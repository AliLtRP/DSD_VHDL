// megafunction wizard: %DisplayPort v13.0%
// GENERATION: XML
// sv_dp.v

// Generated using ACDS version 13.0 152 at 2013.03.30.17:54:00

`timescale 1 ps / 1 ps
module sv_dp (
		input  wire         clk,                     //                clk.clk
		input  wire         reset,                   //              reset.reset
		input  wire [8:0]   tx_mgmt_address,         //            tx_mgmt.address
		input  wire         tx_mgmt_chipselect,      //                   .chipselect
		input  wire         tx_mgmt_read,            //                   .read
		input  wire         tx_mgmt_write,           //                   .write
		input  wire [31:0]  tx_mgmt_writedata,       //                   .writedata
		output wire [31:0]  tx_mgmt_readdata,        //                   .readdata
		output wire         tx_mgmt_waitrequest,     //                   .waitrequest
		output wire         tx_mgmt_irq,             //  tx_mgmt_interrupt.irq
		input  wire         xcvr_mgmt_clk,           //      xcvr_mgmt_clk.clk
		input  wire [1:0]   xcvr_refclk,             //        xcvr_refclk.export
		output wire [3:0]   tx_serial_data,          //     tx_serial_data.export
		input  wire [3:0]   rx_serial_data,          //     rx_serial_data.export
		output wire         tx_reconfig_req,         //        tx_reconfig.export
		input  wire         tx_reconfig_ack,         //                   .export
		input  wire         tx_reconfig_busy,        //                   .export
		output wire [1:0]   tx_link_rate,            //                   .export
		output wire         tx_analog_reconfig_req,  // tx_analog_reconfig.export
		input  wire         tx_analog_reconfig_ack,  //                   .export
		input  wire         tx_analog_reconfig_busy, //                   .export
		output wire [7:0]   tx_vod,                  //                   .export
		output wire [7:0]   tx_emp,                  //                   .export
		output wire         rx_reconfig_req,         //        rx_reconfig.export
		input  wire         rx_reconfig_ack,         //                   .export
		input  wire         rx_reconfig_busy,        //                   .export
		output wire [1:0]   rx_link_rate,            //                   .export
		input  wire [839:0] reconfig_to_xcvr,        //      xcvr_reconfig.export
		output wire [551:0] reconfig_from_xcvr,      //                   .export
		input  wire         tx_vid_clk,              //         tx_vid_clk.clk
		input  wire         tx_vid_v_sync,           //        tx_video_in.export
		input  wire         tx_vid_h_sync,           //                   .export
		input  wire         tx_vid_f,                //                   .export
		input  wire         tx_vid_de,               //                   .export
		input  wire [23:0]  tx_vid_data,             //                   .export
		input  wire         rx_vid_clk,              //         rx_vid_clk.clk
		output wire         rx_vid_sol,              //       rx_video_out.export
		output wire         rx_vid_eol,              //                   .export
		output wire         rx_vid_sof,              //                   .export
		output wire         rx_vid_eof,              //                   .export
		output wire         rx_vid_locked,           //                   .export
		output wire [23:0]  rx_vid_data,             //                   .export
		output wire         rx_vid_valid,            //                   .export
		input  wire         aux_clk,                 //            aux_clk.clk
		input  wire         aux_reset,               //          aux_reset.reset
		input  wire         tx_aux_in,               //             tx_aux.export
		output wire         tx_aux_out,              //                   .export
		output wire         tx_aux_oe,               //                   .export
		input  wire         tx_hpd,                  //                   .export
		input  wire         rx_aux_in,               //             rx_aux.export
		output wire         rx_aux_out,              //                   .export
		output wire         rx_aux_oe,               //                   .export
		output wire         rx_hpd,                  //                   .export
		output wire [7:0]   rx_edid_address,         //            rx_edid.address
		input  wire [7:0]   rx_edid_readdata,        //                   .readdata
		output wire [7:0]   rx_edid_writedata,       //                   .writedata
		output wire         rx_edid_read,            //                   .read
		output wire         rx_edid_write,           //                   .write
		input  wire         rx_edid_waitrequest,     //                   .waitrequest
		output wire [4:0]   rx_lane_count,           //          rx_params.export
		output wire [63:0]  rx_stream_data,          //          rx_stream.export
		output wire [7:0]   rx_stream_ctrl,          //                   .export
		output wire         rx_stream_valid,         //                   .export
		output wire         rx_stream_clk            //                   .export
	);

	altera_dp #(
		.device_family              ("Stratix V"),
		.TX_SUPPORT_SS              (0),
		.TX_SUPPORT_AUDIO           (0),
		.TX_AUDIO_CHANS             (2),
		.TX_VIDEO_BPS               (8),
		.TX_MAX_LINK_RATE           (20),
		.RX_IMAGE_OUT_FORMAT        (1),
		.TX_MAX_LANE_COUNT          (4),
		.TX_POLINV                  (0),
		.TX_SUPPORT_ANALOG_RECONFIG (1),
		.TX_AUX_DEBUG               (0),
		.TX_SCRAMBLER_SEED          (16'b1111111111111111),
		.TX_ODDEVEN_PIXEL           (0),
		.TX_IMPORT_MSA              (0),
		.TX_INTERLACED_VID          (0),
		.TX_SUPPORT_18BPP           (1),
		.TX_SUPPORT_24BPP           (1),
		.TX_SUPPORT_30BPP           (0),
		.TX_SUPPORT_36BPP           (0),
		.TX_SUPPORT_48BPP           (0),
		.TX_SUPPORT_YCBCR422_16BPP  (0),
		.TX_SUPPORT_YCBCR422_20BPP  (0),
		.TX_SUPPORT_YCBCR422_24BPP  (0),
		.TX_SUPPORT_YCBCR422_32BPP  (0),
		.TX_SUPPORT_DP              (1),
		.TX_SUPPORT_AUTOMATED_TEST  (1),
		.TX_SUPPORT_HDCP            (0),
		.RX_ODDEVEN_PIXEL           (0),
		.RX_EXPORT_MSA              (0),
		.RX_VIDEO_BPS               (8),
		.RX_SUPPORT_SS              (0),
		.RX_SUPPORT_MST             (0),
		.RX_MAX_NUM_OF_STREAMS      (1),
		.RX_SUPPORT_AUDIO           (0),
		.RX_AUDIO_CHANS             (2),
		.RX_SUPPORT_HDCP            (0),
		.RX_MAX_LINK_RATE           (20),
		.RX_MAX_LANE_COUNT          (4),
		.RX_POLINV                  (0),
		.RX_SCRAMBLER_SEED          (16'b1111111111111111),
		.RX_SUPPORT_AUTOMATED_TEST  (1),
		.RX_SUPPORT_18BPP           (1),
		.RX_SUPPORT_24BPP           (1),
		.RX_SUPPORT_30BPP           (0),
		.RX_SUPPORT_36BPP           (0),
		.RX_SUPPORT_48BPP           (0),
		.RX_SUPPORT_YCBCR422_16BPP  (0),
		.RX_SUPPORT_YCBCR422_20BPP  (0),
		.RX_SUPPORT_YCBCR422_24BPP  (0),
		.RX_SUPPORT_YCBCR422_32BPP  (0),
		.RX_SUPPORT_DP              (1),
		.RX_AUX_DEBUG               (0),
		.RX_IEEE_OUI                (1),
		.RX_AUX_GPU                 (0)
	) sv_dp_inst (
		.clk                     (clk),                                                                                                                                                                                                   //                clk.clk
		.reset                   (reset),                                                                                                                                                                                                 //              reset.reset
		.tx_mgmt_address         (tx_mgmt_address),                                                                                                                                                                                       //            tx_mgmt.address
		.tx_mgmt_chipselect      (tx_mgmt_chipselect),                                                                                                                                                                                    //                   .chipselect
		.tx_mgmt_read            (tx_mgmt_read),                                                                                                                                                                                          //                   .read
		.tx_mgmt_write           (tx_mgmt_write),                                                                                                                                                                                         //                   .write
		.tx_mgmt_writedata       (tx_mgmt_writedata),                                                                                                                                                                                     //                   .writedata
		.tx_mgmt_readdata        (tx_mgmt_readdata),                                                                                                                                                                                      //                   .readdata
		.tx_mgmt_waitrequest     (tx_mgmt_waitrequest),                                                                                                                                                                                   //                   .waitrequest
		.tx_mgmt_irq             (tx_mgmt_irq),                                                                                                                                                                                           //  tx_mgmt_interrupt.irq
		.xcvr_mgmt_clk           (xcvr_mgmt_clk),                                                                                                                                                                                         //      xcvr_mgmt_clk.clk
		.xcvr_refclk             (xcvr_refclk),                                                                                                                                                                                           //        xcvr_refclk.export
		.tx_serial_data          (tx_serial_data),                                                                                                                                                                                        //     tx_serial_data.export
		.rx_serial_data          (rx_serial_data),                                                                                                                                                                                        //     rx_serial_data.export
		.tx_reconfig_req         (tx_reconfig_req),                                                                                                                                                                                       //        tx_reconfig.export
		.tx_reconfig_ack         (tx_reconfig_ack),                                                                                                                                                                                       //                   .export
		.tx_reconfig_busy        (tx_reconfig_busy),                                                                                                                                                                                      //                   .export
		.tx_link_rate            (tx_link_rate),                                                                                                                                                                                          //                   .export
		.tx_analog_reconfig_req  (tx_analog_reconfig_req),                                                                                                                                                                                // tx_analog_reconfig.export
		.tx_analog_reconfig_ack  (tx_analog_reconfig_ack),                                                                                                                                                                                //                   .export
		.tx_analog_reconfig_busy (tx_analog_reconfig_busy),                                                                                                                                                                               //                   .export
		.tx_vod                  (tx_vod),                                                                                                                                                                                                //                   .export
		.tx_emp                  (tx_emp),                                                                                                                                                                                                //                   .export
		.rx_reconfig_req         (rx_reconfig_req),                                                                                                                                                                                       //        rx_reconfig.export
		.rx_reconfig_ack         (rx_reconfig_ack),                                                                                                                                                                                       //                   .export
		.rx_reconfig_busy        (rx_reconfig_busy),                                                                                                                                                                                      //                   .export
		.rx_link_rate            (rx_link_rate),                                                                                                                                                                                          //                   .export
		.reconfig_to_xcvr        (reconfig_to_xcvr),                                                                                                                                                                                      //      xcvr_reconfig.export
		.reconfig_from_xcvr      (reconfig_from_xcvr),                                                                                                                                                                                    //                   .export
		.tx_vid_clk              (tx_vid_clk),                                                                                                                                                                                            //         tx_vid_clk.clk
		.tx_vid_v_sync           (tx_vid_v_sync),                                                                                                                                                                                         //        tx_video_in.export
		.tx_vid_h_sync           (tx_vid_h_sync),                                                                                                                                                                                         //                   .export
		.tx_vid_f                (tx_vid_f),                                                                                                                                                                                              //                   .export
		.tx_vid_de               (tx_vid_de),                                                                                                                                                                                             //                   .export
		.tx_vid_data             (tx_vid_data),                                                                                                                                                                                           //                   .export
		.rx_vid_clk              (rx_vid_clk),                                                                                                                                                                                            //         rx_vid_clk.clk
		.rx_vid_sol              (rx_vid_sol),                                                                                                                                                                                            //       rx_video_out.export
		.rx_vid_eol              (rx_vid_eol),                                                                                                                                                                                            //                   .export
		.rx_vid_sof              (rx_vid_sof),                                                                                                                                                                                            //                   .export
		.rx_vid_eof              (rx_vid_eof),                                                                                                                                                                                            //                   .export
		.rx_vid_locked           (rx_vid_locked),                                                                                                                                                                                         //                   .export
		.rx_vid_data             (rx_vid_data),                                                                                                                                                                                           //                   .export
		.rx_vid_valid            (rx_vid_valid),                                                                                                                                                                                          //                   .export
		.aux_clk                 (aux_clk),                                                                                                                                                                                               //            aux_clk.clk
		.aux_reset               (aux_reset),                                                                                                                                                                                             //          aux_reset.reset
		.tx_aux_in               (tx_aux_in),                                                                                                                                                                                             //             tx_aux.export
		.tx_aux_out              (tx_aux_out),                                                                                                                                                                                            //                   .export
		.tx_aux_oe               (tx_aux_oe),                                                                                                                                                                                             //                   .export
		.tx_hpd                  (tx_hpd),                                                                                                                                                                                                //                   .export
		.rx_aux_in               (rx_aux_in),                                                                                                                                                                                             //             rx_aux.export
		.rx_aux_out              (rx_aux_out),                                                                                                                                                                                            //                   .export
		.rx_aux_oe               (rx_aux_oe),                                                                                                                                                                                             //                   .export
		.rx_hpd                  (rx_hpd),                                                                                                                                                                                                //                   .export
		.rx_edid_address         (rx_edid_address),                                                                                                                                                                                       //            rx_edid.address
		.rx_edid_readdata        (rx_edid_readdata),                                                                                                                                                                                      //                   .readdata
		.rx_edid_writedata       (rx_edid_writedata),                                                                                                                                                                                     //                   .writedata
		.rx_edid_read            (rx_edid_read),                                                                                                                                                                                          //                   .read
		.rx_edid_write           (rx_edid_write),                                                                                                                                                                                         //                   .write
		.rx_edid_waitrequest     (rx_edid_waitrequest),                                                                                                                                                                                   //                   .waitrequest
		.rx_lane_count           (rx_lane_count),                                                                                                                                                                                         //          rx_params.export
		.rx_stream_data          (rx_stream_data),                                                                                                                                                                                        //          rx_stream.export
		.rx_stream_ctrl          (rx_stream_ctrl),                                                                                                                                                                                        //                   .export
		.rx_stream_valid         (rx_stream_valid),                                                                                                                                                                                       //                   .export
		.rx_stream_clk           (rx_stream_clk),                                                                                                                                                                                         //                   .export
		.rx_mgmt_chipselect      (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx_mgmt_read            (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx_mgmt_write           (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx_mgmt_address         (9'b000000000),                                                                                                                                                                                          //        (terminated)
		.rx_mgmt_writedata       (32'b00000000000000000000000000000000),                                                                                                                                                                  //        (terminated)
		.rx_mgmt_readdata        (),                                                                                                                                                                                                      //        (terminated)
		.rx_mgmt_waitrequest     (),                                                                                                                                                                                                      //        (terminated)
		.rx_mgmt_irq             (),                                                                                                                                                                                                      //        (terminated)
		.rx_vid_st_reset         (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx_vid_st_ready         (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx_vid_st_valid         (),                                                                                                                                                                                                      //        (terminated)
		.rx_vid_st_sop           (),                                                                                                                                                                                                      //        (terminated)
		.rx_vid_st_eop           (),                                                                                                                                                                                                      //        (terminated)
		.rx_vid_st_data          (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_clk             (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx1_vid_sol             (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_eol             (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_sof             (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_eof             (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_locked          (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_data            (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_valid           (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_st_reset        (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx1_vid_st_ready        (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx1_vid_st_valid        (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_st_sop          (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_st_eop          (),                                                                                                                                                                                                      //        (terminated)
		.rx1_vid_st_data         (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_clk             (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx2_vid_sol             (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_eol             (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_sof             (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_eof             (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_locked          (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_data            (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_valid           (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_st_reset        (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx2_vid_st_ready        (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx2_vid_st_valid        (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_st_sop          (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_st_eop          (),                                                                                                                                                                                                      //        (terminated)
		.rx2_vid_st_data         (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_clk             (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx3_vid_sol             (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_eol             (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_sof             (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_eof             (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_locked          (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_data            (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_valid           (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_st_reset        (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx3_vid_st_ready        (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx3_vid_st_valid        (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_st_sop          (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_st_eop          (),                                                                                                                                                                                                      //        (terminated)
		.rx3_vid_st_data         (),                                                                                                                                                                                                      //        (terminated)
		.tx_aux_debug_data       (),                                                                                                                                                                                                      //        (terminated)
		.tx_aux_debug_valid      (),                                                                                                                                                                                                      //        (terminated)
		.tx_aux_debug_sop        (),                                                                                                                                                                                                      //        (terminated)
		.tx_aux_debug_eop        (),                                                                                                                                                                                                      //        (terminated)
		.tx_aux_debug_err        (),                                                                                                                                                                                                      //        (terminated)
		.tx_aux_debug_cha        (),                                                                                                                                                                                                      //        (terminated)
		.rx_aux_debug_data       (),                                                                                                                                                                                                      //        (terminated)
		.rx_aux_debug_valid      (),                                                                                                                                                                                                      //        (terminated)
		.rx_aux_debug_sop        (),                                                                                                                                                                                                      //        (terminated)
		.rx_aux_debug_eop        (),                                                                                                                                                                                                      //        (terminated)
		.rx_aux_debug_err        (),                                                                                                                                                                                                      //        (terminated)
		.rx_aux_debug_cha        (),                                                                                                                                                                                                      //        (terminated)
		.rx1_stream_data         (),                                                                                                                                                                                                      //        (terminated)
		.rx1_stream_ctrl         (),                                                                                                                                                                                                      //        (terminated)
		.rx1_stream_valid        (),                                                                                                                                                                                                      //        (terminated)
		.rx1_stream_clk          (),                                                                                                                                                                                                      //        (terminated)
		.rx2_stream_data         (),                                                                                                                                                                                                      //        (terminated)
		.rx2_stream_ctrl         (),                                                                                                                                                                                                      //        (terminated)
		.rx2_stream_valid        (),                                                                                                                                                                                                      //        (terminated)
		.rx2_stream_clk          (),                                                                                                                                                                                                      //        (terminated)
		.rx3_stream_data         (),                                                                                                                                                                                                      //        (terminated)
		.rx3_stream_ctrl         (),                                                                                                                                                                                                      //        (terminated)
		.rx3_stream_valid        (),                                                                                                                                                                                                      //        (terminated)
		.rx3_stream_clk          (),                                                                                                                                                                                                      //        (terminated)
		.tx_xcvr_clkout          (),                                                                                                                                                                                                      //        (terminated)
		.rx_xcvr_clkout          (),                                                                                                                                                                                                      //        (terminated)
		.tx_msa                  (192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.rx_msa                  (),                                                                                                                                                                                                      //        (terminated)
		.rx1_msa                 (),                                                                                                                                                                                                      //        (terminated)
		.rx2_msa                 (),                                                                                                                                                                                                      //        (terminated)
		.rx3_msa                 (),                                                                                                                                                                                                      //        (terminated)
		.tx_ss_ready             (),                                                                                                                                                                                                      //        (terminated)
		.tx_ss_valid             (1'b0),                                                                                                                                                                                                  //        (terminated)
		.tx_ss_data              (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                 //        (terminated)
		.tx_ss_sop               (1'b0),                                                                                                                                                                                                  //        (terminated)
		.tx_ss_eop               (1'b0),                                                                                                                                                                                                  //        (terminated)
		.rx_ss_valid             (),                                                                                                                                                                                                      //        (terminated)
		.rx_ss_data              (),                                                                                                                                                                                                      //        (terminated)
		.rx_ss_sop               (),                                                                                                                                                                                                      //        (terminated)
		.rx_ss_eop               (),                                                                                                                                                                                                      //        (terminated)
		.rx1_ss_valid            (),                                                                                                                                                                                                      //        (terminated)
		.rx1_ss_data             (),                                                                                                                                                                                                      //        (terminated)
		.rx1_ss_sop              (),                                                                                                                                                                                                      //        (terminated)
		.rx1_ss_eop              (),                                                                                                                                                                                                      //        (terminated)
		.rx2_ss_valid            (),                                                                                                                                                                                                      //        (terminated)
		.rx2_ss_data             (),                                                                                                                                                                                                      //        (terminated)
		.rx2_ss_sop              (),                                                                                                                                                                                                      //        (terminated)
		.rx2_ss_eop              (),                                                                                                                                                                                                      //        (terminated)
		.rx3_ss_valid            (),                                                                                                                                                                                                      //        (terminated)
		.rx3_ss_data             (),                                                                                                                                                                                                      //        (terminated)
		.rx3_ss_sop              (),                                                                                                                                                                                                      //        (terminated)
		.rx3_ss_eop              (),                                                                                                                                                                                                      //        (terminated)
		.tx_audio_clk            (1'b0),                                                                                                                                                                                                  //        (terminated)
		.tx_audio_valid          (1'b0),                                                                                                                                                                                                  //        (terminated)
		.tx_audio_mute           (1'b0),                                                                                                                                                                                                  //        (terminated)
		.tx_audio_lpcm_data      (64'b0000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                  //        (terminated)
		.rx_audio_valid          (),                                                                                                                                                                                                      //        (terminated)
		.rx_audio_mute           (),                                                                                                                                                                                                      //        (terminated)
		.rx_audio_infoframe      (),                                                                                                                                                                                                      //        (terminated)
		.rx_audio_lpcm_data      (),                                                                                                                                                                                                      //        (terminated)
		.rx1_audio_valid         (),                                                                                                                                                                                                      //        (terminated)
		.rx1_audio_mute          (),                                                                                                                                                                                                      //        (terminated)
		.rx1_audio_infoframe     (),                                                                                                                                                                                                      //        (terminated)
		.rx1_audio_lpcm_data     (),                                                                                                                                                                                                      //        (terminated)
		.rx2_audio_valid         (),                                                                                                                                                                                                      //        (terminated)
		.rx2_audio_mute          (),                                                                                                                                                                                                      //        (terminated)
		.rx2_audio_infoframe     (),                                                                                                                                                                                                      //        (terminated)
		.rx2_audio_lpcm_data     (),                                                                                                                                                                                                      //        (terminated)
		.rx3_audio_valid         (),                                                                                                                                                                                                      //        (terminated)
		.rx3_audio_mute          (),                                                                                                                                                                                                      //        (terminated)
		.rx3_audio_infoframe     (),                                                                                                                                                                                                      //        (terminated)
		.rx3_audio_lpcm_data     (),                                                                                                                                                                                                      //        (terminated)
		.tx_hdcp_akeys_dat       (56'b00000000000000000000000000000000000000000000000000000000),                                                                                                                                          //        (terminated)
		.tx_hdcp_akeys_ksv       (40'b0000000000000000000000000000000000000000),                                                                                                                                                          //        (terminated)
		.tx_hdcp_akeys_sel       (),                                                                                                                                                                                                      //        (terminated)
		.rx_hdcp_bkeys_dat       (56'b00000000000000000000000000000000000000000000000000000000),                                                                                                                                          //        (terminated)
		.rx_hdcp_bkeys_ksv       (40'b0000000000000000000000000000000000000000),                                                                                                                                                          //        (terminated)
		.rx_hdcp_bkeys_sel       ()                                                                                                                                                                                                       //        (terminated)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2013 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_dp" version="13.0" >
// Retrieval info: 	<generic name="device_family" value="Stratix V" />
// Retrieval info: 	<generic name="TX_SUPPORT_SS" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_AUDIO" value="0" />
// Retrieval info: 	<generic name="TX_AUDIO_CHANS" value="2" />
// Retrieval info: 	<generic name="TX_VIDEO_BPS" value="8" />
// Retrieval info: 	<generic name="TX_MAX_LINK_RATE" value="20" />
// Retrieval info: 	<generic name="RX_IMAGE_OUT_FORMAT" value="1" />
// Retrieval info: 	<generic name="TX_MAX_LANE_COUNT" value="4" />
// Retrieval info: 	<generic name="TX_POLINV" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_ANALOG_RECONFIG" value="1" />
// Retrieval info: 	<generic name="TX_AUX_DEBUG" value="0" />
// Retrieval info: 	<generic name="TX_SCRAMBLER_SEED" value="65535" />
// Retrieval info: 	<generic name="TX_ODDEVEN_PIXEL" value="0" />
// Retrieval info: 	<generic name="TX_IMPORT_MSA" value="0" />
// Retrieval info: 	<generic name="TX_INTERLACED_VID" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_18BPP" value="1" />
// Retrieval info: 	<generic name="TX_SUPPORT_24BPP" value="1" />
// Retrieval info: 	<generic name="TX_SUPPORT_30BPP" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_36BPP" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_48BPP" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_YCBCR422_16BPP" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_YCBCR422_20BPP" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_YCBCR422_24BPP" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_YCBCR422_32BPP" value="0" />
// Retrieval info: 	<generic name="TX_SUPPORT_DP" value="1" />
// Retrieval info: 	<generic name="TX_SUPPORT_AUTOMATED_TEST" value="1" />
// Retrieval info: 	<generic name="TX_SUPPORT_HDCP" value="0" />
// Retrieval info: 	<generic name="RX_ODDEVEN_PIXEL" value="0" />
// Retrieval info: 	<generic name="RX_EXPORT_MSA" value="0" />
// Retrieval info: 	<generic name="RX_VIDEO_BPS" value="8" />
// Retrieval info: 	<generic name="RX_SUPPORT_SS" value="0" />
// Retrieval info: 	<generic name="RX_SUPPORT_MST" value="0" />
// Retrieval info: 	<generic name="RX_MAX_NUM_OF_STREAMS" value="1" />
// Retrieval info: 	<generic name="RX_SUPPORT_AUDIO" value="0" />
// Retrieval info: 	<generic name="RX_AUDIO_CHANS" value="2" />
// Retrieval info: 	<generic name="RX_SUPPORT_HDCP" value="0" />
// Retrieval info: 	<generic name="RX_MAX_LINK_RATE" value="20" />
// Retrieval info: 	<generic name="RX_MAX_LANE_COUNT" value="4" />
// Retrieval info: 	<generic name="RX_POLINV" value="0" />
// Retrieval info: 	<generic name="RX_SCRAMBLER_SEED" value="65535" />
// Retrieval info: 	<generic name="RX_SUPPORT_AUTOMATED_TEST" value="1" />
// Retrieval info: 	<generic name="RX_SUPPORT_18BPP" value="1" />
// Retrieval info: 	<generic name="RX_SUPPORT_24BPP" value="1" />
// Retrieval info: 	<generic name="RX_SUPPORT_30BPP" value="0" />
// Retrieval info: 	<generic name="RX_SUPPORT_36BPP" value="0" />
// Retrieval info: 	<generic name="RX_SUPPORT_48BPP" value="0" />
// Retrieval info: 	<generic name="RX_SUPPORT_YCBCR422_16BPP" value="0" />
// Retrieval info: 	<generic name="RX_SUPPORT_YCBCR422_20BPP" value="0" />
// Retrieval info: 	<generic name="RX_SUPPORT_YCBCR422_24BPP" value="0" />
// Retrieval info: 	<generic name="RX_SUPPORT_YCBCR422_32BPP" value="0" />
// Retrieval info: 	<generic name="RX_SUPPORT_DP" value="1" />
// Retrieval info: 	<generic name="RX_AUX_DEBUG" value="0" />
// Retrieval info: 	<generic name="RX_IEEE_OUI" value="1" />
// Retrieval info: 	<generic name="RX_AUX_GPU" value="0" />
// Retrieval info: 	<generic name="AUTO_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_XCVR_MGMT_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_TX_VID_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX_VID_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX1_VID_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX2_VID_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX3_VID_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_AUX_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_TX_AUDIO_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: </instance>
// IPFS_FILES : sv_dp.vo
// RELATED_FILES: sv_dp.v, altera_dp.v, altera_dp_phy_rx.v, altera_dp_phy_tx.v, altera_dp_reset_delay.v, altera_dp_status_sync.v, bitec_dp.v, bitec_dp_autotest_crc.v, bitec_dp_clock_crossing.v, bitec_dp_cntrl_sym_scrambler.v, bitec_dp_is_gen.v, bitec_dp_mac.v, bitec_dp_prbs7.v, bitec_dp_reset_sync.v, bitec_dp_scramble_16.v, bitec_dp_rx_8b10b_decode.v, bitec_dp_rx_aux_ctrl_sink.v, bitec_dp_rx_aux_sink.v, bitec_dp_rx_cc_fifo_mc.v, bitec_dp_rx_decoder.v, bitec_dp_rx_decode_msa_16.v, bitec_dp_rx_decode_vid_16.v, bitec_dp_rx_deskew.v, bitec_dp_rx_dp2st16.v, bitec_dp_rx_dpcd_regs.v, bitec_dp_rx_dpcd_regs_link_services.v, bitec_dp_rx_edid_memory_16.v, bitec_dp_rx_gear16_2_bpp.v, bitec_dp_rx_gxb_cont_16.v, bitec_dp_rx_hdcp.v, bitec_dp_rx_hpd_ctrl.v, bitec_dp_rx_mst_sink.v, bitec_dp_rx_pixel_fifo_double_16.v, bitec_dp_rx_pixel_fifo_quad_16.v, bitec_dp_rx_pixel_fifo_single_16.v, bitec_dp_rx_pixel_steer.v, bitec_dp_rx_stream_sink.v, bitec_dp_rx_sync_status.v, bitec_dp_rx_training_10.v, bitec_dp_rx_ss_align.v, bitec_dp_rx_ss_audio.v, bitec_dp_rx_ss_decode.v, bitec_dp_rx_ss_depacket.v, bitec_dp_ss_audio_fifo.v, bitec_dp_tx_8b10b_encode.v, bitec_dp_tx_aux_bit_ctrl.v, bitec_dp_tx_aux_fsm.v, bitec_dp_tx_aux_source.v, bitec_dp_tx_blank_start_gen.v, bitec_dp_tx_bs_bs2dp.v, bitec_dp_tx_data_fifo_throttle.v, bitec_dp_tx_encoder.v, bitec_dp_tx_encode_msa.v, bitec_dp_tx_gen_vid.v, bitec_dp_tx_gen_xport_clk_divider.v, bitec_dp_tx_gxb_cont_16.v, bitec_dp_tx_hdcp.v, bitec_dp_tx_hpd_monitor.v, bitec_dp_tx_idle_gen.v, bitec_dp_tx_measure_refclk.v, bitec_dp_tx_measure_vid.v, bitec_dp_tx_pixel_2_16.v, bitec_dp_tx_pixel_2_word_fifo_16.v, bitec_dp_tx_pixel_packetizer.v, bitec_dp_tx_pixel_steer.v, bitec_dp_tx_pix_data_fifo.v, bitec_dp_tx_skew.v, bitec_dp_tx_vd2dp_fifo.v, bitec_dp_tx_vsync_gen.v, bitec_dp_tx_ss_audio.v, bitec_dp_tx_ss_audio_fifo.v, bitec_dp_tx_ss_audio_mux.v, bitec_dp_tx_ss_de_gen.v, bitec_dp_tx_ss_encode.v, bitec_dp_tx_ss_enpacket.v, bitec_dp_tx_ss_mux.v, bitec_dp_tx_ss_rs.v, bitec_dp_tx_ss_steer.v, bitec_dp_tx_ss_wop_sr.v, bitec_dp_tx_ss_xport_clk_divider.v, altera_dp_phy_rx_native_sv.v, altera_dp_phy_tx_native_sv.v, altera_xcvr_functions.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, alt_xcvr_resync.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_native_sv_functions_h.sv, altera_xcvr_native_sv.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v
