// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nA8Y5xdJO3fbVCxszJDGJF85SDbNGf+riKGEM7WcNAMYvd7yUH4s8NGRO77TuaNh
mo3ig9UCeheEn3W/SoLHoiYfrXVf4TUJCyn1oaN/qwaHzgdeOsYdgZ3SMr+niWBY
veh3DctPnyY+KVA1K2Ga8AyZ6zlon2NWJIDBFNYKr30=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7488)
2ao1o9em1Iaa+YZLiuuEQC9LeANuyGMqBKN7y+iJHGh91H/BSI8RJNV2B+HOZtpz
XLx0FZuz9SV6WXA8WAH71tsfU5jySOgqqYwv14C/rEPvZ/TMEgmAfQRXWQj1gN30
JFQS/Skdpwqy8lMUorQCfnv4LNq4TInNScFNO10VwegVJ67nJWAYcd/0FEvr7hoM
jLJIzXsedVAHgNMkt5gLKbnL2bwkHogyuIUm3CsJWlgI1zCEeO4whVCOk+vVyLjA
B7zo3pP53XJMDJYHawXZNE0NjBUJmavD2tETVfU3gjb9Ji1Ek8w6n8zAuI78ixB9
Acqep4L+zsnvnBDHjqXb13H+Kv04oMGktkxRZyzaLAC8Jn6kBIMpw9KZBoYDD6pv
Qsoqat8egk1hLBujUzUP+WurdFLVfZEZWNa0X6rzjKWG/ZsCZGzZawKZVkSA1ulH
p96fYnI6lYZb1dWZdeu8+UmS0+yTvvQ04D4uSHPL9JMFSYlZ6QAHxEQ90qhUO19k
Y0E/iZFES9foSAHidnn1tqhb65xRw5NRww/jONoBcf07DwUWJaaza93niFsv9H9o
YEezPMJBWuqZQx5pORyedIEQFdnEDmYfw5hpRbBubb0s+ggmBtEgoot6vUilwaVZ
ZDTzW4P+8j7I0o4SbIWernEWL+8W2SdXsj+rnvwQSnsMYWR923faC/ZWW+ZjxVqT
GmnP4vA+B8E0w2GDSwXjs1dRNUpD0wp15IiAC35CyjurnfyJ54UlDzbz6G9lH57+
Pc0A1CBEOR9z5degw5i/eUUjwnT94sxcLrLfd1Rd79ZFJo1GO6qW7fRTGYfTxhon
85CH54hvtLfaG+I9YGAaOuYd5YGenRcXBZshiizFqvyqiEhPSjFUUZ8/xLU1uf9Q
C9bcSbFz8N5cgt/BQxeTrEmddJ9bI9dPvbegzQRexK4LouycXutUMa35p9wArbU3
NK4kxF/ZbMoyrA+p881K5j7LpWKjRRcUt0u65EJsAOVdnrslkbcQ3+8u4wKMSb4P
5DjUP4xgBeAyzZk5y92s/H2TTO6AukeCwfMoIeMDllQGEh4TiDrbmAIc3OE4dwG2
CZr6msOdzQijN32ThOEKKYIGbzS5PElkiocWoVaHtVJ+1CU/Ai4TIR5TqK7ZrpgH
gsf1YsHkRKpczMsUW6oN5hE5ooPKjVo/e+6ivy9jGd5KaC+Ardh9lwGz0lxrLrmM
1bWwYV14BnKomTQe3JwgWqQ4KpD0QOCduIGwG46/SovOmeqIKb9F8JCKtBt3ufHK
bYqgfExZIBYS527ogccivmHjLD1+Z2xCmBpfdjRnvnb4IBsUfCGAIvNAn1ax2wOE
67TrRNcyvyENHA0YcpJVCf3jgXpmcyhOGPBgzWNZmVrDLB6CAqZR4tL1E4Rk0aXa
wRR/LPm0XbX2vxw2zrpJoj+cWtsRgU9Dw3FSd89xQ5hVGbSiuOR+AdO3GM+qELqn
YEKB6gIbX+gFcV2h6UG3CllavocWN9guhehSmcudlixbt9tgRNQqWbVmkUmViGpC
qLV6K0ef3wonjnuJG3t8bT6PxsPUbtAhxNXaNGMF8obQPsVSB333yGnYv1/3SGMK
dInjapEnfasOB/SB2pVRBmmk+uO07JZO3OSVQxurrp6tW7+6stkiQBtkWdHm1RLk
bjURWlaM7Y5TRmHALZvgbNRgvJy5qkDkXblqw3Q4W1xxlVIhYmE/3j6tA65BStor
cdGEiCD2MnJF+IgZ7V3bbrixmy0+0z517QPfeqDLw3BSgcJWpBv4YF5/hFH8YFxO
UFczDjEV4zUiR58cVHdA3kqmNs/soS2BQWA1rZyY4EAS3uecvdQoM9nDimSeJmLC
EV7IB4bALnVEuJRMz0qjMvahYm9u3ieNZIVmAvBB52AqcPdIoSVz9yUSqtk/Thf6
IiS6LyFPxk9ygsPq+Q2bY9c6kKCEY0nnVf4QYmEagMF5qYCsgg1znLk6V0ZdxJJS
1FdgINUBgHdzPjmbi/kr61X8wa+kxHeuqB7v0iFlxmVVfyqEUaQ5hX+rFE4oABnO
ZnUZk+0uwS4Ckf0tD1hWXqiW6nZ82i5Uj4+Gw1WcFdYoHmVv/7eaG3VDhbt04VRe
2u6pZCKhe2yvaNUSWfjiumuoap41+LNnmJYtRHqWOQLdphMwG2CcgoJVwa7ZLGB8
Nb0/7j7uy8fB84gIwTgqXNPgsh/lOWiHnKH4XlahP8e8UPcezMkglJMtuOz4QePb
mz6PT0KZUP5W697SXe0DPO31e0r8iryW2epUWdSox5rI6plQEPKdiqRix6Ta3Dh5
6/o8faEWtIX2f5TNJBfmHkr3Yw5ueMZ7eiZLtcCc1Upd/ve9RnmFE3aVBfc+z36O
Q2+sEsz3xwW7yr7tjWGNNO01jLLE5dVZS7qdPmqAlETbp6zL145+SquJ2qXmjnkJ
xM1zXzdUz8WOcv0st756Fuw22oBWZ7hiFsx8GqgnImINS3UdUwdLrc/QCJjjLAq+
6j+dRiHZQF2QUZDwUWLLn+tLl8wtSg9tUn0Ni1oEqEUvkiBWco4eYyKk4lDsR3tz
++sF+Wb+gJKGWl0LTf0oOEfk13pohlYru31vYk5TRiaBDi1ZeId2dPOO7pRjon97
4Vgo+eQDTrpfQfuHD0/jKYTK3aHgzZh3Nm3RZMnn/fCUdOgyVRfq1XxIRvB4qA9C
yijCcLhvJsS3orJIL1B4n79jY6Pa3I7mRIKSZVJdoNr2WKGMWdU/9f1PQQRQ4qUJ
l81++R+KIHO09F06WyifzdEvjtKh4qYc515C1OtVPxjzBfbttd88XQGLDqScmCSf
ZjJ0NXmxgkEC0N5Dqc6ANan6PrIw3sOUZLwOOK3KJmJ9x1hC6yzXfiEa9KCB+a/d
KgDuOaNuo3VfK3wu66PACBWAMTZ++ENUJsAf56CyfNPXWwZ7NEuIHRc7P2nFGPEw
JfMIncN5IdOCMjwKJE5bpMnVSaPM/ZHwhMgTXRt9gnGn1vOHUuQUlnnDD7LSAWk8
0NH6lA+t4Ka6lHieXkqghF1JmCvgnS4xudWAX3FZZ1efA3fSsr+ehbidOkMjFDid
P5l8IBqZQBTeBS0Q6pXbUVpjrcU6ZBsvEWWF6u4Mg6YxW2Vqznfd+lxXImchXSSr
gxfBdosPIDrZEQXgUesYMKemj7XPAQ58+L6kH69pQ3rIsnSQRug7Yl/h3PwNLHdi
1VOIvIc1g6X9dHRWOCaku958CSRZNgGTXLVr8ET5WR35d+aAp5aeqN7pjcsooU3h
dM7VbowgLoHHAzUexc2T9Hh/053a5FtdiJoeqTHv3l9OdpUs/F5k/ov03EYoAIxK
35tE3qKbUk3SmBbh7u1COkoZjIi2oM/Ib7OlPPLxFD3oTb99w0kuP1N3xSMTDGQW
3CriA6x3qZq9GoOJVsyneMPMZnmhjyifbDrmMzOZL86mu4kFQjCFR4YnxAFK1aGp
Sb7SIFPj3IcGYGzdOrJEalVQ3MTz3MMo6aDYkhv342TSgn+Z7Qq30ELG0Pdvbt5A
6pqF5cM21rhazY+WDTzp8prSfitPrwJOC2iI+Q3QmODiQTmAet7yEt1jZgWqQXNH
p8jJ6tsvUnH1EJBm3Dr+cTH1z+qFTeAlIX0+xjVc+G2sB4y3tHktooZD6H4P1Dp4
Z7Uda+h/+mkmoF7sdILhnaI1HFQB9G2MvQsWTbK9AUCxdjKo9yq151H1srhtxJXy
1mBLjPliMuY4QaMi1IB9+1SHC4oEh3ivzClW9bQBA3zhqgJ0MA4Ii0WMGe9NMWFm
LIgyuZ/zWOhFOv3AouJQE4/YQY940IEaH6OHTNneZhnuZrzxeAHtYAuPIXYm3C9E
6PwBzZKH0m5g/ILnRICix5rxJ/oC1vQ5JLdBGdZWDyRD43Hd8uxy0md+YBgFMxA/
NsUchyoc85roH9hg8pYvGHzZmsez5Z/NWzfjyamUgM7Hmo0BbNCV8rIgkz3rMwGc
1YXC0/buis1EijOUo5ZfotWmjXr9Y9ySlC+GrI0NClAC+QZBBg0MyedOMmcauC28
wnnQjxD6hNAvm6jW28/h6s4VYYO1LLTcI//ewninMOJ6jn47K/3tkvQ5kYjhxab4
be94s2wQL8BJXrlO7+lU7i6GiD1H1AArsAuZOq3FCnlW6xuwxkPlt7XM1BVFlWVa
UB94Okcu9BKoFk4mJnrK7MFaKv0f8zgdB7qVvZ9yM+/z/Qzppblq9syBLOx+kMxU
Nh5tyC1tS1LWUrH5lj781oaLmgrQnerGxCY7bBlyosThWa0Zbmb4teG/0Z/HbwZH
jQDT3JQlQ+UkOVVTxpsPkybqm25LAbrUqhTDCf/3RL0vvdMHB++kh4mtv2gn/bO1
NEzkIakL88n7D6m6oh37bfNOJArC/EA6tdUMlIqed9u/TnGu3zrj5kJ3AAozLpXz
ZPetU8SGiIrNHeGJfhRMmj02tk4ejmDeHLeRuMzOOnkBle4g8V98NfRQ9EARcQoF
SLQOjiByS8qRMZAJZAD8nsTSk+oa3ReQI9NCF7v9z4+wi5lxmWgQ69GIVRZM21K1
4ou7RN33gGWQVc4UrDL94nvMbVR6Z+bSNRt7FAiOrbT/PCabQgS/wp3qN8MTfXpq
LUI/ANAVwyay2ZW0/ZDTS8pBgD4ZlvTZcJE2pMUPd8ryZtECnn88Cp0OcTApELIu
yquqL3be64IpdBG05CPop6Dte+XHc2W0qLqe0IARfDwSKS5/P+0n1LxcNoJQMZe4
wWo3ayGPcxLWQCoRxC10m/PdQxlYrgdfjAQlk+NotXqqKC/ax1MJjHWuX/4ZyWkr
3E9tRdsbSCyApFS+km5GpqiZJuiVf2ENcCYfihc8vpljY15+O3fbSP94qTe3PeSV
Vx+jYq89I/3ftI4PvdmvtBG+hdO22E44If0W4IJnwBjEOOc7h+aRk5wBE1Qu90dY
6XcT2bboiGIHXVjdIGXu/NHfuRhrSZkJYsd7gUeUi92vFx0CDSA6+T5O01WU/ur+
9Grggbwn/piuqFc2EsLD66+rLsSH5ClpyVDhRd+kHAWVpJPoWaW0qbmk8ybMILaA
qFO6LEIZcbzSuokvJYW2MT88BGotMrPZhfGdrc1zIJrkxEUsQAXYBwHnrCm69yv/
YjC65CsE6nHJB29QzfHH8ZAKGToLWVcJ2JoK7OOzzJxOshGpDHrlEV63B4U56jqv
axyqbdFI3iNa08cLYsBpArZsMC+DzmUWRm9Ie3HtQgbsQmTstk2MIJhrG4P1lsJL
Um/f9j2MrNM/GTnnjs2WRHsz1bmMHCuGyczpiQhI0qG2PHC824YYfMvPc2rOQop6
tm22NovtTy3EgpAGj4mT/5Pjx2KGIo28UQ43Zne7HkRgeHqhdtmbyhKGJ4ie+CFX
QPls2vrvYrnmZHstnSmeXKTXdQrKTNY4ELk94TVP/VdYTLs+6Wf01dmkeX7DGFB3
z09fU7qAYfwHkRfbCcOpyknQyI+WRr4DsmN83e723g6/bofKFYzWWWEW3DeIVWfr
h5bFO7zlXn6vss29/k5F6lvTLV+O37aMl641q0Spw1OuKjRiKENixHZPvlpGB66E
nhqaJGjlEMwMgPzq8fic9wGMcXHRDVeXCMAWuYlg/IuEhG0h6IOPPqW/6nW/3IfT
/+uFx8sKUyF2LCY9Dr/Ay00ZNEj73KNga1qUobcod0ZDJUWYE3mLbRpxu5yM8FQm
IJj5srTAMVUXbVKi/zSQokwyn8CsSmnSMspFKzOKkP1dkr139wY/EvJDnk8wUPzR
em+LaeFZSZUzML4qWQYaW67yE8ZCaEVfFmGri5ziCmTpfBNeFchX43yAtGUHwYeg
gnTbjgoPaY7XT5OyrizxMBm47/zBhgZqf6Kp3D3dGJV1n0l6uS+GLl4BVfVBsbMs
U7yE8Py9RctBA/rhqSmBOmvWxCQbvN/7WxvKX7XfpDI7gx0z1hsomgCxWxhoqBkW
7jnQYQd2HNF6wkqrwbW8gPVr1hv107/HiRdOozQS4VjkyZ/Y7C+A7NTsjlI8PDaM
YtmwDyaQp0WYP69bgj/k9HsR28qJadnyP/3aEIdT2FXHrNjsDpYvlCb79D9v0jnc
zoaGH5+kJqrX3szqhXtt2cZcbDCCXae6XqCveSTPKYmXVJeijNx7egE/7mPhEM4U
6F8HGf+it1vTiDQiompNo8SyCRJh45baER/Ujtd2YwSHwD9zkqDHwi2HkdCzbrdV
H0EPegUemnj5SVMuqaQIPhZF0orSbpDhJK9qCIShrdChnL8v11/3TrIQ8S+Zeq6k
+UqoYIA60u2atD4y+869RPWf394Hb0d61/TsHQHL/odLu+n/8nCk9iUrTR+Ed5vF
46O81S8Ej+ZYrvVph2t235HIirg1DAs0Kq6E4ZcxpDXpvXH/sJhW51xER2OuXnlg
so/EFBZ66JXiir1weClhtZTijp0s45cuG77niiCtSNw4ulLMpVRcA6YhYRKUSCW7
PdM0BafVXA3o+UXTHv6fcwWKLDf5nDIwvYVUdWOemrIxcIaJ+P8CXDpW+02OdMdI
tI3+2f84/vyI3LQAgro5x0aZTln9jOxrjiFm47L9lxxuw0L99EjHH39y9uwOcL+S
umeOUTlpq/RpMQmgrm0JrF+WvhlqWObaVicWBLS0e8tN6p0f75rmJ6rRf6mnIeEF
LoJPK05EdEXBV6ERyTvU3My+BSk/pCANE9CJlQhLMu6lzQGozWCRdb8p8n03z0Pe
9x5wjNlcruno75SruvsmqeEZ72K+D0nCpqZI1I7zeY2SwgDxhBNB4SZLtGllmokZ
lx+d8ksS644dYQ71q6wqYb+PRm9c3ek8hIkPjoXHxnwKZYDgsQNW+bt9N357+q1c
uxQvkva8RoAr36wk1gD5jXbEC1Oh41lBu9XbaluAi/hReaDBbqjv1AMyIkX2OGW3
8FgIVNcb10yH8Nu/E6Rayb/kZ8/abBuQKdfovZ18d+8TcjGFif7Jvl4/jPriLYJP
SY90jdCv7vINZMpurV7Tq0Zotc33MnFKC/zn1FZD/+bFRK8bf9qaIEq2evSTiQQ+
aGWIkU8i2iQ+xrzaGuJ20yjYch5pxvBOXUbyVKjLHBo0cDDqMyX54oWkyKYrBGJR
EzBgryQ/L4XpId2O6rYZrzKm0uXAhTrYi3FaFURaXlfvLMLxc5QYRuUPZYDRmnaR
bFqWZjmT0Otspte19PapRoumMtH7ofZ77ci0yOICuGwrsxDIZzIRQY0lQ5yLOD2B
o6mJLl8KSrOg3KdaxykBqA9YSM6qicfY/hiVHR8Mmv/gtYAS/mHHezAEAAnbfmmO
HPpy8kUKzAfMGEDkU1WzQl/C+2QAXd/BYo+IVTKxR/Xa0siIVV3XyS2QlTn7k5Ta
5z0iu2IHsjTBxH6ieg0R8usxQE0gFtCZdiGt7pXzru4NXjagRPh/JIV0GqZVFUvF
N0dc6mX93aAp2gj+HHykfDijkm43eQ0GP1p6v6mTPzvhjWsu/n/wHnY2jmrrZHNV
CZt8FWYO+w61G7eEIPFAAIRY8pnIcTi5ZLsuzyqdXmNXg0xWP4NKbREOw+XWDLEq
P3qW+SB7cQnUST6B427intGRlMFB+BinlrF8MYd2b59fFUJalEIi5thln2tLySsu
hVDPbkOO8LG908PXmOWdtXKY29vU1Pyr+jc2T/Y85o517TX6NpM9eq5X8slGlLwB
b3QdjLRnG01rSmynC8wXOZKxHJfHzy9j+GbwY9pVcHjO09jEe6fZmLzmEHpjj1JD
BXCzlhRqUNhfknlVs7Wxy2LR8JR+BEk6H5X9fg0alDlw0JpQKaqXRwrlTSm4tcMa
odO+tzfVgilspIFmkdVk/Mj6K6HPnTB44p5NmgKxhIXRp69SON7NnSQdQL864vGH
fg4u4ZeSYdGq8NyJDrMpdu0U/0KVqtvZkHzik63ZW+VahkBKhZy0eDlvspH1mZuD
IXnU4BvXmNciIlLmO0h2x9C3qDtNNLUlxvn5pXRHjCzE0gGYUkKyeJcXgoqJNzO4
Ff0AApmUEYQgZ5Q0Q7ZEA8KVB5gcPaRH1SwAHfoyQTirLCIPkUmU11Z/NZS6dA4S
R2hNFj6xpbE7xjg3vTCiGwvXFU8OtwJ9jkZvhsUmrdTEg47q3LH+l2p7nrupBUiu
sCioJxl+rp+1jZKWVaLxA3i55ccd1zw6/eE6rVmYoWK3mkALgKBuNg6QlziEL+tM
tTRVuteEhbEg9DLrTE/uWHAjlZHm10nDp7lYqXoxOaTW4Mk8I6UZjxsprGFSIJAB
qhuwGcIbbjQBDjWJ/YgkNVR/URSKMYKNqXkpODdS7WBSZroJXpxaynpydgK0qFSm
gsBFhCB/L9mj5lb6uQF0m0hWOd8vH6t+0Ld7rbI5mrmJaP2octKXGSMm/ls19B7P
D1Be5PicVLv3z0gdRZVdnXLaRKR2PSyXmfwT0MXfvzKubJcLE5wkk19pwbaXyXp8
QquCTaxlgtXGVoTclbfw5EMcXtgFjP//CWQg/sOhLxfbwhm8KGfgEm44r/qnPq+Z
MXERga8+QhnsPHuz8vH2lg5UM8m9zrwMRhxlsjFGKPtfrbG1rS3nY50Ld3IrABaO
1TGKpkqLWHQeeZk3nV9sYsJDyn9f6xIq6L5d9jxy7RRntnSRl13zhQCqsLlHph42
7YncW2wE03sCEBm7y602EUMtowMinPXW8YJOAtIFs5n7b5OpQ9XHdi2gkjWp1gPQ
PLONQooYCONn+K/gErkOGTkusdVVjoe9r2uJ9l4r24QCRckofo62bttfJevV7X4Y
o2VebimXq89TzEIsC6RJizVEvCKfWeWS2lgKHZUZlRDnTQPiPwcwYfa3gzDIq0YT
FswT/YkcEKrpZdgIPDiu681DwiZXxQ8Hlwfg2JiHw4/5MMobODAR9d5XlLq7GYxa
9HajWa5Bh/trihcykX+BkTcbvvPesH+5RVJR0H7uChlY6AhEgOWTVt7C3AQbw6PT
l1+hLFy46sRAfpiu9rq7fo10gUW6cGzg8m6Y/eeveaBLIsdQi/OBTrzzMtsrbw36
2gRVAExwT0IDyfLiSHhUg0NAqqtwx2/x87IfQu4Zimi6lJPM3iDaCP7S31nFp7/T
3bBktePhEo3Em3ZTQsUQCFBNi6sDminKLyLyris7mJzCcEdBVaiq+AjaJUUxeuIS
BgjmQ6482qi5rgXVETYqk0WjegfMr8RNE5925W9osm9j09WHQenyV+5BN5HO1Q6Z
AHm9XIklumlGlFlfgXvqwnF2a04ZB9TqBAfycpAerfzMHZ9f6WJqwymWZ4xP08pw
Ev33ufVFvD3GjFG6ucJbnK0wkog9/rsRMRSU0EWZ2SF+Ibh5mTkM96fS+sYaBqly
ksDR7tGrTTfPiiz60hrXJtmsm3WC45QlnnTlFvk2vopA0xny1yZj5xeM2AGK1fYL
40Zn1gXx2vI9hHEZTUNwZtmSgwrKFh56wWlwsWqILKqGBuv2ELYvqz/xoVFvQUER
s4ed/Oh5puTT0FKssERsi6NG57p4mRfibjaAEJbjHtVD9Bz0gC7OnA8rv16AfiVI
W07o4T9kvnZbDI8gbTebNsTz8P9+0A54U98UvSudqSIZUvwYWhdwZRBFhctNiYpU
I3h2WpmOdXz4oJhfcW9BuJgKIaHC16gFTeP+Cu00HjOjXZICvbf1NFBNQPKf01C7
r+vPEyyKA1rtxLGvBhLRZDzajbi6SV5gV++FMwu7HorlkXhdsGF/d2WJVU9yyTxF
PbETmgfAsdOqSAR5S7jq4c4uLMLMhDo7wthgq9Sh6FOuBC7S0Dqzw6fvcTPLglY/
2Cu0/62klrn3gZB2eLRMwh1sm9Eo/SdIyEHh5FDIYAhJqj4UpCd3Kqsr5MtHv8bd
Xi/F0MHQmZXHlryJr2QsYLP10xiZ50LsmrfZryLnqF6QZtF722oeUxA+GkXuvU7L
EuD7c60So0J/hjErTIrsGThxZgwpCN87dLJ3ahgEh8AdndSpO1eUgIX4Qir/GRqG
`pragma protect end_protected
