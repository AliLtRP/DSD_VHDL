// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rt/eK/KdPkn4GIYSVYaC/PKqWKQe6V7rTDb3mxNfTxUNn0TskraRM5RIyaJgA93F
aCc8/kwyAnLrD1SwvUSlnMyMaSUWhJb4Tb82XNmzELSGZYgBqQKqMNIYgMYoytod
FTbghXZjnYqprNuhewaQBfHOdenQu2R+ImMw8WScRbc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63984)
JO3bGyIg4TueqDUSxxcX37f07GZT0wIukkCGWXV5dIgEb2kilWbJMnoG8dixBhOr
vn3Zy8So+ufbIaFS0c44EcgKpprkXVZcWdOJ84vKyAaYH3cgiywFzAU8eJtulVO2
glAwioUbSY7ROzwT825WlJu6iuxOpZhVUbxTipVs9QrZMjYnSmeJNXVezGsqHYYy
JDI/PVz8DWSUhc29wp2Jo9nnEs9Lx+iiMPASCTdJYY0tGzw4+xgRZC8i5gUNHXOE
JMXtfhe20q9EmCkfyKo+g3f9UoTI0Qz9eUibk8O22XekfZ2tPxE4CmI5546anfbg
nHlvS0lASefEf+8M6NZNlfaL6S//q5K/JcjRuqggRp/AkBrqKX7dZb+E9NVzpUKs
W4QiGd0NvPYWBKmvKAXu/xO74SuqplD/xfYKN4iGSryEA9qfpS+7E37SaVj7FrxG
ZX7nRpucTL+72YMgFKUt3FAkx4Fleld1tZNHiAPf4rEDfUTAVjTAAs86/wcySFK5
sThVXZwYJIxy8O8NfeG6YVY8HKUNtEYcUwVzaPbU2FOMHaRZHpyRziLpwhJ2bcXf
6YApP6xb1WhSMAFZqnVr0/bH1l3WamVZMmUf9DoVMVHs/s15aRFX4Iibjh46Tt8C
UiURikkMTt7nxAn9Y8z22qe50Gf3QIipjhJn1kPq8AOBCEhLj1jbgZKYiOMjLYct
2wmsd8xjQxC0xBnX5kBsiJrQvwtDS4wr1JxiRqkbDQfrluzfRxzN24aV0nbfEPQn
SdgR7XRRF3as3V46/GtLdQ5ng8r7JSQDS/xDEaDJntKvKeWgj9zv1S5T2DICkhXX
AmNorra4IBUOGz4THDhvoCuEF042Vlx+q4uNcn4ZrmgYsQVyD7P9NX56MS6ftY9s
r3Yeu4jF6Sn/R/u54hBWtgZxvkBAhjLZL10CeL5pe3N8MwDnb98uP7Z6uFLEn+jY
8bq62CEr5GtP0R+3p1psVnxB66pKyYSGwAR+qbsHFwNiIEqJ3za57VVJQnBEC28q
1ldcvfi6CdEWUZn0VTwk3bDrnvXgdx7QQorD1L4LfM3i2Tt0Ks7qDWeXkVcINN11
uXOGvbYb/tVrv5iY048NG7oaEPn1qPdy9C07QpfrmAhJiyu46R23lbnea5gUpfhY
lTBWHYOE54m8SVqIWno8KHTLnaWbCwERTTiCCQ1UjrLUmTBpNHBx1VOirEwiBdyo
WliuvZokp60q1Mpd2HOKPNozxh260NLGF12zB73pA9JwhhYJ8c3EsN5ZRJPxPEiX
3+K957rJbtUIUS2xJuG+uNZw7bte9EZ/OBFGd1tvjCtbJBXXersWbyO8F7t+W9R+
AbKzXvXggzF7SIIvAb75tRJhKiXWgmodhooOC34jAsVSKAYlMalQ4TpD5+vSKV2E
kH+E2oK6WzE39WAEb1UednCC/FmDVxDePC+cLdoVfUmXBd5juJSZ3Nj9Wy6tF+E8
S3+OkcxHxa/8cpyvBl+LY6rJeKeb1by8gWaxE2nTFku9QxaO8tTQgq/XCzCmpXGz
gPBIFa9VplHV+1vceknGHUjfW25AxbhiH2TFbTfXYXXf8bXO67Zufug3827WUqEb
OQDzpfetW5JXtp27O9H+ZEhXfoNyWx8s2j6r7P80p6LJIXkl3/EqpiUIIEzrhMoJ
GLOgZ4YoRHuYSVY88gNgPOUCZ1GRXGN6v3/XaK6kRRy1AfYlwjShairrGN9L0673
aFI8+7SpUajIZKrKr3b7VY/xI7H5iaf51wbDyI0KFm5KEPVM9Hw5jajgoByEMA+m
X1xn+dIbXmO1o0EXZN0UxUdUx4Dtfszf8Sr5+FBfWxeqOAvOs99qcOF4jpFtkdhs
kH67S7TXFfJ+gJMaZKPlXt8P6PCdRkjax7rMrymCGM0Xes3eOyrOuOFcUDplBAsA
bHH9hmDwh+tlRn5rzWQWNwDRU29zdBNeVK0rK6YTFtqVo3KGOVXU7a04mSMHcvVA
fcYM6uUmw5vv0guKVlsAKWJYhz/R0KDpOXhuwQC0758OybbUtc6bpmdWYmePMQqP
OWPcyyVEBGbgHa87qh+3zT6OHW9sn9ANBoOiy5oVbSjDiMealwGT+91L7Q52G0Dz
PLgJVc4o1wjSMfa+hpYW/xkp3BJjn9Z+/y86hxxRsZ0ZOGnZI34OxHQGNOxtmT69
8cMuI5uMdGKoVE7tghoNht9w+rIIEl7Kjf7er9RSE8Bv+Gx6yJ6+4NSiyu/9AM0e
zGI8CNOkxFLDZ//ajl/gP2xYD2OkMPt2SAJoQrYtaN5ZjDJRljazWIu7LO20dJQk
FNmsuNdXPkGrJ+H3IMx5SkydtR2h98crE2g+g+0+Tvp6a5Pm+95+ae9IJjmsA6WA
Q80WJqO9Nnn0dRk1AhzkdxCQ/pNXATPazsA2HC5KnM+x9PZ5k9GmfdsylyPpfa4w
MyRSX7EDewM83y0dUZILrV/4ALY5hPFBObchF77E0TH/65L5qcHHWucIqpLsj6V0
ZdHEUMZM1A+Q3WlBGwioIIbr9fYIF9MKmSH/zJbODRW/EV0lwIpVk6UkkwYv7DAh
Vnvd+r0Ph0Ou8YH+XbUMqKSO7kaMXM0EyAf8dQ7epLdYUhYXDcobSl4oFZHIOlSn
26cQek7BIBYNb4OLzyq5xVRMLOGvSwLjP7VoqVdXDLipeNkiVThL6wVKSsEL3+z4
Ye2zn4MrhS/l8FLcrBmwHuxaaI3FBG16o5kMhiWte9v+H1nAw8NokY44B6JqcGCT
UYajb4fyvn+FC4N3UeRVvOdI+0cxqwZiurf6wJnZXP5n6LwjvKMTSqMHX9x/fakm
hTsiQ51mIpeKTlvPJY9dh8KM7T2AJhIAjcdzQ44TvQqBA/b+9n+BpSC4mrRPOpDg
sb1aI4nGX+/jrRx8qmuy+M+AZntFwvw4yL6gkgWr5A0e7p/qnjGmTX7CzJtZDBbM
FAqz5weOGZI6COA39/+5z0HKXMwGbbDxTgME0eB8hClKShtmX4MKWkV7iEWcyuID
S9en77nL/kkbEeOkrXnMDtHTjO3QdHpQgL/PaXGm7X9RiqeHc/TH6D+i7+9Uk5l9
bbpuAvEkgiMQCXOCsnBoqen/S1RcismAWrOofMw4T7PkElta6fyZGPVEHTfBhqT5
Zkywq2tAjgmHTu319SpA+g6Vlfo2TQgnniIRKOFzt93l58g9sWZnKOt9TE08DnPM
mBhKYSG+de35wi1+OUHZhYfrz4SWmAC2/c1buX3/J9aRd/mpPDNRZ1xuHXxEfPIG
JV3W6fj9fszLegScJ2WP1Xi9G5K4akeXaW558tsmMht1y19eddPkdu4KAma/s/4I
UY+Zn3rPPc+W9K2OSLT9EQoOIxE9tgQ8TPjfKQ3sweGW6hmVAj2pjT6rPPIAoU5O
K6dXBCKR57BWHWyOXnofUAbD9lDP5sLiH8yfa5cDk69ktubt1dZoLEF4oBluPZ20
J2FPYfczeKCol7NufiTIpWcmHrfrOHARFHVoeT0Qh+TQ9QyPlhA1+nQS+SMAojWZ
MEsJKvVSbvSf8hkgf0+2ce15RgW7om5hULSreI9nBEXTWB06E963O4nzcBSxZSdi
DgQ3lwhwrNakxDmgdog3/fazxDrI/NgSRgpqK34ydNtm8Mxx+93AlKiFyArUqLQG
pKw2tEGj0lSfjQjUMJUlBpEfPKXyJ3QuxvAOrqFZ+0FpJG/gPFxsTzRvjPpHXuv4
Mkm2vcdZIkCmPR37QdotuW8W85TZ8ovwWDwzQIFgKFpcsRpkphCkkQSu2B1IpdHO
EAYeTrey0VKxeVvch/POfDTZiHUv+t2n/AYkbAZ2R0Nceee/YFIgc02sRKGIsZCh
DtJoAkpp/4zdYDis2ZjS1BFcx9pB1MDlIk8dCoh+Gjwnik1Q2ES3FNgCWBsUjVEG
IrDCSlfoHIYGj6tUZq8iTbE63N1NAyXBpVBo5242WehZdNc8rHjXPSzYSLr/x/Q7
jGzPjqsmDR8MfdYhg35nDupsYlu1YgoRpp/A3vXhzBPt2/zADQvatzhNEJoJam3y
dgE7vfKVJhfD0vKUuqgzh7bUkhXPztJI5/CfHX25pmw+2aQ6A/YtldIzLCX2aq4N
hFGEZM1A9Jp9TqnQR7gcrpDqkHPdDs9XCtaaAsyrfv2tI9jQI+7ZFHqUZrX5b/w7
ngosuElyr6YsX+f/p7PP6sW64Eqnm+BqwaJmj6GHYfGZHP2NNT8grReFTpjw8pVu
ZhFWeGdzWfSkcuBsS42gX68+udburUMppecL4cPR9QNId5b38XsFMeOW/GRocXrO
7Hj99nWEVnejviP/C9Qeb6V0SRjeLwkh5obdwU8WSboxJmAcLgG0pf2kKwKzIP0a
aSQWjxG6M6EJwTib9BLINsqrVIA2XA1juVo9m2+FghNJWEU5F9aAucJvhP0oS4xW
GASt3A2/4AHO55bY3G0VUjKeL7pGC8VKg8tsbaGcTjvPM9xzvPpb5MgwSzaXH+Mq
hBZxwGmKQn6vSy7pRaq9jPnDgrD2PYq4IuOwaw/+iLsOueJNKCKb1R+1TfXUy+jz
Jhql60ZKT9XDcqswTRoMyPKA51nrC0Q8kf7PeKbSbRSppUjY+kQ6kIi7/OeR99Ar
92wgKBeTZ/IolzVV0MscCmPe3ja16VZ3mLWpzI6oiMWCwtHiZC50m1kVvsa0Gf67
wEWU5xCP9o9pMIkUxOz+tS9FP7Dck0vU7zxnAI5WA1DUHhi+v4ojtB7bnokjrupu
U3dfGC6g5ABoFWLFPy6Beu7PNhP9Fj4Woyu/xG2e77CK2hMSmOzDf5NyoK9JUbD+
A5ax6xc6iDTs/TLnbzpbIuKmvjOY84I9Vze2EaY5ltY9H4X3CJwOUX/PKZlkjplu
tch1cpOF57cqWLQDimwNQnuc5Yan99TRRlgzXAJZqBo0M0OPsJTzyBZWEjTKg/C0
gMht5ec6aMY9EEk73egCBQmtqL8djMAVBxgEEUI/rfGMzmuC4qMVfG7ukn/hTriq
aBlbujZ2bgjLNvaslIuLUlDNGHGT0liuq7WkSm9tLBfaN7FB05lAGBD4keqZOYS+
LAcLqLWAdplfdg8jZJW2gxA6oMcmbemEonO2jSKk9Wv0LCW9CH14xJiNuHgSOTgG
bEuxbZPWIf3DMUnDd1YzfzQU57JDEyJA18FeDZif5o0Rpva3zpqSYAmhhyVDgInu
pkP5Aw3s/FnO1bwylotjDR5Q7tJwQbtC1I5zkzs03Zjso5qzJmANxfrAkdibO8Ni
pJimM+2AMH38NNNPOHWux/YlCEM2jb7vK7KcaDxqwu800UPRjoAgKizYZ8n6E6pJ
fuNvdo1xGjkuiEuJWMOg/idMFaxCsfd7p+HDcveNupDM6qqO2HLyZVmypburHzd0
snvr2gAhzFIm8q6W1AQHLM/NIuOizT4xTfSS3X2h6PFBY0K1wN6DvApHWaWofB8p
658mGifWgYibQPmXIQOB9Btd0osdwG2J75xLdwfmERXj8zpenuh1O3zlhEIR0war
265X7gEJ/212E8XQHcvBX59PKzjb+L+9k9exYYJmXmoPjuiHcmWOzlU4qBGUxP5O
U/wqTBJZiJn7DhrPvD0cDRhc9dUU+5cVcYDQAY4Km6bE53QLZie4eHweieKY7/zy
nrWrymTxrV82GRYifwgugXXWIk10bg91JlW7OsMLsh7jHvpeMftJKW3ZPuVbjQqk
KSaSodjh7ZZmQVgPhnrEhTAWOgY9o+uTY2A6+QsVE7P3BAZVFuzViCHNqUQtDLGt
+8SH19zVeWHX5XMGa2eL1LruM7j/luMoCOS/gY68h3NcJtWyh+otJCCk6m/SMEVs
qoysPYgL+g1EFE2aqdxkMrG5yp1gliPhzGweDlmOZIcn2Ao4VYiEvL++ls+r1fiR
6uaXbkoLE1JGFLqxPxzLX8dNtvMYr+auZBybkJPrTDhOxtRpcNgeeOG5+yXKCERE
gSqu9KCgtxatiZDIjRQRr0acNrFNnhJgZj7dTgb1HbUsvJBfuGnPQJy3/YtliXdx
wloix95+RqAiVlIvfNMkZgLf5IgUjZ1fQexl97YolE63Zr6kU9Ew8rAuKHreN75M
gaRBdIszrXMQSMpysocHbur4bMA38hn+ULaAzx2lttVSD+gxvWjpG5w7yqj3RDMe
vLDrCxdOw/RvHREZyHkTOA+cJV+/fiM8TNEYXV1ItixP66Wu8rBQNhZUQUpRHQw5
Wtqt00QG1EvwGjLcbJJsYNvyCvZtAOpFdNdpP5cG995kJOzi3gjTMVBwq2pzEz8l
mleM/GD2J0UhYNowbb8akx2K+qDeh6dS/sBsybUSshwRPWPuX8Gbeh4NIEIK/Y7q
9wpuSbEtyfeoxC/4lcnCyfKoR0qTOlfn1xVAkfoHQsiunAQ9QH2VKHmPqfm2vsf9
5WV0fMUxcXDnBfIjM8OsDKATB3rJIg3yYJ2dzoBOfrETPStSNpimpaxEDJgkcs/B
Af+ZcjpnJTM7BXyRFlgue7mm3IEHuw+02cnVEqkyI/Uog+tKKEXkNLg+hw3DEgnc
HCd1iub+FbxQv18K72TmmmMNXw2NhxOvt1qS0rZ8tQ+CAiwtz+O8hiH7giV96nIU
47Ot4Rk13Yj9885uJyj8pcLBDN65Kl07BnXYGYT9zJrJZ/J/5CqC7mTSBUs6X924
qdTgduFecq15wZzMG8oNfUxVtrNoqcx/JSH/9Mkz5G5Jp0+U0F2KcbddVzD+n80v
7aNpxUD3PcqUmfmLhLAgkZy2idjkfOmnBxDA0ZAOPGLclmmUJqQLsgQ1J7VXeY+A
YRWl1u2vAONp4eEtFiMd34+FLP81Jip5cBeXC0gp/m0dsCsENmlBTzgp/fYgODH2
pJBu/yXxDm7AeH++YDDVGAXlqUhWEJDoz6CxAgL2o0PJn1FuLv4dAG5g11g56geS
L1OBXh0B1izRPr/IzZjZ4DR5GK/pwRydOHCl8UnwwW3h4nS9gujFZMnSZnJ9ROdV
E5v1Z6RBdjQv3Wza7TJA+aVQj2hyElzoj/FaJJ5AS81QkrPg25NTUGlB91cn0vrU
OXlKpvOlAxVqLP6cWbOP8HGVCB9oLPyg9Z9UkHXB8ZE3n0z4GKrAgIpqAEEmOCrU
1cVEanIBvzLdjuomDxdZX2ArhSwghEwi8U8F5fglOd5I59g9NkYJa+iri4f+bYaz
8U2euR67IpkUq0JxB34DJQwH8RYTGj6qJiCVCVQGTCHHFftIdspxJX5JvtmnYIiL
AGPVmIQNqfZMFf705LteBKq5E2t0VSqZPWyzZcklne2vYhb59QwhXMgB7Iw/dPsv
IwI/UoDBGnzPu4R+re3aoUddFOzmDoCLN+lgV9mBzvimqaVoSXwgwprkkiVY7rgI
eP+qNmkCf4xLrEFwUVZ+bzReUmJ4qE4O6/4//gXOKFYLBJO+PimTJg9ord9Tvh/6
o/alTV0qe0rGyytKV4JGzr0R6sx28+tPFVl1aiT+BnsZlHV5Xw3zDw/WdP3iezMe
5c7Qv9si3BLI4F2AkKknmuVf8P+A0cWBn0mg9Ssj4CY4p5TRwqvulCuE22KcwUpY
CHBZqLqDJtZ7RdGOdft7EbkV60u8ayYtCdF0jSnqXR7J7k0Qo0rxSfkFnsYvyqrl
2VJnreUalG7oACnZWvmrgFTY56ovez49Usd4gcImRMQyOeOcH1/11U2kBhATl+ol
KhrLn4y2bFC1nrVQrUgpUsoQRGFHLsd9UeiZ/VWm1vKLSb4puW5fs0iWa/D7oAEU
bHAl9I0TISZupziR16a7S6UTlk3qLa4zYMvcr5ECpnYPSiJQqdWHs4g0vhTcyXRW
c4ZhCp6pVHesXMehY6iK2We+ArUfVckJvAPFR/FB0ggWROCtQNiMZ+wexARUCKhp
sI4BzyMUCki/iV97wr/aRSOofGrSYwkwpqAdc0T4DarX7/W21OFGDZ0Fb2We6eYY
fzaqmJrtkAmg3BjCsGlmD1Jlq/9ypb72B90i1oen8STTIxMZWI86P7Cs+OBmwzde
USIWy9dWyj6Q4lxC1EFYMrsNzvxQ6oF7HK8opp/RiHzrCMDHk+OBSTcEu31J9RcS
po9HdAUnWR1dkla1YIW+NxShhdfUCTqhgnascPKMoS+f/FT1v9yXpO/TkFsj1M6L
ZZScYt+WKQVpGiI2OUnBRDZLbO/OgnX5i2LUAAa4chL+/Monofa1nahzI2/qBkmK
CWk5c2o2mEp3cJnbLrntJFus6GyeNIvtE0J+7PDt+AMxbSRvhEX0O0Z6dj+iMT6t
2YFmwjEp24EuFLPA2EY0cvfklqJnatGuBQ7d2Of0/DTlBb1curhMMH1ntK9fgDFy
CvHVUi6uBEVYTDxXZ+K0uu5VE8TvdtAIZeqcVEYIJIRIihKXe4BK2rBS1aRjMMfd
asAHIFBe117OBzsPIRo9pIYxwWZ8r0hhAlXNmcY1w3FMDoTyo7p+wefTOWVFe+XJ
UoIdnDQOOAAAFjcvWyaxZE1DV6RMdWUJnEeJatLDdpevG9oBrB72IiyU7cwApmc0
a04+GrJUk7XDicags+F/PYAp27BLXn8sz5Io9EaEIsTNJgTER0QQwGIGRa1qX4NN
/Km+W8eOHO0o2SJraZwMughjOVsiJPEN4fYLuDCpQnuUCU2pBo89pMnDJSI926RV
s0+lolubjVmS0P8PGxl/1CoX5AuWiBIegyggZvErqPdZkE6Bz5RR4hpOio8hMu+g
UEQSexI1c0bTiKCeOzGEh9Ya/wRskqKSY4fuY0g/THw/vXrrB16dwslE4foH82SB
0hVVQt9m23+30HRHHKSH07jVXTCI+IvckgIysBtlX03JntSEUPFFYWWlvCfoQcdu
gVJiXGb6qH7W1eJ7zmtT7Qx/pGhE7j+S3uXXbm/5JueU24khONmt57h3prkj1RTM
KXOp2vGTkJEMiXA8TWtDb8idZmaXX00+HAiWQAS/xtsguUva8dLj+DrSJE9gKyWL
WDaO3/bN8JpCv8DazBsF+1t4IPoKQkIVQmULRToJObc6ilqLPtoQ5YCNTDaQqObo
FXB9LlWH4DMQQhzsIp22KS5wZgiq3JgZwh02CTvP514WXuRqD+18Xhe9sephTheE
bXvy/IBxyLmLihFPvGlNtRPeDvTXgCeqo1CEdgWvHN93Qb2HlQSB/oBg0xtdnmlZ
Ec/d62JUNPk6dbDanv9qNwjqhLky3F0MbJPeIkTR8ZhsIjemHKyXLThiC4/W+QlY
NyJ5W24+NhB4JHnV07v4Ayp3ttvhXXgygrwfAtDe1SfWuJySJ7/FdgMCZ56RWUhX
K6SEurOmtbNoVVd5i9eAz8xySWjQuVHFetSjciLJgp8orUQZNvRTGWtzJbSPlxBM
1iPa+2c2INjJebd1pCCI09nVz9EZbcdIs6ZDxIc184Iad6+i8T+PPi2OynmKWIhl
tVxEeuvV/10rxOKISbHXgzh10LScsFDlBWyv+sgCNTJ9bPpU7Z8gkft31K2c9rdT
OUXfmzBD0t6JMU/nJa4tuCDe0MTHdLg4F+9Wz7waHwZ0O0T+oC3xdpw4pI0B1hWv
4Hasr+Ryao3i9okZmeErBEqP3FRlKA/G/kBrbbSJKpVANodf4nvURG45MG0ssmpP
w8RVSFMZTuTjKRSpk/WMuW/IRQADCPwWLHXZzqy5cLFxIoVYbwmH3HXFp5Z6s5WJ
wnf8E1dgicDH5IPEdbpRB9eNKOR6hs4MzqPy8sDvo7hyCGIMRXTPYawCCAxAtIRf
bvHyUf+MMMDma5TPgzuIGdZvGIy+sgZ4uSy0FGqlAGOibgNFgy8svlphMTMAZWUC
WpYXMaRXG7Bx+plLs6sZ35ZOm2fOVeeBapsS6jl9nT1UujH0g0VG7QmL9MdndsGy
A6wIQQn9EIZgWOokefvVZmBqRIS8fOBwI+oTh1+zJFxNab9ggR2QE7lQRORMCopD
RrtRWxnWZiC3vTZBEpVWZMUyna16+QcrBEmwv6/+VbLDMCRcuXB/GR/DGhgG65iA
DjIvwMbapqX6oiw0wYfP/gmgcgJqLHcMnROwkym4DgjgV3Dmuw/3qFby5Mm9/dF9
NBXUgcyfgqx67uYniYPVn44mIZEBf4cCtwTORkBBiZGfkV9qYC5NSkz1E0bZYSb/
nwnsKHNMQSYcEt1qFcu9d1S+hus7/qMJDomDA8QpSV1sJ9T4JciPRoY2DZp9ncZ3
xQabP60IUGCV7cMzs0s4SU23Njeckh/TzytMAKBnT6m5+qzI8Zth/Umd7vVUvG31
LjMHqBVsu3m/iHQbXktl1cm4iXOZKLqKQl+iDghob9/E9GOS801HEg2nl6uVsvP2
rsjaxGh2txmw8F6XJE6GNNFW7DEhjFTVSsmVM9ZzeXDIGbNqc+BWL9f3miED4CKJ
Kwz50podu4Hoa/1mytTmwotAyLe2YnmqSJMo5m2GNEC3O8vdf7gxc8eZ4mvV/qR2
hAA/TogRhw2jf4fgzWcveRJOX/dpNiLMHKYObdw7IdLISgbN5yiloMsXx/jFjzbM
7VMs5h12+RiVYlZvyraMsYi0CIV+XTpPCCf2ilVCKquf1DMskEXjWXPB9YW5OV1W
+5c9d1laj68Rqv9ziQHhLO0uaNdD5ashkCXB7a3MwqfY5B8sISIel7rKkp83GnI9
yOhH27OQ7Srk0ebki7ZG+lLdhTZ0b54k0nrjXCaJ7qWwbZu6PPDIAV3CxRyzH2yq
Ydrl7LOb2sVWoBTi4yyzOWghqthK8rHBQZy/o1Es9X+hJgPhR8wqMD/IfNvfGMmz
YUc7nXEFJZ1Q4EAumdt8/ElXk/h2ii6xMt4KsrkES0R2Nt2cEtmhDKMeLArweNAR
pNVGDkmcEmhw88CRgCq6yiDVrSV3v1m+n+LTaIGkf5f3VOmbkwya+2MIeuez24Zd
KypaRmzNkHrxPCKfht1EGWYNkPFWK8j30Y9bhQEn1cw3fQT0kvqtkduJuMn2tDZx
go7WcEPeDFNh9XlUfZSpWNUlBuXL9sWiXCksRXjXl+kxjb87F3YceSB2j+S3+D9k
/yxAjkQbEAZZyNznYxDQ3X3e1X9bhd4pZRjNmXpGqG6D4QLRTd0RS1ABoGBEa3OS
zsJja/wafgrTfnQPZ8+glcQ+f714cKknXC71nhXXRG616N5OK4nxWt1B5j1P+cNG
oKk6/VIX1jl0vYdG1q3VORXzbBYtIrRIFMOg/FK684kwN6/2SOOkhFZZNlwvcXOx
jhdD4ayC8WQmu/8unZHkmBdUqhWqBwU5Kp42P2rUVshpEuh8VXu5vqrd/OjaKnqD
/56lZYDff1Eq8ecgHSb1aN2WkXQGnakmUxvt86Ms42D4OyVWp68IZ2m6uAt3dtC0
g9RwdElhP0QRo2DDGKI3WA7U/mHTvE6GK3SsT66LtYZcX+ebmVM8H93hYydz7/3h
ADVhVGMJ8Oc0am2oe90HViQP5xE2NUFXpHLGoHGVCsCbyxy4qIACA14AdWbukO7K
/OvQ2iYw2gwx1oMxfRjtBMJaPYZAU1x9qVSeeyL7kTL6SsiEYcMI3pnDhzQ1bnF2
udkooN/axn2Uhwd/p9oIaCAvDmdKA+7Jjy/TuUll+pxMaN5+Op0v+eUICJkwOdhd
d+zc9DjJKWNPC5VAalwcId1aqUyQLCtzKjDj+CZjz2wuHCmDo9cT2pIMockKuz85
le+Q6Et3HC2Bs+Pz9823sjVkS0wPE5PoorZ5ch+bSkBhyAJXOzQQthkgpsLJKHbb
iphGiSClUPAvYUrTJgbRawUBh+TXhEn2t/zielneuHVnnzv9JXI/0Rynwdp5PJsk
00qiW6uhL8NBBgSmyuN3IYhMljy0fYsklahmfEaeHVoGg4r8G2QkQVlegjosKxfu
PEzf71xH79zO8QCuCEJylSIuBrCjRLXF/6Bw+3ztY0vMXfN1307UCSKEaTbkrjR+
dkydOFzl+Jm060lkpmD282sv9w0d/gwSIRMM7KUzTnNrrP/LGO6LnDMfoOhbwAxr
jcwYsIctZDvHlOgbx179iO+1jdPK6IlL8Hj7Sv5X2w5IOoc8J3fkGpwwL4yTnbl1
9jKxV0WernqBiLM8LBy35yjWTnREN4j+G4eby7jZx/1Hk/NB/o3OsBITXWF0knKe
uw1+vxeyWdCdmgBVtrlib2vb0NVyRT6St+WbJtrLGlEcN4SA+Xke0/fMamgR44S2
WIwUQNwIkIuxU+hppzhsVrw92im3fqr1ObhuD1XLsop7B8CYvBvJpHtMkOkCgmJd
sFtir3qtdnYxfvZaMzSuu11LjLagspTFkrdVh6pde11xABewWuwvGkq2A3ETsIE0
0oZ0NjKp8TdghVuyNm6Z/B6eymKCugz0RzyfMSMaWGTiSY2q8yjcvzD32XMnE2O0
LaOM0OXwOHq1gxQn8Z5P9R28oiPn5K4zZmkLTQY/+Eu736CTzRyH7I9nn1ZcrNU4
gP+VIgM4K1yFAT7guKSwdfiJN1JwvsEW3FTmiYRdhFTVVsIrfOrbDsJXTJnfYBKT
h2n1AzP2YffsNCOaOXPHbvZfw7qkGyUD5h/NoaffQ/5uw8SubvYGDmzamLabwX5b
CvaXmiALm8tj15P01e2j86ynlV1GgzHy1xXnsecGnpBRwQN2Kz4YHaunELC3rRWY
/947CjuMjlnPn/BMLI/zSD1HkoBXpOcFCCGEIwY3IsjRGOd05MCmL+OzMXMCSJ0b
moLQ8VQ2+J5Z5tj+UTxrfR47IUg2cw1x2wIfVrQMo5YF2QJMhu3AhAsX6q2rBE/0
QMGJZPM1P2TYRbV80rwYIVkfvJFyTNoVK9IHYa9qygsaHQz81Ruk74ZC/aXcZDwG
4fqcjRTNULffVCXEZ02CYd72+DTVGZZo/R0xrWfdypcY0D17ZRY5zmH7G7YibKzZ
p5QbCmqx+kgy7fNrTmtKCl6MsEa0CpWvL3QZWQaGHk3XhdmG7hVF6m4L1EUlqiTz
WKQYaCUa6iuof3IR8WAR0kfQnLB9zfmMXJw2MSGqbhUxqeu33FQhLQBeasDX4BE/
D2r4D8x3HlLMg3fjhcAI0JYyllU7QD2QF4L5Yc2LFAOiI4r5aFAgEdWIp3yLVYRR
6AjjPMNmbqi7RfB15yB7lTuJ2BBfj814jJG0MbBZTd9mZ/zU1SH8nhHGi7merNxs
P3Keb5rHn2F6ghjMWTtiCxXz3pxsqa36FnhtBPg+h38t7GohwXC2RZZ/XeddlrWu
FhJ1qL8n1QDl1XDWf6m1R/vdEh5Iy1ROroeGgJ41dQVQrKRMZAVuUlOfH83g4V9g
sFjw1H+8f9SzIjPA4lZFBt47fk9zvvKqfnyrdKii0TDwV3rQGXbrmqYK8eQdqQ/m
hXpAuHNda+tb5wgHNRwJ8ofRxG+C+bn7KAn34hIWHU3wYrLmHGuc7OhCJyxJ5w/c
9RMejR+IvCaFZhU03sszRJhPTB8JTIiRDJBcgTPNripIg2QuJM327dCkZRVz0+9a
4LI2NtEVtd9QqEAn6kPkj2h+fPuvAIPPNve+Wz/IpVWTJH/7/Tq/BOFhOFaAQ8mQ
kJKXc9WypI5kDMQk4iZ9VOXz/VNbcyUZ7LKfVhjpX4YPEBEnY73F797oLYToTgu2
WpUBXprjaEoumB/287hk4a6hkxrJXuTMfujupgUO0AmA/HnN01mAj3R/+Jvz+ULS
wQ/YN9sKRj6bxsS7p9osmPFuhrEUXplc2gay2cv23SX1ElYuqIgl8ZnUmaBJYu75
dVIzkJuj36xaYSvTBHowfetICpumR3cVsjjQhNOU6njjU+yJVJMM07Tv/plgk3qt
rBAgBF8Ky9BgnD4QVXlM/c61/MPv+4vuLyR/6mtwqTwrDbniuc8NHPIlWvasKhjg
wIRocB8pafEPatvTIcTlDi0Cyw0ODmV5K6htu9r46bbsbQhsIsT1uhpgSZed0bJ2
geD75W9Wm0+fjoyeWGCCPtFw5G1dmJ6Qe3l0DcCsomQkin3biVee4YWVDWX4qZDm
v6WtS9c7VePqVifUSSzHk+WaMukPbZRJ/0/VBbT28y6DxBOuKMbZccYrAM4WYPOV
X6EWUvDhAKSozWuvmp0NulkfA3xmlD5UCyMoqKqJo9bRbRj5MGv2cVdtleay2CKm
BsyH/t8SBdA0ZufhDe79AGec1F5NRqTsQauwUNDB4nPUMaP2gOfLIt+kgqPxm8BM
hh/zEEdgvNLO71YCki9wi5cXoYNlxjJSW66dQNhpguNNoYdevaZtM7q+EJnq5DrH
XEkzU8moODjH88yHLCAEUfQ7AVigpUHuGkj2PTbTFH7zsk56bAPpZxVnGAvbj862
WCKAjEXhX3dFXtdd9wJIi3arakDFe1uoY/S1Jm6W9fXYMl/BY19IZjIF5cQRNb2p
22dQd7+IXNcVMkoqFOIUhPXBXxsV7mrGthb1bC3K/CJWERC/4nicKLIPHMy2f3qm
W2udy1k0DTmN8rTEshaDlJaQILbLTid0gzTZWKaki5Q7GQNZODWZbpcv4S67elwD
DCaFMy0ciTVGwI5HtcZZzIPFP/ZgFWSAjEqyne9wYPRCx8Ix/j6R9pjHRC7KZjoX
OZVwM+Tkbu6OdT1wt5lhILWRjgDdnaELGtGswkfRuNIESzPRGIdoINQPTw7o7DE0
owT6T9o/VLesMtBz+te6pvMsI0Fk6Qq4ffGqshd0MjZNazNweSL0iMai7M10gjdz
07RFesPr35PKaYxtwtm2+kP8o1CTW3702CgRaNKRLjvpp94avtGR7H6COkwbvmJw
kPb/aQV0WkUFnp0EtOAus27ZCyYKzJ1VHWjr5rIcmCEtZ0JuGYThq8KfmbXfl8Pd
GwXdIIkVo3TFEjgJeCPL0f/Wb/ePD7P6ZQUQvQVUrLJiXT1qWcffKTuSVWsxdy8X
a7oE3Ezc/MouuKkLVXlFPDmuNzq/NJav79ILGdD50YHPv6RqO1pFSO5JseIwG6a5
fIqC6F/ZYW2rLQ4C49AvEKK6ryBcVmUtg1fGX5alhvKnnCpapM7PdyMniC+yGtra
TePt2J/GuKKL3tGz2DN7Lg16SnFTQ0HI3jw6kHt4gGsQG0HnTZdkF5P9nWEFyxaP
RzwhZ5A55TlalMBIePnPUznpJGD7xD+mZdPI7iCixK2FtzYeVbodRYklerVHSdLI
6eZ15tMh8kh8Fiz7v1CBlZ2vCZZKm/TeOmqlY2mnDEMHj2NYY7ypt7HL5LttkTQw
ROJ5TzT6nnDeAfdn22VAYKFobUvj1WevEqNwgTQEYPPlJ7iYn91vHPLds4un0rAC
nFhgeFj+JiLk6Lpxw4CJNx/XWGcMK/G3BJ9JKS2GlmP/lzC4lgsqHpXxBaSiAsLo
EFmneg6Jrk93QgrxKglgpFinhgl175zxoLKnHaECBWr1JNrNtyUJ6QjkJ3DE94kx
6iUQLmOEPscUBPk3NVr+d11v8N7yiCQy/kPEyKgD0JSDDM1sjvdGtzAv13FKXgzC
bT/urCxM6CxLTrcKmzdcUwJZ+Wj2H8EsspXfGkjALVCzxIjqPDfiX0+N2j64AUfo
6IUY5B4B30arYKSavuNaTKKdLiYrif5N6TTasWmkwTUdQN8fIA2e2e1dCk2m24JM
O1ThHG9WNr3D3g727RS99r+SnCBIXBuUBLp/0LRF32LE2WwKbloMnfAjyoFUz2Nv
e/83b9Kqog7l3C9v1jQClRMu8nTedCYeSnlr73AKuIkZH3MVPpOuuCT6iIgmMYe7
/ceQEPNBD0LgO2BjzeHRD6i2MkttTapkNKWB6YRjq7BCbk4A3i16NEkdSLJlDNAE
u1mIh00bkOWrqW5qgOUKoI0IsVdS97hvZAUUtA4LU8kW1VYwF8LrsD91d74zz/3q
AJevsXAr5irO0nk/r9ND5mWE6/H2buv8cFsXstghF/c8/sLIGaIVn8tI1LUMCOyR
AkeVX3GO5OmV77+FpzUADeVo5Mvm9hv8is1+r4Y+T6uZxvzR95DLmoqPFss3VVe3
wI+GwZ3cO0FEXU+46LceqD+9CKCMas+fyFFkRX+/xKOeFqE1SCJC/W63QmDsENsp
aB8qIcPbcistzWfqZSWmk0w5wlfr2Kcd6QGUbAt2pttcTrngHyUYiKhK6wrjNzux
qP+3UJpHtRxHP730tQ3GA3itoOYL1XCWv/eM7KeqwF8ll0zOI0J/jjuDMXWLBH5N
F/KAKVePcjZUm24X1fHRDMzeznDLS9ePtJTnw01Mm/ciaHdivA9emtujaulL15US
o113L1XUMVXiR8SD4KRF8tSfaXzhygCW9/lGntUWhJjR62S/nz9NOIc+9QcwXQgv
BDEhJMvZpznaM/yifRNMNUCgviSy3AbiS2up5AW/Wx+DRbXjXvbOtxyHD3IS1Qyo
NvEH/AjaTpaDW5Bi+eAiXZvPi1tNnkTDKhwIPQhkSUGMVTyz1ocWykYmM9yLSMVy
ADEoS7STrc0s79qTj+ibcWUNbL3HPptMOFM4P9Wv6AJ7f2+alTHvltj15XD8V/8l
Ztn5wTI57P16rHgOSowNemybyXWJBksjcBvRl2swxwRz/H70t0S5ufHBBzlgjBSY
kfLSxQtoF9LpcHEhrLi225z0+BUMCJhByYXCLNxOUcI8FRXSHFvAILKl6TRKZkZE
6ksZhIfcu6/n8oXUvC/H49nqmvhN14Vdwk6czd/kNfLv9ZOCLm5gAkD4DelhOZBl
FKukyl3tjpOQeD5BxapYRnqahDdstobo2nU1fTd2AHgxFHcmS9e0j/MKWpuI1BNp
A/qe+08XJdMcxBittQ557cWNz7Jxz+1kBWGTNQMihL7YBPSF68q0NhKJLfAOqdnv
DCVQ4bHfxUQYfs+mNG3/MQ7Q+un7rBFEY/l6tP7Ph2JOKbUC+ek33TZVjH5RB5e+
4bRe4z+9TsN8JE5MI35MEnbC+odHRfUv9mweFssLQ7Xtt9k3L9T2394iLbBEGOE8
OP6RN1x0zKpDuUFsKE1iKS+AJ+NJBO0AWBhREGEiG3wfz3tjeC5FxrGVN5E3nU9Q
edVf6wARgqlq9ydduEVyTH6uk+I1z1jG1gl5Flpwl94CCqIh6YAOfNHSGQM9oCeW
OR4L+ZXV3w/pW78IGADFb30C/5Xxwdy04nh0fuHiMBUEHH9yhkzsIsGd26Its1Jy
B6JeGhw+8Aqappd+TM6e4ZaWzwl0eK+1tJ5RC3FLogciPAlZ6ybKqnmc8jfbDyc4
i8F/+0bbIQrQPOch1n1n+bIi0otsgaDLVzg8jeE7IUh6czlZ5nDTlupblmjeSWSG
GP3yhyCZ5f86cCEWC9Tw/yXTWfkF8c7YbVul3CfruBCBAPEI1wVY76kAkNd2fXj7
huslakj/thfSOER5fgGKM2/A64M+L+Z6B1CvhNYxUlC/lNxkBMPjz9TIKcFSS2GT
QfPfswyWSUYUAch9DKrpFj36LbcI9Auu3V/reM9dDKXMQoEiaIgWX3mYKx9dasYz
mNmfjlMLmU80LR4d9KTgncuEMfKyfxWVkc+TPd5Buke099BLuB0RJAErdn/MQfPa
lmzXRfJZeDhXrzXxrSEd2beVvqWQMTJoG9EkNBpKK3zSrTU9AM5hOlgUf3P/QLz3
1KPVMiuGfQk96P38ACPWPzPuiUo9+Sv+ePtA6xbn5Hkpc9kEbisQ/gI3M3xyTBA5
1WOQFqLmPsrgki6CMuOVnrFCb0QqxJ1oOxylkcHMINxO2U+vEtQhWF3ySiB3pAcV
FmvG1ROPny93hwtnlzNEJirny8xZDdBve7khvTfN0c1xULA6MoUKVyc4K6eEjvjH
vIy6ludktDadDyEUOg3LA0OLm85F5k57E6wi8sp1Q/hK/ZiJEyC0nI9l3d6a82hs
G+ZA9OUUP3RoVIuFsrGEq6K3e7FwgcTCqR1UPWok8ZKg8q6G2WLmyhw9B3Pu7Rb7
11T8pogGTZNyWjWT2zpmzzKuE3P4HkK2V36FJpSPdIxP55YUwMbXlxC97tEtiBTG
rMsGYY7NQ+AiBaC5c58yvzkRuz7F1dwPY6XeY4Camph6kRs2wbvxUKcgfLWcz/7e
OzPhOga3cc5puEOddA1WfMaUZ/2V86wA03hExrI89rAjmSFhvS/+tIfzbCDb+xTk
7//1JU7bmMioPyjaoEz64wNfguS3SXchH8UTEIF0w2qrJ2ALBqPL/ZUk5RSRvw+n
8ZcbF/EPu6Bhm46tTpAh1tkrZL4z3F7redR/HMQFSIcentCzlkeTkLLcQNE2dtX/
5FIQ3Kn+xOLRYqQc7naQLuhIulT8fyVuvBjcl5/Zr+k53svar5qub/Lzd7s5TeSt
49Zb3Dihf+H8gXvXI8uZProQytTHB+PSIeFIblgcwP2dQxtJSOdB3IB6nUP9ZgdJ
Zxas2ujb5Rfg5Mwvd7Pm0smcbLePk5EQMhGQtC7XCqNaXKziHTtxy7POGxTn7sbi
3fmmSZhnWFr3sYV+e/a62Yv7phL9pHUnm/jahXFCn8UjqldvdyFo8GrSEChntonf
chpM0DWzhMZSuF7DY696zPBugrmoHBBKp9VE/gkZOsumZJAjMEShMSzoea5WP7Yg
datn+bNV7W2TvMQaZpd/lRh8cD8/pwjws6SvOonEW4UV8huu/kIYNWSLjR/Pb7oX
hyPbaYj+O/xYuYgYKV7YubMkGyRwahcOU5QeiAZOP7V85wBt5ITMZN6PynoOhWYL
VH6IFJaeONmsxnFkmcMx0VHQ3pD1RYw21O3M6glQIf0IFLVBlPRFBk9RcZWXFuHo
2EfwHt3mbo7NY+UCBEa3v0A04c14i/rVQstaALNtp4rGmA3/EIJV9qghLhkfquoZ
4XsFxsOUB2p3byEhRZiOy61+ZM5j4JkvADVSP73250sedYDLMFdhT31KLe+9lGbV
Yspk7IRGT/ZjtGrIL2QUfgZlVDt5G0nn4tHYdp0FjS+lFnaCkUKfmTE9ke+IrrLh
sVevE/u0Nzo7zSx7A9HapbOCVZL86Q9QQ6fknkG8sY/uPqsU7U+in28txrj9ToWO
l9mwNFHM8CasjWXaUDhvLv2AQVJFL4vxwNGeIu2z1hi9k9WKP7RP8ITrLdLW+Apw
IJIJW9r9iZNdSiVFQGMOff0Jmwg45zekfdTPqchnu42lOGk8/Rx1gY+RCSc0ssKY
/U80r08kt8OHpmbkKHmthkgCuTd+gEouqbcG3IhuLBC084Lo5XOkBqSD9LuWxUX0
w4yCS0njujFSz3D76D4BBJlyjQ501qf1uV3GPsMySN9lSaIYpHV/vMYVpqiwPwPN
jY0RzoutZqBw//fi573JINH/pT5iS6v5mOXe5tj+ldEUIRQJjsVYP1NMUz1MeYTR
8epBn9Qdl/7F8bittIFut4+60ebkoVrtU4CpOmr1A5ZbOjhGYfSCfbrB74exS0Qk
w4aEEJi/YiKnOjHoGFzGeryudlVlgqWSKiRoUDHfXCocfZ9Iie3YC9as4F+HQdXz
a+tDXuHYEvquklYizswATQ8TfnkcjZTUQ8y81LD343w5A1PXlBBNplbZRY9nnx5r
/J/SxodBV2rFxu2BJML/JWnxdSm9Ejiayx4C5nAZzXWF5w51FTd8dcnGwjHsHTdM
L5mHL7EDKuWL4/PPgw11AZ3S7y9gta7BnBPoE96Ec+aN4ebNJ0mBhAVOaf0ye302
Te0qWoHr7gh2EKeHgzDJgU3kA/lylxhu7bbsUHuv6Xb57WHAeH/vo3CMRiNOy+Kj
UaeQ8tJh6LcwtiDkbXuD+GbgtKlkQq6oGqHfVDV+T6b4v3i+2YH8at0m/EzRevvV
G+eHNH0UEWCLkTJ9MtxKQmqwWOLxceKnzSYUALi8cfYFGTGjQf2ziEKglKq5Q+Ij
5P99jaQ+dEkEEgHGtAR6kEhqQdKj1ADFmSHE8zVdnXhzeW4jhURfLI/FXll5jsQB
M8vgT3I7Jb+38BV498HP2FfXJFrUkwykE14q3mxSfNqkY+T4+WWeDQBIjKpbYqNf
LgcLLg8Oc8npc3kEQ7aV+X96b+nAIyWlRc80p2YEEASvaCqb2UNhoOPF0TV+Ctwj
1zoIz9X4tuxChMUYL1keJ9ZNKTKk9DJzgWYwaVW/x3QhJGAkFrx/ApXQ4dyiW6bn
BTo+J/vzOYzrVALm3s1yqGWsJZTT9kln7NINd70C9whstWBZnwdWiZC4XQSKjYe2
zbHmGaHZ7u/PZvaXZAyKtL5bdCrq1I5Umj6x5ZfijELF0RVOuZfs8E10SyQuOrPU
L7N7DKbjm/Ox/BMnsrOHwZFAILfqJBisxpsogoD/66X5fwklCDouoQ3qLmenayj7
Juo/VbsIlnzPAkT3/GdfxtJwX8YWEAh08kQDwjQ/ZaQMp4TfC4BUPF9I4Hn3Ykii
9PSmpzJoPO/RMK9es5SG+fSx10rO4vQdeBizZPQ6uhfY+w+WNotS3g4gqSrbv9nu
BoD30PGLfO8/JPvO20cqpNf2uAJAi47MqXRQugW5H3vwJY4sZZnV1bPtaENLkFnh
wVAcTb8pR4S//kGlnWLvAyeSgUBLEPY9FSb9Vcupm2PCCFaJe8H2/0sRpdgCuxlA
AHg8xKrZ7Yv21nku0vE6QY66AN6q4IN4P4hEm9U4hsJyCMr9E5tplXRfdDKOEr5a
Hu+5jPNr/V1nvj27lWs92ED4gmwgKpu7Qq5ZUaEVshsvBBTlZvViLHOCOlDmTlaJ
et11gPUM2witHgeVlkaUtch7y+QW+tXzAYVlGo4y3c50QNWfygPKaHHdvU7MgIGr
VcGVdOQFeSwgeaaUFGiIk2RnE7iWKoH7hSdPK1apF8F/1nr8bG5e0vSgq8y3KcZe
K55pOGgQirpxLhTuHr3kC6ep6/YVrl3eh6DPSMEHT3bmmB6h4ZKsSCy3cT/grV5D
oNxFLw0vS4TIiSPpBlCCUgm99KQJ6y2Wqyjqid7tRWtT7/C2MavGexaDg58SoATv
ZH75fZehiVrySq3Nw6nWgzoVIC1kom1RHA7mYDYiC5/Xv5BuzcLyimY8c8e1h5A4
UzO1Ght96WFEcvVpTP9GwlQ8RyAwNjD7YJNPsluHo6jlkADnYqUyQ4BcF5+bU/4T
+j4MCS75gltt9MFBHP7l7nlj7RUPc+6KbaKCbD2UoTtlHHgiMju7qd5bPDlt/tWS
GrPIS1tyj7jmomhcRcL6a92ZZDazcqN9ueghqP4Qqq9CAZ3C/N/nrcTlqixHe1b5
/s9CrKH5vpQwOeRvrLp5bdNQnKjz///V1b0CPo8qTSQD6psENXRuUmVSUg8GW6Aw
wHfiBy5VOim9h6HBYse+CE+pi0OMLd7zEyEH1RWF7DwH8gbqsfqgYIN7/JE/+ng0
hjEwh7gyRkjaKmH/zCwIDUbE/IvReqY7Cxm6Cb2mv0xv2ZvGzyyAWW6OUJlHcILf
Qi952Qqbtz2lWQb5RRhQq1oYcwjo4jSVHDdY/f5hy7rYRYKElHxp/HiKanujcO31
YCriUkxgPCXNJKuNu8/mJpwXJF9gkrHT2bh+7wwFQ8pNV7dmhc/5l3PeCBzgLDiE
3XONitbSGXb6djIZZhfdPAwnX/0fOWctM9WzCBVD1t9afrtjrvwfVx+zoPcdLA0W
1ZtuU9zTtOSiYBOQoYb0bv0nfs8F4bl6Iu4a1///a/sKKcYkClyy1gAAfjUJ2Hb0
/gHCKsulfr6YQJ0GKLE0OQb/6qEHk8cApu8b5W/wIun6S2qyOSxuR2ne46USI4zy
kpAA+XGlSVVuSTwnTzskm54b8+DefNoDIWaVmN0wjd1DMft0Uq6X7rrIXC6GutGX
ZErsOEk8gw46D5/t4YSG3EBDlszN63axNp1JdAYmQs19wJ0fjOYueEN2EySIPlA8
eyMOr+WBX7xeim5ao2Bq6clJrPMiwxGDASrJNkm7AuR8WlO8wzM04bYGmUXATb95
BABfzLCcLQ5LdGRbBNT/QUxRvLFiJ7MVpFFv1gGzw1EbbD8KvagcgA2DhwzNWTMz
2ScTVxxPVibo3jvUFqGyAb+12mwaIFxygra2Obi2JeR2WdDq0ztfduYezHHS6x+e
awpNI3UViXeWCfVHEjoiaHHv604tFIKxy48ymaqrsocnmZAcRWZ8IPS3H//MjFrT
+d+XImtQj0O3n5wBSpYHn47omgRhYKtH2+ksQWYnLVheY8lY5ZW4OULxq75HuExT
hz7c+Ps2ya7f6AKM0sFfzNsojVDx+UeiGhsaDiGRR6MUii+eTECachIH4U0q7sD7
RYhriAqiHa0RfcXO1r+VAbGo/zASfMtrUscFCtE+RY09Y8JZXEhZqR9ulrOmrApO
lQ10j1ghOc0FU/bR2qoClNFvCOc0oejgnctiUeA6Lhs9xrUWTgAjYY0LXa3/MU8r
Kp9rdOc7RX1EZtSh3Mu9JX/c2SYEyxKi7CFheVsyy+br/J6Kh9JpNlgfdNP4O1Eh
93aanrEW0OP3e1EWtlWxShmV7L9gQvN2h1Vi/nMEB+Uuz0G/u15ecBlLeUqbj+4u
YzCQlr0A046iLyKfw3N+GzCEyHIyDXenGE3pFNZTedy3r90HUT25FK6lx7AdxjHz
U2Z8OPXCqseazoSjsHo2e9V+sahOPJ6xC5ztryb1ZnOzgH07lBqLhfOi/ibV9lTa
8htKrJj9GDtsUMfLLylklMfkibCkQOI+b+oXTS5tQclVeB/kSDcC4THtP4xSPDEp
rkoEaylJMFrfoTLxT0/8r9IDz7D9eOc2Wu/U2JW0Sjn2GAPygHaXtSSBLA4gKIDc
5WfREi8rPtUB/TR5gRLmgp/PPgkhygw5lhaEP9yeAI0oidgJgMR8Fn0AhKYZdHQS
Rr9i8DGdyOYUrOr7jImwd23TR7MQL8sAhyR/4cyZo6qv34aUXaRQ+FDm+fFhfRQu
KNeQGG7Da0PYix/UjN1GrG+yn8i+QcEqAK5XOMCOA4j8m92WTDJfX7C2/dyPWdJL
wz5sX0Qmg3iK+FZ2SMNFQEMo3FxAEE8Q8M+oTJnahsp1tTDc5cJAitRgbklNeYmn
hSTjMyNnmHmzqIXaCZM4Bs7y6qTnN3qy6OaJjoBk2M+RR8V53qd2gFTAB0cDz2lJ
M8OirL9PdVXJic3o5vV3SYOYE12gy051uHX0qcHMkKvF8nkWmWL9rVC6cSXboVjv
Ioq7K9A27Q7QKyLt0X4j7rByE1xmY9TpZ9WmHZ4TLQhLg0ZbWGY8NMMjlRhi0h4G
3pSQKzsomB8eIychO9RAoEna5org3q6zCSoIz/OxTTjwHTMwlOBE2uCc2/r41iiT
1YaRsPUNd5YCzjSaf6utncctEPVgvHvMSA0UUWmQ8SQNZi9QmWkfBv6b0QLb8IL+
W2kzfu8BAfZZ0WcQwDw6jUplTK9viQF9pcVk6WYtQKQZS9FDr1kdSHtocvMbn1IK
88z8EXYM5dtqdoRbHCkl1nYN9oM9akJuohHUWRpHcwL01BeGkoyryM09dLfpswJ4
bVb6hmBsGIG1M3pFyBIIAM+xHG24U5l591YGvqDgrnrlDak/3e3O75X39k8bAMnj
7MKTKBq6y67y0TKYw0YbAqrU1Ecdtw4hFHvdpQt27wTNB2YrtXPXssFXBlFx0sBu
n0nKhzUmtB8MFb7i7s8gc8BpXmDc5uaj/i4v8UqS7T5wIwjATTMqVYBZYL+P6Bkx
HOsjD3HmBrUWHYFi7MeuaXTFYLdfp2fEm9igQo7lQeKJ3vKy6XnkCC8uafvjN5Ry
6P12u3PlnMax7QsCEm1gBplyAABAFKBc2Gei8YkNxXZpUmGeSXkp/iNGlZaYkRHy
040gD0m+qfAjEIOkGnzLKTKevYQic6HRA5AUW13zYwBTwTpul259VhOxvvPIV6xi
0sAjrRCqxggQeVCNq5+/y68lEbJJE1f20PhRRX4bL2g4WtDdZjFRd2Pr3GnAzkOb
AlAi5nS7lmcWLl44fDKntDPTr6RiVlld8kibsmLSe25J1CHbKTGplwzdZvGyz6H0
ou85EhzzfR9oVRL14Mwo99+JdO3PTxAW8QXLmMGRyG5si1UWeXK0K4353LheGb6R
K4Mi4d7aQzDDf7erdu2Uk+nT7Y58An9lHUE7jzI1gBrbQSV2lIgt3n1JPSU+VIoF
kBo8mkdjbn1DyoUNjyYecemffmtNZjmWeLlSZX60yj6jN5gW7FDp0jblkSH/sb2u
lB9SX31hYG0MjuzvGfIaWZDCUaZY5QaJY6mAIzMqx1xKUapd4p+NoC6J3FVOshjV
D9d0uvMA3ZJa2QralgIervWdfi3vqYNFRJsscJznJIX1U7EkoNo5FvE9es1VcvxQ
pUyvrG/RYz0bq7URblT3AaXCUeXTKOv0KWpqWd12k5JXiOB4aPsmgaHOXX+pz+4Y
hDYQ22GrDEhf7BA/95Y+dczwcXZGQxY+o3mzazrITfIMaofb2PH8uqvwEmtgG9i/
On/HL3pl/yB5C1B/2nDVrSgpMIqS9mfz8XRYNIIO6ui2MH37Qd4PzXGnIJ+nyWzv
iRQoeGBRYqxZDxOgZ9cqeWDD5aQ/5Tw4SqDrpmV4S//stWRFzPlbADBqKx+SxGf/
Gmhg66xNSvdV2qiGFgUo4Xd8tIfPlCilwVRLeXbekOPLjYDoN2lacOAmETnfjbos
5l85QR8HVctAEHXPg3dLFZRksuHncRuTlHnk9O3fVzF/Joc7auBaRGWOGmZuxWkG
xSzVB5a4JP15gM/JccCdmrc43jW9919E5DHePGoezfJ/WuiyssnvStrkeF71U0TQ
OrDfXpx4VRmiUqE+TFX5wju9uTkjr0jRBxyzHaY4NBvtq8BecnXtglZ883UO9PJp
EyohMpGpjZSpCXYExdnqEJt+KsOviVhFVnXw/y8sVmdy25sdpTFwWEUeb7A/sgEa
erGSJSCFKbe/ZLQWy6ogxOqTwTUFqabp6RU0iDhKDJgimQg35Tp7qE9oVlK69iiS
/t+wBzTdA1Vqqd2DC4ZvcW2cfp9SUAv1ka4fKA7d7xsOeTZie+fuHp388l24nZXj
cnk8PLPgmz3OF0WKgxaUnzfbReQxRmljW+Lf3T8FpkzvGt+fGy3BT88sbA45jwIQ
BsSu8TPm7Mk6KPaJEB44r5CCEPWBFzqFGoURszHXhz4pkycZmgRok9gVBm7204cc
DqCAi5B+E7WeKJ25D2KZh45uu4KYYRT8ZVpn+s0xAcdD2TfMmTIWM8WGVuWTKeFn
klU3ldnNdlmBQ8PIHnQBW8E8wZgvh3KFcBHwL/SU3kZyiERAvNLdwhNZlakdVOq+
5AtOpAF9XzGQAheuz4xurW+XxXS4xNbJLNs25Jn/Dptw2PlFk5lo0ZuvE+R0sqva
J2MfVNtq2vyuLiLBviEH48JJe9qP4m94IrFl18jgPlYt5ydjyhs4tnE22QquEOJ+
/Z1PY9xDgnHvagTvYKgL2d8zIlVDkt8Fmq8gSOJkwnM9Icq39qQTp1DaohRpyrjJ
Bqxeo5HeTuG8qLgqg4InqLY7H4TnCTbM0DhIkMDDbegf9pHH9GwjK5tLogpW6oTb
ZbtoORMDYcgu32kHntnyBc0qf5k9cQfMvwrwP/yQLvWoEoJKV+CHGBsA1/Aeu++G
7YAwwnDn6tdAMdivry6aFDlP6ZxIzPhMIDBql6MSzbwbd3BTcD0CUL9yf5fIBMa4
g2dz/WwcwDMX/qr0kqPrKhgBwhCRam3uwYo+KzdhyHl9USXzRgXIAZgi3xtZaR1h
nbbXG5ufk5ZQ+/04BEYioJqaITHVssIq1sRgICO+67595F73of6dCx93VK3+nYuE
KE6tk4zBzH/JeLY7vSDmfnIhb8TsZ5JheyszqkvVzrKbjRhsCg1YSjbEZ8GnlQFF
2ANkykRO35pb+rE/qbE4DufWaHI6EAfq5hbH9UuC/sVRtEv1Qls2wylimZbfbhdW
P06OdfP7PSUdSQfCipWCnAthqc0iocnu88LxhnaoAIsxiI/gMPdQ8P8WhKbYKFtD
3x7XVI41mYETJ0yvxgwHnq9LBVdYZBWoDU5+mbPHM9zBDISTxhW1XC9/RuVofgZz
uikbKAaMOFmANjRB739bFPZdwfTbttOuQBZXr6TLCPVabPswzTU9dYDUu47YZGHd
XbxYiAup43NA4x00gNu1qtD9pzHghr80kDllGg9htJG6GLcsVpyny+IHN2/AgIX8
Q+4/5MkQnoFdovqKqBI/xDpPfA5OYLVEzp6POFvo3Uh7/JG4dyVX7BXTnfzY6h6a
1qhMyD6hxstNx1Vr7xl10jpqP9R1czMEJLTZ9HeiQp+Di0vtN+e9dJ6/uDHdYbll
2AxZOJ9EN+IQCC7Mn99sIQDovBQc83/H4GHkMeUFRLOrSpdyOsu79owebjZCj1ap
30iP3UO1izbP3m24EsqSoebv+dMbfx1Acx+0jeVdNaXgJ+YrMcfaZl7G+bMYE0aU
YrDc26GN18bwQiBYydWQHmIrKulA3ZMNSJ5a7LGIiU/91S8oS4ILqB2sE//ATq8a
vZjln/YMr6YP/pvfCip8rbfw4LRyB2TYhBB8RlFMflGwRSZNy7BtBHvAJJw5Nqq2
uFjJvQX42LyuViSSUFaligHxDn5cORKLFKl9BN+SLCac1PVbB7pFQRg7gLIOWjyI
hkC6z5TbNtl3fWM/BaVH+orHG5wII/c0j4GvDETIuAZrgHxQbSTbioToNGcKsu8D
NO+5RM0FgEH/0+fWMv54iEVXF0YFzr3AP7A7QVrZjXM56Pdz0jscwnlt0I+uDBmr
egzhqhVIadkN+xty0OoMN4zAwKQx1Yn2EXta0KPMeMHMZ5Tqv3XtaqCWM73OHveX
bmJizMzRYAwgGE8yjf+cLIkuOIOAveSmPSX5xVtN0LmiUtYt+X3Ey5qddd+2nH37
Ca/815cPg+NZmQA96UufG5UjQ1FQZmVX4BesmY2Pd/KN82bNp61TIB1YK8rwulIL
pQv525W/hy2hdbI2ce6Y/aQ+GZX3+9hDsm6+CJ0hD9uPP0C537p7XgIZ1+XoHJKp
QM4Z+s98RANGCJ2gdDDNRn0q2oOJXrqdudFRuI7UGOG+m4ILrF2IMM9EBvXGxY2g
vsHUf1ogdB8kkRweSSreaYvDl6yXJmtpirVpY9+G0rzpKPpw9p2mxZ6r6s6lxq85
wuaO5tdaqDISXXTzpZ8RRpOYeLXoV53BCnykezzB1FbgBOZ55OytqMcb8VBEM+O/
Fs0qhBNzFuDGihQvXHjB7b2LGWrFwGYW05RROwnC33KN4kEcqBb+dXtS9x+m/vIi
BgMK7/TuAzdvVIWCovuXwwFkFn32XG0hS0iOOiB0dt+v/9e4idmEM6IXQfc9icrL
KVaeyGyuBU8Ovz8LOCkMyX/qqI68YDrZYd8KcgV8Hm+AVtnHRiF76lFaoduI6l0G
99JCEcoooP4mHIe+HPbGTnLcDKp7/8jxjGDexFXVWQ29blxq964OQUlLmrH3/FKj
iBljsEY5rWrxp58efOn81EyhLoovNuIJXJuOXLXE25eVr/v5wjix4IlumO3NPWey
8YglWGq7JbsGo1WPaysnnyqbtOYKQalhoI1ZQsCPErowwnhS1N4bYR1/i9gv6uBs
Fx+0137vj4nVrYlREx7fzE1619vY2RUyRAglwmsyRA4Jvk/O7fH3O7yPeJ6iK5+h
BMV/fuQnoz38qjXkO/+GtJMDlfpKbd93D4Dnz3QAYNaf93oqPl5WV8NdyA2Wpm68
oVHORe/p9PI/XTj+Qi9DHrCCQbDOl0zhSMzbx+4ruUr69ZPDTZmCQIeC5UN/N+oo
yiNUXM8PgOZceerrNVpJFNyQr0YErSOhGN5F+HEz1cr7CGQvCTlULk91xglzvWNS
p/mHFzYY9yfg8GnYsVqGk0jgXxIzRcBpW0DQbjvio+GZFthDZBdIOaLvDFzR28IN
WWyHjaaHR6mq8BOvwb60GeyDlAMJ1WdiScyRXl91aRFGNiqzA5kM9BC8s5XEEvym
pqPxwD7VFx6LNL4SuIZNkklKMILd3EV4jjpVLeCiU4tqIPb9ivlm6mL4oyg1ri71
ZbaCqO278z7QlX+swAwX1lcFOSwjN06U3OVDxPoVwmkQYhMJeRBE3h/+W0yS5gSt
cg6KVJRhpMTXD01ci/g0/ZS9FAIIe2XAcJqycGxYd8JCX8Wv5+jIbbdkMFCR4uwc
ijL2eg6/I7G7CEIF6RGiCmoSyqxS5Lg3FJjPTQi0FgGjMa8lI4Tgx4EIIsysFC7u
qgVuE6YB5h1LrBFD6SyJwbWMCFtGQNv9LIK9s0ixDHJhx9XvdILEFnK0ktJH4QRq
4Lqjoyi94Jth80+TuNDwXgLG12zw2kHAi3y1bdNNcTZ+9jq13z5EK31z7DmCoarV
5GsUzMk/+9vJS4gS09it7+hBJMeJnrWpFXAnG5Rh3cykwOuJo+r/UHoBJ1usdfVU
cQiXDXr0rokXi2VdRGVwxM9nxV4G0Qi76/URB4q9TZIzNxgiX+G7enPhcEx/Wccr
jiY5atVgtdJPtccDjIMlTllkL4IBbLTW7rwT/1+/HAd9JdE48+aLFD8Nhozrbusx
kE6nMMf5RIAWqjqk4gcjCjuW05yw6UMf0S1poHI+Ug7aBNE3gC820K7kZs8O5yKq
hHQHgzN44PdjGt6oskYfWXl3pcotd8S0cQKqzX6JTZ9m8LD9eM3SWi8esI9qUlAa
K/NFvesZ32Oqz8WEObSnjkoghUu6NZhOw9AiISuuBpvvHL+MvzOMv8d/AyftVIX0
tRBWWahqYg8scphbuOiyrmM1yHOU5HZq5COkwUpeC6Sm09W/9igO1tQdfYFK0CNi
6oeE2VtT/7jMJYJ98zPTVBLJW4jBwS3iSzwsNQRS5N3F6vRN/ScV6Mh3UALG4C7O
6xRvem4bQYRTg4qzhh4XrSZYmFSKPFgob/nGNwUzmy3o/QSFQeISYy/bzAhaCN5Q
hu7Wuk3CS7j+FPmMP0aHD26imqPZFCHEp3bW7xTk9ctskyPykuw48lXha82+tl0v
odkATXZh+TvRpGF4DX4sE8HFZndEtQTcVTsTBmfFthN5RcO2l/zDrs+NZNJ/LvlI
DevJgtYa/V1UcR7nLgsUi4c9393dC6CCnv3kZNEOh4fWTNqIDBmAyAS7K/bR4o9z
alb/IwAogm27sZzi1HDTnx/SkGsCCpt5KB1akF1TY2SvVylflnG5B3XACHG6ac7g
TOOf+WLDQ3P7a4t7ijBSSCT99rM3BBJQ0Emv2JoBEYSmGDL2jX8iR8WaFN/CTfCS
KkqPbPIsGK0fjEYlVkBpU8QE8SNHZ15KWb16buGXZHCN1zJw6kbvwR5//wUt0ipd
hREiwDR00m8p/GGZT1nWT5m5w4bYdny90OY4qsUVRmk9kmUQM89zVmaOheATgwsW
jvK54cEmuYIhrA5QQjYZCz+1poE1grNmG6rzArVCgXoVl9bGjLgFZ5dIc4UwvcVF
WjYGhXODtEiEmI0YeRJ1CQj1VDv9y/KMdMOQ/b4rSIH9hzTpiMDpvTzC5fVE5fMT
yQ852bYHQSukrpI6kevh2lCGpjL38JRzRhqgI0uQ2gaVwwIIhEUMMqnVb4X7pgWK
9W52N9G4Hp5ut74DK7Bl9PdGU7kJT5tkm6d+Ud66k5KB+T+1Z2aHs98nFpPq8pp9
aUaqY2H0zWYWg9NcYisgffj/XOJQVPDO6yOh0PFIBL4UK4t3B9RGI924tnb5azvt
okSrTbcqXwSN2pD+at9gJhKrt+ujEE+VuCO7EilSFh6/DTdjKH5v7PyERgmOrTUc
grrxx/MNUd7yW7d8mvHXxKqrQXO8tNS0MojUMgN2ETwQhmAWUpEZVTQxePHWPyPO
r71fC7cvkWc96z8jrjuUpwjRGigCBtyLjBmY/hNu7VHuKY1JIKEuJR6vE/7ytjYk
LbhYK+ZcyM6qjCa+hqkslECPasH1JMpx0I5wnmNT4bIf0XdEk7ZxIkFTHKOloM6h
8wwS23pQAPKVHMzjbdQyoyKpgzR101RL64JFyAS3fw7bn5u5W1jCv2KP5e0C40fS
5q+tLXQWvzm392nIUfDY/K9xNzRa9QtEI5Y8CKUdJllbK4QmtxXyu803E8r1fPMS
KNUaYXE4R3Tp1+8hO7apTwcHNtwoO8lR/w8SHnsqHy/+2hiOXEBn2q8qA7OzW/IJ
xp4/Dpye/oX6MP8SDSbwZ/dR5x2RLkJUMbDATBCiZI6YUzM2GJnDFCgkBA94WuVZ
z3b95jY5OdamtN7ZwDWtlY2mBPlUX8E8ijb9FAq76nXkeDJhpGOkSUbTjdWt06eb
ub3jyeL7tNwAqj5Q4VHP2t9bHnWKcixRLRfTn33byldOb1vfkdRmg3Vlf4QoA2Q/
aiYoFPx4SaWZ1sRRpP3HhdXk54kDxtytE47KZOJkDiwtXo+esfZDSWQO02xIU/1u
Ipxxw5kAGWFTAb/NllOF3OYCDby7z9/7ykcjeKiCXuvA2ODpU3RhkmJEUS1XMMJ+
3dE7ovUv7q5cKmWtvNVrMfV4BRhMTbFwgu4p7oVxN0Xg9sQ4AgwkQUga/XvUAC5u
+bOckmWY+5aZ+ngfkr5mPGzLNDu92WK5LF0tXbtq1eTFBUW8xilBR2zrFsBLpDfc
XJ0M2vUQtRtted20j+L8sPwU0wnfRbmvaXbPY+DzRg1uWe13WG5Bs21Vx9yqOqLo
55zOkOgI/x9gmG2/Klwx2dXrEfeHTMjctAEMfRyPGV2KtsxJX/tn8HF8RFjksr9w
8pPEE5Vql9fnjz6+YP5VEmV7f2CxibDa//eEtcJ1aG4IeJ1eblqWIhBJXF8dXG19
P8NnwSQZefVNnFh7B0SJaXHAWflO+dkhj7dt3DhwnP8PBvGsvui62IV3eZPQop8E
UiSuzFXCwju3MHYdJYBllj52s+1fYYLxHH1fnbwQOIMaf61qMs28FjmB0EcLnKje
QO22KFe8vsmFGRZQoxn00J/2iczWiuDRy24Y76dN25zNd1GV4RMdBiEmTJwcBMcv
HiOEfW2RmHj2Q5WaAjpVbbN2tkXOmbhxRQkuVL3fcDSTfsYXBRXNWYZMIoh7moBj
ZysOcawq8ht+hHnJJ4cU16aFHoI/e2HuOF++02wbdPT83Oeq84t5cr+uV8TTxi9J
WpYdpJKx5aYyZdSoeHCzAYnUdqaT05nngxoyBUPYBsOxc5RkxA4DAOP87EoFkgHa
MG9flDzVHU4Sfr6WqiSPWmKL+DVlKdSaG+FOf8BLsjgEEMROPDZAYaO+ZtKHuktt
MmUJZLby0yRI6O0Hkw/VI0tgGu1JAPpswv11DIjsUlAAFNxiir3eWuXSrCYTynvP
5/gnkkrLkvcbwPN70VhBIX5uOZJaSy4F+Y8WbQw5NF6kNUKipGuOsqc2FMMn40KR
l07YCA14k3sGS8akL6QFEXuZsXvnHqhwAFjyDRd2wMNGbEwcsEW4/9mxou1j65QG
5ShCIoe2VqENOtGnjsZ/l393bnNpRNVELz5KVQvIjsio1qhXqx0WLocDiXb2RNtu
JRIkj+5Mk9i3ntrfosp8idr6dxstUL83s8k3NUFIZ6F0LDaoi6Q9D7FffUOiMHLM
JJGYwZXfMa6AdLuZfEWwBB5mSQhX1X5kUyzYWQl1jWSr6dVRkIuyObNrnyJ/XMnu
fLg/3Vt3znp9lTGYQE9cLXbwI0/InZEioZE1p+jKrubfFkjRzjcs2d4I3Fx8tKJi
HE13CwVu6vnvbsyj0VFoLfxC0A+xmbTxQfCaZTlbpyyCWUlnmGG+v84T0L7ObvlG
+qfyp739eUtIQaBOP5ygmVK3xy1CPcPne4JQQi1/z69SogP0MolpVhbCgZWSDcI8
+Kh58AnpmnRFw+kO4Re4Z5RUqZvR30bGHjVY+6E2pLVhrAcBEC5ture2dD/+Tlvj
9kGaASwLhSXbbLDWyyjbdowwY/Gwm6DQ6p0aKtZZAswVqgV/6Xhr1lLXk8v7vAQn
kF25cN37ynw+pCOry4BTzn9WwHkDkKLebTOMyTGDa6dCqfLIDyO4DEOzoG99YGgB
Xn48OCk+WnVVwS0zVBIy54GOpyf/F5Ha1+wkurDcza8i+Y54E94Oy2J5d+scGgek
Ih9hv513OmeVUZPXgbNWtb3TQjldsC2mP7gDbIkZSrL9eQVRQFYotr5erWBk64RO
nxhPqMsNmBCisjSD3vYXtTB4QTSi6acbDI4bkIPEIAGTW12/cHWGpNcw+2WaPCMm
0dvBYjvjHzqHInuUulfZVG4SY2YqdiojDeAMb8svd6avlZ4D2t0BIW1OBv4ec3Vi
wjAly5YaP0vTIu2kFo9XDVcCCfvFsfIpBMWeT4Sl3haxb+YJCJyhe0fiwoypBAhM
xceTFSk7j2khCy4acZnzdmxllRupSKaQ/MMSgroxRrHnhwbPYccpbxza8WEH1HKI
p6bb5zz/gAx3eNs4iYEUP73dM4zufIpFtDbPtWrlkc9kZUEBfiqgHFVFmDDPKkJP
kT4KgrpRuk1ybxBYsToeuBMOos5JqfvK8ujH/hqtX9O27GOdc1jNPv/ibJ+BMj1Y
qlhCiB3b6eWppFWqAH2QIwuxGgs+02L3OqNonR7rwwu51cs2krjCQ3tOpXXdHqFU
+vyc9F62Dla2PxeZ9va02oUVnHZI1tMmkN+SlrJyqEo/x2/UQ6AgQCb2wL01xNxr
53mh8ClhLjixBHAnwsnGcpeHdbVVXgE3B4rM48eBsobPSjHsdFy0Px0/Io2K/FjK
P4MUvS4qV1xQEBeJXyq4KCy9EgVSWS4502MfTJ7QjZoqsPMQ60YkEFIcJtdnpDHR
f2Bc6/24ApAoF7/iRGci4ZkNSCqJBPZqBhXZSYWpPiGgV/J20UA/rFJwh2la4BgS
7SCAEMaU76/lcyD83zgWCwSlauxIrBtxhCZOofXuiowyc1+wD61KMRgERTu5hx8O
cf5SNln8vu+6xsx31QWjVIftO/cz7njgYtWg4/Gx63BuGupEMEn+wU5KfAdwzKAa
j/i+N9KtO4KmgqRxuRHGsm0eIriwqwITVf7h2Z1fKoTt25cMeNe+IuVn/atW6Sdm
pYTyz5kfuaq9+2N9s4xpCZf4joC5nCOlyqTAsFCVaR8FcotgZAbVe6z3FdIRLVMg
FfwHT4S917Eoexu7t3Jr+cI8hcjQbcjkkasuFjM1yRFAHTbnxSd5ihvZDqkPWogq
ucnuT5uYlz6Mxt8nnnPkBvBBM0J/GjIVKGqhDYFVPZMbODEpUv5Z6cReSBTzHKew
VBdSLkJGSXHWHzPbXcyVb4yhHI+VRLEBQtuqvUgqI8AddsglvDuFM9gAJ9e8Io/p
MWDtJk2C5fIX3zW7iOQot2dOr3AafubmO6r4pKNsdlBfbxOH7yCRvjV9qgR1FTfw
djcrpGxOc5yJH2ZqtZ2ePyOR5ZjUWfNufX0FXHEbhPZWDiPJsBmt7oT1ZQMQHrSw
BB36NRs1Tt0DbFPzPSrK6iSoKqQ9Dm/X3UTTqaaH74H5pIrpp71H273UqzlMrViG
1qa6OmAGg8/6+h1GMUzcKAHHJ8Ora+ya4g0h0e1sPdnK+xrajU1S+Ze6sADbo+t1
F6XWWYpePyLC2fp9vPXnS+CeUm2vOaIysWxkRI8EHhhkOvjml9cfJSBoSjYygT2d
8LOnXFV6qk/xq8SIQ3VRf1sA5CcoOBGdDwatVicpE9VgQflH0STVarEvufMsx9Be
NtYRRfz8iFmxHvR6gwTeZ2F6O7X96PlkQTjKAniatVON/RPrnBO7lUa4HK/Jrm+6
0/M7dC+j8nC4ao7qsuy9ixRjJdf6sheD0OpOOvt+Ovbn5UDbKG40llcPpr6YycAM
IsrC0K/IkArrx5bxJ8j4EaNNtGFy/wCbH16zIYpdNYaGbl/8KzNpP3J+HFCfZirk
zLqsBWq6zf5iPn0SLakO5DBpElt9L5jH7sTAwWwTvXrjcxQfhnnHlbIQr1ZYsxrF
LcS6x49Xlqv5wIHtNyRwh+08JDudrdpNWzdGUp+7nIESltHSzmwfP1pzJu2T6Q4o
OoixThdG4jH/Vl3XgvUSc6Yn1fQfqTPjOqeb8ft8gcsLd9zeSuI0Fr4H7ZYBM+YP
TdzE6QS96Qyf2Sn3Q/mVvDeJAJ/RvRLWwvr1SvW8uOLpfuRTstf0WeOOZuZuj2FK
HqBxNEY8mwJzDd+wSd0VAMSXPWDXXddInr6kwt54k8VakWAKZ3eliLFsFltlOdgv
1Uv9hio0GAXbVW4dW2S6j1EBK7q9GEo5DbxbbU/5XzFFsoOHkg9TmVYrrNBoxn5G
YMEwDzlBNBKtkHYXR7n0CRGBVyeRbogMlF5a3gYHADbIPTEcdlGtWm3GXPxp/vAF
cZh1A6LYXUE23hnM2j9qILdrhH8O4MAGvJTcXceWOIvxbTDIM2MNnKKoxaaz8iIo
PRnmBknJE1+npwwU4+2vcAzdo2HOdNd1gJlvnvzf3/ixMfJFWC5MymbPkApCwlHz
6vHnuvokwHy/T0kqed1FoyukiaQsfyoOhEvdImvjYNYIQHBzeRQpRhQLC5YM+Lzu
05cpdjY6UwL++N4tJbRzUb3UXJYDPBUcbG/XeH7dUx3O7xnq0ZCWzuY23sYd8qFV
3Nz+/7bTeNgRjIqGTiNbG+LQe+L3rGyuM973SDvYF24YIsJLvdaKfJjzN0OBWzEt
m7u8UgD/q+omRX2JNPzUrurhIQ1iJE0k4084rEHUdR8I2q/MENbiV3hPZDklAM00
8uiifshh8VGuvSy4a4CBBt77akLAgUoajBMVQTAq9yvzaXLMLGk8Z7eocnwUU3Kq
VmZTAykSgoZD6gGHNTVVueI+bhLkXt+Otl8OlMX7Xw4kq9QuCXovFMInB2aXLtrg
caxqKu2XNHBPSD1knwkfK6mdus5yZ7IUXdcYbOGKYjlvy8AiEoljwf+F4de19bRn
AVAhveZCCXAddXi1Z4yvOZTSUEKbnF9ecxJbqeTuuX6wWxHBFLOldtgjfCunqI5z
sI9m9Dcopu39pZZzQUL4wqOVuzGLEyLYYwOlI7/wWppgZ0tfZ+G/CdhUqhDj49X7
2EAbcO7OSOMsw4m9JvWmjyBDrr3YPEtj3gj/RmbArB6Igoyb7AP13i46Bfkd+Ya/
ZotmRGRIGM/7gEy6iGsEvTwq0TrX+LD0RyevRoGpudozWX3KK2ODu8b7gW1qb6Rv
JsM+17jAymYAZd7+BEe4X3pAeGZiOMJnPJyqth5F411ddGll3he35dQc6zBcIyhH
Ro4cDKi2bH1Ziyxf+4zcsnfFnZjE/tmMn5lmzL6outhau8xYRau35UKOdxh62VMb
d7OwXH9FhkFrXAa9cZXxq7SKHFqiV4KUu0hMfE0uXClejStW/6dnM5ZYU4YEPh09
YAuE/37QRAu0PfN/KxhSwRIx4oVONIKUlMXVgEQj+CwtVSx0sJnuHxpztVDpzupR
b8arh2o3tiNXvIrJDKck1C6GOQF8rncWpJ1iG28m5DDKIpojUISrtLwRN69Yi5f8
lGrnmH8o5OsvRcH7JOmt3Uw/c2UwOl/b81j9Xzjudiuv5KyRTMfgmhXOYPqnD5kF
BmZsy8oqYibKLIPSOlwqYNClqNhvJmpuv7rE1oqqKCDF/bvr46fT+IoRdMLnrXKk
ySjBk+5v73LluXnoCR/uCHOutsyREw3o3WoHKVPlmui+C7ZEqUmgaoidPEdOt+Wd
ROKIpVg+qoOIjgJLJF7Dm5vjXvoEV5YPgtVEkTp8KNfuNsYTG5wfTMKvMnd7JV/0
fKURCDzjV5+A4e1G/NldlojbP/WNIutnoYldn6X6XCvtv3jPW38vSJNwuatl1bIZ
whWr8jwrJlvd7yyg6JmsnJGu8oClx3COJg9xwDRK/u0Xrp65/H8juKbzMpNqBSbl
hB9Q7lR7TzPPE/GgPydVFL1944ZGXJAXPQsB3E7VdRxpWMc162p8/mRfWTcuMj0K
Ef4lA27l5X9Bc3IxmGc5Gx5EZxEvQB+ZxOBsee9wcY5g3rupjGuba1QDmRrOyH/r
k+qiTx+2OuUf+QUzsFbUZ4sL2c/Rdo2193AobPbf0jNtL4tZsmEhkjOZyBKbfR+Y
e1z2axVKIvRFsiVUgELewmiiNsFMDjFUZIDKki939+oBtqR7BDGnSCD4m+zDD6O0
2KQYUnYldoIIzPOP6ztdGFC0V/0CCs5i3Sj9v/vHHJPtHfZ7TpCsMXFylzRM0lZa
k1EwPbicvr7eRqhDG9tskvWCM6fGgJfEnXqFExNjc+DaLba8cqj8Bb/vF2pC21mO
ui2tQoDU5x4Jalujl93/zYKKUfHJYAS05tlQIttqyEUK+cWyCugIwL/pBIM0/qjq
SldvnOn4+XanvN2PCqSDQHKj0rPBAVLB8/GmEv6pglhRusN+g7xno6Khp33P7zIa
cEkYlugbZor+56VB03HgiasKETPiFZ9J40GG80bROM0ceYmZ/7GGL7pt9QUvQgsZ
Ji8HqqiSJCDAT/+cnZiH7ZsEoMw4Pi4xCISh2mV50SLizdUXvQiU6V8tIMpv0ub3
R3T9Mc2p+UqH9ZMyThOItSOYEC+pdaagWAika4dmoZjOyE2EKGEkJfhYOfWFhj/e
BkWgsHW5sbA3JyA5D/4EEZiFC7v+YXFTFQo6TewlscicdjT9d2y2f45nQUTN4cpG
LTMt93fKk/Qt6DFbFcLZNptYXUjJmXzN7d3fenHStCWCKZePqrAHWmSsZqMRfF9Y
wdvJeZwIug3ec7nOFnaIiptO8UN8oey4E4CuDXQO0bzkzlXN/SRi+kbt9/2zWYBj
5qktsPJuWoTm1QETgSWr0JM7x+538TkB/j1uu6RUa3Kijtk9rQGY8x4Mn+s1x/de
HhdDps0PAbdWdjbIfxyVXn0Bsv+lhBZIA3NH40GNmN2qa1lHMT8JPvZFJov6WsBz
6RPzg4ivHZoBA18L4w6xSLSmio5SllIzG4Kct7WoK4wHWAFjabcERW0GlTZcAX8Q
0W7/0nVDKorp89SuzzHIzcNxFBlrd/nq50HnNjvGBXOWCGgHuxpG61vrYzbpTGk4
XL0PJ5pPhTev0p8vBy4A/qpHR2OzWDPULTNp/5UjbJH1Trz5SSSxB9apemvkreOG
/Tvt9TuTfC23UPI9KnOhDZe9ZEvj0vQpLEGM933IYL/hDjYuptNEQwLjj/MfqQG3
TUe3U/gK9XsuNYiuBXbb5IWa4ujA8N8sa7/1TFztEgvSEzt8ZxUfodkE05LvDaa+
Jm+fJf5Bn2gbz5LLupXECpZFuAOFt15VsEAdcwEaZo2hbsHBkWXPfHyr8viK/UKh
oLKG/tpz8H6q3DyWBWuxbUy7jZRGMQZTymD6ZnWMXKmdMyuwhlvnl5TP+cUlTPRo
AE2F3L+bFmH7vVhIbf69XvMGvko/SthVA+1cYcC9jgTI+JtyhVmwJQMfoTAwJWHB
BXWB6fKPCGqIuOgLF1muRENeaXuWcJudogHGElzZnrode33o2Cs5CMgPNwLTN5ef
Lxsj8YqpHgmv4gI4Syt3SIJ2az8QLypjQMTo0QUmFxqKP4f6KrXafEf7mE3mTQXj
Itu/5P341yLqkYhF3JerEp0lkGiEvqG/Y7ZHmPotR1Br89d9zqEDndUK8TIAkM19
Y8VF85plwYA36jChnMVuchJIII+QL1Rv1SeWTW+pv3+xSUd0G4HpcFebnVDTDzfj
yXjBLdzjBKv/7RWiZZUBDWoLXZThU50cjn0JzGmDG655/wLsg2pYpc6//2mWDdWn
Cwc/6fUY3MuAfp0aHCnU2saoeLmZuY1HtqFmBiHUo6niwhDmcKvHTFIWXxx7tBOs
CPVgihb6wJVUXRwG5h05WNLSE76IsKSpxpmtEQ1Y/zDxxH3K+6TNmouas0sJfpcr
ovNiF4qOb6u6s+BZiWuiUdbStMqtqheZ/YRfqekyIrFMSki9PCSHt44p71eBqj4K
kvGbptcMC1Bm4OwENwHqhkBr7P/F1gH3FZ8VGkUd6Kzcg0lXwb52CJktAELHUfWE
T01Ls+Sj7ZfznKQXcZqkHKFPFX0SCK+1jAd2Onhtjnl1p8CniHPMur/6s1KGuE3A
IYW5lge1lpLmZUysmXYKu7XSKw9hGpCi1P6vbMlA5tXNRM/nPH2PuF1w+qCcKJFh
FxqVqKLqn+4F4UfIEU6toWOXI9FGzrHLrf3Ohwgxew1EG6XjjmEXvGvturBtU2vJ
2aCPNAflV/Ia+d1c4kEqrBkuzHf6oWu5uOvH6VEP51amaPdfyC5xm00R7roZ77aY
6XhtAJIIAR7n6xAFdPbftZE1IM98QE9D0LegCDf2ihNAqWFbBde5wIDe2J7S52v5
XhddcnMiBh9VmLaEvI54RuBgApH5ekbZF2Q5dtFR3HkfqKdusnMilgh/XPZYSAV1
6ONoDDNbuZ73oWXtrnaWAdnr4JG1FYUGVLiJUp9VL5U52wmfe9rZDHaZKcLkpmeQ
6EAI35q1xlZPjwGIvSNEN1KVrUTSc1BHJpMOGNqX0Urvaf1CjN6fBApIPoP21yNi
U3cfGqtCwvHhmxadBmH9m6NQl8o8fZlkQNBuqn2+vd8a5Xald5s2bTYmSsSKiiPi
8mMl2ZhT0OiBkoCBolmiR79y31kF0Hy+cNZ9DUfmGU19RDHUTDI7qkE7VaKiwE/7
fddGqEev0WnsF7xscUtQ7izHEW6ftK2EW27f2F08xWentlRHYGw2FaFUUTCgoXxH
AbzP8M1dC72kBd+qfq5fS05GgZedFwHB3XGFoulkYdtTeAlAieROBCgEPYJ9+Ddk
8mXtlqOagwRSmF3VXjmQJHhsfWMJw5Gh4gI4eNRxxDQ4gmS9mq6ByOaPZIdhV6Is
crN2rMK43z1tB23+7LejB0z2ii5h0vW4xhOXCWC50WVNnZZgIEfjoMKiI096JCkC
8IFpnUaBQ9Lb5u/9Xkp03LRx+jPUVMYo8kZj9tpCnorqhpGeQo/ee5AMqCH7r4d/
XSq6HNStK/7F/ENm7UBL2iLyiS7aK0ZJxMhtArkrMv/ygb0VqMDwKdckiWuyPehj
te9PVYqb/0gCvq5fOUsDxJwtNwg80+ZFh7aGWuQyrDtdHGq51hV3qwpWIyzMCtHU
iGWYM9V7artiwrt9NF91g51DN5wNWG4UaYRNPq9UFulWyh4Z1Z4NOoFpXxcfmJcL
2qzwFi6kCAaNOh6GHhqsGF+Hd2ypxzKa2T8uuDWFVCAwLTpWPjfWeQOgs/SP4NRG
/q83MBQeKzclxtA7Y3gPH1lPS3R92Cvdp5+LHeUkJ0kmK/9JXw3tiGv1DMZ/PZNq
zJRLGuC1JOITYTA8r1nJqvBnI2klIBdOTJAfO6peIJQNWwr4cKThL2DLIY5GErzH
nJLg+BsnOQPLhKmcnB1mS1Vwvy4/w77bk9FnRwQT7rL5JvzsGzC8D1w8xGDYoJfk
Y7TEk3ZyfzHD4E7IfLVl/ZYvxxbwOxFsiqAyPQnEMNv4f6RB+kGc2UCT4WTPJVz/
Afa2CEdosRXcI6Nsz3JjpWQVuE0x+4pvOXkDk+jkKvdD1eeuPT+IOoOgCiiOhcpr
7BomFOq7WUzFHMciXBbIM1KaW3F++bgJZQFghEx4KgRRGNU+MMf90Bd1leCUXC7s
5bptVqPxvf/XNfu8nZQAAe3rFrrBlYOPqFShovRUhudjhyrjtX9My3Y38Uf0rRJ7
nPmnt6nCurx4kU9RcGfhO6PoMMoWgIQ1Mv/0VQKvB+MnhHMOSxAHwQo50hhygh0s
vYdcYQgMHqLbNjJiEqkPg+c8l8ZS3uNae8r6LUeSQ5tUEebyJ2hZuhIUVy+9krEP
eyRERVJ//UJ283uH+9huSY9RIi5rgTnzbbNPMUHp+/S+yHCipaM/a6V0bkhOYhbO
xEUS1WdLhAkvvcAK+Rnyu1XCOSiDnfDWGEL1VC/9jE0XsrguDgvcvYLlBNTCHluG
MpJiFI4krg9nga9rjqH1W4nOZIY4PNlcakwCpLx/cxgueZpYyPQn7+9p4ESA2X9a
Lh04X0kfrxSf94IaN3N0qE117wYKvp+gncE5rEH+b9l+clcayU+7A+5FwCykyWVB
NOVENz4BOSZcv8UCpQ8PI4ThSTDAXo5bqW7CKcz6+IuD+GU8Cf4hgxs0ThYR7KWS
5COKblV6yyznuQjayHQhaypRd0f9ncUbGe9GfPGMpaY2uCEd87h4Nn92ZJQ/BOM8
fmX/uIXVAJHHI+ub4FlMz3SKi803e/QVJiGogz0Jii9ErRe/mJiNYatJR3INKNVk
MxavQSm2NtZw3/Iu4/3CIr9V+/yW2McuSEN089JwHYJScQTnwGM/24QuGTyi4owv
NCSHbBID//RCJLW9EVluHqGLjEp3JsG724+C5WbaiNpImEbCFELghzykUgLSTmvm
KU8k8z8JzZNgNMGve1kSzgxENWcu4eR+M4kH3G2Dq3gigh8pkF6XHUPGOPrDkABF
Wekm8bvnWdDN3NjUQ6fBeSUT8SjUQ/AW+7wTCtveAxrvRKyOWpKzVZrX1cWKFen+
17vuPTeGjbkw6yeZNNwiproeFKaHSrp1nvZ8GZCnviDczyEkWJDoBOcp1LRZqR8Y
aQyWL3qcjbqV5KyPeFQcljT04/PnCuAYKfyForz5doDjZo0hNJj8P0Cb0z/vMWRI
WKfn8BB97zBSWBu6KQFcqoIX8JUDG/M8WmHt/IONGMTiyxlHu2k/9O62mvt104SM
CVq8CKKtu3KKyvWQI0vtZ7ATaGtmljLKa2lZ3z2tGYZ/ibJ3mioISGjOjqP51/j6
FjFEzfw6XrJfGJomoXWnEWRuxIVZC0DbAbLjFh4k3GuEey/RSUlP39zm0Mj5eShF
Nwnne8wAAtP7NP0iiWAs1zvzBeqYio1/AisbJwiATuDjxKarPKgF3z5KNgqfZ+ky
TOb7s97+GoWWCpmDwFoAOTN8DneBtCo84Ir+/Egm58AmF2LqOrYTmRZw4AaaV139
h50mZSQDtw1UgfSj6gywnXrM9CYhHXjC7Cl0sKq4uLpPpesSjNq4oPGLerMNoGak
RsxzwX/mS0YjWbglOzGzc5yofptV7qr1b2ZRtUWPURJhg3b1krRhCW0sZ7Isxco1
BUBi3vpS0m96K3TuJH18Nxd5dqtsgwMZtldg//SwXmYUXUg399IiWZZaX+DXIL+n
6wxOoa+yBk6DUurVTyiMIuF6pHZaQPn2Va0aRu4DjHlAdQXq3sdyuHeCzhxYMcQY
BXmLIx9mIOVnfanoqTUaJgC3LjdKZqec8Y+JY2RZwsds1CPyd3QC3oyM/hbLV5QO
fxIqUroNGcYzwdL2anBVRhFdpUeP54SKRORhDjE+cmLb+jaAMT+vML6pZAtpkdjC
iTqSqVgD9lSYX5x6vZIl6a+spC1Q6HVJa5cbLQDFcJfxkGckQ4oj8fkYQcAWTGJ8
OW3AWVjGoX/3R3M/rJZ/HmR6hGm6OhC9bWDJ3Q3PVagTpAcGBqwE5doQTBGC3mej
QxEtLKZltnIhlTXOqOtIjZ8fJ6zByY/c8YpDY997ttHWUQbqf3LBH1h3Iq1ZpsEr
Cvw7BlulETG4Sjeziyzaef2xyJE7TGTDcmE7ePX2UoR/M4EnbFlOTExhsg8mQbdO
VZ+Kz/DF67YduoqpmGH8z8FdiVHkvGGoAyu1s4eT8GExJJ+N71PAq0Sz4ggBD8CM
dEhv4Fef9WLh/x6fKrU3+2RZj9KX0ZkrVjydn3n6rb3PwTXOrWxZWCdmVN0A6cK4
To5almP7p2ps9bHzyUEn4jzZynJSx9c2SBnJV4Eb9BKmEI1HnHSoP7l3Uf+c+nRA
LzQd8ss9EAu1S8H8cUMloR0HCmvUeHo1d67psIENtGXaW1vpq6XVXdoCvh+v3wl3
QMqZqAlHIPU3LAKWU56Da9epW3g6L2f0NkM/dVn0h0LoZsQYko2gKTQ3ry0JK3MM
LHzMfx4PaomOmyzdpUVn0NTffAJdjLBu/fhHwl9p7rwFqDlYKDm91SIHiHaydWYd
2W8BOsc6PrjiZZLA220UXSdO+o5EYC/K/mWSlNOJ/QKIPCHdAAYLuwxvnh+hDQpl
pd10JmTTIg1BmK/bgx0Zp/ujMwk6YymLl0XiwVg1Xie0N4foAWG6J+Bmob3PPy6T
xO8dbzPJvjTgcBHMf0iQRmcJtU9r2BN9+F+lzHvpTxoPcqPEFQQCAXHgQVVnNQQz
J2ajohnPriM+TZBCL7UKHJg2aLBcLCtPDy68AhGgxS+5fCDUKzbXAu5zvvhekKsi
00Az0pslguDYs3CowDz4moFlOSLhv1rSMauQ6l0NvRhPn63BoL2EBIA2Mx2j4gfc
PruLuR8x+2y9bnXokgB2Pvy+aViytPXDKO/tutsB1KusbIEsaG2a/TCZXvgVUWC4
l21MrBMbRtYGOFb7a9B1om/gGV0wfNjoh5zc++a4khDaH6S+yUSrPIVwC0BAT3Et
DT+BEjth3RX/FHJLIXIFvuWEQEkI8XDVRmLrkq0zNDOeSgM1SYBUbVpBPmt63xUZ
bmjFhRN0ZauDxqXoprAKEvRuK3lbtD3P/NevJ7WLfPgcQAySBRTuWFwGAs2GI1p3
xm3bDcTuITH7sVshI1CGOtDRLSLLNuph9HZOiEjFWwN0TbzxglJG3a1uOrQbMvNT
kmjkqrA+wI3GxV5rgO7iZITK5RMXZ1C51LUeie9GaD6ByDSGfDfJ4tgVYe+3PR6Y
iLHp463oFNgLv2BMaFpCr7K5Lys82C3oBN9VUbCDufWU9IlhNkZ1RMLTPa7JmaX5
qHx+/UvXVOl5kN2TBYwmeKK3gjjmfQ+x4Kc0seqsT7YkZSw06ODAoa2EWUya+XoP
OgGgFWh8fek8rLoXJHHRwV6PqPS2pADulP46kOjWKc1CnjatigX32bR4vAcqF+I2
ikgbz3C1Ax+9tL8dLSZy8Z7KXwJ2PRMIuavCJa0jOeqp1P18sFG/6yowwOZUr0w7
Ze0N32XmrieoSkczvzr0jh/rbwg2/hEQnbGqTPcO5hgwI4B8C9QBGT2PWRvx9od/
161ZeixHzPIV1xzIvndvJAKzMmZrSLEy8B+14zLtue69ItR/sPqGsXT/yGGdRTgz
kEoz1hVkG6Zlkpp8zWlz15KQXmPxutGOSU/cccpIWXHPEm1jun3xAWYSJtpx2jzi
ScAzrCrFxZQBNTJRq5RoRd5sg1Nwg3Kdfj8jNnDwhdf3stEQXaR7hpGMsqsCKhMT
XhpuciMuXi4DyXBuIckMl8eMlEKXwrb9jSISQt4TCNODxH9aK4+YctUHqBttIVIW
X0GURk7IFYnaR8ds0EKLtq2GH22Bue1E9GFTRhSP2xMzf4esPNloAKN/Joih7+N2
WHoAV+QLNSELyKQ2zoutXWuTcKscECAbefNMs79kxIS3gQioorTgi5bjOfoGAtV+
hAkw5Rwpswv2wR/4g54AsFfZqSZKo4HqL2NMD+0hi0E1RhH9KPeesRb2ljsxjuRE
Zwd/+fwFh4EWqt8f7clQ5y9DQprZXSiALivCafQHW2Dk0awuBFBE7i9drZdA/Vq/
zVklUdsQ7/hm51VaowR9WMlZHZh+E38hMYnJjD/dNFfmm1G282oTpA9SaMiw+tUV
dWyokNCT6iujsCworsMgJKIewKpJbsTY1UL3caObjPrDoEj5JohFaJoqFyEt0swm
NgJajdFzYW6qkeAlVlbpl3la0A9QncFojRhmlLoWVSXu6Gh/nROkPYstSH3gdiSZ
p6MP/0nmsOT+YKGqaKetRZ7bdvGVUvhnK5jj8e8RBuY3EDsqtwmEymu1Zq3kOobc
kFeJtkGb/JWKHKouScdwRJnxLOOjiLn5iVQ2Ufzqr+QnKRVmdu3qb3moSIgxJwqU
KV+C599+no7lXzbpeGLyRmPjGviHj7rhLez2IHm2ijI4mfgjNybYL+r9Tu4yuQ1V
INZHB/Vk0H6/NaAidvfk6qmD8Gk+pZudqmK9R4uCjaOF1Xqp25Qo7XvKqdYkL8s8
63asQ5Jbgqac+zaWu64bhwjIn98SgvzXh1aJYtFTzT7oYu4fq0Fs7fgzVt65fmtL
FfgMUKbljY/tG8MGsKkENuyIRSP8BU9Im3k8q3UdfHpYdtlwm831sf6rOncCPpij
7LuIu/WaRPXRPy5vS9yFK2xB9Ue/4Y+SiDfW6METdeudMtQcF7NZBLUPoKeUAmoj
Ha7+ADNOj0bovhJ/Ue89q58pPECgzK6ax8Lt6rB20w7MlRxhlSwj3QT9a9VFxVzP
DSPl+31hX1tBmUnCpOqeEyMU/ALNf88noLQ3tHOm4whYk4Hsxy1ehsl/poMPng7r
OrwRl9q4QoBaeh5i9vV8O5FQ3ejCFKkNzA9wjmsMtqVrr3fbuamakEen8YY7+ATk
XBFWJwyIkMl06Ja+WiN2DgPxel76x5oyS4kFoEyBD6aluMDDYMb+fZ5R+uKf41Om
Zf6stwy+Rn0r2ZwsKhfJMOWUphjIzQJ4SauDPDXbTLpOHw+O7NEPr6x/O7LTcws4
Ze5UTOv98NPaiOVUDH+ZpgPW3sSXQBYVanlooIfjNFjvnNI6z0kPPcxrBFWfRphL
mB17Sjp8JhUBz4ZCw39reWh36/sHDHKtRJmtrdJsR47DAuouggwB9sdAKVrA804I
MaCn5gsTOVBcZR3m32m46g8DSNlWJg5qdgjWktiXbUqT8Ov+hn1LQNASi+mk380R
zy+RrMqODp1UpozC31pNhBP1gZ6PVS1QHl6oyO4aFPGJB4t5OVsGElUq/3nV3iRW
MxpavjjUShzB01t0HQWfFjt9glIgzJ5bAmQewlzXtVTdcGswULlK/zoROUpkJySJ
GLRzVIqxkQ7bpUZstS+Z3NYPZydNixQvJKCxMcWfGXbUaz86xb2af86BPw2rllbh
yW1OvCVqYQGqZcWa5P11+FAFyXqTijHwhipRyMFIevlqD3eM5xBiIGhYYot73d4W
5beVCuqFN+HRDhLe5m/FWcKjbztLd3eYVDf4t2QyhYE8R2kcnto8tChTba91dY5a
PjcveycbhJZ1thc+6h8+LBTdtS9iKZZucd13AJp0MJP7r54G3eggoj60QWHkLbTn
a5Hl/KiUgJ1o0xnlfd/baKi3FEsuDCYYVPYlfBtdaYHcWizc95SFq2ifVPgr1h2V
Os2sS+qmVcx6kt977gZQ1Hp8B3lMUIutaISX5S/lYAiypyNtgBtOLtIO/xDSGVBf
YIQlJFa2SeGlG8SFhVNtDED8YpLQLPQqkhC2W15z3fppr00R30cvultjI0Kl56hI
3eSZvByjwh7t3CkPAsvtCdNW7jiv/m2x9YTKio1unIMUJLUJMvaYSWghcZPH7veu
R9F3Fhqjo0gAJBEa3DjCpwrExbTQvwl+3pe3E9fE5HOm0umLZ9M/DLH++1yS+G/X
8zxXmDnAMweWrx/L+QT+QIA5EhW/4XGFt7Bu5+8HjTtjhlwW/Kpng8pbo9AlgG2g
WYFLlk7EtP25UeoGFv4cJeS1PesdsMtYqQ8RbloI8pCS6zBXjRURqS43Shu8aOEy
DPGUK/fWsGTwm+0unZPPOHj+uAkX68DBGBudytuA5pg/rI3g9c9uDZ8XQTuNBMAz
UKNjcH+A6c5FE76k29nJV21fifd1+ctMDEI8QiA+sIUNiJSwZY1oHmakDHdMsOoK
5VJFtPen8jzAvsg/KAOa6M+XJwIKROCVgXOXRajYRQX7z/x8jgJ7Nbc2wep8LmPz
oXEHUB4y/6BZDpokUoGnnlq1jr3qdut+pLsUTPsSBpMgMVNPCo/4aaxtDNm6gcIo
FRG/c6Dkr0jYZLCTT6Y0ozB9Ma6JquQXHTs105al65G6jNE1ECz7/uxxUgjZ5115
lFeWNggQ8FitziAri4sfh62JEZ2hjtdIQG2+bm6LFqbhP0Q7HTdGBdnjb6jnVp94
vEEsDJCJc8rTHre1WUNqajVY2IM6Ulh81P/hVpu4oBjl9D0NKxkSRlHxoxgEWKKi
b5i0nWoT5u1GSj4vwFwUaue0QtePAEX0KJP85VqkWNJ0JcU332aEnX27vCUFrL5v
Q/7pnT6iKAWPkhyjF4PS/vJ2sDh/z/ZJ3OIDDFaknlDfO7nZwt0BD44iBbuyCCtY
LYrPvG0Dt5N6frUwUgPpxM/ILTNWlMhQ7cltU9CsXQrCunE8SKaw4AMzvqCYfDwe
BU9fjOSiCSax6hQ6VmKBmypWSXthmy8yTnycrfTtSCLkV0F5zJL2Dc7xCsPwcMGC
ISmZkkr6cKaFHMHHvgwo+LtDvJ/+53F/MCk5tq5UMwG76/od2jGJZTI5RyrmIpbL
9WLI0fKKTVb3rBD5A16BljV+Nydqbs6I69ANd9kfQYVFPw/YSW8NToGhHM+wxZlE
VurVCao9GbquVLFzl1v9YShvHhNRQHE1LSwo6mSBmjlsy90Ci1mBa3K6xDxG2a/x
KDurP1Djm0OcjkZxGm6IN3Y+2q3L7yE9JBiRzmBESPxf5cLUaa8x9hqhnmEKCYg2
ssCbJ3Epa8uKoZSnGrpbcxW/bqBzORJop7szPKlD0bb34/hcnq1V62PJLWKEFC9z
09YDbQ98rgUkotLQKiIKVtyaRVnTvUTkjj0xohnjkHFFt4rvXbMSpAFreUSx6s4T
xBgqtr6onXX4u+q222dSfVlrwvvPY2tzJ2k8Wj2Kjku6wkGywuIcNUV7WXWGllN9
kph1O5hLuIh2fXmlw94lEvvly8a+uwY+DB2pARZvr/T+Z6i5tC6g8364u3nlLbJg
5wwGTG4d2NYEIl3y/LyqwcXcUWA3xbzw8ow4fXW1mGrCpo5fj1MR1f1IQk3CFkAI
lWuEau7mlQPoZGCtaxrJta8frpNkxyVwKSBmsXM6UKssx2GMuIRceNuyP+XavnTi
6Scpc+rPprBVPBFJL+H7d6EaYH7mt4cRWJsB1BJDz5TReA2lN4LuIHbyHM2adjn0
xNSRTEkkrwpgIcI54tEYeSkMB8VOYZZ8Wjpm1YXJcCn53jDBtak7x09c1JBrbHyh
qMY6AQuQgXujZ43RQKJXTr25HHdfsDiCjkY0gt7dkWZN54Bxmq0Tr1ztd7J6JjLS
py6gkR3SNDKMTFut4lXiyvSFcQZGjkdtHXRlo8CoZq+GrolEklinhvw3ZbDted5L
Hrq0JV4iaMZU1LWB82GbgMI4on2PTou4inN+e4GnwYbhBEGCDCqRsYnYES/ArCIj
+VB/0mldxWlwbsxwZdI+835+/8ipbHXXJa7+4U8HkY4PmmC1P57AMOajUUULs1f2
wBaCDnFnb8O5xoqdWJ5E3B7OxVFCbm8+JPmIdqT4iV0PWFaWGTt/MCdgqOJ490jd
kcrhdFeWSfzlfNPWdqVxo7pRiZN9KdwXIi0WUcWHMD09xgQBf6rHh7HJnh2usj14
Zt2/KcunAty/gVJ86MhhrMEgn5kwBBiDIeQZFKbDYnwAU9faaia9aAend0Ngtozm
oRq/wyoqazaKKcs+2rkpWbuXUIn6dq2SpFC+sXCBZ7KuV9Su/pDU0VSM5bvQ6qvT
9SqM90bUIBzu9gj7NURilp5IZ83OpvJ5MnvllOjIQQV+XG20dhzW24w5b6Mb7btd
1hVzFWumF3ri4KuZYh9OGq00GZaumZg2LK4Onz9ucdk+JIN84C3kUaU2YMKwa8Mu
Ns2sbGYqm+uiSpLnsTw/jugLtGz6MLzs25hKKq7FERD9/75NFuNYUWCmVtrVB/0p
AhpX4s+TOhAwsKDM8ZwMnoHAxwmzW5ak7asaKx4nXKwE/ocAyTWrOaTngPQTvOm3
g378Nu4XgXIUfnWwxk9RUlnYHy2tMvcA+n8eymQI+oHAf7TDzOpQQjvD8IAUm9Ia
30DGYtAoyUiZqdcg583wQ5xRBZ6t4538ynFFmmr4kkzHUCwt2+nIemDkB0/XqUzB
X/jsB8CrWGg9Q65i+NrqKqK3UW/R4dX67podhrOe3iUaWwWXhBmt87tbU2MHYk5B
oZW9IIBWFyWgZjcT6SWmiUtY94GrMD9mq4uP4E4K52fFVg3BSRwSIe/2AKFPpizt
Noa64HongHTWlXl6L71bP1vr3BMMvuOjFct1M6uS823enJGVvpNziRaxzFth4YG+
W+bHed7em9L5l3iYxVOjndDwbGE3GIFPTGlvgSbSzS5yysyQWFhZnUv3FUs2ADkz
qaUIwNaq7p/FZ60uX6y17ALcbH/hA4w2ugEeEeDQNMyhTIEYTDcqq5JZYnzsS5Ki
1oaIYuLUR//1ylG8N9jEu4zLizfrB0KsVHzPRA+A+ebED6FuYo/FvGTQ3ENecnKk
MEt92RwnMenvN3q0Zn2HESsUHGB/CsXlFKSTJlYE6guF/5QCH9CvekZGIdh9np8l
Idzh8PBCiJagPg4uCbQ9YICwzpNlXRQ4IIEXKUjt2gt20Vh6co1iREv0LlSrMYOW
4zS5FMjLhgvouZVmqfwTbVpTtZ5YKh95mEnXSNWT7RJwvH3H260x6YAjZwy9UweG
vMlZuZgaTh658Q3oSX0obYS82wEKwIKRbrlt/C6hfwlXoREao1EZUiDFtV9+V6N1
ghEfDUBgS5Ncm0eqdvaqsx0ICPbXMqSrwDA6jTx4Q7utpgw/5HgzpCOnQBM+Afid
fts23/S+V47IL8y9THMdAy+D6GccAeAHE3tmF49WKlqewGsbANFfFnB7eitT4Uf0
CRVQDZix/Hzs7QlOPnVdkxDqs7Qe8/NLd0UcekQM4DngWse447gk4gszZGJ3N6zS
dk/A1IVJWDzmU80IPQL313Zewt1oNSbmOa7oyJx2Yjp0jy8Tr+b+cE0mBPUSwzdS
LM9m0Tv8g43zDJ/dQuxP3K/7R0Dlq9KyYP2WYwJ0ZDjBZJpwJMxRy+qV9ty6wPEA
aG8sS5vBmM9J+z6RtnP89d3Ei56ansnHRJNmxwuPZNOgKBNQDAM+VW68xsMzTgva
N1rt/ALhSsabCpz9X8UcAlBvsikdQigvdieT2JNhY72s1KWzzcqGUexSaBAs2srV
ndcYl+XXtXqn97X2QXQ9D/xiGOJQ4KjY/39lgeHRYEvbcFeikTxYEK8Pa0oJtFBt
ZKuWGFfHo8wFM3pG9R049VKYIvZ5wTnuUeUZlWPjF2M9lFVCWI/g71pHHWAcYnv4
cqy2zck7FiuAscfKaeVn1V0JL6g4lgBsfcW0e5+dSWIcs5iHxmy1YLoiHU3u326f
IjmAvDzt2DCuR7D/737aPP252jZrI8R2VYQnDZPSQH1Y9fmi40obe6MfSbhrgjdI
MxqEou/tj2PB+Mp+VXbifJQLn1lB1QQ32ehjhSB9Fa4uLGv0fOF9k4UGKirkWdfX
iYR2LNTiCEFJtBpsP2xdFbmvCsOmUkWD79idKX2tYNgsfBNlsyLb1FCUo2mx496I
fyNH+lHyi1e5FBBUkKpnm75UXSsPsubK9R41qOTCFne0OkqfxWhGKj3Toy/YkRor
JgYnH293DXpSvO4dwiWp+eh4lkWizluwVApSlWwRY1tx46R9mMrdrMhuFYsgNtLa
IoCY6uxeLW1hi9/uRWb8zgaRUpwRnVzDCC0veKUUe2wU6Voy3NImMJou96tD5lbL
1pmKtlWHcmZtyKvJVTF/iQ3J/DGTCG6ee5mZ/i3eUUkP4K2ln85X73zrLZjtLsuI
Qo4vWtD2ccZmjdQI75IrKudPQxCXDwn4hBIBlPQLMYuZoDMvYNO+S1MAm1iSQotp
Ju4AEb9hgQ84yFKoV1fbdLoyZFt9JtRpHJIa61/NbfdUx7S58q6GSiZJGyWyRhSw
IbJ8Jp9S9FBlUrp5XlX0oPDMJpdS9vPGMy2LU0oljd0l/wDog0brEmQG8+5GU5QA
jiv6qacEK3Jj5n7MyxvdbGel4HodyoIL9Ymafn5SndGAg189kG8sNov9A1Qq/sYY
Gw2TDeB4Ayrh/fU8abvRX3PQnE0bIIbZkVcqMtevFDQAbl4zervbm49e0lCfxF4K
xsOHfcWp6Bm39713k7K12rCJXiS1AuOZPi8YvyysQSJ5NWMYTiE3YlYJ+x0DNgMt
JPWlgv9tvvKxrftX2tpaI7DRiJ0EIyiAFhwZ/xF1ykQelhSE+xtfW5F/kn20mYmw
4RM342+eoihpG035aMzRhr0tuQWoA61ZJo7axnfABRT0IYJV0Fdfd7rwkVGCunhh
2Wvht1YsvcHRg4ABDfD1reJ6gcXiLIJmn+kUN/2d86NNP2YTb15zGE0kfbaYfYVG
1zEBNcJpPi56RTObjamMKYEclcfuc3z1bKnIeeGUoovybWcRrVWC2fjGgC1UiK1R
tOBAT74lsfhYlTAjU2V3b7VPGCUjuJoBlrWL597pNNJsj5gUiorBMIYVeRrYYwk+
ygWvenGgWKofpoxYt9mlBeYyTjgrq3KD+gDkDUlZ13aQPx9ePw57DXs5NkDizkXr
vUR6QlYituXWCwxDV1hPKSiePjgWUw68M/wd0hRzr19X5q7nshzeHYb98Afp7i+z
x4ta4BzrOCEvaSe8bVcqfo6T7hvR5rcq560tGT/sN4GTS6W3KA4XusVWhrkyjfPR
hmVtwL4StBI/+b6niTZsBsT13lO4wU2eoZrlOkt+vnExKMQyASecIYKbd8Pb4oqH
0S2mvrM019joYRs5k9BJ32GuwA+YISr6jW5e3EGT5Nr+NAkMrM3XF6/q6kdDbmCf
B5EGfduQZIctJ1Tz1H3KqNxxLhxMmbD+Q6WNrmFtTPlZLuR0EOGAHjZeoH8DRnuK
uYBrAjNXm23jT2OhR7q7EPyZlLPd21KfM3Mz5n3aCZng5NvrWRpZUKCIu2JG0fF5
oFJHmq57nY8w5W6wWMPTDVoCaQimc7ATasqbjQoc2uDaMJ2xugZQt6UChhTI0IiL
ixiLkdsstm/Zcjo36fvahg94JQWfAGWuVTUw33MPhFRGkyt1SmLUA2UIZbV+X5gI
dlxb3p1vd1Gjp8C5wsH+5uaR2Y958YgyHwQNljCTYKNWlm24SFCLmdPCEBsq4FRA
yNv+nZ+g6yicmcDqGz8jO97QS0GkZI9tnVklyDuqfUKF7httXeGJ6EIqmzDa9qYw
fLLcWY7W+yDf3uMFwchhwwqVU0R769YWjPNAn+5hXieJkU0bBFl5D4FXm6KU0T12
l/cnBA5KUSUaP1n8O3l3Nrt4SvvNolBNt3qF7tSd+7Pk3fby9ADu1apv4dymfERc
TN/+C7+3atb4xnLn+ismbSGMSHbcSr8LIHPvlc7akgS90HvmgNtJipXbGS+UmSO5
ioIhBijfOoD3PyYnp3b/Y15UUVIVdqAwTN63BVrbQ6gjXmmB1Bkf48ROA7t0kq1J
cuxgl/fyiZweZ6T6FZvEW7Vf3zFKBgEsXEvOpQjqk3rnzinnYDPlwJ1Ozh9pAQJL
dKKDBl58QLI3BkJt/qbrGbzohrTD0RsCwCW0bHybgsrZWFJuhx8bCBeJ1MXhuk1n
/147gQERHkVVPrCgIWhIapNts4ALHGToZ6jtRf0hEZKoO6n/mmEBOlnlhf1ieGPP
AWog6yCYTMYA68neuRz1t3B3KWZsJjxqhEO6NqoboWiDes0aubPYAPiWg/uquM0C
aimRexTs6dnS/JL7hnn8vsg7dpfJ8w84lpOpb31lOX3Pb3F7D7IapYpvpCXVv23h
LDFEIWg8UhP17gyAzIFADJIAQjodj5skree2vMjD5G+uKFAs7YLvp8tMz8PXIHkx
ORUOmp8CZAl9TCmli8ZfxrlbW5+Fi5St/cj4ZZI/V4LQqDS3l/Z6DvV2x6xssDwr
cxESVpYvAmCVWlLiwIUpz6/tygoneN+fA4LVaCfXB3fUtPlSdBgqIxEmhooFCkMx
8MYrgA/MIeqnWbQcYc+iDna0R1/Qhc4LMYNVPRQhCKbyl4UvIOC4nzIWBd2hxk9B
hMUaUq9figTjRR9B0JJEf3rXancZVyxBhNLUKBxozmYrOU8LTfLChb2yUJx3BpZB
DQg85lnOH4uXhJnFHaRYEvtm6m3DQ7w7h+UynbGSLy3/dPP4u7+lVlf9vyu0o2YC
Anfh+g3boft+tc7hUiVBS/KQE4bNnqyMDXKrTjbRU/CjZ0NkCZrBwN3kdVoc4zL/
RzqqTBVVpz/r58QP8QEF9CL79QIwFkUuDw6L30ggR5Wxr5NGoIX8P76wDnEjBK8n
R8btx5A3VhsbgH+KD5V+5KodO8+Tj2ZQbTyCPI7weNInUN1Qo7o+239HNuJaP4T1
KwAIvlb5JdafvM3lqZH8PrmhmJBOkXaMJr5uzd5Tt78T/SGpXhxm/P9PEhgcHxca
i22zycxH8mcbHq4xlmlzFEXDFA1ICfglvETbtOiNoenC3/632tiVDaiH2pNK0DAI
Kc/p/U0eYcQOZtOuXCLxP42/d3BhVCKaAAqTSsL8nZ5o7ZmcBd+G3uoEnr5rcCi6
7+oV7fJkXG4nDlSzcOTf9huEmOSQHHiSQBSFXTnGdGvdxF+Ka3AqVUIOn9p1kFQ6
/49uHRyYQUhjxQkgNUwkoUClRkqvCR2VVzKGLrlPzUDiCLnNcfUBE5eS0TQ6wY9x
JCnXrbjifcQeJWVt32sRAFkcjMVNbwr4Co5rFjSoGVozTwDj9NBe8HL82S6ZWfQ1
vpLabW+5leZIVizUmrPglSGjXLB+JONCI0mMQLbFrG1VmBvEbHdrrzWj9GTNLJfw
bubB/YYcS3KIZQKfM7fB0gBC9tSnoy9iR21P9OyLtMaXqQveVvswaMj0JBW2jy+Q
JCT9gSO6uTbZTxah/yseHbWgkKrCcC1H5VU06wcM8e7zqzQHVYU+kwKhj4RD8xNh
bXtUrSuQye2ElkyNuE4xOmC7mo0xkNEkS+x+GljheiM1BY1q3xjnpVMq4riuCfW3
c0kFCogype26/Kw3txm7jz31bclhL6QoFNWAkOvdyg6AJudNudCWl6kdocv6bVic
YhpOFxY/i6QB5U49LpHxDYCMytrcmvQKTuawP4qhC26jVp0GmpVmKuJzFd4DZ0KG
P94lLcDEDDpyx+1lIhC4ZVbS19gevOu7D9PnJXa8UyMXjFvFMbSKVidswCD4i0r+
tPM2g0PdWGmnTEE+atp4+/fPursqO6V7+I8excL05zmg+rGdk/WagL34gulyQCkX
Z8gIq6vJf0jRNJT+yHav131dzzVf0OIlSTETVkOAowo9w+urKyDeSkMEyNnRXI3S
mIwYDfDBgnADWp3fZ4CkebzeE2jxdi/zETtxTNkgQ9XSoLMZtig3EpZ6/b09H1tt
b/czZR+0BptYntGOGVu00P9sS0WdEehx3U+ofuNr0o8eHU6lJedv1KmIFYWTc8Ym
8vbMWg15VNxV8zwS1igjkNm4SI5XczrhaMXwZ+i2d+n3z1dB/FW9uNbfkUv3iSoL
lCSc4k9FooX3ICrD0CxaHdKVNakeOJnwHKiJJPJRLhHdxJvNUTAwmdo6sV8akdMo
giS1QZLuo3ljO9wqR/XaGQBPvlF9FLHLwBHSbmMTilWfJd0Q0+KocXDu9PoWr7zT
QADNeUuZ/WpDBGQRQ8lSI67a26sl04YsT9uaMcbz8FPy3dLCZZv6iCNoRqEoym6s
T4yseXrMq6P6/uUmvGm5WvzR+5H5dD2pkKS6P7D3MpquNXryozIQomeGki1Y/4+4
Lv/WH7lK4HsN3Kpxh67eydGbVdGOlCOljbeXXzU7lddDB38jiCACQp3rPEjHKJHz
2KYOhNXeH5L3qaF4aIEir/oYnuw0dLVVhn35bfFyWGRxxwN1c0GQfwy/kb6//hb0
zQOzSRPbIM8pQE5tGmo3Gp/A1zhWkyuMPXuH42XGG1j//B3rPr7S07HARHEuP9bJ
DN9at68ZqanIs/1zWhCwpPd/zXg2hUrlXyOheZ5YbMdS5ooXuUZFWRIcJRTO6W+G
9FgruOuwoj4z9fBpYKPYPn64Pl/v72CuIBNVp2N0DyMeizURbBt+zycmym8UcS9O
bhYK+XfHVk3a8wpiwAyy+OnrX3BVdGRa2WiMHwnxROF4t/EYiYUmsPNnlCW0+3IR
6VkL4r1653wl0QFHB9pOB8OX6TvOO9lyFm5H6qcBGlS4w7sSLCe41NTSF9tfVyoC
qc7L5U2JUlp987/01cf9S7LCJixbCRBDE7waFjA46icwjQ5tnM/y9R1sFEpDfG14
MBEzBj2/LY8XiHPpNtF2MM3FJD4e0U6HK1QQnSfD8JZ30qyHOvnC77dwuGgeTEYz
0Lxb1O2MFumBsE7ie1Ozcp9AmNa8VJf2moiZUmCFNzG5k4opqWF/ziG0SbNGrdSH
CbSJ579e3loiiVeGMTHbQoHgECcG1Q97m7u97PhfKsGxpNO47+pdmHeSnk9bGAsR
tw2iMkRS4a0Q5cWRUAUDPCTF/Lhym75jKOAgWLcjsMzaVk1rgQYrO7JLsCf3eFEA
H5kaKPA7jKvswQAqbqygMvvVRx26K6MUggklw/sm8w5+8PHzrdaLM46OdeZJqSZ1
TJlr+uFiXw405RsrLJK9+AA/xukifXhYIhEFp+6dS4vifaQu1jIsqgjnly91jBWL
jLoQz3W/Cf0uQor9FAEXEXvi4OK9ubZjNWMU0zHyjfU4qTNFtdtRdLvs7v4H6diS
8YwBdDXpf3iyWJfUtnqsyk/C9ElMpMnCGbdw/apJ0waKaVwF+jKTPN3kDsitIAuj
62Y7+qx63WS5HTVuaBBwyInxcu2BPKGonMTgp/Et8joZ3I7C3hm8uNoQIY1bdipt
gyWMKL2QcLDa5M3KtTF//AkbRnj1Z8NfNUMH/FVTqU7nKfHZFYSc2ao/PDYOwyvP
Agg9EEYdPMNZErF0b2j3vVtW0WNIqOfsxslm9cICwDf2UHJB2wCxwPhVE665i21A
oJEifyaASEqVIEQ4YVzmStScaX5KdSBz/v0GKOWKjtxtJhQIJPisd/2AHwGAS/XI
FWOZvPlXx1NM4zoqMUIsRFn9/S21xOIO8DQfGs5htf0RVs3d7EtDnzbEr7ktAqai
ZyfouginPs6DYWgmIHt0U/+2mcsRxCrq1EiLl7TAM50BdfXRHkFlvkeKSFeKykfC
7BaQVSmMoZnChJouMX9v12nXRSwhLX3a47Wk7DuywqNZFEymdQjYEWeTOQLpb9Z+
FOE/k6CPBxrgYly6kmY8xqV3wZ0KdN7HfWVsIorW/tecRqQdhmhncHQomqvjgyqx
HUSnu8549ls/rM3PFl1qHVfdA6Zl0aeGvTJ5ei6CUMCdqm3pQN5y0zhCzeB90qiY
TNQJfHmub/2CYmTB5Ebb/oqriybTXUMYO+bFcFpUg6zeVyTbVcQOC8on0g5kIVdI
urgIMcQcN4QnFDsMpacUzThB2slEEFLvlYQRpFcjfj2niwpz6YoqlEsyRpJHBgCF
UXM6L2t15fTPhbuL+ZjkhDYlljTn3XQcSwvWwrWS4cZ5XsTRelNGcqUt31u5Wncl
n/T4edRB0J/yOQN3tHQJVum+/2F4uwKPIBeJPAFsbdU3NrU2/jECXBIkiyWihRV2
gQ8l78AnBUuSE+/eWPE2H5oVWgM54+K67afJWLeSLFG28hcCpvoGORw/DTpiwAgc
bxRVJitA36dgqN5yO0YHL2Pn1h8UE6tifqLjHTAkRBzItv3rzpMGCKu7NjAFx4kT
PQ/fhehOoEjAalOx7964LjQG2Mqy/k5NMhh1O0zUKJvt1YSEBmaCMZG5MujKVZZw
+U6W0A/a+hZhwPMiZ2mp8hv+yGpnHwwUE0+Knz/koVrxEi3Dmv5qiGo6QVDRKUQ+
bTNR47e0aCIBeAIyssrDcRyGBi/wif2/4KyOyBYcIANjzPFBQpMa445djZvNNQVd
MjjCT+aSY2qMaZrl0XsbMIKv56j9nIy1MMtXIe+uxWtBTWl41r9jVJG/vrsD7EKc
cuoW/kUV94PCKvgCNpDuOaHzzQcQM7/svwagt5svrhc8XRMVC1ENbsqnznrOlBV7
OajR+Ro++DQP7NqAeOzcPsd3jUQMS4I7AzFfVgTdGla+8E4cXcb9uQE8/bHEasbf
m6KpNzJicVK632d0+Yt9S9tALoMkpzlbkLPyn17OAtoCFp06uSEVMQkl1q1eoBaO
DAsQJhpJnAAxT/lmTyvMo4OwKzrnUb3k+9aG+kIuPLFk3tp1xhuJbt1jpT4nOtQT
pFSG82z3QDC3ZNOrsy40HmHMOHSDZgx/7aYDDm54vLwYIDw3w35f7paJIU7s69t9
a4+1LQkDWcq1RnWJodLQwtIK0waPjSywPh14pzdqu4xUPV7sxTONGfe9ElfY/OX2
68q4sGz9ymJHTygt7D3ooTrJBorf8Ob2ddMJqW2ZaGtSaU+JiUJCwbNOJ7LhcY7e
vWFznuYmrwzHfSNT8a+G3tGlBmpwtFD/MbE5a4He2ep+ubByx144izmD2xnIXkb0
9I7g7FL5Krp9AjD/wCmEeav4m/TyisD5X6jvePtk2hHx6fDR5r3t9Bc8SwI1hP32
kIUVRs+esBcs/8xQVWk6h9p20jK+9h/3TIwneSEBnLb/+ungVYPllttjjMTET1Sy
jWR+EJ4hEo9LEA/cfScLVN50zg65BHg24XKbk3dH3caVYNnX5CIigUNyTUlRzyCM
W2Ybd6boszZwBNqhvnYXrBvgd+9g46m719uVoaom/HI3v9r+3aT/muiFrPaRSDRT
1Jzpz3vT2LeRbgGR2MPBbXkh86IcC/TBijoWuByXS+QQQ8M3Vb1X1v35cXTe3+Yd
cWXEM6ad/sL0DQqjDWt6kyz/hhAKWj39KYSMFJYd79zyDA9F3rBFx3NmxY+XROWk
Nm84jAbUTujZt7iE56VJSXsPJEFX8N5oRPmx/TO28JhyBIy4IaHXqW3txPihBLfz
p/DLaW0OC/Lo7m5JnRCTR/9f2xBuKlWHPbSjddrlvfl3rKbtqMEwRcmQkyHcdrQn
0Y8JtXeamCBlC44GOoTNfz2RcS56iofS2giuVQuKYTZVvf1vSsInPH+EyLgj71ua
+cqMqbKhFDcPYRlOLpLHZUw/lOeAuut0zNpAh3+gImY/YBBl86fmIwnekKh1M7a/
lbd5WuvpSPasPRa6EvkzNniTYW9dWZX43qwRmELQlfZhsNLjx+0Z8MAgMRSYLK+p
ZDHoasujrEckAQ7KiHKe5HqFjVvJR5POQbjSpL9ybs4IqZbPpOazfYs5Owyk8xSg
wrLHLB898bpyNkCvVz37GJcOiXR2PetPdAuxKebOOjbnKYwf8UtbnhkGyaoBsw6/
kipGnzigvI9G7ORFoPe9cPQ8u01iaKOpi8Qvhfj+3Ep2lQHfrMZWnlHjPH7PChqV
nQB7ByTQr/XSnWyKgnFKEb59SC6WRPJafNKkTAMQ5Al/PhNL6awPiS7VtP4kJTqZ
tIbv/Th/b0SnO43UPSJX+HyrZ8pH+W9jDKX0KHHIpnckEaV6fBl5IWdxuf5rr4fY
76cM4WRkKkRQU6tvdEPnz4d4SJTdgRVGlSz/HuFHJrDR8He7LSQef+CPLFiu78ih
NcLo+OdH7kOfqZG9AuijgEGwO1hLj3CiXj1AXIo3Kuc3+6fmL9WQSjzdJUusWXUq
snZC8t8hPDVQYSZAJCbSgDHhpPo+/BlhvdSMjDNxs6kaL6u0knNBGvxQKCoRZBgO
DFenHXOMW5H0UOF1htji//3/7ZQSs2rMkRn6Im0uka687A/BpSg5JzyFS/Wos2C2
Wk2c7z4I2H2Ndu+b5cGYHFwOmIoIVcjhZnroIpYHws4T4J9mMDlssT6gwMx7VUVf
6rHCMTGHLMsV2ChEKxT6WzxYbzKDjvjT9YndSO+Bfmn5tt0wg8ULrf6iFGWQ3kmd
GOKltcmo1EfIrzRnlVM8xlMUilSMfdqja/v5SK06Hhig2ZsREjI8NBiGW3knbTi6
Tod8qWu9P7TlBPrH0TrIoe3yezkxr7zKI0rBQomugtm33P7xzgt6qKe/oIEbmW1x
123KFse6mqG/wDmrdTJgpZf6x27c2bvgaG+Hjx//m2rYnyIDRn4xQmCBnKGN00/r
qjXrLSmg4/H3j6Ccn1kCvXMKwbHNDXvDwd5qC5ova+3hbXUxwsR2wkSEA06VsC16
qe0FnhaB30z9W3zRBGo7dLlilRXiX/dexYJfRRp4Udzho2aMinQsgwROmVW3Cl8N
owFASQC4/h1bC4qNxxsf3Nd68urz1KLzgwn9DjgaNxaisYEz8kl/Dh8H49zDdIQ8
bWoFxR/k/JgQy6J4xKFqEyqfYRqMLL5rXQrWdY+miHxx1lVg2VqjAyYUdRYVf3u6
4Q8eIUk/pQJIKVLp5Gx/GMw2XoJ8W64rueYZ0AaqCvNpj3/F2RgmF6E57UF3WKmF
H8iY+kg3L5wGltCYuNb3ooNWBOlQjPfQ2+YVEoGzNrmQShI+e/GKfSYcYH+9WYil
a/N0b02MzH4bxvRzNL5h6QKl5VPrEgUCI4QAMMgMlGtD5zuFVAyoI7UFAPwGjldz
Z9rFlLFUiEcuW+52B8Ix9ptWwLb2irlooRyKiWhsMVAB/hTa5orYa466+qGV+vyW
dpG5vH7p/LxyEz0NrcI5ub9/QJO/MyX5p+jSq/EiQvI+XoBXvLWJwHJ7HmO3FBol
VwulJhwaWtKh8Zt5ErI/M5CXmkoKR6gu4nfmA+AqPidPeldgf0syrQkXRagwndYA
FF7qSDFcFvY6WUzPuZln959mYeWPp+nkSd9RmQh/XFj+rRKcq5aqxlpMODg8G2jS
6O7Z9usubeynobwG3g/bIkQsFmHGv4Qbo6Zp5VseYZa/qDlaT46CZEaC/G6AKt/I
JSBiu2ipImgARIuRVm/KbmsD6bYl7aVnGMDmxgVZf99gX3kusv0orlSiXh6tgNWF
OGEhxMeH8/cABd15cs7zU6s/XuePHaTVDAojNKZUjec39/QsYnOeLWMwf0iLUSc6
qHRxLdffU8FT744AXD3oOfhfeEFZOtHlDOD3+wZORgrUHviYmcxRYUXi5iegTdDS
JpNVP7tfYuzaf6gzYWM1z0v20PHhaS1j1PL/k4i0o4uErstrR0AKel014KvWJ7oa
wecv955RACq5KIKxQalqpqG1cARvvhxDmfGKVQbIboP6rLSCEjdyKQpj1tE9M/SA
ZVTgZyfNr1tDS8W7juICHAc92095hmLIOkDfrdJNhjFJDf8P3t7GZOYQYQLHcs4d
xF608a1Mv8Wc/YFXUCkeoXr4KQGHnJACPVxQbtorCCyL/MNwVd3S05vbBBmVI8hY
Jxjhxpyjb6ICP1YkFtxEos5boz7Ax0e5tVqxAzrDN9EGewZWjMinxDHFioyImDCZ
4PboMXABuAJ0/yB+dEuZKrHcYMv0ZVJj9gnKqH+Hk19/60CZZScCqYxy0oPgrtZR
hOfRRxRmWaeAT7KoU92g5ljFntr5jrrb8ktBiQrZV3CXpniXaMdUSZZzDOUQGx/N
liTiRzYm6e0WCE7a5gvzkV8sMekS6zuT+ru0uR+JA5Rno8MFwwDIfO1cbM6vrPJu
9tofDUKhzdumOticjJmQsloH7U1br1qpV8vPx3AdIa6RivNzH2sio8nCRWhvVtCc
1BruRMVRP2kDFVi95ZARBv7Qjyi/D3UxvFtRcEFjrk7kNyprqSrUc+GcHap+3l5P
gpq/ycCxvZK3BxcoHH3j7VLkaH62Z3ODqcJB3xai56OWgX0AIiYpCvaK7fwqycX6
rDkU3DkSuD2uzD84ynUY8h9wEY/8RU3q8k/Cai4uyrwiLdHYWLhzObB1bryVbgMX
dAJzszOmfecaeB+n4GRCV+5u3zvpmT8rv4wXzGATAsKAGXDkNvtkN1wEq0SleBng
hcxjucN+Ke2I3t0smqxKBxH0v/x+zTcb3V19JnRIYokXGRUse0GkXfDniCe17q3z
ok1L8dU5u6PUlihTfbCsqe+o2DHFgthcx8LgwHNXOdjAcsVS4d7bsQQ8tFDVk7Jb
fDKokix00IoP8N89lnwYJvIEf4gnCpDaxa5dHd0/D/+RzbKPqXtLTGJEpMtb9//D
5IdHxmla26yN2U3Lt4+WZFjn9I1pp4mpbQi3C70Au+/G7tEeGdXGGyMYdfyHcgS5
MKnzH+tbZiti7mF86OEL0f4I/wmZBsY6hOjbqzvokBZ6Ok0YZD8AG1rnpxf1Bgsg
1sFHxmNJTjC8mFE7gzRP+rGgGCj2sL7qtf8qPfubM3xAbK5D5qWZy3NQsgAYudtM
4IQmfTVydQHTegnn0jB3+/5Lemk4OYUTCvbzfyqbrqAzbXNP/LcZnxYaIDpQuVh5
1pHTCxHAjOjt/NKjPk8lzBrbWulaLLtn1d1qBJV9L3JPwgkjfcU5dWY0bBAciHTd
E4P+sw79MXEXySvokThQMd2Up9Z++esALq5bLBicpVc74+03rZB075bbwEPQGv4w
AnNeZACQahmM286/KPoISAxXbKDacLUQBRxFNV3e7VFZTBysvTyCe1C8Vrg6n2a1
q0mf67KFk9Q8v7TvrLWf31d6yKxY9OyQi+5kmRBhxMi7xJGlPHWItTbWRPfV2Hwc
be98G2DEQ4GJmHbQgAw4MCDeQVdZpBYT9rdqWkML42GebIFhqxvESmj1hr1xYoU1
rstadRNfsP8woRefWWZ2jWC7j7Taevqj97R41XJXJdPH6MTU8bdmYEMdVywuMlYA
/VS+4R93wUgx1IHAQPQxBAxfvuNsqSu0fEO774TgJwSTYlGyUdM2saoaXZYPaqYb
BIfYGdd8BrWkc5+lcknQ9JGBdl05Hru5Hw3hatG1ZQ49o+8wJN9i10H+jQu5LW6W
mAKnHFILtNh4hpc6Jc0i6D6PpmG5GLc70D1NX5g2rR2ZtOrLtzmwR3R0lNGG/6nd
d9zv1aiM6X21z4kfW0Qyxy6L0ParbJAlXUQ5FQJt0l3hMaBIr4ET2VYnUAsDSx7S
5y6AWhAKzCl2SZ8R8Y18aG+CPX/n3WhyBUFbe7Sj04Ba4xh0vitjAJBDHD+yvzHY
nCa7gjmv962rFqPWHo3M76bFfFIP1CTKP+MAzv0mWvFOJFGBf2IEKMC5AdFOYZlw
6edZALNe+VXMqbuZXzcM9LguMgRfYZENdC7nmFxzvri7T4cccTL/tE5TvJzdQqK3
L36BoYyTPitnTlINnRWFWXhwRwhb+LiQ2PGM7T7Lu97ytkBnBZt7qt7sS7myGnMc
XWmWShHE02dKRNNPHUgCV2nKFEb/FtvN/XNY7/jQZDoKPm5miwGuyRkxl2bQRWmM
ikW9FsTx8E2knH+T4xOKQyvff4ZPsoa5e+Cer+F1I+6J562tF2zG4faBMXGmtF+1
Qvcrg7vSY8F2TMASoIPfO8598ZIXGs6OeAmz9p4l1IJk8v0/TzQ5s7HzSbrwee1D
I7ZUFbQNcdQUzFvi56adyCPnc5BYUAlw2CHhA2C6MmRnKoxJYx5ydufd6RIa/pxw
1uzl1LaDKJ3cpaEiE0EyYTZFzFUXQH/Hr6LGBANNEG99eek1XxrD9odpD9dAtzgu
CqjC/cPMJAoCrqHp0aim+mjEhxmQkOyH7+WpE8KrRelS0OsgSDz76pUJEVuw85WB
Wz+ZOIDWVc5j+vpAcBYXMRFJHVlNhwPRztkvBVa0j5hjUdpzMh6v7kIRQT7FKO48
h67yOUP+KXpesDLdr5a2jLe+TMPOazr1jY0Lx8EEYKNncydf0mteNlscMBT0dfpL
xyLvWTmKy6ELO8QU8SM8mP7C5KPqwm7aT9ffw+6rbHe0/L9WaC5Q1zoDpzNv5JS0
Un3AEaMRNKNuHiNIywrAQHBZjem++xgVc9xbWZWbx6End6rXGGL9PvkHY63aCNLH
NLIIETzMjXo6NJqZPEhttA/NSR+pm6zmK9nvIThkmdEzSKP2RYifG9/BH/FOpqKW
Gx7sXqB6SZR6xE8ShjNYB28uJlfgrYON1kBPaOxPu6LX3sLq30SnpxfeXgv1tuZW
vyKEcK2kIQxRrflSBNisjgM+gADl52eNIAyVkznBDzSbIn5d3Ox9XMEOT+IcUTDE
WVpivFGglFVbBHJgKXX/ur9Lk7MzyOBWtvWqNKxZAqvJ/2qZTRcT2mOwfeJ8bHL+
H1mk6xelxw/ET+LoSAL0Q1WsPDjLdnRTbCyQopZMrHUcsEQI54a7iXhP8ittCxwr
/hGV5rVQ3fWC4roOkKIprlvPKV2JxbuN9kROLiO+b9Gh0/NrVgl463wrJIfry6Lu
yYY3v/EjIjtc+SissGnYTJWoZZxFV0E20gQ+TNwtBlsFca7qPhxoWH7fBR3ybc+3
aMo2bxQ3tEdQFEQl3ryktXw0TAQp1DgSgYyDeHIClSkD5U6Fu91UtWm5Bp+XZVTT
qcZlH8br/hWjoG1klg/uPInC1BOOb5kXtI4dE/2AHV2vP42DpavkzxtvQx2P+P35
yXij8YEF8DmX432HitSKJq6EEGnT9Ns6BX8KU2/Tp0olcTlmJquJPFGjvUZ5Sal9
Kf5Zvp8w16MEy1AGfh4rxo6B3kFHsyG+gmdHnmwC35JBee3gLI1/VXEodzAF6aix
aOowoATXUAfFaRlTl4pP72UxaG2Z1QxPdkwv4ubVFRRRR9Gjm15ar2O4UZqLu1bF
QznoRya6RnWSkw1Tm9YMo0M3ZEqv/cPjLBaIdhbjrBhumlHob8gPzr4AlHt0eByK
a0hykY7KEEo5WAXD2WqHQ1Y0qxk/PU6VR8YVt4Awilk0sM44AfnAxRHTtD+mY6MH
7lRVhK6lyqo3WX3pubLvE8gHcvZC8Dmn2UTbwWV3R7xrBgDTG7Qk211MVTsPI4bn
i6tkr+fudvlU342y7YqXJt9FxbW8vUYOaYkEEcdJhztCQrFAfZ+gOPppgGXnVxhi
WllKgyP/US+80LYLD9h0PObmkPrYEXhb1lLvoZIbdFvBLZQcmh2AxU9r0M05HXV6
FML2hQN+OpTOLBBoyRKqmZrXBlKcCK9iPtUFaZnS3iPyDQAKTbEIA9f4lPnIwVJK
vgjwtJIUaZp5VgZu60AzGbYB6SYxYQFEfaY9Aok/gqbToG4T57wBJEXrSFqefRXd
SOtANRx5rfnkiBg+qQKSMqKdd2qFMcgB5tW2OunaJEQZNlZN0/uBSOLIaSUtwcGt
hwCPGMQsNqfzcQtHPKu9i0U3NR3JxMsC6JiZG5K3K3GHi6lYSjfFV2w0CuixzfGJ
4ICE0DpDwBrWIGULN+AEOHl3b0YmG1vnhwoFME2a33jLe9d14FBnUwPhLP7QggY+
EkrhmYMIBQRFW3RrEHEtmokSOCEWZYVM4NQfBQMvAqcfJNVyyo7MWkmcD7vUC+kj
qAaHQ9JzRY7jbfHWfowZhfEnWl15CQSgn8zWxNnDlOpdXK7hHJQ0sZ1Zj3hSUelB
opDh3Qc0jsh1Rv3/gUCVnWepdEBg/QYvlfWVgoswAfKQEErbKSn+AAISQopsOjjz
+H5FTeVLxB6u2wY3ORXBiHhfbTi+M54J2ksbJfchPI2sTxH8puxPOwz0c1vOKzek
YvJMtcesIQ0uCUiz01yRaYI6AoWQeUDcz78EllE8V4DzGflu19xmMXZA9mjm8a/3
9B3eAiBu/IJZiUtHhgOyGPHhVfA/vuooDcK5qvOnfAhBiHWzI7SqShinuM7wWybK
feC7FLSXJidNdQaEWY9lqzNACtCjLGilwFZkqapeuzkpv0CCJAyjYVyKYcjvohxr
HtDVCCKNbE+ez/5mODTVjubxeWaVNVgFMgDkR3HyFmhfZL9SGgk0BKcgU1dkoslX
Wlgh2D5B1do/oSHNEJEv2LDbh5l+45YyL0GBHRfpT2X41Mca3OIYP33k+fyn9bKo
8M1PMakVyra2QNvU3aF8o/LNNaJqj8fpGmePE9LyoFxlB81xHmtTeVAqPK2k/iW+
wdzIZIFVkkwhjFJYYRIhZHIE70Jje843e+qJOEOFBMnJHUg2TV1Rh/PZ8ijyRuAM
yUWt6PndNcDpPMlh8shKmtnAsQO5bh34wXkGP8Bg+L4q2ElS3tF2OeKxQveuh5WL
++sjB7qipdUOJ8h4jEfbC+6DOmrE7oskcAyV3OOl7LYz8cSOhIbsb7nryHI+1x8U
5XYTV0nm00inP5Fc0A1ObO53IdwpXX8lu8brtOrzagf4KRfQTL+7F4X7TKEEKbvS
biKZ3rtSe96dxbyUalSzqO+APk/n4bb6o2hiknpSQ7sThxl+3WyvEvndvDRSaebc
nAcZT24W8RjYwBpk9UDti08AeYPPtoYB9ZqTNyo0bxrwHtbI7nlgQxhvzPxBpWxr
I2lANbyuIve+tefhingwTG4CUZ49UVY+d8fmCfxZNln9rhGb4TRuyTPRRJ7OJaKj
+422joIQifJ7me17o0mZDZfOELx6eRImffAjwXbdQ0L6RnFHHTruHgrUw8sd/m5j
YpjwneY4LXZnwftF9s2I/WM4QWenSPybVjClDzfnWSEfeAZvWL/pb6q9KUDVSAdP
/TRGV/vFB6rqK2IJyGab4LW6vJrwNK+djJTQy0g91y8STE2vq68lbTd6nQ9w5JZy
j5+QHPMUCSaH6BlZaxNNguUBBqxl9PZQ37eUoNq1VAJnoPNAn4Y/ffYY/qtxsON7
nSAKHF4fhCc/B2EbuaiYKO5cGAx2zeXIxTX5lRNDc0/0U81A0k8G25VcHVDJcvku
1rCATGtGjhgCd0x1WaDsYOlkWHCIPYvBzdQOgx9JWp/tjscQexb7IfGQVQ/8pfHG
FsU26VhOGo8JXQxWMp81G4fTLVo8Izw1S7/4jbBhkaCdV5g8gwr5ailx27PL5rUS
4Lesod3QQP/vtPdzrjsgv6yMjreoi4HSY1Fb9183lf/qKiuOXjblLZQgNgAUaija
J83bzABS5G1snoxtKKM6Us3P9e5fHbagcC/LzpGmAbwuRDaSRsi+K5KiicIKLVL5
6JyIVpbSoSFrgLYQEQm20x47vIqeTWnTAiYkVhtW2vp9BfSy976Ko03PkpPaNteJ
GsCSfYBtKqMYd5cUBf5aduPXyl4KPr9i7vI5BDjmC1+8UFC80SmQ6SfKpQtH8KS4
4sgEuSs9XPMdVBpkuxlIiE0vdmNvQrgFu+cRz/uN93XwGgkUZk1P9fuh0k5Z2+we
lnnYrvEfjjlhNjJynqdD+ySD8myAlDktR6QB6U2BK08wMNthsRDi1RUz9VbrsZuI
voWVvfVg0inwYykK+NYAbtqHmgtN0BAAzrC6K2b2APFkd+PI8LtegmBu6PSS2tf6
CHc67Nmfh2oZHHu/OL6VbrrT7bhJYOO74wbFCi1p31BbML02VCKiYdHh05CJqeoO
uSypqtm3wR9dp3d9d29WZVBh5GFgqkY7uXYnqrevkdIs4nHCDZ+MDxwh5+cL0cXn
vZZ9HfPmsZ1zfuNISleabVMoX+/x4DoXqjvVmvnkye7epUUOG/gmasr/xR9e9Rzp
e9bL4W4fC+vnJ5SB1yeVdkakLjxxj1ooHdHvDVGYfW6Ox0M0ti28jAyxVSDG0ARD
aFQIXGLLQWVdWep0ZSCMn2AWqCnxZzyGl2dRjbUGGULZm9YXIUevquPg/+0zaaLe
XRcfCvtmdAkTd25XXhgOG8NXh0MUKYpvazlVq3KYeIWVko3L+QWAcPLthmGCrSRK
TyVAErUHNaN3/6IubRQYfybs7vnTUcSCbFIN7YrHw2AO2VqQQuNicw0BtyNf5iQD
VS+zfGmzOge/9rNv7X8KOceewuhCqcfqb4E4JffpH0wNAIY772ifHXwQoczwJFCW
ZNraXTQDEmjZiTSy/+pf7oDr/t1Ex/R5eg5um1IAQxlf12badGpvGHqI+aWWMrAv
JnKFo6p1QuDeE4mRHtigytjwDU2Ord18bvLiqiYT/QkoF6uJiKzrZkuPMEuH1Y2U
5W6mufB2IHmqLS2i5d92XtbzqUj+JtDgiTP3gQSJV66AaANTO+FBux5SnqZ8Ltyl
yONFvtObBbMq9NaD6D2JA8aTzI2qboBJ8ZkPdVOk3YZQp+R43fymU+Gv6sIK1J4h
g0iKPzAOR+lqetqmKYZVLdMiut0ujjro+eGFUz3OdJIGBsVi7LxN1RMDdo9UYeHm
lzG9lxHaQamDZcHNzSKJ2HDJllPv5Dr6FFDYmN79HykEgX9pIdEc+hskObvRSWe+
4OkOdvDvEf4uOBfX6Axfduel0a2U7IyMnegobc51XOaxiU5aIvqNvGohwZ8dN2et
PhtU8rqU0ZomxynHSNzvLh+r4FEjvX2CrpZj1rgbr1GGs/pzC8nmuZBwOp/xW1BG
mVmGuwtzh3OIPSgwn6EoVz2tflrEDLRBzwz+9H6xENMKwVMgApk0QTSawrz01yH8
MTpj8Z4Bm5Gdz6mNfNnnyRmdrWTUcX+khSuezqTycL4b8wLaYt0B/k19jh9tiHBh
nDKnaBZS4K8gOVFalKPqe99uTO/pdNGiVqLty2+2iQW460+mNd2l+bLV4h4iw+m7
o+TTKjbY/z0NF76MFa/SR0I1BAC2NOIv+tA4JOMb0HKLpzY3RES/YbDl4Tx2fbp3
qhjXCazkpSsycE0fEN7kqYNmBgMShKJMFW4ezKlHGA/PsIeUN9TabXkoDOOq5d5u
by7rfP5rKmQJlpHJNZz8ojT2a815ekt2wkPVv66WnwaM351N56EWrNM8Z2rYJ0Ge
TlCWHgvSknY6dj7Na2BvDnmtMPHcDBtZ9LCsQVJ2pRZNQWUD0IC19IuWeNx9K3cO
FQsZo6OJXNKrnFyBOMBJ0kcvLwMSlanm+l2xolt04qKOfxobVdE/IYFpXE+PZzVG
Bmoy4N3XQ5ZYWhscwhu8uaI1Ig6LD+6tqfSiakvvO8lamovCTlmvbO55qM0DwGuU
Vg7bM6X0T06oiw/lZiJfRguUH/JsGbbp/a8jIWufRNcvHvKsqjfBBqhb9awfurjP
L2zabr6dgLc+wBfUCEfy1zcgaQOBg5Hhs5eHBkQn53n/TbprFQ33ki4ZWEjmOTfW
gqTD2Fe9HJx1OgxsvWlqKoWASzh4KyNBO3F3qmZg1NVBguHL/CmynEyyzK4y+qAY
AjsaqNSSWpt+cm2V3WBLwxqz5iDKOh24PGepgInMaQaJ2lq6EiFkOlIiyAezGkPq
g92v2zj9r16XtWmutqbXN0E92/veAV6G05n4DQp4YRKEI9IbHzq81Wd8c93CtOyN
DVYsiosralyXr38yDFXu91HcSwjNWZBuxDM2L4v9p9dXYrJVOPsHfrH8c0JbeDZw
iU7K9gkqhm/CJTFWF+74JmM7oC8deMWJOsXv7Fz3ug+5oUh14liY/7yGaiLYwITm
aO/IudqYMWm1mfO0cmxYlUFGDCSGTXybyamx8HevE/S2ouIGWwWzFd5t3g/DIeFq
VNoKjMID4J65BO8BZIGNoS8NfuG/KMEEGTigrodFvog4yI0jFSP8sIi8WmYKHjZ0
TgWMd7WBSBYkd+JQPrrHLSdgdKkPAn9w/FtqRPPrBkZxDVsV91ptL/z62kprQXjL
4eNJxKTQzovNSlcmfBlIthiSPDytYVJvNi1Ox+IRqwvLHn3VT5cNcfQ9melhw5tn
PRTOyguDr15A8pC/oURiKSJqNPjH3b16ezkkigJddBpDNuFxk4BmN96ZE5yUx5pr
9MOYg7v+l7w/IxRQPQiplgAZxk+gFmDBElrroRtrBxjwFeASOCBUoPT2J2N/cgPw
RMiRIy9qEMhHeAg+ZMgYkqFudbY+minZ5OOZ//88i3buL5eYR+2bA4hsSPfDSF1u
x+t+pLvK5GOpKIzNUNwCJM6nME9XKDCiPNwPl8tKL58RsgnODjkb12Ue24emlEX0
uEYGkktjImY06qy2oMzbK+T4zVLY0teggtBzdbIZKZQhGJ9B967PYL3T6VvXWlfT
oBtnmJ+UP1qHxU2a/KFIJgQWkEdTfzMW0inClBiVDnoS9WIgN4LizGuS6/67NAqZ
L24/ANsjKpPI2pf7+SWmbema2yY+40CBTgrfAn9WUY1zsHmOn6YW8+L02I4vieN8
leelEaL+vw7T/T8Ys47/BseEawM+bICOTmPdnzEbyfHAxsbvWmNusSuDv8WzDOa1
W89dAC8VJ2v7uw1HxZPngnfW1O3s8+GUZwzw9Nb1VsgCKknDWlPMewmoJ58hTnwF
UvBu3V3R1UVm1ALGHgjOqMGCOr1W+RciixlbA/W+9gKLkurxkumAKZEfLDw7etHm
hsrPHoWfKTo/Bkl4tsAkB6JlVYkCB8KQIz4hoQu8Tlm6BUrfLfFxTfn8sW9eQaXD
tj4AuwVQGYG2fG1IKrx3XbjKn7dIeepAKJPk3dEwAJWT2doXbhqpEzbV4yTT70mW
lhrWFjju0LEYVeg3QwC/H+hYmq8dzC7BpuAnY3PShvH1CanPoxGeTkUz76TlHkUV
rQFWv71r3Xo1TaZ20xdmMqsbwGSIPlDjYduBhBVlGbzZAcelsJGIdRvN8FnpBzk4
QD5KVGAcjPESwrbIaJu+CQ+/RudIc7V6oNxWqOlmepwoyLvsYFbDwamRUbrgmCZE
xe8BzxJAw1yccOwN0TLHOeH3DCkoIbfuunLFnT+pRq65xY0kNeDEOigjNc3N03Ho
AP+crLksZwyezWB0bNBuluPBbmneLL8kAPt2iN+IBYkUyqW1gWnmbQkI1mpyEt9o
EyWFvULmzgHimLn72hliM3cVdXPuWZzestE3jA1+ZjZYrS26TQVtRb4+Wtqn9QvO
Etc1M4BYWm1az8jRVXYhZ2UvN1c4BvCxI054S2b2scRPPZlDcLZMlqYJBzGF4Nkx
r4t0q1lw6s4xZw9J0gLYxzpqOMOeJTrIdZslKwfetWR44HKU1GuboDtCE4EBHyuJ
eqyFae79NwjHDktteL/jflKKURvjEZEucc10HgDUkPhrFRfsS+v0sxz029URiQrd
EsUZGvEyjiB9ZRQTC7d8Yjx3bgzImahPYJQCnrRjIALvM8zKLrT5qwvTh29LujKu
xnvkE6zVOk3Q6i64LKYtlaxUV1jQWysUos6z7D+9HwhqDeVRDitOryAnR5Vx5FRA
yPU4tlr68PZV+PQMOQGawHzYogCDJ4alHxLwzOqd9kb/0+HXwduP24XvSBy+EDq8
SiA7pO+AHrrWgwpb7fHSW2vTFBon5Cu+sEsezhv3opOt0t9fV7Py0ZScREfgytZ8
XDs6HvPKPhyBzN1PHEXMh5lg81yMiny0YkbOMOlqcshYtjN3fio0sxrL0T71+N9R
ksEYnVf8aA1papUHLLZHPIe1qXwKFc6cziuz76lf/anEpDqDzU6GruDoxozGpz/o
CSwEW2Mo7Kf7WPFQrFI0tmt/R6ApCYyJWJV1V9Deh11elVxXxBpmb1p04Amv0CyI
8yLUIy7MJiEdHndLNekzurMsueFWwAd0NaaZjMzKraK/VGPLECwZdnE0HPjdnZeM
cXiR/0xvGz8DmBy2pNuLd3VHGNOW/2KxRYfzv/ukTzvsxsVHT3/bidSzGP9O5pqF
ErTuwfWwNd22mPMlsuhhGE9lfEG5rPvZP6nIK19ek3G11L2Jx5M0brLjJY/MYHNv
aKgDikfxw7Zit0EaKj/7VuyF9BrrTlRs6V6MD8jfDegYjXRR0O7KwEFgwYzs+zIY
R/6PYJzX1OGQe85i8wG1S3fMxgs1gBvzOMF5YlsL3pUNfxyBkmkiBTYa040Q4l+K
GQpQ/7Mwc3xJ30RllODMUpoJIpuel0LICMUHX8DJwZiZsjDY3iDpg3HryT3SrYQh
EN5ySzs6uhCI5B9LyihV+22ZfgvhNy+6OcSObZre2D9A2+OtKSGR30grpjjN09B9
MUEFhPpEbem5z99X2JDFSqa1hbu5a/7LePnIM9XvY1yJNRGXQMcIRwSY8mYb1+lv
iwhsvTO7Jotr/CRtR8tYVwwqdtAQXXwuHRar8FTQ6sQxhqUCHF5O1D78yowSK2n4
51SGxKZthbHiAPOTsH/KamOMfT9gU7g9R+F6LczibHIz+/LJLHkda38QqDC3mFWI
s7gmzrPWzd5pSu3c3NLZaeWXLswZXypdWl2juBqpJioSNI4I83Jm4gInw8ws+Vyd
FwTwM9rRyAVxIJez8/TAsQ0f9sXPWlttIP6xzu9nzrxuC4/Wfnf7hSle6sZOS5eg
2z7eflhe4wcQxfZs7Gk3djdXRETaaY+33qzLkWnnOdayrVULVTusimFCmQEfQgHu
f9x9rwxNqo3tn3rTzf160e+9J2Cv/4q5eQZFuVMzwPleJ6lB0ckmgRFO+uGz65Sx
WE5szomRQl7geFuOx+KBkgAEA3geRH0yZd8gA32gBtv9kOv7xZq+qI2Z3tU+h2yz
UN3bQlfSL/nhTGPQW4BXSLrfhqn6EIHt4ZzvKisGqKfa2bbAO0sdU0lzBy3Ho4Ox
H635646MRTKQ8J4V3ZdQVULKmm94FRFv6Bhmwq5kef2mPjWYLzoVbOXcHi84gA+L
TBzhVJQn3l8C4jyWcJ92lrNC8lQQt/wDoPagxX3aWNxpnjpuD8Zj3RNGGsIp9gHV
30TpvJU+TlQD1y5LrABHfSYhrcHSzqf7Hj/qieDnjU7yXJElAsq4ztHwYogyZiLK
aHHtG4bvNcJ3HuNXryXVNlq5kiJctrVAE0a1q4UqdEYlcXeVQblm7ZBFMCN81jSG
0+iXv81UPWA1t94ceqckNSiAAF6AxqD24oF3vYlitzVczFM8llAEc5WKkclJZj94
70JEovLrpvzBaNkkeS3Wfe2/2LbDPNypRpZKGwJCXtUyyF4KuWQa2jbYgrvGJh/g
IfDHwPCD6Pj18IZx30D75zUtYl5K6u5ZsvCIVUAZCVs9Xo64ht+e5VFiAayyX6Ey
ckn4DqJqXDswPYsUb2dgI8zu/poIaoIC3eYGHafEERP9Gryx8s+cUOI9sky/0NXD
Uwx9aGposUQfG4F7bD79r0/5vBDNQugylwtcYcyHYRfuLbDnPyhvybn9Ufo93/74
4Ds2wgDKGcVv6xDjYpajCYKJbalimfTVFsUXlqDaWkA8sKiDZM0Y46WEiPTECFHn
wURs72Z0B720hyKr+EWk6InLrdAMVQcmPHy4hLK3X7IHS7VxW81jbf2Vs1eQKpRu
45r5XdkpKSkYoW39FF+Fb5B2C/GIc9TGJ99zQuShtloB0tUzLo4XCkDKmf3k7kOj
A4jVc2bEklgX/Rj9rcCh5W/0CJgzRG2QtTemewcwkQmHpnxrwD4JxMWtbHLg8JHI
cFOAHeRxIuyX9/bjMCn0gc43aNd+zeiCvrWHVl7O/0+Ws1EwRXYVzPK5ElreyX+d
AuehMJkA4impxA6+2uCmTnjBsSTO0vypznay9aMTrNTFPgAifBsP9W0pKxjEycl7
DIfClwkPSOPCByvT1ISdXG83+XqrGgObs4vcSOM/bmfNQkNQiDMNAuLbFseZ9k4l
vRz4gr11keAqDIuKqui6bnNgEeuofk793pf3A9wADSL4rNO9rcWMqnH7DVy967jA
MCIsAwsG8S+GP7CKFMI6AupVv7ZqXWrm7pAGeJjb4vHI8W7Lv6tcVvNirG/ahQ0P
AZf+Sp5vylAAv5Yb0Zu0s3vcgAP6PZNUmc/XdesxGimArRTRPOEM3pZX5Y7PkqIT
eC7IOcCLwIkEE9EFmO7jCRVqQO2iAc77QUH1uFc9N/+g5CYWyoomCh3p6ELNAfrd
RyMHYSGnaGaOO9vL2cXkXNxKd+0PuBRY+vBHzfql3wardLB0DuSwPzyYHOqtnjSV
8HQPu1WGF/FjMrdBCGZ6MFgT4I3VEZkCWMXO9DsJVVLiAf9Qo9OZp7WUbhRuuUeR
wu1HcEfABTflrtlQh+TAfSmOwiim+AJ0nDPqYHtKHkXE/EP6avYGatio44cAg2T0
w7GPfqkYGpWq+hhT80sdLjDoQZx73UvzbwQCntwxo+4b7DwUYKdrhqPbfBfd8txQ
hq/ns0rJmJR0LsGqwSV8jU9AhlmWyOqeukhkxjKm62D7UW+dHtVpUxPKHTEV9jPO
oqwkhihHBFkaxPeMFGygBiPAFqG8kF8fElPl9luJsXbT2+5+lHDsuSl80/mNHW4j
zgmA6yAOWW4vQYKlx98o/2TK/LCaHCBJeGrLYIFCOqGOuba80HAIme8P0uSjWwuD
QZmM2OPJFyLlmhwlmV/ai7ygN6pokKiAPUx1cMZg2oHCd+zdjF0/JZN05lZTaGhO
e2c2MZj4yPzfS/MhRcvs2+ict/Lsmimk3h/UkdAwNF+bnK92+nbd6AV1BhLd40CM
hgn+Kyk39yOrci7bjUsztgNt6sabpZ9hTPWT0BkP6IOFWoyBKWulegVohjgD/cQP
xDZPIlZBsTvBogfCcA3pHNUy6nNGsS0L339x0Gg+jDbHb0JsQ5NLrwrOEuXLsXRK
EbgewLSKn706Ml8F4HxIFQmZy9QPopaUCbvmSpidGoy+EwAkUmJF7xQKRzAnNGXK
OgI8EaRqQlctAmsUhmoA2FvHrHfCjlNCdJ3PexfDQomptozn2SpqPlKmPzwNxD7W
itFaZyEzVMM2XqrwA8Lg8NI7spGDPzRtVkObxXdNGX3E1cbLclmn08DNwDx+DElK
szOjTor6129AE6J3w6qCV8BIqYiL0+zzEYf4Jf8dGnJsiLzTlTeY5EH8PWl4lkYx
6g7yVtkZ9I1j/BShgoi/Ugug2+JtaOMgYyBbJxNMHrRfZaW43jKUa2o7gE2TlkK1
SOuXsxW25d5J6EWZzIOxvoeq09VQy1JOh6Yut1Eb4QTMT7e8UttHAAr65a+NJ2TD
YDZSaeeoJ+6EehTApIV/JBN/mg0dPNiiLs0Mr7p28H+3tRcIGDfBWw50f4egO/yD
pY5YDVPRvKAbYimhhIKSZxZ9/8Xl68T7lSzEvqz8i7rWN9Vtx5w1Y9QxzLwVjCMr
SsGbRlZSIXOJANzJdayWgvdghItPb3xoCH8y18sztKeajoWDFZtwi3DylKP3hc4F
kR2iSiGvQp2vwcybXNZYwuRgIo5gNFYZjAuyDWZZwMFbqGMmE7GRM5+M0KZsN0PR
wVqz2AKXQFkOrC1NiCGxsb7DwZitmHYY+ns9vE/a5OFxHTk2ngv2KOsbIWIr4EKs
Ju+cS+ijRUw0Wg6FJ/eJJoFJNE+Gy0yAviWRYGsOc0hSqEEUNIQRP0TX61ThtuwN
y+vwMa7zManR7j6bQGsRIsEPnC96cV/u6bLpJvZz+RcxXlwg+HpdfBa+Vtek1LNB
VQNI2kHX3t1ZTv47ewTMKgbIua0WD76CqmKsUMCNdvF4S4OFMenzW3E8qKEoXpQ1
ITVid4GjTeQws4gdjAzpyPwHJEVHAW+a83spT5iD3+hncJUgE5wpZVi9Tg4NiT7m
yy8mry8zIO9nANmjjQya3undMnciLEiN27lPpPAk47Pz9jTKHNa2dNtgHFFHmibm
w1rRiUj1dzCWS2oQoedRahvj7ReMqGY/2FTL1JFp7KYZtHG8Mfg2Amw45ENH54Sz
Twa5oF6bg1aKCIEC1ulUZqc3pm8SQ0eccB5slUOz8tTqoSku4gJBbLZOHzt7ve94
Fl9kcwitB8oJoSM0SmDtokytgwceg4ll6ZObu/qOmpjTbk2MST5zim+dKaGdT3Pe
rgsPU489Zgrkb2NjoY+Zxknrgm54CWr3MEumKk8uc9xClRwmXUyuDwDvTGUT8RQJ
KSStJResMD8m6G15kFdGpk1TBAFhAGTeA6iSP71h2Zw7yETI9PwPYnc7fzy4Cusv
hX6doscrXxbNLkz7A+Jk9utWr/ZBRRSizhsZ34tKzCkOHwrKf05mc05J5Ldr08pb
YPwr076w/lFrqbudwyOfO1stWHcT34mZ2C9Df8z5CSIHcU1APVhbnIvjiWWVTkW5
OllDVGCt63cV6vM/umkq+UeSG5VpWcRtDkDyMlzkIx+33HXW9sM24CTwIsvq3oLC
1oSAFwNvvVo7b+IcwEqA+br4h0ZkKLYICck7LLoxCDidDJPXU4RrdxMy3wXcrfbH
kxEfrNe2W9tUSHgXwxiAvy5lfSWaYB5MlY4Zt599H3ojBfSwwqdPTnWZQbLYhYw2
KqJPO4t+M0j3MLQKaC9pS1ARbJHzBvtGsUVFwpxA+El6bzXfrtQ8R1WaT4N8yMC7
Slm/KEQc30ZfjBAdj2G06+0/3jKbL+O10LwCr/2sd4Kb1nzNbglKF2P37Nj4FZqc
pATo2wwGRlKbVPLb11K/gkDeFo6wQRe6lk2zlGlYG/N42JQd29vr6Qb6fheC3DYt
9kvnhnBnfBT4XD9qCBukAHbMvr7okDnoGbOxjvu+tOqLphLTY5J9WFX1jXO0Mqih
YI0XU4bxJx58cXtqZPG/Zu2PP6VYZJbf7rr1mlGKCAwre3y8zRgBnlaFFbiLseP5
nfSlDDZxxt7J9E3JqUuYCROAkan0PQ78tr293Qa9yENfu/dpzOyhRq6ajxZpzm2W
qfEsO8XtsEcjFcWqB8KM1PveAucMk8E7SJ/Q+6T6euut/+kULjO97Zaw1yEjmgu2
78YfHdRG271BsoBv/ro25PmdnCsfh7P2YmCBoLUlgTdgMqqh9tzovRm3ps0ZeniU
UdRjo6AROeqt8knau6Ay7f3zCLfoLl4lv6z3kdpqPbhqjI9xTFAd5Orb7YrFb9xR
wFT2oymHtDheBHC6A+GrdI+4CKQZ6d2DmCQFjBSCVYruckUUNsgpOQhcWz/aS7Zg
fLc1KgvJyjThbWQLuvCiLBRqp/iHAPX0rQzmyoM9yxx4f4kMdYFOeilXk+j5IwLd
tU4JPWfgpifA8D+JTqUihxR8NeUcqgXQPA5sJ8SpOVLerM6AJKg9GoLf0Hg0112V
tqV3Km/i7k1Y6CDZuTU869PXqzg0cTJhhl0hjzAv/82UuKty1VnPcUAZ9/zfy0SO
+bRKhdkioYZW0tKqMmjkrWQMoumZvkej3jrvzAx1m6VXZzf6naq1OataPAQRTyH9
a2X6aBlnvC8niGAVSaqerRUoM5f19Zgr9NnBdz2v6MOAvXt3GGmaM/ueeLS9y2E4
u0mucybSt4URGCPps4lSmHq9ZVdFYslHkJC7FTRgQNCSQ+ZfJ7qDqxi6f0jwILDF
pzQUVfItbJ26xe7i97egYOr8NaqKXwOjFA4FuYntIoEyVDn3juk04msi+IapllM5
GTIxd2HVrI5ciHkvPXar2ZU8przAUVSDtz2aBB1OYWZBMe99zaD7Zv7wGQqquExy
QQRJEHgtf7oqSjF/yMMBaNc5M3tCrJqGpZQSIW3To1OKGVlF6m2K3kQqDo/e/RB6
Mwleda5eWcRt9jzdEF9R4FFx5ff2Nj4BnhobRweL41B5/WvXoy5dOhhk+iWAl3vX
7/w0LGLJApQGHa2Twyic4lzfelujuRt98OfwnIUre5P1NslY/pcfE2J0QuovXIlu
LcSsYsNvMHI3Gjegs1Ya3VBXX9R75e0/ZAaLTIe5BsFHG+Whz8ylIsSGOOpLf+fs
joT/82P6dM3U3Uz5vrGoOOsEIENgFh7E0eMpbIUlEq1W3enBXLGIlaO0Ud27vbz8
wnfC8v/N4fm0Z8ydHJ2ern3x+vUsAvN3AUIMfl+eNCH08S1slMXdjOVW+4zuhaWC
7hBoMZB737f+93Xy8+Sy+Fdr2/nYADAyVxrmplTk+VOCl4DUe4Ak5CfO/W89ukh3
tOg6F+BQLvFle43DThBoab7+bEJxNM5M2OCdhxd9mGuUpc+HU75qBpYRyjDJVtx9
iiyJhrQGOF8+7Pfbl/5PVzRirxZI2TBMRyS+xDHqeMnOrepfiPFpx1OGa/Eakisc
oP7+8k+/3IuYguAw3cl1zkUVVxNdHARlx/r0UqosG5MN0OxzBg+EMS2jhMuO6m49
OtYiXlchQg/sEtA3cmuCYlsXEzd/O5coeWNt3Rv/aDKia0zjk9Pd0dgIKUhOIHR+
As/lavTWemulQ7zoIvPMex83nJQ2knftvMaK4ELQ9jrp9NueBj9H7NFN2MeKMeqY
sXrhVRdcNmPlfz0f9HNn5/fDOnuM0XMfhWQRwTFx6vjkhIgRPCm+EsxYiS1zCtgS
MKbgCbeBT1Bt2/Lie37c2wlUB3oQGm3Nb3q8C0b8uVXCg3Pwh2EwQcmkGX8/yGli
90xpADtpAMlHNEHbBXZ909vg7GJSubj1WkkOQYU8lpa/PK7dgHHDsXDynKiS6kEN
rZaEvdyF7Mjp2IGVKrijD3o9Zpn6Cwl0uZTv+dur77SXr9WcFphgZPKcP+Cdyi+X
rKx0CCr8oCOBlX4CIOfLVRfibRn196d+4NNgbEYXPEkOyCxa3pWDflKo43ZpMqOJ
m9jcJOXPFQl/+9ZFIF3lI3dtiZZK1AfxLbhbEAZWSAuLtDr+m029HVsLosPCQ0ID
F8Dq+8piozEPjtBYfs2/UZnFxwaZsPSXXrrnx487pEM5WY4AhN2hrdYvZPry7TZz
zCIblZ9xmCgIU4YYgDlgrX0b7TJgj85iXQABHyorvw4ypn2JnM1KurjACt8dzCrm
3tPi4TWrGbT7baiTIzTj4tU6LZtA6yiqjLuSoz/68KvSBoeF5n922SszEzHUk7HC
OBap3p5MLuKTRkBUyxv7r2LvlH3sxS7Q1FtwkHJbyxyfU7VI+hZCUHmnPKdUbABd
TTMis4u5W7U718bx6+1vQr+Jp8TeIk3rvvQhivwRMseUPvYc/wCFRAreC3kiMSNX
ozb/6TW2ZUJGt6jVk2l92QjpG2X9tw1/cefwT4XuJ6wd9IIYKDrOSp0X4HzffdtD
ac5AuHrY75CynJOI4MaDJHPxdSBrgh3MfodVpHaKwyHw1H+UP5pr7RX8yItCnk+6
egQP7+6DefxXQrlW4pxuq2RfEe2KPCPFHaOQX3bdQbQZX0o26uaa4MC/hyx4C1wD
K/gDD3XjNrmL1XhvTZDxNYF/gP9OdpatWcZKUkVRjPcorGQN+x94ONpFZJA4vez8
9KtnPtT+W/LMwBmTQktucPBCIb8fJfvThjWO4OgB21XxHYFW9pdDjGuobJpp/Hrc
p4/afRxKKPvBOwDu5EYHpgXrxgzVZ33VMO/n7z9fzVDAbXgHJKwtxsMW1c6Tzj5k
XbGLSuzw6UzCfpuWQgWa6brTo5Xnek7v7Ez0AVQRYdpc/W3UjtvALsEhGIBLo+oX
qVpJWbKgIwirId+3h4lAqMaZPcgEAjm7hpcTb5qcYu6jWCgZxMLaGvXiOaV7zOXY
/M2Wp/cit3QvagTx25iZEYZHocDMixiUf/d8KzsFN61wNXrd+xSC5ycL5sYC9cCz
zISdoD+ysvKQxbYSwbgR2LMRA8oBOy6dV1L/mNN+l2fUcRiIFikD7HZFSmSmzPgF
dBJar8NEjey2QgObSwSD8Oykh5Leq5fsavyGbAKFMQx9jYkK86CUoCiylTBwHmL7
aoswB3ITEQh7yTcSc51FpK3Ry7B3j3G2xpu2G+dhMS13nfuINqEYDDEGlvIn49Pb
wY7xAp1wgpdWRrOcX/UFGiZx+s+fWwsyQ+FqlBWh8rmXdSmeVV2XB3xnwlo6fPJl
1LkfEqzaXoYMpfi6TrHRe92XDYOAI9H33KRoVHaBqhe44TD1r8bMbrvwST7or+Sh
SctDCBS3U57DLV9fz7wA91TkWyCzswTJeEyzpxrwLqNRnjD79C0B5L/CWnLa3n0E
4Ab0QoPtfpYvMGmS5dMzN40swDdUHLpEJTdl8Aw5lW5dkYHzy8p5IDetxiKM1rD3
+KBEGpVoqs315d7RA5AcS/FEzUgo7ir6fcqyjAHVNYa4xmM5MdUlPNrRqPIIjIPT
bjifn3t0smwBzWkArsG+B8nZ4WW808GvY9K+aIhCzlDdgKX6E8C7w0vhgyOdspYm
7ek4qoiK6NZ7qYoNTq+t2auqncP336vW51PFMFr/L2c9BYrJr1SS2ji68leru8mF
Sh7sE0aZu8tQfDXWM96uib0FgENFkCU/rSgxAGVEsnPXjM3TdntbYFXnAM8srJ/x
oqZd+AaChslFtpg3nM4hGd0l7k7jH9EqFS5Js9UKzZxia0ZMpLBg8riMP+tyuv/O
8M3/7ydW4UTH0Am+EZKUPraFxticA8C1Urs4bS94yapJHMtieLZB9ZS2a5eMveBQ
ge4K/NbOrFLnzx59N2H9/+1X7u5WKLgWYv0OTyE8uz4WczY8WDuZCyrhRXTvsKh2
CnefWFsoRDhSze1NYdlTRbFBuamKFCjX9Pvn60H1s+C0pW8nMKvW5C6vABiOKWBH
qq9aAqfSqw2zocmgyTkPaS/64RQv53S0F39Vt9WKVexccbdfSUDzRo7m5e617Bf/
QgCdGUAeUG6DE+jz7a8hI5f/uBOJH/KFM1Z+MAfNJMPufdy1VCbh10lFxuY59ZaW
N/s5jVo70ed+6yWZraB+W4Qpcm6HWWpPoEMEvuqjhc11amiAIo4LCKw5WuYGrzBT
RK8di0hNKzgXsUeaJz6H4kM1VVGfnptiDbg4ef42xYHXRytaRzukyANaKO9kDC0G
4FwF8+UQwMR3Ywm7ZFQmjwPJ/KI6CJUJLcOP8HybD1m6sPAOCcfXBvOBsuVaRk/7
+9L+n2wb+mErd3qhNw5rBkBEW9zUUApjLoZlBETzxZWe6aZzRQUU2/KC1gPsyLEF
ClVCXZcCFLgmEGdvBmAXCoRGElTKtXTEgaODWwsCHHw7NdTE9t9ZEjLu32neE7+m
PCyBiIvHJFQYI51YFKEEdECKtucImed0nhrVDbFmQpygAU/bf/+A6IC9vjzqCfor
Iwp6n9AtAnQ2a8g89ouqU+uQCrXB3kUVsnqjivKpjhlogoJ7VW2UK+jqENNKfuHZ
1iXdpc0jMT4VLC89Q9HQl9SyDP5WktTvNStLd/9jIgFYhWBdDbLtGHzFKPK9fTsK
iSeY0v6UmY9NsEbLJA4oKYru6HD9+WzkBhfbZpzeesKDnhw+hzRRB7fTxs1B2IAt
Jk/0RrELZnS1wKiBbXwgXpBWl5lqyPK6un6Cs9XiRBbjpCQ1vJGykJ+PT4ynmYLr
V/qGdTjqaCa48kM8ZHKXTPuChwTRPuVWOCoHG+ojR6Soa9/39e987WBAUefgglzB
h6P5IzFPaDnH7seBGMltvHY/HLlt8RIxnIHnT0FstZ3u34KUZlAyy2rRLF0NIyYV
R3R10HMvTrtwc31HrzXhXSlwDu/dcVN2dnzr3OUdupGKXh815q2VV43myvV1VUhK
YuznhuOxO3KeYOwulny9lpud9d7ZzvjwIwha5SKsk2F4kYQh4SsNxUJssFzmyHAQ
0h57+IlsT0R84MPKdEWQqnitWE01r6q3KaqucUoIjkEbCS/7il+fcwt7nAOkKMKK
pKvGr9PPS+2DbEfH9vbXW/rwVgg5vXNP3F08v1Q7V/gceCPEg6P3sd/uBbJyIRgR
TFTqSCrOeJT8S6Uie5/lXmSUyrw6YiJp+7M/eYBGELjQvZm4cyq7EsmCsMLx7r+z
Skpsoam1vySKJsn6C60dYcG7k7s/JN+a2mAqKaprvLV25tamqSM6B9flHpn2jLWu
at/q+Q0Ae0tzKkj/aKjikNJ44gDMbe+K5Q/hUO3kuBtptOTFWYASgQQAEBNpZweD
PkkGgoT5Nb4H4ICLv5XREQqeYxC5+1ab9sq8F7QhV4sgUGySCwPbcVCxuZGHQ70g
rqM8hjyvbGggWFW75Wdrs8ffNp7aRQAkeN26U4JaKCKIMwgRnfUlwg9G3EzeWN8S
eb1Hs//GD0P04KrPRVRplkIwXAKsf8KbQdFv0MwgNZN9UPeqHKUsmptb6m0nzzhB
VOoNvN5T6XaxIIREsM7Fu0wLZPPyQ3K9UwZ8jI3MwqyKlqk9Z/zeQ9iYrnQTWLPp
enDB3aVfQbaOYJwd6A5KYV+HAJhTkq/vVCwY5e+vphIlkTfSrOPsI4Tgk+Nk/0Gf
4Y3H0cwadqPKV+pJndNZsJ7Uy37gtwQeLRqAAu7kAtD5L8mfGSpKm03VPecHWpS/
A5fW8cX4aIhy63a/afHvhPgiu83X3HiRto64n0vmrc5gyBB//YUVawVfiqg7iK3G
oa2Yc1iJ6gxh9ZJREF26FQlBY8v8/eSDGx/jUU+NsvlWdNsx47hSuci8SEB1hDwO
izhHvIoufap7qBXVDJaQ/++asNCQ+baBt00cOjC6KKK16cCButJGuqx7aoaVBuqa
3qzw2Kwe8gq3HZJUFveDWR+6V7jd/pYWIATFQB6mcxRXMb330UBk67ggpal9hLTY
NVQv2k+eIdJo9vTqRA3FpjMgh50/LycTDH5f78XGBCBdG++Ih2sGPsuiKnCQpNCO
3Uzprw30GSBJOTodCmW1AhHiCVfD++yiqUS1sqI4h9K4qHLT/kTBa0MsqPfOVPX7
Aonj02K6LS3ganr07S0+hnC68v6/Q7sLbObXDYllBVvgYGrrz8lKALuQhIEe2p51
ND71fB0ORfOP0bpRTXYInf4i/vukddMS014d0HPT/WxA7RD/MSSKbLNGhUjtEK6U
nBers7pXQtJz3pz9iMWZOzEAlKPHbQQdUvMacCiU/om7UzCQelB5t0LyhaTQhrCH
UGGoARmLmzu0yfDUKjDsuM9pHs82QshaRRF5wamPJBPJgbuSv3sgWByjVfWfKGOq
yA39o6EnsUu3q0ej817k3KqjOBY+HKIUvofOt7IsmoLTk0Fwn5W+J7r467kq/SwW
+d18hKlrfjWZcs0eIYsFJxNtYcMaNQXpeEu0QjJAg21y2ZVVi7oHkxoW0ZOtEIgx
Os3REwR0kSl0v5TVdnm75zroRYCV+JK6bA4y2GSJAhfqR/ynPiN6QTLoKJgs46LJ
beASNTFFBxjCX5ybwWW7qI3+GcwHRMP0AIZcO4v/DSwxlG9Z9g/AE24jPJ7M89Nn
k0sfrkGc1FSGijX4jlrY6q0gZruEhdMGz70sTM/ucrl2V1NWUbsavpGXVCpeaCIH
0hXpLykDHJORcWCabwp6dhWXta5sZKtCdf8ChXv3Q2wZGEJSSoW4aQz1MQ5n22aa
jmCQhQG7+F+ygTyWkUzYWtecgT0z6/DVhK4e82addiou+E9NZBg18qgtNq7e+p/J
7U3/Pr7EUw66EGVdWSlZQ5J5yKUZ7j4vZ9bcMhMzG6O+LqZOzdepcuZNEcBOMXyV
p6qSBX1envX39XYxcisMh6QZ86KTWuV64BQ6sK2xztUN3SO01JEYyMkbG6M6iagx
lyPCzQ98zPACqKyGMC73tbALyW59q8WFcm8HB+I+Azq3TOs/1RtBwhU1wbAxjAGz
bc82HYF8x1JawBbSB42+kz6FPC9/rWznwu+GsAkOpLTziLsJa/3ebx1q3PyXMNhX
jp1mXnYAEx5iPxQcuVTs+DgjUqFxdQXn6Flem5DAzwWUcVI7BvU9BhWPTcBIysyK
IBCLZh3B16uq5+ZMzDK3lB2nvoeNGFELhSxLVV3Og9OtDcvWqjwZaSWCHtYhAHut
MmOE7jbZ9sGF89HI1SmmDj31gspeDaDlnwc3PO9x9UeOTruP4rQIKqZ+o2hLoikW
ugtTYzLWtIloJPyRk48+lKaOizAENltbVXSa5aYQxf3OsPp0Pa+GTxRxisvHRdAC
FPF1qgF+QtyFappMdrIPljDwHYuzoPSBwOW20S0Vf5K8M/paMbkmGU6l9jZzEa8g
mm6Ql6FQJ4h+eUBLE+YNAhh6Bv1NaV4hap/fsQFPanNknapcs6VOw+d7gqFTeCKd
u7oVDP5szyNJnqx0seLqlKZUK8oK3RVlMTqqE+at6EttK4YxmNxPEy6wQsVt0iJy
8bdbUQKJYm6uqNWwgIlQ9ReU3t3st0eMSuMTw7tFPN4m/jAyZPFtFZOy7BFRwMyr
6EZIAh8z6Wa5lKIuWBQz0W+BGBDUwlvVaJvsaf59PPV09FTQDgz3GHGVh5dFctIQ
+/zernE96s5nUIq203zWKZ7eG+MoXpjkpDjdTIyu60hCkHoBcTnmHsE70l2RAV0R
3XXSIuCVl21t5ye5aOlA0+e2OtMEbDtyizohxT1F3QOLql/eyS24Vjc0NtbbBsg/
Zm+y3QSOgPl25+GIrLC/KZzjaYYDItIMBvLdH/Zw9NA3BTUIuZ42jnMYs5OP4zzQ
KDJ2duDZjmTeDiwg1h7ylrs6j6X2uTqTYpEpnIe1o6xjylOuOd8r0bcfVkoswk0Y
CPU94cHu3Ip9LIFG9t2SDwwN2Iz8WTLdWKBPGNbx3LTEBbJi9gbAQqRwPfNQQ7hC
py2mOH7r99b5XYARNmohq4YjEDg4orfc+X1LM/CXqvFILW3uFBBGOirtnVna8OAH
zyQbknPpeufAPM7qX41oCeg1dA9Q5eKZ+nmd4AWFoqImjBj4h4/7JxiO5+ebq6BP
lBGMiW6reLGgLRTjZwvt2nTvXUMoo6pivPsT88tfELFzzdiVDOaa8IS/ZVzZ3vDs
B74z1SSMp/x1jgqYJZkbTa5KKjfV2GxxXnMchkiUYtnhfRMYO5hmBmENcDRY/TTQ
8j/I+GiTznIx20Fg+dj+7RRASTZOK8lnkKzCSVtfs63/nc/N/4TcDzcV20JSnT8R
6EJsxTToGtwKQFzIKUjE2E1xFd1rWE0x07aiL0kOrdnia8gJ5AzoFWkiMqsdfn5g
F1w1NHKHLV4+ItW/go7EsZvIqyZhuQsPETe7qY6oVK0cmu/t6FHH2mMjHjcMT87+
wtgVjWYq0PK8z3ih91HdGzaoblXkxhnOGhG4A1N82c1PQ/IUTMw3cQqtvvUthbff
HXf+8ayRwvlZHErX3e6uLA0Y8n8fhfqzJJzbqwvCZhS/kZJHsNePKJioUsgtkxur
GEuEXL4VRjR/y4R9NlJxiCagLVRT6dwBjaCVVrsBB4XICXf7h9BHHgbT/Fk5vh33
ucVZJNBJaUdHgomEqdnGsKZB9fjUDJGy4ulfchtrx30bQbvtcQtifDClTZFPox/+
hC/bEk/VjxLu6wBG1ItNJf5aNqW9VRmedSooBWOzo/daIOoR7PKnPXWAociBF3i8
RDHK0IURVmaRuxnUWR9sq9R7y5qYHSWNQ24/pDpsOUbT1TM1jYik3ya0dvLHutBG
5iMzIoBEW/P8RwG/wPQ3wF4Oz7d+diDDcM2dRHHnwTbz7Qb2f2B4I8B7rMttExNh
OODkgN/3RCtktckqrNVongkT9fAHOd6jbRym9JyTLYot3Zt6xbW79Hz398HztJ/0
mO8ilvuQ5qD0WO0q5M5wLoTqmP7KbYjPART0f2pppqrEFHobMyAPflzN2QqPYhEA
bX61VbhgWwFNePjrio9klQSOBGimRKcs67KaVotatJR7fu2uSxYusTlaPacRbfbX
hZLizbnTKzLeCCWVRpWxgNPETpoxCFvjsDek8tHl6KpLYtCx77rwlGlBLqaEaNGP
BI2+iEfKDyvn0R3pQUABdZN81EYEmTY8uhXtIgawCb05NMRw3F3xWfArEjbG8EJW
A0OrJ/MLwsNm7VDx1w8q0ZDZ+rAGqSHKNBKobx55y1m1PO478xped5a13wxJeHFl
TOP1VeLeGYt0pw4w1rdXzBIfeyOptbhOCiLXwy6Y35hE27SOxWveI6XNouInR6g7
7JD5fcz1aytADXueGAjOP/Qkw0SqxbZC9JkAIGQLabEaJ4pRUCGpEQc3YtkMT0X2
nXEf2IlT/9g6/Q1SW4pzi9wCUVA7weZ2hFr9Dwgle5b1rNqKw9JWz0fsErrazpks
ZXGqxpdyBpKj6zqQmTURTBIfIusAPL4danekwp8IKCB1lI9GSlFC9m49yQuo8hdh
RjazUi3ogu6Ohab+9MldZGcESIiawEeEtol6nsN1Xc21EEhx4WLO79FfeKI4YARG
iC0lGZHluuZGwj3a/kB4x8L8GLBlsEExHW+zFPJzySQpmLv9MVulSLucPoawk2Dv
CEHnFmm2nJRDGQbJqalk19py94QXm+iKuD796Knqmt4r1iZLcbrUk+lfRQUGb/ig
Gn78nsydEfwDkBWZWGvuHUz7EjYqLW1vmVAD6ZYnd3V/FwdBlwKHtawec3L9g6Fx
hfGssWm6SqCNj3LShyz4vEsIwwAnd4dMosGFnWntIpCUTiDbB0Afs/3iW/kDeNxP
/YFFMVEYZAMtEap9xWmycrH0066iD61sDJ6BM0SuU1kWmYllZiwz9rD+xSbrP+Sf
HzANVU3M4keUoCBVF3CfF4Op90kuxJuTDaZgHdDLB0C3uD33zAJP/fEQQ49LhERt
i9FSLsQMQ5WTuNiNTdF/1ztItxaeTcKKwpk2A4N7zzStE/kehywydjVnEv3b1uqO
kBoMrAuzrNPbyzYPA/JrKBCUFFpHua+Z7SHOBn6JHwvHcJWY6OJVxklMNPen5q2R
7PmDSCFEP3WHAGKRLqU+A1xhgIboGOrzxWCecNs51me5Q/TP9MhTVoUYMIbxa/6H
EqNuVQkgi4pYUj8zf9pnJIwKWJNHWudYkpRvElQvpqATwTq27Ci03CCSa1HT4Mp8
QVrhVf3HAu/JdbXvpFeQQzwE0/1WCko1VLptLMlKfc88IVw61nIuaGIjeP8fRXfR
aRUWni0jVYa2cNKMOqmX1pLBzrkefGkNCBfbwBCg381KxTkq9nR5TuPcTluwHfqV
IH5xZMqa6b7bApG2w7Ki++pDnMFJ0Vd1LNJlyAx5ly07W++D8KeoDNEQYalh7Zuh
C9oWXHkEmc8Rmoellmnsfr3wd18nIIrrOBR+fuYYwlCO4MwWYprOnt6yHwTiiJWm
CevHhsvKn3GyxUCYdNTA6BEExGmyxD8/+1gUA2GM/zHb3k/9qZxSehW4qvVUR5/O
HF/lF9ydcXDLN5cTNuD8b9n9E/9oQt9EXsPL4TQ1u0pOo+d1u76lhRblBk/vXKjr
Zry+97z8SUPXg6VSAyyYBMLLZnzMR/zIwDYLRwPuneWCeAU8fhxlSo1HSV0IXqfD
Zu9rSP9g8mbHiEhW3ZgLoG2iirV4kJANRQ1SZjfrW/lYL/g05S4QWdBPrOm1/u6w
crQNQJD1t71Doek8DDkns8WfT9JOdlkHQiR0ssqJKQ8LAobUsLTZ6uMgLC7L1ySL
EnxL7bpywfQkyYCCGWoR40UIbYGmqM5lTywZErbqD12owAKVo+qM5XvyvkQSXuS2
aj3Xl49aqEqr77ymu84wDZk+nVrw+t8WCv9e0Xuqqy2bkT7fh9LL67DsDaas2GU5
LAGGT9u7bmVqdFoJ7bhGI+e+Ade+nDP4U+2GDEqoMmTqAodNVR61QYA/Pj0d2y7s
evvIMojwM06G5AcsidOQG7T6n5PqOqd06eAcXEERK7I5/CPv0nol9FsEpqvLkqiW
mdIC0n1P5vOh63oTt70OYmPLz084IG/DB+/TQ3z1nedSk9c05lcN/q9+87eRoIS/
KCY3XEzAtzUYHnPeyNWdbqc0IYC1/EWUgUk8kAEw2WCmOBbFK9WgP+6xpF9EmOXw
n/UAm20W1A+d5LF+pzKE9VFwDWdQxgSFa/gzP/Erg9sXw2I9r07krM7/FoLFbEkp
+Rv6JJnEUpM5mMs7lg6GjJG1MAhKP4H/Mx3WXsnn0NdM09KtKdx1Lj/GwarFSZFY
RQ8TmMDrl8KZB124dPx+PZWYXrxEQGZNIeztbkfhaEWTlV8pwj6tQJpjbSV5feNI
I6IbMaSvXSdnNZnfVXsFDBx+8MIExV3nMIaQC3cJZ5mySWqnREe3275Lxb9dafmt
JAS25/0gpUkQDn01+EhPldYyYqoVejhNNETPBMBc6Qc3OxZmvcphgUMQ0mxQRhqF
`pragma protect end_protected
