// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pQ1Y9gBpfQN3BtPUkOEAlAPpWNuaNmi+C3iDY6lp01RkwB3syXfITwCTKIhW/tnO
Y9a0HlAvMRpvCcXrjBn1qNjIBUYM5r7hdqF1ugTwQ5gtQohIpCZhn8KwvBXqQ91v
e/h38w9W204z41LVADLMCbgpYjK/FNDB7sune02Wkbw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10528)
dQEMzv2MpKQdOnj6WhQgu4JWQ6EHVsB+9uhbB5PzF2/6ss4ZKE/rSBTsnGfyT7/i
w4U3p5pRaRsWvNBNTdSV9xAjX3aL05SHPE6SgXhl+ATHhBZP5L4oMvTVTMe2VKQA
UNN2k4Xi+xpvvdHtvhuOrMXWuc4to/usEqtD2l04YPrzV/BHomm5RkDA1sIf9EWl
hoajBszEN5rcURv2rFSurnSXhn7ZRpntb/cCHXmqhpJWOZQWkcE7L73rbdh2kU/p
Yvk/w20J5+pxBX9zc8Xx/n5ZPfblPJTk+JbwnSN7mSavhV++7U+JEHG4P9Wies6F
IF5l3e5dcaSzi1hYE6QV+3ShHTraxBExy8mJYLzo7YIM1lZ82ZcNRWOQ7jUNVr5/
3CCgdDG0id9FY95qDONxe9tf8TMqEAM8+dP87xj321tesn7DG0qHW9gbvYvhBVOf
O6Lp+XZDzTNjCVZQRCe9MbXhw4CJEenwBGgnzM+tkw16zeB4Ll0dVWbd7znDt0Ck
jkOGZgAak1EY0DiK2Zt6iHubuR3oYd0Zunaa9GgwLkG8+JDAuqw1XZU2Q9VslWsZ
PDhdU/1kebxzlxoZU2MP8GdVEjOCsq27uEz+x2Ph3OYz66owZgIyi4auf0RiOo5h
7HM7FdOrlA35934VpPqs8F7c5VrggWxOJYncMlOLY4sLGDvdQ7rUubNdca24cKSD
B7835/fpjQaGieTDY3Otdu1VzUbave9V/KEXFEMFs3Na29aTEyb9nQowwPajUus9
i6TtSoygT3hixZpQsEm+iSR95YoI94Gnn3nlpHDk8WCxAupSKq22OKC2Ei0dPGob
ffgWj1CHYWNJTcTGB7iyYN81gr+HFmPPj3vN8ymBkSadi72O/f0WgmqzDyPL2+ee
tgjYmVBEblalYy0+4AoCrV0ci8YNSjrLnBgj5WAU3SM1C7qvzIAkMXApDHzrP0oH
R2wZgup9PUhHOuAWhfqVBASQIG09Y5D1/M+fxo1zYMP7XM0KC7Imitq451XZdhCB
SoIjEClbV0vqoPCr7ORDLnkwE7R+Y57RU9b4FzyjgWpIz3FHQvb+2e34eCZBKNw9
I1/xso1aiRqSvO+5D5E07Y5JqVFmWBAG8wOnfM6MnqXRM//4bI2ccmOn4M8nGhWp
no5GuWyx6kcbvbi4rFQ8X15q1fOT9MT4ar/QATO0VBiiea5JnTGsBob/Ego8JrSL
GRxEagyfhJVMGLnClJ8cNq4qriQFOdbbw3gFf8mGwU3VhapVnQsOp6Pw/J3F7X5P
14TMDwR6B4Q50FNaf9WQkBa10MlVbRKnlmUw6MHgoUYcogPyUPyYyF/PQ8K+qWwe
R8bpdwPUogAB7eSEWO5C1jBzHx890djKmQGJwZdI37fL/rO5FrKJXGUtvyzxZ2Sj
PMYakTj5LtpkcrKVsihF+f1ywljtkCgzeFAjJtn1mQ4eys1aDh0y2U/tcpSNr2DE
XVetYywZ4yJ8PjSS+Y4A3GjGLlsdI/YKunEpwA9B48T84ww92WCAj0dfFjpnJdhB
IpD6OtHKJxwF1BupeEE8M6HZK4bv+KhTVnrkpvzIWswO5F9YsPb0GytM5Y/Asrm9
511ZRH8vhAhzBC642wWX2SuwJzkLuLkS471nsAabRXAMfZPrSaCpFNYllDGQfMbg
BxMNxc/XRG/HJPWVDuMUWyPLK+gVE6BRKwROi6uxEZhRBrXicxpmm30f+Pe+2oQL
dXSxv/W7Mz/3DeQQuDW512BG2v2LizW5S3dAxqbLKlNCnb60uEjw3okse8c5xPrd
ibfPXFHo+UW6wp5D/MCdaEObxoq8K5iVqZzjeoGqKJjTLgabr0Mf2akTO0W5tDeW
pJzU9sdskzc2W5gYHCN8yOlt/35Y2xy6pZuLZCFVbXbVsDfcLBOfBqpbuAg7PVKz
FayaeMQJJOtcY/4WJEYEAqHhb3kMvjRzwaA3bACuofpWMfrk4bqV3vn59tWaZJ6w
WjX7FsHiF/fS0h/6MK4aFl2prqGhnlxyCYrnnVCcTxX6k9bSoUU2yBgLVBSKd10M
m15vNqx8OrONHBRTAGIxTEE3G6fEN4vTgocxlBvBc3fZqvlYdQBAG5098W30AEdS
OHXn6oP4JW2kT3wy+PpryN0QnHkYLldWukGNHEPwNwNooJL+rVkJDIImyqCdZkmn
2WY4coS9+hNkcFsTeB4VIFb+5lOOghntwu05B6HpuHO02SUGYTNtBWRCs7/VAb8a
q07BRCEeAkLQWPFEpIxvN75X7kOXdHKuGrVcmFUHZsVNoLZC2JI2cQNcw/8XAkOI
2d/M3u9/9K+laI/D3JaRXGhTycXTuRU9URuYMCEzH2r6QFU1xywkAQ2GlaMIIQUX
wPaAYOTw7KBU5bWZjKdJgngyhhyfnrXoAyOQPEIijIdS2eN+mQPC6X0YnWwfAQSi
ndNUup6vucw888JpSvzvkTxuRjRTJasNjfFB2wtEYmCI0AuJvCNoTnl5CkHAaBRn
Rl6vKJVvzBY6MfMhPszMIUMi2OXgFNpEHd/0T1QDm1wrQjDTqwGr/icxKuWd+xjG
/jsvYPLlrnEeZ7kwixTLEWQfj1dvsfLOll/lYSr7mtkVtAj1wfLC3wAImrKPIOF2
QrVL/45bNSl4AOlSJxIdqd6bN2MIeCfBs/RDHzyfWN08zzuHFQ2F4xQUZEOs123p
X3qRus0ZEcoIXUV6zj2mi/YL9oJYV25+TP0Kj06Q81hY506XwxZP4wzDXvCU5MhR
Q//N2he9QKCNv+LaabihRYsBw/xEcA4B2jWNooZUiL6LfqTecTFEGL2uuLMgkQyD
7n2WK2MrTvO/GX7FEQv6JRj17PpI2nk+xddaCJ+nyb8NK/rf4smBLKWiAGsu1ITd
s3pj42XVH5Joo3VOA47PRvkc3hHSa9dG+hDrdrw8okd6bBQ5ysTBo4N3yaDauFlR
WNwj0ZRtED9gAu8r8oplwaONsndL/BmYk8nLfFWDP8qCe4BKHnDxn+Lj63QwBC1r
KUAeiHHBallwYSt6OJsV4g3r+ApIaNv2hbDhSjkk1Kd+3WTy7uMbAjZLxnqC7Krh
5OCVBx6mn4hhf3Rbmtn9CMwAgi461xFvkKaiPHvB36h+40z3MhyzM7jjWNG59KKc
V9dG/rdEZRLLLnDQlw55dGDlEhKbVINFriCGbIZ4QiLe0qELYhUTbMMFfKbe44nz
phkDBRe+PeMnbyW9UtSc0YYknmgYNsNb5ZJc81Uul7GLjHFs6cToYh+G4bS1KOpE
6EUDp8PxW4LKHsMNQIW97+GJ8V8XuNMUaVZDIzoknSGkH4NjoRU/wQKezaHCV1Lf
k0PhkjtpYMivZi/2EhJNcIZp41/rTHy7VrKKwmpSnwFcO4MYdM8/bc+f6/hR8ELU
tIuAvCdWDHxaib0EMxqHfqD1/S4+J4h+hHQLgzCsra8r394XjKE61Ke10jvxMkwn
8jubc/mD2lTY7riQykjxROnx7x3uEicdO8JnGyfb/mRWu275EX3aKQleon6l/emZ
PBw0vR8JjbiDpogJq4W9iFdmo5BxYnkmXqsB7G4gq8Z4fUob+Z6FOqGScB1IOY5d
7qQHNCrEHbJDErSlMJBgicRWpaTSyXmNaX9mBOuin6rii26m4ScQt92S4rUgCYTs
5YAHUamTrRn9VdXnpW5yRzmN63dwH8/vBQrYcMj2qNC0st9c+MVYVTuRESrDpk/L
EiIW12ZZG4p8/2xayNdeI6Ci2rmAyggziDC5RdgrhgGHd3aL901IaqBXZBgg0xL+
whRfTE90GXh3IKf5ZdliutziGCA8c0j5OfS/IrvMOshHzdxJtF8BLwLF6rpaZgid
p5xJjmdQEdUuXBsyNLsGGx86dAW1I+pug1BjbGbfrofm+qO3DmN231icmzt7tr+y
7zKxYc7miNJNTbRK5RHhaiZ0qqlv5RodbhY3GShhCCqk1jf8EXX051KLGnSQnRV9
ob8KQjb0jaMWyas9aYRf3iS3tlXHWDKw1YG4y66PM0AiEakfh3TvL8DC7f9SrQhq
aWidZd1DIxBhu6EAHfqLc7ZAkADu/MbGufQ+oUNwygWiaT4pV2/srks4Sg7tOYLK
IRnpAS+1r1KrTU6A0qkZSCqKjew22aQhr89nV+4L0RvXfzi3bGeQTTLAuCRa+kdB
atQ4OLw6sc6kui83q8b9okyqI7vqoOALd65MN2DhdXAQ6idUVGlJ4z/klJktlVjX
MEnLtwKPfyzvvmB5Mqm9kWrSN0X24CplGAfEYNLluW5Q+e7kq0CmSlUWf7U/Trv0
aAt1+ab9b2M/nBT9H47GMaiFj+YfI6vIM9IxAioOm1Cxi8+s4S0Q+91j03JfJNZH
/H92ZpCh9gqJPp8oncDa1OAaFXeJQftmykqb99O6OpegoiqFBe7FIjtE6XKouUhd
HzFtpFgSWRmv/lsHA0PrfBqAvThktnUI54o9LegBHX6sRnX78nn4JyQTVk7rXVio
TE+7g8f/nOe//bblRUURGb4Pdu4a0OOkV79nBjiHMew/jlTY3dS5GyLp5qQUoyTa
RpYXXj0NRBecwOQwGAWT+ShRTKH1+Fn1qC3GnXQJ4ORdFwJTd6Q7Wy6LtPJzDj5K
fjNhMRy+Yw7dmKTJto7BqHsPKfSrbG4hAW6ZAjX8J5IVrU9EyfN1fYnYHnhCllav
N8XRTWVRcpvQ6S7UJgn+BDR2vAK+oBosYREOBkLG+YazWl6v5RHTwUVgoVi2mQL5
XPnC6+GDftL7TDgGKl/WFYYXZHZ0DQtowf5ZzE6WtplKpSyrdFalPgPwUcV9wfkz
5eTPkwICp/7IWA9iqCYqLRew7D5IQ+BQVYFxRQN1Iw0Z301QpRfJwKBFLeprud7M
hZGBnvESV/5jVKvUREzv5+Ykj02hHMzL3xB9taxbyGDQqtUUo0Gduw9OiPY7QP9g
00Rg3xy1b/zsUX/Hn1GqILHr9ObOdePa9TNbposMWPzRomLQD6t/BVe9KEUgLDR9
v+1aubItYHB3pZa0jdcso54CW8lE7SIXqSZG6wQ+Cf5N1K6C1PjqY1MwEasGb74j
PIkYjGKt5/wBS66a8G3Lf/WLeI7nOj3vQTVmv1KTZ0ujOiOU5Klb3CQS329uC2Y8
OxdOYPhapIlZFEeDGDT8aYRXCf+EtS+GUIi7zWvfnejOknIiEvLv9ELtE7Z3ALR9
or3P3thvaVsfrNNy+c1V5kUIsFD+nRoWTmA16Ovnisk8g3NpzhGrac4XcpRHnkAD
u8imHeOWBYUd+SfMVxoSrGzetrwQOf8VV7DOtSdn8IpZtI1i5vRRLidFEuywzsUO
WVOpbY4np8Hi+lrcjkGpODKCAsd4M6UgVbSmKefq8D6ei8e63TU16tQznNLTvMVZ
PwfpmS4cCG2mrq7wWfFfVcaCX5SDC2RITOHaigWaJF5D9qYpKr9ULe95usid7din
JtzKasSBqj/cY7sB8hlRBNdN3uzK7HrVU4Tff9Bj5IJwlmBUyjYmy9meDTi3Aevt
epA33Qm4gROcB3EqG04rWlB9zI6zHJZhkc4CXNsA/HBqnzuWcVH/V74c2xyLsDkE
ws+V/jNZjKor+q89brEc4tUD5bJk30NsZl9ZxJDwFzgVFA+ENT058T+TgKzSB6kj
Es4JlELwLLNo+SjPGdmSio13+0qvoBnbv0HFu2VflK3RGdDDc3X4uKl0dn48NKce
ca8+fZy11JbUAQd6PjNU2SjWY4StyTNUezbohsCGpTXZY64GFZkG9wYz+lxsuJ8e
WbBkxcKuMhRP2LZAkobgMTdMM7rRXfIrmNSj2t8PNXpSOJfF9dFL6/RgotRPIuj7
s5v7aW0bMOQzKv3UtjAB6VIuBgPxAKqbRtntqXhRge6BroWTCoiOlsEdOCVEI1DY
j41Xn3PzF6XR30Ik62UPudDJfepEHjo4b+Sq7BUbZrNyYUzbULznUwiIeoQ5kOHe
VGmdc2jFKKUzgZKpgfPu6EWx8ZZNf1m4wsccXA5a9hE8qnHZvXPjQ8zj8N8BIyL3
18z+QUTA72VtZPbMg6Yrz5/9nrywmTTg/XSZNnZHlTHlXPKjkM1xavfsuLJV6JPd
75bN8oEtxapCsUSpibYJM8XeB8xipJazdkorkNGqWGZFd9FcA9qGSSjYmHOpUvnI
7WtoW4zhebXsSe1kCL5qHokl8PYUUvaeS4jVmB5yzgqCiOnc6nnCLG3PtePJVNGl
UHXmXm00CvtQTW57yemoqb93nvkrBh8P77pTzn1R9rAnpz2ovqyviSqWRhPAQkBq
cRw5li0z+TdsrOEsvG1AnCKGH0RUG6kGkG5lC1YwHxOiic3vNYdXTC0XLHRkFqQT
T14vJbYYG0iwhTBNqoP3jMlWOqG7HmTpinkMLWdoNMdxzca0oSUL2PYGnTzU9rSQ
6jVWLmNSOkNxnQD6ZqW4DMaRjBoqOm3DZrVn0Qd+EMG+h9Ccfrs5ZoHZiOtvLi5g
Oncd+ukGVfTcX5dd5ur/a0GQk+l9IkvYLkaWnbW2LenYysFS/3dPPHkGJAIYHlj7
Huy1VVeES7AtvSqScmgOtLibs8KZxE/O4SK4RzLxxYzbGDp7G/OujPu1ciG0nkeI
pUmroXtwnYqJMHyYhKhfQCZvXEwUzQAdIniYwZRYNbYp+/S2Pc4cQSiaREKbB+Td
rJ1vGFEWuq8kFT8uxhCySSLS4aB8FA7L0JDnMCl2DqmmgviPWXvhhbbEa+m+XGlg
kBH4c1rjjsKf/fDQdWjwltPakWfOeywLWAEXI7mn8cBArMGlC+rImEPVVO8yDSmG
hLIzgVHP7DrthQGdoRu6onzcKhPDbV8y37LA2jkhAYq2kOwYSwoyDNbkyBf9EtxA
LCg0L7fDGCyAvBOdK+q7g9SrIrTVk7iIfwUYL8/ujbHRqJcfxddQ8u/cnesl/bpg
3y88MdlgU4HDXmDJI2CV2MnnKyFl12MIDKL4F3WZ3wUkRPnDye4zE+/PjS2TGLfl
93NjBGJFQtnHPFUM1CjYx8gvryeimKw+645NqazbCewQiEDzrPZH/tTTt5JJsSVH
/pH+2RtC9n9AExcDunApkunOuVaVycTVOxwJ5sOV763oT4s2xHSep8PYuPT3qxzP
0rY0IHYOUq2RrqEGja5joCmaf9ORfqZNkLlKOiEdoY/ASkm5N2XJteVVzdDfs8jt
BzbzS217qDBmpQH2OIWjerpzj6uAMh8ekELjzGmvAy3Ax3RvcLfh/zwA5F6vz7GP
/1l7QQ+HS6zqP5j+X9Ibpt6Iy7mj7ROdaX73C4Pq1V3TNJugRk5fPmgouc9Q0sMC
uwt7ur++ddjfrTBmChuexfhE0eKZWFKC5VCcxf0rP8NLSSb+vTFPUnyYoie/81Xd
NKw3XDYr6vfkGmlpS/JBR/gNFVT+ViyEkIsrn0t03CLbEnWPzbxtalbQYU8Yt1n3
mMqT4Ux4iMUDbcbQ/Ky1AhCEwyqfCM8rZK3tciyOIwU64BkXaFG9qKMHAfHgxeCt
rxiibn/yICktI5m0cir/zClPreyXU/+ZJGdiVOYeUEmR6lddK8ncmwvrPG6/ndXJ
jswIwVuvpoZkRbnObTQamOqJYiVkf7UqJfkiDcq4H70QJ1I1QAg4q8TNkQWr6qjV
hPcEEE64itN18W2qCMnODN+tHZ+ab9DT6nvmDkyvt1/6Ecz753raj6NHI/tPtMe7
Zyp7i1LGPnClL940g0Zpz7K86Xexv3+aK2XGOLQhbg0pAtoDp5e/5hHzIuLPl1D1
+pgmfcjvyCnjXJeLKyuomrJIwHyqZ0dLVLaqkt6Ukx13b5EGEdidctz5ZmT8b9hz
Akb/Pmdb3HPRl+Dd14YzJTHaQH31+r+EBOMr/iOhzram0PfAFEJCyH0qV5Ean1Gj
RPk5lr195Hfmh2L/XOLpEQGu0phQE/tVSfmLBhkNd+lCFdhvAEC43EsrV3bqVlVj
iaj8PLXiHj+pene7krR3+LqfLpFAxF9RKQB5kTUoICEZ5eb0Bf845WwudfE+8qub
OwQpu2nGCTqvjYKHbUSN6an/nIUt8wA3z0d7JQrupzy8pPRiobX0s0ZJgpP9Gps5
vPATXefrh3qVoMOXU7/6YRv4vQAIoxMCwj4CBncKHuxPXK22Ev7qc8YbhAsd3GxN
MG+tMuw9JvH5CARv195WWpzqv1SpH0i1Gzdn5q7cDmvrhyyDUbar5rr2YNZTsZKK
HuhZ5MQnemvguK0Ej2yD2LQ5SLGYQgJcWIYIhJo7PmvcKZdBRGNmVMktLkavbihj
KgvHkE/QDxcncZvVhwJJ5WdEU93/2EzskyNJpg/5uRPjGG7UscXX1ukjDNjJ9ZuY
krT1LYVo79+9O3m3d+NjtHa5TL1SjxFsXYuGb+b2rBNiXRMw1xe16ioSEu8qHObc
IB6e7X0n2AQdk4ccOfccFFrq59+4a5SCVhmdgCdq3VViq6P+m4AFAGNf3RDhKmxH
8ht6TFtnxMk3ovjHaqyK7Uon+c/PZpdX6AoefEKbc93ehTPkaJTGVznUUUoU+hcb
T1EAkdgiok189RRLe1soCuY/Vx7eJ5l4OALSeluZYcYBO1X4dBEiPOQBQO3AzNGS
q3n8HoR+i+btMtV78t7LhyKedg2a/Xysu6MkopSAPaiGHn8wOu39xbFCFUvu3HfE
o1jUosJrURvyJh3+ZsjjkaaUNh0fHH5VfxolVjQlFAUmc2568p5jui3VoKlCJTu3
7cOaBBMCX0RSx5CjmL5jWB6oDVCSzSTMfywUW2xHES/G7hVbSJ22nBgdYDAmMFJ7
jvI21A1Nitw/Jw6ShQBk0ujMMrcTl/kPOFqdihMrQh2z1NQmuK49/9f1zRdpez1f
VhQHgoQo2fw8PaqugXsawCACVoGzJVlrzznycG92Ma/aogxfwvPs5YZV2KP5Uq+Z
RHJ2ZDtuTcb8e5LVEqGaAnS/+cnZxuJEeu3XJPbYz9g3SjBYrEHc9l3HK+5sjX60
sJtJXcDLsciCiJPIMGKSDDzlSoQqvBIVj0u1avd4Dosgej/JDQk8RWjG1cSoNl5m
kazr4A2+NTkJcYc+73xe4UgIcvYWMOIG7aZPa32kMGTk1CyrbjeDRJlokNGNwESG
l9oGfCK0QUgryrOpaxDiP1q4GK603lfjsIiXeKtUDgf3C236hOM2/5NHbVOfNXnQ
yy8qo6djHanAycQes7xvRvyhy+ZqTrNtoMCjfZOR3P132gw8ONhdk1gctNPd3Im8
F3xf1JMiiPVFeJql9MoNJ1GLw27U0k3DM0GApU1BqNNHiumiQxHjhIjIDj+7wZBp
Zsz+yS70j5w5GNWSOEcEo6P+7vrMDyR9DZzJT9zdvKs30tOfcldZV5RSZqwnCww/
0KJwgLDtJknS08WTZIVvPWeKe39WEmqe+UKkdyEh34h3IDjcpqgpu+IvXYixjaYw
P/pjdhQ2hHgYnnWBo2ZXDTbbXAljY3x+/VfpggdR+7nfqoXCEOIG0Qmme+JwqnuD
RHi/2E+3DM16EJhqXpGZURA4yOcDlmZiFPpSH/s5cFyLm+EFZTqb2Nno4g/MnZlq
7KnmT2p6yb8BPMQdE1IivakRfcUBDw60zMCm67FFzenpldprbn3qMFsZ+hQfTlth
vBzzIFGd1O+i+yggDQwiZSkV6ZnKNqMGrzGXZm8ZGzqK9InuxfA9/lbFrPv4f4M7
WLOKLeumGfYU4yEp1JR2jPXAhLYy+xcfYFJCevqUMirjf7W5c0yTnVeKdRZoFzLK
MNzVYjmYieF3OkXUU6g+y0jXxpNBpouIGelxQPj3LFepCNmb4Q0tmxPMVXpXpyWK
fgLAsKG9XG2uw5P14nLJ1CeA/8Fqx1ENR9zXK72CuAStJzarcJulc9yYI7r89UWo
wooHB1ZkxYuqV9MJ0cnV27b4DpRNaMs80dItHuCjRhU757+F9ak3j3tt1AAA++e4
+bnRXM2wpEMAk7ojfIR3srOLTiKNXkSUn7nHNli+faPh8AhOGE3uShS7Uyc9yTDo
7xlQ3DoBDRXdz0VEDyGsEtJlTMDYARhz+uG191lO+YhvkYHj285xpEsoh/B6PmDo
tCa7mGQJ/BpJ+HBlz2eV5kJRofoMLMtfLw4jK9n95fzGvvbMiM+KVUplWEGQhJZb
bYbf3DxampZAM/PYMyhIZnfEgCeqXmUcs+AS48ymdwA3ThwVUg3w3RhKLuIgzoPL
g4Jwy2LkkgRLDKyw4gKOCoxPtQFzN2NId3iEg8yW52TZ+r2Mq41Jx41yWoxlIytR
/ZU51DEzwxRLCUfB9gC0ogzRzpBZkwAxsP4fB65dT/yFsyLsFflmxYLnpKp2ySq9
j8VCNR9K9Fqgcih6RxkBf73JIRp44iPap1YRF3qY2wG5/CbISPhFbEcy+F34kY3/
Mz2jE5CgnE8bxSYZmu5f/zG8AvxEasLUKP/bBti5yCnGMi1nTL8LlmKfvL5/KUKu
PEylFJgsGsqBf7tK590DutHZg6eWfAlFO3SoLZwKgcM+9xD1+nMvYuMNFRvkdcW0
UWhCESNGh43ehgUU1aUkLytT+jOWcdKKM/TAPabga+BCUMAPNmkjMqry1uG7ta0U
vIoRqVClNfpzTHP4DCjum0aHx1o6oMOYjhPmqziQ1ey4HXMbEWEizd7flMMLdgwk
Do2nkwzEP6kjNxtR7pCyWQJlQP81UT8R5bq+D4NUw6+0hR2RTchS4kti+AJpsKjU
/d12h5kMTO5hf9wmeERkDtclkURVyUEvZpK1EL+MH6Wt67mEtH3AOad6fWUgF03E
OWIZ9OFYm6AuNfw4TasMfhkZa9gn4SnlR53ZK+2cLh0jsClfa/Q/FhVR+XX1FO3P
JwWa6lHkbW7urfHkYHIDCVJB5/tDC1dn0pU5hIsR6e5d6X+HVRRmpuQI6jIQjkwP
h6LVjbCVGMYajcGMrKvEUVRcxlx89aBH9PP5eaWu0wESp9UJLUf/aCnVHailw7Uk
jZwF3cbmhexWaTmA0jLmxml7XAC3n0zfZTAShjzGyg3jA9IK8Wx7GGUOhUi8H3yn
Xkv58UgiEsUYu3VvSBemeX2SB4Ylg3Le34tamfsRUw84NLfHrpTlNkFH/kjBcdFY
F3H7Mrk4gs2OUG2Gl99IfH5SK4eHkV60Z1cnD0WKU9KDFNwBfPNyXUDNsZkwunxE
7zXDBy7SGgrZ3ZsbL2gREX9dX+Uw13fmbwP1XhmjdknNHsBKu82eFjKFh3YQswwt
KAxGu4MXXYwc9c9GmdRlVX0Vf+t0hxkQ6yx8gh9sQrljjKqJ7Os/ChMNuwNfRbvM
zaZo1iySteg6DB6jNmdtB7VHkPWfNc2i4y0Kgy+Gh+Yyx+kEj0v2bI3XuPV3CgJ0
f4HLAfxZArE0RTE6O6vztF2SmEUKO1r6tZuzl0Vb5zbH40krYktFXbK24Rm9flR7
cDQf8ehiYgGfYbPAZi0/UeCld3OJ0xBR3gECSRBrIKpxX9BjL2qLwrmCxZbb34+F
rns3+zoLbFh2sJslcLIdfGml9zRhn1x/41DNvU1WaRfXTbEyJ8VEGv5CHPFhfBLG
1E5K2jR1OKPtH6ysK2nVSil7BJKvCHCOOdIzPXnSQ3iKTlpHeCDolJWd5F5LhjX1
iZISbRYI+C8+aa8ma1R2mt3WTQKp46TS4EWIN4SCc4QbHjO58TyzjeYhx1DFmeoB
PNKZjYrmiH58MdAEulQ3dHusix9Py0tixBOsuBJoNYoVru479/PSwu7JaHM6BWvF
hPtuIYKFVW2Ul4FOrcXsYRLT2KBod/Y9lCzUs/GppP0dNKvo6X2YKsTktRxdRdQn
CX1IA3dM6iMxB5zk8asgE5dzDAVCg+nl+dljXDZ0bsNBEjx17JczGvoYTjGy3aO+
JIl9PJ4uRZisUi1VIYxw4fimxJoVPd+WB4zHT2U58/nqyRehNu8R31bI22qp7kBW
9X3YpyWClUO+j/FslQaPR4Sx6aRYsm6JhbghQc5KsRemIQtDsS1/9xZASkXko1l0
K28ZHAVKE4JDfz9k3Jm8FaQbGtVbjj8aqIy4iYyVtwFRWS9OvYeMbfnrtufZxXsO
j9KaMLihalorP6yyCg6oRxkUsqhG7HPLHwUJx+XZWX6CKJt+Jf0zHpehukmjMdbB
5m9LPYW7jsUpyXEPPP3IRRFiqQsQ7D6vpYHWh68yeAzOmZdJe0jWDE6z9AT11WrV
zKYe0/BHs0O2lBvjr5SQu/M9+KazNQopsB3TyDa7++wnzx9WkK+Q0Pkd2OG0Fcjp
6FtUS2qpmzjb+y1iVf30gXHtjbLJCp8gMDaA86FQ8Kv2/8LBHN7TJ0G2tgpa1ziE
kIO0g7l9LuI2juu+7t4R5HSAi6wyzsJiKs51grtYun03S1QQmcEd0Snhdgfx9S+4
O7Zgmis65Pyppuou6NG46YpyqD5RhLqUEv9stm8+HsNwV15QIa4HzJSDyPreMWHK
J0oQ0htjJLtsBShD1Llq4todFEHdxcNkMa69P6MwdSXmnCmPA8IiRn62gBeDtS/P
OmsGlpZaL6FvFwqYRkNuGcHAV8J7oT07CeqeNZ9d1dZYeKvsEVa8eoOjPrOkJ9+y
kYBcDSTeKuEWOvU+8HTEhlALonFQPh7lVyYeIbTNttphxZjjv6S+Y4Hf4Jw5Thqb
CzUeKva/kVLhHAcxYdVFiQQOyhqwJ74hnUeMvXEa8nrsjeqyondQB32RCelaGSCy
RfG85i1k4rxhoCYdpsjqL/HDKgl/JL6zMDGpszW4p3LrtX9gBfXBUzskKgHFVokl
ux5HjeNdyGTJKtKXYFnp85gJwoW4y0yxpbIa8jaehV2c30b9UScNn0DibUvN6w2R
iWrzYTA7gQnL6qXCYM8V1IfNKipPqfCYynxtgfgnG5faVx002n5DeMNZx2JHLMGK
0dth2KiGR+PocxhRDJcxI9kGPFJP/lF6kxfvgJ9JY+GgZ6sNhe4diBMzzRoFsnJu
n09gSXs1kydDmt99RWmj9T0hKuVPBFK98mf5W+irA9Wr5PqebO6/eSy5fFcyYQzj
SMzLc5NYDp2oRPFRjcIRk/9yK/entCk7zUFs/M3TQCACSY99Mb6Mh6k7RkSlPYjv
eyySVZxWdw+19WzhPU0tRu3Yb2tPFdIulfnxfKkRlnTxwFNxOL6rG/Ds4Q48HBWv
DUN31VyNxAi5k7c2Qp6KyPSYfJ34V3AGcpZlYETJ5zgdYz6fK1yNcHUtEl7lCtWT
BFEl+NglGN65UFAGkhgAeFbeusXgpels4d2Sbaprew8kiJGIwHmV0bl8LoIPvHCE
rgQ7KIIVZ5vboTxFoGmqX/BMBhyB0ZmOpSTmAZSkzyVAMyp3bRFDcU3MGLUA/Rel
27M0GQS1gCCK6gPZsAAfWWIsB5NjVVq1GdsscJrsipN1kzd7Xr8CAtc+UeeFF4vF
M0NY8ll3Uv+cMo6aI2gYfqBf+EoeN/+inFU6oX1HKHiRGAtt7hXKKlgsBu9vkPkT
2LoAoNv/O7eWPTgX9Mg6nez//RuCFfnSFwxsbzwNh3NUHgNPWUt22t1L8wwrsQ9k
mezLRJrpLBHDecUU3SaVsW73JoITPPUBKYdeZ4UEAOqLp0GujvEhiZ1kQ8pspUeu
wu62A74mCZFaE+6U2RV+7NfzCSOBVWpzBz3pOb3UuM6TiP33aInUUDoX/c2hOxq1
W0VF48eifNY07l++1UGJm7+fGEM+V20iEeske3HghF7/t/+qB61/sVEQLZL2cCf9
WoCf3HYRT7p+Q25Nz5tVFHvblSrNAB+2PQFNnXO+M+08+fprUfJc7bLttZsUjRBL
mCBwQs+4eHYbU+FkSDWEWbcoHs2jf+Oz8ted7JPdEXas9IoJ3R0nt7ZP+bmrflOy
MZlImZzPxSIuKIglqX5PqyprrUdtere7byoWJF6Djx4ats5GW8gjRSSZBajIqN8j
hdqyaCEk45Gq0UgwNMekwxYBzsuFTpgzgdxN8FdYoQM4J/TBJrrfrLJiv7Tzcxgu
mGFng1Gcl6XO8rbKMf3vU03g3+l1vY0ULqk5rwAeC+3KwzrvwPUQHQ71ZiNsnIyc
mP7gLQwa9D6m9/rzZj6SAA==
`pragma protect end_protected
