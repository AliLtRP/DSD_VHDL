library verilog;
use verilog.vl_types.all;
entity not_gate_vlg_sample_tst is
    port(
        x               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end not_gate_vlg_sample_tst;
