// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
maWO/0Bq5RxGRDeehBaSkXybmDmTjeYvvkcIF+OpuAANvpybXOD7Tf9DGJhEDeXpWKta+WFTVC8G
mu7FPyqO42sXM5J/qqG8V7vu1LpuvrcSkkCDAAg11mvJ6nlBG/Nj6jfMQ18Ruu4TAbuOAyFILtI6
SgFr8I/xGZUqeA0L4NBY7pH38I2SD4UYX6jjoAD0LUdEtSGpB3gy2LTC+aAzqVudgP6FfW/thnND
Irz2A7Qv1GHj1MfmLNM+w9qu/ILcrb5JEsToqTPlAIX2Ajgu8Ef+KRFiv4y+k8yMTN220hjiZji5
z/+sOT8rim8JnuILDnXhTdyubaEFlSshM5r+5w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
+9H5M32cAdCNFVkRlGxAm4kDcrWgAzI30qYOwGilYFYkFzPSFlTBUlKundDcylUjCRS7MK9KCasx
4J+O0ozIDtuKVDLVBEvHfecrBOFdVOYQTRLjzFZcclOPdELIJjI7OzYNq9aNQ7sC0a9iusCyff9J
QIhMTIfTFInQdUCGgJqW+qwMFQPjSrTUz7lQar/Fs58yqDsvt/VEOFt9tf/48vxg2gsZwBSGvRNE
cUu+cCQaG75tA3S/ejkZ0iIlZtQYdxsNBcSEiIowuHjDmM3GsxsVJ3XXiSh+zMX/QmDr1IbCkio/
fwaMUQ0hfJ359Ng630Wab9Ljo5ijv4ufQmWyrEH13jTOkGT8HxcmotnUWjfo10HxUZ1W/dFW3U6x
UowvEZAzxKly5LEdiQZl1GELQxisvywku54DBk0BKSl18C4GxjB/+YZhHS5LT3sQq7ZfYJo3aeXA
Yt2l53IpKr77eKgPjGdDts0caC1DYadqHMyZmAPNnUYA3nahX/c82RknaRmlxjVPAwnBy/Sb/YbL
3VWPxxEtCyoz/mKOpAz7WbmyEMr0KT/CtB3o0EXFzSdBChHuw8d5PqmitcBcecjdCsplwSAQ4HBn
r3zV+yyiZYGdeFxfnvV+MuCWkZcC/TgPa51doNpIqV3bq27wrTo7lnkN8+Jb2yuFT5JS6f44ZPt5
daP2lTd2oMQ1qY6vY3RHYdGURZfPoxlzbFfe4EwI8ocLA9i1UU9n/3DKLsGw7w3exJhpfaixER8H
FyTPgvTLY7xoZCf9QjNgh9IgUdSKtQpxIDt1X3xrJzEEFfm7/vCgWYMyJA9+KQDfaYsG6lFIdOan
K246IJX5qOn3m0osPQhnBra80lSt0rTl7vTFRdlVDdNvc3nDJ1n6aOOcaLk/9wnA7gY9gcb9nqws
vMlfwX6qPwgJS0uipFPoEBFoS0k1rG0rtrHRg5bMUiRUHG2oPDOH6xV4mcwZPZGUVcgVZV1jqQcg
nHenuES1ZHRUvtzJ2sW5rLOYBgzfoCZ8NLeUXKhrjwfxuvym13iD5q3ScPZs9Mdf7d0XqF7qfpXP
YKcuNO39zPcaGWVLymOiYdXNc1LJV7j0zGFj+/Ro4mfQZHZ9p+3aYdE9URA7KXxtA094clSiei9B
vNvfS7M5Hk7rEX6vjr6fSI+PJZAVOMEP+BEcpGGp6TF2PEEmFfFL4tvrJG1SeHjFD4zEpOOz5Xqq
NU+cjuPcmUXqeDO+My4YkcfcNpIGNKI94s4TsI12OW3eTyGw0QUF307Es1HZkmWovFaNwGWzrSVv
9VMo2qBIvtnYkP1OdyD240eVMm9CYa9J1V2mRt/EQgiehYrIbUs5ukUuTMo9cl/Xrna8gd5MvS1n
m6Kf5EX+xtzdrx3qNtsOXCtKetEymnxplSA3sV1D9jNozfYKvNa+6IeweyC3XdStWcWbB2zJFV6b
oDPzLFg1cQRkTi0KczgQWmics+C4i1fp5uOAv2cbBngRq/7Vx+MRGAsjPmJqfMFhQKtqGtM5jFoD
6ErFAreacBqbY+pKP5lbNsUjiqvFnjLBMVaojSrjAXUhrb4BGMp7MmKJTmqOforQhDtPJhIpQTFZ
STsZc959m/U5r2XJ0Km8AZZtX/mfetp58c8E5zL80oUElW/PlDXDzQaYLDXodUoqqvCYQ0luvAO4
TlnRGIvlC5nLDTJ8vJ72Dvl1QYtnzYjyfhOWeOnLUcB06XZFvNu6wijbEK1Do4jgl4xZ9W5vQLQu
9YGmfhQTWpKbpynesQwLA4JYKNI0EHzQPucTO6vJGSrzz07pEfultxpNqmxFp9NKjDJ279EcMBBC
Yq7QZACBBcdaNxwsg7K+YlIMrnF1XsNtjlUOA774BCrlUvQq/R4A3Xw7DrCwf59dOPPs6E/ZO5GW
zA5vh/qREHxCRtion4gxbbl6PKHBFpbdne23Ki6Ca1PUGwfla7//8twWOro2gzicwg1b3zo8n5cN
iblDB55xUM6dmmssqYZ+4EVZ5OwhLwZbU2MKgAVoXrACycmAV2lt73M1rjbWmCLQ5MPxVGlRFlVv
KV3ouOFl68k5ulKHMYLaHJEJXj3es1R3wVTdvN93KysT0525koynY0CYpp0N7bzQriAF3iGrstg+
n11lMYWMFSN0Y2bGcfyh9Xgst7HCZIuPn9jxmNVD9eQfxFg/w6VXzACI+vUXkd0lh2M6Sr1UGz+Y
uBN+PPwCByhW0thYRFdJEn4qUmg1ziAeLS5ccvEa7grw86k5I580NCkh6dX198Y5E4jhXnHRZSnw
SwbpoZTPhvn4LZr3GSWeBBt1kX/ybFUp/f9vc1AwLx94jOtjlW3xs4+M2gwRTm43g/+ViAcnv5EJ
xrp2G4cvId8xCqRIWcIdRhv6Ip9DuirhKubCJw14gOvxkVbMXfWnBzmiPQCjlFc1b9Uy51jq/9M7
rPM89+/EPqvvkLO3c6DeYA5z1jFWX9hMQ3sDQ9z6JTRK/bNvWNXGG8lwLCq222AUnwqYn+6zw8k+
eMevEToW2c9G5DwF/FIoZgLAMjhMnwss9fl4tZgS4tFtnwYwnG5RJUm2dit3WDvfIkVBoE6HzW9r
dGan0wN3UTuHFkTKv6CgEutHFV2roiKqZN36xX+MaCIkJFxlapuKT12Dkf8q9Uy0s/oiRdA4pLOw
3EHRkj4nNNS6X5h8eOS6EVEMWxNSWRRJNo+LrnEufqJwK64Exx8pW2gd6DWY6M6Q1o1J1x3oQjlz
iNJ04SSZt0aDjAicaMRYf0dyJRhDZPDEPb8PNX5iy+ms3jxikcoM5XmxucDqCi7dmeoXthT3x05n
W8jqgl77l8sl1PROHwMVQPK6M0MpLX+fmAqkp9QHldQ9ihy8NdaXGuxrhNSTXCAHUTufsgEsUbhU
j4QWqwKz+XtmWgm0sIQYsqo+INL44GdCciOE2aOibbsaq/K15cxcoWS2AiArU2bWe2XtvG/hKPBX
Sk1Q6BkPp41dTQzExxQRO71CpTgP5i8aZo06kjynDKlvAkiIKF5bu1C1BrOhbYXKzUNYO8uxAA0F
1qR4k1BstObMD90JcSVWerqhHm90ITxakeYdbowu6TUVccGIgyK48bOap8DjE72ohaz9RLIbc9i2
5VkWdSoRpqtNGppHoYA483tJgFcjg8kqVzUmFKjEDyXrOJMDmm65hFc+nN66yqs7H2lm90vgNK4O
6wSr5PomxXLtr+3CCEysDrhX8dlN63vDrbswuL87379HnBPZU81OFyBXNiruNTPo6Bfu83zpthU8
7WbEskALV+/RsA5tu+c4+6XEPAXNCqWPCFZpeu5IHPuvcuDqKrNnJ5XR8q+rmREhy77dvrRC1gm/
3h6K4t1zZdvUc28fKocODs8Kw7icQ3qIE1WMpmL2uMFmv+9h7ANbFEDzrR06DUqwIAdapVEqw5co
2TpRDyBlF8Xl6JdQzDP6ls/ctQk2oJkAW4Ec+G10tN8jc8lOshIFQQXpO3+keEBVRGg75wrojJ/G
0bpdbCIcZcY+YZHPwgHOjz8hSTsU3YUocKJ+vUer9qlm9ETJnLI1rQHDEyKkuQGXYKgSlMYePNji
xEDKlTTyyoQr+sJL1rn6q7jxXmXs/3PcTLI3YwwZYMZkuZkqL9XkBSPxvFVjebNNuuEh+bxTBQ0l
49tOoXDuQ5m994Grhu0H8aC/qMjVmo43z/KiUcMwXVhylYTEZrq3Z+ou3D09Su1sNoynRZhCy5Ne
DCnthzuBg1ZQWM2gKQVEvItqPv5HCHh1c+WfJmWhngI4YV8eeL4eUJmd4Y5cCpYCq/5Hu9Qg4boq
pw5My70Sk/qK6zF5Cb1Y1rS+rH8LolO4KFUbRpxi0cbUd207Eyx+fs/vimVsHSUE0es1i3H6fIdW
bqmW+eQ61/xBGUfR9Lf3Pwksg5PNzvlUvaBsAAz+WkzcUU7dxZH6Fz2EmWJBEi1YYGuvfaV/XYXE
lDOmAvhlW02k4wQ1Z/R260khIo8zOR04jsof5H07ywsAIMiHxQA3sikc0AqaGoEjJNLoIeRtsWAI
tEyPDdC6uI1fTl6ctGFjgN621SHe25n6JwTvV9km/9eaWjBlVBBBTUviDRfyT+MBK4ACtVe0pimO
U3QFHHyxkasc85YlDsS7j8OgYQ2WQp41LVmKJZIWlDvvN0SbrYIlSs+rkbMTvc4olX1mbln5iY9K
K7pt2SD85Twhaz+asQMp4YrWECJTz3qaOJfocChx8T3xCWNZMeUFiZ2M95lYkfZQZNqZUAN32Yrj
ojaTrlsIkEdSHqU7rZDET/TjjCeuf7bZ8nkqQTQNX94SjzaHyTeFbwK7vHTS/I4X2yXZwNoeV9xL
XaRUoXX4eIEAekF9C/T56d7Qy7rDVzJ3KiO8Zvy48gR0RvhLKHGJzMQcodyCAAfO7ip6xz9un5al
kuzDhm6aeoPAvgKAqwVNCbwgWu4bcW65NJmqIveIkdY76NFZABOo5z+H9vk8CeexVvVohpf6kwP+
/C+JxenBNNCkB9PsZN+7LEYDbFG5U0t1OPn3zbJqJ1iq3mSD29oMLPi69izb7ETNCoukI0xyewR0
/jAhdSHgE2slq9bbTJab6LTaU0sbnb+01xUsvsYyR1zqJFPWuHkoLDO8ZYDkDgvfap7DSJxJ2Ir4
+lgiNn5f3DCj7kyrNaZz9cHZr0KcWNwYzpWqf5ig9cxw2F/TmNhhRIa12R/+V+kiC1ssX4gWHxEG
giKa3H3+bA0+SuzbGQipr+6VaX+46Rdfxzh9XEskws96DBC42gkkmjJ5ObtZbu5f1x6j+mo32ICm
kXGmwSvqt8otJV0HxlJQose3KJXeC9Rm7ayHQSWMewUD0qXR4KFWdUzZbFXb4Q68N27uiEgz1+TS
zcGQGytIH8Qkugdb2bRKG9Ua0kr0hUbkB7knJsDt8qU3UpalbU6TkKA7wLcF+uOSQGCRVashRBei
7SWSehikgiCp73dyPngH+2MpLKt//bHQyRXpfrRrgnEkgGqKyUhOaXaRfDh2dVBGomMxrqc4dwyU
oQ4J2E4rDVW566NznHG7jCSVT1d+2ReLXkEKHQg/7Kuie4iLYV2QipwegNDm8CB6BmPCGMJAlkqN
/b/VpR3SS9kd0K2O5/Ue59yUoYMKEODzrBJAf8kgYjo81XlUBfJmTrXWDr+3uGG6R2OqtbyW5x6Q
OoJCSlCvlf2pKlwCARHQ7SYnGZ39dA9/8WCggvsnR1PtIRKAEM9mBvUEf2GgjaHCeb49TFH55gWO
gZmeZhlBsiUiRWcQ04bAYR40pSam/pt9Wwh2k58VUTz7Iqt5ls33IHw+3mmJtn/PkZtoj6Mq+zpo
gFBeTsqHyxKmjUmOziXx46bHfmg1X86qzOZQQVoiQ9DKBH1Qe70fvlgs1pvenW9fi6JYPBNAZ9FY
USnV9NQIyZYM1xF7N+fJe+2JmkN1V95h4xJ6rY7pel6udDd8W77DbBU06AowaXyPHMdjiu0m54GF
kGbkcaXSgVbayjinGPtP6vxf6K4eyZZ+cpqYPUp2QZW85cNln8rfiJA0uvY7qIn/qIL7xGgeczuJ
U/mu7NvJA13KM6Gmz4Zoj8a0gir+Yp6ofT2IoqKn5hv14URpj9nqNfeDBEu3KJ9wlYkkuIfFxhXT
zaSRv0e9VZIIZB4pvcOKUBobw1k6CaHP0IXC1aZ2pFM2O3VuLxp71xKQasIibkN9mdQRMF3HRUIX
AhqIeRrwpAMCGiwhQX19PmCLieyJ8T15C3JPJ3EwHgWhJ8f+IEvCokp0cxYVP8oiKlR4shuTbhfs
QeLGU1Ju/n3oSR6tJeJtb5sZDEPSx8dD1NamoaqISWwl/RanSzq5OgBCg+agQtkJN9L1srA7IJ03
aIooV4IpPYboCvTEqD8V6pFwZRgbYy03bqF55wXXNpAytpHjhvdAJsu4CXhbWdKiaDDnyv/aRMuh
8/ITLUAtqKJ0gOM71Np6ll19unw0wmTajW9JAMnPZbG6jdAoYUBBVcBpTtQnWT7SNvtVla4xK3te
OE2ScJF443Ur9PKjxyLXKQqNT2vUDRtBeaPDtj4Nde7o/Ie/I9ISkR4UIXRKwi2QBRvNtyWbAsqX
AFwGWBjufAD+iFWT95jcaXQ5jX45xW4iCWPukW2QdssGErOeDNp9y5iYt/Yjy7L749g/YKMzsCn8
/b4iHKnAQqS/RBTVp9ZSecmGLpNND5RidwWLe2sh0knSHkVoczqIM5v1MvUHY8rCZnfKiSceCHE7
pcbcA6KnDH1RRtsEaSm/1GKZ1X8uB7JfzbG374UaBAoRgzZBYMW1LDmHJ6/uLog/cN3nRsm+X6b8
L6+OFgUP3YZ+wiNIZIHP0hxSvqv2X0AgcwA6fW3NImZWbnttGlQAsxCmSRNP92sXCRBSQ+APfj5x
8t1CZml6GYKVlNQowPF82ypVOgox2VTC02FM5VCLVS9nTBwfES+jRmeOsIHHKodt4mo2cWreJB75
WzkclRgn5gIwIbMmSHjswJ+xLb7o5NCqdcRXxhrxuNLztgvBKDwRQNi9YBLfMjmVRJ7n9CXVHP1z
qJ0yO646wUZBTKEsLGFT34v9Ni2/B1kmuOLlNdUNzxWnOFh3XLqFRemcPYhUIFdDNWuD+MEP8Nrr
FZB7x+wGuGTfwUfsvD+Uz8ssS8QVqKjK8/pGziWSKHIr+DuAtWsl0mgASTlFmrpzwdAvZroRMxuS
Ubc1nVTcIxHFQomHxV/+g3WruC+YRXOlL2RYgylWW/VlYntkxNuiwoFE6Jb3L888Qm6S1qqnWPH4
T0UtQBM0s3p0pJXZ7DDI3bMof/PzEoUYTijA5ajPiSqZKy9krX7pTc972E+sqTabXmoCCRYHtvcM
jiqhkTFgMxBrSVrd771rWM34JA5jgs8KcRS/o0VUEcqR4LTqAtoM+JB4ZzX/d3OrYUrSECps1zZd
K7PBjnlOhlzgDSH0pmtP7towSqLRFtk54a4CiLj7fvwobydeLQJNh1tpbmh+AWvRiiafMR6+PaxQ
rKDYVp0btmZ2e9Vxd21mDU7xEdEoKVIpnNL8Pg6LGq72cvIDIbN86aWHLqrIMqXLifHq6w3LdkMv
cgVw9eRHVQIxED1DKmSxP7JsR2RJwTEwKOqHE8uNWKWh1N9HLgDLdzVrheDhcahG9mMpi4tQUbaI
Ht08R5KIKWz8oFLuTCcOigzEIfIqgPOK5Hi9VcT/BHZsjG2FO/STGlcjHC2MvoNuaC+y/VekSkHo
9gswZNWm5/aZHtG/piYP2x6n3UdxtBWbFmOLx43TnWIAIzS1KjDLa+k1j/9QBrSWuSuyMF7w9/2/
QJqjILENR9ga/+vQcFNVLDxTJQOHalzqgJc0uYFJR46QXA3+l1j7kc05VcU3Gbc2qLKI9q0nzzlq
/X1YNMdAxtYIdX7qBUhIMY73Fc36uel0eklNgiz3M/YwVijTq96Tl2R2MmSZZ9ouitBtKPGEfea/
wT8wIaCKdtLes4ZsXj7LPrxKQZ3V5+DBl+J5FRW7cIzRh1hxn6XA84pfqkMUuTUFw1YJeP6Y9/Yu
BbReNQ1qe6p0vSMJtkm409ziYw83rSOBxN6FJKK6cv+NKwWx+TPE87HohHjTTnwjf/rq/7Wndtvv
0ujT5I1EenP7x4NbTFUA4HmP2T6x9bqfN1339VVb8p6jvIWwb7Hk9NhdAghrW/e6QiKhg66tEnC8
Lq4FY56VaCNsNraXCB7e8CalhozQLyW8jQNm781jOiiGLrcndKJWy95WdcfRZPnaKcGCXlW8Pu7Y
xirPli9d9MEKWBpDBhSZYsRwx2ylmV3+d8UEWLM5p4AZtG9P+I+fKrCOHP/6jsxdhFenLzpvBizr
66QWVQ3KOlngJxCBqe9nKGbP9kvc191fptePjTE5bnz90/pzfTsnySj8+XtC8XxvnY0SHKC/bLFx
Vcnck7TRLhUTNmHwxkicE2r8fkSVZAELwKTaKWFUrSx0JtbA98RmbQ/DC1yVu+xtdGT0XTIzWp8x
LSUM9hr7ynG95PyPZUbftNHF+aJ8UmCIa1ra34p5ZhCx6WO8WLAS4KYIbPMdQ0AQnZfeuf1Pavll
9E1LQONcxDuZWlPALKQAanXzzCnhSdC0KuB26yVoxgID7/sccUR+r2w7FoNw3gc9ziJiJ3iMXNvb
eq56YEr2fl+FKLcUT2mChAUDJLrmexKZmrbzTIKsFvmLqHxTq81w4yDEFuxqGJdeyCsTFnSmiOcV
pdwOTNs7WlzI4+Z8fBRZ2aM2pcHl+GgjlNZmEJiowtpb+i+bgvBkjNBxv4u56ZSpQr5EcdRXdi7/
/j42zUkk22vhN0XJH6EgnzM69wjM0t6EVgdj+tkVXOJ+vPo3SEbABYF2KKR3X2rzo2N+3cCZTU3+
N9ovSl4qjk5xCg2J7Magv+JTr6FNPklzvgGhoK66qN9GEpd6kvydiCxGnVwZDpzjSBN7GohoAWj8
pv5HoN4nwjMn9DtkZSv90etydlAUfQtT7PoBly0h3Vla+WyPTte3iwWIEKV3msxdPDT+imIGCp7v
deJLcg/NINUNBSzRX+oE81j9FgAJJEpSQ9Dlss0hKozZd/h5Mb/ujdosqqsyyu1Gw4tEemTOOkSH
yaPX7dYxSqMifZSwa5fx/XkAv2Lf2tDXf9q0g5hqz8aD1KIfctVOFLSi3D8893B+B3If2AcTBcV2
jtHQsOOveGUiPu0MxnROjtj/G/Xpdfq/cCQz1F6huTMI7TLwzCFQJp0ic8ML7K1KYIyVu8/qNLJD
AsZHUJ8D02D5b1zLQNh1bTzmxsQDQhn2nI0oFa9aHGhe597exQeOtMhkfl4NC8Wqjk1KE+MkFEN8
PqhhXjeXkk1gt8kQX9M1aa3bDY2BZgfus6e/NA2Us0J4e3nBe/Ht4RQo4Lg2FRpRulcO5g4aJbSP
4Kvg1OKh+ogQvHR5FQhMS5NPJ3FcT5kaNSfGv5RnvkiZZjv7xSZSrBXCaqI3hMfDNXwn5xeWGVKK
t/kcg59dPNNrbF+VKh9+ywB5X/Du29D2zmHVp5D9zKJpUNB5/eqnMgWV/FGtYyz3AiCMKklQAJKD
gVEE7xQmQxP90/xOMrcyWJBdVtAvO4FftZeBMpkemMayJU4UOFOyv30SkjNxJdH/hCI4E0NU3IiF
ku4vciX+J2IhTFteqCNlfN7OO8jwnjySHcc2zdczDBuxm/QyAHDP5bkAc4VwOELYIHo2TYodC8+o
lvfmkyHlLcDES+Ne0g0ZzQLTXwNtF8RD3e5ZnzJvgYDMSP9rbxbAJtp41OAagLb9tuxz8F3rJfOE
IAPMXoJcE/XK1/XvBA4Or2MyDWPdwG4uLtGYsIRY4p1bXIcwY4FunChDiQYD2gL2sXQFYlKxM3WO
LmClIaAt3ytaMEtMPnFCVp4GKCCN+ZJ1KDZL32DWixmcR2JO+zSCgYnjG7yFS2GmUudFedMMPCHh
l8awphflv09GR6dOkXczSNRnZK4hRO2iWUPwwYWc3aOmyxVMDGvf2IghO/wBZLlOJJZCqepU7MX0
dF9axNq+3noCyp5ALV26Zge63hkhGZMnQK7C8N866Nv3u5JW5X6xQ9uVhUCIM/hBWNaPL7g++pZL
//7QOQMUDp1xgs9KTFDPBs2XKAkbTi5cRoTqYhcskxpYl2u2g3XeZ+4uUwuTIRy7LRSRwVedsDs7
Bim1LeA0EL4uqJvUZz+TSV/RENBX5EJ7jCLGkG7HaJASCocSm6TXXsf5ST5psH6r6B4VvHbRTBtY
ScN4whvNnw+nDVXc8JZde84Qb3s/VxWtErYH0R3PdI/GbeBrLJuC3QEryW5ejhpL5x7ROeA692NM
KjXe3q+3m4AKknQGCbmGCNUI+igTBcqIffiWUE9cFtopkJAJg8wpereov9yYGBZ8Txt6digMveZY
NeT4CYx9gLU2vUAfsFjpJW3TBKVzb9oJD3/6PlGQ9vi/W0yh6vAG6IOYqovcvTPgoB7pzZm9O5Vw
SGv8xAKbaneuIJ9zF6YCwZ5kN01ZJQr8u3MKK3bkbML7BZ4sNomrNr89/9fVW4tc5IiNGMK9tkov
+oDT/gXfUP2PKJXB7WqHqamdaZMw40+4plI8XxUlFCq6Z9CAM2PHcTRMwPfnHX12iool0YciB9DT
wqvN70rc3Uc9q4kNkZAx1JMcQA2sZ58e1MCsqhEQ2onhxEJx5QldXSL/J/xNUIeByPxX7XJjWW7H
02x8SDeKliXOvAD7Ji+9FLtGecCP+7J50PDrKMkAjTqKMvJ4swbi0/UhuIj0f2iy1FWDazIrMJZb
jHZPS80x5qXp1vrzsVNL9jKFrZVFHxwwVg99OZO9ss5/q85YL/cWAtNZurX5caXCZPCQFCpAw20n
DMQshc3kF79GHAyhuqd+/dHbjb4LW5ERmtR8Zlohfur4L9FnqHE2eRgJDHT4Iyj7Snepev26jgE=
`pragma protect end_protected
