// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XeRIq3ymZycJlkGGsq4sMcXwWsQxKwP+4v/QlJiptS9sDq11ThvFlz4CDA9T+Zut
u1LB3LqTCCD+IuCQod4i5HXGBIfi6lVAMbZGYJgreicFcJiTBxsqMmWu9dV8JDAl
tcTtK0YtmUEUqWBpRJ6B9kHkUAVyH+1b3rATuvXgSbU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10352)
kCDICGgZ5lBG39Ivgi/PKXhKle/NOAf4CpoVeR2mE4TI5dDHYDO+xWl1JfqJfuvM
+DuQbZaMBZdV/xWS1Pjtet2tGGR+syC+7B2ws5AZCrpdE8dOrfPiWKTuoqgLCWOm
KEwYJ0WSENVzlRF7wL/fIQtZTJvzjygxNMZk7bPygMWu4HPv2STsayAy12AeYT9A
GYszMsx0U/qRQrK18KMrX5/owQ2flID4b7TX5UyC17H7yvRJms4xaCVLUuGpPM71
oHK/ZeyLC2NGHP/vwpFiTvQ3il6dvHlEVS7hdMO+VaOq8Xf03MDFEdsG6nTsaMDj
vKvPwTOlYB0Xa+jym0pzmG7+bXIDq6x+oAqESM20yM3WvEbeqcK4JUcX7kZdRVFK
7HKnIOqp4rD1t8EhvBw8mMO5n334Jb1hhc3m3D9pqKyfqkeLJNzcBKrKCYSFiwSI
ilR6+WhCuriIYlChTUmru4V5+Lk2BK6dyJ7gGxmjdosWVqgiz99Qm4GBVszGP0SV
h/taK1Qwn0LG7GK9wlJmBQDEenlBjsaR2h3U84HypwnUMP6Ljjc+F27KB5FYQ34W
kwpmvDzgQNhegkdnaA0udcIgkSyyVCe6tJ5Vsqc3tMC4IYClYwAYvtfG0dITz96b
p6fQ85mAZGtZToby46vv85yi7rxi7RDUwMTfmhm23xDosKLHYw1bfD3dpWwG6k4x
JwANUzdF4aZqWgVRoRv76KyamuAIxIalvDUVN89UMQzU5jSCeT4EQC+f2JyybKEu
f3gvFUuBvU7UgughB14bLze6FRB1ePSPp9IOapGKBwDhXxV9bT6dv9BnjF6h//8/
mm04eN9lQl5VaGR1qc/Lcynub2gLeLiuN/AtJsYFH1UT7PNWg16WnmssZKBC/fcz
JLjFru94c+6ywQSWJYdtAXLwFW5pj9wDogfiGn44K7GYI/eZw6jEbESXmTB90d78
Zd/xFNupxNdDjZhtv73pjtSXjtTrTlNbxaVrT/6snOgqkpVrzkyRpFOfHuAADa5h
H3c8HMsRGDEa5xXBtrJNOpgVb281E/T8yHn5UVjwanIF78t5mio+Oqp5OpN1SykR
dLT2s7mptFLXrDZMeRUVMv/QK48XXHjwrFKNcjTTFI4/vqh+uvFIaPOWiDGniXeA
YhWSCznasJYD/h5wtYvR9peNo6UNb3A20cKnNUKPCyGgz5CKgxLB9N1rj1B6uX+k
K1evWVNJK2q0D72dMMircKmxJ5/gwjN9xW2dSZId2xKMx/HrZnsS1IY6/JxhoICx
BKg2j/HFPUUuB2XYmw6ytctxiCNp15FbPl1XHfNMhI/giJez+6ieQcLcAYTIEE41
8YFGJOjbw/M+fGWZ94GOYuzCovVFQX84ryAaP4JEjQ/LRnuVMrHrxiehlBDpidgR
bOCK6wtR1TfjzZ4lLU5d6asw8xwP6wiG4u/iI0712pG7YkUsL6RxXnkzb2HPUso+
K9hI26ukZnMt6R8Br8NYmMPo/EA0ufcP51cMh9sLepjW09TljpWTgwQwMV8EB4QK
FRJjaI3OyL2GR8f5E5aYvaxuL/unoLUjCGkclN91hds9eF6t0wEYo2Hf7Kx5KwgS
zUPvo6EVfWN/UKfW7rRnnE7+oIwS7nXbwp5gtoHj8AyHd94cOpuX4Ljp3GDTYydz
lnmdpySfG/wQfQmlwHOmCcjtolzf+RmOJsf/aN5cjtxrGvFV1vNuWTz4SoLSArbv
Cn5giX/hNqku/LA7IAbAFgAEz63bHHkXOTJAGMR3hwB5WtNat0pvmFxC6j0TtErc
75ugsHA/BRlyKXtM6+2A/CiVCSLh20d9VO7s/5Y+2QQCdanpnX9/huhwMJPZUpNo
T8ob064nTWst7MmbP8xJjZSIrc0afknH5Yq3BAWcWfZlyHHXMMOoYuhaLEQ0IDlr
GyJU3Mm2zK9Ter6BdV041V/ZwcIB9jo6DxFjs6tPgmdrmuirxjP+CIIP6Mm9VYYF
jzkSvGEgdB6xt/Cewsk86mVJff2HdoegddhK8PG5DfB9vwM0ZfivZKq2KlQMu2hR
9JijOjfsr2n+6ZiS0RZRnS/zbRn7hqLEZBx2Xh6RSbmRBx3N1Jbwt6Pgkrvs+KP3
u7efd2dQgSD/TnBKj9WqRlwbzykenVWx6j9pZroHRHY+f126x+Mw2qbxlhrUbhh3
xTS/DJa2kJomodX4KndEXvQg/2Y89R6fXLfakc0eB2F5QI/X+G8wcIFJqq7LraAp
GTETEjkq2WhAhhl9MsUMfRNXwMaHNMiIWwJyRjiK7inGI9r5EeUMGqbacsg766m6
VR5J3sBFJnUAOsOl+r6c3Ov2anzmW/91zxcy86K114f/1AcXJxyzMjDneOTGRPjO
nW23h7tCIdec3WZ70dypB+HiAY37ssWD0eXTFPAngeBQAfpUE6zENEjD2alKKHNp
0DQmwmR/O7nCatjUYz4vyCpER/7QVyIKBcJi2he1tpJjrZeKXMi9JjewJFZt8/dt
bEC3U/dm7Wl8f9nlzk3WpB5SI7JwGlTDpTFZwa3AXCRAwGh8t7jYZYX6Ry4QmDYX
8+DKywiIHhhXZiwaeMWEHziy995MUhpnafrWAkBUVlvJbnnyzSns88mbkLt0yRke
W70PVXpjXY/meo+k98xB++iIwGOIpPlFxvOwrgy7ocF8z6IQUgo7HLx1vMlh/DMk
Qg/S1we/E50fnbaklQ3yi83b+QSXplt6589rAT/RlEGLF6mEio4W+SpIQgIZuIg7
m2xDLeeW+N8YTAs4T5e74sKY6x/z5TKnOdzuRHe6brCFcTvIGcxtOWF9oTNFaZhJ
wgmqzcjON8ja7RBoOmj9gNKe0JFnEZMv1p2nbVsmKsl4cyO4jp6JzVqymipxbbXc
RSX4hoKN9Gw3E4xaFBJgGsoqYfCnelDwa7Sn7tef14SJYxUEXY8x6NYsESwlECCX
hGQn2Dg7sHImL4J1gL27W0fEoTj0e/B1OsRXJcMzhguWCwKzw9d4WVRg+G9Kgl5B
sy/w6XhdSMzA1AE0byHyA2M0a8Ecpz0MceS/S+X2gcnpFbYXdwTWtdZn5L1vCmJm
L4/T9rWIttq5Joc2ZcMuuE9+sVrfOl9S+nOswjPCxh0wI2ySwqF1YM+d9dJV2VMb
WYFdw7Bm1PFy5TQJrYWYR5m9GTdzE53vHKlEvSWn3hnoyOUAYvhazsmMy/w3htyb
SfUOLHNQz38EbyCfdjgPVCP+4ozm9+Ad82Q0U9AxXA1VDMTzf+GSce7kyW+9ik2U
XPz5jqa/bkdSKfZTlkn5H9yA5AHoKS7fNP84lh7Xx4eOKBukrAQRe5HyrLYSZ1E3
eO/YF4HUHY4CAXd7FhChXjFx0qqIcKTi+Bow4wiNiis+WIUvonvaxXgpKNAWeMfd
9FD2pDLnAr6+a9VYbKs4EDDQnPeNkZTSMLf3jcIYVwK4+0c1/olKhiN+3zysicoy
RcqsGtBXdh/0UANwm5wni0gxeYuL48iDpw6ltyqXsyuNVgwwHR8X+5NOCc9+oqYM
Vx+ckS+UNVwOvadqUNLUosoWY/sW/NEtrThM7ysfMsmg0BH5Od9Y1kX64mUs7RPd
H97J6dRUwIJSz5VzyEfi+vJFpWCF9eK3c9DSSZb0RaWzo5JtnYivgCSIOXo5GYM2
GjKntuzxZRtM+YbtgYkr0y4OGsLqKuqpzFc7OOT4E0x8yYGaDaV4XqJPyJyLr8eV
GwWxzGNyhcmiDhrs7wnZvZtkYu1QxJg4J54lUaezumjWPnmT82EXuONhjnoagPSi
EY0AlqQUq4KHlaSAV/mbPVcH0CZr5KJ+R6NSVDBX7/xzm3DIi74+xcmonSaMFzuQ
RCrX0ceQ4NkQgz7pEhJo2V6Hq5wpW0G/c7AabTkTsvCtW8xUoDMxlYtMiPFrHIU0
oA6kBgJvYwF0tbTiPlX8FmSnp8ZHWTIulBXVpTsxyjtssaKeY30yFAGqIRkyuI21
yqJtTyT8BJ2NBve+AhwSGCdF45o1RWC4um5bqTaQ3DYCrjho8REicMpJ58tRKKxt
e95PwTaAlgT1g1X3D/1SEh66meL2/wu431o0SML2axoDiN/jibSDRxoyduESvIew
Mf48Xojgy9QyTY18TKV2itOv80AEqvcbd7yVhECdtbFmGMm/8ov4IJ90iv4C+FwA
FDOu4+udesf5F6RTq7z1rByeT9KOXFJUH2rT7w9pHCBhTOFPWalL6TUGQLjVUa5u
kOn2Cndgdl+VBgvmRpxFZ6zOhMioUHQOlnnWt6941pXZwrd923su9gxJEDyQ+zAA
LjhWrdWSRSEzvhtcZtSEkKU+guHPUkWCLKcYHCnAhRsrtyDbsGzgVPkqXMaLQnUr
sBNhpBNF0LvR1hWdowVF9mHyMP9fgp/j2MwTOh3A7Wh+XaMisJw/hGVup0NgzaNe
KdM3LyA/Qel+ZQBg5mZ37fuCcWMj8K8AiVrPMagB1T6gK7IpFM5F0UmyOye9JCq3
rnBXhTfphjn90ctHlX3num0+3SuEKqxsltfgC64D91CvKLyzRCQz/F4qPN10990P
M7tUV8flGOVnEnIc5XS0XPXxb/2NQ/F9wq2ctGv0PVwkC3gQ99EqSVB1fHJ42vrA
qafKzAJGN3VzAs+OxAmt3EeyfQh9CXJ9Q19nU6gb6ZpvC5+q5GWsWc7y1o0PBf94
fAbZkSDc/lNwC+Wmg6AdWiXOqOeD7Q68eGK2iE0j/PLwW0nriVEYZTZnXCt/psLm
Rotha2Csgl6MAZWrTaqpAI9eaw7fwH2YhjEodg7gJ7Jz9OnAIe4Eo+4eKDIBw8WW
oCNMgRs4DSKnpFwpd8Usk44n0AEwavVe8udqPERHuE0Okv6mu98cWRn55KhjWt8r
Awlc9OCaftS+PIvAhi9ryXJytbiDEsaUO7HhzIRxzadoGgGsZ6ifQqcVktmpytfi
G/5lsxEg8fPqCZbBudrDIRcBS+OQ63RKC0Jc1yL8G8+WiPPZLYdemDsLZAus7FSZ
OtxbUz5pl1nBG+iLYQwlx70+lUYxhLw6cQl1U1FAUW99ApHI7zwIhXLecIRyWugO
FVZeMxWo7oZZjgqCsji5TTj57zXUOKRoQnSeowH9p+yiB4CV6DXuBsSr7AOnRvmd
PXKSfcpnD8MJ/B/dqu+bXpa32vbWQnta6+QB7tStSGEujQKsxUNVzf0DaP9QMYRz
T5fV9GVEOH4ew+f4czVpHwlq9G/Hf6lSRL0XwvJE3GZafv3gFOhQnfMcTJiZLsqz
4QWcBIVP2TNYxjv5ExSfZkyJrRf7pEgVoXGnYxm37ZeF12pKkxaJJCryxOYw3PPN
wyEC2S36iTzkhsRtpSHL/6PQ8a83v7gcUOw0DgksDKTR6DVJ4TgI5+ci/8xMf5tk
UmsNKNGwKyY9rCyJ/S1tJjmlDwcrEU21bpBJSIWZ3cnLuJXOWfz7cAYPInGb0vCF
ckXky28ss9xCQMSZzo/OaeT4F/7qgDXFimhbcf69jvvRbO6xo0Am9kZDQAOfGuad
B2MBmI8bRrvnG7FocwtmPU3DmrNfQeooDhWKajSxYV7dbNsvGGS7Xe85miHM/eQP
Um9OQn75tBzMAZSzQbW1/mAmipNkMBZ+q7mY3A+Zw+tUxhIV1qQihRzNklF5mQsY
Q5edDfNroK7vG6Cs4eEz0N30b3NLoRdKykRwuAu5IhiB9v3Ut+aPGj/A1qVIbLxk
RsZ7RlOeo+Enf7FxTcmZWlFKQgU8f3Oa3BGh3/oY12vJe8utd7viIGUS4AowdATk
KdD57MU3wTtjy6vBA9aYZanGUaSPhpyw5pYRrhh8lnf/E7Kllh89OOav4gUppCen
OdQDlY9h27mQrmaS2ZzFsMWCb4OwpLCEr2k9sGkz5LpTVyZbzFrymyiRWYTOoHKK
ZO6isH32L9Gwl+gvFVQiitpz6PsGD1rhGEHDQI45fE/eKDSaVCeG/gvrjRgGGfbU
g3NDrY1yGzhJp8MpNOEXa2ERks4z/KLzKfYjm5tbo880a2bM9Jf8Nbg1CyWcFdAz
jjSpMBXlJ+0NNy5vzygMOU2fuwEb+fYQjSMV0wCxOari7cZ8SiZHF+qKc1180udf
+maWywmQjk4qUXjTzBxPRUBNoouVvy8taKfRa4zzP9AeE+C/8dKEAi46Qfn4jH94
g1RcObFnUefBGW1rFoJL9e30LkYSMd0gx7AGeaBnyYhZBWJb/sE+CXqM4cdXDjdp
b31myCmuSUBqOxch0gXMihLG2DSg4nJiYq0NEIxHCnRmqpOp0GVApaA/Azwi0ATb
y1g12cfcD+3yq0Y/lsy6md0MMflqx6Mew63oI/ybtl28RjWoHIokcN480d02W1sk
aeqLmoIxgbJpZfYnJLf5Lzxztq65ee+i/oUYMisYWt93/11qSG/RUmGgTMx9PdAV
LlIhto55Q2QSJ/qJg59wMkYD32iqtn1tFavywSTMeIWDo5cnDfeFl4gYO/xdpuKF
r9WdyblivhNxxnIOsKdr7/Eh3SOIEct+z8qRNuJ+A3/aBBLctjxyGTOx0aOrjWCA
jSBbK+o+P+SrkOuNk7nohvx+FdahBcoGuot00ix1k3OE/Fjr1oXmXBthRhBOPMk1
xqbA4jlJyKNPIlUKtWWjfXjm/NxepRiJBisozXIaFeW8ssb2yG9HIcbf881PPHBM
ed8MJeXgjQZRSEqeTRvcxW/rOV3YX8KX7p0oqi0Io3heJLViDgB9qqvBAFrpz3J3
awO14PJoFcXxTNBh4ogrDC7DN7RAvmqaomoVY/zW+qmRen2xdNQpcY5V2SUib0gC
T4CGuBEJ5iFKNJlwwM1kjhDseIdxDJCgfdgeLPQX+YQ3ahJnE/6mXL9DtxOhQS/v
wjdFoLJtuHiKLMf1EhXwpTQlHf/BZ9drt+K6yREt+2oOi1f1QlvQJVIds7GNKh4Q
BLabKnGoQ50ZeqZ9ioh778GCyyHEW6E7WSreY20AEaCJv0fg7785eeW9LWWcaeP4
P9DVTzbf9FKcBsee02UejwvYcI07kgqhjtQkYayf2vZKdBk5DEkAqETAMiviQdVR
OJUxMl74z1yCpd/vAlE6QuDxjIhStWHyWIGx4ZCd7spGWlMrzxEKeOvJuYnt28gQ
H0mgxoUq8q4N5PlGfMgJjBRpAuRVUbYzdPW60/yhbDVBeHpuFEIIiJisKsV23JHW
+DNfVnN0DC/l+o/gdWvqwIw/dUSxuc3R+E/FRHX2cHdWTAeX660adEShhz3qHod+
rm/Y+2YaIFkNDp2A1vsdGdF1Yo5Iia1gba8EpBJQsCK7bLeU3Ca3Pqhf3//vhpWT
AVGDu62M9RO4VcK7YjDzSTuNcSFbJ0M0CEJeC1kSMaH4ZQnDSesV+8BAhp56PSR6
C5UM+Jfs4/oi6kVy7uXP7SxsjP6vkYK/RYTGQEoYY7R1GodpiIZUCll7y7pbpO0C
u8+LeS02kKR0oZCJdPJ9rENdFuKTM4nV5nE9pRi/oTrRNa4MOOEAINJAj9H5ouel
ijosFkKj5SZmpyFO5aiA58RRaaTbmcVST7hLexPDzxXB27NA0vFsO4g3NYfda4IL
e1ulPcwTL6WazJ4oz/SyLcTAQWk7GjwWwH0f+7Cg8x/gsdh4KDq/Rm70jNAtDrtS
1xSCTELzBcH9yJ2XsJCSHAqKJcRo/kK+j0EXP5DtTaW6b7iTeMtZpEJsyQpoFpZ5
nJUkn7SS6z+H14KUWb5o1//f9kek9y1bE0sXcYiGoKmEGKWFSwQUPshxCryJxT+x
x38/udHfSLsrsiDSczX+n8wwNj1ImqqNkHf57jvHIl0IiHMG53pQiE60YvtanbNh
5PoCg+IyYfd5gRjuDfz0k2TL70p3Zk8aP6BBCaQRbEIhQvONXnq360i6Jm9y4ViG
ANxBKx8Kzsm5mEOzMzYHLJ5709wb8W5Uj+1cnh+sjOEnWRRJ1710WEOv+UzZD7Sy
S8az55xEcGzhmgtk52EuWtdkvtmAwIy689L4qbJhma4TewKDdYTE3kfW/4CsBRXg
+jeyQaHsWREwosI9p1Q2ZB2vbPR7Gy5jQKt31vJjPzUMJBjBQppsL6x8VWgthWqc
MIZKUyjSZOudq/lC6QqC6q5a3Hj8KKIOH9rMvqS8FxTwnqFB5qW9pHacRMegBBMt
Rk6PdyhGsolH4UaD9kZm2rT9RYXUeeuViYvp5gKaTnceXSP/9zTDW5IQ7BOTTvW2
zlsbVUqZlVpRXufXf2wxS9t99v2eTNYRkWVWAeAcsCTC56iuccr4S32J1gHAk6Oz
I5kmtz7DcGja7lkkiOtgnM2LcK9SflzTFkr1pqFMhxBlWkhhTI/mAHExfLmTBsww
lCASMLg/77IuiJ1c+hPLim53k+8JwBn1jhvGCnAyMgifzGBQOwVb4Evz7I/Lrdwa
RTfy6uQp0kMuad0NDtexfZdTJmIR6FSLpj3dBiu5f3tfi/s2J//l3X0h4r+hkXL5
mP9K4blqPZk5kIOFXviTWzLzxu4c12HkPSvVuiJyMunPlmlcrBuy5VkUDi1+5kGk
3eRNjmUTzZun05M5vEYwbqik4k/IQf5Dgmlfj7mucFvj0wZolck6hsXRTzQCjCQT
Qk6jcGhXentMCR2dessL4p+dN4Q7G/FEnxbt+JdtWyeJANl4psO0wyDv0gg0FR/R
k+57iVxDenP6qm2UHz8upTY9qIlL+xdxUkEsF1lZ1ipZlfhcFQAVD9hcy6Tzz4Pa
o/IGser36rgtn4DTlGKv/yjFTrSMTqKxq3jws1ZPgqPgPqeiw3kBz0jBOiVCb7QU
ISfrvLNu9n7eSW2mwdS7SKLUtjySDb4e4PaSibx/sCaRQvXiOl693uhMUSD6cJ4n
pCIoqPbT6I4F8n0SjAM7Ikx8N4CPVEIebegYJx721zvP8+eYL1c3VwBTO5Nc8Xz2
4Kgtwvsw/3sSCck8j68tarhiqK7VlULX6EU0RGItaZTfu98517dJJxXoNbYLjvE6
iqF1uElc4ymuagRjN51agjdOw6/fsy6Ll36DMl8aCzP3+7G9pDeb5Dxf2/FeHMaC
Rlb1dFbdmnKJ48+hvmtoPYU3HKQ9pxu98QYt/VAM3ind8fOGuc5TR+lCtzIQ7BfR
5DSzThmLLKoj32oRm4P+502oL5XY/pNxVvA6PJgLchm/6wPYEATxonGiVzyCcpax
0MtzmJR6vSUv2mia6GOJo83F2hJCb9bIsYnSgBcfdgjGjfHh9Hwp0U3JfQNdEg4h
S0cH1301ujtUi97++HzyDWO2X9GrA7TMhAHBUyVWhMksvGMaVRiIWaatYBf/iMmn
dCxGUIjFZRhwj80h35R6Du+Lmo8zMdT4wCFillgykVL7IYTrbQZtDrMxNuzGb+x9
kqa5enLWZHrN+84fqFEONETzrs6tsImGj8Va02hMZEazg4ke9XFdEYhdRCgRzTgg
7xYod8J1tby5ObIM7u4u7zhlvAIb8pZFgMoukN77yiXAdfqSLkutC8BVuvgQzLxe
UFqlnWrCIJw6WYUxrWcqLW8PALOTy2IGsLui2ur+YcHDDlSfmNJP1G/R/YxYnRFG
7Q7l/7NgzdoroYej/Bsz2OF+4dqUVddPRYgEMQuBOgfYFqcGjaEtFCcKGGBRIeaA
S2UHwXHhPVTkBqrnCnee00h3zNFnoP+o8MbdZOF/Z+8NCdVcQ4Afu0JP/TP08LVP
P3+m47f8xWcgMbQNuuImBEd3SIq7t1e4GzKZDrc9WmRZjLF49uS51ZBgXvtWZDA0
ZHkalNMsuikfFYdDtZFnnruBYKKUlO9Ahz5KNLu5GXBlSR2/slWdl1ns+LSgvzsX
85+lRK4GNM6BQcfZv+pQ9ZbEfA5qzJAqutw5dQzA2rRMJEgIPMBP7eGKzFyXimU2
C5zB1JQ7NfjtnzFoTrbsCuDs1129Dul2ZCAuhQHDoRDF0GAQVo/HbQELN0K2xxIu
n5BKbkEKUTZ4GEPPextVhPwvubIimAhL+jldwg8x0CwH0qp0Livg2fiuRQ53m00x
E4BignIUNk5HLIa7zdYGMcubIFb6pHWXeIHAUZIaYsxSkjO3v9YnD4nqUG0VHtmC
v8MPkiGIDCjunzvFXahtr3kFOPxH78G7mgFG9bcn/nwGFK4jLCqsWb5E6YIucb4E
JzaAG/yperHbN6A0RRvUe6nv7/900OKSPhr3tA9jQU3fkxDGxstyFefoP55kfI/k
ao6GYEwm3bD5ido1uRePxrNS6NitAGI6Qbh6YP+xSFizlhttGggdXitRYo34zrsy
TGiFoFCRmXqENWpkCuBJp9uPoleDVYFST4lffXP71y83ea1HQ8sCbVTNJXpIF71G
i4bOREltUxG55/uGWmNzL7PQ8qp08rfa6SObKJz8jEqrHnlfb6lK4jj1QU156c7W
RSHJivEdO5OH1tyX7vv8a4xn8UJM4gSU7aferss1Ne0+RquwMHLGR0lPL+fTxIlg
oF0Cx0fziaf5g46XiJsSJLBCCDJMLLBtgl/1dypGW3slIEBuxM4I8IKb3S/JYpzE
BgUkNliXqKQwxHlpFk668tIy8Ts306XX8fIbbDY26XLoBLNKTB6Bqs8/NgPqmbTd
yPGdfTIrmWTX4kzBDy5pbQ7RSRhqITNatOju6nlz7DJvueNONaiMg3uD88n1ddOP
veUDnZR/XlnueVGExT3Bd9+oV4zSM69QF04EcepYaVy+RYJBpe75ZWhcrrhZEM3W
/iqukb0FE8XbEMdGBe3Mqh23m68FTKNYTOzT+Ws4Ls7MaPb74+4dclrxLaHfrsx2
5CCo9HT/E2rtNAR7MaI13NCIxVncR8BDuYBBO2wzzO/p82rA8NpWqnrTQO5XZl3E
nW21WIFFOYgjafb/+BynZU1Pw/K9sIh+LAT64CE0ttMh2khdlikRH/oHZvWTIskm
eLIYTNOAZzczkhtOixzCfnn/9RUUKRMG1B3DM32kWRGnSQ3cqY4QyLbwfQEM2EDj
1rBuTvok+VppUZAKUtra7iUHxKihMkoLIEa32KUm1EDXkCdSizpC0PF1PMogUdPR
Q2dUKg+9gVYQ3zvKLHfixV9u4ZiVKaez90I4d3PX9lp+EyYcXNK7G6BCkg3chmd/
Nai9UIWAy/c7QwuvExWaVWbYiVhwMNuYEJCqe1t65nLdVNV2+nX6w2ePlH2ffZe1
QfHhqWtiIu41YAqhI2qCIFrEt8TKWnTdNWiS/y+Q6Vq31ykgaKC041yC94muEe9s
+aPYISCzjch44dPT9/mkbeQXZvXk2nHY9S32vNISCw3GjwyYEJze9nugLLzRM5Jo
FNQQc+EjFdfO8wtfIbvkBDVRn+j5XuyJ/OJGC2qzVoTHDI5RmuQdXgis40pvF/N6
CuIDsN49wqgmW2L6vbT1cWju7PsGCySRrIZRmAsZOyDPUAb6A5io5O/2Zb9pT2Ja
KM7/c5t7zi8uzvTC4bbyTGiZ0tKZLKrH8m5ZDfhh+DvYdNRqOxnsGZFDfF+TBvF+
rsXp/63vNDzM2z7LTvMFNupMCQJlfwaTFel4ryNPDr0CreJlCPCtA/kDlz8uAyrQ
tnZHW4Y+mp5kDXj2FgiGCpCvZ+2HswCmIRnofP/KViqOk/GXawuBjPQTkuXEHbl/
7D+XdE84EFo2GjSXDjZbSrvQ0AHtmzmbz14nB20CpaNtyojiJsNNRNTKKUWp6OnJ
IBVYtakecyKv9YEPbpdCdDUaCPOIu8RhJLIpOlrzlWrqZj1AWCr/11XeCEAXdLbf
WUQ+kn2eMb/dgkGuPtMD3v6wcH/ENh2PbeNEbJzLZclEn8jQOs6XVGsbQa0pmXBx
tsuOpiJrVOFuK+tlPbb4lRaX/Mdj/nI8MWtL2SJhHPIVYWi+ielCAG7jKTKVKzuG
YV/MqG7LiGB3kKbHNcavnjRHtf5AdiNKAWFW/UXtbq8KKl4Ffwg5IZYJxczI8Mv7
D3Vs6DdF+SrEM/PwHMHGFghYsluTFGm/gtVG0BlXXPznZJlPE0NLIA2B3iB6UOCj
OgjKYtQw7JTF9BezT9atizAhTlhElMcQGDXQe9iijBRpeLKlvT9XFv9X393oFUyZ
Al17nIpMp7739I6xe4Iv2PCrcDzGV/W81sdcCg3QPGSZKuw6FaKVVTh9RQc9km4X
/q79r6hEjwOly6moMY2fYwRLTw5gvEJ+zHZzLLesap5Ua9OYi5CaxpGJr0qkftxT
5+xU/9bJVOwZysDKfIwjcNVJL1rU1HeZouCykzJXl7mOcl7skm1s3slEaL/MndNV
4uatawKdQZUli6BnZN6YoI03ud+8uXJIm1fbYjSxgFGF/3k1j7pxMxDMEUEk6JMB
+Ywv473m9nSd04jyxKSiAKtVo0584vxpYp+zVL+RbY+vYU691l9cb8ZUxAR1R4Al
GWg9Srqp7080lcOr3zSojiywHw2vHqJFm8Sg8cSnV/TCpY3KAT39fygHpBEDy0r7
fRxm65owYXuXWsurCOFwPnYjomplWj5YjWYx44L+cauzkFNqILQ+xu35g6TQ6684
WW2JixUfYbiOeu67pZm2EPYfPierJ7HCbN5Szu5X1id634tt/t+UayA3hoeTL1As
euQtoRBqcQN8Hlaic8H1ZByb15XTEX9FR/D/pIjQq0tOCA40l/SMk2uRxWquy6BW
XqBA1UuTxsu7oKuRWGqbXfiXAFVeO1mQ+vWKQPct8KUr5VqDesdqE1ZD0o82nE4Y
5ajUUVBCOBv2wnFCR9D1QSgMMsh1/JNwNV0IhAiems6zbHqAHF7OBZbXBjBcs6+A
cbP9IlaFY2QBBBZrHazUhnjGjkc5xfgPlg57dpNRolYpkt/cHy9FTtH5VaWYc1y9
+Nf7uaxyeaPns8TBmoCruDKbl2apRbnTkWMa+793VrBTdI/961UhHjzhEef6p5Cv
eA6atDumn4uBjYHJZBhG/yA4rdYaIsnoe5mYF0hkeLf/x6x+abNbvL58bNXGdBtL
UTR4rmgAORXzQJK7qcZlIw06YyGRAuWZ4tjZ1VMUfzOVUd8qYeaP8xU38cCHKvTZ
6p+Am3FkA+6W2kPzr3J4bX9aKeCUXL/YHIiEH2DSdDzuEOS7W+OUAvTVvke5vp8n
1veQYzaK2Fu7yz68B/0/RpMJyOTykVhqQTDXfortMk8AnF9PjA5unf+42QGbkHVK
fSmCi0sZ2VOPK0f8yp/IULdCjs0fpYxqaZXrJmlbiHW0MYon1LrX8zvPAQZ8ncpe
mnAfO3TAHkryAn4k9C5W/HnKQ6+I2jaON0VP3WrtqzHVQ3EMcPXkTh04yNf2tXWY
vx3lbhmxU9iytIl9Pdoa0bvy3z3vu8kyMAWAOnzCwJwdcRCtbhjMf4OcXVddT/wi
lz+siryEj2voysuZwFaq5Vf8X+rUVErIpFiV8O5L2tK1Rp8fktO0MWbDSssc6DjE
3xzaGe4uG4u4fgJjHWokSTRJ7lndAa99xF1trfXZDBoqixN0QeoqF7o3I5l3IZ6c
pgEB4JC1P8yxuGM44a5PBN5j3QCICagEqq6+aOTXfz1IGarSo5n1FY92CSk7nxpD
+ibVXPWgfply1WbnCvbAlw+qVzEjRHzzwviAiZRK/oBzWNrGUI0Wkw0Ce0BMQSHE
nOtGBOfCaf1ZVwGxv/Ik0zuNguDkiqKt5VuiErfoyNoI/JHDw0weUQSMx0Eitm3R
15OpzNEr1R8vZDtCa4QBfRwleXXP89N9ceZsQvtxPfuSgHY61aihH5usP2ktm0Eu
xq17Tjjr4QEVHLRDC+Wd7FkGNIE2q2Kn3wFUNFZpVRsQKk+GXiZQxPz/c6w+PqHP
6jjNwDb+hTTngSOz6rRrVj6HqOIJ2CGTtqTTheZ+iZc=
`pragma protect end_protected
