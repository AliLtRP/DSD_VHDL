// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GOCfIhS57p1sH8jreTcmubbsKLB3vSbV7b0ljDXXhhWDppndaE4qfMjTtWG7Gmr+
Oi58BZ+M1J6EhRCpYJYrdyk3ctLqPg71TSQ4dxt8sFhAGGT7BQVWBEl+qdPn3kB+
DjwuH5VaH3+c3tSW/6UHE2u0fc4kGmoCmw3+KbWedCE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 86352)
dqS7n3B7UM6v5DQZmzMFwqLhJNHdeZMBUXDlM606QbAzqRYZ1KamyA8rJdcszdiT
CpMUxjOxXxm88s/IepjyvMvxjurkG6mZflNC4MyxdT76RyAlmXGGEpNUlVvlFJVR
88Ja19SrsjVoas97iWv6m8uztMYmvLWdqrbbBqWzMRrsTir8H3MLler9aXaVKz6Q
FNU4pfcep2N7d167t6e12iBfvtECPzsP0Pyh44ITNgoFvYsnUZdtU5RBfNMs3AzR
/QAl5JWqoJ3Z99nwxuuSF1aPub3gdYu3RKu12FyxASQ1PnJ5MSnP2+bgllyHYP17
VZ1Q2gEpgJmjagSXeqmQL1zoeLf13C6dQw6G2isMDWQt+QBfvHcDi023M5Fc4m2N
J21Ecbi9MUa0DxUPF+2cDBo/HHPwpSG7hPFs4h7h7Vag6gE0uKN2jPWfckDLOiYG
WqIaUSxT2alWTq++wnX+B1DyzbUv3hkUmWJuCHVnu7A62IXSG/KQCQ3W5RmPyzaB
vTCdLHHNapIPD/aIwwGdClbnmlZhXdL03o3n7aIFl8KUKH9BIkq7NYoRYvgp/5tt
uhi4iu+Gv6Kh6uRz4AKfoFMtpFg7ct07FWFJeugM2BjnsM95T4Gu9EXQyCR/B/qz
qlhoWpC4GWwvfsNFpOMKVyLn4uqor4GBu0r6BlMS2ru3yWQBcnBAo27I6iFxUq2o
uZkP0f/QFsw8dHmrGCPSzsx8zkIYhGISGzz5amnHk/XhnQMVXR34/HKW5KGDHjsR
XCyzSzuhAG2j8GTCPksTZgN2IKk0Ex4bVF7/rjUnsPmc7RZS/Quf0vTOdNpSAyBq
Nycd6gAvfurbd35gOG1uKqhUSf45KbqV52wazWjVF5ZGPIQPFWMEnLn1N9RIZ5Cg
V5DBLs/M4aKXAmxAEzYHz9ffxye6vIfWIlHLrRqPbjM8eDjzeZ5CLhu8uw3SfzVJ
RqttRCYgHGkYg5BoBJK/nE+sHClSevVePS8QlGDSNO6WakJa1NRbTWxQCkKhJ12I
No8sQJbWA+diPujEjoHmQwtvfii74gG4Q+6c6ZlpH0aN0GiKW9Z49QiGze/G90nF
hQjENoXoFaK5hWnKHlV33jbq12NTxkCi5p3DfOH0mEeamIbfOxhWUF5iZBnBfdRK
p8FBc6LIJp/WZxWSW2nFhXpJj4RYWGyyQmLh13ypqgL4sHN1Ge9qXFKoOmghajI/
7cfAvreQ8Dw1HUHsIYdbqDpURdtOLze8jwoJzI3okEcK4bzizBKAupBj3QTIFyDo
UX3/mZ/2cgvXVZbL8hUVPRyW+7V6enXTRzLbMoPlmMepbFAD/KMgkg3XE9a2AL1s
X4fnATJhmsK0o1I7B/+mfTf1QQzlN9/8c5zzQF1OETu29lH7jT5sRRuWr7O1mG/U
bKjH1LeLuYbFbwwHBtysqV7Gr8n2h2Y6oc8FT02webqq4j72BApDy/j2NhCpvdTm
ULhlw8b0yv+FzPnuuwLPQkZpmwPBiq5rKK6fvcAtZHdh/aMkErDZZ/3QlSsGnTqe
cNiiQcDOCJkh8JT0eglKflN2h02ClQ18MIUOiJKMHnfk4lufDJEo+bTPu4UWPnWc
p8CJAzXNvoW+e+BoPQhNjiBnDwpOjBiMdd2A3iE2+QFyD51iM/sNVBDT5ixngxVw
TkElStwrwCigEIPCOdaM5ckwOd1/9Ju0/O9ivwYI/b8IEdjjoZ/mf3K8eg8OG7mr
u6w54+2vUDt9ylZVFDraHkNMhqBlE7RiQnneSc7ODBaouGj91CccfT2le38IMiGt
0M3qSanNGJfdqPw37mn90BfZ+YyeI4ogk8lutZfmARIUFff2bQnfZDQvWQjlMfc6
603a3+qf8L+GDneOxQfM+ZoYf0/Qagb4THd26LHtZ0Zc+jAY6nNPpsSnNxWXUk1U
HoS4VaIMyFg2Qpjmi3LOgw+Le6Mlw6mjOy+lxl84ZLYNrQWBfHmEhVNpMAX9kokx
py/9M33n7lgyV9vkfCSjVU5PD9MvnxTZd0CVMbffoEnlU1sSY7Ku+nCtaAaM3S68
C5h9hwRNehEHbreQ7SexwNJr3cGHUEUUUoWnawu8EU6DpjVMOgtOaetuR0hsEig8
wIWThbhfa3GsqS9T3VwRkoBujHpinYBOZyXXP4KlWYFO5h7PtoQrQn+l67O3qgG6
CIs9YO0xFlLxaApZPASLv/Uzt73EmBZxOdJ0UQEKYzbqf/5bq4N6X+5RFzNLXTf0
K4VExcGjJj0C5UH9NavNUkPsbtSLuRVP8jGc6ORCkprLO5gOJ6Bg9E+eRxQslcqL
OFgwsLoKHTH2hzvosAt/5nxo/2PP6/u37mRslneRKziAvLgxCRbZnQyWKkmrPvOI
kHUMJkYBPGtLCWqtsVmlPSwu1hD3xYySg7931C8rbJcTKFmyxfcVib3g4qnywLw9
d0tXYYzlHRq5+sxfUWARO9BMpo2DOh42+JlyFhsHKJYXM/F+RN3Vizg3MVweOFaP
3fl4kmZxeUNdOeZBWsk6v+g/Lv8pS9C6UdQwsNTOi7xShrHRZIkX7QAmb+hQc9uh
ZKME07SStFoPWtOvfwFVSO8zfyuN+D46vchIwd7LMQwO6XN8T/19lYLMal84NMAz
cJTjOm85VMuItpkvWcn8M3gq/4jpJeK1aHtRLvhG1XT9fGF0CUTXa7FntdBBpfDG
yl3f+PeJ3gBY3LnfNGP+6OjTUP3nRHkbwp40oNTTj0WitdgjsgoE/K5KPPjYyvFr
TbKRWL6M7dP79C1LPX6s44VKn0ThOm7GDnGznoyL9sxM9fA7HsbVOf40QLbmFiI4
cNNPDSoh1o/DJyMV+DL+mJaYUiNM9cwFHR3kccvJnRCwj5Yc3vsMLEfJXxTIhKFJ
O4Fr7zUtyF1P+gxh/c4irfaGRxTBxkHPd05HFkUEUe26zhn4wSSFNUz4VsLYwDMT
pldESmc3G53UGz9KhB88VtHbyCiQbIFf2wmlDso9lozricX5mPwz/MUXffDlC6B/
TmlXvuFHbOVo7q9drP3xxuajJEFNjMUoFLXp1pcV60jeFUVYW4zko+FIsVh1pmtr
qRydJE0SX1xusJIdEI7WMtb68NVQuvxkhXxiIs5u86GS02OkMujKxSc5jgCBaEIV
wFMdEgYCQalHfOb+wsZaOXcoIAc0ZmhlsSyjkxG3Gn3PKhpK317CHh5mX/E64Zrg
lt7lLMrbvyAiezQbfWEj3+9qi2EqLLw0CrpuwCPW+jrCVqtKZhpfOHI1cE/033hV
0oPN/3SnjwCIPBWpDqD/b9koN47Zxv3xfKYP8tU0/El0ZWRWjcfJQTUusbSq0bYa
NY/E8Z6cNYWhONTMTkSRjqbDpCKAW5J9T0yTllgwo782Iu0GY0QpgG7HyngWf5/Q
pAj7xh4/2eCE+nwShmWmdzqLWWbArLwHL73f+NDZ5aqDngOjDHwuWtR5jA0xdzZZ
432DWuXllGzIefsDLN+RWNKTtzYpkOwzYCqqGupkrX+41IPIcTKYqm0v18UHez0C
X9BY/9rpxbhBBlOT+kdewrhxhgKb3p9KswAjEyTVp3+3mTtkYma5qwl5qU/e6vxj
VLi/Q6GPLb/0eB2UghC8FAbjZjh08+wlInHmlJkcjSWV4cssmmqz6HMcBYZCSz3N
F/cyDT4kDcN72bVHiL649g6XllB9MnncdlGqnNQjuAuoFTjSi0ci4WNdOjUQAVJs
I6vGBeiEMWcEyx1fIKD93egmzdTbai1psuo731cm+oAVpL44cOfKcvunxswJh7zF
28Yarwi6Tu6nu1yZm9vKneCjh7k/3hape/Vqzg4VyZ2svcC16sv3YNwmIYRbIki0
DksqsdLHnumJJMi/mTCbU0RqN7EBd91NpZj+aVtVREdUFDfT25fT7TueOnNd8xBk
vAQkQJIeYJL29eZjzsEKYEh4fpIjG4w8p70lGx5MvFzbmNQsVvu29pIPq5NZOc/i
HA8a7Jpf3UiEsWQFyMJ8j57H64Nz23aHF+vNH/a0VQyq2qEZsXFDVym7OnwII0tV
hC8OfVB5hCy+syXqroSe4leeBuA/0KTnHVi1jE2ZgAcnu7CfBbOQ4XyWZFEngQPK
QEIWp9q4Opm1qez3k/z1d/sPbiXqt7vr4EYcRMZCncP1+gcqNl9h/3tfIIHx5tHU
IQGcWxO+YxkYtcKpcJc82xLLWmgj/K0DN4KFanLYW6+x4uxvr2LJYS3cQsV1yiZV
4cRThsA3dtSOiYinF95Pw9IfQPvF3sZZgV5yjoBP0MnPUfv6WhSz6Mw5eS6WXkS5
HcTVsmU2uNJ9mXWB+0r9bwaETkndocBPmjyFqi0y044TBa+5lidYmFly2ZBT9Kjc
HFb6s3kU3c/dDQj+gUh3yuCy/483//lQT8wPue5iFJ4/S6qr79crzj7cc1x9SPuX
o6Oo2pLH2MzKV+q66DUhWWMDgOip/oUt0p6uhF/8z7cXiqrb9Gq3GtFZHS+woiFL
OoIsDfrgQE/VXe8Jmu/1bGKLovQnmO+RFlUbmvx+GXD5T1D7jMFnd6uG/0CqO2i1
55g66tyAi3HIPL305BFik34HZ/EIrmk5iyrDAvW0d3zharZ5xMoThs2xxTv7gU/2
P1w5uDIw8hjUWTzb5dmJBM058BqI03P4rpO+VGOuZgdVYvAFQhWB9w52oAzfAF4n
ZAylmNeXUni4G+kig48NFVee3cPel0A3a0li5Sx6NxMuJyKG6XyAubTL7Em2nY8R
twPLg85bIIvT7HhSNyKtAYNxB27bWsGeXGjB9+vgupYqV4F0tKiXD/EJzaYSYlb2
u/wt324uYoNYRS3/aWEQHegSSauXkXnReHrnCTRpghl5g44ETDaGSG1f+EPFDyvA
aWKKb+Q7ZFuiCW5lCUZb2royKccQ/qqXUGKc+3k0xa0Fc3jfo0+4NfQmW0+cSpwf
cHUBN0Wr/vbAhRnNw40Qfggo4t/dmHpnIi0RiitOabNTUbXrELTCBQSX4izBI/DP
6/uyAHZgrdW1oHA0J5FWKa+PiNyEdlMBFy6lOCqc+1cTfqhfZgXuR220cgS/RJwB
fQjxvf5q8SVN1ffd606rBRdXXRagK31R6YYOElcCiw+IMvlTpa3CU31pR/tc4rsp
a4bhDynT2qtgETXZ1mOqWvIp13ZWVjkf4/shQj8nNUNOlOOctr7y+l+nHPktZw/X
8uFz2B38cTfqjic9Mv5sXM0J+K94SsOSJd+8InaacEjSgVh8n7zwc0SEJU8we9kc
z8hlIYzv9zYmUASeYgwjY1oaVOCi75kj7jaofkFV69sBHjkwRenzLtw+lPNKb7EA
/9U2sNHe+nXhyyIbXHMsoMeIm5XoNUl01VFYHgiUA4unDPo95yY9wVFuW/3g86Uh
LwYbMI3nkhxxBfmjEN0TWbYSrSXBR2aLf0+dbpt8vNzrCdrQ8aGnkpuW7PRyKdmy
I/lJgDdCFJjPKHINnr9O3sJfGlp2VZixi8BWrUb5zvpKZzgciXLpMVLBxGjcDm88
Pg5pvBF+r2fC9aEDt4xQ4bbeN03k5BhmZNB5C7Tlx2euIIHDbACe/PJvVbIzyaIc
QCMQr3KuNhP3UfKntJ5ei1cAzy45QJsxlik4qMM/wyXl3cJvJYaacc2L9orlLUyf
sKkEGKtUfgfBRWzCwtQ9d33yZGTPx4HRONBs/dwCw8KFrHOJkBIESrP9NJ8xgw5d
bZGIQHxyc22jPJ3g0VPCj67v1ofWw0OsL87pKs8KpN2ZseiMGFAVcJWr0loyEEof
ZWs0Pnb2KT91IC21PsH/XHV4tmG7kAWhQkJND6pjP3GXiSRQyYSPJJYw7KFlAt3l
6rtAKULa1cg90vW5WA9HIcCKkpVB25P6TGOMFZD8pP/7mf8eU3QbYMRFwT4y8qpz
uALi8UINq8R4ESDstIMPWxVkP00j7sKCc7vHCqAK0EaMgi9OXn2Crz4UBxbc/isp
L2wfgB/mZF4E5A1WC7uF9Z8v3vuT22j2cPktGK9QJhBXq7fQShCNIwhNwiaLihLR
dQF9LFM3qIKMwlklNjwKyrp4LdIksHgtk7fX5/TC7ipdnWCDcizn3X1B0aOXmnkl
+lCX0uWDe24zwNLJ+3vWRVvf0B6S3UAnMoQoApGlVTqITePLlVRkIZTMzJ2Q4mAU
qUk1yTGfbhLrEtT2c3ziqy72+KQ7W56UkHdy3Juet4Gpn/XWOYgZIdaA6DlQdn+C
m/HthL/KojgUNBwmqHp1d8LfsEAiFfi/v2mCfhzhk7qR20pFD7sR3NM/yJEdKsPQ
w4uUYZbZundfZ0BtcIbkaD64ZKndk12v7pD214X7+hUaQtKKBT1+WRjSkpOLiiYA
s10c43MzmRfoLqyaGIjWFfrAnELf2iDYSXOrnKfAoz8AU87c9HTopFTZZeQ0TFNp
qr8FrgKxQwHmKT9Ps4/Rc7CNeVA75+gSOIy9lEm46UG/oqqLpLXcwDOV433qm5fl
lMSowfbc9+beQLUYZG7D0z3Iixy/t4QX7ar+M+ee5fzLGBSbOQy6kcI5XKh2HG6l
ov77pE9F3Xe+avWH97kXS6U4SXqu8BXVGtX7KUn0hHIvMQtdoxX9JmN61moFdTuv
xaMZRJT4p2V5j1+1DFY5vjIpOn39QX+BTWeJkDXodGuicYUMHrmVaR2CwdPxjJuE
iBvcrz7Otw2u07HQgYFev8lbOHEKfY14jWiL0VWw51NkULQsbrOUZk0v9wyJx7aa
ji+I31DDRpxubkNeWDGowzt/06powjdU+hT/VmVFzelB35syRmQFeqQOAOAWcE5s
ZDiQKhfZce6PoNCLiQMdTSF0ZCdcry0Sv8xneN3JeOpw2j9Kkhq+8aBtISdettFz
TpJ6QIFibn7vD2cyoB9fWce3qQtESynVZR+XE9KAb7NofSwc7JdsnLb4KuByZT5w
5wsIuJ9wIYFeYnOpMCVVXeM0b8GYwz1U1JGNTt768vg3Jt8uwusOcF3+/TIINRyY
Y4YChcnDiN439jJIVPQTh2YE/VUpzm83itGbUTpqn8kHhsldUAQlDQddro0CkX6U
6u2e/I+QRJi/y2otAm3E7ZiRPo/mQ74y3s2gMxFZrwmY2L0e1Gi9a0C7qxwroPVf
iB6KYxgZW6oT9SQiTiOjdVpH71oKHb7PhBpLrDbf282Z0Vr/Fz5Lr+dP3icp8bul
+JVtGxWXuMABV5fZspd1sRVgmLcu7kgXQs6jaS6Tf71SIq/UTr5CwcW//G4etZMN
XlzD/qjan9Ogw7DJminhir47xMR37raUd/ewhN57V7SNm6mWnTz1Kn6DFX3mpCYk
dOPzl5wEIvwOZ0/8d25lSZo0TG9kOc9TCkbKlebEKKovA+SlsmlyAN/El+36tRi5
g3i54GbHw5PVIMk4PDXt1Fb1OlBXRLlNWbf9+ghRepAEu2i+2N0pQ+o/iOqgR1YJ
IHfRu3oY8+LkjdpKLeh88rR4BmCIlCdlIKp6NBcLYh56crf546SHvtlSKyDXFP6Y
ALoOyOg7DkCu7y57RNkCbl7WPsa4qi3Asqvv9R6gJssmcHcypJtYQHVTz7gU+5Tf
ZDM5PcU8XnjqtVdthbdaieITj4sUBwFThY+yaUdQIwJfx8YdbN0r7nFxcnhLJ6Xw
QG1R+zytXq3+RnXyzorjTvLdCy9e9s8ez0SgNwcss53q7LGMRTVSk/MDPie/ocNC
ITt35Wu+xg4q3nMXuT2nCpuTvZ2lu/2ixK9OhephRHuCZoS6vDzccuKOeZr/UWDy
YQDF6Vdp2DlpYYOeOu6cc6QP+mqdqjt5JK/wdGXOEoDZjSi3qLtR7uplysD/VgwJ
dmrDmS797r4Q9LMo/RhL9ZUmyl7e8hc/S1FbD53Vp8YmZgWDUIugmJGliybZiRDr
UWygYf5gyZFL4Aw0AzCdrZ7AMuf+PsFA/XabzF7QcFqMLJ5hX/f1dK60YTerd/fG
z3zzwp5mF2V5lK3fhc8e5owO7mDi55RTH3PMFzQNMQh9/za65VYumwanCkD7KlGu
8MdAN8k19TJhIdW0OvnW+gnwjCi5Yr+D7u7fcwgBipZ7HBKOo9NW3EDdxjJZPvc7
IYK+K+BX4iKCY+jUqtIsHEeZkweHpT1PeCVh/3tL2yMqfoz8AO/Iv4tRBftjPfTf
JVTrIGsHshj0koA7reosCW0pD5MYF5Yoqk22mA/y9TNeHvATPIhpCCoigX7dK8VN
0JE/2NUq5BaSPuZeIl/TGt9bTqenlu0kqaR+m6Yzxl52EgsZNtvWZNWk1aYLlyQy
K/UrGSjJf+sRCV21zbYyuVq3x0YVkeq05kOfqenBv05Co8htFETMiGqEXHzm8Cio
/QNiK8GQzGEUEDHxBc9Uz6L2sWcuilCRsTcvlLe5RrBV9+C1m1wSvLNLLdcMM/cP
qwzE35zsjjLUJwyiCqKqcdgJaQCMLEbgmAc3huDumsfX+FQG9HXcTt0ZAqK1LmwN
SHrRrlogksiMwsbL1mq+uhSuIHlUOJS7bDQXqItRNLyhU4X8p/qp7cSnJn6Ibff9
+KZIgtOWEVnvPgvctiQYcQTnEpHVyPHo7lYkSpZ13dhb4wlnRKj+OMI5HjwwQGrG
eMGGAklerZwiNTG6bYpHcgFGQ+OOpQeDjdXxlJndG6/Ec5VCU+ztTObA1ekCXGxB
RT0SFGQlH5PtQ10H5l4VklNpdXn3P3hlVY65/j3InSSZf6JwX9qg9WonE6MTgNd2
BOJG2OkJd6kU2iFBfbJKNE1xgzzjaQ53EV3t0UHJC+eEKm8X7f81rMSU9ZpHCjgE
iPIRqVrJRwsxgRJUkec8eRuu+NXMiVT4ZTe0Otpsp0KRuPseRwqpGrtuXpLO5uje
kFWaTlVR8vAD7lQMxG/Upt3Uvb7JSgR9VWeUyaqH5KPs/13Vbkh0p9sZ78ESy6Ww
ZjIg5rwtFUvrYiJP/kp3byff3MJjg58uB/Q+nSMw2Rto4eSPub+tTrlT1NGvXedQ
6dU1gnarzlO7JDhgwSPSDoGkGGcj4tNvD3xb72Ukb13KXWP7gkP/6/AKebYRBEqV
LeELnWCwdv/4TDV9vGUeaDAZBhKRAqk0SakQG/GWcCJBLINoVpW9vSGIlU+/0Vo7
9gp9NXMjwOttd/iw/Qb4Ukqw5rwLol7aRITSlOJsvTfpdxu4uB8RfBmKu7AtreAq
aX0yqifIFVhNbNYSKvLYgSEOEfJ0cxhDZaKJ5tHQzEXJ7JaZM6t65YhUtL4Y4n5G
1Yq6Oca/IbE+8Vp8kyZyBRvC1w9J2naOwljpxF/x/pj+uOAWGKZXgqo8fqFs8vVF
mihgPlu1Dtjbdb4Osj4odpJ6ovqZjfnv0M8bF5GoV7uhizojjSMXEw7f1i67bz5t
iQpVl3MqdUKnRtW90sQ7GIgM/jmeUXDchCEswvm9nmvXU2rYn6rWIwm9iOcW+MiQ
euhJuXX3z8kUij7nmbdbr7d9bHUB87nZkZsZY9+e/NCsPJUW8oug6Ahxq8bUMBb2
J5mzcPCxvpdJkbCYAavO3wkHzvwoCaq+EX29mSGGlGq87o8LZsC+rtRgdrNe18Ro
ohC/r+K5bHkIaOiy2WPeMgKeDEMS1HvaKMgPATJFRS7nUpJUl+4zJsAJpxionusJ
T9AMRpKymZhuLHwNV5ntuuFLqvY37Ge5StjTvfZu4nr5vaN9pbgBLQ2CLQCrWJmt
8tmynnZzSYIE4P762ksRxzzp31u8TvPFlyrzfht+EzXMhur5IT2NgYiS2hkvUb1b
eBAX14v2IcGXgv6bF4oz/0+40W3rMFWWE4yeesqETqS+J97nV+wN1dyM+7JS4+tf
vLv4RGAvfNIONhrAzibiCrpfnmyyjPNZaGTaKxE/8neplmdjyCBdFpwblhuonyNo
V0WFxMF4sm2okPVQIwXLwAsrzUVulCy946VAKdvjwVMc76xQXHRNdOJbcUF6kggP
kt2giPBO467MJCdOsrmsST+ekcqKuweYkR+U9CwHGQxd5ihH5HfM8wVSqdzno8Ut
2Il8goOdstvtCuV2cJ2ghrfTSsffOa2TX4orlkMSQi4PVazAtN7VkomMXQdWq7ml
+tCmyPrvryf0quBICLEGyPme0gWdD08SIREnmp9MHfWY7+aLeiKg+5E9otTfaEW+
G4F98U/7uslNXYwOanBhD8Kq1XBCI3FK0WZ7LgSS06qgR/2QEv9hOdqzO8a+gOfS
nPVclnEJJNFKciuFh1eo4XnvzN/xQvzFyJz6S9hCxoMf+nfdKgv5SG8CGkeYtDc0
ODr3hcSn6ZyH+nQo8VN63r/vYhJllgw2NLGOJ4tRs62GnDtZqet+5sPM5Z6psV2k
mAAfSKSJTGeL3KH1uGEIWuWEHyFwJgeq5iXLF76xXVB2UynQUNig3nC5PPJMVuV5
QpcO8FuF2lKJOoOEyAeEJFJFv5Ess47bOH9C5SfpyfgY5dhX4Ue45JWNX4o1f+4h
2T/uRzuXWd4d+U4Q4IqiNBuBDwQWFNtpcolAbh5wYJZPzboSs9fqSE4psteQCHot
1KM224LrCf+yOrw5p4igGeid+IONTVr4wAt+1Kc49hLub/ciqs51L8376f+/AMvR
cJzL1jeGgsq5d/WjWlSCcJIXdd+DEJafcgaCRpoJrgM/Cr5dXpF17x9684lEQKAx
LAdMQeNLDS1sHNt1eHgKQUHypcsR4w29N5HGpXK27st0sIvJ8tmJZBbgZ2iO6HP0
cRM/VOHqKmjWU1XhWlYViO/sFA77qIMKAjacytU82T57u9CbnEEpfgyQ65V7MJAK
ILhfgSAiIbEP/eV/sL3GQsXu6xTJ7/P7CcjtbMpNaBgm6SZwbsOcopKmzY3VhvKX
+SDfpYm6t5i0AwldrXlZYnhJB9NyRUE7tUtXYRBeqBAFp5Z9IxmGj3o2ucj+88ko
9Spk8lb1IoON2eemXty7Cg43wyXe/eftPIDTBgHITQxABdJ/XLSKSbdjAyTHzDyn
Q873laQ8w42w43gXhBbSStoy22HiAzpDoNo5UnWWKXLsSNuBAUXlpHYt4v1AJj3z
SoqvoBxcNXZsCoRQLuLG2V9By++f7MEDOCfIT+eJ2rT4tWgVblfOjxOgHctsOoe4
6wHBOkhYPS8M0mdK+nfNmOXB1/FlmtpWg1iKXqlzmQwSXE/THobQUnA7k//66BFo
UqzuvlfnyrWVOalMdXodSvPopQeNoLeXCHqqoiGqP3bQybioTL+9EEnxi50C8YjV
9FS/FQuJHHmk1e+FuQk/9TEPnB5VwKArgkptcn2X1+wBt1e/7y8j3YIxgHnAeN+y
FqryRlBQrT/7nGqg50YoS8WDPWDrAYSaPthZ/8E5luKzdAjmjj9hrilEvdbJwIqr
xHpwD1KCcbfCDmUeOiN/sVEGJsWhrnvxgS7yKDAF44NRopB8m7ElCZyQKi/G7b1k
MSH58loDlj03W1GIr7NSe0DJNN7/dYw8ZCWgb9iewLQPzo+2OUiXTzd/InZByO/O
S3vxGUIbxQNPFQIh8VInkqBdyg/tv9qLsfwhnevE7f78QpdTXEPgS2xtdr5/btWs
N0PEzhB5BRlDL59YD3VEDxlPvwzdNrdnlxUzOXhX96JW3EDtxRWBgoYOVm85TM6f
QbAxSO0v6qqh6H00iQjeNKG8sd7vrWBLofZXpkU9edLXj5Lj7v3/eWoCbyGUHY0d
GNXOVQiQfnC+4V+blyDYGFPlVi570GAPIRNd0VIkmbZM8exNTWHCF5n3nXoC97IY
B1Q0itls5gVFzMa+3lmTBoxvPq1FVVNbvGFY77upVzrE9RdgY9S0AMCgXrjclT6c
bI9vg8S/z8I51TotMbjbsY8IxXzkeH1MrAJJoKul/+y/9VfC97gB4kgAmT5t7ts3
bs+uhIIebrQYE1AkrALDjCl3pxyO4cV+ouomuGLvQU1i4mIxE9iWYkJnZDc9cGJ/
/J//4wuWMcPeGXbRq9sJt2BpKk6WSPAQaKJcHWKKFiEaz+ngeKyQRdkI6geMhPGk
hZNg2UTt3wPdiHQY0o7NgDTlTRdl5kMs4ICjQpN4U4DTpXg9ByHiHEGLWVtjHWxU
6aWBVPBEFOWHaHD56TgSK66S4wWRqzOQ04+YdHHJhWpAptO3hVLRFeIl29myT2x+
lIMi+NlnNgMdIamc8lf1FuVMHXckYLpC8HAMSkoPUyvPBLnmKMlhrflDQebIzQfK
94Er4O1xjYkf+vtwfNgCh4a9aGBDhBDIbkrRNkeLT+6hexB7MKTZRvUzcRuZ9ZHJ
HLpCWQESbt2A7+RNRuR/pxr0Q7+0fhZgaHRvHY3o0X97W7CZSJj3AevBdacpY9+r
GO39tw02wzc5biEN+cpvCof2BopjwcsoxtCg3Il3NKy89E8PKj3fz7cmFfNu6Vpu
tyuMPsRksQdSElz1zazaqUxctYzROyyOq3bL06pHtP7J8F1GSJ7U8Q4z4YGA+i+M
TZKWs6QZJLOujNUN8hnxvjqC6vq9BIhYvDmUE5Wz/A5UAJffNNptiR3xsQ3kwiWu
7MyhnFhzuRytcfFGTqv4YbXNJ++AsoGB3kqgS0uds4UlgFeYgZLDt2qldTUJtdfV
KgtLtD3xIGL+agqnnOr6Y7rCvwVEYTc+dAa9FEoCz4nO4yZdMpNC1RBXq6iEEDhH
KK29O/SJFkgWpbANygxH7GpjcUs9+o5d/I/yOqpEVbnLZrz9eEUn2HXVIVmDHTMr
K7i82HJ4qwcTku4iOyB6yUp1XZaacY26z+3NrIfSd5qhE8OaeAStxhNnSpXMnmSl
lOy6mWRPJBscf6sY+kwxy9laAoUwEHJJq9bx0QqjYFd6cos/IpXqoZvx5g3qEF0z
6q6dN51o2gZbBiOJa1vECwal/r0Jm9XWbCpg+dFU5czVhOzdL/NvBrTb6W+WUcXi
ufoi2x4Sx5s2yO9g5fAeyKX3fru3Pz8U/f2wRdPndcIVr2FU//lj4nQ4B3t8fZ7R
+W89Bssywu8x0OieIu2Z5nJJcw5Ngkb3ppML9ve+qG4RcwkjgOJMAb8Rc7Diz9F5
5SK3SvNuGcdnTOGYzvY+aY9lnMBq5MbeFu6Gmb1KpWVp4FNp9D2Aqp9DAZ2QBu5z
OAhU7v0dTGNm4AceQieflEegpjRCsLP6iSxR8YT8SebQNqcj0uHx9qRwmSx183r4
nrABRMkNI4wzSIi2OCu7mtZHVUtelsmXkIKahyg61e4NyNibVVJosU8xM7oqXTs4
TgI4qRa3O+XI04RV4ilZK5AkIBBDfrxI/fiXkPU/YT3/wzPDThGf8G2MPvkUPVUJ
Yzrza6qVs509gT6SlT/MihULI5ThQlMY9RgcHGDHejnR87vv/1zQZBUv9ig6ylf4
N6ZPbhnL9yjMNyPlHpDAHrvIPqsVV9XnepwLSoyijmMXr/WyMbFovEyf2zbeakEG
vY23mAq9HACMU4WtyyXVoCN9RXu552N+4vVcZNuWmitK+B5dJU13Afmx5IRF4zGm
LzYX51KBGvm1tYeZ71RiGi2SH47YjwaGLhdxr9XWmTo6wsMLxzAZjaJEO3Ek/AqE
S06vTRQT0uQRi3d67vog+OFN8D9Wws88vW+O2M5MzzJDEdQW5VShggfsro/o+xhD
p8PegNQfW5DBC0M67ShEum8UICSsDFF47V/ovCgEK4sN8JIUViYOueHaJiNH40o0
YmKIg1mfk5VzQQWXYsgUBKI8fRWCwBaBy3cswauE4041vBV/IjSdaqPmwsBTXPj/
crE7ioptWLdi9XNqT+f/9NCC7Ik8+iwXOtR8iuolSweQUYt8QNSlq91s5MZCjh/y
DLBUj+tjHdp9CNVq2lAWgewzznj+yWiclWOyVobwv/Z2UvFXKRC+ObVhQdlEgRWp
qurNqgOwx/Dz8dCRykWD5irZ4V1jI2PEFxLPZdDF40VqpcP0/0/2TY6C0pN+QGi6
182RfdruVfPC9i9C6X6Lx2KFwyeV3TipBgf0zqnXHdEyad5YXRh5x/PSelEe3xBe
3G5uCJ0cW0k9UEVhBd1hHArROauZhyihQJYn0xKda0qZxdsRGG3AXhuiGJ0P3G0/
PBFRHnsQAcTwd/lf5nEt33LgPSSD9VRTRIfNMpvMBTDU6aCvSPKTEc0Y89NL6lT2
DD0IGAdTxvW5vHxPNyzSplgBdJtKXVGjqm3SOExYTyne+nYmYS6p3UDFGgLc2fJr
Ml3LqmX+juXA6pqzWRFmc5a5LN10Xk/NZou/tN6hDXCdcapd/jY+vIv4bxyEcHNS
8jNHrkcGkdojxyGubf4D8rm5SyWdjGvKSLQsLHYRCRjb742HoPRXlS+/Tdq9OrXR
t0o77XYfvo7bgQLrbQNx3YkQoGI5s0DgNRyxGN8+R/Y+yeszU87ZLLFWcImbqqep
iMkC7INStSUYesBpLo5Qf8NMQHi8I/2JdSIFuvbj00NF738CB1Pz0ix5b/xmCEpO
JXKVYuBvpJLAOhWhiWf8XIEj5zE2apCrVPnddSzAYtwhPhqg6J3t/IroDh4JOBzy
dKe7rmwKbUPKshr2CSBEQ+mgB9BeNb/jC1LnCkLIjRVXlLuLvT5CfKP5w5OWrhu/
1+VcQgmL0GwehnMtCqCCAcDeyb1cqYiQMPpN8NfQ9mkNH7lz+cpOIUBQe5jWlGY4
0HK6mYJaM2YM0HsQeaUcHzMi8TDFQ/MfMwdWrCh5Td5IFwxtNBFzBLKUrQdoGgJH
u72pIb1UDktlL6NOM+8XdEHooxst0epZKJV/kX8577T2n66w/UpqurkjUqMqOhGI
z+MbwZjEx+pbThJH80SzAe2vWiBvTJikv+kKTjp/Xma9ppRJG/LWusjHhv5qtymk
S5JCaDOuOAmbtoXZEhoo89iLMM9LEWjzxxzDdlLIMhJ3jFoUXNizJ+8aLrEsXlW7
C348T9XtigfNsIh8YfFoV2758ifylDZHc4i4KJYgxk1dCEVqodvDwhKeJt196WcY
SQgGxUT6cIxkjoj0PqmVWmO9kApIgEnk4qWfnyTW5+2Jygb4zRVlEK4mBkkrnriW
9VWlOT93LvRZ2GZMoDn44LGGrZocl4TFevyY+QgW86rbRG5DAXWuAzA5vnZSf+nr
xMdMaf4IDocCKgDcQfrYs49yJr5cZU7nQCLWQr6WQmaAxDJhgBH3oaNyZXrizka9
5I0uTAueTN9a5ARa7z1If/knN4tX/W1CgBFWM4lpZ6wMteOMoVsMmB1/tAlg1b/3
67X4yp4r8lQZiRKUGGCqFw9CLd+IlLWtAjqmA2pLaVJYfJMBhXjhLUfb8Vx8HoRt
XahDGO4EW6kwuQOA5zPKat8b8MjuV2RVrxL3y1CDlfGqvKM+JCjBPV918yXGCqRk
MZ4DiapkKwl+sZ+fC8RI//lbrEHZxN7Ti3THS/Bd6WwzyFJrof6Ru0F8KtgOxS/h
0BpO35AqFl0ki3IJyRQUUJ2wyJZVVj6BgozrKvvowoskduWaORrKkXzrh5EVzFAW
/FLt0An6A5bfwBodz/ybSRooH6VXPySvntaYf5Kd3r7vALn00LRA9jY6IRCSSb/3
EMXuOEmenoIn8aBIDIFafXL5EZYY4Kow2JPelgkLSr+2xa0rhgxZEksFZbeNCzmo
987hOdA7b1m3GJnMTM2/mMitqF+FVrkHOF9ilDVrl7qjqHpONhxQVZlhcPmvmVtm
uvtHJOUNMNAx5zMailA6eN2M8bwZiPmPmDGMF+sjFmmk1h28QwBqcoXLGmZN357+
30009QI1u0mFloalY1GfPNijZEUi8wccrD3DFwk6WygVa1M5dsb6z0T33r71c6al
0t8BmX3jNNpG7IREAxQGuvJav5c692mHwPVkrTwj0xNyJHNHJisXapA7lzrA1VKh
1qeB6AzFUntYB2c6FCWk4MDyAw+IxT0ONHxXwNCVvcNijLCjNM1PHiuYIcwAngTH
p6eX2ejrtvOJSjz6K8EPKERfMkqYR7XkRBwgAqhgE1/2/PM3ZnHLR4OIAOOlKjb+
vHxwfavwuRitb7jOaItzEzAqmyBHgBs1/Gtr5hxFy50P2D0Vi3GqKU2ny3nwOIaF
Ox8Rdgdgy5inpx73hXgDuU8hLOUdtGAijUnIASL0iZKHfttpBBJcZvqARdcCIW6Y
9CtShPpZw0LMGUHOHb5t0dyayK2/FkJR1mr7kkfU51OLVxEIa7+w3JLNRdhTcQZy
YB0k3ZZv9E36FG56dZVr0XGk7WA9g399X0A/JvmlE+n8dO0DpJr9gAsln8AhJGRu
UncGSyIFKEgee+suhtRcVLrv1udtZ23+Bit1Z4ACdwd8QrP1OTCXFgifi9PPWdqb
gJAgHusmhAgMgDxHFy8fIkVQIGNBP0sfVUp1D5UowoOuZgPHUcTT/9SL/x8Ancg5
mRgjvcMXlu+vLzKqjyvXF7dVnQUleHE/owI2oGgpMJmmLxgLeN6U1P0lNxRKamWx
BHGa0WAwfJIlLHRqPyt0yZ+4d8iMDXWBKqsYoz73wLcXrwUTBpfH/HdJlpTOW3tk
VHGhprg7iYPz8YzWk6A8Gf2p+xT/Il3dK7VgPV9waOVLpOERKvrZEtmY4RSRmzaK
SNGEVeJ3CBDQ5VnrqRyTrFqDOjZIg+QSs5qlBQH/UjvCoxODfHSwlig4/7wiQfKv
wwZ8GR5C0A3Z1FC9sqUPflMHsT54HYLcb68mc2a73/yZvsJcRXi/DgqeU1fty+NG
U7EyGhkg4tleCLdYYbZokoNDs65nrE360lMhWVIvQhxZYeBGxa15MJV04Uj4SbgB
/W/lGlvPS9IuRSM9vCLyNr8chf9earNTkfVKuno4WQ9KUbqDDedTPfUtkf6An91M
5osTpvOKQQVeSSTSlRfgwYo+dVvvtSsEGfyI4Uc4ydwoCLyJ7Reu+1qtWFapy24p
SZcTkqqveI4sZQAyRDQfuF0iCEQ/iawEbcMjDT6C3HS794UbEsQXS611EoEb7GLl
nilCcqx+/At1dYxEXLN1uQzAzFYODPZXDnpq9P11US39pbhijCh2tU500zjaQE4t
71Jyl1AM/cRG70PqJWLQZTrJpnp11GNf7YuuMzl/mhqgAHVNGlaBDLLVdI6cqqYa
kYrv1vraLVYB+MAQdZwroc6kww8XAinXrpfj97UhWqqS9z9wS1yN2y7OdyXPSoM9
8s5diLoMVqbKWaTMUj+IHMmEIKgF06gL+WerpOLWw6wCNt/5t2/Gcg5bpYwJrvZu
09e4vLH2NVoNphaTs1qY5mdx/vMACEuntNRzkImjckHRTlvfaPlFWfq5rhdzAYzC
XpzW0UoRGmfbpgQdtC1ulyvopxBUEIEyAKaR0LRLbtZfu9j6ziwrZG7DC6xDgwZ3
QdINV3KSD6GDV0TFSzIn1RuGQfntluD3Gs/IUjLSrjLBx4IlYcLsUxwJ07qhqeVR
MXTIRKLLX7lemnRHEkFYWRBIqguyMhXF/57k47SqJHtA44CG5sY3SxGaE8GXR0a2
laokxzb3N8dhkp1/lN3KLlg0Mnh7IkP+w68lHoWIG+2NQHJMX7hhLPv5I+6yHpIf
aDb2ZnlHbhadBLr8CQzJtQ6I53si+Q8wKfia758Y7g+FGuRtMDx8QDYXL/bkMLPQ
zyoo6552kJb38tCOLYnirx3cfg2rF4GlyRWFf+YUoOR/CP6bSyVebI5K92YEPvL1
xt+/+2GsHo7yQa0u0NSe4gbTWq1GDCrihFQ6tJpiwKhQS0rb8ZUue48a3PI7AVzS
dtFQsaHLXQtkkLowJhvmrzo9MDlgT5/qtrAqbQ1xV26s7e6/iy6M/2WuFkO/nTyR
0+wxL9tbx82nTsY4kwvWPxrURKoBkprOjJ9/hht0nHJdhm4IiA5OGxSz1XBEIiDp
xeX3cyU5lJF3XWCsOKPJsFQYVZr0PGkNvu9n2shNk2tJaYGx3e/8f/qh5fciYqtA
dOmZxVrIvSsFykfPNh7l2Rlh4s2H56/1MWPIAqa7b+3S9Mji8XFnR7it0cjCuCsP
8MThbsOn4kDCe0OtP1KAL86ZrHRi7ebf2aExOptKiuvcQYlQG7Y45BaY0kbT7OCG
A7D4NOqdD0GwlxwEZUFpqWHSvVR8hJWAfmzgnlb/zuKBLDHy+ZLhpPRZ5NYYZJve
6aLz3GAYrzFqNcwHDeMF7Y2XWg0ksKShSghelJQCvxmFQwPwRHk493lY5TxHV+uH
hJ/cnIpNcXvlAQ1eACivbhZ6JPBMiZfI+HgUbxgM8onSrWWxskde+AQmNMvTth0b
ZKUSNPu5QyDr7obMWmMx0qhAPSo3rmbNDyU31Q1YfSiS5a+4mTBAgdIrC7GVR29v
Ne5xhhx0ZYTofHy39Z+lu6plZQSMZCDsWOXoaqwYw3g2KBEca59naEAAGysd/T1f
5+A3qLL2ypX+3ISI57EbMUfw9T9OXSzxm7kZwPPJ+BPfje+idgrerN0zXSMQiDiQ
6yAOORVmUTU8fWlYwd1p+HTgraSF157ejBgHMjT6mtvQOA0Y7U87434kuOr8lyp7
+jQUNkF4VkgGgmGJwUTMnKN0lFXYq7MBoARidAk4JPqDtYJta11uKpi3C7q7yZsf
RLb/jyiGy2w0Rhm2aRHEzzyOhcFqjf7TviBmG+DBGTHv/90hNiP9/ji/s1KdhF6G
Uu5YJrOkem0/FTFN8CHq1mXYUppxkwiHtDRITDHwZgp/VQVTspmzLV85UZFmGAlE
pZSf8WByPHTXRy6bE06KnQQd54dQfRI6lW6I5ys8IvHnzA2TZyF2WAQhHUWeQVjo
UVSWvxUYC31tmHv1U9UyINRZg4hTgGqjpJtNsUqxw0FtWGI7UCCPpw0iesVeNKV6
yg7mKaK/wTvcXTiNwjfVibTTa9nCsK9GloR2coPBqiWhPCMyxSe7KvSV765/IVEH
Y++LkcNtsryVzmUh4RMEbNAUEdUUC9xq0vuTgJQ1h8pTywT5Lo6g4VSes9+x11OZ
IjEDX+N8If5Zb1AIGZsa17jZVnq921hkHgAi+wMSzWdzzigNoS7OlFBUXD79SZyL
S0FP3CY8LR0pJoUCzs2b36Vc9WZotqqSyuqlO6/0dzMV3fx9jXUz17pbrk0rJTiq
fYLBsk/spvU1st43FoPjeZ2KqDR2nk+DQJg4fT2yaoYF1Jbr45OoaBaEEfdOheRS
103LSoXvFAeGOXuyf5haxD5zyuXdnWfmGVipK3PFY0EWhtvWufj3zCN3t41CpJD9
1w20HB15mgOWKCKq0buw2Dx/3o23h1RKG2NnGnl4IO7/h+bzazFpYc7kP/HWq+o/
Mx+qTQiN2QKbFDpCYhd95OgW1zkCS/AeQlE6WRqgCUtywKhOnLgUD/rLDVeCa+T+
J09esZYiSbzNfqohkw1O8v5lf7UAU3Z2aAdBKdpmtzcPRn8DWJe2Fbl3RKE8hvYM
E+dUozl7RQQTN6MoVBBMkG/VO5PZsqUQiZKAbAMHpuQ8gOdI6ohqC93DJvBQ9krb
gGX5MPERh0zQJvhtE21b4n6JsDtl189slrtirTWbrDFdKeYWMl2ZVkqxhDV/val4
w0HSBIf+RW3s61oHBrLuL48gRaO6yZ/7rd9wLOzqJEK0gjjGMgbzVOjBrzTuDvko
0fBg1KPzp+Ki6vMPqFZqvDzTShArEdyuyG0OtEZatVVZGDHzEpKIRyhp1eT8PxxL
nfnnMgKO9I8eHIgC1dm7JVNaEq37Lnp0oheZvgq6pnlUe5ApR/bRATW9ZDJYylvI
Bbd608XZccOSpyQgIj4083zpmEpYaMumvVbhRGMeMdw8oDL06DxuWDyXqQxQkYFJ
50UvEH3YJiiU2wT4gsoxBgYTXKv6kABu7lCddA9A1Xg6sW3odWGj7onHfIjAXaSh
ycCWUFvCfmtJoSnGGRxG5G1VunmtYWpxU8jZIHawxTw8whX8JWxK9XtkEsVPY85g
STBRmthCkPlAUp5Lyx3L0Iyx8MbcrLUKg1jI0JKgZs48dlaBSBhiqeGSFlDfDiUM
J8TUpO0yynA5Fjt4RZyH6Ef81WJLaJTCQHxkgu7lYt9IfrIRcdb/lwb2i6LQzuOX
jhXYRfvossWRyF1nPFZki5o1lj2hBt62qrtcWia4tA0Ab3+bLjYAuvjzs1ucs55Z
6T6IO1PmVQ/DcMQpYzEvEBOp4uf69qeBPL4gpohNxfelZya3WGlIojIeM5gFXJyF
1s/q3y1K5XdsLyW111Yi6I7yFmmEjNJfZo7HYOxhPp2NIPEdK1teno3Dr9edu131
FbJxrCG+UsEjGfVYC9BNosQjXepktDpwYJ9I0etER1LK1lwnzMzJ3Gt5uTye6qIy
mpD+H9G/OJn0jIzdG3TfNSQYl5VDR+aWSdfEjTeBp92zkmMx8Mc2Q7yXUrBYW3JP
tk0OOOob1wjINEOjvhLqRKOw2smLSkEOuBEmN7ewAWTmEm/4ucW+ISKimtcogdip
V+aN1bRjz8Gkmydq+Onl2EmuQPr4j6NjFLuh8OzDA41KVEuKxPwcJpRI5MZOpI8t
1uMP9qdAwfjXXB+KOUcYtAKupdmZdeiECVXhH1LXjp7+/SNXnodN9z2X8bGXPA88
VA38zKwTIkzfrY/owfl+uqElciRS3bLuTrKdK4k6Y5d5dWaa584vlM3TrrL6FXsT
X6FzjWR7MV1Kfi+WfBgjAY+KGBTTUm8DjbdJbW4EHTcPSsEjpMjK3wYi9nZYBiWd
cse9kJhW8S16Z2gRsH0gFT54FqRZc79C1ByXys+6VRpVE2dLWIdZqrZKnRByKP+K
w/lAaXkXZ9kJ+bG479F8KabHDioibp7iZ7+lLeg13ZdndcSZOOe4i9xjYPTjbxpw
eB7Z1CXEHGoLfeecEPN+raSUD+yBfXf9fn48lMc3S7vsWtSmCtB3KWrDwUR9HvCX
FnADpfthnSN5XAaIptvtVMBHe8cSNqsieN91YrWtjilz5QxLaVip6xWW9CTO0OTs
Yfhiild3a/ZZ8FUyTnFPtT3nQRoT1u+1Vo28cpAyKn9KydN8Y0uiK+Pqnbfd4228
sq+/vx8fNM1s+fLzmG7PS9qVb88k6uShPRCFIIs4smP5na6u/KHT3aYnH9opXsbQ
MWEcYTN75I5Koyd9WwsjmwQhkBjDdV26WvkyrY+K+2y/os9JeJw5ZUaCmX9YC92/
acMR/Ab4BWgomcvI2ZPvsAiOASL+H1XfQeh4l7EkzJWfl6dfmUGzI2rm1YMBsRXl
ZOPkMW6OBJFxccu3i/RO/W9KjfLQKgPiHrrqtcYwI7JNxJAsLFHrcB8aQ91hSOsP
WAjmCHPvjp9R99wjfmY2Sc0gfa6NwLL1bnufI/juoPsUjAlEvvyW6NZn0CfQPocy
7Y+yoQbK0d0I7GHf39Ng7zU8OreYpVC3uBT5Rzh8SqGN8zZO2Lvu1Jl7W1bVElnY
9Wm6ogY480HkjI5Xee9QODncFwy8iWkV3Iq97Vm1M1PAvsI0ziAwTfubgVPq2T1z
ujseVTRRkCtrX1j8Qx3iYKJ8TcpglHJW0wohMTUVEIIWX+CQscxLvQZFdZX4k9zL
jy9pT5wz1ZaqMFy+YJ/zYC0OZQkEgD7K8pGyBBFE854peg0mc5XJL6DGPSgva4mx
hvUQpHNn5S95YPpA2vaIOQoHPb0ttZRnSG1kW5qOYO4+h7IA9+0NMUQzzHqg19QF
hHgri+gb+3Ijp2xxNDVlBdlAQB0mlv6BnN3SfzphN9+ZxzJqgyQb40Ywix7oR2Hu
VU8JjJCgMfAhggqdNl0svENeTacXLnEzVbRJ1kiyrZeM2x+kMWrBT4qP7kXJyWpr
nOAG4zQJ46ALrVmNfyuEcuyLUDwA7PAbY3VMWmQDdxDE8dALPWeHY5/8dcc4kSHE
v1s0kZ2rYarfco4VRooQ6IkQ9m2leNLJpfEE+77V+btPGAoRq6Z9Ax5vLtAHoJId
cUlCIV//LlMYfzQmdrAlld504apt/J1x41MsS3CJ/hMM7bwKmym1IYmAqInPj+FI
oyOuy5I8hwCy6SEkxZa9AQO90vWPuADBD1p+uLXbz61wKhWWT43NrwBcQ67+1EgT
OCYvE6MoReoAApujYhX0hs7dJYnBCed88CBIaIAuJRUMpRs0I6Z8vmezLE4CHchg
Ll0Fung/htZoAVjQukeopmv1QU+0msUbE0i/9SVaeKlzVMT2gIPj5zHeM+l34Tv+
hZTQrwEX3/2n7rlApsFV+Oblzi32v0kq1O023opsrL2tk3BI6zXQQh4/yFcd3Vuz
MbXGga7ftIK48d1uS5oGmFXb9NMzlx43EZxVjnXhyEt7lC04yBU8+BOgsMH6f3b7
CEaLsp7yM7HLYanP9MfyrOzEBrzUZXbTgiU5IF4DSjM8JwgSJbDTmz1mgDQWwHLf
SHFpdPIGScRHzHkT5WO1sDQk5/3rXiX+ja8WdyI1fKtQLU5fHuAagOixecri20ZG
b7wg4rEL4FOhzY1PsBewe3JIIQroFLSYPN8Pvkz81y3myPW+HiDyR02G5OUR/LDN
WQ5O8yQcJhKKVEfohIL2Rm9+Fg0DVSPa/rqiuyVS1krrzD4YMPqdszf/0zuST6FH
iUl6O7+pJobLAO2mZRj3eSXE7qQJMPZJazgndZErdVPtqm8jKDS1laWbvgZBwPa7
q2oDRkQEQM8rMzQBdJZPwhtc2QifMttb4Ahw166MObBPpkh1cgQhi2Bf2VoZKP0k
zUkQ+DB9S2OfMd3Fa7p6WS/iP/fMOHNBMn7Vj2ZCKl/niTAIEsmoWUOeYqZsjNBS
Gh9XNtK28eRpfzb6WX790Q8i8Cek/ysEkDzUkQEcpWj183DTYRsRYXOSc7oLKTPt
uM9K/VxsEz0Ivmcc7i4yyP5+Dg1EEwWwy0CtUOHRHL057TuKhvpD/ENucwEkX+WF
axZ+T1eVb4QfMVreLRHKrueiKsfJcquy2Ee34jWKrQCveBLBgTS82WZMEa5v5/uj
LAYgCcuz00hDuYOJYKmpfVhxN/bTOYymr6T5N8Hj12DUGGsqTaoa8D68IjTXtuOh
0uvHwmiefRsvVO+fBQwoth7H+FRk/Ev7UaYqZw/ojIRmJxEJ6CzYbLZdqQMyOJ1s
3qfqJcWjpp5mmOvmAPph3zKSTYNvcNRJ3xuL0+witPTn9ApYrGQZcOBy2QYoWWuZ
vWkez2Ucw4ZNs8cRGzu8Uy6K0zpFi2qKPRmFmys6LohqVhViXdxQ3UolnfF2VUEu
mKY42SjGMvZwtqYh0EWfdN6OX76yrDHoGfxjtLG/BD+Hs6PgOAod6LD07s9pP4rv
VtRwd+ITw01SC391fbbY8El6pp8OUDiTOr63gL8QiMGAn26vl+NX96YUhcBL5JUs
ZQ4VoWwRMBEDk8k7wxf0UiU1sDqDty3hLa905LdS+c4xG26e3C87kvTgvR7K0xTR
++TZu70RrGiUledQLayhVr88GXJQFkb4897ByYnp+bkqRG3wTUY2CNdD/LMrRyqK
0nUmg/AJnMZo42mzGqTy1/DyjVGkeiN/PkE3B97+08Q3fbS8GpBuw/dgckELYwwZ
trtGVXzjPMNIlNyVDMi6kT8+lgeR+kX6AD6aMTXl84xA7pqkqAzWqN5rx5Zkxm2Y
//qUTWMGRJTsRaOVLvqTInLNqaNFzT04kLCjFqoKahBnZy0D242pcCZUb/Ul90C3
tgz5wAaa+Qk3TwHn6RJPfkhQTSf+J7qQg60OIA8CD2Xz7fFIxlvwtQMS3U21zzmM
MAVfySdtB+n1SWS4+JI8IpBoDzsI6uH29pwZKrtLNDmGM6Yv+u4Pa+eg6fdjH2KS
RjCQYt11Hds8RFF9qG9u2iWw6vn8sq0O8RoGaxc4CoDj44uiFqncvS2rhfkW4v7R
6u/QMUKO+K8xXe+I84zcnWzLPw1JQFEwX6xP30uTFi6CtttXVkIyhz7Rd9D4uh0t
ntWn4gw6H06zfoyZtQNA285OrALfsYbA9c759T5+vHHFAOj1GYPUFKpJ/MgUD//p
222Bx/ogttrgCmAgjcffwQdN5zVw/LaZmVKKnmk+Y7+TwR6Wn5KS6pqrWciKizqh
XpGX0VugiuRadSt/jPKyPqRAXCRiHnqPHyTyIuo/yntTKlx3Ic0Q6YYfimI6U0eh
lpJmwKIr7c0JLDjmxhgbVaZVkllzhf9Y++KS34RAYbFXLrWBcgC6BPt2uzj+LKjy
pFOULJVQN5e6zc8zewlBzdw4OQnnPeTLwDyRTG6qzITnPfnzwRO/9qMlZAR4f01w
pGoQu/jvAxKMS8frAPuNCHGFXiFRrE8ojcF5zrF2Y1RTnkRQSsBaKunY17SW2dV2
uLh3Qz5+N9yR1Ze/B/cTuFwrjm9eOhwCjEyfyMmPFWx4rj+S/zqKk1zMAraAE7RD
mHiQ680ZDZkzPavqTQNIi76QZr3/05e/Hdmw2TORa/8+AMl6hG6DSgcrXZVrIlo9
4DsTFgvZk0DlxW1xOU/wwcPHz1K6sXDxPnBPYiGkiTm4sj0sio8ikJT93BCNt/TZ
agq+7fnvO6GIb1qyc2ED+8NHGUZx7wHeKA4i0jWex4uYRI7SaaMJUe7c819vUfCv
Jy3BCbepUs5K6epmra3BGeSZKO2ajjsoTq2+6yKJNnNx8m8w7cMvd7NNiPQmvC8h
1edHcjogzphYwPe8vbqJQ+MPohzgvCNHqUuTwhOwIzP6zRL+4V+08pY4mV1ebsx1
z4wC23toEoWaJzo/U/efVHXul9IfVMdEpQZZnovPAsdqk3cEs0xpyblCtKkQhycA
s8R5vZneTNVBCQfO20tbfldIwU1+sZmjpiqNaDPotWCyhaax7uwGWs+2Iyjw7vSS
o0L0y8p6vu4d0afv/a+zVqXv/7ZnNx3b/2U257fJRsaTKxIQa0EY9bRFNMMxO7EJ
3sduvUm5BPyywiuTHDkL15vIvRCLO/ZJ45zMJWNnaGSx/JeIDlWopKgb1JO3Bavm
DAKbyTEgFm8cINeRAcw1dnFMfzKPQUbB3nBaPZzCN+tRJarIcGKDB6/a/g8lyThf
RtCJzBeNQqz4wMOolklEnFnykKRHNM0OBLXr72A1CiZOdmasUJpy0RrxG6iwcG1i
k9Z3djUwyrMxjCbGG0HJna3dMH2wz5XZ7Wo8fUG4lazetqVXwQSFC/Ii7MNV2H5R
cStCeOGX5h24lQpyFQmtH1f928lYeF6/XI3SP6uXTGdU0rnpaOTzeFIQHeGEGBJG
Prw5Ef0cM2IuOYmD25+gwvE5H7aPnudtWeT//DPjEl3GBokbHE5qz8JYXVoG1Dhn
YiBeZ+eEv11WIH5UQBcVFIOGr958tdnP8qFnp+gZed9ZF2HraoArZ7c/V9X1cDx0
7dfz+2+6E58aOaBXdAURojkE7BvA/9DHZE1jxWCDV6AB8tKoXogh6UUxfr96Ayih
1yRhh5/KoXE+R/sI06QuK7o1ltUzfx5qbLzvNFfuOFm5WLz08TfaZT7XTGJS6DBx
tTk7WXi5nYrnANr7QtgFeUUBlfTslqztNlsS0Nv5pMWTyrfQLvd0ngaL6DifSiNd
v5sB854KZKoyuPUhyp5eN5KLUhIhyYz6vPU9gHz+GNcIVau0ndavngLdtDuiuvuf
nY7yD8cLrTxiKd7y9RKK0tTNqCi+L70jl4eKHpZylF1xrIw22Ck7hxSIjnozvNwP
rMpacao6lykkM6gbCxhc24dQYooPNqtbhnX8RgK7t43dq/8ZA+1ClL5VF51NKsj/
ZbBoSQgqnqtqPX868tdIircDoIbButzv++R+In1p4qu69aEJKwp4LUS6qPt3cdQb
n+KIQbEMAip42CSB0eq4jKjek0VSp8s5QBqfTXsZBFLTAVS8VOmzWplxAjnVhPi7
LXRJO047rJMbeYFWxqlBeNEBu/hA8aczg1dp5VpdvCcrHXTrwfNczLZ6A1tMowvn
D2JUdPSPMGtmuFtd5xWFoctuj7myydx4FWi8+i9gvsEl9/jrP4KBoi+Cc1io6ifS
inomOeMvwGK2HAhfRDK5GrSRPo55YnA8t+YKzNQSEx/M5sfQPtiOm/SrFqCBBCGr
8IglNVUjMJyZO+/upGbG6l1w7L3WkAsKNv5rQ+/1ecrQxRkZjjDsxqV1hshosbJB
opd0ligtlV39jOKx9ob8Ovztksz9FuF+Z941042QCu7gisV9i+Om8GEwqyDuITeA
ys8ENcPM//6lnp4DQC1hC0FMLQH238VsM2j7v7jYTtUfjPmvT2nnP7YiOL+L6B2x
3E6758LG78QSHqCMHgxjEkfquRVBQg2IXFK/92Kh8dG6hXlN1Hl0ZiFbzYgrs8Pw
rVV16JGy3ef7H5Y86wkUgkKSjsVvuWWj4ZdXkuXkmyHUrxvQ2tUE2U1LPL9/DbNZ
BYvBSwyZly2B8KfGXBN+wJhBbF4E/dzjqP9r3+pSnlhRGSY+Fpb8hcKTJtQz0FIS
OVMpGIkSPos7WUwKP05tFFpYiCUFNPetALNvKjHFlIgLTCx4Cngg48cpmMUTotLV
98BtYLsIc+rUblNnjHPfMj7TcAyjySrLFbUDV2WgYYFVV6PifMTLoVnMaUJJ34F6
k0v8fiUTKPqLUKbNHo3k8QUWWaKGIRcrQcW2O7rmB0pY003dT9LXjJCdwtyhtFMP
qi5YlgW/f46VpBg28cv1swOBbFLT/T4zaYKXiwZtB/L2hNPhaW4OttXr7cFx2q2g
rEJQ8WcVKTbriFokwstOaFJFU2hCZVq3rMH90O8XQT6pFn1Aqp1ZyPTUJm6KY0VE
PxiMuN5xevoYdy8PYU6bayNlPwE77lnG2cQMq/JGfwfzuTJTT/eoE90AthGpjBYQ
KRL9+QcGdgz7ED1uFHCk5VziVTf+W1sCfslkCY5rNE6NP1k1a3uDBjz55//s+PJZ
QqDcSJ06jALs+qlvkErwPdIkM/b39jXXjtY5YuoUMGfX9j3GKzRSzvMwc5LNs+Gc
LatZSQ/LkNxDStVHZeWh3JxcAGPVn0q4GM0UIDuaeLXuyxC3Aul+ot5mvK1zXkvS
OF89WaEDElDNfCTM3IYATYN9dox6DFO0gluNVy3ZkNsGua5vV7SQOgJ5Smz2P9mk
QJ9yjNfmOO7x7HYCGfNkg8u2PagleWV1+luD6w1hFpALZHJv5h+KX0i3qE2Yd6OU
JG3hiMLdkeWbnpTzGiF85xq+i43J2eelwctwdln7yP1Jps0xr8qO4iEcq4oLlv44
4+ZlUkmrVAmGA5BfoeN5f0ueD+pp1iuHvnICK1uVSC6dz5UU8yDPqr84KssZca65
axmYR/hfHwE82HDaPzkHva3YSCUbuKZ40nHaD6WdP2PcOY+bYJxrw6Liw0zCDveX
9g3MS06zNlp5NQ4iu1GH1FU1qNEKDzNQhfEV5X2bfrdKr+PlXmhLHNwBrnbjFtb6
C8fdbR8kjBLi+Sbnh898PUbZcZL42UJe56hqafJFQv+N6kqIiFctXNeVIsazpUI2
5wodlMoQhWCcAHMKotLoNCKu/3PQgHsAK8gXsog/G02gWXwFTEoNivyaQaw2Nmjv
6MzcL3NKfmBHPuvTwDp/OqgESsxv00k7HCYG8FX/r3zwkPNFBE+7rhqwyxkFrzW9
dK4udNL7xE8sF99viigfgKrFDT8GeSPIy5mIetEfHVszG8W9nhpCeCmc04HZjzHf
KNZjPTLx8AD19NCtDPtSX90elj04GBoJIiRNWEfp+cvLaOboOox8WQ3x5KNEfBv5
l3sxJlChAyXDJFgSn2LiZeP1EH0YfLvAs98hSpoJ9kkZaTJyYElGVwtIacyPw3Z0
ys7F2+4EOg7oGqmXUasHf/Ih35WsLQBP+3vQgv0bRKzA/cnzB6kvH1EXER1wG7gD
++twx/k0nlzGYJBbIv02qSQJtrLHY/6a5cYUNf8NR1jLdj8y0vzr/M4jBf1Wj7dy
SYLgug8DXCc4x3DpB+w3YU9H9Nc5RoM3rb8UKblfBwPun/GBxUWkM8cZBieAMPjQ
o7lO4IG444kyOE9Gc3GaAwmT/Lx6O44Snido9X+T3Bq6LDaoGRtSub8WrSZG81mr
q3/SDaUDbNu1c2GInCkzM/DRUp7qColKtebKRE3qcoYn1RKNldN9BvzhQIt8j7k0
8hModU7m+dBwajQ/gTXs5PrLeg3M9ND02cAiq5fTOH6UAEC+Goa5MhsvbErnys4/
FWLTedcfZ6yP3rIN0aF7gQZh8wOOJBjppNYHyqOazloEcbh++XI/lJXR3ivUf6aa
TAG1CgjvKczuA8Hw0xZlwI9GHmR+hV8LJY5nJawU7RjZ5d0btxBr3CPBCed/xyKV
yMWdBusipaTK2x373aQhWCLPXAh6XfYmZrbvSmEOfxPXpR2jFAW0eETJ+fIYrbi+
R6TUF5DykSOEi+DMIevqRDmv1DSbFRQx7YmTRvUvnb3BsZkrqvK6IAh6HrRFCXqa
MwGBA9lWTDzpazBlniVoVuEFTH78PBj0XUZE+7SSFNvvksO0//81ikEuplwiuxdn
L5XC4dgnip9Mbgn1NsHhLP7jAwXj3kyMReP/f/5qFKcKWyHYiAGjp/xOFApfBYc8
/bx4e9T0O8o2ZDzhve1iKM5Hq0mOuzF3DjVJvE4oiXsGABFP+T6pAaunF2NAsPjz
hDtPxnWFUbVrWBjKg1+spXiaPQ+mIpdo4nS0sPakW7xBS189tqbChC/qg8spLLVx
Q+BNmi5xIXJGzp/3t52fsznoQxxlBsRHiYf2ee22KnTXhoDgnUvQa+QB9SCth06F
nU5WMbEow/5G78J5GKiKXnbGpBKvR/fpGwhBOUWJ1Gh/LRGiVXPSUSOkX+2zqJIt
0lmOt9su8BRWe1KOrwDiHk1AAyQOhg6gL24Gam5gn1+6g92kPXGPVHi2AQsHpyqM
+hwvSb4TbY9xyNNx70pX9Qalxjoy6NOPzy+fc75cwJlDfnsPj+BEe2+tvPy0S01d
Sujl6OOekq2FP4jqoPwvtnQ0a4u/CZXbZAuyx5+OqzVaFvDu5ApfR5iSgoJI9qTi
bkGzeG7PSxZqqF7GEIMlsCwefRMuT0uZ3tHKjoVje6+UmoydRNDNDjXpsArgJGGi
7tV7ozINwoauFrG6+fNtDNnTW9v0i5pvR7l4UdC7o7xy1jnKpwu8p5NMlPhGwTHx
Pva+dsHjvqi0RquO/9k6kiL3o/17oi3evEhPKB1+aopVvCJXDuOFSlgL1N0Og8gZ
XG96S4ccdGtPvp33lUUaxh3Q7j5kfghqcJA5dGe1JTvTUxWR25QxwVV2cPBpIOcM
P+vtUarahD9TncmW5OsKXiqtdd32no7+EgZxkI+RHLIoqsYMm6lqX0eNdQ30LONr
zYUk8n8rRARHJpsKSoJ3ld0rqAMpp3EkB4UvZ54tp0dxRfGXz3jsaz2ndGz4ttkC
hb4pm/PCoYRiTQnUUXFtkdfVo3BfN7x79EKI8x+NbeBXnnIQk7CMvxA64qkH+Ltn
T8VAQUFbCcHnQX5n/2a/8d4pUwVaqgelua4QHS7kaB1V9+iRV7T3FhAWBg8RdbOv
SBPDfehr5g4Al/NFVbQCTljBWGEGGC/QQNAvqAt10nWK9ulfVxAD6V6P/ZmP9DA7
LuORzPJNKd2WhE+ltbZhScMiQW8sArWs3qy1K0mbbq/15Gyi1/fgEovBnzkl98HV
VW87YS/yhQy48UCz5x8nLVxeSEH5xyKWLMK85xmuyARJDPlHRm7cg5RM9rJiE4MP
QwQ4AkpuEouh8kywugHDiJEeYp5WU+ZtQ9rO2p3RAdyXu6SsLHvFz1Z0bIRHH0V6
TFb11WbOFg0c03uSTJPNwyi5htF6KKelIk5yieRD9Q3oWXYbUnRAIFSOWZnjC4Qh
nfy//YXZkOczRHo92ZXQxpMpxOP5VAZVWHXr1p2YcOMZuqQrm/mP/2M4qsccLq+P
161oD59vMXYNMDT+cRiBQTzCx8EA30SzxZyty/dmxvibVddwGyoiL9iZh8zD9qLN
YKlVrHaDkK4iE+0Tl8IBxdqE1Kpd4AqTVSGo1NOdmVqxyizdmrRMxo2QamTYYbcq
i3N+zel31rG0rj9psEaF+763/rlnVPAz08olZRzGgXu9VU3zHWad+IHFrbeLhPm2
sV6Au6rcCDXsVFgPyWFmNK3JeitwQ5IrqTz0SiJ7oNBhmq//wUktH/cUtq5uk0l5
H3Y4mM1t6VE+7Dk4LcgjwnxMz76x/l+udiWRRvL0cqVbLx8Ims4paT4Oh9QSZC6L
ssdUEHodL/SZhA3k0nQQvh7xyAHzS5vFVl3sLiFSdzAAA4/SyWkzhWdZgBgqztnW
xVmm0K88olRYBrCR1fY8eFjKMYiuHMzDzGUGbUKqOTbApHB8AKftBuye0UJA/HgW
6in0yFwfMUPAm9sO+e3CpUxgE21pLmSYohkGL2HE9eJx+MKTZW6k6WQ/RIFc6xYg
F5La4N6HCly8XTav0HGPA7Wm85VlfXNm05w86BLpjuWeZZzM1BpyT4z9uODP/rJz
eKGO1F5QLhgvl3vVsaK9RpxklsqBPJ/Tr7R9xWuGMv3V6z5jrEok++//h67s2PKd
cdvJg0DAnsf/wVPmlip9PEA8ciovpSzGM20Go1gSGygXuQA+CYgrrDvtnNl6Yjac
4LYZeKuDECX/ACaL9jquqOntBFVd6hLJ8y0/duwLJZSIAEa1afR/zJ2p8bONvWlw
xwEs2B4C4nG/1hnMS9CGsbm2m5UmmysyfI/1KO+sp4gTBfw+MAkuLqrXOS/lioIC
C3AJ9BdaMrami5pTVmEHsgm8BchM2PvhdpIitIWxT/5oyQz+MHRjWjNqFGXWHt1B
C6MDkIK44hf25WV0eA13CCLBeAHJZPeQCMxj5fB637HTnruem22q7S8xL7k5lVfG
/K0cXemY/w8fKz+B0EiId2UuC1jRbJI7VqfPaOv0kua46veWFSaWrnqbw+ukWG57
ndI90OKjnrTIWcqCR/YuveSb01JIf1Slnix+88l+djKxILtp+PNnNeuR6kOjDP4N
e1xzQcYxs5U54PrutdVseMjgjtgfQ66iG6n7cH+Qe1Uo5hfYBhRzhGcdUhOZUooN
c1VuenXCQFH50g/VlZuuZgU7ZeOzSjVTBOFrMApOpIf1h1+ZAgh/HGS+E2c+f/ws
8bzSMyK7fNzGTqrkd52VP+nY8ksCbegzB6ELFXedx/37PBKctq3V/ROWmIJDmmU8
PSWNVgOsVZhESPFYvS1B7kh34QHXwsq53yifYe6IjMV7krb0N0m7fomWAd3sDn12
v9EC5z/WNebcsWWt8ylA+dPc5lotvUQyPebYjZuT0lrqrsnwFQH6CuCZ0S7FEbDA
ezy9PHvkYsDxchjWgBgmaNq2XsG2wD7mw73/9Db4g/xAs0ijREYwHlsgJG5rUMpJ
EWsjSvE7loAkADkLkmoQqrJouAXiQMGYWVGvZYSvUPTr96E9Dk3StqEQ0QW6Q+OC
kg9EPcT/pSpYqVbwel2uUFce26qNx6xXnokiEBW+nmaTP54BGkCQmexUfZgSnWN6
gDL8Kgg5dWzu2w8P+TOlXmFXQ30SArHTvTghSYLAk1j1loKSBiMvjoed/ZuD2obA
W3QU28fBtk/WQHgR9hhGd9/HnbiuwJGgP8PGjf4kiLk7/f6/vieKzSXphEyNJgHk
p3TTX121OS2OeLAS2JJoLcqpWFkkeeZ9yjU+bzuCJGtf34RkL8FwUxTL5g0TSyHk
+koyc3B1o1cIj2Phgb5Tas/GIwUdqw++g1/2yE01u9CvFxqjr6jHj+vOZs14jmls
RfOTLD7wnQGihKmNqKiiyHCkerCZEbIjLYHM80GxVBc4GpIlnCf/5x2shR8puj5h
NlFOEyCkUDFsorhHPwRAI+l7r5xx6i/YZmd9C2buLlAKi1vUlFIMoiT0GTpth5/C
zgZiSh1ETcncceOkLc8xM2bqyQwJcZzp7hxRHIiIB1HpaWjs4I0WZhiuYTvRPrXu
iDav1PwQrCNDHukld1X0n/6Ka+YjkMQ3Bnd90StB1rGPusNBn3C3oKv/zZ2uiEtM
Y5HpKFrqPGkVAcb2gIM8F7RMx8kjY2X0ejCHdlDeH676HASeQgKU0Htsl2U617OA
e6zy3hWvnw0UZL+FAApJFpMJcAuI6o0Pn3Z8hGtaR9keBF5O7gMVHaC633FIUNbY
FDEcWZzYgpuF4tDXlPT4G9rAmDcmqMheLuPavc0HJgwv9rPihpOG3eDj/weyAniC
MfUPxZGO5fd7hCjDw/dTK3lYWViw1bvzq42YN6QO67cGyFB9gY32qUflHaO9YTdv
x3GjFHqlmKtg+umEeqVkxrJiAcwAOfFcR5/1N/ROovqqWRDOtft7TCBEsNQo++Me
FZRRv2GBrgW7ltI/jfrnIVy1MsLxCnIdzMQPzBkkNDDYEzIjaHEdk2j94+/WDAtV
Qj+zrhl17Oy50v3UrRNfUnFKgvjOiXlLdPOLFdCH0daRN2v+5xaqdAGKijdHTVVZ
8TSIja3OJL/jDVFATwVLLRXv7oA14TIaJgcQSSQgnQBndhCXrsh3xxzsGZVesGbR
BpdCudqIlvhcppM2xeUgfgGLB0y8Wze9AwXP3CHYeBk8MSyofJAV068lhrH2DPyQ
hfR88aOaBueqZombbR91UhcIw5+2BTtwRe0d8V3mgd2H+wycOIEZWjq5fneTx9L2
LLHV0vJ+YmIG/+LB9OsyZWU8+slyYFsKDkeJtYnhw6nZkJBP1PQii4PaIrKIGovZ
YrkQJN1K85eVNUbdR4W0uIGWXbjuP1q44Whm3Fa76JzLmrXnrvg71DTsKqLm+DXs
iZjZn3rpHGqBgwmpoHQjO79LqDzbexBDwFXUkCp0pxxIxfcXtga1OQwldCJ5RJqc
DLQ0zpYg1REggo3ONknyLf0KHBQBkH91XmxowhzN0iUVWR7bSk0FE12+XpWb93e/
vfJJbepdGTOHbYOOuK13LrJuB2IfBAtO8m+z4V4cXdWf5CPpzBy6jtMGlhbXiW1e
2EfCWR00dkTpl6eIC1Mmljq+D3nV3n6m5/0qw3Z7xZ40Xw1Xzh0MInWXaIi69ecy
kxiluGo5/tLRfv/FfkZA6YssmivCHjeBXYmRlCB6BkrVXY1FJbpM2mRJgIrC8+So
RPVnpdJ/Vr+IPgKanzp+4eqF6p2GEq6zfQGa88NAJ2yazv3itfatTCEYYZCcq9nr
Yi3HGr8X2BJlahBKKKVmet3G8qshsjVCPoZw+uSQSZMjGX6ATRrW+khUX1o9N4bV
1rBeGIQtf0J+PHg8vRywzEFmyt7YwCmZc8fZts4NLjWDd0BJfNMTfpKR5Nc9VKGt
7XvDfzltV2jZRRIU41lRRtmK8Cp7cIaInaNsEHMU0a/Q94i3vxHyvFK7EC+9N4TJ
qzeaqnVOI44AckHsKm6EJyr/q0NlnbHfY+ZFvmrCVG3MozDcn3jKC2i0DIYJ+qSn
5UXjTFfzUli7S5XD5CuUqioad/YjCxR1eK49JsE3V7kf+hV2rjQ1rPDv/RzRYmNt
ZP0NJakhSE5q0uYYkmBbbsrnFaTpE8pXmRPS369qyIutLsmGVRIktx54sool4DTV
oE2UVkhG/DcYV/MytkfoYV1aTyLEuA32CPFA/TasNOd3AeExsGdEkCZbFDyyYnWC
ot1Y05KsDKxz9P2+j3+HXeGS81HF7p8LHn85Hec2am58lILJ+zXGZIVIF485qKVS
g25HeADy72Py02HkaUd6vlSeUMCAau644224pPr7hBbwmi9DL6Q0mvSpgNpN0bSr
mSzBEYocxh2CsoqGTvQ5HVqTgaH7Zds7pEuomQrNELAzLjfRfEcrwLfCmrUUT1uZ
7Q/fmEjXzUWaILWMVBWVSSbgp5vtKXPIuuViUnMKcaBzqx3V7jkxfOMEJOHIV/2i
G74bawwTWI1ZFcH5tWO6XerEWx155hb5lgynxcEK6ZWFnM1r4r7zdHeU5JuWcyKP
0NLAOfim65KhoTmkZjWUgkyF9OTCx/qMB85XNzy0MOBVeEfA0iQdLrdPHESuqbWc
adXKPQf/Rc+oRVkyPR5JiL7NjqI1Lucm2eLmIcoJwwlzTwfCfRPlXYhRx9uWMqRM
fzpGuPa/WbPEFBGXS/JckRFjGVKwaS8IMoWur6jXjUQVQ6eOrRTP/1Avn89LcsCo
iTpQCFh/YqAtBxGnDOKhBxwYXXGHDYMz2GPliWOEsZcki+IMFWnAsLgCVYE11ZEI
nQ7q+tHSs+NlQPCSsBU94yG3zgWbtK3vEPIhYp7TGIijko3Y7Z+6bQ8kBScddBHn
bz302LMaET8EplhrnT3ePY4TrTIQKop62OYw3wEDrSra4KsPcrJ4GFCZdQQfq4gX
dLQnLMpsoHLAkIpU2XQb6a9EBY6yJ6b8UMTq3eOTXiYTZHyZKQgCHtHDCHA0p71W
83CNnJzCZsCs2ET1N1tNIHBFSKlSXm/OUqLzIvh1fgL5dmve55ZSzM+CLhm+VZjR
4WKzy2ATUU/k2gA7EsuSMLNUcZTmXe5+uZu8DYxEu4gOS9QCeHFodAZRdunqwcMw
fDzs71kMxeI0ZOt5wQy6BwQCtkHEfUVKFK4Hnay9/x6gTzFVP/Flp4Fs22mRHNN5
3D00/BIUh3rgFO0QgPmNfBoLnW/ayeUKVnNmx/v93FVLc2ORSWZsWEgvPJxrwCOw
+8pBwZ60at4TKD/Dz2uj6OfIzbEckExfW/T8vqr38YvSXAO0jso0ddOu8PxhfhXC
Z6pRfsTCdY6n8yVQ/6byX6CkK6AGNiNkWLw8O8rB8HZFqk4RMfNmsICUNvxdfsh0
Yuq4LJYCdRqJLOfABM8Tuv/bp8SapHqiBYIpkNXeCEwf7s3piS+GuLzDXlUaexz1
oMRBM1xTlDnp70SKiQSIvS2o7T+bPblOnOH6xS99rRu0mh8oty7DMlgHk4oxQ3JB
1+36YW62evhoHJ9VECecs5w4JRAT9JuZlPnmPxXnr2GnkrgKZ0/ccfexV+DSa/Gi
zZ8ZvYc7OJkeh0lUTIaj3aqLa1m9Bf3i4tgOaQ4h8iIg3qpO7goqADbT8IDAKrSa
AeqDw6Le2k6GGy3zqQ1HX5yS4v/tTx1Q4THQpHE3gUmreV9AhoNjytTd72pfbNmJ
QCDp/M0FxaCDLvAik19z8VzC1LLO86CRD5wMu3d/Vn855PwSpdQFMD5NQqc7YPNx
Hbj3Orxz5E2kI/g1CuV7WAkAfGhLBqVDCB1DfxOQfeZXTMyV8c22+pblt0F+bEBO
DpSu0YdiDdhX/LFZ777aCN/SL58EwiCBrsYyDm/0dS2EiKAE7paYbgJwrrF5ycH+
lKOqsAPMJmWRNBzvyFQ4onapQI5bz5uIZ9MbZczETkgYyCXI+wGpICe38h+VUj+n
JmxxQFDX1vhWw7d46bWEl+z/7C/mzxWhTDBnlCwpZC3wLwr4uTkDCuvhFG6hh5F8
fFLSNFZuwseTfrQhbOhHDNNLnALSRZOH4iwQczu5lAAIIU4qKbjHglz+tk+w0gek
j6rYCQh5M6we5bHTlTGjrBDRY5XRcXMSFyv8X75isHUDk/dZETSI18FtWcdCuJVv
rUprPzG9sVj0ABDKyqXjfiiGZuQwfNwYt+U91afIpMHcX7YmCSdlQTLgmveXECvF
O5sickYJ8Cvu/u0xLbeW6LLEHgm2qXOqPt59kKhVK/IbmCsz0yZFfXqmQ8xW/AJE
73rO3kwA/AWslNRCWkN7K5Pwp6RbG9phLfcJb9IhNmGj6R9UuD7cNokbqZyrP0hN
sigmGD3nJ5QTM324f7TAVE3KM2ToZtrXKsbXy/djGX9rgna9G4vO6vKNqF9jYGka
loJDG/nhXKEpPlsIv25uJyZtoMGCqwP4gIdCQEC9nz9QuXfKjllspUubrUuKMQVX
Z0qOzDPnwSYoZ6maW6L9KQze+aLhFWKLBwFunzlPEeGrnuhtz05+0rsszPWl7y6P
QZdX52BYA5JT22ntww0pQb18MTF2DGVyoVAAWU52n0I6i382xQyIaMr3Gxo8w6wG
WXzs34jDN3cktgUqJU45LmMuDQ6vMi09iLeybS1hKIuJwFBVdG/7763IT9Y00lA/
f4Z62/cqyzKBfxx6g+GiJsr1j+ZDSG+IHnGHYlx5s/PrFGwxHAwcQM4UrhAvTLLy
3RSt87RC4Mhg6zu2eejpznzUs/jqEQXuKEP0gJxSnxsqens76U+uYqana85OVm5m
z5JQG7xMJ40GVpU0njAsbLSQE8hhnRi198/sNIbIAxXhNfJYsRWa+jKZxBUxLU5L
CI2RoJ/GvyyVDhbovkfbOmWVoldd6BiLAyTDjNc3lx8uZpXic7HNZNQ6IJmPq6an
mLyhnG5jvmIndgL5dabma9FcvXrpfnzoBl6CmflK1kwEsUTcnoldjH8iIWrkmxm5
9QpyuQ+YNwYeodmeZbYlqRjAqS0VUEQstX1zsgvscdDowxHAhhKK181DSWH5mEbT
3pR1v2bdYMUn47yeLQAuPfmwOVKC56fgWS4yIqa79ZB3T02J8XfFkJvdBIvfMDoC
ok8e/kKdFVVuv3F6X1pFeEsYBw0JwIGJQH2gt4YEzY7wthjxsTip/EHkO0MfNY4Q
HeVQxDObbywkHnuugLpIdB4iWexUprt7IuWyV8s7IS49ZCToZcLK6I0ssCrbrqJR
0DWDUehdg/kA7FE4y2Os+iyubBJeUP7dhZakSKLMdJFGyunnUyDCIwuilRZ1e6Eu
P5J17cw5dQVEvG2Wm3e0XQIhJrQGGTigfChv4XEGk1bLxeQzLe+waIuSykjD0aTc
pht1jCLA/Lv0icDPB2u50wq/r4PJVLUmKkM+mW03CT3Ojgb/KXeFIycZGeN/KrkA
6a6jgl7elxG3pfcvLig59TDeVPHWB8ByuEE7t9C4mt/t9Cxt/KgKRF8Kbe+vlxhi
lQ4kg6nZWkk0i/e3NWzqvbcVVYyFc0L2K8a/o56kOll5kr0uo/7WlwotnUoXjaB0
caDp5x7whB7mNLcO/hk4NrsKYTXY1hpNybN592gpi4N/4OZU9Jup2JJFXbI2plvJ
Bzo03rR/wfxO2Y4x4JfiBEJKoKxRhd4cbKt87GONs+kGvfomNP4KF1t80RG3ftET
xcBvIFwl3/Nj/KABra6BJDfQxVScgfuNizyNNjl3/qJU8xjhfYzxGe6qieHXI2T+
rN4EBim6kZ7ZS6375JC/hiZG1DB/dBjVltrmcwXyQn1odTUDZ6vo9BsIO/GqSLOC
iyagp+qR2Y0VLqTMUH+ktFM5uBPd7ENG53hfYWgjw4QYR+DE+qq2aJ8g0edQyqXo
mCqT2lykuSHP/CKQWXDrXSd5m/6LXvOJAZrgT4PXTIGfjVK5uui1sjVkXA13fPNJ
rNXPxNC709pVbLDUXkO9TLgdODuxeuxJmwjyvLJXl1iE0AaN+lrAKoEIJXaMplfF
1LE5ArQOeupz6C15EzHHPGs+JA4qJpRKlygBmlEnDwepDuQmtNwyeib0AL+Rm+5j
2cKKg6F6vcOETcWoaF1JdAIDM3C9J5/L4SSj5tMn16DH/XH7Iz7e6xAcm2UKuoHo
W9RuRnhcc/s1PNkDjMJaTxaZ9F5vXKXqYcNNvAYpESD0ODhxLOfSeverXg0kRNZ7
Zb+sz5zJc3eb6n8qRZkM4xHY5xHG9cu8rJNiDVUJFvROKMa+57oYeMERTAO0ldY2
HDR3WRWasc0p77MYB+y4jBQCmXg2t1gkfq630vzIR/Wx/oPMawYXf+1KWAvED5go
NzKC1n+aZK1L/u9h/4n2iycBBusckYrwFtsS3H/61ueBDGeITmizwWC68Djpas0g
+bMfOhgecnsOVP8m4gzRZfy+W40zIZEOrR5Pkmx1+SZrO+qYuI8Tmr1CTFrMnK44
qvLCOC5bqKb8n4moLWJJzfIkWjH15y1MCmMHx3XCkbYv5mKn87LSf4OJVu3GBSRA
nvYRKaJ6mkiqvDNjk2Xog1dsWW315+s47z5KoDGXxD6BekmGd/wHzBRuYLZTRUlV
y1v/aXgIsF0TQaqM86abyyBrO0Z6NVZuqezuj5+h1UNoo0INz6BoMWhjagyH/t43
5OPH8bPmzmL6MjWBa6UWKhVkNd3+yjC5xDUahTPEEoks0H/X9VrVPWjGmGUCg8VO
m24b9FObDpnuXbsYnaVT7h3NUQZhjM+S2CHvKUWGMNtsEkJQI68ZrqENsRdEDa8c
Z5AkgQOYr//wessiS6xACyKDzEJlcQ2wAzy6J/3edYgjCziRZCpEGFoYvVPKrITq
kDYY47cBQF1SM019CO1fJuFWb9uWp4LKF1UGh4yeWjNr0uXMFQscB5PYLxUgisQq
clowLqcDvDqCGKnmzfZ3S0anlN8qAVqg2amMi4VjvkopNmXgA/S1s3TIQDw+RB3R
t4AkcJ7a5fNXTC2GOe8N2RisAGHsM8rsdNr8URXf5V6+3bLfrIOejmlvefAJYMvp
JTsLq21ig9H6fwXdWKT38L0ojdR8tbNDLC+AFbKa79V+9dUDNvTAwHN6vBkRZyJu
fjj1lTmtCZ6A/Ua3VuA+/VCp5IoMfSbpMk6EDwJGG+RL6y/lbXjS4n8Q2HjuJb8x
ETT4zeFJTXR3ENYZT0/OUCIV1K956swWQGgBuej6pfyYAoPSv2h4ONnbWT1v2Iuz
b0Ifc75Oks5qQXVBCTkmbgLlxIT//PYAsb+iRI/vgoL4kKi6RCPvWs8C+H8NRbAS
eEDgzFzbw14Bez3CX3FguUVDgmN0VkSgyKy6y1v34TryXTmLBbhMIKfGymQbZ8U9
i06K9hGHYuaUJPvVBdgql6F1AymZTwI3leFiuVjoeBF+GyHIYooNYpQYDSx5FZuQ
4K7vN8rYtWj9bvSIN7x07TVHBhs9RB8CDFj5G1q/mycpdRDjXNOBSNWyui2qBUIt
48t0sSq/tD54AdcjGROkWOfgIYTwOxZd6wxWIFIYBo98Wf2o8vn7VddtrX0ICScu
VC/i41uCdfQ3i9RGDVMy8nNAvoP5/ge2f1wi9IdUYIbGmyNGyNCo4siUOPorTTLq
dKg4BotD5RKX6vPeWOpf81APJrfEQmElUyOmZYpJYKZjcR1FhbznE8oL4MrrDkE0
nPR6SzxPxs2+czbSkagzRGDcv4n9VgvN8cJs/vy3CeUvPNKEEftgQX8JDcL38et1
asWp2x4CK35Y+5FqNiXiz/JNZIFAdJNHOsXMEqg/VtcTJ2OID6xujc6yr4rGyXf+
OzWoTru7H0+GFLuh0H2AD3UNUY66f3nBPmuXojsZJpJ/UUmRcjgb9jQekSqTBnbU
Fs/+ileT4kNbtcIcc4moN0e118XrlMzGeRyrsg/dkcj1UVXt77N6fPAYGRE9KiIF
8Q20sWlfhF5Kefwimg4cUlRFH8fWjQtsMwA1MeQJYYeyQ4lUIBT8rK38ZjcIGKjo
6iilbvejwLbiO2uvWg+mL56PVB7SC/FsVc4bW2iYy7N9/xf0Qv8YuVbZAoXnmy8E
sEiDQFdE5GYwBUKwLeWvpnXwI6+2HhsORmjRbUuZA+n8Jey4fcM4t0BcJyE57gPe
VJUMmyy6v9Ab1rj5RGN6pEF6seLbUqCi2Sp7vIjjxuR70C14PIqprcdf2jPNhKTU
sVT99yQx/ouHDFy6cXGz47d6kEm9tzX3HsxSt851Edji3N/PAEFuHgJFTmNaaEPN
JQaQGcL887tV/snMvtlPOzKzqS7F5aXAKcEhi+flc5LRvgluRCKWPo3TECYgdAij
QOnqhH3FJhH2Ph2Tls5Hp7FbekNb6E5lbeoDK9gxvYtvgd3SWLeu2JZscAEg8W4l
jmLaxG5UcybiQApLn4qiTcjAg1FPJNzHIv6VuiCE9P5R544ByChU22KvEH3ACxAn
T5KD7d//QJ6Qm69fvXpeNo3bsQtJp8B5oijZHA3AJzZrvg5mxMqqhWy/u8k+41AL
exodjDVsZMjTjbq4RL/RzNXLTlmafsTpD1qegB/HH+iY2i7kROF8qsKr9MaGQ9ho
5ij6OiS5oaLsEPjRT3l1fP8uZL+Vwp9iHhAxurwG1Vz/Sa1no/FlJcdTVu4EC9Qh
UHQn1fCCAYAsYlPFF/Bev4rtysh6nl+3Ye4RCfYJ2MEccrwkK++TlCCNJ/q0bhOI
peK9nPt7l4OwLwgt6PaRXmhsPgJxyhxYn+/A+RUgS+z9z/1M7Q/HaICOkR7mYqSd
BNo6pKuQZxGtAkANxBOHBnyfbPNLiP0ZWEsLXFmJACCi89IjUkoXO6e1OtJI81kq
/Lko/MviJmafBZYaQn3vrBVNgoFx+31qWpLrXiBKKBQ36/b03ZHsArock8uGRZrn
Z6VQW2QBedUgEcPEn/OvYqBU7UEaX31FCZGyGne+EkJuCOUoQ+BkLSg5BiLHqtiE
frOGzAhn1AHr3tUFrCuMrMfoMaAMDZnU16dIsf7pdlkdzevKIOHiMcH4Gn5CuTyG
snekbSDeTGRMb0GnogcjCU91e/fx527YMTpC1arrXtONKhMYEy3RtxZiLtOyEwtf
5WtJQhWHrW00Dvp7/i+6Tz3o2wrXR0RnQIgIkWB+0prflOBQ4UBUAIEXlENQEhyi
pL95wuT1WyqO1K3JMwB4yVUPPIhLbRzgoc0r3p8kkxd9AwwDX1NbrEiBKg6/Oc4h
3X+joYa9PD0FPO8kF7NQz0U3WfOMBTT9Ht9hAhBTWVCq10kIl/N2bRPogIkGw+0+
LWk4q8VsSpvQbtDg0B870wlqMsmtFCnHgFgHu3uEAJ5ue11mS7Y2BHFEUDhkm0L0
1Mc5xl4OXBvXI6OaP6pvifq72Nxs1RPPH7b8MR8NQ3qpA8AK0NyerEtrMI/z6ukV
FFNNPWwIumR4E0W00KX0IpxV0p6bB7+Uy4V6GXAXOs9t+GlueTlCXCxPTgyqyGMq
O/kqii93xaAg0Mj4n3Lg3fytXtQmaJCNF1Bjo+jojiF/iaHVw4hC4frXYKbzjwgC
0N0g8F0eCKdv/mGGYR+8QMAoLrZeXbf5LIfWik1S/1dPdVZfEhQBSynYtBbDPPcX
AMwWaCvuWQ77sVy3LCeqv/9q/NLbaASk0KnzE+LOHb6cNx9ECSqoRYM8UjQNL/+U
LwC3e1u/FWABFf/HggELFu2AcL6QJFHnu7NksPZ1/hiXbHaka5m3IPIrr3fc9o25
xX8asPrhturM5blLApqlv8p9JA26dpH7GVxoajBsTBKyPiyRHpuvLq8anM2h156a
eyUhD/W/bQA3mhA7zqKzJNoe7xyOj8RnI4um/k93Z0GD10BxlBy8sl4OBou5YVsK
YW57WEzo0uk11x0124y7lnylAZMhcbXw0NC4STxrK2KeJU9kcOayeEtnPx5tg00v
6JVH5pjxyhOUFkHVfipAC/BFCv+CzF90EwQgcJPaPJPAc6a/vk0Fma1BQ8hQ5ngO
5KzrLvfZafDxf7D2lPq5oZp9ZMZN2U5wQOutNUP3Hu91aq0jJ43BWQ6RxhM+bXmS
ss+ojYJKoQtCvFAK5bP1UMM+6DktSqJ1vUt9LVgAu/wXbMgrPVKzQFzCKBbENOMa
PzupBGb5CHOZ/x8KfotqfEc9UJEbNjj2jt3euvYyz8aW5GdwW4p2/1Xshb79i5NI
iFZnz4dAFeBacPgskOJY5TmtYpQ/bdRi1OTv++GodzpRV08yA393d+RLBxJzSs9I
WrXkHB+0xGCVnqytyeykqE4Hyckce1mqV/9WjlGRWISbVPhUItAb2Jxdt6UjdZdV
K5YtdsEge5l/nNMrk2/qYloMJvaCqkWK1hWpvLw+nPZP4PrgoPgdUIs30/HTceTb
/MMmhuj74FpG80n1ihf1hELsz7NYmpADhn6dHyWKI5lcHIx9rHfsPbV0JTRcNjhy
3zS98zlUxj70VvN5ayC6GTz8CiHplj75CS2u+vhcEXTyAu4iN8zOlf5isq+tH6RP
edyJfPWG3Lg6KOp93x672M5fozWr+MVlEFjQHlFEPSeo2UHEeeudWVnBxO5/h1ZJ
jjrPzMLbtt5u4pGeKKxW2bvc/haserCif485ROiOIb76liVcQoOx4W+ZKo83w62d
enZVe73cOF71GgOo2xNeB0Nn7oyq0Ll+sbJhYAg8ATlwjzr4Ukk0Rsamzj/S8H/4
mKjoqUlIp1ffZfx7WlA01zyZ0ZpD0mUJuTCUXovn9LEbg7tb6YRqtyeUh/m6qWB3
pDQoleEZkLDnfwrJoZr3EbRwRmHNyzkzPVQp91ehO0jdpYpjESlki9jWKoZu/ab4
NtefhVgxQXCj8q7IYf+pBMzr6mMCPr2r21aUKBGhlwVruc9Docu0ABkZworl1mFq
uWr3tlcEy6DtpMWYd+8UWnxWoZhB4ndLMS4nUYoZ8lN3laAJ3aIWAuEPMwZkS9qc
PlOdhb+346l3P75fsHLAezH1I30szfcHtuWwmkKcDRnu6uM+gRV6c3xr3+u2o016
E0H6YZvKaWxzhegRoZYWclwdYZW2KlZ+LLaXH+GncW6KvCdIPBnE6Gooj9DZGglk
DizslVchVM6vvS9qATqFRdgv1Mogym1rSyGcSG8AQdTCdkJlbd22M0MA8DYzXFkP
fcCyYYmbJUVsV1eIQXaAj5PyEhRU7s5NXa9u3CivzutobdxageuoSrRAKmozi6MJ
gcal3wCTztgfmSGheBVniVjhbySBg8de0yMkH8fCC41iAzJkcCn+txtiy0h9nP/O
Jfhfk4eYvJTku6bXH9klGp9ZbjM0ZaRhnIZSkfK0IBLl8L3ccGXIGN8S/5XlB6Bz
+Yuoc2lCT7TbkG+YxZ12kfH0IA1nLfmcEQDa1JemZfUH04CSeOkBckUkEn+zGDVU
t5qHcTY+LwYUexXfUgQJ1gR/7x9VX8JQ6Cf8JQXgs6HY382NRx9To0RpJ/cDpgz5
oLRIwKVE6vBsQlLwdiX1LJsGwNHh8Zk+jnKHX3jffkEw5N8ZE8c5p7C4Iog1Ueha
+Gva84MpvwfEhkiY2zPsy/TA8b/7baCO3ab1s8lmr0//04Em1QvcVPmGT4UXKxac
MJadl+KG/8wniSK8AsNS6LhSLLNk1SGiZ3HiO9BnoczSugnx/YIRIifrP55SLH8T
dW+Qq9DM08nsDZG4kj8NYEkIxI5rZl1jIpBEVo1CX5EjbL0GNo80czshhdqgXKo7
Vw5wRHgQUdKxMqYUPQ+D1KnFpmsyUfh3x6wx9YQHh9GKQ9ngRt3p2LW2BSC8JjT6
6Z2Pc/j2ciWZb08wGrlU9kUvSOYWdHqHDoXMnunrKdzZ8dnT4Xc5e18P9L1qose5
1fugOmDbBKPSlsn3nmEf/6MRh0Qrz+/MofM+KJYqKhnjaJUzQBFkaa1U+bZeVm3T
H2TrS3ru+ZjDlXqxf0lKrbFr7fuSajf8NnIQCrq2QyzfT6mV1bZwaOczDo8F+xp4
Qi90ds68sfB6fI09mDMHWFreTDONMkox+DZtEXB8gXX38pO/QrI6/dGJWvhS4tMr
rrgCxrQigveLOOT0W7woHBP50tELoaVXAAF2OS2dOcgMn2rjErlzZAVxXhUmKxvZ
s3iPu3LMUBI8rwhcn0UAb7IELYcij+ByIXBMP286Hjr92sKG2WgqVzUoGUCuN0iz
Z0F9lVbh6aQJIFcReSmN5qI+R7V8TZfoCWdHNKTRWN31gqRhRCzGKFkk2rUyKk8G
R905G2/aOLn+G0JO+vBsSe/qy6B6w0qW8s4pm6GgP+mNyi6Imk/pZ53QeL5N4fUv
jC0wpztKakkrk80taEbsAxJsX+X94ObzL+igsHyfz5v41jh0nnF37glANIzh7Dkq
XTivY7SiXsk2bYIovKuNdYLYU3upL39QvIgtBMuctwPf+4Kix8MLtj+wIKaDiaif
K5Y4iX+0jq1kfxXxJZcLmk5p7fj6DjoPeGjZP3BisR4O5HVHGUsYLoMLA+MXFF8L
I5xFPmREfBQ85FKa7tqgELcIi3NNbAJ3ASlYXqhn+LhKS39Hv2iNQ6sTVK+ho46c
kNef7tAq1v7Elcu9ujm8BZLeuMZiw2gjM/EQDmP2n1M+zIp8e+yPmvPi+yBIy6Pa
bVA1Xi7AxKlrcKGDKXfmXNHegC53Y5ywCR63PKviywVdo33BMkAL8Bordx9hwpyp
vVNHU9lYsodM660bjL1YYcsmTDf4ZIh9oxurat0BpwGCGpBqp7zMCpP6vedDDDYd
zHsRtOP3tNxQLmHlCq+0vuRObqvXVXYjtsAXCOQviZRSaZmDAsg4dtdOr1DyIzXJ
9Tasl+zc9zjtjvBxOK4E1aF7LjbcZKJ28df1mkWklaRARw5mr3bitoJI/rr/Y3MH
7AUVJPwSijT44ZkieXKfLtdAp43exz3qUXdGqpOcmzcu4qU2lt8vO2614K2CsSkQ
nqEmF6Lc0Ncz8aERlYyNlSLMsxwg7rgnJ1V7nRIaINqeo5a9HsnLz1BR5LrWZRFZ
nqpmuMKqQSs4d/JOwftM6dND8MMP9Dj71WZ9kvzH/n73Cq0VBmyHldhz4B7P+p+L
SWZKGgdDeNmSKSqweJcFQXmqSpr06cBCAb2N4JGUiT03IoGWoG1b0QDtbONDVvVt
zANVU/ViAt3xuiGBiHS01U031Sfr5mbkcSv+Ozh3P9BdclOe9gbI9egJ09mp3L8i
/bMtlBUc8FvlC+B7e6O7MX+BlDVAqIo4y03H00J1jVXzzGXLuu1urAs/6Nyx0G9g
Xc/kpsKZA+OdtsK1jTP0oEwkigKFNCO0gOxquvIGPwmjWTnMp9idiprjopp4x146
tzqBGpYExgyc4a5KFz5PpERiKeyF3AujruuOHG0MKAHQP3SPyM6Y8OjYFT8bdK0R
MSJcTAm4OVizZrKJ3J6AcdQk+m8ipfVZci6Zgm1SR714WGu4/l/AWvMDl+VeWRpa
HSBqpvULxIk+VPkmfyJLpTsZKcz2lqKu7THJ+7QeFVK/WufG0z2Kdj8uUAb38Bfv
T/BI7QUdmiJ59wZiIVc22tlQ0eX4ckBeUFwCOIT15p4gViUI3KezdJEpIyHDhzQU
ozgviWEdXzO90Eb42oPhABI0xPu1vwNiQPxcvOdQdhhj0mt+lwxW78j7NyNCYOlY
E3SLQqEAc/dnqGQtfrqN/5nPJyGEfcm3YhTti2wZuXmy6cw9iQag8g+vBPHDs0Fl
LCPnsAwXBVV9nY01a1YEFzIJGi0D5lhdAuXNRzcFcY4OtBErvon8qNI/4Oyyc/56
AsXFN63AVJgTmycHfOFakXnV5eb0B4ZI+PsKUMVAvyvvHKEPRsiCjIGfAwWnz060
8Lm0qFDVA2Nhiut0gOZI4XSyg80MGYcjKZQxLFGptpcAZTHl35zr25FIsFjoNuLq
P1541QdBKXq1+OIZpR6f5B1E/ccqL4eATiwWaf0vsPeO5kUrc8ny+5efNtzVRw6P
vj4LEoZjeyVIzyHYC+rXktC/rep4Km6w/YZostXK1WCcsCT9xu/r1BjrSNfCR+nQ
DUALdLjDHmVwiPmO1FsPrcLL9f0iyvrh1hNVGvMaYNsw/9CgMSIJObbJ5FoQnDwZ
k5l4h8tskrvwMmmb2tRDvvW4h1SzqFh7UDgVqaFo5uzaxaBA7XhdcjRRkCuRS3XP
tmDuY1G3ap7ZF1L6WTDxB1QRZvE3dFuLg/1nvU+b+h7qETsy+WvDHZknJZGHalyk
HPSjw/F+QMHpARhx/FrE7xsH38aOoD3FEZs/bXrg3KbkgqOPjs5uPwuP+i/j4vvV
nspvZKrSaQ4hkYp6H09f5O44BiKpSt4+om6Rt5BN0Vij/PcK5JUH1HTfzKLLRPwb
kPFm+XV7Ugj96bd4aT49K+9mZbuobYEn+Tr16vEhyg/DDz0AH0ZHNq4XcbRhHwJP
FuPFdO9662DAzT32Mf/TjVDbXvLljvXaxV0U48deIianYFeAVHacwcnzrrHyGDK8
AtR3TDcP2k1oR0VgWRVn+ntl7B5u/KD2MhloU3cgrAP2pX/sKkbC7l13ck/PfPdi
Ll163rp3EZ0EQQ+DeH91Cb8eb/Ie+NCL3n23G4mAxua+2jxbaxxiuGf/PDARud6N
P9cMJY+nxyOiBL4RB+uqWQEeLy+gVB/cEfIYFjuLbC8u4lUQqMz+5SKHOGKfrB+s
4SrLZr5CKut3c29lDbGEqJ4GZlNWUKX+RVHrMcVbaDsikaOLUN70PRrW86uKErA/
4uOj3NPaxsFXe7kG6ndpuh8yQdq6H63BfUkJRd1mk4Ry8j9/CV8E+mNZb0rn7q1L
35E0+hDU7dvTpOiPNZ+RjrYp5vNBhMY9ghBvpSaOtFfvkjAakQNUsuS8JTkVNUew
AT3Iy9Y2/VfX1wBM999jbohETNTFxd5OMaYvpw4zBkaAjSRHqDpdyQSB/4eoaXuG
MFePInnTMmG+FY3R6pKLUwvKC93DiF4QLLjv0bA1rTkfKT0RkzqssQBPyedAwMAs
dvdnMcrWZ6Pxo7f+uW8IBnykU8cxl6Nh1p+0NmdeaZ4TYhT3QTea+yEXeKsy75xM
zf9mPTBpmgDU/s6n6Cm6o/uLfA8oiJgpmsug2LW3gcEZQLnfuO5qBrT1s3FxOEPo
EL8i4UaboF+u18PFcJG1in6W+foOw3Yx00u2pDex2NuM0w4DJJcaBsAlxbddT+d0
AJGPAl2/UeCJVcOBu8iEEziXCOsv6AqD1gMm77SzyMiuivMBAr29KVeIi3lvaI2D
Y2QlrFM5G55IXHd2o7gITJCTNFDZ5ujh5SofhyJJSdqbCzbf/SfUPnRNAFPvLh4Z
wCpKAZfudL5FVivdrg1huxGO1bRVkHRDH4HVjLn34YkCaGlUJHU6P2TuTgCsu54s
aBMnmtlNt+ulh0w//Y0s705aaG+9byvwZgalc4NQpDM093UYT9npwWwcKrCyKxro
HbkA6OwuWD1LEOZVm5QCrvdpp3hnp+AOZHoBBGBXb6Laou7Huav6PqiAz21MjNmM
38k8n+IhYoE4ELwOWN0g83mMam3rKyITmJzLnkKuCJG6goAd9H0Uovo0LImlV+mH
PJsd3SSiJ8WoP5EIhjCZMMGfdHA8tvrAuJI2DRNLCfntlqHC0t/zSY4N/AuF81/L
rKfEeQMEboTkjGDUBKQ0dzI5E1lA7JTnFJmdxBONhAaD4Pvmy+Z2gfxnANV7OA5j
V0OwLTxhsO7oiPvLfP87cwIV05XAZ41rsP+z85zdvD9X5LR2ZLSAphD+0eWZU1hv
67BiNgH+WsZrg/lCDTIO/XLnt68cWEyGpbvFtvZX0z9d4kU8pw/OCnT2TS9cGvia
3x1D5TniXU1gNGGfcB0YbjRxaqXmsJPjbOHKlO8Or1SGCo9R2MR4dhUZMhJYbBqh
O/6+Ry1QjsT8yLxkbYKbtIR/vm1BVQbERmWX4dAAvzo4s0EEgu/ln3G1bpX9krUk
dmVS32hvSvdgoHWt1Cja0+AXWZDNs3aZVVVq0FsRkgPLetAB5GW0++mZflms3wDL
g9nhG4MbsetCy9sRs79tU7axFrGE6esEH0B9VciMk0xBP6bdrISdOrJgtVnOey3o
deR7rwK0m+u/5W9/xZ/oXBo8y5UMtvxIYqU6uDtvyAjUNgsGrMtvip80cUjn9rhG
36jHgbQwfejJfQb/XZiPSSr6rHgTt2jyAkN/6La7CsLcLDgz15w/HzXFCVn2IPwv
wWNxxmBhZa8a8E3VPJkJeZ3x3AE3BKKBR4tuPvkZoW62mE07O1qIxg6LEb3g+xQE
F5Oo8S+f9vVOGP4Lm2C24GHSZZ0F/e36uuKBYWuHsoF2GW4sABLSoT/bvYv3g8o0
PaL+ny4jZSe0zWMz5mdytnvEnRKCuzHVnsbEyGhiemZUcL+igBMX5QsjqcPSlDFU
frjImMm7764oN3tlWs5zfDuFOVA7jnIfj5zWT5CXB9iGEpjWbYe/fBDIU+2hTAEi
jtDiQga22kuzi+uOgJzxfrMvCvlBtoXdbo5zTEPN+tqPoPEJveme0nLFZZTpM5vW
3yFOTVzGlkvSuq1eiQPqn5zh4T5G50FYkEMFzZfDBQ51U9G2WFPy8cvpyoQzvH7W
Su/9t1tr+NLO4f0hTQh98EstMPqhqCUtvLXu/pUI0KLUqE2BbK113dLTDiUfdqvQ
x4uzxec6KGnxBCC4VW9GGNZzLHV+NXvhvoV+tzrjJ0nlHMzVSFXEvUelssB71E9c
cjxaeGl3GM6puiC5l2+mQohEqdZroaoF8O+CWcLC2U44McZ85OSYOxFmZ5CmO0CM
XGCc9aK6J88ftFbssX5rg9xE6TFSkiaf/eWjmNwL7UGiU6+nMVVnJJlqW610mm9Y
w9cz3TRmL9/NlTya6sJQ8X7LEE5JBdIZ48RRPuNLpNQOnlBbior98OIdg0VE8RKW
FT3OJg5i5+ZlA3l4lwhQEU+Nqa/Yilb7R0hilj5c4TCr7YM4IEa5dMoSSVXiqJLS
c439sPr9YjIZSlljzjmYxaZPCwymA0rh+H0k3Ij4l0NZnv0n9O1mNrDFgjrXk8vo
aflUpswngqkImbHEVBNP6WiAXtlROW5owV/5pgayKQYM151+GIh4i1vHgxM3hikM
L4TQ+r9zihJJAHS9yV5lGyJYdI7KxfllvoAUZTOWqV432pg0J5AfJfsJVPHFoEOk
ROoO3TBy0ZhdEyWoruKQVp+0m2N5DnhpQ1FwdSyMymHnkoUNpZH/ECZ+zkiZvPfN
zIvVSNtHMyVmQzbCM+Js2kC1U4D/5TEwSf2Ezrh4oSiO/F2+aJiRN4XLELl9lqbm
cM+jKrkm2VEdIw495QQTUs6Aq1bwrY/pZFSsEa48SjyqlvZ/jm8836UTVX4j0w3U
dj03EMyDQEtmCNI5K6t3Tq8jpi4iIaUlW/27qDQJDI9Z59laI/3Zc2sVIQYwN3QH
k90SrauY1orx178tAdrwNhRKmnv6ODekcMXsrbC4lVpmhU58sfI7pUOeg4MeRZ/v
C1pJDlQ5neGlYhgEEEMuONU7qaz0nzv7Pe6mjsfgMdlNBE0EWDxbujyTmBW5j8T1
nA0ZrUi1QM6bbD1UCtI+fR1pgyAGflfmfZIoTG9vrCsCiZdfL+f+CiwmLHJp1P69
yRUKJq/EXqFrDBD2fIz7ZGw3EgCIZ9V+SBsPtXiZqmJCT9Devl9AC+BdDEYfkFN/
y+eImWtCo+YgIIjTuP0rWOQ7RXFUmQDn/5q24RaYYBl4ZQrCevxKN71S7BcrqvSf
72PPRUoQSG/xKCuNU6IEu6fjS30OYHGuq0/1+r7LE6cvfs8tIlloTj0NjRBY3319
MHuL+8HC3J+Es552jbjYCOY0Kkw/p7LtQKAFIGzkH5j4/7F5GP2PNas5Nq9vXkXq
xytXnO9lF+83JgXzOYof+MOvekYya1Eolu4xO+QZ+tWMoMEAK/jNTuBJAdBgyRcr
stftN0uTnO8NDlS0Mc5zDoDNXLbKIch1ICQV/7wJHU9PuJG/jQq1EkLyK5Cu3BAt
TNF1txcW0pooxVWKi+C6TquekyUVZ80DJDdmFJeBudU9IRB913PakXXjeiDLbwtu
sJHwhWIhLWLAo2UssJw9DCE7sYn0DZEGtJbcy88lqCNGzn0yO826Gfs0d2z5Rgnm
1SMRjuM8KbHEBiSKmWrq71i7A4w/KxdSwjxS+VUCgpmnQC6dxMbTY7H7NpsXXfup
Bmr6LcfWN1z9H0KgMmNSZM06NV3nBPTAn6a+FSahib8C1acH4NaHUnPiaOS0gPQQ
2oS3qQYydX2ijWP4Agm8dySaveSYfnRb+N3pq2rBbJho0NPUqOdGDJZSqbw8jVeU
I8v8hwzS7tUYkEOLJMCnzvXDfYbmS0B3NKu/lfHgfXESVipNLG7pO/LhoP4cQZtK
4pj5JVNZ+r679gUY1GH77rVU700th8cFPRKWaqMRc4NOswFK5sTNgtiWan7W+q06
0wMfZZI4ZgYk1d2KEXCinFztuKjMdpn/QGJriADZoE3Hw8Gm5ONGMB/ntoDPY81u
pK83RaBaUQCX/6T26U88k3fnL++tQ2ccbydEY2mr/6WGL15lJb4hBcpIZr+cAcaY
9/D7c1S9CE2ChXSbtWPsM8CnhQ1EDUkbjcKVxrSus/m+w4d5cHgJ1bmaqkRsgXUE
TjHdUwmOOOy1XvK6EMdoBLW2WF/kGqH0xqLUf/GsxZGbdczHl1QKCRK4s+XYDBDV
xtYJVZGU/JfbuME3dIde5g6VnnNdwAfZxZ4LdilBwvoT3h0QNFQg+yqcY3tZnFO3
GMz7sn6mH+48jWv3dMl6C75jEcHqr+ubzce+tsa72YyfnVGx/FShqOxkQml/1iGi
jYFb32XB7svMc6E1qlgcVbipKhoDrVhFkn8VKsWyPS1E9nfquX5+RkoIQA5wh1xL
6Ua3TusqgtsJyjB5quTpADEQwSAk0Bg0fhhTZ98w68yHQUkWwTv7wmfUfUzUQra4
JZymmo1+BmiMUcND8WcijHl9T0PxoSht/C/PfQNrBhQ7MwX80jTYvflzT/Lwp0BA
2diYfhOm8p5MJ1vng7tCMMJjbVD+TBNdLv22tf2r5CY8w4p3oNcybeIsseRhCDg3
oRpg/7N3CCTA8j/HtUpzDciIc15xlCQQj+lDRg6BcO6sp+vIybGBrZc7C8RVLZ3H
/NoWLBhiNS4AJHgT1svSRQ7dyCKKPU7ThFxPxBhH8PIsx8dKCmsOW9+Vzj0GhgXA
uNkny3f49Y1W16bRT+0VmStLKbLOXBreoek7IjfhpCnXOKdK7UpxxxtoO5H/2r46
VHv2r9IcO8MPNyZ06p/zvtuAxuCB/QCPE8dUuEMxNJVNpWWy9zZmKzAyQSQe41PA
BUQ9Yjsdw+majxsnOmQUq9g4Hr8bSwpUvf+7yxYVDOELS02kOqi1WuhbcZFFZt5q
NvKzyHsFM8IRO+QU400lnkFZKdB92rOX08+u5I0RiIWdmmW7LqBNwj7UpJHkoSlh
w34FWWXJq3b9jFB095ovT/Y3FOMukyk+4FcsT10GkeS26s9HKLlwjjOvChYdWVoT
MjM2Jm1NlO3zQUuiiTW9i0WK0f0kSo79arUm/p3/x1oZaZBySmHOSJi7EFoDH18U
Vb40UxjU2o/STNGuzVJLUIz3QJtINazWXzWPFirfw3FLB4kfR+rXzqh4qeMnUzMt
jY7WbgYFhoh2xaSazb3aaa5UceJrlKNXzMEC8x3O9jOmRI716BPWbBBYWL9ATfel
hdvuO5KyW9uuRXRezDfqBdO9XEjVrqDnSuW49/HRRHFlDgfZXxxnSNhAeb85bWKM
uDsnIWb6YxYXKV8ON2OMH6bFz4PbttQ4tcIPccfyEgtQA1Av1WutCp03CVlUcd+j
7uTZxCZ7VofyhixArwBAGxlAMTXY0Du0fMpNHKp5rmQ9Ovvv4lk+BjO1s+ICm7cW
AXrtoXdgGXSxDZbUUX/x30ikHeshqbjnnIqqiGC+gltOpfHakQEg52xkkjus+xWv
kUUN9kEYuyTzDM2bY5udVyMg5vL5Efh7FG9cAgAvRtk/E51r3GFTOu8j2elbNBSx
40869b7SGid3KAObmXbU6GF7a7PqGEZqeH9q5QuIRt/v1U/juCqYgdC06oeHjvPr
A5WvMwBXW5xjWzn1vp7+f0MCeBYGXm554Wk4cHPUeBVpfBC4KWd6VposkbGTMd0W
t9aQO/gCBHup/+Oo9FggGohAXu7Swr5b/tygyr1nKuuuv1i1sUGFEjw1lWSi+TlS
iLKzfbVnplaiNBGFkZAj+iqFyKQo35rrd68CzhHASgdbx/RivCpFTjKWJmjQTg5j
tjxSqr4XRaXyshmDY1V0P5gut1y2XBnZm6dd2ihXYevoF8CwBZwlnHaC5TYGPqD1
DG6jLvmz3jMqVe0NecJJt4uiRCymbzfD5YhZMu75tGc++68Mr+espMmtdtO1+ipQ
HHyvSfr64h26pApdnlcllJ53m+z4wmEDObeftJeD7KyW7b0LHeV9yIWM244/DVdd
VpuMp2gUrPOT/2/0G8l6c7ATIDvBRi+PByxwhfJYT7G36IwWGSKk1GXr3k4h2Nca
HV8FPeoVw0M/vV1N+v6QC1v4g73ZC3yBBxHpBbigK/jfdDTdsw0dLCWQwzxvhOS0
QqTZwn59UUX1lzVHWjNW5RUBTcAUH7vjhj2UDGlNEHFmvjQnEHop56sliyW7JCoD
Dpo4nPhHHMymM2cxhijx1Vw/DLgEZ3OP3gqjw3NpE1Uhu1zIFLkMOOkU4NCbZI9m
dfGQZzgn9xxJCClPvxxW3JEi2fWlp+kS8OQ4IPj4QLE8/PKItUcDbJrttk6jKj/p
8Uz0oQv6tlOG8EW74bkkwcw7j7zTTtXQgd/zQIBb6VK7cbwJK0NteorQn7Ix0OpT
nOqMCtKLzMpIatO9vX6W9J3+lSF9gxmm+0qRyZ9us9O/GtnqbcYpLyRwg/KM7VWp
bTegNR+QNCXTaZGD7KGhCh42ILuApjbe0h3+zFWa+O02t354YRjgmAtQzZLCbgrw
vxI6QYKAadnPZvzqyUnB80TDyuavbmUAmAtk9Qlv60tiWVUunkvTgbp3bIKS4NMC
VIS4kklUblykNmqPukmfuEr2eTxxrOmaZJGtu38KT729usZNYzirHTUzAD+BF+Iq
nk2DOsIfBk34lN6Qgi4uGUnc9DmnummUMOg6ki2ffL8o5MfRTFQki1ODZrYq+VA8
BkYinQkgFlBMtqrtti0A+lTKagYVQjdkqHf8hHg4xidlpq0ym0j0UHviU9oMKbsE
9pL72wvqeBJa7P/okA++9YP2Sajubhqe2oiHDSJDLx8IrBtsuXrTPuY4ECcQeRQM
0x/p6qXWHDk1dgqFA7yvpfYJWbk3+6OvNokG99EfIHnOh67M04pMSTUQHiVuuXg+
RKuzoQ8Ti7UIWZ4P9Aob68U9zFNT4VgfOnxpJ2SIpxQ8Y3pyK/2t3JsK2ftBw9fA
P0+QIDqkyi9IhlcXUB3wGdB0LbHsAJMURtjFBMVQKc1/kCJ4VKqeL0wys1Hsy7YE
TTchkdyKKIrOoX8XVi+xRXKXb7prZcrZFYV5ps1W0yrkIB9jeTIXyRSaW/F7CeQA
RjHbjfLB2oB39Ks+nXb1OIh0n2qq/fRpUfVykMGmLwVBTtUvocq+7S21BfhBioUM
O/4VvD/Zp3UW9mmVSl4b+ExkkUYkfJxt4+8TxdhtwvNYmGcmskG0soEiRbsgG6Qk
zNMdo1HrDCThi+6AGAKqqXKHg2YfEc+W5ziDE1SRGLaPJ1eQg0xZ/NVesjIM46aG
U4QOyrpSJnk+6RgpKWL+vZlwjLQ8AnDXXfFipKl4lTMv0wMkTfqh/h1mzi8uD41e
J28uOJDWvJ3Mh9p+l8oo5Iq7w0udL0uQrDWYa6XXsX+TGimW+n04V5IDJ/HcbTbv
Dq51GZNpZLgvQA7kF/1/3OflENL+jh/wETypYfMcKDlkr9TBhws6A4Wg/jErkbsx
5pXiYoxu5V3uUyFJ3acrYcI2vRFcdUOmDQDcRkDiiQqtNnlWMFtRhrGDmpOt/Gi9
rWkztVTluWBuZ++biwmti4Ga8UpItVUxcvouCVXRjyXOUphhrA5kNeS1rvRahBVK
1/nnYzW/uT9zWC8Vb7kQQkvzkBZdhR/FeZyIQGVTNsS/uBxwtNGXcssSkwNd1An0
cQ10pEmtmnDXHA0dsIA2kXvndeAfMsTyOCfv7yUV3+PJAxQGY6y0NPyfRqYDwMyL
f0wQXBYJk413rMgLqSa6Ic6SEor2oJ7WuaQ8iUlVwcYWDE0vwQX6XOHGZonESrN0
QP5HFC4XjNS95WokhKkevq9aur7HhP+uixxIXp06v8s2p719euDktNIyV8UoI2hL
4RtIa368cEBqGvqJO0NoR4Zs1sPcDagQxZDFbKAzsdUZ1XyLI0i9fr7BgyG4N+J3
rdacz+9dv3UNNxTCvLVAqMwH6+fF64TTkykh19zC2cd+m0MDNm3T25mUo6XOWVC7
0XZXEMZ5nemHuwNjA2PgkIAUR52FMJ4a9Bn87DG5F/unyWEL24uAZ4enwov5Bsm+
hFayHRAUc700buEOhxc/Zf4CuL11T98riW8h3niI+XPxjAE7u1uktndi41Pd2/Da
BCSjdPtRPvzSQ4N6OEMnt/ir0HP9INi6haoTFPDG75gwBeNwjmS6IK6D63pnMy/7
qkSilxhI3EgdjHVwVK5OeVFHy/SeZT3e5+2mL+kYONiIth2c7C5eDeaaxGIVvtm/
gHFXsGyr3tGNckIqqubvyeMW9W8Z0myL7QxVOL1ofEjf0+enAu8pmeixqZJcqDkd
o5oxGh+FQ9m2DJgmixeAcrxmKMMvzpSfPqgPKFFOhb8trZ8gSqOu0C4goMFPhksZ
8fJCrzOm3VJK16mnGtGaAKnvU075MWrICrE1t8aWqkLR1k9RzelGwViwOL+5Ht/1
m/Nmj1mvhESltgxElF6ATLb36pfjYPVtA/a32K+QTdFpD/laSch8HNq7ZO7RqhQp
VMJRbLD63LvRDzySKqIk2pblI3klAtXJtNzxr5MLzBOcZPzZNW/nv2KWsN8p64qK
J2tO1Irb3l2qn+z8KqY7nPP6jIl7KEvX4kZRLj683T1Gayfp+aShAFxsumwHawPS
kR8oPV4IcQ7OhZw0PzkzGSNStX7v7ljytIcznqWxCPkFieHgOaXfRwoZ+DHOee22
tRoYZxEAVmqQgwvTSKM+Rv0xJNlpg6SC2cdN765H5m3Lo+pT50tyfTd0L+IwZLDR
PMoRILkYw5KmQ3w0QnivshSneo4DzRMFdbUT+e+3bDYdxkSdDnOdXY/5qn/vzypd
mKeeYXSuaHPQC66bC5dDST0QMlHULQcXkqU527EWWEGE27SCkzljR1gdN5KSiRTG
5sm8n2i5yLrYmekhTvB4Y613qC9BgjlcGWBHYwWgjEi5ZUksFJNmZLn6/95cfuhi
nwvo7PYDBMVKr381zzbG1tkybcMqr769nqfREL8T/ZLhhKN0b3HGSpWOV4Yussl/
EPx3pqQg72srPD+6I/s+R4uP2XRDOYTMqXvlyLTil8PJdlzTrsTIEjrcd45KE/Ds
Io+yX+4eOLaeE4gM2PrQd6I9OkFXldpezRySd5K6i9RbgsPNlSYaal5PrBJpYe0S
NbvBvCHbGfuuGzVfHmAwkXFc+64L2q2CikpKMoHzhwsxqluJWH/MYoHdi5zKO+O9
BZNLEJW5oX0ethXaeB8B1ilvyIMQvcwQIuNgiQ5WbDNcPJSijHmByEw7HI2UVODD
VOMWpF107RPweywRE+luP1MnOugV45Zjl2XnWeBv36JD5BM/QD1imUMqBiqFYJ4k
j9cv0HDx4yU4aZmCJg2gUt+h/BInKkN/DQmRNx35BA46bbfF8bzWU67IHkxOymQn
oR9EUv96or2mvEruejXD6DfKFiBhKnLQkDB1fTIe9q75uWoIeUVnXurAd3qwZm0l
7kYutJqE1Nffsv/Z1K0e4ixhbhzwoXYH1pyP6Zcd+ep9xeCw9+CHfQPjcSjOxE8g
8ugznATmuydUUgSZMRWBOnv1etD0B9Kmn/Kr++N7MpbuIB5MfFsaIFjYkJLumuZ0
yZ/LwmJYxFq4cKotQ0WWXnsUZQQJ4LOgLWdnBU7QbHXMNfUmt+ohusU3uVF39e+F
EfiC93IJ1zuZNE2sEDqSrYQlSy9WWnnd2XEk0Pe/sOSh0NU8WKBWyVrXdT+M1SF7
EScyUEVCm21KjEr2H5w97Qvlh//FooCBi56z4CXjrauSIDLOsfsWtRYbXGgtnjAY
CvEoUvM07xU/v3YL9PzRmWTzOGTwkShd8vAAGz0wEUbZXlWMd0aY6oAWCpbgnPvV
qW+k+OvM4dNdJ8L6YUcE4d2w451J0RNZCWi/AJC68TQR9q7KnDF7BknNLWBhnF7U
xMux54rHBWQvyvCJfw15wsX+D8akDSb2a+zhuc9R7aANtdGzmdV05X+ayyMUWr+x
o8aKvW8mYE6Iw/bMgREXOViC0S2BxeUKIDKDVAPsso4P8xySQAEjXW4E479O7yfK
NK9Ss/WIXx4FLrr9/PXkHlbk5DZRDXrLAYImTapHnIHQ0rAlgcvAMlfEbT0KJz+6
ClwTogLG6Qo2FspMjzJB/3MFLKTuKi3akA+/6tbrWCWGmcmhEEA8bY39NFCQRRO5
5uPIy3/zJzTci+v/lIB6oMXMmki9hojxnN0A9ML3zUAe0SdwY78p577DPh0DVs0t
b1/+iFPVcsNfuMzylF3LCU0L0UB5XlVyU5I0L7ASjHp+rsDVIJmnyQYh+ojKkSFQ
lcs+X79JGqF5DPODNOZHdCl0xD0vDecJETXX9DZ8+XACQqeiUlJE7gPVzYD6Q7ly
2jGM6MApte77E8FcKjZz/HxRJJGancKeNLM1pNjxbJPeoq3AX9U0JKQdFhGm+Zk2
2bHctxthKglTDZJaYOUKTO77qZW/lOkwvRB/Zq79+KpqRvoyGbEsHmQJoiJHUSwS
j8ARHNUYO8Td2JC5uiBexb3DkZzbhfmpbuz/X1gbNVx3FDkXtCcpd0HzmXP7y9mY
V1k3UWwzA657i3OMvljHl2gxxKB7RNbdiyylhqRuqrcuwbOoK2ZQhlPVWjCmimFP
AQfQutCjrQuboXGu1gUSDmzJzZIc2wrqhBomx7HfPsbjmnQl9SZePoRPoMrBF6ZS
xyUC+BR0Od2dz0tr9az7a/xir329Ur1CJfOGhzVDq3n7b7fUHUw3pPIUEJE1IRi0
KR/YsiSYSD366Od+n6bPSW5ksW3cJQJ+rqcQ2d+/Lq9wphS0OsMIfrn816ztyEPo
JPztEXAtqvymta+cj1mNG+l/ZLrrUyZlzi7vFQTofO6/KdpAVTX7EDujzWU9E33A
aoDmj7/P37tqFZYS1c+SRcW2unXuUwWMY/UmQmmzdENQYyfX5R7+dQ6I+Y7gqkLD
cTp/PGRVJpedRsAwQh5VKiM7+6Bm2reuKnPZ3+h+PSut5mn6jp3kkd/RgB7PEUjc
dNyN/zvk7YbAZ75URyaRLWonDKZXPt+wraENRskmvvdvS4l71djvAZilCp8LqHiW
bUfLNk9e7LCqR+gZicCLy34DqNMIpRqlx8cTkqbyPzDamqrnM5sBPg1T71/Gr1Ds
VWrAUHE395SnFd1x6Ld+GEraBILToVh1zUUnv5v1jqYALPRaUIbo44piHVUwr3aQ
fCDegYGJFdjVOQ/96Fd7MTyRhkMjMJiJsdrtW1EeLTGV4zNVj5aDUs8teuL8C5/f
O3TYPp+lHA9IPlko1LXAjgI/riEqZ6ErywzDRqOOaX+PI3pLLFlXwbaP4t+W1Bz3
WwdgSAl1pzULiIrWll9XPFA+uoo2UkyG5bMh03i+ybvlez2I5xo2O2vhoVUOftZf
jcL/CdEAShRgi/z23+4HyJ/E7Kodb79eBmbGbTUt6P+59+qhglHy1LjPRp/dISdF
xk5JqxC/jUemin1LNz26iQyfizbcq4UnIRZAg3dEU9gixclBNMN14Gm/gN55F1rH
LjxwKJE3e5wzNQTSnPaJ7YtxdC2TUK5s9lzTMAYIVcaKVK2U88vcRPimeMGCLlhi
HHIHgHOyXdwYHLBenZS4Am5cHFecx61VcPcZBuBt1rQlieci2uEgjdkITA0p61W6
TlkBf2wBQjGZdzNHj68OTXvIe2gVSXWSfwATE5kZ9/etRGA6AI3aIcnkeBjRPmDq
9sBr0tfsk5lYmamz8v8A9KnS63TvVOfnSHZznUl8y58omK5T5fLH5EIKmaH6Z3Sl
IM5XXTWk9rUtLFU4Gtac1R8HJavGWhSgorHH7swZ9JnoxDYyFUSB3Pvb9Z/EM521
n3vz1zwHUM/SNmu2Tv+gl7JI0e2l/Zr6FT+qTL0H/i8mg6it3NCOaNHHMHRquuR9
WrUqU8CaldpfgOyKZDSfR9eAU4lRUVvJUsuw9SSl2/jg37nKynDT6VgXZkFY+ZHC
J4S0FkuZFPf/VzXJ81W99lbmt01bDFw/lv64Wf4lu92pFznwXvugxgFlwzNPRvku
S/dAzi1Y0PO6Lcm2Q+ExBfoHI1geev7goo6z98d8agLQQvAWHmJl7QFK80+qZHZi
WtASZKZL7u7fedDI0KR8w7aLa3oNh99SnRfbi1xHaGwsXt3sz5uUV616a2w5EKZt
jIKB5CVeLfxyxx2vrR7lAh/4QHzVCxrdsv/iFiWxhKn+65OTp8MKqp2w6YlrVRdM
KWDSPvN/x+iTeSAZyM1sjEd8haHPtw89uSWSvHhJaaPxJ8firVvN+fSlHsIvmFI1
zBqG0k7zr+TTW8paII9PM8pUVtU+4OvIOFfRkLTISi3qcMw07YMmVXeAnU7KDHSW
uAVhcRrWgfF0wWVV9ZO8NutNOZc+gf8EJ/j8xcCQVwYtmx7en5bbNdOu2qUamyRV
KYp1ZKuuZfpHmgFTxLOab6FKRyqi/81AxIdSNRp8kUP50ZrvVIf6mBzL/SkEczk4
ldj6Vh2S5RT7ndZTWmv8ZsQDqgHxC8A4EQo4JBetO0FvzRHI7UKxe+LFD7+wdzmW
KOpDmJaImb7VzOrCEGzZDaXApGcUYyEzZ/DGkWujditnHTLGA95mH9HpAtLrSJAn
r3dCMWF+N9f9QOn4buWpXA/IWWsKmxEHqBLE87x1yTm0GLFD1AimBbZptI/2EPYn
Fk8skPagabGORj1c3/5pizLtHLUsxU7/gGTVRrW9xGxPS9vGaTBJVqsvOCw3MjTM
wMIvzieqRlh4qgwWXMx/tH6NFhWudRJuTdvko9CYI3vEkq0PRYEHxSXAdHe7oJ5T
6G4bX1umvh4acINS0CL6q5TidtvC79suL/8qF6RezP1ciWp+YuexyZjxnNa+pJQG
yvR1XYhNxYAm2lvFmj1BiYwYj83/+OGhX2K6+SVQ6UU3HTptyRv7UPT0fgcSPibp
q/mc6q8mOJo7mXBRfs/f+IdLNwLBu43grJ9evOlBRlmMU0QSxRT9QM7nY2KqGGpK
p65csUViNFoL+7xVzLLSfO6dSyktLUamN1w8mEoNQGDBXfw3iGP+neoWZkBuo0tn
IPqnGog/yNI2b9pe43jYb6KkT1PY8EMeF4oMeGW7Xc44xGmT+nTADLtNplPknUop
tgnsHVdn3Iyy5j76KuyziRp+e7UCK9+rLBY0KhcUWHxqO/yG0lZfc0xt4kmejvVb
4DWSivVfRaXC77qJQ5k1FEKxl6oOqv488e456uLgPwCEMuvXQz/4HT7wu55ITNVP
/ROZzopMcejUk6/dEJ8JlkSmn8QO809lNn3Uw0OdIHBSFrFxNfFj0xdZWwA8cXeK
f2nsDfN3cEf2Ozx3qtzI/2PBUi/J8er1v6CX6KPzYM9S3iD6jhKnE/SLX0XHKuUI
FNATcfW2PRrFMMCImxMlV+OIgs8lggJTmCgbYfbszx2H9GkrFz7nB4VXY44f9sUP
N1fTvfPxijNGfgvw0o/nXwDFsNurMpr56zO2MCMwPe51jBmgGkQ93WJT9tcNoaaC
Tkxtzfps4yA+aJOxgChtRZyPRAY+EfP3Rg62nPGs5unrC4UwK+Qcqj3i7WwiRQot
M3bWvWFlCESp1DzERcel946RtcYkqdzovBR6HzOB5tYfHkpPxpeVAa0IxeP/Qhos
EEcIGKSHbfudFZXR43a8GuZVrev6KiQiEVHVaGgN2oBc+qoKHu/zLV0JTZPJq9A+
rb0rDlCOD3Isvv2WUdQCb1//Fz7rNmC90lYNEtiKeGRZzFL9UUDAoC8azyBdfDYb
+G20hLdiSl4YbB9+J+UWXCGOpNgMIvwkF9iXB9xfYA6EcHaZpBbj35GXjHu18EC1
qDn1uydCkQGeeFtZzenTOiMpfT+JjtRwcPnoev1nB6LOlT0jXNzSO3AtioT5ryoj
CKPK8mk2wM5U9FoD6/qKCtHjHT3vxYq8Fx686aTtCOFXk6BhXcY/VlKsvO+jX/1P
tyJroQN+Ct3TmXWoCtSPJhS20CaCvaurciH7JABJnXK2WtUoaPFWGbRMENooDkDb
WY1J5bEBhu0WEpZgCafo0heDIDk2QvvMgePhrNKXOeaO9EJOcD9TRivD43wgiir3
ZRnJI3niXqSIKvz97cwLw6umFb3+XPji2uV9/faUXdFqIu+Wb6zZSbX3s0q6tRhG
yjxY2LUwn+HuzdIqZ75SJn8/o0IrKI0Jy3gbe3DXrCZD/Vp5gGJz6XZ0pA9Wdud/
8AyNrSNK+ly5i6PfitypIT3USnRUdaQlMLBU4pxoHJsIjDcJiD7U4H3JB4Lkzm/D
x6k3RagroO/jzh4Js2bS88QgccbNtWl48lw57izGI2lhqAPIRIU/aV9BKJP6wUZ3
Vgq3S//FTNNQYQdYWAr3xj02I27fbhoyyygDPpuc0AtFcXzeQRgxpQP0vJdl/av8
DKI/99KdDZUGjYnPVEybTi6Or/wj8kJhyhiDbJoXMPZA0LyKuG2V3cj27rwJI7Ka
FCSpidGdCZOXywAy4R9r+m2SsG0Fdqcqs23mZI8aZHsae36dMSciuElfO3u8nFd7
UtXFi5GbRFBHQ6sQf6wLAJDs4fPTfxu8TBTF+fDwIpj1SNzDMhJnp02VyP1Z1oBm
dYP+luaAtNe3iCu/eNYZbi5LmhlFHcYWpFNeJ5dV58k+6pepeMTGqpGQ5zIQx9Bb
dSzRF7SG/IdkY5tgYMuhtYzrN19qz4GexnWI95K+qvKrdTnJcq6ZYfQDQIX0hpft
tszj2O/0LBDwAOkteb8GttzROFcNDHtBNC8cS8/mNTtQyhEW99vILQCrpT0JzpWM
syfMKTgAFM6Ql321ioYPCfhPAwRHcZMjZ027g3vCaiKcT0O9wveLFeSsOg7ukgwQ
hNjYqeec1w/QttuDzYtZFcqRJtYJQOwTLgp8Lyi/9XlTemsTfb4HRtkBO7gSsDjb
3CTentlCBHKcg3V0f2Lud3d8htN88HXNy8GMhdv9mNzkKiBXA6k0SH5E0hxGWNcG
runsaQN/izpVYfTjbS3hsAURP4xQkmGGGQira/HhOYQ7kJv+xsAfQy/QQxfP/diN
LDdTkqmEb93FcsovZNXT3+TTLt1CBiYT8p3Bzqb7jgAi8J4jC9T7Gq7GtULpZjNo
JwAHFWCcA8/dajUwx8cU5DVdb7sEj9BldjyZegS7IhIa3/9++rOwsPA9LMRAYWGR
bOfj/EKz20haujsHsWeJcvCBSbtEMNmBnSOOz5PFKOxTP4K0wWgxosByTo6FsP5k
i8IFHlBCwwNL8Eu6u7IOVdHWwbMxCDqGvaxpPj/6hXyA6Qqhs5Ty3BF0qkjwqdks
BkooWn2vRTY2VndEdWn05Owgo6Z/rfndi1KpWE+OF0K30OfjScmud5JboYv9Zpxw
lk/BkGnWDTzeHwdf0AUtZ02itb5G7qTw5gBCfROx1cR4OZ6eOE4QOah/t0UjlnWo
sSMddpKCjAjprWCmqJ/FAn7QxgrZ4yFh8FaE8BvnaFQre9Duhd8wbCCuL6s5Q7L0
e7u1lrMVH3IMJBDbnGdgytwa2JIP+zqYYIc7ucIRB36MxYxhljTtXgeY6ND4h/dK
cRnr5fsMfnXPaTBCS/4uB/umttp9GYnMYqZntWa3PRXWMNV2umObTtqphgE4bWKx
mYAmmVWXeh0tt0hvJAcWhM31sj0bZrQAaoH0jjEPF9/GYbuJ9bF7xhuiHwxSHGP/
9TA/29yccqd5WZA7GcCfmcoPhxXzzLYM1Sg57nqs9PCkFy0YG0ZJ3ruVeUy/Zj3u
AH8KhvonG3Phv646jCDyLV3o5VX2NQTijtXHLFciBjjc8wBdEYDqKsFGOktL1lJM
rmPBg6eN/WEiMtrHXSreQXZ7PmEC/8A9aCYgfY5XxALA0MUffJzVt8TqPxHWfDiM
vD7/qFL4c+9j2OujgLZz75wvRyZAAmbmNZdpkon68ryn2L1/Xqn8+V4lXEMTmOe/
oYuLB/jSLhDndCcAIdomlTLCh3oV12DvX4+y4I3U+G0qAyD1sNl276r4X3u1C0mQ
fmJQfWwxjFE8XMemqt/es9qgZaCIzmiMJDPAJR9amzPoptflVqTXBSKA1+NCMSXg
UnD5VwIl4Q5bDcGKMaE7w7QQUl6OhtJJYH3yCtRBiWSPpLrMNQsr+19Kc17Dnxmw
pEgIZ8PlT0tt9/15oawRXeggSkm3vAPEXVOwJrYuiNbxN/kqaRsosO4JCVIOnyfD
sWfRkgQMB9psGjFwgDHon0XfxFcx5q5XlvPP1eJYUvZ1idiqIQKgWwXp+kHCPy8I
EBtw6h+egKr1b51ZTlHu5femCXqQwVXLwFgENt2yP7YRGa8Hu/8XzIsUN4cJfmoF
Cji/cMJkNOq3i5ziPIxDjj9tpCKMht987XHY1CtubOXAjnqBPTOhSS7RZOddfHg3
ikxhK5jU2RbxX7jZz/NGqAOJNm87xm87zy5dX+aP62sIT3IHvILWCirxG5d936Vu
LgOI+OPyupPoFkDr6dNW8wzf9zaDHQyqDJyaKs7nuNBMSuzLOYyeejFhd1ouaNdm
yr3lD2B7pnbRCyqyllFOkI8Nph01rai5HYIKXbDv1wm3qEbupRgo+dySZq9Z9uIT
Tg8d5riWF/qVaF0zr1EesZPq2CToni70LJthZc0gpqQJbmrPpIG0coTqePCsdXTZ
4tAdZBa3zvs7NqTUWBmAYRzjv3iiQ7cXAU4pEk+pSZ5UudYItYE2gMkxqJv0InrY
GPaXXtgra2K3VfCu3o/+9FjsI6kn8xSmEgF7uXaCyTmlOWmdGjbfr5LH4reFRyWK
LYql5BXtNI1zO1yOGSIKitbuzd4BaEsh23Arsd8fVYtnFfNF99bK9yxBEk4E7/dJ
XfZkopjRF6Qe1iWEa+4L2vlXINsju8DC2X639ZtiVZRpiLvlm4Q+ngdXNq5XDAW2
140EYn7RPJ2XWUO0XZmi57znh29vsrGCmJEpDbvjbd9jvPYvurqa6nrCQrdOP/eh
9g3Hzyj86UwtaDE9nZWvuh5+ZufqGN4y7sjuRiydRS3/U9SVIaYI9hh/ezggkdU/
Oi5ZpKNKHbOQRPKa8PoFTmba8mj5WwrNPQ+U4+Qx2ENDF7PA7s21oh6PmuekD6u/
q/pMB38qk5t6ioHcujBmvCxqlo+wcFgUJE+MnjlyFz86KOJDHPXEQ7ErsVBU74Up
6J1OiZFSY/P5MIsoV//vYIy1fv1MwW7dmye+e1SAjI/3ZPDEswQwNHSOl6lk1G+F
z2ghPq7tx5+/CVjEmQdO4ETOv34jYTZVbBXyW/PWKQbg9W/nJcGcChCty9f2poE2
sJYftLJ05I6VDypNUuCXcSISl17/eH0sQTni6iJXDImfHrJefMVmXyXgIlqOOe0g
uPxEhKIMxL1qXpeiEwmjZ/qnafyQ+XnWyIfrii9hqSt79Gr97gGYw78ZphQVEuMn
yU69IQtKqk4ORgTDdIZ4Hn9bKxFR5V+bnbQh7dy+RPD6s1/VL4NbYZbJTlH6Qppc
hlXk9jEyusiff56ED6bWi4osa1LVzZCV9khpo8DRRy0oDtUFLOblYZW8Ekvc+vM9
WZrbMj5TVAN3gALsEVamQAwtd9rgxB7kaiwPkSahamk5DBHeE1IHMCSqVDXP/7mc
SrhhHfMRhmeJBujfV0OUcMahoEGgqd9vyxfMygZF8Wm1J42qE42do9QUTupysV9W
G2nicjpv6Z6o04yvSGK47NTX/W87G/527+S9pZrYbaCgUzMtzteQUxE4WFXrnKEu
GaZOwAc6l5npCKKNy18Jpq6KsGqADireB/5nJOv9k3BW1kizxGbqgKdALxevxCqY
xAtHkL23XKJDUmeBQgru9EqirfLBmZ6aDAYFnZ5hbsrwSzzexJvSCOC9jXHOErOw
j1O3FoV+wu79HRr+QIeU8OPX9bIKjxhd3j/Jw13UW9QBl4eH1rmHIG0GjKuRSx4Z
D2v9vjw9MZXhWa6HUNeO0B18vC801Zpvv8v89e7nfk+XyiWAnwl9bNAU103Q5DpJ
o0XCtuyjXDXA4zIWL7UsHYX/n0hEcDz7AWpAqThwaRWxdKBeh6uzEA9DyxQM7Hw4
GMKTSuFY/qXWoZAzb41DnpxFD+On8+dD7g5gwFUSqqlUiZzyO9v7PNOZ4AvuTt2N
9/6faPxOGOOYvGZHF51FWf0GRVsXhn+brE2wYNuRj1GvuDbYw5MmP9JpIPWWfcjt
L8/yBYS4AuNlwnWHcyobjXNlSQ9mkwrZj4vITTbGiopu1f4qgk8jvx+idJ+ef6xX
P5M7L561LQLGocAxM2oRTQF6r53WXWI9z8qiRn509hUqNebCDYnba+WhZkBKdVvN
tVVoYJWb7taccjYoSx7dBbU2ynml/UCaKq4zlHdkIWCFUwn1y6DBVfoU6zTZKxKC
kq/irXzbooBqw4L861usJDuo4Vp+yXA1YvIDUVIezZ52y86OB2yGEU75jA1/++2i
l40DbZtLu7zeL+FOF4dK0K+9HkWfWpX157eODdc8ldBbmc8jQQAgUaAX3cwDELjP
eUSxujz5tIHvkHMUyrO/0J0xQBerCCqIB2WIKAabT91GxdRM8hy5fwNmK0pDpqc/
HxmdDRK0iw1SAWwlsuUSGH2zMwfmLOeQIp2GY9EQ5b0bi/VAgo76wmrf0A/7QNhY
9PWY2e1pNag7Z2QiuxM3IamsnJRG28wjVxWHmxUsApPZK9yWpDStNDpO6FGt3301
TSmALObw+kSOV/tZwz1A1nkq/yujeVQspYSpiB6cWlwFfa5TcDgFGEtIpzcDCHP4
QAKKGWiK4ZIUQ0bM6bWdWCsBw5YXTAL8AZEB27n+VvNQ/qoGSmsBYBtcye4Xq9FL
r2L+ZT24gG41sjkeFcjvfMOoth0V8xpSx2low5GlK1JX48+Qwkslhf2WPO7Gc3Yd
mqoM62IKtrxbDL6Ch2mIDyLfcgKU/0t/vupJIxoMyDCAJcQ37/pjPbZeaom9nz/n
FgzkY8GTqu2Ya9Bdg25NGexG5NvgzgKjpPuKdJ4t5t7MkJHUZeunERVq+bhJ3fVY
4XihiC+GMbJ+3vWZbWfKg6fMwEQkOczMGlVosHfIYjO6wR4bg4A5fldgF2rIcnV+
tDiAsUSxrA1p/XnK7G7CEyWwn+44g/QPBcZsKZXtka10widJCec8098g+N6HhSPO
nRqEZs1b/HJxmlqHlxr3SOE8AE7uOmjD3ogGasZf+/0LJsr9A5jer6gFKtm86EP5
hDheNVminqE08FuKoWUPhMaTqGNiZdWGb/QBVwkEvuv8bWZGmx9vYBdRS98xXQkd
JCtfLeEmIfwOLVI04cJ9ulgIeTBYZSE7dxYZT4An5QNiKG4aR53rPEmgtZhubu+p
71Hspt1QPbbrNbYNXqszb7FoHWkrQXuhDASUS+qZHTdm5bUNeAzlYFQXjZ6XdAxF
ChHguKr9oxTCluznpZUHHa9Mhtq4HOvDbpHLmxeZ653UT8adNe6hpAByp3OApG1C
rfgH5CddNYEggvLDWbBzzM5DzmqqiQ0pzdpdEgQRfP2HQ4zNwdgg20PXvI5iGeNV
RrVk52w+tIBHTtW2/Zr5Rj88/AQn8qoblLmH+nP1J4fKaYcWMH2TFpkjlQYC884b
I9JBHyDgtMoH72Dos2dU8lotGummpXZWbhfF2fJ4i+LfAppCOKYY7jhvyD/IUB6h
MD0IfRP/9wazYMAD5z3/lrf3Z6dvRUqWplocboLMnfIEXdQFsvK98QQyu60822VM
PLL/Thcaw60qrr7gaKF8SO1em61cpkInq5fQ2iZZxDTraO8bIGfwJ5GZz5blSjk3
Pr5NBPWYmFP7HHR+ORthYv5tZTBN9crZHPINutNgeckE5Z7Om+lA7N57Bj/8/onq
VAiRILSoc1UYbw8p9W7/jwnt9FOCooTXqKRe39LdqvevMs5b5MztjXLZ78XDR6D8
jQf/QQ27W66QgDx4PdHMIg7ic+i25qEZA4uEUvDD2dLdeMUDbxTmcI5BDIZ0a2yS
m6ydYYatFflAvUPzm5dqCmmwCvWpieBbkj7JH9X2KXymBctgtszEzNXdaMegEiEj
h6CwKfJDBrPFgmCsb2yYN8F1TZci2Hp991MfiLTiRosH1Z/ttGFNx+Pn9gkYLT0N
IsO0z8DxhcEl8EmvqtBuqWHRJo7S7A6zPUvxSHgEd8GTYo8VYmpceYI86CMN77lL
GNEGnH3Av1i7gXG1n4uz7yQ71eENPGeO6E0ngmyptc+yJJM/aZOwQhStTWuAMCGh
k1E8TUab3UCmnS0pHv2lfQ2ElMxiY6o/wRH0YylQVZOM3kXUkeQBsOPBLoUwUe4M
vWt1WcXYsMbLRTPy4qqPzoFOXzRQLLajKzAKDHKla0ri7DQOx7z+IuHOlyAVsarT
401LxiNu4fAPQnM0fKjsB2CzconCVms8jumEmIKXGJUZd0si04nfZBslTKQeOTVa
bCNepqPctqi/tB7TBjKg0Ru3Q0yOinqe8Nqk26G6i1T8lIk1YLTSVzMadKGbJmmz
Zst8pSdMa+PotBaRjzepUAXhalmJy/R58xh6e6BA+NDtSzsF1OgkKnOUsD7UDdbX
QalRxh0Vxex4kn7ClPBMkRsk2WjfKZW4j2Xpc//H91IXorxJWqbFEtyRmg1XoDFj
B97qbQJHtobDwMh9EoQEm5EGJ8XAbpUqiXFFy1u0L+IuxmFrDKo+gVZN06aL7HTF
KVLLYDZBLaB/giqu6KmZ0ewNaPgAViQu4WL7DcXP9B+4udvI2103pvERLG6vaTQA
DUXHQivvjCD4tO7N1WanLQWu/HBpCskaQt/vK+/MY9wgHQIFltFGEm0jWXQwDsdx
RytutjdHBheU4AXh4y8lqBUAqZWQaZ9CtbLY3+o6JNa6pXZ3nXa9efz8V0G/28iG
leICAmvC8PxOdKwfrtJgOPV76bdnDU6aEFVXcHnNmneTLsEEgEtXWT8w1p14l0es
y9YebAgOo5bG8vc1VK3ktqgW8KURwJbFezAjpPXxde8zlC89oCgtexKq1bDduWWU
PL+jJQwgYAjj+uQEvK/O2Hn6DOniPjdpgZcCCdaLc+cbl1isZkITfh1KsQPwyGIN
2zxuxxX86m5wYinnRztvOZof2tuLlNgUk+lNdYikO8Zwt45m7YuvqRp7MNts/8Fb
UKUMBycIYxt/pwAyGHX6cSKaNnaEsiQMGhiMM3ArCXVnS9XDDClRw/mCo/CJqMQV
RQuxC35MgdxYFUJJCq/SD/sBDtOXFf1LpTsnzCYxv1xAFsQ6c6QyhPkhxZxQn2WC
ugdD7litnWZwhmIgukTHQ+EkzLz+Ze3cx/lU+Z20qzbIRm0Ypcp93yNjzv+qy35Y
mKN/9f/o3NFEzKKAiY8G0fcUnT5AjQS00WHFzOQRMZmGXelgzjpwo/NHxD6Wgboz
eAAZeEYHVkdOgMzyFfQfZ/frL1PMeQnjii6iUQIzsYNIhr8Gldh0ZvQXcgXaTxCz
w5WPoHOhgXb+8wMa9SU7QOpz+o3wcArZ713jA/rg0/sD6X9rJolPxQBrV0oVlOCo
jOCTKOYzcSntcH+vKZzmwwGVENTPZW3Lu9XnP78Qmfy2hdik3dDI/Cwa+JvJkNc2
/kUBRJvGRz6MoQI3QuRobxBHoigK8/4ai5/e//fMYdh1swjnwCY8aF3dFLX793oV
snOuzIk/y+Vet2xiz+/xNyYbnDA4GgxG0SUlDxwVMj1BNrU6JLFOf+/lS93iL1OS
9077wO6ARUqy7kXRhVN5+5BeXSoCn1jWmf8LvjtEQmx90hJWIJXsWzJS2h68HvxB
6LiX8G0zWaH0LwXu8Zw0HD6cdhJJy+g5fQ1kiqYAO2TUUY45f/qkxbXGa/ql80R7
5V7ig8++snYGc9HQa74ytxgwCbnZBh9wupHc6toLLsOO9skO+9PwaR2GSZH6VWIJ
9dpOQg/QuHjNJAFVVoz7WAmHrheFh9JMN4qMMFbwr+Ty4HsAYuscwEwxjKcDco6Z
9aJqzBteJrMGm3fOMvor7nZ39nr3P+JjQUHP7K0k9K8gz5ogT1rR8jT4LSfq8Zxt
LUYKXVV/x19F9vMmyOF7N2xMJNo2J8hPb+3ky++y+55YtAVzd2NpkPeEjoyUMwva
/hUKkswIwcZuk79WgLQ67VwZg0SNYa1BrOm9JX7Wh8ZgVkLu6BXnL4hO/q5PlkQ0
2wK1K86Da4hKxbR9RDrIBZ123vquqF/VPyJZmfHuwvoWfSAwtUGqMq/cXPfxoxx2
wf6Qc3tGx3hyegwglheR/D8Go8ZFae4f+AQghpt9I2KWh+Q6Omf4le6zjhg9VW86
fsGoPkiASaPZdufc+5tnDf0iGMOrFuoDjbT0C/KVFD25DBN2ZU7KUczu68pbmQKn
VJa9IZ1zShrCyTB9o1Rv79s03d2K1AE1VMg9vo84eqk+sRBTMsqmgXA6YAPmwE+r
CgBUJkXf2RBwURN+nuHC1R/P07eQK1E+DrsngoO5eRRlDKVh9NzNNkGTNliyq9ib
rUe9oFEeqX7pW/w2R1yJ3CNcGylIB56DeDBcX2fqCdfeXz3Mq/5xriV2CeOf1utf
EXqsGRpyea2T3F3ZJhFHp1GyZJxNj2CqcaNzQld/pmlRCpfKdxe4MPqtQZVdN2UE
WbK1Phao2bMxhRKlCFWVMgny1TLXZVWzwuvNMKvDKnXbcRkAqtC2aQDEFus934kv
LYB00xsEsYDcS80mbDgi1z2+gTCJz0+JRbuLthjIlYyqvu+SuYCa4fjuhv9z5BsC
3RhKm7QyFhRo7R0htat8hUKoV6qntxgyUPxLbUJtAHvQ+hw/6Ti1rG09/K7A7gT+
M+wsbjkFNY1km/hxaDLQEA+yrcTvMpucOd+6LNE9hVv/+ksU/Z2vTRbk6goPccGY
Q5D0FZI3hlgh6pftqVQwuh+L7IOEhr+dk5PCfKLkZ31YKVFDHTAO+lvVPti0cMWX
Wbzax6V3EsYBVJdcqiYlqqsd1F60v4goc0Js8EGcmLKO38cmNYGIO37ARcpUxqNg
2F4ivJ+dNfK64Lj9KUrDQk9DN8GKDY7x3loyWsAdUeP3YRFUVN9+CdXXYZVPSTFj
pjf0mM3LQ1zb4EoSPfCUBZCsOkneyNuQpM+TlhXwM0WTW3TfuEh2Xin6eIq431cg
CTRZYMgwCTpCgIbbn+s+ncgcoxzrc0ifCikmvGR89ICTsYkqcGLiN/sH/EFPouzf
Gi3rIS45VPAPMQ+aczRyW3XEr9imh0nCXItdZk0yHNF/isHQM22G8dzFcsMcLyUu
lT/N+cLOJIjvnHOGvKLWm1fzFgYk2kd7ui/vzsgXiV5sZjUw/1ujnKI9uaY/D7uC
C3ONNSzghMHYnykuo4pfTsZ98x5LkODDOclZMzXh/shCuz6O4KED35JDhloxEfFK
85NNfQzy0XMYqxRpD9QExbwB4dvny5cW2kVIjWu7UytECDifFMiYN1rgictdph/B
7eKMBUdFwnjVDmg8L2pwlOZyPuuZqBNV2pJkIzfh+n01kyBFyuFFWJDh3Keq0KiU
yV+dAEdQmRlpH7+r5I2dHAipzGrcInF8woyUljAZMTq8MGHaNiQM1kw4KgkUXs9+
xknziirC2/tv9PUSiyvqUe2kbgcE0XtkBMfjYvOjP5PgFf7tIVvw3QvJnTI56jB9
TCpZfruYCOz940vv7TJ/uMsioQ5lrV3B07VyYHUiIdRHhTmaR/L5Es1pBd1Xox2z
xbTyN0pMBNHPxbE/1A8ietuyymr2M5nFpb8hwZzzVLlZ0hsjSfNakHjkPD7onqyZ
UG5nLJ590hbZmLY8V3BXOPYbcIhFwKm8OLKKUrFyAAFyuJ0Uhlb6rfJQOXgrjtEt
v/idGdu3q1yF6OfgzpA1csVeOPzqjV541OvmZLB1ttdK90C8UkgOKJq3E7m71ujN
aPXgg+OW+pW6OBG8Hr00Zn20RZu9VyTEShsdP+uzOPAg18Oo0T9ziWE8VI2N/nwM
w/XVKyjqr9vrbzR3xVkDmSpxgTF442+f49/S0+wlZpEj8ZLrKmcj6uEec3UYJ7pE
iJtG+IgxzbHbp+dEbN3SH7C4FxEX/au6YsrzjSNQRzbF4GnQYBHE0WpnEpb6Ud3Z
ddKuulnkVVZi/v2vJeY6LHTFNErx+ASFvhsKqLiih0TlBmffk/Orb7Wp2khdQiic
pKQQ0iEQYN8ElC2YBFVo09b3x8dl8WxRKWPpSMHEi6boEwQDWop/TOBfxOCz/5uZ
fAo4G1K7G3W7xT6RJFwkvIzdaQHlYibxzbmVcbWkCwGcPQQO31bQjStLlj5Ax4EW
6W6ako5wh0mHyVFJB1BJ5IvuoQtGGiC9MwVjvns7ekrV0zUWoZ+/K2plLNrEIpKM
+dc8uVKQnvBulUmG6/ev8I9eUoqkk1CaqpiWPPuOTWaOQ9HEqHcLOLsOB4IOYQaV
EkX+E+XnYjVGbHB1MIBadhvb0/YBylp8s0QDX8iPc5w3bFeWF8Xi3BgCBwr444vn
JA9r61foubfuIO8I/ANDO8zsdygJuUO3BZk9ZvPFwTw/NYcaBTll6TUYPUt9N1Xo
GKAE4LX/90mqLbjL0H9r4WBTwj86AGYkjR3o5C0Npg6oN811/S+0G9eMCsveq2D3
UAGvZeIXBK16jMh/31GhknqwcomsPUK9i3wROGz8A5C3v25g9NKL3Cee3UbFzKe6
VBV11fWmxCjN6kdsPSxBueciHCVjUJ9tnmsE5ZQuO+sYoab8dWlEMiHIOQwPf2XB
BKfUWpDICo9zzL4A5RGMkoX8ChuaegSOvQuSvSJcFAcDS2q8Tz05fXdmZ8uL1QHA
VtMVqJpkdsHnzNwtx7HHik82kz3dJBsvmNkIi4JfJ7f58GqpG2l0zyyYGO62+o3+
X+PO3KN1ZVLwOwdkpUqoPIC8zUYWf5b5fPg/6ymhyW/6lGXzFMckwTYUKQTBLlIz
UUpED1rne7aK4Vongqa/DfyTMwLOZF8R5Iis/U9GZBOZ+cSwYzldW/C2np0zHnNF
NgtYJ2IJuBPOca+cGXZZHM8FX449eC0dJBPs4JSc6LsBteQsZScZvJ2FOn8LlDPw
AW3z2kzpPDBZgfuPCSXXX7PwHeJBNuyRTeIN50D+k3Xq/yTayM0oV0Cd1kpg6eN+
qLulluvgFmaAhvN90i14COc13NEvoo5zk8G5nFvQFqmsYnFyj7k9Uw3favJttvWw
ij8GKSpuOBZt8qNQdlS1YKYxdzS/qJRX8/XfiFiJu9/5Yyd3d8bqsaJ1QJCfVJm/
DxWhTu1pNSujoJxZLW4HWrI8666UYv6D/mMU1pOiVxd2edUKgCxCjXROTxUeSfC+
jKScOY2+Agmvvow6QMuXUJ/JS5T61KxOIqUJoPawOfkaxCFew5DUqUMQhZHYrIgf
CrE+iZathL6OW9zhelFNqJ/LNbTZt3r7BZvKWIpVHT28PVrrS5SSlbAkJd53JOoC
b0JzsQ0TWrhePVqKWuPXLyNNqNC+Rdqsnilk9P+ccWy6UPTKBMS3qHLAH5z2dGpq
7pundOrHgQjSh0XdxX9u/itSq1EsxcvK96lohi8nkhwCDokH9bS6r8ztY+ie4oJN
5IWASJgC8Mdx5MmaCDP2qWvHt6pKcECFzggVeDEA4ABxjljD2Iz90f+0CYnYt71c
b7DEb/J9Y4lgoP5vpgIdiPRsbaYcyPpTlQ6FEWtVrEE7P9JDH9U7iA2mWVV+ySR9
HgB8PdEjCOL17doIGCpHfy6Ry/3bOPAkPlrqI6l4IP5Uj/yIhPnLIX9R0nO8yqHy
GG90sppfgcdgQMGOiITPzbjYDn1mjNDEw53x3nNvphZKgXUw15ESdcrunXr2HtnX
/uNXPUVJCe4gbZ3b5dJGLwTN5Jdbw4eNQN59hqBjaU5BX1RIFPWx/oHBGRfQh+JD
Xuo77ux6Oi3PG+UtQ3DlmPQ9UDFPTP267bBax1XALbxajEO6+75/7JfBl7m7uoKr
xEGV4WIoBtUfIm73rDXfrJTfIUbUmp0AmWbu+RIUJDtHOlqhX7pOCxfStlgKzIkp
sKN0FL9L7GpCgSh0ehGb9OifOTyev03rAaAcKUsibSCXBvWizCoq+zRf1KKCM2Pl
3fXTQzl72t1bb2KhIA6uy7SQWLx/UKOshTFYEIjhuVA9ocmj892JewtZIRnhpS5e
N6RJXZS2nxjEHe+3Nw83tII5micQfIRUPvp8nqj3AL0ymVKGqw2uY7wRmJzMmFw/
PM3shwvfI2y/rfqQYGKkLNlHtxZnLYHb3uT0pim+tP6z0NgqPc1IkIa+Cl2HdolI
hecxSIzMOYB3UhdzNyh8EmF88kyPMUBu+JF+4p3tqPtFxYflcFynNNRIIp61/Yex
ZKiGfBWmxcgDSlGaEjg+F2PMgTkhFKEEswi5DG451YmgxptunPzqZngeVb/5U1UB
ie56051GiQ2bWM2xzo49rVsf+HDzgHw/zph0Mt+daJRVmF3naKPsLm7JvUOUURcD
jhNKTSCnllu8hQc23uJ5MhyX+tlMt13BJcriWMhX8vL3iCfdHl0xbR0HVRTWfRjt
T9It6y09imKlRKntaWLlUYhZkiDdraB4OALGHr4y9HfIOjeMQ8slEweGVUzklzRt
ArKwYHQlotPmZLsnkkF9A2gdaYepwZUvxS79lTehNr7q2XhkZ4Kxvgytx/Utc/+y
b8yFM34Mon7uM3ibaQBDrjoc4N06Dx6UeM2QyXwbT+lRbHSUyRWyj6tQI1n4JQor
aeo3VK4thuUyxVwHg0RdmcPAp7CXYGMPBTjekSMyvlt5WCrPrJzE3ArjTkE/bZ4t
2tx1ZF8dkXSIsXohYBQUBnK+wIYzclRqjh5aQyPxYubmjKhuT1B/1xRXLBEY2xyy
Og8gzg0BcLQej+4nRyUlC1zojnJ8+t/2waM4HNU60GVHaDh+UMKM7R32nVipXEZj
UMuHfrX9m/Nwi2AA9SNx9MiIqL9ptUYZAgDURnjhEfCzkfnIdoXycKKxJSNcy6YG
bI/qoATnLXkCWotrx4No2UiF2ehkH/TDn6o+AOfsBm3NJQuBkw/wHwiYCoW8GPl9
rK8Vfdo16Uj5aP8aaQrO3v7zN7c0Fmj6RvAWtEfzch1+H8QcrSlnsqAvuL3t0hQc
xwbXvnRY4xd57bcer0TGnHfHjhsyv2H+eLlihasnjHiRJ0hTGx9Gz4f+ivSLzfxg
Cf+dZoSvwaOibQB7rk5RC5A79yAtTzECKWjwHBUQEDwbcFd+bzU2Ra44KbfIMRyZ
ZjiSXeNKvND3+mNuuyo5ypq1C7FS8ojHJ94qo4OU+W4siYC3l2Uo1rpNarYy3r6z
KqZk/i94kLmbOJruqmuTLblEGUz/hwf8vsYLoA9fZLg+62mKbCyD2nEJt1BhyIE9
/vXECDRFnUEer1SF1IGKXmdhKbr/TWctuqLEEjFEZ0K1iH/QbkWbcH2OoqgFfo1n
3LTFW5+R8xaabJSLBNhdh1yO38gL9qjZbRZNls21+3Cr9rEYbewFXsjkUSioT7d6
rAAKQ3O220lNlGU57XK6S5mPncrXNHlUJiZCnWmUWqOt6U1qdw6tq2am3t9JsZJz
/wnWBzNVdiR74RUgR+JZqz2kJSY7Yq1Tc9m0Vl5oxqn0FFXbQTkSo3NI4rD8cEuV
KX8Fc4DJN4uml1Q8OuCVyggdi8nMiXoZBZQEjfClkBe/yRsxE87b1RQmGQ+iDeQ+
5Vj1ZQ32PBgWhgFGzlbGOnuV9ALr3RRKccxnj/MqGeDlb3HAeX4Ay3CKxK9gQjSe
Wbq8Q66WvwyITl3pSuGRjr2v1l4Szx0sYQnR1A7GwNmTT90yCKxHnXQgo4zqlYgt
XqmoKEwTvBnete193ErRqDz30j2rmF8ShAWjgk6HKynYIT48dJquUZv69Un05FVc
+aKUrCvSn+P7JFlPT2SH9E4VkPOgvLXz//6MwwmDTbkAIPZdJCWA5sIYTAM9Qxtr
XZWobozRbCnmF4LJcvh1wjwC6g71onTVVqDBeIYZ6DkHoulHPUZcDAMm2fcEbNWe
wWhV29yjLKVS6Sm036DwzcBdzOkLW3mF2OEd1gHGq/ZEbiP20yZ9xZFsyTRtTAmG
nmczL/brYSK1LWUkkDLrRlHwrXcFh6AVWIohXJhD4GbShK5cviw4bT8/Ylo6iHI6
IdmyvWCjCjcLHEOBW+i6trhS0Xs3Q45+5Vh9QyzCDXPa/ZJHenyA+25XXhfrNc6d
BCJNXyK4Cdfx8rizekdJXhels2HnuAmQ3sLF2qGQSq+EUuB8rOX4VRH6XhyV42Bv
b7suhGz3kgCK/VJM2H0DoHzDA/Qgmq7HP9LaQ6WB3tfH5liPD7xMSoSll8gi7opK
ndeiU093vj7XM/xZNezlBQqkXBsw2VAtor41oeGB7eRkg5TM36NSudQ3GsQOrBCH
amMKmX7r5GtcY41/M2Y/VkUhg1R4ejDMauik8QD2VYsnyilZ3nKJiBWfihRVF1Ql
UTTyFoc2V31CSKOrWI8nW4RKX0KaU/qt0u465lip5gIR9YUSEqt3mppx3pEwm/O+
0xS9i4uIovLhJpv899DkZzw2bdwx4DQFcNbl1epImOU0l675oTh+mU/dEFqDRq0p
wa6CKfzNJ7sMHs651wMur5SzqEpsR6h9svMnGuLwdRV/M4sY1Ps8k4lLnbUH2OhX
I7wIZ6HRlIWbhsRMY9EwAsJ10uEUzisaNf7QsSgHpz8Zh9pzvZ7recPu3jUm+w5J
EFnStRYltUF6KeACM9FiTAAN9C1InFmvuejnwjC2Wnvmura0rluFIGEmV4KlU1hh
jA55ef5SP7ktyOHRCOwFcMEhxlL6rcdPB7+nUJ70WVgsIuyW4Slc4u73d7G7O4fL
g8do6QNtpZnkz5h5jc9cOIo7Cl1KRHcsDYvRasSdelSBViiAKtH5vNbnsGu66sx7
sDtxTQPQFidQyo+0GlvNpvJUdchWdrKy8aUvG4+6Am+tWOz/hURVpVI79CrsvTmH
ZRcZA+/b3B0QISj1Pg1ZMhP6zcAuYU1NR6r6A3F6/wOb1LP5x1cAWAt+uxSuIDRe
BOPjcXUjzVHauIaRkSAmMwf9Q0wNSJk9gT91AIANbKNNjco+ezODx9z+JyFiGKE9
RDP02QkGNg983G05pUq4YwSmFnvgGjHAXNuTpTGGVq5CLaMxF5gIxzJg2m5hViCe
1QHA1MsCiiGEjLsp3yIBw5e5fa/Ze4TNDU6wzO89SIcR3uPXhJuqaGsJlrzFrkk/
DYnlyq0kbSgVqXtk5HdG0/ZSyb8lU3ls/npHG1RAWVyGVxVgYsw1kCpySKs52MlV
3TJgG5oePDa9s+dE2AnZUXC6bn1Wjt/GCkIhrer1oWVRBizFlKJU5rY6h0l/g+7E
rrGR8+JMqSWNkrirX5aJTWiAfAiTlbhYjzViTmBixMb65GQym17BJtmS8cf892Sc
tiP21DMO190X9e3HZxJXNId9sceDfol2smRu2Uh4f0tVBZ7ZLZGHdKSVuI20cISh
3OFey0ayCwXhM0Lq72QdoKog9axrpguqbcEHWovnJ2JQWR1s6ZZxMyAiMHEAI9fQ
iS9FYyjRsPNdr+f9bsPOpDarjp4Awqu1W8pS5rEP93iqJfh6K2lS28Ud61238OUS
o746W6493QIiu9JuLx8MR2E3sTz489zR45BCq+T+PrCfPOTxprZG/Rj/D34UaMaX
4BMDDkz8TEQNDr/46juH5BwsQG/l41Ik7LndCM9iL7wnUASMe5XypK+n9EhkumDn
ZmQJaQK3h6clPT2j9UxkBLUopNWuSE+Uk6RXSk98nXEckjOVhfAQVcgTnZ2gwdgQ
wqrmhgi+osaXsd1hyPtnAXpNpd2xaDNM0c4NPAEi5ni8PUZbcdViAdSKRGb2xTfZ
WSw3bmnFYjEnSW7ol4wcNDqwUdfZ7m9noVniFS8yLhStylp8Wt5EbyrGAihyx+ub
Hj7z4GWUcnvfEA2FiFNy0+j4sbRbzMWS6MoPnirtcMtEPUrR+oAKmiBehB35DGyh
7u7kJi1IpnV+Au0AvFiX6j0cACit/JiQq9yMfxTUl5ksUtfAvJViy/+YYIoHpvjC
84KXH863uiWIl0R/CcCIumvDyOn7RFqjatu57sPyyYrSeSonspR+DHk1n3Pf4yR+
anp0VNbOJb+YCN1k3vEgHI5gikgNR9ShkaH2l4Z0PjrtqLrHWkUDbA6kPuApz+UW
AzQcPwXGu4N+DJStMpErD1XiUieRI86N/k2tg/fNZ4MNfX7+B7iOsW1C0kKmxJj7
PIZBZyh1c4N4ldo6b8/WWAx/DFTTfNDj18oRiNS+xrwb6g4sbVtx8f95Y4XDdBoA
L9Cn4x5ETCGvhU3v39IvB/igCFB1huVwPMzARi9Jq5O+NCWxkb52n5CXWJd3rsrb
7mWFfskgajtD2cB7tnPuTrXGSBUWN97u1wsyNI6QOVLr+ya4SLHLYPrmzblJhNJu
mv4WuhC3USl0CfnTSd9PO4dR3jBddC7Tc/xVLs3r090M8XobHmCIWCifcGdLaId/
2pedEDR8eqx8HAcgViSV3bwp8xnRua1PYhSw1p+wVrx3w2bQXwfuQUrLHjT63rkc
6oya2qtiDJM7PdVo1zAGmbieU8M5pbvWVZpG7h8IsPrWpnokK52W+UD8HbSrHRWg
6/0Myonf+XcSNJjx2QvJwTsPtlU7idyJp7MBifhdhWRTGLYzxAyfkZiDLc8FKN2T
whJ244JZ0OdqifASb2lYR4yM26fzzdeTYJ7g0X51fJzMWggtC4HX3csTZ7Lajsms
TY2c8re9YBTj5IrZPG+ibP1h8d2nMfRA4X/Plsc9dMqSxBxu1dwZeS9vIeIhn0mC
deF0tZ5/DCQLKg5xiK+aXBBwljonAKP4I+XRv9Dt3J+8ofbZAM8WAN+KimaDqMO4
s/tvBIZGpMnu5G/ofM3kxrP2/PyWhFeYlkvvnXt/QrZ6Qm+HaEKJ/3AQFvm+FuCD
FZkp7KRJXGYfhZ6pQkQukDWEliTT1uY2nZs741OCvQ+DZCl6WZbr6VqjFwLBA3aT
TdprDb4Wa+1a+dkAbMRNwrT4M9B2Z5gt4EC/sFR6LQRtroh+07gUOn/GDAG98ZFE
ChBqKrxJ195jJ2JVVWHc4HCMYfukO7KhPC79B8GCYUSs+r/4O8/j2EIvVYYHxBDO
Oce1WPdaJP752pIid0boNTIiEBD9bZk9uNoeuKwc84kkrB9eq3kyqWKrGK0uTtBA
x1sih3oGeG8JCgI3XBSQb9DHP5jD7nYcCssDtcdGAdqCX7gtcHS6IYLFkj/ael4y
ZVLuCFdcmrE5WTXzt26/rVpyiWJSaRE2oUq1hzJtTdsoGuhSJTjF2M77Nynuae+D
bN57dUAnmaWF+ntiXQXUXLPVwcDLr1Cc368ZSyQ7DxBG7jV8+H9+5hyzruzChq2+
/c44b1RiIbYJ7Nj23Ej8/eCRQprWOFDoubkSwAKm+NUeFEbyE7G77JMcBQRihtPO
fGpjvHgXZytG+76ASe4BaPlvo1MMIn6g/dE6YGmCErWaqCsNxCVZ1M+H1r9tIhJF
HdRxbkExv/Q2YaNe4FaobQzlsD5Vdz2K2Msr2kwaI1Kq8deErW9pGo93nLrlw/O3
mwQODWl8UHtyCmR0t0oX+1N+EVVCyZTlPqBcU8A6RHvxSSn/Wjzmx+D9zdn9leTs
sE9aIMIC8BaX0SseJaEg0a+g5Mz+ooAXfch73MBePJ6XvoCNrUWZb5GyHABE8b69
LHfx1yrosCEIM8h6+ZIM8LKCjL7iMFvPsj3zwZaP+naLBmpZWvxvjoRVM4Oi5okU
MrEnQKfkIBbETRM7Y6VsVqZKCoUg4iXqQxtDEVmwYmJgJyr9nUlLM19Di28Wzstd
DO0Ufe5gWK5+Lo4kGG5R6EtKEXfL52lx6y4H349DCfl1cYaOrDyxZ/nW97AkjIXF
/rkMNd1RCzIyI8kLcA4XmSAGmepUVlqSDJEJAo/oO7N+AnjnsW05gjKpRk3RWKzB
Fp2rRM3d9CgBNP7ImZCcAi+Jd5peh3UUo7ILUtSsQgUcZ7wlnrbX0OdZmriTAECf
17YCJD0tPCRXaGVpLqhDIJ9gjxf8/tCfia2FuWK+oxPx3tubMc8kUBJy9jgYmvZg
69HFxSDRFDrqKuLY0EKNKERGL4NxfQq1FGE+JnznCwSOGA3w2fb2BmT4du3Qxpa/
oCmmRet89/dSSX8u7ea0y0OmDNQ4qL140NBJItLHzHhwkTv74rJLzGN0XsRnXIB/
ZWbkh/cCTNjx0PcQFUF441x/hFCFd5ybbPd1r/GrxaAQmEv/S7gEbYtlpLkVQg4/
ch20QEn1YVwdjTn8+xBg4bgnaExZbjR5uWpdYIXXcMxWyHfdmX2LP/f7Q7nwibUr
yBhecUzXsrPq5MrDNa2nNuYrjkvEnnM1AghkQT04ymcgSCYhe1mmnduDxuKrMMAu
nm6vifBsDqAey2kyKx5pq8ryZ5bq5ohDEC4QouINB0YyHycJQ5NJKwgBAPmR5Gf/
RJNRJW+5CQpT1EwN8X+xChlioJtAakOQ0D12F9I/4fSoDWylZalMNElASkxfiHM5
Gm27VRx+YEPIQcoJxPD2ymEJr88o1QqHgomYDNYI4V6TSNAGJT6L0dSj/qj4BPVN
M58tQ4aKIJ596JGX+eNRae/EJNAfkfO/wewIkuQRpyfruKZxnGRkF3AxqYG9MdMq
4K0VZxTDHSPcUb6J0uJSAeMVsfgr2gwbhY0JWDpRd6wxPPIskfs7EnJWz0YmOEmu
V/Q0VdQRCuAJ2x8XjGAALAdCz1Y59t+ngTFmJ1KFPwRAqyvOFTy0lY2nET0JSW09
bPWAtbHh7rvz6DS2KPTu0ODG9RwqKhuZVf41+j/2SBE1Kkhzsxt1XhyT7mPn4lWe
yEVQ2dp6FvkhtfUPfarfiYdFTTZ3eh/luATt9raE9CCs7QC2EXQNkV3eYv/c1MeI
Bc1tN7533/deDFSLa0Vjy+9+epsL+fRJ8IC2j0sFuIohoG3FGjwgX/tZTHPyavF9
QUlf/SDFOcg1jeYa873qhx02/HfkEmtavaMdjO8/5zlfaaaD0PtmZM5iptwjMVHt
1pGpB3Jsm/L7j2UAei43KcdM2s2SGd911rSIx7sy6M9FuupIsVDdFatLFy1tRGyT
WvxqkXGkqySXL3NrsWZkS1gS24C9K9dCz/AmNrhGaD/HxXZ94od8VpJDgxsy6mge
a3CK3T2JULlwGJqSgKlh1hO9cKPe+slteNqrl0C0L+ZzsolHMqUy7xA1SGS/loZU
InmyGor04O7th7DQPGz+BpczW7C9C+Ncus7P8BNPy9EeawwbYHIkuird/SxqrFqU
cNTi1+UwdVHoYFE6yyuUQ6EQqyzYPlmIgHl0a9EaJDaYiCI/pPZCz9WsWfwfn4Dd
xMLPydBIG+ZEx4y0HbaIEIVA/x06mssUxXubHSAlFUAy6CdVnL0z4gImRjNfFAjv
Ct4Ih1bJ/YIDiHxij8FOIty6CQhlDSGNj6CxCW5wxJaLJDJbnYCH9Sh6RIiP6a8S
zWxdYB5xLTd6pSEC0YKZT7e5G33Qf4LRdlRB6dYGGC6dnq58u+XFqQ3D1IQvhVu5
qAIfat8mi11IvwlxVfbZSfIObkb79HnICCH1edOAylob4EaLly7sTt30letWokOB
rG8bcU76+F35BVX8YTh2autDiAbpSIJ+vD/yDy6uOHnkotIbfcYPMrLbWgpUL0R1
1btr3bgoXgSuiVh6L+Ae3J/y2nOOkjXQW/iVGSDGOQERFDaYSSEiNDcwC1RWdXKW
n6V9BsCPP4MJNw6gLHmvpV3Ix2J8qz5CQYK2UIfcktzyHIMOE7ADT9KgEPordojO
C81F+nL8iRZKXkWW1A1uMihJ8mEdJ2UOnZwGfO24kuECbLdL2fH2A6JGp0a9wMd/
LrPysZtEvWsXS1hADVz4E9EPp28eNJDtPPtYCglkiUbTcI9iN8GR4zuAvBEK/tMt
oWe+/hSTuG3egK0xM06h9rFDTPdF1zQh3Q1J7O7+Op0ZvapSE/fwkHEOhFlFVY/9
hSU+8lyB7o+Fl4pfHUkHkHM8p/YzkuYQ9u0nfhwv3i5y/lco+3roQUycl0m/OBE4
+oMgcDKvOmqotoDfA+WQ0BGK04+IFFhSvXx2+PSJYbuhtNsydU2KqHgieJrgnmLF
akRl+IbiPphQzNhw3qTmDQgsg/Vi8es1uX9e1pRVWHL+8lgcCOqFcXAvDJbBMTzm
8Y1rJbCBCdnHn/9uUEtZ6Hq65Q8LI+MSjktmaeuBnebTkxZ7DIHIe2ypRcMgQWcA
h0ckDlgA+FUhsQ7yOv9KRC4abReekFOm4NQMV8YZPJYmRVWOujCFEbguv1RHWd5a
629Ixj2dl3VyW3/gk6niIeOU9xvezmX8OFgxgIg8IArqPTUpQ2o64JoRCQ84K1oa
OymA009ajz3eeEv7ulyZTwMpbdtCu0Elp9Y7wnP9mXAn2HUIvC/ipZkVf5ndNGJS
r+wi/vf0nbchUlj8sgfutvzKuvyKaePtnvucRthxdPxgUynCJM1ehKdwexgf0bgS
aSCpAnbMAT8LLWqbThFPoePzbwlhDqAcyEKIR3SiWd1qu6scGyQk/QHAisCpez71
RkfXGL9RqeSS38S+WDppKCr257Ml7p2VZgx+FNqEOyr5E9HA67dHv9MLfha+Isyj
MBDciyIJ549QfCdkCulCLHKArLaejMiPYYS/6+FUGxMA/SJb6HTyoz8//8VKe+kt
MHvBs7I8n0vWGRZfG4M2jNhNZpZA/JQF51mIOMzYQV6yvk+Wgt4SEAV7xsPkiC2W
UHJNBDYzYQmwMRYe8Zkx53voVADcBVYjTP1wlh3G4ecIrZ2hn+FGat+S9ZdtmGUc
E1wjyhQIeuPGuqJZmLMrdkpjqncVwAXEadXVmh8CXN5Bza3HMsBiFTcbida7Hw14
HYDAAlJ6Kz3gnYA0oGKI6qi6MCeoshKf+pTrcf0LEBPcnYRNtPUxfKXGVPVT5k8y
ZshRnyE0qF6XBcf0lirzBp2QtECd/Q/BcoSKLHaIEVMlSbbFxXc4SWA9N53XjKkc
lWoOma8X/JaKK8IDmbpFs5dAc/DYqRbBMPW1wMBswOHzQS1kin0KHNBaCvavEYzo
WMG1UtefeY1OOxhnqvE0XfMiaYgaGOaWLNdmhepPvsLQuEUIjvsrf51b/E3h2K0M
7rIPD05flfdzWrRQdPpbpXGgHEYYzYbuhV1VsQg12uOvyuxRWmJwdhoLtgxiMffz
AWeXXP0iVE+uAK2gLoBq39iS0JdGkDzC/Gf2IUH4sHHZyT0t/R4WEx5z4nebtae9
mcKvUHvgaWrPf/D9SeCisWf+yLsg1nk4aLdP7RJA6CVB3ycHLUjDFuw8JLupLgY6
0YoJkrSBGjkqH7BYtvVn5LV0WwqO6/bDoAT6wtzF6AWSz2BQ5m9dtQ+luvHmkntd
BBRQRR8R80nBrOfwt5eF/Cv/uh7nM3Ry0pCoh2K5O8lbH96Nal9LWSKqmAecFiv1
WUZxOIkHkpNrnAWh6AWyXO+akjNjYhzEpbBNTlLfhmI684aRv6CLzXUWshF65thK
sdQN3F8VIsq8KQRTRsifxBCC9gzp99yKCSQHyY7Mbi30tmu9z+0BVy4X1kgH8Z7D
bINFhh9JozIxI78j74EcpyzC+Hr+Kx8BLocsHY3DExVcVH/F7YQTgm/l1ba2tbNk
saxTsV336vCAwt2x42v25fAwQCGfCRVUsVx/u11BJ6j0BpdWoX29GESOePCOiS2O
GChCwlWXc4XWt9HoZJsVdG041Ty0VT9vbZ8NAhjEjLXHsPm5HPtjdD7mxSAMXTmW
v8bU+xQzmxNviYiwFj0extK114g7hMd2KqyOx8dM7ztGIxVisBw7cvhtUkhOP971
oVFv25aWp00sL8/tJGHzrJOeX9vSHZO+B7LU7yxHVaM3/560WHBMNPnKgYkTfnXr
npCrlMxkhQG/XO8WCRWj9BPR1hhH1QUNrV9zRrovvogwu6S0LHn+yLgC8/okfb14
H3MRonZPdkCyWWnNneVGzK0REHlLQFpGJB+VOS9VeEMBqPm1M2DnAAWoaSLbAeXq
fwM/HfR/LFNXt8Gln2FxAqeQVyEnuQP0cLzkKsZ+n1+8CgwtiH5cxObEDucSldCP
3p5slAliGQC2HFOahu6yFeseWAQlKeN7LMid6f4FnQ/osqYuAL46jz8x9iNzeA7d
RJsvye4rJMGsvWidDwMtDS4yfNUkEpeAEgx7SIJf/3udBeSr/z3fhy5aWBAgHhQD
qp+3dl6x90f/6+Gx/4bdq2S2EEMFe55Jg+BRMwObS54K08kSojJB4LzA1eanbYpD
vbCavMU7FnrV64frrvcy4Wm9IcKEP+NE3hSaqa45fIiW1y3JGECEYRhpZC1iAUB2
6uIOsflzB+kIRSuANf+b1SINiknIT0nuXyp5AkBnGBlDk5LiRsaf3X4wz2N2JsKT
8Zn5oXFkfPRHbLElI7Pzv+a4Hh4o958bB2OPBwJAIHGSziMY7KPmWY/bfAmB8kPH
+X1EackEwxNKr/7oWNzjfqX6ciivnXVnLMOwoCPSpcJZqOznfDjUOlQu9n/Dsc47
517XJApbQ91uF7U26iRur4zpjU/wHBBZkmAhqkKJHhTuubmzbY9oOSZJLVN7c9HI
6Tcwe+E+ZTrXDMHzK7tdBhuOFV9Zg7833ZyY+u8nkhD5mAp5poT4euwQxneFjE/W
gPDOEYNZhgg5/vdeRhABiWez+vJPYhw1Di+BJQIQZyZxSsRKsEPRRPcvjvV1hOsG
OyWw8x6df+bIS0fQhmUyTbMydKSBNKEgFfuSM9i9JcqUWE49JCT07CMxKWF/dNlf
MxY/OACM7bUxsa3BpgUoQWqQdzR8yA9m4xaj8BsetZvmig/5KmLTE3UkzqGGxU1R
m72abXw/FJziNGyKYtvsk3UrW6aAXoXPr+NuVlCI8UCM6XlP6Foqou7BiJIWfh9h
wfD6Hcx1TEqqUsdnVC4+uug2KqUyD2Bl/EhWqBPjDHSvlJjgLzJMv7+KGKblzMlJ
VdQEq6Y73B71yNAnYZzsF0WwNzTJAU1U6hEwzJLqViYMK8VDKMfd3XOjvfRZYKHJ
7Bq5imOn7O1GM6aftMiU4EpJpD/MCIHgv/ZkZxXlCqifjqrNLLX3bQimJaGPy6kC
s+P4yOz1T1fXlOrah6ZeL6PvuvJnUP1II5RQgZE4TH5Ss7Otktnxykt6zX0wh3tO
Yzv4xpPc2EF7ZS/joZRvACUm+gEEhruTXzfI7kqalTIJ5RIAPdixs2pDA99xMYEo
2UfPe8LCNaU0uT7HgWUZFBsCzksiDVYFuyrhzOpBe9owRc8dVTl8Oe5zP217WU+L
uNnXqUew4njDFfv00ftkolqysRT4dX8GlndFp2wA3UL36Ac9eqY8tO9tQSCXXcCu
0+TX49eVXjEwnqS9f4CCUKRIyJhCflercvfoK2dl6jtRpIh7w9JkWcHOCTHw+udi
aMS9sxsZyem+yNPa0u33hpbB98/kQNHjddI6LxLtzQzj3Ku35I613gVuNUUU7k8U
HbGVjh5Dg4GR1uMBmY2PGhLKd5ze2UU1iQr9zo5RIGDXyO73xS3uWVUeZIZFV7MT
UcrVjKjKauSKZRLQGCp091uhRwIXoVvvyO6FnvWlXu7vo0aD1z3eu4uDKOcchKBe
IX9l7WzgHcPcwbI72rhWfuoGLMICwSwd95xBeGatQZ/q9T5hUE4/6/CiqILzxDVX
i4teugz85QwUXfuKAPBo0BQtcgyr0GEn2mnJ3w8bFS6IHgl4t/6cFAF5y5vhh4Fu
ivsIYLU2rCEBL/8YhdswzjvbWBnkoI4/1WsfUwL0RB4/GNLsdOeJgljjmuAQICon
w4TJzq+H6yhad1TSbk+Wx533oU6avvD2YPSbVTWxwCVVlzirCFRHsXNVnHVmo5ln
1ZbgJr/yN0TRrI/PCi/TeL5Kv/VUucOOUFxSTKIJnhJkOTQhcAz0ItuUS9iP/bJ7
ClU0RjTlikg2VBeZfyKfYdWz8cmnCm9TePIknt6G04y0rdnhc7omM58AqNkClrum
UePHV2n18TQz4pg/ShijJ8OLM4H2wW62FRDlDRX+OoR6LGZBPUMDx2i1edl2QJTu
ANe0W57euELj/hkGMdmrTfY9M2aT+eNyuYKzb6lxANrW/9iTm4MskCUT69zzxzIf
s2ciwNqeL/ITOMj5AncciFk6D/vPbT23ix6qVL2VKqdiLd5HhvHKVEQQlh1+tnG9
P2o55deEwGKZgginkMOJNhQFF1mZKzYegslfCmwT9B6OIx19ALSIuKYxV05xCMDf
bhFtnrAXARAJV72arvF5p3dGuhO4/9m0lR6SeIgmBVJzZM0O9oBUeAfauZQfdiqL
Qm/VGsU8OVgN8POlrQuQfNVC0+v7eZhZf1P5d8dH53oy0iTzCcs8fQzq7LYVSD9N
dKuM3Xo9/gZXBnCRiOUlNq2ZXSxY2bRX0HkbpHbiJiEri2FjV0rN+nEesnROSMwf
j8Ntnpyfvxk7xreFksePlfvpbyBEslBSmnREbp49obuueWFpX0IwcW0loGVsWFAH
sb0G2a7G4nTNEHU5mLGdz+3X17FL/kBl0qj8wD91sdl6ArG5oSN3Nb8EId8xEedO
vEgSvWSdiNfQDLWihhvsMBcuA3B2lo7gv+d9AYkf9QQr6VSoHVokQNjkG/wVVyc9
Tt9tGkwuTJCk46D3l5M2EpcUTRa/CdJs+NI4nUReUgxQM4v+x7XWWJ7bHZrwL712
MfCI+Py9/XKseUZn4pV4U0ZAYwWCDZJnJbvdcTMOXrzDxVA2o83AEnVf6ds1mbhi
nObmyGQGcQlDRAzUoKuj6u2SVy6mBO1o+Tztm983OkGozBeCCNIZq1xfE+2buPuv
RnIM6fAm6f3/ua8OpuXjKXS312158gH8Ktrqnb2C6+dUafN0S5tD2W7ffI7EnIVn
de0i6cYEDl5mOCEar2AuqgnO/npKTuw5rvWViBzH9MQ06RcKsRSuyjLAi2wjXZub
twklYxufUk86+bi005oWg7OkBa8y59+WyUKBLG9U2tcyf//WqdcYjLQKTDdRsJ22
sYHTt1hqUUmT9j158A8ciOicgGqoXPju8lNuOLq/ngx+Ml/qVWVZU4AW+jjBdJeQ
Op6KzPcC/KSEpi4pUziLdHRaOMQAsBXAKn9Gp+NwMDC7vkocYsH3dapHWrI77jpQ
yoAeKnI0qtGsptnFgRSF3qGezYErDCbUuxrnfc2bP3meto1EHLFJeEOxZ4wJ3S45
eQRnTqjepuYZ+lGz9h7wm3X6NMQZvXDpO/yUUntK0VcWSZ5vingieH4cfrD9HaD/
XOJjVc9Sg0MkF32rYbUKqX3Pg5SOQojjJPShW9zTCMdoS3dHQQIgx1eNwYMsu39V
T2o9v9+mT8QjrVh5ZXB6/rkUDxKq7ipxf7AWQHKx1kKLxWZWP7RcPvUXSqgVsEdL
ProF7PTYiVtP+PZE0hadlwppzwwvHO2nvjI5lEIVWU92geLHtIjitDr/X/EPMGuu
LtAWkakSQEQdivz4dCgiAl/pe3L1acIA+OTXHG//fI6aKT/EYSB3ssABBmA+3RBa
nChLM244KyB3XokyAWGVl5CtADmMzQ741XqJdBJJAfpZOzJHGp9XSZqdWQq4wiet
WHjfsykWy9Mot2A120jN9F2Tw0+dQJ+lmkLUC0mPGAr0DeT1Q/LJwSIpn7Orji53
7DGgErq4isSfNYSnGG/yMRyN9RVKCy+y/wvJHkF1wrvzWqrrNSzDBZM7u7h4yfBD
CAjAKtEZ+CXhJk4VL8UUP3rGWvFt/tj1sws7T1/loWwTExC94Lp/1s8ldtUfUsUh
Gj3eXFboZFp1N3kzGp/Cp0ns3yMcZ/VltjCIjgv6/qUk05JM8nPnoto02Qa2hddO
SRCQIBnCkxkUbOWyavgah8QvNAwTBwL1TEc94zu3Tu4jPVjM1w0cCrR+0d4L5/oM
qcrYpV6RDUCOBIrWgLioCmg/6BaDogmJJYHqDZ51FTyuwnD/O62QJQ/mqWRpntxC
7gePE3/qxCLMPMHyQRYcSHtw1fXhzC50ipWb+sglJqjM07E84o2KSRB4Xsqa5xqx
9HfK2TlnqxZa2lBG6jmshh+yXHkpHoDOpmRCRk4L/jsdBtjLrg7189W2CytzqjJJ
0ODDO/nWrbwbyUV0xJMPnXfwVHgQHrRHAdkczYf1PlCuwgHzQU98rgXJU8jnQRH8
tBhzi0ax3VVsgbmexHRRIm72vASN9RsNFyoJmkwD0fOISYaqAaD6c3zfQOdTEuQw
FmKyyzlgPNGReWPFdyLkyqqW+ekFgrfn9SZufQWfKlVtugRYDLkh55+9jt/VKqMf
a23uGmOVirWgu1YFRd7RRmY9t1Bfkz8G1JJeoGv+yheehwRxQtIn9k/E/Hut0TED
mnpGc3H+wVi0ovu4BMKQO9texJAFssSfWRtWzn0jqyOksLbEd2L+IsleRmd753rj
H1DHzS4l4YhOZIwJivUOQNifSDsZqJvTubrP+16DX9vnlROb/uj/2dg7nMqG0MYJ
McV712U/W3QDamNmHlc5dvjnZEzJqYGeukdgdV4z0Y4Jw2hatnAUWifJIc3QxRQX
F7bOZTzPZWvR8M+0/Thv0qe4+wG4py6AoakiZEMC0KHDGhv0kHfbaR6K/bL3Bumh
zcW6TZRnFv+QKNE6z/8duVJT4o+MEfpb48VJ/49eURRZV5QdEiR8Tg/WpF+zGUXu
4t+9FThhrQKaxy4M9B950DlmFgFYs6e7uRFyms2vQRnWXGMBox0RfeT8L0heMkUO
Wff6A/pcIh1gyOhLIGpfX5v35MirtspxbdU08/fHvMFuAd0Qek29dlDYh+oUsn8X
Udj25KL1FRlIRRZei8QqZ40qdWyoRG5+6uqN9kvjtsinckhfSEteZbbGxjXzZ6yB
M26+THusOT/Px0nlxDVgNagxENatZCVkzGIw9rhXi3Y+PLtDunZ1qb4fsY+E11tW
bm1k6TPosvI7JR1vOOLfxXN+niId+F6E2WSAxOFW63RFWSYKMA0wTmTyAQf5Sm6l
REkegdmhGT3hOMpwGY1INbeE3RZFhTQLkDbRSvKgQIwGVKV9FguwybwktXNz62iI
2EUFk2BVaKu9p403+Fe79mJ0t6WwlwwheoGeV0jK1/tO1o20Ul/0r8SnhJ1hUj8C
2k1WjxkjRXbz2bJNIRYU55zpfd40aIDH+trTNmQno8C+jGubrJf7Re9vde3lGK3T
K2VQL9CL1NOkYpjt3d6cZdKE4PNT6uO1Spz9ZlRIYJGa2XaawzECoHYoEWWNEqFJ
yYVdVreqiCbgIWmxjWoJoJ6MZyvm+NiieyZaHmOMogQY3wLbRhYMGRde4VS5Hcjv
JLFJmy6ovvUH+Ru+8K4q381GU6nzFYikVFsaIKxgQ77Ng3HZ3bxaNqh8Sgnd8k01
xDwGS+lw24+vS6DGmzcbicbdJRimth61AW1kzv1VIzI4r0vd6/25cHZddMgXqyYT
tZ8fwhT21o9GGioJ8ojttW0ilZw28gQwxIGiLwZmVBL7Eju/lYXa1xH2wK4JBVg0
Hsi/adiwqKwl71zRa2hTEncZk5UxaceuPvKeclYr7cu6PAj53udbF2UCHCEJ615a
yKkKvbm81k9TFBWvGR6JMmqstLmGfKy+sqx/IiLJhI9x0f9KDw/RBYbQ+8T7LfLn
JMW46YL7c/DnVlAC8D8eDJ/qjQwmPSbWbyyU/giL5dMGN4aYveeA1cMNr/XXq1NR
LjdkQz41Zfcl0kWRI6naWL/j653nxOqsG05zLd78gUK6VTQeRwHoE1RQpBKViyNT
YeKtLM8k/bsveAgHucIdJcq6oXIaDdbB18nK1NT0Tynr5l7aJS3QVAXH8oT2U0Eu
ZSy6FuZDjtzorUM0rgNPN1jqrE+UgJSaCN4jETjmKMxfBAZKx4LKtvi0QXMmZKUu
w/giDGgSGw6zRzEKrHC7W4gBhd10P9qAE0hABX68vti7f0dpLfwX/AbBCbOBqnQB
qGLv6+LLhlg9wiw3EXEjcUNMFVB15MSn38Lm+xPNd0+b5odial/eROX1lj6i481N
MTf/9BebZDU6CHd5uckBy+CkKQipVW1zMzEXfh2go9YIaLfuoDq9oW1hfEXmpRrW
lKZ+TU7js2JTi1CLmeJLJrpJ51M9NCVvEYaT+5aTXbtAEeXccvykGn7O5BHQI5No
st88jeZXSUX/uEdr3kerZCVGeunaiTbjTBD1qcKDK90wmcC3Dk8Gwya3AK4B4DtA
zxOePDQQWuxrNK5ZCyKJdFN7PY2bIzOCfwRIC/0KfW7uZdiif4Z4X27Dl8w8VNUN
WA29nXULs6z0dYYbdSrevAI8OyyoeKw5n2f83ENNSStlA54njnrrync3Hqd0kwvY
/Ft9jiE545tsWXNziLDpsPv8CuKS99HQNP4fHlLHH9eU7I7JxJEh7SJRMPJvDR4G
nfVPkbZm+AJxHHwuEVi2e+ns+H7PQYOHPbCXQWIe+oiPuv3LGGyxkF+EsDPLnq0f
QqiAPeHJATYb57GlLf6MHhQyq595P7yDFqBfg4jg3jY/Fdc/1abXVcUQUHpH+hLS
gQFN63Rcse/mZMpPDAM9cdzg00Xn/x1dR7OuMLssjdFpIIIxkVlgSTs1jO26td/4
3W6bA5nHti3PCMMZ4X/+P1YU+cr+dGW09TFotE+DVV/iO8s1SeIBBlnp+xWHmJz9
4bdMn5BaQXzNPXw4DMPIbQf/yu4qdL0L3+mkihiepHF2AXdQflmms3QxBsWM+9c0
7bM0ZYJF5fu3c/Fi3XuQddWRNKrFMTr4SHKyEgkKcKGgg9sBi9EkNNzZqKUeg6yk
/YFlfEwaMtNTwufnZJDZXGTXJf2xKYAFFqQRU+HhkniEy3rZlyCVDy1O3EZM4DWW
6KnIGxPczYFtzYW4l3I5WpiV0I0dACGW5y9rRhTuUBrBn3OofomzIdPkTZ/0AuGt
UeLKTaJjDzGfeKSqygnnw2sULM1d393GyS+b50kNtL6hgGCwrzqQJNkeoyuvGKLQ
2FJFhHe3zBhZjLyk8EtQIJ61x5dxmrCpU2CSk+0lMdtZLJykYmGnPESYwuyCjF3/
7LnYDcjbfuLxC9wKJU0Abt6MJ+WpjI2r2OmM8cn7w3/i2JC0LAE6QihAuoN4AMrr
bg4Fr0whj23XQ+4mCP+w/z55+sUD8+vXmkGEqhznHjVF5aAsX2MILqmkNKFBoGIb
ZWvY6lD8nUxZ08hKmjVQu1/A8nrxgdBsu0/1+8fW71CjmDN5xgI8Dl4UuOlk4x2/
t6SlnkPA4qFpSsIjuGx2QsBuDSMEXjBiyfXWREF0v2gsmhIzjBMgdNFzmHqVcWKU
ok1oB5EXqCx/tO/nzqTHU7TOpmsqfxV0oCy8i6s1egzjYJZQSRH7EimrnKhiR6IW
kmQh/5gsH26r6LgPj4IUHVc6cAle3VRN2weAnNAksC7XyMpIIgKtUQ10QSl8jsyp
WD2Yjo0N6qFa4kM8TNl1cjAT+RVGtcU/Ck4V++sdVPCk55P5kzX79BZMuXpgR1fL
3WI7oJyjMStTsR1CVCwLjPlbHrvqc7mAYQh9Z+3sf78FIi2kVzZ3CGCQN3NcZ5YI
jtQSqVDO8QvzjDLDJYoidbfJTIFXczT3NVP0f1oGoZIUce9zHuJ6999wSmR3TUpv
URYeyEWjWLt/mWzXJfdLo3bzn2Z0Sl47g7UmJHlUILdrtOqteDfcMHESbs+0ij2q
5e7NNbhpF/Id5cSb7j5zOX5inbiN+MW6OiRcbN/6gF57GLBULvEk01ItssaV/Q/z
e2V44jt9KBAPEwDuaXcpr7eQQYcLUvmY+VTz2fGtkG0nNmuAjB8sHx3m3gHzUq6+
vcjBV15bq7D0SJyEPrfOLJU2utolPPhFCtxVxrz5Cr+jYKuhEat3d9KEKTHbyoIF
FK80syoLC7piWFfyYMbTbg+PmSkS3fF/tVMgzdKY6EY7QSWDypKHKyqDBdD0Tecm
cI7rVKjRmx0n1qnmEBtUbD7w91LTFidhrC1s4rwqnPow8IcDoKUtaDE4/koJCi11
xl2NFAEybGls0JLoE3R80hV97Q+heLjm9ykRcTYXhYMK7s3iaPG3nrscw8mM+rIA
54pZug2KM29r2AtokOeXDeo3tMlMmG66ilookBQnVcVUdyOuLqmAsNkDqwpqJASl
b9lRzyGGwBug/axKDqUXuS4PpZ/6p46Qa9Xqg2qqZwJaMiRGWwVNP46IDzvWbZCa
s9Q2rU/Rm2wp2+EpMfQv2cusilcRAKtteNYHhh9Lpshb/YxQrCX7OBgY5JfOSJqW
cBoVSAhvUrzdcabwvLZrHnn0TJ/5lIwF9bFlTQ1Suux8Y6y5GnFvEzGLF0g+02tF
C4B4pVqpmK3vSf9DaxdODhwcYzcaHcoGNCBEDbEuwhm3FyUraDuInzDrPXytGt2K
DoaDRuia6ehgPP7O7FECi2EEWl63thyaeH9Jig0MWRcJs6CEC0q/k99GNlTIhdik
PaAAb51KB24bhtV0AohphU9znABJhb4HME40evwL2Zv0o2f6GlnJ1UTqLLGeRT+V
lZKa5xTN/Kry/Kn42KEE5enWchNxiCFa3hdwfmRJYl7o/1VVMU+YfX5PPogTxzoy
NOIYPDPgCfI2EbpsWQY1W2tjoZSKGQVmZ2Qo26MoE+EhXSjA2z3koTrlk7KWmKQq
b9Gt+jNYNaz+BGkVfEbK8VnBgo31JPkUajYOnlrHwBQSUwcwh87CtPf7uAErnqL8
qjP7zb8Rcc8VWroVO8YlRx1+bOcu9jQMgvxsM5d7O83g6YkpfvS0lB8PwGt3EaBX
p3v/GX2Kip8LO7W6tO9Sp4VI23m8WQiu1eTd9SXbTlht5Xk+y9wliiMhtNmwZJ6Z
GxL6JXlwE+Nk1E2Kk88DluxOPYrdc8v4fjTygbPWapfr295I5raksMSLiBytSb2Q
KCa+zuF5ZIYUH0iAbIZ7LxCCWCLyZWCEiuW54ZjdHTYQehW93Wh/8NJPtpsDPeU9
fOsn4GyAvAFMMX+6HyjRKje8Ba6r6o601XCM6oMPkmdFrJmZeQo8A2oibX7rr7ob
QFY9S6K803QneEhtxhbU6ldO/0vsJ0S1+avcLnSkfzc9bLTWf3uolnVMm+6u4fGY
kuKIZQ7cwRKuD+q6Gscew1tdiLNL3rNSs+jKM0pB+T+OoNP6QkhtYXC608mFuAJI
lcW8o1L0nTprTZYGNjJb6pxe43Wd4h6YCvqry9TrN/YhuLWBnxXLcCyQnDwyzwVB
AFURgV/8TEE+jtT2Dch679xoJQTn1oE5tGCujfoWCYXmxLobe5cMrlWXNSfVP4ON
i1VwPqMuxSOYw13j8X3TQBQ4DIfgShQ/0kzELcrOjlSO9XPIDt2dpoSrq6RI38jz
5CDGz4mWeKzHiaKXH2nvN2PQORLhPIIYT+zwO8hp/ilr5QV9UBJXi3uwomr+omQD
lYw9M/d/gg9efgLyow56KXXuCxpuSvUyg8Yqk/4gjMbzE1Y6HKGtZ3C2qxymmNuL
huiYoowMJzPnG47h8b/poMaYm7tPVxrEM7AnE1gMLiQWlumLb29XzllioxtEh+Tr
TuC45rBPzEfJDzMBQ1Oknjeqq3D5LDd7sawwGcmxtj7RpX9wSuDuO/58VtUvAnkL
Od0NtiuDolBWmBqBJWs9kv0mNWYyUXEAzOU9uXvVH2c6MqsmxEbzpBfWxcMRBseP
MMtp6LdP0vvgC4ZM0Zz35mBwThMEyFDxpxknOKYOX7ARjWTlz8lNTnSzberU8dPs
8ld0vnvItVUgcewqvglswDxICQagweb+1yk7cfKK0xPWENk61mpmxyAo20cYx+PB
mT6O12TdwqitSJ71dh9u+ZXAFQVY+zkDAeQn1pWxs1ruePDq1JPjnXvPmr/OCi1A
pCLRWVeqfaLHzAgOjV7Lph+6Y49bRx296fUApBsBfGwGn5dG3IoTnsEjHSPn/nvc
ilVlsOWHDzliaa/1v3WxR40l8P2R9APoTP6WSMB1tf1r7rHGehTkGKWGk9fcwvEs
/F/p2C77p8N8hT0k01Ow3lhi+cM+UPBxmrsbbETdM+dR2jdekjb4KRMIDNXy71W6
GY6CfVpFRX5jrl7WZEiEu6JbQjgEIEyysV1Rmns3NvbKqmos8jZw13Gx8MgmF5JV
UEc+L5PrTVUmTPgn3ne+Nli1X5ogNj/JquNDarfW8WeJORVbYyh0BDhGLDJNUs/t
/Ts7lfOzUQceT7MdUUtTDeU+DyxKJfo97/iGpK3BOsyRqb+DBsc2CpRCbhswbsrd
k3xRQ5Z3Kf8t0yZucGZcAj3kN1WLV5hTkzBjjALgeoslPIPC7EDrsrpViqM5t1/6
s9juyP/BF59zpwxy2crwe4DsUul40aGglLd4uYj9tLMnOqPN8Io56skJeZeWM7uM
ifdijPuZHH+MW87V0QpIEdIggIWahjxrTYZqflOImMMGbtQyvS86Sj6V6yJqYshl
4NhpScR2gVH1VWxoN2L45/iGcbfxYtz1WA3OElgh28yP9bkYd5XtMi5FHZdn59nn
fwQ3YRnQl8ksoN0WpptsVepJRnmTh261hp4Y/l3kw75qITIJSDLst5jHN7GurKCj
todnWkmzQ4M1WwlST8l6mfhkccbnoxchhP558bBjPLPC+zHvSI1sKMlIwcyhR5Z7
exHiF6NfKOtID/pkT+URKkTuoB2va4Chvh2nPrzx/tHYDvYug8WKZCWg87iXmPr8
z1o4lq9jXQMOfa5P0Buke4yoXu96yMWsYf+wzeTDGDPd6hKDjCADQD8Agb+/xIqN
xFNjl1zo6ZTKme3LMrRPN//rFU98AMiLkIArugR41hw07SNZkGgf2Iwr43Ky0PJ8
Phkcp1QbwN+8l/+6fK+k+HEoP5IPsxpb12UKSIY0aAZOxiEww9QaKLKz/Pv/3wbY
yauf0YZdQ5/O7FW3DpcdrbK/wJ84BBt+DqDtZZjN0J1h2nU/20XP9ClZuMNjDfzB
Oxlfb5l1yj4ejqkPm93iuSUc26jSHTIsfrg9OwqsAgHd1O6BHY9x3y6X8eUKO3mA
mJ41jHiwkxT8zmxx8EEUnjhr8lyeVgHnJBnAGPCCeh4/yrooQuwExDxx7kRmY50u
9mqOKoDuisIlNQ+xVauRuYeZQSIiBI/rT6pN5V1kBrEUFV4ZX3CGGRCOmocZ7vhq
wKpscePLXSJTEK7Itualva0kEOuESvpcJSIe94Frbfb6NJI2bR06tDltIEjZDv8q
Pbn51MmVJ7B0mpx4/YQ6ofYJpLaOtgUHJxGV6puWdUirM2oMEGONCo+3d1ndqKZD
0BQX0ReuMC7K/LrJTkamxEAXLN+enSIjXE3P7CI5fzWShpDaVlrLXvZXFGWaVYB0
WACMxadYuCCAREN2x4iuNBHtRHfUYOeySyyMXsGuCbpE600BJl+IQj7VyZf8KSwE
LcaPf6QxdBqBHa+6M6FHmL4ATyXHaODLuMkXyd/9oul6uaKMqZx8gI54fbHHaOWu
/4OsZLfVxEMhK3XxWNz4EfGFhHILGINpHjZBxVUd35LmFMen1rP79WD9sWGzLGRB
18nwBvfEzyqbqwx5yU56E0LBZAyrdpfhM7V29GHJDiOl0pY83nNmImuxnqZDapSA
x8FvJASErCe6b7VJeRZDLd69atToNjzYlEcMFN1z1p3sD+4vi6bBsQJ8GcqWTUrc
RC/h4KsoQY5S9JGJitITK33ezY2Ax4IfaYf/GFS+Ii7X7cymUodLe9fg8AeSdStt
PpMwm6Z5pXREu69qlpYJ+sKTFb3/eyG0ljkuJe2GH3RxqO1hnK/NoNCXB1NNt8JJ
l7OswJq6B6UMxxmhkpKC3DaXu9mWGLf15jWZJiwYUaUBCESHeQIxVPsHE4igv194
yJHNBD/n9ddcHKUIuTuuCEm1rV8MRu0dO5HbERrCYF8PVjscuqxw1lHTkzWCyau8
JnUrK/Iw6ntGGea4Kji2hnpizCQ9y4zrSInk8Zlm1MI6C0Pxms3/dL2iiPb1WCuT
57wQiVad9EYHbCR0/SAdm2akjEIsSc7wF4aOKn6zAvBxu3KzMnMeVjGzVlQ0qc7V
U82Uot0FXaosaQkf3jpLT4N0qkBxybBEUvab/g7outWbeu1uHY3oVyrAgtH01Nw4
xH4gwf219Oewv/LJlZH/IF0eslNQA3FVYt45jxrkMPp/TBBF1uQLfWewhliE+G+y
bjscQzkDzteAUuRqjvoWucTMhCdn5GObvThEpbj6+dQ8QAZJuijgy3sDirRV44J+
9wjNkOD+6LlcqQdkp/VGLNHdymichD0ctu1HU9XZsJ4hUhVAGSuaB6qFiFFD6tQA
lKXwX3RJsU4jx767g0Ju2QFcZ/UYQRgpnWuc4BnV295weJUQvMa1WmsdaUabhseu
Z2WaBpiZwh0bFxRNqfxo3qa05zL70H46VSoPiECeTuAHsKdJY1rUyS5zN9xsSxdG
wA1m5TdsV7TCE7JkWMjw/tNZSucBtBj5OqW93M3F1W3W5HQ+tR2aRMMq+YYzu2C+
XWC8tqVb3AziUHuGTA2s1ygo5ZPce7CZd8EX30ATvld2tUxJAi+fc5vVyskMt882
A8lR70tqw5KEQs/84vtx3Ds9H7CsgVXeqRo14TDvVXn+0DEtq0wkaPHzi5iSFwf2
454X1TFxjUtNCQ3pHtnGZTkbeH0OXN9WQEQkPeoR5eD6/JOVvJEpwkZP8ioXAqc2
EBEDc55flyn9bWVxtcoAyKprTS+8+ekmAWwss+GwVKtxt2HrE9tdQ7HkgIFQB1uo
b9JoAyOtZZjIi11yNmEMnCVlVqu1UvVGlmno3QOy30U4lui2h8BJevQMCQo4X+zq
QRgY4z3Syi1jsifU8yX/FgxnhrCMK7LKGXHCI06K/6nrWxMkwz+OmQBejqspGh3o
ezTvsOq3uadFKoE4Lh7qJl6rZYuRRyI6vv6pB+3BzHSqNBMMHc539i1pOUNKbSK+
qhGB6a71pWCYEx0BgYXJ+9bK9FHdqSUH9cXghPFfqPB35KS2VAOURLyFlKiZn9W0
fVT1dR1aWSe1bA7A8Guw3YXevHh3G1GPBTJimOVCZC7znb48bVFP0ZMyFc5qdowA
TqML2hbYCz+rHdpq11WPZ/PUpmF8B375mAXfTLUji9yrNan6kN7NHzI0krH075MI
HOnxkL/riHgKY6sd2F2Zr39boPViXMl44Tn/Eutzg5tMu0f8TBDt5VOU06aomm4A
nQjfoSt9KZWcoPYTHAnk9Ka8QyrFp7Gb3FkqhRWuSkQHYUs7ac1oru0qgxPNtXzC
ypazDeNJXQ/FbnqTEpWA4pTBOIDxvG+x3sJvdwv3Rs2i52S0bTHvoFsRAAb/ugNu
tMhxG86aTPhHWZb60V8nd+kgKRA8lLUbnjxeWVkA7ZqI9HiKn7U5NdPVZ4MchEP4
FQpnliMjUeb6idhULGby4C4MnLAdd+/JH7QPQyfvgVFBgenBu6zy11f2RCFrrZG0
8E/HesHj6KVWEpnLmzDS9GWG9tZl+t1/0Rx6LRhorCJI+wLpuyvx0M+71NwNXGQf
vrN4mj/xP8tJW3Gr1fHJIv3MY6Lcr5uYQBji1iX8KrTIAj5cP1flf2P/menerGwD
TOEIR/+aZZTbGFC7x9jzex5ilTGaJSK6BHdLGq2PEBicwSeYHDIP8yWLXFrhVp6M
ZkD1tLd8XBiI5oVSReRWYTb5GI6PXX4M80Dmsw5ZhRDcfh8rdQ0Zg4cDJCHuUB8m
sB4bjxaWZbsEy9mmH2ZahTcW8WwKlWTl38RTbBEeOJy9iMFZL/Lf6/VsQlZos9fW
blo4dfrZV190sEDRtykAOb25BzWz9ML/AnlylAwMsKptN6EbDM6m+BAbZDd1yEDp
2CirMu1Sr9oGqv1Sko3cNTXSEZjViyHLjN99TxFmrL3wErizi4VTQXmPauyS+rvI
wqf2SAXzpcA4JX5OBd4/PVBX/ceBQZcVE//JTkPydyIXF1yXqYjbVg9biPT6lPw3
Jl46kLopPmXCIXPSvrFhgRBVCmQkGEoUBRdZbLL3RwJ0uul6duCe9RmfsQ6jkBtq
zf9wbjr4uToFSEMkUF/H3VsbffDv5Z1dism7QvZolQclcOzKwwXosomuG8jvxEJj
L3/sddXv4SvApLlN91fXHNl9eDBGZ6emT8TXbvEo/FFIlfP2c+DUVc8KDhc5JEKZ
ibfe1/gT7ZYxeJwHjoeV7hMnIpiYVAA7I3CyzmmKKVV3YBqAPvoujhOtcRKTfXpY
o0jx2n3fCNW7R5e7WBrY0/p54ShZxKAXzEjjk1fQQmRxG57nNOnMiUzt6el/Zk0X
TfdU8U77Fu4nPgOzfODW1ZCNd5UWJB1Zjdo1BAEVbeyn6QsKDPK8yPvn8nIa44CA
rf9ajS1Ay11MJUO8s6MfNTVzHbypVdEdqaFmu/hLujt6Etn6Xbc5QGwR4fNy1Ty6
tOQwZWossv2IwtJ55EOTNqTgho5+cIdilRlJIWrVzIRtwwGPoJU2U0UlgpkHXNdB
jcoUrQ/fzlpwiOOG5rPCj4clc5Lzf77dph2CYE8amfpY3QzvCxz+BQPT6s/bN23Z
fNZf/sLJQx+otSprLOdk+lhloWw3isk/nnaxUKDglGC7+kHri+HG/m/HOfGMtJsO
gxiuBLnn3rlMu9lnTrtQsih6Y2ynE4hrLHGbHtJsP6oD/E8DftuqIF2KEBjexZ4n
7U/Xx4F7VFL0MPhelJCY43HNqBa6W5t0Sr+8ewrBBPgbrqgiEwmhZDTqbg7T2rNl
OssZdUYwv8AGck9RRHFMkWk7Ukz3oXWnBCQo933D1sJHCupmGY6ai0mNCXHJgzkT
L5wUBxcDxbvXw+vfxPNxu74CfZqkZeE9Dr9OrU4hSJvOUfBZL8nkxgvpuzZc1lH0
gGeFMU1nXqLR8BbR6ex5moq2QCW2d9rtnzDngSHgcyOJK2Y0vgM/9BHZmcDh/FPt
bfeg5VaaAfSnNqFzyNv3FzRb1DxNOrX7b+a8bZUNF3NdcPF/u1Zsoi8QinRoGvNc
k8/rYG7gTDOnE3v0E4TuQZuiYjaIaVSaPfAbN9nbU3I9B2p/72+ESu1RJ/iavPXV
qwF6VvO31cx521IikJBSnHrjqY3QTQHXM1YJGK1oeSVfQr+UTRyW+Qf/nbSa+TGv
BE8U8CwZzV5OmjQq+I8Qes815GtrYhbc4FXdm8KH449d8xcj7JzCgYkhYURDfcjm
XrXSee/OgAj6q9leqLqXPP7gu5Fhbk3UGP7t34S5qVcFVy7nNZ2H1Nd8dFP52JBx
cTMV+LEn2Ts+VOqnPBGE5no6fGnfk9AhZYhi4KeJ/rYbKre4E8RNDWCAMgqbP1g9
+8NckZbgEy8UdEArcSUM+P/8juN2+MB2WY9F0MtC2a94Ix0qDinYtpyNAIyEJi5Y
As6wl/otcbbNzmHNC4JrdZ5q0Tp6kd1xaj7o1dG3GJNiyFDOjal9QjhUSiIXSI+A
mgK2Xt2c7YyT4IUJffvu38pcP/SnbgNIUt1pU0MMu+VnmR5amT17SGKFTL1N5j7T
UbNe/lp1xRWymWzQ55rsMik6t0ctClgzRk/oKywcNANRTIrAdP+Xk66hYoEgBDBC
Zr9TGHH83Nlg/OsiRM2uRqOLynvZZfcpiW3BhQ0CHDDm0x9pVJDezIxn9cUqiFVb
cX83D1oowj/Uxt28enbU0fnf/97K9Cy1amLm9nN3vGWKGEVE6VfGuXUDmf0W8lEm
Ki0Uq7qEnt8Ghywekw7prKtWAXNC2nHylhkrlF1AwmHsQTXL8KKYaoOUtKhuRt5v
TRIF4Q3iix52brrjGItkBOy0ocIf8lZ22gnO0Rql9V/k6s1aTQSavkJ/rtgElwSU
9n0WSVaS3RUiyQPnigNAYNQhqVyC/4rieIZqB7gXmzmiLJx2XvIDY+Ho3VnkHmJA
nmCLZvihK8Dwv/lC8XA7SfzUOvPbllBwwcwcGgpdaBr+WKeCtxRXH1l/CsUjyCJH
fqgDoAEusDbO9SSQgnC250OQIMfMpPFqK8jVkpQT+Qd3UJnipE0rCRO872P/45RC
Fhjpipc0Ki7/RAUzfVFolbIr21l+XrounSYHM3cVKo1EP3p6pvwNWS6rl/TvolVU
dINqDSCOr3ATNapSOnbqL+LdwrS7tceTZ7o/KQnrtjAVfQsdLH4gO1UuSABTAPYh
7yam8ER7Dnhaf9W/cmqpRcTHN5Dw7Ht0Uxq/JA/eBsIeKnmJ86+VIYiF/fJq29qA
ZHBVYGCNRXSoDm0WVkOevy6z0nbkJXCvHd4W3eQw6JTmENs+VKp/onLwM/mqxyHu
zIvOGOQ50nB4yn5ga8LSgQKnxU0NEzb17zaKRW/Zvqc/JpEFM2IUakqbucDaub19
vXAQ3FXn4z4GxFHjhnBOrgoAYxTKzC9hB6WJQpAXBM3o+7ZbNCrjkCcYcTfqXwGz
F7NgMkqbfgMxK9wfmCt781s3gdwVYrTTlkeIIeJjccrymG3SDtkl6xdZySChClm2
/ctmRL0tQ8bv/9+o0a5nV5L2ChVFq7IIIdrcl9M6rNnHRFHkYtilslIpG4+xljc2
nOQVcDL/+dUJSN/Sxk6HcbVo7ZL7OdZJXJ3f1nZYkAM/mQBoQ0Wwj9FjTqC/LHFS
+5duteEmTYwBIQ6j8NR19FkGfEkI8VyfCsdWjgjaMEl4YGNogTLnfr11DmH6LPV6
9xgxGd30cveNitA5fIRd/9uC/b/GsXF/yuoXMZweB/mS1FPMu+eKwLzCYZP/zDal
KdVL3lJXLqV1YDmSCBW8+dgIk9TJ364DX7JvTgl10f4Js6j59/2FmQ21JiKwe8Po
MOVaKvJkzwKgVX0RtGWL/xDD5Ddsp6Y2C3WQz+sJ1yHzukzYqhWAX2oNrnvcqm2c
DLTH+w1hzfoVoVzggIerDr5jLDk472CB4jXA+xk9fgrYJcfPtLgULToQCnZmjusi
332B4aaeMBpsX9jv7zbkNxM50QFc9PQVhtGiz8RPwPtKK5u/cKnWkCK/jrUVrXyq
kvi7le+1HRFafMnlRKwhOHJ6MWGXh5mw0HP3sWRJRPPAp2OSl7QU1iIdHyxCT6hS
fUdt0PIjIyOE1uND6mptW5Ok25zM55ivRg93CH0Sn26en8X2tDvRVDHsMtefUjmB
6zO+4m/sxbdFet9Wb4gkOF6bvLLu4Zi75aQun5mOBBoqFA2DJ7/kVbCFB4aVmRqb
WkWjIBUatO3HGaVMJJ2jVdQAFBjggsXrgBEZDVFDjJDIA35TPKZjQNUNHIbEbWIt
Dnybc5XTs8hJNgOkI8FigHhW869Ihr+KV9GyZ/f5V2ce6/G8q5vT7h6PUTbuFOU4
VRA4SBHGj+a1BhAKqUdxw01l9Cv+0lvIp9C48hjB7l0+xkhIkKZeImgLDXoEzjXu
MqeoTOnyu29UufUcEznyzOHOU9G1PbX819uYfdFna2hk/GiIwnIU0H/FM4G7u/Y3
RwnMr1h3wQBAjWGW0vZkNbVIkEgIKggVZ1DI4zzaKZmAY3jcIsDGXU2OHSduBv91
lC68ILYLMiwSwpcz3P9XLrb5TrsJ5UIvVp7TktmLSzerubefliWhNT/yv4iUy/YM
CArQptC8iGeJSvpg8sCpDX9KAbCV1fXMMnvA4n3/9KXGDEH7m+P4ctuGtKMSM5cI
paHD4E0UJFZCqwaC8stOa96T9YvPlT/wt+PDOhoIHoioLZ9hDkt6PqE74dwPLtRQ
uDBUpMvfq0A+liwHDaVBZOkXDDVp7Sx84J3iCcGiZF9ZEqQCAQS1C6P01iNx8jwb
n2n2JqUvB8Cg4RQh7+Q69yBurwdBLqc6noYocNsYVNcEC1hiUjnd5iiV3NQO/tjv
7OVsLrxBz8bB3ceSs3+1fNWUCXuNEjyALnUa2ai6BP+Q9BcJsK86SIzqJGHV1bSX
FX5kznsEbt88CSUlrlNxsoSLZCfY3eb13d+DUuKsk3wQwhL4fZdnFOGoNB75gYRW
4lNy+VM8VaeqvS3MzEppY9P6nmlgl7ZiwgNSGuwxnWuCiqpdxpP1BimVG9psHaWp
aCcuZQAwHHIlhCohe40nK4QkhDJXFULOkWjM2Q0pW1xM8f+MKtWmAhv/swbxxNXl
D8EZVNX1S4AMRh0AD4b91rG9sldmeVy236cC3rx9hcp2Ygo4PafIUqzDGk75YQQK
CrqLfWOD6k0aVff4FEWfn7Gg7PFycnkSsO/vBcaNwCcFl3cE4B799CHRKwDXrG9r
MnfjMCEbDUCZrBDkm08J6UhTrSmynNDJuCBEfNWLeP02w8MA7I4M8pRv0DU5QxxS
Cqmy5UuOFTJCgkzzQfDiar3DG42VkA7oJmKfWf9L3SCoyqUetbZANUosbh/Hh+NA
OFJfMw9e+TknYsiAx+Wi39tAPX5fZtHJ/ysJCo7S4Pdk8m4uOvrosvyTwKcxVdhz
aOtp3LWyqNsdAjk09J/9oCu5dGmn9ni07/5PzHEW4D+R7SnTISiF5PnZclEfCCaR
V5xWT4yF03ppeUA7yw2rwmX6mBqZ1jQISGaeIm35XJGsVXdmvb7ZUME+2vYER2bI
841ZzFg8Ae6+Abnd3Ox0QmVH3dMCaFokrqK8sBItPlgyV4dEz/HE6yoBNWdnFut9
XVLteY53zE4gC+nx0pPJk3Kw7g2653zclozOEVf8ri/dWXfbM53111XLd7J+eSWV
XrPFL/lMy1q24MeDRs38dbWK2DWTm8r6OcGMsAFW/B6GSd9XOALacWXRojQowr9v
+cE+jh5+1Pz0fSQvVntHoIx75HxSn3e5oEpH4HFeKEhfd2jphqR0JKdu2tYs8deV
nP9/YkY+Wuju4KNYPh1qPJi9cNK04xaQrttl+tVHZh0uQ9PhPJCGhJaONszdR756
3WJoCjbow5YEERQy5rNTZl7UzIITw98Jmi/wDdF4Lf46UUBIurg0xb4huWxGXfW7
X11ffjrxZUQ7nOm1evY1tJ1w8Dh14E4DYmORb34nO9Ui/G1L2vIVJ/N571Pu5rFH
XhCmBoBgnjA4qh08jLbFRN1iiB7G6zaBCrjiO7FPrHrZrig+zEzNcDCpZdgZGrSO
b40q6gmzRusDVH43bu8Zb6s6FexIiIvnBKyuLqKVBod1CUqYk7k8oKHIV9gw5giO
lynLREktWkPAfu8bgJqAgYqAgghv+srZjppW4ZheGMJ90AIL+0VPtusSpNo2LwtG
SC1poDdZDqXj8oTNXGnOJ/eGrXd8suvsRM2VCu2UJ1W/oMSOD94ePcfcm80oxxQ6
KpkMqN/IRzwPPcbGVmJCzx7Jocv59fboJnLBWWazDtsBXGXNeZfX67M8ysUF2HYW
XhdjduxoCZQ08XcVB5KhgjxFcwuyINHtIi4lugn6Agd6A+YeW/cwU9cEplXVJJI7
UkAHspWh7WzvmwdnDWiEkyKTiMVzpPSPmoS092/IOmTxoZk1MvtiF+6xMHXPojof
59z1m6qsB08yWOBDozKOMelZq2QsdeHtJ6pg9oMphIQ5BpxZJv76bsLAlHQvEFn7
l/0Jie6+TiG+s8vOFGrV5ZBuMD/gfHb8REMzOv/sUeJ+YVljWL8BFfjq0n4zUnvR
bsFoHN/1N39+i9dFshD8e60U0T/ZOj9Y7Cg7fcQ0MvdYLOFrSW1GCu2i47+Np7VL
6A356cXxFH5NMixmxH9HFPR2UsUX4Eeit7qolbFmn1YAKdDFZYHA4ywTrWgSfX79
oF3vUnnitQDR6+Qe7nguTXZx6p9y+bIjUPfWnKb8mUnHj5qZBV0s1gX+gzrdI3wS
XssrR0fKZHBjuXP2ZeG+jP/uHicxDRpy6YBAphPGe4vITJmDag74aOsXv2XoGH3U
stCwDNY76ocgAD54oplkhFYoE265/Ti4TdOEdvPFwPqgLexsqlsquT+uTNS8ZRPr
lwqP+opYJawuJmPVMeLO5akyR38ixcJf+a9pvc2CnwdmEn5DFwBdlbDIagBH3bfQ
nMf1NN7MFr+pe3T9G6v4bqcy3Er1U1FAtjfEboqHxhNMsVnsUx5akoZZQjMSDZDJ
udPsPL27Wu6Z7bN6NyR9T77RzH/1gtyyzm6bV0EyqEGPI/8QbBf20Sr0yu02A+4+
cvjcbGqudX9iger5EsDuEmSrp154UtdBmbn9OGc9pox8vj7743TdJchB0CRYeqKK
P+lETgLk+JabnuuMEXtnaZ6i8LsiryYO+pBg3lrTef0IDc5nxV/57cIsy3/7cI2Y
J9WDD1YF7VSaxnftLnal5fTvk4BOhbw7TbuIdXJQQpDXS+qaxWuZp1RPkATpzOZ3
TEBqKD/KPBqY5rlzny7w4AFFrCB6fTEsG52zGpqZecdz2oUgIYu1tz6miqwOBZi3
SJAbkny7SKiaJWfXliG+kNbU3vKKaiK2EExMcXbAimssNnT8ivXRAWnwCs2mkw5v
VSIM7kB3/AAH4C8w2Ei50giUQyiqNP9uRFIuTrX2l4hdAv2mHb2yMDXYIuj6TCYu
yF4ACOyF0HNUAhu6lf8Hmr33w23Ev2s8evB/AXzb6oJvXccFOhiqBiH5ZMUHYWzd
WvhKks5ccJy9tbia07R1slG6q32mUQTUtIwh+LxHIJfq646cWppmk/qrmZH/YNPM
HCkWWn/SmMGvauVCD35nDvXHVuZYVKy7ceZRelNpl3f+zzovccELOFfwwoXjO6ct
eyj2lzKA2GA0wSe3yVNaCjAXq0jOy6LqI1Gf4Z0W2X9gd59rB9YHm5MGpLIUZnkt
QyVI+gRMOyCsCcTCFL5EZflj/Gr8IJYD2er/1ndYB3Fh4/+11FMe0ZkvkBwRVnc7
ovwHgUTWB2qU0wRDGyodqSSfhKJSeRWejYtGTBVUU8WH/Sh9gyhfbsUnixDs6biO
e9q38oHbY3VwUcUvdBYGkgOyqE/ta6pMOhYzvWZnRFTL/jjv2nvnDP7ILEfVFh+K
VjlnB+3NU6+UKmo3x28rYWromwKWStPlhtH4IpVliRdgC5lhL21rO9O9aAl8uvqe
aaX7BbqhFlEGHfZwAtb4kfTZdwCDVJn2U1RTG38DM2NMM8soe+OPolguuUJk21wx
7iQt5PPDZAy48gxt1JVRMGUP6Jx3UJJnFqqTTPG5Y9KQYg3FJhShZNJXL21hzPxH
BeyaKt4Fv6HT03H9HRXqJzGjR1sR4gW9O5HRLxvPoOfZwvrIvIiR9pPVsrYJ/xSD
KQIbaw7+SsPE/fWo10eYPKnsVF+N5yObQ8mN2PLHEdLRf/kMYb+2MeqiVAwSauu3
9vYXFquGw3WL3+cdOm0KswLmcLlOma0Q/bo16ByzII3HaRWbeCjEHya08CC6zNpa
rlv5mSg/45MND/V+95vQrwrDvUJU81OCjohvK0sFcKhEzgnh9h95o/u8fl85y5xX
CSzX3MTd0dsJE/3t3ZcEiJdH2xn6K4STieLeKLCcD9yhbHV7TJHyzIiAQZZDiyvL
o/CmvmazLExdiZqDhIrzH4FRJYcEWepdzZEYTDy5W88IxAM1BNLbBSMBmaZ9Vz0q
1UuZxuK8sIKEg9n0iOhHcnEIdPCPWBbyki+SuDW2lYTC2WMFAzgdYfWWaOY2tnfL
prF5QiLsKVik4ZPWgcg8reyQVW91ag0MXvBX89+m13TC4uI64f6jJhKIhZIQoe5B
KRstEe1mi2IQdjT4MoNqYAcDPZWrPqorIz74I7Pj87YGXzjkjcOmhs3Sw99FjQM2
ZEeuXaDTtTsDqsLyr1KcQX/K4b8VI0yKpsL1XqPzZTGPaNOgx/0NGT+h83Y9AUvI
0LFtKOF5kUDVAlBjAdYcErBnfcxWISDL26O8hhs4veZN35/VT7mMp9jveiGceMTF
nXZjWbU0pLNoBKVB6n7f2Z4YeISH/IPvNaC3i709ZfYRJAyuPogKVd2UxiyQRPoU
EiYjhYz1R/k3xforM6I+9DuB1J29OeB4Nn//n4vUmaOvk+IKnYjRRWJlyz039u6u
TIC35r8wigtisHM2VhHO+w6dCwneXm7Xiy7J23P6kMNwfM0EwNReWQTuAIT/CMpv
tvbHzGhLO18kwUDb0ZNMMo4LQygG6frbSCSciHYQWFaLpne0uPz/qhWtsdDnB1Jw
H6QByi2bEbAVOrrPq4fZ5LFeW3fz1c+LzyFVkc4/VohPeQQfGTDP2jgpM/AiphHN
4RRZyfkGWsXRJMu6QT18iE3jO9q8Pz8FPKlgAeFdvInMZ+NCEMdtobNrYFYJa9Eh
z6u8OYHOnbu46ntcnoWB4Timv//eJAnreRqTilNnFANekiU3Eoi5Hzns1qb7kHB6
ctTSzb/vyZMFVMIh1uB3jpS/lTcZIJKC7csefQULo0nFS3QA2tw9nvxmAeV7Da/N
t7O/xMxoPnpA25n7ZZCyXcyEySKGDDGEUxV0gk9tSqDZ7sNXdiu5EryyHAYuKtHg
siN++Gj6EebRTmzORKDcbmMjwYULG9ZAI9P+PWRMwA88vFdj1zDl4EcrtVV5kIYl
mILpmZmqhAPtiiibYJ+oWHc9PBWhZVz24cVLsQjXEppR3WSxN53sUopE3jGzUlwc
rrBo7bdDCHG0xvKveHbCmXuAD/P6uRU98JNFlsvRnF9Hg8wA5nUHEsI/tDXDVCCR
cEA757F9oxsT8jy5kvKh4iUtA3XYjCTczPsy0PAu/M1heoXUYXqU1Vl2IVxe8IWj
zCdBc1Utp2tx35tsUY/triLetiD//8J34tcu8+FWFkTSi7b0B/FRTpeWikrfT49+
8WxhLkOBmlO4d8bmQP47mKGYeTgyiiJF4LWAR4BULkEl1+Yd9GhyUOxDytxcYAVR
c+CkAEJP08czrWK5YuUcIEAHghy8xyBFEtAkrV+Iz49nq2NGuVcgQ2Pu+6Rtz76I
J4xbf8DHpPFiE3Sw5okhXoyTkceLWBa/4lx4xeFdtbp8RimeGCPSvByqeRZ5UMpU
BN/EDwbt1j9D+w26XC5lPc2YVJujSLjnlE8cm0kvL1RKaBh6LeplxhzUTAxE4lHx
gYKbbogSoHEJfynP/6qgI4+/X2Tf+NQfaJjB2JW7cckPKlMbiyqzxpOza8HA8VqC
IWApuHCoS7jecIYHGUEx3xKF86ODTpzTPkXlJ5xYjMzEreNosOqRw4s3G3Xnkz+p
mnbwGZA28fqTxydFjai5g1zDLsv3hxo/GJzD1hd865AD8ojOpAFtVZNPlWIPen01
3y0zz+W13vjQYNZ6y9mUIG/MR+eoHUp27tmkjjXNXsJOAIohJwRy9xHQlpTmcd41
t55b69c/Ot8r+YFI6c6DFzEurNG0Pxf7xPTCFd7zBHrzQFnzvN4DGwvcGJutPJ4R
Ld3X+DKhA4YhdxAK07yReVcw5IHHWOTCnXJAt/KU7K5+gTIvAHZ4aRWFHTWqWVfD
BI8CKuWH6Xobne7XFPDztYTabVO4tMaKg68QOWqXRKQUOcAlW/k/JPb3jWL3eyvi
2vIyvV8Io8sROMdQXqL7vsab71KSIZW90m7Ic9y0QhPWU27ZaiZm9G8lHtrhWOHs
CQPQjXjhSy17j+2imij9h7DSYFJuewIsXW0IGd2T1X7no6rJ3e+ixsASN9RQmjr7
UOAY3EydX/pow67KZO8PGRTMZvMhubPuv8zg/DNw1gPymvgLv9L/IrV1CzRekgBT
rfpW38ubl5ceVYgm/+xYiDw9MzMpshgtf5mdosaXNMVECnWtIwognPWPqj3r8FeC
yOwKLuUNTyaHTMP4Y/PpoXOQmlj1sgvdh4XBNBZKjnkyLkLYDCxqRUPzfi1CpfLf
hM0KtSIXGa+9izI1+NcUh6gLIM6fkWsB1Zf70C97/sIoCHQa8UpJqaCZRXQbxRvR
6BUMZlttUz5IdQg7gLuyrxFhqAHR/NzCS5WH06CEHcHi4kvuVNj9B5TdLJFuZ1A3
MSq6Mnh3IHzxeZp7MGujpau704c1e9Xl8wpvQeAinBCoF7o/AFikaEtyoIW9YEDX
M676Wh6eDU563Y0cZTS/5sjkrIws95eTSJ6xUqEhRa+W9JD3XhiP/CMhJTgXzF7b
SkeEye4IQRx6GTPqTRv0UokKN2DozqElI8FA6ki/g18jsaD7UuwYvzkJdfK/DcG2
ZlBoqoJ1Cle4c6sbuw5996ofzoCXW57wWvznRropFZG4qckK6fNsh5mmryUKsRUE
PQQ3VAOHuXNFlO/NJgMUPv+LjgHKjx+tsc24xmy15zOIXypXyZ6ZQWiFn4THPCLl
PW9iEhIwhzxPJPHNi9zcTwOdOOI/OJAWy+wkdRpxMaWqt5YS56+3WJ6OnIbCCqIZ
yabtlP1CpOUl4ndvWy3ZuAQS+yMkADJeRAi1h1t//M0FYp+pmpVFz0fZLz+vLaMg
Zps/TNXFL9zWI0D6vqWNVF+GdaDYkA56NZrd4tBIGpZ8+GRnn19cm5QInDjXbHwS
G11cwHcIJsJYUeaAvoZ2BrLX08nGAkDUL+6DOx5WQfvkBbl3qw/xCMxnqHAjhMb0
DO499htjqe2JMGfOe7ZTKG0sb9TO/0dEw3h+ZlIkuGXc7i/+sj1Qt4O5UzCzlBx5
c5qjNhfCX9+QqYEiIEhZk/YOpS6GQrOPBdqjDzJmBeUtHcG8X983dacQMnY9QDu8
pMSaj2rI/c5//6N8ywdy4tPi5IgiPNoteInzNK6U6CrxdNzIWv9lsrkEKvaJeOZY
ZfcVxuEresOyjY1qM985QYJ82CaIDPKPwTdd8iE0ril61zUzM4zZRJ4FXRR9Wmh5
mdUj4xRYb9wCU8Xn70V0NrhLy26Ry2UZpxYL0rDyLHrLu7D5nog+EYRHVaHCFB7D
DRArTmFjEoOIkuwdsTWoQsXksi9nybVe6IhsFk7ajpDidckIF08gWy53s5PpfHvv
cKPtbB1qsLUVDA7a9KY7rWXQN0YSaYxZn6/pgq1eWxgyoW/ZTupIuc58l/OeEx2u
j6UoypabJIWG0/9DSfx97g9HHwBt10WjUwN4ubMb0I+mkj3UPdTMZhiLT2jmLbrY
ZLqYP2JhzTlZpY6Ld2wKGHJijj2JKI041hphUjKNocu0lNe0DNoMeGdlSkCned3M
krrEPX7e2XbNJ3HMhMQeZQrhx4BbHRVWbIGfnaqi+8twwOu+k5znPZdWqeTm7lfB
gbqb8kNZLKQ4ceNKUkd5A5NOY7uVCkwkF1kH9pijhQD9Hji23zI1z8sJiolm428h
Sphl2+E779r0CRm4wp8f8ZiEmCrjf0TXRQDRZFwFeatbdz2JrpkwjC5kqcgxzn0P
8m0uN71itJ1rl1t38JZjiSCrzecDgw/EZLmT32h2kCbhYQG9hHGYkuNNN2t9i4VU
TYpVWlbTGImkEz0ssviG3NbRS7AdmfMoFlxL9vwp7KHbZ2CwdAZSMHbagRBV7zkI
XEJhMGmy4aipRdsYpoEdo07HPuNvDGTj2vfGjtcji05eFgkaqSIA0eKtkSs0kUXa
4/95Lp5RyQEzFo/gVae4v5cnhkEqtpuuMZ/glAP61unKX7HCer5KVrxr6Oq1Hoa8
MO27xit+r2w39OOa3jS5Nt4WpFpqDjVvTlOu/yGiADA/8cEFzl5GPX7Z63KAy46F
zCJ/JV7RM2K5K3oZPK3KWj8zP/2+5rot3v3eDtjqbizRwEah/rZOrhxeryzc+QE+
hvboVFrYdet3083ix2mC2ov01igpMIPXXB/hY431V75vC9Fliyab+u+rK3wZDPLc
9tST/nedvxPn8C5a7bSlHXJyMSIKRtXJnLXED0yDecKLEJG6lreb2ae+Wr6I9UYX
ov5Oqzsv7NKr333lLXt3adFpTyOSulA5mPr7AD/wans2UzercfXCsupQ/QE7yNBq
N03qBtxIVBpu0xY4jmeHhOVlBykqGYyw682vV6K8rxdj11ock40L0/MsqktmYCuN
n+psc9fujHPmWTsZe3hxu+qjuqqNwfT27NPvXempWpnxvLsqot7Nc5rKNSmKHvbx
Qh1fULx/EO4vDuCRZMaZCGThFGYxS+9kNHJwkqZH4si7gx7ZK62RK0CU+6bea9OU
Tj2sPKkBl4n6kpVNA+WW39vv/jr89Oc08a2RbJmJcNZX+aiIZm/KL66WGnkNX9sk
KZY98LIJ6EhbBhgsVGNcDzUiXW5a+VNmu1EsLPApiTyhUVBM0VyKv+SJ2y1ixoyU
hW8nlsAW+S56jhOCJY4GggzHzvuFkBHiWFej6K0AnAaw12qqgxdA/3MoTj/4TxqT
VMr1Z6J81BTecZ4K5LOx8tuQBQgDGF6FpMZymMl9O8lrAzJRbB5EDSxArxzF7Ipo
oiOMJimsGsfcwIU1nNkphhIuEH6uEVCi3AaD+nZDglpjaeR+xHEPzutp+ugXtNCr
kl8RwhE4WysPAUWPUrunrVI40VnqbdERlmXiPJmcuMCebXN7cxPjm3U4IDypSOzo
Fkly4DXXuOumsDVn5bu0Bhqt5Qqi/tQsIa8durNJG6AHV/NrYrZtpV3fdaR5sDCY
3ch4Wkon2paX8gFjK2ocsYS4I4FrSBLJ4Bu336XAyc8LAa2lSPGpA8tyACiwyyUP
0wpNd7To4OHSaqZVZeq8A+lH17Jw9ccSX8sWcC5DXHhklpYzWBDmdORY2G9XyZuY
lbv46QWjbYZg97AvlxMJ1MPK5Pz3R/mlYqvonTVdcFdNqtiLczJtiqxlkMZTzaiT
xJ6gg8PN33FAwf/QXBW+oP41RRDGX8SzSO+yLciLgrFU66VykW+LXDqfgtnSadSo
a81307fRbsFu6cyZKog5e3UH7iMR+eLPWbl6Niaqk2ElL41uAEpVPA2u4df+kxCX
SibopBuRK9/gSyrvIzZsrDeJWcKW9BXa6R0xsxIfUCyLDzn2nwJJlm6hKSZU4CxC
I1PVpsIvq13UE70+0B2jLibloLY55uDwSWxbA460luhiToD9nOSJ7ZNdfMGNF5/C
Y2vYTVYp4AUWy8fDn80M2J+YnXuInQab0tSrjbxKRBm5Aa5Hw8ydGSt2XBo4CbOA
s5HiAnIxR4Y0hbj4cZSgr9gzzS3s7JiafjWm6UBC9Rd8X70QRjyKz8Q9fFQ5oN8e
xMk8s90ydgJ60o2ilqUfi9E5XRBCtJPV3g/8JV9JpHDjRYgOs4YOW7f7N4eFCoTi
itJAa78L0lAV+oJcxSCfyD4b+EZYtmU9hGHnywscQ2d95t5VZtk/3azJ+m6dbl6N
4Nai3JtCFTtdAX+iOnxOb9378Tq5mh+/QuZ1muywnT6xlJQx7hrAhV4U2aFRiZ5t
/oX1nHiP2HPBO/cZTLmlUrPBEdV0kz0XKJ5vrzHMn+2cj+m1G7Vh5V1k18pltGfU
cCYGOzO7rQCp1YJ/vY5yAU+o42zzrIVOIgSyBujA9dd9CXxywj0BnX1U1EYJQXMb
05dudZCIXwPD+7COKMu1zg+/wRBZuBfwUOBJiD+Od9HQQCjmzP6C6UabQGW2P/e6
USwH1acKZoQSzGuh6iG6zSTSharmgNh8ELEW6jMYRw6w11KnTuPceDyvaE6V0lG4
akHyt8rHb7DR8E7/E1KIIixhY/tnj1ZgjX1QA4vN7j0kg9zwb0b8pSXiCIQUWaeg
1Gvbmj/Y+JR/oPVZdrlcggpHRBYLD0xpgS7iFEK4kx82Tr/Ff9t32y97dHNEwDXC
Ic6Km7pLk+niy/Q+cM7qD72XN8FenWGzX7LMydVhysY/lZsMbjY6d3/jvIyjKFg6
mFq1TUJRodWZaGvOko2/8ZaeRwK46B892vSvM8bZcihNTb4MmH/sJ63kx9f38VSN
0siLfWDua/B7U/JzHpkxQy8JJ6tCsigV6hgz1I8voUfnCkQ+du76O60xvE0XjpdJ
2p6swlQxUaemqD96VqHkYvQcB1mOq5W5gbmC0zn9BZbdGtB4j+aJOR3dtkQkJU07
QNHpswqiqTQONP+95fSPJu3jnvYVu5qQF8JOAKQHbzStAT/trqaxGE4Fg68erM0D
srd73nlY7w0U2ViYO4Sl1T4aKJv/b8Zs37KA6Tr/Zl0tF7f37cxZXogLBAFZTcff
3fKoJMljrIjoLKe9S0QuKMzrZ4WztQCJZHWPf9J3jlsTeu4UXB2dE6pXKEabw57o
KGtA7vjyopLWa2C1WN6HV/kHWZMJxop7dR+dhHVtZXZjdCRY/RyxrYXNcTpxNn95
cLFNeT4gklN/xeCadK1/wANK5uWpni56xzr6OzDDS8nc8HXoFGlni4pMDfLtGfVr
BnMggKmT6WGJ7klz25eR/UYocb8dA1/Ubw/O0UOn0ZG6AnQqV3jsNHc+2bg7B3tl
AXQ1PLOVF/PKXj5UY7gpmtGYR4q0zpbj2qX+omoOr9lB3gsDFCi4QeFKR58dUXOL
0UFxy2skAV6o6/oDNY10wugEHLQ5NgKhVmAoASFYfQkTBYz+NT3VcZuzWVoC35j6
AW7Qr2ESSeCBO3pJX1zMdX6COI1sCUgv7os1gskNFvt/6T5Iz1rULEC0dVqyT+m0
aMccmXz3yEmuqLpeNOE9wNbLxehZGhayR+/TqF4C5L2fEcPMLlK8Pc+iVsWHbjcx
O2it7uKpP08SN8kW9396BqKtT27C4wKfzcetGB9l3cSOLCOVNGhhik7LpPLfLyoq
tvv0MxXv+Zsu/1ue2KjZmnou+eGkzxkT38KXjXHmPqxj/wwSOJvXgtlXrQXVZ7zV
ekv4+GemfN7hemsiew1ehpmrtPSoJlwWI2BiF2AH/ZxauVyWMBC+d17F0VHKM60C
VyXshhJq6ZTInEKyNWSNsUwQhNnH/D9LBoqu/BTC7BbM9WQiPcqxtBCNfd0VgtHP
cVAOdOugqoNo7Ka6CB+jCROzn6O3SRlmnV4mZUllmoesP2CEBHx7iTILDxqhEEd2
fOHy7H25nSjPFafgNrtjxrDViqQe+W6xyoTFjLTFGNNo6bitceVxKLTVFpNMsbgH
MaESOsN5WLziFzPKWsGHnTH8V1lBYe2nnCjFO9otXecVkF2qZqQITRpsplO0iWRq
1m7kZrFSkyBKOP3Z042xClzYPIw462DYBxHV35wrqFyllNC+hOJzm0HWrUZYfRpo
feWpn0afSKvBVvX8UrYq+4EIw1bHDxNZPLiTgdTqD9HtmJJwdGTD0jU/qkNBsgix
SmhQbRCxFVPzSi5mlLgXDgaEZR1S5YICYDYUqVr9mjyHUwdEjgmdGAXw9RVinnIH
tkcrIlRu1OxF41jPgKHmEnvFGJ8SHWQCTXXztYfZlgON/+S00y+G1RxQ9z92YlhH
8bGE1uK73KbyBoEWfuEQKqg1U/iwP+vkgjR3e+gnMryIBl4URAWoXGgTiUtq4ZR9
OWyxWOs0H8DG2iQBjCcLNL/Askm9IjI12pnld15ZPj18L+LQaVzd99w+XGBBY9gv
bQh7pog9Qhu6akPAA9rh1YbYrp+/5N4MH4aHFe5Ge8EWrYlcv6Aa1//GtpSlr/7z
6UQw434UUUEF8zFaXyraM0YEb5Hed4vSdcOOtMQ2k78HDwgG02o0TlbFenCFl1Tv
QusEKe1iVGJy1EV+JLD3FGh0ejJkOBFiNiXAGwgOvbz+o60BHwr36xeyOiE9vDLu
LI9bu1bac02H9K8ymxJA/vWmCMi7A8DuAyeYHObrCbwLmFXpVsT7Kxav8IAbEPtR
0XpuP2GqWNfxB246lmkVhfoIZH9jUY9F/b+UvjcTpljTYtjI6FnGYcaaDzkFfsID
kKjTNhimaPkKdOFY1DGdk31WBosDOpVTEmxqOtnVx55hPN9Qjzt7BQtXzL8w6196
vtsCqOUlrmxnSktOVTLdh93e6ylHQIcGriVRB3zF+Axoa7kwAIoouEnkf2W7AeJq
zUauYrBVg7Xo1btUeGzXczNkUvF6R+OncBacIy21LpmKb/XkWkJxQnL7/G/yzdKT
jOnsy4KpfxwR47UQaTRv/ZfvDWQMvKj65TVpGinBseCm1RLWOPp3uhUWEyjMpWkI
vTZTkQuxFqgjESKlAjAIefNS8oYUkkIcl8nH0Skni+CP7I9dTDbPNKdvK5H8HVtR
nci0arfY/FJU3EMGLg7/4LSf9icplbeXQ7/F3DTrtt9RPT9fqiG4Jvcx5plKUDNM
2q03MQRdCfj+QN1yze3zoo/6sf/hFeumun2KUykrLJpVEGAKOaHRCpakEBGsh08g
ElsEqNwalafLobmx0duky4F3LD01pg8DkaCXmAe6rARWe/JscKpe4Ze8vd5zxXFb
7Hg7iSQNeEy8B0kYqra+pSeJC7pwZlw+b8sVctzfwXkNvbf3VH2gLLxhMfDfnkxE
MgErLqzLB/mfexmwRRdZUEy/1+3vsZYeYtE3EVt+HXfesFMnhA1nsckGeHSRima3
7F0xPAV9M1xyTZM0HEBQqZ78Y08dJkeogUrIX/s8+JSdGVaEmM5gqjjGQRNDsyT6
vhiPIkk4TdmRXcEgzZyfs6WunL9vU5YWsHTSgBYvwH0wW4P9HxNaGeuBrssHcvri
Sy7zcsourVsXpVtaXZ4bePimLGkI2EAPuKDu1R5nRTZL5UK6l519DjfeNfQ/ZwZP
yTvzD7i+HvnMmh9YeJc377dDsIWrDhQ+eJ10C8hsFcJevrf0u4BKcailQ3krBIT8
WMgDfkquWwJbHU9KxoKTxaRP9reB2Wbzpa2/+djM4rtJZpeoW7bED2SejSxRXLTn
Mv8wZnOe0uVSD7f7xj+UztBFKO/vqCtyCXdGlpdnay4BbLt01uSrYv/aHz3lApw1
Ca5Iwyk4hjMhTuy4CPoGoG3S4cTNS6wcGjNeDaYblmjSFqKf9d37GiGp7xyVolgS
4YsxhehJFCNoDqADb5aBl7RPgHhTjtihIL4JYhwtfJSqf+ikKllrupkUcZp+8aTP
kqwdLVZ/RcixeE4AypBJwRg7apu0gWRHsCOgXHj9hirTHH7zIcncjfUvM5FnjCzA
ZUIRmQBRiqRiIMt8yCYafnHpIZVb0mtxBWL6o9nBTDzt+jUUANgNIrvp/+pmEIR+
EFcoC3gDkLzum5hZ71axFEZgL/uWCGtto3NfbCTHJL2dxEpxvgIYjhlvBvZrPIGF
DHgAX6/EoMruUZqCEypinESBrpexs9xxvX6py/IJ+nC9XAmXTlpPnQBswRDitjcC
yOa0pfFUk5y7Cu2s2uDNa6Iuxya/iNz+RTzjSZafM6OBB68fN4xo6KK9DDZ0RjGu
YMYUAcX8fYdWwJ/YcO7g3HoxAPwEQoQNChHyTRNZJkBLqyteWFqn0Vv3baq0fadU
cTAjnnLuYlQRQBj4Pi3cRGYCQL2tp0N889E9Q+ZWOdtJkjUdpcXykgNAOrp+JJ5K
ZEL09mJKlRv+goFjEx09QhVd8Cfv8bBb9fMkQoMX8mQMZI6gT0ekQZ5k2aRy7z+A
OjEVduuuRDHngKP7sAga2gQmTAoTKUVIJk+NuzXX7EPfdUvnpGuORsGMg6S4MyNm
jdM3utVRRC1+yr2tLJ7b0nTrqwNcXVM626e08tzdLNk3XYGoMfinbjn49STAGYZJ
fFTwctik8ghWD7nCS6G6qeX/GkX49xLEUX6ZWvc+ucTAwX9VMSMH8mvRHDmhVdUG
0AnfG8PMuNkh4fjGJC+06rVGvlYdAU5/jyahsH8wZfvy059tuq9Znj6mdagkEImE
r9VS8ejxStCZxpBbzfEVO5msNLSNd867Z61X4Y8E+uB+BW5s3RFJpF7iA4Nocq+7
unPzCI1Kn89OHScHO8e0w0nkesv5dqoiJA3AEXIVp6UinrGJIxnj+7c9PR0/RYoR
1ugCBbSUfzHbgg4H5CtfkJDmdIKg9m/kD+vlFdo3ZLaCEjGJ9BqbgKABye6UeAcD
qYVhArjB8uH4jJjBlcx/TRr9t1MNcchxVyXKbAO8nVIV1MqS3z1TRYHUtpC0W7/F
kv45OI129quSg2+SIT7LBwbuSvgHZ0h24fTlo9qGr9mSh1I9hLQb3UHekwoAaT7N
7Rwzn5pBmdJ/5N4Ai7arQ1dbaBxZJPu8Ef1+4ZG2WyEa5RMfcYWCld2YqcSyIhQI
O5i8iwKBRYMbmBVGEb68xYeMYokI37kaKS8i4vvuzO11RyVQ2ZPp2quELWTx7rSD
UXuJ8NUGSoQpjggAB8JXyGsNUBUhnyo+d54Ck8xWEsfpp5Kz86rbtV8bmqKra0Z0
aDRMSVVwe7HujaFTCadgj+8PpS8FGr5w1GiKS6DlWSUfo+/Ub2QX383wne1m0PHF
GZ9zvpTzX47twaHRg0JziTfCAoLbUqwCiO69MqwZHOHk8lSDvXTvGTWyAY8ssdsr
DvKb+TgC3J+koIUZwoKDU7ysibkeh2ZzLVCYQmvHnY6f4KVeKruZOzAl5/Fc+g9c
hBodXheaVEGNMv5spX5otPb0e4jEiT4WGXiT5NqyVi3ABLsE/90fBB1lVS980RbF
vqBaTJH9mwqmHkbvW0XrgbCX5R2vaXO8GgvMQAk6wtcn4imee9B7cmQaMsT1/wkq
hiSQonbTTHbt4jjeNbgOYcS6u5e/1XP1yM/lRpFO3OILzk3WUXlcAI2/vyzyZV50
VHSIc9v8KyiPtKmFk1vEq5mqMbcGxiCY6H2SxDaeqO4hE1udPYeR+i3zSxIbTBA3
WX3gREEXSYC/M3R1TFs58FYIWsnQEQoj4gJDilCcyXc/H2ZT4ZuHyb9cJ2IYK2oy
jCeQ7K2BRY2A8BSQy7DMF+Zv87t4lLc8GEFrpjutnJvzp0+5ZIGojB19iYYvLRGY
dbNauFMSyo1sD0+3x6xtfkVGJKuJb/IFX3QS4cwEWVtjFEUL78C+usr3hYtE3lJ3
tYw53de3xbw5LHOrwrh81P+P5AMZQzKig40pdKNExkd02Zd8ojPrMXJWE890VQY9
+a1yHIBrQuA7+bziS1cBYGpUtjf3HjIKCVrikgKIoxltA9Z3CoJ6wW4Tl/O4FEZE
711cd9RFRxJAuhICKR3D730Y1N9EHVr1Ws86qm+TFfcSNqrLGhjmlutgVDL/Y0lS
v5CgGRPepPO5NZBiP1y6opjryagBOQoEb7WvGeTmPPTwNlE5qKNFjDvQjg3wWbFl
sdde6Oygx78ycVdtWlu1VpGuTE1L+YEp+wbaGLU3gtVQ/hS1Y7jWfXbQ7NIfAURm
eMyV0G7WWrmjMn7uNt4Sk7xYdKbMZwlttB64VzDrkOyb79RgNoOrLnhcnXaYIVMH
bCeHy24jv6QqnJc4r1/ngTKxiN0iznmXhYNkQV7YhpkyRwFiy1A6xTivol4HAWLh
na1olN3cwoMY8SMtiVIchCTqpe56ATENKSerBY5nx5leTWqXvlXiOT+S8afNh6FR
+4C3CodkckgT4lBSuI4oetAciNFMYQ9uP8vHki3oRIFzh4vlxW6Bn/26Sx9WTQnM
aG0IivSql2q0jjCCUZVP3gRh57KFQ9WzmetiJvBgScR1M6hqhXx546DZ0jK5x1pP
gXo6JvkHIvoD/uc7S+lnmcanUvQOLvuUo2vHU1Ns464tft6d6tc8lmDyEkV6NgHH
KBlD8wnjlTkgiKaLCTKM9rJKW/1oAdUGKc35ogYd+dpQ9lT5FStjYt1v3nV+PTgS
`pragma protect end_protected
