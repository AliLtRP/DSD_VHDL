// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YSBPVJC+4WMFjCA38E827waJrtrpHFTmAeUAI/vT+HeP/emAYf6UIs43pSyPbUQ2pjuBROoXl9Wo
x7HjNalgWsweEn5elcSTXSWJNhjEpo5NwLbN2nYpg9EpuXKp0ENf4O9g7jOlFAyaHzbs/QaPxG/S
In7fJXqKPV9nn/7cyOIErV64IxDtOPEFt++tYkCGx8RCU1iQEuQhFetJD8DIwa5rzVA4kxfI4ITh
RmfvDxsD0YzL8yNxFBowAaKCeuI9Dkh9x8Y+GrkG3AUhkmHHjaEJ7LyeV9mIqIBjx0pGJBMq251y
zrfqc4FC/hOUmmJkMkOoKXA39wRvuDnvG3oUFQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
HbsVTCq0Bj0Pnp1Qb9vbPZSXeqbj4qJa0tBNAcG5MiJcZV32XgSjGsTAeQZhll+jA77gxi6DA8d4
E6lT2xCC0S23EASXL5S6lVdFGKdpIkjjn27cVNdGLsyuy9IgjYozs26u13KqLk1mXcFw0cWUNlLx
+65mU16lOAF/URqUoT651nk8yKS6AgpVmQlQ28i7snvFzN5NEGyE5OxnNQJOPHcQoPbxbWsEtg41
TR0OWqkPztD+SiHca/I843CvRWa1g6vrPNmjxuJEYCa0sTwl+NmSa8f9E3fSzcHidD2R9SWpGV03
zk9D02QTmnzFuKzhgvVfrhNbeBiKyFa2RXn0u2qZicEVboQsZqaJmw2oMaBd77P08JG0Y0aHBhOd
JDe1VX49h4uD5HtVixPfzggjEPWQ9tji6hwxUy9okGUyXSR6jBtT2w3UDrP/syWL7tCeCnR6JSEM
uvzzRXiixnTvVKqLOLVStmG6dRKMhqB/TZjqDpCqr/adByFqpplAmpWkuUqEOnFwNDAMYmzwneNd
BXOLNKbU1m1zPUZwxis+WjaeUnj1NtmEFXXeT7KA0IO0wfaFJLBXHINf3i77whqfCS2kMCIksU+h
bnLBEYTGDY3TpIDjTXO38fY8pFYVLEYw2MGp0DvtamCPjtVtViFFFFPov4Kny4dTx7Ju0mF678ue
9oQ/jZnfa/8hDAud0WBIOa/D9QInpUzS6gYP7SOm7j4xZ24gcWgmCKy2VTQaXBuPQ5EIsaA6KsN3
k52akLlGmeUZzR41nToM30TxdReTYxcx66L4DqNd+fhzigvhn353QGqEs5+BJMHUpGyN1hH3T3lB
Ede61jRW2Z94q5DoABr8wHiwNtV7mgl98y0kqIuZvKt0CDqnDxR7KHwMnwAo5OmsDvdkmLvbNNSb
FHm3rAlPx3OaztJmFjcfhvMs2OHsvwSs2nGkMl+7F4hOCQYt+f3jIlDCMTlkrHUciAsT2Y3TSHHe
3rZOKzylkzw6C7UtDYWGG13pFb239yN3SJy9vr4xYa5k1aTGFmVkNV2DHLsUlu3EhKQuarKDVqC0
VMLXT6gL1ohrOFRSKfwPdhZieqFLRnTqcHpnxEi1MMjOq6+UZclAqYYQUz+VtPBMqumpj5hqRYan
IkYQJxPwrDltoGVM5BdM3Bi6n5OY7VFW4cV3odAksKwwu+79Sk4Rb0ypAVGFsnZCBj/qBJpfDGlA
XVkLKW5w6SugOxg5e2UWwn54tABc+/FGYRYHPil6JVvV4E+z3TT4Nq835RvVIK2BSRHFLa5A5Lds
6Mj6Fy+wFJslRNnbETDai3+zN7q/iaOPNATbA2AP6sRk0A+FLFcL2PjBSQa8OQTPyG4r2eHOsqkW
+iWAi7aAoyH/Vmef2AGqd86A0REV6lLhoQNR9UgXczzq+AbWjzJPzBQaKjS0rL762VCCsf/UeB26
rU9ANl9uKROXOJcU5DibiiyCgUWWkn9QQcB/dphTf9gGek1Wet8m//d5AQNoXthEPKQ6dweB6j0O
9omQWIu7O4n+434FKGpvWgXx2OuKsutHji7Qyhwibj7LRNIq+ETk0d5p+BOz7FDKV6sYknTYoECB
TNizHLB339rkVP43yTy+i8RbgjSq8u18MyBflK/mFE/zjOm+8d9utBz/XZdPpTUQqTkXmIGoJCF9
aDbf4VV9pRZvZdUBy7So8kjZmI+cyhmV3PlJVo+3RpGNihxU96MnhfzpjojCoC6mrffgi4lHPnhl
MQQ4Gm0ByF0VsN09KiNWcu4Ec078PS0kC9fzmoRLLlawQWvNnZkHW09jPPw46z57DVCfLwk15GzC
WZUYDGeG5PJmmW3H8IpGQem2nloVnRZnoOKGbPeDQJJXNfiyYAmWsgt8wIV5msSStIjRm7MfH6VL
czSm+8phsqtyQlKMeHPNxFWP3ZyTb9kgITMGA5QGjuY4Yb+k7TznIyLXzcgJcbOQQXhNBpIraVzV
vu40viGLJlaHVD6GTzd7AupQBi8gui1AZwUaR0K1cXRn+Xca3Q7aW/0aUSRVs+lJPi4s8+oROpWE
BFo9WrRJjc1MhPtYwAgqN0raSjyAlUIuU6Cw9/daGnLjJFsSh0z2/sZMdfjynZDRbAxE2FjLauI1
BFl4uQw9HRHqtAaKhr2/N11OynGhddqo7wMwYaKHxlPtkPB63KXV1eWMtYncXBbtkkDWI2Obvocr
WpaxN8Y5QwKhiuawbsPRQfaqmbwrinJvPQbcIq9tr3uOJ86UPKV2ZXnskT+RG7QxcfeMUgEWWIxo
uEOzQRfWGl8l6SxJCvFTzmgZ5Z7EvQLvawRP3Bd92hDZ6xF05dGahQOgUhj8aNG99/7KWXPKigZ5
zIGRue38N3fRF+xWyCOkIkGQTK73G6GY0tnPJy17vGuN/5OrzzWtD1EiIZpRUdebpnzySVecl9zk
1XuQrgDRHSHEdZpqcIhk6DoWuV6fSRgp0rvgq/qKaVrIp7kaMWjBWjYAPVEEfS1i4ZyEoUkV2Gl3
PGbHZMrQehVllMnwAHPhHCuHrmJl8Dg+j87KUWKiOT/C7OxQHkaXSwg/rCgQJgUyOLfuS1hzLcSt
OXvtsINYWZ3ipjzrSqccF7H4MY46sqcA1z1nDthqjmrOX0ri1gUVxNtH3yfJ/vPlEUwbbBaUx0Sp
zbFTfJ/AAxT6uc1wjI1msPg638RguQ6T4abwHBfTwFDdZ0KKXd7M7/vHpDJ53xaJ8X24Luz+5mfn
pUSBfRZUUx76IfTXobtuHsEJg9xtEK4Hg/Z0FBsQ3bseceE6cR1vI45smdViHyYOFlEqtV5KqZcB
2R6EjqRdHwpcmrHwe1MKw207dYXF2df/CaSHe7WkuWjg4GyxRxsiUj5sOu12aJCB3fLI/rrGoO8e
FcmleJm4PqRz61NIytorPQNZB9j5PT/KDi+/ejlvWoj9VMKGbfh+sRKsbdocDGxV+60bfgmWmVwz
qIJS9Qkf2O7v4eQOj+gpg2NgxqXVHRQUDbMN47hGxQ2v+j4ry2BjXSro9Q1EgGKJA45eJvWrwDyE
/L5Jf9ZQcCgEQR/3dQbPctjctPaqTviC/YOB+Xgw+n+2Wvn3El2idUztePMn4DGF/ZL/BhKhibmU
dXLDolyb9cHk28tL89qrXM96C+RiIDFwKVtRNaVa5Iy9GIlYc/Fli8izJ9k/c+g1f2ebX7n6YXi2
O5ue0N9pRsKq5nvzi3NcVV9DAxRSjUZ3B9QChnLk5IMDuT8Npit0/dyXstPhVG/gWgCsOiKszO5m
tf+jQZ6t/Y+o9uPFjFNpPYiZgAFxLwG3SorBC7TW+0Lq34dvk1c745SOAY/f1TeRIF43qBXagdWL
/C1HNeWGtPEw3HdX2UFcW25Phw6W18CmQ5u64sEmqDdNg8q6Cr/6TWnNU96pxyZfo3loJl+UtPVV
xN9w11uUQ3DdQorfxIg6sIkVwea1ySFFYNpNdvxwY9wz1I6cNewlFvXTILhYixYBwZ4FqgeGpv4l
7OhwV95NniVnaSzvv3TWhA1IvNcb5wDOAHo8w7L6wnvug1VrgF0LndhxSJUqRIXQBOYZMWXHNN6g
zjmHnGsz8WYqEOZMx9opf98r2IRZjNpaosYVOo7rR0I2d011B4hmn5dEmD3j81eFQlak5Ypd0yDq
EEd2AOloc9w+d04+uhHENzK8llCROyPFdVVa8Pcy+MM/MfMzm+uFHJw5+Tjo5KF1BhqJkEDkAyLW
2rce/Sgh+csid2o5VSS3MYXiH502tm0phD3q3bMFTbelMG0G4K7Y6aKLTYqGT+K5DE2eIl5QODTD
Pr0VT7ZjW5X3nHyyzHd9wF6DBZQsZq35H/NgNP3lhXW0qrRWyqfoO9WONhqJup4kLbRip8hfx7bB
jaE7JdMyyEH3Q1XACCHjTxiG+DnXwZpn4f2tHgWrlF41APPu8TcFsF9NpotaTFSNhuGmf+xOW3Tt
3DqXJRRNVfYXOiZ/2Z/47FeTLnC6IqV3ofmDcNon1kGSamJuKSKvo8UBhZ26VX3lnbFscRv7KaQF
l2ehOrH7LeU6Ptr1TMlGZX+cBNiBujr+HoL6e+HKvtsDjY2d9HOrqn3Tv5zfimhF7GvfOPSnSEtt
9am24pfVrohNJQ7LEETKNx66QuFxIOnJSoruCOHtzVDPKnu7s5pWOQY7xtOslYz0sAjNwm9aSho8
59qD6s6a8H9EQeAoM4y779w3RHQrpTQAFlKBK0+SCmjoNiL+emYxM5LmLpBQ2F97BSfppY+UbMaw
uaXRdzR3jjrUFAmLZqV1V6ITm21PDZeS40E4qPVSxniYpwpXdSqzzSMkrn8kfyhVIemSVA45aKRj
yfTkqg6iLZI4KGIRlRR8mNcp282fZ/+iK5nAXa7EqaO3WdRIfy1tAD0NpfUTf/3DweTNoHPTO7ME
NiYer0WdsFGLisLs3Ur/+xw+IUEgNFmwdTd4t7DHv3tOhZ3k/0F46HUt24T8HuzMnZJ+H8opDH+I
vaD0i9YJxykSsj1voJRdUHuETXPVLSyNiw90kZZS1FdFB3bZGA73q+qWGftOJdBwllVnFVu3nQlC
xM5FjUUfF9wBA+VYp45+iP4I4Flpu3U3M0rW3C5bRUAwaK/ikttk+tlZQPg9T4X7BPYzCc+kIuW5
gVT2V8VMy7NqsiKQtWxDtFWaUHYOfPDEM69AkA0orjux78E8yYAt/13aaB7ovyBVPSsFvaQwJs78
+xqQQk0T6M5HQu9ipgrxQr/3lLq0qvs3h1C0Owetmh1cs9SteX8c+4rdXR7EcS6Z0m2nB1J+6DFI
fAdCObXN6JAXSyEqmipBe8QR6eO8ClvGYv73NqUdTOjU1j16J9vOap3DHsYXY4Mz3Opb+xYGSq9M
XDHP30kElMUnOjLb2qqm7cTIfjk54TNvUzXP2PoiPKBpgIRzjFuUlUw4bV3KFjaKSadbzOUdSvH6
X4YUFLFq1BcD2exr9tSKch0n+SgJDyIJnOZ7jZgxp2mhnrO6PVasYYalOMGMp1lX1+j7Mmbq4dII
nd3Fsc/hII5V+LGOeflp5rc7p/Aff+aRClwDpBnI8fKvVWjHFdRf1BcdavVOPtOarw8/lOZvAAqp
Eqp5vwzi7oNYsC0R3y4X4EeYxoeDgM8rFwP2MdhJXKehtwG284wSt31iGH+pH2jlqkxchpj24iCm
J6HQmr+hhYkurxt6tMOz2zIza9MhSRK1Tu49VXtKUm+D2GCiXGzmMUf57BSSNAQ0vFQoYHZnQziY
egfuUo/WAk2z6eIlh3ApMiXfJ6BcilxzQD7TZ34zUmRHNuYm3Nui/D6ot7mRDlu7iOFMJb4Q8u0n
cFRKvu92+FbGQ8G2Vb6edq77Jcsg5vpw//p+rzdru6fZVpSvnz4XMrB19lm2Q4rn8pjDlheu8SPd
7Wr6Z9ibaR87GyKIUqcaGzbuCFNGzwmYHeb9gZ1GrocrZQ5JDskwc6Fpd3WRMUE7QP4WURmHSRau
d6Dn2CAChFwzYlsizC6X/rKvAZcyidGQhfIspJEuErxdEebRW1tH7IJGNOPl98izp2vWgzhiifRL
rpH9MWJdnqzqx+dbfrphXfGAOQgHDYHNHEevq8ZXEpk+XHlAtR783KjVsBYz+I50mbcZVTR+UWZY
Nf5RuzhEsG+NiRdwqQ7fYZLeJgi8yZa86/5Fo1SnLrxacGAFbsOVKJdxXkuzjq7TSF+3PR1jO3hJ
NPmGUprGHkhKlkdlQcXG8LyNfbT+/yCrcf4FV/M6M9DwybHpP1xOOyjZofHLDn9JMa/gz2RBJGc8
4wSgmUVbw4cBAUiXubcnnXg5DFlm8rOcuYoDjRB5LDYVrXbxI63yKfamkmJgGjbspyY4Z9pDOqnb
+VapceBKfcnZwS16WTjj0jsgz0va+sCK5CMsaUHme6PZgELODXeW5FEBDYm2NND3emOayUjkJS6X
/saCIhAuqtUR4P4ETZqAMbOGPEzHM/PwSMUuaop1KOc5wXQF6XxH6CDFBuYI48igPBN244ALtHkZ
/gyUa4Uxr/wvKljeqLz6NAPXt5KU3q/xXcMOmC16XmTbo1agTBR/w8+eBeWpp2uMRvXUfJfNbbSQ
VBFvwVGW0fdmbAhsCDPHPpSE/jMxB5tvwvKmdV3vwPY7Iy+iibPNyDtcFLvum7n7AHV/lZ/QX3V0
cKaEQaq+nAoGb4Cga52i4IgP3aR4CDUbrOQDznFksjB61HgcYbPII6ENmrPsLKrHazZxiHY/5QK/
CTJ0JLF30/5Lu/n8wpGNidFYZsAnH2BpOcNcIp6RT/PvZco+1GVgzUSdLCT1CJTNbXsZtdCFQuOC
iPobng+oKqOPSeYAHGdDWjRQk0WvCJaR6Th8s/c9ck0vL5H+3WAugx06a5al7hfHCZQfzsLLFwZp
/b9Xu9ekM40r6Sx3fNLlduYGWKijkHTmwIXUpwUFv+M4X+7gMctWbR33Jgfz2QS6ziqgYqLQYaCE
jVYLBSnF4OBhhbogmcg7np1yGR/cHBKQ+o/ibDFvDzzs32fMj3uMnja+WjAeAl0RQMZb4j8J+BB1
iNYU+80NXbEEtvUWRqRIIyj9oY6HFg5KcvKuKTiajySo7P/DDMXtv6eeY3cghsefLAKUjc++9Ysx
Mzf9wgcPuLCF7HHjjH2QF+LVmEvRlt/jOsqwlcW0YAUHoflEC3Dl0kRbOwjXbIk+6oOu7Cc9M3x6
1UNtEX5dghCLP7GZQToLb8vP2v70GyxOGVZFgxiUlQxjMxlY8XLNkwTttcht80f73HJt9uUuM7qw
LSKZ2cSrGyeepJDVwu4m+6hNd7fOO6jrFvvATq3n55Ma+wxFP8YVwQrX71Yqag3UshQwibWtywvG
GdIa9EqV/IWsmIzfMiEhDP87Zh789LifrDp2MmaPZhvFPafHNjojo5d6E3Dd7lOoW7/M+pt0gPry
Hfz9tia/d/ZE2z5qKq9+Nuw9jVcz9VIiOsOX5VMuDMqOfLnSwCu6FM0k4HQIRwER5pzrrrimu6x0
A4Gz0NdyVDItO1UdEYdbCk0VqfFAnq8s5aBXh1n9rvYnhlOaQYauJp7pceKbOF8IoEhWR+Fxq01z
dryYBMo5UhwTTXL29EwD2S9uAcD40wWMD5sIlr6RnLI8qnUX6aBwjLF5DCqH3mBhUam6fhWzqUN4
pyRHUwuyUoL2HknYQfQrJS4MgiIcg5j2hHvx/u56rU50cYpSTqaMqaSse9ikhZt+LCCiXeLuVHYj
kHftZNu+TMIYVHapOT/DNJyvY5XHyt2HIKPdzJT942Wbo8wqBNOHB8Yge3j9qHHXNZHo7ioX/SLP
BVV2IPdJZhgC63+VHehTtf9U2hxVoDoXE1y6sF3puME1jtKmqS/dDiZN9LtVm82a3RW8GNKrcaiR
HMLKVmMnpOczJrmpnoMH42nM3rwPehuoenZux5nnSfcI5p87GIkNiKsfU4JYvKaiLbvsjlWI68Vj
QTfX6bNxBVm/KYlDorA7B8zd1lZX8manoR7YaEqec/+8UpIgCsUF1UCCtSYY43b8on2cCuGyhQqn
BGBTMX9rIboVoaBPkEdL2tNZyZubHfLYiLn72UVdQ7g5JC4q2Urilof3tuCk0X4WgQExaffRlE7t
Dc8Ssx5//xR+OCLSBkQIlTvxXoUAtpeM9B0iAFI9NmikKUYn3rf1gnaedf/OPlkXa9mYglcHQsQY
beNl1KzuuJnyL9nY8zdqtWQh7NogllIHUbcrV5raQyJunSNvEkNhY3iDhIuaTjJJyvwoAQYz0QPc
oD+ikJGwcUxj/dEshhgwUnG5/Qq+mD7dr5TnNNhFFzfDdLwK2v7gwKKHWwZHV8hzmiWBp+2XhRcj
Dyq/IPkh8ZidmKIXdLhQQdkPAPnDy2/EgZUgpdcxWKIlO1lD8h7ZWUG8mvdHjNiH/ak1cxj965s9
NuXpxSj2z8kSgrQC3M4cktppdITKSnDzrPgWUQKgENhNadjRSFDhksu9iWA3haRAyBH3/YDkyogC
mOzZAoVED6lqDVeWKMyPv+esb31wsu53BTB5hIPrHykRvNjcGtPFa7SGdI7ngXnV0HvrW6I+JK4H
7uq0jTk7+bHOS893vuRiglUZ9LdTL0On9QYmwLgPV3xm0wOGNSuO01b+dWjVZ+Re0GwhgPgQpp6C
0yseUoPW0Ssr20/TriEBFa4wpWDXjzd2xWcgmEb0IXP6W1hETx8Gq++xf/Q5ryJgcpBCAlVuHWS9
LlJDp0ntk5P4i2bcW6QxeG7Ng8TjEW3tIYL7KmKrB+3zcZQQK9bgCsGogR/og0LURx2YTmAsfJYm
MO/A9P4meXNNfMSPb/4zldJPWKrL0tO2vJSCg3HcyJ7vf/2YATo+0ez6RE6xzruG0gqc9xfPxR4s
PfOr8gjEFGOEDmDgyC5J7CJMpwL/ZqJyKvVa5c/wRcdbTSyZxP0LhtG289G0lZvOAwBMGBsBvYAZ
p+RynQRMZbWAUuCifnx5ePdTh2DWgJpFG8zNjEw6z8FB2uRMib7PAaTWA8rwfBD+Qt/Fszzd9vfO
Rhyd+nEGF2tQxvn75PFCk8ggLQpMkLbWAzgPQ3K3u4JybY2L1PNNgUL0ZJv397vcYWMT03zHqUOP
j+LRa5mE9MBYV9jOti0kmOPyC6BBl3PwlzNDs8hLBheRrq8ZMvxifkTtL2nYoNLkePfc1xkiBZEM
hp1j+X5NkxrCUk2MtXT69slOM08+eGKuraNlvEk9Pa98ECVoNWNJ5eAcB7DNgI6avznpMPDDwuug
6JJpq3oHQtdg8dWmz4sdqDe6+U/jysRwFS0V/g8NAQ4VUVJBWYV43fYJyMF8d43vkmBe8FoiHmUp
dfSLWre32cE9LhyrVg3SKkaYeiv56ySQBhZ1wj/EOYXdtUHx2OKalg7BLuLDgI1tqwjPgrHkN1wB
v0KS9Xlwhv8qyMEGulkgTTCltUNh8AM8WliB7LDZQyA4NDK+Zh3tnwfleJDCY0eSWJQsdiWBeS37
BnLECjlfHKS7ntk0znpqixazlb7fG7PHRDW1yIFaKUktfkT4qwl2NLkuK24qo0OCbuVEz9SNKZMv
4HsXDdR8aW7A3BFK7CUXsJst5oHctgVLo+uWm+Mg00kxOKOxU/YC9nrbeaGxLYd//HOQ6r+bBiAJ
/Gr4QFdoYI6xGBRsNWJWlkqlaADclYGrNmov+F/s8fWDZY6I/UKqwcCNLkv25XT3gHuejjE4wXXU
tF2jxrBSIksVaOv9rWiktkaT8swJb2VIYUHv3/ehuZRM4D68DRXJCYtPdZFYq9h4F7NrtTCIZWE9
A6tvOJDYqTPEmry1RkOmgoUBcqlE4UwY6TKU5b3cqDzn0TKHZx5KYV9waIAS3jqW5ZZacxhZE02R
GJIvF0LRRTCJBUN2CbdcqWsESLmJVfnDsxvtbD7C/lg7oncPM+9E2G1D9X7iHL7v4A+JHMULf4EW
3lPG8B7z035FMTgwqdCm822v8hJF3+6sPAgZLNi//8Ll1S0BT3NHtxs4eyZG8jRJ9Z8/Fo80LZE7
xIcJs7i9lkn2TrWTXQg/hh9LxjQQxftmI1Qf5K45aj8ysuHmDOQqbmUjtn74cZWr/oG/pfghHUpd
WcTTLVoqnc5achRJiK0PfqHlGJ0VnwYGGL2cTSXIzY2NISJ1RbcZC4M1iGyXSMVxAGrNmwtnaQ7c
UTTSf+iMqGbXZe24AgV/RlrJCDi57lgdzh0n8P6laEEDQPey9OIEqYxwxNzuaAW0fpY8WBbD56qO
thR6drx7es+Mr8QtPkAPCVMpyVW0eauPz3YQUbe3o4X9LrmWH2lO4OjhMZEGtNfUymkD0X77y/MU
avDWgMD7pChjRZj72G1suBUcTxybnTzWE8KyA0IebDYIdp0Lq2FiO9skWftN9Rb1l9kz8b4U6qjE
a9OARjTn7xHzA2lCcIj4oYWA3voy4lV7eArwgx9gTXuAF+8WVzCTi7O5LFQmfTxXB2g0xwc8bWPi
IwOOwluejQDXWQJAryoDzD/l6RMRbx3bcLmyv/1H2MEMy8JOZtScD964iik1Q3pDIVI0hZPQal1c
3bQZAnU/Se9hUrAYR6h9teERkGeXJYALMvcndE2RPER6aV8mWTJP0s4pukVx8j9v67GiCPxtwqf8
wQBs0fDBpjRXUXYvXK03fBtji6iXbCFe3p2mz2JZFzlXDn7k9p426PnUCf4TfzmJGlD0SUB4r6sQ
HW+C4FPqCul0GmmBcnFUO6RJcEcwa7emxF0GqFX70VNjsMEjDjseMmTnIT+TNM/IOnI3ekZ8K6kw
N0Xzy8hW7s3CcWj6iXYaZZgOfExiUxHB7c89BJ2f01/MAZUmRG+HTo32ssP9OBacP2i0pLFzkkRF
XSoC9UbXJixc2vm7suBqhNQ+OTiFE2b6goEPjwDLEEhODnna8rrCV1zAm6D3gQKQ6yQjtrZ4N4ss
FUv7O/Yw2N6pRD5QCxYgFh/wM21CQT6dK6Qg5sr4fNX8+U1JGn1DJ252o3ey00CrQbvCgX9eYgtA
FJz40HL2cm036vRzfVusvz/fjgB0dVlfHUcXO2DneWGBh6yMMnXtUXmd6YY/Tsjda+TqH49mksRJ
BxZjKBG9Wpw7lemFDJXR4Ef9tAsJbCmJdo0N27YjkgwNMrLxLu2uhV/5bY40/bpmlD9X/IbR+YK6
HzodYrEi2ohiMZ3R6nOQZYOFmDRJeX6WrH2gu5oUXT1LM5BKb8n25/88h7bU7P2jeEMSia9if8G7
YIU8Z5UuAg275W1aIq5ueCFldpRrqFnbqYc+FoKfTzGvZ026KHyAnrQ1yvvReZF74PReuD84ZT5q
a1b0RYuNv9ARUYVVIONYxiNiNLolHy6J7fTgE1K78bB1ptTuWqrURFarJ3dbZ3kye4BHFXe9msFn
cIXcIiYuuSZa9gVD0JWXrXeK2nM4UDMo9klWZUUsPoY6OQNUwLQJMSXGTIOXWj2Hyb/j3YUcyv96
vuAjUN6KsPzY7R/HmNDVu7OILLVvQwguEoAvUt5hWj9u0madiVP0BHUFp6mo9Id7zO9oEEXyDtA7
DSKGE/KaHNVpxHYAPHHL+irnuGigqxgPiEcityOlN1lNcDBHLDPr8v1rVt1E5VQ0SS+y8gJWjbNf
BMgc8ixPCdjaAw77L4xWmk1tKQMW5IXiQd8+IPqBSDs0yPsDRcy2HTtgoUtaEodMUUszo/rXEhoe
SVWkdaP/eTX6l0t800f2H3YNFl4nsxRF8vNYnqyTOHbiIBLfpfncpUBMjbTKEXOz89XZprLLVy7c
iXBzdIHW3ldDEL2MAoWGq3pE/xfjStVxbmMIZYd2eGehwqJjMyklqU+yKNuCCKmmumils8WnjBE1
WiLAlR6Jq4cXtiJpnSVElPmMWPZoOptdbc5VShdOcVuh4ZCLUJijdhqSxhSa2BUbSNf2SlqZ0SJv
r4baXtO8FxluqGZ/FBsV4ARNQV/klxhcgjEARnV83sSlMRMLkSnkwaIL1ZtIAdVowlW3acjP89c+
CAXxJfmm8ghqfpfZa5JzKaI3jtgJh59wHGcBzRAY/NwGBKpG0CN7BZiXYST9/A0JWdYioc9bR2E6
4GqnRgE+JwjkXKLAy8D51KaBC//JsYRUNRNaS/6ZRLxgBzgvsXvLriF7oIGz9cf0HR4IzT9x9EfH
DQPV9xbdLSF6aS3TXZ1Wb0QnhTfXv+/LzEOUPPBhyFxYvFkTrkSjKXOy74CxRmQ5Cae66iU8kSe6
VyHREuPs8WbP+WIbAzb+mDvspoixpEiAhdW3qkp3KCTR2sUb4tp6xWmb6bo8iwNNKFDDvp7KzHQQ
gqS9wdGFByAFHR+CVtBjF5EkUD6epayeuZ1zYuLHMhR3twvk97foGroxioKtDOl0eXADUrS6FVb2
8KApPvnNb50X1PTUG95gYaKowrfYzQj4cXNp7rEc2N/8T2PpqOW3qEMQ1p2iqOgFYmk3W+EVnrZ5
5a5XxGm0hR8dLSXVDH1/Cb8Oe0Q5IgQVBi0eXx7xmpX5bzgw7DDhx3/ZLyvtoyqg6RWczgE3Mskd
jOrNkFZXqZbK1T16HOFWulf+XXG6gMto1KZK5hFxWTZvwT98jUtumE389INkPzSIaLpjBfyokIBd
gy5TQEpuI9JtuNl1oJO5rh8j1TUVUPi+51tTiQnq/wU9w5oYZ5Ve/xJUOC7ARHbdPdLMdW5qSl4t
Velaeg0aay+Qby/L3fXMuy0XqGS7FEwynwgl9Do3TYnWOdUGnN2VVBr8NoEaxkWeFgVrI386B1+h
hmfFvrX5zxOy7gzjoqLXyYN0uK0pkfrXzxIBNHITzSQWJCcg9DuM4DsKhig36FHAPDe0Ln5zXaWQ
0Kq50HjtP3MA5upon48fVDg8JZkXQeMqk5STsoxM1D7kMVYDvp1K7Gr52hahNpPg3K2s4Ku67KL1
gGZWr8NjHc/jbQetrUK/vL6rN42zZAXizbYnwj+9aTUbIjRjMag4q+aig5HwCBlvZWAvA/ZblYhw
s7UI+jCPIa7JEwW05hHtrWh7iRHRgrUseK+0Wei7qfutcH68jUJUs7WtLRDro1Ou9zWk9s83ZWc1
Hv1AWglesjAFZSCxYI1McWzE0x0l9+O6hAn9I/owjAsbUn7Nl4uu4z0R7/xhJgjBJcC9pcA//YI4
VWkKb2FnmyvIfHH+nQDdAjzQ+etmrw3lhSnoLjvl2pDNOclwzJLK0aekJrvZ3AmvnPWOBgrkCzpj
SOo6e82H1h9YWfGYDaci4Dyfr85x7LtZ8tF33D6KF3eD7Q64roAwe/q7Ok3iztMQJPPxIJi4gAX0
4O4UX9nghXlu2ijVM0vVDdBDWEUHDNJlLlpUR6O4B5K8U6258uLu5PGUs67vqxdnPagvm8VCm9JJ
pS4mffawEUER/0KVrUYzb+qAAr6UMYeWxCx5hggCDJ8seQj/IjGoPwq+4VcePjjzcEpQPB/aQLSy
6YwAUAlObqMqfUDQ6KJazka2mmUqvKlBq7pUILl/PfiG1t7qX/21kLPhhtqaRa4zzh2HRLnZ7bn9
XQQmHkBv4n32ghhZFgjoIxz9NcoKlxS7kNW4FYCgm+OkjTDakcfIFzFqfF2cVkfH+QSCuRvF49j2
0VuAT/9NoUp4E0SbymmNtQe5VQoHlYKQTU02a/xfjfl17y64SEgkpjtJul8idOBOCDm+NY24Bd2p
MaJsvGlytgSwU+YpMM2Nnsz0QpJSE8iKl4XUmfC/HTh4JCB4A+xVWHJkS6+2ZHcI4ZDWWVhMe2Vb
vSjGC7H1Zyzhibl+LLeNJfVVJY/I7x//8MBkprlZa8VBb6hX9ndmlSeDlg1nXncNLApx5lByi9Q0
bvxd5BqNM3dZnonQDVfm22tsaHrQGSBKrCfaiXTYL1Diu/KxTI3KrLPR4yicprHRTheAQ9xa90Ac
o6PPG1OnX7Rz1Y5pWrISxyu93laG60fy/Mfn0h7iWZScBuTEu2MAIlh94+inG1d+WJl+ttbBbYRP
tH/7Atpf3/kswCRFIYpXqaSvptq45oPcOzTnTDd5wPCunQcyjgQGDjay1YZ9hnxm01gDu4F+G6kZ
ybu1j+bEAAqd4rf280CWbj2DCB0+/b8QQj7elvf5Vi7jlLsonPpdhzxHrZ8BQs2zVGpQ5nw7Tuta
1QEazzMEFbRQ7Y+CiMQXzCcM9Akqfv4nYGPlCUm488TqVU8k+zNanUttbabgYtMeb8MNyLcDFPh3
9qJeU9rCB/5KipdvYU9ecAqZp5CWp65uCZh4jE6QRDqAI5kGGlhvJVrKTMtxyVOfA7v2XSQF2hY6
cxpPDgLb2y0/FehEoRoyCiirYkZthc4wEqz1y7ST+spsWgDItJJobYd+F0zjdeP1IG7oVQ6fG2uR
lAzj7jcZOifw9GT5JQ9zxO+3eWWicaWa0GFNXKmk97OCCkzRuQher8cfwBk/VMYw+xwr0hB0SC54
63fbhHj7Op5BEaE3bWwButiQSJXJbRYunlz0oG26ZRV3s+fUoukIE0/akifFEkqX642Q0CQDR+e6
jC4IpkxeiwEMfx21uPa8uqeMwifL1Ox9YSXMfUgTEgyvcC+cbwNQJQid1JSqzNJqZXdalVSopQbS
hrzkA32nMqMuZfh52BXPcqkcCAscrMdvrSwl1fXZcmtSDqqgxztOQQbVZBBmC/Scf9IBNxLdTwYf
JVA6O+EbWuT0NhWpigu6fYCcs3clU4tRo2DLgigCum8zOvCPSEPvISu1wh5k4LXU8JRD04gFPcGJ
8ezFbg/Ymn5ecOClcN8PV9e1gsibDPfR99AJZVl5maYS2TxtNxUcRhfjsOIF10LnLgIkg8nykRou
VfnDkTMSJfauCGqwd4q7wMjzyGBJENlpbt/ittjRl4R9NWEgx0ZfNecXQcmD0RHcFuf0+PcaDItg
sePVk38rA7WPZGfn9cWU07jHOw2dYXaZsMzIsOM8Yfx/nRRfy5yd7Ooo3CiSVzw+MthSu33sbmSD
2kMDZ/wVh33HAIhXfh7hdYsJXEgzhZUEbEgM9kTkqTBznD8uJGyAD69u3oklzMvSAa9J2CF0LsyB
DA8Ka9XkCdgszdqdWLS5OJ1UdTqC9OSTxTbxGjXGYRNLUMSzpQ3uaG7VCAYBVJiQnbp8jwui/Twg
7BpTaN96mOlkrGq2BVJOtDjlMU933NWLMA5isP3CUDf03vEnxhfLXRRZwerlJUFbA/Cvi2T0RWgq
k4LDFwv343BFiV9uKimY9Hjy4HIIx0tcqasM2tsY5dPdptTsoahHNnwp8M9C7dzN5XR4kcjK8QU9
8TaGipkcXNs+RHiYrPQEdp1YfW+AOAdQjZ3etGRTYJjQtCcg/ieb9FQniVhclREmD0lmInQ+yjln
Yeg+hvsFBrI/2TsjqEY70wJ/pPKBbzkMAgnqFKEsNtonsuSwjNTdP93jbdKw4hFBhOCipkOKSisZ
z4KDw7Suneg7o0kiAyA06YgCBOqC8eDxcdBfLC46d9fU1QKuMCbzN+aH597Pfw97RMQh/ravq7gl
cDJaP4+P6YlgVlPWy3PH6wxgp4/d4AuuK0y/Dc90Nfx+ruEmvowjiePJt7nkYr5dJYGhWx5kACQt
PQOcGCtH0hVll+EZ7kUWzj4xxMDeNLyt/ELkY9yBIJkY8yY+GZbvsnBkOqDsA40cmjJHp3RqZei/
6x+aVk7QCBgHWcLMoet18+iB+EAh6Iob025VrlR3QR4k84AQ7I0KjmUAQ76saV0r3f9s+4yrFhcQ
EygD7gxo2IgBQ7cA3kRoK9ZMgCi2K8I9hx9MqfOMxtVYpqQDS2NN5RoeqYFBlnJyNj3LIuABBCtz
PjzeuvfqiuaAU6wnhPeImVi/vcl8O0MT+jw+15pRYYnxNoEsjKoA/QPFbgT+mXS7pAgcdPUYqO+/
w5qA/an0LlPd8PAqDhKaKXT55RXEpyonYoCedWikxaCehIbzswzbQXHu5iLrsMo+2ZOYBcNrVtNj
vpGZw68aMpzx0MScvA6TyFV8BaNW9TP9Uwu4/OD0Y0umjAVmd6QeakTBEuBN42WWinrn76bwPtsd
l7kSkrj/SNYiqDBGBSTHAVAAds9+Or496c/TI87Nu9aQqoCiNuQz52iczS0YdxcsXltDIOJ1n6bE
xMIUnPJMF1qJEoX055vJHBnAIThjAClQ//ZPtPY1Rp0Xtiykw45IiogiowBW4Ge2Z31loNte5X6Y
0cndzV9ocXYDPd3ZggCIPUpPExOKHbDJr18MXSC0hw/r/AKWAcAeGBYtJbqwDX6dorOQSk0qtCns
T4vaNYEGqQS8+HiVKQeqToY6cuNp8mrGwKVhU4vjwrdeO9PljfZcK3t/P9IZO1i7FlHYHDJcPCfD
jf8pOmkxKC3lS4BRE1yqKKSZmVmYuEGWLNuqnBX5zrNPKdxXHZD1rxcVTTrhn2TydzEnf0ICn4FX
g3BRJj8q6QHh9881t2Yyh8xTX7/90ZItfH7Pw4Qjvrgxmt8ZmbxvwqHN+R2E4xtA8XjZfD5ti5Pb
j0AQAK6eNWdtY1wqgoaRSZJHlbLrNHjzcnlWVy9O0KODph0nfa8tIz0o2jUQgIZA8rdMjA+kFA+u
vgrXA+J90UHFEmGNF1l8EIKK5WgWxDTFm10Q0fNycd+QUYGE2ZucxjeBTAhavNHoEU4tzlVZziug
7sQmfjYP0+ezYrtI0BHz3/PQ0cuR8lXZk1VAUJvYz113GydgCGkp48qsHuDmyG9CddiM4xLflBx/
9f09iRfu80PBj7yy9+Rt+1MDM7/UZO+oj1jksOrvO2K+VCc6+QoBaKzpqqkcpoip//QZQKC6IH0I
sk4ZXZ3CkEuAmtU7tS5DlZssIoXcg9dcgeSfTmBPPLLC6QfkU86voblFiBdjF2X1JjQhZ5ijtvAM
jPeJQNo+9eqttqIIt1op1X4cWuRgoMqDPNiZeBvaP11rBuP2ajMnsG7S7jR1wTuCUJQlz0eIIMm4
OTzwC7noDGOQqfZsEP+W0HAtF3O/wgUsNm4wB8LAHxxLQXBfzOri+blJR2Ege4ueRXfIhv8td7tI
5+zLRhYv3Mog1B0OgZ93IKnpW3mWhfWjPpgM+/PWypS7cDuov8QJr9vMq/KqgKnv0htqYVeu4TF6
Rtpxr/0rwvUywPON86xv9GXNh/fNGGzYxMYehgVVTpZTaMf0005cQuqy6BuEB7JC9dLB1vAGZUHz
jzsiCeQXWg3N4mjQQhvCi16kZ5r6bzkVctxh2cmOI+WMGqWjigscOw1XANeZxDr7dNS/Cvt2zhHO
oMMSY3UjL8mAoT6NY0Nc3LeYiEyqDTm7ZfaTWjvf4DcqGfljggAwEN5lOZ+kUVPGQO7CyULHzfTf
s+Vrcw11r1Dcyps1DDIEr3OueqiteJXaiyUyz8YnFHEtP4uB1ZApagmf1FfhKXBCSlS6A2o8BJtF
bI/yM0RHIVym4euCdiw5Qzv7yNYLT0YxM9rY4vdUYtB44D2wjtdJ349hMb8Ehi+d5vGkjhxwE9d7
aYy4Vt1M0fsah6TM6ydrg7V4TgjHVyWWOR9OfXluwR5pDffmNDTDVOFa5vEUO5DiBmvPtCetvxsU
WoinlllhgIGDR05FmOorYrsiUzuXD2cyKtRvHMqpxGUrVXZqDgjsn8EXCklM3yxhRLIGJvkEPiiQ
VZavUfSgq8I54rH+JJpsvmvD9tnPLIkhjohiOfEsQJayMa+Ae/cg/nftqoi65ndXaDbtbiTBnh/X
GjRVkxZX00M7NwgtO1enithc/K8+1kyNsJlWfuHk9fL/ITdmoN5TN7sR+Ri9t4rsMvJ1sow9TFHi
qSqWXnfw1LuEk+Nkromk1IGoVjRzZfE1HUO47iEf0wJlgoWh95w76JfvDPeNhd0JrupZ8wm+n7Us
GceBTFQoLdDaIhuDRTNqVkkv47D+5QY3EyJQKhwJ1GTQJAEqperMRGh5UESdQum8h/0WwM7LBUSF
F0UGWcTILKktFxi5LQXP3ZtgYbfbNx3xCAcCDRVNvBRzXXhDTaoEzgMfRyw5jIWs8WvSOiD5eaXs
Oo+u93euJax88ncm9KW0wtUsNS+YhqqFeQYBGEVlV2KMG7t1pqNV/Awozg+KWI9YgEjAUbcfAhwZ
lGMSW2RN+bSpHhllCs4LIaj5uL00WSqn8ebXM8Gj3SaMcULPEascG5om/EZsXXyMeCNh3Gl0O+AS
pSXIR3PEuo31KMJG1I5BGwrkd9BKF53bbt7cEV0hfNrq7dFj+kn8e7fuAC0bcatAoa9j3w7X4jPj
2rkjIOdNibLhbDXU0J6EBFKbANZEqPN35l8VzM3t020SspPoOM2tJlrm6D4Qx1sKDnnXm8w+9J21
4+jmhImagIxcTv5aSlwgy0utzNY5b7/AE5QYi2YPmnHJ/OlLQhEDmmFYZnWteLQZXdVbJv8Bey14
wzX7q6Mmg9Xi9R7riozuqrfyeI2ydt8dT32HliIqW6JLeuI6SJQ1H+v7dja0aU1I3U32OOnCC63D
MxdPERbRytfpEtNChNtOw3tVWW1hYH1UGOuk6ld+KiTnjErQEjbw42HVXMR4v7qApXCHU/CzcV0/
5f/nVn8MSNseG5TsACt5zZU9BOQMJZep8cz3oFTrQaT6VUC1jn4okhVJde42R/FmkzUruJ/2o0wR
os8/mCFGijDsA5fqEFJGYB0xcSxWfVRKEkLlb9R9cwPcz2pTIrLVuIDixOwqlkOdN3p8I8TINfCV
0JGGYWvqrYCCn87oOPbOx9q8Jn5qRCe8/qpH+fjeG9IBUYX1YOWTHzjGAvMvDsEmQMYTfc1CCGQc
lN9lmeJ8syv9X2NxBcguyx9RnCuz0aibWKoVqxat4E5zcMv8WqkyXEtEI8PXXn90WW+MsDqnP/QJ
lEMBI8S8t1VTBqmPqdQcn+uw6yeoMPnyyk3RRpwxG25Bbe81OL8cSc0Z8FiSO5yD3J/EW3/OS1tk
KGxwdGckBGfv5ly4MrFfs5OGKRVdm1lP7UkAKJdWq3PJeLR15WxhZ1d9fq8ByF7qZeoHszRaobPS
VF1JXLgQlvyl6AOvm38VZbeoUlOBsYGJnoA1USYdZK7MfXW6CUZ+cUbiMII8/NF8B6ZCw6Nmmqo6
CP0FN6hrF9Hl5L34UuGeDbodmCdfgMmuB+QU2CIOfJpfXUvAN1Eu4iSt6ln854BnFLhh1bUlwkuY
oKlTpwyzWM/6jzKBb16Q3CM56iIiT+1fqtfggooaTMkxVMue7TGTu/VvDASyrbBmF0icG1YoDG/8
6F9DpbIEcEPJXuZPx72KvLsUfqZ8fGrsFqTztfZPivDF+m15GrnOk73qhO94wNSDUUPW4ixlqhss
CIYXBbWV/RbYpgFqbK7fy3vPcZYWQwOJ8nKUMcIjiGQfNdBkgC2vFJy9RXIE0/8+kvueS7aRR/h0
7KKk+HQ8DYKImLRzeLaUf8DuCeiiIIpaAICVlH8Isyn3ED+oxBz6PfrlhVELTHz9alhFZIK/30fj
jKvWJUxU+w8q2pCSjLjqxOmhhYu7uzhjzMvV4drHpweThAW9ukxHb2H3xSQXizJ0/wnF5FVhNMoc
6rZONKBkHk7VGGSyMULXzwcF4y5cSDaVPttpi10AoQ4L4wJShU0PHW9h877BRuWzLZ0Ad21XGbqB
/TMyVmA1aYRSa5pAepo79ygHGaqIiuS8L3i8lpS82XPxZOMzuY148HWue4Pt8HUgILQrhpnS3D+a
hz7njPVd3Qrlpi8OzK1tlMLKPU7B7QzkKWHc5MQhHUCW36UpUd54WUwKqQKmTm8+yKlo5aD1qkiL
ts7u18ITpRh819Ls8HnIe4/aqoD5GjW1rZK0cBDvPikEAzdQj6oudso3a2KMRRvRTku8pYamp0Cu
st3v1BHveVbq5YnaYRB5s0i9kszZKJmJK2keO5DlsXhvXyOI06WfYZeCRo5mV/+r7zM7/9DqdxUk
VHuJ4G9R+RyAepbHyG7tLruEkicJlQHIOB9F1f0EnjQ7B7oGYiuGes4D/EdOus46RLuMP+0iHas1
UI9vkRpfaFCnyWfXEilRLP7JXr8Py7cvnhz+rwtHNLjIIsXtLEj9hrrHg2v3Hhj0Z62wc9yE8vaV
lkxpcfIXz/v7rZgJDBpm8fLlE3cMM6CY6162eKmANK+226SEcUBQrtbqi3B0Z+SFTBM3ClrNLy6r
nL1DQ/XMV+5Fos7GsANo3yXErnUaHpmVBYBOW8eYCAOp9Q2IkD6FpRZnbBCI47Bjwa9DK5MMIpWc
bX3d49IXQ9jprpyFeWyWGsF3wMQpeuEwr17cdO4Gwyo142TP6ftphDdQIKzsMPkj+FSlPJDKzxBO
vpERF0RPoP2Py5OEnKZMBBoca3Ax7z/eM4i4w80cDuFGtaYJXm4z6XRaN00hbz041x2NRP/DXcxw
liMu+K1Odz30d/j575PSnwgfX3LAIQwmzmTu9LiiKy+cYIG2zSSXKG1zTdQcal9gzbq8msF4tfef
tLWvqXD8p3lkvcsv/Th64iT+0MSnzkytuRe1ZZbY6WbEhkbqvChPN9G8Dgh26AS0EfQLetGTi3iB
53g95zvL6Nplhcs68x6UlnpHdnrKsYfO+VhurH7epYuhKZp97/3kENxEyH0E0RYhSbMjru/2pVvR
L24OSqXgpBpL7KOLkvS3m3nCZ4qVvZzSFkyGOToHrmS2QAnvgKEPvOWuP0CVJ7cMABMIJhQZhz3w
r8DlNQtsmRR2iGAXzme9/cr+Dt9WcJ1U1ghvhKaxlLdTzSrAiQRi+m5wxlbB4Jxz5q0ZDQOR5DkW
guAdwqY/OPsW2RF00JRIVbgzaFI/5+OPQpic1PsBNz6bj8S1stHLBk4S3JSjD/Lrs848TEGizIwi
LicsSL5MG5axxU/dqZ1deDNcf/SEdntrBsO7nE64beCV5pX+pAn3j6HKTeZE/wlIn6FETVUtTMsi
jsVluwW1F/Eyqei7gN/JDnXVQbQBglHvACae2qv3zzIJgNS4ZXdsujzUwuzCiW+OWkrFuQWS17VU
B7ybwUpb8Qzb08NJbbVxb0+IP9aBUB1J9LuizPqIHzpsofKi522dREPv88vrZDTm8muSe3xJ8GIg
CCU19fw6zHJcQleI/CmadExE7qFmtEAckL70udyXvIS4TkGGBpVU08fCURHRHQZvPiGusdSZEGIG
9VNUnvpSbV3G5bDznTXgaUmdHrnMp1Ru5E3vnegOQBD3I+e1fApQpxHHyGN7jTivrtHjXnkAirM2
nlbcQdjw9gT5zzC1sty4TIWf8A1aor24+49snUbIH+AeOmLXJSNhjWptSn5GNKRAtiX+essu8TDP
kcmrfOh03AZMbRV1skMuHjQMT3uccte8OiAW2gJHvLxcvmoUT3Jy3DbeCSSZh9fjUMT9GoWbW0DX
ayZfOof4AZZoZNlhAYqx+bJn65eR7kBGgGd572lueQsQLd9ms6fZZGnurKXEkJmT8x+KPJTjV4Qf
YRHi4ZrsGm8xBz2eYUuouVO0Ws8hIV56ZDx1++eblGDBR0HubOr5kHaYUGW8o8KfX/LPWkIF2vZ9
wbAuzpWx6CS0qFY+VeUOt1ifJ3kDVXVlkoE0OZteZ0K9dy8pppftGSzDPTUEpFKlEkt3821FN4J6
eg2TMf/AZG6SfsFoXq2A89jktKPOextX/KNBmJE0gzzlOZ1TOTVYnKa72hCt4n9ijaAniyOMOP8t
JZZ6Q0iduqjFWYgOWLlvm4EAQYk3jZIWlhdOwkNW2sbp56aq6f2s5dX5AmpoGTp4rXs6eNIMITrG
YARYzJJFrgq8kkIoffbxoJQiELc6pUiTZXBsPQeBcU4X6i7W3mB0mLRHs9C6PmwookAi0p3Colo5
MwhlsuE9f3y9j25wVkfusWds2LVN1I7shaNS2hXQRSytivdLh1X7xpTkf3LBeg+tTIUeM5iFffTI
oepDiM5JgCgeI8lsLlii7MILcaluRLBTMQg90HlNGkacCcmk86BQsGElTZGkS6c7pnoA7B49knvX
KloRjF9uACmdNhJH+pFD6dM4qaKw1H2poGllWiyU38QJoU9KsV2JUxJmNw1TUcQ6PChQRVao9f0q
aZ173+IHLenGBjDW/Q==
`pragma protect end_protected
