// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qfQ9OysUGy64nlmzRM3U2v3z5e+s07tX8WUWoPzQRs1np+VupdjO8iTyI1q8/TLR
eZ9enDyvE1yNdFwWW6M5mmrHf5FEOSbN+v3KqF254HfMdNAtPFTnmDsXMGCtbnpo
6M52nWNKZs2A2tj3V8/e+GAgwJDDkN1CSe7Wr7yO2is=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20880)
JEKGvErr9MfIZhIYZmlIMpRqvVZ5JzfsueiTom/SwecubEul0KF0QgLDFl402QF3
HBqiAVsiPXZkybI9lwwRr6LDccVlAFB7OpLc3SPjewZGQjzF0hFdXqYJt/1zf5a3
jrRC/SK282iTx8Ks3JN+2LMbvcdieeghBpcjc3KIg2wYsT7m0tWrJOtGQFejaJxn
3ZmDZJr1w9nIlyo2NKGkBRa0B7SoE0zBQvKzhPH8sLrFI884yDsFV+tjLgWK0D4c
QSSP/EBGHLUYbH0gY2PZwfQ9/jQLCFKsBh0FneC7JKNLM2OdGudKr28vg+EIGj5V
3LjbPifjcfORRTDxLPuUH3t8MCaEph9XYmrupRj3qkBsIlW8+QielV5SFwX5Kfg1
GxEQQjP4hFY3z1z7RXWyuo4QaPsGmtGY1HjEsNTR4YkZjT2HSEIMmJgrkemqKl90
Cx8ZerlKS+301cDDxoz4DQr5fMjcud9x4szgPmfmH93nFpobn7i9h21MmHYq/4x5
Yday3cVMrBaeyaMVeRiwpZoTCnDBIZzYjmmGpQZe4/mJSli3zAGVnfTLmpm8taBD
JOgy0M8U1rvYLwoKYQNIoBfZR1GW1VhqSc6cPZcLtNy5+szs3qyp23eYK3m9Vcyp
xTgmeaiy6qxmBQPMJnZkV73lVleKMQUaUcHg2OaFpdydNX4+lbaUEKDNuwNa5HOd
pe5exM8vxygcAVDMGloYl7OViBIJIYbbaAhWBuYSYMzoZyuFt46bVnOV/fL6p9zN
Ir/1aFfSLAUiJ+rd/pe6+8NAHqTfOhJrUhhZ5VoBLkccB4COL3NptrD8ktidpFbv
XxaEtyg1AanDkLTJYKPH4ej2n93zaA+Ncc1kZK0yD7DJLkABI26Wtgw6MSUxO4oB
a4siy1m4qccehSV39r2xWQ86SWc7WNOARDqKeTeK1Bt/f84lQ8No/KQ6nml3t/DX
e5Jicu+vdr83p6X/s9UL2PSGcBbewXe3VXm+pzcJtmcYzbymNcSynL/Hul0dwMi7
8sK5ijZwLN1fZbQ/QqNb+f9FkSr37eti7N+pcwFU1CWgMlHzFIi2BfKmJjdPNALa
Tixc71ibtveqWI2+TKpwrV1Yn3blnOmDGoCKAOvRJ6/q0W0K70WkWVg1QjPZZpib
bCRmOUCf6wInPJXhaggBKMZLfv9pxFUoPurEFsgwT7KxNNJ/gPmKHxS0/Uw7/yX1
iO3RzKFnlBNTO7NDyLkr2xuEAEE30K5elOLV25EXOTnwLQcVt+mFvvewaUEw1+e2
K7QZgAmKvz5DCBnvM2Bn3s3E5oIk7jqvLyqGkj+5QnAciWACECWKgfyrbEgbftW7
pH04mcJzgVIUsPBI3WceswvH5oO3HQpnJIrsDyxXekqNz3lcCFUUxjjW/WVEJzH/
iKRX20oC7AccNmdTT7n+GeEiB2LtxtHBaLx5S2o6Hr9XepZMfeQ7UGDrHNioTIp2
k/JfQUn2LlhH8aNEFlqp1VAlzU9INpH1qLh84/ZsECxwWIEIz+fErf9X2OZ97Ktt
GULl1Ey1iPQGM7GhTWZD4Zbv3oDdncxkgkJ+b2vGcqBVdkQv4mXDwJdCtTz11Xfw
rEKdaFSBPfosytgWjKNEDvWqjZ6lhIYg4akEj5lZjyBaTPp93Amz1rCkJKivMXUe
wCGDw6RsizkEtKVMfcYABpXRskCPOwxytYePrevc80/HQMrJISiwVyq2kut/ErpQ
qfwqzfrVbsY5Ar4afOx0Q85PGIuh3IlBWvcmXyPp7ZhNOMwffu4w+bMI6UFDdOUq
KHgXr/OdmtJSIumrELrpDk82MovN4UfADwf3g83xeBnUbG9HUXyP/AgUtpEeDZgD
BgTbq2EzJnddo9ScVy/H7sYo06keJRp9w1QH7iOjtPeFfql4g52Ep37zEFiG6g0m
lnqIvN6n37gzP1mC2knC7EKTvfEU7Yj+ifcCmOzw//ZeK15U6eJPL4nsvyAhE+p8
VG/aOrqNP4yiiW4CSGrlJcgilCEXxu323u3Pkpn5RBDoEZe1ni8iKYCRtXTRHveF
01rQqeuREOpAC/j7fK12/kdAtFyuKraWMm9MJDfXktzlNsTg55U+a6mUr+PXm2kN
KI3YfR8c2aXtQe7uZqXk5oAfDwO4lYs7ZsUy2mQjdRvhAtIGLDciijsQeVjBGmx1
IvivhIZkmz2U526P0Vgi4cqWbqbg9vne5cMwM3CpD5nC1D4tu+DRE1qgjI15blIN
nZgWWzZsYHjAdNvUjIrnYhN3T66vALujkKZh13+wAlf8dT7g+GNK64LmyvSe/EyA
028Qo8pu0PSbBRHFfhNOVuF4/E2nmaYx3lTPWY28Xye8oQMOjDbA0ERQaEHfkGtQ
we5VtQo4f1dvO10GyWeO4pDLH6TpBkiKb+bH0v5SzZp7TRD5g6v5uPBcN7Z4FCxe
qO1HFz5KIZqZ/2wYLBqI/q++3OljFPbxcRgGK/xwCpxAA1Omb9py9Q+PxHvUZtfM
1YPBkeRYuQs4DcMSuZfEEu+TS+Fx3dYgTmGF19r4M92nzyUvqHIustkFjU02ajQB
6BQhMYqn7SRuqpLbObRpCTxO6oCv9ee6yOZFZ8DKgEuVwRY3L6bJJSofK3rsRnVU
HBZ/7/AErApnkd8BcXSHhaTDIUprTwrbdi1xDt7EZb63Jkl2c+umGM8uBvsUqO/l
wQlUWcLw4i/d8SHmVQhjn4by3Pou1Xfo3yAhN8HrmOeBYJR3MrXDd6NOrO2GDiTr
oQmGm0xho6n1J7Xl2WfhHT2G3NzhNi6pppsiwH6/W+8RuF7Cl0XQn79yNGjQeLMy
RzdXWBehRPXLBBXZh3HrLg53mzoWJmu/sNXzD8jZ+YRSti4Q0R6IUlhktbsL6E89
1KnxWjkX+/CDPRoiH7guQAdNM8lCq35ilfD7GXF10H77XumSzLQdBc+QUaQCPQ0R
zOVXmQVNHyEQlHiaIclYK/BbGkB3IN+5cagZy1upX4ke0jA5rabQfNFJq9cOkK/9
Xw4cQ2KHcghhcD5xmyzbO6jNWUGO7i5sJDF7RTuU0F7kJz/bqMo76QtDb32D2FEi
vSRnqxn1Nos+QUC4HZcQ/eM+odKyFMzOX0qOy/k2Dx1agwrVlaIjtJZlbYEQtKXr
QtexRvZn/dj0jjW+aPk0KDsSx+8TDA26nZkVZ1+y2TcMZ8PmI4umRuH8z+qA/SUN
ECNbJYbUf4p81Ln6VpzbLUDlejVKck4fNmfkbJi0dHOw5CIXTSwN3Tm276Gd/Mk3
AtX4Tw6ENxzottU5r0Crus5GOLfpgsiK2+u0G73HPnEETTRQcvcEIL7ir25KUwmE
+bGBMFzAatx9z97LnAxVzcx6ojSx3zWEmPFM0ApxrMIp9sUtOBelSUbhKEgF9uOP
ynSlnFXxteTDd72PY5sPKhzFuLZpQDDPPT6UjQcs2cpreV3PORD5nC/NUEO9Gkh5
iauIB8s6T5OZvfE5+Gd1fAF/4mMzrnxhR0+3eMiVdUk5AdAa1EFnlcPuNII9PFoX
9E46tV5DHgWmmZ9XORmJJUFUY/WNvZkM65lDdMDEUOWhv/dhOJa9JtgbvlcPpr3k
BGlAP7WCR30dqYotmEtaJqjNcGlpxvC6Ethe5pBdZ/XTESCwrdbzbHhUcH6tRRXJ
6Bf6BhwuTU5hU4z9f2w9qX8dM/5q4/AuZ9Lf+g4IkvzBIXaEQyTQq4ajg6Evds5V
9iLYMxzkZSA7UWIfjAsl2iRRmZ1s9HmOHLYU5rzWLxN2Yo8NjmEaQzk/yyUbE2WS
1nE3rGp3yYKWmxkEVmTzO3Bclcsb99YEyRF0TkSX8aUkR0An0BZShkummnd8LqJC
Z7OJbotfEIqYhXmKrjuz3s6eOkI6Xs3E83vBBoMZv6HY8j4huSHenKCYoyA2xS7a
68kcBttPgvebMNglyN0KNnpWXzt/RQQxGGPA6hPUEemMfBzOWTISgwtRpJlctqou
cDr7k7hjio9KnD1FFk87ZEj2LX8J3ujQGoFdsCw1ejxgpjQrKgPMO4byBDdwCmRh
L00EsIXCg243BJrs5/MVvbMWIf6/Btaof7q+TXszjRlDTtGOMG6NeVq0Y8zspS9o
NzcX5vaI/OMd7ylSFi3+Dqbe/O4JfHQeS40ZoKummOEzn1oB0dAC1f3pFKeEqm+k
ZsSOVs/cfrrMIv+/goODaEdmYfNtyKJIVP/K3gS23bvR//Q4DQn6AQXWQX73lRik
AiI+W6uopbOQRaMHRkkiZ/IU577DNa2Fxef0Oc/Gtu2WzvSCB5MVukXcZNO756aQ
D3J9Jq500Tk6obNd9rwFz5DCqOZA7ctRWD7qTzkS7O3Ad7zzXi1TrnD4ImiMorGf
gYI+oDEV00aDSWpDXqzOItIX69rq71y3t6l+/O0gWqvFKIApu86VGFixWgL2xWbT
QXOekWgw87VkFhirYxn9dml4juvIRY0cF43EJC2o1tQ19vOcCIH4h85tsdK0nNlL
QjHtN2v2cLKXztJIIRTl3g9OC2dO6Njyl0dceAKkwDHHyvtpyu9kAgHpxODWrk9E
ebXcoEfA9mYOCG+ia0KRYNitWdI8r7mVzHV4TcJ+VWEn20eYlzD2TbN3QFm7AxxA
kUTda4+NQ4ZuWQw22NuO+bcztTpIc3dZBojoKo7RyiwcYPPPw9gsn1cHGaiSq8Zr
4+2LsKdAvFThEQeMCikMrkT+aIo7ibXPWT+6HQpkLwSBleU/4pa7WInLjM97294o
94NU9u7t16hRnwj9G2B+9IVu6qe/+jVTKpt9kEOAqwtzT/B5OnnoEuXtcM7dKLbv
LMmK00wajDP5xV16u19tJQXqAKZYTHc5yUKABWujiDC0+zg09WBxLPuxRkif35bs
ZA78ncYCNP7OGixK/9Smck6csZJq2S6PvTZ1qQI78ga+UTYkD0FgfD8bELCj2jgC
7RLOzZMLrbxHaucPUHxWINsiolPfoiIM9lEu+pfyvr/ItQBBBqY81hCgLvDXzi//
TVhKB8qDA8lql5ua3kCEO8Ck6LU5cJ0zSnGizydIS6cuziAsutr7B27nUTVNahzD
RH6yjuVLcBsV9tvi8Ur+iuV7w8Y3Pv7Nxt7CIhh1E8eI7zcHoeoQ5cGk3XCfveVm
W2vLZ4mdRuuabn6HriqCdD1m8SIvFbishrWw6y728mZ0GeGwke9NK8aMpE/Biymx
ai5r90IMwXarD2vrnfIJwP+Y1CpbDHvlvQ/wTaGD+/ZXHJMJJOTcjl0Mlo6A18Eb
cPDetwEGRAt3cTv96dS34cLrPrDO0IaMJ0vx2fXs1Hegn+V78pUh3/6C8hn3rwmH
x0YKoSYAJhtyZCZ8Wpgd6bgnwI/N3oTTIDHLvkTTzjem252iQifQKMlrwBnDgSqf
vLrL/v0tBR4ABFqUrfpn4QLvdQXBXmzxWa3sQGw8EwmdSiVcisJr1JQLkz2sgNGw
YqtsrHdz+t2EEx73hfNxm/ygqV19XTUXAmIH4cndEMd0FB9O4g8vamZmZq9QqRtD
qw+7gJNxsvqj3p6BAuKU8jX9D2wI/vSeiKHfUN1115YZcV8Y2ZRQIev5wsxihifu
BckzzcUMINt34xNsa0kDrxNnYFjiLWj4hSsiYR84YL0wd/ng60p6eBNAkQ+VnutD
G6z+V/QikLaoU1+NhTsJmGjtal198f1+nKVniQlfbAaeEVcBe/+t+js/hvaomg+k
Em20s8XSftpQYE4l59hhgp+/+EdFAVeMvbz90a319xx4nmFB+ZKBvjC1pm1cbckU
rBFYOVDIho74wMnzEfMjrWrdB7RI7dCtsgMIfr802ixNWFWOYGhHWR9yktM6CoyA
pfVB7oDRrgWKywE/1ISkKnRm7zmdWpQqxAG+dmrrA1HmLpjYcOAcJJBhg2qMDxcQ
WBtsl9jdEO4t1lHXB9XxwElOmo1o6bjCVnhm84PPTngeDDRjTZv/ma5kCzjUyy+F
qaF+3Vi8uLwEkhdwKS9n/TufMV2QcF2vbjVXKkMsmjuJOBlJQHkzR5ihrjE5pMFt
J3gVoopbCp1HnyqSb5+TC5U1kBjtEHeC+V6opLMb11MVTxzdh8M3VoLT4HFbO4Bl
n2M8aDKAytmZ9rLY3F2z0lOOhPoyPMh7DHJrMiZ+jsCEPDNL9QNICx4o0FODpeVx
Y5r1iEgdy4ZW4G0YJIhnCgE0eq5f+1Hn3TPfG0xMKsCTj6srth+7xeVBWPO2Wm3G
jSVlaRMrjWrybg1n/l5TjVNgFAfedR1Pgc1/M2cZy6M9UtTJXtikDemoohUAYBC+
xOPad/QX9SgB5es7tZdavtle/BixKPrRQFyMatXxcaroUMh9jm0ZfujeourOynle
21cPXXtPFTJqis8MNRai/j4uqJCK+eqmxGJwmtdgh5cCuSfCo9pVy6gnRw+wn+cd
eDXngDnUkhEQ/5Gx8HMJ42kuHuJotUIcR1b02hQweEpR4vk0eep83bkWL+sJJAoV
Ic2GykBCDAwrDNC2ki4L9iDUB/9Gw5J7la9hcBsZXRYsk/gANkV/sQdDReMeF5uj
bkvaoMz4tSayS6/QOYkCCKuMW2Xueci3NABkO4n9r9fUsp5RYHhEjUHpA+YWwvmw
nZIDxxrsvu2vGNC71kAbwVR1EFVI/ANXl09J7KP/sE1th3afM+dsX5HnDLRNhfRl
oOhfEAV3BqomjWb/tIQSmipPPRIQoJFO0H9x2JHn5w7R87NU+ZnjmGYSX6XwDmpL
2MHJ01m3nlvKL1bhHRXfmSmWvVruPaTjuOPB1T3uM2cQuoJTT1RTNL/1IHrp01zC
jHC3CGjH/qsIw9ER0lHpvl2xzYss1++JXSvDeOHyf4N69eu+UBUzLO7CCSXwEcv/
6eNmkXFxe2mUW3eprSfAfgm7gAAG2SrHrbuyOpn6qBNtK30KvoE1gndsybZxRhJM
GHsREXuJachMtyCP+x+Efzdvqnkb8CTf3vR0A5hFAIcRZa2Z/ca6lfqcwAFhBiEd
XUfjkU0+uYneAEWWk/Ibfyec8Ef6SycKqE9Q4uop3j7nItUobZRiU9cct9ooygSj
oUcGL7P4FO29fCGJKxxaOImOoc3OpynLv0RvRlW5icf59L5KXnXtlOQgfAKetEeB
LVXIN8C4pYVlZySluIQ15oFqAM42FwHZcmJuR5iBtzBoD0YevTbcpfSC96SUkAJE
LdFXTPJ04hoofYjWMxwSKn4GUCPrUMVG6HgRveyNERkcsVjkic0BCekqwK1Y/116
xh7dPednlzlTXlFGrWZ1fZiJIMNtYCuUIZ6aRiK9IoS/JqUnLNDedxPQgBnL0uCV
96YGgcqQKrNWNw6N0YD+kix8SKQV5MNdTut2S3FU6s1IzAwdISg09H+3JachS2NT
n0VPLvnfLTGoHOM9zE9XA1GCRURc+g3KfniBLyzGxV7Y98vzUayMdrzJOzu8X1uk
LE59gBULz1Q5neewpabr40TOoWCw3SYMRAyCU2N/ymyMGTr3eiPXmMINwDBm7frP
uKOuxS8yPCkInQNfH4NtFBFWrBwJEfDW0ipxP46Ooml7Lh+R2y4jyUUfTwgqdKbR
yAUvlwMvuQtt1riZbsigAfy3328xMP2xRvDeKhkGP1Tt4x9SoI9IejDcIJ07nhXS
1sfi8+c7UMMLs7+aI/vNKqIbYJymD2KI8bPh4h+j6bbUGDifXwEB9MxlAW0nTTjq
N7zi9pWK51Xg0ZdoNBIxbDHyOIDekOih25sPstkKYMgUpGgrvNqk/dZmemrpcZvR
DDRRDc9j82WuL5Jmp7HnTeILdb31RsK/tHnyKq99HzlZFc11BgO04Jyqm/Fy35eZ
j3moWMZPCkgBr+eRj8WAmWelaRKjLGWlwJAZVbopOIZLomhwvKbtFDqGohqAW38I
Uf7Wx9ZRJCkNTP0afZdwFQaA0CUksLX4k1gq0aJG0sYvU00EI9V4wrfqz/W3sT5j
iBvrmMU5LiviYTAyK0bT9xeeeZ+TvE9jrMMkTYemy7rkgXjGFqVeanv0yKu4XUIV
H5eridUXfLKLTk8ndNfz3aiQzDgomsdoLgg+8fgz8cNLWJQ+/JuNDM822JZfHKHq
vCM39eqlbLcbmzee9f08Tk23nKi7kCcwxt49OPSq/iI+hO3LMnQ5JTtvcgv8137v
znd3ST6DMLZYqx1i1DH2ITQfJtXzIZ1nlr+W3tSB/95tFHCHiLKNw4mrxZ7+1btr
/ly6ZitEakRLkcbJot8vkSHMuHu1xQrKQNUslLIj+kwy0rJ8hZIfKJQ9ekAL7qrR
rlNhEam1zstTMTsQl3MJeMwtJl0PST0L/rcb7DmaugMvsQtVNAvqEj55D6TkZenW
CTArlrFNmgj2bbNxIPwWSrXetK/QKqCcYpCnsghYI2biPqFo9vR6cV1EoKL1e3Sz
ARUhfuG3Zi3VZx4DsAW3PsAd0gQFo01R9xGgVpb4btGmlI95KOnKjlVnJxE70IM+
7udeBtWoRdQXc6KW/CqXeO9kOtV2gjj2cSz4MdVkEeZdhoUQRu3aco73cpeBEPej
qizVNngEMwQtJRedBV/8wUs/LbsBuolCW9zOxogInGoC6yF5WHMw7AzBRCEiPZJ9
coiyRVJshubUGXmb6MzNKNdqkbrn73li9ChKyJ9X5k10odcqP819MAilxTkyvqXc
P3iQfntCR/KmUXk0vvbF1+E+PEfLKcvzWvUXQAZpKTBDjZLHXFjuGDElQIgfZ9i8
8BotpnIzPMFSNGwWWN7kzK5VrrmKmT6jdMdtXKG+vi/PSREG/Muq+7xo6MQLJmFD
FXoJCPZcYhFR7mqzuWEJ/yxBLHAIX11Dn7UZkaA4Ss+d3IqbMc9evmZdXuiKC9Vb
1q1AfH7OkbIvZBiSHlbFb1zv2pGdEEM22I5PVoX+lU9ThuqCFC1Kv9zBJ3SuTqAB
eyCr3oXzN/oQI5EytJgJFNuHGrs8k+87NP69KFJxw7BXA61X+l5aRERNOmvWODk2
DMFlPxmtPo+UP1dvRG876cfY1Hc5up0RSdC4BVPIJSpBGVvXL2UvB5KLXtEOzw2t
qVJU5V3bmLOSFi9gD3+RlMfK/xBz/HY0yC4QTHI1tBnEjdHsoTbl6IWYqQy6O4v8
k/I5MLgTW/mFO59IjoyMQkfMd+nRgrbyUc7c3lphBtSDX9kvv5+OYshtmX2ASK2F
VkkuCnewBkWAnGlaSPUWfUXhwP22+2XMjYkIcnsIJMQ4EtP+SdcBxllkdx10bSZA
R4257PBVfVbSBGiMUHH+Y9abLzL5fV5Vhlo2HCnp+/wS5YeeMSH7WgjD9wugo4qL
OQka3zb5Hg35ror7AI1CLABOH4KBS7a0QCnq9JWiRl5a1AcC2kserWu3GCgdAkzX
UXHOh0KYAanBwPcmhh2HtAPFuXo3tfHoEFHcc9rIAGOUT7YHLrKQqCwRv6/vFbV+
gNgeorG8mbOFVbqIy187hsgmo6koWpUWKmsRmd8KSSpqHOMYgtL8v/tATOyPOpfp
Yd051dI+o60q5LZlz+Bco5So61SVEIAvGftvGlLYTu7D5mZgJ7l59ukT3Vm+RBHj
M+levamH0zfVvAWRRfYK1T4SIfP6+4P5CvdS8K97knCSByfU0+zBy84+ut4mnBBZ
qm3ccxJ1xIqeL4F56a/LzYP07Y0sJOM0q0I/yqk5U7WI0NuIuC3Xp9eiyZJiFwjK
+CAIx3VJ+4b3yMScdklHIx0CT3YULoViORXPqgFgg4sl+SRCKFzSsLWJ2PO39GKq
FzUdDUH1cSaV65k1tkBUBgVzLLbW+PRN94yMUbiGea6C3yr1qnoRxSAX1pmfKFve
c7I4/u+TXVjxXyJoLaRbj7uO5JdQxbPkEo42Wf3wjjJZiDdZNIvpH2zFMovWMKFd
MH5yHM77/zjTeTH+3tgZD5DxEW4DFLgBTmviFm/lxJYzBs1GbqFQ1ETQAfPDfq+G
GCj47HywD+914LjcsD7tTsy5FNVDk4G5pnanVSgnvIkyNSzmdTTdAq4GFCUUGG2C
55aS8kGvOvHCvvRzRneRbEySRbOACsicy2c3IzAuM2wWjo4469cPVVFJZNxD8K4C
W7lECbJ0c6L6aiDTbPg5oc/mSs6bKpeicW4KhAnbBnI22SSvq+a6gvc/FEgLx/4p
tJ1ELn3XJXBhf11aZ8Lr+MXDg4l9LiM5uxvqD9QYTJ4rA9UGw3EtqsMdR6e2TXEX
7QnxhsKbml0kBXPa9Ryw9Tu+jR8PODnqePCCIksORvbZwBJ1xh2Wdqjk+20AQBz9
0AZLin6LBzvyg/RWa8D/FA/N8iFJcNyswYXAPYYaAHDfUwOIPvdTK/Q3WIUoHlXQ
nmYzh44Keub2fLFd4nHYIAte/AnwROK5RACnFTJb4w8gwb9euH43F62gNboUiseb
RmMxk7vBPWMKNtWnq/ZjY6o1GBwJvfDr0hnKdOXtAM5C7JMBsZ5kb8x3HnuYttyW
aG9Ft0Y+mMpR6FDjynyrWrqkNf1scawkUoOZ9ETmboaGmuBMWHFEQ0dEPhuZYmKl
UP3sfRPA258tJJglU+rbNyVeGbKpLu093fXvS2o3n79eZ3tDSR4AVlcYIccJEJjR
XvZS6osjUkJhBeTDwMF+8lbwTAUivSY6gluA4s7jwq++n32l250fCNl1hGq+uFiU
gdwfQyXIqShuaZ0wdz/eaDHHu+R7GDeihBVXokK4rWpaww2OWO7mhJlAu9Oh4sB4
4RGYZIJXBX69knPVy0hqnJjFScfQbKic9dNWNvNFG6iF199rts7J64J3bhmnKH4M
5TgrA2AEsSqHRZAcXPh6VNOIjaA1sCQIwwBbJkDmrB1H6BQJDgGMqkZIazN75fAi
m/EDHTwb6JEDSfUI81G2VQCwHmO5bIoAGwoEHM3o33K3pJA4CiusCYMlSzJGasl/
PIXHPqOQLcK+UZMsYLH6/4nS1tIzBzapMxRLArWCJKzPZGraG/4UAuMgz30Fh2/o
e1oeilFQsZaIHHO00lN4XvoQlB/DQHCmaUE9nVjNKnq3eZNrtns0UjIkpnjMN0+a
SLF+d4SCPILqvBpC9j0IMi1OF67JeYJse/bF+bw9/GorKMzP7AkIKcTDbuubsbdS
8kEsIw8423huNgrDra+g9Hfr4EirQlGGqu7lHHts3+r753sNE5bCV1zxzVLeKTDn
RJ9ZrCG+ROf1C4fT47TVamm5yXWOI4pLKn3B6NBIi8ZzxqGTYZPuKwhvvt1h+I/d
WrXB4odEUOahKJQNnUfwiXa7tDliykxYVYc02G7dR/RcdjCfR2D7tgab0G8eerRq
cndYuIjym6klAthfK37c0tKJ08GmYC3K3YrRtzwdpoWb32dcYY6Ool2IFooFBa1U
W2j5Be1HKAZpbFZPbJkmrAat3ZpbA2pwxyxdpVbWKUF4LzqImc3E8NoyAIPYedxN
00J1mV4qNIg83BJTjwJMD/3+cBTaF4zce72KVc4+apBXe9hDmrKeIKUm3YGL0hhz
1/82Db4cyQtu5RIqKE60jyPw3mzXfsvhog3Vp142P2mqLUrhDH/sjWELH4/bxX1R
MSpmV7ZCQyRBvzCTFMMVjpwD8BLV5B0c/pqhsk9WW2Wl0Mk0B0HMBxWiFd/MzP/G
X0h2g3G0g331A6b8kSRnTp0LsWyUwkiOt00G5PUdi7gRelXq1vb502VYlpi9jtza
UjqSe9qKPI9hfiMcd0uOlqQUDqvokPU2TUCEsIcKPztSlJXIIqQpKQlrKpOjcloS
DcNU0dCXRPYZK7PiBzqHcEG1lnXER7zNC+MhOF4MUOifQIC5L+SpIqOkAnRInrNh
islOhGrAp+k25xiAclZcj9LUJltjbKmRF314b+QXmKQZ/OmGhSnkOskfBJF+stPy
7WXfSVdk4+BYnetlriA5v16N0M8v3AHwhOemD8D1QTiMbzcyAw84BLI1w9FCzZl6
FfBPejpfEUWiWFAuo1FEJ8FalEfTsrwTHZg1I2PftKQVp3xz5kyANXW/eui85876
XfddYKFyYoWCtqM62FcFSCR5ZD0hi+iGapBu/X4kjJnUDgdo1mlfvLd2YDVXAmsf
haucdK29Irktv7hnDxe5cHjts+KKe/q/7LgpGKkTSuyPtelaMU781PmnXM0cE2iW
BzGFayyXnVDqKtddwv3khunU0pbWOg2KxD1Ffh4OON7FKqFQpltW855PVtEsKpC8
QLc/9R3XeajLGCCMDGlEApfq6gmaqMyPTekW2aQgMqGC22zroRUHuRo0MD50Icfl
XVg7h9UqY9fq3ZKk+wWKXrH1/FXi5y6tE65/JvpPdrkztH7Y8QBLrK0k7UWMiu52
CsXSxsrtG33H9OnUC1zvUwzVk+C5mPh+Q33bcRr6DtlIIAh3uZWnVA5LmDqIcadu
XZIUtNS2ic/RzTjjXYe3f1p+1aRZkcb9EnZSMN99WgY9hqB4ODtY/fVCVJk6Xhb5
Mo6XAJ0repojOgixHy1E054PUhxAb+q4FWxSyiToILR9YzIoo4rrqQvC6KktlLhs
JL0CYYO0bJAN1ENoBI4fAT9gOgsR3zZdLto35N78kcfiY5CRtZGgoJothk90NMIA
8Se9nlGwCNCZgZU9Ro1Li8+WpTa1TVj9KMkaXFja8bDlez+qlOWxGHL8cKND0L9M
UDwRe3fZgLGXB4R8bvmnuzJUV+Q9iI1i0U0XhnEaT6XPCkiOs2w6epx7GpN8C/kl
8/AQe32rmOkB1Ed+1OLvc2sKLXOjLVxe08GZNre6YQxel6Bkq7XeIKfnWJEoTzRR
GW8ttmakTo/Ii+FAq51D1cW+rER78FVgpkfBpjrAjPTlMl7ZHHySGW8liRrq8gyo
2B3BlE4B5gvK8u7R5+Mxq1hUlEr5xpqbPCkxu97LJj1XhRnHRHlJk1ocIU5vNAyO
KUYVJxg97AW8GHLd9v3YdSooaFkumKaV02gt+dkUmYUjtESnBGvPa1Cfsl5PPe9p
HhqYzJfG0vee8JufHMlDU+bXyayC8Pe+PBxPbh5aV//6BuGujnIEhwyv+iw0FO9c
evXPcMfz4v+p9igAcaxd0PM/Fe9jm1Cn995u4DaXvm20bsiUBVudprYXke3vliZY
ji2dyYvbLVnwURexFrVqctuBf2OIJcwlQ9ubo6VhwIITQqe+Ir3yBA31tX10AvBi
WE2Y0Mtdfhbz49bJScjaMLBH3A2Dl9WWR7w11W5NY9GzDgzeeYnkMCRk2X7RHC9V
2JHcAvTRiFeFiKqArXmzXxnSZ7qc4FUCvfugogyecMKR0tmdhfFf/Y/G5Zcfi3O4
jzdm2SNbOtPGSUxMjV8rYJH1GzmKu9sxvmQHu0SV1yh9o5LJioE3Tuizar/sL7UJ
+UwTwwgBY62FdSJ9B7+rvlin/wYhFnC3iyXLDxdZVnCe49WXSy5yTBP5z9mbtqQY
jkHfUBBRCm57IQwr+P5znIC9JYHECYOmdF9yTz3wNsTqnoZiFr4QGG3Gpu/hMzvM
bMnJlwCkXL36ExTi5TeUKsvqOpx2hUeEBL4Rcfo7oZ7k1DshppaPbEgIfVOU+ENk
KyTldMG+1I8A7TS6XSwq2wwYvs8GTVaSpywGKwpMeOx5z/ftFLj3xg/uydrAOqeX
F0GlmgeNigW2s4+Yf3nbddq6iPetm/1DcKgDy9FrmpERcV8AIS5VX41oHjLGWvwt
J7CHSgp9ziyIgCt11FJaOnLb+9CqtNwX97TXnbK6UR2qwRK5uaOoVx5STOYZo83m
ymScERMJ3RrrZG+ytPk33F3LhOpJAn7PROsYLEik1Iieixahs1yOnMRnshzWbAk5
zF2pat5DoIVHHYbCTgMAXUSJm0DFzB7gt9DNPMVvSthtnhpwPZI6i35/0OoqlU1B
zX6DIUfbHpyyS/v+QJcHEtbK+HQf8X+EZQmMSipz9foz5FzeHKVVeEMuUhDT3RWp
xX84thODk+z4hSoN0fsKj1CtojTV/F3UDVtdeSXpIlKRl6SZBjdvYQu6epE2QyYy
lljwFmbHL4pno3fdUM+JRlKyl0wWQ0zScCdOUV8+AzT4ud2cuNQSEBWgcAsGPyrc
4iAMOHTCoVvZI++DclVY4+Gc0a3S4C6Y4+M5/E+irS65c4d6UpUKPzuLm/k/pQxs
9rcUnBmTwXJ0CVfarPte+NOGi0+S/MqqqgY2Dsr2fPytH4SMW3yvsut7ejeZRD5N
GrLYGeEqEpgjvNBgTICQSrYQtuIlNM7R0bhG0STGEK9Bpa8GLUs+lbotkGb1QTOZ
h8Mue30h7quMAO9w17H4gBtLFMViYpJhPvWJMNXwq1Y6pAP2rkEYjbVaE8taBw8W
CnaEvetLZkRDCsxxKdKtcwMXO/x+4PvLdyCYpDH+TNx3Itf7U2y7EpmsRjVqVi9+
8PsmFXWkV4TlihjIKWdxbJne7JfXF51suWa7qoCrf/Al029YbtV7rqLYz1BwdMce
6+rfkhVi2jSKlu4JatYIGXNvmOCJQjPAPd3f9/x4YGFGO8Wo1im3dBA/LHfcxJrF
ejfZhInIlR8GZ3A9T12cn3Vqsm+OV8+cPTNkXkPH+n9hYlWNCPaD/rPV0FpFQBUd
xV0NNWTkC/i3f5BvTBBsEhawtYXKKqfXTiD2v29jBX37vLI8Mf3G3dy/GGZ3d34v
vX++zW2/knwWPO+z+0CuczjcqU82ImUf06IKfDow9FBbYnI+8ZLkgrAD4PJ8oyMG
XjCwV3oEAIoDTZLZr0US+wwHmwzEbPa3fTqlOlhdwUJwIPWgycJT4o45qoAIK5or
2KqCCaPaDavMPQ3tkSDprVQpdreaC9Gx3USTE9fK9OSOnKFUu5UKNLpHt98UYjWu
Az+hHzzL6a75uDiLiGvge4L93hrTkKfz/nzQ4sD7TqmH76/IPi1U6HMxyE4D9nMn
wd8WpZoWn2NRXGpXtxWPybbQTizDY1jLGd+p5usyc6eY5zZY7vQt9itNFU/pPnoz
Np9yxOdmyKrCZ0r5xg9Fvq7OMafZzXLp5ceT4ImWIlJYm0GFafrrZE10OHbPSu1L
5L4pBIQhs9NwgcpEmt1x3F/4gtRPO8GuUNBYMMTFcNFBgS+rzzPWXoTxRZFS+ply
zzxtc95N9RCwuo1tuwGDnqPpQCP0AuxUBXPo6a+dnN4nF+tEUKn9BwaYmWLluXT2
4/1t5XStVd2plEQLhuwt8b+9dmypz0SFbVAA8oxQtfw4PIM6d9FYFSPkhQNb3Ihk
Gkkoir6b2PU3vE4ib0VaXV+n7aDiJijcPnYobU2k9SI+5pjbdX8wDaQqC3rl+qiv
WKQIwf7d+ltk5yzdNy+SzN2HcSVrlDfTv9La1XxSH6X3ahJrRkvuEyGuz5M9pgmE
sZysBVnFhx4xASdqpBZTpfuQARPi9T9fWC1VRGT4fCY0dKyrjJvQkcZeSdBgSDD3
c2o63KgFhvvuZMGqiuUBD+PbXtnT3pWI0JR8X0QkaLSciqdt5kF70UWH66uWxrzP
tSxXTntYC71CzCPOULNI9yrsZ2B39Dcvmo64tCRG1HYwcPr2+Hz2V2a1prZ55vGH
2H5OMOEe3oyGT7EF6EbNeon6tCiFnEsFkVJNTyfsiqVMNaUD5HCH7JUPQQpj3AC7
FUFay/S+1wK+lbTcO6VTa/5G3xDjf13QX0GVJBXMbJkimMkbHgQGnv8LXINmaGvo
0VZip+DiKGH09QaSLV1yLrgbCNyTzXYYVu4yGD0cYtUawkLsqEnrLyB+C7GBTll4
D4+u97yTbNTwJEP6liGxfVSV0P3EvbUD5QSUM5MmAR65h7PtOhf5CJiEfK54Xgzb
8GaL0RKw+MvuZcif4E5RPbHEWf96GSR01srGeEw+MVHzrO7kRzgiaW8NiqdWnbRN
dMuXku3rXOHxgYVAfsCZZrS+XaJlSqZp88UmTomF9V2jYVo2fUf7ItDltL628n40
W34mem+rjpqrzBnw4j39LRRSCrkht32jfvRavFkGcOrwYs8u0aQLpFCHHghmgZog
uuLJC3W1hG12zC1+POWYDVwEBLFU5izlo/JESwxWllTQpCNvxum8Z9KZ4gHTgxSb
WBGkfYVIhUu0Gm+A0jV8cT7WMP1O3ii6qSca/6zWyPTTJj43YbMd+WwsTkYr32Mu
C5a4kjrnacSHHPP3wJth7GjZkMjnS2ljy9mnfTgeIV6wAinQC0/MEixw/hxwX/WO
auppyYwsfWFuIj5b7ZS9U/H+VeL1U41ukddqtG0L0cdH9J2ElZAjhzBO2uFplSUg
hbC1OUBmIIx3VO+2VxTmcXWv8is2wLN683GCxZgA8ZDIaHVrj/F97SDs5ZWNSUOc
MlYxJkuO2BTX3jE6OJJr2G/CI4g1qdlYDIygCwoEBKe2X/cSxuB7osWDafoIVGlU
e6s76R4ATT52EqWGHrGFPD5/94dqt/ygpGoM+WS5g5xRME1TxGTOeQSyKfTk0cKN
uvUrhngABWalyVriXK4a+3yEbbRnYuRt7Y/y9cnpyyyTwF7VQShfCvE92PneqlpR
WxXBgjHt8Vg9XP+VfKErmRy+CsDHJ1X62TuAVuToHwfYm7ItVlo+RO3fdYW4q+qL
rLAcf3s9aavXkHJYYy3sof7J1WzcvmlDbbAtPsQPQ2u1r1C4J5h84rM+EKvGBiL1
WR8UOL1LpfJfZrdBw6pzYcYRZY/XYt8J9ZX5XHgboHly87juGt6nZtoJOp1eAEor
Jal1F/RSedVik7YS7grf6mA5HbCrI+GW2pBbBM5VLscESacnrzyk3eu36tHaeZEX
WcgR4ag18Pw3mKK2fu8XRtrS5T3YGAvgqWV8U5zKN9Q9hxSUv+MWBJiM50bomjGc
EPoaEU+2cpSzVcaO7SvHh/W71TRiTdhr2w7tYqm//msZ6/kvoBSfBmjTsy/r42po
YalGl07ZHz0ChBMPIbr1hjPE1P9iv1ieIMK+eESGhpmaKDDVA+vDitqRY/vyRbeY
/MazIaYsxV+wG7TLwmwmd20xAYrW53qDDND6LvD87TqQsc3t8WSFjf+B0Hx5BfVK
A0PmTICLQltjRVIAVFqH4DvBsXNF6p59CElPK++SQ+87MXBvjRLHMAjKgmyjMzF8
zC1Uj11ym7J0D0s5qojoZHwC9BI5bHr4BwKSmsURPC5XsybGB1Q5mZhmcrWBdTmt
Py71szU4hpR66T2//1AFV/OIgng3jaDxmq8BYGg7yZ4CPRkOeeL4SZ2mDjPTBvWd
7k5pKyfNRg/daZ/VYhGZJHrFjcJvgR/vjtMgrRfm0Iji19+3NwEs5qBbqRFE8FU1
Udv7rO3bMvntd8ETRG4jcRqiqif3/S53DKHGvXZ16WeH01LUYfZwvtRXLOJPpcdv
gjXrz2xT0sMAd3WDWKIr/3cX2KR8iIGBtIH9bDBvFiyTVbbzdw7snK80O8HMlWpW
RoW9hanWk6de1urwxL3bafolC684KWwf0wsX6gkNzPyOeBfOBOdbRgCyKfb+KWPb
ZJ7SiUJE9HxSy9ELcIMYNe8CswyduAhY8YWx8GKxs8s5J95KYw45xxLybwlJtj5w
jCjz/hyiJ2Y36yzHdO0wg3o3URMwubIpr8pk5H3LmDEGdHC2HraQCxlMsCJxh2ta
/nCxVaCExDB/7refF9OrHsGUlKKg6aMnduj5T+sMDA7s3Eik+2+cUTRhwfJo9kt2
NGRM4BwNztgAYhgL2jmfCtxU8rORH5OXoGGAj0qiQoPXbbTxTgnyFG9O5AZpeoMU
8Vktc5wDQWxOhPQjsoYWU+CbIZiudKtW5NPqzzd0cIL++MWzD+XtUA6rTBUkHp/H
lfZvRQSFuzudpBsmqThSedd8VUHrhfxE7O5QuaH/dYY5tTqwXBJgHKhOi6IULWfm
aNSBpofCIiEILtvDxjDPBtvgHeMHJUiWMeXtyArygZoo/cesSeSMROCb7ELdxMmE
GYOYkZevqcteBDlXktkJ6SWpzsPr/XrMGUzuRTa4PlbpCLl2IXrNSLQZlHAoBw1l
6z44ojBBfA/WQ70+jhR5cqmsCo22V4V5Ep1xW6qXb6ZqPCOgD+5dK0OKA4nbzhM3
hVLYsC4u1e3fSaUq0fCQHxYV43fEXt3qNocr4xWL+Be/DFpNoqe00ZrweynYliak
5xFun9JOGzMDW8NjVQEEISqki1P57sChgv1LdWeo70uViHY49rOPaxCqORAUqRcE
hisMzF2p1DUr2WQ1K/j27WiU41Md8qMtG+bsbPoJB0s5FwTMCz88WprefGn4SJfJ
DbcRcpFqA94vUoA4uqQ/E1r1eJsnAFb5QSN8O4Eq3WLVB5Fm9FtzRE3O2C+Tjm5O
Xz+7+w+3/03moCXWbGmeHNFYDe3NHc9qUnhGT8ytgz9wuAJRYyoNdmQN/7auAg+i
MlFGlb/UXMFGZW8LMHGfAbZKeQwn7W9YlfAcKt6GcHZ/VSLRrj2TKz+KXV8eaWXv
Abki039mHHOGktHPqJm+UHbt+zKB1Ebo2exsoJ+vqY+re2bSUz92jE6v3S89QoFy
1b/6EMVngPfFMVr3NaEm4+1AaEaTtWe3cBE1HWcwwBBa3OXkm/hMiryW6UfGFh1s
PeBEinQj/GRacRAvv8p46zFopnSjXTKwPyPYYhTVESm/MO8/PhZ94pfgMGh1J+TQ
tX/Ss29DeuzS9+7Lz/zB3KyJ3yP51N3iIu5fXM2zESKH0q3N2cyu8h/1RqvcyZ2I
WtLKt9gxLjLYeFsHALZG2kasn+ntWGeiNnB92UP6YyacYUOJBkwkVNNWL8akCmQ1
8Ibk4kolNRJg3vaFgThhnZuwI9FF67Sz5uzwgsrsk4qEalIcEEMOz0K4+1iUkfZJ
vdRgJKnNAsLbdnqeuoOx/NKth5l3bnVaMjh8eBHlzy25aGy0AN/ht4U4NSxwCKMf
UT33OUucTHwhNeLKwmuif2M54F2lTBeaaXajtEbDBXNlXofu+7qr3comuTcUMlWV
lsx+tKND+5UhFi7hzVemU4zeaqSXfOTKEsyXyne61nhvS9QbAAfaamfzM4qcwnRv
5rHtva6n/6rr7aN38PJto+Efm4jKVCv+wTrjX3UF6UcPn2Zm2onKDQwGPK3iGDa+
38K0y/fEIfEuHU2CkaAr9b+116EcF9Db9zWJcy/CR7lrzsnlscK5WyK+WJ374OPE
OXLBuuddDybyluAZKiSQ73Sk4BoOYPpvzykIx4kxbHDUIGkUsvPz4W2ri4o+Pawt
eoIzU2nxfPMPTqwVAm30Orofe/4Lzr33ipMZJkaGIiMNdw62iCC8q2hjZ1zY9oAa
5rfm/ZjBIZ01yPlUGjQ3ixhCfrT1QgO3Opu48HKUlhR9eSV8zrxFdzTpHZ684On9
DM6039DjjjHBHj11X5mGpq58gHzhHjo1NZY9Yhtyo4v8s0wF7/R9MkKv2u26wkYT
S4vy2rbp9dHITTjXL8wZ20LDv2wJFa3qZtzC+6EFJ9ROUzfQ5wV4ujElbXUbfx8H
jrED3rLyXvDJL2meeFHo+FciulDl0ieEu+pTFc+nudMnHA3Syp3PxgGyQoMLPk8P
xBnAvBY6HW2xVx0vG2ZghrvrYv64OvYGVCbnK749cH89V0Qeji00SfrtTpRVhKTF
h/T3zLV0eRQR0HqyFVcWNumra2vxTSn2x9Bty7IjjN4oR68rY0MySHbQCinVtBui
EV38yY+S3s5RgAlbdS5XpGlw8xKRXtrHfNjDsO5F3YUJhmXZo9IEbl3FlgACgrwF
AqQ3d/K4dT+nD2CYIxcOqCO0bMFpe4G45Tko0uYltm2QjJaNTcAKqt3wTBaQube/
UfGkAeaMtVrUc2n4WMxIhcm+9pukUGt5ecKPi9eWPa4NlapvePIkPg/ga2v500er
5/XKDs3O2kW5s3hwQYNtTJuvb0DlTraDEVeSwuzIUIvkjaxrrGm+RrbgX8dup5/e
PHb/NlYmCLfiH8ejcSspeXuSAGakvF5ji0YIGk1Ay2Ebyl/nGW95GJ7A5W62mWym
CK3/ND41Y91QhMQp4TwX1FvVXWebUbUUgdeF2uWhSc0WdOaeIRUjaYHaLG24dPg6
r0ybk+70gamSXrLwyzWPjUWqK0sEnn81FrHJZbEfJenVqUsJ+Jq28TElI3exPZp1
wXHgO23s9RIi0xwdvRDH9FwU9T1BEL3uIc8JMvJTJsFukGS2jT8EbCG/DcgAYrVx
VG76y2XuGxsHNXuL+ycPedsD3lUY/OjCikeJ9IDSzGhQBRWqamlDxkJERWzoNe7w
fvzi67GbR4ZHBWNQCkVE8ThDYWR9R7Nl7nxwK0tVB+jlpYFMzfcZn8HxM96nyBdp
dfnZ/JnBb8gr2y7iK+abbbquxk4Szm0m1KV+LEJjbHrfA5i+PpA688H0/kp0a2nn
vYXADWDcqNfay/3zTLyDK6Mvl6qGX74K7KSdvxF840jOewu2DuGCzRMHMEblqQ4a
Zf3vO6/0XyvAUx31g6JZMpaNl5wV4kPx5iGjzkqv/rmBk8J+CqKhvGU+demG3VUU
SeLuoGXRWwztEajH94SHfgqgHUHHsuiaeYz4CFXnIuIEDkRgte3tPiq2cTNck9Lx
4vVBsUXXzbvLLs6W8E5sHC/83P2LL8RX2TD9viGTUS21o81jOAy4VxxL/E0XBb2j
lmW36M+qe9pcMYJgxnW1C7f99wYiNyXZIgx/D85cbj6vQQ4ipDjB/7yPm5YEuiLb
A3LmO6Hv9L8PV30Wwn5WLRr1imeXEP+T76nIaSUbRq7MB5Pcin5q8eKsz6O2I6Xg
+6/y3xgzdkEp2mWaEEKaIIKPU+sytOssGDWdKZ9Dm003dHUi7z5UuXGH59cA1O6/
10VoDft+MvpZVm9njRX1n+xzHtK0amAG7u0AojzXib+Ngc6NGCaEByMmCTfvnDoG
Bk4MXkd7XxEyEIRDnhHVDGzH7vfRzirvOfvduNO0sSp+DEkn8N5Pbe0tgK24TMjI
ij0NEfqX+xrUwyBSnyGLGvwAjTV0LB9sMCptBomIlcA9xHl2BSaheAyEmbp4Jjib
nMbZv88OwWyYaE52mbWB3B2fXUVrCYmN06hwe7OGeIBFV/ojtRoiFW0TjSkpZCSl
JkE8jGxmzADVNrpc/NCY3CD7QO6EZI14r8q/h6CqNNu+rbKTTAYZ2fSrsa7WBGeL
q5UYKgU19sn/MmoMBwuSrlKkBGeqv0sISObj8ug2U4E0X5w54co07S83XCBkNpM/
ARrH2XH7ArUcui/BAWdf22o7HoIAMh40TMkgZPya5lb2COaWBZPxKssRoU10/kSF
RTk2fcWjXxJho/oQv7cHFOblArAGPDn3DYJRha921/8lLGoEDQOHAwz8vALS4RRJ
HWK6gQmf25/fk+w3mH+ef7zEX+60yH9VqnQ1dS/nOR+utF5qvwpWwE5JK69criCo
hsMWHM6aer8gbLqms9rWgadQ+tm0JQIvOvqabeBj2c+9JMYFuWf4STLJgdnhcLJE
PfUFl7OjRmBoePk+dBWiv7C2hT3ZggNzNA7LYkmS6CqfrwmXY3tu5XYwpXlN1sTZ
LxXuDRdW1XjKLhHo9lR47dzUdI3T0tuBvSQDIm6sj5tmx3nskLVaC/SclCjaRr47
0hN3lYagxmV/SsUzqmZmRa4oUbOjTTtDTL/fTGwndQ3Crn0PCwzZDLuGSMHUakK3
AXVoWhYOZbvKQ5gZZ/HMZewNgeMXTOPQBLuQgUILlL8GYEafK/x3wO9bFhNhwTE+
7Ep9o6zUbJoZJ3MSRK5XdEjlKQ6Wwytawmr3Ozb8vvNkwhW5Om+PcZuLMkwQIDSW
V7A3xklWLpRkE6GIt0hE/xf4lhzKJVecxdeGN2HhvB23ELbEY8MMiwzfvqQm9/UQ
MDkOp5hUk+mdqXUnIV7sKG2sVqwGtYmlPWC4XXGs7UgA49cv5hgfin4wBvCe8gXf
lcLr/S+jJZJDaX6Fj0lvjSE6IzTPiiW3BEDBURsh3SYmfgFhSemnhamHCparjF8G
CfFPiDIFOEC36ggS4+kTPiHZo+xtPHefUr+KPI+/c+tJTL+cz259OJWWMP/jfKNv
J1oiLu7q9Net8Xj9XYfDX7HrZj/RORr0qJ0M6eeWkjVBwP0DxCMQlsY8i1BI41Ob
4b2ckSmqmfVZDuJV4/dzHSy1TiQ9PfY1R8j15YnEszYC2PbvtPnYuCn4cmqa1FZ4
VuDp72ffAQH2FU0z70nVATsZBIrcYZr8uTbaa1R9prrrz/nS25ZWJYztuoGT77Nn
jX5lGHOO+ZR55KVOYp8wY8uPMOpXDUi7HOyAcOO4+ODW3axubDJ1Lva9+pRjnNNV
vMMAg/WKW2pOkXpv5jNgmVtEU3HfPp2ltucZf4ZoEyIrolxGBVY4fu67HGh6qE36
fmOj6SCR3bNwDRqUBmRHl7IVFWDU6O9j5KwqEv+LYRd7XDBtH+k75HNhWDZHcJam
H66VuWW0bjqRZ6hEtDEI6GRVt+SMoxToGlxQNuxt7LbOz9AZn7J1NlhztPBlQOIu
S1Kus58wZmLvB3OSApp9jH2IDCPcLgp8CH2ev/0oB4Jw+UHezRUQ7qCqVRlWiyaA
aXt2Dr6bwBMfKweMyGADjOgiREytK5Do8MDha2JtHBxmgAN49QzR6kYrFSqOs+7B
hDQboUkaXuqttk7dCyCH71Lg5RZshrn0kz72Cmc8gzMy6t110Tun9HwnlNKqsTHD
KABAAM1yBO1e0vSW7qqQeljsL18We+jJpIfQCdq4iXrsV6iy3by8wuKwKqzafk3U
I78i0xKwjPss3IrQhUCwqrKNBVJZ0oXrbcVQb9Kdx10JL2F31kS1VLX8QL6ITcc0
Y83gbz/nOXnKREepgkEU2yBf/SLTEuvMyMI2FnnqDv/nmMDJQIgHwReAQIO1uMKH
+H+29gXe+NAujhMqS3FhN8IACW3dL9t5HG5jjVVrzxTp2L2a6U82wyMJA0peFeUB
JNnHzyEyYAICM2LSlGGddb+UaJd8FT/ggjjjXwpvRr3oKbyad9H51fkX4VnVa5rv
QnExjxrrT0rTM0OdFBPpaYlvu53SFd+UY723Xvnlv/BYRIghS8A5oK4CcFtEHCFq
mRY7dyHQB3WC9R0jPQ/nZOaEEbCOYlifJg7E5Q2tdNA3lPu65Um41/8SJCD38CBC
loKSPd/X4ItbqM6WAVictxcaXMuNy9+hhaUGvO0aTDubYf+EivgyEBSHuVmtxO3T
nwLLYSgnN4729AkI5tt7vtVixT15z5G8CbFChOTIJPVE4kEbl2HraKdvkJ10WNjK
x1XgUQm1g7pkBWzPPMJjIij8lmxEEvKuP6WyACKpbeIOusVmCXTQAbFx7xcudR4z
oluWtrtzK967/9GxA63B5WvRv/gtd8BGNriVcijScWNkOdjrwLJU6jXzehM+VDKD
hsfNhJ5HtuLnkjdx7Sc3pKcskne330iJxATAH0fMgQ3bTRJTR0tl6r+sHUp+vC6o
PsEeFrTVSMqzoUlvqb/kxQWbhkUtrNwQExerTDyr95scvyyt2f+KRhbW/enDBbhW
boE1MKNVjFGi+lAYFd9oHDGFResKcrmi9KqYCz1q9F9gNprZjVvCV4KmReLLUYrC
4S1Z2M0TV2Um+zHAiDfr7oYQ+kQjangDiGgKlibMCxWIlLUSSLXG6rxm6tbeSxUS
BwwyVIvGL+TSvm7A3deYtje5x9BbjboZ0DKqWgJfjcpCMie7fdWUYOUkyZNIqol4
aj/x92Y5Z9tPvLLibtdIsQLUYosFQ3+yovZzHPaaVxPpVNQUdH6uwIxEt/OLMVrn
BRYeZ4qCeU+kgnu0jlUq4DJtAXqTSnK8jAvYZwUph1kMKI644QRBVwpZihvjqrqC
WzMHjEgmQFmYWR/EaRNAwQoguy53574y+yydMB6dNllojsCc5II/npTK42qnzfVF
lkz79hrDoxCCE6Qd9ciR/m2/uys9tukDZFfKhaPA2ufFaoOKdd1+vTzl85UQzY5m
9dSUReRWcrIB13kdBtvN5lSrZQrDZTlvutJDDqcxtikbAXdCljumJF4ogbbX+mSU
p9ApbgJIesaPabI3cLVqlbgYkol8kdkVtg96Iott9xtToH4RVu+7w7zuL4eQQo/d
9MO++vvOLSBjKTDWqahQmjzV3scfkU7NKhB+Sbb92CilupSrFPgP+zzX1TFShJ2f
TsIy2lq9gokt1vQEvpSp4px393D+btA3NakudcV7qZKQlV2Z01xkJGTrjPUZGNGd
b5JOqN88kGR+/cyLJWObmhPnR0E0hjUmtJIsJIC038+Zs4bWxVIcDEi+iU3ZPUNx
unuvRmkjVOw9UfbC8KU1XLbwghBLGevKklmue/WQ6WM9neO0xojJ7bISl2IIT0hc
Yt5Q86G8dHnWZDrZOdll9bAQXbwRD3aL1ZefC6lYKynj6omHwCCZEfHfXH2Ha2nl
OWDpxKV5XMEjZwr8lPdZG1LQvsThnRSFSR1XjMsbWqkjCZ7OEiAk4yq38dhC+BgD
ALZkyZrMxtd9TomADjLjyVMwuuCDmQhilI5thIc27ZZsTH4s267uVTkPUyMXV0eV
3QL5/JZfoxoE6CCTRg4D6H9y6ybdRgL5+1S2DLedACB0EHR9fGqQujXwCbNG/5x9
N6ouhJvSb22QsqMmGQuaGUKFrHWp2SHgKRLJMFlFNi7jzSnCYV8/55wn2KKgwzQH
9Kl0XVQ8c2Q5nK8BKBahgDTwQTzEsV7xsbDXMDE8zWElrjCz4eD32w9zNpg+C+gy
e8/gQ3W7NhhWy6NbTRBVK1DkfsiHd2vqoSrLyPBxUUuG+F4euZIjFZR6SYDjnCXc
s5dwmQ1MHPRZiDL+9lXTUuhABmvsq01QpBsYPG0L0JdgIaN0caMxtS1EhSpZwhEO
6mi2uvyCP99UmRAlHO4ECoXSqahBPuTYkb0MqOI5h70FAr5bhlZSbGEBhG2fpfUE
5yUNIWPI5s0n5o90b3wc9XIbuDhmo4dao227L+TKw5NHWWM6MHV7cto0BI/rq9FU
i6oCyuSAFLAauKtSMSNdrMAiu2/QS+mvw/u7b/6jTwAoTh/GpXqMqhDFrKxeNS2W
wGGbIbTPG/pqpwNQIIsI8FgyLJzdp9M8NrMUVty53rfpeB1hfw0L/YQld5sIKW4E
IyS/ZEKhX1SxyUEnm87KhEYwb6tW9vD572MiSTz+MeT66bmGGk/wb+iDxZMWoO1j
g82lQy9y4w3zWCFUHWQzS6cT/7VhA/SwzoGZCfosmH36UifallKyTzP3tQB1IP+1
jTqhcu1dw/03Q5h4x3xtqN2ELKmNaMaXZLmTdHnYf/vPL0UwR3qu4XdlVprGULVU
oP2kUeyI8oQ0to89VfT09NZhKsx8SHlHjAkl1tYHIYAPUuWm/S0ROkzMV11paXJ8
6IwrCc911kIPr4pHl7TniaFoo01fZoaJqF8x+hPq33OgqdhoQwGAUKrMob1tWkrP
rXEwcqLxfQ8kEnp75/05YnTJKXyLZClQzQimSlSFhkJoJhL2J7Ttvj1T1LD4FD0F
64AJWNLBth9yCZcm7o5+79qQP060xyDdeoE+70D6XB5trXf+++NBtuDfQZY87dvl
qsYZ8wv1QvsS1mP254rhAo36YgPxLWW8CNiDpgeYJhaWWWzLVGeGz7ZagJqgjMb3
rPExB9OBcdY6Rii6gPz8olt2zpEzl81cB3Lg+BEjriPjG+Gl8Kya+4ji/mPe+tLw
w6Uu1d0N4mDehWhfjyGHZXuufBHDpcvaaiFHbJv4Ar38oXgz4vSGh4r9IBF+NgaI
UZrBREQ8zbkZ+3jgWBDck/MUx1pVQeg21LWV0OS3ZAa/zzQH23MihxV825xJfBly
dRmbjGQ4PdGxKOf+bXiv963k7kpBHs/NQq/LACjNVvWAQ7sxd32TNmJemyVxOyNJ
3M7GqWRBpGjBoQoUZw44TkiVyxUl2q5259RXyHczKluzsydw290GavA5fbe+P8lg
Sxz1trs4HShT8kTDpx40gAPiaSd9yire9UnRTlI4kNS59sYXyd+NThXFfQ5hTJ1Y
h4wD+bpaIIeIaO0r6LyZJ+xdcq4HVEhoi86K1ZB8oAKkqxokbm+tbOHcVyT0Eo/b
bO2rsDpXe32dleMiHzPtAMhdeQgW9DiaInXeLRosojWwim8YOuYYoKr6D0Kq9x1X
PCNThWEVbcXn+0qvXskRZ9U08Emf2uncfmPfNaEg7S/vLq6UMQLVTORH9e9fxDhD
S9trefot+SRzMkNYjf5Ah0V3Jzx3dY4QPZC4lqZQv79sT17rY+vaKR/qlAs95W3p
t8o3zDlHkkwDrE7Ek6+QQSBY2Jzq6+4K8vhSrwGaDxiPL2/MXHTh2f4ulVbD00ZN
BQFJrfSK28G93etmjccHgCO7SeG1G7A56PN81JC0/IOjHHpp5l4ZtaE4v+vgv5Cl
RZ6r7fx3CYiv7Mud/pV9SSEEgyBXoUyxtdTvRA/vzWctKKA7XJoiN96eKINsRQjl
GRgsPpYhvKWpPMQudSwMKqkgpi89aZaAO2h1OGkuWYIYKjqS/zCBh0U9redSfBQJ
koGiOdRobxLaEoZBV3ACygyUcLu9BOEZbOrdd1H48ueghn97MY+rV4UIe6jTAk9z
jWv5BagoSnVonNNrv9qxY2nxKOCgpu6lYal7TONSXJiChBpH6LGmcyvAxpFmUSyl
4nFDV+c0C6tdTuBpanOYqgJI/sGVI6/+D0Lyz9NW68BkrMj1KW/61U6nf9+pAYbJ
yjKL30GlCUOrzmog4CjHrpNpgB7yrxHJOx82Y+DXlkbrQuyUFiTc6vE7ZKbvLrgB
+LtZQuRA1ao2L70IEfKZ4n7UoZ5OzLrc1Acvo1/G+t5SuBav/P2eXn8hvVvb+ldo
IoFMhORoyHHpaiYtCJwAB7TPlpMJM2TUg3a07z7XyYaoRg+BLTu53iAWqOWOI+He
UInuQZELXDgPZPCn4D04JrxVQpi4Fp6Q5DZQiDNrC1kne753UHm5BdoQEElcUm8d
ZIkPpbzQ3qAbZtF6gBSwsV99nAJnm5iBxIQz9rN3zpjG3GNCicN5nr120/E4sC8/
bka0TY7JTgoTG0GTRlBw5+xWUdodta+XELgyRyceooC3sxRnFyCVX/HHgXfsUGDy
GasumT4AiF4n7DQr2xDnNbf7ECmJvzyzai8cFTF7NWTgO1nuS+A1TN7E/ndDWFfG
wXZPjj8chHgIMn9pQoI00J4d6xxsxnaAtWP/2dHMZAKRGpIilKuJbMn/3aYulf/k
t0U5wFfs1FTkJGbr9+omTInUFrdEI5Q/UbrvscdmzqXSgh0gEWpBVmAWI4iFG1xF
elcvDvp/QcAhAow+G8Gb7j9v1l4uUvgmUqYzJda0IjNVSwG8jSywEreANTruDP+g
FSIb0FxOss3PLc2qS/q3aQ6pklrLSTK+y+N7dVVPAAqCHk3PvxwDtcihC1xH3vmO
UwVBhU/VIKP/AaR+x8Juh+AsWvcVnpIXu7Aq5bDQK3/Qbm+MR29/row3oXFdFKq0
X+fvEoNEkU2veu9DTBZMM/8fHwlwNiXgUuADZ7Awnm3APTJcHOSwmFuUI+IT1UNv
IMu5t6UJbOEqVMSHQHj4YBcPvvVQnm4DjljCJQOmqZAYKx5bKp8NooDR5zVkiODJ
WPbkw0FAp1LRU5VvdIbG3+JFz1I7TMUUgCT3+O3PJzfj9o7peaO2euJKmSsnVJdR
GByWVY4WiEkzYrTTymh+JD/qN2Q+s3Sjh9xNf9Q67wQF35MM9rL2HKHksPmyGLIA
8O5wVwBeyn82vRUEmRK9dXSb/CPFEYdzQBlnv8G5Khk/HXgh5QHZgLlA0DAXAIoH
FYcj/YbYsywqOgnq0GqruOwcjVaaOY9wLoOQHcxXwB1v9RN2MBrmUWH5tti1uYZj
2m26zDct0aeakTfejgC4bkH2sHjsm18xNfd60w4S83X3F8u0q+fv5gteIbS2nIzO
`pragma protect end_protected
