// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AXG13nBm9rUeeosjtBx5rEsxnTT7mypGdM1DrNO4q1odCGYtFlnYeKZ8J7C3OLRI
Al84NV7tG56NWSPcA9DraNCcniOTeAaNHX68BatnT4LpGioYIXyQACa3DFlSXxmi
Rr4cV3X+S8w1gcrTFxsGHol2oThkG0Y33ZRp5vh/qgM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63824)
0+03WGlaFpC4vb3G7rgqpqAz4Gz5rQMg9p4PArE9WaWeS5p85nn/3+HHi3qRw0fM
uTStCocrph2tnpIhuTZ56GTD0tGyqu3QmcPXCT60nx+6E0ckUtieQ5jgGHlAAzO3
UAxW8MO8ky1cRpknXNrbVPNJ3o+SLam1zaRVXR8RHTHhV0tyCp/iX/hq+AWkG5uM
1eTjIsNWi0v79KTHlyI/hhfCLRf7xSci+7y2M8LGKqttUUyrl6AS/OC+tj/V0N6h
X953trQPcfy/ISRg1a2sN2jigQdg0LqdD8zGUwn4/sVclj7PNaw9m9pqDouU5hj9
pjamsMXNWt++OvHusGgLXPNvfqeB/Hm3vZUfAAznX2yU0V9Mt9zVnvDAsHPbKPPx
08Ed4KJ6ANmlzX+nG6ha6qpn1SsexoipP3h/eM+hzUXLtOmfbpz9SW9vyfh8p4uX
Y983AMxy646Yjep4yU8YSpLZ63HCJudqDLoNJqlBF8AKC2RRFTILlO4IT1uqT5+D
wAIo3/uMg4r6Kw7pr/6GaYKoPhTDayZLqHNg9URRjzioFIJNzz3TR3hyBcw9Vl6y
AjeYuAIpar4MbbCwj1C5CUhjsqYRVJOBxUzmZBpU1WhljI/yEx7AQ0WRYN6U9aH7
UQljwnK5GOaaHDfCVcGsIyZEhf7LYUwX5oloOPy5iBKBhIiPg1NMzDWFj538Z5+U
5jCfRGKKu++VGvGi8k+JHj7UaUkOPhMc1P37uUlMCw3gAd+seTFnfnQ4b7Dzk76i
DG6NUV+U1BSv2wjYiadI0WKdgll6UZoMUA/S2T3bUn+gu3Xrb9dPd+2dn1oSoS9s
LV1+7IrFNlrzJTD4d73/gy6ZyzX+brknP98y6db9hu89YnQl7q2af4qnayBEQ8+V
Kk0jzJV5hdEeFbj7CzXTPFnHq/IZOZsT6NAy7+VeakjLP3RsdoTdb8mS2x2fUu9V
1u0/FyKd9adtHLzV73HvC75lnzIYkpgFWrKc8VNNqujtORET/W8GRvnSlKhXMaKF
CepqH8lmh5UQ9HlbAAbzUoZsOdGQMQOV0c+cgIa887rhGgZoff94B/PPVA2o/8q5
w9qEN5o/M5xG5EEpcUmTw6sLFvRlKcMG72bbGR7bZS5niZzWxLMKE+M3XJKulCDp
x7P/HOmLMCxnI4AAiNnUUSwCYrxvQNK4ZBOvV9xLAryRDKCs9yUjcqqf7AlepzL3
i29ZfC+5sq1JRHT49p/k92lUgzCxfrwWkdQJcfzUmzt8Nb08+aUGehvBAjVwA7WC
9QSGwZ0lUCyDmL1p95KTjeyG4il2sDSKq4uo3uFHdVXlPioksTjm5AYIOXawLdp+
heENfEjVQvkhQBp4NCQu9x28CqIuve+yVjo65x7yR5trbZO7flKQhDPBeju2b/eT
yUpZXFWuTjl4gq795t8ILWe6d2eO4jpV8FWnAhclAy3ZxNDL8azX7L8V7R6ePr05
zPohYqNgNgKnV12HhE33xzbOOb8uJQUSJqsbBaEWxJWpX97KQVqLEKs+Du7T5n3q
TxzVj8xw79F1O0Lp2eacTtsu/SgnhLIKidjnW1umRgOzKWm+UKr71jD+50tBuNR/
H+H2RcaY7uO+vfm0tP1adQVy/2FyeNMCH8PRVm0jj+LggLDjnYpbcBPBR5Vnigfo
3xiJl8SpUTOI7MxWNJaRGGF1teJ3m2ZoZJZfDNOURcHCnyIqhOHk+5vbpqXMBT3p
ymVS3sV8MK+bi9CPA/NgWDfgIoWHwaaYX05qnic/dW31fRMnpRgwr8pocjuDFDr5
UUg53Dt5b4EvCZ09NCgtStbD2qcUuzuHwdbBmAZwZmYK6SYGczSHGmLImsV4h8U7
HBXId2FdLgiUKb+/FQOIVEOOMv/kol0RjvPTd3qJlcIcRJ5MbLpjL7raf9s17ZSg
cR1IVn93bLw+8jRN5bfyYqBwLNMPhHhiXqqdzuNFq4kuZMRA+/cGI8MU6eK06xsK
ahdVKX+41JT1IiQmcEa3mVkq5mYl1z4OdR6wtioRqggDAJKKrK6KJKgOkW9RMEio
njcqEdb+W0+/nE4IlcfZeA2vga0AJOevelnTgE6Ze4O2O2MdSRrnKwPubqJ6jha+
4l+vPxzQDxqXOviM9/zT7e2hcHVbskym+nRJSNmIqfMBCWE1TA8qDCSw8bniAjyw
HnS9UhHfjNdSfzc18S0+O0Cxcp6Vn4fvUwBpbT12o6uOZLZhuV7BH3X7nn/epPsh
IUAqEZaHEgETeSevEo/46HXp8kSq6h8Upd89ZNRekuDJEKxo1k6h3MmwN+KLLVym
UJq89dTb3kCJ4t1pq5Pp28tFEgTjvNIzjHSAmpeoWMN619xcdjogjwTmTwzg8lOz
MmMo84G4i0sXfLPMSveS233FZ8RuSegaQGN7WElzS7O0zMnjdTnU+J/O3CCoRU59
0GXn3dVRpbCftDzqOC/lk2ZnYvvtIU5vSlbQkRZx9tlURkthy0iJhGdEeV/OQ/ku
IjHEggv0AFonSo8JdUUjeeOMLmkPNjt7vcNtfXc3tlXALhzZxd5yCYWEkxap16JN
Aphr+bOJPd6dOYjBrES5DTxpMX+oKgEA5+eJoBibPbjoTE9lHmPuzRkJS7A/kNy7
DD/fTqXxzr6AayVA05RPD77I3W1IyvecFxP525ap++bnWNo3iC1hdHoNRpgi9UFS
3KNjTKuuG8tWaoxGR84SAkNQbwxHKU/+vLhvEb89yAH+7dDvIAvKcfEDSpzofnBs
3phZ3h+MstOXvy2uGSRVN4h7IxE9GkSkcA8Z+7Jgb4ZDxpZ17t/+7O044Hv4yGJI
VXaLFvtTr8C6+hLvHrQQSpg40w3A69hLPM/H26KDdE5vdvW9yWCA5B05GqCD9YzE
JJactpHHShNbWBIp3R2bbEIJV7+2pB16wFkxkUFk1RVyNguyyPizEx0/rSoXyoOj
D7ruld8itW5XBCCtGjHrtfCsliuvVrR2hoJZ4VJ7P9vXXjnUW+FeH5ybIQUF2u7M
q0tnLaw1G1MoieX2jHr5hGkb90zd+hDlreZE9NJs7d3BrbwmjBYuJw2Skr1F+ZbM
kB4NpdVjekfoizNprZ0DfOppQuN7lsjII4dKBwMcHZELCnpYXyDlzzL8qLgrUBgX
v5crK40NILru8QLyw5cAvUXnsL5cN3GU5iCWUJiJhIZ61ce/CO91eyyAJ+qkisfj
Kl4tQEjwlqUgYLft236OBmSBJ7k6VmvW+Qd59nV0g1+BNBaN85r5N52z2ZWudJpA
MuJrFBoFYl4nprP/Vn5IGnb94aKM6EGT20IWOlUVr7S1Z6yqUyPa7UpcD6+7S/gy
8FtiRlV8NE3knD0W91CZ9tPRK7YrsAQFE2IzCj45Jxhu2OhPlNV2GDk52V010AMU
ivLNYpb9hA3DecFOLODFZjpy/6MVBkPNs8++jQE66vXY8H3H0mB7+0vfn94JrPqx
MPXNKFzQlpBNpZW9Afnv6CU6LGysI4zWIozQWoTuS2hj6cZ7pPsru76X6W/EB9lp
ACeuEj5qgTmfxteJx9W5lKdmN3NkaFpAm4ywL9sQ6DrH2Qc3rlcRolLaId8qsMnb
6n6KRz/BzFkK3P8XndbqBz4zcmg3auX1OyiVH1uR+gNL25kdYZUO8qQUXCiii8aw
EtqMrQ1l3Xu35frMxoJ/hVsuEYeRYx7mfJK7y1VrbdeqyKYEJtGOa+E1tBT2+35S
pHYnnDNAXEG3bXJUOwHA/QN1h3M5HBA71uWcw2oJWevGwWDcg++OWmU1n7VTnEbH
bp6fiP51QSxZgu6bMphVb+lIl5BYNyJ2cjYbStzBLhI7E4NUmQBYufk3GsCfrsSt
KdKtYV4x3r2gMTxrDUV/oVhzxX/sYarpWPJ26EfB4C/BiMWX8CGWZqapP6dKtb8v
kPiavUBRyr3fwsFAtzEaPP9g3W4i+n5DE/zVCXVw/WpEUp7NQACYqs6btyWRpBg9
/mwRcAUvd+tQ7L04/6ipNAPNxUEFF6qQyZbkiOu1SQFVa0sy7x8XxFDyr2zNLVz+
u5eRZPioH7t5uYdatDGnKN9YGQ80debtXBtP0Cm9A+R87ZJXXg8/4EAHkWwtB3qV
VXnDWP4c8Wz2w+U9U7CI1fpadJfmXg0uCM5ULaXtC5tZ6PZKqBnDYlFnZ6M90N2o
dLEzxPuID3RuJ+TqBDxywS0ItWapau/bJO9fvAq64dXatMn9U7/YONkU1XsblrFc
bYy+o1J36HXyBKxzsO85Lfr/Yw7PfEIPKliGxZcWcJnL0cPYItGq9RwmGA09j2Uq
CVouxC3MHvX62Hw03/XZ5RDPx9sA7uEhuC4B0oTY9pXAIoTsAXoAkeeVQD83noTU
TyA2fGNDJPjQAlyPL0F8pBos3IBaiGiWUkVP7axcjuPTGmw/H5aYZcrvUcNtOGCo
bCCPK2C2iGrBxtLyV7ZvZ8SKtegyRSWGlwLDbdhbz+G8i0EmDAyMwYN9nrLCdgPr
xmCCy7ZQYLbgp3jrX7ikDSXNYxlWlAK+oEpAA6ZbeAOnojEBcvA6mGG76eAncTnU
45wxZVHNWhvOUfxUhGPFT2F/ZW0bZi2iOm4vWFJEpw28BPUGBObFoFYiI4tE+15T
wNy4cliUCr92JnHYMu+C0+VF0wX3GpfEj3jq3a1p6gvtzsyg4kePWXdfyDB1KSfu
u4PNYtEnDbLJ0YEuVxcbDB/B4tEnn+JDLHrky+HoxSt+MEsSxD1Upghl/s2+2zPa
8oDHYE0dHOSIdaBrC0Q5rMMoiPO+1e1b3/kE8P+ax2XgJxIrAsYRy0zIkmRAlLYz
63gXZddkhZgx/sB80PQiyq7oHwZNcoEZ7DnE8iCdcGRwrjbmA3bHFbpc0aaBGwwa
nfViNVTScP5VkTo4HzIwoRnw4cSglvlcnxv2JrxWKnIbxn7Gq/KpgIZQvxcAtbiP
lAo/qLdS26SvOLLvFGDgocwuvsChDmTd5nsOUAIXtCsZ2Df2vypGFI86/aLSZoOY
1cSVtVzupokwjKmmz26CIJk114z6IkEVx9F1pd4kXn8YaNuRve1nDP2fwOGCLl1I
K7rKV/2WXWkhxtv8Ky/lso5HcYHRcQgiRJiIpVorGGaYoBTxUiW5qM6WeiO+LN11
zPICIFdIa9wE2djRX67RWT0hEykra9OMUbsQVEDLvepcXS5BHa94i+ajCVnmVlOV
V8QaVruHqwqF7p9ggw8DCrzfGTIKCqIz50xbXDNQ2VlO/6t0DQCe05eHE4i9GBQK
cb5M6mn8qkj6gucZdGw7z76EppujRAJzU+Kd1YtkDnwFfhS7Juj3qnQxIJhCkBij
O0MgMLhAJk6+tnt8F516ri9WkYB7/rIFmx47LC5NrbVpLttFgWuGQNBN/81jpmQI
+Eoh9AZzPCaW8fyG3ZoLQHHKWg7gLBeGKiahdY8LYD0Iv154cB2nt4Xw/WX1lPNQ
mZ66phbKA+petlk1Fyg41NJUh8fCkQl3bvtOup0bkZlZSm/CTduxNrKtqwziDuRx
1Y+C7TsGWb0mFPThf46q2yA29MukxKO6H1qG9GkQqC1Jlxl/PMnP9CUvZGOzZIBW
vbGDYk3IXPXWw8R1oywsZ5Gmy7rLTXPccaASst4hs9erh9zBNhFh4AThw/FpqP9C
IY7SQBgxVQx0AEXRLKW7mEAfCB0xw+b0ml8X3rSjOLKkJOC0wG24uiELQETAsuTJ
MmkGrb6T3cbUxM2ZAayXbnVjMKBTVUSaqaNCSPntLZu1gDX1wbzkJKNCJrxYUsT+
Rt+yrKSAxtvVd1NlTJ8xO9k1pjKxydKgH8zIPOOc9JzJpO/YuLBSJIOqYnCxbykc
hGj+SONcunWQ8QSydFBPPmHYXC+MYRAAFPSUanmpJ61CRo/sLcgNqSS4UVpeRHOx
MeioOnnB7BiadjwIqEui3mxfJWoKDqeVrHwyU+Pq5yWTnjLuuFM1r15aa/ugMo+e
gtOf7USMPSoLknB+kBfSuMVdiOH3cNslP6txoju23PylziutZ/Jpy/S4UzfcWR07
E/YS1aBmlW2dZHpDpX8ZZaIh8uIs63VfrlbTzr/jdS0ZuwuiRDNvDa9ESe69N6/N
nWfiuaMSHytLt8olvMziUdqkSVev2w8fSjqHEe2nxetBozNED9FBj5SD6RH4ReBm
xRviy/SAN9N8HzoXjz9gM/heKCCmWFcy6dO1xmlnHm5zeygVb6KIZN/WsE8sD+or
d900In98HxIeR51sGYlx4BjKGqoyGOJnO/7lpp6LfN9gcbGV+H+3xfmYgS4H5BTS
YnhCGo/+Lj1cb6sZMI2CHvNsGt9PRnCCnScND5b8jj3tZhpAKYPlN8XDMp0Sjasj
APqbD23DcyJE5aZG6wjF4D8uaWYpxhVRntdEy3EYvO1zi2lCyuW5E2tVSsvxibyZ
sAU3wq3aPmBsHIJ2651wDTGwW/tOhn+grcMs2GGIcuEyya6brLsmQ7krClJHc9x8
a08hXWQ2TFoAdQzNp/XNuw7J/k57MsLmlCn/71TrotxDkGmXeU7XsWzJiAtSD4Lh
W6dkWhtDWdbp9b1CdJUDqhZjKJqPfzUPt5QHSPhrfoRpYB/8pc0uYMsD4tAfLDoX
HSuYBMahWvWVSatDGrjgxsmfB5vDap5ph5SlaSpMMxRBo2ueLVuLxOzLjIdfIX/u
L1z4ieCNTKIvIj7CxlCvI5FkxAJ/g3qW55Mnc/6svRXUSor5h05+V5wReb28B2L3
WQ8EKIevw4VZ2QFWToW7kEmnLWFJOcjch1UPZ3P5JqrI5y7PRYYQoWlpWYWK9akG
VqhETWHDhRxYbdmVmL7AFf9n0IUrleFVWInOaqQHVCMN+54zycOKEgP5IiRc9E/o
Z0DbhfqF1L+UiwnG8Bzpbxr6RAQ4OBCFybZANyRESxab4ImZ8xC9Z5DF9Xj9QkTr
zwXDuPZqkbjDp1Roz5OY2uUKWp+Ws1I18pQL/klX94OlK3vbg1NwHU/rV6CSxQB4
Al13y6XJnQxUOQ5k+Jd6Mv/rJ2szn7CHzZkRHofiSecpmlgNEsVACU6Vo3k6kW5h
DzsTVhWwRqa+3TS1UYHKapD5q1vchtxDXchQD/WpuUSOD32rCxpw5ZQPxAHsaZOi
M+QruXqHDJkyhUiM+AyjAtYwmzTG8cUpK3dJBCM96pzzAWAR/5RCNI3/KbUiZIOG
5zPkcA7BcoyXef7WCYgeyhOh7OCiDQ/Bja9nH7pCRnzmO6Se04+ChSla5MD84eHe
bYhiqKarmF/3lUnEMObSYCWEZWrcP0F8Ft+yj8nonDpWyRGNGUTw+SBjm1zfrnOZ
JI3ZnbfZf4BWtZ29QZ7XXMKuKulqHpwetn4suzTeEGsD0OeFwNcSZycqa3w5FZcd
E9Vzk/gl32ij4aIOrQ3sHjORfZM2hDws3YIlfuEmT1/0gn0FqrmGGukrNbtmoUEc
O4qC42PpAuszI2sFOany+ngbcoUk6/VhA2AKAMB/uYLip/30Qx0ZMgaHE+XpqT4d
4mEyGg5CmF8S/PKhAPJ250XtW0zw1Uxir75JGgrzrCuq0eDSXjUZsVh2AtG+IxG6
yubhzTOLivmiEV0dGtzkqsyNklUDdWMbIFjXdfpx6B3DJZgyQ6Gf7b7V0udLOEUd
aLb3RD2PIZyTH0OUOdUjtBYgWj40mMmcWT/7e99Sptoz+StVvfCwUWMSiMqUl6l8
qBsIka5I1n0Qqqnkwj+H2U6hfXEY/nHRb52F7Lc0cD0W5aXExaiNJIPY5SAu50Wb
LWk8nuZOkdnqc6S6PyzX31F7HwHgZom9Ja+5RmXZA+I4fFCUgO6EWfRqJsGCz74b
+lwZzd9enf6uDTIsL6KWq29CU3ZJSMzAGOBqKaemKAKZmEmNRqcPAo2kNS9IhQnN
Rzb+SChWtfvBvdGJuFP9Wxoi1uUBA7XgC9bbLLT9Za55NmMP2fqg3F7WbJg8SHDB
1qgWWsOzPJeB6BZHBtIk2QSkifDho6gQwY7hx5gdJ8fqnWcE2jegvKjpbtxsvqq7
belnV+CT/+jPSUitD6eGmAlVYtH16pidFz+3Vs8HMeqdASzD2zteIGoswT75Wz8w
Vxts/qfsTI9/a9VBTNrGHnnh2AY8fEBZVF1m/5n3TtQYqIATBXvIX6u++T2/qULx
5gz2u/Y/Gaag9k30ErltMYSrOEpDdMfCxuAf/M3yTyE+gM0uOgwe3BcB9QGTVBbS
J2hgaOJ1QsKfRS1IYnbuhEOzr2JbqQrkJNT0kP3eoNMKZymhJW1aRyR3y3zVH2Bi
j6pHloDUDlZSD08ffUMPn9NtNmMkZVdO5lD3rNHObv54tFEcOCsSF27Ks3CPV+op
4rkWZuVnNyjPT7Cq7lmwbIEicT9YN2K7kHFgRB15hcrxgPmEpkRLvroOP8VoS9wI
fxPcGziCeFsukE/5NmLATDRgNSwGc06Tz2oQpou5yggeghB6WoecUeqlYr7dz/DX
18gXnuv/hWFszjseLQpzi5rPtUIJTvVaWOPCt0BHZNES05iIISJjxyJc7o28ZamU
e1RPqjfYoeOrA6ymRk+HO4oI5is//ltkMECw7lBmOTSaL9rxWErfkSgFJ7SML+v6
M1Xc3uRHx72e13w7lJPsNgAf08TVGq7DpBgp+2luKiA2AfDmWclz/qVFagcnMAft
0wDUpQsircFETjcy4bV1F6AgInSpDFkaJAF4jTkPaFyzLtndd8vrFX3ndPzokt9X
pPapHb5L6s0NLteW7Ii8/ltpgaYuMHsEOcoXcLGPDdE3wIm/kScgBqBLMhI729yK
6tKDq3QiRRDXz0hksOGz76M2ilbosZtQqo7Wp1fyBEwZirleg2PVvCo7bY4b0f89
1b0pnJxBDo2Y23VB8Q+8V+zP0heHu09aSXahxFtQIIj+QB+VO/6PPNwAwdS7225x
4wNM51dJNMyoH2zNnavM3LOa3aHcb+Mu/TpA/w+1SLHqoFZXdFujfi+VPxBkoRFM
sQgWiRl9jpT5hGkoYJBs/8HU9suJTeOvBUdrJ1ht1bw7EgxVJanzESBWz57KL0Zb
V5GjTavxv3zQp4qnfk+pfeVZWO7rIUr6g4I8D7XcfqYvdUu1fdINxAzMo2ytJxfx
AvTJG+gRxAwqaPGuCAu1ClAC968Yw7EznBFvjLzZfrU0PZiMsg6pL1e83/1RQiPn
oDNXuof+ovUn+guNxZ/vR3l/LKZceXRJnXYu9RKJTenEtp4tGvRSyXHmv3FtNORM
K/EChTfOvH0GI6jn467J5CyfBGBv6cCE86W8rv/Tea0zJNG0xn9OiSp+ZhpCZE66
D6KpuqvDQqEzJClIZLCxnNfVEgSGyA5JmVz92m3WCsqUOVvsnipQjrlumFU5s32m
G/sf1ynn+6BTtA6VKzV5+S3+H737piTUc9H/WpPi4QZ9Kkaiyl3j9iM7TrP9nfyW
BvdjTNVXybZgnvV946qbukfOzeCl2MHgaML2+osvPn0tdWlScL9TI8ZC05zQDsUS
i48byA5YzHlmNgM7QbuBd480ckZPEju2Xe5Q/655zOopEHOEDDHAQGsmASz2Og1c
t8BKmY2XCYQYQDOBziEPygDetB4mMMSPpBmYOk61SQ8edB0vzdf81EOdO++9d78E
Df00YumMIZNIUzrtl4HBmKzmibgoleGx7iJL/JeP6MzvPJjQS3p5n+jBWh4OqnYi
VFPQds2jstyk6f+B9L8sOtSAKRJTQuYVfTeUtbpdbTg0GvvSQyJTeUTwtTCuKHP7
s2hOnfKhM3zCEbccsJeqYhHxtWEQIzxwZaJDAkX0Y/XWie5G5t+Q+9OADBURNasX
F7fRJp/4jaDkcM2u1SaKvO3Veyp1uoXooCv5LStS9cjijuuQcgcNG5t1/gxKFHzG
QHeLM2DTE+fPTQRzS2HcNeT8aRj2DMkmWm/U3fwFlwKof0x/66pzoF2pQubyibYy
pVz7nJH+GMIzf9LiyWE9LoNKvf+YOchJRhVc+75Hj/MMZLxXJmQ7b1hLnYDytBa+
kUTKF5lNsl0fFGJlPCfuZuoKsgay/AyIPc6rOD97TbgYGTjFdbPvX7pFVkrIkkNk
8P1qrUUpISjUGtfOuHp+7vCACiVZ/o9+Vn4rqFaC29/OvAeWYTzBL8cz0FRGnxLQ
zzDKJFBNpB3Wi4DWdGTIhcqFd973dOOYFRNeds0MExAjR+jBKSJ/o7RTqtlyoNGy
7aS7jY6Dg6rhm3AICfiN1mpixJK9dHiwAGyI6Grige+fkBq0yQ4BO9vj38U4rzbb
cuwKiDoifVdzhW4tuGLhEFfQsDV4HFfAhtAz6EfqDiuAXqsAoUVwQggJqt8DE7Sj
OMzacm4lhyS7i2/LYkBQ0Ixfs97Ogi3TEWRBPpvSTkCnXtpdOCBbPfPzypNwiool
e9AeBcbEFrvbveqPO0bN86Rojn8kHCn7WSpPFAbKapS4lPzf0H2GgTNXu0bDAM/I
Tn7PO7E8pQNFVKH2VXVoNkf7NnOAov6FsT31AFux3cKbPmvqX9544wOKqQtsls8L
USN3v1esE/Pi6zBuLeDYFhwU+nBZa0I3nP2heawqUwiI2RXJ4kOeIhoANqVOgrCf
wEgzAUWTfmjkPnp9Y3TxCFTvDthjX2GmZunDr3vAuX31TeOThgW5jetVQMvoVU+0
CulQCash9jo7do3hlKx1Lb8P5daPLcjl9SFQluuC5Lqy799+1t/figbqkYO20aKp
AaxfO0hF/42jdWL/bEvldE9bHOR5Fkr1JtAkgYhgj9ka0+DdzVHGwdS83Q5ctwC7
98M/C4fZ/W2rw6+9gF7X1u5aIP5Z5NJnV4W0CqphrJ6z3BzdKMGd8M8s6VudI+to
oT8HganmjkrqzFinckcFMJxV1XPJdotPMIkAtCJkACGFLwOB/NDC87fDYi9IAqhi
myLbE7G5mSc5//qEJDpKzc0i0RjvVR5oD35k1g8Gp2BWY1XyNXrZzH3j43tet98j
UMuq31I0jEmZ0UXrzprI7Nn/B3DsKzvPr/vxYGZyOw6KzTpBCi/7GGl5g0xZSua+
ACT2zWVVXanQ8FduRwGg/2uOrkLE8Sxmd/4C/UAbVEBoy/Ol9PVO5xN7WHhX2CXj
Z1XlVo/d0GfH2XyBfCTD7ZpGLdL5wdmb4r/j6lDU6mEQfB9xtvh0mdMnl+3UWhx9
JYMbn7R2oDhyytV9ePsoE7NegtcTBv8DMKZXx0tT+YAYAfHRQdveL8eCuAD3B/hm
tAhVuyQQPtorREzf29gbagwNORN9w8YXNYwswB2PaFDFUsO3dFv0QALPDTIJtPOB
qY9dfMikXNtwua5wHIUSfl/7K7K88W4NgPSXlC82rVdrPc0MsCtkCcD3DlI+J941
4yP/Bvg+PA6TG9LXs/YqD44Z9TgQcJD3vMfRWmZd2DQWS6MTrPup8zrKEm5vlx3T
CHg8j5pTTqi70sbK7h5dfMLwuog8h8h8F3Pe7g46scYBdG/IRM0k4JBqm4vBjoir
/4bNxG/s/Z1t8Cjs+vqtcmNIz0V2XNoXZlfROGV3HxRdRRpF9O3aNeoqgh7udhLS
Q7XmNER0OwWMndUft1krPzojigKdT+yXu814WbyQKDfJ8XQf2y6IxUkiKdL0uIPu
p6o1PnLTRX2YsW4ODQj62nT6xajSyC8Mn2zzQVAvLbTI4WmDsgg+ORjXgsQ7zTdd
csvTI2oWrLThWGqQrupwxyIElGqFtwPChAcLiJTlr9tw0grkn3CsJos7UFtk5l6R
Y1tFHyWT4WJU9RrLu0VnDlMbRkALFxSzzGnWnmUnT/6Zz0dPh1UP700udib31JVq
h+Qt1LXw2j0ohIQKPnAKVDG2Ku1nUMX8ir+1y7IsZD1x68oPqoSKGEbxnkewmo9s
FlYfE0w5XDyl1mZT5OpdFuj9wBmC6nPMbmb1jp8J7s3dujWRFVod1lMyTpGYanF5
8hRZRyEgx0gK/FYLLItDU9BgfN1HzaqBnp6DlH7gqq4KrUlVuMdmkWRt8RsuNcms
McgIMzZPpDZegpvreVF1LIyJpncIrqUbotej7LFxgIKHi2P1ImVsKdPJRS7U+xNi
U980ZEl60Go79aaL9GdnDaxnVk0VdEbD/9L6MWgBf2AzsueDsnoo4V5I2Ih4fdj/
Kp4gfZT+Ul7hgw0sOAtKQ2nnbUdU04rucWv33c9thfAzbKx4E6dHMkcYIzmd6CnH
YujoN7ZyPJhsYqYiZnePX9QpQ/00kr9v2Boilyr+yARcdfZe0NFsTR0pM6CTRQc1
w7kRIDc4nmLWeQSyteozKff2MtV+XfRM5QvQUsF6Sd2L8PjBIjDJ24n8nePo+fbW
7nqT1t2C1/usfLBbY5YQf1+pTZwKWV3msMj5ICR73nfVa/LyyeKONg5IAwGGmHyE
FBXt914/IJ14qq3SUZj2q2W8pgSiYBKQCZdXHdwdtO8bhYqlpY02mdeZ7qFK2XE6
CXHebJIfoeSJHbxmiNZsK93RgzqfPgBt4fI60o9eKj85jck/UvVInOcAiuCA+tvS
u6kdudb234f4RbscwenuGhR7HKM+zCtGQIHdZUl4JI8Dl9v1pnjN4+3sY5Ojk5se
3WzVG9fI7DndDVSx+aokyBZ7KZxKZQtO6eChuXyhreP6PFx1pr1/ZqVJe+Tmbb0y
vCHIlj/2BK+dP2tqvPlLn7oW6K+3J1IJZFg4rrZ9E7lFbc4hcZtO59+D5CMa7sVr
J9QbmbXQKyOxLSwwr6n23ISLl1s4qTtwofgZSQpkdll0NI5LWGWSbIEbvQCxKibd
r/YUyyueGNNGEtG77sulQCXi9JHFKXc0LK+6XpLBvQf/b4CKARfKecPc0S8/IF/X
jU9TO76JlT0LJY1OQ+Ova4lLsAWWMsuC/x9ncvnHOmv3rGe80iwIhIA1orWHcH7b
8SD9vjnmvMRsFi+wvWw84JepSh1qHTmH6bZqG+WbeyzNTsCXzxuUlpDnBCEKb/Dj
BHRhebAdUkCvB1/sI+4CSGFGe6JgDb1mVNmAPq9Mu8OgrWoWXcR9uKOdBH1aqUkD
iP8YsjosTyaqOuuZ/i7oEt0uXF5rfPSI6DXCoNdiWj7rWrR1xfFQUaDUKxaxYBXy
DCoFLbAp9OYPyuZbwXVqQIIwx6v+yOA7JNpmHwRBHDVBin//m0k+DCxAn/AkJTwo
rRRSPLmDeRVNwApnO8ek5qelJn8eiFQrbALIzukkMiDiPK6fx8A34Qe4rR6W+fKy
IUSJKde44RZ5KxYcxtCxGlGmN52Av7ax+jJ2nvx5MRAQUtQxbFkI39uuW8vO3Fpj
PLHc47Gq3QeN5Tp5KJm1u9EzGTlsjkD4sBVg8YkgvGfksYrzZcVgfdmlucCEfIZp
EjokHBjNE5dEktM77MCMT3Qa1QFe9R3jlpRdwFN0PnXygGJ8On0R0B8ZUfotb3/y
yWYvDxrJKT2EZHgPK92VBtBR8Ect6Mu4UA3tMCuH+WqRGCLKeJ0wDWmZdolnAlPz
k/QeQAZLEVRHS72jsjaranke6gJ9uSt1HNvjZljq3VdLjV+xd1tMd+crLGeqgNr2
6zEJ2ofUjmraIZ88UJBdw8ujigPeIbtzGz9m8wm1UBAx3LIaa8WJzHbPZSLKtCue
T2lPBy8EO6WJoT1BkrHu+r3GJuQF+c+1mf6KGoAUPN7DWKcY6apyw+aK3zUtDGzQ
WmJi7b70eJj/B8UFP0UMhZ+cttdymAQ6VhUPwwQ8GCBdAekEogKjQzcA3BjtmFqd
rAzklOYForZXt7qBW/uwc+yEoD1L5oDVp2WAKdQH15a7k1gJK/J35lPjwSkkYMTv
DtT31kFnR+OidZhnv7hwos0qkn5YbUV9EgqPCBikbKcQNLc6znSpGHdhgPvOvrrU
MOYfvWZAHVg16Hiz6UgRWuCsZjMxqQkimMbiidir/Kfq/TY01Gc0vWfQUCdPVYp/
aHJNbbDqcLoPwJBkuAq7CRiaDdCF6ZKE70HWp7WgMzbEt7iKfXtcIDP6C/Xe7cL6
eQ3X5gpb1OFFvkCJ7zp3YsMk1DZoqT9ZSLlk4JQeNLk4uZVRI1q/O1dTIB7zPdvV
81AoZcdcolqSLfkbl9tfSBcO3hwWrakejmNmCyKe8kBcEF5n/jgWymLt4Vj6OpIP
xdnAkhd0XlZFqNxdnZ9XxfahaVQMflseH/tqImFACjwn9fyA7N8pjcdJlRJhYmA0
I3Fzerhmd/6wApxR7rTLbxheDazhoaGCf5fgh6pE1mJoA1qCIVJTSel2xtfklD+4
bnwV90pPDJ35/e24eHsexKU3MeWXEpV/RIqOiOXrcen0iNRnfgikjkJvmBbu7yYd
bq9wBQEqh2cwKXBo1NVHPQye+so7q7pgf/91QbzjF4C5yrOG6RWK42y93tLmLorx
sv5WGovRDb4dAvuBLnqYtjsnKEZqjg4c6czYUcwukWK3xK8NoE/bTiare2sFoi68
nsFp5sZ216GtmDYXtwanP2z8pvFeI4P8mA1HtgrAcp9x2P8pJMzuFXzEDANp8gPD
uJyrYnUt3aXWPpXfi0TGmt9rhiNxFwpd1HS+sxiZjbBe/Glo2iqe6qKxB4hwd7yH
fdmnsTgqpZ4/X+SqImgwCt+AttWdu2wFbo8A3ikC3Hy5k/W3FE57xk9oE+FsuuzD
Weo05d1P72FHJDtvQu49/6RAjxwsiUD+K4+yzhQpTI9C4Y0AOp9p0EMhqotGNctw
IwQo+v9EfX4fW9txkxINzXO1a3L/2xVI5WxkCpttsH8Qn0nkmJS6DaghVD+MHch4
LihksO9/5FCv36TE4br4bv85oO4aYM4XRqtCFIPCC1bnNRrP+KaLftd7m6Yjb8OO
i9R+G/aAuarC8/WNgnaGJS7zHqmdZK2RRpM3+din4ka1lFrGOAyXvkCbPLsAAYx+
20Dmr47/5f2jTrJNlSqZ6oMKDbcGq9RimcMlkEUM6YUt0mstMH6ulZrxWpoUqp1j
gNvj9jeGcqSmsK8UFbij3SR3WbtVKvHnIqKDNnYnGe2MuLEWPYgc8PMRMx3nijNq
dyu5OZsPW+faVr6RjBY/YB1yaXhzHL/obFmEN4azyEzJM1L51sdlkPX5mvkNJOqN
svggUvZlHc1TeeEN5AWFeoFwXV6sgDVfxXPr3ra6+KjCeWLLqJmrE3fYZTYwj9L5
HrCGRQZg/t4eXLVTiAl7jo6yRRUxT7SgWSXvZSATbSwYmsSPrs2ETbmNnr/hQPhy
RTUtMEsHEgLDo3EmHftptUX0vx1r8vXOUXx2e4wEnpRSjsL16MIyycQdgPPwfUmQ
69TrI9abgU/hsKRJAXJszy0k+ES3i+sp15ZKyWB6AOtlTJvkrcYrEJEjB6I4UWjN
oRKt5I7vrjaCGsadz6mo0VW8gqHK62DykdJaePeK9I6p3iiJmZmbSvV6n/M1tL1k
20IioUFkSpiJIce1BG42TSzo7Z+u/bDBFLRcv9OqB2Y+4MRDRhDea6DJVXuQDve8
1OKJdzS2Iu7Ss34xq12J4bphuCohkWJtD4tFCKZqSdfrC3SfACUL+b1OQfaT27Rx
5ZNb4+8fSBBuUt7bih5wZa9HHbC2KhiR4GYdtRehqCawAPfk8ocG7O2rQMk1fSfc
ETSpGFBuH88qEhsiClHEohm3/WqfR5scAUx+3agIBsgUWJOZnOcs3yJXmw1DXgZO
dIyENXcWR2cFjclh2Sj2XyYyojannnQnrqRZVIy5bRwMs5p31hnoaPuvKpSKPpi2
tWbo4si+s8GF/PCSzNEPbE0v7cJRrAHh0eVV8b8TcHPwawuKJXMHWwgXpkwUTTp2
zaw863xE8zuqSzXYPVxPXpDbh3YBjXtt2aRt227VfpTSR4MN6hE+zIk/xh7sAv3J
1QGBijJqWXzQvWTUjc+6plpfuGtZULdovbn781YDdwMO6sFDi7t5zLxv3ZQhSyV1
zEm9JBT7ybwUwHnvJjFXZ20KWccdsDvuPQ49tE+iqAb4Sn2Rf0KkUOE2CyvziKC2
mWSLRqmAnTBkQ/fGmfUZOk8NHKkJSzkbFRWRkoFWzVfkW92xASppkaa7U0q6uzX5
QmZUoFonCfNTfJSdh4OVy0k4aM/5fmt1fofUw7PjCjZa4STJkSX1neRPNWPsM5TX
ZqLoTqz6RYAKeMvylz1kQTqo3WV45T7Dp9snxUjymYxIDyhFZKDUpljGzecRwo/F
YoSL5jaZ1E+2LqOtVcQf2ew3zc3xCJB0zNVMOc6MPc0eIL+30pGg5jFITnytED54
YT9mJPu/9rTKCTXXtziD0M/K4lDHV/Z8vBZJeBPqqM9Ng/PW9BlbOr6vc2TD1IWy
ZvMZe/cvSCAK4ieyVVAQdAy7m7Snra6qLXPxArU/Lem6WO8+AYR5dVF9hqJAe4HI
3ynPJTNousvwc6MbZZBI1gI3z81A94GqQEG1A//7ZFs6hFMeBcTzztNHgddNPFcu
DARIyX+1TWQu4FVXxPlNnb7qvhKfyiqZOwXXHFUwWov9tIDHy/uGiIEC/Cy2j8h1
m3cM0T5aRyFTrRTQO31gbn6xElEA9jxuAhtgj4M1DFRuQ/uWU0yueqvTvKwEwEYc
FQuLGASQOZZar1wJkWFIilpZpVavdYxW6q+KtTdbm5e0FhCqkq7XNGM2zAGXt1OR
uvTcaZpxbLt+zwAIqT5uLQB2TaRpElx98q7FabHcLuUtpzBjMiW61LwaunXMfs0F
MaL95nfXfwDHCCxygwOJHlXoUWUaT/IgM7qjwxMKRlW/Q7QRoldp6fnIVFj+FVfB
1RUaWe9+/GdrsU0V0ajuAcoevvOKnRjsxeYjtEiTJESllZAHRwUyu8SJSj62B3Pa
atn8SfFSFiHe3IZl24tpeixNjhwC7PLY9UWv0K4A17e+BSKovt9kE1rPVNLFztaP
PUfGYndKdfc8V0/QgC1KU7NsQUcmu+K0TGvgj9TUZOQf6NkeuRj+qBpUHyQ0BrCV
F4KqluWFbsnWNXeUmEw4ZR5lbB9N0om/ZQxzxrI59HtQMpWX2QS6ga7vE+pOLOQb
cdMFwbhsVfRJTMMDJNOlOoz9w8evcATMYqQGn69VTuMMxAOtInjlyHNjnq3qe8v4
l2ASAYfQpkdn1oV4XZqrWdfSdNRBcRbGWoRLLYizbnxQeVcxADb9RBT1BXIAOpC6
frTi75DYU0d/9QXM3hcNsdlCPwjLyOmnYFHLhwWp5Qz1AaEhcRt+FfrSKQzhel3K
y3xv6gOn+WpLG4Yzn4fz//W/kQD2+bUjy3ggIXtAy6aN7wZ9w1DVd9V4eZJXKY/H
Om12i/CY9KWBarsxSKbmjtiMNW9zabdgBRiXvR+4KhwxlV5ic4MYgKIPYThCddf3
o2dcykJRLX5lyx7F6lj2VcG9YThuPD5HBE0g6LMNi99Jha8OAYDDRcZ2TxsSgVN+
C53lFPQUxHRcxYzFFTeMxNZg3pXxoWiUOjU9z9MMIPXBgeRmyS88eaKo8XGO0ClK
GmCz4Cx1Hnhx0OU8u9d9lwQFa95vERpQ/7s3x8E9n0iCy7oEnolYzRU1NPrxxqs7
o08nyJwwmPvkLyuZltmz/hRnGSVsi1I0KjR4mnyQkYSy1ijQjU56SF4ZqZY6p5DG
UjIWFeNmTCW9Sz+H7Bkst7eu0i7T6rT3YsFeG+zM9PR3r+6+cXmUiGn0pnTriRMB
br4TX21j83OCD3xp7Gp1RNuFP2faFIl8stRM/GHJyai/rKe7flMx5yny+iJQ/Qsa
AdzhBQrM/hv2cMgyA2NkOegOs8h9KAR9RsaE4bNiu3TtPkXSQY0oG5tftKu0uRA4
nYWpUYjOTBvYZB5P69KjrCtwqwr0+++h4z3FZj4demBB4TXrVAPB2zZEsICQ0QJw
44tcgakFBFpL7rY1xqdyylIKNdPuzoGhrYKWV8CSjXNLip7bM2Gq1ugZPvchiiOx
XBmAiiAD6SSnsxjebPmRQQ//FlVf6DSRYhsyMz1nxt4ioR1ANtSyg6jDcPnY9N9I
duQ+1ximvwAFLQWz4ADGwuswadCnIk+10fwvyozJWLZqRrjawHaU1lmN5EYrryfM
tjcT5GErKcLsxcWYlWp6M+drqYqeZdjmL7KQVojSEQYwLULwITCeFPOktirSewrI
RjqdBZrL2XX1rjdTCz4ma3o7Ap/1XA5/G0WJR3kXJLeCgQ8U2dx3sFJWY2+I/F9A
WOLq01MsZNpJrZEgdHotUn/xADEQxAfhQwTX67M4whYQUibQE2FoP98f6H5NY598
0IiplFEKpmgBj43RM8bkLyt5uRNQYEqX1zE6CwKdLidFP8c1e6k9inkHPZ/w/0Fa
XoiE51Xm6rEj0VMm0RreugGpPwE/Gs6hhyTJ39Kdkb1wzu7hKPRcnPVBR2wHdHFV
fs9rl5E4/o2RCQOr8h7GLin6S5yGwD7utqD51EMozMIeK5WCX+wyr11GVU0T0alR
Xicth1nHb9SbW8F8S1OoqFFWHpTAOzC17yMMzOHTUkU+dAAJ+RzLL9qdtSQ29zxO
ALCtqWrKHJAnXOJfQNDVd4BVJ04V6bg1XB7j0qIycMNJENQWfRfRHXf3hxMgqMKW
a7yiZckNQMGwifXeZFUgD2hEzN59C0cNwZ+VNsK1l025324Pv7he/UFUYhOxq7iR
wecBX4LESlM2aPu7sKS2CsAGDIT6A6Yb8yUW8A6BwRykrUiurhxPdA0q6mOkDDsO
SOEZMgn1f4VkphzoCqN956+SPqLaOIQlohOs5Yoa8tLeAvimFSzcozOOfrcq+zZ3
+v9kzCAklwTFwUv2/+5T7oADzIlqPDtTjAfrNrl+8XaJ86TMGaa6BqfzC2oGwDNK
6KOuxzJwlIHf72ILr1vXPSs2XJW94trEu4aJuQQJEeBhfPyWZt810XuqqdHm3k8c
onW7PLdSLg8DotmbV43Bqw9ifmDWO91W1/MRfiIPfBdzs73KRp/UgG43qPueV/uS
5Mrth/Dy3T1mRXlotKb2EBGPSuor1VRsYhcvnK6Q2Q2tP3tGC2qSvAx4r1aAVbIq
MMSIwJtQLE9ma4gYjpgIIsFEk2gwvpZYru42+S9skGHfb+6fD6S1j6vQOjSnHoG1
ZEA9xgfhM4QCDuFEatQ+MHPPYu+/ZU9n/v2uPZMMxmYvGrENl5wohH1aKmYEAwjr
inr2TF5+VUeUVRPg+rqcDt9LvzkJool1FRSwdCykkT5sbUiVrVNn5sQv4WceKKSU
IVwMF7GZekFSazGleZmiI/cvmzOb+vHzaDMebTpnP1bDvvAQvMjM5oZnDGMSu/7P
aIuE5rndeJ0WWK1OJVPI4M5kR2M4iHedEv7FGjwelCqENl0Jak6/Rwd7qIxffdZ5
EGX5yqK+OVmFyEwjQl1H3RiuBaAuBAa70WBAdXF9wuBLXkCdufBLhrb77c2Vwsoj
0iqEvMPNmOw9pmfLulqUaGdBXmgRWgAdmxq1Zx+HW0BYQ9692X5/ndEcOIl67QIl
EqEeLYPaaWqKo3fXzZ19VjNuanQE1CSgkuNbVOseCI0UbH3XQG5rLAPEVpUvMluz
BuFlc5wqYkXJne3l8oCoXO7mDfbygI1UWxdkxBNEHHg+Ca1CLmkxwKzwEmrJKJ8e
3Xy+3+b6SnwuAKq+J/xvyVFV16SoQzTiG4zvpC2E9t3z7sxulmPeYZb2dQJVRPRV
EY+YHbFo0K5aTUv/guz3GtHXVrn4dHKa9L+pELrduwObXiM9OqjA22qp1hTYpTMn
YRYY+GJIxxhf8I7B7v1zOad4wzkTtJMvJQxR+zF4xiA+S+ZrPpmsxhH3uMlnp+7/
Zh9aLi59RyUTbnPnDJBxpcARzH02WpAVMPh5ym2LHa7KsiVBwMJJYAen5lKThhom
XuiCilrtVhPlUeEC3VuLF1whdkpfs/TSY0BCtTvSn2bkUrooyEMSVfgwBJ1JyR8Y
P4Eo2qL9DURsYd4p8Wmwkkk9T6oXuDwT6hztAl+U899foZZV9C2ilRdSw4Th1oRk
LE7CQ02hAMp00ZnCVzVZloFvIF8MxQOD8QK4blWHLYdT6v0wh7J7UlAP/WCAUnTr
3zAHnOXUbA/xut5zDfBC/+sUtZ+dxo08draPmenJMNnPazDK9PTuW5aewvuUQZSL
1uHn2x1g3l7i+YxRSsLQZA3SYUTXojPkxbB3XTVgthsRSugTS15MuNDaZOpuPkXE
G/7wX7HSF47s1q4rICmDy3Qqp34Ibl1Zhus3o3Sr1WDTOUB28u5utc0yMZgyBSwc
1tQpiqtyPMatH6MrT3NC6LWtY2tqYjRaIDW1+jYMzn9q4l7XlkwQ+878f7SymiUq
i7X05X0LldlXbygCa2ab5o41Ks+zsYTm8xVUP2l+bP2T205iw25fu/0/8ZDlTRou
3ySPCwk8fhjnyyb1/cvqCwS9YeNmmDm79IIKprMqcxV8D9Zd/igTKrKHqYzHe5Q5
Il6+vzsuF0hnshO7NNq0jyIAfgZkIRHtnA1I7gjMC6MxxtrWPmeaODAIbhZkqeot
gzfmOyC2nLkhYF0TO42sez/Z0wU1GaFHT7s5e3aChnAc/pLT+5fN1yJU222/ahD6
U3G2GY33DK47tqxmgDXO+2qqrQUN5CnfBMYFSIIjpkySqRE//aG2VTz2OeiZlHNe
wljax73c43C0R4Jo+wpzGe1L+aSRS2x9U93013oQpaRP+NBZz/QsjjRVd0JWuUmy
M7Pe96WdSnPlZhaDjnrRqhKNLMLgFk0n3FJ+edWTscl0uifZEKfSNYlGC4xRVCa/
uG0PAMcw3amZuACLxGDgdiGwlxA2yNdB8VOwXc599KPnem2f80pFHoe4ydRixID0
okjp8atZki1ScagCBqxu9Di5tGSmsssRQCwdh+RQaw+R4368vOWNoAUB1v3iGL++
pZeekHqfIz9jIoQWVzdNKigRLEf+P/Izc40ycWdUjf9e6/KkTQsDEcy6fEy1rMQ9
rL0UC81azDtZAOLeIMdMhCUtFNWJmc0+8AHrTaV5fPOCuNnP0UyPYak1UESRGodV
zndKHgSoB/LqbtSPcnukELkAZ9LD8cYWcuZehfgXCMwlU4K+PrPpAYPHZihxuIPR
KXgryA+18oti4jxVyWPCMRpUw6G8zzcrcFjAPzkNtEXMIt62lTJagRlrpUkg6W3k
T8ksBm52Spo9fKTwYuszLSmyJmjHkTh8GQdytpI5SbKBCNVd2+LyvYG4GiyUR22g
9oAcxLwI71D16a0++oor1HZ13v7Pq5n8LwB262PACuJqYfdzLO5AEyBj+aW819sh
vPt2ehsLo13Jozc3+zbwhm4fl37lJO1GPZsgErgWUMmydn5Me7X9WE2cWKteYvep
Eh6CSaey30d/8r7z9uvxoV8j1pxmrhLFjs/aMxpmi89QfuYOLSYkyUF4Ubtewp1V
riCkYChYHrJVuWuh+geg6kCjqw4l+JgqNJzxH7+/YCFaucR1GIKN20ybHV/HOvew
tFEKS6Gh6DVu+BfhGDYRKohKY/EK8rPYkIBsAu76aWtpNnRA1NuCreGMR9WJOGoH
nZL1XXv+DsmBI3lI0t9Raftzo57MNY/vyUmLOOv2Z9VlqSqVP9am4Z9M3FkwONER
Cq8LqDZo+FlZ2+Sv0TXNLmFoah9fWTux2u8HXfF9OAzu3TpX6Oft8o93rvlVYe1W
DOPbtND06uLVPZNtdG1j+2ZRyYXcyBep9+AlMYrUWh4fZLCwWu2uPrIxa4iYdD/O
QbJe2Qw8xloxM6UNiak1F1JCjExNKHKL2EDfvhv7d501Ilxh3YPzI+59/J/0kDJC
Sb1qibZAcuVfq55r9l5tP39ab+ihtX2g372K+T5j7sEcu/2QagQ2mTrtNnS4wD/Y
vXh9lDrqnE8Oo7NyKahaqeoD/8DLnz+Rv46/p5AGb5DpFhegHYW3ax5fqQ7SoQ9r
IycUYuX7ty6Jdes/nhVc8TqSV1qVDlZagwYYiffAqMEdAFypO047ivSwHw+30t5s
ACf2dn5XFxPWrLHimxfHr3sLJ+Rnm/+ClbbTui6xvZIR9f6TijYejMNp7cTDvJt2
8RyQOA8LPaUsLY5X1BtusYvIudOBg4SjbHqYMdU/siNbw298RJb7G7LTzfux6IGB
kg1oP1B3wJ3soqwqICYA88ESII4QNXOToC30Di8Try64h6zRFewrajt0E39GgLNm
vz0lcLR9SSBQxdu5bTlJq3MaTwMZUK6pJShPzTlr5MBgpWKYcw9F/0Mt3MTvBVrl
Kz+HeSfD2Lg5LsxwJzALFq0dNydMjBgzr12xFH8WCor6MNBoHD+aFxkljr1eMOir
xGglo94aPP5BIbujL/1H1il5OMqLTvjF+SknWeICaY2F+7MxTzS4DQljAhPLKw81
FAjRhrDHueYWGeQNTlt2s9GLbe8Y0xbhRPmb0qC4mQpzyVHxnn1SLTIARDRr/+WX
MgFvRTSWTWC/Zz7KggApcvK91WsNxeSEQ1cdXZQWl6/sryFqC5u3p9IWxuqWRavg
8EIPCwEUdIq9LrZZZK0Ghh9wi2itljzd1IQ9v2BhXFoTXvsS2NTWHHGZExwhH3xD
DtZZWveVWL3KbnlnECOYB2y/VbLUPh1BYVi7KiwWdH+FYP9ChBDcsjRv30AwOVXh
xiBariGEqjd0nKABXYmsYBV6imo4UjnBLx5AtlhW+rZuAQ6tOYBuW5DdwztI8PFo
VZ3XqRMzENzhG8pGJVYLNQMvoOc+L/ilq8gDoqJc4SsE3UPZws1Ut3XskTffdwG8
NzHCaXPTpGB6IBjjtRpyPdz1FXXGBTJGw4xV9MuyaZs9Tj8onK03eTyYj7ujRSbU
CWaAYVU5nTV/daAVusQfaZDfbgoF0wkBiDMp79UHiRMFDw4d+KzB40sMnpzhnqNl
9Ryc1xsu0FqpHraStREf70kDJHRlkO9sWY3V6I6qOGC678+NpTl4VtWjHq6Adrp7
Nvuk1V9ROR48JKshp+p45AkKhb/f0/kXxaYh51WI2mgaIWv31256SneiqAXRFO0V
tEgYjMGOr530C6zDEF1FHKCJlZwLp3eIMdvtEx4nGggWYoTEYyPt1YvKYAz2FP0I
tjcGa8WzIQFS1fVGT8BXR2s1SnMAFUfuxNzsRLBIUnPQLgQ38qLNChM6WZkXq9YR
K7TiLppToGAHOki/pttOB70GK27ivnCS/7AGUgGcPShhlTpXiPH3CkOxViJwu5iY
UYN+G9140oi0BOF67rxQSrhi646Bd5OpgZth3NJXKlLk0ljtmbvIAA8U1GFYj4+K
dbWjzZHZ11//aSUOH1XGqV+DURZpxIYR3oQSioA5kDaiLrVB7AHSNk8b7ajB0XnM
FQ/u7RNMu9C8mz+rQLE2CZEvS8PVPhnehIWhOsce3qjgydGXJLEsZIO/pCY3L6IL
CBbKEjAZ8Dw9KfIAkIPogiZQlERjfWSFsk44aYsq3BDWsw2i0jGaWPCm7aULrpib
QCORJM3plIOxxcyABgh9IDFUP9s/So7H1q7QjsbZPhDa6GhZkbzxhGWO7fw3y2tU
sPbmTo8Bb0NwXgJEEyZVMMRhQDOxVNR+J43PUeeRJ29FdZPnUaWp3aB0UkJrUcGs
N8tO5cxHPJbgtNrz+pew9pcIAczxYNC7LfOTYSMNCHjFOJQOSNlw5QE6T596XwX0
Kw0UJlcUSJZETo4iIIl2FyvU7ZjcSRUcX4Jl8scOjUX6Q2Ur3GGwn0+zdudTaF6Y
m4vcpn9F20wkiWjVwEWpVdI0o1W0yzQX0o7iQ+HDC9gAnrFejcQUnMWlErCz2TWA
H69f8dOBXOCEqK0n/sRjv0Hwg/j5QiI3qSC18BajAUjRf8ygN2gZyOdZIqZxXSWj
bhsBY3tNJITrbD/Q0h+ldj4VELHmf/TkeIowG/pVli4Rpcs74YqbPYp/EqcG4Jmh
GwLhh513k/+GooXAdD0DB10FAg9miXXvNVIVm7vDK2eljmNiv8Sw0cgNs6xGLvbF
ehE9+B1+q3FidYov1KT0IJiuf2tHh79560pFcbhbpA+4oJdM12Lu9vNX32HY4Lo9
dCntm0/aKHNeKiIAqes3jHQLamJw+gi3+rB9kVAwmSmU1HCgDrTl3pTHuBkRCEY3
L6+aOP1v5o5kNE0Xx5cis0jTsZTagqRprZ5q/zMBbV0ME1T/Cxncgj+bMhPlLrXG
ozFNkyYsDKfF3ok/rkyUXoGtaeCfkWBDb3IwrLKtcQH38OLPtpw4dj4cn2EwLHZ8
qbFJ4egFZAoi6Wv1/Z5u6sxljy0ot6mkcvCK3LSebMp6e3SAxL5m/8xRrbNib3Fb
ebQAXQxEen6NXLP3Wk7qwCG93olbDYTPTFg0GEjxVobruO7OOKsDRT8VWIbj127f
bWoUBB1B6sdua/CaWey2eHZ2Vi0Sa1Smz+XOGpodIHik15KWx33JhgkI4f/J+OiW
Va8+fG77jl/2vNSkTe2VEeOwILGCqKdjfusgKvuwtkhNH7/uTvW691mpl1OR8QIu
J/ot+TV2kB9IkkMjwxPIQ/9gmaxcflPjnwnVENN7kgc60BxaByefPDEcokPCILK4
1ofGV8H2QroLhP+ii+nt6TKo2mSKEsq11Xy354achVeyQv1i2Yb8s56pN9uqCdhX
9IMr+B6JHjGuj0N8kfq5mfoB5SCEZJWBoUuy89wSbURjvosGdCgi+cRH5W0chFMW
rYro1oTt5b0N3slubumkxTcucoB5w7XFmLUtsNdMW1Wt+R1One12n6kpICpQeCfT
M8xtkj+8tBm/yTUonnG1j9p0DDY9dxpP4V6/tboCXArY62PFqIBi6lVwlyY37D/B
ZER7NvSssK2umaRd4ve2is9cogBu/KbbBmr5d6CdSpS28MR6SdBr4j2p7MvIjmno
I0uSE1osK3WLofPriyMMHVi4Ovp8bb7DfcSx4teXY7GxG9YwehTqRDZatrUnZaP3
lGn6/9GtYCniYAID0xyKY2GoArR1UzMmq8uPSl2r9cOqy2bVkr4Sk2jiH/EnlZ9l
SwnrHdaWPSxzF8f8I6Jb9EiOiQTpSUlOB1yUV9BcVvvh/GXEIXERgjr43bSmV8rr
g6Xr1G31CJEh2vt3+4lo6qoJg9Y5BwmeM+qz+t9YMWuUP94PrjXxPHrZFVF+N3ZJ
X0YQ/mX0vvCHpgJtBhiD1BSkRCmLbduiZ+nFG2snECRnH++FNK3qvF9XGAxRqWgO
x7rtGQ85yrz3PtQ7ulRbCZ6GKgjIAsHrRrI5XkTCVWM7K8j3nYWDLt0JkSmAGRYU
IEgndGhd42lJ7iMxdljLOnzM8MaceABVyfLxzBTMBJdae/vwxdPM1LMw/uKx9TXE
TVcpUlbZNU747uWIRttKa2ZHAU8PZB7XbZhoiA6kb87um4kPKeGI8oUGFC0sfFgb
CMtMNrBF7MRMNsLTQEvAThhJnIHJoax9Juh1cfark/1Isi/1X3DOOxmPrGu/Kjig
chgszwM+cdNOuSfvA03fGoPqGjmdyP/QFyLIWSFdoVNT470v0kZAHfQxAX+8ink3
btRf7Uxb1dF/rkiwWpDs6a9SuCZiZ/GQ9mZjfpB9QLr+lSbvDJZDeMg85V5AMC8w
hGhvWPCaWdCvzjx66P4zWSOUclGfzUfHFFBa9MYx2xWigea3yuL9d0JzI4utYh5P
1HiNFovzwRhCHRhh0ujqSeE+OCGghrAbFjmZwJgU6mr68uZn0ogCbTtpou+SbhgP
xFEliO5BoyvKKae+07QD9SkszrhuwGtWWMYEQrRb/+1UZU3IzsnfruhHi0L1t4l6
0oyfQYVY8IGYQhi04fhY3kggW8pRrq+/CdZXayzJNjWt8nLtFcUYqEUxC2kZOHes
9QAEMdE3thPKeM2bx88ZiJQa2BxOcSs/v81oqlysFTTE4jHVttId/C89BhXP1fnb
ZQbw8OKt6gHzeHB/4ga1IBwoXFPXMA/X/vOJe88WlhVUN/Dbjvzlka4oNDs55N04
JVBPdK6nJxb3yAW6fOtXrGlQA0Vzjh4SCCbr4NN4n6W6SAdeGnbFw1OcR7qfVKT8
vwYF2+FWsF7Oq5FA9wswuFYGe8C+FAZRv7hmE8AJylC5LgG4lxgWqa/t4Msx1fdw
2DVIVHOz7HvFwRuplJv02qUOX8zgEGuLP5LssvvuYh3QLL9yrW9ZzBk7hTM9qbCA
q6Tk2vXhXSaSvy6cT4C4vXCZpMIazXsH2VZE39evIWosVqWHDufShqGTeDT060Aq
LV+A3sGW3iGSiGEfp1Jfr1O72dc+LWjq3HSePNAJUxeOHavzXi98KVw5nb6PWgXU
2atNJP+oVwfaVvm1uIJfN4/KvVnjKxo0wkJv4OQcp9CUoLxY/tsVl07ryrYJEO7O
ovhSckDw4/5O8F6GtunpLO2tfw89xdiHptzWlDsOWW8ZTOug70NPw6yyTRX6/T5j
uBK79DrkLcB5mTVaogwJ4LD7jFnbL/38Bcd7X5EPqgOa5Arwk5r6BwwWs27z5fZR
HamMYzf0aNBj/Fqm3j1JJSZxyzZGegepxjMTNpN78fPOBZL1daSNuhwrRdGXX6hz
n1r2E9qDi5V8tX4FYIDC6+QxpfLoxgvzXKq4GwqYWYuqywNqNbW4lRm855bKlRPT
wRUbZ0azdVlAuBbe5UWDD/zBtNhD8Rf81MLFNUTbP+/1E7TCLL314rcC5emwAfBg
YAcJ0R7Wat++lU7PexgIZR0KQdlUBjSnUGKofFs8UQlmb1HFWqEwj7p3xnnIEysI
l1/tAbCHkJ0pkVEFhwj7RMO8H+Rt9i9B+6lCin69WqAZPlYkX+q/BhehTVjHrTOA
k3Na/V3gJx5C99admk/O7nJKvyKR5DPwlPL78iOcqtYgvJ9WTyjhQmEnZK6I1C0B
iVvfEtTN6cOqzYrFWEilgYKqTqTuNCB5+Qcw4iZp6nouv+vgWv7Ikewr12uaTftE
zE05k4eAzAZZagkVH9FVnJikISWI74G9+CCEIoI/UXjRKp4qEgeHT4G8VrRc6fzh
vS+JRKE9rdcL8IZ/sPfcd3M3mkeYpLl3TzVdJC630VzMRgM+EUt7qTtAvbYXJfjs
Hp+NRwHX2xLPHKSsoWs+4IHz5QCgXS7nZ84XhLDrPVeJsqRBzPv6XanGEEpU99CM
sHixB5jHgsEPnnEDjZAKyO3+5vIFpQnV9manmMLpT1ZH9+Yf4iAL6ssgB3tFFQZL
mwRxf/KZK2kn8/P6fO3E+v6mS5SMLhtOlNq2rXjQ3eJojgmPjoseX1YGPJyDj9Dp
VowR8ZIZA96CxJYC6XVl1BS8fbTydQchuYUeUBuny8t73VrHpABCaUdgDqrlvY9v
EyP7SyqD3uBaBifZHRnKziv1n+1ji8fh+y+K4PfCiDLO/5a/FS2GmXAhn1NPYG6G
0o/sRiCZCNGcemKINh5UMolH9AMVBReNinK/TEiyf7gpjOUrrfP0WoN7WXH990m1
OgCQc7H4ts26fplxpGrYx3XSdE3vixWYcBhQ4zMYdGsa3rkEOPUMeFIHvuXPHJIA
hqNQ2kk4f5p35WmLqv3pOlS/+Xxz6RG0tR5gNXzFxuFok+qwkoOKc9qyB4C4UTtw
xh3NmvBF2YxExDM8BzmLNlyar9fDHES5cZVxXQIQXxQZ+rReDcK9H6Pt5lzU5GSA
cAqObY3MS0vbt2u4gfTYPLXWKa4w3YH5Q3Ql2ZtJaxKka4LNAEvuAwA8jlWAiPFg
SwwzTJvWTSPWO/ayaKkvh8X2ZFQkF4Xt+JKPNX0fwLOj0+qL6Pnrrpp5zzPuGzF9
1Ed/uSOH2VM+20KwhbRtcEMFvF4TabxyW2pDpNlbKGfmqt03V/TL7FOcQlROlBHJ
XL5z3Al2H8KHc20aKrY+6U89qC92fupnRmpMPN1rkbvKy5Px/o3wua0tyqQGpJYy
LbEQQAUG9m/yj/JY4ON7/GGXZnJ1C7JLsEfW8QeENfwOWw33j4j/PeEidpQHl6Fr
Jpw2rk1m26iqrgVYySsrLAVLrBgrZFFQ+4pzx1Aj0voEVCwD9skRfzM7a+7IRAxJ
pOamoUnPIa9ZZc8UJPR0HJSUbGNJlpAiKfGmjpYH1V0n9hIp5pruG8YhWczziKgB
+smmam99viuH7hPOlddg7TM7ng1wAIw/V6BT8pMsXh1+K4mTlc1g8PNJQIPT9MQs
b4vNjRbrWpiWDtx08U1aVtvjOau4SvCn0NQ6aiqA5lUlkK3z3AQuel3nTPVRJxdE
Uo559fph84bB/lG5wpLu4HJOHj6iXZ0aD+mOHMblYijm1X3nLbiuwV0iTF2smmiA
ndAVjcq36/oO/EWrok2R0NknZgf9QP5zQtbqVAYHbu3FBHnMrLB7EQ1eH+FmmjUy
Qg37zi7MCkrIJikxaFVUw60od9ITijfMrzUTomGp5FrTBxsINJxNcpGPsldzd508
7wUD//eyT8VM9Hv/Pz72FJfGxSzGk5GU5GzHLzZM3M1xgjcJO0Ajrf9+Yv24kivB
9Cwbo1v5IOUj42iUhIRvTwbnmUYRZX0j6xFXE8XrC6LvNiZNNONBH322d5Hq0/v1
6pfI3jRZuRWj3EhjD7OeXfXCEOHrcJzi/bDr+8GeUmyf05qwgpghHYM1JLy0Izdv
eami7Lku/cwwkvvH81yj5yKdqNLYyoII4ppGB6ST5VkYS0emafC/BkrBBKTlCpFH
rXK/byQPVosRK3rlSgSBFhq223GzM3FofvWmovzE79OqnGifFSV6pXW3FvMPnUKk
CWkPY5uJ6bhSLHTmX4KdOhxsVEOROLJLdv8gp5+e7x+7rxNqVd4ZV5P43EQwcg44
sYljjTIl/5NeQWWPkgO/HLjNT+TBW0oHnO9jD60ewPKjJUy89z7uy/FcQxSD9S3O
oOvV9LkcH/ptJr7KzSp8KWOicSUPuQy/1nJjh5AlAAJ4xW5PNlX3Yih1Vg6+IjBP
UzpAkvTz3+xNQLr3kIf01pl+6wDRDlbz1143ELeDYfBLNrMyYe1a6homw/YPHjhb
TYjyftI+qeTLQuQMBx9wdhUSDyA5/WWPMWR87CGdR63sONVlS2EiTdwzQBabcHLO
6c8wVXOydvnsa4wrH8x8TT8N2xJc4AgD9GfTdAdFbE8VznIJc5TkaKUgESh/IZ6i
u/QDQ9cOPw6V5PBEXM3ysOayWDCWIeADOxNSvt1RriLntNK4jXokXwS8OyrC6Z9a
Hf7+FAI1AH3T5afgB3ch9oF/CFKbZMA55mrvep/xN4Be6dQLL68Fw/nTdXDXDwjk
OVsaTntG9ybWy3WufMSDVnw9zegQTBV6OFZ2Mg16/FtGNWNYTOiTVNC6/3wVectY
nkdK4OdZi+jI2OgrcNfLwLk6s19ba+cOTGTzJYHSYYGzd+8MIhyST5JcCYhv4gnb
Pkn4itVv+1bj87We5nznH+ae/7s23k1f5Y75KVv7kTJOjm9+ohNtUynBRa/lXcu9
/Gm6VFVC1zVdVU9j3TaKEGqChqn3dybxY7GvMigc2THQ6vCK11XRCgELvxh7YQJZ
H5c2c9mUXiUkVEVrwLkhLSB7NqTPtDOzpIuL60Uy4VxZJVG+aEXW3MdFEzh2SlRv
HdfMSm0dhSa9iin/ewn1+QRYBLzRSDeoa0MFO2XJA7Ui0EuDHqBQfRCUh7TYduxF
6n/ArUdFjfYKK4uUzoRvOEsdD6utV+Dm/an19AAcXfVJWnCJBNQiwrv42eAomze5
73bw1J3c8ohllaJXbjpUfoN5Um/a/MyUrDDzpTkUct8vJw8iPgVf9xdNM4+T8wi+
GSPME6MKnSlxbLYj+IiCIDfLdjhz0qV+UowoDQ/UkWnwCYmVTRLBPL85RSuUJTTF
XVL+ORwtPXZqxMim1UmdfXFPjmPYSAr3SObSbh4iYG3iPvccz07chFDWMJBCGxMx
jw0x7AsO3O33N2bsfVqr2yWV2hGGIjDzkmwTxd6aDg6viokNZwVrBMLQztTxU3oz
at8hrrBEBrifSbPnwriiRa6KKHaE0nZVOjIZDSp4ZI0uclunYJ+MguZmixYBBxo+
6s2j0o+QIGMEvhD4+/bBlWCO0n7d4eOidVgaAS3fCdnF+mP1lGpxgpBakMFfT+G3
+ITGIE2+NvwRUEHoqUJydQ/Ve/aPSvay0FCeeeJeuvDnJ3yTMr7RgtBoeJHAZevv
qzGNxpDiaIG1JS0psrJ8CpWZK3s0FfbRMNyAxk6eosAeHvFbY5/80RML8uOnrnCS
ve7IBAPqFdxfRo+6NP/irgsIVe8sqYVEpQuKvH3cxgIMneV2XDJo66xowChS2uN0
b3qyIq925LQ1XcEPSe+SFw6uRuapvfrCQLvEBaitSqmnSSwIlcmsGw07bg+WU0K8
cPHew6+5OnVSPKB5H0dNOzI31nui2Tsp2h7R2cWk2FGskRHk2s8IIRD/n+3FhVnz
AB59hlUYvPtKyVCdWYW1+Q8JICgsbJ38ZuPKql2ELD/H5Mfj/B1P6PBjDtmwjBo+
ICYQBSUx6OVD7Gch/au3mB+G+OT506a3UkE4H/1doW1Cb4TM7gBGb89Yhb4LiOSC
c2u9k/Po/LZZDVlYDkouJv3+9OyBBfPR6oNfu3LjiEUBQmpuQ4owr4MthZnNxlsp
bu32i8sEDe0Gdtrr32iiWLw2P9LJA+ESTkXgSVdyAh6RVvSEVV7FJRwhN0zP8ten
UKNwaIQyX5H/bEeqlacgr5xZ/ivT5DFG9rneM8bl3pLYg3UjfHdNTI0fCLoehIQo
1bW9dF/L2Lmz0XsRPF4renZGLL1paHSVjDC4nmzRb7pLiD4FsfT6BlPBWXMggpzX
QDWHWNN7LD0t4ZE7cDkXEYq7yvg7xxGUEbLO3KgtIFS8Khno34zg9oiMRCtdJLSY
p4PQorjNM6Pr/GZTiGR5Apn50rIgNaksxjXywYKI/wS4qVHxeWTDwlFByKYDJL9M
3gPB6txHxpxvQ+JT4SwSYY1TSuFyH97eDaZyWmmYMfvDhaQaMFgaRjUK1d2zazuq
qoQg+jjRtSKajtIiXvgfcwCqK9Db1NHkQz6xIT3zj0U2iliAX3ZI44L+nMzleQug
uywLNOg0ecfslsTeUi1+oXeAdNCXHDzWwB5qzb8VdI1vsWAdhjEVrjMHnqlLk4qt
qtKIpLvJY11v1tsss0NaDivF6WdQ/QqucXI0oop6/1okmajukkF9y2Ub7S9La05L
63vwnEugXP8Zuin8ZIMAueWe95fUhfrLUsJRp94+Yo7s2Wgth0WAQVIsmXYQ8RU9
7BsF6P+zPCZsuzdqJj7QJqcUu3PI9YKxYl5R1HnWPYHKjDejcuJL89xX8Ru4fWmk
RmBwfdqEAGJpRIXdtGn2vGSrZ/TfeN1mHq8Gth1aX/32HZEJY3sw9gIh526FN2kQ
Bnbo5p/gYRwi1/1vMw2aTxfe1/KDskLgBwtksrqWB6MpA+AeUhJcuxuAvVQQ4Aa7
3kQnGTpQ7lM+KzfPbWsWtRUSxX9OCIP9jJ5dOjVa87707S1d/Z0hjzRpg9KWVyvf
hWf2Oe/OHumXMwa7cFsqvitK0PtNWJwY06rSALYpcdjO6DT0svqB4Fy1VqQfJQrZ
4MP67H20oVrS93RrPELUxXGzOtoqxGg/tlw7Fr3g2zzh9oLq6JLqMZYQfAJBuGaO
fPw9FdOVF4kwaloEKMh7O8zhwcOx0kbfwREeMo68n6h8ukaWv2DCweUaW9SS1qr6
FhCAkltNrPopCipeyJtk+rX2FtCJ8jUZyFKGvsyhCg4ofPG4lnKBkzOYWZDWXrIX
DsTdN0kURg6LM1ocWz11A5DpP0eXgmBBVr55VNVdJqO7GJJF56Z45xBfBbNDWqd+
nk54yZyLSixvw/tEoRZu1JZb7M0EtswzP8dBTRnxLzHzEc+BtLYY5Cf/YQ5IAS4P
a0CExTWcnePBijUdndhDsTbWOEVwpUVd2HU6pwvFQ02+m8MJOqPvWs1qrPOsZDUn
KYwVofBLBE16/saB/O/aejDOuJFCyDvQIzNCNkOs1esbiAhjoJ76Ft33x5AbhvEm
UyLjnGe3ov6SmtFuutvECf8/sZPUfd43ssuG6t3ZmHthagBj/TRZgwsndcjtkAR9
0zBpJ/ciLhDxLuHnMqw/Bj4ySFCacE+hT2lg6QYHl4VwrsaTppICUt0DJmZfJwx4
mwtNxdlPp71zXmSJnw0diFO0n1RyM+16IBwDj7Pe3+EKDvFb4nK4DWA7wQaoQhIU
HoEv6Bcn6Nx/9XrrbltSE+Gi2Ub9oqhnJgxZuBG8P+5/T5ZUgploUoxx+8aQIcSJ
IKskhwWyigojy8A24kuIP434y7iZ5yLHYxt0SilrsSqbOIUEt1jJcBREhf657Bup
vksiH2DrWdz1u5SkpJrB5OE+Bdmj3GGRe1BV6GFWDvAKtk4byMpqpiloyMyakhrK
Cg2VpexMo+fo2Vq8xzU/+cryZ7lpgcB5Q+DjpUxzkK3ivsJ2Q36zkxHIhZloT5ef
KJLMhOr2mUrZI/nG+hy9U64VVxMZC2ahTgnRLjBvdR2rOt8MMUrkiUoZTkbNKIHK
9c+ShdKjkrhriBLZ2LMEiEssQ11VntMmyK7CiaVg5xz3uxLaH36ReIByVUf59nKg
ce8n6i+4pHLo+ZBTu+bbeDNJHZY5s5mZUtSfFDkPu19v5jBLR4BJwzf6u2HxXkwT
RnwkyHJ/RlIsXqC7cJE+62EiPEM/6/vGW1h70adhauRzeEUM5KEygcNq2KQ/q8dJ
N8VAaln8W5Hxx7EX5B54NlJGwyHYz8BXC98LdxMU3dHcsTzzncnhzh/ULoRCI33R
cRWM02/MkQ1u1QzHBM5yTnzP4bsLZsR/8Ez6BcGwxC2sFNvk+qiqrhtU6FDfzERZ
PsYkM23/OPT5dTZDK8a7PgqVZpcotCyx3wPbM3OuhtDRDfgeC54IxsuHQ53KrpzK
T9WJ6BRck+WerrV3jYj/2vQA5nz6sDOunqKofTyk/CQOFWowN23Q3W4MLN85EnMn
hOA8f/6lSc6M1DdtCIHwPjq5vwWF0nYSiwA+E3FU6Gz0gYy7lhZNKb5voy3sEpph
B4COccFN2sOnqq/dtpFLkpMRx5lZdXr2/juYwozIau909UWutLaG7+OdGf1BQWtS
eIFHDW+xn7OZc667aB3UBpS61oyhsMqgmrP0AhefH7YuDXvbSMPfQBe5+Z3bhMZd
WMFYh9iwtOqrr0aT5ZgCxy1DopFHtqMiEEmI5sqjgYkKyOnzitULVNKfXd3kgvyI
lVy+sJHDGq9bMPTAp+0YBcMOWUGF8pZ+bQ7j6ZpZb+uIxbTQ6x+VDskaTm+51Ilx
zaV6Ec6XlNu9b/oMDBe3dviFR9MxbalwOQhMADcX17O6O5YrwtJABnz9NIb4QLrE
9iqs4ZMwk8vk4TvxCyZ53dOvIGyD/lT/VlkZEXzVg+wFe6OQMZxT29RrS/+/5l80
yyCohIqNt3XB+uQf4B6M2cAI6/XkCChIVkaKb0GEBDjOajtY0BJrA6KGRJs7m8BZ
xc4ur+e79lLxXYCJYpCGVb0ocMnTJsQO+rkdryweDqqGj5jpVQclRfyR47mNNwAL
moVlE90hCHJVOxLJL6rqUdZPGT5afmRafs7mkKA7sVNwTgwPH+FfOmvaQDmZjd6G
Mn+czFQwnOWXJyNp5Rjs18ChlCQmrlWmHItcd9yZUdod7kbdZ97/MMRCXUk3WQth
zQr/o0rlpEjEib6jXdMpzp2ainihSo0Acgo0VxwGq1q7aChA578rVcn9ZQLrXTDu
w28+5Mw6vUeBVm8VZQUQOe4YngVYWjr8qkjePd8RHjk5pzc1j2SxL90I6iDGr8eH
pAiydWwg2aEbF/je3B95qxNDJndD//EdZT/cXfcanBFSMG6DrgiXpwgTNLHkgp46
p5N57UYBIAGtx9gpXkZ8uzSqOg9RSjSqrA9UZQZ+in1/9wfV6xAmlo8v+M+MweU7
jFyApjKOFLYNIXds7+6fOsmG3TfA/EjFk2itvpMt/k01ay5V8SF3gRO1Xgp36OD0
tgXWyC+K8KaQZUAwMPQCyK5pH7ZQFRKMts0wNlyAw3kylCtGWAzXqr8WLfJ05RLg
yGGI4n/p5CmzMe4/E/ZMdNnMQYr+Qj28s6EnTaH9PnxY4OeKkETQf+V7b8EoLh3j
V4LIa3flMuMl6DvlG74XlOBIFm6agTbXdJJ3tduo/tBx6pVPfFCnlkheIq2MiKDk
bbdPZPPyq/jGwfeUJ95j7owNyauy9B2pVjDtkX09723DEMoJBqs9YjxJZeNdCtUO
r9Ocd4VZKyCl25B9ZxWzwKkftcNNG7QpDobF4133ZJxU7cy32wxCgF7DPUIC8sr9
CVhvon5am4lzM6frrW/6rc72rDOb4IuQKuCPKGkxi1U44HRpgonmrhjE9bzWiwlB
bDQL89BjEmijZXBtGNoplzCug7mD8QVGrR/NWWVx1KBN3/GPUr1ykLyuFqc9yIPq
Lm1nI/XJfXklCWpCSAu+1RlyNKx4a7E78fqSLapp+Jclj5yYJ5Bs3vTPzaxQKQe5
y8n8tvTnTT5xB3tOwwjzREfm3erib3FjLCLipjj6DBcMT0r1IyV7PxaBYEJF6OcF
s+3VMBR5hqXOcU5FYKM9ZyatjFSBD2agcC/nDJEXTYTvI9VSIUaYLqfxngMtatMN
Xa8XDZjGwPEfHSw0hMGR5xnpdLnV2p7FUcnMMofExu0qBsJqnw8Jq46ZvTNXAeqk
EzuMqLzutgpHPFlGTbM1KnzMtLEgQxw+pRsOdzq+WyCbc3X2JYM6I+YPzTHtiq58
v709otkTkpPUh/1FzHIj7eojcvxT8qND9Zk9QJxZ4KlA3EgktznJrn3i9Z5IPFQz
ss5HuaQPgAYqMxx68Vbwj50F2lMchH3xts6kYRNoypREaTq62R+TwU0sASDAQWeB
ihRvqvv3cMIbUqgxz1L5B17EbsVggiOC3+kiBFxB0OwzXzq4Jw7BAeUQ7jMaH4VZ
LfrGxyqazuwKLRLSF8nqvxtxUHV9ElveRVqmP6LYo/Uc7FEuDVcaGJABJMFckVwp
buxrgLiD0jEHYcUcK6xojZWyPzcwXCafQURz4gUk+wNKds1qFHHAHrenwHe3gNYk
XL3wkYGwK85yFgrc0kA5stllJu5Z2XuHuOPvpppadM+fhzuqyv7Bu7qyRKmOyL5M
N+S+Rf1bzyyeKXkXlqKT3FHkby+MgPQXHivY2iPwOkScB6CNmevx0cCA89HeC1TD
tNtJ686ZZLTPkVBjjvTYyPE5h2PRpKEifCV8DM1HNZpr8TV3ch06um/Uhdn+SVXy
d9FMWhTFBG/0BnPjiDy+TBr5XiymwEFn6j26wmhsHeLQFxOIQIafqbV79H08AHx2
ZTejo7fPCvwFtwDAPP8QOeqEUqB1x4BQrzlcN6n13NMUwtfxthmV2sevlwDQvUw5
AlXAkW3jH7HXgt/4SnczLHa5b9/8i4n3nF/kUoUkjMni5VWIYIqH6f2qDM84AIZk
Yw51NULKt2ol0EzN5RYZ5SZ5RASyvNxj29S3vPKW2GMlm77cJmqsysHC0ZlwJLrD
8DT+UxlHw4fucoif1hp85TR0A3WOHpxm7pIIJWTNs3AXptLvqnJtYqJpyOaINyZF
AY9qVqUjy56iju+5y1SFNCTbSMm2ZMFaEs1bY4lBU1d7WCClV01qlexTFU2OZNzH
XUFaPI/PURmCYpJvRtp8iT6as3PLAXoNUbqG/921kg8DWEN8BOGzJIS8HuKmxDrJ
Zp9Wc8iAVfBDcfZ3f9ZwFVtdKJAUZKZevgL4BJoPjkpUtCyyuUA7SUwhTxTRAUx/
zo+4FGw3jcurkhs/agFHmvgXt+hZMsezFRDUfm0iegrlM6Vf327H4BSXXEGDz5Gu
qGbtkcZ9kUDiE7Jzwc28cV0S9FpbstMpyCkUoHb6nHTdq/GY1jAlrtseDuN6pmyw
tubV6jAAClTVUHHLnOBRZ+tPaj/uxWi45Ak2sq1Ja5XDGmvwu+uSR8A6/xeCEnlV
Y5I7NTS0jk8fSVlgPrZG0CK9UfJP8rRG5u0Db66ool1pFzrfN7lV2OCaom4G65Xm
UBhQ4fn7TLlG13A+Eg3yvQN4Q0FbOUOAEo6R2hofXKKA3qIjJJdvoDHiRjlzCaqj
GOaaCBN/O6Ay61OQ+uVDH3WP1Q8uo6weKB3mBofpz7+dwuUILAGHKZnG369oGMbs
600RB4bDz0QE/9btiw1U0QcEpbmeqLQdocgK69JTCPzJWwzwctkGuLR7Q90BGgw1
d9TCvxq+m84YBK0JKqCOHEWS5NgC6ON6exAOu+9BX6O1jx9RVcgcjI74akV7B8dd
WsDc+vmZAQaQ1u577EfcljKjElvgwI49oTxjAkEN+akVz4EzKanQp00/omKmH59F
r27rO51ouBHxmCRWJoQF7fdnLnZq3+eZBGsbV3uUK4Yi2Ur+R0t1PxZIJCTbzXDF
CNcknO/qKjw/6CgIFkBM8Wg0TdR49cWM0JJRH1nkvQcDDxmFmO0vmxkSo1qF+tVb
pqeG5KMclKU6UQ7VsVak7XGIUvGenTo0DLrBzOwMeen87UppBR/W2vA/Xm4sRqWQ
li1df/rDx2sh56WIf+LznN54WG7vZXCPhRYiMET7VVeEyZ79FtlR5Dd0aXKi20Px
DXfux68e4y/HaxqGqQYBKWvrAXBJgyMOwT4lF3jEozn8dVssk1rdixWNijgE7v1W
2ufAkro16Wb9wOCtCUdieEZVBKeoGjHna28AbWBXTFq0FYfbtNXsdkJBGzoOfjZm
ZgkWS4V/qR8zPWB2oMbZHMI4yNNbjs6fSdCsK1zBgblwD/syZv8eRtsPYme+uluc
FyLHEm5IvRTBr6YB3hvyXgQuDDopNvYRBHZVz2Qe+M3a0oAjolnACM4dBM0tILWz
7DJtHQEweGJw7HSGzd62WJWhFho0a8Jyt+oMZ8OE8wJoi/ygJg1zz/4lWm+Rm2/t
2zSsrrggRzgB/k99Ewuv+nBbH/CDAHyCPB9LQXozObEKL5lbAf3dOFYHi/xWNTQ6
4YPuf3JS0cbYzjibp90stEjDcl1SzTx/x7JmvcpI2kCI+F22xt/FM0nh/BDBMbzg
R6SIB5zqx93+YgOJ29u9RGUKKB49LUgcFjZsXd2bLDmP1RU2x383ZfZ070GSkG6O
ddwwA53BHSMRmK2XkkiwWFkeH/eUQek+CeqxiHFLkR14xNO77moNt8/Tfqeb9e0g
93Rsv6ZOtIUo1O6xmyZ4GwP3Op6eNSLVIAsgi5C6+rttADbQlMwYOYBNtUu6FcRF
buq5fyz2Hk6VCE5Uijl4hLpsTRPqpOXYKhHREVlCTnjsjS3pjlRNozfuN11RFAZ+
WngPflfJ0ues+r2viBMDh8pqlvlolHQHIQUuhQknbS61HNqSrejZz7FoulSEljoA
eIgpBg+w0H2xgZo8k6FmCFB0oy/hnb8nKn/Pr2K4VDsYgM3W+mumEk1ZWH3rjkSb
8lkLfAZlG907TRS9NfpsKcm6mxytm0zlx78JK91Uo4zr4TYxkOek45+80WD+MW7j
bNjKZfB+poTPlpYwOuLucusk9UUx1na7nHOLvfxHUfu7pT5X14PLZK9wOIKEamh+
sM7KFaYX3xhQ1bciiCnBQa2ljqg8Cp5FM7t7/NDDDSncWjYHIGi32zDF5HZMe24j
KxbYVX0vt5AcAVZnpBiLpRuMA/Ho15re7Bxam7MWrEd887rylKgiDxiVZqablSWl
vDVrf2og6PWaLobuHi96D2ebT+ll54sZ3Ui16hs1A3bqoXF+yH5eVydEOMjLjpEy
r0O5K9vo/TYjIRrsrvG7E16ENJ815X4BO4qiKmqnprWQlCmdZmaazVwmueO30nDr
CGiOabAifQaSUTskaWo5UKNS5zTZ3tUm7045eolKLHy7dIqTM42crUPeg+iB6SI3
XAJ9jrOFUGwz5IprBwCFU/kpQyWqndxohmPNlWrOf2N/WdcYassfdFMp+LKQPDPd
lBwnjlNrSGZeYFAfrt/8MV/T9RfXctQXDp1KVt+uzLo9uw15BRdFWOLAF18uOQx9
IghCqcTxTF977td6l0ku2xK6Nqx90LUHdu4VJh/aJauAwcHTD0nEkOgHCZTH49KB
8lx9q07s1WPGA/N2wZo415Hfvx14mDmHkYqeM+OidIFRqmgpNvZ4eHKmUUPLDhry
7gCoKStGgZ7p35CpXzQ3jp4DtEJt3Q1hCJX3gYJvQZsm87cLNfP83fpEuOZ2qhNr
sB3G/TwT27RKHg4OecsqK5OvhA6UA4qTcJfl9za3nrYhNx/OTFOtMAq3+jVrEmUi
DwwjaaivKjy9eHIzkmOwrzfDgQYdkLc2t4F7bcYiOe+cL9JQCEbDcU1z0dmKK6h/
N++AkTEcAZxG+9awTVZY0ULFhpiZ0XddLYptF5SqEUAXfoqCPy3512DRnG7iEj0p
rBPig5gGTofVSG2gZHDOF+3FAwBoPkq9yMwDTJeb93FzqR+fGgBmGDHiL/HTlP/E
m+zdf7VBhbqIYTkXpMP34CdB2KdmGmOJA8nbRtxw6zua/Inv9zGzwwjAiMEs08ww
2Uhcz6mlIBuAJdu82mGd+xwVj6ZDPa0u1bIblevVEtGCMf4BxONp9CXpVnw7jaaH
ca81d4OcLH7mWiSFl0ZQzMIql92YlIbe1Nxz4ltuWgRV4EjdO9m+V/SFpZM25aXJ
qFpt4fP4Ef76Wd/8pF+/UhrR6L3BxsHMlnm9NTngsWgzRYi5YuBufbWK9kePwT+m
uIEsACIffcTgfaGw5xGpRowdexZma4AAQLfFInaO+nLDFtKFOFQU+ISg9DMA1D3w
d+Mt8FXTP/q8EsfwKv3kNzFSh2OuYiWSrKjzktvCrMUjOMC4IeVdnL0RMBQqoNrc
kqXFwPixow7wIZJTmddq5tYh/egv5Esb7tc4Qj4qVpwHkMGNbHNUeXt0tnN3KhQE
WJnV9gDIoCBDse9TPthhez3EAMvWK1l1iz4MO04/MHValbA3Tng3la/ZCswIfrcg
wsixgUdCnIzRVyfU3HhPkb9K0xuYiMe16K0rGd9nWgB8s4rQ1sYOnzcmSuxW24kv
Q1T0/23GRWgmnF3TSlPjS265UFx0yQth+4D/oqEiGf6n+wQhPdxDDjOE98wejPk7
0EOGucxIdGteutkc0Y84zRyfJelrB61iEdp7z6lYlPaTwwDt1r6XNR5DhvvVygb3
pRvZ3A78/mVLySP5/K8l6d+k4wIXiCGr/hnMQEXFcMrZQO48Kh0QVzF0udkqsdBM
07DZRvjjwv6dWw62ySP49PK5ngI8NcbgZFW8iiJudWHkHdzlUl/K3V2HbYfR/zxA
yAxBK7m2NlrNcU4TnrbO4Nh7YKZnBaRezEni/1TA3MpLeYGCPHxyHnkzTpOWnnIw
Wd7WCXx9qCshUSwTT1qh5jbZKt4mgyLmhFhlJIU/a4UlWxzs54Gu4xJSar9ONlEc
Dewe7/FZSF3vycTGG04TiZgeZBim5jZdl8gcVVV0rKcg6ONLQOFi/5cB8UBh5lPo
81gI1bdL1HogUdZz4FOrsZ+5BJixDZ2GD1EpWxc+RDwM3jzY5oQ74qcO/agKrsqM
Ad1nsHgY68O0cNJwjdvXW+y3bGQKzs2WhwoJ8yHQ0dh8dhWjn/jiVmMGQtxeuPCo
BHiFHyx20sg/jQTw7IrQtoA6A26NnAc2/WaLUIu1LYBffGUhUDKeE7pssYFbvNBV
7U3++AFlodCboG/ImVnz4BXc52namqYjMq3XTO+ZUhofy5flfDELK5MYoHQ1tWid
kmiryYMIuqJkkMNucRq8AgOjJmXvYgx14VyVw0oShjkxXQ9woPeIxFgxGOuAGlWg
tUgSKwjWI86mxyeF5nOi+lDUXq2iqR+oJ3vM4J9lxq9tC7lKYZTlfn5SEYGwakGs
hcIPOD2Y62R7IuJs3dH41f1STh1I78glA2kDtc01pHFt3K8ogo2t5gADTQNh1aJ0
635lInzVefZQV5BmTeCZ/evtT+vC46SJ6SDxNUFaHN3IFQBmu0XhIHlQYRmGAg2v
p1I/3vMHSyhde2PcpaXLAaCgNWaXAcOvXHgVHSO1XsX5EHjrFA42iWDeAyuI6gpG
8aOQNbz24QAMdeSLxS7O+Yb3H7HTiIwFgtTuuz9qa6j29EQB0bGwl4j3jVZruiqr
Tyqv4uHokte/AZpcZ260THHQrpLo8TlzI9U+6rJeCLP7CgC1jaUvVN9XeTYBBwaz
/tHpAaJGM97DREGTKrdPoM/xta7a76fJ9GVICsu766MZF6DOka3eX0cpwIKN3BXc
nuq8CcjPtRCzpZsPHvW9dYMwSuKPGGzH2hreVtBKKHI4KvCVTbnd5m7vlK96XT8W
kzSeyEucqeRxDlwN8XsWz4WRe9rybmK7zmxQadR5ovUXXwsc2khhbB9uGUsqmMK0
8rFpLGlB+uFzgFNC3yzsX1OExxgwfdh9qsdDwm2FuC9571+xGUnAwaksAHFiyzeM
An4ady+tUqI3RgYaLtUWynfZRiXwRokEPSOfKuRJKZm94qX2OfJT5U6h33vr8Gbl
iD+/jPyE+mTiT8dEdvzEMfRAUvDpardmG/x5x/YqzRzZRBftbMdiRNm0batj+i+a
9GmQDOdCC4D1HnjwOoIqfdYSTvCcUCDoYruJ8NSl2dBW44IgqdskJEVnCHOyDOqV
QfAPDNKnZnG/CutpJ8emkW0DOREj+7qS6ue0aX8tUs/xo5KAXza9n90T5326mkq/
Gc0J3n15uFQlxBIuHUugKznXTl6LJJT5nBMvVXJBU23XPg8RmluDLhhpubUVGr0P
na+G25b7iz5HsY+xic1MsWS5O+1TnLN0YOUCP30qhwSBa89jRDFM7IwmTugJdq78
koh7d4/FzR+F/TcvQAKmZ9HwqgbcCfy5WD86hCYKmfHdc9uZjTPAD4SRqvj30vnX
Z241Iyu+9b7tBYKbuB7oKAFYoh7nRKdFQOBehUsJulKefC46WpAUt9pdrfJ884Z7
cAhFhLpXdlvGFIQkBR3X3KVbEgdh24lAyb6y/SBuUMri6fEpCQDpCwUjEYGJUX8T
QLnYDj1bzh6ok1b/vyB4P49OlHRHbUjJhHeuvYCg79dsTKSKyyMpueoTGrkERU+f
9aOtSIclOWzLWgdbC7dQbiIHwuPzOEdNQknKiGwYv+5w75iGElhyd9twFRoxvnPg
NZ2cifnX+Tj6xO/mga6BANu8R+JYIpfUkA9/ScC/aNhDpMygnneIrFOJTQbigtZy
V7cgrpPsBOlcCb9OHbI6YKNMXLTSTgPpREUCCSYWnLUU3nTlLLMLrCDBcBqqRGN7
KCl9blbftrjp72gstwgnnFJ0RS5hjKHQBt626NpyxXU1e8u/71/V3z00fOouD5Dp
Ml3qnWtbnuhwfIlx8ibVhTGrz4tSq69FmKdf/gxYDA3rUowNrWG8+mwlZf4Bcyx7
jdD2G5ZXnxfDp3SEFjvKcZpIVR7syIstGbp6rttpxeq3Ckqj5/IdumdpoRH0mpZA
0ktaRvgtXMKBEqhBzqY2Qb5FfDao5NjeeaQN1IGf8STogF5MA69mGOD0Iy97GCgj
sT+7BJe5rf+i7nbEkZx7oq4Iuu/IkD1YXirM7lhvj2vC8ent+mKpa2VWHtShIjn1
/2iAZK2ssROno36D5Y35IMvRdcCwAKp51kxwtjudMiSj/+r2q8BjiC4jTb4guT0H
/xyP2XquIlBaRtD4iYe8WMbZGt+ZIR578IY4KnsZSE7Z9vDyJoyL6LVmg7gN80an
nqhbcud7JKseKI2EJgjgB5nF1Yfvy5ypKGK00aem2NTCfhLMCsJ4gJ8/1WYBMx0M
kv0hVsVDpKUWSx+SEJY+r+zgvoJQ9IcDeY903FB76uPHf5ZbesL0tj7EcZT2+hBx
IYWCT0cYGO2jhLnkLm+AChpTS4Uf9v5ovHDcjEOranfGPV0cv+Z9DOrqdVbk7LhO
e5ZLUXjl7kCV1QWkuQMt/1jfegND7KWopdpWHNzi3I3Wv6GanfYqIk8DhajoNkNk
NivFi1FgIg+9wguNRVdIlA8Cd9Sp6x/NwS/Kt0KYRYnvAx9F+VVxlKamAAP+qSDg
TFVnvTP+ZD72bhZoiJ5lrVg/6KsFgC4El3Krj+JZ0LD+LwqcI5FzeMJoGlwX4zHu
ze+GyYrJYe/tvpJO+KqmcPTwC4ZoF0B2OQJqZpKbCZN7sbtD0G5C88Ekrqo6O8xE
YEz220WjY2vw+h2bz0LZ8P+d0TVrXjqlN8N9sLsexgxiwme3epcqbs6SApNxGsG5
gW8VUr/TEQ2tvXdOOgsn8ym5KKbjG6k2UvvHg9kpfqaQ/h8X6QXJO/ddz4TjVYZn
J9jBN3EFHbhfx9p57PfqjrMZIsKjyzHb/xBwO505oFKf29lKVqXFJ4JPMQ0yF6+f
sTxORMAasawcEFjTgHjJlNlh3yTdi0YpgSwpBa3wgdDPcTuNLjAnoERzeFJE1w3X
S9Z+2+jLx/l1ADotk1+ERutfguS6HncKEOmSyskvBVbKSvuFb+OAGc01/r7ogCv5
ofOcHnWl0iMX/l7XVFBZDVBqLPBQI5Bu6Df+eUstLvULT5iZuzXThCYvoMXUG7E8
MsDIBIO/X3i7jEfVLt6Oq/TvjV2r5ZYJm2EzV6sKsfGjYpg+JwB3hMVzAQOv1lAr
HSb1yrhhYyILvNTYzxa072yxI86fZ9crZrGwBQilLzwMHBsOaA6eyFzlAne3Mj0f
8QvVWok+CFadvpV6pOqMCiPXKtkk/BhTRB3I8nLrpNETasAagpEHo49verCqLv1m
W8gsbu6NOJYZqOlxLIEJv8oYGH0cENnraHr25pbVsaIXebbT4641s/LN3+oQtwd0
p0kRx+8eBGXA8/4r6fubcn7WmbpZqoRM8PoJ4stiGPwD57siKijzUEfWpPKX1Vu8
DnMYOqJdNS+7LQUmQ9lwXzT7j/IUKyp5LqrXz/DXVVvAVZDmrnDpmgNrCOEkbFPE
9ha39zBPYwKBvUqI+Kj4Xen8GY+ALd0rJaNsTAcmHgS6wHts4eCM8i0bbGVgqPy3
dhFVNaOxCAdw3CUfMAV9LIl3+HAGHbyQt7PtEKKklh3G7QEJbF8nyVpl2Y+hv0ip
ItY7m4qVVP3X5feEFoqeA/ZcwtYFxKpf7cCXnms2NW22AvqMejND21LaB9hLR07a
DF1JpVKJiekR/FNXpSSDQQ5/ZjUO73xDjnCEfp1m5P2/1II5IcApZGyKtVbRFv0f
5JaWR+0XjffBhEtdYwWDGegonchwto1rJZyMUX1T8+U4haRc13WbJj7FRDb8uP9z
+wT9bLQoZetLBrCp+LZUXD3rrayvLcsiO0/NzS9uIGk4f8QAcnyYswC5yieBXPV/
KC2bK52+EOZL3RFURQloIKWWt+6om0g2q8nEvHWA++Z1HUbO6pVMV+2koQZhTZMb
C5fH5uS1j1kJYv9N2eM7IjpCu8Qwdctb5KEs2vFYMTd3UqhQLjRD7H/7BTuENP+F
9R7fLSxY1Kew26yRX+Ok0tlIXZKuAZe1haC69CO48VfqS+EM82y8rwppTqdVMVvw
WlZj64XPuuLIMfUiP8kdAkMkP1ojN+B2RH2NvrJaR4QAMlcIpy/GHc/tT+nQKPyl
5XhkGaDgaN0OVY8JjjWhQ+NmfJ/gb9+81paeJDoyh2zjUTZ/2bif0X4kvaA+TOnO
+2RWl4KxWGHs7cdv0W1+ibTGik4LVQX3PACNxA2peLp4g94hqZtRBZHkqSSfMsq+
42WFPDlerQafrbfiXP9k59nALfWs2IgmvJZ2IN7cjwkM+85IXpewDCCjE5yw5Svl
+l8wYTasvxhGhpAl0or3T0rZfeaSexNvJWDXjez15J1Ghh9NCyKGrfYHplOk6jYg
H/iIAhmVYbrnYXlHa6A2Hlwy2rhyULS6rvcyoS0i80rXpigoxelylhKS7JM5BcVb
DfTFDATYPpe9ZsW9L6eGQxKaiiAZBjN/rw60l0dp3iWK53nVN8EOrREDrfCsNmqu
uYiJDqUbIZUTuQlhOcvl5FvjkQF+xtBhQj4cZZALpZyRQpiSAiIR0jPVPtdLRO6N
s1aMqdQ+PTaUvJ96XMoPX8TVn37kJiVZ4JGh81/kiIF0Dk0FFkblwcKpyf0J9lmg
kQgcNAtvxVXg9Tg994NlPZDNIR09JHr/+flLZjJ7EZQh+8N5Q5B6q9rk3Of7/SdT
xwzdNTr+hePtIh9Y5vxJUD2HkFJMEkkWoAn0yYxqLRYPizal6iorT/pANan4eym5
6IZO4dXOeCAK0mpFS1SAUkAxsldu9+VV3nEG7spvqxKI2XGcM+erJ4Ix0+vfmIFK
qbzFVxlU7PJHc++5sGI5p/nNsv3ToqGZpN1ZWcoEQnWgBIKNQaEEj16VDVSYWqjl
CAzfimQSKcKAjPHM0BovgLxZCM01qt6zJ8CCMkpkZDAydTwht8ji7Ffx3bMPmbxt
2ydFICSQoW4lpVoqW2mWglimaAe5L4zY3pbBj6MNCMWNachCDbPTJv7cDjT/R4yc
LPtFLUidK6ofXW1Wf5R56NRRyrz9BDl/U85cUpDVBzkDiUeduWjLXiDQDSwJSVDA
LNO2WcvFT7RNIQawQUh0qqko3f1/oZUu3KH2vxvsO1SJ8sqjhRBeTcVtSrqdhujR
kmnDVKe/rtQTr7cYWPcPztz9gmi5oF6Y+d0ex/pdWzakohapwgcXUD2BJcGfWwsJ
RW4nnLmBJM77p83JnKMgBMe/1YqaB+hSv2RebNr5T+W/YVIV2roiFhGjktLSuxgh
WJTEOn5PREGu+O4yRRf6EbJF9CXj3F21eK76ct+idjtkRPuI5gG5B5aBu3kgyEXO
X9XsJBRn3RPl1FAnCIVB5lN48HAdF4xvRJj4SnhKdt+947n18roZqMTVFuAixPC6
l/h/woL2cYrg9OxQk+9IU7CeB5S5d/i3/URJwrt6saBAQvH+ieOmRxjlieq/9Imt
8gmQW3gwR+Dcm2CyCrv8E74EfZIdjKvJ6whGpb4LRVjCi9irlkBAHVxW8pMWj/Um
hppjfor8qSxFApYjFttpHdhQt6ZY1Cz3S8fBk1OBRALellBpAhf6Ke4gPMoIfgwC
hRDOk+Gw04wSFd8eoyrwvyTwl98Py3ucAKMZOacw0EkyuUf0qDQAQ94Bol1WZ52h
6rhbXkZ7i/siESnhfcTx+0XLuNYOJk3yxG5fE6PKsS4yi945Uz7/jzAmMmH3ngFH
WssxRtvjp+bYwPvYodqPU3X+FQEfBu/xpwZwm9sxp22FNAs52f8+VySWCe7gVE5J
WDshgUEYTE4P0jF1xSi36Di4hKbvLGOsiZtdJeV25pIXugRRE6UvGJmN6msZw4Jq
Kg+ALWum6Z/DgKGpzFSdV5S2v/D5lwBpd7DOfPmNt8i/+CqY+I9/ROW4W+pkDBuL
it9TNspi7cFBYBVV9Qw18nz2ThROG6mNzlqumdTS+20kcKLB7sXn5e+ih/oDCnQD
oPc3YOZmL6oQrC2a6GT0TTqNbOtB616Lc1YUskmcGwDjsol3b0M6ANyBshldCAif
aU5lwdSjNVgOlUVunRJ0219JjLOEQBKpUB+X38iKSPR80R+PzxPXm5cLFyS1eEsc
cIuY8epzEu4GYjFQJs7VUEAC5jRUAXfq9uuqhbZNLzYFqAkbClSdNoFltiX0G2w3
/PnPwgtkVGymyEWALHEtxmzPKuQwb3sgSQcDc9RNtYcEG9fPoQGEW4eLHL5EmX26
cie0gS/Lr09UkC+29GSflbZ7nuAAN74dBfKQgWFWGSXq86cjsFFfZHCxK/LM7Evb
S2PTfsOES1/nJjF9ReWDbX27HDWKUvIVUDoDwFiU38PRjQWFpWwdbfWAwElFqiBW
auwMHV1pEd5Ho3cyLeAeWf5DOogbT2qLZ/xXxhlFeD7+ljRMUXMGv7UWbSgFp4Tt
GtxANNQbAhKNmN8meWWfee4963Lq5Cn3y7SDwq+LDm3iURBEa3Tg0OnEtg/67UV7
vJieQCKgqN/2E8/C9B5iaVCCkQuwtElmoXRvuZrja0sKHF3AaPJwmodM3hxEVLdU
iQo1lqCLio+E6Ae3RKGYbTRXQljqyxInjxRbCoBxv13MOrriaLkPsKpyBFvZIPon
jarFfanNIXq6B56qNI7dVVYlS/+sWzYDh0zE1z9rKsnt9OTyE7TNt1XhHpDxVjFs
LONVXqeGf1L0t5q99/VSxQ9kfG/ZyHY0u1x2GR29A7nmfxc2No3dzGzEbZW4JxyM
TK/Uvf6GhPvH4i6eQoKI8lBTVtu57DnpYX5l9N/LIlRFm15JVKuPNxmt5G4Nh4FK
z/ptjbGV0j3EItdainiXeuCoejTWsvTBrSUbNHv6o4oXHLGYVa1eHQLQEPYz20SC
+H0d5vTo2TCAZybPRgOjsqzm7ZOypJOQaUlc1b67KbAy4Lnj5wvysLjVXgt5TNaf
H5FbRqusksmFAjniFy6+8Z7N7dZ7XPCA0lH96P0ncsM8AgpmoX2J9MqjiuCz+gWb
+H+80wU13jfVbsdE9Q7Vx9JPRcKX2KuqpXuzVcUeCcmXYTw0lNcFa8ZOpjHbpgsl
SbNjXuwpVYb1jVaxpFLvbzzNrUHA2wUrjM5fZT0gPhTTLDRSkuHGXxkVhrylYiAB
V2v+AEaorY1ZMZ+DpoR/vG44pdJlosadQHF40N4Hv8i4P3tVvwqvfDNVLZ/zpdIc
kZbjmr4ZEtVUAXMOwRftwKZfQessecbksRI/z7/PA/KvbgEmxZy5O6HS+bNyRNuM
ACkaXN6+shHrGY62vGcYM83fXki6PYnulxh3B7sqLok60VVHZRic8T+IodepJihA
MqIFlT2Q5KBxyx+Wduc/n4huyseC+y3ycGYzfken2rULAiSPI36LRmo0O4DThNds
6jKPyU7gMQrn7h//Ji+8JebBQwIWLt06tNPL4+XUhF8E8E/yACc3DiCiQ43NuPUS
7oIDV4aRtdBIny6HGkyf/Fhn26Jb6ebkOku+gf3yTO0lvB6U44DTghU6lpuUHre1
qVrHNn1hTrqTYHvQSuNpDopQy8De+cH6JZh3CkhyDITbUSUloKAO7YX4iIGDsGK2
1+SMN5u/To9Fk+f28Pv0eCqulPj3AEoK328OdHh5EfmDLEC9f5impR4j6adeXILT
ZxjHTbaLIvu4xcuFhtnFDLkSTcxdojqMe52c9jwvENSroDCA13QRXAFf9DkQNf2b
yniVOaMhaAAJVwtvk59DDgh6E/eM04AHz5MTOGUxrKVDdh43X3IKcK5Lx0NWgRG5
eIXeCBe6YCG6kAscA+ZtSXQ6WY/1p2j2Wn1c/ng8ZcSwT8OCz8JU1S1z5sNM+6jd
QzCEZSMiZP0yLUASdQGOc9z2P8Xd/86W0zUMhSBhl0SNByBOe+9ilVvi4Ro4WCkC
DPKSbn28cq3H0fVFGXUm8+CgayG3QXLZhPoguRuFs/+qaGHTDVCZi+fBvAQiCzwB
JMhVqwX29F8JA5GPQotKspQhB6BQsuEYKlAAHa+dbonWkdUOYbX2G+y5OpAHYKFv
a72e2QvFqz2fxf0EC/ZgqRWhPrIcqXL3AwqLgPGiWc2fUgbck1qwcZQCOZ9+nuh7
dVjOUP2gN0miM2KlHZ3zfteeg4lSiQe/GuXbLE+DXfbidL1+SjR70X7FZMolYbIa
5mU8kSljRK4cOLdtSl5IwwirGJZebiN4pznFSz64lFSLbIzsTzrah6mu3t8Fgu4I
lew2erdren65ETPfQmTm0NrLJYGTvYN3rs8QpZnDi4zIICH0At9yBeuyqc6BRzoR
xUHj6dRMPThiaY7zzGsph8xlLG9gCA94Nk03n+vUBAo71pNwf1Af/UWwHDwcgCvN
lVDcekWa2eiQvimcvrwdeQvZ3RUR3k9iGzmMtQ7A0J5OCzxNEzBoid4o9Cta5uxt
mS5CVIKh+0EXueVJzlX+77EctrxVCW4Dj1ejcdZmcOs4sMfzsFPeAle82LRpXVh6
7cJa2rGUxT1LHALcu3456uqqBCe8e9AGo4CinLGag7snecg3avee48YY2h6C2TRo
hewHvw+Of950TB8n5MCTZrlem6cQNEt+fQnTA9AYnBvUx3J8ZCatjIjozItCEPxt
HraO+n5HN9hclSrCs9Fuh8zBgulBJxmnbHrTKPktlBXIyLRMVsr0wByRFZJUVBpS
BL68+QVdHHrGWSZGQq7SB9XV8WYmMV5252o/B2AVJ7/AnH777AaoVY745ZYqniRz
zakI1dh8G9RItXmuusqNjIpSCAwid7K3p7HyNISnUk2G3fMclQJT//5KvxN04NoP
qOCzfX/f8ePqU8sp26dqzLWHs8ejqdKdxXzgkVCPUljmutet3x7VHV761KYOOfg0
Xw466Q9YdWvvxJYQ0G8vfh5gi6+rkMLW1aU/foc2UWF9hElRDEq7Qhg+fE2sWac+
ct0LjzvKPFeIxVtNFOZ3LTlBPzTKNFABQW2zs1v1S8XG1g6qA8wYAompxvEmT9lr
GmOKOEfsZ+VoBn9nWDNugGotNOeU1YYluNd7B9FOYo9jg/O70oBtaH2tGe0t+6+a
WJlPyaINrUlGwc1ylyPeB/mIjK3ii0f5BJH5EiQUiC5r6/stjVXq/hbNyVWdlAgH
x6Hz9scEdZ9kGJuItSiBi/zXq7hc6UqQAJG2zB2Iw6yDGG+uBlP/1OyGylHTdTla
cTqgAt8SxBcWWldsIKUnvt8EsKFQpO3nTedJM6wFMm3GMMrGIfhTnUBnJvzCk/g+
uReNsg/dlfNP0x/ksG3FhiPbAFDiqZQIvrkJZ9ev0HKoC8h8tkRoZKEVmr3qBUpz
xRR+SymCIlC8dX/iTQfZbSQYIEyg73qtVesHtvbnwtjYUPcRMN1UztDO9tjIT6oV
ncz3VaEqU1pqEQF8M5FXPuYr+SN8H7QsgxwddN7TWNaIjxIlsByR1kosEPHd9zOc
s4l1vzuXz/sdWAZGnTIXpuJ79KwWINL99R3eb2e70ru8JDA4q7LANzBWQ5+qvS6a
hDF98vRjZkRQvj/jujLx9bCPUO3k0M05rNQSt+jpCOS7slMCGtdKaHjn1PkBV6zU
hoHoee8qU7ZFRnUQbV74hjuND6gECgF+cpBD5t9xZvlp4Wnpwjvzy9jvhy5CNLCh
cKuUe5PAOyL0JqtX8iniGTEfATQLffqRnMaVoyKYR/lXKu5uYRuARNt8I384qLdc
vrh0l+7t5K9hMxXhYqmQo511MOkw6VKJsecTDEEVBqWBEEYr72FvU+jY23MOtud5
GCq+sQnYaCXo4h72/1hdB6SO+VtYQjEMPJ/Eerzbla01OyvroCId+C6rEaqb6Tw/
e8WRBbjA5Bg5258+J6y6Z5Kmmd13nUamXOqelYIKiTV4sHOvtxCHu8MrRmtkJPGl
iqBZ19gGcydWkRHYIBOBOaSiKtA5OsUETlJgLWhCKficAjbJJ1VI2zbnYd+pEuZO
vYBgO7i/kDE9WVXB1ayvw4bFY7Y5I8NvJPL9sEv1RBqfzreb+IfFn9FdN1RerFIb
RsLA5ymSf3X2scbn1zBEkDgw5DbSM/cwfBgVRpScpyKxIleE1qLsW9WdmpmExb/y
ouncUM9JdqeEWjzt8NtrVGkXHTFp2Uam80eCAyCNvRMI0JPNlAb0Fr2wWLmue7W1
h5xHiJ8qAPy4BBonIkPDG/9ZckyZB1Ng6HULi4FXbwBwwRv0egQ8uJjAI3psXnn8
HZ4euUQ9NkA5iAMeQ2am7aAuPgqLq0Yj7WasSKl408atTlbkbGTTA3OF8EIiKK6I
XT4OlH2l1BEwuO8OF48n7Ed95nKSSsjkSA0/Odj0NwOmVIA+EcqZ6WLP6LuS+f/N
XBBlSbRLjyQ8y+0+9C14XqTASSglgaw4/NowxkuskAxEkHEJtqWxXReWxNRLymSw
gi2h8DGpfOWmggERLcu1oDYWjJaiCYwOWC/seBJWEYb5EIZo/mnfcXiKYL8tE5px
cwmjAiAu4elb6sFVPDAF7fPJNGbw7nogXJe1fmln0j/Hc7OAkuyjOZyk9I8SAzgW
6JduQO7tzqfTLRtirz5zBljeSgG9cUEQVap5JvblZGmkpJ6V9vpQhgX1svQuMLzr
XQC4KiPIGYSUEUtLHkgzPpxUSlJMcN050rRIwEuU0UKm3Kv/xr3K3WWeXbnSz7rH
icBFXLCKgWZYCcPr++dQWnITaHQCIGifyjVsvwip0vQDkyspR5FwhCZq/XuaJFLg
SR1EcsB9xCRDhB238mnGDVmVeU8JIgOY5yQrfUlz0hq8WCaCiQBOEjLahDLt/oun
OwpO/7VHGN5SQe48lGbkiFeUmAQtTqI8S524RIbL9xLt2s09aiTPx448jQliTgQV
1b4PZNRapyWYUHsWCW71ihdNC104OgCkbkSiG3uPgkCK+SA/CmjoDkmLiNKd0bwX
FMAPx7MYPzlPPAxf0RdEzi/w3l9nSRLVdPq5lxBvCwkxP96F0N8vqFUdeWqsnmDI
TZ3cr5DS8QBW3YsI/yZ6tgtoDp4x84Aghk+LZn8t0UE63gWfV9N2tvCJYGsQLy3d
bwXwSxaZj6lcA/E1dz5rWRorhsXt++XrxCsJKkLOkW4QyDYPoXzmSwRVEtMZJmow
KVLmpZIlWcm6ss0IvqI1xrIvboNjnU9Mf6xTeX8VwCfLSbHhL4fFTwMhIjCDbYZp
sQMfXaqlB657XIqQoc3ocrjhVlYraujmQlzsOioeJWxs0GaSdIEEMAHJj0y4byE4
p1T9iQRB+hjmjATFnr/55s3pOiuZOOg++Qlo1p9vmtzwIwXFBFbGHBRlbwwD/0Lu
L1H1qa7cdP4NNCuAa9nVzVbxUtRT0D3z+9LuBeKP8fjYWV6kllwUNT/OJMrSCEPC
KSUN/wFTYI/knvnOfE441CcWqhgUs1lkhbCFS1noVEzNOQOiQv0ua1XFXmX3Wv6c
P12PtWADk/QNIh+HdKTNyhadwkgD6u2YLiEADqVHwBZmcxTnTu2U1U0QLmMiwf4K
iWH5p1Yd1p4WyEKt3qk24Lg+xy6oj3sllAw4qXBjy5AcsXDjbS0OyjGj9NpGzImr
GCHg+dL49Zfwec1NHbD6DmooTqLpYkoLPcPVr2ct6AftuKw12Gae8TTyp/8LoESA
0HYQXYgnsh5x2+gdQus9L/OsbPZZNK07GMC3s1izvhuh/axQaF0YB2iTuHhP7Jf0
t4/3Ajlym8304WFlU+604USXMzfJghkNNFuwgQNF0EYlhnpcvRy+XvmeRkiYB+W0
3XXL2U4PZC1JxfV3J5K92rU704E6WSAFxuyJRLhc33NXj3oAQYKwKhsgf8jzGbqx
W4TNYE96GoMa+YoNMHaxYsYj0hCQB1T/3PEBvmYFcSlQTzgJ8Kp3nugiSv5X+Loq
oHCA0bDlJXljA20iG0k2X7HVyso5OTlRT1qQuh7TtQE1H8ux/aPo2/DfSEHXqnFF
lRKK6HrddfVXCHm/F7qSq90JoaISpLccoPGFvEdXFcwari7GMeiw3vITVTB8hyPq
f0yR+SRotZYLpxt6GXyo8KQWZX9E4a1UcLkufWNS8LieBAmJDJYHqI3xcl+XquW2
2/elL9OFAW+oAQEaO8Xq8AgLjoxvbfLMF0hoHMJ8qGL3SowGUxaJ7EFGIoEIi8hZ
bYN+WM/uXJ6M/d+tWLRJBIiLVB5aqKTBg1jHILgO+OjIeSe3ScGna3kPUCvURAfM
cJOPgPWzjanQO2ExPQo/JSbuu4xLneYhr7hXN/VBqYDyAOzq7BInU8jX+OHhzsAk
8XMHIIvSuVeU4wYiPN6eHYu8wQLc9Uwg701sWxsATGm38RYT7JSMrvasMHNu+pqJ
LuiRTKZuvuy3CS20JBuCHezd8mMYW8IpxvIvj+Bq/OUuQP3Lga6QEYxWz1dHUcLq
NAFn13D4vTPmzdcqNdKoUGYAncBAcOazv/VpJbSfGPbW3+qzKYnPWsN2OD3nGV4A
Ev1CLPQjjhBMc3JzIbTOaJrP9eMaDxPERFWjVS2yfJxUO6BEZhCVxDFdVOLPSfGb
mNn4jOQbyNTLQMKXY9Atug26iylTAnbdg1v4b/B3t+i4sbQ5+o/aXJMIZdobO9B7
4zURuEJd/KJrCxng0nBGajx5f1EolJJhXNqHGk3WcJciIZw2SHd6CMl97Ad6Kx5a
ZDFHL1ltalfAez8MBOGnwsImsWqPxysuxZOe5jRbdVeCIMcDPv1pp2t/Ijf2/0E3
6JuHCkxem2WMLtIS8HecS+iomFDboApavq3FSbRsmiVyT6Ch4gLi0KHobXSyOecb
Zaak5TC8azjj9+ztCzEYQYORBmGuztTuUmBnTN1I7Usmv9Mc6wTS9NMzoRSFgjI+
3vFGQ50BdrzTsUHiXsVkTbSoHX8tJ/hv7FJ7elWKXc738HKIBYZuGZ+fOQXkwKyN
g+PuintC1b1MPWdmoFxLkX5LQ2f97XqpZ5sIUgvuqnQyV77yk30MvFsWi32SIFMj
OuAEfIa2tJDwrlbRzPWvegW/Cj+NsXeN9I3dGW5YEKbVQ7W3+hnasE0R2wdGC25j
7pKowPWlQhgdzVDpZ6WugNGhUAwJ5ifMRsueSwU+7wQiA4Fvomsez2Oj4cNJUYbO
KPBEn3VfSV5nMNKtkBbqudF5V+/UWWqLX4bTGk+mjzfsA13AVSFj4idQDZlYsH4a
/ivJtkKOAlu6pyVGRV/AzhNRVUkARpGM8bO5SolxrQBZ0rUYqCAbVRWHtl+CHRFC
YdF7mV1Nq9rWeiBLx5IkS9omS/CLztSZc91C3VMVsM99yq9iUeFGUnAnB7dH7z0E
dO6JIyOBL1OPIJWahbGp97A+pu+vfiufr94wFeCoE58YwxfvjisYWr0yzcpkNe6m
vWENPqe8zY7szhgHhLBGvZYjPJIS16qONqn2Ji2bSbAziNctqWhtouWpxoto4ksJ
iRPaPvX5uJy0Q0eQXWIOY7hoGWop9Rw1Cs6XV73t9mMgQJwLstVGQj+ECZsZqfzk
wAeZ8KZNfAsiLHEieqUwE/0H8Fg4oh/SrEHZ2n/6IdJ1HhD+T4awLhcNEMmpV+62
pRbyP/ZpOaexpFjUN/cnpRRah5q5GzXD658t/m8USb+ODsRhQXgOUXfk2FnLjz/e
6LMEUY+8MJVmUsOpLnVLz0PgIehOuZOp3quSvX4aQJjDfxO62wxCCGjYnp8pGGbB
ZkgitcXAKrQ8CZil/GZ+/UGwH53E/DKpvEWJDscliz7ZpcPofS6sPlGT3W4+KUV6
ngSllYLVIVNbNFquvSYzxLBVvxzcWO0Xdiy/U+ntRPe9uTsNqm++JDEiaX6WATSg
PBtD0Wgm38zxYIbLKOz4+G2hVyw8WXs6nPxH7XrDuTL3NhDOm4HznWu55hjMdeIp
iUfw+xaApoT9z0gczb5dK+QZ+UdMrZOUAtUamSkFrFHnC/kkLv9DDB7oFOWfi+7e
JvkRxBy0tdBhGwbz+wF+j+tluMQ2BggpaJAkRGAMu/ZfZpVLVR3/UyxfqOeEBbDW
u9owRWZCj+z4IpSWwF0/ZTsiOCa5hVOnQv+mxM8N///UVtEMaJNK2mhxZ2C4L4y4
SX6C8YCaMq4ZbNHCQudXFHX/7JGI0GfX5nXqqLyt72I9mlWuAKjlVo4eflO/MhXk
JmNP/y1H+NtTxaIeXLVQ+VM3mmj1dLO5Nsoj4C8x4Xg8sIcchvspHECm4UgvdFYn
VyL+uIrWq/Bs5eB1jIRkcqIYYlKQLj6QHQJWoMiv2Bj6YnvkKsr5xmlMEjVAAqGK
mQSHNJU86hGOGTlXnSK7yCDbUcvH3xZVNhJagTAwBOOroVWK7YK/dvgR3vo2kNz8
1HNRe5sodlbrx7jGFX8QNiis87sSgjC6LlNKfP8coae3lrGYDv3sR1SN18BLvfv+
xp3JlPSMDhtwI5rGI3QVxhZB1Xs9E4h6YZk4d5pyeu3xbpOhD3rMPqydh7R8SBJi
jCy80hxQI/mRzPuu7TSvfKKk+rQrDGlJsfnI9GLNq1LP22X86pA85ZwGsYizMfVM
W4jb7iBEAVEA4RGvELMBqMEOM1db/N/4nh0BtPb2a4KzAJ67vaA9GGviWlBmbB78
39zELPzdMXulESa/1zhiRmUiQdVGkhtNg/1AKKWbW54KOkyo72NS4DeiosSzJlpm
YOi0WbyfbDdWquKQvTZ2ztDZn9d9L2cLDSxKZt4udcUWZCyQbO8sXY1lH1kF8uf1
Dud7U9aG8K5kD5OJFH5Rv0iStMAqJQ3yioE+j+OXyw/MaBcVHVdKlo2HHfb+qVX+
jSS8jT5mmA8sWwvPA/pMIwN7TapTBuGbW/59dsnqr02CLR9xRBzYNAlhCWEtK/tK
XrCQBN9T74Jmm7y7TRlFuP3qFpxk0jaHEWlDQKF2hVNeLt84IZVC+M7uKbGkk+oN
4FgXS4Zy6qLqfKFAgowx7Rf/PkqMyVqF/pYPOyOuL5kGulxGnqy3qRnPFr93mVKj
YW2jcBJhwATWOasopAAhsSJTgsx1s5L1nk7+zfTuUK++3rjpoWpsVvT83ZEEJGRo
3pnCub2YS4cvNaOx0j3YREy2IkXPiN4OVqGtGCE/+QTOEw0pElvffEKxtKjBYhWk
EQVG+qc2gmtjjODIvSfWUPp8y+ww6Utaw5e2Ng/2lhavwsUACEaagj0VbPFH47I/
meBXPTSDKoKL3G5vjPFB1Gt9/RLk1NzBEYwjXrMW34N6/0hp9aUwqARTD7Dz746y
/hYCftFpVAYst4rtLpW6+UWaMbiwS/DZeqw5KblP/oThJpuYBvFSCaFIoUdP+94f
3FtEXz7tX6ifzvQXNbHaBabKBHKKQlSK30V4bNhhPI8l7/YxKVfC7m/htG+pN3oG
QGQBktUrSmd18WYKixaYJN2Fkzr5lmYAAt78ATbjQITxYvjWD36xZS2avKmzh4S7
foJQqGEFxWbsV4t34TX5VAqFx+q0Is+Et8EJ4tyv5Dd2NBa5iM51wOlV5BZXg3dI
cJRLjwIje+TicnRCtU4Le54l4KCPz1d6re8NmLpv76QuZ4St6d0ydFRsrx/Pl40+
jv7jEbDeCtgDa71IbACV5yeYPwt8S/2sM1G2PAZhiqV0/4e2RZewEt2og5RlaEcx
x8xFBvGV/dW6BTq6PzbN/oke2JhKQzGALPXwqgzwbmHFCcGMmxGiVCZvsgepsKng
ww/HHUw1xvsw3oJ80LJkeVKMRzEnsGbVlpLMUEA/fl/fIwD7wTGq9PC5UrQ2g5yz
EJ+AS5LdvpjvjToizra09KGSuSZzTqURysMZLZylIR/+5juvMfGcmLK3O/dh0gtb
0l8cG1AweAiCSxufEbqcApcbs09HJfmPlzeUhvfpObvW8GXzKrEiXUYNw8wb8jWm
rxwM9oXPpFSb3OUAVWBxnvi9+UOPFWEg4mjrWCpHKHNg1Voit0hzOYrD1K3T0/pJ
JwwD5NYvISPRjCrdwX/kdEb5lLlSe+MWPAW1joKBC64WQvWgUUe5q1pF1y2bVM16
gK16HoBrCDXAxX5aF7dlgUmbevB7YbTojej9sWMQVWmMcXEkZoT8i3ErM/nhV/1I
8ceNxPpWvKllYV58+FjbDxl9DGlIOvyjw+k5rEA/g5115BFY1QxnmL64Lzua9Blp
yexq1KLFZZOdDy7zE43BZClr5elb3YhrY3rF2Qj+q+UwH7ycCL8pAHNAFhB8miyd
rktt4ivvoabOL71V9Pnz830uLLiEIIEBPOyWAkM2DfZAWdgJsXVO1klY2CUPj+F2
qB1RAPx6Wl8L2JIEZUlif1PgTZ08mMJRdsuEkiWvLukVQAlRbSEcGW0nQWVD5+KQ
+E+LeAaklLfWXvk0B1v05CWn6v/NN86xAhaBF9RUuJPxx+GeVABkZa+kjpemONFQ
F1cKU9/5WtEEC+f9I04ei3K1zirjAyxOXdxuB9P8RF5PCgYfWT4LBbwbvHW8Fz5V
Nv0mDCgd0vByZkYyVF2t7UnX0XUurF+UEGp1QkmPaYME83QGnvKjn86W0qcbLkAt
WlsyGHxtPeP4MXH+rUCS5oWjsEH62GCs0DbG1zXt7awNcHRvDGUfgUSK+Sz3D3WX
1t/EWJDWTSMAJ9WwcWEBe/GXReq2KGxbsOi6ao/z9xUDzbu2VtKzo8MsCSbt+Wu0
xoW7riPBwm2vVq/m7PqjovqQ+FsplE3IkzJjNguPwJnz+rCOIMktZ+CYEQkm/vIM
amHNdPGXtNCMnWE5UK+zDHBKpV1SnOczGzd8zS+bTiueSNkKMAOiVmFpeRrLCrRE
g/YcPpgCokyz9HEz6+Fu1fkWJbCV6kkaGlqBYYlfa7PNEbih8TsJr/PkjJkSthjF
Sp2gp3Z2wfA9rqEhOpkFesRq/1yPJDbb+G8QpgRVZ/PuRv9TAO7MVwclFFO8ECC8
SdB8xqCDVZQKUWV1dOxEpIjVSWP9jifbeje/nyUhMxWh189bIBzKfDo4hi/XpUfV
KkUASp5KRbWgYMYx0fARRNUsVjvKcDO4dtjbpzvkyY8GdLQMAhM+9jky9Ur+MXgL
dJGV4qMbgWeOjbDkxugCCvqYKqMBYrFqfLprQh9aJVrITpUkPrV2CZMPzYfNPgjY
HRNHVAE7rrJ2f/VnOEhXbMp4G2jvwMiZOjod+khzTgmfHLfoN88dMiqbw/FQ/YJ/
g9qYhnkY4d1yLlSpjQZ8cGmeRYqJIyW/AZruss1p7fAVrvO/GhY6eU8ZsVeHzEfN
3fjwIishr6HEKrc/+sGS8Pn+6J2ZUsHXFP2PrGnpgL5jKlOvsekk1WiqlhXfp5o7
3JaJkGPjajTY6rKFd2ZzscEHVTImWAmSo4/cOhy44z+GAvOWxIqr7dV4eHgjewlS
Oc374pRJb03fqT/MNvDPMTD0bLVYpt7okBj8s3TQ/btsUVFYTex/FioB+3uxlJhQ
zWCmOiUFaS+59kYwdRJlJ0l4Yx8UWCZJM+cyMFa++QB6pWWKIFI4kGKz76kL3zkB
vbxVuap09B2igfJDfFECHLM4oQERkfryUtPZFcp5a68m47EoGlEUJpwICJJNHS9m
rDG4Tg+cjNdK04s0AIWnxbx/G3smT2Rr5rqBlmoBcFxCBhHftOXCtwEIgCxd/1a+
WPV4iGsXbdAEdXliPsIwHBTO9h3MC6HfELKnZmGK37E/7ifCiinA0Z3KcsqgnIYv
r/b9Mo89i0IXwcOA6Iw5VMD+97WTmkafp92G6GJlKjqp7CVhuiwVFwZR9GkLGMDl
ph0Br4EwRt+vng5GFl/Ob4hh1V69WFNBZHpJR+S5PXUwaBDOVrxBc61tW3t47XTM
vopDqc5/GMrIDkWG0RQD+qVQCOyV8jCUEZZ4NVYfBxk3mmpvk3ThTzAXrEx/sMAv
d7EqqKBSjbYdKUHkzKCUlyCgiJo5djd3/RGc4TqjMKkkXAWCN1daq07mD6yT8e0s
nDSr14I6LoeSYjCWv67dWjQSKxenycCOMIsTjPijB9pYot+cDEYQQ8ZgFt9nFn+s
ou+jnZRkVg1so0/lcFXumR3UT17w97iMxBB4qKf2H0KLH/6cu+hjjoApvlZKrp2Y
UxNFFKoGY8fXhmfH31UcYqtHAMl4htv5dt8roX7ESCXCB34T/9dFoGeeP/eaLRP3
QrDT7qxs4IV8fCnXk6My03lpBYnzeWAqPa27rbw7qzxrUQBSqxG5/QPGbC1LLRSC
1lmMn+D/w/GrLX4MjR5ENcW6Bi51XMgjVsjzg9BXALW/LpH9rDCTEke1L3S2qZKv
YFoKgSBGJm8fV6lWNhNaO0ImEl1fX8g63ikgHLCn6P1vfMUTyypa+oOFBhV7AdT7
ts7NGyPu52T5tuU8TaplsBhm9ONRbbatqBHDfLy9II4W69DcXhP7m4bRd5H9xecF
aOPy9Jt4moJ7fjblVvJrF3mpdAvjpddRjjJawLzbOaLpysOaKTnjGoQhJjdq8Zek
021ioTS/ra2i9WgH+/4h18gHreMWiMtita0LUGNaijbua2iXKM/sjovpsEXOaIYR
EqtGo7u5ECq7qK1Y2p5A9KF1oEbt5Qqo/bzQXKAYY71cCliqdMLtSwQws+55kCv9
jPowHiTupIPfkbD+T7QgLqJOmNWSETmr4ir4hEhi6QJJX9B9FBO/ser+KwnTLzBY
iikB1IrZTQis8yhgK7oh9iT/gDVMlLI5k1gB7nafryGbsi/ZQas4S5qvhZ+QPoEl
Gnk2P4qJMvq23XaPthNuXH0vQeDKm5Up2FCUY+KD6Pm0sYMbSHNasVu96eoDWoz3
RwfHbDbbB3eD5T2IE85iUeElo8iKs3bJYBqoAo/FdYHU0iSEkVGa2LIjKjkgfwP3
Yy3Mzdw1N2udtNMXq0mdZqFUUkKFllfEJ9HZwZF9VsDtaBPCEPnbNGhIjGBBMo9Y
MxHno5gCxGw0PxfgXpUNOJ7/l7be5y6xHezITlemeVAzdke91WVOHo3gDVbV6r7n
Msos8GjzXkVNL/saTHLO+zCwVWaASereDXCjHZVeMuNQetoSj5d/mVu28AxZM1sD
lzxgoxleTE2Q5apgpyNeg2Des4P0ciZJ3GHXWcCbM8xqozNn7Isz3qLQXuWUI2pk
qhBM6ejsnFo7pw2ihsjGb11PzLgsv7z1C8bHthdEtNpmQGk9NhKsZ5W3B1MWlEaX
GII9aA5ntooFVdtb7QF+8t+mS/93TJm9jn+rF6KkIVVotHG84yeA1Ee9BLA06LgM
f90G1CO9JReplJTILZQzXJ07U8FSKoU74923J+USR5W3F0jRIbg+7yWMxJ+vB27Z
u9F4EpgP7zi9lhAn0Wjv9MtTzktnNU9PNZGgHyGqbUfxSUlW+ReNn/YtbwE/Ocuq
Pdat3E8+ikIbAXKOVC4Ekr735AD3F1oWMziN1A/ThYliKsD/vbM5EV6pCfg8tTx4
jomqJFFcI0PNN7Qz18RC8ixfXHAN6wrp10BveCrNL/xe19fE2C7KFFR0SuzX5COE
C25UVz8MpbYoUs8gngehjwYY+XsQPuXMvnn3CJgiF9wWu9VcUxe7YMPAhOQNRD1e
KKnLp7ReuWgvhBKk1df0T5N4QzvH+roL4SyeGQTaV8o/xvk45uopHIjggU22mUxK
8ib54xnWDzKLIYtJ0BGlGu0yai9is0sMli7B3k9zIVowrF5/qEl8DD5Cr/wFaThw
CuevGQRLizgxyy6IFWDsRvI7QovzKHiRZ2xBFKHpMgPM3iOnncuH13nG00sVJzyK
Xuxj0Wfb1LsSdb0bC4P4Ca1ry2PxKInt4quufxUivdBYYpHz6HzvjVfoej1VWW6X
WRiwW8xWFqFPzNGZiI0lt+ul9RuGXl3pVS9/ujmpWYKDtayEzg93GgADKX/4Wtvo
CVs4QOmS8uB3SJ6DdkB10X69Pg8KGA2zPolWEFr9OCSazFhAkLw5JCW1QkpDzqqk
WGbL6y2HrZNKJBSSveYRVGZn2oO4D3MiUKUE43JgU3xlL50ccooL2O+TTdlQDtLV
oDswXUaM4VPoTQ7PaITKtL9LMPv9aQuqACJnmBGRNHU31cX2ciZj/O0JKQ6qyCK1
GkuYi094Y8GnuGIZUIjB3tLbl/qJv8A7ToGaiQ02uDwVOQPStuPp5QdgQlyem/ut
6WDmTWDzjyJSKDefa+uQFbadb7DqAxHxioSHoGl9jt8Dy9sNdvai4sdkJqWseico
ymP/27thfwGzgLNXWa5VS6MrYyfCtH7zhBqnVhQFSsyuWTM/iToi5+fZvh2NOK8S
79roBqbOWwpr6XEIkFmtxFND3b1Mrq/gJzECE+eplUzIJXCAZEh8Rt6cLicxzn0x
n4RTVltNBPkhtGZLI0wABgBPZzc7YrcOUoduKjzwztd09Ms647mHYsJEm19njiGE
LjpKGACtL+Z/8S4VVxfQnpAkBbIoHIF59edsuznAW6IpfXl0dL/8UTCY4Ri1EBXh
doMvHuuYmJ95p/6yaXnOqVetKQsMmPlkfEDsE4IAQl7pg9AuE16kfvFjc7lH5R6A
xP3bQIahaJgvuKSWVu5VtjzmiwNNutN9dEK6m9R2agb4zEmMF6PXN7RcdtAQTuiJ
18CDJU2MyyM33SbhYyz1W2jcFoEDtButfI6B71BkKSBWHvEzoR82SQOFxQyX5d/z
5A8J9R6mciIJQabrAtcawkvoEP3Y9sr6zw/Y0hA5gegZb3k8XRRl4KLn+fxVKeul
ICwxQqeVYSaj8W1hggAtclkYMuHJEbs6V+z/9apgijaNiHflQMQFLUDaI0LqGAiR
fLykIBmYEgXhqgpN1JGWxRyaKA3qp77z2hS7NGZ6FyMjrutrrPrS5EUJOcFFI8Fc
tL+8W6PK/CP/gy7UN7LzNUXJ/0bP6f1OtSbs3DaoBAEbTH5XbyexdVn4pnldgFGN
78lIEqr+r5oqgkSeXzbE/n8ZT6zsSec95NB4xdadUiw8H3JlboUOa7d7x/LP9VvB
9ELvRSrNw8foWU96CS6SoKqhmvs42W7w8w5z0eujaKjeCbdCk86S+AqKtG3KT6dH
iklZmaArm2M+bXI8ojoSQq17TGg/+3rLk6HjU5Qr5guLAkV9SEr97+YVRPQsxpTs
8p9KlYS8jbsQP1hdvPoUi8Vw8aCdFvyTmGF1JIL3ozjgk6UldwAFvow8lmpE6PMA
fEafYAe2jvmDd1uxkbdcyzynC6jSAbCxcjPFfuq5UmcE+G9irADxUdQQP1xyRjzw
APaeedJrjxDmkfs+f/MLmBUiAM8JT+pAzyYJsiRx4pyU/o1VFQxtBwWDNAqbgFnG
PJFAJsMNSQGx1m7i/Ch0lA+ww7EZNHojNisiUJCeNwx5WYKNnAeE/gINaWuh6x0e
gOXKjJ9LmtVeGiIvtqdjNcwrnqwimwqX2AoCKgKPqEbylGI1hUWbf62vicnFA6AF
nCA7I4vklKrWHZxULVKyviYvdUq2q0xCyeBPmv8mvUFHV2IM2JGtciyaZSB9xsZA
Se0kY8eQG7orzIBCfX9laEQfVWSh9VWck3K5EUCY8Vw8SHGv9hwd9kTWGPPz9ult
LbsGWlt+x8rMLxyfA1uSFNRZgaep+XV1RIb7kggBZVkJbcVnnjFe+ehCtO05Th3f
Iu/G/7CKpWN8rDcIFG/TfrISrKTnEoWmKrxJnB5a3BOtCErH3QoGND/z06CXUJ/C
kC3m6wsDnnxDZBA+yK5arggsInmZv5W+Yvt67aj41/XpkVcF5rBjAs2a4FtciTgw
t/c70WOdxu7z8CxKPwYCNzN+yFOrf0HLecy3IjrhDZrTdXBHPf9zPZaQHqDSv6ud
51B0es7g7w9q4XZjCLMLcZKr9cKOQJcTmS3U8i5lEaZMOOy8Fp7xaSQxZIv/9t0k
eoDOrC+oqol8It3f1P8TT4RrP7XZpIY4oev1tjUnewuLSwaxI4UYl3MpL+XJskMt
uanWQJW1ROp5xlv/E6/jUBWdffm7EdVIReNBdLaOD4NaE5XudDQoeEaBTNlBz//F
KI/2gNY/56tmLW8zjmWJ/TWfy3EkxiwzEo51JZ21UcN7giKDQTbk48xqhM7kgcG9
lvWXC6hyyChenu6hALyV/JlWiMDmTOImEQdM7rvg3KEVu3u9pIkiw1/m32/qioCk
VJUgE/2/gfhbqNGMxgputDhBPfRV64OAKcaxZTzqJgsfuDf4B1mfAWUR4No4JV++
T+Ct+IBOT2267J3kTKgwTqLnMjYsvezLbAgON4UEDkFmdnKevtEIe6vX614JnTjj
ZYF21LP31h0K4smXJBSSRGrWjYAK82r/7cF0YithpUxP1G+xcxvUdRKUYn0pCubd
FuhLngmClL4Xr01x6M0i8y0cvA+Xc+ajslE2jCUWzMsF7c3dv54yhn1DO38F0Ukk
OXUECgQ8eT9XvjxbbXF1zLm14+bXSf/KPwDU3vFX/JBruGVxgWe4s/5TSBPuZbL6
bv0XbO1rKKPvQfRx4KmlAAH0F7h1D6Fw6UYFJZUiYW2rEeXdF7/oW1jWv8ckYRtg
xzlz+SaqzLADfl1YLXR14fDmIFopK766QsHcKNiC6NIlk94aOVkQhDh3O/8e+Azc
k9V6S4rf+5aPvL9Y4S2hmOHPx6nzlZXOJW9zVkgNFv++QsWSzbN1B9ah7NkdJDRV
2vhBSxPVXR6mLt4NkvpOWiYjKGbFL2co/bwzRNjM+GV4P+HIn3aMC4sIBAA6le9H
7MUq+BqvsgtP+wlXleDGoTO3so66kNli/9R/C6TrPpsjw/A4kSUFc7cdEsDF8YUX
T87R4HFoQK/3PPAUfmnKL9JjKZBFYmFQxao4Fern3LEXPIOK+ubCN4f9azD8WrJy
J7Sa7444ZQKB4L+L29O+Fjdwl9/tMlwZ6x7gj1Urx9cvoyxqkibXTlDX+rM2HEOx
TeRLvxQXobG+oKYDvtwF0ZDPXmIwQz+x57uTxl0Ca8NugfZdTM39tjtZlXm6yFLO
g8xmBf8PxIAMkyr8toZ8Ptb7WVdx74nRBjHDYU9Z+3zdncVksPdIU5Zvt+XZfd2f
tu0M4u/V2PtN7LVdSqGSzzIpldbO3agGiqUeQPI3vJZ2xZWb/jMFpSVuuzbmRHKX
E7Sd58wdNzbaQB4ENYR5Gi+zoWtpKY55KtpdDpf2hirjxn7YWd9chHLIp6KPY3LS
H2toUWi97Y3WxsNMdG4azCiwe7fjohDlD970tq07mxroWfM49L9FUjAXzpZA6oz5
UZfqkKW923w0UYjlEGvofBP/EC30OOwJN7rBYm8E4QQSkXT5+jqnCQjnnxJKFgld
+i/FYnKIXRtByS19y16IAcKqwNKZQM4+E4pJpR1NLzfpQ2p4thOFJWqx2bsXKiE3
0l4L/7mEBE/ddVI6reDHwd130cj6H7PJM0xmxt/d1tp/16esqCwQOi8VDJIUSHiS
+JvEJcE8f6AXZblmP3A4O0hEnW+frpWKtH0IfoUEIf2/zmV1ponWdtuIB4SKsp1R
/b1IboqcI/0RC0UMQn/leDG0VXXndJpt1bNPJpWBcYyJr7o+B0AYODiYjz5BcmNF
IkGOjyU8olq0Ck9jV6fg91Tuqgbedjhxyh4Bu6t7zXRA19ZZiNp8Jd/CU1HahoCJ
pbXoLDwh+FRqBUHLB9w5lX+vkN56N45pjP6/mW3dn4LOoNDrvjtt72viLILCl0Is
mLCbwZcgVd2esygHjr2do4ssP1Nf4qXM4DCmfXct3ZpIjWvZudKwkJaYPa6pHXM2
q9lZSuztpIwIqwolIZQjedILV8Nb5/bM+T+xmnfPUykHVogg1Ql5drWSkJSGUKZj
NYwAyUm5eQAe9LBycAY28j72/N3tTQHbYi4Fc2oFj/7V204Nu/VJ+lNZDjG5kdfd
F96TXzttOgLzzDPZj8O2O+S6q6i5PUXIpVBqbMDbleBEIbTxXD8zE3V0vPqZ/g54
tZqONlQdywHhypAkkPE3lr1dTQrGRQZcUck0c5utT1l81IbUW816q/pPGv3piiuw
e8vj3ewYMLKa6eHaqjYfiRft/kk2nBr+8/j38gj2BGhlDGtL1NZW7Ls8s3/XCIF0
qr/FaVTs23znmzac98TqY/9hHr+gfWyT6aVjhZ93G6grZDW634vGLE4xnGBUrWgl
VDWGTnr95TGVS5LQXqV0482S6rdpkzzgkGEDlROJ7bTpfQTRBUxkiVDFW1c8Cpp5
YKz73xYQpCvGHrudGtZAfC+Tm0qglKpUv5mumZ2GeGEM+90VtEOaJu7mqHXKdstv
GlSog8EPuK9d+8nJLCyVdDkt/oCDshqFsS6NOgrbJvBg1tU7lzBCxz7/bV2nEN2/
EMbgucld9ZMhPPlVp2IzxDJBv3qUbLmf0nrBcIzWavP4sgpvca8XLZFcHfG0nkBF
o7+UvQuEGGUXx6yfQ2J9TuBNI822H2YrlGph3jptIZtkNSalilGBE9yAvyR2OUC8
HmzeenMwgcgXNRW6cdfpMglqyjmtd9n8l0zKGeOHfIvz8QF97VxKrAk17E/xagYo
zBYhD26mOtJs52ja49zpyieHE95+lM0VD1jqMDq1d0SJton0eDjZGLXqqmXs2qJm
Ev1P3bBpsUEMuowKiazaHtJgzlYubKVVumixhP12VdJfquBuEyUc8RAmkvpzxfRV
VGhzGerJGKmpVHD6+uD18Qj/kiVx1q7dPFsf+wYECl4/cR3KPEfmwP/OC/JShqP6
JS7sHUEbTbFoKfjYn1AE/KgqpE1PMZ/PsbjXldOJbP4o/GmGo37sckjQuVauvDiS
Ke4K/i81oa5oy+k0CTU7KLQmepcxXs5S1B6ueN4ViCIajDQDrz9WoxGGBIrktYue
SpMe/KKYm6/rO1vzHZtYja2eK1OOe3Cd1tSpNlXPKITCoXQ9MJHxZVNsYDO56SHh
gzUskxbORpHOqSTus7UWbD+mVuUCpdIWdoCX6CUCqOnDR/5Py7187M3ZvhpQPIYi
ZjubJHw8phOEqNssRNaGd5WqHbHzrO+MNk3xdO3aaXZj/jcW8D5KCcYx6kH1+Gbd
56BDtRbEXBai4V0y2yLUeKrcU3i++ZnaT9pT9uNexYsbv1CUoGEIIXOgllVkOHMM
VSaQuKIpQekG2WEFtf8fB3reC3bWjpWmJxRk5PbjHsG/Mc3I69Xi9JKGyfC5jOsL
lJrA3YLGzsYdBIcbgUkuiEGvPsKlXDmDILW3vS7nL3z0AEsBRlT5eSz4gQlLM13C
Q1x0LkyOEG33pHCC4WbPnQDrToZXqq03n+tNmTkyS6beZ2stPNaJrSUiYvaMjK83
KFJvQpu4/Mx9YxB7/dkPHPlFzpF+yO4pf9WHrMFi6IZIyXqasOR4t7KHkCn6WLvF
Y8lWaMYlPSsAU/hpmkAT4izVrp4rR4uLynqn7ynUO1xrs7KDRgiCJipHV2B9evZV
2Sq0aK3OE1Jb97+6sqnv+Fa4KDp94fwvMxtmlliUa+3KhiuhOxgyOI7UNPmbKKli
Kx1NZlmoRhyOzu2tzIwSzBRQBljaRrmRlG5YdUYu9zK8oSBomA+QcK4zk3PnddMa
7DW7TEqPpN7EzZy3wW4c+M21zQE+u8J80GIlwxWe3ZGq5hmt8LvGrmqDlF9Unegn
Yrv+CGJDrJuoALXKG8eXfM1oIsDVjXzF2kD5xctuzX3o1RZEWuY9ghAuD/hpdVV/
1DXyCP7UZmllDyjyUCYw98u8O/XwxbfayUVH79z6MpEQafPKA1xeqVkzgKP881Rr
LWcNN73gMPqUtfx6Hfu4SOHCOYmlnhXmfW6+pBoUaFLXGjtKbfGISmEhJ8vgaXkS
PVIz6y4zFfI7nDwaMfaAuh9rvVN3AUIActT2W60shdebhpMY+v1nsYopE7NZdmZ9
TYafPrTD8UBIw8NgTaub8WvmDhwCDwErzAJp7xBW0N41jwgfX6crdmYR57wgb4fs
JQnj6edRt6WZDuIF3i3BkvEUNS8BEQSTBNMxA+pl/uRMhsSGjXMtEgGD/hhcw0Rj
D7OCl/xZTS0HGqui8A3Vrd3NUqaQzXus6uKv/IPLnfzlro53gvr1tmj8dHpPacRK
XqnE0zgrHFY5Qci6secbtexAIq9IAcJ3fnUAXBsDLCA5p2yNpO+sNJSOZoN0hwEY
a4Hc8iAbfcr18kdZgsHriQ4r631J/xc4BdPnyy5XCXCVlNayy1pHSdJsEVHMxo/y
RGb51EaBBa3K36SHNyXHj4d/mHyZDVGMWnbAHyY2SWglYSGh4AJMme6/SZZR+ITW
nxaApy35vIbM1+4G3xpwgQDTIJSVD6PlKaN0WlcQgD8ZSk6VKscVJ6mReyQAw9Qd
G+K/TqIZ8MOCxaKoW2GGndvQtUO1rXOBMi8i5x8kftCAriOPHdeesfA5NSpVIeFM
Gaxv4NHi2LFn0S8tSBJpF6AMXRi/VVXSbobBblZNENILQHedHf7woehcf9kkUzEC
MLM1g8RHkO2MtOd1+N+h/tD2LYYCOcDr2HylAxrQ+0xgOvxdTFxRetbqAWwktUMM
4NyYXGbLRKEqRM3Md4Y4aOEbvHfjZ617e6x/jNiRCR6c2jnM0eTjM6UiGivnCh0u
E5EtxftRRrXYg8r801vyIuAB5ITN4VKi7keKdFjAbdQoLgoFDPK9C+UhOwZwwEmV
Q57Ldc8O2DoeGQsOACW61/imukUD9shW+3SUCLtc44CSeYiqS45bbm4gV5See5KH
mNcWvW1mmeCTzGcjBEa+xE3wbh2GHggEaAubpcy++8eIJ4LN9x5MPXIbHo7nM8rd
cjnTbdrF26+QIUIPX7WEJAn/vG8QBmlxMpqO3CMJyQ8wVaYsjq9SN1Uv7E18ilxq
gvLxLkQ6aMAuJZxsOpBtKHSfINtlxRfSVzTw8jIlq+Rivna6H26gP9hQ19i/TI7p
OPtACeqH/AMDaJwhkaIM6xTPpvLX4mJL3PxpLAN/Bnl84hOiNBswqtGpcdWSQ44b
oAokJkAhQLdoDaByknwzFV6Jln4kjxbo3YVboViIuGphYbxK9AgCsg1glLqEIaEY
c/1DrjsDta8qUiu6O1npKCRAspgUxKdCYj70ik/Uy5+l8LlwlTxVHU2ljq/pU1eq
YtEFbC4y2HWMmNMloKdczbxlqIJCmfbexTLet5/jaTAtomnxzqkNrV+pJyRqd0MG
nmjtQsIYt4k1Wz3gT4/by1qiU45L5dKvjvzbzEgi9vyLguQzn61bUrUDjTzxK7bp
AD9KrseUalZX9kJtbtjmuOlApK5tOr1IHa/W2+ziZ88M848ZzMiirNmcsRxYc7MC
TypWbdnp40t3+vdLDqSmLOnZUJQsI2J3sQRlGBNdcYXrCe4Wr/DwxCNV2mirDHTj
Vp41QB64uAHZkjlXBvIoK9ThyZiLAlgLLkOmvc/O/NN2vU35IK4CIx/ZXakKXTz1
AcjeNGVc7lm3M212zdUkSrY9HShKcyzScueS4CPFuIVkvuFGqXOF/n0HmuBO3vOW
TDafzF4a5MPwuHwWvRG35PJmNB0eRMg2Dbj5iIAhbjMIljk3fQ7SoZOpiRb6mocm
iOyGDQ62ZYvfidUPq0x4j3AaxDs1Vp+z6GjbWPpBvNMFUnMop5NrbGPI/72oILfy
PHBZPIlLAMg/EOK7xfrVrxDy21d3+erxLd4cw0rhN8MtpwzNxwPgtEPvtDeeFy/J
dmpajcljvFZT6nug6KYQJn/Y9TZaWON9MX2n6mz013P288k4n16eQ7iqyYJp2Ruc
+IefsYYTEbg6gcTRO9rlX7PHuT6jaPPGrzihzVlyZlzrEUHzfm+9Rhjqmi2uLA1o
7ARqKFx5CTgRuVK4Z1IiPKDn2j2ugQV/JNP4E/x3BE5sQu30tcS4P7ey0PaISbFy
qeYzZgtuhN1tuRAFWntLiMhNLFrOZlKdUWwDL2pxyK490l6uZJa1iE+MknLN9D4X
yaUmxVqvOyN2i46S/G0vkJRLnLtMUn8l9Q45XMED+E049X1AaEtdZxzXwc+d6K3p
wDF6rHG9PNeqlVRx8X6nHqa+Pyw3U8S2y4uDcgFSiDVf3XwCE8yCyerKxFYrffLZ
TaPDVuiTq56qdDSTD9UJQrXvMekJwkm8JZHREH7NZ+51q00rtD5Vmnw8g6LuSFae
N2/QHl/0yPvhjoRF0r47WMs2nIY0EZUUA8eo2cFy/msPI7yoHloWeS1Jkrp8n5DW
YFwST1OfyBvm+X7W01gWR4ffekwhtpSWZRzKusA/kEgQRCsgtWQtuedAZD0xDVOL
yzTp8bQLzMqjfwSocYVqoCsHyUM5GNB4VI4cotPH2k2wWUdrcvpQp/roxbFjabml
BEvRk2N5pdEKlQ4fKpclnsJ3/SyVDgII9nEF5BMoxCeDtXkcEMhJgl748/RYG2qh
K/65cFaiKaDLKvBUqYEV1X6QVQbddB9/8L13IQXnsVEvtzn1kl2hW4xFLOLfDio1
8bE525s/jatALmtcWhKWLAQgapKWtBrIhVpBvLpEDbrtNviQlwnG4f84WGpZml50
r5xZP9uxrjZf2eB9Qn4LNmi+5HWCOq3ExCDgj9rVBDJaa4dSNIKJfmUrudsn9Nyv
YjkxDqGp/DIK9E7MJ+yoV5peLCKg/3UTbYYZ7txNPJnNFqCb6MHm1ZiH90zzSDtZ
6LE3V6tA55OXzueDGRpb5xrFaYhNkw7IxM1Gx0/ALOM0/23Byw7/6/wOUv72Zkdf
Zr3gthY8AVegickHB8bRekojp77So4hyNpihvzbOHLjZcAEMpTHWMwWNDarmA24F
QrxNbZQZr7xPkaZAOstoX1utRz1jSEBtxlt7/axb63dLMJyyUbirzdEkvJSY9rFD
35NxbqtfwS3zQM19dmLH2zxNTlpKC/yyBasf2NGL5kWfjfvK+y3GAcAL21OK/nf7
Sdke2xkrKQmvo8hritWvgCLw9plZjwmk/P24UOrAg//GXipVoYsuBq/P3wYVvJ7b
9FiLUNH0rWV877UYCHInlMSr6yIGJ9oWsi72JZ0J0WPAA/2unihQbp9uJnm/IQPW
pC3cMt9vMCqAOBGRmOylu+dO9myDWcJJsL/IRGoKieWdN65jBvOIZM9P90Hs4kxn
qqVXiEUON9jS3VWUATHDMeBeE1WfP9dlZxWzQOZ8IhLDgUYfOHpq/K9SYTrJFgZg
BBV3808da7Hc2LyzqhE9wzeaugWbY3haGP3V6zV4d6xc1SmnAxu9AHNdxQvTlkml
AcG5unt5Yl/1mi8NxRqU6/SlEzHvF2pdy5z05RpCU2iJP8d8Yz+kbqKJjntjfISl
tDNmlbmEpKrOiKHxb77uT6ayawZTeOEuoUlOmgAD0LZzZw7RVrC4FX1/Q4BQdJ99
uXlfVo+rgtx5OIcX6TUsUYyrHnV2CXL+sdgR1PDmvNbipPdVs/YSz/seTwINl/gG
lBDhWJdDHPdybDKgukENTQu42Fq4ecsxrhFLBYeYhXWghkEq7CIUQ4Qi3sCs8pcT
RDq3aFySSxhlmCXg9gQNz1wm3ilMmrZhfAOTFHKQC5XQ5aiXWzgWlLdSTfyP4yPs
7+tKDxoit044R3te/7jqkb/0aXGV9fIxJ2UtqodSbDPkph4HPK1fv8/GFmTKgOff
xDAdTw0qnUQ5I0SQqaIQgnAWoOFHWV7ZWmFZ4BwUslgD9Kvjge10l7Qy4PFP6i4t
ySj/U7nI+f3IDjm+PkAXC4qMIe+6bF4OoRmzs+930ry//QooajJERqSjrAjjvg8c
Q0sHw9Ut0Hj5BvOoa6G8aUPQy+77O9uNsgKPkKmvX5ZT4ITeAbHfMJEgMJkxxqpW
Vxqvi1l2q65RZkoJHMfQut5WCmaIqOUOfLKXdsef2UtA6aVnN4LK7vLHcut4eLkF
vFh/m/IeFdv/9sBNPYi6H6a9NUbwJ+cqm4kIUAUMlLTNP5H5Mx1vAdYZrxHsG/It
2WSOgclsumjlaVAdCduXM9fCqxjwr11jDT12B1jZWJt/BQQTqkpSoq+BUJDDLhCQ
/FJB/f7D3RsfsPwK/hlljvKRHum8IWL1v43U9eSOFnTbHqLLdRbEVqGzQMMWqkHg
Te7Q0+17ZBhkMqwDnOOMhVjJ1MAntozmUDU8idMH+JRoXPOZFpfgutXBBpMNPRg0
0vo2hbcwPB6Dtxusbyz0CuqeyroTZhaAokKCkCOPJG7o3f9CdUqntL4PYtelLe5R
xrZLszkRMKAybY8vSkaQUL4YH8nsTK1e8F4tnpKrfK1dJMTvhF5WglYP1i1faS/K
PuOztdPM+9KzhyVABfYx6CYYAVNvH0YlUETiEjFCUtUgch68/nzYdsWLglhIRXP0
/TyiYgR2IsveVJoVJm1uMI08/9RS31y5pqIykD+hJjhrJZugi8nQJsL0D7PLR2ns
B+Ye2b71Ywj9WCGndcakN/dyKAbD9POB0Zb6gMyoJUJD6a08ahkLdBBqD+gYNV9v
HttX6bp5oLT9QwaWtIzMzQbuUkI6Uo3REZkm92s85/KZZHPwUbVaLKWfjT7gWivs
YJ7InjVDLGNjIS2kCbEROSW3BndmeuEU1b8yRAF9R6d9hTsE6uFC3mc27AYH9wi8
74T/fBkgF1+pEiIWLsbGAX5osB+orB1X6IH0JwW5KWe6JU80OIj+LouAfIZ2Or4x
FZXTz8GhCJmpdWJFWv9cj0ALs1R2CAcKfxiCLlFON46NJzY7lh8dEMtMZVEEq1Bs
bwvQWuZ0sLrVUUrGchNgW/M4hthl/+IJ1Stz6k3i4tng3GpSotR3RXY38FD1Pl/q
5qKp0gF4uOJF4qnPhyyV9CI2YqxLWbxZSvLRS2sDaeL5OuvHBZ96GcWh87gg/Efl
xQk11xiHUK03X4x835/5fACdaeQQBs6OnFNcieBcHt5L2yHHkr/MfOXWJ0yzoaEh
7nSGuCUvzlMAT3W5jFssZ/C+KOuvc3WIAA5lVbyWSM8YCjx5ZHe/U+wB+edMyjl/
oyXbMAacC7wlfbOKftUxWtK6R/xbAb0x4QYR1sDID7zVfG7JRNgG/DRH/r39XwmU
jLmecm/Zmi1unGtUQW/UMxU7sRdRCGdi1YzYj3/MpylhZfP5sMlE82q0LknQZ/wH
QNo8bXPrmTXeXImu1PyqJ1NMgEm82blbZRusqP8D8COljJzGGAX95bGXqJQBweNr
QIQowLiNNZ470fbe/u6cVTu1xGMp7zw/pWPPIIg9rW6H9EbTOlmDBnsa4RVDEaZA
LHkl1zFnVOYbQmxR/ggPy+0xTlvrg/o/Cocb7Pk6qbYzm8ZxFNhV1kMoVAI/NuW6
XYJz3KicL+OgrizeRISUHpsDw/6umKw7JCEYmN7ABbByglh+rkk3JGrxGCt8tQZK
9hsvLi5BJW0ePf6I/TOywTrPTVT4XTd9RIVCqSECW3xMNlTFFPA9Z8O/69Vshw4E
OQKOvuJGdpl/zmiunu9mg0DqGE2FiA7e4Q2fD+P3OWWmBYp7r8yz0Wk7L4B3hg5O
VK/mmIP2neTrlVI2n5wul4KUWJiw791LB3KHy940bbCEcd7lwwh8Akf/h15JJJq3
0DsCMKkGLpveYKlHnf3te+iEtgI5YPymkzZU68w7xtvXUJGC8M0MhEtGZaCBjZ5A
tgU+d27Tzbo0D++Z5YWTPeM3HV90OKvqMyj+OqBLT8r1RToHjhQla8iFwquVJ3uu
z75DLEOb8BvDSaDY6yGMKQTvuAnvyfQKXreGyoYaVHCpYhN9ATi1UtF+hg4n39Fc
v7HUfYyc3M+q8NIZkS0YMwv1qH2fILHJE/X+MQOtDMmVaeF6WU3uR4vPJXuhCHeQ
086FD1Ffx7gkkAZP5QnZe5zm5ntIBB0jtsh9k8CHhN4ZfxqUZK7179QA/GLByP8w
zHRMX0zT3WeZWzHVDOq+RcNEoRBAeUY6gwjRUHpYnI5cZSkzxN7ERlRuFQP8slDE
oluin6AkDNl9oHhjTMVgeaSexQyzVS0eeGoUTPRAO17QNks2RVMfqo0BG8a8tv03
BspVhMSNQ7vvMzVn6SNhpclZer5f7MyKjh9lIa2MCMjk9785no04ULctbQ6KB+P2
u5s+YJIono2iJN+On9CcpA8pWsWxXZBhqN6FWRQ2DvSEC9aHpxXLG+Thrqic2O5U
vuIVRJ8m7V6SsWnEuysO5fF2/Sm6Xshi0jYjJ1ahlKMCLCXjFo+/7buL7m50p/hj
MkbN9cgaDTC/HzfVqnbEcX68VLbim6FGTzNrBo5ELkgQ58pNp3DH9GwlOiEbr0zO
FGtndQ2ot4ac1NwkS0bLFAI2HhfrBwJPmCkzLeS1AIn7E3918RddYb+KcBgFckPI
SA2P4IVNuZkjC9Q7Bt8d9Rjm+ZBQy54mhu0R8TPcgFuF/asodrqQdD8dDR/sgF8O
DtC3lQWGcHlzAfS9DOt4Gis2bxUdvx2YG85WOqPSyzRTG7K5JRpk8U1Ge1BYBL7b
uQH8Vr5IjP3T/EROmD9MYAv1+oKY2R002VpOHxuuA0LKe34VR1mEnnVW5Q9Pw8I/
8jGUkgf5urplMNw22mXRHlsrAUrih48C3RKryQV4j7Umx+668dAHUUThnLeanpVC
EHDkEIuleQ/QBxnnSh88sxbUrtkwzstsIYO8HVOcTnPqUpy1EyC9wqWGUz9/3pJJ
oWzgYSObGqZN2bSJWybehZphzAoDjFJvWsIQ1QyCuESUpJDALMaTFs0g2bY5849H
T1KrGURi/cY2wa7WP5ef2+Dzf+cJMO7WLlz7qEj1BDg4MBWKSBrDLXcdGmdAfLI0
gu3dj0a8no6qcX+e7R55r5qJZ7JfFH9+kuvP2IdW+wSO7NFTkBaxLokysFMnSY3O
KxPMvpd+vNR85hEyz5sHdJg6qAWuWczM9Gt3tx3eTRloIHz1K+991ry1uVINRy/y
7lE0l+dmMHTnwlqPXiLWO9CV0VeFU7k9ZcUNIZBztPNV2ixVx+BCTijlFn4Ec8O9
+OYM4iweH+/ZpcKMPcQOakCLExSlovmOT2R1G5A55gdE/++PyGTwF9j3h/qcIfwV
RDIqxgq+MZ3g+yjZO1XwlMt5tf+3Bo3sbOcWRVCaVn3PyVMl4bliJYnBC8N6dRHw
4t0QbDYQ83c1o0I9DFVu59JlCU886zDBCGE7xWQA4oYpLiZcY6G5uOAqZmH8HSz/
UHX0AJ/lHjX8hTLqNFt65K0D37asAk5kTt4UJUpAIdV1UZo3/Jnxs3xjlNIWKr31
I321aeuyI6WchuSpq6DTPhxiget+OKU02ERUNUv7jFvnS5qL/riow4eXX+bVigTb
3zCMcaN/BP8u/3nj5k70sHNSjfL4qMzf6HLCeO3RLEojA4Olx5fsi740Lb4ed2qI
DtFYepJJbH2IN4OuHmpIXPXel3HPraUA5yG6DFOB4U+qlXC8noLM0MnPCOnIeZdR
8U0hjLGSLRczH3d1ZxmcdBx8mDxIIhGR5A++bqCJ2nP4QXUK1wXZpzJyaRF5zV2q
cnfolLdUA3UHd7opfrtLDKw34rE3aKAHYLCplH+kHIe8TdftPArsWv6tG1XOP2mc
9esWJSqYIaSD858W3SZPjvIjQFjBDsc1yVqedQS25yd4ahjivludQ4EotRVR7Irg
eSAEvrHR8wUOWk9Fs4sXDlCUTImQqVxgIp9iiQvM1ObS1c+nUwczCR5BPZNathlO
pDo6PPur2BYQVE6VWh0arzgis6YpLgW8sdItmRK7Cka3J4RF5jESZ1Q31mkA0n/0
bSghIGggUQCv2+3O3VDa6M7nq0V+T3sg6ktEV0322zx42nKygDrDK+jOhKdWs4Bz
MQSShmFYqLRVZo/wE9NSNl45g5Tsor0wP2o6AFqsVORtiXnc71YFvoqSUBKm/D/r
otymcbb1dtZgLWShcYxql6Ppr4N/IO/NW4GAiBFag6URR1Fl7Szy90aHYudFFGsL
F+D64VjGhHpA6PeIK/TDec7Vny6e7NLBzslp9atM6VqpsEE8J7C1wF4qaPhv66Em
n/eDDD376tWd1a5lIxvI4YG+P8O8cn9EjPPR1cygNYitNvIExRHIdlyz4YDa5ny7
Kc0S285vlb+qmHVKaPXWtcaLj1JNAwua4Prcd7993T9L+JtXN69oS1gKjnDQHcGa
+znTW0P+9SQ/JRMxtsJ/bbzseX3P2SxgwRvILCmM4GNp/C+mw91N+M+Dqfm+XmC6
iuoZoUwhRGti3fMAwSYNrAY9XAgTSfk/iWu/GTVqz7S/2VnWlASiBewhalrNHDc/
knlajUSe+eR7aencS7KNPaqUHBgOC89Fntlv9ASv/N5e4xuZFMr9stzpU5pXRDgO
YF1u3dS0wY3p/u1LXijF7iLeZurIreGR8EW6CCii/uXU0cQajZe/rjaptyKzreJJ
57Kbv4j2bj+EGMqTZk0qVOEhPsk5CAjcjUao6l59AHKdYkUg2pCp1JhRau3Nyd8o
A1Q77BEnBvb4tuLu/Ke7Q5fMOINvr3T8g0KeHhRDYmTDAiqEK1546c04/GDon+sk
+XHWRv9lUF1jSGApAt1Gtgg8uDozjcZ6Y2uCfgsL+E3lG8NqY5Rt4OgFd58KSMvk
w8cjtjNoyVifV1wvgWEnZxoGzjT+uSboHQiXsLuHQiYVqmDW3p/Oc0KLca7jrLzc
dPzZwAVDIkpTi2QRm8sKArtmRbm+SYLxOC9V8Wi1LPdWjo1KiVVcp+mnQ9amGWls
i9Q1HX5iEdMTYfhdIzrjOjvP0m2oilrv6RnuT8LMeE/3j2TCV7ib2tezlhR4jXCv
Bfcg9JTi+zJFoUUPFfI2Jy5anD9fpeimba8F9GgTSq7W6sR5HCQJQQY6CStg33Tm
efTkH08BvZ7gRtV3/sVU93c7MhsVsr4Qcn6/fwjn/9ljBkK+Vh1afZSHqW5wH7dU
G8M0BRUSfX2Fz36UJip0R+/xjJi8OkYUWQEFdZ4V/e7PfzbH25ZXDJZUpbaNWGZO
D8bK//4Ept3on92p5JaVAs8KHM0eYiXi6DvDtnAcgQF+ss/PaetoqKgfBoCaIG47
36u8ZnXWOAoALzhZhNkSVzrwcHEgmZnOzuFgQB8VhRu+ehfsrSSL1loOl8HCGYFP
w3ExSepRocpMwcyW+Egi4iVFAsjAoryShWKKEXKx9LE1P/bC1mrStQsN6AZNOlnM
lQrIB8I65O/T5YZuBtxmajl8ToAQ/B4YGuGfKmEI4k701BNSg1gQ5Y0zdY2wLo9A
I1c5mheVj1V6Lo2bX2Bb4C7wQZKflYZATTBLtW4KOGFbL/h1fuC8Ww0ru+W2o873
QWHmVnatXCTwJnFw78JaWis40/i6VNlVQm2dwjvPnrGkKrtaLC8APToODXJAdnV2
oVIA0r4BGi/2kLS2ivZLye6JVvDKn6TTE5O0LO4fyLC6XYuTbbHRQtKfT/M+WemJ
E8xkW7AknG1KES77Jv35MkZx8mlEs7Qsm2axYXqX+K1K0ZY1VSj931euT+LoNnLd
1vyfPSYPdqqJOL4XOqRR1iWhCqpY0FMYbh9YJcYuKrIPXV7S3VEiUIqdOwd1hVry
wnX5LVHLDkBPyjoYc4+sOdjmLbQOMT8jGb+islI2/QmBzfGih9srf/3vytBvKZ8x
3V4pcBqrpAbC5t1rFUSG2WWlBt7UoTahbj2xVvT+4hWprjccocqFa958jraU/Wd6
031MHNjW9DVc089OFGR0uAbGtX0wB3OiBJRIHpHlHajMdaQxDdJW00DAATsUCh1R
6vRxrahOVvh7F+fBzfSf29luFjW7cveGk/Wke0q2CeHEnVJKeMaODY7FIYR8OABZ
EXU1jsSGsDzciecn4js0TzSz+CxvjeFDZn2qEYZKOUt+WyrGvrhLq+ey38e1rhKg
/H9cMkHJFZgfej/7D780djjoaGytaeKJ8GVtDjEykrYMdxIyeLKMVhTXDQKjvYFI
/0+VAdXGx301nUIlIPCXI7boeT1kPEUG9dJG1ymQusoMLAp4cPineT4ImzG64gBH
l31s3iCh4elOa29Rgw4e6Kagx+FRbC8NkK7wP0y1Qui6MuWyXLf1jWCIUgsO+OE9
KPzCaS1RiiJeg1quz8wWQ4+IMdXAZcfE1/lZwwN30ocDTMS9pETdq3DKxG2rKW0j
tRu+4GaXuwZ17O6893roBRLIWb0/iSkOI6coOhh/fNcMJohLAO4M/iMQfUFTgzu0
ktmeWZt0IEqSMhxgY46/gEQpZDz86Sr85965N/edsBwIj1EZJkmRhS2z7kNJk26Z
VLFPBGVX7VpQdh8+EsVAB3oxrkq+HSJoruXTPbm5P1gfZ17DgmcrlnGMSA342/ic
IuPgdGG4fR2huMQBDti+DRdxpKlijZ2/pcsm138fXdiDbMOkrtGQwKXdfHkD0cme
/32yqyFRcY5MxsLz5EqvxsyStsAbie8CVyUVrVsOaQBBnXGERQ7uhQ+JnTFvptSk
vHJZkuRgU1H30IjEvjSyztKkob45NkJvDS+F5iT/lFNYogyBKlmq4VObeQfx9RbO
BOWUsc8B0xEOsPoTK6nOOcGJzLRAvuDBAbkqg2/8yUvS9ejNRSxRyoSuqBKMBr0X
63f8EVqXvtepFt7FHAZWzSp9MlH1QDvQJKXmKZsblYiDmf89ye/RLL6NHnC3ZdvL
/Xaltf9676BRgffDFxhdf1T49zldcdOOQdPls/Kn0uZEZ/QCl7ww24vgxq0Zl69w
wwgxIEDl8fXmCr5miW2/LUY89fwx/rly2RYzn3motxnpI4uI34RtSofDnLcoQglm
AV0Mi1HMWjP6kGHDqks7koSQcuy2Y5ZDlqzKTyHD8MT7xVdgTv3jUi6TGxDmWU/H
U+D5C973N8owuMBdXgn0lfUjPC4C5L+c0y45xXQJFYelWlekqly+ijiHctZXrRYD
tehiD2plPqKXwVXT1FeH3Nhcba+mGSHW37xauDWYcCmX1oUun9H8f2Kn5H29/hew
/c1n6v0UuM6aO6+Cjbcci7ra+5l8PTgAs6OpGuX/hOHHKLc2zcq9gieu1tAyXtX0
xcnI1xd8Fw2nG1sC5w/Bx3j36s4+WoBCE5uRUXeJRXIrzIY5c455xAVVwBvaICYw
F5QqsAwcjKB0l0b6djv5qILS79FvUzqRGVUsilohgmJROr/lFaLuJ4T2/yfbvIaV
SBrarVlv2/Xff+4R/k+BvRsx4jDcsDXeH2uc7OvH2wP0GEhJS9sl6VIq1bUtq3EK
2A8yWxMqzk5vW1RCjpJxygMz+uYdyIM1NcbU8QrVdC/aZEQrtwaATuh0kB5TdR9n
suFD7dAEET+9z0R6ehbyxYTukNm15D01a2q4CliSxDx2/fgaNRxyoGVsoqGQ2rBo
yRz5TGf7czBSnUJLPtsGwtPLdd/84HNaSxJxTRNRurW2ADT8tOqvdkjWvYPKSrTw
24sQhyeiFOU5vHepkR+I1TAmXP/F6vP9RLQDlXLsz+dfISF23GZHps2vGO4H1q/k
hDnQAeY81j5kkft9Ijy7H13Te4PXpY/ZHH58ETf37Ah71oaHZAei8XL4WXF0kJ/G
yVTx/3lZCKq0lbFDckFo5O+NCCpQ3aMjkH4dS9YgP0wkOv71OAm6KY3n4dVGRNwU
IpefRH+3Hzxvi2lCok5Y7fEr8hNEYfOb/m0MZFAFQe8S+4seOcloQ/Az//rOiNyt
rTP4C6xmj/zNK++vfNIL0aVehflyurzJlQoOw+8up3TIUtcOEgRy9nPVDVKc/xKy
XbWXE6X/vj3XdYNFYKvCZrs6LS6ELzu7W16p1TaR/MSwtVnMCDgNTyTS2K1z4WTa
JTtUoZDjQVl563n+cMSQUNjgRPiPLFu1/H5oweZhvqY1FJ2l215wqZX+LFDD9CrX
InOUDyr+eQiZZpWUA+nYUBHCNmve27dGt63xUyjL46Fnaq4z7df+0VqvL/BrXp9+
Gmv95z58BAKaTpmshdFzHvUSyKLA4Zal7l7/1u2PWT6kYEkaqHf7sLqsIDki6wya
HWkQ0SdFy376Dv859sdNnbNFgZKZogtmHeooHrJhALP6ZFPLSxcwauCOGKNrqrrS
WIRZ4lO/ec6d3xylqfc4xd/OXDu0xMjL27BFBhMHIefjH3UVzGQK9w8iW0L9D+AP
AH8/MrExs6AhEtjUaYJmTIuhwEzqRGx2Ev69wa7ECNYUc71WgcpG5u7QboaXyV+/
IlkybLmRFFnidnTebj4nEcYOJeWWEZOw9wHPrtheX8T0CH3iRuQ1dIa1UXyVf6Vc
HevKboreiZkQXSsuoDE4y8lEEcA1yAbygU25/+0e/c7FA0/9JasshaSv9UGhnH8v
1q87yt0XHrOAkKh1hCvZwfsaA+I578wRJY7XglYKJWibyMAelHEZNvi7/ZaTD5UE
8Commlu8pffqC8BwrNb+beLQWsdkLkAJWCiYr3LXxDf5vzQSWhJ1mRNoPwaJeBEp
4Mm3e4oCv2P29O6G8pfXAsCak+RnTpUYva+gnbWyrdMedZ5knIwFU7osEp2U/k/c
5yMtI8A7A0FKMoQ9brDJIxA2baHZ82NCac3G6NBiJJc245I6+OgB3zgdCR/3rNKs
EdNNPMiGRhgrJvTMM2hKQyiqJMwJh3W3+e2pGVWhhQ6uB3RFz/RumJytGtgKFO3Y
YiGqC9rBUqDLDMJ8eW/n2Mbd97g726QTu0CSkt8ylGTFmumXFnzhABeMTCDO/Nt3
CiGk+XVD1kbltC3BkwoX0rMVcPhsCN4b3PG/Q8BI73qGHBzAb2DyIaXZ4Gn2aG7a
XEucClbIZkvtjuLxmQaw7PPK3FpvJzwyH02Nd6YZgImQ/m6ucIbc3J+95f7lOt6k
rUbzm3KembfuAjNSjTwdtNPcJ63ziT/FADPyHd5alZFHhTSonf2eJTYWvjMTF2dS
Giniamd0fMi4/B30m7KHfkMGJbsYiK5bUp7T3V9mCqChlMaiTsPAlUQAq9DxU0ZE
p3TB7uJcfvD4lJiKfQcSCMw1lrXmhujG9f+EckbWBHN9zaU917Hxb2Zt8DMNQsXU
NtKRD4WlvZS8Bn0RnGtLW4xyk+IiejbGzzuZAignKQgrR+J3W9/11GzgC1vfCpBm
Epn9m/NieI8l1IoD7LZK3cgz/FsROrBfsyyxA5xBhCTxSnxFqiMAoKI5C5mzgagE
BdW6sUR7/KgIedzzL8Ep1O7WSE2B4FoKqzNz6pH9D7lAnsK9a2MIJO1SzN4o2r2f
XRuczjCv33cg5Mu8gE9ejLn4wlTf6z0QZ10h2gUQpbmPljleNClPkNLrRzHe6gqg
dTxcgX9+8WCCbiTLas3bUjAzK5f3fTrDS6PTyj+6GM//u6iZPcci3zy7xHuoiqkH
4OMaKqoY/tKutj+qcbh5QXJeMjEyxK1LcnAbtYHHAWyPXzarehruZYp8rT2hBMg+
5ts78i7E0vnEMTeHV6vFIEhc3CR6holoG5jCgdZj33nJ0HTL7MKl9LZKlFcWFp2P
788Mlg/t1j/Z4mwZIaT74xPUGbRCQpTJMB3A0oywJkGJZXFm83T65mrwhlBMxNKs
Q1A9bHvhBZO8gSWKsSg9sYwjkghysSJnT7C8G5juuX3BtlWmrdgF/11GlDNzABMA
u55PdlILG3/4DB/ZxgLpGTmQQvM8OMyQwSETKPvj2Bxe/vL8YTbxpCgMjZye5cCR
uZ6snYisCP3c81I28xdvhTHxM7D5L2tiFbos5C7hgDrFbd3iK4juGgtrCmjzfJOX
aWylWfSh9Cn00KtPREc75rn2HtLAcDTeFFE+6TWUXIx0DaqGWdWNyoKEZUkVgtOY
wEY6/bY9fPxZCrluk9qxgIZ/tilhIJjCavhBH9Eqatu3CW+U+VUEGS9iHO2E+RrR
tqDQn4MuXJpLtEP304G7XNSWisR+u+IWkO6d5LQ9uZk02e264wdjDfOLU298nCNt
N+fHq+TTaHTwSXT85e5VBTYQCqTG2MEZ8zTou3BH1CG0RbH1r+THQ6heG2JHJId1
E1hUR4a4oBUh2jWJX5CkDAhr6nVe9zelWer0LiTrR5B5j7J8+WbZtdMt9aWYL6js
uYxL0HCOcKmxaR2VKIWq3EMhm5zJcRgAtZ0WBYJIRsZhheE5ZSM94+VWW1Xd97ON
rQf6iN7ro2E/NTO3mF3siIra1iie8KClERjZlmpF7Fekrd6EL2QL1gHltKK7xSlc
WA2nZK9lgJeftf9sEB5qRvA0Ype2aPl+H8D3OudlV4nIvr4N8ZXG57fcr7ShBX7T
FKwWTKXZw7IHkSyXrvAIxnzB7HwVQiqofSdXH/fOrWaLqLitcA27AqjS8qHzEtKF
8A1B567iJnSmg6kmcT9s04gmKRjojEso6WeIExyXkPMy6FENKop+0KSgKe2iIrbk
qViQRjqjgT4sommEN6AqYfacdHs6OAB2eTvs/O6zPpwQAqrPbTmil3orrmp6IErA
8Ny4hlTZLze7ANrW4EwPmNWRDxNTlphXdPMkK4+Zorqfh99Gs2Xs3vfbtSRII9GN
wXLSvzbn+1dXc9jV18uzIiY0LbhpRTTEakC9PVoLa9j5iWH+vaQySTcuZNnz9RtR
s/D63krFa/QYoyWvyRaS7/sjIrQnuaGoGGFEe+GfQ1LyyqWnxe0dHWYGyLPlcvJB
5F3YJUBEAPSMaJdhmmRpmLuukYfEx68wFxgnu3qh6rvvzyUpXm8nV+HH/4i/72Tg
kBVFb1dbnQ8G1ODuAvyumozF+QHO7FkOwUa/+6SD7+AmwovOyS8KgY+HdIZ0KeVk
N6F4UVDB8IdT9OVtDLH9dc2ZTJmTlELI23rW1ijbKdvt3Rk8mFJNQjbBiJTgemqX
mmWwNbpYuvlM1ha7zEmperaMfK+UhgEZUth1Bm1GDGx6FREuaTgqaW2tlywwCMVi
utY6fIFmbambU4+saKE24jR7Ekqu9n84vlGSjmra/YnGTxOFup3OipPYPKcad7ZS
FZMUyMCdu+qV5S0HLiwj3hASinLB9E4tUPJM+i7vNAn2OM2+Uh1ynjoYo+Z288Nd
vb1jkZq9zQTrW34+BKTO2BkDFJSHdtmYeCAPWg/CeFNoA2ayV9nhh3qfuG2Kfj2s
73DuYS38l+ZKV3cubQDnrBnXO+AizTWAuaiueWI9KDGh1DMYN/IfPkmkt6vB79bm
juMt2nT8N9Q3kvfZ2YOVxT8AsXRJEuvLL0ITvfHmczo0JPshN+uR3GO0w7xZ1gFi
gzdlxiZNDC8SjTJv+lruKmL73EOgmxY4smYkoPoN6/8sWfI9i1uTdeO4Fx25QTVD
TjZijHx/mC6zg4yppLcitcW4FDLWsW/8LvS+ydx4XckG9tcJ335fJI6hpYRTpzD7
DJQ9+eiPPjztt2Fed/eakY3t8N0p4EUqNrZUt+ilVxwwGUJxh1Xj+rwQXnGLEfN6
5kFEaK3O4qBjHyG/Ad9+VXIcfZPq97W+eaUSAIchoWSEjuCDhdLxjT59vmQm7e0n
JDiYbNj+QDAM03faVGNHG0k6cRRybYSLvxziYXE3vWoUdqOZAAzMMgDiz+g69G+I
iA2+Q4+zTUMXJBXRu7tbAxKKccxCBIytJrQXyApWRGuIwyv63p1MS/XJgfZVoJVh
mLgTKAqTLweb7xqmjkwFt67XtBLkXZM55VZvkr71VIQY7HTam1xWwO+4+WhhjNbb
+MYsm9PpQg6P8miKah77fpXsoN2z9UQnxhJuAZRA1njc91n1KPlPXUGGtXau6Stl
88J17nSgUnElazrAwvKGzGh51Xo3xUQXLDbZIdSCDaDki5B4gcGVcVA+RX1u4Gu7
i+LW2jMS6GdtOQTVPsLv30Q9Vh9QDmusumi6Ygy5mPNdUX2aQwIjqq0SqHVqtemg
lkaTgQjyGcW/X4RcrN6dgs1GtKU+c3U9myfNiOz+Jp+SNj7Z2QSvto1/3TkJtgkE
NZPWwcFYznpSORRgAstxwu5Hddxf+URe6xNhvO6umaoH/8oew+J/geAEs0XuRyTO
Rd2GIOrJigOvJdfolGIlbmYjYoB7uVxk0H309ax+cuVgxATkdgJ2x6Q4IAs5isa/
pupcWB60cEUN+X8XmYTchiVzHO9omTWVxsSEBRd9Af3ZK5/lVSxHwW5dG6rm7R8r
ljMytwtf4XBDWpgSaD3NJqKb4wgn/ajPQQ+wuWk35Zn/xflpP2W9Kg5aCYUZk1en
GsXvm/jlzUZdXdEnJf5S7eqpJ4wJcRCb0jE/erfCoyvdpkRwyJziCc1y4m+9LRJO
09r+bjrrr+4s6huif9IX/1aT6H+UFQQ8iYsSumE9fMruEBIytnRxSZY26K0dybTe
pVMzTI7loYVBWCvhM68eIAiHXbbRW3bAwm8ou8CeiEAXW8ZSiuRlhrK/J2LIDvRO
9OSGwBQkI1k3aaVGj4gwo4wHmbLSNeSXyW1ZOF+q1zmFrtfQoLPdIYNfAFbq6Rm4
Wwmtig/H3Ds0OItVtvUhUoDApLT7gKP4y3imhv5hc12bj6UGHxn1Yp0mxV9NPGEh
Xi0PpzKoXDR8xAhHNr+9WyzyVn1KmWru9ydT12TyQDwX+xbNpYodtgy55oOpe+nw
tiw2iTFkU45/+aVw/5mjIOWcC9B8pxqYgjVAGxhE8sbmL2c1mWcKblkAeV6T+TQv
/eznLzmOj31Ma3Q5ylwQzVk8vVocCnrzPTbzr2z5KX81qDhatLQnm3xJLgJhPaYc
3ES7VtWjtFUsw0gVRYbJeCm8KxSbK14aMM/D0+/cnQ5c/0yiWqNf7dBxuC8BeoRb
C35MCOM+p9sP1B10D9JOGyYD5Ls8QXdlTlEHB9rz39H0iP0J4mul5+gatjjA+68G
pq3Q1KKrA3dJ7OPtdYA4X27+7q22PgVy8Ya7ScHWKJl6kUbKL109gxtfE7rKx/7A
xArqUS0hUYt+7gLEoRj8rNWE50NXFO1lg8gx3/hzgRVP/9SlEaSNYXULR/zjVNYL
TzTwQdmnPJFTwSxdEmwMUPZShb5G+5S9iwF5/htUlh9OP4CadFbojmF9dRMv7+db
fmEeJpKcAUDeTYz6YD2VuXHBCDH/G8On/91gzeNtsWWyXLXOkpC+Wp0esZdxzrDk
+D1Ioy1iC7Vz5Dy2Apq6K6laL51+y+wGUuIYuiJc9ccHYUKLIfh09ETL2iUBncIq
0vE43IJhZNbesT5n03rV6IoVUnwmm8LiPXSa84jXgOlN6zelJ0r6q26TQE+vpur4
sMjlC075uL80dk20oZ/WAwp/WHNtTu5qqW8kFFkh/00kDBgZ756PpnoXYRCuIBCd
5TGBio/skmUnUhhGx9O/nB5eDT9Os/u9gp7paSyc0nzukQvson9IV4gfs5bqoFiF
rkFSbc5HUAecLzzxEC/5s+x0zseCWS9EH68PCvWr0LewSUbH4LfgRkZ//yWI5NaZ
ctkJ02iG/BmCtL0PNsv08q9Bf3f7wkKwG75b2hfAxm9nICsi850IJGdfzN0nXBYp
g9nBQ4MTMec2z0dMlu0HSgZp0IYtHcU3PT3GChCC+TLWbc0S/tdy1xj7vbQtKuqV
jYiFDpTGD2F6FHgOSLjsIRz53HFwGx1RN2ad8BC6nUbRcM5Mr/vm4Co+VniA8foj
/+GqBmVoYMacFgcqSpbxFPJm04Tst5/PublhfqEqfZf44iJWph2ktQf9IZwBMPw8
aGcdHJS6d8HfQMZ3vSDwJ8vsyVHi0vtEtoLSpu+8+GvQLQI3DESJGmEEAezAJLVJ
udebMw92IHaf57P3UUJf52u8+y+Gre4LAlwSJSNmz/5wn8uLOnUhZzG1r23gtYcH
8FCvSeOkJfxGbeucGik3eVTys0lSx5dfN7K+Awgqfuu4P9uYMluZrWM7y6l3Xwmv
F1kN1pOr2UR8NrsOPX4y436JgyaiwZl3jKRLmdrmgDQFQrca9dC8kfSGG7c0ieDp
SppR/j+7mtVVa8oW0bS5Aqjz9p/CeIcxygKwmw7Y3BRY16NkfjNoG1dHjSlWxKRH
w3Kg7fd/o8umdvwdxfk92H9WGhyvCfM4yX77sgqdO4iKF+ZHx7anqNGf/C1x5D2F
n+bLno00ShVk+RbkTdH5jGomcRGt7glgGSHv5KutsFAZEK6y6y0cRcVrtuE8UcOi
4+aGCshKzxyHyPTvZruSIfAoB/HgqKsxonJjLcvadEAPTDVaxRunuis6eSKQwkEV
J1uXicfSkEsB6D7MmagYPJEi0qbG7DGobTjMQeRfQSSqO9y7qjJS7VqCaEdpLc3J
DAnDku1y4vhatnTQKMV3eARmJJytQi6711n49/CnEm4Z3eW8QWgx3aiJB6BN0XG9
ZGBDrsT9fdH2/QDhDxu+i1Bke9bj/ERJLMZxxR0oQ0u/oQBKA1gUgfe0Ibt4BAtD
J5thQiJ5OgAvB6BCLlF0h3eRM/nG0pHqSNf0Yj3VHmac+NfIDzDGhYqSYBrTYZmN
YeQmZVb9rprWGNb11xH4oqEZbNmaJvxcArmA8o+lY0UGH7VPBnwj1EOaWW8PO5u6
LVMw5WorYUhKs455IB01g4JxxEPE9VaLNbivt4s34SGGL8oh0xh1jqtEDBQlO1wF
+WVPu47qlvgRpC+nSG3uFQjBMcad2qoRyx05ubnA1eSvcDsopX7yuxxOz7DzUeTz
4xGqJgDbYxBG263ZoktElPqkyqhNd5sFCGyVG/jPZTPsh9c+lTVLY9Z/xtG+Q9WA
YFDc3lJHXuLlW+ChbI44GcDQcnc7O7BNWvpTAdnZ2gMhSXZUy+kJyPvTUCd+T3Gi
2uY2JP8RipHsFzs4WDOPtnV4sw3UDJTooiNC8+5GmxEAac4GQtjjdCMIPVh4cCiT
tNKD4YJVCxyEEhOrKyVgTlnkxxbBI0gpahmpxq1nNmnyLItIwah6t4dlwl1M9yKn
B8c9mrFp/ckTcid4aENO1D/yYenkPD5YcPIFHUkMwjXc/ZM6MnQWXkLpS2H/HUdP
PhkryOu5hTp7e7Ha433RSkchSdj6LIppKnxym1gT6RnPcB1HqDFote8JlzW8NGGP
zWj3t1aUt/NfSrabr56yBALr/SjRXy1aOn4KuumcGD68eV54ZCDvQiYjm4ZyPdYk
B9RmIIT3dakU3omOj/rolrz7CW3XVx3i9Y6ayIitRO0Wg2kxEgs2NbrKjLRQuML4
uohxn4Xov38zJ1A37Bfb/AIqfxipmxyRM1U1/mTblYgMJyNh4VDgrBwB42ETMOnR
LhhJmCvX+858y4PhhI9sXqie7DAv+RTJk6P/e7fL9DNzlBztsZjewA+NaZH/La7H
0tOzokEb077X/Ws5IBqnmg0r1AegzRiuIoew4ymvvV+7JbYI7Ww2MCharUh0MGck
3Du1WW1Zug83XReiW3K60c6TuXucQRh1CkAHOnqBmvmurEeIAPZabe4wpse5iS/l
8Y2jYOs7hQ+3cuLERzLZSs8OT93u2sKSJdyxvIv03OHxvr7IfQjttOmYy7G1mnDR
2K72GIqHgbIaFDMkUIRk+3lsjTejCti4G6gHrXQ4Yqw/jfGsFyVw6vZ+c1/qSjPd
H2VOXxvI1N8j54j4i+T+7HLclASnIMK9DPziEnYu5rMmgffP6HLHM74NA1lwD2yl
0R8zvLOPDBzsqdplu6PYPFP5kzEubsBDEKWDvuO/40LLa3/kenuud7Wx/9e/9cFm
45GkKe/g+ufno/FLNAiyL+ZoWPB3OtVkOoGStlvceqdUw4/2LLZkf5oS+SpQp5S6
nfXpr8wUY5T5UZJF51uurtVBjRvpuNmMd3wjgekCLE2t3JdoH6VOXKTW3gsZSWG0
5276cUxmTKaMJDiphTJQ92Kw9SnYJdapE1nM1FmpByhcdncCc3J7Rer4Ym3ta4St
XVUrshuz8PJ+D1KZZd30os/OBoI5IBv1dHdcEmx8FA5JJWAXFvJwuaIe+OOqfKEA
XkDXC81e9DN/9V8sqWzAaLKY6YwaN7jM6VZloxtPiAO9nN7Nw2WDmTi+5VmcSHWW
XJsJhvhaIXUzKcqs9UeHQYStT/sETHOL1ghzB6krkrk=
`pragma protect end_protected
