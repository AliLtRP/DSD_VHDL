// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
A//PZNm4WauqJDA5OnNykZqWrjE3FIK9Wdoliwmw7Bp8Y1+c0duzV7980sLAnqZ1itCiy1jK+KRf
fMbbYaXVLQf7yk0ItFd+lfYs31Q09+mWhAi8BV6l7/C0tx8+Nn+FZr9eI2OkPJkAlwU7VcJWu9n7
Qdi3RPcgn2D5jgNVxMMz9sX7BEdTVF2pzC+IwxTsyVB6hb4MoW/CGIFOHIwoHdt8xPjqNpKEaKDj
7ZvdCriwM5ruz9laJpb6HHiA+wj+2f3H+uZorTLbR/YLxKVe9K1nNYz/K8RtGQX9co752r5BHA0X
dDRDULHesWtZ/7MF/7mqQsp9o4IlDLSHJ3yEOQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
dg2IW43nQqbt7LdAzgh2/JCkzyqxvE5Rt99wXT8Zyv6Pv0S/HayNyVnZg3iwiaSCzhqpE3G5R39Z
TwdLbcRdD0oVIEC70+g7cI1H5TmX7k9gYiFjqXfvYj74vK7h+L5zcfttRaDK+8dAVz2VWJhKoSRX
DMUPzdr0kVUcD9DWlVUODONCurcRHh+7ybGIR8apg223gtoZ+FqJ7qznBOcglNw1GjHTot15E5fS
twY/9kQqroVmwFdT6sIg0ZtSwwyxOyVYCckTxwd3VchHGiCWlJzl+Fqx4dY8EjNvg2szt8xamFMc
LBzrzSbqSLILmTW1vfuQY3U6kf8PgG4KckGuUp4N5JLuQrzdMlxifhLAclpYOdtlUl+KV7I/FIIt
luHTcP3RPpHGnmAEKB1jBgdCj7N9enk4yoOXrZN/JUdFy93pdutorGS/Pk6dWmxwGQHKzpOZCooy
0HwA4grn91CETChkqOndWAxOzVTjQGb7lMZAnttQMPFGFHWQF5qKiIcQWzqgzZxP6pHzjXStRJhX
XQVcXcLXMOKhq2ns7HIAVHmhuRVYgjH/UueReolE04/CKjydWUts9728NyDRO5NAdTLGUU0caICP
0NZaT4WazkL6dSwDSc66q1cRVXQGUNv4b5DUsjN81zAvAkUrkTRVjFFRvjSxaSSQnSwWvFkt5yVN
uMndwkvU9CqS61PJe9mt4WAwhfz//sDwrrc5vzi/JmC+K1nYIho8RCsmVMCDoZ6xdRKiA6vD0CkJ
ZMjl0aFxUgV/Eij+tkgRIh7S0mXrMo2YEt/TgEHQwGvECJafIC0XrEbqGIymGSoMqko0oMogQmMp
C6jRuRpmulxnVhZU3R8lPg4elM14Cx8ObR7PMKh2wzfql9Ba+ndelE0FojUS+VofCPFIV4XKOkj3
QOTahNH6/2ClemkTWC/B3D3oIHTYcpO/Xychpr8ME2Rz9KTjnkBcREg87S47+PojhQXW32L3hm+E
UiBbi9StloPyGncaks4oMA0XE+QEfqkwKayVoSUtxNb2VdFQxeQB59vfazRd6Gr9a9wRnU8Ro8+X
G/39DwwvI/iaa8w6dijd82kPCZc++qnYt8prynJtgYGx1EDwGUCGQ8kRix0Ky+p4TfC3/RjyJGk/
kwl062cbU6nssEv8+WH6RgEEHLiQp+eS5qzVb4KWHINvVMH0CsjcUMwwSkbnNOrjxxwoGWNYYlHZ
wYOxTQZdrovMhlGb/vMOxu6NWvLbW5GZWTIvQ3SJI2eyJEpOY9leYTwelTeJf/3QwqxcuSBnT9eZ
Rw9DeXWsUi/pOuUtEgKR63etEl5lSTijmO0n6jPc7hAsoQGnCkVaptPi8iXtqG1mUI/s4qFr9EBZ
GPra/WlZOixSy2bZWsHuSxs8mx5xrg2Bt3MrD8RP/pjFOBzzUHK1BjgGS4r4lqpb04xXxTy3XjiH
fnHIqB4tL6jqzCDNpI5nJ9Qk/AMmxK2LHLFCN2qd3E+BSuVFjZsH3M1puMnYSRV79Ql/XhoMPmos
gbeGvwSQQI0LU5uboagbizhwWlVCguJFF4V2c7fipNKS2uIJiGP2aLs8Vaq4cYRNVTkWVuBeXWWH
WrjscQNpLxuU969eQRlhKx4JiMGBwnST4s5yzX9S49RQW/n13Z2OT53nBCZ0TkQG+B8n7jdvEOpl
h6S3AqsAhcLJrgamIB/J8tZlxf1zoZmXhsv4AUMojNPdO4h65JoL1GEkPz/fCG8OvyxBv0AA/tN1
F4BoM9brchHY/aC7dmQ5mV7q3Q7IEPGVaHZEbY48kFkD8La1iK6gOritHcRJ4dLaWBHU5pFy2cek
JX9DlTkQEhYxczBRWZRvKPI9moBnj1zPIlx7nF21+DMSEDAeC7XpmYAsBPg6XKfNRuTEGsRtKwZu
dBzd7VSxOxO0WCcvZUPTrUTmTBtf8MpIYZme7NS5nAwXP9mSX4xtZcBjIL8Eo0qU7RRvV3d30BfO
5knoSQZP266jhnNljqUEWRTsZE6OtPnwHn+7KttOs83JkYUqc87A172NdxvfMb3nhmLvkPF3Hpu4
4ecu2nzrcgMzgybZu9e4wnW52jzqxIuusA5G8r6BarJGXQxv9OJCHzYtoSA0+AptdYKtkpm7Lj9d
PEGVOwzpkgdFgAoqmGnU0N5kIVaS8PWZbwOtkmClitHqQZqZyPZfM9EF1Dxgkgu5PzqdKRYs7guh
F8rc0znPT+8rWHjjDOTMel3nQrsbcVbTKlCeTnJZWY2pC2hKpUxb1a0uryqMM6W/g97bF44qc91t
vAgRZc+ni8fPvAtJsqc2ROYkk72DIP4okkBoDvYIsQ3mg8/qIiMWspoq647r0x0XAQcpQ3OvQ+3I
wPg0vM4sh0hr6nQQISV3Zbsq42TJHaPKsUGKeEPJZXqXo09VvZ7Gd7CxDSmw5RnM0KPAU8POvmxO
40+vl0B6ZbXBeLFOYIFEcE+VjdJSlVeMW4JzbidI1EWpoMbyF3v91eHG2ayzPRg5nUjqaPiOuu1t
zdwf6bFn+q9UStOQoyR8jUl4+3XZbY+F3K7cRzv813UrBZUxwmN5QfGUDVQgz/GZ3044euwwn1e+
4obYHkzTGff78SASeF89ILhCqOq0ZRdFGzvubFUz8KmS83fOJiaiTYfk/Kv8+2zlmT9OPxQQ7vZj
4KcWZ38yyLKgyYtENxRdDRTSeaW4kl96mVsS6UFWisF2am+4ZfViLGl5ciuEehFIIfhipt13Bd4X
Sp42vToh5qaDxyByHybMCkDp3lhjWyJjP29+vsNh4xH7G7WiQGK5MSzTUUPxhk8byJYq1nRim2h6
tXGJOFkjuh7SWdk4ZEnqScCIZIZWseDrtBZKXXchwofxwYYngSnsU1pU+fntz+dFE3xyr9SWN9ty
AD/jAX/t+y6zPQtUDbz8sr2fnuzdou0vfYNnnn7Acbg/jGxqQNaIoR+2O/ARoBnRrkJN7Se5iS6B
p1xdyxYV0WGnqr8rXyuxM3pctFL/48PE9YeGZ3NTMaCF9cPTC8M0SOMfO6N+4NVMQk1QMyJwWxfq
4YS21S38K3fC87e3ZjFJlnL7Ns1tVYM5w3iQBPXbhEjbl3/JYNWAtke7Xr9BtMUKYSNpnT0MYMzF
ocQ2j6ysY8e14Gjif9vXhtlnTE+H227qeLCQdmuB9G0rfBHcdZyAZhUkfRAVgvI87Lh1WE8DaeQo
aaD3DKDyLn861yvswLP5KxAk7C8SjWV5Lrg8wsor04cBwAKar40tHvNoGJrZmOCWDczCH8E8E9cd
HRXaFhK8QDBtqlNKhnXxEVy8yVNLHhwTjUcmm2nb5S8ql1Ch/tNzp8z6g2vRCflRA8rWyqvVDahF
zNT0+nof+XBRc1w/qb26hJcB85e4me9k5E5xrKlIoCIi5bd9MUXSE7meopcf81xo3lX7RqOqBu45
XBMTodWVMDMtlot7FzzBTNkTUyhM5DKQN1c8g56bCdHyZaEpFBbYGXjf4zesTShLSVrMRrT7c23h
KfGX8lyc64+lt8PJJ6NmcKRmnWbI2ObDxaNedguUFSccZsaPjhswHdsYet2QwWISKry+2sfc7XA6
t2pTMIX0BrsimV5Q+Xf1j/2vIkkEqgixvEhvoseXo7nftUnmpmfdwquCxomAUGKR7D5otc1ePTjc
+IoMVK//s9yuf1tyQiAn+BUBlfbJqtXGTc7iKw4LKRp3e0ujz8EMdQ4AS4aaZHeJcyfibjX3ZY+c
7IX8sE7VgQ2wM6acylbXSCGtgVlvp3pbhQztRH1zTTTePZKuFN+qr3/p+7zFCLOUYDb20ri5RNIZ
UAiMy0CCwJBRSl5NCe8Nl1Lpw3ve1LxPv4HqbLBJaQAAM8XYn/NJkUDFwSciSCppZ/flhoekKHXK
d0T5/nhPLipO8Eco+H9+7FMXzWnZhn/1VDEYDamPZ9tKYCPaGq6sy56KiUj5rL8GBNEVc6iueomu
s7dFqrMes5AW1w9354bU1Qw3zM6sFDmKSB+3UMQIhNmvegszei6SpXUZOeMQaegCCnZP7ieR2EZS
tCpYxY6yVOVy0fEDoilNWWy5Ej+cjdy+TbmWi2qanSqGPLqRkReuhjSddF0MPAwCRS48OW2NmyKx
IBE1xu4ppP+cUStjnUL0VGHjF0T6wlNkmyyYaXQoFsXUFHa9OYpk4MYbeloyL6HVtcCYcmIk/9t7
cpGASShrwWlC+Gu0wcG6KbZT+Ad6I6O8aLx0BzBrYxr5y1AM/CBjY4924pqsSFST9DLz9WgQgq9f
dajGWoRy8OC7yqPSnMfTk3Eu/Jxjcs7+yjRK8aXxfLT8hYmbZuWte6y1Y7oVmTczpEhnKQGQyoj4
qqMB/jh7wXwuBSs0HBydmAnHxLCmmDVmGN+qIdVVraoSa0CKvbeX5OuzDhNqXcJ1KIvTFiMD3xrP
3WYETKUWOpSRib8MT8vDTSIT1KDghWaxOsQ9HwtdumkKaUP1ZBvd5d44EB3G5NEmY3sidrgwa13E
naBAzLNWnms4DIAvTc+nZ1RDQtV2PlDfm2Tc87eR70EFQMTdVp2EHjVP1VE2XyJHBx3z42a+ASXv
zIDQb9YBoH9Tjo7QQqoZqcMe3TI5QKL6eK8Amk389TNCopwCIAoTeT4g6IeNuHS6pKqeprOccq7T
0Juf20tGz7ZUe9hf6cjJ711rO2o3386nGuVYnRDB2ImbfVnrrOQmRBSp6qLDpxqa6lqAkMhDo6v9
FrBc3c8oJUYRzo4DXOKybLTCAI1eyNGYDeVFqAGRMLRcLrk0D3f/ylTEwXQbNThGulTJioP9S7Hr
bcliSV/rp1DRzcLf/ve1Iz1r3O67R0DUSN4LfymttR57ug1XhdY7XsLY1PK8ERhZ9lRFFpMrU5lj
rUhzb4JrKk0eIrAcw0BgXLKx40d+8hv26tc4hmZjrT0oaWG/yamCrSLzZcZK6eUszBW+XAOmNjz4
SH5Z9bM6/ZbHk1qxgFilx9sl9qFK5HuF5kgnxwErVaY5nyk6nS5IVaipJVeWdVfQmrQC4wEizvNN
JLIDaZtSFRHvEEfWkvqDWMzUVM4HL37Nnb+RgKNAX3qFSJJCCsN4e9M6KZUmoMqzueixHgHLdI/Y
NDEWghYg5vCzviZf5QTL9qTXJ+QXd0f6R2YV4uhCH9LwscZpMzQ1cOxZuHAjzKJjwJbRXc1E8Wu0
WSpn2SbhOE16dXCVpQn9TvDH6i0f+FHjd/8fOtoKC4EQzOIxc5WUA0iIcx1j+3hlEfROFSrOfMVK
cNoC/nYr6giENo0E9XsSSOn4p+YinGiR3ElWqgcl4O0cfi8J9BgeR0S5CzI0Gtq5Qgu5IJIhwph4
F2P38X1R3EIb9/TQBQDv/wG1YDn18lUDdyzSc2wmogD2GdELf9l/xQMppQNkf1Y3ncUewE9tNi2a
yjGHtZ4Cg+rsLGa99DaXDDg17qUS2v2i1afTIP45SJkruIVA9pfuAWQsg34hYqk7gjdNZXaFNDkx
0B0gpa+iszjBUOTKYffK70HLPCKmsMdTgyT8y2sthKlNNyILlUYm64BuUOapRCVjQFJUHUaICDnj
joBFIHas1soB1qwcd1grUiinz6qD/bIhMUlvj0S6vMmUDQKb7GTjKBgVOZ9oJcNaZpNkE8ZJxYKh
VhjgrCBzAfcHElcJGE1VSgtEwNWbwtY1WrZ03P73ueomE2xckCQNz+Gyw0Y7Y8kQGbaHg+VwtQWV
DoHL3SBNxVsaf3RHEmJLmE8y5jnUZoIQzSlLXLzo8m1Y1PSqZUBt3Km04zupcLwhxPZRY+6Kgpb2
Yhgp6QEIcNVSp6UXjlD8IOrShDxdvpYFCOCCmHuZpDr9DX1YppOo7bE3E4NyqunoGxpWAblNue04
l5dtdnrX7aSNLTYtR3W08CIh/6MTBVd+JH5CZnbvR9dTyPo9CT3raMiVWPmCqNEDGnYW4b4341oJ
B0pFZZtctCPbPVsl0NeWbka57VApL7VED6pnjJFIcE/vFYEyD6cWFz+Fi36GEXYSj1/PmKB/9UIq
L6W8TtKqH9DKS3XRaSXIbaIO3ROfh0/9qi9MphsEt6wF6osVkj8z9VAPnDs6ldY+ZwEzFEy2zFgl
Se/BLW6E8dKyvYSLoRZRiHLuDCP9wbum46W2pJin0d37G+4W1g/2nwm5dnP2/lCifWmbFqbXOoEo
6b5BuCjk14OhMCMIwWxTLJ0vWx2XjArhN42tM5f09qcaaLW3PCJALJU9ZBevu5JNcAAk67jc/mie
JtcsrcVwCewDRxm2D+qsN9Q8qTZp1d3rqJcXB2tRM5HYV5JoeYzxd8dobfcs/UoKEDSy+6lVtDY1
BxL4HdrsCuF01zfFnRT6qmgLQV6u1m4XI+Tg+GT7z9/+IWKJK2cxRgnLMuCFH1YAyLArbm//70Lx
x7uGUbdxAoBUeOVEJgAXgqfIwIWhvBe6zWQVzykdfCktUW/aGtKi1Zou/T5kOid4RNieLvHqWb+V
BkiNBoNeR0aGqVzBausTtBPL7SHyiBhcrV0bQU8EA+fMgZRQTA1aoW/NIslWD6/NTvPfMVp1S9H2
+aLtPDkypTOm6+USFA+DavPr9TA8fiGvvRI0B/yHnCjGFn6fNW13XMj1WPInIFMrP7Bfe53BC3Nh
fGDh8lUr63NB6YojD8o1gkf8nBPZ6WgKppx3MmDnXvpya67aVctON6tIZjTc3U/HuA7uphCw8h0M
JorVyEc1pHutjODV36tS/O6xWBcYX4vVTuuos8pKYqnDNIr30kQSyrliDRqmqiQqdvcUDBeGovN6
7HtF8iSqbXjeNEbcNrbFcfalfydsDkVYX14qDxI+Y9bfp+TVP7li/OFv8FA8SclbLLXN67QCqW7v
lRyBpxo6phMMjqaejoO7YqH9cvuXQU52sbR/BxvoqHogFNaWxsVG2IB2i65nwEKCzbeWkR324Bj5
FoWr6+P4kvoEsSxM95xFj6WbD48bqaUEzRFruAfKdppHd50zv8G6QCTdfPgA4LyR0/F7dgH1lAWD
Cjn5QhgIiWhFCO4NxdpdSpwPrlahey1ih56rZ3IEuJdVhrp9EHiwzZpVhcpGh9NTzRLZw/G17V6Z
+GdXQOeHHynC8UGV1klf5ZGZPEcNentEly7B4DrcZYx9pXcQ+rHaaZ+q8ktngxmiC0jVlxGIKLgF
5iYoQcCFhZnLYHemcTy0k4R1PisLs7+aY2OjcqOnOyA6peuqglpMkw/OHZevcp+GDqK5gbrxIoVB
icwa5s53TiqZSUnVaHaoue5tQ+nilaK5tP+QSyZbYmg7dR+MnEZUhGMnAwUV6tckYPndFFiwW7pS
Dc8ZIubTQzm3MgZPlZ8Cn1roQFGzKXSh4MSktKs/CqTLSZ71pPkWZDqIbcmRruXBq4c6fy5wZFZj
F8v/xVgx+Zcrd1iMat9FCzHK17uTVUfDjC+ZLNib/9Cb0bCyOJCjaJPBuinoYdawaeLuRvuO2VYn
tWNDNzBnJU+MRfwp8x2rrfXGSg2VtezIH8xcG2trGZ7O7YVbhMMOVAFQf8o2JjyOjFS4VqLPQdbj
uIVjnBMsXEsxxkHWLhTSnt6AHys4ZR262lZ+vbIa+PmP8dGMIi2kGzt90U3Y9v5li8cldGjQiqz+
uL6OIgwoo/a+n9n/QRn9mpeo5RLza97Bf3cOxhbdBFCRwfYMmouhvTGcOTB6rHZLaTdJT0HI6chK
znaKTL4IaroqscQywTRDvqqoPWIWGDLlfjxcXI42e77w2LEG5nctuLQnHvi2UKe8mohuLWlT0G/X
Qxj6Ubeub2A/YifeUzsoMYMKdMwovUKjc48uipso0ZZ14VmzSv/5G81dm5U2RQxlkK2Yu+CQcmu5
ZdBvOv+gQcAPZtSHeDRDoQI+/zHNPnDT4m8NyGdydgDwywId55RTP5qLqlNo/QddKuMWqISUoKAx
uezSNZdbbpb4aR8I/2Z0Ws03pazc5vBGXOhGZSjXlPCxAQ+gshtcbPoaGbRHCjyh5cFa6LOUCCPp
L/eYMPdGVesI04IEJLjY8faaUjCA9r2661hl4J9eU3dmJtpRL89sdCuCMXumAOu+nmFNyeMqwPDK
/6pVy55HTPhmsQJRGpQASK5Ndysypc3+LFtE/SJqK7pFNW+AZO8jHa0SoJU5jOBWbvCYnQGJTtnd
POTXCdLZSpF6d69zuodueHxCPuQBtBYDdkRHzD9TCEztsSB9cLKt+mRl191zpxWHQNqkMHThkWLE
kFvr6blBXJp1yoveWnhZxm2yMA4MwRD8Sk6rpe7FBcfhuPWqtwjQcVMIFW+kSW3UB8n5Tm/KPn09
k7XgSHIZd6B/FgE+iunFATXRZQ9YHmKzXMU+cogMzNuLgWZKcOxyW/TXLDGdpesuT3wbVn1gOepg
PpyRUCehrpwGRAIBVjAWXc6lNzAFSdjB+hVsfidc5eXxSHtiDaBmWhc6rqXcCLkQrOUTrGKaOQRY
uEnupAHn8YusRFW+99Wc9/+GQIeuAtAB0RY93XHTGDEvwx31P6lennS23VI/mnH72B1bs3QVrhw5
H3MZd2QlH/OAX4jkxZm9joLQbpCRMnl4t6UZHuYbgtGmIBP0ID8q5GTO+vqK/gnatkFZXpdzOXxK
fBNNaQmioEm+dqqD/uXszha4Ev2YDtgM5xzQyvyMQ2CC5NKqJfQVG5kdPiJcsoRusNCMelyK3G57
coX3WZsrHBnBnEIB8sEFDBoQjq4ieE92jH+nBJejJ+jVoL4Uqgpu4mEG/pnmLUpEKuWWFCQamyaS
BO3R6JLxsNeCd0+SZDsyzgkmpv/5c3L4W/J91okDUD98erYrs36H42cKzCnR6MVs2/7LZADCEm/A
zher/IAr7sT/3EfDnIXJnxTkuZl6Gooty8cWhizJPZdYlNkZk59ifEAnU16XTJYMDdeXZ+bEgyM2
KDmPumCKTqT8M4uUoEl0prJcfQYfr+1871dTexHYu1FfzhwtuUXlgtA7aMbCyqYUr/SLW1Gb7g3B
th/v27vkjIwIS6cRzZ6pI9h8DSpl2Nh7PzQj06Cry/d1x3KGOifeauscewQC8NsAFvpzjCtWddJa
zXQ7KkJmGPeYzl8SgSllIrfjt8G3UM5Rr5PdwiLH0bTGBkKp6mYrlfPZXRoTrUh4K+iaPSIk86c5
Xnq0GnGMqwvJkpS8Ltd+EQPfNtrADJCwEakikpZSe6P3/PEUitaF5Kr+BcaGvsWve08sTpo5kFrJ
b7mNEY/gdQ/mi+VWAo1ep9/+gItd/z3r11Pd4d4yPXQNpmW7TPqYkwlV3lFdtQsnLnLQdZ0hIRCn
sH4MmxUI79X/Xi7O7pmEw+NtyxEZ+eqn/V/00DsgEc6/iAoKyyjDiiJG467iWczT69NGlN/uSQEl
Uzi4cwRWsUYGkAjXcOvDCa9zeRFhzYwqLqAgI9zSjdkgV3RD8KpafIDrKFilEk+Pkc81jplvJ2hv
WxGAcUerW3H6lHjhaE7NTa1kq1JmNg4KfR1SWhxDhhpnCIfIly8mzrSreKf1/BTbGEvY4PKQlFnO
kBVOUvJJ44R784+ekcuU6aPcvA/nj+SKhPwGbu6PCeFpN5OSGxziPvTgT8EfXum0WhF6WGby8ll+
RAMrk3casyAYNgOhAVVjBBulX+//Gjhzv+oSp7nmBiZBQqIYzOoSvvWDBsz0oA0CnT2Yii0HCTXT
okLwhE3ozmkXHV1eh7rdcyuNUUU8Fx9jVQC5PXg0Nw/bxdLdZX9PSvnV678Ss1o5UJS4Nz4E+tUG
5rIR7/HV4gJH+67cG5GZeLu2IjHjiXszNFGBc4dU2U7EtWdHv2MotmgNAk+fhN+Fnr/SNfvK1tPL
jHMC67K5AqwPxskdjfmLZoys5KbLifGUSes+B7wtu4szkdRFEnAlcq2hUJX/W4aG4bkPbMUVfARS
dHetecaji/agErycjd/AlHyI9fkuYi+GBJUj9y9u6/4kZ0rnNiA+2p3ddA1w1QXi6IX8IsZxi4h2
thcpSKfq2DGEZfqtstgxSdkUna5K/tMy38fF4IVt29KVBjvchegnknVrp3UIgLRvvUVEtzlElaV9
W770rTS4cdVqV8WwDgR5iq7fluw3wJxtsirp1lN0dTAxQ8sK7T6ktjkK2p5FA20MuVpU3h543Kd0
Ykn1HwH4WVhumaThJ77X4gxrI5BpcqZJDqriE/CApSg+DeXD6izSVi4xvZc46CXBtDfI5mWrnbgB
MzcrfPon3a2z68itUQ7UkXNBGeLys52ohIpE8Dpg3WFhU107sfgf1wwmgff0bn3q+QqU+5HaTLjt
nRVkMskbqpzKFbsgzjC++yGoKRaESnRS0N80LjJGYFGYq4gA3TRtWfvGk5BSf+sK13XtZmCVh98p
1c6lsDTRncDkr0iVZeEv6AkEOm0ZJc2sk7ICD+R9AkXDxIWmDXrOizERRc32o1ujvhgRuNOJKeOv
VL9twcuY1AhFnr8U08G8n1pHO3voiG2e8tLDs1W4L75TVeQyNX1dqcGo38WlT94jV1qeMrHxEUTl
4p0NK0gTejdunf8RbnJ6qWxqbd2LSLz7O9TO6joqwla7pZ7JMcNRcIrN6YFKFVnL/YtqyXujFkNU
9DaUJbstydyIVCqilDYu7Jytqr6q86hm3w/3oOcYbyZD5EZ+t0mFexYCqHWBw7TYQ8GPSAHRPQ2L
6HRI88ZjVc2W5WPuIuQKnMRgKop+iUbIpsFKxkth7NcpYaGFUZLl75YsxDTs13XDmH7MzM9K8Ep+
PDTeiFCfVbz2+wUnjNIlzk/J1cRE6NhVQRGbeJnisB1d7FmWBlagHmdAxcMlI17q1NT8rdIcrF7l
VOsy68Myigp7knwQKnqfg8hSi5APn95L/PEhkYJ/kq9RpandbP1nI8NRgul/rhJZ8g9XuRP4qJr+
Wt65qLRPtTVSQO5dhIhOqdyozMiMNSOoaiiEDKfsPeFYyDIFXRoYXwPU3hgbmyU5+64KZyM9whTX
EoR7h6OoIZhRtGs/UxkguuKQAu7tDGLBNo1T7jrdeqorXEj2yV3+DG28H8HkkozRowWTjKcT0MyT
gdZLa4QxuDNWh/EU8bM1VWROsH8o4LK4432FTN5IaGTmzC9kdtWe131vYFRI2KLppxK1rMXy2k6h
halAMrGDfxRJggV6SuQTW12Qw9EX2rHy4Tlyl1nQJwgSyKGV5+akkrz6qrP5DG2jNjyF3/XnXtVg
d2ZM/IuudU8Mj/rX2WKlZitC0jiZA7rmj+w7GvqX96K+6r9ZRbZwsBFSHQvrS/uhwp9u6a1tPRVN
wqrLphHo+iv0Gt7/GJapLVqCmQ5NO035ntQ7MJT5HfOrV1PV2sUTgnbCy3Daomg/vdE5LxA3QPU7
gy+sWdugK3VuBKjDIHqstCt4rb21iM+I+AWQ4neVplKhRSsHNo7yl0JxSgOa8xNdG9ZZqPJyRpkO
bFw3+bYAdzrBU0kRuO/Y5sFYL1NRFZQfpXAlfkicV6VmRzzgUyRHa2WHUz0WHY6SbharXU37yRCg
c62YslPzvODsYg6zhPaUX5vG7z3arTj6FDN79ON5XW6Gf1gXXjTvMGB3GAwgKNthelEBtazmmURJ
ETu6bPlSSgrnM3qlHa+BJT+dIDbH/YBcxzjPs9nM0NgDsQ4v8yOFB4bL/DSdQJC5m12yusxNOhen
7hi4V4SLiYq9jqSvL+uX/rU2EWfJ6kxyAg24cZx9NPKDn1BfryVr/xLOq+tBc/LalCwph6yZSLfD
Htn1JGdTc1xNdG9zEl5mV/+S6WS8umjkmS2aJLnEmu4DcUi/6/XMYdA2+hA5oA4wFZlgF0PrDkxc
OO2QXT4Oi16gn2bnPmn5uGWQFIGDSplMIWfM2g/1OqD0ppVJGCc+7T20doj/Nbh+4Fy0NV+sMp94
TppsHzC2q82dcy1UugYrQH011tWjnlEQqn2MBNqkwsFpl79cseh5kSPm4wt7773IhUkkoNUlSFaL
3RsRMgZynEWUQlnbNjlMSbqlPwskxGZ6mjHzlupHp//DL1nUm8voixybkxZABNqVMAl8mEcwotvQ
uJZZdgBXCnlvnFJAxHPd/L/5LpLMJub2d6pv7mLhd6cGAXsFVZmctCCB9iuj4vJ0EoipDWRiY3ec
xRzMXKocmuMa4SjGNWC7F9+EdMEULs/Nh7F/mx2zg4WVD3fQAu9fNJvcA7Cqew//YNO78dFao6tR
fFKN9M3srFnYjYfdEZmXkxv7Q94SXvihSFq5Y9XIJhk7zUgluUpuUIXl9jteUXunm+lSmrDyDxY8
am1+0GkUHOV218aEp09f1Obm0eV8gMv++3UQOZ7DiBoszFRA2/rrtE+9gSjlRzSwGeAXUy7Nzh+H
E/lEGLV5bQNn7Y/7XSq8N6Qe20mTCOiJDwy/tUod9y2H3K3eW9nDaJkhQnpAyL67kY3uk8AHvX3b
44mjf5NFN2iRaJa3qFz9v+Enn+48DHFH4KJ+tq9V5ofVzYQf+OuPgcsFaPBM/SHyJpJG7f4yS9/M
OamgCYsMjRCL0F5i5uxTewYDouIB5BUGMxVSZGgEmYty5/ROm4xBlphDY3AEvf20ShGV9wJXzk2Q
AFVt3nqjtKAxv4LuiS6qonpOtfr7ge9VPGJZTFwUmmTSKzmU98cSno9o11KKQupgGJzN1K61m06w
wzQcK7QYVbarjmut4AYdi3vRHgReIVl3x1BbTkKcjEcbJoB1lXkrbmWSRsC5BN86XZsEnsZ+YBBr
IsM76Vw6e5zzV9OHzjIC/SZtvY34s9rBRyjooKF20zKBdqLfBwPumEDwZhva+dOBhWQgTVuDafiy
0hfeuu8SUr8RCW/u+otaYf3s1+qR7a22/YQuJcxMUqzM2bc7ottu3cuk+GGwVePhGOVXZML/ubUT
Y4BabVoF4X6EOofjwRejoOJJFil4NH85cD1rZiGOzQ5NcxN8EtAfQxqIXaqe7W0oHdhyXQg0AJ0l
IDR5PiV3j7e9e8rXchMbEpLHfCyKJHJphXdZP94BYqvdH5gz4ko5mgmYxWM0N1HigoQU2IiSjLM2
w7bbQpSZRRFYB8vW7QSmyv3BtoChkwI9VIAhCh9OC3w7MY2sMZ0wCTJvmhhcYjuliV37tFSoGzCy
FpTBc8qK0LOM9yG+0X18YUHAgGfH67IiDl20lHkLVFe0a+LJzWsrTJhEASewhpplPVBVVloXj+4f
2RnrjgnVl0/Qq8z++eaa5YdYNyAnv6aArIWMyBe/L2YxnzIntGmTzGvMer9UgjUWhHvijCVL4Y7N
46dr1f/QTS3CwdPjK8NiWP0qQ14a89HbaSd05njOO8bH+aeZB/LsQLOrcyXVjeZXqu8an0ddBr6N
PnyyE3CpLGP0PxqWHXX5wKmXECUImnTtCYaSXnPntntpvkVp6ygMw7EEO2SlzhfR5hf9NVerzIVO
AxWdHsD+hvuAgkeWuSqCq2cOfU8oPq1WhKN1ei9EhgGbYH4Sy4Z157GQp1yld16ozVlXxi1AX0lA
On8Q4z5rhgIS/DE+64oDN+0Cg+2f2+ybHyVRZmh+3ENq12pWADiLFGg9yJJqz8fZJgODJ+ZbGuPh
9MUXR4Us7uwJBKvId+0j7qFDqf4JqistSwFR5YeoK9spZyQPDYkA7ZDqLLlLyt1u8PrsEjNsUa9g
LOnHy6oGvqdjBmBeKZjO6G9Ybc6CaYPHzEVzGnxfPZUv66mtRpDfr3We+WLBG8qp1IFqMXeR4mLp
WmsKDsKlz69a8hzymwBpieTm7wkey4Ruh8KpFDsRs2448kOP9Ql3A49BKZU423Tx40QwcFUKIYmL
CCeAjMQ4noqqOSFeCiuSlIpT+cEzSyiQVD52lAwPIbc2Vwi0jz5rU+c6HUy4E0sYPOe6dF1XOGA0
6ONlPuno2JQ4oM+sYSM5m/hIhnIYbjiRhnwJ0qtqeOUYDBz0as5MQngKe4VxNa4v4Vx2RG25odw9
Owdpl3QRJSzy9KcWP/KtRLos4QY1xHTshpD38QgoFzOf9LFs2MyXLQvnA55Nnp0rwGhxiJ7W5Ojm
IEzgMJqHdSvrR/Zw8yTATNeOhltWa5z3beVXdbiD3KGOG3MsCx6tVgPn0Vf+kOAxdfUbZnix/ZIq
E9U0Kdy+1TrmQ60XNy0Cg6xlYo7O/U5gwkKJvVjpoUMM24cQMEn2nY6zLhcPTIpqNYrpHy0T+HH6
r1iN6+NLRbFx7BsKwjaIrTMqCsr9XNGvI4OjTK5QiEiR1L4PAWjFFWNQn3EDACbblRwZ1bjGdTP/
Qc4Dwo45NdccPbrSj8MuAyineczXrztpAFZMFRJL9xNDlq9ZDfDriDhoxVqi7PQtEY/f2baYerhb
58vzX1oMYKt0gIB9SXvYmPRxfp/AYVD6eRoVARVGwLnNCEORaT6v5CIxztDTZGJr49bPo5fon2Ze
rajI4lg6Z/8bEIXG7w9HzLhHqLySvYySKaBzX7TqtXKFLGthmwpujZKL6R2Sh/KQzNVDREhJ6mZ0
V9ovRf1cB0wtvAhO/k21YIfrqF4D5VOb1Pu6rQep4wfJNVkYug+TrW7dADQdXtdfbmVYvx0pmqO0
l6xHkhseT5dLXjMYeORRb61SCt/kfBDS+VBec6ZBdPt7PUMnSUB94mEHI1jJF5jeObLgUpPW64NC
UVF0MVx+vb3utB24UszCnRzGDsoDJN2KN33n+Br7rFkm+QCTRoA7Oy2qIN5nV0I8P8puQYwq4pQQ
W4oJyPhRT8W9HIftmyeT7DUkq7AeiQgFLOm0JwnJizcRs3GwtRb+EYPdLKJ1rPHy2dF/JK+NZ0Ss
ea23Nx+JLX5wu1BazZ+EO6LQFSdnwyT3CWuGGtGJwwycgvbP9l1GFN/Td7tvMJ7XT6csS3LolzV7
9E8dpFMNaVGTpha6bsXhZOsXQAFCx9R6fmRqxZ1Vcb4TMX1qEDoMM1PQncbsvz3MF/mP67K5jPyR
A/i1FNrsVVOeYzYnAcd6gmIn4/0UwpJnhzhTefEaSMFgDluipHe4HR96QXHF51NBh5hmG97JaVW0
uJq2mm3KGKni7xpal/mGFg3xB7bIeAoP11jB1GofkstPXZL4ckpCQbR+lyZwU+gxeh0ME0HlvT4L
abK+uh7UP+i+gLRgCG6qH3zNhUlgYDVdBOW/HoWqejw4vvCP3E57x97G3+HDeEJ+0vjXQnCw4MA5
pXlSODDuWi9Yuypq/7Aj+Byop/D1UXRRcR0gELfUuLWLWn6xuQ0DuZGVl2m6cHBWWenwY347o9mg
pYpZuZD9LkDjS6Ck6+5DifbqzDQ0b/FVb/GIocIGYDub0VyYH6T2nexAw89Dw6j8EmL8iiogJKwg
q012e2bqK1uk/GF1O1wO4Xb/sCloePkeZyjvWzCED5MZfCYikJhOHZ+ITGBbqoWxqWzsG4jIMcX0
dzbPlmOT66s9sfyy8QpAOReO+nyC+ZnD9ACZSkOFo5PpEWt+lWaPOm/cJ3HakQHZdBrr9eFo+1yC
pXegbBFh6SOdaSQjCvPBZOYUOpLKTRKdKxi33YC3VGhnVW6l0PNFd0Zm4x2TVj7RMJrGnW4Wg5ER
AqoxwlLkVhEdl3TWmgX19L1xpNKK2DVnApZN7jFZtzlTIajH/bA+xchmBuMzYwIotc8TrsF0sTVe
VH39NkErUCWlB257PsC4ZVWMUSd36S+Dse9WlYuhQk068d8XgqccDSrG3RXqXVgMNf6s2QG0f16f
2DXw/Ce7B20MWIwlar44+um4rDsBn57vD02Ln3JZhPYg2yiNzx6aSYvhaZ5XBQMuwA0iUPDlOjyz
4IGiJ/Xxcbbt+OcFV7xWFLHw5JTGZ2hCROtO19rn5atKUWBceSx9AJjEGuFgyV3mo9VQJDcTDXSB
L8BvLP3GTSx49Xe3PZR54RcOHymevr7SQ3AOjiNU0pusWjLbt0VO5YY1WynuGuaXN45GbY+GN3gV
/pVLHMMFKCl57qw7zdc7+XcWOK1kbwdOlQqwee26i0zw0oIS1ROAJNx8tPq8DoKh78T8X8w6swt2
oGVsOxK7ivHrsPRzvuau65GVq4rJDV/cSryLBN5m/O9sZkz8OzEb7a54lBptIv4JAHSfbHuUYWce
CMx3fjUcO+veBhVNV3P64f77yC7enbKQ/yckB5KI/byZ4+OBXf8Yjd2popTzZVu4KxsVEcJgssUq
3ov4/bUMiHYJEPdc8gtIU7alnnKQhx2qGaalHJGzXEkoQ1NvEW9bE+Zm9PngirWTmTW7HPpfmaSS
VCI4tX3THizpIm8HSIWcw0dgmrQkLEH6uBQv6TMwcIuYm3HstcXMVRI4XZGYTWHO9xeaAdoEaic2
+/Q+DC4E8E4trpHcWtvMx5CPdXvC/ZJRjonshF+FXns/Dk03zX6ZzMZHtcmskaj0coZDRTpsclNT
noLnclfiq7CTmCTPmHW8hUWHG6RP8a6L/p4rXxRGZi1kRXnEF0w9w7CjlcTuXH1OZVpCTePmnsUb
aV2wDVOm/XaDdI+UqUGZHfrYpcqKT7uEw7uapkB1jW+ATJ5J7Gt+ogL4l5LvoKPeVp1NB2reLzFK
YkGMtWpeeKYjoprfv0dOcKGHTYPXqMdO7PQ/fIQUBk5VgMI2GTF+t1H6A5mzJ47VGk/0cu0ImlCo
r7CXaF7HJ6gxVF6rpMQaW0wRsv3+JNk0aNemwYW2wEA1esnramrXUnoghIcCUlNLVlDEjhRjSAbe
8TInLhsh0ppCuccmD5N+poSfSgyWgq7rVvG9Kw7CjtUFh4/LauRCbFig+eBJlDu9RcUz442DdQWO
7nsvCNOtbqR9u9/3AcGDbNwFd0vbgimxN9CKCh9qx3TP5EE1E4mCaIk2OD8N6HWyMz2fn3mMCxZj
O8ecDoGEQBWgElLL0HVLHSqOmDjbMTOAJ1h+6RX0PQ1MKEoB+4PQaFlDnIR2DAVKbcPok6b8v5By
3RV1+IMBbvCWGHu6FIwKF4g4ED4OUP8FOn4v/fmuzk1UgOC3V4pPzUJQL8aL1y8fcxadkOB5fn6F
j9btVRux/6SNVIb2olXaNExalGo3FyzT5688343F/h79biIZpW+Kczgbkz8saRAm6Z1ZYevxI/3r
h74zCwyydHVcUYdagkoT2BfmVw9KMhxVLE246RlH8cnqXnIURHNM6/mfqtUmpkPQR4kSDZsEh6Wn
IkKZHhl6Fg69tsukO923KEOL+C6g5ftJA0FiLaamKfopGBWKetiFKaeTnkJUbdEZIItkLe7vEY7D
RfP4/t6A16vqOfNnLV+dOT4rMpT04//GsOLZAhAL6or1ThYE5w+YngKRKiAsLwVxLj4u0+8iyP6g
JbNK/pY3uF+7ETxlmCqE0BHLplp1iuvtiHul5cczEIoKcOqQtrWqb6+sQm3fmldFqlHedWnj2P5e
P8AHd2Ecuih5tl0zscnqO32YRGZYY2Cp+5qpsFE0yK27rqgSZy9Z4cNk0bPXYiVKk1KjyoCo0nvZ
zBNgNIxK3WJiwq4ekhcG2glXZnWnrmdC/piuXGb9qwgcuGCNpjWTn3VoaPgtyFOKouaek3qtUcMA
HjSgMGwgo36wJwbgo6lxuTqcOK/aCXtaL0oUUaIaqe3ibCBiQR/zI9W4XT+TiKPuQYd8XNHBbQKv
avigMH1q4eAHL6iLF8BOkmCRBDIekcpUQ9YUpWQuvDgldYBOfuAyqs/EtCgqj8k9OSxip06jw6eF
WUO15IzlgY2kyPw9pPWdpNdt1hW/1UUKF5iPDw7EgxVSTtixNXTGb3oSbBS0j43XmK+uMEgDH23g
7bC0EcCJuAkLTpPdSV/zq5TEl5JkwRRqrwIf0mq/bbqQLahItBUUGN3T145qYN/px5+IhRY+oP5r
M8VzVgX161xRfzLi7PhhRYGCo5aIWZiOYE74IzZslTcEbDjkRIxrpwiasAvY83Xi7U3wf/uBnJA+
U1NmbwLCBnjmGDnvTlEbWgstXptuAU+LsPGpM8JYTxE4gJoAM4I5c7lnH65J8bmjazb0mCAQY02d
uQFv+WpJSRVEFFESWjciKqZFW/7Zpx2rYsGn/mfja4Yf23OYR5g1bDFjHDA//CQKETGafRumnYYd
//ugzwZiM7D0po/ITgN/j6oPM4AuWQC7VHY8PfD7/cxdeCSJ4y18MuOGjr4Twfu3Tm2VUg/hcJk8
uZaRt0JHDNCDOZyD18XoNt9nmGW9KV6LgoP34uYos+moBSI1De809Kzj/YGiepTpbnFecQbms90w
If2V+tOJYcLfyWpAvSpYJq6OPp84Z2gp0rf+hTT0xXpKFJJypyrIlHmkKHyCWRVn33PNNenr9Jlr
b0gEdervrtuvmbLUTzRk5/gFCoTu28rlfVxJfeYaMgMsNubaczHFTvbFZERi/XoEONGCDxcOI2Hn
ukBpXi35gX4UyXy+LT+eCYkobMEOG3Ra8oY/SbWu1j1Q713wd+GCvVKeflbwNaSXVn0olBUnYwcZ
+KPsvjC/5gZKMNC2z6AVIrQijmCTPjS5PnFv7YwLr13ajC0yVC/RksE4/EJSMOiXHKmo//af1a5x
Ars7Ej+IW6UjDwYzfMmcIvk6vYRWoZtKImUgjxxHfjTPJ2RKPp5aayKom5LLGPbBGTMJsHpmUePl
9Coj8Cy0q71AbHYOnRPQnL5zA+c56czigkoBoTXzSxlpH/85epmgH7RgwnNHZzHw1uFZZqzImXCv
gWEtzV9yzC4xQTmru7iVKt/4XVGNHS95pcoxBI5f2AexasD3OIj/qRohFi4uIT44fFEpHLfouH1b
ivdJ4VehHxQlMkj5lUH7S4rLln9N8ScXPejmPA7DrnZ0NwoSODv/TRjuZSvXQm01G2OzFexA3r0V
/UxHBp8mdfD1vefhNKU8yX4Ev4XgOra92zTv80M2kNRBFTBVZ+CCqXk+6BqtIfoUl/FLcJfV1QG9
0iyjbGocNToqDEhhe991UT4efC8RKaGHA4QAXBEG76pRMolnwiuOW4ymlaIv04WWu+zsDbM1opkC
PIcLhYgHzkbVKpnPfKBx6T84jKbH9459rFn+43rz/eudMK1DOTKwAaf9+IhowQ+shVkuoxAAgzJX
OmfJaSPfisNZTeq34xEzlwNhC6nHQxxHdnbqS5c6Au1gsa+iM3bea+9TPG+y2MXIWmFhI2raw46T
PcY6pgAPSk7gkCIMDgwMo4PlJLkGqRWLmeOR1q6Mea0tUeyfq1Jg3ihPBQ/dcnmTVODifEpQoua/
87EumVE2uLmqKE+F1UQJXPcx1/gaBl6n8fJwrTJTuyLlB2n6VNQDqVp62vdI1FQyJw+CCXjkykNW
v6D49cUn4D2h5IIjc3vjmmvPTubLsIrdcDDoVExwTao7i39gdoGTbWB7D0XjZBAUUCRPgC5p/5aH
ZHdiUiCGTjMZ000Jbt+5AArFFERBuTrAs2LJadtKB8weujSBXTR93iFUnHcSq1+m6CduXmxg4PDT
mELdJBBHyALkPWU5o1uvouYwrZph+prPnNVjxpr2kjJwzNt4MjzjquXXHSIZhz6Grut0P9KW1GgI
Cp5DbvqTeA5fszh1Z5SUMzdxDiF82SUe6QFRtI8UM/UyWOITBEfsxkZo/dyeFYtzGSB7XgvGXohE
JkLYQFsTqbOtu23jZBhUxxAB1+71Hg0KS72Bs2zKpepep37J6Cm9PpOytSfhsZX8pi2gtATzUyuC
QbkCLyE63bFhyC4GAHEV4TW7JI+3zZJlpLvPDfESfF1t3r+7ONXO9zy+1vcO/8JAHhe/+P2p0d6x
HPDhRIR5/5U1K9ZHEbrL7io2jYxa8ORvf5bkI/xl3pcXaehibYbZDag/6sZHxu+B/3F5vTS6rWir
DJA08337+iHA+W4W+sdzskOOdM19BV3WKYpQJZHobCas7JUYBCXkxOs2JDfbiIXreeVx3LmTxCeJ
V7HlOINYvJt9SIFi9qHW7yi7ZXlnStncHrLrpqDvwSKeomPHgS1hUNBTUQlOa/fMZRR/Qyw50fbk
7AgiYTkqKyZZMlFCqm8Xduzfqhp0gud7QmtzWbNtEUwQszTytby42vEOt0BfX8TDWZEjr8ddJASQ
44Mv3Np6p00xodErQQYYRen6P5+f7qL/v466fZ6sxHYht/OfZTjmyG5G+HN8JudbeeiDU0RR1yUN
bKmr/j8Yx7Y8cUskd6kDynVt8+AhQKomZ9RvQXkMTrW8T00xu9q1FPeu7owkAPuBtmcnU/76YIF3
AnF/s05wF2j5SKSFRS9C7keWIWcTYsEvmHJnTgdxDjg0tYfGjyGO9fyZHwlpdNCMnUTo/3YNGNDj
cb4rBRglUy0tgOM3Z0INF+fBeAJpqVMOznGHUkJkBw8oJEBXWo3HnIAkFaWhYU6dWnRj7wnJaJd1
5Kcj/li2f+GdLB36liKVpUlsvEXafaRD88c/iSRcY7gjIr68Y7aD0RiYFuIXisLwSCVkR2tiMmFn
ulHiu93J8tqa2VYju5XkOmolkJGyK3wd30hduxXf4K0oi77gblefdVBsnbvT43+49cQuU+Tc8x4g
1wGF/jF3y5rp1TZ0cttmPP7SmSXYD/bBkuc5I/i0PHfgQER62GNEg1gDimxJBkl4XONcnYs+xNaL
UnuHUlZfY/A9tkioomt/njqeejRxcdYXYZo7hpEUqLNDuXInEeef7pNuulO7PISDl8JO69FIM23m
tnqBXgxWPe/yDTzmJ658YRrFM8ZT+55WQ9Z5htjntuGoRMO6hjKKXvw1+uUvPFctYGg4zIfZ6pzl
07wdMU8dmPuH0xloF+ODN2LaOU2AKLOwOvyo5kZ3662Uzy6C2mhJstLR8I9GK1jf8lyYc8GqTflq
fQOsJI9m1wEsU1Li3RI0vpa5xhguv4ckdu2+9JX7PLXtOThMiLjJDTP4FvG5dQ2PTwfqhiR2mfaD
NjMKP1W8CoywrplwpVhyNpJf2PdxHe6RFZRR1TxIOrs+ztjGNc1Kk8v4KsxhrcIyHVbZZAqwnvYT
6oxmvgnerItZSA5oktnrP3d4eokAV8GWitB2Y0YION/RH7VDmTUlZ1CaoTvqCRud/TcH1YJrv7mD
Z55VVHctkXZOQXc2gc2CHIybXUf3QvEbIz05eJrP125YTrCO5Ir2+KUDWga/K2jvupIElm13g7sL
m4KBbSsTZ3sqjULS4cly+zzCLYwjPTmkgUK1MT8wGpXzX2mvqW1PXBHdbseDchrzRfjJEemruos0
PNO5Mfb97G/Of3PtXo/oHG6Csj2WGa2aKNY7HZVAtjyohLRHMLSVJzEf+eG4yWL+iGUHlAYHnqcB
IVH7RkwCekQ+7HSSaArFeOnojxOZUZcFSX6M5TONkG8uk29UpAEBM+/oLJlX+tv3p9/raZ5txWp0
lLp+yzrKsWZKayljTHhvZfDTXgqI8ApX617h7tKXZQs4aBELkFLtdrRu+oDMShmKdtpzVllMlf6O
L/B6+SpPiWp8j+cwwRoXoXK8LgfLveCYuNBn0RQKv0QomIU7bC8Nzr2BzIlJ7oLMBhq8IX4+4NBx
osvfIXDFW2ETVX0QCxLtbUl5z4o560HNJKxooTX0gqk6a1Pe5fBQltZdLGYrmizRXd5AR4LLz5AK
RupGiy7TM3vsGZne8j9PkYX65liVZazy7q58Gqp4Nl5hGlMYkYNqJM68jiNRPL75TN1gCCDx2jdd
4NU22jArsDg/2NKPyQSyFefiWhzJClbGF45o7Dx1VGwQVWmZqt1EQNLSmMTPDB/IwDbz/coY+gbA
QpcnsaL7KbQGIBXPnvTmodRRVVqffUjigoOqEXVf6dbzup12ui8nacT3ZEi+swZVqIe9VJhV960/
wlr/WEWZGCeA99zSHhhNjC0CKDIgXSpB6q4oUIj6bN3BPHSHj3/iaUzztthB7jgmM15+s+hy26uj
K7Q0kA0a/GH8DVtVw/Kwlc1x8xHQ1VBj9UnTZAwRJJ6tFTOiTnZSXmsSedJUg9MyxeLWE6FYG8iF
H6rKJIgg0nfVPK7wJIKaHF5IbbnftsVplsQgRY20OGOAs6/VuJlfjmBhaZghh7+MUI5hNtR6UZ35
Kh/1V0IdfntrpX9kSu3YAXqjcq0JlBGAS9EHpGLxlegUi/hHYaB2+Ro9+sIL2xbMJBwc5QislF8d
8PQylzBo7fxiqJCWfQBkqUx6cXPq3dA/Ld7OpcmumX1Eqi0FgPyVlsXBHEfiiZ7ps8qYSXA38PJJ
m4mbVkmclIDqvPpEO6aoSU5BBb1hgWp7HR/4wgtdh19XPyMDvZx18lzhA5fuYPJKLQ52TJT1z88N
pWNVNv6ncCFIx4Z70M8IPlnwhDlQHT/IlES2Ts3JsYaJO9BpZz6sXJglgEjJ17f4ChwLeBjld5Vx
EroZ3LNCcpxcmvbwBOg1wbqoRlo8V5jflmbhO4IMn2gK1704oYZvrte6yrX2GMkZMvGasVUQipZV
tC0kzlXb4jHjHX2dUaXcow6mSjnwxJlepHwaE+Iq1HZRHJLc3QS3z67SDXO3t5UKF2BRVmQIBApG
YCYiCBgInyc0LIa6puBlf4iNYhWlODYwexAnIv9xnCjqcFpy35kvbANOAWmKn7zn4pd7BrqheL+k
F4cKUiG6njEjIE7c2dpTX8bCOExEwBxErWTtezxLtYbwMW5wGzIMzftImbuFwSe9wVZhq6KX9I8b
EqdoET8U4ZKhr3WpyQkbaICzqMyvd9Y0S2M1o/8FMHF4mQP93jsCfmJd49TYG9rh6OZb7WeXowbz
iR6Lbp/L58ebDE4mljRZTlPvT3W5BXlL3xe6X+GQ0nFRDwx9IOoB+fvwF0GNtC8Rrq4MDYozKfe+
Yya+NqCqPxqIftCvls7BGzDmcvDDex4mZiMZ9RizblE96ZH4MjwWuclBbKNTFRTASdZoLOYe+fVf
DuRj8rj3Y8eWsIsx/snWpH5jdJ7pmo8Kz/NYeLnh6AwkzoS1+DHU/zCWbRK3YGPH3dqxvqHAVk+V
5nxYWj0tivL0KZwXbpohCBX5pSruCu3O17ESRUF12zF2EQHXaYxMuOjPBanSsuKzYDsryxhN33ws
wf55Erl+q2JsFbQ1ovDS5vGenxb0Q+i4MZKgHISTFeh4WuRqqdVAmWHL5IWfZPPp98dSQSQhj7kN
kuLb9K9YkJoE1MsC8HFDs/iuk97ZSH9Sp5poddPGXuXjGmU7+E4dniVD7krnvsONJkZmweWCL5SC
kRlX4pqpm2/mPqh4+BEgiX9zvDP3AnBlpFGHTvpPLk1XUv0vmGky+pW9C3KRzIeW9wfsHUfwhHQq
o1h9ziBu5mUorFuUlnokCGNwRB0H6OGfOcuHkEZOwqtAEC86SiVQNxHtD7WvqtPiXPhUYV/luluK
LR+ifF2GDt8UVKtg0iEih8D5nqoFVniGbJoF/UNdmMgzTMP7nvUYLQrqkgBodbGjtIiLOdu+5WXM
TWWWY4QAtuRGUWkml2BwJ6Q86NaQ9j7A2DhnO3bY325tckmYGjGJIlgFWmHmrKeQNQbn1zAtupA/
zYFlYQH3Vu1cCrMnXMzNOsfMgLdD8FdRRIhjrzk//bsmN/6rdtVNFktRe9wLeSfjW3vK+khVukXl
uu2IZS9Aj5spiZlw/GwUAq8ukC2uerrJFtpTHKOT6Jivyeyhz3SQ8jiaPHXedmpKcM0VE6t0/HLe
E+Lo/CIKOpLA2iW+ep7TsMOEIbfn2SR6b4wB4s9sDB0SHJKI/YGzggOTsnlw2kKQ1NkvRxzQXNRr
AyH9zjjdCzj7ZAOgs56/nqW6o5HQSlvC1lJWYbLW97nGWt73+DcaiTjn3ZdIihW1enDy7kjSt7EV
8RMhYl+SBJCT7p9AcLsZrnKlpSUb4V++mG3bon99Sk5djTirtwmK470snigRTj79+NrvbmLGiKXJ
hheB7HGBLvqRp1t0wpNf8VTWvUmEzGtoXgk9GHZJNbAXBGMQs9S/ETQTa0t+I98JueoJ6uEVYqRT
cvKCTlZW+vUVDjrVGDPEd1DUyDSQuUF4rdtsxxjMxX3Gb4WHV2DmFWI0iMqF1N5A7/E4Ox/sPxgs
9WF5lj6XUsSGoFhEdxEGp77SrkYBo5O5hoxVq2LLqqhSIsnx3OIQFYwsjdQDul+jFwbZniCAp/tw
wll17T2mzAWLV2471TJeRp690YxHHfhfEPhZ1e0oLNba7MIKuQAdKcul59VgRLIHYBaRKVNfHKRj
MLfZi5xauX9ROioKgDyogfUknO5DEfRwrkBRo/2A3he/+ONMICRZui8ZrsS7PFm/ZCGVVk3fP3Cj
YewCNxo9JIy13mbmVN4Y2NE8teWRzk7Hr9EOLCCwuUBKWmaFap7dm1uJjVSPkySaTRL7UfbEkdWH
gc/wBHL8SCSs89rC6NRm8FSUi1LjqF54zQXybuZHui9fBrqr7uCk18Fpc23ZGy+utQL3zxKJx4vo
cqClaQQbL2Tlw2Pk8HUbXSmsck/oE7QaB6J/QHbefbKLtTzqpYzvJzrM863MtM03Ho2xK2SJaBw9
YM5hJUGjXgA7u/gcIYQx9/5XAjleQW2ci0BCgEhWX0DgOenoeFGkftl99wEmAyCyKuNrGimVq6G/
dhu+dnUox58LafV1SCeO3SO/PPK3HYFlZ+Ymcl1l+Wpuu/3/x1oDAfSzn4M6mVa5Q7OAlZtRGIZi
ZVSYdRdwsRFPDqHH4J3A7WWN448zk8IJn2piJTxcYkpPNoRqQMuWx1r+UvKIN6oL3w6AkbuaKgGK
4nbsPGITPlisDUftSzKCMRr8bgecgZWNWF8l41YjVYuvi+QkUiUOUNlAcxkGhwvX1ZqU/Iqpj4vh
l6SJmP/hq7ylSt5Vb2ylGkoJqFcOJ+x1kslDFBEYCCwvBkCBZX11t9tpAPQqMWPnGOWmsjQAfuq4
vwOcVo+64dGJTw8bGpkA1WPRJbX9kJvaeHNC33aVsJ3Jyxq/EHOvZzfw4mLEb1xW87rqF5sbitc1
IU7MML2fTAn+4esAtaqJ94RQ2s+zVbmy4cnQbMTyOAhxAQqcF9u08uPGK2jFhIFcIoyDJtfC3t3p
IKpuZrKRDCyRmHiQoApEO2q8VtuLo2v6VpV4LIEVYirvNzVMje8oFbSRwwCfNRK8sh4Tg0AZbZo7
85GkJYx4+njmB538ZhCS5cXlx1hzHuUGTsSvxE9i/GbFDCY35CY6hRUpr4pLNMTJWkWLFW12ChJH
lvIRkkG1ObJ0OpkKJ78k1Zk9nXsN7G2Ra/4wmoCt/hGjxsVqHI93Mx9MBrbCBWqCcElPtESEGCyW
CgdrHlR6AM69MiBapayVk7lpN9+X6SDRw4BJOV66ahPGVCrn1A+qqU5mYw84ysSscjAWtBN5LmzS
tx0O1+J9mMnZifEQ5TkBH2HHeImS/IXs32zApi0SuAb0llywTRVrZhOoeSWt4pG16N5qdRqXnLvk
lxQtCprgpMQ7jxdP4+y/gcQspXK6ua0oz8Ecd8F2s+hcMEDF48nmsOgPeJU7RGBhQLiRWJhGuhR7
Xh4NdNM+hv3QKHHf38IRJuJeorUbLJkRjFaWNGqCR7We6pCHEV07gMJ4TaO3a97HFslpfmMWt7SU
xYgnP34Vwd06uVknNeIM4LgDF6CKfhZ+Fyb694o1YzezqDIAWJBoZpkpjLxHMqFxkfkxmghEJKuV
fscSTd0vzYZoqtmf7u1NjQ2+5hyxyKpVbUBUi8YOOzYX8pJ2BTKB3Xd4liFtKnM7/amdQAdn/JeI
7esdG/ncXsEfdnQ6x1/5ztTxrMhC0672STLY9Y0xFmHAM1w/Ku7IIVGMYKf4bprGsf9BhdArD9Mr
fc0dLOp5RUHFnSRz7R8R2KBZ26JY0DZ8mPa9OdBI2387qK9tBEIjD8rFs5+4bk3F1Owlczlisfw+
1D8JQ1PqEpD3UZqXjcDFCv7UVjriIWCAq5Ranf3n8PcUtgWGRxigy8mWMnUlRXd8iSYrlek4DwCo
AR3c9hqo6N2nYaJRdqP9GdWYGbnOSKGkiLtedmD+zPRbJtt++1V6VlgfZ3CoypccJJtHiGHfcNvg
He5wIwvvywpQ9mRJRalvaU4vngkK4AHM58VdnLoIoGha1eeOF/FsG0FhOt+j9OZZv9dI507D5oQH
yMXyTBglh7K3eV7fBvb/2LuCMzctqtsZxKEi5xzu+WhJ8t0yWZXSIuP1VFVjGQh2FIRJ6jfpPxUx
nGPD2qXR12tHTvVGWBo99bNlcyQtQCucW+OFdJ2krwH/gu4gsaSce+xu7euThp+l3WCWGLCTr30k
RcgnZGIgQ/DpgxkrpZRN/rfTEM1ikxldgWzn5aumgLJWG0dUi6DWQj62966jAKRWGmzSSKE9Ii+i
1ghOu1UUguHn4wYQK3yJ3qHn609FJKEXHP/yhU2FmkyFWPF2DRw+kDZISF+ex3vTyHNQ+JFRFbnn
8muxVl00g9D67G5lb16p9EEjynhu9j1Bhvs6yZFBKNiUwttnVbE=
`pragma protect end_protected
