// megafunction wizard: %ALTGX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: alt_c3gxb 

// ============================================================
// File Name: rc_c4gxb_tx.v
// Megafunction Name(s):
// 			alt_c3gxb
//
// Simulation Library Files(s):
// 			altera_mf;cycloneiv_hssi
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 10.0 Internal Build 152 03/09/2010 PN Full Version
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module rc_c4gxb_tx (
	cal_blk_clk,
	reconfig_clk,
	reconfig_togxb,
	reconfig_fromgxb, 
	gxb_powerdown,
	pll_inclk,
	tx_datain,
	tx_digitalreset,
	pll_locked,
	tx_clkout,
	tx_dataout);

	input	  cal_blk_clk;
	input	[0:0]  gxb_powerdown;
	input	  pll_inclk;
        input	  reconfig_clk;
	input	[3:0]  reconfig_togxb;
        output	[4:0]  reconfig_fromgxb;
	input	[19:0]  tx_datain;
	input	[0:0]  tx_digitalreset;
	output	[0:0]  pll_locked;
	output	[0:0]  tx_clkout;
	output	[0:0]  tx_dataout;

        parameter starting_channel_number = 4;
	parameter pll_inclk_period = 6734;
	parameter tx_data_rate = 2970;
        parameter effective_data_rate = "2970 Mbps";
	parameter input_clock_frequency = "148.50MHz";
   
	wire [0:0] sub_wire0;
	wire [0:0] sub_wire1;
	wire [0:0] sub_wire2;
        wire [4:0] sub_wire3;
	wire [0:0] pll_locked = sub_wire0[0:0];
	wire [0:0] tx_clkout = sub_wire1[0:0];
	wire [0:0] tx_dataout = sub_wire2[0:0];
        wire [4:0] reconfig_fromgxb = sub_wire3[4:0];
   
	alt_c3gxb	alt_c3gxb_component (
				.pll_inclk (pll_inclk),
	                 	.reconfig_togxb (reconfig_togxb),
				.reconfig_clk (reconfig_clk),
				.reconfig_fromgxb (sub_wire3),	     
				.tx_datain (tx_datain),
				.tx_digitalreset (tx_digitalreset),
				.cal_blk_clk (cal_blk_clk),
				.gxb_powerdown (gxb_powerdown),
				.pll_locked (sub_wire0),
				.tx_clkout (sub_wire1),
				.tx_dataout (sub_wire2)
				// synopsys translate_off
				,
				.cal_blk_powerdown (),
				.coreclkout (),
				.fixedclk (),
				.fixedclk_fast (),
				.hip_tx_clkout (),
				.pipe8b10binvpolarity (),
				.pipedatavalid (),
				.pipeelecidle (),
				.pipephydonestatus (),
				.pipestatus (),
				.pll_areset (),
				.pll_configupdate (),
				.pll_powerdown (),
				.pll_reconfig_done (),
				.pll_scanclk (),
				.pll_scanclkena (),
				.pll_scandata (),
				.pll_scandataout (),
				.powerdn (),
				.rx_a1a2size (),
				.rx_a1a2sizeout (),
				.rx_a1detect (),
				.rx_a2detect (),
				.rx_analogreset (),
				.rx_bistdone (),
				.rx_bisterr (),
				.rx_bitslip (),
				.rx_bitslipboundaryselectout (),
				.rx_byteorderalignstatus (),
				.rx_channelaligned (),
				.rx_clkout (),
				.rx_coreclk (),
				.rx_ctrldetect (),
				.rx_datain (),
				.rx_dataout (),
				.rx_digitalreset (),
				.rx_disperr (),
				.rx_elecidleinfersel (),
				.rx_enabyteord (),
				.rx_enapatternalign (),
				.rx_errdetect (),
				.rx_freqlocked (),
				.rx_invpolarity (),
				.rx_k1detect (),
				.rx_k2detect (),
				.rx_locktodata (),
				.rx_locktorefclk (),
				.rx_patterndetect (),
				.rx_phase_comp_fifo_error (),
				.rx_phfifooverflow (),
				.rx_phfifordenable (),
				.rx_phfiforeset (),
				.rx_phfifounderflow (),
				.rx_phfifowrdisable (),
				.rx_pipebufferstat (),
				.rx_powerdown (),
				.rx_prbscidenable (),
				.rx_recovclkout (),
				.rx_revbitorderwa (),
				.rx_revseriallpbkout (),
				.rx_rlv (),
				.rx_rmfifodatadeleted (),
				.rx_rmfifodatainserted (),
				.rx_rmfifoempty (),
				.rx_rmfifofull (),
				.rx_rmfifordena (),
				.rx_rmfiforeset (),
				.rx_rmfifowrena (),
				.rx_runningdisp (),
				.rx_seriallpbkin (),
				.rx_signaldetect (),
				.rx_syncstatus (),
				.tx_bitslipboundaryselect (),
				.tx_coreclk (),
				.tx_ctrlenable (),
				.tx_datainfull (),
				.tx_detectrxloop (),
				.tx_dispval (),
				.tx_forcedisp (),
				.tx_forcedispcompliance (),
				.tx_forceelecidle (),
				.tx_invpolarity (),
				.tx_phase_comp_fifo_error (),
				.tx_phfifooverflow (),
				.tx_phfiforeset (),
				.tx_phfifounderflow (),
				.tx_revparallellpbken (),
				.tx_revseriallpbkin (),
				.tx_seriallpbkout ()
				// synopsys translate_on
				);
	defparam
 		alt_c3gxb_component.starting_channel_number = starting_channel_number,
		alt_c3gxb_component.effective_data_rate = effective_data_rate,
		alt_c3gxb_component.input_clock_frequency = input_clock_frequency,
		alt_c3gxb_component.reconfig_dprio_mode = 18,
		alt_c3gxb_component.rx_cru_inclock0_period = pll_inclk_period,
		alt_c3gxb_component.pll_inclk_period = pll_inclk_period,
		alt_c3gxb_component.tx_data_rate = tx_data_rate,
		alt_c3gxb_component.tx_pll_inclk0_period = pll_inclk_period,
		alt_c3gxb_component.sim_en_pll_fs_res = "true",
		//alt_c3gxb_component.lpm_hint = "CBX_BLACKBOX_LIST=alt_c3gxb",
		alt_c3gxb_component.lpm_hint = "CBX_HDL_LANGUAGE=Verilog",
		alt_c3gxb_component.enable_lc_tx_pll = "false",
		alt_c3gxb_component.enable_pll_inclk_alt_drive_rx_cru = "true",
		alt_c3gxb_component.enable_pll_inclk_drive_rx_cru = "true",
		alt_c3gxb_component.gx_channel_type = "",
		alt_c3gxb_component.intended_device_family = "Cyclone IV GX",
		alt_c3gxb_component.intended_device_speed_grade = "6",
		alt_c3gxb_component.intended_device_variant = "ANY",
		alt_c3gxb_component.loopback_mode = "none",
		alt_c3gxb_component.lpm_type = "alt_c3gxb",
		alt_c3gxb_component.number_of_channels = 1,
		alt_c3gxb_component.operation_mode = "tx",
		alt_c3gxb_component.pll_bandwidth_type = "Auto",
		alt_c3gxb_component.pll_control_width = 1,
		alt_c3gxb_component.pll_pfd_fb_mode = "internal",
		alt_c3gxb_component.preemphasis_ctrl_1stposttap_setting = 0,
		alt_c3gxb_component.protocol = "basic",
		alt_c3gxb_component.transmitter_termination = "oct_100_ohms",
		alt_c3gxb_component.tx_8b_10b_mode = "none",
		alt_c3gxb_component.tx_allow_polarity_inversion = "false",
		alt_c3gxb_component.tx_channel_width = 20,
		alt_c3gxb_component.tx_clkout_width = 1,
		alt_c3gxb_component.tx_common_mode = "0.65v",
		alt_c3gxb_component.tx_datapath_low_latency_mode = "false",
		alt_c3gxb_component.tx_data_rate_remainder = 0,
		alt_c3gxb_component.tx_digitalreset_port_width = 1,
		alt_c3gxb_component.tx_enable_bit_reversal = "false",
		alt_c3gxb_component.tx_enable_self_test_mode = "false",
		alt_c3gxb_component.tx_flip_tx_in = "false",
		alt_c3gxb_component.tx_force_disparity_mode = "false",
		alt_c3gxb_component.tx_pll_bandwidth_type = "Auto",
		alt_c3gxb_component.tx_pll_type = "CMU",
		alt_c3gxb_component.tx_slew_rate = "off",
		alt_c3gxb_component.tx_transmit_protocol = "basic",
		alt_c3gxb_component.tx_use_coreclk = "false",
		alt_c3gxb_component.tx_use_double_data_mode = "true",
		alt_c3gxb_component.tx_use_serializer_double_data_mode = "false",
		alt_c3gxb_component.use_calibration_block = "true",
		alt_c3gxb_component.vod_ctrl_setting = 3,
		alt_c3gxb_component.gxb_powerdown_width = 1,
		alt_c3gxb_component.iqtxrxclk_allowed = "",
		alt_c3gxb_component.number_of_quads = 1,
		alt_c3gxb_component.pll_divide_by = "1",
		alt_c3gxb_component.pll_multiply_by = "10",
		alt_c3gxb_component.tx_bitslip_enable = "FALSE",
		alt_c3gxb_component.tx_dwidth_factor = 2,
		alt_c3gxb_component.tx_use_external_termination = "false";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: PRIVATE: NUM_KEYS NUMERIC "73"
// Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
// Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "2970"
// Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "0"
// Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "2970"
// Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "37.125 38.076923 39.078947 40.135135 41.25 42.428571 43.67647 45.0 46.40625 47.903225 49.5 51.206896 53.035714 55.0 57.115384 59.4 61.875 64.565217 67.5 70.714285"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2000"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "N/A"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "37.125"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "148.5"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "37.125 38.076923 39.078947 40.135135 41.25 42.428571 43.67647 45.0 46.40625 47.903225 49.5 51.206896 53.035714 55.0 57.115384 59.4 61.875 64.565217 67.5 70.714285"
// Retrieval info: PRIVATE: WIZ_INPUT_A STRING "2970"
// Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_INPUT_B STRING "148.5"
// Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "None"
// Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
// Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE STRING "2970 Mbps"
// Retrieval info: CONSTANT: ENABLE_LC_TX_PLL STRING "false"
// Retrieval info: CONSTANT: ENABLE_PLL_INCLK_ALT_DRIVE_RX_CRU STRING "true"
// Retrieval info: CONSTANT: ENABLE_PLL_INCLK_DRIVE_RX_CRU STRING "true"
// Retrieval info: CONSTANT: GX_CHANNEL_TYPE STRING ""
// Retrieval info: CONSTANT: INPUT_CLOCK_FREQUENCY STRING "148.5 MHz"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: CONSTANT: INTENDED_DEVICE_SPEED_GRADE STRING "6"
// Retrieval info: CONSTANT: INTENDED_DEVICE_VARIANT STRING "ANY"
// Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
// Retrieval info: CONSTANT: LPM_TYPE STRING "alt_c3gxb"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "tx"
// Retrieval info: CONSTANT: PLL_BANDWIDTH_TYPE STRING "Auto"
// Retrieval info: CONSTANT: PLL_CONTROL_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: PLL_INCLK_PERIOD NUMERIC "6734"
// Retrieval info: CONSTANT: PLL_PFD_FB_MODE STRING "internal"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: PROTOCOL STRING "basic"
// Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "0"
// Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "6734"
// Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
// Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "none"
// Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
// Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "20"
// Retrieval info: CONSTANT: TX_CLKOUT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.65v"
// Retrieval info: CONSTANT: TX_DATAPATH_LOW_LATENCY_MODE STRING "false"
// Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "2970"
// Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: TX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
// Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
// Retrieval info: CONSTANT: TX_FLIP_TX_IN STRING "false"
// Retrieval info: CONSTANT: TX_FORCE_DISPARITY_MODE STRING "false"
// Retrieval info: CONSTANT: TX_PLL_BANDWIDTH_TYPE STRING "Auto"
// Retrieval info: CONSTANT: TX_PLL_INCLK0_PERIOD NUMERIC "6734"
// Retrieval info: CONSTANT: TX_PLL_TYPE STRING "CMU"
// Retrieval info: CONSTANT: TX_SLEW_RATE STRING "off"
// Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "basic"
// Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
// Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "true"
// Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
// Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "3"
// Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
// Retrieval info: CONSTANT: iqtxrxclk_allowed STRING ""
// Retrieval info: CONSTANT: number_of_quads NUMERIC "1"
// Retrieval info: CONSTANT: pll_divide_by STRING "1"
// Retrieval info: CONSTANT: pll_multiply_by STRING "10"
// Retrieval info: CONSTANT: tx_bitslip_enable STRING "FALSE"
// Retrieval info: CONSTANT: tx_dwidth_factor NUMERIC "2"
// Retrieval info: CONSTANT: tx_use_external_termination STRING "false"
// Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
// Retrieval info: USED_PORT: gxb_powerdown 0 0 1 0 INPUT NODEFVAL "gxb_powerdown[0..0]"
// Retrieval info: USED_PORT: pll_inclk 0 0 0 0 INPUT NODEFVAL "pll_inclk"
// Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
// Retrieval info: USED_PORT: tx_clkout 0 0 1 0 OUTPUT NODEFVAL "tx_clkout[0..0]"
// Retrieval info: USED_PORT: tx_datain 0 0 20 0 INPUT NODEFVAL "tx_datain[19..0]"
// Retrieval info: USED_PORT: tx_dataout 0 0 1 0 OUTPUT NODEFVAL "tx_dataout[0..0]"
// Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
// Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
// Retrieval info: CONNECT: @gxb_powerdown 0 0 1 0 gxb_powerdown 0 0 1 0
// Retrieval info: CONNECT: @pll_inclk 0 0 0 0 pll_inclk 0 0 0 0
// Retrieval info: CONNECT: @tx_datain 0 0 20 0 tx_datain 0 0 20 0
// Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
// Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
// Retrieval info: CONNECT: tx_clkout 0 0 1 0 @tx_clkout 0 0 1 0
// Retrieval info: CONNECT: tx_dataout 0 0 1 0 @tx_dataout 0 0 1 0
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_c4gxb_tx.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_c4gxb_tx.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_c4gxb_tx.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_c4gxb_tx.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_c4gxb_tx.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_c4gxb_tx_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_c4gxb_tx_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
// Retrieval info: LIB_FILE: cycloneiv_hssi
