// megafunction wizard: %Audio Embed v13.1%
// GENERATION: XML
// audio_embed_avalon_top.v

// Generated using ACDS version 13.0 156 at 2013.07.31.16:42:57

`timescale 1 ps / 1 ps
module audio_embed_avalon_top (
		input  wire        reg_clk,           //       register_clock.clk
		input  wire        reg_reset,         // register_clock_reset.reset
		input  wire        fix_clk,           //        conduit_video.export
		input  wire        vid_clk,           //                     .export
		input  wire        reset,             //                     .export
		input  wire [1:0]  vid_std,           //                     .export
		input  wire        vid_datavalid,     //                     .export
		input  wire [19:0] vid_data,          //                     .export
		input  wire        vid_std_rate,      //                     .export
		output wire        vid_clk48,         //       conduit_output.export
		output wire        vid_out_datavalid, //                     .export
		output wire [19:0] vid_out_data,      //                     .export
		output wire [10:0] vid_out_ln,        //                     .export
		output wire        vid_out_trs,       //                     .export
		input  wire        aud0_clk,          //       aud0_din_clock.clk
		output wire        aud0_ready,        //             aud0_din.ready
		input  wire        aud0_valid,        //                     .valid
		input  wire        aud0_sop,          //                     .startofpacket
		input  wire        aud0_eop,          //                     .endofpacket
		input  wire [7:0]  aud0_channel,      //                     .channel
		input  wire [23:0] aud0_data,         //                     .data
		input  wire        aud1_clk,          //       aud1_din_clock.clk
		output wire        aud1_ready,        //             aud1_din.ready
		input  wire        aud1_valid,        //                     .valid
		input  wire        aud1_sop,          //                     .startofpacket
		input  wire        aud1_eop,          //                     .endofpacket
		input  wire [7:0]  aud1_channel,      //                     .channel
		input  wire [23:0] aud1_data,         //                     .data
		input  wire        aud2_clk,          //       aud2_din_clock.clk
		output wire        aud2_ready,        //             aud2_din.ready
		input  wire        aud2_valid,        //                     .valid
		input  wire        aud2_sop,          //                     .startofpacket
		input  wire        aud2_eop,          //                     .endofpacket
		input  wire [7:0]  aud2_channel,      //                     .channel
		input  wire [23:0] aud2_data,         //                     .data
		input  wire        aud3_clk,          //       aud3_din_clock.clk
		output wire        aud3_ready,        //             aud3_din.ready
		input  wire        aud3_valid,        //                     .valid
		input  wire        aud3_sop,          //                     .startofpacket
		input  wire        aud3_eop,          //                     .endofpacket
		input  wire [7:0]  aud3_channel,      //                     .channel
		input  wire [23:0] aud3_data,         //                     .data
		input  wire        aud4_clk,          //       aud4_din_clock.clk
		output wire        aud4_ready,        //             aud4_din.ready
		input  wire        aud4_valid,        //                     .valid
		input  wire        aud4_sop,          //                     .startofpacket
		input  wire        aud4_eop,          //                     .endofpacket
		input  wire [7:0]  aud4_channel,      //                     .channel
		input  wire [23:0] aud4_data,         //                     .data
		input  wire        aud5_clk,          //       aud5_din_clock.clk
		output wire        aud5_ready,        //             aud5_din.ready
		input  wire        aud5_valid,        //                     .valid
		input  wire        aud5_sop,          //                     .startofpacket
		input  wire        aud5_eop,          //                     .endofpacket
		input  wire [7:0]  aud5_channel,      //                     .channel
		input  wire [23:0] aud5_data,         //                     .data
		input  wire        aud6_clk,          //       aud6_din_clock.clk
		output wire        aud6_ready,        //             aud6_din.ready
		input  wire        aud6_valid,        //                     .valid
		input  wire        aud6_sop,          //                     .startofpacket
		input  wire        aud6_eop,          //                     .endofpacket
		input  wire [7:0]  aud6_channel,      //                     .channel
		input  wire [23:0] aud6_data,         //                     .data
		input  wire        aud7_clk,          //       aud7_din_clock.clk
		output wire        aud7_ready,        //             aud7_din.ready
		input  wire        aud7_valid,        //                     .valid
		input  wire        aud7_sop,          //                     .startofpacket
		input  wire        aud7_eop,          //                     .endofpacket
		input  wire [7:0]  aud7_channel,      //                     .channel
		input  wire [23:0] aud7_data,         //                     .data
		input  wire [5:0]  reg_base_addr,     // avalon_slave_control.address
		input  wire [5:0]  reg_burstcount,    //                     .burstcount
		output wire        reg_waitrequest,   //                     .waitrequest
		input  wire        reg_write,         //                     .write
		input  wire [7:0]  reg_writedata,     //                     .writedata
		input  wire        reg_read,          //                     .read
		output wire        reg_readdatavalid, //                     .readdatavalid
		output wire [7:0]  reg_readdata       //                     .readdata
	);

	audio_embed #(
		.G_AUDEMB_NUM_GROUPS        (4),
		.G_AUDEMB_INPUT_ASYNC       (1),
		.G_AUDEMB_FREQ_FIXCLK       (50),
		.G_AUDEMB_INCLUDE_SD_EDP    (1),
		.G_AUDEMB_INCLUDE_STRIP     (2),
		.G_AUDEMB_INCLUDE_CSRAM     (1),
		.G_AUDEMB_INCLUDE_SINE      (1),
		.G_AUDEMB_INCLUDE_CLOCK     (1),
		.G_AUDEMB_INCLUDE_AVALON_ST (1),
		.G_AUDEMB_INCLUDE_CTRL_REG  (1)
	) audio_embed_avalon_top_inst (
		.reg_clk           (reg_clk),           //       register_clock.clk
		.reg_reset         (reg_reset),         // register_clock_reset.reset
		.fix_clk           (fix_clk),           //        conduit_video.export
		.vid_clk           (vid_clk),           //                     .export
		.reset             (reset),             //                     .export
		.vid_std           (vid_std),           //                     .export
		.vid_datavalid     (vid_datavalid),     //                     .export
		.vid_data          (vid_data),          //                     .export
		.vid_std_rate      (vid_std_rate),      //                     .export
		.vid_clk48         (vid_clk48),         //       conduit_output.export
		.vid_out_datavalid (vid_out_datavalid), //                     .export
		.vid_out_data      (vid_out_data),      //                     .export
		.vid_out_ln        (vid_out_ln),        //                     .export
		.vid_out_trs       (vid_out_trs),       //                     .export
		.aud0_clk          (aud0_clk),          //       aud0_din_clock.clk
		.aud0_ready        (aud0_ready),        //             aud0_din.ready
		.aud0_valid        (aud0_valid),        //                     .valid
		.aud0_sop          (aud0_sop),          //                     .startofpacket
		.aud0_eop          (aud0_eop),          //                     .endofpacket
		.aud0_channel      (aud0_channel),      //                     .channel
		.aud0_data         (aud0_data),         //                     .data
		.aud1_clk          (aud1_clk),          //       aud1_din_clock.clk
		.aud1_ready        (aud1_ready),        //             aud1_din.ready
		.aud1_valid        (aud1_valid),        //                     .valid
		.aud1_sop          (aud1_sop),          //                     .startofpacket
		.aud1_eop          (aud1_eop),          //                     .endofpacket
		.aud1_channel      (aud1_channel),      //                     .channel
		.aud1_data         (aud1_data),         //                     .data
		.aud2_clk          (aud2_clk),          //       aud2_din_clock.clk
		.aud2_ready        (aud2_ready),        //             aud2_din.ready
		.aud2_valid        (aud2_valid),        //                     .valid
		.aud2_sop          (aud2_sop),          //                     .startofpacket
		.aud2_eop          (aud2_eop),          //                     .endofpacket
		.aud2_channel      (aud2_channel),      //                     .channel
		.aud2_data         (aud2_data),         //                     .data
		.aud3_clk          (aud3_clk),          //       aud3_din_clock.clk
		.aud3_ready        (aud3_ready),        //             aud3_din.ready
		.aud3_valid        (aud3_valid),        //                     .valid
		.aud3_sop          (aud3_sop),          //                     .startofpacket
		.aud3_eop          (aud3_eop),          //                     .endofpacket
		.aud3_channel      (aud3_channel),      //                     .channel
		.aud3_data         (aud3_data),         //                     .data
		.aud4_clk          (aud4_clk),          //       aud4_din_clock.clk
		.aud4_ready        (aud4_ready),        //             aud4_din.ready
		.aud4_valid        (aud4_valid),        //                     .valid
		.aud4_sop          (aud4_sop),          //                     .startofpacket
		.aud4_eop          (aud4_eop),          //                     .endofpacket
		.aud4_channel      (aud4_channel),      //                     .channel
		.aud4_data         (aud4_data),         //                     .data
		.aud5_clk          (aud5_clk),          //       aud5_din_clock.clk
		.aud5_ready        (aud5_ready),        //             aud5_din.ready
		.aud5_valid        (aud5_valid),        //                     .valid
		.aud5_sop          (aud5_sop),          //                     .startofpacket
		.aud5_eop          (aud5_eop),          //                     .endofpacket
		.aud5_channel      (aud5_channel),      //                     .channel
		.aud5_data         (aud5_data),         //                     .data
		.aud6_clk          (aud6_clk),          //       aud6_din_clock.clk
		.aud6_ready        (aud6_ready),        //             aud6_din.ready
		.aud6_valid        (aud6_valid),        //                     .valid
		.aud6_sop          (aud6_sop),          //                     .startofpacket
		.aud6_eop          (aud6_eop),          //                     .endofpacket
		.aud6_channel      (aud6_channel),      //                     .channel
		.aud6_data         (aud6_data),         //                     .data
		.aud7_clk          (aud7_clk),          //       aud7_din_clock.clk
		.aud7_ready        (aud7_ready),        //             aud7_din.ready
		.aud7_valid        (aud7_valid),        //                     .valid
		.aud7_sop          (aud7_sop),          //                     .startofpacket
		.aud7_eop          (aud7_eop),          //                     .endofpacket
		.aud7_channel      (aud7_channel),      //                     .channel
		.aud7_data         (aud7_data),         //                     .data
		.reg_base_addr     (reg_base_addr),     // avalon_slave_control.address
		.reg_burstcount    (reg_burstcount),    //                     .burstcount
		.reg_waitrequest   (reg_waitrequest),   //                     .waitrequest
		.reg_write         (reg_write),         //                     .write
		.reg_writedata     (reg_writedata),     //                     .writedata
		.reg_read          (reg_read),          //                     .read
		.reg_readdatavalid (reg_readdatavalid), //                     .readdatavalid
		.reg_readdata      (reg_readdata)       //                     .readdata
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2013 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="audio_embed" version="13.1" >
// Retrieval info: 	<generic name="FAMILY" value="Stratix" />
// Retrieval info: 	<generic name="G_AUDEMB_NUM_GROUPS" value="4" />
// Retrieval info: 	<generic name="G_AUDEMB_INPUT_ASYNC" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_FREQ_FIXCLK" value="50" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_SD_EDP" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_STRIP" value="2" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CSRAM" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_SINE" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CLOCK" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_AVALON_ST" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CTRL_REG" value="1" />
// Retrieval info: 	<generic name="AUTO_REGISTER_CLOCK_CLOCK_RATE" value="-1" />
// Retrieval info: </instance>
// IPFS_FILES : audio_embed_avalon_top.vo
// RELATED_FILES: audio_embed_avalon_top.v, audio_embed_cs_insert.v, audio_embed_frame_seq.v, audio_embed_sine_clock.v, audio_embed_sine_gen.v, audio_embed_sine_lut.v, audio_embed_sine_ram.v, audio_embed_input_fifo.v, audio_embed_hd_packet.v, audio_embed_sd_packet.v, audio_embed_strip.v, audio_embed_control_packet.v, audio_embed_video_input.v, audio_embed_core.v, audio_embed_registers.v, altera_audemb_reset_synchronizer.v, audio_embed.v, cao_fifo.v, cao_merge.v, cao_avalon.v
