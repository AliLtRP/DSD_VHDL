// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wf5Eik+xE5AMLyUJ3Trmc67Q0zne3AIf12qSlGnWPDfwgwQIDSfxTcPlo9yBbCf4
dUIQvp7d7G5l3zXlnxG1gF2TmUqWkYmMyccU2t9S/Eb6xn0VzfjJyImXD926+/UK
rqCPC07PUgJUnXxWnrUXjj5Jn790FYhhmNMZgS75uTM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33056)
FAJf5SgLcRFsOd1Ouu/nm3loH6ialLnEERCvwYfxQlkz6Bjl40+63I6+SWrY7PcU
MJO/1ps3X0E0STbN/dgWvjC96jUUe1leLUd9YGt89SQjJPJb32KcTJN8TBL/H3Vz
/nIodQugSLo4HA5rTo7wjbXOxy6S73sIDhDQCNAgsH/5v6la2bSejklxLNReanVv
HOpOUtzD9KYDSQAWA19Y2XcKw0hHx9qQaRuW39HuMKFVUBDdd4o5A8KTEX6sSwEg
1Mv7C2Glr5dv63CthBWsIv8Wr2PqdgMWu74u/oQTji0eYUCYSLDarP+AypLfhYBw
SM2t5+z9tdxTv1bgdlt3CrWZMnu92/MeHhyFEr4YxIHGmXxNRNz4+SQYkNRx70zx
h8Hl3zn36/Sh/WcIFgcSDiQ239d/y0nxBsVtGrBnu53XU2ggSwFAMtU7lr3JOKUz
mVFhs/+F/2iVlE8PwSBjcqHN+uZWx7QGQmsQ8WXFD5K1aJXJ8G0Ukwe9RCs5xJ8g
lxojbOij6IPAi7kwzifibYkSFoIo8Zaum7C/l9soKg4v4dtqN3hcMeq0JrkMVEyc
L9MJyc5ukgut8M2nOGqdmWUzxhxyp2rg/9/dh9kABrAnb2Jqj8t99vT1YoD4laRy
SiE6aBYqDI/MDfoNvWgJFNktjP35bvzQFt0a7zZuUesJuB8f5cv/nK2rhk030fpm
gyXPQHkJeaeBBdTVq3BNbgsZwMvgG/i5/23ogOF/fWE/6xFWhXzsCV652W+Wxse2
/nK4fsrKg97g0/WFYgdtBmFcxlBtISH0dMtTuWDFbmv0GTFj4LPF2zFeZ7Tk6yYp
EikzHdyaLNL7SCeI56gK7d8BDraBau+pKfKA8fcTm/5eqIMVDilk5SSbKBBHE/g2
r5lB/Hx1NOs4hKZOhIXXmQz3tr1FGYeC1in2Q8kAnATab0d8O+CCoAEqs/4GnkKh
8YMiZhDRLmKvdAE0ItLvxGbw00RlEGpBrS3MZDc/ALp7WuYgVRJaNLjTWqumHCle
al9EKFd47kyyfbzAhpjNmu41x7qOj7D98dj0f9ZfePgk6xNM+uyGijfr2DC6y9K/
WXwzb/FWUyFyu7FgEQmGwbFQAu2KjmiVB4SOp/UyHX8UqN8uBEj/6yRv2n7i884s
McVohA/Og3opkyA38fA29yAqz8O1VkNUkBucbJwoDtVf3P9/bPGiypZG4qu2zmFB
BmRQyFpMp2PNtVnbU0agYld6tSBj10VvrkKxtBfiZHluSGMvIDWXMlVJ0IEZwjmc
xuiwGFrS0IXp1d9Qs788v9OLIpjQ/0LqWwRPevELiEKicR2cWIM21YegDHmj8zGC
Boow1p62UzTVGUsZId+22nidUVluDRQQv2UQYwVeNmd8CBKtb9faD0mEN2EVpnOB
vrEIRmpbeurEv6jDmR+CpbD29AYV27iFK2PjE4lzmZ3gMHaYYD4rxbDE1xu0rXy5
0hsmVUFLzo8VB8FO+Fs7lLPJJTZ526kR9djD4GxFnQHkxNHVsxSAWbw4u8up2fk8
eo/xKGFArARGsONwvGq26Pbl2aK3x8FM2265EfgL2c2r3tEV3JVeZWpINUVRSnzO
lwRndwftdZ35LUE0VPpxAdu3HGgzpBhKcmVyreT1bvHPvZWtPSCNn9u47eV1btSJ
g4H23BerrRVOw68uVQ+FgCvFdVeTRv7H+hCtl8FOozfxsd7UeeoQJ4e/yT5U4jzg
HKjspvVmXGHBXh8qN6fnk+GUZzdWUhbmLm259d/XNikDt0QZZNvRu5i4QM8uaZDU
L3lKcXUYpEwGo6B3qJWIfX4rQy0usK9UjbKZp2w2Zj2W6zkLuHwADtAk+fsluCdo
k77k2YIMnxlGMDyeondyg2dO2QqzAKChvNCgbeJ+N2GQXnfQTxR/kIENxBjFZNlm
6W6Bow27jNtkNARX+7kp/EWT8Z6xLT+MSafCb3N6mGdJCh/VH++Rsd8Qd/i+/osX
cbRKlq+ljJyXAg3ILoZIrS+b1vKmGpVzUzLxU5VbeykE6gw1XrvDcPU2qM95fiRk
xALMsA5/yfSiIwGgVg/U1vHvOE+LlBpF0FZkijLkevvgEGJJqgbsf/Bpv8LXwNce
QbEqDFzhf/+RoXyKkNjMOkkee0nKEnPyW0/SS9p8i7gGCz5agcjT5dUlS7iFQsdN
fLqgNnxD792UW4popuf+waXL9MHrfGTyiX310IrlFmp+k1ke9UXBEvO8mXzU+VVu
vs1FTfg+IBD6K4zatJk2jhlQOpX3xCadd4bpvoip1z7oL/1JxWQQsYzaCoQpBgvK
vOQWAMi0WxukyqdDAAMWqyXWgWTE05Nk8PFboFKOjcDFFDyQXOpZONJmi78r9JrD
v9BfVzgF6qMb04SKGQUGCtuW4bPc/k4fOHV77Ev929fKo5JKGsP33clFllgHHq78
ab8anMtlrLNjzb/lwWZi1fPb2/l8YrsG4C7zFp5+150HpVtlsidm3hLDbwQr6Yr3
YN8Xb2F179RXaJZttRQTUgx0UeM296IGifPBkLFkp7k7zqdOYxLJ4D/V7cbpqBk3
GgIHi/nqEmuW/HSZgK3ym1OCQRGr4sAnI6rQkHX/uhlRnhlKInJgtKimXgP92KCQ
iNFHsR7tI7YN/S5GH9XqM8ZCO/ooa/eS61Yf8mUO/+HsUq4ST26WkLu2agfiUwF6
zTKX1bavE6ySdCvU+s4731Ds9ld2mqVPbhdtQPj6Fsh4S2X33I9apwoQA3z61maE
Uze90EmlCeQFZeRBXKmluts4PboRaGpDV3EUOsetobhY+dbeiqBixXe8D/xjfpfq
FfcPNSMWsDcVzUodebjDzjRhJ82TcTUUOBUB3yTPu/NkNKy/wkiwfumIrB9tWINa
+TUYCGrp8FZQUkNO+IvjTLAI11EKVXEraA2K15nazkOX3i8KAPdHEKbaJQl24BYq
7QrSt0eOeWyFy7bqCXNYF99HtcNmKdcIDlOU3x1o4t7dRUDbGME9zhPuI5FBUhQj
ynTXnNBtcUjMmORsgKMYtyheEQdcfSnNcDSlAN9/PL0d4rgzC6Ch4ujnp3qsjzot
YgkUFFlXoLrCMkMviQ9Z6cKQF0g7sSslDSyYRbqFZGPpJImIcJDk5eEMFHP+6Fe0
eXHvd4Zjvshp7MLLa7uUPe9Fcd5GfrHoOYxwXt1YylEu7vpYrMN0HVsfKjGQkogk
kt9O3BaXEIS14nhcFNGUAEGU1RSqcDATbqUyxD+7eE+aG7TdfGTO7GP9La2kRVZt
8AWz0t+IhRTApVO4nOtqBAXLq5GcQPhX2KawIPLQbkunvn4NyGnCrjJqWKnVTnv/
AUVn+2SNqvYKVePweHnwrHF07IYCnUiCz0is1loNFFMCI7V/XxAd2WhCGRyGSXws
H9NypC8nUvFCcv8ZpR1XdEZnNhuvobB2AiHYhxtASghYPu8RcZuCXlDMYHSmBorj
f3W28A6dZThV4KG1khDEvTlh2kvTUL1pEJEU9rh+hH/ekTBqUm7mb2KQ65Jz3/IB
ojk0zSDJ/u+cXN6zczaFj0Og6gcO+9kNL3P7TLI3EvKwSfj9g/ZgHnIKppmLdDCx
GS9mu5TBPJZS96y4l0WX5lwRd4nhI7ClDFRnz8ZXNv88q3WzE6NwjS2uJWJI1b++
P91+EQ5Z+Da4HVNOW/dKbwPdiaQ2NIHPku9hwXCWGFqeFHXTk98fSq8S9H8SEflV
hvYdFsNf/u3iadJByQu1mzKaivKx+yTkucks83xR44zPqcXYGfOyu2cBuojFAxdp
58+kCmst/skOyzAICZ0hYw4ve6xTRN51e/iBX9PmhOG7UwoNL5sTkN+1f75Gwlz+
qxL1X60wWqSOW8EDFqD2aSumVK1kk9F2X7v8+sZpZBDqX0zFQNgFAWOCRjL+9Alm
QSWaWkTe5pQCoBVoV/tNhRk0swlmfJT8OZONVviJ9lMMTIuEiDhnE1ilB0Qb1QJ3
t25zY/EOZlPJWLlZEvvyMX/c4lPfjwOQZc2GIW13DHuHS71B2gJJKAu+dOtmRl4j
gqxuPm5le51gBEHCDYX572o6TDCTDEA0NCnkpcpmVKWQlMZcvDmikke7YESdl5nN
ATdFXKG/saNxH++75ru68fCwJ3AnSrF3iBWaDANOdtYqN5oidf1yqaNGMIuThT4v
FFGbzusToi2mhA/dpHJVMxsvQ3FzY8U4ZouMX1BFa1Jv7bR5LGeY8lzjJm50Nd/C
GyzUgaS/lMu3nxiZQKRemUJS+403DnkUzDWupNYtsRdzlKPs4PJETgjGD1QBPpxh
AK644S1LhqfhaRFCUIkP4FUBYLiaMBqXLnkjKPRbAFAw/M8GWlpQZJKwgvvS8et2
aaCJKXU3bhEV/VuCuVR8vy/I8l1pPqW42yXN8KBPFsnF2RYTdjUvuKv7sLFhqpTN
YT0Y+575ZkW7NdXabsjNHCoYfdFL7ptUCBw956CVgOIISaj2LGx4JuqMqxdG0nLb
LPjja//83lzS4xyp7vSxsqNQT6S2NIHt8Ryvx+knyOw0ClEStFh2KlWIFD40AxGz
jWh0U4coMefKBQAxWl9kjiCgJYc5DgJUXSz8KryJ1gonxrjTyJE7v4Io6L5P4raz
xx3H2vfOroFg9Htv3oRZePDs3jhkvvmgm1zivmK8IhiWd3Bx7MwlqQIz6oWmgmz1
jncJLpp13UUnhmZw0MKSsRQhlSWzAZpG9/5KVktfWzLin+9SYpALOh3+sJiBbobP
/8pZZkveW3vpJcAPL3dIG2ammc2DWzGJJNgs4RQMa+8+mAW/3AyvmgXPnTARlWSg
3TL094llykzaoK2CoCWqsuSimwA7relRwiiQmSw1RVfI4opY9FYZRQdhrNHjmGxA
JSvPJ8IM4UJoSuoUT9NrEhB98COngOC8NHV/2TyH1Xq3cYXxOl4brmoF9gX63ylD
eZctmLoCp19LZdSlsAw5KkVkTs7dicx+uPDqGJLqMfNylmYtfMHI10G2xpfWQ0ni
jJFGJnIB4OVIHEHzvSMz+aW6gBNHp25w3fw+YUs1DRO5RJWyeo0WN9Er92HwDvv5
6y3JH4ENmcP40RR/ZDe2WKB6H7PqI01fbFO8Zf02ATdTN55QE1alEZOG4zokPoHA
9EzYgX9fDOpdvCTnUPruv1tEZKOdQvRJJlpt/Txx3ujHy1hJGjJ26SgPTPs8XpiE
3eXMB2nLsYNYdDGOSASFRSp4nmmxEpC+EKtmq+hmJXVoRiMETZkMyLE9IngH85GB
5nFS5PeKg8mXcfmXgbzZE869GFYPzOxs80AOoi3G10buh68hbwL1J9SkJN0H5zYk
vYdbwwzTb6jiRsLXFycmCvXNwRS5Nq5M20KKxNf9ayIeHLRD7hOkCnBj/Q/xOXxb
A8qq7teVYu4+N9Vunvia0GZw1Mo3c9pTbc+pz+X6epVs7Y3w+dN/Ynk1GEw4M5jx
G5ZYFKxbLmdgKKNqWFBiLq3ZJlKv36N9M+SALBu7+FUwkMDqxbAYdXEgJEZfdMzd
jAtt1AU7xYoDLfFtH+K0JHb4EyUAooqSKpttHTUE8rAgR87eWoUqWmrGVU4CpFbo
xE9amCFVnpC28tlcW5KVc0u+wCsqIQS8PJCBG4bg1TKcw6XQ4jQPSdf+IYuhShV9
e4hmlBHiBWGJXGDokWTFGnaTy/w9WUS4AvhsSn45Q+ZJMwIeEu5ZLqYdqAWimA5k
eoLeaUFCQM3cwpQYfGFRHNM9LC3RX5ZpPbM3Wtraq9cDzvFLo8fCWB17Elc4f47K
Kc2z8DcAS7LLE0DjaKSTxH6yy40Cb0CRcEYmNTyl/dfLhWDOIUVeDUDDTT3ImPVE
germv0U8swVO06GKhWFvu9GAjIT6YKp002RFYDO9tdypQ5FQyJMjTKVWfRVoH+3f
2MdFrHRewSkzThUajrpaiCW6BFHcgo1AG83rJpR4/RlAPsaZSmqWa7g/AKOSuUSe
JN2bF8cSxfg8WS62FYXyJ5KGWWZIwo3XYlfOVLzzJqBU8m6dQTPrO53zjN/DnFXG
hh3hULYqWGkKCt6bfcgeQYT01lRSXjkSE0iy5O9mYIkDQoZ8AX0NlCp7BYCbQN/j
pNUAUiN3My+t7AhFcD4ZxfVps6BTFUeXU9CKnMPi6AVhzepOb6s7wBzRyu6IYiGN
dHD7ordmBAhBvfyync6kOauAivCIlUCKvDmykkhqoNhucrzpr3P4F2XsVKLrPM33
oBcQLSDKatC7OcaGHcFs+DGV+KjUwm2uXUhsJ0Md5//7QEffH7Z3GrG/VMx4pspw
+0N517wJEOjKMH/Mp4u1jAo+ci4/0BT78YTYhmVRbDt4JdJsIGgli4W2PnK0oh/R
8GzFVVQz3b1Y8INHCuLDp5AP1u7jznsWRNC1eej0v/rKo8V53XKGawS0Gu+v3o/W
cLyWEOxBlHx9jKQR9jB6x5Z131mi/53wnPTpjHyHXNSauhgTSBehdhJtwYuVWgrM
jrK/62+gm4B7gku1UECRM1EzQCpkhehgydpKZG3KkjN7rlF4+gMdT4lryBQoZy/K
jozZ7tnvspMz7eTSBgraauZc/cOuFSji1HXc2cuINkcbryIkxf//7nR2WfDhVDGA
kQm9a1yXhgJiAncU06Vjgzea9mvCDvZn7YNQIgGInSvCQG8qX7QzP8y/SQcPsOJk
8qi6bs+6YudEzcQMnpIaJ5Js0WMTeOQzUT/PADfmV/rlAkX+NpneWkIHm0tywL4I
uhuz3gSLkBrloF8S6EpSd88YKnG2RdZkc0gczcolX8aI/4zcRZovToLhH4w2ULW5
zOhPjV3RrmaM8+/fd/Wj2eqk59sIGyk00GbUFWUzH8b0nQHg9i9AqzJqJfeNa9Fb
tc69J1yt88tpTuxIJDsz+EwdX7Ge58799rvHehQkZdpUnBE3f3kzHA78Q1CuFzGw
CrvU8/+PPK/POX1A50ke5UYRdrMkEgk4Xyj2K+tWuvqHbArCtvlIZLpKFLmQkA1p
Ef0ttpALFmzMaZtG/F54TGl/84npmicsnZD/GsptzlxHImBxrS2CV9wCV3FRFmRF
JvMfDbS9qjdu1ldpqNaE/xcQMEeOGD4m3qWBG4J4XHrsUh8KSOmHNyCBH5Y34/NN
rIUh+lG6FpiJ/eKC5TgwiHjaIv0CCKhzGrYMMmFVlGtex3UP4FjDoe73El88/jte
ZrumlEJBM3UH/3Z5zjpJn/vBzTu3wk57wm1iw9APq3ezFSCS9eHzUNbXhZgz92z1
Zr3vF1y2zbaAGojVxTD/ofcuFOQw5iD8XKL4HX1VgPXuJPhiyDGCSCQ350zmYkzK
UYUiRvIhtNljcjWfjL9Q5MBgPCOpLYj6CC2jSOVh2S4/ggdpA1bM+FRpsN7PkSO0
xViu/NSN09UVKhNElJ+ZshA13qWGRz05D8UHaPCfNwvezEcTkq9vBfHB4/MzK65f
TebeHpfnbdAec1dMIYRnSMMgZ2DztJ8w9eqbxb0T3FRu4U4YD3DFih5YkG2rRRKk
qcrsRYQbINgYTJQrYOAfa3cQ4ii9RiSUOTkoG5pr47W/oo/w8TKQIZtIv48JHQxI
Kr3cCzqBLxyw/7WbcfNUPqhpKwfxdE1AZCkTlUJkqffBxTa4pnuLUiLh0lRcqnLc
UQ6cuCniW8axcQL711OlLoyesJx59qpv8dtu3TKuJGLIj8ZBujEntWaPQB1qOuV8
egmk9hMbS+ZoYatehWmFjmtzBvztUEOWtlVr3mgzAxwKkMSlzKvCRXz+2BbDidRE
pRBG3WJLvHjUORR0VhniUsUSK8qzl1yrTAX6EheT8uSKPAe03Up84tiVbdDV8HcO
5Xz89s/PqA+10MCdovTS5iVfXoYkwYBJu4hH7KnNHe5wr6F+9SRru1f0uzpEHeJg
2OILbMUi0eLYYiB9L3ibWPswzuyJU2t/J04MKVy1bJDfiToRJfj8mvNQP+TEdpNe
/f/VnAfkz7eJ89L04N3CddBlJSzFLEkOGb3lfMuX/yGzYAfzlUGdYvARVqA5kvZJ
d1LDxXeCUA8fe7t3+x35l+pve6qahimBqd1Y46K0ILJQgsN4SInLCKpsfllAoIq2
YYzV4OVhaEzrEUxnm81CeYLppXk6xjrm0tMjfBBx+X3uE4xPToGKS6iyASOLrI9/
10IeFk90QO8S9YzTLGrA1CJyvJXdGgc+MPmzfLMuaj8Nh9VhGbLoIJzdQzXT5weI
v8mVZqsdG1YTqZgDY/kHNHBB/rJXmrUccYwC07FeODA4xpOkmHEXVQRE1eGyzlzF
MMziEsyBH7lz/nrxmohCr8F/LYKh6cyzv4Qk0Fvg1Rd+z11CSOS7lVSigVofhumC
EEwxsdybhS0hl5HGp8v1xYYLunyhPHauiftC35ACRvuiHzJmLmxPbMbLNLcF3kWh
TXf7oW4P2u4pQ0RX/a7T5ui9bFmVowcFrdwgIeqA5rHUSZ5KFxlqT4OWPKd3IsZL
AujOTyuZJpNa0kYQJSlnXB/3YqgCsxnPhWAxt4LXJZ3QTFMtP9BdukYQWca3jR6h
TJmwWYIz+C0TtHnI6I7bmVA2OwOwGibpqMEk3uYoEiq/j6omCjQk4yodq15qbiNy
PEO8ZrZhH9nFjlfw81FVakOAYVTF/ow58I3Ss9RsFRcH1ji304aAUAQvOWpr6KHb
7p9V6SFVIJoa3Zu4xkUwny8QiZKVdsHLlOcSRKUVzlS/UF4oU1T88GMUpS8Xo5vI
L3bKlhVedHEWRyKFbBUmFOREvZiMkerbU2zf1p0DvjPlLv2u4l3ko62lmAGwJhkC
efZhTvr7d6y2t/GkoFEch8lRSPmaimyLzNYaSSRkDQee1JxbmED5d40liib8hbgi
vsrRu9wk5azZZG0Z53fKDyjU/Pd/qgHG9avP34cM7ZBsH4bEoWjU1KbmbBHFpNVM
Om9Z3WtEuZk321BACXcuhYNynS14LC2c3n9QsnKOnTi61fUDSv8nF/c71S6EEPb2
bny6ZE2BZwZlFQxBYHKHNJB94CeWirlPXz++bwoShXlIQJ8atNlPlKCjUiuvnYKZ
AYeQ7X4MS9TNG1zOXPLfDEN9vXs2GyO4SN+X28TJZ6Li3tSqjzim0y37quVK6XC/
9x/pLs9hS1hEp3RP4foIB2tHszEtdH4C/w14tWkwmrMghpXJZSP0EKEQ6Pxl6Xo1
zWdHFz1gI4tpYtovK5fZBbkYP1u6OJ6woimrFmHCqj595wYIWtM9QmD6+DYvMT4K
AlgseHTgLnGZLzZqHISgG1aOnGrMUeGOcDT1oDDKHfZ2tysKr67WL968Xw0stlfs
/WlG4/9GoRs2kjK7hMuuIRsbySoKqlw+OaNtT1Pcw8+9AX1+he/nxALNeKhxZTst
MfM8LvlsbQ87rKw4BuLckgTONg6MgrOox7at6sNFJaubHtyWCL09VrBUakDLPj7g
4ag5edOvHzaPet7bszRD8LwABS1RYplNbhP088S0b/gq1SDf41rOkm1eHS8jr/S3
4M7Mwi5UGCbU0MT0SqM8/6+plgny41vmGYZAhORQCbqh/1Rg5x9Kd0prsWmc/QIx
wUruxHDOX1kp4nDnE/HuQ1fYF7chQpndBHha9Gw/m/2eXf6ZdJXTGya+CpnwRP/q
d6xlTpESwB1w+QjzsEijxg2AsnWZtWziVMpxKC71djkFVYZcb20NciB/mvbvBCoA
mHE+YitBOI0Iz6l25TYIH9Kuef6XxhkFk9zNRV6sLu4oS8rA7QWn7j8CNQq2/QvS
ZbsgRhew5wDi/Sj1GeWoUI/z2r1o9hDAKGtlEQtzqd4G+FOmppfUPEVEqYCXBj5Q
LTJIbzoTUS1HmJtMhatUkuxX/7/7IekUCO6T3uQvhFqrIEDzUDIE6MwjYQLb4weN
GsdQu46K7QtjSjFueMwx1uVrHz4fIE0gcIr/GoEYm7v3AGTAPCQswWh6zcbc3PXS
1Ee8u8Ti/ByFBO7PyWmHvNBHXuEK8zw1+D83Od9jqBCfbLmtW96M/naN5gQeORsg
C4lSFmr99C2JuNE0Qrqyuf2aZFiHaqjr+6DSlRPFILT5o2v5bebmjr8t/w5/PMX+
ekHbiMNfZ5AnxN3i9hmBBLKXIgoJ54Xbh1hci0EQdOSfgVlMkw4q3IR6yIdobXYL
yYjvkzzFZS/Kx4GiuHKN/Qom1+pQYJBPKoJJy3jbGOWguWsycjj2slNRrDcheNNZ
EdZxNdwyKzTEYH35odIv7dwd2eSkfmszeqHBVdZhe1gm/aARkKBqEp4ymCsodENt
FLDRbL13MaPCAo6l3EBBSqzra5k44aukUCW27VLBuBZ0Y3M32ENKnFYx11+fShCj
1C4QGcrYczM3yD/PnCUJfEmorjSqkpkSZ5hUU8lLFfxGvCgFp84KkYU1CN2K8Hb5
ZF+fyiz7cuuTKqUsjS+a6O/U7EhV2rbmsVWr6pfK1UFNRW2BzaKuN3tg5o9EBA6I
w/3AVqd5eGyd0DVP3Nt/G48XWeXcssx3IXzzEejpfT+o/OL7yghRzyNHr1chFQKd
ypK3bzjHXgJ/dQCpkuJO9kY0PtFy4tj4xpIzrPygSpxZBiXT6qX8USPL6KnfeLc2
0XGwKqNCZcX8fZYNN2JyZ76+pXfEv24+I0w4KK2pq+qmbsyA3BIOANPIt7oCo0Pi
7bL4yMFLYHxHPIp0gcIvDr5vUu9odQ9g83IpvC9iNjh4TyzzGaZ+itP8UZuAXQjx
H3M39XSYPOwzXak3AjMoIOEgYe3hsvyi30FqMEDyavcN+Cnrr0Etf1Cof4s01FHs
fvR57zMRqO35itQGauO6g6a1TmSUOTjpmAPvKovYUSexaPminUYtIIYSWlG9K/zQ
HIZwmmfCdTwYKDtiuujVPpTERvW05p5F3vQ4MlyidyWOFahUWdFDJzxZh02/ic5H
pyCnxiAQtDd8FuiXY/+u9/rS9u1bIMS3iddbQ3KwWHwAOptVgxM6/S19zB5ZVOE1
khyvdqThPFQYJiFM3SgH0t/bnOlQFEx/FF/rqefB4ATFWEbIePWOSucHLuTqADm3
gzBRG7X+DxV82WfknC1SIo8RwKQJNRvV58rQUXbL2fmUaa4s2jm4yTfw0diA4RiY
8ZxsmY/DfDYBnljlbKaC6Kg8HkcIgHh+gZjJaUcGCdSLNEgSCFI6UJHpKbZHKVHN
RjGwx8EQ+hBKegACBBQ6YAu4a/e9MMIrISZVyTF6YfhPub1kEub53KoW/oOn7oqL
xR66cbWTO3oXRIv1RpYd7MKOIMn4vz0mAKIk1Z3+cNgaBpIp48U1H0EWqF8FNX2X
JLhdRWz+Ycaq5Z6q6RxDkM0Q/jFO7E2KF8d9ViRk1VEUH6BvTDovegA1c6pVo4D8
cm4ay/DpBBUBTiypKDycaP+/4U7QzXtJCTYAbGG4RUo+i1pSczV436rG8afhepky
H80uQh/g5S8Zn5biZ+xZUqyiW/YnPWqsHy3myw2ou+TlVUIcQIZsUiq+5rWeXTSj
3TKcaly5vFMpJ43XM9xcnjOCzOC0SOu/wxTguDeNePnpAPaGDQpesOqkXa1lay/Q
X6ePbI/fkProj+VyOEv3okq1dO7dvgtHd2r8DmWEIXsS1/ZbGvdLJyLj2WgMQjMU
/0WF/KQfu0rGAF5OgugsZc0mH+zWhfrAFoB87Vt+ALfrlg8L1iX5cQUJ70/isqGt
p3l8LOdsbPA4hPdspTI1bZWUKluSMvsXWJbf2l4JI2+13I183xSjcPH5CK3YQ7Om
YBlWwFNnzSTLiY96dsJXFDNs2gpK7DIsippmDAu29d3mbm/KIQF8cFWPSfqfdvdh
ZvcWo0JhkixIFIUxkIP9UnWIlYjauVO8qPyK8DFSZHueLToU6oZfN2Xl6vaibg9c
VsU7cgACNuR/txK+KqDUvxBNtlLOVtsmesbJGBzlMsEzpjnK7mQFXxoINOfp5KA9
SLFZsT7CV5sXnNBu4wykTY01tAfCYZpnZNuUSjLnRm6q4rFTxTBhKazMWqv843gs
g037dXMawZ4rVNCuuKS2Dt2KghqbABbPMipX619kC0imRAlkoXPJS9XXys1njlto
CUfuyJaURxNYa8F8kyCdxoiL4V0MHnQO0h+Ih/KlLrdPhF9JDUdxCnhrQ4WJm2RT
FLy6YJhmhKPIJFbCD47s0HvuebphZjsnbPra3gvaTgAeBwRG8zKBCm5mI08dU73t
UBRtROiFrMYJ+H5+2BNmWpCvmNxuOouNjlCUFLm/FxDLv/L2kIyfnf4tAGPzMNhw
mznLauDhKzi+1uzSFgiGKZKkwGLoywQBhb3B4jk66U+vvBxp8qZh3NyOf46MAGjR
soBxU9YGnj01lFw5zNCrLJ+mtkgxE/Rb++/UqOVVXs/ZAMbOaomXOyINWxIByvLW
vlttoCeYNv+361hrG+2PXadiTu9/CkWsgMFh/9tzfd8es7rhWHxC7R5rwqbrBPKd
TdVaf13W01DD2Xr72KuPa2Ov1ozifdmCwFgdysgS2KlXR7MzVZS1ACOPoSzFpr4g
y3PULxs4NGXmYkJmpPE7gRVvtrjlVSgTSdgr0hyEYGU0pu4FDfA2K6IOixweu5BH
dGOmksMXeUZSxHCC5RVStcVONksdf/wA/JtFwsVwdC2tOdsLDKu1VmS5m9BE6Gar
e+GXm+UAOOSPJ9vK/5D86pzIBn9nrB2lDC2N/8SZvX8QILO9JSHagNmxnnJlO22H
zO/3IFIZnx260p09Y0kwA5zyEYQnn6+Yf9PgXy3LORvmFZ26/3E8fQYuW5/V2I3S
s9QzGlbO9/zhNlmugJQXWo64IOq9r3CJItS6sxBux3Pbu4AmHFZF38liPFHNdBq/
DozgykYYURnMe0eKxOXEeehgtTc5zXKW6FPrzGr8pdM5eO9LMq4pCcca2pQSHaNn
1XXkwOJ9Auwp1H11Sxz3GdmqiAPYqJt4xYISGi3/pG0VHTbSwHUrotFdt7WC3CUk
WngNi32UmHjOm+hYMUsDCftq34FwEFSnKT17AJMZxf4oT5YrWj7NZiI2mudoTgF8
jzOYiucn17S4ddunIHIRfv+KYsqnBo9yvRSx016iFjx6AgBgDRj1KdChk0pJCLEM
zmpPkoZqfWuv91YtJ/5vEvljGklcU/ZOR8X4zyASB6he/oY7TyP9zIIZmOS5NJtd
l5ABJOtMHaPGKVRnubxmtE0aE0/uPL3eZbgZPeHTPfSh2Cs7DjiFqHJ/PrwmY2/0
y/Yl8Bpi5RumOKQw9Y5NqEEs4fECgvfU9N2ecrePjzSXT/vo+eMbzS5gafRdmU/X
fcZaPo/2v2YRWHiJtw3aV2jamRsYcezBpcODfE4TcZOefCTx3Wr21yguP5sHnGra
/Tn/xlsYpms5Lm2JuWXZR/4U8kFTKaCCfSdZdyq5kwtNCLrjfJ5sachM1IFFCeEm
eXgTxZGEHNh8oWmjxEVnTRAq+APDuxqovDOcJgwryIxMU7CS+Pw9b8KnDyXJO9WN
BALgdGCVVCZMdVTDtyBiuQj+G2FNoX81BTiX9BgUMmF0ROlTe1DTMi7u46m78HuD
MRG8fbSLjvR5RSYAZ6qLZBn0HL88o29Yy8e6ULhqGV3AUSzEXiu0Fo+/lXRd2H3J
nPo0JBYMVoxrldi+O3/6U1+50+NLnjHk3X9GkJNQrwU516MeEewF8k+mrvlLv1p/
hiTX+kmmI0V4orWJwMlo6zXhN540zTcw0tuazeAPrx36LKChXJxU26MrtMhwYqkU
H+7wMmWnf+h2oxIylYoSv/OVlVeaYGVKeMMdaPXcGXKnZYnNeXx7OJEow/xJ4v7e
IhsOIJPPBjeVVdrjKL/1EpRhRHir08tYcVgkAPZrWq0SyvN8oHp13U3tXMiqFViU
Lpwzj1jaQXWnwYWeDLn5bLgi1d3DeC9JjabP7RSyd/IsowcNFC9yinQu9HVZTzgD
66eKnGGAwSBZHNtZsk7Roccv5Q2oh/4P+1q+p3X17g3KpLOgGV67bXYmjFqfb+Lx
FUkmR760p7el+t4DLNOBfuw4h3x1sEHGgNrEe2J3rSTATmy9Q3l/HpMJBRaosrsZ
8zXhuEJRpsnzc1w+vR1gedg1+EuZMQ+HoMOgBfxcCs4QJA7i2DsT258ybOoLAY2e
cCfj9D48ms9r0qNp/w2SqJReHDFyM3nuJfwSYmSd//vrfCJ1rXpQUkNUKsJH9U/W
MYebKa3JvSaXgGlElh6+4jE+sSMFG5H7vOIZXiln2WfvjY1PZ6VXApH2nFJ4+Nk0
z4T4GAUZio6NCjybxGaMBtGPyBQ2LIhFr8VAC1T+DjbXK4eh4NODnjPW0j/t3eNc
wrb9g5nkdX8iD7V2E/DlP580NmJ7BgzxyuVWjaHxCtRNQtzl1LrpaMy/ANw7Tl+O
MwEt5vhN64/+ji7htoQT8ezSJu2lezbZfbUVzAMAMjXOCLjJDYdk7pLKzloGoY4W
IG0h53pPqFt3/2yk9mVGE15uJV7pwHk7bLu6QIvBOlWXm5lpVg8Ih+ZA7kqbaKRX
6nM0B23OA9+FFXEPnfx3vAKrJPq7sr5ptkljq2LIvpBL5jXcxO/UFpfVLUPwYN/P
OWmsu49AX7Ul9GtB3jN4r1ythuJ5A6hx78EcYsMIWVEtsdmSbFSJV/5JmNdYFmMZ
LCSKKfia4BzInBxwS6OA7rAgpyOReaAGoIgDKcd4/pvdF/Fjpfg4YbMy7zU+HAbI
4U4T9S6CU5TPcUxhRfpgx/Xmn4wj+1A5qssz/RUrV3RmLHI0VcWIgPT/m0swVDcH
1isLCF6I2qTfMi9E7uRf/9zR0GgMZQZV50y2Fzt+6k+htPrUYt7I0YrN055C0wrU
QlZpEPryqkiqE4JTH1N54/17dtIET9ksYkv8BFHdjWgU83IJzTTUxZftTtzz7lGs
xHTPVGV2om5WUwCCIBF42mRbHESgz4lzv0WCo0UKTmlFVhdeFjRNEumA//JGG8SJ
400vNZ7gkisNgTR1Q83snSeFJIcJozyS+Rvbix/WF77kicPlk+SJKqlVD0Ibg2X9
RIHhfgot2x05dNrKEtjE9w/xTqrPLELqax9rCsofwRuBv75jrOkI6x3fK9kWDkys
kpRn4OxnYM+vYzC4SXvdDPlHnhIlIcg24UDOsWIcg4RLy2/7iIzeM5XIA2W3ZCWn
/e24/ICwH1nOgKoidFBXr+jRJuKHkGREKM1SymB7ybuXKn+2fMSFaukOxvTI92eZ
jRPpjFvl5+e9g+xcAwiEl/uj7a+OoiVJ/VAoGm4GZjeopMtGWxEGLn9+BpWC8Y69
/+mhUY/vfoY0yBZg0IeYvL8TjK36LJE5DnEHk7rCFZ4h8zmKcy3p6d2z7G3Zkp8f
B6yWWEY4Qd2xAWAynz0CsweTKIVpCf6hvotZ2GM/Ef2pezGAIcJrQdvwLfgYETdO
GDaXC/ufCH1a/LvmqDEbYlAru+4UwbyiVFLSVnXgffFGBo7yt6LGCGBFsK0nnMFm
/ruDwFmE0vXP/HSWFlyCett28G4T6ZMnTO76bm43jSjvb2G/+CXECvs6sPeCqvpq
eA9eilZoOsZPxugVyFVytv04N40hBMvD661UnXIL+EzRFPv4tP2PLdu5R9HDI3i7
S7nSpoSRbEAAO+wCyhf4Ph8TySURtw9CwVn+N5O2DOkSY+r9GUXz0bAZn2Z31V2j
jUuzMnSTrfX3IFsaVSN1RXJoTCFq9AW9mw0WTp55QlNbUxbRxH1AyeD3b3SoDNpA
oEix3gI0zV9wcBNlPbGeN7UD6EnAQPpOVnTOCtm0ycbmWs5bF9EuV0QLphqe9pMQ
kFXcNgLErMvzeoE2X3wSXYqipxTydEHiUo8DiQnQaSrs3t5xstXjkR9dJoMkdrrw
AnlnNt37N6X3N1mdJ1in8rUoE6d6uzsF1ZX5XsT0SnaTuOA2z+9U6V5nczg63fly
/Q9ZLpzPbW1fqNwO1wrqSUxxDa67ngQpOlAgXDK/VjcJQ/v0svQcW+R104YKlBPR
b2emmpKyjeOkUEkwBXZo4lv7R96HFFiqsptWuTe3X2uuIJWB88S42Qb4YkeMg1Kq
fsf24PYCwk3RKw2yf9h0DQx2B/J8CCOqpjpVLhr9D+cBMbenlvjPNWflB05M5Mib
JEBUB/vbsVJJFKvjFB9JZLmZBXHN8dkNTn8TV3cw5L3vva8qTm7llDOWAT/k47+Q
VGw15MKpGZhKcMvzUc0De0ifFXqDNd5J08DSgb2ogwDF4fVAliwAKJ/anLw4P51d
LV1ClmO/I8XscKF6mfB0NHfHk8t/EF/fITceNavVbzKnSUbtQYxed0HKeiyCVxA0
APwAuNL8Ycp5DMfizsSQB3QnXqslM45jnyCj/KrqsEmBt+pYPmifl6V06inEERKf
qgbEeGGoFyWzl5C9zgfoFdJy23/hJcQzpMMkWzEFEdZ2iYG9KyaBRpJbJBDDwBD9
PJ97NnQOkHiXK/lkOEBGGokGejVY52lFsFGH9SccXgH5OZ/6e9+WmBUyUXv68VKz
P0yroMw1k78U0VxVcQLGP+SLK5fpQsgU5yt2XAgxhGaW3UQUz80Z56tnBgHFT0lw
SsKrctwgN4rr2LdV/srwZhNsAG/sMFFOUo3x7ra+1ijFUkWYDm9s/BmNnAVX4+XU
S0NZJyPEhV4YTvfN2f+Nokw5dzPGAt8t5/8cr9++wjB4d8FPEEvHP7b8NyQCjfY7
aJQ0rVy55TmiMLElHQPvCPmdht2AyIXNX+I6o1ByIjxgXrlUWWIFwgvihVy6PCQp
M6hpYw5tNeQqUdPJfXi38I0aRII4rp7PeRbfZMNxHmZQBZm2kSVRFtoLMSBfypWN
D7zx5FvsKvLhV4bVyMtTR8bsnjZJP15gPhKcNOaOEh35GjYFTakYbJyO6jZDDHU5
+Pigl/B1kOx2xk/FGBA4UnEPS5tAiNVGFJ3V8jqO34uD4RiQ6ptr+qmeSraILB8p
VRPO9g/W2+RpctZ0ZfjNdD8f7pg8SmgQEaAlkLmGTMCAGWDlA/GNBym5FOlVaHog
yYVncIhVGD2nr+wwjg/RV1VPNnmaQUjXrEY85PpgPyJFU06RT/8iOTODXQdpN7mW
/bhVeRTODKoUgGeIh4pJ1/TewAoxRCB+jyMOSI0zh9iOSPPlAIqDjB7Td+1aqQMB
FYFhR+bhNOhC/+9O43x5JjP50MOXCTrKpDIulMTWNubsmcmrJls4/4zhS0n11aOn
whl+YiXHrntMvq0tDTYawSFzf9vNTq3GHeSFCz7ohJzXkajb7rqSWW4YqN9BuYeo
dTgCIFnOzTK/dgNYhO9rvg8g0zXzoJCOcTh/W+N+Rk0z12WwQ+WHn5Mie8WEuA5v
2m/WOZV3NeoVsvuBQPhBsyqbqcwy6bbKXBQtx3mRACn7vJjAgj/G2Re9RpY7khm1
exaEuiQVR/1iO6ba9QGK0vnUEXVgdG1Qqyjq6w0JPOuLr13SEkoIb8+Msw8QghBu
C3pG2NFxiFPtciJ7XaRtYIRes9ZRycNbLKOHAX+eJxGhryAiOMJwp0dzqtrP0ga5
je0FkwfaYsjobCIpdzX3KUJwTMnSoFNLKV/Ub13w99LWHZ/X2OktzJd4iilhPRwC
A0R6MsF512gJ4qdQhnqvh/W274nsznI53//S54L91wL6RkhTagQjgpgjSFEOBdNb
7hH56WqKrPAjLYb7aNu2qQcxKPHebEbWO3sOpfquhZxRn+ARga934n5+f9D/dR7G
pddRjDc9hbX6WIRxd44Ri5s/CUc0SVFeKQ5ZgHZilSIj68gonOzS5jcIVmHR6/Yr
sQmbKOec93roi3bsis8BpZKzTWbNuDE7+7hPL6mW5JjUNxv7at5mDCjidEsLgSLS
me1CaQdsyJNizzrq/bUh8q5MEOA8dvHoXuSKp1tUZC+ETw48lyDRb/E1WdnLG2+C
PdfIN9+dDHxQdpYJXvXlp+yuISlpCdRjsbT9QhOW3pVd+ZJdRCcXtvf7KFvoQ0Qe
w0CEs1WTwgvpsoFcMTvM2UpeADRSvz8JfT/JVS/hp5lsj7hjlY6Q9NcFqMJ60mdy
c8yy19trIqb47VsKR2V7FaN/mMo4UYmhk6yAijEbpniT5SmytLFSfKJbj7DQMscE
GpReUPwJ12xNneYR7WdYy4ZXm/QV/tYTrGA6ivxvAsp48mTPT6dydNtdAd8skL2/
IFs1GEIcdEm6855SOy81y6k6cpLg3N2YODZ5etGS69gZSbNNmcNTsf8Zf0iycPg7
kijVG//3SSC3is0aamjOV7U6s6Z9ZWeu6uxLlJgr4V80vyOP1AnqtO4lvdVboCOK
SBIH/FgVD7G98TjHskeTZsoU/L9w55nSEF6x91WrNQ6N9Mt2GKFg7uKDjqlokImG
O0c3vmjHdJqNAGIlrniKaM7ITqdhjJmzfNOzFS9DN4xYxoD0XvwV4Mt1MMbmNgV3
89C1F+02siilfHunjA6c9GHrCDfL0HrhNR38T/OXCZ5LkcRvLPapKWGYOcfgRFTD
ZOXewwL7XPBBdnN+SkR9dx6H4Wfg6SyBpiKBPzTi1Gryk/i78sZUEFenbrxfD2Y8
Wuwmb01BxjNEe/wraJTZ/VmAOFVTNo0SKY7b7qhhZSazk8UJbhjhqiyGvxk2eGHV
0ki6SIiql5eEJu8egBBjJunxSL8Qv1Evnri+Dc9Lqdm1u4jx/MEuh8GHWJbVOe5W
YBjlGx+vPW9/QxxSrOOvtmWuAUPxXrTAiK0XJCfKA3048NnKbrcQZ55fVVGfvZVr
JpnX9Q3Vd3ZwQEycQ95WLIbr0HsdrZBInG06jZvGDws/oRErx3LRBK6aXCQGz/jv
BPvRd8hkEj3kMnSByoU1w4GtSsfZgibm5vY/G8/0qz6piVDDRHtjDAusaxtMYgHp
u3w5DFLXWA3vaYTR8tFasey1HSiNTBufaK9L51Hzb/+VzSm5IWvo6FYfxTeLxLYr
G2xQk4k9QrqT2q7hkqwiDtkK+66WrvWzRcScjrtqwsiuHwliw6GToLaEnmM2GIlr
CiwTSB9AM3hXtL8tAyhvjVZUi7vn2p36OGYn/uzEeIuWYpHx7pSsVPzYYoRNg0rH
GvxGbwZyxUyFAW5nbwVzzfRS9j0Sls0mi9/yM5c0MAh5H5Ty75z+CWKaON/amJsa
NeuXWttPsXjAYZFMlxgBwx/yF8r0wYVm6glK14lzOeGjYe/It4G64UJET+LGhpGI
k3KzEdGJMWRrcfwWKeitkUZB7L+9fhKa0pbwF/frw262yzOyH3XKuTKiCsUsUvb5
Z/KTF6jGgeKpM2sBBukIKU1wVn3Plc6C74xhT71AIHYY/wGrH4c2QmyJvet8X6r+
LruQwf4x12f4dPN947OIJ3UrobDo5OZaxf3MHdP9TG2SVD6Cnfei/nyj8ia5Gx+k
EpM+WOKocg3xefIGEMjFT/AZ0srI1+N8+NUHPhBVCBYTY8NuxVSsY41IiFFour4A
DQF4Cp3zNn0fMpDA89wupPpiaR4kAjTtLluQH6b9FeKfMHL6p0n8aEix3prB8mM2
217TSqduXXB74gKkeXMFnfr+fUJIjUEE7PoJta9Aze9fbtKgN/Nfa7pwo+ocmZf0
ii6fYA9tuDa5TaiVGrDOlI4aoPOepAfeAOobCPRfTzYbHocoIayNQnkJhKKjjSzP
Yt8tDkpbHUaHaL8Hpj57q5Y+r/7TAVtir7Em4jjoAxqL/nc3f/0/4aMzigXATJJS
Tlcn0gVxEqzSKfGGKBQ7ks7GBYTXQwds0XtFYgEwuuU5F/G8HZ0GzDDlxwxVOaOx
OoR8Krq3I6PQrSstQkMQE5S5Y5JlZbLLlKcar8ARBksH5acR3DgGv0R4CQWgzgsP
NgvRoT3t+vHq+yegFBAGegXDb75MqiCALX4qBWqhXo61vflp+rXXXOU4kDh1kkUw
WaF4yf3RIC2rq0TSpaeZPcKii3egCexr0ntLV+fNsqCmW21HcJyb+WTtVO8E7Sbk
tolueDL8Uo4/U5bYgMWFAK80/ZIOA1OqXN7WeCo9sytDKQG4fBpiJYDR1CdX0xqo
Vg+bTq7aq2iSk3oalS31pUNGZSW3cCjqoVzkVFDGbwUnfMWqHTlHqXFc6VwKTrEE
aPlbH7Mry4E6k5J4Fmjrw8pz7RWTS31Ipg0SmZV7kv7/ifURADsi9b5TS7Sc9tTX
ZtYDq6ExJaWMyoFXx2hJsOV/Hwemv1maXQhOu3lwyBg8gXyw95heemM6jocVjouT
XotOeAsosdaa706gnRIxKf2Yn3l7Wq74eb+X16iLyDLOZ/a4l7iMjasIyPAM6cTB
W/bcG5wvdMUx0wBD/VANKeXZW+hSVzxSH/jRsGcXqnF3zUgnUK7aWVmOma1IDzWp
n2PwJarL0YDKdYaRx/CRi5Y35ORmIJxApACsbErJ28SaM+hYlTMqV7Bk8fo3PQz2
oXgkktxBxcFThR1dsgv0Ji6zx6vthXLfROu03a8FsoMMwR5oVZRSW7FevnNmiJOt
pCvyzcitH2EZgGWj5aqxDdL8shXdJonPtDmscyOuqv3Mgl7kYvfMkoSG/gXNNwPH
nIrfqW5x+hRv1FsibNHc5VKxVWzF9EZYp99VC4W8IUJNjoEFSwgtvUmVbe6aqw4L
kng1PFK+fU7yqGK/shHFLSwGmIUuksCCUsrjsWzdXrRkERFTaIUkgX8mOcdOOrLR
pgvw3D5b5rynQR+tpdk9opciej8sKZraaTG7ZPTAAhjH/YkCA9L7tDe/ekuddwqF
OGippZuT12zRMXNk6ggg5GWVwibYu+bjmsLAcuGX5/FWeE0z5HC+ylvxc31L2aEe
tQNcyJRbWolE0yUw3mfF97zit9HjlMs7J1aXAQoOWbDuZvawg9LEUI5kx2dvhoD/
eqMgeNyac9bQ4KQ/DV0COOKMcjsS/6vONwLzMHpZSCrBBc4K6mLIVHCf8kcb2aCY
D7wwImS/BkVYosMOQGoeRA6Klb8dj78P+e+OsIC1zK4gXdIGnluys5+dmXW/z52c
4EJG7gAWJdTr0eqEsijgsxBuo7lL0KS52uQylgcrzEonxI6qN2a6jZK+HR6/Z4l9
J6bII58mJOBOaPbVw3lzZq7VKch67C4SEIBKVzo/2hNA2a6uJtHNq4zO+tp5uR25
kXEHRVui56kF1cQDGoDG552XTGg1/PWJaxfqRBo3wzmJL7wa19aCwMT2KCSoDTQx
ISxiIWMlv3WCFiV5Of92xftxl/wDIb5Aqf5pXWV3XGG493+/g1Lm55FnEw/3cPdp
f+Sg5kC3p444k2ViIzR7qgY9GdBAjws87lchL2sQVtwk1vIUTY0cEplyJIjZo5VK
K3jys7b2Z+hR3BGJYeyBTnn4FMB+nJQb3wtMhIz/WOFLEQ/rKQdO4hNB0aXplzs2
wl6BYaoTidIkwMuIf1wcTwLB/oXhWnjixhb9us5Q4rYE+9nY70wXxtNySIWroEWM
H6ug2hUgStr0LTXZD9ptms+GGurS//GqQBRFiCzCxeycFdQZNIvtWFAUA3CRgsQD
No2aL6nIsILXOZx9ZntExGqor5bYzSiJCZdQ2HEiHf4bRaAuY2CFjYkcUWQFpIO7
ytMr5q7olizmfQc1YC0XQTb/wEaL3u6SJpn84ERj92008JYESYICt79QI1HzgTE5
yXv2b1vBeGYmPYQZ09VuavhCpX8OMHmgj1lHmySgnKGC+31spe0JKsZPOcFDPSMu
25WOXStLQD9GKMwNzwDlypqDm/K9HAU+ukcjToQA93jiSwN2+YZMB7zQzwu02fLS
mIWuQ3rR6cV8cYbHu+xOrp1oOuyAsdc1IdR2TOrJLroQOHVDWJEscZ5suGIaysXX
FUim//56O8E25p05gWcC7S6EYEZ8qhwMSXYRL+yorpqPhiHiy+QPcB7zXXkmNfVH
mTzW33/zIkiLnwlPovawZoQcWRGXDMkvooHHm0k9C/uC6JHfamNQPafN9Ju2zAkh
i4FOrMX6Bb2BdU4ZjsuqPLshPojYK67EkUiqf8SBzJPcBE3K9SVre0mhuM/3nm1N
gNoP+CJVF7cmSjb3iu7XSZbu/NjqHKvBTWQvu0hT3e/J8gPt3MNPuihMn9JgP/RX
Qhg8t4vmyL3nOOVwGGu86BQU9nQaMSGSZQPwV+RVjsPSiBS+OCScsxQHXvyE8FHy
9qCGH95kQBT7dXfB5STvoYGU4DdLOa8lfONRdjOHF3fWJCrTmweZqrij+22kE4Zh
I4+es4/TQ4ORcYp/fqKK1dj7Y6ZhWqGvMu23Eg7dwxX+/ykGOt/PxwxVd8V1eULe
KieW3kcA8/qHxQbxSwbrr9iZipM5Up/CV81TYbYyqbOSU8vJL6Bdpw0t1Bdf/p3F
AX+ob4svOG+0l3hUQ0zK4RoU/hdzUJi9ohtf6dpFz4bXRaT3JhHeWee3z4b0uq7O
g8yztzbsChGGkZ03ZNrIRdlbJNXa/1CXM3eLP8Jg7KBWJZA63mkil4zoeU0fCfKl
uQEA48aFIuoCt5AtAOB9zFtB0E7MKojTZ3NgAlHkfWRgBtBUXGnmnCIQQc1rsB9U
ptCzrz+E6lziYU9EWFqToh5T9P9xZQF3dX7alOB9lw8OSxgtzhMDOXvtT0HYTfk/
/pM5brJOJSLtYy7keSjhedZVBDRJdgOE6AYNOkGt6txC0SPwePITUskWh1km77yW
z7Mt8tB0maKCjLYtch7eW1Z1MTHXeO1cgGprKQuPBTN4dbdrXUaY+D1hhbDcbJbZ
VOp8Aj+0yVo6ujnmsakjVKjmTcCcd2b8mW+jtfkjAQwpghZcQJoCq7Cm16dxmz4M
o74CI2z0omopEAtNosPqgNMCGs1AL9KYKgnYOpjF3cYua3UjdSVKSgcqmq7kbZSl
ntQ9nROg3aE+BjyUIp4fYwxBxxNywyUf7bhJ2EryQ/WQ2gNAR+3Re9FM4S6cZN5C
LS8aMAsR38qa0B8ePMOOuo0ktA6h96+3BD1yFL4ld4Jz9BY5wH5JeGPnTTiYokUy
Zeap1JJTEd88jQj0d6iO/P6lQTxgW9jrDp1z+1W0iLE4CnPKKnP2kXUZYvMmjrl2
Z/xIPvT3cwxWvLE2SjrQ3cnhvJAiHoQmp1HqYPs15uYbU6tgvO0xpC5PETR7YZsn
EmIKJnMXhGNcFwL86sxgwzjnRImkaGgtfqdtO7VKAwAOFb95Llsh8aOiXJKpUIgt
HG1HfyMj5xNRjNamHAxy8lvNKTXxskHkj1ReRb8XkGSWVoA8lQWA9WaQJkG7Qb0a
h6oWt7lodOuuTDSSOagZKoygFa5FU8AJSIvoVTTHK/TAU11AImHdu1IzsOESCjb8
t/6JX6FEDEBLfifWwZ/7133zd/R6tRrl/IFqddtbsWdYGhiUwWR0jrjT2oxaAhKA
t8X1XB95KqkwIgytVvcSK4N2fvL4uBjvOxBzWc9pVOf6wBzngUdIh4C7qX+ivnJ1
SHuVExWFut7PqX2G3/QlrcOAuHWj1tWQ/TOrAAPB56VGC3MiwsDIp0JTS9wPCulC
0Gg7k9NihlmPc3RkGoz2PH9aVFvAANVqRmqOFr2eEmOJj9SlLUndE7oxeAcxVQWk
i4EODK0R4IgAO2Pa/VddSBGvghZVFKtm/GCs9lgscWqrXmSntaw8ZGcqNrxwwP7g
cAZOie0GTGDCVy2iYgSiUZEqAH1s5ptBbFu5cZjGmxQ/hQMqBybPAGAij6/4vy+7
6+t7/CIuFo6bF5G4EoAujWBdGMOoU/WAj9mE6p0X4GQ+xzo6fFI7UZH3xN9utk47
lyAApuKK8Kl4qFxes22nryhqcX0+2SS/P0Mt5ZaaKXezJ6MhH0brK6Y6e4xPN6lH
GiBExEUimg3WCftc1KPWSSbdBivfOF7I+NJsJ2VOI022vlWE8s2NsxYIWioEGzFq
SCPPT8n1IeAmIufcVHVTsGXAG39lnwjyzzvfy8IQLxlYsbIH2cB4oAZcIyMn+Eaa
+ksF9/ZSZ8/eF1fnS+tRgqWz4VwV42dRalO/Il3ht5rNt66OGd0xugl312k2cvkC
QmQoOu403s+lIBsVq+WhErmtnGjmnZxhgghCgbp5/dx/ZpigBqL9mKUCSR7isPbe
J0bOEICYvExxAX5RSLJOGS82GMNBLqlHKXf1VJ5+vVjyydwohnLDnk+SMqmKTmhC
CcpxfR7YwkBw1wWd8lwOX2F+v9CtL5so/Y7AIijGkirirTupysN3BII9dMFi3A4U
kxqtilY84SiLL9VCtOVEpvJ7zbytBerJp5hoE4UbO+wCsS/6nl5/LyMIN56dCNWj
9oHNYT/dxpk34vOEb/mysfhk943fZ44bIFqdySDbYE4e+hY2w63H4cXkS+iQoJFi
skIN9GmQlMTalv7SWvpwdYk/5JxfQiCE2o+1ddcdShMvKIMDgm3daA3m0Q0zJxwS
/ssKrQfP6c9xtIVjS8b2FUhyFiIdhMkvknmRsSiKh0PGzXms7Zj8R+5FVkDk7sZ+
07ptZBjG/BcDJuaOVmesjYwxZYFXN3T6oSJ1kxswCsrmuCy+lLOPnJREQZWev9GF
bOlRHvop8gplmtUc8djCe5c8ZVnbi+edAd9tRYwZ2407SLrqGniixm9pDQ7GXRQL
0njr00wRoT2yu46n4qoepIv1xJ56CujqjHVMeFk/711vzqkKmIsZ3lYr/5TqnZww
tAV/qkqEhP9o+baBxgJS5V/ftxkv4enVWCioNJUfPniSEnBz3XTpSd3QBh1jhK2K
gH+kUnl6kaWhsI+2jSZzHlhwVPyyIs9LMoD3ls9WWefCv5pBWVCLZmvYFKFhDl0Y
F+9KLBsiMbL0Ii+wlJHUWcuZ4k4+FgdwE2oQ2r5yIU+GjZc+VV5UJUM3OpSEZeqO
KpLTYqPUNypivErH6vEGLxfDBeup9yo3MzUxsk8NO2tSupaP1pe367xIdEAGyU6h
SNr662WgpDOX/Y4HH3LRK/z2uWcCyCxIKnWgXvPi83jLy4wB49QIolPwVseEAl2o
iUOLAe/YFSILWWWld1ScXAN8ktX04NK2524RI1/2g0aL39IstVwccaEu8u0BpqDv
P41EStAX5AuldQj3+nFAZ0DK0L5gFcOQJhf5JIbTmfKoy1AOMnNqYUzxPQahrReh
UiptD1E2PUB400vJ4q5AmuNPKchlq0HNae3dVq20fqjNTwutgmak0gMMfKtN+ZY9
Xc0JxGoaCu+D6wfI3E9WWcMdaAFsBBxIQOlDcQekik16VAl5kLEuhCYTMgBE7LnN
JfxdYaDw0p2mCQCNCTieQlB+waIpV54rmYiLsqnj8NFxzxFvq+F6Ez45lhNk/bk1
81JdZ4WBrKFGNbh1J2lXSs7vU4wczx+QwwNlhzgjbi99b5yEhbLLIueWtU6DYh2O
ZgCgmHsXpXrPvKD5hCDdNcFxUmYUmj2s6BGMmB0xxVxer8C0xEYPNuXH3qHwhayv
vqX6eXuBJFC2lzMD/TfSNBLpdDY2PJBQvO6hbOcePJYPCkxm8uhg3tgP6QtovYRD
ZOKS0ihXOelGV8n52x2E7ZfzLEUsj0NJjRtvHFU9pO0bXy9zRsoP/9Lgksjt2sGu
gO3H69yUUOFjNdLKtiPDDTsBjV9akPBT4i54Jqzt0NyM3QKVp3SmYVInRuSZIduf
+EOR7boitzPGO3FYMoL19ZFIZI0eDzvAUMX6bUMlVkUuDGSsS0vVJ2FZGVQAC8yp
uIC1eudon7cuotDmQ+7F/9fUSeUoPkUpy+hH5zDO5uOjYaLZSJZHIB4GTXhxgHNU
ahFDWilBqYkXt1KoYGeRabFeVenZpJJM0GymJ9EI0zHO1Zwrs6jII+GoiXQ78iHW
/i0jnJsIZLrIoHqxAj9kLRGO0YAZMW3uJya6eG7ZQxhLYuw3rQXiui6AMB8OlwCW
pfJneBd2/Bg3/1GWk4urBeO3f1J23ci4qvNE3X4qYlTOJ1zHAN1Ivkzwz0Je81C3
NxrL2XjzQITfxvl4H4GEZTpQofuuxYTV56xmIr9Qq4LGIqztk4bB8j8KufXm2+VS
Njt9eRoo3q4Js5jgnKOsDyKelrotLutKfGtPT/13Egs2+SxVQ/lnLTG33JRe1WwG
HPnP94Cyzq5mhKTU/F4FuGsS26eWaL8A9LEg7FegsPqSLwAJTy90S7hRU+0+MHpa
53VePizpji0r7tmA5APO74YW06mnNhuEEzis7gBl24meS5vn5uEGDSkEZey37u4U
PS4HBZPmxXUTEUYfgyQDiwTYv1Pc3iBRryoVDo3hhGNMVAr0jR2By0ZuHO1azpsY
p0Yl3dfbmxEiqyDaaDMsq5r2U2T5AknoIASzQTh8LFK0tBZviTcu/SsaICZeir/B
6LTjZdfjIzHXW8/LaNf/QOmRVxIcS3zMN/JDlB0BDYJD6BJxYat86WSK4N+HfkuL
a8wbZo1XpPkcsCrMWIuEkil3tGLpzPrw3vri01rM+EkHAMldrAfvto2kVvtLYcvN
ZbmzSs/JMEKlNBhArcKW8PHCUmpTbkhR5b54gNzQOIjeee/XyKqDJn9EkicZ2IHK
FLVMr4n/4k4DgFxdaI+33xc4YdP5fSSuzzR6fO8tpLIy4O2LAjYNjUajIANbhLb4
/s1LI/F06U9vTMZOB4r0eV4TTp++e0fz9K7AeGFvJLAiWi4RP3ZNqjsiQ3gAgSaV
6AQy5eEYoVeUF7QoKyii3EzUgHl/yoP1o5dp0/yyAs0LYKJtYbd3kuwhK8SI3+Em
f6O8eFp4p3PZVfAzKRFgBoe7k5GZuM7g6JPjXHrqSA+FUTY8vcvQ/k8rZpIl6iNL
dggqxAtkCvLT4C7CG2FaHMiCLzOMhJt+ZmHVFYQRb7gGR8f/ML60OdrCs/C2/GRo
iasNxV44hg+Ha1RDwHdAW/kwJdUg1F0x0NdhmwRZLoMNPZsyMa2pJ4DM3LR29LHl
XJB5VDpdazWUfSj6f7xlpGay6poUHzE0Q1c5KPpPcdF8l558WZ3YuX0fGix8xlsn
pByD5Gh6+ko82XGyVi3R3r3Za0Dxe3VLDXOj+yLfUVXYV2bvKnFPrWiifuWMXGzw
8JSFmk2svoyKodIUQLe52xr2+TgAGMROQMyKc1ygnnJcP7coMBoXzZmWp6XaWMyk
/PD65Di276HzCndG56HzZ6XZdPJcQMzgeU3cGIQA6h1n1qkI9CUwwVKJ0cUtaXi2
tbsliOuA3eQeHpfyQVVoR3ITCpicOyVTiQ7ALavOyI/azSffPk4iSHBA07urf1pw
1KzSjsy5XlxZhpjM2bOmoeIyy5RkV4ssj5tmw4ekgD58hXA2Xo0ihv4PRTXGUwjd
MW6gKQM7xUU9g8PJQrxDVzTuQ1xWMaq+Yy+ADY8lUxLhiT8k9WCSnVfSXpEQ0gTb
DwsPs5zlsljnsxIkvgY3HH9rzWtRxklsqoJCXxKtWAfdBX3tju3WfpPJUv1hHNPf
VDIfdjlr1uheZyYeL5GXpNz85JK4dmPGpU1dhyHGMsdkD0gwGqjzLfOYVnunyDCJ
KWa+I81xvfk9vzAfuBvszU9kZy0NXNJg6V2qv/NxbpVWDyd3JqqvcUJdMHwlVN38
PbBjOFiHFQRopw0Y0SYf1JenLVzz7zUxO5tXLXfvrZCUt+CWNAQEvEFEHSU+SU/W
FGsQolFVSDral518MeGGOJhQA01XB/RA3Mdco34EaltorTh/d4qQC5j2Y9fX046r
m3XNr4ODBTpPsEcIhzjwkO16VnLi36ZaeUOAdt3ZWXqC5bN+49HjNBgGHomk3G9G
AmZqROGBjMsJrj6IqJkVq9FhhJR0TTkrseDBv/yJcZitRKozy1fBB/GSfFHMzSL/
M0n+3GH2RhIdxd8+YdDDchb0dPxsfwwjmT9cmrOSQdP420p9OiFGZO0PEfXj8ptp
rTCCt/+o09yso1juPlnqvB3aOGM6s9OP7jKGZI+L3d+/tHlEcCcSDapUync6J/Vg
L/hYxg1fHCApHRD6BKZYwicziTVNyb8ztCyYrgQ0gSqCNDInDCsM59y3KWFQ6CVL
H2BK0hTsDewD9jXqWzqSxnUP1MQsgT42kQXAKyxgY7whDRqR8JxXhSPMrXxHxVTx
937ovndTYz++2ym9OVdrzKUThyhOecztYQVstDpiCnrziDkbHI8KRo+qfBoVtq30
8F5G+GNBJt+a8a+8lIsKRqCGxfIaM2mdpuH52HgSjSREMV6tYH9K56pYLUW3Qwzd
gyrREyVj50D4+olXpfMaZ4Sqf/R8NBdvXhxGCHPFYu6LxDQ7+GrOpra4in8vAuKI
+6yYxpO9XM0ytfiHMOOpPaWQo1bO/swmoIucwpcMqRhnbu2Ck1P/DMAadWmcI8nD
14spbGh8NMhuC0LXXBgxsJRjp/Q4RZWvaFLHteV6tERXLOslBqaUdmvBq1Nq2XHH
X9+Sii7sBCdPpC5HkaIpzMhsqWtXnq1RPheWYk06LHm89BMlvc3kGwRHwvm1VMni
P9XZGOGNOjS8TFPzVEoTnnC/Q2Vv+Ox14kgdgl9taTFR8Ulc7f0DiTEr0CPLWTvN
1jZBklHA9z+77BBnUVOD1jmi+lRDgL0OAgP9lWlBUD1XLP0csmgpAPZiDJF0gxnc
lxpm/YQFtCb+4xOgmD4dbCrrJMTcl6lze27knVuc/Jx92gb2sfGHjhhupYsWu0FU
ln6Jk/5bXmIr5TmcmfuTXvPhB75UmAfjFnNKI6OA1pYN3qaUMAKI3EAj9abtFmys
IQGmxEUDs6Q+lXjNTpc3FoOU/JJQxdPFSHkeRk6u3OGe3/wFoNLggygHXiYe5Bfh
liVYWQoNUgD38RchKN7tObJEBeEOJh9wRauOfY/vmqu8wZUCWpyRdXfVfvh7FWJw
HbZzRAGleGOIyepzf60DzZpxrOe7YrumSF+PCr4bfT72W5xQMKotIvaGClNkzxTA
6SmPT14Mpp87YbH7eampZCRxWNhkCyFuoAsw4lhFFlGSvVbZtxqUndwGh3uxuqYn
7yzRCxGH0ptKsoUxhRPdKKBrfyuJo+JlbugzaXKFTIghhkPvF6jjVvVQq0eUk74s
k+yUWmxGqvl9+HHdUbelbenTMDcrLgQPF2N92kBgbj5FVqSOaMAKe+D22kd/BeVh
2171ZWpB38o+ODS14opLjyjoBxLF8ws9wlYfdHgUwBgjmfKL4tByCneQBFq7V1jk
eQskGtzLhMA8xxQfO2fr2nzft3HDI+htFGjLWdFD7QHS1Dre9FjdRhxaEOcHGe+u
Zn3mjQoql7oh27RCHbgG/rWOzOAQoJ5ol1kKgKdwNbX4GJXy+pRFO58vp2SYXP8u
A1SM+pZ8RfzifIhjdamJJutugEZfWiACgf/UGinXwMNIgTOJIWB0cyhSDXw7odvP
x+1iQGn2y8MLM13LdGMTxk0vpcTMLmvhXT0xpnK617gE/ueHJb6uyIFZk5xqw/Dr
yubghb1YZJsI/W5wC6oN+CvjF9yiS0rRz9wx89GWsZ2jMrJ7rDbV7VtnpyLaw1sV
zfPIIZiWWS0zGhrzPZ4DyT57/C/6hbSBBOt/fJEmRdWBxbwufOKPXa8eTrv7JK5c
PbfOkBwRopEHu+1ih/Gs05kbeqOjWPrUf7N+Sp9mWTPr3rMlvXvm2w7gLacSSubQ
LMK5/IYXHxPDE618ARnySk4hxwD/5kzNE+T0BUYpGMtaHYsaktsJKamiuxJ4ePtt
pKDbAu/QUwWLoxABAVrWtG2+XtEfalI0FUS9jVnIKE39Dwho9JKgNFVH/jo17n96
FrX2kKAF9ZX+3uqPvtrSH/96hiuCui55KONUaHw7P5uDsnFdKXKzAj++leu2W0az
kwtCquu75yGYn/FiWZkHAs12RaR6s2otUGKlN5yyhtmZus7E9gFeeYp8IcHSYNvN
vFaJfOCvM65ps9wMp0Sfqe8Wd1tKubzXJrqqqsJGnPiGBf5XlAStF0A+8YYbT0Df
rQMb5Voqt8zYGjzSMxxDVAa3pxaRK4C6bihIDotFMQu1n18li4IWaTDz/jcfWO4r
/mQfhDItCrjAnV9Q6fZ3Bf7tzsEPeyToMy0qB9N/AkUOm5yJWWxUnkDQoMKe1YtD
0BCkfjmnmugBuJ4rS1us1gQ+f/vU18cVV8uKsNOPcFjLdTlxXCEgfCATTGKQtMHF
KqS9tarn7IisolCTmuoaEzD+T1HEAN7rt+A155VmSPLQb/FF07cN0ClpGSme4yMS
ZsTDCxaZt3ItujLVcpqf7xTcoDMgzK9IxsmkH08soe1HYBQgkB/T1hEeqKdUh/u3
emkV51k5GuXItbfgQ6oG0jbOEiz+tXQfH8AWwg5Oq0ghQDx659Z31uAjCiUUiipZ
zweXuSLB/nQgt3OLC0L+cer973nfo1kOvUyT2e6L+4zucAxs3k1TFfFCNtpD2Nvb
Hx33myiB1kKWz3qtNfl5xCWL2iC7Q86BaS0xpBGPdnw8ZVwlSyjK5ABNTGCDj13Q
qEGNLHf9C53oST1iEemzwUxZY7cpo215dog+CvctF9G24vR5mmDToLSJKTh544/R
iRcIKflujPQrhCRwpx+H8vXVJf/8OkbRxF0DshNrAiHGl/FwMbAqMLZpouUWUEHU
B+YDfOoUfduGS4Bf9CYQYc/2QQNUMqfRZacuHCw/t/TXnSKKQR+PnYgqv4wEZCAL
E3d+dX11xpy1CIc0EQHBwOdzI49pylqrIzSwMkgzxMlqVQSY5aFXCqu05dVvh32+
TRtImn1xPL/CFqX8RrucrlXvM1R1G1vNKBM4HKDCmyJsrFNBmKgALBhYxgKlpmgh
xsZi3eUryFZy2xsyoabVOLOAozJH4dJlqP7aXBHRm+zr/nAJ4hUfJHlgn3v2LFwx
GtIxrYYr1NTeV/mysqdiXbIq5iRUWFB69Abfsit7XqEhkcVMrIe4fd/oFSE6Pmaz
SH9cpWqUK3vB2o7dQnMnBSrT7tQA/j7gZgUYsdcxpSqFWDOdBEj5SLkaCKd2esRV
UyFAo2pzSXYarwOiWRAG4/nxK5QXPIWlE6+mni8i3LB/2ACbpiYm8Qbzz4y1kCBT
/a34/X6QTjjbVdUGTU9nLIh1Li/M5BFIpBiudCtGfrhfh7c45BauUSsHKCqOb+H2
ZugzgTGP5STJ/DjetE4wJIq4nruFDVVxqGo8Kh4ocmliQnEjxtJjx+Akwb8Bg6N/
kAaAHdqx41SYzNtH+Fs+P+DLt5pEUVHnUaEF4/OMNqDpstSXkBCOs49ZRyZIK4Dy
fnLBmN0gD8J1hUKRyFxpm4X9iB/EmRDcoI4CUrXG7ekHLPXAdDEN6WjcJw4MiiYm
p3dqiwvPpTT/UAkVQshIqeuKJP8i2FrIGnd5Cq/SljOA76Vxms9E4DMIY1LozeVN
EJibUTY3qdIfFZQpRseYTrEfaYb9FNX/gL0ScIBFeoPdK2L6zCHGUMk5nffvVSWq
agevtQIB5RVf0fvQsf6P/wrZJoURehX8tzPovLPMg6xd0WSTm5UEKp7YRbhYHn6u
zFV8/7azCL9XZZseqMTJ8/0YDzET+iXCc7wt+P0dEF+JjfA0DaNs9StGukTi+m2n
EGGxlAAmJBqreiWZsD3dGACR4J4CuUF+jrEC27vrN1xbjia8pb8JRlNHadT5GeLP
qCo1N746hQUCPu75+pi6nZQuRTDYk5aXqbothwUZI0mdBfdIjfvyL99YA2y85SJs
FMF/uP76LmQctCGogqyr3FAkFpym9Qt+SeU5xhrYkK1uH5+vJByYukGnN8jo5u8/
abeIRU1YebbvHc5OCWfp1dn2OYEkitMCiPzVhDaNtuGsLjaWo4KKaVTLMxj9x3dX
/H4KbbiS+x1Uv6cr5QFJ0oigdbgcgbYr+Sd1IgrDAv3+Docs691465kWxL6coYK6
+o88ZZo8MzXVg6EFprJ1a3y3xsWEgv9g/SbXQNNybLb11b9oatxYNnWrp0NojtHw
3zDfus9iE645Ulj/arDdN6O9aJMv8c9VXEgGD7dZ3CTT6LI66F6SM2q4x8MwmaRq
W604yXahh7LKMRKs+yqXobcA3eE9fLpdsre47QnyoT/JOgdL/i+S0UeW4Ce4tbAO
BdFML27Cev1Zyl4Re1xPfGGGl6JqcJdKavOeOHPwx9aukf0aW9PJIITZcTtorY6C
DYlYg5l+K82N1SPI/PL4mkLU3luu40O/yUCcqGMTCZSI7gVV3MUtsZXWSBgJBeAe
oM5vBSskj6UrUP8s4AtKralljhVnHptIZmftpRZ6OxfZS5cxT6bf0qAF/NZiMmt5
SCx25PrNbDKoplPHdvAvXNqQXSnsF+rz4NVERiLQ8uuhqyoSV7U/T/2JwyfdnK4T
zIqs7LznJScrkAXvaUShG56ARAopA2PQ28n+L48/RzBUcaqhub4fHrsB2HUW9Bg3
jNA5+oupEcegoRDy0XGUjdfRMg9r0FL/Ve6ze4ubS9HjDMDBkE59jLPRAN11VZet
OMUaSoXyaWbaSo5WGbkogrPlouLzc11v/wgO/EdDno/hppGUw5Qx8XrB+vfe3Fyk
FEENQkU6tnsnjE4n+gh0gqqIlq/BZGPhpGajdQK3pzLb1g8A6n9z4XRmqO5DwFKo
wtnRkDGlieg4gl9L5sJEKD6azW7g2sgEU2Et9NWvf9MlFSlCrmuFb6T7T259M0Kq
cA6idNUYBaB59Pst2mBOiwsOvZmUqb9X3RZ9kdbkA50PQYafmRlFyVzMDEUQoACI
H14YcrISXXOS17/qruBwEEv5k/i8FoPbsiBoLXNxBDgQiQqUQis9MZiehxZFhtAy
s4XcSGBmWlJn/51lyMz2DkIZEYI9mg4590hewO0ykw/OyqpiPSegaGRd9Wb7UxX5
yDi9Of46W+MVLQzpBjMBPYtdV1yRU4xfX52gE8PS+PAqAVDoN0dIzLAbxrKro3AD
rxw1120El0qbx0CS0pRaw2KHX7isRVisdYW53uhagO2KQHt2LeylDehtnZ4l5LgT
p+ZNwjQie8kRIQGprLP0JAFc5q+RsmqqDR6C3Es7YGu7oPJhqRMctYEU0CopQ0GI
ZZveNnVrU8sLb2V+WGX7VHDEwf2c6z41uTr9aQjQrtkEUDzrg6OUxnGnyFQwon+O
tWpCr4hQs1DnxEcH6KD9GjqpML9M0SxfEgiwTqTWTu+Cu7x6r5AL2BR9OgNMyxOr
shV9jJVzwVXnxLvni524E+Es9XG8ZFEHjtPMvJlZLGb755s4KR3e2SgP7iAdxYyt
4OAJvMzihuXMPRCYdvWUXKN3mp+RSsrhOX1mharQykokwHdusTQ12sN6fzbChUUd
cmHf+Q5xQ276jhIJtSy7gKh7pN9FKi9YMw2jHtLrQDDPfVPK2YaNPoRBnlrbbMrp
FOTNvJadD02z4BXu27SB8rk8E6Owdve4XF0TzgSxzrmzrcCsGpiJNQbflBwDx3XP
CG8oYgJeS9zM7D0+GYk3rnK4nkmnHveROHQhkoIWi6ATpEnFrPbFrp3tSO1rL/hx
e75xTG8Z0MlPgGDoS+i1Xq48RyQi88HX14T279/sGwBXRogt+DISBokXaLKI338C
57ONZ4sTYHvQGVn/bEZCCrHcr+6UGpsPWGhdmeG+pzDDMArG5dI56WXeJy4ckz/l
SiqPcflUhWcr6d4dMRmQjlEuRy1M5n+tQuXqN+uHo+7RPIzhNgInmzxQ3DPRpLnt
ZHbDefolhQX0h5Oyx6y0GKjc+0SeNglxphnEaWYM5ZRtcKnkWVwH211Uw379Dzv1
DndeIQjVYz7IZd7gstk0qmjWIbH0vuFZ/lyt6oD5MZS+QQcJS4j3vuNRLY6Hfz6l
qt9eWfGb3CbRuQe5Ow/Bne3x//dS5wEZbEJ952mKJTBzTUZ8T6uWFRukb3Mdn2qB
l0+rWqIssBDFskAKB9OyvBanUayqsVsHEHIPgze5Kyn1pEsFSZlpLgAyYlmnmB8z
ixXk3KQn40bHd9TPWazFaU4xqAGKjfI+ZiYygHrlKjY10MB6boMZ7bbKHrMRdMD1
4EODzhlktnd7K2+wpHbwAGIdpZjZTZIk+0sN9Z2h7u9CXo3htwE2K3OWSwswmRjc
E+W5Obd8xP6hMuiVj1iiSnLSnDZ6e2xaX1B4DH/feKuK3BDLR97r9/ui44DIDjsL
eBbgddxQr6LEQISjXuHWW3kyu/z3VbVYYVSHqtTD3WHy/li7SpWKoptDZl2LCrut
LVlnmI4ppRosqCrwxdS4zYdVA4qFxZR8PlzDd3MdNNqiXEjxejdcezBwIppRA8b5
NFWgQovq0KB4nsCFN1bxobsAfVyc+RI95XeVynSy6IFfzmQgsNTVrfukurq6crAs
qobQWC1fFn1QQ1AfbHn+lVqEI5jaApA1I+0oL9wr7goYLJuCuxb69cHHvTziWvgK
6GeIKZaW7ZtZZtaBk/DzD6asSXnFKKFxTIsb/VVB5i/OnWt9gHm9qugLk86Rc3A0
AezHrzmidLxyo/hQgBm57MWT8x/RAQ+/q4F8Ly680+ZSgXxIShdJ+S1QpagMCgO2
9mNPkV2F65nUko/OBCIumTD/fkhwwupswnYB/OxVbJEMm0xnMUYhMnKMbMOCHHmC
cjA/DnQ3R9SrBTKv5GpshHfzDcR0JAXiT8wFsrcxE3jHX+b4EAgJEzkI12d8FZl1
mlGdHwNnj2NgFSCdaX34s7n/+h29mI/NA7arJCsHdnZn0XIhLz/wArg9iFBuLfJY
L+NvAQ/d8xGVH+GCszavFAWljfdr+vqnDk15eDIK6dM4/QxwQQe2/C0HK58Ts6jN
IbepG1tDvwTkf2Z4yMz4ypphIeLHs7P3vpVgQJcRDLDqWpfa8TxGUtNOwpqXeLiQ
9/DuuFHgg9bJC2Qtse12e2lmZ4KesAYemnu8jmfAgn3h6ZE4q2Pg8kphpMLZdxLz
qBW354Z+IQkL21fhlRXnqwQr6nzCJ70iOSwNjZJf+pVRIpn3+aPxeVfxXuJPjf5G
C/9j4REesdaklXd4vo7NCrKQ48+ncPEFCHbC06SawcHafKC9nkBOTDp8+vaViw6+
QPxq44A6PfF0p7G+OccpNRmy7kWiTdfE25ietSXeJIfsxRNv1ZNKgeLiD+v6eNZq
y1hOt2zht4sXV7klX/MAzbgckv8LdfMKfRuro1U2R7U03eKSJPmd4YqadPIVIwvA
5z3rwxagibuZIjdOmDyCKlotUvoF2MHi6Tgv8cBIxT5JRL3OoNj5/9MfGgKpnLk4
rDinW4UhQqfbRNpXuk7boeig2Y01e3aku9cSvXRqX8AZpCw8Z1vrSokJFztGfF/D
R/QQImDjVxmdkpLP7tyUCfioqJSjXpsyMElwTcs5PiuhuP99Cu7jHOdKa+H2Icv5
oEMW6WVgGfHO6ruFZfy5Cfag5xa11feyonJ5gc87ochLin9nFwcsg5EGVIyJIEs/
BIM9eU3nVeYB55KJSres17VPMC7ScnWLQav/hO736AO55MuDRmJAcvqSWk7pQdDP
xCPgi5y6Ley3jfG70gO0uYSYJE4b5XmxYUA1EFpw1kRbqdj5m6Y8oZ9Tn/SaW6DL
H1knwM3SK45qitsPQaf6yn0y2ujyxU7KxzXel77vk37Usl5MAgDsky242qtIhGzC
XGvFS4dcAiXK4rdDJHOB0ADX2ZnZ0Z2XUoYQ2de4ZindZt9iq/GJ7lJy6oaXN4fs
nGoyFTUxTIxEPLS0ayXLsirCytHtls0DQxy5md0jFIrvoEUpYun0Z6zJS5QDU6BB
lWeIzED5+h3dOESM/Orz3K9Q8kDr/uZtiODZLrvkEhDVd7dodSZwMSOT8iB630uz
qj8awpRXEV1tHvGml7TjWUW+hEhH9vGrTgPslBDR38/qvCnszBj2aaMHTAbNwhM6
wXJWePQQKWdseahd+Lt8N1WWbp+7Oz0To+ldG4GVDxbKbyJOVMtwCxGTTToAAK8E
86ZcX0CzpUqGhWs4WDkCr4PV4RiQVemt5UVuuHmDY5hz/Uq24BK7bgCmoZxHk/7H
/QECoLYd3C1/iDEs8sxAr6tKcmlm4aKoJYgJWEq0PLHoWpLSVj8gsxXBEylwFO3S
n9zaNESqnbWhogCZRn5fsT5jjw6k5oiyuhmqpCFl7UF1VG5q9mghgSPj53Lf8SeX
vVxI1Y22ufaHLmaoPdR8GTc4dAhpbr5J7MszTJGDmJdzm3zLcfOdmwWNCeSoEKv/
4axjQUPTCfmkXMg8IUbjROhPxAtLJcdUZ+FmDH/J1XbbgRZlE9m2QPWGvq+C/kqm
+SdkWUtPSpDcjdJTLcozvQdC0Mwh2IFeStmG8kq01SHu34ov6MCUlRlYWsJ6WxvC
nnqKAY4cRaMGkK684lDReHFXef3uZ7Ei45g8HsOHsg1EicTxuM5J3E0tdAU+buQ3
2Qp2HNbV3igLNoC4ediRXhcKv7UTnLRYYFFJoWzj2puO1Kk3LNbUGkzL/logGEdW
cXFkqxmREbKt7Q0gT63Q06PAZqcX3WVOvBwwvNcwil3Ksq3WjNZdEMA11h3WITSL
ythzw5lyLlHCnfCQUmfPYrWr4yavGI36fChHFr+2kUUg820xH6oaxm8plN50wepi
o12xAd9AhdPTxEqZ51Zb7Vmjw5JSZxVc532bGrLlklkA5w3a+w92Y3JYerONDnkG
kdqf1PednnaU01e4mFQKNeyhUtTEjmz8GIIzUhrI9G4BLHaju4iNhfOCiVM4wbKk
mFxWvibY7jTkIQQ7KGWTIK8pWMddlRTLagp/CRs+E+G/n/EtFAgqTozjQCW7au5p
TZI0/Zb3uZJnX5bjAjS7J+DWt+mTJ1cAEl1etsh9jJ5J1R45WQqOtWwWM00vn4TD
D/onQL1hNDCxrDb+2+DtKHZwMiT1/UzkUd5bdG0eElgN2JlNjqe98Rm7llwZwE+q
dqcXzQYYbNbRdKmHxqAuUWFzTh1ICzbEnEcoCoyWz70oviyhZTqpR/StYflHS3fF
bl8GGlsV3HxVVmjwkKAadizuG8HD9VYqffiBfk0i5yaco1fAOdnu99VKAqYUn6oh
niD7KBO+jQo5vEa0Z9zWwBTx/aYtGiUjo30JqI+/HctsokGcJyCN3EIh1i0vd6XD
993ftXa2hJL8l85cSAcFAamcl6DD+PDPQs8P5+2RWjDy49aGeeGPopw0K2XtjAT+
P8lqMH5ixlyc0JTqliv7vdf+mseLnb5k1ZEy3lMgP8/WnrOI2+C+2FP40UzW1/4+
4cxd38lYEsXZfOQ+NvLNe28yCyYNGhK8cCWfrylblh/Jt+CNHkAyvT1CTPP99RWC
P7ryHzg8t9LMd6Cfmn6A+ZO53OT+VISBSjjUybv5GvAl6CjVRbqsgtDz5APkgv1v
SQVFJZtSiar4gG93J7iM4EMJK7nCNMQWmm5IZGfHTUsMKqFpOSf6XLM8lYsXy3Ba
RXdriDlC+PfkhDi6ZK8Q9KWgz+BbkZ/h3nukeYIPjn+eVih5dk0n9jga+svDBxuZ
PgpVKfw6J6ulRday4LqU1RnXrjpFcl4eccD9eBZIdvt7z7HETOcPKlsXuCW3H2F0
vyjgeZSAaY1SlX6dxEMuhZxF0/qk36zFWRFbYhFl4iLgOl1F8dhI2RTVfwCmU87L
i3klhPWN8PsLT3XQ9YAiKJsNfX5bqsIe7soegfSOtub9Qa8UCXjvHNs0e9YU/9oE
5PpkdocEYP7+p/PRu3ym0OLmDEFOVVamWpv09ok8ljSkQsQhf9h8zwQKJnbdk2l3
efrmFJsrAW3k3J5EOafm/af2liQ65rEd+zDWzG3x44bR2zNRPeE2RnaCMZjGIY6g
47tn6FB1e9GSKgjFqtuhkI3ttKKBzepfiKcOPj7uSMuWYAX+6Nbvhl11ykBiaL9P
18c42kc10oNDN3rSesQ1lQCtTeAwJ2dwwbgjemyiqf6qKZAlFyzFUDAvVODs3mem
7tl2wJH9JWeAKEaj1+4VGjjrSJeItGaYNAIg7jIo2yXDA7vBRHAuW0YW1uxfdBdB
UtAChnLPAFkOgtbrEh3lw5QFBQSYA2y5AUmqqTPI2FX+uRRFceEV/6CdmUxBjgWZ
Rzywv5qNZSKyUf2vKR/fBAiqXnEv0mWQ3zmQK+VqPK/qCyuzhFRYVsffZ1oy74/I
Td9rSwOkk4M2USYsBxJiA34Ta/jxpZWjdKQGHkA6O0zYDQ0vj5ruHnW9w3cTUF5A
n+EkzBpNgG8DDUnxielRqVpg+1p6qYDgmLxhd/eDeigiSleDAMqrrp3DH4x9U9Tm
lGUABxX15NEgLDcVm7eAC5nIcytkkjnkThVplXwK5wz0pAiSy4c2Gt2R9cgBM3fW
d1NjrGzkoR9YyCS4bWl6tgmbYzFu+vXFDTiahHZ3cJ9aWGNSSqnQsaR1lV0B7e5f
i8972ssuDh+UKUBdTQlJni/MPUfndTYlh5B02vNN/pCezGO0WCUQTmAcFQdgzhNe
XD03I+7KTYj4TRmT47WYN4aZD6U8Q9lhIiDhKQlRXo4Rf4+DXQ0vA6dDddyByRYS
B8I5k5o/8ZTpCrNR8tYglLygpiOc4C4ADA0ffFFoB1GFM1spvRmtx8imJGgo9dln
EU8z+5nH6o+gu80/waEpWYHxwIWaKOwBKZqJ/5bnqDdCadYJ84pL9cyqgGlaIJYY
Ui7UumRBHnzA23OXm7OgnARja4EFIAIEFYt1LebRyrCzkZ2PKQezvCTYp3qdqS14
eHEuOrgzL8TfIcgDcQSiY3PCTa4KKt+oT8TOVxtIKtdIk4XFKYGdL7y5430FYJ+k
K+NT+jHPKVg1nfitBRkkqv+7/bQJAvTLLmnU6mhbG2obe/Do7pXTnHxfPXBnKh7S
LQkPHLvrRBqQ4jfrTtMTxgHDd7aRb2B7gMt0rHfMYePxtI9NxwjfbTOfIcdOk4Zf
c0PRQ6dTutwWdLR+50OJt0M+5/LyVg+3bmQZQSDL8Ak2jtTRwj+lgjI8gPpvtTi8
ruYQQOaNzf+upjzM3ckjr99Fe2a8CgsbrbnzoIp+c2SVXimBFsiwgpIa+KiG1Tb2
JwqPPW/gmHMrekgeYjDrm8RR4LokbXdbT9/Ev8YzXhwupiKAl7df0RHaYXBZmouY
BMG/t0br/IQ9DvjuxXfPAH+dxRQDxyWnBO7MeMgLeO2H3lumyJr1VA+aE8pYvK60
fBqebpgSDme1tnvMNU7uBVgYGFWRhy0tGibpfDTLq7cUO7Ll7RwoRrHXe+VpRiyz
ebtshYJtxrWR3LgM+7t9opUv7CxMoDwzO387tICL5wefeh3+DTjw8aW5a8IpDMuw
qYFhk6QDogGWDmmUg3gFrk1TmnYiZSNZSv2e3kbLeoeK5ozKs0ImYydY1UJPm1AW
m+50CW8mLI4cPJVoZHLj/pyhmVwkkXrgwfCGr18CDWflqFOuvIT4XfZhHXSec29b
aqybUk1pdmKch0e1tbygB/NcAtYasN7jemcI2DmKCewxO1k33X4sNpXYDZsiByIU
O0lPvOjRKlwgiZsmWBRLl7dtZHetFwbR45M0stGv40nk58vtaZxcKJcS8ZydvumM
kgEzA6hVc7deZ63366ERgYPpHLW/iRoGi4mRZ++Ia/gAsRrIHyH8lrvYmj0qoDr0
9Bv1GijYVvT6sTueVSCP5XzDskFQ0HtO/v8PNUMUEyi5B2IoiaWFUVwBJYr6Ip9w
bpfw6PItMavM2P5WI/XxXaB5PJL72sNyVWTq7QAEi0NMYjm6rV9BF1qh0TjjVgJV
II5CSQS+SZrRA7jM/S8XymQAQyBVngw5RdQlz7vXonaw04RmkTeuqEsB1J1LBhOv
WmLdy8MR+mRfNBzpojX458HQrpfGGcp5O5sXUq8jjLYkoIk1jGgo3bI1vYtKGHAc
c742f3M0zmzniwwxE4tKsC+15SO8q9Lstl19D4E/Kx2vNZI20qUR9UoIQCsbMfWO
jMa29IgNZFHvHoLLUkQxW7CCURcuKLF/fW/iSBuO1vxrZ7NP738nF/0zCEnB61jZ
vLrmbUzhhFioql7f7lWluLJg/XKGzhzaV2eO2nBf8MhGKakjSQ98PslyRB7JBNry
1SIGAfjx582rC3xt21o/ACFP9Eq8OF9G/I4Z3OGTdCncoB5r/l9lrtWizFcz4F4z
XhtQRl7Y2w46GnqoxWQtw9MMV7KujidosZkgs81GAXYmDzPbVZdzLxPPT5flKFZC
eI5hCku/TFqovT7a8usKNq31q5V77MFSFO09+5zlaghLtKzSxy/+3LIbaqkFQTy+
OgKlHHDn1RN+sulT1RFBskn0e/cxLaK2+CpVuKoS1eERKkEkkRiNZHr0feXjxr5l
PH9ABotcECxBW7WEYS73epR2clpm5D2VIaAgDdTGixc3Q9xn21n6eaD0Z1Hfd9iY
72L/Ne0iFpR50mGz37cqQ5IVOto0u6xQwegEc7vUdmB4frslIFd7ecetWCmeA9p0
npjWdHkyaC6IavP8Ig6ybNN//UvTlULBeEIOxB7Vgmi32d3+O+6hJeQpZdssHVwx
LqHIk8eEsPbvJHYDQnozjNehNrf45vEsanLPXVkwl7gy3fXZvuUZMZ+ByVyiVCSF
HVgn9lhYGx33hNN1qUCdWW9KYWQ9h/3/eyiYo4IlnAqf/Sj20QXlY0DoA+rBIP0u
paRabDljrL1bqcsZA8Y321sEbvQobjwiMk/tYfho+nQLhWLmw1gE3HuoArX21w1R
6+QMDRHwCDHkQTkGF0BfnSKQF0tCO3tXxrplZ2H21t2FglDUGnPpoAoomQaWn3TI
Lg1F+m00YHQKhpwZgyUen0jE6NbCWx3Il6ko7ZH63tBBO6bIGNRCAmEnjHCP4Rvn
buts/Ed2fweQrvl+hmJd7nEE3/UgaV6nCIG829T5QSb4J1n/GNg6huvtI9we+3ov
DyPjhsgRbnU630rl85KY3hn7qSYneeQRyGTaaa1katA6ig2FTkapqgXPwPnFzjVE
VAyZ6zfJ9v4+SKbcdiXMdDxm9qEe3JGPAaiSNdQEaJyIyzNSgLA7gKqXG81bl4zJ
VOvMGOZ6EtfOO0jS9Cdzil4vfY0695dqcct7La3nwCIyVY/khutAtkPDGp7x9BVh
JSJDKk8tj47zexRW5iQdoluizNr8W8h2fkAneMdJ4imMZNqw2+JXi9jThatthJDQ
u9+DWWBYIjny43lUdxAxjW05ZuK5UUnBD3z633xNK6wXr6qMpZP2h1P29emOnFQW
BKpy4PRbbzBqRM00qjc09aMUJyGVOB4Q8DZNPFn3Z3SbYx8HvLa46xPoLDZC6Khb
tRCACoqQwTOiEvAtQIFauf71xvRb/piiuigVLJNgqTlJLCuTm+5jZRAQGtjuON2j
YkfTBIZfZDdOyELDZldXdcYAjk1VZaiUCoVU54PEpwIQWj/i1qe0HrfZLVQn0jqi
1M5ylvakMJjt+NtLErbwO459jSO8EMh7C/fbMlU5cdSHDyltnv1vt62QGETNEI2f
Pnh2rO60o6hgeUkmZwvwOpPaWdF4dfyV85XoZq+BiFdr7Hae0F8ZY5P9YPr78jL/
3G3j8m4BdJFZUZv3iNDWOGcIa3UywlfqKTFoYLbdtrMirJg1m9st4eWXm9oh6qtU
Vry/zmB8xV3+odM7syBwXlk5irHIIz+6J5G3Ggl1UwlgwZL5ZE8OLr2tZijQatdx
stbF6ut3fMrJIyiQzR0jh1lf5qkGNsXw70dHIaO+LrgXv+0iEYzWWOkPpuKBGRc1
a/E0SF0m13oFzdqSfrQxJipH9mcFGitWNoBmdk0K+3hK2NlAN5vU3DmRycA6X1Jh
IcCic01WK9ie5lASnWlsx6zLHCEcY/ObPd3ywM9NINJF0T8jc87z/ZKrBfBmae1Q
VckaFCpLjhJ5DJmJEmhHKBflSDS2EtdkPiAEAVPdC5j4dbzYoHaHaOzfwalM/HY3
Zz80/1vEjwHz+/uvx2XiNCS5ucbaYrFtkoC7c0B68+/QePI1H5qvzjuAKf2rjgwZ
jAYOVyTzWOV5PJzZH1LxH8sZSN3z/Z2sVbyZO/CIZNEqsDv10Ce6jIdhJT/B33MV
/a3gL2hV8QM5sGkgON1sCA8RU8jOEXhRSvDMfOPZtxkWZRph66sFK0V66tBiiOjF
DmChzBWeruMotREQL5Gx5cfnNFx0TtE67iGeSILns5NWiTpmZ+fvy1jUCFXciFzu
Vlc/9WYK8qAeTwBnuRsOpGC4/pdG1aRZYtSZ3xJZW4I4vQ/K9IOD3pHs1jgLiUY3
wjhpK2jd8gc51ezNvBkIV3pzgD608z3oxbm/UMs0hVkptNQamtGFI8nObTSFac6k
V3AvZaoAmqcEg+SrygrId7ZJwn9rFxM49laqVGSLWwbaILhiLtUUPPpghVrC3E9X
LyvrQNvZj3vMjLFnp3a9XaBkhJiIlylZrWVDc9Sa7bvxCKozrOy97hBFMS4F1YHJ
DIoM4wAGcs8u2BjK56b7CvrifdrBH/1e5flFFtY+lbJwuKgSfvIZ2PGWOghC/u8u
No3MwpiOU+xpLX/iCwK3Imx1pe0c43Hw2Md77RkhOOjKfvm7bCQEn6zv50S7JJ1c
I5x12CmZqfnsnpzcXyFn+dx6eG3MXdfqqafhArTZ+fZ9x0UdaZh14NgB+oxY1bo1
hRfS0CMXa6E52M76kiHuaqWhYOC4WMpEA9pTQaNa8tZKC6e2+Z7LmLdqYiyVo7ez
V64xtL70AxksZhugbbios1XUiPs06Yk/8IKn9g2MnsgJJL5bOYoG3gOl0CYN3LHP
3njdnnj7tWcyKND6rqGfpUsNWwTZBqUN8HF+OgzVR1Y+j+8v1PUTdkL1ivVVSDWA
a3qLVnQkXNwl1gkLcuny6s8K66KBsngDGOCIFIw3UnEFvBye8CS+AbZxbVr9KomO
bFV7JAkdCW4veAOzHO/EIWWA2Q+x5sBMaNdhRRI2gUoLTI2w8mBx31BGovXgvXVk
YnMhgMVorsUfW/cikN8+zhLejfQCJjZGojP6m/siBy7lJ9VfRF9DHOLIsTm2e6V3
XEXVuXiWPqGrYsoq/B0ouNmrqBIJMELSC6VzxckyYhZFzh9oNuc9gpVi3Rk2IftX
4K1bjt5BQcRzWxFvdPyslh4ibtx6NL2HlQ4cjik/cJpwHuWsWXX4lXXjGXgZco5C
YVdHMuUCkwpvU4oLZCvtmNOJVqtuYbm7T2G05QMZX68X7agAdsMNOpQzRDtZfjtc
qr8r04ozQQBRxR7GB48r/5UoN+UxYKZvRhRO0rLUW4zri7CbZgUm/YjHbfXj/F1n
pkXoFpVEK084ZglOISBl8PIM3JwrTnNZhg24wCk67LN17aEfA9HuOhqH6TsaNsEo
hxqxtuCULzloulq+R1nrAHoCZ4K4tDOVtZ1+OEBehQ8f0b9voOeNbLUhpyR2ff4W
TsLinJstMi3Rmht+EKLOsm8XGfJTpCPOeBQOLRV5vlLf+DIcAxkv0aq3ZJxIqdSa
cTf1OyHTCB75sUQYpOM2zeevOW5eetnRUdMykMEx0A/kK5mHWshamSwDaNlgKFht
sfHj3KoIcHNAGsZ0RHLRrJdA8oDhM3MNtH8h0Dut4E/8RF+CmCXZ77KR2lKclDEW
8CadPfBwSxAnkH04KiN/YwLNefmtgTI9awmS1LAYwY7TdZR8xSzgB7h64IU+uDBp
fzu//lFYNw48Busg/hpLjl2BjFCLB8QmsOOJa0kiprJXFC63YF2gAYkkxsAnmWpK
YdE5dnqRBJUUgnd7Ry2g2QT5uH8xp/qh9vsnII7/54LkU4/zlnpqJKJMfVx0EZro
Dc+OUb2wMYMBVtDWwkJcOReg+ee4oHBLFjDcJnWnVVIyU8BbUcuLObWViBClmqGO
n82ot9uIsbjZtrZsJVQ3VyTfVpgJ8D+wnEYCdsK8+YhUfA0LVCDRAw07WxyziaJe
Gx0M1w0Qlivj2GrqNAgXPbx6KIyYtGAguBsp64hGcqnfwFbIqmktO0l8fTj5dlQB
UijFf1LQGfnbakiCexxlCPz84sxu4ubDsj4vQN7igfqXGA7P0ZrQngGJvbCrztZJ
Ax2lGI+OZpMhv2I031uHijrCgDl5iVfBBtdj+i872hjMnrnSOmI4Lf4/r/AxMilD
4qrhU9E5umQNyQvxwIEfXhFpIsvx2zhUCXqguBY+qfhyLI1teewO05KQWvAq+QnQ
5CAH1sscZKaGCVovHBlBRXDTVjHf8TWAJWKA1zVN0jF9RuGGJkn5lZNyJNJBNHZW
ipsj98mm6jOi6Gg5B/k3LmtGnYcbpGxFUr/eEFspAi8=
`pragma protect end_protected
