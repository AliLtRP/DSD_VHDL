// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y/t5jRh/C6iXcu41zCYmRXYVlimOJmhurIAPFCTs/Kh0btyuuhWR8gfy1mEJAZn0
xLfmRtMGrATNaJXOcto3DxrRVwp1EHehow7ZG0xF0Ht+ToJvFnMnp1GSu+plFB5X
kKH5nZWiww9bIfqD7/S5pwn6CpwNfRBQ62pxjQl17M0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22144)
lHG8AxqEWfuyp9BkSpeOsQdbzYHOOnJfeNv/uy1n1h8i6lqhtwWWeT6vY0XloCxf
KJnd1UhGUXTxxDqKutht1AH6zORvXcDdmbupcaJZIcqrntLRUir+bKwsZkhF8whc
PEF8JvCSUICsG6xgV89vd2pjjeLaDNsLKB+hnJ1aQqXHDSuKzelKK8glD3qNiaEg
Oolw3UlLMGCy4/ZihJP7JFZj4wmbyFwHHj9QGEhjKewUdC92igmSclphRflQP1WD
eb7iM6PR9sXmYgQWDpDdtAucdmYnjpO2pyZWkfqEYmOjKB+jUFOxh3si0AOz32h1
YuszRpvTqEuvar+qFFHUJOm7aiWLBHRixaBkAoVpQQoooBw7R/B5teT6yJK1pEDB
ezhhRGsUXCuhdAIvBQd1ncwk29/S6a42OSfcJ4S1EhSMveM/QSfjGUSjnMXgu7bV
NGmjO+pQlyhGdRgeQzBEopFCgxN4DtzxkIL0+vtyxuzjNG/boSrKQ2EY/O+8B9Kj
1/CIPBAUMGt1dFsP0zxNgMky3kOPLQa8+5UokTHncQsVwbJRdTnZlWKLUC/r+A2V
sxIbiV0xTbsFYE6BTDlT57yUpfGV2C8Upub46vTDdDeWM0SVUBXzlzvGnZqYIhDp
HzAB9mjKXrvgYUt0MyWWyLmPPPmxwSR1jltleBCkuheoqMCTljHnXsCsVOzvTL0H
8xM3NGdQqfeP4KnRlCT/NpBWWnW9ylGxZ2FgGl9SskhgzzABjhjJ571XXPweOhPU
c+CcElPR8a2fsFSDLXNv7OQ7LOsV52AL5YO0TJ+m2oishZlGdsygk4CAFtHh6pF7
wqa8hx+WAo39uwXnq+Hsl+zHWdQTkpBV0vztqLutytJxg/gYqok2HTDShn5QOzd/
B7karzRsK9n+o8ksQkqpAa7pYtvnVz4FBwq70bpmPWH0lXZNbY8qPUYHsvwjrDRD
6X0JEYkMGMHNP2YHKPd2LW+OywcXKcRzJo25XsFMlj7iSj8Y565VUXtfTeeFSMrV
0RBxrAhEO+n2+xgPWRUxtAnWskl1LXUEkryTMmv8TOX+y26yhP8mQOljsh1aJUSa
Y/M/BpqtQv8lfRJ7BRnke+SNQprJ7D+4ajxWJ3mahbTUClc9glzZY9fYhl+iZfZe
qlh3FneBzzlhqWqNBDXr+Suc+jz/z7P1OPkAMfFfdvhZq7FhBlE5gCl0POkaQ+I7
dN4KylsnMGW6qc5tUjiRlrvwbwktc0Ax6rq/LLF3niYAiWadJTfOrYCvLViRi8Xn
OEXrduXGQm62mK/HJHZhveHB3IsQZ5lENywhfvmonZvYwEtqg0KSB7wL9eqqan0b
qI32TZ+d59yAyPRgUU/4D0J6trw2AL4jeWHbSNMIM9Gq42GjzVf6EB9Zv1Ogncfh
CANGA53AIoZcJY67/VIJwwrcHNiXHz4iqB/Gl+Pq3v2Nwe9LDwkY6NlgDa//msJH
xEYSdz8GFItTl1GfWYbWSfE3MCi6rRlZWkfJD1yhFCvbh/ZS+jbOyKjidqr3XCZw
vQTzbZcMT2D+GHqyYONTC3igZ4PBcVRtrXDlQQtqZl4n3+qxaPKErDBLBAcD4qDD
jFs4CPkzjQ1cU5/DUlUFfv7B/yzt/JSp0ZmO2fWEKy81ynegLq1H707/QenOQEax
sdrEI+C7XbzgJgsiMR1DFDf4gvc41c9/6zx/JFRTgwpj39hq/oweSxkWdoEs0E9C
auz8eNw+x2WcihJDw2NutdUztsDOgQbOWCjT4aAILLwiWFetmDnOTiK9hdQPYkKI
PZx3q+nyBTsGqDZjMgh/wG7goQOsXJJebTFS0nylKEg6nATAnp9OOPIjdjOE1cN1
kbO/uar5mDu9prziOGzK/DZwAnxAjfY1/lmj8z0vRoW43zTyH7sNhOBXcqNhMDeJ
yV1M4rDXBmWI34OAI/I6ZomysK58Lvs/U8hUxc9Y02FtV3xbYVfCDjmXhN8WkNHE
mpOk9O5nE0aC2hl0Rtb0wEqwFeEiIO443OuRVfpWO5A5kDDAzWN6iEJcu7hTz09T
qLRkZ2VOV3zJcmkRaez8dYq4IHd1kFgjaEl9p1U1scr477/ljmBtr+CWZOgSuirV
2Uj1M/bWhVeDCso1bh1/C1Z75mDTiufEuIdyx2YkU3ZW4ClVTjES8M3iv6gwgbJc
GssXufB3IPZyEyAwDelc05s/0HoVSk+kBp7E2RRZPLNSiulMZvbkk9kjpqPmGajC
SuttFSlxptKcA+SrIaow5HETjMQnTdS9ajp1kdvJSlBMWgn3ZjbmptYinbSR7jjz
ntPL+aeyktFqtBjeHkUSao0FyPnFmwORYtD/rW6zc1Wda5NWrri3XNYO8KfLR5hx
uHJnbNU8lGtdggM2N/B8qufl2d3MV5oi0LmExvNrxLkCOHBNx7RSHkXBFMDFqNVF
ajkj+NJPjhRjoTIruMQiPXlDFm2+VoaPHRu2q3oZ3jNmuSIqCi5c1AAqGRQ+kvR6
bvE7PHmakoQcJkaLJeXMdGan7ZwEVr12dHColBzjVIYdLz7bawBs5KQzemLbkYRf
NcAnBdvvT6INrc6Ivjl0rGzvKh6F+Bq5qgdMLMaem6XL90uP0EhMsgQp0tBoLw8D
PebZ6Iie2YsqvLMllKvu+ns+nqeI4+Cu88nKSKSmP95gpPvgjbGc17uyT2v1lcqx
1xjv+QsRLtAGq4n8Kgw4Je0TRPa7xmgLmiBqLNh6qEHBw+mrKkFvrWdwC/T+VsxT
1RFnUH1lq1lpBd6dUDLUgbdkmKe9ovINKrRJsBzjtZTaOZC7WUxZJ0w16TdS+P2T
7hwsmRfW/Wu3ZdKz4ZsvPCiFfp64uMDUv/znAZVSsUNSk0K6XmB7ozAn6K758u2y
w9RGbt7lLXLs7l0oOCkRl+GjTTBzc0Qkb52LEAZ+kS3D/jH6zpPtX0GZF/V62W1W
qHWjnaq76Q/DNHFqtDKlVcS2hNOGJhKRkI5ZR99W+dVY9KYA1AfrxQqxBwysW6qZ
8+ogxCa9/nQlCXHJxts3C5kek21Aj0LxGtrUO7sNEQtPnvNGjuvHg8hd2oJ+J+wa
s+VVHmopqYjE0cQM8EoGIHuB2AZZYQNj43n2FgMvmPUmeMA5dA3bmvH5aSHI2HDP
HGAwPb5y3dYd4MMIZsORHo1jJCxL0QNOcDRy2yloBf0C6kW+KhxV19Dc4Ea1NV4y
rJYPEly9dEDiXTt1TWvPi5Z27tYTfSJu3OPLr9lQiDd7DlxGE26NgEkJ6DXO62Ae
Z3XgNH5UPZmbr+Ci+XwUJTKoySIFgrvH9kKE36YFpxPmu3HDutDYdJJuzSfxGgFo
uzZcw7oqPbLpsnkNp4ABfs6zENK1PZHGU3e2doPehLovYTL5miFGtSvchPKv+kC7
7I4qA1vBkux0RD70AO6sJYcjpSTBo6Wi1cGsHqfxtOTqvFOPJylMBEAKS1YrEyva
gAAtwRCaMAFRCPYN7+Pqzw8Aq0xxX65z7fX+XOYNMSFTWtkxVq9bOpi9m9DeD1BM
ieaynj6C6oP3TxPKey8k/EK/hwR63C3EAcZ2wJenW15lapxBywxdTijwSutz3DWa
m5uaGlR9915VPv//akvPfNZTNnNnd/BD8MEwfljjrabPDxTi3MkNFzw8Hs4eNawR
KU2SxP8cdgMrehmF5WeZhNOBbSI1u9L4hH+taE9yeiuuAs8CZHdLG7EOGY+mpH7b
L0pRTaLjnuKYknXlI+CyD5DqINc9yRbHvb6NZQ/JxEka6wqaQq6UPgXRcVwIq+cm
EwCx+nV2i42dhYbiHb+cJhVmjZMvOZPI+oBUTHp6QZr6kDIwSevxxrYovupPQeik
SuCVtKReFryVqnI+EmJPA3p8+oBnRGCIxGZpBMhhUPElznnsf7zt8YipI4waIJb9
bOxja/ucT1IzRikVN6fNxKonUoAXojnUfhSIc4l0oVNeY+IxQlsW8ERuh8CSOXke
7ZLLVpqink8TjurBStnS3wA5S9pvuQCloeMjfl1cAWdna4Kvlw2NAtSRXGjMJscK
B1kvZVjcvTsyGHuZ8eVmO+4tpApyoi+fxfgcVm4lfg78gu3lbburMK4Gkp7Rpq1c
8nP6K4To+6Xpukv42jDyKT48HEToyCkKeVoUNo1NFem0WDbhQoMbTNOxINWw+bMc
zM2QlGjr9t6vZ84y3hDCQUmEOqf2xFvy6RMQKz8jSuWpYmZ66tl8uZ20QSvcckas
dvFSABiDhcOVwrH46e+iz2i785n5ph4X7tbe7r1cpZil4hhqyktQWSpwR6X4Px9g
nEKxTr0DhU1gDvqU/NpJMF6MjOrRbYYHeTZaIOEgnaQe18vy/4A5zjfbtWBVJiGy
TCdx/UfjFiO5epuVjmDIcX2TTOG1C2aRpUwdg9Akut56DOZgqRIm0UG9P37U+B/8
/Stv+FvwtdJO910K/NaAT3iWygX+FvoY5tsgj8RJU62/f9MlyFTf0TbrBEyTnHVd
SiHqOVPDt0Q6dv/58N8JF2kTCeAMGpe+wyvz9yAiBSS5UVBuV1FxDxXIYrjNFx1k
2Y/ufsGKsSvzmfolYKCD+mwTm0kh+OkrJ1fgXYRD3+gv7irV12iPewjVg6ughoJ2
R4IZrjNxu9CSTFiEIPt7CnTR8ZpwpCTGz5cDWt+79eu6sl6PlfNrPO58AYv17IOv
JH7te38xqdR94lPb7Llr9EFwXgygpu3DjT8PVRuCNDYz85hKH2gd6B9lEM5UJL06
1GkU58fndVLbVpXVg7H56cPXRpd+R8/IIzbAtLP4n7QoDYI5fLyMtMv+7rQ2ilUk
9W5ziWhJfGFcbM1hrJNH1kVdJW942eQlUJWWk4vGC/MIFuBjfu2a2/vZZOuXnr0h
ysvfyOtAIF/c3iOzzqcyzsEQ0O6+diYGS/uv+9qSV5i5rIYbqrAMgCC7xt6Vv5lF
F9koN8NdvTfFb/d3T1ECN1foo2aKJ9SAoVK0H2wBIu1J/2y7W3hVQw10IvBARklj
Gkzoy/0VVff47B8rZoFuk6A4OjtOyfSv8NzGpP2ieQ2z/DVMMa3RjzOyL327DmbH
Yw322L4NdULei/7oaBpwXlplYapkOK8kv017EUmUg+o2XyLq1oEAU71jMW5I7ETH
6yYay0lkw83G7wZ+X5P+fXwnbWPvkLQsICcaigqiNm20NWwnrZ8om6cRb3mVXXyz
OBbjDHfGsEUS/jE9fwRVMjmT3xAy7DRRLlbWxlbOtxthLzDxPkAwxCijTej4UdRZ
ed1PrcqVij5v9SvH7qY/H8jXUI+MyritFef7ZY/O2Ih7NKl11dUBClBUOAjCp6Wp
2Bu0EbBMAV96Mvb5Fg3jyiuEUu70f56qtkGtLMV18+6JwS8dto/bipgZNoHci8Wn
Z06qdheC+kQ4v6XdB4BjJH+0r4UE0Oh46FWGsCnF82SaL3RMPXRb6wweBoZZlc2+
+AA75+nY1xznYm4DX6gudo/N5UscaB95BGLpxkasfn2UGVIjo4/YB0V7Ii0Ru8Lk
15y3G6ZNRLPybPXNRb8murhBQA5cxUrsD30hBaoIGprU5Dgly3cBBg+Qk0WVZQkY
FEv0NbzLAaeOOC3LsmTTgXGis2p+zAJkd/WVzl95OT4SoLvdrQbjo6HElLlIk7kN
KLaJs7YqqK+y5L288B5cMJ+BwTUvO1d+ubLOP1sGMD7lx2U2dpKQeQ+l5KmgaVuR
yARsE17In2AWAEw18PStE2Wy9ZdonR91EUuhvW1//b9vGbJxqvWgny2NzvE4hpQ0
1jWCLkoprjX+xIxAW67xc+bPYApr7+FNHNq3wE6kldtKhXVTURIiC75e+A+DiFSW
aeaypYsMD7TlOFJE8GKKBaqIUn12heAvvBIdGzntqOkuQczpp+XfitnAB3qXGsDz
0RSNZGLK9t6iYXIOMudsMOOJyVvTqhXGeIgMrY6reEkztXTsPbpx560qD0JaVKgQ
Ghl82qTeBNG3NVa8xXIrD86fYreIy+rIaui8G5oXkgIh2LFdoT4RnB109O2B2pgb
B18LbD0tkzcLzPUdhHXhh6si3Qy0dyu1+U8HM43OB3tzk2tu7vg7rT4IklTV1Op/
qCEUdkI0T9Ho8XiS7mawl9TGLBCYgsauBAQ43uI0cstkTMJSPmZMYTNhz66OcGXI
3u+i+Mr66+wgB16l8JMNmnrN4TimoAACTphwGy2EKWnZHDI9Zs83yLViFNj4g026
UjOu2gx8mcoVsD5zgXzPRmvCaO/4qRwiUASkHBrSfqh2Yy034yRFMVi2OOA3s3+e
fzYBEK80jN1OEcFRCJeU6kDRXHZvNuRQkMp10CvlBqRkbEKU1w/fNwLppc3ElUSB
R3R2g18O11vtBkB4ziWXICwPNiafaTxEpVoxJxwGJUu15SwPkV1jflJ7AjWkF5WU
TUN/JHWSH1bw7CwmT1ccbaBjBr7byk3WYWxd8Lt9gr6jVpcGoa8BXhJ8gqqxVBPI
SpL76+utLkUqlqN7A4kVA8boRBn0SKCbu+lehmApIxZTz0+jfe4jpaBmbM3PYoYd
YtpLw587e/Tc6j6yN9eukIzKHFhAEPd9UFZ2AKVsi1VA1E8eBvcRXEVH96F+/fPm
gXaULk8B9hoGgnYUc0mAAWaEIuF15ZwgkBTh2efNHW8ivn3YPn7SyZjjfKg1rYDI
3HYO4/+vZ/Fan3h+4FVguRgDV3VQSDaKzvbFq0jEn+8+JdwzfLfp1ywSk+hum3Xj
TiFGMuTSmQBUinTkGR3QIvToTVbLH82dAdHZNv9ROWVI6WXsoNOjG7MWwTLDciIT
uqTTbgoCz9yz2f185sjLgnIk6Y/ZUw+bY+ZSjSJZOxyf2subCb71qZTPlN86zzkb
Ag0NrdS5gTvJerRI1PHjceZCMDCqnXpKMpbc4nR0oWIQpkFlIMR5znN1bPlmJrp7
I+foMn0ecRT+Z5egmuc0jU35+x6qdj2ddi/+tmf5s0sthzbrqUyFd64LgB+ert4E
iAxZVyebi3lu5SHYuQYNpMd3KuRIgry24CdCe4DKlZz0XsQ5IPLGDY/rDyvHJGXS
xVfEIcOJD00/i7sU2YiSGDs1JNZjD0M8C58gxAAG5w0qTf4ITDp5Tl050tAsKje/
97TTWrp4NlKgGbYqVUH7aJ8kMZVGG4oBwwsj9vbiMk+fTRaMf3XZ/rvntc634OIA
ffWX0IJiyIVjQh7Y4FxT3VzSx1emwfdJoOyEuL03BDdr6nXfkWPCOBvuAvivOqAs
f4J2PYcI/ysCSsMJUgNS3Vk2lkHieoIM316dQxUl/NJdsE0MJU50PYrwKatImTio
ozi904Z1MuocHN6mB9zuetnSFDYopGxJI4dXIE3vfYtzlfhBI4Fj/tlpp29oPTiq
ZZJdHIH+oez4wA4snzigcBrSmkAyDd5bVTOQyh+ET+rT7a8gSsj6PkkGcdvi4ToS
2w1g5pGa3I9IEjGa/yn2gnnlrDNNTg1gq5jU2/aaRiZYwMEwrXHb8dOiLE47Bpdd
wk9tMgHZNipwMhN89o8qrj9tPBqMym9almWKlCqPLXvfjwMI3HsHySK2/7GYYBYp
VyEASrGHBxUFcoswvb/Qe0JmN0Lyf8yX/wA7A6yQprV6g5YPxdehL0yziqaP8xkr
s+4H5PO3YT4bYOVA9lqqt6v5dBzJpR1d5yQYhIHctgh04szRnt2EejaU13uFb3nK
DI1wefWJRsy8maWD5y4leMDdw2B2KwI0STQq0t7F4tQDsqI+e3a4RS5fXZqMx2yx
SGDnEN1YdAUzqfntuOpx5dmNz5ZXOzRi9HfIuEyXaq90AYqzQVPLUCDFoiVzOnRT
DENwQDTcOvRoye48PS5MxUG4VnIyBVAjtnJ2rHXwhHD2epcShjaTY9xfbhwFG+gV
4xKnTl5n0ZGfs895t4PjhHS1lA/7p+cYPxZwS94nlMM13mmqlvMPQZ1uloF8oEsf
osCj4AzIpwVuwsWKWQgwnoOObGm8ay1jSxwWktWHp71soAzulohnjoN4YNHjnQSg
s4ESKvJ+B0T+MC51XF+sPyJUYBfH0f0y0+6bbcbw+h56H8xTVIP9H9nBbveduXCz
kM5ZJe3yQBVenluK+HtXAmFLjzEPEnhQMCPCrwYqk5ovWrQ7jtvnT2iz+S8ouRl5
UdOZjjFyRMgLGbA0FPuvT9vMSRgWoYoOmboorYHiCvgmi3kRgdw+wVuzf9KY4i9/
eD3YBIYLzitqI8karIRzQmUrcjBKe7QRWxZaPREHfGvsGcsPh/BZYRxft5Of3ezs
LjQkIgxaDg7qHsJf7pXmyF78m5Br6NZUW8y3zz6blTna6AyJFjqNlK/vqO+anNjg
eh/eQ+4VTIEUFZMcFaJ0vxxoAJkKA6XAIKNJev6BQZYl9IrgMpygNnKy1aqdHGar
RuOvVRnb/T0FCwPXIuYkpOUXpatTvCouU5B+Nuw5aAidFwmA3YWaRWKfPzekEW4f
EGwoXOpyrLpZvwfbHd/9/M3OFMPHRaBIyCG12kP9mMFP8JJ0jV8E1ANoeT1sB7nm
kdVEDBssgE0Szb2vYV56udVLvd1f0oLzqdb/kxt9GmlRgWi728Iopb5KnU8WWhVE
Z2gCi2xf64VHlIBn38zFxi+MBpp6JFqpjHJ9xQmlftFWCs26jfGfF1DkOIUTskng
EglsrKOOkBg4paNxUCaQC5cBRPDQJv8uj3vq0GQBnNeNS37lWXJk7GPTXrsFojaf
PwPN3wDn6ntHcIToDKAuR00zLfFZxNPAje0msFiu0U2QLOYWRWmS2vEHr5qZvMhB
2obO/iNAKz8bk4NVhZlHmr7BsKN/ATqdmXkNUBvpZs0SXCAZC/egjg5YQX4fDSYS
wqjcCIOLLEEkBGJQPJ1qBRyamc6kf8Hxs9w5tsUARBurwEs12Fuy0WdD1HDiWILD
/OJ6Hxb0lrhVNYEqQkAofKvMnsRWLP4iGtgdDn7CZuM6rPGyXU5A5mCrEW9MtcJV
oPzgfHJzre3d/NmU/C1QV9fd3wfVfSpNbOsLqwS5MRwDrG3bKyuXLW7XpkCMWvnO
24gWbrfUGgprZB/+wLZSS8LTI8X8QWiYMGeze1ZbbTfRqRzXEjY2UofdePZUGmt1
OREH08CRUQkEHg40NoGrR2hEYCYo4AbtlN8xIMtVuEF9M4oWZP7eqRS2yoq1mVOV
ixzVLy2E85bZ3LZnPGAYynq4Vv1TPkOCoOwkFXVysx9VhbCu13L9Gp6TWDL+WOmD
tjjZwOK+Xj1T2lt9MBXku3XRqRKu+UJVjABDJXkc3+vP4eZUhpwtJ3fKpdXlLxII
jdFeJQHUncsCztZqT4b0zVMkRqTUfBxpBDg6ryh3IDdXab91WZG17CpnyoB9RXAi
H9QdE/KK9Zw26J3zBxLDPE+KcPFkApXLKLeStAT8ZAW1DAjHS3tj08dmT3PPS6wX
wqjoywdArMKmSWSYzIb0sjF1/rJG0TmrZg63KCdcx2ViNVuzfta581d8+RnFbPWl
93NGE26Pe0INAtGgHiiZQIJjFoEAwnksV9PUd6vwmJ2zJ2nc0J0Dyu1w66GZ9lAN
xmm9xTasxGrNz3AwUyNWsXdb2+5npLQndzvsNYDoTGGQ1VRMKWb0Z4+8zGrtHOM9
N4drDtSF4O2OSauUONOSBQksmdQYP/b/rT028vM8rxl8pc5/ymFcgYiTCENlTJo6
QNf21TQZGHZDk5mYzViwqkj9uNG03UlvjQJoA5KuVxvxu7VqM+2uFcztENU/DmIu
xwQZQpo1n4m2cxPzR0vxoOvjmjDwFJehmyJ2a2/AjDZlMJUt9nvmUpB52JcWh4d+
kXAxWlT9NAQYDaKV2OShHoHke+rJ40xEVrDyfFZJ39MPQx71ty7v1C+IEx55vta8
cVaP3hBKTRjqpLuyPA8yCJrGH64jMxz50tPcV2NnZ+/NZ8bGP35/boeFff5IKTlh
zW3DpbvTrJh2KQSg8kIDu1PQgTvIuYlR2YsuqdPsO0sGn5NVceSe+BAmXxflXfpY
RKEEGJWzGCOQZ61Pt2sP6xmumr17QTWL6BAlbR+pb8gYtAp+mJazCO7EJ41sVTOj
Ly3gUuxS1SjGDsn1V2m9cArzl/7WSSTOm8dth+g7Zf576f4fcyFffCHyQ41NYu1R
HPvJOMs5SASTHPVswugRCotHDBU8DRMtRENDirHpl6Xt1ofa4kFVMD+1nZPmemzq
HifPKjXCgk6p6l/Vgu72xn75qH8jezbe2upwBPjek7l7P/7tw4/L0orQqFjHUcpI
/KgMkDdF7/Q8QCoprHUCZgUP35HvrPKdKpwCA9yjgpuszZRLBGvrofyygKXywHDy
SkBz29XUXPkbbV4PO/0Z0uXXXL2SMlDd29zJeqqjRg2iLsES+zApJzshsN7TMJsX
xQPtA5WUiuNhuo75PN8CtM01j43VTk8cyqSI6c++1K9jXBdhm8bIuqin8EvRnl9B
094KI7i5q6x4n0dxyzgQ7s7vDsmf+RcHpV4uYTDnSh1JZpsOvj2f89QCaLyMvwcV
QeSOARz/vkhnsqiUyRGhWws/fqWpvov+mwBT0cfEE5vVWInHriqJIRcKiVJGb81I
5x2lLLflAtTBSNRxqNe/CrsdNBbJqi2iDGpvO8781xCvQ3ZPk8h4VbD3nS+UMwms
5hvFnlcMwtcKoyf92aszNwxTmmus5ArdqvoRCcwnCkHk/ZIGwiA9cPX95xJ2gfTQ
BSkU5Fmq0hrpTbP9z7fIiC3yNsowsUcvGGj4+JupUgNBC55XgoXvIGBqws56JID4
nyBvM6i7hHjngSHu3Wydx+euUk8BxMtRK2RzNoKyEoRQPfS4uzpCTAj/c0CcP6Ar
Z9B2ogs3i6K3KygbDorSEkZIJ2vSGItFLn8iBJxuSDgkTchiJyhg8wKb4v0C3wSS
7xijf5fzXwZzDUDw8CWCPUe4/cB1WbuwHrqemQ37dXLNPCXQ/R5QXhFQOlpfKYoM
O7fOiTwftPF9XjzCeZjt4DVazn+Xl505KUEGrMrzfMncJsWrlnj82pI7PUabUVJO
8RYcBpCGk0dQgG314gp63AbCNNoc1OdDOxYpYD9gtpDFyCVTAq5GjhvnS7lD4QgR
BWKJ9yU95FDdeJwltVuz1SajImcbKI0tn78FA/5k4YT002ylghNCPcHH9XCFoCQr
FUACnCesoA58679cIPxQIw761HKAlxxFiec6NvpoaQgP4PhJUHZb7gnBJlwrNcts
1oid+YmmpkxWxL52uwP19ubO2By6j+4SbtdlvF8m1kDPKxltsAVhKayzXJ1+fCjS
BvZHHCd0vyGaTJHIda/i//jfe2PlZFOzidfjvnlq3I7EcLC01WAIpFbIMFh0Dqc1
VRX7V3v2LVTklVeXzQMP8xT2UB/qtSoWsTCx40+PqYo7kBnA2zThrGVcHXISkaHm
Z5fyqBhX+Ad/2SvEB3jW3gvebA+WhkNglO7kUvKFHLuhMSaNrvpfiXXuPlR17IiT
nMKYCLcHBeBb46UEL4oTpiW36VgeCRKqw9f+rXEeJHGZptMVUzbC3gcMGs+rGhoe
ykxvVPo205AdCw23kQosyrr/+29v33aL8+38EXEQfwtpeFypb+C/2FpP7hQLQa0T
pvZMeUfmZ2HZbTW4lL2SxpIMW4Ki97C8Jh4phNCSkmg9li4dPYVTfbVpV1+D/73s
D8fiu+I4n/Vzt+NcAymYdnU5XbzGti6wvAaGU/mz+7s7bk+zW1mSfUzZ3WNUpusl
SEFenTW4nhdmE8bBPU2zZhnGah0qFUk3DIc6c+thyGJSRCPaSTmKQR+ZGcajKSvx
TxoYfMvbLsuer9VpXsDAZXNI/u9QjIpn8SoT3eguC1VnTxKqth9q45akGMiMcEb9
P8CYuYU+NePrTTJer/cuUdbNPwuu6Bo8IfYGX3QqlUtLy71u3pgxd8Ystlw4PT0U
Vk/w+Cy2C5udYcPrUkw2FI5iEUKb2hLq5/5aKdYZ5QE4QxVB1fWd0uTv6D/8M9sQ
JFcAbob/k4MzYjOid1I/dwJS2ozJwUWk66D7Bt/1KPyszZOq2izTiXIydMH2DC0s
eASae32u5bVl87q7H/7chkb12O9eZN6zEdAPUjZYYGq7Hk7H2HvYXtZ66RgYI3mT
Gtr5JICjd9RWYyb8pDj3q1/lIS4DZxUq/4gEveeJR/s2yu/VRqDfAb+/w+27Ascv
xs+4uDQF2mFgqwzVRre455knYXUAwVeRmIcU93ZrwI/KcANcOmze1k4cuFkZqsHL
hSP4ZcLO/E80BSJeJxaNldjjkTuGw00ZcitTXtB9/fUsZsyCApYEtakpwY98q76m
VErqNaIIS2WEFnw8R0b/xZRLCv4hUHf1FQ0oK76IEp1tDnMccuDJiEbBjixxFlfu
JCqMPbYkevRCA1FH7dQik9gAfKhHUUDcq/9R3h5sPCcvXNKdbm+ncKCe9BkYDSji
a98paIFV9KXVirVjkzTo6ZYgEthIDKbF4PFCyDttYGO+zBTNENO6IJvqr+4Jbo+F
ZYU3BCQVPGTU+HtcebJZdAOrrcDPr6wFddqRcUJ8j87LqwMWkytQEsDplX6gvO/O
biR99d0I6Qv7wxoPAwKLV0/JE1qM0b8DtxYGd9cXoxz6hGqrPius2QWfYOc2bxUg
tBYcP+8RszJilhVC3f8LV7LvGLryDM8NTuexWMPmUdLNPnJNfB8gJwMXtTbWD4PN
9EyA3TIAqxaUgjrYsGY4+afnfG3RLqvpDn6XbI8salO6euUaNy6HOlHEJUXds06X
ju3tBCITb8F0TLZKZLUbmgzc+IXNJbSjCyszjsXZAzgHrIncJx+I+MfY7DKH30TT
mmbeaXsIp+E0O3l4gSUaONi7WFA+Toih97Hw5rS+nXnSHY6qCAZAS2IqdPzXn3/J
qruA0/jrsJY3U4GzetADFxeDHrM7WPVghUM1hGZgxfVkK/cp2X4NSZOiwIj0dfZg
OesSNQW9DXhAiwA7i6yQaUt4KkWkkKQQQN9sx/fnoIHJ55DycdUdl0Ttp8hRIYQ4
kDz16XF4PrqIaWi5IrbdQMQc9ltcQFLTN9Ps1XGM7GGBQheskkVMx9Z/PORuF1ME
ps1bhSWE2YBlDhj1jTn+7POO03UiZnu/hRHWawRAsBvUQ9W7LdraIwHBdcVroe/Z
I7dsAVC3YpXFM3vfD8klmYi7QSz7vU/5+wtzuwrm7kI42mDRyouA5x+W579u63qr
luVtf5edJ8AmGN18UotFFVn1IUsMii302YDr+G72VbJ904bEnkm7Te9vYduPz15Z
kSXDtKEgliWpTP8k/3j6Of0KSz/fn+jJXQLfVsvRKa3QOBnMIfc9yolqeHZZNDDN
5rT01Wz24wsl0EJ7U/jw3EnKR+oYoWfPIbcLIxABV9vJvSuaRA736CisDsioZQp4
L8QpmaNEYewMYxcCDmJBFqk2HK+jASKXBNdUe1ceuGmqrgCCEByhLD805UPTmFs3
G7iEQpQnAkXonEEhgWryC01eYm+U6vB/vuSdqKk2N1N5fEuqLyOullTkyeQNoyKb
DmAvqpppfwzi9nPD5v4XfMlpV58XVSSoUmj3o2gka6ChL2Uuymt5NWi/ULt2rbTJ
FQUCWa8mnP0/uZqU4xyh1YiTYNzavXHiM7YQy/1JeWZbtxvKt5CJDX3iUC0VWzE9
iiRLA6Jgi2YAjt5PHaKNspRLlKNuBbaY2JjvpTxlR7rIWbH0vNAmKgRxGmMP0rln
Q7rSBboyWtIc64+0j6MpHXUftxyNmr9yyh2/VjRcqTisqjdwPTawrNfLHIWPqMk9
TdP0abEDACGhRSK90MG+Cn3vfIYm7vGKvu05iQExR0oVX6KaopHdHySYOjtHLsjP
+mkS4/3kwgKTUJbzOswyG5bPChna1WBhAS8jvB6VJzisBGqwYM7TLrj/yX2q8NX5
otvu6EsnmeZHyyvS34Rht3aRKSDLV+hLydqI/uEl1iCMwSF2f0dvYGkXcgUtBnXk
X+atKRwrj6hx7NwfXVHKC9DkOL6IWAzrP9D3X5AsHj+fiyRX7iDbPapwRxJcaJtj
tGnliEL4tjHv3mspdZP7TGLrOYBe8VPqYwm88ELP9ZwwJiqC+zFdm+X42Jjbxpxd
kEqFEyutEd3Gbng/TYuj3yrUIWhgqeKO8u/58e4TaujdWFkn4mfsWBuW9gn3LclP
793WOkUbcPMX/E5cnxIqjzflJ/8mbLy4CwLD06PLouoTMyxwb2/FnTTwUdXXmyYG
8/nXeKe/GhQKGNKLdIkV+dbEtex/FoA+UTlc6e+rHJzJntxluGDePxzzE5nW6Csi
XeflIErq1WAP2bo5WfYTaDUKkq5k3z35eggAuQeTHd6y5V9NK8MXUl4UVqqAkm2O
RL9vogQoEkzzPsNbzRiQApuB6luYFzeU6r+o8dpkemrFqqK58rytcFJJqdCpvvN2
wTLa3bgrTQjIixgyuSgTxCdndIYdG6vBbG0zRXfAJxC5osTDFGn6eFyrzElUMJBa
p++vi08pRmC2i6YPe7xSX0nEcIyDE7A4rldSZvovHgaoeRf5AlXGrmpz+3M8dOAB
yMPby2Qeqaopfn0Qal7UpDMrT6A6ETMdWwWvTPxf40hXFfrDUm1+5fZqR8r5pejy
/7bB9WmL/TUffsM6r6gMUFpfTo68DoIaYRwZwrjzxV83RLOYfsKLkRSgDdUAGObX
ZbEKiraI4Td5dGGUphcQzvf+X9a+MyMz74IptZXIHr4cxO6p8tVwu5cxXRo9cyLZ
Zp2lSLu8dgNKgIwssMsz/6J2d8tRYQ9HUTkmpLQTS9Kzdn02xrNqkgM7xHZ03M6Y
x8952MW3bbbPoQy+b5dBk0gvhkwRruoAB1kfIsYqtdkYEeHB5Q5ix4RUfWsM2meA
b8FZOFDLW8HHm21AKdbPC2GeYldoqkuHWdhdfNk55x4eZ1Zf+YDYUQKVw/butvKz
AQLbRVRmiMba0nZeI8yKVhh9cVGOmWva3SHAe5tGr8SPcVvx+Okjqf8t7K5aHm1N
gcPKUSOByX/ksKJzhawnoGggQR2ZLAhLb9iRl/i7iBOXkJFhEVmwgFrtK6RzqA5s
cPcPGZn99nJQU1E11iESAN3XncQL1HAyV7CjD+92wvgKij0nFB0mWoPZtMExDa8m
a8s9b3VpE/1cNiz9dzCpENFxC7nVqNRediozUhiA+NoYOqxzWjujAspAnDQ9XaIS
cAd0bSAc8OB3M0QvbDoZN4Au976Qmx+54KDfG6v59QzC2G8NzLxcyDsLWrzqu+FF
t06Z1DQlDN2pTPHCo76qc6dAgkLiQJt71PtD0EPMKS+Om8AYbvenI1CJefMddYCg
dcG2La/7qN9QlRezp36ftQ2mv1jmXDQIh4MJMUbZvBsyfZ7PvtRTYT9B8zY6+HnG
sIGBtT8iPEEHpVc0pr6V50OG1hKRq1Jv9SQmDavp9mb+JjylxbIrpxoGTtLIwzuU
w7MoHI4i9+VLTQY1XvTuYiYgdR8IoWXLH9q7CuoO0WigJlmDSMnkz/y2wnNhXkbd
PL8P0JVcVFZBnQeWAx5P9Q1LXPAxQ0iWwh0203ayrB+wNCQ7BRswXvXMkW1SBTal
DNv8kdFrn+LcZmPzm6Lu7FKgtkNoNwHmZvJQT1fMqR6hFz2Zk335OWsZXuBF4J14
7fP6l4TFlRlUuVKQVewMm4v6g6ehDupn+FgRHG0zCfHA8qby/ahvtxvHrebUevXe
zWbSXODtA+tqnvQYspcTOf/gDp4hfyoXHg0zBCyT/Zj0eI7pjBMfvw3DgyPDKS7S
B7wTYDOLfG+c1TA4g5Cab6OTnjkBKWtrZiIQFjfjiwbugfTnIwzsvj4wjTdErs7c
EYIOM20THoMwGHkj/DP9ptfxagPmO5o+G+4G6JnDdIxlpLv+0k6JdnKlVf5Ox92M
2Cu3rs3OLhAH41SgMavQrWNuagSl/5bUzFrqix2Frg+yhOKQNhAb3XecwPADV6QK
iQuxDncXzVuWPU2S2gwIIYQXw22jmvuZEHNF7iOrMxN0oypGQ4vtPWjx7yT0MqAK
puJLLEvhiUTDiIj2b0tZfY/y9TLHxjjBauDaRVRbHx4JRVYWJmG3Yrgh4MCWD/WM
O+vDPgq4bnIPVGZAFJU7B0Ti77kQphnwzoNkwnoQmnTG00aG/YHimqXAKCcIEsQ+
aJBS+drcQy1STYC1eHrlco33N+FjOvWOOu9Rtum2q9Z/qcrkWT0ELt5TQh+JzVCZ
gbCZg3GL7Rbjm88EroODO0IRUoyNOHJFrQIxEBUV4hxEKnR9j413KzktoJFoEK12
v+l8Fw0ms6KpknovURevAuuHwnR+hn7ZAovx44PXKbAuSIWasB/hnoF1tqX4eHc9
XE6LD0D0ojpbe9+bb8V4X9WbPtzIqzVzhYOarFiIy8s3A+P99qs7J9+8tJcJagDi
31dp3I+svlQOJCALoazCPlhr8gXVy0BcynQeDo3gdPkBmpDAMHjsl/vPJ+fkYsQj
Q3MF173FHOq+2s9vQwYiv4twJ2KoOGejV1nRDUZm83B2Y3YoF6/mkazCf1UbsSTQ
L1jokcZlOd32MopC9fi0cfLdXo8ya0Xx86WOCLlCGBqYJc8OWHAJKrLSJdygyfZf
e5zao0XsCqmyLs4xknOemJV/HUeGBkUj9nCt7eE25SqyWkta25T4yeaL/dWBdRn0
yqIkuz/mxMOfklp4vCZbo9wwCVtP8ngDcsf0d+9VGO/A9gNO/V6F+Ez2azP6+sZX
fy2tO47p/jXdrpnjtiml8X7iLreSu2zp+gL64rQG7RElW6cBiEysHzo8Os2zDaWh
UTEcVzEGJrQnlZYWGlyVmyf4b3hreLF6lw5t9xLNpDEfSDz3FAQgNMWbKnhTVmTs
pax9HDfEoR2fHf/sR2gUc5/nxn6f+Iw+HgA1KRGi8UUKzV0UF4TTd4WtPoRKXfy7
tmFDAL3d5TRyhSEO8mLtW7G1Xzm+DdA3439L4oo5u0cUra4MRhzCOWVGCur+LsCy
CfU2amkPPuKrldFvj+jt5PEH/LcGHRb1kPkSSZgty9vffo7gpAhvvuNCez4uCJt9
WkkpN4FXw9+JkT+bGcZOdofNZt7i0/tOHxKrWn5L1NXgN5FWNT55DdbM8aRFk6c8
gAGD1BJGvGQNNct3sx08CqU3EjpDtyky5D6ruH5p0pKqqXDCqFANyctDWGNNM0Oj
mvJ7NTyeTs5myIKTiLrJYZYE2Zme0ff/yYuymuI4CkteVyYWuC9SCbmc5SAwP86S
Odx9kgcqJtiwOl/nCJlooIcJGd6GIrRr/JM9wmhy+VOZ/GLsdB24xFSk8JCeFJOF
3DmqZ2s+pnYOgz2wdgggmYrouJvsuDZ+Rkm3YcNpwC4Mf5w4u8UWVqH2Uztd2/59
rIjDal50AYw7xB1yNAm3sbm4QcWWJlhc/DYMofCUvlZdjKXd3Y+gthRpO99SgAXB
I1bwYsPwi8WNctn2ENO8UPWv9YIY3RPHy94ZvldKQtFN6u3nFdJGB8KF7WfHp8UO
I/AfEDRTUJDylXBLo42AfTzFgOtdR5lN2OsrZ5N7kWEGM3OfJO3EStG+7zbAF+YK
m/3QQkQXdPeqiHbZO4a7eFB9WsyI9tMRxMtFllbQ4xd5ReERIA8I28ySOYaAgqxV
cDGaTB2xFD9GuFR+GZhVc59oqI1RaSMTD4yUgjPWb2R8d9VvXp0A2RWOCa+QDbSQ
8LbCClGxF0TQMFm9oypNEl4Fmc7HeS4j6qv3fvs9TDJlAOfWhtNH4lpoEJzFHLVo
/gyRXi1+Bg8VVNZEqf2GyDdg3H4WcQITW0p10E/GVn3Z4NzCpRBcbTLGby+/T3be
lZohmCBVwnjm3fr8xyK9ZHIY+vZ+se9R+vKz+srSsuBqDSwkqjzYZIFKhLWp5ven
G9wZArV/GEPXZStyJ7Ruj6txmhtCAjJi+n8wimiIcCL9BCAQaRF7n6oeiLjRWXWP
MbtZkulHh4TmgK2TleIdVqxKEzR7Pc+A8dt5Kokr4lsn/zNMYK5rRylWX7P8eoQv
ejNsc1EsuaxZPpLgR5JBun+0s6Cbqwumvc8w13eFdqvnoggdEog8KhhfYcMZH2/4
WZLyJK82fbWqPfKxKZypTHdztRKUXgRXBZr9SAwROdSvw0/StuP32+Vhi1QIfzQ1
b9kYPxp094gin7wantrtSe32KGyU83xUDrhhyfGoivq1bJ8N2o4eZn4QdS91OwIQ
nSbBidHRLg9Vh+o749hkh6lsHitBOA/JCTAr0RhujcvKcYexD0qHY4kH03dS/LPx
HPFlIwuLkhkNhkGS5r6WTrJGALJyukTIiV+oc94tiUw0O3Hw4bd5bxz8z315Qxqr
28JcCBQ32uTEpo+KlJh4i1Nta/MmRA2E9cQ8zkXMRCt4RbxKPlDQRexCO7stEDqM
UDdeBSsxAAqOIlOLWJl1ULdBqkx9ESnANF/ag9NV9FRF61iEP82Mn3qTCYghpYOr
1H0l3TT/2kZ6hk35Duy8uL4x0N8HG/5AEhBrVAYiyKsLWHVS+NU1VT6Ec2EBfXve
xdCgv79vSFhhvX79upvae6tEzTaLt8JdIsHjnVowRsywn1OUJKEwV21Kf4ffnaY2
ezsPeaq7YLMCg+2qmYxV5jo90Kqx+xoermXa3d3ROikWTzu1RGMUYquPn3qNhA8O
l5c3H1dpHzWSgSxx20y+NehcBFUeqM6RJGnBJv+iYTdB0BB8giblYT2fhOOfncJ0
quZdQ3Kjy+c8ej1wwpLQTSYtOo2Hp8y+zyJeDhg1XjG551YawNmHh4R++x4VBwQJ
G64gCwwY0sBazH7ZGKPXXO9d35i5eJbIwnxrh1x6qbWuTcwpFZmfPNq91qfzqTYt
yfmmPXzOdq0Ba2UyvLWzmmqERgX0qXe6DpdDjnG3i3DLHEoTbeGyUbu9vTdjlj1k
0oHKNaigL9D47eEXXdcns2vZNA7NsnhcOQelEXCO2f6zqE/bLudFITboj4ciP3nl
5bx/DNb2IMxyorst2tmIg3kuPy1ZbhHfdR/9X5wR/9m89XjzBhJy2X5l9KxrW3aM
jZr23qY25LdMxIfdoOsx0kPU/PnVT6SQmJ9O0ICGjtuQTydMCSZjeVqSPvswEoqi
5AFGn1Tb/L5I/HutMWfDfVA/AZH2nG9YxFgJynnimXbMrSgvfYn5gaewP7rUmYy7
qHB7yFZQPq/eHHomRxhdis1KnV/VC8c5PpmG/rJBE/TnWGm/D8LwoHfP6u7E+D2Q
Nfbg/WjyAG+UJsAqO0H44HVupaZi3gPCilfadSnSgrrlVkGKpV3JUrVDaKBMbSsk
f7Q2IPERUX0B1Jt31jImaJ2SJ4b6/yG17m0p21BsC1aXqxLsysCygniNFFkidWJM
+JJRlKkzT8sL5KHHaN/FRvW+T/NjGk6amY81NMLJNdb7bdD7rqyCdWY+yFzgieM+
lA/XIl6eAcet5oec3ph6K7Y5Cwzeon9EvXXsTgHSA6V5dXEl76+DuReJRPInqK2r
NRGrm59DYQvtrF0MbYXACiauMH34O4jnfBREvX7QqQZEKVzJlzger631v2laBV/1
8LZuRH188+DjqO2pj72doEVSgahNKi1mXodCk+bFwE4EVyxvDzsS/Fh37fRzc/IA
tGQfPjgIG4nws7Aptg97otOV6wqrG81BA4yvvDEoH4hjPfdMMAQcv+Xd4d+sGdY5
x3mws0PsCb8462vQRMdAOigYVVXAbGrIfymt3Pgo/VbXVLnn+TALwELRhzc9Bz4Z
mzvuWoDyxLr8W6nNsZbYZahMi+OlMYcOm1EHVLsHkgN8MBqQP07rTBVfllIMVw45
Z9SREhskVqE304V1EHXtAp6bIjCusPsPT9h4OKdiLHzXLJchWRbDdEammlsrctb6
lAUmXiOBQPD0F9rjMX+0rr6O9QI1hfwrt3s9d9s4DQVRr8Hkicdrw+RHxN6pUB7s
a6nFDsoxMMn2YPLazrVlbhdHLtcdM2ZRhZaV8Hbim1kY7Dhnhs5MnMl5BGGwkHDP
eYrvOIAjyfiPZUa5Ir6n8qDHPyJBtfNdnXqwO5YFXtbkK1gTYy5O/nftxQBkaOBj
RhaWFImldCZpomppHfgLvd6XsK9QnCNtBIq+WlYrKWu//YJt2Vq6wA9uW8HCDQqJ
CK1XZEWKvIvV9wtW+DmfVHY8uBIyu+GRx6P+F1W5WcHjZMaNkUlXZZh0uuRzjsSM
CR13fdS30nyyweuEXbFTfQqls/dJ5IwPfXKYO3U9m9xE33F7nMcOkC7XiQD2o9lr
o36o/WoyPJptZpgsEtKTE77boUusoIjb41I3nYQMIZbHkqKb7OL4l1Ko9JjN6eof
AdhG0HH0Zce1yBvnnhwNSYu0fdXXAMP0Ba04K0JMXiOC2Cc0bWut9s2mlsQVzsA2
+a0aPd8FgDaXntWpDPi0He/kDR4cb84DWNUN/YzrPBu82JO24FLeL7ta33/t4Nen
rOtLOOc+vo6xVMeRd/jo/grnra4VF+hvutP+d1F0tX5wWwhyIfNaLFeK4hO7H7xm
7V+lWIFoO5avpxn33m/xzGbyqdeIxG3wRLBSzM32TMt91v4AFO3J4Z8GWi+bnHXJ
uBwh0mNrda1sIiF4IcuAGkUyq/iYs4S+kYQvMCcax5h/8pbTZUoDErA2ovaDjCsH
5BrLSvssEjASZwsfGbUnLBT29R4bJEqEMKO96dHGlzcW+aogO3BqA2D73mxw7viH
xjDITANrPcywXmlyGK2Nl1OiWevnF1fMSEsBqTEt7Bz7zx7ckzE31J4z4qlZhc7W
qLQNBmnmSXCjAmawi+ePxKYF5/YaX36Kw9+rH6ChwZ7yCIPlTrAgtCogwoxJCHX2
UyG5m/58Vg47llZA2HUc6/5WLY4JGx8o7gdDFmze59sOV0Kvfhmw8Had/57SDAtY
GXbzNsnoGl83HwthdQmMnkfTt+/sphcqRI2k6HXB0mq8z+dEdx8qr4fopcWY+WBd
7Q6y/P6AR2VnND9hEtiY6M/Vcn/e7z66fqVVFfBajwS5ZrSNKJSkEqXvvrJG5x7f
i1wdPnxTyl43jvxNt7mAwStap4Ij7Qj3FuP/Ygr6dYUuPqwisi0aQQGg47E24XqN
//A8sbxur63UUExWgNctXL6I+41TXOvbdm5hqZFkFw/0r3U0FR5/cpu5FAHJIJbT
ANpqtJ0w04n9TV6LIoCNwp6dA7P7LE16hORsAOXVslzvs7YHa7R7H/3wEuPtlrpx
r7cRHBwRcX5zmr+2xUfnTMD80ZZayYQTi7f+g22Wc9FKVth0V0+qG2UymwrISnFz
Non61LO/7fumCat8Itxo2uYGZ63KX9SIpo/jnN/B47/W3saxzTWqQ9AuE/ttmEvj
Z49ULSEVsHLTHod6MS/KjLRRfIOQH1KyY0FMz3AAkPX1tK6J6hVw2CZpFZSvVyO/
nfjYq3KLsojqWWvKVBds5KXOc481AS6Izx2f3KLjle/3jIRsAkI7g9OooVPL2tAf
lTj5/5UmTGH8Ww+tUkOfFZ+Rmk3GbHzV6DeGcqwr2Stodk9aT8izjKgr6TZvdLBL
TGA0m4iSb8xZDvKyAj/3sKbusxWlR+f1CclqEe9PuvtGsNBWpe2ctSB5VqAE92e9
bCYUtG7ozfkKzaizR8g2CsH/TuopjE6x+0t9GFyBnYRG1MFQx0Rw6yGgvPMtCP62
DQGVaMQ3FIrXv90Ay5DTje0L7oFnVOkvu8cO2dzX0eR1DsX7LO0Rippp2g6/yHUr
VfjIBZVg870bAgLh0rOMNrbZO5d3uwqYXllHJaOTpStF2bO50sReoEV2aCP++q5P
UUN/1ElnvYX/NTsJVtGF4EC/3gkpcLv9HR4TlZ5xZev/FYz6gfimC+eS1PTCZ+5l
fdKN4sfxzwFH0p50UPSGEGyAcOBjko5GDEYftpiWFdTvN9ZvKDYbKKm4AzptmFJB
mee0PbMQNa72kxjzyODZjursevVNIL7BWxvCIBd0CHL9Qrmcz2TYqknorsg+E1XY
1y04V4IkY1nVOxBeGB8D1Cm7pCSs7leenX3x8E6O78xTMdPm3qICcJlmmnKXCYzn
zlwywkJggcOl26bTYn4uvXIfQUxrbcxZXMXlkIvVYGM+R/tiHV8jlSoeSHJJBvmH
Hhb7k18La9X3HXuJaz0PAtWk+vBv+F3NNCwAUXjrW/b0aWw9ys2PJ2NwwakPI0hZ
PniOLvMIhs8brEgbp/C2IoH+U9rzhaaewtXDnHZJ6KwjDBODI5AtjLlPBzKK+67e
uEbimvu1Sk/OJxLj8rtboVbjULPCVGd7hou6BGyz5/nLaNQo5E9MZhlTcNQ2XWyQ
wZ0fnTI5iTdT+TBn8heTBNVa4sXR8dECFFSZc3sIoRWBmepROrRuGkk7WqLfFVzU
3E+0upVlGP5OJwBgF11U2i+8XyChRafC9MY8vRft213tqU4LJ+vipQFm9lfn4ASX
8fl1vK+tmtSN//J1DmA+BD4XBZzMmHObQMkCRvWKklvrBsm32Z2vHMLnxvBOzhnj
TsZInAmBjqxFwdwBhtEPA3OdF3Yg8mqHs5Uz4pPTv3xk0z7/CgAeewI1JOs5horR
EuB2fTiYiSEB0zpC6Ooz299347Vhp4hvTiRo7KlH8rCkRCi+ZkK1WwVCEfQzjOou
of6omAzLopsC1NxK5zBd0ufNlpdeN04puxk7qm3KkxOk+eG/ZhBfcmGo1d94vBoj
Vzv2HYBLlSv2xEiCR442CL1QD5FcXi7fRcK0P7jWdpPczsjTRyHPGGisSlwDVUuk
2yq8X9YXaaj+s0ENXMfq+qCA0QRGVVZPCRitCHapzE2oftHOFGwCDGEuPeneqREv
aXjVCIPn5xTekvX74sZ2sxEHM0K/HVSQR/uPTlKYxQOKkUR7B9/lXYPNZh+qEKjo
+F7Ob6SNsLKyORcyLF9OsGHoraT13xfzZiZcNccXWzFjKT1fbNLksiKWUybLkAwf
G9V3ZZQ/PCumvrord9AbuZlJo5LtQoEM7KgpSICRPkBwoe7puNO3SkrsZ4MNwG/S
NkteZtfx35H/Gj0CiEsjq2maMBC7+m3sLMAtNSDe7q+kVgWtfLxQAQUh/NA/juu0
Np9NANy9FR0VBJ9YRfsa9F6jReeJ47u5XeNiygN827mKJ4CFd4VY4iuD7gdNrWU+
2D0ndVn9AjxFgo86WFPcAc9fF62GV/nG6zyKKmYcXqqlrkgqVQ5cYnqEvx1Viodc
E+8yp+nCpuzT28kHX3qKT+cWh6tmtjxZ7Ve5zpkN6F7ODUBprgiQH6S0WvsYsTEf
hKV1YlfiPupHBL4QQUDdkzC2tG2I1iGiGLHgVNLG9dHPq0szJo3Aj2+zE7MbEsDG
aPMOcEmA9+8ynowk80cA3l0HEnP6PCVv284DZ2nEQGDNOTy2ZxMcX6VgN+ZlSqUF
5hMXiKnes6XcblcSBGKcuw1BiPxdbLM7OmJ1uTH1qAWw22vx4qVsbzmF3SqYxo7a
wmKrWrI1HetWgecpm0AbWxJVeF6EamnnKPptM79DioSaR4ECL/uvmW4622chRVXB
y2BVX8ItaNlT1M53a+cd8EesM8hsrkhFboe4iZs0M2ILLCUTc0LPxgEimP6qTP/W
NRvlcLLh2qmgcxxaE1+0m7yRUYf5kLz+GyNyy6WQJLX85FZjM7BumShfCAlLiY+w
6naQMXOckJ0jw2dtWPhO3H86kC5eW8r/nqWiG94K2X0JzgqElH84euztGukvx9oR
sa0737BzM9jI21GniAkFZvFeSDKJwIw7fYFrEOl1IdMl63FP7EQdVA+3izepegje
Sl5/zRwr1AYKhPS0meNfopvFZl0YjYeeWszS8efO/fdGL0+CZbj119TWP4YKIjW7
+n4jNICoQYqjQi2fLIxe9Q4RVW59gqmrmtrkj6fzsptgMk1sfrwjZSHzZakpILrx
qOfm1mL25S6y8Oy8mQ7XVYHf/e7+cFEpP0KbAL8PImmcxtgHR6PYjz5Q/58GAKzk
RJnxDUakV5ErYJgpMjJGerSdcoA1+gJeDd/9tBU/jEoQVp66hosMljVSIE31ffJI
hSxsPiQ0WQiBMhdDGhFpFfkffyshCgh/lLNeJCxUydOubVquyElH83wlDk7dHye7
Zy1U+gC+fpjOK8GvRpcHp0zvlMXGSmD1zEABnQffHLXRZ6qJEl41uBUcT/ncIcxf
DppUQKtbDoD74PfdiP+HdVPt17aAd4tffimmCmzqtgWhq7sHNk5XP5XFNDbNPnnM
jWJVhihO58QyHzNn4t8Tow68O0KA+eFIgGnYe/nRrs47h9wdzZJ65SOKQetBuvoK
0vHAA92S99DY8ySnpzXgiM38MnkyIwnCg1Fdlx9DsysvQGKqanvAGSKXwOTzz5Ih
NaaCz9o/2+rw2sAC2MdJDfKIxD267JNCW2wN98+kXU9vCGaFALoCcnDzMEx2MPrO
STTpzDgP2epoVRPXl8Atulvm6MIM4tJxjXlELlA6g8cvQelpN2UIUxegJTSPbQl5
OnY9XExbZfzYgncQVa9DqrMnTCAezugIpRB2vDo7DkCsW3jWodsfZjM2YWNwu+gW
A0suhiwKnszEnNk/mgYlLe4bhjjiaV7ApLIUxWM5ZWOxBTMrEWrgT5d6RKWrNCfh
P7kRH9JTjYdSoO+mJb6hpM1lXPmJHS3fBP+CVdbjCpQBpYsTiD0NpNKfLnuRA9tH
s70IgMw4zqNV6nxpst6DBIQ0wOCQbWOuUKSHZhD+FICYdMeYs7sqJFSOdtb8oL5h
pUWv088pLf1qSpMDH2JnoGP9X5WZP8Z+RsKErmmLaOdZurUZTyuw8DJhva+bBvJP
SL68XA6GtLn0tT1LyyOht8OHY0iMfUAt4g294iGG7C840RFmXAVVs3Psd2CN9HYb
FjXEvlH7rIJvaVA334jZeuRcMbtE0tCGhBP9RcDBiYVIE4r1kLJTC4yt1znUZk+G
du/Ibo2OoBT+05gus4yJMY4H02nxmC8Mne4R0qjBUlMENOKrnZar16Wko7gpwy/N
lQL53uQ5IzCGXSI1fSwCxk0l1+NBBd4jNIh5MQt8s0BdGhizIF+F1gSIZnHmPyhW
ulzliiNeEw24oDUNHr7RbvFqIS6IBqSiPUAXT+pcbE/G5fJ49IFAFng6DIPMBWYA
OCtLBuS1qvuDT0ZBWZBtwOOIv6bruKbknnuAOcIc2hCYc9Pi3+tYzFVkIKMfdaWt
+s3PloLXnn8LlJJNtrqy8Li68ucSBvPVWxm63tLk0O7Q3rB5T+sRCLFWsKKpZhlR
ZKn3T4CF1v1Lc5gYaA23ZXGIKVJCkvWfIg/MLR4+kcOgs3bBQb1jeDwozZt7bLuK
iA22tBMazUTrDB8Cx5a8cP55ZIJXR0AP2bDlcEC6UIK4DFqs5B5c5FU6+r3UFGZ5
prSo6YV3YOZHuFIBNIM1Jk7QL7Z9B6oyGB3V/aTjHknM8EW5mChp/E9c36V0EDRL
QXpABXXKqf4+2WAzbjU3sM6LhgC3A5kpVdFr1AFqbWZnYLx2ENM41BU9IJ7Y3gpF
Ev3PrwFDSjUwRVqj8oIqaypnvw8FedVRep9eIyHOA2HcR1AXS5xtE6Zo8ZgIWEwy
V3lG4U4UuVxpS9ULROTxeydh2i/mG4TslX8RUqC06ndHP4RX8C+GF0tjTALs+Ev9
dxreHwGJAdw/cVsgJG6nHSyLUbKy/mdvxsBpwhOgiof3bz0dxH24Yhy2G/z5VAxO
JGaLSU2R3HPAnEZTs6Y5mxUYrvNGRdMuGTcUoi1Tm8bGuIAhN66rjSjT2POyRvZX
AqtNzKI9RH5yV+qx0UzwFz7MvxiQiiaT122Rpmbj/PtGzbTIwx0GCdaWt2M+8RaU
vWy+UvUcGvAmrJlPHAGis7dcnVwdVXorb081MTlEavShjpf1trrRVBoKZ+DE9uwE
Ir5wP5J8/l+DGfed6eAoDWC7w9kPMaR3dvrvlm1u4ml8tPQYYFTENqOhRSFEFA5g
a6ytmqXe78PgtYveJazTvY0niod30LOL7SkBYWvqwfA8nx41I4CDp3beilR3PIjr
3nBP/fvN+Fexj6Yl69z9TMiGpd/gL42nk+6PO+EIYOrtmKK3nDpkqykip8vid1NZ
VRS2QJPDJQSs/eRcEOShYMU5EjyFmPTdTLY5NgkwSVHo936VkikNfU3k7u1tKtXc
ffp1nvWd8b0Y+ae97sJvyaUyn2ggQjLtW8Wa9wERoTGiJ3J7iusPncl/FiF9l72I
CM2QNFDFl6kXo5cpFufagcfnyoS+pdtB27xnqm5ONX/YpSy/xIQWm6fsE1b52gSJ
YXldxt1aVHszi5If2bI4T8au4oGIQegppcKEszGLr3wDAv0oEWqnUDAfLlryMk1v
dEQj7tqOTiLVXOVY3OVVZJjz7zC14Hwd3iZViCLXz6lrrlzjwABGV2j1W8giJr7i
Vwqxf+Gh7UuEFkNnDEMxaNxYWgEJZkW5siFURdAdcncDPzo6l00ULWdrRRmpG1aq
uYhmgHrPMtIN109s85aqQbSJOpL2gnahK4R+JyjmX5/vrg63EDzOLSl4digzhOth
w9DnROApuS2DQhOWllexGi7BhwHO7OuhQHQzQkMgCiJxhI7NBUcSybILaUOn666k
7wSSIb3psPz0B/QnPa9vlg3/de67LhBO5SAElwseSwRC7UN6vpySx/qFnWhvSAPS
u+CSH5KhrvqrGDA/8Ov4E74w5D8YfAOJ7YnqJzgDjevZMhb7A254fWyFut0gFCJP
HCRtYyJHEa44+bXcvobFeU3V6UqZvMpV3gS6wdSaslooumtun0VkDwaJbgrpUwCj
vm5BXtbBgORy/MrKMm11ABJX/WbShSgi4rZZw2FSco0LRRafPunRPkTSuwz+WztS
qiTap2/Eo2UhK4gzFcLEY8kDNmCL0YV96SUpW7DvEm6PTOIkD3QAOPdYLkR3Tbgj
hytY2BveNDbgK1mrj6CQ5MMjB4FPzYzyTDPk1nvOacu9/M8MVSZt+3ZqtBb+AItw
H6OWlA+aeYMIty8a7AxH0MaL6IjuiOJOvPn807PsmtHjBB5vZ4592RtcBlG1/qzY
QxZYKMvXq2QRt1v+fmIhGt518upl0UefaQNjrEHRh7GnsTz6aFI70JUW72keGV5Q
FDvzjBoP37JleawK8PtrDOoM7f/7BgVLFZgOoSDLNDEaUCBgstxUXVh070yKiVYo
4T7tC/tkzWnsIQwA20p6/exBUfAkaL+udvpbmpCT8cddoAwjo8sikSnGEyPX0nhF
a0EpsgiHo2WPYfDf1xR4CZmNLupXptWH1jqG4ERVsHfURAEgyx3pz7JgzmjcXEsK
kH4gOpkkuTRLP4Ho/vSIuVRjRWHmzBfIsqlGjVo+9hx2b6hTBvcp4gsK373GM0bk
L5A0D9PlW4QncYrc+bdPwnn3J9Vb2c0aeg+kzyPWxQp9eoy45FYy0LCVrSe2vBOD
fuAjcDF8Q8kA1sETTU5DfXRK3RgR5bQQgWmqkRfr6zFPMvcRkI6zUTl7LVEXlUSb
AY+hXbzieNrVTS3g01yDWbDPJvx2Tat0yHWEUT3r2j6fe/qWh5azFnZNrKqdK0sS
bwmUfWrlZGjDDGaNNyz8xb8KY2fnQ04WtUunmaHTJCYyElWmCC0ZKG8JG1GfEOoI
ODj3LS6Ce/RQ5Rlpi/Evfsug3uA4Kg/EOu52QJTDQaXHlXnmUCzKYqSgf3LmpdUl
Sw2ZR4Pd9RCcUM4d7JFZWM6Gmd8CkirWoCwb3VNSPDKD5RWcgVIFbJVeoa/UpC9x
daV4rxyFgwH6k3Gsc0oIie4wc+y4kizPktnWcHi9SMaHN8ti37UQ7oYRfLCHsO5/
Z5Zx+S5QdAj6xld9HdOZZ23jAgYE7uiSr4408qRDDgtMJOSvW+Fw04TNJh0r1tg6
JRh2FeOhrjkfSSBoXu2IgFuG3NRAy88TvoDhSKlsGiAp1PoFOh74GsdeL+gaqRGO
ATrGrAX2YZXjCwdIgw2sEDQobsxCFR/IovyL9r7tfKgajcVTz+m7zkPnL5Wp8HrY
zmqdqoLhZYLb8cplqpD/t9Rf/YBrbAyirqSQAqV1UHH5aX72KoCzyhjOsFmi+v2T
73m7LFFkAOjKZpOutgVNuJ6MLQsXmxoC/8ZNxLmnPbkC9Wu5TPWjXX9+HlKNKmut
jSAdkx+62oIZ0DnGnXJKx9QhXiKShQEUlCFNY+pMGxNEnltMtAxetUGBZ89Kr/vM
scoVjozizVpIw6zXSIHTurJTmFraq2TEl7Odl+Pbu0EthQdJ1/5bLu8PsOUJVQ85
eQksOyUpU69Ohm6gFIdxBudBovbrRgHzgSiI4NNayos7ZLJpBwxMVZZHXjUCgtv6
wbxh8ehgoB5/btpx3xBiwROPSndQKZ/Ixm8Ei6ZaH7Vy7sw6Jl6WlQZm2aFly9Gy
e/30IvXbVFB+6lzTAJNz7LPUtBQLHnjs/7fk7Vx6IT1Xc9wnxMG4bL9v7Y327sSv
RBxP2kG+HkooZ2sep/fshYQqK3Vr+uUbnfzc5e4F7MXuxdvCg1TVAbGypuy5p/oI
oRGllgl83JBTSVWGbtftFMOMEQYXFCtOvEjHpWpT8f55PcptOw7U4plGPAgGB9yN
97S9BLcAAhUecp4lwNsviA3bhtokD6EcEDliJOw7k/bacouOXOATbw5AAW3xTKjr
cnJ0LDw3s9Qa+hanGbBJFi2714YT96lqrTSfob1UXbmQ+DHleht5tMI1niNXBgQT
z96Y64QCieB18aX3HVLZ5R4GGbOE7tMJv+xfnE1P3F64jJFSjSvVKktKos+YWhgr
ZIwFEpgWRXjPUNy0eMJy6ftU8oR7pIFbwlgMh4Ko4U9S0zVUayOK2bJN0sa75Fl/
Xh0m5gczybHuvBv4wQkF40aDyN4NZn67ubQ91zCxvKiPyeX8npL8tJogMkgugbLX
uqCMvMv1brJ9fRAJeAiI9zjHC8AK+lvgack4Kbt+lGJvZirvTIV5V2XFc+fPl+7f
QwpMk3HViwUh9D3UVmKMLXLobGQs/ahLYWYjbqm+lheumGiyKXsKaW6QEyC8uyyU
lISbBUkn7h7lPk3UACI9ifH9exj7qckjTYbpCIPXN2ZsnedW+yJMakqh4aoYo6BI
uCgjQZonLpoFC3Bcq9zVtr+1ftIiom0B9mMMFSAqakxSB9TL8B4gZUrhcAw2kIek
kQznQzpHWQ+PC68emrPTpZBInvxDJIT1npd7jY0ayjZpoPHWsyrzhOlRqLoPVpii
XRv6MDCJK/gHimigud2iEWkj4Wh0uYtxFre7kN+BibyjlrCB99xfDBYitO1NpgL3
PKB+UsiufYcG9xsu+isLsrzbV1Hlf99fTbohI0zi8nIvfp/mglxA8+Z9CGcdY5ZL
arHH5VP3xRVZPbYua1XePPS0VoR/PAQXd/YZRksnoQxpUDz1jEz+Bpbn7rLzDdmY
u4+yQZ+tIewZiz9c9Xw0okpTz5iyIYMqu+fdfCmwT3+1uzYyR4D/+RuhtCNo2tLQ
bKJmtDQQq6XcX+ztU/UTkp/oZp/rYpm2Ylam3MlcTtK0XsG47ceXvqzMt2S6Nm59
sdOEuqcRbZ7FzqFEuBleFQ==
`pragma protect end_protected
