// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
QpjR/jffRR+g2StyjpqL3o6iU0G5Zne29fjQythot4n/duTcnpLY0aZTbIOA4XNuWheaXZFJxTkM
I6m5poAvq3X7RiOUsR9otUij51c6ksfGe1gJzb8UQhz5LJVE71ZpQbBmT7Pjvpput3ASMzdAr3Db
LHlLhcC+3zY69Cbupf3nazobrHC2hMzNxGro5fpUsyej9IrmbP/DaVp5J7QPf3pkniR/U2vKERl7
rlJUxyacjv6T8ZZXHz/dsrofIFIoNzJdsy8yLs6apcHk0DTYZ66gC5TQP2ELlK/umSb0OMPw9T9g
QBVyLMlhUUHTerir51n2ewPo5VCtmXduRCldLA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
W7yVjDDA9LvIfz3dSKWi0oiFMehoXPnKapoUVtp7LqmBnTPVriSsJTA267db8SmX0bI07+HSjb8u
YLiAB0DhAcGz/j9zckETm5NFI1nllUrVC8ujODJFRp5OnDPgCkOSm8HLSjvzQMzKudgdGzNfus2l
aen5egb0HFqSY1TKLtxb4VYJLlpPOHFiCo0aqyL2pAJCswqFX3PVQQsSjFTyX/XnL2hlTE+y9tAa
/G8H20Vaz/6AotT/Ig5QkbSNrULlNfZLxk9TzlDhokgyl8CV2HbFbfQ/WaDohgAf5D0sX61QuPDG
5t4CteiPmBlgbUTr5TWvBVW4spXqJtLpoRFXVEK5FZ93BHhSRwXTPufeFT0APzF4neIX5+t4mTi4
4B+wkFE5/p7ulPlfeJmJKeYWKCTYNh5E2G6IuVapIOq4ApOeqgKWAPQMCOkoUXfEb68mbHY9ommG
ALaW8Hj3+W5daSjRC5VtlH4H9M/GBll1Y5nGr/kyzsi1JRJFyohsOgdMP1lc0cHoO+t9xaCchEh9
cHg4KJgVxzzZF1Om468eRQ/kwB88c4YRdlv3WjppTWPPyPBL7xsjJRvDbpdMvEX3xdWtPi5TdBK9
OeDlVXcrZWLuiYbUbOnxqm/KP+Vo+qpljfg/mCE0JKKnfN68ODksPZYkablWBj9yC9T/+KGdNci8
Mmu0QAIfeuVtmuWPda19/PvbWuS+94gZ1eteL1qlUBbDxWAUKugOuS6jzX836mGpgaWTRuZYpwEg
S0mN1dxV+ql5ijebb47grYi/DvQBcYvzCAEUG7jBtIXog5NFbla42lqSaAvy66liaMIW/WgLx0Jw
lcAqo6/mUKw62k38LtzDuB1EJWS9QmcYj45RrFTULdkAVTJc+M/ESMnIJ3G3/cZwQocGqtiA8KmA
jSWD5oYXHkvQPHyRNtKBkXria5lLjrog5csgfSaFSQnYfUIDLWm7Ich+IdDPlrFnHa6+CAIuTm1y
c1pY/EOdIgb7Wv8hvD15RJgo+Xx++GRo0/DtrSEtpewqygFWCb/rSlO918x3e1OXdtjnkuZAraeJ
ifnEAgddFMFKElcFobFRWiJrFUToL+XRj7bNimTeqFZXg/AHaNL3WC9WlgwdbhWPqj/pivHLjZCm
Aip+153U5p3LL4cMmzvoUcfuZswqm9cBDyt9apCqKRGUHEx0IFQ5loayzALof3sdws8gyfJV9mqn
8roZVVcDaHcS/TMLwpzmUbQfavGUBTgkfp2oMA/rTBHtqIaqjAdku9MYfu0HhgEc5RowXKk3odnp
0/g3Uqjvl+ahDiHsec1Mx8ol7ysAencqmxlI2NiOy0A9Hc52LizMkHuxUuPg4oK2sJ4fvMCXKz5w
N6URfBs+7Q7VBkr31Nhpbv5qAK459Vtv/a7SlVPCgxU6cbxfesml8K06kifQ6R6QCYzui6Cqv/9s
fGjvqmlS9SJld+NfH6nhZAwOpELez0/6oQBYirMvkN6YihvCpZGiic6E1c3ARnxcpic9oPWNEThV
rtOABJTwfi/vk0We5qDHyeUSqKfu9bqU83AzoXVSKoVzYz533jz4MwxjSlkJV8p0ffPlShxj1mlD
fuDKZzlcwimnhJK2xUc+HTK7H/AFhb9oa8gwexWZ4e0ziYYVujk5OGp0DGA6tfoE6KNOPkXUD+yz
btqt8Gf3jqV1r2pmd7zIfoIK19pXg4kgVIo2I4BlRbc+wPB60MBGxOQwoyW1uXrzI4nWOXBXAVuh
zug3cOotuy2+gvXG4aCDEPkzdt7AgDkuviWhG45zfH34N9rhg3tHTrCDn+DMgVWhHbmIwhnE6Vpg
/8af9c+tRAtz62ByPFmVZ9Ow6UfBZHtbb95ey29an2IWiA+RkxXg+wmkbQsyt4pMhjQNTdons01e
eMiYHrAFzIyUb5ncW06mp2l9DU3fb6rTYy5JZQGF2fBOi+VYkBLETQThHDkvhimIuEFawplxLjyb
NT4c34i797LbKnCpN5QJgm4Zt4bGiBo/u/zQN38Za7SQujdJAoeuEnUhX65EcNzRLEdPClmR7yF7
mXcuXQQqUEG8OxaVwCY/ADWe7As4ijTy42ifgyc0NqMc05YuTvy7Hq4eCZQEGuYmaN7rcWhioHsb
nK+AQEAZUhTekNfaMHmXBI5M4OhpQ97H/rtNkbDb07MVXWMaIeghKONeC/o0vyB/tkbg4Bf1QIPu
Wkl579KoxAF2L4MIEX8V5Y8szwLAxipAT/SsUHIOU4pXkjZdj8CvS+vahjR2ZqSDZk+v0Qkrwm4n
s2MH5+DoeCxwiI6S5V/EFiQvk3rPhUliiAJ66kXW3qdqigVVO0ebN6V2C8qch538M8YbpyNC0cNh
SHn9dJ21p/k9mfiWhPnI/enruciQrFjLAW5Pw1+8FO+UTuKiu0gK9/uvB8ivUhgjwvEdF8CMKexb
VQPc/6VKx2+5iYfAAiLDNbWn2wxRrflFflAhKKfrzuX3nA9iuhR98KkfN6Wh+UCXxCdlAYlbf9zh
c7zMgc8IyDEqY26aG38OTUqtpMJBDMdn6icm1x7h5mIGEWIVYNhqzS2oirayd7skp0kUf3iTqnPn
K8YRrgbdo7Mp3GrwaF3BiSeI1sH+55IGdrORbBupNnrGBBlnOc75FTrQq2gSHuAsfDGkXZX+eSrZ
a8Bnen5lQwJHpnqWzSpU5ScUFTzFTrF29YwYTLzZ/ISwnS1qGhFkhwawqpoAwC9y3mNT1d2MXN2s
FoeNgeMbg/Q6XgZDdnaUPQxQAcQLFyeV4R72nSf6x2GH3lR5uFampGm/PXLMnXFtG0IPY1CrCl4F
W8lKR4ovWR9L/2NnFKoKylGuoVOboXUqUsIXx7xZB2b3rOCM2/5+BRgX3qrlG5nCtT12BMjEZyuF
fTn0NJEGp9m6M/X5VvSKHvYs4Wq8386a9+A6bv1t1Ruuvcz6EZugzSvAk/jZq/kA9acBNBPKcn26
cFkNOhhpGSIi5rrNs67nR13RsgFGKN6Fjgtw9Myr78ChOZ8K2l5MZ8nNRP1FkOy1/ETV4ocLzdMP
obn/vyohzn9jdX8FbA41e0kChU6sQcErydBoHFQCN+FpErQ59sIy9M0+/3W3AWAJzObXhlVQsAoW
85F4fzY82l3bRDXSCW4dRcRkHLeL0+uvS1sF0HOenLrWWnoV4BbAfxV1IYLMbkRuTAzoBCgECf7o
iLJrbMPv/0zxl9/9pIyDp2mvPgbVdesqo+3ug3IZyDPAwByCTCN9TdIqGlpl3owlNVjHNiWRP7R+
sgtjpDNLjPIemKrBxC6VPBxzpf9aikU/zO9Z9qHisg6KVP2vS1gxDmZt9keqdtFhVMeDbJf9iF0H
SKr8/djaCG+Zqc+lO29jc9Nn9HGqvrbhS8KwdxdYWXrL30CwT2Uy1Pp/FKcwPhwPZXbvZruDhiqs
S9Qd9MvWlEElCwZ8JmXq8P5/0O5X2kyxFYgp6y5Bvg12tFqey0qkG9Hk0PSacD7tHsqWGEUr1o0R
MLhO5JilaORiMz9gxp9tD8DwdMPTItlLOpEq39Lx5kV+eZlVM8gbMkC/UU3NgKAnWumbpAQNR3sw
JDaqvxYS55WDg33XCJojfX8cnzWt0/cgrdbsazblMaFde7HrLG0LoAOMUBlW+uhn+v1Egezlv4YR
RXnfI6IhzIftCMb/4+zZsChnXM07TYIiSlUDsNWUiZr7+BqEIFblLG6yJ1n/4cN1vFTfBm9RX+iI
GZ0gpFWe82xn16RMp+bYIX1vfnAJiRwZg7fCbk+U5B2ntBirB4o5bFpxBcA0wlF8MnMft/rYdweZ
M4+YqUuH9eIZ8sTppys6xrfbgxV8GBgP4BjZw9Ugt6rMwUkFbkBr0SilJfAxwXIPlLtLlQRQWFEr
oIkGCF5LycpuxdPQ8r4S6XB/yDkgm3v1BuxyyEzdHv2wCS/4EkcNFJh3WXcUeHMDzM3DKP7OXZv9
PHpC4jmNX5jYUcLmi7Zd24TtfPoogmftIMOhprt0jr6/NWrpcDiduCgLx+BrvzFP3xcPGu+spwJv
AMLP+OvDvQvMoO1WXvdc9lvQJ60Diq3ASL4oqR+bDg3PIWwzgwyoWuNvRccD3CbClYCogALzcEfh
OnWq7rgrMljB1UpSZ+GSI+XnAj9CwfUloeTUeQYFB5OrR1I/6tzUTG2XFWCoHQ7XK/lnUhLulxXi
fe/6OIUKFgMaKgrhkdN5bsJGsTT2dOhBTGZODSKBa/y3moODl6ATZOp8aa2bA1F9FW94V4r+TNaV
8OJyDoRvVf4f3lxncA9N881RiIzEw00oj/xj49qDsVsXRKkqUQB0lO0wWdv36dziYB6q4TLhbX0c
6TVsa3VXkfUiajSyqBakwcLFoAdjuB7unfvMwql6ekCBuaHM+OGAU9lkrENp6oj3xf7ewhJpT7pI
W1vj2/QPXuJsdFFBMDD2xVo/01o7N0HPGEhieIUiPnVwCkzFJ377tQAgM4wlYwmrFJ7D+UQBxLyS
kuRZKdfCVKKX0eFJc0erGS2ZN+4uoPzz8bvFNxYHqm/8mFhTUDXi2bFet6TCwMGNwu6HFRBb75Et
U8gQVUfX5NE+1Rwi68vlVlO4eSdURPquuBbeZEaje8zeHay727VPHIOIV/99SQwD/DPMFFl2KbW8
jqZC6Zvbb3EDBa8lZhePuR5AGuIMqaCUo+UKPp1olnDef3MR7t/HTpEUdGgVQtijHPDq2k7FRADk
+XggOR+BC45d9du+qCzifAOAptGmmJMFNsBBIz7b0FjGV5TpjtbPR2kiXqI9jbiHtloEGlfxknnM
NfsRMuE/xOoKuAPc6RuIetd6A/VOZkLm/xEJhSKwFtu9WRAJ+yDf5e9U3pLoGfKIx85vOcaEVCcc
JkWcZwbMTbWgUATBzwNFwQvh3ge41u2xlLP69Of0A0kB7WnSs4aXRn/JxcNp2txWI3yV+kqVupgu
uTYC5VN8qMbeyOCMjvNCHiwDujn//p0x3i+FYo4J0iFGUCgQwg1N1X/QFHSTsWpoAaiQEIqIF72p
yZoeTnb11aDjbnwpi+RuXUJXqCxR6523zyN/X9VIH2qyzuKR4aJd9u9mmR5CkXRd2Fl5GaATNr4v
dcUy+B+2jr6E9vKSve4Pd0S/gdJNgO4TDmDd80PhNeBr1fSp1XAnNx7Iyj3ENimP4P2L26m/oX5z
SQz4hX4pEVwMybU3i9UtyiIiSgtJA1agirFTCK7K6PDEEGyVw9tiEPGfVjL2Os3NCyZTk4xwUYJB
G3rH8fZuJo1dmXzjTcoc2kkDwI3yjspdJyeHRMwAfxmM4hmBHyFthU0vQho9BE9jnGNAaoayNiYy
d3DbIKKHaydlaFYlDpki234go3Z3aMWkFdcUOEOrYJBdo5JjZvUNrN0bIaPJWtSx+Wpv+Ti2jLdx
axSTBNhYt/I9p/Q9SCQp6jBcKGIPLF3vIknwU2OYof8DHGnHrUHIkyYMh6cvq7YDoyOrM5sQN8zY
hOyVi6O2+XLdK8S1WirPP6Qki5j+USJMGyF5BVLoU2LdSegV0nHRstBYMGrEGwKs7oiG33RAjbrk
3J5Zt4Idj+9GoRK+Ug4i3iD2opNPpS3+8+50P0j9r0P4aL0mXXUhC6dDye5i5wWxHapUZjOrOvDU
QdJpC3t+SsozLuM48FHwUFz4NM28m22ldsDNqj2133KPIWe59iGHBYhq5PXXnUbyldKeGUI7exKt
9STdrL5gefwcW2h0MzbM/vp1pbxOj2o30i0Y28KV+oE+TuZS6CuI+lXg1mmmfuDVm6nMBwSblBZZ
fZaIf8NM/iL6y8LlcT0jnToCZHUQF4TAM9uA8lmJi/Uz1vz7fgLT+BkTYKBd5MqxqR5r2paN2x8Y
mR7Vas52HlmWB1q75ejt+Rj0LLQw/E7HF4WDdJy278efE/6zfTEhskD6hdTQpdS9wiistCpggvbQ
pszCkwksNiQzJsLv+lE+zk90FRNb4VTq/EaMkfVwrE0Yw/4mDgLCp3eRQiUxPSuCutu0tMx+eTaM
qD1Bqqz880IWidQIYzItu/9dkveNm/vzQWC7BmNQLqD20vxEAKflkRDCz9H1ogf4de5dEBXQOIeq
q+484EPsq+jVY4eB8yqrCvsWc4FwDe0zdEixqNq3MdWCElfl5zuq6ivvAqXuD+aC5SHUQ+Tz8qJ+
i9UZayxxvIiFNVMRLXq1MGSEUQst+a2HWvYYBorUXQwaS8ewWzCCPDKlpoXF7Xnt5pMDLsiBUTXF
oy9o+Yvk2jRUhlKnXK71K/demSqpbhwviEIzlWGV/gefnY6s7vpHo931gOpEowz90u4RFamKqyZV
3EhqAt1IvEfhoDseecJpgwsL6BZ24HmIfU2xKz2p/88nhvkCDJqMZOTuR/yKB5GzAwl5qOgSlX8J
f7BRafE0rXDiyfUHSqPfcnaj6wWUyJze27y0WdcKvFUqNdj82uEEXam+1yPyivp0oLsV8cag+3q1
JcOUMsiB86ZdD8xmwAY84tjXgkuXJT9iW+SLrGWsbliiHS+pNfbWHIqpJbMm9TnT3YrihQy323Zj
9P3uIacY8SQM4pK9pWZCl1JtJ8peZ7nriFYj09BM2LadUEMJP6GLav2+ZLz92/ylU4S+xOw5o9yY
mDwgz2CzgHLwVUzgkLyh+zaqioxEvNB8vC54rTbcMdxAPwnsZI07bydZADiuw8XxIv6aJpNTVHpj
KQfSeHn5NhifiU0SpFwCVqJUskoEPGJRV93T7sW2c/nTIorFw6HExQii7iv8k0EWZWHRnV8jfqiz
w4640O2bWm5E/+e4h3wsSgbcevEcV3iYyvkBrMDAfCTVgIQF3xi+xjNsmaZEBBi9cKURMUrLg/HJ
DeLa7dAdsT+kOGdiRb6MWXJCxRzKAf52doVPV2js6jTFJbGSchJtl+yMLlQRIWVkjnHz2Qx0LwcJ
2muy6egNES3RUkJ3MiFSKahDnRbKN0ma34O5fyyfP9+FcVDyBBz8miCrAtb0bmtAvgHxl424IOgi
eBJ1T6Y/s0GreDuuDqeuNj72otSli3UQef0IuXmoTQvvtVfzkulJQPStYeGP79HF52ZD8DmFZQXq
FSOkeRzlo5RlvBvf7T4Efe+QB/aageuS0Bctx4w2jq71mGb27K9det7KjnNMeUkG3xgBgEZrNJkY
W5SmYTc43ruCN/sP04niUj6/bv8LIaMjI3AzeuuOP4QfUd+rf6a5Mh4mh3oZvqmnL6zswXIeSeMr
jyOxE/kUFdEnPOY8pXvCUM1xFSuPu5aWScqneDchrk1xlAIIOGZH0SHcBie/mx2pX2TA5K+uouvZ
jM7INNNy70PbxAX6pbjaXeKpfkDNdwexy2Ow3YbWLe3wbhCmBw2Sl3DmXEotQvcDA65hkg2dXhZk
1xVz+lj2SbVFtb+88gUMNXha1aaEsWlcKGChkzVp0aMkuxWsZWisgR6UWp5zqoEDn9RmnuCOPAw7
DNHbkcJzJlEW4+RgfYRX72rX2GsGBcfPXn4A616VsB4ZAPdxpbFvIgsNUzFG0eYEV6aPWZdrParh
rOY4ezrNdYroGxg3eZWIi5/lrp0hvEIpienXLIqDqgDizBGeZo5sFtU9du/b2MpN/7pgjGc9tt+U
l+v6Gt1CZphRyskUneXNd4wP62JtPFf43UT7t/RpSNWJi2CnRo9hYJMNV4DUF+9h1JrkmQiAZXWX
joEd7fQaAce8tljq1y/NjZMtGp/M1SW8G6svzFdnPK53tabzN7onThhON7shuPECf8QMX4IOhwtY
hkg7oJrnKZ4g3SlGh4r9c4hDX0mJO9RF312EXB8+jdtjQL7TeaIOjUYuPqKtJvJOVEuyAHNuWPXW
IQ2gkGIl+7THWenM8LH9UN9LB2qAKL/yVyzkA3f4OR97CBhsKElS0FrovHUHqxnmkf9hiiVasnjv
a0Bwh7/bLMV/onTWfpTOdq4uwD17+OI6k9LuyQbk0pnPtNdrnzlsO31svuMOs7m0/9o8NaHk6GsJ
SNCei5ubuErbJoAYuejxM6uRvzLQMCFAdON/p7BObRZdBIat3oWMv+fSAqt+qRUHhhJWggefHNv4
m8d0J544gmiFztCb/CRyYCePtbXu6TC0vCgAJCPU9NvYUTb1C6yTZzvhhirwOpPwAiDte3VDsJFo
3FGNv7F1YG7p41QFt8Rki9A6d4uFRgdR/WgItXiiUCgwgTsJFjI8TR7hNS/a7jM+GvUTpfH2R5Wk
IdnqT/+9zf8PZT/z8LoSFGfjM1e7ujw71k8UDEjKCB4o5cLXZuAq7YjHewS2C/ieNH+F2JuWSYs+
PKG1/bfuou5ZTwBLo+gPSX+isUXwJ7oBD3/p6wPZzhlukTQ/C6Lf/pZv5bPNLp7uyDCtea8ZUPrT
GICFbQFE7URDOSu39ZZe1iuSZhiheQ1HHTH1YVesSO/cbx8VSLfKHUDFLOBEzclfwiHvaxH29aXc
oJMBei7ZWEkMyacQhbOkL6ED6av+ZmlCvgwzirAq9yFdpecCof42LK+wvuT6F4usnw3PjdOQzska
XlgNG/Rzfrg5AkBCA0tVQUKoil+HZI9IT5cgECDQb63sH59BrxSi+kjzay3I/Xs41q121WVVl8V5
wDOgVhjKY8KuG2DO6+edWDzLcB/H5AkrklU2vLCwhQ1dJd5QbC9kLjsCxgIdyRZUNcGI5RnSoroc
+C68u+SroUOMwzehO9qjjbcqdrXFPiaf/Z8cXZJMzasq1SJE3AhmUXFQhOW7ADqF9IUd+9Ec/BO9
i4X4ryNCIW9WRmSSRYbcE4asB89kyWa96kB8RRDtZGJSMtQB+2fHJobHpzJ9Ee4E2E345TvkBDiR
VxcsGTcX+sF8ONtnCtiUDs5hfpJZbQV0JZ0sCS77kjprofVzWJnOffcv3suy2nSUnQBmlviUGgUs
a5YlrZuxd4lpC2dVeeBgxSgILESsOeNJPBMcoWDE6plClC8xA7IRAqqlf4F9jcDXeVdb6isCBv8u
KoLAdqBkoplYrdb3kKdZPaFy0N/6gqReRVXAfwA4BMC9ojASoePnRRhy6U0WW2xHJP/r0g1n0AMg
Vh60s1eqCmlXq3lfOr0udvGc15dqj9Zbm5No2u9TuKWx7eWGQ6ZsAcXzYoboINZb5RP3QMPiUM2F
Y+vjMZQLsFw52NTSeII5qqgkmIaHXxMg03xU29WoB1buwyqGa/H0E6l4uzCBUykNdcG4t5uKaIb2
BjM9R6+5AQC734lULAxKYMnRu3McSVDW7R2NPwCXfrVkLnr9rJswOKCiwlZv3TmLYutcP0uTixjO
cBupmGU7bNgiPqaUu678JDCY2adVBiorZxLP0sJ5YIa7u2c3EInFZaNpyT2FqfaqWcaxx7Wn6ony
VcFLuXgevU25cNCE1bUHeMlOF7zFrpipZPdPnkPXg+57HvjcSutXEqf72RQlp7OBtrYxHP2yZSxF
B0R4Easd/LiYcpU8JDbKMdUCmw33uaKyeu6+w7Tjxa1tpzSM5pE/2rX9tUjQ4cvWJ+D1MHOzf+V7
5fKKfCQdwbpCzkOD0TfT7fYRCk+htOiwqC2OJT71SnYUg+Km2h4kascNGZSzg85Fy9UbQCUe50Q/
tBwGvaMyMsX46ac489A0tNr7nEk+U+vfLpAafh8/qDn50QKniVgOP/NgI6Mtw+6WbmtxtmQCywZx
JUVeqoIEIyQy7/e/61vuAwOggKmANRKYBtmcA8j++iDWRh8hpTNGhW7eSdVgV0uC78PUkqwwcTcX
QEb+IuK0YFbdpusscTYEaoOIlmWoYlULeulQ3CrdkmiVosX/PLHKRJnEkeqp8VPXXT5ASzfOtD7Z
e++yVODrEJlgmC48IoHr5DqNTCl49jBt4j9vWSruZC0IuNiZFosCD23D7SV5PVqLCC1077DM/L7A
NvGQHjeZEuOGdUowkTZ8uiskG7xs59nvrikkcO93lkuurqnLUtuM/Ku60Ko2CWag4xIsimTMBagn
VnZpwYl5AXNwEeHh+uaIagw2HXheonQBZZoC2lk2hFrmHvDlqPOYzShcxZ/RTT3slPRzhymcv1YS
v8dhhHCfoqe55xtnPnuKs9e7ritqb000M/vuQ8b7OwUrpO/rwvv3MThqE6BEmZeZZScMdDAnjrOo
elOY4WdJcZvtMvQ0X2uIa2H94lMQacqfSu5xfDvVHp8GouwbrxzTvNlNjj4XoHB9SAoYnnOgT9Z/
LOGtswv9qU1i0noLAk3t2p6nd+IrRRsdNSFyJwKQWzcr6zjFDK7hrqs6kUoKVPPqfYpah+/GcDCi
2zq9+VXzvcvMHAYrMC+QOzUZchQTkI2PYNNnwvWHlbybHdZ8N0bXTEzOR7mk2GNwI6SwmlYT3o7t
lUHncmc6WsYjcz4Dr0pUKQmK7rJ4Y4bRF9tlz0TKqPH2WDLIEjiuZ5fytxpHO/a0d8P8xo29vGia
+Y7WdFJ1eba+yqJQTCMQhiVDxAuwVXrnK9RyAqYGe2g0sq3yE1SzFCn/ZnQs6l8eUoDXs/TPEW6D
YU9z0gwTVdDFukL0zWnOkWRB44GRHxpxmdbMXNcj9n21NF0W+DPGbW1MdbTfT1g9bHQNw2R/Yb3J
aWdBdKyX61W1iYpAiEGkDVqicXzalTNJFYs/JC/Rptj3uq9ShQfXzVkyCOxI1v7UYmD4rTD9t7N7
4GxGhETl86fcdIxxuOMk8dELA16ptxGQwHP6ZGAsaEYc2QDjOHjCY8jiUxHsOxfN2U7e8b5LSiLX
0GLH2ytr5hXh05V2dre0Sy6mCrzVLtnBuk8Uq9VfSJfZnh+XqOfqqQREf+4ixrD1a8AWNiuHXySq
bzBPGRtd5lRgf61XBNMiiyRoz85I9+3Iqr5wOR33Zg8yEGtalwhuUuIl+u1HRJFVPnN/gqvZRBGZ
syTFTiFJTpC7wpjakrrz9KdcJ2WGRdDd10ztQpHbiGQiP1K//EfMQ3PLCLXsr6HFiRMmP5k2ZhkC
uXc2StQxBfmM0iX5uhqG/oXLVQYOxUkq1+atjngeuzFPtbvoVcH2sTtwQRAbu00Myp5h36Nk0kOb
40SmEWTkA2ma4zGLa/XxB+oMURHDe4YArzlhwaA7gANRa7toeHoJXtp7rtLiEz8a/Z1dIaBgrUjI
7+8WOKPOL5DQvGvNur9CaASVaCmXlHXacdrEj478UP/f9zE8mqcaVzDIHEScRbsi3Dul3vbcp6I3
Q6r2kt7CvaIxm3bFQIZxrxwqL32s5lifF+PQjSCfqYY5KXJSSPeoPzCZ6E3FQkWHQ0Y7b+HRTUhv
IIk5XeQB+SNyFJjLcAzYZ3CfC0QNClYiF6Ch9W+E06WeC0d78Fj7WOmyCLfWO+vkPkQ6PGbmU0qh
pds6PvYZ6n4wjauMC5VmqiCSCza+y52BW8AAFHIAgamOffxPreVSlWubL84oclr43tpYtrqCmMRj
4KTxdCvZNQITyDlsXVU7F++H/+ueVDq76amIjG+b1Z6h0Tu59u769yqAEmgb6/chNVWbqrDVpSby
QbLinYRQu57fZtlohz2VwN4YDhD3vV7sDUTj+Ll9VoZn7lCdGfsslmKLjEtu416M7rEqBmXO6EC6
h8tcFI/URjZZuDayE5t4cYk6wRfcINxzfhGt5a9GK6V3QW5/Y7WKeY8gpb7oaG+mEgd74PGXbJ/a
cvaZ4gC4apFTJEHETm+WG1TV95yRxBpmstXAp+4ilpeHMCQMBOnuknVclp+3s86rS9ClND1vUptu
2Emk3Z/wuLCkWIHU1vdlEf3yJ3gk8RExYr1sRawGDz/fvNojfTL95P/kS+WCb62BIJr9wpb7M4Hs
UFaCy+Rz+Yjlxm6JSfoi1pfRag+XW+ng1giqlExhbwPX3TxAo3YV9eVjFERF8/wIBN+yoMvgEBMv
mb2U/oavb7FQbRKb0owCdt/derGizRk/JGHnROON4YlmCcYTCAcovaY6rXAPT2ffUacWNNUz0rrr
6h8LQNpOOTyVeYw+2DSfjnq5Onmw0v/pwbx2cguilvg/LT4QMcEBT8gL9s3h7rANX5aQG9+y1BbD
D+hSSJsAvi9bm5DnwY9bNCvGDXC3dRRl3yONbMQ4l2fvayOJgo6DUh6EBEuYCy54jtJq4WDOPQqZ
yN05soYcvHIabOVvNJdETzSWbjZ7Jp4eNepzABLR4negU8T2AlFRlk5VgKyxLZ6TeIW2dbOwRawR
4mPzc6VIgQhwLzENu99AFTLUPIvH9PGOZKMYJuTODpPPfQ6j8MMveM82MZuXmlzBcqehW0n4K2TQ
AuFIgieFq5JB90BsfWj7RZLW/9b+KfbzMy8WwJ6sQLZp6g1ooLjjLYwmvAZncBLDM4FsXBUfxO92
SmBYi5AWRmotfnu85m85JitSkHILwJ41m5d0KVyzmkUacs2jjb315tKbwvSSPu0xeMgNtO/IWsV1
RhzAyHfmlnNA6n1jCmx1cyNUYcWCLwy+3HjotjiqblYsTETncpoA3bCo9E/yLhNBzVJEm/sFQJes
20gx0hBhfA1puTZJ
`pragma protect end_protected
