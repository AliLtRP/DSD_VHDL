// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r8tlrIRTjNhFYmtzlVWSAQNPzyFXYCTZ+i/IfGeXo8DLVApcnwRXhzjUaDQhyQF2
Zsp6jls7S44ZPt2xmbtkmcg9nxVY8ntYU1atGo+aaIe3GUuAgwznaaeUBcsR+OqM
Y1xY+ptaLhLaZkTlStXKS+ccz3AN63WxaMXyq/gSNNk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3984)
RQZ4CK3VQNn0oq4RyHUyzF1+UaKn0qkLEI9NOVEdPIRCmc1Slywi69bHZUESYCkF
hXkCbjUIcCsdDojr1MC7x0SKL5U+np/G4o3zNTQIhqsawNtChELTTVWBqQTwvlxa
A7gMdaG91VnKLWf7GcjYCq5vNlsIqdLAckRjrZTd4HD2RVIp1ZHxhjcE2i5t0oph
byfKPV1V5jIdjAoiys6RPb4GunQrjJIJ4Nb8eOzjh8W5GY/iCUr2BU6gjLjZj4MP
jrQCKKoV2//Y681fiRfmsh/KK5ZGVRXlvD3AQgzDj1dC5kFRHTikHL6RGkrN+TWZ
8gYFovHWzf7I1ce6rQDT/1ufJSAw6GCdtGAvVlAP+CWLMFuGWYpSN+GtPGd3G2kJ
xSKP7zsNM00bi+GbqFH+0+Qh4aQEFqMbrIc3B/a8c41u+BUm2YbgAZuTRWHOZAYN
Qd7Gx6ZDMGsX+qo6XlFuFdbg34ogikQvZ5UfwIrHLoz2phZz9/US/WDhv7xmhSib
MYtvdSfMMVJat6z/5U8GN5VShbaEjOpLgwwkuXuJ1zB+zBbkwgGC3UxL6MvQXyG1
FEYbTp49lv/NWgt43D7AZdzXH+36MSJzXE79vXBkffxj6k5sxfm0Y6NhRjJhYoxZ
4mI/zfZTv7PhUcQX+mrKwrFRNoRG5Y8tsYop1Pr0avg/PyOvnQKMDggty5DSWwKd
SQts2ddAhxQFutu/bdnFuIx0IjZoLcxr8AiiOAKGZZoT9nHT/y2joffJn3KUHK2D
iydhFmShljc3vQnqZet0i0tuIKD08vkw+02jU6zXbnx9Jzmyhd+bb6I8HHdZwikB
NeE4L4rRwPe4VpoTkCJaGKkIh10AHT4yA9VfC5EZcSGL2c12DPq7meWRrt1xU/Kz
tC1JyQccIZdR58nOvc8qSmR4+86Xq3lpiB8MEYJFfpWyb0pZAps2h+j/2uKCyJ23
8Uh9ESVESFOEmsIBFNhKhvs/GQm6a1/OC/78JengLVeCDfBf8/hkB5/L8sV1H16i
SkLn/rSt/7iykZeU7rkAZoNT75tfhXRexZDhtuCKMCsLE/GRyXbZPybl2ojBBWTP
xCvXoN8ICpjRzhZ9coyjHi89YQRAPA6fP+qRiZ/t7so5JCw76CL0pV9AJ3SP5l7g
5Ru0ODA2qn3Wtu9g5dzkoCHmGapBVXiX3EkoHqWLUOc7balIPBdYeQ0MzapVhsAr
O5agBxAS3Q2PJaDZ7v97GwM8OdQjEXMAQZUMxjig31aXrE3LmuWptA+rvrLsoz5z
xPFDN502G680le7udpE1kn6ABDAnKSBkx1J7IyPv1ARVpHprhyvn+hX6xpE4nC6M
mTvdHym92u454SRFNhIFvoBI0cpiT1I8mry009BPSe1/tMr80JiPeVmOpr+GZ6Op
XcdxFzOzCjeykn7tEDD3Wj8Hg1JzyRFjRpYQKgUm+wwonWkHVPIatGNzh119lDbQ
njWdGfDUxZD8tFz5nhfV68R9cNZi/VJR3ckAsCwp6P04pqoO/i5eDpaWxMaCPrMI
1/4zsa0eqyJL8SO9RVzU3WwVd/ZMee8XjyF4J3zBgKGMbMMfSpiVNqgkwdfRz/vQ
SebFMCuzjl/UYh2EEjkQW4boul9OupTA6kSMPv9MTBdXTa1pE7XVH2jUuI5LDMwl
wSlCKiIxBB8Gl4/5kdqK2cU8pUQzPSp6s4OeyJfjcqXyaHcDkidpj0WbS900Ix89
kZ3ljrkLO667QPGq7URxbJBTp7fCRDKeQuKZC4A0pN6niKkGkwJR8Bv1m8eNZOaB
oWDM7xLwQyGysYAu5FJh1CnLUTmkDck8YECVU09PjBOModyo6Lmqfwco6oXb8/Wc
OB8zYgsPlwbCkpkiFlmyUWdd+hlJNtgztfKaZLZk0w+G/EFnEdhExCkpfB5AcpM+
6DllZGYcC252BpekVquSo2bCrgqOA9q9JvaOBtVkMKxaI9ZJCDJLG8zq9SrhGGsr
ZHWKWqzhpWFhJjUVBfiOT5j8F0Vc8Dl9UzrQlx4jz/7ictndbEIusa0T8voWgWCg
Rev4LcErHZuON/XZbYRcyjJjG2Ub/04IlSIN0Mv/9Gu8xu4rp9UYidC71XkNVKIL
/PmbaNMFH3GxLrzRgVEEbtuhw7jAuZtIHeFPgVgXeK6A9tYkGJsdxOK2SCgn62si
sfpjckEXI5NgGK6M0ne1yGLvS/MQyGFwS8/cTsiesY2ZkoCcm+ZtV1Ez1pXzoHQj
/NRJF+esJ3UxPkzZylG/LEAUKyp16Jy/8kZtKqPL7+wbVQbluBVaYFz8HGH9a7q5
atqpB8yf0FgKVcoNvENCarYKa36A5430rBeBGPn8M+7dk0zl48Dr8QIhtaLs5qq8
FdEWq0ryhHZqIWphn0g0ld4A1+fhvNPAUNjVIvlGbIYGKOcDlDo1ZcwH2SquPo7Q
LqEfGPsGzEjJiIcQjxHoR4ENyrvOuIXAACZseyvbV8V0Rz6yNnf/41QzAf5qN8p0
6BFK0Q/f3C792UDU5+pNlf3LBDKaYUNLz3NPEqq6sjnWryOlAWLawYv4oQr2NH6v
nWLbHoV0mTWdLs05aPr9timbVrCh3FJRORxvi/IAAGfUwxt+wRAUkGTkop4/07f4
i4USTo+tRtSZlNGpgRWG3aInlodNEM3BMwjj/qzLrOp3Su5vXuQHToss99DJstpP
wl/LG+COcmNC+Ybch58ikrFdtwuisvHka43wmQHYKnD3YSWAZj3A9UcX2ue8B5Q9
RK8RK1S14n57PAmmScHRhyX3gcEWGAI9ycxGC2mSU8uQFbh5sw08LTx4WBIKNFMy
T1zq+Xov2HZijRqaiNQG8LBwq3YCWUaimzGVdWpJ8dxjwGKio9APINCN6nkk8Wzl
YN2ZlW8l+2tdB3MGC3u6es9365GleVkK5PuQw54Bacs7eT90D+439sV4yuKf2UT8
PmINZxAZErU6LFpBgK0ME8zX/kKkpfZXjTtfJis8AqM5hI3KPaUmUXqCvi5DmB4n
n1l+lq1+1QMxzyQyjTAfc8POu+Afe2DZvjSS3ontAvkiCmDd2gYk+VavNIuH3qS1
Y2n2MBRml+EjtvgW0AogKNp5c2t9pXSaD87P6GJaSAhPWGOxsCvmnWBvfGymJ0G6
qDl+HiXT8ln/kskRX1osMFkfAyWdKahW86/Q6xcIyC4y0zL5G5puV5NVGfiVQoXf
PHcn5FkppQ+VFRUhr9O6CUbl3T0nz5RPXZoAQZURghOBlrCoGQVurF5g+NLuEhiz
2IfAeX0vYXDvGA3jHuM+22mo6UkRpU+nF9iJxntDpyuhqOmLch6dTbpKfeoX+ZHR
0ME8cH+fSdX08YVF2rlkRWFT7t+G+Tm57kgZLcQ9r6LnnYuU1ELnZ0zRMX6ftARq
VuHpUgnYhLxKNqBN5MN8nfXGyhmFw+9zf3toQeSBDMrSeWzso6fBzD/gmkH6zXTd
VUUYcaZReOTwjpmSQwjrodnI3FxpfBoTLAb+3z4i9Mv1B01QuiUQOOBQ9HpSl3MF
5Yp33fdeBXwdDNFEMjO6PjV+8NeErinD5NKVAqnG/45ck3bjqmPxdKZY8NoNI2AJ
uTLv1jiO1MwqWO7MXnR5R4iMy5scvLmgmTUUZ452T9jAnRuWusk08DgE7J9kbZT6
nP7XHKA7PKj2+lghp8Tzut8T5sdXeX5IBb0IgptCbToNf8blYRNK8h/Rb1ftXk+w
upvy49pqH4fJi9MsiCVSCpAxD/vBgkrU1410ZUU7te3DnpPrE4j2PfrBFMmEbPUx
ivKPf1F8DWKqBmvH4FuBJXec+3BJQSsOLemfawpcQhtixaMCpfdnKsBTVecyginq
J/jsEMV5S5VtUzgekneZWTJR9ZqvxrPjVO+/tCSG4/IYSGwKV1UvpiP40XJwYd3K
I+4MPfNIXt9EytBoA70lOxH66F1tOAhSdEz8pgnDZpqYFmPMTn4aA+AHm1+3gCEo
RfJ2LF+Jur8ew9l6gk5HXGBfqwqGyh12odds6Ig6EcJbySPuOjcEkHXuXhry0b5T
eacNalgCdeAvfJZul8jndyJMlO9RbL4kPTKlQPWZqKndYnwa04yV+XlpjsecLyal
xHYZxUUMDuRWl+r2A1Hjup043u6pK0RgKzOb2Ad2k4AWfBQ/icTGarDQkunc5AAm
bgLJVkghc0Np4elD4NGBeiIN74JqeamWYumNPehKaiJ1iAxbTofj81oDtkKFMsLO
vQ8ca91N4x7xMO4xCginOwqvDCo6JIKPZyf+1JOaTi7QeDLgPyqsNLQ8fCRFZ9yg
8AnOg5cSU16FNy208v8xn3tpzX4/zwFR7ubOdMJsu7nSPSqoq55WyjNEKz95S33F
Ls3eYB/SeGE4ooHwIyUqKfUiLoCfXfMlW+ARgtRulHxbgFrK/SZfxsRdq7mHwT8B
yFwHp5f0OUfE3dysU6G8ut/p7nKhcUPW2v2eA8dz7pH6HeFGhRvglBDJTMYjVw0P
4zC0utJHU8Y6gY+2hl/zbVFcV60rIHH4cbI/SDKo1uTkuWzmiw/x/+3viNooRRVJ
BbaqCWHV9CGra6cSiR3F4FdjCuyBaU3DuXBnH10IfngVSinO0gXEnfrASVnAOIiX
Vs4RetgEOF7N+Fv1ofqj3IjiEVwp1sqg04ENvxxuGDFFcuNWKTAVIBYEw7blK4PL
foGAW9HH+oab42ii8+TyvWdvaD79cfE4+p/KiActDqdSkasdoW6gxkbiAnIEMhP5
ORzdPc2FjiBrDWNgUflq5d0IkUtQJ5f1hxep8VHAzVsLHN+MgxK50n4uI0kPhTmo
hCE9QQ0hSJduogyeFiPTVJYrCnAXzK4AYpHJkXLskc1L72moUETxm1K2VJDzouQy
npQICGvvxeSY0wkd3EslPIYzUstHJ6iuaEaa7r6zna4PeOJvxRm2Y+BTT1xNxtAB
eT3TjmOOT1wP4wzDeweKBkvS1LK5dcQ2wEKIq7JUj3Gq7lP6vqjsb8F1Ha0sMJI9
gjkohhFS0ymSAzLyFoXN6jdPqjf8X4VfpMsCQ2/RzTyJRXXTBxTqM6RPIRho8zL6
Sc3qlzUHrbu2XnerrvQ1fE2ZW2KnF/2sOMMQzQBd3ZGxyL7w6YqQv3Y3dNHt+D02
Zel6l/IW77EOrhaZSytD3yni2tf8rT6b8I+hwQxtflvXcr6K8xQi42t5uui4JIQ2
kK3wuPc6uKZfp9SCHFRqkSiz8IQYc7Y5qBWawcvZcAi4kFCemc7fCooyyDzQHR+0
JBCE/QzqxpCBP9Pi87DkjjYj9Agc1pkNxYlvDCia+k2dKgdDT/TcRHTz5Fddxg+I
`pragma protect end_protected
