// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cZPnKenBlx5vy7j4g/DHCEepeUvR7U1WzWKvimpz6eoWHZCKu2elW1uUHCXZfRoI
D0DXj1nG4Pj7FcxGQVH27o6guwowQzFji+RLZaBDDoa26zCnsgteijUPhgnNHlTD
GrSjwK0NB+/pqBPh+dThdgCYyUNMbvb9G8K2qksZsqM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61984)
KDmG8jEQlEtLHN8jiOVr/20NEbMGSdNnVBqG0QGsal7XnmGXxb/j3VH0XSoqTOLB
dqinMHosis2FKGlxzf+SPGcJIguTCPYWTOYf5wd7soOMpri9bHo6lHb8ryR0+dS9
+GGD4sc8ICoHJfz5tqoRwuaheslXgKM2fERQeEs1sRhmQiC2Ix09EJNbQnD44VTH
FGgD++XCQ9/AdCaI50Mru3YJB+lmpsLcNTlJu6isJaQBZhzWYpp7WyquNhRQDlhz
3k1l53b4mn8/DX3kH1sy01tnXZs0Ml/L5mTClcTzdGBVPd+/YgCYTstXq18LguZr
51X0rQ3ODtixwFAwy07sKhPrqpv009pAtMIaEaTsEfGmEApqef21xIf+/niWx6vc
WgxnRn5vWFoaGqMvXA9SdlriV0LI0gZXme47SjCSYuhsnViiL1rEfQOEGZyDrzR4
Q+1lXcF4H3OQkfUku4XzMT29VYJrb81cDSM/1Pejr+DtA5auf3RUtvxWvJCekrwb
3Hcu6+JS8DPJ9vFghtOKmbs8PlYfI5Y4V26OJAi33Yrs9vnBFp8Zu7909YQ/WeaA
IO7B8AwoF6RFjf3/NolIDy5D8mVK125mVt2LqOBJEguDdSo7U4orr0kwHEY5+j7K
N35Cg6LgoSw91BkHoRz0a/fysYiTlDXe26GOEBIlkQUB4A+UR4CulJZ3sCKADq2M
M1ChhZuBBWLtSeGEWqSvyrnUBwW+Lp+O3OzgLvDwVDy9pNsIfN5o7DOL+omF9qea
giYwqdJVg4gkT/SW99j1Wic52yBaa6myrxZW3amsFgdTsOS4whqFybKJAtlbHzi2
qrVPCIXg7zRJ9UJJ5IAhBpSDhBj1ir8Y3BRmzYWeApXYdKkVk1foQw4nm70OvrNN
ty6Eql0YLXN6c6kZLotAyPQfoWmkmqMCsVLjAbMeSsGGx0mJpVzfB5FmW3dC0ctc
929yLqfP5onduHGjAg9a407lj38hJ37dMeWKkamM9ICEfugQTakU+T/8T+wvQ+DM
3HCabYm07kQCVLruK87D/wsoAokcRb6rH9t48q3cWt2JSFWQimBS9t8Dy9G21ciq
6sZHQQDtrsvlcYYuAvEvXf91OXPV0pHHMVLQ3fJ5oC56EdMq6RGoCC+UPpMdg1I4
DxietemH8ZRVX621kGSF47K4UhC3J9twINIY3R5oVKoFJgvd0HHJKefUfmTpp0fX
YwBSjQjJ3j6itx6s2DKApgtDWtfe3vyZ+pGY2NZUBXrOS1xkIVIWMihq7dT/k73Y
VMTr+WWj58OihKTQHihVeQyGJUi6XDVQ5tN7G+ymeW1Daol7XOGn/WWzuR4mTy2W
dcQObS2gMKLdTrBXJtC01+l0v3dVZ8sltasfrvprK++cTDzOgPdKPYCmMdAgmgaG
VrTkiN7PA1NARjZTR1aUyqBUX8o6esWMHGZObcKhaLiZOjvB4YhXl757aan9ph9T
B8wR399A8W/ISQ58FIu3vpJhN+TkThvOM0aVwp4JwADGGMEeeq8yUjykC6L0qbo1
72tZj4HHC3P4lUlpAQT0nBFW6CHP8le22cjlGQVldA2/KKV1PiLe4wS+rFUzpbj5
yc0mZAMZCXys0gOOSEAcMjBSk//cDTsb0cKGZPaLmRBfmQ51uMg/rjZoAacak9Pk
5nVoYHIO/W3WOH/jehdi5Z0wGLnRLsZjpq0UvNc8Asnz7fLBv/dlE9YBuCZ5hZNy
JCeKPJq29M12M2EHhl+XcT1lZTPCkqd3vk4i2jMjVWPGSBv0kBQQHmfbwik/DgYI
53WgN+c4JdhjQBv4UEYVafzwipXCihfIMlMqtUUCqG+4hCb8WfiyyCg0XltyxpIW
rlMtflpLg/LEcWDea5ZGK/K/g51SSuL5/ZjKEwfdDDyEAE7NVi2WdRArrf7m1jup
8puHNJBZA2xFRfKhj864elYSmlpyAzym6+4+o8iY3jg/eYjaRogBxtphY2opDfoV
nqVzEckTW4odr3wMtiXbAhza2tE+HQNF/0c2Nb+4l4uTGnFCP0lm2qfhx5fWpJTd
8nnLF6peSAB0zjQ3rtJFunJu/nlQZmIWBoaV4XcE+k2xuny5AaJCjo291eWQPDVl
SHD7tduaoEpW/KhEha72nmYS2YJ/+ojP9CqALgM3uDH/85W7RFDzVlV6MoeEvjuz
1hClB+mT36s4B/x/Y+q6NjDCnqvG6oBWpv7qBv+Xj5JXILpkHWfdvn0F6tdzl8Gf
LNE0W332pRmNzsb2QTBriMLSymNeRflGBdCntzisEGodsUgeVBbjPRXIRuYrGlL1
O4apbOsseo2zZGam8xrnbCqeQ6L1FG0oXm+EBDIDMKYl6Hfsv8oC+uy2SL3vYdrP
PWiCVmh/Lukp69IkmTVJYr3fUkoH2n0d9/gRYw6X4B/cWUaSzka6bx+wB7zCSCFk
avfzQFIpbUDnu7cyoUZi7ung/CeTYxlOQCA/Z7UB3W9WR8VDJyUCyxEKjQszGFIJ
x4j/vOa4T5b8E1YB8kFV/8Kpz+a1QDX3Ni6Ol+AgLOeQ/GKfQWtLJ2rhfIrLWXnp
p2ZMQonlaokh8BjWMyGI6dCbeVM4zBotjVl+frTyPGt0G29nw/Y+zToIJKmtbFRD
VoJ6CS0JpbY+x92lzgmcL9x+6OSz03sE/uDujKsc45OEcvfPZ7CKQ3hNn5fC5+AE
SmoRUuCNIyCJe+FiVZ3ZQC3iOzV8UAZWmRgBdnbjX1s7wO/IW0kuDonQcPP4moNO
5qm6gZb8DJL+/IWFJ5D9xommhgd7CBoT27D+i5wevPYy/pw2iel6aA3pD4aN9ajA
oW5szDyFKkufTRA8D4CMD+Acm2leQiZal6jBEGQ0JLY73igBYLfmwMzmIcCveDcj
Xdhde5alqVPN7abcMTniNZp5mLMfpo40p5VEByF1Tm4CKBMlAFHX9VAfjpDU05aD
R2bt7Ly2pfqLQXpfNlPjPlSUZYuyiaXIpKfHYLhhvVSCV2aD/0y4OAO9F+1doVNP
S0cpr509xWHzw8BD+ut20tcOelzSGcTTDp65Ex6dE+gAmD5/XVj0l3e1n2QyUMTw
tycGlZgeIAbZk/Y8Kyy+3vPz/NTSJP4HS9GxMTKn5IoFh9hIoefEQyxZ6GBzI1EJ
2nrMKQdApdYaUG4wa6TjuXOuLCkrzXOjyZ3wxEzw9oS4aLMkKhju2IMGB2MPVtrU
DHiNZ2hTeSBJ4n5gnQvItyAnbAs6QKH0GpRT4amEB/GV4LAqSatDzGr6kNTml55C
eHIqncPFxAVfVKkWWpVrQFcciR4ttBylZxy7lztMCPGZuKwzmox5q7kQWPOw49Nl
HcqYlhakkp0KpRKEa2s/P+9ctdutt72mzx2GdX8zH7W1FXvCtYk0wI4xSNSfswRq
EQhLP+cL/vdtF1ju04GhLcVXFJuVHfAFMk8sSrd1YB7WDt5gQqVtdt7FofZks7n2
JSlNqm67Q/6zn2Z33aYbJGsBETRtu2AdGEOL44hf3yVHc/Suk+7SINOQoHpTP6iG
YfPlyS0ZXWS7f23zneAdcaHpNiaFbn/mZAYGI6gTSd8PaMfE0Y3K/ZIpKmOuRf+E
bQUXzw++4rBKJp0iC3UPPcKWvemaNJgh9+itHH6xePlCk2dYa2NW+H/r8ggEZuPJ
0gF8ZZPC9fRa6uoTnYfgutFj49CNUbtrJFZ3sdj1GxfFWfgTRTSnFlcR/JRW6Oee
YiqTF3a4ItFonh+EUNzauVy759bJTP9LbBZkU7J7g6Vh+ZiUlRAasfx+Wv/CkXK+
jeLx+mZTzEuQ6+7/Cce1SO72McFa1btPhxiBnyO4OQa9hyn9IM35yxg5VtCeQSVM
eHgk76k/g1Fx4UCIFk4AwPWsFSp+cRtk23Yvb7IgNhHEojalLtu+qvQB982uta9c
SjgkM4C6TFjKRpCZjDE/7xMjbP3awDgkgl0IXaW1yWJv+K9nwmuQDVr2sGlPmppC
uooBsi2I6B4EQWko05GQQGl06Sx7qLJ51cVk15tNfpwMgi7+mBgyDKEA/Jtd0j8o
o//xC+90rzdJwwDbELqgenfG3YkEkm2zqUa9VZsaPsz0SR3ZJHRsqpIqp5ygHsdW
iyrmWISGgr+eO6uVZZw9QbQdVrsPLRj3IDNQIY1YG21KAO8nD8Ok9yHHc6sjO+CQ
r+AjfL/mzGX8k0slP87htBIBxc/Qh50D5meZRIoPAPJ58TsDvA/iCF80yq3ifDW8
RTK88cbGIv84KvZ3J/Ws8gUH8f6HSpZXnzeRk9dOczXTIyZ0uLPLklUPXa6GmwTE
od3jPdjqSRBD+1CCk4Z+9njGkygvqVEB9qNg8WQhenBM2ZWqB2h6AGDOD7I3LQtB
BmXm2wYS5y0I30Idk9r8sVo5eyoMMgMQ399DGUoEBKuYxN2jiOKCKfmFyN/MTHXs
Ted64meootp0Sl+t6U5gMqwgTAdxeBdjZ+zj7BO4AnQNYQiGbVjjo0nXY2B6eb7k
c2zzWqIQYJxCno1zFC0OMcsfGPFOSSyf7YaWcmjQoAAH9tMEcc1z6MpFU2YnoiRn
njorXzV4T/S4mFbSGLMOVpG6nyGUR3qxYuhvuQFinyEiLtKqjxSGD0PKxvgARWoO
4u2Vt0LIAF1dlIdfnh2aWmQyCNSLmZH1dI+BIPOI8zGNtozuw2NllAuSMsrjTknT
gfNU4msK6+uQFRfj4qj2AnWwR6DqeJBMsjZ2CraZ/B4w0cy8oV/MyaRTkX9T5Dbu
bYuhI4W6It+MRKYusTVFrn+b0UMJPxBpvnktJpGfb0j05g6KLBTf1V+nVlSVV+Zx
mQDSpGnOfOSLW0WEwjtGQvrwhjEb4YSgS/9sph5bOMkDztdjYwBwWh8EtUBdT4uz
/k9wEa5K7NB++6S1fUhnSZS17etl2Wflh23+wdCgmODIibc0mocf+osL7Hvf6lxr
rkaoh9aHM7GekXYxHbmmvYKz4rHkA1CaBsV+mwlbDWrsFSHSSHbJdYpNb9512nvZ
d01B7Bi4JHBS5knOTD2PJ32k9eUEq5XI1NI87nh4ZDHgxxR02sQmoqetJ/FpnBa+
PcCDj5HKeI8QkduGuSAprzoFGxnnI6WgD597n7Gq7VxUpdV778VPjpJu6/v6LnUa
l0FwxUMY2ITrG0f52l9T4QeVIefoOEUVIaJIIRJxZnvGZTmXJhTe3PtDSCWuxNhk
QR8WALF/FRByM6ffmmVq1gCyaQeHU6OhyrgOE/6qLxhLaPyjThsqpHW3wnAib9/t
iT+VUkNfQaApfl944nELKm+uVa0D/sZIM0hM+R9pzOalvrUG8BRI9ZWzvpTa1ouD
RFKNg+QPw6kRLsu6puRnLP1wmrrSgg13aY3mHhK6jZ1CRrrHsvZZ+rXR/5TMuim6
KgTHetI9Ggpvnu1xX/fU+Tl0IrJDYwbYIPxGwU+azHBWUaQarhFBtZeekFekLHN5
GKBIL2ecv/eoQ9Bxu/I35xjZut+JTr1wjG7QREkyu0FVsfOlCWfeWLCm8JyCY1e2
FKfOd8nO5BDVhgkuhATveZqic3LwnnjVkBpLsW7AYglmKCfB4fJSNLK0Xt64Ybb9
t4xvK8Uq2iJJCtWIH4KDxYQDnKdJhXeNy7dayvsz245Mlq/yS9e607c/AweB+AL+
CCewZqjJAPFQ2rkefAtZp2ofKF+LVTns0U90J8bQwBlPFW5UeXAqQTBTEGpOtdBN
8VGGfCmIhrsSXenecwrjwu7qtyOnDuhO53K+tmPpl81NUur5HLABsJuzdLJkD/jk
4qEzPbjNJylDPZKPZJv4BicZyLfFU70oU5PVHCGgNw30vU62lYxTYl31EnXMAxx0
BLhRTLpBoYf1/dDYyL6Bf7LXChDIax6MktlQQTwVAe0SFLBq8CBxWgfWZYy4iFn2
6DwbZA3XZ+66TQd7vyPg18ALGqh34eC0w4z44eU/DgGFaC32feCy7Skt8X7qKbw9
Rw9PxvKZr1E90rTMAghZaR5QNJ3uulIAwcZ0Tp+5pPRjoHpwZEi2OimUhBOHNoPM
3WQN2Bo+OX/OoYe7RnZodb3mYlXvsWYHBlX6lzGnf+su/DDp9abbpNYh7RADP43G
sNH3jmDyqJoi42+JncaO6Yu33SVZjM8wKkS6W+LhqQhDv1NsScP7j/5EOT+OJ8in
e8D+oaEvf+V9R15qhqGnnSIO+vKOPrEcdQhTRr0Rv2VytDmFZBhhZlVsvflFaf/z
uMaRk0Dl8/qoBdEckFWy8TrZ2Wg8tzCiOq3Du3I/GVUxxJP6rFFaTvmw/s0K135z
UVR8qr9xtlovMmmqO21zr7c7fqJO/BgU6xLJIAg5lvaR8CegXrnXANK9pRbjuEle
J3zVClszH/dbzSiLqC3/VHuppB1t6ekNIbSzfSuL72fxCQ9oe+eDVSbr6++B1gHG
e2ctvf7BL3zY8SScZn4/Sy1x+9t8Y2eyRInH4W1h7TWM0BwOZIyzVuThkZ+sVy6e
KcNI8zdYXINIe/X6GzNMORHaGJOWfu6c+gFj27pLVmkDxajGdFvgntMctS0j1yp+
YB311UldEK2CHDZqzA5qPs5FuRpa7Igl+6TFY01jT+QylggVVpijxgw70P7KwSLP
koF5Dhna+bOxlj57yH06bXahhEkIkwnWdyYKbnEdEcBY1wHe6WQAACPZLbp0fuTJ
DeCqA+/wNRpUnp5h7dogG+e82ItupdWiwlC1t4aC+6sKqNMksWDIB+o8+IWcoOyl
2z6fvw/c+V+t75YQXSJ6WWuyaDBdjARiE4I5hKyo9TlybQJvMhjVo+moRCUshOfD
JuepXegT7mVus8fKtzBdx94MR57qcQMpoJ0/EsGPMpws0oKviwhub8z4D5r3wK/I
QGjrUnw6jMz4NVcen/Bp8mOA/wKv+YqN2SJBq2GJVqeJJUoKs71m9BDqaLSZeceX
P2c6e07M3e1eAtF2XhrQFyP4iOBQ4S4JfQ7CyB9TzsSY+oN3ErRxaUig6M9sDj4/
nlrN5McFGXSWMv4g5Y3YD5omvQGJhKpDDEtjNM6Jf0c7prrw97Dhi+A1fZWax8LL
OEDznTmPSnC3I5kx5mrytZInai0pwfY0RlAPsN9kgCbdmJ5nNSBJZ0KZTHvxTW5o
0f1VXfN/3LKDy69iZ6Qp8KIHmKL3mafxGN/4x03tfFAbBYiuDYi81UhqVsF+LU7m
A8YZKdqBeWlluj5JZPpyO30h+e2eqtS8g5hC7EQ44Si6RqzR8FqhDt6uZi3j+qoi
7+MAaLSxF2Q1eX85AiToVmUVihS9tFWgqz1E08VQUlgKcoN2ruExJDiJad+JedKp
etyPMdVeS8WLkgXxwBNIonUi78WeoYTstoBPg1XlDBlLetU9SrWd0pXDcvzNP3H6
hL9M94cweX0Ot+fieFcukFPPM0ayIWSH+45nUJGe1pa/7/I8p46ieFtyDJ7qe8AN
A8ljw4ATm4AZ8rTbqpZpfoN5PeZWNXW0BFDxMQZqEUGfVf+x4pOBRBV48IJGoIeb
K9ZNc5f983Wr6Uqroql1uN71Cj1HNakJug117Y4NnvjpuGJRjtn9weosLmMv752n
73HpEuL0kvO3vu5oJbK4cwx2ocWlyChuAwfYkIkWu5fZmylpF9g5c7jYF1O4HbE7
Fv32hLJKcqaAPFc/rjz/vPiwvn9TBp6qrjpab4ui84gPyaDOuK+WzkEs2pmEziVS
Szs7uyUaksd15h3UnXiuuD7QflkAS6+LZlueWED08NLWgQz8KOBm4zIs6uL2WggZ
qQcZpn7NRVqc+J65YLP0MX7SiNE/KIV9YBnHezm3aqqn955JPIf+FK7s2yFnFD4V
7BuBNonzRUsDXEgZDomfTmYFWRrPHv1NkqQbyTKOS2YepSBnUTXarxvjzszE2cnf
MuuV6trnWYzwWUhG9X36/B+zB/nkvQCYaF4NkSljoaPVpYPVQ+Tbtgnitiw7Lt9D
o6YzA/JeNyE7a6Fyq1kgZ9N7emghu3oIeId5KpU0esoNvrU+YrLg0MC9gz4s5jVD
JJAbLhDX1uPxDYabEB/zHzG84cDjT/yqpw+gn8gQGdejuDv1/CUYcAUMXcogZcEn
5YuphL3toe8ZqC5WIwEE2+hRX9W/I3gUi0/uV6rVixksOQA648DHXJ3CLJJJcpeM
boTG1MnT0pGZnR+5rC4GxxMASZuMUYzaTc7o5i2wI595YtL8PeR7aDCM8H6zPEtp
84MgAA3Q/V12dOrPBWANVBvuFyGpNG6wUT5h9IWYTTAvq6FY495b2ITb+zNNrn4l
K5OUVoKfDEjntYY0EmVkj/emqu/xQUC5BbG9mFrt57G1ot4+5PVSU4NUKlsqSE9q
KUsQTYg5z9tpa7031LNu42SkD37bhI3M/l60zdDmcWd6uheEEWZwukqSFo9psuBg
OT0N2bow4hScczOn6vdZFNS2fTJgq2BJQHpArcPmiz+OXR/jquw5gxB9enL21ipQ
cPipl7rn4pe6rCYPymiCwnpKkAjCvgUgv6/zA5B/2amKCbcmYWXcWf9I2cHsEA9m
qcwgu2UBKYB1Q2GNWDYDajkQHrcIe2jNFofZNLz06SALabaP91XZ1On1sQulNx34
teckl8JtnGXH2Zo4VA9LfVeOsJe81zq3BpKSVvYOoeVK18K2HvBhMlyfe9kIrCg5
TqpfakcyawcrDnaL2qoP/rabedGFM8RTzito1blSd0GTmTT20ns8p1jhviGV1n9f
P94OXGCWmHWWYtzbeEdSnRTxuNWQbh2Gf3z5KXD7jgey+kyKTraZGJC4NEpiuV9X
e7KrqZxLRYon0O+qgCGi711ypkZBP+F3ZVX8sEQNFfhrXB0ON+JDGEccbY/715+J
qE1G1lnH1yCrBw+sw4XbUlEhi5yV88wEKVkJDmBEvZIiIrr4740Mub3lgRKvtmMr
vqryot3tf0TQKwiqHKHnUGaKKpdTRLK8eulF21uAzQAXTWsO/EqL1UPjQ6gvogkS
+N7j09Snwdh1ZBnTKQKr69nSkAHRMH/Lt4Dl9tkyXoiyGUWUbbDfh4mhlFfLHadL
G+R/iGmVVOIX98H9SObIBgVciHsq2Pd0QhzHxRBYFyD08T7fvt3eS1m8kNl6guiM
2efl4lx5n0telTj8p3js7VUPZo1Bj8sCsw8efjeVbmVr/nYu9gzRuxj39ujXaB4w
9u98wZtkhbOkutD0zVefmRaCTBlHHyRJ0zAn6pucT9UKJ+0BYyMH6Rf1tncH5EUy
usLTspc8QuwB4YVyi2jqFp0rGfd+j5qgs4C4ncgPQT281PPSYs9gGq+Q+0Jv06Hw
QScuQHDfiVF/ApzGcmXxy5yCn3rhd/IRxhE5r25W5MBvGyLEHqQ99afLmifeiHwp
x8Ch30CVnYdEd6vpUmMfxYOR1ym17pcXSJsBkPUT5qgOuNsyFlDucktyrbJdJMW7
0M96/s5vOcj5Qu1LxC85Cc9RIei8VW4SFHeP8kIDVLe2G5r/qyAv/2VF7dzAjToO
ivyjSJWfl7ZmwWkRyP7jbIWGLOsfFHrNWpkDrQw28WVM8BLwSwa33Zn+uB2FWqGf
DJQ3jrMkYgEaOae/jEYJItxA8V/Sia5QG0uyEd2CN3jZqvn1ZroDCg6mBYY6yiGZ
Y0zANHXC696gy4D6XeusEoiU8CIIdzlM9ku5K0tkqgQKjvTUMmCL8LBAqoVvpDr2
HU0BX6OCyuYL/rjpvBpFdKVo8HnuOaQ5JT9rVkL+ow4KAPKUQr6xYCmGkWpyqitq
JWRWp75bSG8dqFE3uZBzd2EmPZpCiQR9l3kzXKTu4oFRpp9U9U+7kq/gyr/kGc76
gOy13Je/OXLiFvmvJp5TBpfbDyHlQXEUpVoiZxiyVNvDfqp9EdB8tQyO4BaOyoSa
C2aASe2U6Vx/89MMan9FAS1skkyDvGW06vJurMZCuPSWInGIl981oShp6R8CDHVh
wwux1KFcitpg26CSYkRmJjQb1UToEuvh5CTWba8BCdzdyCHDwzRbuLvQrpajsYMI
VHzbfu4c2hnqKq3FfwO2U1Z/lynLo9cpkKowyTsQoSQtI1hrAlm+ntn8GO/ZK+7w
JmYNLf+04rsKF3Eq/fNxOVQXDc4a2vkmHEF13aIbuwXi29RCVsV0tVGOiLmDIZ21
BYAAXWUlscvjp9R0r/t/4HMbbraMdxKs/gKJlYccs6xqZABHSHql1ojLuh6+0lm+
UUZHBZSF9O9z0MTiQe1gNC+p5p/Lur6Xyl6VDeFQKvSPaQSujU+LWpW9Gc0wNiPP
gY8sLr740qQ2nFiKsIw2pLPTmY3bPhujEWwPtNygU1AeDrkEOFTtg9LVtN59/Hcf
J6GrNmbaqK8QtP9qz+ZAZKrmoeth8HflSTho9eK1K9svOeBHfvKinWqrEUMbGPi5
xRXJ8bQs3/DHghvjxK1Sdlhpl9+jPPRKZQv4dKZtTMz4o6kF2g677RLZ0KAGFNHp
P79xg+8eGqIaNlLrZ+A7H9V6lwaLHgnD/0vR4zHzgWR3+IldKVdyUBrqYo/iLx4j
nDMsrjr03cB7DazhSNgwE5Uk2uQZOH4ybv6Ks8v/yuQ5nQe/BbohvOHcfKs3Hz73
SwRMlm1YqVQsBpKzTtOYwwj/3ntyrSDNIwKVA6TXMWHQW7k8qTI/PHIlqfYA3S9z
oyPiEnaC3U/pAXXsjtrw0Dcr6rukg1wFmBhnfXBAG5n2LVKbNGzuozxF0roDZLjS
SJGH6k3I+qLPjxKgH0ZCVqbFoVz29F1g73LjCiWqSeJLFXrLxGqL14pCPGYL1aOu
Pxx0lguKxk5JUZEiKivALPiSDBRBH6qtC8KbBkvp/8r61F93F3GsJNyqWHjonvkl
WzoSOCd7j6wbHNgPAfYmVIYtKrxhz/Z7VpO3ydnRTUwEdrHIoduLiHB6UDXL+jnX
WfzEmB4CRiDoVY9KGSfv2tEk/0WvsLKVDiFtdFuoz7zwSkxsKKY6QYCHtIdB+hSm
Osash56X1nWka39Gg7xott0VE3fpZ1tT+GPw5CQMeIxRee5oy/fYMdj/PlHdirr5
vdzRnJhBj7tWw0+rIkt3Of3c80snIpZx3Fke58rvtU2kjDjGEVHtT3PYQoTqMajb
dwpyhWQbiO9onczu+iPIxFAdqTEwLYpBUHP+lp06F2/I9+6D1A+U+QoM96eHcABj
BToDl6wCb9/YStxPWD6N12454+nMWvMex0gqTeKz220ArQVZ6XoMMmHbqsGdQ5rT
9y0G8jucZHE45JVytDgb7xmC/nZ3OYZ0OUbBJLn11hclXTvJd/2u5KwXqxUuosqX
+lX1LYZCYpJ3cWsvADcL8RxZJyq/ZaVF9y+zuC/wDhrXUbEdBQiLDqBhx6xcrDzj
mYc+BsAUxBCeC1FuJVRm62KWPxFd8Uw0v6zTkoLggHUS1g6JoepKv2pzEwJ3Lrrd
1kM6wvcwVwraHJcOM4vy8IxCtebgb5oqhB8k8+xrlt3z/hncEXNxPqn3nOQ36v5t
9PawS0O2jqC98llLjwwWunOG0YthX5q434y7xT5bExfeGvtnXb9bsumHG2j41Ct/
1/mQ0vuVMM4gKDv3CiNHQEgit/2z3i4572HVpi0mZ6vIgpHe8rM1HjqGMguY1Yn6
ZNdKV6w1ZsFyTQJQbvSfjaJ3hkI87Fr0+4Kb8x9eC8UhB1WZrjTRE+R/tBjSWYOD
GNpr1zUyLPHeLxvDa9JApK+oWMytSdYkKvWCnS37YmF4BR5CDABUKSv1M7k08sGY
JKK936nmiZ4VO/SfRzZ5oR7pHb90wxyKLzFYh9gGAhr0YGx78oFNCasRTj+zC9l2
ItFSTg0K/xoZagr6NO5QxcYjwV6ARrK17629KDpx6XF5UYwzC2163UbH520zWi6e
OBUCX2iLUPhfjXPjn5gP/M+xzXqaIaf6+UFdebMCEREMus9o4QK5HRriPTpBj2r3
I2BZRY3aEbGD6l/8FqIxuaIkNqlUpSv+/S14D7C1biLNjOAYvc4kCRsrVBDCzTM6
4f5Duz0MJcogkGo/FuRWyousCDqxSmFx/lvJjks3hSpDI+d5Guuul9juwsvqmIBY
4fYY/ZQskDBHpN1vH4+rFCOUm7Rbm1aXn8+dVfCPBjoS5g9CfTs/fchhKFoGNH/z
lXHQjTjoZbJGBbmMovr0MyAtBWxXtfsiSJIwJIORDb7gSc6Vf0vRC93Hw4Mg1eSC
VZjwX3g1ctx1/xae+v5GEC6Vmje04+/s++y0xXDbVf40u8owtRDLpKiYnkOtN95C
NW/SX6Teo1tUSE1oYvPQ7p5KIjV3RRnN9z0TQCvTX7ooPJeLA4JiPYYKQeWbcD71
JI579rwpyrPsP1bcYydpGASqNarZhapVazSq9mSTG1vJh168CHbNmSb04C5mRupS
kxu8zeOG9w3h7eV9UwiDdzAZIvUIFrEV+mBXotj19k733jFBzUwdkNZT0KDct7/t
8C6pPq368g9hisvKYjEURS2XsbHzLnpfhZ+iifqwSrv7+rDWSh4HQywMOvFGFcLp
NByhhMoh/fn2kQmTWap87DzJXLiJhjxc7wGinUcx3RkDAIvMIZITh/88RYWFlXN/
TB0vVGDfDXg8orqJxWQrJMy4aIvuQziaIdzynDzsO6mpqFr6nDAR8R6EJtehIoj5
OiVkTbnkaT05mEH3AlDW/+4lqU3ZiKztaW54TyhGfrov0Eq9g/LAZNiWSqCa+nGe
bSG3K4MFztflEL5ZEpjgfaOSIzeOqWNYeWRKngHoiTgor1p2jAeUwciWdtm9m9sg
WaC6vRggPtaFv/JQ6X5ESasKuPLCVpk8tEifbBptN+E40dX0NRUEIiwz19AJzFFV
AlQb4o/Xs/uW6xSw5wNgrE9QTKsvTafGV50svPK92FNN5HQNSNw48JA+k+UutsVN
iw/IjtvqqOFAxENhhCO5ZWhKwBqnUElyaQ1GPEBncF1j7yoAH4YSdQvyjVj46GdY
jHejR6O/xTkzIGjYCXyPg5vPet56IvTlA56TLpi4fFR0aWB3WvroAFmCtCrQrLCu
4n1RQApu9JfB32m2VLWFuGnLBUe8WB6SYwCjnMv8KAtRIto7vTY90XAhkEBdcLwx
1PKcCudblWF/yxfE4MmXzlYFg4k4LYoy+e1dQgsCcM4czP99ejxVHi+v7/yXyYVx
YbZD0Pi9KiKY5WOSIo+pnq61wLx3eKCb7HnaRRgkqi8gy0NMnZbUVQ59Aq/Wu9tM
yQlB6q0GRNRft0Fskbl+LcCI4GNaaAGZpNKQ50L+3wl839sUJqVrQUiN/GQRpto4
xSDa7rMcbdk7LARSosMXBTXqbO3FE8O07sefd0NAuIRfPeIYMHcYeNh8yLtPZHZ7
aittmFdzDsE8kTHU3V2vRDM0i68u5iZZMsv0hHO53GwuhCDiYJsUgr5Mc6Wlqiuo
PhaWCfnrvLz/7ikYD4ZVewP+6vbTjLHF6GjtMwW3SmcHvpgfvFLSDJGUBvl4pCvF
/4JLs7vUi74y/7oYxmkWmFVlIp2kc1L5Jk3/4BxwutIUJoyCNF4/xx3RsuD2gv1G
Z1aVWYnjWNc9DtDpls+nEDJc/hwWUmJF0GbWWUswT02QiLrYVfeMGRhMfYBA6aS9
LNy87Rv5SXg5pNv39MEWYYdnD/WWFco8lp2OM/JU/IjRUsZYBPxTDew5U+tb4Qxx
TLQ4sCG89fnEKRZ4geE4YW9mAQrgPhnbgsYFr2WrQ/PDmCIQBpy7VEbmIm7lPwop
V2uXaQO+ooOvWKbTFoRB5128vpvH5jScAHZabYyWj44DnqxuEJhr92/E7keD/+Lq
gUIhY3jtmQ+e6DyB3fUCoZ1xzIKcD/erkNQB7uP1W4mbTce06fAYcmnc5L53A+Pj
DM69UiKMK8qwXbHRnvvKklIHue/jixmCnoO4Pn1TrId6E3sA2JtIVQKteXkwJGjq
9B6KJHBICjPXG+pwgrweqmYdqDW5DLgxgtTIrhlHxbgqan9R5h9h+GZZygHm0jYP
cmsQWQniV77FO9bp3Bn6XRHJMDmzaukyvTF8YEKJfnr7ojM73VXXTj47zJKx8qtg
2qjwZXARbUU3SjyOVdbriMTdbvpzkaRnLMrAW4YX3t4Qxqyuwqg2uZsZnxps3yCV
3xwz3J6e62LbcwfTYckFCtOfIY8KWL4kHrgI4jnGqG0x8+JjaMHZSTZm7OoT3sYR
UiTC+I+ADFg/k4yv/if8lrcTYMcLwRluiDKj1YJQ7abedldEiz+OmmINPSoavKa/
tNHgewfaoPy8lVr643X3KEmEANqlZqDK0ZGKr7ZkXPPaF62rTVDm42haIR1PNLVv
LGarRMiVPSfDkRvX6HIOv2zkzM9zENKSKufZ8u7EazVOJ0kGD+JyivoLKAwUDf0n
9jpTAI2SKYxOduuJ7op/Wf0h1scNNiHYCUonLsDuGmf9ntX34bV914cuSH8RGiJh
IGi2nMUjmdJvlPYx3QiqLwyzlP6CMppVy1o5U4puUuEBwaQXxufNd7a7WCw08UJk
Pihat1tjHpZ4mLh1g6+ftUTeVD8faYErBwEx2tfAoLbClUUsx+d8OG19lqy9lLtE
khf0cJnZFTVqR9sXs97JYa5Au0OIfm3BIKdd9MxMCZY/QSyxxT55g5rAGditvl3Q
xfOMsCv5NpN0QpK1nD7lvTG5Z9seFNx3BzPCtrowWdfcN77zfpYLL5oFcIscbnuY
gKAOjoPd87YLvcdwIXdNLVmftDOR2eiaE+EQEmjDiWrtuEHV+Gzd8fMZAGGRvhUx
0S04A/RpZCV0czr6dsvbR7Hv2o7T6nIGxQ7WMwlnD3vffdfF2CinIZUD3a3/Hwhm
qhbC8Q2suZnOQ+8IYifNQ0ax0xKCwCh5OGz1vo3UjsB8mu3vCVw+ju05kIetCdb8
sn2AVqspEhWTanCpBhZg0O5uLwmuHluiemkjK1XzG25KgnJnsLetG51F4Y/xq0qS
0x+Mwt4dOiVybgLk2J17BIUy363gDYYRHUpDoQOWRva8+TGLGwmDolcmAWUtrr0k
NEQ70MhvbnJBOuNpHp65hV72anfU3mufVc/UhUyRd78l66N9sp1bi261v8IeYwvV
U5QuHwLmrvrXm5panMZK8LbLlbCa/kdoFaPQ0UzX1VtS4qKIsUx+2+CS474neePl
kRXKu4ZZC6eTCNTOAxfRG496tdjU7+ifLCO4ekcdhd3cTwu5VAVMSzXLEzUajtHV
sBosx2o9CwL+9bWJC2t/HKMZSpf5KTRwGGqZ0V4tW+1aDiEhC5ZwBueokGb/Gyfq
7sc5PN083sJtLPREI3tiAKavLtHUCMOeLilFhFPgNJjjpvf//0keOcqihqZzrxHG
/Gu/RE+qE+OlCE3vV4uiL6Y+HQJDjom+n1F/zWGp5N3Q/kv7Du+1/1xpdOHWKHQK
vD8siD9KLfFBtdE+3eN/GIZoPNKWtuq9s/eA8U8Nw3mXtBBM83R5CDEhXL0rtbDv
hPxNRMNcgX1pzcU6q+QpLYI3AY+BXBjfNALHbJ6OgFcOh3HqwMOMn0CDrhwFo56j
fanjuHVW9FlLEQ1MGAEDKq2FFG0twUajlb2PDdfLXH7cC0rhUGRUQMV8DrSeFPq1
tTEsW2C+NTLu99mBLN74zZgc9/2qDaRAzw5Y1MdO2Cn55DBhvQyZprVG7SvVWZGy
G6q+ZnV4e9sPMIxkcwD9XzXloTN8s9d/IId+Ln3vsGpLZwY/U+TNMzRtz9Sot+kJ
3iyNL5pTnTnLRjcgTxSFJ7NTfWHWaWwhU0TwAlLtzbyUhQfvtr+MiZ4LFXuusbcT
8XkUd/zqDpDar5sD3FC8iOBEl6efGaDjUgHolX5aALuOZ4qDuCAv6L12PXYwldBQ
Mgocut+KCCCOuqWOLg1g/VUCjdT2p8ivtxDf6uCws2fhRdm5+6AuXtbl8fOzSCq6
JVFb7dxTkPSRbCw0mrbbpOItsRUtxZ5sLooi1k6f+K7IE/NuTbedkqrf2i8nQoka
Y/FzMqdeTf67ao4F5B71wILC5XdD3rOUqw2v6apiuBu/jnSMK5ahif+hBSSKpRPB
cDFrJv3GdW/Oyc3I3VYBRhBZ8015v2iMEhNteUfpXQMvo95DPc43RpVdLsaO/YeE
INxq9p/pwQEVCyilLrXX0S6rEvIWkKvvrJqe2bpCLs2MSEfbv1FvCZIcbTl21VKG
/ZFUguyVp2mdX3rAlXXEc8ACVoiene1I4aHfc9UVXRI5oN9WKswwJ6Y2g7BMs+oa
1DCCjulC5eH75/bjFhNc8EuupoL5u1b7y28u4JzM36hECmzgd2fhwaLIHLBkr9JK
q9mON6AfOvFCUw9lPJshEaRst1vzs9MYWb1GiMfo2nyfj6ZxBychu/+JucMkFl71
EbQQfzzPyIx2i42OMwt3dyNvCdiAr5EDItbQFEba3z8ZQJe8+C2rXrasJXN+kwsJ
Qft2iQkfxB2YoxgC4/K+XzOKjFLVrEyG2jBDpmk2B2VGIMEU5/hbHDm0g2ADcyce
W/XFtwKO68G2JAUsd8lejiE2aR6oCCONlHLyqQeFv9QAHbnXn9Evew+5A07Yz/zD
oGllCsQQHuW84i3trc97RUE9D5oyDvUT5lMZ4QMSEBugf+9S+A6MXJvnVWlJpovv
4jhnt2//fpnneh1+nlxFZ8z01GcaJ6I5MTjxdMMZC4892kv6g3bCqZlM9N45I1nh
1UiLfg5Ru9oIkyodnuySWW78o1dPUIHKOhTqbWYTzaOxPT3bldfiEl8Nzsm3Bnan
ou+H5jXiZO0c9qOet7IE0qy4CvqN2uL0HSMx4AalZ72aCkVjayqpZMveVTvh1HEM
aorIZ52mjNGtTqWhw1RDCPtZ7BJOXvDZ2yEMp88Mg+NuYtSAwqCztr7eG9s2eTWQ
Z56eb+TPlbSvW5vwX+iba2wsdoAVCqP7AU3Q/XcDiyz2q3hFhI9wWvVrtPZxSXa2
Slwo2fWa2apLy61JTBwvFXIpyGLsMMWskfIfXPFK/Fp3QkLP2dvhjHE68k8rqurj
6a9FrtSDcsxnfesdkkVv87tPnDtH/XvdC9I/Lars5m5248uclIN0rh/b5JI7AcOA
XfSGuwAyFHbY3o4Dl829MbNznI7cFpkCtjfVVclH7ORpIjsQvQEnAQV94hSNCEur
UYeNljZ9d/G1UYEParaRYFjonF00Ikt/T8djx+RwkT+Z7w0fbhI3f9o551V1+hLr
MSUI074qq023x9+nSiQ8vjkwuvfvWDEaGvmHTdtFzK7RowCNMBigSeZ9vp1g9OxU
YFWm046T544xvxvP3GxfHlahD5YTIuhDtDdx+myxY7xHhq2Cg6WGEe9cJvwjBPk4
pd0rn4foPGbGt9biHXILPaatvnj/BMxWgN9V2UYy75Qtth9Nss6bnevzwknLgDt/
mFXdoyZYJ55ooEapD8AR8wlzkb57iyClZJf6Lo51N/P5MYLg9I4MWBHJ72N8KHBe
Bu1vMVVpkk7EHW2BqEaX43LH5er5Hum2sukczgHdATTvcLOGeWZL5UhSjQLl2TNR
pl1Hcz2+WTVA6wMYdGmK2LTP7p2Xl6kMjhQbNEFOESdbxTI7uIa3W7217vQHe84U
8xkQStZIVyWKHMDukXjFUlPSFyDIuWYMhh+2hvW5xoTJgJz25x2jjh7Yvwt5gWOO
9XwPvSs2nEUsWlvsyN6hot7GG6GnkuXhGTo53omE5Q/W/IzgbbAQNtSrWyxyyt/W
wAqfDLqra0PMHPi4WtKtXrIatPEZHxLiQNqoWreRNUDdwYhPT4MYT6p+1cmOvlAH
8dOjtNRcecx8NZQAXHy5z65+0MOnTXJRbDXCBJz/nbHOK/zC+jbNIg4ljFeOzlYz
cG8U5O1beeryYBD5MumYObU/08mo1GViASq/vxse1Q++a85KGByDIp5LZBsT2xw7
g0B0Ap9PDXPOxAogAexX7AtC23rsnPXVhJrDqw/3DcXTSgeyJhur6fg30N/u3l0X
sSfbQis6+4pr/Xlu6jv/Q9m6tr+kEpTLD6w6tIWnapv4aVVqRrWD3os1ZYXPHwGX
LImahpqKHY9f7aL15umWp3ozz0Cfxq2oySD70PYXDAkOYlxgFTY+biLIu8+/0PxE
0fYZdSGEHVxb3Xod/OJW6qxKut1N6UAUB3XBwIZ3AFrstRqdqSmU2v2x7HCCnH+g
I8LX8iP8c5qtVqqLy82CKcg2TqonWT/y6os5qF0cqFLo5gvhGy+IedBjiPKpAYav
s+KZli3hEtwZ+q7GUBLl05eZ0E1Q4nANL+VHoqTc20heVrs3zC8l3b2dCJuLW0M4
tn+8y8GoQPKekJeSGo+AF7zJiwjKTpz9lyxEnOKtD0EuJQpBP7UrgyVBYXlquIdi
FiWMjN2sqlcNDK38zrjkJtbRrlewco5eY6OKdF+sFTVYoUwRx0QqRhyzpNbxOa5t
Z1rHvCUb6j4OQndH0/e4vleQf0Z4tq2CWDnq5CyhG4LHs90HWtOmVy0UKAccBb7V
sA+iz6LbQjXrq+oQmmvCfQSGWsHtl65iOE8CcvKfkC9jQiKtdwoUU7uCXIZDeSvI
HtjEnHVVLu0brD8ZSx5EVcPrUsB+8WlVtJIbS/Hsb75ocQQ7kxCkhLGb1gJMEmJ+
pAqsyGKdYEYmaEZGEVkhLaS47fYT9PcEJ5w8AP8FXXBiBZ46IyGtO4d9fEKHyAxO
uc1Dzjp3DjGGfiMYUpgRDM2khfciStG7Q/BUzUOYtyLG9kObBXSK4IQC4BS2YR15
bAk+ju2FJwaw6xU9mwXQ0DKJSRIdG41jdmIHUfFid+2gAyLbCp/6uB0nALbkdZwM
Db5VEuzy9MOvpcxseRjwlo8EsPDjY460CFzWGDsJwkYVy0tDwM3ZbzSwJ+t7j+FZ
nKO1RVdw+W5nNvTFTyua/YqZzVuq799bey4X9cYQVeGQ70gW//VDqp/WqDFeLcDu
OfxOnHFe2XzL7roW730cUpA9PUw1yLLhKbe7paoGe2Cltj+OMFJNzex8NjSXbBFF
fgdz6N8/RiOhGH3+uvVaGMFTaJS6niZWCyU/JQ2gVWnO9egCiOCy4rgg+2gjSMdf
RXTcvxL27vU3jJgRkgUGueZPhlwpOCqp4QmzcD43vlL4yzWXIHx4uYl3/uoh/BeL
ziSLt2qDInJwEYiaOOLL8+6dFyc/BuNVwVVG9I8rKqIj1ZFpUh6KVnFURKYv7Ciy
7uwBsKRFLWWDBo9XDGB5stURxBzu5cLgVAV7WBjItIqKxP7Dtlgh9Uq+sFuk9xoZ
WPF45/1DbFjPBI8ERiSX3KbFVTSS7CdGDkGXJi3J6ikjY3fuBeC2HI0dwSDF6qY4
C+/KA6CxNOKaHhkFcZmzrCJ2g0zaMBoQeVk4W5PtZ2PTpIHHYobqPONupo1pciPE
F2AAcfTDMS5w6rwqbTDyA7OkRQ4l/jBEPAaHXu74NGaqS1jSsYIwYlKqNW99hoqf
9NxE/O6Lzcr7/6yuSp8jzqZ8f52DtRN8UDwUnguGohuNM5Wo2fcUm6KkDdQHOvDD
ISz3cR/57XOcYdFdqej/sYBVGfbY5UBqCPQwSr+8kVcGSRI1VxxVD5wZ/velGUoX
5Ppv7kcW4psgu9dvzElKDCrPxJTE4B0+xlOFEAkcGVbRH8IQ1QRMFM3GovMFNcpK
OK8Fv9iC0dBiIHE1Kk+6nnN0MaGjJxhQAHI4X7kDxe1stU4SD8NJ+MKOoBq6LryJ
irD3L8RI5rSwt6gacRKKlAdp3XIc28FBb3j+QPalzZAakiZn50rgwvt0e+BlYdNd
TdVATSfC4zJMLJVGttgVKwJfMeg+UZbGPEHezD/8c5Qp3KkbCJTpAM/twVjrn1kT
Ov+Pp3SNS29P5iSoGa5InZX3upw1zCfWv9sC7D9jCqEDFL8MtNwzIMiG+f47Y6oi
B+EAyV4ecyO973pFYNUPwoVqQz6JzyAWu7pU1zLpfrRPsJBnjEtLzI0PjgBEC2Je
r8WQbcCGXJZrxnSdF1R0p6FG7sXlL9qUJfq9t7ScZv+5aObx4bS9Oj2FHgj1BVfE
KCoDAiEhGy7jzU6XqslPhsqPYJdYiyY5sZ550eO3qbCprwb9DT/0eXamz1VGadwK
q6KCniZ+yPenMXIohB5XInAkPtr5dHw5zQumLHmfQHJO/3Lt+TlKoOyTh7GTFgAS
BnUx+TAsO5v0a3lzzbs0dxAJY9rlWmqANc6kwMBPTtlZnxwqN22fscBwdpLiWeey
xY+BD9JF6tIERwT0RjxN1k0SU7usdKfYjgoXDNZMhPfC+17oCkxXkihpIBc4T+ZY
PkzUYu4cRJhIps8S6a1Q+JbMKjC5JSRtZOwgs9PUa9PLOynxCP/0D1ZLSHIRzj1b
aHn0sTe1ddtCdAX3Igj6bdzppNZ6NcqjSJsjkDZLP2kspbpYF5dwIpd4MKdf2ZMu
nLfaXhXsECd3MGH0I8iO5RlXl6ggx1X23CWO+YDhPhHf7thGPcs4/zCJmPPelNW8
v7dkm3UR+POnxF3+6Kn13maCi6kOTHQff4Gk0Qo7fOQn0gc3bZfPuKEPry1hFPud
Gh4J+B8VIyUONnpcnuzDZ89aJBEft2StpM5t2dRBsgJIHsvcklxA8NipzC54wPJY
76F6lXr+j8ZANJkCdSBn3Rk684JETTpii6UYPsK0f7DnJXq9AH3TTq2QVnFfL3rw
U9mlmleYoW/6kRRPAqyhi2/MQTt+SCszPlxiumdiLbqK9Cpj3A1nIzvesdEOlihL
Yi7eCfBBHfpjdtDz9fziJvhYTZbDuax+klUGain4o6WAM+69YceVWnx8DjsFngyC
AYiWMzKrE5a0AyUqkJfAtzxseAiiCnpMoTf8RPY8t/fggbO94WHuwMXalojhivkh
dUqgZ9RJGGZUG1SFb5cWNR5GRig/Rg4F9SgYD4OucGqBmMmaNodcGtHIN8tRRmvx
2s6hONYf7tWPQlvw1jZFgsrtDxwLKwDntuCGcDjH781hjSyo2E60B63ZheC9JKBX
+EJ0jZ91x5RKMVi0j8lM+o/bq6xX8l39eyNEiWHw2SuLCsFqNtmyLny0il4DbjUw
YTAA/0sufC86qffO0Ls2UVKNVp4GWv824pSc6/yA95/m/j+7MFbu1lC0F3qfUAEp
0iAn4LLpS02K42pSPuCrrzCwteJduS9+9BpmGMNLSVvm3GTHPN220xp+pJcvxcta
5NlmK1V/DMr4CdQ7zUg9Bnf2AvpPYmpdVnpMc1EKv7COK8EFXGx3Lq2FTrv65au1
w98Bytgk5K/X7iz51qj/sG0gosbEEYUkxNRifywZfMXEi8LHUDJn+BP0UDERojXy
wTUK3+VH09MIRlBHtf/ugNsl7+bWe+3+CvyDOfd9Iues32EsTy+3dEkv1h35T9fk
6QzbdJagpV7oL4hl5fHRth278ht1Gz6yvUrd3xBtwag0a+mu8Tm7BSAa2JiCDx+a
y/OnF5iZlG+4AWwzLpkxenOt2Eotni5Wt82y6iTzF0syH23tK9LsuXJ5EaDIGKjR
99NqelY3jL0zAeukt1Fzd+37dJy5wlZYdH3TGDj7Ae79HZvM6WfyxfH8jCo4qRdD
Nu1FWfPlFavqIv+7YZI2lbHAo8h+6uKNoJQ4jtF2am1jhRzldrTs7Vjp4O9TNTfe
lekSiuNLhWrPPNwTiLuWIFBaDOX4H36ucXIgQUmwjLiXU/cB2WiVg+ywCHx+EPbT
DKEgHJ1T8h/6XVSkrPjJIY6cHj5YbBggACKuwFdM8MSX0OmtF1RCAXqRicw3+tph
uJKukmgNDlQx73ZIUwUGEKFExIK8eVXBQ44vVG0+28WFHOS9X54bAFM9eNSwSgy4
M7fX5YhjFgeke1Ry83yA9f4TSuKe7xpuqnUu9Z2SYa8QOf6U4PC4NGrfdHde2AlM
vEqKubIb/ToHWLCNwn/vVaZ9d1ffR/3vdoThNtLIie2yR0HNAGqBP67hjxGQ8ErF
PzLaPrv1V89MHo/DcucWpH8X3wMpBLRVSlwGzrmmP7we1bxjVaqCVp6qAgRdvlWD
2hv6d+1BaRlnIiWcp48+84ojulJa2MURNbFz25nGD4S5fqLLfC5U/2fya6Vyh+Vx
2dqPidI4p78+Jh2fXD3raCylc8ZUM6sEebqkHQDAeFYYVOQYZ11/Km7nruBjrYHT
Yh0sDI0Sa5upbD41DlHv9/Tq+N1aqrhJTk5PYNyDwQDSi+kxIwwRobE3awDD2Rds
ULoPA1KiowXw1kwimP0rbTJEkcY2zPnIzOUsYeyObxOGjeb2Ni/53nNZQAXUnw8f
R/9dW+HIe12RLVy2ji3FAKrOZpi5uIxZRLKUeK8MzRvuUTslzGMKlaSG4JxFfHW0
llcG3ZcH3ztxYV8mGsQrgr2xRS49y7LCQtqTAg1xeCgbC6V8+C3t+Q/8bYIcfRZ0
liOcLKq8bOY2cTYqtEyJGGax6NYlbMtJtw+dJ18bU40pOEWlNsRLgR/jMFSSaIsv
6ENnPXQinMwxnNtufzRErYD1ln3pO9bV/cGAebO4UWa8vB8lMVo+5i+L7OMy5npS
iYDVSkgt7CItQOJBSdXoyzX5zYjK5rZSVPymqCM3boKOJSB5z7wexmDH7Y28lK04
zDNg0PqQPAg9Ryw3WZBRfz8M/z2xX+Oahg+vg+tH+Q4nkLNBc911daKHaV/9WdES
DH4aRBxglzRArhrDNU14fkLbJ+rj7nhe78egB0TRtF8+J5R+n86GN2LGJHI8pGSc
eE26D1h9rtuuHBuOTIGBEehQhLCbD39CQ0+/cBwuI/1+c8k0qACb8GcSvvhsq6mf
IIj00BhgYb4G4gETPlgqF4PQTBCyKyeOBf/7/1ujYx0+HElVxw7M8RdjCpTy9gEK
HnwMfr11UOsXDzXpqduovSY3EHNa+0pJC3tggnNnao4b+a8U+HEDfZvJpwQseRn5
Vo8dS4IPwAoUGaYaV2Mc5m597DKH3QB7bVTONss7nsYIRf8NI/yqTND9KkeSBk4K
AU0Y+UTXN5XhZln2Y8E8k1xZtCefHiFX2/JwKCM1iPTMparB7OYQ4FUECSP+I3Jh
+rlBWxTeBuQxxdHwiGWLC81FnWXtDT5JdGEUaIFGWxRXjz+7Zvcf5l0ljKKnQpfb
1ZrM5TrTmuCCUdouRSkKpJhEl4tz2qY8G3WbKgf1VsNcwr0MKZhC1N7M+l0kcE69
5M1E2qW0H+tPPn8cjAiHnopSGCtoTjP9ytl8ostzU9rynIe2qaxxGI1we3WDhY1Z
9PU95GKX3hh69+VylWVE/uG0Hq51H1LTebouzkCokMWBavbav+c2Ok+Xx1nyUb5j
Y9xXG6fB3K1+uOhuG1qOyDUfzYzykfTsHpJjkLvwC+C9sYq3Utc8c97v+ZdXfrME
rOS06TWqjHj8dEV2D8wyM1vCSbkV4YnjvCLbTZqqPypIvcxeN9aE5Uu8l+UAgdks
TsISkLqRmT2wbptf48ZvqoqNx53PEiDtOMe6zwPC8WfCpMJ1kizCaYP3n3VlblOZ
24w1Io1FLHg+LIl+VD5HejQzcnVjIYHSvf3O4ifPS8z6iBLSKYHo6S6QYQxS5W/I
M4564rJqfL/nwfdTje1+LfuxKsfhMIypF6fqSubEbuvTu2kSFiZEPpNRjk8bz2dP
cdQ+oOIPvxJCn0MIp8BGmfyMQ3yFqL2uQAtGba3cqZCbHULhKqKUvdiVBbmhzmrf
Ugd8b5+tYbHzmVHdH6TnsZvvZB/tXwxj0i3bDKyoR2qEkGHEKA8XBJXhygtNYDvM
p1kFh/ok1j2faNqhNXS2jCUac1d9hGtixrWGKtQWJQPxMZquHvDPWMYyyqGIGFee
DJN/mgqZ8m74LZP+vgWxXtYTlKGmccc+lImza5opKXaX4DJsXqZ+CWEUeu2X+mRL
MobFE5jH09BXaPwhoCEx5xzUmRRYj7PxXjWCQB0Nh81Ci/2EbXjD24sJSn8mm7Gh
a4RMJt+yZZMYqv06TgevsE71bRKBtfHXadg/j/JjD3bz7P26MOPgCUFra0ceQnZl
1xeCYOyEItrYLAn0HeaFdKYMeMx7ly4aW1lyv7uN21nAFXCH+Y3XGOlH0cr95+8Y
Ry5i5Z3ZmMnh6Nu8tBc6fCLPW64YUPY/dUJvAgSasE6wiJVlj3Bxyytr82a35q6+
eP4goZm9cCGA132YRc4CpwvpPBB2aNYrVxnDJlUwXP9cFtasrNGygNgP0DTFKMzu
aSvVrmKRyhcKnXFWZYe5QJ3CyAyvztq0Rtx871OEWjjlikNXWnc7Tht8s2RSgBPr
3yv9ekcMTdxgw/Gz1XFcGtmeSMN1+bAO6BxFrJPvR9gWi7ybIaF5dz66Bd1YkQTy
VxNNVPkDmNR1MoIfkcoBLx81XmZlRhilvTb/6/bKpl86PLSZ9xP56CN8EKTH+HZ+
OvQ+ftajFrg+Cv54RR6SpJcdN48Vp/Lx7Op4Yfx9BDBbEppd6ASht0IENqhXPn2y
+gMptmwTzUcoBDk1NQSNIHyTFHlTPlzZU/kD53NOODpxTkDdrNk4ivAHyEVi4Vhc
g+rfKVjqKAunTJ9unEWofc728z8ounaE3Doc9TAKBicuJZbt2RwObXqVQaDcg0J/
a8uCGqXXJaIV48iTwPPixcDJXTBoNck3bPmFcmSnC4M+B0mafjU/vVa7+FwIoFFY
O3NDkZy+c7Mc6CBKxInsftStk+4tYPzODFqqZ11XfJFmSwMiFp4eZApZ/im9UOv3
v4S5PA82+sD02Q5GTmKvWcw10j99l3Tc8h3S2Zn//84Rt6PG5muLm/JQDJT9IEcf
ZeBWUcVYVVzGLcR/rs7feML86dlgvvxR9617pmikN8w8K0BYUtkugoLsPQNPXhbe
IB1zlfZwahld/xDjZCC5qHpTJ75Azfmwq8IPp6vDovKpk3Yrekl6yre65J7+Ikdj
X7r2nKkgbxQBynhCQleHZOxNiLNyUiuKD56F0F9DalZSCKQOkHgNSYYb8HcRw+p5
/xfPIA5qldX6uBRgStp7yJettbEVsgsFlCB6T1BKpw4qYeiNDSIDOK2rDAqR7CJ9
7xifXn+wIK8zghVIor4GTRitkCC3PyRiB+LOXn6foVtqofLKDOWpcqe9EJGq3J5B
oRCzp7NPnH6uvssDsToLSCM0x+aPClRxAgBjWWXmoygY0iqGSfQYV9LimMtTVSv7
c1Xf5P1aANnhfiTRBNmhmWDaq6demB/SU32F48UKaTxJg/LbO9PeBtaYMWZZdHCO
UtVqU6EIHKtXyx686+47Ta5N40hzkAWGf49gDX6Je/qU9eKgRn4VPW6PVTcIfrCR
jAIzHbnkua0ra/csOip74VekUn4OXbrkNM63QXK3sjkQ/3ZpHFoVe64pjmPOkuKY
a6cPI2n8+ecz0z99ntvrdcA36oLWuy6d3+O6y/5OTRbqR22d2/IDXO03S+Iu1eHc
nyJgGCvBil2axpgWR6Dw5eo3taXPzt3KcNIW+ekXnZLdlswUyMSUMtgt9hBK269Y
90bk6bOXhArYYgtZhpEeVFQLofb8R2L9ZzoSMSoyVSNqWYCr3em+AXBefnsC2pU1
OwfNKFpPhEDFiEGI9c2PZAIXb7TmgTDykmDRSby6HvKdUks89Hw6r9jUQAVaeovr
bBz4wFUpLV9prDBHIo+/NqH224qZbR8Sw+BpU0IU1eEfHZzkBBqFRne9qLqsizOo
LpO8rrbKyIi2MQffKMHqn3QK64HzsbHEBK/AmSBCNDbV4SMhbgGXdPFkSh5IUt4F
xvz2HWiiipl3ViOyit9xJWHvdsEskYNqyGqia7tNYtjbN7pP5xKxE9BkjOa6Tn17
4Ckhir3iGpoA5cVDItCvr+SyTHsmK3XObI5diE6tGDu/vYtQAE/QiVELox4rMPpL
9EMXJ93/SdbcGG4kLzzvLh8uF2opWdV4AjHRd6h8Vj5yPl9fVouO+yEye1DOkPV9
UggY1Fw4BKoNIUvCPGtFrEVm0OxMPl86VgHucVzRaY/+OHMKaq47CjLuC1FthdWG
Lr9pjGB7U7CuW46Mh4iF5rcVx7BNz6YqkJmpUhi13dejg+NKV/CjofhVS2PYSorw
nuB4nk1gl0T3z95zOvaYNGF2CTp1HSl+nfv925IJxDFUfben07vDLTUE3OXqsVoL
AbnjjAUZRcoyYRQG71vsIVeWy3JeeE5vU69I1PES81gGGgBFyy1c3/metaBTAdEv
9n3ST+Hgyg74ef2Wch2/J3ggTlfrHjcEuGs1eCwITmqpMGeisxOeN0a+nRG0Lm6I
OoIEHsYD0G23gOry3tAoRoExzCssE4GEkNBVpE5uonbdhU20Rbe7UGxIXmIRUVK5
coglq5iVj2bCj72MDfIDxD/75mMfXA+tjdulsXZLs+d/NK7zJlVvVabyfcw8jxvA
km0XyL6/Xel954urVmuTcXqkc4O75ZNLPBBOzeu7zNh0sWNBsk+EEMYyvIO1nL42
p/j+OswfvKcff17yYPRyIx+FtGEj41G5apFvX6hpHePwRCiLVUnmD9143nC97qjM
njba8TISojVhHiy5rNy6H61kaNj1DIJO6jk8YJv71Rd0vpRqJV+2xvkF6tNV6egG
wmQYwr3NUfLUDDxpgXJ3eoyaimnZG3NVEDxIDLTu7Ma9WrSWVRA9/VkDPZGZPu70
22mxuUrGkVnm4Lmhhyao2mD6IP/w50yRo/V8q53HjC4ew5xp1YA32k8MFOKohkgA
YJD0Q/H+kkZw2ESk0JOvmcKMSCDqklJ4v9FpknfYRgO55IbKzhTkxsY/ri6bNa6n
jkww/rMGGSlHwZ1o9LB6D9PDSR1mVkOZ+Zr4+60jDkg8KCj+gPmQX4hTV+JWPgoO
m2Kcws8UvjAxXVgJ/wTecsTbCn1N/Hhee7YxBgr7523DspEYVgj020fLECsmjtkv
PvvLW2tO6q5y830iqj0sBXjEo3EvZrk64yI0oeKjGOUOLVNLBaffa9H+r2o5hcZ7
Mb6lBJDwArXTbNsaGoJMG3fVWYVBw+2fOTRJS/vANbWUooAYYKzJPzuqKlpH37TG
arOTCkVOmBzb7q8nRkapOWe+kzGUJsY0ETjiRJl8M2y8tfN/ILicGC1/coChPNKc
+6Q9XHDtj0/kj+BW8qzfGwKYBH2UjtNZHZwfBgmB0ciLoatHJ+X8vLAIOmfuhmOT
ISYIZ+q/YSGeiKPrzBtejLEMLOdiVg/eoCJzcKSdqUVkyOPwgu6aS14HAFTaRgQy
WCNoUeSRVAIrtHFhJBTYvzFlm4fyo1kzpT5/RlbVC7C1dV6vkpqM6PEulvnp10GD
v9GU6JjeHg2g7F1EHz72Y1aB/SqnT5q/TSryYW3x4BgLeC2fSWqth/V3VfTZAYcO
nMQpruN9C7pzPp6UFBMb9eflyurqTFzqwlHZKnpHOCNFYXKzpOGi0LZdsBDc0Yu/
in6k9tcMKjBUR5aIqCyz77vMalwvuKwgn4LQmjFyt7BPRkZ0Fc+8GVoGI+s3NkRJ
jbSw7iMh5t0/IfsjLPYxjEjIyGhBB/JAMyzeyp1yZVPpQ46nulG9P72MY4meetxR
dAa7AahvrYjQ1QU1gbFq94BRo8+rK94qZLcc7WIXKJcSzPGUCJfu5ooZzxITOgvk
VRf6/fdeLF1P9C90EKBW1NtzWxxXI70YltW3deNkJj4z1YErWAerHOJmy9BSEfJ/
F4DmO/TkXAKeAiVhxjPXgfLfU+SKM89QGxXSt3BmFFTZF7oFqge0DAPvgXkpLOkg
cLQaIXimB9d+hbU4TkYkNt5vFvydSfWBLbIKxi9Imuzn7sT/Qs4Zibxykcd8LuIv
2Y0YcpSv9K+l88YE9Op7VOl9n3vx4I67KbtVmqwPXd+XvB7SOv61Y6T2oE9AhpLK
gdv/3ACBVW9V3oHf7XFwgPwNdVufuHzC7oTPHI3F/s4OvlxJZ4ETYaQGO87/b+PV
0QDIS8YU1vkFXqDceeehv0PEDWSMLIuGCqdXb5wZro88glqOd8ofXT4AuxHBqoSR
sU9OO8t9otRYpFh9C6oj9QPJm5ZeyFJZ0r9sQcU/Z0AxEftRCk4sxJIu1k1PeGuB
U1+gs2B0FzwPhPyHrGogaWnoFQrdOSD1wzks9+dODmgYQpSzdGo4k9OrV2qiKGOs
YpO/Fu66YaQFin2/5+E+PlMQob8H4hG7VluxSQgK+9g4LW7zGoSVoJ3hu3U7/e9C
aJrAJJcQM24BC4yx0f7Z2soYcm3dq6OVT0w3VbnxwzYyu+8Abcei55cufcnPi4K7
khm+SCutQsoLsh/RIeNylhGDbXGjahnyncUFj8RTFcaw1S8qsJFqNr11pgx43m/6
4rf6/Q3bm5me03VnlU9fVW85qP3eyPkUCdKpX9wJd+n9zSS9Vqb0w3hmLbp7PlUG
oADjQYIsP1Sa1RilS/jJ0X4amA84AAd5VJAoSHATpFi3SGEz5N16oRy17oHevJBr
LBckvnMRwuF/kfcCkxQayXioyTNXqDs4i7CDN8gA46lJi3P4zMC9o9DBchXpESWW
l3KUQkHU82gDKhxZKiIs3QToqYPcHNIBtQ8tJ0DWUZq+bqv5/cITEYt4Wu9XSrHK
7AWr7KyKTERBjV2GfifoiQcilS+0r445dbcLDjN/G2cImVZcNVuMcIN4IhFxZ64+
SZOGfV5LjjJ66Qs69ADjbZ8/p4ixb1tgVzIlyHGj5AM96oYCFN8YGo71dh69jqgD
MmxlPcGLahNglFtQod5ijH5ghTejYcvgs17Pj5sMrntoJuHvWS2PudhnDubBglD4
7VNyigWyuCakTikVZRLC98R6eAMi0926wqfwG7+kZSCG8r7FRsAoVj/7ab3GJ67o
lL1rbriQelOfON2KThB8b01JjqUARgvwDkFMiGRSskolvfPLY27dmCT2WAz+FHKA
u+JJcpUVtPrW+ZvnWarWXG5i+dG+RZcRw83OljPgie3+HAG0oEH/m/zhsunCKwhP
VlHyNlaLzDI1GiTG7TXptlD/bLNUldP5cS7Y7lXNztL5QRvqBA96Qu/OVgKXVcA5
aYkHvubfSh21wsoUoUV+PssO9JGqgilL78gR5Twv+jIsYUFjJyuWxx3aF1Bhg/ng
DSyPdbHc71iSnjGq3Spdjq99lhjmWxHJA8wI76S3uVe90R2OCtQoxVOJxSCwOT2l
UO4CCQKFnJoQcGvS8vyYLt/E29a1I7M0mmh85tYdHWU3kHEtLel0EJIg8Dhdih1k
3Cp41buKX6tumjBOBa+sRvzVVvbBgrBoj+8vUr0NZe0PivTbwfnCc1bsMbDHkTI3
QyOf6R5RFN54mkSo18YW+VvJQeH5gdJi45b5pWBIkrTxKWF23ez30Ewop/fhLEzM
9wt4u13VzUkp9AQbsRmHYaU6+fvDUHV8s0D3af6bM8KHBXPFydpeoNDKItzSHVUA
C2R2N0cQw5WAGEZoIsVHXNyg7DOTAt6PAj/t32NRWrkESRilg0f1q6UXsAujy6oG
WHKqvrLKQAITaaOoZ3Sf8lio3uh8441D4uV6VM3Bi/+7MnYGa+Mqg9wTUmM4j8Kg
RxB39X77EqEtqMMTLrMSOgdnFDK6kTfVD6YdcJa3FGrRDXOef8UQbAvmYBjnp53u
ths1DJYA5i6YHBCm1Sd2kyJgFp/7lBbNpaNEscfcEKpoVDxLBKg8Vb8kAx9glm8k
S3WY11PcTloTierishUYdra6+D3tmaBlrXSzegxQo0mKZL4C7N/+68S9XMVvoi99
Jq6sglGvIqN7veK5cZAkSPBAOxeIyJV1obLVJwRaO4NS6saE04/brX6PWgU5IJ5Q
mZVZt6QJUEsxf+VWKJ5GqgUGKtpoTq/IbD3s2Fh+BinewMubybJVVH4KrPePlha7
jVwrtNYKOQ2P+HHGcvmzlkEq07Xvexv3K+mijzWx9ZhNAHhWPvm4RWcuJzD8oRly
tIN4aTQPaCCRmBgtZ/KMK8rqpjcDvBjn/oLRRj58nuCAFG+4bJLPebtlGPW5G0mS
BuAb3RkHw7rawv04Yy8wN9S6sYv7tnmGw/Am3CnuFiVp7Y+/WDT1UNEqc8vpFjPs
oqZzci7qjfVgmpnk7ItaXgS4mpUXUiq8Ft8blZnhlT6MxT5BlIVhesTQ7E5kN9Sb
0vGEes5LUx99FnAke2JHfB5yb7ktdrN0EzjAYj02TakZoE9Jsh1+s+E+Dmg7pBex
R5GyHurjcz2HoYZaGG8sikZTNVu6JprsJxkgnUMnl25lOmx/u7J/x2LyYZHUXHlq
+zdNr0iFewvHsXDKNJ5oxb86UvEfy9yEE8QJ1S9Gj3jxhC2IR4aoDKfkxaWo3uwP
LZVjSJExasbDsRBwRRWgkpnCowUJkvbmraEcz5gy+dLCOUfM+B2DOOz4sgo5ZbnF
qv1kM0Ky4VjPOnwFhwz7cwkIFF7pa6SgIaoBhv7X0wLVqu/dxdJ9ycu8j7lDeING
GQAGFTbOMDuRt9fAozzwss5aBxXFEO1q1Jy4Jw7skZ6SRJn5xenvO3HL4b5p5Izb
Z4gyDVmhkxIoRNhge0QK9CA6S/SKsXuithvqo9afdeDO2hBlyMpblFqqH7xqwvRw
xsMVJzyyiOTPks7nv8cmW8byDjqhAhCxZ49AN4mGxkh9+rBQl9b+wONm1kxnEdB8
571d7+DH39GWDspLxljA8JgvVmzFB3oEMr2Q8R/QEp4m7FuFvcvk9mLnwVK9Ita+
YzwGtqWm7b7EBoH9very8J053/vJpz9z61SdQkA61El/NC05e6Yhb806Rp1QEimQ
zoVnTEghy5UEhGucUuj0JWvbM14LHFMiseSb0EsgUyd/hHJj/wPfGAhT6uap8N8V
/zcVTmo9hoVl/pARS+x1QfFetgFAzvGby+5h4ZPmZuhBC+Mu/thVVm9BczpLLaV0
BN62zU9XroxhvpPPBH9U7uTretdtoADzF1y8ZZQHThPc7ynCJoCcA5MkXbSLIbMD
jJeC9Kt1USL0hoibHuUgicEFTg3BAsjJUcbbX0biy0Fc6zMEyp1clumDpdo6lP7I
/6d1OO/FA119B2TMDzAQkZygZF+/pliVQv3cr3ePDUZKUGxkqQzzMa49fPsKWPxe
orY+66bGx9CAA/OlSCfX2wjrYuMiPWd8Uy9vxqqVdocU9So4/BlzRdFfOBI4LrZQ
03vj0yLgm9JY4zA4wRjgSBQw10biiWmfQZXNLKwxOYs98tGM5krPYpAqelytxWFI
76Brxlr2BVUcLev9f9TxBDoVBK8y5QLn1bkrv8LJaokzByT0swJFrOGYtP+jD+hm
6irfkT6Ys1XfIAUJ8PkPy12/NUX/McDZoH7LHCVG4oG/2Y8DMcHXJYLAXEDguwZC
Dseu371pnt9kT2uC5xeqbQRjk8xBpSWAw/JtB8Aa14Rh8oxCUwRCgp9fwRHNGiXZ
MEMul8EvjCLI3gAuK8uvUxkKNFs4ci4VJ9lSqm53JViEFKwk1zgRHEGxuhze8dej
re/pXfU1A2T56GrB7SqmmrqaI2Ca06GvCKvvoqDEIIPYzO386UA12tnSi2BiEf8n
EyShnkWClYTmNtVYnQGtMOKcs4SKzk9CA7Gdw4XQ4BOw/C6GRea9OOgbC8CixUSs
F8inb7UaNDaJ2Pwa4wHXGfWIcnudVie80QmEh/k03xZ50THH36sv/fksx3yYjlCQ
iDwguY1BsvECa7PMfiJGBKP5u4H/HhgwGZT7P2oIpbbDSL4oAVjiYdQIzxtqWJgO
NSW3yUITtA8JeOeAUJe1PG1/oeByUDacZUrW/jTDfa2pIUeU1kKBf0UKYJyTl8kI
fQcTN8Lfjywa0hcOcOlPZOVgp805EpOkoYNOEu1L3QVwBujJ+tAv0dEc+ptO1HgZ
pWfM2m7XT5QiOnfw198ZuxEVIL3IIYF6JuB6bMm9sbMjXwHCZOhHKM28U4kwiCNs
Nmnh91GPsie6Zmqh7CYlNCZQfe94MvzqmOcx2sizv/kJIF5l5T0kxCHVaO25b/Q6
XoCq0CNhSmTXiwRbigniDECuvhiq//tITSCYDeSDHvPkQXbjEGKuOvDmoaordAqF
d9giwY5fAA28DD3IrM4Vd/i7WefMZnKpNUzqbJwuBiErY5epnci1CmuBYkXKWkvO
219GHHBOC2AH1Zz53QSYrnzYZC8YMzgYfv5SOmXLiN7h/RpR71KO7jZXXaVvtC9Y
Bopj6oDvuZKmm+b2Rv5letHCXy55MrhkNiAlBkuGm6oZl5u4djMNKYq4dkioBVka
td00qPFXDwGjIKV9JmAFHvPnepjHJH9LFbaTqN1aP8r3LonFCuCHq/lMeIS04NVB
IgbSIoXv8lMomXyggspAer8Cr53CBrlidfIuEkpR1vAS2Zsci7DaMcAF19WVNCNA
2op/azMUTBM9SkSAd7ybCFW7AMksF3s+XGgM+Avq5wNAeiq6I6MYSYCjD8M45CGy
8pFGlrg5Cs2Gc5uwjkgDIrkqZKwjhzbR9nl5NHJzt5U7xugU7qnK9gi94Ks1AzDH
xcjxYDgoMCQiQ93Mbyj8q/YEKd6Kgc+B/6HPFQ8o+JndbOP0JbkhpC3a+lEsqwOG
jiW30kvU9NKGcTLM/uSEFAPbExcFhWWghArfQp3Pfzb5fnActoTHB8r5U457y9UW
klAXfyQUbFt6DSNzEd8U4ivz0qBFNjKlPPvNV8X8oMcyJ6xlxI5lwuCeEyW7JHUT
bMNvVFI9/Quj+Dl6DVRi7TYQAj0my7sdMRC4PNMA3nu2V8Wh8oy7CrY0257g33SG
tupnVTRyhqb1GQ4dEOXyLb8r4T6e4wBodoudyNEL8xfySTs/s0+iaUpKCFCiQDFW
g3stK+b1NnACe5kAqSS+X27e7WDbM5llneuXU+o/UUFEA+zkG65c+MPycQy2MH+s
GOYYQhiBkzoh7MDQqlHzpXb4PZTlyuOat5MEKgAKJi6DBzo1wQQXYBbTnrFO7D+k
VPA0zumoQof0JAYjxkKeSKURw4RRPnllaJi+C6nN+lmPn8db++XMXXluTdmXh/LY
RTdUNz786YjtFoV7+1HrdsK3jS+eB/uEt+p3kBM225T5S9OfJT7OkBNHlKkIJ6hQ
iiS2R8S8scr9A/aCRj7UHCTWyjWZ8cH42FgfPWk2gghspjwVU05HKGRABYC6SiIv
zKZ9qSpLFraw/iSfHjbh4vSioPekuDNCWcyZZuROppcM5T4FJkQzjAEyN6K7uGmX
BQXSaWtz21lfQNHgz+ovxPJqTq4RHFbUhGnFr8uX1RNf1zlCtPmM1AWvmuu1ORL4
d7kSgJjZ285FixZOjUv6NrNGVvSO1Nl6Hw0eQNJobXKGoXnRV2rQhsJ+ue3ZgSaP
Xj1RCPe++muif0a7OPUSPmHrImOwHkFTc2bLnTWXZXITKws0hOJj7cI6AH7DyHUI
haWvOQbacCkhpHlwS/ZSJptJNax4j7IhmY2iKZwjpbczBTTzjNziYBTHS1d0XbKk
jd6hhXtYHePKPjesMFYWVSmx7gyGBFyzzCE80ViXfBMOkkwMPdNObLuWe7DKI/Z9
M9basG/ZCxKdpRfYBA07d1csvSAj5J8dazSZ+StWKOYn/KHD/EwvgPqv0W7JO5Zv
3cL26wLSmsBNFRVLH/Txm8aNYZZFV9OMLENnBX1Xw1MH6ZijNWAac+9knkFhLCfo
4tOxef/qjPhZgk27f9pL/Tt4EMjeOO9XYxNb+Y35+Pbn3K6+zeXtp5+3pSSBGwJn
rLYuADF49UKXhai+zNtpkPy2CEJcBghRNY6wN/aEHbw+VOLdNqFh3nTZmo2+CINp
cCnrsDH4bS1Hjivy77NP+ljE8LfBU7XlIyef3PhCHsWvwAvRVyU+axMrPXn8xD/k
gTUOfz3QvTbBk3Whe5Fb/q6nFiLuaNh1wt6Td9s0QmPORs0SC/7hpZFoWl6OQVba
wKZS3kvr+/wfGhjV2l1PWanv+v5USgcF+RagXxNactyfGTPgUCJRFxywjrLayrL1
Zcuei5xgW8+WVI0lRly+/8eA3hzgVZDGuJ1sSrjf/fxMXKA1z/y/s1nzI7lyregM
1k6R/QhsScbXT3rPdtDjInGXEiRr9wdyG7KUucTj+CWVRrhlpL3+D2dGhIN6b0dY
XQENJb53nxPNN/qvi9CSQ2XUNcyHFfuq+oXOUGT/O1cFtusVglNE8xJ3sbNFPbJK
/cQCxk+vDawJFpn2IENRbCEnt1vgCKEbGZNkDEhru5cP0+5GHC+XS91qEromNA1V
HpKp1e/siSqC10jrCV5+6+RsZamGtxS+cwv/F3OdVjGBu5rMU3aPzywrGaUwIYlW
kQUOXOK4aIKdYcjjLSNAUar7XdQqBCZSL1CrQzqpE5dj8eUjjHJ1fZ+Fd03vFnB3
9eJOI142PFtVfU4AHoC48PeAdujZMMRbXOiIGX50T0ADS1eJaaNmucqrTt0fkrov
L3pK5WH+IJQClNUuKZ/hX80re/Tmwa6P3lpjEkQ9QfggREzwQuW6uSXDBenqjthN
B+fTKP59Ai1uL/h8G5arjc5t6Y8FJ+TWXw4Obk/10HQyu+8AITVzhDD83yHlYFpm
on6UqRdSQaS9BHFF1R7hNHgIw1NSDeNASDG5vtlgSC5p9dNWSzgx6vauZpUKp8l6
Ze5CghOThtWVq+NEtzxlh0ZnMGwLsBTIAgO2/kc0Ct0TwGOuACepmYf8LbepT/Ty
//Z6Mq+Ou7Cu+NF4MjHDvMil3R/J+JRyLRaihD08vKb+CW4H9bH66omN/pHd8N3X
1tphkppwGkFOLN+cd2NLwye9sEoi3blHCrqooW5376Iclybyg1NIm9TyYUHXgUx+
geul9m+E0pWDOd+J32gvZG4matiA7dyADthZJ5JOZe6dl5ocsx/vfR8yMj+zYCOD
B50BRrWUucWC5V3UAwWRNTUGO+iwCKRtUp0+O8ybAy5ZVQ9Rrgqbcyw2fFnuayzd
t5GrX0ZcQwIADTo1++3Jd4PvgsCV6S7ObbjyWWFpT8U36bJXThNv63nQ+crABYfK
9mYWS9MkQVR9ZeAuvWSA01CG8lzfi9Dk8JfzBU2ZA05lCmfDPWXpr0tNzTIMTVgx
nchhJ2Ju2HQW0XNnienjW4pkQ1hKOX7eP7an403OXF6xDKuLms87H8Nu02+PQQtg
+v+aUgJA9kINhHogByAMNa3g18LGKPi/cdUWhjVH6g7k5kd8pr4jKzX2ubqr+f2+
PZl6yZUF3Wv2xOEwulNPSZjQe4dl1lB8zznn4eSD/Z1Z/2Z6PMONb5un05/G21er
krx7iHFQXB3VKj92VMUVyoAYRxrtd7vpSk6d5cdjGZqfLiK6wNWYoztZ9JJ5+oww
l0FubkIxJ6sPBj+0tNZma17t8qNtEoxEcNsxJ9W1OUDbWB21ZzUIKsE1okPpCILK
ahclGl4grYO98xWZwhz3KzNnv5ZBz36wQyfqljQr0ag4/OS+o1XvPgyo4Vyr2z3A
bseNvr7jTN/FdkgOkzTSnVuZGk2iiath68HMmWAnZ7yBKWbJCrYjANyMcYX4f7z1
IeFgzuPcg5XNlotOro0VC+eicoqlcNj5h5osu7gzXI3egVA4JTOvwIdLZNMJTSsq
BDzZT8x6nVmZsgOIJHK95Zfl2zA2ndQ22CbbGjqimvc1De9qrYIqElxakD4p/QGY
7/mCM0t/6rPQiKgyyycu6V89O9Re6dGHeDYolkLJlbWIy7Z2Zhr2FAIcH7zW43fe
TIpYOAJdOXL+xJ1GS9vd/LO3QMcrbyGdQPPGlUFSQjH6iW6I3vH8vMtctquyMAxO
CXlcHnM40DwljB9QH53o0Szp6cPBEd+Z2ZhuVlp0vZvw1DwURVGQNSDcUR/Mf3x8
QS2SOD6L3B/f48YioMoUrmi2vqIFtu9+eKSitO9ECngSNIDyQURikZBYtdsiirEI
hWaWj67PsplZZgHvESxsnWxsoO2e36mJjR/EG/L6FC9hCtFLrijtBZePlexLfoh1
YQB9VrOchnV0GDL0bo9vLbmEgkF6tFBt3qoS0wjPME7bvsZNI5TTGpn/CIPEXoi7
FJoljb4vL5Sr4rSv74M64klJ9WTNK1Mdr3j5wU2+RPiHGQakHNAUqn1Ttm3Jv3yh
T44o+8NPsVRisnSaLFmswcdbuajIJRcQWup3hgYz7KBFm580rpenPVD9vtABaMyk
250U2ycsIMR+/t6nSxB/DhcVVADtaVQta0T6qktqYqavFavhYHMEq3IdRJqeDMmc
CBf9IpPeTd2tnU791I6xx9ro8bF9BVgW/vQrSnu+zrCcu3LHBpaKQYuJA2j1jFhy
eWFx2Dr7SA+bq3IdBwqF6xbyX2jPt0COD1V6JKQMrBuq4mKcoVqV8dkHKkPkYSNM
iD6ntCTkqihu5GKS3WhK8BPRDqKwMoL4bJDd9YyUwouwtM5QHBEd87cgGGcdkLqD
brrceTAKYKgRVitbKJyTa/XYIP9LAfK6HGvaGYk+ZQwkOv2dgIQ+oImV4ZtqBkmI
X4vvaCzgs1OW8a9JSF/Ic3QTnIPKKfzcBLzF3K12bXDJyNd1q41dw3lZoAPxrX6U
wOrFEXvX7+AsnhKd+VPAbobLPG83VwxlMPSTzvENoFIpdp3lSQM6qOYwTt+O6C82
BRfNaYRVFLZ+JtU1kSbElhVoKsLal4gvVq8OiW/zAvJ7J0/lB6SxEAz9FArLRGgi
Slx11XHwUT1kentBmH+HuuFfTSJIerEuttssLQyUo1fVfUcEkkvRfa7NdUAOz1hj
r83JfL+9uTFcm2inJv6rLrdjd1njvxEOP5dbIFYXzOfCyHX/MVgEp61m7kkc2xS6
aZyeyYrViHHQsbWj8CNJr68gm6XZTHlNY8ApESjgAGWmw3SY2tYSF8TVafMq/RRY
GjYk7pfzKlQbk2Iwxo3IodvpJs+uM2ii8qmQSAbLQAquqYkBSTdRufHqET8uQur/
34a2QL9FVq9B/pSgcKW0cJ1KEcz4SKBi96B7Homg6X0h2qX9JFTglNPKp7R1pn9V
pOt+N2ILNQPOhlvEj87FPTDC3AC+imfG7WD66AdvDx2RHSkqz34qojX1l8LqiMAu
hwSJTnTrk3jdrlcyhiqXV7A2JRTPpPQkcOKGsBX9KmDM2mPVd+IFS90HAbjaV821
YQuJOsGOQ0dqj4Q7Auzbr2x9jLhx6kLxHgC8DUvaJr8KUK6nS450ThylnaCLeBrt
yR77brYoRaklMyBTTuExb5gfl9b0lyD/RBjSjQX1ot6iw9mVpjbgB5O7SSjYHzjB
sU0IQWA27/OJVeF2cmsKlgzdKqajp69YJi2J5FHpe7UmdhyA+obTOaXzXUm/1ROW
ZHBkT+JD15ZPKrwtDIhcwhF9eTbx1rubf6I4OHu6z8Ol03knxnee6zrEcMdtr+Lq
ZN1FADMuKVZtIpIFUSYZClrmYqgNQ+Fvncs5USWnVnrtvic9H1liyW/di/wCWGnq
bwDgytou6g6PtrwPE2SrNMRLsjoOoeKwaZ4HFOnXw4a5g7WNJj4In/rqy+0KFouL
fS0S0To29GKEplZ+TsE8s9BcVx2vqspqSwmJM9RjmRoSUw1hBPQ80ttXrGrTVwyH
tsTArLjtzpecIfMSGYQdqikDBkAuv7xrcj94wiFOBb/jn5i0iS7E/htS2RE7ZgBW
s3p7s4W85PoIUU8O9XbyhNt/C8Ae1b1Fbq0LoHZ49+Hhw1cb2BGAdAb2/mo6lhE7
X73FsNZ2f6uJ8mo92i2wYCbgEJ4S6/G5wd1Vqeb2nD+ybIsbRAEVOVBH5qmTRUJl
RPuX/cxg/UZj3MHnG/6Z2OBAAP9x551E3mkcisLiB4rBbOKtZg7Jao4oZfAqijuB
XLf1ws2oAcWEUoSUCMlg72fSjpvQ1Ihdnbp1faE2BO2w+V75VCU2s2RCEKeiaNWJ
z0GWCIS27Auz8kAKYt931qfuUYBFW69h68IwSlco3AwgMCm9z7GncqVIDMDPyv9G
Pfui1YdW8lYVw9B7CACw2kWPTFKOObXBGC1BDAEumyQsggO9voIs6iWtIqra2Kf9
/viApQguvWlAw2DR8PJBXNZS+QmyzEabF3DJ/GNw47lcRoilQitkYP2MP5IQb0SX
LdoQuOWCAodKGIaa39qxNSlsIW1hDdY7pPhnFUhD9yiotQMyt3rBZFmkAZxh/uZ/
nMrN3uSbc9U8kv1z/XfbKvkw4qZKt5zs9RNV5CNaEEDhdmZ2U/BamAfS6tc0Wee6
vlAGgNbbAGE5e/ct7E2OLwb9WV96BR4DyNxcN4q573Ymhtha2i+FDct67eVRqOHe
tknuYjnupqv242axJHCRKZG5bxmQ1YdsKGWHjcN8rT+pWQtKw5ZxzvPOc0Rp1T+7
ILE2/JRmlaA8o9D8gXHej1T/GTF7J/qeQ9ipT8ae5rahg7ElN+5sx3/6hLuDrH7B
pKCeqGUA/q/v0ITfgYWmBPWEAASA3kXOIzTF1d+k7vk+ob0GTSCp1WjkoY1T1jJe
AmpgTjiAAxn+aPeCmT3GKgfAQefc39AA0UZYGHcAU1jKvxG2Ckt2t0EXo1puoZQN
vYS0tdDjocywQedWjY6AM1bEG5E6j3MKOCPqZfrmsIk2L92K683xz+D2xhBbB+Ty
Q69u08l906BAV/2J0fcoGqd7PCyT/PzqyQuxUqA/HKz8ODhoHrkjN65PFsqzz/sM
X94i/F+CeCEudvwUA1mHsLaU2VsIRU013oQ2l+qE3reY0MXrBYjIbJ5HEui6IwDA
iLCY2dcz1HIdgdjsweibUIN/0kVJzGz7t7PP5w+LxKKNQ9UFtBIs508PokGep4i6
MlyRl5DZYDHNyql5Uh4kIHb/qlO2m964OPz9jbS7FkfnAL6jyIK5wxKwv3Uqzv/p
NdgEvCw6b6WRkWv5WbW/NrOrkbfQBnQRequjZrYSYIdCdSpOT2J0MrlLhodd2wGR
z/CTi09BeltAySFP1dvcTRZ8A4c5+5WEt9EKsoIYBy87uy3U3rB1NfOdH/1MyaMB
pCEicl5S2xf3PPR+0yiPLaFGs8IOXGwP5QXfMVeYEiDCCxKdzP8zj3BINdVlvhnu
fA4zyoKubbX05KaeP5JFwuSa23hQQvtnpF3Rvuv7ddd9tps2FFV87ZWqFhEFSdWl
hRoyL39Lw5oJ7/sCWziAJY89E2nnZadaKuaWXbI588gk4Io8Nap5BUs4jaJE0b7a
E+SWfNiw88u9ZhkJ5OtpR95GdPSphQZwESmRh6pMJ9XDfqE5NX4cY5atur2ba7ee
GxXjsFpcfb6wT9BTgfImxjWjMOlfliBKppzyEG/4ubkw/0Akkd3Ohttxw6albD8I
P6RJn3pPU+2ZHSsUArvzw+cWdaUT1LRf3mwBtEYEeYbuzeFS4K800Z4UAwe9cw9J
Golfdj+aj6OYv5SFlBfaHPYReQVUHpj7cfkdweYqiTQtdhDkhjjctxxL2RETGBjb
+3aLh+NcscaOqZ31UbnF0pEQ3eLcQNiD+F+Fb3YXJYE3ApDAFLElJI8BQFW3Yw3I
SSY0swiPtW3gctnrezzGlfcRD/iUx24yME4ISFYlw5DKGr0ZdNvJIij+rwrJ1mbp
93PylR2osoVcqyj6kprIeyRZ+z3rKP8+DMqO4aytyTfiFMh6d2guQgdVa0kB8dYz
bJoqcV5YURf35yjAIPTUlaEz7IEMhn2u/fyfcPE/NLlU3FHLxpAq3t3JFlzI1Ojz
8rJ/JJL5mzrOfMzxd8lIaLQ1pTMnuYGvUcgo49eav13+SgcassBk+ysKUzEtWVVX
HuQldEmpZ+t/Rx9RznuxrXpoDeaOAEoTDHA/a/MZoEej/hLrPqMkmHg6Q34/4ryg
4EclDW8rcOMSyyZAyxO/TChOvOtiOUznH1LglLYGo+2Hil4rjmvULW+UxD9a+u66
HuMMC5fOfeCs4OfMtlqshXn7Lec37Ti4MtSz9/ApS3JAhcRVBeNXwzG3McaTsc2f
ublzHOY6Epb6kpNQ7e40vixO/rcUOjBKZGsIezAjJIm4L/A7miRbYotwO0qcxlz7
LwynezVKzgXT0mf1eJoG+PQPsT1bJuYj6Tx+B4e5Ijf3OpN9Djrx6pS0Rl5mAyNF
KQLOcSgXJwFfZawP/BvvpTInC/fFwm066OMzKOXgQ96DeUuNbDse7fJZr8mFBiCx
K4Ovw7O8WadIqaA6aoiopUmPcBuMvSMch14iVqF2LziTsHwhuM2/0S7u8IG0BAeu
haBg2ePNYgv9X5bCxnJmyh2Aut5VKP3B+/i/t0B9rOgw7XX/wxoJnc8MypjDk9ch
wvniHAw0CL6OaaLJOC/KR0+B2ln6oiuoWb/hT1G3qEVam+q7RsWtsbGQQUB8Rs60
OlfKSihlONJge6z7dcUOS2UDJbd7NNqGbnF3R4OiQ+Sc6Cvczyrp+EjmUTcYi85M
L724NM0OslV1rLa1iPSp4NLkOJKCe5KHt0ch4hokA59OBBCkFHF+uTv78S6U+N/u
yaISdNmxjBS4vM6M9zNbGqHC8twj42ii9c5/6N40KiIjr5Jiw+GFanXMG9i9Lrhs
aS7aZ433Vt4LyeYyXPkufehoObyqYyTZV+IDc7m9EieIbQD49fizhSEIH4aoQtvL
fY/KVxCF/MEktaJIkTTkLlHdzyddeZGtNeCHZPuEZ6qzDCXVZCyxZ5gkkL4uSUWs
5r5sMJWkNv+lH/L/4uK5Fn0z7+f8Cq6XYrwH9E1jqJhsr1R9Wk6uCzQ703QQpgWO
8MoRcrYlPpFyObelDqLOd1U/lc4cMK4qPCdcCoEuy6C1Q5f+tfUyKOyY44yWrbir
d0lICw0OiRAtG/opSawJLthixz+s4rjf2pAr4SoU74z/bDChYOqfakYjs2/YgaYI
WjSKtv4j5VBrtCf1bLRI3E9lP6jTdXf54bnQm853uUzdBZCVI4ugD0M2b+Ifs5zV
uHNZFFqkII7ocrL4h2RP1wLZP7JTCZfz4Xi4tbPb88C8SozYrb9DpqG65SS/Vd7P
Itn1Hv4DS0/c2nn7jpa7lew29pjDAkUs3V9p8zq4B0tBNlR1zDmexDcQRy5c/VaC
GKHGH1U0zihL/O0VAfNW8cfpTrsEMAkkfLygPJrR+hEkQvWDB/RC9ER+x117+0I4
LX99QPA6Ir9yTd4BUn2UzDaU/0d2wtvoaz6qHyDRIvAfa1i1i9G4TqNr3K64BcoX
GsFijMWXEsaqUSzZVAXLFgy1eg4u24AUFKv5nlFput++AB1j7OZjhI8ZlzG1gZj2
V56267LfLI7zAT714zPt+DytpTBRF2dcHLDF9jyBlUEodygoD9AJSWaZWLCAR7VY
Ci3Q00j8vE4GkzDhDKvi+lizTEw74DwglPl85e9fZM4qBxB1L6TT9G+/VVTih19s
xiHuERiwfXpCrTPTGqFI4DaMYv2a7X97LRR4QEVa3kFOUfpWnXvsrWirgw4iZs+s
4k82Vc1RTnAADvIeEd3xYXrLzGP9d6eLRLbZs8tBUblntTcgAwepKS8vlllJLylU
FPBmOUpy4+Lq1CpoQ/vA1OPJDb0uK9atlRPtS4UH8ToykFO2iPZyyEnp//CjevVx
SZWHEyuGFAZocMNL4yKMeX56Wxmd5tNpxLx3GckQGxyTDKG0+dzoHYyvx+S7nNpz
9+t3XzpiHkcSktmHdMF3jpoqoL8z25V2hHwbwJJjJLtRnYD/baANrW4F7WhVwFv6
AbyMbhb9QJVCzWoZyLYu9KLnjjjhhXgIXMtntNqwaUsC7GEkOJBDarKcqzCxo1kL
Evc/+MfzLBLrXRyYr3A4qtdBShoE6eM9syltch9e36ozx8wO7uWC2SwkviYK2uPx
ihE0EGNk2lnoelnaA5nYMkr+sgi0pApXhN2oMKleNrVlX4s8qE66QJwIiX3c9zL9
P25+rceAQ4t3H31z53pGNPSt9zHGOicX/b1vtK/HZtW616k7ysOjQw8uZEt8Gsqo
zwMaD2Y2n2eMehVkWqb0Okn1VpRzN0p8cu24/4f4b899XKFgcTP+QSVrD04s6ZLL
fEyzREpwT8UIYuzPYuOozkobYo1m5GZU8v44t2mycXAP1nmhHS5ElPZjDznEY6dy
sgwUXyLF4fyLpBwumH2azxW31ULlOcWo+pCmuDhjfCuxlNySu21hZVd6OpqjH22h
WeP/suca9ayNANTsWIuH5JvSxQz9EWqk3ujEaS8/Pu+kwFlXEcMXcGk2V81oy+sx
9B/sEAT+9AhTR+tjbHNYs7EVcgVR5Szt8JTLAtIc1EgasdgERbHCRB3P7BdZqbKV
iBZ4LeSS1JZ/MsBDxfuwdxggXZ8iHoeonIz++zgZw9TnNMK5e+7d5wNZqY3dbmT8
CYnl/t8izVHZdrQWfnrVSlHbf6u7P10AoFi+Ui4poWrMnf+BSwZ7NxDqIdeHZc+A
vWqDIhzLxqTzD22/t5w9Ddm8ZctdWXq9M3ml5ZK/wS8g01oC3tnIEkID8o28dteR
eki+yiuUsii3So0r9FyqqFqNz2Eu0nAfOrA6Z/rMNMfphEl524m4foS1o3iiPMbx
2l9G94fBBOXcSBXUbppY/y9Rm3gATytrLA++yxdRrPQTrDCwmn/ctkKc+jZHDV1l
B1UP7O4ZUVoY9e5pmnKR64L4dAFhz80W2sftlfxFSM5G+RMgZQ9aPTniO36TlAXa
Un29tPnMMR+b9S1hiv+T/hek94lo3HmddbEGkUHC/CI4KtKH2x1+S4uncbZYYPlf
wS7u+wq3/3iIC7g9skEb59+aKFG9fWG2256nEA33kuq6bTTQifsL8+yz/++CX8hi
WeYVxSY+wBCR40b0+YDYfi8z1NBkXglUWaqD5WnhxtalpKJAhIDEwlwNE3J2sD25
NiCIURxgoj00vdedQWVG3uf0aLdnNx++mbQUdzSc1AFjsBC4xdG0lZZWZpZi7fXg
0533wvOr6vvJRzD2VmMaoZrGkr4crA7OsM6+173HKhp226CJQjNwJAiOcTdMHEPq
3pPJfg5djaqf5u/Jp+1rnqGwv+oSaMEulpApCVmmYwoRSxeZzyvBlrWeeSYzLDnr
zoBTVRr9Eg7riFE5aIUuObichB0l64dEys7X1ZOUb8HWItetcq/yr/fnRX+C2wBQ
WaiMvPhTNToUw0koHybDn0wC8HgQ2EDmFm6zubUGXzCg/Xf3IUKE9CwoFQDOn85g
oD0zm5cQDccO8U6JJg/uExCrssBXtGoYPLttOXCMAP/1w1MUJd4IEz0dbeASPQ8A
zRGtr/qHAVnWSvZq5mJJ0mzg89+hUYljQCshkoqez6d0BAcNc4bLKu40Pnz49i1E
RH95oGlM9LeGmz6iZi/F8lBdv5zuCvh/d7iu/pvvLBNuVNKm0F3RRW7bpHXkGad9
Qg5keI+LlGMWw7VOsBwJUcHZL0mD3q7UCwQm3tmnbOse46SZ8i82pxMssHf0+P1B
vGuR+Mu11kZ650GVIuKgCym0jAZVFp2N8plDougbZywChq3eWumtY/9TdHbwPs6R
yYXyna/i+HAtyor6+ayivBwNXIsa4NUNHhqYjcCuLx9C7lG1awGRynzKbOGPjuq+
tqBtBKNtG8dsAwDBVa835qN5M43gb29AXhUZs+EOtoSLrkqoTMshlF68QORwJux6
exdKzreE5HeTqBk9C2a4+K103mJ+UGyAfFaAI27qTataP1eHQEKwdJYLRkFGM5Eg
Jb4n91IW5JgOrowY6xJ6HWLx+Z8m3d4ema178l/oRXbhBE5n6qNMSq2BdYooR/yn
f2fyNMI26H/4ZkthOeDtAFmDIoTMFE3oxuBC6wQUJqv3H/3SV19V1nuJDmBjJdKn
XyF0c1ROFbwmXUxdqIyE2Dp0DiZpXbT+6UHVEleS3vOYnltgPXJK87Cpq7cs7iSy
o1H6qbpqsVur/3ZE0wVKfjvWyCJegI8nPN3f8cPfrskzAkwfm1cAx4EHVjay+U0X
5t6zAef8fALeWyAVxRLwUqMR5W6iImiNbzkSegK6MZRmoL7xEWhRn8RAwir9iyHj
bbSvwihbKOqRS+hRQ8Wgbhyzx8Fk+jHr+kVuwKFFVC6tSYOy6J/TUBQRer6CfKO3
wjqczeYcYIgoq/wmlCVDVkrDW8GO9jsNgQfA0R4psFxAEkrB9quIr27AioHrkmn9
/GYKqV3VeucOHoIo9Lqguf65SSzh7MGB61cU5v5O9y/FDnpWK/FrF8vUhxV6EftB
zIuJSbAwqm6FmjlGYzjTXJdjiWEMbWpHC+0v/KDtEQUzWAQHQg09kFd9dTTq2sk0
YdnOrLDzP0G7hCJQwpFwk15KVFEVplQEstFF6neocNji2deCCzbKkJ2Mi+q0Zfck
l2mjROAUG24/SPEX9xxUMo/409Mx3o2dLTMNwtjGLEDaVIxPHMt8jqovT1DNAw4F
8vRj6J+zQKlLqVc4oXh6bbyV9onv04HWmOirfLzN6S01i5ppU2p5QGwFf06E6gDR
s1jnu86eC9Awa6G5+FxQtnOjcpd7sgPfFEMWSBnq83NrWZHPRuoRmOsF0uRx2agO
K/xvAcEdtzaVy0Hujk+BXyBELs3SY5B7ner4aghjRHSdrEohrZ1qQOw2X+VGF9qd
OEMAIxXR03o/BXyUWCBQNHYafKxMqNylAisiNIbXxRsI8JfwtHSui8yRjeYSlEHk
r6i1zVPSD2qIodaKZEEik2ZDWazDObv6ci88BvJJLlY4uWVbtQ+zeLlcwIDlgHGY
fSAGZmGX3twz+ih0eX9ISc3M/erPmTNOP8f7Z3qJmfq54l5PCg8Pnxw7JNPx2Woi
1Jt4vyo10ucRoo5DYGsp8oR0a/Er3mVfXIMc/7QaXQCiJS1Ty17lamWdC5fMboOm
fe7SiKnQGYUAlY0w+iwxGwJish5bGJUws5LI0PNJA95tn0Z39vn+eWxboFOek+LZ
UjUSo4K1H3+h8btJ+vnZzggNSFYJ8MHemRaBhldd1Iywc7fehxyDU4ITY12Jgpjy
xln4dqXRPToBdf/5Bs0BoPRJhv/v48Vb9+beOSu6X9/FUGyMJ9F0s7gtN8c3H+Ps
cHvPj6bwssmjf3SEQ9il8e313TxtgCotCHdOgcLwEKM7ei5EPbrD8L6g656OWI1+
iXeMGvIf+2t8kBdDD+hL4UVK6WfpSfYHKW3Gu5HMfbYrGVU02Kc69uUJOIBLiYWA
+A10xruBs6VGON8hArlxnJ0sQwQ6rZ6dCTQKJDlfyqpBW5x1Fka/07D9Z6zJFSpx
/ojMJtEAMnVY7lbrFgEo8Qq75NVv2TUPFAgckyXllUADhWjcqHWbCVCiy2xaR/2y
Cd0wc71wi1x2sf2bPu5CyUXktjs/uQ93+KAgnPCw4ZAXpomqCYrEgYdlrK1M5CMn
0mYhdW7xlsdwT7Bh0jaa6SkQtGOGWyKQbQO7XqK3yn7kewC0XAzBq8o+gmyfTn+F
m7n+vCPbi1+OG0N7ajNNiinVTp73zMz4HoAA3Z07Xvc65qVCM5Hn3mldEmdODEiR
bAXMffdtd6T+90acgQN/XLwqWf/oWx2LNuiR7xhz2uHpWVkE5Y83ryScLlrg5vzP
4cBteuXIkerC4/L9TMjUS92F2ygRmnrpQR2/bzxdq7VjL1PNaFyRzHPsG6ASz38f
NvEXcdVcZyZTk+5XcncwsDKipKTu80a2jIZeMYgfDYD2+K4b4C4+qrv/8V9PCNgv
Af7jtjD5d108+C/Nq4jVLtOxokXsDLdgk5rENEwBP6/9TUjtorlmbhxnYzmNR8BR
Zv91rLZunEoP533k56Hbl+yNxk4CGwzMFuk+4RK+wuOHFys8GJZ7F5Odf0zMSQmF
Hjy7lKhtp8s7gnSr9aZVQ5JOt8MnaEKFzvnBsc7w1xdBGpl+LtoYIT+ELy5WF3n0
+KsCN3HP+qVNw1ecj9AQsN3Iv1yCIP9hNmNMpj1C1c8/9vXBegL04nOlZK+3FjwE
mVNBGjeQlu7IkqUFOAmo+bzZ5B9UBGOR+5RdtGb6Q/zBCKxM+pEc+LvMFMT1TnZ2
S4Bzx/mlyPXleJ6dJt3ZFCgIImVkpww3UCP1xlVTYmLjPSqZ3nPA+YCAvahPrq6O
gdMjlfY/x273PDU3c0u2gW4f84YAvBP+UeRRWdvNIf0DFx1M8VFH/K6VzkxKh5be
oICfF2hng6RFSm7CDSAtsO68CcmszrNDtNrCxZylaHfUyIdWzCjl8rtu7vEyqqSN
Zzhw2eOgV/CcimPDXWuC9BYTrRsSZo70YUj04JjTGqJlBV5LIR4MugLGAklvIdtR
hl8DCr6pyaAiNDjVMRWROSUYhbzbIZxDND2Pis83G5lPPUg1+lelIe4ZM2s5IOXu
o+wMmxYDlUvLRQDz+gdy1wyEu0LmZvKwZfDd04RHDQOTvhSvC6iN4+EGYagGG2Fb
PEfY/jclAQLFF6j6u9NXY/6W9Zc4Xddrxc6dWzfkcPtYeIlFecpyQ1/HrFKgzT3W
IgKWQi9+uuqkz+m3SvgkwpEIHcUdzDAbT1pAbQBpPa5EKeTDMK+Cbw4uJJWAbhyy
hSLfBkbEkpREjkaNUgdeJvfJ/NC+uf6Qdn2DdYtoy3QTiyRRv9dwD+hi6mXsc8mP
ABmZw5UnkWgy3qHG5OQJSxqJ7TzY2PvzvYsLVyp0fo9jEDpeeQ68G7+r/Vb79IVh
EOMkP+1blMM+jr5dz603Xe7nZwXwCpO5y8ANhK5I9oYz/qc2JFuZrbTbN2VHQL8C
+q8xfnnHnd3XDCsJLDFAivAWbk0uZL3rt+CpoVxGkzbFtD453AcxERWg2qFVGPrW
oxj77YQxIrYg1sYbZaisPzBBudIKksi/rELYZRmw7PQTAzaDVgw1T05KhoMmrtbS
5QRYupp7xQDg4pGCSXtqtDkks34WJkjghu+V+UiYyd1LhyDTHwck60kfJaCuGcKT
iJc4xDLPIWCcXml19seWzjCxz/C4GrZNuBcc9IHQTQK59T/ImA+I2aVYj3XVYfS/
fUPEP8z3GqBTmqtkjxdt7WgIzN0MyQ3LnvsDCf3eeBaJgJHlw5wufEUahQeIBqWh
UUsuNgHc+p0aQo87UivpRg6x5X3Sua0AhIf5i/kLxFFFYmCfpWJ1iZ9zmALDWiP6
mls8rcd7+emudE3uM9qt5deB5k28ekmyUh9Ek1OuGJ6RlFyC7JHLxlv/BMubdDEs
CAsycUbGP3MsZJzAFSrXrl5/LeTw0I8tuVwjGPqrQJoCrOL7quYqwGyxO4FsyCSR
bnkIPxHbL8cPwcQfeJrGoxtgpmRG89mqBk18eS5P0go0TPNqm+PPveFc8/a6FSOI
WykuFZ95nJLS3ebPzjQDQbVJqbQz3DAv6I1kOCZ55zK9PBmus5WL5N1EYjdiAktB
jqSmi5Iee3wsCtLlHXtRL8IAywD+PLLQ3N3HsNPOJa+PBaDWjsOguom5ymzc1JFs
x4AfeBT0Nsx9/6X76RzTtLI/XkTb/KQPZT+eufI0CuuYItJddeGG04tw3lyk7c1F
8NqU/htKHwG7oQSK75H84jefBwSl6Ns5rJFfRZoZT6RFO9EpoYpXdRT48UY5Ngxc
DOOAGuX9Qt4YUKbGzPgjj3EurPuyTiYrXXWdu1MUSYIz2KMYAr0MN5rjuFjvS8h+
EEUAdar00b5yyASORK/n5CfEInURHK7hLkP/sJ59Wj884W1fFhH/bc9o4+Yz2pE+
GwlK7ff08IhLVK4rla3F3fa7UyrqDLAva32Lq16K5vX9nJGv3ZJ5lTddUlEnDO/m
lfOpvi3AFd7dQswOvnc3D6GPt+/JAYWwk/GQ/RvKHaI7NI3Do4u9Oq2iegxMV8YX
iy0KUmEldKUiV1Xc8fiGK24p9x0SarUwUT6IIQb2ncqt6+7yt9Q0MIdcz6/3iLCF
lnKYorIzUvNvPL+YY/rTO4/W8huGtIMrZTCK9IOGPv2pt2FetoZz9aTXipZgoQcu
HTbT73t1X+omgf8nKUsCCucWFtOzKSfENn1MuxsWH7gCGzNXT1GbL1v3zjTwUu5p
XZAVIEP3vbhwa8BUqjqqLsc/ijJ3NM/yQDhaP1UYie7S7k2XXjJxMsq0/79pVU/c
MiR5Y+q24DrvjM6H2DRkUJt+UtuU/eEC3xHbLx0F0rpm+PQ3Qzd1GiJF5acYKD1h
7lZ5LUgNbNc9ZnP6hCJa7jeLPQThNVKFuB5FAP3tuEG9hGB5mqa1hpfTUsyGZBMa
kxaC6VQds/M8oaKnY3HUsMVIMtWj9uLu/+ItQ79piJpE5Ak7Pr4QNXixiBZwwUgq
7M32kRomhoTV+Wf/SshB/kTPpL1otmOmrpGDPgI/h2NoMZgcks71S9L2B89dPYMW
/4VWBh0ywQA+BfDwQJNWdVHW7kxhwLtz3qD0B/EzE3bUZNXnCYtJshI/a3UL5GBD
9gTF2wwA8l8aaNEljbql0YEJtcVKdx/VxChi+JY+hdz64p04MwU9g6SrkGtMBlL+
2DvZiTZ5uXXuVefapP5RdFFyqD1q3V3rtJuDfy+yairZzCUN+Mx/hUg7k+xkkgag
3CjD5leh0n3xDAhy3/719f2pwYYG6pE4feNRfQz0xNCMbD0vrvCfSqp8RyipDt1y
pM8jFjXETAs4JfV5oNnPpgM3oqJ0vKRr9desqHouMacANBkv8Qpzgs0No6YbjUmP
FzvxosPfn8bRnXJdPmG+4P5vcwjfQ4xJAkxif49WHaEEiPc+v4UlgqeZmUL5q39Y
nsaQZh24jJMY1uKwivkCNmqC5D/TOcVFCtoN+vpbEdfOsIR6CBsuwZhehcyCYT6n
STHvtoh/IrWzMfybYWfDrCd7b2tweGr5yjzt09fqyqoJB5Dzd/WEKO4ZDKisfl/a
poZjEnH8IOh6oDZB9aKdrXQsCaRpntegbVifN+VL0I5ZszdSeUyDpVRZPrgBJf6l
DuHeecXX/GecSQBO6Pab30Iq3kEB0yPo6j1sP56m1JPl0+g+UDasKnJCjKf1cAXU
B7Q6wPJY7PHm1Q8vXxfLtCMRXeLAl1o4iTrKpdS6KpFODHIXxGLiA+Fx7cFTcLsR
DBc6C02esIjYc7XKdGAsQPpb5PwRQECfjW+G6f3XHhFydypxCCIIfEEL4/XYX244
aMk7BNvSDDoHa8AT5ayKdQh0XNq5Ay06jLLHZDi6tsE5xaenH/iS8S4BSZxY9WaQ
oNn8WGHHCkcJEQ90g+lFLd5tNo2DMQc+piRM/+fZ6ncPMba04aXpxkueRczw9o0D
JiJaQTK1EkEoaRbWm8WAMUBOx++Wf3Ga3XLiok5F/1ImdDz/K+6p7LaAh7aiXbNS
QjPAW8uI6YJ1k7YO/uelBOvBBf5Bdzl/x58TJa8X/OadgLFCaC+7tETMiuKYLyJb
yhNvjBV2itRywpJ6ARlml4aRMe8JrGwlU8D1tP9qsk9gZUOaGfZVj3Fk1iPUJXbc
8FjZBMYdGT3qeqP7MUFXbGk0fXcl8aMAIWeu+v3UaMXvO1UPgGD9kis9rqFrU3qq
obOBHwUaJ093Otc1DuHn4Yu6M78qpLomS4VvgVdJukkT6fI93yFW3WcpPobt9/NB
ZmU9WwQijEk8II+sn0xqnE7t3GXgCW7dByIEx4vR9TQSKJHOFKHmGDqOEZnd8I6y
FfRaK0gQ5+44uUzm/sepZLZbZKMlUv4ykLTWx28S4UfenBh5cW31R+VdM3WBxu/F
bzatzwnZC6gGPjGvjdZ5pz4+U2P7KSja7QpF85n4WLzB0JckXenvpik46w/X9N7a
sPD6MPN1QgtIp43YMrnZyttTu2vgZs24RFjiveofkn6F3WPcVPuqPLw7rZaQWU7q
jHx1X8cL8X7WkXcFc/pUGXI/CN2ezKZJHrlqfIAv9mQ6yMBoIcsnsQ5p6XhRBuo7
wOQmpNK7yrDp2w8e+JzBrjnPxUAGepUojbJ5abE3GgOuAElxEz1xei8d1F9OmlJf
P/dBwMP0ZODNWsaF4Kzna0f9+YqLUnzYV1En+iEemQdGhdKHWgGsMi9Ml+CSUAGi
4pxuGjj7LqhPvqFETJHjAkE/By1biUXs2dgzIpk2lPV+nVY1xRkKhtxgHTclSuzc
iXRTDe7NFLWaluAVrZ+/xikm4WG6itTLGjUz5T/nj1+PVeY4ipXS4043D3po4rb1
b73jr2tlaWcydjTz2ERUf4sKYIKZ5w+L0FWSQ08eHKjz2oqgnsTO87OLSOydLs5t
d/K+bvSpxUq1Bavwml9jBwyTkXN/o60pwtHE8a21IUJjEVFh/VsFsBWpXiAEsOG/
/WEEa4wPL8KRMdgMHJKrxkPrc1rJVTUO9SbQx5oZMDpt4VHNoK17tlNk+89B5ram
VFIenrESuPgu/Gmga5ShgalaZug8TJ3roqPggpgdwQ/7vDIdSneTJmNMeFiWeNu7
KT4S2B55QPJDabHq5E+5P63m1Eb/eNA+Ht8jKHTa0zKrO4StcJcXo89hLIrLa2eN
rc5lhiTW4+PRcWsL/9jkwwHyKIuxKz0JHm5nwyg/ZHStPdfWOdtZo5jtmPRwNt80
Igtj6eLFaPsh0Y/otlkXrtH3572rPmSHUn4lzOCAfENAFrUJBXCSNrvX0PXa0SCw
GvQjkRcRbBqgiMdDnT5XM0JiIOgpBqtFMjobw+yjbAbEkp24LahAEUeddSPUZ9Dj
4SKpv4HZFoHfvseuFlOPJdRYipHusJNn+sDuAXWoEzR1zX53Bg6edGF/pMLluPUQ
8ccWo47r2Ksav4xbV1zaKFGgFxUS55kyt3N7/dHW5JmbugflCDhUwIem8rMxGug0
mxkw4dYDpCWhdf0IzGNJy3f9TMDYZki1qEVc3jeHKissLEBPkbqq+jNY3H2msQ54
va/kHuRqoZR8dDyyy43ezYLiVVOKB7B3PQvVa4HseSwvveLkpB5xGVPkaZXWuhCX
A7AqTCIRXBL6/XKdYZB9UAewoDXW4nPhBzg8ZlqgYFH6bwNh7Y1P/CcKV49nFujQ
HEYweyEnAa56Z1F7M60T/A0BoDOyOEF0+Zobhu/X1HfrSA0pPLFHu2FUThfuQpfw
LG29ZQoHVjFfYYfMGUQ9AD5MmKYuP9BMMdUFKSohfP4YY/nKSQELWg8SsugUPEXb
eeNOg/WjjHnQ5pZTYTAwXPhg6KORF8DlH7ctXleTJLp0gpmPgRReoM8Vbaq/6ffm
aUSyxzRJLxKndkUEsQ58zlDkYIGPebm3aJqt1KeFhp/Uq7ASx+XpCl+V81kA8oqW
QTagh6GfW0busasY0nxkzLZTJEZNdC2cWKv1DPWturiZtJAZCNlIXuLdJrYuqqpy
S8fDOU/kAJhAbYhwSl1BcYh/zWQ68vAvzdsVO30ts/WgmLYYI8gzJU0dHuRFo/se
Nvkq081AYuZe7lgdjNbOc9pGzJk9yvjElkfZNeFvbpHlc8yF6Kq64asewRqsSEtr
2UFYtW7sCnu/Y30jEI2tOe1Vflpo9QRoNO1pK5EKewUqwYRIBr99jed7ModgLGBg
/3L7GSmj+keZ5qwzMaD3xFcRNF/5HKk+HqWv3GiN4bKjKqYFZlrAQ7GxboEKLEAn
gbGY3Nw9M6DwVnmLOufcBJgLFgbaP6+1RDxRTt+0v0O2mYzueMJPKg99X6/yukJZ
3fjpUE/sYu4RaweenjInOqDEQGi8ZfCN5V25mXLWbKeuMAclbmTSQ+VMRPJXCrv3
pXnxZ7ZUG8KBEhJdco6gVTy2lEOYdF+36eOlUeD64y3UVvOOtEJvYrhWFBVRSfjg
J3sMOt5EuPWFBOtmDqglta8/XBYIgDm0mdU3LMqRHdPgaGigXQl2pYmAxm0ZL4dl
zoTtQukzy/4/iolsUmXpmX+PyL7eCLsB8mMX9kZXlkBjFCyj3wC5jmY3blYH7jl/
mafXaxnzpZc6mw2Pc30K4H5L+hBcVNyY3vlq00P4LJKCWgw1IURxpK0oXWSA2RM+
2JoQxDUWuYZH+X/3aOisMrgHII6fJFaa0OLXpg620iCmuWN+A8fymw/kytmSmYOB
MCGddxM9jm4QUkpOm1n4RRmcuVVg4oo56btqFx6FUkQ+uykHo+YssfNIVzkDp7MS
P0ljsABUuzxCAi382AOHcpVAnfj9phAwzTZf2uid09PWToWT5CdSkoYVgXmPqPiG
4k5PEkSTWV7PnrnlL1gBY/xjhPZCI6w1y+3W9zo1YrqGgXQ6bpXcVuPsq1kg5UP1
L6qT/TEkExi2WtGullFyRWRIlpoEALpt6fKOhSq+zJiTmR7IaqgYB+S/ZRVEY8J3
PdP4Glf0DVLLayTQadHEE59j0i07+PqfsBiMAyluV82DsQFmw4rKNys5LXoDwypu
zD+QSZnZhjkVDeQuoxNlwzsK6o5Y2wriIE23wYHInsX3u0g5UBnk3nJ1Wj4pcOJR
PHxzYWUiYNXfcXrUKubO/W4dkP0CPJxc28xrEoUouhQ9Y40B6WQZFRR0Qrn4wTim
TCVg2LVrYuzkvpNGxDIUhkSbq89HKO4m6KbdOjCdcHi1ARD+cT+l7BhKld9U2Ty2
M79zFy64Kj3e10pbKbN5Tm5p5xi3pvlmYjc3JmJ1dRJuc9+KFEsRU4WHIaZ4YSND
P1GCMrhR+o16zJwsr7NUvIvVsAXCGgCFb3AIhbOXIBsnhz6GfW0m50q7/x/KJW4n
b48ohAmbSoMR5w318jq9PWT8uh72tkgZz5PEaWeB5PjGC+uxG7Um4MKWBH7S3zi7
PT7U0KNt2AgMEgJpViZYztOIOBcZN7K/wwHxZEV9ekSuC2UCtzx+UA9q/PD3JCEu
su5yVBhh0CLKs/iOpI+ACG00Tryca+ii7sKEq8tYjlb+HmEpS8CWEgP48asX6O3f
gA3YJQ8U1ix20GfmkvYpagoWS7y8nS98lEf0xoMzVRuekPs55dgeNxayhvDShtRq
al1RqU0jMdHrKtEuUb1M10IBLjRMd4lWkoFFg6NEIB4B8IydAkpaEn3NA1uWRBOb
RIsjEuHM1FUsAVgKwofozWqBt0OQJ/cZQ19VbU4LIC8kjniJLbaUdS0sOAJV+iKW
8nrk9/0FlKqaQLJJEzC880hZ028ZSag0qgBAzGkJoa+5jWlv6tpogW5rNXhbKcjK
Iue0HH3w2Vsr+FgfRDj6J9PRArWMAwEPboCi0dYUHXXb2X/beRP5WrCUijwZqU2l
EhOoioygaZ5gTOH1vpPnCS6CqqL3+InsoUgVlhs/RvD8YkyDtCw4V6723HyKj8rY
vBbUAfmpd3INm4DZ5ZoWEUUJTfj+dtxkpacpp93CSSE0+H4CaZucwSO5AOcgOPf4
UeVTFru+ObrM7AcLK9hnoptWCVHrQAP73GaznbtvTTyb2KW/huxUejiNbwbwiNCQ
8ZgqD0hSk/8OHSeyu4eOf1tfWDbcw3UIkU0tkXkpQOd2jKMvcOlZ5LKNBmanTgqD
VhxZi56lCCbLuSyX95mAGkvJtem1Is/AkTE21xd0sBTWihCs/JwXjKCaB2J8EfQ6
NYf+0tk78PBzg5ftccRt1H7TWqsMONvI4gKOrxb0hybLfXCVYi9fK2YhuomTQX+d
dXwg/hMsTRNfXT1He0haTbHG+y4EWdBQOZPTTj9p8STvFGyKmJKIGafWnANCWvCF
ygWow70/3AOi0kSo4dPd6HaROd4f5j+DwZa5K3ar18wACk3B35oxgOoABVvY4Fv4
Yh2a/UpTbvA4TV2+oR3AokbUwTJXwN9kXIAu5YKS3l2ZNyOykz+sTUUCNH1U6B0u
J5cfV4xN9WDO0eiFTB5fHXCj7dCtcLr6jWGiRHIntpwO7VPW+JRNWw/N6/cBKakl
umjl4etSLICtT54SrEFPkyf6WUZuAHVJ9UxXhDwgKjH1NNlo4P9Xt7K5fZDZ4kAl
BaHxCuCx5iTvZ7SPy1Ti0s8FOvh6/V1sOPs5Pd9RHbMvytAD06ASJV17NeAafeIU
TCf0BSF04SminRTGr0/Y9kdktoeCrWxX8S75ZxBXsHCxJRgEwSw4c5SoiMEFAPze
nmpD9aPhi9q2Xm6HaUG6/FO33J0bpYVHl9IA0w+Qq7DD3fo1mshLxS++m38+CYFG
AGH9LnalU2JaXhsAxlAyI8W5tjF8ePPIDrmfmlW6yLZjIxp1Lw5CB7FFIT4+RGYW
YOAKOVRYqxEOe8ANB+agIjBqjiH2L7uftWKfMI1t+r+JWb4soTnEv+N8FauY5LhX
YUFtMu2Yjnl1aFJKuR07prWTLrXqhdQb+8kH0BH9UmKbGfRR8FF6w9KUtctfVyQS
fkoIV2b3MaQlVhh0j1r55T+7MXQFEqyjAn2AFwIog/sYxikdCfTgdD5yrJQg3den
vOc9VwOVo5KLU2g+BshMXmvQmyvVH60pZ1+IG647AkOk5NrdhRn2pyBLt/Y6HY+k
mMnSevGNwEWqwtUDoArcxb0W7qKh+I76O9o+dlqkii8aQyykY7rPSyfbLsBV/h1q
yAo1XZs60eZ4JeNhXCmlUH/gZSs6VEP4F5Y+ko9wbdBZa6XRyONTgpIHdlH9e3Wi
48ySGjossowCLgpO4OdGqT5LTtiVaULoSRSz324bsrvwa4Yk/wosbevizHFbMkzk
V0L/gNnX6Rxd5SZw7LlCOeViBbDu2X8nt/myYqmZkBlv7D4aNWDdemxcvdzMj/dZ
yI+sXsAR8QrEZouegETgMf/dWEFDzM9DJW9hVTKIiA/Cu3uv79PGlihL8s1nrvmD
0PojEVMnvC6keCPuMvlOAvslGJtnbmw7yiQVaNMWCMS/MbFe9jOAQ1lQak/IIfFp
M19hZvlmzsICYBmLSKKmKhywF26o9nnQrwX0p/EK/Ur7Oe3aaDSOaI5bcyBL5U4L
IdOtEe7WwPFdpreLGtRw5SgymhR90/uML34I6ChjP+aC/YgYdHgACxH1X6crQJ9s
KrVhU49rq2axo0lnkK9xOKFTmTldPI/BSPakb4I8mJOcqGHUk8mxfy9Fi879dBmA
Y+TcBUaFxuhp3blRY5Rx1bmBAHOgHPEfh4dH4d0HhhduLd86kvwAE3qOBl6JBXr1
Cj0ESMWFDuKnPTV2tJ1zrqBiMxvWr+0rK4Zob9TAD+fkS9jUs5Q996RxVTQYrdzq
4EZOsyKRDgRNY+SiRo168g0c6UeChDckKx1W4NheEN80JqONlXCJhccyCGQFvydu
Gv2BL8TI3IOFeeg5zixrq9XYg3/3pReo22hHOux56DpLU8yoxWarTCluOwB0YeKv
Ai9c6L/aQoqo6Bpd62Q/ahvRwoE88TGZnn7nmmyE5qIlj5ODyGsxBHyAnmF1LYEW
6m7573VOX+rCBvqu3x0Xuj04q27YaYQdoXjzCu0fBKBof5oUP3UP7c30hRUQS9e9
vEOI3ZezN64YwyQXSuQATIcA3YxVLu7tjM+fD2MMuWULgAjz+AjeaGeiAhSJnACD
Yp5Hdm60i5+tJDmqG0aPjLRCcsFpLJfwgKeGT2ap8QJ11PiNbDoiqXrz0xN+yYOY
czSz+AvV7tmQsBhpejJkqc0S6fY2mAWOVDzdhy3JYtFhDAKdYDakcC7+rWXdbvak
eoqV8RmuHe2hkeKgzhEjhNxUBPpDwqrWKEK/nMATXPNOfwvOQpEkb05FPeg/rpYT
vdNBaVO9KVqpeX84zVm355SAAKypvJWBWCMSivJZtiyMP4FlpQkDuPXZqtDKByBX
U9p0RLaMMiMtr+q9m47AtaqqNyXCMkNhupbVKxaA3FN9pQClgd1YA+vxGnoAKjqw
dmq7cwC+PUJguuPBcYk46unMxJUUVSJ+pk1B0C3POe9Frjvu1yLYXbAjwRmiD0oM
M/xvm+qZ2YLW6DRikDDZVOjqoWX36aqwYigJBqX44F+kiIAmdyUEDGVoqMGWWQ3Q
/+IrdZxAUg/acwupvuzSf/iDwODykivVtoO7D6b8l++wFzjlhcAX1FpDWiTGHDap
AnTxvXIosdEro2JnNS4uP2EsgPXsKhNAD6HC/OlO/BHB7l8RWeuFrJIR8tUF98V2
Fz2j2Lf8Mu2++Z39tRASbA8EJiAqsoPMVPd5HtpIxNPPCYbkQ+wCTSqeoglroa1x
Cx4qPwdSSgVTnyGZ1mBs2rcU3BjqulH+3sLkhwxrR8U/c/c49Ki8IMLiJNv2I0KM
Jk89aAbUjQSEbCJj2DVvc2lWSiBxItBe6tVBJCc9wXnP6sQT1+6mJShEyfaEPstF
+lPotL7BhaIxnb+LrvISVWReZMuGLtM6d4Uy+jKMBmy23DfTdPEJEf8dtcn+6a8O
WOej5PTY+v8r+38CcyIz3S+WyPcrtar/h2MwxqRLPl9p58lfCTCb8UAQJfAyDTDP
+orNqv/hLhw+/VCvLqmKMGxjtuf2LTezlmVWFtBRZLTeccePMZckBlIhMu/gWtAX
3RO+Av+d871TdMkMSAbVx0+ZXv+bfYpkuxfTvtn3kL5nqxW/6+mDTVFOu62ZPDqL
NPM4Ni2YiYm14mgp8iKmunTcSvF2p6f6pWIz8UAX7jSdeOMsuye4DU+piwBosNSl
RLwdzFt0gGhvUA2Is3rnre5CgnfYxZnOpXAi/ESzlJXKqf0AjoTGPLkHFOren3ET
ITZLS7w+ACp37d+/KxQ/vLLHlIfL68sVa2C1cSRKyMtUm8fZ0lEjIqF/4DiFD+jW
oMF4fX0HBC8jRtldLGgNYh4Db5xKDD9Pni1S4trUYlKFRalk6pkwAlUSXqz0vi95
GMnwY4AT8e6G/cBSptluDQRt2ORFGBCSlWXQl/NudekxjyFxR29TGO/4HkR0t9eg
YoYkKGlPLxOq9nezofHH2k4ZfF45B2cdillT1CR6EGqofiLfpOsN5NVW2DH3mzI6
PIEZWgLcFtA3cW7DI9rGSOYT/2CMC5hWj0TEYhhwNB/wO4LR+l4MY50u0kUKlhgK
iLLU8b2pbPy3OYEa/qKwsEJYnx+CzfKDfGrTppGCHj639kLvivK66RC2mdCsYtyF
D2Y5WOYRBsIV3kgfkgQ8ughf0PBKRAytpV8oRsaZzmtLt3TcOtO5rBqXJWBdQ7RE
nzrIFbfpBaOt/7kS2Ggc3Gcp4sg9mC9uyQAxbcGQZ+fl7bgVtM9NGgw5ccFxoNH4
gwx2EHP1RE68VS0esImyjA0OVy0RotBXi2vS5mhaZkwM+6M5DRSvldi5yw28L6Sy
hUmcmLtAr5622PXT1TslyyERRF+xkk34gAnig3nAcDGHMA/hI/SVJ9c4QndQMTal
QcnSgu2IMsBgbKaioTi9QlxzWznbk0m726bOnTYDl9RWC4MN7Z0Sjm5BQk45GKse
Q6bXTGmIIthjg/68jgnmQJeFshM3ke+QYcttsx7KvSrEvA/41DI+AoBqBEhZaoDS
foguakImqBf0s7OVy7/YNkRXlftGcGoKKDeooBVxOruBtjpskCIzOHP74C5v3ByD
WJt/+kI156wt4T4nuS4Gq38KWDrHG3oQ6lnOGWk2OfucrLVyUyMnQ+vhgj5xdhsV
biuCOnmlOTHuM3XTkPw3+00lOLuIcySl3IkKm1LVIoyBkHzHU9z7uQHEZB+CS3hX
WiPtPQidiUbGfSiw0S48CCVzZ152sDp7rdkobcg8HgN3xUAfb1G9uUXf188Yjnuv
mTsk1YabrGgJWyFKszkXH0jk88tQ8tp8GVShpEWR9k9fowVgSBsD8k2vShJHbHB+
q1bnWO2kLCyp0y0BmwNuyuZ9sF47y9BV+iRPhVW0ze+5hfz27AnS9j9HC/+WV4tY
ETmKYdwn+SZdp4DdRI22PUiRPIh/ut03CetfhQJ8sPFW3RSL9V/OJN+tvWv1gNWu
K0AnlF0JHw5riY7mRRlpjWqc1GUXQMjMjk+ZlPqeaUXhuGJt+mai0+k/f0Se8TmU
7Jekxikm3sUhaJFbtAgp4fxOJOcUGKBEE2KAFFi2G5PfEHwSBL+43Bf89UfLg48J
ENWhGBzALYXcjb615RBiz6QHgNqdfQw4ofUCbhFbdvlq0K18RyQgHnYQZ9y7jMet
bYv7warw9PMDOMEUj8Ng8+WG5C8Tjy86UUn9ZLWMrO72lUHYzlDabFiCcvt8evXK
j6p1sF00E2HjoMfroNMJ87QKeDFZTQtUj8+kmNkSjOJxENtP3pIo7r/xrdQnSyn8
YhWOULslBZg0nYa0mOM+isIf7xtvJFPUyCSsPxIY8y5dtEsNqK9ydpz1Ixgv8JHY
uZmBXsbbghHb1AqVfNDFB3ly2t5OoVfjqXy6VcPmMbsuTDcd+igu+Mr7h775uWgW
Cb2LIeYFG5jIPryX4LXSo1WiX7ehoxM1D8JDxjAyTfJtFmifQjqoHlXuH4rP7Uy0
8xwixEsi9bR6XuWfFQENwB7ZlhgYqhVMvTmDSaEelPpbbED3kV2L1tPRAMnv31GT
y5jbsS4iAiFnTGSe4Uk3ptYsa4Wx4WyTKNew+ZTketWXgqj/ZJ+V5rsDTojd38vg
SSOVvVq9wS69aQcrci5DeXKoptQo3MiX8cQZ5KCveZ4lsXY0u/FJ/Si2Vgzyj/sJ
iMuoiwG5nb0v6+NXnqOGOEYeBS50ejPpSaT6Tp79ecrjO8LekYBvKpHvhLcVfjlt
A4AjWAv4N3tQF9U1NplEMP2ObBhT0Qlb3d9cLvd79NkB0zWMiOqHHhF53vEuyzPC
SQxf7BJlZWvbS/o2fJ2Y9iyX86GMiCrvvzX4rCDMAonplHDTapoNZuiP5ro/Mo5I
IjreOGqxA48IBOUfuvozAZxICkdom8ZtaB/juRKPo7xspJDSlfb5ev1nxHgj3EKe
bW+W0no6k8aZFVlCPQnErP8S0aNZZrkxNPe9iUP+Kfya1mrmTZjyFwP7s/olsNtO
Ad9jl1UR6LCK4HUdSUjCGD81Ay5PcHCE7otWU4XS/+0PzWPGg+nDWzJazDXcA40j
7oYzOTezWnNrhVKyxFObXmLl4j21aHGZj77i3P/0sKdl3LJcISJ+Klq1I4omlu+R
kS8GfycYN2LSmCLA2sko0lkiGui7FfjRuYUGeZkphYBPoQxQiW757mQqeL5ZEw3/
jxVrRtzeYQ5YdLtHFOtxXc9gNtD0l5kFDPQgMKJHzl0QQyE1ASoNl5qaUcfsT13+
TzeHpdJqXPGQgQ9qEi6dPUKnbvXym8mS0CJeapdAe/WSwv7SC81unFWex6+g03cH
xodLGek96Klb7sqg9D6rWBrwMRKRBsufJcp3ckIshMDvPSFPMs49UMM/yP//adXF
6pL6+Z/KIgarvs0Ih2a9sPHNTfvvSNmwpCN5uZcCV6A+MgpzBFV28TGAg7rt0ipf
jOcWpf2EaH8hGW/TBvmQjDHdlfzh93PhRS7TZgH5ZOhD1IJzc0xdbjhsrfudaeba
nqbzL6Tr79NA5VwejP8f7BP8OAbiF6SSKbMDEFso0VdJhvlGvDu+LWPQxPu6xMsF
e90MTWhQPurMgteIpke3OH7+kqHgDl726oFWNx4jJ4xJ0Aui7n2HeCyiabrYwFVD
TeLwbkxmiXdfYJWl5i2MhWWqTmXm8NLyV903vMB4iK7fPUBA2exNZ7sFE1Kf9cEN
sv02+SXoJwLJbpMAMiHfEPLIRir35Kt6mDpDnj/eskHF5n+y8h3lAkT1xzIeNyhU
CCMl2ZGop4WvSZ10vOPhzSAKADotGRmxruB9nKxQKZ15wKd3EBVK8XjBNjC3yr7e
kJMsWrBazfDOYOuOLyJRQCBw5paDp8/tdi1wwXem7xj9blD8KuCly1j2g5yaBVFs
53Gk3OYymtmasXigFcETpYMG1LHAAfMZmm77gFYfkxDg/hUh+wkz4n7ghw5Y8IW5
BSC7L6xflq3SB1W6CepEpV9H5m1cx0pGODIfWfCe4QVHvClPBktJISIgLXvQ11gm
VlXUmBYPt46P78T3QF+9DJecMOMyFkSa5BSuL/yoxQj1tyVmDMM9hg5fnn9PZU74
UwDnXm1hbyOHEl3eEO0QTWo60PZnM57X7m/ANh5m9PsWKmZQH+GaWpSNRw6XUvo/
9IhOIM/Nrh/xJJJOozXseD1myw4o6pOJlqlcfYh4Xmop/lLHP2A2JRPJWnBHBV1n
SNT0XoZVpcn0DFsGSx/A7YjdQPeC4+OSecuDy9LCwipkQTGY10scMxX8ZJ5Cr4C1
2bEWov7UnfNLyjNZFnMoo/gwO5M0BhX4mfvVgRHT9C/KXkEAwpr5ATJfxDh4F7ud
smhpyB8myWXVtA1O1pT31o1KbqAkmlH/eC/+dSFRQnb+GRzc8LAkuQbNVtKYZ1Zz
sTNSHj3d9/ZaXdj3RbaPdJYuivjkX2OXN3HjxkUGKjsLdlmkFXTW7GvnwM3ebgEZ
Vno1Pe7t7w4aC6FhNQaDI6AzZQ/kdP+lNViiuaqm0RHHK40lEromD4Q9yYKccFNI
RJhgm618pgbxJNpfxfF3VU6cSzEQHBghXmxxtmoWwLQtjD/ZuWFFvEGxz/iR6sLW
BO/NaRHnr0i6VZMW8y/ZtLlFCS0Kk5JEaYS1QXzlTr3y0yd4Lq+7/ofeKcr8ntUJ
ZkI/X1fxSrjXKUmrzwpYBHMopUlV7imgiFkg/O4ZfqnHThjcHoPcNFcGf+XwLkUV
FcEfQw9+DzBZjCyp+4Uc5K8Wwy6H9qk/S704WB5hSOQoKmPQhohXn/4fVzcZWL7R
UWMjgWq1mfmqyZmaADHlDQgy5lS67UuZCoH8vPkD6Ez4UJZNrp4Or7w4cjmVucWH
NtmdWeu27qIc+lOKkcOz017WJLcUmsyAkxnPjcCvGyCpGpqhSJEECJaznjfGgGr4
P1U+FnejzKnNm0r/Vzfz2JpCy2cisxIL7lnq4VV8vP8ReUzlroWr1sneliz2MTT2
GNvsZUltnxCkDkSQC2cY0DWjWv69adXjxI/qhjtCnL+9eCFAWFjn8E7P4brfPNSU
0sDRlgfjkeck/tZWWHm36sOmyrMXLnsTM/AWby2jMfLroa/U3FUnenDxDkRwO6VJ
6RZku3arnVfsJwWTErl4J8rUBCw+ev8SyLMVflTq260oO5npLmc0T6hetFc9/CwH
HnDGx6hmO/o2GwP0+3JWkxyb73l4d16bE6BVfF69jj4PU3Q7aHcgKC0Zs+OKTEY8
aqAmvl2RN255SM53sTePTZ+OH1wGuoIngnHLxoNVIRDI0u9y178lq/waOG2zUQD4
WsQUHd2w/EvMzelFztR+DhOBtnrbnSIWbu3MDzOEzIu6jJRZTe7kLv7Dnf74YxIU
vkfqM94WGwJXIONSz+T6xgP+9F8VlIOsDZ8zhH8AclDdoLxvtv6MBRgE9WImoyAx
Qy+6hrHIV1JNmAtmscM7JOQBKqZrpPDaeumAjOHgw7uM1vobX08TAqJQCGl9P/Ks
MTymDzndX8aF5NwIM6MZuJz62tlIvC/X+0u2HJb8DR8ZyzCch8oNz9FT8MuSwXqq
A85Qp/cjBLbYb/B8ZHagyluFdp6j4TuZGmzTQfhSEiK8iezjgoc1XGWA4x4rZn7N
tXMXuA0VnFgpEeOFygUL3866KY3n+9O5tiStr2muv4W3rrGuGYcsfn7I4r+LY3R3
hZOe641hMCtY8CKa/VXO9RRjRCZwXtFgPFgDfyIrx9FikXkisduqYG6mecR7w8Ny
C1GP7YW0D6LQJqoyFEC0WN1rcVqyN48/UvyrrP1qrio+TJZ9wFhTm8DdtL3DPqGb
P9HOjSXz8WgJZ9jI0vmVP1zFpqDdoDVPSStzlmJFpLRkFpzFiZZLr2zQxmYoOKgi
BjVMsC4xKuRWg7Q0XdSxESp3TQDfY1QNlu2NbChqgK7rcdWH15RUalQgIfDPgd7X
A/tYyg1P1LhRCRNKrnr5IjP6dPpVMw4uPMLYs+95V/rrhodBTxf8MXoBSrD2E2G0
BxbZ6qBcubL/TMtM2tlFddvodGtA+JbWIpQ+wH1ilsc9pSvk5bbMcggGWRfEp60C
XglbQBvi41FQOrpBm51JTN+nFYtXjZ84Q7vQE4sAdfFhG4rdA+Vz95s2ry4AGmKA
5EJ5wZUz6l9jwBlWVbWkUI3c0em8hTP+uLpcDCKS2IrSRjUmeMmbFooQIWXypDGv
ZaflXD7p/iNB2VSQLprTQziRWs1G1+ohQ/BuPrmETGimvatWCiMTCuDGeEOIDMcc
+MUMBmOc7twusbkaCUYTz1VWRwdCgAe7Vf0hPtQU6MONmBY3a1k2RvBILzdMnqeM
G4llcsGu72IN/kmB7WeTkyh54mnd6jnIG1SOvCWqMmf20DGF/q6IIO4FHP2aL+OP
yfk3y5kPzVKJGp7XGklXfxG7k2lU0550MBm2BTaSEqah8Oy0i76ygaBIPUvWsYXt
XvZMpsPS3GRH2dKUvsv6Y94/uvDI88oPOxjUlJKTWhKJwGcXhWrO1ueVTqPbDrle
yh1AUcP55BPhbDZsALStFvVJGwoucLilypXqD4UtWKgF06LKkYi4BI3gRWmvM0j/
xzA8uI268gWKwvDUOtJ9AEazK+aE49ZS/fcIqDJL5aqnrnVGg8KOgx57hFIRQUvS
d2f077McXK8L+2vvGbTk/3JrHSrvPWmaNquryF2kIVncV8JVtlabmrMf23QGcEzq
R8M15fCglqbhVc9bD4wpUNVvvDpy6whp2z+1Tc76gPdM+oZJx7J4+d0LDdrdFJiV
9jOi+UsVUit+vMQ2jyCr5W+S2V+baITePYodp7Cv9mBeTdVzeNyuBIjmaARRtr0o
r/TL6H13UAfGAgYptdjmZPz5ImmcuL94Bbmyppz+LUo8utKf5WMqrDeKGSaFC15F
CYlEb14juiaMxoueACt9N26ONd7q+vPlc7x6AuKQHohvSRUTTNuXIXcNgOf0uoTz
X49KOdDV5/k0IkrD6tvZU/V8wB4HIqLiFvOEV0zNrIMsnjah+R2Z5C4WeW9pGlri
oo4kCpR1Lk6rdQLTBn4Sr5Ddb+7tZZjBn9PVHr4lnMYSx7tDDmhaDUTTc/RuccIW
sXLoYp6xP4nXqFc1TRV/dq9Dl91aaj65dc6CIR9dd02hxZEWviLf1OUQJ9nV1i3f
ZPraCctAdFShRcadhIyvc0nAFQbJ9JMv3OcYq01XI6fBWusrRTt37XRl/CXlwQz2
2jRbfPv8IBLafxxvZ79tI7MpP5JNe+mfNu70A2LRty8qyC+w8+5P/6Rs/wMWLMZL
TYdzAvO6g92tnHnl6i40QbSYRhy4ehe0H29xJAfdRnrI5aOAsXH2KGEc9oH93Hnv
JaOtnNnI+UAUDCYT3cGXOv1Hk7Wf+xVMi0k4aBoNmba1IO0qM0apmY4VlomuvoJh
gO/IcKBnM02c+i1B0x1cP6SYI5D8iwIBS/8ckvHciRKQARAd5DFZaaKxFYeNB12Z
Ud97K2H2RoDKtEc/ML4CguNA5JgEq4vK+FbKAXK861NL1+sK+fSOY1Ac/4QK26Ix
9lrBBE/D6Y7jpoO9LBUJ7tKcakm5zNihNM/sNRwJO0yCDzPZuqiFUV7aPi5RUHgb
3W5g6VvQ5PCoOUsfqcs/aleLSX7bGF1dileM3qzSECfJXveB1Fqoo1hJArqa+Q3F
4RMgy3HNoB0eFVhSXuHw1TJt5nzbq6lA8EOyZYdq7syEgnlj8F0kfwSsRhtMicaA
liH/bAEztVX73hAB9QgjLD6nOjisOXFp7lvKfV7fp+HYcJGIA5JD11CK0x3kAZ9x
EiZLEXqSjD0BcRWAFhev2vRLZKPtLOKqOwp+5cYtTaUTDTI8asGL8nOIe3GQsAfh
jRPX0TjA5cZYD0SAeKK5erZJVaqVAroHcr9crPBxW1+V1eoAXLDttocBJ0Ptd0rX
Jj+swzCvwV7V8ySamZZx6QQXIK6fIhNW4AUPmPnd5gjxLaq9w8Q6bwsDgCww+CtU
S6JPsYA/grAIQbhISkUzHRh+rWyAF4KwzJcW7jZdRIOkrgSQgxIWJ3HtFWnFJIc9
5O76x1rVV3fg28Ok6el2C7+yG+jp+fuT/otH03oGtjuzVUzOSKBUBkXZajYk+CwL
7Kt4xtaLppVoRUekBlykLRpBcjP/UUCtMAedNMcOuEPDhcvJdjjnY86aITneZT+z
XqpQZjLbGPN4qSPIbs1pb5fDz5B69VvxST4IeRtHwaoU7pbj7y9+yPkKDb673cUf
BY9ErD5Eq1vnQ9Jpxd2EDWfk0pQc5M7q7mn/Xkr4lU1d1U/P4iXRcjsiFqRYvhU3
AKTQsnPEAYsTgStGFxK5eb++cm6l0aRBGdP+nYd4nt+QazVerjYCFOigUKbxmJDQ
Nu1krFPTf4kY6YvjQyJ66xwT26705TGS2DzWpQw0Knt3MC3iPRzn0vgrpUKQJsxV
Xv/3dQCSoF5cApa3ng9ZQ+sf90jJu5sg7iNKYNpcqHeiWShb+j+hsTJJ1HJFuJL0
pSq/cRG0sX5Du6JD3OeWnDJplp619o4XBGQrAFPc1z+CExzVo4j3GNBtA29uvRKB
10AL7iEjoFbG9M48fQhGdd919r/tVTDH4oJwUfCSdSeq+8cKB8qnKI0vjyhf0eiP
AzSkxk5pIMUB6z2sZFGlHwcUsZIDVmPann98QS6n/G8bhssx2EumN5v7YNYeA9N5
zEdUIfalhYeNFCq4bJqUrfVdruJFYLHU4O2gGloJQcmeWxHeyjU6z4yFA2EWuojR
rBqE2Scr0UZw+gfdOOW9kRdRFcYoEju2oyEXP3QLahK80ZkArcDztkP8Zy2xYvOw
Gm0k2A1I/X6RpsVGbHNb2Osi7Gq0sL206blexd+vqgnSKHmm4fd4oAPC1hiqJzKR
cz4U1RMlsmMPG6c6sVRx1Rztvv+MAVEXzxpaL/2jBqQETJ/lPTDZVND/3krR6iwC
DLDSrC5rrTfdEgnHAcdcjvB03Cq3axgQxiOy6vNBnI5hMjl1iAN84rH7oAj0nT3U
YWTdt7uR8xFPCl1Ys/vT7czwo7U0sELiDSQcsjFDurod9Z1C9r3dc85p0kZM3ql5
W+3P6JU9HO+7NwPYriJrQuZE77iWvuzn2PRYLw+mJqha45OE/4u62i7I/X4sfU8a
5MWUUihbACc8I9W9TeC1CPNyMF4lo6VUyje2GHdXnjerV/OrgQPgDHjaM3atheoP
oJ4XMv8pP39OdsZkf+WXaCKWPk5FU2ylPALdShlwwgmgKS8sqTmB0N/M5SdQs+wH
upEVk8BxYRfvTJ7brDNFrGjloDQxzjT4a6locw1fXihuCeT91uNbVO2hgtxegCdT
XBkxtFigOmxfjt80YP4oiCRQlVdPIZ3hn5hPyrrBHcosBFpXgCaZRddbEEI99+nB
EWC67INkYzOSze15ZsPUKAn3aznPAB2I2gxEQu3uBOT/nJkQGzwIEf0Eag3timXt
rl85YfERMOUODD9MPdb/1uMue8PTn7KTt6btg77uKyXey6fUeP4gV0M2z30KdODg
HSmIwsbNEm4eQ9L+5utTfZ1iTKpJy7mCWmfFsW3BBWSFakZAhtKvJDoPgqoehzyV
uTIfqle6UfNeZGiGS5YNUccFUzTq4/CjeKB0uR7BgEnddeWRjIC9gURyEhyLB7Nc
YzmxXEL/Yn/8Cbu3az+s7FRfokhqtbQg3jFQrHGNu/W4YMrkSSALsIIs/49LfKfz
aFCLH6z7D8dpv6UCQnRiQ+RmLCNQb/hbW5Q+kcjMr0wOmgQYbsQ94zUqFhwx2/SA
tevfyHVn5yDeRPhwDna6a9C9x3wpCB4joUyv5dOekoUPdKMswqRpojYCGxZ5TMsI
gXhMAQEJOoSzfvRRcw6FoWz9K43FeoZLFHI+axcQALI+R35I0PZKK1BgJYZMbF52
8f+z2P8dIR2/1qjmajASm2tIdteh/MzC3Wz4Bo4xVpOhlv6h7x2oDgphQ/2VBGdy
6fKZOtYpkrLpQxSKrsEyep2cSd6n58Z2n8bCGdOITKrLc64F+HdzP5Qafs0+fOZ7
g82JJNd5cXnEfEotBreIamQDJmt4RsgbH0fQNx3RqSNmxueldkQFWkcDtt67YdZV
pD/87WsXryQ4+CiPEyjrjgwDXLN5XtqLhZ/mt883Cg4KvLFR/X9g4lIwfrlnY8FB
/8U+m3y/D0oV0xcMImOWBR/HJ97qjgJBkDEXu8ptbR9KDGUM72Z0MPMdf+gRmWlm
N6R0dOlCgYB/dBCPgOZYT2Z6pLi1/Vi1AVBM86ut3cA9Dx7ZcRnN3RGPax+BBhOV
IYDEdAymE7CHbBR/JDxStQwqwLFMgzZBFD/F1NtymS9LKtRqtyIx8qlvX9A6HjAh
utCf4/EPqq7ye2t6s6LJQ68SpTQxeSkYbhs2vDoMqcEAaOc+EFL1WzReaTM1J/UL
l01JBuuoBlf8HtvFWA3vgfXq4eZUctYHXlB+4EKVzgdowLNzTSrDGNW1ZBAh0a6m
r+cJRdHpk6z3ISxxtFFlUa133LmKowlw0lQCVwE94Po1DtbCMwRp0TYZrgW1wcBE
1zsRGqc0MTMIJzZoBqkS9SACDH0HOBhTIHhouVbso134JFThZW29no5Gf8cCgUID
IXFqYw7slWj4eWLY465daIWYpBEMP8NufFqSA2GqnjUyX4IuOKxBYsSg2EDuFHJ2
w/L8J0WTlsRX+3+mG1IhefSgV0vqRP1a5EjqRbBbEn0RC60jljkMMhCIj/v8SzJV
KOg2QB5XzOGGdBzKO/RxyB7irVOsKfGcieDFszhgiwKqmuPUI8Ea5k+K+cdjWPDT
sm5kI1QVdS6wPHhcLUu44ppWWy64jFZuNIdFPJ7h0lKDGU6wiqI7ndw+EN9buOPf
4Hm0PnT9FTUYH51m24KOzIl3nifg21fMJQ5vrhgz8bQ1By/CPCyorb5OCtMDoc37
cqaGfxml1UsWw/8PugtFShEsS3QDJRJedKgZzdqGdCAiLoezCC8FLd4LJZqZNAH9
kohVofUK7kwPB6aRI0o6X26Zqg2yv+H1gQVYnAO2zFfqA6yd4jpnFz3IJttYgwl2
uAX1HAGnj5222v1CQM288g8DZdvcuTwvTc4Da7fhZELPvjwsSLx4LmW+tmE3/mwD
00VOW20XpZqyyDT9+RqS71sYSqr7NpN+KzhyPL6FwV1eULPWIpCIs6LvLZZPmB/A
FeAzjfcGry9HTYXTnNMWBQb2MdZXkop9wuXgUYmHFROgT7ZfDH3xLKd89LiG80JC
azGSs0cXZHJ4QhlErhVFTOhxffxOL/ZzyWkjoE3exEL4ZDycEWveFx5vJt0imxg4
V1RJ+dOFzxJ8psC3dEOUTxTlyQD3RRHlM935/Ff5O1YQRK8daYnvfokcsuTMlVoU
Fo+M8ie7ajyYVV0PtbdaXk8rUFJyj8CiQEqepPLKwdnbbffAoIQAvUxCnvsYSHCC
oZH/K46UFXdMRPie5iin9JXJVvlM4nVuspC8cSs0JJG0vVfeAnz2YRdayH+LUpPC
Lor66NWwpZq6nnqLY0ZoTAI919fvBPXoyjg/xjysmpjA0irf10aN8XBwr0XdAOhq
Y1VA/6/qs/kqQj0NmGssblrJfgnRNn8vn6yuryGR8BvnkNTFSOeJbZq8aA5IMpxx
TRmfOjfLpas/CHDRJVJ2c2vnhJodarjrsFbxh71K4JvY7hDmucLu+Tf8PXGih/gr
5lPMG0kl3wrva5NUHslt69CiwY9ATJI8Wxs7itonSm45ZiTSScxXr165plBd/NX7
sXolbPz71DVvoBsl+SCDXS8dRZNqAQbnsgSRfa/u2B041YaaRWN3EN1T1S1NTac4
rijAJy9TZYS1WgxNwx1ruLPlRZY5E5V4k5FniBLg5MCI12ANhm0XG95BxJH65R9w
+tSGTp+zQ4dewA3lnqxaClbJ6feLKp+EqtAmH/N0r2XqzkU8B9QK74BoZxReV88V
gydYAIgkN4lDm+wCD70CvrchknKgE7YrtymKlD1xajW9iC9tTQLOtLFW0QnWTs+9
d3Ln3L1me4IbIO2D6+SgcpQULJmYuiDIEx/+wRqf6ByLvwg77fLuvPWr0x1AiBQ4
wgCfoJbkYxOOK0wEeuYE8Qjg9qQ70usmec2akyCxLLAcgg5q2jSBd9Ggp2aa73WC
dmSyIlEPAbBfTNPfNtfZz1cbKMJFZ4MJ/59mYZTjfZbdfopPg83DW+lElR/pDLO9
iwTcCsPW8DdPAwAymZnFwKLcQc80Y8Vh6IzVhdZvRCdcwL/bfxr+Rf+mrMwOa392
UwXsCdaUgBNAuwx8hwLs7B6gzGywqmGu1erLEUeaqUkoQ5tSarP02vwXBRVqXT6h
duI4ADs6JIsP+TlK6ZO8ZGPIbhaCJzDlKYyGQ6BZRpA6SAz0FaKZA9YRa/rA7ydl
ied4Csb4Emx9YiOfvJZOKihrLPcfLUCeHJtvOxKXHVctq9pvXStIp/TdGAlX06NI
mLVBJTGgfwrgYsRkx2amvIqy3BPX7pcWS5bhoSyMygTdFcDWvaSZz/tmnNbELULK
aRbpx+rcq72JRL6RjpAZUgpRgv96lIKQ8kqrS2Et4dXzeIPBKMoE3Fo0oDZ4qws7
A+4Va0CtA6GWSC6fEfCtK8wt07Axs6PEiB7lT55OPzxborGChWeeCXccyguNG0yq
oEzU1ydD0aI7ui/nFOhd+PPOCZrutPhNVVRc9h+xwl6V0wtVzCyGcPAvTsDAICv0
6YeYB6bCd8505RKVjKYhGcnkEzBu2DbKKVBMlhYI/qMErdD76ZAVbBJl8frlebMK
dTPCFN8s7Eo80w4ZnS7LV2Bw7nWvNM6Kc3/0pDm8Kp3y3uDdC4xp4SZhXyw4nai6
BMs6rYTkrWV1MEs56Uq4/fCIdusL4ULXuarAZYE7mAAgx667INqIbwHCaUPObiQ4
ldo0x5Zm6Ogt1vHPUXL8GmLhrSkFPdjZCTgFwr0AQfSX3ndPtgOwuR740BLSsjZe
arKh+zzmfK0reEXTUW8gSLVJqdHJYQbX7mYhaaRd13IOTyqJ07DkI0dGnBDKObK3
5ISApCRZU+KPH0SQ68UTlhLVJo4h4D/7eajrU2HwWtt6FgvneW6xZbmgm2FndT3P
QqTOxgu49GKxMh7SqWXJNhH8FBdsBgniGHpjXBjFzbNi4TQ2Ugx1SGk8JFKuQqKz
YPQ93wW+4tncYParlBGkC130kozuILKjid8/ghrpgXzP9bUl7oMdtK2HCWD7ru0V
VE6sNoaI9kAJDc521hzoq8YMy4vTfjaVxCUrrRbcHJetyioMi3Kh+Xa2UoMdr5Lx
0yAkGNJ0xnNXOKHE4hmfySDm2tpnmJmMPzA0fE4VIs6WhHyb8/nppdIq0GRzcdiT
nsKzS3jcifPYnF8wKX6nvIaUlOwPJgLNzmxOaMw57BN6uy8FvWJ4hc0hMn+jN6wi
lcW4dAcDoCwEIT9XK8ihtz11TKTgC3I9qfjxxefZ7E/QXIkhS9Oicef3WJwccyDz
5VI5IulnMGXEu1DHIJJRk2YDfNURguMBsP3PAGhwiyzeLo/DN61HEfDWq6f2utQ2
YwrMYps8jzEmOVtKKINz1DVnir360xjasgO0mAzmXxiBKzNwA4FMWz+KXtVca4nk
RaZgJq2akNaDhMENpUUi2Htz/3Xybh23VSEkTpi7wG3QT4Oy7r1S5HF+gB8/1ygu
nfFW3jhaWzaLkNWUYoF/ERPNQcpC3qvBrR3xcO0TYDDz/fpzLKIhckUO1YhaitgQ
RVvHIUZff5w0z3DeVV1YhE/HdGhgWJ4hAJBqNhle/nmRcyVYucbC7COaFGlRGyJF
7iwWquY0KUx0tREu7Fsj4bZjnr4aQsYFujpWt4C4M+CLPb0OaMfqNNi75wn2rqzO
6rTMH5Nbsq6nSPCdLyMsMcNJbJka/QVKvWqtn6/Ha+tco3BMs9uaUFSc/HwSNeM0
HUccjzdpFlKEyAUYACnQC+z0hqx2LUpalzF6QB2KJ7Qg7+rttlPL0TtmFeV5Acnj
/8oR4o8i4iYPKxHHxLKFuUictKot/G4jlA7hTFY8hgTF46pNOsgAO6M5hlbRjiGG
cQ4nm0GSKgfogi5pa+hDifu6gT6erddsMuM9xYqmrBQf0QXWqsiEcX7decAEHqov
pxZboR1I8X3/Kl5ei8jDaLEjLEycwDncX0PRRE8Wxj4gSErz0bY+TIzRimi/QJVm
sNbnrrdXhXiBQcbfkl8b3IKRZbeC1LKZXubqwmdPBOaZUSMF939bDuQpA2Pelcwa
gKpAzccR90WUMxreWyA3NQMiAuvmSW7ndVbTZV/cXAzcdS4hF/YZ+uI51dcDViTw
O1tEgSSyqkGzW03YlViv52/9vmycgWRy+JkFkBOGKdH8MnQ0fMoh5kSIhFTkGt8Z
89tp5FBHi5F330674xHMTde5i1nGkQ2IKj+cmS9q4dB3WwD+HtoRtcFF4+vHk/Wf
WLhN2nSS7dhz/Hy9OHGqTuiHngbBgpCDLaQ9JzsfecaaOznjouBi/Q5aURPNpt+j
gRdtH+ctHW1IpIjinjlGgj8troyiAEWER3STjVwK5AdBVOkkdp6f5eTVVrgACYnv
8wAl73J1LhNrtaFzF2LdSiHE+qdN5iVVBrMntQZDt4NEj139pKbC7HwqiC0qrZQ7
s2AGJ0iduPsxpcMJIE6/osrNp25qsxObnz1GVcxtTCAJZXK4KSpVY8d1LUCkwL9F
zLlxkOvpj6BVKn2uBC1lpb006qEHP4KNtkAk4HV6sVeJi7ntzx9/yvpwEb4XpoC0
QfERxM9JSMVkNMyOz0w4GDsVkenz2r8VJr6pqmTdpc5NNvk5kpb2cyOM7CRnkJ4j
hhDxrZwhZ5fn4MSazsryf9N2S9Jh/z18+uh+L84urbUD1RuGDQYYgU02HyuEI1Pd
bVysWdI26lxPj58Mmf13bO1Wwcg9HH2zYaEhTbo4OGxjdpyHrghFr7BhRDPuDNr0
0EBkSl8+BxmagAFYE9e2HLscmBGNwiZph7LxhOXKEywUHCIWDzBpwG0WiXnOqgAq
z8Wg13s8kIqRFTvXXgIPNjdvWCO8+il3JOjLxBF3UlfO1VKlSDERZPSVTFWwFkmi
YwWd8hYwBBA+w3UOUCu7uD6T4U6Ujb0ywjQptSoSIbzVhfh9R0MfdYfczrMX5oTK
mWRkYviIAlyFYGQeiAsWCWa2iKMX1sAKgS2X2iRuOJchwb4Ve1dJClIRmJf0Nykg
CgAZsFP0KL1cuSiYnqffJnw1bpW0eDiu19WeJFO+N2qLn7pinsZI6xh5i43AjZHb
5rECmh2/3lCpf76OSgBWkW5Rpk+cRbmQA3COyPDusgcSmDMIKYuvNaJpA7zt/fmM
YGQCjGXZG24jLtM8ng8r5+86Qabc9grDnOuBSAfLImoJ1akreXftA55EOaA8IPnd
dr8pF33u6IoYJDQOBwtx5kxRzPxFe8lz9cErtHIIyUOdYFVMBTYFAZAgAlThPeUh
BW47PBn+OxB4QwZwPv15vAkRju6Qp1L3GAif6mbWH38aLXs84rZuKPutfFqq/A+I
7+1hxxfAh8Pw3fHbNE3PAxbkfZma1ymPa6ksw59i6/Pv2076ibwEsWC3y/20TOS6
luaEqHHrKPMOHDfJ53t0QT97Z16sdSIUcnOw1f1QBsRI3cyJYjF1hkM36kQ3yfhe
fi729sKCtya6cqagJ9fNjhQxOYmfUfzSxyChJ8T/sYOihFVy0XuudOeKDwYlLptT
qbmmajNVoQVlUswBenXGGVFk6JwIArL/WMJlpjACWbj5gpbOTjwNZ6mjOPOkZXXn
dpwIDj0SarFp6F6Xpb8fZu7Qd+AKYAEZHAwII50ZF18bsFvTuxUhQwHZY1Y6w1U7
uGBmPk2HfMKZOy9XaY8zF/YGKRg1kLppq/Mer0WZ+MkKUtwuIqEoSxPKNN9Dd7D3
6u/zmc4L32KsydPVRefQsYwtsbjHh0bCrSF/fZgM7oXNajv700ccDri7XdwctQi/
+NpwSasAOXqYnLYjldkws6TKfTHKdtNRHnuaE/LO8nrY8FRHnpkcWo+zXkSuf8jV
+9+uFutKb5Xu5lW00KpSyfhDdCwDfr2b3pbWov6GR0Ov7TNyRm5d5Agje5pLxkct
IRHEFxuEKuoQC+vRCcCLRhs2d7wFwpAb6W99MPtYrVXCX82qIp0hx+ezlpScjZGt
KLRfgxIj6O+mqsxyoqwxWWeWzQThcIntnUorYxAEWCcTU/rRCHUfRGCx48yKfFQ9
WJvaG4h3+ES4OBLxhus3UYP2gwv5hNP/75qobgy6OC9iTCEImxtOoXCtbp3M0xw+
35GlSmvxPjl0rIf/9lPJZxUudnC+dMIU/lSwWIcZpdlbub79zB3K/Bx+deZaBJTy
pfemilMkxYjTZA2BXHlo6INe350InTZLY/ukLSTHSQDj/EV9qkE4eH7yho13JiX5
ntqgLcHV9TT4SYMQIduZDBfhLkHlauc1cj7ZFRWqQZlBCjYXDSYXKfLyrfwsYKg7
iORUlLZc+saUXOvOAD55FiK3TVKoYuJj7a6Cl7qepkC4T2Iq4sn8kCcIksXBwOc4
PI/MktcNmjVMuo/Aa576eSvyMGrJuipq3CGS84hbKTleNr+5dT8nONCeAsB1rPBd
e/R5TwC1dI2pvbcwGWQftlPuQZ7NAG9E54MYyjuXaJKCAJdRktyLFDph83wWUqs6
NbMNyPKVgDPNTXIu0luXm0AzCmU9w23WUzr7SIjPciGW5t+3QKxsL9N4EqTKeMmV
r0aVLDcYyw5nvTPYnjhvlv8qR06MoKLro3R9Lw57g8Zg9M51sq4gt9msUa+mxGQQ
+hCoWXrQvkI5uXVdJUC6CovtRv9OKWy7U3sj0L3NVYd+slqIiR9MDriqZP5beV/N
X2RcPGC5/MAEfcr9dCFcNvUigQ8gZ8jtS5bo2WRdE1cPXdCrh2bIvxHarkMlYPZ0
7eJsHn0cNagIiPsp9r+apvF2u8BXeISIVxVohmbECYsU+q21fWt+iu7pLSPhBeg1
i4O8oTMEazvf+ffUn9AphOBSImipPJdYw/LIk0SEwGKnVn1VOm8pUkzIbMWpEbcK
RdfSnnXlJaSgZBsZm8XU9GUGPnLut4UHgQt51ZOUXWwUrGQesPcxaEJpm7YJMDsJ
F7XDCQuy+UYbCWQ3XESN0hYfQ7jYpGMSQFopTamvvbiPzDPZLsOmUQdna4FXgGAM
7c/a6npRMYJdUQ0PwdOnsrOKBg4kpYTGftI6cG4PnN8+OSXkESnAxvSSTixgtcQZ
QkComKShkinOKnze9wTntvaqs4cYDYzFIX8JdPdwC7CCkpwKh1UFZQqRsgB0IFqu
kcPN7cpzBmXmlYm3zc7Nvjx3M47g63IavXx7kTuqyG04EyL+71rSDI470cnAJ88j
CKhEYNLzWDqsq7juxQH3quMN9gY9RNZQlxQimqWAnVz9zvhx1/JR0xOaGWLvCODa
Bd9LL0RpCmy/dZRe2qGAZEep0hYh3aHyCoh8oQnvEuVi3oapZOnmEnxeth23qdRO
DM24m9ry7AY4FFzneKNxeXvKrLCuuSJm2EXpa/mfHcCtUszdF/Yw64NL7BdjdqWM
YuZKn50YnI5YNprVcZdNgvnqL9QXSSCPPrJfawpN3WvcfCsOkt1FfNZaSGAX2kFe
4RmI10RbG4yrUleN9aypaRGkVBNt1F72IhVUJnYMfe5iiBd3aOLwTHA60tPkIrPw
VXKXVflqsHUcrovRlqSFb3DougZJr9exmkovhxoWSHOG1vSPFic29lZeHp1hFrTp
m3tn68nVsU5iKUeRtK2y6mJ/Yd+imMW1EHwxABoojpZxjFT2aa4vsvqcbd394C2u
NEo6WQMYLb9y+FMJ5HTSJsEo0z7hXzhuvL8DuBXTevVVtcKZ9KASGyO4AQ6XzSEI
PtGJBqUFyim8cYFO6rT99CsPEKcl7ve381nME5sOT0NjZDjWsWLKoxfwMk82kvOn
rzyvKowpwPTcsEaltj4u0XhWwiW1GDoBTxuv/7Q5zrqJeLDwrr8XQX3a6gWE9Iti
U2SNhmY4eWvT+IjZqFrVd11jIAoZuHmmAWyxYKXmCkgA8gYydzmg7kQVZiYFGZOC
rTOLY5X5ENFnDudBwLenUGrAOYDoxmtoY7qGymZLfY3fk14XmD8SAFxqsgRxtDVF
72Nc7vZveG8wFoX2MGZqNcxJ+TXa5kecH6IMFrBU6APNZ7ScidI4NiRJn7TaNAA6
6URNaAhiQjoKco1z1eqsNCKLdtME62SsT86HWN4epyXkW/taKaXJ6JNceylOrmzw
jWHuKqieWyA86ON3X7r9iPA4L1KMDRc0c8qcYvACZP9+6hS790LXfvyZBObzDnrH
mDiB5HiseHvDnVG18HlBeLM1eL2AIyAsLxot9TziUx7ievSDs4IwK1a94G45IKE1
GofCVv1oBjV2nIB3HNd6oRi+jR+h9hzE8hdnyLdpdiqlxoGzpzpD0M/jtzRAWYmX
88aaSh+Z+sG/WnUsdbuQLYd07ILaT6zoCJPjKTFpTCbTKhyNkcpC/zBeFCuz2JRh
kXA4BooCNmXgmqmwOJ2Td648upiP6lox+doVss9WqPi6RHMKea9rlCwk5tKfIbLa
M/42X910GxWWjgmFS6ipmav5DrvXLZNpwG8i7Z9PzaBUuneHCE3ybI7xTioXJ7SJ
+Xgaftw69OJfB+LeiqCF/EmyYfXYBtufuou2JDS/KNEdP2BbcgU3LtobqIWD3eME
c/91pqMoqyqTqBeQF3/xMxRCWgZQYUSOYnBJ0oCYHRXm0pLsTzNZoTWJ6KrRuFjy
QFmiWCC0FGjuvGTLa+6IQ8ZCO4BEAzBhfTefmnVamCUdGFXofLJswc2mTA1eK2ka
fbpq5hwLrIDyvJXeEl7o9jEPqbGFF1qfGuCLCyTzW9SoByaMqEmLSOI18RXfTS1r
hBSLGsyXnasmAxqgAjGal9mkA/eyHlD8HNx7Ps8N3nvdxbuWcnzzqAdtFhGPbMFm
ZFOwrkdsr59v9utInlo8MDNqVRRIWVyw8lHjqrOKe9qCYNzoPWo/qYS08hGfGID5
nkGuRiuxQRn8aKReOGx4oP9XQhrnaRrwnfDhsc3o4heW0kKussE0ToFEbnPM/qVS
oon1vDqTFHWpaeYi6DnyTxRRntdjc2iC8KfuaiFGeP0jIS7yFqseHBTZ/VZ7YPmz
T2s4j0Ypvud6zcDbPeKOBq/x8xkujAX4jJPLEiGALQOz8i/ddhepbxh/mJtSxyQl
u0LbsP/gfC95Ldy4KyIIxhU3Dp2APzkP0xkOrACWRzOLLVXVctH4DOZqB3d5T262
BeoFfYXEBgyYluYPNywUv38lHPP2YOsY7RWFSTcAwQ9De9PIp6nfApyiD5ZBd2ii
bvZdMwlkqliZ+/mUEll63b3I4aORoy/OroDCfUab57KZ8IggwrsP89CTMIarGNGk
UvVZbs2r/TsWKA0PA/zvPFy6rirOWLvy7FFVth7Bmgoat4ghyygmejCZTxmZIL17
yuyr3fvaqkWFsqHKF26ZK7nU0yIY5mzs081IHa92XRUrv1hA2yNG6MQVjiLnP/v6
ueHp0j+N3mKE0ZKLPgplXvwivhyhnNu9R3PFzyExE1qPSMWTvwptpPNwYL36fWee
17ho1JNW04KMVtQcMBk/3gkTTO86xWmYLmzP4sqXCwy0HWMeG5lRLezoBnD4K8GR
cA8noaRxnjwex2fkY8LKWS+qFnQ3BH3TfrZ2+22QqDXt8i8g8a845zMOdiba07DL
PDb2NZ+0ZhB3WgO4F17Bbvys452I7yHTDTF7ZioeuPv2jdoGWQZR7CmZ71+aDu2t
vZaEZTVqaw55zUv95XPdkArA7FV9KP1AhkbLLPmms/1Omj96BcyvmZqzsoAqzlkW
SrFAUvmlrzN4MeczqwkulOTH2eXEfAjUNK7IGxvvs3+/STMivyZjnCsQozT1kRrk
FCIaN3gsFMMqQYHUnMSUA+Zb09wpHuwA8j80E+Wvr7HVzgK7zrhfxPgvZyadpb7+
/lyd6Qe/gsqlBNmtj3hyb5sWRCAyUAUa7f3C1tCLI/ntgZNf6Li8sEYVE8bTgjvF
JZNKkZeS++ED//MsivkW3GzBvGu8SQrAhDjpI0QzNBcgT3Mx541fYbcWTN5VO9fy
UQ019adFl5J8t+zaUUcrIrYj7WhmoMt9RkPILB/j69WbCNo42WG/OHJhuyT8yEKq
IVdvqt3vU7wrT5X7gZ7eYqbOpQrfmuu0wWAfRdUhLfUw+pj3jkM6jUUU4fSWEMTT
oGcGLgnpdzdCtsps41c2g2+VCTMJ9uqCHUDFgTUhrjGKz2ifuuQnC7vy4mC9sywo
qFrraEuoL1NZLs950KwQqXU8Eh5TGM7d1rmx+bPon3i//XUigMxZPlXzAuSb826r
85ZFqfNwBHkXi7jhq3YLmQwudX02Z3fa6695D3yYBV+ptJ6EhvGZ8PnEVSOiwLGh
QHupnkvS0vTmi6YZnrr0T4cPXQTrQQVIlzgOHdjQ+XKd4LoPCn9SjhaEJ8ax0eSJ
Xvay5FP45lB7CbN2DuTLdsEyVt4jbt+Ins0xmYElWsSLQ0o8VYTvsspjwLIOGku+
YUgT3d2KaXmgGQrd6LUzbZrf+JMhOeXkTrbiBTFhgfV76+rtNNvoFL5DhFR8cySO
tOEDcE7/MVEmBKeptx3IJOz5c6CM7At2FjXvuMYkbwS3VYPONKqYh5z8bEz+51u6
IcDlrljbucyUfRab+EpbDyP5/Kz/TwEMTxvs8XRmmuHiTfY3vLzRfuyuLGuDhy2j
mASyDc3aWKciha4Mag0Lc3wsD6ruRJYuhOVvlVJYIhLacWBX/hrICV8a9ECbCm2y
bOKgnFv5yfNAnG/N846NNHYPWaBJIjLMDq5iLSl2jTpe60ouoIbuZ36HuZm9Y/t/
8Rn5fOBNVt/hQPec8EJdXSK6hzhlrGwI4Lylm8KcXEpipagPM0ypAkr90PFzuoRm
NH0klpbOV7ZO9Eef+Hzo7tVwybt5lnm2xTqAIBxN/zYRvS4qdJramXgC4KwI0Fot
8A92/IELOj3v2UsojCsPyLnu2X0zUoUQ7bRK0xODPcp1GBiclQGw6JLoYGk77dGQ
f/vNE2S/YYoV7Il1S5VbeevuyjEWEsbVHx9I8M551Givf9f88nXGdczsNfHZM2Jg
/Pd8jVRILkmSaa0jQdNIq3G2eQomEZM+5BHvCGKKYu67rjay/AmrBgnM4spaCq5x
Q3Bv8dATO6tWS8LWUHgrj+hfiSpoj1MNcE0TqepAXLppljakWpxGbQ0G6Y0PIAqg
wbV4JclmW5B7l6jTPvdOwAijA0aathIkK+JDuZq7OvEluoPgMco8HZuLbxZt5qqQ
909mktjaHrCabLTp5DNXtrLWGkM4RhhzDIoXN7SdYwHr7h+Qn2pcpcV0R+7qZo/4
uaiV+loro1UN+LstC01fwF6NwbrFAYNFLZhF4tXbY76uJ/hNDLBQzFnSA0VvPzU9
NNX1aziAJCBXsLQCCzHuADOZZfy1YcpIZsxzJdGsmMIjYunjXiWvL9j2XOUoGo+P
eujHiM9D+G+0qAKd0yZrxC9PeqM10t8Jm+Q/bNMoJN6Vs55pO34l1j3yYK0UHtHX
CQECFThCsgkE3+dpTWUY97OGmWhkztklVlTj580y1J6SD8aKEZo/Gn2S30QAczZl
luSDcuqQYFuVr23XOTPQDemtvqUaNGemWtq0W5WOQHWxCcGfXBl321xJIozs+WG+
ODjzuqjWNbyghOvfxQ4/ZP6xrj/MyKrpEdD2z9uatq3VgLf2PyVEoa1BLVvGW23n
DeL91dVm3RG2n8DdwRwp2WBoi14F6iMT7wlZJXy6HkKm+VgW3cgbWjl9ee53XVFw
1UNDx5fU9G9M6Z7XX5uvY3Lwino2HsX0WQKQLC1KgUtkLPyuJlBrOM1Cri+aKbWu
bEjZZAxPDVYD6cTMZ8qtogmWHB93Bq/ik387cV8TryYxC6Ky4Zq0LstKi8TshcSa
j38l7pEEiQCI5HgOEA7mp46g9eS9X35d8oMozmi6kiw/v6B3u74BbeDjy0SETgRp
0gqx0EtR7xHWs20xeHnLa2WBft03b8b152LenRSXk1bzcDgxl50mNfSku9itSPH8
cu4Cu1Zmv1OZ+tl4yMjGrcAJwPnB4vDdCtR/GL3G0eXYPbhM80fsV2LLeaWK/mrw
ENJaObZi+15tfQVTXIB85lNJfGqGGYRsIftqa/xQ/LEAppM43BUbaLLrHZgovVbl
9bBT4xrRvMfRUdj0hGyYfEg8ZHJ1nCnEECi9LcDQ3lAfwEpuWPWY73dTVeoYQT42
VPnzuLPZziP/shg5p4l11dy2U2HinmHMq+rzl6WZKc6DxxL5eXOg1JFqJ8Lkcp71
kOLO3tfGKZ4r0ratOkwlqxiUurvQkqPiDs1TIM2AJ0ALz1FEMyxjy6t84yyj2jU3
cPKIH4k2pmDlcY06Exgxr8LcPtfu2zY1QjlW16PPrYVlnZoRiLao0DarKJBLH8Ud
NLAQbaH9RH952vrTYO0HBqP4SGmjTLiIreNK7JyMRlwIU2WtuSkL4D7lbXAh+b53
3fbLSdaZWV/OZFdqiDnj5vT73pD7iYYykKOEFK1aDh8ib9M7uWaC4F8BqWLOnPkj
fi/Q/sT5IpqumuLSuEaDDlJ9PrUVww2Ls2H2LsZkiwDbwtl9gy65pp+2nKW+ZVvX
AAo33LfMwjBmFLW9owmIxmGBFXfx4GEJmCznmVsYoeYdUyHRZqK8J+EeBaq35IqW
6drUA6EZZxKbZlaFQm+SQWWSmchPtK22dkRbGUf5RHGnE/OCQ4akfONCsx/cpYo5
CiBzQcOAuJB/89naRj7hM8vq0chsyq/Py0mIY5RLAJm8Nz9eCj0gwFWt0tZ9bZkr
m93AgmwmKXz1TvBLM4zhHMwa+BYdQT/x4740ZrFEfpwxEmT8sKqWRG94P9PTQjhE
/jWZ4LuAjopCqKU9drrmnYJkrL4nrM1gMOE2qpogQ08AnfV0M/xVzj5D9CrhoBIj
Uycb8Kf4LMDXATutcnj1U1a7hZatzw9YN3MYB0y2+S1KBj2dfFYly6qZrmxuTmav
Y+wGuo7YxZsF1+3g7BLHTBjfRN/XVhUKnsDPQ+vj90fmXi/tGATlu7cDPltHjBjM
aRVB0RMRpnW3B3oXx58JG5Y97Xb7455Gw9xTuJKkzMI3+gnROkg8pnVzZjAplqVC
fs5e9UgGHOx3FIf5zQzEu6alos8AdVaEqY6gT9T8W6lXnKSGDUfXyV0E74WazPfT
UqPG1LXT0dByMOKuj4MWJj4zMbFsM/FIPKabKYGCKkAk+TYcbXDnudo5AYiCVlXo
pAKjIfMr4y114VHs5CXPZVTREwjahcEZctp/rj4Nnkq1P1GT9SX7dfivXacygIfl
Vg+GulCmi/jfIa0LMzbK+TqmRsomsxKXOL0Rq9Oh0V8hHAByJn+i8CuDr8H6aRUb
4NTvFm+jiyUvj/cHLRytP3zaf7Z8/H1sw05NYpjan9LPFSk9G95prj9yYyozsHuB
xCkQ0VmJDWoV6nclMnH0AoHutYgaDaWFR/dtmdUTEUYuzH3UCNVOT2IKhwsI55vN
3dBhJ3jZLnSwHWu/OKaimQ2OBX1LguCWQQ2JhG8EOP0kbwCT2e8m1YnQ4sy5Fg9H
dZXsHMi2mDxxfJYSZ08JWC59v0ACLUmOV8KnEBHBTZRRYO7b/khqwXs/LHe3a7nH
XfFA8eDroYpbiZRTvVPfjoC7vWYbm1m733YoIW5llLhN6EKE+KVasOPod61KDnWB
G6VMl21+im3EIihJYAZDVkbYvBYo4w1eUa4YcIp2zqV40BbxN0ElWYFgb8m3S18K
/V5KJqUaZ13IoZEPMim3JZQ3POK3h9CZcYSRxoWNfFF6T714SH6WL1Z33N+O4nXx
R66lYyw5T7uABfuMLluqtDFFJYQEyoce+Xc5JusV8u4JjFN/0t0hxWYkgJ4zSjZN
1lKTrBPKVHpb1T09Oh9tsjqvPWX7ae/S6uBJ21wnfcD8vwcalrBCGX0Mb1oveKLM
ckbqZmRnf545CRXb5tk7IK0HNN6EiNhlQv0pLwTMdXQfRbGrTcxlly9pAzvxaAN5
2uR6Iw4SLUgCN4SpZjAmK8k3jDBIRHX+gyo4ZlPhqMhMBw5We88B4gofy8SAtmcB
LhlCYGREHVOQz3Ye4oPlEOVGQ79RQydy+83sb7xKOaNwNiYDbzfdXuFt0/FeQ0VX
/IZiM9mFhINZJkVzhct9dq6DSb2mba02/jUThfCMYGplj8SFOUPKClAaK+F1xLVa
raE5HfrZjvvQM5Fokril6TTEuNqn32yTF52dFZEEq1bJutSq6gSCZDtv2+Gk9ZBn
U1kfCm+6OsxaahaC4AQ9NiDyBf2oAlCKTnnVIZif18+AfD9cmecMQ9syJIST0C4x
n4p7dAfHw5cENJKdDiACb2XSqIpT53yIfAvbIBGJewKbdoqpyqmutfkhy49YtJC7
/wV20v/DHM4d8EQxlUs8NGWzgCf+xrOHl/RGQedJ+NCwVlIc/RuyLrJqTRnFtqUh
B935H4zFoLd4+qvmKZA7H7jlax4sUBLXxbw8tb7Gi+wNIvzxEH6Hmr+wCmOYG8K8
vcLY4L3/trlEoPXXx70q7ECNVW5eivp+/DtSX5bqHVZ2fbk/NIE3JMAVLMqlvJZf
ICIa2HFjZ7GQTQ3zD/PVtXgK/Sgx7kqke8oKeJcS5VHRwKb3exAxoxVNpZNCf3G5
PD4UtiCuvCcpBXlsHGRAIsIS4yIEYLghpzj4pbUusvmx2kGjBvd/w9OED4TeGjpt
IDHekNfGXX2l0JbZYGY7TboR2y2VDnknJ0UbJ0LlfCy27TmTL/Cmn81B+mBAfR/A
IIBzueYdTd+wb76d24JcTzKz9n/Wi/Q1ofxjul1gzwD2C++MgRvtsXQS1/DMktfC
B+fnAF5SB7YYY2Wpy9MP6iIX4Mxm2qdr/eDStJLqA1WO/ljw4NvWWCtQMK3FuJpv
QPSmngnymd9VqluzWrParT99kMvChgvtTYsB0cOd/sfxVhcr0+p31tcfy8M/kZsk
ofNPZwPCTwhO5cVnYh8X2H9eacI4T11dTe6lAjbDUK5ewoorKrzKY0apdw3JAiHt
/drBXocP0UK0+aRDAoHQSeT1HjIMz07Bk8RLE0id3zxD7v8wUslmdx4m72A1T6/n
em/IAlLb9HGQjznyNPkvBC7SiJm6Tcz7/abt4FiY4HVUyV4lGMvcCiQ6XQtucpfX
k7lWVkofG6jSghwOHuKhX6fxKPurdjZYmpZO+pdqvRFt37o6vqOuazjsKO0JGYk6
kvnp1Gvbpw5D+v7wAiKq8plZE4eCf2c2Ps7SXgBStGa7oP/fWpIBiKUWbz+FF7JH
Q1LdLyGVJLsYovbph4AeKHWi2qopN2eUv8ZgaMxsEjveQkY2BuI3UJOZw0je5GRk
JbQgaKq8HjbN+tGOIvvqqF4w9NnJlo+LERh7aIg3oV2FpvJeHN5jluCtrTiWKYHa
BwPyiX3PogpMpzX2nuHzv0n01NtqJpX8V6N14BAGZkofRKbENrDc0qwSCoA578bj
uJyde738bwvh7Wqn3R2A0aRyn14Url9dulWfG/yYjBKwM06rjXrSb+l+O0Cd2580
rK/sVIiliG43eYCICGaGdY/O9KxwRiTGwOt1YNP4nQPOCb4mU9fL1qY2BLBTELha
pvwR/A9kueEOU+egEElBOToYFna2GTcSs3/TxzzWnHzVXHI4tIPsvFSw+bRRpfvl
6Yq+9b0jTNusVqvqjgxZIM4AOZAooz8qzou1FaWXSXpwpYVUoppbuEWh7UuMUpCM
k7YSXiEG86ERUsCtqMtKFlWxBD80AMXmpVlSUYRTgn3hb0sWxSjpEQUaCbf30VG0
FwP8jhyzAuZ24FjIPgFLT5bcslCGSH/XZQZ7uRbmyXVuAltk1P8w3SWdeySTfBGg
9kQ3xvY5tgVtXX7Zb6+n7VWY2+kLwV9US8n7yZAT6v1+daD4+cu6IWVFmGHKKQtU
90w7dftxJ7ZDUgzRLldhYunyGjAOXDM7Qmrjs49cNL72og0A/IhLdn2yt8gvleME
bAUhMOD6rK1TQQ+jN3tCj5Nq0U69ZtVx+W+uLxQg5RkgbI2eSKxi3x2FhIH+S2QX
L3SL9mZdei6D0+c6xdr8rXjbiRHOgOtC6xUR0JdZAaUqdJnZnv0ticS1VoQ4CPs9
QmxWe2VyY3cZxbe0Natsl4q6rEh4l2uKZiOu20AUGfRhqQGCzEToi+XQbDvts+2L
HPmpwyzcFv6przr4w0Y4h/YBvDF7YybO93W5JJsyJdW8/br5gRLU+XcsXU4EeJpt
42Dm02Zm49ZdmjneDO73KlNFXNYL2maPnIGfqo0RX4XGZx/C9AAqFgWGrlBjl98C
X/9RQ8cEWwS1tUAHTxI5vHSRnJXhJXez8BQjlGtDMWc3HF7jS9+JlggDopVOPRMh
hKbLa5lFNUQzhwRKG2flwiSCjIVMB/FepHbnx4PMUoL9KY5ovPhPggaBumVpfEc1
QEbDzL22HD+kTHweK5wCnkIkadAVWqmmpkTKqo4KmKrEwtdZq5bFiXPs3J9pbQWF
6NnKQWDTGKA1gmyf0r3l64OSbpCwQB8QmOrK+sqDgF41BQ7OUpAhsUDCfqDx8h1m
AIINrbZ7zZ9ligKAiMH3FCHpsMLNykOQVxfNRLwf1mK1e+E0OUqs9G3X+zEnMUJJ
HLDA26L3iuNbIcWLCShpnUFTUqv8Eemq9N+xZGIZmL2ow4MwrBcP7PmlysLl7GE7
hKXO9794rQ9DVCLyTo5kscB/lhAPssC47S8n2WghPPO5xHJHvsddBCJ1qxZJWO9R
bK5UmuFsLel3exA9bQOLmg/m3GDV7Fy/LcT7ZBQZHgRChm2usYJ9E+28jPXadsHH
jch1rIsOrK2+z/67ZZX28tjSJNPNaAxVUOveA/efbTwcK0jZxuKU45EcM72lK4Tt
TCcweXyiOTZONKzuUFxRKa9Oqjl3I6NWQPI1wYC3YsAuwEwauJ9tUunkJJyf7ie2
mHDD4QMPpeVQs53QTUXr3A==
`pragma protect end_protected
