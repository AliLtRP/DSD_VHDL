// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gQ/Pqnq4Oq9zp7KqGG37Y2ypBzwqi4gPhMKHjuRRKwV87l5FoqYcQQis2HINSJn7
MGRgp6+yvVhRKGXoJxn3uoK/RIbkKpq8l9nDSuF0b/3905JLrdr79RSWLfspN9DT
6eQATcdxHCBHMPG9bkQeHITAISZ6E3AWaWE/6hmWS4o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18272)
g6K0ERu9ofW4qGHGJ5el/f360HsGbulIAjVTwCb8HBozKwKtKLfY4THzpeH4pqry
VgHCqngSmm+kDmfpK8AEKmVxAqBm+N3L6mZs/JhPM3IL/MNwSU3QvllMCs7zpjdG
uD7ATe4vuw7SFz2XryXrYu/XgEnErHx48jvVzN5yUYXY9foh/yexUPLJSnmGgDeW
HhbGLMR/3NGz8VUjoIbCLiHdB1jPUQElUTU4DyZ4omEgKr5pZbexLoX1SLHDBbxx
hG64kMwNb3dgyMMY9AYMn2TTC5tb6d1U8ygl0vbQJqrNsG1vVNJsQr1gz5byN+kQ
6HBfYuM/sITHXqpM7kg9Nte4yX9RVMC9zv3FRldL8Wgo7oNnJB5azICgfV60KX/U
xN+tucmWlMuDXl77djFQiNuoUq7YFuobRtktgFPUlG6vfBbhwPvVNvERg770WYm2
L+RlZpSU6W29FKN5bjdQnXHcdArJ7IR/NBJj9iu+nej5CO5zWBr7PY3BaBTECzOb
IkXG//Na8+bVZW54Pf8o6WqXLvRZBsU3gx3WuQ8gIhxbafzWKZvLX6SymCJK1njm
Ro19NYguDLaGW7pXJk8gM/N77sUbyxhvDm94zUhnBqJSCM2eqsilf8nepSdrAoQY
o1NoIX/e+9IQzNSFVrlvkOQoQnOKSxA/BHWQTiWBrxHeuM7xqKA9eLCjfXcwkpXl
dnrdhvlHLzsZmooSjzi9WDzoUKlA7RqbEHoqCGBKIgf2vY+qO/j2YIaPh6aO/gUn
jrbawkmhbCofpaJTSTCfnOTUiiEjl/Ftbt5eIr0ysu0UR4wkD86OUO5l0hYcSBWk
VYpz5bcmzJkAOSl2sUkt3LelnD9wWEMQ0QaGWP7Ju8o+l6VnzJAB5fAXxqQZAX1m
cYd3dosTSQiu70kiTO9HfFwPJQiKZAjZpTSng/ai2GtdSVPlQF8njDrVhrXhqUPD
lYgmeL70As/ps3gUS4+izdFCztCXMPbvhaVkpwC8iFH3cAxvr10UTTmupYZFJOFN
RLM39EdiWPS140/h9DGeI+1dBeGTEkt3t8YNvBBEc+FNaN/tSPj0s5+vyGC61WtM
W5ouof1iKqC4bDZ4tuCILODsL9Z1iTG6ZgnbXtAK0+F6rQOqEpvV50iQTqvxc98I
J5ITYCFV2O2S+OliNwIhxQdw5LY0IbGU3NZxVDl6fANS4028MtBXsSSKRS9wnAE3
e/VB7/QG42hECnJi0vf1fHC+2vEGipGP4IDL3nh0n6GGZURfvm86VpBoEiclA5yT
lZdYsp7Fpc3MYDA2tSiM0mHl9HWt2KM06VyW6lpfqM3wsrl1z5qQQ24JB2qLXxS4
czf2M4oVAEU+4l49opN/oi8NwPqk0k0IdA/sO7QJBLWQmSMfgaDpngo50b6NwUb+
xrTyI+CLo7TbVpT6dKiBvz3W60HUSNSTS/NmroHhHvi7zdXgCUbJjq50zAUptC+P
anAO4bCJIIUBnk3e0jyi4P0Z5B+L3ptdG8oc0YFWVoIYe/vtDmSDePBda3GfNGup
dEnoWM3sd4bGhdtB/uvl82nwPApAdKrgSYRR1/qSk0wEsepVrE0Rtmtz2sGYsFzF
7L6LNOjOYzpSVrlddglBvA+jYWPoAUJ8fqw1UphX2AWnSvmKXAK+Q7gVA6/rVRXz
J6srKCQDvJlocyZFYIWBcEP81kDrI6YjkNIC100Vd6PqFT0XLzejC9ijfuit7iO3
i7VF2RAMcE+sQfX0aimmfKfD3DFCFZtCCmlJMu875dgvHAplsHueEPbXGCU9fyoC
BVdCybzfrXlf+3dTqLBNXWhrKEWuY4neb34l62ln5bbYCpaD2uaIIxFWg3utt6IS
+tNBTI2b5oKH37IbWutedPTmDWsKZ+euvdtT8YN8m2WttCZo0hLtzcNjGxd6tuAq
th9IJTZpaHG0bM95UYSTgX6ZGh3SX5QNd9oYPPx8lplCDQjA71lb6CqGRE2GT4xP
Z0p4OlpaivDjpNkd7M7AZfJMy4oNEJDaLP3KK+bJNiEhemt4LR1llulTDimUlaPm
6pJVL+lkIQOjrnjxFTId+t33Wru/ulJz0t9PF9DrobYMw01nHFDw70WqRdKcyxkH
44ZfF7xL501ZtFicxcpttKRIERpODRLZJ6rskXs3SNtJ0Wofmgg2kBoTR1bluNUA
qrM/En5gu8FbPtYM17bE9O/rvzw3nb50tiNCLqB03m47oma0+FwIZK3urxzN5z1X
yVePOF/2aZ94tRAcXz8NKctaI4xECWNWMI0lBLlmugFNfTeEP94iw3I4sh1wnAcf
T8VjcxjygpgYA+m3lQ9j/GyLe/ZqHruBqPtph7FobH/ajg0PrlsSLVGhV06IBOxz
/4DFEK2OKpn4wtEC1qt5ygIubOsB4yTmaKBubRj7c/znfNd8KkGeUTAsWoR3bjO7
gHguTMNCtKcP6cAsT4ooOJUn9XVTHUXDcA61O8xEpvjQn3QAPHKrKDS5KQvphZrL
Cztvr83ba0DfRIxe96x6KZAog7PhPwO+jZuGpYzeBY7F8QALo6Z29STsA57LNfu5
vZ0o+eEQnio9+kXuMVvG/yTUv9NZVTIqnAKRumY2Kngf+dPpcEr8JIF1JAmZ6d9P
JfEVGvT7/8wB20OJ6W9u9CH/ML1/UHpWeXlDXvLWTvc/RX4Og2EoObhgql2ahjKG
GTwvj6hDxHlAJvfnHTXLsNAAisvNZLKvcpmPr0Z3ELvKC7+adAlN3HJpnVVzlZAF
wNhAU2dwRCUuDXIhhbh5CJzywj4jQTmlR4wy1yCKeRuP9ov7dHYm4s03MgNYxk+u
U79ug/k3U5yL2Rv2aF/WqgPlSbNKSAuW+00+y3RAlmJr656GXJ20qE/EXiEVbacM
/nScAC1dLHtzhfNgiFXqVhlM6bHxG/O0Xzz4SE4vQCJGarZf639X7rxU9TCc/h6v
o4jkLfs6T/tkGWZega22zD83lSxWbwsur5pFQZZdx3R4PHRMsbjY4OFnPVLztKAD
3UGfYr66k45KQ0lx+aFKSFQCOKc+CvPWtWWMI3vD5s9v83NEGDDMm0dUnWZ43AHC
kjmzUU5oHJtwgHFdrRt910qVFjOUUEr/1aQfncrecyvWLxlN8iJm5++PZKlff3N/
oJYmm7S3jENTvBG96pw3Sg7/QQPFLED75CzpCk+s7Js9Pxk2LxqH/LWcvXMp5P/N
0jLTwdHlRlM4z03BEbhMFmv6xz3S+nNkY5MbAx540nuN+OF0VWKFLezQXd+nsxke
DZSzxR9Duxa/by8KTf62tWoYkZ73gsNNH4e3b3jG9TNBl+WqCUCO79aAKFNIcwGR
BOJNIg2Hex7ZsjPipSJVLa6B2G5lvF0StzBRxzR+Okqc9cUeVlstLkZMGlYuXcv0
NnPMIwAcoMQNV+KNUiQFiSUTVfoOIeg1rqmCdIAfyAeKByKC9gW3dnYjn1DZJeRR
33YZuH0MILNuoethRsO5dKWuNdE1Z4tWwg3vXs9n/wlYzGEv+2g4DpCYU58lixpu
uAHrt9YLyeWMVBUXEd7tFgOUNNQPgltsu5/lN7EQPENGZ1O5FmzUuEMTfdcIK3lV
9Kpk1EhoyHwu7sn0vvOueiwQgDb/+joXZLRm6VuYuey+4KUyRmYEMPCh+3AB+8xj
//PtMEaqyeuEoXJUjJw14DLV+0HMrmnzGn5WMPbtvnAHQ0dtoayBdpA5VzKXrEuu
zlCPVD1dmmDG7b/9AqSVMNHC79pLFJuOMGoGSeMWHfTFQEX2bxvHY2IvsNaojYqQ
uVpgGB/IZBXRk71J8gUSrLZJ3KQpUxbzljGDMur3qlqpbLU9L/iFX1StqMRz4cti
HKy23tLAR9nnFsC0BKEdJ8GzZcJ40IgIfeGfqgo33+NONM4mh65Mj+5r98EBgpK9
60jEUXtnZ/FQ7mY0Xv21/NbNPWcIR3K8SCsNUnxtDEaKFppzPqT+1hlDwMl/UR6F
ZBnkUExcFZB9hhtFBUWvpZjcWDO4/EF3Oe5O1glGkrKY7NMFkMrLTUhrUbKake7O
eAQFge0PP39K6KWUpm8DViAy2Cuutx3x3VAledE3DMk1ebYHFgScin15d4Z33B7l
648JdVGpP2ZepVDQDlmxJwkhrGHD2del0m3CvYT7mFhMifedMaaBtz00dKnFya9h
XZ4c3AM1eE7+k7TUWpDyWCRaVYkJpD4dJHOQnfxvSuU7sLZk8/whk1SukWbFOwML
cyCqCmZJSUBS8KNhl5yI3oAbE45a0M5k+nt1BgjoYp2ChKxpbVUa1VfitW/F9Ftc
/wfQr1hpbW4V+n99SU1Q0/6mmYfqnF/47KxEzNqBXRpbvhZjhBo1oEdfYw1dJJFn
RJYuF+fmTum2qGX9SIVWlT8exhvxHqa6iBoXcaCVeBNJHYx2qVrW13J2ipULACXU
gr3+xx/tdtwW7fJ+22sn6Doyl3SfLbz7xzT+ag21LgAYJEyN2bEwqOshspYCLqUi
qU++FcZkfOkY+9jT9wnBNtR1XQqqByr2a19dIHTPa5wVKwg0LuqIMmyBTNSnpjlo
vHnjcZncDp+eotDZxKIlNd5dS/q4W5rOGGAxi1XGoHwnLI+l1C+203e8d+ymY+kd
v40b9gNDTYo2zVfxDIn0+U7+SnQo3/2HM1Kgb15syon0ZiiG5WDFnQP2kYnasttU
mJCQ6KQcRzyVzHTnkPzWZoxI3GIhciJQ1qX+e5217ivGy7yz8wC+BkcrUwp1dfjW
AasYoMZAHBZybCjTRFMaNa7MT4/aQt/Zb61CK3DvnWjtYCzbogyNoMKzQXVhxguJ
fzu7TH8IQW1/djKSDSqHuDv4IagDt84xyLv42qxVzfqcKKqDTVmup73E829MXLzc
ziDiQ7ZljcLXqJRObLN/B9SRddKdBqrqN+4Se0yiYhfrq7MnQilqXa9be6kSEn1a
/ygWPwLN3Xvhyb6k5DLLKE5PbwWRLgBsK7j54rZZLSM3Uz1fl2vMgg8Rh89yEX/B
yWC56k67kbvkptZpJtyA3gmmVBBFxB5oSLDI4EHLMM7ZzPtvITL6yySjzLpHKwqb
ycPXY3qt9C4IRB/0ESOtE8qxspqCor9EA60O18xvafVDLyP/zp5cJFj3Pppin4Ax
FiDNCZoMJBfIvfFdTmO7mHmg0NcoyLDVS5klDCr/3flzD4v3gQoZz5N04u0SUpQL
1W/1PMZwKJ37dULG5pXdnktnK0Fjrvr2GaYgJooGgvgSVrtMmuHiprDY7RhDyuSf
YpRct7nsCgL5/jVhdt2OeIJSfm8Pprov8C1HyExFZtsP6A49+rq346jPOlAYxysK
Aafzf9TAV1VnKqKmscxRxlfbS+zxdAJ1j4qqlXFuL6vyto12Si59wf+HaABpLsMr
3QF1atmeuONMi4/69v/l6RsIXaKPvly1NKaiInNvV4FtzGhVFtV6JIlEJ6+qK5cL
TRz5BSNTutp74cbb9HU3AqT5dMRXwrLoDGEHAYE06NIzlmf7EdwaBMz3ZD3u0ay7
V9709QH28XA0L4GqNE4l23SQMp+5pn8NsFkw/uUhtNrfBY+0+cR2uLHKQXXgnpR/
t1GGt3MYR6EdIXqggXVNmHB97wzsMoHpoqOK79VMgNcaTSmwscOQS0CMJWzW3Ls1
IV67/SYKC8gzYppjF7vUk3sj7/2tbptfC/TyA+ecQuAgH4/xIm5hwZvFQ0eNXu4a
j6JB6GBxpfj8UOi0BAJv/ZRG2yesD8h18W/obaOD8Fy232uDmr9gAEemcKJ/W+SH
7poCmsWIoduOn9Qc3o8Y0LNDDgGQyOqkMK71wwZm92dpVwhPs3BpYijxAtAbwEqq
ZZe7O6/VaOwKFIKz8jR/qsqNfNeRdEL+IvowH2oDs9AMNDmCYjg56j8WabU3hoWU
eVpcavVC670GTPjT0O5C2adhjtKSWARIQox1omFyyOXSj9k6oDKYrUNCwex8edha
OVcOuIYd2u4CRMV/fh2DpuH/CYTw//UTrdIv8h/lER6V6jdR1pB9QHN9uPdJg+V0
yZS0evgnawbP6x8wbvVn3e4lLrli5agi9WdDSczrJ6cHxyWgsFSo/+kpdxDnaXgW
SFigTAWiloltbDELX73oYYmGfs1dyq/stJysXKruZm6b68YUn4nQQ4QL8p7EINs7
JrtIPqFeWVYHHywackS4k16+e0NXzb4k6ApI3QsDZ5svilb/MeE4Fcm3swsO8+tA
dQHMgnU1ZGzO3qxeMnqUAHJCyZ8PigSwsHbuVHJC0UDODCrohA4UtWCKjXBWWarp
AKf/fjnOacbLDmVmU2ZuAcoeyz23C+0O7TT5vVbxMnhXgx1ZFX+sxBiMVlIQVVQf
ox2JExH4p6kOINzQUQPJyyyj5zPCvtgkIU1m+lygsK1wpez00n3VMw1UBQ3LP6Zf
wMApz3gVUcJZmUy2mg9qckwXO/eOlNUPYVbUUeiq4NEUrAOUD2g1rFC+MS8tcoWw
tX9AWNkTOqw8MLEDKXhhfJxdCirlgc4qkTlNnMD0KujjGrzry30Kpn0hRTZCcSyF
BbdjtL2PCRckntQBva9e3iEiH5xbW/ozUyQMUTr3wimV//Ih3cRXXkpBcpfNbgLz
9kGt13nlE4vI2Q52BXBcd0c+nBQ+TiT0Ay51Qy5JFKpwjY5BZWoD3ReTEEgaac/6
SGSlYagS/rcm3YzHvp5PoENodO91zGxh76XSTgnPLwvV9H5gSUggIqr+0R+EAoBI
rCAjcJi7BDv75KaGM4BIh8k4iETGqobTzVXHcngX2ptTf78PKaRsOhgdq02qLAXP
vOFBRiqMc1qmouwojo0khL2Vm8TTiJbX6Mba3BW11q92vaKaQ1SphDjyDX5a+Oqd
4azAYnepHPXRwYYFgiYrO+eJibF5m+pFzPR5Upu86+ryNnj055hFXvDmLrYWvRjB
Octi1QzgJvWwrbSvYwMzD59b1CFRp+X9egpuf4dELCg/9uEanvO4Q0MH7lVMto9k
Wk152vkZ+YPFTLYiZJDRrrQfwWlx+SkTJOBpDzNMcYeE+8dQ2DrF1I4txVvUxAMO
gbbp5QQ1nGuoB7aVg1Q5GnO2VoBxWclAoMBTR8yUhtChz33FYzBb/9vpzzltrax4
QXzugPqd+MFe00pD6kdaKKuxTT1F54BW+ZKSOx+VhAPpG/ieXky9x4f6VOX0Fvdb
yr0VS9DRoNkQqKjuFSMTJrHaYcv6M6TaXwrN7c6FUx1/l48RBr/Gh/0XbDPU530q
SmpGlH55lo5isr7gqIAl6KvTOQgc6PgCOI/Wx/izOhKY99moSUfiSpcxIRu9r1OI
qiYhrO8BIgNcSWQMXJMgnXYBOK787PrJa71gmmr8GcU9aEWoD8RHZsemEY4v58Df
ty64u3KYC7yXCZGAuUhoOLkIbWUGnAV+stsKW1HOLwOBxer/JtaNvEVGyGYaJEAj
C3j+m8Sx7Lx0zzyOyULEcVbeyZE1KEU1LIqqi6ADrhHqpDBMyf0VY01uG7s8C5Ms
b94Xzbiad7sv5lgVCKB4pp+JHrcaJBi0XhqV5/me0BihoD1lAZnMvpK1jUpMcu9L
28oUDnQZv73o2P5JZlepFj3Gt1PlkniLk1cQvvZnHfZpw6s4UF/RFSv9p9yB/PgG
9jdjmLHM2pNVcUECMCG1WVgbDcTnf0rzaRbOiIHdHNLv7IaZ7F+zqix7tEMhKhL4
+db/Vjonc1H+jVpfSJZnuJytgN/sGb8H2zHgW4fbarvKlRwWZRz1BtkhCxXbaRNj
lSP/70T+9HepSiXF81QpMtQ9kAQl0oUbbxIU/h6paXnN0u++uQwTuWgNLxkHYW+L
h6jZaW+9RScjLFm7Xp9QOv41MeGXbsR4z10qUlN3+VsLRVYM0PSY7hUjojh2KyUK
a/y84nHBvC78WzWg6Eciq1zv6Eh/Vw6QrH0cYvfSsXT4UofCiRh03zwBsmQqA2Xp
g4GFp0E1bxjPlOvpibRutdcTDSLmyKy/dbWPAdH/uCtdBG5N104lo0nmMl4ohvjA
WzdVvNYcntNT5u92//KkiFATQG20rdlG7s5PUUuWeKystX4lRu+ujeKkErOlfzHa
uB8NLgRVhMbdWq+CCyM25Oc0LoG/cSD58dQOSBpgYmwcu4cx9sXwp0MSK35LXQQE
ufXCs7/inX8Yd/pXVBvIY7nTBmX77e+nTOr4EfM5W0BsW16Dx1576LuzHOR+dZec
f34HbBTSt4aK4uvxSDtehzrefOFavulSrjIrYa0gg9MCN8fUgB/DIUrSbP/7anJq
zp17erplnwFpHfjb2kVCswYu4KsIKcwZTKsr4esUVVX7u+9+qvMTDpz1E4G7/QvT
0uk/klARgWveUqc/BCkJ9J70CIZVb9OKZwcVySnP7qu6qnEUP/JAlSQUXB0Kn9NK
5YutfKQ96ovNSDTaBE4rduwDMYBbw/fQxhb/2qbLIuOrsZVUVAt38t7TyF056juR
Ksi1gX9uvGdTHdiggI3yp6ecVm25oReiXuI2EpZa57EzQTOb0IhQdUfFChz+G5kj
L9Bphhrim/DEssmEZFJg8+vGn2AASiIh+jVtjAdN8PLjszDt5YMIqCVJbLP+yHtJ
1xsLKmD9MJw0Fgw6zATFxK7FbR+JeMu28gkk6KUy3i5Lpgr4g5s/niMALPgpMaY3
K0isLPEMf1FIwxo3sYzMJB8ZlZ/fBYqBqMd5P7MngPnOxepluRS5QmhtPOx4caki
9pmiqcvXueIS596NILKxu4xz+NvY4WAxqFpr29nC8rnEgDuSIz/Yf2aYKN7Ld6NL
oxemvBmWlE6WNRSlIw7LPFu3myXF3LjMWBrYTxoWkXxbCkpsCzAcu1gRAo/cAfP7
itxKRHbC830Mn0+2uTJyUDZCgNGNZMfhgVZPbt6cXTrtiEqAyPFVko8gkeXVknMG
ygbVFL7oqXHRD3avZ0DCPP2SP+6p6pRyKQGgBKkkKbx4q1P+voTSiHOkqL2akzxQ
JRIRASOZBHYjMZ9P3sx4S/pp8J0k4OBEJ/iltAnFQ45o88ufzAANqSPwBhASm82t
SoHiL5CJRK7dVUWMmzrS9C+jw4nLQbMA4N9CvekqKOIVB9VITnO6tlG6QOtUxNm8
aozOHEXnEYTV+9B32d+ZrtAqMqilyy8UmgUd5K/v0d3uE2KW1DNF4KZiN+AJRhtJ
SBSZGURQs+dMHCEjuZINLxKNOEtHNrS2QFL5ESypw6x6PsWLihPzwNOclTQkmBa6
OrTLroBPKcnJ5Hsexu7tVI7uVfb5raVqy2dygiDzhBlFjGa9ru5R0OHJvh4pml+u
O0xRS9Hs8OJd/K2wx+H8nWr3EfLH+Q2rb+gunzrs5Xnw9+no3Z3nBnpGFcEQY6h1
TJ/ds3wMtLoXnP/bERtkMGwSR7VqFsBEVLCPo7SLbZXBh+pBf+ObJA2TbTct3/9F
b3kQzjlpbqH8WuwguLzhMmSckIOUs8CcKtFpwqCigfUDCoXWf9bEuEO3tlshYXBW
B+tKNk493Kv9Yr+UW8z9xfF6fDAq0rfSGeUXRTB9wpCL7jLFh8qcvI9A4Rj9ztlj
czRTqVuNFAitk7wOlhIbVSNxi73WGmJqNgGTTXz94rsTqEN0+jVZ43dIMLUllA4Z
Up6BVQ35+8eB1WGkHherJIWkJ3fkJ82XJuXwHq1suIVAz9OtYegUrb5M4QXJ/yXa
NIJug5LE4VVL1shSMpPMeShqMr3wFe5WIzrkwnA0JuHEGTsSGWQZSUXQ4oTzIe1M
m/BHgiffe2MwDg5uOfVFNnoyi2eUwpbjXkoUpnENeg/Cro2SfwlFjXO/2MTygYAL
4LjeIXq6OW1gjBY5jLb/JFnAKUhVDPG17M9V4VG979Snve2aalOJ6cDDc4zheVQt
28u3YcNCACzk7rkh6iRXdf7iqOMj1T5WNE76SOjCdP7Cq8K/U1BbJdyStVfO8b16
2ELAcAmVfvC++7RKfFFo29hKubtKax9xhwH/BMNMBozboGTXpgRHxcc7a+QbuUZt
vVxkWye15yEFd3oOU4qWD+GUfOFQCnLGx7hpVvqdOQZ635NQNgTpTjO74UGKBVc6
TB0jhr3fIC3QH7VnJfomAJj2K0WLMb1Cr+TTErawsKmRyS6GE2pVI96xF5QsyWMt
x9O575EB8cItCXOkDw185m8O9lryE7QB7r1cmSYvGYoaPWIoBIOJ5YOnuQBnMPuS
PZOtp05BbhBGWFtCgmGKXwhJE5U6t6gaVwIwtrpd39cZQTqEHLVvk/bqwcfbbg7x
0YjifOT2EQ4FjxvHPECx9xcHOtt1vk9PSS9De0VA5HH5t8VxwsNpTjFKcwo1S4pF
4PUdFixXAugcOVz08pu5Rzq/EvhO+j9IR5CFNKIcC9CUBvB6MFoiD+uLGfR+3/js
Guyi/JTS4a8yypAKiPgH0gP8GzULdsyqFzcT8rIXJ4pG9jZxZO3xAHcHRjWM69Y1
abxD0K3keOXG1xZXqdIyNWhM18ziiJrlVwuKJyRW6cjxBRmjeE4CjY+IS22E99Wp
KDNipf3AloLZAP7bidYpXIOj8NuQZORNxgkfMm0q70xuK96FbQF+O999cY3PLCke
IDm9mleWtUoY0fw85AIdD1rYQu0lM8XAfYaaSaWL0wGtgXPh2ZxNFn+yp4xHjt79
HppDVQBsx1//oELr0lfN/B0AbtRZg/a+4ZRmYgCD1n9mNzoA2X/OWsaiiZMdCqaL
fpAXajGOYH32y7N1BPxFXPrcbLQhAPF031vm+Lyfyvxj4PgF1soXGt2+f7Qj74z0
tLgH9qZ8OMKjUTzl7Lfs0pqOanm2iIAalxY0yEWjQprnXVBPnRqhYLroCN2Id7AQ
wX+LPJWD5yxzGhhRwB+kbD4KIrF7hf2jxrm3jpMOK/IX1whsHiT5ag6RdBDMQ4DF
CjICLIEzFq/r52W2BqQu4ww6rjFIVGvCei+3DCcWv6ghaWc5616gUuKY88bIMpwp
48OQ0QOzYLxhzEaCS833IrX+U82z1y09djIajYdqkSZB0nzlKJs/9+VbZ25/bPhB
uX/9uF36ECPECZHKdv+a+g7qskCOIM8PtQB1BQCzYsMN3JLnXdJh+ixk/2hQlr3i
2t5wcxdIBoZZAiZW4iVXN0B1LLeBOA1Q7zAQq4CkI8S7z8HTUH7onX9qM1Lon8nd
1imb6LK3nALlPZ/LXiN8Vd4q66gZMlQUKKpaAabaOMOM60X6Z3VRaFj6qQglMmNb
2CzBlqZ7kjtqdotM4VC/ibxlNb8D+ifLyrG+kaOrTLl98GEg1ArmwoETGmzwJc/c
h0H9Z7Ko1Ta+mlVzks1CPgSkN7FMcO/Rh8y4ltfXeLIbazsX0m5q91FmFFUle2vl
YrbIMZANWHLtafBUsREQSdz6/dI+MAwreU6S/gXfT2rrvd9Dzx1hSmsNb703sx8r
UZGck3tFisQJItioPvCjpSfdfxvHqz6qWuR4Ral0ZdcolG1p6fS5Wy2onULqzZsC
sxlwhRF1qnYpbJzEBSiK623kfM06aqFXtUoc3hXmytfLQq6pHYgzvFAKS5H5g2LS
5llxeU1Ls3dEwESWYDD7mEGsdhXpsr1D7Ic24ium4N9bM6+xzr9cgCESUW8d7bDJ
P0aEiUHhANBR0jzUpzQzOHZgMKLbWsEPGFHhNvGrO9suwMvV4uFg9tMLTEus9RZB
SoOJYLdtMi/pkQX4Thviu+gkpvHFxCpxTSNJTNE2cRfArNSR4ntEZPMsFOZKAl5T
8IhRFHCTS4z/+AyuCm+QnXdAs06cqr9OiKRNEz6FL0+GuAAhQYEsGzfVEdPLvKWG
9W91Fm79r+14XRH+cMcfvSGyQfTomVgHlS9Nq4fBaY8JCt/0DBgt4wgGR5hsOdum
D77bTTjxytydRNSqVDATFPxFpgv1hL92KYBVHqHX+4U7/XO5BU3nGV4SJZeSf+vv
UT7aDE3g/zw2Z/dFUU2/VNo05ZWvu261jZhOQab61ZP8E5lXb2RTbSI0zABPjqCa
53S7G+5KJrs0jSIMBrIWAQ8WuoItW9xkvw87wgfZxaore1ell3jRxiVsQSKzagn8
FlDpQcJVYvImZQmoo/WUk+2TXIaNvFxgMpdmXAdEMLmfcpfUFUgVPkjcIRYpgEbr
L/jbiuUrJBVd87B5ObsCabXBwVzStNko+0xK8iOXjfJbHQrF1AxIHaamCFhQZG2T
HxJXQpT5en5xDHSAwgh8OFXPFPGvxbKtYodiBSLwj9o7Wb1dnub9dIZ038nYbLew
ftNkjNFIMqDawrsPaQjEZ9mBwxlhjSUBC0uth3yhi61+7K+w9P4wF/f7zZUyfNM2
hwLuwJ+3or17fJG3/Znh7JAQNw5fujNRDgFFYQHOjRsGwhhyUooNuYtYmmXByVjB
Dw/3YlQatm2cGLZELJXptvI3pkHgMHzaqQ8bWSxugv91NVOsOgFp2pQx25iFnEgt
r29t0YfQUen/Gv0uGPEHWTlDjePWQ7xqmek9obvPdr9aj/8HDnvo4Dkeb19Z5Nx7
Nni9mA77HupmPKeyerBtWd59+35pZkBC6S1hl89SAlvhM4wNSYd2NRAPI5xqz/op
A4i7zJAQiDEQrKtUOfPxeOOu4C54gUfbCfKJ0BX4Hkc5XJgGrJbC6A7tep5OSLLN
dJQKj4jKv2NdcXNR+JWdEKRuvcCztL6c5eu79bb+fMS9tshASN6sLZ/sBmCk7gU2
NfVfuvXvaDPCfq5InD82SkHVSwoLe5g/hc2GXJvuaL/Q5izPRS+tLsdJQNbfRDcU
iRZ1YMh/+VsVmT/3byG6o9edUEsADC3XiEIa7IAX3yE+9pUAaDvwd7+Sx6/ZLx3y
NBbgIz/YZQYl1lusYRFzU7n3ak9qOcTmZDraT5vc1HHPgCSrua11ijtzr1Ch64av
rxjCD+GQBtt20YI5p6BynLk4uLBxlpattEZiDmjE80F5ka8Eawi+ttkOMv3tzEpM
seY8uGqG22bxODVdBjoX54P/cMdD1DZg0d2fhfIT5P6olTy4x8cC7GBC7JI75ibL
28glfZA7iUfLPmte53cFi/cXz+5bueTHW8V59zgnp9qY0uWhWVk6TJOe/i5rgk53
gzX2Rqi1g7ptif2Ggc2xrdtJt+Q/HHA9RgZc/qUHps4iqmCk0FR+cA19Mr7uX574
Q2vwxnCWN1y0G1VtOQ7G1V78LhbaGVDXo/vxAA0PUGnPrF/NDO+SMzd/tthu1zs6
JPd1kT1+0brI/HgGCL4OqFmT9lLZdYVoRMiU6mjB0G95UZ5F/zkkqVJ4h1uXillj
nleHixcS4FYEYeLmAByWS45/Ws0zNLoLEO0ac53bUNYbp9TKPqxcoWD/vvsDBN68
kvuhTZ4Yx5IzZGxcPDfXh/vt66G2dGOzXZE+kjbp4xGF1DK5uo4RIkpFBltH0Tls
kfBDZLPuqeb8xsHHgTL5He/wBT6DvrMZ3o6LrDQ3TJQcKtd+7/58gh8OH3ht+Cs1
FtmbfhwkP8dzcuxpG3vP95d+f+1zhjbPQRJFPohaxMR01y9nwhPUtWLV58a9n0N3
aLpYI7UCeLnafWwFq79g7pofzvRkoYIZ1YTMabI015z/5t6CQ7QiqWb+Lx4w7kNE
/qudE/nQ/WDOhhoihVgJfmaSSAiR/GIFL5auWhsr6l6nNnLl9RcsVwXQ6Q6GhOxc
GWfXedQbPz0Wvra5xiCAhBL4J1hAYQU3Y9b1Mf5OJrqXKA6FkdnB6lR66dEPRxSZ
x7+/MuT7BQYT49NnKpx3wMSkp8gWiFV4kh2aybXZ50vMha/ehvy5gRcpzl7zuS+R
ACV50IKQqhw+1sIygBX/Eyp22u8Kwb35+z7gl0m92cJwYgUtuYnH3y4t38YFdSGO
9VufOll6f95T2rgtHGU6jn+R1YDnfBWjtoaDaqgrZNi0xPToQJjDIjXWF0VMYTuo
2mk7Bt6pbcppf5K70xL8aQ4G9fABgfA4tNP5maTSMjwLCW1LomG+ucYLXVlhIyux
sNtQlG7aPtMVVazGHYlr+iNJskPwYEE43AVw/2R7Ey/JTCKcU+ja9fkge17t8OMQ
FrInEcBscp3sguwan0hgllfuj8zb8Pi32UZVkzDWirVWRVRBoebOrKrVLawI88B8
iMnd9NOOJ0SYW+3T+qYdAAtH1inY6vc1E+hsBX3ktK9LkDCe54pBpsJjiEpAjWVC
af6lcL5bxOBqMbqF0qGVwHcgiMYeiAR0BH579lsIPFLv6Jaf+H85tkYKhmPxBZfV
5pm9A3Aa6xBiFZy1v14FowKdCiqPDa0MwX2RA6x+3Aal4vgkIgKwepIVocq3mBg8
TncCDa5z2fGx1yhai55CmRLuW0jyYWirz7O4bxB4Dd/kUUqTeddGmc8WBKOIiZcR
ozBdFNMWWxzJOlozopiA+HeuDavlEKDg9Nir+82mD3MkhAaG0lTQ92k9ED8S7gxE
dg2U0qPGmc/GFlC1L8Ic8Bytct/eNkxODkiqgOpuShhrZSlGpIaR/CB03afUWhK7
2IyiGdUPIRyYzR6DZu/KXKe4O6FTzQRqx4MyP/M6BKArRcEf7/2dWz3aNk6YqO2x
Ac3DNh6nxhH2YdkysM3GmqK76d1RzsHdvudKDjySewKbIrTfRqWy4loIY+WfAgeP
bcQj5BbmdU88xfQPkKsFTMg+2nfFIz4HGvd3a0WdPpDJ2MLB+CJn/MM8fjJzyqm8
37WdOm6BCZbf71Vz6qg7Uy2z5vCrOgEtkWN7zm7ZuY6vpHyyusrIHD3a7mZpk805
jupUT1La4FofzqQcXT2YHUoMk/PIQGjGxgIEJzUKFspnXRCg59Pndw/CcyRiWpjT
PloykIcHeNR6+D3HdIY6Jx8zz0Lm6ROdMYlU0afFTVtGzVKr6wcSPfcz/mSw+piQ
yAjRj1ihE5mpyWGTWX8BbQegWQwR35jEQQ6t8W0qZdToUx6x6rv4fkOM9fnlPpcq
6WsApxkj/pAG1ZKGWX9VJ7uqg2hBESFtd0xNbu2kQA3cDYm+t/oiyFfB/tq1YEK9
kOrJ3zR7QwJEFqOKwdnaAlEtduI4phEqTYleM0ANkh3SEtH49D257MyrBmDiE/r8
Skb/C5sWBAmiMrswvP419/QSP1gNThgUjs3FBIzix7ehCvRTVVEUz3WYMrHfl6dS
1izarW5WQMy+14dNGAHx6UGgQAmrI8H2Xin/coC5uAWWUyA5UUm9rB//nsjbRR9b
x2rrl84wZFI2iuifsneqq8Edcbe09iZCB/ReUbcqe5l1Q4pfR2ON6qJk/YL0MVM3
Dw7kIW2DZEXBpv6KXBtJZjUfGC8xmtrwxqvGd7Uxi5/Z+IR7j26fYjpn6sz0ahUE
p5sUunQnfgpLwjkivVg6I4yoyz9JoJ3q7kmjEdRJlRbivQYpWFqQ0kUt6tb6daBg
20mthLCTudgv/rewkoVhdsf+GThR47CfUKfbCRfQQlh3sC7w/exzzoMmwegxZwvG
iGq4QUOGf0Lkt6zWS3/REfidfGk1G839WL4lDEEtwtaZoNmXYm5NSlP+31T7Fs9H
PYAZS1dVa2FHdluk9k/EFm3P33SYQMZ/cv/yrIISfAbVdy6bcbiHGnnb9ONlkjdu
dYtisnTtqFV4iMsssoSBsiQ5colGXsp1GXxgE+kPOIPXvc6TlUyQa9CRSbAidmD6
2tzBsUuge6n5J2huxbwpxfh3hqPazMLbcjh0Ayez3iQtjgpsoZ8cyPgB77RZggjw
HR+tpG5cEZiUK9shUieuBFqQf140myo5WOK3Sq+khRV+4AQUCykXQKACanq2cx4+
RCNK/JGMr7NBggtkYZd7umUfHgcCMC2FVfj2OSeW6JS4NUzjoqGaJxvZB9J5lIEb
m4BJJIYMlnYV/nIzGhrp0u8zksBFe5KhuB+WYOZQF6u9muMz7tfq/ui0MwBiXyns
GJxSbREixDNu1tRv/+v3jW0aCZs2k0L+uYDm36YZg89iRtK6q8CBjeCdtFIZj8og
9ZKe9O+91YQdM5SWihqXXBhOPohZWjqltGAfeTCfx1OQtkYzG6UrgXQiuG9LC1Lb
25+ai4THSUQtwgz4CvepLdgP/BK2gZAQ6m/tP4dDlVnXPbqKoUiyP7yJQ1CTo/5B
ZRMZ4d0rDFU8/JWuWnnLhsYw7ogsfjlmGbtxqdgYG61X55X+KtNzzR3AXwQ0HFHC
OUDx57SlgI4t+56msWvW0EBw9gOjnpyNeEdSgVsg5WKwE+liMrjxia8g5H5gpx9R
QrRglcdK3Tmyyu0GJl8o27fgRed8dJmsQW78G5XGkuDrS0RGL4iPsF+lchGlYA9E
1JI0A4LlLzNKuWJl/jwz5WwaHvopL99VaWMzoW0h1RqFHcMsnKYodc69miW4JTjf
Cc0GhS4vQwTCrtKiBdjiqn/vQgjSZWUq4m8jz7Z1z1WziMslk7LEyQ2ukPKTE9Pj
n7aKmBcElxPLAjo0yvIpbas5xuiYRRBcHXKxukDz+iqSCiqEegssCXmd2E75cjDG
B6/pBvBEEXnorJujqTJyHLGMcPv4Ijz3Vd/MM8hCkHYnxQPF7btv3yj3zejlvuui
HOUUrCT3X7mbPWU5jBm4GchcoroQaH2sGC+ur6d+WPaM6mFCtXEUCcAKOsVnpgkF
EeDFOXulXF6RlJMq+/ye/OoMuM6qanqaTmKrYvTOWcRH8xItav49XIlejJqQU/kZ
ra5SZt1NbVHX2tUu2i6EMJ5cdJZU0N+khY4Valef5r3mmghnkL1wFrdDFM6DL42L
gnMl2iIJ0yrRVTqW2i+lzh+bD6aiE8Pe/FpWXwrJdgPBBLh/M0g+8yNAYA1A26Wm
00D7FDLyNwYjmgXSujQ4ZeTdPBUqEgGvhRGpOcDSswZvO8BSjPwlNrqGRh3Zj8+h
MgVXs4FB/TGsNq6+JKs5v/r7b16RISl7b7FwZ+CUsIa473eG5EOPVwwcYE8GZh3d
Brm7Ey5veJRXfCqg5viBhxFZwkQzLfDn49TCsrv5ztuMKQatRj/+GAGbJ+LnhwwT
nNjwRJE1M+/7HJB7Ygf7YT3sLSGlqHJ5mYUZmfmBOUYU5KH49tgPaEaD+agBBWWQ
tPplWYb1jC23I9Cin/e4sjF/7Ba/GNnvT3m/v2Tov8D/iQuKMQK9lD1PxxcYSlMY
mEj2utzPBk3t4h2L+VpJWylb8INmUucG2e5L0nPcVjSNOu55GRVmQGrnFJu/z8lY
JnT6EaELxWOqgF6oDVsCgHsbm7p8p3oGODVGy6qFC0F5pxvGUgTFT3AUwedoxKQt
WCg4kkrzAROE9qXSm3YVi08nB9hw4dOQh6M+8oZPlUVZ7TVKDgKDC8t6fm24n/85
E/9xLnjdZEoJtHNT7ngk2voMLJplqFsS9/C7sa6urFyI1HUiDmDDy3a+DW3mnY1S
peWdEQwrv/5vMJ8U54tfsV+UourSpvtVoa1U4n8Oso/n78gB3AtI8npwZjkbk6YO
qD2flfKMRiFyff+YrIV8y4tqgqUKw0sKePhg1iZSx9QsPaESJURB8k0uOPkCw0LC
EGGULgOhpt3ft+rsLcD0KXo5/Pbpos902XTp93ISvgsTteRxlEllrt2VV6+aKcIT
pcOdTIjsWoCA/X6pASlB2NIRBUb6g7ZXftygxevHRofpu7tXvgICO3Zfyr5CvtaB
9OMRiLePzmTRCfUXGZUrxC+p1iONiDSPUx72sigCPbwU/wDieaq5d+pzjojcYW3O
E9j6B15LRLsKr5WCj9WV1w4Q2HtaoaUQblYcYTI3oFeoHivVmUIH87B99OPMLJ7R
OlreTPKCLsX4+bPtYMRguxAjTzacG2T6pC3kjw7o0UKTpMXIQPXqVHfIzipeaNs4
/9iGiJcKX2kishY+o5J6iQyrC+o7DkoUM3IIrzdDVM4aauKgqxgFtLahHyBOZAT7
1oGH/tklB9YKazGL4p5BC3NkueBl/s3BWc81f3oHuOSrqAPF9+M08HD3wIliSPZj
D3oyEKu/JgTcrq9ILnM92z1ZjRn1tTY0duWTG50Y5GhEw8A4Vrrejk9l6vH1/eBL
zqzW20jbm140Rc9294dcebxzL8uGoCyWIwh9UFO/b7WJbtH1FLGsRyOQE2+hYFfI
WRdip/DXEtJDCI3QQAmdy+ahEJD+yq+KRWIT1mInhBFty1gzzehlhKa3d7ROGasp
n2pw9cQIqZgraR2osyOGLhCmzcjQLmZQyCawYuHaNkYaAnqjQxUCyuCB2kXbRrsY
Cb/rr7DUaX9n9OzD3nMaXofvJnyqWMXbjw69+J+js4dqx3c/JRFcFfVlQal/m5aF
gRLJOq0sWZrUde7WYURD6QRRtJqql/51JCT2lNlkkeFISD9jD6ROgrAhkwIK3Lqi
usHblyA+CUwXXc8CpTlgsTHrRVnQ7QjqoOagWR78/NBQQ5Wlik9MCYfSC+WZPF8N
TjRmlel3xlNF1oP+bAxE23lqvx0z3BJ3UMXU7bcF84imFwwacfBxRGRXQvjc4u/4
YwzFCpr1c7UIHOawOM+wruEjWLtQSLLOenhiBT6GAcoKrNr7g+Qv9snH3PDaWqxc
/Rgig/otG8x7hd5Gdbvf+9c6G0zhZz2JVEoFcnCz37/7ABq/lAxBH06AMmDqTrM0
y18CuXsKq90b0EkySvKgpwT8lbHXbRKKWXTvkYjnXjXaggMueP6SbaeO15yDM1fs
fjEnrN6k21bvdR2ucTR/4IJ+FxYgcUeDBq/XQTM3H7g8XjUHknM8EChCjIHWi9u3
eSi32VBmAtkhuge84Kdf11DDUU9sZzBCwhcuiZoJoSTvqeu/s+jjoXcfu9fJBx0w
m4lwhHwqWJxWltsmVwoe5fPSb5ddkbDfINr68+2dbAi8Bu0KCV21xRsuTWq57akh
aYdvLik1hMmeuwdCxEEzQnYypdeN9t0m6IcYLrxZzqVDSmftQU+BRiORWbN+Z6G4
yih+jy4AQPYPeznFzwsuidJoIicb/03DC/ubnFCfUK571w1hLmw5q7VdGUxx0Ivv
z8qZauyne0UuDYE7KQb7Gf92K/xQCaeYVMuR3UrebBcklr3/LNTFxPfiDzc6jAVA
pEb5pt0Py590bhWCr8XdOPSXi9CKBqY+8hvyrxQeUnma5ijPcMiThJpAIsrun9Va
zdcuFX1/+2uA15JXqm8DfASbSKtu9ytASwBIzHgu5SxVmcWHO6AUswAiCxCezJIk
jDzYsRNhxQ9nbIqI/vnZS5IdV1zdfAwwjXhdN/VQdYFoj1uA3ROJDUBQgil2Re+y
lGZSWbku46jAOIY1L43cnQDn4RfigTgaGoRkiym0E9kTNwsUvL7phG1Ooinyl25P
KbDoDe3Q3XLPW3AEZJc1TI33ECugNr+izFwGhggjICJRenNEAnvZJ4d/sRXebANS
kplYu4OwDfcRV9xQaYsb4s7doPpifizUyUTMN3r/cWBb2sbWjAHHn6Kkowrfq29F
RwuvHrCIe2IGtXHXVvdK+gfjLSmC4Kfk1pF6gT+tcR960JRe7Ky45kdNnHqw4sQS
O4zGr3wlroUCzKPeipdDdoL/E0d3HSXUlRAo7RvNX3YS1zEgZxa/e8plkYjBQ8Mx
PU3UgzlBCKb04TireO5UfOEw3g9icy3LtERdATiNwQgsHtlUUskFLNWDpsi9V16y
WGXeUbVwJ9njDTsZIwf7dFo83eeqB2q294tRPdzowgn9MlAAe2TFvzzPpw7aHBX6
3mcanjV8ewa0a+5lO/OIJzNs7MEDCsxa1sTDCy9tV7WP8Madv2RekE2wFRH7thuF
sKD6EU47rznw/ROj8DwDrHOIkqbDAo1/R1+o5+tBAD4zgTxoi5xBfTA132chP5oE
mr8zfjlEoFysgX0408IUmleV0xOeYBBCcM8SHvOsdM+2O/WKWm9Upk8GrpQeBK1n
Y5wBH1BPn5Z44lGdJMYG1VBIbX5uXrrlM0B1E0wdlTSmpaTiVUaFVHxkqLpGIgJq
YAsKXjHVD5E4Jb20Yq4rEIwHWQ8WqXc6T7V0vGKYBt9mvFG+ejp/PjbMQYZYDtUU
Bv5UA8GTwozJxqekTltwPEP5OfGXaxKyzpLUvwKGKaGETSZ1wjwg37fAtKUtu1nv
xgp5OB5oh11WosCfL80sizQxI3Jcvkl7SICJef5MiMD/eTQPTgxfDLmPwfLrhotd
sKCsZTmUiOOhIlGhobPoPaooCmwv4FeLCMGreLrA2cqIG++cIhgyx0Z5Rr6TaaYH
Ndgi19ewAlbW1g8SAJgbBmc1Np3rcPg5S6Od5lMqOyMDjT+hnQfd0qHv/A8RvHH4
Zmd7EZk5FIZUx+vGBxzIPT2xjFt0AeoWVYBX3jwMVsB548JF2Gxzc5QIFF43mZzp
FjoHIQsO9gkFlbPaPcQEbpAlO/PdykqkKX8MSHNPHu6wdHkuap3oD9toMWhM2g2F
DIb1BHZPa1MU7EzEMPRKO7/SC8BFCrueoNrqlS6U1xIN8Yv/+nWpF3s6J0APOCad
NpNpDBxpXakCibyBMEcQOSraZiGk4vJ//7dAjrAoLJHNkSw6kuGrzu+HTmm+YgwY
CmCJmvv4PsErPOVLl/cmtfXoAdFTzsfZfZ7ajkCOxehPyQDNLaGlcDemU+A/UO3w
kEg3BLz7Oa1hwiahd41uTxjDERrNEdlbIxZuhk6ZXPluokwPtF4uNVsC9myocMHp
uXYnBV4ihXwPPpO+FHzPbMob2QlBYzh4kNmEGkWtjfQuzEbBE/OKVs8tMUvArexb
ERZZ27RqggyiJ54zXUR7n3HfvLgm3RSj+dcDlTiOjOjRPLu3qSAB2PzCaT0jlkeE
UlhHZA2EFMt7xugOe4HF3mU9D9r3bcSguo6ivP+1EKwlTqdCKoz5Sq3Q9gaEDs6m
Rw7j6rqebPl05LoncE0F27jpFQdMYoPMkBUlTVCJJfFBJRZuzACAu7DLl2IiTi+r
EV1MschnRAxsHBCmf5RTlspLwnhYpZDWeggY8MT4mawGW/AnJinsiIYNGSVUMmr5
aZHmcs+WUDlfXGpFisn2Sl3tQN8kGmMUZLqBYkYR1FoGM6J4UGBd5Xg86sRLz1w+
xAgRu+Ltx1RoVn6HC52EicnRIBWHvthaLQlX+KgidfX/2wzg/aHS/iTqAbezy29I
/g8mZGTWg1m2ySemIFnQsTHhU2CEUb/OEbjRIBA1aVOsKLufZNYbrVtlE6kFQ/2L
DQ9g3Bn0wfrv8Mwu+nffHoDsHKmbLlFf/fknej5/mWaMCCink312wWPmOsxzeo6U
kgSwHuLdIkn+qdE3QiXdgfbSaQHp7wHL/AVN/VLDRpdwdUDMKk2MfQqU6Cjss+pG
2972VgeB4xfj2iE+xOMhiCaVsx5DgE35LfOhAatwJkp8NVCjYvOzXM4FJOsisMOG
fYqhJhjBoXEFw6bVLkjtS0EpYTODCd7wZL4dt7qRGNxuQVC5UdBbTYEzClP72Ls9
EFMKYE9SCflAeHcJ6NaW12ANe8xrmcSc6++HBa+qgLlzYUkyaC1j5HDAhOEBLX89
JyyzMJQQHCYdMzw7RCYb6jllHI9CpT1/kZrD51q/QgKHCGZHuDhj9Ok0Q8fyVYJS
rj8Ycs06A6G0WHd7NMY66zcecyVbfQmRvknbvbBt3lQSUwLP/3TXFeRgiwdPEy5M
5vwNYkDddNkTOSogpAxGNO6FQ2XfUmfTioaRoyZbh7UFQ4z0BLBSGFWTqI384Prs
HxAQiGEraP1MTNNKPiMlCxCoX41aarwn5FYa6UYNQO0hRR42obrMyvTngx3ZgK0P
8vWupN5H7820/GscTpQvcmlY05EhZQiCkmR7+DxHt4XVnM5Rx1O6YuIw2FPi0cAV
fCjIJI0OOCIeeEhMwOsEPRgMxzKtd5B+4zYf4iH15efaUpoLA/CzmlH7erOMQeQH
j8IQyL+3AmkFJYUy7C5NTM/YV412scKeox92YXbMXm7wmOGxHZPJXB5A4FfjVmJD
OayZUZefLk7k2nlWnCveep8DfG1vcpqr4AFsqjwNWS0Y8/GHt5ODorOsdVsfYKyI
u+X/g3iG74QFndZmg1HBKySW1+ENa6Nmi5KjSh4fG6Y4nfoC5gKc8CXzUIuhPmX6
r/tqYhIID3XJofPyUJcJHs6ucmoZw2io2AIdUhcoAT7FDFZePvdh4M0HydfrtdWE
6/r+ni4TZz+sBJkEVPTDQK1x2ooiLW++XbIETEeMAKvNTtzCEE6XYAFKBVs3U8aH
ifC9ShSXo6DMknWB+vGRwudtb+nqZRk55B8cUNeHZJKTiCE8hnbUgm+GIBEPWfx7
NX6F8M26NSZHW1cxbkgldSOl/sg9T/Ra5YuM29jcqQC9MWnPxIIAI8UAz/qVRjn4
hdxgGW6MoQ2sw1L6eos0nKH+5n8VClSFYOJGuinWGvnLUsiFEeTloV2kv5iqtdc3
7lM3sLvr1Ak6HH128DzKy9QeqEmDh79CGdusRmDRjcfMc9MmIHc6fn2c3UQH0G1G
FPn1yIpVQfp+f96c49SpEwoFlPpXZK0+0PTYT5+srdWfCdw01tzw1zK97vfn3dTf
MCNe4GHaB8o2X//Ahqx2LG9HziCpmmOnd722acNKwyuice0pBq9ptnt/Wo0PaJGC
tiqu1x8DstUWc0jz9sqMEy9QRH/xeVU+G0lWZSeJQNYridMDncMkhp7Wl3OhsruZ
qyn07OmocK0A4e6tWv4IekPPZdEZtVIDchIUXrytNTNH8+WLJySF+EGPmMgyC5J+
TPMT4mfY7DXWH5MD8gimw0T3iAd1UZs0T4VV3kRD/FfDsZ5YD+VNriewT9kdjKAK
ZtUou+VUPHWl35ul6dPvyd/V+Y67enDqnXPiavhtI7gbb1Ez2VB9UbajzD73VdIH
aEC3tRkabQumifUQfv5uT3vs02g9+80r1bQ8EX0Az3dZsPe5dXEqtS584irVSz69
DMCidzDtKi5N7PcDVJMa21h6TLQapLK/+U4MMnezIJ4vBgTTaiftzF1vWe9o0WBU
Rpr7t5G5lvQjTcUblMm0LKEnho/txqpb/JyH9MOEJCUiDVKIhTZWbrb4ADnh5ZMh
leRfRrYf6drWHqQR19GwYH6xfnVOqva/E5e08v2UeRmgLWLeK2Dg72OO/kvf7YyW
K5ATMJDDuS9F+hahLA3UtrUSrkm/RTPdQgQLIrtpc6IG8a1GD8wVNPXbf/hvFtHZ
z9niK6eLC7lXvnVAdZ/5Amy3t4HL7CMDG3nAZ2yu8uL7g+yZjMzyWusohPVeWC1E
5X2p5Kj9lbqjHBiMoACI/6OfY80sKfVheQWvMSLjUui19OmP+n9pTrt6QDkxQKjF
qlb6UZpXpCfQIxBtzTgTyrDYqzx9ldQa47FE3/2TkV5kAOEVDeiN+rInnI+bXLcq
S3zkAEo6HgJRCTfk2p4zGEl9m8vFNuL/U4Ne7qeaALIAj0TRpQHmM3uRG4YgQa4b
FBXdnYXHOniQzIUbjkB0FWrIh3ZBJGe3/BrVJuKhLfDoSN2gf66Gl5K3xUwr/adb
0X2y6Wur96e3n2LSzhcfLg3UZf0WyOaYjUoUeArg4kcdaDsZiVi4B9/59bQ/WS00
4OwV20JF8YihrGUGCKdXomz07+SYxS9NsgWTYMJXicTo9iZjXTxS+SIobUyW/xVz
IchZWvuBRDsFx/vQQ126xDX+tR9HkSDpCqen71wzhpDC0v+AKt6etgX/qxlcI+d3
Zd7nNB1pJT2MdqQfTFQBfYw0KiPLlaWFrKeON5Q3y8zo8kNCNjrcULa2argdO00i
zG85B+EtgdqjL91K6kmwFtXewh3fzbXnSCTGnQSTEaAOfSoD2JuC606zpuWCUa3T
ncMa/rMYdGF90mPrsCB3KSY5xek9NN+3Dy5UiQkDTOJEfbgC9qgvsLV4LUiw2g7c
wZ5rzmSQ40pnEqrucYbPKTDMvExa5W0mSUJ6RM5lHl/kEG2kojj7i0+3bSFAD9+C
qLkSkDeRjE3/o999Ig8gLp7GHb/FdAp9DglFZI3QodxSN/vceeOOHqHzRQfa55yg
6ft0ReynAYf3mnUBmnETAYDZf9lM+AU7JJF3aFowdjzGrLnNGSPQkBYWeVse046l
jjGwK47bIXjkrnr61ebqZfnTVVcx9gfkNJOroPntrBccXP1YQ9DAPx1A0uROw5Fk
UXEqf1droMBCNjI3hOzrpN3xG5X56GT6tZ20BTtv1CyQfBpBcEBUS9Qbvur/C2R7
Ph7cxyLfy77HUvENCYELqnUIZujLENgg71ChrqsqPEH378pKzIRImqP2dYp7Ve9k
tCzMedKvwamKfTQYoBRdQzdonmHo0m4ZxVfBla7AhuB9BpCJ6vWpt0qvJLM3gJuH
K5c8bpClkUMIxEkd+Z0sqD29KWj4N0rWoYtRgeTiJMuD0aGiPHSrwyP5VI/oHuJc
8zgiK1k2YwTGhmgNwuZeulRDFECnGkHhDBAeqIGOwaM=
`pragma protect end_protected
