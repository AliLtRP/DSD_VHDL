// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TZqQNIG5uUkZQ+2ADl51EMWgp20rvxkZWTloDcvtlBbenbj4ESFdImRovbGpkX8E
npagUDvcZkULVUUu2rPKvA82XbI8/aMnwRy5FgutvbuswePSxubpfe/tX0HdqtIx
b5r3U3WIIGSSrysWI9+5JiUSwcf720Q1qNw4u/5Jpus=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7328)
lyRU/zT1i8ipyR9rvf/bfFmDagCAX05nC9aaZ8JaQkrtjR/2UhnE4VztDid6PMRD
Ehp6WEsG/sUJVarhdLYvgeQ6pZX8k8k/saOrBxeKdMuli/l23qOwX4Q59qLXDfsS
wO92Nu2jKvCZ8DsowqFiKHGt9LyPgdaCiit9X3qst7J4UMc4SY7g0AUt3EdHi3MI
+T+29HMLER5W2si9KdXe67nS1rJoy6rzQRDxfCxMbRHBny4Q2UNCtYWHoDKg9MCe
yAlKX5cp/8gHwnVg1UbKEX8VC15uuLFd1Wr0pfNENLLg3zxpd4/kAsBZblNCk/Ac
rZfZb2gx4UwTwKNQvS8vPZLA53xRVnXW36jABCYqICJ+EI0kI6/AZGZW+g2dPLA1
5bGrQEL/OAmDoFeJB0nuc6dlPVkQuRbuOMuDkVlSJPWmINeVTH6dvHCLB/kzEnBv
39j1ERAIJo65a++FfFWJcQMR4abAzMtH4KQLW6mE6tj19aUpZPQ8KJ4H/VwhZJYg
r6wTdTQLbYy++rp/OF0aS9exZmnQ/PpVAXT0hvLuUjTK1EygXvNsvvL4Lwf/eXHW
cuuaXlwxKg83o87AaI2bAoxD20gkiA01Kec/3y0CxAkVO4D7iCCpRgWKYCh1I4RX
jKd6vXX9CdIwmePwVyreZXlQH3JQV3oLzCw+j32/O8ybFZEJEtwNs9T8rUmP3r77
+jJhCu9N1UTvpHJXiefk5jrORshnaJMHYTBf6Dc3xrgayjM3/NmBpffSZ4rik0sn
NZ1L7+WlFd4kVo63QFM18GTLZ9QM/5t5OFma7SDraa2s1Pb0daWVgJwYW0wz2HIt
m/Oa4+iVtNXjbZt7bmQUHSNXYIF+Ha44pFCTA+baK38hP4K5hXqY/WhDYh5vBw8x
2gLI9Pw+xnuic14NAtcS/zo7kymMIJFW7UAdmumQyF5U3NMAvH5hVDMYWmVGXF2e
gNFtXXkJBL/k3wJp87ys9QE1adX6/3Uyip5FrsLio9fcj2Ceg6llZWHzxkZFCGIw
dKIdsLZ2N/Fzs6UtI/6lTXEfEYH1TLuYI39Fht8e5fNOWPkcKg/t+SC5Lk4GX5kw
0RAL0KvlGIoDNvLFxb23Fk9Ks4ELDAlUBCqKap6m3NsMp3W+u3ruDRS29Q4siCdN
Zt/ieuRrrIlWqeVF1Es2xWGbkWD3Q4mlVw7fUJr6LJR90LGEzEf+mCQf0W+an41u
0+VlK665/UAaXm6YgHpqkIWJgNela5XZsKpt3b8Nm+PXXjmSC/f5wBxZL7K4pLOB
a/83krd0rlD9dhIBV0rTQbFIWtOFUFSe+PtIQ9Zky30hZZuTJjj569MfNVtXRbvm
7jJhOtQPOU9WebATHWQZoPhtOtkTHVehGeotUE0fVfJuNIXtFxv24V01vgbnFlGG
P8eEHSvU3jOkivrtirpfkHB7IBKofA7qz53JqQacBajWIeOBkp+0B8iSAGxAtaG8
WuLtCp44/1E68iT5Ava8y+4oXwVJQqZ6A6bB+SmBGSU5y/BUhpPsI70jDAyj5Bo5
HIf1EoTmfOnNAdk65pF8dwKHhaEikMBaBvQTmERYnS/cluU12weP+ynAhgFFlu/q
aT5dxJJEbYYGQTO8CuiDTIIFluXYc/q41mVS8goWRee0JkTKKdOcYS7nSwb6bd4p
I/NFa6zyzeYSr9/Uqr2AiE68lCrfMajb4EGms9Oc0jve+X5Xh+XJpKtCRAwKBo4o
zXAVcAyE8Q5dDfnB2aZI4snhs9f8HG0JKmYWcWv3GVbmOu6pQrBjhR45edbCQHSd
GcY35WfAeNj6rygmfD/cBSm7SrEOUJ8lz1pbHj21L87ontnh8S2Ak/saf5cQ0aDK
xgNhkte/YWxktkYUnxqwn3vT4srjeoWuSSrkL+7vsVo3ugxpUcX2MbbxR7meIEji
+Ht3UI2UMpyixYA1Z0J7EFocROp5m53coWTvPiEyR2CNUtzJ+kFk7tjVLwj0Xr5N
0Bd2T7pkUcxnyGq5GBFSWMRyFuiNgEy29yfY19Cmq5sF3zdVTIdgWFm9IQW6Qpfp
LbKc8x/CGayQDNFNupFqYXuyUJHZX+6QEHHrjb32Q8PP6NPsqIymexhPpIa87fFl
V/ivUuhbq3R9Q2kpl/nMoUPaM9rUPoElmvxBHUiPhVXNWSJctuE0mHVdsiDAOvtc
g3FMku4EUNDzqOXx0ewdaRK7eoJgf77tthLKk9sx0Nx0u/ExmJWmCXeKdG4fow0y
V6ZamhzZFTc+IcmKoYQVeH6Q0NEe7kfZvDMPhOh8lHOMkYZPnd5ag0FMegIR4ZO6
d1W7te3y45Hmz7DqO4JJhrpcZ4ysx7vlHpIOv87Sbs6T1TQhPiNQC7DDFsUPMBnn
vZhUfU5oB17mZ1DG7Lw/re4qOskZObmJTdIqf3qanR8CylJ2z+ZnjXBaGYvwHNnP
iKCrlHjsS8Z6w0SygAYHT8loEj3OaZoGEuqupeCtvKNv9GQPdt78OTbjfvnFqMgE
EgfOopvyCObZ15lHm6ICWl8b87Xy4CARlbfagskjuWmX8VoP8iMvFF5wgayrqG4X
2dhUuinCK3Vmqlnbyw+DyVpmu76yNWEu8ZS2OG8xCUsyUXVdgH1dWcHfQPUE7lbA
6wxL333xKBbaOg2yE8c6anU4dy7PeCqU5NDwmZc6lFCPjTvzb86HjpQhLSWaECim
kbaweLlupW18kJ8ux1k+sPnu/UnviPhXjOp/ASwADNcVGU+ORarHfzyTHLY0fV35
MsKQiCEz8eeuH1Sb0Z/E64mnS4ZEcGBWxN5uglEiMWcAG8CXybYlngwP0iuWYdZB
X2l7K/7UoZdayyaD+SgUqK9tFMIfvD+R2grdQWpSC2xhN589tkTvqb2X1bHvVHFf
Ckxw3CIEQasHdzCFR3sDRwCD5pknvoAKstqdM1dSZe/MGy+JknqEpZ/QVcHghk+A
lJl3usBgGLIoCG9MCR2dVCyFjHkDHMdB8rE4Ly8hXQWtze04O8OtZ4LoA1XWG2pt
b3LH6C4Xt05Wi+gL8Aent7KH3++hICF14/R/L2dBvIP2GE4fqgMjtiuQdUEEJ63h
AqsukNEFIBxt8NT2nDhqgRLUtOj489wDVHBXXC3nggGaqtdKEhC84RD7pcxMB+d4
kVvpW6ZCbMfHfA81G8MKzsT4PmHP3Vm2U+jDkPkgijyWL4lMAQdhoPRCik/zALOv
yTPDSY6uLzgE09+jfuwHA5CahdssJrrq2aAbW44PcNqIQsqwzfjLRJTKdgsXZsEw
APm539AP545dUBcvXJmIwDf0icYwjbYTdYvTqRyPmonk2DZvBWmmA0XgEnsb0MZs
1Bgv4K1ejYwayJTsHPDjheAuMqEgZqe0+N4MlgS6BnOq2gFrh9J6w/OEXeN9BiRV
7Ei+ERqY291L8DMllGpHoMZslfpMgr0pDVAjcDhYN6RhRExfxPXNHM0Or+wQucSw
YTLZJc6O2G+ox8Mx8SiL9ceLsiktCeXhctummZCJTh9vHG6/loXUyOB1DDTcP007
8LPQUSLMpmwL0Yf08gU4OsRhoznfBFJi+/zUmas9ZRJCjLOgfyb+YAbVfmsmBNIf
LyIHewHRRidsr8nupeCpnHpNbrI3pmDTCDLTZH/FL2NAfHzHhKYm0B62BJz3VtCA
f36mn972ZliQA3G/9WNHQc5vS268T90n0u6sm5oHkVS31i2m9PUIpxnrc7VSRQVs
boAH478JiG1vwpMSbCi3zVOYhOPXCWaVhSDhfYCnVx2howFSSmEuZORAsGjCP//n
KGv5CNQ3dXkljDPvbBnAUDkf+JFCSObbgo/9SsKTIXoN/lDpf30GDmQz2+V3vRr9
2uKsNPfIrxEUeG4toOR7e9Ltw1EQ3G8qZ8dc2G3uC6bKXaX5R16Qzm82NfojAYkP
H3+79r7BnTDYPLvmiLK2cDr9bokA+BBIE54PyQr9CrWZvonha3MdiEhbK4a+eyga
/yoOeMtMzlvcUDPMQmvTLvRqhVfM2NHMzDY95mrjzjtyOCbdaqOF8QBUDSByLUcT
lWONI6IpGeCt35St3kgQAoMNpZgDxdba/veLEsvOB7qxB6UBoyTu9tRj3w+ARCUP
jccjSQetgFBRS84biyqmwDHgpvkCjcD/u0mtW36gvwZ2Zpx82CZNiwGMsCydAJu3
HRB+GuBOIZjsiNbbfvnhWg6+rIW4gH/ao+C1dtvbYvFB6Qgy5L7JH5ZK38NH9Fct
C7ri4cchH8KC1IrIOwHK0/DUgBGWIb6/7GQ3EVhPo2U/wwLLTsVTMeKP5jqfMthc
kWcWCy7AyUJID5j5VxHGmycAiWhGsf04+oIdcDtMfpztI8sDb7HFurXKsCoOs3gI
BP6JN5lX7LXZbbGOBcaR2lt61ybyH2dlKW/qt7YuUNImORfJ2ylxCTRbzujhwpT5
JEDxkVL0IYA77ohmGiQHJwWhXnYAeVLGCvaok0v2Ss5Sc8xzeJ762c4akahb+opM
XMiKXcgAyaTKEDQww0i5LoiR0xApCp8+44W0oIw9s2kdXJPU2Lr+wuYZcYBg3uNu
qdY9EqtGFZ3VHyV3WCq2iLHXFYkv7tzt6MI7+k5eQ00S4mSwe6jjFF93sJ8IqFsG
Ac2v7baB78xZ6kImV7Jm/pJQFTiNZaOrn1zWCZMJXzYQkFQzyvkHnQFhxb8A/6sH
n056bBV5GlenWYoQ4iIQX5BYoFm/zY272S3F3TVMp4Rm8uOhnqq+EVP7wnQEOblY
HCpvJKwXMgHgQsJ35J1eJ7kefyBooIhGMDH8Qk31qD31HxcplbGQASk9TlWyt6Wj
2pKrvSWqA/qVNkweyUtyy3CLae1a2Og7RhT5pgovqYGklwAEC7hStyGO9yT0Sb8H
MRlflwb1wS+9X/HJasPCqFQQE2dJ675BFh32KJZCYl4VbJpgdWwugpNuCUQA5U69
BF9IqxBxPzvnP2KReTR0p4Rc6Fms+eiEnDeJB9XleLYbAUWivUzFCkOIc1eQab5O
fqUD7RDom3tClPC5Gk5Wag7GuGz+D9a2qp3Arb9ctzMfw1gT84hTvE9eu7F0Ot1k
xaXVckEf2eeqfeAidp75Cljv81ANPhrsGhyFVRV2akj432Yf91ZMtiIBx+qndDpn
tvauvqM9iS0fB/3AS3V14dKBzikRucv3iH3AIT8nS7EcwnbtRLt4dRLdhqld0BkQ
DPxKjpEZn3EmFUjfcnYpgLg8sNzJVWkduIeq4KMXpHHVqMb3lbBW/tDkDGPUknhp
N0E7PGMaqKC3XeqUikFSAwSB1GsADXgtlwyx95+3va7LBQyWtQqfDNfezOSvEJNr
I4ZlEFUPinoIzn7lvPzy8pQb3EldbmBObpsw8dBZvfi0f2Qx9c46dGXFq/Ay/k51
3HnYvAh2fvogNhZNTh0cUJ7i9ibAxe4m0T1oP4VI+KpBUnGT7qSJ2dgkf0KXrkoJ
uY2OcjVqjNh60355dPvTPlg1l2usRJ6WmGD/nZiJ3RKBurW3Gug3XhoD1fLiarlZ
JSKGGsmkqlfYvaTbXHW/RAAFgjx8HXJVpPRlL/AttaH87x4R7OT/V4qOg8x4SKhr
sA10cO6hE8yStSKXWhDVy40PkKGNzod6BrOFl8HoP0PMIo761L44796MV1JfkUW7
yyeYkeMSSz0Sx3ytX/gnC39d0aotfK3gQ4KpUhITWrN5e1jtstcoC7U4oj2EPU2M
CA3+1sFdLCUzEY4LtDA9TgP7RGy9BesiPWGP7+KvhR/O30Oy0Js/T4snl1Nl0QiE
3K9dCy2VFd1Vv2C4bfc2m3T9VtNnYkT5WGL1mfAMvPgejdzG5OvHiV4XBFjKCRlY
Tjn6OJKkC2KTYavqpgZoLR7k5ZnTXyhtcVjpnJNUi9AazagT3vOhvrzxPra/7Xlo
xyovAYv7JO+JDmCjFUwcws92/N7XMyq9pddZG6cU/hSm7PcM1apTWm0b2L1+LWXp
X2xH2nREZtk5yUKgm2/nDmB9odCwcKUGAoQIiCDoW0v9G21rKJhL2zjqGXkakIAC
2Wg8HCNaYQ5PXBDpRx2HDNfQyW8bJWJ1HLf9UplQZvrq+MgEkn5VSRqUQ7Itng3S
iXG2urgFiLz3rnF5idBlYHBMwiR/+qhEq7xH12ujIh5SqNfAs6ZOEQQvWjUXD1wX
C4p2aSibofrED0fF5face7UxCLjBK8djZMAf+Xo7dgF/QrggY0GBS6D5XNE12G4p
ZnI6/8Az054VMlqeifkGf66y4g3LSceMft/RYQeFNYrk3KRMZYdRXixpKFnm19e+
wrj/606FsJAdlICJPT/1kWFRCPpkFz8fPCiQrDEhBbzV1/A6npbrtB3uSiWWADan
0agphbPY7fjl04KXqD4W/YrV01sIeb8rxsTdKfkA1RHx25tcTb3u4+9qqXjZMUbw
ijmffcm5x+Fr84xf/OcuFYK9ezEvMO12usZXcIL74R1eAoFXAexGTHPnxDBVNdsX
WrVp/8gc37pOKV/6oZ82wipbjaphiFYrjDyY820281ULC0OYKsFSg/nXKt2Srie0
1d/eARl6paEnSvlNiQZ0XGLdVRDbbKjv3ULBK8NEAMdw3DutOtzWnlVE53nn8w7V
0Bn64s5Z0Oui8C3xTf0BXoyysy7tNu2/pjwQ4BUEN95uvxeLL0jccxw9U+vWZzcY
UnfhVvt6iUu+tMzLzmEN5oo85uCpaAAuCeaFrqIuS7122YKbaSjUZLz19zyVw9Ns
KMJ09hLpBXKkLUrTPxfmL74L++hr8X5H3PJ3zas/yRfPkKqTqYbP6sXgCt7KWP2o
BvIXUzShG9Isti2tposel7OTHEIgJ6riZMqFrR+GqkaZexp3oCYd4PogUKhBV9Hs
FFJiOMAi3+NW9ixuMTu6CEpxCMwx8JQir/83E/0B94PWoF9CmcVhZjKIWKarGVWq
Ed7r5YKrzKMFsvMWo5y6EJKf9d0dqR5Nwy8Xx7saDW93sTuPKUw3FtnW3PE1vRCE
8NB+c+odJeAYZNidt4JD4QPot6RVVj9+FwhGA1sDJ2rLO8w7QsWO6aHpOAN56rMz
pyVRxDnUsggFoYguz6A9tVq06/g3RoeLQNWD2oqKaYHfsTaiHW7kkO02TYPqsO8d
73kwnfG3Hv2S4Q0Fx0oHoyQvosYonkmJp7yqETEOL3MeWHrxpOr01z2Q9OAyOpdk
KcN+B3VcRmMG91QL+1AD7Si/J0IUaSHDFKdZ0HYqgauxHb5g/6VqBKlfyzHhDZv6
72pWVPKNaIpFV0HoM3iib8o6OGSnFuP4RVuXSazU3tXD6myZKKenqhtYbf8wau2A
wzPcY/WakVa4vKZKL9Zhr1Btc2iDJtLAL7aN9LFY7FCsJ+3IAkXaqZuWBF8kuSQ0
f6jh53TYGJ4KxRE8V80jcCQVYjf4M+10Ly+hkSLAtKztHNQK2lLeN9DcMLVIwcp+
LhWcARPKqnn6GoRQpp4H492gBu3rFp8mD69ZVDpPLxapJhMd8flbsbxfKnzkAx2T
iB9R1CQyzLONScXEVwVD5R9by0NLJzMv4C30/hTS6VKBZ8CiNSic7fmXdveL6Rkn
tHcPzlfBfpS5bfNAXJ8Md99WyC1a0tUmfyt7IgA3CbNXrN0IJLLl8DOTssXqIT6L
VBAxr8qbVd5qFg2/+aHcAg7DryP7VnrLEJZ99G5/NYNDegoze+tGyrUiKb9oZylp
pDRODxJlxfzw6+s4SAmryEwuYmLfCio6XahYhQBMz5XKB4mDdPYLbGPEIV6fN9WN
BDo/qG0TwLqccYZJbraHvhAoopenbGFkOrkiw7X2ciny3jW4pindzirFXhR8XG3X
APi96tIMvkjNAQ/eLnyGXlp8Sz2+ZZsOcC9HR7LFpXq1rzkWI2DM3f0y2o6M1A9j
hS5KwTjRhRSvdbJwdn/Epab8iD+5G0A01mpf5DxqEu0eHO4IsZ9ws+Vaf1kfYKEt
Kh9gFpufuMd/dmuQAFlryeFdc1Vq6BdzCXi4r42xMLb1MoBZZPrBfo/vjMPJpd3A
quVXEcGkiiceKM+35ritAKCY4Zuglw0a5oPdxIw0pkoyikCgZVIN19VcZ0tDaNDi
jzZOk2OePF731SCLIzJvRSn14Gadmd2Vr303LmWPxMSUxQNI3JC9sB+J4b6pK6+3
BYOHHlOmN2rovUfLeZ8hdgdzrBi2HUYvWb17PuvGM5s9W8YYjcR+ltha5QXq7OZS
mBLv16N+Tikt2UUN8s7tjbr0foH3Q8bW4Xxgs2+RpqpKys+A6WDTkoovtJ/gm/YF
1GHTaEK5jRarKFnx0TYmUfhO6YT30IYkza7c1uJrxPjOgFrWIMFVkcSlQP1fdVFR
Zh0T75dzrLM504E+QgmsSYO5HprYQpxL4wBnVcYavKoWA/2sXNB/SK+yLODqcIex
MJIcROQ/fHTXEAKc6CCad6zHQGENGuxJzac67U1FxL8HLEpHh6bi+j6LaMdGSlXT
2ccPuuXg0DYCbO5jb0GeG5MTCO3PzgS/E2BbK0nE4DsgFLHD6egEU4yR4LXLkvpZ
wc2wlxIvqfLh7+IVBZEANxHDS0aU3yiUF22EgLQcOgLzA1N4MQb1EqVYVG0E5+G9
8hGoEkCtjsyLt07saBs2eMbVUPNNd/LvtQOBEW5hCixqpBjLrJko51zgXvsZWvhT
1mo+D1etALoex4GyKepTLxJ6pe7xOHmgz2mBdsYL9IpUnmoWGgvSJDtrEW66DW3L
lbqbweW02B60zlQAdR+GFQ6+7VJMepth8P0LYWjJQ3pe3XjI6/Vz9K3T3XaqMgh5
JhTFDpqJAuK/VWQuQzmUr8OMdIYFP67A5JBnK6oYgHHmRd6l96m4tbQvWiwQiOCf
68Dted6CvFHlkva/KRUyb4jKqNQ8sjzEDSu/W8NTJVtVl1COQbBfPwWDAC4OIE9g
1MsBS1Ne/qB67GWydXCMx0LgNY3n5nJ3O18EOr7u5yyhx2jTNkHEfowdSLZMJtg9
oZtWH+in6ljsJukNd7v4JC2b2HdKtkBiwOB3UdVuim52X1+sqZGb+sQJounvRf0c
3NOHKvz2eVNzSRNmHeZcw+6IkcTE88VXY3fOrTtFFng/1Iy1wkvtFkKnjQ/0NaO/
LYHJTZZSgAZ6YT3CC7QJ7lcyHagSj9pyQX+u2xY5S1dNg2yLtJVfsgrPQeGd8PAD
++HnXLxrHrbw4LCq8lQKNyaJ/cxpIj+vKYt5jY+txB8zwpZLHvs+Mvabd5HMPmf1
xE7kvpJ+Rak7XiDPRMeYJ9ZufYLaNCZPIGozybtc/kgtQ3cfmyqP8wgeCoe4Ixak
hvOIqeWHofDYZtmbvfxlYBiSyLlz6yWxARc5eUugBzAfh7edsw0aldUQfhU51kBt
cw0Bjt42p5KNLvtKbmso0SO5FkPATNu3igpwP4KTP6FruefbCcW2VlBLrZEXr/BB
YvgXyJfi9i1MAAXjFgxScXYLvsykd0LTokSpa11abyinvYn8LcZeDluGbdfAF9Ky
FrgJBHXLFpp0gphcd4wAi4pNhKErosRSRe7J/D6kvGNrNbhp+vCqF7WoswI1hEoJ
3zUvW/QERbZDfz/9CxF7PL936SqicNvZ41nNWxn1Njw/cogKNYyw+/SHRoZCaPy8
Djg+9POuLTxlPWRTdWuj9PbvsR9WewdDN6DCm2XkSq8cjjW56jwWiDc6vurLnHy+
rSmMslpFHwag66zuZ8mM54StBu5lWbdPhViiKRdGKCRDgHfAFeSN+sPmQWm70ZQo
pi3xMaoLIHEYQQoQebiprNCV5YQIHVwkXX0uq89NVsc=
`pragma protect end_protected
