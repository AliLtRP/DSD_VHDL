// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hd1bqY2LJdVZlKD/CUMHDrHyI5R+CDgXzNQ/Fmab4eQWTivIZoKU7KlhthszxZ7b
rdEZed81HhgrqtVzKhYpd7Y0bemO6jKHgr1gytcFbiwvLZsFX+wTgew4GAagy7SB
DbChfxY0ExUvEVddSuDs73LVeQdTClBNdB465IOfwIM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19632)
/igW80p4ksybZoUu4DqhcuLyO88Lq/3CwM0VWkS9TFNjhdADygzzRnRrawBqOQaG
wEUv8znI2REsb8qKIXjLXwCnG6y0PzNnXaImzoAJZRV8XW82BuYrJfpiiJPppPnH
1F4Ue30btPgNEztCIj1maGN4J/EZ3SVhJbO3BDmbJ/WwwVenTLYPO8b2inL/Is2i
LdJqt3rL9tMgEkgIvWndWGHHcqdLkXJUz+KE8rA631etEamuaDuynSOSnY2tbQHc
3G79pC87okreQgCqHSS9zElMEgI6IQsKR6PMf2N07SGevsb0ntt1Ji0LjVI26ysd
WiGCpz7YHe2r0fn2524dq3yjHrdMaIOXB4MkknVzxL3yy8UjF3RiX9OL+Eph2TJ+
eJP/VE/SZZFQU6chsckuOCM/m8NRLrEJOQj9L96Q69SW/0Kdkx+G4UB2DxPnPRsw
JfSTuvhkq7F9o/1aTwL7JQMff2LsWM5Mhu85z1Au9tyFw1uIXspd9rkbLgF4WfO0
ZkqP64IFkWT+wfCoEIWgF9lMrQyxEBlTy+FU8pItAFPV7WO9ryUL5xPw88b5MJb2
n/SqhmO4NHlrJxPN0hhemGaJG4x+RlOzqB1t/36P1gzTf97mYmshnHnTQYJ5XbOl
hrXhvPcyNoMd6zVVRHZJCkdWblLHZdoMxr4v8JVrpuDyBpY/1MMVTQd2BqWo5K2G
LYlnVPv0Zm6R9fZ/0dcJCRWl8ccrOxDOR33ThpzkWp3JmyLNFVCwJwP2T4KaVMoC
5rsz8DGraGBXcb0x15hXMGP+NcusnMJkhuKPC+CJFteWQ6d1F9U+hhPSdeVtZO8A
pLMd4SlIowEuESPRBllVhqodbhqeRra7Z7rUYnVG/nGvRw7qrPwbpsRPJpT56wsW
4ewTE3paxpjwvF9rVXd4+QmvU3W6uOMp5KRhSA9oduzYCZf13p4+QGZ8idjBIAvo
+BLuGqrWmt9mYBfZUXFZrX78HEqC3FKdJ/eRoI99BPngaKzJa9gBeUUerZZHNcS9
X3cCBURjrmx5divd9bdZD6UtUGoUFf9ubs/hDarohpuU1cCiI9KRdJmp+yBdkj9J
AJz98XcdfJNylR2FsGTMugnUAP9d4dDl2WLYz57dUIIbRQtOMCJxclpQlyi+jF9B
q271SSfSYBeV8oeGo9m7oe0dFMJ9QH6KVSUecK1P3Y8MuBIZq0wFCwksyCkHzWB4
yjOAOLUoBw+FWzjlL6qXBN0fP9/zWNPEJ1xY4v5tYc96+MMcrS2BV2fP8uEwJLaW
knHjsnm03194MLnZOAKVxkDZigCBxYaDgFeBNFcNtk/EC73UytX+qDy52l4puo07
Bh2/YrCom/uBzi303DZ7Q++xxiw3nReoXYatZrbz/1ZUoZV0jxB6UpRO/QuVzukr
Y9o8OtQGZRV9PfT7mGTiAGKw0vMuwK24+HaMvgTs+VzbIQe8GkAZSkj2iR1uM6jY
yxClGCnCmXAUs6St9fOXa43RTXVmC5UEodOKUIEELlqoe6rdUjqs9dCqGNR6mHSj
iv1NBfToG5z4KqJykSqGAGpWjcoxG89HuNnd5HmpttE07RbZHkJ11dnWIXIby7yK
NO+jaWN8yKiMx0As0nxLhiC6gqjbmOek9TCJILuFywDF6uPn+FLPpjrqUgpWHXMG
tk3s/TcRtKBTVgxLRTBSvAwCX8F3Cx/ePA9Lo/tY9eJwcKbigWc7AliIN62ebUEv
o/bMoi8T1j89so2iYRx03Q8d8Y4Vs4Mq7PQPpqikqVXEehe8PjHDs3+aWMN4ceu0
EyJUQliJARJLjp0tCsPpXAR/Ibj4lBUdvCaY+aCsTnduKaOvxXxF+kbllVS23h5d
C3doQ4kINd48nQe0BXkxKjd/CsLoqKNCLbo10kUFEx86AWUhW/HkXqrkEE5RC8H/
7iWH62sgvk1AiSXub49DMzvqPFxunVYFv8j6fFbuN3h9W3Siwx3i3CNvmyIuNjN4
hfQw6xe7wJhufE9MaHi3zpuX6Y/93XTI805tsdY7WzmwPO4cGMfTOTalBlmHVKGH
nG2/zZ3YHeVpHsZcAIPmkhBPU8VD03UpXHW0883j+yK6yfTO0BRIxgWaFvERgqyM
AO0yPq+P5HD/Jd9ibpyFd82OBOU2cR4dIv+JsmTJU6EMr3B68AI3TrbWIDT1FSZQ
rAurg3yL5J/yhjt7IQNmgRMxcQLp1u7NfDneAxgrxm2I+PTzSTKz/jAOJ2IJx0y6
L0TcjttpLROHrpyajaT6wpv/dAwjB11QGD+WM93GWdHvKD6ROCApsEQIRMDBjnmO
lal8zAcIxrtmD1hcTnEgFkSvAqH7MhLSWzeYJ8HyB/nohtzTFRdivVi4FjIfQ7Dd
R4g3/g/xp11IRvwcGaC8J28/AqsOPx9u5gW2qfzOsZ7KP5gfGGDDW3lDpK7mcTuz
wZYBlzTAtEVr+/Zu8a8UMHnwibg2xQz0/+sG1qinz9hnLq+BM415J9tn73G+csFP
Fh//6ySuviZHEyPNtPxTt3YreX6fRilFEkBPv/IClXfViWb2iQypcdsEV3aZb9hj
3LbPtn0dIzEpiAJPJ0ctCiDdtpPci65VsvuTXjkUcjWy5SS6zXSHyqnFHcn6S4VX
YtVOs1TGGy7YJbq1WKCZFPaeZM5FYI0LfCr0WSKn/NiJzLkMye0bV4tJ2fCtMKOs
bSbgx6ibr6yTEfDn69VV1byJAa7S2d78BB8oEgvHWAdrdkDZL+MoY7J4syR658CR
X0mzdbZPOjy4hsn4zCp3BiHcdeW1LK2qEPLum6gP8yL9zbwrvUePKdsEozhAlXBW
SBkv7pmzyZOkDR2b+ygfJ5QvVd+GWHhCSMGDaWyqXRNKOebUgVP1z1zxfS5uPUSb
xgWyKVwxjEyj1M78WS6JPWpvc2VvRN7t374FLtaFXKqE1oZcHg1RbDV1gUbfgIHc
giffUEOSF/OB1a0clp16SKyDPdXk5x9K3uTgQfF/OQFGWm2wp81gr33jAnn7jPdB
Io6BjGxjf03nmn78UHGG/TXhlsXtUOikHb1sqwqAr6qT129FwYsJoiJ46qmNmRGN
b6RK0gii7Gpg93iMJmz+ijleBQBa9aLOLR4CZf8AE0Z5VzpNVR9wPx2jkGDBb0Mt
20u8STQcCM0NoUpfbARyNbdpn8WY/FwFzbHgNsGx8LRExpJWpulhlnX5feok852J
2HnG8QIsTqfr0/BK4g+p013pueUVfAM42A2r5oDPwoDSwU5PRjgY3S1CyHPlLjsX
TzzHZtYqzZ/5arl2dtPhSqzDuNqa+Z3gGYTugOL0hr2/5n7FIJzP+D3bWLvbZ7qW
MetZxc5EOH+j9pvCi//e3eHoRYa8vE4fB7m6BghgM4hm0QNm9ZB7v9dR7g3iBX6U
UY8cgpBXc/RFfXGUdrMtKCi5gCIewgokAymyV2akRvfOtNbUFDyAxqQKCEAdAE0i
JTWajmO3eqrMmmV/lCkhy5lHWByTlpKDyEXspuF1BBmuHQ/S5uVU/3lHmHJjk1rk
khZWshmrV5/SJ45wiKddvb2uIHiyWns3X8vH0cpCBRT+FKo91Bt3HFM+nzdhEWnc
YKZSGgErVIYSHLm4axYpRlrSEVSaANiPCmqcdUnDpHPx0+F+ns2yvtbYuhtuS24n
ldTij37tZ5DyiK7A7K8YQstOkDQMzrjczEuG1SMVSZp5tZZy5Rfwu27AxiHyOcbG
Dqw3CuCoXx5TeY5D76YVlqSMwKN/ntMOCikctsamZLB+uOJjPB+69osGBCfA4y2c
9jTsYupYzjUXJ8+uV23IRx9E6rj7gMQ5pzkJpoRTqchTgumExiPcrzSNhKn+OiqA
bmYj0Jc1QTed+ero3iyDsD/Nd7dH6PBpsTikfAX4lOQGy6qeLDODJ/BRxgQes+08
wIWtBRXazFQUzERHDnE7ItiHbefCidQLU7NBti2XQYBsukCzDC1ar+zgiLiVKcLL
LniXmvlxMA2TsGCyuPQ6WB2Ihxoash7zb4oQ0xBV3lhfdm+Nc6rxXMVw+YUu27dt
7QGVG6kXir/JKFKRWhUmJbbrXdxHLR2H5XdqNzjx78swB4N305e3OC2PikoNX/yI
txmauOyLh+c5BzLZBAxBq//3h54nbiiNKQDeM80Ki516tU4nN8ucODVT2b1HMedj
e7V/3W5gzPVrNpskEH9y5on24XNXq2mkp7Zbmk9l9CidWroo5R3BMWpNFn2E0qri
XuSMisUCt4UcX5AuW1PSOERjhjb1tmHGtb7WN1Wfp04JueQeJ+0IIUlpIoYH7hft
0wan+GxRa/txenCXj/JlG7o97wrnthoR9kLYHXB0J4MwzajY7xCrJ51RnrxwkbPA
l3ym7dIC3FkBuWjPCHApfRvZGrSjGfng2yYiF6DqROxT4U1Am0FUzXfFksqK9BlX
Q8NzWuoHpTA8D6S3XN1mCDA5lJ3bmSW9IjDbrm2guONNvx9gP+na6Y5q/H3U5qtp
qzWhvoLMU1pJTL65ZlcuuE/OXX6HKl+bEEYV1oJW3yibhF4Rl6p6Q2nm5T5o/oNC
2kLSmPfTuf/wX9fyFOSc9Hp7MEo31neGQnmeU2r+OkgaGFn/bEuzPcMXMWX/kNNT
CICw+BqfTNh7dPP9sQ2aUBW57OKgqo2vs+Lw5Emhv6itHa8F9I61OZErptn3d5zC
x6jSf0hOP8Uvgyj2EqDegsCYlvy1H+x8+Z0aZpxZRnsJn0GBQdAvzQ9h8bu+/t3a
7IuxEcpjQCP2AQZeke6uKkaO4o+pzOXDqKKckzp48T+lbiOoi9tacMO+Yi+Wlv2d
NWECHch1l76jxfihSXC7d3T3mEJ/Yu9h2+ejtrU6XFNskbXT3EQQ4RHk9rxJ3GJ4
t43Wg8OQ+fczdThl/LDaIuWOVkMj1kez/86X8mgXfeEBL0Qmff03NfdTpEQLBNMI
g/HUTavVJrrZp0n5RpwQxwvPYTdFWG7ZwSKZJj7T3PjbN1M4iBlKht5c5sQsHk/Q
NUMs9hK2VS+1BXNQnI8RilDZYTE7FHgjAC19KyQ3Qcuv48KetNi56aD1Ac7l8HGC
3ou1n/UAtVzGKZ6+gvkoudl1ihmgKupfNx69N2pCq1X7Gi7puOGab/Kje0pZvvg/
A/eWr7+/NL/eI3/ZOx1pri+HBk9uFgjitzeUpY8aDrs+uUBdZBGDBi3VTyQrMA/V
g8NRE+ey1OTwHWKwcXpST0ls7EqMlIyOLo3IIA2ukWSrl/klfdnaHEEvfjWbweS6
MZ8V6JNF+N1NGAsAPdRB6JJRx9UU5vAI3p92IVIbWWV2U4lbP80RRuFrsyel4eV3
NKKG5L9In+Iz/v0TZHQOCajVfYTFr+J7TTD6Z0E/DotilO/dGbrWE9IZw13UyokC
qT/zmw2OJIX5355ZGf4DqhVlf6kp2I1OLuIBvIBTGQSIhgcPazecYw18iYLwQfBv
dEMdhwIqXVTQS7dDb/tXaUAkogAvPFNp2E3UIF2SCKu6C+noZPeCm3HunYWeLsge
Vyddw/1Yh2iLD9C0t88bazuULOJ0ugN7WTzmmqFxyovXKZ1Fr7Clo02a9FVEmNZn
unuKIdawa96T260xLQuWhGOkMKiBl4jDAHa6kJwKnQQlRK/djv0AkHppi4Ha6UMA
Y0cwGKyXg/f6hT1lzyHjPDjBosFiOskauPEEMvNzousEfTFLhafgnWFL9yPOWGm3
gUVUJHfkKXn3FFjUGz8CWf+qt8+gQx/gPmmXIC9DLuTBXSxXtKh59S2mGbkgyD8i
UNYT87rJhTTUbgZrO6/Nq0EEsfm7+hEKlw0/0eIiL2lh6q1PxoYPRLNZs7CrvxSh
o9KnIvKvZc4hTcrpYzFvXOODXQRrG/r8B8RY6n9VFwcams0NYbUi4F3lc1tENgAE
z439XmBC+qWEmhbgs1HpLsf3C3NkRe7JJqK7Xddfn9EDO3f+eBF6klZXXCSdvOx9
YQrj45S6UDYCCbFxSolpnESUxD5X3aHqWRwwyOMSyOUDiQ0gq81ZCGnCWWtxkq5C
cPhNr/2x3fbOMD2+SyD9wQwCd6I8eAbFenxDQlMnI/94dMD5u8RpiDevGiVbTsAM
cHmzFWaqnd1mqZlu6ZTuBtujGuj2zTF4nAGpl+UKmQpX7Ln7p63cD9KWFhvS7fRx
VBfuAge/Vvd3/8IHV6jhz1ERULm4RHwo+ZObJONFcB3xgWvmRn0TCDCL3xs15cJg
J8uqQJ+BtyhWyEgqxWnuqTJGvc/gOX6Ww3UQ0NFVT6u49z0IJrD3jz6R7LVx2MK4
Sz3h7iFAuuK1rsR4ZF2GQJ10XGnBzu3nQk99qA5xONLmX30mOjeoPqe9tsQkYAQ3
mb41+bhEA2cqrjfCgSB/YdRFwWrSXhKTjwopajm1995UzLmhQ0S2CIZY5TZMrMh4
oZjof6gc/jOTiuTPipKgtcr1rbOTVl65mJQtaLGVASGQEIK9cXZUZSnstaKgvI+1
UobDG4Oyv3H7TfGoA/cIfu9jIRusSTOAeYarMJNdFIybDtlrqX3kK6++/B4WUTrE
08v1/A+yPBwBcd6tPow/f8m8NRxPxzFscKjeuyUOMHW9djio6O7bFSgFD16VWfYo
zco3X48dQBO5rC3JuvwZal/FDABJJGRHvf+kS53s4nCe79iQHdFo7H/da5fr3RLC
osUNBi4DKOrlBhf3XALwX15zH+rNq8a+/YZf6kYELWCDbvUHcEcCKJJX6YLEl9eu
im7YnX4U51lU8PGn1EBJMj0xKgVbMMT6a7lnmAsJ1ZH2+1qQaE7KMAiAR6IsANQX
dBmeCA1BgyvlQpnnkkRTfM9Wh6I4HaUhMYRNZiaztcjiqwVVeynCbP2e1uIDsIQ/
piUrm5soOj/HdFxq2aLzWvxU/A4uJ7uC845qBpyCS3QVXFs/KQIppqXRAKE4wcUK
6L5fIZaSLDNN8ZrApe9FSMcbUeSZiAW5h+D3xs3tIt4BrhXp6BSD3EuBDQvt8RZZ
0hUCdoVOiJABObuLCcebMOe/jUtRT9+0EXxnUJritllLjI+uxbNPWQt2ku3vFgIu
CJRHuaDdleAGo894y/6TpcPLm+ICcWwzV4fwm+KsVh5UsdOlkb+4fQN+JiUkY6K+
V6TpCF8VEvMtq4DFSzfzUyA6Nj/mCx0QMLlReQxuBXHYVDwVQTPKtSLU+e35PSQc
jF/maZOeKmFqG1w9QmwiwYDk4sWIMfM8YyWjo2lhboD2ZxjWN5XsIJ0vsjWjC/dO
/Yd7MPM7DBUR0GA6sdgF2/PYQ3JUaXkT3Og6gAmaSMEpqNlf+z1HOR6caQa75jdm
z71LoDdsgOcIFcznHacGwIgyeWrGor6lpDdTSjOX3LqFajuCle0GsfggZ8DpwFXS
6Gbjj8r4AyoaTyYFiHOMM1ptt0ck/cxp1KaLfK89fuIaWX6s6aZYIpE62ngiuC22
ysmcsdJvIYXBNfmCmfRaOe6KewHoIoqAJLfbKfyJAc8uyTdSxcMbHIZIB/WKiy3g
ynqMIVAxnT62A608Lzyk+FVADdGmBh++Dxin839B1jtx1yWBhZzSoiWY1tUNEKrF
an8dQuGYxTF4lxgjFz11wc3x9cipEK0u20ZEyvayh9Kl5wpXnIdVlsn2EBVjnD7M
xMhvhDA3bcOCgnBrg3wpm5lBUIajC4w9azIxzUGm0WXnDOuMT2qkP2+9udLQH9Sx
yC/tLsahBjpu3yoFS70aMv1vua+BM6fte24aS2HEifmRhSkIrWBQDLDAX4q5ldMf
JblhGhE0T3OphZ9ez6IoBy6hWYUp7j1CO4OZDFDJDB82LXpfq8m1EAlxPhx1Vig3
5iuTKCE+HETNYF1S15WvAggLttrAS3ZxW/ONUJt2uwhbHpTUZO/IEzIa6BHgoCBY
YscZCfVtsNksDnyK2y5bDaxKIbQQZUMKqHP6vON+bqvPrmydrbaz32ql3XwwvDUv
R7ip5X1ADNPqaG68/ePcoaLXtNo6540shTSmfccVkS4YXzL970RpSKPSfmb1YkAX
umqbp8DvpICToQGJUtOCGgEa1Ad3oxl1e4ilDcQyAkD6Ijdk8K9h2X2fZG1URIuk
7VBD+7USQIERJj91vXIlU0uq/QqSNidg+DPGN5XzFjU0qnh/AZTUIeY39Ufz9/EE
QKHyD+jMdvhUlsmT8FOTF0ISi88rgZse7rJVsKungQ6kiimAKPOnxl5k+9tRshaH
QLyHHu9d9pZnbkqXg3tussuWtYRmztoTQaooi+8q+cwN1+ta+YvfF9IFLMRylo18
/MaDsLJ9bhcIlVOEvgHpLn3s4njKXpZSs77SEzWXj2y1XE+Wg2Yln8OmcZOWdDB6
LcDbgYgyoJU5pE7bIhyFxq9va3hFGPVmL7ku/KX/SM0dwiIBZtC8ETAK4rXsV6n4
r7cg35sLipxuPAmARTHPnbno/KvkcNKTEpd4Jq+t73emIrygUhDAaYn9Te772SFN
t/F7LHZIjoH3043Y0fouxnJ30J6bA7+nJ8OI2ux6UZ04PgKwljLA7qMAl1z8SS9Z
jB6GMAf/TV5BlUi/TQLcQcfYo67X4cEdgowvSNkjIwSx6HptiwmTczf3lVqHk+EU
Gp0soJ8xLAK1QfeN0G1B4FL5D9HzVRf5gvmN2Yqy7zYHJ/EFSRhshIO0zfFRVuqV
8pqZ7dCpOcwlIbOwd/l205cRbPU9ZwCjQS6IwXw1fxe96GAXp8ZJqrAuDepu8e7l
k0NBWvyVfhh0oGG9VksM68+yIHigJZeCYA9dUnQCWMNkbswXNjJNu8VwXOq5ixMx
VLn9qQtDEeiB60rVviAG3KAnt8oQr/lMUBGFuDuNz2s4aXOXmWANDVnhHNVNq2q3
zy88BwgHxS83n+iNMd6QqvRTjB3HXUt1fR8Ez1ylTk/BghfoxVdVujsN0sbBgrS0
vhxGwQHwPuGVW9fQErje+XjuiQm/UCT1KPiP9+O4caFj/xaXFsqEuevmZ1Q10HgK
dO40Cs/jttd1X/Ogg52XIDo+HmFiue70Rq/MmDTypBdM1qhVWCnesTi2+eLjXk4G
qAmga6iQfB/JYRi/mMADo8NVKbhkP0Wn/4GE/oLGB4htuegSl2bADH04W+KT3UdR
t4n0puQY6Lx5uLY9BraqjSlkvVt8qppckKnJnMHGfkK9BWXGuKrDX3m/vd6eXmRy
687RT5X6AdLOA3DLZqPP+lnSp1rvwVIZ2fhErG3Ycbj4jTTYvFeVAvhhqKYSA5Jz
Uk/1DOss8R366+OFSYuPDTds3jbxz/aISZQ7hj9rCYADQJV1IwKOGuHCcDqDuCwq
ajFm5yPfngomJx2TPmBoqm54MHyBddY3CC+TA7MUsA35dr4adjOnfvPikoPKgqBT
p6Rnsf2yp81TmIzPkzN3/clmwS6cUSysOWBwcugDlVvmxPnU7ThH2VQhV+iktIsm
A/qHaQMKL0r9ZoztYpJVhmlssaMaiznEvHzN9B6VoQ3+D4Nr09Hm669S6M69Tki9
ngf0SuFnbFeqmjHPRl5zNrOnZe+rq+hf+tlCzJk2dwBC5QNbP87ffCC7C+lV/evm
3gML5gytCrfaHbMfSPsztm8U9i7MS0eZdtH2tuql4I5iol1i5oKTMoXDDtXKV4qA
Flmhc2R7IfjpuLuoW+YOtOULFaX0OVroVmvLOiGAAn1MwP3xYPz2fC8CBM59d3gg
x79J27XSOco+NWUB3z5csGBGpPDpyyiWJfQoCBcVn0F7t7yXuNeJvT5q+kL5JC0q
Fm7fJ3sxOfj1B5HO2WRI3NVd2JTErPjdaTZTuY8HyKbCA6S/AxvYPIXhOuZmyrQt
Apb8sHZ7mlalaNuNLf0B4QERjCzkJzt7bFVVlkz5/Yap6xephu3IBGsd7zbQL7EE
42ODl1ypWUSncW2agcrT58S9NJrowe91GUDSgH6zW5QxFejsf1KiMELx6LZBQ666
+oJKszdUONo74pMS6YnF5o78tELTx5m8aWp5R3eNuTF0kd+40HmDvUWUEXoyWOmR
5KZzOh17Mt1zBNoosLKeJ6tbVIcK4V+px56bJjSAFQvbedLSWc1ZpGsDtSO34Q6M
P9vbqXiRXVMN3Zi9vw300+tCMbiOj7HponQfWZuyLxCeGqavgs1BPCm9iPXnUx7F
Ugx4CWwf7ZEfhAg+3z5TjFSb+/WTHt41YJ5FmCPKmlix1cJE98Dur242jSl9icNH
xvW0omhNnsfNK4oJzc3MIW0zywrR5NIJ+ViBwx7qagzXQ/STrKwU6UmURT13Bjw5
gTbI5SU3njc6O1UjxkzY9Yo0wHYS550EQjqouLbZs3M2/E+C76eMfh5n/hwaCibn
ziP+6h1/CKc7aXSH4cv8cyzHZb4ko/s/OU4POGMLc1z3WUVVSnpxAcyPKpGh0ZEm
B0uX4G7AhZjxZt1bgqwHr7pA6s09D83mCgIa1id2CkvdkTsGJQZ2xxlSHmgksSh2
SAqpnlan9002gZYOkBKvISi5H9mlxEzcWMS01S8bhTovFPaTQSDmbKlFo2VftWLH
2gj1+QSrlhiDjULl+wOOHCHbW3i7/JEaBxZuQ/gyW4Jy6ifZo0XC/+xXX3TOe4jV
caxTm1/m8HjdR+wxnU3NFeHXdYptB3od8fEWG53oLS5jjD74NxOonZK2sVNCwxJw
gNLFuXAE/J69jUC15RY5ngRI/0JxGlr8mCirOQwklJyp/nlOOn65YDu67eFmVbEs
cGVw4mgjGVPGpW8v6xdl1gWMxVfMMdtb4RmiIYp2xfYeDoYRrs+s/qDI5OisvfCp
q+GZ7GiDP0rc9VtDcs3kiSyF8K4edUWkpjPMe2h2cxksDtqKMEmSJmg7/6ehQklO
w2HfuDdfbfMwCr1VQyaWhbP9qxCc3nabuYsZSBAmPab6hl8ksv2ZiTgYTdaykU2J
945s8ISwF0Rl8yPhFv56fuBJvzRrr9eN9QQKwZJjXZqyaiegnqZFL4ANfMxFSYVU
aqXn6CIH4wLrYeofKjaxX8oJC5ZsZIaHJnd2rH24uEHCtzyI5DTr57vfD1nf/66I
EyO+92pTZQQINGweLHNTZAWHkIEXb2BbWTsD5bU49cWoT++fS55Q03ujb59AjRwW
bsB/6cij+V3PJT1zCrXGUwXKAhPW5t8G+kkM54Io0a31aZQiykdQTqkuQyPPNmVU
sAgj97Yph54b2Gq080zvibViwuxYiAKb/c1VPZgGfwZhxN9o1lKkFut+sEVBj2PL
foan1KvTOli+qQ+WJZ8lJGd5WIDVH5G0faSI14O4knRHDjFXm71nx+ZcgwDkNL8Y
3MCmW979Wv2z59thR4o5RlRbXs3A8L2G/NsRskEpfix5glNmmru3a6p9iNQRCx1b
Q9aHHvq755kIQrlWSiZlVeTuz7OWGCrfvaP9p1JzT5bS4d2Oim6V6vhA/rSkhUtm
8QvlppGNGvRDJ2IXnDdWOy43+IlBByfmQ8xeLq0LJNBt8YqFat7LcfOiVd7Jbprf
mGS2n5J4KAFIaXWp+KHam3VCsQBEe2RvnDJnL0zT1wPLKpbmZ/o9+drXSv99KJlH
WSHZRidWY6RgTxu6PmA1D5nSYCAYE7uxpsh3vwFWYvyoCgbS5EEytbtrnaiY3K+o
j6byAKe9Ki4iywYkjFqCvFPOW4nFrHkFqlIIAbrIcCnoqW2zqhGQ8HLyVIrPAkeD
Z06s+DqMYPwP6LvAh4YVaYiYyJAYPpIAuuqlJnSKhbpKtpcCU8M57IB1zmE2vyqL
e32MGnc3C9ww1NImKXEh6KpUjLevFhlNTqy7HU/gK/R/GY/5tlAY+PzJV6ioL/4j
GzDe7DWSXGsiotRXDctFlvFPhntovVGev7FQ3TnvlExwDteZP7ogIaQzHjMja7yt
x0n1EfWN/QzsnEK5ld9bAUBqpQ1lN7gnFSZ0Nr0Q58KDrpYCJZ+npVN8EoO3DRxf
SwC5f6FLJl+zceLgvgH2a56S7n4Gx1tHY0IDb6uNJt7yZ22AVt11GxU29pEgc9nW
iOsPqWMOXaG5rLfWkbSdBt+1bXWYlGKxem7gBE0XM4LlAAMmWrTRbWuMpyOi4SiT
PsO2y4PzbcdfaLNS3D7dEzqtJA0h+ZhpgeuuEiclXaWmXZudJ8JNjlDCcCvbFfgg
O0keB/9cGZ6vYzp8BlNmpgy6/Kxw+ooXYWpqplwG6P91mzdLVE1kKCubaH5p4Db8
5dTFVGS5T0gGrVj/0Z+sErheEbp40p93R/sS0DWMEdP2aCIOanL+aG8N+2YYAMCP
xtRJBo+/zahRSkPATSFI/nCEoxICYvHuLO/MPKF8E3QJ2DPWCl2YeAAeqmKrsR7d
p8whUlU8JXiNXS6BWZ0a1K8WPQYkkw7F/RpHkPhmITS8P21+mskARRTWXIXQ04gw
z8bKzgZqirJdW9gFCB2THvGWwECddGYTx2SHk9Rt0MugNB1rPwzf2INY4VlIq025
wnfG/wazRJiFQPYDliiYExF1bxibAnTHPht4RgSNyMSbtCyDr9Erm/7yscjZk7nL
izDB4M2iejNCprRQcBoOSlJl97pnSi575VRKVa0JEeiUzVnVCALZMXzHHiGpHVzG
2E/7uFr4YrL2NujoOcdNQoFLGzIREiY0uD1u4FTaUzKvHrexxyFh/qGSfoYr2k61
MgqmG6VvFispNRl7wy36lkruyDIveL2IFnIpLJ6AIh7kDzUNOzXoIdkrfAJ/MtWW
QjOn8zUCCvgwy1bOL+cQkuOepd5hRPTnT9kxS/y0dBhLyZj5/++IuZU5CkFuFVQ1
0xZIpEDl3lznogVNN84G+u26JjiBXXtvk7W0puhAH89L3MQLV527DI3OGIzfrpFV
uLXL4FIph7it8CwYb2eIakGdEWztkdXsqz+o+e0hUPC85gWUibVKOrEbBBr7hfXu
GJfYHNspNaAiMCkG0Url4urbRvkUm0B/ZhKvnfswbNwrQWEXOhfbeLMM6Ry1Gh8v
VVaICkzx3SL4HGkORjCI2NmbIJJvn/QdKjDjcoDUR3ilhySkajk4JVKjYaQYXcyK
KX8Kp7fmVehGKlSiu3FQtpWmt13OQSEBPbAuiZ2qmfraMe3zlHeDuOREU2WiUoja
GtS10CHIp8yS9si1rQkGnchNe4ZWmU72xvmjyFSkDfHAfzWjFPx0QsVDwLx9OJe3
DXCGyhTHOTWJGj0BihnYg0k9xdGQZCXzkqEvtPxKVzgxEY6v3g+KNcfxtHrTx348
lUeCZ+4Q/1IsEHLMPzCHkB5RLaONSuLr7AUUe1lEgkU44uEqSAyjF9X+Nwe9FZ+S
XAp9SXPPqB//bB0LrXDvHOoT1e1z9noUOm94Kz7Um00JCy/9BqxgQ+OmxZeD5UzW
C7W48ISxXuRNd49QRAF5cpb9QLy5WRmlb2WlEsc6eiKIcHYbO3PfLiB7uk6U09Xx
DI9XqTg1oW41Lef6xgRSlwpFJ0hiHotklB08mhPOUihvIVS3wGSr7xTC93GIy6vo
ZGhjx5eWw+3qTPHdGz5I0uHwdcu/VKci2KoJBowhGQyqT8ivGh7pBFIIdVFqlcFd
7bn86VSFEb0QI7QupKPAY3i31XYSdHGOLJowoGcXXpdQWOf/mPbGdoPuWgAr3eF1
/OHzkPiSz1kCfOFUw8S+Y7GNycHUaAp0TwDzV+l8yf5iOTD5FNkhHbVY1oRnH50M
Qwg7rGfy0tTdMz0NbLmZKYijt8ujohLGLzKVV+NG4pj2frnP5V64mnqIG8v/OCBM
aFnvUG3ZsHXJ/A7RtbwATB80LbGkiZ2/1MvAbAfyeWtAfhZa9hufkclZyRIAPPOF
YMbK+xIvQWyUWeDYlEVLWG6lEntoHM5B0zUGKKiJeVdJDjhCwjEoXNpWjte2nmc0
Cshn71A+IZBaxQDTjbhYPA5/LpO73AxC7hZRcCcMAtOUmO0U0/CxlPlFUQUp84Nl
nAvsm0ievmie2SKmHL3c+Gxejf4u6G2XLXQh/oKlRBLptdurIq0dNxoZUnui0XGL
nsXcJ/FGTZgfJb7YY8SBxgy0FSWFKdsNifnD3x/ZyqgMpqa3AsEvz710Pnf9gY9m
96rE2ucLsSssGjQCWgqxPHTdYH4o5Jx/8cEVPBKPOXrqnQeqgsmqOQLMClMwPp4M
z1yrRmwVaMerQ+RBfnwjPS/mzoaZ2flMuH1NiuldHq1/J/GVCIQZDboDEDpfOm2u
GidlNuDb5aY9s+QJzRTRvDYRxveCNhcnl30pZAmst8SOBwTDOtqpre6onWazEImL
5FiU/vHou210xN5bFXOG/pC+Kc+mevE0Tz25blQT2N9iqL/j8vi/kdmUbYki+tw7
/8i0sRwe/qXQeqz5aBo7jslqUY79UojZjgrdSjZLskphpCqFtVidbdQuTUbA4yNQ
CxtIVndJkkVR38g5JaxrqTeZWJrr8ZgCAdDh1pGf8zqaQOFJQJFMMf5OUXnnK+un
kziZkL8dliemSN2GvC65bjuZ4pE7Qm4+lILn2er4EVuGKhxjTNgoSxCqshZzSMiu
2BWhsZAn1PF+Td4hW9ZxZaPpkJD9LsQCGF78BG7BpbcRS4xZa+3FtPsGeZbeNL7Z
3aBIkEphQsOcgxzxbNYMv0u976VOPF5os2JQsnOEgt36sqK7YPmcE6bjcXHOEyul
3nkxd1E/ZivowE7J9gZusWMs8F8jRaXfbSltQ7nEaY4PcibQ3Hautt1txzqcBWOh
zsl3FnHr42nVuXEoECjRKNiiSuX6t0LL8+IhJj/eh+nUwqxYDGHbs3RMBzEEmAlh
lmJGF7kNoz77uT/J22aFQyVjEwcmFY3TxcFRy/JfT9FA0O2aW7pJEsFoadqprsZk
mtjoD76lvEXDdoaTOj9fAWgUJbffftThO61hOWUhk1ZlicmCV2EyMG+aMoErwoDr
JTTruJ0fCYyX/uyUoP/44yGcKMPnPCLZs7idClx1lQuQfklDYB8D+NsNxQfGvasj
7Z5uTOMCKBV5qwYIdB76xcG6lErKyD+FL6lwzOwOoILjjzlz8uC+tFgHPCMFjJJl
QMrCfecJlGx+11tf5RPw2GuWQ2riS1f89C2PwcxnZVNClPwbmRxY6QuLvzkDaVH8
fPm/c8h+LbaC+3tDkJal1irAzw9kIZug7RoNczfyi9v3lgdru4HpmUZZ90mVGGr5
0lRucN40XYSfzjTP/tbXSYwZ1PF0FRoK+yXsFu2s9anPzcxdD8jGsDFxc5vYHiCx
Y21Ju4gjPKe3C18JB27C0BQLgfdKrRnwP1kGtrrGKtNLTBeGg8okHr9PGIwVQRlv
z7ZNSytZGJ4i8WeguWRFYRnjoy6UtbD4otAsb+Va0h2wgWbXGdpda8z/PwbuTpg8
eVrILNP+4kNpgqGs6MZF6h5Hf6mEHG0smj2zxZxsnUaSTa/FIj+grUHcdmWGBNdW
Tjdy2J8tb4h3fvuX/0K4m9x+PiIzpCIQiWOXAiLQETMRjLh26GG3NxjeBjZVwLGt
TCtwJL/ANfROiVjl9etU0bpOt3C2NDeYICrdjtzz/m7pa7lrdce+a/ocuFuw2wSK
p+deJN7sqnImIpSzqQYpwvW2OlMHdall+R9wj5PcMpiyhTPIzvTZ6ybiQitFz7qq
ec7/jEg9AdGUF4CcV8FgJZ5a5iQ6loaLBSQ7ElpbONUATzHQQ625WjEokHghMYTw
J5kaYWFoiDxVzUYXghlg1zj/4fEFYvJbumGo83xNia6Lqg1Pkc+R2PIe7ptzbQsu
l8GYFwAvbVp5LNnRf05cJnS0rscDURMlE/phVmdr7m65N7ci7JW5U6NQd84FzUfa
2/1qWWHO+JivM3gPCk7jHU7L2M9h0GKm37XXq775d9ohy2B2C6dQEEzn8xuDSFSS
wHmapJJhN7GVVev06gRLBbtghfMiPiacsIE+Yad0xa0+I3d2Jk0ciC+J1ev3q2kL
IQpIYFgNj9m2Zgh+dLcXsTN/nNK0fjM4yweG3eoQJB6fHf3n82yfCPXMt12kZrkg
aX/GlqDTU0biifFzyvehFEr5REfwe9AcBycOXt4OI5wgNtkQzMOvITpXIs78Q978
EV5gfkRJDmlCHkHMufQC5mJM3jwyghGGyZOOxClON8UsDVyUOqLb043NNoV48h21
P3XkkxK8YBqtAsU7bvOYKtbGZGZ5+5JumihkbiT/CwZAjXLqMis5/1c23ljQ+Ler
ijnRnZG16SpmeRoGp7a4qfFbuOXfP+nom4U7I05H7z7A3c1TX0ABCjsRFfBim2S1
+qjr8sp6WQGhwDE29MDK64BBSgTZMyYZH6TgVSL8KFZZx81p4pVqtyok6kVWW4PV
5bLn/1/WgstpiPNFRY815ii6z271dgVV0Bu+KmjaWTDc0ucWisfb9b0kfd0nvyfz
eRMwrehBHzWcY4wIqybDAKnKJwJq95+SbE34TLoXbCloraN9rLu3Kn/ALCRLYnMn
Nq3q1zahtWaGm9p4vRZefGUQWS28GV8lSnlAH0rO3IKRnvlWuQYNnyIjlbxdWc0n
y86O1sq6g2RuYI/EYwCMTWQmzvLKYHUZ3e+l1vwkGajuiOuUZXT+bR8mrtYFdwCt
bs/ist2VtPxBggw+bHa7O1K2moClEWbDtQ9RYayPGBDETJLfpBXHnmDJHjnGkkx0
iBSQ4So2/YCrM7HtYyPhfmXqoNZpCejp7Vl5Ak6R2ghnJ1CpykM8ouYnEKHcCV9j
mSrc94hqgqDhGY+DQu2jyIcJxF8AUw3xJdZcYgXyryeNw0Ov+ns/9nTXC5gke/sw
hNivaooGPOl+90JzU53aPKQnB5n00LwaPiwAOSbHd59sa5HcM0rW54coYD2mVUBC
HSK4J8aD+8v2YDS3NHnW2uSPdZBNPhD1Ypet6fsbW6Uu8NsXyF5Pv2mNxwYBukr6
PgjONyzWe4xFqoxnfIvEw9JmlxhiRphptT5E3D2VC6RDvAhDrJKBjHozoRVpBvTf
WLmOQ96SsTj4XgmWilk4nJl8F4wkkKg4OvpAm9ZfsuTP/6rTmqR5JqfXwd4iLslm
cQ9N/QwBQ89+ICJ5BW8BGRSCzQ1EgrdR1sAhuY/kJIdntSo9oW9fg4af+nb9YuIq
RvM8GGUqN9MQzMq4Ih2sSdW2y89q3YaAvlZKjEDhVQ/nfFl3X11LgwtvpG8uncDD
RXrqYfcgIfL0X2ZqwLinzfKYYSc6BVSH6lpAgcStLkyaC7ddKRV0jDGV4uwByQCI
6bTmZVotiHxn03U+iOIXL7f1S0gPB+3j4XCqhzBCXFl3KUHD9ljrOJLBJgz1EeP6
E7njGSLVrKkEBHv6d3xqiSuVEq2+9P63bDEocYsYhTPeNzJRANGhC4denFrHyunA
foYQoxaVsmRT2++1XcZMq6Zvec9K1RmX1idxizAdk3qPbx8E/ydkzUNMI6iCwxH9
hjpD3cqDVQRUamQt0uTdbRAJ1dwymbQki5FJfLIPClg6CzZxqX2KrahiWq7zfpSo
/w2UDTxx7Zpt1nKPQY76n0Rf8gY1bhcqVyS7AyrPgRazTC+Pjyk+uv4X3RCoq3wp
9oLm+0pGcPwhhEo+ol3d1XThsM0XRfF0vSyGWkvlZ+d3FFL9KKgmGyooJmnHm28M
XIR+bcua5CldyTx6CqWeH8VCRO0U8gUvfadnM20F1X5JCs+KEyIULCRyW4/w9JEw
EgRk6tW/CrQaYIkBwp44qh3Y4TTF+NSSMLUlNeNB6vbBRFJrj+zGevYfl3bfAqea
sf1Kfm50v5W1VJMLrv3VXImpU0BBShFEsV7V7+YupJD9MZPjHaJ45tKUD/G48CNG
CPyo9AXHc+Y5n9E2o226fRxywbCcnp5gNdyIe6fzVscphX1fU2Kl9IKvthF/JoKX
w4kHLnUpX3/gm9hz6SsMaifLU5oD0TiYaZFZMd/itSTHzFNds6KvgcDs+LH61VZK
rFy9dlFAucNBHyjFBI89x18aLy5f6pXT85McNTGw9sw2Oe62HVENkPQ2T4rpd4Jc
9D3pW+xNZz9GNcsvy3pveu38S6gZbY7vyUNBnR6NT1n/2d0mgV5TubGg6XiywzwY
tI9TaRcd0Ml++qBPH8Ii7spbKXNF6cO0vHoDZ77WUmqZxDFF5LdRctXcM9HWNevy
CpzqsGE7vy43ymOMPZtBtF2bbFtee0d/etiUL18vFM9w+1io68EIFta0t2cNx8Ps
EIjAhJsgwjd+9xvonmqEkE8k/R6lembV4Z30KhyqFdNZbTLVb0xDnpFuqatCh90F
rrInmQkVDIGEA/suDPXSbPBPDlnZaqDUzmvOPvYw+bndr9csDUdyZ2fLgpAx7+Rl
ibH5COH57CMYxg4W1pjl89+AUXgq0tdcEJqveaZUNiJDNts9wJNJftm+BGwglGT1
VBOjlnAnEXJf1kAWkfBRLMjByWga7x4kpD3CCBIxAZ2QMdV696ZiiMDgMXyUvtrT
vFAWlxhiuNXoAzU1PP6xbGul3hq5lW+WthMJhoxpRZiPM4P2v6BcuaPeHK1VJdX1
nh6OwuOdSawRkGwZ0irX2OKUZGEnZOVBwdapVEgfAA/oT+WPx+W9BUoiRtDaOky7
SEpRlWIWu+5ikb+xmQdCrrI3mx6W1T2dHCq+mH5kf+G5v1QWFtjDFKrUhxtQgl6S
5Fyr9Q598YXIqY3gx4NwXcru6XOtbz5ZNb/IUp9yYIZ9RtsM2PGbtbOF7TQU2Bpi
UraFIdEs1dhU4+jbFbLZWMO+4fz7aYT5bhMJVvHLroUBzEHVIsJhvQfDonzMx0m0
APO50LJVVTlBzuFCB/898MyiruZcyse1/jeGRAD41syTw08S6zDEaG8uUIdaDE1f
+eghxk55tjksbqvPrG/a3g485jFlDx6R34jFWqpFvhjNkKvlSfgWHjCvYxonMkjl
wdAXUiu/UDM+vNHP4FyQhkF4YijB5WeaiO56jwYI6WFjpR04OMpdlAZMc0sbkTJc
xcUo101cP1kNwkryiECGmwhJJVPjpfPACjmBZOz/avg4FZ0sFU1EJwcBFNihTfzp
sPDDACQOjGg4gkESVV46kEdVLgxw1Ry9M8aG9YibltbdjgY+89EKtM7oSsvYj2n0
imcM6Ph/L8oQrxKvKJgzziNi+KSYjpU60MsqrDCsewq8TRcJecN5enLKkuTV/j4p
xQDdz8vSAL5YnyGvAKPMMdeWF5EVBxdQ876PfyglTYIZdcvXEmqZ6j2zSp0NBMse
kXkT/f64ogiDNrA9WrzCyLTx33Mpd0TLHsNp0/iQDX4bDPtsPDNG7igMY0JoWvZ1
s/Rd3GMn5tFLj8IhWDTDPj4B8bHVOK6vdVMo7+JrJp0rGGKJ4TpsR9hsOVPbK03Q
ppYVFTPe7gAsfFF8IpJr1tBoL2zsUdPSW8DedKEuo9kZuC6wVGl20oGJS+/HruZu
MaZMRQz5gCtD6xkDDqEhgrMdOvjDPuioPg3L3LPuvzzrhD8RhKuJ5fPt9+csXhtd
St3L5S+M76oMm3ZOtj/w6+8x3w8DlzvMucwgxW3icpdG0D7zVDqkQzXCb64Ygd9q
aWyb37hNak0xSM0HMw/aDFkYw7nHB4pVZorMLtWXc8cTQdUTV4SEWuHpVr9GXkdC
UcfzGE0yWej12mI87e1bUVYeegP2gX6XXEf4whP17KxbhwTD8IL6RMPV6VU6OFJ6
kqEPAOL80+pcB6bHTqlCFqa4TSHCAHYEEknEo0oBFIJqfRDVRgZHgj6UBblb0IMB
Loj4ynG/Sz+VP3EM+5qogt5mxcssqEj0ssn3NxzQRBQcgZFOQ9/yaOj3M1FjPv4H
3rDA/HKks2Tl6SMYRGD7366l3zvrl7JqkutuxaO559PT6hxo/KtBJPPMMYU/Q64A
fFVPfNIvHiebx1xFvIAIc5cp2YW3mEHhwQJxr+r3SPPu43b7lB8MD/Hod2GS6M9S
ZAxmwtv9hcfkTAIA9XFv/YzSEy0OK1xpvJDsdD2DVHw1CCGD0b3cPXwvpIl3Vn5y
eidcLKeVNQeCwYoq+B5wKyUd6Fqfu9x1tB0mr9GtmSMov0/zVHMkWK41NnLX2kvQ
fjnsyMrD45CVSPiteI6nA+iO9hojLbzbv6WautZrcy5fUfzxLgDgKMOeAPbkIaQl
+xvXG1vRkioJ0HyJ4wcKTvXLpoahW3DJDbslKoPcenMIkDnfQ4W7fLQyEilBo9ZC
5bR+bPh+Ni5irvaJOy0o2QkCKv2jlQs4ACwfw0hab4oEpKVWTQHL1bM7gxHZI7+G
giQNRhqV3V+BNrXVOvqbZcfowizpB9L8ZQGJRJWF+NVGb+zgKl5f4dSM3h128E1Q
Au+vxTCxLzJGXlPCpe+PA09yWgwy8INXtnnh9/ecBEd27wSl1POj6/lQKf4TugLD
BFeqjvqc/N/tp3FbTJ5K1EkwAAGX3SNLuCLAdJ2TRtt8GPOfo9G4KEfwPajLWKjl
ZzxrRMxnR5ZC078xk0YDzl6X0Smx5FwKcZykJZ3KUIPe5dIUqZ66IAGWL6kwLNgN
LT+x62MOIkgdkUQy6wqk0kGq3+TMr+KBd+GcbOWKZ/yad81wb8cPP5DV0LSzmWO4
3rhc0WvUvwYyk9r2xRYHqcYFf35W62Ca06ijNH0JzsIHjK0ljxJIuhoJe0q5Npm9
SRlu+WjK0kOHxeodoIyCZQmubYR+XQ16g8lGhkhKDAQ/KOO9Nt/fmT4Vrp8I6Y0M
d8C+ReJue0+ufSqE4Z5/s62i73mGdAQnA0vrejxasDxzzk67zuyRjGc56bRWO0ha
jOT+tKswdj3shWGKEotmTaJGbv4F4jP/02eDfZ+K9yt6L42LyUa0KdDLfFgdnYJz
45BHKf6J/1g4ahZ+y0ZnQ7bN1834zCMbFMJBzBjzseVvCdXzU4BrRkIORQwxNz5y
GBpNtM+jVSmMfPFzzGOFghS1GJxfvjqwsO7YGjAs3Fu+47wDCkCXQh1p7Zqgy9Xx
BtCkC9ZNOgxPiA0B8UarXzaPcNzKme0EUHgP9QA3pDqzSA0CTifeH+NgrZzoFB1m
H+6iWFgphQsTTHMQY5Yy9Y9bPjLAqiOUwE2nOEtDnUG718XfKHPcGbLjsspvri4I
GWPFQL4ku5j2sooZpeUWobiVVBj93A+dp3yAlCmRpIVvJtFrnm7EmVRsi0lhFkH4
j4RUiTYFHWZJvD9SbYfHT/dU6ubCTfzINiD7xjx4m51eNKSGGT7h1j6A7FQ79vRG
LxzkpNYEPY7fLx9KAfvwOzyYYKzS2x5BnTNWKgToY3uBpoeyC0jQmR00it4p+aJg
oDzNb9KGB0MPjmY+ZEpvTSnJBgQl2J2FVT4Bj0kaATZYCj9yNtZrYLfX4c6gkuYj
cWnMpNWlwq+HTAlx2hkohVMS6Zj1WR78MWXI4zX9dQ4/wuKdWAUOpjwdg1f1cHja
g0g/N4qlG/KNNn50YHIxmsTavUB3ST1sM1U2Dj8jfZYlHkcD2LZC7bMQsmlO9c7k
F9oXjTaMnNnmy6U35BvQriObcxDY4BXg3ENvlp1PUN6d8xRIYb+iws+iJkwJ6r3e
uFM9CgEqQ5VXiKjfz0wUvHTGUP8GaYy3QDg7JahJvt6amYKWDk2ZLoI/dfNOlEwG
3Ea0ZKIrT8s60JRx/9r2KVIY0J15YxLam8Og+LRZbw4t/RfOoO5UTscPnXyKWjH+
/HMw3R0ofi1S9PxSnobYt8vq9jiPrOTgMqmoaxdMONTxjVEgAc0XKLjoNAmeSEl2
jFovOSxgIe136F4JWqU6CTT/VsHOoJe2dr3DltpOWWzBokB7ltrdBZ4/ZkNFKs+2
ZSaAS2Aq2Z71C2wwHgfpvzpJ9NW4vFmDJeYIbUimCS0l/BU1W5NjGSO2EmfbAxIm
+NrHJ8RZiMBSEDfWqr/6AO0X5qI8sBesSnJ1yL3cR2JKT0CIAN/Man25TJbWo7QE
jwrYpdutJCzDx3DRxjdwdgzOBxxUMFAgt6nkSB8vHcDaD589dFr4xj7k7IyNCHfU
6T1jAeQUAoEZZfwcCQgwkRD1iL9mSwLwPVFA1ovKMDThrXxfUJf5aRABRjZsBGmO
lOEHGVHcnSbbe0S1JU1WWnEACqza++7gYUhCB/P9Sm64fvarxf72zWz2LUIm6mUB
EtWzZ6SSHVBpZCo3U9TWI4eL8wjbt9ssNlCm/YGeKXhdhWNTZxZctBk6vmKSWZoj
tNZiIiyEzA4QqOxPVtoVKOw16feAxxGyYowKCUUuZjr2UVf7zJ8pwfqkNRqVlQNa
sYtmXzMGdZukx+4YFXcaOnP2wHuyndc43gBPK2hWJRhwm4z8KmhFX/tArmGhuNOb
f0JK1ZKLrkD5Vc/OVwjXstvlNabD1kT+gmQMxbiZp0b4OHgrgvHJUcKAnVS2eGMq
heeNxxG7NNb7cM6gjPxl6Bns6LsUogoWc8oSnrRDpVmiF0UIu6HuZcysWKdw1TKz
24+1nALCQe1m/IYBuYu3ScCOb7mZKrorKc5ZNL+e11TnrbzZ585S72nk3OPhtwBa
E9efmlNcKwsdJlTmZGrcqtDbwK+UHK/1hK1vsuAIGTCRUpUYiv0xgO5xkVM3m4Zp
+H+RRAlFfK1+GvLrU99jKzp+/VSEg4I3VCXnaz3yroZmaeP79vEUwZyqTEAtBVV5
chMoSMrNRccnAPGpCngGXw1oIlSKKHvvkZcaDQiSFX0e1Y7jdYQs3AbmHVT8/3nh
WPEU/NI4WUNGGFgr8AXFajwKu+SoiqEeWHHFJx1WqyR9VJE4qpqCPgRKZakSYma6
7vFIDRFAaPcGli2QVIfOGO3KPsJzmGUDZSyZJpIaoK6A33WWb+dKzdsdaXEaI79E
n9X9Rgmb/RB7Y2awhVPEgneByk2nVg+g/MdfnHu+2HG8O2cCABnFumNEB+Sk9jYh
9/cijMUfCnkpl8M1IlB+3EJvp3vGHCSOSUbhuXSQ+v+Rnaz80tinHCnPEvY6CG14
LvcTmT1BKdNkGPVUEfSuil47YJlMKIUSZ0NxthWAnCZDt/GbmYp5b40clYvbxI6l
NyL5CS9tzDAPGXG5NIeLcc6jXDqkW6HhNcr1TXfpSThpp28gk9QynTmtq5QN7X7n
xUuc2HwehcUuGXboSFKGIkxaBEnezLZMY96d/jG19sIy2ZcibXszpiUZj9eqZlZO
9eZffpCkUtZfFEpf70FatnoCVUKr4/GohXP6aVLNkFBmauOTspVXhpDeqzMKFyq8
FeYDHIPc4zOFaOPR9CIg4bdFFCSmoEdgnqDkuZ3FCowySx6lRhJlV9E6Pp5pfXWU
eCqpa3ebyGCitemUHqvQjzTaUd+4hCoRy/o9hvugNw+nR/s5UvZ7/3v+afQyv9fv
5ETTMY2wnbwZZqFXuEYbHmw98JsXJGiJyj+u6noJ4BNwUYB27j0F+EeEzvHL7Xkz
7fH57bxo3bm7Dtx5CZtqxIJTtTy0NeFD+v/MLxHNUASmEFeM/nNWKNDN2YkMAprh
bFQtXjxoctdNJHGKpoHGQ7N1+HnNGdObvdRiK5blCq83kdjU0YoFHn4BlUEvEhRt
/8EYW2g//sF9ZviEILrwupmaWxldvb8MXu2H0idzf/7t+aYC0Aa9gjfYorWj+q4G
lXhgSjquaWZ00wW5j4eM3t4AppU+J4mjQ0xv9U+xOLG+dnpaip9V2aCx2SL87hgE
D8CMOd45ERL3o44rqNmNQ5t60VoBWAkt1UZ0olhPmGRK9aNxHk45qYOKXK8ZGgxv
JfxwEBt0JOLfwY2cjZCFa4cCrE1nZ9MY3RACJahNjwFZvRuretmPo3Jy/WJE982p
ypHf4VV7oZXpkKxCJWocGh4yTQQ7gXMn1KFrpFB9qk1E9UU9mDMyu/ysuSt16hJX
usVihSKR+wC+RY6qhutChkFwvLsJTIf7noKISTfnvq1QCePZuMa7lyD+NwtImodN
S3oMd+WzSPG1iGXO/fPTnzXZ4PShBD7/fyF6+mEr/pXGcm4sFkBl+2eldD6XUXmE
qqEheqJo/h6wZKVsnz91zw+FVuOPvni4yHn0oX7FzCdki3AlU47Zh2e7lv1Als0b
QE3jScA58jI+zagdU8Z6gnvNxQbL6l6mzilL/Q6m2akIW/1wGnY0+Kd2zD1yTShW
s/8ksfYz8oq3NO9pL6+5W2X79zgJ2ctp3Y73QJBO9FkJXnnp6sTQNIS1xYE6Q8Ac
cfN1VJNc1q2BXxhYWnv6emffpkqSJQO9ncwzSBBfEdaVl1RVJV0I/p+sO/v4PZM3
+8IvtdXzGelaCjf4+s4pWZBPlz+xncGLKZaBi9d50EgQxKP3AFvteoH+Mzbx+/4a
Yq/c4sBr3IpIwHMJ1NiJ8cYViDwbi1FbL/xFVR+qZHBMEFmL43az1velHGZ9XkC7
Dmh+yGIY5IYmqw/hAU+TwDPEfxzTsvH5sGknQu9BF9f9OHVFkWtNAQsVGmbL//jG
UjnBT/OZFPn2DaA0BvduVoxaJxdnKH+FehKfhtz7XzL1HgqE4rmCaqiVSPxrjXkX
D/Zyss6yTrzPCdPVj07Fo9GXSxXng9e8mPEruGqU1tyFfnuer1Cae0X1FIbQaVa9
AF9Efxog4fVN6P2Bgt4rpbMWQkmaB3pK2hdOtP8k5uyfo6oAWU6AIN2p8+8tZU08
cwQj77V3OvLMMMo5QAdxKf/alxAHmy8IanSCL/t/cNzJYDAizZru4ztYy4JlUoYP
HYihvEHMTbNMUyQ4tgtD5/+w/XnF+V4AwIIla5mCTvK7q+YhFl1ITkQwInU7lliR
++Rpzv7Dp9DonpM9FyftmNMnYZ+WH1CCZW12DnM7NRisG9VAcs1dQpyWQKPSfebE
4O0cN0EjfSOpv0607+z/ebc7LO6f2QsrM0nn56TeQULjCVi6EzY++drJ0FqPNIBG
iTNqTYm4Vrda0ugXD9MxRyQjRTbTD2JRtmfgbs4Wj/vhDRH1nT8/L46d60Bln25Y
BUrn8s2+rHWorH53uOTX9G5lemU8BepVZiT0OXSCjEr8lEVvqCEPdHwM1rwP/YKe
11RyFdd3xsDMRq20tqvGW9VDu+eTipSD+S0vFZZ639bveHfnFsFoIStMR6SjSKFh
AqWa4ZOCN3fm22d6SbFpSnbHSWNNBhv6i9FPA/I66HABOn+/F0iIHOm2Loryl1EZ
67UFhbVIONG1EUyevwsNkJYrhEIJ999pTWkHVh//GCeBm7OjE6gBCudJncn149BF
UBteRMfEtQxGoLxDH08qxfGVx1GDOk3lfamoRj/ecARJcmmJPldk1SaToDr9gbmA
S3KX7if90p8zst6GVc+1kTow0UX37xJONC/fm1p7Pk3VVADenQxPDO06lAvqGN9o
gz5wmLRpQXe7ft5SPauOH8KjJ9YTSNfBJ216EUADXmkvkYW548Zt3hakEZh4DlPS
M+vyyIrWVzBt79J+q8OQzRUWqBFBAO3+jP06p9GQyg1Lzeb8CGtzIXhukHlS1bEP
AwM+nAk9siEforMi0JZrnnakkfu1K1vAIXk29yE9rlzMZhM2+LK7dtHz+ySHrJka
bquE+8LEQvrkdxk4sNE/WrPW1M7O6r24+Be5vc0wgzDRSwK3ilNSjaQ9KP6cH3nd
EruxObguxvrr80mCleimvEQvtfsAuAzV6yyz27MJXJ51P8k/9KsqncqXZj4aAGCQ
du9nSZJFBe4OEy3IJiC5jYn5Sx2YWEMDdFwLbmOEVYfvLQs3kZO2Nau9/MUzmPHW
OgGn+qd+I6SOzI+mTtKr4qTvG7bqc/K2DApUpe5L27ol2xAb23Chb8SxEKbDWk1v
oECdXCooz+ph8utcuOhRKiLnvKMC/6/3aDnYrVNVTPWeywFk3N7CYbRnGi5sadDl
oS3SVy4zWeOx7/B3fbUMtFg+ox31r8zveajHbA6crma8SMoLhwcS6fP/U+buMWkR
kC4/CrBrIMr1EM5tL0cIiI+zvLBltNIh8pxtgQ5tRIxoH3yq5+1SEkxozSe//Z49
IOy60LnLsbJ26jjC2e/y3sDOHRsYGptTzrC/rJSSb9ahALp+brH+7P6xUkMeMdx9
iHCiFIgH08M4Tyj7r/G5N9Ow5/6uU0HgDvPBrkl2NKL1X5D3S/4IzGIlsPWI1gHj
DtDpT371hhRHgolRDo19lHbVtvvvHwXyPexwaw7PvmggzsbnrJllR7JPTS8MyyjT
esEeTik2lNiYAqtIZNpXCkmR4aoGmla5BNcWErBcZpW+ka6Tax6Wz5wAUg0Jo2x+
pYq5BdcnDrOL63XFkm7JLsnb8SPX10TYXfvZMMja60uHmI2cFhqqdmgaGOuRpmTr
`pragma protect end_protected
