// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tv3tgLt7bXYopz8U4gNXlO1pKxtRMRjZRM1NvX16lZlMZfkmCYN/XRTaS2Ca2NcF
Ucu++qwdqjao32uURgpl7opuEDDkoSdu6/DmbxqjasgR49nCqDOXKfQXS+goVToS
qMngt/ucDeR3zBlwMF2DYoO09uSEYlZ8pSmFIDztUu0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10720)
mprpwxdmtyPxpNUATyEr3Ec9Rbes4SbaNLMKLzuL5irKwiUc7/pBbAZQjWpSm5zR
GXBZJOc7Bk4VaPmcUy7NuGl8/BRRZpbGZkecYEYn5Q355PGX/x3YDAMTP7AwQf4x
fDb5/AMJnKx3RD/9Uq6p/gXhGLqZ+faIWYYtLlimuRJEY4PmLKIUDXEfy47hEDdw
9EVDrvYS7GE8Z9/qbHa2/ppbe9HAtwXHs2VOPYNSoYSqYsMgxtzs+YTdnz9fOvJE
BegmaVZ+RdjgJ+DBnnIJlTdhjMqBcA+GcNWk3274cLEco2umzecGQ6y107QjE+M5
xJ1pcw/xJnB18r9KiPbIMz7PKgyRYjvukT4VbhttIoQvn6O+BevLk/ldMRhaWIDd
YRsleDEYsh/ImsRwxyBVdIoHQpLsjD+x0/V1C4GI/TXow+cEaF9iaR6BzG2hlgWK
OAmAwvke6hICdzgqUL1RcfM0DNbDUrn7GLiJMFml0pJo4jQnXEa0HcDV8XKpu1MG
vq21iqueRLkAbrDg0WFaI52FRcW8DBox6XaCO4ICwZt9l+mQmLzm1gL5bApU4M4i
+Ro/IDGPTtmwL7rfWod72Yyw46krzqnctcrc3L8hn+7GgeIWQEDA1gQ2FJR0DcDy
d5XvmuE3V7lMqsKX0OU/l4UHiGWJHVQax263X0Q8b6VeuCzzqcS1PP3hTtPUIDdh
Ukw1lzb4tP29CSXs0ZWOeC52rbk30cb4jqf94tcxbhyfHDbstk4FUVeE1M6rDWBB
cU7J+Qs2mVUhntFbyUhVH/3bYO1HSDdBLcIe7KOU2tzN53CY9pcBFc/oywVRImkd
GQqBITar5nOtLjOvrBDTWWRE+Ni6bLawEhias5PbWcXCTiECAukzWoVhTxpBYvI3
S2oJB4q2x9A5Jm2e8EVPDHoQKLhypBrLwOhCXLPuf4Z7ZO8CFt2LAsR94QWKbvoT
SjrhDHpH1M8TPmZZ+mnly4xzwCaLbrJQlU43GxSJELOAmKbsqB+de6gmxl+/0K/0
Q7KFyhifh0X+M0H5XDFBGvY0B3ETB7cUfWf0HZ1j3Yn62setKhXtL/nL8v3iSZZL
CpsNW0nc52byPX29eRX6WoANgWg1caBc1H209eVt29Djy+tfdw0Pg3YWqds+jVIm
42HBgQ9rd9pBp4HcwDGz1PkK4FFIJb5tWA8IvW9aipCTEh1bRwEsxW0xzCRxHuEL
RsUgp9gLxSHxxoSSHDGV5jtWPAjaMj00y/QJQ2aIogVvPGz1WjkncqHHsgO8g2R6
wRY6jsC7Qkfvzyj5+xReX0Psw+QKF2rbre8+TXLlMvXijRQEMWO2LceQlvpKLcup
6f45RQ8CiKRO/Y6z39FIOlM+ExJdRme6vtUlQMR9uHN6Jse3nFuKqFwan0OmjnOv
DNrm6/gYzPhcl5fJHzMoSHTZBK35Vu3jutP6/J96cz1TrKZ+mgiFbUSLuaRgNY+l
qwQKRIFH1Fv+Ppb44AWWYK95uoONoIB4wHaVioOAulWqeWh0NZsjRwtoc9GMtvwe
hXe0wFOokZoyDsQTaG1OOvcXlZmCkNQS+m/4AUB0AO0cV8RWxTUARWkd8lCUa1uU
ifOUC2OkDxsvoOtVTvZ0E3ydNUIpkx7+07ysW7iyf3Ix/IwO0PUabw5Zmuv+y63c
pXZ5rFXw9KP8/wC3VewDxCmlNotOnK7jP6ROXMZoyMc9tDNw+U7JR3rxySX7dmi0
6Xc6pi+btG7qn//ZBh+h+4MTHjTPSKIlk9qE3zZCatKBo5yIOL5gkD+6I4ELx1Hw
rmjfw8HG4ZTrjWFmTb3rK3dRJa3m9zCBpuCIVy6MbvmL6LAheI8RkcBhXuS70ZCX
Tyd1la+P0Kp3eMIQW3ka87tbq7EKyYyHO+Km1YTaIXUKb0U/f+lGkVQbl+CHJpcG
Fak10IEbUDouINTSvV0S7aHeB17fvgpUbNR779kA/ozfrzTUWhXLQWfh2ZHUWxAN
DsXreBmm5ueTixpqsPcz31QL5fkebrpACAGDJRV1bmNy+D8EAOmuVVxzZETA5WGG
u3yRtqQy2rapysI2WHZjgFU4CIDwdmQJPgEPOcW+vndAvROEYTPN+DM1NhWR6ESm
Y3vTR1rsUF8W5KSDjg2A/0KrZRRKJF9lzYqmFYvXQGd2NpPpVTyYAgDy956vTj+D
Hq+fMFblIRZo94S2MtOMROzvwcjmBW2YInlzSk/1gPX9cWcO3SaYOdEocGeTNvIa
pd2yuogjJJHEZZG2FKzf4Mvaxk51SUldGjiWzGbW8DbBB/qFnHYUIL/2qHcnDIJQ
FhzllZhHnf6nSnmeQg7GhqrwXsuzDaN/0XrDUELOjgZUPOWavn00VUcF0AY9pbe6
oUl6+H9x0DpcEIGy+VclcQJi8m9UdMl4HydhTxXh1va5Wv8ClrttZUwnL1Z7s/t8
LsoUmCxdj3W6onfMJpQpqyaBpdORx+Wx5pamJSOKpfO7znGxLNnT5a2VHmbu6bF9
R/ArRoT+Azp7VMOXiUPDjRrZShmLiYvhhWVEqqd5wliZ7rGuRq8uS6HQoYwH4/a7
1JSOyw7z1QpOrMIzWmu/utOFF1R+5Ua1/tI+0VS4pSlCR8PlSJf5+PIYII/XFX5w
CwOg4MSjE6HRdj5qXHmdqN1bQrdLRcnFyKHdrD5HshylqNlRpzP9A9w0Zazx7yVG
v0I8f7scR7a4wuJi0d+ff4WvBQsb8N0RhGhwiY6uADvugbRZfCzLiJ/pE5JvA8oZ
motovyAPodUN7W1PoOmEaNaTdcFltU5LGQ99WdMkpI9SBLOFrTrM2Es3CI032xMA
E/mUtHXnhdikMG9PS/vx9xCeVrFBsHcl8633muMeCcVCPkD5srpxV6b+CdFDoRw8
LLvOdsTEQYUB32zPAYLva/XEwft6D5f08u9p+h3nPUsY2dgOcjKVe46OlM1bPits
fgszYAXnb3k/OwMELctP8OHD80TnjJL1XJ8y3OXJzNWL8RqiK1syLUcWN2Clnnd7
3cGqbVI/TuFygWJhvYiOtLMhkXW5cAdrZzVE0ARI2QoebsNbij0EwwyJEO9ZnztG
4kkfyrk6hogF/u7rsNfdgXMsrZ1Tk0eoS4A4qjQHBkwVTEUdgiCzy5OpNGxCpdJb
nI6ZwqtWRipC6mq5ktIyxILVGXjQ2W2qFixB328Y4IV5U36NBCo4u6WpRX/CfQuf
XKMubQgIyu176PAvxik2LerPq0MZ0Ld8uhcrxDbEXTrbPPyjbY890MEp8sKqhtcC
S/7iQ5aPCdu0scXb3VQHnZzIEaRhpkIlrJmk/kjS9mFCY8Wt1o6nn8c33gCPtc7C
kLQA4dp8OxMISs0CEY8ShL3oWE5mExRFeTZZKgSGoHIqsiyusfwUyrqIJ5jmI3B9
c45SkZSc5AsBah9E6NrZhi9mVRyV6q7eY1uKO8zo0Faoz/NkUGesIkRP/Vd/XoHs
5nl48+Px9qNOWcN7YzgvQjJI5rp7J4dKwsiVCvlIuHji/P7QOBRo1WBOj/zBK9TZ
VG5jKlBYS2w98ZiYTVMJCfsN/lJwoOTpehp8NQ5K//ZIrqCD+4YS0As9F7+eDs0E
ps+RX/yXNrnQgm0/f0QLTR/EDsEH2f8oxSufYvHDP7qxfDUZJ60lBY+g8YL5bvST
d01n9ri+/FB+Rn7BQNUZEZPYBeE2BZvbV/xpiXOGAvZd+qCeO+H9qDyDQ3Mh7b2b
9RCLfgFPqxz+svE7i7iKDWTprHBHcPJecYZrQE2NOXVu8tRGw6ANGRArmmubWANa
iNeoJu7LuGUU/YNg6CJI1v1+4ER4rrz47qZMcEOkZPG2s1HxI3wmr8Le/ROvFWHU
EJ8XFF9Q1yVWmEmbe56VCKppN3PuIXm3u1pZI8e+vkAwM7Ww7ycVPIsCAqQ46NvU
z0ivqVJhnfEHx1X4u/DD/4E3SDkGLZS9jW6ejdfdgXEI+DW4LAh7/u3Ffm/bwkFX
JeTwyVOwgPdM8k8bb3YdvrG09HdyZ1HKYG+N0q/fd1HWkGrLxuvdmSaEazjoggiN
JxsviPk2Xyvi1zsPVysdzXvaUUqOqXVFF3qjVprWIy88NOUV827UoU9bJuP7GSdL
ouZ89FbbvkktC54h6oFXZZE0XXQ7phld5vJglo35HulxMQxslUfg7GVTpEysX2Uz
zQIzOJ0bfw4H8rXrU7bsSjUx4QU90RC29sXKBk/H63gnzfyp7P+0gdcrTlR7iy4Q
2FjDaTON8ugIdmXTHUxirBjc9U0xbyf/GVc5TuXUKp8SwnRXSYNZwYmNodpZGtK/
OrGlPMyyo5j51UqaYphe3D1Bv6hs94rhc5VhZE4S3XrL9rka4NBzBVSUKaIFIAyJ
ucLmPwusiNrtDphsajfqxJhGhwWXrGkTZWra/v9oEqrdbDIUvjLjakL2InyCZyyi
0yN8dqFiC9yZPMaZQGZfqmPbQz6KrpvHdAmgquwMgLMLP/WZNL4SruR8mhXVsafi
amzC88SBgEw28iy2vZuCLA1WcYsr4oiehDXPq1JaOQn5YJ/ik28Ox9WMEXYf1YIc
xzhztBRezoj1R3dHAxF1r5RWDTIqiyJG5Gd09UJan57HDHn9NugU9B/o7WjFF4Nj
0Dqr/VgYsjdjeM01d2u3q/r5TVvsrBtQREOalLbAR9vNyLd3BTYMCcwQEu9d52uh
+SJUmkun+n055aR18aK2pEFMnPjdor+AqqLKG6PrmleWCOgEUnZ6EkZ0DL1aF3q+
7QpyZaXxnkH+zQ28Y8LpFH52TnULqjiYhiGIVkDXPm5YYPfr9yVCN9S90P2hJfo0
AogVltapFJfU4Dxk5ggS0CpLzjn2Ic6cbKBN/SLqI8TT30rP4r1JCUTpMdcx06MY
LkZUJdLFnpI1bPj734CCNotpjszEks61yRUhyqS574zkjcxDhkrP0AZG13RIl/Nt
ZHNHX1VBPf7UoumpAbrKJUlOMEw/cuXE6Yj9ScU8XYpRPiYgvH2kkN5n7JAe852i
PFIvP4Ue6ASlM0oQ0hUyxPKJEZRV7k0OR8wh4CKmf8MzzASVBiYNF8VuTXNWI9KP
ZUqcRW4xneAmJm+wLVY7c0UMYyT8ONzG2WLPMPU1XOgKVL2O3HPm6/+6pMCmvUc+
mnIznZfZSUGedX8iry5Yicz+HCLrKKiccHQOJrZbkp+8H1lSUlPhlwbPX9ZIAvo+
FM9XiIjZmExQdXVmPsNapDxmvyP8/dobEigMOS5zC5a0pEQNrvX8enSU69gKHVIZ
tI3EwySC1RJ7AVRAwqL//SpGM1Gbkgt/590R4FD1S7xOPW47mNnmEj5vEjA3Y3Xk
fiHARapQJEp+4oITxJEpQTwXRiMnJCtUDFAKM1kNNoEikGVottJ8kZPzORNztUaI
i6kl6HpBaSk4S13AmGeQb80R8bRsagtzlsvCihmGx4Ea4G1kF7OKrgQnPtD2o0fs
rODUq8G+eJehxnNcgH4j50Sj0np7E6X+B3Tpl254SA8K9OO72TKTeV9ma/tZ1O+R
F8OEdQy/AhX3PH5HTTuTrlJ4rOFJpnpl0MY1V3U8a/fsL4Z5l8wPMxCltoaQjrUm
YhUQ7y9jlBM8JUblwhipKeTl2zPT4x5Wh1xX/8XGAfmyPkoY7pIwonNX/HYredfb
/vjj4c2C8es1mGwr8n0OsAnIMtHAWHmYP3QsCAryknl3Fbyf/kIjN9rjSpKhlGb9
EMq1eFjvfxDpcJ2hM+ZEAy7x9HGBlsGxayKneZPegvQCSbUfwcsDsV5O1oT0D3yG
vrK9aV3x3TJezO/xSGm2wySMSo5A8erw/mKvMccGimO0CDCB8GVUB650qnjNdRxa
x4cgO1dwTv3Yg1fRN3T10A0t2JCqOSPSYF3CsXbu5WvrlDW12W/wBgIIkrluiwGK
CsPT/u2y/2jS2MMsA9cXlDCqxMXOV6HW7kX1zU6xBU++LxTM6ipnhds0hFG/Pd8R
UE0S6s1abKjYm4uIQKF9/hhWjCGRyHVuDC9aQhxixOksDNOwOHP2aJW/S/3ulQ86
/XcL6EOiCClm17NblPGql1esrgeSM5w33Kc0XxKOfChSxAQ6LcKEBVgO+6BFWdRO
oVrOX0uy9CJA1S+FTs5dKFypKnWjP9WEzbu2DFkxgB9Ld3+U201OmZnx0wZso9ro
YAsrCFROf/wNVByM99AXVcRYyqXX9JL/42cc+Ke3k8bOfDJzL4lksMS2xsMVtUL7
iSA8S2682TFEYms2RLWpkSwh/JzZf06jxUVwsG0NA22KNhoHl/w0J5hilfxZcstj
gstq+YosNJDU6a+R85fPZL5dOwzj8GYDarIDzkQdZxb6IC1hlt30WncKZSjmq90j
Nyp84CPFEfUhyzVg7JWu+8v/PEaBem/4R+W98OJ7jds78QBBiFj7Fufkblb8Q4pf
AqxSBjrXxZbuCYGbtq8IX33ohfK6wzzO9OA6sOsEARcND7oYee7SIgrYwucZMcKq
u9IgsQybdB1gAJY2K+3KngNYd+w2H1TVL52AEJF/aBrUWbbJChZKCV8IEFk564QT
daLW1pkEVpplZue5APeM0NNOl2tZygYTb1VuA/jXbSx5r78zHNin06M+WDb+kF0M
nNXD++OVjVpylOpurrkj/ujVmfwpIihN33BMVROh74vOVtVaaSdavVeIWjPb4Eko
9HwT7XVUHt4gt0VOIYdjXNC7h41DOwz2ilfHBMU5Y4bM7mEo4uGpgvxQdXwV4hg4
vVUzA2DqHNkaJDfkIEanKU6k2UvfRiGeYwcy0L/dny8gTIKNXqLmf/fdHinbrls1
WmLwBrkumHE9tzRywGZ0o9BnWCQWOkbde5zBsRd9F0Yc8YCTJV2cNTWga0b4Wq5t
tc7Fsx3yITH7TKoknh7lGQAvLNm4nt5IGQzdixr6bsGQcY/E5woUOG/bBYIX/A1t
PWU8RTAC4YIGRxi2cuFTdO7kk58mKymZRlrB6lQ39i3cEOQLRCJNwYkfusllVQJH
Hgi/Gw3ss3JdG+47TaIv1rqyg2EK37sqv7WLRQ8SXHK7KZZ3tRLoMVG+HS1J1MAp
4hsbCJ0ALByNvTr/UmAjk5oMTFpkgzk+VO+gNIzGXDhWJECEgVVaPWl4FalEah3b
xVYYrch1KLUuC+glhS+TQFIlAd82Z+EO9IGsFXz7oiKObcROOl1/LJjcjxOup5ri
qDo5lEC0zJG4p3WsfP4GbOJLNtZ70vDTL0vqzAyNjpIHgB2NoD6JMHINzZZDVAUY
FWWwOrVPWC0Y7Oyg3fNgU0xOfJrb4uQaZW7yGstgFUeIs1ePFOLb+mOn29qv0WT1
BiJQrajKDXyiaY7hZKFbZmhx9l+qndAb3zdKyFaWINLwAx18b9tGMrCORmjwP9Md
oZ3YCECcxHzkRlfST3wKqAB2pgv+u+ppPRY+BH32B2W25s8bhQONMXyRuLra/xed
jvVY7VS+pcX+0o9z3YBXrBLr4VyQ1L+KCw3ig3z8B++D2nyLtWAi/7vcOyIzzH8W
oZ9YWtlRPhrGCed+uBxe0UwyZt14+jYVSOK70IzJKKo7PJicvs5aNq2V3K0s1d1u
QMo971Mu/8av+B9wFHrMANB8XRGZw38IwLSh4juQh705g+qV4MWV9T5fOdlYMC//
F1iIZ4AG95/CL/+hTlnGZ+sG6M6ViuRE8wODc4P82+mVBod4YuvuC0YngjkJB5ea
79gz0XFNPGcLYOjL/2CQ40pSeD4zUZWgX9Jh2t6janQNPMJ0THPwlZ8vF756Y+yp
WNrKhR8GJNDgyn6gEB/jugqNWWjsWCW6KFySMrieCmfoG7NZaPgIUlbajk5Y6MPW
Z0lH0QjPg/BHp/oyLkXvgEcOLGPsTHnXUcUW0moOH/oGKvn8noMs12qeiVVKd9K8
DIq98uxl1gdbAHS73ocNgHhFBbNJHw6bWdXEdoIuqK5kdm/RiOJzt39KNyf3iNGQ
100OjfRiN6wpUok7smTnCwgf6jpri6TwePbxiURfOPG8q024GkRnW1kmzl1guKE5
R953YseQoz8Jr5ypw7YXdyAqigzlq2e1CArvrp8AqxFcB06HPay0lHv7loV3b4Aq
q62n7ok30N7Urgzd6jtVH18o56liWrCMhWwPryXALTlZdWbh3K1A1e+a0Sbw2xdB
cDWO70pYYRo0huZLeKO7U3t04LdBc2/9CxqE2AXs4CM+l1c5S8HPMMiKqJk5p2hI
Z9o8hN1EedZxKOYlvHFEdD2WFtNGi0+q6KUZ6WuElKImfa4wEWzV3ABwmq2MlHGx
NA2tooEF6vdnckPRNwN164B8fn+4rT3KTb9Txjhwg0AlJ4Akg4ZIpMV5WHp51/gC
AuRqHHqVaWXxFxh36LfMm0ab+kN4Rhc4h9MAkubfvbqy4qHD5UmVfPWPn2sJ8zor
kh/HnA7PN6zkFHKiqH+zwPvX8LVfJBzXfKrSVtIYePET5DwDaudE+z7c1bs0p75t
veAxUNcobA6Z/5wxpuadvW9YQ39cZik4eL8IgKvKa5gbeGXHUJU101K/KU+J2lfo
hUle3ss6jtx2a5NdzM/Gtb8o+GtZuPDsp1eNsHhGuH9ZSDcfm9nGLhdD3eOIvVCz
WJg+JhfKlmD6pFZsgODR8u8A1cR6Zaek4c/F4RWzS1ZFKZDZWsKtn1JJMOxkz6ne
YAysqAJYX42QsXxi32upbV5dFa/MDCGzzR4SJZRuuR2yvZsyrKnjYK+oWMiegcbm
viI4vJUF5FH2YgTJEhNzPgLDe2CfsiuUHC5xKGSs2fPO5s1q7NnSqWPQDimu+YxN
MGjC36mz+UhpBo/5/zvOlbjfXP/Kri0oTGnxTsBtRpTEa7bQKfP4f2j18vr7LCha
JqVLJM/d+h9HV9Hk/lT46ReQ6e1CkkTniJNo/M6KwDyWUmush7bwKPUC7xy2w4HI
NJqSXdi3ckdI2MrSAcHqh4ItZw6+vTZMC2Bgkp+BMna3PjZ8xoVyi+g5ltxJ0jJu
3Rjt5tfYaVd5FgV2x1ECmeYTzS4rRS48aRJ4X/+m8zlReW24CXqVsouti6yBZkmB
Qgg0BkaOBDwiQWb5nGEYvvGK/7gB4k0F9cpkctS2Xx4V8xObvV/FhU3xb5GBkPTX
29AERc4VCFMPYPA3LlM1np980rxCe0lDHccGS6d7ZlgDYX2h4KYUUUqg9L8fR1mg
KzMXDrC53G/04qGn7kNQK6xzFY9LQ/LhAv5PvIsnTcKpZEYIYF8mb/36CDHIGSVK
ktb2kBilA4kTMZkhYo4xLZPGo7yhwbs/eNpAmFY3npv+LsTkZ3D6SIJskMuM4sQX
3MuDH1Yybf89FAp/NRyhwRjux43b7OxCmACL8nV5GYcSCoTW53+JkjfQjpWiMOB0
2psCFhHXlHWDUEvWzw3RuUViqWtSDxpuW00foDXoSIqV5eCa4IaIn7X6alrqOr5H
1HtchjoF80tixHJRaZe5PygbqQ6blR+VeMJl6jDey8520o36gz2WQ4Gyt/BTL+EJ
i21kUq68wpeb6g/59HFOoX9e7TQdhOVQ6SZGBThvOHiXo3ImjFaSyQ+HesgEVWwt
K/VEkhhd3CnAqEBSgMQuplC49auH1y8J/chL+CmGtt5mqwG3EEeHghUWrkvVKKQr
eJHLPAuGzJ5ChemK864NBWUaDTrP9QYYE/pLcLeTjtGvdBOgik2RLyNJ5keWl2wG
k+xQDt2TPyXEmluiIH23HgRmRZMgVR5psSr38hLIhGBmUCyMbEJiAY1ydWCFQdQ0
fkvaXWXPfDt4+Gdlpqs8RhDwgJFtZ9l6ZySXKmrg84/ZjARXDoT+HcsiYuTr/+Zv
GIRjA7e2m4Fwy+OiVF/Db5h1XbM6K+PJJP1C4LMufgvPvSw9hO8R3RgljctlKcNG
Ql2Plaufvu1w3P6D2vSLMYmtSJsY5ZUKh7IdGF6zXBnkqCrTkfOQpnk6J6RoSR/2
W0cmgJ2SlxhB2queB2jwFhvboQ9jazU6OW+/8JyUOMcvUoUlswGT5rPBhYBUGWYC
7o2M2lZfo+L2uMmBkRdmgBMZwFKDMGOOvxvlaeeL1Q9C+5Ms7eEtu2qJvbYwNfWJ
klkKdQTLuL4p14Zx2YfHSapaYr1fU2wy9t9P7p0a66Y+KUTQqVGb2usMQqR2UpG/
3OCyt2vB1s2d+rK3SWSsoF1yTzXqnJuKnWECNRHOq/9ngqlZOrH8GuwYlJzQp4nE
iOra7Oomq4GO92+JG/GXXXy7MeW8ToH6trAPS6/x7jn6gTaXlEvhHrINxKQouXk4
5KmEC4auqxqC6Q+9wOL9zIW9pWU4yiIcTLQU0lfzWQOraq0a0WD69k5e2gBbcotp
oUUDdaDqsCRbHKQW9pnalbmRNfsmTgg3zFj6FTtvN5jmQVlWtF3fyPiBQM4XPEZj
7FCIbKdKcnpX/YERCaQr1/bXqybQ/SCM/OLsRRP5IMQA1lYJ7sK9yTVO/1DPqzef
zV2FzeaUOkjNYWy2KpBlEbJPDDvipDVLTJr4OUN/B++7Hr1m6tNt4ouIulw6nRsX
qzSm7czDBusTNo1MXyNENU2qCgrr4k3rplKiXtfUfjmVjvQRJWoFOTSpWCV4jZFD
YT0pB6F+uu+K2LaQY82pyin9tibwtJBsgmAiQex9//0DVQhfVmMgiJHzEBeP6D/N
4fJ+czUcgB6heJcmMLbncFYuxUCsFjVI//XG6Ud25ZwT0kPQ0Ql9laqc/gJUUmBd
VSPa1E4gaaQjbyzUPZp2Hgj1g8+pmNuaAuz9wx7pWQ4CP5n+joKus/03kYfTL+D8
VyqVJIYkYiLR9vo1zkNuYTYQZkViNnrolBdTfAec9E+yD/8+zEl5kY1ONyFuJbug
Nk95xVUo61RZCyvHdKdLpTpU7cBgfhw162VjQ3WRhYesUA9eirA0WamxDDdZ2SyA
Ml4OKdzlDiJhHxLtQGma/dzNETSceRQkpS3sCWrcRZf9cRCK3U0feihZ+Y3pJs8D
8OdEbD4dp5hJtf8S+CutbJrbzY0oYflJBn3fswDwulQZ6vrsfIOcDqT173h6W6W6
HJNTVRcKL/PK4ScYJJ/RJgjwZizpcn/mZn9V/CM2C9oMH96SBcxIy/evaVakWS+F
oVc/GSjsPBN0aGwVTi8K9MyxhnTvh0eN7zqvFdLqRk+AEwRVJ7GeBHPF4d3GG/2d
03oeZe2U0kWrPNek7zdrttCP7+E8hd/GywZpysxhtcgjB24Rs23nwQeALlEUPfOa
u2iQ9Hb0M+m/Gjs9bIokT5uXfnFiQTJv+2sQi1EVhCl0IZcGkzvDL/d9euOZ+ir9
r9TqnILVJhhE26OONKo7qmAZLebO2GDT73cjGaz2w6zfAGluLjaWnX2eFV1wvdDa
g9x8kqJDIZuqvfzAAUNH6ZxNGXQmm5OE899YrwTI8e1HKiBshrQEnUzRDm4LfKi9
H0MyJaHdRJpoAlLvbJlYtoBEtvO1BgwRm+Dd6/gZ4XNMNOFJCANqWvKmpP8SAvDI
TponOzpyuPA48pOBYYds6kNcgHO+iRXOuIS6+gwSxzchLMG0X+TAkvCGj8vn+SWd
Z/bf+ywLvbN3PGmfvnju+I6dPIYzMpLhi0Q9FNiz6aJTNtn2Vyw0kwiDlrX22iPm
pYWfJguBVrgMs1aKnXPsTZxGBPb7LUUXNVFozX3JcGeyNltacs5H9myEWDVlkHgm
ZxDdwwFyECRj5iLRcihdoT9dfUvv1ZTrCi2DNGo9rS/nkbDH/3vCc7NL0iWgM7TM
YwGirROvUkYty/ooCa1ph+Cb7noKjoQAYR8xVbYhNtDyLLEddzrKy44oM7v+kNal
O+EVPO0R9brruhXHRuLCdJTa8Nd74K+w16OjbCPq9Fwwzh9ANM6d5k+HyBITI62I
yby8IGzov9AsiZ8Om7t+4EKruoyeZdCCscDYk7IlSjE2d2dkNua5SdYFTY4Lwnia
Ho9vvpHDem6hhnBCSuQfNnPor7u9LUb13OH2fq8rwirviwAlszZU/czF0ujC/7uz
v5CEEV7cLBvTri0YaheKV0h2W04EF3ndQq+fXZgL0znAr8WbqISnsPf7NcK+QC2r
nwvAf5Yfkgo2WlXQDshqYOlyMYO8yo5abbiIJFAgW3Nrs4jWDqh611AcXN0Kctp2
swOf8jyavelYTOQ3idwZ9s0DhwG5sBISbKvtIIwaBh5/SfPFo+jJcqsX/RjZGGgr
UKjEoX/uo7xYe48mhPuVZ9f7UG1lGOPC2wdt6oLS/kwc+O1Okh6vpPgQUOnP/r/j
s26RJwNZceHfv3pfOXRseVEG0CN9lkiik5BbRkutZoZ2sl5grWilGIZpl2bvMtUB
OwE00ragrlEMTtfgCasS3VNDTUx+gG53TEvGZBdwBVzBYsOpn19IYQqf+9yVxT4P
R0JoJBvGtbU/YCfMU8I28ATb12BuSq0lGrfXFPvSNLHMF5piY/lsREglrdIEUNLx
wCJUPrP+1J9W+4eC2QKBqwOUy9AaQp7VfP1rnKvKncVJ31lVUHkXjXedpZDn0zV2
c709rt/QxgXNoUWBSdyIKhhbN2MPVDJUH2hut/dNqNLuEJ6ZRtGS96Emx13R7t78
iKeLKEl+zROo+0zkfukKMdJHrMWuW1IGTUv6gRsalWCG33xW9jvtQYTdB+0dtg0X
ThEVE3aGqxnUZSlPN/p/C0Y3lPx8ZvbeTm7sE6ElyEwKNXM2hQounTthNXBB/W/s
aVqhGv+aIh4s13FPLWuExLZXrp26FsxeHRMh6HMnBOR2OWj+VC7yRrP/jup1rh1X
r0OeNvAIOvlWct4BF0Kohz/rsVmZv+15puXqKOdWmD+u6CZcNsK/qA55/SJ+at0a
ypJuQ6E1uo+y8u88yZg2YEaJX5TV2kZIdujD1heLwUQWAnm/OgcifQkiY5yXO514
5jLpzRBsx9kZku5yjkDUQbcmoFaCSwKTUapbJitNubw03KfQ52MFweFT2PBj3TLp
Rd6RiWe5gZf5SkgLMHChUV/HMbS+fmyCQldM5AVV5EQXP9y6rnQfz++gxRHc2qOT
oc2fVHRbBHCg8wqhZy4tt09JitpQ9qqvYtNOlxJECWfT0Q/8LIvqjs++/pTwc7SH
dTGG8NT109o3M2YfXfhrOYsJw/FLQGP/gHbIdD9oXLNRD9kxdX/G5wtdT1MHfC75
80J9K3/icp/juFt12Do5nZsZB0DzVARhYvUoBnbyaA6B4pOy8/w+XmH0iPWTl31l
9fijjQYXQiToxvrE8avMk8erH+8IOdMnwAocYouJ5FI01Rx+yhSRYO67YM6SkRHg
jUhaBp5SE4CaEqBR0DI4g18ap89p7Eom7lk1ZlePar4l9UY3mZ5bHWgTANQkKtim
b00gySHOIlUMVR+Ugen4k7T4nBQ5VrDQd8fbKPdgwArmRfnehXTduEuxDVdH7kQU
xFoDncgKlYhH08+/7eXb7EgIVyCCIVjm2u99/nTbdBtwzdd8Jjf1cs2LOieBvnoA
A6/rgckOHmCUCsqt7z3rZgHfNMZvmrfGdhHSISzJce+bwqa6NKp/3zA47L1orsPW
OA216jISiZl4ikQPYq4zaj/O3NVUbUKAkxKMCo2xzaZsVmMh0ktjX7ScPJFH2Vly
lM8fFxldzptAHZyQTTXQurafHnMq9K2EtisptDJqNUqvANsjud7M87Kv1/KPBwgu
5igCARFjhuDoJYLi9pIlNNKPOc8BwsgkqfTx91pyzlKtpY9uqgSQgXLwf3ldo8Et
xAJS42GX1wobCSUeoTKr2f5lwfHvlM1+8z8iYNqqwhADnwPkFHRfEPJ8RwRzbNoF
S3KfGFxixEPzxo2AJCM1q9tXKcopLcIIBGP/u9+vgkJ7K4crArTT5s8DaoTBKwHL
H63ndEay8fNxXZv9469nSl0Tm59ezwBdS4sbBjO+LdAeR7N7SP+BKztr+GuFeFwY
Dv7vhnkMJWlv2Ut+QqbiEPqP0RQyyH87sHWFCQlaDyqypIUjg4BEG10/7NrcpTDK
Hk7qV1C78JU/3QgWuzesWX+Xk0pI5nuje7WyccwKjIxEBTPlJi1tJ4qDqHMQrdHP
X38zV73v9Ut67SYx7G4kQh0jh+jeOZDAV4xTHSIYiuePv2/NYrTUarwnni9w9mtM
I0VkTCU45iPNpgi9dSTMyo5fed3PaqZYjjFpmLpWr/Vh4AXb0FjjUBSPidk0nsL6
dlTUrj5yRGOTJ1/xj1vWwfRxan/8aAEnS2ffzSQlgjAQAT7nBW6VdPTwJZvkC449
rpDZh4aqZ+zuDDBMymoc4zFcGISD6Y2fVGdQMN0G0K9EzUvlwg+BYWQe2zXqfzoV
BQ0oFMxUfXiTJOQJvsWkig==
`pragma protect end_protected
