// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
M/1e8KM4z4EoWsIw6i4+5Mt9ddeSxq8fibU5KVKzcM8Pf0aS+TbwZeGgeNMLtv33cUTIEX8ylQBO
uPeexHXBkUnePqBWS90GsDhbbD258VSg52JRuYIo4uTLr1Its78E+iv/r0MhtC3a+25CpzuSns7h
UxNVA/2YxieyB8ECtAkz+isg8pGZf7rFRpIepTfobTKenPtH5aViUohM6TcW1swK5vK6lpehFUWK
Uh8LhkjRRVKmsnwpiXD28tobdY10/HthnbrZYrPJeeY6Jtr5yZAqwt18lDLLtOLAdX6rMWxTQV6d
KXEUhnS+8I97zu08sQeha089G8VkoYgRVkRABA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
UWnST7EfaqWnUhYC7EpOoBF0SXcuedpWgFjdfaN7ASyQh46Urxh3YnUy6FHmaWqTBFeMP5ikC9Bg
+3wtQ9mV1a8VMXywLQrdv8Q4FbCfHvmZDuQBHtEJjykZRGSdCeaNqpS5kwMAKjHBoH/fQ284Ohr6
IPKGs+o/5QPfJXRGo8ipVk5iEIK7cp1ZmpStKq6sLz2UjHSHAg06axiuPG3FMNJbmaqJY1+pg2Y8
g5ffpQ8SZAugvEbC/iA909AuKFZuBwGcJKVDhJ02smT9tFcd81An+jtfufBacC4ZIRrLsKWOWGbr
lUdafCL/S2XhEqr1Oq1m8cN2BLaN1/6bj3rG68z+1out8zDGRv2S2AMolhd8gU4481yyYROf96Bd
CwSEjT7dfFomGIxErhU9/PfFgVNN3FwPb4Yv0XG7g54b7NKmlcqTC5OIl6R9NeP794RdvgCwnTal
jIqcB5RDBQjP2UOAnE0czhJLP7D154XxTmkGkodpJFihE+6k36C62RWDM+e5qdaq/z104ZNCfcEb
UWtVud6T68dlyZS2Vmkl5PsKr4kh7Jdpe4gytSLhXm/By8CpIfDLiQycVX1GluM1YuvM8vBs4vgt
OAY8xUdmr+7Tnps/ugmh6OtwFrtJNoEhcJLm+LicO97eQLdagbT3hbIa3UBo6V7gUDeGm2H/mZA0
InBATsIw2YEqm58LAt8A3LKi2Ke3oh5wo9eab9207SlxkWnKsJgHDWcew3W8UH/qdZOV8WMliRQx
jOgJ2U1EHawLIFrKsE/RzFSaLyeoxoWu7nELj01P0fFNUGqRQ0h80UnQN7euQTBB4rKKblSqEkhv
4xH8Z0VRjK+aLrOCqWCtQHYLfoD7/BiSz+1rCNuxg6eXbYaLjinUsY1l+Jj/igt2Fj4uiS4x2yW+
9CLm1Q22nxOHPl7ISpu30nHcFwAs5e8mACLf2MKcBpn44Zeh8MqUD8TYpnpRexpH1cp9Tlj7lJku
IRLQpSbKJ2IS9FkzP9R1dTVVlJUlpB36sFP25PWjoDxF5oN33ku2gaJr2KNEetEXW1MLS3Jlkpu8
5EuA6J1l1yzbNOj/pQwEymnOjnMdDoQPgSkrObOeRMubxcO5aBBJy2bVhf49ZnYam7YuGhhTu5W/
IyVLB4w8XIVhlwn0rdFmwunWyFE2c3sSeJYyXAHbxUasYfNAwPp6MS8zlkG8DFqJ2AZGSpxk+fBD
AgQD/cdD11GSgSXZqosibrnG4uWMIw/NMDQgiLevjxFAdkWHfye+l0Fb29qkha2gu2AP3k2UYwgg
+S7su8+pBfCT2yRhbE0lqyqnw+7GHWUNStMxSSlig7Tj/2jpDIdUc4opQOMGOmNE2WQ/1LzegPO/
AmeWxQcmLPVQCpT5ipWiXmlv5IuDFDlVMdomNkBNP3+89EB2mimCpCIxifLMsRNecDwyOFJ5Q8iV
2wRc9BpskfQqsH1vzBWfUQ9XzUqiV9P3MFRoOYvyVCyNDVj5kVbzty4uTBvXq20VDklVKIBNprYS
6uDHQrYTpwG3jID55vUEBkDqjxccKKcwTFgdeifB8DQZRWBvRSFyHZIlY0VJxQJn+IvbJ3k1s5o3
dvlbAXMbip2HFxdUXW5xi1JkwX1+NFHue9OUn88Qc46v7v4jwDWQYiC5mJOgRN9V8HwesEXoJPQc
y8SKUafScyz4nX4SSH3GQ2jxHLO0nzW8Gv780oRZccrFVoy85p/dCugqf2HBhyF2zj5od8FkdBRM
2v0erInVNxnMG1KwFBDUzwd9AR7D7KJAHI8TCyOWQDaJ524Te1XfRoaJu32+q68JCi2dKhys1xb7
cMUPI6vi7MoONkbOF21kAxUYnWe6qvcFTU1HztBQV4tMSJmP14MR4nFxBPGAYChscED3FfbECl/5
xnuPzs3Pam3ar1aITlB83Nhe1saU7/gg1A5a4omXQ8A6J+e4W/AuRh0yOr7AqvoOrvLM4aatkaL/
NMVp07C2sRdK9uBvY+2y8xrSNTV3gcL/rnLzvVnv2O4cOZlFJJTMrmbRgHZ6PPLg+FsKE5nORFkQ
E+GWC0EIf3b/jWkyZbaqaCM9GfGBOuoBpXmA6fD6F9Zc0HYvoEriofSU1aRAMulyf1ObRHEjuE5m
shx2THQvgi/5Z52OmnzI2h5NTRq1MN6zExJ620Tpf98mX7Q+kzb/4QRAXMSldOWldFcsow0ZFIMw
ZpxI11fkMr4yrpusVrcMxXcD44LHOXTA/yG1iYcaNF19IxSJxqT+s+5VtH81Quyd+SSATTcvwIKX
b2TuWF6aoyoEUNWE0Cn0kzGVsZv9VGdNdBehBrdX4ekGjUfBgAlR1PXD8jHLFA8hTa8pjM0877EJ
YLvQABVOr7ighSNEmnlEBbZLsQ0TU6577wuLu8CQgzDiOa19KCkumt3sfLnnzrKI/cleRGMxKYj1
hQdwuvUUYHe/Q9bGKXi7ewYe8Y7gjcyMg3OEvI8R1uQf/PVVDDK2d9FBjdH+53A4d4WV9cBuulbe
gC+X3Y3SDOcjA2KbYFg4uGwLa6DE2NJrytie3eBOW9d8eGIIFPvfqjA8nvhabkQzZ/BOa+i3hcjz
8EEbMOqYZCor2ZuZpPhjHj13UJsZv4Z6PaUtfX9Ahnvwo/xfO05Pb2hvAAj1NE+4XTUoNigvuFCt
yyAdYKAN7PHnPIG7kB3sDjGlrlGwn7Zr7HVNfzFA8UakTsXaofD4MVSNPKXpDG/nAzkAnX1SYDk6
yDL8jCdx+Z/N308T+1mAvUekyirb1ayuBMM8PdrDya+lMtyHi+GmwsTdjP8ig4PfSqPgTC4q6+2y
n5Hl0qeolrkJaxgEokla8Pof8HFCR0G3zDpjubm53n2vdfNOn+emYFMgogNhlGZwIRqLzs+MAohe
siIZZKHYOtQvZDzTeX1s9lSdXsKfdqTl6eUPP2ACy7l11knIcpBpealL0xoLYGfM5euqwArBysuA
SDH75L32IDu48pBf38rpPbkswpQNBJ79FjcfMTPNhnVn5DDgbvQ26JoafKMsROvRJ3a+eV2QvK3L
B0BMGhGH1pfNJLObrpgmsyAqHl4E+ymUs2dTZ42XIitmihX9jF11Alzed3pLYzITBaJh0OCVfpEE
9PXcjlDcUfpoPrxp6RhKxYU4zYcwleyPXGqJC2Ewk/WCTWBSAAjwcoWI90nLvkIKFlVBdoIUjQaj
pOdarKoXZuS8Lugq+RrduTyC0NEziXIo9BRgFPt8wxAMJAGHZEOOyM64yucRBvzn5etP2NNF80Ee
Yq8qej/mu5KLjDTksFi4Ur2m5mymWSq9EJpQTUGea+J+PzX+hQWchaGsR+hmXA/IplfGT1wNoWJQ
oDDqCCQ64h0VOkq/BPYnW15cq0os94jZCtsBWvWhQ55shoGGnoA5GFnQDVtvnSeSNU/UaCgOK+jW
vVEWdsXkCqscVSIB9vBRkOsHxwrB8ftsL8rM3w85o6PDYxlXh4R8OyyLw7sWSgyDA1HF5IaQ2KXq
UTmhJTbUf5IslY+flz2xLSI52FJqncAIvqckMBIW1qLbkQCrZ0QD8J2IVocSvTz2/l431j0PasTe
vZQX85gApXR7eDFtVcwGbf1gKcs0dzrlQ0Vh642Hc20wM3rdDTMrWmT0LqT1Rb0anYB9NocK4CXp
1orUgi6QN3JxEhnUPLKcaUbhh0bMY5gt38LLe0qtc61b5uPsRC3hXjM/TvCeJYNXRNl/kypO31xR
xI2tEv+79OCQjgkMOwG7Zm06TlrsYZN/VzqCTuYYUozonZe0/5DxBQjC6S03DbAMTbqE3E3fMJrt
mPu8AD25ofl+UjLcu8BtqRibvzQLwokQ1o3su6ejC+Ho3XX0sIBZM+OSIf+AiE/9yseyFXeXRdoT
Sa+Sd0f54uBXbCfE6ZJ71Pb9bqApkXMbGxkT4R+1j2waW9xbylxn8rrJh2N7oPN/HzAtZlGNZ9S/
csbBxVqixDhaM2muagsb1IdRBt1uKFk3igpnEg/+88XIAkaR7APfvzfrc+W5FoONZV055TlCQvXI
bvcMI/2nnVRNNZwvOud5MhxiOWetFUdX3PuMWcxw1htARH9YzD04czzIOfW+WD9JA3thaP1XrbiS
Jb9NzF3q0Jh0TErKisrjd70xG/n0Ok2ohDu7uNX3ZoEUjU7WAYdkp/I1etOOzxdVXdl9fK0BiOPu
DM0NJ5Ho0f9i2RPFOjhl6b7/DU7ngcag0bwoMkwuQGSJOZ4QZbczecq7ieQd/HvTd0EalTWymN4y
bTzf53M5tC96Biv+gIMeWECevvLmst+phKnz5VQOjzlJkFEUwru4pGyD3Jzacd6BV4AA29izkUvS
C28mS+xkRS1b++W0dMMFaHn7s7gaGgdoXiBKGyd+H7DfPaHiNbd7BKUvuM3+vMjkVp/MO7NREgTc
H89HXtYMMSqySC4OXo1jdU4JQw/c6/5h7cs8xcAnan/9ytpEaGECk8s967mdx+2c8i2K/2PX+FKo
fwukDW3KtPODI6GpGmlmgMglxZ2vZ65Dx3HRkxWKx8vi8+ktgHUAxUtB2kZzmJJ6E3DDdpA7h8wW
4os/5egAJ5UmgNYAAXvMzNi+Ib1rP8xtlOg6tDLF+r8z6JIfzO0xFiZHRcxaS/q7WP42Bh4DiwQy
Jt+2x8pIc5L/Dl3il7jLsnWIFijepOYroIEH6hR8zD1uoqKNa9KOeu8aBVf9vOJaU9mXBeRZ0NmE
MJjifAgga+Nz0yP5t7ypq/TwvrVH2J6cPQGfZpjJzge0sufLMi+X1Skb5K8u8zdrEixtDpCXRORI
dy/54qSZNQKUZhMpNounRZN0sFHNz24hUqvYgcfc0Une6EJpaxtWfZ3otY4uMUaqUQ+il52/3oEL
0tVG62NIgpTvmNit9N0iuHmsjpyMVYX5nGdDfeo/SdPYFFQOEz8sBUpvjQWXuwvQIS+2wwTMnkky
tKZN7QcU9Vxsv3+Ao5ckVLGwICopA20Tj6xQFVmSDvshbwVjHG689DS9oSWaWzjyvx6ERmFa/ikU
neT5GfWebUR8A/AZPiMptkSHBT8yUMuwfMtzSnlXIrVt7Pp5NPp7HblDKafIEOzRr5tZveV3+U0P
6BkkuJpo6M71zo9ZTCCTmp7LmSlL2evAsf8Ek+zphCmhU5w+42SEdU1LPpljGzIj9gHJZRJaO/Yt
tGFhqiYhWECUjO0epyqhqIf1DH4NL3kvtjGJjHOF55Tew3rLS2zr7l1dfrVyo2m2KpLlyOEdyvaf
HvX6AJzY26zCKbX5LVhHj8tt948S1qeJZFpiMAQKDmkBwGy0vy3QfwG+Vms4FfKsjloQUl7VMrQQ
n5I4mYWDgy+raPWeB523SHnH8KjLIhZmVjpMaladxHHsDfMYXNcLcEEYSLmVDHD15QFD1R6Ysc1s
BUul3jEH3eNswAAWCjN70hz2dkKHo7Zb+1EF6xfQ0hK0O9fMi4AbMP09DuBo23tSOpEhnqFhvLP2
GOx+fFw9fH3aYXjJS7GslDA1kTcZTkC2EV6XKJ83jW5R5W/HnZPlNy89SrwecUO/awnh0H7YuX55
lT/zzjMQKYeAZXuigs9DCropSbrurKaE2LNDSBkweBVwmHw5q5tnfseAt92YxHR7F/AXNG30XHfu
y0aLqmWfr8m3jWsgCO6jx4R6NkggWPi947qPkweZIlfWgpcwGxCNtZ5U5EYEyXTI7TrT2icRxsJS
dKVwqJaw/om4XW7r5kAwGdqb7U/iNLP9fYfgVfoF8RMvLqjG0jVmJWr7ziJi8CmhoFBsufI0LWKx
NwBXmJX08gp9hqMyS/SnrzIXEg/sp848yp5Byfa8zUQsx9ZYct99kzLut3ax3GjaNwWFhFOQleC4
h8gjRi1G7wtgw792YSEwguCJMbZDqjIPb4FbI9eoAa5Rj30JbrrvaEzFg7w0beTwjkuNAMdR9IMj
0g5Coh/ZVdap61ArPUr9IOdS3yW2RLdn9f914mtnUPUwnjQ3Xb86nrAC5Vgb8XkJ1Jn8kxnOr5Bu
o4fE3xNm42RL7Hcfzp00V3z9YEWL7I/hkrXxCLGHHPkE4m1iQrZ2A9fbwTu/O0/i7qCyLB4XJxMy
OFfO+l43y7xdMcwIzyChgm1X9FnMzt7YO2BGe/IFEHlj95JUnC/5oujqreXkQGCUDQrLGKi8Bsu7
TirQjIIzs6cwJSDv+tObTWRpIXnvCRXZx1yfl1DLRA5ldd5uIkgmslg97pjHDpTERvZGno05eVHa
1uNKw59VUx/Cj0tE4ZvHSleiem6WpfwiU51wtmVtbI7CcjjymP2W7UNJnNKIKc6Eudv0xoUyPaMM
ozhx+Idcp9Yb2UtMcLcG/7S1tPFQawv0G8F9F2gke8t+vWA90hqg1r+kOWXswEAHWZt0Z9NOueFc
humMEQ9NkgXY8rfHbZzjRrbD+q2ay/0qIPVBzEhj3OsavMSr+aYAfg4RRQmbk3bjoi8gYe7ls/YQ
xHpDoj1QQvfJvcIu/exqqUSE9iRqUEmcPf1qerE5FrRS2zzy2twpOUD6mgeoJ1FWEczBvYut6pnv
d9BUveLmN5wpU9KfiFzE2C1uqruVgJVD07t4rI5DMc0ecyEgsrCTQ4AZP0hhOMp6LAmIb4uxmsxw
VXqG+Q8G8VAaVppLyEN/JyTC2PWzEwih8qoKhM7MOUmLJyOFjIFAJQr47h7cIvLIzErKu30Vojd+
CQKP8Xkuvwntk+f/Z14WywEnv6dsEWF+UKO3uEXDK+cD5JRUqnzVoArgyIrkmbcixY+Wv35IwCwV
mT8SnVqqFNjQtC+m+41wEfM4KFpSCZtTHA/ysppy3oZBYfUVo9bNObF0eVHCepTEEm9AZkVri2vD
s/DLMskBLQRP3kCo7YzePCaFPFjQA+xNkkN/ijzvBHbWy5WvA4NDQhGxZT22158v9R5xrfzYwcC0
2+Hjjrq1nIbWTYxfQ2nDHjWbcy+z3OISt9edeJHmSVYzOSTiB+FtOpVqJY6XaDXvShppveVSJQ3N
H6PurX51vS7JG3KxwIdHVQ4skRa8wRaXEHg+6aqvc3hTpf+0LTcbGrkgKLZzAFvHsgwBB+/M0gZl
CIdkxZVz7TMtqZHsOATNbcJ/RppoWuPU0Pg5I8D4/A0j6z+TDReKW+pC1gYDcFLF6BANF0nWVjDr
1tf1a6uOggkyYgBYarOo4QfXgIYTYky+925G6KFVaZS5ovA79H+KeSJ1vPwoANCjygvlpdT6U5JX
aSO/KbAVy+PM7XNJ31+mIxsZO7WWjoyHfdbdq+Hdcdf7xWo4Vqebx7uuhnjFqfwwkOUgSRa1lRUV
Kj84vpAsNbzGjeFiklcBZk7ws+a2KDDXvD6mDoaHVNoaXOaUYO5i25af5wDxnKPOngzN8X0zEf3e
Yz3pGx9Z/YNUGTn78FFJF7kkZXIuoWBApqlBAKT0BetfzkpNu3hPh7lySPZ0hQ3j0PRn9pWmRfar
oEhhyP3/wHq30Jf2sSXuRfKelY0TS8ie6P1hmm/jPjobFg2xmX1PmqBx3YRUhzLTiq5Wteaabv5A
yAIDKY0sDUXIdQzPHsyNo/uIVGxA4BMbjW4/cbrUtxFSfkKPbsnmrNJdO6qtxhwzr2Eaw0sjyvae
graG5THUmYtSDNvzmsehRI3IlGkw6liCvjtSEm6ElDwbHmCsGwFFY3UDQ2MnQuYeREyj0yUFyxgA
G0sUkBLOtrJK8t1aqoTWUtq1lUoQ+acz/FtCpfXbEXFOHUGbdosun5DY8/Oip4uZwdt0z/fv2Pcs
Dhjn4H0Xb0OujYa84ZjZ3SiPGyyAlIxatLEb4WrrPQuXtuaQHTmjsZkxlGcuLsqt5pdasm8spYOK
lQMBo//EYP7yai/6yWvn6N5mKl6M6rZ6+7s3gZP4ZN94cRowA08Rtlc+s6B5VQjveKTQ35b0KhGA
XU4QuirNlfcskmVnnzLUH9iq96l6TQaZxkNF2P6G57U644C9CULcQ8+F2e49vB4GFYTp4GHK7Qtx
IKsj+upfRe1vZ065lclsVVpMm5V2f5ITDjXaYkZpAlPqrd4VjwaBYgI4G4wwK1x4/zxVnAJj6+L3
lQDpP30HpDWbY1gTlD41TLgnOqjfb51x07ZZ4Oj7M4A8dYtrs/i9g95A2ZtWg3O7BW263kgSbVlr
SSvFDQJeRXuEvLDnQ+NWZ2tLyv7yGfwcs+XQI+UtFk+N9AnHVY9aZ1mCDuFqdvXYlbLTOPlhCHkO
JtnSVzhnzlFo6ddgxTDfZDEYzV16DthEKGSTMERM7BcY+7OyP6sE9zKzM22vjYYV4dZXgQXAUXh+
bGFNrW09DEXKtKgx3rFeEUHzHjq/ryal2fIak5XYKrsKIzWmDWzIasRcI1ERf11igNMeM2/fHoVQ
S+BXp8fBVx6gGhXOqLuTeMs656G+LUPgZy8SvQJWQqFYFR6dDCBCEVwjy84SO/Xx6fRDgcHpJMB/
TK+7krtQdFVpLfKmLTk0Wq7rp2+Oma/YFAaMlboSxJ/yF2DODrNe9M0KWmsejNGyxgVKYnHPKceK
QCxqzLlDBMlAJNTLDPhe49iNtnmFAoM1yx7J8UkJZhJViB/v588j8y5kTv5kGRx8r8JNpzJH6Ala
tI8VmAVsytCuAr21XgrjImflWvLnTPBsjYCwmTmyg0fvDw6xPnEefr5DNFLwn+ybgRQRl2eMShTc
KdPBPYD5MFdQRCIO0GxQ7CUfej2DYEexAVlpOJb16tqf3Ae+nVsfVNHTxCWSit07UdF4FKKHOtFT
8r9eAF1pzf/zhltFqqrWdqQs3qF+Pl/8w0fFIQ0VghG8iXh4+Gio03qjJms6zMhbmlyeZdAixuSu
GUJIJbgFmJJbBqSHtpjnhyAotoAXildrFkRUFr+WmU07+m0c9bEsPZoJ+qausVlUVsl8iTFJiDKc
b4gsU9cMPakSOdvhlcY8NXqgbgsVebHdxPBUXk/M/TbViNJOLG9RSVQBsV0MYnoBfP9sVmu3H1JZ
UT27GeWptxgLJ7LAiTdgbQ1aUNGT5/IKVg3rcCid6WyKxa4VtACRoVkSqu7ENMDVvSjTNjvGitls
hPcJjf0hARm5NIqVgcq0TiiIhcSEiGU5YOWuXNukhaAaCqVmxcqCEupL0HVlNnwwYiX2SgOMsBqq
zqlx/A55R5dUYhvtzCxYjxV5RigM1xhpSK5ro2G8vCEqmXBFRVpNReOTNfGwypez1QA+sQydnBfr
ALVOmUPtGYvZzzqS6r9GIkycpR1L7JtI51cD4Fyh2/mHGSxgmrOWpdezRTjFMLJ3h2/gHfvSmANr
J5C5JGQvcJybpuHXcsxcISiu9wN2r62cXE0f8z7FX+TIOVpHIkKSNI6HIyUR6jlSPop/2RQoftyN
vlekNIVQKzTn9DWqzibqH8dc+2dKp3vkkNkGNNKSYaIIrw8oE+9JL7MVFiJQ6mm6/Lisdbznv/c0
jV+Ay9D77cpbs6FYd3O+nniPHyelAD1mRVJZQ74eersAMXscyIxyplnPkCuhuHfVI80gzSTuO9ul
bYx5Pm8gftq5G6kaa/LTXpb50CCt3JcUQEej81eI8A1HGEDXh8TzFjJVv2nqPYJCPQWsGYhEtmZ2
BqocaJWVYj9gN0TFYnT5Z1A5KdOf8yIqEQyGG+uEF/09b3EkKmfwkFZSApV9K/A47ITHyHyA6tMl
/DpAJlHVSBbgoGo2Cbu0mQ3HQ6ZtR7QttdKGwPDYs3mD/ePclFhyvQH+7AVzrwUFo9sT5T1hLSz6
2OW8mxKXzSlzVlsTUy86zkhQ7yduCFKgZv5qKRfyd8/TEAoKicHzDM5qt/IerKtUtNxcA1BGEMss
FHrSqK5Lb6rXvEVxRUJWCyVP97cEYG3tnHAz8R71UHKtlCJeI3AS39LXWcw3CbjNZMs9Vj33VXgl
h9PyBNA/AdtL6wz3Fjd6OlOGVrWX30obHsGf+ZocXPgQBkk3godENhAkF2nyE/wWUOzzuqUFjX/W
i1blBOhKkd9z4Gw+DADyUBC9d9m4fC0254YrD/FcQnnpqCn2j+7e3EAcz8y6H2+FYGav3i4kuJki
tfU5DaHe6mrGl9ECyJz8K0z99wwKzCtsIcoK+9NZ7D4I+Fkje/69d/JQC0GrBSz2DjoVeBoQIwgA
ki36m1Do4dtrwzxKIv9Bn8zcg7tiJ1Ry1GKStWPhtBrYzfYW9EJxah5Weagbcu5LTCms1Y1IO3KL
fgqj4MCbcpzJEr51EzlkTVxmuI/v7qyoL9S1NcjgETL1Zffkib/3FpgFqvwUf+2QtdEbnEUbJG80
otmztOtFZvAT/apaSQVQMSzma+uc+ZabXV7MHhuxn9iSFSV7WwPwNVVnh+ne8hSEnIhEL9qRuIj8
lySqaMtbTdORlj/4HYMFrvN0SBR47hULTdqEwprWc8wHKmer6Ry4wlH3/4UhsXMleVB3lP7dSXyG
7PNd4qf4M6oMf4KbfrwvW9NgPYSZcdE2dN5XhtDv98lmsl8gToC7/UrnhF0F5T3F5N+ViTuWj13k
/6YjYXf7hPXInc0LfqZnFMTJuZqz+z8/7TaF4/fzFaTYO/duhUsa0UMKKA/v68xJvonrl+76zcqC
4KAsK814U0CMJKazqyjZlB4FbTKekBjDQOTOkgzvQ31LzjviwFZ6vKlPtI6xwuS1+Vkr2jD2mZbQ
6gQqqJlRSNPNDzTgHHFOqfQSVFalcqA1qDebQ8lqMipv0Ij10pJZNEEppI9Bt95GiW+tmiA1OUPj
2W4JI/ys2kmS2Qm4ALKqs6BF8aOxESIRz2yIGms5K0AyFMxx2Y8nR+x7W1xXHQNGgf3ryV0cY2E7
yhgoW/pOh5KcALCnjh9ylxJM9DlzXAkNtQvLKNysksQX9kAr9/aBMcz0mmPkIyMLXbYXshq/xSIu
otCNpdXeIu6RAL0Ov1Vq8CKDNtSiWVZvz7gFTDJMc4z7CvWBxxhjs6BCQTVtzty1TS5irkp3E59A
h2whdJjCHemR2ALLjuh+GTEoWpX7Lz8Zbx5zL/TZPOMSHaSsbYWFMeHudodEOdrrD+FFCZpfGXzh
W+tIEZwjAP4ai7NSBKFusa/Jce3fYD8u6kijXr4op00LF7WJAMxCL5euDd4PUwpw4JgQJ0KC0+ik
FZAYFaZJi9LhK0KdhrnULdyZo3xVjarQ2CXdL2NWr8CuaeO9GouvvuIrFXzLKw7HbxxsZtJwG7Zc
OOEpVbyBluP1b4ixpFXVzh4diYG46bOrJH0Y8JZ3fTIflPB4+zDQunyBnkQ2tgy25enYGva8tLDg
L7GfIJ93wBFji1pEkasbGcB5bWBiGfNBJ/jo9k3sC5foA/3FfF489J/2KAwfDphnHMOOYlzmKqRC
7Jb42J8YfiYpejdY87Jq6hv+DtN2Trr2QsZzJzzx/czM3gWRqdzof06IwrhA3EWUfAeZUWXuEEmE
HvZXvknxf8ipvxJxNzN5KHP8XMICPrbK+CbFXjz5JKwg58WXI5R+A6mKJDA6kS2bj0LPv49RsFb0
UVLSMdvme9mPxbFskcAnyRMOFchlBW1oATtvY+xGR8hsRod3UpnDsYWCf6vKJYzxvcwoO89qLmT6
r7bJTdjMWblk40eVyl+zdu++fwu4/PjrHHKkGbCEqtUcODob7S9/1rwaEP3o/NacNIw2HA8YZN5v
spIy7beHVB2QvCwohBus4O5Viz6dBxD71c0nv6ld96P+mIr0FTunJirX11DnAvbR06nxPGti/S1j
ksRBtHNCqCLwFE0ygczbiwbYtybBXcLInBMsTfXN/EvfNnwBz5i8Wa8MJ5nEDsov2HCdZEb1SbDz
sx3PbSVSQblWEuLid9RLxoqdyGp5ii2dxmPDr4Vo6sivt1dShmjixLrF6qWb1/NUgdXkyq4m6oqb
89v8rfH85Fi9dRomKPW2hMeE77l/Bb78F3+zgMoqxrEc/MTsncJz0GnHno2dfy1dDLNo6SU62Kv0
P98BISXLrCsvCajDvkh7NZy8d5y/n3g9hTIfIIJt/cKDUo1ayP+Ry3kOwNrZ3JB9DlNJbHNxcCHZ
nqUTEndthJfLAvxGJMPDqeAvU8na/GiwP/rw1TU4F13AfQhvmOfPisatt58DMRUHcJY4XZsiwbJs
7AZH4atsVXHoedgoU3SXpboBcpxErAgeRCHrAiCStbcRPeZh8qBUYeyzd5ELDkkVk5GhqkWUTbpx
66VnVMNnZA9cPmfCz/EtQU3KyJqHv+SKePZ0Opy4zALr0KAYXb5FI6zFtda92hIXIEiPWxSypK9a
tEWtue7/wpXT43lH5DqOraz7BxvRo/eyrqQBHk4nnWT0Vd9odeY7F7mY1U45LfFBr4xY7Um8VjbI
XerWUZQC5BbDQ42VSEhJqpafb1mqYjwty7YWqCC29JPaQPP0QFR0oFdCZER+lATV3j0xIZvrmLQf
21cmUTZ3ww7MgvMRoVXtenMXV54gYYSiHSiIzqywo7erDBctAcTBNhXd6zLTvmX6ovk6gZlBrKCT
G6IvlU4z7tOjOIoyfF4f7fdQa2uIbzvpQl3hJHwk77934MnYBRxwHlE01Vxu/GltPmLKaMXDFder
Q7pGBIIC1PVtpIkfAvupAfU4p1DMkbx888nZr+vr0dFBFsMjoSRABETzSLh7D1ViBAJAN8jA0QeW
3JnsAPVqNwLPhxY0Cvos+e3WyCQ/MOhucJ56ebvJtIX1/PLtEv6nOXIp36B5J9DyDaIOnkmF+Q/0
dXvLlYc/0aBJS5VMxhTTjvr/zoXSm9G07XF1pUQIWa2coFQqV7IqMkCojrPtaWdygPYW1iWa7+BT
veQCiy7+NdgnE6rCh8XSSso3xnaaBgPb5nALBxhCT3+ZpWKyoInStPTjz0PJKLjXDnrQD5PQIY8C
H0Zy8lL70WAlRKzCYJ2q5QlIc4gCxX5QlAgw8yWMQMqwfSHwRwqn21DbM/8n6vVTqIX6W6UpYEF9
JYGpKCdYBUUy4CcC4IBX9ARuh947KFrBKQXJojjuv4YYx3J4n+xeS/GeBof3V10vr/DkIIKqZalG
/6qJnw02J9mYbKLohMV6d0yZmh3My5W6Yty1rIQRnv070nxkwNC1Dstzym7LjI871F2ho37NdkN3
QYilU01+IMCOPGCIcE9U+0pnaKewxextDoigw4DHyJC+UI1meMWm8FJkIoB6Ozek2Mhq8aaHHCbp
FshrqmeUNsLWIiexWVgDEePzIhtRvrRx6Cam5nYQCwmReT5dYzIOQnL9y+KFsaxTeJ3mP+EWG+HT
jp2aDNEutpqmabHLWx+evhAZeDIn+qGRLlwSFyIwT8Gr/O8hIa1WbxcDFOeKH/dcqvLmYTS3nCCJ
sBgRzfa2x3E1eEmKhpuAN5sEcY4jTSv1QxXrPdoh5pkWIRYblf/9/EUooZ1Q4i7yHI/I0vFZwxjO
zMLEm7nVZ0PKxK2onraAn38xsPufFHlxoOBxVegY9j4oYkyV0kgQcgkITT/LCe+TJZfyyX8Vv/nE
bTVRdXoIs2FF36fTWFmXX8tBOqyiN2sSuk/hct7jyfxKFsWDijWLXVhRNaIbrP0XKBDs08MYpJ7/
vxh8CqVVDnA9YSDjyuev2c/jTv6AdHr/y7aFZ53pYn3uD2mC5QWLBfvgPHjGAodZSl/1hqsfd/7T
myYsKlwZ4EZcMM4LBZhBNduMsjQjcVGP6TstYEmN2vFzq9ZhhPtyDz4w1Sf/e3awpz4NYGSNiA09
g/cya4LL4JnugxD7F/UbQ0etDIbvRddewSPbQCNwBt9hOruZxDOU5gOHZsKLwUUq/zXN9Q8fcBcr
kMZ/QtlyWx7HFzUhq0a+/17eKz4HvYtW6DdLJFGpkCYZX4tcJ+zoUpq83DGkr8fn5gsA4Zk8Cxeu
7trXrP2A1QFPoqmGOjnRXGBM6Ukm5jX3Ry9MMOzyHxraps9ls9gZ7hQcuVp49rPL/t5DWFTi7iQQ
H3ke17ABeeriAbXS+CXNwJIqmBskIc0rfz3sFz4xtotxvD6HGFFaB3ngGvIAKCFy5KoCrWfpMJ1E
R5fgLSrNkXq/MtFSHetSku1xo6TzjVmZYy/6r1n5JLI02Yslo0iQcw2fnMJaGklF5vdtW0RXFD5z
LP1anYwpW/ufnqaKgt0tYq0/kHaQjNlDNU6z/hSb2qpq7vqk26enXIKRmb/71wdXdQ2goiJS4r/u
T7xZeTwaCWbAUnboB7+64dmf+5gdzQb6CIEK9BXGgPpUqMQfT26IlWUSvi2ChmnTwhRJKQ5it/Ri
fPbDjok1IJg5fcxXimPPEj5a5pWS6QgrNSoKOOEU5aTbdxJFp3TiftVR9XF/sgPXq/KiwqpcW7H9
CM2hyfDZTlf1Mk/kXfB1J7mVbKA8WOlqIftI0xZaRcepvpX9Wu4DIYXuQf1n4DObLJDzuZ88q+Zd
q3OEPoVr1vDBlPs1ZwbBYmgEOm18zHCwQrdN36kCSbqpQCdPvQxPRzBXJYL9MZc8B6133x29d9oP
o7W828NCaAy9+uX6zuI8wSazBMtgypfFbhmtrgM0XT3/QDOrHH95weFEx8hciPuulcRxcRSc8yzL
6gZ7GqfyS2sgUs4W61LcUCl+ZI/STQXCtUhURzC0Sd2u5PUFn1TvM8fQ/W6B0jhC9cqnLeWJT9gh
y+6EyehwUYFUOsrtdKxm0nfPXyXEhTju+j65gKih9owA2NDUhtzn0yVfwepa25P42gb6pW2uZqG/
15CZLcBh+V4NNnK+4ZCfAPSnpCkIRWssLPq75quFPlkewTh8JM3NX7NsbPIzOZN4Q+g66kmgRe+v
Wq4D8KQadK2n6bFyu9DBTYKCp6gUBTIxRr6coMi7gGzV/bOfP7QpWa3/q5S7N7fASHEivHUSNDOB
JokfIM59qQziNGoaXrc6HQZEcnRDQ1Us28CPdBZZh483mc1UwnCP6KwZV+XLdyzNZMTWHNXVdRLc
b2ilZSEaUgto5qeDeggWhftwBqVDVZ7y9nRjwV8tCawj7r1GZZ+mHQZYxshsQumcov15de6lcC2d
tJArqbj3/5KlgPfpKzx9SlLdUieOWK3J1KA8hRb0tZdDU7WAxb5NbqPRKLzMxC2VDy6piN3HpLy0
Qd+fiwWmQiPAhjWMqg8l/ufVEUAIx02HW1hGQvPNIdL3U7Ye+OvY8f+8W3DMuB35soBPYYjaaAlq
mBnPZ3uP6DW6vVofa5pwNB7GGoowwkqkgB2fYFQQaq9ANZo+/jdaQb8k+8JzPGZ0q1dgg+Nw9MyY
4Q0rKTicyuZtlYaBOowZ6wyLcWBwyPT/7OP0YJp1uyjzGcdcfCnyAWN6d8E0z10jGauZXCsXPNsj
XswbdTy1Nbe7fvyUao3PRmzEB4Ns8m5xYIA35SZRo9qsjOHjtmLkAWrxucHyx8MVD5R2CRVHhB1B
QE3GdLhj+I8+jtrvZ1YhgkgahOsRRmvMBTOqMlkk+HccGpaotepuxzTW1llAzel4TrkJ26X4REw5
RxhR/DbUBSIHmtIhLM+NGnzozfEeIDmhdzf4XgpWEPP/TTeuTGJnB9AILDkrdojmyRsF9psMKCUG
vxuzH1zoKNyJpDj1lldi577CgsO/FonAwRzYzyZuquJHimOmBl7pqgtF75bdqBu2T5nLXpl6nBpr
n+4xsicvHkRQ9gzEoCSOjA4WnIrw94HEFtM7+1wMKsq0MtCqYp1+TKb9l47gCTKYtc6SH7hxk78d
e2Bejp3b/yxVbJgMKdJfnBuB/Q7E5xGJcKKcfNPtc69b+w1nlUNXDZwuDj0E8l9Lr731b9TztxVO
0uR7Y7whkJzyBbcEFYMmrSn/S4t6uV0cL+QKzzIQ9K1ptS5CwDOA2xGoBZ1hhGbsKMVCeRfL7Gya
DIlhkEzuQ5CVb8r3tOFERHpfN8nBHJsmkLEd38B6j/HJnVZ1YlSDebs2osjc4aJanPaN3sGTVUhv
H+3dPBOriPJ5WQJ4CLalfz6BxeFXAHWzZ3DcAXBYqDMC5v3iHE5fmQh138aGT+rH/vP9+KDn5bma
GNWNbmARgmsAUUO2ffwsaKUhPDxf7i23b4OR4xqNvV5HYPgLirN73ixvsEkoEnP+HhZNeFfrHLeb
0sV2tCP6m8k2q4WpsGzC7sP/ydVgN8uXKINAg0TSfor5JIRwkY88481RdhZCFxKpPMrm1LAJcQTM
MoJTnaOwun0ind+f2ULqN4vME4xgPNA41z9vkWWRcqS7kCWE6/BB0gzeBr8l8wzZvGdu+3umqeQ1
kFJgWYQv9rz6XIjWgoK6yAaSMEQwL8ql/X29IkmpnQXe6jMgApQAY3j2W6JeJbrFSKEtDWFQrziO
H7HOccfTGhndI/b6nyO0wyxAbQ2oZEkjLCYl4NcyZTDVubLPV5cr94laZ5y1WAeDDs3GJwyC7fKK
hdqaqE51js3QGG3z4sX0B5tHb2FDSyFvJlPCMKRlu49xbIreG+a0O3N3pPQRHwQoUW19g4tOVST2
2u7fJ1D2REXePyW5BZAIyYtcdivegbPQP4mK3UZI6/qwy3n9vTGQsdO4eXeQ/+HdUQactOVP8MfC
bLx1Y01ZyP2Lsz3yKHqH+SIPWfhm9pFsnIQHJGg0iOpCoIX/5TcTNPhr+barYvJbONYv6jxQ02NB
IRlojBzT2MwzBC8Tlf+3QRu7Z0zoA5c8+AXweO8BuHn/jK7TSLUXV50DE6LVpMq3G3Wg358evb56
jHP37cJTTJQVEUouHRq9i7X+GWIA0XJ4Mliyx16b1vkfpl7Sx8ujOuSrua1X+VWmiRHNfZgQr1x+
tpbmfYxN1Jp6cdxeQbxuW/WUrTIOMt156GWa4qQYTdvbXz1TKw5v78U4gXG9A5LxYpL67/aSiGRK
XIADmRxT9EWlK4BuUy7XaSFC0gunyBbhcPyDDbUhdouTFdF9pPSW9j7XjGLHEV51QFZ2/e4fQwTy
Bed/Xkw7kEUGFFQGeFH7avCaN8XdWQtFGc+EE5cG3WeA8auRQTI2j+xYICm1JGyLXpB0PGrPwMRN
Zy4qnTcpY4LLW01ryys4Qi4506TluNNfQQGGIuLIeYXfaJREijiFVhQU8KNg5DHM8MvkJsd4taGI
kQxCS3hEwn/Fwe3Ity9Xa1EB2bktDjwselTcGlpES0OfPhMGb8D37+eR8ffBX9XyR6umCg4FLfRL
OjzmW85JqBn7qB2hIpqr245xbPg/3R6lA/pN9tysQbEm4/IkO1LcDcgo5fY3QYnhW4/V6f24bDOt
sn/tHSEe/4pVp+Kic6I4eCN4GJO/zHWCWxjFL0utf/6kLtD78VQq7VM88M9DDTP+N6WHkvvyFVE2
vz2ivZyC/3+ViAVDvSjZCpmhny4271KqbVykBlDg2U2afd9L1QoSri7E3CouhLV8he9Yx5dwZ2NU
Qr2FXiisFkWhH1pADV8S7BQHUIUD6dNpFH11+UXNmzBdCpLfnFLvI2x+pBrRY2lCutas0rfOGhIV
Vkq+pBhwpSA2uRPajWbn6QkxVk6Egrb6w/Vq9YEUWuViDPqNsEsniF2DSmRNUKcEw+PBQXKX6rL6
5dp8vmJ7jDfETbQ/pjRjkciJsGrK0tdoMtGfikS5HOkIUohT6GuqYGEzY7dDe3rzgk0VrDtZlAlO
JjiIlBwMfyBRLedgbNWlcCkFFAQ4LK5/BnDjAJcunQBDod9ACO/r355MmufhcDsryS6HntOZMkaE
zG5neH23hCv+LAagpxPG3PJsGACPXw7bHL93cqzGKtSY7lTadlKaKdKMeLYr2xNZE8l/2a7nEuUQ
VtyXseQLdEH27aOUxlCOUQCyAgVz8Rm+x0ZSMGn+5dYG4coguIp7+3U/fyHhmZUzHXGrIIYQxaE7
CHFRLL+5uBPio0XcSnTanZLPbm+JRrdlGqLChmOGC6XHO/BWVA4NxJi1xFFDP0pjrRsV6IWuWnnA
CsSROwyEkP+AiN/c0QhOYhvCt91kTwIZFEDv2bt7YHnYGron/vtLJ9LX5a5B9l5+KvLGltA4tzVm
Jy94aOli4UNijw/oPlXC1ryDDez3IYNx/p+3/eEhrZG1G3S1vHcaX5/CbSJ14Ak2RTCiMEzjAVIv
g/uFbCDS8/wh/d60xCA8FFKQBTtkjEUspzC3W6INlHOKKQk4dcAlLRlpslIduIKMIw2NLeZq1Bpm
7OvMlkmALyzqIWFbbKPuz3OE/IPHjts6UyBiLg+TG0cYkWSiqGhJtV5PhrFQFh2AJcppbe0TTtbx
XHmtQK8M3m3FuVcFlEGPHguufzhtu6hXE1+Sh5tp+MN/UNwlh95Lmpxsw8Mr0uGucDEwO9r128ir
CMdnGXXw+G3yyyXEszq3r3ARjU7e9/dKBegVmEensx+Fkt4rqThzeWB4Q9JNvXNxXnkcbzKW3ptz
r+fdh/DD99Km1zdlmTE8IUATEHS+gIX9TauWZ61DyX6pS30aHz1fvsoNXMQPfvmPl8TPIGwV+oWU
jpD4L4BXSkxPg8T3Z7X18XVEpn+Q88SXoEzr1AN7osF7pS9Jby8mrPJaqzYy+r4eoTOUbzsXd3NZ
hpnSlWVIg/HTH6nHv/9KHSD+XHPN3UyUW/j5ZIK3kFFv+Clx/VIkrGzteJ+/yIwHyTFlYsJExbu+
U93PY1uhGNUfleg8jIpBcWwt4ubl37lkq82IGU8rCxt4HiJDs//bt5Dd+yK3crR0aEgY/QyI3EIJ
lF5nfshOVB2Kv1j0DazO59jvFca6ktVJUbTtJVwiwhVDB5L8bHtnFx/R/VZ1Zo5Cstv97PA7SFvU
qBJgwTkwHyXxYhKmzoHzuu2+pHXob0mjq20GC1cpFzR+drucIBGvuIrS2DH9925ubAamZabsQMKJ
iUslDRqUOoOcyqjjY3iVGjxbFZne1DZ39iC+8GxGoE+Ianr0Ueq1MGV8RIKHNP1E4/SvPQnzFAyL
++U1mKkpTUwqryeouqpT9VrRv4D6ozSX5mwtxe0KsOWakhpgLzVbiJ3uHK1+W173ieFhnUVaOJEL
ARS6RzUYw+fYsGnG5JpgLx9kOc/R1s38mGyTJ3lQ8qtf/soO6hlcIFSzWhMZGujTIoO24Ne4mVjX
iyPE25HMwKnW6l/78JguZ8VpozdsT4mwQKjl293H1geP7DU/zbhG9NGO3fZWLKNWW0TBQoDxQtWN
OHUEQeqIpWTw6oMqSyD755nySyvjT7II0ygkjQalME5O+6WGkXbCA+8jK/oJwRk0go6UQRLMoFhz
g6VCQAo8rIGkGltabl91AMoKYd1ohUP5d8WTC1dYSpNmJ6DgxszvaBrNm9X7byzwyCNldwtufKqY
2URLPtcDInftTuG94yASBP6HADycGWca5WeX5CtjmkNLHWlGIe+Js4UQeMwwjq7oIDv7MCrqNtHW
OcUzuMXNWtjdTIR68a/eWjIafL/TYU81VyiKYFO1bC/D2Y+uE1UQ8Umj3wTJAt/gd5rHEgxtA+lk
lSXtNDzEdeuobeoDD+3bqPGsKtfMXovwE4d5PcXgQc6xZcIXfkOhmUluulsSbkLhI1GgTCQyVppv
Mb57ubM+UTapHJ+ExOuqN8Q6Z2B5IOqz8r7/RpIZGNa4kj+vsh5vQOL6n3zrZEbLhEe80an6rxzi
pOCy89FZ+vWlIH2e07pyqdi/qJC+gY0+eVNdu7PvppetO72dM2LQ4gepyajebs59yd5oE4LntGhb
h8C8mQYML/b51I1vDHiL7RDz1V/f65D+rJuhUFwavoRP24O5u24C0qY8AjDzP3j3Jhogdkbpjfs+
m2zAARKZ/Wl4kr+LBan+4kkEMioRXiPvuNWKkvSq29+mkH08GRS4Hnk/RAcwXHqjCOSsC69JI/HJ
8tt6kOTw+3rLC/axZtebtbIyvzH8jVN5Wr85iwoC/RB0o5zDqQ9GUAPFg/51foghG3c2t20upPHb
w5HWyT7ZxoKveZiVXuMhsqe6nT/alJWw44jkAgIxW533El+00Dzl4L29aKyiYuSMwoSEW4xd/69W
NleFzXwv6LKBq+XFRJfmTSeWnhzJGWTtfwqfYfHi9W82IBqw1eydmW0rOXuoHJe/qFUHVDgXYJxR
lTuFPGtwAjBqMadYY2wuavX4kNj4WP/nOR/3+Bggo0zr7AMr0a3t+0EJxBqpwnncx1xX6Wue8bFc
EFY0VBwhGI1ucE1BYYjsk9MiHjovd9n1xPdsgaGvS7omUyI0SLxIShfYzDH3GDeff7HG3MEtAm8C
aDAxAT7iFcFsSYjEDii6CA/VAS1mbz6TMjd/gubwEw/cN2cS70aVP3FwQv0mNdsmOz7B2PdBa9d7
/+qEFUhhn1FjcaGXiQ+Jcjn68EURWasED3qw9ZOzZ5KrKnCHvkEkjThWmEudadjm4NhyKTr1P4vd
FuIloo05M5ZVrJiZdlEVWoM4thOi+UiAFVJwoILIR8ChPxkPthiJqv+0nZy41CPY+v5ktOmj5e/V
BW28lozJKd2Vj3QMaQqsP4QTEDOQOCpw1K35Kyn6fCIQ2ZWCH4YG6EJZsSIGhj0388S/xKoIjMlK
L5X6d4r9ouFZoySRH+6cfTGgsmdLuKRILyqxwL2dX2vIyLIj3GPGJF1UIZpvZNzvMPK3pajJEeAA
Of/SWGMgMcs6o+6khgsCiIwz/IW63p5Mf2PNCCecR5OzAQa0R6gd1FSaCcUBu7IWdQhTF0psS/Qv
snyWR1IvAmr+5drbEWnd/DSeEwzkR/f1z5I2ZDh2j6k5IuQBK1SY3dmSNvnfxKUcP7YP/osmJlfx
j7k/mcSbrV669CewksbgMrtHuc+fMHnWQ/iHVaqum9bSnZitL0f3ZNFwIk2L7uT0xVMWyy+z3iwR
v/LRvi4q1hBPEb5f+u4grifAYZKghHBwomQHbgdgsbn8pqGCZzeeti1xmNuuZC0aV1odOaZl8pLQ
JNYwG7prkxWx3iEnmfPiVvZuggPhblSdaZSEnjHt2vB69ZnvRmVVeYqgKe037EJAlIg5hGjAxrFo
qipcK8XBJmSVWDXxy7W1MW4GMUj1MgbxIycINH6j+6VY9oSWNanOHT4fb7aEaiZ92fqEQAmA1qZO
3uTbA4Hivqlvw6IoUOz8LnQdKp/WcpBc/ubEaQ3toLjAZ5tc/R2H26iqb7SaPZvWEj7SoPAcg+BV
AOi+hIpA0FaGKqUo2803fJw6xsFh/7IhXhNVFlskRvLRBPP7LlC+5fZqru1TVi7KTAFQVyCsf9f3
8LP43eON4luJZnV/0bS5nfJnjpX3LagBm0qzSfA28rXAcX0Q+ZO7VUwYSbeMogi0cFuf8g3OOm/z
81upsDL9wAvDEuEW16L4tfACsZ2AAJnACN1HvUUfcuS9MJgnn8VTxTpKYmDDCTkieumAmnNcUKYe
8OvCsttxOHqpBfvIzXNgeEHajr1JVjANwodd3MvQyHNwxA1p9ECLpF+mtL50xoRpqF1M8PxKMrJm
FLDNWYBjdo8tpdKf6aD4bMv85kgpQmIstMlfpNCc5ILeffwTmZ5MLsIA3o8kJP0wtkzIrrJlAgV4
+aZOHQEZ7UjQxjg4509ida8SMrUtfvxQMzd7i7yJmR3XL2J7CYKVBhhJV6yBB4vTiw40K2qqJ31X
9cvGd2/+qIiJp1OkRXYG8qChnb6OrL2R6bPeeBy1lAxsIo0X5+IafySn/ZBU+pl/pUDwi+DIAaOD
dNtjtQxb/A+/OJmJqsjiszCNDDur650JAuM4iGCPjE+Ha7JQPSaNXUXkPSUNxhBQNlUWbtp0IKLq
6KuM6Y5nqMGFxLTx/08SyE0/JAEG7GYNz+0UnZvQxlcNvGvdPKwNKPBkfF72z3D8c3J+72/+EjvG
DFs9cZ1SBd+9QMTvYw5FIkkPxAEacOcvyILT4QvTSl80AexFpTR0oWuWlB/lvEf/JMz+xdctT6Is
bj9r4L7etwNjfTILMe/vVEFYAGQRaj9R7ml5qE/AQz6YN8AsyKW7fEB2O9dxE8VVydZswkpOC9/I
ZrOx7ySe89fNfWCHD+Wuh/ITbFGBeYs46o84d0BuO3rfB3YvrNccecY70+798wseoObPlHYaYyqL
3StYCqzzDcZI3sAUWqVtvGlTLUv5DtoTMxO0o7EXodFcQFVIkE1CUPKvotWatGTAGbggwWUUU5iz
XrXAZOXmpgAAO3p7OY6FkNsqK2wohpP2MpvsIWizirWOV5Su1SQWwL5vPyIEyghz3wvCsefUknMo
2qieaU0XBN/Tszp6pP2e8bfgRAuOyl10f3q0dIoxVnsKSnWv4bLdDzZpLRu0Hp6q4hIzgM1Dns/n
B2MiUzzzQYIynHiqRKtO4WXVBWwecVCkaSOoglrBrRjJlAwp1aGlCBxplaN43flAAlPdPVYagkNE
LIbWRqH3Jfl6YNP2oQWM8gpBDVA04sNZXO+ko9tkPxU+Hfz9sXcIvOzfOkZWekulqnu8U/sICsUp
/xbZlMGa/Ju8r3jmfQTzv+Dvoc8MHTzDmBVn+guCMpazAxkQAdEFIaVhOVRTW5moYOEtOP8U2dKJ
nfx0HFBapB3/iawyJw0DgLKhxGb4TJLCww+hz/bQB1HKnn0KxGi0MzxqhSXc0Z+D1hPEr9ZMN3Tm
E2sGG12BD/M7vkE1b/t3C7hQMqs+g1BsuvhWFciN2UNLfy5Z3+1KDa769bubEGGNCGnaZJ7AeeNS
hYh8ibxROoJpKC7L+3UDaGn+1oljaCaTn+VL16erMsMwPrFKoWtJd+Ec0HzSYmJamxM1i48M92QK
/101Na0XIGseHvneKUH8rB8TaQK93kqp52clAd1N21RU2tS8R6vcX36kMZZpGPyLRatz/qBVJn2B
3IYuuNchCGx16oOoU9iGmHS9AeW6SNoTR+pNSa2KNajAjqqKjIdM4DGr2/Zni3Rq9fAfJER7n46p
jxncXyDG1ZVlO+6Gf8e8LoMY8V56489DLYFlNFTK697quVhzROIh33/J4rcERa93281MVk7f574n
St/uiPib95wCqsoq34v8+cAc0OeKA0akIYyOl0PClYmDAkVoZKV/IrUYW2GgfKY1IzP0szQuOhEB
cXX6ALiMFXhRa+f+gWHD5/sONk7Pdii9Iy5682JSnNbA8aMwX+xD8OkQNTjJ22+n/cMy10s1+lGo
ovrGPCzsIjmJIYPCuyXAPahbQ+pSu+ZtutO3eqD4FG2R7VGRFUeTzlrnSXsjQDEN+NRIT4jT2F9H
bV1P9itOzbK6vcULUiAaTRL5SS9Oc5m0IFQkusyS+1DDCcvu2IS3VcS/nG86c+oJyai6D4KoqTEV
InVNEYuU2xOpxLcShDLqJZwwTJTDBXQXDEBLjrLqmsp6BwnEMXG1/EzicQX0Smx55dlDwAltFOQh
zpTh0bif0Dsih9dY29l6Xg3Bp4WyjZXuYvYnenlK3XW0k4RS59aUYc5gGUqErBz9oO4Os+nhzhKZ
MWK0SYZhbY2e+N8dx8TcTMFsusAZW/rJt5pI4874x2luuxzZ4QACEVVvF93MK+hOziefafy47NHv
Au2C+NUQNOmrfePm0LU6cSjVD1eYr80PKB0QAGHbznD4NlEU/8tjHozAj3I8WA+Rn+ThdcPH9ykO
dig9hhqQ//1i8Yy7Ue8eX6jfuYEtM+kulUMnA1eEaHoeMXbthOa5GygIMT0NgMT8xcRJ3njh9ekX
BocKdjubD7TOQz4XQDo6PRCNZsLDK2NxkXzijgQwR9AuLpToVEA4fATONO2aitqUX+Ltqew3oacM
swLary4uG333QRnTyAs/Y2pc2lDwTB90VCTW5ESiHt7ihediUBsl4+gCzp0QxGQ0NTQICYdhqQzW
2e7d8nO+p2KL7WFB9QIJ3rt7byIvOHU/qVpDxwFEnpbodGqLdU6vkIp4mYhgDM2esqAHcUgX6wLe
mi5+TOdr0JCPqnaB8MWgJLX8LUM+R03rxzVPCt5xHp0IP5c7gTy/3XNSeTdfYcdcAQegZovyZLWa
P/8OUz/6TB1tEZXHG9zoQzXCDkVwx/leDpAaZv97IjGMDhs1zBcP1qpLHGu3R5IH8r1xAWKFvykY
MzGRSo7f3+RAcw0QHgPSfTyjdhHccVweIfg+z7fbeLsFThHzslsTySRtaEsBGm7Okc1LVj86qONb
/YIAXQ2l2JHO+yQR3lblrR92nyJ61KiC/tH8kZ/E+Www3a60xknQWf5j2gAFaAxswl9atgN5s8fI
AAtiK58PbD4O97I4rIQ/JeLPE9Yr+Wf4cz++4/TvgRsk6/4PnPGJ4THqpntcxadRZmlVEZ528FCi
76b1wOGlHVqaulig9iH7NE8hGOhfMHoGv4a6pdk4VogjqQiozlN5dJIwK6U3Tzc1Y2mh3JWXPzzl
oCZyR/2HgsCNpU4IAbSIYe2cbb8DlUeQLVQeyb/V87yiRltOXCGL75uOakt280Bn9fevuXADhtmr
MGs2kdkF9m6LUJnrmd+nj6OeAgqPS3HvDY3mkU1nFPI9SAlCr4atCIt+43rd2r/ytoxT8yVRFR7A
1kuO3JYkRjoz0OsYAbaZO+TIiCvSIy6Mwq39SC1+PDLfi6TdumkY48W8T63pnCDDk3iVW9wqA/B9
AQ6+3jfzwUET1MQBIhueVAN9EoXCEFAnD1yRkTm365nlbZyS6/fYCCpd06KAdRmuzmpUu07hh4rZ
tu0VzIrspiW+V+WNQLak5o3SbGzb0X+xrFxE2/O7eYg8QswGIF1r9Q0tDhteP+ADqxruK+hG0Xsi
EU4uoeTRbHARPr2ANdzmrg7NVfGgqz35A1w5wEzjVNDLplRoqJZTEUe7n5vjAkzT8d0TQpvH0HQw
TjgIQWR2V+A2hm0r12FNLawHGKefhLpXvwHcbvD+MQLUM/HdC6m0HEhxmsgAn3h1I0mf/ssoP8Lj
7S/Zufww9HrYUrnG3oRZkivxcdKmL3AtSYDDcC5Bm62FdGy5mlYPxaDUKu3sNbdQmVJMlTJcXYku
0Kmon5JeTGCOV5/6PWcyDXblr6I38Z9gVX47LbbIxn4CR6HmcxMK7+sh7KBhxikCQNU0i5GmDGmY
CTJ/VKmaD/5ojTGwMnKlZdo2v3XVYVR3ywKcan/MpT9ROj8mHn9EybKFmsQ4HixKb+wlXo3xWjE3
VLea6WRKrBVuWhi+RsK3CYC+OjOos/AY++h/SaIvfTb6JcJuWzg8sO/R8818ga12+uvGOgy/9aZN
cy/v4JB4dkVXf1ZJqHJ+o70abhmBZQr0IX4bK5UrmKzea0xhaHNFlIq00QjkU2xOsEUgMc1y6su9
Ktvsz0/rsuBEPMrikJEG0n/+qOr+KHU4u6U2IlpAOtMkmSyrJewxLCub4f7tOSFSoR46Fz3/I7Jt
340nQ0vFRGhddoMnwKnlJ1d2WT9fbXXn1WLPW5KoJcX91QwdxRMM8zg6tdPEf2TDSao9Lx8j1ZEP
7a6HFilxm+RIQToXbUwBtH1aHCqzqTAHoyZyfk0mKWYdHku70ZvnldvcgBx3PJrBqJHiI7x/SVdX
U/H0OotHJGT4erfshVFbXyL/bkaKmP9Q6xrOGrsaXOz5KlT/khvZ0RvLEI1K8A5I81TRqQNBv9aA
fhlI9EGsJzNZv/Di9gM6uiX1qEYMzvEO1irakdhu/dmA9xNt0Qo0haI890pov9NQjKDyDwOIQKGj
zWK2k6aEzO/qJfcK8dwSeAhOG6ayInt7ydP/HeOpjuI5n8bY+ahIjbbdn2vuETGJtlMwp49WQB7G
CStkV9k60rCVbXDR3Opqd7789o496Hw1mGkqz8SgSgHgqjxpklT3oplymII/Ghf+FU35N5bbT0/b
AEM0mDs0E13Q/e75erRROlCbx5k9l9a4WHdunQ1YBhTw8C7H7ShknGGwjpz5oBrcXCgfP8KRWEX0
RzU3qaVjSYuS1VhrKPrB+mPI37ot4WkykdvZdWc+jlFYqGPTzh8CWRObe9hFQTVUZSHJDcIH2VW7
EEOVgKx07WszAPXH31J8/VSJi6OysAay47sG3xzdZC/1fNCCMefifWk/xjcCzn3jk9x7v+DuwF16
UHGAdsJjTIJ6PUPtffZCSJISjQnQPHhAelmTFLuOCQrgifjLrz9r32QGgaG2Eu7jHK+rVKdxSqk2
pdEjXceMQtmqEP+UeE8DWMh33IjX/do5T9Sa/UYxj4sevoYDmBZ8yrXWVcojuU0X5aZ0ZG7syzM8
BwlmfdHWkT+W7kmbBh8qA3Pq5SMc88zh7cQ8sTkOHwTIG/dVShBIQaNCyOwywMVjy+C2LU+pWNOz
OlCb44n2Xvojm9Ywg4JpXrXSWnnG0YANPkZjOsYSlks+VzWtpQV7VrBMFIVnYsZYzxLIXYPC4LT7
lhTLYeBy9zF7+XkngPgGwGFrhfygRWvKrPX9p5cVMfmEz31C9qBEkD+ZHjfV8n1Iami29MT4YUY0
B3bF4qBUiojWcduzTo5c8y0scG7VFQk/sHJiXkvXD/JYHsxzemiF7fgTglmmY2kKBkk4dvgtVuev
6Qv3LyV9K6xS2Whyt8hvV5InMC/mzEuVwD8ht6hRxR1iqTTS5e/vl5AP2QQsQFijM8slUJ/cQVT9
FckIlmWRp3nMdtWOTlqhresLtFQ3i7R6yGkNX0JXOJ6MGGcpUqatXxezING5vPJWsQLOAQqCHpCS
2BhQibkT1/yuDLq/Q6PScocD4UP6lWbb7I2cJPHsVbo6ON/VAIjl7NPYOmqCxUmQ9n8mZUr6Esoz
r2f3R0UPPUmSPqf35eLiqU25LFr7UQHK4OADamQcEzmRgZLZluO5amE6r9ymXldI0d1TjBSE8Oi0
26iPkKHHz/Dc/ntZfUrrI2s0Os5h+eDTaUEN8Q0opJJQ3FKCg4GfVsh0NIuOnLdFZ4oxgDXLZXhc
k5n7oM8O/6f+FpnbsQLJ6az5x4TU6fDymjiRN8zVjim6B/YNSXpNKMyuhJiE5rgpV8yZnvnIulBE
CFynBwg6EzJs3h3BOMafiunjsUu2wpSUx36wOlbHm456BLaT8a/hqgkIseuU/oUbiymzTgqMW22u
5aUkTCU/ARXJTwJC9DzoLJgRXI/1E/k81r87zkH19lNph0pWiRe4J34e5PiE1ogAsigv7M4vo7uW
QKor1hI27eETrl3FUv15qsZCKQ1/rQ1oLhFwPJtdQUKEjuWXmm7dMf1c1OnTRb4jMLUYh5XkSPeJ
VakmhqA2fOSKnLaQ1eWE8zWuvnMkisS+ftyN/kp9DURbhTuWIlJiZhIDyn1GRFMw33FXXxF3qOEV
2+VTM8EzJFpUuTJkM3WuKz9Wb89tcqxvune8xBnrtqi7QPH/ov5CPhtH1AHjJoT27QkvRJ1R5Mlc
lTYF5ZhcU1HOeoegOx/E8mwfhS+rvtR/pT2Ji5V4IDUvtCr3Oj+LDZaK23wa5L/ZjEFxAyfT1S7o
xtFbDu57zftz//2hZeUNCeCR1NpFrhnct9pbd1ciFSaPKNbgGnxvu/hSjGwU9KbRJKmmSwxwmeTE
8iwqcrf/pqjuYcXEEQKZP+KszXcTDAGXeY3gZw4BXS3u2EaYkbg95ikk94RzwzUyrkysIOeTm8qF
R4ICe+O2ppl/JC7Gqbvf
`pragma protect end_protected
