// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
n6kY6QN4Vnwb41OiHBxZmCBH1XFFZQgrCGY/p4lADFOmqft7mYNOoJvViGz8GUzkOt4QkbcxEIvz
KmImRR2drtCF3MOwqqTZ7KiMfjaxzDMs3yZflnCQlUOKjyv6iyAlUDlcBvuzrpmr2PA14v3UeQ3z
geV4oiNMXzhY9E1soCWbDGM0Uyux0Zh1pf3PQtOGsUOQjnHksVQVxB/JqhJNTS/sA1RcwCYom+ue
PDoZmYSQOuFhnuUeypWJjS+txa5sZUagu+EqaxpHZG5//WH/CYxEm3BMxSVOUmrMQXpNyrUkcWJg
0/XmvugjPaGzeehlZakWp1QmfXupmNyAH0pMpw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
wKnbF5xj/xysB/ujoQx0jrWS3xtpLQM0G8NuJZt28wl64sVkDPz2qAdBMALCee1VotZWgHf6ojgu
bgf3GRTrbmIr+VnoYF5b1SNftf3+nI+EvRjH071VqUpN2cwDY63i1XW7BLaUNLA1TY2soJcyD5SR
zBjMhXilxAzCQKM05jcyu6UyZx+eEVBR5n+7PXURFo4ycDi3QRvsoa4H14TCnLgfka/bLUH32WA1
bXxVw/0zrg5OLZsX4najeWCMtCbNEJiTRBR/0rCrg+bNmmB9dDYYQsoAuxDuYknGM3FnyDHhkymp
qXPpZoX2CbjJvrxJjmciIeis/rPOjp1f7+l9wwl0CW6b1uu05jnTYPzlCUJSCblYxbKXMt95321D
xIccSV9RrRIw6LPMwNravVoCZfFTEbO6mOt1TmWUZXHIYIMEJb8eHJYXkf2786WxR8vwmCxsEEq4
BX2YR+lrc5NKxw2rcaWvHB5IvXbksfhV52Y5br217OlKP2qSotFtPxPYVP4CBvgrTj0BeinT8nrb
cB3ow7dJcd9cLernpV4d27S9IE7s+SMb/KjxAiO0mGSndQHt2J+nC8n1OfN0GyaVQElfGd4uh/Cz
DJNhLj/g6FArVX/jn+izk49kETnW+QHpsIB6hffE6NevsnAozn9PVpPqe2nQ9ekVRJH6HQlY4PSB
FPzQVxpREUfWTBwBF+7q2NOyxq83PNKKdScchyeR2ig4LqMZaUwrxssZcSYAgnfJLwRnvSj0a6/Z
gViYG7K39+wWGT5zrT7IlUfDkj1vLZ85HzkmPVCXmkavz1UHYoGA6cpxPPURDhFV6hOsNtLCl+uV
R2tUxhKAVA44inOYtZHLkk3+M4XHJVPIVzXNI3+zuTfNdol/KxvQ/PmD+LzW45BuXCIIkU2ZKMit
gGiUqZbMg0a1lyWmipJh5aeEuyK2dnmFzZ7V174HAUn5Q9sjChtHtGbHe/x2PlXzNv8hZACY6Wos
+/h9mITcZndBfNnjHKzjDb17ehsX1ZKEavGBECRAVXiJVB+pFpxKXfM546uXfHUEPgJ2R0wgS80n
VbRjLUm9CHFMG04EkL87zyV+ISs6ytoJ+q2y6wR1QP5/pGHvYjZkwTC05sFJhBF7u2zLB1O1+Gz7
caBZmI10WKASf5x2zrD6owpiluvVj4jmCPhYeuYSDjMwuS4Q8Abwsdy6I9BUSu5Zd94HsC+bGJKL
ac8e5OB2wtOqu+86NMI/tXEGM4MLU9N2oq+a+p0T8jsSUyoU9kCS11MmDnd2kilSe+WpTItK44mQ
FdPOfSCoVFIha++jDuDRGsjfoxBLjS+CRyk1xQbuxEa+/nJr2HTCC/Rvh7CVnOz088RMQS9YIsJo
ltJ1y6s3+WqKvzMeFDxyb0zHviQegp1TKbFhKHcZq+PABRdMEmVjiPNzTC/s9TZKwhCf2t5/HAmY
gpIWv5RuD6NmE3JvhW353juYR7Obssyw7w5M0hN/N/7lA1dWFFkn1BTGEMS2U9WH7aoRa8SYIKFK
2iv6i5t68ehc6O5HZwGZF6PY5QHy9K3bGNlvk3tM6Tx8orIwH3IOBP2mWFSUZUcye/qYT3uAkW3X
ihpkbGdu2WHNDdw5EkMfz1AKuKmQTIBvyHWUiJ0Rany52J/TSRJuV1c7Gtjwl19GJ2189NyFq/3t
zRrsI0f6VK9mBM4pVbx1VTmiZmppF1fG5vFlNYWdAUoM1l3WqXT+AvHZAlFt9WSz1V8aZcTUxhW3
u+qcLWvEAi5MFQSOH7pQwVNllUphkpjZzM9HQ2kPj5Lh0TLb/99s6bhTKKBdjkNTONU72B6Q0Cc/
UQKD4kYBmMCpsczWEzz/xfk8eS5KaZiyTCBk7vpHRvcd8JKXxnxG7h6O9u3TSvYrkdnyKUsdiIaq
rBiGl0TqWbsHuP8TK+X4xZEdPg7skYBbV+XGWvOfHacKbXBGAx1LNqAx1x694U+mRupufFjyTtUC
aA+Uc4etyyzVZsxS/0xwPaPFkV+o1oZqsVYH3gt7d6SRcx5EDijFcou1+cYZitp/Idjr28DIVWlG
a878ObifRX4iHiu9GoGwaIzszC72gYq+KT65u/EPPUJsGL6rWSI59vgjhv/zA4Ft68GdHu+3RcYk
C1R79oL1PwOnp8xMr4JPTSg3sWkO8DZYg66x0WTMIdPWYJEfnfVlLaH0AYe9w6jJPI42tfdxbf+c
9WBK+Qj6tBZZFPIrZ/4yCwdWJsAd6E5fQLYVjpVD0aqa1yWoJwuq4lukNKpRKC8MIPIMMPpfU39i
HgqZMSjn0Tq35J6FDzr6d2Q44zJQkgvPT2EZ70mw+tYEURU/yw0aofuvoKBhkp9x4khjC2LmrpJ2
8clFXIUQZCSEqJu5VbBR2EPH0CsGfEXiVV3vaZzhtKtGKdb8PV61gy9bmoFgBbsoxVviLpxGwwK9
xbdTFegar/TsnybH6WiEf+XJx4dT7SC2w9+Q9OsLV+BnnPFjb7+KSnc/mOEmHxPCUJnaT/Ekt+Y9
cM0ToAh7G2P5nQRDd0fVaEQisPZOPkJqqaGN2R61Vy1ReSBakHVLKhQV04HvWN/CgY0LABecGOHJ
AbawkLN4s3SVJdj2N+vwHVkf+Hrc5uJANEOI44jmBw2xgCpxEBvWor9rYiJSKxJ2CEsML+EWX2lS
cZ9O3qMzdkurEpITHonKNkr2ikRtTj7jE3qv0mRMWA/gejVICzK3rHswofu7ttmicygmTSaIVtYd
5ONZVGZODaI0+xkr/tKKqyzBhUTqBEFSaDNfv7uMoGB9OtiowfcFXcwN3NrwKw6G6lMsByCJsVkH
iHzKoXcylO/RVf5VqQniWqq0aqgHZzNxxZ1ne3eJJdh0U5jCuHA8cGeyy9m00+glOLEt0xg0erOr
SmJTDilv3Zam+9VkjazLm4bk2gWyp2PSZTlPWgOn/6FeVmheQS75AriuugCww1n9TH/uLvhRgFdI
hMwLykAhSYPdl+JCoyY38yvQ0THTLFti+iXxiW+vjVLf/6TOO7mx3aZMfrqpk3Gjmemeu9Z67z6D
PmfVcTFp6k9QgUf8ihuv1EkF+ikpIR4bA1yL/7UAVQz8EeyVM4pNdiOOM8FI1YRF0dVf9YFRZyJI
Qu/dOxR9z9REoQmnrAVNx3y+VpG5L1G+b82VLeYL4EBaYUnNKCgtMDhpf5GX/S84vLkHrjohefSb
BCp2CL3vO3THoht2eU0OHI9N1snzW6BkvUVIG5UI+NZVBLhaqCbLM2ranKS1DRbX6vFySqJPh2R8
TDhN7emgziPFJKNvElS//T79gYS4RtRstoSVOSEVX1Z5BXCczJYqGdI07nv+SBzPhm2ixBUlNdQ+
RmeTUfHCoC2mfZk2LGRDJDaoOZaEduE0UFG+FA6d1fGl48crTdxfKvW1W/w3+1+Y0QKXubGxuJ/n
/2J5vrw9L0qQyo3WoeZITvrGSpLa2Pr43lI+cAWcqaIZ9DhAiA8iZ9iVwREbPMwh4YQK85uLNJwr
qZmgMfsCe3PHuq7GQ0kusRPuObytuMXRMSd7L+6JT+vCscbwhiLzcaw2QvXYm6dsriYTbs9CXbMS
7tr8D1JhZPC2cSv5fSm71juPWCfGFaoacLoDViw3XNOKMEMZmHDzEIqirc+6nPlcTRcjna+CIQfm
o4ra/r3ml09Bcad+omEP4lMxtJ1efn1PpY0nHZ8to2zc6GW5/cTrxYPqh2M+jH7OXUlH9fRbQIpo
gHuV+kag0PnRsuSNEjSgnIOW8Fjn17Yr0JJq9sjpSrhVVCFS88/+E8GWEqLjfCXQgCrK2XpG2fRY
XyBlAmUESKHZH8jowBIqQO5D2WlJtpIgE/RqM+f+6lZsbIVZ9LQf9H++h+as/umYBL1n0HboGYqn
5dJHp8Vkdo4M2Gd85hBTVDhQdQMzGoG0C90nhXghG+/uljwCFGSZ+2AFmI2VL5AHem353kzwNqvO
BkKab4nyXXQ9zSpl39FBwvSqwwE1AkQlVbMOG8TEIpovjeMaxxBBrLtJRX7Ahy+suv5GABw58JwC
QFUWTarJhBKJvUzf2KAyh2aBlvUs11V5/NL5WGc0TQnW5nVMWgYsQ9Y5+EtTNYjkPwYNf8BL+2XD
mnn93ajV6cbMBFvX/mJm0bM9AktSu2pcHAN0EnBmb0pQe+kDBpD2IGbm4v/mvh0RGaqTcDAPDH6i
Ae3VtDNPfZ64DLOkb7NcQlU3OKmO/4VWbC8GmRN4ekJes1pOsCEIg2DrE288u5Pxp/6EH+1Djg6O
Gc5PlSuPm+L9Zdr0iUBGeerWOdwjra0qf4U42pcbHUNT6hXbJG1BkL9K3ED9ATavim4c10tZg+DO
jAwyvVTKg4X4GgZqeK3EGl8rRl0JSkSjsRPkYyV0lQD9bAd8+WYhKBTLvR1AMJTmejS1CHiHv+9J
uNeOff9WrJOnnwp+ybmx45ohkl1KE8Fd4H6/TUQ9XtACL+3aOYeWXLfPiraPQJ8udKldpV0Qz4R3
C8ogRlE1K8QFQRQBX4asOUdWgtnYILNk+17sOJ3rAiiLYbCesJ3p+7ykyKZlIRWXvm6qnPgn+JOV
zODb/ipqH7+H7is/VLH4Mxdfa1DAMP88g/N/DZ5mZsQjwlozEM7dcQyufXz3Ky1o5NkntaQFc2tF
hn5eFm2rDqem0b3Au0DCWqT8cpAlYRbyPyFBd87FIPbvHUFMaWn83w5yePypB6nDCT4UlB0rufAr
5RzydW2mWBHnZM0ZX+4u6BwTkl80YpDYUOwRcRe3wVy/RPA4MXF4xG1brgXBvta+tYHgOBvs6VDB
uXKQfQuw9CUlAXHYvtnQVjh9GsXAy3MP/GzzaWq+zqPT6YS9jATO+WT2Z/t9j/PF3By+4VyVRVLP
/0aIj/x2iMwMP7ZxyE5CtRziM4HKqtIX+A+0KJ7d2sP3NK3vZnf2/dluCx6LoscXN+wes1uR316m
tnX/OoRkym0St01dMS9FBnt3rZ2i3/3J7rnuK5y+XRbkTUqRB6GEMkX4sJbyjHDm7fYISexPQSx4
d5tMP3oMrC3zE1rdn7tbK+qR5gMIxECf7EI7N1z+oGGe+yaqV4UGjRn17Z+R6tIihgmiwgCfvpp6
CK48CS2OJhl0bkIv5e9d6q1Urx4OsYXcdDwOlVn/UJjI/T0QkCo0L63+OQDkwsweZglIED/KKp9L
IIDyqQ0IsERee52v6LUByGnZ99HCmi3G2feo2Q86w8GqJSHGriCEe4nnmXDZPNUT7dA+qyUaxFKd
sss4uQmouIZU4J7r1iQ85Bn/WH+8oQlw0Uyv6BCNfOet0OUFtajpvVYHmYUqgGhhJrnO/+V48ZoS
ITGaa/BQOWGrjYTQgUQeaTJG1L86k0/QdaiBk8h46EH8eCFK/rhGPtwhnAkoqGgAkrA0qKo/YCn0
mu8yoSYbPDZ1uDCUiW1/k4Z5Dy74C1sLVzXshNX9FCX6qZ+9Y0tPz7KVLr0Vcuyy1HHttIHaoBiP
1R/BPz5Ky6VG/QmTaVVR+ul3DXXyrb9xF5hOnI0Fklf5m2+aviZ3XmodFhB+Swxs/1etdZxyqOt3
DTbVbC0zvUhDPXx3LurdTeOdU8Z2nt+FTwZAYCT2fqnallfqj75ZMV/yY5UHPQnFPbIF+TwKmPxv
zXwdaN2CxT3OiSgAXy8jN6CIkGgjq0qiFntTztm6NhqBoO7ktDWpZiqmDW+sMr2Ltlay6L21JL+v
MMH4qPprThg5rl1Uj+Fo9M8pGeGX5qplaWQ/wpw9HMJvsYs+fjawRzbd8guzKkg6KZPwCOR4NcSs
mQQnOrCR855HJh7MZS6MXO0v6+wXvkUXePs7xsPLRyZKOzSr7sSfSFWrVQTw/RajiKSUMKyVScO2
oTp+G+UMYc7kS13AGgt9uv1zsM/wQZX5QBN6MD7LtPrIvfiwZ0R1Y3Vq/rgt967ZqWyL9yFQgV7r
8pD4mb9FAUYO5McE6oFynyVMG9TETWM2fiR/20FAMSu7O6zrT6GIAn/4wSKct1hONBGQy1YTg/W4
DX5cLBDiF06dqLudrHQgNoFQN3f9cwhD+2bf41/6K21A7axCzpcJhGXyqafVFdNWC6AAebSBXo+K
a/ewm6ID4/YuLsRr5KY16laKifsTfAlNawbX5gelHPhmTToyU2F9zKY8UmnkCUWjxHKpyfz+ABQ7
nF1LXqoWAnb5wI/uE07X3qPF0sQ2k6C1XFFo00kGof5ztyev8+KLEukkdNQsRD8uchyG3ybpHaTq
QVACMqHgv6626UWAwxiizZwFRTPyN0o3p5P412q2T5rhwKlXVaXXLyRrnxrrtLohi2Eei4BPL2Vi
inQ2M3lxY3KvbMpC/IrRTJUtG6dJKN2Y2RoEQhQBd0BVTB7TMQHVFNMXAzDrUDKgfLechqf7GBdN
EMzHvVenLqqtkVf5CIKdzfDJmq9UXZgWt0po7MFjhVxfMHESqtnIUK6d4aEaiQQrGVeGxHekdinn
50ll6MDW1y8kClC4evBgX34fJ9VhzfC7IQX0N+r5HPgiZxTtXTBWIr88Sni3E0PXbhWYKOIGAqhP
ksRhOM4S6a1zSeNtxwh1/F/UdGlxZBdjzk9xjYthAB4rtJoOQZfLuh2WY3uKz73bq/iS0pi/KKHI
tOpBcET2pB2goUqwJPvyDm0CzT+tJHjVxTbQ6QTMa3sYgu2NlbLTYZtnZ6+ERyqraM2Gmj/garL3
NoV/WHSzwWgUfZC8nQwf8EPmTm5L6PsHaqyE5qM6G/KfAWK0S33HUO5z2DRKmBDSZJQPKw3fLiKs
iQh/U6WvyOsrTMAwAYv/CzvCLFVukSXEbmkZShkZQTaeu4N/tRa04HLoBUHZKFn46hE+nEchE8/g
BW7miHWlr9FG+XFB+y6QdJqLnFy9jYoFvoRS+dnQ9944/QcB6MbF1w/5//LdNE9N2wIpX8jlQxAy
nCV9nhjSXDQHFpaWgOR7uoTO6cVxgqh4uZJesVBSmsHroFiuy6uu07cxJalWnhwGMrthBcE/1GBL
SdfQnCntrJ0VISmkgYz7lOEmObphAugxrY2glYTknW9EWXCTiPht2N4IIZLxPLqtYdRVi/3B0jy6
xlGUDTegFyadswj2tPboGTkMYOiJT+dUcrb6ef4YMfoZVyj+zEOoIJsLy/dnMaQqzFj8FvNsEBNo
jYDDkeErx2hceqOINmiqU0ipNX7XdWjeXhRU17q16AjhX3BwElB5OfDjQTitsPi0Fq/Hgd5YFkbz
pGwJkG3CunoUaU3eXwKOR30XqQIz55jhK9D14uM6cV1UsKHmFFM4Zd0AVfAXMZ5tyu6C7gmSzPLK
qap2H4vnh0/KrvriDB+wUuEEfpEp3eOnvZV+NWKfFAg1mxO251Y5rez7SOUjfAuFmirhfghEJONr
oyVfJJR4GjyWGE8G99JR1ropfJstpjh4bwLPYpSWzK8xTFYcg4Y2I+sIYPkM0QWP8My26sjlBrw+
yH21Pe79XXWNZsq19oxP8SlpXWUzcBFfvgscZA5wcUJ+9KqHC7SiXLMbCTCXUG5/kFWsH4FlBzBB
IXgnrOGpslA9s1o+4Ux2FljYE6FyEII15hkMMbCmitogPQFIrh4Bz8HRFZiD4BqtuPkpdbxmNd49
70Iz7hF3pceZff5tfBq0o4Y81X2Ul40u/7UZOUBIRVUCTX8LJTwEnz341uUm7/gUAQgICgpilglZ
EGkjGSnGuLIDGhADU2wyJ1sP191cRANojziiqu82iq/mIjSY2MMRCDOy8Fiw6wcFdrBLoEO0Tpmn
Z4WwOp/9Afo2l4pVCvezhaELGai81Ea12RwGUz+sdTt3J87P/gIYxHlrs9dQhVWWvqqZlcmdBMZE
E9bAmr4VFp3easa5QXbgSTpek32Hb+CbYcRekgol7tS/P0uHmhyAaQNMFHPnHtUggLfbZMHVhIkc
tIsukzIWphl//4fjhGq7qWEve0Y5qdcaHO45PH2gB0f5DzBLbTAlO++fJBb6h2DeNpNyoc13gHMM
Qn62+KFlcegc2YLF9751BeQyESrd0E9g9Z40jaJs862tzkZNsh0aIN/xue0RBo9akdCkaL2gBtYb
IrzQVhnbH0TzaG7oSBPA1ovuhqMZHT8u3VrQU3Zm4DUcvrTUuEYgjbsPyRoeb/dX6ezk7HKp62IA
74b909XhK4FX27MsPy/pcndLVWd5mExJFGNtgPTOEi2UUrndYPQgmgh/aTtn+zRc1g8NAx6EMF73
hmUQ+OuFmV4F3KTTTr08cUvbVa+5FipkdKaBoBl7cVWhiZOmVBfpjbzkVGm+75aR+mvlCCDJEugP
hJIfd18oDUTQZzs5rkVQMrssYvoeaUUQFu8cu74EGaI56YMZ5beqb4WCPk2Fse2j9L7SqjqaqIyN
tN/01TEVLfXb1VZJHlkw9GjImJFGxbmCcEVSVEQsAMYbhMvuFiPV/rywX43iTgBMGVGJ86o9DCdQ
3KRzNv0AHFYxHuCxlQjfmVplA15A3MXAE8wFePo3SoVN+1cQbVsWNb7d7RjNsJElI4GZhPD2PpMk
SV1WRoF3KuexvVAFnK38WKoM+UwlPxVQqPC0lHTEXfBT9ZjQ2ACp94s/Mz/9b1ig/9HOUOq0LwRh
kIRhw//bx+x5WrzcGRi/y5UOV0ks1PMySNGNmckP3uF09LAwgsmfMTOVcFRKpnD2xuCG0mjgF0v9
/KZutJg32ZPC8NcgDk13b/dw+s6wGs/6G5vofCh9vqR5GevHBTTsl3P3pRBWgGVOczn1y+0Db+OJ
vGUp9SBLu/nQnSXSY8Hh/g0KpN25lhzk6jorWPLRnNjI8TI3BdE6ovao9s96T+OfEGJorteAU77P
OQafE2XnY7vm4W/212JqziI4Pdeeg7oRvvIPk1xZTd4/s9T+aZNP+wefKCvqVqzRVejBN35SW/fn
3Pl0IuspTiUAE9M/nfRM7Mm2UCTfdgiURZmSu4Hcb4B47TC8C0ypXy0M8vcwYw7zgGmAQyOUqUqu
Z6kdl1y8W3Hhx2fM8zjYFyp6ls4DlK/RiCQWtYouVaOqW2OmB5SM51Dl5OwQNQNnxXR+80RNKGYP
+SSFxB2p8TfM4nFfHYHxVxsczhqK0sESnPWxEEXz+oGx4Hb4dXCzL6+LHDu0+BtT2sCZUJ6kG9n9
r2usuWdZGFkWH2nYqgthjL0GCH7E47Bfc+h/Cbf/TFTQQ4g5rWawTWkJbVkpTooAGwq9tHrEM7/i
PYqnsCRN85i3+qvujDISGqsqDg9nAZOjrIbtoIa9sY5YwLEYqCdtEjk58hwrhLn/d6uRfywKhxVZ
2MkC+11iKXrsqkCLKdfDCMgiNFxV0YKgZpZ6t8YNV5WbOCSdcsBBXHD/Al+Gk0OUCXtB9cMMOGVP
KsIe7ASgO0njzg/YssHPIwQSaU7Z4qTosq4YSi3gyugzY+Ip83dKp5CKvD0tn2Wg3/5GLtmHxxo5
vMZsN8bp3p0TI4shqPkPrgyybZ3+4YaywgLtdrEf+PUIr06EUdFrWkU/BPJ7CyLulSNX5993EvCO
iU/jXWPXhLYx0e2wXtglHUs7NtbP+ie1OISdH5av/lIFcbuGDh43bQvqZY0jhAetatYh6lBjGU35
WILDFJM+gtiMERlIx3iZZ6ztZLSHzwmoNmIFm415vxvwQfikyl4Q4h2GDStC9+xDIAXoxNnuS22I
+jnOZWvOrDKE7t1+xxH/VUeb9r+E6Y7t8ybS99lQ0GJebehyU4MHSxCt0CkdCD2jn7yjdgUYAIRt
6Relm6Xpi7WxZlGDJ4JIfnN9nJFxo8WS+hTVbZE32ofDutONa3mEhO0e8oReT/0nsmefbMi6ah4m
lUmiKC8wgf7zpAfzMzgbh7jTnfpgjJeJFwYfS9BD1RBpPKV1wxEQFQYBIVMkXTZM4mRRo6BG7KQp
WW5uOKIbFvTvStUJ+UJMnPxz5Bb9A1dDxv8oXKLn6zUoSprzj1Gy7lFf2cjGpf+t1cjfvntcVrGn
oVtHyB55GLc0wGqaw3pExkT5SLo03ZW8yizIedDsYESE3Ab3MBd/mzStePiFOuFMaZSAVP+IQq5w
HqiR8tuO/Tw/6GwMofsj/baDphShIvv3j/OnJrn/qiFVCqhNtUiekIPyvwc3sv7yPH0b19x744+D
ly0lsjYw+xVshIzzm/lAo7BV0q1vwpsplvddsj379dyFoJaMLmtTpXpglnyjhBu4A8l9W0sUYG3K
kZOIfSSKvKXHBy96tein04uMWYA8sP57L7SXfZksf9+kRiYHVDvvTXiGgQ6n9tYA0pZnPLlRQUoa
KifOtgvnbgOJ3arcw+TrgXziHl3dfV6rLSWn/KiMVs8gb2KIqm5A1tvTqo3uJNN6v7poO8D16mYp
rKzPD8ek9ipjCOYX6qgag50gTifzC+k9kvWObtOu4iAG97QybQmz7FYYnSz+Mbl3tod7Fs2r4Pbe
qzMwLP4UcK2ViQc+aEv8zuQFsFtLfzc0bBZEJZC95xwB/hXHLcBdADQ/UQli8Pfm0V49xe6Lx/Id
8znZh0r2RhozjT+fkN8g2/4mbux7o/kzF4nQziG6k7uREhP+W7Lb0e1N8GLskdgEirntJOucuc7N
Wa7DM809Gn99IPSUcil13LbKyCn8yADtrfHKRhS5RV3fyea+wlhChQ0EjZUDQ7Jeee2ryNBJkyRc
92Dvlec/qfpu6zjfvNzliGfUklZdNfufRsvnhXEFvy3R/2IGv+BEbod5TWi1jcsC7tTStAdouBVL
qifCoOyJLgK3Gum7XfMeyRh3vSyTJgySYRs8c0ZWwUGz7+f6pJ/edNr+Yjta5CgKc1ZJjzj8uWYq
118j558IzLsMp0FZ5O2ioyWHuSFKEsN+bOaRWr5Ny9SLweE6PEeKdjYDWy6AtX/WqOhfp3/O5yq4
0UE+rp7K4XgW2Pa93PkuUmuDzKly5G8JPeV9n2e6Zu/Sd3+kbJCz+6LUAcJ6rQgXYsaR3EbtSQUw
p1l8dguX8Adp7x88XkQocxhRbPznAbnRoBRYuzqSFdix+5alpeXTTnwYNxu7TqWvbxHH9XzIj/ry
uMNhXUQxrqFmxgEPF4YkCotDWQuDV5SANaFGDIPptY/6MaYuhrPfa1jQmUzhlLJDR++C22Q/OjDB
cJmvDydsIaQCqPbPykTBdvkZZIMZGNW5LoAhXbgjTuarCkTTUy4FQqCfC3ONtO1d/7s943X6JgpO
Tu+L6CmTG7BSuQmPjG/pCssvMiqimsiiO/zwhHVdPsADwrDcxg/iLQ/o69gLeeqp5+Rjplor8/gF
veB4u71i+nIY6/Z3rrD6RV/34q8rsDOSP5UL/McEswVkp4yApyAkcbSvXiBQds3JYrC/kTydIhbh
oTmPJkQ1XzrFs53+qJ7FsNOThHwPRLFIccM6lhPlD07myqVWKaskBTwXu8QgmmGW1YA6WH1fEvOe
rxf8cgtehugKuKQgKz0FUsrjQDRCIJG30ffHaAOSs9NUtNy+RXdokdjba6cCsw8V8u+bw0DWOC2B
cO62K6QNqXbK1CbzSF9PUGyDL63FNrKM5btH6H2DklWZ26bCz2Nl/igD+0tsE29PMOkwS8LQ3fWD
u3IN80j9EE3ZlYcBW1UhPogp6ILk3LqsrkauuUyEl6HnlaMRC7e71//d/WOw0RklDuCrDcdCl6T5
V0iDFj0ARY8tOFMKy6bvpvSe4sj/AySew3tyLZXRFHWqgsjr/ZYZsHKhXKz5VPjprTnJMjHT7JGL
YIUzCG7FDZ06sTKBa3rj3lhkw6xQJVvBLVkrgWmZ/o0sZzkXJOUNng99CnwReW48wBqPbtloPRhF
C/Ovo6lfX1K1msdz0TQaQlspJau5Gwofv486IJ/BL2opCLuiuuxwQIoYCxTYLPqMJRQQp7hlQdM1
ufv75yG/3UEYodk2zItnBxgNs3YC5oYnHTDvdPaXui1TE39YuVRrCR8i9U8SJlXdnYY5ahflPkjV
J1kLpmmqariPuS6oiuGI/WBxsWHh2GKHSKmekPPYFWhdEQbWZdlRTMXkGZrIYllaDzbPCRrFs3/4
XJ5P32AVA80WThpBNVpiaZaV8ZNd5Pb5Tthl08CvfRVhEn1AVi0omGrzRk78ZiH8Xr5/GqthTaOx
qzsRv4GekuWh7NxjxXhwnu0LxHiDITkZFtMc1qwY5YRCf5mMQb5tsXmM7+Ua+bwXy9Cc975K9mWa
fRGSMMBwRx2kBQHZ+m040GsMxpYb+g7QrFxaZGIr10DgT9yyA7owxCexsUpuQHjeyKy3z1l8rkTS
oCtlqu+23bH/Hcmm+PiXiuSnFedBumKev/K2v8JeES7sNjnplIw/DEHR+LPj/wFWk3C3XKhb2Pp/
KIAi+lHCHREUvOmLOPIpZ49HkVHINxMCReYpKBg1wosdXwsfuN/KD9Ora2JHlhJTioQGHLLQVs2b
JvqMQJHKfjiehCV9gOBYQIi0C1EKJccgrszlOhM67YG/xm8BMITbNVLDdyv7KZUmYKLB2DOBgw7i
jEtV+UKSo1jDaDzDiZROc3BHdGOsKe0RjNKXg3tp0mAaT+SB5NKiWAfJCsTuc6AjxGZGSjWO/nXB
dGKvFn9GqdF7L/B3eDXctkWnAqXo1DFbp7UqApbdcD4WTsXoDYzJy/acSOE1t/fMAgKESPKxrQNn
R7NiDUy/M++tcK3aSRrwGwGHmS2FUHepwqsGcWme1ewB4r/H2BIIjNWGh6IrqSW6Cz9KELQF5jxq
YuJaR2H9Ptt1fwdo5tgoLEX3hTZbkx+4HL1VV5XZm0bLA/aecEQpTltr9JHr1sFki3HB2/BPa/Xn
T/4EbhUSZU6PSiL8uxxdMBvynDvoB4FX7tlAmLRx5GaQBDNoNkDDWG/xLOHk89mEqD565uW+sYOo
kOD5O3vnXsa5a0NFJfMBs44N7TGYrYWEX60r7F1OhAqj9vWa3wiuB+gAekLibHD1nPGZHRPShqlG
Gr54PiBSO0cCAigv+JmdcDxu+0ollza9LogNc0P/nQe1PyEMgY2lSPx20yoQFWRWHxbSHiYCVLcD
EuBqTHA3nzHJ+6N9cJC0Ls6fUK+USnE8MeayOBIDVPUKt8X8zGbcmHGRXL2WO8mPhFPbLS6oKWWu
xapBZyMlQjZTtE8rcRSFzuTSMKzegSKc++xzLcVLemtMta2QcvUBvsIJo6lhcOhHkeI94Ip6Vm51
KAjGrGoCfg4puff0yU0KvucD6Ea/SMpYfAsQ4zvSWsjM3gIiTm8n1OR0qZAWYnjvilBXgWd9Xn7C
cBs2pkriRETJ9oJOvcFtym1j55XaIOUok9eNCjmmOjM8DSKMmLfCLul0tLiRNPdWJqA6KieBSDJD
/79e0kYDfB+Fxblb4+qxRwK40N12o6jCFnTtkFlBv2F1+Csrd+q9Y9+xIymAuE6gRpcDgV/PmNF6
a1w0Mi18cAvZxqVaD5clC+alAoGXTwbz5nXGswt2G4LDC7l+/8oaqz8fC9FiEK0LklWFb1ZjWnvq
oKPecokv8C7m8RkYXL7gA888+IdbL/ULCdRX7leO/nZTfCmqes5gf0zKR0L8MboY/oyMU4WD5c/F
BCqBzDopE5m76hGsktVmKAcKDyufXACz4++CJNHyEV4n7WBFypNQ7JzU4HqoMRoYNm1/ZlaI5x+V
ridRplVTOqRbxCkau60E5NOZsgl4aOO40JnHOK9RsOTHkBl0Eafi8DfQR24BGINsVqKD5hctwnqZ
Ymzznhsc8OfNRF9ap++si5b9BWW04AeD+ak7Uafd2pdu7p+tQY8mI31gwC91TOHG9EZkn8yz579H
IiWKSK/Oa2lo88u2Cyq14Q+HnhJaY7TR+V+t3wxqMrlY8cIbOWXDQNx/qzWxLkGwA9mwNyeNLSgI
O1PoJ5uKwEN1OCqI/R2bLpQIAssbDeJKlz3LJZOmsHxtD0DbPVx3hNp3PTfaKUcv1Wbygf+v/21e
rrnkZk+OPH71CI3A/K+C9GrHvGw74n/JhmZ+gtNs52aTHfx797YvIZXmWj3KBisIe3u0xvD0Vv+B
OzEMGVJZhxy+8GtAy1SMOq+6TXqo9Z9+fi5i+JYTYxyHu12iMFSF7pgK0tpeg/xixIfYi21B9ZYY
/yLeSRRXM0sBd57xuZT7MVQb/c80QjDSSXITpWpA+2xPgTKK1f4TXSGWU43RHeVKFFkNroQgnNsI
WyAKx+dOBImqCY1ckXrnfy8jZzC0D3vt2pZSjJTHHkFtqIr7oHSQDrci7tgrO+JFjHXCluMHU536
Elh5uxLB5dL/bc4eWctKAT6wMQmelVu3tZgjsCRnHkPSz7QicmANgvLado7RLJMXcvOr5Xp3rZW2
6cw4AKJ10DQIY6xwyj0STLQXaemKHkNOm280BVfyX96VqWhWXjNluwppvRitbGLgU0eXJ1YaLdgG
sIaeQybTotmt08WHzR3KjP0IhYUW4LUtiVlM7zhmnc/s7DBq6vo6g94baHz7xuOZ6GvqVVu33Q/0
oMy0OXG+dhTBL4+Jw2NlxV0yDhsYJpJF+vymaZRxcbafI2t5W7xOrAWUqvsJsMcZoSIp/rqf7W9A
TqaIogRgByNExQS+hq2lw2DMX0MKgAbTidVyMdd+tsrhM3Nbbzruu0D3y0dU9tquktL1Jn+uHTCJ
lxXEReKXgdEwYSS8p3J5+HYFhlCnqZplyBzN8bvyY0FxZEdeFdneMLLdr7JaSMCXtrd7pCdJe3/h
9TSqqWNIqjTf0OmE6Nekblk82wCBHuCy304Hpy3boXaICBbl0YRNYW5zh5MoJk05RhGtoabc38yi
wwBXYC5PSmd/GUEhosTNWNq7kn/+7EpbgQTgc1SQoQj5jyGe9Sju+Mow5maeuAbnF4cA8ZynQ4l7
jwpYzKt/ao3jyep2uFcsRQZedPIJCwxA/p0ATKYOPOofvUtGkVW9wcYr5Tq6npnhSSDCKLgas4Xr
+VeQABJX1O+6JRS3D2pcoEVypUqvGXcene2sRzcxxVdl3tBo0I+cQhEUO7MhWsyH7c1zx+sO/Rfo
YS5lO6FEsUBTp8kt94T7GRVNPgSuvcsNmuSQvJ+IIlgkmATQRKJnHvkOySaf9Epd5SQnBxxRLGb5
lF7/zBa69GG5BQTdwGUnBrty7QjVjVftsQhu25YAKzrqOK9sTTqcSOSMIuKWlzngbUS9WzUFUfRx
sQ2j/GSxRLPjM+qXm5vMIkrenGB2dXZ04xPwutJc1k/7DnLigQT2LcbJVp9LK3Ti0cAJdD87c8f0
9ber04jZAvymGVvMOr2ubERIoccCexpcFAWAJS/rcLwbqqvrKnyPhrr1kPOZr59k3wjBSH58ek9L
HqPBYgdR3RJK/22cRcv7rjtPcq9UHr7J6czrBvxFAqb99VHo2SV9QiHCzXT5LBklFDNdKMWJvLsS
vEAaDJA9Ft7XXAOvVoyv8KwD9Nhp8bMew3CFxkxJrwc8dUN9libq4Gs527ZXb49cZIF4ttDhF+jH
afvhz5If9qVuVGxcYM6rFxNELSFacqEsv/Ophd1n3Zx16ukl1IOVEjdL0rfc3LZ+IarGIQz8SM+K
7hyKRkFH4T32wJfaqhx+2fkP2Ob/Y8vYl2MoPJhzxNmODjYwsWRWYc04dF6VSPM7vAkDaEQegrRn
2JMVyPkOmtQBsGOfcSY6FTbf9biJ9z+gf7ymnvT0hQGBh8BDSRex+C7qh5vY3gusBQ6EyEjfiI1s
sOQB/at+SY17g3lDtjb9l8E+0toXXmPaWpLc619qynxpdzyIkUEKk6ujMFNW6AfK0jeFu3ee3Z80
X2XI6f32nuItJgjK2XCcwPB/QGftGWl5yQuN1G97T3Hvp1NsY3xB/7US9tBgTeaVOc2RqRI6KqxD
iWCZoBq4zOYURjWF9nhMU2GqK8hqY70xIUaLOE4LtMntWsnlvSBXbRsdr0LV4nUdt2yr4cnH1OiD
Dd/KXi1wQ3QypMyUtxeiPq8yI6AxzSsWbJgesKTFg1HE/LuciA6JNuHfMw2VXT5HoUDDWvjBxbil
yCUT0TwShjCkeZTdTIiifoGVm+P+kLDyVGzrAlffTiLNCMq/FLiCMarnN56f0A/ZtXnSz6SNvHOD
PetjpKg2kuMVxLy1sSagSCy3TwJZgX7gYfh5OEHtOxI7h+ApxiPxXfdmrtRS1FbCIjM0lA5Z5N/k
jVbpN43hW4ueOu2h3jLGHkHiV6Bg/QI44Sm/0oZaX/BzZaqMQmQIttY3XOAO3efkEFRxdPMxJIdb
iu93Wd41+ieBFYPwyhfNevYSi5mS+GtQXrOmCR6cPZruIOdhrE5C/28eAVtubMEeVIVS9epFzTRW
lRLDLa1E4CkWRz83LwC7XcCRdvNZ0WhncZM6GXRMU0ImJ592cGAdg70HPAF/dJ49+N8qVPIewoo2
l9ZA2spb8bTZWf4h1yc69gWuef0HOuS0QQ3w+U8InwjfkX+xvrBEsgXIx08Yh5DsKbJIOjfUcDZu
XBqpW/P/BYGB9wSxk+SIwCcigKUqMJ3TBC9EOmwvpU0ZjLN5N/NdpgSdkGRV+RoQKHxqpJiOXIgU
/4T2ZVikOq4Ojr4vFN3s58Da0qORZND943HP7lZhYh+Me/KJKVdFBm4p8qKuZ+yg1aCueTAM14sf
u+qXHqmBX3n6nWqh30EAYhCl67LxAvd11uggOMR2YLbCL8tCqDMXeaJzlzlaBsLq9ijh/92QE3je
ibEIajn2xTgGExE8cTa68jdXS5Xb45KCrcJPU/f+XxKKJGwOSQmJfrVvSFjMJLNOzFpc+VHTDnp8
eDLWC+8c5WjFKlhLk1hovc1qqneU40Ya00zapCibwh6hXPzQJQI1VFL97RGwClhXU8GeLVZp6IbU
7EbfuShdOMmsDijWDXtzzq28spEPafUoiE8oz3cTPjTxwUvlEPqsHaAGGyBCJkLRkFxgTnEtUjbV
40paLuKREmnc0rPsevlfntY30iJiJZhXuCA7ewTKNUaK9t97ry978EAO/EtpBCHlusD1Xs95is/f
ZJzxaoV1X0J+dRO7rNXx5fKGjWQ2s0Sz1W+I8HXVit4G3AHi8bkkY1V0ju43qtgXsYDkS0DYJ+2q
oVt4WAlnXZ014WDIYpGzNnJlM1G45eHkrAMSjr9GF35RCT1XXySUzFmTb/70EXm5Kafw5NobfASV
1mSAoAFZCZ2vMsOSJ+IJYT+XMyb5aSZ4OB/mOGnLC1M8uGuSkoYHI3Tdnn2jUViXHQb2NoVOOLNG
0G12XAf69iRHzlmBIWj2ouAgPpBOjwG/n18paZxAIOH1E4BZD1ThjK5VFtI2AYERw8Z60ue9tfSp
pJwK64a3kp1SScDZ6ZtPY2p8it0cBxckK7SsnUs+1cW35R4ZQR3uv0ftD6BxQ+dHoV7SbascVZGB
8mY8YpiOestGKzYCHc4m+87Sjx6ufpJmq8e4+ZBOuNa4bYw8xf09VJF7QDQQ8HD1D9NsP9CjEFiJ
+HtAmXb/s3x25+qZo1Lj/PqpU4ORtMO1QmDfL9j6F5AkI32oT4ggGDYbqTzxLRgJjynW8+eCJSdT
EHsaELo48Hh5IbztrYDiC7245M1Nbu5QKBhOhrXgEKgaohmBj3Bc6mt1Q0o9YAMhEgK5Tdei5hgv
eBT5LBNVkvuExvPEYhujSstDA+es4vFOOdZ/YN41HYzM+TiOKfMyww73cGJ2aGGJWWih6hq25QYI
7pi/22w8Q4bvPZU/yzd1/q2F5l5PF4pL7Sl0Ts+I7g5KsjP4IfCdyJ0dwoKFHhhYF6hS3T6yjXSl
cRMsQGdZXpY3a1jrGGbW1U24ojYUPepcKxKG+V9k9gTuP8JjCh4hEG8e71YWt687KK4umSyDxOpn
ezKQE+xQadoNtIKvObeGDdwDosZ27/bcXS982N6/wiKrqkTOprmDQzKahxLzzWqUiyRQSgXEQF5g
v8Ykdomy9551HIYwAHVpjG9epoN0DzcagDIm7ivImwnuM3oZ6hcLkyeJSaujnvdPPE13WUl3MTvK
1QuVsMTCj05NVGIR8ywba+K3EectHXwTNef4SjfWCpIE3WCgyUBhD7IDdDF7T4aVaknXYLAirWMA
oetuhT5KB0/bOI5IuZM5WBXZorXPkhbl4UehppfEeELtfTZPEJ/tHj+e/uo3EABdByZN3kEX31Ra
JQ3umjDBePLlbwuL6MBQkZym8drdcg2MnFIkij9041FFJw/e+ecTyqkfELcKLYCuF4VUI+yKj4Sn
h4ds25KQiI1g35d8Elmaq5bI324Gf/3nnGFbLRQRxoo9SfrJAkkZLrgH6DiXQMjktfyniwqdtQNo
YLUDD2Si0XtouRBAkbtlnHFKzcZJbSC0DVJNe5JSbB74ns5wLOI2VInXFDtWUwLEZZn1/W4pf1ir
x15pkGvpHcH/3GySyWS98YuM9zqaZcPlkI+8dxJ+KRCs+hDg2rIdPR2Nm387w1qeCmKfaNtnlo8C
p26xKv1PGoMZExWZy0KVw8b1j5qOSDc/WoDxD829CDpCRqWOTB2rLuOAXwI5dFd+3CxlLomj2o1f
UUwCbzEzMxAw10gsWJCy8rHPkvpOIvrjeQPpmKyRtP0TcWS0BJqStDJnOAQVa1oYAhEVnUr2Jysl
7GJEaJTWdkFJFvvsC9FLnFmnFwsRH9QXqPsgFZzxUEirVgXhsDXYOmoF/U1/vkKgpQU+LGTdnYZr
z+xBY91Q5yQZMvR/3NgzA5jW4lTaH1DnezeDxWpv7UURJcErmB51EfAszocxIxeJHBy8mRyq+Cad
oUl/4cdtMbfmU8iIur/cwCBpGetaXjWVKPpWc1D9ETqTS5QiqnS4lOluSkJPcuvGIApfg9nXIc78
I5WvAW8igOx52vVLoVXANlukKWf4oDcCn6/2dBkWNTNs+3KXYQIGCP0A+PEjIvoYWrHvb38fZ3+3
75e8Gm5mhS1EUXy0MbrcM+52wt4wOEazBkEaqjNfgk44I5culI4n3YjOlwlHBXCldb+dCw6rLenM
wBv7kYcBi20HYtDVJg7+nKxW2qxbJETh+BKq/Z30ZuJDxco12ZaJWGXD6/CI7OSNs8hN1Y1Pq15B
9l0i3I0ikiO0FnG2TNTLaOQHIdlQw7gV7Z3YroJ1RGSl4VGm1iFLBJUrD5B350FIuop6fGaalI+y
yfx8gVu3nSYAZ7FoImJ2Pf0QDEo4ef4EDwX4inSw8hQiPzwthu1/sKFHsC/CCp/RatCLZUOehAND
oolj/YCyRNkxspqDVG0W5Gn471fE4u9lNaLrNyL47um6iEmd3vMYehA4hHxJB4mquFPCyRoSUtD2
Otz7hKFgaYDFLWLYd5cIJvaR0+TltxqGobJw/PCO29o/vxYQ+z4VyBUat6odqDaIo0mERh9dpGKb
N/X5J04VazzigiBi/jPTdt6vT6YXsh2lcID21JuLIb+BtJx2MgheDL6JeYXPIYKcwzDz31VNTQY3
WQ1dEzytNBCE8oUWNjCUCHeV5dDCCbxpquwQgbOjUJjBbnHCVFam28l9U4n+mxfmV3dI52X49f4t
iR6/1yiOmHIaQA27kCmXd71N3PI1H+s80RJbZTY2fxsmYP7jlKrxIdK1sQqAXIeomTv1msJp2bZF
wZEETDmQh/1M355osKtXHGsS9tH7pfjnNvmO6V/LV9a6okfBVMJw4Vx7uJ92gRSeLGpgHFv+5rja
vG0Q5Cn94HPrSBzjuoxTSZDdeI63ZApVbhgZB1JO+PUWarO4MFrhIPNGSBBSUfl7/4BVopBeuNUY
AADzDi4vDXLPuh42ZudabdOCGwKyPw8x2D8yEv61jeoC/NtHzUt1q9lkc9y+KWXb/PDcXin+Zrh3
ugiWc6DIyET5wphXTiGbCL43t8RymJXOPC281k6/u7Gau8aGTYQtF2YGcLq4Xq22EUXIwW//rnjT
vtTyAlqKdfVhWoGzGq68G1lWxC785kg/YZSI0A0X+5iS1qZEBGyuTgEBAI516ZW5iTAuTfxSL5Dg
V3mVTW8zcBUdJDOpHFxVhB1N8pNDrk2JtpFobw88yRKHt96lIvr/ccQerowCld+cXKI3uifh2ewl
txCz1XBfo3/ryBEY3SOQ6HgWcARYrzBzf0SRUepbQI+I09+i1Hb+FuFyxKK+29FjMMc9w3uG3rEY
ySd5JFlTKpMmpfEkf6XJl9gajH2qY2YjZu9DTMP2+wHmWWPtupuvkkhTeN/HM9AGJH9MDHg3/kux
F8MT7maFahcmsoJXX4cB5hjKdAWWjV6DjlkyB4yMsHduRB1ALWx9P2/41pqjaWUl+QHW07bwCvhf
/Le41EbKdseR4zYJLdtgfNqDRT2++MX3/LagL6wEJNbg53JnK1kUsdAhWoRm1p33tr/ItUM3IERN
FNsSvqlh/kmq5EiFqO4kjFFR+hugNGcwVPC5Gth2QOqf/Wgy11ZlNJaCvTW7WadIu60csLKCgmAh
8HuqCDNIL+WdnMTnlNqmkAr9FmP7Nxn1FH0nZqYTptQsf7zmMZOozTxF+xHeX2ieMNcW19XrxIac
1rq2rJ+zeBxgbo4Q2aVjJdDInE2TklehIUYYL1w8x0WDJSpOoNwBL8vOAKtYcIyJGSmBeYvQ2p8M
0TuB/XoRVhB7LvGcFlmMxGxFPa/JuBZzWoqC6JHfSNVhwB9HhumJlCmRelJGE6vPEXEZRWx1Av6J
ogjM7CeUTUuckZiXVp/NRxB+9cDdfB0VtO6Rwp0cFa/VwpvCvnCkomScCaFeOxkLmjbe0yY9RY+F
ppEcwtoXHRyBN5bC11wbNyCBFXKhC9VFE074L70tjfAXYndXxhEFkUlCaINLQuHBcNd77sdWpxx6
KkoHjHG6NgAvU9hkvxT+ogpYkj5X+WorC3UTo64WUSg2Fp/aHhCekIFtYTovA/ZVxODeMKPK9GKC
hIe107hUpU24fblDHG1ql8f9hIwel7OcVk6oIkR0MuCS4gkWwHyj/jLp41+UpkRT12md/koQFaQc
wo6yYHVb2lIrC4kK4mcPinw770x9L1ImCggfEYQAV1nkHI3Nil13u8JEKlzwuzCKtyTHgeA4v9Vc
SrfAWpDYxbAok0xF/AqWHALeGO1bFl4ZwFvEwJ2fg02hpLJLoPqpXDDZNiWV0aDZrQ6rX29Fe3VR
ddQ1ofhfNfBTkoMbg0brdGay3lfZTdgk7rhjqkvditzFyB37SoWMLHFKkosNpo4CTNc3
`pragma protect end_protected
