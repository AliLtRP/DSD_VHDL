// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C5HZmqCRu4ONkBNJMcY1YyFdsNqBdJh+yfIm8akx7qholvL0E0LVz/4prLJBTdEV
QPik0Vx9N324bbaVl7tRRVM1cgXltim/eSod3A+fG6SeS50RI/roxjQsKQDfcN3J
hJwhL4whz2aAcAiO2PTuHfsmTE0FzZ/xbL8y2Xi4BmI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3504)
usOVQ9lAVkUQdN0cNSvvGzfZ/qYVkg+EylI/mPpIBJprvoEDT4jO/lt/Je8YOe4m
SG1jusqPbeGb3QfTfsuwb51M1/gPSO07K2T3qvd0u1SvEIX5pkDvdAbbNHMXSOUr
zcHCHmxOA2VWLPkARuJRKSwFbG9y8CXzGmSdvCvoqQs3edeFUqz2M5IDNXUPiCR2
yJqTWPMfvD9Hh5p0HdCECU9XFs6ww3jB14t176fkHRWH9yDfuMhUFgoAK5hapN9l
ERvpvp5Xg8FAoQJ++hvhj/33o2sxod+V22S0ODqgVs0jp3EPCbRcyY4uYYbCW9Ac
KkqNOrGqpfcsZ9OS0V4oQkt1obCCsKL6MABKyWSz71UtwbcQ2zLsVWUSlnrGsQu6
afxJHzgBNjYUAil/wmqFUkplt0x+vIXYVVwy8ptGkz8Il2kl65TS0VbdHQwwj+Jq
WyW+b44K093gTR3EaCtNP03DRNdTN5Eu6rFaMEcBieuZHYSCUb+p4vYgjArSjg3G
nhQZAA0vafQlALCiOjWlT6HfhBI1KUwx31o5aze6E7xpoxCDFtI/5ZgcVASPOX3M
poPzPZRuaPpI4gF1E5BDOEPlgqx6rKCrprxLfeaihm5VHed/SWJUiVc2v6BlzniV
gtRLzWZ6hTdLKWN0K9AF+7WjvlXpgiYsyPKuzFtT32YivukZRgMGNOHQxAva5mwC
Q0av++vAlsnnbI2ZnlnwfYLGGZLi/c5MnwTgCPBj8KgIwaEAZ77Y/RxMSSppBD6X
sZFFW9fAw9/OdcKGpHGgHcjaFrMahVGMClLIuTYbB11ELyqosdHltzgwT/VEVLqq
vLBRFqpUwovRu0DQlG5rmUHhFJ11jK/0Nh4hEVdSRPWwy3sGQiUoHw4g/JtbnXPP
jkreAX3XPve+JNTuSdw+/cLglklhaMfmS8tTUPbiIENnHKm58SV8SIfpoTU+JBcE
uzzMqrY3hZXsdi90pWd80QYVkLFluh45AxX0O9QD4RKB2kWUrv/rIimOQ8m+HwJI
+WBIiVHG3cxByg299Fu8wYCinEj/D/uVuW5vvKF8KHewvqsT5gQ3jh7WiOzK2hH0
j5noBoJs09GU7hO0nYru+nhlPv32kYgVUYWLGuVL9rYTqZwq8VoaSkEU3bfCCYLl
xFbE6r/Mvq1KtY9drGaFyo2FRPzMOsOxd7IHs33l9w83fsIACQtmJneYt/wNIXSb
ie6xqv95NRyrYbuxk1m2AO/cxpnYh3j2gMtw7ETlAE4XOmfOl2ecZdo5hDsoN+Si
+oGzdlCo3ixHMKv8Nwkd5CccZSaxCDkt47hm0i5taXgrb959pEAorUeaT3gQ8kG+
cA/bTnEtzuOG4qcWJPUoUjQYdCKegGbtgIZt9hBOWJJvZONw7Z5EhtensZ80LDaQ
VttvndOXfQpGP/wyVqQGdny05R4uZw9+2OfkI/8R2Pgo97LVbUaILjwBhDSrof+B
9gQYklbizaYHjnQZr2D/vhRSgRQC3z/u80yEJ3YNGSqg0AgNl1Sd0dKfltAjKAAc
DWnC+IwCb1a1udyRK1xmgY6bNriCW+j7FCtUyEoQMP6efkNlYWqjtwQplUkFd7v2
DYmPr5cg1EIMei2uQJqs5n8SmqWYht8VrsIv2yuGrg/oisiWgWmtQxeKGquj10pe
I3lOV4juVoeSepP2lllqMbbUAwAAW+VDBdh7aVzvWpi2u3Rn8H9sykdI/W8dMV/7
j40JVTIEBJdNxvgOf19Z4iCPfdb30OkNlxzxj2yoEm5KNz1C22dmuFh3Gyz414Wc
g1IGIsOmm7tx/ntcxp4fQnxBlxfFj95Ty/pulHcHIvIx+xaek9KnBTCfSNoNsXfX
QffSr1OUyds+1meUwddmY/9g5a9ceaIbGXwe4Xol20TX865796yveU/Soz1d+/qs
MfKxqNLUCExO1BoEC1X/uYdGk5fVaFG2ivkAgYEZfoNa+7J7xhVfCo23kXhkYAe/
bufsEHAt5+ve1YiJcnBaprtjd5oeaFBmyjs3cZTueF3Ou+WJn2q+6n5zeRg5gJ3m
eAqaiO0QNmVpJK1o3VBE4zGlFfDZRsxlPgFUrO3vHRRSd1SnlrezRc6f5RaIr2JY
LMKBIZjeAz/q5UjZtcdEJFPzG787jvJJnEokJp5lUZQpBG/dCOn8El1DmbNgIa+y
WsIuw3SMvgt8Z556DxeBN91mxOl8rbOkKIW5syAgNzZc3f5fQtkgkNBzRvTW6wiG
/2a8cE2ZWPu/MpGYdrrLF2mJ5KtjnsGFzY9qcYI38h5DKPz3Ywd17qeuFqu5FRZB
11+o2mCbDQVzcc4Wuviy8rRPDQWozH3+pZjzBo0g6Ycojhr2aY0m6qzyjfsHOmvh
+OC0F/Gv4Bj5iZU4zGVMDCaZEeaU/sQku5gqeK5Lgh9kx7z6huZpj0lyqleJ2IA8
gz5WMTFypOJb/fzMUakgynCd15EqTGZKsyin9PkccnVKYxr8dDEDiDJrYYgigwYL
iIn702Qp+Lj2w2PXg8MO2d8LSoEX4fRMPvy1AVnE+XcTmF2OfwldTeALy267V7QG
UGkYMJrsudEI5kuNBZmI8p5z8+aF1mW8BQe1kIBgnTducP0PL4NcvovjP2Lp8Arj
vyPl8UjwIw6Nprr5L+GTXzc0spk8+DeyELk5jRQC8IBSr+cKhI15KF70zANp0+ng
Dz3P7E4/Y9eo1cGQ0WnaR1y0pWhHvmWyHEDD3z4cIIQ2nvtJ5IZe8k5HiFmecu+X
qGQ/uLp1stnvbmlEr/i/guhZzywvt3mlekFSp6BrDqmyXU5SOdU1TTm18AOo9H8s
eKQGFbursDIEzbT9RfCsOYRCe68rEhU7d3XYTjPw1K8sHtwUMRp/fo9TvkDZq1xL
jLcO3HPrgc+oGglOzL3FIn8Nn+Cuey3E/iH2KJiKZRaH55GolB0j3G2lYTwjky9u
q2DvxKryoMMkLt0y+9nQ+/1dt6hoNl7tU01PeWcnhYAA0Y8t0HVNC+NncaVF/ApS
zEkkGaB/egu9ApVj75/h/0aS7NdwrOjKEqAPDVranIusV9ArZFz97FDrKr6w9JQ4
AKPeE0G0ZttGFsNYs96W4N6Oh/oe3/WWXJUgPmrVPFqaqswIHvRtnD72auzVaPvq
Fn5dC4JGW7f1Xwzs4g3h1cBiePyY3Y/Q7veYux3d+vp6dtqupgZREMX8Noo+Irow
m4q5M6EfuzhBsg4Xwv1aH+TqMOM0UDVh7m/rirTNM0wsqWZaTgjU9ApO280b0Zoi
1vWeZO2BaJhHJwM0Q/E/hYLtslMdGVtzDyIQqseU+X7kvPQkIfkm1oNCNW6k7KIw
DAu2vSAZRjPzTEln0RpGTkx3IADR6yVTPBXOTZ0wRriOYK8zlTmF+Jvk5Mu5868j
hQnwUG861C6cMLMRyFK4b+alwUep/kPtyF07oiWnAqoGbCFQRim3Y1Ky7htY5A7t
+jTBr1MYNKsYD4Vt9yefWEOZN/6iDMogS9gMBnoSV2bLWrRnDkHqBMUvwMIxhz0U
2FcwKd9veByi+QGfc40n1YcvZ0vT6iF+1bhiowK4/Rt+MNetvoY8XxWj0EJMHhSv
H2gHVZxglcR8m39c1ziKNpZEqyMjzXkFjRz/h5fsdzTayPu36awaf0HGh8mjGswd
yyrLlHVuRI4jAjzKDztFp3WdM88u1IhpLxa5EFyONiRaLRhHSBS73jbOaPv9G6Ew
lod2SpJAMWVlirEHUElvel/PqVqqID5tdX5BjEoVgWCWPGD0GVWDsVI/5ZDuK6RA
Agiiloyi7liq/cyM5AIGm4Rup1cOWgDH/UX6go+Qes3yxwGWO1iH1jKG56A/mqLB
VLv/q104vICkDYNsThwg0KpIVsmo7Oqee49107tWL+BWTypnqHfnVzki3C5xfwey
8nZRb/9fetIYeM9OMRrLFvFXq3ylisj/c1m6O354AUsXaUV2cl6xdd9DVeSKXeYo
IjEd2zu4yb9oHDxfWk6TvJezZ0OpvufO74PAeY6aW6iL28jqDWwgOG1xRRjxUbXe
KIFZKdPHyyGLxa5stFt06pMHmmqOANtdUHht0WtmWLfjijEWnrv6qB1kpG5ygw7G
rRpB7yxUbrIsTw2jU6F6XBpEqVwNICoFp5l3RebfsBoyC9xftDG2CI3KFy1cYOsX
W4NUYbNX7Nq8fpN/DSjZ6+gehIrfJLbcnU6Y6gxXHXQEBKVecp0mZUsntEnmcakc
MC35Pv/Rs7dp5U+lnUmYQKM+6OD/s8sw9vUR7UWBvDkgg5qQjrQu7YJhPrTJmFLv
/VIYldMoM3z0fvc/24AJX240aSKQO5reWXXO9zt3hCY3XDvf2tA2BJy7bj1LJc2d
GE3v5HxKD+YebZkorKcNaV8U9O3aie9i3F228bmaCr5G1pfUn/so6B6mN8m7nfyD
MUsdWwzRBJvA9HQU+EDceUzinF0KWWVvE2Bjq1EDlH5H0n0cMPI7ms5CKpM7hBXA
0eO2a8w9KZeiG/LGH0stC32M8SWwxPCdqd6Nd0HZjaV+W/oKx8O9M59eqsKY0uUl
iTa1jMlnc2GlmikA8hnop5HPkQF3Am8SW31M6Yid7GpX0VGb30qaDvdXZznJikqn
K30TplW9JaW7PpVy/vACvhVM5l/r9SuYscT5f/YxsanqiAAqUV0x2sOUYUSnVx6W
`pragma protect end_protected
