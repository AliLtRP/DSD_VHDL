// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P8FFQX0SCwJ7mW1UGFd99x4Fi4D+yZXhKZaUzuRfDigw9hH+p7aNtFgkjgQyWdAo
WPaeHW5bVZfUv/R0BHazq6ktp9mtygezVBvnIPTEuDUPiIMiHISxh6U6lowjtqSe
4yLjLNQmcPnBZekL1Vfcde4r++1oYZjQYC/0mzxsutQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19536)
0yjGO/ui5P2rpdOCPLOZCna7X4EdQw3fr+ALKFHCI1gGOXYjgwCQ+6IcKOtPGMFm
tAJTr0I1OIJYiDDf/urkIA6gSlf+s3R5bFL3LrPKjrlpq+g2kXA3MSl//9DrQYiy
z1C9yR1wFQvlgOxTVklbJO4xaFISSb3XzM/WwVPtm6J4+pQG9KXeFT3DMFykOoCL
VfYb4dns6ZjXop5ckx1Vh8C7rLEH6JTNOd0O1UubxbMFTS4n18zFXmv0eamvmHe3
ouhuAtAuel/X302d5UoWwJxeY/l6mj32088712wPjY6NLXAYmrUiA9teXpYR4Rv9
yNQLLX+Oy2A1vYm3oCgWcXCI0nsNIDsNtuaywrLz2A5DnSy+JOT+wiapudc8kkri
ITtnS1MTuJc1v64R6p/hRnmdTSsFqRXrgB+LUZ0g9zbdkZuMM+vG/4qcB/csZoMZ
4azt9D1gbjS/e0kzhXyxADLEkSOIlr+iSg4UHcpCH0/2fImmugAWyIu1jTswtN+F
LVACY3cKvrlUl+hP3/hPBpdVlkMCADVZ7gTiOD9SEonJ99SFMZN1S81S0QpwM5JZ
hu7EfCg9EyCWJwqxvVUSMwKP7HranfG/WAyCXVVS7s+K36pH1CIkoAPom2mMAUrZ
8tOM29FtjBbi2yFbgIzddXTBP7nq5et/yQqCs4Vm45lHaTH9lXCFPWAYXDb8J0F3
cwex34oFrhY7ce2lgqHUx85HLxccCjPdHx+yhYOvIRrS4QVdnh+3xfJwSi0ljtqz
+NvuJiRpsmO3DGV42qBQ6uEeKbG07LekQsd5WlqPJ2tfqxJGbHig9NjhH2MfuYl+
GlpGXjHL9NavvPL4Ot3iTuTUXQcUQzAsmT55Lk+4n3zZqHvhyUhfa+iDA1+e0Car
WwmW+UNqEwLhKjZI28wur75aennG/avIPdVFKu1e70j+qYL+ghZPbkL8LEdSIBPH
jd3IuY3oOloVzYiIlUQI2AwiHBR7lSlfZ7ORatwWwvglEWQl1DUO5VfKQu1kDQlV
C1zrHkdkKqYfnjI7Rw9xtArObbNMovSB23uEGQ/rsFBgaeaFFabjskb0Apc6n43s
yrUYwofQiG6B8sy0yD3gbjb3WYrfgskZ9PASXwp6MvNmWUk4A6l5iW05TWMVDo6u
1v+giVvkzUBwxh1pTeTq7AP2fNKn7s1JTvEltw7EM9MLEhFEgw8dkbi+1pMv1un2
n9PToV3A0Ee8YF2wHtxGEIzSSePco4j0DiBbjpErJE/ZBxw8joSwE1tZ9dm2BoUt
laBcYjk3S7VJWnhWUspoYuB9EMn6hTCLhk/1D3dLmL+5wKH88ZF3lk7Gu+eeJrB1
pq0fS1CUAACh8ddZKYoFKolUDzehQpFXo3W88P7FAQ1wUwYwiseYXEtcXhYMEzNJ
4K4HY+HQS/qB9kqGswSAvLhv93IEgnx924vuCYgmz2SWww+8DOt/1Pl1FNyXDCKb
+AIJ0jS2IqzpfxPsGtMvLcxtHsQ81ePSok1A0D20KztatFEZLwteMlCYxSE5qiWt
odr5lxOe6VG9TWzUD/vwnr+aFy40UXB1sTqZGHzRlsTG8DibmV4RjSoyKlTaVFU0
nOjMSsubZhnitwBbfBigNjmjITAlM5ZkbZceghoG93jKxUQsic2fDHkCv9+JkXqs
jwFvRlbxHY/ZQUrbRfh0/xWn6lWMGtU8+Vwr/OGwIZfO2iXc9IZOaZKE2dEcnF/5
aMfAsWYQTydAYEWMaUln1mxmsbfj0A4AdGPVpSjL/aBFWiWYYTcpF5+rF8o/hrff
yt4HEW6iktgAtSU3AtOGFTWaavBXQSZkFzBjZpJsOZDr63Db3pSCSS+LgHBYq0ur
eptPIehqo1W7OunqLQduM0NVkC0Tqrlf4zvb0P7DtvRci3ZIuSrJzWVQ9dXL0Oir
RqHdfRPW4aMqhamv3BxCDHmoCNeOEGqDl36frVLbq6VPmgLzoHokkLN8qVIfnwtE
8ViRczxiDiqtLNS+F3qJZFP53MsyT9k9bRqJwSOaBBoBojeMBlnpTgRqV15RG+9l
t8CFOMQCXRyPx5W/WbcZwIhsjfDoO5iQIvRYhvn9ZTi1Z+tLqWH/a8c7Lto8+wXI
6gHhKvPaToR72KMqa6neKewDvN9vGl+MO0HIT2spzFvXb65iXXb7793KXsjE8Wyq
evVzsumvWoLtqtuR8KLx2oO7Z3e0bCxN/rWaqvDy2/HpUP2HlR2lw6XjyzXQfX1c
1brcIzdGXSbIRdRqQ65v/q1id1UJqMZ+HE0QkZOwvn2VKzG8hZ+OIO2vcjf1XRZN
Ae63M9q5hjNi5uMZ/oVitSUMB9BfpcGte+z7eHM1LNSRIslxkc1mwp3oSFmn+Kok
aIE6+vZAfAJtDVz8a9VWSvi7NEtrMVrUs/X5p+c93Ajvj4xDWH3eyE/tijEE5RCK
XSIrHf3rpbje6NE0wZd4rnBCJF2zfqzwNlAIrQ6zrZTbImtA9fubicSnPJKywUm7
17uJzClzpS0yGEnG2c5yI4zFVntbMw31Qtkz8mQq7rRKD4iW3c3eg8QwF0WVCEIf
PS6Ek656sDcVAnvWhQz2dzmgHrUdy2cuPGXBh3BkbifK0R9pqNt8WdP8cQcm4ga/
gcqV9HRHhCCexV5bKb+/lsfufU5q9FHSG2MvwyeWH5Go4MT1VpoVdJaopLJXw7bi
uxJ/TayxApdyA74jvluS0D3MVWIpzLgoUZAIjWhAEVkxjdOSoC8VV7sh6J6O3FJo
gO1H84wU6OKplJ3FzfpB2I2CwT3jZYzSzvbQozakcQ+wzMEmw+PcAuKE736/330s
fqLV866KOGCjUO/uIiDDdwFpy2xDbjRkHYQdOjz4O3Cy4jWoA+J/NNbPoGT5TNJk
yEGnJ11nDAqsQyGUEQiWdf6Tk4SzKHrM/kz4XUWxkSmpfRw6GHzOaB1+Yebzblye
qpEBf6L7zzR3iiJZArcVebREPPk2jlXtqp+gHGKMs+Z/okH4RcUYie5ZOQD85Kem
h6+iTzg6cuLzn6hQbsJlD+8JJOZ/lp18VusjH9/bgBC/gBqRVCH00ER72nEQew0T
F96HUTBu5LWuC7VjoB7QQLUNIrxzb86tAfitSpDfZ13MNldXuLO+XIglTZyNXoO0
MjFhcO5D/tvCqwyk6u0/tUhzmLei3bD8cLYJGzLpZu6BQDRt95uBLfjT2SCgF4Q+
iEFn6Yf5fOmNWTQG+f1LXWNdNL9/4PVR7lCWpNwpaMZR0gufe/ld+VAGgSMhmZ5z
l/yXLjCwox+M/7e6Le9/dYfA/e2TGy8FQOZ3/kz/D6WP/NfHXC2MGcj1BIc4jyR9
+lYBDr+v7FKNEkWWa+IyJoZ0Cj1aTq1RRIF3Swkg49lELzECy8OMXdkbeJWDK/q/
/x/qDpVzhlwVVZhfRGeL48IHmVtszYIqn1TPavfnCM1QaBUMnwlm1k+A1fGxggOt
msMEN4R+WSCjg5i6ig6kga8zNj1RGh0AWGXnTYSa98yLk6fsVkEE8nlKoK09GcZk
PKeIZlkaCOfe+XYSHqxbl1GIwa4XImNY3FeBQzpZ6WsXxepy6c+pSoWNJBJ/dTLN
hECEIYmJur/6hmx2/buOPMVAM3OgyWQwZdoV0OL1X5QfG7nD7b+ZuY3CEs6lGpVr
WO+q4XKRMmulr+tsIWIJBj3833YFyOX7dd/YwZbDpNK0+OySYz/h/GFnY87XEZAS
WwQ6U6FUsN2BRyfmNRv+a5dgpK2XWWHCZOI9SCzNhxKT3xffmSKtMDcwTSHbSU0+
0qtksNz+8wZWoiski12Q/EW+HHx7D7QhFkYxjeR6ZVDsp+EkfQyuGcVUOgV+TY84
Rcet4MeY545+omjk1QwuX2h9PYSN51c8l05JZGWmgxpJ73rpxT+kbIN7FZeQCN5f
a/zepTCdlav/X0d/sEtlskmZ8RfTTUGzTfynxPnI3n7XccJkeWRunDT2TUPxO+pJ
cUP830Qmhg2OWKyLP3kF3KSpE442OpoQMEGhVMEwVzhMZRmfVVTr3ODeiKZHBlUj
YTffoCQHcYwPV1v5zFpeJGBT9HcG8x+j30DIrQGUkcjU9cue7pRab+jkdgCqHncD
Tg4JY+IvIKg179R4XW1pF50wEgRGpahk7/O/DXAfdBOowVnjhH1IWwXn4F314t8B
kBkRrGSk6i+CCzPiYJvz3bpvW89v009lb9S4dy+fgHWVAbOTrupXnVO8hP78c67V
wWB1L2Yra8CSlMbYL1hLFCh5j7Mscc9sxjt5M+ggBP8n1Cdc4jViUEShANLAMih6
u4n4afn8xtnQwfJAJxt//qR9nlqPdOyTqtWqtSsxUJBYFf5MMpdBLM7h6WE8i4gI
AV9F2k0WReUbuaT/lQCRo2j6USR4ppbHuCp4XvAdOlIvvI8/Xe16KWMqLuY+pAox
SAJq2cRuWhdtYuvbmyRhlfjp0MWpxtRVOPq3HLObPcoy4yQ+B0/4dzruYiiB/evy
lQvr9rabUxkghCvc+hw/UAZrQ8ZbqTSWKq6H5tQEgAt0jPiE72b2Tr6flxKpMr3t
DA253mKBe4mlwQK1GiLO1ISCdkcFPXNoEVifZgOvcMJVGoiSv/nMUOGhl6j3aUGm
0sEd/alxijBRdUxTr1sLolvjkwzXmnIBiQV8UEz8yjOI8jXxoz9okc8BXcQfkWVZ
zpYMtXcLDyZoAYNnYmXWj43gkQyY2w2anBjgymd9hxcNA1z9kAx2BvzdhVS4KhBm
pg2rwV9gwAuZNeTPlxqw0EIJdgtl5VdeRhSVEiLy9aTdtjz1DGItvyLpChJ2Exg3
kcxKazn48HYJ3PZnuiQQjTDjlVw+nN4ukDr/zQp8YVlnDAUD9KPBUxBZKzrdSz60
GwTn7BfS1OVWuAmOVQSr3ezV7CgMZA2meVDalwjEes2o/Bv36L3eH4kSlp5mDO9p
qB7sjpc9yD5PflyFUtdvefHtmPejT4RLPRS9qzvY6xVcvt1mtmKPB5a1ng4kMWQl
Q3DaJKtjBR5ZTvOub/1WLYhi62NsHN1ZrXjnQcw10LWK3vEw9dexc9JttRIA0bLL
hVZ5rI0tJIliBjMPhHSTm0lyN43fLhHvxrcrLz5Dp6KQXcQKq02B+IWC/SvlguMv
KvG2NEjF0I50DdJoPU4wZOdfqUNL4j4AvK9aLumQB6HhDT58MCU1FG3FCOrN5BLB
T6VbsQukiB31Btc7lRWws09vh2PlG86nSxoH9yYOaNrHJZN//hKeeDpV62ntvRtN
2FF+kLp3fNo5dIS6MnWZewEB76ZY7hixCNSfhq7ogyFcSYkQ030KOQ6oVh/fA4CV
RH6i6qVeN3KPlxH+1eIkNeGDpDa9dB3O1AOIXamNi7qITauQv3bxscb0eBik/T4N
fME9puseEaN1YRQdFAE4qEGlTXy/p3+g2EmGfPHh18/HR4fjuCjdgw41gECKo19b
vFaVl2no3SR33oyFPyZPlHSOr8kvwCcqzRX2jVCHt35OtVgQz2IPfVt0lk/k/h7q
0XcWli9yuQei7uioMY1IJMgxJ/YAzCXYovhVWRkesxUvAMZFxdALffF8+BgA52as
ZTlfM0d0UNpXoCTtIk5n4BB2eV/LV3t5b7StWAOSQyNBq7q3harQjDRFn//NhIwu
AMnUpxCrCi5Mshngi+mZyLIMi1pOk00TOTKeVTPsTbbiUBvvNK55zGmoosyehVdf
spjq4plrKcQ49HmNzwAzmTo4KAVmy9DI6l2P8+p9kPRFZa1jkLjkwG0FuFtUdj27
jsWJgFsL/cqajA8BawmsC1vgOE6fkrw1hHpRh/+rVNP3IRS3wjxmGJO4q76rDVGj
IYDEwMdLR39xxRsz3+YzCHC0mC8PYcSDKBYV44zgylLCXJnkMp9hGnuIYoGuvAg4
iP2xjN3A8cIl4WN4icuzYY5TlJNK0IVQnO5LBDU8urXJr73WT9y1G086sJsQKSC0
AYek+APk8uDlkbw3GQeFOFYc2r4a3aKJOge5adKfDgTSZZADu5tycRMT79tSnP3j
uCby98sePz0lZ+NMLfRA8w+DPva2+yIkIk1HifEMgzA7nFjBy41nQA9Kk5jFmf/7
Vl+4QkIrfa1peGqft7GmuYYGCSoa5a23/NP6aGjZyXbheExnn2UbC0V9f5+XcWa2
pVCsU6OdIZOzNmFiNbtQFvabFJJoHSRGjUMlO1t9cS/DBnchV8dkVR53MFtTZQ8S
l7IWffVvb1EPmtswSENrkMUdflgQQ5nrlI36nfx7bA4XI5s21dvClQYxF3BHowOL
5fY5St2NOPAleecAm8nDaug16l2G4/6bJ7ImqPjWnzrXPKiza/ovvbXw41wBS67E
TuYvYsgl6zPpDxorUij9GQwSpr+0e4PDhVuAdNR4URNDZlUoGkjgiRgBjJ75VcYC
OY8+qTORu6SJY7AvxEUGDhG8Mx6G5kUSrQk2dZr6uC3fOkFEfF4B7dZA4SoWZ9E+
FwEbaJUjzNGQknoltFeo1tIQfui1y4v+KF2JPnYogzAKLXuBexG0kHdbr4HdpIx4
l049UiVLjFahK2B0g5XNG3qMzD8pzSbhfqhOq4yC/Ke4b2ix76+8eaIt2H9AayfP
lE5LpRYaEQjX8xQB+ONkXzdC1KXKxd7QKc3hCVTKsIRjfOq7prdVeifUIVVC1AE6
P6+XvSSr/EdVo7omM8gVh6ph1v/k6Yz9Rjgga5wTQU3UgRVKZw7d34yduTs2dEy0
V/oWxMkEz4yntXTQSjEX89KX0XnLnmjZT1QffB36ipuq1x5hM/c7qel693F+3rcO
TxUmXR4hKklxEn1JKQrTGMTfthTvwutlazBdEixBvdmqISjv2U5jEhurMEvBXJ2j
gdOL0RG0Yu61tR7aGCp0rBzCEvJ9XU/P786sG0KmuEaSKtoPyQ72lngCDGVEpDk/
/b+VDOl4OR2fZ3zIvw1g3STn7XYwPDBH6oCv9mQAUPdLSAK6fHrWQ+Pf8E45rd/5
TVhcvSQATFnwn2s7+TfvbLL+/RZAVa2RKqGU3eQ/U7Iz6WMM/eJrM7ThUpfJ70Uj
mDQCoAUYfb2Fw6sR6SrE+y3vpUprVT09ZlfucgPsG6HPcEnCkHhSlcXv+/6K+arg
i6huQqfZNBr+lhKR27G8xDetQGQD8Ei4QabT7ejqH3AG63kOdtayEdRzhZk/mvVT
0l4j3kPU1EnVCVlNVShGPHXwdv+4Z8r4Mp4MWSdW1uX7eVzbQKVtHsH0ZhTrijkm
655tFr6T0xRWOfoxM8ZAbbqFADATuHTb3AhQokdHMDVKF4JBJma1kDC9mYaW5cT5
pDKCsyH79YGWbENQEvrdgf6YNH8DDljevntdqFSUB7OyOtMRpm/v5NAnwJaLvoD2
V7LZbpO3LyKwRybyg1QiMcBoT3627J8gWzCohAhV8oeGM41l4HE0QweT8hdotwnE
EIZLjc/zq8iv+nE1LZ5ywAM6J5M7KzN5+XenNECfZ4TE5r9tDcRwGPFkDJZ9pCmA
O4hiWq1WcE80RjIM5kHfIjg/+GJGzO+Wzhak8VAxu9hCbC1fBYQcqK6lAOiye6MP
Vi0+9BlK8uvQHIku0wyZ6Wkb5GBC9HV6BbwOkdBIAqJgxoGkKCMFhXU9StLtXymM
bcytsBCMZa8fSMq5GFsfkHmbIF9tPeYlsSOCy9OmH7YzVwI3NtH7Px/+/aEYOT1I
lj8Zp8ieYtIKLbqPlGL8pDt37NH5jUgmO3HhQDdvKPYWgb/eemIX/H/lYJMjOe3N
MP/Y/9jlokSY0E6xhtu/KS0v0QwQUpTBX4+ihZT4hvJLjoa1asBKSO82ZG7cfrxY
moU/rgT8VAsMfwcA5cqLP5UCVHIs2xtDoIamqYVL4MTFDdriWis0l2KRV+h9Ode5
bCCAfu3Z734Wcn2Rt3pZvJnmtnH+6sT2t0xeXsbo4KE2t8NF6L1G9tAAg9qi0+f8
6EpLSgo8zecXcP3b6OIV70+Gh68JDW7C/S1hv3+Jx6gRA8v4V9i1QhRpY9tzp5Rj
5lMb74StklzzzLk80AdDItoEg74ysG8lZG41ZDjx4+DDxfvtsnxvWXk/3XuNo63D
gKDeNLduuQhzHgqwnRLr8LndGHwEAyopypnrh6hDXqabcffJOMr8dDy13h0x+p6d
EdQ/O7YGJoD1sC3d/8CfEZhcicF2KRk3E2ITGgKnpmNnNwKl2MXYtql8oFM+/AEz
3tDDJLEQ3pIG1SjLlsHv+iSIWtQxsT7/CkRasgUVK3zDfFCqEK0uu6paLswgY0Te
avT+02ojvjLd/T4C3oYwnmQCu4AIYyqHUaLaX0JkDCU6PiKjbiS32Z7TmLIe8/5+
2mawjjuuQXvpSKpyKe/Uu0XJ+oxOBEIJ48B9KgCepX/m1Vi+DeREpWgPTz3C6kKX
vww4uA1AvcjbBp44BPg3T/55TItsf21LHsoenf2ip7NDh5PXmtCupvD+pWlHKQeJ
1PubcdYTZhTQygSIWM9DtZGTW/cMknz7HZjkmRH78RM/+NPK9X330IvvBPh7AaWv
5tzkFjA22ODbn8s8VUIdmBsURpOkl9NHMBI224i2RwNloxtxLBzsaUD2Eoj29Lbe
mCzzx8E8pU08RXNYGREBBNG44wykS3lYd5RW9SjDLGVb67ZDBB0tt/z6W2ru/O8e
YIDErC4wezb5xr3Ij/uOlDymgS/LF1SS9X2HR3JQfbVXjnAwTwHmh3O3CXM10e6n
J9NToyIlv7KwCzOCTCyC8EMyOrc92Bl+QFECosH/sKE+bM/frYxBiXIJdET1GJ7w
tjnMLjBh/0slT9vxUVDfJrNycJiA3eZl4+45HCBCJTuQW0XcJdTCJyUjD5/7y3gG
TNQ5GCZhvx1UXRl1dtGWrm2ml0Stn0bN6e7nUNcePOwUon/igA+CIgApkoBVwpaq
xuEQgwH99BDhu+huSErXUeaRRUug721IoKiNyMt5XuyurU8Dz1FY2QmHtFsvaCDf
AqEsQJmfwzTPHxaoW4xDam5rdjc2QUTFdPnKPVzx6nftVWqLAyHvVcEzhYgjYcAc
Ox3t02wntPYkU6Mi8+ZGm2GX3mM0mZZxk0tIbZoXtownO6tBC9lEZFcu/+53IexA
k6xXgJuV53lDWjMx2u0y+DNaFj+cB7uuqJws3R3vqOFtedn3C1vHPkm7wlW3ez6c
nKa/6V2VrmTkQdMVF1kwQ2sEgMKk4VWzWhyKKs1qKlJrMBWBTCWUPDSL3Ch0c1md
Z6RgG8IRzqvASWPHGXXxcs/nOgdjBVAmGSYJy0Mf/0dM4MDcKVvpO5vPdG4+G3Lt
H4yhghRyYKI0ZmUvdEhAebK1Yh6sePPJonZeo9elw4hAzHf7Guhp8/dccFYOFicM
3pm9heH8RHx/az/OPMrPT/lYArN5jEslE7dZ2sCltL995gLWonTKTU9ZLfgAdCXe
kniXA/+ENxcO53t1gJxM4+oo3pZadHL5dtTp0WB7Gzilt+h4jVaWFvNw2E73bABO
dJG2iXdYC75kv7fJBliY5xF8K4Rdd0aUISKYksNDoxWlpzMwVFPBiV6jz3E8DcBm
2QYvdczshfSmeEOTecdhcctzpQTSbKEqCYjwakMImwqViE+U3BMijBo1fYMP+3GU
YYLeuN1d8rMGJ7RFS4lRdCAa+cnaXI+4W4sChZ5LygDKqNoZggyEQFKkk8TKvAt3
+MnYxJ4Da1gZNjVydYK8MtqMra58grHU5MqJTHfoCGHR078XxGPHycpus/9m6Dog
gAQrXs6+vv1Sj6rwliMJe4uJY0bugatPfO2y5NWL/l2uaivKzaDnpWvDOTxVv+rr
Px6TGGQ/yCDzboMWwy2iC6fJlR/5pn07c690DbiVo0ijyCxO09NYMG3QSV/tORHp
Vbs8OoUfr3uRToTCaoIEFxs/jH8mJUp8P8VShd6juejW8vFrxEtyUfm3QH+BOPTs
nUvj1aYmdcaWXAt+aWwrOKiSS+l9FZRMkF9oCkk600u8fpS4fSjNz8lTDS9bnmH4
bMnereezVAE5IkDLtkLzmbYxHsrRc9SlKT6ypErljJx1mvJYcpr+iASLCFEIPjFt
7Z2SvS9K+d1QzsbZdyJJIhqNNF7YY0Dyv3g7Oi565m81HaJrK72QOB68duXruHms
B2LTcdQzedO6AiPwaXMx3n8xfJIhQjjdMp6qq478ne7E4NyfSxI4eJ/L4xorbk0b
VcQ58zlj5S45njB14IFJ463lANiyz9vkuEkCuezi6JxnJWsT2bBvrPdTAfgDG6Qc
O+eONo8kQagxR1fB6Z6GhVfsCxFmHlsqqm7G09ToUCSCRtXAKdO1Q5xKZ7F2vHyq
59qMdzP/vgn6mGFI4ULsqakWYB6aWHAIyd3cA5aM9JqaECXSsZ7q/074dMxunXHl
HGFPvB+L3PrjqFa6wG/2Pv/auENT7e7NQ5bv60xWcndWue0iTsd1YTfKBBXOBdoL
zGlJ2nsSnP3eZ3WNN/p9A550XHoXT0yBR2vSMGfcppooTJzPnIfDedOB3H92bE3y
M46WhkDFykcxEyo4zGcLhNvmflYkBI5c23Z0PPLh38Ahbfda3fJgZsdRds9bd2LB
R//9fbxm/vhcBodzI0w7iqYW6ZTjsbZWcAjQdo2NkPlpmXSnVArPTvIHoIznSrqo
O2hN55YzcSjPs8GhnMrVewlqEBMMIc7UZiKEzGN4YuXMWvq9fL4wvS8HxSi3xDyy
ANspZzA5Z7gjrLa+7wZCuCktpKLbAFsBm3jp4VbYMSTQba7kkvGgE00tooeGKrfv
XLQih1QeBildajhxvTEXOOe1V9br5CqqTnYLAYat2hp0umlwCN020WfjP4UKudFu
4TD26+eWlLwOkM3IV1SOeLxEpEllGszs5A6Lmv8K8iuNWGl+WcPlF/LyPflzFtZa
izgcyKmhhOjEKt0psQO5kws0WG/adYn7CjYFVwcIsE/SCpRI37/gYlUTApdrGBk+
p+E/EY47DrU3gLVEXcFgRXDvOlDHap8KzyjGllo0pHQNpe7H0PAlK4paL5ZR+oDG
uJGwyWAS/SK0Ld9dpt7gfJqwrpyOPqEIt/g1xq0W7esxSMs2JF9/qodjEyvdZVT7
yNN4MqZmS4lUybqBhJtzJugFxgl0oANGbFuiBJfeyeB03wMKFFV2PsTMm36SsVZw
7zkY3mlIsmS/WJJR5OJl2mSalzpGgdrliRQ4FVwbEQJRowhwV0SoKRiJ90Ppfk2Q
/uBfWLPznfi9wUi9HODp/7wfSVlze0iawdsf+jcl7vNdRSH9ex+ELwSNG6+cmUdj
dhvj01VyOx6QX7z7m1K880OQxFq+XgoQ0VZDIA+p+5VJro4Pc/xFHTdPBnOmVwyN
jDRY+xteHD2TS+pCQWjys+ddyL7SY5C5n2sie9w/jmIsq9dWVlSXD55NdF+kI5mL
riw15KPLuCvvG1P4z77mr7tvWGqjXhrGokyOSg6qwg8Hm4my79myOtiYe2gBhpug
/NL0tT5OcvnTMbI4OndV1UyAstN0hxDAEBWrbV5wScDnYsqWss+0YScxPX60H4av
LunqllkHms6rJbd4QFeY+Gjl+PCz0/Uv9F5XZYIDg9C+KsdLk+4Wf6pEqLyTz8ve
KMDMQ4JN7C1ney8APlSu28J8FioYTMxdHDIL2WLCJ6DbettMrqvS6wveOIFXxgNt
eMatfQqazFz8Dxiff/oil15FNehi+p+/yWNyFnMN/Y83mr6rBGq8MVpZxiSgpm5E
pRjFjq4oDDzj3wlIYeVdFGheBBaswWPdC31z6qWv++5O+qEhnfxG7ua//FpJmKIw
5uvThcsYLvs/oeFlq9ZH5pQDLpcgCvJhOVrbaPEiz7TJ4rl1bzEJX5tguZancXq5
KeS/vmdhVYguOvga63jc024lTJOmlZQKzEPzPVL9ABgEOyZHNINHT4RDNk4gSZ9F
NJyUHFpDsDJUYZCQM0PEtoeD4DQ2yRwEXffpuLDMqwe7v0SaVNerRZ/hp6/Rp+YM
XyjM+TrnlAjDdG2TGK6fkLYOtRroLxTbHrUKll3C1pX/MfesAjTnbx9RZj5Z5A1L
WmH5PYpNGZpIOsvAIdBt8poiG7cOos9LJQaK1UfbkGeAZN2e/WZ6eRMG2pXyCZ5z
vxwdhMxGJw3slPhwRxbDMbzS9AbpPtVt4xxOgX2IhydKqKk3YYpThGLT1iGc+h1M
1+vQ8xRIXG3sS8ctDuap+QJ2E/zgp7GoxUOKm0mixOZHapFPoA64i3bgeH3ESSyU
KSSNsjsyGUSIAKIeT7FQ1Cy2Nr0rfCDdvAjlGc57s6S2498P64da6JLLOskkvNNR
CD/6gYflD4fDs/G06Z5ZSlukVAovT2iRHdT2oE1cecUXX03QfqSAKtP1GUaH5j9C
ddEyzB7/iDPXZZ1FuMY9iIHbDh+2bM5syI0nIss1DDqayxrzo6qIR8SbfMB+Je7e
VGrA96t1mea2fT9P7eeOIBq+BmNZoOEWC6D00p50M5ytQjZTnKgSahuSeEU4HsWI
O335agmUeFjoGNI2lx7asY/wTl/5lfU7gkOSuL/4kGSzNXMB/g7fBX4QayVkGZ/i
J7FDQ4sjaihHR3eMt/KoToUv4AlWOYJljeJ/MCHCFti4CFjT+UEfKYMHOLbYvdgi
vAn62qp18Ld9bhx+0G7W16yBvtgKkqZvHtTPeF+PPCnMUQJ0UFNM9Iz0PdH+DHl7
bUs7LOdpZWFxtUsK/vp72mgP2+puk6IAhS0v1HIe+e+x88ci7X6KJZjBF6t/1c0Q
ZSvB+6OCWx3fPTztsjuDotjxQD2Q5jcj+QXo8ttrQU/gH5WMVfXrhfLSHq3LyPmW
RFdz6HawNQua9r/HOd7smTJ6hEO4irGegRxdYQ4qiGCrBkLEF+DKDuyLGbWXcMSn
HrmtVtxKXyDr79ca1j7xRXKfq+s23iuNXWf62hW8vP1B5+ZkhPVLcHKjNLR3tfsm
6FyesImiK98r1m7J3FEWFMpjHFQBrAVF9bMnS+jMRb4cfConpub/kz0beq+WUowh
ZySYwuZrMjWKtj/zaj39hsCZRDM1rfjISPwZ8ttlu7MaTXZk875kjmsMjYtu7yLj
rVqzNstgu9ZLI6janokQNM4SVI8yLDtCSJ7KPFsdpyotENnJKz82FkzHXjA77z0d
Lm/QuYVu3lj8b9vnwgqnTV6C3DAePiApmbgm4rxQCbzX8YFePEo2BQxb3r2uaRH/
D3xJ3bKMbGENixB/7jWkXiLQqHXsp+/G31auyQB3a2utw5OECS3Vdjx20Cn8Ln7h
8UjQOdOvvdKM4stI4qPgMsPxX7hewisPYRI9KfsiUtBGIm6mqlLInEb6VICNP65C
wUqwo9MqEWAro42fiHJXYiiYC6uGN4BaSkYxNhpZ26tEWT9TMxjsIAoYFKi5R2cx
q6c1KH+VpODjf4FjnuLPxi/fXHgyLenlC+zBK32fi5Ttf4GPpljPzJP3tzPzd3Ij
ffo83IAAVxzihd3Yc5ksKPIZX33D8cFPGefNRxX8T2Z0wxXUmABAghhraagvWebE
efJueHHwLySQ7FdW9/zqt+tuaXdZJcW6FaVgQKebrd3kmRseIisxcQY7jf3MzqIL
TX742Bnp4KuVVLSTPkZUtIor0G0IJFt5QnteR+rvgtYVe2paUS7S8Hutmwc2jtf0
JL67QIJVvNcGsLtxfeVPUrlMBw6jOQ9OyWRTjRLGfqT3QWTnuI+yEOmw9dKqZF0c
MrVK04PyTBskRbvCR57yLzXfKwLXG/Pkp6Nfbv4eT8XXK6pcenRd4phU93THAzhc
VKP5okfuOIQSPt4Kwccg9RU6rrToy0jYldutlLZMuEwk2WyZwKTP4+OZjwM2yA3d
jl7PDfHIUQxojQM0GElkticLtHYpuSDLgTkmzIabX+olL4OjopiNqSddWQmpfPwH
Q1Y2T07GHAetpi544ASEaobErW8A/djUFBmvC3gb2kLqg9v9TE7UYOmSdC62v/DC
sXovfxUMlIa+RUsxxeMFBcGF0dohZlMiZl1wI0xggeqU+KmxFkeLQMXuoGpHRAUQ
QNjv22x7SeLV9ZuwqM0FCqZKk2BP0x4kiz7/3q+KXo+xDgyivbJLkqEuBvF8k8el
l3tPBaLgA9NVElNrmd1VZ0M8eJpqcpp0I9H0C+XK5ap0rnd5EPQVWBT+88zJvu9J
tDtwR+2T4Sq4DdMB/IhbLBLa6tvfqouKz1zMSVP+ZFMV0HKeqrIh2b4IaAU2o3N5
2yVoO111nvaFo3V7uHS8Qi0l8KPB8iTrKmKu60Jz8JiPchTt6UgyEhc7MS6mp8XZ
5CxcJmyRg0CwF1jmhS9jXchWmKwNbv4pdfjL9m4bDLzuRwBUyGZtsk6nya59oGU7
p3gzCRsIIhSSSsQIQtM5NDD16Bh/vu7olsSJvmZkjs+JE6+XmjWro8KI1mZDhrKL
FUo0/KUHp5tHR/Iln8kBOXoIowCaJYnjObxhedrV1lzka5bCssCwJgfEGm/Tl/bO
GzbiIO5cIGk7b/h/6Yt9LKB/Mr/MqbK+DUwdloch2huqySfM9YSoawPLSlEVB+QL
dKPrOasq2zEB21FL3VnGyVkmkuTOGb/34uMcZpuoSBfY0Qrre7xrHs5LVXYDodkL
QZ02q+yc6Wr3cj0xfk3zVHdjIuUYnNcSny6YoDF/INvg7RiqTjCHzndXxl5HTSSL
KkVWLrrLKnrYa1v+fXRTNIa7jINIrVODwxIawEPknJ9aX1nywFMaE5npH1ZruWBr
P1Qf5ZcIjb+xczuJBLAuxQCs8usHdjEkzjF6zXi9dgGNqQWttVpWdKshadIjthwm
0zKSpv+7t2c1YiIlrkQDP8+E1j3HUZX5+dBzTPLaEULgR4KU+SvO3975xCMDQ4+I
gLKeVfClkAdOIGTpGNo8Cbvnciba3xZFV1dkOctT6sluhFe4Lbn6Pm+h/63uTt0r
e0dWxDpN0KOOfRJ06+hj9wxDWi967H0KcjuNQwYlxPZZjr4TBFbt1evlIfazAbKr
LbuVVMMnRsqMSZxLTdOlnWbjADCFBD8uF7K7yCjxgh8SMisoSB/99gX8JvDGOOJU
TTaQ6TkBGYGyJ1PQ2Z6crMVUUj5S9e2OD/3tC2dovDvxXtezUtgCUjiGJxZ09Ivj
gbhkNj/UJomeiwtEUQHloByJf86vdIljQgFq2/xSP9QxYbLqkZlxESQ9MZmHeC8W
HwKen992QTkJ8YBkLwbfqILY8M6UArWaH99lL7plX+wDJnKlQhKx4A+3vP16d9Pa
oyti5pZYybLBGw5VdFeCYqDJw7PVsnGYfxU0AUOhzNKbOL/z63syvNAL2oTKRFCv
DTuFEzVayc97MaerYrfxjxfKGFamBfcZmvMNyA8kAbH3O78pqfSqcj0tjCLyP3/j
eR/qXNh/1vfYMccT3T7KGsyKJsLSOHt6YV07FRz/LY0hK7QBnYZeQ7E4l3mgSSp7
JyVpsJudiIcLouiSugStYTtFGsBlQ9lB365Pr9nU9ZrOutIwDGO63ERmpE7gp7f4
xGyk+1o48Gg94dVW7Hij09st2I2/wK3IHmtLH1UPQQRPfzRDeuyiD/BjgC9FEnFY
zdBV33RKOvunwQXt2DmxJYn359jbRoOxFVksQdH8+4k/S3seIa9Z1mOAlCl9L2gg
585ohCYJWhqHc6aSPxSm9BCh0CFD6C912FAGvuJUZvTc+ns5WYTt2140aJXXlCET
XBCMgvxkiY8mX3T6gz18m2mmsOApFaK0JZ+9MZwNA19uUyNPFfgXuwGYcaluKmaC
tHzYD33lynNr4X1eGVwSudEGFxLkERJISGHGzbbj/H2WLNnarhzJPJ3xcn9Ji1UQ
VuImPBEOXeuqqSX22PfGZl4WSg+FSRsHoVRsIZGKoxjFHwgx1nsu0/D2PPndi82e
NFFv2V9uZFJYKi7tVC/1z3Z2dn0WFlNNhM2gffdbuEo+GO7EuutAgR1yBIKPp8JU
uPAm8HkBwjZI9ybtile31byjpfT2Tygcq6YFnS1mWbemvh1pKHm4mKYRratIwuBl
N18txhhDjSyL4/h4vZ2qOcV0GbHsw8FQm5LfeiR7L7ysJoe0/3H4p4C/zTsVGNjz
JlFzQPJdei7b84DNTGwC9F4eCsx1N0Pa/ojrozr/ibjw+fotjbawUDqRaFSrESbV
ZeINWQ3VM3hJaBJUbFsVcIb5b3AE8B99IkspDkLkk3iNrZGZ1nlM5jJMHHV6VHmW
nN1hPrWJ4NiSaxDMtKQGgkU8Ju0wjbctUUhe3Ppc0+VoUwhhnesUG1MJ7H1dQ2Rk
ToKvu+0Wk8qHa5H2RSGRgWozSVnYBbwtpBwfsM6IZtrpbWdL2CMaMw+RA1kwIPq+
JTCK9Zgkat5s38MDCcIV4aR912PbRuruati+kLDmkUBdZZ0hsS3MBahmJyyglzYI
DS+i2A/tCqooH7tkPJJLAFE2qKHfRXKnmrjmu2x8e+u9zxepGrUHCPLDyU+CYDiv
0IxjUtSjJh5+AYjc7KkNV4thYAuNl0RRT1rwHmjC3Ytjd9+mf06aHNKDv7gj+pXb
8DYQNk53U5JeFCPRd2tnDg5mbRfy5QC1nO6oaTaUUEXHqNC6gEr7kh3fKcY/vU9y
4tdbE0mbgZahq4/McdHPZppc0lBQoa3w5qNoAElCTNsMpU3hG9sPB06fsOumbNNj
tzsMiivRo4MGGEDF3lAqaHKby4TpKQs4JBwkGHRcxZzOQUhyaxRj/dU+Zv4//voW
L79n/GibdN54ySMq8nzGs1pXCZpMRiYlE3FgRxzS4TEnMUtHfee5FwYLdGpMcpkr
8p4HYxuOXtsMs8/+rqmctRUb74xnQGI//ZmFw6NXGgU2MO0bB4bQok5Tz/p4kYVI
rvaxbuuxaI+5VkUPXLI3drSiw5kDi1WGfodUTo1y+QiTcEdQrEUIxFPxJtDSb+CH
HTXV7Zwv9DYqmLuQKgiCccW8cWJ/OTEQLj30Y6bqxlZAzvsuwvQO+vsalVWIENTT
qNyVEKuUVzGfZSOjaftCphFyPWkb8wRP3M0poqKjEgvui4rhFBjVWWlPUbqVkBJY
JFncf6x3g8oisxAwM8MXms9dlRgB3+Cp2hkVNFoI0vtv3iAkUvLqZ0NdH4EMr3/Q
bYo8xhX/lr2zvcpjKJHF+VE0PmT8ElBiVcjChObGbsH0iMBmw0I6aaeb1V06pNsm
sAWOPWSC/afeiFAq9CnlFfNii+ZNE6XfSRCRNavr9X+ELdmRj5O+WuYnZcwYrTJK
K9/rznSjhNfV4l7w6/gMCUwI8XMrmvHUMDxYGefWu3/tV/9HZhmlXUFuIZw+GHVI
VEgOc5OlMRSmLfnPxlgLG5CL41UV0FHgRMhYfAehWJVMZn5Vy1eYmjjMCMUNLM7t
nyPPKs9tYQOUaHE1HYK8JXfeLu2n51mvfGVF8/PgptB5dxp521dUTjSbg42V3q+p
tIzTXkMRsvAFy3m6774ooXkr/fUfz5VZTADwIGHhux+BtKy9F/bzJ/ePkf+rukKx
IXP3qvone31L5t2wY5fBBwSTYEqLL/pZTm5y0jle/GJLsU78k1qlLFPY0hqZBuiD
VXyNiOgziLCMRA7Fd0IHJV7FfqMhK8jNVr7omNruY4MBQjnBwo6Kz6YGn/Qx6PFz
D9zegvVTBsjHXFmTIKWCMfgNOFvqhlqElxn2kXCfupEjkeh7K4f7M+boQprp/qzs
CNTpqHBVcoS1owFgnN6jA/Uekbo1a9LlzBtJJ0XaU0WnULLIo9nOoWj9M0YLo53c
tuEBB5SQMs/8wgfjiYLZ3HEq471mXfqQbGBjwoISn1qguQQbtsIFLNVjq21c5cJZ
FZ+Zth+UOOhzMyoy9zUXihK6PiyXLuAqf9ckxh39V1arH53HE/TUWGwuqhvDEggL
SoWssBM4ieT+N6CgrAHKZ5mVlBXiAlj/8xxEuJaY7vf11lf2/glwGCY1VGR5x4FJ
idz8y5ALh/CxQyeBFI+HkfFzJBYy+UtNTqpvPjzo/+gGi9QCDNodPWBnsNxn5Dp1
XJALy311rFErC8pN9H0TJ1jCPkrhvsySTkQRRTEegafhXIZcpmVzpz+p9Pqh+RNX
VIJ0pAs2Zf+jF/Lyv8W90AgREdONZoxFxT7Y2ulBNChpAc2IZAFUPpcrJW8r/2UN
F8opGt04CS6SpmD70sTpeRi9m504clZ4ktG/uXNmnhAC9QVftmTjBXcDeL2m2ng7
sLg72ldwPnKT4oOAin0K38MrSTL2hXNkJYb2yj0NRx45CRGaIhz05d+yUwjB8fhX
HSwyW9Z66SbXdv3XzSXqCjE5xNBGJhBUaJO4I1av7CGTL0CndBYw0tLOUl37K+WO
+C2vrKvxky2mAf/E25MzNVciPtGGUtznQWq1wKSlg3jLrbrKfeUqJhw+hetuhQcd
x994lvSelS0ln3ZWiKJ/8m8jVzAM7g2En+odezYZgJcywrHDNUckwtaX24pOzWne
xwJsP80p4x4HBlr+GBVy7QdzaKDNogRPq1esr+//Kix5GZaGXqDCxmt6GTommqUJ
IZx+q+ZoplFZdUaU7KRq8X1o5dJy+mRcyGZjZmi3TgvOlc5mnXF3wupGbFE99Y3l
IgZt/VRFxUNh9kR0CTqlwyW1arwEz5bF0DW6tOoS4YZYryut1mbH1Yf6Y6QUIqTJ
YWM+DEI4lJnEqJW9t/0vOlq/hc07yZOFJuW8VflZ8u3CizuRyjye8X3dLDhw78pA
uQ3c5f6drJBO0WQdXhuVblc5Ymp1Y2d2233XOXdLbiXwaclDR+vGhyKNjsZlpXFW
S2jKNh2F6OXWhh3tTC9xnDqjHML9iNZJhDLwD0eu9Jl80/IS7TwL20itLF1JpmpW
GcqnxvHtyoJN2KOhB3dw3MWhTrDZVXLllFz9r52cb5Prk5berD6pVTwpY+9K5nHk
Cg0cQbgoYx8LaHnIvvw+xMf+81h+C6gv1HfQ4dy25lbswN00oGyXqbGHBe/kosZQ
b/3tE5CWnQBx06jkhoATmzogJnvDvKrhKJvB6uXcU4HBvCL/UAxkDN58eZbahWIx
FHr6QAHNfFR2Vx2rhVFjOvv1KoJFOUhQLckvYhM3Q0Vyc9HBjMs5XFVzrxL1qQwa
66ptp8cvzkVEzHVip0TxVvMrDzOjKW73sEj8/nA9vmAZrQXU9to6/eo7DRg11XWp
jgoQ11zBzdDXTUIOCxP+sW8aM1+HLbXLK01dCE8uqmFgA7adpELzTzBOjHxmGqC2
XvFJvR09Lkuv73gOGAP2hSyxtl2+XL5NuEpYMutLIn7we7P4U1JPN8VVEUajebNP
UEAoyoav0xHFqFqZPoDd6qUfOzCuEYgbIy9Zp3rqSMm+14pScXgZxZQX51v+qSPU
FCNrcnBv1FLlT3p8d1sNXgQ5p80CNL/hFvfEF6Edm4JG8hPHDCqmnjNVzpg0pwFe
bvuPFUMBdBysOXHM17kxOIPG8MgpHN60Vn0ohjj/Ihhjv8HU7AiPVgc3mN1bf2UM
kiEW24hlZampISLFkSgJPrvL0JmNr7dDgWgT27Jb1nXmdaEa5Uda3f2bPVCwpMmO
lhP3TfPZUA9V8YQ4LsUInp9fuKk558bY+WbEN+gy4m1ffFCzzW/jEJ5NO4MYL7uk
Y+sccN2PSGk20htdiZzAJSDZhWShvy90uGYCIy/aH4cRNnVAy0t4PgQzCPohbd2y
Llxub9G0ug/HGgPCFJ724GWZtZFgUVFp/ChhBBeQePq8TiMfKYyvPXNO+IXWh436
FLtxMHWInaUBUgjVajqdy5I0+CDaOlfPZUjmeQLsMLR+QY6IXnmK8h3y9tVLDVPl
H6N5EMa4m9aKa9+tBTzBYWiXmb6DAHkteGwuymEbB5EvYYajtsaWOr0dyQaMPbKs
05YE+ae3t7MlruaHRGi9nxiQs5vu0ifB0kD7lxEHup3smYq0hH194sU5wc5GZ97y
Ku9dmPvSiceMs2N5QXWZp7zZxHlE6tiAEf6ZNft0O+0jN4A0mE+UJ1Q7rFMPwMFV
JxGXz4JEsvSM/wB2Rf8aVeTyQ4AQVADQW71OoxBTJYfU5e1YDPo18lpHG/4657oX
gAwuV2N97/h/HXoaclJFS+KYM9uAFxa6zrdL8ZyIT7/opzi/rSwLgepzMUbWivsi
QGMQNnpvYzWERu/BnVcOhXmMFEjw+NELNv3/Apz6zhKulMU+oa2tqfnMR+ky9OGY
ga+0RcCJXomSK1C9tEIi/D81lYMGiinMdC2OrLnq6AUzhOQgWuhqR0CobJsQ3pjc
28pF/3K2AIuwwZpjLJuoOCZlU0xeZ/LpIrQreIABEK45+6oRcv58vu15VZ27TOLw
xRurgilMrLXC2/mrFhmR5UpXdRvBnWnGHIgkhE/IrN0B9uegL+B9C6CanpF3D25f
09HwqF158w1y2sXOtR+2pM5dxPUcBPkzphMEhkhiBK7gg6isLyXva0VJBpZN17Uh
5W9r9HAGWNwsU6YVZdCU1P5ifmTpSSktC6CDPzA477a3NRqZcbtX/D+ymqYqloUh
jQnF1CqhVMJ6RoOhDAin9J4U3WWAKttMHjcv9npiyO+tfC/J9NSD0PPcwLtjHXdU
DV9DuYWlZIvvGHj3Bomg0K2J4Vu7uM/cP1AEB9zn99kB9W++x1hAuF4TJhhaibFU
QwfXT2+TLljns6ELbIBsuglqPG5zG/IKmKYUMt2FGEEQgbSvAJv9xUNPQkOGk4qH
qTuNT2C6fy5GJtj7wbJcjDx0aSFldQ5I8HVozgCf1BSHYBeQhwrFumN85xC0v2eB
iE/pk0LMSC4MJBF2l7ejj7yy/xlIqAQHb7FWUYUEHBc4ApwOHGLeWZZxwXlrBZF3
R5py4Ltb3Nh2J++PTNsnySAR8pKqdFNEPLDKwjtWxFAOYP0d7ZAUvmlEoHEQTYIC
xoUoQzDaQWjPiNAsQSs72qCUa6D6M5lKDkCScdzYIio12BB4kEc8+laZlw1tia5m
MsFMMgGMfaaQuwU43xOI3YphQ8y+OQofG1pnegXBD6zMiRclN9+WJdYiYRVdB2zF
8gGc2nzXpo/bL5jlUzzi2nyulNvxyzXDtOHad1x4vr2/dJxgOoO+thMeq7hLNXG/
oAquIkGyihGHmcwbnmXtzZKEt+6wbC9eYj9IJ5ym87SDvguSDWd9CIbFlJLsvjc2
MiUP5FtHk5SQ/AsCFN4UkyxTskTpvFTC2SuUG7HGdyWAuQc2N3LIBDSeIi8XeiZn
PFiLBEb4paQUeSS0r4s9SlxgCmS+ZJ49/DFQ4UmbyAwcVPnDxj2pfIC3dGCwd6oR
DrUuqMNvVO5qhZ9dolwRlPDVLeqG8jtl+oY9Z1WYz5XXaaylYxEavocONV4M/oaA
rD2QVTfX8kTjGjTEWzDBYrgJ86Z80sl4IWCLP3RzRoRmB+5G1lAXweT8t6xujsq7
Up5d/i80Ibj4aYJ5pc/jgQ1BjG4XateWS9WIDj+rM97yDO514vcARXN3gdLCOpzE
T0j1eCyx7KTasQsGbGpNt19dL8cyrdUf8xTVdtRw2DMUqDQxBUKZxq5jHPbS6lpd
115SrLw8foUopuFlnUKq+23xOE/2qQk1wzSzQ2JaLKK0fFg2FDTtY3IuYLj0utgX
/xz8BJs6bdcWs85OYvEN8RSQVUGopmwnrX6u5ulJee2J8S0/do7SXVEkfjXJhUeA
ztaM+fjQAStN9hmZnd9D8n6bIRmIMuVwEPOEsHjdzzwjOFou/VKuAyzaC4bnwHuB
O/2brQVCW8uvPdeGrey76FfL+KGCbR47/8D/VN3YAQ8SPbPueYRBphmvibhXmJst
vQURiQkMlvoGFomYmYkVNC29bbYQ/qLwhhbHLsWw+bY5HXLrVE9kdHlap9iJa0ob
tqiE8crsil4Ei/KPiLY3XEv7vleBjmXQnQrTplBt0wJWrfjff/voSubR4akrY2x9
uIc6qTn9Sb18ndHOGiPSrJKngtuqd+1fwNJRlJUhRF4+QCv2flhXEcfDvfoZmLF5
Iz5WY8xTusogTjZyPjDP80Ara2eJWDdgtUaEF43Cjbtg0Me5hkw+/+NKBogC5Zrp
BUAqepLlFduRGDpT804nKiU54CgXDgRgGVRu6DChmdkuCu/V0Vse/MNN5ZV1IdRj
w2StTbh4fVa3y13oK0M5S0oR4SWY+ijyor+gJRVj1EpEu8kiezugMFbsjVNbKex2
1S1iCyU6XLt0US68NorNLsWVsXXqm53cEEl78/1Va84JaJ8jZnRWsWc6A4OrPnOj
qhMSlUX/uVb+80aS/8MAhK1fM+X6D//ZuV4XOdL/1Q8z6YyfdL7I1JVAi6CLHmFW
cOpSb+5/QuE+zVj5zHmcDZkXCrVQ2KImt6pgEuBTJYcbbR7BYCEYH5vvvOTjrt0g
FggO0St2+og3Gdn3kzPlYH36reXI7vlPrHX1BUHQwaduolWozNhGLd2DF9QXVmw9
FikAXS9DrIKVnBdxtWaRRBM6ixW1kkvnAiyXmLFGeVYFyRXznbSZdTuRifJsPRln
UtS0O0GY13G2zN2wWpyItMo+o0aAwhSXspDVGCpejUtrPL93E2HXcvpwCa18UfVi
BOx0cv69b5Z6Jv+jHw+kAq9WWKtGGlAdX1/3/CS+DlyxLIeMeNZgE/LENS4GZ/YB
bCga0putBnO9b5M9D1li2z51P7vwQVrOAn0ASrgPq2yI0svJX63kcRPqUzlwjdh/
QifFCEwHocDREU+9/T8IEZyxMnGu3WAUtZaqSM8xbTEOdQSl+vzAxPOCN82xQAX4
oBmulueQFRKL30q993LMTrkhv12TrPDrstWc1FyBu1s5qG4JzNL5VXyKeokYfE3I
j4bhpfS0OMPaMszOsvcdVWy+Wk+QpluDabeiqP7+BjHdXnpzmvRmxeqiER8buCot
pwMkR0uNYkqPVHEbZiWPmzT+b592L7IY80ww7fu56q7lsljs4ALbb3Ew8NzLpYrD
96Rozz5LdTsKKGy2lVnR+e7pu8bmlrggTJpBjF+dVIDKauo5jEfXnFyUDFndr1xN
Htfslo0hV6cMgULYE+44FZ5kNL+SHNdK/JElbZPE/oJ8XZSfC3gCDXXtJaRSmhey
uMNNLgFeN+yNmjFoyCPPgbyLzk10i4dFDjRsV6XGlIdM2FA+uPqC1Jz15yAHFOLA
QHkloGEsnGdYU4B0dFqsXNTzpZRAB3OGNEAqe/6pzb2PrJ97t+1q2zOpbYS5AS/e
BKGm+Rw13txo5IxysNFU0YqdKLDdz+U+ykZJ8y2ryPsfod2uzeMEleKlHdfgJfzf
+Wa8nIfT36gg2Fssk+xijF8B2rVdxE+3mRaVrIFWqukA0s7PSDamBtUqXnLsHr+t
S3csql5HxvtTWOCCxyXpmmvL0mhc+EfTgwcG3ExmD03gtPy8aDqK5xbltwWpsJId
+QS/oLFTQEL7/WWOsvIFdE391ag7egSqsGRih491x9QZHWgPmGJSSwi/BHPYJ9H0
5YukRtk5EWoPw2aEQcsqhRhCMJsJUG1R+2PIojsmgCn1BDaDZ8qa5aJ0XEITz/U9
2ajXmzlQjKHyt0SioBPJ1dRws4gSYycbN7v4MUmN94Gyncqz1VamLcHSaT8OOtRO
2adYwcHFEC1iIx5jUP8xSVbwhZYrmRDiEjSjydC9mD3iGhS9HGH5fdEZpCMfuuQt
vZMgfbwvqXs3xgjA9PtKi/AX8IUmxHXGAoYo8UFG5n+NV7uLBdz3dqRce7cxa73k
wQAP1p9dkLAPCKK6xA2CmGqA68Er3gq5+zFBOZGmpWQ2npOJ0KuJJFMFQ/PLEQw4
+U24ax/fbq/FlbmP0FJ8XdjXua0I8+yzpWvl5t+G3ct6TjzHh03WgmNrLRufaYTc
lenbM2pm4/YL2pp2lV+VF5HRDarNgYsOiXzA46SzvJvh78UQUXn5HekyaJhFYMz4
XcJSPlztvZhoQ8Tf9rz9MAWJlj10AvEYRHEljrvyj2u/EUsycHpxJNwc3N2SvpKL
UuH6ULoOGOOUcbipfCDyHQl7maamiE57Mgd0mQbKu6B1pbOtDmEdXfWKRrKd5D2B
SYNJqRabfRuJazoXQviAwM8I3LcFXwK7PjmL6zEEoe7HNjSX/cpDxVAUPfgz9bs3
G/WcNTosEkQSY7XtdDr5HfKGkN3lg0zhSRcihJs6sHHJkEdxeLcfiOm89Z+4Nso4
4LOaA9rY8zrZmK8UlNvuHdpihb0V46rxM8uN5j7CMz6bvH5kODHZmtwJj+ZLjv/4
Tw0089gLjHXrZ33lpUkTWC3CSQF/gUNNMq/4YdtJsnKUJz7zulhEsE84VDsw5UL1
/mz8juuGP3tcmJWYgCnw8Wg+kKKTpCvv9pFi+wkk3CZ7aeUsRZY4+KAfv60dTQNt
WDk+H1Ga5G81fAA1h4THFgFhe792OJHRV9kfo6Y0x9Ys8wDQESwjDSTzllltAs2n
/nmbK6dlOqyScn3ibUJE4mKfirJEQtFzTb9YKq2G821E0FiiWk7BqgfLgPVtVjGy
V1bPpWqb6fe/to++OXvjFhkEXrNWBhTIYZ7hMsYz68/VCVPefDvb3ng+LiNIxzeg
ycgRX0K+9PzUWb+DZJ+CjIelyp9zVEH0HBtwuw5+tabDBqlyBm2LlvlluHDhTsCK
z06uEtLuxT/qhDPPDAeeNANpno89mA2IMRs49TTgoZbIHHRWdABuGSYO3Q0PqGxi
+6cRH+muQqzj2t0L6CVVDT+Jir3AKAAIw1FQ9Ka96IQVCNYw8Xoxk2MAY3wyW+yF
TshuV/Xs/QuortQJeoBY2gx36qCIBWsLzgTUfwoGC03HavuAPMu85jj3eKcWlVvn
zzsUShxmQp5n/Kad4/FQ9eN0PaCRXAghuhURU6ePC2WMRQDQEJzAa5kM6akHzFfz
pqaU2CjILBnu//fm2caBKwVGSkeiLNPGG8ZexYsful0PBfjzwZxVbUv0nXSoOwty
TaFnJ7aa4lBiy0IEohJMweeMDBhEfNDJT8YowhSylJKATSOsbFySZDWO8/pTSlEk
77dC09mWPBtfGj3UYcbdUwAX6/f9VaZE3k8iWlaEzEQDpFKTX8oR/fC5l/lObS9C
HgZiD8x5xG3bBiKfM/mnZD++tjY8VrTRaTeYgNh+RibjBn8qLBMiCNVfq/8MVImz
u3YDaObR3xcvD3YMGLqoa+AmB0c+8lXyRIYgsjCaTkWrPko0qoVk4o5jTS7atCci
8EBa1mPvUMb19UcfSHJKK4EU6Lj+ZK7+JM6Y6pRMfoGeMBtji82U2gKxqxRh+YXA
/9vS75ARgvggdVakibO7/urXAvd6/QLXuvV7Xt3ZXdgLZbaboVIFzXE58hGcrf2P
qE6w51Y9ajKJ156TkUb6FcoBiC3LBmeLUov8cfgSo67j7PsNud4YROCMWO/8BMFf
bf4zafpjq5MduyWKjVM1COaOd+D+8+Ludhsi3Z8JvD7RWR4K6S+XmpJ1IImnudjF
oA2J+S8Ug68el1sWIecDDMddCP7AAfb7M5+mLlgj7jMe6ep5YXOzh8zs1+7nnr0m
cFW+j0MzhiZSD997OPNzJqvBWRtKE5JWHqx1q+rFL7iX4K2g4MEdX2TTiTYVYNT4
QRWAWvKQihOClyRMyydt11KORfaDF6mlY1QxNbvP4cSMBliJyogcyKpYOnXJg1xV
ANByN95u7m+RSIAhlDvV7C7Ubl3bPUlMTs0HndlwbhLt66spq6X7bwDpmRXAjVci
BjMQqCcM5yNFYNt3vAea8k8Kb526txihpQZCvTm+lYm8bCmSMeuFqRMYMASx1dl9
pjKNVpFf7IHKoZ02Z201O3skq38n27aMDQybRWsq4paFe/nUTuZ7H7HMDonOmdOg
pHBF3FpJ+thiEFkSX01OIidXWm/t/+wXSDND+xIEdvzSgfpw5g7jXRJx/n1p5TG0
WHmPVBCApdsrvvNpJf5n42KGMegsWb4wilT1z7ydNB1VB9JsJCMxdc63r4ZRWEp5
D1AYnjs5421jo/r50fccvS6MOei0hYI8MNdz+/VfbufWawedei6IzKmQLqr90Lwc
/e2Dh9iMViMCP4toRRpHH/sw3wWhN05kWuqobwS9UM4SHqE8IkjhecM8cOMUf+rL
`pragma protect end_protected
