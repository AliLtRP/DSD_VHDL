// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bIpRRSkx+iRgcCskA3vrWJ9v3OGKiyruERntqELX+LEmBoK5IiMthc5nfXDmgbDajY0Wo8LUE6nh
7sdY9uhO+ubnkMw0ZKA6ZjqK2sdBdaAi5r9sNSvKL3gU1fYkQBWKc6+oZAx7Bjorv2AQSX2fUXnC
PcEk+4/ZNcDLMT2IfL1hlO0Ax/L+sOSXkKsc48RkijvG7iyuV4jbN9E9IicHL5fPyfUsGFxP8BL9
0sZghl3b2RJv2SxkrI19PpyXUc71U+rR+vjL1g5ROJTIW3Qcx45uR5t+WhdFtsngU2A7JsFJfsb9
WU0adDKvcaC5ZctYE4RaDcjo3IT/RQIOcTrbzg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
r0XNPPTyVMbIObH83u91rXi1ktPwHsYlUOAZgFkEqdvvZv2bexe9JDRdHneIlMxmtUyn+p/H1SXC
1Pwiqe14Wf/pE1RNyDaiOP4cwF5JHASPmMpGjV5MoHeTQNQ/WTroDk5TEe8cl5CpVg146mRiBrc/
PyI03icrhc5UxutLSk7imCXdHxoBVzNUMX4qqej+6WaUWILd7JfUFPkrGyLIFR3TeAREglfMOTWO
pxerBuy/LnNNSFVeZtpcsuPpo8M2QEdy5/4inNqK1n1NRzGmTi3pk3M1Tl1KVHlE2rJJNjFlCOD1
Kxca7uRh8/WUSLzW758ho88uUolCctzsPSQ41exAig8mk6xRcLBxYLXj+0OohGzOtP577hncfDDc
JZonJAOnCQnCKbJlw/w73y6EE0942E2eJrLeKxssUxi2qK2yI3Aq9E4hHwXfnFBqLSyJRrK4sKRi
RyUHAqMwXBQUr15NOtTTZfLT7tmHg3SKD4JqBDG4dfVkfis8eACtejDxwqPFcEyIaAWAmLBOlhlc
q4453Zw7hw/6fzHnPgqhuJdh4lHsx1kOTtUiNobzjS9+xQFupVAxQVNfYcLOicKhEPAWX2CY+u1j
nC2qizl/jDaXqqCwa0hlK81ICeLqkBRuLPzoC5yAVCLf91fB+TDZYqVLKyL/NN0+KCrCEQfbK8E4
9BJ0DjiMfbiTP4fMqLsRpjoN3eBDfqB5ll3IAj40YnDgRnQFiMnZU76eWbFj+4g4bfHZtsborQN/
IIDRID7AiK8g5xBvVxE4HOaHK/rqDixwD8j97O0IDHzbu/jD3GpesKUQOfz+pMrT1pW4NcGpkj54
+hJLN4+SJFNynxRDBfLTfDbZuGMpquev6MD/DFwmecHEc42xGC+f+VEAUM6d+ZCGCpkBmQY2BnZz
VlUZh80Vt+IDRk6cMuSfDluLPoxqzirAvoTYJ91hCMoF83MBNZGHkJs+oNyKB9xwne8OjIq1nTJp
upq58N7P8kSU1FlQq8oS0YiqlNG4LLRJ8F55VLPDDFGyi92M8a9R1Uh0+4I6MUFMt3+KrtRu+ZaN
L2kL2BKzX9LH9/M4KBTkjlsd94Y5nbSigMXKkO1ERgv9csWcjcuGGZCXrgU2KlxSw0D3kuss+Bqe
61CRGqcwYQyzVAxzZrj0x/aR9e91obWpd8+LQ+NK3BsAm3gGHCMFpUDsckF9X4bj0VHG1HGjUsmo
5t3eGTgkzJTnip4R80nCq/ukTOhMsfQG9BXrxR954hXZzcsDfiZhRcpQ2YC8psDCQ8NcSgTLiclG
up8smFDiR9nSSczv2B1ksDRnnyKBAOmRGK7/QWNGSybmodZUdjOavAviGIg0/vcINe0cbVVOYAzA
jfLhOX7YP5XA3NPRKepc1joPKw7Yi2zDBr/eDQR/ok12OFORf5MEQTmeE+wXjFvcpLP9aZ8bC1Du
s/CRPu8Q1gX/oEbcTstCkuAGGhZ2RJ3hiWekYz07zfXXm+J3vabMBmzJQXMrUKxyDZ7OSuOrm141
ydoTYrOCpZnQJrn3O4ucrvoFsOCntoFHpMSYWua6+qAWVtccX6wrbFCh9E2OtTl9zTficF0AcdIB
mKfJtdnhnLgQKm2TjN/NEAdzuqt+/6Pj5vbIltMNHiDwPotzmXmk5aejQsG5lBcBw4VdDQxmGhUE
j/0pxUfbELn4oPZl+ls1esmUPRmNwUPLT0Th67ov7GzaN5CAcdKa9vLWfPi282GuLAPE29kVajkW
EspvVhDtaXpp1S3Qvzr1sg6BOl7EsJeyT+sb2Yx/y6+xNihFXzLY9d+enq0T80J2DHw3XoANaQHj
p9pu4JtrklGZ5lrVXKvk4K/fJQK166Z2E/HZWPbcSoWFxOBqi1hQGw5py+78Azmz0lNe0u+qRgH/
nYWGg2rN7D8QG7ASqFrnFj/R0on8JjIMVOG+Reb3OnWzE5eepkuVgb1pffZnzEVCKMzpxAqkPzIz
zgyvaDnF/GrN/TViizu3sSM6ClWxSrdfnOmGL2Ey7T1ReDlgYWP9Tcz4dke82f19z+KooUaQX6tZ
+9phB0sqonwx8ooniJCXxlwJNaD8LTv9UAZRAcuCAh3u1csqg7+UWIMIcOhxo02mYDyPtgTgqiC0
xLkLhmZhxWIxf1BHnbsVHewMl1l7MNJrq4krvUmqN0ZNreAsvi9WqDoQe9L92UeavY3hnpPT4tIa
WCcuDFKbU5hI2PzrwIo4Qchd4wmWjqDjZtmd6YrbX0w/3yckv5O7ZXue7IGJn2bqRETXnX2dHlRS
fmiGBQ7p5ng5fdtIB0rcqo77+tzPZDWjTX/QusxDnOyfMvUfjW8AXUmBYlIMsOeYTyWSjQKb4YP6
q69bi4TDnLbyyswFlGysvh40E6kpo9VPhDrvN5bDQ4TVTpWTQHt5HQV3r1JBQAY6NEsZ2SVv/g5A
odo08Xt7dz2WS+U0R7dLJ9RJFwN9rV567FN60emC7D6I8RP3YekaTIIZcsT+MCadZASHlU4jT8Ig
b+2Wzc17PgVFVaUff1mYsAJb0oQrDDhELM3HoCv0uiwekbFr43/lEgRBr60cUmResfIT3fvv5zGk
f4TSLrxJ50lEic2wf+KifzvSHf0EpPMCgA6NyJujhpfEKFP12UaUCEJsBRzmjxu3Cm+cXB5nhqtY
ekfT/oj00gEJgCwuSY3dXGFZ1fIOKpcKSuFJcxyZzDSJiQJNGtBerWWtkzIPrWPeQYwwbYfQdYX0
gwuvEuhZvBhPeHECis5qqwB5M+auSIFr8gftqSlPG1HzAYNlJtnTEitm4YyWbVlKVU2/d539wDU8
DPKFfEj+e70mDuQZIEBgRkGLxmto/wRa4u1YFuDRK8HRmG+5TUri6iOqBkvp4RkKxvU4Nqj7H/6C
s/Nr5acuTFOdvaptyeUv7tyMyrDkx7ip4Upe5d1wNyRtvJwT5cjX69DTn2IRh+yDVocI6+lPlQRQ
D3p8r2j87i82Ef9fANu0qwimXRyJIZ7GLXyrkJct8jdIiBO7f7RYlut4ZcAnpX8HZo6KAfvMY+qG
r5eQ+7lEMHqWN9ENBXI6YnTjlmId23EtbOsK6atuP30dvjWRdCnzz9rFdz15hmB5GkeIC+r+Und0
AfV4ilX2DPacZyzCpFCO3QoG7uvp327UnKINfxvrT0SZrSZZCJlL1LNBvzJWxF2ySlQNpzuPC+MQ
IcY3BVHJPCJoH66vlf1YaPRC4aOwKLIr6l+jVJw/l7KNbyYQPmwgZGpeWB43GIBrYZqBzRfJWTYl
TVYoNKhlT1jiP+szSYs56Vmt/JFce20HHwrnd3LrLMa4c0yJpG8jw0Nno6o22BPuqcXsCbBeAi+H
Qg3Cmf4GQ5R4LSQev9Zj8S5zSs0nD8nVZAUAo9+alISqdBvYrIdY8Tqs6C/yD1/WC3Y0wr/Ya4dp
iZjebZPv/r2PBMJaBuX69Sj2WgtkjgzbcxLANpoXix1rvR7V3zvu765vkDO7GHsS7p+WVuOOfRVf
YLKytSm/t9vD42qxl1KqIMEuHey2ph9RxQ9RZLz9H69lPKoni8yVxk2sHNHd4FygSh11fOoCH7GV
Yux2deUUVTEe0e07Z04t+G/wpvnxcaGpoKszHFC/DqXGkh0rDy6hsC0P0fTZL18mxzjozRDbxWIx
68D2jT5UFHzsH+Nku57iyoiDSy2C4DTMlb+9gP7v/9r4MExHT5cxVT9YS7oZD/SJ6dFnlbbjLdRq
+hW2C41hK0jOevaAYc5dd+N/u3LMht1hEXqDyzb/krwYve4+5o2rTmSi4NT1MVAVZM5eDryowGyS
eGhf/e1V2/IzDtkVC/D+5rBNWrsRgM78RfLGop+XVAqUvDVSr7+oZ1f5Kn4ECWnn0Rbglho6EcYi
MOKBfqZFueY3DaNc/pIY+0yzVkP0IciuqNqPH2/qX20m8UkDwaby+PCx4ZZqubEDunPxFJDgiKwD
1gaJRab3KLUq6DA0KTy1MxraZJj4UVwpsaZ9r2gLMq2TMrK5unPsHeynOjIH8zqS0QSaoNBT4WDH
/FRaiDYkIRsAp+04IX3EFI6TM5GOTtbmlt3+/AcDpzwuqO1ZraM0i2Rm0qZDLSOsnrYTrwwZ0jMw
bOYlRg+riteDuw0oObu5+d8f/5i+Vb+oyK0rmBRuA0gcLQn4To63D0rED6dTLomg3EQymHgLzbJC
0pUxkLffO6XVAdol9BLFYTeq1lSUXNq7sSo+u1RO+yllKzgbI8Vw2/KAQKCH9eoKKalR3TWOkK1y
pUXES2c5M02bi0x7vzR70H/QYlv7ug0+ok9Gt/1e8rG5E5dwa0/XKpp3uQfNmsw7DZCNh/BFeySG
FKm6NN92KnjJ32rOfKCYb17gl8UNx8iUFFpxeDMqdn4dW6ZaT6tAwpKUAbuHrI67H0sjxWp1YL1T
hjyQn6ubxzkwWtMJ10RNggO8LoLZKZj1hCNj9cHoSjXTmijNk17jTWNCv6+x5VtvDHX9xAaRofF7
dS99nLUbO6f89MpaJFYCSSXqWcnT4kNwrN6A4FjvQXb4COa1YsEvzOSblmqiIUT+IEVmlNMt0eDK
6ZxI+kzD3mof83qwVCHAXgFtE4tZ7BUKXbG/g1GpolE/4o/tTMKdT5ef3y0eOXqPA6OEgZsNKQYv
2Ir7BpsspKn82XZqulMY2EUH+3NX087LX+BYTBasGJhz1i/YN+bHkrvFcH1Rt66pqOGgcQuzKfFk
pWSguA/CxvsRlxvsV+kjELx8MsXpzWZYC2Tk84KXCCl+NCgkW9omc2wTcznHXYwzDMLL2VZ1PHfO
EtXrgMq3vMxtm8/VWCO4QCQQpBdVp8jlhWz0f/i2Zb63F/qFeF04P5Kpb3sv0zbbSn0GnR5dWknh
0vRWilPuFHh+QIXyaGKWC8Z4Kx4jM+5ddgPqF66oSY4K9iuwH/rz0MdxxNkrWnIyy7bh1HP6GCwB
f6mp2CGdm7yH6TUWbdrXh1tBeNk8krPQMRy/XiTZQSSh9hdLx9wdnEjR0z7dYnATFcaRbURRfWpJ
dc7HTGl3LQas6XROwuJ7hUcCnX5nwa8AMYO3fnSGzxdgXQlVVI7L/QrJSfjRixt1uZMCPgYYodDO
iEHA7dFtpTKhtuWrnaGnMHqN8R3REaI6RQIUKh9+pWxdSUj92xHJr56ngZ57SeOOcxTIx87dOonA
tvd4ooBMEaxj5vZhkxOCOyN0lZe0fGUIBQFQSOxeEeI/AiQSrIcyIgw62O4dLe9V5lZzx0+lICZv
jHF5dVxV90gIt0TITI8pp3VlvYnQALyZSOLrEZdP9Sh++q9ds784GlSTB5GQH5cQfIEQDFcHPz1W
aZR6G0+av2RVMjnMsVLFNCq8jm/UtT6Uci8jdOzjmBy8Q7gJ3+TJ5X34ncLW0fKpKfyYOOAZzi1w
/Kr9nocDiNOzqxHK6L2RujzBMhDZtv1KwWZSODpgLmSqRwTqtU9mmDSCOYSm/gOQ2T4u/mLWgmav
COFuAKeuKFQbEQp7VLpPm4QGkJtNXwPUUne2gyr83w65rA09xSOaftsfqs34nBEIZBpf2CS7Dw86
Jj6L2wNGChN5NS9+U9RddylpVrdtOHV2Q/3Y3yxmnQhX0MR7BNVRU3IIiiaWv/M5yadzyEDAMQNo
Emcb8XOO2OeWrSnMFVPJFOCAPhkItGMkR8WXFQXhmN3sfAtdhYE2puGnpX19sz3ym8Ou6xrRGWSC
KDhrx/8Ad0iFKg/M9WPbKA9HagHjwejR8CG+Y7z2t8vDETUJiSHxrLcX+ZpUljTKT80B2HClxApU
kkbC6OiGXC7Y2QcUOaClscbZMSKEy37kRUQc0YQkic5S7EUT699PrmuWW9Iab6XZPtg9r8ck2cX2
PHgE4cfSlAcXWrM5fp/gjgyTbz0MXWrLr6PZBUcpA1ofpHwecVrhKvnd0dEbc0ywBZKEe8ECkYPB
NZPb2Q6BnjGTCmECPrFIjE2cdUQq8bEliNEzDSA2mdnra2rP7WL4PNemn/mkenJNk94mp+46Q70v
OQ/ZVHkSHY8WoBLJD7vJNNQjdbvEdhqzZ++DZxxXSCneXcK42JgipdAboOTwvOhUYb2DgH8985n2
mRBV1oqsldfx8klecJDwf5gQl0KagH8Z/P7LNhb+PpSO1N3zXQ4c+NQ4vvas7J4kkUAcx7cWqQYh
39jTRhmMPOS8LF2W/626Ozt/Cu3xc1c+8RRuR9986IYh7raYjYNuYupfsXqN/DtgYWYaiaj6JRvZ
uiXaiC1rpjGohbXO3lLloCZLxLrRLXInOyYlrDHuvBu+44dPxfxizG4DmK6IkivcXl2eNfy0FKq3
yVfOpYnSXPweDG+v2h/PL0RnnuPF+8JrffHXKzVsv06+mVm2woYYZJrCRQDXrqQVUD8R5jvtXu19
ezpzDXXGaDLI7IA4J1rKiFoW2O+VPbss7DGIz0U5fSNPQuHHIu2lfZLWlKdoVeIV7M6v6qbGWEqq
l6JHOwgKAFtcWaS5ELXyMA3/+epywF5W3d+DsAgrk0402gmNyRoEKFdVgLUCN+zV8+mdIjFZmQZy
iT053YKY7Apk1yZv2kvqSXjIUEQqd8E5CyjaZyAf5cYVj+g+ty92OIElL6dglUbRVDsnW1BPufo8
+8NuqPCofVvdsVo6xI1pw+R38BfDlxb1aZ7+W8HqUxurRHK8hTlTUAAY7pswdgRdK4b3vDkgC5n7
IoCUADYk/xhQZbj19C1ZtUinpaIVj6ugRVBtEXuzZcTlPDOZb9cc0ZxlI8VG76S9D+ZN1en7xbKp
Ztk0y59PKWABvijc7XbSSrdbAHTgINJg5Eqyj1eENJsAyMybmsGLiCjdVSu5X3BhsfLmPmznj8Uy
S2z8ukayutETEqwjNd3FqldE3G8Ro8SAzqUGlnrKJ7WJ7LxoEcXa825eoPB9+vtWBtnRZiZSC9is
wOB9kXfbnlRvnGtgMv6Uz0DH/KyAsYiKFQd7zwnaL+3qC1yI9m5qKUSpUtWkvAjriJ3mLrXlyA3Z
E2mQUbF7GXqOjKs6oE/O0LAUOvCYvOdQWent2qfS8EhVZa3HoRh/nNbn/mNf3dq1twFeorGaknp8
VdmYqWn4YyWWtwcbID7Hu1cFHqqvAGIWfsPFzIwEhWYUDtRyfRdZu2nBoyDv5HrkEk7paQ62SbDo
JQfQVDoyv1dElvPbaKV1JHEZknJtW9CxjMqncoWJ3iMigP/L2lOwebYqjK3Jm9gEgmre/UwqaTFv
2UxnQUhTIHbSrXqU2MHNWfFGQm2oAaL5ULG1ECzLTa/9fILVKtPgj2s4qSWy3HwQAD7A9XcTFkx7
UL7g1eKnjlq3iK6XmltoajRdoek74DvJ6GEuIsEanXCF/0sw49DDHHKy5+u2b3YTnUDvooJQO3lT
2xCRL3Vi0sCoITsQc2Gu5ZCb663tRsq4oItPQIVcPVo3+vMAmg/ubr+MzpEiS79HFlq6kbZWzCjQ
BZNRadUWgVG4HaJgIEH6M9xwMNwVTPoM7ksGJcAzbp3OdueILNse+1lkQQ5XJvVafOmifbBSXsHc
CsMSYinuOVQfIlUuaaBICez3u66GT1uUSSmu/MgG37GMpVLFJ9k0b0ycxvLuVcCHIe4LJHReKxti
jnNkBnTLsNjakBb2boPg+lbdrXN9R8TnhWzGanxEjXXzQV3RPOp+djVV4XS1EAh8KZgIrlIFPA1E
ifcvBEILub9nK5NJ5MB+dklI+XQHZ8dGpX2a8qszijMoIZiAGN5/0Jm6W7F5fuRoMAeB2z6VI2uL
48Z4KF3N+FHdxAERrRi5ymdLkFGyWpzrKZzDY5bcJ8xTeE/Vw09vUNIwMvrSdY48kT0LCTLWgias
Kt39YpEQMHOvk4+U0ljq27/51aZOZxAhCmWt1Y+Tio0+AhyNQolIEt4wopsdiwmPFQOW4ZUhROGa
yD7E/B5N/bx/LCiF1lujKK+RRQb2pwIOKJgpSLtbD0CnNgjoh0ZRfrN86maWgGSYogN7/Lb/Hbm4
1X3YuqnVExAOlKUbbSHxzmfffU8CEf2YYtMSl6MV0LX33gKh5XDo3Xwx+LUEkysp0kv3A9iAaWuF
GsrmMWKeBDlvG85wb5qwPf19b1b6O/N+SJr4OTGfK5LYxAv+VPZfHI4bSdwjrUmR4dTIcGMaUY+M
9A8wTyG4QvuEx/f16OdYuNLRfLUxkLG9eaaXIm0MZe4rtJfi4A2BtlUaBgvhET4D79VpmaJUojto
LksCNEqkLimOd0G4GE+4K1s4lX3uK1APxEkfJkJuuCmhKjCyXRULt1TWv+MUyQLpphmrwghU4B/T
vVfjNBP/9JHunId7nfv5yQ9tCAbPssV15/R96qRLAt5c+dR6Gsr/uOfyhroQe94tlMp4FRTbHzfe
htiu9geSc8kwA9zMVLJXP7JO7FFzRq8KsadDN6lSrFYCI2S4kcq/A4XUUjJVKvUfU8B9SNkGG8Rc
AQptfPSF7mmI0qBiYFpC5yshmvx+bBdCctPAs5Do3XanaihtyBbB5G4ihm8FzztLaUnmcrQMDx9m
bPS5eg01KtMiXzf80nUg4g0yi8syhXb7DNABztG7hzAmRVL2xadBZtpT432pRH+UyTWGMoIgqUfr
Ap9O0qG860QZfuun6YXMce6TYNHf0Ln09bD71Ru445em7TtiYh2pABXlM1oPYOuXTA/1t2kYDHim
VgTU2AIkur0tqPBnuhxtag5vJrbHdlvHFqZYl0iT1JblLtd8H32eGoTZLLCy1tBcrQ+QRw6gd3Z0
0R0w0xJgO4Gk8xPrcjSuy1wToY5cyoOsC1PaP55QrxzeTQiM4zxp+6dqXXNhY/3nuSpiORsqFN3D
c1/WuXbQ5s3sipB0Z9ziLsfR3I5TaAYlWNthFhfCGR1lwoxGqvSrRLMUXzauh8t5wEVpdp/ww6Qa
QBNUOPFbaSSJCzh/E7u1mcoOirPvXfY0qPiiumKE48rfsGIMQQ+q7+gjWfbcijCUb5qhIFQRdMOT
9AjhJNnDb3+QeoKLR//oN4y+WsKuZDJAa1Rb1j+fukfXMFfn6a6V0s+jxKn2EYj7Aq7FRdQDdCwq
GcMv2p7nJhNN1t00NibOO/lu1fZKcsJn32BZ84R/TI8AjkqQbtZsHz6tfT6/vJSE9P1eX7IzcQ1H
qrfTxp+lqfquRVeUUJZhUQ7w4OmvU9nCiuhiW7VnTxH5vVIn20q9ekIzuOFueJb/fV46Ga1SA/1M
08Fz968ekM7ADC4ZPy5tooxH+r0ChGTVnQDDermin1LUjqH/DkkNH8hcy27PEPfx1se3FP4V3kAs
ovQm2vzAmKdgrfrl4qz8GPQhefRIoWDxoGBVTc7004o2u4gu1VRyznA3AheVNfZUMI66X93l8Spf
xRjurFmvUXjvDoqnxATzVZ6WqIKNu8oqczZZTJ+22XjrJJUuuzoU7ZNkCHz6OiQFtf+a8QgoSJU0
UNrqD/1733pMSmPWVYsZ/HBquKY+Y/2b8+AzZ8nNYPYk3BficsSZ/5+9ZlMujQty1cxObUV/YYcm
Bz+okMg5oa+Yl4nslMeIlZoKhdWpjJILq/dyEyZHDfydstWi2tJH25NxwgIODszfhicEJSiabGRD
5tkQo/dV0X4VKVqMuywF04ibQtzuHRQnzNPWZ1j/OrcHP1Cmm5f5GxuUmTPTDhcCeQYX1vnXwInT
XgwPTdHN1Xj8dNY9l0jfOZbyIX7MIG8n8MKSUE1u1dXxThPMMzYIUgz2tK/BIMS5ByAfqzhvD3rD
mg8Vz6V57jM0R7iGI+PKDyA6Qq6lS5nsDurQXPFxlnbagtUZgnFIxXb9yDMj5tmOmSOfL8vvAtSp
7otflKdltD4x+8YOVhwe3AS7Db56fc3tI0xL42lAYdGUVt2T9CpoGqPTLXp/gIvFFQA0wwYhLxt7
4hQ1tcEnkLavHyCEMb9bTRhJS2pHjLd1+gc1sQPYrXa8Fsur+rN00XHe2PFEVplwLTpqMPVoVIN3
A2B6z+SP/RriKYI2ZzkS2X5bTJMJFcq/rdWsck/12/rbw0spaVPLMpBRfAbdA8oSV/pl1PDAC/zC
JuVPhH7KlA8ej8g92ZwAdrBffI/UDpBi66U6XfN+/Z5LtUWjeAB1eQ3s/x94VJeVflk9Dcrm0MUl
VjMAnvX2YDr6AYpeR+q1OP3gGUj1WVwqAJOmqU+dQx6kgzLVtTehzQ8gjHZruB3t21NmpvmH7Irg
nIJbRbflXDV4nJl+rJgTmfuufLFk8kWNLxpN9tLCeGPz023K5mF2U0s2+CeSLpIcv/Ri5lUJ6UTz
46mi3OPCRgsiGxv2Fe4la3oxrVJyrYYoyRkUuCpQj4txmdukkwDj8Rl5IErjpykSQRYa3iu1Z4Jj
PD6p2Ecm6Vuo1eQi8KiAkT4xUes55DP2vC8KtpeN0BwyuejYYcZEcQMYXWFDESO077tziIm/8GHt
anwfXEIPZrojsda7Wm8ErvuC01jVMzbHemGxWOwedXkmQ+AElpqgO90SpkVEqHFR3iPShwArRAQ3
+lNZWa2tD5whn7UC0Tso1xr51NBu/Yz5FHjqHoOAj/F1JsKR3ZCOo3EwxD8LNP6cnsAENYoVao7X
ozJ3zkpWyu97vnNpc026PMsKY6kUmOGLjlhbfkDgjm+3ZxhYJzygZ8V7r/MXiTgcLj5Y6AnA/nDx
Dtl1qubigvN05x19t5zRIFtNJ0j+rHCggreFu7G2fZ3o/UuPOgQhK67bZJILma2i5hUvc7UdqNZj
L6FHLAAG7IcditV6QmQ0E0m/qqw2JOuKqVtSXm+dGWpTwg+bkDEyaMHiBRB8yR3rahjIm74QyuC7
5MLb4YPgTpMpphGTvFDJ7vx4F+jAb4NqBefmTATR+N1cB50B1kGfcWrET6aCCXbb+Cs3a2rNzzeE
hkYB6VslGGR1HQrBkD9HecToPXU7OmrmCAIIfRyq2JE9e4C/SEOlxHU8j4kJH44rPbVXZZPbkGp7
e3Ni1PJyRfw6bpnjeUP2XeAlUPWbHXB2/2UL+4vE8fCn2FIXTOgo9A10AmxbuCWqJceBwXgFg/2S
dlB7CDAD0e5vkhd7cCJsfgJDun/FP7cuiWAxzyuh1vAvjzssc4XNVsHbSmfyRCwP/ZBLnPSC+dDY
zP/89YtBUD+gNpEEVzq6thPjKBXPGLGOjHRLk8PyMGn6iGXsBjXBktkaJcG4BiHr2a01nycmIbpu
1q2AGK1WoexP1ZkDw6Z6PMPofo/5SEFBdZoFpuPcjZIiPEyLpaeciCXE9jo/kSsWjoHGeqXHpNVu
JHoZKwO4Mb7vfmvEMHWqlJnwT48KCU6fAlXcnMcgx9D/zi/vFZJ5RXHkSAKYgPZuPmS35M+IT6JC
4dqvFXA3excnhn+/gmro3aqi4u9Fb3EcQQ/+OVZUQvbY0Yov+uHk4GFaYzJiZ6PD/GZvkCprq0Gs
WYyhg8fYMNkq/vy7L/VF6Nih/64SL6MWoyyZAOoMHJkLosl5/Ow6UZ/deObV0Ofxib0qd3+hMZWx
Lk9Ymc3mAqHoabJmhPOE+Q16Nnvuwhpf8u2k8XZSqVV022kgXinlmbeweh0OqzFW+Sigr1Gj37aS
t7FV+v+1XQGzXfP4yNB3LgCqnYfed1locqGoQWGxxzTg6kxj/LlQOA==
`pragma protect end_protected
