// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l7/ONiua4YXH7S6VfUBhDiN5vDJVFRD3Zg0i9NkkjRweYF8lBRCsieJ1TBfeB1Gy
TNSV8wXU5KQMaLzzPhKkkKuJ2NNaakLh84QRM5xGGxUKDzwe1SAcKkcHxCCGdWLp
uRj2RPfqNMjg8P811M3MqsK8IJNzsRiX4mfh62AR7GM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12560)
fpkFeJqTXiXH4NJwDIlv4k1CeZHumccyZ+KdnJt0GrIi4M20WoU0edqRg/gFeEBC
C/XGO0AlHhnIPSy/ZaYvgKMsLO6bjWMQgvzARSe1gYvlSFH9fPUSuAr3bQ1rO+u6
pt+TFbEX5XLQ5B02ObkjXA3b9lgaRNvv3n2xOgaWKZI5oIpIAJuLp4RrUsjS+36l
F1VGw0q4TIR7elTIm35bJh/M38K158f0z4eA+hnPe34fDDTYyJRQoqyesNUL9rB1
UOtvo3/Q0DQgMMUw7Qc2oSfrab3H4LvGPMHMosU63Lxsr06QJZgvrdia8mO9uthy
rZfQyYfakl7kkKN99JPiq+4+kKbr2zkXJRLjjCq3hOdCZyO/eOmcUP1cVJ2KpSwp
rhULVZstwEYWJ/fA5zXB59Q7dXGlb7Rt3Yqg+pUyXiTkqzaJf5dyC8H6CI2BKEoz
WFO54GTuStAkdmLEjiJLYC6ypvKxzCU5FuSFCIBPKQAhEuIr/FZe3jWr0oYlGCnl
xGQ27GPwhX/8B+zTVndCbDX46XxENv25l+QPkxxJ1km/3TyxLFx4DXDA/nTnALEM
L06yYj3ekr3swKINYmDgOs0FasoDedyEaVDLjjMkuDR3lqen0WVVZpBHiClCbpqD
hiZu+WmHvdxt3HPF2/rv7AblsEfy7/5ffRaDTn3/5XCao3o3Ua7CwPmleyxTIypC
6cSDFsA6HX0x3Bj5f4IJoSsI7kph5TLrdcIzLbuIJjt6JcwAlkpEZ6YsFVFnkkY7
KG1USYnVNtVJT/p06QYO2GgHb4KtBeezfTSNbOIALHTSM+WSWVW7eRP1fMQMIlRT
HXEpFLT6sGCxMqGNUmYtthekEIcALt01AEC7CA0g5BX5JgaXgF1BBGKYY/evNWsD
hkmQv3dbRwdylmNI+g+hRRVVdXEwvSIdwpjoK/MV208HU3mkczG/j90MfsqD7CBT
szi/EvI8iJq8KuxKONs6NqeESiwlTX006ZTvL7xCMk0trwLa/K1LM+3FjdQBCA4D
O2DZpXWdd+4C/exO+qvNz/N6QNTciq2JNEtM3XOwzmTebyRSKIgiu2uInYBZNdFp
dN2AreQE0TYyW2dYwHvUWsuDAkn0ZGFOPvpCl6pszLqdaO2Lu2pJGodozU89u8pg
GbFxyYZ7m/NfOD4Y28vmOai2FHws6BeqJmWxSSulLSdcGHmsLH7VD0rxuyoSVE6+
84jxCIgBHSSQK7AMLAF962Z+3AlWhl9oA5duqvZzt1gHeBYdQXwkbhuZ5SA+1YLe
ADYS4J5sm2N0fR2JXngr7APn/jChcD0+xw0zLFZevr+7IkxHEweYf9IBVpZZRZ1T
qRA1FNb85C+Tsyk77UygQX3M6lQxyL19yVgysbx9q51CqdTtxpy6+8JBvabcpt2N
eixxP/VjPOizOEbcyeLlcgM9+8E597Wy4/4flxNgSvNFWdNL2EBl6Aaj9ubf4rQa
vpXyx5+LrG5/XQmIKok8F4nooq5CxSklbPa+d9DhgaSaYkKhe8moN+SZ9FNypb7w
v9ZUNzq0vqLSw/WTUk8LvPGBe3K7dgfsAVMWa9zncGc2vQ8uo6A0jUV6ybbyFFJj
tXqP14ESWZ9tgEf3a0v2TUSpYc6RAwEGnTz0ueaunufxKNjEGYQDW6T91cxPe4k1
91/+9HK/+LotNSMg/DbLn1L2LrrhHybbAOaMnLWHgFY9AnXPwalLTEjsDhXLt6z6
r6/4F9mjpgdM9UY6215Yi5eHCUvHq44e5OjqGFlMoE/VmRrxCReZr8nLPe/2O/uA
mJi4Nu7H451kg5QX7xaaYlh/jO3FPzJkDYhG8VcJw6TKE6LIwXYWpK1QK4TMrMoF
WP1S6tOGCywBeK/SmPt5GyB8ZEUap/gMSmQDMTzavZFqpQz7BkDe2Q/rw3VrHbyX
8q2RGj6TVvfejNILkw4h5oG3zKPOW3ruV6XakqrsDAmhpG/5H0qCm/wd89UKPOIm
2oEZ2+j7s+oKZ+k7TXpnt4RfT1GFRUFNcMHWqd1ufzlvcBJ/zdDYmSI9BAL9rXc2
KPsjskyBaWlINCsue/t6+TBWby6GJ7YwqEjSweVVTzkQOvtakmFcvynrM3TvcM4y
yOHie622B/r3IpaVzQuvy057o/6fJXNAowMjCiExfp10YM+RgPkiiYvGJSgunIA9
VmUml+rKj5qpaob6rUBq0npxLhd9fNx3oXAzYBz4tsBKs6MsC+jLh82l+EjDWRrn
0FlOviWIqSX9DyNVfp8VoS6SF3CPLB8pCPhLY+6ICkUP5+68JGOrge3BZ9dRbIS3
FYQUcEds8Gdl53/JKBEhq8CyvLsx6UJIbxUta0Eo2ZZLdOzRKJLPTbReEmitYiuB
XykU7iWgKTtoIXc/Vc+urlRU/0PvwsK9D7s/b0PcwdFwA4pPbvqwOyAmPsbaxQaI
5j1mOeHcO14da2C2yBhWv0YiexhqNMG0ZSivHMCNMO7Nrm6sqPD0fgeX0wKN4nTK
dEWs53pRiN2JcVVsx7rqFvBZw2K2FuogW72BRUrz5N2vP1cj5RFbBD/nAZIa63M3
rCiRPjFSm7XJJSyXELFX49TjEtOhup5WTN7BnAQ6Gyx6w8lNhr1oTht4B10zTau0
49PmGGrj3T/Xnla7McdsmMLUcIi4AFuca8UepBbI+Gj/awJCGkx62qJXnQ75b+9j
DAIGWVfjzgK0qYIMfkhACb8HjcJto/vqpIGFp0AHmHE1pu/Q2pXbOXsSJ7efgvry
YDUn4lXSdB2n5AkVBz9T1RL1ok7ckUmC8SQWFioP36l5Z0x6rXv7/BMY8whPbD7w
i6gjaS1zt/jOxrPpPCUHElWh52XBU3dl/AEh9ypfCXIz5gF3qP7RziMGfGznjUHo
CO5bga+etPp7tUq+M+VKW/Du+iiwfQuStTTTGCSJPzT/z1FfEi/cSWsNHAWlP00B
d012aw5VO/bO5RXjLj0lDaYbg0E9io5f3Hm7/JIIbGB53u1pAoE7awrqyfoevtV/
y8GgCXUwXD9RCU3n+K4epZYPpFsi/7FPjuF8nY+pSoSFE0oRCPvbCM158Dao2JmK
aiPZcSM3+dSPEuY9aig0jZrlmB76ARJhAclYT8aMcp9Zalt7/p2eEJJCWnBwKiZU
ZVj4Ko3faWkVOo+/eZYFXvivNDwZ7WShbMW3ZtasSV9QRw/XjjwzdLGLG2gy//ch
NRbGIBwwFjZM6KeKNx2tyrvotnfxbimNgQoh49bGIaoVvWCxWfaacScWWDKtmD/m
0tv4+/9TJlt34M0zq8TdTT5J+vONPOOxp4smZO09aYSvuEtf//Gd9MRO/tZmVa+G
QXwgmPcogQOQJkWnyQFAz+iTbRB4hyHfs902N+17QAKiReXuFsrk+/Ktn/QQMZ0S
p3+ceC7WJhQE3bSFzEknwdbxFbxcYv4tH9fh4+ZdaS375un5b7hiOUNe2GCoJBBP
70tlQyI/uqu3R11jeWhlheo8fKwD4vceZ9+L4hQYmlPb3SCu6sP3pbL+qZ2At+Qv
GxQ8dA/TAZdpDzF4rsfLbGNNNbt2D+PsH3eNFdKSqFp7vFCvjP89iq3odgXRIXcW
pRsAOiCEnxgTbabwkHExjL6urFjiSuO7eh+f/xP+K4OnGVnVUnpqC7MFru9usKhO
O59ZszTRbLnRTTmKtT8REEee1qqNytpt9x/qsxixPviaExjcXwPn5rpfm9/5liAt
mOaOGugewbw0YeC2wxULUvJBqLXUOe57El5FGndcXovBi5fRPaMi9X8qTtggpMx6
tO7I6dqy2xNZwRAd+sf/CP2eu4leTabM9SPyuI5BGTsbH74zh76Cf1hp4mPFRSS2
ShBbe6PCFjL5JtG0g4j8YvyqohTd1w0knmcc97Gpm57wW4DYbj/vgZ6AHCYiJXct
fIyp++hPWFpW6EhUkecSDCvpJ7RHL/gPVQEs7e73SX96Svy6M8ZWZiz54Qp52Wi+
dis10ELMZtH+Y1eh4tr5lQnNydmy14cun7i/LDJr8+pU+LlZXdB30coRRiYMFFU3
Ky/yr/sqUJhxUJqstA9Rgf564TtcyvM9h9UKxR/uQ4xyJni1lv+Q0jv29m+fWw+n
/fW2rJvvuMC7h7Nr+H8lja5PfWVgqld1UFQFzGx61ORp4M4Au1kXARHnJNfRTcu3
uB/IU1SzxOt6+3g8CFWcUkgIERlsKzMVI6z5iqGldb7nB2EoVIGRAWsHFEI107DI
Qzp3IgbEm60l9AYGmrXkGyRtXCe/NHFCc5XIDGr4MownoPZmsEmcNTTHLB7IatLH
pEwjSkeP3EXv4OkZ1Ckq9M3SxU8SmM5BaeL+crStCAYapEF6JD4utAa2T328Qmbm
x3TbOWIZci3skyXBIwTSc3XXXTo6yts+uzwaio9RDYF1zo74BvYmq6YtfRUZlbjY
i6sdgn76wIKtjzhEEhHie1SqrSelPX6A8ZhNbg+CGxYPdyTZYmlffrm/gYYPeLvc
SDrfd1oGbMm/BpPFUgmv7hXpQOfmvaZlimLYK7hvej6RXRJclCASIQDmaSbbB56l
CfpAe3DVNfLdp1Wub0gJVg8wyhCn+dQ4ft8n9+UYm2yz9rdKb6irYaS3Mdc+zy/j
2jqp7sYta9xS9CU/UHyTHRXrBtNrGUIxzAVuLG0Fs5XwGhCxvyBrZltCZic12uPL
QChTeleQJO2wPE4eSIuO6NwnX1kftnxzlJ8FVeF9n2ll9VcLd+MrIOGu58/GqPqy
gjy33bTsI6ccChNh7xdy4RvVopfz4/opCEd4gRS8ON3xLD8gCS58gZyAbK+9fAz3
KJiMIasqleNV4ZhPfa03fgYUN2bdvdgOL35aVbKnQ06P6Ndn3hsmQw4k5vApGB6B
GkL80o4vGkwl8NsJHlSUsuHab8+CDg/wmF/Q2zoFXi9/WATrsT2gRK5+fVyLYX3a
qTGU2KbQ4FVc5inH+jezKtjXYKMoMiUyIDuXSEq8FJC+bCQNxB68jXp/05g64a9k
tFugoSMBCa0JipPTD5x/r1ndFdgluXuTJLtgDIbRSzHEVNoFoUoxaOgTZioKT/I+
QJFasBOQTUjhqHOM6hjQ0UxWOE6bcHE6JADIyJ3ATnbMFLPiWA4cb3uyoGnAKf3V
TMJ9mIPe2iNQ0hE6+Aa4ZS+9u4B5Nc99llvuXyJuHfq1wsrEf+1Ds8SnEUUy2fF8
CqqDPr1I4hMCo1oEtHU3SXSIGZIpvmqUW2X7q0f883sYDadcjjuy++IXKampvU6b
4ZuypuQQnE6jq54v/Y3hnZ1p2ogwiN1AFje1geBaInV/lgeSDHDTteHKAzMUwwYb
bXBZizoSe68h4mrzIpimLT7ZCHgSU9n5jRfkE9SaZEFzEsWMz1n/pKuJ6HAyUANO
hRNpThHBFh14136i8F0rITI/nvEmWoETVAHKwcEPA8RMbLJxbPqgB1PEAlGJcdJg
L2D5nxneP8mpGTFhCs1yL0CtMTvv3kapaXNNpEBisbegtizmWPj2REGwPwrkWmw1
MrY6CgXLm0uksQb0y4ers/+RS2Es6g2DYNJVUnC91XBYZ3t0ofMOoaJoev6zqV3c
FqCpUwkKMhzs5zoid86UMQv6NZTltBYh0iYyu5UJNw8XJsJZ2FrnsdWGPcY3X91f
r8DaaT87+RfKxTi9TEYvjUBkkTQ0YD/3HoVVEcXmTkSonBhIbyYkZ5Qt2BnJTG27
wuBh6zM3pgkkdRkDV+kZuhiku03nfq4ZGi6Zy7MRNZuLqAwS/6ccIp24WcpUhrcx
K3Et0288aSpZFsU/6IQAqRf4nrmnN8pY5KDW/T9cJKfioHwDNZDXamyjs8pULoRl
A9vKDeJ5MpJuPbky5AFtj+be5tV13egRWqrPWKsbKiVx1W/PWgfuAxsO2CsZh6qq
98dz9GHgTEsanWluC9po8j2JhT/Obz93MvxAZvtHI3rJY7vaMKEhu0m2NASDXsuP
+CO66Z2XDhekGfgAlF5s03HDeborZFocHnUqoywBe4NLqFGnXb3rCFIzPsk5pzyK
Bi7v2TEXYb+wDjXzt2z2CFO4RCaOjIy8BszubK6fWs3SQWYrS1EjdrFvg+SSQIYC
GKO1iARf4x6T59Pm+f3qr76ECe8E70+E4aUzwnajSc0GtCASMxp8W9VygcZtsolE
VZc3nLnvj14O+W1sUpTqwH61c/eLGoGF89WwfLRg5r8Z+XYxY6BfGQ36n0Qx1g7l
xF+5zu5EyD4JT5UXFT66JjxJzesx9pIFfua/VY+QgXrzle7onOMnLzXbK47hqBNc
oHqOKbTJ6Je1TO9p13zmUjjVRMB1TGYrihjtPNRoRl1e9vSPyQDRnBvQx5exkotL
neSKet6S41Hk4n7qwiG4JVVGUfx9MnCVgrT6DjAJHQcpgItszzGRWwxhc10z2SDB
1Dx35wkNEyGmhi5qXD1FtVUsVT87gRq3h9CNw9n0X3j5p5MooOPWtF2WrPELD7jc
z6xDp+dKgyme1NaRcrcC0e9NHv5i6eGrKe3tU9vCWf/9ZyANc+CLDgjBP8qbMs5h
NRmMAbubKa604v2ucSAhGVTEckoIsBRQ8/C0/VvyBWUEpNSf8kbsi+4QlAMZTdvu
K72UfH75oSTmB/3NM7VcB2r0hiLopanwh8FzmdE2kkIWkvddH7EHYBql1iBRKjZP
xQ2zPax7yW0bs2iwpbsw1y9FaHy4XkpAAXFd3H9VEL6bbpSyyMkF0FnCy4t1wz3d
ZDVpgTXiBuoViEUkFyKs83gsePzOf6xrUrgTbppXiRa3R8CeNQmjHda3oN2SX4Ve
xd8FiOK2BhmoWTcs7wLSZ99c/xnpKUifMmQuGMdO9+MMfKMUw+FtX4t8F12ZrHq9
rBxmu2jiStBzLqOQNT6TsrwJXZY1KUnDnnPL+wqdHrJTbcdqwYclgqe78SyoXBG1
Ge1gqNzejodeL31yCfUmZkZYsdH3th9u1Ae4k19qrMRUTOLqBnia2cwU0yL6WLqC
Aw426CzsgtWZwqqxFfIco4pJSyGQCHqRCgLPYX0ptQum3W/JLM0/9pIlIRcOzw0b
ytVnL/ktZ5Jwg+zgE7FlRsGSxI2hnct9GKjyPA1RMOwvJWEdpKqvLsug54ZvQjST
yUwErrLvFyAgvrS0YvzC55w2CjuJLGK1+7KAm/EpNnWsEhozDs+/VibhD4XbsC00
phromndrTvY1sbm0NJSXFaXTDhcwcUbSCLRCE2d4C1CQXzbqV55tELmbYqRN669w
AZFxY6BsEpOPaT1ehZPpaoCuBZqC/Z8GiuhyMB6T5GrrWgWvMqFc+gVCCQQr2ZC6
5NAJUCVOyKHOA2/K8OsTGr/272UU7fAONKSfUiTe5um9B5FXLU8KQWW/Pg8Qc+/w
+Wm9reQlhaWClk3wTKMX025x/AVb5zwaEkDB8k0SITR2qwR9C17r2CIjwDcXVUt0
77sLZCv1cLLsHvSEy2el/SNNB1RucaV2xLy/1fJ3ARmyGxY8qO/Y3YqtPRw004Gj
178jXYLbLdM2iApcjM67UArUJMMx2ETm5M/rVRWQPcllbUgRJARjyhv9iXhG1q7A
eQhL6WZrUOAnZxI/uE2CBM0wFda+eaYhdbvtUacdxDiCWAoNHkmu+VvlrHUKBTR3
PLLq8zP7/Nl9znRkX0EvGBZkFwuPJK6c1yx3EhryYr7NN9KzI1Fi1/zkH0lz/XGu
uFQuFylGYQOk2YQIX1A8GboehqKdA62spek88bCg23TY2IPfIN0Y1pAxnvu/nVcc
36DthomYPKrK5eBF648oTJbDvRTsz5Za4HVxS62RC3SZZtjcQrk/Y0ZIG5gaexPI
lwcKLjQDfyzqDY0avOlke2ZUWSx/1uGWXybW2ZZ0hhtA1Y6pJMf8ZRy28EJclkKO
brOPsixN8gXmMOKM2ujsIoQudbu0xozkKuOJPQ/rWRM9X4aSkF6q8atIcvtuQRp+
PXWi7/oQL1Qs5o9WkThv5GOwKt7O6YCMdwotosQeyUQoUuGquxS/cygcsKK5Pu2M
Joivp2f7vDskKxKeW0yl1rx8lY+8LB1RKc+5g1uLC15GNE/OizWiOczo1MFIKVOw
4CbvFCN55nVkTMN71rCc8HamyU6dJRE9S3iNz3C9CQPa909426IJl1IB1pwIAoSQ
4qtCmBAmtPPdUZtGIw8ww88Zx5Tq4MarK7us6PWCk/HtSngiwMdLoiY5Dv3ek9k+
xxEPTDj7s55u2ktsuLOBwqUs1HeCW+KowBr08tME7fV+Np6pxvNHi7tJEQixlqn8
y88bjbC5uNRgtsx50DNplBFOlg2Mrv6pdU0tytBYkEZyrzUcNxYMJQH8J3N8buHH
BiTS4RMZ8nFQw6Ci82FtPMvjUsftmYG6F82vMAo1QpEAZL2kO/KQpp36b5p1WRM0
ZJlvO3RwmHEFS3aZWNezEGuTkGoG/kisDeWre0aP0hmPuTBJESD2oE7xxDTzHI7P
PpNoHvGZwPUihmhCBCr3Bwxt0cJfKM5NYmtNCJyARkyNOmxN9gR49RtzCpweY8Sm
fj7JFlDlwONqi2YUgzMEGy1pLI+F9zg8GVx9G7U9RtDrJlGQkOXFc9g1i5uBUj+S
11RZHeDVlaBEpsJZNk//jAZw/77ITb/V0e0oD6SRcVoZ5PNcIGTjZnHdI3KaEdIl
Z5qf+pbwQh+RgPXloYQDqka5MBG0S0dGCOukMspR+DiJblKWIUSDoz48on66l2uy
PjhDCy8X1aYWGR3OzJLl7Ya0imZioUVJ+CpUvdjNvoruUSeUDnVkt+jV8kZEIGRJ
HsjEgoV7TPOJsoeQhPfCYDspe6N2K8iGlM93TILA+2nI7MiMQjQN0d6AgWmJzHEC
/Lz+zvY4+/UTc4J0AeD75EOkWQzdlAT3Ya6uA3o7ky7YxMRlIE5ODS09BpFf4aaK
U+dBys09F92G/0ST9Qj6b73R2+IGkRLJqcBtJGDrIfYv2HXHgZYJGoDpuOO/EJhE
MQU2aQTVxdp/L/y6du9kW6Qu3Si2Nq2NRDraMZ5CQTcI0U9O+Za9ywEiRP+5o6lR
5rBiv+Mxyuka8FWM//T1+RyFgwJFhoNgf6GGOYXIj/r3niFUoVXGiK1aIf1FdtkW
Fzn40eB4sKkuoDiZWHOUWfJ6314DrHrXqHyTugn4dl+eFgHcVAQ30eJ+2EbjJzn6
l/4hDU/8U4iSB/0TT9TJZPNScQ+AQQpBzAGuOIWiRLAUBOCfxhi77q/yInELi152
+t1+1sn6ZmLBVTB9tR45r/eyQhb1sRDZWOgmZqbYg9LA4DU3nxIbp2E+Yh1NEQSa
xU2Ktk4zsJ32jOep5fXIj5+jHB6jeGSJm33UkhMPPOM7llFBtJxtqkUBNtydkmQ0
ONGh1uOZ+4QGjjQ0gef/pKn+RaIWSibIRUr+nGXkhi9/fNV5iN+QhsusRl4ZI6FY
thBxFse6gYqOgxDPJcWtbRRaXqEljXAmvI0ebJChsYif1bBPWrE63uhfe2u4vIlW
yqoyB4aIwxJmh5T9QNn2AhE1BWdjgJQHiB11enlzgMAcl2JwTpckYJ7TWpDIYY5l
MvU5bCzQdf5crx4jy8bugkP22UvGDI2bESGmAovUuK4crhl7ebirq5qtW2WGSNfR
rH7pB0ZwUiI+ODLemcIujojmVhOOKo5fh4KkD8A7IsfQwSJewiAEdMeCr9Z+ZNc7
KAp/sw11ScdOknIn+92PBgDq8gGlFk3oftNvIm/AxtVDCAQAbWxX/iUnxjlOmenL
0cnJLU04NV8ugs+XdP30K2Xt/SwDwTD0zSu+2t8zKA+KpvPOLzdRG0S3I7Q6BpSV
wNyBCz5iMyFkqDJ+aFt6eHViDkKFRFHfU5YAWLgbdfLxybCmiEBYUXH/MDpdCc2X
ojswvpZ8oSIEREKR9a6vSrESUqi5jcODPON/DuRFqH/9GVEsQX1W4ZS4hwfFmHKb
CHWj08oxdxaTpF5taDOHZg43kjWvsQcSKD5kjWxS7iLlUwMcSzZZh7+ilq+6LRKj
IH+59PDiJgX66aSzBJlNWB14oHZP2q69+vD0QN4N4cDQw6p2EQTOiU7LVRKzbBhe
FI0EiZNfTiv74drXCTNKsJ1lYXhYXUT3sXUEU9QupOsuCprX76BG/WOZD0OVrR09
5v4t/V6YPp0oinFBrWmRp3dZKUuZaquG5bGHl/mfdHex9M4e0/BZkWC3fJzFWal9
YHjLmRmDv4R2ELIhMv6HptVT82PzVlidXEqRcGH6v/MNYejygJyismd/iXfn4EYh
Loanpc0cxLiULFdOLtEP7I0JhbAqwNI7LyMfbcFY/zUTYCeLahRp6SzKYWhfijC5
7jbjq996HgnELnkJ56YZpw55yu7W8L2Zz7ROrO5hHXY4J9X59FC7dLiC6pQlVgmG
8/mYIV6vyQ5O2orF+f6ssoQeDNLTD4oUZ6hN31dygl8+9TAsasJ4716MHH2dhtql
FvHr68pkbS3pYuLxIzofw4LvHVtAKFsGg7Sab49WmfTjtqu3OYYCEM1jHcixdJzu
HwZNzc1KgvJgBatW4wfbRzqt3S1MVRpZ6x0bKRERVtI41qFfvQQmZceaR6Q/YGRA
TRmT3VweNdPH/zDYL2wbxuTUk6TjU56Oy0KtLRETyuW+HiNsNUHgPX2gN4XsvYVi
f9JiIwI+VbGT3pmuYycRWsDpfTzxYKwRm3D2nbX1vRpUG8YsNQIsBk1EKoMgW7SZ
F8aQzhJC4A1yoJEiIA6LQC17NFS9qsav2DYc6W4nOr8rRX1tD9wvf9Rltn3wisTw
J5NgZuxWeD7Qk951KSoP+ZVassjUHPO7XxvdZS3JcQ5+y+gQHUxSbwAtKmityJ2r
SgjM/vZLx9cx2omR4Sc3cYo5nUuABAiy+OlCcac8KMA/iB4kztz5Hg8QYfMn32H7
/63/Q0brxVJEptqy4BN1/yP91lgfffR4DESfA0U66voQZm1XNZsoEZzmz/0+mZZj
sORWTwr+W3dO44RRedSF64mqBqRh0CB2yWTQoXZPUrOwpm07RfrvYCvcWVIi+0Os
rEuZ2uzUvNSffEf02Fp32bJ906y1ZBx6d6v4+LlMArQupJHFwWIF3WhU/lPF9YDZ
2jnNc6EdpioNScYiPWdzAFDaIM4LY2NwR5vKd2GvZ05JL51lurSCUnK1LANI+bQs
0r1ZbEG5hX8ornuKZ42G7J1qQRdY3WK8tAm8gYoCsV6qVtlnlMiRyhfUTzTm2s5t
BfGUAJr0NFWuGhDTPkuCctY0lh0aQH/S+abwEOsSdvYv9Ri9a/FlpMaBistm1Ev0
yMe+8E3qnA9qPTp9YbIkIM73CA2p+8m27Zw3QYcGXYuZhluo1Rudvugyla4NrTwA
+kB1A4CL5T3YE34WfgaJMOxzBHbktOF+MJVLbaqXGwX/2LrOvEGBpNgDxM6dVtWw
24gIgsyxV89x+6ennB1lZUKgrfU0eBJ2lpPWp+r0Ri+CnrUbjVeEPXQjOV89eKJL
Rep6O1EO7tHLvVenJixNdPIUSPdtpYaJuI3i/9WTFp6T1hsfERQ9zSKakPdvKNSb
OesnfwGdyNiVHR1pL9uL9kINpJGozOcDYB6LOKbBF2LiO2vr2fSTfVjaJqpj1OuC
iqEcaXSiAzrNXFjBbbFcI4icxe69D9nyPn8NPegmuU8r021IrxvtlD74L3kpcumW
WlP1zzuSttdwX+HTpzYUiY/rrgrkSzglNfE6bKepXGIxYYvxQ+ypPMgty6jHb9hw
A5o0sCp98vs1yy643GU/94CadtBL+ChapvXgHmwDhI83i8n2bmtORjt4J79664+Q
PNIXGr8Jxz73MAIiXrp3s23kEZBo6Tx28p5oqHhLCbLExHQryKDVTRce6la7+lzB
IqOIUzpr3xxHhq6Kce2omvSnEiPzrj+hjqvpvWWQawhFYiedHfDHAU6mZ59+0N/c
7anqLUCmoHD/c18ns+rwBPaofwExgbYv/VbJZfzewl/uWbbYgih7SczpmUsJy+sS
kg4ps+u+ZoGbTv7K8q+Ieskee/CRQCgsZWWgPb0Njwqo0zeQ0hqTcLV6hZII9Zit
dEpXsfJkp+msQ8JTUAWRXl1A7D58FO5PzG6347qhk4RpkoF636qc5V+yrh2zbiX8
KARS+frPkDnTsxLFMfwuRzIy288zS77VrhBHm2SbgRxpVRhMGZ3eCBO4465fEhG6
YKqGUIW8N+thfuolYrmuQxc7XDgB8JJlYb7sRVOUgVrjWKKDsKoDWTipJLeHnQmO
kj0tgtSwGOj1cgw7a3vnUSbTpGOSlTJ7MSLgr0dfWzHC1nYAmnDzYITOFS0isPiB
aahDh16q4Zdes773dVfuPohHGbEdl536i0XJ1Z8TAr6xiqD6E6StY0pEIJj8fheW
KcXQPpETZEOQbfev+pBzSMiJdhh+jqf13xygMT+F6ILBBMz+Dh1IUTajyTb0qSJa
20MHvk7C/zNnRrhGy29VdkpiX2bmNaaMpD/zkNNnaFwVX3+U0inW5guBqhKaYL6+
WkeWF8xb63RTkjx2EreLPtwJobclV6bzNuOoeRj0M8dX90u6m53UAwyTIkVg6QHn
KVqQ/r6c0BZ7QFLFlMMRA7p6n0T9+ves9SjscxhOUlMFmQKrjxmcyqmhMYVAqkyV
+jCJZQdZOYrgWBdcwUsMti8QdlaMZUYIbFaiBBBCRPmevqvcFKv01Rw1rJGuAd21
4Rsf7SyFqpeDC0tLD0GkkgGZW/iOiW7ORxHp2wyDvwa1wpOowf22ADTyq4CHhjjw
8jKhtNh/nsGKdzYgcx88BE7RYYKw7tUiiA/O58SIuItexYE4Gn8CuazlqE9AJzSq
RoJUyB1qir422bYcOamNMv3rWTpZYLOc+A3rx9t4EjP3SuDN+yMbHe01/AWly1Oi
He1VaggveFEkAMRuUjS9LbGGOJ7DAdDLEvLTXXMmg7GvQ3xY9WeI0Hb6xemImQcN
sknzYugLqSTEBL08+zv/2bmXkdfIWtKUP6bdDFl3Ysh8EMG2mQJfHmgT1W1FnWBg
p7t3uLg/piUzOztHYtSUqilQ7pyUIBUFE/+C6aMVOT6vyi7nYF72SMcTPkKAaSH8
VXwVMnesk1iMi7+Rahe+39uTVYLGdEPDhKId/5vUIKlzK0VFuY8qNFROuaKGy8sW
QkUjoA0bKiEeMZtOHLBdUrJ/nNucOFob/0PqcIiytiPNDFtqHNlZpheFN0D9Bvzu
vtaC92SsfCMJCYIBnPLkoxQW808/KEG1LX/WfDK9oTHSxGYpTfz5UQaeV/brfInu
/WgpAvcVunVrPJf1lHHc5Df2WU+NlIzto0TnQb4takC62LlIcTTsD63oVLk44vfG
UsJ4wsKYEDBN5DaZ7fCfL0kBB5KiIXj1ACGtzUVACWnfJFDitJYuINLnBezBcRCc
eRRSFhuIPp7wN2Rr5/RxhsyI0w76Z/Lk0xTMgAlw/TGRWsrlseLLh7j8BHcj+BML
gZWeVOKTxcaaAC9+AWEIzrY8D7fFTAP1fGoKMeUAzmNAp5YkEwIyhGe++g/UP8Ia
1rJhTPyozcrzvOQSRSt7OanCpg5ptoiX2Mwb+w+FpcbScmPV+KTF0mGYykdnolvI
M0qTzyk1jQMoXLioqRotRxTZVgJ+pmGSYZ6UumIY2Zgql73e80ykgBN4uxKgAVCx
/a/dXOTwOmyXGd6dH2DD0bXBearojUtHB83HvuVdVKRy/v1Igcqckjv26YwwtQq3
d1zDE3t03QDnjtNN4KdHStZXMz603drmiCdPxrueIB13P758gKzU2wqWdGAh7tow
NRErJrVzypcJg1pXNyNutipOlSFGb8vxN9+DZZq+XK0tdToOsclF+qDhFEFiOiKn
GS3BZOm4JRo71sQ8/bXOfOnRlBtcOAY9KGqK3HCO65kYdG09W6w1XmihdQJrx9DC
Spz3TTj5YVbizXS6vdGGVYex/cgp4EXOJuWpLLr95sEf/eJZ2vVxmDBb2ceWJ2UN
wvB6EStnhRguK6GaRw5HgJ3Z9l2x2VUttYl97AtX00LBOUkd4M880kKLHuyCLnAA
bj8H4ViOWJtCqlS1Qe29p2KueiL4W204idqK5bfeit3cE+zYEpHdGc1e7F9iHwcL
/H0ygC1tjKfPtpWHCEhdlE/o3Grko3sW3X454WCXwZdKWtUhi9dILfDOEY1H/xHM
44HallWvcH8CJqU+XhVqqMAaVOkCBQw4NAeZq9YsT1ZBZ/yTNsky11cm+0RpicCA
dSskikTUvapvkwCenFTFlVUT1WLCKSHKIV4SbfFsD17CC+GaGNddB9KkEIWjh8Vg
3ZvtICFs7RcNSjOPgBs0SNfRDRLXmiDIWJ2owd9AyEaWfxtZwZif9bizhm3ETZbG
lRuw3cIf4EAo/5RgRmlJbHz6TvrfO8CNqBZqgXzOlKP33AO2C5CpN8NOOuk1WcWr
DpDjX8UURX6btADv74bVpixlSqu5slOsMeoJsMcaG05GBG5oVzdgESUljuxCzRyz
f18hajl44akE/Nzvx3ufKFH3r8pAiYnJnCbU3qB//f2GEuPLttVdfvR3PTfBjOd8
8TTkur4nGt4rdOH3fWSyn/NiDb7Pr98JAh6hHyi38fmzCHIifmCiYbA0TgpiHjIg
hIZ0JbTXhxCWFYvrNCC3EC5acfAQ1uGUJOVtdfUOpEOb9erujzB8Dc1PxcTp/f6L
R5SlgjBTqqZb+7yiflIYc3wCLSv4HVh7oVhAquArv+Bw6XWocXessH1FBHm+6qdE
T7yz0PScigOGZSAQoqp+jF2LxhYKWNxcafNgpR5l5TwzXHWOeW07DYtKdGlO0ARp
mnwxD0tKFZJNopkzXtqiOF7J5cQ5UxZaxXRRf409m39SUTTnm2NERY7RGmGQqs/e
QUDtm1nIytyh+p0binB+HqItxC0Gf8590CwxvCGfVVjO77EMDmwNkhUn5SxAEMft
WctX/TcbAJsCxUDDE7L5hQhv5zzXx7xRvvXOHb/XoUKr8bCGcXVQMb4WtNVcvZ4t
jGc7zXTDz2Hg4zQDCqBxVRgUVrOhJ8TJBNw6NtM0MNF/RlxYSoJOVSwERF7ybWZ/
cpT79krmGnIkvBg5rvbj0ngZ3OKK16rf2AX5D6x9ZcIoARml3aIyXjpupV+6e0hg
rB+1T2UwQB/h9F44/e9q3ZYC/uPcXUISWBeCyFXotMdq5DqwSsJYpV7wHeBAZ4mQ
5RMN4p1lnEiQXXgBnoSNST0U0teTRyQiAHedV5zk4ShmPKSnIlknSM3oC8nJUCFl
GoJnlwLKI6vmgTsXvW2UqEa3HW/OoOWYO/mvhqdhmBCqgTiLaC92micUSn8fOC90
d1RISNlhS0cIPvfGiTLK3nmyQkzZiZHNjZ1LmZ8wkEabftkH6tKgL200T4MPvaRK
NOImr8OF16Dyb1TgKQ9gswnTQaqVVxXHr7HuM98lqCDBw3Y0jSjUrB+plE+tCAdu
a7S0QVQZrMmRyJzrB+sO8rPkyxuhx1xML/q+DsPeyuf/CE7XH8Pi+3+G56XKU25s
PMWjNF7PAJlkTosxk0093Q+kOpo465XADEJaFffDIuynIQG1EdtFD4xUBB+yLvii
jSFRNl1XPhtwb4Kf3klD6VyrDj9nI4hk0AySnDLQWaLUYU8y+oVQ4vh9PL9xkI29
7/GkLP5ZK52dm1ROmp2lxuXhSZIt9sW1k9wNRl8iOgm3VYRwlUdknLDYqh2Cx7i1
naB8YQ+K+X6EUd++GeivY+TGUoBz/VbRujF7rAl9gID/36k69MtkW0mTo4IqNQJR
lOO7crhqeKMXJNOLz6elnkZH+INm4Myxein1W09PCwV1dgcMFlqFWYi819qnectk
j5X0CQ523GgV/2ccrP+aU3amPFZeaIDhyA5HM+KLJ6r+QZvRem/AkW8RIdCKkl9E
tqE6uBzJNT+KCEWRFToFBMznlZDUjC8NShjkkbb6y0k7hLfTR6+c0o+YpZmvu5ig
sYhSWQeiXajmef1jaHbCNnFJp1X0pAu3AYh32t6pTAm7cPKOaIz9cLXKF0Q/MS6S
8jozG1/EamCeNRVmxmdl6+ifGe3sgxUF6OcEgi6ILCIuq5bSqok5ckDmA4Xj7BC3
nJtW65ks/e/PUXm0yvmuBsI0fW3xbYwcM9TxcPg3EuUg2X79ZuWoKfCDGOFaY57X
OUEVKssB5My4Rz9y/wzT9P6AjgpPxYeGO+tXbKg8n6IXYpHIWXyTB+0zoZsVUwP0
niveRHX8dR9WEA8ieTt8ctw9nQW83EWdS/yzkzUiiiilPiexvZCrKq3Mt97wXLZs
v606RqJMn8mTAkjLCopwEYqa8HbPIxowdNpHh2ZQuak/Or+CAShKV1s0CmAVtep/
BGM9C7AY6RRNEr+g3srQkTHYd7D7qKOeGQzBpYmjhH1mbXeEDj9/uXQgKg2zOIIt
m6n+2ZzK4B+P2OQPKyQlh/xACfrZefaO0NyUSEyi5zZt73FyvozAwu0hwo7pe+p4
jw4Lfwx+VlbeteNyYLLCw3K8HCyQOA+JwVuhV+jOyc8cReeQeOCihh8RtkPcnFJ5
wB6peu6+cocSNyAv98eYlBkw/zBmT3tccR/C8/C7xoh60aExk5g80yWwOgpF9TzI
r4tdqQ71ER5P7mGXdRnCmldSR20d60mZHo6iOCUwbNpXHK9JNMNQPPTwpv6IfnW+
u8pQZJLWo7iMGRBxhlBpv4NiCjAg8rSZr/x6yHtnORcz17ES6tFGRu/I0GqIcoQX
Yph+82aqSk8SFYI6j6NxBu4q/3oBl4x4WvUg/yRPjFQ=
`pragma protect end_protected
