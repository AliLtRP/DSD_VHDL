// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CplLCfhM9YbXZOIe3BkWAmAgA/4XjFzm7ZFX0oPmXPa9u8cxb3IQzb2iwlHg9iTK
N2Q0Ehp/Hqm2NJiqOqJtX9LTTsTdl4wq8di5UUlMvGBbpjQjpSDpHjRgExq4Utjj
kIAzf7jK6MOESjFI8wNj0reAnAQGdLhAKC+H+yyY8U8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9040)
ZdrmBcOLvM56Jxj3w3zH3YqxdjuHP6rsNwY4vpOgmvtw9YWyU04BPuL/FXNszIVJ
s1yf4dLtYHPKmY/euK4vF6sE0BhyC/76LGgLzUkZdFhgsE01HAzbi/V9GZVD914t
Bxyv8wMNYzQi+lU/2U+go+sv+EXDpUkz4xTUB9MLhkrUCoxmWvg1JNUwnUSCuRSJ
SY5KglU5a6xJRA+O4jbm2av6/6RkOGSGkpjBfPSr0Ko1h8lXJUDzYPm1qQq8YU3e
Uxgdtkrn6zS8xYH7cGlwBD9DCRIv1DupzXLnSj7/W13HYv5A0p7rDyFKAJzc/4y+
3iBNrN5nuBKiPmqqU12xTUVCup2pVb2O6X+CexAM/X3MY99ieR2A6+0SyYb9VAUs
B78C2c+QwOQZrAxDQzrpzkVGQ+16b4ONTdnVghulH+9zMt288ZtV+WWXG/9V/oWd
NbnSBUUNQmZfkCABOGrGhpWzl+583tzRQGVTXr6R0fQB47T3T92JbkIgiTHWrGxD
nmB+/ADLoF+GjgW3fTWu1oqb4XELa9C0E/jcnWPQ63QBvwNmVADmSueCvIywSK0l
cZ9u+DD0IJaLILece96SYIiyrs4i6RuFNUGEgTOyB4RwiBg89wlsE4xRLUuHeOqF
lE2FzZu3mXPYgyHCkno3AJSNaVf88u9b+9hzwB8yDLIxr7TDehIa8nT2sDdALO+6
s4REuv8ozS4dO20gbGfO7r+k5iuFqSs01rxuwk+ggjoGzY7fTRSG5SadQqACnaxO
nAhNp43G/gpfc2KW8tBpVlkdQwhn5qZNQgDsUgy6H2ByhdwEY2JzvtYOGhD0o10V
nkV5rEoiExv8iUKHDs8xpiH9qvybi4VjpI8ZpJzPXE2XOGCjoN09/H+0A1cysSgo
VVs018a1s6ppSWeOVUkjmt1AIiI0lTvMIGmNEskKfEtaWMG9fF4P3Hv/fD5BAV0a
Y6iEJBFb35goaU3eHks8lS3GTrZlRfi3Moy3DIxKTIKIYEeGjNOiiLhHwHxpS7b7
uD4SWW2Q5+ArSfP8Cgv9hA1Op4PFVYze2sZZpy+1Zga3rVNmwU7EizinE3P4i1IU
toRljSpAi5TziaNr8RWD2g975OpxofXtOvaguIH8JYERxkKMbeWv3jNn5I6tuHlA
FJyMhAWkvQHSjOkUtlXgpl2ofzRzU7pNJviUNE729ALtQ/Oi6y31lvwOlKgutufU
IHYIazTwKn0LUR5Bo93az0hXacL2WK6kyTSsmieI26D/uK2DGbGoCIu12B2+z7VX
Kx2DNNlN9neE0VBYpEBi162aXCEJ1/JpwSfQKERhPxC82P/mDL3g/n1aNKlawwGY
4hNB6rtcTfI0CV8yD7d/2OONV5sb4Gp1lvxyTgtQ3XNYyG7LmZaC6r0Bwq3rBJXJ
WLv9Ne6F72l1P4eAOjfiNGoO+z12XFFf4LBn6QitAAD8Gbj4ipX7GhVibLaGCIuG
Ue4coV/6SpIpYe/NFhYIuXmAd3FcYva7gxo2pK3wFHv/l3ZpF5qQNfeqM+dexSr7
In+OqT5URdZeB3dU55xP+cv8u4lYJUR9h/Tc4sVxkSLBzyV+08pZfNWKrWG4L2Ze
MtMDKIH5nIJaCNw9awlblcIvl9EyAmWTCNjwlKmaTJFDwLjBZ/pyJ2WsYAEbBVHK
rLqO0aZFMjredRA2GLAwjyXA/X13xIE9ZdY3rZqE5R7Bd1VFLlYYhYTRvImtL5uE
+k3YhvyAaMaBpL1VZxHds0Y32pozoo7hzvNuEr3/M4wzcg8RVEBz3zEgt+oepTHf
d/OLWkxC4djZr0jflfRI5e2kZr/OitVqpM3bceF85Xn1BH7uXtUwAcYBfAQphL/q
+N9+Ggeg6AgLMerG6r4TCl8MW3VYbq6IOI1+uyh3INCSHeq9acyDb0B3iCC3tTAK
tlUnKMi0LxH6K0Kz5zOXWgLihvkqcB13gRdsQoNGgCPheuK3nRv22djt4ICbDXe0
8cOwZoEun7ynHYsuVmGAqiIQtA+K6PFUk2eny0Jiq9+ffpLXy3Q/lowB1YOB2NQO
7ohK9DkHul1FmyZyOB7OAshL3YO5O9z5WRVWqIGqz0rgQoe2/TXxfaUg+xY/GvTS
UpWqbPUvBkOGkKJFi9KQxUaNnK8KJB/DYPlB9JDkhnS33GIYYpFZNLUibLryg77y
3/U+KTH5NuTKfUNfvfjNT6rt1Zlg/7I28aaVxdiCfwl8H/IKVphzPtIFP3M/i1nB
7NWEqLjiC8fonxzXtX8xm6rZCilk3I/2zfTcizN2P10SHP0UOJViDCF9JdbBvQMC
ocBwycfp9NCGDArqyzSnUp24yz6s74kLTLYSJnGJB+2w9Q8vlmUiWbcR/bl0ngM5
krqLSPAYYo+V8BGZNINXwMYVOC5hhY+44Uw0kn6mYRs7ltbrNmVliG84KKL9d0g9
SRbxXXvWgBFnVnSS0NckrK8h8MNl/1ytppJBvJ9IwUONvHeYopRpBFXNq4mDTL64
WQw7MKG4oDeQ7dt6wkfvHcX9ai6R0xNJ8GEMnGBKNLAECNBBQCBCZAvgmi9emWBo
b5khIDCfyFbYjTus/+9qmUivq8+5sYRv0rrZYcX9ybkQT8kCLu9eg6k0t7goAnvZ
SOZHEuz2N4BqgODA1xyoRuIyaWYB48Hwu/Vg4Njru+rZcWFqMBJgsV5rKHBkTIi/
HY6jlFVF/ViuAUuyAGt6JtSd8hM3s4Ll3m2dKr/t0x73UcNp/IfYUzerN2B1esOn
E/euP6VHFv+l3xsOgJOlAmQIxAhK9efGWyk3eYRyZGqxKisOUiO8dfsTIfs5x6tj
FP+oWb/sdY3ITqFkDm1CARBeNx+CUtVOd4+2QfFc4hVax9C++Je1s7XoNcCU+8yy
hrI8QmUObQy35tQxerMxEpQx4jQ1GgvA0SjHNwwYrFoM19ZudTWtkgWhPcUrXZpN
csf+qvFZ9BnXiZBCnZHWjZM6/g+YAu+40s3IeNwTItAsSngLgFQHV52ByT556w0X
oXuOo5Nr+4/S1G9/7r4Ol1elf/Fu85p5LbB3pAhodiseAa1BVYAhYDBP5bh5gKQZ
8K9Fm8DzJhR+P4JicPF7kmGF5MaSKcgbsWWe+C/0GMeBebEN+JHQxn8trixaFYU6
i1zgqlSw4nmNukZ80sMiooz4z2CO8VsYd3AAowBRDu3vopEXsl5rgkP05bUl+OQh
++DWwR+w2yQWWMrSTEyWLdFVHx8m0TWzp7BB5kNQqkcX6P6CLiVbQh2e6ViFI/Ot
2M7KBZwHDyC/nAOhL5ssx4fMK1nvgRIWHf3OPUMSw2BDLbv53AmyGXcXRgwh2jNW
29y0t4s7ZpAyH+9dzEJmoYDEmi8ePlkiUHXG/RR+l5CYlRz7yOL0ynE3TGcocsaj
se/LkgQ6Tgua/qwR7X6E/VERv8RCJM830sdbBXPoIxGIwUgDFqPJuc3CQdnVK3m8
Yj3B3frpuebrtghpdlnq95OOZ7EhFYQZVxTAnXQ87UHKlQkFqrMc6NDP6M7s171l
2kqMHwUec8GoM83Qtu5OEaQgMlLwZuT7221rH2OJKY0zzFWvXo395hg8sKOB3Ld6
aUwqU4dbvtOsxYM5BQP5iRvlEYBKEYOqQVDpWMFFYks1OixZjFc/0WZIffPuclse
OvrPSyJ2uKc7PPz/vWDkRAAxaznVO34s+DWJojbj1IPnoXLjRw/L7EjZKsQ8EFUw
Cj6X3ZSNtnBVH3OcCoBGUyEV/f3GHYTW6jC2WbvZEMPxVMBUcZxB4mIgdhFDCTOL
yw8WdhzTWlUU7wWDRP5CAft46Z5wKnBIZuZrpe1L5VgSO89DlQH2yLeWcs7C3R7y
gXTN3SVzAMsiJ38YFx9jMCidcLOXfgiggCKcDiUiFX03R04KJoHNMGjZ3nrpAM2i
IjPDxfg21g9lloYSVbFYI2iyV4uPRZ6N1CwWo0kqaNttxE5MsbXN6FD/Ks6Ww9KL
leg0G2lw8ohyby5gyqIa65A/ZemKIWz7dJryUGTaEaKbP/lCl6VORIN2mFubnw6n
vpkOnvlRbnVGZz4+TNQcgpm8larL3H2U06ll39bhZEYtmf0dQwq2f8rpXDuqpOuC
4x/8MeuJkoHeNgNaJFlZ3i3bIvFFtsERfXUdCOfDO4Es131dvB874Jq8ON0RYWAB
cMuiHZmEnNQfA2zJ2HCLxWQmetnZ6LGSg266ypTuO4fn8rWu8/5Fr21o9T/fzugT
bcaI4njE2+nzD7gKrKhjl1uGBympSRNqBHEOkAyIATMoiVoL529wO2UoQaWyLEKJ
bKRKkNnyzys1wha6KFBv6KyaPwSkQB1WgZTJM03ylsach/c6VjtiXCfPMVXCuUeT
2GNTRMNCE3uFw+00Uc5offe4y4KnybV/AgZURqSH6BUKjnIlWkNGxismrz+0OOy3
hES4wJmMYSsHjrovUCNlp3g0qnQL2wb/Xmydzr9p5j6iUi3U+ettNRsYc17BVnCa
Lfxq49f1rYRYMlp5Sx9/E/q7yc2eaEvMvXDuIkQRF6AWnBpjP2gAgcTpY0QcyR2z
PJ4hgP2WJy3X/RFzakA9s7fa9nm04tN8+/jn9dThswfjzoOAWh1yKaicuTfuGrYl
l7usWIp2nqEtgAES0iwMhTeIOL7vM4EuVQRrrxZgtCCvliEhUZT1AoXmZpgJ3Ztc
b1dXmSC7uJC0F3kcYgn4kUmiA32KsKH64gN4kWtsTjHjiof20uNQ5jXYAU8JNFDH
8gDmarFdCuFvDl/8tvjs+OVNxSK1afg/FZPShGcGVY382IQJOK44RWMIjOaV1v3B
rBH2kMaF7S5QnXrL8Ilftc7ZnudwH7jlLIRYptquFXsUJZWWvaerLh0ckq4HPZpl
pUbXtIvUp+8xT+qcian5FXl4O/Ta2yRqxcLfOniPVy9dDnQdGlMLmOApJ4ajbggm
2zaIWk6nGMPYMsHXfVaSqy4/gjpEHEW1l9pXG9tUdxrt7iE57PvNRp8dxfQNLgd4
Vn8URr/ZUhb4gC/m4UgkFpzvUjeATy1OD1VByO/L2kcCwF6VTA930oGhUjrafGPr
tMHSP19H5IO31aH5jP3O6JBQEERgExeglSOS/J6q7FvA7Nz+x5Xr7Ny/S0X1+w+d
gVqNhI8ul3Q676v41+lpm9LJ1vMDw/LxlUzu8Ol4tiPPS12xlF9dKy6X3FDntEfJ
3ac4Swva4yHTfRlPJH9hP/AL4Tkl/QhyMP7qrqMYbAZSsfvoTmTamq1WoyZQS1wO
rKDDm9eDdBkuIg2OrpmJ/coDkbC3J8AxXbzEMZasGjwqJsd+d1ArAP/5JFwgxgLv
iGH+ll+LWLMirse76EFaJ/yHoS2gt3fTDhocUWXa3iSfQ+MEwvcUXmlA1PPrEx8b
aNvxGfBAB/swcz7xE7bfTJK1N5NA3B+KlAi415VrAJhf2T7GDv036iPW0Xd8hHM/
KaxST1DaawqPLqd756e46RVot0g9EnYv8Vem/8waiF6I9QB4uQNkwV/vEp4H9tpi
b1/4b1jKJXYK22JFdbH2mE0f8gxkqTaT/CVYfZst7BLdvWG1IkTAwkuYFobNqpEP
qPkzRyjPN2+LrfHfJNcB5OWtWCCHIayzEHkhy+g3tC8TrYGwkPaLMKPgIbNK0PQG
Fg+jIqDLdF/NCZ7ZPJe9HMHSXdRaJt2vcElfqrJB9Dtqe/z6WbE3pPICOjtKlvCV
/fgLGRjVCso4gIRwDDLpRqc9885JJranT/RCUjeNQbGjbcCzL3GaJgly9dlV7/KO
zNCAipgLcXKgDNao21sGbwN9eLH8bSZ+DTU77EdSN3NeOOJiStlskUAkpIcVb//7
CSj2i5CRiVi0IkpE/AKH//rXZo8v+2jA2NzxAozyBWWkKLCei1p5+ozrYpY+0vMx
HwQGSbYQaQXovG5b5BncYIfjQ6yL0Xh4Mw6asrPJ4rf81khPyj/654SB+iRyfU/v
nNRKwP7D7miSOrSh2DBYdfLFg9mBqUhaxJMF54hTb5IQwjBUAC2ZveHlm8T0x/aP
YOWlxeJr+HALRwqQ2bnnJM14XA5Wt67nUu44ZquUqfXVoS+8rZH70rHobVsJ8XxN
Zxo4R5jT95Qg3q6v3P2FIcXdTqK021QY2CRkHl9c4HD5zmVz05gUex+MR+P2Rh++
Ou607U2iHLQCyUIvSu1DEbJz4u16nyDHhdIwiNjljv18IpIVPJJE2dz57xTEYtqH
+skZymaknvICZ/cWLdoEYRR2ViUv/+IiXpq8se4tHQbHyTTZLd9+lwBUqzU3t73y
qi6NLfIuzulIHuo4JnYEAa1sKOvFnk/9/AnvOnrai3rAEZErpFknzkUa2ulla1hH
nDqXQePJZKAIBl5GZGPSImXq3wSGP3p7eJ6p9I0syApIHQgzPGAfOvWqhtlksjWl
xU/b5rRDHVTtPmMbpu7UyDWaxdahKm4zsNg1WsrZgRnY9s/bfQ2GJtixFO6JqY5w
xuWKtqBDtE58aurgwKvlqeCnuWsAWohXT8LzA3S+0u8II44OVEgvxHD29SEUUBlp
L083wjAYbCbaczHt40PMfQl/ipcI3Ri8vyKCQ4HOgzd9AzIZImKdsPqoMgLvEddK
EtMbFhpzDJSD7aP7jsl7K8Ojchto/RykiZZj6v/n/MDNjAPxfgjgVLOkw5Cxa9sI
iXm2LX+JN7Lr9pO+fFufUjqMQQBILJ12BQFlfKxd8b5hsn9uqbpalMUfvwzy7shx
wnQtxz8bs+jhMhHWsp1Nz9wusA3DddQwWMdL46oPnpPJ7un/3Omr+RPTNKuF4Sq+
rY1LzbhEJ1fEYLYhoRQs97KwodyPhKv+rRgz6GlxtBOAQEWjMWu7KmHcaBiC49kk
+LYMFeJ9RPQAymTn3++3sXeRtdK4gyxraQqV+DoMwRk32PQ5SfexdUcO7Q/O5rxq
BEE42/rUnbnjHXrMqOHw69umcfPQ7sBn7MVUFrV90G34IerEGNmOP/GipJ5Iu8dq
OYnIJCmXV/nunKwvWx041BvHhQ87bKThoxU80d8gryBAIPAdyqvcTlVWZw6NJckl
MICwxLZMfMaXuGKYc57VaY2bFfF2NIhQ/lEmF50Mmf075efHjLSIbiIalzM8pDfd
OdbD79Y5ZRtQMsOzd7y9O1cG/TqfuXdb1pVZZUnmUXY1UX/NX1SgYOIyvYPKSrTk
GNGqOg4gKp8KxHE3DoW13gSpDNZoru6cc1a4iyfSdb1Q9ovqLaanMPJjGfd4Kn9j
IyzcUh7TanVMKuZmPtjtlEiK/p2uMRNXXY7Gwx+2whQUOCpZy+5ZobTojNHUHE3k
Te7iLUhi5tEbnZTkj3wb20NxV9ZGQ/X3V2Vp7tAHOrrHSDQxol+YCOchNCcMjn3u
H31vi8pPHGojFdzK4ngOLgqmqOfboZrp+Cki6/DUZaxauOAJczsm1TimhkLE1pCB
irYowXiYxMZGCjT/RxdDVYp5tpk3URsZr2FHQRIZzxAVoQr0U8wFbVIU5unT1GeL
AjpvJ7ICe0zPzivfvWJGLTvih89foZybMNbs5WnUBjLJFnypC0nPneCjyZdiAWd0
Him2GFQzLmXZI3ztRkv6G8wTY76tUnaxOj7prAx8PjjYcX+jiRhHlv5JvTx4VBMi
Vv/IOpGrQ2EzODTqeZoicIKXji4orGaiFPGUGWjkmYNyGn9YbQX5ouZwJVNpG2wY
QnL+v1v71PziKAAxJGFsi8acsTbDxSHNJGyodSbZGhaLIWPC/v/Q5kaV5NW72M7r
Ir9NKhA/P1syk64nkBeRAzXU2O1yGAWh8EdfAbpQclhJpmNsrDVqyK1txzeSojk4
pjl1XQPabsfnPqNUr3qriJwxfRIbA425rXUdyYHgFg7CyNrHYK6AIwf6zl3GOuNf
Vn1IHFuxtnGWUcCQrlRnZ6uqAEELPWbte7fSq+5zQKzBbylEQKTIMOKnBBXZ0NF3
/KlbiTxriMtJ+hOef6cHsGWjtBujesE1fngLAwz8h35Qv3xsawX1dk3GDzRfY6ya
AtRfONqAEqCAd8oqKaW29VTEdWjjn/iXnn7HOtChonxqjjMlW5qKWN2d5gOhyiSL
Nc73CR7MOVK8K8MAa4rXdW+nQWuraRQjFnbS3AGDVxTFzs9hpzRSJzWAZW/e6vbk
D+NIeUVxe4Aq3k1ocgttppCNLsPaYNFD5j8gSvcLzF5360RBhl3Iky03qMCAyg67
SbsCQAra3eIGusa8ievIt1rIHb0cFIvQWD8WHmbvUntSHmhNiGiJQ8Lp2f/AJtMY
WWZEvNoFSG4NSeOB+5qxCQJ4HoVwHawtPY8WV7/VhPCivS9M/VgRJe3QdlCHv8vl
wXHA9gmhuOV952A8HdnFo1IG9KwuM4CX/dK/eSSYNS8HYe52y5hdCtcUYox2Nqyz
aCNSGbf1p0qEExD/1g0FucC7OzzqsOvULW+G9TqqubhJZd5aFO7ss/Da4ykPdhDD
1xdHeHfSGIv20pVQ5MmHm9yv8tkmZHFLOq8b1Ik6pyxvPW/b7L1iOywVJP+6BiZa
gVXzwJL29X2e2cDNv138xS/NdqO5MbnGTONxqIHHukH033Xa9f6wK0jWb5FFoOTb
kvFoZfHFsYIhSrag3mGwp5xnEl4mT9kzsd/1W3/GycfL4PofZNtXSr24s5Lp9xnD
QozLLNO1WEudtRyPfrZ9nEfzMV6Yo6D1VMPAFVegs0xuhfaVXihwwd16yVtJvzFC
PSnaCZhQMAI9PwjAam/glhd/7I6PmpjdOyEHN0CJfQ0XoZ/EV5K0/lxKn+UUEsq/
MiZ2+BQCLSGAIeU6eZ/YvdxO3nBoEjXwFFOw8Md8Zow2WIluUb1iFDlYXfFqKAjH
nSz8mKBL/32dwaB2yFI3P0CQUJ0F4iZIROxP+wmI0UI74PDTRHdNHJcDDHv6piyP
+QSZ/j+dNWj0AMtDkEqKMd+p4GpmdHSpS2qNi/59B/UfefZgXp4oynw/6QyY1/IO
2JifaGb8F/7FHhP19vLEU/IhTwCZOlouqhmtLlSBEXKDdEz9Z9HU7zQ3N8P1H0Am
k5j4ondKfjfGZa+DLbTt0LEaJV9XPoPDiqvYP0lXodw2tvBrzOVns0kp0n9kCHTw
qJNQhTpRaTeOIUtIJP/KFMb9NJIesP1gqmeM8UDbZ506mLbyVFfHgSF9+PjLlO78
AmfPhtpjiViuZAyDFS4gaVIbKViKhsg0T/g3h6X/XotFBTsLuU39qHDf+GLu6n50
LRtUNdUp1X5wjlz2xayyxM2iuS9Jlb5786qr5pVCzj4jXUiIy+XXxzSHiMzDynPI
9633ycF3r326/K1U4RkYd3z589o6HCYmsddf5dmih75IMwdRyWf13o99L4+4qN21
sl4SpNRwbpJXBu/g0fMttwkYPa5f9M52pmrLmKkVfsPvGwGzAdFvAOwERaULcWgN
tn1EzYs9B0rWaWAwxPu3gxHth0SjQv4rXRFU+JRnmmWsEVNHF9VElO2Wg+V3hpDA
Yk04T/DwzD56bGem3YV0WZ0LmfqGi/XxkBcztOI5167xRffNyYbVGAIT0vtuWIg0
faR1/mIEewXhicI8vQoNcyrYz7kecPj2VcYwZQKGyYmL9Iq/YqcyTuM/oX3O2zq+
Eon2M3T4as++Et4ueRv1nXAPMnJLlPts6e1OKaom1zZugXuoSF7waDL2zyf6vk9t
PlbMw805jRXZo2Dz6wMWHO6csUg1+0W6AFsaCW7K0PejKPSD03ZV338dLo0cCMc2
UGhkKYYyKiDqtX9JUnbdAla1Ep343Sl2W9uqbMc/5WA7buwLWNtUt/JdGneZPUUj
e0+J1UrkQx0cIlkG028jJULg/OfxnC4VM0lVaNhxGidMwQZrCE12yAPiZrWO0jDU
/VrnPsxHhUX66cj8dNCYEJC5tDAFvHrdTjxQ6ROFWO2CjCpokwI8SGIG0RXHjL6n
2cSAz0zflL3K8AFE6Jowq1D7imi17TinizOs5SGcldWyheVSYxN0zlTKAxZ6xiV1
BBoKZOlpo1LeBcpoAiftGiZ2anfX0O1UNKlWXXoRA3tHV5hL4FKYf8Xwf6ZoP9lB
yDUyp3ko/yjwiPAz8B9b5U0FvKUfoQx2EYSRvRn8QBRb80Fl1aYYTHa7SSot5l4x
aLzZc1tivMXMKOEF5VDpInlth9dxByNDm/UiHVXsoen7eqPM1dj7C0EwT0NgWiOT
VSEexxnfuusFZv0dsqN8hWsZB6b2inXphIZT+VpjAz18xMsKLYSIOXK0p6/jJboz
j3kSp9wftpcWHt4S8X7XlnWXssp2uoCw+dQWt2Zh51O/M5yacK6ux011cWrNylKm
iMeCaSVUrRQpdt0ga4q8jUQ/QYl34B4LIX4HYdG3UTrA8EnXBLa6XWR+htKW4e8+
lA2VE+7MonE+15gXPwjEblOemvx+eQ4P8dTiSNN+v35DxCXqNtvUtwPykeKYJcDw
6+A20VmLd4a0AgOv+djCreASbZW8ZII817lXCLm0Ugu6Gj6YsDm2endXScPlqxiX
5u/SeZjgCGigaQDLNZhPfG/DqgzqQMYn/bswz40rEtD3TAXKYQrbIX8bzL4c4jly
jnCrVVDNSwvJIfe0IHnDM2BE9hPKrnnpgJ6cOWYvkWh8VyJ1Nw320H2wyw4po/LS
dijJvyzU8gfiN7DejehgtQ3XnRdyMt+n+FB1QuW8gUkKA39LTsu0hw3p/c3lh2Z+
B5SwbVUgYyg7ilcVxLFcynJbBORyp2UyhM6wrpyy8Ns5JSYZHHx7PtPj1Aoy0tYT
/wJNN03IekcyO81iq/d3+laXy0UmBMtOTUFRGcUUOYNWmvOYgfBeZKZb1TGk7VqZ
MzGTx1pI4a8sY/wunrBy+5S9UK07AruuhFontYuaO/iNDUazGIBzkBNwmDu8ZMtB
oyUGtLFnSx5DY+SnxpH6I6MIOKBOrHpKpS1VqmlXcwfsaU6k1y8DNNZ+ITu/Dfl4
NetXzmNKFJ/bHaSh/2g6rE0fQHQw7i74UkauiAXCKarj4yUZXCErbFGOlonzcFXs
Xj8A4znRO0eX6EyJI5FLK/GO7kL6a2nGCQL4xcN4NYn0irU3Z0AFWS4TDaTTEvDz
2D0YGL6gOIugSmQDNHmyG58FFt2MUwgiVnAqM6m5FQSpqpVVXf7ekMn7xudaBonj
jqhqaAdRqCD/dEP0oF6ORxjVeCjSOLix1o/PlTeKpEHiA+EB7QxRQhYDyxUDsSPa
bFN9LCADnaAnIbfJ1xMY0J3IbEr65lGHz6zb3pv/J2867ATWwm6mu+FJt8tu7rf2
Gq6t84FNHgrGKK9A14G2d8S27UQ0DNq9es0s8QcS0ONpdMcqWgIoGGmC5V/LYiBk
upXktXhFBZNma9u4cofBqfy5WHM396ty3EzHFC6YWT5oZFEcIvtoTXpW3jtWMK9n
XWTnOxwdm4kkP3vqrG5M/8rbN6vx+V0FIlojMM1O7yd1orCpHwhBX5Wsymauk9Pk
7KU4MCgIzJc8tlf0lM1qyI1+UteaSqCtm6R3ORuIwdoBx7v2BRmo17Esu3FKTsu5
eJWOaHhzPXAlvJoSFDBpe/mlGiUN0e2myYfCEYiC1x+7dp0yk+e2/Q6LTffckPZo
NHLuthTIxsmnR/ezgLcOxGp213Ifm36SogqDPmaB7iFR9Z7x5ZuhpuXIh5J4q2as
ZgSLCeQnqJFG+ZjsjKWYP1XpjrOXhN62iUDs1Bex7YLKRhSbpwbLinRq2klOysIH
WUDxwLxn1Fexdv7+q2qRQGw593KCa8OFIcOOZhCw5bRRx8lhdaDn58xrzF9aPGqf
d/tRYfa12KwiVQdlx78QJyv8cp6USFSlPaiqrljlXGjYKOtmnErYeNAytFk4q62x
FzT7970WBzZMpwwjmivjZMuU8e15XXxWtvTPBIA2rmGFDd1HiRWmu9qKlSqCdbDE
xAvq6d0rgWAzU0W5EyL2ltKqPcyq8Ijjz2wROuHzKWXkWLGpKjObgOojecTN5RO+
zOEDF4mPsb5J2RCgl911bDeFuy2JDgU1jr966PgngOUhWgVl76SZA9dKW6znWhCn
F94dA04RL0cHaGlJZwCbHA==
`pragma protect end_protected
