// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DsqKMqts0yh3aimfRg4XPgP4TCseigNNtQPEDZ0IWHHFJLRCUeBUhuOKxSeHoIdh
DZWfm1eNBiCgakU/Bf9B1+BiDYeLxx3xNtMdXaGO9Hlo2+xjjG6cW/CNax5GHu+9
LEOX9pDaDKeeWFcgV60mKgKo1IudKqBMFzEQgFd+f4A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21184)
ZDDbyxiNlC8N6LAm1fePzz/Fqf9j1nFni4M59f0yHnkNcQbJ5VXlRLUv9vlcFk3F
NBwd9u5qABWLMRY4I1jJmDk6xUJYRkro2OO4riQWSzqOuEKAi+W9FBdWe5A2ac7S
+/IO2i7C/j27rKxALMLlCfpxEF8Di3zMQlnn+VDMcLvXZQKF1yByAu3W9AL6ZkO5
TvsD1tkplJ8hHF5dtMyHYVtg5UBPwQIIkbTeTVXCdG6AF8YoCEQ7QSkcJlZNTx/u
3vNZKCp89/096I+aSLAJMK3MGGzr0V8JXjZyqkyLxRtmlXcwlmr8rP3WaCbBaugC
PkjvtzxnUtf66k+bIfcQtgC3NzUvods4O5IJ6ukoeUP8I9Ze+lcPhtHaYq6vlHY5
x4l0GOQtUUj0K+731/D2xdV7ZQAmlg8gROtdBusKLTXwu96UVQNB7xIG0puRfMh4
ktxg127euL/gsn1qbGpgDoWg5L6F/VmfuNe/uuEP7ETlGZwhQ5PVROQ8Q15sXvM8
fZPD+9n4g5KE0TyDMxSnTJpmFDRYZOZdswi3sryDTqY2XZr5ebAkdjtSqFWQulcB
+NwgoMammre0jHYY+xnunVZREfiMvfRxx2pHkzXqWFs9zNbQ+ViNjrxFsicVCylG
ruA5y0lrgs0W3y9GCGjRjxa5almmbjCDyGhyG3PerwFgjnKMgICnhcyMXI+OQ9h6
r72Z4BxgSJPYhERydGtq0JAQl22FbpkrMzJ1NgdBFVSlkmKLyANnNURligEcXeTw
n79Y1ST+QVy+Y3e7//MSRPOY/9O9r+RPEG7PexnblvCrx335oA2+BDeko7PyHAlW
gNnUZ0TJQYlhmyAlm6uSYaIBpplJm8J/qNqupB+PDXyrcXcr73XjFEtsizCJtG0m
UKXfRqrb9YNbMfK70rek+DxOlyoB4PVy0osBxORNU/RhfehQxORVme3nfKBkI5OF
pEIIuvWxxdGx7kjMHYfE+sGIU5K5snbps5y47vdIEy3YU5RakI76uT6T76wSlWme
/ciAZFDp+czO6xeGDVrsyReiPw81qJEwfvJgkUHW+mmzZ6zlNPXpWPJ+q4zFU4Jh
IYXC/4lr3wHh+tY7HYV8xn8Z98RVLU3Gi1nwBt1Gl8fn+WexWbEnNzwOgyTlWGJ8
rLx1yzWJIQizRUMBc+qXsaNeTcjfPhYECtVqwlbyroowlpDw+T87xEWDryQRMswk
kJJA6DHb+XHjFITw7TH2+zd5PERtAeH7LYBVkf4sFpYTIoHtseDFQGTBot9qEIY2
SQJJTsmLUvdhnVxBfFPyWUyL1QcGMqVBp5Diql58UScd1Umhe2ooeMHfCIn5r5Hf
cQA50sI6Zrhy7qWlAySRbi4U0orTXv6uCpvFAw0gLcRw2xSCyEd14fweCOx82gAd
evkpsVpE1SQE/26XWvwXBdk8pCQju5CHi3obME0c+Mc4uvApxLydd4Pz+//PK0qk
a4WEH8lXkG5qA0qeUKWcqFSDIIqTEGT1XcpH873hiH3KJQ9fWg1aAgP1hZJymrQT
wTcc+dYZoEf0QMqFlNjcqljdMPQRouBOX7PYiFuw2IFAHnWVFed9tm5I1nLVM8ll
jJiUEk6aDOwolSDku7FlbRO1LEOwyCczY8V0QgMsIlyG28jNGs3sdHLJd4WW1KZA
mLqNlpQv+gS74ddm37dxKcxLWzN6VoBHLgn6VAnnE99cWRM0mVEb7dLMLisqnWww
5VBijhKKXJX6qW07NESyns4K9ja+yU4gwrmHl3nutWL21Pk5400JDT9bxC0Iigfq
gaqA7IL1y+Az08raca9eGlsr7caOuuA2ZXSpPYvL/ByOsKunIhsMsci0NFqURyhf
KE+S9PYDd+uQNUX/PnkE+d6F0D0g0GhqxxIx5Vw94yO72MvOMqL/kSDLAlh9qsjg
tJO8AZVkxjY0YT0ZL/YmmjY77boU6XQy45nTxFDre3O1n6TiVj6K+trCsvVSZUsK
1Q0dSsBoWzvzDHO81Oy/+Wl4sLUbyEGsV+BwC9m+E6MjCvzhulrgq9VftDRCF1Ep
vQE7vtrILU3YrHeCsf8aUR74x42NqvYT/eP20fv0gbWmL4z11fGwXMO+gs/j3wvq
U4Z9TgwYqnnxKsy4o9f0CiELLwoYJE+VMZo9ML9PLIWnGI2hszn56ud5ilIh/VuE
lZEK3mUW7/I6HjDSgk2ehKrK9NUfWexGqcJb2Nhkz0SIBITCaQW8d7sc8qPxZw0X
z58MKEfA08C/Ket6OwuiXWcOghRJAdMRosR6xof1UwZv/f9T1uLZNXUBdSa/f2//
B3ypCPTEp70d6MmVHVkhM2vS21mTpNEI6Yo32tO8FCgWJm1ySpFK3Wn8w7UbE4kO
jO7H7gLsLSp0Ss8vxg835p2ezqZrYXvedj3Q95V0OIsnPeifultZ/1S9WWqiXNng
KcYYZmMVUvxjVNgYBQAGNDKhexi3tMALu/L9S6chL7VdfHIV6noaawLQI+e87m4T
iAionOd5BTwMbJWqLctGOIutUKBFrTZpEv3eb1rY9zi0EWU6aCRtxg4dzjryayZY
cgrHRbba5aiIvcKA5vhYRHBTrw+8HGKgEfuZUjl1L2TefxHmPcbtcQ5Z+2podUJ9
B2fXvDvGqy1g9uYvv2cawbVu9SDUGGwMBlM3trI3nGiJQVGJeJ8LVbTrwaP30NDM
WPYUooOr1BWWgz5QHG3NnrgKTudd5l1W3YenxcIjQ/6CkHkAm2R3HRSdsnkNChit
TyuXZFZ3wP7i5kBndzJW1Ey0sf53Zjeim8mt8gIF3d7AbePog+VdCllQqDGkLALP
9aIePepQTEW/DMg6kjib/DHnNL322Rqjsb3N+oAIpf3QdlnHspoRUoPdgQg3xSHi
LLeKfl1PN3QRYKfNVy8Rvbrs1VvuVRhz/WsNR/4UsvJWSQDyb5F0CSLJDIxXcFYh
UySBgBiqcgcu7XSb8ekYgBRxwucpJMJLuLcXXLzb36beLPpx2GGqw8BEf03KC8OC
ZNcISE7qSBsRkY9uftesOzQWce22AEgpYbmPWBzv7+ZUGG66na41wVXE/JylD7mO
XRxbIVq9TN9kuieEIo1vxk8Y6MQQjazllH7PSxRlBIhIFG4+g95dWDgZ3+UJyEXa
a1thw2/jJknThAW4f4hNXHivfpjgiGmGPw7ZlgaLC3oNJyru2KzmccCaCqhpSGbh
aecYkhurXgGZIjGLI9cX3U04L3XH4t1xI0zPioMEvrWxCtQxDZHTDzF/aIQMszgV
bv1PaGUHEF6ey7erGeXaLTG0cDY3k1odC0TsOR1ZFfWRfs7VyEba/5X3sWd2wgaQ
oLI8IZ63bhStFnl3bEmAclGlT+ScaSmSEJ3qfXHZlUYNLglj9B+arJgSPyr8h+EE
I0sC4Q2WY8R5N1xJyVKHOLMR8PH8go5l7ZTkT/Gxjf1DPkBpeb/sMNWa08tUXwvF
7MfON4d65Qen7uIvavw5bHKIpP9PWPZhES0VTfgQIGjiLuJ5yomFrd0446f4EBMQ
/0SmGWCcG2F9qLCKRBlLk3M7fPkQINoKUXrVFzCNEE+vDCSzU41OODly4NeS1erv
Hc3ISPsRBgQwMY0lkgABu5xU+kRM7Fe23wnUhJuq0dAfGVTKnwAeFDfiH/DG76FN
l1iZjKpKd6fhFK+x1xeGtfk1QylWdRV13BHT03WizX2WgUqnGKW0frCjJ+Q/TCSk
nuzj0lkSs18xzWjfsN3/wlxThB66cEgpKLnI3WY2BQ1hTc+8gmjBZYN4Gr+t77Dr
2mU6N41SqFi6nw0g1BDSzi7Ct3Tet6qW4ZFibLjDdSWyutmPX8U2gUGj+4Xa2rXH
L6NjD5w2OpayhK7fvk6qXpGqqI1glSDK6DAnFid/KkZhdgQ2TFgpgIYgYH3ce9Gy
0a8nNKx/utyTaJNMNoJmqckAARRp59ifvW87/Bi3L48SPLEVSPhvJpW1R0c2gvfg
34+PwZ3SnYgI4e5N4hhPgA/neV2PkOH8nM11H6VbtAyyeVVk7KgdTecAyvsNXENN
lc9lp4ZS6C6IWGjdYucHrPzc+fi0QGLUWM/opnqaW/+TX0IUYcWSY26jAXn3ywKP
dhV5fjXEx1QdzPS7w4YkIksjfl0n7rLC4heGzV2DDEBIkBdq+qzcLtwQPamGmez8
beuHRfK/6axG3DrgVwyD31Wsvm8tbmjB/abe/l2sCizdXQ7jj3nBVuGPp9g/Gjm/
cWIL2m7GCAdBf2xyVUpEY6CD67G78N7Ed2PXlEiL1u95/Gnro+eN66DBgaNwn20V
pEuBsgJ4qzPFMtdyFICDmHJJPxNWejAfNqrjGk3m1Y1HoCRVczcz5tQWRzMJHn9b
HHN0s7mNtQLM5TwA+j/hhix3y11VHD5CaV1TTQJ5e2WUoAKRJIVU/YzU9AKujX6E
ZDvIzm+UhvBm37DrE789xqhThur9d2lNRV35ZrC++VRx//8pFApsO+gl8MRVkCRh
XA5n2a6xJFsZxC854Djscf8OrUSrU+i/k0n2QnsV3teO5Ps6lM788KZNe2L54M+R
3HW3ilPiMwAcWwcP63VBaeTqwnHaUmy8pfjnp6moUwy3LH82jwXZ2IN+9x+Pp00f
6cCbq72I/xYSiBE1mTa4sQ0QcVE5ePtjgio7VtIZWVUtIAwLVxr0veQoN05sqz4a
zYjQ/swifxD+j4ZSpl1dPB5Gk6Xg4nIXNWdUvGM6fl6Rjn4A+9y7A7p/fQM3H2ll
9bPZvug8gm9Lpqz6tJBimJDrUlgYJ2jRD0DpHF81S3fY/AnGBqOYLYpeG8DmGv/j
5mC5VQgpA8HsYb6Za2eyyQdkaxJJuS5D1IG1tD/UnRXW+Zt/SkBqj934sbeNzH8k
PL847PeflPCvmTpIY1GBarlfigLon7dRahGO/vxq/dD5ucW6y665MMHu3IMYK0OA
MPivQfqNBCEJBkgh5lmGOgxNMzPkDqLek+HlggDfbzgCArDP8tKReNvdm6z1fPLp
EJP3vlreUrvEBw8iRWAbKNu1Q4Wid9x4MQQxYEqHvrdE5bAVnGWmpTDKIRf8Ib/6
P8VVe3Az7Pqv7EcfyjVWBm29aE8SYgmcDaFtwsZBbO3IIhiG+yYag7ulVENPxsah
kVGh1LCTc40TqGfpUtaPCPsBziLKiKGgzZCwhDdQXHUsSr8X8lYixHQaCSVDXAy3
DQpKhMrS6OXmE3R7H/Q6zqghnxHRILOBOP/HmBdnPKLfQhwnTGx1GMKQIapOtq4W
vfePjYSWYLOMYtOxoGypRiAd+Fhc4aZJfSIQMoB/eTTVBY0uBxO3sxdsEOJsGuPX
IGknCStC8svps8pJOIk5+BQYRvzZtQ6gfUnyTjDX0Cvz7cw5aYk+4+ULp/IvKzxR
v67axf2SgSDid45EDnuivEoI954Lp8gNHtKa2sqM/qkMFpw/ZiP+5PzeLcAxtEEn
DcaO935FbSOSSSAz8a1TLO+kKyWa23884Oin/5+W6fzWSjDHAXsj+rDsiERX5EQ3
JKhxxAyPZMpDpK8HSGgmaIQ9+MSkBlk66sgk/MvVAUKDy7U+MB4SVYlqhnpLHSTI
mlXTTGh/np2klaYuWoXqaywDQO0+mKbpuU1VJ69lQADB4vrxdTTZsLMYjRb5AFFd
AF7zvesdUvBnBDMapvTFNWC1oJy/7EuMnAgm0g4N0R0Fzv4RwEH072LyuN10bPGA
0HPZOX7J/Tn8wRz1rD/AZBY1fOytwOg0emHJXzMs99AbaLwKaNgx1I0uIgEj1QEq
dBQiCq3cdIgWs6T+yNUu78JQMpPju+6/9uOIadCN3WnJW8r7vOriTe/Ks2FzkwXS
LGwa2ZE5WnaPykhMi0/OECgNr5s7vNbkD14J2/l+axh19IVopbbAeL6tjiFVMz/b
nGepuI9O1XO24wXTEaLM7EsvboS7zreFGAazM6p4OA6OgxekgE1GtIubR/KVZTl9
ZMfGiRgPeM0bDHwcco4kKc94BXYCej5GwepBD8FbolKNoXw5lwn3DdiqdNiLRWLf
3lLw6zIgCEg35MDVRJ6V6hlkG0Sme/LK/3L9UtXo2m97kcD/AHLa3jqTfwia5TUe
U4abWYQ8MivAZpSmHLdeHP+HtYfh41qzFfFYBv2ixZHZGbErwH72tj9OvReH4eCp
C/JwzKxLeoFzE6ieDdk1iZZItGonijG5GES+MCIaeCERo6DRymytPKW7qTt2KtYT
CHBbIo1tuB6myDCy1WtJRaGn8TTXehNkbdzWkqq0Lkt/sdm1ULSsG51lH5HWCm0t
rTLyKInr6Zg9sYR8EnIAnNuvWgf2uix24Rgc6FkA6kXKg38tEJGX3O0jWG9YiGA5
LQLUHkKUxPGC+XL3uoMIE/3T0VowePtLSvd/euTR2wG+L6qPwe7ruqg56VUDHjlw
p1kM6Vf820UohD5ANcZoHjg6uznttMq9yNQnxzWMntwSXQ50zLS9zYSLeGjN+9rN
ews2Dc2fOjaoVBFLqZIj4NlWnUNHuUj9dUzp/3ChvsfmpUPHOzd6zbk4/U946ZQE
X00PFG7nh6uu/mET1D++TqD71mkiFcNwtjRyMPjuC836KxT9r+YuVydlaxBtlXSH
hCKoPe/27coNsNwctNdJMZLPMbQSeZZH9Yr55F4yh1DaHhf1sBmXePuS3sUMjSbc
rF9Ja0zV0q0TKvXRH/VJD3JvpSFEavOTY51qU5iwSxeIV9Q4e8s/7xDBCnKCwkys
GRDgISO9HaujnGaHOE1jhph03uOsetTZovrUe+Nt7fq3DYluAbMyyn57ZbkSNsLT
GYNDLgCOcegUeKEsc3hVuKi0utiOkPky44MW9NpNF+pPFss1HDyajgHljyKxvPS1
serq/edtWWs81b0mmEoas5XWHRb2jAMFJ6AF6aTJnCInaH7Nh+sivKnnLZehgkVg
JB0ve/vcX82L1flnm3gk/6dp95eUTVyXYUmwnq+hZvojYjyhUU7uY4elt79ZONWm
Un3obVzJ3AcGMWsZMkuVm18GUWJaJt2JTtCcJ3q/YbOShfVcd5Q1AH0PNaxLNBuJ
x+wr6q/qeK3ABRC5qrOOFLnk20Oju03nAwP9iOTScabWP/YZBDCg9lPM+pnoVLhE
UaZoPDtRaVQmzeTOYDGNG2TUGq2ElwYt+e1lVIdTzijN9EIyt4WV6V2OMXDSFOE2
QYaZU2I/Le2OJvIjyC9GBcLxeW6dcD9YGCNmU3xjOI2YxUiUNANdCnMmSW4ePmAo
HBgJ1GUUq0spulJPfkeT1TzCmg/zoRG3hbz2NzqTTVDyKarBMCmgZJPNpkHi0V5Z
F5zcO5nMgUzTdB8ynCHvfT5aIpOSPDOIg0FFwaFt2yup4uvG0LwKWGpKr4uG+l28
CyyKPqMfs8KGq9lHR96fy5AXPsyEiCbI+6FIfZdhN4uzHgpbh/+XMvDztj95FPFu
jvV0aHQOsWSrAR4q1d29ZGLOgslXzv9Erkb0CljQULujUnbc4wh3O+zOsBWQTBmY
dz/HCxU7W77Gbu5jSyhliH7xvdbhhc0IzaJ+dZk2ChNHfp4cg3Qc7Xq746FjhsLC
UNt9kVvZ1vsVjnp+DvQpsqVAQl3ITDOK25F7sDaFJ1u8masxW+lO2eCGc2ivSeqx
kVLWhxuYJXDwK0jPUMh5VKB0jVK+Kt9CJdksxkyff2AAJCESgpXk1WKnMhlaRY60
blo0EQatNq82qkzPR0FEqSWXB/J0er7mb+8LBfa7iTfnL9LKZ/CuKDbsJB17NjNa
HpR2LhFPvKlKAAMM+wmzTwcmVKOIPGVqgT2bnlmaUrwJSOTO23iHjF+sWZfYLlpv
0F8w0GcDqXmXtFL4Uy0wTGfhGHk7K8AE0TCc39zA77H/Jd3Ch8wI8eRCbdWq8mrW
GiuXNSDCjZfWrwoHqN9xQlyd1FNH2VMvFjVJ5eWakObbxFX/moaSwcMxQS3BTP6D
iKy+w6dwD/l+urOf1VsoBNHHyisctzlZoPFrhOZtzy3iExxVo2sEGm3C8ZJaKWSI
hR2SRFMyyFkBU14FwLXU4DEmAbIuzXBWtexWgSJnTKqpueUIlN0YJDu55PzB0DsF
C7c0SkbImaLWuKA7HESJU+J9rj5sG6mQG6CSmy9fYKVvUX/eu59GsZgVKwIzr+Ez
EYAaaGwfemgP2IrmJFYRLvP2+0t3V77B+ck+KIHUUswGp7AsQXoWwlEa2mmftFfV
oiQDzUbedxd975zpOuK+JlrzevQOrDXV6H+NHUopBVz5ThpjPRiyfwplGjuGYy6s
9fxlOHn3Z4ZQAlLJ2E/g8m1PGnMSDTdAVp7MzDDesDmMaOB/rTIPLeDln/igKpjy
Lr9q8Qi642fO1XvrPaYWhHaVAYcAV5mxOWMSke6Wg5jtquJw48BrYDAj7V1lns+x
21cZ83NoxQ5/94U9wRoYwDomH+ks2W9y/srCCq9sbDn8f7NtGDkABTfeSe4rWmGD
Q+2M3gqtXwO233shJ7fWFigKAoOE5HwiG43BhEkKoKHTBS4OxaxTInxsDmbTgYTv
qIPAGVhEVSHUa/RFVwc+EjUOONx5olx/oiqExzL4wpYtVnQCjmdDwdtne843w1Ii
j/UEIAvT1UW4jbTMwRCS789130TgLBDxpJvo7nTXZpXrxBx5mmCMCTTMnXKRv9Hu
SNztxKCKzCCsljlMKiFW3qUkAlglF1+0p9Ueq3Nr5vWqXwHlYSMnC4sk1aJaf6S0
/RYfJVuka3JAu+t2TCxBho36Mh5Tv24ngdWtPhTY9s2h6OCFt3jgjbjyloU32+NS
DUxWJFh1WDJz4i+ZYDnFmSaI54oj6ffDHspxyN53bpxT5C1SRKWpR+zK4ZOHiRss
X5UekaInLfBWXB/ATOqxKxMHq8grXtT+SLxg+vjOuyekllbcCmUujJghNF/PzFlf
x3X/mfWVHs/VnkyMNRIEbtKcJhGXzAbRTtLawsC8XVNX+kiyfK+f/zHGGjbz0upQ
nbkw/uYPizWFegOisBE4SBTQlXAm0+VYAaahHtYSQnCcTfOmFQKeL2EN9mWZ8agw
NwMjBjd1T3wveccsqIjKfelegZjso8Y0C6eaGBSwWVOY/69RwAq1zSGBj+1TAcq6
58JmF+SzlsEhF6p18Cyp/e5ZAIehrVSHgwEALWG3MW6Nbm7t7STnpX/gETWDULAD
5cw29haL/GhqEntUINB6yrrEbrB0r16VezEhf+NLJzVYtAa27oMYhPNbauw9Xywt
eFDXbBabfc//EqXvC1ynzgMTFqv5gl7Zoot+mjuhAU4uciufzRmSeM2OCH33C0zH
D2tiHZa1HvB6uG2cXtlUobikWa94WNjMl9c99y7s/K94sgWiJ4QvRV4UfOONddYx
avgOMO6A/6xJCXhoyDLmLWO8O4suq6jpRTX7S2gzbEup33FqMRvYgde08covUTfd
2tq/paLXd7BuHTAoyLIwKlwPidXgTuqYa0r3mNA4ddUi3gX5Y7kffibIgu+aWHjd
2YqnaVh27UueMoQFJbjoY/a556Y35WOJoaSJPBSPhcYHVbTKKXla9sicNRiicxkB
96V85LPFBxFsI+4BH0TvpQbr0pEoJQtIyOMjg9AzM24z8qPs9lfUXBuMoKslJKD0
z7AYxIwZVJbID/jj6g36wqRUpkC6gLm5MxmL2ycq0GhCGeqrEEJjbY0NMMiDZC46
TXICTOuiLR3P2o5T4C+Y3h/ATVH67cPRHwsz0y3ok5l/0rRyFrIURhaEuuMYvREo
lUpllyaR12gCpVv4PX3WWnOi/DewbQCiMq+AaS47kxin/aIhRdXnDoBvJWMYnZT/
vV2Kq6xlflRkYluaecA53XdZvlidCgIeDhcQalhcNUoWv/lVTthmyxaIx2CONtKD
eTtSWcDPkYKZrrLmthZF8byO1d2xTUhFaYNuAzT3284Ya1O8klCbjADlEX9adjq+
ci8yhD2D76c2YExgFUUcDZS1D3amoiN5cXRbkjm5db4GLf+J8HcGqiQUMebpDQWv
qq5hdb5Yc79j0db/Rjn33gc0HwFpXvDMXHjQryN8iApn9YaAX/8ykkbJDDIVDFZO
N0YKBcgECnCrjZ7T4qm5QYTAGq8N8aiSl1G1Rkq6pLwEPonGK5wj6ylsk2IOof78
4cw/ds0Be8DF765lMS2NatRepcqW8octUyJZWuSlkv8gF++dZo+R5QPv0P5PyFHO
C0sTfSqAqYDEi/8r6AOSZkUItYyAH5Kx5bSTMC7GZ3nmPeMUKdMkgINF2kkYKzBC
tflVmyUrdRTDC5irqgiUpfWSuMggbSVBz3zGnjZW4YSGZf0xpvsmgD4JLz/racbL
G6ZMlCpHQ0kn3VokLq03TghnL+qWB7Ntxyh5vwywRHBFyvBptveYVSuMYNv7ndhE
h1cDt8c6vE7OVQ9WRLuep/yptfNul2DeQ2MmPG7v1FnbdRYG5/1gAOxO85GQTlLA
pmmxfPpGNk+foBf41VaL9SBaNDO/6du8jnJPnQo/4odMjixEQmTvWIc7dp873QVF
3GstTgBAxsC1YSNBTepCnu0Ji+EU+o9FCJmz5li+ZYB3Q4K+K4PtzwdyJIlao18L
qXBegOYQAE4n30elJy+6whqvvRwvgGBRfm/JuEW+Ea8JwbUBUVFlY48DsFP0y9Dr
OXfFt8yTjrOmIK4Hl/zd2/ToaMJejyhtGAkH3eS9v/R9oduPHqYYarWjLQ6qYMEN
ChrDIY1vIX+yiof2rqf372HSHTvYrbcTaT60N8r0A3UAY0pNyKOFIh7NB2Mcogxl
YYrYRqU4SV2Wv39j/ZVaMNywZRC/+caPbTnkkSfnHsj6Z/B7HsW2mukku6WpMqnF
EGEVodZrSQmnk4zlMntE37JhIxypM/AogrRQJpcKMj8FCnM8QfCvlY5zGMWRCZn/
DG28HOrZl1SwP2I/faI4ZKkp3AY9ORf3LvZAd3ZHnU/6gd9YdGFbglhq23RirEj/
QuhZbU5uGkKQ3Q4JfhJXI210pZg+0h/zWnwhShZRhQZwHx+ZrmZzmjbeGvMduw48
jd8v3CoW9hk6+/bVoFtSpuQqWu3gn703AUlffc1nmYfuow4VQsudANqOUBGYOrNM
n5CN4mKIuq8jDrnP5KQNDaAb07qZCXgXb1Pd2HwsL0Maz1Ai5dUXdMPHoeRP6ZF4
Ext/W0a50uCh38jfH6rgDs6FRNwNhAQoeQMT6iYAnxeUAN72TD44aMXyMaHzpb07
jaYEzL1HhV9B7m/OVHGMszKBgyoWR64Tp5pLeHzgB3VQX3Dh7wHXMIMYqALvXcd6
EcIvS37iJ5oGDAJLgHIm2LrSFlV2jHLIdE6Q+L2ZjQVf7bGeKFBfJQ5G7dnM330W
KRV5GE0nit3kHjnWLSdK6db2WYo5yVqKVGe9BSlG+Oc+V4DN4lN5A45rwfFbDTAN
0ObTn+NoTtWPEp0gC13CqklA/s9OWQ2dRVqfmJcVbtDAAAMazIFgJmhPFnI1IjF/
Ka3l/FfyoVBJdvgBJ1ONOrYRk5ZIe32kxYbte6FNb9e83IZSGCrp6BHiphJca0nA
VvG+iK0LJ/Ke5SdY3Oos9I96xzWxk25tQ8PpFUglu65aLJ6rqZOXpR0w46/WA2iC
QSbSmy7C1m8h+2qglq7j83DLNlWvQFQf1lmDhBM5GxxgzBhFxRRV+Vl4hy/HA6xg
nxPYH4+buYFaiSt+2iYtoSn/q/d1Q/UqG3RxCd80V1UkI3ZS7yVFN/7HAAj5ZaBp
FYKKhRDOSd3tZE/Pm82DuihWryMx714d6qguMmCM4bIPmnvFDdp8WRa8us8cAT/k
sWgrrQn2BM/gxB6sHIcUUjg00rP5Csm65ta6wcLHv3PplUNAaJrnfZQsPTnmqpfM
w/AAe6OLrXRtH+bmZ20e6r1018aWZmcmZSXD2GCYvoNTbVV4yCEG4G6eolbGoHwn
T4/JhMSjqRTNCtB1XgUyRCvrzhEVlI7DAbVkl2pswZN3JNsrYQtK14qTIpbbTJ/Y
4pa+kAYUvq9gplL4shTt9IB4vyMECLSC0m3nTtNWP9+rOk75QFlMSrQJsH+U+lTb
MqtvFKi7WIe+7/xrIlZj7eWLw/CZ28L0/UU0GgsSrgNr4bg0rknJ0DpKeqSLAo7I
ggTzez682/Sxu7ktzQIdO2l4BVQrxKBkjknD2ktixoHw6hNktRs8hfMauJ93vYzF
ZGKNDHwch1osN6cvCAf8fKOBWBOxNKUrOHJAl8Lnzin+bOAOVJvIsOlyuy7Sph41
PVgY60WprmdCVsmIlHvcMymM8/hKIdpOObytFjA560ot1hTS3JomQzq4SjN+wOYb
lykG7yFiw0aKTbd83Kmm51yoBnqo/CRSBZ21yqhDEtfYcEW+RKN1TY7E7FQIDV7t
txUl+HOiafYlR+wqgsIM+Hr7ow0i4Sl6ottYgim/9Hljq05oJX/1R9ZushvclZJ2
ZILaOP1HFsglcCGV+ZXKvkNfEimjeNHzRgwevafkigEHdf9EvcafXf8Q2VYQNwGm
dm/aQhPQraSN/OSTmsaj1hAO984iK0YZGdkNbqrol6n8c4gBZnwa0wmQzBwAgnfn
PP2AxLJsyVeaixcvZ9izWpQEJg/jBQdstAnePsJQPvQJp+Ho5eZiv+iSjltZZqmu
vduv3X7roG8c5hXjx5OTHTu3iF5AhF71iGBfbq7xQgEkQWvUovg3rC2wTN05qySD
hUOcbqnxq842GzGQD4q/MKbrMOP3NHpNRq5YbeJSS1D+sQ7n23zHcD9s7+N7P8wy
zRLGDa69Oa4LfUKcrZPkG4qoajutX77XVprFKZyXzpzqGvXsi6ADMT4zmaBA0Mbx
KXpgQgKU5LRhTif8vs/FHtqAkmeaYxTY06c9jMPEK4k83K6d5mcsKcvI6Mzu9Iix
ec5HG24oYTsyacP4n8rgJEOgCs4BAxqNaQAcXmgpTUNuwDuWv7lo4Jv0zcpCfUjc
kmS4FxgWcRb6nDx7bhZQkzzBmaEh+iRkWDSR4jZ2bXW8+wQ9zgPGaOTDOAAiHpT3
7D4m1i/2uEPvJOTVE0QdoZD7kGSTaBtZ9MhBuCxLEsNUYvkF3xvZXX/DSG1vC3xY
Vram3KVYp6LeDEHMGqGmS02yLRB5iONXcxn/Eay6STJokq7kbIhiQ5OioN/wWGCK
f4ARJgfZemO0t8qFcuETPrInCUC/fxHW7ChjI4DdFsJrFt/T0vwiuCYhODQKFut+
TJ2gV0sGDQZSXA7NZ1MZZOM7bzD2lKbOfVhpzc6FiGcGr9ghpORvkU7OkERtAAqx
QFAzZpqLbbCJyd8YSM8mBECsbm632JWhbNM7SJ24qh/3RmhW1FRBmslXzj2kpBPX
gnjQyl5ffsr42IDfv9PpC/phHH6cbX61CrUJ1Hb6g31OpJJALsXmx/YjHfnODayG
y8w13Kh+oz9+/fR8xxISN6e9batlSDaLkYhbKf1wtEwUMRgas5+EKxVIRkawsbwj
JtgkqAvBsMnRv6+79DMYi2VO6kxSz9PN9K1KUSbv+uBXF9AhoMYE7VnfXR393mdT
9ZR4wsslbSGbOugR5TgSPnLzD5RfRP9AX/u1czTkZ4A36AaCHhm0Pf8gS28roVb5
nlUa8PDKHQL0rLqGuiGjXx94twVcHbJcbiOWQ6bN6nUN3SJyMXO+OD4Q3vmtCcNJ
NSCbBsuh/hOx3H4Xkeus2ynou2I4ePUcocCA5+AlkkvwwtehnKVtSEUCf3HENqD8
p/iEh/IGJbh1dNe7OtGMEWzIjq8xOEurMxtsTgz3JjsQfwcXR83+MPRjjcMU0UlZ
7dc+wtEvA3f8KVZtbUA1jG8AlIKHjwaaQnjfSh3XGWJWAeaJdnPwSTBS0RuQs/EB
0tCjPHVvFllZjjxLyX7MsEsjZjL+X4Af7vMr2iHaGLJhyy1PIQjidx/voCo9D6LK
9GNUrxpDBg2xsbx7eVXJFMkENo/Y8EPUaUdK2UTlXiK7CLj4ROWdIYefWCgN3TAl
mTLVdLiZ0RmaUk4kRYr8PWo7yzi+jUmrGQzOivSSQdQ4Ahu59rd0YuF4BrAlzx5Y
yWeHKirxiO7GP9G8sU5fed9wZw55Dt+TBxLqqaVmI490LajcEoQUi/8g7+RSN9wc
uWy6czuNvlC9N3rtr5/HRpz7d3fHXtK7WT55WMAFN2XIjPwW/vCKY+35HkG35k8s
szCF33KOdZsC/MJia10gC4xFW/joYLIH0O7440/vwVVqrrLLTSCTov4+ovdyVgZs
80FNfTRAk0x9QoJEcoK2s338QIf5kOzX6KpoqQNoCmeMqan7l9BNXbUrZBVyjSPE
zpjvYJfz3HassVT4EyYXfhKWW9sME48/oa11LKE3Lcs7W2LRRYIix1esF5I96d4J
uqX67QKQnm6f1LsrVrk76+R8n0HzqWUbeneerKCYXssfGGbyALzXzFst1v2RzeOh
EFp5tgz84TLeilImXlSYAnpXPoLFMUdtn910NEF8ebI9Ov6hoJvJuiE9H995uT1T
SYNDf5BeIyNq/qXg1Od7pOHMjmXxNlGkBtFXxT5Eiihhl6aGzplSI5OtCnt1jkVc
Sp0vIE/U6XrCE+CDeIDjxYbkwTVdFw5kyF8phljGiiyv6PTtyfoltDM/EoXvRse3
2Q9lgLsDit5bfGoTMuo/jNAnJ9GgHZwpDOFxm12jRFrTvg982JkrNix+9PkeDKq9
hjYaDV9QN75dyyG4ZKWmHrknagyC0ZFP8jdkAYtvfO1y/DuMsbKnFYJc1z9f4PBG
eccII/2IaLZMF9/ibLuXI+CaiF3TYYYNZkfoCdx325H30Lti1UvsxPkvGSHh6hsA
414J0fO25cfaPzypWKiOHVs7ISzW8zcivmjL9sXk+uDtYZ9IBAPhgXwsVxLARlaP
9wJN7QNf0AKrBWY8pr5+yeY8y/ms/MWc7o9BxiBpqaDq1yqcvRid4rVQMNrSTQyo
wWUMsGPUBXTIsszmFwXv9FZaCx6llbSUUvlUkGCxHgV/CNDcHT71ecz6LRzqBmYt
vfi9CMxBIL3pb3l3iSD1cz0XYhdpyZGUOM6ivJ+3y3P2U+/kk43sHlfTnzX+i28f
GcENLqZC6nBbdBl7/3DJIU7LxdKzuvXel2FtQ88LuCXyxOWxe7BiPwd4cNmfuwQM
SR91AfOvNCyIOenayOe/574VWD6sbxGaP3ntjR+EKr+iJePPkHwdqAGmLrFSa9R8
RLKcGHSRkTwxYnexC336ZRtydqVHrphNXJBdo7qGggLH/NayVgV9IIj6V39JQj+p
XTopJ6YCOMC/YVewu8gSmKAcTTxWahUDXZerQW9TKYps1T5rg02ZMxJ7rqYcjUmR
x5Yb5lnAYFNHMgH6dnpsTjjzFo6xFEjK2BCXPycqVAs25HHlia0vPJiU/MRPpqTS
H3LRn0rh7xZoSFtJV103An7nrbgqtmOfU5bOAaWUzmilffrgTjakmtZDEnXnzGjU
elZrqrITwX1osp9HFLubQToHs20F8vKY8Ga+zgcOPWmbXPF9yFMppLvYGPJXEf5x
XQzOTS1LRNYyHqbfRr9OnriYfEBfMBUX2sJWhVYWaM+t8J544T8m2mXRj+BtF8ZL
s5+7hK2mPtMBJ7eohbr8DITAgfYm0HUtsfFbeIy++Nkp9/ZfD7H+rueEQ0PRaiak
Pf//qv6YN6+knxcYnwy7PDeCRCzPZFEUNiZw04LvuejRefD5Uovko4x2gJ/WROIt
Hjv7fDtFiQ1NKzK0zShUMNRaF+zjtp2nP58Iu9H7rUTWD/Gkol1VIK0G1v+xL9/l
kDHBZVoVOO704FXMATCdp6V8wIQs2k9BzvGxCfMfF2z3IduZ3lukhaE2eV+vA4j8
nxRerLiuO3vK7Y6qXowcKloo1XcY3gxayNfajqHuSSg1qxi/CSaQHFMbU2XHpuX1
GU0BprSwpGBW9sHlgcEAxf7oGXFB9jlMEjih3uKN8a26tbAik5s9JJ/TAVjRBC7w
wYdnBfQ8JyJJQepZp27jOAVmGiLDxppBokrOA4AKmiSQ8ZLrmX5biuUrvftQ21LF
hZzWu0WXCMy2aJT8e9/hAzjNhml4b0txkHRtqU2VRH4AUTH+hxg0cB3humtQwAab
KIAwVA86THWktp3N/OKCSPBYGAa7R2yo0xdWhyw+k9GRDVb8LQzLybvCTzrGAz3H
W2Z//hg8hr//i9O9z1dQ9kTEHYcxXwDqAv1tnemU9GdbYqH5ksM0UoHaGgVdX/I9
Fp0APV2EpXC3JEaJDYcMrXENrnwOY3qdhKPuxqMIN07ezwOv0oFMa9pBZo85Rs4b
oIY4D3cGlltehyH9WqBICYAf84be3Auun/dyXKg37srvD6IJ1FXofY00a7LcdCdd
N4MSf1zyVwD1SMsKI9SZjjFJa8rBr6xhWHNhCnP5rkjfGRAAd1TmuVSbDqFK5Cmh
qdSlkCrVNqmlb/Z4OuL1aZrgzeql6kKlrOTwueu7lmALBuGcYutR3ZOhDKbOqxgl
U8+wpZLDa7c72sMsZKXdd/CD0b7dNMeLv7UUa3GX3mqknzrRGfyClI27Eb/zlL1E
W6+C/DIiaj/+hJi8j93huY3XYSR05syKn5iJgiDHb+GVeORBInXD/tA7lLpQu+JD
4NGgh8Ur8kxxQkvwkeX5MLYvBsbxpOYTsiSgd1edNEBaeVRlwj/tSizAkSJcwGUx
zu6Tsu8trAfN+1NA97tJGERES9Tr1sjQ0sXYUjMRwEC0Z7OdtObWDOWzyTN948cB
XLtBqS78NloMkweBZooB4VNeE+rWcbgkhX8iwMTjWGuJSkFLAD6IA7NE1sChLsXq
fR2KqrIlK7T+F2zOtuk7gaP/RjpMbF5h4CHI+PatqFW/Hb/GzeDsbpTghHAaVn+S
iqY/J92/uMo71Ha8oajJ3H6brGna3UM1ykcEWwGFOIhM2W/YSo2SH74J3MWXHZRW
QS63OaGSVIN7JvfvAlsB1iQq9PYW1kcDiy/3sAlF7giz98KOQeTrN1wZ4/+RNHFe
U5eDSyHgFIGANJh+/HU/9kosi6bdY/xW7JNWwRqTuJyo0zXOaMk816nLg7+WTbQA
SAPfMmjPYhh4EvZ9M22h10sAbqGCvrFOzyi7JvpeoF8LTbZJ10U1/Vp2UVN4+c2b
0mbp4UZaCoeZPPnUf7Zot/5aSRQXgqgGW5zrXUVWjZEuwbWexPFOEkbbVDI2k0nh
VTmSTW4uWOkNzLb80lFRx8azL91fBaECGYO22EOdMVHnxY/udaypTD0e4q9EGBo4
iePPWAlkkKfWG09uFt+y7M7ULsLQme3BPqb+1xKzkNSyu4zRBsnHN7yaJ48MqHfl
wodfXwwH3MyStMI0pOE84yp7Wp9zctCkBhSQHHPWRiPx4FuxvQ6xCj7YO+4HmU/e
zFtMNFrZZH5VKRRJEEXBElOc+BJgvH8+ouae7I4E/67M0+6gaJ3dDYaiQRq58FJe
1yuyEZvVo/gGDIzYUN8WBnhg90yD6CP4/LKjt4PliiqIjj6kE5x/e1YSXTYI64Id
01qdOFVJWqF44RS6fD2wLpm69KBHA/P7ZYZbkcBXX/AOZf6UwPTsSX+oeJf81+r1
syGFcu5izq5YV7XNTRUZ5Hsx8YKD/zHB2HcoSKCbnc0o7vT/hmZ1OBjgWtjf82xW
80y9oF8EE1PnsfwrzajhPTHtoWVP0NnWApFCan19fsukkvztFhV3gXPoGh8HJAQa
arZpWfx256WJil1IrO29HQUvcEr1vuvJoWPzIJzYoDpfVhd3a+wBN1whzkx1G/QA
pczC8mRkIzUoExvA4iw6S7OSHff1MS5Gg5G8le/hqlkXBxXyIOzFgfCMnnblTIAd
ig9n9IEn/R9+ja4yLoLBeHhMyHZ6nRAM8UeXr0AZ/dlXEmgEUqsz3M4IOs/PW5+P
GfZqQiL7rp3O9z8BH9d1H+dLCgfbLRyqvoj9rAKAoKlmMJkKAKMIKg7hH8wgRb5o
hiFsZhAGK7peY/KgZ9sf1O0lS+wjNPvCwnPfaLjnEngh4+Qa7f/hxMaTq9WEy+kQ
5q5PVBlDmk4EDWvlLifk3+lwAONKmI+DpRR72KxO35NOAW/EbIBQJ9YUQC1HtkUo
PTOu3k7hQfyIjrkdicXpui3Wwfgbm+VyyiAtTYNsmHPliq8qlQ4rZKfiVQpLN81a
UjdBP3L0MfVOdbe7Sy7e22Fv3nD0ONWx0bZrkAOoV1zpd6SQ7kAc1eHGJYazw8Z7
p5DSgwlQSqkDRJ3kfFGLGxyHO7TIT1cEddphqbgX1znIo9l0SU5HQwZTS84RmZ0A
ym9/nSTeH0ZkuPhgeOCOYpK2ftmd16soYxHo5KEWZbgMDvWAT6PNNH4I+OlLeocs
mJbnVZDTnq0gFN7Y/96FFpkdF/6R6t/Lh/XhzG1BN+Vg+hWonn0XU9iVJ2GjghXm
OhN9j4KDWcPdwhXefktpvhdghVFFXfeZR+5+iwQDNRJBOTKj1vE5cq8deJ7Q70Ic
hw7FJuVZmMjfPgfhRDh9BSJSppD3tJ4FS81wq9afqAIcRslJWb8LBNnHIRmB0Fou
QivZJRpTjmr3q0WDm7fmibyGjnrouP6FpLZ5JribOhzr9mBi/eAWKamoyPrEOYR2
mIkr0Z5DWceyOOzDpNSOS00KpUPApIw0bHsww6gRTaQSF0hOgDWGilpKFB2/hmD3
AMh8UEcPhS76uHmyjkBDIRjjPS5AJ8AiQ/+qPe+FaM0Sisv9hfeKIbesGozL5Czv
Ebz5mz/CVcFJbSIAlS07EALbd4T7mUyaLpS6CmtYxg47L0GfWxxm4lLHrmq4/hf2
Sqt5pFGl9sSaYCKgDh3CjSiKOt4ZU6B6TJceVZIJFPCWL3i1BXMjzMTlPhJ8+pfN
EKAbKbLVVw5z7t1iife2h1hNcCAaYvKfodJ4JEwByjQMBQ8ZqcpZ68/GUKo4EtMC
32Jb8xiZ8+tRwUO2HOiIXoF6K2jHmhh4v/AAIzQ+pWNc8A/fduytqWsYyU3ZK31h
I+aSq/JoOPCSFj5uprN8fl+7rN8d5a26IISOuJV2lGkuQPtefOpiQ7eVT78oCoYx
Ap1NJNH6NLffYJF3hdiw1Q/oYOgQy+pXuPlQ96J9n8XFaGIxE2zSniAP6cqaTIB9
mi6QB0dBt7hkkzjEA4nQfTtgDwuPiRqELhFnc34d9tpEWkjhXQM/mcUvfDT1gHDD
YhNfBR4Kzf9F03hVOJtFofr/G99ms/mV3mGaQH2jtqsmpalDpCskt6Lr7nYr/75b
ApKlGC3UUxjLOy9wASq7sRHi8T945REu9Ez0IDeFtjQZMr1WGFJMZVf8eQPc1eBq
fHwDgcJg3iqZRsvcAZq/4S7AWfgo2n62mxs0Dg1qhEbUFS8okoFiPZwWqlYL46Jc
SDc9CAAqInGNP68+C2dkyb6PCJr6wdtig3ZWsN/stXxclgLG9scyFWaooPjirp0O
L/aA2+UfnJxBNHr5l3ZOiqtkxV8uMEvQk4NS86KjSe3jZf2i0MUvQF4afbJ/GtFL
Nxk+6Dp0thL0b0hIHEPnk6zO/QMhpUhlKUze+I7tv0geqoCJcJPnI6avc3zHt5rc
6+FVPL++64fxiyg0Q4wP7mQzzuiu7UTAMZFcvIwoNkYJxogJ8CzD39OWkVEp5PUQ
1tlFaic2BdqmnV4x7eavd1TVM6yZQPRpZQkIcXYEFPcXM/hlD2oHdu2lZ1HLGaG/
kam/JPjLTZJpjD+xFEAB0JEGhDn3NfeB5RwKMVZ+KOW6SA4UrZE1GrTTr/7O9wM1
s/55Gblq+nYw1J8cxd6lUMzd3iI7XyTCxNVbAgiGrjAzd8Hz5mikzKBPLyP4aoaY
JlcQsmN4BaVnhm7JY/jnR9A3mZ36NAI9YqcGxUvlzIJpBOmT+v/Fcx/XqQ1HlAgP
JyW+ZILQMxSzZP1ee/uZSbw3TLzdu3yjBh9yNnFhep6tA2x32vHap0WBzC7yIxig
knawNZZO0WAS9jLFfTzc2EyvbSBXPz2gJAkymLkHlrvbrnbI5zJdB1I8/Ji6g6ik
ddo962uJ782U+LKwXLekimgT7WlSg+SOmmoXaXSjW+aOuKjUeXA+rKxSW9xShuzD
zkjeaVZbTqWbZeEcVn5hxLManGrCDIHyfWVwSjyVD07PQ9smbvziflbVHK0srpcE
Brd9P8MAX/QVNwjOXdIFlj5BppVP+EWx5DwxEo1xUkuh2R9Ti5jpzQvJ+dE6Fehj
fehYzKOTgMipp1RJuGA9CEX6NVcsPL/fGIU5vMAOshyM+gUlfHJ1DONJSt/FVC1a
TeEjoSDNjp2xvdJqSzWEoXsWznzJpCsg6Zl7V8M3yB9ZQHnjFHNtgURCqMKMe36O
4GiaYMoQ/y88+a8c5iit6schyOmUauNTecFjcAQbsB2SyPx9lPV9UPSNs05/T4io
zG21fpZKe7bKUY99x1PXKa3k1rjf1QLSS9EGI/3DOeBhpZKC02NRvsKMcRE2jfeA
fYO96ptehnvdef99EbxH9C70I0hrIaVonwm6Kr4XDuChd3x82ByWu7FUAScksaN8
cCHrq1f3iGqyEvHH3dfpFl8jzMiIlN1dMq+CHRNdUOfpQ14SsNC5PYuf9yMQzqPg
JSedo0BW1iOQs6eFmVip67gGDbcJKrOvFXGO34VDHoo6OsdD1dpnPuYKJv/ZruA6
C4ROZbuO46dTiK7GehNlyjHy+djcPmC10aU+IdMXRWwW5bRXUZ51gTXRUVs5PvvH
xROrjWg1jnuYcSdXea8tbbDfBnuHHVWsOas3o0naY6NUwV4tBY62NgQMVLv0ji/9
16k8006HArMJdpLL5x3Y1OhAn6ky+zGvxmtT65dwQbz0QYcxTHLhznx9e+R7oPfx
bDwP6AUJ7dWDgZlAXOhEMSMs22GB58fM0JQVL+zpN2f4Bx9/5k7CLDnIzhs/korP
pgmW3etQWX1ETkli7dw8CiBfS1pvLV9xKVejhkHswTz5pqypX7qqVXj1vFnWgWIi
FCmyj4OAUlPMuDD/Uybnxiu1zFyX2W3itLdnkARg7y7h39QkxQNd8Zq2mH92jfiG
Gg+wsgHTAvupTs5X2y/kLFx3QprFgXn9G2IDcx+MFQSJB+o30rAkiaolzBIOv4TU
yzOWIuO5m+lyTFm1F9tTK+rQtAk2GlhUidhXYBSWn1gZ+h35dZkZXQhwusDqL66r
i0CZqNmfPNOoK95NhhZOAJk98tfhfXITrN22coqUSFACIey6bdRktjJ0i4d49QLP
bHeYQR2QIIsdfqg90/Mmft1I4RxXwHbCHMdI50iTpx99ugjmFix82b8h/kB3MsDP
fS/rXRKEaiOuMIJfkiRurHtkbG4o8FEBn89XkaO+jn3RycfeoDpo8XraBWzewLJf
ozqzIIGXMmEmLGORxQtOPU1PNUAfGPYkeZY7Yf1MyyniwMsT8Zz5UwYC/8AJaQUG
mrnnTiideiIJ1a5YKX5hQM/XDa8MEEcPQ79UMshSObYfiwI1FF6SFm3zqH3j4626
5aAxBZ4N3r73Z7jbG6o+AYJiXY8j73jLWyQ7+nApCzy2yL0JkU2F1YYHJmjtNHgl
mvZOO9Bw6BLPqtx2ywiGPqDAhK9tz64eylQLO+/x2xxtGtePWN6t/PUJfKr1qyvx
zMvmFXRkVReQfNvEUjFFbLC6dGYhYL9JhpgnYlDunixm0YloIFV7kgRsmOZZKEC/
oLKx7ysmBVauATfhDuQzQxAEcXm5m9dK1r+8wlXea6ri/7256wFXul+HA0p/TPiL
rgwcEqwSvqSn5kVZ2LHbdU6RGVe4oJiaMSUqOSiMXuYffqb78C0IUu3nqE/wPtCj
8PGUmeomLGhM3Jx3CQJIHF2tWjIHGbwTACmpuNl4xdF3wt0uj1l8jbwHerEXKZA4
cyCAXjTDLkTcISQR1oFe3Gz2Mh9g6SBtHhbDIX50HhymUaEP5pAW3J+4fQG4bbXb
14KeyrO8ODgbj8DUWOAj6szSbKlysGHTwbC1tJC4HEAC2WO0CTePWPSMSg8AFKJQ
lQA68Ns+M0yDlNrApZy8xfJAJwtRcStf1LoaLWb892kXH3kV/73rlPL8PE3XQBpT
oPFWXnxioLjipBa8JGUS5UR4TAnofVzQ2CdL27RfFqzOjGiwI256Ue9V/fje3bn7
RdMXQV6HpimRZ3V000c76z03XBKlRjJ3quN/e4UhhPLTGeoaoLZpqJVnoWpQSK+8
+oxN1aSefDMmN9uQGyw2Ct6TnaG3u1DBPbmgwwx8aL6iTIWYvofDVwhqTlI30rxT
E5YZYocHEUZhhqrp8hU//lG9s/7/ZlCnRJDS/tEX7O2upHEjSMFXiOXQ43MTjPow
PQRxnK8tVT7S+qzlTmeJBdU4AjE/Y7E0O6rwPdNY1TQO2k+iI4VdTvYKWi+yJ6i0
EuudXaw6Epkw1bvgaUfAf2+atHOZOPBSsx+VMbVdsC7yBtl4neFwO4h4Y0DmgKLd
GI8egPHtgp/LUTvHykWomaIZJzwMOXcKt8zVGgF047MS+nu5LncFb1OPV0FmJH2J
Ync+xq+eicXBX+rpblGe3cuWnGnU8isqwHfXbjS/GZoS1/zFK6+zRonyShX2+bj4
WoVV+ftt2w96xEtczY6Ul/JskRI3s3/hRjslsoOW/XxnIE9rW9qeJzYqfqF50PJs
gjAxlvYvqQBfLz2bgzB0zGjsKh5CSuXCeUnqO3p3O+atMSeRLEOBAT00nd4E8++d
GzuSvq2+MztiuAqaqBe7OB0vMgyAL0rI1MdyRrZaYprbPMy0WlQzHUuVFo5YbtGI
l8aTpMZGpHastQgHkjt3v2CfeJMON+SdkOZRImTwPysNiENw3MG0c3zy1rmbeK8N
BiznVEqw7sDzBxgKS/CR5+Ym2vf08aknyOEbe3zarxfTlVQdUse8raWpYp3JU/cd
mgnTW9jnvlrHnSa43qbV3OLuKivoYOgVmoWRGvdZAJzsrnqNVe2eriRiqdXCUZBM
IQpwM5cl/A8rrdxPQcYGUKIYGLZGkhz17rtOgXijjOeegc+GLlpo3YgwCcxRPkz+
YgiKJTve1mruDfYnY5y72tcfub5vGV4IB8YIpB3VFoSticFLVY/bmWefs2DH77j/
rn+ynrmtnHyWbt3j4DdkV1CL3/5Xnd2HpGAcOKSqSAi8h36JqWiyuDp/y5gT5Pkw
0XWBYArlQM6A5V3r+l4okAOynuirzRcL/y8FoicdSK4rl9Yy5+AzZPC3xXOEtMs9
WsUAW54/t4S35nyes5APo3S69NiDROVIECwOKWy46OEq4PcCQwcp/Ev3O1StKzDV
BdeIPlsBXbDqCMMCRjSlUkvPOr4f6Eru5dW6juhyuQsKcr/zq9EqT/M0qMH0mLUy
zuddGLjhTSncAeLBit8vnq3f6tdoQnBvML5giHrZ8ZRS7Lg8r3/PSEGZAHTATotc
9AbHYhF4191AvukkbQ8A82a1kA9EMOeG4eU6CcnYHWqpyeMAg+NssOuehByOuLXA
TvGWt7W8EEPizBdX7ebYvG9+TJ4Pst70+M1t3KjjfHJIZAjNGS87ct0DSY4VnPV3
xWGj7BZAo5SFTctqc0KdZRX0oplqKCf6hsMcQMMhmmDAN8z2l/NXwHMbyro++cuQ
eSd2mAjOHie+RcshBd2/XsQx8bQToMcgq1K4McJGy67q+zXL1WvuXDT3uOPRLgh6
7Oo0Kfu6C+1bmzzZwW40xQGhYOfXr10zQfEJ8wkyud49pvMywlF1w59HBbp3yu6z
k8ceFWKFqMaVP3b166Xv+K+xZJM9LBWZizi3W4vP7DBwX9AZwCF8+KzA5EJ9Ibdn
ZNx5lvpn+fD6MEnTpjOMIcobtEZIGYwajNp82PEiDTXIOHU9od0JKTN7CXQ42B+1
3d5GWM9ej905QgJrdws/VQz44dCsLBK5fI7d4YXKRZUoh3p7qW7Fp3X/6ipidBvC
BAR9aOrINYBnu6RWlI9M0SBiio8sMPPTCVsRaopFxQtcxRiUe4sCX6bOXGlFdA4n
HuxjCUSuNxEoIVpI0D8eZeVyYIswt8wjx1ZfOzDABPRTrQh5e+/NTGz7PlGB+uOv
cr9pEdfOze6WtYC0Je/d/PggIzvb66M9PN+CzxrNU71hEzoCdWHv9qodv9Vv3lF3
7X2BXVmILeBpm+F0+1WUr5tZea7VUFcBA5WfWS1YEARkcRuPIjzE+IngYhq5yDeE
2a4JE9yvGDARSkkZAiRpQwJP/j9ytBSp0bco73LdIQw7lDBMGAqRO5GG0v24qeDf
NY3bjQMwzmjpLAJsdPQqe2UxUtFOatSdwCQZUzCLbfMx7fA7cZZwnXk0dOtDu/qh
PegGEblvs8GboZAS4gcRCNIXQqiGtdtyeO43vVhq52+D91lT6L3zgc//7BfCiF+G
JQMnf+iLHsduu/822VfdjniJ5uwCdgR5HCiq1egC8UIeltd+VvR1ACieiQQ2fkH+
Dl2f8A+e2ZOQxPcp9MTbHT84Zziv35tbH3RUVzciUvMLqt3dzPVuMru6Lu8+ZnvQ
Dk1pkz0eUzLqQUo2orLZU860mMYGswi3LXdLC2MKdYTq56KHq9gZUJcKgXZfjoQE
rKmGiMiCpd24IL9TrF/QSvidtPbjACOBPRRHDgq7e5+Royl9YTyPpwm5ZQSyMVgt
YamOOnPGo/4xlptcOiQOTonQKsVLQjTajx6TrSqhNJ32r+HzYAyR8PtBncHQz1zE
ob1aMDofMcV2I5pK3F3M1yu/60p16JippoOMxTQJFr5QXrFlA6JPv36PmbnuBi5b
bsmLzrV++qLctPAntGuKpWoxein+4i6H+bKAWPTeK/+zOUR2lz095dP1pNb+NbuY
8eD1Au0ut9KApklV15LTz1eg6tARInCI75iHqgHXpBZuROKsnxglpOmZ8H7cQ/tK
5z5B5MeAH4/6qEhSFPjUURXoNAchhnBKDCtftU3aRzMwIUAg5n05iQKHYAmWT6QJ
xhvv9JXsXNo6Y4kkz3926wqu/NR/tUTdBG0Pstut09szvNmpWOkNxEZSpYC5B5SB
I23+iErXXD94J2gOV1UwEN0yRw4QoZ6KI3PH2EJTRu7ojQtx1dOQFT5l2czm5Ogv
zC+rps2w7WYf1SVCD9bcCLaYvDQuZHVvqPunQf9ytk37v5f/4uPSIC7I0GsfZUBB
fbotcXXswYwBoFOErZo5RvjTGlLTuPEl2X0O/V4H88mB6LsIzKjbfAoYUgA+ezau
lYxg4YNpngruc2ObMaINL8WiB+zeRGw9aFWElswKzkY7eXU5RnAF2XtfvqR4crsg
BoSUfPZMhXXq3wCXCcedihMOvS3PSVuZFkko6iUrem9bQP8SLVntByHlQs5oMlTG
ePPSESkeOvL1OpxBz1VN79KhChZVgY69d9gp9r0C9AYKUxor8K3rmFMOS9Hbh0ow
eLOqJJDS+YP7NVpNLxHmQZxk/5Y+I2TZjTnjrTrt9YBxgP5Nahz6SGP/tJarDiuk
5RGoo1ZKVG95k+GUOqh4KaZG++F9Pke2GgCl0GnWDbx8FaTgY2TZ3yCkfBFUrL2D
jkrhe/2RQzksYkIwA5OtkfLsAH3ru76nFVcyg9NBnO4TiCHTO+nD1JaT5ltPoVx3
8po7/934I9lg7ry8ig9/wyqo8vsq440+mvKVZhVpRagYHwG3ZxyCgC811xCJDUzZ
F7cDkEpJLJioDg1vZHlreKbQ3xSF0AmMz6esJiHL1oLMJ5MUyA/rHhhiB1Wpx1Jp
J3TVT3M+bu/J1AaQrTP3TBg/P+d1yJf5gGIextqKfQjqDVSwME9t1sGNQF4Jnp1g
kET5TUgFsarT8GTyBsBrWpSWWHf2IlYCd13KHL6fR9Gs+3GK74x7cqQTyvxEnrWs
pixMNWtD+IuBcGGvVCcZ+FOuKaiTjle4pzF5lqPRPxSYBpNza3mNwj43yUxB1xNM
JCsDWcp7S2gxK+aHtn7MSi6L6sctDo4cbYX3ZG8Wx+DU2sCoWQ5iLY20mr94UCSc
S3kNUcMiYhBXlUG65EfOVDhl/pM3x+isrLM03T3CcQbVvsA62qOXxISWcMzwKVnd
GrtQitByR0S3/Di/T4m2npqOkQV7c1ZIZUMdN4c3bu2N6WnxVWE9Oi9udIVmEf+l
6p8MHfYbUM/LJg5BKBcDFAdJUxLHS9wq+JQl3+QKorFAHWhEiJLqDDqwREJV60WW
Fm5zExUm4BnY1uquv2aF/bSUg8qvm+xmQCZ2ju0sfoEDFI/JY2Dr38ye+RCHkN8E
6sL8kmRKDIAcRY3rGa/2FshGO98Z1xQMMahWiRUsKcWUtvZmEkb3tgBnhJPHUwFj
erP0kxOKmZOkfCqDemgl+dEVDrdfArPgK4YJoU8wc1Q+RkQoelyoB6qkmVKQRLIR
Qfvq/QTCrc6MRh/HcgCEar30cvnH1RcG9bajT3el/lsd/YgBf4QPxct4+xSuCuTX
m28waHfrdyljwD0TGnBQpfxFXTnrjrE77r+mNZqN4P3pZPHYZ8gUw3tHjTzDSL5l
0OeF5vwBihXop62w0QNebg/fEY++z6piDzrz670vcGFCXutoHD1YnNSfpR+juHE/
q8dpZvQQ3zbeXls2o8wE6qmolOFqnVq+g8zIaSaCBJ3A9wEPXQYO2adLjhoDwcwp
xonkwk7zgdtoK0w69EULoBKxQtrj8By0lid6zdrFzywaFuUSJuVIcsjPm4cnsMO3
cj1fXktsR+6F2h/gee7Bbxre59N/c3dGhrLpILBT2GiR+fymFTv7kdF2B4SQIcPo
1h46wEqrtqcGGMzpa5bE0ks1sFQmAMxOOb9oXLevp1Vv+24jCsmOY0FnhF70+Am1
NUiSs5pf4MZCTo5QsDZDEcA5OACmSmhENaYMkYQ/C4QO6WMV+anG9KLChSSBa3R6
XV3pGhdspjsagWZ05b0k+XXeLHllpKE6Qss4q6fFAUj5K25P4fH55Y8fPZFdCKm0
c30gy01/3eF5Ld9z7/cqyGO9p5GvQoLjuz3IYb/E4JkpLGm5gS9nyOAaRuI+Gh8u
GHrSIiNPa61G5JJGOOrE2B3777PmbrBhJxOGgXj54/GyhKKSu0az9d5VQt0UMtMC
lh5hbsp7TB/lmNum7gQKckuzDF9g73OqNUSaGS2+AIVkA6VJoEWJi6/VjMJljjgd
GbEV1VIfpJOyID7DodwrwgXcfmLMnz+Ory3tWa7SwM/Zwpv7NB2rJAB18sUrwsd2
3AyZiR3F3xBquuVJoBRiBtVsjROeDXNPHCq6J7y6Jqcg2bIVgqLHmBy3BJekG5y5
FtJFg3GDpmEz1MI75K8SY1Cr0RWEx5FtbPRlHY8O90KB8g35ybbW4GdUGlrOBPCU
mMR3HoXzV4cKj2pnZfRcbYMmgMX8YE9mYqu7yrhbokTwJE95N7DMNcHTvUlNoq13
BAglFDHpOCYZbS3FK8ODfCxrBeKrZHxJvYXoIwWACcqyE0xh4IC1v1BNMMwJjlb2
LPAmYYVwwZKvGxNJPHxUVSvUCyS6QI4hY5K+FbZpOToIuV0wG8E5CiD2a1+6Yo3x
SxGtmPf3Fk/us1w1zPaazbIl0hCK/ZbgmJbQnWEWEFnk0RE9VOsMv6z2jgWuA7Ly
oYiMePO/d7kPyprnPEeAx6FE2/YVJ89SyZnKnph4hV07aMhUCqft7EniZvowHP/t
7T7iV7Ci0ByE+OqubMSNw+z9rlYiRGFHxzQJEnlybDfJSD2itfE8HHfNtwXUUzM0
ncmViLkQs8G0wOPNeGWu/Ii8zlFrOOypWqSSYoBOdDS+7nnBOZDtNaefq7r/simh
Z1ZWgh7Gpsud593b/DhmPzuozbzt8qdOWjPauARjZHYkr0XoHyx4oeng9IsCMuNc
mEaEf9YTBRt4G0dZgnNC/n4os6Lg+H4NMXnnXKKHMl5k7w7Z/O6acar/+rfF0PYe
6zsZwAro2MERrwOzZWpsUjGM+JiC6bwjwa9G6Vguy4FzHDUGOOZYWJ8jrc+SfoCk
Ybr0wk4T7YL7jRjlp9YYSsgIuBpLUwFVfGcZTUHAE6SyHEBZTJPz/NMIk28WWRTq
8OE/Y+QP1nid2Cxc2lu5Q9dpuHKJFs/PuvjVMtUtM82dK5DHSA9DVWy0o31LWOK/
sueDUltp6Tmg7sYSiqjTCO8/U8SN9STvDceNdWTBWPyTu1OQjGrrF+sLzqvZiYCL
owlSY7fLXUwWz5QmRO40lfYapQr7fZKJ4Y566eM8QH6xw/1DYyo3VdZmMFfWlUL4
7cuYB8X+dhVhr9BJMak0dJZDiJ9YW4+BIQqAEfw9xCYtItCzIij7ygAK2GsPNKNI
bw1g7F7AqHkSkQ/dfQ71zA==
`pragma protect end_protected
