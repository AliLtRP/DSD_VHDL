// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
tWyo4Pj9jhYya6QidIdoaTb1trqS3uEOxFgrxK0Bv2e5KjpU8bKRXZPY3g+ETERa5uJH7KWs5hwX
/bs8Sbs02MdrtnhNZDqPBbBG5lx0RfLyBM3wO6ZwMnfddnxhuentlWk0SVUEJTI+m8Q9vIe1QTNC
6hwc47NxxNa4wl0fwJIzP0EykPOFOLGsb6cTQhYR4gsFmGTuqZlalddyl0pLw2YV6vZXTL5uENNQ
VGWra5uGy8DNN1r0iljxbEgi+CZx2vkUeKBJ3LMbF6VIFcSe2QD+Ss7srCtvaSQ5CmcB9qXRyCe2
hZM9vDQ5fQqA9/Ju6dEdo+4JqZrrB1CmFna/1g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
n2SUIpc9VHp2bJNbnFXMzRWj2Hq3XI1jgNGkm6TrewefOzg9hpSYBaGBJ3aRX8qgh4xC0FrNOwHq
aTn4G26OerX+YHhFsZV7wUo2A11jWMXb+SsNy1HJbstemADFAph85QATZZLUDw1P7Vf8SBrZZfTE
MneWFLO7XnsQ58h8EXaQfE5EDP11kjgL3g3LvwTwG5ctyCUC0oaC91/fO19rFGGjh/wrEaB9q5eO
DBA9BrEGpWgoUl/Ozfivb5gH1hTPzpFilOe8ISNsIUoYOojm8KmImx5FtJ97F/kXdd9TplKzv2M3
wM8CFnrfh5yHOkp/+JcyMs78GgmHTB9hGf4fYdBvrunZHqmvUImzrPTarGKnC3FGErBr7GO+ZXbj
AYA2Ky32Pho86hlOpu/RlcpgM/2e2FJtnlkXxYfwuVnOuPg8lg+QSnj6frOAontYHAKu9pa6/w1a
Im+tAhzRkvz0PvtktkVsgGfVKx8+QcsQCtKJj6dJ9pyOEoWD6cfDjYjrmWVXD+vf1JH5+p9367Od
ojvhiw4Osmcdy3BF5fWvbc1iQT1oYH9ORu7A8m1tGAEXyQ7GlqxBlwDkn6NnxQkLfxHFOknfvLcV
LDXYVhF3SWDs1QBolxB7KtlZLCvln8Rgk86W/VkS0elooWrz/cuqWWSmDtBqCg2OU63fdnE7Nl5V
wBbQHpzNshbgY9H1my10g9124IOC08uOxTKDy0579jzl/hYFWltktxgTFT1+btxvO9OLhbT2Oahw
o9hQzdBk6RWlrHp1rvF95kzDJztR7YINe2sZHCB2mi/k8Km0c52VSEntj5fPxqVRB/d31o1Topov
6Y3GeksbugHYsWHViZwY+zmehfxQoHVgoWv8eWMmrISCe4/6yy3fjTmgxlWqRZR+7YideOKRfnD2
0g5ZdBWU+wT6yljkz5XaeWrB2Q0I54KOHCm+CY5HmYnN6nn4divsAF2waIHSp4tq+Tdac628oEF8
pjs1+Tw5qYlUWNel6p1xDor8PQ8gI4kejCSTc/xvetR+bh3k1sNrsb7R9yqzGkVclIH7o03awZCd
YkJE68CVWST3twPLR2eGGY4NZdCF0JL2LkThIZqYjJbXdwNhYYWRCPtI0xk13wv8swKjtALRQ75w
z/Pn7qPJJF8yqZl/Tg1DYUx0u0RSGzq6xq/Dzym5LyJ92+7pcojNVi+3wqebGEre9l1AQbqJ4smN
5dG6f0XyIbIswPpApcnZesvjq3Lcw6oBqLTtxhYsX6gZBQPqvD1yaudflseTNQvYKqVlhaJGN642
sex7K6BhSAfgXvGmXqE0xyADNxtekKhoksp+/H/LhnLj0FZFakZqQz46md8zDq5srz114C/Y+1Ki
/ThsLQCNcv5dpKMN7HNvuLRgtIc6kpG6mzRE4Hpg1x6WqSBjn/woTOf4DNS26oTNvF34Frg00Xqd
FO6v4t8a7oK1fXAJi9Dg9gUCtp3qfUYYFbbqo6f0OirDLL3tljWYoHc2VrPZ97UfQMMCyasZMbT1
1yUaK+sDQJ47QfyU9JvYtPFK4N+6f+zhKAKwi6AUJ/Cc3dze7cASJs4hsI+Xkcoe6G/IJxLPGD2k
8+56JiTVIwHuNvxNc2fKM86T5qTzGjqgbQDclK0bDaDu/CAl6FZXv81xryrO2OG+HwKLBJLZCa1R
0M+AH3F7OptI9wgWQHeg/JY7jIN0uDTXCk9KMhiCox4O6Qq1b6QRks9IYkVXmHBTZ4k4oZcORQS0
QFNaXCoHHsN/qOxncnxBWpBCbegM2Rmt5Oj5J6RZWsDNQp4KMyNrkMEe6x2NPLXhG6g23VmVmFyl
XtgOnIMGdtIX0sa8S5DsSC325r7LBoVsA/fVllz3ynTl2IkaPtm2Ivmh/+rCDTibElwxwzYLudCx
6oF8+9hDAQxXyZ75aUm6TzRjbVFNYaBdsTeWmx8CkQS3yV7F05rxR8ke8E1h1TIG9AdK5867ivYw
7LiNOJyol5MjE6WTarG2ldLpVwHOxZ+U9NozWU1yg7j1xEDbun9MNn04CFSRt0aIDD9xbW1kjuOE
MzFaA3twYC/hAnDIj9lrSRk6WoY5wYvdzw+hyAPFzA9VSihZg6e7I0WT47lWtAKg6HNjN/cUo5p6
JciPU+8CwH8IuJk8M5+Fql1TOaqEng3ihL+nNZH2v8KXBDT7w71p4xSAT224fzHZZLDI593xaZfT
T69rLXGGlfDrYyMY8bpLtFFqomBg7U72RQZ3jjIuDh+GMpO+Z8j7qRFlWrGBOel97m9UlASCEDQi
+grfW0Q9AGwl9iV5L28UM2GLttbM2sqFT73aFm9zYGGlkEfoB34XydwrVL+jBdhOpqYN4SR5aZvc
bu3POztl2pC+zxOqS0BF8hWb59aXjqALruNRnpgLg8+20B1F26Cn7zEWvyehpjL4eubkpEuO/Ok5
kBMnm0hFn4S/ZDkLy8FL4FymHNqA8SsvpWI06OznlIme5VO/ralqgIeGVZBez/pjK0z1l+c62TvZ
Hz70jXsE8SgWrslW4kvE2ZhIvSHGOhRAJLd/ia+NwZINRHAfzucNAnOpAHfmtu7I9DTYdnfAzti8
N4HCPGrlecfu52GgdYa7LlbFUIPcJWyYYkVErWRVTwfM0jxSlpsF5t4yipEb/yd0iVDnLysKKUEx
Ljiz4ERymSJvN7sXQgOXz4b7NlcpeJh85aG6qGJFf14e4A3V/mobSgXiJQ/xztij7Y116LKWLt4y
sYJbNPZlML/KoeHOzHo8mZllrzg57Ayya81VexkTbLzXt8C6TrdUSrKUSN98yoB8lb/LFCcJ7x4d
VRX/hNoqX6CbhPImKC52stF/0EDrImT8KLg9bHBMiI7y6TEEpMCIuqx4T6kOwujQvgdTPlwXCgBU
Xbv9jF2bTDmUKi9U0QKFgMNOYsbhsFbc5uXspZKSNngXJ4b0PUoBu7tn1yNZ78Nl5nfSt+LF5cGy
8JhoK4+W73ZrW7HuLT77Ekrb54Cfz54cv8NsgJ5EoUM9shpPg34murPCNakITkj4c6RPAMd3W7iN
+MIy0qMbtettwZxn/rHqBquoI9jdwPl4vj1c3xLZIrM6X3AFB620tKsXGdY2jJneTcvnX6mjYDGT
2NlzQXn3+kb69Jh+tCkQIfP+r4Y8Z/ChMI2BlB7dCjwXWY7/gGSLHRxA6Z2DbHW7NOjWoiQuT0J8
Oyg3KPtIJYrclT6X2BqGUTjuScqGXyhyHOyGaFUTNdxANt1bG6lVOmm16E3OSJSYdADUZBwmcTMZ
2EixyBSDci4af/ITHSWf2aTDjF55ZPszcpZO7FxKNxjrpI5whOmYyLFJsTGZZPueVhaZ3b5tDbpW
yvb+HYtHCgHxgbwRyL1vHA4HkygxK8iTdvlZztlTKxfFVyExgTCDolIlpMJZKSeEc3H+HWHY3Y4Z
eZBSQYKlwXzEwsrQ5AMyLUeWGDcU6DrGRZsALY2X4gWlfCFPiIDLjL1DL/2wrhB1KgKQZe+9+eBd
arfe3B1zCqz3/3P9MAbXCgI6y5X2H8Iw2wgGV1N+oLPeQoCop+D1q8PmaQurgqzHk1FdEFVzqIgE
c9uJF245RyZJmp+PloCd2QTXrGT6kUryyrp2DcjEVFy3UwGB2T95Rt1gwf+b0YAajZ/NBrfxmUbP
zfFsU5awmxcKYC+NA52sxp/MHi1rvz4z9DWgkXG2appEeK+7hh0SEhVek4kC2nVUlFOP4qe9zlTq
3Eh6iQZjg29lrL5Pi8atNw/DucOn87FD6xxNq8b3KoXwsewmmsXmav3afNjOECu/XNyTQORzmf5x
4tX2BecIeLluMFCuIg8Eg2QQepy7/naXIzprCpZWruwtZGnfyhrWJRRAc2B+BE60y9m8d/RPhOvC
JiIAeSAoG4Fih8DxTo3zsOsnjbtMT52PQrCMhi31ORIkb74s+sxYnlZTakwm7aPEqjfysQ69ophE
m5k7x1BGCBS86MxT62VX+81vNz0hoJ9ZbMgcYwzjjB8m9g0DK9W0g9yIOmXWMIg8aP9mq0FguR6P
Fg0toT/2fVgyMMxYwcvkIujiRWEUGTBXAm9/W1Hz6MVuQUT2vtnUxQ4B16jLau3al+LOK4/1HO6L
9J84v7Om7yJkaaTQTLMlKutJ3Rndc8OF2QWCVfyqFzSHmaMyQExsKTvWWpWpr8ODenDDKF9gr9x7
sEp5o8DVxPou/pYNpy/gUvEG2rushb/LHoFCnC7qeb1fKljCzCATTgCSpnmRT33l7gqtvxm6xmFZ
vJ/RqkgixLlR5qbu4R9y00OEOar/sFv/jJqBlym+lvigJYXqy5VIGnbK34aUDYuflA1jY+GOl72/
JRQUgNkc8HzaHYGxpSQwglq6bQ3E7/zmSJQ7m4unb050MBOp7S5ViFR3hVteNV67aBl+3wXEuygc
KtSvwnsM8bu5Zg155D3tgLR+TBfsSQhQ8Kc1qm+SUYjx1ASX0qfZjIRftKG+L6BYMNr94eySmwpP
kRtO+l0lHf450mYOFuO2Ti6cA3J1C0Fu3ReEUel5fZyxBGsOls93gJ++f/ti+t6lCpVM87MxOJPX
+/fcUbEQOZTjv5hBtRwPZgDtZJCF8o869jNbDBxvY8jgllQaO1hwFY2jOhVTzLKg0qG8YCJMDn2F
gmBzpy0hnpztZWqjriXOObAF3reZMnsfBcHFGwlGW0G6F2XIOZtR/pKbIm6qy7s6cXhgs7sWmG9a
hhvg3/hf216e9PbqcB4eMQgrv2zN2WbqAeNAl2Oa/Zy7GolnbTWYngIHjYY1vnWluE2tAyxq0Vyx
vaZ16F58Lm3qvlPFGpi5TMVG0Cgerckvktg5OorClTcoXwcv5OO3vGgDdDlZRdq8BnIY+zPxVLRl
rKDCHGwFzmh7eymAEKhzBeMdGzXET5RueFM6is+Yft5CXLllFE1JjzjS2ISDRWGTMimMhaZvS201
m3dyvzE3+krQDWhouK0JZxEg0srn53FHr6ULodLY9jr0hV/joKsthlaWvWwWNHERfJPGvEBEgDI6
ZMcQ6R+rIqCQDAjMCrKrfrnD1vwxrREdcbnhGTfyheFFCL7HoCiayYAQ8CDxfElLxn4L78595TZj
hnufPwhTTaUXR0JgM6Pf4r9xycLo+bOGv/vkxFpc3C1TMVPK9WiEI+vd1x1Rg5Wc2b/BrtlGbkfW
4r4EAMzL4bAUI8ziJPNLWHm3CnbOY5AYWfWz+t5sergTt1SIWhRSZGKXoTjc5V2Io2mcZZrnj60A
RhnSYPKS91E1ZBHcPW9kpMKio7Q5HjuxmZzinO6TursS41NwWgq1zFZWw5St15bfAGUVNJCByvBM
4Ka5bF3ulIhekqzAxffcQbEhsd3Wa88fHvqUuxPGeL7LdS3+NN4o2KFoMCkhyPRo6OKUWobKNZxe
AsNGmqQlnPidth+r2VZUIB2Q1ZEx3TryRa6jb5vZKb/CpYlJLcHsMI5EmgfokTyXD4qD5VZJuYAC
uFlb6uevJJQ+gEjnw8iEedoRyMtuW7oJWbTiGGcX3bSzT1GsuyyVFR0AJlRsGucNztdvvrAav9EM
iQ8EjD6ok9z4c9rhKAsnaogi+B6+N6I3xQwV21pt9l4o3DF3kDo1JFg3xOiJ68DHeHfd2hJfehyl
niWQipQfU5ffG2QC4t+Gm7IcsHQWIl/8esFINMO4IzxfYzNHl3ma6cggn3y5CQWfvLFKcyt8KuU3
/LJbXngs/SaY0TjOWJSYMFZ+90IHN8S/xqsOp9xa1czWDmgZRFkSVzBq7eEXTjzqnsq2FOKWnF+e
RL468FFC4cSpSuoeTg5YX/dqzMIO4NB9PP9M2TDmf7mAWW89BOkdfWqKDUXFnrrHmdtPkAGtd4/v
nl7aFuyw8aIUhKI/Q2ivVrMYW0j4uMsVYqoPNZqOzoEJFmvlIG4Yt+EVGvGzv6Gu6qm1aSpJG/P6
BQKBbSnLgTxXxeYxb937iyFbqp9wBcNWnrlY1hoY2380b92iJySCOpTigxDRCld8wAkJcwZ1ta88
Fbkp31CZKFw2gkckpv3aRIV6EWovvUb6I61bpXt6PYIKeBVD5qHQn1L+mRqNV6pu3B83MPtZqUhz
shIpGyaMiJ6oaN0lXBJJqdYbtbRdwMrfctpYS6iM9Y9G9TLxFKFVgfQlJ4Iik7q9b/vkN9JY7OJf
uD1yEc5KLDWaIaaSrO/YA9MtqUVhrjMr7kLBdObyI531SYzt9KlH9iSgFpWfeZukIQexL1bKDe6z
BuRcIJVB6VMx67VAo/M02D5xbsX3NWDje7ZKryyNmKWEv3j4A3jbhl+dHFkxkPe4XZw/GuXUQ4Bo
EmKPX3xOQGkRi28e7s2OSsclKK0eRmDaPLPt/IPQMHCgCGQvofegrn6kxekIllKB9UaYOhIPOXcm
CS4UjyzhiRXcpp4elEL04xEafSxfvpMKULy3OGuByzC7Tg+S/3Kewoh0Bm6jcRfvm/kpQrFEYZH9
1NwJlsyyRXf4uJLgCE6BADmelH2/dHKrgB4SS7EfwIERo5ifV+6qWCKca3whIL+c8vZGtu6mbQU4
Yro94DXOQYwcoIPVEltCisrne4glAC67JpeZbzd9oQQxFYKAgX6X5+mizgkx6peEiY6DaVHTjlB5
7aDwK3Tj0cNkb+UkxKxGDVQJgpVzyPTIa7NG5TXRRkipJTLO0281w14vp0AUDm2rRJ1PaB0+p8z/
iBv62Ss1kBbtsK/YURh/3KGQQPqSvC58/ubhtQ8n0j3shCiGt0dpvw/7vboMfDmJKxjJvqty60XI
WB7IYF4GlKHox/tVYEPCXClcdJAwULrjrCqivlhDxsauSNUPdrslDVLyK5C18a9xPrgAm97r8zxm
s0F9ylVkXQGreYsxIgTOcAbiVCsc4VIVTrb8Qic22ffjWcVlOdiaLG/QrJtsMOcTn8BHZBtel8kj
qK01rsa95YjFz8Hg7gX5MGYS2CcRRd89AGdiu8mxJp8jA3Dfh18PyZMq5wzyyiJc5UMk8jmePWhK
+jvEmjq7A/Ux+vXKwCHoLulNt2Cr9YF3ktF8v+EOsyE1/hsKbK4cjSDmUY8PXIsJWkgMs0YRCZqj
HHdBjmfrwn3JBzStvrhQkjKHuSntqohbmq0bZmOfQtbNE4d4mRvhShm8VjASteUJC+SijX+XR8m+
hqaIzD3X/ifqYar0DO5L2vswo51L+2D7g63wrq1ZFnjux8D22YIKbKun8PAfz0Sos9hOJUVxngqD
3ZCWusWb9JFDRep64zYDoVPgYU51KAmFLxwiBDNJP0zNLldC7VkY0EadMoIRoFe8oC9QtJNU+oLq
QFHBXpYV923PqUQ7Hij/spix2Zzy3RIhpQDrB3+vUZ1VAqzqUVuogkI9juF3q0Y8EPTnA2yQZLpq
UhEgrlsMlFeG2vmtYxDEmYkfX70Kl0q8NWtHQsvmCyYB82UeUe+OVuut/go6ETSL9IemK9MvkaON
Ou+YR4+nAetQuOHHFk205txd6aa/1xApFo8CmGQJkBgesUe8VD13kKXRfsokF2NcIjCEwigE8GsY
/G6h6sRCrReoC3HbnG1CWRCv9EUlaZHRpx8TSlsvs1TQZhR6EmdToTnM1Pho1mR3Vc+0VlELFFXb
+wM96a36yJJi0FEPart30OOUakuqFlF7qXnlZRpa8gZO2nuHHM5jvoGjIDGibNShUQRWNlAMbr00
ZaPDedHoMHjndZwZjyEUpFGUyRAexnY6ZdmLeo1ShSx1Qb4uT7qq0aD/mk/JAOl6af/haH3QGqiX
lLMErNJKvTyx+ZdkHZ0xjfxNp86YHblhqZl7deSH4PjoNd/IiqPyMAWBu9yEIb2RkbkndCTeogJ2
xX2PMAvu7BB0M0wqjsBYUYajE79CaWgHeaePT0hQdlQFYhex97drBZ7Rrh4V/tkARdLQrHudyUDe
2vJXGAe6KnggppK1pOMxuWFZUffJUZ4afTG7L25b+oDLaQHKKdNRiiRwxKCIfhifZuXdmZy55aDY
J0OwNLJ6pxEgJ/6Qr5NLH69IwUt2MBUE9uNh4c7M2PajOhRJEpL/ffdZVH647xFqQaY8veGQc2hi
JNmxkWy4oZwSA7QC0KpByLZmwYBsBhWTamFSnx0dLPN+3jdIkUgQSYTRCs+f6aQPgmg83F+84/eH
PcKhUlILlICnZq8gdPbh3Av5lJxtdCpd682zfwzpSDXQaBh7FVkUEcxk7g9NDlqf+c8jhSW4rKsh
UqWwCWx38O927WaPXlqgA12105txdcRSVW3YzyZfK4YLerIwQaTyKMgeOQu15zk0ZGqahr45dPwU
s+54l8VskM3+ROCWMoNX9xvDaQQcIz94ZbaPC2iEkdQikmu5t/ZRqp5qlJoNVHEEFuSmew9rRD1l
d4ejMdhtsFw4sEADgc+llQ+hUFXuTNgOTYPT3UovLbTUNKgGpWbM3zKgwknh7xtrS11jhZ3TWZvN
Xp2hBb9XAYWiM04E0/EvcLQU6OFwnE7lQInCU60pHZ7vTRpAVeUK/smXkJAltgrJjRSQyFJawohf
QeqNnf5SdHiD+t/yt5uW5LVHWdXWrgaUJN0AAm+uwIHL6och+an4WjBQEeuvRoCcZc7dr8lEr0P/
zK4zNptJlHTzoS5Xx5EMxxqAACs3iIa4bj6PS7AzXsnkJNNFuOWY0ueynCKixKB46ha/1ekLL3XE
5xr53VrRYDwcQO5DefOZG7jw8/uEd9zc9MWaE+Br9kEJBuS8GqrFzfiUK+vE6PLHLRFQS245GSqp
bnEyrQk4R/6ULHgFW/lajQcS08fXAHaZMRn0ZWLP9LWRZ4q9ZbSTVftmgYldp3fXZ5bi0+YFwNVf
pBaHR82GOXaYJyFKMi6+CvqViw2POM75Jg0L0K8PI9V78T+TBzXONjEzuUAs0tlAMqaQfF0ajlwl
fgxYrtStUrEgFEfW+JCKBTA6I+9aXuHdJxnrYdcwNgEC4pl5AMhn8dDEzz+2Y2Tq6k3N0ywxZq4B
VhzmTkfNXg6lBX7F9YnFI9jNlj1cgddNKNU9SDkhIhXVPOMdhD+z/NNGWtJv+FR5EwlBkAmsy9i5
iXaHa5u7tPTmV79C5MvBEIa0NFouaz/ZYeI/kD+9xMN7Bri+yZRIfV3CwGQ6cxwlzNH2iFrrlhxr
eZXThmLZ+makpCipWNhbI9lcybDVncR00v47fcemzul+CdJcG5bJrMWfYNOcxkJ7YDRRY+8xvfqH
BjA7PIWN4+ox9kTkfaqwO3FV6xonJELJeiuX5yAJpRVLHmyY4wvvNV3cpOvQSEeK9BADQLOleP3C
bPL5zqjkzZhXQPZpfnyyL4xpMBJNwDT3NrOk6jVR80ZqARWRd0lIm/qHfyVrTBTHZZvW0Sr+Wdvd
/UmI3stypra9CIC2D6IsIP6DIPjNlU8PkIzWrKpQ5oDYhZojCZhto7nQiHrP7GbbbouDWQAGgRzR
/zXGSlYgf4+3UWqp4VV4Ir5E5ca46DLUvsTy26MSOOULjra5vq+oUtVjG7n0waVX3FZ5RVWtl3R3
AaOnVem0VhkY7KiIcH5Un5KMcyPMuGXBQtVFGQDhofcKb0nc6i5XlIe0iaa7pygk9IXLqpNBO2WH
0Bn9NA0K1OMSc4oP846mjycqll5FZSFKghXP+N25x/Agq2nrn6RscEp0Pee5x/cNh+ApqVr1UcRX
lvx7TAvktAqEoOz+KrsCWXeVi/qzFfi86ku93P3gzJu61A21zBednIAvpbMlg86XiAY+2nVKnDJv
KjG7zQwiVDQBOGukADXxIQOuQlnvZAZ2MZ2weUD6I/x9WLsZpxqrVOyeGC+VkMAACVq1OipZ/fvX
BKt3vsos0XdwD9MY7nyyDEVdpJ0L1xtfuq+MDcg+hkCllp/lalTPI7PxV80wnynlBfTpSEb6MF+T
PI8vHVuMYMxaHJPoj+TycDJ9HGNZwNUcO+B1aCOSZSX8Pn1yV1nAnDGHdNmoLYP6nfMbJOexC+RP
POdUK+2gCUVITqklYmevPw6VqOp8dqq8b/ztOsnvQNrzTV95YgRp22bE38zWvmPEvPZHEndxKDkv
GbZlTWJ0hUhT5+nxKRTUR+n32HXdN0sDWwR5PaWpKQKn/OIaCswz6PXUjau324eGA792X+K/qrZ5
Fo//LCNAKwnPk7dqu/tZhmXgtzEV5yfem6xOGMmaYDfvnX+UgRppEy75eIKaeQfuD5cwV/QOI7yX
JbJ85QmuJhT9ysuZ4HpmSDFvYg4UrJbqrvmo21iJNz98vnKWR/jQ6kqKw2umokMh321cnYj9upuX
rgrcrwRYz8i4Z2miXsF0onMzsSrpp3fXCyBskkW41Qzq8kB4GAbLhF3zm+s/l/dZ90dNaeQkGI5C
U72PROrS0J8FL+7fxNMJJnITfISedeOxCZY9KsPbl2favSPo3J3rRPpskWpsO2m+L2ntRJq5/lP4
6ErTy3ffbU3hrVVKnYzKJCJ6FFQinqhcD/qs0Jvxo+1fFtG6JFckgyxkqdAw50aZvxxQQYJSsvN+
dsCvyM+/SyzhxcbUEBkOjPtHV5KMI4cpewA0DlpDcmEyns4F6JdhMvctEOGR5y8J9v3zXGJO+xXu
wWAM2j0E8SzFcBoShVzSLWlGFUAO4xs1eYGYDZt0kIRcE9g7UcOwva4qJxT93f0DgP85Pzr3Xy/W
70Btof4zodgLtXC9WIHYp+WjrbLdZIN8TjSZT0B3v+tgO3v+XHNYosQu5lsYEW8/yCW8/xMxW9r4
z2ISEw45H8aMTWhbMq5hYNKinMJtZUPF1ktw3ZJZAfri6ctll+Cbs7aMJ474/A1VARWGGccb9eWs
fwiFIxfF5q4t9seUEiUOoXb+5oLlUrzssqPKM6doksso/Hfq0Nq7Ua6pDqRjj08eNPd+1100RFAq
xMGGHNbrI0Uw0oc2/qHY3CBCnFgwCbjX5ugZBCCAviWyVgcnDH/AJemD0wqDEJPW0H8bPBjSqs/h
UYaxsFcMFbZpUjKCWJDD+nvZESGPnVSjFfxVSlbg+VzhY4LJi78X6qUOcYYJVwsmH5Z74BpHFSa/
K8Gl3zHQ+5RK7502begAGCYgX61ibKRITameT40WA/Xr6KnLZ5lDHV5UKvAdhmXMqi40rw6SZadi
xRhi+xE2etwueV9JutcsfRcKpXKZoFPFxl2QkW0RVHTkQLO72kXsEMr70oqtVq7N8Vcyyy9iKZw6
Bey2vjt1qvc517xZ1J1vsZb6f36k6DzA4HG4qpWPJj1ngLw8Je1rzWBE5Zk9q1VkbgKqWrwcaZsj
kojIIZSso2fhvZ9QwIbr5m4WHBre+3l4DMl6krdWj25blhAiyGUJOSvdul4lWcUez9k7vi7Q0X/W
gThHY987mB5ECwbSXUxN0XhUXYZWvVK4LQrBhSux+V0NF/f6ccFqwzsVBIUt8eLH/ECfe1lEeoSD
D1FMjF75EKFe/8stnzykmggf6eeJJBhtFsoBroFv8OK6L3dEZrRWe5XL/cVjsgjJZEHPHTxXA+MB
fH5mGOJzc4UjJefEmPMIqPTUFljLuRSIrW+c54OeQS0O72K1GdFCrcXO3q6HvKmvs01L1538HHo6
ViaW0eQgmORaazIf8qA4hVivbrjObjhEBiTRSCYEM4Xt9ipsnDAsZn+LCkay4xXHVNG/iOluQKPq
Op4QDCdWR5vIjURBUUNKh9f6MHa+yh1Cj6k72byru9I6kInOfmg7WFlgp+eES1ACk8yA7vr2cN/m
KkQ/Xc0ZYXKq+Ojc9WlzhuFWZn8xD1GOal7gEDG7QkPNJ90fx0CaXlPOnAPVgBOqTDrtsmCmCUfS
Tc8kwpjlG+MNCTqbSn8ZBC0X0lsKLU4yzhpsbDUVWGLQvXtUR9PYXlk7cdRz1UjNn3i+BK/U5faE
kPBqKmHeU7JreHQweFGP6t9P4EWsVmJTYROjK4Qe2PIPVEHPgxy/L2KIFfIlidjF0Ev3gbXZFST+
kTzg5ktudpqmncLW2hpEYXmvyk5h1RIx3ZreyPA9xFCZCWwD8s+/IwXfOYVa9+ViYdowqApuSNhl
vikU5GNgZGmCt1irmAV6U+21EcPhvO4GAYQI619F7ABAvm+84iCC96f49wIk5Sm3Qw7RBnRe72Tb
VOKifj6o5zUf7vgH/dsG+Eg284WIqzoZ8W12DFLfDFlBp80OWPSS6CmVrnnL+p9yKQTIwzyYbpUB
jr5DJtiG5K1nogUjQj3jhKUR1gLsqe/y1OT8AK/7r78pkUeU6RqYTrOmS/fwCa8WOxVtbLfj4XTC
vzxsMnuP92cIxIYNQXYtiJ82GlPzrCx1TvGir59QYM9CYLczLEzQiGJUsEBFZoa67uJrsBwcw9N7
N6rFHMZ36OCtyBW81cc+FfJOS2Zj8XpORbOFwzyLKk4JldRxHKOjEe5QdtdkA5nAyJiQnIMBT/Nj
ktCX/OM4OKI6aCNvizi2bj5IVY8pQ+0T4vaKRNY+se+Xx40iEWzPg37bQ2p1Oef4qCd0OwzeWU45
8LgpAa5wZwVFzt1j/meZBkGU9rRL3hN0ZbayXJiEUSl65jh6wkA3PH9VfOkPFXUAMVDzhkwdLcfl
aVAwPGini/oqXv7Pe/YBCE+MwTO8O4lt2F7O5AX0TOkOfpNGgMUhJjmOqTxful1qkALyQmBFINsg
cdQdIfxHQvMtxLnvCdwjSQMPgD9ZVxyU/fj2SSNQ3EWKBpYalmshXQ20m2+dgOtw6O35PeobnMbh
EqmzXltGB1KWIy14PGOVMgScRV8SsmpNtsRt1P6JzlNCqapSjNTC0+Sboil6MHs/YHs2mFcAgfYG
LsCjCqsedEtS/kPQcg4MdC8it0rVGG3Q90Pm0M79QVvIBw1TBu6i83vNGS3sPiN9je+reCPw3046
DQtwf6yhqw0bUvQ2j6jqVicZGZj3bHDJMxKHjTrWbj9Y7JYemIm4pt/QrIukN1PNwCk2x5HjWRXu
gh2HFB/JRPGTYdOTSnURLttkIy1v+s6D5Sww0HNpEQ8Xp/UWiHdZZ8EBVok4NWDsGvL84E3GjbbT
8dGD/ySS0lj7D/kuRPMkWkV0+llULjjF7kHib4zzOqhLH21QpZuSHnMLWPXI2MafR+7R7hSD3gQW
I4fVSEz+HxkHIXR5vciwQpdbkN/UF14510pv4/upbEQLgK+iurlhc3TrxlGtaxyPoe3F+TCJU52D
OPpYdtTxy5b63hjWii2qd9eAv/JXjPJp1L0NDSmZxF9D0+bhwoZVYKBJ9ET+PKO+eb25qhIZ3EvD
auwwG+xpr8cGoc3mGmv0uYgHz75l++OdJ1v54jE/W6G27/cRWY+Il2/NXhkhFe8I8BKmeYH83YTD
2SL5bL9ICJ/NgmX2n4155yb2PS/Mpl9B6udDiaLt+zrSlp5qgjhsRd4Wp5XyqPfaKY/NKRfVC2sM
GazxcODIUK8TkR8i/kOUhpyaei0j9sBGlXRrn5Z7HF/Rj1AwOa2kCSnqZZOhrWdAvD1c+nUSWGd5
KWFR+uWYs2bCubKaicyQnU0P41LVpEKY28HIJBNGq58OB8lvaaymfyIISR0d2yeV6gbn7fjdJLAY
Vrwl/Pz1XfbAkVVNQpQuPtCUY1/jXWVqsxyPK4J/GAbqTTlSNJcki2ah6kPBsXQi8avtFXGenUhA
GCvi3VjcHuTfGEZyonQsoTssm6EYy8iUOl7lq9n+NcrWweY1YhGDRi3POLHTS6JyHjbGhlpccEud
B+zFobQ8vsOBVPHwVL3bX1gaOUznvJVV+A6+PoFuxj5DgLLn6NEtkPX2O2GsTOhofOqWrFuOHwqw
IMVkxOf53RFFZj9Gr5JybLBVgAZYdz3Y8NIEQqkrY1sZ88obn8jFAxveCBp0eZjvalhcxGqgf3gG
XccvJb+vI7H+qeoT9IjzuxPo9HGxvysHB7JYuNnhspB/iMvjYVZItfGoaE8yjjRdHRi+Tp+m31ri
sxOV3S1axd7cwb3tQRvxoYLs9PvKmD3yhDCuljSH7lASI26YmOSb5UDfWh2jHazgs7L6AN+i5AdJ
cfsnM11bCTEsv0B4jbK/ptMFi65/H3gZpvhPyyqpfsJaFVd2u8493os1vfFA14BpcAsq5W2g4pDh
HO3qyM+/KnzCoe9qerWVt/82IwzkqxaZA+bk7m7JQJbBHp9GUSrD+4VYU6U5gDJySeQvP+/0kWIT
0xro4PBMM5mJC7l1JFqmemVXQS36bjFO7JHnSNfwleHYaWjZGK2bx+dT8gON13ozeUtqklHXEuBp
TVuwMStMhfuBEHNHzQPTBjuwG7N2D4dVEXNiD7W/aLHmW2DZgwhww+56o9EMT5VhgZhSSIZm+kfd
+g30g4UrFJ1T/rR6Y+h+UVUVG2XqksDZSrhbGidy9zJVRDFDGP5OW13rzZxjTQtvjKuFVfTx+abR
q/gWZi2LotxyZMjsGMwgO+ww4ixzbIRLwJ5cnJYNHVnCC8iWpZj9+iuQW3lguhpzbiVaJ1qEcaim
fKXimPviE3zOvnYYcyZJzCwZiETK7MTKJlYoXkTXGJEdugvcWaVfxUoXs3o6Blbe6KHOZxY6MCbj
ZCNooDfn2v6o0j3kKKVVxP76UjHOTKWNfN1meGnm/X7x9U1yiJBUbP9xcWAN6n7Fi+0a2da0pMbw
SaDxJrcXryNqGXvKmeleUyQ83y5eF1H8wYTzIllTK5asc1MjrXCKg0B/FGh1yBHbmA2uL+jPe62H
MaIbEzNOTYTWDj1xkfhe0u5xJK+OloAZ0xn/1IGuOAxT/dKO/56v045AwLLCNQH2LVwbQwGLAHJJ
7MTepdiNgatFY4CUpc/gTaslbx1LQyEnhMaY+HEG1Q3hQ8Lg775ZKPyk4/s+4fIKHHgfybaKepPT
XreC7Fc8HQZIPZnAN4Hq6gG+tkSBa/Fmm8WedWniXXCU+GN1PR7z2AMVl4ldU/5bMQEQzg/LrwMB
dQ8BgvpGh3mAbOSEUSpR/3lpVFO6misxOOfJyTzhuMLRyqgqo7WEpYyLgTtoY044QrGOBUA7bYsv
zGd8vfNTQeTTPvG2f43ytJPOXO0sWjLoMAobgSqdBn4TyGXx2vSUo/406bwpNoE71fKOOPCZGQuO
u2yG3ccndLI0pUG+UoCDBNQtcqpAxR+6GKmsg42hI5eTMx1yGluqpUUFL1mF2f8Hf58nVgEivQC7
qYSFb6A3z52DmNUJ4wqJW5mXPzXRQRUYzDd6bzrHJ0ZM2Yz360T0pBKtYApfvLpN6e2JK36OVcDT
PfBBczRzDUPaCwsmFH9V9jC/eTJQxOyx0ubGXN0OP4Gu6CzZ7/mOzuDwQnul6MDispy5++8hGywU
N/TVJEZ10PHInOPCxsiKpsLY0/f6bylGM0KklGNJuKMSkon/oYl3lyDDdnF4T/nVe5hjUajGib39
JrqCW5Bkoo1TazP48kWOqJ1+aTtMmOHBSB7E/jLwftPwHK2TDPCpsy3ZDNJAK4AV+SDFouP5aJbc
dtYngGrxx0izaxitfbrNCtQAOWSglNexlwDismAJ8MAuMv2hk81ztTdgoCezOQ690QCqJxK6Q7B6
FnfT9Iv9w7ipMfoA3hEGTk6NG7lIxXCvfNpN7FWH9IuSu3IQvNnc9x8cZWUixYrQBNBpWNMlS2h/
U3Q+4qYkB2ogU/tGBGMqscCL62p2jTVZ4NLEfhUR+1Gsdkk1wkGNQbnFFtD0XRIGHl3FdsWQDusA
ty7v9pHvvrvdwkNit080unSFei6OhzGUDDzs+8mTI3uer0zgF4OM9lSgmxO7p/fvo49c5NIXwVxI
psJ19gtRJnspFzYYV4tvrVsfmVcNXZLYQg5oDzQ9Ai2JvIVY26uPEcfC8GYpL4f40D+9OJkUVQ6+
+MfIBg0lhbYl26DCGklDBKFUenQH0ZUNW+l9uIehoxv52QJe/+3wiRHlgOVQ92hGZLEdOPjzCaUF
PkVfs1ZT7J8NBMSUce5hNW4A73dbZ/xx2Rra3yDQtQychPiPpgExXnH0kEdp7iB0ryziC5Q+37rF
CqR3x3pqnszIdk3iNOkDW5JDIYvyPz833kuF8lUsjPkHwPAPVa138bfsmk+3CKXGqT2f6ftEGY3n
3i2EgMM9t+ko9TdFxWh4JKkijQPQDX+Iti7Q6QXiK/Ay+kVlA5Y/D4CQrnozmam8OAbhVONPLuGk
j70oBa06lMwbXL3f0v0Lp+4yCEjoMi3eCUXCGHY82bjXOmJQdNZjs7ZWEIGODoYDwmCyVtbNbd1x
Y1uAFlFxvppCq/RXQAAwEWOi/ILJOnf9JPkHHEBqzQ2m0XkpUIdr0xDzRdg1asVzuoXiPO5rfzOm
W8UoEUN+9hTFmvLph3yjks5YzQ6zBh5GV7zmgFzeBLmfOhaVDVlKbAByZE166poMHYUQhIRD5rrm
1If2DjQV1YLuaLz81nSQTUTOVDKlBVa35JI5QqS+vwbB1O+bsn30h6gcPQ3eqPeDCxT4ZOv8olnk
hhoSkOh0yYv4S8Xj9h1gvDVGkITIDSTBMmQpdDTTiPPmPVuYL2HzHfs9bkvUyJAw2hQoDHmaKKLU
BdP/imQx1wBY2mLlgUZTSXnFR8YjSS+OrLv3usht+KCnDcJmaF7PTzrIKSWzoqC8ENglKJ0QpU3t
RB15sZ37kFyePKL7swZGN6fODfK+yqFL1m1RcKhO2xz6nJugT9Gn5P3dtr9guLMPUM/l69s+TG8s
MZASLw5/c9lUGsUrTKGyupj9BFPiF4xhyHL/BKVTyEO0iW9NONxBn1uebZkbVdL/byTX1pj9lqXt
pFothPmLzYr7QrqjIx3LSASn0ysvWU6WVZ+o5ytQc5B21xit1DCeQzLQKHGiVyAckSMLcAcTKzyv
LtRTSGpSMbMk8PQ53aZcKT0+hHfQq6AwMUMQ1t2qLL2KFcop76zOpwJGygMbVcuDEI8CiPXq/qrO
Rh0D1fQzhlGod4fTPq1kUhM7wtlWXLyq5JB53pPgwY7xafpOXJ6jUXT89BLNLvnmibt2IwDS0MOS
pgKoZ6gK7tT2Fm1VR5M8xZN6DGdJeRDhO1E/ObhAeBf31qb8IAT64qoTt1px0W/l/xff52cmphpG
j0PQdg7SvFbysYMuXeF4BMbvfXGVVVQNv9CIHnmm9uSRlH3BE7rc3SY8nJN+1TCmB1Q1BZvw/GrT
q6mXkt2aevOR0kSLwKuptCC3Y9gkZcfcKC8MlmNw92Qk7xU5f3XPsdmoo/67O+a9egIDckbJsvb6
QyjT1elOm4582wvBjC2Yj9Cm32QNknZjrHB995PvuEhhSJVjbg+NKLp9LLt7Uu/22i+tt4EcYhPW
31GjTQ3MssjhdHzHZhfLlP/PTcGEhi3ARtJU9CHi3hA+s9vMsAGkmptIMKLXZR4ZOW0Tmt9l7RqI
7hO5k1NNohIpGJ1ZuqYk5t0cJ/iB3lOAMaccHtd6ItBwc5k7RhZEHmfULyAsYyby1IA0XbQZ2NNR
SIsvYcm6rqLlYh7VLkWeKNJ2hSSX3E5avKWo/fHrV6tg/kG20+d+9ZXnLlA74+idOopGd6zWNDwH
vTo3yLFhBguDPKlUhtJT0XJ/dQZ4iYepwwTD/13BuBazyaNZAXHw7i1eGs8JZSqQUX266FDIUc/0
jdn6jqLVT7VMckEzGTbS2/HAAZwkm76CI/smJDuBON0ccbu2m5TPuo3sSLNuR6SOcbhUjT3r3ARL
11L6ku1sRgcwEchixdsd4Dy6MmcycytddcV3WBBnCxa8+ybxZO/tvaOcaakI4/8R0aEcNhhq0wuN
cleGVBFWZlRAeP4+eqVFPeeIF0dCZU9phjCmcznD1DvI+SzL+pQsBv1/YzGL4Xuunf9hv26QewYU
9Bjpo48RXEoyObFjTAI7v/XMz/Jt6w3+G5eBSk1XLvZMAwm3/OBvc+24rRnldGvaFAXxH0ZrfpnE
HE5fw3JjTwzE0M8nwqCpoPISipSHuolxhRzAbQLU9lrIz+Brw7bR5SuS48WUU62hWmLZyZ8FQhDu
7VaX4NOusOQ7DLq5fgxauJhGywrjuBBvutuYI/nJUxasH6AwFkQI6uvWlfHRfbMROE2rNgzVEFfZ
IIh7xJTXQCyZ7sjS9+X1CoylLE1YindFxXTneFA4gu3ZP9U1PmphVI0NVpxZqn7zSrY64/G89E0j
KURionpiVb7dRXSlBQ+IxFzDDK+BkCagQoH3arFFMPXKHvWQ0Q4gqiYaWeqmjDMoOLQu7eawtY+a
Q+x9p5SoTAZlJwymcNaVdCS72gFZ/vE3kjzwTXWz/lrh2nLiEue5D0hNlsDf0E+7bRwXZNo6mfRo
xwsmrfNhyPKhuAbeTRMxW8hTtOOF1BhwkUmycLAwMIhLKVyRJ/WMS1iLP9gEfq/speM00n32m3Dq
jC8m+piS7X6KvONhJinII+sbda90iOKQraKGdbwezrL/mO3c8rQsrwfX109YOor1b0nMOUGna4iP
dvwyERLlYHY5e9JgobkRjEWvyNLzVeFFwy8gj9CUfSK7NWmU6Zbbp4Ydr4d1xrcXbQVgWPbtUMMK
u5lq1XN8qla8SszKjlroE9nd0poYR0lPcAEiufXwSL4mGawVsxGIETaQDuhD2dr6+YbAL210iDXX
k1nkCa9yZb4rTMHtw0fBv0vJOX2r5hzG8KFa/y9njzFwBgvj8IqIE87C9+vLryXio/hGUFyBfDrY
5143wgU8hoHL4txaHvE+EkDZMmhV4JEowSZ6y8obsrjYtMovgbG8uVAf+GPP45r4NPdXQX8z4mwc
WMT80EJuXB13YLbRfXHXs9cXPQzUghR608P7t1R/B1DjU+PjvVTuAMoGI6wPt+hogWiXUScSZViE
jzUjTXWk4oz4zQCF3KwGGirld/aM1BnSG2ccWQ55rQ+2OOvHvAtKfMvvpu8Ctomi3XG3sBNoyiER
eAWviHce2v5MYOEUJQqQYhYZxTbrR5sISMnkQNxrxHWxdNh9USO7LdvmsQ5SYOfaeMQoeIo5binH
4Ewh1RHBqjy0B/Sin1AwQq0KziqZ9sI8wjuwB4WcB+OhTCSa6WKfyaJZOoT/wVeLgPDn3h7/o4tU
CCdNhq7WtvwD/gvbsQ+IGul+DLyNolCbALGX9ykjLbyYZw2VG7yYU3Swy2l9DlLx3yKfuI++5IaZ
LQhreCzNJO0g8c1j1Oc8xeoiAUZQvO1t69PVBeb52LdJhK7pFHwdpC54Z2YSl278Vt39WDIwrnJR
6a0RbbxjSZZ+cPbebIXe4jFrK8W7mkLFS3NL/MmJsvs5DDUQjmfIjJjsuJfvIHpiGMHC83WSRRYI
eUuvNQvoCILlc5YUTscEU9LRlUuokvJm0REintqfB7nMoCqMDcQMLpoSH+rELF89b4bhSIIMf42l
65Wa3rwKnUt20F2hQYgVzItlDWT60stKQ68kMY/DeIYXspDXFiiHyuMaCAIx1fY8NvGgBm7d++q/
FTjpvBoBhrn10CCkP8tkkDgBp1Y+b5Lq/ibpnY6MsDaWlQh8PCbfu1lvDy07DtKiAjv5jeKv+0hA
80hEJQtayWwP6659b30au4aoPmNsITCJ/vgCpC6jHLlEOjnXz9d6jQfK66iqiXo4KUiA1Db7f3eO
hBEtbx6W8DiC36sbRyphtfb6L+jVlCNHTpZa6ekKe9Qp3kk0cUPXc2YHmSaHB8TgGBqG6I3IwmXx
kvvMvAoSTnACDCkl+5mpS5TIWqBxmaj8LAY/PwHTwIfae7B0qseP0Chjc4kl5al2z6pwGmrMPmHm
0abwXGne1c+0ASl8PC9u4t/KR37wcVsLVTV6TmJw/fFR8xyCT/6Zc85YSbW4SKntNm8Ja2tAe+mt
NtuMY15yW1eeWT8VkirDBETv+MmdnKRFqDvGHxHfkJS2qJPKbXjq3whtp+i9EMuJQLjq02eJgmDW
RsCMCyv5brsqn4Q/QRysvvAd8hZ3UaQazBPXpWxOeBqP3chaLapHL2RaGcvXsh1VfE7P5TegLiAb
vb7O7HwQioln8JKUn3q7HAuigxX5NRbCJqae8XuSGNQCwM3r3Z+zdDjnrp7zZe+aDFMTfiyPcaqo
FRcIa7KMhE9zOvcFhqZZiZvlhVG9bj+QHkXWN0jQinwwOaddflntuFI/xez5L3UFb/h4xn/iSwdA
KfYP9awVnhj+Y1VxtLkI5ITaG+AZEAMMQLI0PwEIoYipKVEXyf/bRT2RGfeUrs/aOt95l8qvBxcT
WYuMZHmm++Dgp/QZYe8rJj5rVlQjwC01piNPlYspyN7mY6nintpzYs3JxQi0fhwb1LFFhNv4zoQ8
5ZSOVtYYhifW4B2Kso5BYbTjUhTL47yMS0VQUKFqoi/kRyUO/4sBFNjGUes9n5XHHl9bV+7JjSqu
1VNkGtKtLa+LoRwt0M1Mfwm/h4G/mITGyIk37AcDVBONBieSJ0doFth8YUh0xXagkECcJv5EDv/L
ufSurtsJCFr6lw8XsgOQ0QFyWsrOPFIJ60g/ko91RLMe0G8vpraQbOJxy2lahH8jnfvJTAoxkYqZ
72k446YLsw37jNySTJIGqadJ6hvCWqd0KFSozeuBg89uiKgm/DM2UO/0NNw2BuPJuziqzMoVjAWr
Y2HVxTmWnW3EoxLttXqtJNt5ZEikvKR4cLLMHOHbvNFytnw9JtuSNXFqa87Ngr5rBshRkIboo5SU
L+iE98Dkp9e47etK2Ay8jVlGwApIt8JBgD7nZfmmQTTaZjpdT/WuUnsU3EU0a541ubNGRYF5fWto
TlDRk/Iv1vTyP7/n7WsLYiJ51u7iWgX9MI29jMFSw69fgbacdEqtsO1B6UtWuVidS/qVd0l4Ssd3
ARkGR3wdr+i/3M49NuNrfeeEB9EMFvdwGj3SeYl5Ox2HxMFmT74Y5zNY6SZt7kSmV0MH45ePYTjA
e7klRojootgrlyivZjZN6qH7/bREKMB9MVRrZnqnW1aNG//oFs9IGY+f6+uNi2O4Zbk+C7BbN9ik
DnOzlJlz7zd+rBU61kDmz5IwTH8yIVmNAFPrhB4AEJT9PPIAnFm7+xoi8jlVWRVC8ql81L+FGdOc
c4cZ5C4AubbmehwVoZhCfgFwOa5inEGKQYWsBpDKNz9Gb9DME9pXSukyCIT3c00NXRdz2Kxr6vCv
K5SL2XAdzAveawUhmjHWrD/b+s1JmqbtTjBCkkjBcM/Y/atDQmyH1WllmvxRYkS+jDye8Icpqcxg
+D8EEkpH2bfoZPAgUCwwaa6LMBCczWsDLUqjnGVN/NGXm2/nx1Y4G3oY9OeAFLeJbvaSPoh4jZGf
nIJIu+9yNDPjvePTXBCrGv7/pxed2+NaVijtfA6PScFWef8tyB24l5iG41yosg6YIxR2hidi1lOi
jJiw+kZpKDlKzj7mVKqMVKGQprzFUEh3og5ue3c/xCyjjh/Mn/fRiEwr4bsRuYvC43+nMZk6PHpw
U6ygL9UAbSY4gXQCwtA5tO+9dXILf5daQO1LCbCw1F4nKbD0fRFSYKGA2afahrbaugmbQpHEGq9T
96FFMYXOShYlZD8+AphB5GCykTMEXKj07KZvhONDg314RNRhPsVnpohh8hQaGpBbxtWCWRmd/wjJ
tbUCeJTUtYl+qFx1cfFYoEQlt8SzUqjsyX4vlB0DXCvBA3/SgrQX6GYvQ90wUjmp0pr6RbuV0xv1
BO8PPZPyk5+xi4eU4KSE037c1cRRh43pL30u1dZvl04iiC9b3ML+Lme4OyfdXxr339UN8Sm789t5
N/y6D5BRzgeFdu4pn7Nv0Ywakhkb983ebx1h3cM7jP9ojOyH6kLtfBN2bhNFPKYFQrWbghMxAudd
hL+3FDaBwXYjxNcFugECy0qeJYdWOMfLFwEyHEKl9gtsSJfzlX3b6tTTVqpa5cAjT/AKXngoynUD
sN5BN5SzsYPrM39x1w5lNMQ4OVRBv6pUTRRJRKDYmKskmEIUjycAur8sIAkwweOFJ7tfH+rbcy4z
R9Tw7JFKBJEjlD4Q2/CXj9XfTw0F4DWhTUJ0xDaOf1bO9mQZh0paqbWgST3aaAC0QkxnPxNaKOHZ
Ft21JVXOIoUtGZtCu0T6WIxIFgzTqxRe1vt/sRGR0N80Y/Io6ZxtthjDP6w9qbw97F7nBnvNuLOp
BDZ2PJJtbwrZ33HR9jD6BN7XPjYEvB+jIVuQLnyuL4BW/7yiOBriHmQI9hARR022JOKX6HAL5Ldo
iQFfTpQ3d87UIdA6EUzEiMJ72FRzgAsfiF/Bv2MIBSxyk3UU759JrUBnvZCl8+XpLTOyMutuOAV4
Lnz1/rwlgEmNQzkCeozaquRZieptpjHOT49amMh1nzHtsyMREhzyRRpeRHqPapK3lNGLzMF7Chyc
hqGthyj4qAJIaU2B8Kr4un6wo0vD8CB85JGskglKfQW3EFKT4reKG3ReLO0pupf8YZ6U28yClvvV
VjzF2NXkf14EXfm/L1V62mtlfl1l3kKFzPJvRmULf9s2rwhG3D6Y7QYP3uy2LhQtbYQiyb15EQbx
pySQ6bseDdtWAOV18gzU36ExDadGQmJId5DnwbL2lKOw+d7eA/XJx+YtLd+jM7BGCI6FHpfHNZgk
52pPqPjJBDIYjTevgIglD9KBJ0eGP2Pkkzaq98bgmwWKMTYLrXvTjfJgylNiJ/BWQhqGogi1pIXa
Mbs1MGMwDE6SmMXzcCqyV87iBWqPibH7sBQBxmVraWlCQU44hg+TnXr44lvRuK6FrDz5Jsh9a4Ol
nMsNbaQiXlxWsKoUPExW19qtxSavN4/Fj162FQUePAd36s8sPQ5IWHnYEEov23BIuoNNuxUHIfsE
uLCT2gp+cd8iBCODFPb/NR/Cre8e8FE0xL9laQle8xuRqelaZUmmfTWJ4cMKiyyBPAxdABRCptWi
GretBq43zw/TvO2tgDJcBqlr3SZxl4K2nLtxWiYjHcUqiiHcqRDPFPG5b6EB4oG2l6fZVR5hKt+A
RRQ3QlO8J6/fB6viHRIIAWFBdmGdsG7d553tdWfoRkc87L6mQInsjShmSSUQQ11Uup1m1o7RG2on
a1l0yqJ/W6P/1qAyYwlBzAu9iFfOcDkKoiQrXdX1Zy3pDI+jNQYYeUnClqwmr9xiY3F+a5VjLZ7L
J/NwO3jNaPG5Kuy5VnKcLZA0wG7aPFzrb05kFw4OA5VEfQkJJYj7tHyQBOkT79H8dkMIAa1zYzdk
ZnueQOBFUg+PemETnspOPlZxCVhmjfZKv242xNeOY8ioJRKVW4mvqC+qmme41xwzzxvFQgh1QlHl
LYnL3hMi2GCQf+XIT2zMbIUQbOHLucX3z36WebiF16GtGGBTFzbwxu+55PrC7QOBDfUxmqHziSSz
6B3dj0X90M/dqUP3fyGvncSa0jMfDjtLzDgQJ54Z7gvpMVIEy1+BrGxduqMhDjYhwChaapqsfjbr
ddXvme3usQ90Qtl/xmhbJ7mBywAkP6c5LEogYMoTwWa7kIWVJHb3r4ak8Wb3y7RSnp5So2E7YEq9
6ay9rVYQ963t8kVff2MiUslDcgg9sWhSxO64/xBtqKqUJCgTDDnuuUlwO52Kq6HTDrVdUS87AQL9
BdIPDtZav3mWqpqmuzsv9LOMPrpQulwqtOm3lv7E7eyjv9JatrRzuHL2z9TwAEfAUbc2oKY9bDBP
HtWa99wdz/pEN6NCLwSXwtIsmB27gQDQNZWKJyHldz87ai3c/gD0pKvikXZy0vMcgOL9oifjxuQc
PMuamkJkfpt4noPbfwsAKhxs3xHAnUUyR/OeVO1DyOZRGOM9K8LDusL1kXSXjNGhK4jNfao3GJZv
s+s+IGRtwF8h411vnG37pRdc2TGEOaVgkmBFjD7KqGlzu5MIGsZpkIkCn4GNoVcrSh4qXrsc6mSn
A2/3ZTbJ6sJtNWXW4f4O+j8gx9rvqYCFvn4vQJpvvZekTHmxNXS6ycR4sHH2SLOVCLW7YLxtp+fC
Qo5jAFKcJs7IUMWVmHJdJ1NVeioO+rEnwb/5bd4S76BsIoICANl/3umMJ/ZQTNsie3vsi6hwNHYt
A36eK2lX7nDB9AdTPByQ6QipFaZHVJ9Yc0byeWXexwq1aPxj/MwhIFqj2Do+bWEp4MD9ryOZubZQ
mH1jFWpOqkFt99cAi9QxUeChuYS/wx1VVW1JywUqZOHZp3fkh7Kp3K9jG9+fZFmH3fT3ujRvA79H
TUNDzqOH6anymnmiFTzD3OJ3lAxDGudbSex2R/G9k01E1f49IHHiROEKQP2bqit1FB+e8QPQDpbG
qYfcIPMn+F9kfY1OR8waDepzKai5S71/K/wvWXKwPvYLNAUcCesfb8xW0QAW5iexqy7PWI3UuCus
QTxq/sj/lpbRCs9r1yYQ+T9mPlIaOrJoS4FCEUBvheT75ZaJ9GNIMGDQGpR0GRqPGrNtWiNsD5J5
H/B9cWHOhWX6s8D0M8wgNzABuSbr5Rs0Oggk2pYj0FhXcXeG5ziPoYgmk11bZynBeGdSA3IZaYXb
xo1Gz8HMG9IElY2NhPDF4GDIPvbUcOugiM50IJGxF5iDYTDICnw8kcYfOESuoVNQCt+3HnI9/kiu
P8kjDCTHONH3l3XggqyK9ESHXKsVDF05hdO+jof0qk0dQyFUdaODNoUIH+aUDGQLZbikrYCBYk75
6SAf+cOFM4Z3drgV6XQ4ppHEfVX4ZXlSa16cRoNJmTTZxFrlGA6WGcPqZGb6Ls41bzjDlJHHbItk
8xH2js1pbtCcqAPc50/WZUFDcoIgcftPoaPgg/H8oQtPnay1Q2JW7SVYVafs5tk0diI+qr8YO+Z8
DBYLdIbTDftdUlxiA1UjWCOpVP5WmXHH0wmeoVtZZ8k+BKiWJPlJb/E2Hsuj/ctYU4+Qjn0Gt0Rr
WZwquqvVzwxnDPCXbcmPiEJwLctye9cXkXI5aeM4Y1D2tZrD+wQQCkWNXG1zTckNQFg6/H5TU3PI
uMQQ2lkoh74H/MD3OTBeTHF94cS6uwSh0tt3USdj5q4ZHyzYMKhL9BvWn9c1ANZRgL1kkBVIR5Ky
M1N3pbocfy/jAa8HPSk12kqhr+L82vXKsNobf0G+7Gy6pUQSKBkGJNxURI6aVYCf+iC0YytW6y9f
vj01oIaX4mp5eaPh6ISo1RzQv4gAyHTn75EwyJPUUfR+PvxFt2W9hWa8IY8S/HCqW30KPwI8VUei
xcD815B8BNzXrN5i5ALIcfTw4O5kZBBvzHdIKSxyzqDEDqA179/xA7jKUuJVgdiN8z8QXRBCeAja
wQRVWVVQDkkITXnZoAmo17NmEk2JnWKnnhouN9tE3NC9Yavc/w+frlqAN4JKbrLF47gAFn1nTDez
UTRSW3OI0YqZOQ7FOQKH9LsNjtGKP64Qlh4Yw3AcXVy1AqYDlAB1qZRJ8UQkwgrDmi/i7rN5D3mu
9MgAAfp50CLPcWHDaHdAMfGEDMa6HWqlLpmJa0vOImQChjxc/Pci4bzRm7qpOCBNMnKoMy76MjVs
JeYPjERw3e6RqIq1jmHuehdG63xtQBCybhyx5fp5oTdau+pLKlTjn6uWXRH1lVx7r3O4Kuf2CgyJ
Ed+uysRm64RmsR4IPP9lEG0hy6zEXXsHz9U7eywhkaLRIfIsbNieLo/GPe4bRZYQeo3RTVHrBpUa
BqxJNFR1Wr1LGCcIpAYaHHSVwaiw6Lip8jU/ZJ/J3rRrJUvnLC6l/NaEIrnMOgIGt3jcCwgisXay
HT3Wo4Oja/Wk7HuGtTXxZs68VFYbCWUPqlBOGTOs03T3fNobR5N2CJVrpuBQCWvmSQXdeFDgI1zo
fCDZCbUyF/EdQN5qhnEYKSn7VoijQ18JLeKvpKqvg/Re/5z4s5PLz9EylA4n6S2+SCCnKakI9U1S
kzm5/PNoy8KwC4qB9syW6LhAdC3Jv1KQ3O2VL2FRyky7EI65GsWAf7nDWWLaj9nA5E61DWhdD/RY
722OAcSoWewT/GhA9dVsFKQViKGjsLaIb/Uga/NIDIlC7D13r5g4+SZ8+cGX5hB3zT3Lc2bs5Tdn
fXNl6i+Ari538MxYIEVEA15zA96VqDHaFJRWnZj7s3p/80m9RbwjwqFJn8H4LU+EXgBiCb1VMxLM
UT8a2NlroMbyiRdnKGOqc+frh1I/xVZ3aQumYXOXxuo3k6Zjm2EQwfpJJRXGGEu6JrA+Ky84zugt
OblmspfVtiACPgJpxln9rfqBu1wXdqDdxrbUDnb2pqxQjvtRD7+5jSc2dwx7clVRR2wALkPFN9iw
tm08s9HUsHbZo4WMJS/0Qjskaikar3ehnXMZRqoTmsflc46OGC2t2UpvhWFdVA0YMEgwBt6F30Uy
JTuNIUkGHX2H5PtutLY6f7MWeUfCGW+zXVI87WPg9j4IGsg63DG/DIIrhU8QArnSpvLq+UpEU9aG
FSbNag0FNzAZAmHD2yEBcAvrM6DLirGWk5OqMSoHQ1MsUVnXr5/kkeINgYa2BCMzksvBa9YJwym0
So0FvYN0lPiV9dKytNh0zyrcyUxPxDafJ66JTrTLm9EH6l/zu1Sq5YNr7iXHpbdPXDOMNC/lkV9v
GT8Yjoi8zYo/+ROh1/NLVrqhN0HTl0yuaPqasyjhAbG1D2KiB2o6+q9SID90pmypkW/w7as7ceyH
z0q2CF+VGUbHxSGcs+G6E5vSQDhA7GZWdsQWQkImY4nobfbTP0/jzATZmB6YLY61UM+AWTquWKHn
Wn+ikxt26oRIomQ/bG5fcNg/uYDos3/saK6tEybkngXIEjW9nWyMllQz1em4/4SvBDawH8cdkiCB
iCJb4wXmK66shlFpZMvuRnLswCtpDgu1lsGF++lrLpKB0byz4Ke05TQ2rb/ROifWgr9uddcZSnMC
Kf4FAoAU690M18akM2TrYsKuSZHG0flMG+MbJc/IM+N0OX+wAj+g016CH+MykeNKUAj/UzOBiosN
5YVdol1V9c5p9wQ49RgzuL1sFbmT42SuHsm5y1z71vqYpBL+2MH9HGe5lGi/KeseZTZdHFCEgUMY
fF/2iDT77iTre9zXq8OQxi5fotQFwWngRhYPmB/n4JhsyP/OHSy2jVj896SR+K20f0NJ+sNKjEa6
KnshWpMC1dZd3BXEvMcAb6L9qT1j/6+nLsuG1kS5cHtru6GHW1+mEO9WBkRJCGth6A42AH7NalzN
gfewEGtroJoaL8hxZBzKOXjBIfQjwtLEyXUjhA/JviGuPhdMZuVzA6Mb976odmUIP7SyH+uWnwiy
ooqNedqHdjWoPu6u5Tknliho2lBIPFemDCEW7qlklT2C+Ixq8gdS6Eewy/t9TzeIB1oU1BVCHhM9
ZvL1VG0w/MT+UidkfBD4BO28Ty1H3MT4oIURkBBPuS3fE1rEvsnLYM9SVpdeFOUXrF/fsrDsvgFF
lSVrHscqnmxVfvRfTF+lY5jxW2MISUTB2pKVk92guCK8WcJ+L/bC3u+HlsUDguTISfab+Y3zy+Jk
n77tnuTqcNumouxzepY56nCQ+MWJmgAP2NtwIrNPSpAaCA56FpIbUjSs8bZtXrJvWRsiNDl+Mtva
WnAYAAvIW1d/BItTuFS2YwTN86cn8zzQv//dIVsisMa2nIYvOmsXP0NzMYrIpTVrl5x1s1/JETV5
QB+gRH9LJSczzMIDXRsMEuiAJZLIkqwwBJ8XnOoIGgIYgsltfRSGXnlLsgJtEa0ntv/QLInczYXo
AX/DbxS7Q4Bh8pllfUyDav3bwDAk/PnrdkkUrwKL1UR1QWP1d/Zi9gqqd73HEJ9dDbVysHWwWpro
Lob5MFexge4wtVLVeWryw8oP7+cqrWgl74GpKFFXc+rUoHj8GvjkjmTaPk7qjufwg4GxaTQlWLMv
zywtPnwuonfVkcQH0SqLdTEYJQH1o9OxpVD5kIpSHYFvOz72IVdfcME/FvAqJJWZ66TjC3TlmxAW
+k1P8TvnAK0OQQlRTark9i9kGIZ+/G/F8dtZIhwsbbWw5+zuVQTHmqFO0555U6GXLkWYnepzqaZc
rfMJthBztJmoVpS77JqQWBx5AKyBjuQ2MLl7YxEjWyz2eUP4VMXmiNbUjeAa0DGKB3/L15Azlbgr
qPOE/4POi0eTq++Rlyq44xhH/s3xOKT38oljAczVLtGCp8Rr4hD+O3Kuk/eBF1iltsPrnUjfMe/r
mjAtembxtOMEYhiqynJMxUFTDSvvRjOPQ/ZBNh3hSAWadZCgVVpTn2GN9HYyBp9tEymvMXRbCY+U
Ud2efNVYWDZxn57i4xtyK/iS0kdGjgJCKN3uQOyfiopisUd2mfDwp/Ou85RLy9jbGtoPwRIa+oVa
OT8pKn3wlu7/RBB8Eq4oZ5W/St0f90fLyZ5fwx66G479TZQd9aEkfeCR9OX1i9X7+L3U7gtQVgJc
WNKJTUCvwwv0WGT8lYraIC+/GzYYU5N/cfAi+bAqwcUAKZ5Bt7fYwqurt07tp0lt7HaEmfMn8tK6
vRObcGrR99o5tigWrYHT+/hHexsXRqbfbpCPjMgA5WZs/Y9uFelvO4AqXfCvYF3zuKdQg0MUV0n9
JaBLTeDhoBYnC6rSVdSu4i2G3jfr/6ddnXf/eMbA00+HWH7LIM6fl4LDAcOD5fwVsPf2lJWE5w2Y
wi3wh5TCQkcZ+lye5Z0gxJssuF5EOYbUAB2lZSJsdByuAdVRIVlNvVSM8fHI3wur8VL2nk7xGkKm
Q1p2eqP608PdeXrJaz2lZ89rOGw2V8IXDv5JoKQ7+yMqBvJBv8fZ+dQ416aH9pSXowqnToCothJZ
OEvqHaB+/FcwDLAFYHBoGrhvxsjClfM/mL2oLZ8u/bGVFhPoBSZ7L1Cjp7hHIVMkoWY1B9UdIUSB
KHhc42xyjwpPnOv0MawQHkd1oY7z4/xT/C8mG+lMLjwmexglAXQcLiuVHoYvwQRKTVKgQG4XOsAO
wpXHo+9AaXHjLikVJBQo4qNVsraSv99GCtq/LY8APrn/hPrmPNGdlKy6Nwac61/fnyv7N5ioWTCR
cckf/Xa0Dm7EJUZsLB/NPWDcAgbAw5KPdOwMjhPn6Tvp1mt6VCml8H5PUhUN4rpwEGNsUWy2D+wZ
ffrpQ9cxRRiAtRI+dhGagRvvWVRfCzFa7CuwFZBJO8fCHe7oYkxWLcISPmW/K7HGcZahCAGcM1vP
G09rWalUGVDkYNCfHn3YYSpooNfzjnjQfcpjDtpgeBMI7Gs1yO+Ucx8P9wgKhYbd+fP80d1vOkTG
gDZpcy0/YEDz0noJJQHnGVROynN3icmFBslqWIypHUkFKkDCsLtT1Avc/WWWLA8llXj/LQ4yC4NQ
OgAjIf4911C6XtoS3p00IadhV87qgZR5YW/XaBynylut0zniVaXpOUmuaAPTYnhuKo5u0hsk5vrm
CN7NTRgaEbr8gWe6Mz52L8DgNuQ7iYhu5BKWgVpt3x2L7aoZ/A8B3/JK7rZOZ/J9N56GmCbVyoJ1
D1RdvtPdxNJyz4P9YzkxXztroqqzM8p6mzMmSJluErSoHplOn/+NkQ4XM8fKsJeNiuCigdB7Is/o
ZVrQCI+fBwZHH9DMdRHNUAmvV15i6sT7cdo5kxBd9032SqF6dvVkFbWKnDgFcns9QSADjJuIcm+I
XaQeQde3ueihhBucAKDXf3uUBIiQHehqiiBb180DzaMI7nMKJdxWLAx6nhe2C1ReXcYdSUITv9Rq
/XYFH9b/qWrwVkcNRtQi22mGXfMOVKW/DTZvV/VJ4+4gvdNPvzJn+rgbKs7afuA7IGVYsOpeFpc2
hZ85LaqMRWKjC/dvMoENbxMW4lvpn78HAH+Uedh2PX28fhAqLKhitZxpNWVdHodAKiko3sZWLQ+P
FlGnHghCtYWRT7SFIrCpfrZjGi65gpn8+avhZqEOhwOGGNURb0G4XXn/VKtL9IlEAQv/HYsf7YIM
aKELGo48c/xhrWnFlCJ5plzWUTlBUtL/vOVVVwI3U5t6FHEz1s67pJHfBsKfbxwb6CuSM6uv6w+w
uZiZub38l/dNjFBCFZGyIxNhmPGVBSxzxuIyK9aYEGwUhUeHZxKRrI5QblBipDoGQoG8fMXjkdoi
r96y5+vEvRUXJZ5JVqGpjcJgeW0qfvwuqPnEXe38eh7+3gPVjBFJHilBgB3ylJIOBVp4evIEOB5R
KQ2mZuxY/CLwUpu7yU7xPG8u2bvndARaBQU4PqsgmgrsEoQWhusY0Oi30FhBdyEUzazTk5DZGRDj
/NErvGq32aDGiNNRuIYEJJVGUz4dgwnlzmKuVkDqfmv99qB0vNO9pI4WpCclUJhWXryfPozQfK76
5efkGDEDpV8r/3vMToiUm0v8cwPCu9T5AC5jGQr/qY9DgQmbUKPGjal/dOmz7VTMRyaLem8EDmJS
PQ1RasmMAm+ib9IZS5s22cUPTLosYIjatvBQVFvW24V38Napt/ta1ivq7bE+K3vRbOtJqRm1QesE
D/kc7vtgdQGC+e01rKN0cXUa0kf0yXPnTaMo4FmlDDd2zwCG3WFclNLF4MApPd60ln/d75meyRq8
vyqDC8skgm7mn8/iuFMJFMYwoFqXDLCt/VBvpCae98zYlVenQVACtcm7QgKRijYZLV2BJSjgfnVK
AJ7l9vd1G+eWJrDKjjpVFO6vgBP1/+GMU2wxZ706XX5FyLzlOlzOcouseENwkfSwY/Nmebj1sPNl
rgMuIpekJtEZq9Lhs28YcFb9XG/4a9b3Q6pAK2eRNETNO5tNYcTbMcwg0RGv27oliE6vibHfKE3G
o6wAfDVg2k6/yvpQdwKUlz2bTN4c8ddYhimbMcfdwF3Z8xE9Yom+Y341c6gjOzfqrlTwn4PcHiQg
X6smiprGzh+RurvLAovRFTdBc7GrOamCSvzNILF9KQ77WuiT/8aVx3KRGR/P3i6O1WCSxNePwOym
lluIyGgRAXOS2wIS0Uely+ePwLw9x+Q/lxEB/v+R6s+S6guthZkDhHQYlJtyQNm8ZCI3QMwmkh0/
Uqd0M/FvIEwzVHK24oumZQkVc3m3pg/7koCG5j6luPD0fhcpNlVSG8Stlqx9OyjpHpeQRKmO6WUK
IxWnCBebrCefewSltcdykYvZC/Rwq+X0puG2iCh3gYlpbgaUJBDxP5dZH867bNne7l2Ni8QKe8vQ
Ui2Kxk6dBKE7IsUnnZRDSGtZVJVuxxn0ieJUVAW0a2OS1q/L2ssxSBtdEnhfZqB6ArHDSeEUYtkt
fAs2vk/prtZrjA3mVhXcrVHhXqGHBxMu27vyp7jFGCdBMxGuVcT2O4XQcBFlaLELXIIsCn/3Z9OK
ji3xkZs4v4sUR56AAn3s1AJMx34zsKRYP02OoJZi8AcsfVJ51cD+JMxqagMhK+RB1fpKxlRGw1Ey
gDC+2nL7Kf5IsDIAQnOr1zZKITc3Bu8HtLGbhJK7XHMfFW41cIbu9+k6Qjn1hbl6s/E40qGBgs68
RYQxNxnKBYOGFiWSUlMkOackT/oYdLLro80LvFXxM9KPFX7z+Sz0dpnm2QEwpmWKg7tKrDftdyZS
Wf/JWPpAIloZmqkDv9ckQV3t+N2q7nNGxFvWg3IPkWCvRoDMd2WtrQ52Xz8WP7kPy+MIVkYzV545
Cc9DZVHLzwoQUhBK3iXqi6XRMO3OiwIQo5sA4PoqBEHhzGsmg7HaNv+2FHpe7fezCssBE2vLeVWZ
6HvLGEqZpbcni+BcA4NgqRIJeKDYfHbhN5WGjea9oizET5/uoB3fGbtTSt4p4MldNH5RADmInPfo
9b9Ss3KiXZp5Q2f+udEXyCrvsTdoZGcPviEXeoMb5dYBgFqxNZlHdXC4CcmVAlI4KLD73rKOMtyI
cM0hJWeZvy6ECGdv1U1IfzgVZfuuaUh8Ckj81tLtZ1bHAx2+ghsoe/UMJiedtHRf4EDoh3bp5c2k
ydvoXWdsDRtCu7ji1K4N14NAcZxi71f9xyUjBFC82SWNLaJBoQhX3C7G2ka9+iSAUyxO/acxSvMl
lPk138IpDHFe2FbwsOVHyNvP6RAKjrcTIQLeXZ9Zr1YytXP2njIeHtfRZcXAcjdASZ0R++aXx9RJ
5vNiBdOaP7VzQl+b59qODADdxh8hqyz1s9wBthfe8IsCp41qHoGw8dPOK1hagwmuGm0ex0TlZeFJ
5qZaK3+ZK7cTRnAPLjWa5jNQha9hClqQHjhnf5id5XoYIhXhEReOQs/LJXCPyGUDthMahFAdaEIn
wyO0UHsxdTTySImIlcnYbN8KCXEZCJ48iDAL83z7SohWtqIFYcWrbIWu0/8N5EWUcsLKQlbx07YB
IFmyO+IREkB3MR3Et8VSsTzmKSEy386/sMLGTqJni4DgtnxT3UFxb/q4VYICsCDTIm7LfRgTq1gF
PsJgbz+hBq+KQT6NuyB4kkI5OmrSo096qRVcSbWSPwKXbCYXfT+1OPupCbKfyzxAFmtQm/7RrAdP
p31IxMLPuH51q4XtZmi0s3OelUBczO6s8gfmc83rt9vmMJjmSDYi/kWZ+vzzMbF0sT0BXOjWsRkr
0hcm4Hdm1KbB1tpndDuKFQXhbeHaP55sqvV9sMtc7T1Fzvbbq+jE1W4VUIWIptKUcWJ99P//pMV5
fGg4zBD7MSvnFmOGqhuEz6CLHkdHUv2HMIQ975zBNkNJ556KWT1pUrnGhw1tzlbJGwx4fYsl0jsz
jth50iXdZSthBGLsPlkCq2tE4nSQ2zHzX21GIOrmSdxw2F7wRKnvw/ymUL3BW8H2amlzkb1b8CuK
to5aqZtwOSZpQkxUiHBIFzk/eB19SrYKTiiTmTc9aWRkv2kz6T+gFBR48OIk/QAavUFKxbXgyX9g
/F/Vm8OEHTiteh2WhRxZr8CaTFyQgCQ7ya6ac9dFC0pkbvDScB2IF7goVWYtKSosThXsq8TJuZLI
r+i9LOgHbhEMjR8pxgVY3qpYI8U7XVyh2i8tSPhWaSN/cXMUht173cKx4AcEofh68oN2WVilBHkb
fKKHzpqV89AdD8iIfyt7OUwWKNXbBsuIbudB3Xvl4cfSuHZPWcMUQhkQYJPkk8EQnSqGO2igsJSe
1HETRD+p5Vf7GWSs9QSzzxTAB9B3frP+khhSE7npKGMqVAaUitvw0jKs/LewjG9BbkIgKRuWJKS+
FJIcuZhbdHfn6mGX9uFhjhymtKNz7DTLS3r42hFVg/bzbp/QOAm4z5l3dNycPLK3vUzsiNBlFL1f
I6qEzEcxwlGjOtLjRlekpCIbhM4ZSwG1FAI4OeLxGSOGIMo9wow2GuySnpHEdsjvv07tHAiiTJ1w
VRzZRfAaLR4K3jBAmwQh7Ufi4+ssELQgHOS6g3sN6R02DWpmE31eU8PmSgHSMQHvdHhEtjYkihXW
cuUxWJZfRc7wmFCNQ43Qnwjpqk2zEddYhqUaqcj7Ge7SEOYYwWyQkH4WMfMVTopkC00ArvFEA7bm
Xlgy41Ua6VhLSFrcbXsRF+2opgIMv7+40TPIGJzAjXr45Ps1gHn6VjnCnto47MDqXFl57XaH7N51
Yl1A1UMfqHUTS70fa0Yg9tWPjwJ20mKjZRlLOuv5wzdgmNLywmmdduDEMvycIQnjQWABFUPRGuFF
nk34eZIadzJLGvUiDYYJd9bVsDSMJ1ZC01DQZLqc56Fg95MPGszXl+ojSKnm440k1i/PL9EDiu1T
9XH8bDVQ3bjM7OtUD/Z5fOYnYsk2K+CYuPDvsj0qoG38aa+0A3sFa0W4zGt3rI0Rg6cm3pYbpFPS
g/uuJI5FLJdDHeZ+BrTONiI7FlfFMIF7kVp57NRtHeLIARiKBxnB9N8e00x8iirZvrXJhZYrHqRG
gFKD4gjJIw2/HFD7FGvQMLqzdfTNpmnacdDLhoYN762xX2D3xeEk+EoBqsVRnipuLz0EMPK7BgTX
E9dM4GksATy6W6kMwMBjXv1k3MBJCmpp3v2jW9fgqSz3hizgX/SMzrZBhyQj5kMV0SGfsEtTsEkQ
mu1fK28/nCiVOyL06ofZcdR/U5d1HXHQjTriIQd9tybKBwbtGgirS71Y5N9z8bE0PQPiCX4Q5Zxq
fhbw4LJDacStoFPK1aBxMXZzceqS5id4hjCCqemPG6K/vq6Sl1Z7KyC1BfEfyciNFkasoSjJ4vhK
buyG4IdiYn4pey8g8DwOZ98X3wZ2OhZBvRldUe9LB5pGPlNOmns4e8DSz4q5LBs9/kkuO84suaaZ
04On3GKgXeljMOjPlofwI2MMYcVfNYirQFstjRZSkp9lZxmCdBMaSc2Sqr0Z59aHQzYvKLhYPhk2
mYSzA64czK2JcrTdgwg1dN0xynajvm1Lx7k59omeGhdd24RfJ3TK1dlPRaVkYG1T5hQdSjbrZWwc
en5kRH5F0ml/GKpRrTBQfOvPADT/iYBCXwIgdPTVqx+yN5DGRxUtEPUIhVgQ9/8JuXiPvJ1ZjsJI
bj0lacw5pE82nCBPGB8SFHP3gwgXCV0ZJmbWuPW5V1zFqTwMJqG/xu/yD07THQ0oJfNmIRqpH0Pw
7roaBVnjXQocBpaXyCIFMqoctAsBOx++iL/+ugSHwpPjkjC/05BIyuVNL00IcK0ZccBtCYKm1Ld7
J0h3oFtwgQEBCE3NKMC4WuxM6GJGevBbyFJy2Bwek9egLa0vXiIKzssRlJ+h5IUcJDsMdaCmXD99
avL026ECD9c6v7jk4PlWzJvYrrxP6Oozrb3WfkGO1Au7JfzLlqYIJqJCr4ro9vqwqnumWZh8yLXF
RCvcKjZUy2itEu8fQmnNCnrViDx9VKymhWTjs1eDjWk9bMkj9LhMCb9hOuZFX18f6p7xnql/1BYj
wCZI4TC220nVWk1etenkNy0ICszTJ1RBVI37SP21cBGyPgkp53VwJBPt8yAP044mhifmdYjTsj98
FqbuXu2YqwZ0WjwtTgF17wle0LMBjuSKEiGFjdzh23uNjeO1qylJMBXK3VzE3/0K7lt7H9xthGwp
fmanrK6PBgCc3vnKOsVsY8tpt9vF0sEJgiNPIuTR/4PflbZlvOAO4GdDs3WZRJ5svCTdHVOgKB2n
BCAmdC3Fus4aLI7wgSdzs3c2yoYKG7ezidWRIW0FxHENz7aEeVsOb5ZoArK9wesGv8W8cZ6Vt3v+
p9tiKqzAeJTI5YXW6jxJxDqlmGHbjLdDnbZ6TEkz8+ekFguuoZA2P+j4XkT+9BnJEDyinuHaHEzg
pBysrObNG2nFS1Gt7VBXIEl+0CrqVbmx3K4oOmo5O7g8Wl0m6ukO76bsG6aghDd1nqs2Plf2NsuE
0rY=
`pragma protect end_protected
