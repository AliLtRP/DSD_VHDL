// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
r3d7NfCGKbkmLpiCZ8aCOczjvKy01yBwsPDGOzFu8z/drwvhhsz5md6qQspw/DQ/opL9Y8nKLetc
V90QubhXdqBZ9vHFxlPWEZmodZUAlk0aMln9ec0mRmZcmaUx02H+hdN1rB9/Ys0qcLsXrWVQMU6P
KTty6PYyx+2DqTnxY+HZmB7vNwNB716aqTa93GRoFWes1mK5CFt9TBMjqL93ZbJxkIdKC/b1ljqj
DsWXG3/jsnq/VD2dpQfDyJvXXTwqah29OUNViby1ZCszT+DwnUROVU9b+7Ue7rLj+TMnYpkLz6sx
2iLsCukZJUJtEIjk4DrbrZyOdS4a673wT8GWpw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
yeYGfJAORt84NVnVIz0LBeg7KrwFMenKDLCD7LOmFM29Mh1wQRXgkZzIatb18ab2cZur3g9nug9C
crbRsIXGtICuOpYTlGIdiOhbLiQxluAhLD4JETNKS1Pu9dzyGODWp1HxUzL79Fh3YxSefQ8+k+85
KZyrmII0YlxahcbHfKR3L07Pcn7rTQEF2U2ahkm/DoVjdc5fJOeZYNYW3Vw3su7ERsas4bd38/Jz
T6TurrRjMw6+ee5MEqLymzIf+tSAB32ImOM17jXQha6OdlkXM0k43m/cFEiHNvpktS+4tHknITee
KfOSTO97IbMlwwI8CXWblNA0EU/HbSFiKI+lX++F7HbAQ7tNhBS014GcIwLnN3sMDjuI0fuqzlFe
yOKbDdNQuj9UYcDun/EPyjy69k3rGjaC/RJX2F8UWh1XfPngO9YF+JXU2nMYUtspQZKL21s+TCRz
GrRHhK/Lnq2ciW+3OixKDLdynj+4w7zah5bOfsM8Vx47FQNuPvGU4lTQuYQChNTEXCv5f6RV0OjO
oCEY6T8HUV4LBHUwwS14we4pQ7xIzJlXQYQCjFzaJ+J4+rwFgEGHiTjHDz2lTXy6/qOdupQ859Rw
laDxqijmSRtRfEu+EyPxAzxIQt9yQBDYcQZoehBaRH0uWVS7HbIZWOFEjoNUTCs0CPwqqXozX+3Y
1d4jW5KAdkYR7qv4EKgowT84caXRmMAxw4tQ/vZGZM9p4cHWeui/7YZMsT6xtSJR+tDIfDKxqpo8
cwLo4EIF2xl7jt774emuFocniEPcO5cDhfpFX5zASoMRqbaIyqUSmZSXNfzhGmlEp4ySXcF8olbN
KSmIT1HwRdYaoFL+63YyM82/VPfkgvxu4wsXlrrYtNTxO/mv96iRYz0S7l0W6exAHsa1wL8Ohy7L
90+kCGxr3pCuTh293+F5iGX44lANRLAotcBk142Z/qkUGSOvtbAnmo+MVq8iNMJ++jqPLhZmXZ75
EXrPtOk15X+NEPYDEl9XsGPwbJAfQ4ddOLu/GvrylRNMRXNGghcQgY86R9E4h8lS09TliB0aQxVD
g6mmNs04niu5a5fENWX6V/ELypAnHoauLZNdS38iQFGcgRvFQcdSRMsXYWP6BpREeVY4DXzSNEYF
idNkRasPg3/NqJGJCZR4iDu8eWEzUQM24L2+7OD/1L5rdEg49XXebK9CdBnH/INWt/VUn+pHioeO
5lhlJab3JQgUlc6u5Gq11zsMQIiHd4K1/7dNjj2Yj8jn3ogFFNQgBXVVbMuepWeUrcdsmmFvgtim
Ee0CxPi0y/hB7DPeBfSwU4upjs3sWycQyEzros7EBAta+HPv1q+AQoKqSK6FQ5Yx+v/bwtMnYB8X
yRUBSQJk1nQcXlQnYGU65iQFZQIg+hNQb4ssxIX5GtWZZ+hiGVben8NSfOW6McdUPLvoQdjOTjw5
TFjyeBUk1GXFpXA7hygvA1ErCA8Qhm5gzUHQcJMKPkt5wt3nUq9r1Sf6yTq/rFFAK6qQdbvv5oIk
bX6VITgZRsteYH0Lc12xV6juQTRXypBdNYmiL9cv/4fPmWBfdygDZC+615WNtd5M69WKrPKbsX7C
SaDQPr4izlw1HRR6iMwt3G9lCcieTyuJOZ8wtt3aO9O2ojdHB+OcMg8+XDwV5YGF0lRut4dr6J/j
Wo9c8WiEHJOpMb4DaWRR8q+eQi5F0nacrv7Yh8yu9mIvE8HWt9SoSMz1lGr0VgEiESOWftn2p/Wp
UMbQTNDg0Km3IFGYAb4Dpk7VcWPo81MaxnyLCtbH8MtusnHhEwnLREjFjvgTizTn1z/5q96z33Ha
qTN4JfkuOZKh1cwFlRs3GGc1d+F2AHuG94E1P6SgnNNDF3O8Hz+7W6J6WByT2QjS7kiPgO89i+ZL
uHbxvoyVnVlxNubJ2NKGsqKuIJNzGVCM9Ap34+OgKZCY/gt5NIpPf0dE/Ckf5xIHEPoMK1wXSfio
ltpNG/staQqr1O4Nf/HDSkU36v5GH+AxFDAVTWbIMgm2RNgd99ICaEQeKOEgWPdJhz4gDYsUBa0E
bs0/QQFxUwMvzwb4D4pR+YDvgMo6WugDqzwJBOqNteHcL+VgSwpRgdRfTu662Gvi7/ZM1ucVEFqM
Kq6K8ROMVQtDGcyn/YqviQaf5pDHxl455v/L1a8OmMqBgGnsGGOFpTjYEhvS3ENCGsRkXJf9Qtpu
9RcE6F7IvZ/gExSrv2p5x2X7V/QKYGtI5XQjnoMHEyA9MNQcH1Q7FKDnS71oFEs4ZtpmvMNPsrDo
Vc2GuI4Ffgs6Gzc89+lltJgclYbjHYW/GFZFV2CoBv4BYv1qtOr5XbGayn7QKwZjyQ/aP1lqHHmO
qx6WCGVdrZ2Gqbg8N6YQaLcGAtn+H/gZCuF6jyJqi04jYM9F9+PcC6T23Xd0HDEOdjiLUwMtDtgt
OuZHF7liftpIUSZwls6Vz+PUOoDz/EOvcuHI2J8VyaPpGCn4n0hhT+3GRxN8f3TgqEYW82befT2a
3UxG/7eeEajLrxu57SDFHbsRiNTI05bR5RiDhVkWT6NJ6CPPSw+xE9XUdAAswn9R+nsrQSDUqDcK
P0L1smpbLWaPmi6P6wtbXif7fd4vpcUL5+6omR77JTxmfsoja0eSkqeHF67fflSQdBzoSsKDMSEW
6f/9rx2XujPyG2FPirpbSuk5D1rffylXI80DP6fY7Tc3Eyro1mWWmF0W+eepSBy2As1Jyk06JKfk
9iFWZMfxCP3p85ETQw1Ea+qjVYXyQ65daN8gQrIYgtLji/Y/gBaVUaENQEtonTxtpXPnemcFRrKn
+oxA6CvwrICLe2MgVBuIEWf+NizmtVpyHAbpx7pv+E6hUGsw0yW/+h4+YYOK6uG0KoT8aYvvKPYi
6XooRdVMDYqbJ7CDl2oS9dlrnEdM5rb19XKQWjGperSPC20yMSgjyuaOb5x/02m8LYcez00h1dp7
I7CZepipGHvlBpGjd1MAwd01yUEfpVcezL15kCtP3YivSd4OEUSZLWjTDfKdUr/5PKVmMHlDTc72
xzp7xTemG9MDTuaH9YlW+L/UfDDdCTFZQAp0QBZL0eGkO8iqkfI/0aG7Hn7iy4ToYe3opOiLP7ow
LOQ/Vm+iyJ0Lf8dbW48yRahwiuDX3Sc1CoU+wHRS05vZWTArXYpfp/KeBej3AhALUGFH2HxveCIt
gvyH1rO6BdlRhQX4dvU5PBturwYeiAyIpuQjBFmLJRnyUHSlnb9oDkNd40cpIKGvzgFK9nTR93eW
xRrmu6yKCrE/FSR92WY74KqBnW/cXUhJVCCNi+Dm14S+gmN/+SObBquF7HhlmZRkUAmyVSIh5BJH
OLg54epUrMa7n2nQHLq6h0kcrJNh9IqR97WzrePQAJGLtbY7hrIgtoaqkuYqo/RbAr4B4sXmoZn5
wSlfEPHy5QDJnYa3o/vnzAYc4INb4T1OnBllky+oxB/t6Q6axGDZ62KIY9h/lIShHaTyL2Cgky7m
DLBFDA1T4U6OyIxjtIl58E8JXK0GDt85l4WRpoxNdRiooc8/N65eFlfGaQazDFmFNvCvXq5rBfa9
MCUaMBwB71YtSbrXZYYDE4cvcE358btRZCo7ZurY+MdEebkyyo2Dsll3qC5atfeoeYU8POH+xo6+
Meby0eTod7A7KKJhkMKBjyD08sCD8+wwGON7803lE//9QhYkRWk5/QFQ5dUu013JC3ZPi/GqqCCO
yqD/2U/AhIceV066mSBFgzVjpyo3E+0h+jkM3KuwQgYGpUdK9tO6l/DRLps+FYDBYJxkRL6TliLx
I7rTlKTnEaGMUFzIZlNGLf6m4Rzpmbd5yQXv9eQX/HXWtshEwFWemMch+7PadfMy6uiUojdt17TH
VV4NcqElT0ecbgXpaGoM7m2am4q49C+dC0HbuoE2QuymzHRxazCjH0fXO/SbJABrU/6a1XSRSdBA
7cXEhTKwqcj1yDaoqooUZ1f/WbDNedSlE22jA7ZXynsQyKwwUKsDy7t9LClzckwF3613N0P6zjLl
p5iuCB+AtHaFgdOjflHEsES5UT3Mg8ZuXh+nYM3TU3cF/eBNiVv0vHd/sIYLhjbmSnA7RijtEGWb
IP66r/3u2CPrJK3ieEcVNewAYcBv88aKCOJtw0ukqLTjXDjSgv/rZ5Rax7A6Mmknu8SCzncVnXQE
c/WQcylpn/VnAKMuWoqc/LzUhJpYmNlhdKiChHSo1MhZdOBOWLVzSQfSDIgRPNSpuhXABZP7WTQY
p30kMwHOmmpAN+M5AZ76FBNeBtOsOUTMiUnWUbWTUDney0S9cQZaUl84sG986Jr3mmLjKvNpw57D
JqUktCYJ3Ut/LimbrS20SLBQwR4KCoipkhwQwpx1LTJOm88lrYK0wU+sorNQQrC2FQeyHJA+OaWn
1s4VoOp49OIWwNM1VyqHUoHiIBxG2Jau37Gw2WDkEzp5OfBfTJy0qAhOBsvCr80F1rBN1iABJqZQ
cwjNCnt9rgOQVkxyUgap5DUPExI+1U24gWnOBzNBzsrd+HjxadNrT6dROQwcFLBRmP1OL5RrrQMh
UgHmni/nnmTZS0fOlRtjRSyasaoxj3SXfn2eKLpWD1sA3qVKCkj+87eiEcwAstMyJphFNdkhcka4
2zN9MS8DXFDeRP6Lhn3Mtx0hMu3dVYQheZtArENoxyUgqRLJsrFKmd+otE2Se7tUCYNJmZ3fvYnb
N6sJYjN82qm0IGVAb9gF7KdOs4Mp4rDMlpaenkr89xI/MauoWhD8o443XDPEGiH2b/vSbsGtFbvf
e5hA1wrDr4F5q07ZD5HzuabvvuTqyL/+ja1pigEO1nGYh3XR3Tdv1W9z6My9Hbi7ljA9/AHt5vP5
CjBguMxIgCI6KmAwJ7TNjprSPwe8YahAaKqFA6EZzupfZoZIRYkyBKbZ51m4AVJx5C+ulwy4XLh9
V4ZS7JmJcEtr4ar5akzq0RoSKRQD4uflO9gD9c6PQRQMp5N/XyjcBCNdIMHGGA/iEdvmQWKCHc1y
lolDHnXfTsJX7fcowUsoEJihPox94neyPtDJunZLtKZ70pVmf8F1fT+a2iqUAhf2c11s1b6bGko9
wEvXU+GeBe2dev6oFL1GAq4UA4SW52AbzOY8WXhVPsxuwwxDCknhENMNK1dHXk/IQ7JCdDX18EVH
BPPxGsat6PddRigzN2jh4N+YgsdUjOwxbpFZcN+DOyKqzDOyQ9+8kTQGs2rSzYeKe/EcnN1WegRk
C7UoP0Kl7lvL2+6FWUr2/zod3YDyzipHsF6y8pWc5n4KWlQBzJJWTFzUaSvyjrmIX9IyWCpBaOMh
z4LlXxahxYR815O+wx6MMTvUYZZWPhFhlqFScJEQCTHO+vZlsghmjOXZbheQpwtUDtwhlRVGB5TP
RVegT+uHDK8c0XE3R/KPKOuk0wOFal9gbqG0KHoBL7reIdxeG+T4cxEYyrOZzI0UP0zwYxbQoKuw
guoU/2ZigcCP3+Mqr3gpoXbUpDhBn/3Zrk4DWhOF9EsTUBvrD0biXREMvJ0AFDbv5hhoI9b6c/Sz
LEuasctpNGiaBPPqBSMUXIQuzVW8mH7+Hbd/Uu54vvVw20D+jesEiyqzAfbmhM2WFQJxHrDMYN3F
ph1U+JbBw4lglH8dd9oDMtXCdGC8PT2b7K6S63DnEULRPWHn6B7gDIHf5YVKoaz+pPycSRdnANod
Bf1Mub93jYzBIeb3LkNodaGoWCOWc0fCadacxT4m7xm+Ewx7TdQrZ2Gia7BZaMpmqNJJCqS+mupT
dPJMK5E98uDDEjb0cy3Ijqa/K+pKjrPjEoZ+N7jbAEkG1Jp7QcScOKoUzV5zbhqa2UjfS06gPpC2
gC0G5WGNcYev4FMySI4QkMRRzrQsXPAQ5i3O7uk8DULpZLpgN1hA2d+3mg/YRTTNg4N09J0fW4S8
OMnCwuV5JCcH+VNgH0j5DKW/4p+WmcirhszDexa/kg/7oZuEB7243Y2HSYoqY8hhx8jhh+mufg4X
aNM4BSGp0dajTSeMCVfbPP3Q9r+jVwE2br80sMcoznW4pwJ9dqsKv+REKrnPTmkxc1Oe9lhwNJ5T
juISh9BuOZp7cjPbWxOG44zPODr7irkgnn+s9zN3TkzekdfsUTnSWYbYfJKKqGyRK9b7cgcSg2LV
8Uhy6x6jVb6aedcwl+kujadEAiZiubgPe+Uf9Tm+wc8GfmBWwtAMEEN8kVRL+5jk8k2sFrwI9u0v
0QSlBpAORIdeg/BgnTzF3zEVCnZ46okxRGKDPHUzaoIxRudzONSmK+2DeWCwC+Vsst7fDGc7AscS
0WUQgC8ogc0IBl8HIhI8XIuxxPvhztFtEUYwqytItSenZn5YDfx2KPmxCJZ6t6j2v5/JPak2GfHk
93rEvSyD8HGvCYM8CFBo/BnZJA5kHEjz9FdTBImg3f0/BOTNVBN2x6Lla6DdBfjHi5ZeCA0fcj0N
EiaEUCl5KgWHkAncESNKO16wgOQK0lxmUOA93R+yTjYCvpGf7omVWwbm9eHkvTtw08Q/ZGlheC8u
+FaO0aP4mMtSuNDNKPVUEr3sKS7z7U8dZ35UOWlJf7wzNOfy7kKtD1iWpPfDf1wmzhxkj7UOm+5Z
knVSd6XpotrsyAPTXjkxkoyaAF/T1mi2CX0iMpC7qI3PhOBTtDekut9l9RqYZc0jBfKDM8onR7Ip
6Q1FloRF/mX5mNhoYAX0DijG5lI/ZR5IO53j3xsJiv3s3BNpyeSIagZ1s5Os0VvK6qN6kpEbo9rD
IY8Lae48vydojb9YPx9P3eTXCATIWHRBokrfn99bhegTBij5M0ltFaO51CroHI9ILfwF7qs9Vjcx
CzDTnAnULUsg7GRXdJpFKQKGx4yosGOYJODWjvMaK795S8yTmYBkrr5qtnk9RyTa1E1gq6rbe23e
w3rthB2vqM6/N5XQXUSen/VhmFLQRYQZZ49XapGTsiHkY/58kZgYUbFVLnggb6QMLbRGwhzVHx5q
cbWF7yhU11TtZENTWXhT0tFIc8FT55PbimhOjL5jpXyl2DMTugMabyPkkconZhf3Pjaejnx3WdOG
eXS5Pgr/CWlD+/JC7dnGPTarhl4vXgBu2CxsVZHaGg7j2IrEM4+W6fSVLDc87oDC7PZinFPB4uUL
RdO3TsQkNAhI4lTB2fh1c1G5Nwzo/mMmF7q8LcCvAT8OTyLG7X3gE4TFc2F0yxLfulU9fLL7ybkj
y1JkMzfQfILPC7xZfraHGUO1D7X8IXOEhn9cAw0cKevfHik98pxLKqs7FY5C+MuL5ghNEjaQUhmI
jFslyJ2KcK6rZRrDfE/LLZ4NLWkcqhVuTnd/6VNrr/TFuoJc8LGxWJWrIlqqlIRrKv1SOpfeWN/A
7VBRTis1Fkwb4ASLnjZB2oO0GbfvBVw1sktGC7B01i6z3xT5HiTWg51BabnDqiCeQWLNlB2WDDmk
DsAD4nGlxgAQxSZOqPUdwO39AkhZUdEdFGfgUfRC/aFIYZJIGE3cmKintaPjS6OFW6Wu0ULFN7hP
zYDB5O9gijC35u/jsRxMHJoov+UXWWsLEzDFC8l96hfsDAjEi+H610sFgQGTOafNt8ml7+GR+Z0Z
BeqZXkMBB7oabjA3VD3s2nRjepdvzn+hEXwoWsZyQuctOea7jNNQXll0NsInzjagNdQp6eKBVgIP
7GsQoeSZFs64Zvra8ob8FM3DSWrlNJlqtXumaW6eamVqimg1C+hUpsqnUH3LwvFa9RCjzr7hu2Qg
bvVCGZ57P/yKh5UW4urXwyOAUw6KNPSedcR3VyJ+404EIOeGFCEtDpDlBeF76Cs6PBTXSb3HJ1pl
PuRObPK+io3qoKOldTOZ44JamWWZ2GijZbNk58pfCKXelQw2uKW9I8wyWuP9cYBmdbF0jx7K1FiL
waXHBkZ9IKrmn7PXrXUxYbHKAm0fw/8AMFghm4yb4nzic/QUKBoJqBUVseNTZ9e9iLZG7z+reRM4
d279AjfhhVrJYnQuz0UpyoY0G7Zz7L4xLi3OdVyelcu74wsey4d8fr71zLWcKyk5/mbNDzsBckcm
n4fBaHM+bYuxmanSTQ+OutommO8/dmfoPBhVigN+eCYAwMado+jQlO5Dh5llFAGouT+AASgkeTbz
jzOWZ996AgMkIEz5XfzX70l+2hIFtG4NVG9+fGQNPsGtk52zQr6hHJ1sETqtdOfqggM7I5xJV7OY
DmR7LdvDQcy1tfblRsirNVvql+eK9LvVHBalmesb9On0UNS4nyiR70D6H5ZHg0Q1FV2/bVW7g+ar
pspW8thwozVR4dJlLVGPWgjsDIwJCy4UjaZ8Rju5NaMyhvXbsnPzajaB/o+0mVhIumcQ+BJmMZHN
emWWo+si5R5iyPgCukti3/bycSjOTXrrbaUMg5rRj/6Jd70p0oJIpidekWK+Fk9crBW+YjJo4ZdO
ptPc+DNp6ZtAWxzNZJ2Yh1u5c1urS1uUNJ5d7YVdQ+kOVNI1F7KDkcakMm4XqfqbFpbFaJqzkk0o
pHXtwp2Ap9VeTXEnZlDSeu/PxN1+33Bb8XDRymyfLlDxbvdEfIWjFF7iOwMW3cgTXKdKXLejXi1l
g8UP6Z9gtQGm151SF+bWCY2ty2zNpBC3745pUxW2X38Ab3W3rns53WBJ6NPfslM7TCdhuxDK/Vz2
SykB9usBOYnbonJs/5YYW5yeuiBVwxCNp781h/DTwWZFNEf24RwvAPfDIM66GhzvKQTtIFfCHQtM
7O2BNUboDIsFEqxn1qjUibq+0zfdOtBr3S5bXRpe2mOZuEVpi23h+auGiQNhgdfZavPfwouNwIcx
bxBVcKQ7AKZS2C9Y3bklTTKiO2jug74tGYSaf2TlidxVSPxr+c+GW8gIm/qTJ/JD7ojFUW/wtF1Q
1dLaaI4/ufUxXiLsFYY2HITsWqKqgkhfjflyKtfxinawuYpbo0I9sgJJNMxaquwUJPL0lMp6KvRb
8SZSO5z0UvFcQcXAGweTDpZ5523ZiQ4H9tspzQR84kngbELuoQbNdeolsRUBaeVqX7xlVDaclLhF
1s3lNeAWOyOK+pSA8qHwy3NRV3N6GWkTIJ06FJEsqDBrQtv1jeBLSVxTV53BGtCGSkLrCKiWc2e7
U+0tC2BOb2cAMv891Z4ew8gApN+f2iFiUoEkrdZbyzgogL7fq10FEX7TZZNdg9Extd3iq+gOMdRe
tNw4AU9UkXnxC0XpC0xjwqQN1sMMUdzNwUTOrs8Wg371RbNuq8BqmBMRVs/IlS4hN0L8Xr4GQp4k
jrs7dgstVJHMPdTXRwuxAu9aD41A5m5d/7HgUNfztwM/fAf+USdxjubflHLw87VRO/LVxZAf+d33
K+o5+spdTddnOdm6lwqCSt1YMQqbYtRtko44Y/eMVBlU+Ef7KVlW25qnncvh7Y3TqhYuICA0I3NI
rTadDzns18Cs+c4RuSN+64tfqjiPAbR22nHE7k10TWdBDFL1qNrbbzoIMQ3Dcgc/C2w5zyhTr5Nj
+bl+NQgBATnA5qMFlqByDNsPLBXQt3d6xvGiYoHPDxhy0imjBeh3rsZbt9cc+ylSYRWZMpmm+eHJ
VbRG8gDHtiNtk0EhK4s6+ezE5FOYhhf5xV1xD9sIYX8s5ycEcXMWAV6auVQ8Cc47SmJQ+HhNrKkF
pw9RO2/V7kTXyvwRWNAqnQr4XSsElBAFVAvbxr6w93cdZftEqj9xTTBIaNBjvv+M+ScT4LlVhTdB
PC3BTmAYM3QdKUw15JwMJfaIYMHjb1kqXDbtmSBlZxB3x9d3wZfrocnC1E3RMD5No5pnSajPBy9q
W0pcWFH+OeMTEhFLt/ncBVNqSilMBUUFdNwiS+OQEQ3u4ET5tQV58QTE5Aqe+fCwjcK/IPFdU0fY
+n1D9yetVQ+1+WYgNG+/1mz9yfc3I8O6oZPpeNgK14qqGkVapVDd6rCJivejtAdT20e5zkNeuC6g
cfteDPJ3zuGknrJC2h7F4R/MufjZfEQuOgxQuKe1h++ClLIWtYmQu12Mklk7q1XRv00uH9T8yzc1
DrAC1nSjtigkumeKzrCHlpf6lDRB1h9+NpPL9NwuiXY6alyk6x8eGUK0zNhKuhMVtcwBJ1oSPifl
DWuvEa10QxSxIN1p3dlcLMXwMKp7/9VP8ksrGxmc6ru5WCsqV1qcmeAFUNabMFu0dwwOS0u46IUe
3kZQ+yHG/KBW5GGh9HcF0b0DPtxT/gQDy4WQROWugtqW1fHSBzO5K5B3r0B4Ai1gPgzpFR1Sb+qI
4w6d0om4xy2bfxYpjB+GS7NaUZDy6m/XomUXDRs/O6Wguznd7P9osK18c0eqlUTvsIpXOo8hreF/
npayiuMDYq8r/YV3lb+Hwl37T9Di6hjY2c1LdF+kginoOmvyk7TAMgI3pKLDJvJXNifufVCD5O60
knfVFQrnbbz9p8QMGYDJzgtJJT+pMEIEpiBvq6MYT0gF8rMU5nLmy/qZc/fSLllChn9s8Kgjaa+G
vZ1yj4A7VqByqVwoio1BY8rnA6TjFdvZXaPW34BD1aCcxMLgWd90zhTWJL/TY2AUw8wBbqzVF5/S
cGB8mBiXh0bsNAteNyJsshqBVuEDC2OqrazGCVL2UItvEkRLIIPG2/0lzh0qJzaFQmZWIsrripdR
YToGvWIIDo+lEdjfyDJGgagYdxJArYsWaD8KZdlXkZpbRTd8n15xIZzGBjCwbjpnWo4iI0l/G936
wFea+yrRpXxChSjUv/tL/MyG1ZuHs5wR/oVTTcuyRc792iCzKpynCsjFcFEycQVg+bLSN4I8gvgM
dqaok0SUBhgD2UUunzhcwagoTk20kJJk/cxhEuyerxHNl4e8OKxvjVI8VwziWkWSr0pbdSoKO3pE
r0ABZEh8kIx2iTuvnJMPpg80Ux3kWIa6tsntlLQv64or3qQ6eiBIQxyeVNKHjH8D6b+ZbTnkhtwv
gWLl1PUlouNPB3Iv/dEiGD2ANO1e/9VMW6A34U3zJrZcURt6VugjFlR9t8Yk26S4Ek36Ii7DomwO
8zmQ7+Qm0Rh3dwlUcDXRcUWb4pRKUlMlzJsg5bqVmCNhoJs1mh+t2X1AOJjireWqVeQR88wSDCcR
J3dWvrjTtya/ZS1MaTUCnFXvwNDXiRvIrJXRlqnhDVOQyQ5ZffwgEvFa0WqcZ0RPP5Q+VCOK7N0j
au83FK76gYp46UJ0Aq1fh+lohQ0RJnUfU0yajqgNSUT0mDNak2JN6I747pJaSnXH3VwLmAqnAlPg
4+YufhbNQ4x424/bWIMNrLjDSNjzZPeGeLph9+oQvN/279rl+29imZoi51MO7MY1Orvk23mzZIY8
sMtgmuvXhwWim4/HIi7rQjeAomyFN1susyQm3IcWFV/SOkTP2CuuJMJPCQkxN50csTvJHsRXRFFW
im9gSLgkXpSaE0UGUScobZ9/u7a0NFUru+JDwMHOSYBgRLKjEPWsL6oqkZdO0xMy0fkCDF1yaOrz
79dzk7ri/2z7K0OE6MZ6P9cfsZrLToTo1QgmE7Nwm7igxgbNAbNTaQ1vBvndQFs0Bu0JMY2rA2Ct
M97HIpyHfoDeoscWzdu+946rKTsijeC2Kpn077NSp1NS4vGqFaMcbY0v9rCm+hJH5efyYd5jQjWk
VCOHIxmVUKAbvQ7ydD8FSDIM5nk2e91+4ctDVmKe/nn3ZSYOaelfX5NBWLZAgBOjanmYfdC2VJog
umuX57i5ls7SCslXFaqAFrLxITT4ivjGx3HJ5axUiPe1BbzEdm3E/aB2Ar0UpF+oz43nXoBaRpGj
1m0Pvd1vxmMij2GF2EzX45o8yFhB58yV5Kfd31ohc2Cv3BICyT1trZ0oxdb9TFZvnJ+XCaiuYc38
2yt4qPkscK6nyplMLlWPA8PZad76wbvz/KZ8l9o5ncosIjbLAcsPf2+OejdMZMD4cPg9MUCd8FS2
qhfk9JJ8Aqu9rzNclyisSh8B2dfaFzNDHrebKHt+ulQi/XXUSsXOZJMfXBfsgRH2rfuZn8cDy6g4
QQnamI76ZzKYNmTscgTzcKLF0tNOSIT0Q2lhXNbdFk+tTml/nJC670KIX+0ubgjVSXuOMvb5WsC5
yjG+GRVzShcNeByK3TK7nI3DoLcssShakN9bpvlRrgK2aVGQgcWppFJF+sI+tezQ5tgRHoSZl9+t
4FTpat4i7c7Dgy11pxSmyohkqrqV4yar81Wok2BQpeClTivPY3DXz21b7wB94ME/+st+ooE6mvl0
rE/fyK9/+fLk4NcEeA8Y1LhpC6GjIkEYOuSp/nh5lLQXsZfJbnL4d6akYf/mLKdbEVTszuzCktPb
cTOKsW0ojLJfkaKbmHTkox3WJy26EZg3IhxUb8fhV+zMKv4SvCW1nXixRp0AGQuuIpiIIyihhDc7
Z+1ZrSa1MjjAMV3JOyabETkSFnTeIp+WSIFpC0T27JL2Xo982saxpJ1cntCHw6Q8Tmf2HoTTEyLI
KlU3JQSWU5+j/KpgSRyXUKpABUpLXBiMRSx+gt728B3UhraebNiYV6Fb4ZpNgjtti8/8xFYt2O1n
LeYZ6vF7lTmjQCXN+hhLHe8r/2fO5j790nNuuIc656/z5yttGk9lKRhLCAVc/vQbz7uR4x5pAn8+
BZac//lFit67FAqiQXgXv0LKAAaKYUDeBTnfr1s7iLaOvFlFwHwRpDwhgZqJP2411xvWqOQ5bvFD
lstCajHQw14ODmdIVOzRpid87secwaVDmFwpvhQo/WdH9VeBF6dl6iNs9pAImrVNUWoS+qOmsZAg
DnrTY1NBiKIdvuAq/dfp5KoIB6l3suxGszgVl0v2DHqOfYt35+IflfdHFgQDHRdl3uDNPaqoCcyr
yqFo0etK6ANdo93DZh8cBjWzKvoR3OYJpPKldOiw2Zote8JDE/xZyWBNBRkW4p7kTcb5adWBf4dT
ieo+CnDfmNMUDKMo4dUO8YXJiHFgBOerl4OC5z++bbMkmoKnHGQ4zGjfRD6Ta5HfJR7tmOcseKrU
7Ux5zqYKEVAa9PlWljm/iBZDNBSrsuf8+W7W4LxgBqnyc8ZN1E7f0s8YzyDlQOo1M4LbgM4u1Nsc
BwLjWj/C6n1j8cYYX+qUc2OWipbyjRu6TnaqsP9AruvgKRbmV4wWG0pJzIHeg3UPsBRvZCMtlY1m
ZWnyDjvRrG9cTYMLih//mLZS7UJ9MtI2sd8kd7qIodfLOP0M3i5eDpwcBBoV/yAcBHwRksTBRtVG
Jlss+GrpHiZGjhC5FMov8elszmHGQoXWwZdAGcvx07osemSldqbFCoyTkmJca7/k8QrP0eYIBTgQ
L9KJ/BBJBLGnR7sdH2OC9NjE2cVSDS1jFxw6KeuDcVOpkv+YO0dSto5OeHACTEbPKH3/6DBxuxbG
4sykgn7y/6kL+VCYuxtnZlG7lOgHLMYhIVD5PKA6SM/QXzMEjU6wXIzApurkjwZmYhW8i3BtpZ8z
Su74cpyJHRSAX7gBWN7b1h3L+LA3YIxElstxVn+WWBODNcIHYyuV7gCa6yusgCOVMDGTBEbCQPZJ
rJ9BuUYOf3IgRUXDT9BRzzlJhWcMbqQxHyyYSql9etJln9/+A4N9gf4G1zEx5CowreSYvLGIGWW/
+OUIO+AQJ/EaUwhJ2dMIIK9pc8/LCGYizQisP+PypaiiKvwWV6OPl3ha/9lW9iE/hXGDKCNMLFhk
I/NinERpcXyCRS6NxJSS0pR9VwC1w8ZsF583cqM4lXqfqRFhT5ahG4r29mtvKrTB7shwcEEceCeW
v7dl5hk99bo4LI/RzHJYZwQplYcRf+P3JAeyUC1/fE+hqJ8AN8U5UBDBH4ptWxn60YPHq8C1/hiv
EMtP3uy+JdjR8KfCO5GbTwtWVk/sCZAJSdXDrahfT9GWBJT5YTDSZvctIqZ3weh62XcAX8Y3dAfW
29kvJTlTWHG9Kt53AJGFDBGJgRuXwIzm1/lpUxhngIdv7Ohl6wm7eUwBI4O2Iq14Tancysg8Le0U
1cCdkofCPjB4X/hFX3ggBlbD++fL7LKSh38CQ+MOFT0iQZoeCGemcqfSzVhdO7QwlRPD9cLcB1V2
wBBoiZuhu+hByubvUG+Q3fuYElP5fE3BuEM4lVzeUMk/EAV9goIc79nJ+oPTW1H4lh31ZVoBIJOS
H9hF7Q0ComQ6PLchxVOqmCPicbmJDsFDnqoWbZGEKm7GasKl8iPg3PF8OpT4to/GWkywT3r3Up7c
rh3R8seh3KT/QtWyXNam7cAg5QuYaJo67MoISO/lKttOMUQvnufK7Bu+0hEPtBoQjmWhKmYh2JvA
37VIpo1lwfY5GYuMFemUdZ40eak4PFOHr+v8QzSZ3q/UsmUzIh+gTO2PpWocU8K2KiztLuTeoseC
gW/0itwqs4hTthJsl3b4U1D+7i4O1dAOdtnytEo9BP0pttE4Fe8ORKteEQZnDXSjaMdsstH4OyM7
U3eME0uuaAIQfUzo+DbliGZydkhGPcOm9nRtuE7Hmz4c0oVxyzQa03n54rjG4FDnyXVo7tEqIav2
JXrbOsCUjlQN91XcytFEQQcOIQh9o0jwicBMzEK0HzNwlGamqhKtGlWotNnFE47Ii2THn2pAUAtn
MfmSKBKWVglp/fqrweZZG5gSmAXjBmQUd1y52MKvnV9rWp10GjfD19F3afvZo7F+QfI+D0NX/XMT
CNTZNv7x4p5PjK4DUolZ5+xH9ZL7wwzLai6nw3aKELtfABs7yzqRfkc1BIU5blcnZ++juGnHuQcG
ILi0b+EfmyqwraUcTNnzRR6zJSS560WJWyDgKk/TCj6TnQ+C0r5MeGqUvjx/CSDMLZrjkWS7FmZR
/ELdTltve7IJowxtbmost13ZDwjaLbVQq+QcnJSDrZKoNSM0Ko/+OWnwNEueyQ2ob8C1zYLgWcP9
LPaO3Vku8DBoAdedG2eaBTG+QdaNjEeUFgWnOn6w9dLSBiqgqqTAbUS967J6Nk/DR7b5OT40XEMd
xOw1lPOWHFhffQEjEBZGSJcx+GdnDzjucGrQOy6gUBc0/WtGJwNx2rAMLP2hx3RvTuVC1+O8e98x
2I7G4wl2lGdPwMezWvkuX0uzbnuSsqJygZ/7Y5wpz0dAXhYYjMqdWzOE+BzvpoG+XAkkDh6UHdmV
xT5E3FgmC08OzyaqD7R5wcqgSN0h8TrgrxsxdZOIG4bI27VqZMCX24joQex2F2nHSvVjdGGip2wi
qXb6izudDFnZraiFyRtfAfvYJ0ev5nk+HeAI7Lz3gHSb2LQdmVAePXM6V/pWudA6YFn3YYL/MY0g
DCiD7XOeCUYzFMD0d3ZPV9F939ZUaaFfFKTaZB9a+pVq6YoJUvYq5U8scP1BrL3OmwlJ4aYvykeF
Z1dRCQWIYFwHdL0qJIzR0DKjujFKhE+4alqEsukYeRQWiJY9rN20kPnWMLx7XVgJxBWp9b39V1tB
CmsAl6Ci5NlnAUPNQ4Tf5KDi+jjF4/iCFnhiGITlzhYF3flxDJDdQPiInqWVeGNDXrSVOXw1TMDZ
d+ZTx6VRWXibjTvnB+A6ImEn4sVe9dYuEmKdWJqP/sNLh9mkzzG+dVNTjdxnC8ER+8YXgRdMC04P
Y2vFVgOZJzm5ZMqxnV1juE2Xe8RlQQW3F07ZDD4d4wn7S5uBubj6rUL8GyGEnzV7+nYx5yNd8Qxa
g2dUE/ueYFawzuQTga/eW3VoHErSqW8d09IdsOAwWEN5mCi+T5iPcqBQu5egJJabQ9BfYfIDpTU3
WXj8uUGX1ZTgTLWL5zlri/dQ66zHSqnnlvgzXMk7n1SaErgrAXD/Iuh82RZeK34+FpZniUjRUOEO
z9AUs7GNZaOLTE8o87LBtGN5UkcaZOoMMqRr6WORG+Z6XLw+puz6Zd9wD+QUEPDCIxbs+2Q0mzDD
Q5wcVrMeuof/1ImSzwZF1RI5NbN8xfVjwZR9YK/RXseNBaPr01cnlvgQC1z7APIZ2kP2hehlv8AY
1+2uNaHuCXCH3Ye0NBJ2OGbG0ZU1R7Uv0DSTZImnZ5UBn3NO5pOBrHUomG7ow7+cgMEoQU62w4Ca
YKXkiMshxfQR03hMMnQvKurCzLCWFTh7eHTM5R/fbf1Gy8E8DFjUIvediDIHvHk70ew2bwp2/3xV
tf0L/wjyxSEMMKbHX6bpocwkQ5LXq+qSanwm7P6vJwXUfREUyjdsWiObSz5l9hoBLhLCI2U7P2tW
yqZzc20fiTKxHaX+F5yzkpFcnSfHhmnGIBx9pVoARdeCBcGFws2gtIAaVnBe29G9AP9Ki0cBBw9p
IgBFwveX+V3Ys9rEODvqFVsCiipezVNuf1D8nd1Xe/n6+RnQLRHZ9M/LDJmFKB5hqBeGcrB+h9Zw
0P8+q8ml/j2wQ0qB/1KtrVwvffiSQRmGP5hvtLh3ti4OB/dLUuYqexq44wO1UiAs6cYf53BvMIqn
y6igZjjV7jDFoeRIDZ7/jBJhGZg3Icgo772xzQ44DpyuCP8/hIxRZyknA1X6h21g/+e0wf2Jx8cF
K10I5f9qNel6aZ5dqc7z5E7/4dvQ2Yw3I8LImLYtgCGcbhbeGx81d/ltCCwLdPOZpelxcMm7TYn3
H9nJ4DoKnwUyRUS2rXEERASOOqHiKQIR/vj6jcipr9jkbxrkdb1VBDV0hfkeF8exJ37NS8sAflgx
asFBRuH/vDaY42TgC/4os8tDrDMPhPszLobnz5Xk+obdrDF9AsmDr12mjVfLP5qer3VJrojlNqCu
xx0oV8fNK6uJ5AHm9YjjurjiFoyxV+/TngHNvJT9JQVM5A4DbrGR/4O6osAeKgH6QKrDscPKts3r
MAsXu7Ia1VXd1Pe4fvEJk53g4lU2eItZ4P+G2UFWP9FQzNxaElnYdsVjo//W7Cecns/K77UoUoHN
PpJdI1YXbkZqQEEaxnsR4kYyE3N9OoEMGsiiSWbp5SxFgE+EBiaRPFy40XyxjkZW7Gzmq1yZg5TY
k0UTA+1u1KnXLb+2OYTqnBgsO+JhykC5PfFdbs+YhylOwuNwljf1H3xJPLcKvRLi+VOyO73EsbDu
unxyEpE6yvQHkdwUP1Tg2qf20gNiZlNG0gRtGnbJprwXe3WGAC6vZcA7K1/SMCjsdDF9/SWDoiRM
K/Stiz9oY63C7bNwGsDk8WaJdUuzy2PBXcMO5mlHnRqW2azyfFbt71MCkqql6KwfOMoPoEYpyDk8
oRsrzN4l9m6FZk2dBiN58lJ6extDp9Tr8obrVckwy4v4wL1a59BxpwIXXj8aF7cmXa42sq4N56B/
DhQM7444wWH/xskPCrkQR0JgJA8Bz3OoYVX1A1T7zR/cqXrB857uQhhVWMxW6jND+fatSxnvsmMT
zIh2BLAZyvotC4Pp92Js1HuCPpE1FyjM2w/TTOezSjKdpuapAtCiY5audlZ6zeObL7dWd9ae1Gvu
Nl6iavhx7IgZ6mVCQWhIMqSk5KpGiY01bn9pk1DKXCb8FEfopw18bcw2Xet53N2tOg7kiiT5RjaG
u5eIhP/7uDuoeicNSU6Yt9tXKT0e2h0yKQAusn/Sy/8NiH6d0D6lSh6FUQHJsVws8T9zR3ZdTrHS
3+/JCCiiOPb+3/Sdg7drlIu26W2fIcHGIyVdhp8hc7wgx9bO1k3YtA9aoB9zQd8vBLI7pdYHpWnh
b6j6+CuPowlD7ilCV6gXimu0JTj3X06H2Gm6NJs9tU6NKl6Lq8T1Wg9zqN/0PRYePraJLDn2FuEG
NWJqrzqxl2OKbPPjUo2cS4DfpOSkLTWYhm2BI00ysYXHZCpgMQvxoL0zb46aIKM2GX4++gRDIT+R
ioPVEaBhKQPxpL2ezUB0deIkKZccRsb3GBgvxPp3JIF19c9FVjW680yGAvGeSxNRQVlh2VoQhroV
cjw10VJa2Zjxu0WJRwTnhsS7taAFwDZ5RVe2FgrKjvlqmIpVooLAXJKPl8+KCtwbjRrzAtbTeeu/
FCr61IzuK3Ui2WpXmFBW9ghTDMAD2CewZwWG354XBv2HRJvB3NkzpCxmRLjVfRMXqPLIfchQpEtj
nFyxgdUGIRrI5SC7eN0HKBDyHgQBBUYescTcGtZ3CISbMru7rgK8wN0yb6WjtAAiAXAj/rHyTikU
jGTao59kz3xt0NMhpluLFMKFucT/xocrOvyLHxu+KxmU/HGSkOsnLKMQRFZ1fOFAKWFHURweGOIH
/WcLMX49F8VH3pjPi+n3IMQB9Qveq8o3hqTwOZZCr3aPntzj6CPIdHrSGYmfFShWHVaNHf1vF34n
YKQmgTGk7DvvXfta/NtijFWxySO4Ivk0Z/Doz0/z3YVPjrUui46FwqRtVJ3EbevaOzdMWhgyd2YQ
SAh7Cw+xj1Nysm7c/d3Ccr/5CD0GObwebNhPOEiQwYyFz+VAISEf2Ep0JjMw9rROT5XtO8V1YK7m
gVCgKPm+OM09rxBbEMA2kmx2n1kBT8HEU5D9PVCbSLQZ8+jFIFzbyE+gMNHptDnI3P/VATRPel0F
wJOZkTBDDS7+AUx0I4oOpJfZxP2yvsuY9sVC0a7TgNiARRO2hgejZtcCQ0kKETT7TWF1AvaWqs3J
mfgGawEYxIdndLtfor2920DZIY873Up949MdsNSex2SvtY+EN/8LD12r0miAQZO+r8eOkFO7xyxe
g2rVaV9UefnGLG5/GIh4h9lTlkqoAsyDwKOST2ka65EFdbIhvMrAvubWowDoo8lGXY0kgRH2RSLK
GqkQKbtnZlV944j0sQIM5Gqzr3RNHBLL+t6iwTaZqFGIZ9iuxws23+rVPLIvJ6ZWWhIs52kcMp5H
p5f+tXX/dRcCwP9FAgjsyKwd+2nL7qPWFWAXtseIsEIz/ve31OlG/M3M+lrgLaFgLy2+3XrzjNIf
1k0tJfoLkR96NzLIyELsZonX8D11zt4ATMc4nGwfRky5JlH7s9+2DFFnrKyKWU+SIhQkNy8heCob
n+Tgcf0gLo6RMMI6FpE11swba6OE9dlTcW44FWIalXkJAq5V3nyFFHAbwMmMnASyNGVBB5Hn4ro4
6SNpboZG+Sob6zKnygNRJRqALweSHc1GOl9cwnShloo1SS2t2uCXLBv66YSAFSroLCLamR+7WdeA
tXBF29YcTp9zHpnhr15Q1E4tTX3VWiftSjTSZt9pfEQt+XTKBOvBzf34RV6r1EQn1YRiAZ5M+7rU
3yLynEt0R96ACg8M9NdaadKLtRg8u8TN527KaGnfIg4QTE+/8wo9ETAheN5E0w0EFO2QldO/TKU1
xWObiD+qYBFPok+6tfKLrVKXwOliyy5wFSA/qkhGqVIDwDyVHGTKhg9idA7UjmX1oI+Qib6B/lxF
Pk1I43PxoudKlkg6PMioCsab7ZvFkFZGqGGb3FhHuYWNN5MvFPCuXAPQLdzj1thGfyAxNWyoPUNL
TQCAg86goNfxlKaQz2DUUyIjHtP4guZdmrT6uflJYwE47As9jAp/tlsxwnIFg1wkhh3cYvWB3lpO
7LNfYYwn5l1Ks65SZBOA6BwD/64H/Wh5eSPngqRi8J6zkpR97kz/hVXTSqfoWGI61C0XiEWm30F/
MfKj05gUESOy1tKnzI0qd/pjpk8bbzg0IHrStohZ/RYhQySA8y+NyOGU4RPyjFYXft71f2DzI8ZA
iX38mfPqlSRsubYyzGL+VNWPvsfxNVxh0dWz+lmfHVlMJJk0eeUUO1oEudR6VNgYSOMIRpRDcI8Y
vx4a32ouamJYBY1oH1MtWhMeufEl9oLpYPzb0klQ2+BkjXxta4sFocE7dwdKCfeESY2GdwpsDMzB
lZcjzNPZqyNngqgXA38eGdErdeSOOmP+Fv5QV9NJJpJEGK7Rh/wqhqpJwSCtV4cOQQ+L9vd8jkn/
HVRyoBcqh5IOTd7sXmZxOMclsSHegjFeRuUz0MAzQUULlu0aM0lKaiUdj/RQCvKQXY8Jc8DwKa/j
leJS8VHC3fzJDo74G+/piUMWTQZKcZMrBAXhfPXHYJV1GeG3gD1xoUMV0Z2VkSW6E/JbIGk6dvJj
BaUe2q8U/3cBYwvZWJcg7F1hxAE7SbWOlBdeJ0/sMrs4POxTdnSI3QQNI0206uhvSgpsNhKiVla8
IRVJAUCrKz0mnxCQpX/OM/zBa9BuEsPlJBePy3r/pPXtne5pGGn5BsM/1KXM4b/Eatr31+wQMbPm
yfvE0rUaDv8tGWNqQmR15m+sEEzQXZIbVd4ADf+nWatYCU3dsCeWIa6S5GxSShgEm7GwlGYXTonO
D+pYD91bmE+IZvJZ14ASVe6/tyFZFgxUfiFDCV4CySQ2hudJgWgNt39AxyJ+F1mGHFsQ4oKmYl67
wo9i0yQX9gIgGvOvbpUXtRghHhkJ9aN0UMzYv3ID7/qPG35EG3TYHnwvA34AsW0j5FxPnx57rUOq
LbS6v08wBlNQEf0aUMf5gJYKjtNfKK+HE1YVj6XJ8cJHuX+HHWzc5RHoxuXglvEpmU9mhimBvHlM
0WTwPVXSz9uNCCZU3ISHSPS2vzhx34F++/HsveiEOSkGTDN5bQs/OaoJvpOO9Crh/Dbn6F0i7gTI
PpX5y1FdaGxbrWscXVxB/5Dr01BO9OLMKhN0X67HNRI2ggZLaEpJxPxaDXAziCCqreN4D+YK8NwL
a3uWdVLoNMFAnE9kz9vn3xj2HNtPRsXrSAqBIt02Hk+W3lph5mefthD9qGt0kJVNGZNRpf0AQiEr
YVZluqbHxGRXpxPLyMiK/Fuk3ij6ODCTdgvvBdiCqDy6bu/nGZW7BzrWJqgAl8Y7VzUl+0Vz6ol0
HZ2SWdFSkEFnbD8JTzZfp0YbkSa+SAMpf50UREoMqa4a0zDv8/D8PZoEFubdD5OAjhPubeFtzvFD
trayALBW4igllQLOwigqqHAbP+ykN+1FEQavg+2/GbddScPETIrd2OFagvD/a55DooPccEpymDl8
kOx263JaZ6hDSMHpT5nE1faDl8vy2u8bzdFeHfR+UxsWJGtHMv9YbD2Sdk7PXGHp5ECrHvsWX3Kc
w+mxh6BhX4t0kQj4eYTS3VVRBVPARX09gOkmJtCTnobDJDx+F7damAtOla89TBXtJfR+DfBYjLzz
UzhWZCwuzyeSjZkHR/bRPq5y+yHYxFEJe85JQ7qSpuklsmgLEg1DMVlrPohAJBpbnelp7hsMygzB
nLdU5gnSBbBAN/mL1T4DxrGYVhDc6Ct5TQAa1wSeCHuiPUF9zXcXPUiaw63ieaGXaP0XKT5j9XI9
95JY+B6N+plWq4PLPjUlS5HhKWG/nLG/svfjUc16jxCCAHaa1rdLg5IdbU6o3MJwWyGUztZc9A2z
5HqM0B085wg251IQGrlRFJ6sd/wZOhrjTXXGI6IadSYvDnmLUZ0GyocpSItSsLeXR0t7VF9K8O/r
K56BEFPq6liZw1NWr+VCR+6vNNi51NK89jb7MJSoUHJDbdLIfbr7ZnmNMOnjqq6HpIohn+UA9HJA
afkSJao5GT+hFpR95PwaWYaqvtWLcqT1uSyhDGQAjtzpykGMIJk/fCYgELsUBszrwOHiqDad
`pragma protect end_protected
