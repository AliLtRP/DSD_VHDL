// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SxQ9b142YAasvZY70+fvQPuTpdA2DIfvfzYQUBvLs4FpTPb9myhMNA9iHJdRj2Uv
M1RffyQwUyC/RT0mQ6F3x9uiYU3W8MWXjCYm232MQg3EXBfkSCd2flfy3gZfQ8o1
3AuDTTBd7GiGWloku5561RcMJwvmwX/fK2PgYlkjzA0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 56240)
zjp3yj2ZSvHcVW7/KMP/87DdRDRbtuiLWo7Y3P+BKgEokYmwiOYuTxLVuvPWizNL
fiu7Pf4NLHj220B7FGfnkCEIZxtzej1jq+V4qVwlmfum1nUJWJQMN7bA+91c02K2
Ox409DzSqrZkMcBSyxmxbsdbY7jkgUxsjIjPHkRN0MpRBEH+0B+4l48yL3idLazQ
tlVKOS1hpkntv3IxucO9AricaNNVqsSFZW5VaEo1wHT8oXo6M/8HYebI7pvqNpoY
NPZPKEmVOC/iItBglxjm61kXFEYl8Qf/vBcSYKX7nMNqAaICdgZuHafC50iyuZdx
bKySWfRgmbPT7l2Zse/dMGjmeCNNBO4+vYLRzMzJtZR2p8Ew11CDvoTxQMpM2BuI
RMdf5Nxgl3OkDfTiI2+2elsFbXkBonx3voPIFL6r0NftP+7QiYch1rTMH9k8LW0M
2yqZ0YusObqOPYeWnES8tBvGRnud917LgRWhjDbjdp/V7vr6kxIZs+Hx3gBc3yCj
EHF7bNxgTRk4coaYbUE1ZNDeIWgpkm9mKYQNo8cTEIYO3jFEEd3lWEZiHl9SerKW
UnYXYngnuEpdPcTsqsjgqioJXI7lopsSfVlUJSPItKCLRg4GboHQb0bKfx0ncBDK
Exgp8qqyy8uT5Olp7PU8X6dCHZIqBAC6TjySCYkZ+xm4yyuw+jpGPJ0NJvdKTLOe
VzXRLWY0kaBQkYuTHdX39sb8k8gn8HQnN46AyeIHAge29kEyliz/32MHUMVjCfLa
R8zmul9ZDIAT5burxrZLJbZt9LX9KHt+CJghj2p1gX0MuOkHp+nGZqNEEtxkFaC+
+wVvkP1f8wqzsajD1WNYKMAIfnQATFmAP1Ur5rprDk61KQksEcybYhE/4+1OrWn+
1yQEC/Aq6CVTVqBEnuul/EDKbtwcEIOnSHSsc4PmapkgdVChtzf8XZXCDmL1ginD
W8+yZMSdwtF8ZdZjAxLAHVrlnNdA3mv0w0zIIIEujaxQ5A/jIj4WL2q2no6Ss9lQ
R/W5IlPqqtPdnN3Eu/IFb7Hn02L7XCTfUnHuGFxtWsNrxqTqv+2Q99eSGjsMuqrk
XMat55wihBJnWrBiPrV8QOSkjikundNlAQH8po5olbYdfdFzgHBKB854Qea2IncV
0FpegB9CB0AkkLcLw/fuPokTXMiZ0a9Qkvegfvda8TT4TtkBHf/QVkIP33l4AQM+
35hBdqqnLQNNdrapX7aTtrVKLbMSXkJwG/QQygq8wmLfrud+e6y/TmJSVTmZL8wp
Q8a7SLb7WVwGxET+kHj0dv2MhO66AU+MRnavetpF+7TdiQgSlNWwy++T/1bgEWF+
sjr+0Fpb8HR88+oK6FtVfjKDAS/AAnc7IjbmJ+tdRei6AhAvJS8uT3J5REriWqZG
0N/gLzfa7iO9A4JfGSOYjpJ2wltNul13Xlc3WtXc9bphdbzVe3AOjDRovAkWJlyL
S/BQEoq/FRzK5QCMfJoXd1ezooJY1P6ghWo8Zs+iFYuoD4IKf/YeI9qzsz7QAN8e
ADIPad27EBjy6Z7Vqz79J5Q4gRlUeY+nB/b4CvRHiBgARGTxUHI5AN/IjwYCccD/
aUve79DjZoeNl2oo5HBmi28AaoZZfGNOeVh/mvo0VBJjjIoZxDhv6f+RScaCuvLc
5sOzIHZaNKTdeWukW794dz9pr7GXAkBOHlv+kYQBCxLTQsVTfSYdt1lb2s/QEH5a
S7MyDLbtAX3UY2Iba1AFlRBxkr2MMTRBJmiTHGhjy8KPkaB4Gx0WqXYYmmxOZiq9
p1FEvu3dK4Y7LXNh75SRDqG9YjMwWHjzG0EWT6OPRcN7QdnwLveJa5sKDngznad+
sSjDkdMEiosUZrrrVC/UMA3QCZGFm3b6Feo8+6WiwbULJ8pQwNjQtw0DJ98/kwsA
9GkLrtAuqKHK2/x+1cB9f+Od2pmix4mdo03xtcO4eMZBkC17/jV/o1uOn/XNTbQ1
qNm2+1SbEuI82d7aPKnR9leRRB1hoSUn1+CGZmRoFxxzMm/w79n2qWvp7PRYBJsh
BbrrYh8IpZUcgQWOHVcUArzgfLY12OOvZ3tV4/l9HDnTAkk3rV36Ob3u+k90UcpQ
zv0fHkTb+3V/gB4Je2sjnMrJ/UkEHfARz7+VTFCAXAY/ThmkH7bxXYFYYVKNjdXB
wHCNXKHKxQl2wOUEnOGIfn91lLNDeteiKT6HzUaZ4+kHejQ/nnVvD3H+Fw0390Vh
dW6ytoURc0EQVc8OxcDnOFDdmnY5aY1v+nXruSiS8JrCwCUFeS3Mi3+83Ni2m0KM
UvGcbxgUhlEaEipZoo9AT6X6VYvk/RN6z4Lv1XcrrIsB0Y4Z3WxQgxbOjMiyqA5x
xEIjIPCHNe8T6YUwXXJS60ZJ0WSx1RsvybgFToYYY1FG/wFcD5vMWQy5VEDEY742
qgosYil0x8sbgj2ewqvh8SyjFLAPo+6/pArowmEgM45O0FNAw33fCPr5yAAlzk0h
uEAdfQ5C7s48ySzNZb+/QKUzUQ1NJ1I0cRAZrQuLA3CEWj4gnYK+RQbCNzhcZlze
pevy3kH+BbwrhXRDYgXyh+vvGgpXe8/0ysa8oDmqK73Fh1aMaCdehaP/27pbqU6n
2Jd198O2YBqotoklJgf+T3l2cV4tNHAYhdO5XAtR3OGuTSdemupiO+zkxl6BVWMQ
mkuWtNU8/nvNIvovKpWasAQgGhMFduIfU+/4Wal7AAX21FsWQ6s0WLzhErWV12do
kv9WPT2mIU2dy1KCKvCXZPUDPIXQIckxq8G/Fkv9h4/uHS4L4WJgw0H1K7NCSzpp
hVjchjulJ/HceS2d95ZI9URrY6PjmX+g7DF7QcseysnWLjpt/di/2zKY7X7fOvVm
KvYF66DGLbjpmhbyhkCeWB20+hOKbxOii+llhJs72rZS4P1fskam5QzqKVi/AXvB
VFefCiTCN91pGBzahImjUBd/5LYU7o1rgXWbKBaojRFNuOkoCGF/bWaZkjqHEq9u
q63BPi0wISKbLHD9XsUY3F5K8K4QEiRGpZ32/obPZexFoI+XZuwX1W9jKU4BDPd7
V973aaaTzXpdtOhoYKonoLLW7zLT88f1N4G/PWRf7aFCdd1ROHGq69AUvWOMxNxk
3rQo/UykQnDeM2M/I/DyY/J9JELXz3WQf9Axe51DtqXNQicpKZQkgheE4uoI0Cd0
Ha7vcybb4/zbQriDDbFbrUZmlqz4wBUl1AtT7ttRi2daUHFfvBXIznj7fbr5UZKj
3xfZlHI8f1MPa6HPem1GV26j2uh5x0Tq8r0q3/Ru1bFix+Q+cmFRU2Jp2mjUcakM
vTMqnNUdVCgAe66NMdtSsTK4RpbKoEUEsH/WNrD4TvU5vm2q9/mm7MVjBFxYeCLt
R959XxFTwPMnzxik1FFsWGZOX9Su+Ki73F1arJFESEoVX2/HPrukW53k2ofeKs2H
xrmzC+zcjVzBijMEv35mrYJE9n19KYiNCNg8YNWKHodmxc7FT/H0f6tsUWACHN1S
qyC305+gPGsMQl/cmROva1G96AfIz+HAOPLa/HkAB6v+SZfoH1UQLniAm6M8loaj
7dTesl4i1IP0kpzToTu7/kF75Ts0EM5l+cYfcvo7CW9tsLnBbZ5Og2SxtL7o7gfX
8jMTeyq7WQfEI/jxItJlG0PxgRfE46NOZOJ04R7UZ+i3kHHjmcPImrLtaKBkjddQ
L9LppgPvDq7afZVfTamHoyuPrh7u5jUyqW3l/z22HsMIAnUXIr87LeprYVREJXCb
eqWrZQkPZ1tjASBZPZcmB+/sIeiodcwlzPxWZxaDt75XqyT7HZxCzHd9kD9DklTg
ajUYUgR2Ho2KCr2Ob0JZp5OAWI4yLIpOYtssyMcq8sxMSLv5QXkKyT0rJy9CvN8G
LoPYY85TxtIshmqkRs1uaheYhmci3jwBLEd6dT6HDhZW3FNU/gCqWowDr0qaDtNf
D6gGiWTFg6W3LVJT/1vfiPkXBQToz48LWGpTKSLEaZ3XchajmGiRA0TdrmjG1f1Z
rfS7dHO6GYBaO8enQGRz2GSIfgtTMz4wVKlY/l5dr+zSAiA5s0hoCboGyfP4l9UF
HFZcts+AsjCLnXx/lLkJA8ERwL6Dr/EzpTsZHZMqO5A/Zridgsoi80j4I6Dh0e80
mji2af8wW2w955ikRAIl5yN/xd5QmnTGHeKNGariB+ePEJ7d6VNMi8rjSfi7LKyU
4pg5brbxcRbgmtKgW65wPeTJq7WqAYkpScq5w71opR/ibEXbabjkwUlFamIiSjMu
+3nOA61sVj5aBIjKnWs3V5kfYY5Cn+yfW+ue9Sh0Qg8iQaOExumuQKePYiyG4aK2
CltSMLQIdj6UFoVqWzQyr7D+Gk+GpHDzyQMnYpYSVfZKjDMY2OP0qGL7rpNh3PFk
3ndzVm5G4YITJ2Rf3Q8HjDqUI8JUvx7zxRrx55J+1Ts6tMWePuMfaSiWOik+X5HQ
qVfSSS6aCGV1p7PLbSHSG5RmIathdii1XNRbO0V4kVavBLpqWX5PyrKTj8B6K2Vp
5S4+kGs/d4GavxFaT3jKDf4NkNPa2pY0s+wKhz2QrH+JLvlWMQ0jELHxSA8mWT6j
djvYtzvzvtTfY37nmH6u98VAWmjravww5t84JzbJmpedEa94BrORbo+/2t+is769
X8BBCKVKq02nw/fQcR462OoYf6AU5RunfyOc2EwAZcS0umUdvCXTuMNRRwcnyJUq
72pyXKQ/pTfhCrRQX23L/Ye7s+klrY5Hy8PsVAxBUU4eEFAVwambN+QDrozkWDy/
8Ma22i1eIdHawAGjPZvZmuO0VDx6hRmYskMqee8qJO3q1AD1HiAecIkMbdseefbC
QSUGlhSjqgHPIdbcQIBeaLScso/OLjrsEjyOIdg+ITU9zC3dWShZksE0wNlOwGg8
zpwcyuKA4EIh0e/JPejEvC4v8DVK1kRo9NK3rxqxfYFj0xxv0vhzev6Oe1EGjkGo
OxPcxBAEyBRrvgNnYj2pmat+BUloX3Tfo+/ZiqMRISGKhQA5RCa20QQTGhbT/Eb0
u6V5//nwebz7lOiWvM60xsp0F10m9U0UBJeRZrE7BXZEphss6uQWb8VtRBdCYYnX
M/X1xyv898rfbPPdsIlGa09Gb3/aCsGt1QDvy7Lw85Ofbzoz+I6L3nwU1gNRXZOI
5zQi5SAzvqqyFJvUjZLeryhbxspLw+uNAw1Gxn5FZcBRe1G8avjR3J5X0m7Cc3HJ
Vgq/kiOAueVRQdAiHz/5nnRDiiBecQO4f3IIEXbrGo752tBTQA098jszlVvE2YXQ
2n4TaHKsmiFeGjuL67yEsLXC3L4as2JQi6XjBMGzyQfZslBgo+TZI3TrKzA0sjBf
sVetRX9X+schnaKtzGY+QkfAijuf/S28dQxX4tOHrhcItNgHm5AZPolFc7Eh0veL
fzz12WgxV2fsMxZR9tC5VU2ERjxylnhrIR54CLycb/4MjkZPhJYb+QRkWY0aCEIS
RFTndulYiseSbF/lfdKGALvKOCHaIFSRGuZD3EY8CODHguapWTZqEU6T3hPg1MO2
zQ7frytXgyPLEpOIDsAh2ZR2bK5/YGC8l6S5aKtX+jE1AI3QXmbCJrzfQi+t4+5j
Y8cwf0W2P/JgiK5fv1HAlThsAtxt1Xz3T590ZiDEwgGFMLAC38SB+ukHETyB/rJ6
G3TYKAb+MOrXDPidvo81idtrktA6zRirBJXTXqSHB8Ox5zPvh3R+5QdNFQgSNSWf
GEhLAX6ubR8MzQZ2W4h1g5DDtoaE4c0i8qyjXfgiuKp2FUKgllEjy/9HxMOMs1hw
O0a1n+xCLPTx4m5Iuy6crBa7pi8gGoYwb3+ErH/sYRo2jnQ+xa5B0ABXZFr0FhwV
r14yLY0fID/RAzX3kTAfphwq6OftT4aKmOHQqQ0RVFXr1rY/04peq6yjWXCep3Eg
p62Akaqgg5znXbTIzdLC2FVrahct84fBm8XGOqsP0FmJ9IChaFjdQ1oo65kNF13X
n0hiLHOc08IVTK10LMv2lB/JF1axGde9YAwEzD/Ogf2AvV6plH5+tJhwSkYqkn3D
YbcXS5/WwTlCEZcbnlEpCBEhTgkcjMFPf631CShbp4CtK8QEHo3md5ho7qtZfCYe
CVFZNWu5U0vdSluiom/908ZMjssDPOkqfePUV/mRomHpzyb2qp/xpRNGd0PYYrNN
jGCGlStnJVl0NykhbT7Lwjf9I2SAsVxpzkbCubIncxi4orMoCjdfkdApKUSvLLob
rFFvhnJLn2OfhZzOTiMdVyVS2CqZoC6t2iW0LhCjRZsGgFbbzaqjiNsTLLcJfFi3
405Xz1SV59Ot+mCpKquvnCnMkXb6QYPjss5cI64gmnzmf1wT62xURAW1LxYHgH3S
+t2P7IeEpVy1iuai5jT1bOKXwWSOYozM/ylpH1sMuBImUFuqT0kyCXRCNgd568E+
JtaK9g79pucRr44brynhk1r1ISXp7YptgGcfGBozXFbSbDC908tfD5ECyR9GUqHi
uhr9g76It6uynFfazgiW1JVEnpnHUPQRufjPhwK7wCn75OeL3oMcsudlCP4p9ITi
zkaKxQZc4hl6AY6nZEOYpSu4alea/WtA6byUTNpKMg+9ByW/Xy+XFC1vUCLBJ7pE
RFm/TfiR0q9C8oawxsUdkjcbO9dFx1/YydtP1qhaOaG1RrOwuU+IZ0e1tJzWwjHU
9455EbZ7XxfhYXqTvGmSretFmMGpkJDWnCZ6uXJD01S2FdWQ76RuLHwiFADZIfKL
p3+wmbephoXqsVCgLIZ92mHw6Olhv68SLLzQThTZDwRcB3KJkAKXlEusfg26zHH9
2hj/qtPGjQ3QZ4McnWMHOa2PbZRSxg0de0uaC2HF7NWh4Dwg/xqV0LHU5b1pCJiF
/DFiJquAsXJ6pcABq6wufYkCF8n8jxEuXy/I80oF2DIhoE+di4jRx2+s+yZZd68z
7S6bLz2qkWQkqGa/0TEWtejSw6YBlp/T/WD4vK6Yg5Fz7HDyoPvzn6/qM5q+nf7z
I4coUTSFa+NhFCnn3UCEGze+qytt3nqOUBmvQ7GjLVCOZNRtY7vd86TUasBKopzr
p/RLOJWXQozsiUnuqRRFILe8ORs4cJ3kk9mgfPUG+Txs/zRpQz4sAWPD9p6dZjMo
chcnV1GENkFHsSlHfAtziG5tnjtCIAOeKx3aPjNB67USmNpb1QL/UOJ5Z+dNvirT
qJJlzdy0WX6FqulPQXRtvXA4gihqCmFg/gd7n6sjoRcm3gAqNQBhPE0DhVMiu3YH
7AM71sWNtKQcZ9qb3cbW+2oC8JfzyDbw8tUafEk/nUnFHTBoFTHQ2gCqOX/NDK0I
dPz6iPPLJImCwQx+mQ/REh/jwVyHH2sUzGNc0XZUu53cAyihIrrNHRnXa8OnyxZE
B+4yvZIe1koeRMv4dEt/i6fpKeLdX6zsaNmbq4KHfZGLtKsgyjgb3Hl9JMNVinQH
+7zZhKRXIyua1S8Sdv4TAkTOmP96hue8Bn1JUXsk8r/R9xkBek0CFlTMb9cQYoCp
yclKSPpDzlw3QGeDC+SQSo718cekfn8kMatz3GcGNINX7vgJSl7BSxeE+tBomg6+
olkEMGYDwLsHQcCVBrA8y6oYG6Mk1I2WBBxw4Qm7GovYGfowGkJeo5h4AsCDsW4u
Gh12y2Xtx3xdVQH+u8CPJl2IBFFSnyfCaiKW4KruJnVQkBVB1tLZbwkJLyhnWuTC
WnxPw9MH2i+mBnsO28NRYjkRcRxet//9OfAh8CaG47tEaa+fpCrlCFddJ5+ZJjnp
s38ibM602JATUr8I77GNhANvMtKxS2xBlahzvZsdyvYxkQmYcCCA3SmRmila/qpZ
dkkVL3QLKo1nWY4gawTYGFGbv4tSBYgl1aaElAaAK5gvjHVqsBUhHtdT1d7YLAS5
B38P4slaEoodfZsHkZUsZvXPoce9mCEJLfLtfZNk/pPaHmWuBR7KQ1dhyD6haPOX
1/rMeqpK9zrH79HTJVVhWzJe2FgHEgMoMMlAyZJZxk4RaJ5p09/MR3a5WRlQPykK
lSWXppoUbCy1Ltq4f8afCfffif7ipSGWcB0hohVdXPJCUb+pL37buOrgPCOA9iVI
hljrKM2BYXEO1nsx14BOay1mTUPSYXpaVQwiMLRzZTWa0FooDio02ZIRMHSShN9E
DQVJnwAlxAgUzGLhCllS8o6JpEqzYEeJwR9q4Y4N8RGVPmbC5OCnCkpE12arZAJN
Dn0kjREGifD9M3HpcEL2ZbI4Pw224yoCYv0Bl6z2Jl4j0nSm9pCB1hlblZzVV6oW
K4mrH+y1rBryoM0k93Ru0IhMPDfC1QVA8U4vVN0y5oyQnxEYo/3KgsmFb7kdyVij
4FgpDznYUs/8YiJkmFdNHuRp6laQwenBui7QTt7iAc5msbEo4GKZkVLTNlBF1yUo
CajWpIxe5c9BC40SqZQjlPd5pL5JtcNhM0r4JyGvENB+9D49DLNNGEaFfB3eSxiv
cf1gsnKvoXcNKeuVXYpnXDC0RT2bcY6iWceufW17EomhLndoDjd8z3AIwr30P9a0
oNNehHb5XqMebGpTcD3gwIzsWF3Ow+5a2jU6xe3Ob0qVISHUiCXagGcg+6CCGA2Q
gL65NZQumsOryXkEieGrTML0f4MNIXhYA/yLk6x6fmQDjjGQxgeuSr0cUUeSrf52
nfMjYy1F9XNkmpZtuM7nI28qpbh+eTWfJJTnwK+ZFfVFRumrVyNlpgw7nyIyg1AX
ExnASlKo/3ZuJnxBJvEtNfjICWIj6xvjTvgMt0ZmNa8qskkWdu5Tlrj5b2b7Olsn
fLF7CewpbxUdqxjaf9Nk9ApLu4G/o9m5rFB/MOqLHnN67c87PZUbJRO4DXAvOht5
pvp5gmVYO/nPWC0GbuC72Vot2Px7ujIqW1MyLRw7pTmXPWTNU6yglnpx8pv8qb92
/7polia9K8qQj3Yr9jor94cLWZDBjLu6vkUzX2zHTgo9K1hMOedbwP5niieu3+an
OuHuTzFeJiHG2D4WV67A2wAwXfh1bBLIsoqaj9aztla2pJ4ZC/3VH7lVYXTORnX5
MZ7oDNJm7x+iVlzEZpRXbTdUc8e/2AZrAYVBQvWOvEjKCOsUgJfs3aGx4Dfr+fPW
RxKKpualpv+aYRyrths+u+ip+6ZFUPM01iovScESiMk2mvia7RCU55vhrwFItHgy
y2XJCHAs2pM6r87SGOSnZNvupWkWBZc8Tnwvob/9/CLz7hjRz0gzOzpctZKcxLKB
voChWKq88cZGcAMTFTK0/mjDKyZvFR/OzpVKeYJfG/8QX24DdRX6sAqUFayf4nBb
tjW6nT/36Ft4dVa9zOhOqUGZ2i0Fyy4ODNweMW5u2DT7LtBUiXj80sIKoFhTzKuy
hXhq5AW4o7+vPvCGrVvY5rSVqSNfzCves17Z2uSuVaKrGxkJWlnYVNxE5TnM5Hpp
DF5ksdfdt77iKwm/e+Par7Zr/5ASWBva24z+RsUph/3U2Yz3vHVOszFyXIg4lMRl
6PYX0/D3l9CDWfEe4oUJLGtvcXu4qVeDAEMbm43PjiMIcf+4pUwaYKgQFbBwoTEU
Rucrm7FIg7UfjE6qxj30xE4XrDcQ719ZjNNiX6BQPs8U1vUcmPz3gEUhqJBrXdLd
nazdO9ghvHM1o591xFru4z5rmBrSrjN09v7e1tZl2U5lxDgD2OFEqG71dZrCEKmJ
nRFjkgxTLkg+dK+2Na/M7ZCagoRlmD1PxMKYwbuiKA+RGIqvli86au8vz+LU4067
nCd+Yrami+79m2GxP0kE9WuFvt6ctrYps3zpa1sWytcHxxcrETAWf94sK8dC86gP
i/EqY0PArP0O3jIBQZ5WNwIFljhq2WnP38UNvwF+sPTXKUidGJVyHVEESMSThySC
vtACQzwVwD8ibOWXFsF4PldoW8qOGWDjtJqH2SuzzvnRLi/wZrzTtjgeD2WR8mtB
6WUmud9ijN5hAa3PSwAAVF3S1w0HWu7RgUSItSEaUoSfsCk6aViD461uOaQ7q4iD
UsEzxIBbpec4cMwC7TbQ7sV+sbBqkkJm5Xg78OBrQjq1eu84+cWBx8WTd97R5Ttx
q0twIkqUr1b+otBvedVuHw36On5Mk9r2uuwScwdEJkev9wdHb8NVcVNO4M+t/xQp
7ZUpVnLjfxsDxd/J+tTXNkcQeVmzopnDMoHJqinD4e8pT/YY8Eyu9ZeZ5oO6+gM0
cceeq/5IeuFZOM1r2nA8ACVvZJNox9lVAjhX681sHZNgXESv+HWh1kKzOzV0z4Om
sB8TBoMhfmKFYKKM/1fL6/ZloERLNIo+6GDDJOjShzHbQp+VQES7sUCmaeSYG15G
myJJqWpiCCyWCgRQT/yCHAzH83EeO5lTwNfcpyq6kLbd++ymHDXvT8KXT0Zo4azF
4hWBfQ3pbUpxR/LHFrFqY0dQtjbvgGkY/PsAinC/Zp0dqRB6HdjWSu3FBVK4AFQU
Q72o4UbOnyxNxqTyJ035A+lfr9PNRBUbazwj5GgKqWxDUlQGcyukNEp71x+pdoXn
v0cfbR1GA64mSxR3Yo7qLuvGqNL1f2h/B6jwkfehewLEavDPUDAzRSPouNpBmf14
rLjW3yyG41VqlptZEPTsBVM8zboe/Lnd6Vk+Te7IRXD7JBWXhBiAvLwPRqpRlu3Q
Wcyly9tdiiZ1Y05Nc6ON/1nd7eYJ5ZWnsjbfKduNhaVNJQKRaRKvs93hraXWP0Qa
Ah7JJS3K8sSaw54LQfY8DuYPDaUlRqBcu4DWwQXG7XdOyHdVh6EpxJlgUR1mEkN/
lx0MnXHFDH06lw7oENZS7nFR4yML1P9rjx/o7YIcJH/5uIb7jTLuWdSUopfzcZi9
34vbNXImAsUeWh4h4F6N0axRR6Do72O+PKL2WkJF2JPPPcdb6FPTxeHziUZRNI3A
5OI66QkDpafku7yozqSUcbDJ9UHoivvOtUTCXCmP4TVQlU1/g1WfyT9NLIYFvvG9
3rjhQVIRedPGjUdFniZqD2gWSnPUpZHEYxDV+smUFhiqj4rU+CkDD7b95ZCrLyBt
T4nk1wBM9F/KUlkl8rZNsUNlMhNCoy1h2aKjAZR3+Y3FSy+3lRnE108UYguUiFy4
jDAcyZ5UnyAFik+qzrU+Qe7PqPBiltLiYxfFzyxlSFj87phh735/yWGyHVlphdSw
Nv9MPDGXm9f6tXtQlHXxlW7Mf8X0/W4uoIB8fT6ZPZKg/Nuv+J4oMWOIxVCezgW2
xC9JTLxwuwtIgpwMvg+FqFcKIAB3wLQfdXGC9/evfwR0/LVvo8Ao+GxP0DtWYcDo
1DdAxxkKSYi4II9wWzCVNYRVb3PUF8Xc5RpQttBnSvsoK+s+sZ7r6fLLt8mP3v2I
fOFshwUJTV8IKD9UxSkoWORwfMPnM4T7YHn69Z6Dz3ugFNgHWFRBXDsIoa+pfJbB
E++y9haJxRXO79jGV9prYEuVwu+UeP1hxyphpAr9VhNBltDj3CvqMjna8iIamB+T
QRPbB/uJ82+sL/qPm90s7CT6GA4LMJzh19Cu1miyUdipY4GknVkv8D6LOJyc7uce
uo/oR1hhyS+LQy1ExsD0mGZkv0cPekTSqne24a8QryfIFQNC7KOagDqiZFJaljoK
zgPmnlOcyRdaxx+eAtP+BJFQ7UtTMi1F1/58GQPq1BRk24sZV8qj4aSlOzIG8siT
EIxiLBri20V3YgzQyMAnsjt27aQka3WQQKGMYYKJDPlXnJ7BSOy/K7j2j7JNr6H5
5OBL3+NaUaDraYRaVJAYYEuwg/b2kwDpAVPheFsvU70+IiGvT4KeqW4yfQkg4lmH
muahRzFnq8U4vnp3pbMVEwMx8rXyHYKd7EfMpkMVdrvMjiqE3PNt4/F7KmKP7etj
eO6/r055kuPAmphZIBfj0VpyuWOQPVeBLvSI9GARsTHrFKctLr34c+04AfnbsgKA
z02IdokIRmSaMzPj46zu5ZhT1W2thUEYHozLBhS2TketHwbPNVcAw2WMfacEbFi/
1tJfm1axyJIq3cX3Brve8wmXg1YCt5W6Vk/RBVFKBlpzZ3JidF+aXuuc5J0o4aND
owZVWH1yOkeTYwflxEggPedKI7b3B2vJMq8YdPHNzN9L43lq1KmZhqHp/hoEWZNy
iU0RIZ2QSTPmGrf2t3PWG3dVtk4FO3JmVSLL/5NOkwE9psZzDMNQ+dRtAuo24/+l
EL+8DJcyYeLdOl0alqV7Iggiw8A8YRTn96ph3Rf/1DxMUAexiAwC3nVH4kaXavbw
tjjxYOStJE1aDvywqLDjZP6s+hsasICo9lhxBuWqTFu9eWqkems/tn2zW5sn6HNx
NXjgkC1cH2Ow24BLMerbgyzeCeyzBlKYm/nLaASM0llvY6vslr+6iNJ4wrAm6pVU
kbAItpa4/E2lXCtv9ci8oXyFQTHiXafgLrY1k2aX21MkOCsQecFhLydlafot5WLb
eadXi9R3wtvFRUr+lf+8uxdppntWMqzcQ5/dWtxWxexodVJpqCb/kQoHvd7fw7hH
PEiOchcS8K8jtOVg6wKcpTCSMNA6nMtajkDKa6nN7xEzz+Zpy8sSMP00cOE6ueQu
8yZxvNtYOkI40b3VxNyEh0agi4B3SVW+M/zQzEH6ACo1lxeyjD/6iNUfX/SMquj0
d9HcTi7Vo/cXihQoFasICih97WzPTl8OrrgtOLhMba2rFkC/RZD07tq46Bl8MlUX
a7hCF8oiVkQO3GBjll4gcV9dhPwqvdy9qeDrP4IqrEp7afjZNN1Ij3ZipXzabVft
7q0Sj42DuWxBurXzVx3FGt9D58pxcHgo1precTfXW6ccFZyjeOAbvI4OQpraXXyT
pZFJnwo7FC5xZf/OMBNkul0Cm97zQTdFmhXmhfWlZtvguF4pC9nymXWQfCM/dIAy
WErR3j4ufWD1vHH0RRhitmwUcRhgIueIIaX8YLl4Z8N0CTgqHt8tiwBIqgtDPnI3
bwwkZC6HxylsND9CQcVMr01VuCnOAeiorzkUbC8j95P3KlHXYBOdILsbnW41wcqT
lXhw2Pd3wvxiaoMNl9HoumUsuoLO9c6fLQBhn62Q83d1Lo6nm+gPXmkdHi1PJP9s
5yDpvEppn9fzg5VDKxuZx1YV3eUKw35gOFwNnOj1vbnPZ8m1l4W7hFOGvi768zGs
gxa5gqp9bNwiGN6Hn5zWQ7ArvWD82qEvn5gWQ4fZ7tX1vRQfr1EoQeTnGV7OI6Cn
pdl41oM3jphS12O8Qx7fE58dcI2jdkQWaMu9PD1e7f4+e2Kt5MnzYh/a8ZvIC3ME
y+RP33oYItABMk074jsF13acBD+on47YFBxSXXlIILeRa5slvJ1s1r/n3onKmd1S
9BbDVT9g5nDjM0WKAb6aVJyXZhHtkJJR0rY5+m+DwT+uhXWMvzCBd1ddL32rwRNo
7X/ItnCZstF5/wYuQaM9BM7+hmyoEpoh90ye/q16p6dtJEXC4l0sRkiXQmZsvxH3
F8eGAAmz6/s1ycgsAdFWVVTOq8sEayYQHoIZ8mRzxVQYXc/fQKkns6aSQoaKw2rS
W4BsnPFJG94Pt6UjfomaL2TSbjHDqkOF2keOVkKb1sLutviHb4ndp9pMEGMzzHz8
z08lzsVaSLn0SY0FSHp8zfchQHBXxMAYLH6w1PGZvxqjSBl/MDqkfAgOV58+oMiH
jxZ/I99q9I+YppyCXEnWJ38RKmFX1ts36lGpLhxnRNg6kRTgwDsEBMU/a2jB6UXC
CtLLHKX/C/VDvKXQaUrem45+NohPwQkls4wP5DNkTPMI/QUQWxkiqAolJo8TPw/G
UECTGCiY8p8meHHUehbDWFHJRaf0Qa1OwjBceZasSIFdSx5mxprE589QazERDpg6
Wg4Tbqv9bLX71IWX2lfyiPVUfEi5n+KxyXxGbVhRci5yGj3SbdgQPIs+X0xyE0ne
IPX5u/EcDDdJ8+HrOC85fgZqtYusqOvaf/n5q2qxVuyGtZcvxQuQH1dAh8qVnKcy
yzJPm+w83QE8HhxJoCfWIPm0OQ+XHLiYxY6OeRKxXrDlI6mMBS0bwLNdzRReIMR2
NLuEaQM3Kr6H5bDSdVzcMk3ci/w0JpRc0BeINWe7+VZz+q+daZNjAgDYm7KzHkYs
RmCZ/jvDkBBNy31O6edrGLNO6UVdGYSLTMOaCfpUqehLQ11W22rzwGS3P6EA+Ibf
FiD/e5A6t2WrfBAMGMYlct4/5GqfGx3CsRPq8ruYwzYGf+peE0v52npFjCH9zn/0
avYaGPkReMXxogijrhiex/Nqzqw+7Lrxhvc7xuLKSTPwU6KEbenCHfXPUsNBaFmK
g6OkaXffGZrCNo50EkDJRbYo6yHqpbgfzuxV2O7jJXwdgWri43r8z5H7PHe4IaLc
imM0fjV7NpYK5fyHauDRxnsSWE+WaPzQ6+pIo0fQe6+IS3qsAbW9ExuF+euWp2UD
hesXlB/syRf8nagEhA4nVqvyihCjP7bzEmjk/2qOE4RnFvNHQuTF09QdztDK6CpG
0rX8TLUoLflBJdrV0KBcqnbgkQGWoa8afaaENeJxvP7LAXil5yZ5Ya89xzGcpBwF
Pa9nzXbUOxBZEDVtT27mYovNx/LQwyuvDcqUvIf7qxAvWWqJx19+1Q5g8HoJeULq
O2gigCF3Q6+uTxsVrOEBIPCqZZDZHC2+TqlCrOrQWz9eiIXsieQ3WBzF+PBM1Mur
QcHrsqaqBR7gDQ+iKhPu38xgUtL1N87Q/2bS5i9ny8VLtdhjT/e4GUdWp17I0cmK
2VuelnTIp3Vqve+oCRLF6yAbgB9VYD/+LWCukQmYKMI5r2uknX3CKZ3hVFjgaqCi
FbUVxzG9xu5moIjhktCNULd8HoHcJodWntigQvE8Adv2Lgn45KOdze42EUhINsZM
V1uLZ2pA0KfrSDJolbsX9BjBCK0jiJWXUDeD9F0c35beUFaLMKAUI3KCjW1rBFrD
i4WmVh8Tz5hHacRkr5bX0x6cR8F0cOxNOl7pSqMeyfGJP9Gf1D0q/I1J+9XCdVoq
j2/8/4hiwPexf+SAmbrMRxbJ9kw71WsXaAe2VwPpwxiOXhiGLr1r4odP/bskP+Gq
gs9ugyQfKeVl1pKlHSTa/74e8KqDHsrP0ZpXmgTXbcNELuMv+2dx61mfDkr3iouA
Pj+LysaXXQbBt7uVK1CGKfMG1UbtrPmG3wdsuVAKyTN853bOHFHvH7ZfhFYzs13b
yO19AeD4490SXsgjyK99xyDVmVCdS4J/Opfk9WirDGGjNYEjcvfY0w4d0Vb2RFEt
ZK51c+cUEc/Vi6wRDInHlATUpm60rmdEndIj9e+8kE9Ybd/r7AOW9g0mJTwVXUSy
fEv+2jGBVxxNqiwa7C8td/FTZ5c18yAC/1c1bT+2PWStgeMQh7CM42Wj/ySAv0Im
xgK+ePEtQJs1YKMBqJfFE6wVxKslfDa+5UWAHGYyazh1sgOqblfT1IOsqptD1P0Z
BJdvjQUxUNnYspVbCPkjY0agCHOZsU7y0wsy/s91CzKyeSDkDroJu5jRGdmsXL4u
rfppy7SMi8g1+6h7MkksOzcZLAOhiSi817M3278TjdgFMSRFApp3CUxhdRRHxAfP
WCeEgK12m+E3G613twF3U+BsPSI6ftXwQmUK4C3FTS2USi1Xkqy9yEYrYpiJ5doV
iE9eggPCy1nQ4fFUN4IJJlEYj+syz6CBNSLaO3oVExwfxGCKhSQI18eSo6mGDpXu
38PDGpz1JH1H8zXri5x+6LXMfj7b/WIyJB2dyiiVSgnEV0NnILPIqfSGfMPg3Ygm
HxmbavOywfQDPojbwP9NsL+28rxDkz3OLXryzcItL1z7Uzag3H9e7d1pS6yU0OKu
R6sMFicC9ruzddqOVtZBUQgsp3UMNluh05x8v2U/pxVPjqk0Gym8kvJ4yaYZpnML
3IwSXmreedYqqj9cPW9hcjAmC00/ZzgfYnwLJWdw7ogHYepY8FvqP+XI9LTbowf+
h/pFThcp7CzmJY8xDnQc3TE6buSR18mqJLzph0qEyS67Q/03BMDc+ZK5pHvcpHlA
feT7Ow2tcO8t1zmlouWcdFM1uuif/dUQdMgGhKp6LxmCZh2UTCuo8b/ZBdb4NFWO
cCgsjfy8ZBik8VZU7622Ouf2dd/19mTXIIRz8QvT5/J+xQR51m52xCrhQSYjeXc1
feGiJFAySK7EtEBh1Z+d4RX5lkrORl0lWYYTg8qYyTww60/8b8CGRSjJNRJHGcLu
zRAYvNB/NC0jZ0bBs4ebAVi4HJVaAbC5Yr+t2ip35KKQTTBvJCuf2qFp81LhG787
pAIc6q/9zDu4tT+keJ9o7RjX/aCKEG6pqQfFMsAd52T67c7BAh4EV5I7amYMuawz
BBKdkXzpAkQJKfkN8f6vWjC1lBmTYSK0d9AHdJieMpoYhSfPlv0dSBn4VYRQIwB0
xUw9WbuAOCRZyWwnh2gXV0UywW5qIkke4VX0S53LuqtNvYZ9t7e77Py1wA7H2kio
3V5VuEQ3yxbUF4HFpxt69xcXCppx1aPgufMgW7OwdrU2w6sel96gouTqL2rDpYzg
IOePI9sJBXHjbyvukVuFFpi3hjl5ASfvRk7ThSjda0Makt5D9TKYSkwtXMPYoWJj
9cCp5YFdtvj7syqxWcjOegu+TDMkpJiivVRUnxgeQ3llwI5CKORUupHW/gwF7V7C
JT+thwqBuCNBCA76Jp1H1rAZhXRdpXH7W0dKZG/8Tupdq6WU9F8TRf6Toi1nenQj
/eBjO3FAni0Q6dvV304lZ1SwJyTbBa052yuu6Vo0kyt8qFgy2VIMVICTExXf4yNn
NJ2XUlpVKVC1U9Wfesm6zPbi2TeKOHXxYvEA0fGLbXo5a8rVK77e7CziYgs+qb3O
Uvjn260OvhYb/fv9DeLZU2iSj+JZ/lGLKXnJIysiadqb++5Oq3xNg2UvjaeOzIN4
5BUs9IXvb2L5Rcmnn5JAnnesZIx2aWaS6xM4Jbv1HqFRgwoXKT2/kdHG+qW2zSKA
deZ3Nj8LCs8vjY7u8xkYwdvF1oUBtjmlMtfvhhZOBUEWKPlkNL875yuhlR4HeZ2S
WNO9y4SSFo5HQW7z6sL3FbHWfAJQZFVhIBRPaXCJ8Uj/bL8hd8E7n1Q42Y443fsD
d1PhjBXGz1GYUVQy/r/2Zz99wty4tKoRKaPVIUy8M3tQ4xz/68ulNaAgtzu+35y0
6tDzenzv+UqcaCehnAiBfY2qysbyXZTvi/nEX0a6Htrm19+4x70zbknig0Zj5BSf
vifmb3fiP3jV3monZbE6axuHZwLJszkvK+u+i0OTEbSHO+O0EFCo7a2hSzahrLtT
B9UvenRa+vYm86TECB9952kHZWZ/wXfKCwJNC/3FxJTgTjPrppQ9I6XcbS8xkJHq
6XWM3ep/kKJn1JDVMw2N97QvM+MVWeGrfthx8vufjtgUlZ1sR52TVF3lh3ExcXte
rjbGy1savCZMHXJ3bSaUe1NXq4s87eNvnw1acvj48ACj9XJhbkAuvmLq845+cB+i
XaSfaEApuEnruN5LsNrZe6Mu6Au4ie5FaMtqYdH0ZicEO6jWXexQOn681QYcjUMx
W2Ib58l9sfSSpXUfYpYTJPTzpo9qSxd+YK9kaGb08y2zn5FFip7qb2Ug1zcELZlc
4C1xpFVqbzzPfUJ4qphMosKkJJYEIP81gfCyVqkn66i4UPjuy1U7Tyvki02wMrnF
8otDm9Mi7zNBriPUVY/tA0MdWbH7ljMo8liRgpdgpHfsufLma4nGv0Ox8gygU+uZ
+rX71ZHe+0gKay4o8XA9pw1pp+ogwBoXBzwSMzhVLyxKPsXTdeEk4UiJGsi05YqK
YnqfxPXwQOISrHNoIi0LjceAw15JFB9bDqDWq6OKyDV+iMTzGVX+NLBYmM9tyfMU
Jho4fc0yj3TG67c5KUzvgFP6PLMHlgPOEQw3Yj2LTufvF6Gg3TJOJb6m0SV2is/Y
bZpSmjyF4c7rFkvTpGo/zg6DFMRZ4iVURPPdvovxS2UlkazEhuUEPptjudafxmwh
MhHzfpu8jF0+f90cRzcwyVboOz0lJ1O3JDlDcu0sFApMGaaxMpnOe0CiY7Uxi8lc
da1yXBqveiuV1xA5Soo7Scu94m7AfUChjiSvcyiy2zHXQBwHN9RCT3/uBfx2bTfW
HIKe2nrnF67TYFbIxuIzwXUAXcvn+Mt7K+7bdFHAXAG1a9vjZYgBhCZqpLVrrUL+
izvymrEV6iU9EqKkKTVbPN1fDeA9G8w7tNizP3HROHqmG5GUq6En26pvWn/lpuGg
/h+m23AU+PaI+tOXfTGy7U0C815TGmQxEx9eH4ORrhTD0QvIlzTE7I3ukifVdgrj
EQ3NantV3uFe6Mw+PCs0L/fstaos8Eyrqq5oa5CUv6U2pNZ3nYK/FuaL5ya+WMwf
DQCwbzOVlD4SY9CwQN/xQ/e2z0/cU20KmTrCuXWdlHPJmeXtAMFtUU7fV1088uE4
sozqXwgk0QTazm0N6EpgUNgVN5H2JyP0WyEiuKUxAa5FftHKkGQ2uyQs/RmIef6t
kUcVQEfAeLhVk1bZToxUDKuONt2ACn3W0uLDHWkE3TgUjqcRjTv19iIhd7Lh1FXr
aJuhAMYPg2TtZn/a+DoAqVBzRkZom8uB+D8DssSAJrTrjOFlh/EldC4ldRm/xwTn
1P1xl04eUh230zM4UZ0MqD5tudGz8TeD0er8AfsGLboGy92HGjlWUBUX04XQi0aV
eRZArKljo1wTrdH9VSfnEOGraOrnDm0RLn49k/7VH35yKjMbOcK14FLwlIPshOLV
ZVJdR+fNXrSJzzzTYtIIMX7IdJAqQPbpUrVsN0mAZQkRwsFqwOspiRRhKKE8upY1
oOV1NdssMUvW5qbk/f1FISNLP+TujNk/DUAvIm/60kQk2sR9G+p8bwUP9FX1a3GA
QgowvFw/0PjiODjipiVOiysrURPua9fR3Cf64eKhSA27Rjrx2I3vSzNe/h3rVMlN
6XYWiB0Sx2ysp1JhDP8+O5gpFjMAaKitDt2n6tywDEqGoQEL9X5ogB+rsZUljDVK
NsS/ENQnRB2kpHUdrU2ER9k/c0IynajI4y7DvvupVcPGfwK0FVLWU9gD1gJn8jmI
NWlodJXU3qA6HLj7RZXnJ2MWHJe12AVP2QnbRFCOsA507gyirQvOy5XWyGydmCi0
tjdQyojH2rsFAkr6KWveD8xuwPnG0nJSk2QqASCd5pM8OaQUULOolrSB9qzw0Zly
HISzbSMU7nNKvQXr+RknaVFVoHBRXdWmY3ilQ/jCsdLJzPLhpH+hRUTQJUEIGc/K
N1jcyNegCF9M0qW0AUbSY6uRx7LAPwHMT+CC7QgCxtvuqTys75f5o7S6Ev+uHkRw
fCozGvP4szzX/pxbOJcsSVQ7KcACYKa9MRalVJOenQFgtLuZ8//1mN/t90hQzmnA
AfThtg6NTS3OvTJZMnxC1YbBTHhFyi82LPdS9vLGEoh29qA+YcaTh6TpK+AKa/4c
cASobtGT9Lly1Nbqn0WR4KINsIIezDGo5uFpVQaALctBBZTIaIu/4czB16/JIXBe
NB9oy3eSpTKYkGtMRvnzxsRyHS2ofEmhfLiDeV309pXn3WTGrHnfGIF3qBDRS3UH
HCcU19UQg5DmeQEniM1kpjGIoG13z2Aizn46Bt3Z7ExMC5yO8YI2RjnEiLMUTeqd
xh7nQ0mnLxMqQB44O22i17XI/DrISFckUD1xzWdlQxLCI0q9ggOcJulzNxizP3C3
eqYofF/1gJnkbEhkiXcuHHwLzcLeChddh2+mZ2I9FuL7GXHQekicSLHXLB5bQnFS
e54G/860UcjM639bpZBLu7i09PrCuH5B7zwJ8knuWIikwCsmZR1AJutov3mSU1P6
awfyYTDEpyI5hT+qZhYrx8PpZx3pOvlxeq/J2sYrkpnpEf5F4iUSlzLk0XLgNrGs
X8LGVaOPY/X752JOWhH7NMiuUgXo4j68ue8/QGp+Kl2AgngyL3WNawQfRMtC2634
ULte6fTeeUwT++MBIhCCC9HftTtoZko9b93MI7itm6VN/IAa5L518WXcVaOeLZCA
H86hwM3x5NANkDeTw240rQ5732KnRup7RHtsusXgcSJdsRmv74r5sc75TaMPlWW4
PQEH5y6y4HTnB9Ho42mtLF9SxrEDLP1UQv1o8OLEzVh6gJvUPzpKBd3+2ZdxV5Jd
1Ha8WI9ihaEsmp9OsLhtyWQG4IaXymjiyZlvBrxJNBfpTp9ft5b2u0zu1Gj1EN3R
GIPPH5E/hq4AtQSojvXWpOGT3zc9gG35SJiuOyCmKhze9VVBUK+aLBp32adgMCxL
XyQWHw3WhrzfTORsAsr7pfoMGx9ctwRbJL162ROsRt4MgGdEq4hw/KGVXIb4XKDK
ha/lQaJ68XVXUneuugVEhvjGX7DBhOB/2dBsxmsLdsr3QqShEwYS6yn2hXn5W1gk
TA1rajxds+IMmliCA/PyaLcoptJDroqzVxxb4gi3HbrM5D5BZctPG/EcqqXA9HlP
Z1AcxjTjoqy+0Wjcxw0haxGSXgieZjRJzAzuNCZtZ112rmUqzqwGsDy/9ucpvDoT
qjGkWUmL84nKmsrbThNMaeP/agnEMl821efJWl5oLAW+oqOMhtDaDN5VABQ7k6Qs
UvlRWBjV/DDXoxmn0wHwcsgQ95ho24IrFDROz2KxOvPIYAFuKvSFKbcRerJ67Flk
c2w6DpJslLzBxh5gJUUnG02EaBjLMSwRqFHOfwUH3QIrqRIbdDIg6kSgO7kdvV8q
oQSyjbuqGJpRkHY8youWIq0fmdzA5Kvl4kH6lOykC0MTeAiWIQFymsvRn1yQm2RC
vlccXcCO076a7MpDo4bxzVy0Zzvj2RauDifrdup7NIrDACchOTlS9ZH5hfGapKdZ
0ejnZ8GjLPdMeBuXBh+O2n+8v7Bjma1n17I4h7rkII4qmHWs0IEeTuR6TuRKN6LS
EvQ46lFU2x+46bkYsloyWHkX1cSfSBa/9FRLm9lEkhO4qH4BrtN1Mt3rHkKg5kbY
RhcHYRjjgf4cDyPC44NvTGzlHZiA5oNI3QFJjmm351kGJkOmD8ATuT/50CVq9mME
thLO07gghw4hWSI3PkAP3jEr7rWt3whDlP0NXaifgLUf3NXzip8Bv3ODuxMuBGLm
ipM/ok6/GqI5vV7zOET2DA7JXbpmAq2U7KGCoKOijapFydvoyfMvnR1cFAAocHEt
VggPaN2ZSrvRutvZGpQZSx2/v4IruskOTEMZi+NxLSt1CQ9+mkCrxkAh3wxPDgE+
/AuN9TUtsDWv6R/JJmOPBXhvGGU2gLamRbKoZdX8PdJlLk7tV+zQwyWCi8veZaFE
wQX6F5EAjLElNzHymt+Xhhl6Z+AcMVv+4D8qkO/XWWahMbTDhcQCHz8btwGbgqEK
7TMGDbLDScrNW4/LSbyP9ZSbgSpJ49QhOOLR1cvQWKj1BnLFtUfQqS2JGMKndRsU
jhDeOOvGw05LsxgA1hiVIa3aKuzIJ+YZCT7EHOrxePgtaDB2krMTMqYWJ5zvR32A
FwZlk7eSm4v+XWGx25apJNir06X30BxTF4m8OyDifmoig61sN3YNGbQzFjXOtUym
zzCc52W4g33PgXw5lbigQ1+DA36Z7csSGmOHReHnWzpoxWnovSKooT4Bn8W2o8Fx
dST33OTQp1Yjy1fJJwZE9GOQCmgy43y5uAE3iugNO/O2RfhqvCKKHehENJJRhcWR
JQYbOKCXQWpBK2jQ8uOp2FbIaRfoFUIj27jHP0gfjECsFJkRsYWIOfsPwGQLRn3E
7v6tNkra9Ivc3cvebPzyIvL/w2JbsfH588kkzZzDj2vsZXuP8As/JSUvA+KfSV/l
ZamFbZAsFC1WwGxU60lqvqAARXvwhcJhsdxQqHfn2YeX/R88hW9GLVXoSxZtgBQ/
c65QKJ3Qupm5enJsVsLfjdo9JI9wZuLQdrz3ddTXOT+GW120QR9svaJsB+nIN3UG
E4D76PAJJHFZff2+VHXVLi90NGgJWWW6yPw12dpECyk8+DNcAHDAaSUee0EsoAFU
rw/mOeJ6V3C+1AbWVCvp3KdVlKuuF+5ZgLbRQJamjXMCOlzvNUjAooje57Pq0YpR
gp1iE1puS0amRsJbxFkKtUAgJecH+uIoiWm0qDLQzlHJTx1DcOkKUx4fsV7dWRoX
/w0sTedExwXHQI8Nn46VIMVIsrB/pFc0jiC6qGvWqmt8SHtlTUdf/DrHUzrDb2bJ
TLVndV00EOmC6ysJdOv5I8F66hPvzqI1owbLWAZ/xciIFiKhWG/Jh3VIj38MzKjw
0KVksv8alPhxlRvCAlnXOXeBqZN/dGhcoinABt3b/DNgvg0VELCd1GcwABrAYCQr
c8u8dYoKal0Vzb+c0ujEjqgihbcOf5v+7CjTakjsRWlOiC44Y4x3cEJd00i9Qx6N
FKeltz9Xc6e/gOZG0gwmrBlq4X+besWGDP/RnUfxYOzeI51WCu/jVISd0DgGSInR
89MkpDWtYG2p6SdY0+JTuUVzZ6eAt0gMbMA+hb/x6jhyGnyMuo+HnTQ6cMyLEULc
rEj9XgV6w8DpX6yr4eVNJ82Oer76vwXd4CV8g7hEFCB50V576PQNXQpy0zy3t5gS
A4ZqFK7blB45oA1XN2PVp58/nSQCfKgzH96seQV4lXespjESFOotbrRAG3dlC7ST
DNfmf8Phq51iAUtutgKvvWWM4Pv13eQ5dO/pVaZkPYSUm9qyEMXDjd8N0KzZm9RE
/x15X+BYkpcTJvEvfXowU8Qu6YTWU54H344YMC/AfEuz9gbxDNPb31DL+C6O7fso
evAzq+4WC+kHoW0blehD323JpSNiL8fjIynfSSOeUEi8kPeQBIg/X6oidpG4HZa7
Sk7OdBgSpd/fnMp6PIMF4aveBem5WGDXOok64az7nwIWc3OBgyiHqG0P1H8lVPw0
ZsmXqllZJtZp8PkJqULZnOZJqmICQ4iBQLp7YqsQI8AVmLC1Awbg2vzhSC6ddNuG
nmH3GM49X5aieYDPTjZJRNmVcXOAdRIqY3Myp07j+j1r6QgFtSFFx8HX+dF4Q8yI
2aL+plFlcbQIdrnLyBCNmfx/jW7ZmLD2mzb7y0ANFwm63kVVsdEMqc2REOM8ubk3
MFs1epwQS/xidWw9rEvBstrO/3qB8hfIJM1+v7L5AVaXECmRgG65MiI0jafdhKkK
KCfVOF4Tc2QJz9h8JWcjwQhMYWZoE58r0+1RLyBsW2qI2ZayqFJe8O3cYE25KWqo
BdV5z71NlhP2T7VlpbIHqMwUVIC4sE0p52nilfdW6NcsSWTqWIJLNnkpbybMzezV
wQhCEoNRI/yS+hHaJEBtYqwZIiolIH+5IZXEh99SqabHb81h4f6wq3OBn1PVKozk
hzMpkeCrw5cKkFnruPr3XrPWWyG5sKhH9ODtOIMaeP/zgh3BD2pRsfcDJk7bA1Ym
rCR7jttGa+6g0hXa3YmsHjZgoWpe6xFwJH2EPH+JRgq/li6uARfI9jPX6hbPfW+7
QsAwu3/cc/aZttTe+FpPrj6nOyA3ddISTL+GMnqkMUPOSI7JySBsafUZlsJHJvJt
TVznFTrcbxbQpGA3VJa5paZFjX0EqZFV4ZNkGtUehyX9Rp7x7hEWP2GbF3DCgYXn
MW9zwY/lA7agKmp5ucDYBAl4rfeXdodmLt3ICFZ3w2w3SdFZO+mO8Qr893YzqFjx
e0Jl+G8vk+jO9lKjLno3F/n4ECd9BUsBBmFjdmhNHr/BZbmCpSxWY6AnTRwNZlC3
WxUB9rWAelo0zXbfFJWt1Jev3z5I976rLVBBkpL5pEzsnd+qTvSzlA8SpQwgGCxY
rotLI59pEh9ja1EUkI98qYCvjyMhug20Ix1Sxzd9PJxKJRRIWquTHHfmcX2DRHj4
+AQsARd2QatrcWVcL5aUS53U4UQ35K1/fSIVmfPcXUnHetxKm9YOAmJt5FkSuKCF
Cl6e8n81lkSBcQVnfd/2w+mIhG+xJgJuF2gANCO2J1SHhoBbCB6RZLCheK6XGazL
gN1yzOmpvWyhyDTLwI878LnGJei0a0b/smPzEh/2LsMqcDJhk9dHWbWFuGFYeWLJ
AntZPOZODdNkBu3oH9n9uVl4Mq/gOZI5005M6a2gp90ov/sHRT1yhB9U7iHrtqzy
IOeTM8qSAqNz/6GoZAJo195RRxU+lmc7JqB8a8KLVxzA3u9OMlpjI71ryvaCVz6+
vMDPFBVQIaobJG4aZkwwQrHrC7a0KJR3lfJEvxeX8Jj0yz5z0f4oV3SPsTsFkUD1
TSXF8LKlBm1wHWIaRE91VciYW/t5QF83JzxkCBedhZBNF6epGvruisYkQ+UmhjbC
gildgLtV9z/KlvgLpw2rFLCSbnI+S/sy9+Nff4y/YeQjSAuwIsUDw/+XExevkFr7
ePdTWDMkb4T52CDQvWaj1Nc5aSmOz/WhVJLCFpFVdPbqEeLpfO6hZYY+XQHyzGiY
hTTRu+fhEHQCmNPaMcTt+DUl7LURTakfehLeXwIqjC+99cWfNY17i2ERXBhPKC3S
/YeBJT+IKq9Bu4neSQIUza7wseLc/5zsLhj26/qmSVDc9tt09Ot5/+tezHb3h0Vu
MAogrydmisuihwLsCnzQ8Q9qhV3tFWktq15vQmwBf4hVDS38nGfiLHwoY+zWD8HG
khWESMdxKiX+z9XrpaqS+IjyrXU/exWCINe/WW2aqStOmrvU3EGjwRTqwTFL5vSN
kqY1aDqNfJHx8H6Ur+p38kmIOGvjFK/Kl8Qsgg+XCQxZ7Jhhq3TlAFj0543Eeit/
tLjVjjUepeZ/l0fEz8IEgVBw4DpZcKaLa1tuk8vZNi7xab4Mz7U70jINjs6aySgE
ZEzCOUbFLxX/ZwGkJyRlSRooTlEu6MLt1sjw7zlnaurQ5gsPk2VVVSNhaxiqttTv
IzSYeQm/GsEfVdS7PCLQdTpvQR8oN+ArKB5pMcUQ49em/o5yHBBvpUhkhwE/27/q
lIfG6zJ5066u8acbubpee4TD6Rc1mCuf8/pFpB5g45JCxxQrxEWHLhx5LWzfxALZ
J8UAWiJkr3R/J6J/JDW5WmweP7jhDaigIcGrzGQk6u/5omX26EwpWJJ8B0zM8IYD
2DFoQxz7CeQCTJ76S5D4QNpXz5eh2FNanotkHIo5E21WWyN04cpzCJgRxznc0Uj0
O3kPhXRLF317jkWmTO5l5pWJoT4+0ooXq4qOp5YZ3Z/exgA7OACR+fkhF1bgORaO
nFqN930C8n4XSO2zx7oJ6gPY2WsOldhCClC6LPGg0ZKqT9CBmORvPn46EZ8mX5UG
fVGBvyeY+Z8fraeIAQpz5jR09S7AbsVousWEutEW4LWQtAUaEpYvbounMfw0Y0Be
VwSFKvcHd9fiu3un5l0vZEhMG7oUJS2Y0iHIrhbPWmgRWF5OrzU19n59t/gSAPki
fZr400wbzAOoxSRizMHEOskFksBUc1CtG/zi/zlYVvdSuhx0+H41YycbOr2rySgw
oTNzl7kIG73uHS+rJFLLEG17I1nMLth1h7NclPV3R8CktVMOcsOdKaYGU6AFxpfH
Me4LRYqFi3xjmboA4bLrsSgun/+w6X93V5zQpFYSloX41OWDcScYBQJKIvLRGGZh
sfhR9yVo86a5gqsKJnGZIwfVL0Fw8Rxr8mAO2UThPE3cP2UnI63rv2Igb6svMjSN
mfVmkjkFa//J8pPXNFTB4t/2bVtaXenOrqjqhcizqtyGEoGBbgkjWLDPOtviosri
DuFBiyeHqJck0HZRXkY5NNGXY+mEgjH1dzGVndaVzP619BEO/8HfxhlwztmbUUFj
ayeSdp5iHRvoEqVAAndFsLqqB6rtKhiVYo/NiHPPtkcLcurw7j5k/37osABBreVJ
ID1FawyNK7LeHySWjrJIgMvgRE8vCrq65GQgpjcUIYeUrcvjWVdej9xPR8oUNc0F
8XbQ4q9hr2ez0kzbH39sNKeYWoCsnlcWAnpKd9nxwymuxJ03QGg9JQfAfGjGWmTk
Bbwiy+46yfO+bhkn8uh8mQVRNFIjamIJiPaFoSdV6PUZCvfNxhE8VFpcwtGYWsBE
ekU3vhtnz2AuF/1QcnsqTkcKFUNz6PXUoJKBjreE+ITnI7KmxYLiFl5tdpYpOEIw
jhPBIPOHaEVz6Rkt7jWvX9V1geoeIUL8kb4igwys42SwamHW4Gf5EsYQbvg9KJIQ
aRCTVYKXKkehDESR8J5ACiofzQFe1Bp+VKyFNoRcCUbuxeJxAU4HBGRN+lZlzpSJ
4iFaiuEto45VS8vO3cDSiHkqN5tIJNUZHgZMqumJ3w/xxPT4LYaw6bhtS0GS1Jj1
B/c0P6l5OT4h8akvaM6zUF3D9leOxuUdi9PTPlTTsEQcrnC22WuprNStb20gjQkL
oTF3fXVr8JX3hcKCqFRUIRDzPJ7N96MhEEgBZf96fVsfc4UmhyFhlNHo6d4YBXay
j1R1LxyltLWnhEVxGMMRDa9L25+EdA8skM8v2LAIHs1v4apBcu+9DcrHEA6iX+ep
PS/dnPq5hfJ/jvAMgH5T9CkKglt//jj4/TImoIuMdtmS0r2I8o2c1SKekRH/b0Gv
Gm2o0MSBMJgq1Eb0W3E3g3g+3iLoGV715NQtMQFm+Isggp4BaFNrrx+37ygJVdHe
/JVCaJGLSa1wj/BKJbYSqJeuL38o43p9jpocqWhAwuFBl472jkQYDeYgWQyvL3vR
ss6DpVJ3hWqBS7NmW+kjJ0y7ZGZZ4kXla3sVGcpYKpvi7YupEdJbOsdvuG0XPkK2
t62dslz67td0jmpkd9jbh77QbgWPWrW0P6blBP+0KGWi45LourK0d9CFVYJoswf7
yy+uZaJi22EL7J1uVhKcXV73H4l4M/TBqedg9jHLIE1KRMy5OjTr25HuzEAdugLw
kAL0/oLL68g2LFvrlgcUzpGnqrpQY/GTqoNHv0O+f7ZNHal//dTTWN8GBOEDEWn4
7pspA87vuqLElQsX4awviv0nJ2ntcs1LBCc/wY1Tp7I+BOW1aUkrMkT2+xsUHDDU
KuBg+if7bfo8+xX6oFhWWN4SVIXqwCa7iz7kn55vWv55ms2GGCcCz7zUcIfGSn3t
OsaI/dgRCRBZWDsgyeqbqSuNxS9jWmVoOh2zmWdYgrOm9s1XZkbIlWQQI5d2Cduv
qD+dADUUZdDGS6Dbez9uqgnZpYtdxom7p/1TK4VspmhlntMeuMGddhPBWDBDWlZQ
nIM57A0xfys3NSebSVraGFuNC6G2WSlhcHzN68Zz+sJRsJFmaMgjUQ+1GgQvDpiT
GbYaUDbGgfFohCPUi26BQFFErRcbWeHouOiXPXKNyKRqHImms4MVFJlLCnb6WMjo
5kqvmBuHCZZexlnCRkEA+BxWRjqAIVFMlBLsbiOvrAz+vXAetX7HC4Z5x+Qx8s3W
hZESx1psGfz+vsvFi2n5FFkcYUdoj03GtVZCnv5xbR532glgIY80vmwdwa5G+n/g
uOWUmRJGs4fIyK5H3pWrFi9SCj+eC9R+HcaMqGjgU4FPr6MZ0GofTCYHko00yX3p
O64zqm6o1e+t5KA0HRckonbObmd9gjLvkUUCk+mShYAg0akSVq8PdR5OPyLlAma1
RfnePtS+8z0lEd83oSNcttR0PglhRJJo/tiOU6H2uVB3CzIAkbiwkp2t6zi5BcSM
4K7K+7sgO/g6v5UqoP/cgIOhr3+emXrHw4itJbnNW3TzgKnGciRmYSxfsJbz0NtL
A02EcB9NJbhE4+mRfTR6fql2BXGRxa8uJELavXM48rtwDVe08+ehDFQyB71TjW9C
hyvsFOJfQYSB2T9SAZZTu2nX+mORE8yrmdLOo24r/fhxjde8j/si87Us3WQ+cg6i
ICw2/ZzaEj7W9E1zJ0haCUQDmTqRnbaTkoYIaUCMu/iQgA3Lr0nXuyD62VO3yY7I
VAkiQF59z3SJlinTtiZRssEwkpFwS7DCZDkkEIiETlV5p9lqNDKeR8nuzfaru/eX
12Mapmp2ESn5rheYls8HfiwO98y4MWUAdI1hSoDUCUKV3AhPsijB4Y0ZYdxdDn7d
Y6A3dT6XZQZjuT9/DN9jFs88iSIwalab+vgjhwZSo6WHyKcCpjzBCZv22GaeUBWv
1ygaIUN6uOwia452A/nbOXW4zyGrxIyI42LCy3IAIb5gUb8x5/WJa5kL4RrV2DMQ
Gb9enYiUx3BRpYvG3Lk6qwltP2SRQHo+iWh6ehBHiRHcyoQ9H4Yw8kqyTsMVHS4h
F75WVKStoYOZYFIN9VnLeBelnp3/3s4sGuLRL5oqNPDcIA3L7f83aMJN28vfHpdg
mPLZSro4Ev0YO1AOYAL2Gj6OyoeHdmA5V0VI+gbbsmUxiQb8zD19UY4OnEdS62bN
ECrS82/1PH2tCua0c1+a48nJE3BnuuNy1HPVg6a3DF2vpFd7sGGvRDD2tr7Y6q1s
rvaVuCaR3fZr0eXjQmzv84bD7A5eJ4gFDPx7xM6KQAk+54QFzOcyGGZg16UAuT6O
YYzQABeyN2ujR04e1FuLjzHrUS5QIj3uId7E3PeOupVIlzEwRazpXT/JDvO5NO/l
c/XuP13DquB+jKpzNP4/5A4+uOCBW8YKweJHbFARUb1tYDgNLSnXfepjGkLT0354
ABsSRM/WyesChKqWOdxMrLZj5qc2mv3j9VFSF0jsYVlpdFxTmq8WJHyVUClmaZPL
NAwE5lBnJ82MPuNpQh5lkJMZZTnL2HVrCabUKQvD57arqjT0j+GacJSztpKmRjbS
aSLHJedy/P4oDwdcrwbFsjUHMLV+7RPTSImZLFXXmNVQZWmdSRem7CvsSnLdh8Qz
1qjpVa1gBP/dc5ZzVdMh+AAJjJqHPUR7FojapQKbxyt+hzad4775g9or+4r9Cq7+
qNZ+zRfawB4v+ro+nXOwEjdUERwAO6hFyrAw4sgX6DUGJXBsxxPR/JZQWGn14E+S
bbJVjU0QrzxETNUvyshxCyj+itcLlf9eyjmpBfZo7hBkd6h7TCWQKjljuu72jsN/
Z2o1pKMunIJYV1mrMHIPnjdXbwlJjSKqtxefZmry57Qkw8bg8Z+AM0ttMzCUsH2b
5JHYl/9E07x+l3rEFQ0c78maAKsPznJ6Qu6uCNlgClUC/dunvFl0PqfRI4++7NXy
u3xKriRbKHhApt7h98lA3W/PffJqJVyemmJMvsV/rPVyYdOBovKqRKXuPtKVMQJ6
HP4OcKr9aaelAluGNKxEhFGFqSbbU0jaiFrMndX8xz7N6dRhy/t4w2ruRXYd9sN+
ukfZQj4YnBhazQja6nwppcaIiIc6r8GO+jFIckNTn7JoaHHoOYjxTh6PliR3pI4r
+D0O0b6I+w7gnj1GrHMaZ/d7DTj/fV+RZF3M+k9lM1MfhRlyIqzFb/4yX26dpvzM
23NIVNjc5FEwuY0TbTeP4JtKS4auDfp16+0MQBZPLMB03E5Olop6bp7pC4ZzU7u4
a/3vWqUAb3IHVpHZANmYIwmd4WTP4mNNRwD8Hza0IHyrtBJvnhp19Xr9GOBuiccV
UxaTr/BrbQ5XxezpBHVpNl2pZDVEcMNUWGWZr2I15m8yJkyXxXaBDAA/76ulQ/Yd
0SIaBjnuB5WuNcFU5Vyl+hV33Y5UrM1Ul70QsUeP/NyLOy9jGIoE7Q7ezGx+bz59
s/ihTOqdJC2gbb8tlS4gTEWYpQNPC9aOGZLlSI7mNzx7xEAjVW6TvsnYyr6KaI6P
Ff82C1P3Ta+nWNvkNOtEK1mYpTzPGQkfMU+nApJg6HTD/MQWdB/n2kFEzq0Z1FUh
LHAX4majkkRtI0mVaAHjdeUA9UMG/PAfn5x+XRJ1pLMdxw1FuGW0pnZwU3/6a/Kl
HJ9skyaudtgtldWaTDo1Ue7UxPVRMg8HNAeA72hnZnBnotQqdF02LXYZ8lkNZv7E
CytRHxspT+aBGzGYu3TEBbE6Pha2GfzzS1DEjlmYzYqpkM3BRW/qbFUQJalA1yz6
O4VG98hrVNN0fqI59iJmdc4o7PMkYkHQ9unOVErs+AM+Qoi4g5B9wlqLCMZKL3Os
2vZX51v+JaooMeNdZe3wA+XAuZZZKH5HUf8OEqzsbEnGYoeQxkA2UwgbRkKXudm5
ijWA2GwqHFtfNZMXm4xYSknCH7eg2fxjaSiBGL2ejl/RVGnhX+szPvdLrwV8Qxe4
S4Hlv8DhIfvaRpwr3OhJS2RP9y/JNaqHhvTx7RIxHji/9D7fFKVkGEC0ouiOMRRr
ouXTESEYtWcEyP2JmBiQEl9UoPUIlLY20Y8j350RbnL+KtuJP+Iuyka7RZhNjvGw
s3cjVb6nORmisNAz25aqksJd5vCSYEglwPr/T/Yr06jkCnQHiOvKx5x7+FdROFP4
+2v2+VMIr9AAKY22pUqqd1J/+t4Y23+62lKX6VBhIzs3+vMRFdck27g9yum7oHLs
IcHza+ieACaLStMyn/JWJGZsefZg72rJurWgZzMBz1cEY1WzP6ayclDAx5+B3E6l
T7xLcv58qOMZXJTivCTIosT0mLcjazx8VeXY4kfolXHtIGxC60X6gt7P4z4OI+d3
1LgyLvCXKzDSIxQ8w5lHOI+AR99YECbcIyICURTX/yVqiHNBrMKxYkvgIJSDk1yU
PlMiB+tAhbs3NKcGfJ6+foP8W7k9jma4nKXoLdgEWRJAjP+NcTXuOuP0XyHn6O9V
/V3/04WYB0uM1uTvlJKIZJeQ5XV8kIEs1dPkZoz6XY9FMU0DRQkQ6f13BxxvW46y
DW+UELSoK7oQKhhvSQ62adAe5ZlOy0KRSxfTr9KlkN4AWr/XNKa3bhE1HRX2RM3S
LJV3Selv82tdltv4JtcLvXmy4Yg1HIQx2a3iU4W7S2Vz/JlInlbO2TL7DShYXzTa
f4OEH7vLlkdvQBY1fozaj0bx9tr798mw48N3+IdIRPPOe3FaefBDa1CQpg9evK/X
Dt2gzj3x1vAVu3ZWmispPjTZU5bSavPFk0mFKoPww86J/MSjXa6/VtFFn34Q8Pv+
Km4UsdwyQw0IY6v4HAaMpC/NUw5itkuJc2aTuGDeRvl4E2nhXjT8TlIvSysChs1B
/32Y0ISKLnMqnHQVA6PoOTjr0WXRXqf0u2E8l6Ycn+atlf6LfkXAu4hpdaybsKbJ
4Z1f5IzBG6qI3aN2Rs0Mq3Rvs9g7QcNpcCtOpCwwMk0dO5mwCh831v+DUrqpIEez
NQT8iP7joVvuol2aPGZ3r7pkn9iNypzDHQMsi1X3/IFdF5dQvbLPZ1lzyFpp3luF
cJYZYMJCx/0kwud2bAo/cxFRYkIV/w9Q2yCDnkwvvFgtdbOcrIX+j+Vh6HQhM5Gc
ZufnYQ8hbx+qUZ9bjVJln9i2zooU6UYbcTLAbl3jBRxs26bzFAxCSlBO6HKYP13i
A/oQu9l6j1wtaDwQbbG+K6URUVPjwSZzdoXFlBfDvxnW1vhFB+ViPWX4tyuGs/m3
7itDzlztePB0A2TEIxvop5JzsahM1BpGd8VuPTMChR6qm8F78Dfq0CKDmR4x9lgU
v2PHTSWffzeBp48Zv5iGmQypx2Iffr3Qy1QY79Kgbq7V/hNW+ANKDaBxdHbGvOe6
6QJSW4OLFC6PImtCZanXaus2adqj6hHdJcuTEBACeSY3ZD7msF8JFmFaHDJDmmNH
aM9WycwLec6U8jUDroCquFwVLjTEUt9w/rY0nI82+OF/S3hxxZkoNxI3xRynvh0d
I7NwDOF3P5vaDlp/BPaXEqGZ/DoG190ZT9mgGRNDRbGr6Wd11PxQQE71Ab6FBDze
jQVhkXyHDpOqCRTyZ0b/OKQR3qT/gbWggrmw3jDrkmfwsVN1Jr91B3/NFWolEdS1
f72rgTM22dc2IjEnrNOV7wCbdSvohH6kdTJsfQT6IaZF5ViflUtEEzzRxP07/eS4
4inrOgbPrOxLkD86hWtk2ssB2DpDBVXMZn416kBSczxmxJGpKCsrM3xmLwUyhZOq
HW6KwvnDqd/g+ZnW7hY3OjDH9Ie/8xlwkZb9pIFollckbHu1oNMeekrShWz4A8Pc
MAge9UggVWs/7topm9BQxEv053De4addf0/fAPITq10gJDlfs4A1krUhxs+v9the
ttsoizIlWW+hwHOViLCASocbQkXMzl7Axn7wTwQE+kdlDsvnlLT9gQ9QYawgyjsN
njcEBW2QXsljvz1e87r+oxzIJhmAJ7t+yhavgDq71PyENww2v55rmb8hzQsgzYO6
KltjGInxuj71M5eMbBCR8sKuMWUHmmJ+zmpK7bNqbbzxoZOzTyrpZW8rmHilyXB4
rx7jC2Er0diLL2D74CaWZFgyzXizJFyhzx2E0ucby2JryyXfZcgUMpbtFZLS55W8
kiHxwYu6bEaxJgu6BxSwb2HFA8vLlwMQyv15OT79ZkBYpVCHfzLEGkuq4S/2mX54
6XF/20QWvTGYFupZLxCctLaHA+TlhmTZ2HOtx+b/UK+9qPw0GdEmsJY2xhFp2ros
toCDJn8aFLbpn6mj7EYUuclSFXKNAu/5RTyAsg2G7kPyi3vGfXkS6yjete8EAr+y
H2a1BPklTNQqeN/l3YuofjiicFfglz5NNDFo3lrmksxXerOx/1ZiSf53FpQ2Px+T
hVVIU52/wdcFaOD19wvXHM740DAjYYC14r5UMuhr7WyAgR8EGD5yjwMHL0Dj6dVH
vQV86ZI2nCt/ZatjOF7ICy5OumZvx9vR5Qfn16CP2W3fxiwgSURXSbNyuHOG3vDG
v4C3ZSBrbcrl1cPxlmdIZE3hVmxBpe3Zuao6Iy8dIqZYzYT9vpSbIzFFKJATgN4M
G8a1e9RT3PvB16eFZBbGx/p/5YuwOzsy8zkqcKzOppY587mutBsC1CjlrB45GPTd
SWskdy4udCuWfKrI+XGhR5GFvip/eSh2Tk+tnQwPNQ1LTQzC8aZLstwAGfID++60
K0KYVE11HJXEDOBoWnPQMb3NqLk43kXaH+RuOgC9OZkmyeGUiH94pGSRyS032EZ8
/iADGJ3a3pqU+5upfYjiHMaD9KmXJgVk11RiiBX57dwFIKjUh2fKz12MJmYv1fuB
iIML1JJAltelcsngGpEaKVbZGxyt0oyjERnrcp/48MsishjZxtZslhgVxrCsd3nQ
i01gcZGQ67/KqlhE2RmVXZ8UdVguRigRWocOxnJU8ROPGHDqGfc/VQNE76RquQzy
kDAtZGXkSb4wbnQDUUmpwi3R8DNWxp8RHljQTzW5vb0Av8Ltsl4EIqjkp8q8A3CM
6Woch5QQclvpA7u8gYx9CoMZa2SBtLvaitsByln5KKc73PntV3Z137sSdtqHNmHG
yx4ik1olkoWfkwbz9VEgvyIz00rjzcUUL/EHJZwJ+9Lc9Is0VEyd1aP+BXx5qmwg
R9s5b/TvwEFcPxZsNhfr2nYmQA2Y/CObQhAN7G4l5D1Q12JzHGlNKnS0IaDY2tpZ
RUoEyDPbP2xM7wChZ+rupMfzsZ3TQU5+lwzAddF/0UOqF3dQViG+1/QHTf/UD2Rn
E5/MmFnsoZ+8NMt6pGz3wSrnKGP1NOfQm4bWIhFYlWD7UBmFOr0Zy5KknLKFixRz
FHvAV8kYXjtI7AesC8T9rx3iz8TVvCNF3b1ULdpREmZMtKpY70qS5hIb4mKd+CZf
KliqOqiMwrWID5rtxrorJwr/x8AfDPUjU4QttSspYZotTbm5cERpmL4spACXcmWk
PzC7HnYDffEGseMLkiQ6FNUNh91sSHPDgOW/Fzu28zS16YIow4+oat/l11ZFFvOn
C+bw4ygpbMGc+GmxBXwahABZlx1yeoylZ/U705j+N3h7u/AC+eODQMDroT1zd05a
h1UW4i+8sieMnGRZjcKF+pL+MWPXdhLhEToSqr5aOFpc9+soFHVN9QyEj4a5MM7v
kfxrc5s0Js9XyCQphS0t6JeNGBmbetki06wPDbOyeaAbxJeVGZ+e91XEjFvhCp8R
BgEzsP8WBXzsTqvT8gCqcS/klL0OSYizV2UO7ehf8CAhodpYTTYW3rR260FkU6Bp
1v2ThFvyAvvGlheCOgqY1Iqp72D67ppXEPyVkGRc1e5+wcuZ+GdPPvk0GXuTVMso
5cKG159eJJtFfGmUoQEZRqzwKma30hyPi2A46SnsGKzjyFgcjVUu+mUbMdS+2kki
WpwEALEMyPm8LObeVNY7f8uwUL1Zgoqkkcssh9P85iyoRv+PG76FCoysFmxgnes1
kCqmuRScYTi/4r1PEDSW4d3shrnA0FY3b6iVD2Wc4HQ0LzQg5NlRKH/vKaWnFDCZ
SXI43jzAfJoDkETa4plsgFa/EdmN4JjKq1M0BY+sPHhBhWkXd2+yuLUEY+VBasYM
sLiB8AOk/E4Zo9jCutK6tM9Vz74mKz0iPcQ3K2xCmhMbAEBu+CJSQLQJWm266JcS
kZtgAngnNPf+fd4psCwWgw9MMnrUsxPn2mocBwiwiNFkat6rbWful/lPsl0nwJiB
X5ca9Rk0jYjmhvhq6mElSoiuOPbBbA/GFOg7+MGMJtTZiMvKBfZ3h+e7jyQzKe/c
TPWviaZDYOtC/UbFFV3vlxUuVK4iLhXO7ijanj/RWF/ELrPAs4tvKAGPhFbd36Id
VxZ2tDvsVf4Sr22FHEYvr43mwk1G14DBA0nM8HhKRikyOY7EK3leh/WsS5Q60v5M
h7UR50/eLczvZhkEBXfIzud1kydIIWcCKAv14+BppKINr8MrF0SlvZAAnhBh3ItR
pZzna4rf8Gb8UBlfdzPkoCDVZo1ffA48wvIG7wvpkg755efAbPHKK9vWwlaA5v+W
riibCprwMy4+pmB1vPTftMWQmVwtnFC0srIBWktwib12ZPG/gNRDJzo/aldLivYi
cLjSqqZC9nZCrTZsrWdioeCbIGNjjCvH8u+yDQjdY+d46zDViiqnOV5UskUKiyJR
qV8Mof0bgBQMRujBWaNK3ZLbZpRsSzgizyYb15rJkHAFLH6nV4SQKJm3Su8QD6DN
Hgc8/F4Qopk0EFLyiN8s7qdPHuAbpkEgqmDp9cJ+Ivnn3WsrIjAN8fFIn8IV1kzn
2YYrBesQxv9FsTS8r08wq/NBi4L3PCQAee3HlZpM8vzLzrp1gIX4gIfV78WL+KtS
S1b5OCzg7sgAfS9D5hQipkLbhvNN8o4nVqxiim0dDRbbvqCNdoA58RD8Tp7nCMO9
wPrz0INuNkXSzyVMxWjlp471FPOBE/l/J3kX/B+gmxK7a9n4CYa9Y9HAe3675Zx6
PtSnFCdclFSpRw1bh4qCKIfZMspuEvxZlJiUdhC/uKc0b1LZGlslJ//bxVRTny+9
ypR6SUAmHl2rnSPZltYPSIP+lOLlWmBXdL3QFN1wwtOQaSfkbj5h9lWGu8Gog+EY
a7LfdXTOVt6SjGcrDZOsMzTY8SZMDmtVXpATqiGb1d9cuiwr/zSHQfOqNCcLvW7U
egQpN7oJhZJbcU2yAQqqzGL2w2meFMHPYcq4iwqnZM4QHjrS3YAESU8NjsVHSHJK
8OVSEv26+Zmjb9hgHUVbo/sSOLOlRBeabSccv5fNRNSvJzKl6bGIkrdew4NrX9Dq
DFMk97N7II1qkq7BuaxxHwHu/mh4FEyB1KO0GWvM7BNBYucGRSudLJqfCjKS5Kic
i0qlsBeUScZ784bKqfDnf0gvWX14RaI2x91IyzG8htcOJ+wdGKRVkImcT7FxX4VM
69/7FPz8ofbqaxP1IH6ivTJdCbujMnHOAt4Vn/H5CAk8382tnn+QIY1hCjIn467Y
AhC4a02B50AtvYzVFvY3WeaS/cfCsBzC2Im2djFQt3fPfj+meINLQ/V4K2u08TcJ
ttMmwsAF7zTqjHpUZIXu+A0pa+Kz+lFlMEdeCYzJjtnBNIaHF19sRTOKZUpejbxd
3rfKJLpIAvDX608+Y6v+QJWH2o44O0xp5/FLa9ibNJPPsNvZPa41grKYX8CwuiR9
tKPLj8ukMKPqDzNrvz1pqaD6VNJRv/uA1CkQzUOZb2xQHxqaBhES5b/3mQOAL2I2
KRfmY2phjfZCkfvvkZja36th6OLOB4aC9f7XSDgDPbDHRStjPvkwfZBbgURsKmYC
dxHqbeuTVrOIME5YidZTBO2iVXiYbj1JC4bR9ini2ENkGWi/rOudbseqL6CUtWUR
7hfaRNxAGKtTsAT3xFO9VHr5LZtzemzdTm4pbHV3j54jXsxLsCah5Utm/qHYZjRj
n23l+mm54BIQEZbGNFsCeSqhk4oNRJ3mmUddpS4rdnX0x0E06VAQQyhb4eZdjJif
Ts+L5HYGbavvlB+/yCW+Ytg0ukGYgKNXqkayhIRwrpUQXqV2Db4E2lXNEmsAQo9K
zBdC+p5w+SU/GAsKw2RUf3y3RueNwDdso69yEeHxuskFLeHJsMN8Dlv0xt22LQtC
7/1x2wmHdJ3VTYHOqZnkJ554QyomTvugHgkuCV9tjbAz3zEVtWrhuj9NwdRtdXzA
9GnQoBx8ti2TjkavrnsD6kWgICYEP8MnIH385xXyfZnPmejRiJxEcJnHf0hxZ568
IwQ7Pa1G7IkTW2Nn5580Up93PlSWsw4PW+LX01I8MtxfXJyKdeobtC93OFAoYzn/
yDqA+2e5a/W6a7YqN2IsbjEh+IsLRV4HVvo8woY3DFSVX+CJErKJP5ZmfQXOd9+o
ClAT0iETih/60Y5ydPvKdWUhFRI76SXtbD+/JyZAjdBaCTwlMM3Uj83+HdYZuyzo
5vmWjQFSPGiqqInHJ/sQZOGEnVtetrDlGSW1xwxTl9pHhGWGnvKOUmh0uYrQIpKa
MLu8rEhSNNenxnXf94c4/I5m3xaSUH2MrpX7Iq1xubNtjJx04PqXcgtYDG0lcDz2
sVBxGZjhC5saz8o0M35BmllFYmATrAkOeQVG6uHUGS+HuYoYGA5DPYqZ8/430/Di
M+l+ialkLZGD5S3wHogvq+xz94YJKzhvCFLfQk0BoQYjqvonAOOLfUNqnLimp8g2
wp6DgYGurX4p05YCeiArmRr9XJ4YsaC3shWRgCrW20qNJUizw6dQYaNEa5nFua8d
H2qV37NRNiUODubUCduDmwEmgW7DYaWXpF+gdSAjmx/5YJGb7RxriWBqA77K/94Y
sIaJbp/frjTn5W1f+Pc+vQ7Iad8G2H8Rj0t7CzVrzRH4alrXvPE2BXv6zSZX1MSK
AmpO0d1ET995MrZ5gVHYzO1C6T1ib+Kg/1J/KX5Tj3aNQOMCf28pCNI1M6oWb1S1
NkVIFfo7/u9WWeWBFhhVxglsDOKC0S6FuxUQGjs7/YedfgwbVvZcvnihI1dYfLVl
ltwXqlDnVENz9blx1TghsiF8dGHqFX8FkWbYCxLwRdqgzZGzWdRgJxhQPL5bhUdA
kuVxA0MPN/UAOHdc3yKFhA2jkn+9vfzLGaeDXGk8malAD2Yo/HGdRdwhGQzSjKzW
ZxzOlFRj3G7KC1T4va0PlBuy4cG/7qQuySlCiuFBScUyY9wNzVOnQMLeWH82IcKv
/SAXtBxAxpwXTVFzzFwQGqGQx87b/FKK9/O1xNOIV8JQf1A4+bsxBCj51OXMzMm0
9BNC5G6azdFBwL6DpK8k7KTiv8Skgvp+q6H0K6eFVPcustyLlZGayQ4BHDq00+pT
cMqA0SkmeTQM0luCyaBcY2od1RbzP7lPR6+O3fJMKeJhzzontGU7g2K1TFXT614y
tLDY7WCxvJWZjq/cO4eoe8z+iCOcZZmV+F6ioB5JB1XqpSq9to+A7BoFUg1qbePl
dZSXMB6Ms24807+gayRSsGdJauwHUK3yvmPMBYgexOp/2/22PhUTEMoJjFbDZOJz
Pj6r4yi11PUOpuWawykHkvnUM/e5KAH7bxtTrJjP6zVFtrtG31U7byUBF9NGBJcK
feHkmGXmH2OJMHI3d09hR5rHsFXK8EXbaimgisjxvqM9I18MJI2tcHxba+wIxDlq
umIWu9K52VOjWnubeEIje5w9T6F7fk/q6Q/BorIIsbvRlPZVl4200SulrlUBvGCx
ajiXE0DYvpcsjdjpl6vjPP0ydMtwRRnIfHQm/weow4z/hCGm0OBI6eRzes8QWnrf
rw2aVcZMeLcSS3ZqtvGLtyRyt9TowRZqvIWCLV+fwyAX3XFOhz+4Q8novzcQYuAO
GXyCcsMQxb0ew8bpGXj+KZeR0UMW8iSolE8GgnOUnvwhagMhLG6eUdoJhwvPjfw6
/S/wHKIiRJl/BsME3lEFbYqZ7+HthQGZZ6Io+48oAVxLxZ+zcy6EduwTQiQ5la1z
M/2a59TDywOSNhrhvTpzWEbQjkGGFnCLB1o0gMpAeR+eS7r5r/Xmwx/MRxMTm+ym
P4gfGM3wZUUShMGj9XoXRELYAtObpUM7z0k8W8cuUqvC24iWXTVfg44RQtI5YNaz
T/krUV2V9+kHbwpxWB4ZQmtxEo8Lbfrs8eGKO2ctL3MLRhGVLi5mj3q0/Ko6CWXK
2nfyl04+Ranb545+cCeTXEs+HhnBxjmuBHecYby/kaoo/fzqbQNq0z+1HmJrHZ5s
c/bSGRLibPIXmNgQL9vUkGO6avnsiCU2cXswdwQSDPVIUllgp+/kzWRSGxBfzJOm
I+9dBnlwaMWONDszO5KimRhjvR2bzVl9dpOx85HA5DYJQbNxACfprQmxpKnMpFSB
zbst4GkjANNC72CJqGe0UPkf8EWzb4hShfxL84BevLUzUt/Pxjel6wNG9QtJ21MV
hOqdW6HO8fW7UP2IrEKCsOAyv4BZkjuNdASgVMBalw9kitTHKMDd7gMI7+HqIFOu
wbuYlqcd0oDQ8Nvyx2gk3odN8IHNhtiNWGloot6q6kmpukntQak6JrhjLOW7BWBq
Ov4VgaiNLrioOjhw6ehDfqB2GJshgRRHxlnjpu9TmfLb5X9NW+aEgTlKGWYB6m4a
Yd6jYfSUqhz4StMLdIvbTfU3xKCw64yZSLDEtsDwZJ9oF/e5okhlo1VhT4iB/41J
B0rHxT8AOvqy+1U1dxb+N3Stn52Jh+xM30mmyU3YwfRZAnZfc8yG/bnGYMRVq5QW
GnaN/WQMZ62Uqv6lifNJtlg7voxgfnpkTJ3AguRWBUf4zz1lu1kh2EtenCOQUjK8
Esv9M1YB35oxfcTVRap9DBFFPNyCkwo3nrrEq28C3Ry8tzVjC/K27oQ5bZoKA6aC
lcbR5DQtjw9sh1cfeDSsj5oKdHQLJPMmXSnogeRG+8FUbu03/sJUV+E/TIK+xqbN
PYmpn8SthNqAh3hGpytyTKGVWYL9EbVqq2af/Q8t4R459ZATH4X22sqKCheq6da1
a2aUxk8CpVlA+RRV90aV0bii1xCG+aEE2x0dFiBe5Z0YHFPpxyi27JY9fJ/l29nf
p9IZBNdLiavUhSwY4l3mSVSJSwCvsCgtFqH49Q+dLJjtsm6MoVSExia/NqmnqHRj
J9eDzt/+7O271krlNqC+262u7Th+5PcX9TBBWR+9+eUqtjXCCKhhWCA8eF848Ff+
adi2gumZXyWJRf6n7xreB/cRTTGwUA87L9OHeVyj8BVF5fVSKoy/KcGbFq9f0Mvu
CcROdCDoqkU1NFUeZNl7zVaB4UbQUZklkufuWrJeI4jEQyd9iDx59Xo5S0y+SIRj
T2NDNGO23k/VQQKrhqd5yHBXmjHWqrBUg3sr5mR82qeDBkd04naSWeRXBYUBrgWU
cebItPqIIfgDG1OB8oaJLE/6sUoAB1Ss/mA9aQSUy1e5tOAW8e/RwAh/7bnXfd+M
/HQGRQPd5/hIDPQj+oScavPkPfSahZGWVyWK/r8V2N8kDJkYxjirDle4dvoffUCP
rW0jn/nbIxrs9jdbNjBzI6qHTZ99csdKu2M3dEnzCCt2b8oum+FpIrc+Rnhp90pP
m6fxvNC4jYEHSHS9kVMm1w97/iD3PD+OhGNrV+oBnhGnkZ0HZtv8sk457vPUydpd
4LHY60vCbU5Nj2uUr40z2AJIPS9uJY6ODz24ARlyNKuHewrDmDuDt8NHeL0xrbzJ
F5HFAOGyxeifQdbzQnrDn0SmgUZgub5MEOMCZ76Ahdx3qxvvadfLo3AOXYcSXNqf
TUSt5tCfsweUNOMIna4rCwniaBn/CfiJM1yPbqHz2j6Xq9KMaoUysTYF+y2OeH09
y1rWB5ik6y2nYQy9/O7IECbeLBMr501s08fMEpDb2+qBsJpJXmmPJYidKWRfutrW
GR9LPAiubmDgBgwwdCIhKEKB4dZIorX280CxlAs1sDAwLIBHwVW9tzZ12gd95tiB
qRRNP7o24BCbgV+/4EeG0fBi3ssVOtHN6XR0648l3rnEj6YfTeDi+cgRhs5QFUX6
WbKDh4RjyYldhAN23NdlR6VrxiH7She+FM1Jrjezb5Ihvu/rNx/OSdHfJQa76yoP
qEpxOwEuB2BwMNcSd+Laf1NotEa1v8cfKemgtgMkRewW45lPtvdZHS8fnZZYHyV/
ezA3j8nF34Li5RUsa8+v+/yUjLlP6GiLRvoYNBpxxAuqYqHIIOj1d240szil8vIu
2IeLZki/Rgseusf3l13AK/yydYTcUXYJfrMi+2YiCx9uRyo8Mrfr+tMJxhZ+Iexb
+VUxUOzlRSmE7kKDdQ46Ne6VgbFlLTfEc9iGudd9fKD3z/tRXUTOA7DC9vqxd2cQ
vqer0SIvnlVHiy39B/9ZOAnSl1kMgBYFRkjT1z0CbJkoBkq5bAjBAbx5cRwjqlbf
Q5+g8cNrTUfzeZzuWKYU93K4b3lmfIaPX0KH9dij8mt80IS+5+mz9nR7KnSDZY46
W7C4nnhX7XRchbebJctYVXEc95/9THInWjpk2VdVCNNKrtx2xMrohzklr1lH1RkA
iJOATfaYLf+V0r7D08xCbv+O4tuUKI+DOtTbx+NhvcPOstVUhgbbW9mqjLrz9uC/
ADQ7QKDIdQjNkmudg3zmxomDKP1/4JG2a5jONBZFnY6QnPXkLBIomw0SZpoV/OT3
AokEEuqpJgC4564un75X6iMAkObjUbvz4BbSn8vjWPbRhX+RjyTH6IqK9dFy1JED
o9YEv1SpXqwg1btEoZ9vGJ517UIwqKNxfJ20u/pswTUMHJcjkEl6GzYNHFPbe3Mi
NyER5h0Xrh+S+H1T8mqqwly8tI2EDE89H74bmqv8w8GyRQdzreZhTKlzWuCkaet6
JrlZIoiLnJlvVz6hmen7OvGD4x9e3Jt1vhcUpPvd5/m54B7SeDweFEq+fV4pvht/
3cTUKCZ4n4cK1FupZoFl/r+X5bQTE1/gKbwrghiA2RxbiI0Ya0/iKC4eymNgJLs+
XnpZp6fpnqX6eoZc94vg03gvLQM2TmacVOFofvJN+PGoTsVubG201fGNYLJsM9mJ
OSQgQq6dbZpKTQdMQvTcUJ6I3lYOmxkE6fIxopDCwwMZJfNpPQaRHdNYjb7zz/D4
PLZpk2SVGNX1yViVWJ2bZINB5URUF7eouILZYeQnbA00ypc76tpdZe9BdLtbnRz/
+6l5dKT7XCiB64SdPqlJoFDMWT23I0Cvui3NpgHBpRwXA1vk9g5nftWQWZWlXdhx
4z0dKH+eYmgeGlJfEUbAgwNJvCK+kITCiAjmRSfEsb6P3ugo00sIvC7iFaM+CG3W
Tq4gAtS7Vy5wy/+dD157/QRdqDlBe0ItIm8XGQAgjfmpb1ZFNwAbtiwlYA9HP3af
yjhjkzkrhcgPNwu64s9XF/sGLfGit5rqWhkg2Ng+UDSgQvxe2ifTeGwttUcAvOwz
Tyfqcs8vsWwVgkZkmwwH7bwmGip2wH8eWoIz8DURugFhQyhKuLn8FIvAw0NcTlAe
qr9c9ld4CYmev1G4IO2OKTsXEVOab0SFX4rrfsaSQFU9zSrD/HZqQBv0WyeKjbWI
KWf3A1ZVVQnVc+pTCbAZW7uLQ/mQY/Qv0yAGy8QCsJxJdnvJ9Y14l2DpmwhzalWn
QjqwpOBpQr7bjW638WuuPgM/mxz0SFtWa07UX7i23nhuVOY9qZLgb4mh/ILc7q3R
S/9nhnGECgGBBKagVNL4KQE9zBoWy7HZEr2bo1A6n0lM7t9hg1yhKrQ222iTYIGs
WxjDafs+WeVuRcCrsT8SlLOTBFc/JXAlKpLcAlmoYXj1I55FbUNWPu4+K1jwgMGp
Pzi//dv66n9WC7g/h7bmPU/858AvKSsn1RYieS+U7nGc2Ws9CD2Wl3D8DPOjifVV
1f90HZW1k6t7zzNtIGPBBAymzjnS/i/wMnKiCbSjWjH6eJEaX543WbZk64puu88i
A96cZOYK2YyjUMvsl0qViwXsfYapwP7yCD1eghmsxqWabSbnyeV4OFNyz+JCy1as
p251jqwargS7DfK7hj9+wdiv3cIZ+iz7WbPlqby5afc6YQhtMPnrdkxrQwiZDxOZ
S3A+bsMA3+qVC5cSBjR8St3tug9ZmLKJpnGWX6Zb+Ze2iWdmsT8NkbOovIswqZog
8DucGuVthY/bCKp1RO7FgujsZF31I9jWo6CuFPBFhDfZ4kjbnhlJgjxq6WYdWVmr
6CgGqhfqZn2jyR5ab0xQSCSCG+88bjQjAfhNJsu7vQsUrO/BFOUsLb/l6nttGB/L
hCMjqLGJHFyRwVLPvZ7w/lKuwemEdVo1DVLLUgWhYed7RRi8osjKMkUPfLGnrWju
DLSpyGHfSE/edz/OfmIS9uBOjq3eJgIEEqiZIxXCDkhBKmc1gtDSumTT9cbZt33v
qI9a6muEfS4KbheFye7KkWXC3B8SUjCi1WgBERdYSIqVw/O5LKv+z84h7A8lLgEq
OLrTpiiBI9+oCGw9eGCFMzodAo+WvUkrpZQ7wJnq0+d5Lf2L18GcxFzLzIjAYWoP
+Po4Ml2Cka4N8Z4ZeTak0ALV2qGY/v37+Og/TM3sBboPNkJY8J2UvRupBr0rBbBK
PXuW+R617ZMQlziv2zQVQk/Dr+L+fOzfVBlabpA5MZYk0xDKVbHjP9AkQg9ZMKA0
8Y9YljUZkxqXuRRFfc6KgxqS07V2heAb/dQHefNDr5E3K41/iPa6h4EVVkcridVi
f6lsyBntj1UaIBXNPYxM/84DhsD7gcT/f7CI/dhw4svmRT3sri/+9SWeSfSP4E2l
l4+U0EBvrzdN63n7KoW0UGGee6lHKzW412R0v91Fcc4DcJjN5nQnqdlQFVlVb6w8
FxGJaX3PrqoQhJxp6q3ofW+Vc5eZAG7Y1lmrWadrPGddZYUiBkfR0142/Llp/HTM
O1P6LSH+BEmhUSJSw7URTQSTgOP4DQ3/w52xe7NQuXTbzYQSh+TOi6RsZcWfvQh2
ImbBVRudL02CJT89n0pYHvAzU6P73VGD5/dgH1psb9Hncj8MEjHx8ITTaCBOQNYf
rUztyYCUgZttZam341LIPCZXFkD+V1/hydCFfOjSV9qkDbQEFTQmC4buaM5qzhjV
hvijxiTo/VGNnzfFJJnQTKM7zUJ8LXE3cDmp3wBrNhb+6sW8z59kAfo7MXJ4U+nR
yFAl2Jk86Z3UBN2ikV10wYNg0DKEYRaFy8pSeTW7vicfPcFMZrrBGZkwZZQXVac6
Y6AsLfmVgTIIdYMew8tR2L4rLEVQZX++kMH281V/DS53aTe7sCW9ksOiSQ56R2wk
AW3UOUq1LoKeQUOQ4o/41xhC/h98Qaa4tCjJlTM72qXkqUWna6g+vq6W3CHIq2Ec
0XiAGnI7iQqTP+BPdmYhh/Fp/wzDSqK2oUMIrIap1fIgSnjbgHsIgKntzY+sbHud
ldm9XlL1CInyL5F4tDHjs9LXaDx/mYuGeuhomJT1hnk6j4mMDG0ksIOz02ayGick
GmWrQTBcTrgAOeKcwktZMCKky21vXknfXvfDMM9fIao4CpWyxR/xjVHsubxmLWcw
GDEYr8OMU5wvtZ7g6e+VVYS3iw3BNh71iMCos3MuR6fnOx8H4EQm51GJ+Ikh2GhY
haiuxo1VRtGhhQFGq0+s033r/cv46pQWlYG3TRFLgfNj7RZXfVLe73+T2xlJa4IH
n8DqRGWYodvrxFpV5dPmAsz5iPZv1KcUklDSStThu3eIT5U1yUdQTxNsP7i5dtkl
68XscUNwUC0YMCHeHqOtNnYZEMZCSUwj3qXl+LKOX9uoxyXQCuDbmORZDc2xjS8Z
PCZ4sR4HE/DbTM6U0CbNcIVs9Oxama2yG8pTrPlhQJJBvw4z2vqiJnyVM2KDviPp
/FUY9w/Qh8UiHYz9ar6bh43Ptx1fNIRiP01zumdHWzmu9KYULC2eHoyKtFDIU3K1
C4nYQqgoXIHoICasiDI14KX3x7VqYNh2fYMURKIIB8ba5n47vjyoJI8MzZ9cTuIw
vjAEc678UWfvgnZi+fwfH36pim3MlkIrLj8mA5emakxcvD5O8BRTYuRRo0seeRZn
4AlMX5wN8mvDVLkyBccbGYjRue/is41QFRr1r+PIqGjBnDPEi6PZqTIRa61abpQT
VZOi897gIy0z+h/SPelqLoq4tCUzr5ewk7TYIWBigLf2VaRgZ0hYyA7iFXsAE9KU
OOP69k0FVoA0dvNSoEq9Zti+DENULUCG5g80wq9Vs9DLD90MLmfeuSlc/a7x6DwQ
oLONM2sRZVQOEr7jFBjJkxmt3neUdm37hPGMJkh6Bu26SPQUHFkAi7py0eVxj5iL
3SZ/ZxpB0YFJXmTTEaW7zfqK4Fh0bQUNZXvwUcZ8Rorgf3Q990R9GmTD4hwRK7kx
pxXvaafUGB5212PDAiAmEmSmjTPg5YfOZ+HQk4gYgjEj29Q8MabU4U+EemzjvMUf
If/+WNOyk6MJ8dxLgH4tebzUh8zGUC4eEbWAjSYw4dWxmLVOoHNrObZMB7Hx/2w2
WSIryWsNKVFOU/+kJQOFHHN6rOwJTsi2viYosrY7UPBpc1j9KDw/dzzsqB8SAM9v
3Ex6taASqZB0mt+AFauiOi3YWVIEpDct87u5WHXJdT/8O0Gpwp3IW8ZtKYeqejxt
tq8Cbw08nU3aFMNz6HOlgqE4SEI5cEFW3mcXszxe5gfLpFcgUchXP6hazJgOKu+n
dZHLOMKwtB+tAMzktRL8UwyaSMcFNdokzX6jxQZCxuOpijeTLJWX7sGNHKXAOQ/s
GJrkKTIBGAHoNjIJA88eealvglfGBsnX3NsqzMXk+48QdI4NBff7p1DlHue4Kdag
kJq8bL6meWClRFvGADnNkw6WPmn+EwupXPzRI8AitusEoqfw1sJhG/5JX/Nw9WaI
xTqCj+B+jau62+GeHTatz8C3OoKEXwD+B53j7k3DJJOpPU3I9HWjNYxLABXisqfq
ZqLSJoGYYQA0jgEUUuowUkXp37Lz7ilddD+JZ9J/pVjS1SyQrQlEYd+Dp8aqLl+r
VsFAOieXzKW3Z4HfwCVzvTZajthsdQS17MwcNKwRQCBU4XyB+S0SAae5SFzgVH2l
oDxNCu6NAFGR9lO4bsmwOkIRHUsGQpFsCGQZdgnKi0Kx4Nf2/CZ81rZaYdW+fFu2
8OTpmWSXY2w8HrtwokUSZRpd4CpboyP57AajjUgQaATMXwu2XMSYkU35lbadDiuW
/FO/hy1s11MG9mUWp4ChDzYmHPQhrfUY7BIRGSmWUf9HlZbI2tydRyYJYZt+j4L5
0MQ28fs9p6t900mdDDZ/KyzMUeRMY7C/9za9ifhi0b+tJ9MRwPk++5Q5ow/G5hjb
2y8cF2d7FTB9/mProFNTCLmJe4/F+7SvRrVkv3O99419SL1gaSur1krAP20ZvuBj
Hkp5sQWVNZe2nOzI/AzDR63aXk0R4fbrPcJpCf+KOv1mJ/IlJZad7dg06f0KWvkA
Fm8DNmqijmMPeRkzjpeIOEpeURHNy/5h+jYCp14fP2kJjI/Tk6cKASAVS3TDM5Ry
i2SOkIQI1iHSHPeW3AH6j51wUB5Pf5BRumAQoff3MoUWs7B6y9MTjZR8f7Ze/FGY
MDGW+MI9FVHkuUxGZ7o+N/bYNYeU1bg6mPudHHuHbPK6+aEN1WlSV8JidL55AU53
hJXjtmFn74J5C8EyPD7IHBER5DGP6fJxxRcUy4mssAHykeOsVV0RQbKUE8SQgtFX
7xDUtELInnjpMq9gTZOr/SBy6AdvbKHNx4kyjHlf++MIoHtAVQ4KQbvhJ48nagpU
JpvAkTWg4Ww1kFkO3Ipnhe5d9+8Jiv3WkP7pekHABWrMxbt59wDSmj8e1wJH0dsO
CG+llc8xlYyWfzdH8zwiQYcfbSJ3/SM9qp9RUOEYqpy6jZTRcL1WnDU6qo+ESV5b
3f97zM/BQHuh8BLQQMIQqGdxPGPuOH5dWE7vyhHfKfnBX1Q6NO1wUDLhQUqfcgVM
/y+FafNipBkRSrotS6WrUIJNe2SCXuf7g0bEPXmEidmTlbPfS0rNSlnJvrjC42b1
XSPikvMNFc6tNjT0DcLR+U2Xw+PN2d46lncB4kaS6kAimxO8b5t5hVD0C8BriF4I
vlUvqQd62lsxikiyNc9rpKQGm4hX5AJRF+1nCsOwAoXQP0xmJEvu0eT5QTQoRnp5
WUHALq7KUpoSg8pf//4Z9bW6fL860eT90pVClJEvAtnO26xPd1hWXV+F7cII0jAj
u20PUTSARNzRCgW6LAi9eJnCZamgLzxb9J1VWID4PevOJc57uduc2cQ8qBRfif1n
uhFzHFd4p8fbATAGCeOfDj1ikUxu3829ERs5VHe2M4B48ArknvBJ4KDg1lXFVyn6
KMlb8lJzeCFt0T6udPg1Ix7jj/fHgZt4fzhXOuqkYaikqiWM+pzftZHiLeLRZl6T
7DfJk8sssdhmqOiKt2kkUxz9k4QAp2oiXRhdR/dG2o4742U88QBm/5VuXDucldHw
StTtDSIkvXX5E3T08rrpj/hhqigFtPnqLsTv5JGTIqsr48AOxbuJOYsosu17Q5mD
hDjObRIYXn7aY/4XPcIuXq1hjKyypMFEyckG3Ltq6pj2T5lHzwk9sPeg+f8ZaPEy
bBoyZbhJqom6Ix8haKEmEu6Mr0NhEN7MMv8xMbEq1P4FtZVY+5VLymRwWZ/wAM0G
mA56K//tfIyab/v8cMPiohvZGnwaJ1uXt+aN906X6oUwYQbwIS7t78YeEUqEDTWk
6rs7K2b1N3RDZ1ti1vvlFCkYujatycBlQF6VGjr015zR0+7iol0iQwXjyT09Fpcn
MRImsoSrnwhQbrne26DB/9Krva2h/fRmRWKahhomuFYwf3P6c+QYreM1Y+2W3Yse
rs/cs5LbAOjLj9+0S0YDW7AoDC+ggyuxN0/qTn09fEg+UDlDC3hGcmGVoW2aztWD
mF8Ja9STYUrRr6IE0AMF7iPACuV6/cvFvRjczlqtxI72IoZ/UvNDpB9A1X1XIH0T
jTWbpkni1ehxiEjix6KLgsOokYZAQS9Z9qhExe54FF12zxiWWY2nC4GaQid9Kdjk
rXCjFnCuYd3Ov8ebEeVNDT3C5IKa6fyQqTYeX/ohYStNYXpNU4ReHOFgt50Lzg7N
ZP/B3iy1YteQlCmK8RYHQ5SGOyLRKejLG5SD7JDAHxhxxuwYNQi/IjeCu0aZSHzH
4XHnuP/KRqaylvB1/I5WPI+G1ddBAG/X/MUi9yIiUeK0jdFZprqbIigODjfKNBSn
aCxDHEPQGyd84r5ENzUH506h6PaqqPO0kXJ7ptAx9vqBHLERtEx8RZMwrTovmUJ5
VJtRYL/yzpaY+YhQ1UrHXER2DJCNc+3BgEJ0qmzKq1o3Pa6gHRfqq9G79p5WJivN
5Se5GLGCXKfuQFYDUTV+E4QwMpLhFYYRbxYAoO87RNuX8EXF5YauXExvVcCfxk7H
HHOpTmiI8yLTVF1wRuM4gLzQKXLmzJ7E44RjzyC72aQ/LOrnZJDc4i+XDeR/Yesn
ENMx0y8C9u2tIY6acqmq0oPrBzJ/8YIbiMyx8gTzWlL5H5vIxfbr1JmReIYhZU6+
+ZrcxVgnT3CaUK9AfWAA9ku19vNlRtt9JgkQiAl7cdeU7SrdVB8yCJ+HEiu/9YVi
DBh1LQJDfKhT6CuTFViJjl8xx07OMLrib7KpLoGgj1yy1+hPpJJYfsmapJqqiiq3
JubtIdc6d28rfcJC9a5w4Y3osu7+C8XW8pIiF84wJcrwoX/+zMlmq9YBamC7W8fw
Zx+8d6sPwFX5IQB3p+SjH0zJ/eNiS3deCmir5qdArKeDNZ57rPGu6Epcil9D+CtI
iA2/giHSs8nqGfqHDCm6SVvo5ADjefG8TLyfSAaqaqb0uwF/J0fv6INKu0bCRAXX
V1DYdZ/KTAnLiP07ZCC5o23KYZshnb2MVfSd3Lu/nReqwHnaBqxKvG05bVCvmrdo
YuqBBy5pkIRfa1zf6SRw6vx4Fnyo0rEZV6ifCgBwhzNh1I7iogGJHieSpvk9ggtY
G3nUmqAiOuAI9iMrdiwIxYo1AjMEi++xpB170ddBskomD8OA0WY0t4dGokg4Ol1q
sV8O5eWMqhRhMx6xmWdhs0ZsFhW8iPqG0uQrrk87W1ZMNf8RCFjNCANdUM28iSqi
weLZRfjM0n/DULh5wB3mhDBUf2LMZku3Mg0rcGjWrDVJq8ZOAXGd/1Kt6XsFYMhx
xUCXXeFNHmWjhIq+JL96bH+V5RK2gV9SsaYipNttYpo2hbab22I6b8h9ZTKFPrf8
bvSwhXCLKuGS/RpXw4+xsU/krjV4BTxtFcCmEhUrzgHcEW71evMsRMyzFtSJQkm1
RADmuup4zK8n0NreVdE1K/n193EBy+bZGERvL0NAA/NKVrCf2W6shqBxscmMEWuc
2M05hiLJSB7ihzrFzUgO6mGsn3Rein9L/uUpwSZ15nSk8baXSUyFudGpyxV0rdAj
wIbnVtNXPgRD+ywkqdFUqoRtaWGtcS55alhys2OEVnnB4yVPncVJf4bUJbnwZAYM
650eWokBC6S/9ZaP0pklMhMlXNDf70vHkOw+bJj1ZwX7pjltCFeOIqTRAoo4S2Bb
EYQaD6XWXYOzBpSGjUn+XiDpVYGHRE5QAcsqZyGOp1EO9KPibhhcQVq0ak5L4ntx
ehl8CAY6xWukqf+QTkusb4SRB74y6xRzwy1+68T8WX3NvZJ+B4qWOv6z0+xrPOdF
gxKcj9Wbd6yy2BztMylaG53IHfFNJYzL7tZmJUj9MQjdt1E29AEuKfbfkXP3TJsE
0ekXDe3uzztOwYNsjiZ2jV9/V7Rv8Y32qn4TcHCgSCMyDh50Am/5nXp/SD4FrIxr
gFgM9FncBl8RjMQJjoe78ckoFUWW1d0/DujZCV/tuDvvjBvQ3q/Yppj84/asVj1I
OAAHe2CmQwtv7Jjkq+LILovJ3i9V8kIviR9TsK0w6mZoh6Ln266LNsckQV6kexNI
Nyu0Abt98qgG1/qTzthXt1ZEnHR/N6THwH40LpEMg3nhhMay+BTR8rx50RoINHg6
tPKuB6jr3MdDRcRZiYaoBpErSeiH/1SX6aS2aqZhhcISsFERYRyvbSXE4dHtS68A
wpdpuHwt/ipvalJA2BTTsIZ7VDAQP6oqa87vWIvq+IxBB/H+ZgB1kPcjMmU5NSnX
I3Y9qau4A0bg6DrcjqnfhzTYCaB15AcMzEhsxAqtLi9dyFtm4eWnvTDEXA3t78D5
ZAKcnQVyb/S5pIvpx5OGPDzpudqDJtwWVkxSsLkAHPTrx8Ani2YZVNHIOXv/Kgx5
p35sTtaL9rxLZ53wv3kZ1CWJJ3x1Z3ccnHtoz7NcND1OVg81JxP7pr9kCLRBnrnQ
rxo8t03Bd4WW2Lx3docIW8Mj6cnswe0dlvF22i1Uk3iiHC1uwEoO4xHVrcr7oIaR
lXEXJ4CMiuUVbaAa4RLZVHfSdYlk48/YVALiPa9CcJQiyB1L7DZ4MxItFD0V8S/8
gnVLjuutBIxfDc1uHUoqNSmbEUXsIoMInxrdPDW8wHQbqbIBsIYJHAZLF3rCY3NJ
uJ1fsrjmHi5kcFIQu2hxBsUKr6DOLaGXliqgRcuVs/lo5TMhFmlOnyR25OuRB53i
P8EgV9UH3WXYtjbP0c1Dul4w19Agv4UkjTsb1pVLfRU1XIaME8CiRQgh3rYRLpxe
84oEGb2pNVuxY9yZ5JOjPT9nnPnXawCIQ/yecyxSztdHTdO0g/YSL5RTxtB9+GcU
lDWjgj2pi3qlLgIKbngyYFf/bxajdzuAM8eOGsrbt0UPR9xFuGJUwaPKMetHC6C/
odDFPlBvBdrkAzt2ZPnXtpkymv8S9jDlLrN/bG7ckNpLkf35cyWSErE9ePEFotMN
6+8mcBEGBJ3xiXWe7YybduN2qz02DnT2/m2P9A1Ub+R5g2YW1qKneJT5vTG8Njde
gvh/6Rhy7bD2ox+WiQ8zU5C0+/mirHxJNhSklc9H2DNR0+ZEaqAmaO7XaBRv11F+
0SO7U9YkksNweVXICq488Qr5IbKzBnh3PZo2dqju44lryHK3xdqXFDh4trrVY0AQ
bZRRt3r6YqSWHTz51tl8Um5OwNIjsJe0OOEuw98NYvZSXW7Iom0P7TCiQIthpM9q
bv1Uc4+Y9V6r4JTZmwTGn1MzHtXN+a/Yp1Z5u2zQ8K8Pi4HWK3yLcOz1y0Zqc7oz
4d01IR2X50xTPoQR8NXsDnP473rOV8/upsM0AYMWLwrCQm/cp76+WvYdPMLFssbI
EDGY39KwUWpaZgnlsS5g6AaiDSb7bm+MfRohWqOg/gsnoU4rUDF+PGpUuWERMOSZ
sTbQO7kHGMGyZWamdLb5WnJUORiPPFg3mlcZBgIBR9CQ/r876HWL/CQ+5XBxyzQK
4VZcM74REtqSlnhQImSnjjDYXJH3OhfVN2yjhNIGZ2QxMShHjdViXZ3Sq6p6MvXE
Awvdg1Euf2kmDwGe7/diGSwVXyF1dSJctbuovAc2ibDEs03Hmjd19KjeHErpRSzL
5edJuUqLpu10Y6Rlj1EVRbXK7WTU+BZ36Vxg6v/CtL7do55bCIupO4ZG5k5StSIw
o8f9egDK0rhr5CtRCvtw6Eq1y4wfFt/pXPO+cqbSm2E3RmjkNXTFdWuTc+XkxZqT
XCKzCGaOWHI00+hZvZgDiRyJLnYe/u3leYqMbT5EpzCZwxo8l5iRYqDoQ3andh+/
4Y5HYCn7iXDp2ot4o3ZOAgPYIRH065a1wNG2ANr0gXKS1Go7VZDz8daA04zd+p8/
X3zSgBEKybXjyAmD2GXQp28nbN2/xUBhrsGKz+cMHXaWxEbzkW/UdsFGnFGmxn9N
P35TvDAnRkcoYlhVKQKvrG1XcpTyspRg2RmqW+Qhv8tGCjfZG/Wy47E/etR54ThY
WEKUzZecfs1vqL9N3Hqi6Xz8h4/z4kWgkOh0k5oUU2qRw8eMF2mIMSV4m4xQliEd
5rALXXiKgVnPhItDeMlE1vpTBqE510PIwxsZR8g/bRgmZZvOyF9Tcvt7mXNzdBI9
cwz7iB6Sm1NSAifPmEDQPl0SbZ+4w4ARNGyfWZ+iS8+ApWFrTdqp61R/aTMT8JkQ
rfA8VUWjk9+DnnUb4IS0gzVW8gsOTKrjxBo89JkukTDMivT30vOGDRx/POUzU8Af
YXYUVT1In4QWC7KHX2qWycPab0b6ljqLJXpHNa5fAUC9kpn06FqAlfAb2QSft+p4
va98OjOxgT5SDNOOS3chxJY6u3A5GI9b0T/BjXpyV3lVi7RUQAAc7/HAR6O62qru
d7Lev0dnixlsgH150aLd2Lp6BbMuVsD69wypJXqISXPzIq1q2tvIcuv61WqaGYjI
2Gr6e84vYEzz/4+y74xv63wqJZylx67Y1iY0g/U4Plk1TBbfe4HduaFvxlcrK+dE
Tw0ivq6GHJNrow0u1icvzYJRUMWZuuapfhZ81LU85BSOBck2c4auQkGUE1XryOrf
EsFPDqx9dvXOd1B5Kl4OPjpZZsD3IrwoPr9ypPX+aV4sPNONFibsIHPd9m39+rv7
W6ze2B5JAA6vr1He/PRbmnNv/rfMwz36HnybvptBOQY4W7AMqzNZa469+bQTJqww
bAyEwj3LSY11yEFz/MEmRinHZqFHhRNrF7RS26lm++J+6ncf1lgBypOVMijxELqa
f74DytXO8XFuKvz49heSOk2IleSeHphIg95cv8OMUa0fg3W6hqsOQ7QFVdKPg46j
wLohE2gUk2oSyg3A6uyxNG3q6UohrinVQO9CgR4CUsnx8CpiHSMNdwzURzdt8p6U
ahEjVukh5H5u4kqn3sJm1/9Wg2utZ6SSpCI0HvY37Lcc0sLqASLaB+FxssHQSnIl
NMreUfBFzBy4HCvgo9SX++B82p+OKmvHt3SbWzi20xYk7pK011WqlGIRWQyx9DEE
uxKdataU9XKJM2Hi7K6mTtctliQEKMOxgzKYDRbRJE9lxSdO1t1x714F0d2MFFY3
kUjOsTR5Ee+dZA/o2lXb2TvQPFKpBn+FArW08EGOYcTl0BnS2osZFzC4bAhjrtsX
oABpi9DQdqaDdS7qDBBAhAlu4jOErvETVlFc3ySfGn5MudqtDqyBbZub/5DzStNy
pAP6wSEeOFT3oYkOc9uz92kgcy1ql+N+UY0MXxIySw0oqwLXes0eim6Q396/GFsC
g8L5qkTVdUG1+ggNqpL3k0XnbldhJVwKEALaDGs8BzU3zi+mMNZSpbC1kwcqegeE
r6YH5FlsahoUeD/PTwzcntPWouNcdVBGCrt+1gFzCLxLPUXkBnmWCp3FRi2gpfP1
0MmDoIX4JPAe2kf8IsBWu0lgZa+r9KEMG091yo0GF1egSLqjxz1v+EeTTj5P4z9c
F2xK0N/vtlfTkXs3mF+U4LSy9th3diBMDpvEtrUZ+KfzZWdbVTHToSmsalDBUJmP
7Cj8HRZNhsI+UyFww/ZMXIs9J4jdxWTuc9W/FNK9oup3yoHT6urhHRZA5Q1PgJTi
P9sh2KN+532IlCV8wR/Jl6UfnI1m6Sch6jmewYa0PsmwpBRx3T2IcmyJClkv8tTx
rX/O2Bua9t0RtcgCcIzPNz8w3dzW0s7s+Hkj0ictEp+xcLu/VrsLVIDexSNeUbla
34ALsb2oxGjyAWMC4KYmlsMUz6xtUMb7HEQ/7ErxWMeTfPnP9xTRTSH25PagmCLy
YoMoK2YXZ/r9M1lPn8+ErtUj85mZauY5UGOOrKxxq/+MUTbKP4jhulV/ebC8K+Fz
j/m4UF//+8yDSSHtydm964m1ppub0p8vhptVTq0jo8k5xTo7LX+8zhsSHAEMpH4F
ZiZjCCT/lp7U+5Utt7MctcheJY3PRnbmZ0aWrizcdcnU9utqvs1/nBNnRSiKUIgi
Do4d21CPilWLwoTP4DsiYRvrXqDffvSzjI51Mlnfwl1KFILuMJVcMbhvpvU00peT
rLm7ztO6huAVtVLuWWOogSce5J6+4wedQDDsZxvNtETh3bhNZLItC0RQRYpNniU7
bvM8O77fryems/KiOPN8NsBtCdgMY8x6vx+BRhqdlaienO2jpCKPIC7vnLl5ik5Z
30MJ5dIVM4wrnnQSZzrVJo1ibsIZLcQSbyLXy1G17L3ONt8hEj8GZimBjwAhj/sh
oPZxDqBhZ6lYFDFnWcCHrvlDveYkxNpovCqe46d/6YhJDMBY2h3EOYSaLW9ilISo
/9e/VbyZ7uOeGzkfAYWA9y5Pf1V93JP8hpYDV1DdcCeIQefCkXZF51PbW6sQmIcE
eUuma+BOyb+YTij3UiVlqV0wN+fPJPDIywZlT4PUKjdzyrpEWZxdy3pXDALfsAXj
iTOr6M+HbLjChjSKoj/9CrfOkxXM22XSVpKEDd2oBNnZB8b/FOIjNqm2L4bkdaqw
dx+ATzAUZWl5/0DTk4Jzxwq2NeQUnoQ8T2VmR1PSb7G4U7LhMAlnwR4zoehwk7U/
WGSYcZekp3VAcz9YFCsrSklh/S0lAytEWX4AreoryOJGIW5b/eMJ6zR8pTqNRQY7
afTSY5o+8KZIahQmS0d3HBMtc4FhxMTf2YID1pIKLAftSAsW+LBcIGMZUxkU0cNK
sCTix7rJJ80lGEHTZ+dt3VJPkc/sD7BgHxgR91EDxZ3SVWMEVs1iaoc1PS1V9zHG
in+HJg8k7dO2zFOj3u+F+vrU/xka+1q5htmBG9eUWA3+RCYuSh4ch7EjHGwusytt
JF9WFEs2Ftwr29BTO6WTd66ZJXcW6SQqe85FlGniAqpGRqC3grXNw1Y+EQpNEvdA
hh+LwjeViqRc6RbZOHYIpXRrW8FALBa8IHwH/cZK2HYeL30d97h88DO5ZzLWIzSb
oaZmX8B6pNIEGtmkzrYTSRd/8ywKFS9Lcvhq/MOGT6jvX+BLGP/5pt7e0MtaFOAI
3qlhE6pRF9ptCVMTkbMGOmC7KI1LODaeyZCsSCpPyRxSxnzPBgQtFw2HOXYoCXyW
K+myqFJeE4uRym/MdVE/dUhHnhEfAJX22NsdxBoiBjXuH8Suwx3ewSISdQRGFs7u
UXlz3OXonPj9FNo0zAzLRHY081rYciECCx7BUGeFYsU9MEJgpQeEsyPecv/ZKfUd
cx1UqdLpbWlM1+YMyT8yyizzr9k2aARSsccp3Gn7FWniRTluYBk5CpMPuZnMw6Em
YslnUkzyrsCA3w5NX7VHlxRXPoWgB+x2FwrWs0kPEMMKYbLYnFyIgC94upsIf5Ah
L7KCns7V69s9y10MmGoV20bTC98NAWAWkvAd0wZWNsdHBQadbl6bO9Pzqm7+cttw
Z/rla3F2rMlADdYvOrf1LlJv7kvo7E2Mg+X9KxYS4YdMh5blJJGrjt7BVNHCY2eS
WJQ/RbvR5v1k2uxL3QniesnuDFBRWT8bKutJupgWNwS3GxW/NTq9peNzdgoQRk9v
aI+g1tcbXCfeUCCmXKIGGU1lIYevaHWVSGyzcMNWwdLQ0hztv6KLTx/QFOjBmQGh
t2HMLqgg0Jn6ILay1LzlgAwN9oL9i3Qs4il8zPCi0akKyyaN41gfgqdXS5Wr4W5m
JjdXYuDyZ3ZTlMHCET8MRwKPAxiBdIAP72Pbc9xw7OW72eaIPLAJw7mSuF8zfFPr
xT6HlwCkiCWKi9+zb84lgHfef0iVNkn9+8XsiGy+dMffGpiVbPHH9q6GdXTlmyos
II61bV3svnBx2/G4qIvB3ge1+RzVXz1BcF6Ls8mFXgYOXiqMnWtabMV7cZqZoQpL
RXWo3h6ScpDI3K/ZP973TvWfkmGqxRbdZ0YlqwAT2rtyRMdBjBXuog6llJ/UZWN3
iBXUZnWlAcC4n1R/ECmoIG9m63rqkg6td3HmEsK6ucTPadCSwgc7STElXdqi0nR2
x292EjB5vdTdZkkDcU7ZxrW0XvkmffnakEqDiFK3iSsUtlzlvKALce1AzWw5SLU6
ES0ZNvxjzh+wxiXxfccQuv70/aTsLRCbT03NJw8I/6RZ/iC9ghteAax6sQ8vwN7D
QuoTjkmdt0YpuIUrNaB7axDtXle8RlXAM87DdH5rVuYG0cthPjgYLW0ch0Ah09JW
+GS62f1/0qRNkCbDFQk+SB1ovmWKXkWqRjb8m7jQ9PNT7R8u7AN0VRK+xDGLMVfn
KKj8eX5bF071CxY/vhvILusA14NVTz1TzLNXnt42yTn73acHXOmYlSzNbPOXx282
Bfra+XNEY05CKGk5qLETll6By3BYopEtDc3TjGOccASzPjxAIh1EP40ZxEJJbd/f
+vL6gvCxWZQyFBIn7zrmnED5xEBtgxARBKyeNWj7mtpp9LPguoRLbHzW5gsG8wFj
GJIsltbYODVqT4iZAbEF7/1ZD4AIN+6JXzmY6bRh0YNAVSUQAD0Y8NN5Ls9CiSdx
c0zChAbe0hcXHlSODbtiFfzr0MacNzhjLW5IwCq8Ao99iubfBFo9rBLZoUThsHkR
c4S4ACx9cWkl/s/PSJ2MyLYBPR1iiHYq61Ca+qXKSBP1/eHTCyRfZWaYWqgaLN+8
HYcplbvZt0XJzplOQ/jypIzlROxpg5OWc8LY9/SmhHQGOn5EVZ9/gax1fgkCqr5D
UhND8er5N/zOuSuf6cmzUuLoPApKUDAcGdk+agq8ekszO63VtYhhk2c7RY+fiHO0
QihadghqryQlR8bqKkA3z7jRNnp0iAia//SNIiuf/bWDJ5TnrXHcQ2lj15qVzH2R
c1240KwIPZePBpOExo3FVQ9M2myLqUXgU0zJCm/vbMSyi+WMLhPKVPCBa7uNIE1/
N+JLEV0T7j9AisiVvZ8Tm/csCce39AvIJBP0mh6c22oPrkoCH+BohFS9y93g+3O/
CoRZIssijl4zJ7HUthQb6uMSEzFn6mU9KrJmtSRbaiSU9ekZbxW5CAavcOc7xLOt
0nPpBBI5RslFCJmHqpLHbPNucErQwGwmP1VygNDoDRprhze6ofWoBun8i7WZFdjg
3S+KNRiesyqP32kzMvt7rCaZJumlzLCmvt34eIqKuk6IRnDZPMEWTe7DKgUCMD3H
r9CXTalnXjLfBkQncjDyWN0Y/gTyt6aj2YSnLKPN646BGq56e91a0j3oVW3zZJNa
MZDkC8OjdQGEEprkDK+X8NpGgdsL79WAZDbQqWXfY3lPNDhi9O20nyIxyUhdRHDH
kgOTQrPLZ8nUE/CeAheKPXLqqvNK9zYHWgUuiZlXitwcOFn3wCeLBuwr8DFOuzRy
amYG+GsEZcuu8MP3i+cDmabLi6Zp4E1sZDao0KlOJ9nZjNoGBnh3yFOdc6t/PGxa
97Q1R+uvDRL+I9JnJ9WCAJZ3QcN4PmKKGHqXnPrdHjcq5JtWAiliyMwdWxHHq97A
+aHu6iAjl0YYUWOuRadxA6rA/1vdnhvrQekKYAcSVoLtFTTTVGiz/iFmCP7kdoE4
dj9eMpEzjgGnjZ5eZ1LlNO5fQUgF/SCS+CnQ4BwzlhfZUgrtP63FLI0pvltbQ1mf
zYw++/DpyLI8V/98Oq7H5o382+14s4yeabClMkAOMu604XBrtzRszPbCFyL5RHH4
2GKNbLsOSgwpVpKGC2ZPiCHcPTj3jjpzQUPzMey90HmEYvJ0rzcvbdZiQYRAzSJ8
PbOObySgBG9xD+HirF50ACLQz/uEbJpiUsvVJLXIu4u5zeryERa3IfHEMJqEc38x
+BYNIra+m4z0WBbGXa8kMULPfCddYbDUypDBx3ydHJuzQ8w6tTw8DrFYoScDdz2a
E2QlEMiDPRGmiDSNFU8RrdwBUijjoqga3N3HK39Q+FdKPfWhvpZTTLoKLG2VJXAe
rMLYdTTM/i3IJjrw+EH3Z4LR6duq8qSStXKUOnlrkNq96dMxGdMbO8Y+oNQ3JzmB
Uaxc/0ZTI7jFcu77S5K3pt96taJ1j8Tj6OXhLRvq6lI4tivWGPg0cNUSTSi4uLqx
gqQglrnKPtim5gesrWykhNf3l4xULOk9NEf0DkA02NdaYL0CB460D2Ail5Teavtw
8TEg0fvj1xMFee4RAqjGiusXGkJbCDWbOkEEwNfIhRX47DpGQEhpg8KqyL6GnroG
aw+6EGse3pWuvN4CuXszqC7DJS9Ipag1gPXfm5asc6l9nv6IipHvVlgL+sEr5fIZ
LjT81bLX8lyAsmvwrg/eN4ob2rDkzQxoCEzJBThHHJJ3THP+9BioRtXn02tjoRkF
fIJDixd2E6daDmmuqey44kWCarg8LhSEbai/tj7zQ+odu/PnPD0frrwxEgOL6EsW
fmdo9HkVtTzpFQxDXKhP5RN1tcCBjXqqpfMHddQc+fcTGT5Xx5F1S5uBVyqzNN1j
c4CgpRbqeIDvaQ91o/hKTe3TRyh3LB8wgTt5L6YAWkyzYABrEqqYDo0zM3r+73gv
VUG+FOq5U2IcpaVa11icjUi9p0i9CyU5F8n5twp3e/4xf5yJHg8zhSEgw/FHiRZ9
o/qohp7h8HP/OdbosPswYdjWH9S8wEpic2ukliHRTyXVzEV0Nl43Kzd8Y2wItiRH
NJgr4IiwMu36QiO7JBHbm3guarch5VLNOSFyv3PGSrDqtyTLHNntz8rOvSl0f/hj
Iu4Svpw3ZuKrzcfsxgAjAq3Zx9Ic0RRh5iL//vWUuL+toLr0BDCXxhFzmZ4hycKJ
I8dHLqJgBzpqspZ5dg2PO3/SZUqG5YosFXa+yBDrzBesFE/7co9eQcjrRzOFzNbs
zcpJWpqbhN73pYn0ZyLrdP5qYxiege3kMKl4oRYP7goapqgICGDjUVhZEd+uaz2F
ZrRlf8mmqb0Gr92ARhMzwgAyNqcZOmYNzOvBwuJNex1XWWXsTRTAurQoFU8SfbFY
6zCvmwoEhjwSCjixk8r2BG7jAesYpzuJm4wFHyifLVkqTEVjVub6DhzWs8WIC1dT
qLMGH66+p8QDxTtn271FwGYQVieFvQS/sMnKH2vTJrWYJbfaL8VceNr9+RZxEgBD
BHcDcQzq9BJGYBMv0ZwaSbLjMd4ncWUfhSxUYFyZE5cHkgp2VlOrFU9eLrrLjHWG
BGs6utbxcNB8D/hVvgwTJdA6kwEdP85jv+WoaDJMsWtw7em1H9kxWbYKtrGqD2+x
5ntXdeqqt1lCkLd+/iDzoMwpPXh6JvmpDwLda+iSiDocJ7Iz6xlabdeOAWLAkE1s
DRmmH0UUJXczmfiqu2dKGxIHMFRCmvOfXdrQ31gb0RBWBWIef/HVlXPGLztBR+HO
Imseo5Ga5oO6pnaYnllwOh+CjyIQKlFOuhDjEfT5YHtH1QPl2cmxlo8FFDlFNhmP
/LzBwXkWksXKFeiOjFxOB7NbMJ307tpJeozSTC/3/wxLp+xLlKYeGeYTyiAA61wC
PnvAdepOmwkE6QsBarzdTYwjuwSLsa/OU9W8cE0gm6w6RR0DB637f8wxcRnsSkwR
FgzElNMP0IjhQG9yOHE5onHdevxwjeqQ+LecH7g+Tu2mZHsPud31v0QGW0jYtqDd
yxnnG8x+IHKFpBfRmjnoKCW0L/xqjQizsmpU2XcIecj06f53PGDZatLf8HTZubkk
TVZNnCIkNP36JVH/nlO8tR0kHWD3bUAHM+yDRqPIyo+iET8iPCzDcrh+Wuh0h79B
vRx8s3aSIeR+k1EHCNUzzh/xh+AtQx/rSOU1hpOqLde2Qqhem5eJaeYXD0XxLULP
h8rxpvKF9a3do8atNJU7C7IYeHTfoIcQQ+gOSJ3acPo1QnoG18GGYyU6zwu9GnUg
J+GOTGW3jeAolraMNb15Tepq6p5+vSui81WxiF4MjrQ4xqS9befNTSAPWmOHwhWn
BGlanydt68MDMnl266DrUF1WCpHVZo5tE2ChBDRgo8CKXMhnJMK4UqXGI1EnL9lt
YzKNaDpbCY+hyEAYMkJSE0/BexFGwZxt1+gvLvgyFJj8C9aunkCkC1IM+CvHTzLT
ZgrUDtWDkc4kzyerjzqITHIP5Kps5uBsF8PWUigrsSaG8nKNLsuFRxFCZ5Y65wVD
0bDLHg8yYfkoRqEUVkwIPj7Tu5mWF6sfBvIeU2tcJ+8sZgNCppxtfkxS38uGnd/G
g2zEIvbkuPqce8+4igxmHBWvC7FvcYO+yCfk8yagBzPwq1cXvAZWZBx34a3ugzpr
LrTg4qVE+i7Alx6BlVt1cJQocUMpKsSHT9na7PaEj5dlurW4Dk1so9JAW2PWQuuh
UCy5VnsGsmg84Oiv20m6Ueen/KL7ZCWWc1r9vsLiJFEwgIhQXuupg1i+J5f3lrh7
eqbkTE7TIKK3mu5gMpo/ribYYYBYCWth8jvbfKNI/6yCBs7ulvjalKPYemTawCNW
/K+1alPuOO9R2FxdAVqVwUjDHXPZPsZQav28WFghGQWz5SEmQDFe93QocSIiG+pz
wTB9hv+AlAfqrIP9pE6uhKYYVuSx3i5OEfSr4S9giNmsmZfIlp0ahErabAPWvXnz
V0oy+J8dDmNL9nQ//nEnUhUGN5MC1npcGN+C6IJPYjcRp1MEB2sUo0oC7klFdOPc
NvtHm36HXKNCAu4SqyJvJwcHulDz6YCtBpqxBOZJN45/FsYFG0+bxhjzWt5oulrD
NfNVnsTjtllOEnKupP2sv70rbVLPdIMFB3utGM8W5+RG2kty5LPJwvhPY9Q5uv6P
xM8ioxxUhQvvd2SIeMNHgHXklBw/tP+qPlXIumHsiUzptRVfMeECXv/7h3FFdp2T
4gtwbXR/NrzWGM7B+fq1EghSkDNlahJzKK1/OTumrzvhlmgfsAAgZmDho45X9ErD
BpKeckImnLcpkxBkIOtr6XScWkXLImvCEEmVrcvRCSqEnByWyhMITGLH4YDAR++Q
1Ir5hICHHYBP3ddVgBn43C1jRvuNhi027uixZNPZ5mhpZFbdVxWvAL2tgxHxTRZ9
MfuLnWuJIoTK8DM97PnP65wG2jCYhy+9I7lumpzCFtreqf2FEZ3nHiJN5h8z4bwA
XEf+d9vD8Bm23fMc/K+DCm8YF8bDP0ra6aC53kfW3tkmSzeG4XUU82MAU0N5WA+5
6AlpBaMf+QaQHiM2yaijwF6GoowCnVawtEOJ4hWUEE8/R/LLQFW3C57PZBsbxbSO
LesSV2Bn9oLI7U6tFm10m0ZPNiXOhtTaoD2NshchjaZ4DbLh7eUtw5vjlcON3K58
pf8V0IQ74B/qDLhwhGXfFHIRkZoNzm5KQfyoSzkQKVB6AX7mfzXOtLSqgmTsPxvX
uKETQCl1LNrgIo6bUwhbbD7/hLmX3G96rhdwtRHINP8HpNea1vxk0GPa/CRTS3w7
YQ7jgTa61dpbWbPP5xxw2hjpVyhY45/Hafqoheu4kwjsMNQlwsk1K75rrFb4yaZF
5EQ6spo/3wJQn9GoVHTPSR9poDaaA862DsZ8x0mO8+foa+7PtrlXXrtvVC68q4cK
YH8iKazpZyn1l4/WWomwy8Tg17K7AsivK4/qQH9Lesi0O4IhNZ4eOvQNlSv/3ApV
0mCTUsEVOQ5YzLny8mS6sFIXO7cx652QzCuMNWi4G5Oi5Bq2X8/1HLKHAcVE/A5I
dz3O0coIFXusGSi6ramP5DtEuOPsF2CewMQ9wbwD8b/I5he8oq2fGpTxAjW05tGY
gtO2dV6sihTAQt7VP2RszNVM6+Ui0fPKKAHO15qchzHce8tw2hbWSMAPk8p10J98
SK4mW7hcB+5Gw63L/Jq7waPzNb9F1JAnAv7QYhgWzvRGBRuCoCtuOsRXZOAgjY5b
AplG7d6aMmO2fisLnq/4RtmbW/NT7GyK7uX5EVJqsVkxEgo4XPErjMQ26Ke+KWuJ
O/0KEXh7pHtxjEablbOAtUzTRzNYyfiiOYwVCaSg/TCA/Uf6+sIA1GtHKpPVQniw
N5Idi6HgL78qfscqK06zKKBgFls/8B6wordT/RrAxHblHLNRoMQMBsU8UYFNFR51
a3tEE6eleap5zZs4Ifu3xMmbrds+N5NiJRDGNCZX7Xqw/ECoYRAmporDEtyiRFrE
V0DSUWofW+32jVMiHy/uNT6YHvVuX+H+z5CNZ9yJa1dzYomx8iIup+Dr9QVV+TQ7
Deg037HS2ujlF5QH6YuMikdaojMLBGVHETieXol3MEQAcmTIKFHr1wtuVK9U1NXZ
4m8JxgiTM7kB9szF4q5PFt0xoCvrhRNVMZvkLw/q7MmNYYAp2SNhQrZSf0Ncf8mb
IvvOsYl2WaLZTQuBj5fB994rYWOJUm3a/JVEnRkqXrK2RIAK7RRgtKyg1qTUXAPy
iNxQju538Bl5oFW88tiSkbo/qJUvec2HoKWg185JhDcweN8GM9p/3U9gtLSx4afN
5EA2f+zclPxQq6xfE2vXISI9vf5kbNtA1weyo61lAgKfVkaF1GYAXCi3fMVT2HJL
BlIwbY/F8yUp1AaL1QhVNCc6LvoliqRy0T/NVjCgkzAyGQtrNUx0AmUgj1rTO3Q9
h/I+Kl3Jj9vTxc08bN2g4WkBgjAjE1rEzk7HT1RTNtFqg5A1AGP7n5spK06221tV
JpOfoP+tzS1LqbHU2vzNJnZtG/PDMhS2DK51x2sjo8v9yxWtdpKnhGxMNZX+XtPB
URSyBx/8ByQCb8ghzlMVbAP+2H0ZlIVzpg4C4N4M4grZe88M/T1kiVnQaL4exB+1
dBpxalCZdiH4OPznA17kgoKMw1X6n/6paYW/r8DIxrAi1l0/3pwER5mjig01Wn0h
ynfh9LeGm8Lb67II4Vk2SrGvqFbfYa/ZwydWrzpvnazyJkWoV25mI//Yh2ghrlow
JQMjn+0xOZg1/Tpny/pY8PkRdA1rHUj2y5qPzK23i5sPHelp9k0bC8+mnEyeFs/S
bECA1jRY+P/1pZfrmV04ullGaL9yF0InrIA8ly2y3+OsGwyu6wmFS54yw7wr4C2o
jH5mP+3IMQXFHl+fzGwDyHFlc2h4Yz7epJP1xEbW48s1nINjWWtTmfd/LKEE1QXS
+REzZapQdInRRwAZC76296OyaC7u471g3eNQUsmMp0M6k4o8Zm8k/p0DeeCOTZip
I0MRiiW8IiEtPfOWh6QTKIaJN4tny0wny33ChVHtH4hUv5J7BFYqYg8mki+Bduj7
FChiwbMUkUksDiUgp/FsIBhtNbZmfTc3qbniWxuvJOxBVAqW6wx73t1PZ03nQuxF
bw3j/Um7/Fy2XLXmTlaqQia5S4St7rQjB8H+/CvFe4jHdTYd3JmNYatP+Z+843E9
jATTSGUv2oVDsQFOyaZF4KZlu3VelxSt5uso7dMiXBFJBs8/HgTBm65NEUbvf5xH
9UfVVUHTL3yZQpakNRlDfXtCB9Sd+c/WkoahONOzCjVAQKp2KkFMD2FgaTw9Ql+c
/pGcXBhBaCRIsEuUT+PO/H091RYjyPjg8TMV4sL+NurzwqD87lQCKKmjqulOFH5q
Juad2RNiK5gBRivbHDyQmFcBbZ3A2/CbM6+neRf4Utw8Nl7yx3Et0gneZbUW8ToU
/tyQt77VQ6cnkUw5MQGbCuX6wLiZEO3q/xQMHZ44a+zi43bdT9J2Gv5ZUKQ4sHC3
Dp0ZmgGKMum/tn7c0H8fTKEBHBpmurEdhXFUPuhTAAKEqJi6FAxJpKzSkNFgNBEX
tH/0BlPZUSY0p1ehu8BXpWLQuSMebik4RJIQ5ksh/V3qvefPKUz2plmnO+ZjgKBr
3LwsTEAkf6v0cR423GdZTPyGEqKG/XsOCYBktrpKuox3aSSL495xB7jIWmIyD6qb
ZzouuTHJVNwCGi/IPzfsZKRWPfstVc4Ztu9dudtLYFWl9DlmMQ6kMGPJOaQ6ppHr
VqKF6FonpttDPoKOxQyndHArDp9dM661Zbjrz1lot1vYJNY9S8xca1WDKy+6WD+p
tH/pwb49YXpu0VTiQ5xOjj5sOrsBN3ORAhUnPtZVOCcI009F3hAJH7/FVN7WlKQW
97TtFr1NkDkLrSlMolv5KgvuqI8dl2fSHkR37mVitu3Wty+/yqr7l8O0S0NYcso4
kJxQ9o+LrJ5mdcLy1kuAPGS3kWuPb80zv6favyyPY5rLDayXlRCXhC0oEjpQYkgr
lnrJnj2gTu1dHX/lt2Ar8iomX/gGc7+72q/ygBjMha62kya08aaqZddISuio9+IP
G6qYYeoO+bqffqctbWvOZSsfNEyNX9aaRs7shWbriPwTB/tkdE5W0McHAx/yC/A7
Ofl3Ta5lufjG/8s3HaZVKsZrZqBGSjVNXXJ8zdxpX0Qp5haA+tl2DEoI0Z0LQRUA
Ux1iZMG0SGyXfZ6kPhYW64HVGVaIsBNyjugxgE1f2smaS7XTqiZ62OEFQJ5UhsSg
qHwl77UYW6jPZX75LAhYdDDMM72reUF/GCqwkHMCCEME0udrOcCqOy45i2FM41PW
/gIp0pzMAN6XXt2GHc+F6/7hkm7gxYKapFiA8fYVY2iloIr/syfDPHnGsSyh2QYx
TD7Z6VjuDl6A9tSPCs8oAQKfaSAddI0QsFMWinelikhxRM4M17cIEK8yvGfMubRJ
WBtDqlYdZMuXPOe2XMREzBG2MGtSeDKZsttqgPddsVe4OIuUhYS1ZM7VAxBP3rIW
4qBIHBSyK6o4bUyvBNW+j2BcXv/2of/ufUTeihvPFV0SkKd13kESfJ1/O0bmLH1F
FPzVpMivrkdFPEl4cUT7S9aJE+CMXt8wiTD56OOiNMMaesj/7ejEXjOAHuqho2vR
F7F1kvkU2RxlE6YS/KLuT6Cfv4UDLILqB2OXFWX4I846Sr7HuXqrYykI6g+yKRoG
0wDcWbdXft8/DHbZ33V3zigPnaSaUodekSPdIrjkVDf5L9fW9lOCe9w6i1rqyN3i
2y5wDQ75WnsnBjdx6YEC7w+X7APHFhHjxQt/fS/0OTL9S7sbmBWAYV0YC9h9V2sN
x5oH9+tJCtuNnJbDLetb/OHPUnaHNXfyzVeGuWtZYyGCScudLIqiRsq+3sAKf5Qh
uU6AaNWxhHzarXrlwh5vNvzZG39YtnFSIMAlc/7l2T4Hhu8ZN8BRl4Ia9JdO5i8X
3JBQmLT0GAql7A01KziXdi2OczqkPIPN7mMcirzOZmOZZOG0tPSFv6dKHC1m6zC+
98l+7Xkq3hge4m+89nhd8t3YJHVPABIB6XQGZXaAihXwZWpESwlB/8oagMtijDPT
Tv+EO/JlmiogCt3bLxtpYDG7xzlYNHJB9KRA7duW5UnIsdvNOUo6kVanA9LLyeYj
VU0fBdtSPmx8pSCp4SHzGTMrLXnEFjk0q8M9BObXYKdCTVnnj8I5GCmvSo2DhWxA
oCigp0XZIYmsBXgFwVskAnW0mAswuDZHQj+G3B8/Frf+hzC81JM6I1dZlF5Z+CpS
UE02WWBoLr+n4fbRIcvJZDjEFjB0qfZIN5T/gs8AWrMQ+BuBhwXe2qJ4I+DEan1L
vydF1vCx2CVIIYrkpvzYhoUPvZABPMUTc7beSVIv9NBP23udCGaM74sUDBICCsdL
q6btScAL2TLK//EjjOIs1ku6yxCQqpq3Lv7Tenkmdu31kW73cAnq4F7PZaLfC1G7
2qWH1TkjcZ9OhNWsSQjDCo7zl1W/LyBslJWNduS5gRDk+/0V7b1glLo4Td+cV/JZ
Lmay/mAexBm/1A2CJKX8yFEcrlCpMUH1lc6/KaeVErOhbcxy5aoXo+irCPZsFVdL
J5TnsVC9RwLM62xOV6zsRnhHPPoe26SwNnnvkNJZK5bdlqDKcgTWaUPLMf8wRqw4
+blX9TQUIUcNi9ETZ84Jj0riX5p49w6mdXISrt17T7stIR/KZIh42qcHrUZayfdz
d/G57HTGTT3CBbWMudqrlSc/gn6gNrOCQ8oWjcvUDq2feTEkuTK5QFoj824pKFhy
d5a2uM4D1wd1CItofVTStWKPw1ijC6VL0RCDeOxj9M5ZeC1wvOfEUP6pgk5fNwkt
yvS1EH/rHowFt5IlAaK6IYS1xahFI1RVe+5kM9pomyx4Dur0Kly6oSHTlGedCbvY
EoPek0v4gVmhKlgkxPiMTylujUUzj+bfCcy1aHFGlZic5I15990nUngwi2yBUGgM
qbFdZUumHF1MpyZGgs9LHN+UInQhXc4DJv+D3CbfpZPvP9o7a7gAjReh43b8fGtp
kW+g+rR1cPCU1ZwD/ZCIWW0NDfbQwsmMflMwRO4ZTs3iZLjeuXwnx/YRE6X51YV5
97v+apCBb21pG0syrDQEbQMQQFIPaG6WypQ1uokaGReO5NDkjY6aiwPBFDiJYX03
ATDvACXV0p+hDwKvaVrO1Ydqdd8CL1aGbf52tLP/6B3EzX2VVfmXNYyYbxKnJNdT
PIO1uB1lykiOh+EVuYrtUmJRkmBBoQPphSUI3OHQqGy5d8m06L4eUPEXqIU41A4b
b0KgiAHSrLzQVN+GjCGr+naUCuwzQUY+vc6o+mTWYX0Xu3733c2nDiYrWxTezDAj
L9S+WI6rGdVMwcjCGBbWLrBwUEj3izQBn443l7scTxONlQmU+kh1FrhOlDYZNKuF
sT1hwM9LN2UGP57Nr20J/qCjYiYG8IVydfBIiPCgCqU30OU1HVH/DSiHX0pLOAoR
oVukfgu2JWvvNXZSa1VpwNZl+ICpWbfZcrEnlr/fNVpljRoU8Xtq7YGcn9PiQsxN
suSqXnJ17rDKeXiUJIzn+HXlf6Pgo4CrtIPUPe7QVdANmijvEcwuHDVWVNU2s7OZ
ax2p49Vk6L0Vghd16gdd4h2zjRKbg3NOJ6nOi3EUg6V04HBQBLoGB9dxaolsjHCI
4WCQLosJDGCMgetLQyWuH2ghEMoKMQ4grGcpzB9NXjwg27HgJ+qA2d8oG73ldPh1
zrDgbaws2y+gVULfQs4cjZrTlq8s+8RU6ppy/A1x6nGar+gxUKBzqYg7sBq9oYo0
3Oehnl6oyYsJBLCdrTFkHAwEDqFfomnCUu+Ybs/hHTGMIASg+IrdFAc7DhvkpsPC
BAdNq9NKDkD9BzwVL94Nb3FP2ZGP72cv+M3v6r8dR4vQg/SoerHcwWareS5hpRU1
C2XIplumcEFh1Dib9LwgFOK+PB9wAtxCgArbkHdYtDjQ5XpkrmLrVbcaZ6BeFsXz
5uWXVrwLJLDUzXLjAMNSKodBOQ9mm8rgyPwgrowPjpnURcZfNcboLynwU/IHVglm
I0QBAzIP9eLMPWDusJQrdDfyRapzQP0niiJIfnMP7eu/5pPN8j45viVRHa6zEIsZ
wwc9udMk7p0B48aDvYjdWfPqLOlTa2uY+s5OD/dowhRgr3LRkhha4XcqGOd+esNB
xkzsUTcmYtviI+njT1x3kuGoYzh9WPbmSNftJjRxXEOx3zjgNLr+vaxGqRVrZH9K
HEWeu4JU3fbjrlj5nM7Z3SUJ8hO2FmuIiZgE+KuuCXi36tw8oGwCeJqc4Ip9hus2
rfY6oiiJwaLYzGivAN+5YbgPCogDWpNKUTQWntGRTTWIaKFeJtA8PqwyyEolDtyo
hfQnwxIbgIjJVK2Px7HADayA0h/MNFBOpOlECZqu6m9RBFQCx1Ep4b2HDlSDtAm0
mfjk5Ll3A7wgg4gU2QonKwjawfb7ew4suEflgZsbALm2aHTJq9C8EgjQBiEVvz6i
Mex8Gvo3ZYbalB24hfmItxnZeuvBsMAgqr2DFuFWiWL6s+IXMe7MPwuZwt1likRr
8NTL5xjKIvg2LWwG50HxS9ulqZYjILxIiiUNUxz1tYjYbbpXho3iM2iuaQGFslJA
clXvSDA7U5nGKrQPlS4nMXCxMHRvAk5odOILYXbJDaJ5QmvIuV2xi0CFFt9BaQ4w
M/loA/mdHHE25+NFxfwGQXolw4TvuQRF33WHstTvGYohf4PU1rnt/42oSb8EBMj2
Zo0Y9F4QRbfQaqWGj53j9N5nac72ZsboatQ8F3kfnSiosUl7Pd3dwpiYdwUF8lms
yc2FoxjnOBqqc+r2kX2o+AhQiJVe3jLtvkJwTe3U+3aI7a2hHkhOcoJ67oPBaBoM
ugjY4ddiFToez25CbkTcASfMbLXTG/oplzxAzMNWZKjw97MX6nfUiDXMMDIGqG4v
Jz7eSlXz2EqwAhJGLPcmuZb9R+8x8yoiRgPkIhceluaNf5y6lQhkbvRHPhBHsviH
Uu2kh+H+JEC7lpHQ7NBIeYrsOC2ifuiIor68GAWISRhDLdfYolr75VOxGCU+fWT4
JVGGPeOPu3p6SPvPBrKVaH4MCZcklkp2bi0xLifOFq4jYEGqezYwjfygEZSPGKFF
B+R1yuHzxQnfJnRJKMVVu3IhNBaM2Fi4QazlGyGfPkukDn58LQf/paBbE/bVQv9l
DOp88DCgVfdJD4g/eNbFdHJQwn+YTA7F270XeBjYGachykc/YF0891FOAMAGV/OX
koTpL0Kh48UhleSq3qfyN0Xci7MOmzHNu7hHuj4nVuk9Lwmo52BFOHYdvalHg8ov
Y3C1tZnzoM5PpKeR2VT6UgrBe3L9+vjhO8tFL8ML8WtjrZq24JUwt404Nv6jmUfe
kfFTg5z5OL0NnNOPWOz/hNu+LwDPYdjoSRmRf41yMDA773feRq3wUKbg5oPL18mC
C1WDP+yJ/Nd6BwWn2fgftBDT7yMWYk5SlMgp2seBQOAvXRKEflTJLlSVH2gfD1od
ihUTDbjaIH5+eo18gfp932/epQ8BIIA4DvXt02DPA8wr71c2vXELcwKa1RCN8YZj
MvE/B4vOUzkPCWzX7p1z3OBuSpGAWF+WnxEIF0menJB7wxjZSWeLshixGDPPq73G
8Psqc3AlqE3RvDxSF2RP/1aNijFCOUSqBxVtp/Hz/MyxUI6nJXLDPvNWEHm+XUj0
CjxgmHGUM19sC0IlOuoNtdW5CMl0YTk6h8aeGYFtsjtbBpKlady0BWDf3K+vjFsC
h7nWHeTBImapY0NEj4CBLeUX2cS/dBNwaoGcFUDLazXNdllxUnlap3Q4LPrdqzVi
I6eMs95bSCv6XFhEceqtTwGcTALTET5gUwKK9A9praYINcQgVWIP39M9K+dpaJRZ
16I94a8FxbXyhh89F/+yAuadI+Bdul0nD7sLCKJEeUwJemHXIGmGo0KNeBhKmYfM
K1YrRdWyLNwvZBZEZqGRcfosoFlVg/04Ith5D2SZCMrSTpvzkz8Zgc92Me2+/f4t
5p7npjerZJsRbT+jx/EluHf6OTupPxKh5+JzWAiJrQ3Qx2n8EAAfRUf9vn4D1q6E
9vTw5esY9nRf/NDO+2WEsbmQbrVmipfVccQldb7Ma18gF1Gj5HuMs4q5JAuA8oW1
arA2mGXpJAliF1cUz90GR3jO+uWyWD0XyUFuNOtj4sHEN2GhUM49wVAvc0tJ/XCq
W5YJuylKX250WaR6SXhhN1C7s7Ci6N5HsZ3YYKa4ORf0Id2OBtV5gOl2AR6p/Dqi
+YC8fFp4Zjz/oJ9uMwLQqpKcDWRU3A8ingEMU7vMY6xdgUarqKNw57vMIm27Z7eI
5WLVNQF6hvYNvUl8LqG8cPJjKZ7gQ9199D5X++/oB+pZcX7ipL4dlYhQG35jyiBx
1rUSRHYljE36JrEYYYhtVyTF49czS43WR+erxemru8rSMGodOxhcQzj4ExLZb4w4
HoevQQL39RpmHw2aPsOtahV1d/BiGbVZEw8GCZfWciwLLpwfkMwmtZ4zQE4lMEr5
ae3XJnVWOerexAva/6lFr0OKOu+PUUGW8bJxRo9DaZQ0XMyn2regIytaDUMLL5T4
sI23HHSiQwmN2k0F0ADxXDNh7VxGjBtpeiB7viAS6DpE+E7jvNHHlWK1twxIIozx
BAH3Pfy7kIQs35/sn2e7h9Sv/SAormPTBVxz93tSMowQX/UdHkjtd/dhxIbbhOwA
e/3lQ9cRD6Ae3nmKXSpk6vQf0t7p9+vCXXxanlmjuza5GR8j3OyQLHw0bFR5xVRw
z/D2vQ9+HAeFMngzRpZu/ZFKCc0zPGIekHaRqeHez3xxAqBkph2Sf3djZDk2b9WO
5B/VXs+J6iA/KAtani2Py6z7Fx0AVYZwcjWG4gryHGZFqLayOvj7ja7P9rX2Wex+
5MCuTcS5qqZWPNksRbTHaljBEAb7amzd+bZx5U8mr0bV7tzgdS3F/OLkhcJdnMXD
KmmxWZr5vUgjtHplAKpaOF9o991X4Uqg0sPnR4uRNixnoZw4mNGC3SH74H4vEOKz
nRlkz5scLqjCCAX+JsW3PCN0EnFtaOXgyByoZjXQE5YFMODGOpobjk7OhWq4S13W
+vfX+x9/IkNzdcG0gLhtFDy4Gm1wP3fqymEwbOWpoPO15vJDtrtC0cIQwAwpcd5Q
b06l2jLovlIg4pCCpzOTLnksadJ2n7vNi9wROluf9IZZuUQ2TIhSaJYOqvfPg+gc
+AX2X2KMQuRjNZAOMbb6aJo95nX/J6MCqRGBVjopEw4QaUdXNd/7GOl3c5xqfo8C
VmSz+R+RYjYI2EIdGR063eniQoyaQfTXFebRc25Nc1qIVCnCLd3WlU12bdDhgXKL
6fLkxWn+AD9aPefa509j65hBSHVyr18U5ChssxIxtwUxxHOOWNYVDrLxRPx7vyh2
VMaj72FaHTQjgF2IQQt7cE6UtPUk1Aq38+BwKwWTLCm58WOrDR6beujmInxOPFBB
3VfeuiY7gUJklFqP0HevkIDFgnHEC4D6dyktVVxnylLMkJ/QhQi9j/HlnrxKr4uX
ArXHxmNLK/T/t1pqppnXbCjRTspukWJu92GYUH5F2jSorTeSAuanqb25+WXUd5Ua
BclxhQgCxoJ7k2/P4VT1VpK5xvhaFGUgO9P6GeWyhcR6nMhbnSNBSTcTVK41uUYW
Gg+OHyyBwiMQYH6SO99SINBj8jqr3p/H6j10A0p/13bF9qzkYBQYnLblhi+9FHwD
hpmPKUnI9nFwUxT454OIpfaqpZVBs/KmAYUgfwny85zK5bCKMfkhhXpoBeYkFG87
luQ5XsDz9jKGOei8axbOyNIVEWt8reppdO6Dl2N4X5n/7fjNON6EDsggnDlUgT+7
kXBlPiqEm/3Iceq4YF+wI7IZuNkxwptoE3DJfNzNP1+SFCvU/lrg157tACw6he84
NMr9LuEsbYoJfB1JdaW3TSR9Etjrr+RhycF7VztWD/DAlNYTYW9tV39l+TryNGNg
OTGLVKXKfIo9ONLLq2ZkvJm+nDCA9lsoHf+oXKFbSKZpr1P+jVcOdle33+BieiIg
SoyIgO9U3cjDbJnOqe/c3/IgtxvmfuvGTJ9YREi88OEcc84prv5ZBCytnuz1YcZB
Pcx9Pkmp+KCqSEjS15zEZu3+SLyedcugZ5gJqgTncx9fHs34MJ8hnJW/ks9FcYZ1
f2X7s7iRkwHg3gKW7+/vB5RXMSAwFo56jQ9KzzHdgHcaEZV9XLfmkWudI79aCtW7
E3dhnvlN8hbpI1K54f3tDUCjSSQApOD4Qu7KfkySUfTHaMf6JbZp0HmeajYPjS3d
VxggSVGTaNQKKOMxFf1TklkfuHjs2kojJ1oFwCXhNDFBkDmYWTgbfem0Lry8MuZt
cm/E7yJLCgMCEjby2PJ/HCZvHPpi2z62Mfr2CHvlkk8xdz9LpXqMN4/21hLRLUnb
Bx8vdWPvUQ6Bw94E7umhX+OxFL0BTzRh2fzgU5rVKwQh9gTJu/iJ4LXfBCpo3CSD
JLpEFExa2HxA2UqqTPXwkeSoPA7f/FWNfZ8x3Dcuez4XX2B9cnuw/dY4gIrDHGl9
KvqPO8JMGEOJvzDEFYI7+UUCWDbIqhqsBP8V1ApypPkZo2yLCtxPoEQWm1GZVpa/
bIFfDayDkgyvMR/sxva94ZMODcWclN+ZfLb4i+7pvrAua2rZCslLdmoZoNkoy8iw
ejCfsgMGXNZvZsPMTire3caTRPPfGpSvq8DnUXrtlCY41NvT+gFVYawb9WOZT2vw
uZPuZZslPNInAWSKAwCHa7Q+qb6I67yiKSEyqhBPuOtT21AiPIt1JzN4JO+amV5C
QgsF1DSqoimBqvbn2zqqIIIfIMOJYsC/IjVH7Tb0k9VYEU6INIKAx19TZRkWzgcG
GfDodJ08J6OtIMwlj32VpN/qwZ823yy8hHO8nrsrnOu9Wd56V66an+vprdCnp1uJ
ld23QXVVmBCMolvbyi25hWNTHcUbyAns6Svg7T+oAstvo0p54aj01MwpTXBt6XZ0
Gw0YExg7r/0irvVAhJ0cMZhxP+bpq+z1THhppu/uLpTktodmh4L4PpkNMrIfIdBY
yIPkJRPXK0vEPUjcMZnJDolbivIkPAw7kMkGGfHpe2DB6G6nZjQrCvOe/WYvSpNB
V0LQuQv3D1Zqz9Mc91kEjW98lBjVBjNG4Atj6RVpZU58Of85RASjxW9oCU1dSeNs
IR+O2wQ9Qdvz8gVwrHyg74xSQn+LcsB0v8KGkxCgOdYItYDSu1XSFMR3DT0/ULao
EJDL0Tzhw4I26nBK/rfU0qRXRXQ6HwKnKsjbuIiJgr9h2lC9+ZxQQ4DTL1aBQ5ll
gVSQ4yctVC03jwdo/vWJ0nYCIpXHUZtgpIWbx+88SSl9nySW3NiXHECzJGrN5gGJ
GzvHgzLs4UvlpWeZzZLq2h73iyzp9uFIHDHOwvs6YscrGm+o0fN3nyCSk2/S0UyK
exhApRGW26a+GRwad212gfoKiroH6Ydnpzz+Ft9uVK0OOqGX+YK3IEurLf5fw8fE
ehnp93RCrjsuPwr9Fd1tXyuQfdaigbwj0eCidZahVfTIce8bTMsNKWiRgkmNYABH
M0jieCvcdpsMtqbMhtLyBWSaqVYzkpU9joMfe4sum1hjusfNCd70ytjoZafIDAbu
Bc4snmDwJV5ZEqUfAtrtzhxR+gtVBqQgYK8WSPKO+yFMMyLZSt3Ftc/ueTLNuBpi
NbooxzYBb0O/Sm7rLn9RPGub9clW+OLAeTjt2TYdC4kpghi1hAwMF+qKPaxsoKV3
af344BHYIOL2tSLHBpS9NUDSCXPnodnydd6Crw3IxN8XUWG5Udt5LBMqJkgXXhg2
v3xkKd7+g4FQQtsJTW83CGHOKvo2/Ulwjlr31rwdzGm/Zf0J2CoKMbr1Atfaix7H
gz2QcnzrzhpvpoZKnDN1oe3M/vKuV5KS90+kGqDEr0IjdvzvLlKaWok42TKnEOn9
aTtJxcKFF/7L/ohFhlDhl7gj6NOSNCJZhFvJcnbjv0ux6914MPpjMRgN2d/2+zD1
WKANychPta9LV/TAfucl/Jdr+yEbgLTl7vy8/0/85OM1fftZV4aV3913dAAOYLzM
6IYHDYafyX70Pwb+3G76oLrSh06Raej/i1IapdBPSZOr7T9Hzt/QgyoTXtr2eipD
j0XKXwu/fKvv43zwkFiWUKZzvLlsTKSE60VZlprv831p3YvGCOcZrJLsLby0dZ3D
Q7i6L4hrP5MHb+R76oQiIQgo1Zafb7nl4chqWncYFa7KV+MGftUrZgjRSbHjy1XW
DxObgnyX2xNEfuNXmCHYOcjzvRiVEKaofWTDxB96aP2lZ7Aab3sL8LQ+bStR1jI6
1YW+6HxXe/I8UCGgHmMPDmKy1r/5npZApLp3cPp7CO6NwLdk6YJEQvfRI+m5aWhQ
m7WEaVSCcicypqKWU03khw5GgKsEhvOQ/n0xPVVIDVJP4v+y7mqAQ6HbevnWlJoZ
58I69Y0fHPj05FBMd8Smw67eaKSzNfPhU2B1THYTWZSTuSKnxrYEH+0XrIY54/XL
H3LE6iUQKbGTW+QAX+I6l0xeoNn0aI+1uHftQHKlizrG5z5ml3wmntRqyDd5pTsB
MGk2WHgXlSSbFtjMqTCy6yeig5++Q39oRPdnRnwYvWp6xDN1gvZ7DGvJvLeOd+42
VyX88xP78vlbAdoqn5QJ/9r6/BwT84z0f67+4hx423pmb3M1AI+kVheast9gyuT7
TStKQOqlRFYEv0K5Kno79FV267Pl+gp1D5Kt3hhtJylLvL1C0v1G78Vfk2iwUiWj
gCdLzhmNxQqpsAfB16VLun30oiuRG44moT8c/CVYbZRpV1We+QDbUjsOWZ+HtgCu
nVp208F7sm/iHwNlMpKpMAaA1ni/+euM3dcZ4L/AWBW5nC3IeuEu+TNWY1y1HpbA
eEc2OaNwj9+1xcdTgPs5U4qt7O6GL3ge2CQuvjlbX8Ibw8pytR0L9Sd7FoAPxxFi
Zp0yNkNXJuAb4BZPLXg1AAXQA6hPXbt3i6SDLJkROj0IyAC6U2rb4a3fO6E3p6K4
ze98dy9uM2K6OrX9lFp6QSuZ9Xbdw/VhoJQK5QgCSpEcCtiAvvmpAOBigk7gWQjN
2S+lEJZy39wUeZpnrAyOiWjNrHADkLhaGq7ppGeG7uvjDfps84n6apiUp8tp+B/y
054RWNqUIPxQ744mgKkJJxW6fcuXMtMDViQlXBYrIyM0Mkt//8QPND9cF9PG+1JN
DlWK9ndzcNpiKT3a4+mP37WZRcCRcIgOyyDnfHYWNYiTYovf/afxvSChZTnTOKIH
cHKlkhijTua0oLGhH6QsKm1dNUrVJ0T/9AmmCNE4M7xfRNB1R7drFAZXgSdl8yTP
3uzWbuoSMYEN0OdxSsXLrTYt+7ulI7hrYGkbX104U0/QbZLIcfglZMP31fpwhTZC
YHnE4duNwOZjKghVPkx4qcDBi4o2PnwJTmiGGmd8LPwbxFZkzc89F8QmrTxkVoo/
DkS02F/DNGv5+jDDv0WSUA3c0C5Do9R1scxrRjSa6YymybNiABO9MDaQQAmxb39i
1L81KHoVb6NdLSwAL1vP+ST56b0wow8qMWcL4aH5zIZfkwR083wsRGMMElcX/HH5
zibfyPS8EN7Sw7Aphps4kdWiZemQ3gTEil5GQV6RToT3IOfwcW6SBsw2PKX34nJQ
f26oUc0vJhtN009kWY9jT3B/nxcT87bTkb84SL39k/P5+YRhujsePjDIz3w4WJ0d
jG9iW/ccAKGsZ3+zCSaYxWyh20dx/pCv+m1VmZ8hzz83o/XqR1Cfp24WEP9inhEQ
nJ8iI4ysW0BPr+xvI661YYnPEQnlysKWBZ1wIl1mlXljMUMVhFqcOjWVE904vaWz
bua/UFjwavLz2IWHe9vjAw2hN3qdxf8Jz3nY8KyYtMV/yTH2F6EOKjKjXzev9Srg
iN62hW/5b600qWaENVXTyfbMKycyjMCEy/ZWGcgzo86lvNWBxy0K2lYKEL2T9oMm
bCQqSI27KL6kQL03EBDmykmUqczNzHwfxYvUdNVtCBgiqH/JzV4E3tYZ6P1sAMoO
FbYC74JAjX9KpPLxTML68n4g8PvFdI6zcB3I7BWjwPcQg0dR7tcBU6IRubmf83H7
UHxMXUcb1bGy/En9BfjiK3EqvaS7on1H2G6qe23ec8e3wc9tyysQUl6rMLq9IaGp
GcmatJNsZN+6ZD9Mhy/iNEsZxsDLtKngCGPn7SpeUAbQgWz8C+jHmXhCShglzbDt
xznjcU3s0yoifHoKTjw2BG2ccJ7ktI1z3imKRtb/ryQL2CmnLtnQbZowppV6ER0C
EPrOD21pkqVAQVccCLWuyAPgWX+ahaIPcz4pYoTfgrwIy1zZAmx4w9H5zcoAVQXL
32LBSTRnKTRdDl8YzR7xgqieb7WoG8zVF3/4zFGn3ir+/OFTn/LLleUoMJp34Ebk
bpjiFRpnWN9cTBDrUuA9ZJJNLlP1etQ/547kJ2IfNT4puyrMCnbuB0Ztf6kLGguP
o6tyMtnkHL+7uLrXkYbZd/lBOjB5UOL7J4paLsngXlPUJtA9kEkyNP5reCey47cE
EJccP4E9vVP6kftzQDtAXb0R4pPbFLVN2cMjHJ78/18=
`pragma protect end_protected
