// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sl+BKKhqHTnF2LUAxcxH4HdSJAr9IhjREAS73ofjwj+3lUzLDvo+yro6kwv4jTLd
4+c26IzQhleNexpHicqW2n/lVx7rbaZGVb05yAUgHIpLmk+5jORlDzAp7Zvp6KEf
dOTAk/8c189GCBiahsiyn+JFG6PHCUBzS+nX16IASJU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18848)
2cDRgz/r+drWulcPJE8+u51nrK7J6KfViQ0LTWCVrmG6xyP4WjW73Xo2aC/rSwOA
DXAiQc6ZJx9HkAY1KBsuv29ozEGLznFqVhrKfX/4THts7pfANmvIktDZbg1bwwzy
YLVlE+JHrqxsZnUVKVuz8ccHj9ghl0Eg/4wWTjK/Y9EF0RjXhcxJhLeoxXNfZrFr
Ce7n1avDi8sMylHa6rKU48BWZvMoCEl35DcsPAV51VL345Fd4QNgERWPq2agPFfF
9WPVRxGXhtng8znU47NABVaP5AR4O69KDeN9tDcfomY+40HDSDXrXPBY8UEKH0wO
nzq0DZMgz22jSJY4BuEUZu8xKI2+oSFuORGRmdWTBCrNm+k+miCMfMAZp7iLm2ey
gHd72sDh12uiolPEmg2k8uj/3DgavB/6iRN9k9fD/yepV+g1LNJ7UARjVDFYqS9I
58qyKXqrjEKRbIASdzwHRdVmnfWaT85cYZkINOUKGfuDi7HpHGmjbcNmPBnYExLz
uthkN3M7gxoqE2HiDLe/wweCBZ4yKU8fwX4q4EtfVXyCSM5D/fQBSHff2VkvVlNA
NrXV/wKOiwSwdJFRbjkcc3ycTn58v+eZzIxV/uJ6wVfXo8FH8Kgw/V50R3fHU3oB
IvUW4zvhPIkeXqAvhQpddLOQOm9JSJFnXKtnBTfyxaAOOx6F/875xhXyovemH541
3VIHEYszIP1tHk1WYMifYaNkm/9J9h+4ap3geH73O4+nByW4weYBbvWeOfvT3Lo1
4r0jhXGpLbRP472n73fBkhbltfHIAq9jvqP1Eq5lfAElOFaEuMJzql+B7ctqRFnN
/WuzfsCbbZHdfr2KsSsh9s+DUkk6JlteuxbKTXQFm31Gvqfsy6tzksLgo91AEWTE
LaLFkSUjmtAKwnklhJ6eHjWyql7ZqET8UKIeo/HqlYbLiOEbU++v/kE6GD98cJ6w
+FAlpWZyGtWjjfE2SIjjPDqTZ2/0app4YUSekaidmubNpcMBAmRi1KNp4Yte1d0V
+o8O7g8ZyHhiwBp1ykw/V9PMDrupa5BoJEmdwHcfuYTlFOytZw4RPNGoXnukS1i9
XMYVAejX6dtWRAG6RiMSKfBdcMwu8DjQptavbtN+5I/kSgsLj6T/PWK9WK1Lh3iw
5m0hEpXqK9dO3oqKQoMKt35PswarVSONugKGKUPpsR7Kj+HtOka+SAUrhw3k80ed
dh/loPy67WYTNo3E+MG6OhmGdmj/1JoFGJrWW/hCwhEMxBhVpQ0jwAefrf6orkA0
owck+QW9V2V1/ONdDFauvpWrGsly/t8JIa6enRufTXG7G+34prtOmnxxRyT23gIk
RiMhXMSqPjmigTTgwakg424SZF56Us7BjTdgUo2JetBlggWkk64i43SnGRYtrKUQ
hJ9jg4OdX4oN/2ILoS3KgQm6S+pPCjNgMEk+WvnBB4OSZJ46gxQsEBpVmHzYg/et
Ba73Fv38PoVMLq3kFG223jJuWxPlA14zZmv5NAwJ8K2QcQbScX9Bn8iBlg9elK+T
O8ue9YxEp/2NgPEMVlqeSSgvjuGKM6yZb4X8TW7zzS1SSo+kriwXP5to41nI/OUA
oSLoTM1SBaRotsW6faRtXIFIHkjCIADYs7S06Oukzt0T6XFfwR7oKCuarkbi3tJe
371H6u5x6oY/XMESBWsvlAcd+zmGysVjZ8iHb7gtXeg+4803M4Rol/vNkzMdUP1L
2KW5hVlkF1ILjIhV1VKerirx9YnFseHTfNcYJsvdGimFnF/9zxAFFk7qqj2A36Ac
n87LkapkoGefcx0wmX7CIx2qkTJ7jE02+my1GTB6Nf4QQnpauZXUuTkvyCZsz7gC
EFbTwQwD9hsGzVS5PamGLgVTY3ewz2wTFPi6O4ugNgAyl0SCqLKG05zVtvudAqrh
R7SxHRxklEFtohXnX6c+0USn3by9FNJA8MVY97lZDufm4Y3F71486SzXmODu9cRp
rUpXMgMWhL/c1uQULClrYXRKlgZDZErQHgqQsTz/CJa27bpAbKOEfFQbpSd7L2OL
uod6Z3K/z5gXTgD0qNgKlGq2Lu2QkU22kjl8B212c1AnMBwopVOS6usMC2Mv2z4c
lwNScP8tfMeSGBYXJEZZTrTn+m7H0WTYhARcnGfszg95WLTFacErZW9YQKtjkPm+
HD/zyfvqP2p0AcNK80cPxJJ4oEUW+RCh0R++gGz7oLlZFZL8v/AvTlXXBag5zHJV
26ZQIrARJG2JH1AYxowR4Y62zqSitoM9hbMGWZkeYPJ+rxMMTiuQ8R7pDAgACFPe
TQSQEL6ScITTMui5HBf7CdDSbG7AHX+3gHv/tGAr5aejWuc7ZwAp+1iSIA7sdtz9
8cdh3dQ0nOC6mNzlkOF6kmK5Y8xOOiM0ObQeVwrMCF/vroNs52MMKjPF/vSmeOGj
0Zx3IolL6KNYMG3HMqrjf+ofRoAXv6dmdNDByqzbvbVg+2TNdzfBwfQ1EHBbnQPN
eEfKJOwXhXMgL26VVOkyLhRV/V20Scxk6KCu/9G7oXXnXlEgptjnM1a8Yr6ns9nF
vnlzrV4dmXEH0GSAV0blBk6uqLYIIiGfp0lAAQYAGGRU6yiO5t6RQB/4lyVovt/f
bydGmJHUUWVSYgWVhxy2G2Wrsgu6MWhauP29C7yvquHSlnEpTFcMOnGx3qdlsoEJ
aSY+Ttw/kNN+8IyQicjQ6T1k/k6RTr4TMjvNcSxFwE4fUm8t5u0+vW5V49ASWbTf
Le+yQ5uBqWBjoFFmdzCsYwJdh26P4Q5saKDhxEHq1q/Aezwv33+5owjzyy2oELB4
qWXjP1DcBJbn+Ilu1ESdGFkJDrmEFK8qlowtI0uDjPy8qvqoXBgoz9zYZxPkdEtf
SKTGN86APRj0dVqNqG8i8Qrm0vb0ufyEh4P+t21bbk7BWvKb053Dbm35ZrfBbC8x
VhzkC47De6gZujwbPDDb7LZLPfsSDLAc2sTnQHVLyW79EIz8AWJVWj48y0JR3F/Q
MLp1svkj7U6hSRDzvCwcxeWk4nGP9XqI+imacPHfDObpFzSalR/s4ZWjkb8Z7xKi
ZPz1ZnTKL0x5/bo+dwD+zXiKQu/mykJTTC8rmmNvZpl3qq1Sx8M5g6rX1rh9X7cZ
LLpAG+maP55YAmfdtmJ7guTVLFVIkYV3wz07C/B6K64uMA+rGZOnLTHcW6hN9W+F
hnEXiKzJBYGHVEDaZgcgxKjfJY66qEgGEE4SpmUIxL6ZRflWuuFN242aLFigqUH9
MHj+bhmaUCoIZtP52DX1g20FKEhnTpTVBG7MuJLyZp0SKALmv0DUmDv39qTj5Y66
IktME8PzQ9eCACnFexKytfYx6LUKVlwkb4/0F21tMNlkk1EDJP074Gs+NbtIwMaN
VwMkAkN4TRVc8V7Q9L7CdM3rMg/FcysYogwXQUsIvOfuJu9Hzm7sdtrOr2OqRQPz
DF5iO1w+bIOiWgGZauyLPv+A//3URBU84rjTHhLCJeSJn4L+4Zu9XcHJagIFFHUR
Unl2lBAV/4ILTphK6ZgYgCpKy5X1Dyoq6E9I4DfXD4Lgmnbxc6gmT1joRPtq1BV9
Pp1J65J8yNbSFP53RCdz9VLOuvOFSmxgXtGRX4P++bMmrgSRGJVp7cHafqqFtRhI
uQImxFOZKZ4QOxW96C/nm92OywteKOHEX84y7nFFZdJCVk+AnBlgaL8wEi1IdA88
rZTM8tlzoxVnpM3oOKcbHZr76lJLDF9Bd/IX2YzbISNrBqJxGFzysGEQHwn+eolf
6l3xyn1x51U+DI2LYPFYqaxvDVNjiwraLByzHPNM/sHuPu6iXn0+jmy51mZJCHmx
C90UJp7MNPHhXSQuTTkWG4MG0vBNdO5BsrLu1Ju3L/2sADOD942NL48IFkHplMFH
4ZWdbuU7NeGauSbAsmx3OxFpUDud0Ci+iSvSGFjS+oce3YuGRfI5b9V6tcShvL5P
J2G9VU+KMp3IDfL5P9QGaLdaKBXfLfI16Kl2rsWSN+R60/8PlC+HpJ41iw+gVPWF
hvGzLdThABiwLTGbo42hjDyAWsGQ6HY3Zdoo+CHbr1Am/msZ0RP+QTXx61VwdxKU
fsEOPMLIlVbl1iL/hPJGoVi1vHJBpLyq0/gaf+ZGnYAcVOSUBt/vdvdIgXJ90oI3
raNBTY3NnRKPG8H729xy7RO3HLXRIDVUfW7FBXvajAF+mrYOH6UFXMxltIH7HnGC
H9lfm8cc3BahThE8OghNLA1Oro5insx4d/CgUbP7ZzhFw1RBoUMzdXHBVtnyyLH0
5SorJuD0dqMnkkZmL+p+CaBh2tUpWvVRI7NQv8P+VHyV1SaVkQs93Y0pPoexnnaE
XJQ2pKq4DzkUFFevrswLuExqJXpuiOllgMlnjsYnlYZTHTkunJvYV/XVuqUVidHa
eSBFA+Dc5EFAOdLooy/0BuN4M9X8Q4O1Jfvzu5Vbz9AjIvdlVeWRK2h6BxAFGD/9
8wINBo57yGTCodrpCB39m6DGs5WEXGT3+8sZb34FIpWDYVB2lEv2qmzZGzcammxG
SVP6TWe0N83giFy6Wght88eHwTaTc7ERJYWs4UOE2UCUuSvTUmSs9Q7kO0wbcQy2
rkXLHq3f5XXWbCLLnrx8PmR/70oAoHGu/lq3sMBBbUu8r6DizOgBCxNi5u/Tl7Y8
D0FCuIoHyrrbNBvSE1RqqwxEWU+5wxdGEAc86ZmGCRbKFr/lwCc2lyrI8ibsU8ah
wvZMsV4f2yoChOycWmB/ihxx/dhylR7SPtZhHoacEkMtS1SVZlXFMb4DD5pRK7rq
TqBeU41RrPmFV5+fJlqo78RAsGTEv2sKt2dmcdnvpn3OhcJkYwuMqNbM6uuzDu71
56MdJy/yUYbgeNVNu2qwfNkLA/ZJAAsqDlys4yX8LRGU2R4Wrg5yRluXreATxgJH
LkVQ5lH8BtbYykJb9fXAhMSqtNMxNe7ayxv1VTkiwXjPDTjj4YERsmUiktfjwsx5
e2nxN/DhYWklAmgF/IkCtWiLz6NgJp3xzT4B7ZdHnN9ulbWx71iToDKCMzrjm09a
WioFNptZuMlI6ZESA5B5eZpb+b/+ZaCS4h+BMLfLDpLrdQflte8kVIAWItA6ksU6
Ytws63R/Q/xXJv782RA/Bash+3/0wYb5uh8NR04JYTIpKC+m+TdxjeDwZBhfZbUQ
QIjJRaEt4D41fTvmdV5VnztPFUcLeUIx4LSQrxvSoa59E79mWrQV2UzfQ6hAzyIZ
f/skyzN5l2mi0jyne9cRHfKLTKKQA8PQsEpxdT6m1lStyhP8kyzAhaJjXM/EF21D
fqbukM+xj6xrTzyROPVshZVXsU6mZXDaGJvNOCWcQFjJpMshxxaAIaOWdEzCVuLb
CFocLUFMT84RtG2K+8G+QSk1Urc9IwCVfKDhpdzCh6u67YHz8YdH10fuAapb5U98
H6DrIF0qEWLCVA7koTDI6GGymX9MCLIZZeWZHdi5z6KCO5i6hFUyv6NnTTkIeOS2
w1nZdkUypEqQ1XfCXHMZhTFWcwAwSsmjvdnEYoRDTorRSpi9IAVRNqnWc5sUfeJ8
emjLpgcSiCo7BZIYHS/ET4qMQSvkbXRY4fwf+ulnvI7sVvee9DepCtcG3lnPcp6k
0pUTnZ/DN8wQUoeuljegZTCFqN53B1SdqthWtagH1Nh2kOnCXeJsUBQRNzg6S50h
Ma2X4nlh8G1ii/YTqQwKbEzWB3fw4IGy9EP0yP+1cyez0OKPd7WlS9WQ++QX7dX5
Y56o9buWbLyubaQlCie84oitcp9b6L42I1S9i6bjwvCnDDV3Q4vDYLTm0KAIIUjE
Jqn3ho7Y1fy+j0+ejWwW+YqXLPo/X2VZeUMEb36UR0gDvZYuFv9CT9j0zPvLFSFz
0Q3R2t0AMJg9E1WugMnWoK7G7K1ZAuqSEMduOTUom6RJIRmYSNNA5hnPHbV0d89/
sinCP3aSEZuNI0yPv2FRAmn48jFzHIgfHBJXmwga2S9Rp1ghJ2tPopNe2s0E6wDr
wz9SvMxjUC4sHt6orHE7bRECNWSg4NF03vJr7OFpnA5fpsRoIVc209dYNhwuDMDR
SBP/2jfbsbOm3hJ93NRbf7LW+wRBT8j0Jm8R0b8wFUYUS1zbF0YZISbErymXadAD
v5Y+r09aKbQFEVR4LkYCZVZYP2Lsd21y/uvdQG06zbuiht0hKwTcLOp3BSphmcvF
bI0664FjjAiG+lFWpkaX1N73fFez5ZPFNgyp6Ev72tjYU9qd0Vxtaqhax+VUnNgj
NGvVqSWsXr51rjLaRLzHObvDH9j1VVxOd6pmU+0ZkpiAjgO8UHWBa7/vbJw73yin
9eRAPzvrbfpxETQTuqh06KyPTRgFzuDUq5cpBeNx+jPOAH9Qfew822vcINx+4wIx
odQWV/B8JUOGMeuZnzpAYRmrCTt3Y8DWr6hA3cBM9AmUyLqMjDiK3eSbUZ6rKRLv
+93VQRKK3+BAs1tXONHupAX6fY0+xSplugCaixc4zsT9RsFlaQ2adwr3zgBJzJ8b
21Ajae3+sqJqZPHX/Pl5JBRvr6ELZp1FV3i/MA21fKqBIYahuLF5TGqqLJLDopdV
SLra2k/ePtj+w7mwSg4n3NY3eopJW4MJ75zKPxyrE5gbu5FdaPRYJDTsuZFPP7rM
A6fZO6kNfh7VI+QSm7DlThvOa6xVBQcORrtIbznWZaORVNKl32l6zsZVwNXaVMOF
MKcJJsld+1s8dtpfqQG4cOKmVlJPDOx4+Namj4oAT+NA+LLtImAgzoNMQIdOPT7t
BZrIeGa+/ZdoJPEjbYxVRZ0E+qHp2TgQnvwrfvd+6VvrZpFeWHdVHAvGlrJZ65Io
0PHtt9CvBRGBIbAXg85JpElnqPSUDwJR2b8XRde/BG+V6Rd6D9xzeI7rjJvCV7Pi
CD9WtWcT0wBxdR0R7IEpu0/EOd80CmI1KxSpYxU40qyuSpvomBh1BgbvRe4bYH46
rLzxDv7p5pGuoyOe+Dt/HyYFbxO7N+h+ImCvMeM+rVS+eZuHj9CdURizZU4Aa6MP
waOnlvhA8MqbonNEGMq410jOqYykuZMv4IU7PG3CSOOQ59ef6xamWKlTsg3SH37c
pJIQb2ml2cmWD7glFtHNr35R/Gn3iIRELx6IKu2Y3P4pkwYesDsIG+3DNdmRQqzm
qyZNvHz+usiM9BFGVLvmIJ16/ouqiIxfb9tkg59nvk24w/7KU1NgAdLTo/Wo0tJh
31rAalCdl+7P3jRSp3sm5PfbOCIpk5NBsSrua5YV1CQS+8xk4UT6KgmLZjj0oeFU
vPF6Kmqjf4VI0N39rR7UMWdVZul/Et0atDBxwhbIfyr179T6hCUzjVnbseYo0VrV
9z5ZN4c2ZjwnGbSB1g3wTErRATS2l1PCIKgA+CNEexHBI2lFgHMWNXWP1XWeyDAW
H8sAYPHereXwMefGuTH5W0WOgjQhi+DW8gDein9RQYefIE6uqxX5XU6fjIpVVu6J
mzvh5LaEtyCxMmEcBg0LHc8L3YssvavCWZZdvxtcgs8bpMPiv5zE2qWCO6F6I8F0
KBhjepVw9P33D1Ni6GyyQJw4WLCKWfcTXyaMPzeij9IekrQXnJHnU6BBZ8+7H5gs
cWsQHhBqU6ihXctg0++m5lRNHKWM7Qm39b2iFpanR/Ce0z+cb020mXIAx90kJm0W
au+TiJLmi+H6j0L3JkeCF0A+K4wkeAmagrcOWNEy9TcGEixckW8w2f+5PDmCMipL
VLMQ51ffNSKcGImKJwfCz4BeQ9S4lHS1/WuoDoSAjlwqyVAj9BYhyNQfEVgrsDXT
Rd8iZPLpCF39xJQkMDtsBMEZfOMaDFkdXC8ixIE1jDxJsn79fM8aDXZfsw50P7Ld
JKNfhj2A4IUhUj9fLJGi1oq81PSeV+O353ntWWbnvCMZVttoNF51XLrd2+h3NyUF
Cla20YvhBpzMLhSzp2lath7VN+hUOVzjiGJpFySW5KuBQGl09aSkEZaCCSXAiFU/
M0EoCRJeMxxhX8Z2H7nr7+2zAMLMw2696FUcq3DXkUj+zqYNXlulTmdUicE/Wc1W
PUTFpvl0jT7w9ZNyZgr8/rEzqtIHL97NEOlMxc5rVRBwzmROIYa9ULg+ac+yRhyn
Su3DV2uXZTNggFn6Rlspt7xMyB5IgZwbnFP8qdtd5Qad2K0XGCLrDqsyJoWuvQGp
RjPSM7ykX0PP3guZnmamCM2P0BoYb8+Zbm1emY/CnLncx8rSSFAVhslav+ez9xxZ
2BlEg+GRyMG00oOOodTqn7AvPXRnNOCtUi0InIe2NA3qX5XGo7F9g3nZmmb37ZxJ
CY4qgiMEaf6LMM68aWbVuNVYkLbDnXoAIGNK195mCG0UESQhb4kcVnJMtite4raP
vy4b0yYMXOPkFmzaa6kGb86BGSvQbP5umHDujQx4LSj6nv6vGp4tsRAKH2K+PC7z
Qrc/1bLgZUmtfiKWMfBCSv6p4G5kXoqgONw8uVILM6X954CYTZrLzMjHwvzvGFgi
QlE00eRU72lhBjld/gchdFQTzxJEB1NnR7cNzLCouWYFVLzqcFUn4aBi7UfrK998
j2X0ad5KVHv8saDCNNFd9uibhdJOQrEgWlsleS1carYgi9/ZqyGC2AwZJUpEKePB
tIJCoFe1hC9iFFYNUOyRKqxQeQfd31X4NMwwQrRT1mebT834CQUsezqylpM7ZWXK
p88XrEmSVrqo0AGfxlBPjhfpCnQ87pF2cCIDeh47r3dRUWFAoy2zGqxAzYnv0sEF
W7m7Z34+GVP7CEiVrEpQOBjV43CIN+8dX4uo0BRgEhTNCYrvIrhqUSy+qkoza3dQ
Wa/2lfmWWqkRoRiGOnshUaFTm2YydOQy6wYMINi4HGgR6ABqT92Tmdt4mBfipD8q
V8XzL62zm2LIlXJ+U1HeZVO3IAk1z7cnlz/vyIrr8p60RmEiamO/0wBC7F/Dg4pw
9o2cUMCG7XR2KOYBeooqCuLPab+4ny0wc+aAeS+/EMIoTssFjXFquQoTiiUuEZ5H
Zl+I/ltxoQM2X+cvLmlf6gWe3xPZVjwDrIX/imQRrE1aQnunKNgMxBeXLdc1Izcv
STuvbeocmlQ6j/OmUt6T88u+7UZscQ4fsR2ko7eqCCwTpWwRpuAFt+2LoEfkz58q
hoEmcNsvAl88D9LrTRHphXBZODc8K2nq4uJUEQmIxytZHUQ6k1HS2R69x5mUmmbJ
stgKgC7VcPGcsmz5He7lMLG65B+owHNGdSNSnKGwfQBPnSMJ/RkefKl8shtnhPdh
rVdGb0SchQAYMr7nz7vg8qnPtQvtmoryWfDh9tb5P810KL//xZdq23mGGxGHcrYE
CjPgvQg2kJUhObtMlDSM9Joezt6wJ6r3Xtu1Pjjg/nnkJfU3WtaTtGjAK5ke3Mz5
NGUl744A5vHysSrcDVvd9k/1avRe4CawMThMUK/K5Xk2EOBMXLv4EmEbtpMW4YBE
qpSMo5Lyk/tG70aDYSVulFiI8j6EQGTbZJdf7laAHYoC3idmNwUd5UXHDZOlSdHN
yqny04rsvW23k0Z+YUt9V/YbwAvPngItioENmVrHZqbN7+1IVM9r8GMBx0iuHgEz
QyUFO+iXKUyZjxebOpPayJE/8BVF9tIUPQJHQ4cCBdL6SiTaEUS5pMMJrVI9g7Zv
lCfUOZAji3bMrSzungeQca+cwExuXWHlKtna6mL1wWzVRtrG4ksxKRlEfrVUVLsN
RSM35w+Q8+JPDuvxyKBEN8iEp+qVoFZdYTrTRjrLZu2dc+XbZiogpDahRkkK5YFp
MgcejvmVyArqOwxserDCxrKLp+pF/Tg11DqSEflBHNo1qeUvwz5w4Ndliijn2wSi
WCifGYKrxVXGuhXSKAzpy+MrZBxdOY9mXL0kB1x/teBYDBDd0myIgTfvV2i6wtuC
hib9vwflpljC7qqmZ93oDp+KmQSueWRImO6BbidVf8JarRe1QhvgmIfFRQ+1M8CW
ReEAJvkP3RemVsM9b+u6RIS1xJ5IhaT3VI1hpZAXHKtx6rHc2kC9d/khuaAlcw+K
EOahsMg2m33aHTqfznTNOCiws4YoK+mwSMJI4JClfYInKaKQCYIePG/2pzpgpSBo
5xeXF2oNxe4TKIWHZGGvGImZ94aupsmNhdQNyQu4I8EHkp0hSfyXC99QtradmiBI
xblFAf2ofq2Jz5erGinKamxvGSFM9ponqYHfmQSr9k4IjqRV1lnqkm9YvyYrHEEQ
zO5x/oEIlIcm6JhIM8XOTiL8Z3SS7KRQMbpv8w8G6C2UzZSdKWis8KDQCDhvY6I4
YZeF443xvR6WSgYqri9s2oSFpfAhPlm7514HmcEDAZ4rmr+/dUFIl5LE6GfxZF4H
yaE7501POuUPK4vBMWMwXwBvOhIcqOSTWqRYttoPENyfDsofOCQhdVVdifrNV/W5
sy+nNDPdbzxXqICuRVCw98zdt4Kf2nHaJR+BAduA7VQzrCRAAB18MC+6N9LBPNRi
hyLhT+2/kGj377IYgvHYod8FLRzNvC5plYsqtaEXjM96QE1RhSttbOWGaGOTD1YA
fSiqsRTmrxkVo5HfnWrluFQsaeGxiv9ClRtmCASjsoVd6mcEw5kihhrePkZHweX/
sedq3dXgnZbUnPIl3p+qQGOzDa3x+nSy6BhvIRxYsLbx+GXJfA1Tb3jyMuwF5XC+
/kiUpGf/+ecaVJEaHDy80wsSgkrBYG4eiC40zUrXRhXZDwOuLNhRvzri4eEeaFwe
+Itel9CVU5sL8DYJ16kq42wfV4H0V2mMqjdNpoSF2IZjFQ1+RoZ269rZ9rgOXMNp
qq8BPEbbGHPMp7NLIxfFBQMaARC/BYXnj93Lroj2A9+1rboaf4W5oYCyCevaeJ0k
13ynbwmRWAvl4rpcIOj7MTAHGZvluAZidfzJjBN7imo0UkoJGHXRCsetVmnptmcY
P6wQkzcr14MA16RzHAkJMi36Gb3BOFHchM86gtHjbOZgYwbOb82AcIAxxH3LBo3e
MnjWwvNm/sz02PwgCectENSG/UJ+c8Qjp/t6lHWSsUGrz+ZQj1F6c63BAiKDh6+7
ZwJ9Nw7jdze9s7+vLGZ3YVxCYilW80s8LK5/d8RPRVkksBToi2WZwXE09kwnAEbF
1ccxxQL1ECO4D6vFecPd1tBoEGJKkK5u2CCat/Dt56adWQRYtIh3jdB446Gld/p3
iM72q7c4e/AX4Xt3mL05x/ZaDtmE0uovt+Vdl19oi0P7dCuaMP6Y13KUHTlebGrq
SKYegetKj3Z1cN6kduxSYtLaoQZ7YiHkdd6AwyPgx7DirjzFfi6Uo2p0H4ORlKUy
qCwI+SmxNK9Z9BoP5GaGTk9tz9iZynu1oq+l9V+XsjtoF0vKaeLSjEffemkcvVk8
Mhve1Kv03PLF4EiatFYv/lBl0JHtkk1kPI4UF1s18RmXYkPAZrazi43rBPhKFceL
04JwMd6CLrW3NfruF2t+mN6hrTtcgs5GChuHLF7lc0PuodrM/uKaW8ib6a/mq6Mr
u6W4nRiP/eh68pa0D7hwSYybQvo6mbrFW/1eknH/jEscjrpdbi6jk0Tz7Drq9cD2
hZbtt9hdzEZ28BZf2w+YqutU+5Kqe/FZFwPYDk8zh/rg5wVGQYQqVTA7N/U6K4LQ
zBQlURA6zBwAzvorLP4Iz9+hor+CwoU8a612lfQ62EARdZk++7YPZDiH5xLpYi/i
KitV+yQahKOrff/jmkDF7PylhFD3H3Ja0kOa88pOckXpzEgYS+ZVM0LEAucIRMa4
WvbdQt1LFV4ZyrhU0rfrRkmvW3Yj/RHgCc8/+ocz+S7Sj6ihOQNojn8+IblQCenv
5w89AiEniM6X4eOyAN3/gc0XN42O5YAzlnbCfVGYgCDQFSoL7K5fZU0MDppY8gNb
rUddIcWB76n8gqp2U5h6fFcI0xTfz7I4E4+u0/ilZXQDgeEau9yY4o5rLZdhTtvJ
0N4ZHYfeETSJAhfhNsfd8hP+cRlbgLNd4fq4eBuatJ94Nyldna6YQ47qBfv6LZB3
FUAzeyy5gfZnYiCEz4fDCAmlaFh8Z9VkGpG8DNN1vVedsf5mFg/riymXzjhn6IUB
29m2nh4AkWZwk0M0L5mOU6GWCBXBIhA0rlt1fQPsFIiTJiSH0AbAToJ17O36jhIE
jIfJN5xoUmlLz9kanszHhn0s9qLAbcMbwPd7YQdZVVl1bLTgn53Fi+UW47w0mQAo
pZws6zPvXCpyb8uQ24PFZSagE+Qc03jiXTfu48AR4iV6EnEs6SxgIKYvCZzIQcya
HDkfUs+17KWchM3tAgCQB7Ji0Grvt7WL1QyMmqMzu77qVuPwj10HITggXkn6PTBn
x3+XL5/3pnNoOb2tDRcumR7/7MSE5U4pDO6qCrfE3WU+vPJq65CsBHMlCnWfy2TI
CE05p42HUdTuQg2sl9YvqXbKt7xJR5t5GqfOqVAdP5eLzl083lvuphGPIGw7mEAC
tSxDw9IGQzzrvgNXX+RaCpteXPbnhQd2/KybDCKLQL2Mhb7t9fF+cFASKHZP2QyO
vvgHGpr2oz0o5dTfBUqJu+pxLr79h8WmdkCL5Sn1Sos7B9Fit+iOFkqKoslpnlm3
6OBZexeTe4kHNTv+NQHn0CmcDZeSaYdWuNBbinyeApzKPk18R+YluPuNsbGnhUGK
qWLEPEikzdU+5OFAivh6Rnpw2VbZlsF5KIDS0XC/UnpIwu1iHpGyWnnEEkFHqUuL
stu+Npb4jzMqpr+aA3brLQrJAgQy1+V55Ti35f/YjAhPGR8sY6RQfAZBqq2zuort
3hVa+roRVYBhroos1aSBnbTvzm6YajAj57kBnXTrk+p/bo2xDKJuQtGGsTTwRR9+
JC9i09zbjtycu5zP47Oyx+zMMQbYIXtZZNVE/S9PUWGUjinYid0bOSd6+ZbaIt6s
p0oImAOlcy/CbWbTcRlAJirkputh6YAffv+JGWYsBTKrY6OPGToGDZPtRdVUBFvF
iqJxZLxA0Fbc10S32RFaEtSjQR9OPKC5aIOqDG5wZGr7yk+uMYxNg2LcDg+Xk84Q
+klzRGeZQul7jVrobHwQaTdT3FoecSuZfwzqloo/2JnT3M8zlNT5a7ngZ2Z8DQpX
khwvwFr75i5nDv17TU3OOI8HwfCX+jRPqc2ZzpLMFPN1Q3WgHu9Hnk32oxR5MuJD
W7CL8IcbG/t+oeIUGWIYT7d0fmwkXr69uzAh/82Z36I9wfnLkD6RBP8sgVeN6DLr
Xl5+n3wPCDd1AKqVo2I0C2X0ZqKd+6NBBv95WXSdLjvEyorUXUkyb0hRobjWKaZW
mIXSgda847bTsYwlxe6wpMb/KIIlrc18zL3WaUqiKwSyURWrdPm8cJsB2qXv1S9q
GPDrw0ngxaH0DXf4LDO51gmNTYsklN/SgtRCWB9wftY3dR1yegPH9zzbL/uvm+9n
U2jnKdt5J7Tih0g3jAUkWVHZJ9JT9chVnKzcjvejCmXWdkRm4J8HhU91Ms3pFJbq
aQIBnOwHaWXrYw5AUTsE2OeIEc00f9teq+qr2u3lX8cQ4D561UAjxVzfaHYugPds
aDVwvKo65qZ+DjmpbTkAqhQycLPr60A3Y58waf6k67ZTKrhV9RtEbl3oWsUGDAdm
fe59uKSEUaT8OgEzlJY9BGHAQBQEp/bKg/vyilLD9kFDlG8gsbFZZJ+aO+9Kn8BR
7XW35MYXYTH7RwBdGopwx28vEOdPOtC5aD/wjkPlAh0T5RZcNxBFt63HwDrKcnZy
FkRvQMIznIQEF/6HEPNv54M6IfoKbXfvhYZ97lh1kqlP9hEZPt1Y7HBmdDKtZgxI
/0DFTFgaJU9sdfT8WSO13sDX7IN9ZAQhj1KgZyujZJpcUJP35tZp4bVG1E8uw/lm
O2WH3h51gfpDvA2UFveF3TPZw10/ab4vXNn/LjKqXDKMTvxNhRGJsqWS7ARBIAlO
XZzLIdvKhMXYnIX5hJ+UAst7cD6QzoaSpfDcAZJrfluIzYTVJgHhx064WtbYf50O
s3RuPpXabG5C92bj9vTpbUhHxnRUWSztPhazidiQ8Y5gRYeor04v7kNfzGAy4Q6d
LRqf0VsQd8oOeeb2oea3pE9LFLLoH39BUoS/Vs6YkUxLLTzja/qncKQwLyJbsA4x
4hUFhAZNmcDaqzbP7+2KwDgThfCO4Uz9v4dF7MQRvVzhmeybLv7nctmBbc3ywl2N
sVoMPQL7xV1oStS7P7V2yScZfoNyV++5znV6uZgOrvyakeSKSHSfhnSIsTDiSqPr
h+Sx0pJqTnOt2RTsfXzK9/QZ9D7+F5+bPB3CTIy66TXiL4AY7aAbRcqGc2N1DI5F
vWqvmITlVLINBzQvRNOTlMXbvl++10LjSlyDWT3N7Y2+lqb9zz9sEqxn8d5cnlsQ
T+jDVy4aGo7fLH68OBFOkTfQBRvB7hcYjNwRClSyOzT1QaXyBizZeAgYsIRpqFKX
1EclLICxtxcdevX3Ooi5QfuDt2SmmJk4Cc+lig9mj6izJTmWl/q9iKBJLSooCTDi
/GSDGamO0wQHwD3ZifxGQuLktYhus0hgtRMlM9/Tj65j9Yyt/Nr5vpCPsbMBrSMa
nIBY0mC+DDL7M8DtoObN7/RzVbTAxL10rXPCRY+nmgxDSNJ9t8fMQoOy1R0pxae7
3HujBMIek1+VWri8mwuM9vAhgUGJ9XQLY2cd3GIiWZRT+8eprmNPGy5L/JHiZ1ZR
GA57QAJq7wBiwKz0JdFubZM0iG5J0Cu9B4A1rLUAh5eul2HVhTjsL8kMgo7BMbk5
j8+MUjk0m2C5o/OXMVaCSYKwp1jqzZ61xtCvYyPdY1z0RPrCCN3VbCcplnHR9am3
jeCTubjv6oopac8wskgIt8uutSdOjFzBLnaPc4xK6A2kaAaMX+MFejRxmgvC0e35
QuZX9NRtM46z7LNEzKQMfEXO5yS66VnbYF/5NZiOosqv8dFCuyTEj3ftYs+dJmSN
5G24qAt5lG0xBljBJb9qX33J/1pmCpS6tnLleSgy9su9xqSBqtoy8USr5QoX6WTt
JzVGq/l68EqvL/BVHzV9Flu+LaxrSgjFUKbOvGxqzhkUI/+TQZk7xHT/edcp10Jj
OUrbsHhHfEmDqKqMnpZYYj9xv3YprDFuVz6GBgRW3RZ0Ec1co8ayPN6rQPnaQ3Xy
QaHADFvWGV1m7SMTWE9umAkRA4jSdpL+5ww9s/i4LDr62wQ5+g/rxD3vSvp+wDjB
7gjQrZ5kpNOdxUiNVutZhi3L0E2zKgVnLHoElzhnzPK41/K1KrPYnzKlWzDfOHhy
H4uEyrUytUWt5gMuqhDwERHXbAOwn0AdWdsRiZpGdAKwd7N/k8lrrxqCWS5JFSC+
R/OqbNfBythO0M7rn6ZgnuV2im96ItnKaJ/zW1Oz22DJlA0MdS40jRVKNupPNK89
Jdliy6JIr60FwMeb6lAiz78ttv7AohppKdsfPVLWmKcmME7ZaamKtFm+s9WPebR0
P7rU2OYSqmHtciKw9lOFz7RYL/6XL0dU8Yrzxsc2zNbwllZPnZkswOQ8+cStiUMZ
TcokvJTjQy/MJcjNV1x6D/DXNPpcXB2YbHnKhSew0DA6H1LDBQXbQrocV/W1gt+1
VRKzEgKEX5PhG9kioga3d4ELBnkkOnhKoduCyyHzyNdFKCn17OdOz4dOVl96+GWH
FGMYoi30w8PH2yEsxlgvs2nfrjnPvKdt5wvEKDHe1+ouz7QttYLzoUlorFIsFp62
o00w183pvSJgAFIf92cjn2yLyfy+AJgXsQIM6kooIQqKgbCN5xNCe9zKzoAe1A3O
VWQ2cHEtKN/VtXVn+glJqZSGfAgyB1P2yic5rpB2fKsf0oYKO+J7o/HY0silH4XO
QctAUGFhm3ujhc7CFgsT+lJbkEAniM/UXScJ+r/AaWzKEpGdSxe/Cx+zXmdsGa2z
0hhCOn1qbWfVI/yvkN6pAaiWbMTQuizYb3sCuyCe/f/256YbGr/V8hg+rMLg/HL9
8YQYcRfM7yyBkC3B3+OLJ0CzGMYHQX0jaHHHij3IFW3IainhnPbrrk5PcpAZm8SP
WExl+dfv5lmdV/yK1caO2Snj6N4KF8mjxFPnQ5la9NJBK77keIzERVrQcAWayUu6
iD3lbs45dZeIbgl43m/ZdFmDsdC2NYNFoCc1E2fquofxSZ862RjGKLprjCGk/9O4
b916dsxSDxoZYfuYKAn+JACIf5JlN71Y9lPH37jRTDKvGWvpARxp/Kv4F0uaVVFK
5Na1RkbleFgKv2AQgQp59PE6/HU4U27E+KQ9kF2oJL1xZhuoBva/ZCZUVjnYX0av
wGnsKitvatfCJm63PUlbE8nb/SGtb0DHy5DdAgtYCgn6YcWo8o+M8IzLY8H4waqz
vG/cbCkgEPibd3LA6vBGT3xSfHZSB+QIcNDyAXh0TjlGYLQWHQ3t8TLsLRfS4xLe
pjsHTlgTA+jd1Q8tLr7C9Ek0hORlACzSvHeTX/ddXb4ZJAyw+CEgrax+B3s3nLyY
w/jVpF5ePbHpZNph/XBC6QJhXwFSKSdv2tH9pb3UzU19PT2BoLQnqXwvJ/bGr4cv
Lf6s8q3dbib+hNrJreWBIDC4WJ0wYoYG1JB2hjghr22m7pmw7q74ieTPyrfJ5ovu
hqsDzGJmV+Xzwlp99AIMubIxgZS+UKc8eeRmo3mkc/mF34b87r3rmR/pjKRMLtie
KWTEh9FQBNTQIQU5oOebBSPXMXYxlSvMWg+wUZBVD3405yrD9zD3jM2W/k8Em/Ls
MZzxjwyjaa8W+2W2j/t0oe1RBweTLGsb5K0Vv5OZlQtsn+FOd9sG/p3BpdcsIivV
kwncDOj0fqIXMcynoy8nPfOzqi207rId9+o7Mu5SFWeAhZcP2Z9qflQhyVxFA4U7
pzYO1cSFHZ6TRFqef2roiPFzBc6ZaoFjgGvqQ7f8OrhDVWeJUiytJPojzwP73NS3
zCgtxCJuJXqA93/B6aPEYWD9rbUTa2hsy3xMXzQEZMZBZ6JLpdRNbr5edyvC4mGS
8S3zBmMioQH35F4UXGs0DawtEVjlaLqA5khPcnk25n0KFEpWmHqnS/FZFPXo+m/y
guOalM2g4VJ3//9+6H0HZZpEYjnBeYdcubs1NNGWIMD3sarfX8Snqev4+rCmE2MB
rUfH+FWqrrt9cANfVB9X+vjhesEBWTdO+xogFxTwsV34454sfemR/1OApj4QbZpP
6Y2URU2hazKDBE+INNpKAuyHmDO/Flem6qkuInIKgy4fhWCasxz09ErrNPhn69kJ
6EFd8OeSmZeQ1feC1hRLdmAe16FnBTsT9DlyR+Pts84g0d8txYwhRaGulbfrxVOV
htuR8EJwLJppIWwUOSGT5F42NNwE5J00hVl7Yg4H9S3XO1t+mRUZRCf/ESB/xziU
84TkHQqNpVm8ylBKskh1ndm7VN1RS8Qyp4rO7xcnQaCK4N4trZazySa5Qbgs74o8
SipabmQ6FUXqKtwHTRd7wjBOvnOSew1Whoy+W7KzSVVtXMzA6yPWnOgT9YbkGG1p
3e5EgxRO+JB0T2fe4op6YU0iPtEJweau8vyoqF1mMgutbdIicO60u8GNIh1tZvZt
qqiOuzRIk1o6ShbgNLwvF17Xr6Tpn9ypghOcqYqP7/4bO5xsixUYHbGTgzsxxKUm
gJS/E756kXr5d2L8IEcvDY9bxDRg5xUBdjv0gKMDhDT2uPk2lr1c8oZDOvuEtcuH
WabaCaff/IH7mbdfrKnNzhoxhICrVOGUfKk8pCec1p4d6Glwdat3K2jPyjZCGtE1
iET3QS4kmm5oEWFzARbPuPkHKvn3/BzGl1wSkfkIjACa0vvgeNAEPokB3SaS7UHi
akwEJN6RUhbDQ0x0b32ju8V9UbASFpde54WtGtt0hAE0ylDeRWV+9mJDk+f3XklN
CdsInWKi5EXQvxCRGhxTJ4D3ISNIXaVhWcgKYQeYTAmSP5/G8s+meqQTmeHKDmH0
Tsd09OhVnqpcNNLFfm84vskGg9Sr8P7+tQgK9CQfQymTaB63uL93w+YhEFEowOp1
rg1/bIW90xQOtjj+dLvnA5MoVFQOqIzMJWO7EjT/a8sPANkNTMumJzg1uDutAJZt
E5GA11Gd3tSiA0RWrSE+7xOBCZlb/vn8Ks1MbpfAMCJuxyhBym4Lgb4mgTSYRsEx
/IB0GpEtlN23fPMowfewAVp8Ko5NxH5wqIXk1XMuGpbsqhvmKF8MizixDo/X0dek
5nz3/ueXFZyiSP3ufHB0xiLFGcbBKPfZcsFQhmMoR130qmk03IPepyPt+ERr59ci
uB7hjCe6OnT5daJHx0CW1z5Smd6Y7gmNAZvHJjGMmyBptuAnPn4ozI90GF3/K+ey
GBJP/Ou+UJPID0ML4deUYVZm55wcCoa46IzXlJ6iyaJVzvf9oiHvHQeT5ovTcGls
B6zZcxnD/mXHRUd/hL7bvOMqnCMfFRV8pEAtCQjbESkTf3D3mIcw1ZMmY93oUTGD
QDl7KNpq7HfB+aAQ0Q0jFThGh1LNUwY/+SyW1zwuJlcHsaIoqoPIvthxL8rOx/Ta
PIXLxXmMlE3PV4Hb7Y7ZyiXloS7ApRFHo0A1vY0V0msBXghVi+sapjbQECLuU2Wq
GsAfxTpghFkxpOyq7eRyqbT04S5yy8paeDS1ZygjfQRrkRBZsomLPCrnS2f+pVx0
jLm3KzdInagI8nx7T+/boHwM/OnY6kHl9U0VErsq940bqKAP0HwkrTrtNbSIotCA
LM6ZkH1nGK1MV5V4S6jsOrvTXjGGhKeYQ1wIvf94yEo8pwswA5MPfYJUtP4FvIRd
rTa7RE8+QjujE8+F10eaEglrSevHWbdE4Wo1AzoTqajp7iuLVIg0n+B8ITGF2qh+
fG3/0cCelzfk3Nj+kNwQ0/xYnQ4baNOjP6MJcgQdjyospw/Lnv3BBPFpiQUxuGzW
j/O/LMzcKIkLT6OntdMp3J9wULuXm7LVempFQoM3AVwZZpV0ovJzhr3w/X3q1hdi
9vwwRLA+RKpZFEfwJufJOscxalWOWn4N5irAufm3X9q3a0I0btavYq1la3B7UNZF
KtxFBEFQ+MVdCJd35Grn0SDAvT7tDOOEC0FNxuzfSXFQDr9d/HlL11baGizacpWj
nZQugF2fh8Ssg2qvCZiFqvfmb4K1OL+8JQj0Zx7AVFymC3OZ87GJ2kAjwSlNi3X/
gf7DNmgXG6d1q61cNag/eUOTw1H8gPB2341w8fa/1+wOVkYij4EdmgBqn2XoW4Mu
VYdBGm+XYcMLnxGTpVhrsX96tjHrgGV7ZY3Rv99iInKKkJLOvmdUfwD6Z6ORnPuU
hwnZEvNEw26z/+lWkrNk54J6rAc4ravVO57nMp0R/ZpMSmqMH8ofRpvpVuscYekN
FjeOYT2giWwsZh2mMN/rzDHKGTUq9RRcRQlkxGzEkCn3ki4sGvcoltOvq94+Pr53
lUQSiwNv14QEpYghmu4Ub1lIyFIDYeLHuEW7IMchO4uQsQk+ZVOuHBEgm8pemu39
qO0JoJipdHLL5Kpit4YVFHrGp3VzDzfuIVyu6kFok+ToMmM8tEMRXwbizDTcN1el
g/iPluTBIQqUSRjuBWFOnoN9ft29qCiIP48n4ECi82WTLpmTUrlxLhoxF4ahzCx/
9dElNY8etnMrY4vPZQ/F8oux6P2/r6z7jXS8WmwD2czHdxJ6ALyh1jb4apv+MRiC
NIJCDICsQrOrc9YV1XkzdeSj23wZF6Z0L5pB7QScgM0hNVqEdyF99QWuqfdCWX2D
0+7YhRWxnoHb2d50BZDkL6oUV+2oWjB9ztAuWN5InJ+P49dsEJTjdfvafMKC+9/q
vZeKLINiyhA/BqqwBYDxS/rh/fYQFu0w7IOEpeN8R3ybteZLPvj+5Pr5o/P1J+yt
J+MKkF/mPLYzVQn9J/ztvmueXd43A3KSLT22CvG8fTOAq/85TIV/iQiSiQU0QGK4
xer268/nNjRnizSSL1Vgv18emD+GoZMgeX5fKsjcBYy0dgxd48PeHOGC0cLoHOy/
F4vcSHZ7Gy8vMbxa/ZNdmwd/gMrETVnrKSy5VYpB19QDgVQ8QekKJLTEaSV98Rqk
/A3oFM4T0lwF3zEYNARRvuwDW590Nknsu8lXIWr7cmG54vujVNO3/+7F1b8Fz7VI
eGQ3qxY/D5k9mpaD7IQ8+dsZlkY3Ji8N7JgdD7R5T6lCT/FYzXJCSOMAYVvjySp5
hpHD6t7trFumtvHoiyI4zU4NJnvsfddnbU+tBi54TTeCTF5FRwQBnH7SrvRnxrK9
DkxUtu5n3JAlFuJUcA03mPpkNoPHWGI0ezqKeBf7zjlYAvlmyZBZwhHlhs9WnRn7
lp4m03qs2yH8hQ3mSPUk9jbaoF+RZnz2Fe77pgO3/kbXmuHIH8T0vwvIbGzsFlFY
Tkl2OR76T6cKh/sHXeYmBdybyW3DsdpUUAVxtKisywByjpYOM3oTKEUJP/sLmlZZ
o7JVi4WisLCR7bzsYt9XYQi3BS/0lUx0ZiRbJ+7L0OP4hUHtzElc6wcg6NYYy0Ny
wlNsJTiluT4E/Pi5SlNDbmtB3rl35NdQtkwKo/M/uBRQV4mxKu8EuklLe/5cP3Oq
HpBnAC/1odnoFcVYGqfnqkAicl0NBeBnGJO1SBDVTKjlUqSrXEJ1792NOwzvv0N9
yWpAQN1HzpXBrcsjKEg7ZF7X/Ozzg6vAM8bP+SDGTlPzZvdoXL6CCEFNeXWxMql+
ThDetgqjRBSBawP0ICt3E84e/1kk23ExWavj4nXNaLm5cHEFqfW8wqakMBBvKKfP
EiHi0/4/b5Ixme0Zk+hvOXhNYnRlFSRzaMzIBWstSNa3yHqkxYVbvueLS0P7Mv8Y
m13RdUyKSk1EHMP7D1vLMpOGKobHrd0PoiPdnSoAdrc1qdpy8lqKMP5GGanUhi/p
T5oBHbpjmGv4TGXdLKaIAYRkshiq+N/xtlGXYPVZRrCyNPv+OGxPKWIdH4pCdaWZ
CjWYRAyCWP/Q0ejSZT/4Rp5tN25hkKo/RCRo+uOtxG3Laszs09c+IJxogUdMc5/j
csW3y1HsSgv/NAwR1tw0+HJyigypdnchUpDuRw7wOEB3uGtJWsHSVTBdR7kvK4JI
RkrwZ2n05+UvodpYQbP23uklHMFvrl8HqZXLA6cA3W6F7blQSmrzSXn91sv5aLq4
BIcnJE6LICaoHJ50D2Fd7VmK54/Wi8+kb1j8MMhD20Y/lApaqk4Gb1+fmj2Ckmon
0t5v6doeM91SG7ddvNzZSLO3jk5n4fxQ9/Ddf9nmpsXXwvZwXaIsVPJzoomMNPFp
5/iNbFUVg8k2wfjzVqSh6Gyn5QadvCwgrgJOyxtSM5NVNxce3RIzn8nn6nz1UcMG
Azp6OyKIurFk2hDLBPpAiAtxrah8R6A2ITv1lFyVypLUwq3fHhnMPHgm9QeKmElA
h7l0qCGqgwudmYWV+696pczX3VExrpi4ktxJ3SbAgkeQoxSvGjz7r+kARY5cJ76v
q29GW9er19+/bqmNbcTYd+5PgMIjcliTf66AwGdxhd+2ZKwKHwmxSLPK4segMoQ9
ROBgcQPdgLg0Bu7PwFhStybXG2eFQhk+I2L/JKlCRN0Ny0IhBeJWX3K6v3jxo7uG
83JtyyVg2u08pQfj+kVqA1VfoJsHwFhAo/YlVcu5OQ/G8l+R2ePtktip7DYFIiqZ
U4hkdaYPEe8I9fZgRplY51CVDe8c2iQ/V/MrlPB0svL7l6Nv8DPgP1jmDinGzzEL
+nmjKb2InLnK8fLE7Ecv4q2335XFJs7wmS3rfkHzaSskUAgbeFDiXOyjGsdhWXza
2A7vYokhizde20uO9PpoXKeNdI+sMtIOdmh4g2hkO9UV/3bN4M86MneeDtJ3L0YF
dpTj79/xMOZLU15GDThlkDgL1pfAE799pGAh4RRXMI1ipVzsJzH6oDbrZ6QKkbcy
MKM5moLY+NK+RuCRn4UpZn7Cq1amQ1Po0rTV8g5bHitFCjzCMVealmfnGi4YqQT8
3Xllp9O8Y1TW5UJyqikZ+VyX4JHr7P5SeVrYGBewH1dC1yWqC4EVCoZguHxmP+e2
BlI8CnI01p+O9jJ6vuiOItjUdZzs6yqGTamdZuCgOu8bK2qoSoHmPT6bcX0kfj5Q
GzfY8y7uhQkYJksDvHVr4vzyh9LpSqIHnAzBzZ7x0b22kmMwhqLRzJH+td7eHFQQ
a+yb95OlyzfYeS5EdiXYH0ajvIp5e/CrNRJnG5rMQ69dutrNaA+rZCtfjdYytu+V
EEUaOiCQ2f3POY7X3X/yseKZpDEPUqa+Qw0AcDiT1h5MelZV6yvpUL4MSeyQZz+z
+2IgH5f8HRWxUJLv/RYfJ1ga1nHcAhh5wCZaHTKAZRIHE/dfXFEhtdoYn0+1QIAH
Ds1tgjkoCj98C6FNiH33PSLgSjfU064lcygJC4N8Lwhtg2FjeAhc5ZnyNA3c89ke
JgfwcfXHL4hgPfcxaohvxENcNBRPJumdByLylENo9aO7VklRGLPArKkKm1fHyuKa
Pyi5KC0krskHt1t2LXWwk6uzravfZC5CJz3ZDIIXvjCHqWQmkqVsvsv19YAbPEXN
2qVEsNnDF6X61ZF9d3gd+6HacFl258wkoe4XzpGdwnKEszTG7HLGg4cNmzPk9f4y
dL8GyqDKSWrnuBoNQPkPzZQbJaIndm4f/QdNWC4+cGNI4WF0YnhO31Z5YOGuCowc
ktBzbrpuO7YPA5HOo1K3YRHAuBlsetx1U324ad2uphH7FChp3GAkThtXQmwJnUfB
mEWTVMvySkLabxiUobzbJ7mTJAzF8vLbBsf45+DP+vBOQBHRiNdr6TdquEWcDy1W
OBSXHijHQQ64P8Defyoe+JHnkcgzeR+mLgDC9g0OVeTBs28Fpfxdl5LuUy6UBV02
g5/pyOECFaTMw0WeAz/l5/E5qg0q6enhfofRSizCw8PSMHwNfw948302KMBT1TuP
42CzEjIXBLino1LxDld8fmmAQaHiL6ytnMaVXpVIKCav5kZ8AgoqdUlRkUl1cn+t
DVMFjUJ1QNkJcft9/JmrLcsrnddtcDJBrlqMfcrq2Y/FFLytef1Br9NG+YQxYuRD
WyW3tbHbxEukaR6DyFtQHDldNfLtqJiuRjRg1UYnd04idlKh4LyvzAEOHUAWleh/
esakWH8qtimnSELYP0O/ENfibM6fiGs1mD3MDzo+R3zK5WgLDePQXhwVs4i5fr25
A3x2Sz2oDqadyK5rG6HI7lv0XjTuI+yWjeB8xOefR0Jwk9D7qpc0elnaH6hqIB5/
R02GnGx8BKolWvIh91TOzOCfOez0OkHpN49kLS+65FiyiSCz3y5JEPukzlTou6cP
b7kO2JzB4IJ2abhiRKbNESRhRJv8qiNBoE0z9BvZqFfdH/INtNBAAOyBXOg5QAu0
dQZvfQDsF/mLvwi1Mr4QRFnBeyBpxz6amWpYjI6lauOfOJWnvBH7REP0kDPVMxfK
cIl4WC95d/7LqbynL5qfZ+dfWJkYCb1w+ViuuuLmGpZdCwLJeqJEHAOL79xfv34c
CA9IbAAUKzl2K9/G0WyHCllkaD+loEuoF3R2jrLul0stBJiDmpmPAokURAUMZ3D4
gRgAPnL5fOfBjXZN8Ipln0K6doc8YK+RrGTNkqTvdgtgEvCQbQokcqxMBZBohRPr
HENbq9xkdZuIM0W07j2wwyRM9CUW4nJAFotvjMHTffQVK4h43nMIpXg/3rysUon0
CgHy4dg/1ndnZQxU8B6TA/9TAq0KAA2UFzdLJHhVZUQu0Rl839RQxiVstwCoWMq0
H001ap5AJjxaQB7As9/CN6o3Oyf8xBwUVIWqL4Jic+iUdjnbiPeYMCa+eYTX2hp0
b91zZjhRDjMFFiw84tHyQ29UbUBKp5qEkSppxxuNxa9XPQdqsfs99ZRsMOZbnG/c
GtsJkbmGcCkq6INV7LdRbMaoSaaljEjzjjrC9Ka8ZVnjqDs2N79o8nyOmEO8RTRu
72hDohEqVp2tA/KXM483Nh9x9ANOB+bc1F+Re30ZKnfUD006G5M4YtP4LwXxxil4
U/Lr+a13PXIMQVSOygBsQVfpRpggXLJK5ckq7ATX0njLtHFhY+pkHrcv4kQoBsKU
GFWwmdvphvqRFXbiH64l0WO+sIK+fQx68gwb4alZC42YRsPv4ZaY5/acYSsCILqi
2WyeL4CCAHGUG/PeWnRXNH41JMLl0revAgxhhbKyuxD+kBSeQUv6VKlIpWqM33g3
3wy9p5e863RYUgTSfdJ9xBhngOi+ZHyoUP9jdy6U4ACMJ2aK3s/m9Fm4I8dO1CQ4
PfBjLC0/sDedtKOt2YPZvNuW20SCRCpIukJRtg+LYWhLW2wVHGBXdb7hF9W6fA6p
Fgp6IOhdxJSp8oT2M/S3D/k1122dUYR7FuM1MlJOqVWFJ9B2EqxTkCMYDghNVAER
7e/NMgTuT1KxVfMZaPyaxO3Ycm6k5fRHxAFJoSRNoJiCmtf93nuN+4x/TulhAT2Y
nfKrBVxm2pbuZHAjsiUAA8vBAbc/QHrJFNk4FpK7pQO5Obax1TOX9+VEuB9F9qCE
rSoPTt3GXr8Ksw5FpOEcgrpuRvrHhss+vUqqvnbGrGbt6Qg1th8jPyZe9+T/bmwm
Hf7Z54UeyiwBWrobZX8jDuQ1nmEsEw1GJqyuHCXnSC2v0OqQ0g94ukUvaDkOxYp2
Zwxiwoy4yawJ7O0LSeP2TVHtzkFsQ/JfrObHJSqbSUOin50Z7+C9YLKO3l/112RQ
/qs3+ozNZezWcyNBqVijCet/x3KzdOVoZPLZ5LGAIyEvZu5ee57uQn81ieB/yDO8
vukByRNhm0PlCGThxWtyHz7KldY44UwCZLrrwjwP8/LM7MwaOLvV4QDq/Y34Exzw
wi7W2daDhptz/8ht+AJEEKAG7Jovm27BS6//XkssZy9QhZKM6qZuG5dtGcVTagE5
esgs9m0AMJ2k2QtMlQqj1k9HsVpdBn6xTZDkcEFrNhdkXeqUrwVoxHrL61AXMM8Y
3DDXUv+4laBWba+6dPR+nMoEuLm0t0koK2kEVa3lFAwVM1UzdzIMX+reAQPC/VEh
izGrNugz2tfi2FQNtL1CH93V3FthjbhPEg3Nf2aD1eE=
`pragma protect end_protected
