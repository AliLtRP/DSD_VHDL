// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
FcLXuUbBnl6zMvACQnUv9GL8mRzbZ1FktVMUXWhq1snDrdrF0efVpZ925QsE1Mi9BMKOYquFUXMi
cZx25PqqtRpu6Mk4jRYrXbl5hyZGKfNwvkisiJ0PI9NM/lNLxjam2cZt7HQjN1x3OfqADPdiFTV4
g8UFhqQYgp6QVE6VpZYclc49KEKb+JxLI7/UronjNbqHueYvvgGCTePLolX6tdLkoyIAh/n+6uwI
ztzz7XV9a/OG0+KufPVOOkU9v6fkBNk2AOAJqEayTXf3TtLKScD3smzqXbh1b6OBSBywas5u9iQ0
AGk3ki2GYyic138Xl4rr3onSKHgWqwKedd+9yg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
GwT3Ibd1YLhiIR0nsyFIAP/5TJDqJ9baMHzx7L2SYyv0PUlru9enycX1xsPdIdTrJtIgyV6qhC7A
2omH6L4zgNhP6GkER1ZFzG8EpQXueywXfxxkfn8QoNEZoZDXmCFQ+hQLUYLO5ivPMaLjadEC5Ycg
wGkL/EZxP+iRglGauCp3z1u4wnS70kosLT48IF8m4yR7ghfnYXRTc9zkXlqhnO70+31xaxPuxjsc
At2i+Y9HXMESAHRY12/DbLvJ8r1VgKo8zKYAeQXi6Pt6kouIVA4ZGJ2gSYFT8g3/WESutRTgpiyG
f9/LXVmGRLvdsU4fJRF4I7r2lgxoPuXMqotbPi0RVzXtBgNQedh307WF5USta5yyRyC8D9de5OkI
x5q6QCbkdluHQCHFITRqgP8UqPIpchINJwdQnsKm2J6faPqZ74g8bBZ9iwut+IPA+Iy3MpZohwLa
EdEoHmsWHZrF4DTScpv9Ul8i3gnLH0mrhNorzwdCH9/xNq2eu54DnCq8LPpyS667t62r1A8E+Jqc
0kUoFhRzMFPfW7EOeKSm84lbTC9poXb3pAwhmd91rAxsZA75AsBTFscEPzJGEHGKigK8sMLu19pB
Q4WXXAyuo4cBxpU9VR351njLN270/5Yin5nnf7yMKUVBtK60xNkbkOwfS4Fi42IofvJy13UNfBgl
I8FrLUAbIzAIMkX8rFPQhygS9E1IIFJBvYW8CjtlWTxySAILSWTqkylabUhYtG0Lnv2PcTo4gO6h
s6LwSvzQgvdicvYXCbfjtECN1dm1qgsGoeZtkEf5QCRj5w8rXmNNV85Ft+Xs2CmYvMnuhpXY8k8Z
e9n20xa0dwr429QWeJPwGtPQIOE0s+a/Q2uMnOQSnvdFxwuUQdfjKu5Ts6AABhTtLhWAd9VKeFsg
xJDnnS6CsmQAp5A7d8jq6waMX3sTn1xAXmA/H8Y8NuXCpfBfjX0jyX2x77gGwf0UAMfUTKzz53Pi
5HUIFRB0cTLOSmid4DMhjzbsIkZgYFyGgVA8JvZ+v/4YQNLUqr5mftffQ7ue8lbJR9BQ6zKQuyfU
EsRUA9jS99zH3muhHXZG0CkMpO3xTqW6DzXUjXNBLRqBp5kHC1/qT7aJ7rRISGKdTkcom9GTeUYn
pcpsBzlmlRgZbJNPZ6nOJCHSkB0opo0TriPXpKXRJaeyNno0oGCSAoDx4VOfC+wqLWmgf1HKvW/v
tRBkc7ZiXXFTACtIIMmthRC+R7wxWLiOC63EvCxfQVe0tXCe3HRmLY9XRoZoq1Bxx7rEvHb4mQbE
1cQ75JgP+hGqBQktAnw2ItoXkFoJ3JDe9ZjJVqxpZHZCSmkp8BfeIsBEvLy5sGDxrEHmdGOvn6PH
uWOabS8mSzZHWFONjQzZo2zh8UOsPX6u2Em26giDS/av/kRtujf/IGgU9JZd1yVTSkni8uPcnxze
264V2ZfMs44xNSfRDFUxbb25k9nhR7Ydh7sNZ58Tlmvtfs+YyBY38kL9sY1Y8C6jC8bKVO7Pov6N
kBfUs4hZf0anNxAnl9PI4XQHPNyPsn/o1cRFaw5NRD6+W/zw1FLbe09K3yPMNBeJW+p9zuhij4dz
Tr1bcrINdKKoAnY7N7yxTy9MgDqKDU+QkZhEO1UCc6WWIXG6hKPGP8bum/AlkOCz3LF/B/LWmtls
08HfVejqqemYvpvlTAx4EuMV0Jl/J/odX8aF3trQS1ZTFbLE9Y9c9nIRFR62lL0YM+G9dHRRwFpf
7lwfb3GWUi/X7EBqK8KT+PcB27p9HakOaJYN7nWdWtOP4nPUObae2oE7R5ZbwZ93l23EGrhcknhg
O2yM6K5xSveqD94W3BQtYZ5hUKtIuB3q681vGUYHDquy27skObUWelzxOOE813hMNkNPG0f7fK8L
1whb5xN8J857jaGlsOvRTa/iKBKRvlISlSuUpoxsoUgDjTINmRwbOas4RY6anMBpZvZEeDvSCkpB
9cEa85qNMR9hGPeLa9ycEjwFXrhcl2LhwT6d6QcAz/vCxFDjgEIvWRusLTGFVhdbx8vwa142ZM5Z
1MyYq4vl1FM8Q3HU9tiQtlCvZY7vaZv8eBlbLyktO9r2qWqC8sIdCkQVGIrKC44jJmz5PM+kiw4o
BcBGUhtedRj9pJ2dVaA1THDfTb6ZNBFGHVzy0XCqA3U/jAHHFsXCnGAoLmt0g1yqT/HBu3Qv1kPc
R9HjZCWsRVxydZBlqa6oknUaQOthYVOgP7q/qqnFzfIgA73wbI04sDNxh0tuQUYm1j5SzK7nwN0R
3Xbfdb9H7088D/N4cuA3R9mEJVZdQ68F0TmjZw6tl6C0EF45FjOYWbx3aZM7W8tcfkfNbWz2QNKV
y4ob05dhOttYYuRN8HMYRB53+/1GTv8jAewqLrq3QPT1a/GNLB8nbzYW2fMclC2WF1x+wt67q5yA
tKpvl8797T4cDcER1zvXiKgc0Y5o9VGaR0rrRUiOvN2LJi1VmkCWIf9xcTFzaBQ7bXmUlGsOKFlB
kOEs+kw1+umTsyaRJ9EnFF9pt2/M36O9zGkT3BBacixu003Vs6KWEXKFUQZ46Z840uv6HTcC27sf
MOMAkpIvZuB30Hclg+RY2+q97xlaJeCarfr7vkFHAMNYLiobr8edYrYYNI2JzjoBNQ3zWmm+pCbD
fFheVMD5ooc++e4d7vq4ql9yFzbAKzyacgjYN4yJbt4vlJnYmo0B2ng1nLEMX/AFjttlne5jz93p
5YkB3gO//qK1TM2cqEU5RhLnFZB4Bnmf8+YvN3TJUmY4Gjp10BcMEJuR+OkDgkG68OxTsym6aa9V
Jj2NHmQRLPdY50bzK+b2ArfuENsNA4/dzgcr8pmlWjoTKdhhznfTVdMDsRScG0wnD2Nr9LeelBS3
0AgHuLOroVe1muf0SeTkg5PLFYT1iRMrZ48VU8SsJ8+iu7QKawKKCV9qhcyizfbY7LDW14Lz3HmU
PmOBlqtk7xbxO1VGf6mePY7NowF+6ptURNkcyZhEG1/qTf2lXIQxd7LDYT1KNtW8DyACPjYIaZp1
GLhWQR4IdQFifwyUdjH5w7V5+hjIbvQ0BgHG9ePGipQjP4y2AJDbsiFqQugAQ43q6ZOiPQhxgjpV
Le0PL6jAOLI4z7GXcccDRv4MCSIaTOcajrPfXqldhQtRWR0xwE7r7pIcffR/RfOytfOuVa2P0Hl0
MI1wjV5McdRwLp1Knyhr7+nvG8/D6J3Yweabv4bGELdUZ5sJXhbgdImUMmx8gR8pjq30g5ZqNm6n
/zAvxL8H6Ciyc45Vtm1ExPckFP9jN9dMD0VJOmv7JK0RfJhYTC8xuagIE5b9Xa2FkdrYSDBr2bXI
ln97d4WDHkylIHd/5KNw4MkiwL+ZjlqxOoxkyheJXfhCPZya2OAZzR1zmIFinZmYB8s4DGlCiRep
ryri1LSljkCxN1PFqjuTDEb55IWMXzO6qmCBHDQUXsCndWpk2rPUE0LDMqDLYYNRcLKr+7QIoFAJ
+Pt3+XW2LuqIdxfuFBIZ+NW3T/UFyFduT55FHXuCKpFzHq6ymhkthvdIlgOP8DK7ETX118DKq1cL
Wfhl3f9ousZStnyxfYmiJklIExalix2l8hMAAckvjBpfRJTh5CY76/fsoOGLsWxiUmZ3RJ812teJ
zaQI/EBGKZuZlMlTXR6WJPO8B0Rk3TVGkVTEsZj7qd03e6uC+7MfA96iUlibKqffA+OyM50BsoS8
bi/5C6hdOJmCh8T+9HPgChKy+dkCd8rrKqFdv5kg+eWYaUPnN2sYjj6AAg4mBQ1jApK9zwWmO1xR
zqfpVdKOjkWcqcf5K/axdNmJj1qX3vov2MudttpaV5UE9AuuVq8irXIjUxYA0sdxHp4fRk+XOwnM
qFMshUCCRimxvpqMe9Ih+/S+7ry/xM3X7EkrvvFotOlBanA+9oA8uCSrjOWSIKJqWCEgcCnvUmJo
HoH/3Sp9Ktdnxsrrt3z6/prwAtFHAtnXvj9qcdkIYmUrGon4KJLkT9mTjL/DuysVQocxIcc1t5Qw
oBs+8IJp4oW1hbP0iJmQ6aufTWwiNKPv4VHFuZi1P2WoJyv3PMs6U3t1+V2Q5tBBz4GMfH74Oeym
IOOw3dpt5TJGb4+49iVdUMO3aE4sKdBIRjmfweLrm6+yNZNFbVjoy6Q6XRJust2b28HQcMbmB7Ds
wu09cDqz6YCVyWCwfTQaok/W5eIZ0P9rYi6nsdjyd2Qrdn34k+/OBboFff7mXmejOc8Wv00U2Tbm
9qihKTxV9Fa6OBq/mL1JFHMbY+ooOM9wW5KTXTrlEXIP9Dujm9GejAOZAu9WjicDOnefAmvraiw0
1ub0c0N8aPcgdZ8xiDTMX4BL8v+emSnpKsgRTIenHocfKDnX138XQIC34ROLW4DGA3vwwTBG999m
CSWaOpXfT2Qq9aMJHDXUT41HsRWo4RS88kERZBotKvs7JPDOyLq1YeaSMgBasXurFfpV8bm1aUmh
2surlxK29pBGCJDQ3PXveuHhy6L+yMescMfBa/HkEZjC3teS8lHkil7o3P3Bpa92sZGQJjRIDCMH
pUtUfEV6NolSOE0xToI5LiA+Cpk2p3be3Kf8LUeddD2YlQjyWr3SKhHiwaIsFgrL95Q8Ht/ZUNlV
K7CPs/b4usrkDGIiH9H6PYz6OGiocSWI8fhJHwQvZi6AeCKlvUeFNilfv0hqh+G8bDHuvSBZWott
+9G/CQudKY8fEzpq7/jEOCL7NjNNP0yzYbNK/lLmRP0upmAa/h6a6Ik9ztT/MUBLv2e2zR8Y+YnZ
ZVgakk7b3RGl+HSAGgfTTjh2Z5FkmjgKm1E2Lcf0wZRCzw1ZBScJBF/uyfZkzcG+KUfXsgM83WEm
ACfsrokP5DbUL4yFKfAYMreEUCNXneVTD73Z2EiHis+2TE4pMAuuU8VvTLUxa4QJsLcxEIO+33UD
bmtp4eHJ0mu9VmALO+h9wE1HCxlYF6Vorpn5oSpYoSJOO96rmICPscc19D7pdk5gbUOko0U6cRyL
irfdQwVksjRNCjgSaG3agRoxbm3CyPbOVGpdlRMT3RD76W9Y4jdv3mjqjMop+YGSz/zztgTYnzDV
6mmLzpF2jv+F8mKfG+a+smBrj30CyUD18396xbr6aNeYdSkno9YNNmxyD5eHeDArgWtAo8cl8uO3
e7tzHAcbnTqBKGSR0F7eG8Xpt0Bjp14ymLchHuCQaEYc2IMtftswLLL69M+QDn4gGIsK4e4Ql1sk
R2gxPfynOeZScCYa1KRM4mU2eIhaiFZ6KkSWgM4xrQnOHSpkvsCyxdFGItUrqXez1E5nDOR2gNkG
aIOV7OobOppkoqF3ay6IXa44tCvqb5TbTq4YrT5xm2S8wQu7t8itX3T91FTMDWU1iYGny0O45t7m
1FIFtUm4xu0Bxaz6qDg5hguxRh8fWhfR3WzhTV/UlohK3vv5hnruH1hqWpjYixJTZWBaY27RO7J0
WtVCZfGCuNdXgC3IbZ8TQ7skQ/mE3m0B7xI6z5TGrNfxX3kP8KBdwHMPR/m9T6tVTRQvOApmSHin
AbC/1+KWDyn1kp2EJwdFyknMOwNiCwclA89oWerVd/1nYYnxT6mmH/HL1fiohCV0DgaaZGfvbwX7
ga5uJrK1ZrBSfedoQ96xKMw1KO/aeNbJrB9jGE+XTxzGb4yfQrIhRIsabmHRRBXUwAd9viuwSPrA
nBzmk7SZCwd9KzmpqIc+6oLIoYrUYh3yBYX6mp66XVI7ZPVYKcAIkzgOobM6yt2OoKpXTOjJwZ6h
43gVjef8u3PivqxaSoX6gSADhBbUsZr6E6XIYEoApeNxdxGNhSAfVXjOu9p8xf0wwZpelwDm3cq3
VO49kkKd4imXeRJfsXdolNQYBLN/uGuIKMmTvrLena/guGu0VtM+FluiYz4wTA4M3aAatFLx6wSK
1whY+KnBp+ErG2bVMnGCWAQvz047cdF6dWt2kW7dkyYUkh6ugevRux38TTMBX7dq/7yAqYCWjdps
uOXX+NdSBU7mTFfM5lQEBqkrQwxw/tix9DBVPJH69ZUL3qQjJEmZdizKF/YbU3P4DJSJop6H72Tf
61k6BZu9C2gQoKb207i9ehY2L5JBncMVAmoHnmcTFpHmlRPIAIsiZKf1l1qg3vgZ/InS5+xyBAwe
jNFX9SG0tuKdrr9dgOIppQNJiPqHC2P38DmoN7lSyMC/uKphrp8H+DcF93Tj2beQ0H0ss0eQS9hE
aanqizXelixlOgr0+r4VHXlb4AoK8uixuMmUtAdKrvkIRQ3i54cZWaoCMPdg6+GivCoYRGv/sqsr
XYEKptb2QqblL38XMvWyZEUYxOjzk3g3VUJ0XN5yHECXgucBBXv/PE18JrefS4WHOCd6rzEnyGMB
yYy0gNrPkuIrYwZ2CoQd9lJ6VzAfvyX9gQj9+66Q9K6TjvWI1zd2RqbnYd+KR14zkcqPVgoXz1u+
aKIcpZfQMmer4s8sWRhMZ2nkQY4AHD1Ix37uaFXpHe+FYDOHVZCF5GzV/PXISiqgwui1ZdAztbz7
b0CnhxUu7kxnVUBWnTQuQ5yPLpZlUE2ECRC6QwjtxdshmZKIMawiIgAT2/iW8/yK7gn5gXB+4jsr
kcI+QnV7QNL1+zht19Q2wm7OpPy/1qyEfxd7NpJQQsXBPDYZQfUo5PCaYQs1oHlSeBaqbLYI7+ee
sV/vq5Al5D7nsSTFGsmfmldttFcm+MxYMwFxXKF0TlyOcvYHNh6HmK4CzfkbQY6p0NH6iB4GF/3c
5npCkKuKm7e2dLPlwPm9DF9BBaMchCJN6jwuYst/66G9phwXg6AFA9arb/zlTaLEd5hqGQpmw00X
Hlwwof/vbbU1mpViVKZtkmeHgnidTQAfNcGjB3BeuI24gidx9Wb/cqxwx4A3zJl5X5VOjp645/Qp
BqxUvWQo5lYzYLMfRB11f+V0XsNaFLq4pcvpWB/t/K4fPZ+hkrMLkkYL0xSh0aevyjschRhoyv2x
rA3U3zbwtvs96a2jM8PVflwm0NS5nAYSd5ets9qB1pxTvu8UYK7nZAfXU97013NgOoXce+LpeAS7
1JgQ4r1cwFz6diT0NasHgTSFUai5TERScrFVrl9L/0aH6tkRBU9kxPPS2UAF3NGIv5AznzoVNReo
ceY7eaP/HFoD4MNpO6l8pyILwuLteCInhHc95hs4rEdyBwbv+nPzrzwqk/1OI0FawO8NyTpYe6ih
GtBNMwljDSI4/LKO3FjkuREEXs6tw/xxwSlBjC89Ef8YoIInOO4I3fnXFoNZdQCBqeMC+kUtK88K
NacqGfXbrp1EIagG1ZU4oqtB20jFmqUtHpGqtHSQ5pcp/KScFiS9kn/SlcKtoVVHIO5GxmZMYvPb
FUaj3kge5Z31YpET7vzZcNJIn+Uk4bmwLAGN7To+1JWqnEfyDAy546QmvQaYfT5pWC/3uIlhWoPv
ePwex0Kym6rhEbWAzi6RqKE4/f3wAk+75PHssYQDa1IYmk02SrqZ7WYd18WlQYcxJURAc9esE9xr
br2dVVkvbygL41Ge/8GvcF9LJLYmTPrmexRCU9KRAxkDTzLAm/jgqR7neJYiwWnRrqyYWSPSRaF4
Se4RMWvPcmGkJZI9BZTLW+QIeqv0KYqN8Ibk/y5cLMuXoKeoyCCK/pYCpVgMkLPhvruF9H7cJ42m
2I3SZY48f8n3kqLEvwm5Em3/p10BzRwLm4Llj4WtIGJesisazviOQsVFpOrfc4E5mKvi/nIrQ7f8
6suwxSVTKN9D/IgmkLli7KT2FWTLJnoNl8XglbRlu+dhDhay3RW5rrm9MvH8LpHu/ia3DIsSxuVy
Nv9ZeO5unS7Pr7xkKyBd0cKC+GqGB4FQbtUEnlvUYJXQ67Xe7aUpo1NS9en6L+BQ3+mLN0YjbrKv
53qAO7PiYsMXw/qlx2yoTwAYeXH9Mqib7hmazavyrOO+wJnIFYW6wk4JPgO2S95xxF+gx9wLa7J2
MnVb39UeFT9kMeeB1Ks4eyOm1OqFz5tBfp/Q8yAnJGzYwM8Z7GU35QjDv9WMi817169P4vNbHr6S
P2PDFKDEj2OyNURJukmrbbN4vo+QrxiUci4LIZPKcmQweWABB6mr/qDKGbReXbJQRZUk6XQjApzE
Az7E+pLDjQW3IcNT4qc9NO7UT5Yv7sjwpJOWUwmEXwbfd9hhVz9jSr6LB2SQARmYyFqVEl+CzcEv
oJBD1VglkYjR8Udbue5xJzYNYJqSb6G3z2AD9hcFrbu+zI7haHUxHs2B6NAUp6R8oAYVOrCkQ1ZS
lc6DYpnYxU+IfhMSjxdhiDzMC0jANhqsNFVWGJxRtSaQhj8yc+Mm0hA9UfBHblMtXmqbqjhopTnn
UmzQgRN+7XdgkYUbFZaOmBkD0xFhGOWhDCijoBQhbJi+A9+hlExcAiDMbnPOswpbZlDUEeMLJY/W
GUXonlzWulya/NKMycxYIQYyZXQjEfkNwnpxIu/vSTDAqKSJu2xcqDd+g355eN+wshDDL0OOlZ8q
xtKq89B7VBx29SgGxwKUtGEi6LqoOuxIXW7BxFbYXmlJUhtHsOdLwebosFlCXdC+GvAbDIYdhxU9
1uGjme6kcXDmXsBMWN/UGz3Q+XHwgeo9dQVZeSAp65mebq32YQQ+Qu7bV+Z+ztnU72xsZaMnl9Un
x08nRbbJmwJoeJbmUHSzfTUw5iTRNv5FpVIv8oFxCs2YYCjK2fd77Vabx7xNdkLVmkyR1ObJ6ILK
0xPrhi3zsv8eNBXH6CYtI/A/RLGvcVBSdlkSUuFlRAjd46ZI8D20ejUCDtVEXyNx58FiPWWfvbg2
nZoS/tHwwlfpcCw9ivCnRYHqSYw4YMJdWjjDp9l5hVdMLMxLM7ckUt0OU27am7XT+a2wS1novVFT
VxFjrKq3/zQQzVaj29w1V5RbDmIJReQmZbpM7QBBqpRsFRO6qgwkIGTpF61afMMfjh48Qh0Yd6L2
7uIvdiqN4oOMO+BrVVnSl/Je/ObqgnITDwNvJZOvrNDFj+qAEl8BPiXe8nH0umm7mw3NmxwdyYtC
/NRKXyj0OpUZ8raDvZu4Sp40pwhTNkAWaMqzracm0UW2YM/F2KmTSRSQzAPAv1x7r/ipPgSBLwTy
0YzWrUXVY997/hTCqENLoijI3Un19PkU6znMZ7WN2dRDxxiljPmMVBEJ+eKz63Lr9TNZ+PbdwADL
mqYRJ3wkr2YNMp1SuRJLRoqwI8oh9439WGmQscMMbbgB6V+ta8jdGHD4ATHsPM7QeaApRTQ1o/FJ
6sMXXRTtx20pI9fyzjg8TKFLdVyU7KBXPUQ2eVGNtiizqTg5kbrlSUzstohpSqmZyjsIoz123hyq
K+JwO9FABSkHMhua5/nYf/kKmYHcXq0EJb2+zPq915zFYrwwBphtsQWe2kSfjLxw7LEnbUJNLaoT
NbOJw/4GchFVjidNW9aHqbUs60QpbFqARiX2qU+f3xQ22neg/vsW6RWkDF3zmGm/Zf21OEkbY3ld
JBBlQPhSPKgyLohcnGW8neYxK6/FIZA5cNL051jgbcA8cTA1zZgL+wsTpiUuKvtw9ztQEPmmOwlx
ob3VneSttHucWuiVe1WLfNzZttSnHr0a8ob6uMEyCV10xlakbE4kSHuyFDDkEQLJolUO5vg+3XaJ
NMT7bST7xB3P4BnJil1j8O7b8EZgbbZN+EQv2Xkg4lZtSexOkeh0KWNZ1NnRgMS8LPcr/xesZ8dv
Q9MthKeEPee9bcVf8AOj5Q73pgsWb7z811sdJznqc+135DjhoJP9PZXMCJrnC0h9dz35eFnORQqj
MkB84zO4aroAVkvBPRtm2H6DWCSCUnYDa85yK9nsqV0eafrOHHFHYXaREfTGUlECAOPvQIy/wQ6p
pZyzU9auDEUEiKMeYgy20Xtq2Ih1rMQdL3QhgDQ4fvsq0+ASQoTMUMW5DfqH+DSIxRvKMfHX7iZB
yXspK2/MO24EMpjQaHKxZY0fvlTcxwE6bxs+ptT5b+kwsvalynycnqNguliDJNB182GjHTVp1bQF
Iv3g2p+35kZm4tzG9rz3ib+n8SbccGEDTIZZG/OIyWupW8+jsRw0UmiMijKVKFH8G/bz1Qlcrfna
x+L+cBPp+5mAMcjBThFt+lp0MauX3zZaakRE2ae3xO01H5bCl6RJjgvBGd/Wt3S3t7TusZCskhkD
DXA5zBX31vK5+EQZq8Pz5BVoZtxkdVSU1kowNSG1cWkPVirJgLs5EAgNoMyH+sxGLhDxIh0ZR5Fs
Fx6wxQDRb7t/oqBhZvJAd6ZA+9hkXG84LrjIbd8YE8taaHm9iD9jC88i7zHpY/rPLYEvQOkjy+V6
XmSfLoj7FyX495c/DvwyxgvzRuQhguQO3bkQoeECmcehA9n5Iq3nFW9ejWm1EpnSfJVI7eCR3vN+
E3lIhFui8NRkmR6jH1nBR9flzUVQvHu4NKk6A63HSzBKRiM+oFdFx4yEqkoawB15Y6fV2NnUSCTW
XL9Y4JaQoYCF2kLDlqjgTK5CktRj3tCAymfjmEN5tK/B9rNYDky3L5HORkMaEeBpBGQL5px7V52k
E+MRTlMK11HJk1F/EXZPayqhn7i9HEfVEgwYN/wcbQPZ6IXEo2C2LHp3/wr5jzGw2TggJEQRc744
Scrd8W5dLDe/BqnhjNr07fYfNSpgrkCxG/UdKBk3irDfRKYmlOktIz8iM5iZ1QQY7qO9hg4oBf0R
LAx9MnUheC6UzZDiTGtI/mu+J27UWhkrbf9kfMDbFqmgIiKRto1d65Macj8mT30C07sFrIj0f+mp
GmOX3UrHC+d9LowfuAg1wwAC4LUoW7zFqUyHqu5xCZKY+eTCUhcBxI6iAtZ1Qr+NKqtqGdERvliS
AFtvavJ1otOTB5oK+D4GshXGNF/gqiLumqJJ0kBIUpNJlIldSISwq5bqN/007/aHi173gr4OMcOJ
F9AKJbQ8MXdsrw5FnSpqqmsbb4mGjIqV2QOI8qDRwpwVfonFkjSbSN9IPCBvLEMPFtYehR2KbxRc
QvRJmIpixwMH/lFc4mPtUbamqeasaESjb/sjHTIQXHn4HuLGZdZKHPoVzw7uKdSncVkmlo0sWjw4
UHxxxdPVh70tRDHCC4jpcTQKzlNHZOgJ4ofBfS/qd+nTSMpFW6WWjdS21+sj5OpKrEVG5dA3UV4n
yCRBJAYTv2hjM8X0SCKPxhQZKg6gB5caMJalGPym2pZysOIAtM/Dz7ryFz2GLWa7whSds4apMuH7
ps9fP60ABAqD9x44PXWztmpeKn6jwgeyMaCvP7rY7dCsCnC00PUCSclneAnVHItnzlmIBvf07Aqk
udDfvlIRt6gbgd3bG2/ht/gYD1LkJb4RYPAXXiOkDTk05eiojt1ZlYkVH2Ri0cyx3gcgJUkleKEA
0KJnao6VQQF+/62PcxmM2ENb+8VWxFcJdoFi3DydaddVbozGs+xxgAhETMn0H+5hEc48ESdZbURA
svzEcs5lblaRECQnAFVJwOHQJIeauneY0duooAPjTX/n4QZM840sDerbTMFl7T4oWzfYQmXrPcMZ
t0wABgQSFehlEboqfO+lHaftpxLJ1g5km8HSFiD2N1qr65nqNf1fRlY6cUC5dDBa0+Db8EtmJ2Vt
HS2V+iBgyBNQD3aovuu5ABrBuMU61EreWU5bsk/7tj7DYj5SfHltif/KfCbCXvB1ZJ97wsQCSCqk
MNT3irUdrFq0eT3FHRQW0P4g7e5fuIua9wkBwuCnX92bSm+l1GYmeZ/HX4RztUxhRdfHPo8dzgjV
DAVCn9tgOW4eOqxmiCv00aNl48cBYyXV+tq6E0/b811CUjWIoluY2jtUpy+nukH7hKcz3+Z/vhBp
16DbDDNZPiy97qgXaWQC+XV+j2sZHgF0z1NxL8F1aopJtx0GRAQTg9vCm02iWXXQJsTRgnUXvMQK
3Rwx4hzgk1gbZk+QDZxCPhWpUs5195y6qNBBDgvbDhQW2Ue/enTaxap/toj4amxFOElQ6g1KREnl
JyH+pa8BO9XhyK7WBnyig7qQw/73AlB6BI1UjZEnjsLSFRnW+302uGnXg9t58Uvnxzxwjwi4vPQO
6KoWHbUNtIpto4TlHTyc8GjvuJ+zGGZD6aG4xNEskXDddPPlfMfFY5uN1g5q4SG5oaqBtI6dEQCt
4XYAOyzP+TANAf8V3rlOddUyCRVjgyUyAgOL/dnpSNjrZjRnNwsHokBiMd+l86wy/LBLNYUX5jzF
ZRG6b860wAAAPs0Idf8G8BQCTmjinGCzwJqnQZ1SytNsT16/vlsAsdiqH/CLrALSgH7JVNqKc/3Y
EGh4q4q6ms+jlenu57bAXCSFTb/vwm2WQiEWOQIdokqdN4JahN+Pq9uy0A+lcVQpXDXoxtieAnBQ
4AzJDmvsc13fDtzWoLLPIcfD6+i0Z7NyQXFMELPOyeKiy9GIdEddzhFvBTxBoEsFaT9y/Sb1aIYC
relAL+vB2n44P4VzMaJXhx/5UrB3ZwB0PpaduCNdMT3oYaAg3OC2qSKew+OyX+Wo2yubRG2rhL59
xuLWJpJkuc/Q+jHZizwNhYNsynkD3+DiSE3T9DpsVW0R8db4Z/iM4eBAIP+/f5Tw5TFSjrym2QfX
UJw3aj+Lc4aD/AFzwgMtV0Y3pv7AIixLR3dedudchLlc+QxmnAqQuOHqxujmts+jkK7eZf+8K/zA
ihZWrR9yPMpLOoSmA2aMQY/uGUbLSOTnMLJr7qSeUn0nw5SxMt9ZRR+s1xrAM3dWA6U7TvAqIi8c
kGWflnbruqrmCi4N9JSUzmL5AFypIooYZoNJq4WiTTiz0DUIcpF8I7pveLJUhDAPxp2mw9u0VCWQ
8NYTLMHpZfeYoLljrSsxWDBBA60w3huid89MEqLxMGqmDnJ/mfsw4o24j3T7ox1R/KMfyQG7+4M/
alD/mZT2BjpaUSrEqKymszwqY/i5fpZdlz5+ttbKeEsNbenA9E+dg4x/LLW8ruwqJ0FOCJMQB3jm
CAy2Uw1mqOZTyTiqrMAm00dTx/9r7Ejv/NNHBhuzRWhXiwYwEulZvxNI3p9ToXcpXJH1mGcAw6Ra
OmOdLQZqxp+LRQEMDwkFZphlt/EaOyzvt90EPCe5D8cw51QJZVJ56a9yt9Ra3OCPg800oM34StBX
C55v4FjHvTDjb9hbRdn8fBIW/I8szr0p0uMSeVsbm+TP+YxNG5vy1vlysG1lyhho2lqp45T4HhMy
BKGV0uoR34IuePNQvReAEnbKQH7++VzQJlTOOx56Ms+ENMbimLRtBZVDegUR7KYjPvrh5t1eU1RS
i2D1VHRyait6zN/yh++VX0ZzqV5q97Wm8+0iJOXDd7ORMJFhVK0809BRZz8wvDk1LZmQgZKWBH/2
HHy1Sl8zSH9jsw93vXODMYaxr3WEN40lEocOZdrUpAyDNiI266jx+P4wZze4l0OcCKwitO9U9gns
Q8mv/O+5UwN6PC1mk+Co+bWKRSonydiKsnYEBFCiLigo/Av+zcAvT3zUGHL8P1bfjO84RzyzMm2u
jYky18rFFgyxmdR8EOWi3ZVFNgFcfFGrJCzC/j/u/RAlti7xTzTdPcKLr4WRIk/LSZ5yPmJaYNQ0
htxxslO58X1h7uFXXID8JBtcONLZVSK6nfZ3Oy4SxgL94Slbn0+AYuCjg7+mzPCNS0H5c0EADAzG
IYQZLZZnReMp59qXnNIQi5IsCw3tHK+rNY1nQVZJKTtxC0x/1FxKDegzDSibLEAZqhgIJKK+Ixb9
PBQSfp/YHhLX+EB0ycPo4/hTW5pROGcZHl5rvsu9xeeqCnx0MQCZ0cEZZRFBBC6JyM2T7Un7FsxH
GQBUbxlvb06ZVvP4xwuKbJto6RulBAve9omhjaaYNipPEl4+ZnqYXxX8DgRnCfiy+UWKzRkTu+X4
nPNDV2/2aVV7WfpvZnvTJJVY6eABO5PRU44h39Am32PRNCjs2QpK7f9aoMWk3X2017aMzMzV3rMg
VEp/QqyqyKT1LnvB2NaPCPkN0QsS/KTY+ZPHMUFqJfgtULsVZ8QZ8Hrl29cCT4nhivZXNd0dOmOQ
8BIg+EjN1i6hlQ72MmmRz7qWhKEUjumRVVaBgZ3aga4T2wvih7U5qZC8fcGFKjBQoiW/wTt5r4Xq
v5VR95ffSkk3EXmycb4tGBkf0xRWGk+Yrz/MlwXrSe2CpayIi3LyeQP8HyubK6brAXjIptlM8OOw
QHAhJrvtSkj61RPHdJEB9fYRTI3Xq1XpoMSniIsHpXdoTgm+XSVFxassvP4A/dwT25DKLnELrI81
hAih6QSs7bYxP2PAvJsT2u0Vc/U3S8LDSZ++51RdJ45XunKn4SiMJveaNWI5BZNTEPe30E6XQp7E
r2OHFrx+yCMsoG1v898Hc1tDm+npVCn+G5Xf3oJNzKyB9NQ3/xzAc6p3OslTqQ09KQxrV7cXyu4x
qIDSVDkM7ifW7EHHXk1ytRloWdoBJMH/qazEwgjuzy89q/CBi6Q9cEfznln0KJXG2nM2Rvtvyn89
Tepv4h3mhTKGMo8mTbgHicfcFnNLry0V5SkXqfJITW4kn5DTcodJFX0Eg5+rYMlsweEFP5CS1C3z
Tke/2P11axc98A/2Nsw5fhh9uHVPr0dxgouUI6l/fWvJVAZxk5dlWVGpK1k9Rdd8ViBX14GeZ6f8
OyXyuObluhBBhBcGW+24Izg5mI9qJg4+0tLW0aBN3CiiZc7tKvEuDvf22lbICpBRbaHXgIH2wdFX
GlSllLxFzdof6jkJt+EBE5UmYFSPZB3ER8ET0d+XiO8A3nXLq/NTgu2KrfIoPDu9PoNF95AIrhMx
rAamh725hQxuUF7FJ0lWmWsHUyUWAcTH7ZHhO+bJ10nlRsSCZkhQO4AqX5sEJchrgeuwlZguu0bv
VcNngY/5U+loRRpTDsqrGbZHh7RMJXJ0l8NUAU3NVoPMU3hoVcePYILriefrA/+jygGftAnk1Uc/
Gm2fooTjRc85Y0zQJtdVU9wiRI1IifJ43gj3Rb9MVjztZpglF1kwhsJrdpxdST/wsB1cTjjPq89p
C0+UkCclN1jfAHOXGhBvqHuBOq8UOFY6b1Cghf4rYz6yMmtgUHzjdOVia1VgNLromw37QMCUOQ7P
+0wXs+b6+izA9afwc/LzXu9Pq9P3zyfA73zkaebK46MX50KzkGnrjikrR3KUfkLhjN5PqD4PHlNJ
v/amrFrIIhNmRUreAOZyoGb4pD+UznXKfsRlhlQz7vA+IYdayydpN59m0S0ZRN1aC+LGFtefpw5S
oN6ot8fH5slt+aF64ePJuWyTiEKviX8F1Ocq6/UxYYGOpDEokJnf1iezNFx+/X6ToYSBsonzrcZH
8OwzOhK/40uiFeeZa+uBcmTQQo9k1+yn4eU7CuoGe5GuCw1YAoRKmTZ09My/KyyAV1YHjZOQYT8I
vwQG8gM7HGNHd7N4u0RzY3N81jLEWClHgGvmCzKEPIfLTnZ85bOHCmAGK0evxKQdGtvlPQSGavkh
DOSntCjoNtyOI8L97Qb6JuHg8S7AfOIEAXlgvhvNYmRyltZOj0wUZ+hr7+QZyG8EMzG203PjIT4I
3CbptBG9R4WDe0SYlHRJOQSBefg+QZdtHh8RFvde9uFz0EhtdbwbwhxFc5MjB2WaPqN6cmya7kCa
xs7knkX7jGix0syOW405Du/vhRqCU+e+fy5xEUP+MmccKWTtGVElvn5cE9Aox2fj+tWrbIChshhe
4gEPAgR0VciCy6YujRA8Xj9RFdqESvV6Tpl/6IE7jTFhCRHaScMLeUhKO6laVtpNoDHAbYoDZ+Ml
boZfdTRT9Z1hlB7AmfVqk00xWkEyGs4MOKVIPB/WS0rbtrVSskPGtyeHa5zQ+vvG+S78ID1eO0nf
vHBx3+idN5A0/IEEtZgaHNIlibM7ngMElDsacsQoxsLTSj6+yiawBgHilwsC2hZ0oZb3nwtcK63a
4axrx3h/liWlGWIYRYEHubVGUmElA86DKWG3ANx+6LusrBMFPwsNZTpalxqWRHMr8feHdrdXEo8O
//k2INGkgjkGluwNJ9o9aZ7Ad93gMk040fOZVSpeCu8nxjv+Qyy9ahLkO+z64B/k2c2qZKIe7fR8
6ir5LIhci6bJnLsRwsNo0jISV/rdRdPrgiReg00h/totFcT+LMOLflqkIrzfjmlCGgDz8s1obo2A
Iy/c5R938mAOkWWl4pTGgdDPb00xbvAMk3/D+U/Z4jNFGIzu4S/OGgwqCYykJeIFs3Sg9TbNwgYu
a+Xs++IqySzibu8+EiYR9oAv10HHbkIc643QJJPQQIyi72LGflSxl0kMQz1+oZtQ4Y8Fn1wZVEdz
ILvedIN/5d8Ucsv2snp+VtvW+yw20rDv5IWmxtdefju15benTxdD0Weic9hnkQlorugYR3OtF2t2
iFtYu1YUV47Zf5t+ukJQyyUFK9ZS8kSiDEVP0Oq/SGsdWbpICXgdBVPIgkXdVTVIrQzJZ4At728f
dkzOOSdBrbOggOq5EajvpWQhy4L93gP/x8LAAkDM8VY+zGX/r+8nl0Saxfdqbaa5z91MFUsbipc+
I/HmHORufYVr+DsaBSrBFBRN/rqOyIa+7apDyQd4ss4cgLhwFkqTOH9hpBJNYbBv9L4LmAv4nFd4
gbwDqLbKXqdZ4sgfjI10X3BE5y+zc8EBUrLkpmQIYbS7oGcJD8w+K7fmRPH0RwNDFeRJHDxRRP+Q
aV8xTXBF19uDbLaJr3KwX1x0PEuL9sMp6ljI+8dv4T5MS4APphjffuLa49seMNa8VatIOxp9CnrE
tOTI0sWvxS/6VUT090rLtFsxQhuPksJ2qv1psSUT84FUGPfFKOGHIFbeH3tQq9DPCX3aE6kOEE6D
KjRISMLYRtbHz2I5lzca19ZE9ZvJLNyenqQJbi+OFs7CuL4wGRji5TFoA4tn7KYsoSmiRVAGmBqn
97BycKP2W0plIIeHpURirzFL2e21FlNWNXDHWruLt9R/5f0wauzoC1k9Cy0z3t6lPUsbqnMBorq7
QjUXMQsYVNp3kDVKY8hC9lmP9m6SxEeOa029iexRZbC/mZh7zq2PLORI0c29M6N1bgF4EmZV6W1e
toMl9Ki9OhORNzhMSz/LRffBPlQ89WQ+B+8ZupdlCUlsQDBZd+tWDOgys0qRBO5utxbGdSRv08vT
ONNLVBcJvW1T8htg/p7c8UE93Tl2UQarAJyWM/R22rW4S1gNTTGaqfgoiziMZfkfaXAcv1p226Fx
Ai+OwK3mLmRrbLHr10j2ILRxDc5o+j4uUwQdsk1WrtozWq2lFt/VcsVcp8g1Y6cp25EWp1rtSlj7
2qiJR/b+aCbJ5UBzrCNIpGx9Wcm7JB2bVrrnjQQDQwhxh1Xpe46NT2puirii2n86PRVWNr27lII6
QJodje7iKpexZPIHs4kOx5FvsvToKRhFa2MS0UPhn/5iE3YGGKFfJxgf4dcCxLSott4lAgAzCSQ5
bUWkbwbBl17Erx0sCRYFGIvUtRwAAhEgyG6JsXQCTVBE16AGwebnoqlCTOz00mU0t7z/0CC9jaur
2laBFwddbCMxzFgoKV2NUIID9pkTfJZSW+A9Etj304z9jCY+0E7diLzCjxNaxLJC8fNbEKfcg4kl
mLNoLcN6QPfTMyWsoa36QkUh4GJCvCK9dQxAAPT+bWI+wQr743FSl97q58IdJG7YSEatRKZRD/Lz
ryXHkwCwhDAxzQk+YDwA1zo2ViGm3FKQ7Pmbv4sRCDPTwZlfh5grG37EtetA7/nvVdaOLk6Zvw6Y
c6DlFdnV9AHMYPHP7e4ZiTp/1FYZpCoPRjTTbMEEWCg0VgXxzqR+etkz20bWrUXD1ZXXvTSMTFgN
zxo5TkrTwoOe+Et1/rrYSgsoIdGwdPeBnHDQhVo2oQGJY6UkiXiFZPECqwGvjysf2ZBIERUNYr2N
xRbhRmxVnXvbyydkPit7yUps/eV9BZ/u1HOtj121iFgfFjmf3MaSQY/ARDQ1uMuHuULf7wiFSz5Y
/GOXkUtWd8oPCLbS74yXYrmevzeldeZGaBw+aurrHG2ZUzJqFFUzSF/PwRVpctqMa2zivNkE6DCb
ENJiHZxsl19hymBnGtl2Aa9FP8+Aq4PF4naCmdFuKWJprvq/ddZGqXPV24j74Zc89h08jqHY+ztP
hfWVYZDute63Ev7bYttKbkvm3GX9pFRPAYTm5ziulWHPz/0oJzTlzJfN6fFaHUWD1pcLfNbLMqwZ
ydJhsCGWv9kcCG4RWGwnSI9keTycpANQypbIeZLAaA3UD7S1o0eLgJyvv638WZUhiFoAqyMMT2do
SqRMbW/hnaEQQQkCOhnTjLEIgk1vfugoBRfutWy59izQWLI+0PJqR4aaaXHRhC3unuWiYF++XYL0
gcoQ9bPASg95/edZA+oxIpLFjm5BmSlJRkO1ib3Wgo80391v+bjctKrGqumTO6V0rWRZVTMHc9jN
WZUMvvn70jNHuyXrGGRl8rsiQ8o+2NGUC1qyJrZ/y+YhUF9KmO9DlS4o5cQ8TpCyOHbNvEdlLE5s
wy+2ttobv+Vv1e7NrA47a2B9sd1ZUy2FpBka+N0abpQxHY8qIJmYowwH7fKKA9CoToT9Z+MBMpcA
KPr6d4lBD3hviIYGLvJP2yddwPCh3+DLxcO9Vywf953bFmfmni0Oh/SAKUe3p+uXaDZQoligNoi3
lPiMLQ0vE1mYt+0W/sE/assL6DTG3lhe07JE5IN2CBtytpC/SF558XflD9LVRDMBssaAdif+8k4n
Y7AqWYEC4lRLlo2GPDQYVNMJUKp9h9npRAsLaJga3YntuY6XsJNfFtTJNJgHjO09WFOM9QLYA56r
pIhrbPYJOs4cNw2/lilFno8qrY1aFXLd653+o7KsAqbSA4jFBPCrgBakUUFTzpmb3GnwKdEQsn2N
kJcuw7ggGw+cIWQORc7+aX4bctai9sC6zG61PiHrla7hPiXMEVzFzLLKe9WkpbaET5IYUDsva5GD
hqnLVd1+M9EOyZQdMbTlfvYew0yfd8atslyhEyilhyPz8IGg0QL5Nbc/8a8Rk6Sj/KAQezskDxij
u42NyGWTy/stxfvAcqEM/ZIU4XHQQGR/CbQRBuL7Mb5LBcJ90KxcY0bQouEOLh3t1hMaRUDhOGJ8
sQrinhuE/nFlamz3DEs9+StEOOqeI1tsIF8k/LSX2bWl1rL4grtqXBElDq1Ob/+nlGZc3mwSNi6Q
5ldGS+M1LXrcos38sa61xi4XGag2onmsEx629x3tqjR0Su9xMmQ/wdkrfD5jSshw5SvnlYCqdmO7
99R5+ca5XeuCpU34Uq3/IDtr6f2pg6LX7agY6a9jiDZINxpR1hullV0DxshmIcWJ/8mPjZei6GM1
Ax/SJLQi5uIPPyE4wpF5fecmNN1v62EJoBlYbE1WLUrQlu7SwaJd1st2atm6Ec1P6j4ThB3pTyxl
jK/E2WkMHy4lA73jewEcBm8uXwHy5MTSJYz8vyhKfUsaRVYe6hlep3J6FkpQUCBdSi5OUNwE5FJf
EUm4eOwNkXdlpCqWsWidnNPN7Jqwk5i1oY8t2Wac2Xo3rYMrCGpPqlGOB9FUSqsdz2d5qqPKKHBt
gbN88BF5ppMvxZ4yc5tgBbnoJqIkEO3MnDRWp7F0ooZD1l91evc518SHKPfyFzw+QP5SUER5Pabk
MvDOtjUc26+IioMYCIHAp0hQNDwW50sPEKWe0vd624EHPbvnSy/NmJ++ygwaL4u8kFVX/Fz//z5Q
eKCKdSi5R9s6aErYfhsAwIiDh2hTSkmsb609jZuLR0AcJovz8vZk4c4PVTfCqo10UfCtf/pWu975
Ar55tSRHtBA8AbbxmsTrzs9lz1Lpxfn6MdTQnfrsl8WCPf0fFIGFqSSBFE/zQYyrlBoQg3cF/Pft
HFU4vaKV3IlOOaL/8LTtP01CsmO18g8kk8o2gBJdx7xPqsXYaGSjHwUPXPu0op8hlF9yVgL2kk/g
NBXe3jsBVPMRC4z/89q5QWCDiDSLZUyC5Tv5NVZgdecvQOOcQPjKh/spb0q1vvHYNaXhQZ7ytUpg
rUPi/ATXwJkDh0jzxsCJFbs+AiuKkMT1mPjswZpv+1lj+NIC5k0uLZuaQtQ4VGNx6eEGYYUZyEg6
5MAp07q9/8R0dvZOXFEXNQD20NLCDMbYlrwAYIVGSZ+x5L2l6mC+MBWCQho+nq3qjrNHgwEW/uoa
dgmgB0PCd0Q+VW9AzVXKhAqCSCGE3196Owy8EX6tK0UXE56XRCfbLi9PT40bKoykcdhUDDFp8ehz
Xdz5RqV7+my3YKIo+8c8zvG4tprrPygu4cjo2hKfApbr2NGeyWtc1QdBoT2MeXIytB4Ny2LSw/a9
epLumexykzhDQ8a1V3xMDgR1G7g0xKQdqfZ/BesY0C8BUwUZvtdh4kuyGUzrlPMhwbFWGoN8oacl
HJ9XlBgA92v7eNwd+yTV2HdBgdPTd0NStjkbhF29nC2wkw4QUcWvuE/K7t0u4n0lQfQo1DFK1/e6
EEvaM3/JAhTPDktP83K1K6w1ZnrVYMaxpdPkPryYHV7mrkmQbqN/RuBNPHULvB0MFUWwo8G8mgyA
zEQTnIlB98fHaDvgFMxxltanbnp4O0Jkbvs7k17VHdn2BGBfGBc2EqrgdCOyP5Hw7LcgE/FI+2FA
Mcaxe0Zc6rc+A6x7+479sPVxTGEeKB/7RMUAvQ3IZaUp+LgUWpGDzbc5jGWPfGSYnGDOl3fayhFc
xMHBC6N2kHxE2DwjNSMpo4wQPZOQU5hFwWt6ivJUalCGSRuK1sAGnsfnWVuBWqcXGWQbzkSAQHFE
I8iCqlgbaAkRiMva4afPfkYyxCohU22zw716tZ8P0Mbjtes78TAxa0KUD1NjRDyeEs60hWwintlZ
ifELNf+d39TZbQPLByGTj1BLjOt+qAqNdLYGy3LyiaEb2q5RaUYDDzg5kwaI3mBPi3nc4qkzY1W3
QMM5F08Q2JG3m8Q3jtOd2pS5RwRRZC+byMlgS/Q+z4gVgkmz4MtXTvSS8y4OKhOQKOHymN7akRa9
Z3onGPzqcUuZo86KDXaC5PsSazWOvYfqVYnlgQrGe38/emsPR0Qa308l3qRx3MvyGeQdP+PO5C5b
0JHaIsS6hfKyq+kZeEbGEMTqYaoqAFNaqW7Q7gqHFw62qo46kXMJeqs9BeqfetBDB38TxoehnKec
Y3V4TKiUNV88rgPN+fjUGIT6ckoJrO7olPjwbLAm7uvY2AG8Tyq2f2t2+YdhZldcI9kzn4HFCFxW
LQM803vqlVhFEa+sSkFNKYP3xyWtP86+O2xZc6++2AYkhlkvAfWI4eCw/3hgiTuRJmADujkBErfE
WI0hA9eCp2lJYh12ew9ucNz57QkZIIKwZ9vEo1H8izg8np2PdqgroNkDsVCAwSCRZW8Huvb8X1zK
dRQRI0fq5fTvi6F/9FS683wt+ia1EzACd5kDFfbQve0KXy5CsJc5lAAAqnIf8pqRvxk746ghWdas
7SEY93333g9MFFMnmcXP6W5OKAw2l6+ljQX6trgTIRMDFqe7Lw/R6ku4n115KgpK6xUscZA1v72w
L46EaqG5/ETOGnC/3CxEoAuqhfX6PcN0WOlazqu74OnQX1ZMMGi3JzWtgkxm2kFiPZQjayJjnfH2
slNdAPpF5ju7pg8tRtQl0/44uIDczbwjSynOvVM6CxTfohd9bRH7bt6xZO3jHMsRrn7IYXGGV2KR
MnV/P/rNR/VXPVqNaEjxZo1sqQkBbKL63OehtDJdGiiaIgVnJ7o5qpzqmw5n3sYW7tSxBnQT7cF5
DDaj7jPSsQmJ8D8XEEXyhATEe/ppffuy73r2Xg0/nY7lljX68KVzGz7JSolDTse2Uw/u1TPmU2sp
giBvHrWJZ3A7e0Sl0431kaOXX4s6twnLVWwMgrCi7D6iEht70/0VSfgMfuzXfwfGozIoy4tSKGrM
bGdP9IUAMjUAOySTxpmNVviyjx98uMEUgl53B1Fzv1IO+D/v3bD+tw7qV+7jWVWoWpcAV4LvHp4g
MRyH6gU9peFRw60XnRbwaV5+frUG53qGjKKQiua9dsxS2HQRLTfb2U4iCCSitnk5zJnY48itYvSg
n1E3S5HvQO8gIQOIt5BlEu767or4htYQwmWyfIrNgmQxU3bDurca9nc/F1/qWLWPIn0/cWoAprC4
R5M4vXGZnlzJICwNCYZdXBFKbPpH4PhLgj9EiKFVkQfBtdrnwi0EMrgZ23KqBChDYY90y1qnE76+
W2jd6pCPRfjtbOVUyiaWsUkx3Br2lby/q41uPS4lmZHXxbvnOmAyBLfZP47M+IxTi3A8iaeCinlk
hrapD/CMTjoGUYCQ5ktcqxA0Yf8DgN7eBb8PuzvXZwVzwVZN5j+npkjjgqz5owFV+f2dYsffCftE
jki/7TrfDyf2EYTr/pUciIZm6++XknbaewXMWc73MG68RsaLaLIH3USnqav7E23rR9g6kMDCtEON
+6jTdhfrbO809NYAREoTTCOetLAjz5OqFskkZu1ZSk085MfjZFRBKOKl8PkkKzcihrrgwaWVTtn+
fzuFPYwCTTa1DKbnZO/G5op4tEPiZ5IjIQmaauB2FqrpRM3RkhO/fP1ONjbDlOmNBWkXpx0i0zbp
tuLj/JdiMNj/quCiCfZtGpGZTcNRH6F3o9rA717hbVeuWtUNM1UfAJ8AL+q3/LTa2lm7MSpsrZoy
oeAzKfT0xDwdORf5Xhnpb/vBNeSECzcKNegRmihNp1A5lS33SMTI8j3qFDAGl4RiCM/FmXbhyErf
lrqzVVsaMNJWTFz3st4LnJ7bdj5LvCa3lBloIEeq7MenVqUUQSrNjmS4vR+FBWJMXvuNx1NylQPD
Fppd+WELzf/3sRNsB0NIw3/GMc4EyYLGkPYitqKXkRiB7zvq6RGhMvRch55RVryhFhOCFzKuvam1
3L2xisk0vver/FF4nrFN87SQOdCFBpIIpVZ623DHQa3CyOxOj5UablIqs9dKQOulnx097+1T/s09
vAdUcihJOkRMDxnEg3PiQ+YNTpHYozVfZ9DlJyR2lU43xYXQRshEWep7LbGpgtRhQ7MUvV2xwsmM
EefrWQbpv2nhj6asSuJTGwGkS1ORgEUr39t+EKc9KsM8U3Xhs8iYxqW9l3CSfounj9SedjykaEKE
7vaqhd1vKqZdtmv5OFvxeBcSQLwEgZQskype6s1MZMaOpGKvvgEu9diNCFKN1NFn2R11KZwhKGv5
oiOAAHkvFvgnYboPpNN8GYs++9keAsNBBiUEt+qiEQsU2V6NT1MadgrSSZmLHnPiofhqgnSkkePU
Q/mrMlv0CAEHQVT80oTbiRykK9AxrdC/+ntLnxuW8uLqnCruE9N720oLuWVsKWdKZQew8ucuQzpp
1GAS8gOIQtGEWi7/IRgiDEg39TYmhe9TUYt2x/BQazc0g5TvHRepFf7h2ltxtgoIHfv9+pw/U0d/
8en5jhvVZyv06Qr36vHR+zNbEca0+LoFFont69A6sk9+ghDBi3dIKnPUKDkgafh1tUH3YRQRtK6S
Eqf10jc7DZvCjbHtPuP83cIJS8K8ydts+LCpp7DF4CcV0iEZkMiPvbVUu+JTPRQwVz+3hj5tqrf9
EN0B/dW5WDVoxmD3DfVzDCr3xC5IbrIrcj2drgw+03SlL2wvBovHzm8GBTMWUVuGiA0zvViPWXyr
GcTVxpxi+uQ48sbNNXx2maLFWTRBPbaNOTB+FOjtjqLE4Xr+7K4Mwd799WYFHhNSeAFCd85WwMvU
S0No7o0WhMXybvZGc/E+F/4j5HKQ3vRupaZyRzfdijoqLHjzbDd5XZcsq3AappUsTVXGSyxhiidQ
vhgg/cifs405wyQkiac59WqYMTu62G9Yqip60EE2BOkQ3RwAd4N/PH5mdVhausO41PaCZpwz0cw/
jk0oKEO1gQ/pHJBm0n3xd8pjz4myAlOldzrM13pErXbHFiaHzfKYVbuyKSMIUnZA9UFVhxgJY2G2
CiDa1mdGtIxbLtJnezhecT2ymQ5mxSpFKai6KyxdHoPZe0Swexge6+e5/deg6tFHjMAzoIAEm0iJ
dIcdjTgAtGiLy3Av+AqQgyywEhGCwm8I5KDWQw+3FNTSS3b1JcpCyJ4jzR8rLsF7CeT8vKukRXKH
rUKCqS0nUwNgBAiBrbk6UdTGA8dsUnY6nb7Sv673rOHnqB/dUqLbYi73tLzM1ormR9286v5sQayw
9J4sjNjj3Lgf2bwPdFYIMqBbj5lVTGAyOwFG2wqiaIGPbk5ra27Qc3OZ5nL3wOHONFlBEwp/C/Ud
jEGmsz15Q2bi6VYTMS8VRxfshy4N2ASfIIYy4vm+5BL3lRM2ig3k+so2+9cGzN5pBHLK80ofiDCW
scT5pohITmKzHyzbs0f9wImcEzNxycmT4Uwn3N1b/qCQBijEvBniisCJrWzELqqeV6Kce9u+hWuG
nuTxXbZwz5mjyRkQWFosgWkeGBtTRhAXA6qUjNHI9rayKsJybj2GxJmh5rL6MWGkZ9vwXUSuYMwA
WCqqvONPlbXJg5o/iT/GL+zfyiXzfKwzGVEHOd4gX0Tg8LaX5FzuIPXHvLXiVUjfJHC6+0hdu7dJ
gdXL5PJl1FsGqqzfPxUIzoIT5cX80oy15ajWzwBzqzrn3LkOYd1ZElJH4mFR2Jvi3Uo7GVFS3Ru2
3MOhwH1gqnxQKEldH9ASQJjf0MmJUYtbBuBo7MN62o1yLaxTYIFnY4OVID/Beg47JQj4+BUGbCK/
P7cgjSezh0KtGKUSj3BuNUcBS62yXM1sy2QpJ6rD4PyN3Ri/mJc+gTWllZ7WzI4y7KAuiE6xP8Dg
bLOqPLuQ65+84ywIsZwLG35Vio1DxOMAEoQgY+XgBMZYf53INIRYqE7D2C1o4ZZFoYY117xDcTx+
8fC7RQoI0inOxtw5Ukw+xNqwahUf9GbPmM7D49lcc0tAeTYh/kLK9TSt2PBG33oDJYXYrtZIj+g8
ND3TJwGcU27XVu8jSMIvngxEIBCDTcE8gdLXDVQ7IwjI7X92K3O0GMnktynfxR/ZYBL0I28BwQae
r1ewIbldh2O6N0Xeq5nBScBwu6VOnDuKMudqOQZW/55Po+08AZIJ+WErqz/TUQ/MUMR5yEn34sc8
TouT0PB0hz+zo+sIBR/Iz1P/m2j6i8zTODTk63QIBozjKj8hh0HVoykuhc5F5JWEXmFn1OCgnpU1
skb2H3OeaUbKrhgZba9VVDF2XyMkOmejkprEDvpdtS9DWlmWxNTaB5snrAzkqnVOfk7UspH/w45E
x51YpP4evNmHHqlQIbRrvcFX8FY2BbfqCFLkv4mqPkmNbNjdzB2mh9+cQJDggOdwqTDdpQaQwJ0G
fInKV8rv1DYF+bKeIdwhXhPyUscqvmdxA5iNkXDhdwEO5w5coiDC6BT6tA24KhpgMwmWwPlyA8RB
cANmO+Xy4OX1fGoBRWGgSgXb5ZttHa3F+IGpIWJ7lak4oNdpoaAfCENTglofb7gvvZxaNKBqaQTu
RQo9Yf7vxDdExPJjxug9A52iPUiqgodlnh9DFlWOmIzq6iGy6KpSc/+TLAge5Usu1RK63HKiHhdN
2erDEUkx2K1zI0h8c83iCc0VhWW7HHyLyQPIi4Nt8LnkUKargeAWFjCkIuZ4ENHFu+Lt2hYwBvsr
RfRJYVbQbEWvgMfyQ0Cywv3oWVY1X6w9KOlsL+6n2BQxUbe49mLchC1HaJ7M8NwKa+GwOqKhJSq/
Qu21SRitO3z7Z6aAuZHKwz8Rx8/ZjaXu2nlikpkyP86FOiFPal7Ogo2pJ6MSjmO/cLgY18+jRouX
OxnUkeME7m6+Sj9kLG62+gIVUfmpgG318pXiJol7mB7ep4KsLr/tMR5iSAIxkiB6/EjYQk3tqpFv
kgFWkM4fM5zkwyffnPmyVzx56UYcdRibVCOTBboJRP0IAn5TpJ3Mg2LsGzJgdArcZV4jVpy1NN2/
JRuPtFVN9VZN6NzNxX1PKY2rWNGJN69Urmi8LmkjXHflHPFPZTBezp4Zt0W2SV3lnGuM8MJVO4jh
HpAONP/KCX7yAcs5i5b2u2Ggp7K+Tr8v0lo8fCrqhXMmeXnQCVsi6C4jX9SsK0bz+nVe9Ulbzb3y
45uQcrD47EYUeQWpLCUat9VrNSySPv90s6PBY8a0YbH4/siertSKX/eZz8Ko1RVZ17sjKRCMUzbt
73nj3XDd27ICF/lMNd1qnpodz+ixwuCsaP6dWeAFgtysm3E0iSGHwVP5a8eaMFKlPJZyl+ygRLs0
Fz0+da1IUUuPxOHu/icZynUjilNWtKeBqDYJjLd0pY0lRVpQL6q8kKXW6wg9QE/lCSKpPiVOrnLP
LMB7QWilPLszP+5f7Xcv4WxZGQo9yQ2IWJR1/e0RIbvchNS8gooOxBJ/PCznP9k8VtwihSnSlDra
UI67IxComY/2d7oLxnzyVVyatNwXNIkuhQuF6OoHAPpe6jD18lCleB+8LO2U6zMXM2XFY/yrj4S5
7awxK8Ynr0yXsXQONHEQhpqQSU4/gfV+V5otTI4TuzdZioIb0fL/hVN/J7RUrb9DVgTPUpCYdq9D
7lASZikTg2DWFcewjtS15trvKfLAkYvT0ke7alUZFkgEfh84NIF7+JmZWD4FDjgEJEiGdBn2Jdn7
5XnZV6ozW9/nOBnqqBGTNH38rIFwhEtQhxYYZ4ACJ+4l/9YSMrxPZ/UYfBfO6043PJmz98t7SqDc
ObIvzzCDPO/TVvlE7+Z35FB4hoBkFS7E3ymgJhTGcR+3SR0GT0rb1h2NmJla+B/GxEIxbSOHHkR1
9Q03KibTQnQEm2+OxOkSNsO30OnuYVg5sWbvdgn2w2FxK7jLJzQVd2psA5gGjhzav3nk3iro86uB
VNCaB0q89VItfCmwFY1dqDK0nTOBuhRmVXvoeq/RwMGeOzi5prtIbuRaTcn9wk3DOVAdBXxYV5Pe
NdlHULx1w9pgvmwo7ainKiar3S696MOmiipqspqKD+4ZT7vqf4CAa1hx2zVTYDlMMvRNuYyzLj/Z
JQpxBiCgIqWSRVl1KmLdEonp9/gTyFI5tQ8FuYJzi/Ce6FiTsv7zxhbHrXhfShwENdbcznDE5qsV
WyklICNRS7XctwaFItRVdeuwZcZuwqMCTQdGFpBO9JKIwXeyOjPNygtIikPTzgKBhMoacaH3IBiG
SuKblQg65YPrHWWgPwmm2Zwtib08VMhSg6M2kI+rl69n269f7oNDsYCR53zS10HRVVQzbqGcwGYo
c6zgfgCQRAcl771/ajrcuR0qPa25s8ENrFcEmYg6dicei4L8P/y6s1123xCxdGMKxJkB0rqT6KJJ
U+MMxhZDKg4uaoTO6RCtI31D5+Bk9hU8RzLrw9Gn9xbvt5+2p9W+PTsg2YmQgYr56qBV2UAdXsjb
RV6FCAL7/2oMUi/qor16ZM6ZvsrhCxVdVj9juN6kTG0Ac7svzBx8AzM0NQdO4yP05xtMZdvhFDay
dIxlo/aNWG0J1BSfPFz9+j3bJnatX/Q3qdRFzZVryys6HnWnKKKtmJLJlMx1I5r+jE13XMynoNwX
Yz0e01JNIF2xpiugGTwTOrtF6lBXAtl3wNtk0GjGB5tLUvtM3M2qnhceejQ7pAieQqT5VsuJCc+K
iWqhBNk+WBojapZlfetAuRwsVUXbQZlIN13QFuyblKsAaQbmskZn4eIRxlpdVPwxQ49wUJbes++o
tzons3TElqyo/ouIPYyYCXGDp42yvvEO+E1UTyqPYTbhJu1BODPpnfcHofNZ4l1L3x5+ez4n6s06
qoqz2ZyhuUVasQmSbV6yJULsMEJuchcBHpTqNjg8oMQvAitCO+76ymDvK6fbcWNKT8uczVEL8oUa
XTTkWiym21tlZxX5/sB7CDfR3ooueZM13TBvOSKyz+4jZo3yXAydT5/5VTy3UeeTnISS9AnAg3gX
ySax2kPUFl5povN/maQzgaPwSwLaOMQuQ5bwzYyRxTf3WQuiv4LUB64ze8r8XQ8pZS27ggCcX870
qcHW60vNhc3/CLaijH/PNZzliHmGrrd5Zo8BhT4yYeO3QMqFBC5xgXarI6EDgl4meSGYliT8w9BA
0d+uDPU8o1LCmdhO2Gdbe2aYvLWkOO5SqiyMMrl7lEDL66rVG+Nv6mm2oFHlPQc/zUcyOBk5KISH
OSTpk0CqP2lhbzuPf7qpSpPjri1TD2T8JkrOtWqlB6KH8cGLxY+U7aLOMtfJfb+Fvrq5Nif5wlfQ
GZyiZGpryARysKksaXsj/44kvtDr/vhjWLVBsQ3YHSn9qCve8wp7/VrUgIzwngXXN9NDrGH88/Jb
2BmqNtgdra4DG5qYfN1yuLIY0mDGWkIterRhMoRi98swSYrFrxJRxd2WkofiehrkNzxR7Voog7Rq
08cXfq6+iBhaohhHnjdMIOn8N+Jc5LS3jQkV8vwHrg5gozCQus6d27xZofwF1CxOp6CxzRl94bUk
DuzYnIDTp/rmVNK+nsHP76tPtLhZ0fGywoguxwzmEel87UTUhegev/zxQrQOuXM9AICnpZVpwIDm
KIkXbeBQxqjKJvrAWTibxW6IFC6OzudJSHewYG+wQu7GbKuANR/VIo60HEUa4UghN0nl4axhLRno
qclwAKzftVTnWBQFDjfy/ygI/KP1rUZXQXPK0bWbeECZ1MkYEqYtDAS4ys+U/J56mdbeujpef6gQ
GfgwJgr8Zo5oEkVp/+uFrnEnunGZdiwa20K7LJY/B7xxWdSEda/cthqne7x6waWybifvCoZC1M2l
nPU2sDsBydusa+2CJzcFjcDwb9/QDGDOyRw7hWGE8c0exX31wtxhcy0e+t/HfKcHnenoQ2voorbJ
yYJChH0URD6P2pHybHEMOxrKM04nAQrgqbYqy3bfSSQ+1h489b92g8pKrLY5q0EYUXgJQld7vgtU
rjJy2dCtLx+3e9RTsY9R3ee5AJM8iNsSwFS1wIQCnVsE/OnjSXfeF9lxMUqmfVFDpcAoIEsg5Inq
Vnmx+tupZzwhB5IoSdRYiUv/ATlXnatjgdXZsmYT92WsxPDE38eI5vWUWrLOWL1BQ2ibjYBu9SyF
a9a2rJtnhVSpgwGW33nooevbi6sS58ChDm+3erCTIjtdjFMNT5GOcwsUpWG72kBz77GQ44+FlDqY
+fVJUSdR/9EOkdHrEqMBybKuxoi/6Xkt1OHkE/r8fAMBakypqwB0CnheZFIAawmMmpR0uiFXXctA
xowbU41maZEzLDpfoCDqrM3kuQD6/7MTTKrsTNoM0YNShK/81NlGMX72bpJsic+feeY5D/MD8kEZ
zgR12/1EnwFGvvfkwHtfWyaHu8+WNVUV++5/a1LTeoTnDR2HrelGY1iPAq7LhYkxL9PqEBnVK9f9
3yiUIosuU9GnQPa/QY/KR0WeTN9bhlVRF1YWPhiRfhA1HnR6pdQkxKrOzPhWdoT8CGGNMbs0wL/2
7DwRTnHdHd6NCzyWMtMCNoe63vZHN/fzBzgTzrvMQP15lfG6vyY0ZJNPhKILLCtf9bHbmLW0uISS
rBK6BqpQaw9Bg5rZsLJwYrMotRVfuXH+xnkXXbIJPfqTvJsPwBG4qoCHtXBmT+rCfPXhQNjs2qbM
X+DNZXH8rfTdKeYeso8q/bcqz/pCtB/AQfe3VhLF5DYFkvn/4k7hl9EKBAczFCcUkXUhmhAbItAp
Yj6/4iHWlL3C+0TVCum9ibYgUHxiYx1itUjISxtFrQCtRUAUV+U99N5KQ24B30TXwD4kkIdlSZ5e
cfVjmFLZOWYUx8iarreXdbYlmMSCi5GB8li86aI7al5WQGpMFkmvDnUxCgmCZjTpYvo5NaeDEddi
+TYtkTA9VSRnr5DvZb9eTmzcO1w7gIsrhUQ/pNgHhfCJbw7DjPNxFEn+nmVURDrXfeKy4u3ORmnH
BzBA1ZP+rhsLhgV4z6YNVx3+2Kd55PIOjRZzE9YFG0VIC1NgNfkpQZW0XQrYqMr2UR6+HmdWMOkq
GKis3gyXknyj9WNYcPInoxGtwrUnLatd/042VEmlKRNlV6SHE2iW+G021kADBgMY+YqjZkZBmrtv
O8MXbGdnsm427JlhVNGplkVsgh5UOJsqovWCJhrCV00wYCJDHaayCXrnTiJhjV4/abTl9pgl7cCc
0mmn2lGMjw1SzdKU5dve7VpXChkrFzQ1R7BimurDmRjJSa7fouoTmXySlyKd9DZ0u3mEatULcA2y
tMQMng1E7EHWrF/8E2D4LzJpF87q/CCwkgY+Z+w/nnob6s5Iu7K5BQrOPGWqdVgnjN7dBGYVttjE
AN7imusqYQ5x8vDtNaqwxrQ0S5QHJ8ePyVa1JGo2g+SXJKSxNeuR7ghhGOuO1OXuVUB+kgpFaiPq
+BnBSuK636/0oDi35mVpGVBmAGWJIjM/KMqwQ39g5LkMnI8lASV8bJWOaT7r/FONUSRa2EXSy6hN
wWWiZ+8nygofdfa2ZCYoClHc8qY2ehaOjTepmHlvvdAbg75yTnbQeo20yRlbQGDP43qNGH63SOPm
tFuqUS6ocPjC/cK2cdqZklkpym8RduaVLP3bHm0ieUiO/jkrmxfjFJs+eZRmvXU5U4zhc1mLI/6o
+QluprNmpxyFR8XNwBo1/S+i8dNyMFsIaAAc+AnU2bIEuRtAc69xHwSuQYshSyw2iMKMe6q00IYI
Oka7dkT6n0lmQ3qvSwBHRRxynCZd+JAMzJJOa3gcV3++EA+xNmQtiYSLQ2+nrTBBxnJBbqLFm6wv
Hf7VZgke1Cb3Lp12cNkK3yUd3TcKe3W5/9Xq+SrygKkv1djyGJAXqW/6OpOrPPH3HigDookFWjh/
8K8i8Bg36cidB70T+csflfkB+53QeheZfNv9O5rgFvQr2zqFli1heXlQ37zn/4V1eTZosrv7mZi/
jP2akfoY0EQXKl4H9OodYQvd/GUIAAlFJJdJDD4oAHcuH1zbo8XXCXGAjsos6GAz3V8DfwqMrICo
/hHXTJ5TLrDMPHrss2eoLTumNe/p6MtyYdILCrmcHdZAodBlpos4Ydo2ON4WqgW/4e4OtK0Lgsaj
zLBc4I91Ddfw/IV+SEM0HkOyL1p369xQoaIkwRG+ryHDmLoq38fxR3FBnA4FsP05Uc8fYemU8xKZ
dlTkv9ZVAyX7asKDaNJz55nc6M0UiX11nvWzcfuHxNul+q8avJ1zdQrzJBXP0ts4K6k9qCC7zomO
U5VrPDvnPCpMxv+NAxTrXEXsZZXB4kuaKFsAx42GookrGw2QasB5hr4EaTW9O4Fd3Bem6Smoqz6M
zrRiPZtpXLrTFcPccUy9TEXPkGZ8Sayk3ULilQQzNXE8hsDiXRmqmw/pjTN4NoLmseQEWYBU2UNr
q1YP6qHuECVqHZEfSH21xKmbpSEsdVZV1M8LDc1P06hXb4jGUxmJBwunC5jPZwMKw5jyC3WkAv2v
dGZweXQnz0V0Ow1K0SUmNvtKnuzRIdi+EmW0Oxj6gCwNPSdp2lGlg4HU8K5PWXk43/Fm5Gj79FKR
BSMMVsefSDzp1jTRISmKQZ1J5TCY2GBOKfF/K6z9XPurhJOyOiMUca/8F62axuOC7LUPibzat/BR
6ZH2DjjK1+Y9YetlgCNq1U7u3G4cKcDVGIaqlBc2lwPBL7eU2jxTgb1WSBIYpWi3x+JwSkUjunSY
5FWpJcPfPJMkLLSbBdS1LHi8LBGif1Pc03w9zTdf6jD4TKuByMym4dGh4hSDqMt/dwN4NLNdxVU1
1wBghFyM32JHsaJWor8o2XNuAy9L/gGmGfPqJiNPLZB59Ygoqbj8fXL2bV0dgiuOpKrOE8YYEro4
U4EL5JpJyvss2mlfFzEfMM/Ckhr3/+eZJKvxrmalsc87kTyZHKTZxuzXX2EzSZh3Yj949KDQsSdz
cltfekNqNv2RipwmlMtcJldfi7WBOisUWcITO7Y7/JX/I0b29dqfkCph7sLBvFtktr6UY/1JyKg8
34se
`pragma protect end_protected
