// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gOK0BFV9PDt+z/xk3ftfoobYY5p9XFyNhCL2pqIxktFN8JazrPCZqqVqGaNpiy+G
i6cNIOwOgpXHPbkx8+NgSSanrJdxma/yAhTxxx/LKAz/VXNVhWO1FdhxVNOd+Xws
k3Oy30bdGL51Usl+0BOW1sfkSX/02yRiYDDVUllL7WA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7184)
X3n6d8RNoeOkBF+9ah4Zq8r5RvA1Qc3TIfA/vzb/BGIoNPcWs4zBYuzCOcn886G/
vZLZCQ56GGiLuHLO4BO7X+UGBeZZRHWeZNgLUIE6oo6YUAbQ3bO8f9Pdd7VlrIAh
j52PriczeoeBu7AqMuEPD1ftBqAGHqOKg80FzCorMQi2sfmvEzF+XC47ZaAtjKCl
/fUkUZDCLCpmwkx61gdUJ2Bc5qit5OwLpA/LQLEUtB/4x3k7PB3et6apTbTGi8Ui
LLPm6GZoE2q0J5MCZj0tvDrUyubL4cq9NwYMd3qn3uEAvHq3QNA2WCxxYALmhsF+
9wuttOd/rix3XhEs71Tq61VlkwOWeSKdBUpSrH81pB5N7A2XMqgoBOYPd3dMpaU6
5Y6y9u7Fa3G6zBQUWiaRMjZOm4uvkiKCzsHpxnKhJ66a35aGyW/WrbfudJmVeyIr
aAOeXhNVxZKS82hfflMNQ00K7656BelQw2UGfqDG9cX0fL7EC68SlBWeH0Rwfuhk
mp8rViJApeq5E73vwetaCT/C6DeKVcDA6/0ba8xZ5A5Il9ecAwa8mz0r3shf/umr
GTPuyJ5NfQf39K1y9u8uMQIsP0MHTAB4nT55LY26olnbloSygNVLw0PL27BnOPtl
fbVRRcrVxK6l7jLPg7neyXk5H4/pJTaX9agyVSOpTs+NHn2jasbF2kQKMbHawUd1
WkdRs/0Jw2JFdH/TeqsahytMeGDpiALi34+u5CySQrnUOcFermOZSIE72zxBddxR
aGz2JWe1IKN8frGZlAMrLm8eKfNnwEnsqj7E5eU/6+hkEuSH9Mc+URWJVTO7gbwY
nvxz+XXWmYDLh5+3GCj7AolIX0isDwtu8IqUI7+Yl04Lb6FSlOknAvZvY1LG7uUW
248h+o0DwfkJ+5XVaTEnc8diL2prasgJvdsidfdTJelhqYY1YsRg8UZvNz+yWlnb
WuaR31fuOzaCy4gcI9xv9R/3rvcMue42pPYHYUVPSWY2lhNf+6vQL9SNDbqn9qfP
hsl93R9vwvWTA14ajj/ibgvBSPct6tpIZBB/RAqjeZk6M2/HZgv44hokfYcHBX2X
vlk8kulJurbZjCu3vUyP19w4rVc8mLZmVGTUMEIMBVOnTfr10dQE8UEUJqZSKM2x
GdVnznqTNkGl3QBdbllOcTqdWvih2QxCtdxMheKiDsCWPPjzxbQ8w/00xhxzW4o2
f/VV12ZJrrw/T3Z7L6jxx5pablZOfGZu1JDlcPpDKDVdkWv5yYl/H+rbHCAwfYF0
z83SJkTny5zyzc+N1fFhZEyefPn8yhM5hlVyb47QHwUjk+QvPow7twHupmQiQay3
5zdgRX5zp38lnPxJ7p5rXlwxLT3bJ0BFm40xyltMg7k8U//WZTgXY4nrMLSnT3FL
bywBcQPBP4m6gIUoXyue9oDPJXVBWAXTYjfDVk8+tr1ea5DYY7O1bwXAv6Rt+PRy
0AUDnhUUm0cW9Ya9Qn8vC6twXD0dGaSCIIOFzCzKCv4xuUKgt3/S8+c8U7ZZvmqL
cY0xf6au85viAX7q6hEcafE3IYrMJsXVmEgmCnuhctsdglZB6vVwS3oQzBWRWvHj
fRWmQ4Ur4Lq+nVEZ+mQLUg9t6hN4EvKKztl167JQNoWkaGabB529ti3b98woQmJs
vqB8JLp1WXg+E18Oopr6wOmkylc3bd77nsE6UHj6Egvq/dDY1eH2hw96odU6OkJn
VmApwstGyK7u1ZMyz+C7L3WuA4OtKBltM9VsJMhbW+RYv3K3Sk5YYEkaH6MkJtPA
wyJQxH71wdgYdJtslJ8ryc32hX0x55SFj11vSbA9vHsluH75iYWHkaSXycy5/3Ru
34yub7inMXkC37+wII1mBSZclrN+bc8wbv+XLm4uYUQP+wVEXa+0dKRdjuHst/2g
g2r3BnxOeKE54HtzJP6R065BlXfZujUmc8g60GI7Tjer43E9oYZATB2NFZwBL1lj
5DOOSK06IHYwpP7VpZbJW+n8/aZ4Bv9Vo4j1i6l9uef3V8AfNoZQhERpwtMxYS1p
Kzo4Tfrtu2H47YZjt5+fZ2dsL9NZR3iY/VaF56gpGSGlQ1M+1gmmj4WK8V15qFQB
bxL6MMJdxwDlfIDSlrQKGgYxD++WMQ89KNVquT4zhOI37yz83n5jeG5eStIUpD8z
2jETSyUEesXYavcNjIXyEonGxty2qEUvhhFHjHlwGTQ64Uj9S8/IVHS0/FN0GoWN
HJ0P0K2CaAvYOoX8hLBRs+ekgTZL6wCtdIcl/7oEKxnqp7meWwqnpAAjJHGl2/3p
8jTxCHs1Tp7sATFi/OdeqHhazgbkIsVDyqYHm8r8oN2TNi5n3Zc14ABGkdHFoD7K
WJ6sBMFMUWG4RWqbvkck/7pf7SlYzlZFjjPK4xWM0nCHZv9rZTmiD3GlboydEnrS
7KkA0CGsbjXqLuW2lPXpq4msla4yBMVhGIRoMRox8rDCV6GHVLq1p0/QbGlanVne
nf9p/OPk7YrIlEfs847gyIciSQMzdRwxxoCNwmGxzKt/qkErT2VFUFcM1oaXJvUo
+XnUjmp0e/ksKJS3n9ipNe8dUZFFWTbaZ1H56Z1K77X04pt6iPmSL7eAga5jG5CO
N/iEgW28/z4G/iODj3Kb7m2ZLb3xRBVAd2wxgt++ch1OCVnZ5VWgs3mC2FG1FXT1
gc+kWMkiNFk35C3DaH7mcO70KlED6w5m3VRV8gx+O54EAQzEfjFzfT0e1JDy1wF5
Z5gOWbRak7vWYrVB4BqeGuGFEVRsjeT0fmG1vXfyf7kClk6VXT/Acs4/V7Kw34Zd
/T34P7Ev5wvRCA+RiF3T9nmE54tiwAfMZsHpqke1LWNCuQShQCholmKVz9OXEFsT
7XnhB+E7zOqZ2I8yZ/422yGZbYPhI0xucMB8AyErwENdMVXKIJYjDKOZJWd03kBC
E2B9sDdDaa4EPimic05dC6klqPomWtST2EjN57Y3JVuAJheQ/SyEEDspU12OvYkE
Ky+XF9PL7WSsD0Sz1W2a3SCY9XCb1JXEbzX74XhbXHTserroSHd1eNX8yDYxG3WA
wVgCr95rGUWElQNukWqygElq8sZObNJPEd7+qnm+9ANBlWm2p7jfCTiAL2YUeDGh
8VcWbxAZ314hjDa0ssHP+bjK5lNyQiWSx2R6sbxJP1ybDlL+u9zWA3st68L7WTJY
mAUVQXR4oSVBzlZynsaxwfEtLDkkRTUbal9wh3RRIRx+FJsy9bm0hAvy5Had3krH
usC9nxJptQG6NuOC+z7MS3oKIMTDk8DvQzupuB6dtEyXbdXRyeJ/1yLCqe06LX8I
GuJkvugU+22wLciqzDhRdTDerrWbTie7nkIEtu1bBP2BWhQNc+2y4xwEzCCwv15T
Ai/eF5QkVaAolWLq42XORpJ9qfd1zL5hFnGRGNpFo2sCrEDFTT1u33UDzPiqXo+H
lo6ar5qp7r3/b/EOXY+8FvQd9qb3cgXFexmxNIg1WnvNaG3bbtILBykyQHyGIBNF
Oig4BawHtLigCuynTqNAofr8QkToZZRpoYKu1zi/zNCj5el2vXhRtYS1zHfDn+lM
mNtbL7EQu+IZyDik7gin61rn0atXZq5lxrJP0iqyFyMj/1DQfGch1p6dW6+AOwVN
2lzebyho2UnpUtqaHxmAtVsJuuJ+859W1G939qWndrJW7kyhggFbt8+3zPFU8WZK
Xr4ZdYzyHB8Wq2H5wQYWxaoaZ+OcWQk3xLJwAeAJemrhYcyM1M/6l8K/pJE9RSBa
RLjrKobhYduZKlpEIDInh8bN45GrH70J+UxOh2CkzoS1p+648+fl25hBTR//Q3TW
BSQNPlcdkjelofWpQvJYByXhc+mjAl7SEg40XOYZ6cuSkfG8YDO+/tIn207Toh57
wIHOxGvrWwnzReEZoCXUYGXCNCZyNl9KbuIBMtCzxXZDl22WZmj2R5Z0Mk8eYMbQ
SIHAoeUxIyqNObpJDRrP6eVvqe7iKcisRgH8HrXqTS+5HBb/FemRsNTdQdijnA9F
IJPvwClh9xGPD2n7+MCPr94n73pyVcUkN9syYzttS7/a1QTXXUqePY+vZY0ROPsV
5FG4duQTwjJqDvjGFdd+TOwY9kBTMjUO80qYc1g2kA0ufrMuga9RF10aPetnl6/P
OUBlzmiW+eUFeG+ByDbZHH+V7uQavwL/quL7i5a7dCTgSd2FhNrzXEtS0bOK/TTX
AvLWcFd+qClzLFcc/h+nAVuoa31E6e++OAyo2PNjnbb2SpyTr5oI02R3IQcmvoCc
9xGrP4sGrJVeaeqCILCVXT0rgCOg7lFwdEEFnIg88KJNeq3ZWY3XYH86lsLoLSbD
179UCH3BxVQ4FgZVheePEGGUlTginZPaMF7REMccEM5VMf6CfmRK6uxXSfHVw537
nJyFWUj1sZxzO60FQ/poi7OXDgsdCuvD/Zcw6x1Hx0GlDMiKywGNyYh9zqxYONxp
KPKdyHj6On09AfD05PsZube6x9G8NTXCcW7HJGYCovpZtCKpNxhB7+sx4csuq7NV
1qG0bj8L/Si8KKiaqn7/EvalX1WO/LqOaMo3NHDygjlMgOB3pv+PoEmXFVXs+wtG
i8qZc/NwzsD2vilF8gKZAoqXGgebkx1koQmJ2zF4AMTJ3j/dcItBvO4WEZkmENse
bKDgmbuqCuYvQLqFzAw7GRBMVdedQ0fR3EkPgRjpkd+Dm/lDeK8fNHBJ/AF/uS6L
zjpJRZV/Rwd6yANBfOqVlRYt695gbr4Ao24wcxyChwW1GRQ2N/5xlmsZFkg7uCO4
H9uGu8gwwTV8H5aXEZIgrTaTQrXijbxDSM0DKg2GNd8xpGC0z0jvxgSgBQX5t/6b
AVauu0WCXXWuQfRC2q/iHaI5tTR9p1RGOOp1WKAIbWmFmqrjlNh6elY7uAuFrN2E
LfucmFKmV+B3b4YbGy89K6iAHVLaA9ylsl3xex5VuRKVqUtjoJ5QHakL3lO51sy2
Nee/ePxR2YcI9hieMRigrCPT1VwSb4z8vaQzBXCIoUQ0f5a099r07x5zLuyK314y
kT1ZNK4lG86cEilp7SKmnJJZEZxuyyAa8rcwDKmfwoT3FJu++NY0FIlYW4fSv/Dh
BYLaiKGzpaurr6z6GkGH2PgZFk4qZEdUJhZ0PFUn5I5yO3QpwJVsYT9UxO9mRC4a
Q0Ke1MuQVY2kVKZwPSY9K6NHKZeErbtCUI40vG4JPAiCU1pTvhnuf+GAjmn2+Wvl
afwG1yy+CvTzL6qv2rhsF7xAqW4zZlAhiouXOiY0xD7HZ2O6kJBbN7WPVChNzbUq
EAkQwnLpMdcE9NMh6g+5rxQDVMrleF37NzPl6VpxesujTnTbFWib0uv7VDiXAv/g
mbR7UO2eCN9XqOVPPgF+kgYuhhu0uANGXrtBNpBS0mZJ4wis+oi3lmRisEpq+HDz
sXvlq0MAC8Jqt0xLhHTpUj7VG7zYoOZmXBz7tzpHbnbWKfNQ0moWoU72IxUBUyGY
2zq/d1IKZdidXsOs7vO1JRC48BuvsvvcIpl3z8dWJ6cDB0nOxF53QZOjOvb+XHgF
R51Yk1ZYezuAHCpWN6oSHhof0ffZi0uC8PFoqoUJ7Saf+xPSVUIMBn21BfGcS5pj
tAFjfRq5DMBBqFhhgGOVrfLdob6XqpLzFlj0efyB8HSt288Nu40mK1kFMv7ifRa4
7GpVvWFxmp0G4c5qdFF/7Apxl9/+3qWgidC4OHos0uZfLlclF/HSj7JTvAMdF6sA
+aOgc02scgRIasAvSxozuImaN9f000gw0mN6ih3n6gBOQMpqf6raNHGvjONWCYlt
jeh5bKftWFAF5moxK8gOmMCnfg0fu8PYq+YFYCV/JbF7NbCGDQpvPkAtHAbHq9dh
ZDg3/FTSP5SfEMBKTkZ0qv6Y7cP1y1/VdJfGmw0WXup/Y7tNsP7SWo5Vp2Md9AM+
PKwN/t8XHnY0SolIEL+vHuF0p6CQxQur9O0iURyFB8BAGsluxi37YGv37JtMM2YT
/fQUnoOCUrRCYtqXuxM3ttGlJp6ZWanV2mFMxl3inK9n3xqRGTTN8dKWhLUkacJi
q/2xKdcGfrWsCasUmEutmmvoCagcEdinFQmzoCvroVcP7cNpsV8YJMud/z2mPiB9
EvFfb03pCKlwqqjFzmQD7utij0xCtY+8/86wy3QUyzIC3P0mYFBFusdUCeAiY+dG
qkqXraqYwQ2esSHsvJKwV6l7lZQMgb/W4vNGRRMVQE/Ule2j8pITTjebwjjJrR2D
m3V+0bsSZf1LzE9lUXAEx5kZoiSPwxh8pWK51lgeHKTVK7jIbp3JVvJbO2S9wecb
qSi8eYn2xaWTIzK6F3wTiB/7/ivhARqvzSgsYugSLGcGngH0per7soQRevMYlb4P
GGhqJdpB5ujfVkzYk2s9F6ehcvuOsMeVUD2TGx+DM9ulIDpDo8CLLJ6SIlauvksV
/m7A4Sacg2dZJH80SGPaWTwFnUCdsCUiZr4T5qB6JvjJNYAWLANAdXIOpduGtci4
cAOzp+SrkAHRmRmcya36LfBr1FY9LqDSE1O5Ac9IHRPZDSBfqndJNLddWApaOsNa
rdTxPNCZqMNCz4YdH1bRN/bTqqO7560YRNtv61Z71Bttl80Ulx4cZXDBO23qDd/k
4XKFBDdnHnLYUq8BnkmId8PvEVyeDO4HuK5fU2FIQFdmRIdc2DqBHLHFldkSKx3x
P75sXvRWIwhM1bQn0yk7zzxikO6LTJGgQCopwxKA5RhFwF8gDzCuUzjikgB5+YP5
Un9RygAIL2N3WifQIloeJTCRLbM8sg8tzIG+RDeYJ4olvZ5DmY9H/9T6qYxY6yQ+
ZYE6U97OV21FDB/95Cox/NuV0QqMUoeVuaTXS8CnDPbym96+eeMEhYIxGqTQCzVG
CxKUz25vStBykADfKuggNCPLnVl+TaJNaQEhEa8aQ51oOchLDE2mJWGCqoXeoRVj
ITxesMdFQ2jXSk3CIHjE/wR4fGuSRyxZGhr50i5619/W1Z22T2r5osgvrU+ziC4G
m7j1gGg+xzWPQsutmXkorExDtMSkvKBwonaYS047MrapvMpjKZYqpZvMg/qFH+z/
geBlHod33lNGJOnT5ssAZbqdxz6tk9LNNMs3mWNFpMHIY54sn8ioCo+NNdh4WnIx
zfMupSQzH94fy0GspOmltVqL3NnbbLC1273phQYGmqnVW5V67KcEs+qUjT28naip
13eW7xW8QtqWIbLIwzHo6sdNszDGroNrK2DB6roN48dosLSQcqIHSzwokE72WXr6
YtR9oIpdZuX7br/o3HT0ArcE8yJm3/HPBCrqOpdQHjoyAY1wdilJf+8ns/Wk/TGq
LkycD58jtHPFwvF/OaxyGDGWX7BITfAVnZgVywJBhfH8mm5v4t7rjgJpqo/FOxvm
STwr+o5ptTf0tC452JWiLyicsZh3WkVJmZS3zv03KuPkQ+/2wUP5Wcty9yJT5wer
H1HyEkuuRdTIbvbH/8KuQSdiFyrbiQCx+XfVS5Ppe9sy/qJ+f3ReA47+nznNYmNu
Jgncg9pMxs6ROaAmdM5x+pSucFhtEt0pDgmIxun/6lmH35LIQAqE9/jgTdh9Y3dM
u066/izOwWUoSI2oQ7ylwgQ7eyurZAOyTpm7bCuDjL9FtqRli0FNMrlBl9AjFPj8
f2Ghhv2NPNXKEQyMZIMd9FveJk1sc/pXSi050dONWXwqrgyANUkr+JqUS6Eg/n1h
IjY9/NCQ+1g7kPsCU4MEDY+CgSMGmcwt0CTa+rd1suWLGpPai+fiRL1sHW0+OrxZ
rNFdPM230FBDOB8d729dip2tR5eyc5ANu35wE9liUjTW3QjueIVy0hhudxI6mgg9
o2Uc3ZG3jP2RLCTvT4Lr41nSXd8K5n/nLU80WZQQE+O1iLFHOtowbAmmIHmB8A1J
s9+LRYOk5rgPWiN6Cj2tuA57HWs9eZtlJ32L5FQcJaBpqcSZqD4+RaGpNuDdkiO6
Q7LEcLisJnrXE7BYJl/rPnXAhDTmnJ4eqhjCJ/EL4DFskdZ48VMEljl2VQN2bGiQ
KJoOAiwQ0N0CUc8wU5zyDU8B6aqhpR9bMzoFomXZRuhzhd+QNPUcbQxeX4KtL+2R
PHXGllQpBd0CwIHbau5h0OQxvInCavkspEFuQZQOpKU2c3hwCmpes+DFdKxwc95g
lHPgCyh+oMaySkCl5B1Kop54grRgMz953Drbtb6VRaE9Wq+abmzN2co4hH79erPh
VVwhWIhQ8qje+vJN2FaO8zyPTbFUvliOeExTkWGd3V1o+ebxzJP4RQCB3Mr+egic
avEg39+DOucxEna6D4jTdI3db4fsr01ttWAi84yPQ1/cTL/4HEaUy7/ywo8HSNdU
mKH/XGBji+CMoUbr01F2/zw3Ise6I6hx8Tdv4ydbtcAyoaMqEegUuI3ZHbDpxPr6
lZ8SyLF33p7IDMiNWHYp5mfq2p5u+CQlUUGntu0xEoN6fR82Z1Dmp/uC8tNLl75x
p8bPC60iYV3b+vmATMp5RI83+lrbLOUkoLT4cqmkIhuUtVTXiyFT/rpbDEHunoPe
uE/lwW3m03HTj/qaJt/P7XBUusCfrkCKXkrUwm/G0iUCNCF9Z/ZKK/Zwy1OTSY/7
1/LDkwGaAcGOBvZHW/Fu6PShSYIYQCRHKlppLvziL1OEnYpgILzOw7XP4Q/KbQAM
DTohST4Jvp3MxXCPRsMrdkN5TO5WSTS6HVd2fdiVb7sclc23h2xHXwaIqTXzBoiE
ld0QecXPpCwordRxh1QbCqGNZfDPjqarEMSFtzu8UsTtayw9RP+6eyBl6m0X5dR+
joddpJbo8eMNR/W/VDZB1KM/xrvW0lqfH3NXVyX7ceQ443GOd6yyliOCP3igSPhN
2CjY+Oz3Gf0Catmp4733Zu6Nm4oG11zuT/JTmtiwLBjRgFiDBf/o67+CPVbzS+II
6GXPcQYz4T1fShNcruGifl84YXkw24je75pJ1F38Ya9cj087Tldkjetkd+6/rkaF
NIJ52ET02giW7G/CxgAT9DVHnribzDGsbaP2w22CO1o3W1ZWU3kjhl5++bD9xi60
nwAa8IOkXZ4/rYQXvRR3rymcf5ye4eNV8f23AjxNIvYMna6bMruRPt+2Q2DnYa8q
enuCjO2ZpdpwMzIlsvxBONjdvEzL6FmsDdu8pMUvvNlFJ3vl8sxMI/MipzfIKu3v
0ertyL7TzsvIL2e5d18JvRwPzs2tXeF7v9cBNkZ5LYmKwStiLF+fDheMw9lFfb/g
yF95zX8Xuw9EIJFWg9B2fQCBPYJzGozhYw9iQoFi3OnS3Pj37h5MFv7e5m0OsAFN
NrFDpdiaPjuFD7G/p/O/HsjPbervpEN6hzp6u2CoMtyQfFX11L7EkENHDc/aOAh+
KWSMg+rNRKlc4pt+V+2K2MAiJTyAwNUuvegvhtodapCF2AcIYpevq6amfbiZAMCz
T3rRWqn96MI/hj4R4bitDYM17685hIgV8M3BIft/y1TJG+USmaq2JH/Bke4mXvED
zJKYz4LIY5pH1ZcI10DM3CqC8uEy87cJRru0pJvvn3s=
`pragma protect end_protected
