// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GDR/py8ZYawqC28jOzgQ/LZBhNdXKOaHwx/w+Fjy2OKEd21lkjq+wX8DwuTm0K0K
2LwmN3liLXh9WxZK076dZNia/rVeYwcy0UtUli4FSOB0YtL2kug91lQeHIz/B8fW
hRmthYQ5MjaPutfVeQOqNgQs5gFw+HzrAHU1aeBDGug=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10272)
3AiFmgYpwoulMoPMnYq6fMMBliQniQmZ/WSYTLch8xcj1QVUGxhMrKG9YqTGgNX4
SHAvgG4TIJdarARkcyy2HYC4XzEz/2mxxnCQe8AS0jevdjLLiYF1iAuAetqrs+iS
LQQfFF6Qx3YB+JJdRlR3r3dkNPk7TAvNyupIkU+hMQg5q+x+YQrtR2XM9XX1qRXI
vwkpdfb8RU1ZYs3zQjCR10qReQO6+mttZ00ULAT2u7ZSkAIj9pxs8S9Qmax6DWIe
X6azTaU141kRUcb0KRKZqzRkEhIjVVUe+UvPHm5meq0hOBNBeOlTMseYN4C1QKCX
2rRifa5CBLSobEnUmDbPfjri8HLW6ohIZFcKs5ECKuH3OQOgUSJDje/v3t2hzExt
6mCbXguRrmjVixU1sxQ9ZfjPPOFQsRLkW/TYFjbZ9ANiZ73r1woU8k8XIHt9/GF4
yHhPEUVYreZgH7PbklXaHfubMABlhKP0mqAHJxMFH7ZQCJY8lSzpwEHdGzOKmdrt
lO9iR2o1/xqa5/bS6RodSp4D+QB6vsuTOqnbsIo9rQbHnspqdm1MujFQvgQz3Uob
j3+l3GtvNte8oWi8lmZfUZwaSDp+rDBMo1b0oQFbcT6IFdgjtdztNa47YCorRFwG
U8fbAID0L8zgc72tDlfdX7EtxgoPmuVo35fg0J2lyQV2xiFH6Yn/rnk02qBRs+V6
fEWs5nMRAjCXe9IBweO9jwIyDrf30DVtBTsu/DkQREFMVLGUp7WqpI4eNV69w3IZ
4R9lIFVeqjWCg0NduLWgCfWp1tyjfHd5zDdfmklcH4lmaJLw7q8njjtE/+sSd0Yn
JNGdm5L4EV9Y/s42kPhq5p+q8tZ7UVWmnSpIlKGtdeOvVtehx1+8ud2H9atPiSYB
WJv1R3710wgLRxlDuCbXOCqmaW+4lmCoWcVxHEtJDMme3oUAtcQ9tPSgqu3xzSDN
ruCKBHh3esTGTDxgFT4/PT0X3NiCSzniHjF0S2mUnoNAuUXuHq0gS7LktrIww9kt
OZ4g4B73VIrmLH2dRcWqX5Jbl2Mhyy+Pf8krAFPanfwU8b9kn306KAQFM2dLdimm
6mw/p04D2V42ivQ2y5FW/qMUi4qlt1EeSy2eJ6tij+PRvQFHvewcZxx+LQGLh040
tfmAKMnfIk97ynEQ236QiuXdgbZVy6pl1ELA4uO42jsOpgBkovG7sNPdMuNJ/5js
yEP2eccYa2pYrMF3BjzKz/lGhvs4EtREA6B1ePLiCCtq4fRx8paZabRHKJmhDmqs
A3RUoai7Ja/KIOfUxu/JrqjUlF7RBfVUsOhvYVazsjv2Mn3kvBV43IBpD3ggwT8d
NreK+SaAK/8+DETBbaLN/KmdU7hUk5gmSh7UmX5OziCK5WHjfdG3FUMMmDtbWW6W
LYxAouzHDHAq0S8e3cd0rLV2p5LmZLXVQsHKpIbaNnzsV6euQWfLYN176iANX+Gh
WZlzsRIINRtULHaskoV9o2GU9CTDjYCnxnOaiZOYrRY5Ivn/TQxtWhYDI1bAa3NL
l8gueKjYrRcUtBRuOHPVa0R+fVycMrMhO6u8WhUDFPrQjhH/rTkso7hOZjmQf97t
UBUf4ccCdfPSSmo+xTOXt4qL3s7PXsALPpD2rUMP9+49oCo0SgwsI5i2OBR7bHjp
pzPMUcY+l86g3tCOLBWgpeIWpqczhXiLJpRuYwrTJIi2bVyyeZeby+I1hrQnWcUo
8AFr1RtE0C2tNc/jpFOnLXKOepU2iOwBSj1PLarbTiuxC2H5uCdEPLwJh5pXJDik
3RmDcQ/Qk4E7I5AV0DK8cxrVqnYp+sgWnyrk8sUyE5d8DA7jx8KWaLq9EsARVGFY
DtuNW2NdxiEbhs5zPXGyffpsiFC8rLdNZMSxmcBFqcVpbkh3T33YRKCHuAVo8DO2
ObaDWz0Zu5LDkLCoR/N7VCQHSJpSv69NF7g8tyUXQPbmBAOiduUMVVrIamOTMZ71
xoM8qr27opWrrJ/G4gbZZQI03wHqOwc5KpOqgiyV1gdRvv0wsiiUNiE/YLUeielC
Cz6gQf1zW+G+tRYlffMuod8PUViFjNoanF5WusMRQ8pwfVriE9UuSiUpB42iGS1k
qyvEsR7CgNQStqj9lz+/hmOMnOGofhs1cOeCAtQCBxET7jJixukjDFlzj3ndW0An
gJxS0zNMLbvsFl5if1wChKYGvRg58z2/Cm3owSdQZWPGKSReW7eeU4VCguqTFnio
9qsVIimSDkUzUMczNioBSnnS/f384bDUOAdFqBtuvbc42lb+3/MWg2K3Z+vLl5V6
754/NBf4PF0/Dzcy9h1mAn/Fgj1oh5vE+Po/VUDftSCu+LGAOOZH0ayTbeC4kEuI
7jSFzwtrKnc/djVyZgtKUtXQAHFVX1sQcjd8wE4M2uDNN8eLvhVUpIFzWq6Y3Re5
RAHcun9JuQOTkwUidMq52MizAVSq2Aie3GBPOtTklv95jvYnvW7PT0JbQpr7cnQz
+8MMN6eyJfZygJ1UGd4E+6IEijS3fec54S72R8asDi64kWNNYoF18lhr8CxkxBpt
w2nEi72k2f3jm4k3BO14aFuuPCRpR+dYa7TCNOaOzt7hx1HykrJcNMHBURr7edA5
lze/8jneXjHuMCmjBHegCQ9bUpmRjXPCkNsc18kVSptB5481KnkVUpqxRijYdqUG
38KwXBXxkgZmJRf1uVFHKsdBo7KTaZtKcB25W/VMkm/GOMgWzUiLL/AOMIoV06XG
0g7/MkXFRbwXMiNbte7XlIkG4GxwE9Jf4DaQ1OpV1YmKp8WFi7EURrCKkFPw8dSw
oMYuJEmJrfNGiVFMb4A8FX/AnjzHr0QPqBgSRVYIskm8XAqvUxuL8xyXON6mvCQx
n/K/JoEtjEG6jBCVuJEdsdxNPQxmedHGCYMD0z6Z/aNPxjsZGVSL3YX89vcpDPgI
00SWoax5iu4ySS/KW4Ri6g4AnvlF1lj17LG9jUgAZLQZNYuxGkGq/K2/5QaT8/0y
4+f3O8BT+dRxia7EwYZ6PVF8mbCgHmEvQv83GSzF9v5WxV10dhEPYgRdGfv29sjr
X8ZZ72YOGfB5srQ8UO51/qU+irfLxTVaHLDVkmlE/dYFoxPFu25CmRKTLEYWRUAn
pVqrPxkvYuyIsXWX8DeTtvkDNOYQ3sR3wrL4SSJwf+7Lw27hgueDHUY4qahv9moE
+dD9lHHuMa4zz23Cj7xZTuOyBVM36+hT/v1KzMHRFOV4cQDwJW6HtiGuWZqw1OKk
dYx1PkQvUZMheD80kjILKpXLQ32bheRisBhd7ypAsC/giFQbca2UD43m1pEMSptP
EeYTTi7875GIHKfOygnNmTw9HvxPKpLSW5L4G6N1VHMWO7qc2w/2yS1V7eaiL2wq
zie32AfgGvVZdz5i7fSVvIPCv5y80ikJqwaqF70HrFIPd/YStHb3tUXx/BTNSlUN
m+ps7p+huGNpE0Ww+ym4lA3Om0E3Om71R385V06T32W2R8e/+IqBjoZBXpqVjf3X
vaCSmK5Igo12G6NsDRkWu4I/Nj73BGRVY5H0VajrHCxSQx4a3V4UmxHV5Ea1cuDQ
uWwvpxMIVhooLnunPCE/hC6MjDdDuiTRhorDxd4V9GsizwRPxqLG7moA4Yjtzg1p
d4ptUGWSxmORT9uHAHZeDCV4+Eve9rDBDL8srse7szLAJ1UDnsMUIcY/3r3jHXwY
ig4ssHv1n02XTAmQdoCFxWelJlvTzyaJeQEifqG61h8LnLqvYsU+knHyZfbqzwwM
S2YgBHNJd8tqc6nzVoGw1OlixHJBi3VfHpFNg7CWIPCifLBW85ZvduufmXziRCbp
fk6plz78fV8yCjd7ZG/tAQwgitDY4VWgQMBU2xDlX1doGxAgv0zwup2IscBs9kZz
OzQ4VKgM0PNJX7stVdJVB3ISllNU1dJdf+2GMHKWHCAXSfbXHUfcs8QWQq2Pgaqc
b6fC6XLxcYPhWPKNY3k7U+ma98mKu4hG6zK9XCsQDGTgdJUJEC1WCKsxChSf4/qv
krtuTmRFvoGGBvzLo0JaBzpUJOi+UELhv4271W9r6kTd7tu61YVR1LAYcf8gnBZ7
fwkdii7rj2bRvLHhTlwHXEinM0eLgBlRAsodR+aXXnbaKDsIWnVw5SC5Huky3sa8
AUP/VqkqE4Eq3HUEXnOG5RNhSbOfUhZKpFaaib+NzzDNJp0OlLg5bBawlBo66xa+
OZBhOK5tZQTIoLB3hXHEfKyWjZ5I2Xj6HgV3zi7pXsCFa1BUoS0ZVbzngBhOFNMk
Adm36jwOB3TmJky4b6x9HFiz3cpVRe6MAD4jPPcpnwUa8SOs9qRkD4zeT/yawrS7
quPH9/qx56iQaMGCBga9LhkUc3VG88B+uWPfHDv62HN+w4ryebmzjxa71pvjZbkv
0JoaFwzpU53Fht2JDWH9afbJhsRDT1mz/E+tzXw9xdpglAu8JeFctVzq++HL+JkD
ceJ1+EVCQPE9hK9sgs3Kj8LaYL4bCc3tFW6wX11KkrBSitRKWyzEd1D71tymWNW/
3GiAy8qWFQRXjx+o0awBwf+W9BMR7DaLfxx9BE9O+lAZ1nAer2MHBVl97xcKq4rF
Cu1aFXiO/IG8GOOkHBenZKWvE3rSv397FYWwIPya+n8deRHcSGsPkPFIjh4HWqKo
xheM5PRnU2v+0zir3eNwcI8sBoDKkF8alHp99kOKI7stnSa4T57pr4eYT5PBwHyA
pfqADu56gwfwnFW4OQZTNGMFMIiqO7sJ0y4WLg1I2fg4LGTp/NCA4Lmf+mEcP5yz
4wf/EQEuCt3+PO1+T2XDpPjDiNHar/KxwooRKtUg3HywTJaW8m/fTElSnwx0JSJu
zgmvioGP7Y0JETOr4e26lUdC0R3DnpaxwZ2C54m3sAcMKJmVMcCvnQpL95VVz8eD
lu2BgDxq1V6k1/xZnagySYMN+k7dFFsldFEZH4vQ1OWtlZ4m4DWlyEnF0XTwOtfV
E5Sw9LhLDcG2cxYQpKDX9gjkQm+nyROmkJWA8wWAhK1qP21sqVCX/eJZ5XTNcTV7
trO+qkyP4Rx+4AqeRQYL8JADcM0f8v1L6Wu7V6ya2dfPIjemLmbegCKmGGudfDaO
3ig6rZX0UmVo/wG42HEZ1PXZUNg/45p3IKRXkdzLO2AM9QEgUIWkVjZ4FRYAoDOO
+yk8tRpefl7f18FcTI1/KsOdyz9zniKdxHFRkOpHgbkpelWXlVzNgRuavRoDZJ2w
a/Yfjy067dNaqNIxoq0W0FTY9JRqBLiXykThFTKOB6bPsdHOMtQSWTdtOc7lVSy2
hWL66/s7rwtb8UuxLYGtmu0QsEmQlvICo2YtqouP7Fylj1PVoZmpQZ1JH9huj8BZ
HZ4FSQfiMwmXziR99TjBHeupKDMrb6boPRj2P5mQ+9XPUFs/G1Z96kxhGpKPENIm
9y3JU2i8f+HeBrfXfwmPd2k0Iw4ImswVOVDR4kNwCm2oEpIEswis1Ta+nUG2ak1t
ke4Un9hu9kkr2De5PfyG6OJ2ilhIKFI1rk8FgtnGgDPIKwlE7rCFKFp5m4l9mTyi
c3Z/ua7u9wtOADSHH8kLfYZIYn5REwu70RqI8poj2ITVjozaLvqUqAhzsLcjwXFY
VkEWHHCdiim2VxsIPVG4v77zNcbkTUGDxKtnQCEcjjQm1mQ9qnE/c9h6jHj/uyPX
sOg3spDs5H+U0Gqr68ilQr1dFqjM8Bq044Z7WDZZ2TRrQYHyLppPRnQr3x0K3iBD
+Ip7HNjE7lkRtI2P5rhNUKScJsKz1cyfLvx4p8Ji4kbr1+vSImlCZ0eZtNo3v29T
nkMXTua347jK/NGDVTNth70H22XRWZCKCwOhfmhKcNDFYyRPxjpdD9wCRz01/28r
NnPQ42P1aoC7eSNTTksLAkuGUsVC1D2hoP1sgp4xSQE2TOxJbCuSe78SnLFtLcp1
kl//oxStzBxgVZGIxjMDHyAE2GEf5HhJ1RJ0rP0lZQLfNcwwprC+zyHl29bZxDtk
ar0/UnFi6cvp72xITUw1QER+R79awdh3wLhCNtpq9VRIHtdaen4Vs4S2RXKLCA1b
CnGjJurfj0ml5wwWu5qYvS/qsAwzcGoKdyMwgKiXir0MqEP9Shrm1FgmXWWHkCw8
EKDcCZvB7VZxHr3eFN0mkcBMStfw7Qm4GIz0N8zyCUmRLfNbS1z9aAw1/qk8JQds
oqA0YVbttGB1VQRqTcQtCkp6awl7whXBChCrJljvsKuXuFrueMppbfcB/Bo3p/h1
zoGAy76N9GyhtCXuhUc+aCxj+IXGeozLAEouSUJgPkkfk0/Z1wPyQTvnQCGpcNoR
3Jrn1Qkp8IiP4KY26eudQmWSgDbBATJHeaF1Kebpu6B2Q+2Cc0GxlWr6SGyzRZEF
6/l/9iKFVBGtdQQOKHGVSoL9lOEiZL5SSnjfZiIKcVULjkuYAjy5FhkZ0MclBqIh
REJZS7bpECB0JFIE3i7IF+atEvZrpq+YUCKVjfLa7/GH2DjCl5LSIW0QV971CTuw
SRMHhiQRhCUEGOYzhZwdyNp0ezFIM6yzqfnpG3MLbZ4A+olnRxcOSamx+vnyHJ7T
KRKAT0vcv2+/TGeGAe//6eAvkx8axnp1H8HUO9klZPsdMRS+6jHloIRC4p0+uKSC
YI1P+I9cWMADthvQMMhaj4xuoWu/pG4IqIJ0geysCZgU9KfBQOug/58jEILI3sUw
6W16KGCKR+/QuwIKGNlMOHJvWmPZJG0jL3EOYUWl2+zCZH813CfkIWEaX8RRCtBK
VnvFzYDYUXwYryPAN2nfRob5m7BN64tI+86eY3DcbSzV55gtvpE2NL7wEqUGpjrT
itT0v1bLh8NxL7a6ly7pDTieMClpZSvXRtvm57Kr56YgemBJC8n8QrbH44aD+R3k
9iOW46Xv5qL0iQtRi7TnNKQzB/fhW925czvoCdrchDdbGzKUNvhAhrSZrT0/WhiJ
CznRik6PLr098DMHcgJ2HOsVx8/IEuqa9rYJW9RI9TfyJ1BOQkll1vsihJVqfIPP
QZUBimS2ovY+MbirMpgPcJUKIyomnLhAHQZ6yAAJRhQmGBBTfGIJApifUyHlKkhC
rh4BehK4X7hQcM0lmLAkgExXJXacPQiKL2ihJEMiIBwBTLZHIuGQNTAIvFlNxmYW
2PSwd+OXKTfFmjnupYPqOY3j4+cH/ipxUVwuO6bq2u84claMz8l7vrL3T9nNQi5n
5AjDfu6dvbUsQD7QVd++u9yncoDPLLQfuMNgT520nXBJVs/3yuyAPlhF2FMXGnIG
Acoy8F6Pqy4Fb9PXlZVw48fEmjmGr6fHMkhynl+mItAkjOJ/gCJcfCeEcok+jhBf
2nEDZB39S9zI7LBXo9bWN6vvckLE2nv3mbM6UW7fOjaZuVzULWNPf23tcu7LfqIx
NSdyWppTrZJnva78IVLQGSpEcue75iVjVLAsmYctTWIuPY97h4eFkSig/bWMeER8
pExyUqDEzOzgGF2m9MPa/02zHAJvRF3zgGouU9InQ9Upel/AHbTc7mSwVRI7s1aQ
hbOBeXG3k3nrvo9Y5be1l1DrwP2Azo4X+Ix/o4RNNmeiIeLjHaQHuV1b62v5iZ+J
ZZGrtlkh0l7XMuxOk+seJvyg3tqmi3to4m9rgYNTjYkCiHM9uHoGFrIxUSpcEQyO
FvjuyIzFLWlbpmNuMyCuWitRZ8mBP3MR6+HQgvdFMAWarxrDBj7SF/FJRmQhX9K3
knxaU7aRSH80DRTfcgCCIRXFkktk3lcm1hLtN7VH/uK4S1viAhQkuUOniTWArkfz
ClgkWmFi9ggr4n3FbH/TU9VdQGIEFgy9ruql3lQ+Y9atKt+mEUbTg7ypfsHHcNcs
HWdImkWsfEX6g8w4sUXSveOtJeOXtxHOuqGqwL0pi/Cu3fKdV16GkFNPR0THGI7p
I+yiYB7ByPIeOUYmVQQ4MZM0RuHY16bAwMLy0jjda34Q0Z5JEDAnjO80vZjucoHj
B5iLZ6T9RycCcTWKulwLmqFaWqWHkmXludSpvkR7z/UIzvUCy3IAK5dcJAZmlebn
5kgHqDyX1FH2fSrVoy+kgpZy5PdZADuFe9j5O/rWCT52/14g1SlopJy8uMhMBDc/
/myP6EbgY+1UE+bxtsbLSbXHxdkm7ynWJSg5vQfXSzBXquRAdZyXZrrNa/KaUxj+
QKFBB4JQ0goXpQiwgcDnSZ45MvqPFL83tYhQQrZE3NX6zTsd3qVmouxuPNkl9nPQ
WqUS82UGhAaoAFHEtME0Wy9ZIOCc36E0AgCyTRjHJyqm0adsvFx0PdGPYW0vYr7h
rBBZcem7qR4A8p36TCJFNhZZhL0Mmfi5z7+uo17FEHzZ03Gmbfogo0IsEIs8aqT1
1jGAT+6jH/Eu9iLw73z53y8SLhpu2nITRfRKGCB5GUJVqGaDoazYfSCzEstZJM4Q
APz5dbyVk5YZ4TQIk2bHLT8S1LvyX4HSnGOVfr6aAojZA3JQuoAQwxktG8vK9N+y
9GuAXWzhNDgiVkf2b4ohJ1WZJIC1Fr4gRqXa1alVnewLghxzoFVh+M8XwVtvTLGZ
+VsiPfAQ9BPvdo9jeAg9mDWoeQd9NsDqwhyiWKh3CVLOz7NeEHjGbmAVnTYr1W6/
MmGYJWB0ls0Phz4XY6Inf05vffLgY592iLlleqlWzIG8cFmp0D4vLPob9c21cNYD
/hWG0Qe1h/cCakB/Xav31OhqNGgYtjoltKBS6MAjx/qCKWyor0Rxhde74cLVPe6x
LeWw28YWQim+RrsQKzKyYaF+vHdbn3Ehh4Kkrsz6rat8h3w3ry5F77pWNbB6oOac
QOKMM0aZnuCRsS+sz05iSr8wFRvO5hLeMEnYfftnxVSbXSTdmmrfQrBaECgVf15H
xx2fwl8pjBmOIAyu/+pFObgZgVvoM4TXSH9s0BLy3Tt9Z6WY3VzJAhd1chq6HR7m
Y58OJXcnPjoJdPS3brtHGp+qjZpulKGamCg3LckGqOOGuBLBgmVg3G278yykg9GA
JFIPneJtM0A1xAVCsIfrA5m8XhZWioIDZU2NUjKVMZwUp+JZvVwYcRFz6iocQdhb
Vz3sUhQDspUPzH8S5DBFlCr2JG0NCGqEPEyWbCQNUxXX+UIafjT9Vmm+LDMlYyJq
VOMeBDy53WdaUKWLxmXvNR7QTFZeXMkI5/L14Ab+WZQ5/noIUIjVKyfx7LreRd9e
Gy+97F5QiDYJafCLjupz+Q0KFvgAZYKnai77Qc54BMOZ4iFTshtBIz9DaX68n87h
OCc5H2mTPJu7fEF/BkxPxECKeSd/QQ3yYeLGEH3xUVsqMYFvbgRrxWbYwMsC4Q8+
+kV0UiMDjo7qKkVn6GxjnW5k4XTOfA3HpUQ639IeuhF8ktZ8T9+N9uawrSi6uQ44
onbr1K15xBkMVCmyzkDZem/FOssczToyGU73UNkVpI+o3LfvO/e0+UvCXAS/NW76
t2SzyZS9WXtWmGhDFKAo3vvai871a+CQPVb38+zWa9serpWsha0vi1YgKmqhtL8D
Li7ItrfYxmeBzv3QRAROmjpNYR5pegtJkTd05BUBUFafd3OxKBItZRbYKVc/bTja
H8rpFZmDeyCtyhuuFI9j0tBjm9ybm9BWfRgKveYI6w5IGsVlCp1TDbhw+L9/6UXR
ukrug2zyJMb9wZIef4Ma2aRPRletKF+PGZJcbi2NAEaYCdWCTEYGIe/fotb7ZcYY
jqnhO++BKfwFFWYMqt/2jqc4bk2qzgTuUVieH/+JLPsd3FAt9pmoh0+VhcQF+jIl
5WW6BoT+NiCyl/Pt1P4+QOuP9hgyrpNT2Ud+rOdrRRfEdjOkne0fNHlZYGcJSlHg
BDz09Zo/Nv9sVHWurRazzBBWiESbhM+Tu1OoB6ATHMpQlb2LYfPnv0uGdk+0MiZI
4OoUgAS3dUVYr0MtZC4uEwjR/3wiIhgbfgUMZltwxESwznUPRQ3XXn9XV868jkgN
XsTd1wroqHKsmL+fyOtoxrH6VVCWehR8rR6RkI8NfPckbLeVhe97UY2OBqDjq3F8
9INuIVXI55rsFMrLCxyqbIevEe+T91eZDqWGs07NqrL8So8Uxtx4nUCCJK9KzAj+
E2KOdj0duyLaXhJME6/ZPh4Aet1FBXBeAr2vRB/+Ft3B9Kk8nLH5YecCpXuX1fcT
4jqA6Qp2QQ1uHceP/xLus9ma3ozH2nIc3ZBhy6QwOQW8k1b69NOJj5g6Hu66hf6Z
6WqRWBr+D1lHqz2Sb2QOOWpO/33t1Hl2aHTEJIbbk8PSYUmv9dERebfEbawseJSk
jjZMnrL07cUj6Att8QNHBAUnAXZcX7gbYojYJLLRtPEKzsXgsieWov36zWANY5N2
zjA+nl5wCIbmP55QqEvWpK1TP97yFL0TdyhljSSjG68LQIBWZa1q+Jij26HcGQWV
/1UXJPtUxaniDQZ6LXED7FbKxIjHM7CU/woUTf057sDae28Zxigu0aCSONafqmpo
prNwIuG/sK4ciUcbfgK1JRHMdWUWBVZakhI9cWFiBN/TEEw/lJJA8Tu9lMoFJQJa
8EihZ+o9sVx4NqOm2lBaycK6z+0ZTkvkNhfBRDkgTQ3vAq1cf+xeTUBVl9nsGYEq
i63OINIGDD6ZRoaca9QmlBLJSmac+1E99ja5u1Cs4iqxyUoEzdQJAp5ohCEKyuSl
H6zy6vQL5LNzGMupSVUrgaWKTYwOXi3S2kIkZXD3viKk6nHnDhma/PRVu1kM9iMq
GTgh4B3aUNkb3GVX8iLw73fF3X6bgHly4I3mRXKsKSKH9AKQzcRikIomyckHFoWt
ELsK7y5lqc+el0oBUV8W3BQ3/B1zQXBBmSPYmtH1hskPhs5IJbBnrfAAYy9sVIF/
zJKdz8JSu+PYF/XGCceSusZ1qce2u+oGdmTjOZ8jS2+GTLQT6ToJ4ZYMGD/p5Yim
qFavIxHGPBUX4GZDI4xp9B8PWW/CNtg35FKOORBvEM58T5pBhfQea8BsULP7JW8D
yX0nQVeG5D5WqmVBcCe5ZPDDKVuSizS7vu3MaSpD0xL3ncV5pkk6/mlKdzSQ65DA
1nc9st7JnU0IWCQbkBBrNaOfleLMb7D9ObNFu3H4HyCJC69lkttm2xHTThvhH7/U
4M0cd0cRVmvPUs3fH8JFg1wj1Tpx/+GZmugCodQqYjd/rcHoSCebKhq9Joeml/bE
aYbhXJlkiL0DRVrkdVrP2sxfq7vWDNFFSgql932pH2O4DDQFuBuiIwPD/4e7DZ0j
s0uWlbJ4dfr0eN95Hmb7/3MFKeXsQjxM9axY5tt9ctywILUeFwFeA0vKqWUdpqbA
/NUB57f8PWicAA8AHbNi8iQRVYxMZ4UlmkZEP0rAkDnaPv9nwbHcGSOHw1KL+pZs
PEPrsqg9F5IsAKd0v58DBjw9SEdWb3Dkfx6+S3mECr6Vbz5nceyZ3y3LWPfGm1Dm
BVc5IEU3M3gg+6EtbQjPEGuuFove3GqBzvvrunEZ0Nav88tZitEvggCoCu8MOWZr
F+FSRhYUGKaErWsq2wr0q7PSMA6nPCMNLuRI49UI97+EbPkxeRvm/aL+9mpt6XYg
XlQ/HnvD09/fJmJ3Jr21qYcw8G+AFBWf4fRXeoJHS1tiXExmHUUdp+EMqu7fELNf
FKf0UpnQdph0G8EcxpguR5QUIk72TkTQY/QTkm0x8zkLuGTFfyJSHflwpH70R+Dh
A2xLlreCTJS6zAM8psL2i+kjLXon7dEwjogriFSUAtfxCnIweq4EMbYpWJgO2ZoL
bfhlPiyscgGnVp7JUaQxFn9ufBJ2mMifqtIdwjoUIi27AAGOSHwrFgbPQKmf9loQ
eJVFTh5jNk0SMmQmI/kHCEZ8++aDon7/uDhjm7JyTt5YjEh3R9UKOidX6YgRxmaH
K0xpS3k+OCEvP13YqSzNGq93NL5M6XQLdQKoOVPEjYs+A0FhccvLFOHspOcVUCoJ
H3OVN8HuW63x8qP2czI9wVGxjfHNjGTcC6Nkf1YH4tCmY9DCxcicKF7wmqhO7chb
n+ynJkcMrulLd4Rx/9EFrftxroKKWf1Y4blgWRUKjLoXzx32TO0EjAC8C1FeMkmd
/I96LBVNgOKMb/6nnUkHj6F7potbJGCP5ZVyA1bCCszeR8T8uWKxAwtlSpNyI5J+
AKpsQf5Bmaist19wTxT8y2yvSppPjod8HgHbjdJf17etc19a/Cu0WXBoVJQK29m/
x+X/HSt5YD9z/kO884FZfm1jUJrwPwvUjI/npgDdLZqjvb6WNbCQCGKYMKQz0cNj
MQ0tOna0UYCH/VdIoynUX571YcS3q+86zb/2LMyqOYGmP08O3is+Q6L4Ttxhdabe
5y+Gh94cQjBbu3RloDZ92HBnEGp/uxWH0J4/RKoOv4We2ZkwsAnP4XouIm9YuFaM
CdESmpylJfifB3sTJAlkAOm6gTmESJDbSdYRxl8bPibZCdRDQFxvLENItla88voE
8MZxjkFzPzl9o/50I5cUQHI8o0vtHhwqc3+gz+V+wspwuN/qfikS2Kl6raYGgSsO
rGVm5aoqvCREKUUPEDshPNZ6p2RQd/oN3MYiyeVXKADASNoMPj2b2TTU6Ru9tBqc
yB3mWCWjrMwbAoZqCgGqzqRLCiDVMF5Q/PlFIjoVyDl1bVzlIGAczSysw11yRNmf
MdA+gbNmLEKeALB2SS6BQe/TbAx9jgZrXf3JaynUSNJPFAeb0GEaq3zl3ZRDizIa
cXgfHhSQ4fXeKU2U3xkyWkylczbo5oh+cNpUaWbqwYEE3kJ0zQsVd2Fkr4CzWsNT
0DH71l1n+8EVmUQ3kpJhcWLN9Wv9cv9PUOMLlfD7HsVrCFaWlLgffoeKDpKT5Wiq
VVWhqEBMv3TIaWxhjCkrLnEK23z+2nY406jxzueE/gjwLySe92oj+MITLyKnBIJ+
ABIAs9Fh6InCh5+cgwqLMKPhgKyHpMb2nF1UeGwFsamxMQddthtCa3hHHg/XZn2I
NNVRi32bDnPnC0ctB/wsXSGg01Zaznc6Bl5SM1AuFZcJY7wVM8wbm1ffh11MVAfA
/jhLMPiYSvgP2wrLE15JCv0AvcAmrAvX6/ALh3o2hb7LKq9bV61Ls9IfbfIbvUt7
3eCf678bcNmjld0tNllxjZK7BewGvF8aB89r0DOgRuzmW2tZbylfpkCsydwT8zG2
kWWHbmqHC4n+OhpEhpWRp1E4pTsPqHDccZ7zS8GqKlKKOHmL+7bHmnYUxDy08dk9
09vWo6m5L8D226yix4b2dOWT4HarMIW3BnZfAOvaGkwI8z1FTjr2sXd3tIrIxS5C
vKuBqwLy6NjnBjT70YHw04rQ9OFV64M1oTN3h6eUVm/Ic4p/LbG6UKkyAbSmWf2j
rNxDjAhQMkdKxhKfJ7HbkATqit4jnRX3nH+sqjbmzpThKUfsHqi1iPMyb5I82bpU
HEuHbmJtj9/VL9dG6pEi/x8ggdVGq4czipupeaNj40uPddvMaVbwEFBgxjQq0WkD
ysnMaCjtOrtGEuvedTt3c64viCdopi+vv72j5g1r4tTXnBiqJA8HBwvEBFVAU7EM
Q0i73t0/yxprxNukAwHYRuIN/wsxTLDBQ9V27C0zamJu33ec0bjSe4O31F1JRYcS
b8i2h2jJpAGjAw9PABU6ZhMmNmzcXtAcQ+iiAh4GBcoVNAeZDCfj2smfAJC6ZCjb
`pragma protect end_protected
