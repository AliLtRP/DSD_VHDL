// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DNQ7EGDsBMm9noQO/C6+VkxVZ3dfhC6OYylCaLSlxRxEo7AMoVmuBduOPf6/C9I4
t0eg2NPttf8lFR++0nraBz99hQZ0buKVDOgrArene20JNjhJ/ZEx/7w+xHeARSJI
JDFx8wm2lFrr8pD/EI6dsVlAcnP+cMEvQijJoFDFH78=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 83008)
GF7tXGHlb66+biUm7I8C2YRNU+GqO7XMcFZl+/lAe4n52x2BvorDISATe9c7uL0o
e6TLKlXT8KPNJtJBTEIchZrn2PnC+9xxJU9htDi34EqJD/HlOW9TOvWGuDpNxYix
AoKNzPoCFvcy/c2EFeuYY4Z+Wul5KFcukJz00DZxjRd18wFPxkNxz2OT42VCQK2b
8YOspAqrdLtfZJWkFXryn3NmG2upNvJ6W0pxHEbBEy/gLe5GOFAkbRHRW6FAuSvT
t3Hq2TZj/C0yOx9Z/UaOohakBCbXp/BWSRVdtjXaz0/pQX5KN/hcU95dY0aqCWQ0
eqXGuxn10DoJJonuMzO/m/E0M2+8YZleUHxlbuUdQdb3t+KcVj/5fjEcRxLD5zDR
9cuMp1FtxrzQccFtQBc3567QkjTovGyfH7WNc73pQ5tHKDttrdfk+5eXoFv1Qu98
RUhO2xyS0bEzCZPSkVkuW0MEGoCamI8PkHGFDW8ejj/TLEDNGILRZcHB9tS0nOa4
0s1JLdLi2H1lzIUskpGAV+2QB3DJpfDfg18TnMghwoWhPW+gVTjIUdiBYQXOJq7k
crqzW+uFKr/2ux4hZheSjxJm3udMcAAhMlRBQveeh94CivaIh8SKR6B5ZYTYrYnr
FVIh7jmn/XAuXhjkFAkBmoMLb75+di+aX5YhBXl1cfwbTxPxZzt3ESXLxIXG8Jd+
HIh4N19rWGMm2kSY1vgytIvP8bpW2Bsq0UC4k4iMctFQuDFO2nDH01BsG99HvVCS
7d7aTu3A+J2+VQGYrDjo1iWuLJsTmZtm5ZLPOyIFhRNn+tR9/Y4fnoAPWQF7bTla
8BHoO61OOEjJq/z6gB3QE64Pb32fGpmVbVmYrQGx3zrmPBqKizudnsrJHCjRcLpu
EmQ+58lvboCgRZwdCdDCdpN4gwv+CkGwVOYWHrta2z32/hlTehRGeB/MSLzqajtH
rSOwCgasore5gx9IKxDy0sbiHI7+T1hVFHdlVCqiSa744fVL56lBFBdBuBuLIPQr
J+yjdc45gAKJizbUZbX2+oBZCIKPLvfFkwqgr8QftcAQuWzsfckVBDWrWQpHzT+h
u9SVyBvxX74gg39maVkPi/co1NBvXshDXr9OPWbCNWjZ2qY7vPm7yXpu9zGd6Fmh
jKwLxMVjWBF35T6ppD9DHylgLtjiU3oACDvSnhZc6WQi++U24BCADKnyLXfNx4sk
p+dQozYrShl0I0DYk+33n3O10PBlz4auk3YA2G8wlv4dq5rP8Gr/0iJIOcLFm07K
dPf0Al6Dvu38dN95hCrwICZZQZCOu07SZQJMiaDLyoJA72i2wHvyJgTwCsMYZiX/
AHj1/jWoPAnVtM77vmgt0CxxOmAZWxm71knoT15ORDM7gsMk1bi068GSkkEeLUy+
qCpIGmbi1FjPHdUln4AeqytyLfd0eHyUA7y76vciOj/b9aJCpeT+zXEHx7R6CoKh
ATfXlI4CDN4+fyO0ywPhGPKGfxqutoefqGbFTV7DX0tXPJvNXzZ2Q0ENRCnY3Ysa
3f3w/9Dkmhfe+hmVNRZq9Sw42hNuHDIJzSH/sm0FD0HgvXNhJfcgIk50aAya0VFT
ORO5xLzB3M429Dao7jM53+vD0rCoX9dqxyN2mvRLXsqMRtRT1BaqePeGJuNWt0Tp
o3hnXUthWeXyCrcMOfOKTkuE4FYGsKfRvuwXw/6Vu0jNTHpWI6jIZZB/P7baZVrP
7TnCe9RIVlXjzH0saMoi74ObRDHs3QC1syVDslDZG+9ZEiF8ywlNc6Ekd4kwZlPC
uAB52zmpge9ZZ2hajPcVaBIOeWNREA9NpBAtNiS84n+pRgmU2NuIJx6NXAdGJxbC
EymW1XcoiqUVfwn0v3c4fRCUzGFDEodmcpDR0RpKFt2KyVeeDFchM6xWFdb4r7fr
pwSAFdOLCRp4QEvyqJopdlnNT7O0TLkZnwevi4D4bkc9FMYhBFCW5NuAeUDa5zcC
95QchwciZJGrGpscd2vkW+J6iYSvykMkXLMFBmvinnaCoq2p7MLdEDHOD3qUy+X9
0m30NvuBxbSzTqlFWgHlSX0vUjcQlZ/uFBQqVLUlbK5vNDUSaU5CT0gZ57TVioIZ
xXpXccNfOX56mMBPEYf/iRKKDXrmvmLFulWvroMlJLqvVL5wg26jfhmTlH8Q6Mg3
RrDu7fQaNFtsKRVICApKXY1wfewmKzvgheUIVqz2IGbF+Pj3xdoetyo6JeqwyoJ5
uLqkfcPEkotTmyLTSrST8+i7eaEDaCGO/1ob7aVpwqMxWkNoM2KQ08cwY35S4yfI
J7nfVyIx8TjWJ5Fa53kZ9MWldO4SYxFj6F1Af2dOlgNJeCA2TxMzDm7Ep0P6aXKe
uOjfV5Jc2s8/qD4L24XGKSDzSNr0UrjUN831qyTM+4JLbkI8X3FNFibauWl3XSrt
L9vFcdwIM6hcbkEeUBg1NxN9q6pDNlrztpMAexwI9Bg2W5uf+H+W4im2rPvh4IH/
m+RYnxRdoYlF7m3WeoC2iJYb07yWa0cvtsCxpDT8jFYoMo928W77N0IgkZrLvzHe
GaysrxXUuIXkPRFpY4F6ujGvjgLo81aCLqzvpHh0lxXoH07IO7jiLgSdne4TEV8m
P34qSnBIxZs/kzuIhKQm0ZOUo378c2cxDqlw1I4zIc3A/CSuOjVosoHs+Dh5FaB6
3LxjJmImGHr7yVn08XnRvu4VYdz+Ss6C0+A/bf2R93OIKUteSnwWfT/kwLW5J4J5
jJTU0Ekk7sP/6CoePXSx3FtGHBXIgBGqvxhdpdkXn8Cg1sn0hV4bYPUSbVtzUo+j
hNKQnR95JZWp8S05j3OH3bqyH9/eplx2d9dnIP46cjNQ0I0DLwrH18O0MAAKH8GA
G8zk0oVfKExs7o8YMhPPtrxyPEHval1nAWioLZAhwlYhaL4WVba5WFdeWwXqYCJg
RK1J8H5UQUz1m4gLx08TbtzF2OY7HqqVkP1ZPoI3T/8DvhmDqnvZSgCZfT8/PixT
fw9OVkVoCgh0I2VxNywRTZUa8UyoQ5jLftMpRxN/1J2PZSKBd2CrkBydn+rlGPcE
W2K9mzOhul6TCGgLhk8/ziNXdYw5NDPu8BKstU5vNd7NF3npmORBdSm4Y3L+GFmU
wqXI/HcoK14gyuAjXHq0cw80ujf0CnaqIt4Ao/HzF/zgQaQPki+Z/eRV/PV0RL1i
bs94LDx8YeHmg5H0idNQE1KeJoUuF/28fSle8W81H1iQD7rSJqx58wzN3WBJBDlo
cAv/abQRu6KnT2egaO4nC/REUtNONiFhccuZB+Js6ufTO/lvasX1Xm83qatji1c8
N+L7a+gbzHyGkpGMARSIMYZdyLCYw037mzEnb/EwXmDi1wwAOzE5fRCCrNPNDEOK
p0Z+bUAT2Sq7pEDR4RJG5y2jTt7xS87X8aib7E5e9dvt7RwBkt221kio6SJbLAnZ
fA7Kd/s7CnY+qonpOLuGL739QDktPFd2hvEYBxcEg/V4aUuNT30kRWlACZHuVwCg
nT8iujjO/WyEns40KQQIjVf26+hKww1MWDZZ3vDt+uY43VrcoyexTToGUOr1JvMs
HqAV3shStVQ/W5FryQt94K1/RZxTH3sunBoOJkV4JQYtTwRlD2Xqf+wGFdfzw7rk
9izxmv/zR/4kKzYf1Q50L74+jWe/rprlfQIP/E5B06ZuxrGoNGfQtdIPtoKI0z+H
rycY8ydbNyzNtPiYGgOGzdAKabdxSyVlscE25yTxQVgk4VqqZbppEC1a5Qis44QB
cDDRwb+GqrEPK1eafgr4ANKbc1Pb7dqJsCJIOPPFh0eN1pSpQseH0mZ/Q0z+XI6m
BmtcA3RLrgIj8YvsNMv3X58jprre+oTDeg1NKTWF8WOcX3lsZhPfvaI8mk3hQZu7
aVtOVTKXq4UvTVKnr5aObcL2X77w7uPiPyi1uuPB+8gSl7kSg4/aggwpZcNffnpt
mz3GOjoSJ8GABZ+HE139of6rY8OL4XTt8pIAvNgoDeCLR27VZ4JHjHbqyXWw7p1f
F8knlD+9Wd8BgKDXOOUmFOYq0ae8DHMZfEJ+UeVdEsbAVBwzg+fRtDqpC7GSp5N0
KgTSHKwF7JLD5IgvWnKJnRi2xB1fAoZoIbALSYdNhDtDInh0pIzIHtYEh21Wgr0K
jgiXV1CYpSNepm24LHqNBVBWsQMXG8N4vOnRGJvrKw2fDhWbIKlrzkFj4WIXXqZ8
/6/1GOM5RL3RdsJPakV0W3PzqlTP2pBYbIdBmyo74S8QoevwRJc/WnZ0G3M9Malj
85fxDtWB56Nj+AYKWgqWd445S2mi7MPr2oq+RyBoYOuv7etOVBtTe8QPRwbMoOfn
Z7lzw5vgyQ7WepaAT0rEdGPhQEjNVAHQ/8fWWvlb5KzfH2i/vyr4mKc5KWGSnDmw
NBFAQGU6iyLxOVImg34xgj1cmdQA/6WL0QodckYA4ZURZLIZtArxY2/GoC7Mvp/Z
makcwgMSqTcQGNfWg8ScCzw9iLvIbk9hhEmR6c/ucTsARc0gMhIk1zwGSpBoANds
Xn5KQH9TL1tusMHmPfrf35G2bNBZNwJ6nrbaVHKO1fIV/y851rg+EFwX2Tao3zbV
dhuxan6lUICd9t4/gJ/tg900b5veaV16nrTvzcdXKOZStxrzN/endQsWNS1y9aaF
/iwXX/+3W/y0tkrzPszh6DN+do/8KpzGiCwPD8FHNVey476izXazYhATIspIR2U5
noUOtq9oJpEH9B/xUY4DUKO+q5FGgX6oYAFpB+1Aeaur+HbR5u6YFcNhMFv8wypS
S6szNhaUTtNwFgWP5Z4Bk0FRbaRopGNSfLdg4OCg+PizlHfSk2AraBwNklWEhzkk
7eIycMDOCOsnQ4gSmFkgcDVqJckZ06n/vmKmBX8RuX6uCOB39EAXanNR/ycW13fo
wdNUmMuRP/vcL1uNDIqOu6qxFtxZzMAT03K3p3xU/v7EI/5nhtk1ShOI/l+9lDfA
GJHeUr87HRc/N3fr3MhSqsz4xbvtVrNwklfp57rWAUuSI8sOsITs+R2DlwymfQva
ESi1ZJRVUrg8ILkUStxPjcfBQdyJDDBSlNpiOiKmSf0k2EAZ+wxzQPUFY96+i0Cr
/kopFeUUOYF0oWn2+GKO+DpBmibac4DnMZTGbBgtmEQjuGBMPTLSN4cyj1ihil+d
J41DbBv2A0mx3DJO5Yw+xitULDLJvy+rB048lYW1Xb6UUiM4ej5nxETrYILF1neO
XkA246/pPkc5iQ/weaPgC6JrSNIIwLBlOSkRCBL/kllWpqrjloHcDr2aJTs4G5mO
XrMhHzA/dqMnwW7B2jv4VgR53tKmr7FpXgUSEM3r6vyWOsu0ohtiqOS9AJ3PPRiy
xS8nbL6Gy0HAC0TsfxRkOR6m+Fw/jaLBQT8KxiJK5jgELRFkJ/jKmLVlVFAN0N73
gvUyyysjnqzyI4Fu3T0FAnBFWRvaKka5Ljn5i7yeZuYHnzFNVKJc4dj9P+cPx/mQ
yUogGa3X8qtMjtr6KJW+wRHf4wbQkiPQy/189ZZohqgRUp2nVywR1fjgcTd9HPfJ
K9upku6NGxp1o5lAK2DYdc/z9UTPjqrMwEqZh+FPIMus+lrqh/RfVkXfj7VHQJzz
bsmlc12o1EuWXWm2lTiZ+D9hS/R6M1PAYCvhNtuIMEklUnQnWPd3GfBboOStSBjR
hWxHCFxi0uqgllppHbyOL4N8aHOAlfwl0mS4Q2nZ2vImQ6tJwPUo0Hz60F43BEZt
vKwTj2HzJkl9kVFYZO6OWAjhkLFbWub+ALN1lbGH5MSIudkiSeCmYJHn0vEYDi6z
2lelhbv8D3rg+L1OFynaiBVZhWq3BAptQSpj8AQ/E1BCQAcRmchfl0+L3XzlvHiQ
MxRDlYcuvj3DyAsJqe8bzmlcNFCpZi+U0Xw4eKEIP9h+DJ4zgjrWVxHkq8F/L0PL
QxxXQEAGTUBEIU59dBBYoNo2e2oeL6WI/f3zO5lw82g7GEA0ZDyfqpVjchEjxTMx
KKh4dFppVY7Jo/6HbavHa8qq3yvm5usDL6pxMSO4uI2tBrQreIXCLwgnTa/g+4pu
Vw5Oc+QnfmlXW5CXffFFHwfyXndYRFWp6IsA2uGKHRPKLmmXGtwIPP5GQ2J5ANc/
xlhXau1v2hjix1ZIIzRBzTzZ7+q4ec0RFgfPOzg6bGR1QZOUs3jfxnoKMsjM7ESV
N3486EZKRPPw/bJZJfM6GAH4L0qu7IGYYrsWXjsAkx8kb+iqW0+7Q9iR2VIr09Di
jYTn0G3oeto1F9If89F97Z1v2aJ7wLYRT9m0AtxNad/qo3oAEePIinzWZzdggwA+
AV3bZTVM0/lxgYjizK8Eif1rFUJM8TAfVbzTT6MgI/0xq5kbHOiAkuQqu3ojcTTo
zSY+2kNbERQWRBqwwCNgDsSFKu006Xl5+RiRrVxccQweU7MdEObzZYlcrfElhfii
n13g7JTER4IyQ51c5/EmyDZIiA/3O/Lur6fDdIx/zSNE55nx+ObOP2vMS8jlgpa+
ZcAmZADn/ShLFjpFm8JXc7SyAXp7FyuowqECLvbAnRoOhuMLCesFsfRl8eyH1HXm
LHmhJesELuVxR2TmB3NCv4T25PSx4lMLDN3gYIFirSPCMNRXjSytUMWCXDgdcos8
K8Wza12pexEi7vXcHgfJuT4kZXQAOsD5OpXiYwhwSUr8UcodN7ygKjnizgezWnOV
l1YAdkb0xPak0RwkaduV3XiuZJ0bYPFdPlog1NC5nnrKYxEMWKc2Mm8lgDlQQ7HQ
94qis6Mm2aw5iwHlgxgCdUvqzzjouggv61SqMK/YEfnkJU1peBGlllucXAJvI0dW
D/ACSBkA41CvPqfxGfbgHkvm8Rysc5Y9RMOtc70Ozz27NSx6HQ5+KS46kAN5k7CU
Wktu1B+glWUF3cmlff0pCKi2vTiz11HcrySYpXcF/3eWApvGgXZ6wImKtcUVeHYj
ndK2XDsvy7qMkie6S5r/25iO6MvTg46UUiq89euq1WeLRtkaYAouCKXXaBHeRNNW
iv/lR+XE5749+Pwi8Mk3P9GNlFkryc1sUTjs8EXvXxq0pcpGgpwjvZDONQpXIJRE
k6BJlKiuPW2nRg9VmhRIBa6q8BRUJfaOptKqaK2sAGjEHJUP64sHrUgxKZbgW2Du
oqKaymY/ZjDvw+sDPN/NK58pyJKcVnO1pfzHDHGE1PQkdagc6hK7G8JjWXnnoLae
2G7i9GEmyBWOrm7qmKbqVf1T5CZOAWGKof0GaS5GLvXYQty7XmJxoIerlpc/Qs+d
ugzjSJ1NC1pP3GkjwnmJx5NiCR9Y4xwRlhXqTLbUxkPaQfY53mdHkt99Alu2TY/U
ndGGfg3oww3a3lkgEIy21zIzyJUr3moHwkviNtw8Rx7sEQq9hiNV6tTzTz9sPi4h
AjT+aNAsRKAhqRlJyJPKgHUxhhUphzrOW5BUYBTMz3ezIcJUTV3yoZvFKaH7zYax
EvsYc+URR/MXWbXnPZTVivDiAnG+5IfjXl0Yy9MdjDArcHTRuOTofHffa6kI9bYj
jG6Cc5eHmeG0QX5ZtsgbIHQzEXxnmsduqSAs8MogXIiFpec8zUEValTnMOJ/W5ct
ueOaDnE+102rGIRiV7vKBn3Eu5Yp19DdGZtObXU1Zng3tD7zES65Tv0JMEwj73kA
yzpKWb+0iWRgEHI5m0y0WtZPGpx5GYbQvlulTtZrTSdPtMaN5jvZD8h4PfAG2eQS
0wSyP2qpKdiR/wWK2m8B1lMP7SvmGP8FdGjZ9IHnFZFu7Xln5BaG0f3bDPLWBOMS
ffvrGrmiV9MIsqYogjfDW3WE60ODVBtTIOPWc8MVzlrDBC5TgCWdHDu7T9ZwTMRw
5L29Zp30DazcCLMJJExv1ezvTvlc9O2LanNpI+bvDvS14XVK5cYOPlXMC4L0jBjf
oIJ2zm/aLwYhXWEdSfAqk8CeYl/j0opGOZJrgrYn35OsXFyvHWyBR/jxmnVoz82v
qFsYcjgm0ebxevgcOc1nTZlgLWd1kRf26m5nNCfHK69sdhVxSE0PbgjSZ04iR7Sr
gCiMTZoHABF3Dz4EVzQVDMvThAYcLIvozzYMT9uYxNZUmfJ+QVaEXzBncnev5yJe
ypfa+2mrPMZ3hK4j6Tbh2WoYYhKU2C5mgGRi45WjGw3mk7YFXgHvmpdXI5ZiP4bC
ustUI1k5GfEEpPHW+scp8Smrgi2o6X6oVVTECP4qoVmMgmwiHOgvyXabO9iBo2Ls
8S53+rwrPbh1XwGD1aYq4pIydmCKw6EZz9Z2q6Tdy3ml6FJo1OqivWt41fyWWH1C
+4JCZcRANn+yHJiIXgu4AM330uQ+a77kjPY9TRXmNXGYy3q95BoVvzYhrUOBr12l
5vjZgYwDE5Tw9V8Bp2L7ksep7o3U/wHsYudNNkFv1X8SgDyApwYhDZ7aqT+vHwne
0qsk4vS/hitu6YNegVjqkaTmm8N0THavrASehh3TSJrfFQ6X8QSmU/rCT3b9aCI6
MdXkO465YgKyrp7t+RtEl92sLtGH5qkp6gCzUIn63Gwp/DXrw3Ums0tGRPlcLIBd
wQjWch8siHox9td1sjW9slNq8PHyFoEVMspiJyJZ0bC+Fy9J48ksE0o3t9EYyHdc
yDEl4Zs6P4GEP4kyzlX0rkLsxrxDXKx1mnMSM+UaZTV7xYCmstPNLNRFgTu4l938
6Oqnl5+0YCZHtoCpUBmwa7UPBvMKJTr9YlGXVRe+qz1Mnn/aZGB5CJ372lb3TH9Q
ek6BMVL1578xx2UdmLsdyD43wQ8AMpB0rvE8sVK3b7pZOBf1IsMI/R2D0QPkpqwE
BjRojiLSwX9Lq4wBiKe3nWX5VV+EgugVjgFWGwsqfjCSPYJi0zRBD9JCxdbhQ3K4
lZwMegnzAq8MeR/9fiBUXRKsf14aZYQv9KwK/klBjbSORpIUkke0+dsLDN6CeUGb
tC/lK6peKS+5ysWmN8kJcqXBWFH1aIMMeMYTFd8+Ge43VUVf4ukrMugQa7LiAOJv
afA2rUCZe9bAas6CRHB/wzjoS1UsldNEk80pbiDJxmnosTbJAOPuVLvmqIE9o5ma
uvTRN6dVY96VXdLISMNKSHEqMfWvx4XBEyjul0cdA35846QteRVuoEHxLTl97XXG
ZuT0L6Rerz4Q4pmEAGXo3Jh0vC/i6JtB7VycsvbYeq4eplcshrKA7hTLkJXFzrze
0RD6wwzeDPzY8mf5F8/zmY+HkyGwUFkC3QfbEJMqw5av3JgA6P3bT99HztqYQRRV
bX0u1lZF8hOhy13icDlW5Qv2EKRIsK/hszR/4QIqg0rvvrinni+vHFU3RWq77o5I
7cNrrsguSdV+XLI+uhprpkwchxcO13r1KjB8YI0ivIT9eRL3A/Lh1vnkLpCVkOoI
76syCvvsnOhTQ+5z9qx5TP7EZjDJAouIUmYSUEDfyf6TrIncf0kjQ2oGS9bjV6zH
CBq5BamIu12Gd89xRdv10jNPcE3HMBix9/0kj6IXM6FDHK3GK2DY1oyhUkSndZfw
yoHxbW66y15u7Te3PUlTF3B6gMZoWvX78iLsw8G/zqEXnQrR8gCyCtbn9sCw8MIy
4RhkoxkuDOTYWDGb8MBNwQlkBMHRWkrDH7cHY0utHfxvSZs1lJ99LyAZijWsnF+e
XlqiY2jQlbuEQDlvGGiuZ0ByVXWXwF7keDIU3oYcdVJcsxp4A3Kc9213MkK6cW9p
p3S5M29n873A/bBiucZmRj+J356RbGn/J+PN5mINN9Ejro+AgOscPHk+FUuO2OCX
K31mh4jL3c1kzULrZ4O39Pul0BZ1h/Drluip5EkGZ9txAQxe6SnZon9dEks9Mo5Z
aYjBFBqjbnNAqxby5p44TQDbyWWLN8b4F/KUpDRCG0CGuKH8zeTlAvQpSHBP2N+X
RjmpsJKufEM7z4esVoPF4WETzNG7Bvy/Ee2xKeQGLnY4Nw5HJa8c3k5Wqniy3mfs
0hk9ejASqpqfjOaaWbkyY/svPrMkNg80bYn/0+GzWH9LRPlUU6O5BxRoZSeIn87P
JckHmEWfGvoOivXfSKowSseVHDb+SzwLofKRbnd61hhQ1XXWKPDXLexEnK/W2SWW
TWElBv9DJE+plNMvDeQ3awcuY9aGBecv7bkRYJi30E6evn6ocG93HwRWTsPZCe12
MOM+VbILXI+8PyidbZqg0hEDM3xzyqwJosg+YllCfBPjGxiUPct3/5w/h84MLun6
5P5vnIpElNWfQPNUmN/mwb8R04bXeuWGxvMARGHoBlsBLtPfLBvvUYFO5oATYl6S
gnrk8bZ7l4tWncLz1asCkbdmOOlRptXRBIE1Un+P5/RwbrGMtVQz79r96Eten56M
H/iEXTWGz1alK1viEmrq8bX/Wzs4NqJWKdr7a4d7s3f8LBmsh5V14ZSB/8/dbetM
FHfIoLMm8XV9/PN8s0NmcfviLHONvC6kh6mh+hqfb3u3bSwn6bucKNHCKW6ikA9N
YVsvJxbftc0zGWPj35KCWxI9ymTTF1lQDJC9Bj9WsNS/LC7u7C/KhOb1BG5hVRVC
G0RHgDZcHIiVBFbUpZ87VEx8J+y4QSumhGy6zqyy5kvRuq2hyhqWMUNWVMCJITqN
IGoanRKwfwX+ztxXlsiL5T92XA8cm4heGoJC11QWGCus8QbBmEy4hxt2LOIHIcLO
mcsM9CMYyMmai3eAPPCC3RSWt6gs5FRwv3TYmLLjoN3ThaWo91wsPD6zUgnM2HG5
CBl5L+xijj13lu1CRRQYqgJ7v90dDROo6pnDHI53rt0icxC2cq7TKZFTfW95vsWX
427htJJCOSlO4hi5eIEHuK2ySMLUNRXQuvShXsHVme2mParnwvrptIirtoJqoeMt
PICl4Ut+9Fq0+pcS/sXYQtNbFI6admLfO2i5ZUDofmEf4g1ufR9PCfb3Mrp/K+o8
UR1F2OqSAAEEJ88uisPhQaZMmfPZmGxmmiOAsMzawfY/Cx8kOJ8OKKNXnSK2SDD9
DKFdCez7Zon3Vp+8IeS3pEX8dES+tsAKcu9MlywmnQjwvf002MlQweVSlpcaWiEp
CzOX/3NfP6rjL5qsaQeh1hdvwG9EVYFOzkQ64jIqxLOfkyZ3UcNpaO2nUyexAHmD
7ua8pvw2shYyPuwx37xO+nQUZBIeJMyZLPN8kBtSpw6PdXn7PlVPz6YrIvDCIrrT
wlbTByqGhpO+GtEy0FAnWi46l8eGFqufR2UbCvZzL0g/90jD8zU/Hg3drLEFaBSL
ge2OReCMzcGEVWZlfQ1Qrf0uuVqCbsVz9zMHujayGjteGBVoyqqDKztehpYxb5DX
gZNYwjrhVFZTuKhkcnZndrrjpJBezfzbbu0oUR1xZ5OjFt5pBOSyOwk+uS5GudXn
V4D2ckANtzCSa8eKzM3Y2Q67gREmslgXS7Sp4M/yYEQfF9qGrb+ZWbvr5v/HCxcn
RHwxb4nas8KSkiGeJy6rbEQq9UoYRIb0pjSLdNt/oO2gryYjomAalHgamNs7ZjrO
TEX54bJB6erUJKG5N+5+7vWqvttQRyJSt/Ba96MSqF7rOGXO2++rId9bv7x5nrFk
fhYevh7u4xqfIM7ecwtsZ8T1jedy9y8ruRUdod31dRCzwri0sbV+CAwwNgRx15C+
XACKfKemKMEjWGCY6mRJMAmCHIUQ8peOgjJa95uYfWc7KxQ/RXfJDK2uLLZnESYI
vVxvVLxaXqETAbg+ZzlrxDmpI/TaBybgUpzHIA6SAfdzJYiSdbRqLdi5DiRk3Fb0
XHvz1ViBEsJFodQn9mWdVS0qEvYrOLfh42F3ylv9vKNUsc5JPIY2UeBYPDEu5R0Q
hyRe8wwPEbqNvdpZ4s1CFyZHmTo8et7A2U6JhZ3kNwWaJaoElNBDe+s3FmQiInoc
7KLjiLvZDVE/FFy/ruLP+aazCJyHkLpuD00Ee3b2Few/VaYbLVFTr4P/QLytHRnG
EWRDdWxe+KE29+mRGjkfMp/QxsjqJsUo5WU8zH7cjJMIiQJ2zTH4lkPTtnxFgr7h
86uxpdw6TqavW6+mN5lHDO4K/RPl00emk3SMd0bBctKPFdNWUQTpjrxkw0hZFPzM
x0mT1fVGKM79gAc+KasijQgZPWftwtiFG7MehdFECYODfKlPS7zN9HJTKz0DdsCP
j6U1A95W3OthrabFUtbs6kwM/op8jCHP1O18MFi0PWGjfH9vDV4w7/RGqdpUdyxO
ITj5MmF4+sqUzTF8tSoaqO93I4lOf90baBvI9xRPXnBcd9dBTkMTPst5wf/UTYzX
pnrl2VXNHV3uVq2evDWeOHyQJKhYWJx9nOfiao7LbwGrQ/7hV8ktLGMWpeMQfeRr
3YX05kgIEvYf/Xc0YynTPcCe4C4CZiw8ojImHjZSnTZIY+ngWqUWWHFtw8EPUab/
VdLocp0//YmnEwj/lLj+esCavni89dRGxrlIpLQoUlw6mDSes0x44Vi10/XiYqmK
0fwKfifJ55wxHgpvcAgIFxxiOZwtMDOI5JQgL6CVrwTDjYTOEeWXtmhwlOYpWQA0
Eb87EH04SBUme9ndesNh/6mAlVeMtkzU0HDJkZzKGmalecERsTEq47kzc9c9q+yf
p+06+6LuRrQvO/mdGJdzIT3lkFV6i/o9cG2QZkTAGpqTLA46e4HGUuL8BkAs+n4k
zTk4x24IGIszEu222QQxTHPsIL2pt7dbAxBW1ad4JbjqHqhl/EjoVXiN3KbJI8pL
nCKjUiKwSVPundKecdJNDWUZRjLP+Qw0/4juJFfsoAYRXnPiCr1eHoO1GAzh892R
JD5UWuiNklA1KoTsAkR6l4WOp1sqv4HjbA42IScJvXCdI6jYk+yBAdQceGm1YmJH
mDJ3pOitxmja9meH6nxtHxdpSJnQjNTmsiYTe3q0iEpMndCfVgv1ssU8oJzOX/u0
4WFRBu2VSOrRMbfieVomL+9EEXFrTeRTwX+nprtadp8eIZUQtSyxzTR/yjJ8qggG
MLUbhYXEScZ2i6/t/TlZ6/sMMSppnx7wrzVmvzMTa9hJCs/H7QNcMaFdDL5MSXYt
lFm7LcoEjkJz3mj1m7W/BAGJXzp838kke7L0z0CL+IAGfJGAYd6Zgt+OUlN96PAZ
5Cqm/u1dKvU3EOuBgcVDANh53iB2dy3/IINLUU336VKo5pwjzDO7RPLeTG2ksqwz
dtsmGYddZ5gxD5RE4BwAfnYJyslN33prxRrpl/tHx/Kem5pvqG36N4e3IAFZS+C0
FEFj24NHPER7FbuSTMxrE8stcCYClOXW9eMNuFbVj/JKb8sbFzT0VmTKrF8Vhc2I
07crWfk6dWKMrroxebx0kFTuAPMOYBJKa7z8qEW34oJgOTXn09RW9tVEaodq7ds2
xAlJKQf9bcmMZ8SEGHvdLhljd0us5Jdw10Hd9tx4x6qsiFVbLRdUjsbNUboOCwPs
nOo+u1WULZ7sjp8NrLJjqjywIW3jlBjeTGMQfI6glc7o+m3VntYktwAn/pNTt3LJ
AGXfDfW4hrB4Sk7ykYwk28MLZSu/YNMvG0bWYwuZC7qGYsDHqpkjEmq21ImS++d0
4+9e/CHxEIowWuTFH3RhBBiadJ5a+83N/shMGKMmq0sFIHHM2ONWM9CsyhYIVzhQ
xu3kFHYGd+0iDRHq+GPOpgyA60xYqTYAqvshdtxGzJ3VspssTAnDsaLx256IN4td
+41AEcmp/vML8mH6YKUzD9YCmjsVT1hXNbF2YmX31biAITGySlxUQu5BOxv/9ybf
JDa17N9w6jYlIFzJk8vP9MhGJT/NrWhWpNuY0PHnHbT/XrsEYwfzho+4rYGiREI2
2d6SpiNtIInWXPm4fRWgyT6m4ceCclPih1Ot37nj5FLsmAD6WNkfkq/dcjJic5pr
xDv9T1xM6WoFaSbsEFApnriyxXYrXg50C7O27Ny6jyDx4vDDA332gjjUESyF1AZg
2W/U3U5Qt0moTQh2HOMsSVCeWO9X4YYDZE6LbnAdvUteGuYMpq5aDF7rp41SC0/q
nn6EYKPmbdTyE+UkglWsfy+0cMluiQE9zC10ZOKS8+K3GJ9nlx1djlvzzph18rnz
kKt3iOkR9quyEfYrIkT+GXbx3Rg8EqI1Zem/UBPaoYWGLT5AXHJUlI9d4kZ3hULa
ITgZ7sCeJVf7AneG1ehQsSOkr+olB1AVsWNXTgLtRzvy6XPezQW+d/oxJ4Hu4Da9
XszesI3vbpTDaCjQ5YASpDxkWKIWD1bTbM+7BByCceYMBkaGR2x2muzG4kDmTie6
VI3CfbAL7rO74oxJMS+ib/7h0nATnp5TGgZ8WlxZI992ym26XQ/ukfJwopluYa4L
EwOJoA8aZqbLS7mceiVhEyJN+nKl8MljXU4ljLcDMpkhxRcfBnv5WGIBXG+Jvp+E
8fcdp8XQwAvmCxLQBKTxzso+ck7MUBvWMJcq+XtMr20IutwSaUD2E6u/31KUw9Fv
xPhaUimhwsro3Kc3t15aDx4D/IdOM8/yZBKhWBJ288yh9LnlLO7FsaL+MxtPKeD+
w0S3xpXAegSCzmwk1ky/O25yIulvwM09M/WhBwoI4rrkhp4/dQTfbIyIaq56kQ9E
YsnzUni8nAIFzBEnMqe73erK+hPRrcA3BnbVzXfRVjEOXrR7Q3ATsY4cXeQDQ/YU
nUqhFF7DcZDzAvcrWd29gLFA2Bl7hkbxnlmEKiQHivVE2/WjL33no7morRGrCupl
F0/+7Y9WHpCK938VlTZoeFqV2Ah+c/lKgA/PqdpavWDvbu4b4kEox9NoM56yW6bU
qRpHyNt7G1BGufL+tym9pUDJRKbo1hu0rQXpWbC+D1RXiKzfN9j5EoAQ/C+F2ARy
uwxoTAeqBoRR8lIBRP+KmrSPa5xPwXlfXstsB9iQ0nCDM5MgaHXRioDdk7obx4BW
A1G4r36eeQqQkVOfgnarwB0YfQGeiFSSudZlr3WYKiNQma3uN+UPeexh5rs3Ev/L
73jZVAlEd7Anp8Dtj3/MlB2RtxgvP1geEzYO90naW+2hPv+9xoE65r1mhP6+ImaK
5UGbvd5sPPknWtYGTrGIa0LPwLP+8dzqUBm/82rGZ+A8oFSCnxULb//wkcS9zrhG
9akHcwRt6x6fteBMnPC4U/00Y+nKua6OmY7YvtieKoiVadCtg5X8SWeyqUHZIrkD
YHIHS514eTn6ff++TWNVYGln3Cf6BW9TvNIx7tw8V37mYz0YtHy6x+41Kx5HeIK3
15voKsYxFKImPaGtmD6VwBvjZHsv78bv/EQn55i4dqFMQ7n2wpIfHZarFFcuojRz
eIKigJlzom4xhBBkKR19ZIcUHBu2DCZ+ZyaN+1c7XZZZyBrLFWxdx4ElHUbSVUVh
mO7E8luccHSfj40vCNIouLl3GjIjqGpnBsTqQVxDIQ1RxEZYQdcCwMvj/8bmlu9P
GY9Q7lov39yBqdPg4nbNC+Juxm9zoib/9crkq6NZ5MgxLYUdbptUBXESnmfi4ycp
0D9+eeUQiNDLeA+/ue7YYzq3x3cRmogPjD70aeeJaGtUXa2IaabNM273aNuTP1WK
95ugUaTEsOXYKVKHHsrBhVE/QMcYDUFSJ/ZcRdEgplwjp5Ejw3hHoHQwrzqNmyNa
b1iavtz0ZAq1CNyaQSD5RJ16IMAcpjbHBpMnf5SmVi4niNes4QkgbxOP1uBvuLxz
h+5PbmWcTFOeozfJJDCsOnR3kr8m9c3TBP5iV8v0fb9iACaZ35IHT95XytPQrfxH
pNcP3cmSW0vXjAP8dRSihJlr8XS6170+lT80X9OskvsJEwip0QGGHaUh2m4a+Kxr
Nx1TlpOED4LU/JXC1MijscndWSjSBUyLVFD00ngN5T2+NSwHmRVuKdxxsew9GVih
LpJeCqOyf6f7FqQ5IQLxlXq/qaNi4JTtHSe23JktezWQ4XEKxgDpEw6X2mOmqAwy
1+rk5GZ/UAuCFVyl3E5pACgqOP1Ltusx8Zp6A0eyR6Ko6iI1l7sj/qTSSG/k96sb
VyotvbzmS8BnluVP6pzXD/NMRhTH90Ozdc/7iQTyAp/qcOGzm3moxJSJXz8h99xL
buuCXT6d3HzS5AFV1PFF03sklADHcf4sgpbUQ6qS7OkvL0Ug2f6R67hfaDG4GPUH
OY+zXMuYOVgcIA3yxAuM8Ke22GUTFuijaGwewr2c1Zhox8lhd4WQQZSensUmh4ug
w1kekmMCet5wE4bip6esWlZF2fiAl0W+wo8l0KmFO4c7ZloW2ExcFlWjHcm+vAYR
9UKK5i+iE0mnByAD/q2nniRJSE6iKrQiHvsH0TLhjaE8bOsja8pKOmAsTZd3aS2M
wixV/5r/VxGuwn9pp4LcXtgT3sN0GQ/CNcft+u4ZDn933lwfl2CKSxMmx+yMCHuA
IPGol/Xn+v9CWeIb+gbGikb8gydEfcZ8kpeEQr62ZDTSbVOcY0KMWut4euO8Wgz1
GIItcmMZYSp1c/mlFerp22dZtt+Ce0tuNYl0GZLCjTTbLmumb10aaWk6TM51nM0P
FwJHf2hkLjqLK1MSihkbZ2w4zPVM/I76mpGliJIRbuDSILmwPkABFMOvcS48n4qQ
HCBjPgG8JA/GGy/VHumX8q0YIgfAYMfuI1dI8ou5SMWzqM36Y/+CRtY+CQQUICaX
jLxEvcbwc4pBMVBe75e4+Qxgbbrk/Y1TNPwepBNO7CPSJUmdByjjN4boW3VjRInL
df1j/q2amVf3NM3x5hj5VbiacM+e2LG/jctPF/A5Xk+9peZTOhAPO1uHCaAFPDMz
6Q9x4IHmX3khniCg+pyDUZziKGfi91mTnBH7Mj4UCFll+tNgxhffbe3QZtJdVf1Z
ucR7yKgApbM4VKgGWo1HBHZKGCAyLEXcwOZD/ezSMNzJ1yxpQhnnaVtZm4DSF95i
B1kl8bIlXDJTSGNPmh3BQG1jIjEE3jNDS5RF6Lv3dJGwpJjzu6KFsb7ziCpIKjqO
KGgh/ucMr7B2FEbspIg2h3B9G1ermrUQ1AdipU9lC2YVdZs+UeGgoX6vnbG8qY1X
8Xqa/hW81lziWYYk22yca8MkfACnvyllfDCG1pS6i3zj09ISim4HaWx2nC+oITSG
ezxb4FenF5EaoY8Rcfg4PlsxxWCb4W/MTK0nRHrHqV9Rxq634SrwOpliY4zA22rv
XcuG/o4UEgbBxtaFucy4CmEMThpJMVNj3KUPvtRBq7JkfLahf2CqV3WGZCh8VeZk
OPTH3YmFHOu2TEn3LR4mBrNzByvmfZ2OKZ9MnngUvalvodnm7YEUgv0l0y2/eM1f
fyW5o1+RBJWkt1YCmf8iqZ1i81ZLXHxG6Jjuo94mEtt0EcivjyEeeOzGoak857qM
eWcLLOcoavpmqvGnpDHbtUSrATBanELn1EPfPudteumu54EKM54R6J6cENm7fCAm
QfchjDZNCACGDtjRsh0cyufVsesf36uPcP5UPH4pXbzbiak6jhFEta03DIGBdvRf
XNSsjfp7riynZPJUkHB1HAGQqrOK3MjRmCTT5/bIViGtx/9CxEo95s/iCebAoj+h
EepQFWdGSUgHehzRR6zUWfKHdjsdXZAlL29Advp9EY3i9y/fVg2zn/yCOWdnztiA
l7tQIQWqa3WuGNgmbvYs2+Mz5bXFckZzhoBTyeRoinRmMnZMMicQ2Z5HNdiQcCvf
A3XfyKJszYzkVp8yIVJaX9hoxxZLHunLdTf4tXxXggPYS6NovNXADkmAOulCaWlX
7sgwA+peDE+QpCL1r8b9eTTORRrKQQbbg8icp5jRiiayyoZ7a3GgjKF8FbZLnxl8
i2iqaWFOnLznRNWgUltd44cOQUZAiFT2XQwegn1iJifMBqdiOb6j7nfeX8i6gCF5
Qg8yGeau9ZFOibsHQOmFwnAIxCazqCvQLF6fZoQTLu55ji9nfs8iz9YogfzoXY4J
Z45WIm/mRuNNzGP1QHhLXXFsm8wFvgu+8swY7pFxZCf8Y7vz4tUH+jBxUQ0M5Ib1
iZS29+jJkKM5Mt/mCbobCzyDkA9pZVkstj0Sun+0qFIeW0BIJ/d3QcljUtqMJta/
sXR/DCLJ+KBCOS1GtvswPTs9mnDXfZcx7rZh1M6G/Qjlie+Fbn7hyfP6HDIF79pk
P9+1UHcl3+pu8qIaz6aXphA+WB+/BKrEFPl62FXQlAqIM6+EKG2D4y4zjNQhUMcD
fVh1XusWmTybQUwv36KcpWgP4tKeF2i41kvn9N+1tpAvGpYDJblgiGiCK/8szcDc
rBAAf2yfFud7tEjJHuyWYKZr/TMkawRekKZ60lcE4M5TmmiXc571Wfb+i8LbbifY
tpyR3239RrUyWZ2ZnIAFb3+u/pFLolm5Ctx8l7KSQs3QG2z8hUdXnstYgurb/hcg
VzX8OO04Izmv/jW/lGEZ8TZWoXQEwc0gLCFXHa/6tP1H9/JXoyo5ZhNgqHtl3HPe
6BbKBSQBWA/kIwNz7NjqRei8VGfTppBUHPy+9Ss4Ju8Zx6Ir5vP5k1C+zfIs/XrD
gW0Ewp50I5kyVDRp5uAZ9jKldwXZBeXlRYpdsmJU1+JdRW0RkKIlYPFl5Hrkhs8a
goQYUoxTFeMC/jncHqd/kY5+iCdYzCMuDyi3iIzYTAfkiTm4Wa0P1pFyomHiK/l6
6mIoQBDo/SWTfnSTj3kPRg++gkBsk/srWzhFJaNM1LlOEBeVjGPy8tK6mrqAjrDz
JUYiU5ZOr7P4gTOOm9EVPWV4O+BvhpimZ5nSmV6LUIkAjMr000fc7LnkMkl3q0Go
Eq3gdW63Fo98LA03IgAZlhxMULaNSN0P6PGdRy3KaykyvUQ4PymUl7/X9ktTq9Nc
eocoHqKODjIObttUY8jcl9xeK/P1h7RJoHeTJ64zMVR5JDYEhFZqw2CtfFiYY2e7
TIXVhQo5b9g5w08mNJ3yrx75kEJ3qfJU+QcdQU6V73F49omtesHsCjhU3dEzXbvF
gxcP/X++SLakyH0ddDMbuD5jTikfDBsB1D4OYtxZ8264G7/6WwsOglpxmmX3ZjIv
xpP+eBAYs2FrsPqUdDz56Ci13mVLgLF+e6r7lwzf8wKxINkKW7TZJ3cwZU62yZ7x
nkIPTw6k9TyabGh88r+5/5nbXjITgxS+wpnM6R+4L1pR2DPify8j0Y5bri6TTLmc
0TfnTTzINhFLqoGbr4WbQT/71uYIa0A2RVPbIVphdLwgmNvUrJNb/+d9gLDCq/+6
r7mG8LMFW5FBclKsTefJdLvj5EJdlclBxgKMHUi06XA5WIDfMqZ38jvgWYBZIXln
bzI8D4uil+dQc6hRVQV2l/qxt442arFm2xt8zGiu4cmsL9cU3VSrLPlqnK2K6TJ4
TGISOPL7rKq836rvS45kHXmppzzFpQ0QP66Tm7PiVL9nUeYJLFCIKqPQc0QQbQ+p
9arcUsyEh4VgxoIr5W19cy40nems0B1y4iDvoodNDIp9Y+U6/YpAco3sN1UTYgX0
m1huzZQ/hne49rGyaPvgYOd1PKZPmb//4/iSdLXlqLolwtar+frPRtDAO5BRQj0k
jOJ/lOxhzmFX/rUtVZe3q54XbBmlHbZPCT31CWUMbMNGr8XELaIfjLhSNbUDW6RT
WPh9NCRLzuWbXIqS5pouRGO4TvJz73TtK8w68Zp/2ScLiqp+vnP4e45DNSnCgBly
F07PSGCNuE2pEryQ4ocgV8rJeWXZDBhWTwHJ7Ko4KXUuU9bza/gCMeK/TJFLrkj5
ZCuq3NuJd5mNg2ykduDWD5XnE3Jmm2e6FWaMNlhgZJYlLzEy+/MzYVElacxz1uXU
Obij2eRyvBhHtU+H3hw0y/XN7YFm6KTlyXuPzrae9JHAo2e1mdw7n0uJRjimXPpQ
80aCqWZPm4FAJcBmU05bZoDwpNgEku+X+rJJKkth8d83wcOP/pHuQAqH9qOlaZ36
y57iO1cLEnuXD6wq7ERSkj1svbdS0Rd9ZUkr5TZLLglz7fOR9B9VywIouWdGp/qC
nd1f4wkVVwZJWyKRTlxr8ngFZAaHx20VCHZXoZ4yKK58RE/kkXISQS6OOrzkfL1h
Dltv93fZFoPWfBUiUeMQY9pixWTGAcCGdjmCyzg1lxwOC5HCHvuXAwlr4D08xSiq
Ek03jBI1CO1w585pl2+jzFnqE/wQTzjSx83z3hb0tw0OSQG6GGIC7LrX74FinO7K
NopeCI49vysLCLSP0RemUQdi9zp4gzQs420St2YyteV4d/LJcGdODiz58wqf7m/4
r8+oBzw0lP1QNEiKjD1nJRjKAWYla5KC3oPBnCo8L0lyjj5xz9GMbL65KRvqBVBx
t2Ggm8MPeBoxflKK8fBeqpC7GoIMIJ6syyL7ov1Wknpz5rRE/BlgEIXqf3KrN5kt
h6QpWKcm1AaOEKF0ZVwKDQmMksTk0ic5GSoPTu8Q6jagcRzPKCJ0AOzmB/8rD7NZ
8dQfE4L1SNrh5jVPDkOeB/dQRqXPtxOiv0aJ49c8nzWpUfRlnZa16+xYCXRpZFPo
TuTKSQEwCPyA23xDkHKR002otAneD0flEI5LUwffyop//GfblAvcCebQQ5kYOkwE
c3kzGcLDszi2NiZDGeuN1/OS31QIJ+jR5fuYYNgo+oso9dzVvghDtmFwdTaxOPtK
FI8EYm2OKTs0ScYDX8Dh41wjO+wHQOVptdNxHqayfRUmFMn8DCJ/gA7W+Ew/i6NZ
IgIoy4mUh1F3UuxvS8/qRu1P++6ajXmH6R2K9RMkmbjx/xB0aGes5FFIbdtWztyn
okBiL2ed+NWty2jVVnJq5Dtc0L/bJmx+rVasdjEhL7HDkGEQytjNhLUeiLRQBlPM
rzR8SyvAMhFUAPwT+C08awzd7xceI4OfXIVdVZsewcxAGhI8Cu2wucotaD9102x1
LZO60Chq0xfVghH9lHgCiWX7s+0AcL7Iwu1a2I7c9SgGajE4C/az2HRus2cee430
oPIsSdYXsdNqJLMV+finLWgBKtg+iRbQbX5ZTyvwGavrs8XnLwGTDW6t7VroCQUY
ZPqQaq2VpxJGytay2WLb1ce8ABinhjW2Ip0BWhGR/NiYXmWp6g0EIF5RB1lpeeTf
1gpLPI+t1Jf3AEVbZUxEBOynnLApi2Ks9svRV21X8ymfPwAgCcnZJKkXE8iuRe5S
TKgXUN19U6vPMBQUFDZO0Fyv4GIm7XXp/1IKKp+VutO6GG6ooyGNxHfdcoAK23Zc
kyVTB6JG5UEiSseVH4oCg3/ToVpXejUmuYvN7vBIStxet9espFRM8gvXZ13Z/yRg
Mfuz/KqL2NRgPmHIPM1HHe0HPikDnRGjHWLYxI0vwLD8WDFP1w4RGQs8P1Oh5Gyg
puj93r0Iz9DJkL8iW33PseJtlLjJqidb5kIm/dPNEjmxjfE68Ifv4uOT1GePFDHp
vEboOjuEamquzDoJHWXVxfou7wes9HPMuSF1Z3d9x/T635aCvCg0IM7MMLFeMQq4
xmMxqCGVbiBY9CB68AKnVOb/rjJn2hZSx3YVejQLVf57Vflzv2akU9wAxLvqj5iY
gKiBB78EMduE8Hp9+8GI3Dk9PTWVgiOsyoSw6DNH4J9CC8FUCOBEDEoP8wqMIiSs
7QQEA0bDQMqZtLsBk6dEsDU211RpIf84caM+DTZEQCyH9X3fCArbAZMxLa1uAmyE
bFBqXuF2Xjnb8ZyepmzUabIeVSLW4aep8KkSZUg6o2Ck9C6S4c/TCSDfLsGehYXh
VsFuKU8b/tbfVJcuCVKbt1qqhKI+1jq1FgO2tud8XVk+kLSbO+4LKPE6tU3jegw8
BtcfpJhOH68BJk6e3yiFH8vxSo6lciO7aqEdA4Nt8wZsMIaOoJ3UxJ3gWFBc28Ou
vX1cPj98JXqiY5iddrta4yvpJvHDkrhqcuP3atgNTYdZMQ1Dp7CLKcS2Z+pvLxN8
MJpVaI2oKmMSOac4Na8YRKbpLZKSaeUVmN8OUmJPdgXGqDgpxPdg7YbkNcrpi9k0
PI+vpOb3Iyki1+TfNJT/WMswdTjrwsYT6slVmug7rqnjYS/U9ofz7JA2sDqG9wnP
BeverlsRnzpjLy+zLggOJKkbJuMsbV8FJbzwunEwlUCh0xpl4ysxuJAVGF7uUbVC
mMVqqmy8p/6PecJP1MDst48CCPfm+p5n6wi4tr6ra55IrR/slVVjgVuT2p8PvMxH
JujvyUJx9/Zk5JGjwsJa3GolkOlk4/3btyo+9nJO0Q0dP/EpFrWja+aD4/gLTmBE
vtuawiax6ZltB5sP9+c15UMNU2IjGHpLJwHAp2Rhw6SmxYMLjnR4NCr/+MDDIwpw
6eFTuUVOGQ8Otig/LDDOZsV8Wsapd7/s73hOXQunytlxXTEdqjZrJxuxisKiOEdP
F7zjwMFK5Gn4/842Pugw3dGBrfr9jR/y7RR2CVRWmNpzQhSJPRUdrxw8A2ovHD9b
J7aHKSPjk1wbpiaAiB/PtFTe2V2UqV7uwBnxBk+YCyU0rdnTknpjr3IjZMwyXgVX
Wqdac+ol6+z1uTDRh2pA3xjyLD/NW8mqd8lk6VkYGfmNdIYZ2GCxMoPutS/QLyDe
SGZoGRPF0PfUfzQcGJ4bl5iDqkLCSNEDPInN/6jSKYD43bQ0qAu5c/yEddvj02nK
X26gj1Lp0mjB06xbIW4XlRlmHIx7tWPSXh0PIPKotk56MUA5dumIoQC6gTEZvviI
Elp6VQiNrKjSAK4L5Pl/U9V39ahAMn9jGsaUKsa3qCMLqNiSprEnB+H4aWhzOLWo
Etjy3WLyedFGHVjyLZiYsXWn9iT3jxChKN8FD43XyIp1iDAf9fsF8ecwtuUjBPPm
FqdkeL6tpNcFhVQoHtpRrSVo5iXK/SmezaR5F5oz0WMPzR7lAjWbsN27QoePXdgE
+edBG8oSMOfDr5KvsVkWTK4cZewKivFivqmigo14xq8KlCL467SK7Xb3tk3MsQ3j
N8HtuI2l2cA/XY1dsuF3NGkebofpJEyris0UuZTuE8VOcYYGUxld1bKGrpgDIvij
rsdslbh8HG1nMaICmpv7fRJ1IWGO0J95LGrBQtvAvfXI8F5LehWuJzi5e3Fu9eoA
ES7xTPGEUynya03u1YiqxyEfsmcLrAnqXIm3uDhTiNDsj6FlyDHgxeM36e9QkscA
3BEzX4wbLUy/mFYUfyyGPOM+5Qgt+0Pi2SdoQMWK/OtTUwdLzQl0HtR2Q7WsGey2
FQJGmKFR++YQdYy91p26sPlpsH9zcbEknajQJjMdJwKeBsv4aviPQfvGfVI+Q83j
IJzqWwSLwzuh6HPgggCAyNGoxqcsPRTqS8hqKxoZvD/xfIhtwYamDTNkyB/ixaRm
mxZQbJloAXk2aeABtm2nmq9HwtKgnR79R+XmxjacRFYjtawDmXRhvLywxfxJ3sVu
sRcgNrtZq2/TsNH6oS1Qnw0tbfpdOD5T+/wihC0CVfUUY6Mt190ikHE1mfNmEkry
5ZmCdBDdCh3NuUcbHoECRkyp6hAio+sxw4EW0asCpQv2eCRslJE8kcm6VWvquJMa
1v9oPukcLiLJer4v+0eigDZOalY52vMF//TW/0BzokBSxRxo0qtKTdyf00i2fyyR
KC40QmzI8PmuM+9P8l5NjqxcI9iaC75gt1f6yEFXYuq+MkDcxOt72AA/s4cfPK6F
+Z43F/xIC0qH/4NWKEN0TrsBpA7gf0kQRPHxf39FVm/EKVmqLh3JIgXtGHXH6XWC
8sXSbxCGQSAv0Za2v62DInWJhfA0ZnfifHrOIxGKfPj2Ln144+lTMMt4B8syavj3
LO7xFVlQkAXinLlq5I5pNMERDJwBkdklRmvEJgVfBnON321Giy5Iehfpnm/21Ptg
DwA8Wsq4kPwSVtltLSNSBmaaLTnshwG9/1T+ms8AlREgIcj96gnh8TDvqbZ0WxsD
xSJsAuU5iAffbMTe1B9qLNe7aZngmCfZD2DnFfWQ55aZSBDozw91I+g0O6zfT/hI
zjFWis0ao3E0tw0Ws4JHP8NyEMQoxhJgue7qHOhQcVGtUUduLFHoTJmD+rqitNxr
+XoEjKspJDRIV5MsqyQ9VbbnOd2vzMddeX/XDKNlMoR+Wq9oIqdrYXi+0a7oD0iE
hGBMJppEhrbouGPyhQTFm/aNy+0gAJnVB9dFJKZ/3izLyjmwdi+xaRD7v6UFj4+p
bsQpa4cOigQq8QbqXmyTVFLQSjznO/c3tEZ0eNquxnCoaNBTZ96xrTbrcFdf6Yzp
8PbeeRv2rPMa1mjWUltK/yMB1PFsUKvlbujKY5Hg0U8FtCudZO4TckuOFCU662wf
gVwjHzoV/WiZjnEMyOtr7ceeff5Ng09gy6xIo7aGv2wwNJsH3/g81U2pIPukeMkj
j2LOoVrNsgYJZ8ByZnGrSBXBEwoDTuQVBVi7YC+JOZF3+Lmh40YecJ8ZqiAFUdjP
ioaNDB0Cr9cYlbrTbvJyJQuDSwUJeJtHb5Ydgcp7Wph5bG+4DMNE8jTqVHu9mCiS
oJH6bq2TPaiUnVfSIYu/XCmS+lJuMrR8Q1B5f9ILphF+MwmL1m8EDmnS+Qzd2C/H
Jh6Cmbcu7oBvujucTDTqsHJNtqjUkp84JP1LL+qEFBZVbB9A7pIahvE46Ii6f0f3
jM53VhjYPjDN6E12I4xO9OqZ2We70FFyNhmG7mhwvPzcMOKIV0ZhpiqED3C4Dlsd
h+XFcpzT/bIBDiTnHrI5XfoSC2A6jCROKB3dnUjuz5CCEXzfU28Wv2YnWCm8X2Yp
OZUdJ9Qff9DZhqfA8dLGOAEgSuVjkWz3x47csOXOZn5cGO780ETc2ks4AFY0a0p6
GHQqx27nYT6AADNXRgmrAkEKJzrbRutrVpcoj38O3xqzZ/AGwhBm8Zu3r+VaCq5E
mvcDrsVBNluVYxBZtC9L2Ook8kxtFl8b6igo+jvVCiMSeG8GU/A4eTAzIaOXm81H
B8/JzkJ6ONiloBEH/QrzUld1SCTAvvQqGg9grHicNcVeL7nIXbFQjvycByyoWS/j
6IMrWf3AFunD2ztMccRJm46Qt/q4+ZHfEEX45xZXQHRvJCfxKUI+9I7xGhpM8z+I
Yj+QfPMjdLb7jozzLVqlsI+yU/pnGEqhep8Y/TMxF+Uu17Wuc2+0c59U+EVQo93W
kb1RIQylayf9nh3umZ9QdXSI2FhVVGnqCIOzYAkIAKVGsJTrBmnLQk5eMYd0BFmm
yussNR/aR4yg6CEMl43Eu8GN5/VdypziDcozbnZhaVKyw2CM8XD0zn3vwanLyfvk
Hltnzbw6PjwaOlsqB6IojMWv1jbetWItxmM6wgp8vh1J8Gx0mdpyZIxybfDUn77a
sAVL/TWLgkBvUVqrxmUTHW/QMvKXl7blEmvpaaIlSX9pwHLUEz2nSVuHeYpg4xOV
8qNkRqXcAPoURtZ00i54CfLCNkGXolzyZMhpCDVct6WGtVYRU1NROGZOpL7ySKJ7
05WHMTnnd2velYu56m6KeiO+A3EeMG6kxzZQvvtIdZdVKi5wsuV1S0wMri3XPKpe
1WbWwB/1znKf9Dor8hlParL7QvH2d2tYibvGfX/yaS5JMFyXlepi/3wx8XqkPQvQ
QTbT5kgPE8c6f6OTj9Y81j1SR1PJUYcXc2c47/LRk6R2/TRw1WhIhEc0JpseFyjv
FvekAI80c8o0vRuHgrT0bseEcNMY5lfcLHg7XuW8RgDP4EaKjKht/A2kW+w2ICZR
m9/5EREzg9U7rRdUIZxVNW6DxLGHd6nh19zELFA1VmkSwu9Iz8TmPdXf62TOGccR
xD1PZqEgZ/yOOVAprUYfj7gylNBwqwibql9IQWiRboDocNmzxGbhOtCQ4OgmPQlD
JqJQ4FN9LHmvbVZ9YXx7H5/KqTCFcEi9hRLRMMsWOqutQXab6xOlGjz9AQJZM8kc
qhIK51Sl1KRqPMqrFTpradGzQZk7xe0PAGF87zfJq9zvVe/eAA5eV7lbBR4tpoLP
L9ODtBUU+hi9F4xdNAcGSQu9oeINHwg+Efekbx6TEsoEAbjilMWTmX6li6DJEQtZ
iT91Mpf2qhUL7xB+s+OVoJuInQBUMQiNPzF547sfvyWwVghTGb1dHaAiClCh1mTp
sk69OYmqqeR/BR6lIxRW1IQSNmImp8f52gDStL/n3V3WyXJ+aK2dAtGIIiKOef9/
gEAspr+wnqL52986uAnNkZf2kSqY8oy6uta06XmVKeIm0sbQncaHGKb1/iFcUHeB
QmHGFwznSsX/u9wum+7JHssL4CEyTWIf/8SJN171mlfsWv/ze3pu2bBpVWy60ga5
+3lAuSQIgwdMvRG9kMKWSzkuCX96bqNh3hBQGVOf0NoRyacYcVZQVqTMY7emox10
eurJl2dIIxLzt7foHIqEUFvCULnJ8Ra9AUONlaV+S4BFr53SV1UESKJQLgiUtOUO
9VIsYRaxLrVDKOBg/i1YEmgHEnfnXd2sD5x3+PpfdSUs/Q5teEjRcMpT2Isyv6ex
Zs71oqNYSobHHv5pMZe0mH4ZQexhL5i2uiUt+wRVsp1E+FDu9eDSUzoq39dnO4Tk
Xg29VqASMm47+HdVucIHiCbKpSlWv0WRbk61d7Hjv1QnGZSOLLxUNgy0xSsIGOM1
77RvfSbiOR5cOatETBk53phzAYkEtTxquYWQfRvuSDJ9HZ3pnxk0zgxD12DZggMb
RL4a9vaba1Zya6VXF/3yXN1j3Z5dpTvCXFd5sJbK9FKtyyPkyqgn13JAnbIZOL8E
HtqAgBDa897b7GqPKWtfQITUEbM5WOF74uwgbKu9VUAs2In2JNO1PSVFLrEAwfXN
LXnw/D/S6x/Pif5sjcNmcY7iAJL8p6kuvji77hwAROl/UlhHccIiT0BWlMzr47/3
KyYWz1ibbdaAC9Fy6B1Wx0f8qWRjKJQIPEfGR97kd5euABNYeYsWneDESxJEe2bl
BPqDw6uhmozDroVM/QOklPShZCeM/QL9rUBP3baMwOErXdfc/MP2FQJgs+jqbuLV
F/Ru0MXeeOp27CuaHSoklPlWYZlPzz34rLBU2M6J9M0RgxN1LfKQ643ISKXUxwMr
uqXspigpVQCi5j4JCax85sb3UqwP3xVYTFzRCDID/ErRubjhj1IsF1ITw9xbcp+O
M1ERAe9YnOGmX6tPaZLdSWsbleYc4GWbvQi1nEtTtlHiOcqPv1ZKvp9mZEF7Y8fK
ftiPVL4q8a2XpLylARu8iZpp6z9HMef9u60reIGizrRZIaIHuXUiNYeXt6KNmr0Z
XlmUCI6coAa15wZfDazqJ2KBVh5/hTOyUw0gh2Aak9HIbpZSqSMUpUvup0NOCdXq
CLsm+dgJ6fR00dSxGmXZvhYGuNt70/x8NnxYu34+7SJ3aITeJFK351y52TGJdMc5
Vyg2qnIRhBbJ1NUr2KXRa3LlDYt7y1zxNzD+H595NYktoZQGApxvhqH7S3tGUNsv
o9lNjHqSTRedZFyr/cC96EhV+TsfXOW5lnvu6fsc9raPTbot1x3/CCfIP+HvKu4Y
ISNdsu0CMqOSf8CIhnyDVlNGncPHh5S1e9+5Z3MjLJr/DcQdbY2LD+2cnEUzOa4U
NeovFzNjfT+rHnqJ+pJerP1GIdIZYujb0TvrH4/ZMMY+DGz9ViUAeOE6+WchChcu
DotqzTfsFPz7exD2OdPkPf4SXww78KrNrcjF1MjxndGUAyeYH30mn790xfJsELU/
TLe+q17Hcp/Ex7Qq4yr3zvzXMFHCjO/u4SBYAG/t68ef2mouvmrxy9vtIVrQbKLw
TufOrS+z362hcNMaCsrQnG5gfUbE5dAbJKe/lruONKZBOeQKZJbpJCR58bC4V8zF
duNGOaz8bsEKC3UWOeVip+oY4kaxgEqMwtgInT0BpYpfopKNz7atrclY5OPRN/Mv
cuPN1ukf1a/Y3PVlhWrUW2iMnIbIYI3B+wY4gi5veqz65nuxjzjPhIaRSLWh3E13
CAnAwUIN9CHVG5Urhs9eeeupyqM1Uob5qM9/bRTILp7p3oRwloJp8viRClMuVuIV
I+shWHww5hvDr9DU+PzuIuDRtlL5PSkUAk6+9FEq3pFPIj8K7Wx1V8pbFdw8pk+5
ZwyQ7WEgBjoGeg13BCTxQKFySwYfVGINyZrEs+/QWRyc+tiQdjvkeSPed9eEZoIU
UNKYVwR9t/k+8AFJfE+mzr4aq8n50fjoASnjWcLtRuDPGULf6/SiSVxb5lE4Fa1E
Th55Oq5YtYGxf/Q8TzbM6m5gNbjhT9TToLrAxKWnBqvzH1TItpT7VYVxg1n6z5mF
IJxi1AfnwR5zN2oXO4vr1TISMANBHS0MQbzcbW0INTcHBDBGIJI1f3rRV9m7Lsc8
anu2/ZhCDBjL1FMd2jKwWEeSLTyUj6VjDwtFzWTcOrcSJo5PGYp5uIQ8HXIuZA2U
vjt9p4L2IbyCG2cMxua+ZuaK7iSkZgk8KUCuKdl74pheePX+dMGZH6Z0ukDv8TKG
tT/WuLmVdjlS2aQCacNKLVvVI0iR9okI4SzSbL5jMAiXc7AsR7oYDmgUivAI8HSy
03EUsSwI7rm/x33seP9ktpurlmU3XOjBzg6xYsHDSZtRhrsWzW2xmmHKF+tGvaSJ
osp1nKUYK/gz+Vx1S31pbJzQEWlJsxA+RKIuqem2r1ySU4/fSqnAqGsAFAz+meRi
bGRrHDevMnfxiK5qHeGps1DDZq6jMuEuM5B2/dtQY6TbsAzq5nSgVSFPuzf/PLtb
4IzcGqB4E0hrRq6abuDSTu/6Sf8Fgrj2zVWhqUNTCxs7i2Pa3Y2nQOsjJJSd40Jm
pfxztqIljzSI2r908vL88hvg1U21m2rv/5fGIO2KDz5zJSjH5WRbCWa5A7rySC4g
tgo2cZVXZy44z3LUguf1964ZS3sj9/pjt4+6ILwoJ8wogMgj5nJ0tyol5iB3/jfY
R6lCtZUGbPWRhR5D74Prb5iop4/dwvo3urcaAHCUJMR7RTCjgm61S5GYksw3L5Yu
t9U/Z4viNu9e7Bie9UWfKl+tUgeyibfyz1fWhFZfZVcGWM5vmii0FFOtVi0d/nyF
zoO1PbFFRWzrYLvhiaA76BSsaqt8qwH8xC1cOXb5efjyI2pNKEJT9jq/CvrNY3P2
0/styOlp59u65tf1YYPMaA3MekRhW9YYGjuMqmU3makWTm+VVY02RKY4gvsuIbO7
wqU4s/zLIyfkKTFnKy7xNqPIaAGZB7En+EQ2m6ouao2ra5N8Fv0jVL2ABLsTFu7l
2SDoyshwGQPzNISC+2IQ587SkiJsPkOeau47KcsbhBPa0eKlcgf8O9eo6UmHV8HG
ST3WPxWP8gcVClDrdUaAPshQ1byxcgt6CgqbdWgx4HWcaxs469CzooeBKsff4hO/
khC8yo/ta/UDk1OamhitfDIsVGF+MFc/83DEtsHcsW93pKI94biqhs1qHt9/EHnL
Aj7bvOCxM3vkyMCZKyf3G7nC8n5xbxAHfCp2QA1KkGFesKkYPkYa/9OZDqRUpjoF
WX+7RJ9obEWOn9tehH24sTl23jgt1lXvwKJFqdnxYBHNbLinaSbt75o0ox5BTEtz
zslQ3GBxBTmPdge7kSfib+76Z2zX/2aXXM4pxzMaJPLmmLVrodtyCEB7J/shXo+y
Bwhjn3X7n8XDTtzePWl1N7a4lNrFz8o/0e64aH1EcR1AfAx165Azic8cja20Ycga
S5F8gPNbPnFnlqgB2IWkKEq2LZDPHzU995+DdnJnAOhpGl0TG9jS/dyzWNhbI2/i
05BTGUw0Jr0VecIVhY/W8ZYyskQRBLUUsJbCWLf7kbZkA1wlGk1A1AVUk2LvgXiR
VRleoGUzqxFAeWhD2I2VpDtdH2ZkxTwZzDyWm3DFscH7qYgsz0Sh1h6CdY0Q+ZhF
DY8amt56bRxAMrFaDSsLaf1KjIE6ZbCNyOoCQhXWDjchmhrqDugaNBePSEcgVZSQ
JBqAGy6Vs/jlq+gHkJ0YjsU8enr5xxvKcQwVPOUK0LxXOBoiguYs9HLFaabzJgzX
OQW0gbNncQreJ65+k56zteKO2CF322Ow7cROfbWn9kH7NKgCHCzpjFyMTa0Sp9a5
8vMbds0fn43qT0x+xZ7TZk+XBgjf1ENz6XTWqW0+ZBGQxJu/QPzTdEi4aodSKGOo
iFqI/HcR2XdrbGWciKIC/NL8x53rZdj8Et9dNMR1/C/JNl5D/lrWP3DF14G4LIvG
DU0QYBoaDBJkk5lGJLq6W+cOOCMGARgIr9VHEzJ0MmrYcSN/KvUvBXozJiwPkfUC
70UGWBpEEupL8lzOu4Xl++L1Bo0LSlCRAkp5Ckfmc1Ol6Sk/qIIjCqPlhS6lhqrM
GnLo2DOIiHD9HwhUQMzATPm6uNp42dWybOcVHWAuG4GEA7UVGVUL53sSzXTp3b+/
uB4PlyvfNUesI7LC1l/V6q3VsqFEpv4pAZFd0HbyNvhA3Yz6NVusziXHWu80ilFH
sDgKd0XoDDwm7T6c/fBLfVEiRYqTt7vQRHjDQ9PwPKe6aS8Hu541XYlqpzkhdIAn
nFRwWUyFKJswmsmVaa0g8zdiLCpBJhPkf88uMQOaGpwdbq3jw/u3YKMtd8T2IHmm
pRZlbqN9uZXFoOupEQZyD/9bd0fUNSfCFfhA/5BVEWSWd9ipooqERXcGC4zX+odc
4mpKzsk6cOR6tA65XEb4Hh0ObIl8csqaVCK9eazf2HBvKqBdhFvkQKmnXPw+zbnA
2jyFZltFqKWY4RguvaA6reyE6cNpjBMkhUrV35kEp5FzQc3srbG4q5+Y54Ai9Tol
FX0X68pfd+zfENBxiwunMHk1K4BaEA5RJyAz1Jr7tW+HaKxvRMt+yZee6RGZfWti
zPTBhgRQ0nrF4lS1I8/7L5le5m1r6k/EuyDhNl1kA5ylbo6uISO3GsYgc9gDU+4T
h/ilXUhR7GpKn/btphttRQnNq2yg0Zebqliw+QHApkKzdrU+lLBbdgOlNA6dB3Fv
3Ix0KeWWN8g1f0ALbV6FbWAK68G+Hy8GXfFA4S2GU30FSJ+Op6gNCY8qCThwgfX9
iPGe15cSOGYEK8ce16l3G1oNK6XTmbu3Y0PHtYHK0sNBq6kPWzn3xd9FfrUdzzgl
woHtOBGD1FRPBrAYmwQR6Nl5YmThsct/vbyIs5F0zKdJVa/TWbA+mhI2nwfayNoN
wZKOury+RqERPsCz2F5nD20UshPWTHLSUS0Kfeg/lKFn8uFhKDidxHPSvHcVOHNm
qAlGH9DXwS+2O1jKqZ20HbWzwPedOKSCsahOXxBFZQxCVkd3qhBaqPYZGHph1+Pi
YeShGz3DjHYbp0eYU9eD+q6JsVEAUed9JaG6C7E18QYdQbx98+0CEgZgE9Ec+0Qg
pERxxuyh8G/x3Hn+fqIddNDEDJ8+/MiFIJJVWO8rflCzhSp22Yf9eEdvh9TkrfgH
ctw1sN3atf2Wl5rrv0IolMTBua6bFe7Bi/iTNyQgFrd0dSWUhibVm+RF/pE/txIn
piT56JrnwTbTN7W5uA0SbHgWGU6GUC9YTeDCgVdg2+AnT2KhIV9tliMY9CYkLBYf
8EmbRg+xZq5WP0Ucfu9P87GPGIO5h/YRxVQr2unZ2Q2ojnDXjLP2ARN2fGXqxFnz
cU5dB7hzzQQIBfV7YtsPhMUYGeY8oRSCiM63TkoVc5SC0L9VYtBcaxWWfupHEys7
7EaKam+4gqE2ps/8VGE34aTub77vBrXw4sJjAIelB6qlbs3kw8BCQUXUMTKK7/78
LaaMNivp1Lo2C2fqDRVWwK53ejhOtn/VYJP0RjOrpdzPm7wnIbvgbeJlumnXcPwq
fjMCoOV/Ch7QKFl1ulNGpyPUtKZPy8KJ38V+ZfLAqjSlmVWOR9mH21zvN3CKgY6l
PRpg0LrXjSNf4UVl2xQ+une7Gyqwt6NaYx1O2tF65lccopBHoJ1vH+DMtjIwgVWj
XFKzVjoTw2tAYjNax8lNg5N4L7YIE6753cUcBp8xKykrh+gc89bK+2zzeGgcrR+9
sp8L0N7UbNivL7hH3ne+cFSGDUxCz7iyTXAztSVkMIMuxq76GhtvV2uKjN+2yF/I
0flo57A97wVv3MOXUJ0t+4zsaJbpcuT5dfmKTCF8c1XFf3+IH5otCujkF/ffC7nk
SPKUFygKrLa/fB3Sg1MkzyqfUUFTBx3nCl+5QZCYV9soM8aXt6iam+Lu+jwjBRuZ
NxN3xgGE0oE/a6CjghJCTZy0eEJFTUPx3Qg9MzajBuUa+jJX8IMpsCapYZzkVds8
bW7HGRWDtxCA38UWPcjC8XdafR64RdL4EjuxXCFy399XOxGxbyHJB6YqDZ82jhpd
F2jtC0Kmn9Oj9ACB16WpMvKBMeR/haiy93obiCQvXNR7Mh4hklzP0XyjRgD8rI49
c5KFFosMW5yvqHBYLJh12swvrZR1lgtHAdL82s0n+nE7V5tUWXBRI3JtQe+Qf0g4
CaSoPAlGO6cbG7hX3bgXEMCGXhmNoBgM+ZSEd+Puvi3n/TjQ6P8k/WEFwVk4f1Sr
owQ6PKPZF7btAOg8tVFrvsG9X9MQtTUtJl1vemci3mBqw2cQJMr54tQEOCxL/1G+
gOnQPAtKszZuJlKO7df6yLhQedRjkWdFLSEcCiN2kcMq3cFosvIGxs26jZxgP/dz
E4RGu4DOUnoiAW61f/U02tjXFTY27OnhBmarGzDOzBaPaVy1HtOLYdHJy2rX36zc
pcNm6gZGmWm2xKvW0wGDdqK2cch0+zE1rM3tiIN183LEFff/qFI2MVCh+SA0SY2y
x7twGttIgfjpuOZrxmidZE5A2y5T1qEEMxmhs/o+UiPnDiDBiSCiBjt+dIwEhIjx
jOkGRxcD1dccSwsLfKc9Ao4V1QEoFxVZg5nMvS7HtSYH0EUCv3XMn7AjCpADSgSJ
Gr7Y/Wjt2g1QBg+8Kg9FAP+SuMAGV3+1Eqh2B5NU/ewgpyLM6hu2ZnVb0rgmm6Gs
oH0TTYLJ5bIyJFEiSYiRaSK0fiA8+vfsjerDD8F+If6CbyfdeKGftzHHRK+GGuPu
6zBY51vwWXsevLbSAMdWdy7hYFER/GP3Xie1weGgGxi13TXJv5VRdoUJNbkvFvnN
zs/dO1LS1A162krJRyTYs2b88ovmUCBk69Z7oz1e59oSXydzGI5S97I7NRSLb9Ug
R76LynKRuJSFKt0BPgXjWCQDIfpDjXtvJFYNoa7dWUDroCjzB0N35Dnk3FGAtR9x
o0H1/WsiVAne5S8KdVmPhfZYZwSJ7RcEjPgPA0AWowHO/hNH4UYSXPcR5EpDj1uv
G/5cvids3MfMgm5Wv8vNRFtjzhhfBRFPqmZzVB1+lQMwUNlvbPeHQJv41CdPdh+P
GuXvNYM9lPmC0kq2KuldQnPd3045SfweqPPcONl4ZvT+PamJ+9rWB4t0X3HG+ajM
J8h6Bvr64UD8sv2tfvXWCMfQCE70r9kKWf9o3XA72aDeHBKv29l4/KH16Av86Dyi
iOYuFSfBMVU3PALkw5bsU5BKOhnGmeej5Y7EtOYgtEb7ta+O+Kd/4QmFzaSvZ7eU
1nLdMYm2YTnSnaYqakepKR9JDLsaQsb/AA3lsO+0wclLhDifUlNonxOVKqsNsUSO
OAaZdeVEH/0BZ2A2Wy7XF+M4kZhlwBbVtBmu2H6z3Gqbl3ZweRJOqWB9kyBT7lrU
Z592+xHTP8UUV70QuvydI4QPuFxdz0dhHvgi/ep7k0L0smHkWGWde/OFMe9BMd5t
DozEfMcLu3o6oFHW4mXW7wRyvo1FlFsEJGE3FImnUXWGptxlAhqlGCXvi4mmE/DN
7mcuWzK6f/XWTgQ1SSvDRn/l0FoVlGAOFByrppy1tNjTMIfvMbvVGO4gvXBbgG0f
NZZGtmWqIXLjjVLyxFlG1xmjYLdAn2zm9ftv0ja9nxynCFddN+2Aih6tA2XV3buI
TJIk/Elo2XPnQ2HiPf4W4RS5YSTgN3Ph9ueAQOfU+QACOB7aWoG7gWD+WBF3ceYp
LvbPX8/MU5LlJk/6F+Ffhd0hjlBC7oSZTbJUs9cTIan70QyXbIcOppQvwUuFNjRN
ED/ITQuF2ZlQiKlNLDy/iSiF0ss9/8AzAiaD5dzFcd9OJ7K3kgZ/d8HeQefBDkml
VsZJB2XQCa6SCPL/3UNAFN/ym/4MaAYwRh5/EI6If8Jn+XJn9BrJbq7mAvuqfaKm
Ss6hZ74ybk5+Gi35xBycM/kqz0O9myNL6ChFESzwVpMfzm7VI2IOWq5wFN9a35b7
Y4EpDEXYSA/ESNmnLdQJxqHARiNO5uLijKLfmut085OE1EIk4+1YW6peMWxEq3Oy
P8q2OqP8JcmD70XsrvADJ6BjpND1ZHzfmn6lC6JydMyRzai09Zfb0go8BW47mfYJ
WVq9ulSQ1r96KJvCM53cDnR2F/8i2MmwdLUFXgVB0wdGcSNsTjuLRa9E7YxGXjXm
LZSquyn1p0BEIOUiNu8IdICDZ7O5VEE85/27MuDqEXN4DcJmT7FjYDBYF6lqJ0yh
mjliAe8ebfuuhspSCcCmDTC7knNuNj3iSUSyBMLD4Khm+hQIKjsuTRyjW5A7aemz
0AulPutJtBvW/mdQYDZWHBJtcNzVwfcPuWxKPgDqfo6iHVjw8CfqA1sRmGsKREuY
uL2K1lYd/wpMdboKHAaPxTZthqMXwOKngXdadD1rxkVPesxOuJCyJaoBAsD+Eg+I
lHKGzRyUl1cTBZjFxM8QyltPuc6gQHAKyDDawEUC2l9qTdn15pn30K+C41aISf0h
vWNJ563y3wnvRuBUfZj2GdkOQRdH7qaIrCHB3CuiuE1SUAm/RDGVsWdzl/Mkhd/E
sMRzxOu6lsyWc+5v8QT5xVqkhsUFUWBHq+NZQcFWXEiyAaPC2SUifhtPgAfm3Ghf
SAB+Y1AM0W0kx0pbGxRiDhj/GNKqYvX2nkJ366s/1dexmPqdvkH0uIfVLaMYLMXA
VwfIb1Nuh8/HRC6TX9+iVxZq+A/PYv75JMTOVkMx61zY4BwwWDUL7N20d3Rr6qUy
5+xvw6e8O68rPNI4fnND5hWZiFWjB3wETZjA+Mcwx7L1h5N7189cIM1vErrCnnUP
n7Wru0AdNnjzF9VOL0XKRGltxzUznTYIAeQKDnnsDMkg8RS2BjDc4fyhrYUd5ZMb
05A8eDEd2CqU9QMHFpET8BnXkhUm5Hy5Ibs58pAx4bJGpmymVoU11YKA6Y1JyU3w
GDvHWRsgxFqMu55tkhz3vmkyMWWyAKpZAelUFbSgQ3E5TPW+KhCq8E9iUqHo3D3x
9Ez2GA541IR9/EPqpeS5AAWJD2Lxqo4EoDHYrmryTVIdifcyFCxPSLFOgUePnnSQ
h/lkzrUQJkvWbj1hXIEp/xh/zF1Kd46Iokob+CJz1tST9sgFsgf2sZKtSqX0iOhX
awwjvLJEhKrqZYsGZBDV/IOfMuRigYV1FnyrD/nb6JyGkxbxx4U9xjnkriSZ7dUD
xbNWsSi6w4X0wXL6iV99gmPNh9FkueQLV5mxbicWo+5SYPe0nMyyJoNhpBGM04KP
vGOFIdHFlDeXpBtuO7OZwiOyiWMdidCMAxZ+CxpPDkO50rlJ1BblmwWK1Bt1KWfy
2KkemIsB3c/nMftUSavvvprrgsTJgFXCkvFqa7N2tJK2tdgLKJbUxaAAYZ9EICiI
XGSVXiSTnMGNHrAQBS5Um09I8wD1nosumgtAVfqDsY7vv6VORLhmdm+uN0Za68ZZ
tf3y6wvAxI4/sH1+28dnBeAYecwLiBkZ6eQvUzPlGFZiiw0Gr/6IxJUgv/bR5Fuy
rPNYmcy17FK1cqtYUCMLnY7hYz7FRrCbgsHogPgurpgX0zu78gxJpZY4hyCP8oas
aR52bRpAJkCRl8w9VZWu5woZRxCLRgTzrAtIouK5JHRF9FyaxpVpb/s11LAe9chw
VkfcFz8i4CvbliJKVKY+VmoDz/Z8cqj0R3+lfJlz2pKO6VUG5bI4IbXVqs2MCkJY
nsurd+iIWVm87EfnC9T0M2HMzKGfB5SEB+f7zrIUy0Y189eM8GAvhXbyOKICKrjI
iM+omIvISqvIAKDa7F+ac5piMms2f4Kdfmd/kZKXkeJyi7/uEFzB1K0lDo1Nvr8W
LGOOqQs2+wvDak/ielz6q71UuEsbTeXKjNlVnfHOYlbUMGanQQpvPmmr7rAexYeP
kR7rflIQRI1+0uf6SSCjJ7hHaDQZtx7yW8y92gUMdC5FuJ4nXSmkK+utv4aJ66JB
6YANIvM//GsIB+7ducLkFXDzHvWq62OAgFtRqtx0KEG2pjGOFt+Lwre6FYDRVWmC
nMC279AXGSI4IzTbVIVy2xgTVR/w9cHH0wT01iE5DxZUb9r3Dr5VVXewLWFpYJT1
u8ZSuTbVJ2iggJ81dZRofZFMzLb9M/rX5mBcvqS3sIqoJiNd23MYelbvAIvGSXeE
NTLFJx5P7qWeGGRi39ZhTpUa78nIF/1dQsm8R/DtTC8IMVohpSYfG+VNz1EN+wmv
YqdEYUZILHUHyQbX9KdgBhNOyMQBlmBmDy1guaIkSW2IBcNoAob0jVo4MimAJ8ER
H7yBO81e6guI06rbcIoZqVOEI2IVCl2opm1zgOaa3fd//Fl81igXt0XH9nFZeTmk
4aW8poIDy77QJVN42swhKJguw5Q5dQMOVcdBwwiIcHNvk6E4xYa/fDCnW6cvVC7d
CLLuMo2a2AENAfryAuGmM1tuv3As0fFvztIrNXAbYMo28dcD1P2UcsZXd7twvFmN
908khMHc+ESh5iKD91DS0brsFSOC9N5gAKQEyemL3KgGY4uQWhITz20HOI2TFsO4
Cv+Qy1nhoTUbV8r37yF5TNHRqKcLb+S/CgeVNyNszlLiacUU9JET62zpAKSnS57t
1nZRcgz+bw8B1CX53/cx5Mu8VDxgHdPpemjMauDW2izctWKPiwEHVmncow0ETTrn
V8iPWknzYrQ9fj+twJOqtKizLoI79KOPqxLd4vXmvvOl5aRJxqmFg1qbCm5Oq7X9
QkmxHW+WrEDHov8xM4X2xwIcs+/LY6f/R14q1WdnRi0ReyG3TnLAh7ikEBECI5VT
Zobdq9K3g8cR67pp5e97JAmmA5cgtc7/pAVeBCKBBf4d1PDGsn5fT+MCxgCrqhjj
8/f33v3d69wOMDulHEcbpQqDmOYS8uWxFWRPyjI9XHzVwhLpGWq3sjnUCrgVUG89
3PBe3ttQET2oxJhqoiNZNpQyWw+vql+7q1JYqv/a6KRUMtpdNwiyuX5TAR0InMOe
+GkdzVPySzTEfMaraj6KsUJ21a5SEhDL9RFZ96nv/+SXtmYwTtuhbxuB2nucjE2I
+odHnZ3SQXnmzyrCha45dPixFkQcIkUDjIIlHqha0wIfUoq+iodxkJiC3YIWiUNG
jUaI2IIoDJzWF3bIv24a7/VQfKWup5n4UJPp8PO78/o78YmwXkiBbnBh1FQDvmmZ
DTy48+2vnwIAAPCodv0TXyzTj5zxjTuAklyXKoIHjs3nDRdgUw3a7qIHFgYVgS3q
/6wqyhwZzb8QGt0qziqP580gGwODZrpiaIOYXoa1tFODAh8Md4yXCJ2iodqqFPBH
tgURYdU9xgPvW54EpNSrgGrma5CNOXknAZ+iuQboKBwSiKGgranG+DRqZ0uZLCX1
Yk+vNA6Zu5c1wBhBRyKhoURP34r5hc9QwlijAHZp3E0jysS67JzfEPj5vdq3v0zT
YJxkDHDtsgrbD+W9Uab4vrLJoSIYpm6lbZfDfUK1TvgDzy315fAwV62q1HDcaFJE
cVP0GzaSEpiPvOiHWs9ztT3BOXskWvRar11+tya/B1wyuverYSY0moEIzAypIaFE
Qyet2W6WzXwPr9NgrA9hBKs2d5ICnKZBbThIWSwny/W4GJmFW9xXdbE6+bA9VWCT
xG3Pqps7Ys7ODcVMlnBjLaZc971z9Bs0tC64MPgOS67+UbEbnWO3EWi67La7nbml
YdDH5gbhFhkRMTSLaq+MSStWFdlOfi+SmhWyaXEiI/pQoH5LqK7d7NDaEHqMTdLk
1fOV4rf4CdIms9lSu/yGULFXKF5yBaUht8/xp29nOj0Tvf//mgm22dHkwpJm3hlz
YRXzSDNgOA3OzmlY6/ghHz5ZdjVEglvuQF6oFQGAA747CA0x2jgU70NxRcvMTCb9
AZ7wS1UH9FNvnm9SOLg+ZOa2Bn6ifIEpmT1mndpXT82Me5nf/uwEcPgxc00btko8
lU00vCJ2b9QlEP7X2su4ta7mpcXBtgALeZO6cEulCxoz8JbcsCPC1BJDMx4Cfy/g
rzPEtch/plqKPcVWK/LEUvpElTrVlRDJIggMBd4/7AxPpwY28/wtm9DQuiOiuIKw
4j3NfTNPR+vkknE9Sv1bxL6TA+pYDS37GQwQRNWN2ToyCCtU1ATTuIxbyPYzl0ui
mWmJGWuQmYd+GbafWjg2X+kctBAQud6d/nvRsteKdtdtW//CYsxoFZiFs+4jysEP
fUGBGSCAECaG+bprHypDkERHFCWLuV/MGgngGSdzQGEQZaYJ40BUaarLgNVs6yQg
8q+H/bZsV2U10iZq9q3NvIaRN5HFoWj5fcqjFcmlSd4K7GNIN/dwk3GZUdCov68V
Ney+C5KZ5jqCTaO4FSc5M5fPxrPG5GzV2DK+bUPp3YpX36/cje7X99c1tz7lZS6B
Qvcr2hzvoRZ8IPdcY5e/sDjqd4jKAp0XiBhtpBG4sJKV4L8ZhEoK6DyQ7+YXOJ7M
JsVCZ23Go3iRR5IJdngC6dBrrjGUBybRUUFY/L/rYGWP70DgZvJrQrKsU7eTS4qZ
ZpwwxVUxRtrFgjx/A3dyMgZjUEGw7z5ZjKIyI3/7Ku9dqiVt6e+t4B6iPQL0AMbD
9K58yuLYC3H3rnTQ8hR6zVMCRb4+yL2idYCxvtQ+CSAE+gIEUMGGS05R7G6lXEID
YxCAaBg+9G6vF8gCOpny8ErnYFK52eBEqaGmmEYQADBwTKsFbbK2jWePoXjFG2vv
qnWnYVS9EVNdMWmoTAJTqPnpruNB+TXYqiZhTvsAt3Ioi4WeGyvln9byObrDGzku
boZWVQaK+f54vcBuxSMZJPMTqCLKuCQuikwpvKOdfjv7e73Rxt0wuhfae6paIf5u
aXI34y2MFsRz6dAmTY6TfDENErsqrpKonc87+5XTTEEqA+toZEcUM+bthq92PeEl
8GG5GHwio7LayuArJnWhpcFmbyCp4LN1AzhuHK7TuXMVq9ExjM8uiDXP1tFNHG7r
lGfisRm44gtB7NucD05EgFViJSsBnUwVuGNLkXKWeCc4O6Kq6kW3xI035dMen2cN
42fY/Yn3eEXtxQ4zEgRZ+sMdTwq1a+g3P06L9o4OpwLT4zwwjbBZtfs0m7mmq2fa
PDQp3JRsA8MLwVU44F1GHMj2Lyhe9wQR20/uzWSUhGtYg1SSPc1QF+XLQTaIsZWo
04zgzkPOZbzY3gUATqp9knEy2lHSINOrs6JBz1cVW9qgfUxw7idhdItIi1lGUPdu
xonqoJiiRxe/Y934LOd+nrfblEBlZKPDLPLGhJNJsXa7BDcKyAiCoRHopqmc3uDK
frIulA4/DoCc3Lp6OKun+ZJo7QBoDqzU9OiWK7udBBQ1nA19+Zjh4uOkxT9Yn4Yy
A82JTtSxqJRmn2tsGq9mRQZm+/3UvGTDuCOz+jKThb5rEUCOqJt65LO97zFOfjwK
K5A774B0ITDHHhPdLazjX/NBYrqgrrXsikKSUor2FidfVv6UnvPVPdtP7AeMKCAD
zR3+cj1rgFmfGIU1JlizDwZvOSAcY4cZMXC1D7zQ5Is+qeZXZEOmN5bstA8GF6y8
1Jd9zNrxVtaJfrZJ+cuHuLCWmP5zp0Hj2BurOUSUfQUqvYmbz/OgQWef89DNQlQY
jf7cqXSuNUa5e1S1WePDx/6IrZ7SF21w2FC6c2lh9NNdOa+WiR7nuNX32bfmpU0h
68qkxc8b/ubXEBxxZN6appilr5mH2uXDGRfMJR7dX+Mw7Bdwhpfgcdxqd07fxtOH
tLTZdKper65n5uVMR+C+WZsl5M14P1zDqZKYxg4R2ccBJp68FghqGUkTJLnqhx8h
Q6U9vZsYYCbJlGDIj9gQIXIAh/TY+/AJdjaODX7dQe+dw32cE0vTvOklteAakHJq
zUneRnc6PJOmaaQO22+ek24GcixAMRgQghqjj8cXcVvI1aZd1y1KUQB9XGUUQNrR
31AMhihmseaZFPwSXCzEuqaJrNkuA6v2qNXcEMOTxtIasw40KHxv3ykbrXmzMXCX
9xXucei5Bl/JMDWqVWEU/Hqm7U+AWj/2tt+NCOtswyMUGHmHB0fs4RgiVRX3iinK
wtcNm82GwVjsOL9P3aG5lw8HSbQWIcDWMfhpB0ocMNf1w6CcTqBSx6WV4HOiBnOS
Vmd7Zk8RgCr/PjjuaPXBROyyX93KGjhYDQbq77UDK4+3AJrCzRigQ8U0k1aLCQaZ
pqE4x5Ak65Yjemd8FC1y/Ffmfvx/cV8FI7hE+YfbiP15erGYB5XlRE6nXrJMKwdJ
s1TZvpbfqpbJ9Moq84aZExE0IHoqrwtLhcTGMKSU6Nn4sndr9PsQCQPExKStZtZ8
tRCXeYF/T1lpkn/2kzyW2dbAmLzjPNsFl2PEWlSoZ3bp4oqCrk5dywwuAz/KykEz
S4YRGy8QdVIHJl+ZT9TfBsKykmFW/cr3C7lTrtPTcbWAgPymEo9nRUc/ZCHEg8G0
w6QChHjDiWB4MIqTH8SC7BsdIfINZEV8Co2iaLnFxFczewXEEiWAF6iPoG+gtGa+
+D2scSOGPYYmT1HE8vVJ8X94hTen8oc3IouoaVHCXblaLKY/cR8Ez0o/e+1avJR9
7S3sdW+MO5IlTy0xbLfuPNwWN10C9h7OYn5o4U14pJ92Ya11gBeMGPZ5VLpDsiJU
yw8ouUV2wwl/mVE0sQTyDmO20L5yFf+LDElVX9yuU3uTIzhpTCRq9BPt/BdI9vhV
MuYd9AUToucyDPS3W1WxIcmPcoxKD6MMkUfBbMAiX2leSucFxrez+XN7OKeyDmox
ek39OmkHoIiEtJ87Z+yBRSlk64oYY4RmvsUgsZXqktYN1UYaFa3Ydh8DScrLoSHk
z7QeMKkZasg9XAowb82C3gE7nLtRccgGZFbXCbRrXVp0TlNC6SQOGO99APgcgW4N
2X/fDDYAvdIk5+D9jzMMeDlyX2M81oHh3l/MPlvgOPQJw2FSldaXH99+oyNBjSAH
Sz1At5rQUdjvpMnVyBzIvTNVCc2yS06YPvYs5QZPnHEsSBNKUE4HDyQjCFTmhyk8
JSHhPnCGE3Px1w8j3g2FovrkV8HZia8wasJ+NgKA774+cainlvieu1sf8CM+RqMD
f+iswOsSq3Nx19/uWGygAddwEDfIIdR6VRPcHTBQYASqyns6ggBjjYZzSkH1XxZd
oeN/uBruAIi8PrJ9SaNdOtYUNOguA38/ppKKZ+xU+qGSh+2Rqt89LTgKFYzjgY2h
xJLlB75Oy/la/kKOCmyxbLbGLySp7FOEsOwFQmdTBMBBAj0MLB35GB7Vjf2XodIn
kQWmiZ2rA+uR4rfolK7GhNJt1sJMOzVn+nSYWwUUPgSUHmSWrVmP+73yKCbYVlxN
Yq9XX/R+CFmDGlwBpsd/fIUbhn4PYpaq+8xdYPe4KdA4Y861gtwPd3URDSwy6s0M
q85+dc1Cny0q3k/Su1j19wE4AqIj746EZ/WgS9S6t8FM/UqJXD+fOb/fb4RiC8vm
e4FrOIac3nRuWPp1qPa+wN7m+pud0OXxvg8Iy/pmH1jObKtFAXSTyRsFnoyv7Q3+
wb0ca368EJiOcIpRsChs9GeH6+USmP+MHqfz60p0QRpjabRA9Zc9bLd/LNuaLQxX
sxzs0Jp1MBBHyNzmwaddx1AYDU9cC1vbOpiRd7ZZo8kRo8ROCtQnKh2vkOO5zDCU
/hHx1hgyPhbO8Ju5hl/EY0U5K7uR3m6BkwLOeu+9Hr0WCVtMv0o2iq1Dtfn+hr9E
z9LnWcMAKTAS9LwrihuMP3yc4FqxYwt7RHeWGPRVI1bPj6Nb2jAsepaY840H8qrk
//ZoQtp9N7znK1sTApebwSF0I+5Cna2mIqtmTo9Qli15xY5lOZ+Z/E0HwezYrwwy
7R0le/OVb5F/lsWP6uX8xG0uoWidEUahIVYdpJr8dNcnfH0p4CFF9FS3m0UevyRi
p9TPfHfbTZFpzsyHjtwPTvLGsS5siiqb5nEZO/pSTkmLQnUebFRajRUUApKgwBEQ
/LoyVcr4na1Rty0gVxLyowlyRniTvqrfofQPh25cUPGqUccGDXit/U4Xq27eKGCB
J1h5/K2r1zLJ7hRwbz6RVETQZ899lS0nTcV/SpTtN/mgxuSzkHVvG1CDx38A4bLq
ryJqaX+Rv6QENFjFuNizkHZTfQLVuHzHFBoHJ/0a/8bPLcwg+u3Rszz+Nib6U7UZ
KQfcU6AqvbqKIwFcLxMLI8BFhtVJv2EBXdHkS2S5kKNuFYQ4v8GTnzFy04Jd45yh
jRDJVR86YhMiOxPQskkfO1Zot9pZrjS1qVZ+pHI20UaWsTO3acOu0bmpSDU0APFY
AjBlqkI+FM8OPM5mA/yw13rcW+DxdTo4LDslANTIbk33UMeYXhGf4JG5jyumTZVv
9kcGROgRUolevBHM5oP6EuHJ2NZOqy4T0SgTVyOwP0RgRvx12EZ6iMwKzFUW2QfB
PR+EyXLqsg3nxHVr5CkC29g0wxYmB4sQw7urpSQdGL/RPxfMmn5WzVbsC+QVYto3
c0H+Lpimb78sBiuUGJzwvpbAryYhik05N/B7Vp7aLc1N1gu4z4F9Ei7k4reGep6s
Z5rtvoHAYW0hdEzc5Pj9ukF4COazSmj3tpmq3L4LTFY5kcaHJma7ALEJbE7auQzf
fCTMfIPP6MYfqldxm67cJl582RltpxxsuHMrLQrj2GIJ1GAZTHLSGX6Sul66O06b
W6BVj2c74Qm2B4fYwbBVWJEojIO7jGqoBF5b6DSmsMCGPnFjhHwL7LM2tocRDwMt
gsJSPQ1oGUAiWFNhI5/sxM8nlw40SMBqn542MbBB/F0wo+pp4zvU5TMpZLfC6iIU
t2I9yzZkQnDEEtc704Sn4TnpFsIIpMeHG02zj2IAq7zXEbddO2MdVyKqXhVtM6lT
zdILxfYERfB7+F7dl3Y9jGNE/9QhsB3SejIEmwhK8Nw1A4n07S8ij26bES/Sxjag
E2bwpWem5zAV1T5TrVvNhKpSnnYpSbbJkC/69RfkXCH3PV46ibC1QIkX8d5FS+KQ
3qQfMsdR/behZu6dfJj7n8FwRIOWoV4z5mHMPbmzgPX3PMPhayBdmzlIDvgIgi6I
NcKZ+nUhNRMiJMhUuKWe2uPyGhgjcye5gCJuo44yutbSQw2DIOjzL5PU5wI7Ewj+
i/jdCLxQdhbVf8DJ4m0VOJ2u98KsxryYDhEky6BkDddMtwb3XsLqxieOBvCMrLhJ
ORx3xt44/jCbTPlGtv9Bet/pk98hMvzOepNN2paI2ik6LRQ8njnGa6IBZbTkMRJo
ZGachwluO77QWREse+rUMjT9/pcc5vp3Z/qj4V3JAhoGLikWNY3gRDyZa5p2I+UB
ek2e1OzMFvwm9hK6KBFtwN3cpq1TpdL7fbuIptKbNchPtYBOsH/BcyDcmDrHTpn4
78kjBdd0uNzRq+UWb++Z7vJH/WbIO1rGFXqgtKztK1YKU5dnPdh5SmzeteESSL77
o6trgZPRW1t5mVwlBxamYZR131jU6DaP/vfg+x6Y5N0ygB4HzM1KMfjD9EWez8uu
4H2c9uH0YyjhTuSj5klys4Gsm5Uqon2GrZhrjfkreClpw0x9szioItFQrDyLHZwh
Pg8ENxIj6Rbb3p6d8T4TzBXyVs2Vllk6TSuPMdwmPUoha2AAFpHvJj85JmFuTJdw
5v6kv6MriMTgkw3+gbwkKfT1B1QbvmCbljDUeTeoczqWnitIs/es1V615NSpX2Us
214iRhoaxBBeMlTbfvBrbmhu2HSUXZTNT43FvKx95Q0roUJ6H+cufNNTJ0dRWyxU
dTVpzwUVtxcz7J3lErNDV/idSy05rxlgqyohKUaABseOXXBZTZuZg44y6C12zEqh
YbKyTtPXaYfkTSom959TDHTE1yvtPVFb/uAes2B9z6jxZVAWX/WLBHH/F2BRtWBV
ipKaMrmi6PfGrrFEO2qKpOgjYAh3FZb4z7s0IFEunBNwXe6c7wm9qoPvo+iKCIGk
NQ5eyHbNNf/qEVmEA4wKYB6eGDR0qpwqxcKD+9+RXXAaaBEmCv18WGfD/vgKpePf
JNOfO6bS54B/NbXJ/kwLKWLyFQTvUI0IeGjD3Ux+sJYpOnuL0Q69WfgVsnPQBq5b
9dyC+sM9VsNc/f3vmSiLY4yim/yBMU4/NEe95g2D8Bny4Txlt9DqVzO2mqz1cYz5
utTETGKYW61NoNQvsBH8z6JeKooeNwlQ7ZGhPtn84cLAfYx6OYqC7Q3rc/DbLj9h
0EHGZ5upGphk92B5FIyp9akFLOPSmMLRCBUzV0tiH4pTEkFKWpKJ7lJb181fp83t
bKw6MZwCtJVjV5yjHp4+MQGnJu005mzEtFgX9u5UxH7Fm2pDIVi4cK7BVmUy4dsZ
94r/CNGauCV2AhprC+A8TksLtScOPwNnkJ9aXeJjK1GcuyQIFOpBHBuhzmKp2oJj
Iw3CFZ5QMUuAqVxK5K6oZXZkZuQ/4FeuCXm5H+YVo0BgzM8cAxOR+kx+VXlbxSGb
hgBuY55rXc+uUA2pQZyznA9yYAV/ueau55o4Fz0d+ijlzGPYSkl1DvGIAn4pEV9C
X8HlJq4qxNWz1mz+jIuDGOh2JCbYgQ37OiJ41m7HIK9qYepBqpbvpFraWJFofvoD
enrtrr/iV2nVKaIHUQT9sj5LKNVzMNsul1bcOlRvIfm7nj3w7y4V1Zcld3IUThCh
NrGkibGNTM9OtRD9e/6OsT14DorvS5/0Zm9rjg/rX1cHkkFiNPmSqG/4IzNvhdJd
n6YbHANQ8ISbhXtoD1259b/u5E9iC1H6K5lAh5lwWDEfW4t6axlq/fcfY7z+QviY
1w0qgY7XNemQZZHB0R5YJhWwcQwQQ99pUxJ0IAY2MFRakIoviTJsz2GZzL8kokhO
GloG7cCLpmtcLljsz2XIxgB4dJ4epMhFRUEwCZH/LAIkn9SFvNjufXGD9liOhvjq
XeKzBjcDV+jZqQWD1ny4VfVVDcv3vh+c3qCl8svVJF2YlxPFgjbF7PIn40N8orYa
ckeHUoIYToVd9iGmKuWAgPasWG1fLkTTYQNRFYs7+QsYWnD3d5PXC0aBn/1gW2p3
E3rAWhD0om7MDt0SSSZHbv1Wid1Gk8+adAjZuFE0cdmrcHczcdVMsi3Ki/nmmhwt
6SDYilMWnKm19i1qisUKWc2C2zTMgz4lEOypHmXrvMFOlcQtegAPqSTe7h42+2G9
DfpI0jsuf7YrzmyJLR44W3BmLIo0FycAt1oB4z9hiEtbELe0e12Gli9ncrZ/IwcP
lCsSwGL73oidVTSTbJkvDoRBEUNr/lNxmyvEpH60nZZc4cJECxgkuF/VB9zNWH4v
3Ja66mZHCkSRiAI73ZwecMQDc85EhbP/PWinrtWtUEfVS1xOaq1XemWVHJg5u2Hz
M8V3YsAwgGKAtxbZv0xw8Q7wWzPp6+h/E+mmyobd9K6cLeUnj/FtkLNMMN5XU/o+
t5xTXfJSDNiuQRPHN8TA+/QKwtW98mpbekkFPb+zVXt8x2ArTwo/SOv8Yj0o+MXV
to3Epl8LvgtAVwQXSUmrcBe2a81ywmun5qE202EElP1El0mD3NY508qecOpqEU9K
rhbu2w9lmnfnp6+iPhthhJqHehgvvaLhV6kuq9CperywMIvfhnZ2FtMQru3bGqas
SNaOZo4vaJTvbk9X3BQIdrf2pse+YNoI26GJ3kc2tqTfppLSp2czDgzQqLRAlsgw
SDkXLKMPOnFt++2AkCsJeIOxCHqRPWNFVG/yyQMWx2odHOVJFrY3pqs8oINrCexB
E/avaw8GWvI1dfJ1P73mnldI53Hfu12LGdbcbhI84nsmHaq1TFUqPKRp7YG9afnK
6yVfVwNMUvNvrqlSGS1zLmsMnf8XIRwFyW4KhrQi5OZSf0ObQfg8LLkXuMu66sHd
/X/teghRGPC7wEQuKT0PibwhxDQHObRlU7p778uhN27rVOtJrfc2N85NCNRdEPCL
jpgOhZqP8Z2/oDfmKWcSIYd0RzUfWZ4eWbgeQinKgAil+GBBbHNXN4qfHlJRn0jm
tlg/Xh9nkBeeY9i6y/LZFTd/nKRTeRTV2Sad8+x9+frhyWTdDFIlFySIQlC8k1pw
GWk+4H7n8Qa6BXmIJxxFcKILDWpwynkkoJ6FBLAYppdWvg5vcps8px4eJCKukbl8
lH8ntuw3h5hB9yY2tbksNgNUIPF/w5iDcjtgE7PXianBZhWOVpWtwVO0AfY4mWbB
YVjai4q+ur0i5viy0aHbZPJRSYc7SHotE9sYnn21J8F6gdKg/IZ9/m+8O8GNp3Gy
1qrd/7rBy9WfaKXvlmE/e7OOyCTmJExO1nNmWWeY88a29riONm2tFRMzjx6NGOJW
SFE0lTaCDcbymzF7gZHkVdZpB7VnpUDa4k4wjlMRGQHCrpfPeaKUy2lAvcBqn2LC
nj4uEAf3iWl79gvOwr52/hCfxn4dTefJ4zegB61CMEyLpH/cz+YfYCKuKfy6Zeq8
Hv+Xxn0tuQr+79H1iVhyqdkcnZxfh+uIXpWL+AoOmqu0JPD8CHepJFEsKxGKlCFQ
18+pO75XHVnj3kFC0178BFbo6ZQRVbhA0ECLpZslRKWXfXjYVzDVXmrD4CfSUIdg
A/B4oegPVJyKRcvJKc3R5+CV0JqhKOcmOLutauATiAQ5QNXhUpwwlVck/SVZwbJ5
0VsGu4LzM7mB2p1AvyTzQgmomgqtiHztfspbixPQ4RHcXcOtPih/3B7lm0zQwycP
rLxSn+nY9maYo/mPbH+uin4dVVLRXpZEnEjzcEMTMYQ1e/JZ3ZBQjZO4DnyW0Wtz
lvbqjVz95s9SHqIwQ8+4dBGy0lsOzpxPDJKgOyumJcg28CCIlyeTQGebzCcQ64Ma
MS0JIZQ/BAzx98H6NSigkWi+F0N7u/5jXu33Cam0zC/7DX4zSgEL1PhrAywcxRY6
iStigycuWSl/g7gzDbN5wsc6CKL7RhhyDJlcRDYeKm8kyCS5il00fLafvjZs0PI2
+2jMCmus1X+h1E0LtZcu97DDmNV7cUJ94m8x9w7KzggfUiM5aWubmvkMA8BcxzKD
3JrPKRadZRtMZDBxuOHDXuIuHY1YQtUBCOYGYFsczvQkJkdAZ0SmT1y/AxufXmxC
OLc5x78hxedLQePLRUxTVWIpB9NEtH444oK51fxaW9R91Vgy6McE1IOGf1nKzXDE
DF0o2w3fkbIj+x2UWzv5uf2UAU/YpmJRDPcPQubBL7sVFBVUrGsw/JnkcUJrJv8T
uPK+aF3gbv1kreeENNpri3jMZ3tlpwp74kUaVIql3wyP5TthznKBSCrZVFKbEv2k
n56JBX3MRaYpnrNiziL8fWpNHYNrEFcqZH7LE5SDxYGCftkVVaObwAmAeQkz81V7
bg7z89WpVydSuglK272sz1kydkRvpJSg0DTLUUPDyBYM3isaJ5xc8hOVi/S3AvxY
mAtBswZR9VuNOJlIEVqqM/qPKFJ0QiBuTORy5o0/iW/h6ivmuY5UAxw58p+Oo7T8
8UE8Gf1dKpEFt4R652YVGGRCoExlzPvQKdV7k4S8uaoyrns3D/C7dGi3oIUMXCAH
w3Abrb4uHw5NKfozOgQmAPQ/TcZaoV1eODkQqb6JBWBq3dyPYonS9aPmDLgbq3q5
arbJXZ12xonteV/LZiZMnezg7I5NsmayxHyjX4uGbKQoFlYyRAJwI4pfxyDcvqpg
KjDQYHqc8LUUA1qnzW4+WQdOv9P3lReFy00rvaTaDQ/8Z2bSKNvWZwDQN+3nd/y9
QOdURvdqyaX+xDr4VOW4r1jalejg7tG1Z8zxbi96e4vAQ0hLeIGKUn9ZoBuYC/01
kxXAkBk4958h9UfQTsvyrVG695YS8Ek5iZ+kzpzVtha+0YubUKqy7nmHaVn3mhSU
1TovfXf9fSnxpRWNaDk7a2owhb8HMFkbCUY7xuozz457QV1hl7q1CcMpVCvp6S6X
0lXaf3ROHhwGbOzYAKlfo1btcXC0vXZzMkGBc/bqPNaX5XlEK499yKmAUuLy5pGI
dPiqmLUhMsNaVvilMPi7xNP2q/otGKKxUFYmZ4ARx8RL0UmnXCKK0yYav5L6iRLr
uBXV1DLs2IOJ/SoQrY7CYQWJPpPVDZWwodS6adFKUWW7tA3SsB6nZOBzRrMWEVdx
jX0WIqCcQFYhngtFnrduUxtQAp4LgJUAANaHRPnw1YyttKHM1rBhuUaeqVGAiqnw
YRIe8Lgb8s0sVL0cBV8wkKCrdXphqmJKGQbiaALMtgJD/3CKk4uDenzP64h9Ns75
RJTAQcCK7EUKmvaPO3vjw9uC542vnQ8Vu7eybn9CFsb1pR+0PnnSmdhjcoyeFwKR
NlBH3ecJSuiYn0BvPaRqLXBaOO9i1xwX51yb+w5DFrFtpGfm9aFHYE6B5vIChWgV
YiHUqTSiolT3IX2lHBnJ+iosEiXNTd+LHi3eNfZFYWsbFWvl0KillxLR6C8EDazJ
Q+5ikLrmYtSH7YfSFEny3Gsw++GzoIPo5iZssY069gi360jtyT5CjkN2lSG5mpQe
zqOSwVCjy7EIaJWuF0EWLP2r8NJxwx8vdyJjtjw22tePJeUGDIkMn9tKNuEElYRz
b1DvxRZVeo5DL7i25L02kWCluXTPxY2AknRtAKEAx1aFJDgJZTSyfE9ZCCCiqdfw
q4Fn9drQsHZKv2TegvWPeKKf37r1ZsJDDtCbasJjocjiV8YbZ+XG1SD8H1DviRtJ
UvyiF6wBLSGAw18zoV866RoeUvgl68OR2LSqUVx6sXbJndTaju2zdLFbsHMOONuk
jhRlR7VAX1raXHzQE60MtMf7ZDPEQWVFAJNYzI0Sa6Gc/q4nc2WmzHBUONSOsigi
9sFJLKpcMKkDErECRyE8PJmzr7GPVm9FgiopbOmXw/i9u0in9emxDjsRdXDq4P5K
/jr+HZM5q2MV822SzbToRqoUJsOMdIEyfjEyP4KLWqo/xMnpHKMl3bFUT4lY3LJo
izYnyqscHJG1RfGFiPpvtQFj4gcDCpJzoZStxv0QQ6J9nUdkkqNItukA7+z5qruK
XoprQoH80+TapTJ40rP0rUpMCercVxNGrLp9EH3PSRQqztHJO2K7DKXL8REKh1Tw
we5Uyja2p+ObAsdGpRNk6lYMvVF5mK6q8U1IxhEoLPvB5Vjl2LMoG0KWBUi9+rA/
6a8C8r+HVP5qBAsh4/H2TVMJ5QXRUwjsNZ7m1KbKnkh1rLCVpiBC1GU25mbrqXpb
AwTevEHIMCYuX6oDGkZukFk1knW083IBB6ewrOZ4Vk7oQCNgtTM2dZ8i81UmlW/X
/svTA8jocqLbKbYEBYfl0YZuO88TcyVzg8E1U5CIKUoJspPBvEHskh03QDIv8mf6
zN0UEJpJNXOFCm+ypzN1st3gqt4wfI6in8pGzd9e9JUFP3HKYbdFvpcAMmlrrlah
nbETLEgJb8d9B3zN0a5yp3i6oRfkQcTnrhsFh+fslhV40XRXon/dc/fgDEzloi/u
uW/7GEG8S22yGAayAOoa+oRRUaq21HapP6RyKqAQOrHhbvAv/OePDbv19lvIZn67
fj0j44tKCHx9fjpygBXR8b7DUZLDPbE8NGQ3qyNZTTBRNtquOQTuAjtS8BYSqw4W
XgONah4AnxErzva1W7KwH1LPQbP+GBuefDPzJt9eBaHGxWqNJ2tbMcys4wIj6SNr
Mj+OOXenUlNSSbSGXX0enc2jz4COjfe7T+wiiHZl88xN6tJuL5NGqcItcxvK0u6D
b4Dg6Eq/YUw4pthrEFJ6wBuUbJhudHELo66c7WFk/KmHnwrE0mJQyxG0tU4ABh5m
C8xSJ7lgl8Qx5pyACZQWVB0hPW3Y8P7N/vAvFn9S9Tf8qH6y3Hdm45jMmDjpe7zr
XVGDXiNZrd4hLmEbgo2aZ/Jvot521iZAMgwg5Mh73NJbspRcozEdT+N6U8zOuU8b
vhB+zZitVdw6cAxxKdwwsKOle8PLhJ4DZ29V525pkdJ9xuBUsaeGfdDDxVSy3kgr
0MkRdGd+wnInSdbzT4Jq2LW1U9eDM7hpoCxbjh0i6zLY5z95o5HlZ4936AhnDRP6
YvdiTFSW9i84Z4ggfvv5sWK/rkofST63nuw2aDHHMIZo9qVU0zqu6czhW/giBNe8
QIHUsmH7Sy0ZrDp//FnHYfZfiSmEDuPdNENwEmsj/HfW2iB5KpcA3HFICfHX1znZ
sVKGiU1n7wJqubZ4YrEVSrhpiVS9kyWxBrReyc78AlSMprzEK+XBFWbaG25p/NeE
hESkb3KZ6XDJJWG0h2RzIcKjp4qgxDUkh49YgsbS6Q+g1EhHvHigUgzWHYR8+c5/
B/3VhCWzfkPUFXjvgFLD7tzp1H9DaM/9DUXMN6nS0Dd5TB3iVLEiyOSl08ki1m/C
uIoHMC9fI6HVh8KsNL8+t4b5TqDkUAWXmtvoGbVcvhydfW8vSbcvIiM30bb6eih4
414yFIy/LuWQRe4OOfN5SZTi16ZvBkXOIum6WMD0oipqwi4wq0tDoiKOsFv4hMBE
o3VIRmi2pCIeAdNTbqmnJ34cQPx12sn7HD0zGVCgIhsSnWSfMzkzcby5quk15pSQ
czUZKhmrR7spUo2EMkG7l2LEMsv/+U1yw31n+dQRH7097hDzZGL2kPzkVQQFTnXY
F4Cvy4ijpPCQf3yAaLlidgWQ8g+ZszKPHrVvmsxhcitkpndKA1CRolRw0Hx+mJXh
nxHcc840CGNGe3KNwJL1T4JxP9arSvAFMHW3+rbjJV1bpP3/Z4nPVHP8FQYZKMag
/zv0JvRlP6odxwNPl2Z4pJoWEEU/E/LjSKXQRL07sDJ9znpPEYutRXmbBga7Hns0
M1VI3WffSxsvkUaf3faLbXYTjHDA2trn/AJMa+Esl5xzRrtH6LI8OHy1fgdg93dq
sO5ALww0gklTLfaxC8rDwK8kOpdT54ubtJ56hRhCjwq2j2srxJeLGSKRj3woqqvF
eZ3XgVsW27tQ/kut/1OXXA5lMpth+wbzo0cuvzZ7QNuUctAYIjHdbeFKRmqAtaC5
VXeHej9rex/AwFCxuEb6KhTgwVEM9Cj2vsJZo2klPfzLtVltvS6kbCJ4k7AAlC+5
ofmQUnUxS7WVCeUf2eDvBqgePVZs79ENRKk8dhTCJza/8hMvwHKvAqgwGcwX/+JT
TMKKXDBzSBFQ4XGTpXqiutdD+B9nzlxx6AZjPtEGjnKuqza6UNAslvZpVIMTjK0h
A7HjnQV+UUQlHu+JC0GUN+yWQqWBJZoIcGMaNkL9DZeBlWSQ3KY5I3Sepjkd7Zki
zeB+i35821E3KoQdFzhNCWa7acx5Sx8C5woA3s1iSqG1Jjiq5jWgXuUrOUyZXiVx
7/pHxhHvbranW2z2W0DAo7/X/C+En32dQHe8DRn+nrqvXSB5/gBjlBpZCGPaTnts
rX4IrIEclDwpHBgUg+M7lq2Y5OAI4Op8LPQp1US2lTLodU/Rb99QjqF8CKCF6JzG
vv0u1L/aRiuVPR+5I0iLP1HFEX7QjiS2XCANx/oxV0UvjoCQMZIhnm8RSatBjV3v
12O5WjTjL1yPl11tJwCbHYlw6cnFKBpDa7jAx9xHrAzhcSgoPOBh/hW7aVxUi0RT
ss5IcIUhkYmMFdmDTovkSWqOQQl1KHgPAXEGcNbskbMLdG8ht8jFMCFOm6gfpg6i
T7t/nDx0Ywh/pAxImyz+U6JlCYU6IhLuY3HSxEoXwNwSVyzkpojZRnPN1qd40aNT
7fzTOGJLcHSSJ+artUqzl75iMTisJ7/0tBcDMVApuLR20yt1ZehW5D8xe4IBddXm
p957qSXiaaKwU67qS9B0bN5DKu427aqbmB5PKDGerbKVsyWRDygAEI1FcqDlGN0c
5NXopiwa7JVheK+wVJVSUVcUiDX9Qv2hSR5otY1PGpgqhIoguGWlwGnlnUxqZpAS
2imE6wM4X467ZPtUNwBlF3Rh128DK+A2wvbzEj6MoCkZBz8YARJpfY+NTNca20sf
s8HhjuFuKrOx7LtEf6zgvM5lEGoBXyDF3LCdvrwd4g1JjKgzCpLpuGvEKTG3SBHE
VWTpvYl3tuE2/3ePQnj/Fgg5dhsuvoSuil78aO2HoPGyTJJRnQs/uWaJ30fc0AOj
pPBOXZsW+v1+e4OmxuJ+3Pq9ujcRbYlZVPnEidqHvU9sYp3TzSwRNE8dLGr14z9y
QuaLHqq71AIa3Apv1cgGefTP4Ax1s73bog1Eq3hWoPaWUAseQ0td1fOW77R2eHGD
v6XGPoSo3vj0hUlRHFwkB+r0A2DfIqAjhPn5mawxZm+/7qG5S7t8cHVl7Ya+P4S5
KaSR8v6tpTFAPqsathpp1HlSTZkMjWOydPb3yxCbDnZZ80ix9Jv4ANXEk4Dnuxkr
IYksBlbiM0gzsdNmwDwYbF5JHdE/VastyGi+vjBWfq/xuXzroHx+q4w0IKBVVYcM
TUTDU5USvGpmzrKoLBaWkTlECkbR/IjhP2IrSynPWnch6O7h6lEiB6xRkpAcOz/G
CFHv2fQ+mlf3pAj+isyu1pgql9GvkvnkvS+iz08YTLGBO8T++p9iWPw8aCLHKsmf
x9qsWpk98X1yCKSbUp6WWZ5fGxo/jeJNfoQWHdCMJLn9dnGwr/22SBLqCgMchDX7
USC5/mBx0eE5DzyRg2X+OjdNK67/KyRBYqFJaocDVYFwQ8Xo9CmhlFBEvr0iX4CL
kYYI2RlnRyfL+rirzmi7cJIHfhtRU8t0EMKruf/r3qFGGp12CvpJ/V2eZtrtocEe
K9nUMoKDSyUW7/rf3RfdyW8OYAiK1vpQMrxU6D9EYAEGQWorLtYbIgZA2wXPJfPx
BxnClMaKfsQf0iOkJGH2f+dYcW9ozIiwYgMZ5/FCl5o/vy6ujNIOMGZ5tMK/oKZO
olroTLhIPisw/9mWRZIaN2jJbQx4AWi7VDIrw8JXCA/74fv3fRJ1h15H4S3YVbFA
Vmn2E995kPwQfssJDsqgshZ7i+MpVkCXi10quES95BMkNzVvmaAOSwjbPpYAcfsM
3WWqd9LzYbHk+ySZ3jmly/AeMe0SjrmHfk85N248ZSI6Z7U6U9bmp7R3pR+74N9i
mYhGFTk8R2Fl3ZfkQb6g+K+dUnJnSfmhAkmWyecbDIGcbM82F/ds2XXSs1zI1n03
2+7UAJiKhO0CE7MDLgLssgOQIjwnF/DHnNq0T8koGoDy0ASc5O0TOoz5GjdFYP3c
6C1VtTrs/J3gfJqTuaaPoIHqnkWArPU/QLttTyWLGbJ75HjVaQNDUGSz1skeWi6h
LwKnREAmQCZDO4O+vb+OE6DRuyCp61MWHtb2SNfsEW/UC248e4at03j3etKBRaQB
RVTp/VeiSYw7hqvccSCEw+WuwVAtHPQu2as5SEBeV0F8r/70OgDDr9B3bvfMxW8s
ObgHchr93UuuorJc1KlkjtfP08CTqeD4GDW+UKpeYgBBGMGhocvXs047UZ7wM/cI
bFyaGES6y6jyRs8Hu3b+thCL1svoct1p4O7qsjECRuBoymtTrKorNzV9xZKDKvtX
0h7CC3igrA+R5FqcF1HXzsWDeLcqwjCXohHOfR+sNBs9VM5Xk6KjsWmxqycmw/Cd
OzC/XyKVyPZzV+ANl13/QR9/7Gz1XvmA/id8x/GCkAGb4sgDAwI4ST3ykLEYvzNu
M8uzQaDqRwaqGO9GWHJ0ZE7TahaCA2zbow4ruCyBIm2E6AvPZ8Dmk/aAzEMcQuwR
Ur2JiXxAXQTDZ51BhIB4FHmMPd2w7LKOfKcR/bC4t/RBZR86JiP3vtCLlFuTA7Cq
dn6DirDKfp819VhqdV+3Mu/c3wrogcV617H4s+KH8VioiFFLoWbeApamC6NOD/qm
qASdGzmH8mMBKlyj5afMmZEXly2gNt8DPrkJ1lLoaVPTf92N0HCVbsjUC2oanxyi
MisRB7XtRThA951nQ/1dPFR6u2yCGpLmM+1mIzK+2z2Fs9xZ3CFtKtJiSohPqNEC
bIIrxcJ43MGXvhwD87Y3e6YHJSrWVolJT0zCpaLt1KbiOZFdRvpTcrkf8I8fAKA8
++tPzWlpyHwwA9l6+C60LqgQhBLJDkkIyBMbNVbCgQc2l13v1IGp/22uNz62oTOq
2IMgW0IdZZbkOt6abo7BItokLMfBv+zhf9O1k/vPCfYsQOWsxpQ1TiY+04Y9HR09
TuZ/1Kqn3e2XTxgbfHJhSAQc3nC0qys2tSHXglAjtg6JLKsH5TYxl/NHhKjEJG4Q
n6xY1FtTPg3NmwYerpbB50UJCjFaf5SK8xSgNGNiHLjX52uUMZh1YrZmw5gOdebA
p3Ss4T0LlBPVcDzZGp2xM6fcGHpCUA5Wx65dorwWsQvBxA/1aUm952Beo8uz3deg
4y36xmPrrXwFRlAi7CUUAJuYT3rrZ+FCYFnvaUPCdbinsFXOG7QXopnAQkoYlhra
TJdr9ZQQ9krc0y7RV8qyyVuV6/CkNal07YhkwNB1iK1yR///3V7vJFLNEuRV5loN
jBFKH88gzt3QrIsB83agwxoQR/FGpRNvZTmu0dDll16/GD72oFUtMitcHkXIG1Z3
VGMZ1skR7nfX1zRt3dKfYZd/v2vy17+5sKGXBOrIWpKSfYs6WtBFQPCtzR+W0925
+5YWfzepmpL1WH8ssEwJ5ySRnxaqv1x1ILpzdjKLIg8L3GAe8bXx8FCQiwta7d24
bF9IoaalU0hvqpmrQ8udzepePUEE3cQ3WUrd04gsCVfpBfyVHFjK6Oldb/L+ZPSa
i/gouz4Zf6Quow5LPTRhyjRnMX21/CuyTQ9yKAviW8yYcK9jxYDn7U831PUzCLE0
MvDXL3AJRYEqWi2eXvnXuTMTFFTJVYkCnnfirJXomn+WFD3fAaI92+LM/Guprn3S
uUrcId98xtebYCMrhgR8FMAIRpd5/s8XHrcyS7OkeIdGgcudvN0kF1fmklmUb744
pICtjnaIISQ/uznFTkkRvK8w9CUbfkxl58OCLBTeX8pSSPNE8MtdCyYh9iHmMcZA
fGp40Jb4Fttf/MUl4Spmh9o9BVc8sgzAFAETjfmDUC5x2ywYUcWXnCHzVSp1cmz7
cUJ8i2rwcAOIAut7X/Wlum2kvd7c7lawg/sG3QWFvHnU0iufjnfLYEWKMBsuOlkQ
Y731OUHXTO/K8P7j3bZ5ivVI438mQi9MKwQnifVxO3IxhFtrodr5fjCOJ1/0LtsI
wrFj9gjzKcWkUQ9a0+JzlR8mEsSuKOfip3CP8xfnJBn5CrXdfQ/tlZu47ghrsChx
51DS7Bwsji6OuzQpQqVVsm9U1aRw5D+XGinfJ4df89wXiwSuSaxIex8sFDqzL9p+
Yu+pTbjOm0iCIdaUMvnJIAcqdLasbqpNgpr69dUFYLT/q8lRvjBrCS3eeFsnjbBx
fn9CnooBkWUa5TlL8y0Axc/Dw0hW9XKp/vBgA8M7YJ7pkaUgZ2mLLD2FIw1oxQEl
Soms0KctR2LerWmg0HDdPPom+YOpj5C1pl9z8lh/HOdh+tp1jo8NwgcXs6b4+E+B
vXTAwENXfp4xWSdazwgVme3OSSfy7mmKyeWXqd5OhNNWEpQTJGarNgAEoEAzCt3G
JM9xt72UEup1gn/2Cz2svyp5SE0C5wF10C1c/w+8E6pEvs5gTzxOAHGyNKlPu3HR
fq8y+VNdIdmF8FRO47iQguG9gdr68mUFCZy4QNcVkyYyzRqayXVVB6frO8q2IbJ7
U+FQ9Fx0EuCtwaga24Z7Ljs7WKEAtk/GHinoVml/oOW90wMaTKsrMC67rchpBk6j
+LbbUIfQ5LHh+fvcJCpj0rm7RRa82kctsBpe7Aon2oLJVhEQ68IT+qXrpUz67N2l
nBkRuANtlZDsDa/5dH+lx/0XFYtT0OuwP11DbX84j5tmKtRyil9zJMe2SRpj3+8k
ipheynFpTmR9O7fwfRBKf21kJQ3ySWKl0pLhLue5S+IcHPMe2wu7G8xUbVRX6/S8
VFlP1fpkPhw8sgA6nmSwrLXJkaSH6Eo3MSu4fsYgrF3iRFHW9jG1YsG/G8OrLoS+
i6o1y+wu6kMW5KJ4W3lIBJBlqGmO4+gNk5N5Xto1DyfrZIWFXCawWkXIQ9dzvmFq
jC+HSMDtRL6Hv1y9t1/OcJU/M4m1VAC/skWNZaQMxC4YjEwnKCmRfzmHOCGE+99s
baIpVWQ8/cgeoolNh4zm9r3tLSMQaL1UG2KwfL8cfWTEj1E+WjtuEYNjct4WU375
/a01IsdOb9+EeOgWuyLa38qqox59bslSL+4XR9eFfQezutAS9rO5WC5dn3WqcCS2
OU1TjPjTyaTgrYoNWesjtxVXwYIzadQsaIFETlz4MwfEAE3EGgb6i0ppc8j9IDtK
4jhnw/ErxC24J4+JtFkUkVyEtQvk/SnAs+DZI5S/2U9wERmLOhZ4kMxCFjR4r+yx
BzHUtzyoWNy5pR3Mw3EXEbqg9E45+wFZNZmSC5yOsZgg8S8YV5avxZtWrD8GTTgb
TZvlFIH1XRRN+bQGfTfzkXLdJJB+VrWfQH8j4gIXCAFhszHvrvfZNiFnO+KOEw+N
CjxFwevttG/7vdygg4sOJ5HHfri4uSxCnBz4BF5KUaE2krF+1nGkzP6amI+Khbte
1AHgNbHEaxzj3mswOtEBsr/nkxDfVElU8VCTuGeTttCZm+iSetSg4OSgsKWiWw9j
wQ4wuYZgOdoOa9hT5k/TlXk/HUUw/dp543zZlW7aCF349NTEbpXurViTk82Dp319
reUlrOgbdLnqER/1kdq0qbs/0QSBc76D62Qi12M55MRNUe9a0RB9HzzYD2yzogla
PpWoqEXc6grLVi3LnWsrh9DWJdP1i4Xm7h1QCC7tM99fxwjTSOcd6Pmj5AZl1uix
2VdgOr/bu2uW/m6sscStOpNQ8SW5fw7sv6sttzk8b8SOxTO4NXaoHScG+FwsTmmQ
HnZ4dClcB/Vj9qJBAuoNQI6ErK7NoRFkPyQE53AF3mE3PhEZPGpT8mE/0uTvCKBY
wbtAP9ai0fwElExpxypYhnYlbJzk38UBi83AJNEFyU033MY1UEITC5k8aaSUw7iO
ma5uEvFxHoRmzeYII8MsUWk+JfrP78QjoT+/MGI4rfpaTtbbvx8Ox6nyfoFDiqvt
1bLyoAtO3hj7eFf8Bob70BYZevlkmFwvxmbpughyd9eUsS5XvaPhpIspUoIuy41+
H+dXMKtWMIwkVx+AQGoWTw8FHKw5NVlCkyFSFb44EPT4XgtRcJY5ltrYv/K3O68G
b8lNmY+x+0n8gGvSje+Do98cZT4UsY82p1QU0afMjGusuTg44pO98NRIpaktZ7ji
8/gt+zwJzFgC2EBh3ThKoswhF1BQyBZV3hEfLOUS+3gYhBPxmsrRMT70V+fUDZo0
wRqIgqPMhlMachy/AriIQYZqCzBJorQihosdwZMM5fYbxCYxNxwaR5jN9PyzOf+H
kcO0ZEfed1Y1ZdAPYT+0YH9KxWcl+6a33P30IdFDMX8MiGvp4f7W+p0E2l00eC6t
XNmVGolzEw/GxqOWU6V6nyf675lLHHhWuU1iaRZKAaiqaAQ+vhSym4Vg4pnmklZi
va62Q2daUH2VxYD5CZeUj+lo9ivGfDvGyM265yE+AnADtM7jL8rmtSs8mnHFW7AE
9xGO3tYDYsKcg0BQEi0dZ5bTEX8xRsspu0753at/0x3+Yl/q4MLoF1hHD7UxS7E6
2f5Y3/8b15u5bLBHZIYa5/6wzeuEZzTIEwnx8KCIKlZWU5RredEWiYK9Pm+m+h/R
IlwK2ONKaOcdKuSMNUp+8lKIc/q7GyVASYtA+jpvzp7w7rQh+aF1phBVkQFUSbto
QgoQ9SqpafL1QKYwifQcTJ4jtWH9DBYSOmBruoc9XKTkhZCPORxO0MvTQo4SycSI
ZZWsJJgddemi6Y/KiTsGh6D2U3RcCoorVbHiTJShDdFMfOyrDi8Nr1iqJ3LxJ3MH
WDFKw+EQEx6Z8+cL9m5eVjjIsNMMHdzgB6xpL7Uizk3BpGnXbATIbse9u8Yi5yUb
enAqdO88sxp+1VeUK/SGLS+BfvGrS8qeB4WWwfu6cj5q06+23tWwDYMpbOa3Y9UH
VA0fahO0G3HZ+NOK8h2fsMxun0/KY985WM5Sf1AHNMzWgrlaq+VSflQJ3ltIbaQq
QeQpfLzwIKLAnp8DRsNM2RwC7xBJStpHZSIZmgiZ08Dn2ca7kppackM5lLMz6rMV
FwqZstgDVCYKV3gfUOe7SEdnJHoHRH4kDb19cDjUALzz8UxhK0J1S0la2cYJY7ul
uNlTg+jH+l1HYLdbh5Izc9mseiuS0ucR42x9aW3+0XynZ1qLmO49by30NcL2XJ0D
bRKMnSIpIIGJZNFRqYVGl3bcWL7Mb7VGrbofUAIJfFMR/qkYZYADoXJCJ1Lcn70t
U3OS0hEU28uFx8roYl6r8XcUGLLPW+YU25kwIrXJ62YHHKfqXX14TqcBMYQmbBMJ
YJrEfz0J0CqTbHftcHOFqWfZuVkN1ds8CwZwVRCgNHs3lK5SMeJmDM+8FHWIwI4X
IAA7gKXxslqSJvBloSTd0JJSUA26hdHNS08+yKnPLzKDdC9mojkubn4mtfcjxfPM
aSC7f+Keq8v+Mz1IG8DcQwP+tay5SjcM+GlKoAeL8oiRO2CLIx3qBtGZYYQmtvTi
HPR3goruWo11L9pq6CNAMieF8my1TR7hzZVx2RwmiSTS7GwUnFcmj591aJXwaDpI
MPsnVoByf5xNiipgCehc5AJvx7/z9N0RiwoNzcHQtEcorgtrVbrsaqeJDCQJItr7
wtB/u0VGSijJnODiOXOyHws5jkp9c6WkCRPf73Kr54i9eMGQ7AR6NJO+xTJNlqB7
QvkyLAQNZ7dUyAya/g5sqKeWG+Lci7AqTldkxZnAPQxnmhJywl79IRdf/Q8eijYT
ld3dg5HI5f7rlNYxJUO6IimnDuRej2butQau9nRnk2ioROPX9NC6xBkZb9vc/XXx
YTUQVOS9aZIu/NuQHyUJ2JheMhIQC2U5PVHmCVzlPN6stfUJb0IzpmwllMXSsxyS
NFnGvNENy0rzBZqsiWr2d67z5Z9a6QrXzY0SXZgqEgToR9WLzgd/gBX/CQTSRwYX
6LvpoBFGOCH8bwr44r+4ae9w9oV+snIc9BPCA76vq7r+PRbBHdNBJtYViDDX2HaZ
Y6qP8eQ053npFYck/ftlrflRRYKUWr/ilx1YVtrST6FR0RvGLNxR5FjV/vA4CSKw
R6ekByNYuVImtrBR8RBZUZfft5A7MoaF+lV/ilHRABHvLuOLEHbK6x4AqnIwFkrK
m7LyJvco4jvGM83rgn88i/NHDc0wcj2Qd4qwztfauHyzzMhc9lNBEzQPR4dhADMG
M5wOpE01W9FWfbW/ucILQd2g9NY1eLDYDDLadSf1pp+GnJBPUqJneB7Oy3zio9Ny
XN0MEgMLQeekgxYWlyKFQNQUAM1fC31CsbYynybE97zHYaoew1/lpvih/wOtizux
UrxgeSd/ammRDJwigGL4OHSNj1icN0/3rnYshSfwsirb7Qoe9H+WwdC1tACEs9lo
ppgju9Qjs3F49VRzKPNSdKERvSJMhAG6Oc5I3UP8i9laSIOa4K1WmJAR23n9Cz7J
9WVBFauxHCWzq0z6A2gaplOQpkqVKpcwo7qnqAmedXAcaoIY4TmoLaLITdzAuhLT
WhKB6E5BfSQ5a8b3T7HyOuBos710V2HXKQL6JnPLG+ZborzeqdRWzhMvVw6GPwE3
QB+oJcTAYP6Yv/B7PD+biCuoz/QXxafN9YbkDyoXit1gb1j72Ujksb/aQbv2xWFs
70dVAn3fx7xLFff50EcbfqPS1K6MZF3narQTfrBf20SPpDAencwmYKTaHxhySs7+
qtLiST0XWr6e4kz+n0d6FT/7v5vTACjV7IrHxcGNWgBALVmAXtJAVNiST/Xpwki6
mErhkwB1tKEat1nrR2KlZ/9WWhY5U9YqHzstUJvZqmpncdZlwKwh0HPeWtT+UkU9
KacdhGBIBVd8pDB2juIGnmEljQ6vvB+XuX40pL+Ekz87t34ZdYbSXwePAeoXsKsw
JXLMhBQovAIYDKlJGH0RPc7eBjMKuePbvX/+6d5TEj4iIq9fjwKCfZ2qy+JQ3gIH
cro5mLqwgO7k0Lg154v+V2zfCQQvNjqqleBLQaVfwOGRmo3sN3EQ9dzon8aGeovW
UjACqMeWEBiPyu2IoOVf2at8YaHio+ssCzSjhasa0+/6nvCRM0xoHD4azTrzBYcg
y70qQ9ZyrryRDlEEySdCePElzG8bhGL0i5aJtfRYtf9AT5genoBQcl1jO1G6hwSp
MxRSkJpRJoaa3Apk7z6RUqU30PsvQiWsePygYFIfJrMgoFTn/MOvWIxWIdd5oygx
g2TA4TvaitdWwNZneqMpWReuFRIFOBFzaSCi0HvkGzu1FPDp7OnrGgW8VI5dHCKf
U3LjFVYTD7j6/6iGKAkfhM1pQ1SV7tTRLnAZhMDYu/DgXCCuMdfJtEKM4j0zrjMO
qe0JTvgTDXmP0FE1OfYKWYC/eAavyKcnMxMrzqz+R6TR/fGGy3W4qLEO4mijfIKg
z2G9Y4EbyP19iNHAbumF5tNRHjSe0gL2p1GiklzBL5Lj3bfKySJHPS9EF6ICEvv4
+b+W3NUH9cBnyse6T9q8UVczMnOwbUtgpZ2jEUG2JlHtWuGflD6w8xliO3tjO16I
kkUA1B1SeoDvwcFs7S3rIYNw9RvJgB+YKZ+zulkBGxgGAaxBUvipkxQgqvQC3nsk
8mjeVSFBUn1QSHMuxGa9I2SzB0W7W+ugke9WiD7VAmfQna3xqPfBpBhXkXVuOAB3
xPNGUCfAxBYL4JCDCBBhHF5kl2FKmaStI3yi3F0ggx3++6nrApD4OfWm8BuEg3wG
2ZeODWKBj4B1SmoYrfDYvlFpe7NKfE4l3MYPC4eKC2SZvICCROHJOc09ZNkb1rU4
/EtYHkTZ8qgFRCUHisYRkwrXPny+4m6AbLO0vQLnVaAQH8qwI7xK5DdWKNQoJqrL
vsuAv2XCSFlBPGOoXhBQAUPV3dL3smsX2wLusbjBjlo3lB8F6tDff0KG6xiJx9CB
qws9HFSDKXXE/4i1BpAFFs58yTJRn0nCDvpkiBXB2pezXPnFNo5i1SgYlWIlOKwU
btl10omTfvnON1StZclQskancy922kZ5iFTpM53jqgRNXGLg6tOiFgYsowXcCiP6
71EwK2rSNXFdYKmYCG3kfr2QlPp81KYKP4tjgR9yH+iTKu1XjdsQO3m6DcwbkKz6
NtxAn34aMYOP39CSjmuqNlnUfk2Xvo2s+s5YrQas3FSbtFuKDLT1TI3nwVUHkPRV
bGIlbRgnRmGB2iDsh6PcrUdZpEkW0HBmqiHvwl8ilHpt7rC60P1rpuN34Jmjl/ry
5dZUcQMPE53AOAn0x82dI2lvhRUs1LbLr80ZOzgrGRpeMWzai5j6YdTDha27wlvM
biGUWABacyxjJDM41imGAsEJA4CR1vULE/Ccdv7LaIlisEucgQrkxkit5lgAIhTU
OB+PGE2Wi4ReexiIFDA65W91OCP9+1FACtKF6r8lZjR9WFchPXAQoEnR+FXp51p4
8UNPkDSzeM2L+At77+FldTWW+V+xqyGTugt5yZfYH16qBLiSiCKc8p4dGHGzrBM4
7lDqKOHyfLoGEhRRPU6oQAGgnS4BCNBMLrvtp2HQDSBnlblGaErq8rIof62YYIs1
iRqxfVKoEF81pvOsnl4U75VpyhlFB0iN4IYDUp/1WYNdxGPfciHuZpnbezuecHsX
dLondZKIulf/yo9JM6o1Tu/9AYBt1+tb9+daYy/wWqadHUDgMCNeDIjQPJ9SkDhA
WU/WInbXpy2s4uQr0ZKC6JRhaZw5ZSBZfLPLXDVHzv7hQx6jmsVyoxzpmq7M6Bpg
vbUqLV6xmp87wlk1ja+/mb89bBh/LxC3UQuhYGLLBZAeOdACREvSm/vF74CISHqZ
nnlzv6o+ZovMJIjOafXhOPayhNi8oERbLmeZeiWp3D6cnNLx1yMbzrI1EGb9l4oi
Xaqz2u+kI84wTb3MS0WwLfnea7gVGMu645CdtYK1LS59LkCv/ZKO+B2NXP9pnVPL
mjRrC6HXNZ/aAbLKkwjDbqf3GEeKINCN+ok4ZkCcwUtgoedO5ChKybx+mUAsST4L
YZRwIZk6ONXC7VcHrHDG1hEz+gIA+Pgknz2DT6PTn7MOhnuejoLUHeb+8J0NArkz
j2dhCmnxQE/GFRcubdmuNsdzJgQ827JobIwe9QDoILCi3VQOSWRmhjO4bSdxtLBy
3DJXS7YUgUvqtL07DxbyOFo13BZXAdsjSxQvO7Iz6r0+M8eG9rZIKX+EsgKETI7J
wt2+YGSHW1YCbtosQTyJYHm6AX3KASqOLBzritZaTyw5tZYuX3vCk8uVesfHSREB
n3lVBuubDk66pMNlvNrpz3zWjB9SN98kfNHuCtEpYpeGPfiduun/yZFnqc/1jF5Q
Xt4HUPtdHGVuFVDCkY7fARYqWGT6JIisLMwXs7Ie8cBwjserJlvWHDC/BtGnFMW/
9705rTqIxu5cDgByRtqZXe9iScaUL+F+c3qBf3VIVNG82WTRm91DwBn2ReMEHwmN
/t8vV0Hi44H4PejqlGL4GqvH4tQENQiBMs5rOkNiGvxfjg7F9O4dE9rN6G8qfvgn
IfPUDYtTulk0BSiIXt8/3sS6Sy6Nm8N/AGDAibABh/RhoQnhS/BSsAGo+PbVZBLr
qvRPDlt68AdLApuxDhQfPS6xGwE08BM29Y6ReIx+WwLW+YG9OX3QQHaVhEzUIHy2
dSsEl1wKrvjqYkhoEPJdShKQ7CTfzhUDQT/EpzS/xaySWJxnYFGw3EP6r0Qr6AMK
+w08ZDYBPN2Vxf8vmpB/QCW/AdjAfLqxELCCfZ7d7JYesfXm0bYkg/mAsgDxAU0H
tXNruDqbmQByHSvn6E+rLNvEAit7ZZJOXpgziZf6r++ASf3HyVnbL9FPfYx8MzuI
/qDQnWNMKNj1fBhAwBd4I7u7FENmxO3CKsZ7tMRxJ81m8ZDfE9si0sVs/oVrxwZm
A6TdYGCO586rpSti++5zuAq/H7xvLZkzq/gZO/hQPnmKSAGGTdk2gV63I4QEYZu2
fd1yV6v+lUYLGQy0hWZ4cJzbz+hReiLAjOEBys38rSfx3C5YdTmtyZ9/XKAJPsyt
zz/Y0K49E0v+oJ1xgrU5dlnb52En94RQy30FT2KrXv8k7SEBje1wgZsJVX+KyLp3
u794bxQRnx5uDBhDiax/YApIH6tdR74KwPgwbrj+Vuey4Mv46Inx0U8lTn0G1mlU
HHeM0Aue58wxeixeqEjg+Lj1RozN4inDM4WM9Lsc7hEm0b1hlSo96oTYO/yedq4Q
RhYgbokm9bmR2HR59rz2KiZ8oOZy5DcxGoF5L+zSA36RvQnPjQiErs1011i4B4L5
XsYKhpsW0Na+BypN3t3S/DZXlFOIj7uSUdX0s5myAkvCHAVHb9fU6mEmAQy271Vr
rlW/My+vK/VgM8tcrgPcP1u3Iots+RGsdn3Dmh0InkQHge9Oiriv8i1RJfKWetMt
qAYLjBzguy5BRLd4qup9kmXw1s0KCrRNcfAfKurAo71vS+UJ7M+dB7LNC7ie6i/t
JCU+dhkteqj461guX8NtBuxGNQ7VPYLayL+fcN+nNaZnQ8b5aTYLIlfI4P9FFOrI
Pv4V5oS9WFQj//B7R3oz04aUEjAtoj2S/+OV563A+HiQ8l3XkGo0z9uN5Sep/k0B
1XoZAXkb7bbg145iG2wO+Vj3Rwte5kBjtNjy3BKJ2kc78u1FTf6glNr7OnGRtw4d
hCW/pfQkvb8OLpipduEbyQMZHuILLgLQXfXIQ6i0Jsi9P+VxvPujTlaBMFqjZcIF
knmCJzlHi5L8LiWFsYZGvf6oqD0e8z68rhvTspkFfyItfhoATA9Qt7RJ8vKZaaYk
LLKHTZEIioY+RlN/uuWJ4eaWwj3vyrOHIkj7BU8dMyBacTvnWKoIH08JFsQNm8F3
kacvFJ1Gv30RqfBz2Zi6U6xM9FceGCm9HQG1HkhI98LuafgYtCrR9bLV4atcaI/x
hgzut+GVZh11olPeWHMVAJW1ttuG69ESBvMuDHkQ4xG8uc9Y4GgRFp3/Kkl03Ol2
RuQPBCmh9mVI6J58WXbfdBpTuu9rfi6fTVHAJ0l64UxttcCicMXZiYU8INoq0gcx
UXsfraqqrRY6+M/d5nKVEOY8fKsqk+ii9W7/8uLOBR1uqD+KDV1QiyXmfYmLYJDf
2jccvyRMNOmhGFHdDnlv0mTjAulXej8QCss7vSZvaX9vAzA5eGLAoZ+TwITAXXIk
POSqFgk6iB2S7KcpogfeTEh8+RbQAJe9j+fB+bXTs0FZ2FdXeFvddqhwqpAqedA3
8pIQQkXeexoJ4wqXcwt+Q/a6L0IB1mkeLyb1wqUhEM3RmoxyoDVDMgjcMYfROMK0
4PcLwmtOEmhTe3cH+WXvb3XqizCEntSzSirS4qHlpZ2uVdTKey9veZnY+wX+qpCC
hflqSlQVDI+hYJ8r2xhk9px1d3aIHUXZMSfmuUxgTn2LxEznjaGLVYToymGe2LDl
7CUfKXn6slGbQIvVRhkrFvI3yK/zeM8NBDiSMjPw/+/0oB+mijM94mMlJfxfGaXK
xhg0b5JbOIwVxhBDScQh7iA33bQBaQ6ShN4FZHZUaCas1BwQs6fbJxMLDwo9EBoR
D1/QEQ9MbV07lTBK0a1uSzx2ZVF5UGwmS2F3POW4iabb5Y60El6AMGXxvqFbMTfq
hM+/bLhJvZlLd6MSgDSpiqSCqNkl2+xE97ebkwOPx3ZdeQmkR07sPZhhK5i0TDu0
AiZOs5D+8XYS4vqb+rUaJnOEvYbeNGbW0aR5Uf+mxhNMBdTRgb9mAUvjRVM8WWwq
TR0bfmq2jbs/t6ab/2GqrHwukofIEfPIrsdpDaHFjeM5UWAez3/RCy45Ey6EvD/Y
Mc6GV2oTI37ipNzGGMuLhyUTO7OOCJq0GC8Sf/xLqTt62Z/fwtX+3rvQZEs7o2EJ
ingbmmwTNLHrbLbesv2S+8WvqSqP4Rr9fQ16NbiqWIQWPtzjogCjVUDKInK1FeBB
UouTjq0Xl+GTMxhX5f9U1wt+v18yFtRc6QJI+bd7oU0q7KA1wFqkZwK9/a2EPynu
vU0YVGEbbxf1qvoqtJrFlhWRLuQT09O+OOSShMMz8V8xmLXDw0RzAeD5r4pZVZYv
ecfZnAQATQWhFkMh7XSJkz/O/o8mhP2PzSxwnBHpA5xZjZDfWlRq4cma1XKyLQiG
8a/MRh217lNntvIX7Ve9PK9/S1RwVGjNRGZmFW6TdBVqRKa0sUwnNBgzN4JJMini
f5+yDUw1wgWyOfAGfdi3ZkydwGOU3LkYkHF0wFrsXdS9VyTIVooTKrRcGd9n10gE
5NsnCRLMNR+MLr/0wG901zY0NNrNqA9PLNw9WTyUFT6cOG7xTLCSpdhYYDvcasz4
JdFoj8ZYnfqbPcidCPgBdtpG3JuoL5roAoTUF51z/eTaGrraFGlzTQvqbLbKb0SO
HrQMKD/57INzdj+v5YE/vCxJMuUsR/9zpvORldXQrzj34qXDlRfZdzmCY1lC7rjw
4jLRUd5RYZ79i/bt1xKaApxJ7aq+Ok/Wn9H0roQdlcVrDN9pf3dkFF/Ut+8Y88lV
kFQYBV6tjJS+oSHkyH4uvW0OHAPdUflZ3b8UPAoxb6+AltMSREGMBoSEPiqpK1T8
QPxiKwCUL3iqvAReo6REhuwleJo4hiygPlNPk4i4DPluvLjNZyTIHighKfd6P0LX
RPn8Dp1SJmUviy6MfR+m7CSVAJe28ROrHKm0p6jEFrkQsa1JcJ53ZWyCBTzP48Rw
EmNBBRc/7c6oCt7opYqgDbYqV0cCvhhlGQ7SUf8EEo2n+nRsGu29fL89ErFMZ2OS
xIuZ2f1vjmy8S/e2tYZn+3onFmxLQVmR52WMbwlX8UORNQkSXARU3v1y1RaFWz/2
xcoUgvSDrNw8s84gIk/DpAiScwhAPqTPzApBB+jSDSrxyZvlfdA6j+JlRWxK65jA
Lt3dXbkoZZmc5SS1RXH2HEkksJ+X10x95ft3s68MmKqNUOJZQfakm1mooXjxCxHu
prb2ge02aKmuMdl6rnd9PjLpZMwM0yNSIwpHbeVGpth7ByKG/DLO1qm7nj9DlH3I
lGo47nvb6xoc7lbdtyLPoXa6Vg+xSFXbeFytTCvK+M+wjBYllMZQzsd3zO+V+FO0
C71BStq4EaqfBNCb8fKZmXCa8/miUX86PoJq+owxoK9UtKu8+fOgT9Dpl0S1TiPL
aiyXCMQTZVpDiM278k2yAf7HcSQQo6S2ycYjNyz6ivOIrb5F+BN+HBnFtns3GJH/
lTqSBOi7CEbMOON3RCDx8aFTWVkUWta4LtxV3YKTwJ4us+vmzeAi+QyGsy++WlvH
kmSPZIl56FgpGuTpql2pKHQuIeWpJOYAfJ8ay9178019H9dV1Wm3ZyLM2bHIQi0V
uecHGMgnE6HI9iUIXypcD3UDskWhawj2a7FzsJ9/CNtsvXm0OAef8e5+cZTpmQ2c
KCTD+gtog5CXlNlfbFYgDdmrVvXaEGRghr/D/5p1Q3YIlKb2PgcyQIukHKjmaMUf
n93bkHlGTIPXrDDkyiyBUami2JcVdC7c5balnoNVN3BP1rh2E9OyzwWnUZsY02Fl
d6Z9+UzlNIv6wj9Q+4dmYcu4bOTblROqD9f68LD4ZsrV9vu449SHy9nGG3JJ6e4F
q1sDqcOBGNRQDrQBnBN/+fPi/xZmi+2wM7cZcnN4ji13T4cTNTR3lbc0DHK1c7oh
oDW7EFhcpKBfE+qLrPQCIEbbzLUt5FiffA52upvzmsSYrOYV8jM01FhHC5psozkH
59F5BtDI47V/PPMQAE3XrEbSnSJxKCvWmdUykn9FGhMmiDhhQOlP1maUHm7sQeht
G5Fdf/GCPLQNQXmT+e22Xwhe6D14sgoxFeYIQhTF8kPyYvVwLdp3YRRVIKuQq4Aj
9akPM/wsKnqv4AZzmXj0FJAUXxrnh0fQnO+6fV51X56ewFfRMJ/kID13NA17fx3N
xuvzktO3hTv0Ptp3IxBJVVZHcPzC3okLfwJIq0wTflnoo8E9oriv4P0f+NqNaDuW
F9by3WoQkbNzakktqRSGH6OuVi9GZ4R3/Vm9FDhNvXRbzBStTmXNi47Epoo5Y0Yb
jQUVgXJlqMNyaLVAt9UX+FZ4rnCW1ex+457ff/A6WKSZmisaITal/84vxlVW16Gb
RCAzx0kT53+pNwNvyeFGHg9Zd/nAUVEFSYNSNL+ZFHITCqLrHPF/TwYMdRp6rGqY
JtG7E5vDI91y/PAH/b2QOoXcahNSYUg3FWt0QaoXKWhBdiy4wnaJq33M0ZJl5+qf
CxnEv8hcY1imjNhuChp4VGhdKDYAwKAAU8EINjczvygKFpptGEaWD4UusdkkgSUR
ahSgjuBD26PTb1Ntfgvg3L0VgelXVon5rgkDxsmLImxYWxaPBeRHc5ih5GFv0Cn1
Vc7MvBmQWKI9a/HS9rpWWx1OihPKU5C4DqHHHXkYaMfW57bAZCGSePlv4IzUQaiL
4PmyuYOr8LxjO0MBc2CB5dQSyR5oUdMHq8qHXCfLD/1GvDI+Hsnpg9z1eFHpEQeV
kXIQ84FpKQevCBmOlV+6f9XjfPJLi2tp58bkSHTgm20RN19jjtpuq8928JM4WwKp
wjJxHDNuiNX5KSpHviDJS3p8H3mSIatNB4hpPH8KL8zNONsMI+DF4zKacqhJ6AIO
mfbd+nWFsdenHk85kCW5w2wJ6yk1AKnq5eCiBWyCtG3W75CuT7FWbXa5XuAzOARr
A58EVkTzMqdaY6JfNw36Y9Zvv3InnPh6AQcaDqzaUk+Ly4jvkI7tsWt1U6leM2qS
cyKgLqxplVuvKwLIHLlaXCMFSEyvgycMahdv5fIq9l9gPCzhWJdcngKWDgKIokFj
Ywy3p1rMnpYSeKGFCwZCYeD5skUJO4WyByWyHY4QkSr9CulnOQk4Ttz12kPlV8Yr
n0glXL7OWpdRXe0V0sNaJ1hfdfFiOZDcLTndiuUJ17dMaPA9CCjuGWhkfLEiAgNt
ZbQWQla69jkYU332AL627xlEE3Ancy9P3PnmHUgln4Qx0leXFdSUd+1MCG/bKFE1
Uv8TXpM1twGOeJzQhtfKA0kGKKUHbtgPtyg8cZiidCxW3pSU/1iHllGxS4K11a1N
qP2R9KFy+Vv5hCbrGAxf9QzcaIoRGERzUhAnrQiS1zO4zb7yVUemd0G8OT01FNTp
by907tvhjne/yWXGVScxeT+kcRwDHz7mr+aBw2pqRnbtxHmYpJb0BbA4RlmQfhMA
YOqvUERI8vagQ03mmg8M6oib3tFOuhsFHGSC4qlcR4xgvGnj4V4wcxdFYCOjqr/C
J1QFDypseOrF78TTLsyqdca52kANd4HgmBLQQWuhNjKTGAa1765THPunr3yYI4aG
MeUFCdXLB/AeR4zZC7dk7Ig7fLim0QNwdFSypxAQKCCOtnd4wGL9Pe2hx89vXNp6
OJXKMXe3LOnYjOmj8lEq9DpE7FkcCqf0N32qK+cmJP0y7VNacVSNupA+gTyFo3Gi
5dyXj3X6e+DSSyAxHwnNO6dQGFA8af7sE63Owv5lxHmPJyDDzGx4fY1kwTTMfpMf
0HW7tk5s4HOtkOGIUqc8T1grJUdrDa/AXVTOORKdFpuUM1LHp1f0E58bVoJlwt1X
G7m+YHtPXBl05Jt6jFaXVFX714v0ZarfeGFxaSQ8jmkuW9VCE63hfgnlEkpbAJ08
mcTLGKJgF1XrUrOSGI1xDr3bGogTeRKnpepRcnvh+Xxsod9j/R/MEzUvZKNSjNmp
gnCvRAHpFMtrXL+2aaYS+iIFFkYpihwnXLTnyITQ1F3G6Qvb4iQtUJcrnh6Gje4j
PFKumKsXIaQ3EljnZoSluRZykPuktwF1afJPWe0n+Nn7yuvk/iJKFMA6basLQ9oF
JzRo+8vEnA3KQ4IKQdGvUQS97gkkrUYq56K04mNPJEcEMIMoXQRJ/hR8Utsn0wO4
TzUA+EQRkspWxEv+7L2ClsGpTC5hVKgAm4wICaZI6ZawlPpZpekSICv0aX4aTWkZ
gsobORXB/qsPiXtaSVYsfV6Okhq63l6zJ8dAU5vtDWWihniOCobk1ekMjAgUeDBm
OrFfXl4WYmxC73j+o7SiL1x3f+iUBsSy5PhTGD4t2BWHkJbhsxGlKXamV4673GQq
W9lhE47A3ZRm7Zjt2WHUYAHNQgGbk7ajaQbOXB0dKdCMAhlNtFwdYWdLKyElEN0V
ZC5xtcqN09BzlaQDM1lmH/LMP8AiWA1LzRHh9lTjba5Lj+1J/ij6UeHbaFe0oBm+
FKGrKmaE+HzJ0bAH3M545jtZzyP/gXsMdEgnBDPk8iCc6Wito2BaGxmWfJyLQnlT
GNpU2OGHSC0j5z77+FkAXEFQbBDnK8q+CX44Kgl6O8c3gsG9mxN2vega+z8wdjI6
fv7DifMTSxGJTsqq+nnjXfF97RJNt85p5Aw+BMUme738bv1QTiMyfZXp7B4WsDG6
AnSGcQ8UDfvBCAbwL4mlwW2N1h3V4jp1yyUkfxpd0M6tRJL0qVQWc67uT5io4XuG
pkCVr/ACbpEBrKihP/vx9SACbqIWtmlJaG/Nz0BLa2XdQ5/HiSw3XMVfjbTzM7YM
BuQVkkx0ZP08Z74FPfMuJ7ebmCjRa3BhwS9gKteHxwlpRhY0r194EunkpaQ9gFbB
fGwsz6xqFtuSTqa0q8VOqwwzpjcDyRxjzFrGO+6RYX0pJAD1aFW4zMnlvBSG+sPS
eMD6B9Mbpzr8P3TEweWnA5sRt+PK7UeOqbpXrgXhXj3RMcBz8v0jVFYfWN+VW3vd
Kj96iH/Fc+Dhm7xiOv6J+so/hbqo8U1FkC8Ti/UAB4FZyiCbcT4KMY4yS2aAtkjN
nBHlx9d6TYQ0SY7Pu+BVpXBJXlaavgSs75XyBROkR9DU16UCkA6GX0kNPEke8A8r
5kCnWgYUJs6BAZtzxNu35C7V9uJVB/3Rp9w38tm18KZlQb3mVTxRsF3KIcaiZBeg
r/9mA3N6Mk/gHynLR60dfmmZuLqgkhhineOT64vb9dJmXK15ngKsa/wihKnsSykt
cZlwiJN3FNcglQV6zy5CVasr4N0vTLcMOhHcEjI5IRwXe6C+QStfyDzUiDMyrPIt
Jyg1ribqWpktY2HdK4GnSAGHZeVNWuO3l+BM9zcQ2XcMFnVmnScp207vhkY2vUp3
BkYU9i6D6g7hkZWByYwZDTJyjLLSW42pzTm9sy/Dx8pL3gTmij1f2AD4dcA5mcl4
cCpjqbJG3WNdYzbToZYSQGR4oDtj2fr1JuIuTDzEYI+TPl8ct0QBI8wj3uh2jsrQ
bxUidWXG9KVn7hulGHkivz6qJ4v0qYGdPsK4VLndNvlPsNJmlhwfVHqFlRVAHeKU
aOCVk+Ad7ILm0sXvh7E1lbNbXbZinnMvxAE85EaeL+pZmu/aJhkaRibiTjj5LpW1
nyLeYAW55pL6TUpS8DgJR3pJH0OjzN4GTTgFwHCSMP256/jw0s2yiNspYds393Cd
1z5VpVPq1li7QiURsKV5BlOWp/c30sG2y71USfQwurR37ks3jKjAqR6NsMCHgye8
YAHf6asfI2z+vsjAtlB0tS7gGJcUx2hkTeeciuTGAoWyVd/LYz/PEdJ4HtNInyRB
YpwB9VQEm01PvPVCGhVA+4Sq/ab102cxb0SxzXcOmofU/xqvUnvt6TqDmp4smP1D
o/Vay9mUHgKcD9o05D9dLRtM4iEsyVzmoXGXGoloT37hl4ypWgDWB09YLQHpo6aR
qTDLQkUujN0uOlOb528Jw7TbycvrsiK2uSFZxLiAz23phK7nZyranLgg9vv6nzRi
CJ2QYnu//C6C9IvrtErhLQo5wchQx24yORAqJURhEj2R5W5cVnxrkp99iBMJg66h
tw5fqe35ZN4lAq1TchxLv4NX0OLXg9FWYs07m21ibbFxb3TaAqZt6uZ6ZVj0+i8P
cKQWiuClYeJC1r969u7mHleszb4fnsa12US6EhbQlt7CuQL8c7qDOPN6DtX/vZaL
t9g5RvXmGmyvOFkmJDX+zWMa934aOb14NeRbdIsfiAEFHZCTmZHjjDFUlEJQ9Tsq
+9zuWWyjaH0yD6AC5F+/aXow6BhuFAFSOt80Puca8yQM3c7z3Nt+fzLxCvvmD18q
JHFgy0bv1Qjz+CQHtQG66rcb0To4Vx4liaAk8JxQmj3S3bhi/wVei6pDPRX3WeBx
0po7jJWOB9IIh+4GuRnZ4fCCg8SoLhS0VOrznBQouWuT+efgBFNGMPGpx0BqOlKS
9/SbtmlRneqAZHqQc0rbu1rraZs061niup9g9bhFA9mrDsWWIfjYOba5yMB3G53h
lJXziT2fAET5rNtdL4QsUoN4EujpR2NNElfs96iKyXLPn/4ghDHA01Olv26GGU1g
I/zuBEaPuIAihsxGFKXA7XACYCMxfE2OY/oiIxISIUM0QJXmjrU0qvdKftJzhP2y
S6jkDHtjP66mxRUW48SHYy+7hHNeBDEFs2dScyC6vBIJpKZdsH/7p6SG2eFQEmyh
lfgp7JwBrxk7Lyv1dgYPmDNNEMD99hZazWzlKqdQFlv/nIz6bIv6csi2PMkbUYiM
rzcAmS38taZK/m0HSXX2DtGYAcdyyyGKaqkerrGWdrwQyIqUSOdZNK88/Qvrqtt8
aW493slXOPrnM0fkE2dIpYDyxenZcEZAyju8zuphZkzhe0NNOFRb1sOMYMyEIcaP
C96QLoa5xcxwEbDozvGerhENNs/ckLnXkCu22nGTFfCGy92XL5YUdZOu0dNN6w1o
qDo7V7aNoYAhZ0Vovm40BV/f/ctlHGd6bOOWhtVPjVN4Er3DgPi6fBOakZxUIAJA
q6SmJKrBV9sI24IhAOuNq8i1zYyJI0dcBcK8GswJ0b7tQh9RpLdIAlnjH3i00kbq
OhuEfHBSvfuf9nkxTIvSIWT4Y1VaSKWh6OFPG3S9ThggYUEV9DN835HsNxrC+BNI
GUqowKZ/lsLT57ZhmkX++jW/bqtVLX5lWg2ftgtArHaODn5IrwYU3YoFhX0zeBEf
p7OtcCviHo/7FuYdz1eqZj92XAMywQZvjKsWVpQu0JkQB9Flap9QtOspt/ne3051
Zo6t89qXdzXineF4pWU9O/cg8e0EPpLAEeiuDPItT7p5vcrhPZRq19barnLzoZsv
q1h6wpNwai8tm/xsrkfpiQCOArJ07PyYekcAabgVvhIR4fvITGA5s4panSwUJ37E
+SufuZcZgpbQU/aU9RSYY+4Jt5psoZxx8X9UEAkCsJuMDPWl1k9LNGk1qZkZOjl/
dTedOXCYQMvEhJ+I0x3CEjlO5+cuEf4f2DVMsA3C59c8lKy00wH0C2MV4udPK25B
fARBWAaf8fgzB238AeeatUou2Z3uGiiP5hhBWNFCFUCf+IeTsKU5u2Ty2p++sIPW
TQF1XYYmOLWDmjzdHvjy61IUMFRrSWDaZHLyVGKPDHOo04N5RjZlgDeW1KgoDsA8
rGBXoEojSqXAMKrfyXwgz2FIS7mFcl/EZrXH3QkFQmOHsM/yRUzBhOo3J0euZ2Bt
Xj0+M+agDwGf/b0/qAQXezlCW3sVLT/LSAWtpbzzobfev0rQBrF0S6ue+c9HWNTk
A+WoW96LUEJI0zUuqD0mNKgf6rKqF2zJW51SNS71tJR3XF1aTqwbheiKQmg2zHVc
VTjVrL+xa4fO5aJpd8811bM4+cGzz/n4ntkEfQOGrgLnkssOCCQgKaa6hzOUVpTZ
FBqBGFKQfCEgAJum8pV28FDIEBIbQZn0Q8LUEBEXb2zIztZTruTP60mFEBIcP+De
hb1msHxsCp19cXYPCwbTjd8JlpjTgFJqa1CPUxapD/s4mZ0ohFQ7Vwvil3YoI91U
+m4aOOczqU+FdWc/YlKqf0aqocCvmFa316HYpEbbgkEat3YsUv/oY+Gv7p7g21rN
l+qxqEuATo6uhYtTtsnkbpj/KJaD1uaBVrGbcq+0Gmkd8ytGWFlQUzvZwVRc+/5l
EJP8Q7bTnoXQBwVVEf/wd/7UnxTsvQQ11A8apB2VNn+wT+/F3W8nHWATxWWQkyt8
VT/+TgHa3SodYMXOkOT12/ndtE9417PcUcvU65n+E7JKXQmFiqWegeXVXgXeAa2e
xvAeV2dWaLqBYx+4zujut6bm/yPN99bfQNiisOz0JyPueqH1dZDRFLa4cOYf6DfO
xfzBUa0MfMR9pd0oD2jVqydDI20obzA+djJM0hQ6DW0v08WGBGcpMNJfdt+LfMtW
YJEF8VNYT/LVMsS3ULLnatuylRB6MIog9JfGjQ0ljoJ9mjUbyT8ezTyowsR4/k+9
8QYvQN0Sn//y84ELZXissoKBydzsMOe3yKvD+YzPOniCz16QVpZou54PlGPgQrcQ
qOjszskENBYYFj5qrpdxzFPUlDWQh26RiFleIPiq3QjcHL3gW0EipcVTHkwlEGhN
s/bUVzU89OEq4U2GnsX98IoFASo+Xg/5l4ibyDzMl6waeJXnypboNov/Ktz329Tu
wSBWkouMZ/yw+idDejjH1xnVQmnrP96XMpDSuOvK8VtE41gPMZX7Ftf0uqFD/NgC
71gKISoFT4r4G4Ef4Wp530Zf+/x7QUL0o8twVyKmZKYjUr+t5XL24TAhowHsKK7M
DvZKG7hxP0XfDbSjIkaucmWGIQyIexPG2VMRVJtHOsbrGw5w8BVf27QTaOR38ZBJ
5Io5eEhE9pT2JNARr3msWroWTxMC0ZKlRpvpKhNWlReNf8lIUZc3sTAzZUVPn+1H
9mHT67ni4DtCVNMdHoEbyos8Nll+U25ceGmT3NJhAJYptsGLJmAy4whR39mLqsqd
UqwANPAMRT44RUNpLBO+ygCERsQ05Hw8lXP4gCRs49Kr5HVMf8Y26TRk5nKBsGoe
kJ90CYnvX5wpyMhtas5d9/DxbWgu30ImBe7QiSU6LpG5np7r61LxurnbHqSen6V6
/nGsUDSMPvJCFSvq3gpIMIMD0qRQOEsys8vPhdCnbyBDRxfILkwOaThFlZbOC5l4
aVvGhGasNnuBTwaURftbC9gkWxuEUlSZ3cDP1yk+Hi9FtWhkIAh9RHietgBa+Fpg
ALMai5EukVXSgBKeCWd0rVuVnWORlalDowmOlWGhQxfhBNUnL5UtPM37yr3VP1/g
F1mJsqM3wiw/evwDT0EOdtG44NvQy3r8/h5l+gHpa8lB2tDmxJEWQ9UAE8g3fRaV
V59yAfCDxWBsayadvAt0kZK6/ZB2cEzhr9JZ1cAmLGoeZLI8ebG69djAUsd3uxRK
8wMkJh1ILBu+KL8j7bpEZo6L93jrdqpkP7PZ9mOSOkHczxun813miKDR5I7mXohY
kYYrR6C/3UP7XYz7fkBBh6+iC7qmrK37eVC/u8poyws+OWnH3yL9zKD1Yky0EDVl
6Fr/rr7gBE3U7Zw96X1IxEPKYmHjnYMADeuOS4yaeR8j5zs2eK5dY1iDm34QI+/j
qHd93VaK8I3iic4I1wXIueUdM3ONMVdi7IvGVc2GcDTHQi9Z285AYYsyAVusTBM2
NSa35IacyDVdb2on7Z8YW3zr3UQxgiP/nUOF0CTzpxOGMGt1iCnzoVh/4VarAW7z
pNDdZfGMkbl4aPBKNBBWIJHFkzSEzJhKZGpUHnF4JoNLhzKd/VsVrlbRhMJ+czuz
qxrdzkJGU3TO6KgDgtz6tcUmirk1xdpnrpt79MZ3bNQL9AUz14K2P5a172Wlqit/
m+8mfIzwJ1AWWo+SMFB9eGLSMdytTSIW8k8aN6Oz5T1BRHZRXfyhy2SGv1LYlJeO
gdnyk/mkN1me8T/CjaCGQXsb57NmWzCWvontLG/o3XtCPi6XjDTQ9L83NZDuxyfN
kXi2OgHdNPCx+VSiwsBvt3Pth5DL4jye8vi7jUZKBn8V1/qb20FSl+9GRu6Nz18d
bJvUmsy1k5QC3rpas8TIU4M4O44OOe2u492tOYQ4LEcr7lozVBbXwT2oTSdyVHkM
FMPWKpXpO2JrR2gY4lI9riY88yU37NtaobRUPb0B86iqu/JcibuvoFcWtAFzNp9i
rrI1E/7DsNgctHiX4d00nUPXIV6c6OzstWXoEqW5jrtcUo7C1Zwqk+afDXzEvT59
2p9HHTmgzgKV+l0JqrPj9sbX5+SioQEWJqr+FnsyJpsxWaii5A74jiB7/iE0ycu3
uvplA2NDofrJksfl42seDEFM5Jrj0yDCNapLHOoCV+HrgnniL8sknQJKxsDuVWkQ
DTMHBXtFse8paQp+WC+4l+o3pBO6f8nQUcT01/NDdQOhDtTN/iNYJ0COWUZw/lTg
ceSAdHhEsRVAYLvC9T7+L4ACzuMlQQUO/3P/zs+wDDBMRHTmri8ljxHrc3IJRHF7
/l9geIZBpRlXm8oeYXnqqFmMQy3L8oBxxfNwDztMjtAP8y0kfGD/gibRbtxoJVqX
aqAqXTvyMso/+RtKwLlvbViSWJ2OZb5C8fvENiIRjNwkzK8QmS2grfzeSSm60DGL
7sxaxb1K0fdymKQRBHzg1qXqRzpgjSDsUqkVh+FyOagovo9n6uxr3PMOmFoDKN/Y
Lvxk33LN7qx6hB7QzHEvxluXVDmci/yJGUkYPfYbaTuP1+sF+/AU5ZtR+zhpwRPg
x9tXYsY32TaVlgpmRT/Gx1dwcRg6Z/GOVpqbm/7YKjM6Ts6bqxoYHnXWBWxLy7a6
NZ1WOATmnbMSLOFXfh5Il37jPnz7ILRF+emG4NRK5/VD4WHg3T0xJSu/W9lNl4/m
brgMZZRi6GAt6l4YsYjUiVyUpLndyB/LPzrBT5tFV4fLNreuQjnb5xJ3yD9UnkT0
+psnkIiwktMaI2uv8wbEdSKFaqL9doRXZGUU+PCNbmgsvFC/4Ro8qWspwDKZDRvO
+KxcmSoNkUnGvWQmHe+Y9J/yuqpTKFK61OCeKM5b+GPsvQnOvJL3uyVzWkjZNn5y
Yh1Z3Vwi0UCHmtWZb3oIcIOnNVdBnhAgYyMU7esnLZlae+yhXE9ao2Pn/Rk6+D8T
8/Yw/ePorQeurxWE+hlr4PLC0lr3TvQYR7iEhkF56sKuKN4uddT+5DfKCSS7gHVd
a+wPFLLF/5wvLGpLMSdUSQ4VLUuCDFaOxeOrHpDj4IMLVowMjpvzxhSV5ZTCd/l7
7lmEzVAKnUjstveBoVhQs977TcwI7aPkfOcnKaEajnMDweuLvz4AZiYSEvp4e5xF
+KZjcMfdjDd8Uc2yknX079ShmiZ1roFCLLWdNM7Urn2EXHglvLLXDCRzWUmcGSdk
pj+xFgYFlT9paigXo8qPBmWrqKOQKQDK45JPu5mMITIldfL2XC81Jt3vqNKdV5Sk
j1CpK4R9UZgobHToymoHIPBti9PEgIY44GyOxH4U20eVmHH2BYRFSvX+gzMc4MD7
D0HnOU5duFfKWEseSOlrcuKsKDrucgyi19nYop0xV3qc6PL+SJJf/05kpazvdu1r
J3Q1nQC5EGCnjr8qFEMfRrgEVgceQMddmSvmv68eTqA4Wc9INpzqiL0Usn7dLucN
LceevvFmP4E1CVJVasQIBWuZLCr4NVDruaUW6tXH4c3lLQwgvwQbikPnatcq81/R
ckWaNEB3jUhIfjz/gfzImJHRdo3FTx1Q+r2v0Ab2eCGSQQ66lM7QJo7YJRL2f2yQ
yCd+b6lynX8NRzSusOkdFp5sBs1TTFf5QrysqgiUY5YJTkKL6yT0MG9UneVHjWUZ
EkPF3ApdIFXccYyke2hDWc8Q7y91Ejn5c671aY393fPTifx0tkhmL6phjzyhQOYJ
jEl+UKhz4m0adhqIlYPXlGBDmPUIWo4ldANg9ZQLNBt6NIygTe/J6qpa9E0rB3Bx
8r7JqUW4foh94px7nh1ydwfiz2/dS0Iy8IctI50qT/cV0Jiw+jrkhgLYvxndRkfI
VIz/dosuvgb86NG/RsOkZycUbFd+nj1rTl112fXUp6sSQtphmRSjuPgqiFaa6vKl
6Ye1MeJMz+9T0qzxY0VVhJXKO8PUAeH0ykDTn2Fndv6FmZqJTwbRT/c8Fd5h+jSE
Ra5JDfKVHGtpQsSRvEJ91SBHMGtTwW8KtSnnBiWI/JT1MK6rgRDhYNKPuuVzOLu2
aj9y130yvzYsVVfGfE4uZcjLvow3pimC/Aiklsbhf5zM4dqZLwWMyZ1dRf4lT9HU
AjKArhKDxeYZRYET95j/vvPYPbS5pg4ZteSXo/g4WXbCttV81aqJtu5pyJCuts3E
BUona7lS29slXknLQvxqvhg76X2OaQrh+kQdAAZVD7M47UVwz1sVu1atxSa78tYS
2xMhAJgKodInbWzTkQ6hArFdOy3tPdmykFTzEyLOj/StkqMAI9qL0G8K0xEgrzKw
czW3xWAneL6WlNpy4GlZdTewB/NKsVKNm+HXcSZ1kHS+vi2I6wBKlwngUMW31Pro
fpYh17pVPPfUFjr1vUq0fZYfYlRTYVND+necWiu2rh59Ez8h1TgICcMFjI0YRnAb
toRdzziXKlxtxS48rFC2sDQoBGSbT8nD7HXgQFxwtAlFUP8hkpi/bpKXgHl5f/yQ
xN3cq8rLrfLKbGm10nO0fjPoayH62YS4Qq+WEQosyynYkI+Y7Fvr7Mn7nzqVeg8y
qnxPOB12qW1IkwliLpuVN5nncM5ymHDbbDpc+AodWp0HhSvUtTBrJ9/TXmAPwKm1
KfDqn/9H72E8hQtJc95eoBjjgEx56Pkat2YDzVdEBA4SsxIggdesTCUI59MJAmyT
etwbqSUISJPlrfY8vK6JWXHGBYfmk5vRW569XWR4E3Hd5tT2UIu+PMX0JwhDBkS0
aWp8lu0gxGyinNH1Vfc+uswmexUie0p7Uj084NZ9oTPs5EIggM4JpZ2YyHMRaN43
woPc1hweGbiJENnCSrToWiNvaY2rwbJDmZ9ENJiZFzmZ8XcIso44g3jc0bVh8tPu
F2LCkXbg8PhhJA+c3HaLesNn+Ofm0c8nIkJeRj7PDObitnLothf/p2iRmXniBFF+
EilLrdGn73sawoGeyJgKHiGEuSHzabAZliM8tl1LHqjEHVrjoND00LBdWuIQUBJ1
3D0u1pl/ofIlKcgj2ppMVqHqLe3d4khZ0B4oGtxHYMzOUjerzE2QxQiRAFQ7ZdH6
6kfRo6wSdN8muLMSN9+83o+pAOUN5PtkAjkLbDgvxYEn1gfJY9gqPpjocjZHpcJ5
UP02RgwhNu3LkC6jnMnJcNkpSgC4zRiR3/3/i9isHL+pHKnAfzDElDg4Pkn4cJVb
4GXJIaiXrWPmZgOsCFLPeZBhJwnJOW5PuB0tpYYkuKvcI4XGYGCKr8xXRUMC3msD
bpqrf8dUq9g9iPSgFkVbHsqAPGXNfNYoa8MSS+qK6XasFxNioKc9YuYJKHzNMzKU
U/Wbc0VHLY3yg0O2EL7BY8LZy/uNdowZr6AWui0V6ekP9Mirng1dOkqs2rRsTFvw
hjcS9fTiMhJLTNdkzlXBDKdSLBZcdbjgCXZVYg1QofY61tloWi6EGztIdcqLU9qG
yf54tjIozve3LiC/1tokS32cfG6FKdG9zOpoEKffNHT8yez1D6OTyrSY4C0Q4w+O
1XuhvlKGc/jZslOgrsSntwteKfvdcfoBevzdnhCyJ40gcnygMCPPW5yXsxEUyt4r
3UW9rMs9u4lPc5gsGbKkboJiouJhfTWV5lpGuNoApuiPSkUgivuEHr4Ha3GVkeGN
hkTHRTZyKMn4UguwSkRVflGBUCAHSGIbB0JRP9JiSXohBZjl6+N+RxpXUdhnhEF6
1PgpU94tXavFk9MjC/akxh0H6Rnkgsr20RPONGMlnRNhqztg8lz6Vleazjt5K6FM
jOmUF0QkWKhCrNa1OXcTccFUDsrb+k/iSGkW//SvV838rDIE4ExvQLHtUIjGGZV/
626UYiv9F6S3UIGTamdyWkFpoNAzeszLL/pUavqCyi3onJb5tcd7TKeqwdJBGF36
zxF6mPBUTmAa0YlEytPE+QBgzXGj4xVdWl2YMCc+rzX59OxiXI6tCXuJMveERJhb
Go6ICXbq0uf4BUfqwXdbyitp2ZAC3uuPCiSazc0cERe8tCakrUiMOOv5oCksOh7b
z9eLa3EzFmjGUgMhcTpg4vW55Cpu8POwXMCiQcVyWjuaYV6r3Y/umFTVoxekrF81
5AMWsfe4ihyWpXhE5cDPbNL9PDbJFNx9lJlnSL/eTfhClKnP5hX9s2yoidCETwnY
Fm8Angracg2EPlQoMwjYbjuutVHxwFoo8CWvQU4lBDoEjhg4/bSpc432HO3opMRg
T5bxiKPH+4qaYqqS2Di+2W3dEc6qUCqcOBNtKlExVjewAnragqZCMKQKGRmgu4hr
1iq8Byo/SPvOgA5zl6V/xE1mRB1Igwq7BljB1jPwD4MAHWnl6684RPOlmykAH+75
aCtq7z8B2L8SNPGVNISMId+0p/KDCtENm3sNkXmiYfOS0sDAQ01Wc+758l5r/H8F
E02RXQ4hqp3JhSPTdSdQrVaPj1cE1lSuq/wOlq5FV4RvQYsrYMgMaxZot3UfOMbQ
OD8Wu6aGWvpXS2HlcLEDMegcxTMF4EOQugrDE2WR9C+II9lkWVWYixWt6JfBRy6k
2T0XalMxuHcUYdZYwp0fRpjR+nMzvfcX+BeYIE46uTwCwENuNugkhpZHb/+yBAJh
yMPM9L0DVXXvPZYO8KhTc5x8/M5nA70xfP3BCbw1BFO0gn0rXHViPk2wJzgX/MnX
j6icMWj4tbcObA257kGdlURDxncz8Py+Rw+eUm8eKYxq4BzY2u/kwb/21s5FOuQi
l5KEs8p1USd2jGHq8ees77qi4NhF8rN+RtWZsUi2GfP+k11WYvPtEiSNz6OJHWSF
GKLf0upEOW3/MkNKv/Aub0NXcVJhnwKD8o+7Hf/QXUASl3qQXFtzPQzbrBHDSCyi
XiPaKfycL0kUA0CmR+4+TOu36llxTw6Q8GZzNIJBqUIBM+dnRJNsbIODlXf2XgyZ
ofHwys5F8FKbK1M1vXA/rBcz6HOt4EhaiM8en/UUjgY+HJuX75kT4c2ZHRdpdpqA
NJ85EWUFF15TldH8MfCUK2/4eGzm3rCMVLpeQTNcz2W+8HCZEhGthxO3d1opbVUO
fjGSRoi33+EECOUXXMSWg4TR08VF4e9Il0LK5s/F9RDAZicwZmCqGmI9ZjcMeqAJ
bU4vn96BcapB17m8hBvpH346fiIFgm7EQbsibVwIguceeYd+UY1fCg6Lm02VXKjM
cqbgbRmzk4a0mYD/WKZQr8ACTJsO0sW6TvnO/aESfpko79BwNNtLQtbqR+EDkE7w
ptVLl9QcHnreQd9oOFPPlAvij1c72gF3mkQGcOQPktj+PawLhBze09UAEJet4pwE
7wpCNvhzQqUQhY+UNlNR3njfZblsYNQClyDpg/FFAvrcRXNXiP3xSldEOx3BdDU4
0nw+1XKvPBXSE3b5Z24kds0A7RQ/783e7yssSmgJcEXAI0fG4AvKRZJQVMRWLUsZ
Jqfbb4aNdnFlaWzdEydNYFUI0C+Js//5FfXwktYv0Z1WC3OiyMXgo4w8BkmMzPYp
LjXoajqpNfWJFaBVgyUCnB7OepLN7bpGbndvTLQD6rr6rrsOBBlfeR5N3u608fud
GjVuuE0gvL3ZAsiVXbST/mK8Z5oZW95Bb2EMeyXpuZltr+jSypAlVqghUK+FNIHO
H9bgczgA+HYMfp62Hjm3NlIMha87fQb4scx7JImmu9xoqo2wNWsshMXpKLiahO7a
RTTecYoyoZ/ZPOY8ZPaf14BeQTIZmUdSncaKjq5WvDF0QZZM8jy9gIKwsKLci+i5
UXVnrWOkL/mbuFNrfc2a3ul2/kRB/dlmNBRnJOFWE3ca8BNOmffrjF1hEUtgrJSz
Cd1xx4twMrXK9n7Y3i7Q3saidBFPdchP3V2+Xx1SKAekMF0TtSjX3jEmHf2jUSPY
0cfjdLRaCHNNllXGcwLLBpegWFKgqZGTGarVfp9LswMBTfbdLHDg44CPLAfJRBFF
fWgk5S3cDzvSMBpFewV4qUq4yLuSxuzDm5U0kUhXXZzkwvuDF0hOis1a33B53Te1
4Pr7TFkWjFuggL4ZIRTNhC2fDPQI34AFR6G4JAkgb4x4wgMEFHPg+HjqgG9RNAjt
huBSltMX37y7hy77tj7uHOBYbhInADrlQqfT3MOVghalKsoNqST4YUvLKlMr74xx
ZhiUDXop9+kaI3TUWwFWHCo2VFCiHayhTp1/6pRQBI35KDhQouLj6H5Y3MUzxsQZ
YCYvLS53QHxApUOJl1rCtY/NJoDk8tfy2v7vtaai5x4ZYg867GB4kNsYcvZ8P0L4
OmTOCdLVS2gbLpTSCu1xHnYwEltIJqjV0kAX2ygXz9Dt74Lh2LcNAkgXwPVH1NXP
PpSsE25nTmylgGbVsAwl5lBMJ6hxAHHiOPGgv5oRvwkHHYGVlSksjOnJFXA/Munn
RlF9pZnYvwVBuMIi8bduir7jTtL1jxTlilOoAPGiPDqgUxigkdvVWcf71i4B5cOz
L8dZTXmcsEA95ZkASqDKW0pfvOsS6f45LeuCf6OLVTkNz+AmW0vJImiEfRtYBAPI
x3nwixmUE4G2WpB4DWqnTHaWxqsKAqusL1XzejMD0ydHGl0HJVC7PTWJeiVzmQ8U
lV0sM+Zrne9/dZ/vdYnYsMw0XNfD9sSejrBrW8kDmNRiYB7UjH/HMlLGiEZI5cr+
aOju0IHvId6B64gahO/vT00nx9til6y5/Wc/F1u7DwA6Em9TfbGc7ocs0Vf989C+
9kcBCxbEvrYpreXroXheXgbn0Xhc7lc4ju/Fh6MX+hJml7h3hgXVZIDH4HY/6z7f
A/x4iacjo7qOE2FYNl2zjeEHP0TEapq/+2thGezLhLotUdI7HQsB+AeJY4W1dtbt
f4b/d8Rrxf1JR8JZkVMTRvcG8YVp6oUsurL/XhpZmEv2CHbZxEejdSiOcPzwST6M
Y7pQYISrWxXBPh4yem0A1T9nnMLBmX5AZIiwL7Nk5I4feznpafTclt99M+L9CcfX
Ao7ju/ez1L89tj9dLQowU6EM09U9bx3IUZ2p3cqlBggKiGsN/TjnXRsLx80Xgqjm
VvdC1hf1v0zkZ19TlUYUO6v04gpnNVJ+9+KVz9oKLIDNnSpIpUxnr1cE1T37tuDB
HVoPJ5WOXgaDOinW2JzDEAvPaf8UoAr3b5/Pd7bWI3Inele3RRSB31AZj99yck+w
2JnX8CJtqaZpEULxqHQrUomfkM2R7ljUH5FLSDzZ1NZnmrXJ3nMbWS5zpPZNfMoE
E8MVsG4FFgHsKAQyfo84naVbdul2c0lhTro+jW+yzXbbXXLkeSeby5GP192AkJfa
H8xo5QmBavE3oPz84jlEqNFipr8tkStyjuTuAVABdPBFtWDwo+8fK2O7tGXgkez0
gOzFlUEDWZqHKQOMgQtRS5zPcu58tXjZkob1i8B/RmQIrhB+my+thtTlJ5qABL34
MKx7hjK4OGVd/LF6HwrhijkKTEwG81An3iXxn58OfNSm0ZH9XVNZH1ZLjx89RkSc
G9OoRl6tCeE285n+ezolsfgEVrR4lQoHY53m+n9I0zz518Y0XpHpxISuDe9GWdP3
mISi75OwIw69j6TYNxnEq97GtnSJr5dV2y3Nx46tdoUhKnPrsdxcKMQBnJcDEXSz
kZ0nah6+tup4ElfHILv9lP+2tUfkGNzTcgykACahlTZI/nOd4blpdnNU0XTgnjRA
H7/YBxFtWMpvQ5K7oJZR9DmVZQzKbyppktLsgfjVV0fvOyUYgH26zPcaXOyySFyJ
BAGHXZrrYSdK+1uHH5MchBVCOAMtQ7lr2XnA/s1KGzGzPTWoAqZ5RA55gGGg9bkM
f+kTw7c95/Qe7hJmHVEaZznbHvuTAA2lepdiZDYyKG/jKBM26VpHz19mausg6G0v
GgJk3/DNqs8LAzmhCg/xMBZJfqz8/+Posf/G+79Nnxa33c2WUSkPghMvb4PMJLzz
tFto2P5gCmYeB0o0/Gpfo+Iiip9AdN+lfh1jvY1Zp2g7W8INnEVkPyuVnh3t8VxU
PtPi1LBjjPAJ16xKcMP7ylkcSNJfMUpH5DIPQr1qA4SGmOW/iDD2O/90KrM9E3wS
uBTQpqQm+62hSZ1KENXvmvDHfrUL7mCWdmsOcyd8zRDbhQrB8buRPYLygBeha58x
jLrlbMI9j+m6kNsu1vLbBMo9AijD+wbI9EWDcnMwz+dqOXC6UDyLtITGocEngzbm
tlj/0smVnad+BZcHrP5xXEntJisdDuIgcQlmy7gPfmdhVUBLavxFMZoDm+NcPdSG
Mh7fzNWxrbUIn2k1QGShlFTZky9zMSBxQU0JPsWVkQEEYsSxFb7d5cVRdBzAvwHU
Zs44SOhrgpivU37+eU0EXfsc1pNEEWLf+4ZugcVSBIBB3lfUhm3CBY+F/ioZIj6K
kIBWyqIku73CIh67EBcnvP3Upbafyj32I8p3v/6Gmt1mAvx/BBe6XJIi2tEXtqgi
gv50m8UuoxNbgRsShSQZ6ol/rmaIbMoBjTRzUEVgiaSN2pbEi2z4WrDNBIKUj8gN
2b4L2ICGjs8r3PiFLZZfem41q5Tu+5609D6BvldGoKazw2zbMXrhEh3lwNjbOXHF
IoITm0s2KscsFt6aIYbCGTzdWOAOOgF4wwCPnFRFK5HmP/gK3bK4PbmkGvQNKlSS
v/FXrioW3XgQzm7ygwzREXAsEYaKK+Gs15Iv4wlVhH+CLrlgVmjQfbTMINQiskin
QaLYHt4+UnuP9aDLV3XS3Vvh1OXW2AKRVe/qfAl0HVF9cBbUj49dXN0VFZIW7GYD
8wKCC8te4NyXvgKkYs0agY9eXa90MYr40jPW1EaR1wZPVRS+F8b91DILbnV6k3tl
AG9x9aiNLLade44HMkpB0ItR9n22zN7sGFQtShyRTF+pKft48CQM1aMHclCj9vDB
mqDRmN+D76N8GiqzhHzJcIwXazkOe/vWIYT6+FtHpLz7CY/9w6Vu2xxLq9gnNArU
akoRvlldWRYeXFz2fD6VYhms8v+7KNGEENkQSd8DGGbRqBMNrin7NhKdicZYn9Du
pQBe6VzoE2dlk4jGoqb9afC6mZ2eVmCAruM3DRLvvoeYtg47KdRzsR7+ZHNkZDjo
+d14sT7DYL2Hwu5N6bUDD0Fja4Vo9/BjYyXAO2ge/qafJGJQwGVv6gkaRkrVfaLo
LJGGa0rqk8x7EQeCNDgWLr27wNi6FjwsONJ6YjDTYTImP5ygZ08rf6f7Fkoerk79
By9eLhw4ZM3sS3gtsUdIQHmqhV2JA1/YkvT7ec/1KDNqueE85b649vEDMZXaKpoF
b+hE6wMPeZdYPZJGqaMYyUYLLjAXE4RwVj1TwJUBtbSeb4ckIwFdn81Bt/rN49rO
Vc0GkCfqHvwuTd+UQRogDIsLdnZ36Ve1UYpdsfME/gKYQarFCIA5CAnJDH706rOA
76sERDVILSbpjDsN4tBZr28jleTSdjpoiJT+SVJC+WA5r7pqKDIa2pBXxiHEWNZa
m6eyNJzVb6Dx7CDVjGZMychFCmWBfYt0InuXjnWB9JWR9TMNjbSZMoBW3ctqijTQ
tsN4t3tq1jH78dFqmDo9TqSZTFGZ2slU0Ly1HHSGJMIbiVgNoUnFWY021iWee6Hg
yne3F5sHu17KHp52EpgHo4S/qUHssqr2OGhddmgHLh+zmPPg+eCLbT30RN/xRH8R
z5tV4fv/6OtmSuo0K7XClngFVwMLgLmOKaTtVHgzJQggOe3Hvvte0yDTaA3c7l4+
AIpGn5CGj6LbJNl6LR7nEwWMYWePweOmsuEugFvop2WadFzmgobihuET+u5IMOQ9
KAQvrsgTh4qlaSBTPGDV5FWvRAOrrWZpzHZM3AIn+kqDUQs6rGJLuL70kh5Q41B9
l05FJevwq1SMa7/GMLtYO0OJSOsSrgZEkbiyPHrLQCvzDoe6c95wVmoYwRxJ58XC
Viz6o2ySC7D2jRT0JJoVGbH5UIE6UN9RV34Xz/4UhfrDY3tSeKOIfn0I808MrWb2
ZLiZV+WuDlZ0FR5+2NMA56ouAuCE6Qh2Ujw5e9PiPQJQKofcEqfs8ueE3S2JlWpd
vHh40Zhj9zzNHmQN3t10fWgddqQaYCtqmslsH4f0BrFDoqB0Fcg75P07cYbQr/5f
N2ENBIEoeuPz6yUTJch+n1JlblaMkf8VI8YIehuHTJjOoiUjQiQFeryMCD7iAZqi
pll1LwrsG3/OtNdLl23QvqoIbXYoIJQHCrSOjahInyn/j8vukLclcNK80J9n51mD
g0UTbgOCMD8Ye2lDpEAUvVtmD4GVGtinygHrYciAtMTSKT+AEMsVCVoeU9xb70Kw
evrcYrJxXrXG8D/N1SIzeQpJ02uN15498vUWow/oJ67UagW8iPMydVqv9Jbs8VgY
WFw96YIxdhP/E1nNoDy2IOoRzUHxzMhu/XrQ8CT3/dys2nllUT8FODuKfsO7qpMr
79shhfBfCR9O0JRvxJGrGtdWkMOwAW4qmxLjprhxxRUNBOkC9yMgiQaZX83IFklK
bPWCIE3d49/scDMymXi2PxU+ruYg9FQYyMqThzgymbL5NLP5by6VcdLPvNnPxzWj
xRI1N/HiwKTljW2tNiUkTUKEgkpovR9Tg6kdNZZ0Gjid9UTv2o+89Cxn1l2ds1lA
lLGOowM0U8nkbRIGpqmnBBZkRTj+HCjTmMsrg1GOUBShMG0oTjBdOuOZlUXj9zLr
ZspN2NR6rpraQ+9ZdKz3X0LA+3q2xEaSU9WXnowv3kiJz12qHotoiQwqXWhl2YAG
itI+LaBJKA+3suHI3F3fKGJyDssJnjHa1lLgQplazJxReABc+/eQlY+SUUAipafk
ltsAK6h9lwELIFEGADHzz8IKY0uV9zjQBGnfpmD9UHky+frk18qt0Dusq1ZMnJ0z
DI8To/9EWl8/FOubVQ4lnPdW3hdNlKBZ5+FqGFA8Z1XGQi+eBskcZx0VeUjLlpDN
VbDcFxfQ90U36IYUdGFzdbW/NyUkAIngaykPsaxAqQAtdcK5FdTytU7zSQyhUtvd
ZcpMzaiQLm4TXmox6eyXCM/90B0MPCkjbEPeuzXtmRNyMOUoFYm+kFjU7OKzWfcV
YKnKSsilE6WRZrnswktiYTSdZG1c6h+Pc1v+1I6o3qTjTw8yVqWiaMokP78URMcW
x/az35hD6qvLx2r99HKFoufrOC6Ox57cwOgLf4K/RiKlUbwUJrZ1GzgOiLDdYhBi
sR4/24lXRe3LYvppgyzZfXrfQSakN0d8QhwZq73HX8z0SKUge799ql1VQ/phgg0M
mwEsfiBNdL3mbXXhLixy46QVLQHEL0mlDrcy+0RzvoqMdJexiEmAE6D2KNhBgq6+
xizX2oG1P5SDJHJRWOUYEVsapbBpxQyIdmFQxRuYgqdNan4NN52eadDIy8GthfpN
tny7b1CxUnxevVCr3ZAm1epFs37Gz3UK8Of/9YEs7pWpb2Q79mUzs7hgQv0X7yR8
OiIhJ8A9apP1El/gK9nQYURTpgvLUad2z2CBpfewtfNAl9H2WMNi3gzTQx8DLpD3
wM7SXEj2q1DkPQSewRgXzmJGHjzpULp02VqrzsqwpHPMlLVbmeR0LjgxBMgrM73Z
vKOV7/8FQCCBC3V9ndlRCR0Qd4StGCEHFRHmmJS7vKhFD7X/VQPZCi7DMAdJCaG3
Fw6PLpucgkdp4G/ETmIj8aqcX2eeuUglymVHbLy/zNrETs5FXUZ15oYOhT7l+hDV
QjtsDb5D1x7CxC2ajug0pfGpGF33McNy3DbHXg2NHNfgD3Lx0WqFgvurnt6n0AzS
+T1uHTO7BCTsC6LF7geCMD9GTaMqedCb/eMH1CNxVourTSjB9t18YZpFUTrngEkC
Uf8lE4SEhS1lgZ8JisXX7s3/+XrIiva0d1uu544LpZKBPICKXougD9CvahEz+jYV
ZGGVx+QUtwrD/hyJO1r4nQ98WQ2Eh82yeeTbmZToz2HqiLjyadYEL3rfSRjdRiyM
9iBzIvVVw7K+gShj0G7uY2y8riHWgFoZk29SHSK+wGOYCFzMD8bYwASFm5Y4gVnh
S7GPRcMhrGfuGYoqICdJSeTgiStqQMncGAQ1x5tdRXvaCkhxzIGH18i6YfbV/kpj
RdWLug/h94j9INNQDleo3+T4mqomNo4TIy3Bxjl0ERYw/lfAYzPzBrcNenN7Z0Lt
zJ6IF3AmPW3JBO9KH+DmUrb1CHBMqxX1sf8pns7LyHwjVFCMsj9HKzB+8o1yd8Da
QAvz713sTLQDWF5SBZcU6rUC0hqBds2YCMVi0e2p/YgMex5Azz7vygBrGq8XqJ8L
OV0HlYufFjKNCY8Te2aMyMvTTAljzIgeQgY/PbDlLNo/EFEHr0PH5oJ6OqP7tI9m
UQvVBiwJxj22leptY/pRiZBQkoTkLpZX024Z6VA4miwXSQ45C6vigZ80EY/ea4wN
pG6cx/kC9ufj3CfI0L9QbvO2nHUQsxBIXzDFOfS/j1Uhi+leKRN4FbFAFq5OSF1y
y5hPQwnFJy/eXGDjV5DYfATdN3Gm+A1QmJ2LrP5dYHIQTYki8i7Cve/6FZoAiIJD
bKh/D3VYqgnbCUBDhi4gjtG08pzxfodv2CL8F0nk88LmuDV7+gNVy10Z3Tz6as70
M7Wm5it1CpwVqVPBHjMqwJLrOME62DQz2SDDb/yVmjPeNUbs6THR/QQd6btemDLP
HoqnMSv6tVVHc8/KYlpCnrFLOvQNH97SN7fXL7hR8s/w6DsOLnilax1RMzsuDc1c
hen6343aKsYH0gaRyAoGwQgVopf37e2C5kZ2fPpzb2mk1NCR32cKc2xEZl4YHZcg
PYdd6tShjdJamav4zt7ivUpADRfPViflcyzUtpXkgO6gSA3zyW8Upk8nWCoV3VeC
aoJzDXioDLG5eDbqsoo0M+0HYnmNDR+rvARY+HGVS1HxQJSPxhpFMn8k8rIm41o6
MelVFVl3uANj/TZZOYuShbbT1p4Q53RLt14H38Yo9fAQ+Mv7ssKYD8gPfVaGsxD3
n+y/Czem27GFOuH74DRZOqiWC//xIZats+2RIEO8kPfARSqwORYeO2I9OccBY4jW
OWGcQaqv5JRnc18M0jtxHTwAImKquC0gep/TxC6vapLTPxIGGXyKGnwExLEC4Ge0
64Y6uekIj4NEtGP+RlkhrzhDMfMX9ngiBNkA8I8GTAcwm223z1GqOGBAPwP9aVL2
GLQjCWStx3f+XyH4qzad6ARv0PjkDCBzYPc7ids5wH1ETbC95xkQ9Km9uwZTwyJX
5AsreCtPrlkA1j7+Z87SGhV4ur8/JeaH0Lgh1RBTziPLESwFnle4uZSCCDTwRYcv
VSECw7VT/UnS1AY7bNYVswRjjikAgKRIN3Kb4sCogaJpO2vVjINzraWkwgYfOYVb
Fp5OonVTOnZOv1lXlhbMJ/kHJDKDniKSYYotCVzWDfSLlH+Z7XswSnxwiGTKFnnC
npYEJ0oV4MxcfioeaUFGKyHuFYAShei6p+LcpGhvu1fBnZcLY7EAKcHE4ylxy8L+
+TTNT6xSi2FrRBq6EdH07PADv9Xj8nVtRYoPDJ8uQm6F00L67BDnOo0r7V3oGsAk
01FS9xj/1U7BC5C0WOmX5tQGlzVFLztn+94POvL+A9dE/aZt3XEaTiBOqb+KZfB4
qHGKrBVDvff51nCUEgCPtSu4VnQHBQ0kUTUSJPfuQW7CLtRME19d5IyjdmO3zyTK
Bz4rYNeHwoI1wWPlcqU67X0e+k4GGIrzNFOAKrpqUxKWqxCyGzCBXeRdIIg5452+
5pVJWnShcyE1O6wPjnZSnQRjhfLknJkl552TOYrYvZ0kBbsw7IXH7/pxwqBhpDVZ
uBaLZtPpMX1u5uyh8jjDzXm1hMJY9tiEE75f0V04A16vTZnFYkoF9bO744A0jZM0
xLhFOx/JMx2MCWY1hEBQ9GHzVsXa+0rsrPSHFHI7Y5KrH9qEXBofAaZ1ttlOFNmU
OhZAF9eptNAHiC6IYZwHEE2HKRMdOu8F2isUfkQOrZ8ZdD+TzemvMicvUTHouwru
dtY7pKqRsGorFU2H83rZNJVc6+kHeuWaV+aVeeqTyDYAHMnNNpGdfbocQ3UZeBeH
7xS0/P0nO5b6n8iON1wptkKgsh+YrGzDXlAM6/csZ03Geub/XCzsQ9ofXUz3oVn+
4pRgM0NudM4MY/+SlY2sKZeZr5+ycZu9SDh8Xv41RH5z2Aoam1XZYvFJxiOc43p1
z3M1/gMmMGFA8QTzU5ianT1PBOMrFLPlPfMfMU3X6H0Klk0aH5tfHhUF092i0u0w
l8iwISVWoz2MSt+TGIzfkQLLbuO5ExV+RwruWkD3YJlOyur4XaLobshLyJLgcmd9
s3RogmG/iQ/I0mOvVQ7yHXhBZYbwKpGmXj2CaYE8tQ1bfygXVUzhL+Fwj2V90y+m
KZ+rEKBBhTxhZltf/lO984xrgI3sVWcu1jsUFlIVa29YAIIr3yvbsy3PF86g3kaJ
Pfitxhm58EYLGdjvdfTtY8Jnt5rDzty8U0Rzp4FF4/dIMWqLbJkwdmQ3gkW+M7yL
UoYlilg0GIGVZGuDhXdqhleulYrjZl4vFcnVhys6UjB4k2U3XRZ88Efnae6sGVeC
oyC9AbD+fmwqRtqf6gkeo3ut4xmRyksAm426to39ewsFDIcPW24FW4+kKPr6puHL
55EoPxzicM0PCumbzdPwnGt0Ob+Xw9PcKgAXG7+rlJqa/3Qvd4m9Lq8IO1cvkxOZ
q2xathXeXPeT/cisNhgG8yyxM2qd8fob6hGu4SyGNhLv4tJO3XNKDbtFnVg3120W
Cb3j+mIvIe8N8bZ9meebBvJLKBNsUPK/KUPgvw2xVY9FSuZkTnkwQqum5WmH3Ts3
M4G4ys8K4F1X56/E/XiAkHOAJ6XchmMOVNyzx+mYaUbh+avjkfzokYCvC4iso7Pg
N0V43ZMqEHeUL1VFkoJq+hslYQnHRyz7w8rPwHHwZxxIvAyTVdSWmLBZglofv9m+
a4ZydP+ts8B7LnehCkNCTFHv3LrfKOMHybcpW6DsPXxKXE3sihpq8auX6KR0PS1Y
Kvaj5wycJ3891kaSyaTpV/piDhHxmDNz4rvdTIumUxIedk7zsfhw0aqMlpcy8WpU
XDfkl5ZdGn4bgQ1XExdmTjMs2DfNsUGucZz4vKeg4hvc2Om2OLKARMvwRPm6PuzD
o+2YKRoUhIhq1vzowJ/l2jHFtHiyWCFXQweiIjodpimAPUgd322wwSvODVimgM/m
L7MvIbZiu8sPRF+ehx2OuOPYHGI/hqHCEMLN7QMJhx4XUavj7MboAQkXRWrgQvdt
GYitq8V29X3DjWHqy1lCcqDY3jXuC3YE8gzZs4o8L9jgUiPzolTWeh4V+OtBIHDe
HU99c36hCezGz6jveM34C6eUmB98u6i/TPRzqAWjNECvVu+XXNNK7I/JCCfWciOA
KLpb3X53hBjLO85C9j9jTdGGDq/zEQDrwShCT10jNbQDjI72rR+crzBRwpyy65HR
1oSpwYjSTKJ8kmY864SjMUAMjeOrtKJkzmoM2lRdMzS+ImM3SyzJc87F5gDZUHGl
GPvh4Ixecf/Txui77hrgg2nagXGIQPxviyB4CmEUuXXx+zNuu1FBOxFKD5YJWxAz
tvB8AC0p2Ezz88cRMA5sAMa/Hm7NPwROHfrgUlNQiIVWm/z+FPUmcdb0++d8l+lM
5BZiLfgsRP9roeXW5JqKEndAbEEFM+IeP0BlgbGa8uS9jYH7ZQDHy8gJE63GQWcH
6U12d0tJ39IHJH4TaNfj8Y/wu1xh21TRhFTkxtMJbj8mQtAK2cxXE64zVu7Lyq9f
aXfy8/wMkcJJ0ADmpK3cKHISgstvOOy9EMAkz0q0EcY/lDvYXMcJ+4HtnsLGVTzv
rSrThLUXbKsPrbyNKj4HowdILC647F6ooO7vtj7a1HgGtrdb7cGHa3vZItbuqHv7
y5HIsZlbnX3j2XI/u1LMCtyrYIuKq0DurbdDPHm6fpgOodCIcxFjdgd3lNJg74vi
uf0SIvebwffJO3QsInap1+FFVtAFLMYOOSIYm2tdj046uYzdV4jZpqqfbiSKP4OO
ieXlE4XC4Jwb3b47PNmlRAV6lmHX8w6okKOdyR6bQdrI4I6aVjaTiILzY4jLdkeP
Apvm+yToY5Vd/rKt7mbbeLJwqQt7OfcEqORsRMNxrvm1JQ4qt1hnyFmph55q57oM
0JG29SXbJyFXdnOfJVehWMQej+qOExNyDJoZx6YS2juzIYC5faAkPX81tMZGFESF
G3VSCtxn5nVlLmhbmgMGVvtFDwgzpjBEb/vlA/9vEaujaVFc8DY6zEkoj5luagSg
SLTz80vg827yNTjOmxgYsAxq8Jglb7v0A2xT3R66iSYi0hIZg1d6Asg1VoEgLuCD
fZSFSAKRPEBeu+rjRSwCypMRXctqKXD6VQe2+3VcoGJEm9zmV3erUMrLynSq8FcQ
9zWBnbrItmcxSyNnDTgxPCMe7J2D0gL6Jx71NKGr4rZve3VHwunIb/BL3oaU2QR+
lJJ8Iv9HpBM46JIzToIrhuQNftRiuDruFZW5KiJYa6QqyX25uW/7dBcbjBPBHb7X
uT3W1QUlIsC/ocVHgfIo+ZnFGy90H278dMG06VM/kIScon0W0gaLofAM1Lio8Zdn
agJe6mYfTf4zW1BAHaKuw49B4SXRuRcV8Mw6Yqer4pHOyiMrhmpTmjT68l7gDNJT
h/07HrD9w9Wlc7xZ86UcWZom4AnfuBt5zuSkFjNUJg9yQYustIUHOy4f39GtImzl
JKUI8/Ykcmh4CZat6PsakU/oz+sIuDUk+VFWjfCUPHUzVD0q67XEEWnRO+tAGTM0
wtrEXHD3TPMK9fv7W5OA1v5bCMl0zrN6tHsvtSDifalPo4yLi9/L3HELtNDf4tbm
HTxSJFpZxiN6jdKG8cPJ1A1g1RMjjiISNz1jQ3DkgF/ETSyq/mRiW3Vmksg3H94t
6d/L58i7JsH3R6EF7rqaVvxFI8PSMwxUiv62LXiKbEhSVQqTw+NIsn1p/VMixvCz
BxemgyWL7I4ifSdmDiRf+DqVlXvuD/Z9dA/r9D62JieR6ZbqvIXupjctQAqgZ8Oy
/2l+cQACXdv0ZOFAy5ZWt6xzL88pqhbMgJ8XN6W2jlsoREIYCY+8UyWx47GxWdHb
MQuOj0pG25WpW7U7xnV4wZNcUzCWJdYw+Y6tIooRH5RvCdTLzP6lOMr6iihbigN8
M21/GMWonRUmsoAJhZg1bLPF/tW7cBezVGrpaV/Al+vzgkwZxQvaR5arzzcBZHJs
D6OzRJq4NyjoZWMuT7e1DHgtLpMo1RqLs30syCgYLw50TN6SiW0+NABYvIRhQwbE
arYMey8PCJnC6n0bkEPfsZ/1IgMn0BTOknysOP4YqOPoSZzKdEyqzaS49D7xVcJE
t4iGOnqMlTKY2Ghu4EUqyfSMEpb3fI/5DT5kbzMCjesVG8Yrd8LLFcyAmljSK+KJ
+Sz1eEgXiT1FGabD8ejMuuuYxTDTajOC4A1pLFMsnguquN8zYzqIMsYsABsJxlhF
asnAJBgWMKmuIkwLFMeH0mHme1B41IxEt1i+0RkMSNyLzq1FpDE/5PmJarsrlXCw
ol4ECqVLUD/i0KyqLuQsDHYFYN4+Cf5R6D6ZgLAD+nrd5ifF+3XZ4kFKwu10BOra
u9TIBpMFVJNnU2z0C2Gnd+vIT+GBLSyy5hucinx5oazx2vEiOxkIU4VpGVTCy6be
9Yr5MnhusaoW2Dwu9jOJ4MCsZ4t5Eh1iDPqtLTDSKQb2hfBRVo1dlHlIGl1hz20K
1v4OeiANcagq5hsYyOGKSt+A8kQ/rSxwywtLos9flLkn1TxAAwGk318pDQKNU2aN
rV6F267aEqn+gGN2MPg49g6l7bzOq3S+n6I114fGrEfSs9GmuPJp2IfwGFeD9E03
kWQlM6MdZ5uy3POUbI5J4TRC+oNVngFSZaTdJlG18mbAkJPde4IL6rbYuUMwLldq
kwtmijEwcVTz5TAHhDT+nKibcpDq8GpuiaY8N0q6Jv9PfZYjYbHa1+obFxbYUNjQ
hoQyMHJ+AY4Wim0exxjnR2E76HCI4b12k84Ludi0UU5Glvi1/kPFBkRXFg/Pw1EC
E4yTxYWzGoS3h9etZEb3RVyDPPH7W8DCct00Fg0SlFPsNGSOCFjd9KdlTnhIrIVe
h1pdaybQs82SpGrVtG/zTwLHcnUhHjAddKD6IY2SLLk41gAaGM1CzvP33Hx92IEF
1h3SKA2F5PHwpXYjpuWilmt8JAR0q1JdmzQSdI/HDswbxbKkc9LxE5xb/2HFuOAv
S/Cot2nMOlBVss4mXxDiKvtxsPXxH+ENEBRAmtciL0GQ2UsNpVS1gYtPQ101weHz
Kok8j4YJenSENzBTi8RntPcwUJcAab7LXMfG01ZiFsXaBgSQFkiew+mnRO9Ko8XM
K5N4ByglUjY3f/SmoamnwM1DqhmJj+wqv2F9SiR8yprqXravxiCuUp1JjQQIq6NJ
dXwzWjjY9jg6zUpAKI9JP1FP9nDuC4GUIZ0ECYQiNvQgU6xE6X4Lzub5KcM2hOX/
8na+SplVn2G0RSUrDR5xQRsWadxdGfRZgE3EuP5ZUdlmwBFM/NT5xg7vHTqM1c7H
cslKak9z9JmfcJkovoA9MEm98x1VaYmf1D/7tpu5GPc4vKmX2DZhso0lJR4RH3WC
n8IZiptrc8/GfeltdtdZa2dXuJGo4ADoQbyNLzzmUqrgaDmBQ11kXGrIlXfDUBzN
aLrDQi2HXacspwwehW2yxNqRlx0cwMxtlQ3GQHdAr9dTlsjIXXjrbo+wx4PE4leX
KI0X7e2KueF+sWPIPiqP8BkLO2MD5sG4cz6sZ+2RnCW8tMvcz1KMIHTuLkOMnAdC
k1oqAz87G1DkBvmkSijwdsljks212bIt/LEVT2E44OPGcJlUIbB0PsE8yt4UelPt
Xin7tZ1/T1msGdI+bfHzuPJDGfwoPTsVWCvQHvYA/8xHByOZ2qpMJRgcyIMmMZpB
yAnCq/F60OJ8ftMVN3sIzK+5VDwTQkIaC6x9apltNYI+PgklWTXFPqyTxrzt0/Ot
YYhxejETWy59y+fPeBa8QMMev2ynHDXyZm0XJs1d6j5f0oUGIgChuffR8PqNuKtC
o2QbmyXy4bfdN6rAO8FnGpVULpzaDcezZrnScMO3fJH4SNAZg5mSX/WnOHIhLeZU
bo+c5i5Nqy4mqs/rlBCju068aLhKDnSjAciOmMWRwnnSSq0OPXBhsOmOa1mOdQOF
0LtOSQSrpREbIsRLtiIbTAiEYpYOxVWjIwC4gXkAZqIJcTJfnVfJ37tSmAA9PvVt
DlRijxmJEyfy6CKA1pQr9FP1ifj3pGREMcOxU4ZPq3jXeLv0AwVFXo++3WIbmQVw
M/Bg+oJh8FyjdWmMVfFzMiitbj3GXz8+JcOozyk9V4tOiPwl+toqzomBrjGyl2um
/n1/AX8qOvZ4gVkW+p198JDy76pYJY/6Nu4+jMQgU7MyNr7QVsVKA+fxm7WHy6dQ
WZzaTcYLMiD0EzsvadY2zvBubCRa2nRRiNc9+FKN1bxCwh28C5Mqxq+NQYtO/7dD
A1tKFSaMQzyw3pSrSxWoDmwndkI4AItOfL/JQqIK5oDg74Sz+gTPCrvOK6D6fj7K
YVH6B891+lRQZyTqXt7IL/sUXP+nD+AdBo/zaC5NMixxxzdEoqnyVOrSylp2X5tk
rZl/4y+QwyHJLq9L0DXJ/5EO5Twgc2PySDypAPDRuGTpDHzYNNIprFKgLGX8dG71
xGdAF2SfWyPOI70kbVABfBd3fqDtB8nnpsZ32sPWdZmY6VJF2iI3MfvBNOUEC9It
B/QSQ2r04H6GCpp2an8BPG59nzeZwQ7IKIdVlmlhyEemFjrgHAWEHde4XtTnZloz
WU8/TWfMp+ChjPHT+31KNMxKltBoPPW9AFgRezCrTm+1vahMIy/KxcTrs3qU73yt
KVdz9UhhkMNcjuG7JblL+XDmGVDSnxzTgC5Igfmh8yPl0SWeMd4Y37QYjew+VdSS
6UnCe79hI7STVknj88zQL+KsmJmLdJSEFWFLBDS+pUixpmhosj5utj6zFR/yEBaX
xjdjEVqflxRwVzzftfLCXh7ZrlJp3wxkbE+V9ndQH9oee4tFPHcU1wf2UpbKLltU
cPkkEnUiaS/dy9rnqPGuopngLedQBuYxVWY7YVyWLI5aexbhIwTz/RxBTTcOEGx9
yaHXkoi857UftjnfDIo3p3AjT54aZPgAfe9zCMplR9dALsGIvxwx0TfPeT9DOUAC
2oVtbB43f9898ljbRdFAPq9C9+0tUnEmNIU/9hPEQdO2u0mhqMG465RaLpPb8dwF
scuz0M7cAy18TleYPmzUGZWDzxhwZUxdYq1t0d73haA8hdW6lVBUNfqH78xDTg5P
XEHYeuQBC5DdjR61WWDplr3cWZkYm8eCLTzofnjtPB7gZoUD0gAr6ci1WdMDUNXx
bLQqGtwd+Q7buhQLsxRz5Y5It9gPKYNycnuXDOKDOyVYFQX9Cy6QgTo4PZIIXY8m
YCYtu5cXBQUakcBEf9HUeBt8GZQZN/0jWK6Qo2E2zolHrdusOVhobx5qmyJCl3iG
g7eaE/2h5u8Qz7CQn1ipG2UEh8irR/HHl6f1na6sfuDjO45xiCH5ftwdSn/xXatn
FFPCafz/hD+134o0pAt3RM5VFh2LvAlBeMic1wFpDVgaPC9bgAMp8dz2JCUK0o1h
BSYped9S1My37JR8EOneb5u4p9L3bR2cu0oI3kyx+Vcb0xdfxpS4VCWnDrB9FY2c
dWnonOIu56ThRV8xBxX8n6MQDwPSnPm4x2FvetUl7Va5aVB7Cq+/995Jp+ZWOHAt
wgjVHZeNwt4SS+zR35wPiJc/FtYnr7LJXQxDTnd9PP8q0LvwG2KgqASJf6vQDPnU
JGryJwLWoD7JxAgIX/hROYghbgHbArQ0badj4bzjefPCFJL9cLs0LxkMLoYWjbjj
SDph3xtJG7epD8B6OciTyVmRyaUJuNCiigjR26vptaT3ljURNmrFnznX78gfNQ0n
M94wZIv0vjTeEKUYBIH8o60uO8QojDn27WqfwtG7gD6IFunD4ChMSWZFH+iD8sN3
wCLRNvazv/rKOpZ7kf/oXloOZXNZkseRhPuomn8Jhz+B0nMg4Axd95I1tTp9GEQq
JnsswaLBlhoBUuUc9LOs8gsNJh/1bRspwNN+4VRa2Ol8aXbAm1EQGMGErvE3Vltd
56uRkLblpeHqh3DIAwR7m7qQhIiQTBKitZzk+MYk3ucuYr3pR0K3NyDaddLdbOHu
qHvLnVpjI8Lm4mFD1y/RShcadXtu82msSNpZC3PQymQ5Ig/xYdWVyiU/7PZSDWuJ
e1k66UCp9pD3z4CqFL86qSucSAED309EFLk+aQw+EIR3W3c57ED0+hjOsDwtISg8
n9ZPJlHgOHNvsfyeg+z4zpZM5GwdwDhr8f8rt4KIVbYPQgb8JJw2UKCmyXvCmuX9
Btgz1hlR08C8W8D8nrFLFftYKtWEvY9hfntPSUCQbvugIVcLi7jv+NkADj4F0t/7
xoMEqoxitXD+bh83dWMfdONC8PyjttxvEWx9Hu/hgdfZUnp/pDE7eCzFD3xz2rF/
KV8bcR6FoSXOvJ/epe0ukbuNXfGXEdhyNEA6Ob0Bsznc90XnJcXpWMD3yJ0OkZ6D
L3J99zL3jIIgM0FB7RgLEN7EWdt+1J5pybMkDhL3C3TOXmoXVipXY9IegifsD1mV
i6L09Y8+Wv2xQCdip8DVlb//G97CUOgS1fHpT26tpS7NHzmqJgsiYUepNHTcYZgk
e3QVtf6kK8IUmKZCSz25A8iM1rmg332fbIN5AkmRmc4Sbtz2Hqy4tHZeuXMx/Gsa
yqxiFl1VsMDP6ljcZLFn3fVwIpfikRxqVuLeA0qHoqiqn7tojbEz6gbDpEivtmqN
IaAwK8VzNkTvWxSBMBE9WhXMzID3GUBHpQ+o7ibSWovgzI2ODqgGHR14ZDe+0MfC
Te8axPtn/vODE2FJpi5Q5Tca4kNqzwEZdfO6JWVshUahN+ETbEEhZEIorbvCkK/X
4+Pkk+8xdvyCZONIHix1r9n4lxRFpeWmik5ZhIQLMXc0FMEMAacbYJhP9m2FurVB
QDgki8oASpPkINXb/f+DdPzkR5GPvnqaDZ3pAhrk56ovabMNi2h0dlDeaB+3bW7d
IAHZis7CFAdihhT173DbcvP/YF7iwCQ7s1eQQE0kKl/RWHJAgTdO7G1t1wFyNjNd
jv6o1Rd7nvEr3GgDbcRjasVv6alEdS5yTpmiy5fVU5bR5ScIHRGVB+GGZTRqnKXW
thiChsbePqD8wtxn6etuql5iUKs52N56YU7qtkBzCj8QUQ4cA6DCkOmfKUfz7mKW
TYkP/Pl3ow0FlS0q5HghJUCnf9P404EKvQyerFYMVbBCW0yQCwKMEHQkjjWgeXsT
GmL3y5WyM2RYcorG2KJwReQ0VYBJOUy2N8ZKHqbWiZwNPfG1pc5Dejs16H8sSAIc
0XnjlRh4Pnjlda8HE6hqvLngUbfCVPecHLCuKmzBArlOFq6H6mLXgrxzHbTNoRME
BteL4cilz9BAzkiyW1rJkYPQoBJYVZOcC51TxqLclRodEyZfjdvO3h8cSQVf9G/J
S0+R+OKZsYhscaiuMgKlq6oDvj43AyUbUWEZbXfqLbIUjmAXaiLd2JgUZHCYPD1V
hW2snagun2aa6w8U5zmD4R5Z12L7gj4Np4DYO1o9+k4J+x2fwpi44L1ZK5YyHaeg
Rwh5aGoJGJcgO1JoP5dgbBbyVlXY30E18KqUvjpY/scplK/XMmnM4T0eN1QiTa1o
yCgf7acTe8TY3/NqxKsfUIouDZhxiDojDutlC1xwvHZAyGcIakJdmC/M/zAEY4gk
g1BzWepSDsqtVoILlZBWH75o6IyQNn/FDnMK7URS47EiPXwSLTOzDgmTAvHRDEUE
zmLCj1kCOa4p8ouBiVqFwrLCMLMfgzCWy9U5wocErRLxTdxWM5+xxgLtiTbPApjn
SDtHJz4FSRL5cPWZq5EvEyQdKM70WoHzT7aC6q0JxKaL7kmt2VEBw4EAq8aZMp/S
iQ08ktk3q5mgktaW2klU5MVXTMUbLPwwbLnYbHZUt8i4OqG0o2Tqm3YywAUi+cSX
qLuPdD9sBApBLX8108vH1HSb6ovpqhuYPKSwsWzvrIzYrPfb27s2haH1WDXLcs1x
/Ev/twzn0rvOiys0FL/QJ83U+4qZe3HwkTkH7zF3X3ExoGCgIdY0rZQo4stsRzli
xTryF/hfAuFteI3aYwriu4CAqmC5lvvDi0m5X2WRiPVkfrbl47ASQKh/x/ukTB2X
MQO5d4bbh0k7suu1U/hyvhbqrkDlGFgf8wWMsEkwoTGQ/54CuYR1yPyJQmEmPcFX
3k06nazMmimPUKpAdZfGR89JXbsgqTHmtDqZ0mQIKm16BT/Imv9L9uFq8DWcEViM
hyaj+8TEL9laKbbyNMXKh5ionJKZ0279+TWfxmDmr7EmUsej8gqgGRa7VAYicw0n
FE19Jo+kvommgfla4Oe3lgHIL8rqfPm4JOy+9TP8oVFLMIhl4AccnietVsHjNg+3
CKqSI2I2bvnGqLNS5kTuIbx+Za4V6t/clEQ8aLMnjV+34ENNhVarQ+nk3h71uQDa
vGQV3PbgZIyzfnFkiu8a7Bf19y2siChsgehL6P1awLbDMnHKtX2WbQfi/w2PLlvn
eACc6tfDRfo1sgt3c3GmIX5puf3adz/m1FIh/M9em7utrEygvhJCVcxoa0HBovY3
o9v7xIqKCc/aablVklenxq/Md4AeWo7AnzDWA7+4qN2iVeLD28jzPGtEiT3hJQpX
w+DPzYT+2ls2AZLV4kcZLT+Od5EwuVVZbWv3RcNgazl9faaBV+bsNVAjk0xjMDyY
tZoS3oVK/jHk9sXRUqKV9TiUUP4u7VWNogYcaNla3KSf4lGwgw7hcHDgFp0iwHjy
MBmzJH5PiuhSUjR4M5Ej4FHaTfcrcuGiL8JXRceMjDBH2eHaBMNHfiqjoJOHeftd
ve/fwYeJD9gs5dqS4IAq4YdS36Al/k9P/lKZbid/aBO2nBgg0s58wDsx859IBA8b
2yyuj7moVyiMgJjv6hoAehZhxsS82R0wkPwvTbOrbK21IT5nz3S2Bq0SmIgCzFit
8p1WFa0IokXMbydhOvr2OfN+W5q8lA/k2/9Yn6/y+Es944L7ObanTyVrtygvW2Sy
iMjRdyi/NHur8ahfILlxj6HEznACkyPGfH2KYAoxdF3+wb6FFSecLlyy4d5QsAyx
O8EWODKsbGbcpp+8AkmhW96PaYaMY9VurKYydsBQngR1aIYD65KuQRZPKMJfh3tV
o4pNb29Al2bavcy0ps6hm2+J6BfpPVbak6K5A77zmSQEeqJZtz9JbslZiXMVhKVU
5LrbCkFSR6OhaOMkGGi5ti/bH2hpTHvBZr0Dt+CJbGUip/qe/X+B7dLLvChyQiPo
8MFwrzqqLdsICww70UsGWP4zrtGlPejkW40hQlko0ZDlqG9VcYYQgK7eHS9GREVW
3mLkEq5PT6Rp32gvsJKeXqAduAJwi1LJcJM3hqctkvtgiJudgJOPd4maaGijtNN1
PI+sYJQYMYkr4MbKBTGJMibzWxs0XWOF/Wimj+7dur+fErkpZXdbCheYavCiRStd
kCNCQ38dg6knEVDOtMChivlzqTEGxzYZ4UOR8nyuY8bS+cdbq5+axbVNqfGhq2bD
BoyhVR2cOfIv3fiNYOMdjXUKIskiJXlMosE2je4HitJOM3Pyeyl5G0TY3tEtfdps
qoA2FNFEkvkaUeYpSxocCm8z4U6dkCAkgnrAbbojxpLFuwQPx0z/3lT1sHz4DAAE
qdi7QRHqYn5ra0vRy7kgA0eQGtBrwSPZa6eQGn3fck4rEbx4Lx5hlytVWEpb7sn4
kFvZCE+0PbXsx0BJXzO2sXmnjkkSlzLTrlWPo1aTwfBfoOGy8ueRNUIyan27ZB7n
rFDp4TX+ev8lr13irfE6UUXcBqLbOTf9ph0Y7WKNISq6b4utRZQWs/zltD9oOWWa
/+IOGvMD493c30yNzrqTIaYa6ndaF/PG9YgPb1u8kuezpYugHjPPfMx1+cj8YRLk
RzKNNEK1BWYnJW6FMxeRkvgtJxMWPuEmdRRY/UCZNwiqkThV/WEf+Icqpgtic6HY
XQJjy2X9pD1jZTAYXQWJU9r75p91+fQtAlXVXq9N0jZx4Ntk8pSzFMTIFchCJNL/
vU5WGC8K81ep3ictPi9Cfmj3UGw5hVaER+lb6AHDuq5uXQomtiDptHGI8lqpSfga
W+l3xg8FggI4yLnmm6B0qVgj4YeKCIQZzKc8cjYEgy0ifneZXmQcIgD/P3qU22aD
xbbGKt3dlu2+4rwbCFiNv5VB8NbkW8N4q6UZEzACF+1l3NLK9YT3zRZnakcP+tle
6LSdrVX5BM5S1Ytt9b66SCT/YLW+Ha6R4YR+P3yCnOMJzFmbBKq3mxIVsm/PaNFM
WXhx0nY7aWGG8383QcTF72pciLKA3gM2nvm3fZ7qKxdhP7cjSpxakZzeJRJPoPW7
Y/hjtKtEQvH03kQGFQzmgk+jj6T6drhGRTm4/RIEic511LLo1LUFybAhQ5BL60lA
J9MIrkw37exQKeGI0foC0BaIrEtI4cCRjVx3pt5Q/5Vk7jPiRyiNysvzlZFVD0lV
OfOMVJ3rlLfDSXQr23xbug99VV429raZS31LmMC/K/SMAmN0QpigZAHIp1DeRvnA
JuvnAu69LskzFxkY+CokArl6E78GmrlVXX4K80hwalsrqwSgZY47QaVdRT8lH1p8
SF9dqJd+le3HdZmMkIvKrZgn3JjQrkCFP+EGjqiTKjavCegxAWj21eOCxBcamr7l
I5mfCAfirW1ptlTYMUZDhpGhb0JDq3denweQFuLgxTnwewqc2Ls1DUzHM9n3MreQ
FoTgU2eLuTKpceVLNdj67BrFYnFj8L3jKQk3B3TcfNLEaFE5N0RCZpXZk5mC3zVb
e8sWyt2H5afX9bqCLW1y1osQgv0Naiw60qqkde+AHZHBm2Qf/4n26lSRUvvhOUL3
FY1vhlR8OABQqdyMbSVrRWPb43kWakiNHL3nB58bWDA7ibqOpOLBqL5fX9VX7ypq
PINOfYpFAWs/J/psmv8d2uCGqk7wKBdZP5nwwuNksEeeX4gD0Ap7Bd7/9kdTop1b
siDnzFSwLR0ht/J55lR+nJwf/QU/87YIeBGDhYDI73KixjRVTOTLUju9N6F6qMkK
NH5Kh1Fpe0h03PAN8HKVjgikuQbk+oA8itC6wQzMgFNxU1jl7JaTlOlx/p13xvBJ
Wck0WRzp4qsfuo5OjDTKtyC/TDGQw9bwo6w6D7T/1wW9aRC08+jv+7v+/lirBwNC
Is2Pac+4PEuWlDz05+/xVz0QWBXVTVlboD9esa51QdrKPoD6UhQ5OsU8671gkyOo
rJ0K/3EKEVPWRkb8zOEgqPFhzTXUqOnKV1h4Q7+zQOsU7Bwrrj34l7E44FxlzYPb
iDH2urGhvdjsLfHcfyvj4ATwdgGq7vmc5H+S46ZM9y+DRztbFG/GoIW0k8z2iUzB
id3gqscFtNcq4eJ9FcokwmuCSKRzzVhH6uqRDgFcjt4AXav1ZO0pbpbTfZi+G0Yv
hLU/1MQAla/uZ9xjNwHM5vvj6xWF5y/MpHfo4gyv1cPSXSef3Du/p5/Yk2x0diOG
WyQBfydWLTINOUyUYdlPyaK0SbG8FZGHMBhuUk+fDt1io7AIeRw9hLreACR4Da3N
JwfIz95iR33gICVt8aTIk6HEowPm7w1Kynng8mVXGTj5QLmHj+V07JCAaqMupH1D
7Jx2xxhVOnF2wXWnkQ5ou6qBB8rtv1xpj9zQvnhB1PnX4/WIitWf658FE/pb/tP2
1RB2jjZY+VHUy9n5uu6MB6LvCa8/aMIuVHFzdXTuEp/JT8/La78CPTv9CYCNo0Bd
miGTwOTTGTXbat3vqkoOMvtnzRJomc2bTBDLJ301auCUgwYPsOY6TfVW7SH1+fS+
OfJNc3mjpRjsJg8ZKBCaSlK1fp/MICFV8Jjh9k8RI87jg+sk/1EwPcJnEovUGHiI
+ySQqoFj7aRO7z8t9spLrQO3HkRB9p99SFtQ17FyyNffDtJ9TeiUzMWKOIqau+cm
5iJZQVDjl4qhwxl1V666Czsq1PAfJ0VlGL/FbQ4FaL+Y0XllCrZwdciOMKP4rTeD
w+MGIYejEWDXaTHu5lglHk8IgNynnd3v1pLJ//BoKO73uMuIu13QmhCubDMkxVho
7YfKp9xQLlx6a3Acv2qfCLSP/iwdudpONUT8mG6xaGFhEkozzV14Mtl1FX4Xg06/
EKN7CrJ2poEGPIDRIsxGIjDPlch4iBnLYh0TwIH4mLrYfqbkDxHr5SlQYcSbAxar
rDdV450sY3TkWzZom0x8dj+J2g/uJIv1VqaZxmVJJrvRCUc/WXnXeGpCWmvCE/69
Diw08JVaL3cdIn2OsZ2sSZJ/6VD55y5Gke+gZRg4gfh+buoxXEiDJ8dSTEdgoETl
NoITqqGxFdgwxpXF6tKV9tTvLM7dZXdPxGlc52kNeHBZu5uVi9jgmAK1rhukxrFL
GY6jXWjundxbEcNMK8M3LwiX/kmD95qVnRiN1ws3I5cUMYQEvBikntZ7Ml/CaVDI
5telyWPwmM0k8VPN4HDXGPT53njsRLbOPOjysTXFOYrKL3D7J/v2AM0+Axua0jpM
qD57zcHHtNyLGfWPZKfZVursWBLbnGsIm0vQymZ0RVW3tDyVh6zOY1wqKfOAZJ12
RGc5/SIrCsNwAnyF35n66kuFhkJ/RHxXnfyTeBxcq4sRntYBmiMjKEUk/gzq/zTm
Tb8l+qMM6rM3Ah68gRujRS9q0NQgNyt7xQjKC0Lx2WlDTHsriTYXMwTa6BsOD6XN
sKLj+ivIJsMP/7WKUS2ZEk/YGc3PW8+LlYUlbHyt8At7C1RDfTZigJTHiB3pbTdJ
0mwzwPr6xpZ+nh4fnLTzS6SjuxoG/PmcOvxYAhfuyY94boH2XUXWLE95l+CS3w0k
Dxf7jSWF5OUFjubNTWAPdzG5vJtYpY6jU0lslazmdZQmY/pbC5e1oltwZPjQDzqK
22Y4wwlkMkCDy9wK1FkfV1WCg1Cuyiw8+pT38jWVc/YO2YqsbZNsPqUZi/obUC0N
Aj4x2JUwrcWyvhFFO/fcONOYkEFRHjAttPv1Cl4yJWYOE1swmSYLj5gng/scZGje
sfS6jrcvca2B0ON/eK6RkJ5+r2Z8Ux5LiQvaROA8TcHDhiC9Bbdvabvei1ueQLUC
Qc6+qpywzGlCsAm0aMW6RbmM44VBcrpYNIpN14FBuxu8Wk8Rf8E9U0N8vLXzi8Zu
VR6380cDDEwik9cJAadJpz+8v5Xosebj1VWFp6QWI32B++6TkGPvMj2XhqGe/yDg
G1RR+DCiXcD9HYpgx73duy3Pkf9guJ7HtxAwRrKRhaGMtTJKLyCOYoyovUKe37fC
xfcEPLKNQOStF5iAGETb9o+NYW2qH6GhY4Go4ql7ZrqN6GY8tp7yVFib/fVEI6jg
C/A8q0FDK8ZtDX6RPBU4ysdY/hwaPV+ha/wtUdiFNdx71AL7jV4P8Zoq/tnugQ05
5BZS4BTmjj25Rzwo8Yo7SEqQLIHvwuXB+/6bF0rIw91aqi+hiNeYEknLYvW56Vrz
jzW2L9qxCOg6NsCxu7/aOmIxXKc8vjl0jVTrbg5WHbWfD3n/SH2FGlansQPENHtj
AErUPN1XwCwknb4kO2pU3rmYcWhcfFE3A1xJBnQ6SLrUR4d7ZOunysAnMoQpZNfR
6G32GteOKLtFZaPBrhjTVritww1YjyNyElqgl6FMoW+es2d+lPwVJSZ+iP/SbBgl
D0Z836AjxDU83iL8NtjCGRjGr8/D1XUJnljPxKvj9m8TNglq6BkXDfTbMe7133TJ
3G9qPIQtHy23x6DrMK9SZu6SS4NigT/P/udDuYsghZcvcrIMAMp0D1dTLmlztw8k
bGu0jPNln7bxeW7YjXe8SBNkFdsUOgqFzRFgR6mh+VvjVKBb9Ahh4jn/CrDdRx2X
MASuWE11wgXj1ppSHxOUr0fkcBal8u0mk6Vs84qX6TJOXYtFD+xlI0jRYBmih225
BxfmxPwFeBdhpmXg5eabuad7JA5EH2Ika9qWj91YzChqr1QTLFyeIlzkpbt1EQ6l
v1dj9f7luyketxS6arvl2qNcioWT9B85H2jpkS9up2Jhb05KSTq354LG6yqoWseT
4IYjvYacL57vPjFqxpoxOjdRTk+5anZzfIB+EtKtJNQl9BhaJG1r9qztnGWiyoNG
cmQIe19Zd4vy5CYGEssKabsj0haZlB7Ds9rNJl0mKg3j/fffCU74aGUdYECUjwIU
9Ug/h8C7RQ0z0ULKhu1jQm+eel1NdF9u7boMs036kWq2CMfJuKyPzLo7K8Ssx1yo
4biNfMLF2cruvvt8AEi7MZg8FHv4krlc788fsnFd8rlWakE43bqL0nQ3kxwIvdJG
n+ZWigqTkxZuv1i5F9YDGElukaCgjjYyF/Owqh0zbYp5+gIDOxxY/QYjF9ruvfG4
5/qAVlQl9eI91cuKs8mgkasLo0ZCnlCgtVaxK1BZX2YPrrWSSklDI6RdmknD8Gee
e1JtZNHkzLveLtqsG4pvAeeb3+ZuN2qf5ENMiZIkXiwIRRB2Jqaeyl1In2vdpSsV
Lg/amhcq93wwsZQwkKZL8Rc9QVBfjBhJ4EYYxrF1S1+0hhhitzwgkRlPm/gKLaW2
bh2YXaA9Llu1g0ahUCelTXbmD5cIoRA1GgC6U4eO2L6rosL969yLCPJg8InB34dY
maPfKbZllITBhjbqZia4nbPR8HpSHAqcoVs78fYVWH0qd/iYNRhhgvHufxSkzFSk
sPfCKWVcuAamjZnuHPxbQYqZHbNOsycF45qXpS7UaLWbRiC+eNwZ9KkLyG9Wpw7b
jDDz6m6w9LnimB9uFt1zb2X3i4heB5YARyiNdh9kBG8AuxOh9if8RCupoDAXyZgq
Ih4YzgPHrGGimRad/90pwmp6sX9NjyjMx7kc2nNLfspd/ThW9aLzp7u54cm5sHi5
gvYNmOknv7bmvOQKN0az4mMQZMApnF8iDL1bvdI/Ge4bmHZgMi0qf1V8uSLPwx5i
udqhJ6/C/O/8+e0UjNxoZiwQryCsZZRs8IaWU7fpxpwjorliuMcBom4vi80pbi8a
xGpF6m18JyMBXt3pjV9j2eoDy59rUOShkugsd8jUOrzOhuPkGvFS83epoUEvwcfw
EhjimFTKH5OXW2p6O/IShThN1MnOJf6gTQvwAVHtpdGnZf14pJ9TnDcvGV+YlnER
PmNndB6Ec/th/y+s6q61GriMTKVeIBfLJ2qVjhiC76QashOo0rCBXyQcMKPnpWe7
g230pzeFeDlutUzdPFhCQQDB+qLvFI4+4Ec4Vp4JmYKRJMvxkzjcOm1fuCFywJBb
t0ohs8i4jMTwCvChX12PORo+r7k0Ur4rhEinKQF823fJBycvR8Jq0J9J7e2ftAH/
20icmlUTssRE9hxPaNXhiedJgLbKSJBA1K3ajFOb2UL6YI98sWN4kEyZshaL1MX8
pGx8jqWVLB+mC0v+cNxUB+n2+EEk8Ygw9lxRbH4vgei3rYbUn98Amc6rraNh6DW6
PCQ4qCMRtADxmSO8J5ZahQgfc1yQi56lqtmtyzRRgOwl73YAEcSvYBaArbnS1wMf
133J8xMTIugErz0ONv+5my+3dPpuiZjJ5Oglvn5b3R5W21jYyPrLse6jNsMR0OeT
AwsrqCpi90eXbyVV1qyCztDEzojywe3Xq3B47WPJsw0SXACvGPedPdE9H0HvnJaH
1Yon2uedcxJ2iJUZU4KKwYW9prYml1yIfuCPuS4s4XAZnYiedXQPohXW1DbSWvTB
5JRxD+TIZ7Bd87RdKEtXB40HtEOizYOKt0r/8a/TXFBfCwiGftfBwJnxmhXQWQqu
gzdDrv+XXUqRINl5x7wxDDQaH+iR8UV8QrW/wdSL4Enwk6pgbMbE9EGzY99QX+O0
6Xv3KDHVum7kXbBbjWYPOFuLZOYmOYdJ2mHZ8/Jtdn7PiZLY3p5KCeoVUuTIj+9R
WRmvTCwHsTEN0PWdpHHirV975OmQ6oee9btswfOrXMHqCxOlMUM/1QPwxhWdJwmK
nyz+F/8okaDQVPJMn2c14Sw9ESL/osAehlzoKOksr2z1gH2RyctPWBqcFJhAsg5s
wcoKB6kIOlO/gfhi0wW2m29dSpihZR0i5vE2x9nNWep0/qajhHCAvK7Uf9U8DOcG
YKGdmfebRI5eAigWMpiwTsuXz5wQwqx/NyLrYPhu++oWzSOAJKaEncP3PjX10bbr
8MZLQZ+fbH7DkVGUsy9qFF2n8uvXWpQnbkjYZHckyZ0rKxmhf4kzNcsw+97C0HkL
B4BaZoHmc2RJc+0KsIztbyusyPnyLRCF6kQze8cAJTlcmHholygOemDY6aGlCk74
nLSLegT6MHwKjJArP3K2GRZMCulbkQfaq497dXj5Q8x4gHQ3EfZE3FCAhtRVu5iU
/iQZOEU2/b3dQu1w6cptkBF1Al9IV+tbWGbZVT3iZX32o98Hj/WMqRAigZtk6OJZ
wUhgoc4BGxcKQ110xAYSuuZ6/OI+PWLsQXjrvIV7h1LrmoJCnhI3AkruUbKQ+BtD
qnslVfqb4coHChsMO29bt3v4XEe+O5cfyFCg02Mpf9qHURf/4Q/TTrU+51VvU1jt
YRfxONIaq/hwqdIaW1rAg6YAYo4j6Gv8oFxllZUWEBqMIJnD+5FhAaZ0Cl6HWS3R
y7yNmmV0JCZGyOx/XBXOxsBYsGptR6ctBxgBxCFv1cCf0JMLz9y+bhpPoj0bYgq3
WamtSvHZv1xVuj+qxf7+XY2W+O1IJ38GBoaiUejLq3BLBtA/STrJCl5EabIw1qLp
u46t05p7bYRD7DByYvf83wGXbCJBXwfoVef9L2UEN2waGSry2uRqkD7uwQyHPRAn
79Q7hgr/y8u39o2uC4tC8bkYlv3codZ0E9Aj1FhFh8yLDo4kz8EANiwoSHWhsi39
8StEfk4jgnF/L0qsjgH0oJZFhVXqhsWTqzFGwY5M9Hee8znhZEmIsNzuxborwZ9e
eO5X3akf4vc1ioZmag6P6kaVaEvkaQKInXuNRSLRg3/Bj5HN+djVroSI4zEi3M6I
J9tQkZom3fGi6tv2jxeu3rr5J6OitaTkb+6E5/yoShrKpt15EUeRGUW2RdbxjOf9
fJld/b/W9BFUvqluCfBiM0n6ZJ+gB//AYZSDo7h5X+OSZNbSHJ5cCk7ACmwxKFYU
w3nAXI3vHrGn6s7bFdmCIwCyVSEfsSmHmFaFPPLa3m9Du3DU6rnga/u5F+DYkeFz
iDmN5vj/6TXFO+uKTgTOWD1MVFOO8IKQLQmHbS6NXMq+SuVudJwmnzXOxBlRHgPp
QPvY4U4DaHMbkfm0uuxJrULy0zA+VOHXnrlByrVNzYmm/3awL+JPhvP6vHnT0DZd
oZmY8I3oytmOHSgX86c2fSUm0iKgn+50OM3amVzWSVcuS9AG/Z8EGQkOGdM+yme3
mhW/n5t1cGab+X2bAdEjnK1OalTje7uyvp/xytMJp93AvvRFjDf+jNVxo0vIKvn7
x4QVwtIFXU1yC1G3yMP9AlQ5SEbrGkffFmn/wru366C0/HiBx10QmQfyx4HRT6Vv
8/QXE2wULklM5eMcjfU+sIcj4iy3aCNOi9VwqHzRF81RGmXr62cNyHQn6T95DHIp
+3Oi7PzXxn7bY1L0S6neP0Lv8izApmd7D1Yd0BoPI/qgDRIaa1H9a1DvnTWuFAge
EyoF3+rDXvZQtABJjeeeDZ7KURuEzAdV1kjkXAbMRthkGs35WNKWFYuRP7nuuW6t
LAb1B1TNY5ceSkzTQByJU2r/QAk7mnh554kkvXopB73JkqW/j1wNEM1VQMvCkjgf
HDZcPJ7g2nFz/0fMlb5ruxiADynalzqNFttM4MuAml2ksjSScrTTh6u44PMiFjIW
XADYenbfbGZ5LXcjVDk5UVP1b++VkkY7lGRmAKin4ADqTFkXdMXBIKoS4CPrm2c2
9B15ydIqctez6f5Xiiwd0IyAmcfH1Ym27SejO+A/bAnKBQx6osewh9bKP9DptS7P
DtrwnmNQ35vw1h9S4tGeagsrzGmXbJ3fhsMLIBtpcJOxiB0UjHZvjWSusJ+R1MUI
05sy+DH2PHvj3gHkreFF5fufA8xjgxp+lpfTWvUIInvFL2PwfrLeq9xMdm/8+5eR
X0TeMkskc3vGa/to7A37WzD3imjNncKMR28FhEymk7/wmPb10ON1D0xbkfFSUAWx
8SnBNP6WAaGATyYr9d0DX+UI+0x8RYAqyLhlUvYbX52GcXw8jZH9qLD+7ZOPOqEs
Wlz18QynskWcBcHiTxlW6tVQujxXkMtEHpU7658xPt8ZSddgn7kWgb02ZPenBuV2
kE4PYTV8y9tpUJSlzsQJ+VYqb7Qt6S5lwjDx6PnLWrfcf2Z5n/dgkD2zZVNgg3jk
3TNxYcBgkPYGx1mnYyPc5DbmyOylv3HxW38o9yMz49CZgAfdSc7OdCia0Tbk5LHS
IYtGfj1HkJjGojQcsFiUJ1AFuv4cvAIlkC1KXndCvjs4v7v3LxleUdJ4sQmCGYpx
OIEpKCzYcYWIdDksR+MwPl1kIJAgS/rUpj07gctM4pwi+R7Y249Fz8FCw5iy3F01
fBgfifA865wPBuzKybUduBvRA42hqwsfGEg+0/hh64JKADQ0sLC4jFeO9OqyR0Qg
HPHugc69QyoPLHKiBVQQVV79LWHn1c/uMghP18L7Ax7zalal4XWMtERl7xkHOMZY
DVbUOTlrEkUk+HBjHoIkBpYJ2xbPmh6BIOtoBPgt7U9bTX6m38G0KlhEr0Z57R1V
Fs39Uy4dUbWDV02XiLaqdMqhBi0ifUPNULhuFTR2q2EbDhmVE2XycSuke71Lq7aS
he6xpU/cn7Uiv0xmYqfi3yzUU8fh23/duZQM9TKKu+WWx1b9kbMCNwjeXU8vWyOb
s5+kSUkqRrknz+3VZblQiINAlrXin1OVi7fh41keRbtcs3Hkp72q2/sUQ+rpm8hm
vN8UDdYMu9NU9qnEJbzCkU6hp3djEExdopaP2Q3nditPMOYWgRfFJPuMuY+WtMy5
1m5YAlVezaSy/DC7kygX9ATacA+mUb4fXopDQYRReKy5zFiRr4kI9iUMZSp/BFd/
wyYefUkrhjikW82uVCZx5kMIYTNtHFN/MJHJQE3fvFZo1X4+dHfBwpuklxyCijLP
lSsZ/pUDsTJEKsZImTVSOLZLqcInKfc7iAOb2h7bQnJdZhv9czGc1yQknF9mkTAe
XQ+PxlkdfJi88duoGGaJ54MDCwJ0LdnXB2vYt30DCIUov3MPczq4KMBAb1oCcrkg
YvSezprAtf2ahi76HM7SSpuWiglyP5UNFfI5vbVKXlVFveIasp8AXpTVRvi3fP/R
TXQ4gx9K7vQ7EnuZKGSO9o61H7ksDUAHe+n0jRTIM7kKDByz+hz/dDRv0xpwLjEB
94KQEdNYTzMQ69NbvoCDse1+PLMGfZOpZk4XwMZ630tBqxzLKHSsIMU9c07ROMB1
Ahj6sYLa6d/nVywqNedh5fUatJnXpNzEBP1xFqrUmKShHLMWq3c63OgXSxL13nWE
tl1Rx8SaZoCaMS8zPYKFoVDAC1UsaOAu8g/0qtNZytxL2rLknVFwdipt6UNRZO0v
81MhrorfymOi/YTP/Mm9MYrxQgZDA8UiCqsHigh64R8tNekR9VnUzSfH+5Ec7cmF
1pzqiDZJxHdss7z7IvzCzKQzUEgNE2Lg6FWSNONn1yo9yCO+BiB+qffGh2YGZhZi
z4P01Hri/+jBCgmacVvCIrEEHnDe7TYlJuvb4FGWVYpTu4DX5ntL4TmV0f2NySv9
gUWVawN98ZWsOedmFOIH8KnxF/96o3Z6c25Jr6hbWvD3uKxcgYZef9Qs1GP1lWy1
DlEQDM0otuu4wUu0prXLfomMB3wQmtCLURWZkyM9ssm/Fisak8RyaGm4+1VMrNnd
0Pjs9DOP48GuaY9f3tFGJ3xXGSO8DrVakugMYzdBOAJzEFDSgF6EOYj5wIdShl+x
qU3b7LmlXzWVtoG5UEDvun17C07M3QKbTZotIsbZyumGs7BMe+3C5ghCDi/NN4VE
5Ikbf7/Yq0Drj3xhmoArBYDZv6ULRd7NtzOrU7e5jTmL9H89l5hvUA14wOwKZV/1
7mjJdaIavYLLNqukKue90w==
`pragma protect end_protected
