// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
q9BnQWHVms5F+aXUDj1gFhmHb/gvjy2mTJWpCMqsNzk+AN+ahhHvKIdRujgmEy9X1wFfnxPgzScO
O58hsd1ilqtXrZjCkupUAKXUK/nt4v6GLY6//fw0Xxu/K3ToIjuJk/WHyxN8LFFIy/36RkVMANn3
VMIsgNa0H31TI5S9Ru5bVSzJTdps1/VU/yWqTHFY5UI8y5H2rwuJguBniacTtSX64po+jolsuOgb
b5N6BMEMWBP2aKTlZcOiKCOM3YXFaC+j/U6HmhrTJKdC0POoyZymq20uNwMBm4qjBeu75XTEhMPm
b+PoVChQ6zTztfCWz2MdYvDabrsCGugXWsLAWg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Ck55bCuOg2ZNEQlF2Mf0reTZD8vG2ZOYm15vj9PrQALoMeDDc4pUWxeaA7jFXdb2x+9/9BcmF14f
ROtbdUSnPjclxawJ+yx6zesl5am5Lms2Lw0R/YAlzlxf1P87l8pwtObo9n/66qZAPhrK3w3rozpU
dPRQYUGVw2usF7COPiIZ/Hy6YJIB//rKF18yEH9LCSa/wbyG+yBk63YvGpbXJJ0cE2ycuzSnrHz2
31+u0UQJ9hLc+uocgZ3rgX5lKzazne/qcze9GV7U/yx8j2XxUa5xWjus6+SZprVHc6BbdSLOSEmO
OmUKY1+2A1WD9o044eJgRiqS5MCDOFnXseb2N9Ol+yV/1QtQdltigyxy4HcmCUO6yiy5xM0yB/us
ThGM86OEFzt7bfah2pfYO+dM7Uv/aUZ1/m3I4K6qzAWCzvYgcF1HFZ+Yx+SAj+XE8iQu210rGlqp
vYA4KaVjYhT8s6teoKrTIL0XWHAMST1kEB0a/94ULnBeSw5OBnJI8RjfiP+T2twh0pcqhPPxMtnu
z4L15VU9ClYf3hemmQaqtFSMNbmvJbN1ZA57hwURIIJPb0iXJ8fybk/lrVFKm01eDDsGVtkMmWik
agQbwTDHm4PxQAwL/zmKEcWJcP4nog4B8xjIDB3smhnh2v8cgg4/O7YnJMg39arAnEI93ldl8Q5s
vAP/5Zd7XZD+F3fPk1YPIVySWx6MEseOOMCDToKlS8k5H735ABcBonA2+jkyNloBhjhH+e0Y2n/N
5l/gyml/XPTD9ju0uZG2NVQI3q2FyF3bxs6vVMX0MOsCvaA9LAeJiRO5W2uCzVNtzljbSdt5ua33
KGh93/i+cSkfuEiCQ3k4ILezNtCuZe8+YhkFLWHgkfEYwhRVYPQhKdet4k6HcDN7LPR3lbwOkdH+
azPmmrepM6ZVdH04pYmbZU2mRvWwaqnnegbuOlIhwqSUiNccmlhB/UNjT6jFgLLkWJ+yV05b4RPD
WymvTnusXfT8SLJaZQ2sJMyQSQDYxnJ/o5v7qxfC2QYxEeL5vTj9oY/XBbahL9Ql38IAkp/aots/
w3KAvUPZ5ePCcmKZipKr8UqfoWMlyr3yixzlH0uk8zsj1Thx8Akcj9wTTYSxcCo1E9Fq7Gra6VS6
CKBiva8hEUiaCHKn41r4qUgPuoxVrsPCbUEFVqB9Wdm0uRkck8+WssdNeGufqBdZ3Ht9wAxznXhy
RyYHzImPbE1dVhXqm3aKCrDB/81qWIfmpE5A3OO8bxnJI3KvXfsInwFAbiSU4083L85sMNNF0kDE
J7RuHHFKtNrsjreAhUZVqo70udve74eHg2xRjFFfGRBoB5fDl6+VES3wWaXopH54UwBayotZaKS1
8qQuqfA2f7VPxDOgcVN64sTjN6IbVvcrG2VFdQsSJfAucOU0dsgwXjinvdYefqcCJHLVVKH7uSap
TKoSGhJqqqVLgQqsWCA3pyJ+qjCgc88qHqVdL0lrstUgwKFGcYNYUldJS0SypMfCs6LgvgdbAu5s
o+ich3Y4dZJaIUkppFR5XDZzk/MQxZflWxZBGYXubUHRWb2EPdD59WhVwNfMPJmIAKDFVks54X6t
2OpxX81fmmGy59C07COnMasSu1DAI7khpIBG7JeZv4RVynSX2RbIYzyIHiAgwDx/L/OoXXTb9BbM
NMaxgqHA21UXVlA9uPFrLTiFCM4Zwkm1zDyEyNUU7aHi1Ze8r/LGY0nfgzkAcio5FOQ35Ae3ujJl
rMnMix6Khj7Kp5eOJ/1mRggoa5/mKnlW7h1UT3D5Wk1RjlKvAYanzouZzrL2jg6u2mTlgu4gWBee
Dv11oP21IrllWPU9270lyKp+yU7NTFO7hVF5R9eT1l02bREODmYPtVIOpyZD9iHbTBwMR3AevzAb
0IUgdqMNakskH6SbeBCwYfmCJhOwNmFR+P38E64DLbqF4ug4hXg8YnYw82nDaMy2SuRBy6cdmZpa
jqa+ZT9sJFXlrnYaHQlNhA69ID0A0kuraLV2Rusd+QMDHcAd7BqP4Sg7XJAcDE+TF/EO79NzYH3r
MG8FfIxoyYPmfKgWtG5AKPs0JN/CPgooWDCer3TRGsysLOr/MT/+QDwIkYVFjp07neTQyoNasgOi
ObARtC/+YVRWu+njxkwLvG4Qnu7li/pGek4Q6ZoQRZpNBX+v8I86CQ+AL5pp0th2gbREfJjbEUv2
dq0rjKQBzkC1tePxE/efAvU9uiTrsJGLN8l3x4t5plf5aYOmQhgMLkmO512Ht/XpkmAzKDw0P8zY
uANySkB5cxsmSDeKAyNGjaLEhfTUhQpRKBJvvwTf8w89bBCFQQjdN8EovqsAfxOZeQUywKT70ejC
FOK54+5rlRcl7fvM4hKj8MkQ5EoyONx9tV7M0NI7klVChfN4xH6DGOAbV0nq33xss4upgLrXmUi4
v4KpArcHhEk9UUeg1dVvl+b+1X3RuT++HsZzrig29Wj5RtgHzAYqOqoOGCGB7eqYepzO8pKC5w+k
LnggBdqQuZLAPK1KOv0lfJz4WtY4KzGME0/gpi+yTjmKWLp3sQ3GOnLmZNF275zFHVUHToks6YJy
Uajao6KQt/k6bUUmgColw8WkEHipcqMVgKozQN59giWkxEou7wSS8NEllLqWVh99mJml95COec6w
WQeXsmUgihJOvlhCep/kKs3eXxAk9vArLJDMaL1IShEm9Qd4OYrpNYPqTeGQ49rEAEk1HnFGlYPG
hShMDN+PxDQqBvqMuhtCszB/BXQ1jnvyC0Ok/lYKQO/ZiGcT/1WtgSiiqC1hosNpl9YiO1dRy+4R
kMw5fFdb6t9cS6UCW+WyjT6AfKaMOpNoE/53QuZB1ET/SVHqNssOTp3pEPSxP6IljEwVCIqFkwCO
SAIJsqogZOOtKBzfYbws3a//ypqJpZ1kx5wNvOsVeDIHhFRzBIzuKmk9rN4rSRFsTh6FkVjc1NGH
coYnl8pb1nGLqP+H8UR1V7Yr0fYb95xUOMezjTtcQyjOJESpg1lN4lOw+ukMrh8OP4LBOPkCW4wJ
j0dYh4mqHhfufq1V4pOuG/jJ6N2guQJZEgXgAWweKqfEW8US/5qf5xdMLX4DNw2N+4SpJHTjOSRz
NdYnEL1lXNQ8QzI+Rs6plgmkpL1i/peF2bIkASA7Hzp1x2ihbFoXu+4O1QgFFReOGjERXNUmozXJ
LKYsidF9hIUc48POjINgObGktSy33NJoTtcpS+gJfv4OTcLu3vXSZGPlOq1edxwao7OCAvkck14l
1xAuTKRbSCa9tnK4S7+bTGp9YX5Xdpk758olNNRMcrlsSsBDHf8e8AuUgBHM/IqQjEwBhcOy5wBu
dhuDTbznAon8eu1Z4SidvkO/m3vPCvm54MFMq5o9+OqW/8nXhDPtvt5MEEdMPYHBoEuukVizv57F
a1pYNV0NweOlXj3l75czV6CbuTfm1VnixX4LHTrEDmOkFIW5JNF7fGyM3t+/mS6pR92qi5m1zPlr
UNDb6CAjKd3+7PcPwKUOIjOEVjlVsiQGDIkpQGrD9H8Zz0vQjwnCGE0If7noUmZImWP3AhOEwUwT
7iMKRSa869KpYn9qTxhlNrDKA7Zf69UpdzuNzQlTRMzrzXj5KfSWq42UNOntjZhbPtPxFIf5u0Yf
Gh+0lLh1GEkES12yXVpV4P3YSV5/ILTrcLjQA8wDG4N5M2RSthNcfgt+CLdF8r2LZjIrggMia3nX
4+ZXk2kNv/8Vnvh6qjt6ynbjj0bwavgHx4w7Vmt60jvE+/YpyGXPEVILJ9INFNPWEkxdCC4+YeBo
6LN9b53O92zYywFg1rlZaEuqNDb9+MriKP6gFik3hlbawmx9Zaet6cmqdne/tqiBWAno54eSEkad
PTR6m7adQ/EsBN1bCdVFh7Fqm7wiJpngGLZtQ5qmWriCiINg9HXTmI2tu3AtPCvEg/EfWsxmTuEs
EOZGQqo3kK5DzeAGXlYGEYrGJu7sbwUm0kTwPJf1fL8HIENHPbEJnCEaB9SUcl83RyY/QyX+t/LE
HUOyRnfXNZS6fezfh4/pioGMJ8AgppSgVUp6uz8cgo7POuG0WwZAQNIoVw0ssV6lgRoYgU0+WO2w
esq8GTPI7JSViWBIR5MeV9vY2u+eV/DstRF+94Aye/jn+gYSgChc6m+lIqkonQjtusoUtY7nMB1w
t04hd4e2rSJ0VJF9VNEb3/XnC1NRChz1Y6huUCH9MvbeTtXEOjS/+DeXWIJgEaWxhW8Vypxq8fwm
fa2wC2fnXNbpYHWYHZ10Y3+YyPS/kqsHZPLGnvquRMbESILCuuXLLuva98+AIgHKAq++lIm56go3
ImcygkP2FEKOGuXuYAyoYVQfpPZNIaWvjVUJ0P5Urwzb+UegYqyqoKfX7kFyWr0yBKjCfFWLTkrS
WTzsnjLU/TQdtEEwAanlnyUkknpdFFuPba24QkB9xvQPhbBZDT5AIN4o83iKgxplo/ApECszk4lj
Q1TcZakrOVTMZs5YgI78I9f941DOtxP1YljmrG38bvbxeacvx6mCrOYI7njGySBnBUKVlh8teBiR
F/1U1qdz8Ztc1+g6BgXBTzSM0RUhOdNI139rm1Ik6WXBsoM+DWnAIS1K5Ve7essyfU5gklZq0ucB
Mptxz9FZE+iw8VJDK5C/Q/SaMkjsXk+keZ7LQCCeyU4S5EggrqWkC1Sfc1p0pFLpUJL8pLlsH2EH
NV+JUYJQBPbxei0jN50YX1+raO/E8WeB/bhOnJw6+TRZ6Wka7CN2rVy/Npb2nmAp+H34cvu1DTuV
mA56q9QjUU7/dJq0XPWRJvRxpiQZtSHkzv6pAFOn2W26ZvOUcVNGAIVTebBmaxiMA0RE7RyBBfIG
8kVDRcEeRIMIWX/LAOPQB30Fh+4l1teCOwfONP4zy3GSC5cmYyzcv7uMgGMVpK6ZEphN8LAciBK2
NmQsQFUWr/Uz8FMXyGfVMnpVyFl2cd4I/oW6wUO95sdm8wY1VwPK27XKZMFEqSbV/vQOVHy9GAkX
9ncw4wq/h4py6QDRKCEjc7iGDSbCanUQKpo/W1n2Y3a2mh6XkG168tL1feti7XN1bTgHLZRvknJa
ABQ+hGC3fxAaQ6pzu9uSSRwniTwetS3mO8hoQYOLG/75H4ZwiuxfKcwrapfSCFhtv3E6FrCgpbps
66SqJc5ICTJLipRtUlfmNvJR0Ccj8ULv3mqFm170q4pZc8VcnFMGFBF9z473oRGijTQuQeAM40Uk
pxYFBxa1/86DsyeRz1lcs1pftt6ah/JJAkEbw+vV1pDT9kwIgjVClzMDvybZPoxtnjNcqLjUM9KQ
BE+/pt6x5mEGRwBfWJQuryeplrGrhr+XyncfITQbsM0d6YPGuKSaX3dVo25VksDgtGc7Mf2BkMrK
7E4l7g7jAZK8dwHyWZ/7HjxtQNWt44OiTGg6hIHwLcN7j4oepo6XxmV0siWSRX6MCmFkED4Dv4PB
nE3nz8o9Dhfm80rwWGWGClhzepRDVFhWLsQgO1hvyQTx7RAAhG/kNpWIytycu7GrR2yYX8qppENu
6iGi7SN4lGKLEqnHlM/Us90OErLFtH4k47Fp4hYLREpk5T8I5Dj8zaCaA2C2MNCAfeR0XIh4toJ3
2ofCxqUJloGCAyKsm1V4nC0gU45DUNN1ZRFZqBrfTXXR2SUq9Gd+8/VwAYr+bpOOQZgn09VHjAFZ
kt1y//TbN/SM/bX2Vsj3eihtKUhINFvqUkFrDeV3MMsyZXr3C0Lr9b9o4pQ5o76fRkZDgjUv0yTw
/7XXHnWRJyHlt7K9jlLxuKpD/xTmyL6bg8/Mc7860L8RR6fXcPkvxmisDOWiAZA7nFptkjBbwoWK
GpPHQII1SKrFhxiA6oHYsipUOyHMArx4hpsut8LOwerhcNQsfb1bCvitnH2EDo7kwq/7a/Xffrw4
c4SDQye2GrN1tFacUmuFhopAc8URdlH8qtJ+lNnXfzkT1CLM4GhAbZ0eP24F/b5CiV8kL9wC/tOY
RQl6gK8pD/+R1raKeI/dxIC5N45WFmPtSvy1GpSx98c0oUfq1YvjKo/6yp3I7RS7BqfBm5UQOAoq
mtGNoATFH/ZzFO9b5QkCwsfC/J5JHgZP5WkFxS/TIgsNpuzY7+itZLvjCMzJoVgEsD8/lTySa1av
SGFky7Tr6wlLaFf+dy4nQWh9hE2e8hcmDVzzFCHjR7Yq9xu7gd5nXL2RoytT3qu0EK1J/V4mtcmU
f09YiLtoa91pWYlMrVZcjS7j8fEum1AQxdzs1gBOOL5134SeWCH18ldQ+JLVg5BR94Wo9ijGxdJH
jshN5kTb7tunaZp0D3o4HgN6CilaatMj28NPmTf8xPQcG2jb1pHRTplurvKUn0A0QhtSmFup9DiR
ymkyHdljX8BDIVWvMoXMi9fu3BTmgrfyKEZnWjwZDTLWzDvXAyiWWFWbfLrxdx6Ss0qFG4BsCcvk
ZNylOp8E2+ZycwTGcauE9fpS8FoA+z29iBxD2j1GamUpU63IPOtm5iSvpbkCXlsqg16JBbAKY2O9
bJbOAjLeGnLEoXynSElyuufFlqaHfNaCP5snS1BxF4hieXPt4WPlZhh5zj/1CX1AOZ5IG8CmHLHo
mQzg817+3PIlbRsjiChNA9X0GD9+xt0phs13iVFkjUuic4inuf5j7rpZXRmR0feH3qvMag66XO/B
46/WtkyyrAInoxAWj2CaeA7erP3rMf1M+oNE0dB2s7JHt63gDfvVxS54B2ZMPkROFvldp285va6g
JkfxRbOkNT+cBm5Dyjj4Z+LSy1qP09RxZkoaC3rHxbKsq0nUcHGUzbyKFIWXB1dpWPrNsP0nhq5s
2crXrAMSMZKF2pbDMeYHxjg+LrUJok7GO67EbSFgcqJM7nxEtzAg+K8mxueLMn4f5Oku8H4KHCnZ
w/Kwk3l3hYTFC/96lNYrO3jnrVQuKICRL60+KXdeuTK9Z/jUz4EIdPm0mW1JvfBkU098y0yocEG2
o7oYe/H9yVNM2YEZkoDg5mFJ0LpzWJCtoPoFd00kVL316vb9gEwG20LYw+2jEorPcrC82t5dNeFs
oRCaKjhwY6RbKOPxTcPGZngDbHvvZxCqV2wbOI89R5ZyTc7DSfffIw4jTqHGEfAApv/ZAyEmlmn+
08oXJ1yyi/XXgKrniZTagBBPc3AsZFf2lrOecQbC3PdACUQNXPq4EEwGKZv35zrtk4lswnvhtsjb
Lt6EyveWEOScWopBiDiPtKAMGrFP75I/t8mtECbNbZ2/1O/2rf6T29iC6ggXYIKv69ezSmvQmGuP
B0pVmEPx1tVfjNT6BaS+Doxq3YDgm1kw5GIt6eDAZQUYQ/503oZLlCnJ7N4VRc803RNXNB6ebH8R
cRyjmTgyHOOWSV4SD6dw7tC+2YK/kGPtBKRi+1qRZ5QlT0XeDoKxTUgbzv8MTdAnumSsj5RHDgq4
ngXsN8lPbImCR//Ew8wySag3CoqkxXLfHM3YtpsSbZ24tmOtweXtI75rwOFzoCcgV412qO0L6ul1
7Z8pwIT2xVmfydHWfNkcBkfe5STiQc2xMoLP+plhV8ZGmr8zSoMhEfFjreVl7u8riygUe1/VYMoh
FCHVPuSXcCqQXn8OnYob6sXJzurp4IlGBD8ofeAW7JjS5PBIvfj1QkO/CmHRpGiKROd2D0gnjI4p
lCJQtHEW3qvomrvgCpZ0cBcUzqj7f5rNKnaXjI8MXEvbl2ZtWkAlZ3e1KY0Fec6ZXKt1q82eIDaq
k99SpXeJXgyibb1elehAnb+prtx8zHLkBO55vxmg3fNNNNjZbT0xwx+xkZzMlNhyaCrEjIYkTj8p
PRrGnPpFFzUUAKuJmyZoJSM0j4cOgK1u2k8cLh0zX4DwLL5X/zaFZZl/DX6jDHduDvdXleWYBS6A
Rt6MQIZxEoYgSFQ6nW9gLsbp1n+urdQMTAUVmQxHk2mJEKS0SJK/6qPxFDtD07AoQ/Md1xt/9L4i
bStqY4MR+wHfEkruiJ/lYWl3dTiLqRE35P06CbQnGT5CSAYyp2b8TxGW+FRGws5nTiCiZL2RTZfO
Zxs1UqQH3j9OtaX14sBYWEPVgxyy4uKq+kOJcmuyIC8bQZY0+PIBuURPDBboLpSkn3DzxL/B3ZIs
IS6EQtyDBIQnrcb8kV99xP61IYCM4zF+EcMjIlHlhz9myXOctBoUxU16yX+qGdNG5+CX//Ia7XD3
0PR6kjk/IgUoQaLIJtjs7o1UZ6Dq/9a2Bwmb1zL9eVm3g4vtm/ma6Z+kMHI3B6Qmvmo1EqyNnjMx
XqQ99cBQYMwy0BANWzINfMo0NoqGUApfaVzT4ihEIuzbGbVgp1C0x+FOqpTwxi70UkEV8vUvifQF
hxIL2j62EAOsjWi8lNjw3tm4ZhZmj+Ts/BJNt1ItWw9gVSHu31o9DOmpSMGBZRrdZkxW5pUlMBpM
fjOC9N/oiAHFGcUc4PBqk9wpAuRgNgfg/DAracJeF15u0dZdDG69xs+g8ziyfLerCE8l7A9s+vGL
kVioX1jlI/7bpXY1bU7uSZV4GH/eZP0dwHHjTzsbUUo3G3WT95wCkGY2lzM34jscrRexXyL7wYJK
y/UnRxogftwiK5YN3p88ksFv13qQ4HscSA/iBJkQwoVfORoi571F5lmdyCoh0Kj/Og+CLVxOurnX
gKN63XZWmii0VhTKB7KNJZEyYNnmyji/AGz9Tx9n55nlJhTjwWNxvAbiOf3P5elMr4wiHvQWORDs
jKGsXEwEiITlkXSMQRWsi0OfHn91MNF1k7NZyejQvjsnPgAKjr1Ee15syEDjdx75kqNWatmmesgv
C/yBWQbBav4s3ieP0Q9pT/KeBKV+BkjZ/Ecr9nnYVPmvvmqNiEDMV3XQdzQgn/K9mOqQZMltPC6M
EST7BjwPakrpuLUqpZPzPu/K9Hz8nQ7/DXi5hk2ww7LYeXhc80oIh0APTX+cCTZK+88aw+bvvBzH
nIb68vM0BDJji3X2FL8ZAlfk93jwIXtbopceeqJtiED8LYCqrAMuD2b3UQg/KoqcW+3kk4V7BnAr
/cZJ5EzDemgcuJEg7FVKDQwRqkw9uBPR7Q4IMcjP5xODE9z1Y6x5DLtMBrLWAUY4LQp3/mXXeAci
aCpANGwTDu025Yoj1kH8EWifZfFReoyaVCEVOzd1ZalfpGCgSTu/5wUzycQ67/IZZAHJcwhLZnnW
RR/rgagowse3rTRcmy7GxIpKd1bIVcYZNNoPvpxaoRSEUchT62cHZqSo7HPTiMD5ygKEmgNGvNBP
52Drd2t0CCGMj0/nJnqawmtOTtmU+FafMdyQf5pBeFwNVE47M5/dvIRlSLRCsxHMpJxI6i28Ylf+
oPhuRYNfBsQI1Jo8ZnpG3ls7g+vvxq8p/xzdTzutKzgrmA3QH7HFxm8l0Um3nemQCVrvawjhs4PQ
RiCsHVS4/9F0h/XfIi8n0CG/QDkW1wkIRJQF+5Ql1dimYEHKgFdm5uU9jDM3NeqhkideTvo/Q5SI
d9CciuuoNZ1aqFgDJ6Obfb26eeZSshe6Qfl9llzbtuEJt/yodm0KLUGm/hpXb9EMD/Xf/cw1zbE4
VkSFuUaKiuklR9bk9ZWFVebNiryYP8mBBFFAvbEIbZyxQD+D0AY9D7jRUlLAl/x7Rumewnbi1rcp
g5mETxoDTKGSYq42uBsEcNQUIJuVQFX/vFOAZh+rpnOyAVaJR7W3kFrm8nehckBHWUFAnqFHRWaC
aJLJUMh3fodm3j23SwgQ6NwyYDiPx+YKI2OLW0w09isRHQac9P92MUjGH3UA0/cNL6ypqWGhSZhO
rC4ygfxri11SkLXurGEonoXZuHs/iDltu4TDWkzMlvUoUKSaHFJmvmSyiWqKL/QqD9Fokd0+cIZ1
vrJ/RctIWdRU8fDzo3jK3+ju64O5EjgCQ5siPe8mXUzT/1yK/k+nzrRatg0xChA/PJqzIIDJym7g
DlEZFgSB622oHFj+KnkiiV6o0Vc/mL4Ain9AtI2rL0+LltUV76JO3/jzTz77wbVv50IMy0QJMRgi
Y6lVie/I2962Ubeu2p5SeG7038txLfDTj/qdL4iG5ZjtV2mlGmiI2VpfR2cRvj0cDIxIxhb7xXlP
jTdBhQscee41Tn5hOsYV9NF697UzSm0JVNI1bYk/ihil65VdT+YoLqpN+R0FwvFO5ft7arp+hsgY
YcbUmUJY5dW2gVi0mKQ2VjEAn9IWmeZVjo54NBnUz4Ew9Rl0YAXmIbxkJcUBz609O80xCi2F+E4w
xHlKAIi2Wnr5ls9Ox+IJ/sNbD6NdLgdrRWHnkspOEO373Kt8wW5fW1Q0HbWcqGuD40D939FBHFya
pxY8x57nmZeL5ORdx3fA8HuSNqEMl+bkgrSJcije7KOexcA2K+GG0TbJMEQ2em1sb0WVXtNE/AUz
PDgUz3WqJtWTiG8ccMvwAupwH45a9pfRWPbUzrlwoO29BeM0jx2OaF0FH30G3K2yIVO+GMQoga4m
ZypcMj3xib8sy20/VIkNGEQl1lo4n9mDkLLeNDQGCr5y7+nY/utEadNaUF1so/AV4eljIjkoLlwZ
u1ewiVZm3o1UoIcRF0XwgxeXltpC0EQ2oPGA1IqeOLsfXPOL3sQqw0/1XPbQYek4kYoIRwKvAr47
z97rVgny5cRU2v35ITQDKfrk/aRI4j89f+ORYYmWvhXxG3aP1AoMUq6LnA9vPgtGBnOO0hUuVuq/
AEoZJ6zd/emuVR2GgRpy/DQY6SLsTADthbxX6ndE/RgP75gJk++FDOD81G3j/gFJIyWPJlgt7sRo
DeoDI4TzpNVzfRKTegHKLtmC2IyW7WiNRoiAvhn80cu3C30rzLUjI4EX9QPFwJNS3w9lvqGFHPMZ
O2vI5GzswWgLvi95muvZoIknRkROXdxpmiNvtF/V8omTk26a01WhdqBb6KOaavu9BKt0D/ooSLi6
YiFYTRhmFQfcpg9U3s4hGpSe+LeifOM/7gFgX0D4jmCjXuXFiZsREiSAppi4u/PFdYle0CYK6xfC
JBa+yrBTAN8QRTUqak7V3lQGtNjjpvUvD0zpYlEeRgQccXn25WlsNYO7bA8x+hsTiAm8yu11VNL6
rFndA1If7Z584dasbRfsOuk1bxlT1k4hPWTOy3DlLsLUW3qtLr7XaekpriAOgZQFKpN+HukYFfjI
nNXacNcRZHTaLCMZaTsBcdIgRmHsz3IPG0SwsW7/Yd0gUi5bRtX3td4MyjC7SmGzBLAJD01RjB22
Y8D/wyukb+FghjEeBXXu+mr9kwrkUAO647YgiyNXgg5ONTo9uA3wmHM/G+0a+ligFteR+WF3N4Yh
yCG8NQagfb9+STKy10x67X48CyXlEeuLPtdnlElFo7K0k+pSMUmGiEWsOx6WrCfT7/rspyh8Xc4B
b2bXSuEynNKCXoqsbxZJUi4D7GWdJUuBcdugkTWj4WpAx48bJi707uo0CWDIV6ebMi/1YyRU2RMO
U5QRbZA9XQM6ZllUg/KjiXINiDuqSGIne8F9E7TnvlN+y9vNnV2ZGGZ//+Ze8s5M89bUbftTUoNb
NL7e5q2DDyFHNcaalmLHh7ZukIolpyXN/ZR5DNVV7PDo/i/qQR+EjNZHeevVdT9gqdpcaL2/8qEj
qqJSpZi58sX8h6bnOCPXEaphxEISO/kP2bQA4uVOPfPEsjlOuSy8GRLfshpoh6ehMNWoS4Q8sEgX
xTarJjsXt7Swqk9oa/sALgYqRQEUd5RpOE+WEhumH9nwpgkxoLUvAO9MVzubq9gE2ftA5xCKKjqK
jzthQVQBN3gG7Jgogn95No4TocYNMBAlKUOs99+1s5x1qMCP/HPCf4jSgur6PfUrzdaLMHzxa1Va
iq0uNnWiE3EMKRrYhG34RS/UbCVpxI+DrI1t9JMYaZe1Sm0GtrUYOXQN+oC2FfoMF7O56Ufji3go
9GyGJlhQsV+d1K7QEOdprkvvsUkkmElLU3Rk/KPhwvNYVqjwhzEFIX74ybHIvB8rAknvP7ZyLIuF
OmPZmnszEeOwrefPJs0ukttSsjKpfnCHtCGMSbqKW1ks7r1GMnJit/j98+ww21Wun4Fihz6aSW08
S7nbfJHqKi2F0dWtGnQr0r2GeCWAm95K+AM1vSY/q6UqbsgYAKI7VdqkkP4E+f1V00davjEXC9Nn
CWHIiqde9O3zkeXmx7f89/zxo8gpmMQ+ZzENpoFxIa36cRGdHFEfHSJ5NU5vCf1g/maKEmJrPNr7
aibAgDzXnSTr80tDPM4Zdv3RhpqN43bxnPu6Q3OjFkTR1mJ/CdBcJR0vBQHN/F84GHdPI3tKRKNJ
EpV3CwCXRlBQojL+WX3vr9x4rR2we0ym4MRmrh+yBD2IU7nWAj6vXLugtMXoDmEraps5iWmUHrKJ
pBnRnqidXuDwLyQnnPrwC5i9m8bsKKFgH94WblnzoYIp7vm2M+tlEcgL0rWiEIeBlrpAKYRZnNsb
Uhp3aF8cJZm0/pkTu9jiwk3xnZ6uCBDAfZ98npfqo+0gPQMQZJ4af8j/Rluq/aWBkbRSOwL3GKC+
TjT6eGqJgi9OBKp3HTGJx17h73yjHfMrsFTfWlgICZwJEjEHmQYaO/CIrTEsvsJLRSrqvPcAMH5s
0hU5g6/QBUi4pB7/MWdeP+y8VLPSBa404GQBmRImKsoJJRBIXmeEuP2qva31i99zJpjvP7+qlKz5
xJlq+rUQqAKpwtIzR5n3z1dBGtmb+XKy2/X2bpMkOeVF8Fg0s4Zsl/IbhJiC0he3Xgf5oJ5HZhVs
nKzxuhnPLpfD2bOdhuV4HCTJUJndfryExtryVE3TZf5hnW4zdGHvd0n5seb9v3mpUZrmwlPatSup
4WwpbTeN2jpRuIbCobKrqWX40UStXv3BHYoFEOrTQi2bGyEBOXv5J6o3eESyu4FBKr/BVIsELFrn
+V1lYAM6ywyNciNyZQqgXKtiEyhEM6dQpZ/FMHt+sQAEvoSLuM556QhwrHYkPaeigVoJaG/SR5Uo
VF34t/2BaqXtJkSILM4C00iA6Uk3c9nAkZp5YcXMwdWa5LD4/p0LVWghTisT0ypUpI4CHFhc2v7I
oNyWK9b0uRCeyAjdnw6usJWAN3DWO9tUOXAWeC1n9+QbKLbOB4D3cnB21jE3KJvSgHZc/wn7Almf
yuyErIjDvcgKyIGViKB8sYttHsFqhrsx0qcdjaLcHU9309ACopIiYhC0I78GbcIkj1Q/lT/RQrJu
QYW48ALbGaEz2rY+NsgGIJBeg9V+VZTzDVioF/13flAnS9KsSpYXo8aBXYezb+kehWJ340U2WWeL
F41wFhRxD/SguKqk1d3eS9ApDnlreL7XrSMSbues38SPQBLSyDykFLB7ELG6/Ld2ng6U2112q7B4
OBNMzIFTTHrFvceXS6kQzAA3oK/+6dkK4FldNa400zfqRLqHdLKV9X1Va9EVOaj8iCYuassoAeOf
pxqCvX55dwvp408TjebCgWdmvUinjTGzmiguUl4jyUpY54BWU6p9wASf4AdlTClrZsvL1YtZqJyL
YSdK7LsV6Y36xFGPnsQyhthi+ZbEZjJ7DVHMen+pyzQc7GD9enQOXY/5oc5DcJabkmolQ/dPAjok
KIQ1MFLJPehpQcPTenMc45HQ99sU8djyYDfs1a+yhgCcI45Zd1KG0f9lj0eEuZI8b/rLVX/JAyYc
IpMzgH6iTZxEaDr5qqRfjz3IJBdQzrUB7p3wFZRHg6yzZGuOgdaQXs8Lu36BPrIKTQmHqJE/qRz6
xX6HaVRerAme5sf7wBF3mANeaczl21RDRTa/Bqts1NIiZtXgDBAxcVT7E4ahiFTEhjYYrcApxnhJ
8JZVdxLwgLLuWMn8Fsxhn4SNloGahhMnPqGl4F6h2zSUXhE6Ibw8L60ZEEt56nbtBQH1yfnlsmSc
b31H2ILI8GDsKydlNe9kiFoZa/GNCfHn3OqpjtbywPytobesaITytXgTjLleROs3qJRbt2ewFO9c
QYfZw/tWuC6XVgcr98iFZuYcVyxQABDbbjHYpm//W4BI9hl/L3u+SFGiK6NP+OvpowXiEnbEJdh/
6qOrt2UVGz3DAC4Af8mzT4M0HOanwjsJx111VtqnkE1S74w5iWlBCwPOLiLCosRJDpyn6PnGaHQo
UZO84BNcxwFmUfsqnzpA6+0feqWRlwFlEdC9F1pvdJ5meWHgu2Cd7ga5yFAUrp7QikSmLd8KalVb
rSU5V67XkS57/t5rcM12TcDFvkRiVelVJj/9wm6H7AlPOJ8zTC6dZXY6qSRFZXzbWDRQrW3Xss1Z
VzF8L0NmUbV+CeRsERV4LarzPTQa/I3QqYNNaMm7EkkzVGkHamHY4jOD37S4ORHhDERwEzIW9O0O
/hKGlurCPLy4qYSrAyVBYBG12ECcy4ckR9LoxdLqT4+mNvgzV6KRysIB1MvSIC/lQiYMtpV9fZHM
IiNIQI6nwLO71W3lfz6irPqRCzvyB9ng3r+J3J3lIuEQQmWWLE3UylfE9LhTNbZVAVm3IhfUYcoS
n+agJoH/WNttEAUbcCatSFxTYCg/HsQz6263m5KtE3bfhgV9y7KftrSpTMQZBzi7DkgMvi/ddDA3
7e+RYLVbDWuUpO6/h+ZPhuKSgMQZvCWl19OiJ9AJLyRAV8FePY/j1dOXjg7j26L7SSax85G7Sf1m
7899awLAkQpiZKfqj2oSXut++CTFEeXq99nLVO1h/d8w54i0kFD6lqB8f1fUzS5HPJG4zdffO05B
R3qLMT+HMILmA1n+yCp/at3oe29sSvKRaVpiCXVS0vcqTZhFUGs0szb2fzxzIbRm0WDJugMVUT+0
gAiMoCVi9mgN10XyU/s36Ubw5d8yx46F8Dzg8PeotTjE8VZHDR/zbpOmI4qbxMlXaOBVrf5NQ7tK
Buxoj95U3t3ZfW3SlO1hb085SF8tuVodU7DmwD24gGf3Gr9iNzKPx/L7ocy1A4G6qKyzmg9sErfz
tCMVqv6wSk4JEDD2NNpNqp+DMwna8Wc9wq6o1Nh1xSBGvVbI1F6meSZQlwCZ97txttIGayPGEKjM
iuQ5F0+eeTlcFC3PbsQWnBzYw/19DSAR4WDkkNDQZVBh26whqHjk6ik0/M59pVkNWO6trieLBYpz
V4cpXHKMfsprhoxP7Kq80AWSG9l1xnj9ck/M9OY5FGJn3jAdAdo8nKNB37P+alEED1rkyEWNwF9a
CE4PI+h01oP6XD0pbP57tNBonIrh8I6KoqnyfIpqNulsOelkWaBHLxuZftrLrx6yIbsKG6W+rjMH
mpr77w9A0Esp9jrsM0N3V5/tXFDmj7KuxoQU8pdrBfGu0b41+ZG6FQRZBka3FLa28oyZdBfvjg0C
sHA7aAbTFh48Gn8TGO7VeEyy7+oMXl8MqE+xB3zZhCpCmEgOLKog9C7LiURprwSLBZvQnfOeRhWU
0LV0P4ZtMXATrQGxgDqRaol+s5onpHoCmITITmMn4aveXP6BUASCe+VaubkSnNnV+qHoILbLJCZz
xwao6bCNuNtb5Roz4FLvQczj9/eObwP3FtkP4WXDypXoh6R+jb5Ps+99iSBowafVDgWBGhUpGzxe
anqsP04E/QGhupGBYzXQbipwQC6BYd4/gp3qtWeRSdgzv+hO3RYl+Ae2hkX7ZprY4fgCvYsEPizG
sCD27GmnjTSTF0Sc4sSb96TkyA/goStgWxF+tU8fxzADi7BbGKWFLoQ/zX7FjSzLdwFBCYcqHo0O
g86pBfTtZhiQPnYCWi9CrcaH/yD5VfET9dnlmxCJ2vY1uYR1m7IeSUrhF+halYkcI+dhizpfRwHL
B/WDoSoy8P4dZpM1pcf4HtLk8s/W2HzlOFDp/p8k2CwI/Kog3Q5xC6JAZNNpVCcZmurQGc9TP3Uh
+xwv7/jfUX14FLUsrjir/nQ6mlarGIstPUbXNYIdyk5Iuat67nu7JLmNJf+Oenc5LfJ4u64xxc86
aaZJlkSXtbFz6NKUWXXG0tvmqlxmG0AonmV+smDqcNBHpjxM39kiPo4KHSN+20YpNtHOG5OsQXCU
eFkQx+LH+z026FMXBV3YngIk0WPKiKQJgpDO+zsmdBftGg4ekyvbKSraLfNiCNyhXheQTYXWTt7P
j1zjL89JybWZYzUZ6tfW590I+gUbqchzWInhyhhPs9c30wDmg9zMel25YgThP/EL/xeUlzGSU7b8
XsoOzfcay9Zb/VMkGCjdnPj4Q/eKeXc/ISGtZ55kKCJYpyngWdVehSHpYjosE/Vv/jYeTOR1KqQY
HWM62jOIhU8C02+kdrV2FgekP7xqcrzNsb2ac0qSnPaVKe0qRegLDBfbxN+7CLcc/KX5TZ1xvv44
SDliiafyi7vKCk5zOuzovKlg4uXMttitCsdY4OUSXaiB4JrbURVvIaRBdl8JhUe7bbgiqFem8+4k
9AW0hNXJynAWslmM6dgLNwigf12OfRf7HbQsb/RLLGBioTsgcyq5+n9MOQKdEfT1iw9LnoiqoCD4
2iM8BUm/KF9hyJDfANSKErzV+ygtgCngVbmXpUOAJnxTgXEnCAjVr/LBoZ8pHy1ajIsUV/uaFq2p
H6M571jFSkWWtPHR4Mau/SwpjuGMk8ES98G0IavPOFy/mRJmcxZlB694tsLESQftLlNx5PhUTiqz
UNTo/lAQtJ7dWSAFL39S6G80EXcsDwE4smFD2r0x2OE28D8dHuL0h3uEqLNPBSlgpK+djrSXfZzW
c4PCKTzuoYyStNpKJM81Yjvm59vyq1SgpE0bDTVD95atn+UANbPlt2J7sUShKdk6a468K09AHr4B
i47mhawAHzsNbgUF1fZNkISAdAo6rqv+t5DzvP0tVZ5kD1zj2LoTrWJ29IZ8K8tHys6FrdYYH3gL
zsRnGl5FLSfHcJP++8MwWaDxYo6PowzKKb7+H3CRwoP3Qwx071fSFk5UMq1I0S0RZqFSqkLd57HG
VrB681hLGQr3cNx2thdD5igOcHUrhGKQNo6NffHRvm2ariVXsXQvrVaMGOv6AfYpa39sdVYRtS/J
qNxJw/s1Y6I0MzvieeXOyHC8tRFgFKCMQdSeLSCcVpGuOn3U2JZD/PCCq+HBJcO8kHRHuSb5D0U7
VcasVjqFCVbJLjAFbMj899B7b2CmOpUv/uLSbs/rXHOVyBlVSaqD4IKkWBxPBJ3m5BBbLq037+d/
5pLEoGbbaBKs0ckSqY525hnBekZviIFczUVIEmjgFMSeBSoJFh+jT/mfaU3693YY7XKbaa5JZWVx
WrC+QYRsV5g5WyyCOb3w8FaMkdvCDjUq44Rgyv6f0001f3y/K/FvlUuYJBHtedao7O7LGjPSMLcG
tdDE+0VhG2MqwpUnqQcXhuvB7f5fnE+d6Q4SrOnXdOubwcgqrfdlUEqeig1jrDdWGwngkKUlMC1Y
Ygd7TWXdrIPH6KxD8cgxr2n+EOapxIHuX9iAubeaD0vT9GYghRuEJtyylBFlBxsphL7em/lOHe/M
EOgII3+JpFeCBJBeiepStoTGW0G39+QVbFa+/9VTe4ndVjibsl5CBz+5ecmVnF7QuVEeHNqCBLf8
vBfTe7+zMSs4visJ55K+QCh8fgNrHktDrmNeUiYc3EiMgPHIg0zW6dz2wf3PyIUs6oyb5uUT6RyW
R5ZkJD9D5eqfHVWg91KCeANsk3Jes7B8lpVIsAJjQMCVRDq9UbzBCX/r47hcqlQ0Bw6hRSO6Bqvh
CqIyh6AJB1fi7RSSF5Hi63oX37/J12k+DMY7YBUJD07QiIFaYrYPRRgvJWQyCdddEDbAnLzKA7t/
qOPCX0eyNlOE9TmFXhJGI8mTRnfmTHS/JqdtGPcidoZagb35Ja7dtk64ZDGKDy1iegUP1dRIs1nO
MXV3lmiyn6GnqPNoktehoZ1MT3ni8jU3TRTyzvWBQD+S19qym0QnwCQoVRH7bRT4s9bDFa6k0nXA
ad23cERQuLaEkZ5/QWMBpn6ENL46Yj0JsbnL3x9gq0ZFfCJvoagS3cjiU7ETjwO7hV4HQvS3jMKV
d7ytQW/YGNHob4gc1lgsxnJtJcm7DbKpK5HHwvhWfr2BJaHyXW7yb0uDQh7jEconyWSv7Cw3dIMY
ek/oHzCIZ8wnNKaXkQbWndknL9GmKp6ANC120wsiMHzafEZZ8kdKa04r+v2CwQHzQ/kLSkUWfy8e
vYKJuHfTUzqIEiq1rCtSmPWejVrX6e9KXndViCTi22ZOPYlCRQ4QF/CvQ82erBsM8BRKdoSGiatg
f67xchRqnL5YRkRlSQuyCjf78yDsqYJj2hMNRa0vzsWCBXlawo3sKWql59YtJEvBlyTfw48wyOCn
L+V11TjhswWLwAjZqFurmRGR7YCeiogSw7Hx4P19gmh/JWY3rFyX0qZg0gz1ErayUPSv5lCEHQAp
QijqILUzy7bsC46gS3j4NRwH34rC2VUAOOaMA0vmYg0lYIMyI1BrmtWP94dozv0lJWO1F1KdHmLy
8ULO+Fzcw9Y4xkdjRlj6HG/3vY61dF0YzX1j+8PGu1fM5c8W/2GV30bRAEh/jrsrTdZ9Mfa3VXqp
4XBpLPjcHlHh0JILuQtkL9IQ7WhkgN2wKXbT2tTjN+qXOUsdYR2NaGhpscPutT4S0dsP2MQfBM3S
mC3tieR9xHHJajuDU4XB40TLqTwrvc1NUmq9K4H2hA12ET7YeNJN6i2JcktxAtxub9OFcFT9zx8Q
J0mKKNK1EHXzVTQmo4WoD0HLjEBsMPOhRn2P7cRKHrgNfmoHlXX3oaMCsrCeBBmDSNd+ZNG5rvFY
RPTOeuVzpt6jh11tkuec1U6wQglv5c4mAz9xAHrzqI+gleam8/fm8vYbJxSw50tcSjjJ47+jfrRF
OSUjBeAGaYLVtFxbgxKel0uLXHPOoLx3h3twOOPDyoX0j+VLxlf0DC1u3EmnB4MCYwlSNAeVtfLi
9y67/o1eCnT7X/j4UX81cLasy6YwoNiS/eABIYTuuHlirzcFztMBXXFl94Ao/x1/Eoy1eCNelcKk
0WXc/ttp+A8DGlrjrpCOy0qTVr05hcrhRjcYPBuurwLu8X3/ZbgtKUo4P4XqYHpcVHK9z4x4lO9q
EG5zf4CjXe/oIWgP+ljaBDXvJ3Ke+DXDWtUJgA+S8tY9AFCj6c1z2Pgc6MD2sFlpC2pORZaSLXrB
Ne0lUlgdRmvY75bqwKui/fUrhD88RNUlBdYLmdD0fBl4Wnjn7dJX2vjB5hYjS8SIYbhJiqdJplnF
AF0tcU2gWMXT0qR94ISnCw3w0951g5R2F+v1be26tJRIxVhJ+LkIegU08GGBX5RZThx29qJpj1LB
hkNVHAPmgj7EgwPSmDosdgNe/eTOCxkVYlY3CcCmP7Do4NgBm7uOAol5nbvPMuYB8MlPsXl0elPm
ESSWDBV+GP0tlHYRPXR+8Yp+lSBxdhkQueKroIl1wapbyKNjtyqXwRXfm1774Smwd7+jbjNgTGL4
fEng8jTdpujSDzhKdpyFhiR4yHWGwSrufKkBrKQbmZJfSqWgAoEFopUwQtg77SJyNLIembiAzmc1
BNgZp0AMEG5OBTYrrZpRcyABfyOMCfW/08MzT/vXC/sg9TrHohDlFDxDHQmZMnzDf7bpqwpLA/KK
tloHWKtc4PHdzY0osotm6s56iuV11SlnyrfQ9ufRS+vacdhpuaMZReRvjTtTKngZW1iP4OBoTyA1
Z5veiw6gPz+21HpKj/zYdd9TsG2OQ/SJgHiuZ9hi5oMeRFQ7HV64cO4fRoB3JngCVC2bUBUwZGpK
i6+c5fxa70OPFSfM0Nol6almc2ve91yHltkMKsL/b81U+fkttoDWC8kPDyfSUdyRt4ggGn4IPch0
vs4sKxb41bOhdDGSebJU3L54gyB5iegiwRCsy8KFe7CXp5f1RNMZXIOonJ3XDN4C4pLJqrTOMAo9
SvkWhbqxGYxXwTCxq6IP1W72gRb9wxaYZDo1k3RbpV3fivWIBTJCMMWpgrwb3HgRD3Y18CuwSaf3
DqwYNrP7S7P5AIVjIVFEWAffPeoZiSvizoY1S2ygbUIF32mR3Q0sIOyqM2+2WwRX6IBw5gUA4/u1
+vo8sOpe8B5LsL+IeUAXM7BOYRHw4VKiSh0LesKMQm7XZFeBLbTwryR+czsg5hl/WyhrcZBT3Sly
xkRFnmoZMHmo7tlbSIrGJjrzPbFqTgzqtLmn1t6yulhlm8dJxaBg1oIJpE+D4WD/kbXSKNcPBeLI
/2/CJuqkzE5wqC403oxV0ifNdpTCDkOgs8umEMt5uFo/DF4jNFLmw66fZVqXtJh1QofBu0Ksq9cv
FoO7Wbi/QqawL6Jh9436srgnG5Z9kWlF1zPbQQbBGTCkog80uZlpudTCx4v5W7qtfZETIcaATLYn
4yPmHMTPW1jk2a3pw1A2pBe7XKuJ3h2Ju2LeVxVffHd3z/U57hTFltozzzXhKaIgpatd8fhvuIqG
b1X1P3qg/2j3kJs1f+R0AOt/XU9HeevlK4+dCv2uvX6q5Ub6153YYS17rSb/BL3WaXxxZSQcUduw
hT9q7tE6h1cNQzCwk9p8J9dRhJiwMIH3OYliepCTgcgYfl/FZOyiPDZXYggUP9NMqXFie3XJnH0T
Z3IeeJKHdpdWRSU23qGqSMC3B53asyfOp9FAIxDhDsA7rmOfH1/r6D6l05SJRv01E5bXqdymxy0b
QaZ9Qit8FxQ+AS0Lyl4AghmIaXXRqUiK340u8bMKw33uZ1OiqVKo9lpOimv84L7KgGFalsdEmccr
OqcI2pkEwD869Vg2AKJMfBzJCIQI2Hq+nZAYnYwuap8ar+i71wpbsFw7hv7nzwd7+pAkNlsujmTy
OOzrFQZ/0kTBySBllqo4Yx537RLf7L+DDDwgE71cp5XtFUmV/rdH+eNfR65+JTj9+JlKVck35Fb7
5qwQytFzb69WeZOM1I/CMp7dtBAIEl53PWjwutWC9Y1n7wqpt+be+y+8VgOExEvLUI8y0foF8Yke
mYizP3Niw03JQJDcKiHtdP2ssElGwcsb9vHyeuSLiwvLb8sXzsyFWEI5Qtp4a6sr+JEvr6e/k3A6
5ATt0V5YyfIcMJvelNblEGR7Fe/GrOeD5a6YPHroLDowxjfRBQn3runN8Ma5UIZQdbpqTR4KO5LN
pL0YOK2IZjRejxTXsORYmcaPuNATcfb0PNvuTO3zh6lnVEG/fyLfdH0cNSkxdk3qclYQmoa5XLHN
Y1tLvIrFXxufV+8hUuo50uY0kkE7ZgxkGikHMTJ2avBLel2GQE1iE7pr2enMp70J1Ei2SSkGBlkn
c6+d9RBO2a4BKgucFFdUAZJdLoSWHiGw6NCMmLLOh74AWroAwqeWc39WfGRNgBj1wDp6cgqjAyGJ
aYOvLet0sH+dMQt1D3yDVG4ZYDdJ2EgIkQrExYjAyNIzp2CbOuYTi0GpUlIZan6S0LA/YJWDgeOG
vlHe/UEZw1innlr37ludqaRnJtjlcAQNMgh5XMgbtSpP9ZtTajSqBVrvGusdWoIlZWopyrNX0uEa
pxXXpB+IRVAvPY3atPYRSUoRbPuCYWyy3uf1P0qcS7H5mGGin/aZ7nTJ3keYmUtylmwQAiDAO1Eb
XJ0O3P4wEO2wGAa3VvadV8HxLfRANogAiJkaoF+6f3wROQE9dbFvOSyzFEJxWLaxT6hxC64VygY2
YzoXOTl3s7iFHN1SQeYyfua/aXz/fSTVkfl/HTT/I6tZIHS0gb5o5a4QU+ljY6ADVIMpqV47xxuz
GH26ZSz3upOERsUTF3N33zXoB9lPqdPnOMN5KV1icDyoqQKcexBtSR8Hoq1/VOgrYhy5I+DA1eRH
Q4PDtWaZW5Cdvx/ZiEUO5STQqZBtGMGRelciJVV4BJsl3IpEQ+hgiEdsiuTOV6BJFUqBXFPfQLPv
/aPLBnACjXom0SfSn8Bmj6eHtnxXdgMkUd2fAdRUIb3rxEEtWBvlLRvCexDw5G1tsdCycUW8VhME
mI7SZKsyDxJF4Q12a76VJs8CSrGJOCBICD6DTz0BPhbPY6BcWMf70Cnh1eO07aCHGBjGPZ4RZwdV
BsLMOjb7OM4dSQPMlj1Is/C+Z8xYbRpG9fKpBy6JwBHAchLwEEgHXzJE6Fg1nHsenY2RUglwEvAk
i0uPDc4KjmGFFZUfl0rjeQiag6xClgLbENZHi6kgpCjpucVe5FAcQzmCA0zpZp7zNq0OGv0G/EI/
f1ktGRdn3fT9CKSqKJyTZvNqWVIr9IHKlfvwaAyTgwsHZgp/icVN1POzJ0rUA/ER01SJCIE//sF6
+4AIkKVxOLmFVdo8Xuf4DEReI12jYOkcPDbCqCoeCHYVWCdcULkpZRVzztAEVT39pnwQtBFfoKs6
AVmjomQHa13E1vQjwI+P2qrwluOwzWbwTSHxMdQwDcvqEWB9p6dKRepHo79tf1O2BZxSpNazvRUu
fk+nbDGsKIqPB2tSw69haFYo9+JYh0DGnTY37MYrWNGTJfZmLlvdoV07cipkUktroCg2anNVluKu
HO4AmPQ8W8lgGLPm9wFYyxu2J44ESjFvwLLzDCPhFWVgBsAr2EVnu6dcURIlfDq3n02etULy1we4
NUjKX2HR5rLu/lVLQHNBzovhv9HSd5I7+s3owosJ7jGkdelUBq9t/2amPc1/RDCUjTcR05B+gCUN
1uaHM/hK8Zj9dY7DzzWsdxae3KpbNmfderqgEW7tu0/7C9RUFjEfdzzUZUW0gH7qNFR7lELip/Hv
jxlzKvVgSHFASDwEhM17KIlYRS2IpW8IAFujhhNvZADZylLbfGrkiPPwWKdS9Jia7JPpPb2PQVRW
FGb+RHeKV9Jcn3kwGT6hoNKqVxrGD7+Lz2BppEhDrmkHUbPJxYbmJmMhXHYe/jCa2/F+qGhjZJjM
3nzYJmp430ELv3pdawtDIT0X1u5PpPHNs9z2VQ9KZqGbf4sgpglKex0zqb/nfaYWfRFt/IWbIwUi
LB0eBjq5bR6RHVbkj/ElB8Ri1N84GjvwudAq8dG3p2vS01OwfDxgPioNsC6c7N42RtymlPqt+LEN
9V1zS1HkwAZoSvxjc1KvWXJcThbGmAzYgTg63LMiICoCgEG2AhcMw0z5fjkNyY3Skd3FRB4jjvUz
zUC3NVKYNOMiepcnQe11/sObTYd4sDCls8/mLto5Aq8JDAkeWDYEuwLwK6N66Cylfr+8X8f2y7wt
juyQHrJchuZGgpukWegJ2c3xOS7tdDcVY+FOhFZKGfh6PQjo6dMl0ssRb31kMRakco6RzDWiadfa
+CQs1TcQ5PPyL41mBVwIBs+ew8TZDko/jFC+wZWwUmVBR4eJ/OEbnQUWfdce1TGq7H7S5Cp0RKlP
BVokaJgCFF8Y1OW2+KnDvkS97fwA0lDxz8Mf3ntz2sFS/xoZmfM+Flp4LqHsLK2p0MhWTNWuqb0F
Vwnn1+5lZ/gEhGgcx46vzYSb5yVMR2BUQb1cNMcZ6O70WtTyjsQSxi+s6bxJ49MIATVQRvGUx7F5
7pBCbbKrDwMlzgjT4NGQjTs2bBsFQyNeo3AZ3CvnQMqJq378sZxkhtdVEpmccPT3RCIpBOUaJS2I
62SXc6/EcY5ljkY7ii3t5iaVsIiuW/H5s4w14I9Qxs1JAEHKxYpL+fbzFHVVwM+XH2BVUJj2z1Er
AeJNM+5FKxY4r0w8XRfB7jwBa1/55nnNw6CfW6IaH0iG599LKRIZOpNPX7D+pAs5j1Iwc0HE6K7k
sz3Qv82XgfzC1uoXspSMWjKDml1w2LA3Qt61G6XC6kyikrURR4b+VoYBH8e4RiZDJGcze68cfPvT
qNBAIjSbCXifbeNMeYhvz3oFb0AwB5IWnQbTWxqebjPY//7nG02IvrN6DiDRQE0g777rpRbPe77g
FfWTTxO3d3tY2YXQdEvAEmVCaCd1yod3T3UJU6IJUkFccTenVSkF+65T6L3nBVI5c0f1DBjt3fsw
VuZYMKRKMINKr7+WM0VQjr33xxjvcN9p6zEKj2VQYJGdck0O2ADphTL16KTbFG7MrsPiSySSCoot
wTIuxy6ET+14NMjPYotzjPv4lQYEwq/yoUOijSGxjWq6q9yo3sb+s6D9zl1Kik3f7W7VMIo756PU
uMdhBRqzhdjPAi3gU28o2u4BLUlALeLv/q179kZ3mcoE4BrMC5SBCba23BzlPUQlbdWcWsbERkE6
2jC/273K7uCTqvNijZR43cTMHJk1S+jomJzQkDKznVyy3sc5y4BFZ98Tke0pzIIXbtBZXtYUA04I
P54TSgKrdq8LWQnPVuVoqR9KBbtLeuT/PXPV8O+pbH/MPmgPvloit1jrW66Gz0VPvbCsVJrjV5lM
IiiFTOAUmKTdT8qdxBBCZDX2Otr+Q359L7zXuMoUiMh9a96qEJsc46aZZb8EEzxLtx+8sT4REX/e
hUHqo97xiZjnk/OBC8TiFhgHihI8L03GR/MoYx/N3/Q652w3gTds8kAkaYEZxlJadQWVI9wOEaeD
joWd2aetu7NVNq/I4lbAjaMksVtbQbBVBjnYWbNoo3AkOyjM+hc1T/GFCiq9Rfq05aJ6ZNkmn4Cu
wYApcorCRlYZwkydsv2EzFICvI/AwpeoaHg5dWopODdr8Xh+kyKC2Gi+AM/6QOV8/zDhDJ5brxVd
tMkVFYCPIoy+IrLvGe3r088zAc0TFBRie5Gs+Cg53BAKFCE3DhphdJZAfkEMEgcD4+RTVCJcMP16
4chr3HSGgdgQiTd0pluquDp6hgued97aM8e+co6l1jtejuLq9k9FwxZ5eYLUNAY3Ji00+eEqTT5B
aR9cnumJJnDXWKIwLGef/uW+HRd/M7tTpiYGibygPenCcw3VoSa7NU8icANqStpIQor5/hm8HuYn
3L0Hw0rvLj8F7bxJn7cmt6csQB7xBkgrrOVqjcwpJNlQ+GmcXhrdkiuI+PTiO7VeBuTcvvL0/M5D
oQ/6vQGaQC4lpmb34u9dfYbuEsTO+EZgZapyEDztI+GIWgKydeDGAoY0cpBMUt7zakLGunp4Axz4
9oztmymWDt0XWieER1X9bFVk0wly7AD/ElHWnMWg57vyhUPVES94xyRo3HDzYNvzpXZtytSngk9b
8MWIULkAywJbalVSdoFosCHeJavdDw3SInSfgtwTKi/4nxKo+2Ov9JyAs3e/Z9QSsANIAh4uWfPD
EOBnBJeEqeWYCR2d6s7hWVDzNJNu2/D3tHbvpCDW9BHQ868Q4bo292ehNWaSIG5qiAtE/1Zeh3wh
aTxRq+e0tujfK5znNsi04Gk742OHrjd/EDb+227AdW/4J+5P2H4tB6rEBy3eo5Tz2Qmq6gsM1pLd
mqTx2UY91Rp2DedIt7Ef2usJSLKYdUc9ozwMwE7xWubjBpIH4EaBz9wB5IJgHcV8cVL87uAthdUs
7ahQqL/ruYdhDGF286RWRrpc1GgpPWRoeZKCeLW7odcwADlD5/BElW7Vx/Lxr5XBY/1QD6uwMogk
Os6XAyRSo4NF1cGTENlvom1VxfDR39YJe+r5JXeNh/880sbtl+ROy2kQMEAI/5dYCJOkYgKhBDvt
YPF16+QwPJE2qyN2Cc2uR5wO8FIPXHNaVFcWNJf0WRFr+imgKDGzZ2iZ+kyINU5uIGFyo4+228tb
WVDwic58TKCOJ3Ld/OfTgM6g9cfvmZXy02vDuTp4mcmt56JbI3JJOjg4g0iHA74z9kSJ3M0gKjHr
9vMfQArD8yd0XW4/u7h1Z/STbMoKarJoLjsnv/YVDVgHhygKUx9D4xBG7+jtwwlfdZqBwBf9riIs
+/ycdKyCDEl2DlJQKyFCW++wNijOfUbmv+jB57skbMJty+tAK1/ThrTLpoXcX/JUnMjMkP/FcZDV
3KDER4u1Q3FXMq28c21AXK/q8RKtCpeMx1uHYI1K+BFABOUhP5nKzecEqtEFdLQU3G30mP44K59b
o79HLB4zPqxq8JhpKpzcuWFOrcgqfLdocZOcq0oXVFOTbrP1wttch5V9eTtb4cyqCueD4reCp2fA
/zH0ryBOR3BFe/Lph4FfmIS6i5VPQECKCvkTsurLWYxlC9RxQcyOHssRqUvNrdVI8VKZhuA9xXNO
MZEk/bmpqJbF7zTIFfo/uvYkZJ2XJnE9S39C+vRr2s8ZEkmZaIT+CMcR/LUQT/2begp0pQkXtASO
pL/2iTM3bPW7s2I/MU9QJRjcXxuedX9Ub76tfTHwFi303mFszgvIiNq1KwZHmveRwR4cI6+XpO4d
PerK8T75kifuPHIKag03mYuWYNNrY7aj82ycp6NVreX/H714dERXlGeb/VFZg8JErdOVAZ5to5Yt
M1EYRsW6JxBGIebjAG9DNMHTRyVGA9PqKNl5TyswTR1Rw1ls0tfkCOjFWS5o4ZhGsRjMuTYDQMTa
GVGs7bOg/YcNkXz+I3o0dzv09zewuyiXOEHLEDL3899FaEqNkfZpmn/HWW0jYA0pDUcYW9tj+lMi
8YfFYparU4/sc4Wxv8p7ffjBJ9SPLG8H47ojGpRCdK14FBQgdbJe4BSMLzDeKT6HbS6nfcWP1asB
y/tiPx1gcgtk3FEHC5NaQrt9U5R946tEGeR6Qfkr4sssVdPJ/LoEm8482Jck6oyallDp0vb9ICJX
Sm5lVr843iMd4DGqVmjNIzaauXde7RTBzkP1ASu1Q2EFQhtQM5jXxLKSUxC0dipIuBIuVDUIkFMV
G1DK8oZdDU8zr858nAhQ3MscmrPQBgJb1TCmJZx0AkEl0x78gvbkv1eBlaupBbFhLjnxvFpCtyZQ
P8/H+tN1X6LbYTLc/ACcRMwrAdIJi6ebiCYud1g9BjDANqVrE3MwMcHlKfnAl0r4LmGPWiux4eZC
KSjWiWUYGmrAsMXFDuL/t7LUDwlmQuU3fKGPU5WkVLnOqi6qteloJhOjCR9cEyMTOzu/MFssBKpK
HQa2+5iZUzRFX+RzTDH2yZg/gHOxJ0RXFy3OI/CVO0w6rZAyYKl3anIZH80+bJiXub/a7bXX1AEV
qht/f11fd/L+Wf2x2zl4NIFkBXnOsoM2qnLrJReMGRjKNtK2QHBosoNSLHvY58iZi3mcyUmQmMv6
DupPTF8+0mIXEypKiDkCVjrssrAXt+xR6eaU8CPCpu15wLhPVHJFUa+Q24JGfYXjvO93iUi8cDFc
DdOMX3z2dA0T+Opl3LLEDXVnitmxns2oUr6lbN+U85GaiPaSxmc2umly+AVc5MD5N/uInNkYbFId
ZKVcH4+SxkxhjCvYwdK6mkVUpQRzqA4RpT5FNRwKgDkNoVh5YH7mAEaNpJava4khULj3uu+rfafe
uy+uan8QBeOMgDPKV934gZRA81GUF7nQGtcEKrHdmFrKaUsBGzy9xst29TBuQmfWATZgzOh87xTS
KU/ATSs4s5dYqUkoq4gRPAr0fqTzhKSamV1eLV58+TepsriiN6NHRPRoPDFdoZQoxuqLFxI1BZF1
RaMyePraBs5IMJa7gVnl/WovZH2a3EWFveOm50mJOKbe5tOduGNO3cpDoDPHlU3YjADi4ita/qyV
KpPg9W2HSOZ4BBRybwG7xiv3t83s1mm3yrmLFyWJssV9ijIxdElt+m6drvpoFmRkEcTP+MNOF38w
ywHBUbnDvO+RbarWVv+YN0zEYs481Mq2Zb5xzRVd4EBd6cz/SWzmKfwlRX2b//lmEgum01rQFH4+
gR6d59oSlaZEl+kAc4Yn0JIN6IIbixZwIQrosMEbCNxnulYyt7PFrcEvuIGv2QBOHsDdGpFs1977
/65y0uzuSVpxOT0RdOyuIow+gxkFOvZvumXBJHeNhpwaXpm44WtecpJNiRAyWQbo10RVN87KNkb3
wuWcXwCytjX0z5PBfUlsXIkP7RAGgbeFHsnIg2b1ZgmJK8KKRZU7NqRFAzWUBsEe+wAnzYY1brRU
Y0FWWkDQCrzryQaNTTkofLDzrHBqSclcQPb1Mv3JbzLAKeMCGJ/DPhbwY6eQPt9OW5TZI/D8WnKh
FXWL0rerwGyQJlhUsU37PT5nnzYRewi52PtX+2AtCn/raog6aulMUncGOzK+wQVxXTEacOcHaRui
6Gj6lxpE9ymwC49DtkXbjcpd2wIno32ZZKAEZU2T66Yiz8zp9fZMdrRNTToYFFeoBl4Oxb7/sbW/
0BoL6q3YQgfThG+z8gIvw9ylXYQQHYC12YHkaBxkGgrXYGV5v1KNey0Ja7Hc8HSn3w/r2nSgfpGW
CO4eWxjWP+ZXWjNzI+3yBnnMRLUR+rXJ9q2hf0+K/Jv5egMGJJNjZlVvQzgsUCxgb4RFdw/TmMNO
7dhcskRvGECW9ad45psndzdKzwtLERX1opq/Qx7UfOrq9sipkDAHFifPGY4k0WaGbkWpb5GRBOsy
KIIZuUwNa0ryfbe8dYvyS6m6G8ne34KITXhmVZcQ3GfNpDNwvFVqcIYh6ztNGcXucGcH59KGq+3E
Qn/nfu64unHaikmQissCwJ4CYUCGQnNpl/uRRyJX6utG3X1ogExqhghPjsYp7NrnvCt6s7GvfOwk
8J3sRWZtAnRg1v/rC8thd39BwLYpbibTxeYS3nEd0Ewph1JCUP30CESPpIQ3yKlPXFEvfVlsKFe4
NPEULRzncfcKC8BRitkBPGRguAX1yaXd0SSprqXzm4UBnNc9A9ZwnxBfwjvKgETPXk0SPXbTX34r
lt8AmbDef8zUbw1pIVsO4OmdiakAJMlaSt7HKhl+i6p7XIRSWI3QYng4UXL4zWmky/DdRhT1xaZb
ZboWF09sGEkHQ9IW9fc+Tv98jV8CtvZn30CJEld6uQlxNpxqnXy1RCO54QbXkwfx5mpx5yWYWpOE
cQu0eUE1HWTrZ78yubCGP08IdGtGJyFt+W8kdzsWJSW+yPHH7sLiO9AGyrPaMcz0X/0a3dPHS9cn
jfQbVBNhIKrTrxrTcBZzWI290yJmk0Kv4Skg1hwU2noNnYsqCaPjUaHF8TyDyBEL4UqX4qjUQFJC
3dYQggFE/DKzzbrAEDzEamPRopbsSgpMlLSIvXFztxlsIHdiEG87j9ueAyTI2AfyEeWaNdfMbcP+
LnjU50qXzzdqqhgAJLPGVOn2c/BXjc/QPsF7bNXV1+T66AYynr524rCoqX+wkLzx1T6ha+gZfdfU
1LRQpk5BwARBLiO/i39yL3avOxr5GW8hPA48wSGc/z/KtxtK9A7axtkZbA21PAKTTIFt7uWyY30z
pvK6yK16X+Z5fja4te4K8yhJHO4VcRL8Sf9m53QgRD/IUmO5qmgdjL+xaRMGC5AReJBz4vZtPq1w
FtyLJ9nxp0O4VYljZQbbU53WOPZ9T8VLY6298BzxJvYuH9VjeXjq8+1Vh2933laz2kEOZzG6b/3Z
We1oxqN/FeqHo9Lwu/eKgxnOcYXg5KNMao3qsbnbV/dzwq4xDXZ9lrhD5Rp67PKROc1wQgO+zs7R
VyPATQlLXBWwQ4b1eHjKuu6ysfR3fnPv29Yj60KOGe/e1XfA1eqEoZJkrsHNeKPnJb+r5ibG6yW0
YPc36wdUpYihkcw+92v9Xhqzii7jpsc3RE9pC1jMccN/HNaudddpHQ35KC8VWalMQzUl7EntRdOk
604W2Gifu0qqJaiE07VfDAuUNNe2UjePz0eqymicic5xnwwKNxWWTfPm03cOIBIVLuKKFiEHet/L
ps53qHkF8R7dbNh4Fc0xldaIWl6NK08hzKEn5rqrQ9BPCUYClUaSZJiclQrZwVBfp3K/yaJ0YfPz
dS+jJhxjjTn7MDolhb3REeFShObXSDunrsmpJPUUVCW/pg7ISw3d5IGM8RvTQYTHpyHFgg1GcglX
6Kj2KtsqiHAwYZYfIsTC4ZI8djzForKM/9jRBWYCf7MChIETc+p2Pd2P9BxmQkJ7bJS6ItkznczP
UUUXVLAwFt0gYENSYBfc3Ndxl+GfO15TVpKAgFAgFqANLfolQUbw2ccbfuvM6geGZXK7RgiM9hrc
7wItj6yNvzyoTYyoTpCRKUtNZvigGBNV9O7Jioz/7Ny8WSrvQ9itAepfugmKlYS89Cc5iIQBsoiv
Nq3Vkt2Mde+D/vZdeBPQ3UUYsv19DpeUyLqQ7ex3C0irrej07iablbkJTY+cVJvc2o+0prAd2muP
7NrtkLD9Prx44aHtPocfIuAKjEQ/VTS5MjEhC6yHaCwfeF0RFe1YcHwlu4eWEWJfhNOmb07RQZPA
Sp+iC02RkJ420x57rlhslhe8Yk6mz2YNjGOmFQoTo5Hhyzp4ut1Q39Evpmfasz3cZVwtUlIcEN4s
ZOhRVGuj3VNXIW5hiD2hKsbuOb42uG3+S5Qa+dM5KGiY2+9Cj9gfPvuMdwToQEl9ACDwWVuGOrQz
HuXMKGZHmpl3qupk/i9ynkUO8lYWGA9RLLxRETOkI+uEb358W6bsFaPHXUKUpQ0AWLxm2j0urar6
f/JvtgWj2J8JC+dSrXYkqBWLsbgNqhnE8uNqAfKH+wt2dbVWC8XQAEOTiVKbrM1UeYCCy/+8QaVU
/fp3Sq+Vm5RKm78iBwQwUZyMLShu8s5xQT+OO0td5E5OcsYl0yWObOYWPKzclXRNLHa2XNxBugEV
w8+QvkyGr3LyAIgp11EipjPEseAtzd87O3ITHGThWb0IkplF5EKOrMDflP9veqo3QaXYfQ5iwVKx
h8E3VjduI54dzEET/HD/SIiyMJ6zFQ3Xc0guCkGrIhKbpUpkSNjco9E6VN/UBcheyK6S1PqQPAjl
xPHfi2CqyDwbNE4UrKfbblEOCOJeDIDaj2Guv0KjePsnnbR94pzLKkV+c8ipvaPkHAJ1y7gVXCmY
2ZkWspjWUKW5/wSrLqZJ3B4t0bkMtWwXOlDdi9sprHgrFZooplRgZytF4YQW4KdSbLPfT3a6WoN1
CuV2QPufM3JCH2APNI9Q+GVsuPTIiOVbTbHRitLETlZrmyhWWdVeRgEostz0+TCU+erwGekAlqTO
IdCeo8XijtbS7WKQzQsn7bSQ0FBTbb+jULJAq8nB/g2nbCsgce/0a52WeErBYGcQpVYbrLR+XHoP
gYO/ftlN6S4hxeFC4HpwdR3PNbR3E+eVof6vMCPX4a+YGSICH3aCOAuhn3syRkYsMlgtugRR5ejo
4l9aHvBuQR2qEIa7iSdr8duo48oQbD1AFoo8OduZ/A4/T6axYzkzxBUZ/Z936vMnqdtMRhcTJiE6
A7jxfA9Qpgx0KJ4rimDFAExT3CG/ztoyHt+B1/fmCJaWKFINkAM5nfmP1AIfLuQdIroZTpuk57zy
oYC0D1x2qJH4y0xa/ka8BTGlVHxI/G92e52gd3i2o7XYvluGblgYsK7qtSZ+o7wPIS+fuy9IJskh
sXLlOw6Uv5zgEzwZGWNwmqx0SPVpBJtUNjKXFaX1mSqsvyh6BKBwOFFG7/WJVjDSSHIVrvSRIkk3
FuJG0CiqKcDT5h7gwGIAZP3az0vS9yqqU1o4trnckAUrJK3np9gjspmW+RMiZYSkO59WCGcKfOLl
QV20+3+TNc+WdRh2XlNZ+84vHM4JaGRZm4/KxnwZ6hBDfAYtnvCOFXRK3feF5b73n3nUmP6PaHgs
HGpZVJmFdTCJl9fNfJkUd66gx6kA3HUoetiC7jwBuTnx5WMRqq3NjfGsHyY+Hia6R5jw8obwlItp
bKVkxWn6MMDYKGdkmpVgRA1BACJsclugLkmF1mt3edgBQFUnz9OHPHhJ2QT4e5vo+Ck8jlz+xBjX
qMT3obV/3mCRVqP2jrpT3b80wG7f8WzbwFYavl4dCHLmvm/jtnhpoQMLa3Cf5yckuYkgONf9IwWT
4B7w5uGoUUVoUGCj9Q+9Ma2qzAo0mAE4s5W7+idXmp9yQ3dw0kxQOeCTMzITeATCvxoJ7lywqKDY
kM8Ru5yPxrxU/aqr4CEdToL6hPd4rjGW6iN2VoHzHYwEYxcvfVUXJ6Bi+M3avwMxe9NDoBO3PDz/
rKxHfG8JIWMu0UxumYqpbrWITYd3mR3wmghtixHvw2iF0qLxDMF7vjwRAnmjHcsfjvuVgwMFoLeL
TJcsSVt3rGOEsktkn8Za72IXwPtWCG6mVBDemdJAZmqc/iCKImDzq8hvRQ3C/mUE+kOWYtjIp7Ca
e5AhrRUg++oqH1fBwG4Gtp8Ntzpjpt9Guz5tZjH+BHUfhW/46gW3Jw99vyxH8PGh+VQa+f/kZJ0L
Z0mKMx7F2qtegOXZonF4sRvSwQLC8zq22ep/0Robvm4H2THDaI4v4mpjTqvFN/Z1plD9tZVXMiOW
VR8oP/ldmyePQxdgnBmPnsXFeDhSqI6tZS7oMAkF1BfgtVyz1009d+0ZwZ3axDDZ8Kp5vYS4DNtq
+WilXHKdGzgCFmSfk8MF/THAGFneABfKjZfvhqTE9gsIGj0ErO4l8CtBdWCtrdVJ4m+cAnDZC17F
ScqzfXLgcKNvBWZq5zveERNytXA6DXNVBy802l105oNbzno4lo5/ka8IUnk7DwOsCicuO2lDNzd+
ib/lQBBaMvtgeQ78q0B7q1LU1EPMfCWjEnHq89HYAT//9Y/H7YkU2VdJDMVxG7oQLlslrAzyYB0N
jGMn+rCGBKZndcFnzLWWZeDbUwCTHr9r/94fFRhobW8OUOJIKvYd7W9InT7AUYudzyBW1+mvCjQx
QhR0sfhkSg5JJ+G0oe29U84YCkY7MskkRMjXlpNn+gUSEByr0sVJS5A45AiuezGSeJAhNG7MDknC
A28udra08uG+kAxyi8ol9gC+du8l0+KJanZtfJWlrkN9w+b+2/GJ6m9lZTTRie6x4OGqPu5zV45a
ZSghR75i7r1bCFyu+MHDA55V6oP8XZFPp/4Kk1ZCisQDdz8RgLv3ag1vkTRTnDeAHjTKMoXjRMPI
o+lsa+XISQSLC9Jgad4fQUJcuICGtBMEPpP69nYZpcxb+d6VS/bXv9JLwnkSP/ZuGvCD+W+Ixt49
lO5r3ctm/HllXwzjtFX0D3jXtKDLRi+aY1FUhQRL0Lvy8cg4g+2FDlSPY8n8TUhJaR2nTTheRnIU
th2xoLx5pwKkYsUOXpR7wR2NrnnVCeyd4FPlzZz21esjcZQtD2hGquKs4DJMeHXN1He4i4L5zZ/J
MHTV7D//zmfiOaxJi98f9h0M0B+PNIrAeUBZ51fMON6oNKrSeyTozxVcxSU35lovzKcF/LYiCt33
irTAI86TKgg9gH9upoi5ZcGS8Q4ZHV4X57+SuGt8i8HLuiBSW3qASt02sQa7I+6mhANFrOMdi8+F
/R3G
`pragma protect end_protected
