// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
komXqsru8Vs0XTZlSNa2dO5Dl4D5EslzsN+jgjnKPL8ogp1KvsMZdhUPHz1vRHFy
qiMDnPD25Ankz8hWeqsrks6Df5nBiiWH1XFelCSFp0aj/e4KJraYP1DYhQEkUpUH
uG2D5mz0SswSEanPNMB7VdVQryivWfy+w/Ry5kuTJcM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9472)
syrJt/bNvRiBFzQrkgVZ3aThcYRP/JOZ9ffP7AcuSkuvRjkN9jhWNWaSOPxIgxyn
xVqA9WeH//ImyQyXcV1rr3uxpoOdiK3GzMSbQWuoGcOJ447BbN8sAWFrVsflsl/f
GWLbHzOPLBuOH678asv9bRyyCCQRvQTZNEZxL64HpeXUkw8SRiBVhUyi9/EyqNEl
OF8GzDuscQ03EiWbWUzMkLslVMuC2qAP6wsiXvwq70Jt4P1bkA3rMzLv2oS3Vfmn
y/PKg+ZW1NjmLGOXHmFNpbfPi267a0iC0hfmYZIYjPvNfhx6+jGs3TDPhffbrFPg
nscedGl7Wwyc+t+bCW5ADkHFM1TNZfAAQADn/E1e0lfUcwFp1VzXXJrCjLCaqmZl
6wPxZPa1Z3etaxyE/XeAvDzAIxRfEGzRxUdjl5vdCJlY4STEOSb3T14/sPEkVnaI
QLoy2edYWJwLnk/K2mQnpmh3Nrb8G1B98BYDcY9cikj+0RUYBOxUr8IEMkiari42
cJLRRnsLcFRJjMvZ4Cc6KB6cm0jYCKHjJTw/xguNOCmSuxKIz4kGNB6jgDb24XTF
TifJ/u65JU6kd+Sr522wxT5PX07Jcq+BpCWSqH7JUQu/fl1rQ2+Rm5YzlKyKfA6K
UhBWYvKI8e8VTfXb9knN76pdpzp4byLJYh+Iuq2y6hET+jZ9qvfpaEC3p3rY35lH
X+JJNNDLPX4/9mKkmR1/6P0MGpaBE0xS0nB/3wL1V3wLXgfnFVWdT7q9hFHFUpz4
PmOjotOfDmiR21VwiTd7IgvaHhHYu9fB9X9goM7cUoCPK5InoAsysQn9kkXZEunj
jAOWEPTLRe/uh9fr9Fy11XX/9udasvZ18gvl0BihQt8MC4zEiq2p+DY1P+h62r72
ZFXuAx3/FM6dVHkTeoUeV2kal7I2iFWk5DqRTI8jatmx4ee9Jjg958M4uAFpe7i6
sOwkORUMV1w8E4qUUYMENlgxgTUtxZm6NL4tGwXcmsbAvC0Sp06q3SK0lzTLtSJf
oDjmJV9QdhymbbzYjXOMYK18k07IzHR6M3ho4l5DwQ2412nEmrRDvOoC1qhV5lOb
ahY+4lZIEisM/lDe77Yt8tY/pctu2C+KY2YHQcd3OwhoV2ERnmHf2214fSC1QSlY
AYCzZzBhVgf9zBVQrpcSmFOhQtFPyCR65G9rGzHiLqkBdZSIzWJ9hmZr5/+Sr8Vd
39OoLVVY/Nc+V6PVsdhVaJUWTnTTif2XZr2jxo+SBwzyypjBSpfKw8PdP93L/86h
znCScXEpmUAP4z5IRyfalgD3htviztawyRt7Ub2WTC0g9yMUExYgvToDUpE4KIAO
xTsL/piwOFQX81yO/DouGFIzOdFZhxdUKFgnbpWoPCY5MnoT28RkrKO/5pQhZz6M
oLRBBFD3e02hlrgSzHsj95Ho9FJavCjdmhmQrr7jAMQ9DAkPeCAqGXdVMk0FKi0F
P6BWgeETxNlSKjynDPOVVICecAZS8hxmt6+zA0khK9SVrVOuti2GtELFL4EV7Dbr
nxTCRoko4NCnCR4kqRjPCtjcGcWl1k3v9iJQLOlT1utKqpvtn4lqnlQYD1FDStIF
CVufkNWaRgIba8224i/9jeOXxDrMYcabkva1VZZIIn/+eOhjD6YVChUn697i4rg9
gghYsCpstKUkT0kj3gmgeI/JfrjuOQnH+i1ydFImkjralKxA5wMNpze3VCtCGbwd
WFVenu8TK7D9otwNqlIt8whzH9WCE3yW+hvQOqZL9bI7OXSGYj6ku6QSqp3AnXxo
BQIN/mANrCKMScYd+zgBn/JjRu2a9WLDb63QiNI92vF29taF+l/QwYivVc4zE0qu
0uAteWYypmlnRzlAqBghCZA+fVUijm2RuHy8vapBRPJgb1TOdn3N+6rSrspkyqtw
UbS8Z2acoGXj0z1rspAHq6EYECKdt6jh1xhXI5U10ZSxxpzgFCZqt+0S2VEAkqqw
Ozxwoa/0LCdQaLvsCi5NjkwHrzsLxEmk0WUYqFdHsvMeLad5AgRQTcD9gDmP2TPl
spk0Zxl75sG7pCn13SZJJpJqOSAF42zzPOUY/pPX5GoqZqEd3TA7pTIK7XFsKRIV
9lgSXRVHyUU4uPHTAJEcEgjN4fh6X0fpIn0gcSq2IgBsf3zH6QS0UN/yDDGBrs5Q
mrU3NAvCC1DtmE3vZlbW+GVPgdMdFbTv3PSseza/rNWYU2cJgoWwawY+smGrHggB
v+L3gtTlq+ANvYUUTEWM33U8+7aqfrZWhl+IYSBnFhSlehoHE1AYHtpJOcFy/ex2
rsILO8MfjzhJ4w9BOFW2S4Sj8zQLSvetdq5n2aHG32oURfFmI84CLD+Je2dIbCMt
3STf9zbWLxnBMnqCdOwt4tkM29WJAN9rrEbb38A0BUoEnjCA6fQ2R87JogevUkR5
BVjK2j7lG5/qA2VDToDXL/t/JDgG6xrn0qWIh7j830+zx6M7SG1c+8Nm9m83sfpw
q4WSmF+n5mgKVlAnE6h3EstRIGr5wvzTLymQRHmFrwvyZGdjV+8j/cD0FZi7jJ6U
PoHY30CM4Y6xqqrwVdjTuSIDdPTs++/ThsW5d/432f9CBX6rlfm++8bM0ppcxgit
Y4WA8RiJHkM1TBbZg8f9jGYHw04PmHMvUqqWYpJkBAByb5dK2qIXk85ygg5tkLg1
lLViWcfJj4Al4gsOygokFwFE+sr3zqIm13Usn82oc1GJy7IzKXnObnutrhR7VctI
Wa7YpVBeoPJzPiKkHf+ZauUKTRdNAjWe6SzAVep2r+n8nOA5sEWd7cChM0DIfViC
2MmEvfqkys4P2pxPUu+xv0tL0u9t1FHafbHb6yQDqLuAODptm2YIg/Fty191JrkB
slt25vvn6wWl5NFEw3qiPX7trlsQAHmTrH27qjtSU/Z+CBhggT4yvkx7v/N6RdnG
4bea63N5mfIY4iudCu1g2+muyd74AEHa9tFPwrRx1N35W2YZw5uAGQBGw64CT7BG
08LlnlbegxzuHcrzzP0/9NUWW5DVc2FutHXjxXVW7mE3IYkeohlzIWhe9ialoeeA
Bf2Lkkh4MMHwerESAxOuVwZ0Dzj42ZAmVhg5zMBv8e+cPSxR9B415fFwoZaPdGtJ
fc1aOdAqCfcnjHk4cP0xWQIC8VKjqIIetm3bXvQT11qn8Af0pZcGDDdaLWiHD/fc
oAhd4mtjCZ3OcQN8VCXaoIHC9hMR2Z0lrr+dTu7+26pJqRmQTT/CzHfcb/p5uIRN
+OsYtcqG+8xQbDqITSvon1vp1Kq7BU5V2t0PUXtAg//Te3wASXNDYvxOAkS2DYQW
uZuE1HS6Jhpq9iagPXL6fUKhUxAJZ0wlLoruaM4vFKSD/NZrRQtJ6LaDrP7FLDEz
lpI6inVFILOvBIVi9AD1Y2c0cZ5qCFK2LRMKd/TD+XfOfXGB4zakvZkESsgZdfBk
IR9WxNSHjAwy+4jBgxrvsI9NQuTkEPj3ZR9MYVsgHdnje9PtpaPVEkOBZ0l5jxUU
rDptWiRLxz2XdXFg8v6HO55VM0bj3hB1PyeLP4LwZ0uNkbV5KiiWlwaUuTpqF5Jk
DGYgh1HcTpu9kMZkSt5+hB3nK9RZ94vwVHHbz7NgE/ReQ6s8QFhSEW62m5jxyc8Z
BtDNp7HJp1tkrU8Fjya+KPvajSYu/JXRQxPAdkQscnsSbvN09/v0e8OFN2laJgtn
WtATZ+D9CDQRseFFL7tmOpsH2inkLZ5f2yiXO+Sc5u5nh9TP3/c538IYqfXcSlaN
noGaQS1tELpADKclmOM2mo6Ijj7zr1g9kGP35cVvcgv9L2qkPWC4ozciosRVdex7
ycwuEz+pLAAzkFdYeIrLX1bKBiFuL5DyJtHNgC/cprruw27Ksr9iJgG6oItmlFXc
xIFtgPHjbG80uR7DSMUlhownL9KhdZFtLU9X0cA3k6ldz46DYkMjGWOMtVsJugnC
tgtsiKKThEGXdCm4hoh05zquJvEsz2GcU/dzLcxRwMdBzRNVsVdxyxepIeDSD0uO
8YCFXxa9Wfmgnm4wZBmsJ74XVsBSpCkHdyYudN04m4HpFj/jIz5AgVr7oYL0e6pj
7nLXKmuyOu7oYRb0wxU1rYLVmnuvUmgJl/n7Fka+c4eBDxZH8MoUbnCyfay8JgOH
MfXGEzWQudr1jUWc3+ITmQIcJdBmJvdUm2HsmwXANPXS4ygUkGHYYtLCgKLXTwA+
DuZ8pB9X5i8ijVZ9QZGLQCFyCohqFxoDcAxxn9Zqfh8j0kfoxspgwsp8xDn+y6/c
UBqdq6Dq5/ci7+SLvYU5FDSDZ5lL0fkmEWHuI9D2h7yW9M+6JWP5cLj8IdRWCQoL
cA6FiU0Yo/6mSkrSqX6IbEqz9G17TyUjNSzwZbaQ6/PC5a0CviJIPEiCzjV7JFxp
Gs6bh3qpzFhsnV/AcZKSQ1Wbj11qdti4atEQedkP/Ns8f8hmGUw/bXKbUwqGwKb1
H/Z+geTd1eHwNysjP4bNlrsb4Cf/De6N/OIsINAkVgkMZUIbnhXaQePEGSE+Hc2Q
y1HDGEXlGH/ga72nGbz319d2F6Td2on1H1QueI1siSPAgIL/n44NHqjuuw4LJyrW
NVfVvD6qxd7LVi1Kjk83iiNia8ZHXuYDE7TYNHhcvbG0h0L2C4wbiIZi1rrxeKMI
qTY33TiFEKp/5kzTJRZGSX5YnIaiVfDzCDbxCSH39FTjs8UWlvaZDYn15RvaYYZT
PRKJNsHwct6M9NfLfkT8tq11IqrDR8DTNObqhv4TFg70WkVzMx4sYvMzJ6ARy3YH
ISWJLbubAbjw656u8zXnEOjXm3+1yn0lo5FuwUY+92kqHurfJRPfS3WmrWGeZVX8
I65hqh101NcM44fokJLWweW3OKWO4l2WUwbF8WdI3+H49Zssr5dNJOeH1GudXmw1
5ViEYzadvXk+JkuKfr9RWEDnTB8g1ig20dG5jSs+nY10t88sJ8FELpnfV7O0XCre
MCbAZDRxLN5r9l7qVW3q2N9X5VwUGkhwu5L19y8D/d6bRwtWRh2F86WGSZeasVZX
ckfdJAU5hY8aC8dCT0H9J5aCSsP9g8jHNcn9fpcxs4kjy+gTArBkRxnmN2kkiLse
p5Ymd9l4FQ7qefu3b7mXgg59jSR+6V6WLvRHvgtq359xSfAyYowmDuh24ayDatzR
ONpNvunerbIbnCdbYk+d/OSqwTK987Wi/qiy/XunssRREdAt/sTzb4ymsUqD5wvh
VTowJlIHQZsuTV31klxW1EroVsSMScuiOEw+CndffeEYtHv7EbWRsA5ofcnv25yr
viNoBcxwsDoX8TAJiZ3aKBSf/AcCKRs3LFT9XFM+wK20TVXnbU7kEjNy9Scz4tf2
uDHwtAYaeoDvfiG7N7bSJzA+aKn4SMVmdd5uEJK8TxHxjtnlwICIDf3HmZZ/ip8b
N/WRt2HvBACwQqSeyo54yatjIftJyplIwImc5zLqxkC5FrSf+AwJsqVmLyoVZlw4
itQPrKQbxZQPwriSrZhXWukbsUKCe3eIKX+JAFu9KLSyjuGfPH593DIc44gTcKVp
IAkGAFJ3nZTPAgGtADACmqRAboQrLsMmHV1bgpXxJwn3X0Z4wHod44zM1prqETBu
g8eygg+6kVF7yO2geNjiU5jVBhB2COsBjoiggjWbPhI9yj1p7KYWsHzNgVom9Dm6
bse+7Fu+WLpK/vtt2P+0h5S9g/MLeO8K/mDbTeAjbKPCardc2qynG6Ay+XszAqpP
fv0wTRclYESidIH/mIyC970lBZTY6Od1UziV0dQ7TjVsxsqVDSTc5OvGrvl+XTLR
cAbjN8jcQCVWkemkK1W6E+Qtb6pvG/jre9iyy/SL0r/jK/5GBFjc+SevxSPN2qVo
Maka9uNejKlgoG9qPTmXBT80xNNfAyXpJdmIfkWyQFQxHKN0qSUgZGTWcUFVkBcE
srb/7RugfDxdz9cExkTJ3sJCT4y8AXrfnIoqe+C7lgoO5qnQG86/Tg8EK1p8rYuo
1T9ailbdNvKRnle4gu79mpjapKuxiWq9FMQ1y/2gXYhzwlrSOtBMub3mgFVgkXKB
YRj9R1afwQKqoIp8aDpX9fVLAx/JmD0p3NB+hx3jULNVXpa1oAsQZ4D33j6g1qMz
FVwDrWmKoePsRS+UPLNLAEkGeTjGWHFdFFrXvW7VmeCZG3+T8hcvgHXLySEY2fbp
Ay4vlfcaIA3wEwbvURfVPZXJ7otBRKNsb2BD0t/CqwdA8DffH/CAUqLWSytexOit
4AqHy1bF/WLy+7bSWsa7RGtWDBegXMxA/IZqaX+OO7TSbTWnpA/pdomDkd6U2Bcm
EVx8BnYNluCvgl93djB77MY+hYbA1MK4X+X+VsbT+41EO0iUg3F2c5N1N7c3z/TQ
TWTmtvIfDBLJtZr8hFBRB8tI6haaNyZwYvy3ONONekrOVQC16LY2NDob5A+8ReQZ
dPpqS7kYxiMXQuvy7SsW8qCN3JEt6KhqYlH5j7N7HyBG2//LA+QuHy+qsMJ3XAtl
oUplXIU646FNyO9Bf0ZAW6Rd2PiD/9lDLG7eTz+53HHZ+4fg60tQ4F6/WWv1LNsU
UmZ1XcA6DUwg2exFfdW8cuD279CuqDSr9YxUxWU3WTAqj6K0M+rb1scwSzyYBY8k
yuJVGoile3VjMmIizxjeNTyGVZexrIKi0QgrI3zbyyLLcEVxByF/u6kMZAtX/eLf
1y+iGSOVOG1NAy1n1aNOFFaf7eR2ZHfHlEwAeNA7/ilOw5R53J87Z/Aap2qE3z6e
1wpsZlkU3mz+uyJPGm7VJZguKXUnnunkNalfb50XVzuUyA+Z9rBWVDvzmQnOEnKR
lN1PpjA4nB4hakYkk1iYiWMNqzy8N1gh7hb+SO+b2HIuynBB4+NyvW7PqWVTrdlM
UW7+PzzbBWzohZI4vH3uiA1lsKHmPg0jqmMMHrO5hNyOow1W1v7VzgJP5iWGsyo7
TVgg249ZqDKzCqKmkJKnfSMgabU7UPag8Tr1h5DMvknNY0u+F3MsVo1oKV8rFrcG
E3PFim1rX8BJXG7IDqqlMMlbRFS03asi59TdPgiToLzKJkqLPUolP93Dsj2WzhB1
KIvEAFqx35uQaCHS6LQyG3HFhRvynbYzOsErpHVUv47K+Y4QP7LfQhzlLVxYdI4D
Y8/CO9sK52QzvXE3mRIOz7CCJkF2s/VvJesQ+CaZQvjFHaL/7Mj0qGPLYv/LimMW
jOPsWAMm8T8MMjJTCR1tcnDvC6ym7O59BjqfwgiavA1akOpkXgSqXA0VgkN6rcUP
LvWotpSv+tjAoMYHSKTwTT8FL9v4eH8ig3a6ut0N3mXlm4oAci8+F+x7PFMK97sn
Lm7kjYoi8pwtIxRzsjQaPxX6hPX8BWEAdoHtpGK8T+b+AGMgsTu6P4sGl4naOMKe
zJaVZHMr1uyYcgSwjReffnzYrN0YMvo3Rcnr+6LMB8YX/hRZaKSD0vNSD8TJPAmR
TT9Nh35tl+NwB1W2S7MQzGQc9UhHl24Jwnc57skLE7y7jlerlEct+PyzTJawzLA0
GtEVb0o/rA1qzFt3Gvk//v9gJw99wd/JhEjr9PDEN9Y1mKOY9JVMeoesYC5G/QAi
t8G8cM6wEYTrO1OeefEZcTKmow7lxdo6/3jSX81OQ4R7Q0Wuty9MVz82L9/iPINe
GYuyS7sPvX0gAEE3vPG/k3XmIb5fDV0RiOyubUfe0565afRAscgDiWiIPgO1dGZK
HwrgWIOi91gapqDmi/s2U7WUXPxj6c+yRHZuMxCO5F6g4NRJUL01SudepQrHX9k4
vXubH02styD19KT7mEpMy3w0Sxpvuiu6srOQVI7v8jCjP3wUjGXzgve2TUyGIcKJ
dVYsAYeIobs/4qLpxP1tu/n/TopCEBof1/meaMIZm8nKx2azV16iWUsoIcUtejVo
8ElVrWP//SqAMP6UD0VwOqNVhGdpavTtiIfjtsknKggG8GsdAGV0cg9Oa7K3mcD3
xEvbOKOn/b8Vdy0PqPF2/pPCVF7AY/7dSKa4IiGozL7JxWaa8hdz4IfCrcYC0fZV
tf+2OfNOHF43CoamHtg3thCO8+NQJXfa7+D9WZsf1u8K77SpXZiAaU4x8hTCW1bh
IPbjnPumnslNKbT45UB1h6uRDslxuWiGHXjQwLYpzdp+jH3sPLADwXDBkwjCWHVY
U6N/+B6hfvUOjLRZ6VjhTXJLCK+yJsjLwzYrfNf9/rW9qnqMr2cY5s23I0iRGaHe
pGIrTd5cJL7vOdqNOS5puuBHdPavT92tXDELHk8uG0Ywvst+nrbrt8YshSLBYWmM
BxFIxo5GVuo5imOtKQGpwZXFK5ohIcf7qS/jk6Foa79L8J6nR7VMXCbVD+RdwX2d
vowOdEJnkl93nc5EkLWGp+DbD9axXLa3zBlrIe1Tj3RNh481rerTe+wN5Yn6OpVs
MyBGALWmF0QdOdoc0uXP6hX0fmoCyL+nqEMvSVHV+YNdXNfWf1uShOZ6YQiTWJf9
k9iGHnWDo2ygjBarfTHl4s5j/ocNC8zbypdt/PZIx7tWWYL4hMUSSdSw+BlQ2q3p
EnxNpwD0wC0xJLT0UuueMaMOCwhktwodfVpSZ+R8tEDxOg5LOdZMDnmkFPSsoxcb
aabgMxARl2JeNySUJMB4rPZhj067GESkKbdXShQZlb4G0/Yxh8YY6VAYeqiwajUu
OkKsjTys0xxCcxv5UM6zwxZUCyqc8yN+hVGG3mY7awM77Orep3ehqCx+OX3iHgcF
gDstHFoIEXBV/XIZCQQf+PDQiJmPF5DPDGjS9fDSjpKVt2hID5P/T0btTL+soI/S
jPB/JQV7ptmt2ijinZPaVrdA5md6cI1D/y+gR28q+eyoGPywO7PDuL9CKYr+kyLg
AGO9GSI1DUzM3ZrTpioC6mCLOxT6VGr6gVN/vrtXHR2DJoO1kCNvJ1L5traAD41j
JuJSQ3Uk+oiT8DI9I7VgC/3lcjBWE6ZUIhzt2V3bkfl+tM8XsBsT4CdaFWXVxuht
nR81Nnfjg9IS0qNrxe+crTdPZSvjLVoW0RD3gwBZ8btw6iXc9bAs8zytAV0ukV5P
j0S7PP7qTHmA3kr14p2QrVr/Q0PcjgDNUmENvtxY0pZD/FeGDsnMrMVx+d+XZvPQ
S7Ze4VSdXE1S7yfhSjTFobVd8Uz6Pa6sWfCkw7xZvz9ppcBQlPCKybtI0+tBRjuN
oiqal9wckcGUAXUvhoXH3JGP0nA4qPYai+ZZKRqgpRpUh0C6761f+wS9eaW0IAUW
DYwMUFkuMl/XWdsdK+u9k9GPfYZ+zGNXyIsj5TmIAH7nAOfpGhPHuGRCxb5ejML5
8HEzFpFLRltas0qZobefbhBgxNkGPztn8lCdhfAJQIthAVS1LWUO7EPVwEK1UEzd
fM29YvVW4WWKmwWAVKNcnaEufvPRMk8gG4cGcfoP6CbIna6oVcMiLllaVk1GrHR3
UfYl+wDhmImzPsgx1Nv+wYcKrJBJeSVg5yzRndzxwrKRD5d0DrOrOSqgPjohjw7w
j2p3YLxUTfJoscn/R8RKSRkxF7zgZjpIwn0e+/8O8gyJpoUn9u/5MOujXSZPHwVd
mhNY4XQcP9ugaKmTEYnaGUuNmLRGyakZYpPjBsn0QR7kXOjtGNY5xu0pJOJx3HVD
/PlSyIBqmRYKdb4dS4N0Ly1UmncEZM1Pqx4U2WSN0D1POiSrEgxBRgcBuUuCbR25
gZc//kYXUw5NFFKf59Xruum+u9TLIT4bABFl2eZj/S1RVYPqtGbhOwxkt7bf7IvB
rsqmi+FRze7MReoa+uYQVRgkaPqc8DU7m4lXFFgsO8cX3I8bM3gWDU2I7pLPi3gd
RBzf8auNHWagkkG2DwFzSiRjYu5I9bWytyr5GM+pwbpEUf4eUfWp7+pQf94Cn7wa
4YG+7qSTxGD0Tv68TkJ8/oMpyGO+GXOF7G39JWp5sVIooscAC2DcAjIB87s3f518
E/VmcR6PwK+vNkwmjHeOajvAtkvSFUffe4U+jLtPVHl66mrcOjIAE9h9ke5TSd+Z
ytKomUY3O18G+49Xe4TGTdT5ki3JTQgOLoQedSIsf1jPYHIaNPb2QfdA9v9jIswy
olpebuTNS/CN8CSigBm6YT9gOjxMm6yXP7S4yhucXZE4XMwMYJAuQbTAyY7ozVwn
wXNEFn5YJ/Y6nlTx/T/23MlCfP9PaK4LhhQdXANu3qqtQjISIdBBBNTZ/BOGQt/8
5dKYel1NXVQ5wtimy2A9ZS8oemZ56wA2fmnOAK0mMiB6s4+E/DJGMMIEUSPyk+cA
YBe6SmkRY2p1tI4eF9N5YzPChaePs4AZbNhTGRWsuClzBU8w1VA7QyABaqqWdWNq
Ics5al/dL34FhwjMb9V9+dc+jk2zB3sygNTj50GEpyyCWZ/0mTlqvqzss7+JHnXx
ALEbPkO0lZg2CNSeiAuFBreR216ie2AE4LGc5o5SFVsQAqDidaZEjYri/jmY9bl1
K6LbI0FhFGrsrC0+UTveG7vhsMk587gHEHIOkwYexEsPtfXA5OgxmcLOSm9gzLLV
5DX8yUvMw5nf1DP1q+eZ3PceBvURPTbHMYXxEKtNjNw+6/9JPbaFI/pP0DqKXSKV
1CDMZ14vLIXJxlmzEwFE5mleN0IIM9aBbB4S5on+TykfS9Cs/RIc29l2fAN/05kb
edKYc0yO7S0JD5qyP0OuFEs3qs14ngHNIZhKnrgiJzVxk+nQN4gTH0tp9pBZVa/h
cUsOBUNsZjeXfefjOOITtbaX7mh6Xuj4H7dz9WXVkL92NXH6gfbqp5RTyFo+27Om
5Vq8eA1hhq12X4Q6XM23/6G9E7xSV1gSVmR/cgNjqRElor8tlUvXALo7DOpmxpTf
gIn/ikPmqnMPGEfAzC+FZMmwZEJ6ugMpXLqo83dEjatzkELLVE/I6DoHkJ0yOFNI
ut0GFnawXPRGWfIMTBNXChj8NWzS2U713aKzlFOxWOEuG2VkO7pD32Un6kMZ1sVm
vVelcpkMuAN9ZZMwI6dwDYMkIMy8uuiU2t0R0GXB6CYTrsGXOHBJfrqZxhirhj2s
JXzwA34/QAVsq+3mMOI5Ng4Kjz08x3exmip6ekhewpkVjvkPABznXaRxM7YLXgbK
Tg23OWBiafekaw1RWAeUwfZXZckOXB7N0OU/VtwVYgOPqUILoi+AfUJ1gEuS6ObY
B8rfa3llWuX+iwofYebPuiwZ5mOpY8NPqjayFsnar8I5X9LmviLxCYfCej7a2Y5h
/psymbeL2OwKI+IvcV7QhIngVOqFIncq3QiXC2MTXN7R0h0sBL3olADNRCTSvOO8
2VJpEoCyn+gPl8GbiS42otA+AwOcwwgOhex0vGTY44o0I9buDinzByLzyqAxvMyl
4309EOY3vybtVsXuX2c9uxVMD0epkv1Ovk754qr9MJX69mHhDI7/vP2h2/pCy9S5
G8g4M8WiriNqzDb2hy/uIJBnoEBVwl+nAbj14Yr5PrDMPQIWdv00JS/TvFSwnnYQ
teGBGMKWAfz9VLK4hnc7T6Qwx0BsYS2580Jw22bWVMO2/AvjcmOvJ7Nit4+Pl6MH
9c+pmDhYaw+9iF1Z2z+2Mi40CYuxdG2WTe1fuhQ7V17XZg3AV3MGvESDCSANHbaR
XdEzcnwRtbAnW8XD9Lee4+nqlL0G56s1Ht2Gs/d8BMqOAYVL72zTmNmmw7akD7/A
lt4VF5RHxGTlAvGXvj2ghhmh/7r9M0v4YFu8nzHGHjBl4eLyW+S8697PhcsENlpZ
RM6YHriYXdnTE+avqYBvUV2PSPQ1tg/AUyQUxnut6+V37vYyDK4snyxdR7QCAw2X
4xKmkVj1PDBMyRoyDPXOS3Fii4UvT2prFtsiGyEcF8+lm2XSjLiU8hlATkRE4rxP
TVgitUcIHsCc8oVU1nPgKRDOCWAIvpEL8GV+BGBiRPvUgp788wiauvps2GWsc5EU
AzBA+fujbXwDBM0nnM8nCgONaU8I+12yeG2ngE6JGOLW8o0oymcKqXffRabIzu0i
sBxZBUohWI+kbcSwFUfAQAa5+PSyOVV5aohkaeZ1gJ8Tm74oudXxXXM4ifhl7zzN
1G9AmdlHnu0uxSBhCIVqhoPaqimNeDHqr5irkwCNEJsBCT0j/kQet+/oXc5/zzm/
fosHxdNCzWzl/oOpgZKf51d8E64Hm8ISGpXD5NZFnlxb9BCprTqppIQR3EI4b4He
4+PSFIhmqendsNkVQRBcHxzEQOhGlgKgYJtNSU+TTWGDQjbhhY8FMcrAsSWmUs00
xkcbTxdkc5VWhkuNT7GKzELJsFUDQH9/BnpOrjKZLYPkQXpJUuNKUZo+t2P9UjCD
zMOM7oWsh92WXw+ewo+g4znzR3ThlfkIMyQ+pGETb0Q1YzgkCLN3kHxO0h3Khyoo
aMrUKmJ2e67Yh5Qq6bHfmEtAndhXFl/POM4OKhcNnd2djQF08+eExgNWZjGuS6+/
51W79EgXb0L88lbj38qcRjoQxGJJ1PJ4CO1Pb2y0PIjLxsy/fZ8BthudL8jfoybE
9J3zy2xG5n2HBQnZ6WH7XrfluKcZQjv7a8l8JP6rZx/ftnjHLTltFJA+QDVvVz9G
B/rN8w4mTrMTlH3Nq6P7Ng==
`pragma protect end_protected
