// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
iE11KVKqo5m0OlBlPuSX/KRPjHoMuY4CVzztNHVOeEh8xF/lNCLL2vSygH34WyNVirma2s4bN7am
LBWQDoG1L5GqpEgm8+5lGUsM3LFbHw8oHzz67K/FElxMO+PcxN5GTb9qM1Lw4k81IMAm2VqCOE3a
A4mFytEw0cOnYyt2nmKfrHVwhalsKlX10catK3mGA/hsaHtivfHGA3eTB9E8qftdMBtFDrG3ZfpF
qYnFjqOXs1quoek7cyis4n/Aa/c9m3PFBMzbmWvw+jH7kUb9yfYGJQRtQXy0dAy3fswtZFOkZGIx
ZuJ9+SAcjTHXVfh9bF4SavCG3Nkrf5U8apq8eA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
PCVBReywFh9CGMdMAMWbGo/+b9t8oy8IRNue8gh7gwXPKU8N9m1rHS2+fkyisBBAMy54gYHyti0t
udskV1EF8dkTtnanVoU6UcpHV5StXXlkZfQCLEcBPDuog8qcvlHb5mS8X6ipPk7cod33J3XWPt9s
we3EZmYHYGGQ5um6wdKOAeLY2n1gfkwlJSySIr+9/4/H8CcPHK/q4ubkZT7U07ff1GvrCyFUCUfH
E+lNLfR0NDibGZjmRiFS0kPXDBvyDwQsTLAnN0rGoxQPJ8aJJYboTtOe4/T0vgwSVhVq/JB9BLLM
IS5C2ncml8rZZOntgrRAgDWIF2K2Th7+UlHGp6kvX1tUCvuSRlJElQD2fCqGOeAT8W4RAUh/fxUX
jsts4x9WvOjQwdyubqmNWomOXSAR8HMbI6aBfhKG3LZB56mRUqOM3Fl7vYrGE6ZLqZbQEtsSjq/a
V1UMUnuqIAEJmCwCnYwQIzz5+vMT7pRqH3QOGVhm4bAf2vEtKHAcn1V2OAf8tWV27PHEe88eHWia
+5iqwV/A0kUKWa68sQe7aH17r8JFgtxts90CZ0oQssWsDvtsP3b/FgFxaFWsQvCOIuaIiXvqOvyF
fxX17yRLLDZaonam91D0fyNgzGXldUXRShg6JboKYynfFPSztFqaRAb93G9Tza07xHyThcl0gg5o
xW2RFgVibRlmTl+xYfUPT9Djoy4HeWbE10WGkFsp29rzQpfYVJV1GDdd5gRueu7ItIhYbawseHUq
r0r2bGgh+u9ZcfniwacXl44oRf2iNHVtqYYHVRxLZJyJbUjwTS9AOZf0ufrvQc+sExeXaEEJgHpT
r1LXYwQRw8PajhzGwqe7EK4EyINz3msBUaJea/oY/2FrOVeYhWaGPLvOMv7hvXFGUFfQZM9cvUPF
KSkOfZfkrL09mwk1rApAW6jZQwqCp1a4/MbUIvYswvBCvWsKMI4ldarMkonwP5treNhOHkO/zrol
FAD9f2DuXC442XfTqkuWkuvoRqLMbtAsYwnOUdkdOEzMQ2DSwps8/Tp9vUyME2YxYcLd5TI30Ska
udBrN2I9u1XDE7puCosjGuBxPVHmS8z/BbnQDpbE4L8ar3+9Z+jRWVKYAfSBvwKrcaUt7vByzf3l
qVcw2IUFbpYSPr0UPDcG5N+xxFSW7SsSiBjMVpGqvHTsvp9t+YMh6ha5nvx74vrmtZQ8BgoqmFAH
SQ2qPdjTXZ01vIreU48H7T1ISE/CiyC2v9Acc3BF3YI/ZsGyTfKtJEEbwirh7vbUgyyp1MzziSxQ
igsnfsIzFnVsPI4R5h6nlt74u3FvzZYdcAASfZscFFDxoLEUORKCVjcUkDBEQ7/hhCsEGwTWlhnx
bo/Y2lLjSEMjTf9bAfnkuZDuSks2/ezJehIxeT8gcCmxEhHkFBh0A57ErG6yJF+L1K9CW1B3Pnh0
e5mWQHrnundPLkMuox2CtX4BVINrylg+mq9VniJBeDsICyS+kkkEkWtN8ErwPMFXBHZ4uwxy0TLe
yY58BIKr3z+3cIZgVkefxU5tIIJA/7vkyRIUHThvreBBPNzBgpN4kg4ebhYABHzjsb0UrxPQqQFP
ruH+IXmfIwuh/Gd55swx9IT8KxSUDwGkGwn03PJo9VlPECh4KIAs0mA3HUJF91uL/HkNug117Qta
njcG0T/xAlUXzdBRPL0WYCqEnbFP90EhvAL5qCZDdg7adX1r4fjqy/ZFbLMKYkSCcOLRo/6jDQbZ
CJ/SXiicYy3cPr+dk5mFtut9u6gm+5eyuyv+axx6G2UN2ndeTNE1qxUKy/6q8xtIa1C9dXuGogn4
QbGsPz7g7r3DqsrH/WfIl5XXsJTCcb44P1gHjngDpuI+BygY91bBKdJiFwfUEvvYfnCXLEDgeCNk
DFRsy+ILsyBgBfIett4tMnLn1uwvAu8HsoN3Jt5EsuhjUEzM7Kf9JSML+i0A7FdTxzDW9WvKsdek
335JLPUG/W3/oqqHx+fKMjGaOton4lQv0lmAygjRVHJ8eN8a39A10ZUBRL2zZ2X456c4aMtTx2S9
vVdIDSykaMhKycEwnQRmUgRpcQS33B2vfnOJ3+fixOhgltTzSdNhEmvjRFIpGlnkVszBwwSglx6F
imzDzcJ8F8OOabS2S5rGTahM+yvcGVKA35ZP8sLj09pqsgQR7mth4I+W9SmdlF6HkPD5L1tXa6cM
T16YZ30jDalOGLG5889OmkW8TGq5BxuDsnHzxtyQjYwqCVMz04tWt5xV4EzmAXe8p2uMgKg0OKSV
reeH/b5ulPxslJLHTlslKZ6J6HnZrjpCXsQdm23HoEmzU+p6GT3+Sfz4Odt0ZDnT7HNhPnW5lzAs
vgoKsJc/n3I1zBA2bbLplF7lj8lnfXBcIjU1ag1eWRRwxvYBnHXJYbwc9/qXTeGJ+arXQKjP4TeH
HYHJAz5HtnyIReqO2761UvdeCPqrnpq1c3QTVyPgEIWiLtI1KflYNzws7qb5tlLyU5MG0ui1jIk7
5MfGvKqrv7KUdBMYvhtMcrcNnp1DXTUMn4LC4n0g71cih5+f2Wndga0ZdGUehe+oaaWeTFk2mqTE
V90QIjLhNfGfh78CuhWadaByK/X0iQ6TKeazQ0+1R8N+37kiTc5weAT0QB6Jf1ssOr3KoRrmqkZg
VkdQhgy87dJuS+xmkJ23wuu2M7Y7xkiq3/wcEa1wMX29FJ8NvUUSu5WAusAXz25ReYpFAArYbJxL
O0E7hjlUS+YLlJRHrnXrAedYaiwjs1UFUyaVe0xfp2QTC3VhUdYF9f2LcD1QJnX+bW881PWF5oBD
7HQ2ySFICHNFG95ZrMi4t6QlDszt7H/eDQVHRieKJ4u/qj5ZJ+FHUJcicbcU0YVcGdtXJCAuHW7c
x9cNr1MFS0vAnXCDyXQN0JGkVOMD2CSRQ+Y0dWW4XzSJw3NKXgA0fQo5yS9YrI2gA4tqF8gNL3Rf
5eAyx0Ro+62zeqI52WcaPN1zo7KD++A4jdMBrb+m5hUWJJeZUpiQ0N357lcpl56t6/kHgZd+Us78
LXSwD+8jWBeW2Kzp0E9bI6Sl/ab4ZGi1sB2TStDkUFxvbuTdgHEzCEKD9qVUzzgTb1FjDSoeRmSl
gFgkUYRxn7Kenf2EeBxDJT3lKOC8J4QoUCOIllOOqdETXfBX+7ydZx7rRs1rMYDzD1VUvGfUDq9G
a5SBmxwtGkU4GQ7rVpRA+R4WcMuvBAuDaMD+b2rUEQTAfpyMhpVGjYEmiytNVkljRdssB1GWdxJb
KwRpxzdS/XfQ6uQZRA0SqcczgnvZ5gMa55TNVput8jA03cvDMvO08Fpp6gAjvBLxnPpmZvzSLUt6
10kAfhD7SoUTdMgsyKwtixJU4/HzWlwvvFwtovKE3W+2fMIUpiw+dPMyYru+jqvhoX3DqEyJwncP
mLRGzxDDCUQRrS8fz01HicIp8Q6ZFYawt7wLyyDLHgpV6pbRsHt3OT44b5I/45geV+FiCysDhndg
/melH2tztBGOAQnjq0RMynZn3hihz/WiIHir6XqsioG9cOr9KVOJH2qXyb8GeDO3rvhRXO+XTaM0
M4NxqDpSPpEtKJCWfPcOpi5molzOGd8iHc7Ja1RXqbOKXQFsuAEwG8wZEGrXLONdOvNGDvyQi+vE
JjqjhCIyCtLUYkEQ/hSsbW4i6zFyDWhztny2UN5yt5Ult7ToJptLJ2y0I6hum/a4j8ACKDmlSNXg
9G/HovPbaq6oPumtRPW6dwLGrIfLb8ACEieVfjEzfbSf74UGn4e1p8I4zhaBgTxm8rndCpmCf/27
DKuwNgNsSNZdiwFBC2R5Z6Ue9IOs8/G4Ldfg1HMzYUAhH0B+M/hIMx18bj4hwiTQIOLWDsqFRtSQ
OHITrtV7ZYQV8HTLyUNcww1VPlHg9CUHy0YyFiSDwdRg1PXF0ZpZN1DrqiHmC+G70jxBT7cHRWCU
hTNz40xvNITplXKuzf4e3+qZux0ytKqPumPd6Z/IQOtI/GcHCiUPL27ZlskWjEN1jzBPkb/e3/a6
fvxzPl27mrFqxXEgmawvR/qKJzYyaHx0Auk7S63YR/AENBBmiaJmxLkYJ2a010xi0+KsJXQFZ0rp
XbArwMn9pa/prKWNUbFSV3Uk15kfAGhMuEZ1ZBqj51J4KQUX09PnKwgooZWcgE42ZCVP1AHkK0vQ
sOYoBiP5VqTFSoqVheawFzdmDZYzXass3LRkQmIhecXMvZ+Xq927wv4c6umsOACyX+OLXtPOjxTh
m8PYhvF9SlQysAE8qPwjNNSn/kGGDAomMLESmIQAToc5pOi5e0LNarljqxLhthdlLfhiO+8qDBbe
IkGiAJKSGGakn3izACVfxBVSiiXrNK+UKgV2/JhWp9I+xtWCpvCXDDdJr55tZDe9DB2FWl3GhuBu
XCn4pKkM0pwmo001BImqxEyJsCrx1fqyX1JYXQZoU85wlWOyw0m6y4jzyQmijhNqwS14VWNYktuk
gMBHsRrc8hmrMqJNIoTgLbZUNzqjYC0epoLCDFkgZzYt9QrkZ+ci9nmxUPUvH7Z7Oh3XgOGI6do1
FT+QR0thNx7ZyqmW277AbOiTmYi/6AZazGICGNc3vxIRZ4mKodPh2XIoq5ynp3pOAt98Pjgo1CSm
eFLu6OEvlKdEENviNFnjqxO09BvytK3jQ/AykDlj5VbfRglAqCey8pB7nUpq7c+krsAVbQqr7XJn
31ksvphUJor0g46AX9gjRU4u+JkMxFH8OTs5aDspBfRTAMRdsVxh9g3Iuo3qCvZv+u1mDUc6ocAF
K5+sqviHMUjJG6Hsuby1ee/U8Vdc2zD7Zyz5PpWyPwR3/TAPO7kLAeL/lyo234rb9nCKxyjXuVdf
OxC+Hl7DE/0YCdcaji3VioSZxMcwHCkKyooJUSf/Tb4vObyNZOx1tsa2hsGK0nMLpEAbOv7b+wGT
bGVvUamRrzN4p+Nmtm+pEi/3jPEtprYWJQWQxUwyCHWFbqNRLybsceTcbLB551x5/scCAPLwgqgE
It/Kjwrj4pX4QjLhDtvIRGCfiHApyxZLHzmRsOkrFCZDTou3u4Yz7yjRCu6LBoXPk+iWbUjfIHYw
Vlln9BjIdf3hhoiwnxa17tVfD4578boWESKPP91kEZ5HW8xKj1JN9/li7WSI4eyii97gC/bolRUP
N9ja8WG93/Lfa4+dEogFLh2nAnEABZPtBOtJYuICMWHGEot77HTzsMZOX0Y5GadO1iuPyJLxTbvQ
n4rNEZNpRMZFu8jdewo+7yyUMit3mlekuvmUTs1//ksA2HBGM5Q3CIHa7XYbLwgpOukwQyjxbyVZ
awokLotcGmZNcyimXHRWGZIuaRnhiNEiDIgxlhRNOu1uUSXQAJdZtjwK1vkI6ZJZGhGw2Xi1eWVn
cjFGZyjJjfmJBSKioKkGMcorktUN6Q23rb7BcAo4O+dN5YOGu7C5AWXiQNKCSrIIaeF8Q/x17bBJ
k8GvZNI2VkXU9PJTtHEDjFA0g/EHh5ErWKDvxl+RTN+puNbQLuJTFF7lc0jsKe22SgSuX/HmApGY
fWKAdSjyDx0eg1eJHCk7U9A4TyvW6Em6ux1Egku4Ec8ECTFwlPmQ9ueUfgfka8JlLuTtj/0Uim6P
bIFEDOXnzd0gCW91A1fQUcCvu+2SruMa2pKy2p0yFdt1seYYPXsAdLao2Nxxi9jc3LQE1d9pYGGg
9qZKyJplLJjnurWOEngmXgprvV3wXFHLjZyTi3GUlcQ5O2Po9Oq7+OIFUol5NHo5V/4+sTPtNUf4
51CqTJLi9Kja9a2ElZ5A/erX2TjLOiMqIfvW/Cuqej5UWIxVEXxAHynPo3m7WPSysnjhIAUXUnd1
icyIQ8Pmh7p+3gyPr7seYHdN15ju+4qJ949ZnU5o054OSIRRO2+Rrt4VfOPabYBj6R4DUcFhnnHc
5gxIfjdqNUVdC8fjIYtm1GGPRamqpbmEn73qX39R/SLYY1f3VjPBf45m45FMAHdH7Ik/EdjwTUog
haJIcIuGcLouSV+1eEqro5PeKsZ8mXz59TDAtGW53sf1cy6ItdC4S9L09AX52va1MXxyr5vmnAJS
jOl1eoPL+zTpQ6HCAVNaLIXoWdgip8jTbLl+HozvLJV2RYFXe+EaBiJ+zZnMm+qEqKeFJlzwtvKo
7+eVNzjuzB1Z7Wx0/H2B0wdet0ZWQy8yNuwaNOy6LINKEEgcBQSlEcgcYmNiPxpRrr24ysacO5St
GfxxDVC2O3Hx8MfFcaS/pnuLl8pEt2vpZ2VKlO9WImRn0rcZh5HG5kaxdg+vOVrUWyIcW+gVbdpU
/5QhrCid0ljUkSC6+Cz9+O9HbdfO9WLSvsB7zmbBujrmnHLRsxUARtgsdTUMPz/Z3K1hyOHVK/hq
p4zjpPaEiOPsfeOIbSKeVwml1WgPWca+y72quZN2oJkBSlIFp54zHk7NqQz0n7UvgMw0W8L+KvjU
ev0LuGddnmjX09J1y+J0dXjn251de5bh4VLIAUlHk7bGpMc+HYV7dl6w/ce3Jm9iIRJQH9ZrMzu5
Uq3XVQuWhWyhuWn/eRPWKA9PNZObI0ai7ZHzr/KApNWSi7VQf6Ky+4jlTx8NWk17bWPDOk+1SuDj
IF2g/90z9D11t9BxAXbDDeHJgoF0WG1nMiq8XlTz7dNy+vFvSJwbhkmw1sUk6DDawB9F49Yt++mM
T/nP/m6kqJYZUsl6//zOJgWwqvY/UHOKXaVKoRpNVmeK5OoOUvfDuvY/p1vcjjvN4Q2nZNjL8BZz
7sWVRTwR8e06+dJ+fkzFKeIxD6jFibgotQ/tuqNX7benWNINElZ7/RWTT540OkbPnufShJBM/ZIX
vBf+yx7GaJzwP1yugfan41xt/WmZKJYxIVFV/coLGZ1S9+CM6GrZS3mhZZEBOMwN9IcrNRr3oIUR
Mpy4OALLCvGfiRphvHhDS8gW78/1YhoQ+0GqqV5WHm+D1UMGDfgbwqPuav3DkDnomOifJ0JewXnm
JgDYaGLN6DvfDySDB5ef/BByT1pGnHHWT7Pq0cirbmdkGcIrGmI83JnBYzUHIkmlDsjuncoBaWNQ
uvQFbCBFCSrnN+zgT5vEOT+F2HVPS/MfX74PWMb1FE/CyQ6zexz/KavVxO4BKMhsXvWT0PFNsP+i
JEVvEAmovYMGDbkT0hdFWGqHShH2+r211ZJ1viT9X+VesT7iymXVgvhoe7uhHZCpqdgmrecqw06B
p00KVoYZF5ZnuabSkZH9ujS38WLfFsWZRL0kSPYCQFvdq6sTJWxgXGnp0pVGM+d44ox8QWFkCgNB
MYOX5tOGp9O/aYB34RkSgJdBrh7gm6Mq8i+Ddmo4jY91ziHZdCvIGfF7sydXf5wjzEyxhu0MMT2c
ZZRh5uQvk0n3RJFGtZYQdvKkkf2xyoqoHSak8DXd6tgxOE1Fn4DGL6aS5wev5b5vgJEbQMcpMbMt
3TFHpPiIwP75jTtKaGqQZp5Im6JwsvCJu50jWM47G9IPoLSl/6/yr3qZOb1ji8u0hOpyT2P61lP7
847g+m9EZzO0kWTICCJHp0v2D2f8GOaY1b+nc59lLPjJvxvxYPmW6A2wemy40a9pv6rfscKnvLfK
0J6bwqd5jyRDQ0qam2OEjJzUJHuwe5Mlz9a5g56FCl0R5bXtjHj++mWOP3frhpNHm4P/NAYTm0Yb
U78eJ4+zgPsyXAGQz5ADlR3BOT1y30otCULEtG7V273geJwqp16t6WmdbfqrV9kmFxX2eWuTZUbq
UeCWOxwg4PEW6yJFsV/gphhjJrAjBT5uhJLuY4QllgI2K5rn1L6vUVClvmPBiVThZ/cVcV44bYWQ
6GsBRfgV87poAEcN0rUUZbbLtyz4woucE3RF/slD/HBARRA1jarMPerDAznJwRLN3OrcF1OiLl+M
3/f1JAPYnaYwH4fqz5kxwZlEFeSh6Iik9uBNGwrNsMLatg1KkEePLd5cBRqlBEv0mt1cHsxZciMF
AASdkQPqN+pHyuDI26KZ6P5IaOV2nmXoifMbdOUDU695tcjn5uYaLlXoyk3ynYxw4iQZ54ohlLUr
g0i2KePs3XifFJRYgW9mE3P9ZxgUW1lCnbegyThYJFRgbgcVIMr0RZNJ/txVnjhhbENQknhwYjYQ
sYzC+MtoJz8uMiieVJpfiasMtkBE9jJyr33wYq7W/F2MNe7oKBiRkmzAjyt3OjNTdh7RAO876ch3
g1kmSkBGYUmlHcen0GBO7RQ0v8kMQbyZ7WVQ+c2Hl/uULoFQUeiTVLDJe6k5UxQ9Icw3x7U3ykqQ
IT4wnhqA+7pr1AagP1Yd7ZxzFXtqOvevBPpONMHZ/Q1fKv7XupGcecT1vs8w1Uqbn1JVy8VIL1H0
Ljd/aDCpehXp4IRQlISxFW9OeRWB3cNycAZfdd3Qnj8yYSGEE1iD1egA+hnkSc86NpQwkFud0o36
BW59JygSnOukpcETCy06DVOQa7IxP2/RvTpNcs03VvluQHwaBcknI7BeKIYtvWW7ghptwq8R/bzA
juqyMkloSWGrC7kb7YqYg5fWC72EN78P8jW+vVL50+pATzwunD4J8LHJu7UmOwRwsxiBfKaBlPQc
c38u/E5xeGBLj3j7Ix8mUsFEnl6EGQnvs6PVvDtSgtBJhfUBzyKvkbtz5Vznzu4sqYUSIAf1YSWC
hi5wcylNzS21JZRfAeAiihVN4tWMT3ZVlO1vvmy9w3TOROP0nZxnR0Kf3nHP5pFoUA2x8DjFsjTr
V4zdMn8i6IOV4PsRVyE6mR9d0oy/BTVWq0RAh7ir5amcCNBzrb47GKl2Al8hGpLgG1p/UxU6jPTL
RWHj5ABG/9DAYTInr/5Jjc6FQK9bAxNHDn3KPUEkIoZ3eJtN//9LGzmnJA6LVQfr8pD9BkPwnfMm
o4OzrmxCElSAyGbjT4bGlaX94Hg75Q/55Hu04cW+DWgap3gkpMnqiiA9Qa4OerMrogZKFOflQkrB
eghfZW0JckVwV2PJZ7LAoV9p6v7z5hyOvLKrMmorX8NkRMn8U1xAc2FvoipRFptYnw9TWIGx2nkS
M3t5FbffnUnJvhinsyIxSxqda9CjOUhHfaBhH3pmdwjNlvplDbfES+/i/XMTA3x2QvUypvhKHSHZ
PtSLDtQnbEYUA3U21GkFgK0rvBtWKpdsPxJ6aWcFHz48T7dAXJ6DWwDv3hf6VjzRJMw+oVli/15U
FXF9EqJpiNJSsojXwq7ib7yALLy6wEBWtJpWOcB40tCh9kD4NcpZXXRSoVKwuymrg18zRZChuKLg
KCKgHbRLKqFProcMqKLx2i7Ci/Ee51FeGhqA3uGSBxIdsDp7smWhgNDQsUOggou8OupK8hfiqLYo
J4B12VOLz+RwRVuwgT8WsRS1w1czFkzhxLrhGTPLWJ+RH0shygPRDWJgfTQKEb7JOWXgFWyLu5CL
CkggD5wC69WU+LNW6eUXcgbrunTjj9d99Ci0ctbWbWx+5RoHcnYLvD57UXNnbcz+2Ekz9NZYpwnS
5AKIsUHStrSVvCVkBJSSXeS3dttUPlYqFS6FJOhVrvlSu/59NbfzG6npRO4tqn4R6Jjerlzqu9yy
eyVe8jsCj4FwGJOiU5c4Y8txri1AunkJi4TI7e2ZN0008qeQ+CO8CciwMFsKqYqzYCmVS6c8kB1a
66rGwHY7YyqHcRs/BhTjhqCsm0G0qO1ZOtOW/S0V7jrI6kiAwf1MSmN5KnMDBCN6magiwzq6MpT+
g+vsqv3aR5xk+6F6sfVXeii3ZvH4+l7zbU+bHbnMVFU+VJNr/OvYaKyxzGlQZMdGlLe/JDYeNsri
wX87/9WO/oKx8ij369ETWFLombY8azvDSzMpvN65bzRDgfNW/sfNzMZ4bSPsPICaPun2FSpXnd/G
5HJm/SsLS2Ks8FudlGgZ0It6fGVIg0bcKmFkUvKfBXzzHjR3xyW2R/GFNvmUO4LmvSBkAnxFSVJv
HmWyU4viulag+a7dyKgDl5cjCmeDpvGs4VEbDR0eJulysW97oVWB3CPHHDw/L/CpoemWXbmZ+hx3
7NMb9YopznlSt27sS0beIk6lX/tnmUZHhFPM3XeIC5a1NR8lba3MYMS24vmWdE4pXrZI14hMZi2P
Kn7DBV+LmQZ18zJ+7GIEcMQgzlzA28TQ7RQGsI4XrVT7I/iOHwGCMgc6ukTwrpELi1MQVrHnPE6U
j5ug/TQDR/r6PcDvQ8Hovsw7SI6XKRigFqEpCe1UOWEUTGYlqXamOsSLQyzaWlaSbbSSrhr7HvrU
C/1FDcbrXx0jX/e4Wb9uR9zf+wRAUHEg4qIo3ZjcR9KnpIJ3mttc984HgEjWwhNB+BLDl+DfzE4j
3VkStzqnQPtEQ2BNERaXzvHWLcANfSOAzQHqPQeZSQ5y/QznlppRl60x9XnrGrjdTYX5f3/it3aH
Nin/zWfTvIb1Q13Au4zsr/BwrukNLkxMS6TM1lVwwDo5cjWxzSsuyEvEnp3JsH1DaQK2MvFFCsfb
6gheIR88Rn2o3oWWS2cP1dkEZwSfHfqKh/45ilf5WGKvR7BHXcDCZltlo0NoxqVsdLbyPxbAYHrV
Tdqp6Y+HcxouOLVyqBlbzHnK2SYYWeCtKRU8nQlF36ISqMeIqwwrFIYFBKZ6O2rjIqQvrEAPviEr
8mnxSlDIPERZH+WndA6s7olmnqhcATyD7uUhonF1MwAiMxDItSIwcmHZYnRQ8k7losDAq71WmXZe
CXvFcI7IwBNob0jOnr6KMc7piKvYdw6SIHqtYy8BZwLIed/j+iWXE+X0CLbrX3OSpcypQs9+q3/w
Mn1ReOqwZLik67upGHdpJW9QOZ1cty8yHwDH16+79HIxwcm+PzVUK5LnbJFPni1RXH/ukxdCTNAG
bAr+WFpH/hpnwRy9MVM1RYsWXXK9T2o8bon4EA4sR79ZG2M4MLzTK14IhUzVQK2nZycZns+32HeU
BjfCOSLI/ZS+U89ne789u7sitCeSpVjILAiCcnt1ru6YiDtEsT4T/Rsc47b2diKG7wHRwGXIJHmq
7Y0FkK7BxqXbETpoxdeTuTc/tdRAOTlkhQK8xQNZOSe067OiDWial0r3Z1H509/GfaGRXDHhPPjt
OicMSE57UjRz8IDAm39UDsu/WdVKw0rNgEB5C3yTdLtV2uoIsjgy/CHWNMkv1jXcjrJvMnevFAmR
f2RDKLV5HyfOMVLVICsZ2AFW+BXVuuk7WdAoF7lRh6uSZvA4q2b2OEjZOwFcb+ebORtmAZ5fiiNO
yE1fBwGYLSiyQVxI1CmXkTYUYy1JLtKtQrAxeY79HIkHcxhBjh5Ga/GbJOBnLPBvGc6tKTZHRqM3
o0kGVu3wxX6IaTfUTCLSkNOlT+maYn0QJf1gwhSex/jOg9Kj4fEFuvtohi3TSOk2WF3eMbY1p2Bk
poyCxftfteUvgewLhkaMRswO7WkIbFt6hX8TOCsiUTt3NJM8NjP0l7bcC/OkufLOvk9f0xPxfuCr
4uOJPrKe1ZkFv6kcAkrRN+wAzJ27rPCwOkEaOzCl/WH6ONPPbtQDour4ejnBDANLDE3CO1rI1XTU
WEOyVUFr3FVBgfCuc3j0InAuJvQv7rwDeAyq+SyAYRweFrCX9YvkSpaMgi9/B55sDyildRIeXVzJ
iQj2xJT1Gm26M7Q8z0yuZ907HytLkGa8I1GbhiX2fb0mVLE2QPyAWLWOhnisy1ottLe152i4DRns
qW/t64I/sagRgs0yjMeG6HvvvBga8qGnuIIanBg040QKOCN82SDw4RWGwJ5hIa6pbjkB2el6cNJV
Z0ZIEjs3pzlrqLs3awBfRHKrLHbwZEs2Alah+4ZaenQip6Hj6dWOu6BkG7YLJB7ziUY4TqDUoV1U
wYhHIsBh1ogMDbzO1VrokPftO4Sxj4oLIOFswGvEXke2zYJ2MB9NE8FtjaOS5p4hQ+LEcy7sVTWj
k66vnofcuUwLfHNYefOUtt6DMVDEesypcUaOhPLwLsv85TqPl3T94Hz3XHONpEXGPA1qDFO19n8A
rrqSHEHqb8j4sJNdUlnJU2YV4nSqWBcXLqNLwVWqzPbesx0/YJkIavA287+gZ47oc+CwuFwDcC2c
H79OEg6GxNLpi+2E/WzzjLlZb2AcJ2ouK35WHe0Y3Gfku42/G4zaKKJFaqvfg8mxOqvfi5C7nw+D
V6cH7wrN6KbXRSh6wiqb0c3ThzQZIhDEmomA3etj+UVrohg7SvBDipQ97ead2FR56MNxw8VBGdV0
3fVzpN3qHMlYnS3bA6dV2vBti1HR5/877GT8WO3vV9vx0Zcgct4Njwj6s3gDPWG6L3FQvQexWIRm
0i0mkoX992rEBwoFynlTl+XpRvNFsJC1Vbpos/qz1fpJUjAyDPjJLPhW6YzhSdwCAo+Eyunk86ZY
zsNRd+FYMl5jo4h7YVZecurZoIKtJL7XmmyeHt5hB/YkF/YqOrzBTe+1T8VWpIjhzOt7dlJvZXDE
0XwyhVCwiz/jSR2X6nOzyk1BSSiVoU4rg8P3IILoB5vd62iZTioCONV5XkoF9JSOs3Bjk6l9lf/x
J8+Jjy9QfAculx3ifLtFD58eZ+xTD3oSLMso8VyE3l50hBr+saVPvlsF0MRU0dOLVO350hgRMoFi
3ye+nt6Yj8VoOvE6pNoR6gZFGLKCZo5Bic++LeCgESI+Nn0g2C/4oPQFlWvT/tqIHJU86jZdHswk
eC657HQWD29ZBma1sNhv1OcJNJGJVl7LdtTsI8tvSA1im9tGwkNY81dJW7ug1CZ+Epj15nSnBSeh
JbCxpS/ybNlWFTr7B/gYJEm00eSmWS2RYEydJ/zwtn455rW5GWfMYoLA1E1cOee8SI5eCUgeTN8y
E4mI//SVISW8UbGSfS7oayZ160ASJhUWaSkH0e5iAwK0wV6/FaHNTFfWPWzHIvTMiu4y7RGwx4hE
vE8O7H13FloY1q2p/WhXaVjZwCxFTDFKXQEfWBOreBbpGQDgLfSCXS/Gr5l2sa5yF/9NCssBcxbl
AC8ZFtPyT7z6NQwhReQv8Zr2HSSQQndgm6OhpOm296rGYPpaDMwJSUvSpDkfaEzwZKnFCtpIGI6+
k+M3GKnJXk/xg1qcLshwIT4dL/eH9/Voopv9pmJiuuRt1UkyPdXB6LL+csTOV6eYW64n4XpYVlym
IwITannEW7K1wWfgedgVq2uKw9rEMLdSMA6PvTSyjkXo5LzjVL4NERiNCdj2rjX1uEFc2ZkoUJG5
/CPLKnK5pmRMmtbWoL61t3e+xF8/X3eT+hUcMbMZd5M6OmBuEaAk4O/PV1IxrK1GSszv5o+w4J0o
MO6UPeX7GLk9Ls+JA7ncDE9aejK6Xo8oSIC2KqgG0kwBxBA3pDI8nq47fcwTn8kbFdDXzBQUKmJs
8ftacehiJlNq+xjMxmoX0N1nMD15kvBd0Lq+WxqwP3yCGCzgW7yediVn3SFUeh299l2B2jYdpLkQ
UzwvrMhOCLCeW9T7xzgHapVe+X7yUCBHyLhsQiAQ7mzhigKPzbiyuYA0gWw69oC4NfiLw6hzDesz
BfxjodfGHl1goU+gJ1NVH7DA7HarUEs2j/lwGGv8mlIQYHa44iKkPWXziujSwPN3SqXT76djTGXv
JeNXJVZA6P3i6J6oSPO5lNFSDXBfYiYHEhnNMxw96NbY5IMHZqwRzVn6sHeRYzo93aDbPCvTPtZd
vpcnp8/ibJf3pbhr5ACiJJaA3UTxsKgTzLK6RnBhPGq6IyOLOf4ztCtn4lVaH4WvQNGuZubC0A3z
4yhTLa2OrbKwN9q42I5xJ9y0ohsB7bcE+hoKhgF77wPCvVH6VNoXiTUjHZ6CH9380C940g19OM+p
HTrl3Q3wn8zin6E8JvBItCN+n89EFuRoJFxYDEr7arxFcC4lmp+3QIEET9zprqdUDTL++MGyP2r6
FL70gEyK1PFjetfl/Ewzhix5fMp8JwWb9GTf7E8tf9CEaFO5wuBJbeVy1rWh0e+PxJgJxNj3aQJQ
jYE6PZDEAUhXQ+pF2F2/UdhRj3zKazryZHoSUp1vFwmFWlElm57QPu/PmL9jQWUQZGAUhOyLFG6K
IFbNAm1zhsJZmY62sYKZWZNv8cgoTMPFhcLdZcNJlNbX/W/2RcaCkyUoI5eX1/8QMocIDI8aas8r
Q5QXvpGfudMAptHC5riLhmMMahIi6zqAzyQH2knV1F3ibsyPN7MBBp/Xz3lQTGAugTVGhmuPWHjE
EM1Yrg6jFkIpUSLJzuDr7W5kTRcxRavp9nWW7sihfvleM6hh2n+oJYKRf6p443P+FKTDE/v1Xuo3
Ou6v0elfQiBZC02U4HcCK/s+clXQgEiieDYKy3c4mpWB1b2xfltICit53WdLy9/OjRecMA8G5hxm
FkKvDjGyH4wLcvaMIxLcMx4DKnbIX2X9HCdJ7Im7ypGgksPE/E81PccC5Klhn4sHPKzaEgLHmjdx
09YXW0QPOt6kUWc2k+Azo2cIPg3eQKuNwSORiNKTAlPETp0+WzrJJNyTaICC5QAVajLilJZUKLh3
CPjLipkm96U7qmTax7OTF62267nrRitaXkPjXv7mKCMor25zKtP7OJc89GZD9Fp5NXA9sp909r5Q
kDp8GFscq2XwJddII336XhV0bMNdzyP8smn6C6lbwR4BPfr9eNlPjrb9VhYx8eESPrxvpzCq07kK
ATJOmYqhKWXVZvVfjjqqGc5pONQ1YSFHL4NyPlvxzLTrHrhPqkcItOsG4CtImBFsKJe3Lzhxctx+
7z87lgc1t9fOksZ7L+PTuzV6slnNYcCyAbsvyiJ8BBwmnQDm+/9T9NWZEtGCgEPId5/lUQNh5q1q
XnVHnZbOBvufrHMl340RfO1Rp5ko7/rnZNXqeB/44nvuQ82mzQYkK86wA5ZRjC99jwsgIBxw2dp9
28ZmR7pxlVFbtZsG+DpZi4ot6JRxfLtBCLWyPgUJyosFNWEXC6moVBPBzd0OeZqgK6+nEFOFnr63
bkahxhfepgVT3VxIoUvjzLZQokoOQWkcmGaY5URcO4fgAuuWZGqoc5gidGQQcMTPq2CaIrmUW9MO
lLVsxRSbnatxhq5igcuDvtwrHXdy9RAQ4ameSiqeFmPbO4jrocfG2Dud4YKVZHVSjKOKf0IxuH3p
X8A1GS1mqnmCrGkJUONw2V+pMpyv90BGkekfoagH662FOqHt5HWh3AUSMVseXdITdfz+jJpzdlAz
qI4CzFkJBBt90uomf85pbStMJQmDC0aoFmfpXQhq+cqC+aGby7Tyl91mK76FyzsFYDyuHZytibwH
BP1TyarSyMs+RnqlVWwoDDBaL+a7gJJTd2IlvIgCAcokBRw8NNnL99yqm5PlmZEVbTs7K5kg9mjA
kPOzoiA73Rdpi+mM6v5eeK980o18zRj5PtSyoHxiZ6mDFgV/lTYh219hNygSLTZAe4IKGlhj5Owp
0u3p93qoRUSOMHGfbWS47R6NzkdEf91v2zJgTeVg4qeIyiUC42VkF69ZUN3r10+OamGPGrTFQDtR
q3IpKo2jpqBJ8qexGBUPgrCNh1GYY/rqaFHFxQnrPU+f6N48IkH0sF4t6BT126Hgi3uQsH9/R//7
TiveIb36To1qpbfr/xfybbonSlmtEqAaKebM5wjDUWPezSGmLOwMTUzkRVhGIq3RNvCm/NTyd3IJ
NT6BxemCMcz2v1JfDgxOdd0dLh30MUdh29FRyu/OJBIftF7D20/rMUplQDUhSC2m39RyN5vvfTQm
omU3hbw0UVXEY1ppGXavrl82jWnaxRao1wjIcY0mmtZDm618WApoNt7hvZ16aJfCJwCAw4kHneq9
7CpN1huiyL5E0nAUkEcBq/zQ2YJFMyY0a72pd/cp+1csSBxFfdvfQ8/jxzA8tQod3WNr8urr+Umx
h3eK+NJgqe/ZYWVwk86w6X9nkmGzgW9uw68MX0LBEDlwIy0YJOkA8RxPtDHbcKmEeoYJec9yBiEg
0GKtq4sX8VntYc1gHX7txRCrOP45/bRroV2kf/Q/rHDLeOJ/sjG02xI4j+UmtyQ1O/bpka6++W6e
kNbtELu9jnmiVNOJ7fEmQmBP9zr7kA1trhwwivMMTlkLGgTnyL3KNk5HnM6xcIcte/QiOTFGACv3
oyDKgmtbiL4Y0YzK4RdDpj7xLni7PwkrKFAiRwwWC8x4waJqzC+D/jCHdulY/II79bsA1vAgavL2
IP0qb09jr+fcwYRiOrSxiWhgUp5y/4Dp6oBZgCbqWjyV9v+1FQPK9+jS4x31YEOHDMhAX6PjvrEZ
ic8Su5K6DIeu2I8lVah1kjLKPU22aZArD6KRlveDCJ0xyCeZ8RyHdtcPLGD5UVgl6Drki2ny/fsA
H4rtN5pAWjraI5UeaA6n1anA69Jf5jrZJgbqtsYtMdfcCxivsOaM8Wbx70I6Md6YpnKFfZPoBu+F
tphbQWvPhRNUrAhJGxiLngeJyVllbACMAQ/LzRZDyi48sbtAltsIg23SVWnQEHwZ9hSApzxHzOHN
vFTRAzCH/FuBppyB+kR0bWv5Mf+4uYExicRIu8gSTCsPYP/KPgnEiBUA7Vs2cg14JegQL2E34rJB
pPQq04t5XTqPC9TcMgtR5vHyUHveyRM6xcYlvAlpcpeXMh3urg9csWdPFqet92t/32Jqni9UbGuc
1nBG6NMMOVDFZbhDVi6Jx0UUAQvqbW9ah4E/5240ZJsNE101DLvYBqvncQTIj/QpaxIMERM1oX+a
WVxjUOicZc5whJgPjBEWwCPe2XP9C5YrzZmp/DsWgxAxzAytk67NqfVW6W+/c5fpZ0Sj8blDW4j1
X+2CxQAR2N8O5YX3Uspm6v4Q/7K0i5ex0mMXln5s60cXtBquILaW2jMXiWI+ldcjMJ0V9c/I3KsJ
vcenYrFUvGoCGWTAJHy0m017r5cpHwwGPKCTOUjzz93vaOMVARrdaAkpUTY6WJZQnOeoLC20ikr8
ymrO5Y2YE8F62gr2z6k5TjYgJM+/Gda92O2omIGDa99eAdbWHQuyWLKOouU7HrGm3RmeO4zMiWv4
xhxlPKGY4tw3bb0cHpsB5vIXD4KRAaMgmJrueJXDeqmEJ2Fh4ibveOHXyCgqFVIRfVwThzjAz5VM
GV9NomMdoVkwfHrJt1v1AQHJLGh9b8joGwNkYMP0kr6rOpVKbAMvYGWAmMbw7ocITZ3m6epB9CH3
inKipRXZhqnn2DVKRz7wNsVKWYmAJhih/QPIwr2BU0BIQYoePsjyQ5//tJkcGJB/9+P82vxxxog0
QLwqV5ZC48NjuO/iWpIglHJ1qZBGUg8mQ3jJvCnfeOdmhn5GCZ3a/PcfDMGSCeCepuxdlTtp2oOn
wWsp56kOkVlsX4Wg5uSrI00f0Ce62h8dZD9bbGS6wXfmEXxpEeA0DD56qXPW5K1yXAcIrXV8tHgd
KzXU30wQNSaIQvBStpbB+uYZJ0kkYPNhSILmCBdTJHqwBgn50ts9az8xSDB1Y7QpKdx1ctzbtpHr
BSrRPdXDYJbIxFfZLfOmPhiq1qjRBBWuDH5FcVk/1BgaBV+JFa9sX/ZjDugxrTU38QwraXoM3SVP
MGRFsT1BzC/TOD5jGBdDiFz8Iq7SOwDrzsUu+fQLQ6b0aAoXDPiuLcawTJrHvNMMpPMYt1SqAHeR
RnSs05yOynkpDo7aFi/taLGcHYfsAvKRZSkLbK3Zf8XHmwgpP2jRmuPJlnpAb8hU7+33vYnI8jTk
DiR/s5li2PR9yghvlf9+LWATFKjQSM0ma0WGY798T948Lssdb3T7wrOSBsobQ74Cl6Ye6WDF7+4A
ofpIboKGPvrjIFd3cxE9/ch133g7SOr/Ebl7x4NY7+fbgF/n608OHCqtwp+Xi99rkIa9mS6RfJji
CQWpeJzuf4AwEX0xG9yAK1evfhjwOgj6cud160w8CkboWrgpUsyJN78iOY/NtsqwG9mAMm4NEahg
ZoN7f1byRwodDZSuGrLkdJ5shKLDSF7kyasXQkgeUFcutGd7ZG5brvbrVpNNm+qVXTrXVO3jSeB6
etYNz/83f+P2oX7Gq6MLRvytz57By3NVLckgxZUbIGH44JaUqUlCULEj/YZqCe+e6BgToMiFfi6e
06kQ3BrC6nt8pIn64MAsyGVx81MySQTsZ7VmCbZFBfsTwQuptJMxfXgCdFmUV7sRKk/dO/py9qV4
+4JqzEF/WaJMo5EvisfoK4GRnXPDIfnKZOmUlfScLvtCRTcyQU3fbbDmdA0Mb8EtomSab7SX5EbT
Mo5nS00AKCY+nP5UzMcK3N6E9Mu0sB6Ro9a0A4PvEHrxL2ZTGvAPqutpm+J9uMLs/1tUq1TwtSIr
7UvXNbX0Z7J+eqwb+rjJnrHcki1flyPHLsKvxQR1zo1JlcriDpBmj/Zr7nVMp1W0gtcxKTixm6hd
1SCVd9HSs/qNyZ4aMaRdKQnbwlDrCrkURSJ6hJj1sxo5oTqBxS5IhjDxqtPP10lwwMMcOEWcv3pK
ePdODNbrOj6GVUn4hdp2NJSAO6t4W8UfQ2QUtm2d02pn3R/lFF975IOl9SwzPBIU+AYcPm5IPBMS
ugbuvj0rBn6k0p+DxzETdYlRsY6MH7ixmVDckVEKwkn1THJUzgemkZSruw3xyiDQvMG8ZJQTMIGC
14USiZqHUJEKqkIBODEO7dSWMKvgly3Y0JjCHlEEJ/4yQ9EA7OmY80hNdZbv3/ynvBAe9RIKXS8/
R/pO52nfEbrzhDUYafqtA5zVwdWaCbnVCGWFnA2ou4rTTWX9BOhn3mCP6pTTogYvtQs7bxOPqU5T
s/r3MIPYpRYppjwUz0Pgh+WnA/lH+PuqEmbOoj0wZnx1nxVatWUq5FxwVX3yzOtluatd41WgdNDG
HwzibwNJeTbUyma7eK01/1TdqAN2n0PwwVixO4dNLmsVObLlSxyFd7W93UCJkcOCUviZ+PRToqZt
BKWZmKDZtdLoKMoTvvuXf/t5A8OM8N3SV5uT7pflOyox5eQ6BC2Ia+Ht0LmHnQMU1DoutcFFgRxN
bIVSQCbgx8PMBhZkdRRycvhVX2QdV+8Qjfy+aEQnvWs8v1AwUpN7s20olIZSdBpKUf3jTQ+GPo9Y
aDIsaNmzFTmfWK1qA0nW5/4xgsSL6suySUgf5YFhk0OPgD8/xCc/QnZ+2OZcYOhXntuIA3PfkWuf
WI1P+EVwxjsKwygtHiWbxs0pykvM6l4UIRAGd0fgANBVpGKcYdxhsqOA6KF5Ml9XJlqE4xJSMN/8
IJyzmR+zj8GpQb1tNmjpcatSYt1lfQIZD50o0vObj9GUsfSxnTnJyBpXhF0/GtNG8U98bQ3n0M3a
PgoqZ79Cnl+bG8awlrq2QQ2zih1Nqz53sWcxqubX0ygY10HHefpFpwOMNafFo9vjrVv1LETpbee9
zUl2zk3sf5UB75tfQymMTAlatGkqZAGwA4hkt/uTr9IE9Vnxz8LqhnuIObqgeleyN6TDF/JpZpCK
8iVPXd+okPkj+xKyzcJWsrdcszCrPP6nfs6WBc41Hk0NitxGuIxibu8VLXQOBNo6MZiV3rmhlRm/
aRxd2y202xD0yddwHrikTHLw5ilqgjwfY+nT6u9ydzOwAaUxv6kv6kvmviA82oRBjsZmpfbq7j0K
YZMP8Qu7ktskS4R10tJE8IWpYFp9/9gxDe5b8ho5NV7ACaQNYlA6ABeiy/DU4duEI0lGRRf7uDnD
+Pqha215v9/IQq2wr6uPXdMjACRbxWUMt5AHPSprIIb4iHXQj/AioOWMnykaXtETtdGQFiUAwkVA
WrAtSIX3bs1OYROpAuCbZRD4Knd8dPHRDLRYd4LUEcuoTzNgep6qggQvbCf7zQHhBVs0eP2MCKh3
I22lJ8hYqXd/cCDwIoXzNNMtCUdcZe40vWlQg3okrgo+Z6wrCP/gNrCn7hwk9J3cWsGS5p4GhLx5
KJZQyl98yzJzsxHMLatsx+eEcDOmN92S/+HDayXLPhDj9YRgAGxDiwW7MAjp3aFQpm6SZfIw2CYz
Q5pNsjj2mg3s38Pz8H7gZ/yahMrKcS8Gx8or3TxYNnOJ3VSkgNWK1S04sVVKETXj4kaKzgCUScWk
j2kmngAQjL+qyBjR2+IS6bnM4pgDixRZ0N3oCQ7awlwR6KIS9AaY4kU9VrWxAi6whRCNhIAiRRKf
mMsO6pIbkmrUaCDNfQI1olzFM+NR3sj67kMVB/5C2+4lGILCSt3uu0DmC+D2gbR5LE2UDiqa5usN
nie7sodsNLU0v5/KiPrwJlf0DjiXpiCBX4nLzeF8hDC20CoAAyQKwkEB1dIjGk1VDfNQaik0Pwk3
ZFGDr7WWxg9thcwDhq8I5RxOKXFTSGkibHW2fQdAQ15J7SxfDPLPQgzECPvu7IL2ATo+DCzlGHfZ
kvU2wfs8j8bryXYngU4oBIren1MgNkXJCLRviTtnNdTAP2dF1hRd+8YN0lO8PcwbkLJD4SfIbZw8
V8ZRG29agewi+kBOk6Pzh9IzT4ryvqdylfZH5u11MHkQ2VrY4El0D6MB1EbyXQRdTxHiLivxAlJY
0065Qu8ThBWifFaaFaJf+ZAz+T3V97hRdjLc5e+FY/RFzvVvd+pxU7ylnodR4e7G1MmsLORq8ysl
t+Q83maJ5UiPYAfl/hVjrDPwX7aKm8aioCseDt+EwRoMsUgqADdrkNLMU778cyQULtcWrzSyuODa
QUT8CG+EJPzozPoJbLm79q7Lj8x2ve8H/y1zgNpficaesRwlwgk1Cdxsj0XX/03yqDvjo60LeCkh
LwOKLUmh+jMuI2ZeYyl+/UVL35ZPaB3Ld3skGY7pI7Z5g7Hi0onTG5+B1/rD4km5ZlWJHVNmr6xm
ORaJFLoZE6/8G8ybZQ+QPCNZoISbeLZie15MsJ48p5KlKEUpmo0SEL7Oj2Bf0zrdKNufBxxkY2/I
WNUcVAuW0wp+3wBNKaCpxBQLZZyILqZ22uqjLlXW4LXJqiFtDRCt/ucgrDcFbUyhhSVCIQGSxu3r
QrB58/w9mTKvfFXM/DhUsC/GXbAw8NNc1lHNewuq+Fk6xoKvU7Wr56MRBDcUQiTe1LEIFZI2B1wW
0o09kxjG3QiaybqVgmiBro8q93Dnp8Ikfcxts0MKlP0tWQaCkS6gbrFcxGyHj4yLdUG6TaE2bzS0
nG8bW8mACwttX8nH/A0ikTnjdzGQFHy0bd5A6WR/75ELNDhezI6sRm4Cr3ynEd3FdPVHguDCA0gt
lFd5nO0PGJLLa9Nw1PHR85V4E4qTet9Li/wMh9rfbhU2kxM0a378BxdtDHS8OJZAHkZVnt5eNVXX
P/6QN4FxUsTQWFrLuFlp9sasoB845ULYq/gE1eT9GnbpZDx0x5t8ENi2Uqd1mGvZ+klZvsH2ElUR
IbV7YmNM0Jvw+Mo4cwrh/jcG0qabNI3OmA8stL6synTz0McgrT/bTqP80SpwNAUaumHHnns32ACu
UjEQQxk7BQWTPmaGQsMqpkenkTEmj71zPCvcSWrPgQ3V2kFFJ/QPPeTZzfx8mHiXraV+2b69wmXR
fgRi02OMo8RqSvMceaEkOZSPO96vVhCsyH1ZI4nH0LEIJ2RukC01TBbbydPalAM0vXq7r9LJ/2hI
zAk08ppVIfpj4ucIgGbkrttt/6swB0UKekXpQqCip7tnlIJns+CYrJNdDJ0hscHbTEkPu+jh1qBC
hWMXjaRUxWuCL0I6Rk+p523uML/iOtsGeCO3ChBmlkf39fQ8JsCRTRObmk0GLGeDNjGJPA1g5kTU
+8wUip41PHadludbNmuH6zDmdo+dCpqj7wcGThgLcFjxSakJB4lgFK7pLONkG12pHxblQi3H7o7J
23K/5K8HRNH72wIaFfe+IUa0eQNXJ2oLXnXidJ9KUy8C4b+ZZGBiTz3Ds1awl8KnHOhBxW/2we8x
zYdo27EQvjAH2818GNl8Ubo41fdU0aGBdSuhKIVuVDRUZyWVQCqw2JvHK2fuJgYidTLKv7MuT2Yr
AohUAgKRd0puWVCCoq6kPjVtVYoN7lrSEtEPU4t76fWmHHG28EevoKcjPJvNOnl89YCbxv2sjYli
0KEph8teXi/yzOvJj/0Mr9niq1bB+07QZXOCy/ESoSwRVPEzFeyPKSPIjRl32q0NshxB0ffOB2IH
c0CzvrMGQrF8YJsYYZZh+o9tIGOc7CYifCbWTBBeCrVwa01C82lxzjdQXAOWyBgu+Bb3D9uyNAM2
The89YXlN2gX73h6dcNz6d5InmwXGNmtR32FRTzMNwPGMP7JfHDvnk5SxcChmwtyeUUaFP0CHlZG
N41EaiFbIJiciaUSrbLKzv0+F2vp3+/kg7HLPklLDSNZ+CaiO5IH5yVN0O0ZmRuiJFAfJn/0Vu+N
gZ56vRW/Y4WneOiAtT06R2tEItgzoBljj//xntAO6yKce8pvWwtxqrJ6njmrpFamVNLbNsZHIPN9
Z2M7XVAH2az2nYSx/uSBc4TLmIIyYrkGAePHKxvKAfST0alOjV/qqtRnQSjy8B1nrU4pl8o/wLFK
zaLr0FPxSgYe7DEIbyYUUOKEvrSF3sILJ8WovDxev6whK2hD3SpOl1sPYJjvFYHO9t/FftLLNsyO
6hmMyLFuMBL2eFvOuM62O9f1tzbpOYcqSHnsC1gZDh8ve4TBwml/V1mUlhrgSxZW/oI2q4C84XLT
wA8K/FAdDhia9mMPh1wLyssaJ3Pd3IvTESp2RtH38wUe3nwHrB+0/iljzf206lB1woZ4Iz53jCTJ
eX9I+ysieaBNwM/bJaiUkDeRwBhAbbsJVHYtxHUXBnPbiCq1tpNZvi13JmDkM0/v89nTC6D4yhBU
Zih27YV1qCz0S1Po0rv0Ot9LRWGWdCyHeQUzTAa5z7ZbYTKaxHfE0UAKMoA2vZa/c+McXV2SVJPz
etVYN2Kj/K/FSADkqXSe18IIZNmO3YYyFeXb/vbhcjM+/2fQ1+gL1yhEa8q04UwDpkoeUV0jZ0gY
EJ/a35h4z4DwDRCD7gwWnH81Jgaqga58vJ9QnS62ST9oI5C6CT+EZKQpuPUcHRfq3n12aEgn8qxC
SaKzAhqRnxLdRJsLEnGzKzEJqIHXJT9W325NPOSLfWEUkrNv2vYOgZPepjcb7QcLZ2BnN9k6TEZG
WjYWcWes2EgBCOuTiUZJfg/gBxd9l5AAfSxuhMb+Qw4dlTeogZLoiz/AX4AMJ3DweysPGyA/oU9Z
GYHuzUD6KKfeGnkSYBqmPUVD4/8+LmC0CqNyldSr7y3sG1DL7JLRLO7Yo3tEwTZeMxTjDh/NiSN1
fR1Lytu61X7bRHxe9YgdpJM98ZjSnkdz/+cbFc8NjaBfHk20OzeTnyv/LIZSJDCGG0UehXayOfrq
hhv/mPHoR7W+gi0fnfgeN0zeWoMVWayl8x8lrfy/eEE+qk+naKvoSbQMz4hJiCE7KPWloWYe/n6u
K+9pZZBQumdJpDAErY3sacM15m7NvOmLhacbPjkSblToErOerm1fAedP4ILWW92wjXb81inyon3L
ZwAgN7N1x3ZgHpG4K2xbziWqNl/8Wtva/DlHgV5DtXCPWDBdls6tyip1zZt+7Ikzp2aKoGjCQ675
dgM9jR8Kjm9WzMuEStAxy4MLJ7kcbjVyqzHBttRHEWwLSVR6c6rt+p6fZQOxYB+YuLosTHpOZPA/
0oTScdOx16Ax8QdPV6sHws/7jZ9SytyMnr3G8svHvnQCiPXqYFhVlxGATy3/jLgb6YtfJ+YWI4mY
+viFYJa8AbNrqTe0WK9ak3T2f4RIj1I14gFV8vqp3r1FzPtg7TBgGGO1fuBmJDVB1VqnuG70Q13N
+6yag7XAqt2TlL0k6SYMbSXxtbRyccyjgUgwUrYTrgHOri/Hfyr7IjrGgLPcl7tWb/kTge/HE+9C
RNAg0J2tMxjpboNzfOfRdOcOL/ckyOeW/CZCmlUUuuZcacLe7XecKrhfdFfmFatd1gJSNJ1SkDo4
g1V8tr/YgaQlBrte1phKjtkPPJPkHwCBziaxOtJrNE8jtpPkKKWNIBVfngvCLTgjtXyDY76SoOcW
mB0LApdglZVDmAN5LXWyslJdQV35E1rH0JilTCtECM32Jca4/EbWplVnSNQxJRAWU8tcSGgLtYx6
Eo2yLhDWHy2BoMR85xw7R00omiNJvSnd0YAvdg5HISTl/iTEfd3xvoabnlkRsb5/tPxd3LAbaAk8
Y9kZHtfY8gOZsex4mdJSckwIA2aFYtduVhpXE8uL6ZX9ie5r+lpXw4YIWLIxvgkraMB42vCtLFAR
SaJKCCA0cA1NNsbCs29p5dZAjkeJ4VDBHxPz29rg7zjFAWTx/Ol1xVFbEqv2db0zD9NcoOrdU10Z
xaXji0hT0yHEG3HD6mGnTQfdvYAbQb56GDd4115ZKBNHYQAW0TohZwl9MTTyLw5kguybZmuvX6U4
UdizVu+Z9GJ6DTerN0C8UQLhJqUacq4b4aooeV31zLIwnm8Rqd8mxuZ7Hu1zlz4ftxL0sjsZbjeB
LthjNlpfRrBJhvoS+q40+ybt7eFEDDQzXV9JG1ThkVJrLssOh6kqS9goSfZXsvY14mWnsXJkXo8d
sJR3N/fDKD2Zk7DYL3FGio85Sk8JCqE7NhpquM2p6FJn7z2NeXejUoYI1pa4s8FoXG6ruqnKwYKZ
wQPnEXDmMetHH7Vl9TNw/kWLgwsBSE2y2k2YYFPYfrF2RmBO4faubrsbHKdfDdFquVF5FJGfIZ6Z
02VPJy8M5SWO+Vn832L6aPxBTefZ6n7tHKcX2wUgL6O6QwRVX9SJPlN5L6TAQLrsHGqpmCnzDQG+
hxObDh80oh6GujW8ZBqWESet/Z4RRYOqyoHfuYDP/FtcT/7R085QXyyKLHAyf8dcK1rCipqx92sN
JLycSbQHknkKLO6G3dhuHnAA+pQ5OsBlSk5SZJylPjUzdeXM8FC1F2znzXYD15L7/8ywoZ7e+tyv
yKLQJlgDCLJaCNcMUDWXdoVugST0vbLbLNdAd6fWjZKmbpJgcI1yy1r59HTjc6ffggNx57oGPAJx
GN8CMQ2vO4QRl59vNlAODc9HZvZ3dy5lfQ0prmeupe31XsvJo3evt/ZLgUBDO8G4sTmuJL4UZHat
gxUuXs+2PHvkWwKWXp5eJloHXz8445NGoqDup553iWTJyM2oKQCult3AJ2UWbijWOJYAW7NeCwrS
5xFPiUQvImu3ZSrLUeSPgRK6Qw64vXOhUKTxC7VI2W7vZKPqyYFAk1E9VeXRmSVQFH5Bl334kDik
hzJOUqsrXqh4SAojIb0UBhIS+G8gcBFmhV5Mf99KfWfXyPvoh9PXz5KEf9AYHh48C6FEt25pIX0R
T4ZNxfttG7sCs3Nk7DInRF45w1lh5kk8TKR4HEuGKNZZYP0AeHTG7gkBprFTkwYa223b2hhw5Iaf
BO03YnK5GJ9Oba/zn7IUkC8fbcwDoqBS/wP7mN6dS8ehMd/na9MWHjJM/chHcGWL0OogHaRUHabK
NQApDBdiPH9LxzsRvs2iWNETgcvDovkwD9D4RCVnqqiscAukq3RNrvOG0h12KvZmYReh6Cevrufk
1WO4wuHMIygiCnLphLexL/R/xMwdIedkuKwU17E7mPWbRTmLXJHPpm2kvmTWLe3IXDFsGYCEjNgu
RNs+z7hpSwitjfRXn+V9xEvLbfPKaDH5eN2ZghiyL+La/taOy0zaWfeWTRlFV247+WA1iTU6IDlz
xffygDX+rG5DY13oI3AWiMkEAF5Wxxe4NdDKwBxlyE6pxS/qpdAes4H1Gk6ql5wbg6WTv9cAebnb
oUMYwQKyOqagJPoL47ElAZnv23mbXkw6Jz2zA/TqGxliy75h6m5hlqbQt/29aT4XoUzX2goTgybD
273LWITCS480u08GBXFPsbtSGzSa9pF6rZxswUsCiNnMTwYrw+ZF7TImSfluIGf9rUWpIjP9FbwL
i1H900wU5Qzeu9mDutylmEgYSv/T9ZIfKqIwfk9VC2NtDpnzmGoWWDkXQwBS5byQchhVIE0Fsl04
nY9QjMznY402hfEJ+dy6EtzCAZU/mJ7bWcHjj1Ofbyi49LADs2tzcVqlYGgQjHxSBTbjEyNQ3JSm
ldbAa9UbwOronlv4OrWSBxMVfjT+kXQnvrRkcPKp37lnHM0qbYJRp1l1hgihzJhCVG3shbljtitV
ePCY/THEuot+bdkhhYZXxqTN63WqPLjZ0X+4XvnZsF95vtuqzQmA1LTezMwnIz0ATyVc46XbgnMP
29OJXDz0IKIbN5QWeUIUAW/9NuVqoQAFuJl/3pXwAG9ubvqaKR+9ViYfxvKQfBJOgJqgEVlwbOBI
ws36AH9tVppuP4uImmc4aXg4926PX6FKZpx6s9Jz0SzdN/GllHMoZr6zoq/6GZO48kmdj4fyfSyP
X0vBhYQwKVMzFFBXQBeDyju9MkMMP47bFCw/CGD3AuUPGvjnao03x3pc3rFUzsoYQWZGuiUML/0s
7npdnJ1qVGPNUR4/IB3C1BNw/N9VGhFlojumviPRvgawO4qv3tqxlaJ8wrP6IViSwiSgM3CvkxL0
M21iQnZIEzqt0vm9XYnGB+yxYnpL/80aClPMLs/siTYb5Hn91z9bIhVK3aG3DkeJPYUQzBtC2Hql
/hn5qpfrSiaVy3/kxOKZ8Gc8f5tzlvJPQ3jFNWiod7OtfwC+J58Bsg4x1nAjXUDIbjKs9O4lOG1E
o9//81U+bJ8WG2odX4jyI3Ps/MEpiTqkCdFBVFV82cDy+fZtcfUmraHO8mK330pYsIYXUQKSbz7g
WSI5ELZQy4OA1pNcwt55S7Ow1mPN0W9IXbnQBs8Iq1a6nLtt53L3BFNEPcnD6oLzlvzpcgj+8fgV
CznobhB2QbTmr2MBdXtelMcYaqxo2HVj6sfizxUXXj5qqbokK1a6eDsHVmSGW+VIT9wYNRkL4/HC
WLot+D2DMMAtiMbLSDXavTe3VWWG4ZLKiI86SRw3QdzN0Z6bhEc4A/2YNSA+oEVfcKLpY9Rtm0EN
jTPombrr9CEkwLBS198weuqaNM5w25wqB71KbhJDHERx/qDxf/M4AZbDjIGtCis/Kpgr8Vuf+cWe
nPkv41IilgGbPNGVIZo2ug3zqMAxT6xkdE4mpIVkDTrcHYs4UoeqHrTNXioR0HocdNmY+n+ZLT3J
QSlAtTMRZn7aYWyJJNPShiAmIWleV+vT0N6OEzdk+W3WTjs6gArob75qlK62FLy3pydKCuZsFa2B
1mm1r095URYQ/EH8tOaI2/pFVXCGltVe0NpQkBjaZvOx2KcEl25SgBeZbDZK+CVnGIbOwVBT+N2M
4n2PqiJ2kjSxHwQM5GLwnPWJ/cCom0nzI/dcP5wY51RUP2wjVH24ZIEtetYiE/EDxDPE+rSgHjhk
QWvWnic9XuB9g44Q0PzFeT0VGt/a0ODzEWaW8susD12Sw+FaIRgpZDUQRySiDE05iH5LHZ5szr9G
3bpDqfp2tNFTOIXUjNdhd4hzh9Wi2ZUWUYW70JDU3RCY/f/7VTkHot96k9qph2ympt707DmsNbJ7
apfcWzSRFdVTtictsvZnBWIaeNfz8eT1hnBrgwzZF6cSoyDJRjn5svTbFP0xfPAGoOD3DXI9blB2
y0JnlS7RBIyQGwlArbHI0kNc/LEfjLc13mjCJ2kOQfMtzFObawEKrOU1e1bjke3t0Q7atg/5VD4R
SYv8V2qa8auekGlNSiEvfFDzgoCDCU+UPs7prGLNaA05qv2janb/qd5c78a5+pr4/hMfdm1x7CU0
UcdgKRsgsfGy5TAqGfJhhUeLXVZsBUJP99TUJNo+uuJ44IEgizBpSLJ5uk7+55LXbhsepAEzKXF2
q5PBmoGEffxDWqeHHmZCMa1SlMVj6fF+Ia11fmRltLuacgUaZBTbKEGvVePzss2ca4gou6r5m5xm
9z+0fIuolySjPwDINB0P/ZocZdRBJO2P0MiqYm91w9LioBqkz18e5rkvnCKrKa6R7A1GVdkHeght
xuc8ABVzdjFG4ZRpGUl1BP20EFMQCo7yg7xi6Y5FFqTEnkJEjbi7qWCOl7WYaej+YgtyH7JtFhJg
5LtLfBVfxdgYYNLx1mLdKfWxAXyLPNJy8GM4wrYXFisgzEHnmS4PpadNhZfMGSku6nnhzJIfd7aS
6PyE5TjlIaNgDzGpiWMAu+p9j2x+K1LZmudouIGOJCLDfV1F7uqBkzZJ7faKh11iO841EIGeZkI3
BRL7R2nWyXGLPrUvvhNFmwrw8OsiwUtU8i+SrnkBjv9f0j+USNZf0eU/Vu45Nu9nNz+uKs61OuCw
hYw5hgAijXXpL0mkLzL4DYAYxGcWQyAZvSnahbtq0cEsNAGi7RoJF5H37s4Y53rqSeT4BtLwiBQj
wj7Z2EYcQNVv6VM80Ndt/Lea9BYcu3ZCnLRrivS22qZMeqgFISTQL9fywPwYxDUD4Es9yi8fIJji
O4jlaJaNkYskbM8XMCyPJFIASNrUjVeWrjq5VYEX0hEiIFc3zs77hO/V4XlGmQ7+/vx0PGSUtbgN
gMKdj5s1F5+zxnXkOc7l3RG1JTQADWu+pJaxAs+zVYIDc7ylqa9rmZbfQK+sw37f5UdEa0Rj00TA
mNxeJmsC7VdrooUvJ+ssSm6iCkfgL5x3+iSzfElvt2YtzRxOLyohKfJ5rDfKHphXHh1sOrVSzhTA
lw6bKVtyUV09ECSClgy042GHp5zcxb1nTDjbcTnp/KHFkiEHyvgFtRTJVSqyBTWWCeCnqOOF6Z9m
GXFo1ssSyp1Zsz6qOfYptVSxxv6Txm77C5xDqVAxKHBw4S8P+W+OI7FkCBCjelWRbwiNix+ohBjK
79TfZLk6tY6+5COBRsa46r6+GCUs1Mrg9l/7wtdVtJ0Irdg6RBnEdWe6n8S2JPEfRZCiNoK0y+ml
RAFHSicVk+JJvR//OtFWVoCdbv4bqCkULg++Bt09FTG7O7Fp6lUAdC6kpGp4azTVyDSAMXpaYIVd
s4bfJCEHGU/fmxp1z5WkEAk9RSTugwm9+d+dGwEP3qMdorwc81yvHtNaNOGmam2gsxzltKBnU42o
ZG7H+VnoiQ2i9q9tsVMEf85EG7Aa+lVc+7QQ7OkC2ae0bNn+tpNoeCdCPJIJIEvjsCcCSahDhRhV
NO1Gv2L/rFtqBT/U08jf1J5vqSVohzsMsY1A5LAhK8YciCdo7sXJ26cLXH+vhu7hRPtnhmyAcolN
wFxwfS279O+/aY5EN59Mjw9AgFsk1/g45LBAaV1drNaJiveGghRCR+0Ug4vD3b7q1p8L+6N1qoFO
IfsyxOKaUVQ5ICAVVhhd1GDPXKCxG52ELE9bQnqNo20rwWURJ09zTmfx3mDGdRdB6CL73yXz+NXO
YyxJufkMYS12CWwaZ5oZcHfFURLBSSfynqQgn70TxSvq/o7hu3BvgHhTgsIv8BDVlTkSt7EwYjjY
sO59OcmhQLk1r+Ca8Rk/wi9ajmoK00ZssJhLWTvyIKlPBL1n6bvZOkZRleUX4M4U+EcOGE3Ks2fQ
UUT9qiu9zTkjVrOEgJFcbRdctAR/6esOpEeAngJC/zxGWGxqtGVLII5LCx8QP+01eO0pBWnck5gE
v2EN8wRm73afiS8Gen52L73717V1Xly6fcUfo6DqEUq96AnNe0HRgkY5bc8S7y1xLCBo9kaOgGRy
wg8gMZsor6bU0RMARfsdHtTRfZvdsMlOVh/DftziKisYGBArVsLvi+6IDwiQiwggEJK3YRntw/ju
/rBNESIdvGw2pq5AtXh5PgLGtBgsbep/l8Lo70+vgIn6yPHs6I571JlimrUvLSbFfc+/M0BZ4Gcv
RutA/8oJD9VuFbyAAIeBIKUuHCvPVShxAatAmUJr3UONPii3qZFjO7EBnTwK+mtBKLvOwCqQGIjs
wFTEuv3xB/AXDWNR07j87/oxpmtqyAO6jyFIQFCfPEP35SW70fZQ/l2yHm6JE/W2s0tN2SOtebyM
2t7+Os9Qn0fcfy4Rw8ONKY1SiYK2BNtPTisi6IEe9nBDfqgKAWdAe0JmZ8BBobB3aJkkA29incU+
5uadBcnYmaX2wTJEF0KknCyM0lnKrdBIj/rTRNcledAfGQmsSL55on9jE1r/NWZKIvMK2mucmO1Z
uU7DU3baOvGXReHOW+j4pJCsSRFNSF3tnqwS95upzsisctgz25Bnln/33YVy0G0qLCwUwha3lkhL
bdhtw7+PzApfb/gLMxkR48hB1TZG0Vy2IO7FDPANsVg00Ehk5avSICgmD1WzhWcpx/OEIJsWmzYR
b1neD69l2c53jfVc98tF0QKbp9g8K2rgXDBW3kbDeCj2vQtp4u/0o8KJ/IRSJ2ehjzd+iEe6U8YS
055Gz5bkXiCFjR4gK4I5ijMF5tgfTVzCwjqIN8bTb6OSgZyJKuqdbxm7eM82kJijUnzm2zC8hez1
2oCRckRD43baI4tqeqoox8uLpDW4hDJcR4pGD1Evjp9BdV/oT3UrPgan2/rP3oFYdmvDBcPK4Iyt
/0USGd4m81WbXv7YQeQm7YLxF0YMvErEazj7n+bQvN9iuR3g8GlCFVVrmejw+ia0VCbM1hFSPEPE
PkRNBdJeQlH3ihusA0KWhcofynRvpdj8NxL3dYi6IikAwaNyg0FHDaoQEbJ5K/U+M9l3tBjIcqdE
kmAw36iJQXVTLoxpmv7ZYlF+82DTjS/laracTi6Izb4CL0M/hoZlG0UxRwn4f7aBCgTK3Znd1Nbp
JeuAJ8pRNr8YjZ8RaBxU69i5Viof2+9HgB34g/oFghxvHQlu5xLAvxMyBpCxotK/5ULqMVqlZJZX
nwIwY5mKQgEPBt2mr14x1eeB6XG6HJMoi+5wvmhBfUY0wmMtcDzI3xLRglTrTFSJ5USa8ld/Ksw5
JL27S+TttvjFKIR1kBHnK9GemMtqUU6cwFK1xz+NSjSeJ3sui4BpUBX/sxOJAAa3IQYpmfB2jGm9
DcWd5ZXV4sjBc+ZpaQ291DwS6EVkFysDos/jiWhOli7HFhhcOlWK23ASEkPR6kFp7KyjfnJkEC4X
M0ej3M/LQnwZHDTeJORVp/u3E56ZbuMXG8AH+dCm/zCdgE1kgQx3FlM4j7i1Yc0EkTl+fsVjLFFL
CIWn/dJn+s103W4OHC5hN3A6HPXA+gb2/2ytP++gnBPAKZOQvPDow9duC4Lrgt0yAcaR3e6oJIw5
p5fBiZ4Y3ZGCP+V0QM8SL6j5QeKU2P2omSPOLdm9V18GdvxNdcesW4VIhFeYInq4M3VGhcRWhCsv
v9CKmkTuI+V4sGSofffa4dLipHd116qgyqD0HYYVxhFrJk4GWB2ijOyEox2aADOnhf6G2LIcLdTr
aqmDc5nQKVB+qn69oAk1DNwVzxc7JTZAiyK4BS3vcXKEZqJa+e0ycvPk+oxBzKXLGkl/fGFbjrEx
vZw5YBeYK7Z2k//4rbbqdMDr0W9oxK52WFpL096vd6Q/OvCUGNJ4APm2lP+9xVYH9np5DEVrrcLf
eK+2FEaqg5VGLQoos3Kjk9uV+VL6u/hjVXhurTLerMQlKK9TbBPnOnCmaeANeuMOTKlQciiewiRQ
+5yQQViYvKrwpLEB2KLsCW5NB/EC8S6ddkAzNUUrEaDRsVcpwCpcblzjui8WyA9D7lhlzqVL++j1
tVndArB2AKWRIavMWZgoeW+i6a1JYDQZ5SMMGqcw4xCH5N0b3p9AymPXlHoWsgjzM1g6Vmlqymr+
P4OCO8GCeI/IaIbubYpG5xL3DDf5v25/xYioPGjFmmoKFfacNG1qkB06AesCAm64inWLiygCOLbU
ODo79oKI93+lPKVP3krnl2DNpqxECRb/VM9D9R/fn4WGO9Uinf1zWutBwvvaAEqLW+nxFFZKLYuf
tq985DoTjN4wjoxl5ynpO3Q+qBpnzgUlZLBRpIF18XF5diaTalHgGx8uqbDD/uvAkIk5vd4VdD7l
gulrorEsiCGjBM/doynx8Mn+fsKl7GTU7u3//yVJbI2j6ybgUdZQANm0JsbRdUkr7aGQqjkgYGuh
9svttg1rIdZAS17XypX4hz4S8QO19aTgUxjiGhXj9E5TaFXzx3Tm4YwZYXl55JP05S5XVo0GDuCi
Vsbod1pm3qHy8onHUs+WcZ9VOkvCSIF5Q/e7ECqhJgc2bVV57qM8jOxJ3DkVN9qGXKLW3UFwPm/x
KlYJQChrAau33F0es47dw43zi6wZHdfflNO1Zc3FDtRAV0a/UQWWF8+KGBOwoaF2Jw3Q9y+h9Uqf
ZiWg57g5FXSdYw+AyUMwpYDICdVWh60lsGwyjjESCFYEUuhwT6DzrttF/KCt4zfI3swlbb640j/w
4O+FQbPGmfNPDHnu2J3iUNwG5bUTHEgRO1GeLtqJsADHW7H144WF7h4p5UTeIGZG+P/pW2eve93F
Ys5n3ZvEGhWAIPIO5FOxm75eG2Q1qa6IygG9ANHom2Su6xiKklsl/DkUOPurvEENEqfnVMA5s5Bn
QCvTVtrCrngAm9HK3LYZh+vun97N8ogYWFrXQHT2uSnj/l/S+L61RsLDmilDgBwXD9kowMmFGdGf
ynSLH47ftxv2xqpJaOZ2PR1xv8qNhnpDXRz0s9TWhEehu3yXeUZwUqZavZio+UgBTZ8162zoPfFE
gyu01un5IFsklMluaOUv1sUxMPLc6uQih3M838pHcAFCCaHGXBxe6WGaso/oEvOiv9qhST/67EPP
firLvfWsOpWzYnGXdok6BEGWeeu5mxx7Caz6v9igtqymaYO1jWxhnggSYcE+gZj4bMM/3zBImq0s
U37tF4ujXUV1J8WySwgV5AMTXZABlFjUikBdesYW0dWFkrtfLs/rNO/ttIEUus4p33usnDVo7CUb
b/zH82zIAnYnpUw0jU9A+V6+kLleLDJt23HbqEgpMNP/w3keyqQYwdXAvQNJ+O2+5IpA53AaCki2
12tQsbjAlK1BC4m6pXB/QgvWodHvL60OyH7ku55lguRmMzvpqScsr/EZC/VRfdbdLvz6DtOAsRce
mwE6ZMN5rNyQtQWKtkV1dkLzRpxwJiUjYr+QFuLGExNUviQjtjUroyrFsBCgILbw1z90z/6qKPnk
oB/PXehFKG33GLejLOiDxbJnPUCwzFYfdtSUPZJU+HJLNECSYKd7zgoDYb56k9myYldOp0FlGiR+
RGd3kDuLmiUb8uRkORNl0j/w2ozZdVDpCZAJHhLusII8mEvYtySb4KzJWoFfJNroY9X4vhjIjuRo
HHxI7aH/4bdHw+Vu3mLjaSVb3aCvNebJkCg3o6kRJa+yU4d2X3i1o5V24R4MDRD9Yr49U8lY6dmT
L9Yp2kIhEOqXnOsm26Qrj+bsIozzXrqrqLcxPTHFQ1iQoKuL78C5ykXljhNS0D+1H1gU3TH2kgH0
YPCh679oyT/YsDNNN70xA3RtcgoGR2ZC+3t/2/0GtplOTJygZ3tP55KG0ALu9hVnZZNqhR6lbUaI
9/V+RgwrzRhoKWZet9LFsqagVvNHCcUE+33FeX4CeDA0C0szf1+d6gxmkIPDvES1AENzf9Z4aklE
ukM1xdOEyd/Cc4jegdtP14MlJDxxyx/xwstIaKUfkALOna5Jxoa5KsL0rIF6+SImJsCMF5oCd7gW
UvZk3aTKmHUYChe9e22RX7f7oVrZK0IhxlVvuB+fDRpZiVeJSoyOkepEddneHsNl2evflbOEO3xb
oPoRHNUf94PqRzk3zdzFTVA0GAnQEsRRVWEN+3TSzLSujKnzZ/kSWp0dmDLsC/0KeGP9mEhBRJyE
grF7A1GvEhKBe7vvjI878X7cAAjX24a/ZoFRkNuRLPInU5BpcTJq422I2kNUm64TxrwD0jYo7vL0
vnQRpxNoI+KpQyL/CAhPT0SLZG17613/uuDgyCayNgA3ho4hmE+5EBRjG3WUhjuaVa8xHfmyMTS1
mMiynv4KEAsmupgN4vk/l+H/H9NIjrPEMeU/LnTQ0ukdVcNKfHu1Me34LklZmaJplNAa1Vlvky69
U+FmTFRSZhA+7FRWE9yDr9VtdnUUKAfPBujWqbwaK041Hle5TdolzSgHTTFPjmd95gfw1x8Eq4la
pmDnrc8YdNcmwiSWPiguAyTsTothwYvwT2410sbnyKd2PT4YXCl8IDktXrVYdfp9mYzvwoWoiZ2m
s40pL7asXAOrwxg9gFOnIoeC+Dc0tllNpCHNk9M6SK9xhI5KDCeMpHMrUwf72btsj7rA5G6tYPPr
Nejg/LCifV5KPQN12TupK43PHU1OZ/QlnT8aL/McDJqgeD2+5JmIn7YMjCJDzaX9aiBfKIagaRR8
OKk9Lv5jtac/E9Yn1nN71gHsdzHnsJMNOxZsDwiDoKPLAZyLNBW7viH4Aa42Kwc+shfV4mhQEWq2
A2r0UlMQ+BE6FU6jY+AMOs4QEi3O7T+vw2bfrIfCJLwwkXPLw2hMH1oXWOQNvH9QhsE1Jzj7P+Gz
T/4zLN0jz+B4oM0awplrbZ+arvdZN/C/lK7hYn92yPStqKYBKXMhZUiou45TjKTFxDkorLvPDKjK
hYq7Zv3Nr9mCmR7TbDHAr1QcSUSwWbTw6w1XTv8SvQNgAT3gpR1kXBZsK6wyGPB4LKmnTRv3JGjV
YH9pRX+4LlmUUH9XNEzp9FNNEPwm+YbqqG8qGC5yNJ2VR9I17ZLhl+MtpkEZu7uATwn3fqzeWN18
7gnEigApjn17SsvzFeHyBHdQoCIp/H6vbAJmN4dpmgpxJfjnbRrKnWhEVfHT+ZU2pCDF8c7eqX9F
HcofquNvhxul9HArEOuYOUU0tqs8q3te2GEzBbrmNUNExOuJ+KILCAtqdvJIFWVLvZChvlrGMUvm
bPlPDw1H07lijt7LStH2ooaonMaeO9rM+dfJNSHlGowEuauFQyb3H+bYgroCKznvpayggyMnlUvs
V1z6/4FF9LeNmGbCZOoKMz13sbBEXs6tDqVluq2GH7VfjHlrUMOSaWzX0amjBzyMgEn+/3PiNT8W
jKAhvNmMaAupU3GfhZJWHvcufu6jY7St9u0nXNtvoYQjYm55ytMc7ALI7eEARnrsvBWV1rqgrAQO
0YJ1224uZ53IVHrA2NU6pUKaa1uWHUHVrNl93xODfb2wc9aGGSObQNNlcCen2PzVkvYsd57JD4Gz
spTzQtyVxnaQ+8OXN1U4yWyLGOkWAHiUoCQG/d0GxBE+2+ixGddSaiGvIPTQ0cQezSUh7GDsgK6A
IThJyAoXLF8WkGzQXyGZP5E3bVGa0zNmlm7X/Rnoi/3XMUc8oxKForN9evl41CSLT5QYry5K0M6o
ciMintSCwwNU3kUGK/0Nvfm1T68G4kcW7iiDBR1XOgbW4zWMc4f0ydg4tGln2hz2jkrFxo14qxbg
lOMN9Ra5HKb9yobLKMXw9ZTC2wxbTnkiTHi2X9rBUf8DvsJ0eoEbMv7bj973xsyBizoh4jJzAJwa
BRY40j+vlJz1CnNAP8cKCS41aMI+yhQ0w6XNvIW+6Jj1R6WWklZz07Z0qMTEm8mASrmPJr1gwqEs
j/pW+rjROlPGpnH+mPqkCfG8gUPh1IuHRgv7MO97EPDmJfD/9irwLGcyDLZQHDhr+oLix/C1MJ8L
DkiHC6pdV2XHbRnZZNPlaiTy84pulmTbDWV625zWMPeRJgDkjDO58+SHjeiPbZAXhGFJBztNKQzD
nXGHzp/elYZU5VT3oxUdbHJ7A/kvGk4TAoHJzzHbRGwidO7+cNIZqFReG2l0EzJ0ajyBzVUX6rS1
XFCxgRihmK6c0JpuN2gWk+1d1c9QI7JDxeippDhGXvpsqJGppmENBhTC5DdBZ5+0tyouWlCMRnaR
h/c/rZw4PCbpELwnTjG0vwiog7Qi0zx+slNz4IJ9pyOj30T9jeDHKVPRNSVRHQiY5b6fwQT8IbIl
AIX+gqaKdZsBDQReCqczmMwG1aGyhhuPJbePvfS2KecYizhkxgunw6aO2FPx81WDpQk61XgI32F3
rwhoob0u3jkixUodxlkWjT/GfJWyt0qSCIwVdm7cHf/eGYjleiyV6fVAIRfV62Binxn3uKuPK5VW
0IETbNmk8wGgCX5oJPsf9y3fJIinIR19V2/NnILrP7xA16nc7N5HdwJlMiayHjYs/Mj8Q2lieyC+
cccdL6pbdh+yuylCvppSB0Jm+YHeFU9IAt/3fxXASx5Zh6gMyh8ETtOpAimAGWMGCTXCS/xRi0h8
b/UAd4F5y24Ca8TZPUoQPZfmJwR6IUIjoxdz79P/amigiLzX4QublI7U3gby//NVt3wSD84dRfwl
543ZW0EpZr7PVUIKAkszEFhTEI45gziydj5MODEq2aBdcqYlRywslwSJUKfK8hKe2S9OrBMIVGvO
E9WnOOOSuX/SYUEP4kF5dHS3nR3FCUOHXk4Fqf7ngTwezDS0n0a4FviKG9uTKML8+UTiNptdJDAB
oSS4fRStHGYss+3GzvZWTardmR4QmYj6/5cxnVLTSQZTaCHtH3EcluK0Oj6RxyX+fMnSGhjeJhoA
arAzaL35Fh+Qn34oSbPdjmm1Gm/UeG/GToag1NZt1y4EBKAlPwR+kweiqVsVRG5kBTCy4GmupexD
pYMO5HeBFgrBe45mywDmLEFN5CWPWcPtF584At0dfvW8Es1ax7UYStsgAbrkoTx4/Tk3P1F8VwVv
79RjzB7wNhe7x0jYo/Us7bbvvAdv7GgZRFM6eWoPMJ1w1t9DvmwH0uhf4quycZdRWAzt9FNwUofu
yzNTsT+akgpyydbJSnlhgQ3gRN7lQnXAqaNOOK7EikSWu4I1aIItsFd8ECevB3buO27eHYocUlcY
WLAXXhCeKL2Kp8+7tJU46VE5UNR4MuPKyjN2px6zsPS28xDPhq9+ti7w+4DUvZ/VQQGATpe70Kll
u4hqhxc9g5pCdBcH2C8DBmXAjrS27OyTX9EHyowPYruMksG1co6Tvayp3sE8y0+TsjL54GMQJXRx
rMjmmB2Pp9uJzEz83zBjMqAvGI00tAtQOj60fNAn5aswp6OuHDivyXnmSUyakPzk80oqloMntQQH
BmpFJarJOo4R7uS05efZ4aA5LoJS7PQ3116ft8U8kv5sd+HyX2/EemoC8DPINb/3okRfL5XM8lFS
uHgwsMosu7rFZz0t/12l2v4uZfS5OnxJEFPzDVQrH8PHNgZs/+3uW7kZdRPemQ0nFUg9xv0S/qHV
zwWrA/m/rgOXRgiMLcWK09jQXLC7Rn6KuDMLT43quQSCWXUGH2Uq5rMLj8N5rFqHZueIRfTGpXHL
6SK2v7E81stYLnIkrQaS/q/k5Lwk1vKdj15cvHYYwAtVNLUTaDQuhkzwPJN+QunstpFcMMhh3sTp
gEwaIxwAJM4e2UNs/Q4CM+UPWngdgdY66PCDchawrqVaWaXilA853nTrU0O87KPyuJkBu3kFvn3X
nPWCfD0eBqbUJz6tunh2fsPZdx98f02dsGSi+/nicPjGtnR6wM7I5P8szcTjmR/zdVX10Mmcyc/N
Zw+mhXrXoNT3fuWhJi26BtS91EQvJjeozmv81Bw2xHSUiCpzxvF9hX9tVnut7z24PiYDxFwBrTnN
tZmbNd/x4GosWDl90cCi42YXTXJg9RXULGipJGYvG9Sc9dLXLLR/zH6CvCsxLGjo+uy9BayRfqsj
qxBzgFNEyykeqqsrZyHD9gDHh8clC2/NhOUP4Hm10iZW4EzRh+iMVzOS9JWrMlQcl9A3mJo1XN+N
LIWm1v8yl9PO/FuDpYkTI63RWTIbQqLeL+N8EU9z0uD93xbuNTqh73Xvr1FHrkb/eORjWcVqNHtu
JWc8kBc8y3HtRK8z2JbSkjOr04fppVfVdZPJZffuf4jrIgiZx4PCZa82mG/tzM05KYa389GdiJHK
UDQLGfYH38EM1NrA8Q4zS5XPN0PfvaZY4VvN9uwL5xcBGoWlds8xGt6bZD29JZGuEaDu9KGaSS6A
yQePqqtGY21SggROe7Ai4o5s76eB4N7dMrDUOMYdEcaEpXg5x5A518dUQzQW3VtkrOe8Pq0a/33S
Jec4xUM2OVkRptUMBZu3+dBpHwRI7lBK/vH6/QM/4hMgD1z7d54C4L/1gYDVjAStEk5hiYuxSoxI
RRivttJS/raeR8+85x4xqQ90sTfRdAAHHun5cA7ozBnKaN7kNtl7vu+i4xSI/MjySrPyn9e1Gbzu
uk7Su+/rrCUJbVg0EcNPbKfM5HPgAEFlucockR0Olm/UdGAHYN8c8Hidk+5XPNw65iFrvgCaEqGx
lAPn7Z5hitZv7viR7xNe1n2mtKlHZB0poFbCn+dRCdlp73IhB/0VpD5y22jNb6NbR53Q8BPW+Lsl
uFUYxM6Rh0fd9D7degSIaitp9RlF6uEpM5y1mfEYavHSQXsK7Jq3lDqFS5LtAuEzlkjGT5G/+58Z
vaoVxnH6JtMghkYP9dWeH68OaF34NgBKkC8GFzqdZ2Bljv+QAqonvLDR+i52BT04o3NgehipYltu
7qdBW13qrqiWmjqz7gpey1SBlwi2Xy8a59pDj8xTVY5ipJrLNm7UVv6VEoEaDuDprVeTcTAaFxxL
T5i+qRTeH4rmvDXoCjPwk2UZH1Wvao17vnyIoI7GkRW1dtMQiqzXJMS/i0PwL9oc6LStoxfROkL+
skZukx6L197KJTfsZllXeonFyTbd29HIbCtuVA/8Yl+t1PoWVieJJxx6sHvdNIa/2qjZpF+Ntd4L
+kTzOdmKHrqtEmv9Jbz2qGRuhNdghobmjsQrqrYUJEq6ZzZVr/Uo3rKWGdXn9keXz+WwZmd/0pJs
j8g3ID/uNGqhQ5Ye2vLUgIB18wXgVmaIU0B9Tb/v8+d4QoGv9mwgvSWvZBiSwFT36Q0YptXGVq/G
Z+JhG9bE4RO676ThvOlvi6Ir8qELwytlQa3nqSHyvGS/CAWbtm0QpyFTdjS4PVb5clcBBjbMWthz
aHTfirW/qoimt/57/OkamA3dtE8vWzfFfNO4Dt/qeR0RCXDwCvqcvWfGTmuefYpus31UlVSjOMbV
2qhD6JyowSsG7w8x8Rgg5Zq8OHSx9WyizY0TrKHNc4jbKs/BMf4n+wtG2cEyEkt8VeqApUh6fHki
ZRkDZD34aaa+kIhW0jJl7eVtbig2m/lWyyewAoHqpyeSssLMN7nZDgBEHowMSihw5gVuqvvn2FFC
/Xlkg/szn8HyVqRryqUbFDqwo4n5EO5rKGxU/ZbTQ2X8babzE5saDl/p4YS93fIsEmNbCMvVS52q
J5hmQ5O0icOJonyeWX8TLWOeFiP7xVno4bVAbR5+NpNaY51/PR1gFpamomQnKk+orOr2664iykuj
QXMuI5mPHVjYhxbzv+vVpektx7iOsy1BtJEUuGFWQRHYIpSFn5fj+uzs4aMcyVdF1yibXvnGEOLB
mi02/YFz+V3k2HUvyofMEf43Ydud/f4DbgTvlOf3dUoVr3kP87M70jJRbhArDdn0jBpc8YvqIG6c
poGHXC5XgcKMyTL29JXoufvW4Ryoc4e5JlWvblqM4pAxJ+ZYheluPTh2B9Z8X6rRohYK0/b3NkFr
ujb8W5i4xiDfGTJTp18Jjwvs0wqNpq9YfHYlBaa6EqydG+S22kF3nlg+rYKejwtM9rXxo5HJaOpW
3lt8uhhkSYFTwA0rUUurEUyMLCiDa0vGasqhEjSDgNPTGUY4w/KykxlAPWVQ+ZyLzUFj6/9n2va1
XZ3AhLTo5X2XAKWFHV0qOj2DGxicZAypyI2E/98gcsoi/NaVUAckKW0hQpib1l8nB5aeyQo2GTks
2gRgZPP33TdPUF4niyArkmfquBbsHqbxSNmAAYrylKCfv9Z486ud5AB7vaJugSdGwE+n7hWzqD1B
EGagIQxhWNTPHCujAHsmZdvswP4f8RXwFfDbcrKFiTWdjGjXrRPuru6ty2rmW38jc4PFu3XZZlzr
DCZq0qlVteC9b0hIbF9G4TdBvhSqV3le5SxvypxN6L2NPj4Vt6kQDweu4eE9yeAgrvqojSxMRex6
jpNSi/vs7GdAj1Lj2+VlnKVWvygFmnHgnCQUUsB98z0hurbU97vaiPtOi3kOV64JTlbAjFQO9LKC
HDEwolMC4Mrx2k5b6lUNMPxxTN5fHszzKPEEfQRFdRhrLDj6MJ9sVQennWK4la2w0vQlOCERCrAd
WkXa/aozS+btOD3iKt6Lmo6rzpGszpiwdj2/zev4WOPo7/Lp284GKzwHf+l1Rv0cGs7JfV6ZiYrN
1JJS7LGktjZjHkqslsnoU6NBpYuecZi2mmoPwlGiG1DyASPwefZq/Hgw49dpFvDg/ZMX9HdgpIWW
16BP6/m8J5P4KWYXLoVIS/cion92P8+kvy2O83swhYUl5nqQRQcDeJaYNamVt3uys/2S2n5SAYH2
DIysv11fSAgQ+yKCt1Dhk0MOyYB3Z517sggn2yZzHiCEUWIw8x5FCcvj5fIa3bGNIdDRVm2Rl0I8
GrarauxsQZc68fBX3NOMftA8BAsDFNPBBsFN+fy9EaelZSHz/e6/zu30OT5R0zvimhDtnzV7bSpZ
bh/vwDyhwHY+r6ADWDBeeS39xFSL6nhim96w9/YMRrkGgr5RXkFrVDsaBMfkIlGiu0u1Y12VskcB
G4nUhN2c83jb2vH6JX/zLssAo13/tU3KVE6vT/8mrqEq0LDsmfwBPk5nyAsmcV9aPCeLxwWV5Ht1
H3ZNRG0NdWm9r6wb5BY0oFUoFoAhXMLxnUY0b5R0A19WT9tApS9e/PcsF02sk2ScvteJnzrFSXZK
LYFZdhbMsiuoy5803k3mlWyzdxy4iXpQzMQbE+XpP5FqAHQZKyoOYwYIPM72VHK/MM0uCWm6XoNT
D5o+a/cd2xeIqFgf3bWLJ86AcIzle5QxUXWkT/mjz/TXkRpSyMTsDH8YuFUQSpIqgN+mOPm6TVy5
mdsTArLrmQCKf5ZxcRfbIBPbgf2PnZ4HBAkA/W0oycCJFXgcZFgLmCKlt3WvB9YtBROwDLvPevcY
E2XM/LC9e5CkzWEJ2/ePtd28Zc/KbONLBEKnkcyhA4tsA+PEOWbqOLLrpiCg4GcbTmp0xytdzvFl
RAa6VgYmf0sXqPSuVocmqvW+sKMI0eBAqD/fnp8kWAxFQotChjmP81tzZPcQAD5VfcNnRy4c61/8
N1OYmHxxuTS9xCTmnqhn96J4OuJEyddzV2JXYFcLp4stzNm+GZfREZVynGPs5qK4AeWlt6divuWP
iFtirifYDe5Kdqo6hlUPwshPGqinEbFEWv/O+iOI3+sxp1C6cFlSMJOGFpU7kKiVLUhFm6nzxxcK
i3gydjcQevyRnHPBn0iapE9iB7YRLIF+2kXogjv3vx9fRsZ0xThGBGXDVy08hHlhhQsZxrWXfWGd
7mOY9uOIgsCgnrZUMc/kO2dSuGIeNcCOosWCnmfREJ6lh7AxA9BNzTD1Oqg60qZqxOq1JLcph5xa
vI2bY9x1CYC57LJ579ixtafqCCtAjl/MCDSCNLVcPdOGCkHbWKsBNfg78FqMca58jZVaU6dIXBjK
8ggP5dJi9VohZIsw5aP3yCS3cpl5pC7Lu1HmBiP+MnBUhe/1bIpsKv5qwZ2Zr2jznqcyK39ITTyr
D9giJqEfLA7XYWcbHS4hQht5rLC4aMWtSQAQnY4KwiiaABW+yTpqIT7lYodHJ+WtTN7cXvW0URM9
xsNEVf/+ISFhW59ZT5MZk6CzKdP1U9/mmQMlejw2dYkRDuYkgc85S2+aBgactMhhOkHazwvD/jdW
7TutlYiV9qfN8r9v8UfMCXzKCtAvSnZGnqH8FZJ5G/jaBBNcZorPPoaubeuK2QYJhbZyU7u/Sfti
oiPR/BIlkUko+OpEtynap6D5+sWnSmSg6NtrcHnLdRxDtIXstJO4VqLJ0P2wAQUbvAU76i+qL5HY
v8HbUHqBDN2en4RkByc3CsSwB8PxaQgSyAI+5ZHnKihcH10BT0+Fyx8V2pdwdSIzxRtsn+L5Hd64
0DgCaLbSxiWhzbcNxw7pg1sJoFA9NSQOERpXw1H3cBAhEBdFI72m8t2YEVlMtcS8LH7rpPIQzkzs
iI1TzWzjCUhHXu0NEBFEzVXXQwn8lQzjrDAhXks5CW1X8TApB5ez6FpytfnzHOnZbk+WrXY6FMQ6
AhFY1kz1SqLhIoOkGFfoKjUsQlvzI2GJGpOzgwx/mnoaWm1vBP5jhWCC/HxRWwzWaK/3B/rKi5uP
gzvJJdvliPECTMjmGzpad8iAOVSCsXY6xxU2XK4zatkRN2dg832atra8SCg/I0rvgw5Rip7z7Lnp
tEu7UBFA7EbCOD1jNWncq2j1hHwtStj2yj7AZuS4mmGhLMO0Epzz4HsKjHceV69bdoCXE8OzGXz9
GigcvE9rGfCdP26A+iY7fDyfxrRLKQIjJoQLBdMPsKXkbNAXGF7K8lo/wBvxcYhoqpVB/vBxVIoh
MMsgSF2a3hWkJLTzbP4QbH5XUGgC6eWzr8eiHWfXBpivI5J7oJ98EY9a4gd3pHuCPQenmSl3fDQa
+OchGU39pHSiZKZ0I1bIlKyF7SQosrpCsLIWhwgFMMVSMZCRQD7+9hdmKmlybgsy+rKUX/u2T4K7
/qJkJoZT1jckIjtKjXFkckCfDgVLvbscFFcJ4TG8looJM3NjTE1rFsftZNoFl3F29Qbls/6GFk6t
x0wBYBs1sxBjzNA5CX5SRy0UmO1LTI2YAyI7vRQh+kou0earVVNfnU6xiFoHyFADuPwbv/So0Ova
rmt1lJnRZpyqNd5JcPgjgcVmsxRQfI6DbV94p6glUWTx1rDEwYOasjWbTVmc+Me5uXqSaaJry6Xt
/+A/q4dfrFtcRIpJF9Q9H/ZekxE160j3aTr+Ol0yjvXPxr3hiBNk4vTDCekXGKp4qucKl+HD50Yk
kzi0YvJE/7H2CiG8bBMiJTTpa8r6tZOHeDpBzvtKmo3CRTSSrU3Ed6xw3Lb8IEVZVDRGQRO2IL8P
mEw0zvtD2iHpLxxgBHa6rtnLHXCBeRe4WUFUwyklzPn1gLR+fl4/ppOxCYtE++6KveqQvreAJfN5
2oLozqr1CLgdhkNgqWg/Q11YOn826ajohqLgX4cuCv2G+7qSG2lQ/VERHat7f+e57UzmodxWrwtr
TC3AWXn5vDYGYzCnEG3AtpT4iLvWTGPkCZMbWcUWaMkzzL23nXVegSRobYTE3wp2FAGYzS46mcED
boMrGhs8tBZe1nCFg4AcWUmKKXFz5wg0lXqTVx4UN0JNGKgo9helEx+ndSODFoEb5L35Ovoda6L6
ZOJ/ZraIKb/hCK/kj2JeP4f56UAS7UJFB8Mbo15Q+3b2S/YmYF6VdPkIb2BQG+DSOa4EDroFg0sF
z7+/cMDusuk1KVnB3fWcx4MxmgTiQXJO5jXjceDxdc8rkIKfdYvrtalInga9D+nnlwlULOetptAD
4vPXidd9np9i5hCqbN6lUB5DFs5vAGSaUCkULTe25SrXYS1rbG4/KveFOPjRtjTjq6UcTvWwC9pA
VHw2Xx29ld8QwFdnDpQkWMBN92YwqdqPsG46cn8EVgdD8TX3vytQuvXkJD/WYqN1/3uUOzImooul
66X5uu3v/Dl2++TEgLS7wovjQHuKyX5WQrZAT8R5h1gSVFtf/k/UJ6GV4IUJDeGZ8V0OKaiKd1VV
Uew7NXGKKMV8gAnvBro1SnGoFDCyvDsmC9InETu2IXnOnjZ5mNhzTl1gYibySU3eTgAY7bVNOX6w
F71Nf9WHSlsZ+7Q3oWb232Xw0rw4oaiwdrtPRyJ794uv3PNb/iUGlTr8hAnDMYLAE/RXg8S+Ldw5
OCIPqK01KcCY1SLJ4u+BW4alL66glgN1tPIOdVJXsa2apN3RO3l1l3AQ5vP4VOJdshMe52ADgY3E
O8IOfPkBpVHZ5X8gVmpiAZN5QYKV5UFszCfyRSLBLSxVds7tPW0CWiSDF+vMhpC4pl0tqp2qzqva
dumczjdkKGpu0Cf1p6w0hmgmQ/fyUmvGhw/wSpBi+dnVqjCgyfSirojw2aVEe9LrsjgX4E3GGxD5
JYgCLXl2YhLmWPrlX6G0AC0ziS6QArGijTqqXoLj0441lNohF+2O43p7R4kwe6ZpjSCOcn9omdLR
0DzBqiyLZd1rFGgcQiyfw0JVuars14XoPxL+k8uL25Aa8avNlRAChTnwZ9q2JhLv131S/aesJpk8
jP7Lj0J6KXi3+fIEQXqjFCfJJcW9Fy84Mor88hdidwkHmQrEux3FIlofGKEtOdML/s2ZKHxTNJeM
MJ8HVwcBP5TGHO6tOD81JoyXpLrUbrE5q5e00YBJA3qmoOWai8Bb8iikPN+oG19TFr3xQfqFpalt
HhsHyqf3E9TuYNXqInh+lKvyYYMPnFk2NiJaHJ/gPrNQLSj/C6aF2S1nSE9FSJUVkb28+D+43Byw
2gIJ7znF53VByskpUGJTAhZlxO85O2yN/RWCJX40lg8Mpx12Wqv1+CwoR+TdRlsocaMfVoMvlysK
KaJ0QAAwL/hdG+VLUuv7064fOTXtzl+hTMN2Vm1N0JIpsjOE6mA/7UoD4NArWO42hOznWQ9OF4sg
zL0uEttavcwHbutpdQFaj3Zr0C7OQzV3MhAVyK4+FAzq3mgAt3pn5BSnoa8Y1z9ZoG6zdf/l5EpG
BPw1eVE+7D88oYN2pQIOjOwOxUFNVzVOc0ZN5VLeZcMEH26qnKww8aoXT7ZAIj6Fp9JpK/IEk4MX
LgHurx5b1tTc3/rlaygimrs6z/6sHxUwWbkea2eVVttr9866BLbOvmSwU8ztN84O2G1P01iNYL/C
yeQEaqg17BphBva3mhi9+EQcpIsYNPnAowp8WJ/8PgEoaSGJayFQguhsFugwceFq28YGQv21tSYo
sGZUKBahrAzT3+EvIu2y/qVLnHKArRFnPFD8c3EFQ/pEqMZCbH8iJOHdSrwj76acrwI5Vy4q2AVT
WR6ylrtUiBOS2S+PLCgo3fRCAjfVAptu3AMepjvyxv6sjrS9efy13bEY5mJGL8szxV6igBFCZBmo
nfEOJr8v9vl3Ov4q4BDFHszjp4emMKmXwKhHqj5+UPLgcy0kfO5HCYUqBRZrJXogz57tZdtDb2Z0
Ln0ObG3egJodIjrkbNztnffU6eG0iPXA8MibktzCNRYBJNcpdD8/x4r7GGaeQRyf2sHEnqc4Yp6P
a+K8a23csFJj8tFAzoVFLJWlDkOZMQluEQ7H9DUU5xMF7NAF8/O/z4OYNw/glZfePKJwCiKvSLFF
vaUSkLJzA4hzurbiO7LkEYCKtnBYokapc7hStgJo4XbIGtZBLbMG5iHtFddj8UkP1INkkirU7h3X
fBj0aCyhg4dASaW8jnSDmaGACGnAPQyyJbuNIll4iNjjnh6M4H5nTmaS8J/m+mr7ouUG1nxawmXf
QF2AtLR00GJHHImV4FU/HFkTPWt/JF1ipmUfLz1WgtDYuQLpQMy3SydhFSrpRzUTNsn0w4EI2l2F
syq4oKgTesq/uD+cj87UrIvUCHTAA+CQQuTsfIBoGsfwdaBrUap8482MsbBPU2pMl6zqO3iMODPa
rqi4dhjr+PcPmEZNYUFvArwWPaASZLRliTti0QVd5L84NMOnTBVxvqU3bLNkq5WkFQrZt421cU0p
j/4YwJQr54fq8D+WUmh4r/bYoUEmTKotIHqwca7JGDi32Cicp5IM3u14w2xSyRAeBiiLtEFMBzgx
vUZ3DIj+SDd/VZ+5v5J+vsXopz7vGt+4V6T046EnrBnCK5Gi0eeShyhU7UNDMpolXJWVDBSpi6Yv
J+us+RiGQH1OqHPqzER1Ww8B2I5+wbBn6FWM/JhXsVfQugI788KVUq6G/K2BrUMPCRbpNWI13uhz
5Z5IqevYp6iK1+K/mWoTYt5A0229fMyom15iYP5h3yBH56+QsrE0ZJyFzBt+gM3FDRUqeDHfNaFO
ULZ+sJyehdQlt+GEv4+Iret6xHoREdNid7xLH/y9QoMqE0HDMJQf3WrwPszy31AkxGrSFEJ/F1Cm
/9/MvAXarHt4wncqNKQ23XrGjSJC+1mgTeC/qX/ER/9/0poBRmeAaV+o6/XYH84J/qz8xZXToXn3
2upM9dPVdJIhC/BDh5ryziGx5vJ0ZhccpIBZjyO2Ky6sF9Qwjo158av9Z+n5zp/01ZCihTbxL2iw
35KOkcoWOd6YrnVmhObT3ldRbNDDK8B8K7pQKG71bx81f+FjQgtm5oRsZP/uUMYc/YsCY344qOVb
sLS9HGqxI2T5diLYcvkvVRl7D0yxVhtpXhyosSR9EtpH5yBFtiWDXegNWrSMazQQ5bWfIQquM4Ho
KWKw34Df1yVfYl+6pFvYdskCKMKlXuaJRiNSvh/cueoKnEWqiMz7NCcMayDNQFHAAVf+GpX0Zjai
pV8raleaY4HTw1M3uIs5H+GbpWKZbvyWdl/7/49WqTmjtfa9x8LE3sQ5HfVD91n7/ASHQ+FVRB8p
tW34AzePfImtHgee+Ydtx80n4ug45nUonqTLSJr4UEQwTTdhileHSa6fgF2N1bSKRsLuI64wBjNS
fKDH+mx3de+U1+GDNH6R+DPbBCqSEaJ8LvBP8yrlCI33MkYLH7xWo/aNrebSHFjVCYRr90XCmQej
BbWfVCnDiBKt0qUrNbkschx1YNfocOBv5QxkrjgvToPfQ2Li8vLu+GUPGIfRRjqV3uYYoMngbD6h
3ZuhP+Y6gvWyqcffZQGzNvoGruHuGEkaLflc/xK+AMaKs05w5HTrt1LgmkOrrypOze16WRNMc3BF
pOskcA7eEZjCHgir/2SVn5uScBH5txPVeoc+hBur0qp5k5Qz2EHIhP6FdgtUO0FW+GtH9erKRzeH
dlUKLXbD3ac67LZ1k7D8YJ7Ae7cb8YENM/Xe31ku4SbEQuF4FZ+4+Gmwl2WNdFO/oqAaIAqVLt6J
7UMnabOxP2oLVny5JoqJikejyT+46Z4X68t/U+9dsMwdU/48dDIowY9DWCFsocshB927fPZmxu3p
R8huK7ZcoPBUnVcJa1Ing/ogFC4uvPfXCoqQQSMR4uexUlaB8cdfopl0GcrW1LheYV6MVLwYP2SY
78OE+sPbLYoly+q/bp9IEvlH0EkOOeb8uGWV0XyyRO7QVVLc0wARPTGgvRjkYJvpqBzC7jDRMA6/
v93LTY8P3Tm+81xTHJ+GpKHVeaHsW+ONd3UlUQ4hRL9y249Zj9+v9Vd9T1hV3DwiAcRMYxzkrLfW
wt4OEIkZgIAgVsdyzFuR+hbSLrm1IrAT8kkN5stRzhCUdfbNX6uTxkjZUwif7k1EkzDy23P0liEE
Wrfp5QVZIw8E1Q0pI92EC//zu6rRwL/8ueS9ot07fQX0JZDmpHJ4VoleeRVYrsUcuL02mKgHiPvg
d4Xa5kWLEzECAEBjz93/gDyz7z+LHDfsT+m+pWPukhJjGyAhcpHudmgmfWAeibtufVBpKcqtTdQN
NP5J6hvdMUm/w3HQi5gAzH5gBf8ymB9zYdD/Eqinh+DofZrJuiV/m+nxs1C5VDGln1m26QF8eoY7
gTAdZ0PaKVsYVziPbWT8GvhGOmjrL0rCxS0uRLCip5c7iQQIQfKxSjmYxqnIPfazjrAujElswhzO
uStndvVOOn1s2QeULHuHRStWT6aC0lzUyctyqChpcw1lP2akYtlqsym71mCZhgBGhTZFiaLv4k0f
oPh2jHw0dqrZ+Ac+Y8KUe2xSYTRSsLyoi9vkOdJF96JnuGc59huKmdRvs7/16iegKTAkkOsQvf/V
U3dfkWoVe5L6Er/Jir91ksOZr7X7oSsAcEv2vllSdzXrnxih86JlYKEDSY7n5RVUmY+ahFKlKGMd
PWdeQRYNrdmgeZPtHkLsm+QYk90wwCvSovr3CGH8oSgMZFL5C1mlmnjCoyuz1eXeSIeERJmNu6b0
0C+eHAtpMwmO28zp95+/m3ZR4TKUBO1uTlTaH4QU07KDbarcIFTxzH5p3jRR/ZY1mk2E5ObjB5Cu
q1TZoraEUpztBaUJWE172suunjwAU0j3yHGvh3oeZoJvK+OtQtTqTCNHYxKIo34//lxF5kHliIDP
Y1vjPWYQOMFv/rBoa7JCzYC04yJItkvjx84+oaALhhsLSKKfLNhYaA4U3D8fPVwnpcZKJ9QoNj+w
hhEZ0vcuKJCoGm6Pxf30iAcfdcqdNorkLKD92omg1gP4Hv7BKB0Xkcod32WHVOixzz2yYoyyf1E4
HN/nU6BM+pKZHWNUP5AtxbO2z3+ipSPieENFslNYZURcDmoL925qykx5zTRcZq8zb7hZWtdX+zvw
CE0gLhGHFk3cy/dTwBzlzsDI/D99z3BUHMm9w3rUlVX2v7ohHCOAqN3ipfFkZ8bDgc3jFuLgebkA
RP5NVaq62tUPMDL1nLcmhhBorBHYUMSAniEuQ85Uhd1R1n/N1yzIAu5NgXLQi3+aimamaKln/4vQ
pZ7MANEoeup78zg0687Bo62JKW4H8SL46y4smc+kV2pHPLjNdaiYuTfXZoF/Rd1jsokvJmBv/U0K
ycJpTh6NZUu5qrujCzgrKt+CcWgENHpwH4HvjQ6hthcPnG8t3eApm3vXHwX1B370NqLur4bdnnd6
c+lBMtzBHQIUu5hgGKzcDNFCdmzzRlccZUSkRBlyGNz/Fs98sV/VLClHWzTO3ks8/nwOvfBjum/D
+BtFLZ4DY30aKaU04tvrNUAmO3JtapO+P5NEf4JurdLNE8kIHBHxx40ocz6VwT4Db4PDWWdsOW/9
IBLJn8fvNc4OHGgEmMN6KfO6LX8/AsVyyELJoiScSnHRWxbFCcOcRqISgJkeVCTQiC4MUtZ80UOG
LDWhIJgbvXEFLcJ4YFrdi8JZjVtYSaKt3Z/FfP9cRkv/M9Bv0mMhztuMd05pksUcE/Up2upnIxAz
LpYeNpJdmd6dLIeBHPXS3j4WeU5H1v+dFXBi2E1/k6xGEO4PiMTPBOhDt0WyLKJ/iebIxhxgDl3G
dqYrjb1FDmvrlWD4C9ZBP3UyBWZWbj+v1UgzMRBbCotA2UoK3sFRWsBYiNqiVBx41aA56YMZZuGK
kGnlud54RrSZFixI47f8oxeXkHlTBEFHWGmSenu7bq1ulOIoaz4wgaOQyGR92a00+coLVqWiYPXD
gj1YBSIbFeDJegYfYi5xR9G9qo5kgVQkUBQVWVOicsWzVUN0EXJt4HYqjUOrvNSCNKGDcY25h/Xh
xHVnAKu82c6UhvoIv/H9zTW3zrAeDyRZuE1jxMXym99q4aDWe9TTqBYWB3v9L417fcLh2NRJTTOr
zp4PRfvMolzJllrHihmTWhjuZe8p0sWhhmeKSQgXrrkPb9oE9XEW4cufmU8kx/D69JHPJ46T6BL5
nudFQHfDHBNSCuU9qnKwcz4oJkG5nzoBElGXlACe+WnDEWFk5d2QeDzkMsSmou34yx4FWLWteJra
8s7WFD0CDzxg4cPNuTuuqNfY8L7Tv59Lp0jGhIfIm4/1/KDY1fj/R86nNozVkUtXzTHWKh130uU/
meZ5gZd8mMtIEv+crx8+ymXZwggVujIpWwiXz5jM7lLEjaJXwcALMfO72esE4mDDRBvEhgBl3rjV
Hudz7akE5VF2y/9CzSMck/X5YlWjvzPru5Lctk3UisJGZcEfylQkoAO6HfFojIB76iQ9S2HlQjmF
afJS7wgaMQPMvpKvwT4N0JuJVY16TkH+vsuGA7uESLKHmp778fIumvNM/ykRWGGMp9LaKJamFS/w
FrjEPxmMgYTJ6WdM46veEf0MWYZ+1BqqzlAlYS+pWSzw7dU9N4EWznnDPMCNwClpXFCiPALvVoHq
uXB4ezSzFOxPMbquI12ovU0mIa6NnNuwyuu2NFMO8nD+TcqE0CdZS3+LQxajsOotZq+tacaUXap/
+S3D1C84TUGQ1vcyVmjH3w91u2yoomYb29OhVOPpm28CVrFNU8ksW79oMNGivRT5zx6IC7Xs/kZK
pN4yeafizJUmi7+MkBSkE2290rr39ioIkbABqU4wquoEOkCXbLflcKenWKVu0RJvVtRzBwuh3ut8
OJNJwy6JIhW9g8mFcNM/C92WamQ5g5sqDz334YbOxrMJWkDd984kA0I+1DGGgwrECv2UJarPtgpv
XmotxlawEmuWzfEC5fn2fdIdB1hIzPcwntmPahYIg67AnW8mqg8Qk6d830L4M0Hydai4rS5DoVqU
GDmFn/s3etQH4aa0wCDgOlGfEUMuV9/iND4rENSFrq9fBR8qoW7cFDKk/65mz7nQCuco5auQz6M8
Dzi4SheEK2sa+nhMPYKaPom4hqu48rst8lW0ofAOFsmwmsFeUP/9JAoMPHlvImOP7jWT35dwcX1M
tAN9xsZhrdyqS8q9oW1tZkcpwKzPANp2erqSWjdobEOBIlkkFGZmVJlOSMkoEyHyeI+TODc7ruGV
7LEDAsf3GA1CNqtXWlH7Kv9jQuMFIgv4U8Uti2hxiZpHIX2YZ7LgeXZzw3Q3lFIan/1dS0n6dJ2w
ofv/Y//ORT1NDPs/grnB32vVsXI0v9MoEFd8arVaMpFCwH4XMmULrNK//NKR6R+sHIiTR7GxvjQC
uQhOhEQDpr5OvPsZRffGpz4CiuMMF3PSFDPCxBKmBolZGo3do9ig4+z2aWboALQQjb1mPGPwRtPd
X2NlekUrNYitx48uGjnpbiSvlCEjXdhmbUvaN608Z7FABpeZZKnpt9otL11iR6Ec4VxINM0p0ATX
WyjHyR7d23jt7cZXYa347eDE6Et3dqMhZsw4bwQi3aYGiLkz6BCbY11oSk6ZyXwWoiiQqugyuldj
96cLcSsCo+wYHcgO91B9GEqPVVMQ+8qU2WWWzNC2VBf2aln4T6iWsHpxlhkA62kegBNB8BujRIvL
2y3AguAqwTqDWxRkzzSqWWESvzhyeqiHZRU6IAiYgyhfJt7EKun3kp82zJlFzNy3OmEeU+I8SL7X
VGHcHmITM5aQS1YCNJgX6V/P9qAEv3RyEtJCV+r0PekqEnJiHhEAipCflftLerF64Fs48O+hV/QW
F65n9uy5le6OmRUbC4DRfL4h2ysmxnKOpMgExPE5Dblr4MZZXxUSqkYjfRhTPgawFtEdKsMaD9Bn
epDRv7XHnEa4k2+avxCPEybIxXTL0I/d+X5DC9NUWJY/ju92wU9d9Vxdh8K6VivfDrRepf7vrR5S
WQMIYLoaZV/MWCwtKX3n7rKRQvyzLcrginX7iimVyWUpdWH6giH7jun01seWqg8K5EHu8eTB8VYu
9qylaQwAbTA27BquMEd2Go4fM+bI4h6VcRYvJf0UKHC/k1PlNiEvw7Pna2e6BtSWhyK1cuSNTan1
8GtgVd1Hxldiy+GLZlZKyfs6iU6licufw8icylbAqCLN7nWclOKfzIQrd2RlozaSJ9XXyVK+Ertr
g+IoaYEbD3WqYZktfbgSA8A2VLaM/WHsBJ/VAoCqd61lR3E+ee+y46Z61cu5KllnPkAP1Swf/hLC
dXcfUG2yqPu9/gbtVAUjlXWbKJBNdEI3PqC7qat7VDxxv3j7Qqot/bYn+IogD+QK4msSuusgFEGQ
1h952AHuSpCXfoEFI4zYMh8y9bBFYlkjIybwE6Zq1Ukd9Drv56psR/gOhtp+duJ+waKdcA68lEeh
SXVQZg8CBt4SEHyulWaxHetn1hzcF9X8tD7lVyOQ/Kzn5smKBiRsCl1T7wTKGoqpZVLGOIfo32j7
J+O30B0kJM80+ASLErizfQHuaoXYwxG/+4c5CejknA9ML9a19lv3W6DmA/EPBGBsvebU+GJSX4Bx
rWbWyo5o2cJNBYBfrUJ2zEOQlvh//R1yfi4OMVfow3KNJnJSfkXpQBsQzeAXM0Ng92rf9M893frZ
P5PBtjGj7+sHYo8j+kJkMcKZA+ctWB6Wv/NGTCE0STtFWc1iDgkLdkKyLNdyRbQ1+M6wjzWwGQ20
3G8AM3n98Ts9HGKqzXOFDFtDaWYxKFPHiL3OXMukFFblW85eJ4RFhXjBaAyXVErNUtCncP/3V+oC
iYIYDHE7tG1CnZ2Xh6oJBqa6+teZ8i2fbxoNC/XIeWWa/Vz3EgjKwrBdxITPsYmr0irHZuvKzqw4
Sof6x9dJhOBchXxVHjUZdUrTVg90RVEwWdm+faQdBWdxJV9rABERa4eIZQSO/r/1RN3F24B+KdIV
/sa7BQzhoi4P63MQxhiq1P4hBV5uFVBSAsMR6Ubs6OZATdbi9ilbTDLS1Vw4SZtVVHnWNYSlgaRy
pg1CQYYpW56b9iCUZmYO8r7NcLWWbdV259RvXKqkiCAz71Wi9CnjAxEzfCD4WNT3v7yWjj3MthMF
ts8imVeUHjxHhwwpF+MtUFdhuhioRVOYdKr+UtCi/3Vk9w668+AHManP6wwuI0LzeceZ+bS/9/N9
NjSZepGeRgpryyhpsHn8PgiJxmEvoI9108SCxP7PVpmXd54JisbvN/RSukxMC5K92AVnlccOu+nK
s5BUu4tNYAE83CIUvD6jwA+QZsfOR1p/j7Pz4ONQdJXCe+/qN1FeTOjf5d7sxUssYeTj0/Vn0PlT
RyXqLe9OR0I5tUwWoKWGvbDrSG42Wg0DRAXmDtc7n/gNnpNElpBHO7Vuj/Sv5CMrGainUxh7DgGK
2RpLcwUQQwzBtEqdqUd/qQmfMkhdUXbG+Fye/hKrxG0etvY0N9mveStKzCS91EKl+LAGxk1oRBZA
m3It/zhxFaNRhyKrF3DaUPPiGrFRrMXZHUirk5n0ViVnkzwhlHo0UpT2XP6WHRwJfNdP6f4+1AU7
Czz1wrL9hkbTNJyzqS0fmGclM3eYSkISQc/DKyNMn3lEeqVow6GoXIipL+XwKfA8VIQkjq/EoQ/C
if8ciINJN6XzQNkIfxigMRXkZh2pom/50YUJHXaowuxaQGfLDvJR5+cHDStAEEs0G9tdfsJmYDzy
r7nhH5GltMkd/9kSTwQFoLTdIp4PO5Giad/tL2m/oPMnwCfDpeJWryBLlK9TWulKgKycnIGiECWF
MMWeJcMDlwyx8anJ4+egIK9Y7aE4lBC3xR38sotXFHhbfRu4olQ5XZcbBW/FbLgPk0ZzL992FJ+z
6AhTNRAbKuIduA7jx0bN/Ea+qGJrTeHGutceMFMBu6gvPUlikIExVcU//fdCu0G+arurl7pBWwam
bBvw88/hWtBH2mW1U/PeLEDtmNI05fLPE3X/K+9AC51TuWSDg/3Y2kfK7mPdmhYztN2CPOazCoBC
yw3pppD0bzY4c5ALEFdy/k8ckKOy0OgRVwdfJ+ebQ2bGv250aWldj4Tc9PwP4EbPKEgBc9a7sQ9k
9YA2TwjBeOSMTuIfigFXtzhC0+EYnGgAfUWv3aoYKQk629Ned7nuvli0gjybdzE+W6QUcXEVP8XX
tPm93COtVnqPS7RODshvvXGFw6284Dj+ANHCAp6FGmRCF+dWI6KGRZGyKVt/0A7NRRu5FfGvIMTo
nBMbNuYl4GQf+oki+wUo67UaotxWNCcs2/4Es7pflRNd+1l9g7qx/RO7FAvd/fJtR0U1XEshhWDA
lZjUH+/MRiFfLfjLGoWJ2aUZYAj9Ns9KRhV5S23RnLOohi3cUkEO9FZMuNUXTHqNDpRMAF9kx17j
10VyrcWRdhQ8hOM8tF7bQ8jAA5usAUNFUzJgvwrwLJ1pI7l3JoP17QHIY5QnuQ/AHO55m8JK8Xuk
Qp0p5PKDTl5BJndYgAHi7m5TjBqCHQuaMAWdBZ/nNZSBGYoEn6FA2SGq7mZtXRHceSHqXeDYFTlS
xYtHXv6+4GJmupDYjAWf7s9cCm7OjTyCg44VYEjtAM00dXdrZMdJ8GBGVHHI2+gBpkJYQF93psl3
CzEf6yo0kmxXypMsueAujmVbWwhW/l4cSy6IIQsVbzqbKa3QyvSsCdxkJtJCVqgdwfpI8Uvk1f21
KIr4JdXKvMCV1cZdNqRrPOsxaGd6K4tZutZEDxj4g6wIXIkOW4VzoTv56ZrA1fzsTCTy7JdPyOkl
kkvgoSt/lVbcKJcPSpCSztCDhw/YQNHp+fJIurazEf2nVyIEbUsbcR8SZLJMDXLREvW/POP84Prw
Yr/39QMlsMOCrNbFzWRbDrWmBvntniO7nW5LnLiNpwGBnBNHkqX5vB7HFUqkQmPjcyEE5fkOs78H
qgCaLyb39WbVI0m4hsB62Nlz72HikfiJ2VDuaqTYfK9sVgsspr4RXsAfkY6baLGHbl1z1cMzRkU4
ABkcqPPhBZqfx8Lxj8Ur0L0xCvyAU8AAJEYhZoxwD7R4di99L1zsAN0VveM54fy6osd7z8llv49q
FVycq//qYmOIm+1gMh3CiqGHLu9H7+08ZNQ99sWi9DeyxbB2T104/8Q+yjrGXQ2Z+PhSe+TybIno
HFMtV+jnJYScLdxCmY9oPN73OiV4j1FX5KtK0h01UgwyUS90p3iiXxY8efmWJdXXqs5D2S1zMhr2
0vALz//iqeCU9+Dk/Y1d3OlQXL/tSqAqV8kV/g5NWfByHj2u4z04PblwPiyaTQ7x6vCgYwpCggPH
f212dTH3ICVeRQx0o/ZThdnNzucxMmAqdEa7zysvIE0uNO9dWpkzAKa0aUB7ZKPjTmQQZWbL976O
6R8tWewVKkzYu4VmaD3wjjqa4CAuMRswgAqvzRexJdD1tub9X1yL8d8rHNNeoKZOZppnWU6HtTrs
x6tPrJi7TO1U3yhr8wwPDIb9+R0EeBHWnVYcvfogwTOpzxwfO/LOsJrH0MiOLkBRJItxXlGgWkRu
zXkucOMWXoFxwWWkVwwjuZH/7N8u7/62ydfnOrRRJAGn7LB3OG/69eRc1gXYOYtiVuOpk2PrjI5l
bB86/toWHrHoxCQAzto40SDEEzV9XVPwm4KzZxgxFri5YkeXQnGkwFKa1oUbvm5mrYSJv3YUuuku
zK9xCWcxoKz0hSjP7AytW3nbdv1Atrneis+X2/0oA8XsT9uufrfWGV+PI8aUue17s+XB+uGzGqg4
HnkBaCvtKdtgKCT8ykcS0ExIom9vEQ4RWh8//NKOITZkwEnnf/JL4RkiG0pMmW+9KBy1NeUb4QPC
WOYbucaC1p0ezLOUyN3NBOpLv7OI+6akVS5ywKq2kS+3ICaQHLSE68GdcwSMQRtqFJNsmJvSTl8Z
0OUSYtp8CUdYQcUhiMmJfjJ6psdt7u9hoTrMInc4Pj48FIpVATpWppY0aPpkCZKlraN+SH7nxoVu
5n1CsT8aOt9LIWVfOJY3I8OWlaBcg4oYR8YlZYoTkot7FFdl0+3Hq8JLlAaQagP6wtTM5CoS9PiI
odLrNUGw5RaGR6xG7H6x5gyU5vPZo8ePVjFISqfNbhsuQUItJlSqwEY57aeMleP+E4AkX4x+6R2o
lfBKqizSJ9Txhl0yER3ILT9ewIPrD0beSQgab7HGL3i+JOUdysDJedagIcm9nlYbQviWWoEv15kY
5MCqhk/SZgPjQ066Hgqeqyy4e8Kgmo20YFP4LuU9H6+kvBaV4VDOMuOhYL2PT5KDX8pkDS4clpUL
PxGoNxtzWxiRobA8jFS4KK/MBVsI69PuJi6ixAGejp1tCxKlanznE81xT9gLJTOjAvSg+UxRoOkI
BnRYm826OOx4l+J1gi/OqAlUZzEtb7dgUj260tJlxgWSnSrb1g13a26q55oTPEBhQyv3D7E1uzXs
YUuN1KjjKPOk7VXAOg37j5kgkbrODdSS0xU2KKq5oxxgX0E+bB6hjzgF+vW3705Wxm/xu9GoE6ht
97WD7dXuqAF+/USk7iuA7fTGrRcY4EmNVtLEh8LTqqMnN++UmA/VnCQ8e9YvNCngqzST+GU3cU5N
ahq0JufqrIySx83Uq9k/3zMWmN+/x/cWQ54SQrgK4QYo4dbifiex5miNIYOKMHpyne2RAfZKQy2u
M9WaJtg4i6TkztloXKwfyJ/F1u0XtMZH6VFjdele/0YhfNFUh5loPlBRVPXRkosBZ9jx7N999JGa
xn59viLha5Fb7jVxgr5Bwy7M/eqWwaAxOY+6O8pW9yKKAT2lDPtUEWFrQLmybBGnAxw9Wr2NG5yj
Etd7cpxeH4LYmEL6nC2hdOs0ml6dHe7cpuELBcx08L1nO5QbDzxWAWwa4Fx8Dizj4T6AZEWvKiYT
IioPpUW4dLMjLnYFqLWzB3K4/6NYAXQ6jY+j9cL6yXIWmeydlzrmpBH9izgkYrQKBb3o/1VMoztD
yawDFqi96P35tjD89w7Tw8+YKeOAM+6ub4J7/GQdHl130EuTVCn1x4sZyy8/AzX+wjF2X6c+WxhC
NNUaiC2AwRFd2ig1fFILttL6ycQ3TTG7Qk1NO62GDEXqvK1d8k3Ojsk/d/ur2yQ/HtqwFMV53P8r
NhysA0HhwiPMJz+O2yHxr+qIKQt8HQmdnOSGG/JoMYrSbWNIxNyFGVnyYHUyuQ4fdo8A+fAU0Tzb
zmZx8eRGhca1eXHC82BP7cnhdcDVdomg+zS9mwF7OCuBu3FVZNM21h3NKcDMwWrAL8d4DXKXTZ4p
k0lnhNkQfZE4+qIWPm1abPwNdPEz6koWX0MrDX71O7ytUV7Y2Lix/7vVF2XfALD7CU/P7j2TD5nS
qFHdAb0iFO8nO3kc0OJ6M8aS5gMBJtpa/3X+ZM0yB7zgrUjre64heA7ITtgs/WTPQylF2Oi07mN8
yLV5q8lg4CEJuE+D2PGziy6TKvyrNCsZW2OmzSsbQUQe/azZaUExoQQWkwFi38F95IeqLVXHzHKq
o6S9Cep39s0V+yTAiZl4mtZHTlgrQl2lofxj5dGM8OfxlLDGyqMg9ECSsMCfQOR3pM5jPPs00fVD
BdK2wFGDZ06hdxFnS11FFkvFVKLt8ljAmcY3aVWh9FFDBd8epaglLHMaNJoCfn8dV6pzcaf1iBDZ
dSD0SgnfC4NlCl5Zhli8MWNjNoJP64onIzV+PxPcxUHa1Y3KpYwucN7OUE3KkgnJTSB4COToPgQG
obaYw4RVv3YzwuJFQJ1RfBK5ADsfuCpzR9dOiXbdzB1YjcsO6+iijvxgINWpW6QBkuF5LQJdwUUZ
yArJ9aIy3sXHWSNq+qQfC2JN9DIaezKrnxYTBJWgjMrT1j8ouaGraBDavQU1+ZPO1ibSOlqJbL5Z
lCm11gMKJezqRitj7da+vDg8VW214BDXuZnmTKjXJSf2Pte0Mm2LfV5pZGvf0AXyUZEab7d8jZRg
qCGkOERGnZaQW0KE2BSb6+BBId+QzSCCZLeRUwrQAe6trgsWiwZYX0HbucDdpbT7uGA1QXQTDYEu
m6mFdrZkAHNi66TPQodUM70TaQGhovws1XqLvWGqnRFalLRcmQkAiR/xuS3FWrP4FUkFeKEsnS+b
ykuecXWl5nBeAK03uFK5QFGS23eE74vJ3sqVXwRMNiPhpd7Kz0+JB/fR/pgh4JAsjJwc0PsMP+2x
gluqRz07JO9crhqKNXdh1bAvM87NKDcfx4o/mQY2HqadyUlJgNReRKrieL3ecZM23VYj/41DL7dA
B+lQV42j1C3iFyBVcPW9RyvFgNKSJ4rdxaDNQzygIuA+33Cy3KQDLmDigIWkbkqlMnaafaMr4Z+e
r1GsFJgc+daAVYsv3Sr5dXBTgve+BYEXxB0cWDZa0DdQBczBhyOjrBsYeoh9NyGoXgKo212c1mF0
15D6RbcLexMBPy0hDBNGPkpvsW8C45195HjX8l4TiIxVwKHl8bM9PMVHPTzgPWIduM3lSEGyIkex
I8z2EzJKwdTrLBcqa+3HlIDot51m7of5zf63giFEmK54tlvUOld8JNmMwllQNb0+N1YYDXoL624+
wmlf4vh2Og8jqs4KtCWcgNBB6wdr3okAl1FU7QCriTMo/s1aruJZVoYf5cWNx9Ovx4T1ikLxVAQ8
c6OX6H80uO8020AEK5j0ZG1+sJpWgbG0k3xrAnWYelz7ZyzO8sO4eLhDTs+x8S74z+l1m06NDH9y
Eyz0pkqzgo0XbJfU+0YDW3iALQWnLu0yM1BOshfaeGfYUbzzyRb/v0eYcbm29pJo0Rt/pewSnGmg
hPcOOBu0EoUOrItDUf0byGYoobZcYzxX4Yc+eU9Jd+wrkty2hH44t1UPJPo+dgd7AT8us+FVOihm
rN8DYJqll+MSaZctS+bs3VDqZxZ4yGXcgg6tkhVk10kHckR5S5Fv0BO2T0/3g+KjnXLXKYFwBl+4
MvxhTXAUCxTmJ2Se90kDdU3EMVuUbfSc58/zBIBg216jWDNhcTCKrs5w7APqULdyQiGutnZ/QjTP
C3E+WF+j6h70vdLUxslGik0vE5LFsFnvxutI6Dk6EquMRHL+Zabd7ymaiyW2vubF4tHkWsmaJliM
6ke/wrEpsAsznqtM7abfdqXQ0rkIoYzsB7q8vtDvqeOUDx0EHwhfgDpjlZrgKOigDNvo7nm6aDug
7ZymmAwPLRj0XopzNw+X8mAKZRp7uGwnz2xjNM9frkXo1EJst4YOtmb7iajDmT+X74Sb6QkGRSM5
iVsXsovxfkhifxBGwPdFMG/m23jRQwfvmXftzoxCx3Y897D1ws7VaWmL0G9yvWzp1E2XECULhywT
nnU7gMzOSE0qSwjHnJlVqG4+Z59YyX4UonLv2syn3t8bFwx3me07ysHDWJ9tSPwUXQNez1tIuL/+
EU1dXHxGwgqGejqjrj+B+RZYehTaLPcdUAg9W8OJS6+h/OBdAtZipSB5XyNXwbeR17HIq5BhBoLo
Ea3f+Yr/Kqtbl9Eic5tLHmARhA65qJm/uLQQeNvzfZ6UnCoFUDQciWOLYpgBn3n0Nh4vd+6RDpf0
DkPzKmhLyYXwEHIf/z6/fh+x27KOU22YrvwgJ73/YZaGgJUGsiR2RS3t+1D8DBMj1M5XhycLclET
1nP0QLVQuy6q+xIKLRufd7PB3nCxm07BhEEa2q5BhtvHCWAMJvVCDwKbTsosPFygAxlLah9JE04h
yN9fDrtPdK6SaQMRjBTa4neL4kr+AQC104I539XlR2I5C4Qz5OWgZgtolVIlchnP2SKFLl2OdoPC
1k91kuPd8Qp0m244uk5knKfuMdORkI1Nbe6A5dLRdahfqP3aovvjdA8zsVjagIelhjSBEqudtiuC
boys+lG94TiXmF4pnEdpPt8saWU/1u5uTM4bxvAZYSa1rHHMsqvGSez5OJ9vXVrcbysbFEB0mNwX
1xXleF9PJdsW1Vb2Vpo3MH9XXRPmifasLQ5epaV8t+3xQu+cKG6iy01t99HqaRMJW54j0PcYzQ1o
Wf3N4QA82tBFh27hiu/F9Bc0uXoFAXp4AL2dQWOsvhsT12eXYHaypJg99yUBtgIh0YcTlr2l8MAV
uVmkeX7SSIjknlbhplrKGW7FMvb3NmR9/riCg8Bt6i2dujZ79ot4YSYCO/xUX2XkOtk+akx6lgtz
dzuDFYDJ5YiZ/eJBeh0h8T6TdIwAzBH4GBMfukKqU5TwgHawNDyZlyM1Z+7WiEkogM702/G37eYI
7VGvD8gWWusxVprsk2TfRUObeQ0FEwrrH2rpZeE8winrStBngrwIxY+ogr1HKOHtaehUdOe33NjA
q/46Rg+4PifzBil10LvwYNhPcI6YOh6EqHfl0xr0jrVPVSAR6AY0dbe/VbSVKxjwLjlxbw0/irqZ
oqVT5Re9m4LTudocLf0yxD4Ss7if9V9dSeD+t/A9R7Vk5/XUjVAoHULYJLe1Mhufh2rMYb+kQbX1
0bF2H2MjLwakTypAs0NlcYgCPBOAZo0xVVVR12IAsftgot5pY3Syf2sKCHj+4chDmjISUpSCIQNJ
HCynrXW4poR6ZXPQhvne6JBrqsCcne02ppS+VgIFiMoX6OWSWun2oXzPB4Z4rF27ZS9gdaygUlyi
d5yIQtPkBamrAit4Knr4pw+yfE1Zv8QfH0nifu00UOHpdSoui80O/t0T4XyBCs/pPKtupPIJ0Vj0
0MNKFV70lBI2UIkrjlWilHUsH0O+1PYBOIflodqLdNhyBFoHmPyDcmfXAabxjKq7YIb42dYaiIHe
eCP4W768PwAa+CUmU/pnokHvQNhxYxxepoLSXSKQ7haypElANk9Cw8bw8B+0TgnTrF1ERb6kFPcJ
eBCWdnsS5R3bg2/fISWnmkZ/3pmF2xx2mDuy0adx/+pXHlLBWqmsVcDc/WI3J74Zn1bquCnpz2Yk
rUipCkIeqxYjxfaACZQSyWiNFfeJ1zcmVYvipamLj9EE7Mcc5grtvD6qEhN/8PVKP2/2WavgRGqm
eZ0AOTx9XbqK5NrVPKOaDGYprYLvN99+H4ePRvuznS04CEGpOaqxepfGRLUVZ7F/x6bjHMq6qUxK
Rjvz96dFY4oOtT75wee8qe6fB/GQtRzZtC1/GT1evC6r3/2s/AMPWLMvHKRV0RaAL02RDfulQMVN
e2WhQ01m4QuYeFGbdAZoQ7Mj4InT6iytIOBBjz9qqKNYAECHMjZgJDuWtC9IrSZt053aWOqYroQ0
J9wSSAKhEUzXxk1PBZ5bU2gTsuRVLGKNQUXuvnfOKVcHxq6AQ00rwy0Z/mBepts9eoo6a2pu0GKL
FcSaU5//O/IJqtyQcv9ZCaEbT/tIQbJdLeVCLpxo6qX3lGHMRCyboeJIjlXR3hvYHnzKPdnbWHdD
T+x2v2XhTCSZerED6pke4F7z8XD4eWRfEEHH5vPYCiq0ny7qtbFQ5UkMv186e5Fho2VWPt/7yfc6
wmvzOA9alMVXoOpCg0dkmGze+nxHGchnvuXP4Xesoh654UhzunxWXpfqDCJcOeIl9VAUslqqmlVt
BtbVodfGgi4gPHncM7STgf56bXdfC41xYsX5XNQjEV6DJo/jRALaG1mu+CahYdlGowBMWtKELeMe
L8n490UqvKBCZ7+4AgbmykkfOswoflw56r68RyiaMsG8+yukhsu6aPus7uPIxJaI72k7sn/94hSS
6syxkg3S/3hPrZymI7D3AyR5L4raOurYZLEdqi+afRL7pWhl8nYRqfX/f2rg25tK6Lhx0R9LcS5j
yhxB1jRF/oKkhd/JWBQz5aqm4Uj6lbfTA22hYa7QFWAPJ56LGnpwf4Tt5j/jVWaHX675b/52/M4l
MEXiU9iTC1BzczTmkGS2Z+apyMb2pLsib/gJYlCoC2Egvby/lJkS5CTBCd7LZwNG7J1YeI3Yf1NR
HpJVH08YHftUXW4HInHc4RSiP06HqAspKiLuqE3SZy+v4aT4Woi7Q8IKsjTqGqyKriwSJyyy+OMc
4rnbg1pz+aAeS9BvAGD+xNTI8T58j1p18vMiXPVMbw3Nh6ID9fL6ZwWr0H1dZ6alRaZ3K454VfjF
Svcyoo7PmFMymOD9Z+9gQbbca7MAGdkB3SKYp0s3F6s0QzVKfCwmwFa3O9+RokZEOmda/xpKv51R
5JCEbGy0+nIBccplGMEW5+3rU0I0XXhb8Z9EvKBkivbJzTovfMv0GoOJ/7Aer9gGChrKBn2vTF3x
2n3VvpuGSt7wPtZHzsevOBKPeN+ynG7ceFzrwbRh9JdDtyRTL+pmpkqOLj1BagD/n4PYvjZxmex6
ccNsM3KqLFtLyo81sBB/eM1NXZRhCc6FFR8JkfdiaSeEaaA51x3iaQcpGA6YypFfj2Woogln3o22
QC3Evdp0eUlUcR8QrR/VwQ6uLlxDmtry+r1m7+Xd9g0YCraQCLhGTw8vhgXf83AgsuVw2Ho7jjHB
HLIzN6MHJl3In8WSdD2nTaU9UIF1L2qgJCPlWkOAhxIDF6e2AVH9AOzEWaqFKB5zFqpAkCd8GeDW
CeMVH3yLPdJRN77WAtgxIjq5Z+xtCxMhQnoz5agHu6Le3hnQtYggK74FiuG8GrFrb+E6AauIYUgM
37OdejyDT9X8qI+ZCtdVfYokd+cVklQ9UM2ItzCEtha+m4GS8Y2FwG6vRHm97JmUMZ5wRmmAKwkW
c0TRziEenmJc3Mr49ZYeqazlosIayoIPmR0ahEaIj5bk64qQxRd8NCl97yrls4LoIO/sJsf5EaK5
SHgHwtR1Djq6qdbzH7TU3n15fd98Te6eX69dE6yjkXYfSzPOv/8sIscb7Av8OmAF5M+o40z/dYWc
a4m9E7lIsVBEetPHxD8FXV5h/az4kBzF0mX3ROi7Mg1ocH4tr90WfiUYVv3ovoiYDS4Wp68FBVSo
IAtxJGdu3skeK9zxv6rkZnQyE1d0Ao2sEcu0dUmZ/8Nbvz4LRa4blTsQ7WDaaXaL8OXbKc4+slOJ
n6Yk2Nbvm6yEdGuLBsRCJRctOgC42OY4Z1hm1hx/+IRFjoIsfuu0iVBapEUxCReBM7OjFp9I3fHA
TFwHsEZ+HXiDoQo2+QXBL/sq69y6wUVu0qAr9O63Lub/NO9yZkpa68jCwo/Hk0AuHzJylPbsf3tR
2MkXpHhpQljVXupARILezb0NnR+0w9AkdIXLa1xfTPe9UdU5/eMF6BO884owfnYfywDc2GLGyIta
HOLbQlLXKeqKHddU03vq/JLJtNNDOxaKbe7zARadw/GvOElARj8X4t9r0dvBrjiGQA+Ip7146Jet
JOV8jT+wPvMK6evIScoh6aK2t3OQIe6axYU1NU/Aduxb5DhHMoPxL+mKFML7+r+EfP4m7BYs44OX
SNiAyS5CfGNEqicRVtT8cUOBKs2hHGa6bGBHpQVmc9vi1xSwvd3Mb1/f2v0c4lv5WGt14s4luCqY
0Ys8o7jY8x1Aa10piz9jFVQEjaZHr9bBWxPIVBJf5dHR9FvGkz3/H3pIXDfAJ2JQZ5krylR8IMFv
TTHTYgbO5QZ3TRd98mP/gqNNU+j0Ds1xreAFwrl93cs5Yn84yMJpIOfZ8NpJfVPcEoVb0EBcvmBq
jtKOS6EBM87YmRXnDeLyrT7NUrRJf2nyif7wSPSBVdYU4tgV/SfZkS57zg6aGnJRbsbFunEDVgZw
tr3wNihMdnxwhmFXIvfBBys8BG7wgh7+byZbEuP/5+w6fcblvd/bZmPUm4LSDn3Q2zc9Fj2R7E6c
FZaVIh3evSlYBANnEGywgsh9ek0S7nyHsB4lweWL87gm7bZapb3Qf/AP2ewsDml1I+hN880Xj6Xp
yngsjcNDjR2oAka5s+K650eCOXiunphtotmtyCiAUTSMibLKVSuPUzyuxU7Piy6aBu3wx0OFf8t1
m4Ig/lk5D3Oe5HmA10csDNzA7ZMUHaLTxXceB1vttJITKyfvcB54/Z2Yl3mzWBJdcVpjMU0ogpmN
eOh8NJxDwzbgsGsng4+oAIN7SRVpOSrL5Qc+M0EN1l9r3secxIbj23e8hyc2gsV7BS1yAV3DuO7f
KCqyD46hg21VHE1bJlhM3O6lXL+aMtV66SbKkYM7tZNOi46S6qiBzuyntd0fpnDC5348haYSq4Od
8XEVkEOmzqLf6VpqS0TQMm77+RSJCmknHpBVdtw4SYpZx4iCGjRPG9AirjdE4JEA0BIOTqdSpRnb
oqQ75y8Sod1/ZkXe0+EOhjLzEPMwF5hanSIf34qYDcJbUejeP8SKquKD6+5p8Pn8Kty8wOJGN3hi
qOZsTlgq+s/vF6SzA/NsVl6mygm2U9Z6X/QMIyVB1lXJ3KbijshEOvNRGi6uyImr2SchJbHgOOpF
xvzz2Oh+VjB0hIzwNuvJCLHJ3B/NcAcXFyMdYNA53sZwtZ0lshNC7UP9RCxjCU38F3/e4nib6X8S
imqoDSm4tScARLoXqLI7rQBM1zcnk2C1m/ERUjMLxOpKMV/JSuY6Gulv3kry74exeA9iO9i7JErc
tcSrUbdzJinMVoTk7uZV19/f/Y71/I8e8b3ioC2RuQ6bIQOuYCSIrC8PxzutnKB4Zrgm1c7Z0LSV
t742rKMsJ7uzs5rh1JnPguhry94s+RPExENIMBNyn3VjeY5Rx2NDeJjtuY406nGh+BIyVurtl1Ee
Q9BrXTidE7Za9vjBUXuTaft49IJjRURHOPqvv4g5vvUHjZEdJp8rzuaGeAposnjLgU8X9fFqc3CQ
sUkzxwUy35GuOH/InGyRdLdwVQCn34PqS0yXEALJyDLyJ80kSBd2VQ+9cecu/3ZedfflqtlMDDx3
p8QFUboNWddSFp0D/ZxL9yhQsK9/svAk7sCsXkQ8Rn+m6qOIEDQ08PTEwNPFCyJzd8McMWmDUnYk
jSHDfv4gUvOiO2tJ+TeiS5tFmmX96o0nPiXRerv/ISj7m+02zM6W7mFBtjSMvUbGExapPZxf5cU4
n9hLlzk95528EcaymOPL5PzmDJG8+fONt2B7DI/KlJAGh/nRfa/6VkjB6xynguLnjNu0pVah3hEg
wiOTOPLzpF+/WJ2twfxAV7o++wXwAozt7d4+4Gz35cClBsa5saY4PU0CaK/ZFDpstU4SPJ2g+fwd
nIeSnof5zLuHDJ8kReKlieQ+4USZLBZjbXZ+a4lhCWVDN9p8pKxXN29UmcPbsFzSoAweMbc5b/0d
81NrtHYou3SiR6ZEDCO/i30WVVJIHI6WGlkir6wXg09YmMFPkGAgi6DjXPqFrEquooE9vLPP/hol
w48CD61txxC+G4X/4shBwO7qoIpiVT6UmHYpsOsieDqkfAJJ9GGWtlrxgiSqChymVAMJ9ht7DbRZ
8HPt1/s57tEn9HfFUjd9z7QORBTwCsLens2UeG3iKvw588aBOgWNScyPU2LuyRMXDb5B5j9sUSmw
9I9EY+EIq5/3Tv/K70PlhLECunN9AmVH/QkR7IiVGkhxk87UqiM60BWhB6Oj0+UZQT0n7/EypuuT
+NiGYvz4aWZIIL6Lg3r0K8GJvZHoor5RhfMv/3l/6symVcmG3gpMdNGJ9Ki48YUseX981xzDjx0G
yzvlvEGHzfx2jrNDNrYcNVGKUWgP1zpkP+zGysfLZ89xklHDFg+At/f0G5iM4rhNiX+8VmP6XBlQ
wVNewld3Lv/Ytky2ANM2uQYriNI/vrC8aw/FcDR7zeEgwm3EbzUXeplTlz2yZYMW64YQ9mtLJd4g
jsyVu0cxIxQI/j8+m90ca7dla1xo6bsrn4f88VIAA74OMVjeamZ18csdPA4VZwUxdTNa6dw1Y4PW
VCmV2FzYSL/TUDeGv3Fo3cQMjWWOYXioqy5+aynP34lqt+gEr2AhoHnugd7IuOhQDsGBpLkUm3NM
fifs+QpwsuRlb0ZvRH7RZjuUScXjZ5KeN6lXm3+yhHjVvWU0jFYquxj7imkSBhiqOg6uOMJGHmZf
8cdZ9SbS37i/BzWyOLzJwfhWR6lkPf8pAhMo+W6y1ZZWHdbUDRuobvYOZaPV9wWKeb3Bj0Fibkt5
zPDDk/HMq3KHEMWyWcS4KYzwIV4JIZ43t6NHj7nrzM4QlUqa2EAP8KlCQbvDFBSV+l4ipR/ckkpg
tKjNZ0r0L87IGuotcFdx+wy/YnUolltOHjeENYJBp80DpnNvNJPKQn9cLUmYDcyiK251uAttNLTW
KkRCPswxdvrj4zbm80P0/wpfJgL6pH5YFA2bTYVyu7AoZVsI3RwcBG9JY6tAkNF924LM2z/xJgzw
Puvtm53TNWRB5XBMJqfEiUBb/RFBX15LdxrYlhPY6oMPHKc+A3VA9bv144r+ngyw1RKkJcpx4z+C
jYoYNACGskph5HkPSQpuIEGnrk/g1ypb/I6wIper0tiIGFeECOp2lzbdqJjJ3y7/1EjLmj8HTqKD
RQsGa7gC6dsruvT0wElEf7nKTeeUktxEIEL0zDx6ZHmYaNAzDw+muMvQU7CY4fVmZ4xURRt9RhfR
b9rLTMBUpXMJLPI2tOL6zn2RcI5QHRtxKWOM1z2V1pSLAGRKj+4S89A4guM/gsJ/oM/ldBWqjFB4
h/uW3T+NLSxgYlGoXU3cz/cbsAiOkixlb3iB2r3sH6cUNY9JDC5/ZYwDguq01X2bKiYDl19lnkQg
9QRuSVgCBpqZruWtG029OgMu5bFiq3inV7OpTvCQJzp094EJbDfquxSh902F6eZtsICXOACB6gaj
ASxqz9g5W/MdTO3QzIQSHmNtHrpVvREbiRsHxYUiAEx/0kqxCzikTY3ZuRWngVvNB+nNgC3oi5SR
4tt2/NhWi/eopFn8909jrTGt3aOQYrGiCH6lkoD4cCBL5eMk12l66swUWhJ8wAo0mzjLcbiIAn5T
Njj0H38wyI/aDTVVVYlZMwYphViTHugsw8bH05y3hgJ84OEDK8NF2z7CgT7L98kqx0HJmLzHjPv1
2/ekMwZQiMzXxFPK85ep7rUI4qqBYwqQ4EuGCQqaD3U1coKCtGrg13CcEebWuZn4xtLcLY/PU3bq
DH3bbnw/Zg3VpFWjhwITwjMj9oHnfzinrPAYgRC8Cn56AXVs5i9hJntEDLGbdBjEO/tYTSpOF3Sk
UPJ1DeJLlBxp7RlMzdn1aT242cGeQAxxL8LeOnLuyiADDc1THp+Cl5uX9uMUwm8QTIrgQtdKLvYN
kTZ3SGliLqnMM7t44+jAa4YCLDqAhdRNC0jB1ohiYMm9nPiMhrFJBWzeWDIF3trDsN4HnMNDXmXt
W2qkYm3GxjJrxsa72d+m1MIhF2wl8yJ6JyQRREg076rtACaHgToWQZY+BNIM2PbobRiVvvjZa5eL
WkWnGh7ql7htF1MnwsLFYFNXOFR0nhNYoVuO3n1lOu48zFs+cbXohRtlYlQwgMb1MSFY7FK6k4y5
xZ2Ed5AiD+HrhFWFaQKUu3JT5pdl2/mpirQLye0UCKYlQsC3XaMGcYWTVv/JHMp5p50KPGyR+/PY
o2Oi1wUmTljLNYDVCzifDnfGqSgMrRJWgyEEiBPckM6GKqzXgkNri8lI3uGEKoMmfmvtvdrJJhd1
d3PyJlqniQglT6L9hawwjIiksHdfcvaxPLBxdlJz8QdFjhymJLveCrqt+IdbDTstl44me+Dao/es
FMXhP+Poikr5A7PCtWuQAnictwv13olxdQ2BHobFqfONKVWmylFFdJyTPec8LaypD0LiFGyUmx3X
598N+H3Nbqsun0uaEdXg79kk9HZ+QY/8ka6YbSt5uumnCcKGBzKsV5+8G0tbtgTrrWRg1qQcS03T
D4jZ86XhJH4DF00rBhSvls8FsagUu+uAWfj+BnOw5mVd3nrewlu0o20O1/lmWyST2HJhcokDUVcQ
Ycaag2yH8k05zQsJgWOTLEO9z8CW+55InlBZAhM2vpDM8K1RJwR5OPe657/smG1S4zpNkknLvuoo
9sIcJwq02YBmExDJIIgEL2jt2j5Zej0l+1ZrY9/UtCtGdkLaiYEVbw8f8o2MWj8S7MQFv3DYUc22
JBVFInnEhWJ/aiAs33GaaWVf36VyTctluq1KD065mOpPf/f+0Xcc6E8IzNzSpnMDNTyhtCkBqALV
62NxArYsx8RRETKrm5Kt1bSu70AcTjS/7Vsmu5z49h9ejTeM9hl5M1fZFkpYiO/K234RNJLCv3bT
EwVvrPFq7fGnAIZFhzmcGCB9/NpXXSaL05+QR0Q7so1GjnsIA1ByO7YXeELHsFR0ySAomU5TkKLt
Z33PsxbBPPXyXsEYZyOldZDVqSQqegcnMKbNMG9AAI5x7BdRf+2LtYMou7i9WJM9LRaWRNZu16wA
haeY6gVdISpMqNPiP9fBZ1GFiTkvmiMHrHV0tqHXNJ3XmVteq6WWUgOrQ85LsQOE79Atf7501L+t
kdWgYQPDi1RyS4BEWoMk1Y5zfu007TN4+Ddb3GaOzhPoWgpUXMmeWInxMJiZbVWwPREyqlk+20LD
HOtx+oi44PlVqey8NlLMB3/pb/ZCrWrOnk0kUcHYTDR+oIrwZ/TVrplMWqX0jWfMmfE00KOte3KN
setwgWQZhxo+eSBt06M+4yyRxJwysCADfhkhoiCuxbklF5DExQ5m5Pddq+I+FmT8wb7278sC/F3c
Y8GVvCAAptNK07/GsDVeuQ4yXibprsO4rjG0cAnV1DjBiuVOiS7U+jFBaOCPru/y5Jp5fZ35IuSE
XRtCSUSzSU7CwxPu2nYEzhDoPwcf8reaixgbA0dYmmlMq07wSpXcVLhlLgBfmj/HFfmFyqczf/5S
lLF6u//XewqkvogLpTYWazylvysAoQJPxvHl7D8CxHU7xGqxAiRYlkCZT1DkMWqQbSbIR7eQ+p+L
f7nZz2JkKHnZ4GTXjvdJwaotulIok3cq64OjhI72v9r3TYwXqrVzVdIER4eRY0ItfioP0DnaqIcc
S3XK+fTI1ezVMC+0hFKD6X97HZ80r2/dERJGBc7kEvQvLqr7huZ5atwu4hlCIepIavb+xbg6RLk1
PkwRhLVPZINJFaaoRANtLiPGVoc9iI5WDgUCj/+2LWlBM+PzMYRqcY+9FlBGCqc4H6HCk8sF34KG
XCO7xAmQ8pVxlYs3zx2hDjVEqrC4VJ/b2jH9FzyYlpLZNWRjkIgISmd9g/lM54EZ8kWPND4h0b35
VOrzHqiVkxzqvmTCoP4AM9pkLyqOpRzPeLY4WbgNN6kO9bzURTfz9JFOr6SGeLUTCzUH7QbTLdeh
8bLl8LdD+rvTUi/46yOwbMcpGkEANSlKuAWapoE1oibU9ZoZEO3z23NcTGjyRifu/kRbmEcD3Azo
DtYW26oQkkEDVGKM4wDw6hEJQvACT+3p1sQTJ8aEryNmMcrARL8712d0c9FmASTOlZkdr9l4tDAt
vJM3YPg9vCxYtlOT6UpATj4Z+A8oWuHIupy1E9FLILznr250uA6IVus0f4bbsHYGeyV5Li9fmG03
7KIXaQsTinMAXgtCwG1tEckcxVqP1FjAoRauvTQfRBbJLIEwjU9WdJftJb/y/9/MKRjFMlxCUQB8
5y+SEs0opGGgnnvf6//NrnligLyOs50wuH7n7uf5MoCT30AlgBmAcvr0eMeMkRwtfrgZHINPSCUv
pOxlgjgY47RKp3akGOzpl1nlknxViJBZE++FULjqr1VE34DOdP54CIWjBHLCvCoxLgPw+eqgcMgY
N1IOfX6eoCBtfQ6RzpMoVRW0Lpf1T13U5yJdEmqq5TP3m3F9kK4BB6CL9dzB+oAwBbM1ZIenL6OJ
N9OfozhzfF3tIrM0oyVYZ+2Fou86pekOMdK5cHP+SUXlcZLSXMXvzliewQ8Wwa1oJAxNyuchJhxZ
+nuZYRqxWgxhbbX8Ge6eeD1ECuKcA5mgwffwj+JTBiKL9zuNqIsSB7c24YbxwYNph17XLI//tLDh
2iPbqV+bq5wEqI0jvB28HNiSWBzzktrd6/L99IB/XwO7yszRbvZknrKDvrdrsM9+wfqc2xMrmTLf
brOvl0qpiGSEOJvaNoVmPnli17kHJ1tcoDikLtYlXfn/cV10+YRDwxCngq3vo+z884jC08YbO4Mg
CO/zOypjPxer7rkJtZ43qMz+J7bZRhrgyWLOeetPUlkblIiO5+9V64zqAwkunG+QgFYLtmpv2y0o
oQZUyhn/jq4Zuwq56cOEynCygK4lvKAB0vV9Hbq8voEhQDX8hB5xv8Kx8Ozrym0BQ3+VHtdnAbNo
6Taq5EIsJL2G4MWoFzhuUuQsPdMDU4OrAtgaJf642JntFBngqheQs1EY4Okkf9bvlI6mKZOFL/44
pKyyr8aR7+IW6sptnULFVJzqYyUkDsYlFPSNgabs1K0IVHai4MUGdwnbRjHuyaT0id+xqJcx2uMn
15Ct3y4ssZ9sPKMZNzq4hpqM2YkAMWjGcjtHHOe2Jv/ukDepuWww2tG562+vFGartaLJt0tXXagc
xNjYZZxWIfRhQHH0Rks7re5YGNNWhhb3SoDpqT5SGPXir+5XPl6J12fT3K0mc7UYM3QN3l91C5ia
RD0k3Lp+NGAl8P/vnKGkftXWfoauvCRLoq8Y0ZpL1mrtySHPtL/w9z/ftTofkTYPCy9PVs7eTrco
B06QOkmX8hubc1K+OP4r2XfVpEbM1yGnw95xTLEgYmrlLiPSoq8K3c/rIhbn4shJNrvjLEn/rPzz
vg==
`pragma protect end_protected
