// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sB75s37w6XCOK0bqbPah7MCLIJOqH6f9m74YlhQqxF9c3w+syv/yqlsPi0hqCIZI
YiyyBBsx8Sd+qL4tz7RyTeDQUKOvKpn5YYiF+p1l1dPPDpAeLigdlmKRGfz3CXsX
xjerR9qRcuzH5ysKoB556+gM14KV2YRJDcHMBYUxcWY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
ZYLYRRN0YYpvYRXGdT4kNXVCfZIGIJQgXGt6QqCoP1WRpUONPUEYbVCNRLIrgFA1
ewpjjYpJaENW9f38KnrGlMQiWoEBWZY1kIJSCD6IsYAIJsQWRqQfNrhQiIKiEFUV
LEVchCGepqlkyFhx2ayLtoOkRYSvNoOXO76YHcoq0b8bPdDgszESY9er+N89TkAs
6xX3gpbV5cxJsEfYA4SSMlxWZhs1utpI68w6SMqOE9BD6VOKPnsvT8M7q4lGgoB+
5qiuiykTGY7gI8nxfUDsrpMewpBZfCgP/KRHC9q6fctvZ8udZQ+3hkkOhp8poRtC
OqTXa6FnOcasdi2WB++yvq36DmkBGl4GW2ZXlDqd5Mgwcca9VWzjCDDyWr/Csgqg
48JcE417kWkHBhv3KSLN2vkP+JxZWNLRig9L0KijjlRGmMNCsdEAJ1Qv+gJtFbeJ
A/uc0JGchJ6qis5DtHkcC5cFwCYUZcsMIz6y9eW5UeTu4OArTzsShGrTWx4XGeZL
353OYkWP9nY01j0QGqI5qh8634XLt5c7ZbDKjseYlKMBTI64ifdwM8idr0f0QCcB
jGTmmZmpF1hUWjN3D4UebPpW1tOlhSFGV29AgQBJ70351FV4xG459hPTWJo52peB
maY2GzQxFwAxKPqG2iLlg5EnCyaHkJwVV2g7943aGoKnVxUJn5PTI6Rhly0HeMYN
5ob19co2gThZ9hGkfQmctAUhSzuABLTq6Irx1QWT/OlZ8I/CIgW6kKGIMIRnfGt9
81U21R2OOzHJt21lGYwjCl32KEgOMwQXxSgUKdsnrXbfvu2XxU8qADcVWKvMAOep
fCQ7hqKCNeaVT7Ekqjd9fyd2Xoq7BfqzN82WalQQhlBPHc4V4vrvN6q5nQ4z5Pyu
0l5gtYQp5aGVvsrwzt823OwI159LPY6WsRIsznFR10yrKZASdumKFaAumHFlD0sp
wbNv2aCdfkyKt5sSkWMmqKeCwz+EWFbsvauvIS1eYGEgatQp01smZ8E1f4W4MHRC
gRR3HKrTIStckpKIKG6JKTp3VsO/ubMh6d7XyvCKU7eVYCz5bBxQDncRtB0kVAGC
/WehygOzozGMlvnCm/XZDmJdFvUdymrd52WqTqd2MgCvB0BbxkSAGlB6phZ9lmQE
51i0YQ1The37c2supxyHx14r9rwFsJ/v8k0MeOVrwVj4hk3s52xH2vAhPdR3GWGB
bVRdi3YNk7/MFsJIRsDIKJ3qGMwcINjybCGpdrH5maIQC1TzsiLxDW49tSFAyFWX
l9TnnvKM8DjKVSqHXuuZnhEXBqXjnhBxFatu38LwOQ2pVfOJbATdPa39e2gE7Rsk
2yYmy2teGsf/7wMeD9+6f8ciCL3X7MUmY+nHciiu0s+QDKi4zqvbWLYzQYdV6EOC
hljOUO9kCFD2RbguJTRpA/SML55TexyZA5PBroTKmjFaZlyug1wcTAw2jU8LUiXc
F2upqu3k4DS6IoIU7vIleMsxmtmweD5HD8UwpSN8q7Ux/XpJnC3jf1s1Srvvth81
HHt3q60eBp1ZJl1embomX5lnaiwx6jtXKPCPZ7RZoEErbzDu6dcRRzxszJu5owdA
44sPtTVLfDcDoXa9xt1/kNWg8jnf/shxFPHOEdEOVvPLvseuWBxhgcLq6vjUuJ5Z
tFlR9smOOCvDJSkm+yhJz2fNgnu6Z4v4G9uKik/km62+H/jNw4Q0cMD4yKND280e
qy8aVIxebRkaGDT8VRyjHoAmuxzjMJObBKBE6Ha+ny2OHZoKUkHZCv+/FP7Mwlnh
QvGgkNuh6DLSKlj87K7+joPaMruGKBKfi71yo0b3YFrqZbd6eD6RxMlhnGNbYC+b
QDwpe/1gdQDe4UtJMUXB841eoVXuzJSUZKeehvwl3ld/z12/DG57e3rojCL234jI
pOvj5zfnINARLdmo4r7rEi1BN6pAfZ+/rxL2qXChYkKjkPkvzlX/CWW5sD+Mk6ks
DXQltTs7VRCi1g7wVAp2/ftJKv1YZo/7g2sg1aaaoGzyxAdIz8F+Q5LLdSXzU7EZ
VfZgpT3TWgAW/Uj1oSep4Bu+YhuiUTNNSGkhqC6skXJv5c+6CriWIKnarzDBoq92
2cAMFLAw/D76JB0o3bL1teWw4SaKHhMYLWhm+4cDpyVPVprbWJ4e7ef2OGLYcx/r
EMBNHV96eOrCsTpalZB/g9sCAiC7SyCt+GKezDsYwbcILRJo719L9if0urB83p81
2T+FSb9MVMSfTY+BDmuYt6wJT2w7ePXC5EkG3P02g031mdEOrzv2ZhV11KpT4yje
RIWztDk2bK8zi7cH4lo/6HXF7vGcNOyQ67AVbogmqiC/ZipqitxWUcZBmAiV7EcC
T9BWbs3K2Yg3Cwt3sl6Weou+Ukr+2NttEbVLOzv7Wj6S2+ETEsP4LW9JblWbiAMo
4Wq5rIS85hzHtOsuuP/OXImKvkdNbadhaE20ibTa0nS75wCDbxLovEJd8OCUbtfv
KZBwOKtnBVSHEoIZZ6qMuHNzYek37g903SYE30nbeAqxClBaqUKNj+sbKmE6VTGD
CvL5RLuocjKnlHsTtEQ3s4UUGKzIfgvUjLjAqn9CtNC3Qv5s71nroEtjJL3KQBEV
A8ZPA341jMcJk+vfb1GmdLRLoMgQMrb94rr0+AleycWS8AJiP7KuQHKqiG4oZXsx
FZ0YbExovLG869wSgqsBMMnvILTEejrXgKTuXLJGp2P6PH6S/RRe0YyE4hKbDmt6
RFv+MMJp40RL7kdDhDDQA1HMZ58rbbZB4Cy6URPSE7AmeHlYvR00MPCtqq0Q5CYK
gLhAW8HBrz69Ig/iwq36VRpKOOQoIkzALAbukVZ8xWepplCk/BTbS52ubBCNzoZD
vfU8D0//qVDKRH5lnniliTY/QlhKRgQ47txzBW782NCCzhpR0ml47+zX3KMX7mc1
F7PKnPiTbEfX9+aO7d0JwjEkUyP3FxEtAj+pNB19I4FR+sNv/Z3qKiNytDGc1H5I
aGa+ukJvkTCKyz2TmiRdgx9VcG3WtjEC0b6Mh6RGmyHNAAn9J78dLCc/FTbcFbWg
9hIDzMfhZbbyCOsQDI82tAzRpfgMS8V3pouF17GZJQPE3XMCmqzXvf36acCbmeIE
kL4yMgczwf/uZDnyU7Y218w3heKZBdGEljyoq6u3ETnhf+yqR9P2he3FpTgeG4nR
k9TOHp9Nht/TsCwyuGsNUi8a3nu1ZnnhCGwU2J0tmq/k8N47wQcitTEiXY2uorWy
SJOxEef2+qKrXD9HHnUknpxH26d4JuLaMSRah4o7rT3eFquaTJ68L+FKUfDHuYB3
22EUDpWo1lcMgTWuMzBigHd/SCkvWBTHRazx2LcSjVkvirHhq2VLLPcXBTQf2NJz
vSAxMCzXXv+FDNCPjHE6g822jS8t8wshGA4XT2usxp/YRwtFafCKfOiJ1dQja6ED
JyMHdpaBYesQkS+z1nd83ugm8jvCcuQ48vJ5Sr3XlbtnhZdPV6zh6kuzKYbdNttQ
NseLGu4z03fuSFmNb2hUYrH6qv66ziRRL7ruCylyn3JU8U/WpqRgI84dlXWRHbIj
VT9VOm0PgCZlfD8hjxrKTHGBqUNoBRxhUbrBQAc2UW/8VIgpWL8kZ8c81ebw5ZZG
FsuDq7HFnR3ABVC4oDAzf/aW2XiTYxb3y7U5VYgXmhud696VCQsOdausLTvhVGLz
era1Km3YnvwGcoP7dGbHgXkeiuz9rndyMevww3sh/QhN239wxbPX2MgkXHvnfFXx
0OcbbLT9ZSN/MdhXlEbL4c818d/AqDQGPbuO7xCSp8tI3Gr9/xmjKCxCDjxR+5oV
vxDW5Nadt2b9K4kWfjEqpH6oDoBbeXxJhsAiUnHjFrO/XEgo59nMFHxpPRN3YITf
OPL7vA9qMvRCvo6i5r1x85gkzoMRua+KoxchSUHSODZ2KrT1pJj+GuijfW7qRing
IbpVK+0CYywiGaoGiaDTw6sX9reKElBvmfwS1yqAe5SeLpuXluHDGVnAjypM45jH
qIh1R1T/UE8Nn4U4//cFqlJIlwsS29QDrBS9RmhWrOKUW1BKdMePk6bNGOX9CyXc
ELETaXKk+xmHzZTst+c+oC5eMfyRPp3qobVZwwGfMVmZjBQEoZmibGkLSA9vwXHX
eP3fulQSMxMSxAKzjHsMIj/U412EQOR+CPSMU+euSowuuP/CDAh3OEIcpRpmZcSI
vNoMNfO7i1oja6vl+iP7xHEGMaUoOa9v0mJ5NSPMhUL6/Rby4xs+2l91OtkE9FGP
P6mUtqRyGWfQ632VkUPEqwTQs9EG7fSid3kRNkkTEXReMv/VYSZQpNl4KcSL5NCP
ErlBeX2GmOi4+pdA1gNXDMp+Uwu104JCajje3fT6GRmXUSzyaOFhS5W3lBSgphYt
pKn9VH2VhJJTdb7zIoLi4IVP4sdAuI94nyfG98W4i5zkKRRTGpRHU/DDppfCKLAH
lrr8f7YwZiHTZ+upnpW8ZITIPT4sC1gdjidkzpozcSJyaYf6Qgwh8/2RSBhaDh7p
cZsO3PDDdGWtD3OcU8HPV8eshf7blQKJFT+m5P26EFJPrInfxolwhZLXQHtvBGFA
w3vK+gs8S20jD7kV0b1hQc+Uq3NsRiIuAA+gb17a3Iz4yjfPOsIj68SjP2dUd/tF
1l+5CC2/oREe1zg3R32xWdRR7f+8WsuBLebJjAZCzZ8GUqhVB4bshZ+SWQ3uQtiM
DzqE32FF4hdkJh/ybw+CaSPYMCm9Ig2HilswIe8DNirZQgveooZivijSXITPS0RL
b9u22CGF2Oxg1m6AvY/XQrOs4ljecPS1iVnKGE3DjXj60mEZbh3h6HF9cHHSMOnR
5N+axsUe4VT8wknFX5gfGndeNON5Ihnd7zDyCksZLILaVHbwdJ44BKxxNpHRseET
TiqC0KehUyhCOPDIJy3DuWF8q806skQlBJCguXl+Yp947sQLewNXhPiBdZCf+yRU
oLIZfpbxEpDpc9K8oIiLl0auRixrJsXqdHBALWmm93vGto3LCniikzkupAcJlDn8
itxLLz6SBtdZVHM8fAWL7iNFzEi+Dp4BAkJW6BlruUZ++zu01KTdJm52zU9eT9D6
kAmQVdzPec7WZYo6/ZWwNaNEO9B4UJffdfNLLx7uemiBHjI4pWNnLvXR4rQNXzP3
R5MMUQrKVquTs090thD+PMzn4F3JvJ9DdaPGZnlLPQHYLQBjVP/rlODAtdeTRaYm
r0AJ1AvKnYmNG4DoLwPonUw75mfKQlwgD4qfqm9MqL6z3p0hO5oyuyh4wNk3hgtA
D0rFSTnIajPiMNeqIMIGcPN42nValy+9tp0h4L7LITkWmn8CW2vKecbudPSsGujl
PEsP2L6Bl5+aYfRIhKV9VaP0T2hHYiPNN9kWI87pDfbMOb0BJ3DSd+9uHUvJ4gQI
FkKuerxJisOxGdviVCmIXIa3Nc7GxvROOv37b4fUHTKfLF9qwwINi2V6eXBfQkla
Mjdw9rA17wsNfMunNiKY5op0zogQhnuLOh4Hqeil12Ah6OCmJYRI3tnoxg8l8AnK
wroa7rr+tPgGdt5i83qTtVwcthwd05CJuKdx6gjTtJ03W8d/vgcS56p5cS45Zqk5
L/tfELKFxFIEoF2WBuctOq8EXq5L0lrbcdqaDvmA7lTCTi8/RjBoCBIbGgfv4bk8
NmSOc5D5AtRkRtNsAnDTu0PJotgkQe+8CoHRnWlHSSxdD40DtSTvdB2x8UXiAq6n
HEa0kXO89iiAaSUq7oADB+UWDZ1sOHhtsr8MPJo2wBdSzJE56Ct6KiAayg2KvPhk
e9q8qqAz3KInJcKLbhgxx8Dk0eGfpBW9hODekboV9Gt+o8Yde8/DysmO56Dd8AuR
P8bxhdGxysrm7X37Ol7hfQuEfLmBXqrnR+I5PK9bD1+/fCNvGUINm5wABDTQY3S6
mBqxqhuZaRHKxvU5MxBgTXPR6jiIP5QuIzZSsZBgjoyZULFSfhAWzOQCKgYjYhEo
1mc9yMiNoqQGYi9G13ygaqGgbI1MJboOxBLNwO341PPFgzNXPne0y+AYXsTUkaKp
cNDJuovsQF8do1o9Ghs7qQqAfWEcmjp3rDrS0PJP1f9ymbfyQwSnBJUfXyrsZP5w
FQmxV2XzTWJgoOPBI8Uza7R58EbjjKAjaogWKUByeuXhMu+sRHYykM3Me6sqpqi5
5gBWNOJB2E1dpkGmT1MkkRIOpEuCrhzljDyNGsL9whI5KNqElxU+v5c9UFn5CIS1
CqMAvvdQtTwptY2s2dPA79y6m9+1gLxleEd1ulsUeUznr6UiwMklqtMeKe7PYtqa
kKA60LqOZkvV7Z7lHmEpV2lnum9iHlRRGEvqvlBd+N2V/j6WOUK3aDkCHbXTPjXq
2BjM27j9A5PT7pv4r45lfkV3Cf3/SS2ZvDfaQPjBSH/oPNvlGx0s+UBPWVPFqkQ/
THijIvQvKlqGIONxVhcVKWfhfgfyqjrmT7DIRwVJ1+ybypAlf8+7chyv4CB7iu+G
p5N9XCeXDP4ZsLB9S6CQiOfk7zecB0o0vaZaLZT+cB7U6noOIrhV/xHVnJjJ+ke0
va2QnV4yn8qbkXzET61uxUq8Zh73uvZXgdZ/lsmQ4BQR02Vc3sZNoaBifrVfO3GL
NYNZ5EAB66Fjx1pAQUmps99msvJX0hg5scPRRed5gpfFU+762OV71hV94NRSEbvf
dH/0vFJY0HDQIbUWkZppBctOPHYiz/ou2+ovxLoZwLvEbEyXdZn3xYyI/aoOeUG9
Fmu/HnODT0QFyfq9ocVeFa7lXT6mxhPLPcYZVUnK4QbXgxztRIpNVm+koh2fQuzC
XVba0VLS3XBE8/+XgtKE48EcaNUPBjYskgimyfL15DfIOMu6TZUW/fFDDmz0k1fM
F1JimWXI5QcgHcd8TQ+Js6EOCxKzbkZwV2mSctsLLzWTBjLvvfOp0FUfalbcDSaz
QgIluE6dhGLEw5tASqNhkQfYMupCZjIaMI/+SyQcPMX6w21PlB521BGqHw4CINNW
HjgqUA3KNTFIVA8i41nJZBgElQIZ48m+i9xvC2mMQUS7UkKdBamVA8/r9PlSy0W+
MLhGlR7ugQ/d6Egz1CvrnpwMqClK9l+OEFQc8J+oZcYsSCf45uPyvos0henykFB3
yMXhNgBvGNsxOVBr+t4v6QioP7VX8RwXskvvzHd4a8qcgR8vLng/GbG6BMEBxGJo
43OvBtE1SYSJNkl6qnHiPhwJnlfwc+XXR0AMI2GHLR4fpYKQRqra138aPdyrnH3H
06GoxhmebuALs9oHQkIMZm1llSCKOCmLA2OoWvXN5TcHRQC/2Fpa0hrjA7DigSZy
1VR/n+NkWbCaGGVsjanRCUgbEHQUnw9RzQIW0cvhUC06DAR/ojwVgKGZkVZ0wYKV
KIzQFFJthxEC79kVbbonfzQdRYbtDDWP0mV4A0b/96xTGowDoAQWeCc/uYqO0trO
UgquWW6Xy4dnIj2wsicudsMx3JQPW1a8trK9hAeSQ0SWfUF8mUFWAyCJWwekCUpv
EjQLlHIMzGQntqaWIRP65U9m4oK20wAfAMDcLQi9wTA=
`pragma protect end_protected
