// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R7v24r9u1ctqogwGyVohHaT0JjT64mJ/Ef6b0kSHN3d4FDxLhrgCpmy55EZxDdHB
OkedqDs8aEbqZfaRxz5aPgDmL/EiKC/ZtoKWFtmd+iorB4VVrojI/nzSavp0CiA8
QUkjow943QWuy4VfxL8pCf4YpkFefWXkGoT+KtYe1ZI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9744)
ET3yHJKr4P1lzWS3sp4N6ijzpX+63T9TSluZLX1c9h7mlWRHd2lIK39VTzrHxYCm
3Bo8pV4ipc9vWyyfjwxJB0odK4J8vuVzzbghKSvEmGjGs+eNI6DYqml7RHkGYdvx
pHWkS+KyqJRgWOxFS7dh3X2f5PhJiXuSwikQyfn2QvwPGdyvj/Yyoz91SkaXPELi
+GAVlrVP7FMD4Pze22dQuuAEGBndDT1QwOmstE3reMUK5a4gl6kOf2Yxa1a4wyGI
c0e61e3Xpsn4m2zwN8fSzMVvKJe0ca2j2Ty+LZ5QJvpsDZMI3PWKhB4LtEP28nhj
MN7PQSWWgKhDLVaFXsisU7hAtJu5kqnOg1x4U9YT5chT4vueJTC0rF9wCSih/O8w
70ImbwU9VwZwH1QNRgQ2gHSltU/gIRzIPx69nZEBnoXkrNqS4HuO6tov4OTIJ9vm
YVhi4A4hv3GTZAfUgtVM4C7JiCfpWTXttniDFsjilbNeT7SUUuNg9vs2/sj9fWOl
uk904C2QNKtTtwPebl5+4HMODd98v797dn9A6GnI5d++iavRLxcscGggB1D/94TP
ZEI26Ee6RXzfFBoUBh4mdACV0eStCr3cgZczz1pICBFw1vvf5Htdt9NPrjbAE6OY
bxDzSrw1h/+f9t161vrUza+gS7Yy7g9yViOMHyz+XqO92zDLVxbdI6b3y0BYkZhC
/jHz49pIt6BE/6JH26pyVKv+/P2Fu01m/wbtWoE00752C4hZ0u0mCTwqTJLoV5i0
Icna9SvLvhZ1zNduL79PlPb5hO6zUEXc1Lw08pZEAntWtQWCZ+h3aMq9OW4HdZON
uc1hfHxIH/MA4ffTm0izguohUW5yiZ6uVgM0vPCjp2mWCuNBai4mzDL294YLmKfZ
hGEDN2NzgYtw4CjmGqtfW3CUrB4oYuWqsPq6ma75iR5VUE2btegrU8FOtL3ziu0N
RivJxeBhAms+TBcvQDdq7xMvzbydbM6sp88DCVCO0Lf/X7nEDwPygeIpSuJhFtmD
ZmP++wRG0tyn183aNlp7P+CZ6D6sAu2me9AXqCtsWcNfR66X8m5nm2LylcAx/I+B
WSZU2EOUOmZqAYmKyTHruqdsps+1yyTnAQqSyG8OS83OlhRPkfmD0Pjlix7KxVl/
kuFVoaN7gROx2y7mmpyW31tmxBiSmW4SzOD5AJxSCXepu8iawEi/WmAO/1P6cLTu
KPf2b3JK3QuUWcmNxX5BmuIg3sSE1dsbbZtCi736LmXM35mhLky7DMhl3qdr6SDC
3bzYXebJIrgBRE9++r3enyZb2Y8+VEBhm4ETdsoo8rsAcGrffcZbWnqUCezWePdt
qEYjDPKLMsmeKN5lxvwnGCTnmFLOzl+rhkcJkumfNu2kPwTPdk0Sw+i5o6rvKZkL
ibEr3TtyDqs9a0BwZjsnRwyfCzgbkm1Y+u2rF1oLmKKfxc2QmJBQZD5t952tZG8K
kjzvl3clLP3CZhzn7qGhW7VsG3EJXJN74Z32WNRHND9yPZHiRtLglHAXXSeHP38y
en059nH1/QM3DTa9lrVf7UAXq2vsQ2XTnz+dYkBrLneLZQv3DuOCB31lBhzt1LuG
Ex2SXuOQkjFV2b5Qn0lz4Ey6yhZpFBc7CKrKh4WhNNbguwz8Fj7/ZHNKdcwejv6S
QeQ/6DuoR6ORNDw3dVkRJh4pWEMRXAtoh/+QuZ91I+nXmALQh/4jiVDgb029lxU6
4osHD6bBlvfJAydOrqUz+vYAOp3VInrPepOwe1mQPKQHc+3u8d5HUkHfzG5F/HIp
dL6IxSbZwtG0OydcB7Ammwzcn+PbFdEo9FGdHO27+//wDMlWu+X0yHhwZTybnpl2
3bqRlnFOjmXAxK9pgL3gda3DKrP3DVmiju6zH8YldkIuAmVFrrSpbRkwJ48xNRMv
Kvi0Qr+QYWdtdjCf66XoMC0bPR/Cd/34khpHvv9iYfWwr4FIuZYcWJ6XROMVSk1g
oJxJXqdqTe0smyaZ1EZVavrY0IGZNT3JGDqv5tEyxKAcseSqplHQhkkGQZ51xiXP
zaVz9VJWjk4ZvWcJyBNLozTy0U/80QkkfwIgQ/ZhzeSdVT+Cz/T3iGnp194uQj9B
+ef4BrszdTucFmODEJfbBWQb5b1eEaVQOQWrdQVPOKtIdMgGM1kZCqqc8mU3GUOl
iF01P38LzPyPqVqXOk4jRMFV2+RZ9KgS+4lYWsZnVGa6JhvDyWZg8Y8Jyz8QsVdN
6iKNhmYNKNzGalNqpB7gYfWrN6756t7Jh2zclFDlUl5TNySRtaWnwxte/jjONk6C
ASSwJTF16m7ytKbvmQJjOA2yryfhC9MgkqtYn+vNOdb5Ui1LT85Bv18aZJvoca4k
GmrBDGkHQkRsTe1cMUXexax3He2uZTtgNbCR5oEAQ7Nu0v6eypGl/Q96eI4vQ9xy
Jn7umP7R/ND3zEm9xqUcdYR20sJiaMdvPriu6UH+STb1TrjivXcO8HqPLY+zRy5J
n9/Nrje+zKTefIXIKoA5hgu8JKqNtBomloWXkzmnuuetxWMTqfNSRf3pZQQJ2fOA
FveaYy6Akc2MXUpxbT90wHXyyD7sIDaor1sdU/GUeON3qz+wMsUBvQZImM8Gpd4R
6NTXlYbZHGclfZagFAseC6gIbHlyg7czigaLTs6oQtgkLDMXwgZKquWwI2NANgkz
FYR70nJHHMCX7pl0Xv2aw4y62oTd4noWcoPSd2Kp1ucQTzxd3bhddPn0g+hBeS3I
iGXfG3pxlKwouxrSicnOe6fYqet63xzJBPVEhohCWRCqVtMvg7/2Jdo4FISejGhd
EhxnZVFLhaFRXiCxGGruM/agsDcll9V6MWYgMchyTmKr9POKCoMZOEzgiTgcqjah
w8CwR4YmS2lu/wvqDAnr+wVpTOdDR9Z7l3NwLcrI+sU8fwgRBIGby3CKMpulK+vN
Da/CQ+7kTeIEyvA4OuOzU19+gV1i9TmpEJxPzhPsLY0pS7yFzN54H/ha87uxwSV4
71tdCqWFEHHwjT2ggOAx1vCJmj6t7i2ozxMfwexmibEhuaYl4tGB/4UuFQa/RQbe
cVzQ5+pLb8Z2i4SXpxXWhB7MvT4gQa7xwIYBV531FARzm/IdeMfMcjCOvrNO/8J4
xQiSQ+zumwiVCT2tA/IRRnyNlF3mx45D/48p0ljjAEh0eANvVWTQuTIJnLTX9/V6
/4FXvbCaJNP/gR/FlwqavVQ/QhgVu6YVcPrcnMx1Mr32kY6MhSPf6B7nK9W585kt
xg53swev6EJOtv7EGL/6E85DKCsefk6KRfL0wHwSHaNHy3ufqw4nCUdSmwrSKRML
KVxdhZJk57/Z8FLlk0vmT60J55vt69qIhmJQjG15WnjcT2wPK/DECA3xybHObgvf
X9JXXvbwtIyFL9UfDQSTzSY2j1iTDbPJJaDG3j2zpR4HFYRK02Fe9ivg8ydYLt09
TEGwNJzQq4726JC0lSczl7XuSaDOXlBHCpyhv7mMrAzIlSNo6vJjqLS2UAJw5mYU
AVCpVKFGyzS8+rglK0MdzGRThtBTQ7oD1BW4QqxLs77tbOFJqa/z0Qi3aEUC5TDP
pUGzc3em94peyJf13lUdYRUDffgKsNAH9S6cHHzMuPu4o8HVF3Nz6T5s9UIejyXj
w/KBAc4CnHmFx8OorSSOYhNwYecixCaB2Fzhy+4yl2w3Xs22/uI1nCedZtnTnzDB
tfXo28uOl/far0GpOCPgv6IDNWmSs/X0TZ9ZcqTOBjs05H5F9CbMo3+O3z/bDpuH
TOlr7/8V6FXvrP106YYbVFjbiNjP0XrqTNlC6pBRkxKrH7na+3lXCI3aLG8lcJfK
6TSlYFJuV/QqaeHuLKv+O30OPjQxKDK9+j7FrN0+4bky0hxWJ/vuKNGXCxYQRPju
Cy2FppyLEUfuP6inbYRJ7YLdRvqYwmXMoY06dvdQpl6vLcw4Wl6rtNoN++UE3xEi
Z5UrfgRZSn+Md3idpHr5uiaALxkUJDO6n77yzWu0wBFZL2IzggBrc2nU9gL2ayFa
KntQDmKd9HlaFiYuq1dSiXnn2zrgLmbxbf8mIfTNSPakAZBVYTCOaWWwsoCiaSmt
oY/j9CzUHC4o/N/ron6CToBtUbA++SskAVwLDYL+yA4mbQloZ5no9c/d99RBH84W
9Yy/bsDSyWfD8edazzBtlXM5N8qHBXskLnrizNIvU+iJMl5dx9rRDkNZSn6TdvQs
k7XS/YGjIvW4gTGYYUdW5wI6KumdidSnS+TgW5WPxXpNkOKWcPhYxqGtWYEK4v+K
/UW759RgzoJrDNinkxHT7wGicLC0vGABclsw45001vhfDaV7FAKtJY/HvAZIaoRO
CJY2UPPRUCV1CPjQ3vLCtZzQb2FbtPyCAedhh4ZUNIoYy1/qApz36dvUQFyMwLm9
L0jvfaPBtbmawJod6dz0n4+riUU5bTpbGccyUFlPK4Gf/cw9fuVZD4ZDuLJ5My95
q9JChe6uo/16odThyfF8Hc87c3+kIZNnOHJjk1lSuY8e5JLIP4pM1YOhUc7Y9MG+
d/5gALxthR4Iif9L+qtTRoIMvAvYy9zRJJnYE3EwLMtVDgsrDkwJSxAJG3siu4ai
T1/OGpSitCDnAJc8SJNjiIjLIR7c6kIoWYJhWUERoxNIdI1YRftQZjnMjLSeRNEy
j2NxT1RZlJ2vK0S6bkXEjby5qPWT3uPnYwKBkVyMuSoMaVDpE6jMWxYnxl05FbJv
YetJ8Yo0LkIoe9lxU3Hs36VTJcpJZOwTqR84EgcCzMvQPiCHJNxRvE1l7irdMaGb
4zyrVh38uzNUwf1gitMqfGsIdsrECZQE76wRLls7l/+laPeWwTcFCTXQcf55Fq1i
7ChlMeGXtr6dJqOgToi26JPbT2I2TE5BvrWYPG7zaFL4y7QyXSK8XPSycDt1v3jY
nXjBjGOgjaxH6FJ5Ej0dyuAK+7kYJcLmtN0QkRFWmcnDgcfRnvmoYM/aapJ5Hckd
ABmcf1rhr8vEPGDiLQ12MBu7vkRdsZfTO2KJeNQ83jqsATJNLXpcAqYExTbD/sgx
5EAVqak9uvph75GZC/iprwRFblaEcl9Fs1lR3jySkcEuWAYDaBvwD4/Fj18wXjMJ
UUxYFqGgXQLuniioTMRpjZA9Kl4ftaMFDqCIFc0KRXYWX2LgUh3iv/5VTSO3XDoH
O/fXXN4lTKZttrW1Z1QIgxAG22m1u2jR4Nac5vjpXIfgvVRhcHWPw72YgcJfImYW
1dXUGIutxe8AHHG2NniXzgcU7TOI66ePz+OC/un+UozEVssgqP9nq3fENJ89EWW4
PsYa1jRSUxx9gX4JxMdJqQPTAtsYHB+L3WuNMYZtW4YG8gh4hjApCVU1FfXDQhIu
Qz5kKBG5oUY03HFPgFFh2ctVxybD2dauSFOWcaAU4at9fkAjFB6BWd+6t0LdCxBW
CRyxYs8KVuuZXBgTvpxR1uHyL8pQvf1oTfTPOcOLY6zLQdHCx177i6Z45y9Imnqo
UEjAKGiH7WW3PzWHNkExAsd5EsrC/tthlfmPq2o8xFvETgHPH3t7NOASSeJP3okg
Jg0/J5lrRoHUbxlJBdjgHfLLKxMyizHTQcRqCx91etSnigNFjAIy4Vkyd42J2VUN
O149JgYrbCJ1IRliEsbWku8F2ozuB0A660UcxZKaHoWRCw+n/gHg0Ni33uT5eeqx
lu5M91TcnrUjvckgmFSB9O2gl6UMuNpmWdO8QtgPp0uH402rqdZ16AxX9JYRKfGV
P9yceUerGGsbi2Hab8Gdx8y4GPZKAEqH4hEAM25QYK3HrsdJlk0KSN4fe+HTN8Kh
6Feo3gOYf5QTpOWQMnMgu1N9b4M64AMkW9tc+NR6hJkHVskJrqpfdTq/rrgaex50
wDz3VmipgiwifKng9sw/fJpFSDlQWBhGlUux3vII9gVdnULToVAL63Yyq4cF+zOM
vmeiVl0Ok0KU5mTgUBFg2DP28SvqElXzq/+0fmJt/U5rUmW/a5HH7yDE0cbOiAYP
YZxsdvQDU06jjV2z8Xu+SNLBaYMJ5HL7usNqKrVW9x/3cvT3xkMlSHW+etu7nMs+
C9lURv8tksO3v+bvus3QFH6skVohGH++ZY3GHNJFLBbJHZRWaWlvLJubNmC89VJF
WowLc9SyL5ENuSqVoCKFJ6J2Je+wEk+sKTHPJin+u8DaODnLdt2a+ZyiMbujQBuM
z1GQR2bFjdOwGGDGh2b517udXbsrgncnBNdGsypW/oSNDdE9JKsgEKrbL3Dp8Nay
dDRLE1bdB6qNkhbW7J0VbMafJH5WsHgM68Midgaxkik7YIQTu1CuknAqVTsT/ixA
FpkEeAFsx7G+0NxYkpzEjGKAzKmAjFGctEsgW7n5uOED8qDt7nu7srCLlZn2ongt
6sPKtxPKiZMsUnvOdr++EvqI7w0KsYFXLXxi/rh7/z07ZA/uSl9sLHR4xuqlfMxb
lxZ+LArG9Wq7cruDqrdgKM5MtUP4OjpyenbAABEIrIe39asYMqX3eItUxLZCaz/b
yJe4/KI78Xb7EfjVtAK5h50XwRWXEhtn6sAhCM0g6f7hh458d847APRBLCeYbhaq
s1gKw0vb8oqXYNmBUeLwL5yL+F0TXtwchHLpcV/1U2irf1IRXoDuyaqauXTAf2wZ
Vn5IX/TYq8XY4TJkOzi9RHZxyPmSdqmGIW2M28nnz+J9pBAliLEG/QiRf3MiiQhf
Ww9Z2njT+wuSh4beKHtVZZCFWZJqb/8K8faXjHF1pzNBFaxoKfLoI3JgG6LP1NvA
fgRqfwqHDBrs+7qw9uohtFOkWvjE0xjygX5q3AvO/klgKfn7DJQDqxFNVLMtolzl
Q0P6vVbCDZ9qOcallU8thyGBFXCyLyVRzLE/So4Z9KbMUT5AwJIaSR9/6v2AlAEk
irJ8wwVLpYyd/P8jmVFKqh8KCo9b1xS46IcuQ71oTaLL8hPp73kUvAuaXKeUfXVE
8npKv3CNUlriho5ODPKmFX8AX6Qm+NqgoDbLhO2AXMgaOVd2iDhhksC/df6zhzof
osFNUE30MC3D7yXJbk+Cdu+WYjpL3x9ou5ioyr4Bf2cIn1XtOImIf7uClemH+mSg
Ve3vZxQdMdN1u5nHbnB/cVMjK4YQ2CUBsLmG1wRZl+Ftip1YKtOrlt7Xq2ii/jXT
9kYhyYO1EjagoMRvpVeC1wuPwcOqtx/aDAU2wUCbAXpCl5i51intSE9ooJaFXnrA
3d+aI+W8KpfnXML3J96AOOGYzhBecy6loYqMrEw40etfWB86sKrkt4bMqnrD2SIJ
66JUehyqghKhoghTBQ2+H9PA9pnpSuXeOQmRELzdPe+C/qsCJ/lc5A0BULUS5YIm
5vgVZaJxcnDlIrQ5NdpKQycCcs13twkCWgy0RbDzqXMYBz4zZHUUB3yiwj1njPMp
egbB9XKNelvkjlp13N0yl5vAmrsqYNBUY/qWNyPitfBSFvpFwfR4+Dza200N+VZq
FwhdEg6yUxG2nkA+xbOIyNYukgVypL10C9QRYHOqTKLIibxoPDtPyo7m8gfF4WVk
Y4yyMMKmdWO3XT44CoubSo1JQIp83x9Nr2qd9SwLBUpyL1/UVtmxo98pVSY4IAJl
qvXZ6rJDKdlTUQy1pXXQa4kw5s3D8TIxIUMB4M4zcTt1XoRqOnmnq6p6rbmAbMrR
GDeYpmKKBysYkYboKreLP/TtfHt5VAInz+XlefmxlLehlWAUH55+DVaYMCmn0loo
sseNBlJFcKFzfSpjNHPya2n0PH6H/xsd5qVRZJxBKTWl5VK+gFgxhqi6dVWe8vt0
3XGymH1lXedFUt8k2WtEd3xRwR7S9TcH3oFigRSzMRvEouKJLo2+Pgs5xW2eoLuk
Ums71jyG2YHZftWEo6L0lUr8PtNrQV5Rfq8KaccWKMaQPF8g/LJ1n+BQ9ka+gyhr
0HyY227gNokC9C+oD/ujpSq4mLDI2aQPNXpy1sXgpHrKPZpVbMsqWfltT4+qAPIc
eMFZxGqckmQ18sfsB1DjDhcLX5wD8o5vzVE+slkTTX8Qalbk9kt4Dht9xzT8jH3T
wH89m4rNgmuhoBt/T2muDuKxY/7Fg3rJSxBnm29kKfavNM0Q640tuvZpmZm7NGpS
K6O6SbDz87YmBwGS/5kj4Wh0MldUs2Z6nn1LNOJ4zcZ1W0Wo13DE7NXcIpj7ufRP
k2hkh4KK6vFHpIgd7PaUE6kbh8VcVA+nwc0XdwGsxvR9BFg3y9vC0gTUVIwiSRv8
WxAIpTFuLwKaaRE9eOEuqopFuybYYCQA6Y6HKIU8+xcVo/hXZPwuBqgWikuTJtWW
oweU1DwU2UXLVvJQ59dF4ntr3IrwsB9IQ31K2gsnE0G0J+znPh6zK9C3Z28IpnCC
YqaWY8Qd2zUmxQOIhA30Eflf0UotdZBJ3+xxoEp1cm9ap04EkDGLzWqcFxMbjSQz
hD6i9+MvayqDmqsgtjGikIgprFYg1IKJRxMgA8abuiVmDjoxFiTwCddOaY8DUyLJ
XSqJjQQAAbLhI0HhEA9hQ9KJ4DKqPPKXFASSg15dIwHuexcHqDB2OOuhPwBMIoIZ
gEHZ7SBS7r9xSc1E5+LWWHcv7vVMJ2GfeUaP7y7iV2uctmhJTDu1U2TDsAmiIQOa
byxQnstBOZfYGNclAOCJnqxK4Q0Mbo+/ZD1MWAdjs2C4GoR1zGMSNxMAtgNeqZmB
LwDmmxDIYFfXkz4af6lx+N1mGvOCci7Ld7ly5QT0Jr9GNr/ZK2NeGkhDUvgnhG8S
4nEglmD3B1p62h612N1lDlSnEr2OBWurEIC+2njKQdWIzYSvIStXXDfbB6n4sQps
JKgWMoOAjqHdUCtXv97WtyeNokPgFRZ2IRCS5Ms2GolyODwT/Ts0HgL0qHx/ua2/
j4JV0PEURPkaTQs5g/TDPl/yL8t4IyxDqkJSCMMJIMhDE33f7tlxzBLydmw3dNJo
EsVf9jSgzT784EmI6m6lEHaN3mxmOqGjKfq7KxBx0L04KhNO1O7ja1rw/T/E5Xfk
/HuzwA0j3CCTYRlKv6UPdnXslqS3A0q5hC2ktJ/HRdMx0Khf3DYoaGYZvWbQY0/M
XXJtV95tWmrf0AZX5FNrCgtPnmJr9+iY7s3/FOKaMu9M1K3IicPoVCgbB5Tp8jB/
qR9InTtQsmNt80C4pWt0Ab5PRiosk/ei/lxCoWyqBfO9TKENyIOFY4lFtg2VVWXB
j36G2CSNDS8cjHCMEWYOZHZetYL2uBXF1rfTJel97QWFf118NpCqGfI7EGJ68qW6
wohA2iKkT6Bs/vM8+rIw/nebCrYs8oHeiOyh7DrrdayPNw4D6pXvLYSAivxE5Iq5
d0JBt9xJSn3JmlWJK0JDnR6rC5JC7+UxMDW6dNc/ToCk+Qol00zCi/D+Sx7Mz5ml
+Ltsg3bfiDQuITWx2fYkeXJGEpvYYz1C4+a9RE0EPAr6Fx7f4ewwly6DldNk8Qpf
qmlEnbMO5K522yoFjNeR4OZxuEXWpxxdkd/2CFglWnjV6t970+82zd/GiNw5Mf5A
HDjCIDSMnKDdrkELsUqnhl71VnPxNe4A+lM9uHDFB+njRU71gjJ3rfeaEz2DjuaO
j1EIi1x9/Ha2Xk6AIkbwser5El1jcgQhvUb/lbENscYniEY3SGmoj87Zr0AzokzA
gay0TgKgMvOj5eWZ6vwYmXfksZ/fip8yp39JiAoaXkycH1wM5EYWgedoCDHI4ZTq
EBOhC8mFbXF4Gvk4toywSAtDYaBxmiRi0oXB+bPgDGjiq6zDQExn/UXpUrt2z2Ea
PotFQNIjC6P4MYYWmU1FS4A2CFVsxSAqL72846OtzjAIW/wYaLbAnQujRTDXHGvC
22uQmRcFfBW2fjXuDowYhGu/ZMfN7fIzW/Ubvo7NoOKdv7e84QQLY2Fap01Hm3AZ
Czqicg6eetD+NlV7Bw9QQRCdiki8rkBnmOoLuU7h63E9F0XhIoOyc20nS2RtidCY
X3GGu7pcWLUqcorlh+8eNgek/SLQ5fd/QAwWoOX8EmvXbVXqFu65xL4mFS/A4DIk
y4ZcveIRue15Cv/Vo7S1z7r3hscvwNNS0e+cB9gp9xK8wi5gexmSZVJsTx8uhsdz
1qU20TzZQWs8YvaaRkZrLSKI3BFwadylBeriyybHbxUVj+yWsLOxlKCBZfVjxX51
uWxVFeH6q3feVNqUflg+wtxCaPY7gOMwUQ1U7EYKhqEZhNgTziz/M8Hvk01N+bW0
8gD1sSAoaC/GO9Tf8Kx09UVG0IuXdGM+EFpKlHggj/5eitMAT+vlnk2hzskKHj+u
DgPuyB44RQlaX+n+y9Wfda9G1rlJoRyDgvOXOLGph3yK/ozIHpXdzjk8lu0sBX+b
xVDDsqpeEtSfx5yjfkNM5FgU/S5GLzEL67d3ZJba2eH5+py6+dhqqADebwlSAu/b
oeZGaMWjGqcpCED36zqmvktKUBsk1uW+iGmM9OE3LIvZ9F2ZgdVqyVWkmTLgZgsh
1DZOqkstTndaVyzfqcMdW3908BQHqIKpkC5jqBCJZA1FLd/0H3nRq8AyLPLXgXMF
Vkri2zNPLsj1mSdsNqeZPTOJSe0lf5Hz2KYHUIWgfNzEkDJiyGGgbt3FboxvsShk
CtzL9ZVd79K0m/u9IIqCpyH+HNZG1enW0/duaV+ezc0bI8+AH6ReensuLav6CvhZ
chV4dgxma5u6k0/ZHks5IFY8t9Wp2IMSPrudcHjHLJULDwXlt1ntS4QL9aXa1bL4
VnUNy5vp+P7DnnhNx5kAFCwOyB5sX75qEwYutHbjOtIoGzMKfAjdE3ELLQXLkeaZ
+oN3lpg8YHwMYLejQ4eUPMnBidXXah7zdf2Zu3eR9/bg1cmJa+AwmJT93/glnnI0
EK2DmZJjWulWh7EaZGyqZqSF8xffjavtkYNPTbBya2pHrOiIQfAnKZqAm+AKPQi7
YI1DOXFnE2UYKDYL5qJ8x3RByIfmwvr0zpjz6Yb6f/vY1AVD773xja0I4cFt3AG7
5FY33m9WK4ASHqEvj8K2H8yj/uWrFqU5mruxF+GmG6czusEphzg1O9iJtTQO7JPz
1udTy10GsDMurJH/HSwuDJ0rWxbCG9P5orFIPG3X9fgpTd5I9kNBI5jiSATg+r10
v4g16pYbOM+HI04R2AJw26E5vEEu555LATBAXkroLPHQDQMsPXCOeUrkqYiLuzMY
dc0NkwlweOqua2n1ICKCUWmu1k4+IJjdgoCCZY4vjs/EBbI8QIcZyt9saWErKMWj
o5tWNbQBNxBtlIXrQQbC8IrbeLIyXngF8S+d5/zAaWdyvxAYQXOJkHxopTlj4pYG
P+vhXzkO066w/TJv2MS9PBC0buTzed1NmIcXxZm3UWHnCY+JLR5nJXQQ7KH5jpz3
HftgAUNS96A21oiVB4bwpyaRsaF0hGC3RTlFblg3ymfwVbfAkp1P0CIKiLhxf+UB
12WjboA3orVY1hyJUujTx7ONuZn86eJ/Asz/OYIoREuVBHzms5EsHKyvRQ0Hfz0v
l3efBdjRGnkYseg0PipB7U+/8agm1Qn77ptY21e7A7cpeALduEcuUGN9T43ALg+o
SPiJRXq7EP7/5t6cMBvTj8dbFQpkSVB4anxsytoz+4K0CBnnfoLT3/346EFdu++S
NY/g7q638aDPHIWpRb8qBZ5640/ES52czoa+GiLyEm7RrUNRZ5DDLdFsgOC9V+nf
YEz1TnxCPl9oh+/+WjAYByvSPz99B+BctR0oXXD5NYlAGvmvw8hCpMbjcFkRJuPz
KLtgb6oAh0nE7Op328dPpfrOvC4J2r4KtWnXqI7H18IwrVZBWEiw1dmvNQK93I20
kIlu7lA67vlHFNnFG2ecsiPlX4hVrpGjBK/B3dN8G1kgbuUh7ng2PvjU0Crx8ZaV
fdSS3rDtn5UGxBrgh9jNhjXI0ayDQu8uKTlnbVmnQX1LlbLJv6SEHqhkjZ0FP2GJ
3BgdMw3+UBYVgKGJ/Wh0ruVlPgyyov+738Puh6yWuC7ONMYB7VpL2mKxfrhM3CK7
8O9kROZawAuVASVDrx58vmEYIxXNhroP8p88OY15JSQ6o9DremVb2+J+5Xw6NTs8
1dnrb3Z8AROMG0uaKAs1iC1MeiBHZWeA0bxOKdt0b4i5ET2K6ngM2r0GQqrD154q
LFZITO9wuduXBcZKorXp08SMF+V9RvkoyZCSgJm7WazTltqEiRrUArfgFAcpQUer
slmcMaV+TYxFlM5UzrvXhr6fj7dY9btjOAPMyIN9Nbm0wtbgU/4LdrXu9XTsD2ZF
Kbwwj2BPQkxcy6IW9vZe9gcphaLUQ6LPG+36jsbxFs9pdogKkzNOr3VicrJTfV29
hDV48cc9Aie3TpFO13fwdCvG0HbNT6D9y1xIzYG7RSAQCLp3vw/eCiF4PZGCueJQ
Lxl0LADgWp0UCGgWLlhjAnZrMsl26ld1ZvLnNYlarsTCO+LG+pJdzON5Ek4izQbC
u10ElCl9IxVLsBm1OwKkXxHTmCg8rEk22JlPcZnXj5t6n6XNS709zh7DJPnUvEvq
3sgujEqNXL+E5wLmOpQx6Ldg77uPkmdFNP2BMg4AO61ppDcWRiXSsrRm947QFNqk
CK30puwapoPdJoS1iexVJJnrtCGlAVJvPNvPCQHT1uT78aRd99Uwe8MWgYa8b5db
drRMhafrdNKQwpsHCe+SidKBgxA47DWHHfK2k5MDNhF2Wbh5n6ldZ/PQOjniRiLA
IxYyJHSskXjYqrQqme/fnc6kyNaokgBCxLsDgJ6vMLaXxCLdqoBcnLWgd/kXsGhy
2dDMyUVA9mG7wMx3atxM4e+EUdrR1xEwFTMt58CGjMk/w6S0F3/t+HaXIBJcTP5z
TkOfCgvwdJe/GvI43D01EYt9oBrS5Wj+KsbqdtA/SbJ6w4Hm6u239pAgkHQmUrXi
abv/bepN7+isrIDrq8MP+T1x86/Q9oPzpLNWrz1EAG6ObQUlERvjzpxa0+KukxFo
`pragma protect end_protected
