// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Gj4cbz7m832K8JPuLz4fXDSboTxIM/fwgRZ5Lx0Y70qE0ciYhymA0LE2M2D/I9zu
x3raTX7h+J5X7dKjqqyrYQEHab8eSijmdyrpvfVhYDgLnLJnWbOe2ozoG/RGqYaa
avqFqsOybOLgpq/Qn1A8tNMm6O4AaVbuIcVA+tAK2x0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48304)
94MUPrxHQi7fr3biF2zOAxGnppK/aRGsZnvQ8D5dpgO7qfut5eDjrearCg2vVjCx
ZViWdmdhycbb0MjBM83LN+tSuNtDCrjyDuEqqBvg+URZUEUQ5UIOI+dm0I/2GGj7
iO4Wfs2kwBrkCzRyPN8qeNLl/FcPR6fdBKQ94aU4EDURewuLahuPtV9dz/wQ6zdp
KYxsmgibnWA/NP04VfACFqkHbgwP6ZqmXoPImYynZQgSKe1LVi/kJfZnh053QU5w
hq/KT3rreHMVlottyzomM+YNUcdXG977lQOeGfJ9Yw4LaxTQSHGJDZLTsQec3m5m
8tgxrMBokJ2ehMrHjidmdbuBMWqPSArg7nHHL5DMah9ndWY0jDppcRMYJrusI5Ul
eHSaPmTD07Cd2Z0tMZehUGWFEI1vRf2wYw9Jwh0gzlgSKIWPO6cIIS5eu0dA80Yr
PW3bAFwThHEdjc3DiFrBG1hx4MP7yQ29gM5YWAu0P0HbQfpqce7Fng7jWyAvVidK
3998fXad998tZnSeXjg4w5z+N8Fkm8N4I2oFOJa0rT605TrxK0jM8RicgiOURzQX
9Iy1o/D+v3V7fo27GAHBumihfrNm7CzVP3VtNoW4YqAoqn2pijbRyQqeO8MZ9FM5
RYjreOQ5etm/QnAvaNfG+rPQl0Mr/p4mpKTaUrBfjcrwHUX30MFsQfaqXYJjdSEt
WvK5DgyTLoxbx/RnBTOBTviUOmtrkHLQWb3JkUjz5R5JBMBhZ+sC9NN3mufOXH0z
l9egDSVHAo5Rn69OtN/rewi2PQUREgcYXJ4AYUyDutjNf5xvRXlA2+uMOE6rnG8G
tZNKdKdUXV6zQ94xShPEm4N0Vjs41gAiXJRUsxnAgNYOqSoxFAdkYv8ry60VwAIM
Pp5LL4010VtCgEIDY0Fk3JnyMu+YGG/PBPrcL8P1nKHIzbLnYYl/w8UmcDzwZs1b
ihbQ8rETCIIKB9JLPR57gAkeaV6l8ERw5rMdecm0kwA12FUoTd6S+sgN+uREbbf/
cTX4fohlg0Km9fXCAyRV2z1MQQzOA/uHWK8TxItgKgEHnsudlC2m8AbnV1L6Nx+J
qk8HiC01U3+wFFtO5RIH7CRqFmaHB67PKx9zFan1OfsKITC+LtNujlxA4HqCjyVt
RTFvIEy6GtDJAvIwF5tmjg5sR0ATLQii7NsremPHTeaeLg/LesJndTR0NfX4Slnr
UD55SPsSKV0SpTx3Kdp5FWM4I/6bEmr6XzWtKB/Rli6dmgo4Z8jbL1twfrqKnBj2
uhjxXqjjIPLdLJfd4aKl+rCVfzejhvduiYbCFuscpoA557u0vtPc6CtsdNAZVGGU
usdsQVqd1uIKBmyHlvwc2gqfHPdGRYHr0O2u/XiMMOaksUtsY8siNUCBu2b0nVz+
TqyBE2/7jLVVV/VrhV9/pPNbrvPgNhGEpXvWEN2kEnM6PXqYahf3wKjOzjZE+fh9
mWXcnYwPIzrl4p4u4i95ivfEbUyCBTlYpKe15z7hnjzBs9QIytJmVShven+ykE22
99CGx6gmdRBffga3wEr23kcjNYZ5ZO6nHXZC7SX+f1GoWgl9gUXmm1/VlFrAiTc+
UDlBQFwPPmtrmBgHDYh9wisQ6ZBO81Ua91mySivKowQdpiGRW2oyjhjntxJJafay
vs0NuUqOCxam8GOWi9ugjEYQOM7Y4b6/DJEf9F/c5x1mt8ZRWykylKJ48je9axFE
7Jf7SrkrEN764A3BlHSMALqzQJ0JGY607lycJ18kHnuPjpj7X7ulukFTNpAeyUzZ
UmdWO7YXn5JsHV/Wi83aw3z7NZ9p/5thik5/JzuQgSVaOB9AJyb0LkL9CjJXu+Ms
eYmNoxqsmcJOXYFFUIbT0x7J6y7UP5Fh/mFhNosaRjmGgKgZOgVUe0agNdhZq+az
OjSMn7yaEA6fPA+achbPB06P8tp0otpp0eh0s1rrs02x6by9WRWI/Wo28qs432gA
GUcEBP9QiZ+u8fdOz6hKCWuZvZL4bdDO/ECjVtTRfRAAuNkkB2eR/H12E6Li/W/4
UhWUWtCssL8tF3MUg+TLrCKNaX7djjCjXXspZ5azlEkPyhQ6d8YgIDzXWzPehJsn
04/yum7NmTmAxi3JGj8Le5cKADavMEkiaKcDBoMTvqNrLmEhMvTGm/hJG6JmeaC7
XhFhEi/5tMBjZlT8fc7S2c7cGBHxfs8WAAEyJBHf8j2zZjRGptWvg9PsUyrhFMLz
zomHMmZrRIlb/1h7TOsxrm6sq8cboNwc9zPqB5sWy603cOeiIO6Ns+0V2AfcFCnl
GBPZoqEr95IgnoTqOsbHSj2p66YkQvNzesEKzXzX0NhHe4/gHjWtRLg0bPpktP07
ZqtK1/I7cSGgHialVfHVQlWsJwS840yGAEfsIjMIQhnafwZTZ+rdWix553w/ucVe
VGCG0jrOlP+mZ6Bv/IhvqOD/YmA/xe6ojM0QrlXXK7oKfVuz4xFJGxNyhfG84EHG
GlmW3lkPk3loIXpUbbMDpY+ekcsWsa0pNhRGYpjOLcJOg45P5L4K7/fsLBZ9vdsd
Wy9YGj6jDrStEPCSz62vE6cJxCEn9TcWFQKc7Jjyl6P6azG8NjzdU0jtHTpMm2P0
Uv4SRkv+g9NBrlDJbCy2TWkkp6RYe62boG7uDtDlEjWtcNgfIO6lE53ZHOIqFRit
TjE4SKeXjMwJoSMtMFCH1fT3Yl8Pgg6sN6BAVKZE4/t1N57Q/+r4IBrT7vozWwV5
XQ4kOeS7sVrcpgu7nFa2P1uI00AwkVl3won6FSFzg6QmYia4CLEf01vpOO6rhVb0
LII+95k47VnaIMpJGWvfoNWZNKrsZVpv+EMoTj5jkToW3j9mLMGyUdDJ8XzqEOBJ
qYbMhdeBTlLlWBqQUW91UHJNUcMs1dhHFID929DKuIB9/omKWFwcsuntMrH7UEjn
TjU9Hyg0ksIitMYcwx14IYtX4N6JQ6J5Umd2JaMGAXHXFCHxmYotWziBWf0qw5IP
jQ1tp9UphpDROXbTQol37v103ELyiq/0beXpy9w4hbZrVj/CZKbLoBtQNCTYYafH
//Cz/NuCpuwxPQIv0iCuK+E6ZLfc3Pang22WeKmPfxEVcJWW/lH4rhzwZyS8+TPs
7M7+D8Bo3Q1ynb7k9uxEYH/6q2Fz7JjVSQxI5/4ijTXGAkMCVRVOXfWBCYTZtlMQ
tPV0gTuFPoqGvtWAxkUYfCq4GNVnaK/hxupAxVh+y7YyVzCrSA/GY+BmXveIxD8E
jHHhlDDD3VhuAxbAxQ24SxcunxYrfIodtURo4dVteChu1xhHm8uG3IzR4iyKar8v
PqOUat98GjE5ac63ePwvNg/HDUuf8z/6A2c4yv+X7adfx5ZAV/HlN0x0QpHwPWeZ
ooKvqZjm4PjC+Z3yZwOr9HoNePDluR9amekKEGIa9QwiwCq5xqT1I3UVX7H2Q8gM
aVFuzX/rqsbRg5e7N9lmZVUOaOlQsJc3Ap5enJy1O18R9UEjsk7Pv9+juJfSzveY
3+U55GfnHR41kl3ggUKgjA0dPnVoocYCtpMCMsc8XMiARepJFNgQmL06lbGyCHFB
y4uN2yZekI+xm/lWJMbXX/OW5ZtO6kiutMOXfkwoK18uxhMdHoHh26vJzFCWnM+o
QhldjPjuzkbuYwojry7iVEJO0/jLyMLQacjV7l+aXbMZG7AOj6VqJ4RAGCr7tmk/
h/rzfoCFbk7Uhw9m5gCBaH5+d7B8mqiSfpQpGZdDm7LcPd88mgUhkvg6XlrtTG/D
81g9xKSXElao8wAhqSSae/piT2+1vhQnvHYRsCz6GU4V3H+PcMstrKJYgLZAnLFr
v1NA6zgDMplBq+6GMOiVrYiR0aMQzCFoHQDRLiTHJotDeho/lamZYfxuv6uv9w+Y
ovgvwHkNOweflDT9jW56P1fYCryc6tM5AlOdaCr3J++XFzLttMnq2JrtQ6FsX8co
V10HOZcT4KUELrz7NdXzaX+dmV7/G1VGktM0Cp9ESAGP53eIodsIgYQlxu5Mfxca
lnjlwA1DkP7S3wg++MmbaT0zFjw3J/8ZDVI+Hg1xiyuBbHq/cEfDOHw+zvpgE1Oq
aWUsLQlVv2R0wNW2SR/kxl1290v64CdE5uvzMJQHrhm12Jhw7SaUyi8HPbG00tba
I835aYjc4LLyZeT8KlDywXxhV8+a888KlZJqZj7m1z14BD9vX8ajQWxsWINa+HGh
hK/eGP4Yhu3A2xktXAPWfw2sw/7zyZNFJAH1l5MZLZsFLaZQUjkmGKvvEzwdYP/Z
5oM8bxSnWawR1TmKh/3cN+41+rxkyNV0paYMjxZ9OvRn0b7GXt9dIja8wtFk3reP
zymlOcVcKl4RosagYPytRmXagxnKTC8pap/Bm33W91w5gTjTNqqzXjIuxpJw0O3r
O/XdyX21wr2tluvkB9dvFuox5xT/EZqQWuVJADm7O+3JJGV/8WMZhKthnA+QiyVT
xq7qTM91ihOWeuT7KLd2jb4hWiSCqsVR5kEPIRYCBgzD/FwzPFOTlKHubTkOJkLx
iN3NZSi3lT+Bfs6J0xG2OP9ZMlgu10sQGIMy7P/+sfAhNfw1k8lo21DrEEMKSlqe
lF9Bo5nYdkco2EkHyB0BdxzVY8BnOvh+Axwz/Q6viuhzVFiqNzjRj67p0hwAmLkY
i6xKkFSAKrGJl8g38Sdpx3Vc5+gclon9pMyoCpBaxp2kgVYOcPcLFdib4Gz7zsqh
J4Q4tnrwS2zn4OgHN14urSXoCHxky2GleNgxcfJiAcOyp3E/LK2JkuCijidMZBmQ
7zs2lmY19DiCeVSn6Xg3T8B1YKE7DNM42eVf62bevgG/CMe4jx1SXAjEO+TizxLL
Cgyh20DtqcT1PJu8xNgrhuabXX966Y4JTlqr/C5TXa8p8IYKVOZ3fk0n3QFsHdfx
kUjf1CQ3CJWaobFbGguDJN9qbGix2NB8aYSb+WqAGZe4NDeuPez/3gGgxtZ/P24Z
GPeHOfEGwv4dyBlegWLYC64SVl59Dexb3VnyH+Qy9nb982EM6UaicTEysQsGziIa
rnkAOgfYqq/XAm6ww+T6wMMRLPS5Jv/tNyLMQKMNIjg/BL18ENn2q6FxCrn2TpB8
dT1ToIaKel89c7ggnx8xYJHjZZDtE8lu7t8BTm43OYkoNkakiVjr+QW+VHXRu4W8
6LEWFvD7wsxzfrFBgvqBK4QO8VGaAmMO3ACrXmThRKsvm5sFdUSqbH/5s/crHT+g
harxIFuD017hZnirUjSYOfr2Rgoknlr7HeDdRe4l2PB45wosq9pW1hZhqr54+O1V
RJNdHlVCOJGxxhL2+2jbwqGf7K/6wwQHtyirTCRqmidveN6t9M2WbYsYMgX7XzpM
G7U0Z93ZB3RzxC+ouoLO9j9TYCGq5m8MSeH9QGNn/YRzWJhMcHgrNJ9WXArWmBJL
yE2nhsiYxBNfsh3+r/vVUo2pblJ6urpovjf7X5qN3TGuZ8k7Ec44ssSmmgFJfDun
/5EZgOyGfft90299RVf4biqVCdRwkVdk8nY+AycHLqfLK0gEbXQJKw8rKsc2RL8c
zh2/FOJ4D/2g4qXi9tkv+zmBB8sz3NRpASG8x0CtKwkHN1sOYA0iAxlD9ky9Dppa
DlS6wTt28PMOy3DzHNSXXpJ4yQq7mybD+9bIuAxBGS3v1feZVdeKx8N+nun55nM/
XEOoFapwZYeZ4uoj1sUbuQ7n0Hq7jTYDuUxkIGQFUL+cP3ocl0YNSRHw82dIs8n9
LWmsDb0NkAhrFI5xnukKcZCYOZWaAvAPZC+2la6o/NKAe7p6DeWmggOt+7nS6ZDZ
mtdZGRzeaYi1j6LMUMSyUK4h0ND3w82sWrLE+hBCxeBgSJas9RKpt1ZfuwXxnsDD
Tb54yFsvK2yuOQF4ydKqNUeQBWirmGGmR3izbO8viYk9XNiBOwpJglH5WFDxFUOn
e+Awllyu9pd+bzVhNpXiTNpjLUoGD3hLZHwzRkYAwVY9QUBVxrwWUsQMlj49B9aI
bQDhD5VxJEisLoi+zAh4kV/bcAtC8Emjs3pcUIeCBD8Em5xsuOngEMu9ZirvTBtJ
Wh1MbgT+ld3khyo5YyGYL46cZHY+Gxd0ZN57Q8dw1pOrltV2wvhjURV7G5fbJ/Er
P2G+vZP6Gvpb3NyUdw5YK+qdEfcep3nMQQlCbHNwR3M3z+IH1djRXvJpZCc51FGn
YXRhW0DA31xDY1DKH6MLUisA0SHjHXCctXbZHV+E7PfXnMHS02Ff84fnFhhtTxwP
Dh64yfNPWbS7YW5zIXPJ62faHYvZSMQPXYBRf8osbUTwEEzLlxiOObEzuYbu5G5I
rH0puhyj9/n0XbdyfjqQ4D561j2d2vepF/gv7Khq6P+ITjjEyMBmitSV+AX83xk/
VTucldYQfX49cJGX8T2TyI2r56WejWzTyuboJw33glAdnAiWPlHp7gEnVsPpclNp
CmG+O0doE5mSgjTsM99ZkDldpqPhpd72e2YFgrnFHudr3a2uuuzv6JYfJJWTDv8c
sXDTffgukBu6TblAS0GbAkKzeI+TVwJbHv8p1K7sTK3S/6NNkh5l6Viugd6Fw5uG
dqK5NclHZbl8WxLoXU/jc051jZONeDxwfH8L3/MyBJsG3OIoE3wC9u/qfF8pm7v1
3A6jy17IMsQO9+3J35mlvw7qy2W+sT/BUSD/YTkmSS9/0eiFLz6WJ5bWhgW0VRb/
7yeB7LUBZQzIx/YicbJa1Zsq7kkASbtGicrrJGhc1pI5CDnRaIv/lbhmiDxwfrdz
d7Q1G+fNtRGma1zrttbX3PyByu3LSOLhny9YcWP67jOh3GMDv3Gd8IhMPeNx5Hub
pBM1QUArz9N+QnmC5GEirrvOv6TLKv6nL2eOW+qSG16/pok8p9QO3LhpUPkLwu3y
S+8g2YnWj6vQ4bvJMgvrXw2MbSo75t7GY2HBDJUR6jjW/wB+1AJnPL5dA7yVJ9iZ
lBSAJw2A8WthAgTgPAzsr+V1RMLfIidT5d9QqpF8h0WN4nbZ/2s4TtenNhfudM+b
o5qOk2V7wdbBb7ma6AqqB0IR9tbDohxOqH4TUfmuGJt12NpptQgzGbngHOgWjrS1
bgP8rB44wbcd+wz9ZnUaP8XWHuoVuxYnltjflhG7MI77rtZS3nbmxgFiMjVCESB/
uvYvYdU1hqFgB84IfpjThM/tj7QCkfYODMsx6FcMeMcoddVeO1no0VQhmYxqAgwy
lmCDPWPTaxzAxfzghiOo/a8we1bzDkrFd707QWTZcaZguqROBLM20Msgstmsjwed
wh3pp7Yi8mLUw92LGqSrlEvygEULW4vf7F4b1gP4uVVbaA1aCbBwv0DsnQDVhPrU
bqT9Rk+LWB64GcgHReO+nbQb5/4UpsKbAiqlA2RNM/vjDvfWFYv7JB7OGmPnEaXf
n3X1ayBJS8sEYNSIZvSrwbPDr3sBSFSd7ajcN7Np2X76our0e92pzzAjzTpXg5RQ
BBNEGhwj03s/8f+MoJpKQI0rscE7FU2fKVidoQoBavouK384xtjLg9ep8pGV23mk
BWJjNikfRUnzCSn2D8J5zYr8yRXsaIoNCMCriOK9rBl+Hr+GUSL+35aEbwScy26z
M90xhf4MOlwfAkZh5eqGCTWm+irO4PumsZoN9YtNaHoDI9Y2QYW/pyM5Zp35nUKO
/eh49CGbXbJ8zf0xvL1wf1t1Ue3/Waq2yLtnCW1I16xnhgf2gOgpBc0FO6E1LNfV
OdRRAcSzLUxfCGhjp2VdvNETY9ggoiy1zlPS3zuWWorJsi1hEBMK5Yz5gEQnnHbi
qWb3rgbdEugvh2nPCPuf14p7/UjF0tpu7MHx30s/5eixWY1CtaAf6n0Qe0iYcjCO
6/BjB2yydrhZJlvkHDEJo14jJXh3zBA5xOWYUdgQblF+fOsjq2kjzo87VxaIBIhU
CmlVWtt1aHi5pkP5H/DHgK6hDnMMOuAmWw0AXo6OitjXr91FgeVAzg5HZGF8yWUL
+ZCXB7XhyJH1ODJYAgEcQn4KRrC/7K/TVUAkUDFezTTyVvavtM81Qq3EdLQuCM1z
O03Zcsx9Xv5Fllb/OhoQ4UbWyUu5st3A8MDuG+tKMT/fTCcyS896nl11mdo9gsMb
o3in4y5j4CNXBiLlFThIupWMuy95YIFxgcbQ1RLaswrillqDTdJMUeCjDuK8/h9O
oXkEPxPdRDTf+g9rvGStIIgTs8uGdeFP4bMADmmmYLqfAPr1utVOpPaOaxauhFEO
t8OGRkzKo5sGMVB3ujZHDfOxQ0JmZtHG5krT2uWqira9V1hRfSyMKOUYhoyV30+7
Grs1PdFv6vKz37mkpAJViY6qNnlYGKVFDA+/1PBfiVz+oGi/WdYLtg0WgkTKIKbp
jpAMQsrb19QBkpiwmB7HpTc2OFNsI/cGBlW7iLbZGrq232+di6p8UeUO5Px+rE2h
AfB54+CjxzpzqTEydRI9UpaExQKG+XexMK+pIV24woZex6qls+1Ogx2/KJslnNli
Q+CDQXi/4mZXgAExX1RQmC2xMU6Kyumzwdb75Nle/t9pZYYbHk4O13WJUVq+RjV1
R/gHWprBnf9PmZVHz28WPaniP0lKMfLARNitaUI4UxYJXW/fTfKj9Yoh+JLtTZrT
wX9GRVWUf/io54uSzlMiC+LCS0SWFX9hFOfW1sk/aSD7gWsgHFIrBQ+pAzsgZg4G
QCpvUQAeI4z7vvmq9MFxOU5Tox90yRt3Xelsy3CVuPqNagc/BPTQDpdx+ctsROH3
mgRGzHd4VkV8qVQ9dqXQtZZojgxviMnfU+UK+8QI003GEF3V6RFeZDRNfyHqGjPr
l3UGRSv9xhw2T/SmRkjsukl8aNgobywuffKf7Xsa9hEuWFtlkRCZI5F3e/KZa1lE
ENKm3kcondxOPNjTekmLTKR8tZ4vxxC7ynnu7kHSo1JNpE1eZx7tWV5PpeT0bp+V
kG8HMrQs99tIDPF2qhBl27zWPAMIh45gzn2tK5j+woqGL2Ce9A41H7A74K22xSIr
DRdoPsG3V1qt3LlNzKNSiloWz8CsQiH0mJVHK69I42JFXXs3a7dEhO6WzTWChJyE
DkY+IaExP/yEu+YiWmnbLA6J538WZ7QIbbq5RoXQ9IPm0UrV4DsvUAyLJs1eHR8o
O2hmZsdEzQH2iiMmpRdGvx5xrcz1G7AD3lxyq0Y01D+e+9qCjQCm/TuCtG1BAQnQ
5fnlNHN921MSDYzCYgasjMcYsXtXNqagZHI5+JY2eJLyI7OUrcBD8Xbzxk0f20XV
1YyzSn+G6Lb56244IK+shSomjUe/deMOY4grmGEYvRe4YsYMSd0oHC+l8sJtIJzD
K9oIRirye6ZfHK7Q809EldXv0kyX7PmM8VcpmGPcqZnOwqwOj3SsxzX85P8AnVsr
OCCMPI1wLdXBin97k83xWj8nFeV54sPSqWUVtJ0G/AAwtOlkaEchR3JUNz6b4Ozz
9EWOSs9bGfNq3YjdaLv6OVgLqMzyHPJpIRSEY9ws6+lc5NGo04O2lHhUrs5disuo
hcLMTlLZG2NKtMiR26Q/NBhUnsLqRDdS/fIBVD8VIb/GIzwnhnIwZT9leUT1ND+m
uhJDwxQ6wUoG5Aa/+F+r8h/wzcbo75FQRg7ZgMRdfLrlSbXwuXc8FJbL3ctPtJNQ
wO2I7ghuF7QZPimt4+8zx5h8qTtMfl5L8NTZmJ3T2FXkwBLlWhtXyFtVXZT01Zzk
Gq5Dn1oqRS9/B4mEGrhLUfpWnLGl6KEL7lsmAqrYFwwCs50XeHkaEjfI19L62O6G
UxTounzyBjJhVk6Dry3oTtSzjHPKJdqp+aw7UGgOcCnlt8Aqvan8+m3JZq7p50Pj
/9y1AZk3vqs7Qpus+pJx44r3ZIqK9nelPM+DgYda/ppHlwISAmfd+XwyHwRz7KUc
66oR8PU68RJq0w92rEeW4ZYpC27wTJ8jR62Af6bkmnXUc7fESvBgjLWS/iBBWvzF
zvcmofHSxQ0WZmIYbLPP6S6BlmiE5D3n179zR9buTDWWA2MZv/jg8fpjymBqCV31
ucAfyHrPEOxdCsPRlopyWhxHykqa3g4OEO6zSwW3QOsoAsuJ62swIjc9OCkEn8fC
+UzxEouJ0f/UMgnMcWT7Z8FpCEiaxE+gYeMpaD0Pi8T9iknZCOt2jF7tUSec5UyU
970KQP5ftR2R7lCnNbSbrMkQe1XkkubfjiqzeUpBMZVPBNlXxPpt7g4+r5sQ5mwa
+M80c2JopLdeGxKBk9N4VCFohL6ubgu6LOBUQkGwDabEtyZ7YaPXx9kG+Ow42VqD
T+pLOpEXjL+zUPlyUpcodf/ZW3zZDsVV+w7tQCKBxnY72QQZKCFeBKn020K4J0ue
7x9MCkvD1/jxg5qZKkhZ+SM5hQAGv+vE5Vr0vcNvclVdY0PLsBuL7081+9/DPv46
plEg4unLA92BkXtmJSiQ0Umh/ubfmfkZj07tvCGRDtHrGbthKjM7/kKV/OrBp1Ez
cx5G8dhVJZItpDYoL7TQgpJqMl9aKnC85U8LGzbBETSaM40fcUY+BNT36/Riidih
hkOExnYteUL/xuGGTRmGlCQhMEKM5d4zuG8OtoELPBQUr/QGPqN9GAzEgeqSs/jh
bztDa2sGzCp9sfxfDjnd+Ti/EvlNpUWzw0mctee4ukupH1gGoTBIHEirvkc9zaCw
q5hshqZyPSpFRB2uST02DjuwjCu56NnSRXLh2XGUQOcFrRT3Ml1JaN0+ERaNyE9b
e706a5OnYbxJyYiuusMOoNYenjwoTek3S4r/D13hSfVRlC8IKMSu0PCdG/U/7O8T
qwJCwPpwRPYZCrF3sOF3x5NYbfWN7nNQ2SKlM8RY5XZclkxGPnKr0UY8ZobXdlmR
/2WAdnsz+pQ+McLrUl/KeKpv8tihKBw6UmkOqTVa0KYytTfBC6lOtcC48tyQMymp
3ut/aAYuzGWVHqjF0ltGC2gIWtdkusWIvypH7w6bds96XuLkp0ObCcuf/ljCulF5
6zX+AJIvItDD6lAh19WOGwERU+w3T0G2JYZFC8rtBrTeF3aqCARmwAlRlmQAZGg3
2rn1hwqbsg4BK0Hx2Y8Atigoq7KrSeul9SV2hK4wKOW55QcDK9rSrrsOy3XwZiX/
SJYkLbIdXXeyid9blRv2IvrReiqFpyVj0IjM50RJ5kqRpegDFXdMcGpls9MJRxOs
uLhOkZQrpJQ3QP3IqKtV/duZO50DH649qKQ3+MONXjSTCGeEy+xjM8Qp+2qDa/gp
p/qRwkS4kwTAeGSWksCyheDX50mSSe8arFc6AVoA2KSvkOsUDILocFuU5i54ofhx
mkvUvN59o1hJOJ0EMVecY0ctY6XfvipEIdZ9EP64BZBCd2mbWMa45pLFO4YPE4+x
N9AGeao4rl1AcBwDuaOgOl1HM2TuXRudUGLp7Uov/22fstI+ehv0XJYDyxqq3TjE
9ovU/aFcckpkqKXxLflps6NiVUkPEg4/I9fsNsCYkSZSLzeRZY2zPHP+yzEQuSdb
pPXpplGIOEkcH1+d7HjvP4oiA3hY3Xulnko4c/alvwSj/PkqQle6Pks27naMWM9Z
pPrRKpXCKCY4lAJD4/wnhJlGIMIehnzGr64SAZR18WjeNKNvOpVmFnkDEb07g2hr
S5B2u3Wr4Ed8/kfjZhbNIopky14V9mp81XsOzx1nbiDrbsERuXGfxGHlgsMQa+QA
/SQD2D7dIEiWpm44QTSsGZI00s9m3iCepxRDqwUuoNMuspgt0IsRJ60DtJXJALtz
ZaJ1xNq0BkLMWBifId/faBbW2LRoOeSxZbEPj8+8arrQRLqY6gXnAQYZmSSwajGP
cSrGawzwjFvOSi7eW90UVGsydLXJ0L/RYwSgI3fvLgHvJ6uu7h7VQeJAyyrhrQQ+
OELAZcZDHydsKrzCWr/ezfEK5fBAoOgsSfpoORmdNVm4+McAyksle8f5aeMLRvAX
0f2rBh2srWreAZWpcAAGn9mzUZEML5OS3kLnTHCtFJYe4bg8hcYM/by7FY9meRD/
CpySxO0uK9ljwFjO7zl7Xuwh9fQCrsJU1gm+xcvBHC65woevhlpixE3hD+7RMTgb
TAxoMMUjnQ6I6IUnPAG36a7KmZ86rkmbYL8O2VlTp/1POTabNfx0o7JjhRscnUaB
dR+6mxtevQLd7Sn1GQ57qkrtUH23glVBIsOEEK7+v78eSNotq76WD3GFO0KCMp+i
l07Pgis7ejCwUFKi97OH8/PnkLGEpSvs7VtiQ1MSTehhr3FbhqttXrjJsCjVyCWD
06bFmJ9F/KOPCerJQm/5VTEuw+hQYEHRHti/IBbGqAc+nbhfyYMwCqnL+cDp20eB
iD1mETA8oS4C4H+RH0T3E8dqGtaLBc3pH4AeeQe7v6Syo5vlnJ28GT/TgQrGjLam
I7OeN4GyiMsxeq8klmFeD8Sg8SjiFMt0CKFyDnoWUZ0MLWj4x65on1+YOSk/hagO
sZNIkO1HH9qgvZ4VrMXNMZ1ReG+qdr2Vmw0BOQDpSUb+8NPIlQCyaKZTGzOyaisn
5D9t/fWlykpL36mPKAHtcszfStzm4xbC6qXcJu4kmjrOyWiNRFPvx2EXWWRKc0u9
27/xy7fzPL3ZbIfyKHOgybLJXpzpyAzDhZ7F4t4tINaY+Np+vTRYQD76Bq5mazFe
zygbG58YcxXp/WtVkkF5H7OL5rlJfSs+TUFCeQDe71hfVHch2mjDRV3tjM2RxCEe
o0ccloycDoXtaTBR70s3OHjnk/XPyVPBdWzvCiFDLg+lVWqxoC28n35wJeitNUCC
I5blicxNzFQeNJ08Z5kdssnCiu3OBaVeZodHYmD9KhMQKhu5nq/RBe9fchgQHejN
6d8kLGYzpaJj161tCryh6hSFE06LGxnleIY0cuhu3uvKpnbybKPQDORdKsO+6byn
/kVAqJKa8kCz5BJ4REvvQ7czPMqorpJ2B73ole3Ndk9jDk4mlLbW7KAh4cfC5mSu
bhtrIJEskd1y/9RUa/4mh/3/3bI6kxb7Zsc7AYwfgNCugFF3R4AGaklVSIEZ9hlh
pdv8lXOeZNEVU9nvanIi713mYbXad34d1v+afbCNIPKUrhxZFkDdLtEDjIQEe/D5
j7S4fedXtVEzQuD+E4E/rYxwao+wGu790EImYOW/9BnntMPzzGTJQ/zXzRPQPAdt
pcWO56lEchYlfEd9hpAjkNig0dh6xypV4AAKWEjhHdY5t1khAZ6o8R0zcoE5vRe4
sYLt1VKFMPFym7N7pGEi47GYu1X4y14ub8SMeuo8jS44ZJGTh8/b0B2++wi1Kq8T
fmQbBPMgK8pJ5uedvaSD/Cz/9jCEPHxnCGElsBWxhN53QjeZLLCyf5bnFs8guBsW
IKS35KB26WYqUCw2OIRem+b5hWwE5igx9IHnJsXxzgJpcVlR184oNEAvIiVq/3SW
1TAg3IYsgEmN9mIDRDkx6fPGb7win4DOmL6UcDAzZhU+lU2fnMZU7ye7DCPqCZE4
BizMUfysZ+nxcvW33Qr4dk1qzBRHF1uwZeCJY8lOJtWSBDfyYMhXsw7U0zcz8smR
WZ1ASwfjzUJJqSAyogoyTlUTAUcJdXAa9Pitp3RcJnRLo5vZUzRuLhEto6Czc8o2
GeJJAwDUiEr5eVaxaKl2+RmV4SdegfqsR4MJWgCNrf8aUoX/J6z9SioVJ/85cJj+
OB3kGFmcRYk7hZngWXpW8+I6Cy5ktTrBGG1fwhIz35nsXqWzSSoY2FswTcZqKFMJ
QDw/JnOSbgaQ6e07+HH9RocBk3KGyoJ5jm3rzuGAKtNEHCCErH6qPQLGNIVdUOmS
NkcrQ1jnQKnSvCubPaJFBRDDkrjN1kpVgiLBSLuYfzTXWGGj5AFb/SFis6EcQox2
SeFn0C2GzuXMJGcT3XobMFXacbPVxWCFTyFlSY/HzR/C7Fhguxs38cICUqBDYgtz
1or2a9tXfVhvT0to/OXxCY6r5X3T+PC8QpeviF6ie8xxDOC/dKkGJkzUEQJZ3r0S
t27SxsrQawCt73mTtWezYdRAKh27Wf3HGR+5WYSUKV9qJQQyfT6gYzl+SQGFHMpC
krdlpNROiuTjsPpHk6XGupk3AcJ62H4E2lrsdWd1idWYUmUTP9TfTRHZIHWH5Hdq
6hXSaq24mcm9sT0C+QgbdeN1cjCWdYUn3z1Jh+n0iXkWi4NsgmTX/BVrjxCE53by
DpWVb1yQ2TGDUs0vPgBKi6TbTM3IhHUWHajtEl64z8NC6qp0AYoRtVrYfgMa/4SC
Zp4DWp6d64+Y34Ry1Xfgm12se1YnawpBB1YVmAOXPvyjYlvQimdITK99+xqZFsmz
34r65uaz0msdIk4Pncm0mViXQRSU6tqloJgexLPbAYp6x9dMX+FtxELCFuixkjV4
X5R9/3oAcv5WrQ23OrKfyAXWj22oMynv1WL+sl9dhCCqQU69vb20YETfRPqGx66U
HtEz/S/w6kCPgXFSKqsnld17Fs+7DdR7Go5q6fgqZf6FsPIAeiFBqnRQ7Qs+L4Vj
q/DfM9Tw68mMvoDrnCNr8jvtKrcxwRr4J3DXJUGWwH3iQa17IEU6mdrpcP5bOsvj
6sf3l7gn/EFEhPaMZy/UaWt3oYscK4qiqmu5L6bPjawyHq2mNCZDEcnS9NEKc2U+
T9zhaU+uOLOWBjSyt4xCoz1GydQi16Z9N9YjKSd/dD7L1Le2GDvAA3nHmcJsGY9b
gPu/FVTrkxqUUEj9ieP+s5SMJvAJkujv/A5QAErJWrksrMXhqUN5Rc7+1VLije0C
g+HpIutZGw1QmBO3yZqsD1YhZvd3BCP5DU0UmJSoy5KWgtYMEPhbTUKoVVoJUOBI
Hoe0jbhHkfpcuIbnWetTpKJMDPMNcamQm4s57iGdzlxjUeGtl+jL4GrcV4mdDTQ+
kgNp5ufz3JlDzV9kEZKB9P9gUPkoOLbZlMe68SIiNgxORNTj+c0t4lA9NrTPqCN1
0WOcGSe3bkAYM1Sik5TAMkZHvkw0jJ0mlZytJPh8zEafMtEQP23yduc2wFUtlvoy
agaRnX76QAI7uJg4XK0jbuBkGOh+8FEdAkaNKt7LTNuRhedrSHQ91hT3h1i1Il5V
imTmdttChSSP4vWq2fJ+XdJJuEfPIDCPkc5F6MA+AX1hOSW25KpeuCaAOdRPP93C
NwsCG75Z3CuAPlEqY+MZybjgtKYI0Vtx8T8iEfzuRzcUoiLywXvptPjxvogxZbf2
axLy34jJbOrwWg+6AoY9weIk1QTo5dB/fBgnDzq4LARf5Rz5tYKSvtNyDeunzSaI
CauiUBHB3GD953/dz/WWZmncphXjGBAJMzm4KygzFjkTfPVZxM+P30eg7swn3KMX
wm7+1BzcXrwPxp/+EC9qcYx9ZdwzUP/FTNfYNpZy0PoVU1l4rtWs37fcerNs6kt5
uXLePDkE+fXZu5m+oTgyFhWsKLAwP5DIgy4OVWvAPHkRk+D16EAyPHlgzYrzq0IG
vYtSPH49E09ywGXlFDOYNartbrJ0t9zq9W1l5YpR+4qo8/m3SOQJcz79K41xpMmQ
qOoY2nIFtkn9ssal43aLCOnrHqzvcUmqFK945PCyUHcWfe6XPUAfGnM0krLwTcx1
n0guVBvfdq4velKFdA94ZXhrp5Q36HbGRubgkQdutrV9SfWS694Z68mq1oNXAAkT
lUsTq1AD0LuLYIxNLee8PVEcY0EtMvOdQqgFk+m3uMTN2IxLYV0cyHA7aISolCeV
f6E45p88BfLpQOVGXorW8m7HwMp2gKhXkaiVsxLMuDmQadWMimU+QyArn6v79zx1
GQNMOoTsBGuWDo1ktS8RyR2qk4V1Mx3neXVoiwF568wuKCZ+w1sjT8ejH1qF6DfC
acWPzX/w73yvv4S15NB4f7c/HloZMnX5PudnbrPjwmZETn7puFJaHoh1CGXAyOCc
fO/mbSQm4qdOsIlzYRYBtqEAhcGvCasV20eQg46uByDIMYL4mBqLbQqIWi07Ut7i
b/79rSqgcZdy5DhEWjHRs7Eqw6+bfDC8AWMNbFUlkWoAKlQS96f5TNyJuM+ZUfmR
RZbg9KkRl2tv4cv2FhM/5ZkvAAVjpMU4iL41anl30mItI/xlpdsOEiyKzN/WqNiL
oLm9DF6fXSQSCSgyMlJyPffRZyT1ynH339Yq+xcUgM+j6H3vf3wiLUKqiLK8UeKP
aU8AkYWyGoDsIwwkTgxSxCitMl783xHt2EKYWhHXuylcKhX7nejnQnf04CtmvDku
V0K4uBTeKmP+gKkhCVrNT2ttM3Cf9gsPgmwFyva0mVBwo+GktR6VFFC7VgPas97i
xT6A8hmFRcGvcEPrrdkJKCT6rmgdiP+7ok/AHrGthL4ziGoXnCGtiVBlXtqaBlJq
imFB584vAgPuN7Yrgd19KCsHqxfqnKA7QGJtfX592gaTCDhO9L5TIIx3mJrTbk/Q
bZjhbAjQX+MbWTrrPoNd9/c0E9WLtXFoCCCA7zs+1gnZOx8+zcKGgEK1lf1FhGQe
Vh6fks5Z37muO56LidlE37WfLv3tNOwPTaRccVLjAxvxAoGMEUzpgbIVlFnW3XzA
ErSueSN15mDd8z7ZVQl8oNoMQXJirqS6DTuINO+s0CB4CLCO8kKYGEraTBclJOcN
paXkZxX4y4tfM3j1FKZVVdRL2ewhxDh5+i/8Un12J04Stx/GqdSPPtCjA3JBZeLl
Vpc+9d2lTVPj/NapZ8ObZ/Xud80e11wscYM/o1yQ/QxFu6hvCYNa62+aaiz1pAkq
YQ6jGjSBJLrHjyGtxUljYc/9cxynGhofHt7zPBHyt1xCYX/iuGuBzfc/joIdIint
1y/EAvZ/RTvTG+jo2ucnzXx3qEU/9hSx3dNVNMjBk85ZSi04ZAUOIkkdSU0l/sOh
nCZMsb6NbDSqeeG48QQRXY5fotb7bMvYSYOa5JSfZezp8iGNF2cQ34gLcy5HCfb/
IVYDqqhMtB5sanVwuyU7r+upcjb8ED6V+yt5wf5DadJuWeKFV5Yx8pA1KtQGLuH0
5sAE+4jYMSqFlVnL6C104WIidbdEVN9cme+NJwUxDcEcA8V9oOudDizZ3JY1jpEw
y4pES94zGXLYJ5EkCa8C1THmPXnP03LvP26vtLrBPIMsVTMeQHpi0wEtCYZm8Q2U
m6XHhVdEqLDffWD/giJ8W1LE7Y1gM13s96xpJBd8gCKW614UWW5jXD6Y3pZtksgj
RoBWRY3TPoiKlrg7xNwKMb5udKnG7Qvl9mPYkqwpl6vK3ThzX8w9bN3Nc2tyL1or
9uGQ3QhzmZlRV4CoSb9n7WzaG5mp7D8N6NdZEb4DETiZRQWd5BewmeMkE/4bhUvL
QPm3i30t+SGDncqbY+FLS/0T/QTz9LTuYq7PqaSJaXVMAYgJGI311uYp8rmMrIMS
IHS5bQ9H2Qr8Ywibb86veCyiMxUPI3aewgx4MEjz46muP701vAYq/6K0752pYI7F
CV3Kt3qhcAsPzBgcTkvjQZE1waZEOrHMKsnjFslmc6hynlCsigWqkZlcYAgHd1Pd
bPniJopIvyUCfCOC8A/KCnghPXt6YrmlLKSeABVGKQ73sI5RMb9kNVowmagh123j
bHauERpdxNTwMqvkCh9SkiOXcscPUOXw7YB3y9QzWt3xzmjjeNYOo9R/ZCQBjI11
kXNnxWbSqv1kmpsav0aThAkgtnAOvu5qCWfEkgVzFAl7b5yIMHOTi0pb5x8+vNX3
SEpc3ePVJXp7aJhLPeMGqlrgjvchxyZ9sKIRiUO72mPeO2DZIhJf+u6MxsMnUAda
H+QZc67AnUe5igjYvRUFPXrcgSM5femiNYLqGwttds4H2N+phXTmcg87MiJoVf5e
JBQ7A201w4pmwmV/ltjGx0hXWgKhBzftl7kaBvler0Up0UBofLOMUG+suRF8wKOn
2BiZiiNpvvlJ3b8fwrFSmIV4fzcTfmDvSYhN72gRx2rsQYEf1UeqP7eMUM98xsQ7
4rT9uDhPOvjbzr7G+vWEEfPNv7YBjVq3cyixD8ACG+fCM05IvJmvtzRnPHEKfRM/
uuqYJm6w165RAf9ZnMaCcnz1mjJDKV8TiTs9CWBzE/efNVPtU/0Hacr7dG1uvgVj
Hu8M8toWdcDEFKqUPOqs1XVB0Y01iLDbIA2+lTHP7XofYj/sP+2ugbhAR9bWzjFu
NH/5oddxZivUfbVW+XDG/pDb7F4JzUvp8Vtr72i/foxSn+ICz0xfCsxsaYVDBKZO
Tq5CwfHlq+vB/hWFJ1nbR+3NLPy3Cr/kU7Rpi7E/IqRLjDtzfwHPXIWOBqYk33PZ
DdxUVMh9bmvf964qba8vXpuniV7D/VSVFYY6h075KFaXlG6n8/qxZEhdXIsv5bcS
UxhnN/HsiSHDVuEL8WlsToqU4AChc89TGH15DkoZeB1ooC7s8bqm0ZegQ89FH9n1
exaqPCWyfFU5wTjHOjKtLDs1Z9kq2U4PxLzWBnmBbrjtPEuaG3lroTyNbA394mfV
XbEMAywTWdPGPDgp2K0UbgEMDP4G3bD7RH2BIRxrvOkMwZjLP3FvtegUNMNuPo/z
0BzWApj6IxdsjuaBlEZpDf2FgTIX+Z4ZRoOfOfMepVDxNkYOt654ZUVSjZZeybC/
SCyQ4Br2H3d6akrTk63mi+WVSUS5QBZ6E80TKfgt7lVzmb9PiBHS+0dt1ewvQBht
g+kktDR05kQYLaRuOtdJ8DBbxGZNuimaPegJT4mf5dgPsgpHhmgHuPd7zu239PuJ
4jxzFvpNHwRzuMfUA5p4EipsAHkBcGnwR620enTCpkU1+EDvueg97vTeRBXB0HTc
/HR+MuDZAzdgSaPYb5r/4JlItY7Awe+eHwFg8O+iqzrG3pbvZC7RTKmZ4f3gL/Kr
UqL+Oz5wya5y+ee4oKbv7QJFxJyDY36Z8JeiMR8qQKK6qrxlmrKlBjXiSMsiVHHi
by0wcCBdDzPQrebx4zIZ8TiFLkOAz/9U9dPwPvmDacHSEchZu2fmG6tFzIElcsuc
QGRLs3QGBzeL52mXaY2pisZrjMNmFA2168J50PYMvC8PCh6crK3ls29z+Ih1ouI9
kwP+TmCtr+0qoVyYywdwW8/6c/CQX/ZQOBUUqWqst+iL1N7bcEo23ZnDkMChn4vc
BYZlnA1C9dzDQiOQSDf3rwYXBI5IGvu23Cb8wq5LPoiHEiw5wTXTlDdIUFuVfQ67
qTdvlNh6nFo1Wzik93ujrNf6zKb/Sr2F+ZOKN9Ed+YV0TY/I/JMcqSep4hWLWr6d
PqaFYAqCjN0kKBW0zFLZO2Rd3PFDMlwnBiGBVNbHs4KlRZNhGGT0VgQ5jmK12d3L
VQIwfi/xOv3ZgfeJbb4VCwScP89l66xzSr7w6Yr20JqzKs6XNHp3hNKLENrZDfDV
Akb9mfbJ+egd55pz9674SMn8w4oQX3fJMLLwwtrUdA7Xztb4LKF1HzSqy/ifh0pC
s/U+Cq9uyyiAhBj27vFrgjLMM4nL/86SLfFQ23SfA/Nd2SykAh55zF3uueirOr65
htj+nqRauqKAaMJzy0CgmzQEqo9Bs5aZMTnfPRVjVGHshJaDL0DaeuiQMj/8futq
jPVhuzIbHBLpVwKNBNT9EHT/L4ovksHKuGvnnhUnL1DcUC7FNNS8sDYJu/Pvj0Xx
pvhMJ7PKy37HcYi3SUsXGeGGnZgWDzUboULMx8HSnGdHrhDeC2jDMrhOryfHkwaY
WoIOJsP5fOgsUqKKdUd5jcY+osCVS4CtjO4FCOf+8fQD8MN2vG2Yv+F1Nis74QNO
TG8F252T61P32rIJjAGpOk+tO6XSgndDjInOvxF+ig+C4tUqrXzmtIcmcHquYutR
mdzZUvJRF2La7rj8IN+ddTMhzHL77HlLyGk5d907BsRE/SD/XG96ooj+pbu6gIqS
QBM27z58vxCwo6JpFjB5arpIBAYMQRLozMgXBuJcdaSrk4D0NUas69wLBQ+zYKp3
uM+SEP003GIILNLnJXFXIYoNJyfHs3E+H2mIlfq3O31h2ewjykAr5i3LN5nrioU2
9g/VB7S//Gwn57+MEFSzUqbl23oHXHOq9c+AzWiEXkU5uBQ4XX1iNS1VqPukiw66
dTHTMs4yHWCHqA9TEm/2U1uP67ivgWz4C7wtq93VdZ3iln5/8MEyVfbqvlKW+KCH
+hZOU9lrfYpTNEpjMIcBCzkhVqoH3NnqQFqvBEXvzjnpMUh+5u665ioQaVPA7wPo
iXuxjvdrsgEgZCH0j+erpsweh3cWN9yo3138Xfa6zMOzo0PzFxkKXvxVp9frlPRy
bxA67ui2KlrKu+b/qdz2DSdZ9PaIkwBxzcj2R7xfR7ufFJzH6oFlkMMWrVPez7xC
KCwojlobTzmhM42R8a8t2CNgGxSWgKi0rgcaVCD6HjoJU+2YZ4UHf+WjZGprP5Lm
oGhEKF3pKnEcvaMY2bkI32VJ/uLQBzoDwggG4EZNCaqR5VpPj++zsndtj6AotmyV
+VFem9NLJajcRLjv9A1+bQ6q4/TFCIiA6+q8p75zIoGrlU9xB/gTwl3451Fzf1kV
/0dkGas6hUkK2IdbKwTau67eo4qU4OZT0PuVGIJnYytdupM7BbqxHtxVfpy5xo6o
k6lyXNCNvekd5XfN3kNqbM50X9D31U24VzxwUrVcO5i73rhDGHq3kJcK7rpdNJb0
KjjxtJdAoHJXHWdWRX86J37iCptewbAqG5PcFE2lyJML/yRpk6wdG1u6wEzPbPlu
4sRzMAeTmJu7Q8BhXkgRtuSD77jGaWFsOaBbWcGZ9JBvcgrWddICKluvos6hX1yV
wSIkg3nGj/Vtr5wlLFgjkXJ+puLjjYDmDeGoUIpg8PntTSVg+WJtHOVilS9uxTv8
ELwmsyTo259rdu7CA46levJg92QiHl6aiLIgKpFTl5Ff1irdgktSybX8i1XE66ZS
JaDRDUkp4SiDNfvHQ0mJcCccwafP6tagLKyUSu6VpU6QQlS4th7540n+U2y1H55V
9upenQHcamJ7EPHfaGy4HJQYYhv5OCnMZSgsBdrrXHU40+RQ0a5B9rH59KSbMf/+
pwKSVCrAA+Sg5Wk2/gXICgsRrjq9SPsAEELIpSfe0NSj0HcEYVlIayeACCGi7JOQ
e4Dibh3vimHk2IN6b8PvzpzHpLv8lvSa8z71D3FQLsAum0WKIpkOommlzMQ8h4dF
yw7sJlAHwl/2UKyMtogY4Rz1c6etBpIa1r+5p1xMihEavUoUpUzJBlAPy9litM2O
cgGd9GO69u3iqE9qCyoD0lW6cBuRfWQIsDHvRXwyD2Jed4mLYEscJFZxvB9UNqxS
Fs1mkpej1FZSdt3aEZtFbHKhVu09FZ6cdyVNyYDG7qmoTpJk8ANGYaFpAeIrGWk5
m09l6nbS0oJxsZIpmz3abtZXydNqbdp5msVHnaZhOxZVihPgNMxL+FRxXZIWxinG
pBCzigk4GZcfNhsjQHC9EZlfV2b9AWMO0b7XJE0a+a0dMyIgIIvekto59eL395dx
L5h6dCE9A3g5QyvxCBcU1mROc8poe6hJAfTme08zRXl/1keYtSHmOfSDuameNKC3
X4cQfaaoFqdybijOm7GvKz9eS/DsTNWjS1oaQDnVCTf2P+NlMs8e/9fda4uc76p6
bCv60RbABti4KThOnDdoofYK6sJL+49oAldPR5RRSRXmddkJPKVlE1bRuQIhR3uz
FPLA+T1Xqp81awUsoohxzX/eNQN0GI0bHZqFLSBws0kvFAR1m7Cn6ZtB8b7CXB7e
vH1mEYRRBrDD9teMU2KVGTNleHFdY0Y6HKBFKR6Sq85wepXUcN3mIMG2g4X4zU+d
dgYfjNPLB7KbL/3yXeo+O9yrEkxbtN/Mla8FtXP0bywPzntYKubjgqQn+64kLTPr
LcpYK7aZxtmPxrAeLBLnqR2VFvmLVDDErnS1E9rHyB4cTHikIyFbuk8WDePU8wNM
cj0vC1yCbzz6qrPrDoza/rvYGo/Ck6amnsMV2m9vfBJlyTLMaI2ANvLcpyTWHIHR
ARumfSVVgH860VVoWCFuZGoAWuy703AlbbzPUSrQNudWbA2odBwj+6zobYAaFc4r
AvIMkJY9zA17fUxBuLMbqU+aqHmRHOMSeWf73I2kcPiSNBbTVvwz8zpg4WKgZEfT
X7LhWC+rb+E48t82vAvuSKj2Cp2LaV5D67Hj+KbQpfLq7Q4XjgY3N1hi9sRGHxbT
IepqnsHwBD5JG2JdeaEKG8TVw/Z0wrows0vt1Z4KA3BiOUPOHiufo/Z1tnMZVa44
h2jTYT5RPDH2f83lJtKq3geVvPSkfnUH0e3/NJocu+/XznLVNPVoRACtqjhTbI2/
hy1QaZpnITKcXOdxRMuX8RG9tVEM9ZGGqWnPKZAMUn5cuXx3avzA8zBi4Egv2bxs
h9jEIyjb8bHP3gewuV7GStLSnZsojDQZ8k3Wmr7O/PpkcmArHTML8pntYkfFyVas
p8NyfqvYuCdOwHF2OaCwNqyapUNCtDPCp051HkPyP3GJHk7IEdg3YDQ8gDfQpgMm
yB8NgvgaiCpwc6KKQfksUf6xiDj/nxzBknQbJbl+LKtf5uD1z91Y18DmjdAo01/j
dV64cTvtYrN0TlwoFDpMYp7Q7cpdnsv75UmpZd7ldjHuwabuvhevr5oyYdz72qoJ
kHsXYZ+tYbq2VrqXtUSBY5REvj+f05pN7GRs/YE71v4AJecRvUzEIcW5+6Fnv1ZP
CJQ7AzSu5IvKfcvuY9DHWhgKmwFOIIM/iAmAtD7eb6zwp/eDv/847hnS8s8H5MKF
OOWH7GAecvnwD+lNNZ0OqPBHkk/9AGWEupQVsong5TPL2ziNC13RFOtKxyfjBz/b
b2Pjn5F/eFs3NPFqNn5IeH7AEWAnN8GcYzpOv6kkdI3T7IfFSs74XrwwiUjj/Zwo
l8kt+XFSJS8KcEoDZ7qePtCSCx6/bOjF4/nEdpwX4wswqAtkQy9dyDT5m+2okhKs
0UftVOVI049GbKQqjUpEvUApBcGJ6YOGzAgWWAqyvwnEHkeQVw7k4WDgKMA7ysHy
QqZaaBhvgWjtsCtIJD3vSabvQpuneo5wMilrsokvBop/ku522o27LdkZ2u+7wiWh
qYGzCBssMRX4QvkqfTiJoVqyFpM3GI9zJH9qj8evnm4p04kOj2Lv5277vt90wHEP
CWP7Hc+52acZjt/7vjqew9a2CtU7DO9smNUHpgeFRAPN0gCLYJQLfy+pDTDf4Ywd
xXBrw1YMmQTgTQiyrDLs6JhlzIphZbnM0te4uW/rwjKPVRIhicsd2fHjcZ3bMcq2
eexIcFlmnQ29qqlRBPh4iBFaUxBjWYhQ6b3Fwp00GjLuwK+Huvrr1AOg9LHN5jAq
r0lui3qev5+I8PC8Tm/nb1XyI8cVCQilI0XLCsKsdtXqtOfTACPFhBqCOemAts3U
8/C0X44oaJv+utPXb+KlXyo+y9iBpMo0Qhf0L+5EQgV7IZ/iJ0SJenMrnwvJk2da
xj+3pIth8lOM1TuljXeRVTlQYPMmVYHOlMEhJ3LI43ullgaubmcH6jaoYn/aCwCg
HIkaDUiwCeIOQOFjhkw4w5fChsgx/+Qh10BHxjvP9BkCOwVUunpn5Fr/qjxqBxnn
R3SWCDPb+FRjXbQBj9p/ST+t7PY4gj/gPE/jCjiX3h5MWNZAFQf09du3wyLdFMxC
2PjMuKxat8t6Ijp0B3p6YQjOAxynI04TtmOHI70nBUSYrhUaA8cI71EWkdbFBK3H
fOBqlIQho5vPD3d9cTuzp1LZgTvLcm5n4SCIH3cteUjreDaa7mfvU1QN3xZcaG5l
4o9H7Ipp0vif90rQ64+qeZRrq0SZ9Qv/6BuKhAA35oAslkAGZdm5+voJJtMtHSjr
H494W/mpfN4fB6UFB5xpgt//IdKlhLf/Ymk8LQwaVXu4kee6LcKD7DWc7aAgCXKg
BAci5NwF6b93KYx1DJkL3imeuQq27zRHatDIdjGjyW6aZsiJSr/z9LOoIoO1mzMb
PdU+3nKwDS/MUEB++v99yLuG2IQS+Ssqaxr/AFOuc5VAKD2krOoqcr+KEocjzpm/
ddqTcFeUMo3gLY8iFVD1L0hxzTYtkY9uqEDv7oSWnu8y5gYADEcrU7b1mGf3WfCl
qsh4Q49yXEDC4hjC733FIHZDs0rKv1/b9AegGqRuavdswMgVhB6AjbRa6XF2y2cC
0iVI/pAz/j8VNvPbucFr5+fokfIHk++7lv+y2wXrevhomcCTu9mcpERkPCyCgX7k
NProiO0Sv5azFKKYZhIcrKvxTPGZ0V5Tk8KrL7v/WHMgX5Gm5rLg6D9qfAZxG+31
R4zOda8felSGYgeF8vdNd0/vm+geAsRZ0BfpLRrM4mcenJ3XZorlN2pelIM72iCg
JLTUP8OXIoGqs6vu6FBeMKSjNj4O5L1nhqDute1+MWKcNHtNIid4a1NGiJ+qywsB
uXPBf1MDI/JBuvijnGrhtwHutceBJnHhCsPa98E+/ER0WMjyQj7VhnF7kyL/7Tkx
KaxPMYuOt91FykbJSpsh57SMeowHfhpr4doqNksIldFQU8YntlgvhyXeXFuPVIh5
Lv7aj9IL51vsA57py5YyoBjXZ9xAs35ip7WtY504k+iLXguBAK5Y0XLPv13yXv+2
BeePAsS0vLVE83jvtIT0IY4ZzeaUygK8hq6CQPudBPcfw1lG/BV6hzgMSelHh5kG
euVvXowkJoq58Foc/U5N4pY6bzlQRdofDNXo3jKd7ZKWCOC22xnMgGts1Gchm5IY
Uv8O53I8RSr81xdMDtQehlrtdEDCXBq1FGSn9f/IsrX4JrcEBwov9nwfIth5ONUS
5WzZUohVJL7aYK3RZWFUIfeta3e+hvr7x+VaSoWopatwxsOjo+BcZqKLrT72CSMS
z5Va0VfdvziMoN79D4cQ7M4S04Q8hK1QC5aBAVjj6Ui5c6Fos2zQw+LxVBgwW/EM
jZdYAB7Xu3gDDx36HMxs9qiJTvjlzHcVDCs/N1CIHEDT76VBww6SgZpWz7JaG9P+
QNqwXGsABPabARqFONF1fSE733aEcp+/odpFQ5VzOY/K0ppkpcidWBv4xlhpUA6K
LOVXdY1KqrMauGMnXfLsef3XsYPZOWyykALtl9LcBWCeEruhkAC2o6XxxlnQfaJ7
VszyR0t4Qvu51IznnH312Hca8UTBDkkvn+snxHAIS9AyyI27nQADbonx4e0GXmpQ
h0JVD1AVkL8L7WUN39AYe+ioIkasSjSGXWIQg28mxw/wIzE6ValenzSQAKngNmag
pxiSMvJPPhlDd3EBhfgGuM3dGDbrcR7Dy0qd8mHVfUcxnmC7Elwh2KJGwYX57/Qu
3clQg1BRIsnKqPOlb1yniONq7TKYwlxd52UZDCK+v4aEeKTkDuckxiQvOsWGeqaw
NmiSv8W1wsx+9iSck4B5JzOk7Rk9gmJP7umH8KlSLHnhGWAaCANYe602FJEM+gLl
kCQ5jiXs7bw5JDj4b3DLxwc4aUs8imKAO2zKaMzueA14+URt292swqIym5JP03l0
GgL/PDzTpEUHDP8CVT1QBH70IWdMIhJQ6o85+eMF8T4/h4YvzTriWtiyQwcGQLuq
ko4d7bWtE3nY6bRTOtx/Ocvliyf6gVXrG02XMByKCQJ7N02R6c+kxDP64tqR5QV1
0eqANBirIoA5a0FIsw0A+nWVHum65X9u0ixVmsT2xs/gB7ptuZdkeZDwnytbMvAH
dp8wn5GxFsIXm/MyLQVYtK3K3m48YmCSkzYYwR3EPvTeEG5AoJ9uqPpiNvDieRZ1
BTBvXKP0itfTam0LCNPn3lfEPL/scut6S1SvDXQcrAp/1kdnKN//aQbhUPv8zkcH
0tdoC6wFyxIOu74xZTY/BUR9XZif8nwk0MILHJW+vGtXboChBsK1tbu0thUsAKnY
+Gw9TgHum4OJuI4NpU1hZEksvPd2VS5II5Dt2BheIQRDjXJQwqS48t9ubgm82UQK
4YrhgulSHcoDVrArmzwg/S79tYv08+bD6jiT1yZ8PFr0mB5A5Sp2dSGK4oJH7VQ2
uQ4K7OZuRlzL/55YD7ZZTdG0EoUAaezKmSLILcppU4/f+/TqseP15liiz4WzfTyq
F0eHLrVkeqnypBzVVPmWodKC8fwDyNoRQrekuUyHUTrKM+Vs0PHPqX+/AzjVJrlo
uBVFb+O9pOIJiOGveMRbsaBxu8irX81VOhv4Qz/jMmJFpoaaG1YoGoJRGBQV2Rez
Je7T4GfLE792ocRgPBc9mbh4s+pKuW6cx4wcHsJiwNMS5Flt+vuDGCoXIXgzgyrx
dsyZjUgQvvgKhIRhQRmKTL7j0E8OEz4SA6Hy/PoxIIMSeJYTpc4Lr2Aagw+iMT+y
gC8483rI4xsRL5pETgBHZ3aMWj+UrMAbVK1zhbBAv+vhmmWl6UFAsz3N4VFI3JG5
Kw87qd4LM75P8J5G5l5iC2r0UgFZfOaZlFK8meCpaUFjMgWS5D0hLtNUE/94S6jP
HbtYX8bcRdkmCvnXISVzfAfusy75niehyg6kLywxnl8PzQD+srGETUbReV2YbHq+
x1+oS87ARwgO/e+w2GrwyZYLArp9TiL5Vz+vim4P+xy4R04h621yZl7dTDIUznij
9pq/hp2E3HMvaR09ficIDnkljUWUj4R62NMxQX0cNxasMPaxShTsDlj7ihvg6w2d
Z4q7jXxzQI7ynxYXN+PDwUqoAvh2+G28mn85thjyJdyAXiwgS2D5KR7ZQlnTadZu
cnUTjqTE8R2sNrpUBJ04W+8tNNT6N7fqoHYEmAiliCkvWfJwLxfDP7i4ZKV8haFa
JxuqctkvmiJhznVmfSMBAmBnt0mh4Fda/dd3Hb8qvtPVyhltrZ1ifIxGZg4+Hw8N
QKCzNS40NvjChe/LDHa8XPiud1tmxitGDohW/XVSAFCOnv8sj/cmgAUxcOkdiJIq
9MxVvu1J/nTnRWKNV1PJh5C0YZG4mdUa4HkFgrn8c2dyquajGzjttCbCqcaubGeo
bvuoXAf3tavhdf7o2VLQmtMPHIGO+d+PSjnCnkbH8jg6jhL5YqiZEMLDglSRscSK
A/MJQGUYZ6llEr7Qz4cKiBrPN4HjIUuciD5m9scbNfkJHesgA66FmWNQ+5N25ajp
3wbmnOmg8HyefemOelWGFMRAiBOWt4GqjinoQnMy0LlOPUuEaZOp8Otyrpr4Jpvh
vpMAOpqxC0u0T/uVBdBB2ir2CtWkYceW1rt05Mtu8tWQEqd8EL41zyLnK/g3c0zL
RWMnRU3Twa4TyDXmgsqc22wqeCK1O9EGBzAFMbrRgVfsTTmfU74Yr4iTmRzW1B1S
cyFh1y/ZuEVjYrgQz4MxIdHxdGEgLp1pXzHmxyk9OnfB/CHL3Ew2c/jzWFJ2rfWm
AebAHEzpzHLkOE/QkfjTh9aU183SSka+U0lDbeHtwN33XvNbehMd4SFfQKQzXGJk
nKBZza2QTPtEbNzR7P2VtF738dykd3Y3kDDYV/cK7Tx3M0BWnYR8cPmmOPTC0qs1
R7QfKBXZvKWETUdADH1gzkeEfSN7CWptvbT806GqUjV+hFF/gnyvKDSiG4lckDb1
XDqmRS00ob5aBTYAoQV+OL5iJCeqdjd/AqVne1BqXGriTBmauX5Y5m+iAdBLdyFW
yyGVQVKAj33ZwO17SHZhMb14wbhvgUwtXKX5WmGEPeR451MC2ZefI0MewrN95ueS
07LEf2KFRUCp/Ih5dFpt8dzyYPiZfvwWlW+OoSFwIk3HyZ42QlEqeUW1wknayC4U
4xm05DeBoSHXUhOf7AoknXnbemQw6lHRuWYzq0rcKd+TQHbpQhKFOAaqFmtBAyMI
XJ4cVmQHzHpq9wCN/4iSz0OLbN5XQ4aiuP8hMxmNRDXvbXfPsEKHITRTj7WgO814
xbD2AkBj2IXZBy8yMOauiNQsyuJlT2827rUEeFTJC8jljx+WN29IomFlucd8ZnjV
aDYWCkqWd3Vr+kLHbetDfqsrkB0skVwwke4VGsc9ZNNJ1zwD0TB3/y7RkGhl84Uj
JJVKNxv/1hEU3s66NMQHHQkb5hF8YTHy9WzMLrJSWMlzNuPv0xX2UUkuFXeFdXU8
wY84hW+XsCeJLMBlXlBtLz9xF6Y3Mmw8a++Oyx2msi0N2X5dwzOiA/C/KM6e6QNo
Etc58KobeqgVBvsHf/tJlS1vpHIoqScPCK9vgQOAEUpo6v7632u5rIJxI5XCMdna
vKN3D1SO7NHxZ6s0biAI1yNqzneAuL/hSl4UF0Io68yat6h5qpmwNoc77p2SPtcz
oixObNcLOg4o824ZoUjqGZCIW5ae8MmQGwl0NBcySm/elr/oibbibsY+3wkY5Lr4
FyRoC6utQsDeWMPPVodh/GWEoFPYekndTviSADpUWWnRgnjpTShhvbfwwUtCTRwz
TQjT8y6Dbm52XcjLoNZQJwKhiwHY8Ewt6sBNC/apNn6cWkkM2D8+5dQBOBKoE8Hq
+5RdsnY2Q3U0S20ag+Uj+DIAQQz+zFDwNS0TckIwQj7aeMhF1daxCH1HowU3V/jl
JkDup6J1mR7CNefrfhgfAQxp3IZz1hqiJYeEVJmu/nixEiqKUb4/vj1eO5tIUIfN
cwVftvWHE9rDL9lu5O8E/S/aOHaOnEaBxuJyHvid/4RgxvHZ5C2jeBbzLGYQ9XRk
Cdf74Hmea9kvuzJlC9pHI67/xrA4sAotaqGYIClMYtHRSbmYuVi6H3ekpLiRBfBL
hyghAZtyLbrGLXS3pWyrXRV0gQn5ujXwaLPfLEFBIO+wlvSDbk7d/FV1YwWHig3X
bUFV1U9NElGzvUN2LsImnlCgv7mHJb/jgQzwd14F1+/my7uGRRqER2jsk4p492Mf
KSqSBoZvA470mw89G+l6Q17rEMckW9UpA0wyqJq7dRIvEPqgyNRDtsiCo7fYy5uH
h2y4R9VxLtGSx3pYrIUtzLf0FN415nfICy4t9DWVXJLZ1j7y0beBenn58o/5EXer
Wd0Mn4GzXFJVV6/f02cZ+Qq8rdVF12mGnjJtEIwqzkrXe8Y/im5rjKbSpCEVzqFp
7B2zOUzDWv1O05xd25atFobo0rc27IBHZ0JVfLkiRwdtCt+F+Yd5avM3WygX9r7k
G9yXZFyoZU+5ntfQTMDvkBjyu+qDLq53YxqNxQWNaIRSjW0bDdkJPsiBItNIbL97
lj7Rt2hNZRGD7l1dJCgw6OBOi62waCGQe4aevsrocRsz3+onYR18K7tEs7qBinqu
rIPcEg9Je5L7mJofLuZTC84z4RvTyJTzUzb1E7KiANhaXno+ifpI4CdOBgawZRCW
60omL0h6E4FcN2HEHZJSkTnf3i64XgGyUkI9g3LwR/GNBJPDhXAn1f+2xzJOJDpK
AjvIHDRta9IHuENPV2L2SHPpvpwfTOvBre5HLj/X1EZKcodlw6XtA+NqZym0ucSh
QktUUFPfgvP0b0bmujXRMdVj8nNsKXWB76zHPgxUwTQel3pDX/dHSJx8+ad/rtff
sLa4jBHi5IjYRRQWlbecqfe1yZn8M93z5EyHni/lRl1jE5gPLLjmVEx0pR6rKe3F
TOWRh10/Jdi+2GFQr0d3+vaht0B/yXoidKfIkpCqe/kT1433uuQKVTrpArY6n08f
7PhzlHfmsA6dlw1rY4EU3kbAxzSYX8lnsIyTReWfJrYRaLGSYI4HI86VuFnNXZ55
poIWo8kX7k9S4IwjsHAe9cBeehWX3a0Jyo13Z47/KQV73QUHaN5W2zCdj0B1CKts
Bj3VZrAqQareVJTDqLAdXB4Xt5lAyQlkdFZHstbOhda1xZ98GYOTtmOnsBFi0P0I
Svq5mFkVkVDr/MZC50QLgqAWK/wLrnvdSC76I82LAHoig5x/O67r3t6lvlq3RPTz
RfCKXPHnTGff7f/aiV+CQlMAk3F2lYF3e12YbuSJIWs0HNCItRL3Gru03+LMTyqr
pBJoFzUIlPauSHwMO7qDf2aC8MMsyb0kl4zyNrzRLag918ybqU9MJWpMd1JQGoYL
78SDS29JgyvvbdZaxrHWW0xHxmtA3YcLW+RvwhsmlHGjGrqirIGmN+FMY+30+i67
SKzgW/2BkYqYzqH91r9VmuwpEtt7ctPArU/H/o63dcEsEWE9qHVxfIfg8gapGMbM
L24PMkoZ+dCkt3Zjfb7t4REJ5LVwSTbsOkfBV0asxX4sgQkwZfWAKFFNbUaSCWBF
GyexbDKINMrx1BJMMPszOPabde4EyiZUHtfP42fXd2aThMJmedwQpbyPum41odes
sumRA5SQQ9w5HEU1jDLkTxq3e3K7jVznLJw95eF/etoB8eOgwJzC7bY0IgX9DoUI
bbNqUenTn/n0TdBjgZONEt++Ex6o1kzRPteFR+UoOIjyoCFPnMVu5gY4nByvcq4b
TtZhtwDVO6Kr1hYC9+1GMxXbNTNpfP5jna+amYokrJgWURM69iGg3aYhI8XmfBYw
b8kV0Ocvv6rrhOL/2m8+mEtJC11ZY+fo91QY0lGeq2ebYnOFSL/yF7T5+j3xQquR
dyDnpHpZHMND8fn74TSHKL0w1JqyORXb0lklI4SrI0RfPGAokLcqbE9v6zig//T6
z2XkchXtSrwkH/QFY9clXQJK8H8poAWDsE/PyoDyfBxyFjbFsrcYPMH1tfAyIUOa
vW+h8W4hHm2pp9L0vW42Bo8TD/E850C9Q1jfYbjFAZWH1GeZTN4skjqnT0TCxF8e
KDc3eeec50EU0vwxjfA0vGIgu8VWk2A44iuxyG9eNk/MZS614fRpkW/O/FzhJZxV
BxVt+cXaHmdiNoC/tu2KmwvlVW4vnu8yl8ezmJ1msOGXM4tsT9N7LmvWViqeIytw
f2SSw2XD/USeJJPnRbr9WLhekEb5LLb7fbFBINSb4EY1hRN5b/aP1V/XCnhxypF6
OdR8KvoLC7E02PJBi7C1waJxK29IFwCrCTMBIfhp7vLrN7jreNwFNkGZAdgutAqb
t5d014JBnUCBYyehYNr17LpPW31Y6zGfbbpgBMwjk7utl7yHSqxRstNEvi/EceCl
WaRrMdWQsnT0B/w+WpmiRfLUJaOL7q3b720Ma4YYmBRqiJngfsiblA5/0mHyc+yq
zioEVGe1M2fBSHy2MazpmdfO/MtIhzQoWqSmK/mqAwD38FLy2Fy5PmQJC8b43Xwo
//EbLG1E06188jO9zN8IjhUrRUNLOdJxftRFwi3GXFTmUuxDiblkLuIvgfxoWjmJ
gAOf+cn9jD8EkHmoKYdYt3oRHm+OdOUttMMQzX6183UbOovhvbZTh8hy/+hKzXwl
WNctn4UBonxzy/KsypmxvblipvD5wlqgo4HhQIj+7msd6CSqOlCpgJ0SUnienilI
WERaOJkDJJAN+w2742OnaACMiduj+pDw1UexD9G5fSwK+SIq3trtquP33mJYb7gV
kYWw9GGh/hoAbxV1qzOSrLVXwgauK8K3wz/TYOkTo6xrlf4iK1gwpWWfEU1Y3A6D
7T7+PK6LyGnOwfudewkoAHscUKcbWguSWSjQHsX6y6GwekPAF3y3G0kE0ufwSNTJ
jyfok/SPg4p+tS+6UWKQBwyL/VH7k2fSQBrx7sVHArrGDss+oKFunJPbia2UNx4b
mImmKyfv6KwnP6ymgyTP4bNBxdM7C7Q1Vbh1sUV/wcFhX6fSJIgtldZnl4S0B+ts
AKJc+HusstOllYCpkEII1dPqz0GdmeOY8BL8VflIJh6nkyN81A8mb9/pe89Rmzz+
Mt2AEDrdapQO+Obbg9GUZzfGyK2lWgh/hO1vCa1KCvYX+YtgJ1lrWVkJj1oEVj1w
hnJyUjEFNh5d0D5y+05NVyK/FAfj8QPUcqu7UhoupMbvFAh+w4FoTCVaS1r64jlw
FOp2M4Qxh3kcY1bk/UoQVxH6MlFFuNSKXFKXhkAhN9OaWZkpN5mhFCoIn2dt5Oam
9NxOJvuQ55aEp4aJ3Azi5MqZ6gBKhj7cfigq8SGR7SZIu5uK2S6Aq3KLgkZ00FRT
DyvW1UD29dplVM8agQ1zLXEGz9HMna+NM6QQvAnEdKt669BMWOP2Zit3DHdLP2Jr
x1E2YYun01Eqb45UgN7Cz6JAUcIh3wVJP/f7/cN9qiS/3XN5FBuklbq9D8aIgxZi
XovCsv2EQy/+14wOfK/ELO5ufFkNQU3r9SLjXjmndx8jP4BCGl0ky2tEdXMynmKl
TulVc8TF9ow4gHx7Jq+7TQ2zW+kkRXUvQybyRugBMBBHlRIw32dnwfeMcxm3We5r
nqxS7N9sHZxlZ2IiwjH01NlPnkMkNuWhln+tzrPDmR1LDEFkMi9Wto9a0z6JDI6k
HJf4A2KhGarxSEy9hMqQZ0d/jwq9dgi17VHeZzPuadUL8C4/oUMONbBqj+7DH8RC
c+n4KLdgVINVQNFxFL0+wXJUPD1d1PZGmF4IHletfuk6EaMShWrhQoKhpstc81Nn
mDhzB2tEFLohGbDnqNCwPK7/aB5f615NNyNSeTZCVcwugzjMx6YfgMgFGl1IhlVE
TaRSh4HNq85KRgyJY5kykg8b1bow9nCN6n6WbITK1Cbyg+f/V/o9M/MH0xc40gLL
P/kNNKHmEhKWUZqFBA6zd/I4PdCmyE/xDPjvV9antYf3y/s7RQ5fy2+TfW+o2RcC
bgTNKZWnjXp0QHtQy1NBqiDgFpYaJ1t74hodnYkd6kxgd4kxG1oScRRAGc9m6eqd
tYoDtFQkWAQxTYB/UOqDSPz6OtBkgNmmWXUfSJ1/xzN/ccTpHl40rgMbz10tPfa2
E7Rlnx9N/UJZix6PMOyCUFzWpyy2dtnaIIXbIFoEgasabk69NnZ3jpa7mXbcvome
VAGPU++tlxG6Qxz9BBy7AIH7wRQOVlY5CJ5Kf0Yj5qHQY8yhMKc5uiadpUezTgaI
zO+rG+NWZVa05N42kXYc7aoLKOn8yevHhDJCb5ws6LD9HmbB5zW0el0OUJgrlFTB
mriIzaNtXbfERTaFf4NIQc/VltWwBNV9XAARgzhZYJazmKq2v6Q3DUjrzcov1hzm
uxI8NNtlWD2TEW8CGlDVdVg+wxbPsXx5tKwmRCrhDvsr9sReSWyMTVXq9KVXCBgp
0UA4iIoIAIgKzD0MQB4wfISfPNb7TacsAIwMRlrDjk7OSuudhN9Ur+3Npi7Vxptr
ixlFk9jjNZ45TuV0DrivU5GpUdUpPRX0lQ0igLaZyFhETa+NDNEUbwxtcvKstSPg
H3m+cIMmqbwQnoq0M8asHNknwobZwYgnbLrOU3OjClPZnkCRjXZueEY4X5iQX8YR
cxYrFT4O6IuC9OqrNnP3t7ESF5ffV79Km9StLCyIufFHZNA8bGSvqbhhMFwX/APe
sPvvmROTqQ9jk45TkE93Ezgb30sUqBAazQTrDuD8YaDFd6aNMt8mVIA3pxDLrNS0
QJVqqTlUZQr05A1VpMnqRdXmX+esaEJUbNMIs4YYIaeJjhztR2mJi5F67HYTPUvf
ECmGMpq0JKJFZtFsqnuEayJrPaNOxQXBhSM4nVz/h/ORthTKuuwxRFBMh/FFhVp0
/HnCvQ3MSkPBlmvtSxYgUC0tB2gq0Mca3NGf3f4VuX4PXOtUj5fkHOXrLgX4XOuF
wGk25+1V3hPKgl9FQdb4MGVKt+8wrFHqGKkvjIo/re57Y2EVdhqTM4G6qU+X08nX
akKmZSco/vqSkvYTuuZWSHnfI3H726ytPmT7DluwS4lUm5zNOa3WkFc8T6Ej7xPV
4idDAXFhfq9SGIJWBZwSFn5Kcl1ZI3BgXbh6PIcx8whKHULmgQWKRo5Qo3+tRNQD
k891I4FvqR4JVPUydh2WC8AUHBFmhbGCoNG1y+TRMOmgN6fI9vsRERi4Oic6w86q
/NWEtzbe5j1g99bcFQOrrnPM7A96tjrUZUg1A572p9hzTr+lfErccKbBSyjwEvqD
ya6Ba6cF60sNLGX4JEnz3S/JrDY4il9nKjWvnCfvsSah+PyjNEojlJHgQiuq2quh
IX0ZJpnApW2oLwSKUJQYjYP9+168T+ElG7f2/x7lT+dXUNIXRMoIb6SQIgfHmmo9
kg2YE3A/tRUWdw1sXKJeCh6iRS9VTl4cloMr9Ruk8ntFXc8oZwK1ia+gL65XoZwa
7L0IIhq4FsVwtuq+xZyMkWlsnCIjHqLUXu5xlxGnAwDXrabXglu5gDQLywro1Rqi
49OjPP61hI4xkeRZvgN7rTvWJAsoS+pLa1+TWuUwW6ObOX1gpMDPISKmjXY5cKzN
jUzMn6/3LFSwimETHnsBsmeBPuOtjTeS77STnxH/VtTQVrk5Qr0jlcWQpdtt9Xmj
CeGX9CMOpIy+tU0Tlgr7VGzIKq0tO/EoDFDWErKdEHOkOF7warwcJ86v1tteIfCq
s/cls7twlV1/hbuxN/2vVTvF0P6NlF5grcQ4XFCSHTW4pYJI1r93HUkuj2vLZuS3
KiSAEhb5y0EdP55h0gPdVi3gXDUB4xTijlW/TNjQ1SvVW5gWckQB+8lV1UG2DjxF
kRZEOcIKxB6Z3mxQeRPQSw06V8tIKhcqGrZOMgdTEjUaXvI4Y1czRWUbvDTTFDd4
f5K30QkxX2gjsNA87oML8cM8jG/eygv6864+SvLq5Iegyy3emEwUQmuKYm6JQcyZ
8LygpROgptkr0o55VxXVRdFtXggqVvP3COccHcFYPB8arX+5hRwxeasngApCGwha
2tgYs4UtjWmTVyUM4ayxNJ6kEKlcJFyWjd06gPnNom03z6QyARlvZEFRmD7UZC+l
+wmiHa70T+snB4WfBo2FkeJHIlBhABfgl/ioNJ3v7VnYeo0WN4/JpiWrCfERE77e
BAg4rGl4OlMDGG5y4ifNuIbg7pbID3cbXerF4uvqaHWrRgFJrqjDLU253+d0fevz
gHGZefYtPDeai7sKr2SOGdprdUcvZ3Mdvv830gCPP48ZRuKHjFnRlCdNIOIFgFy7
DkMo8ndf3cVugiGmYP9xAamMSQtBYZMkHZWQEBb2v8j5r69UI4/JhLGUq2Hg2Rer
S8trwdl/u0DDGWdcKpvQmwZYyewV5Yf/J+PpXZpNgBcMnyK8si911chftj16qHKc
41VoLsGeg8NdR+FJN/aNp9Q15kvrQ9zKheJEuwaFlMV+mg61F/N3Rt7abvwoJj9l
sCq2+/7uzsuzzy31I2mZWiqikdj1b10KhJQi8EY5jIMdz1S9Z08OIvpzmccNkdlg
uKaYZISJmPNIfL8dkqeaUQfztqDK/jWLAcO2RdT87Gjz3MmzVgyyO0mNfGrpefrv
n2twFB19+X9SJ8R12Yio0uC3v4TTZSIRO+kZt3nryuD2iUYS27Lf+myVdKO9v73p
2B9OD1yTUbf6Pb0vhSanWGb5qiUvMuRlrNixV+ITH1MOM2EbyBr2GSqZ+Hc0/JAH
gOyoLY93/Xkdp476ZCSdkgEIUJ4rcva8ZPQGhZwTMOfxn7ZqNLBeSVmxpB75H7ua
cww83LPH9jwz539Oax3NRWJ9PZlyhihYtMMHyw0ZehUrd6X22OisYCto7rY3UkCH
8jHFM9ysqSjYEzciabmTaAiVfKQlUzcgQkZDnNQPiT9473yEKnd/QHt80W1J7MR7
LDpDsrKyg6blo85Lec9D6dGWghzY3gtS0ErNpvv6aOLOLjkyubC1EVFI1fOswrrr
E3mPcNE7iWY+lnQMyEd8fHgqENQ1n/adxtirTB4CAxzz6cUZHKoTYvZfPH3Rh3ud
9CUycrUKSUgwZHVYrshhBavHDpSzMBernyEVgZe7LKpFi4Zx8ZsVvmgZmplR/tQw
3Hl2YGDt2H3kywsMRMRjRKRZpE7kw5uj56HxqwL7E+NDcmk4l1009+OnOLdM3hqn
b81dPmh/Y2RTejH8CceCAsuiWkVThriQFCO9paIun/T2bb5H4v+bn/ALHf58Dnn2
a7heeVwij/M5NOTFvB4LDFqM8zvr4lXlK++lUFraXg3elwfoy4sx7MZeNqRTC0sF
yeC4VhSXLIXdHt17NAsHOxA3cMLhZ39PZ9D8JqrFgrT+mStnzH97QXiIgEBra6o+
UIYycyo98nKTXa1gfMIKa429oufMUa7JCXBGALO5hvLUZU4hxAuqqmg2OG9DmdC9
UGNqy4onSS1D6ngeHUbBY+0mLiwowGfJZn/CWg5HyjYKUVwaMDV8RaYJuCD3+kVN
MniiwJG2s0V4UR/hIS8Q0tmkW2yejPm2D31INvmtiitga9ijDB5qU+zeTIbKowAX
YrMddjm6OnuGxLM5vFgSrLeoWYMkXVu8x2jrCIl+2UGd3yHSs7FWjWfRBCB7KeA9
agbbW3HnOLOiDkql3NK5S8Uyt2wDtBQRGzLluDyVi5dwVydh/KXHEpECUx1op+Jg
NsQijPqGJ0/ye+3I8j78OqxLSAKnLuvdIIGHPEWJd2K8HXz4GoOCgVWWAK2VBzQW
GL80WDzpGRVyetzUIWfwWqfrLJeKqvE/9Pg3PqJjoz0laAOL5+LW5NqqJdszBPGX
itMCXP/41T22y0qRTFaSFrup/zJABGgqkRzgg9n5QSuvKbRfZsyWRISw1ZWW6rYJ
9JX1ak6C+NNqk+5b8mHmKM+bsudo3X25LWHuGJ+1EIz47IPL3YZASz1N5cwahNDi
IymmzbOedKiRv2OIDMvdj29V06vRs9pIpBf7katpNPHIBUiIbscx2T4nF4XWOHc/
26pMAZD0EflA6I0hr0UYnrpRINrTteCwYyj9lBf9ryVSi4Xz/B3lpGnRI3acv66h
RPwQowjsa75j8eG7RVk0C2/i7WvfIYoZe6Fq226R3dPS4PEe+Jck6+SAIUen3WP1
hBpU0/8XZb4/BUKYmajoQ9bbrhXKJC+KZl2Tg3KJyzVFn/GMpcz8P1Th24+7ZzGs
c+jAZd7ulAgMzHFNHIFkR/5EaI71vLMrpTc6pl+oJCTCvFjranEGkOJBAo8PO9rB
lSH7RVbY3TXzy7P7ASQjYFYzwZiAMH5+hcAhrp1pGm1xtfSGwlGfj6vJRUEOmgDp
87stp8+z2DST0H75KPavzFLQ9SMGGXNBOhD/cJtRyDPBmNqazmLXunpwDkW3dKB9
lKmPYaP9z9WU4zVQu/2PCK77i7BQotYKPKRGxAAWSaWH/fHC7OCh7qPsgWQMwx6O
mH0mZ4lK27429zWfmFO6x0j+FpXxAubASahM9bVlOWNowYt0lizCRWLNGQr/fO0r
43b3NUdnHLF+p6GPZsxuYwahUbUrrW5AfjNyrm1H8v5z0DyfaPFWZfQdkRSEl9Ek
fcbSt6oxwdNavT02z1V2/BtotkYCZwWpAF19rZ5L8zGnsNTP9LAfGkrugivfMcUX
14Cb/fdAiMCn0pJrWB6TwFZFGHx/lNVgTordALIt8y8iyX4Qu+tQNQGhL+Tk/MPY
WKSlKIwKcnM0W2wFQsaVYjM7s2HW6NphYFXQPwYL2WEjtD0KeOxzGfMe1WcU6Mbe
L3uyXyKnPmoplxNEClrVGLulwxNXPcU1gSGWmjMcmergfWMyPSfiuUIyqyZC4Q7f
2IIksIaW8vozJDAzzVzFYcHUmRCCpxoM0nwkJ2DLbZ9RDHAEL84d9TxPY/2nEYpS
I3tOH/tI5tCiSnos9kHOum4lLf1C71Dca7PrUnoGEe525vi3De6fVHFBx/7Qfqqg
lW3z8Jp1JjQBFzquGnbhS8XaG2LqDaUCSm5iZFaivw9UUs1XzJEpM4QfyDVIrzWX
ayukTIhe4xVNsL4Jm0eZQ4OF1yOe3FolG60wQvY4uFqs6AcFROuF7F82+hOJbdTM
8f+rPlQP+W8xKC9P043228A0uSU/zQcmCgd5LqNoV0g5dgwazwEkoeKdJv1j4kUP
g64+pH9G4PhW2utOwxEHF8RIdhGGo6Gr0OhDxHmplJiiWVtoqr6kPT1t++P8Ieqv
owqFmyKyurzGGxch8GqpopnPlrmRqa4khG0vNcBZ3f6NTFHDL9fOfW3/afPMNRdp
1AkCjc7NPbqamPGJTkomlr8bsYY6AgofqpQnu13lRrHiFc+Dda8VuGdx7s7trrR8
PjRnOeYKTdT0NxUC1sIOlTx4qZks9d0tS4zDlnQ7ZbENXd1cnVAAFIxE2mbkQD5z
gOr0UqfEtPZFXAYsMrwhyaQwF/F9pkb/Kl+Gs2d8BZaurarIIAoV+ZvzhvgmGpfq
a4AVYFPtI4mjNXj9Td4s8buBglXa0vJheoKvpiVV6SV6nTIjRgySCrIh2Xz4++vQ
5mz/TxMYfS/UQ0Xcso0V7fzh/fqLzyhzhjobQtpp01syqf7munxyYloPPxIP4Fjw
cmEvJ7KCMrc0WntR2IDBEZcTtn/pEhhTyE04CWDz6l+sGgYkYJ1IdoF8rfok7I/x
A4u+30qycbljHKZdr1UNIC4VHBcfjk7DHLEEM3JfDdYdfmgmMc8imSaADzExVOqz
pF7HEjWmjn19+pV3iswP0wXuPSZ5ZQgk9UCFSbNzEOen0PphZ9uiPvej2aENBoa5
ESy9b931X5/uFYnI9XHgnYZ7bM91JCF2OmhBtAq7bsmmBNFqNPOtHvNB4ojLP/mY
2wf8gfYhIW8i9rZ15UNMJD8nfSt/MgocrEYIeTALPokcZ69fOvQf4JAzGnVE2Wwp
JJ5pTcsIXEbkLRA5iCGE7LEzssME4e7YAh7KNkbs78FISCd4hysBbAV5cf+c/iWa
oE5SGmVmPpNFhu8OqDf6/JHk0UOQORuUHif9txlohSkJlqZCkEUVl4jAvCkOjs8G
rU2/LaLlwYjiGHhgDgQU5OFyjHAhyfIoxYP0p7lgMy60gsFkTWczByNfQ33zMeOs
Y07pmXnmUSDtrDY1KC8MFLQ30PINUD2SKqalb3P4a7IZxkyi3ZUBJLdBMSUavd8G
vdxd7aqZAGpKSb7z8RKhMlcSFogoy/sP/Se7K7LZM/qAEoVy6mEFkUC1Y+eWsGGy
IZolpTJ7eiYHEF6B+TiTPmkZM4LrMNEtGhpBg0WVYYhpSTbaOEgMtfeVXWYrX8YM
NxrEVuMtNsVcjSG5fsqmZSGZM00DLIXqIScKZlhk1n2Gr6/Sbgu9dAiXc9GuJFl/
ix8UxMbKwvA+i72G2DOHw6ctfKEJxfMBg94zPCRgX39cfQCxY18ucbxi3dEJbz5i
axLyqxeIwTW0+nm0bAap8vVsOMi2zF98G2UjhUD9HxI5vHd5MlBa3mH/vZiU64JP
3dyAr5U+husQNqLL6/qzeUmd8HasWsgbuPShcZgDqv8Qve0E/WAMCs5zoMIHn5Tx
PhZeOfNs6sKhBL2DKX8YF+1351S3i+Bqoe+I5UefSUmexvf0wNbti5/kDM1o92e2
S1PuvDhpsmv05mzPdocYmn/hZq83KK33DYh2DwmNo/FStGjl219kmZlfxXCXy6CT
26RSMmJje7gNVTDAoh6x4inInNFJypUhTPgR0W1IjGYDspRE2j2j158SPMPjHJga
g7QG0dhy42HeTZxCYwymhvEq8nQryotRSt7UTqbgbzBnNivTByJg9lybuLk3bXEt
fHdoM9Kq7+SpnAgRPGMovdj9kOO0hwdKN3tNYLg+wxj4OyMsVNHwTGeZqbK2Ns8a
GT3/z3xSV+MgO7tVidbN/6V0Mk5F1EkIpM/1j8lOVYqpt1WR6fvPsiin1wDU/BIL
Jb+jTL4SOKAYh5xkJtrnfYhI8EOvTnwNu5hGmqGYhjzG8fLJJkSrBiemKXFbCL1p
txZJZRAzIxONhVijR3+rdDbPwS6/43G5F2FGM1oG0NwQ9s6N8m9DCP6p1p1dcvUv
dPk3ikAG+eZpf64hwaMcVOROgXvOLL7R82vBK2bGn1Pc5NrFJXLOxmEWxnwGXWGT
2hHhGAJVZj95fX9jSq5KeJ8sNHjhpY/Bj38Nw87CczsL78+Lq0JtwaIoD0TMmCpU
i4g69r4dQPX5al2Nh78yjMbDaTBhGtEmUM9hImSOQ85uCz9caBhLUud9TUHCkrxH
9jVGKQn1N/Ouq4RPlBQ2jjNiSraPSl4VKmrnwmuzc08J4N+6M53uyY9Un5SCAh4K
dDYPuFegNMCJDJmiN7Wbt50EnvY86KfiGGok9F1gilvwjDsRdz6oeYXgGxXrjvtv
kjp/Bu/qiePbCpmZ4hpYssPtlPlT3Fu4yuqJyFc3I3N7nWczo+Ls4QQCNn1Z82eh
sMtefCYulnMEPsCRk5LBHde3tvsO9KXEPC8PToTJeDUHvpqwMn/VT4+ize85llpG
30veTAgi+eTkWgAmb/ppjArOdRGTgM7/WB9Lif19xE6APmUNfQoC6DWZPMRDMr00
1YU72cZS2XET2Z1iuJGuphqy7Sx1hAe8mNww/KrjgsPMzQ1O513WrqUGkRYU2PFJ
vdqZxKs02kdrTq9S5LyeqoTOy6JWgRabQmfItc1GEMxYK05N+wfM+lglHuKKD37B
Ym2kvtn90rB68homPhefqef/wutooQ74mMnQRsFgzNecAua8fVfzKPbGS1Lvu92L
KIvzyzZAeKn8r4sFXnHxDTNMMtfkzZl4VaKUyXw8jsQMojetlOzrI6KlOr/EbaDV
Pw5XHY5z8Q/jzsdPlxkPAumhaDY2BSDKJMRYTBKWJ0UBsxNM+wW/oM1pqa8RJY2P
vhFfx+tZJbi6X6+W7laQktWjIv94wItKZRwU3hZlWr/Q6fooh/N7AtawoaIKUQGC
zQkOGHJP+MZSMOMnvH1FBgH1Pk+2vOkREbyqdq8oLUq5tWeDPlE0dEAGOt45r1tS
I6sj8A3sHWwQcyl9vTERXUPbPa1/l9EmGThlEKIAUQOEmdNE+UZnB1sKSgCqIe3R
G8+bpS0OBFcxi0eZx3r5JQZTpBY+Cm6LV5jdWA512FGou0C6MOBZdUH8aHxmlOGR
ZURua9ZMOrxSH15OG7g/hKUowkRztsNG5UGrAQpbW9dDqdJovqpvhaNf6k8aofXY
2+FCkNY38Orp7KTMLAx0m2hqDal02MqQPyhhQXBCVFATZcgQ4daUbCGguoc/LFf1
io/8O/6kWwIABIRyj255la6IPMIwh+BOVqt7MP6OngO/Ch/8JiNs5sq5ROz9etn2
l3dxKaR7607mbThI4BMEht/t7mUj5X6xm+6zAlVqXP7icWzBNmDRJsf1WAJMNtXS
cISXPE+esdYI+vFcMf+ClWtf6niILhkHKi3bVAfotlvVJKbv88uEBgvag3EO2nOC
GMzt7TpFYJr9mXbwauYB7uZOPLSzEWUTUJNaamiQCrZjx5P9q886wrGIekPl+IUp
bitiAD11T+swT5ndoqJni1sk2jeRMqPPoepRunp7X6icBEIjFYWHsgsiuL0ShXYv
VKfefCe/r5C9l/MD+NWxUqbY7WCxUD0Qb/flghBhSFEqMDjLfzrrXODy431jUl1y
RActkfw4ThV/E0kB6yqwwucjcw7Qqvo/z6kgwnMzxVhn+XJimd8oAtts9xmY0QdU
zNCm6/buTOinJZq8+ZHrLtrFF3JrQGFF5aR6EDheDxBPC9nDj7gRUlEHy8WjI/Vx
DnyUsMOuYYEe4ReOaOjHGCcGY3tVWQHgzPiNLECHdYchCfBRGMxmQ+5GpnKWBy4O
wzlERqp/+mONbdJ6k63Cr7gJ72IZW7OIzvNYqrdbcCwbJNAHSVlccc8k+ooH4KhE
qKvQLh6+pBxFdRs8YBKc2rvdAwI7hKw6uCFombO+zHSTLI9OVtL8aMk/6ih55i0K
EeNsjkmoy9YqgOzpFWuEjxnEEoJ1j6iTvlFMOwcQXe/Vcd6VIVhZV8kR1a6si5JU
Li5eSrs4DZn30wnChsDD3qZUHA9idnC1XCyc59MCPmX45vtC9Zgjx2mKKE04Zkza
kw0OJoS43DCY3rPCDRXd/u1/zUl42fFeo8LHAvwymGPrzs1eiDIHfUk4ngng8WNG
ia6gp2lcfPm4/Ox3oKSogzDWsbrqmeGAoKbvlwk2awUiDh08TUb3pKcQJT8fMC85
hgU9JFY118yVdQBnKi8iTr4CkPJWeu+rQrewtsRuhqCHknxkoelWfI2ac6kdiofl
4s7Y4aoMEEnWgX/RQmWi03ZGLAyd5BISy9v7O1nq302Imk+0YVhUs4bWONbcT9jx
hEWh+h0dJgOvk3pX+tQHNw5C6sICc7winf1jR7yGRN3BF02xDghYj/UqKrnXwzGw
5L3nYyi6UZaI4TQDwYPxeCGwWJieppAIrOjuNH16w193B27OXFRGQZBmeJvz21Ho
kYWpK7kdAbAuY1CIM0Dpv9eMoQC7tSZXvRacDJFCON331phn65Tf/S/G+lvL/bN1
HwpMhUEMmMOCgUd06+HMB6dY392P5cDE23F/+VGDtW8GCFy66YE9+6clKmy2bYFg
6i8YEcI5IJxlyQAwzdz3NzRTAQfnqD2VCrwRRM0FQdvu5uhjLVWMRMXa+DLlyk3h
salUWIgeUHcxYKp2Gj12wYTnQQJBkceNzTbr/7aP0N3vYImFZ+oSQe30xqL9mDU3
THqkyXutMdzLNYJX+ab01hqNFED3MbOnQip8nwlcOe9fIrLGLlkvTLkXuK6yPiJe
PmcCGabO+puZ0seb9JSR+PYzoRJa6dFdhCT5euWXjA57JLreBd/AHyHk56NQcZHD
OvCpNIgrOD7VbD9n0NcuHgZP9bt6Aiob3tOYdFfW0IKFcwWP/q1EkwOCm6Kqm7EZ
CSj/4TrKn5Hn1DmEDNRg476VOuUwngnRevBZQkBYY1b/9oI9k2qCZKiw9Bf/kbw1
oI5E316DceLIScA44LCy3MZfzeEZfvL+UL2XHUwuQcrSzS3SdCE+fH6wZjvbgCBB
oRnO4tm9ztX3BilMBjJv6zx3KYWaJUgfAVoKcaMQrxUPpSzRwzevne8S2WIU4FKY
BToDTPU1V8wDy1NsGadrRCC3+xPGKV0EVepqi4StH8D0+WfKCT4QLi+zkY4ZsFqD
z32q9P2z1NZnX4KYX4mJPP/CoXMbbYfUvjm1sYOmU4A/MizueYJmQ5/aI4/1kyNI
UE0xS5tIjy+f6ybd847A5rJpCZTn3ubStlH2v43C3HAIadJgm1U/OjdH37pr4D6J
859AleugJA6haZGczFfGSEnvUuwdcn9prh7QGvi485C8TMWKQMWgz0b+WGQXQxUi
G0SOnEB2t7QfrJoMDoZLj+J+vySml8DAS+ebBPyrpEmPn5wqepwTs0EaIf7JJDUh
KixkE2Cohl7lEjrhyv97Ao7Rh9n7OxnMhSrhCtBIutvo6xJpDiUy53QnagDJpmiM
Uw6oKqmuZKb7e/rch8pS5QVY7S6RRWny6hiGCLvR6l76Dg9YEx8bjg/5qMqDjy9I
9I19d7HBeMR0MZHyGvOddpkexZnIUsVbvmsHoV73U/7Xga0MGIlAH6aMDdzgVZK+
tH72bunB/htSN+/Q8mhzWF859r7jh12/BEwO8Z0ypFNr3rHAoM+35f/vhqjTDdJs
CYiHXVXplL7LQqk6RQUS2qFXgLAzcbwQCoco1jCQVkh8NHowz0wj/T4dzeAvV2QL
XuWfBGBHFChxXfvXGCno01yzuRTdDlKcsCOa+XJiM2zMSTwmFcT7jxNviAtqPbc2
537AEEdl7mG9c9FHJWfmz+iCIZJpm5GaTDeRkF/jSyBOArF5damD0UGd4u+kXI0w
NKukhvSU7KaefDUu4i3IjXzTYN7NEFfnX0xZXzqEEeJ/B1mjOrJZO7lu9cnW+v0z
9wIZuLY2KjuUuA+S9V1fpXY2aAJcqU38vRLN1LkNge8AkOROwZ+0+q5fATkYORoj
ETf/wqVL7G9hmqtpW2OvQ8NQN4a6kLhqPboZsAbWSeZ8WQ+50jkY/iweR0CB8XMC
rjeqj13ycPQrQuinE2T8xRmsioDI2AICt1qbgpoGvT5VJ2W1LBllx6dbwyJ02R8L
4BBAaTq5U4sddn7xICOd94YUL7e80KynDLVA8O3XQJQD7BTPjJSowvX3qiegYE3S
UtRZ+fP/o8FDuneogHDtNA1nrQOnb1byWCYglrUkCuZsPn+KtkJpgUEcYy0Pub+4
t7yP/APzopTnQyyaTh6ac90aIsjp4Vqp5c26lyFNoXMQtvWdt/dp0W6FGQFeTujJ
wbW0HIB4RF3CvFP8POVvgxoSZGrox9wmTf+PmsYwnCKRLCm3hc6NXTZKytX0qgSa
3dKhw3ETK0Izi9HtgoDyZ9jPH48yiqpniR35Z7CvnTaHCDpnHz/csEPSZXQiGdX8
SSHfdN5HsMP5ReVdGQGU7n0F3nrNw/TAjKPmDBz1M2A8FL9ZiekabQW/gpWtyolk
rphGXy95F+Zhae6heWtQhz1W57UhzpMmK66NPzjAY2NFHqnumqDzQeOZvVkMGJ2e
OxSp6ApG6Fja+3Kabw/uSPGbcad1HGVIETYz3snBqRiRpjmQjIF9orbImUkrxv2O
NxblyWolaRqlK0WbkPJzX5Ncr9DABkLpVhUamxOJcvFzK1/6i4enYOIdoryWWRDn
Gq/xD/anOgRZCfnfF8xDHVvoRVX3eJ3/ZgKK2OaEqymruO74ELOlWmKtbTYWWv9n
bs9vgl575jF93+VhdoN0zE2J4WpXC39ExGdOAQJ5tyd/f5x8yQ9KKVQ7QXucEEdH
lnDcho5OaHoQDyjAUlKvJ5q9nLspKwU6+9nE9c8IKczqXz2XUNZd+Bi2Ip32xWz1
UgkrzRezFVFZ+f9x/BliznRxmhn+1P+EC1ZwFiEZX8JWPXYDi2lChgO9kJlT90SR
SprvHo4c31C+I586mGCC4abRj2DVb6F5gZEViBjTwye3HuNfzZ+4nGuas+lEMQ2L
1pBD3CICyJ9+t0zcwnAfF7BGn8LmHs+aMnDn7mDez8BRh78Rr0FsCNMA35dB6GJx
0motkh5FPs24Ob336PILjcu59CoXU/1IrWvRjysHA7/Ku5hyDFMzBTwGKl+/YGKe
+GRSjhfjLUcBoBJwnng1fXgptT5kMmTyhSuNrYDIrD/GRvtWpsSuuS11ev6QO07H
1hx5ZYqLHwzHb7nU70+8fqfULjt8yCzkRCqzF2K/qzCsnkLH3VZHB7NukxkiyZj8
N401Zihx5W8Io/VgFG9JsvQgUO8eIhebzXV5vj9jOLkX1RM62rpZN7NMqJAP5W4C
f3Fkt/EANBg2BQ2Bkjyu4c9coI8JWDxz4KmpUv0fJfAExIX6vu9XjswDNhXfiXK3
zK0Yi2fF/JfA7WxwUPUx4Nub4Y8aO+WlVcCllZmLrLJfm2yZPEXT4GeGn7jVwnz8
B3n378ehBZk+FeSCYhj6OLtWk+34NI+Dcrzv9iI3JKS87PlJTozy46rkDF0hG5gW
OOgCn3szbfceTCw+oe2cmLqVbz9VniD6N1bwPAa+ynqM45x0CdYZwK/9Z++BoNlo
T0zUPw/Savj1ulIXTDnDndrDO110sMzlBHY4nABZUdd7qyflJmuQ/FOn3BoSbKBe
h1AUnPc5Ibu5a7M3juOySfUsr95R91nTIBRT1APvraF/8okmbRlGsgzp3PHMkAE4
Cn+NolwGf6LU3p2JRLRF/HyblB/wvPpBm8pEZFS6UgslocO9Vs8GgusFSP2gyssc
2noJiAzqrjDggrj9pYiduc1YTyorKl9LpPOKleMxTStKbi1LCm7i/rKJgAZqzOLk
iB0Rd8f+IdunFtNj34oWgQzfm7IVpIRG8cWVv0UYU6lCcrcc/4HNZ/OVCXGPypN9
mdIiQxJUoYARiTsH/YT5SUcy4iDfxCjnlwQuWLLr1gmgf+pDQFBHmp8d4LFusbW8
E9UcGUK7Ejqj47P9kvE41J1PPPKIQ6TualiiZ/GsWHV+XfzcMJkETqYM4jzzEjaU
iCEuG0eYqLfjopuaNSNpUoZXpKp4IFQg7ACSJjcMzSP0xe0RPibyb/axRdph39Zc
EcuCJCKf7KrvKlEaVSMQtG8KurGW+0Ml+MSODVKFUrkZToflPpaEIaMjbpaaHSOM
jmGmcRfQ0RcA5oLldT9qQ4QxdaurjQrXXCrDtPq6yBFhLTaAmF2qwvx2IrK+ePUh
sUgCwjal9Qi9Osbizw1LFSKxXz21yFpSa/JjR5X0NjgGbdo7WjSO75OTfJJRgvzB
9dT0d3HJLbap36oW340ze8HqGw/bp6kzjQyqP08tzPwb/FqpJray2UsAn4+FlyT9
VzWKDubzBC8L0ndaAjjX/nSL4B6UkRD5XA3ucCs5r0s/rK95NbnQ16iVrM/3noaG
i3NoL7dKPVM5p6p+Ev7GZRNi+Q79i49sYjD1uGIxpAta73xO0yUHfYSHzVadeZYq
nJE77HSURgIFF/sipsZNVKX4o5aESgxE82LkkIRK+p+CiZcfFXJeuPHg571i0nGB
4OHa0wa/1ylxdIQMJUArGM6h0kmJ9nW85K9jFgON5O2S8ThuHymGxGYgpPbHse0u
AgPqFfKAnwL22nQmGpBK4MclFx6d68agQIF3grcUgk8YFUSiBX2d1uIK/SQUWLj6
I8xY3LC7Q2wKE4iGYm1tQa1gW7YhiDk1U271HHRA18reMocXqzM74WfLgdaGS3Qy
2gNdg4bhuXx06d1pIakMmkdcJTS1IDgTV6tFugbGdS7hLYI1wE4UIqzHGoyftdGc
JoXmOu9AtrL8oFWNqgk9UtRsXO5Ien0ANJKoZtL7Gp9oXSJVcvstir0wcJ+qaZL7
8aJu0px3Z6fNza/tmwhhXv9ZdEBLF4cnTUGgsZmyYb7vOOOSha/16iDBV/usWci8
RIg1LsQe3rKwU7EeIylSz3+x0u3IGs7FXiAaH37DQrdZ9KsfPp3LdI3xef0yH6Fh
S1FLBYJPofA9pDVEj7iTj+tSQ+3BWRjxLmbCKDjyDNBBxJF5cumD/Ac37xAL2fma
nGp+ouWe8FhpFlc9A5M0n8B6ytWeQp0elM+2JLauuU+v+niFs/BeCxpPKLiQPRh7
GRd/Uz39kuP++P7eISq9LwtfUuSl0qKPBjCO0dK/cRXC+gXJoAyg1Vw8vPmx/V4W
lTztl4esT5SK0SNbDUJox8kAaDws1g0OU7y3IHtMxWs6dXAOgbGLDDYJg3lBEfcb
SU4XwTWbceMfbtwRMLBXKUoSGHYRish36aUgscRJDCQSbmcdnqR5t8pS+XjjMwFP
IskBAtepkc7w98GuuvukrRs23rabsEZcg57YQiYh9UqeSXE5ol82p6zfxFdYlQtI
bNdMrcLC/yhNt6JpRFFXcdntViKoKzU2jmSQO3aaaSWF2FVvECJo88WFoyphFCKw
Po/PYGJlGwywzkrEhA9Pu3NcY+ezucVb57QSVXzW2V7/CBeqNM4+QADyN5X8Hle3
3Syp7gM/lwgANT9Pp9YHdO+u3IN1/wCWftzQMbmnmBc0xGwgisCVGZgYFbkxwNxQ
D648WG184ULcyzcsEY4x+fI3ogEDXJqjHLFIdgipcW05qAtYJ1OBFKMU+JuqlMb5
Ow2U6jEi1qBU8SBYJox4tRPSRobTIYLbQhT8PxQZB961IszvBPHjGySsRmuXF43+
nzXZTRKBN6wMB3ehuErWWkWJnUof8vtV82uZu9rpDbBlS3jrW+DM9uvAx4sc2A0m
/+ahLph6qw49/NfRCTLTQW9nmAMiHTwLW8rKzBXKRf5wIJR8o72X7mq1bYTGJlQE
3ZArfj/iKYEZ1U2OPxzH2kvGQOAueysbzyHaPAD4j8zcNCIla1RKuNb6eEZJLdki
HHd/US8aLSBZqWlR/WY6iQQ1/1EpeejfDfH2dc6gpSecSCC/TMSZgk6NSFZ6EvoO
sNPpDtLRF0THJ3WzwvuEWRkZCpnRajilLgDigCrKICIA3QdV9lVY9M/KjU5HSBaN
6ViseaEYVx2U68LPo0M1RTa76Ltrq/Y1thtw7e4Lv9v/o1BpsMMq0DhyxBhwREI3
NmKWiGcmNIzSQvIRXG1zppb5yxfvxIdOE2VL2yYBqtYCJeQegfRlSLB5Ai9NxIHm
TvGfbRvdCb7+kt855NILqt5LqGuTi6m+/tp+Zuq4dRid99Bm4wfYPMf4g2W+OUi1
VW9aOLy5tBxW30iH/02OOz4+sb5BGrotDAsC6PApb8s59E+fwC+FGQZLljh0zh8Y
TGfAJKt9G4tfNx5dyM4tD3XJqbq6FYav6OipUB3aAbVlX3VJMySBMxNSMBG82oO1
QulhzIOWHoSte6DiGlt2dEviGbyu+q9U0xfRSNh485f+vbJe2iO+kBcA+6fl0LOz
pshwy3Nfh+ufCyW3dptKl1+96MPYMDgztUlGFovWK9uIH2Utxlwm/yoxGkhzgBzy
huwSnTmzxX4uHV2hz5re5dYPCBYT3gjG2mv0+ReNzSHNM3Y2O/f4jHKjcMW2x8b3
p8m1kuKEAQZQGT1xEgi3Qk50yFqQcie2eePO5ZrWKK507Abia/3tscM6Y6JaUunJ
jCbL3IdBphnCuwY+MbPXzBy0wzpPqfoQCwBeHQlNUIZvmDFrGJZ+oJLBEH0syxK9
/u3H7lK2YXaVz8+LKtsN5oWWP574bDhhCptag6vDjtOK8M4BJ1Vhxm9r3WXzE6mn
qKc0c2pwyxFzcdWYsAv41y3Rjtyyl0CI0Xi9dlBZoML0pE6uI33G9KKXEGq5ph2f
ftPltlZ6FFItuYmhmG3BFbU8riqasryIHXG8L9gcKlvVDODJUw8/5W5ucZDP0oeK
XOesbA2wBIqKxyS+03KdeFInFpUPWnpUDG6cKd6P8qzStU4KSs4Z1dj3xlmCfZiE
a2VXK8R4/ypYBzCwv81fKyDTfoqqq+ZL8XDBk6WPfhF69AWkDpyflfV1LxQitxz3
H7Lp3MV0t/gAQoBUv/dgSFQLqJWK4bdpeNDoSzKsR1NXNBLn3gDJ0xqdaMBukwjs
KK7U+KP3JTLL8nl2ScZBKB2N+F48hmL0aG9+2o/T3bph5sa4T5j+i5ExNlYS905R
rzlBvW/hPurzWyqPQ6Tzqk6CsCWdzmlCisLJgcLyHuW8RkI69KXDLPj29q6HgDFe
D123uF7B9QyrKczlomIMXtj76HYFcmud97xK49JdYAah++B+fLGdJbbn09s1ZzKy
FoSHAlLuiALbepiHHLWC9jmwdkon5zoXuAd/4seSNxeX9jYcl6Wpzv/lJSPngm+8
5Is/kacZqLi5M2liajWVhpjKfqPFGYW4P1hqG4hU+BaG0aMI4h9AVgJPNrxlomn+
mwhP+Llfd5JQHH92KN+aPPuK5ATdP2bgGnZhnrz2Xn8Mo991+PjKotKB3xCx//CH
HiafUIvFNoEDTvnkIkTN2QUYfQMvftTEqRW5sb0Awa6zjSS3wCjCrADgxy5LCd7/
WaapJl20bXUlhtBnq/vrVFM/hzzwVzE42rNaCvljVEIXhpd0JYP0bS/3SFp5P92P
tEZAdP5CUYJ8qYwTJR896iMofw37DmXxRF1ZCDhg43UQc8tu9F3z28dd7/g+mvE7
EoAqR5gSd55ShO5XQ0JY/+TY4U5VdqL3+/uE6CFHA7J4OR2w9HuzonWAMCHj3j4P
kT+/EJjpNOqWAMHJhiBZtQ4pd4Z97eEDE0bYYXw/glCSUMJQPIBGFK3mcq5nDaj6
tcPYCK5ObU8XT2GUOODuzvKx6lhjqmDGC228Aur4JHyeZrlCsJu9VO4itL/BJtxn
/r/UtuvRjy31yrt3u2DHzzehDnjihYKx3oZ5TgKXgFXPbIeHrpgJ9o6qwe1s/m+l
qCDDKNALq1p1ceeKLylYJtLxBjotd/mIjhur/7g1+S8Pcho62NtCT7Di+Zg3l686
wVin+Dsi2DUlxKtgwkTlZK8QFNecgTZRuXB2d/UIEXCBukjCKTD5rntl28g2Mbux
5r8B/stDBCB+zTU0eRq/EYvsR6QAFWLZTFsV3q++ISWKEyd/NYnyNFN2SxbzcNHF
tskCFq5YrJ+YJJGd4ITsXkAtU/B8qtf3+OLh1lGwj9Fsyt1p79E6/E3RA6K1z26e
i+ceEQQOV1LqOCs968GzO2JF4Mzdd78dN6lIz55tuVmUw4Mk2fIzbzt4JK0ak+Q/
ffAmGP8YWeOeERz4XSUdfWrCfvAo67DTPNXyuvYX2+dYAoHdTWdBCa7wAvF+6R1A
kWIDkaNVBmQQLOiRtwQaEjx/Fehh9Oe268lKGZ2vFganh9dFR4bawBwnAbvRlRgQ
HpLC1Z62ZKiBYrw+hRqZN7JdLEZ8hGfu6ssnVAWTKbdW6dJAIwbhfb0LT8MsCYfy
mMGSZjbOZ5bFYmixtJ14wbxjUhkJlVPC3xJqRJl2inEF9X+RHErklZoIPaJETjoE
NI98pY325fwGbumPqIIzvq5h2Q/3gCLtLbmsK9IXthpeClzndYTbmxFm+woFqHH+
Sz/Cqdl9fPFfy0kZLXGc63Ex9/xgBouxrRwY0FgsmvZcVEhSfxYoaokWGDG5IdSB
H4ewo5MQEo2Dyj6J0ZDgq54GULcprMbK5SBr/zaaPYUBHmtwTjEJOy+mR/Ri/UQ3
fdYWWnS0Z97jJALW77R5cNsXmGeBcGLb7pvuHDT596tXmzkEoCsX6jaftBa75umE
KD1vZo/NvIZ2dD1oHGVUxkxgCagPC4sx5lhRHBLvFaLDxs/4hO7OlE9Q5GMJ+G6O
TBe72HTx2hV/1zAVg8aWjH1YG7BzxC9Z+JmdK2VcHZdhDglioig6vZuIRt9kvWNU
HkyjsLmqOIugEpUmpte/96fzonlOdkWs4rNWTav6asqNk4KKvoXHcnKrNNGl+yjs
q65EafyAg2udH1Bm4bG7CuEwZRDB3XzL/ly+X2N1mM/cqGZ8BjYw2wpAJO3Nc6uW
Ds7CN4nA6tDVlRJaPWIrGCOitOmlx3I/vas/nSUunwrXZkl38yrFKVhmYslb//pM
oD0pehf4UMqm0xns0VrwaaDQ5Nv6gR0zq2pAOJudl92gulwY+XDr75R0mfVd9Jx5
Z9jFmeaXE0UTYRa+zk1+wnLk6vwKPZ5HnCVbIWrwKhv37UaxpOysi8DGoXjy5EGP
MOB9IRv7cyaJC0qxq6BKNTbaatgIe8OcVAnC3ba3PFd/gvyUpG2lmjyX7c3wLyrW
jTcS18CvUQU93iaWncwtxLic0+Wu366YAxFPhnm9QfaSbOyCD/8u9IY7d0kMDdNn
gdVxDM+Hbm9Y97qQLXF/fzEjrnSiwvGe2B6svJaqvv4GeYX4vs+bBlejrcvNSB17
2wJFxkYmW0WjawCm+WqCnCbisGbL2jXRtLfQZlgjnoyupAmz8iBz/0wusiTeR0rj
gvGvIJ6kDnD+TNK8zohPCTaVTS7THLSmHqcf3x0iPBVVxIBeakwnHKfqbNaKAPGA
om7Ctv8Au2q1AUScksb18s9w1fiPxZfJPwwUB6hhpQboDrcwsCkx4Dg/4cK0UudU
6WxcfKC81ig4p0tJFcQzLr0PbBsGEHx2304kEJKOz9IkMa8ooOyG6LDI3HQwVoPu
RKNfs+dm+3+BADaHHeBB9mgjwH1CfJLgSF/IVRM1qqvgnPwONpcXNVNO8bGrr7Vx
ggXMNfzAZx0Uzdqs5asTJvnb+j7V+QTYiyn1NUb3sPPkfFpIKanqrCnGna/ftOL/
+Xvbt0q2DxXmRArnuNjNUWNUMojcqLd4c3lOSLzLFRZ/SzN1w2R5qOHkv8AxNWaQ
fINmE2cqmxh1s8pSDkFq/v7EdSPFa70hy4yVccRwBAG+gpSPl4hcNFxWiVqwcOAC
wewctEReCnCpSfb17tPbrJCFEkP7XTym6ejVd+Vech0A4LEu0fgxFn+5rN3vemWB
Ll9Cucee1ImhPgzdd9OSX5FL8+VktY13cCkkiTSrVeCuwRp0qMPhIhqjNOrpnqbT
MMXglwKXg0Phzc4ri96zSgIDoulPyfaShPGCAq8iiI3BirEfXBW5sVXWd6Etgg1c
jfzAbjBAIs06/OmpFhbLYcav/tEM1JV/VHS8IF8rlhNZJum2prI7cRvT1voA0bPW
JwcTY1S28Xs8xJY/kQZSU3MHWXPytWVjKAVpm6QEHZKz6/B5UuefghGQR0TQuVDP
jdXREZPELARqE7NddQhBnxkOR44IwKpDuvDWkORX2Ntliq4en7gBAGAQ0Ochumwz
fY52l9tmWVK1pVsU4Zed8lNQI4UD3xmRDsN7j1vNaMhkWbzJku2Svj3wO4355vh0
PZB9wvbsL0pb9pfsHB3B68woMotVgHpaRQOpBlxHJLKWFs+99iSjq9YAzOkQj4hd
kB/Ac43j+ZsCtJttFu16A2eN44DHLljHqERZVZex3YjgDgMVeZIc8l7pe0uGKNS5
TBmNXnjADRwY7arRLIHS15OWzxXeotJhrS6abGu5l0SyWKDDmsizy4qHyOk7a2A3
oHH8ZBLlc+eTb970hc6Vbrd7swG+CwzNn3O/EyEko5en1OpPBx22jdeaMx0TpZ6/
ejTRmfYX3n0vXQfKzOsvT3tjcEmBKGOg1VVA8Jpb/cjecGJ88B1gQgrhKf/6I7+M
NZOoVXMm1oj/UtXCGMpV/oaUvtSsYSVSIgizh/hUnMuEUa9QlCHxD979QIFolzTz
D2KGT1ZXgr1fxW9vo4pTkIUWUxUshuMLbfBenGRqk5YruriLfEuevS0ClyImi/G8
k3RhwoPs43gpuWrxWFs7O8b50aBp/A2bUgvBshljZa7VnnNddhG7xVqNAPyXU6dl
8nOQ/aHlnGVPUveKaRtIxYYlt9844tpvCUN9fF0/mcAp5Q5eTHJnZO2SfeRMz1zP
70pnyo6kZ61jqaGcWtAH4ailMmvwj3tJcILKSOo1C4oK3D+o7H4kd5HeM1uVoNJT
rH6TQuFxfhKi3nh3ENSgkMapo+HmrRtqqoj0npMU+oNwQzdwL+vlrxg+f4gqszai
XhMLQmxtjS6ahI18eL/aYiciIh0sMRwZ9ZEgX6anGYDhCMaW7jiPqfHGTgrsAI5K
1gJ0JMa97bbhrZXs+2EKLYnKr4g5k4kOSzULmm8LcbIZIsO9EN6vTXwHWf8YuqX0
M401QzKsLUM7XZO6bPmngWKNPxK/CWo4ok1tbE4FIoF7HHQSgr9Hl4tJlWY2MI/F
/fyTaqBY34FBUJv6+TL6CqCVo1YRcNn2DMA/MvnfxjKsPapf+WVOrNsQNcevUmdk
XTWBJzHbx0Qd3lx+b341wLF1IzENyZZvLSmHwwdALicJgSuLtycwC8zrsZYIbaZN
TRQJaje7qIyKjov5tCb9qmux5hds7V0itpogA5ENsWBuMmSJxW6yYi1mm7uroPC/
VJztdPhhEtvuGJT8eHWNHe9L/eavmYXT+eKj1zaqS4R96VkT8ysAWCwH3UwJ+K0s
rts95F+flP8m+9Ta1/MVngR93czA3KQB6dV5igODQFz4zhk/DHIooo8NeJyr2ubD
gLtMLpmOzoBdX8O26nzpvwXbGHVv4HlDYcqcmVlxDe6EIqvaAI1wtf3lTSs57IJ/
TfVh+sHd5PYlf+5nKvWlDeEprBznNBdU2S2p7hrkbNqr9Y3dNzA/VdEXN4qc051d
HNa2vMh9DBVJB1ctmd6V1U28EcpO4eGhQ7lpv4di338mEWMdO8XXVZaYZ2J1RFKb
r2Ghg/xuv0H1Xfh81iF2SNnZDIwcGSutuqxYtuzV5MGzO3BHDnWA3bSEYv/ZoYau
MgyeoLrBO1dDSNmWHAQximx2fkm1MJv/ys6jKBQuuNW/RQONXqL/Nfs9ctticIxz
gvt3OIhY7oeaUMMEoN6vRxwkwBsjSiJpkaROdqYumIOgmY6jJcQMSAVVNYqgTh6z
vsmhipD7/iRk6IoHbO1l0erxVcskigsLBXKX+YSc35S9uOFs8nx3s8cvCncVKp3j
o1lvejxhkCVPjatQtH6sMN+paFDyJRE43iKdDzXg1DXgwxxbZv0RWyvaGN73pPUb
eBsns3UqvAjey2d2Yde8mpsgMpZY8c5ZHBnnqyXWGHaxGrguzLEp6Fp19ql0hRen
NS4nVo55qSiIelCyfT+FnjczVFVxnTagIipSQxmXi5ILKeBJq1rMJltlvTXY4fwx
ivo1CWIqbDOG9k3stkVnpPOTmousi4xLDniZN7q0l0gXTvrNdrMeFleKFgDEI+zi
jyyCV5bws40gATWz5gzshazRVypbZUmAoOcIQ1t2jTbi3np4vdp0v9vXnZkK8pop
QlzGz2NsZd4eQFM01KXbcOYxL0lOtGia/gHCWaCuxcmjzw/3h5TJlL1oEqLXkfH/
/oPf2a+4awG69tM+5do74vor1yebS+qgzNTHytudtcqbgTmE1iDSd0m8eO4UAzui
KXfnOsIA++2TuhGG85n3GaGF5RkFaY87z4NjNnKfnrCftikkxPb54/093nHWPe4V
RZfek9TAX+kg4hkk3HzxAa3nxM5dmFNHpwTb8Zbs93XwiowHzzxFEmucLWNN4sFl
TldXwu6xNSlP3sXFMxXaFavA8+W89HFqFHRQPaXkXalR55CzSdy8duQK3qqejG8D
y/mZmcqN4AhXXRPIVTBZuQDdqMHGsD+981Yl4+N1XczjlG+foNBz8kcPPRNcVYLG
aSo6Oa0uHXFN5O7HTxLBSLfzhYH9tz9eSLKs9PpNiwbJ3ouA/BgQTJnbJUC7Oc8R
GXmiqzelbOMW43eLCC3JOvRlXwdBX6DarUAcoCtlVQz38DMIF06LmudQjvLmRUN8
pze9y3/tHopl42PnP1cJFBtaKYIlpNKz0wKjWQFQBWbF37WimGB1TYGtuL3Be6Ph
/2euqt3tyXIpbi6YMohvonE8S5cbUinNvdz867SH+rIRfoUOuzOA5aFEde2UjXkX
JOXqnwQXXobasOo3EiFMzjPGuv4fK4LkBBxqTD21/RC0zfKhbMn1OJ9r8fCQ7crQ
yuELrrK9MhrOIM5t01isyQiTiYA3/BqGNR+6lE3XGhtxI2aDOfZv+9xbEa7KHi2v
5xCUx5Z4NZD3uwRcy4uSdIGN15yXIXH0fOwiXD/Nr70SwBZVn+bY59X1AyWGkt2Q
4SC59WcaY1XBU6lSQBDZLR7sLCdxoadnyYCh6PL4PJHKpr3VBPogmZ3yLbuA42Q4
ypYZkxkOPkEtpltWaugqiLWSuzSFodVV0l/kDtDNyMc4qJnSaF9ZqhcwsiX6foGM
h+r0xW8KK6OMP65YDRbNbsouk4lVOgl+meLxfhrPWlQQje03AIn/EzTdhgm06MN7
GCjoAyR1cDygFVp/+ixpzBKFfb6ct9YW24zYzJJE6f8bYQgYjlkNPd3PeSiCn33k
ne0O5+R8gJKePzwgGVqKkcntumM/hwafG2wgKLHCoCn8zWPHU9q2u/xfWrf4LnKj
rzQ7EKSwz4ACZP7OcuN09x3qe2gw4mxPZ2uQJdOIIaFbVk4gXd/iVWhZE7LD0sgW
N2ihW41lusVXOEeo0aM818I3E/KL1cNUA8vyMA99Jc4n85LuFQ7x1ne7vkl0oJnt
Fm1dn+kFCRX7nclVtmX/x1xAadQFwS3lV+M5ggaVKJ391fTLiTHWrduVGb+CWr7d
59lZC6eqQRwBI1MU+2NfPF3vDQlCFqgQZ6rZY+7PYNOSYYoKsbxEK8znEZDGUpcr
UwZhJ/WOSMZTCOtfDT4xuVdzoHld3x1Pm/TAOdTctrL/LOu26sCwgGq8Oc8ENnIM
+J2ikCniS9QFHzqPfOpu8Vni+MbAbUixdiLBdJW8k4jxA8eZ2qhxuEt4WMjhI9NU
ei+MpBtFH+waZNvWhfF/oxdIAJ72a20yjCZuTTH/IeViswxoF+deAK/DlEPMSTxX
z+RVREirAbhW1YkAxhYVQmiHtcOqx0YZn3MeK7L2oxQNONqMbfjUdl4SmvDlFF6b
KrM/BaVFYzZjN+u2+v4MVA2j3jsDo3V0/BKsjovpQEe5VmA474bLxTYng0SOlI/O
FMwrx1Wb+6+qNDE04s075sBduHoNDb5E05C02sJk/cDqdce+nbjmBtGRSp7xXuPp
XOAHAEtfS4Ux8uUstIIi5ddTYTaeV1vlWLxbQjVg+rCnQNIZIWFLhYHh6GF3Gj1o
Fct1lDeOd/D52Y8jQ8QM/GbboiGJL+W6qyirzvhSiZnA3W9yCsd1yiLuIcY1Zs8c
5uS+Kzk+J/4B2O7Elqn4JvgJWsYcxLper4VQF2VAWoIiRRxrn73QErSaYm7WVyUA
PchzTZ3xVY281E59RpHTUwt5p6zfytpBt9cWxsRb7X3Le/qdxy1lhILqO0pa3VZ5
dLrI3HgP2miL3EIm+nzwe3iwIFCig78I31tEOalEf2kW/7BEOt0jSwHwunB0Vqp3
1FkxHKEPK94o8t9ThPB2hiZEeIYhSHOZwXAdB7gJEvm8ogg0KzXOKVQ+vaTSmd2+
x+Q1P2W966tLW0ia5hX0Ne7eJZ4VgMTI5Nfh1umnnAnL1dfPp/ZimaIZfg40RJar
NfbG40vdJ9NZeOdITrF3ql622671mxzc9i7Mb2mkVmvHN24kpEFNIs0XECJmv0JC
QKaiSmrOkfnvMnAVzB4McJOFgRVfpqetKjYBxNsmXIuSyDjbhkv89a/VlsVzqROC
thVEThJCur4vQZgIL062PYGLdvopQsBNgBtFotwdcSWktqLLpisEFsRjdA2bqRVc
CNJMBuFKmLfk9XxU/3d2T8ijNNE8vEIeOD5iaaucAhDvjEW/0TGI+d4UdWhy6AZL
eagYRHMon26QNIDR2PqmL3kE/k3rdMRm+/uN38zMudNESY4tEWUuUaNIWdT7GZO9
FEwQh0b4ZhnDPe1viQcOZlY42uaRiYtUfwDPbpokm1kJAAaPujuPsswcC4voArSg
Zd/Nxrg3t2gPtfA3DwXMJindRZIhvDT9mvmuAO6q7tXEAKD4U2gaFZ6aE58LL9gf
XdrLhgufvJOMbVncMZqGXBg7hPN77254HmsoOmNCRN2QWoWHOL45p2IHI1cFbajA
aJGCdflFI0iOEr0Pp8pTPmFV+b1Xq4mgd8nVTWtdSZUXwXjGxZHLzC+JoKBIJeRI
F4I+MC+acEXkF+ym1bcoxAs1HVKpAUmZHGUYWr9549b5ix6helawJ+fSVJ1pQ0i5
xTnNCVT5w/IMxcCMOBLv3CsCCoaT/wZ7Luy2/nMcocl4xK7xuGTdrxOTiZeLR1ru
owG2J6ThXNxQZBtdYKNGNVMaivpfdPiHIGx6NQXaSzCXuIJK0u5D0cdNQTi1YEu5
DTcrNr0TxfJq/c5Txc0gfcBIwjI9iuZ/xkzlS7lFBhD/w61BGsZwNnkC044WGxbw
qZ88HP/UBSG68Ac+DVN/Wm8NRikA4T4ZgsxIltM34dBkTuWTuT48mPBysAzzoeKr
qGMDpu6CSDbvcNCO/NOj9Dvogc2Yuw0XTPQB75iW0MAy+fZE0tE7+2XTIRooSszJ
N40dCyDFh7c3pWpcCIari6drLiTE/JZ6mJXe5X4n02oTuy+MZ0xFW2EtOXx//ZgF
5R7BRBrvCFEaROa1V5aSHEKY8S5/qO5STQBW26ydj6B/kmFwwq3V9k37RqPf+AW5
k517OwCU8WDr6X4+0BlMO3SgajjBQ+yR0RrM9Azjv9oAftNXW49vIzMW09CsiZBQ
q82zS9laOMvIOYoqxE9X0g2xeVAkLxSVfxYceC6glcwLLOr0fZIcpZp2zxJxrOqp
z/h1+lQvXAJx9JUyUSeHO3EUTd/Dc4xJO4b4fgkGvFwxJxFlVojytOJnDtKbyHY+
S03kHzKMKiXYGhIzNeQOnlO5yIXaApRABlVAUxPfFQkq9X6/58sSOn7/Ad8wpLJA
T3oGPVgHrklA1GVuljMpZ1Fiq1Kiq8uVPUQf1tsmmoGD9LjhWzoA2BtkyfV1agw5
5EdbJ5FSkzQFXyfaZKcqsrqBq58WuCmkN/c0BzpuXYw0tP+IEZbOtM6RlQaIc74f
dcPp4N0l2XKNA07xfGLYLqnqyFEx3/eHXEfFTdG9OIk9oq93+DzIgNdnR8ZYHR0A
gzbVZjaKe+mmpUrzpB59Zf4zlJm/1DcwC+OUJXlzutLRl2/iKIifR5NOkCJOn/Qt
UdYqTbd1OVsE0d4c/jrFWqnZ/FUCpCbUC1zO6EYQef4AblM4SvC0BB3orbmar5ue
Pzly7L8XLU0e4nrO0NQCcrIDF2JIMV01iDKl+YyQ68LzCQiH7OubmSgUKfezt/OQ
y4QHGI/PYlCfv/FOp67ez7JVlCnI+vVvcZRRYQq3Xv3HMFkFtoXuLMtrQdZEJsyE
f1Wko5DtkrBY3hlPDLjybk3/Ii0FpWHtQysAbwhd6AuAZ4dcyEv+l4o0etUlMmYZ
0ZdOZlG9UfXGtaylprrC9JTF54FWw28zCtK0Eszh1l66wjASedxw3jFoqc2lW1Ef
qlGf7zrUm+KRQYLkpsgATyFA34MoejjBVVcjvXxdvpP6lXkQIpa4v/Bb8/DLAdHX
BtpGJbxZFIdgNwyB1YuoRo6hWnUkWl+bP9nOX7O7vvZWtrqJnXuv6GTlkwwvQfng
0Ghfz6E5dRV8XLGhEn+NJybVJW4OEo1/32GalTE6GbDweRb5qYDwVnlHlvYvCiJR
o41KoVycxbXp9gqSxaz2nB6Uv8bbh4Yt/cDxjIevnGhhe+rfAiixvQebn1qGeEWv
S0jKiVnUyoCniqRaoVfeyJruocIPbgMnYnGRbrJ46Pw/5VR0Wn3rS0Gbg4pjxcHS
jAvUpjr2Rv3n6W9LEDjRNgaZU1t+QKd6m9L/asEA4y7GUfgf8efg9oAAih5yATXE
KM6lPBIVOnE8Ro6fLWZn8UjEfCHihYqKSsnMCKYNBSEecIGB88e6cCE2215R6ZC4
46HM0+MpZOD0pxxEgE/SO/mNUnhH9YI51f/XAu2bOYcFEl8+94qYiJymIE7ZyhN8
3VkPZSr0l+ujPLXQMh5vnD6Ty7smnkpToHLMLGbfSGJRKeIa/+PvRIWYrA4i8nSH
PA4m2VB/p5ac1EOPvJyc1YD/U1Xnh7+HQ/VAnLZDUNSoHSjWlz6Pg53MYSN2mrjg
PGRcp0NePSyv0ax6QQoKZ58KuMPXpJ9iUz+ZQYdWT31MXf+lilBWsT6HJqosKEV+
1kZ2txDzCzY7OjnNx4vGvE7aURSUVPTLxg6N4NLEv37skcN6ke36uZlfox5IAt3i
ow0s5EIcExnlsjivy/5Ec8RIhSFlrmpf3Cn3kPebj2XSzrs71B6j+D96wzM8cGhO
L32ePU+wO25+IXSEQnGCy4lkLTunA7mTkGyp751/sF4vLw0AycOb1rlmC9KnUr04
9WS2LolrPSt+4JwO75jt4kZ46/so00WtaowUjoG6OvptyjYLjcnY49j1vqev8U2I
wiDNnhsn8uThRE+qOAIc4SO0Wc7ysZ8Q/6HIzj4ZEgvJl5P35F0IDuynCDtNvfkD
JbuHcs15kj/CvDPs787bNAVg9bnkT1Z48+Y/Bk7tFlSu2lfu9Tm6KY/WIvNq0Zmu
T1Zw2FNGgQKp9Y7gu8caFvW4IW8EUQoHoQCsphrEaXn6pp3psmJejt/7Awt7H/wT
qtL9SQmWDr25dwo6N6aOCsI/3OauvdQLdOJjBaERM+/LE5vp9jBy32OAD2OCxan8
r7FM9IgTe2cHJDf8Nh9okE5zZMjbRdT+xNHVij1hj7ZxRXi+rw0JhbhYZQZO35Ah
Rz9f3iiWvZuUDwLbkOsgCCOGkX+THx5Tca95YSeH7VkgSKPHNXFnctrpraH7ym+M
BdV1HyqzWQT69WVMln9r6SElWvQBiExnTmQyDD4igYXt5cc4QpN2DfkVa3cZDbs9
fbjU3VOHLVBnrIzW0z9Ut1UfOee94vNtSv9jG+nQMdVnCorYFjPXti3DMsNVyiup
N9uxiPG9SISGp9iFoI88pn3UHkbtcY/5GgBQsc/KyxXsopTo9DWyZqdN2z+pPBh5
+ujjvNNfA8dLmFJkF/wuk5BZHF+2cn7usCEpi2uGAkf+kycw2QwMtwKdQ5ePdpCT
ld1x1ll4t3hgLi7ThyREki6noe5m9W6XPCI2GkNmiZWrL/gBXDopsSHhFYj5xv5J
LfscIOD80Bp2utfbBzDLE15Fkck9G+uGn62u4lp1XT17Kuj8OAqBSGymFs8otMgD
Qsik7riet8S1IIzK5BmA1FrYvav+gyU/qP2wkgJor62+gCaKocvBtJF5zyYWIyGn
sdMHr4AFCao6AchvtPWNkRzwUDoZJDxoknq9XKKY0zTzMb5Mj/7iEJ2OVwIvTc/Y
5FmZa//dNq7kMUgbrY6bx5sVgmny4F5eG1V+JaCwhghFl/+LhwVtO4XyryShqWiG
ZLjdtm9g2cs5XMOy6l4VFkKYEjcGyKk5z8GUW+GsAyth+xoqbPiPXTrFzNt2BBFf
lnNRBsdJQEob9en4laUwRD41aNMq8W+VhcB5Z0YiuyzmK+8atZUG9AF6wioTJH8E
XxhGQP2dubcar9gcINVkNZI9ZUnEco0jg325lRLq9gbKkCryHnHYCO6wTJiFaUZN
E9bp19Jdx8/GjC6Unr50v1j2R17SMUckxMqJJehXTeZvvIUcrLzm0iyjM5eJVc6/
BuzbKq8QXuJJU0S3YrlU2Dw6VGATlcvPC+TKRPnCbgRvc5XsLU1lflVbkiTqj2S7
G+5dnf74SZbysBkLBFydiOY14wVtXxDg9QAFIHUBMQhGuW3yVeEx+4LO3+RktWRe
ow7StEpXIc2itQu9EON6bZazpvP+OfMhgxOA8k1xAnBUWqLvlqplyiyfkF7qqxII
wzdPiuArkWPVUfpgjhIxuZh0j0MbT0clPS3MFK4ZnY1vjGw7blc3gZ33PMgu+HC1
UtXxQRhb6wp4KMqe+3vaToSFCR+f/D3tD7Trxj36lw9lgRtroMk+um0KI4mc6dCn
KsJqAQY/UdkOVCuClJv7oIvMy8o1+njO5Xr0XGKZjqcWvVNdGb/gE1N6LHZVMMTv
owd+bU4Ol0y5Da5a0ryvMb8B+laWTrFiuY1c5xNzNnAksMRqNq8pyrqwezilZMkm
M6AB9/3iaY82eTH56f8ehFVj+9uzlxf+PkeGDFHtVdQvnuBJSyoPc9pAP/6IrZPD
8rrZX+jaex6oJlHjs+jVVxOv9Djaj1HUab/H1SWsKYLkgoaoiv58SNpNm0oJXFwH
W/eMBvJhIRdqL77eS0tdlE6R/+ZY/rjEpYEE+Li+xJJSFz8ktzJ57Rukcj6sfk83
6hO9Jm7YWxmAp7PlCdzkcDp7KZMzIv+UfUbhPNDYq4ZvoFsrSXXTYfet8sqkUS4z
D8y7r2LQ5Inx7dV0lbG/afH6cAaY9ageR1NLeGIfF7YanmwwPF72U9u0sjryGVii
9KJdSncR3pIOK0JNSBkfBgG4ipkQjc6J1YvE1lGcdl67rJSZ2Vp5u+MT7GqbKuYw
WAGmygmNtu59lYgkT3wTU38xJheCr9rFmJ3w4OndJkBxlFxK/8sxyRLD3lq7VgMn
P3IWJHw4LdyhgI7djqMvmRYOrRK577dCRfFiU+u0RH2fswLWT0uFhkAALKHgc4H9
EEm7aIXtikY9Z0wTrD0FB40anf8Z18QVBD2ESbd/Db/MIi+K6pQaBctwrb6UkSS6
rme5tpbmbLRThmNtTKQ6jrxMANJd7jS2neIC6fQRi1N3/5wbNcfjfQYb/rDUHQxi
CI59BY8BwzA1Oz2QEthHTmtPuWx543XSJee+nXP6mShDsngf7WwazP2DxY10P/GF
F5o60Ta3Ki73lDfuXCxn7uRk6ZL8kTfPBQS2Z8I3yien4cSToxc1uSrwvPPqVUCp
APoFEGroTBQs68K7lHXI6joXUxU4IS9J1f30VT+dzKXIUmTBqtoVixMN57fbfrHG
n/HgI8mDP1iA0B18eDgzD7ip+kKL7KX+x45Rt7lA/atXG0+CQxNO3HcG3j8HELFa
suZcHhtzEbWS3OZIMjlfUbVjt9tIBb+WottzLWbSldZZ/vew6Rd4uqizSmrLiTcP
9TTrat0C4dlozJNrd2zO3+a6c6JYBHfvRczPNcqrtHiqi/hB2dkVHoLQJrdaOxyy
eINHsLyQJSDKuyJXAB5nbF8X/DjOJdjROscF3ajHnvC9cukH5dDPwI89VhxSkeqb
lpwYT5VDBmm08DIU0R/oDNjX3Rn+Q0LB5X+OAiQNFOcimSn0tVk6dmVuTf93W67d
nUgMHNnfYrzhYZJdRROezhEEAGWlj//bY0svds5U900diPtKNKMvhqgxMmYxP333
8idRzWXqSWnKWbyf43+KhMEccfzsfq4NjO0BhTbLa0TMBr0k8ggsswLCQ1u6H+LE
uhwDWeNAFJ1Ofv/6q4V30LpyZ8eOuGAflgHfDnDSJs8u+rDnb6mEKBYk0pPlRS8Y
WHvv/k1P2Kvlf1FotcGNqhay3CxKRKlh8GR1UmYuEjDCrP/niWVv5+d7PNA+fX4a
MurTLlK+2T1PsOtJ7zQ8yMOyfKAQErf8kQMxvjUpYJyuTeA77GxQAxN/ix+uIcwW
YxuZ0kM52RVkjMnIMqFI9cRVdJ03g657IaXzbFKPq+jbuvLJPU+D1NY2FcNY3nJR
0TUKeW3aOUJ+FsX1MC2cNK6WYRmRxI2cQXdlojCxC9bH5jC1kZAMsT4GkHGKJvrE
3Ey3s0BksXkCFkCX0OliX1VpkN8tcSgpzpoBtcvYJ5SZZizxfJKvaZYUF7EsXq6J
6lmIr7RMMUS74ib/Idabd+Ck2LAf2XzhPfQdH6xmIZE4MEEpE6iEP1hwGTgvvg9n
yhzJeeAnZxt1pZDXVFfHIB/6UkhbIPwKl1kioxm3GPYb9KkQ0gvHGvK1zBodpDdu
HsFKI1p/INav/zMeVRt7SJ6thIAMVCqZt/7M6dXUDNRbaCM1efU0PYIVeYQKUZvJ
8ZDQzJxVU89guNG5YKip1RSPjnQAlajoGw/FbMFlsoKIspmV93iYXfzoKjD/XoHz
JqdExYnsybK+9ejX2JiyD+M0AA77ogocnyucOXkzNUhNgB9VKR34IVdihO4zChix
AmyluCslpTq7CGkyk05xwqe9Pb5rvLCGYXdrk5tXNOqJVy4Eq3ieALyAvYUJm6iN
pTAg6t26Lef0EyAb+cIulIlTffY/fhD5udE3GvxfymSaYzXHNijgcvhuepX0UYwW
lVtUBbyIEwiSgMskozLJMG5L/70cRtunBYXZVYKVOtTtn5n/wTbHr+UZLkZMV/hx
3YE3VQNeBAlr53Cqm5jRdJ1njDYxjCPslYdMivaW5mSRKJPio5GeA4CqL6hwluD2
7uTh9U+e5d3uyFsHJ1CXk5pUI1Hf3Dku+M6vbJjj1BZ69SBGojdRGbqUTam7jEhH
ZudtJhwMpWqWoAeQN8RRM1EvNUPL5hqVTMJ6kc4GC5OV90OhwtNta3dqKapm1kY5
41JNds/jPC5q50FC//qxykzTqU5LpCwJe1BAwNZoj8JQ3Kc8O5qAZlT5FEf8yxE2
j8fgCgHGkTyGVaPo0frMObTC0XqRKj8Tp1q5eMFiewbOU2RfWUtkxjISnrMqpFIV
8+Waw0CdMx3a9/siAU90/Do4WdYcugPVd8EnYc475vMrz4l1pxxngTYomlkIOdlM
qgqj4CNG1T5g1NdeA3fxhg7gFcDjFFtlqpH3QKw3xoyIpUtX5W8+yLfC815rK3pB
AyKLWch5KaFv4VFNXtAeWPFrEVV+Q/w3JoAbE7P5a4dRc5yCDrjdkhoM3dyzbZW/
wmoauXe2NBVg4t4QfcKQGtM+tTAfM8tSkdO1RZyHPdNgHZshK1A59OGz9O6SZdZ6
lxcVzRv+gbdlIMcEt6YbDOu23ALnL4tp4rzTOwgiVfCc8Pi9VyBs7f49ILXLgRFl
xZQ2PTrJ28rAMXMPiapPQ6V+KdWgqsLYxOuDToiKvAl9pFPsUmgZu3mLXabbNxDc
NjfBlJNbFHCyzBeq8miARDhXf7VvJuZww63+ysJuAv5/NPJR2SN6OPE8se1mWpR7
o1hO2TvaKItNbgi4nkmUEU8NAJ7QbMhDw5gwFCI1nF8LbsColxx8sEOUU7AUntuH
YCygHLUZEpQWm8u342Q2C0EOylWFRI7e0nGKnjxbkokHu8UFYlc7MwwnKSL0VVd3
HXMqd0SAtmVA6Hs5aqnIWDWT4I40ZaSBAYkxeQat8xeihiS7B55C2gJ0AGNCMHsX
TUPt1GL+MkRZzKYpMzOc6Ub5wkfrYbxHEyp4mpKdMTiigVM5oZAh8ejJA3Kfmc1q
QI0sEvUwASBTwUYnBTNBYzwHNoxzZlqHkq5SAZbi/h5iUlxz1DBzvraq3aQamz6W
rH5JMzKESHG2h9nPXN1BeNXm2YJfBZ2Kgd8Dl7LAwfG/egvWH9vD+nRPsEkk1N7S
TdLXnffpsgT6pxZFWhwHYLhAWHNiDMtytuFUXcCCW81i6EBfDCugbSoeTzKJeu8H
8tKgr4yQKEAfboMdWcXjQmEo7z6K6JD5NcSfl/sYeqrcCd01iEk84/fBtr/y+LqU
NwiXocSaGuwsTfohZqIWdtbsrbR+4DaBBvILL8DBWyDyjPeqq+rvrIx4bv/hJXb0
7wjYFUYkuxMLd33P6CUCbxbZnIzx4qJok4h5LvtKvgPaPKakgH2pYm80j3ZrSVfg
eyQHrRTOq++NT5b33Xu7IQ==
`pragma protect end_protected
