// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HSK43RX6mMwKdpp1Ut7y8qxenNeo16Fwlr+W7Pn4h6zLD38BPkkzV69CcAxdsHCe
17XKxh8Vo7Imi1q8XKZJ6+NHUCheuGUQ80i+07Vc2TVWwN34nxRN1YqllIDwRMQ4
HEcx0odYNWv/HntV2fqfgaAbEmybtTVY4cnaSj/w+rc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7776)
2YIOr6ZrMqcFIUjY2CJzDtLD9xX7lH+DcBoOXOiP+Jcpx4IzJRgYxAMOfG6N/Smz
fPOjepFgpzaMDgttYq7YvyynORMU8KTh6+frrz+Iqg+/mZ0mvBFPTTUbg5ncL+Ec
iRdikl/fmkXJXUdkotsxwTfThP+fJM8PBnhm8hRQEGtx/3fD8QiKTSUedGaLBuZ1
TU7/lNJ49nkq/5jCRSS2+7OEsgJb+Y8rOAdtxmLi75TBtjgwkCcpX1phto4bukU8
WB1iFQDanx1tQT2KPQkmW/Gm+2ZPNfzIVbnMu5wXp8/pcbYO6eeapRnNl//0wz4U
1ycjwTo38d80QcAru7DLSB7zQ7Tg71bX5vNoFAEALsM9Bb9ug47YNtj6sRFZ6UEY
RddOiiWsOxpO7H4641QVi5iZOqwZG+tlx1SlHGmMefwNx1jO0JKtZLp/8KiixVcJ
kvhrirwlGPA5YvMEfwMMjx7jubYXn1vIMkQgwf36elqenkfy41TDZQ2efcHhxA4U
xBmkXu1tYXLbfaT1iyNx6eaPdUl6TnVtAWqgm/4o4516khJg4h8vTS9OgHT9zQBK
8f9dSv7uqwn+NG2Ab/dAoA5cJgPRXVYHsrW3okpZgaMFiyki3xVU45f2xodpc+QM
+hnOCTNANznZKIaRjJladWJRjEh9RfyZpV5GAZZx1CZrapYJ9fTch4a02WWVM0VI
iRJ87hNuytFd1gLsE5pq7qtWRZsrISQfAtZCDq1zDqwSIIWPc9x123Ycr5kReYSt
wtamyghwk3tKWr+4ga9jV6Z/n4CFHjr1IQJ8U8xDn/v8tSO0rBToSXiwFFr6kX4I
+KiJzNTM1suXuPgrEJR4RBRXDn53yt0k1hxBW1LrRJGUt9wAw6+VcozQdiSB8FF1
HBcO7zHABRIZ0DOFYMLEWGhnnoJfy3A5CRIRtcpf5B84zXuVxagRuSpDlhw2yzVi
ILLD4iu5vTUSf2Jrk2Mh1lIlz6GozX9wmQESGXMe5hUthsLof2b+UfvGoSfoEbZG
Z1f6QVD8TGwAyLGW+rryrId2QVqvX+WdDlhorYMjK/alnOYPaxikjuZLcqNoifeS
fKGR7qIb3CD4P67EXRSxqxXVd33fXBndY+V++A6+8YLWrC7X1TCtldouuy8dwPR7
UUr6iGzMtxnafaCa3u6Z0ne9rmDo/PvAMW40L2gR/gdgqHuBfF/tofR2hOZ6PU/b
01L/5EJe/DjMeXjqJKsfRK+SjnEG7/HaUAYDwqzsN25ZJlYbTdGYaiZA29WFAi7o
6i54o7vASmMPBqC2eXl6xGAC3SMLPUa5CmF7KyiGATAaPM4Hv2FwJSXsoQ7lEyNp
WlrTto+LKypI/VmpiSsrrofpFppVa86nyQjHhM3dDPqr73aHZx8ImEG46keTW//h
zXQNTB1JZr4Q4oVIyc3HE2TOat87988ML9qJcOcOZAWKCANpXYXX1D8iZg1OsX2I
3mXcwQcAxur5mr/szEWXcXzLjktsHfbJFVNCRBzhfZ9FvHWXD+vVeJ98C0gOn6ZX
hWEvdQZiTKhyEL1dGlL55RDYocV6xBisQDYVC/0SKqzNGDPLkAH+6NXAMrmui0xH
LL8h41A9qhW1ciDm9lmPezaNebX1roDQwy121OvP/5I8leeiSyanl201zBDaabWU
CicZGUSokfwmpLfDpVPnhwKm1o+OoWbei471kf+c9L/YjfxXqqiSN3mkE1YFfRs2
TNrGyFX9W+ZPr7Z2uAR3LqCjiNtpSeIsorK/GeIdDnuaospHzquMtuo7A9WdpWAR
GZRVfLZzBsuQth+SRVNXqxcQk0VHCKIiOgT7yIv1IkAaIpmaTs4WB/uX8vINWCMT
/oLpdP+0afKPKCp9TPLf9j06bO0IAYhj9td7zRUsCTHGtIr8xVp79UR1zciR+gBr
ETCMdbe968sF487+Kc/H0KZItCaCNhVIyWkADufdFEmpqQe36BcEOtuyDdmiIbQ/
zaCKQibqFKu/VYy7scRcFhRcncgM6dT4+FyoTR5yMsCsKDQDgccwsT50IFTi92lq
HnpjJtPmh5lJNKrhNRrhELBfkqM3fMvtOrxB0+gUSg1/vhmevCngbt0Agt107QAo
ySVoMxx5oMMLJiTVoOAjz3MqN2aj36nC/KroOkBvY4Q0crA27pRL5FvIJcImKuV8
EZReffxAF6G6Yj2BR/O6Rs3EWQFEfA7eGeHOJZOk1COVOCv5/7uweVtVRDISYcSM
zhsVbPjxDYmAk13D6tj1vJ8u39VNrMsYHIsV8EhkhNTprSbXxvmqbSafj0cmX3OM
BFwpBS5xDtSIAD1aG8EDV8pEMte/qBYeNMlEOdGuvkGv4is2ZTs3PktbVvE6mRKL
U22u1Yx7Yaw4C4UqvuwrxKKQQcW/6iB5tLA3LKsLO+t2M1GeiVJ5dEoQSXO+7NxC
D/Y6cckHdyaJcBWgSEbCtgidWKxav4Fol2vvMOa2xgN8lStLtZAswtqGc1WT1pqP
/MEULr01MDwHVMu8cIvOQj7F15cpdinV5IrR0fJNtwKmJCf9nWvhgZhvY5+xrDzC
6Vd5smaUpX/UQwKaGVFEI6onsozmlseRlc5BXFVSacqfojh1lf3Ln7UFWaKdWbdt
YiFKvQjQ5AFuF/c7z434j++yegF+gPDV2jUTmmGWyBi/o9AW728NCJYE8YZO9khV
7qitQrfU33GAQcWEQc7FxseSMpIDcQaSMdUxdGQxhsuYIfNf7SGjLfa/J8DkiVsk
0EnsryaoxvEex/eEEJOI/qFjAaOC4RMSAAbFrjo28tClVRP/vPk2PrUna5idPHRT
r/8ze9C9DXVpqR1KdOy2ZCaOeCqSn9jSRPRTEqnXMGkFsU6LOQV/bv26mZ9BNoPc
xCmaeZo0hv7pmLeFbB0JvrqKaaXHgyknuuMbtdXI3cdrSpMM8dOXWjhWvkJ+rqN6
Nf+hY0ZJeCmRBoG6jRTZ05BjSz15p+ZKU5NfBTURlu4C9a/y332MbwzlDz+fmsqN
+ydpChbi2G/HhP+kx+AD7xyRQNI1ezcm/+xbF8ktnt3vN0u5klrtoEqbU1D0m+gZ
YnReeElSRmQrk/4D7fBMa6cA3S256p1IAJo+isb+ZBHrniL0DMLB/NIrmwptOdVC
lwK5XaiADC1RNC7NTf64SG6vPRJKKdBuPCakHlfLaYOq80KsuYbCDBWkPCYHehx3
7KXRkQBUqG1e/SD2YaWAeMuI1Q+UZZ7lv/osI4QV0WaSqL+QLd32xrtuxUc1Mc6P
/pgd2Tdh3KpYjud9nNgscaMk5r7x2JNl2qNik0kDpcYTj/fv8hZaqD+BT/6S9vls
1p90uIzMFi9/EyQ6YIkkSGFYS50g+Y+POI+0AgpntHhuahS5KIMGSxgjsHbiX5zW
65XlkEIUOFk2PmmMUCMEFbmYcOrGFjSypqq3FXqJ1AQt29YSuvN6zdxs9RblSING
3aXLCcFBwA60EyMBAp6tty5Jqljjipgv3MPXa75a9w2N7zdnFW9a6LJZJ42/oqdg
Yj52LZJQd3IJHgD2CFD2lD5v/sZ2bbrD2TTu5LR94sCamso0xz0bXFg7ENmzwB9b
DiyEpGcUCKQ17yK+pdEt6PL2BKvYTkwgUnh+5qbg2n1e7lEF8ju/Y6mbqBpP19fD
n5rrisr7sfgCmcwlVAEhU958nngk3D+j5cjMYC7tol6dSc5BYBGiwqFUVadEAufE
3r/6/1E7MIoiOBSimnA6A/tOp7svuNcTxAAYlFmBG/hYhOINiDUQhhON7wTDtrBD
vfuszPm4yRUcbVZL67VPxgumJRAKiOILVLpICf3hyZKXMglap1tWszwHAroNZ4sk
uSWHw3b+kLrw+2cPOr5bIeUaoOsZ8OQRDmdk1oFjWRC+1xcCASCjAnpzUy2DKfRP
/qotJzHxedmfyIWvJMhkSecZBDO9/WIRqPjCBqKGn/JIaDZ6ZqPh9liEs7w2550f
hTxFzyBNvBX4C+OCIWE4srYlW758eKbeU/4KPsTwtDs7Y7AP8wYAHZPEZZ2wcPH2
Z7S2yccFIULPgEyV4MEiQFsZYsFV2evvNU12oh2uphSb6Nk1QjYiqhbOihs0oJiU
sunoDVYW8TVJWYtUx795q2Jw/UNo+G5NJISE4P4811QrLobPurL4A+SMZ0LggszN
2y97Y3cj6beypQhPa/2mR+31dGcA0VOFiZ4ByobarmXVqehj0BhO/q0C+f5h5l/o
OC+r9nQmIX5G64fcUzwdMYqg9ib2gShljBEcKhtH3T1CRssVkNY9OF/SeDmOFlW1
xSk2+aHVD87LFir0H8oaKUfqsh5a1ID3ucP0zJNU0SiZOggOpm6yp+ayJdu00ABf
jNeFluySA9ytV00ZiDiYBbOi1WXWzBmPC1YaowbCEjA4AXso4DqODngE7w+BmEeL
lnIPNDaXkY5mwRbzWu+C3cjfIFgTu1JBopOeMc5KFXDY+0xk+h9vWbftLkrKzic5
mjvC0DBVLk2Nsuyz1UDZwB/i+oofGMOl/9yO1gqrG1Z9mPHIaF7ZBsXNVvdmthAV
mYzRCbpwbBC4uIBUkZGzvXRLHIk5A4iazSBiXpdm3wB6X3H0v4ianvS4tHVomQg2
Icl5q/WnDyhXfc8lSEL8WsZe6CYM8/4B/gFxRrPeilMw4/xaHexoObWHnOGpkqeo
Wv3a42t3frLzmYJ9o5Q0auB2cYvDACXgCYD8EYCRjt4u+G5vxNoNZxquCsDcLN+T
JhB3vv4FZpW56fFtn/4BvwjD/muvymfhyxzQzN+qDaSeyGspCmqdMobDo0AdZ1X6
w29wvZoKQXVg/DKSw5v6qedEcXMzJ13Yb9JJKYmLIxNE+iF3OGOCQhsF2+U3DjRF
t9L9dURM0s5hXB25e6b4FhpiOIRYRXfVyLpb4ZxQHktkGapJeOy3Qt7M39Aipz2w
hbOmibje+ctRZmsKBmNd71JqFfE/t+HbIUQHtt4MDklKWToU5PAm+kWYEp+gmkQW
rFrTRPxJZHfT9ljOurjDY2ENTE2RFd16yVysj1osgQyGHgOmDss/nsg3/8/CI1wg
/rNEoInsm4d46G31SZPO8mVg3EZ7oB5rVzVmWgmEuFdVtn6mf8X7EW9UOUHNhKHd
sqzQyNYz6SrrIEdEQn28Vwkb/6r/OyJ4JbuCAWr6ElU5HomGffW/z8mYnCaqEhRv
poRPjQXjQqdpmXkNzeiNOf4QdF83aJEaXhEhADHURY/EfWzs4P65cy7IOssgvntu
/K30hco0HmwJhigvBO9nJgRjt2Y7jyltFvJrQup3pkwrwAFTJYuHWqLPhKxwij0w
xzRXeA0FX70A45LDwajbjeR02RIVAzca6EclOz6MgzZ8E4mHHZKUSvedpqptbbtk
83AGfGe/31uuF8bcbGSJh8p13/7cohnJwjFPzcn0rxokv+WwV0LPdPpkRKUxDNia
5VQJ4flsK2D6NxuiBwcKi1kG+fETpQMozxJZa9rQnlQDJnSB2rPRcBthEpC8AALa
+6IPDD3Ehl1+H3vkus1yY6Ni+XXBefCJ6OeSl5X3wuE3DO4/AokoSN/rGFQXIdiF
FZd7urBdkAG7hJyCyNZ0b8mLda6oC9kKYSLfpEHcvp0VAyMd7SqB+fd2f/Qk9vFg
mvgHahav5g4Ina1Aglr9nunJQNneZz1aqouIx3wI0wQGx+mdVJkpD19LXb8fpIPy
FQfO7/E1TzcmPrjTNnLskXlgWjfbCXKz9AzCnLY1RW52LflO6at6AKKnv7NmwFYe
XTZozX9/RttDwjjoPtighBNQDrsw38n41I2X8Q1+Jgn5Snk5XQxBxWbfOE45f5r/
fou/wIwNPQYh7TokEhVA7WdXDFK+YiQ1t37/ZhJkNJKW8l6uQYfW3ywudZF7v+Hq
rE0WPT2wgorX0nsZ2X0mB43oPpIUd4ed3Ju02V6TpLh7x3e+0aAUuWXLQFX1gEJr
3D9GIsg5vhZvh//PnDbMmt54vHHb/kvsQ7EPjIc4DgzALW6MRyuIR+zgRBCR3LeM
RSIrnnQUJRIiTPHSMUSs5fTC4sAEHRwmspXW4aY6/zxOdT1BOSdy35I5B9Z6WntK
tM8VZJcV4HSgnoZ1QqgJMTWE0yZugPvUEvlhzOrUoJx69t3EYnGBCS89SP4RvH+q
ex/CH5M/9hekMhGmDuKKo7rpFC4bRQHHWUn8/tRxFQsW/UDiOMM6VaJHbls/jHoj
Ra1KCiTXCg0jpnRsngp8X9qfzYcWiGe7pwbg1RpACwGh7yb8aEuqutzm9kOzA9a2
b4UZQVwlJiPHsa9A4aetRDuAt9yjeJ+zdCLOtXgB5noGyqhc00ZbOMRv331r4Dqr
NuUEPSDxOhq034VgmVVauQR4UhiWXWWPUm11WLgZ1MjhL7IXRZZPtln8ESn7gAwX
6iIvM7k9MsXyxVt8aXBQ2TCO+EyxcTX1EoNKWUnJYHIv3i71ek56Ao9mnjsimGBt
vDoD1dAJNnCkEVPJrOaI2CJpuj+UNW36wvglTQr7udzp0rZPX/nF8QRB9XE+KfOi
DnNyjgnQClP0i6NXUIxRaq59JG9ew2bwrhQlr3ivZV4gDrpFvS1c+Rzx3wgfYViN
hz/PKdzarSWHdFFh8EFDgjBdzQqKcIzd0sJo5oCP4zJp7TnjaEwJjN1Xl5+XqieP
Uoc2ieq5oaJ5nbId00PbgAYShkbN2MYFrA+PFoQ8ON3VPhgMqZRp5KEim1UxtAhA
QU/Hkw0Xya9ZbNKg2c0aZvNou02/YmUjHnOP2WZmQufO6uRetA95wMFikaUhhCfl
lgnxGQhFwsb+6aVv3jVxxeiLSRTVTemv3OwDcEg9eOhjev/4NtMd8s5NJWpV0rOb
lWM008KE7NWEW0qT9JKaZzXDNZJcfadPP07w3RXRezfi3lWEEwlgNiPY0aIbuaZf
hHAZYKNUPs1ub7K83ycjJPZJFi5vNA8EPFstjeGqRGHdYlR6jvAAc6kKq/kNpSRK
ra+tcjFeNMjcla1yLcH5WnhKx/oym0NPqjRcCuSWylQcWthvZIhlwF7CDQpffxYD
gMoNQF6HnZOS+97GYcPqDldasr2RX4HFLvafR9cqSesI5PyyQ+NUVYA8YCb/VrkN
HfhB2QPm6UsWem/I9AbIoTVhysytKSwg217+Tq2SklSsP7SRdC+ZLdt2SlRUOLTB
bV7jBa0ZzrRSxWLXdZyjev940N4zG02PGZMPJw2N6C3rnPtX+3O8P3oeFnNkfYRX
Uhfi6YxJHzhBT0zkh/6rUnhpnNa5JTCj4HJJo31rwgqQVtl8614IxXUMzQ1DG5Lv
NLq5VXfZDDrwDvpOiZ68Z5O1sJOQvG/jdTD93Qybb17eqyaBEoy2JdS9qdyM4EVr
YnV8A/hoFqgbZIN8NT1h5sQQb57iM6hwIDS4lUsJAgGVJ2CJb7yyWdD7AjIk8DMc
E8THL0TwjqXHv8Fx/sH4cLbn1/4qgGAR0VePzZFX+JA9DKPx7ubViiTKQiurpz4v
sQEKD6trY8iyMwIAlYkWC9DR/VqOKr3n8peDpyfAB+tUp/piWngAaiyy4e8jhUrI
38RkfbP19adsqMtTMIPZ9CWsu8BHAhZbpXPCdBBLmw2kMRrslFCC9jjR1wBwqqUc
LWWyHBF2//W3dfry9o1iFQPga9BC9F+BRtKM9zacsxlTIGIO835AMhlVWAJBtAap
HzdiyX93e6bVIpMCxEhDXENiI5rEqEVP/i2F1VvI/wJcTZo3/UaK3tZ74+2ngLVz
nekaG4jfk5ZQI4TGWjfx8oVfT8MjFN4wGRycb5ZR70i7cKoA7iZ1xr9Zyhv2QAQJ
Wuhqj7l59latqMgRKKCpxWO31Hu/otiVrJdt/6ofcAIqLY9QEJozkDJdBoaBboZF
u9iyD9bM1VfnQfhJsJmuKMX6POTYLz9nFeI3LCt0XMaSiTLuChkXlNcL4hPM5jQI
TI3RYtwSc6z2tyjO617LCbsOkUINcXzjMvYOBvz/dQinlsZVR4Mn47ZrzcgFKx9v
dr2RkWKzn3UumITS1kYlrIQUm4ZGFzstXYdiu/sNO0qm/Nc651G4mrndLYDz7emY
6t/Kb93BBn9P38Kgt7933tzy9dFSuhxE5xmeHsKxx+JwrvuLtDCIe264viH0V7UZ
SD8DfovK3VtXpN7GkU43RoB/IUOKe+iESWc32oyfhVUVRfMH7cskd35W+NIU3sSt
2A01oj2PmyGSvk/ACqs02wU1OXrjU/wVNn28OpBUfjHUWcYkIwS5ru3UvvqFlfF7
gAEbn10U5QWFtu/eNIR2g1aAwCpiUeoJv8dz6RVDPehEcE8RgMIv1d06lKmrOa+2
4awF3iAeNkFKcUy58uT+0o6g5htdmK5wEX4bpCn2iuQdfVA13F05qW+5L4PDwhGp
5xokG3nPKNvRxWSoUbK8ZUD1iowoMBAQ7AQU+13DW2+KC4OuHZ5PDWVIn9PvIIf9
foIfRwOlPhHiTFb+6x1cxYKG18J9bZ+zncCLmJsq0SG5+1qjhHHisrdJoVwFPlJG
K3X1FRXGjXZUZhtYODTR3DDfTJ701RXD3fg6X+En4QW6h6UueGG4i0HiQnJudyQ9
BamrvHLUY55Y28wON8fhimSKJzImaQ9VPLGqjWjraR3ig/TXLq4Vd3JK+lAwaSLt
4SfZydt9l8etW9NVtTHcPnmzhXu4JHZcWFKcD1MCg/Ea1jh6HAlBrdmh9EvvhPRo
gxNUdaXeriEBmgcJCdJk7+LwjfRO0huM9ucD5VzZFn4+7UI4+b6auJ3S2KX2LO52
iI8ZUazLNV/dBnwvgPBKNC4ZJgdlm/uJ8gLaUKutUV7chvpWqYfD3kQs8mbkgrA8
QnIyg9tlFL2sGHOq2+w0AsjRe+lSV8DkoGcQJtncN7gT8xIQTc6LILAH2ji0qayH
Soxzpo2UFelgnvqyLBs0B0ASCESVQIpMwFepWSeQ2ppsYlQAWqheoIsEqcXgfsp+
ShVxvVr0DG84/R935Vf+sFrHXwHM28C2AVnzWKHHfpdQTrX2ow917HloxFbGGQWF
LszhAOH5kHsC5BTD9fA5w/0rb8GAIGE38EQwP2vHByNzN4wWcuwH45yTLV4yqRsQ
gQJZwunBTfY8EtOGY3nV8NuNODdlGOkCFyg2L4h6WaMy3CPI/A8psmi4BsCC5cLE
YVthhbK9QnL586VV8/S6s7f8UCQk5J/e1gxU7017SOTvFQ3VS08032bR4GFpOHA8
g4s0kBuX7yeA+WhibEA+3uS5BYn1UJ8xWXYYxtXffKHx1AmUhGVYNaLCUwumFvSv
/VCSCLRnyZLNQNe8Qa+mgTpUM4Qn7zCU1uvOu4JDFIdSWc1w+O95DpmAIgTxZFtE
X87Y3BnK88NApU2H/NdcGo0wxBVw4HQm4Dvgi7bvuyf0hfhJseiUHRyQeXPQQ/j3
9v1qM0+sdKRop8aYAwm+2U+6gpCbGNlGbFu/Gm6y0SLYsywwaZ7VuXqy293h/+aP
Z4CJvv8c2b0lhAzr53/eS0KX0sGVSqswVtkySQGT7OzDx61BgYJUVvLPpw7+B/Yc
1xiss0AcuWZfjmyL0YFu8B7TMekpaVSIxRkgRgiyMZ+LZmQ1cgUJZtjLKGuehCQ5
3RqOL7zFel5xN/as5B/jDjxRFvIlrcfKbnsaYNvY5uo8xokYzcAkPoFXkvn+myBY
UAlHLqHB6lrRARYM1lItbpt5dsTEG3ZfukEuqOqQufFOAxtD/UlC8MFdNnK1G5af
Y4AUfurSXd9Yhh2JJRsQy3S+HasNKDfowRbIfxpWABgJKandp8DoCFIl/oECK7o2
KVJeN/zFbc4c87OzCSvuqqh3zk/ZclhCHVwniY80ZU/XdCBNXvxg5rsVl68xmk/7
cj9FFI5I+TLVQW2We0LwUSyLqW6rEXaYJo3LnKAYhlKs1WZiMB4MRLjIYIJ7MgQ8
OHxyVigm4q/DR1d4f94w4oa1QWWkQWji8CbLN88aUalhVMY3FNDHsbG4mX0XTSSy
SCOmpae82FoJknwe3q/JetYn2Qg7yieqJ0VuCE70urI7V2c1jA2p3PWSSpoNG6kF
Zu09GxPdslf97X7403obsGL1Tf7AsosceYQV5uWVIsFBb/QerQLhRlfxi5qqvCj1
3Z5/U/HFz0c/4mBlnWUYxLfq1Da9a91m2VpVbw9sRtxPhOv+5KuZo3FtQlwORlKO
PdaVLQNy+RUGh5PoYhS5AkQZpqOdLtYx/plhGnRwApCn6yJsjX7P91wE0YKki53e
W4LVdDTIBJaL/lcShzxlmHm1wqSB46SBJuzerbXrTnMbJ1g4GDdKkCEbPvNxQD1M
tEKYu6nPBwoX9Jj86iwCbLNT8Yn9T86tUZ3HtZhfiXfip5D3Cou3HjuMxQuxcdWn
`pragma protect end_protected
