// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IPyihrYhGOF9Hl+4YV7k6+Wk+CXukl+bWaQKaBZLdzBm05grbd00jhpRc2XCyI+D
Ttyaffpg8BG5vCBQ2LHCHGuZFocyMcfW/w4wTJW+rafugliCBalQmD31qkQJlBPr
koR5XHNO+sOWVU/tXg/Wmm9Yh778XgZIH2wkI4YoXBQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9808)
OA0kq0ja+THMKa6aKyF2q/p4qupi72KLyMmLGDUlxID2k+xQPMGGtzIqa+mEWlRD
fRQy7295ZFuc/XWsMURmVdQrGOAPSU8kEVL/t8oJfWJPMh8KtARmJvTGjxJQ/3Vu
u6tuwtPHp5f2lTLFjClsvtsHSWfuSiMlIfiSSRfl/1/rNFcUwqyX7IQ0gPr8sX3e
bYWQpf6Jb6Du2BF67uTvl2opiDwzZ7Hho67qSmK1XLMVkrleowB9bsNnHmlHdNcn
G2OgM928mpOOpd5m475Lq4iXMeyhcH1txBOZheGOplcuctzG99HXd1aiZ75IuOQH
OZ/xbir5eAIc1LUWMrisnuo5I85ImJJFK8n+oX2uFj8MzRb6FaxgMmBEHCkZWWYX
V6jN72X9eFD1CL2pZOmJaFAnEicr3gJjbY6vxmyZmHVSB9jzyir5ibdr0nI3LHSi
Ye1stdM6hzSrSLOqjipMLwL7Ur8U10FSI4/uJGNPyrNUzxocbFv3No9RfudlGIkG
dQzWtuCvQXUtGHVqjqQbQV7lTwlE+TbfXGaQ5rMqbsf5v3YRzTUXNYJ3mUTkC+lT
gVI19WhNwdlt63V8x1IvW8hKPH0XRPp0sumg8i680CJ1YIjmpGHX9j+iuSdh9wpO
fRMwUmRCR+3+kdpPFEgFWNSVON9vyy4GB6d6HQ72+4EikUzbimCn3i3SPRaAUqBe
/fIvofsuCx4O8ymW1cuwOUKsdErjAPXcGTPqkflTNfl2RTozivmuek5D8kDbCxs4
9VpdKLwtit+z+mfCPVgUtWJXeuZ1CD/cWalA3yfmiK5kUlMNfvvJwM8j9tU8/wlK
EAf3dlw6B9PW2e1pmwq6PNaQuNWke2sjJ2gtYk2bRnyA7XXwYe0eAk1zANqlB5t/
leMYq+t8VWiVgkpGkArP/kRu0lhYayiZ/fIzlFuKnG3sihpuNQw5fu3nyI73Ye1c
ZLwgv/vyACIPWM2g+emOd2Ra/+voati5UaBIlaRn+zekoEpKvWGrxn6Lh7D/dHBD
JOK7HYsdAVhMRrptIPAhl/wgaqv0Th2Ahc8EuPE4TivRItXFB58sErsNLHhTIhjs
vodFkL7i/NwENi0NEkcSorE6q4d257B4KgW+881x5bErh9u3d2pbYbKbl9K9mqsc
e4nsvdMNmPMu+kq3WcSd38tBDK4WDknv9g0kaK1aESM9cP3QO7iwlozdMPfTuDlc
YlfvuhhQposybkRPNNSbnw/clM+nfM+SaMF5sWTim4JLkXPwl7gMNA3iek+DDCkm
LeZNH+DD5DKH9WX3OH1d8az5MiFbCkBSZuvu8QcU5Z+ZFAhbIvsLR1jhE3hGVh0D
zaZ9D7oqpT2d8TClVIMRTpw6W4zHGtIqcrams/KymRD1bykG6aqaAUDuesYJKacd
vXUB0vPS/Dy5PQxOzG0ivuCziv/c5Mx3Q3wTKbVY639MDo1wRw/6bikoeSXGYKqT
lRVHw4t3xRqyi4DlySX3CIx+ExAsWVUy2nsQcmB8aBpjm88RkQkOOFaR3H7L3tU4
HuCWt0u83O7TyYRZCGk5JNZKrtNysfgvPpQr+VGOxSk2JeNYpko6XtAysC7Kzqb7
0cw5YdAdMVJaYE6FnkNrggbYTnANCj+sZtNpOYa9GaZBDtJv/I8OVS1qsaLG4tqJ
pkBXrrHOjLmkrMZfQTEhtHBO2+/G6KDK1+t+bYB2Iip+OrPUf3iTlCcZgowR4eis
3Us0XMFhuKCaKaj4Y0cfxZRyCkMilpPVBzbbg61NhBRuqop2NmgYf4TlOVNU1VSL
RO6im8aa/aZ2QB71tF/M002wHMQpfDf6g6A/2GN3nUJ/6g0Iu4/xHeHFXAXbAgi9
EbPHfRKBEm2iYGccIwRu0OXjUfNiV+7vIdCGIx3LfbA+utYqgWu5W3ZWQkcSMoLy
SGv2LHPp4bK4mJ4YCSne9HautRNqMGJBePzVLwKeaBYJoXB1aITDLvA4xN6w6rM5
Ybbk0KsH5zS10jQ3vkev30RQUjjXao2lGGzOfx4zvaEHMUVlAwuON9rgO60uJOP5
9BLiEgkZNys4aJukmFLs94vlxP6ZGMAqe4J8Ay17AZ66ksL0UDEjBTeaxnLKU7d7
6V9MK4pPBWnJzHRU3zYdWGpHnYne3mF53nZFQZvm9c1llPRKHyQWUdpFhmo5s5Sa
/SE93ioCl+NYT2DB7Uuu0I82/jn0oRhXFDV1bYzl416oQDtVK8EO/nld+KQPkHpZ
AsyKg5sh63dvUgFcYfG2XVKxVJXp/QfJ/mMdbHOjdX9iP1edrJCWAEDsI4OTjjtw
byn85OzCloCpg4q+uOPWXhcOeVTy9eLD0YcLH3cR36WNtiKvqCD2u46Zik1L8E42
PeX8Prho8GFIQBLNjxPfwos9ALxuqG28zgOvOdrNvjUR+CeSuEdO0qL6WXqSNuv9
7yFT/yd96dbFIu4MpPESE5IQMo5n7434TRhO71x/jpbyx7L0OFWROXj90e9NNgTg
587fQPH/h4c8SDROCtSqEJ6NNjDR7+HxurfaMpF+sjwcB8KK33Qd4p+CeGo15+6P
WrzxeJNp1/u2hE9IK5XoEcyHWW7N2EPRFCJgD+uWC3bd5CMAS+wUWHJJ7uVr4tQm
hf6FkReCdtcG+idNOYzBqjRrEg+SeoZfZjLPU5mfFxy+sOKS+V/eP4974lHq6xgs
zHf9duTn9dEX7GZ2guGqh1hQy9VVvDcGKLop8v3Vat0rqzC+pwieLGSEYe4j8fL1
2sRkE0pejQRANAcLeUFZ0KPt3BR/2xf8kbtNoYMDvNr0THklrh3D/1zPEWeo+iSH
ylMvsCaloVJWyxMKlyGBRgbzUGU4ScC4/buAOLfrCSwBwzWM0SBU6/CrdjFrdPja
gfLaaLm+5HvL7o4ubR9JWSdfTGLykC2vjCPfGGzcm923EvLCZcI2M72eMp5kqSFs
NYyILet88emgfuzbXRUn+bSDA6VoG1f05JkWgPYGSydYxQAsi/8Wpc57Zz8w2YK3
0CorwF0BQAPVWo4osrp0iK8PhmUCVSWLHefvD9BdB4mS9Y7+C3jS7i3oBTDiw3YI
LuhWR4PpbXlr9grfZGRy6aGZEbgCxQPtlLgTPFBYMOxqcKWb7yV+EfxtB1ICOMxf
dccOhGjIFEN3Z1fTKWR70QnVApLKKL2GDMY3xw7oDeVb+yOTAMiPjnZvPqLDnmzj
A/w3GWM4FUZnnE1Bw6nca9KQaBneofJaDAGyA2436PJ75E+xEP2N7dtYq+MxS5rB
K142qt3WHCtGn1nEcvRw8Y2A/r6QxGQiWVESAboHv6EunyTciDbH0GJtSYxJ0JLP
XFQbGS9R3IJv3ttEPfk2G6VZbWrirQzAS54JlEj+qcCrTBWsaGiJ6EkrCf8o2KJy
dZAUgILa/RYvvweMdzi1io0R6EjPYhDsCJbcYvL6pk+6+JGg9YzCxVFkxDbbUyJF
bXCy7oN4PInwy9lnPbIRbTD203PSSq00n3slz+Idx3QAh1YVtYCj2JA82Z2U0HmN
tftWlmkISIq8rGv7EWPXoLPpLtP3UfpEa9fpPaSzMb1AA//I/IwGEHhHAFHm+pM/
OD05lJUjrFyW1j7TMXiqOvHjKQt1UgyWboYVEWDMIA667G2is8GtelBXkJgKBcpO
halXV7TJq3jVjq0r+jdJqMLNx/10P/9EKbIk9YuCBZ32mTHJxOarySdl02aNOAkU
h0T9tctb+wLk7JW2pPcKLoNEQXsSyCvPe11P0/ia9oFJLSLfhEBzA3NmMnoqp4Gr
XhAzLYoFpD7PCjWm3xHLI8tIHeCHNTdiWer7XBZz0cKi5FuA94Fs7+AXyrVrSJvz
PwH/szkQ2X5xYYG/d8hCBpR5Hp+mVStK7Qr9/CqDZeFJfuxEmQqwv0FeZ+IytXdj
2Q9RCX2itX/i2Sl9NconQ7zTdJ0CjFiZaoIZ5kUEj6KeYtTpiSn6W8br66UPbZWM
GDFulrsL2VUaq91g6aszYrH2MrnJvl547bgKMEPgj0PGq4qTuWhDbBXK/zC+kiT1
Gb+zaOh/wWs64niYmefJexI+0hpiHk89jqWZNxd0aMCp2xZCxE12afY9A66FQ7gR
qpcbX7Ns0BJw83P67M3OPnugw2t3s5/canDXjoVZ+YA617ACA+RHWvaTLkgY0yVN
Yldd46mKuHWf+Psr6IW6hvvGEuiT/TwIfPA1R9VeNccQb/09qUXw/g9GwBiVSliU
HPsYi5zkWvwkCRZ3PaKyle6zsm+zfAcJebl0OgEFdqKvWtqUZMlDESK95h4cgFSR
ylcvlXctzP0X7CEGIyJVXaBlk9G7kUhpSd/oqEj5drsh+9dZFbKpVBuIt1jkKkta
qKmZZT6d0OxKW4f7OzS3nW2fv6Zln0oMCQX8Nq8JTuIIrkVc5l2PpTWL5+aW5Sg4
ZgeYXLONlTPXnRjPRgyXg1oquEKRjH7rYWz1R/9cpO18GrdHe5YfKfJBgqx8fTtm
qsiHOKXk7peBA5Zo+7YQ8giTUxEQOklo61U8AazR5nZvbo1I6EaXrRV/0BnLEQ8n
aTCHnYNR3iTBFSJKP04YFiSRQResdQcPTR2ccDzMJN1nfOottE8GSA4+0cgIP3ia
Rle8wklSuDRJ/zN/XahDkHvDTrBUBEMfPA9XJ9iiTvBzMWHhPqpIew5SRbjxGZpQ
N4DEIthhKoCpUm1UEICK35+GDhxGRxIjFWZ/ZRIKNxNhnYRZkV/kbZC5e8i8KlQh
q8ys1JG5SlZj95MKqtIrVdWvEN49q4n9N4y53d36uvoZqLXsshoRLYZgYUdfH4zr
hqLsFto9Bz8Mz+xPmvVSwJBT6blptc7aWQAe9/+SXkXS8UqK0SYMOy8cUUUOrxUA
nPRSN/qwokrdWEU1Ixf7umtwd8FemUgV9cB9R2CkFMcK6T869DGl3Q7nhY2/VkGj
xZscfxxlOqFKHpR3jcIMVEi3hh9TAQvsAd4+riZDgEo3eBzMy82YxbEDkVQ3YQvi
35Q08sVRkz+sWorpsi13lC4MloaD4ToAI/Qk0+LWblH/OE7x42VsW6IVaGffuqAB
6D6PEXiDxfso3AFygQJd+aAjtqUFuA3TlDSmvX/A9WTSHxmmYMZ/tfG5wNr17y6/
f5FSIbpTSyZLWT46ek2G23S6AL6R2PP6OVIvGUjzDj2BhlkyptmmFibb5sjdiR62
/NMYTYDRbpZ+yvPt1A+PFkSggWUq/ee3YtL1WnTQdaKOyIeE8seTSAwwtLIMk9op
M4sKpAysBPSoPN39DcD2JDeqlmEp2sJW+NTCQSHW6BwHmViYB3ePRSdzF7XJ/BR5
OD/zhwnxfaIbaBMS4uVzIDs0CywUz53YaUJ774GNWj88nxevRkZfQbv8Mm//SRWr
/GAA1v7GiKvbPD8lErrfmKc9qv6KeI/dKJ5FOFA8WbwkU2gewPn2HLJk3Nh3s6kA
78IV26pumSrzlN/f5INapq6cNLoyjjgpiziXo/RvZaI670ZcW1S+nAJZu7Hw4NXg
iw1YE4iA0cnc3MzfOwP5soo7Q9gKScJClf8dUPeZwiwgU0yyPxNI6Iwb1ELeLx34
WpbH1hIN2uEf1cbKFkbfGO337Tx2TavW2hQqrQrJYNuc8UeV6gIrDBSDfCAWYuB7
AhzGQhHnB0NxKRk2K6WRmntISNDBgEREHQFJftGq/Ps2YI2Ze6P1hbs0cab4Dd3n
4QCGd/wLXjYfNMCMwb27T/o7M8O9icLALlWB3pk0Bf7+zI+T4nF+A9aNayPxfg/e
gQfZ/uyg+xP0+74RCpFCfqxVnugkrax1BcYPN9mgPWwNbQjwwhE4jg89mT+RURyk
DVlNx18zCoHL/5VOxDvyk2hjWXbdOAb4NueVAjRQu13QmbPmlpZrQidg/ilReAUF
BdGuPa4fddopXgnGzoDlOc4LYmFnn5cnf36xiMTe1oTLB20ZulXvH9pEbEIIR1XG
IoooRwuw0ZQNNt1RJxmrlsiQ4zCkhQP7YFwFI0pZKGWeHkI5XNvM9fBL50Ptt5VU
SbdN2wVQsI/P5QUU3lqZrbrRjhb8H9RDzFoe4OzkMItER5tmrscfU0YRtGQXrmUC
87euhz+A5edid9f07kW0D2LFsElKEKbbMWPh3Z/BuPBxDISPD7leneMjSuOfYqD5
IWiIp9Bfz5nuekzZL+mbO5/6ESFNZqPrbCXR1ygZI3nFaiGUqSazzq6qI/drDlj0
+VFn75DIHcQuUhyOkq/wHKcLbCOXRB8399k8/WdErN481iYVn0Wg3JS3D6bSy218
31l/okaVnk37kbOYJy7kMPh++9C1bOdY/uTdsLqhJyV01Zrj3/XAq9JNeQLQYjsK
RgIFTvGyuE3uBLuuOgcFjoPy4l5+tD5HrzkFq3ntLphZApQU14P7VnqEa2ZHZ003
kc7ROapVwiL0LGYPg6C9Op/fh2FdQZwclP4jYGj28tapkgMumvWtNWs7vbhNPmU9
NthFxGYd1zfZARrieVut+MEZSh0jSJOSCUQE7LPZpIeeg2zZGkhkl6ueVgNQBJKd
rvtQd28D01VUdAvlek5Swcw/VE5+Bv2HNPxBYEBgPcJyLkTJcRzhmfA6mBpUxph1
LMNq/hAuhEF2RQNaaYwXf5tExKG6RMUimRFb+fIPx/HnMAA2UscyCd2A9fUrK8n7
DFMv5fP2qIA1lL7QjUgitoNqGmsMRRruQ1Qxg+A47aHzmx4193CyVPMFtQpDnK9M
QmPZh6WS211oAWqlbjMZYjKk/iyT0pTx/EwiSZyTwnIX+hEVl9XVNaz33lfFMERB
hODzXTjwMLUIVkBa/y2aQolRLi6o/rK8z23RS59VlSIv1Y+dv+vj5j4wxYbaDnZx
s9BA8Nnr7DTQcQu6E1dDIjN5DphIiXGpkWa8O2SQpC4wTXM8KprurpD7f7KjwEe8
yS7BH0vfbSQovVV6dBqhOAzAylR6QWmDLQbNViDUQBXUCSsXmXJ14KMi4egSX6UG
9Akdq4ipsYtmakBnakCbvAYbrIxZ3ZgAzRG+5SANKwZ9GRAC7Fn8fwsHDMBcFrgJ
cJpwMklXVkMpRKe8yhc+RqsIhrfN/K7c3isTrc11dmBiWNB8x8X6SAdQLckZZWQV
G9umUcpV3tUUnBK/goVye/dOXGqYFiMVCJEmfXzDJMe0uyaFfXOXWoMGt4nYTgvQ
z8kXkCt9+vSnYPFAOe+ZkMr2SGNm2+2WmoWIDhtg9ZVrrrTdlgzNS8wHVcSwARrs
tkriX/pl2gafbwGcMLgL92VBINk06/AKSAOfr4QpoHWFtqz0iKpNvpfpKIVfuoA2
KmoOkLmdlkKkpoSNK7zp9fWSTJ0A4sBLJk8RglFBD6V5R79YVywo4eTr/Gl5hnSJ
ZxffRFL6n3fP/HmPQNHI8E3SwhQj87J4K2vIcLCr8Hj9vz2Wj8Tw4Nak7MFb/ksk
5hW7d0Ymb/cKxiIahTKwGRgXhVKlS2Gc+T2J5RO6cNnTupQFcnMHxZwl+3hw391B
ZzoHeAdhGe1KnLX9WPIaSy7OFRHrYZnH9di+XfCPHvabKwtrmHQE2GG0WSKCoD2x
AEdVgp6vRNccwZF09zCwI55gXmgxMkD5tiIOThY5IRf6uzF6OhUAicBVFJHXliiR
UbJsN/venOSJemAQVFGhjlcT7HdpVv72x1TcFnZZmpjzh5IqD5pGBQaFxZSVmeak
U/HJV/MOJi5SdCU6id8wNf98mJL2SbcOCFa5o4MIiViGeWMXm+hw43tgSYiE7Shg
SlVKP7u2aknhudorklJ+4JVPzsRYc4jFevoHoGvIQKHIEOj6tgfRO0i6aSOQj7Jc
ov9JFMMhkLZJ8YZPtITavcd7R8zGDoVAzHAs1dBp58svGrYN+2cgDJMN7Havik7H
/pbfuL9YCzDMa/4U09+krrdschHW8EY+7h1Vfv46O79gGx5xOYObSeM2bYVRq8Ap
GQRKcTfwfXW0SwMnSM7AHpk32NAr0dC6kj8jOUBRZTomzwVcn1FycMjq7yarpJKc
SokzC78lpnqnabSCLC8ZVIPAHXNydOvXkVkOoPaMFp22XfzNWookcLe1OdHSne1h
X4jvfeGqTuWpWVgsb5j54Zp3KCyCm8B4ZT+cUs18KHAK+DfzrpO5hDz0gnfoy3Lj
yj/7ssyNIi/NlBq9ooKNF5mmZes7DZr8hQZzUyk+2COToo++fjiLGv6klhuFDzHQ
iM5honfEd7VDucJOB2u2a/28kUbIWh5S7Z/OXjGkgOi0B0Z8xrwtpttu/ZqnviZk
rbvUf777Y5+U+KrL42aV36xRwrtWGDFC0vWlzGlSHRBbw5PY0xTk3D5feVdX1hU/
Qw9mixq1Moma1F03C9v6lRrMzAA2aE6BUXUkyVtzXCzynq/nG067DBNHoP1fcWhD
eLbtGCXk+lGVURNeXY4mKmrkpFgT2HZW7TrMy496wlvp6/EzNli1QgrAKVvxmbiF
kZhAvj35CdMQPTfAiiPcH+leKcFdN5bZEDPNkeoDcQ3BeyGPXB2hygU68AM/YOsG
oOjSucpD+pUbtBzwqjaEPXyW2vob8bjkwvMt4Z1vMgc9Ap7eYs/GNHOPCcCJb9dH
zzQTdOoCqJmOrWbluygvSuhZ3xbjCaasVyNL9BKhP/guofZvL5oY3VcWuwGVJrMu
ZL/KyVSSrFTA4oTVw5YINQMcvuLeN4EG7qtXAVPAcJD8avAe8lHAzz0mVBt6XGh4
cFgHL7mPOLiy7+wIELfH+U4EmM9D4+tOVXm4H1LjichDNRGNa3dJQzfJM7HGUdP2
RtCKK97gLepXuOZ4rLJelCBILjxEH37IeFRef4s6BdOamJ2N4a8MnpyKt35r0h94
sDoKb5AXsMxzV6sGsLVzY5OTH9Ctd3tI9/33sCZgis1NSo+01EMwtzGaU5Kyn3ae
iGEfmsZ8GZon+CDn1Rejy86KI2yNNq4AcZC82pIds/EEM0F1KlktlFBdROOGghnO
CYMv4QFVqQl3wlsYCLIlOQZon2kObJ1v19IqKcbmaZqnADQQKG2M6DvDyoaPqm46
Ygnu0MmOQ0rgZd3NzlYLviMqTerP/EJhERP3Ibpdh22OWDV0H5OnjLjKtSdDkMTd
hK9ZIPCwkt7U+ZMOvcRwwTLTuR4j1Dsi6I0tX1FUIDhrZkaPZGAXfUWUgOjVMeCe
U1bQ18pVf4VfeMGB92KKjDLuumzy4uVeXOHpxMLJgGdYoU2mYNKjUBtrh6NqSgQ4
Cw5U9osoDKapfBqgTroy3mPnS0SnK246nXRQ/q73dB3qO+ONFibokUbY6dHNi4v1
nyMw/bvoZGlFOiPcAUkikj9GPlzsvdwxeayL0Bz6bjhpHm50tMVdUbkF/ijVRZQD
YxjKab06Z/LzJTSGyAeNoWeuhvbebHNJ8rKFVxGCT7xuqp0gl5EBz4J+uaQ+29xN
lO11cWfOa0oSFIXu9AtXo94NENkxzUO4/irq+/lnL38tipl60bmgmklte4vERKIZ
BLfqPOdH3u69DpuWeulCQZQPUo3KW/PyzN3fspLcz5o/5DJZsDAGEbFhCij82Bef
VoOBeuWOk2RpohwM8IFqR0L/um7LJNKQ3TZygtlLreoAO+D8CH8Er78JgKq/yPsW
7CXTDgRkNj5eJJZUN9no6I0yZ0S2YyJLMZomuvPCYA7qfL99exp9l7gd9rzs7cTg
gmAnOinNkd3YgsFbNq77koDB9tUdTFYNOJA1Q9RARTg3FXhQaekKzj2IdRzmqKQQ
o9SiEf92tDFHwrUoYmSAD0c4rkQI8RhklVWe7v9JbLoQPzB+BCaLSAvrF2JiUUs0
RJxqWGFJT2U+EDmQlDhN71VYRuBJ3imiYpxQK9vSGbfEt1VwaaU2+BxX9dMdH84T
bCu/qT6N2t3JS/bdN/3OOLMoNyMg78/ET0MPvmimCg0UqPJvY7Ouc93v3h7HE7YW
epuco202E4gQ8ouuRpUmNz7FcWDNyZVxCrir+STQdqasokPTIezAN/oPqnYmGUAF
+ioiwMms7hidYLv+2VWtO9YrnVouTsWcnOp9NdtDBbut7wdGSgdC8gmaJZHLg3GJ
PgLgQeBWc/LsNWk1ju6QtfaDN/xddw1h8Ak/ZxXxZaLh85wlAE+9+HzRHNW20Nku
1MeAgpRa/p9qb1D0U5qmCQCUcjm4sXOsS1lLu4jpAG6Mm4G0hA5H+mpKi6ue+nKc
lpxCjPHssD7Ong2lUl4Wvf5ezvZYp6x7IKrQVd3XX6ggKnbyyUuolNCLPFAGb4fF
gYrZGXW0/U9NZiWzzO9PekCvgswHInp6xoWCJPgy//KGcSkLNe25FjCBvvKyTQan
ctmkJXz8QKmjJMgJXY9Ymhun1r2aOpQX6MTU1xg7lCfnyxs1nQwIBVwyyY4eWF4p
+qxaO3wzAJMK0vb+Dy4+HLMF5lfxiKcq05eHYXYPO5v5FYAGduTHLt/TdbSFTvv0
dA77Jz3fn6mPTOzCMgyP07wI2dAx7lexPHrXe2MzdqAQFXAnibp0qNERxM/mWzH0
8ilZxaTDs+v5SZUZjGM/1JdEzRlA+9RWzkG+Orvv2jO9tx9cSa8w7Mv290Xumwyg
mtDgc3EDh9JohWpX3FW0YLCgecqLpkvlAySLnQYw/yyvvQMjZKq6uNPXO8X6P7Dr
hzdfEv5bKCfR9vcoj8j0YH0TeEz7+QJ16/hysi3ShI60N5dC/Whjl/Xbm5jVG6Aw
vBLMS3sHDRe6/oZMnN+xHGPN5W1vaVXd4+zlUq/y1A5od9vhzMu5uvl6JAWEexIz
Nmbt/j9fFpwE42izQ6ZxcaIbEK0Mb2aeqNdpCbiB7qR7Fr11irE0wxdfwEPxQEGg
mxq3VexlX6PWcfBGYuR822IubyFW19SlhoLvYST83wgtxtEn/cY4pKTfIMchMWvb
juky+g4uPuBJoPOiBxj84oAMed1Vunzhu5eALt0T65IOvm53CxD5m5e3idu5CeW5
vwd7UJJ6dZU9BzHuUyNLoxDpH7Ykhgtv35xmLx1R3c1qZXQilcU02jO6WW8Qu8ie
ZXEhubYty2B+HBoSFznelVo4m5lMMN+hDk4GxwW+C2UgY7Y0jXmmCF/sAD6cfJgI
3eb4Bj2xh3RBTNbIGh7zOsy6LEJN52Ai+p45RQ99rRdd1U/CzeZky/D7zODK2W1N
vV5l+7i7UZqS50QJ4E+Jt6FVtEYT8fzwTv3o5Ro85aapl26BAYn5X3x3tdg8Msce
OfNjsGgvkqfFunJAOccq0W145AGyubeIBBvhHRqMboaHUnG8H46VWNTIdCsrbIhW
fCxw8/BLmQh/Q4kjijwGG7ljD8Sxq0rRxVKAv+sAAeXcBhQcbjmQ94JQc+Ja2c7q
MVhzWDwoojhL8eZdSsYET36w50q7Csm4fvzDtQWEFUMIgqxNRjkUl8ZT7BqkT6eE
GLJNeRDO/UlZOZ034by+F/1ZyeyfdRhsv8zzsZZQVI7qDMC4vkFwzvVvnrlAX1oX
05ZNpiFUa5uWpduJZL6Fhl98IFNOWnEZP/7t7Rd2rYk5rdRJfmK3W8o4F5hwnbmP
q3qC1tN5L845Klz6sRnwq5zxvZTc2Ec8zbqLu0smhco7W1HavKIvLujOGKonTJKB
gAPxfucTFzzUmKZvyinmCgP/co3mnuqc+LMpVPDQUHy6Fnik7UClf3OrjuSiQVqU
uj7eEm+NzMU00ikS8gCDO06/xv7QqQeNdHYOaZQPtEpcGeqab9XJAxusFsXet9XN
Oooq0wv2Dl87VpyeArsm8sgt6YXWsSDg303R8I2hRfNumoJrgsmPr9h/GFVD0W8D
Ozs6iuB4EukugCKDBeMQuTWISUdXMhdzfZf3KXFVC/DIJVpfVf0NKxVhJURcXPO2
yKAttAbCIFnnVajXNOBPF4U0yr62Q9B9CrOKcHCcOUpBg0n9TEdVGxwyGmSrns4i
aMvTnDU9XI+PbkK4UZN1C1f1lZxAwht6e1OnISU5PQmrXntiVDPnZREXB3PKGIwt
hPbUThzjxCAHZWHCf3UOlEdkIAbKxInGonzRf4itBs593+1nDzcfOoHmdJVvsCqd
yjOld0eaB1OV4K4kMhKnrtO1o/eaBBUiY+dzBLpvLF41iDfEynDnbwVzyUPygxtV
1zCWKC+AMyIhdWfcBq4sgf6qnPK+1SyuEW4b7uljwDL3WjbBenpUOvceUxBKAwJv
usidiov4N8YjE3J4br8cleZAe7uMivFyDbtxkDmYm+QueUGySaidyNrBs1QmVeh0
8FPGR6ZRsWH4gvPFk7uwwPrQeAcdN63ehNHhtHDYXWC+NIP+8NnV5Icm23qtw+oc
ztIOZcsirFlhXEmaw6ZAgbL11bZ8zn/XdMV5i9shprk2gHYTEoL8JksWncTlcq4V
4puIMR/ZHt18oCRyl27e7EsMh+xOz5plBbuNgLsIymxJV20AriY90o553hxk1cYb
3vbX/PK9p3x91j1BtnvbhCKVtQiNbo7zufxPHNisQ1sdJvkjwgQ4tm9Jpw4YGw3A
mzqj+VD6AcawaR8LMEcveY2tDae2Yvk/GTBBDeYXNKF7UPKXWwdWo8tttXWRWPnW
8ZwFGT5SBi8j6+dDQfFq6Cg9xRKp+QDdi/D+5l5eP1cc1wgY3sBQFnSvIp7DtZmp
7W5JCSdLqrnYx0jr19z8L3j4hvLlncNz6+iYhdQMx5ZjQ6F2rakdFKwBNtNF7xUW
jTwzzJLOL/+SJ5XvQ1Bfs63IEOF3zTkJPGR75gzyY2qhbXv+hQLvJaEbYOgKeBb/
RVrNJJptzfOI306qevUoP5ATpDi71lPqqojbVxfR9vM7kY2WUVpcSpTCHVJq6qNY
+FcQhkInuM9ltIaxibSvlD2thnaumIpdTJL4i53bRXZTxBv3BEA/erlEG6/98r8U
dL0XEpgB1lvAkj2CPxjGiG8hAGxR2qJ9lqs6QaRJZslIA4Akgztcji/cTp6eygha
lnFshtFpTshgWjw4TcFzXHEEjLc2pTpxGU6gYOe/ISRzfHHYXLlNyvZP1YNV96br
DB80+yle32MkQwxHBL5WS0wNz1LZt32E7yB6M2cexHlhkcHgZzJTPpPYBMYfNQ4L
V7GrmcXQrSikQNF3cbRY+Q==
`pragma protect end_protected
