// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bbncSl0O8Yh9y+mflBIFqmw/hgc/istroDW4VxuKrmgJnz+gl1L8aVkLaevxFo63
Feut7LPlX+ExDlEqNEFgWXm14tbacvT4FzCmZimI54e5ZMjMGniHM2vMrm/xzbH1
OBtx4ID39xvld0cR5hPlzjujOyVLYs+xbJwjw5f4DuA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19712)
XCJ/TzM7tDtphA0hAOF9zDpSJScyTRaJWbORTJ91p06UpCeZKaGO/sDnzyMLqIQr
xgPMzsMT3QWByASrgKRrk80gatN6aIOAMDotLYxKUxz8Hk16UgRNG1aYOrr1dm2T
UyDESG/4Tyumx/+Q56AX+NPfI+sTf+qSJ7u5oMmh/ircTmQ34mDqOYCohmOPJT8S
fuu7lBgxX4/xoDUz1Y+Ph697IPvECLtdY4YRNbw7G3kl4ZCyHbZCcSmmP0qqjFQh
SsPf5BYAFKfGxKg3OZA1+PG9+hk4P6lGthiPKEqqUM7Mi37NEEX5mNW+n+zSO2Z+
TgmrlZfMmaKmIjkwzNxbC2s4T/cMOkAr2NhQCz/A7fTTSdAUnAbxdKUGy28trI5c
WUJ6rKO2qV+lR8F6P/3vjIvWgPT7dmQhbV0tnu4XuvXoB3r/yVAU7qksuiLR4wUg
HSOp3kyGNJISnXUQAbTLXAOue6mdtDTD4GBsvfJYRyDQPjQ+j2/NToCvQj4G3+uz
vKoE6KbqLh6eLPHMjBoyondhgEJrFbZXNyB14xejbaluMGuIG/xkqhYFa06ghN5G
megQAjhhLOgNZWXFveX+4Xs2ouaCE/7gBgPa/6CWl6+6kvVzpPBKPnDwBSnHVV8P
KUQ45SyWgOyUa6Gz1dxnyJZ7wiBvXpUFzt32IIKBwpYNFmZ57QOaZhOlG7l0aPC8
CcZ/Pk56NQ2DC2SZA2fxPn09M/Z4H6Y+oNGUWRyJKs7TPdWafm/lcnBwrZMCZldh
suRtS3p9XMrSnehomep8uC3qxaF/tIgVgcud+GYZgcTQ8b3nMjSSI5cIgzzJK168
cMpMyXPNaaxOL6uV04pWi6PVuFTPotEEJKrNc1ko+IBcGuR0G/UDtrRDjq3Oq2Nl
owKefQlBQe5PZyZVDIgGit+TABGfs7ivCUHgh7LZEIIEhcciYen9F2P3lyXshc7D
GvMkK8rNiH4/sxU2p2parqL3ra5sbTwepaKfb6keSB3Lf29n9fGopPBDjaLRhpG3
koDcjNEpn41grNVweiqd/BfJaPQs75VbktSeM8RiO6LOdpOkKn61+vrCquDAfx0X
H2uCCaE/Vo0tMIUyPSm0cvtHc9qT7LxAwAF764ldvvxAm8L0eiVh7lw8NPbmydLw
Nagg/CM3ZTuHJ38S0iuljFaO73QZNARIsMiaxQQQeaJ5T8jYPXKmrsAQ9FLHr74I
6qSRyrb3nW3uMVIUdV8zLlboF+Hz62Dzc26fVvDJxmpRbBNo9dHC66HWR5MDHiGt
t0Pdv7Z4mrtj1alaGuT+he3FmwhfI6ImBeItjCTLp86iGa8h9Oq0r3Bt0Znouv0B
ffxMY91mGjKFaQuw0HAGefRfI/hDnJw9veluzM6Id1gMB44n5F7CGCVBo/CaW1ht
tWEGeFRPnikBrnwrZwxQTdHji0A3MHOHLWp2+jgFbHpVneGtSxJCCwuNA0ARtyUj
jTiQFWZXDRYWqPwJsD9Czxk/FYPUbEXqYa7Wc/ELOq4VDsX0MNs+1/1P0rSFoGRi
Zgm/yoYvZK3Qw5w99NAFrpuwWfvAMNeBTSQmI+gAi7FS0uqp1h78Xxk/+2hHTrsp
q6C6yxzUVYYP9eOkfMY1eXZjwWjhy8qTvxeBjQGWiD8znfXwacg34qdeEfIwabV3
dcGzrXdsbGq1zh2RslLMRja3S2yO4rEwZEXHfHcu9bs8XE/j6hY19q51Sew9adC7
DspkLOrRaFCgc4+y+E8s6de57d95TkYKeaAZ/nMbEP0w1XLe7hQs6M88FlFRmXx2
/r1ndorUs4tRE7TVO+I56bfSrerJA4F4hiCDqSNz4nZSUOF5Ra24JEGsUEooDPPU
IZT7h7Wyaga57bWZD9JlwNnpmhvMp/N1b9M/C6eaBlGAv2HJb5OWnqZhn2nOcFNv
XRsEfOiLnLUEQHTEAWXGBWVHkkSJSr3aVRhb9LBxEeWWqu5cRww7WBmJjJDA/K2b
l1d7zXoKZrKUR+oremk1a86BGJDnemPPMUFOwl1oR0j8dhvFsRJAXqmqLec4YspS
PbRW146qwQaxBGu0UChC1Vl64kSbTdSvHjU+pEbq3AgwYHmqpNJKr6w2cHTNBiRN
+k20vjWKO443Pt/459ttrf2hNlMKtInr3QduxitaZg2kUBSvOdWQLL3oBO8AQfW3
ELjDBQEJAYjdYf+jJJQX4BCWYXhJJySAcMKRY72ICmLn+YP4L1gpt1AZT7J3SyPR
x8ZBVmf2oamDh0saurmCJ2peR6K0bP57Q3DZsYXU3r5/l3yHnQUPvxSIkBBxpota
MoVrQgzP9LZBXpA4nT4WDkpPm2gdHK4mB+UGZiYgo0100Rj396ju0GalPgtr/t73
GIny+rmoqjXa/ULsb3WrnLaee9Gt1WbuBKOiZUSmpu2P7MtL87p58RUao8mEpiGb
1TOq38ciMHyeWASs8/nnuFgjbm/wQcFbxlNbRFz+CugnC4r1Z1N13Y+UGj9drm++
B43V9X1w5wHqK19OZcabQikVmelpt9mBArX2krkqf+QlePVA+5MSgKA1fM5xKc0U
20ARu/j1Rswp0MZUSY08WiHv/0T5soZhG8TfrNcHRZ+qO/p0BxaW0z5Mnbw7Ii7W
/jIq2ZGenaXZQzwzaauB3Pe+LygPOkSeENceIRAAIm4LnI4wf+QbVjvyhzgfaPZP
52gD3BWJwBjEQ1ULcMn0GIdppSvIP6+rHU9ye08rI+9u3JJP6PqOEJxKnsnPACvM
rZPHbMroDGprkiYfqiEwtxz08zKdn1w5rdn9B+xsCawL9Ch6cjDSNLqp52SW/kqI
0Z6HmjhY8ZxsqjDdjxte/pT7PnYmJD6wfkJ03oLIQnpntZzLuJKM08PV3XxYpUJt
+DCSyIKy0yxjKM3VsXLNOFuOIpeBQhjPibDCfrqIQaCH8kf8IxXOZ5ZusXqTiam4
+iJ1o8X+h1UOjJZqCBf5Fei14B1aN3qytnsy1m+9a2KjAEqDzUy9imeK1B4C4dKh
4poz/ozOKGKxGBE2SBs8suYsvkqQqzNTjtPHb4+ey94ebHPrCslEHT26PQvMJ6yQ
H6EFJCa7At+nj+ShzHnS8qV75/JcYpChqHZP6pRq5NOYbPSaMNklwM8/jxJRQUlh
gUiyhD20Ov5ajFy2/stRXFMS9+vAGKDizs2DwvlkiWZnXJPoLeKNJ83n8NqINg59
3f59w5uEodJ+qUdE8OTDYKlX26qqgqPp6EXAdZQ50dh24hfCG0aAuR1W/9c5V7/+
KZs9A32MgOFmbugOGDxzYMEOZRaNOTtHMSC006kPq+Hnq7J3OtrbTrG3EUnrmd08
xO44BlRLdD5uB/e7JXE0E+RI6GoLylNCoP/YPpkkjH9WdduYfv6EK85vJ3CZJ4eT
jEgSAxJB39HX+Hm9RBsNVxZ0jVtnA4Vrz0SwnhmJqrjTQ2m69tyvE0Xtst1rbO2Y
sIqEmn5Qyf92A42QhlQPp3PFUyntELcS+R1fyzo1puY4P/MTZPm4svADslMqq7Gj
qDdmTeNY4691PYvfgkT5HQ8+YEQyMzKpPZ52bKnei2YYGziIFs7i1Btqq72RA4+/
9EDQnC2cGfl097weSKAF0jXg17yqEZ93nC2X5ruu/HM+GpDdB77iYav24/uQz9mH
JylJ5kKej73kRGAmfx5FLfxjDyQoo/IXqX8mm8sb7akEQwRuVtZPNb+VMXJcqr6p
ZYSxgL8tiRpamNLdkYuelzKn4X5U8V//2tWFUZgLiVgQulx1dovWUWW1pWcWAOPE
sZW3NjUt39yDNgk7htzGTUtCXKxjPoxstjyQyMYL7Mf+UwMCYP6pgZOEwQdOj7zu
0gYAZUEmwMxEqrC2RH6b4QSDt7LfAqw8VcxUBQpG7DetI8WePtcaNoNz6AbD34mC
u65o3KdGad4/6XXCUbHSiaXE2YCWs/D4UrEkL17An6PDjW5vpfh+L+iZswmT3l/I
HSeU/YDeXUUK5gWVHvcAQ7RKhW55k0iP+krEETjEwCuqem9xP/Fc1m3rLNlnH0lc
oFZSm7BQAbCqOYLqPOqB7z4p8SOnytyujxZakz+XzB9+OwFUrN69oSGxDixAjFy6
t4gfd6zFKEgkZk7oB5oki342SEXNO2ueWO2L6ae5UN8Hd/RQrrhr/9nREWImENig
9zgtEKMt3mNWgMDVohg3XBw/CxmlVMNnLY2snL3Exz95QW7m6tGlLTF3v+XZXXFs
doG2XFBRddZyVpOCLVyNsp5RkelX8KrRA7IMxx7jutFTtgFZTVpYB8TJPIqMibGF
t60Xbed9X+MEM5Lz5zSit4qDFQ2fNeRnCd6uRFaVUgTmIkuJlFbGOIvtWZUlsrj3
IM9GyzAnpP56WXTNOb1upXMf+yo5rQRO9sHqUqjUE7AyvOVr/YT6mK1VVOaSRS3A
hMujssbWFUawDJ78KECkasG/ur67cYQDvbzvj5PiWK1/w2XN4f4ndJRBb8DWjRuQ
QPMhsIvZepxfRFpNnqNXBXKc/cI8qLqHTKBwkUVCdQ4n2x5Dhew/AN3Sm7VwPni0
wkpHyCZR6oqamtyYIQ49ZEiqxrRzNlfMLPJzZk5ur2RicMm6D1UnyQDwsRlyLFbo
Wqlh9d/Jy5RoS0RfvswEzEl7DYuSDlvU66v0Y3Hmfo5Wz7cAEWUOUAHbqFgGp1kl
yO66ytOrxig3xA0MAJfKyTH7KqyGJzgdmdnzpsdvx0FD9FAR5bll1i+1G+XlFDQ4
pD1/VxQMl3a2trsEhJEpdgjwo/wuT63wpzvllY6TnmwxvoIpZ04/2zA6rE0STF/l
UX+jktD6BuV2a1bal2YFz5S0j+SowQWLxCZOSuYg16Bn4jdeyvGCa12x11i1zP9U
rkCBIrABjX4A9KEpU9vpe4OmS/08TlSYOBrrE0NSKG39wc1meQ3pP9T3QHtjakMH
Q5lVwG/vsM+r98KBbnkbpu5F3m2os2iEh8VIqEILSvRKuNZY3cZZnFO+stBl2yr+
e9clsO0blzoWV5xLKx9mDdgyTBzrIsrEwt6lHJWG0kI5YgBEq3oqLaivgUhQXX+Q
W8xs1KPjcitRBta9y9WENy9u99C1Q0INDnaC9LOjxAtvGF2qjHdhCn9NfUYS6bid
3otvjPOJp6Nk7my0pEAd1zLDJyPpP+y2+F9OERjzA9VpT+G9veaOHCMJkAJGD3PM
m5/HhchScW63f/oeQH/j+uRqX/Y+nWffJH53nY4QOugnS7B4WrNxszjWH18ldNhW
bePPqhDxa/zOQgDnFk3lVTCo4hJlZdfzsewbtBM0z/ivIRaZiidVzHcGhC6zzUV+
/bVeIRsULXP/TJbbi/VdvTSiTAokLkIWiMtS6FKDPZKP0zJDfop7lqjl6pnIE/3X
kao0yBMa5cDazqI/FjGvF33JdNjHJrpoXIIYeEyIaZ0em0A1wL99rx2USwDU816h
vjs7Eng8SMLeuMf8FXnOLmrfw+qcZC5OULvTt+qvQlVrjxgcl07jMx3WgHs74clh
IWD3D2L8coG26epCb2Qwybzui78qndcSmUMFynkllxkrs5pmvEdEK8sEjarMdbL4
skCgABYYD/wNeZ+VYeh79uMFtEq5Pz9UxRv/1nCcFEZRfv6jHazGx+/bQdZoINGr
hSIeGoLjtluz0KO7D2U3XLdx3sGtv1Zx9T0zKLhNH1PNHjX/640u01FBh/R9827I
Xxfrc0NptDgGmaeK8PhsIhE+umAKiNL3JVGwNQQeCFTP5+eVe6qHdyvqFgK1lt9F
f+InQD5R+eWGIYhjdtQP0LPDXDQkB74bUOMfDJXGGAjFZj5oeqJi/3L94LMkA7fQ
ekeMQ1lQs9rzqaXPWYuxssD7Ll+XJ0WQOuNubpdtXDo4487nW8nUW/gXj35BOFmU
dN/9MOdBA5h+cpIfhdwcKJEKco/tGPo1dgTpsTyCCp7+E8ALsOAKVVAfJC+JUsKa
VwYZh+I2BpdlGaDp84X0zbpQaEtcN9fa+O8zCOdsqLtGGpVJqPxNM3uPVUvMEKoA
xWxSLefhOqpZZYsBsseDA2H14pCyPRQwiMfFaFQvbt5hhmKd9ULgvm0yXGbS5f2d
Rz6km71MqOfqx1GLwX866CCzFQNYOT0CakEdljJ3fpK9I/3wn9j7JkLMtHpeAeIc
3DC3XrP22phH5pGTIITeLmT2FwhgBiGutsZC8xsLy/c7qq4NbPI6673UpjkgLNCl
VdkNKVh6IGDBto2LXCGhn9EN8R9kh1unGs8rmjGH8unxDQZM2kafSotprT6Szg1b
D4QS3K47T12VE+XiKfVpS8WMmfJtu3d8zzHnmB7fmPRCBlFhYsj9Ogtm/ifs9O9J
bm/raNpJv45Fh2KapgZDpKTJ5CzJ1WrAaKdpT4FZfmIR7c/C3IynVn4ilzvFq1V8
aSP5+Rm3jTWQBGPlGBXSX/evq6xa4DjPuo6scz80eNqqUsO6jKaSShZNeVtg6zix
1+0M4Z47wKA344IB3CgYaaKPUx6CVtDU2y7C0zVMc2sQ5RY3sP1FanVzuAF08udY
4SPTm1FUeL/1pVUynC7jPaijmvKVUWrPtORWoO8BswOdwRAJmyk3UWnhqccSS/w1
NxTqkkfbs2xe4lGU90wkBSjDhZtPlZO017cjvgZzcD+miyGEHL8C49b/JXnWtpoI
lfdQdkJcNZRua94hi/6mSVK67Ysn8kGhzRFDGA0j73bZ0cep5eB+DFUTRa4rWN4K
oSbp8QDkW/uWTvD3uLhHHzdUwjwHi07FZTwT1m0hMQfjFlry+tq2HXBbw+3F9MrM
ZWPV2xSHxpxGzPViGhohDAT2dZRDKSRy51Nfy4cK0b24kyoMYfPxy9QIn5/H3ibr
QZ8pZUp1URbCNJCZsTLkqF5I7NWv7Yuv6uWJFWEj61yOY672hERENmVQqZr2pAw9
i86yO6Ra+ELCBUQP1N2QPApqO8IskqGUpyDj1sxBUsSlE0Qd57NdIT697MnHjcJo
UByd3WVTV0IbgoTggeVy1ylBEUQ5VZzfcxp6XHMxvLTdk46diiCS6XOZxb3BHa2S
XwwrHykj31cfDtX2VdGWcRNHE7CMB/NZJJMIPObiCoct9KuBtMcidVnox6CBivpZ
wDE8EE11TRH5s2TLUw1jNmwyDtFw9lBgTVAAxqy5pZuCphQR+ZsEZMniFazsgvLJ
NSommwIkmGZpiCj+zy/UVbPkymcj68egzOKWhyChBoOrd32JaC3CYC8g1MQME1Pl
NDGwBMDz8kQCghEVF1ZI3QoIXCcrHaP3NlikMGzs6i0xAcmP8cWARyTlJ3I8JhtV
g6lwagppdjO1og9mwpQZEKu7d3mc0nELD2BDgnZxvIE5b8MV72BHlTBEm3yk+hXx
loDSPvnjjThVM32wNUemYTbUeqRnJzOWhqvpAYRD/jZEfn/e6e5TvISDcnbR/qwC
FvWsalFJ2N6vLOfsXt+4d24YcD1/6+O39liV2vEmEpuvBm1gdkWQH0EXXPGJZwn2
n+hWmGeK0dVBA8pzom3++SuvH4MUTsh7XdCJr2Vjsf9AuHY9g/VfpkgowkHxL2MP
xeZb0j/4RXutpzrmAmwhsyk3ZbC8xIhhzBwjpvLfHfjB3Hvm4H6V66QS6cbyni3n
MUzNUsWztIFcTMkKUd+nxCpR9VMubQD3idd+wZOuIVgtsBH7uGER1N8jBNyTQmEz
L1URgMzBRq5r3+pg3MqwvhRtZF3HhDJNxjuK+FaIh6LfgIl7Tbxq3BX81/Dn2qZt
Ranpq+RCPLMLTPNfM3pHgkCq6VE9fQB2529yP0tQtRiXHrpL0x069GUn2iscF2r4
mecEd04mZbHkvf4mWD30MyhwYNc/V0nuDxghnzTuxqfThOCTZNYfYF738zTO4tU2
Ns9d6qJQYR9iPcSdALT1ZoqDtL20Zb6fp6MWFD1K5X+N364PMsO6I7yXmD5W29A6
2WgHZrbOvhCnHctF+A+LxgzvRKe6J6eiFdx3s4KY/j9suNhGWPT93q9vpJp/OXVh
n+CAIEUBZYSy6JZiq4ItM6ESILLbMs1/aKUe2XmPqeqobI9r/ZV/29xPg1x1I8cN
N+t6vts5StufiQDwbN9oBlbAoHq1OTGL2ho5SgtN9O7eknbALZJ8vnpyV8Itk6Ep
zJRoEtnmBwgpXPjLDnfiUGaLj5pod5Hy9jxSz/sh0xNhKfVQAIpU10A9ePKfXe2y
DF0Vq6uTgxpgcSV8DONhdtu4X060kAY+vgzy5TH9BQQ8+xVhm/4Y+naNwg3nYeJH
M1+dkMA/tnqUKuRUZyNphGnHt/jxpE19ezs7iPL04qVJXrOTTvTYFSNcRwsX93mV
pxYDQ5fbSunPWAXMJ2Id1UXowIfZ+G7RUGonr+HHzQBXZWBYY3YJVKfuEWpqa7iw
NNDXOCO3MKJTKnVg3ou7f+aMyMm2ah0EJy5pTXGVj9iMsuHzU2qmIvMzFrCyvTle
VEn6BUpkUKeyiJZ8BLUEMv9XqbUtCgRpQU7xKpGjHDqdyDjkpXzMqgspRP5/rA0m
FAVtzdKmK38GtY/w/2QXReC4KTPYg83zzApSA4fziKCWAaUsV/EF3mhJLO2M2TsK
BHOi3ZmtVe7dI1TTVSY5/WuEN64wVBRRgEaT5am78yQBRl/9wyGqa8rMcb0gcZb9
a7Fg1Z5gEDSOJQ3ddSK+XhwJmdb5izMJwHBJ0ssHAKcTJogereqa8UIzU0oyfdqx
0b5HPXTsSVvyNj2m1Jd3NIgQmSwS4JvE5WLLAMoflOvilN3tL2qofdmhqzieI/qZ
+n7MphqcYHvbyXfGmpYYF56T9XDC3PMe0YRzLx5qLSO64dLKFOWPuU+b5P99TmMT
2cySuXX09lSSCH75nDXI9mSIEZJKlKZerYUlZ0WyykGBOj4FQZTvmGeXZpfXBtVe
kcyuE1+b53aO3FBYMcH6xCAKoKU7a5IWHV73bYDDOlRTqPc2/Jts2udZ3YQZbSYx
lS/4IESfRWHXOIZxYKGU9ZCljKoC9Ja8LHbhKbE/xLK2ou0J4rxWF6VcxEmDE2As
Bv9ADCEMvIqynz0EZKlFm9ImLuicy90AZ8zqLZ3TvVzjsUk2VBgJ8dtySW2o66yW
Vgirx/269NKVpmisJbskkHrRejgUN+/+zOY6PFoTn/SjWVwOzuFd8eBAd07fUTmW
iT+O6ArshMYNKUGdOaGl/fQyNpQfGVR7tap/1tVwt5MF774+CF3ShmBGTgXdocKW
0dIXkjKXBwA6mavOgrJnfztaKxcyAGO7DjxhKM0A5XvxzenNHr5wQ/hEZSlPiSc4
DJ6oYwR1V/+r5Yn9bdK9gTCrlPVYcWqjXEy8tig6Ce5DPERiCjY0FLOaM063nq2t
GN9RS/0Cwhq3fjA0Pzgs+uO9lTOHiywaRMCUJdMV5/1pNrlukSE/0G0c9n5i4I4m
4d8+xDl1amK7/n6zHbokTXHJnbM3X2VVJPAwhsYUpW8BUz2mrAklIna/zEtS9BYN
q85Aqiag5g07zY9yCEvlM19ae/wmAFd07dXCziQ/Laqw9ANdR3L8//JYi8KJCnR8
q+Huh+zBDMLAvtpSg1AsSRX6b18JguhdEi2N5rIDNXTyKMhnMag728vLKqEBhZcp
9PjO/giPqDAy9x56jwoLPsxgTU/PJRlV1GG7WuN7qjqjxwPfPrcjfd+x1Ip9+gg9
aYq6kbDx+TgOg4tWDySf7jVHoNO2GPANEHkeBUHRFITOsjR3BXFYxWJyNXHc1C9g
MkW9rsCJgAPScC5ZQVKgJS4ibLTONgKFljRzFyYKpYs2MojCn2+GyRjHLLrmVeFL
XFsrPfpGScyxx+/h7q6QD/bPq9/VVBBGWj/bP9zI67CUrytpdB4yKVg2xBfOzrGQ
X4z/fnxKZeThSkCFtONiS71ele21h51J/GHZKRGDtwQIf7JRYKnr058G+glae8nn
pjCYvMJVFE5NvBV+0OF7nS3WD1vvTQrgwdaaDL3coHgRGGxTjeXYhfxVgz+X4PPr
di/3li942G4zhxZnMekLbMeFUD8/FdoConzfxR+FV+p0zrZu3W3hZcNK9uYDRRwH
VyV9uFAhn8ySqYviMEzTy/35SH5E6WlZvyrVlz0cX3z9chN6MEoH6pAJhu9XTlCm
qUcpPld2b1AmMDTGckj9WO0SrZLSiBBSHLFdI8l2KKVFPHDZd0E6etlLulbOq2Xc
XkFmcdvmro2sJXVx5mn2dPAgiMeawo1eLw7lcGJR9UHTuGTKlvp9IzEuDNXRmvCL
36qLKnr3lIYH+Dpah6ji4kuAzdi39uamQ5fSSzcfGeYCdjWw7it2VDZgrlz5RP4J
aGOWbO3G/7CpzfLCKYnpQCucVcpZrtWURXheekb9PcJ75dEhaCRjhNltqGZAKVPZ
0GMRUTxlW3JMJw6b0tOS+CCDXD8fI2VtSoYeupb39CzXLsxfOJIns+nh271kZB+H
vVBYVVHZng5R08vCfjl5q/yoEvMwxKwnZZ0dUc1LQ6BUN1aLG1NANSxbkZ5jbm9y
oiQe/8b5W7e9PV2XCn9uBpQuNp7MGR0c+4SuT6BV5w5UiQAg5iR2yTL1+1fAspEu
Pgv3TSJKI5tR843fiUy85O2d/yD5/mEBbPe6TM9Ux4jTAIgHTE94suZEW7y01Qqd
Nm9LinVleTwNHzNc0e00KY1p8z3lWhek4F0SBf36mqRNcEopkwNwkEd0uoMQLjIx
cjdcK7+FsoLGHlvX/OKTvef228VBOPbMV9D1LuGvlB0WRXCeEqykIA1wJ/FTDd9p
J9Ma7ImK4U/K99BkEIv1jK+h51di1Z2QPiHBefBfh8G4TB8Sn2P6LzSr9RsVulqi
boRfwScs5zxPwv/3KlEstA2ZvMW3tDA+QwTSgTPpZ6O5672j84O0YHN8CDqtZi77
EyY79FWEbg5WN29EgKqHb/OGUN+cknZMffZz9c6uli8ws0oRRR3a5u3loAcHQBkb
3/MxkG9oYnwRcZ2yl4ay2szK1QzUWXHafNwJQu1ECHnJl9YtRTifyB50I/WPDzIG
rZ9e5A0/VnXtjc5OPFxnZMUg2+nn3ni8KURqDB6KRTTPIvSx1nOcgRhmygqSfT12
0cAC5VnJehfMB6KcmIoIBEH+MdLm3lo708wZEkNbTm6Kl7WBEVk6XhexTuHiVGPn
e1dsILkj5seej8Jf64/VVtUg1gzwRlbFAFNz72Jh9CCh0mCjcQ8qsU01czCA5/yB
8BPZ955JizwSeWgXTPKbTeog79l3vhUiCm/okW3neQ+/+twNvP1NZ5Inlk4/b+VZ
weGMNF25/iCKaMMAkNPmfmfGePG9V9/4wwF69NZHDBHqCIVJORU/mOgsNjZlRbGY
gvWZhGb3S2b802H018+Z2FGLVfi9hbg7P66vynYRfet7qO69Dv1rOq+tsFdlzzAT
rOobuGGDi/jIJNxXejSnMeaKvHKV+yxdE1JjiMTufv1TF4ZXxJHFSxzgB0x7fP3/
orZcUIEqSrBab+XjzgRCQl4I+8XMcqObq40S30s3faq4yU+tIwn8mn0gOUPSupUb
kk/aH9zay+7mQ0v+ixdAHXAhEDVYim59lgALjYwdv/M43fGwe+++V8glsFQ9C7Xn
i4xATyL9tWT65lCuyljUi8auoI3MpwMB0SyS0M/P8g+JZvC7oJI/I3nJR4zcMxtI
woyGlDM4sArO09e13qBWZgMEMsBi5oOV87UQ9riJFbgmQbUXLhryIZmtiyBErkKc
JJTHv/MJEK+PSvnTJketUXdlrU+1IYkAeDCRzR29zh24ptKIIBaqtxVHg/s2N6jq
dE4RNtK45fJWDbodNqSVuXNwdyhxMISUcsu0TYJxPllJL7UmaJ2ly3JCnrOs0x8b
PERR7NNyEJ6srfXB8zXK+nb9GAWNXCWws+6NMUbNngF210kTOsMMAY0lobfhhERi
ZSVAopqJTejLn6o/EIPIP7hrwXVWEHCe7TdT0+/+AdmvUdY7yLeivNHgd32mK5wl
857SU0gSb80nO6bjfJ3cvFyH4XEl8BG6ooGfouN47Z69oF1BT9pFk7Du9JxIob3Q
s8Kn0Wv66c2hcExUNSr5EyVB4w06ZC2lK5L6hmIBg08woS9yOjgNzaJgKJBcZ0sx
ExupleL+B76GBOiipxKNDh3kVp2SAvzm2XKnE9yOmDeq+srMRuo/5EJm+bcWGGLM
vditmihHRbIyot0meAXQ1hrRn89mK/bVzwCljZPJpM0u6kR9qsUKOTrABuj/1GDH
vYb1hT6vLh5VQ3ysPo7qPu8/ZVLE18TpttngQZabjwcJbwI72hvJOUwo5HpMfJku
1zBCeB95oxKG2QQ0egJ6MNd9ubiQpyXfUwcXfXLZ0HSxdjAXNTVYXSF/m4MuLlvo
X+pxGTuSM7Q8bgex6xwCel9Oyc2iqOOt34pln2r3jw5aBAtXB4QYcOrVKG34Z4Y6
U6mCuabZj6/vej41ghfdRuDPZhOamfVcBaPCTG7D5AzAofuaNwRPJu2hdmZ0N1yJ
sgh+iVVi0fYehHY1DPc0andv5k0Rc6PflVxWiGh5Zbqgqcv7lpZ1IoB6QNdQPX7A
BESBXBQ6redWX1Qm/uflgtpRVgbSKXDjLcobjT+DRDu5OHluYLyQDQR4+Fwz9apm
FN4a8ux3D6e84rPw5nKRkbrFfN9SVhQdaj81HCM4GAsS3JBEcF/p856xdzv3ZAMb
I6IqyfgUIHq5I5JIGYO4OjLQnAxH3sOsmvDbo5IhZVJXRja6EUyUbDoX76HE+16E
O9qd4eEv08Z4bQzYCUyM3cjUrlnJPezQT9jnGFenRzd63mHoNv9LbvMYujKbEBC5
GTUpcd1QlLkkrIQrCzTqgrxjQ3gPaks/7qBxamoP9nV0OKsFrVCmm8IhuF9nKp9T
+P1Zwil52RVEjaE9wDwOrex9koJhVvBvPxRHiWVubLwtkYWA3RAgHMr8Yf/DuG2n
79evi1EPn/pneH+vuRj1CmoAvPBxorvZUqY6QLn5AhpEJCXiYMxL8GDLNCTotlYi
9n0b51SIIkWe01Nc8mGTuIaFJiNJ958M9Ty+AnDIN49IdSsGtuefF9NrMgSBCCiC
68Q+Jmfj0mbGM5Sr6BXeFTin169yh0bSyu5jHforQnud8lRdTZojC46OHEr6QtLu
Lm9/v9FsWyb1oDDlEm5T4FYoZez3ho8c1kjp3guUXxX4+2TzGfAnpFC80mq32d5W
Zesba87sIGq+yZojhiYTUYjgpjsv7cuPFu06iVN3facwF+LrnzNFjekLNwovQLP1
bTeW4VjWRBAJoaUMcvwfC7K40DhEJsFY0DkGaI15tcubF0YGWJre9ciwYWwl6LLv
6RRUsvr4kPoU71/TPcNUUI0x6Z6fYFdnmi3PaHO0fCsUThTGIkjcU6MiwHcsu5M4
/9DM+R/e9z8brhzYU2Du5hbxudiLKZ8KVFurvXVMyQ8f1hpzVJ74opkubo1vz5x0
x6p+WjMNMeZ1Nl0bimmGkFSpIHS+UdL+nzxI2hpMtSmhS+6h+94a7I6+y0ey18iO
dQSO8cGnFjRqkKNhFEA+2u841hjlyIIKPvJPXbjX0PbVClmXX+NF2XuBpxvBXiya
GxK/hce6qJUXi8NwYBvZbey9bR2rfndSgRJu6DHlUtytIstX+BVwvaY9GEaHYmeD
NeTAvQ6+UKRwfD7wkQyfLuIBcX06patY/GWYT8nZcPs0AWUAyXZTqAduj5p/NUMV
YhbNMXT05kkoUkv4/zfsxvNacZmna/8DTAtLzdjScLsba5coI/eXVVBUiJdfKJz8
2XpZiVOVOZKJki+gCvWXXmDoOTQILI42h94gDW3DcFayCNv3lYUiLcTQxjOxFeMg
99hsT4oDZKlTW1FWTI/mXbGEEhuBo9baF0Cq0oP3g+IeXPGQnEqbNXw2ATEpGjug
siIh9PUVqxGJD3N69EAvVFunLUOCBytBfz/2dksLYcc7NmcaJ/70XTTUA+NEb6En
skH9Uvd5UKSlSZsMCfOJXCw5zlrw2UhidjD6WlJj/W93YtZdUS2UtvDTlYrLjZTA
Z5CcuBn+lCtx883CWahI++pczb3+LZhvC4CN5repwBFN8yRdVQytVNOWgw7wgVB1
57vPOncLMjn/KLegzjqeSvaH64DtqIeA+8NIP+X5fD7ftl/oYep6W5HAEBy6UB5d
JkjGZVPcllqT0JGSOgf/WyOc+6iNDUHiEi5lxlcRrdJIMrJ+8qWTG/atYKiDw8V+
NAYfo1T1pDdvZZbKU+mi/ZJieTx6xu4bxd6W1UaKZVm5ceU2bSfnsaaW0dT6f5c+
TocsyMMdPPWlX38WnPt0QyJmlM1qB3BsB7Eo+B3FVvQnlW1kU8GoH4sgsOyluNxd
qisAHGSMKYBxlhM3ksiDKv2f/U+jJvjvVJfhQXI8CAuMlicEc99oopMnk5zXExQP
y4YW4wtuKtEUGbS1gwyc3TL3o8YAnGOaNmCYhIPpIb0eAkwyPBTLLfUSHeZ+YIDE
5A9q5Myv+2JRXcCZqW5TtaMlYWoN8/tuTLmAqhGBckDcR2daDs3cEVM3z4Ywfgmd
uIPjk/F0Y3b5V/AHtfXHbvlnJKJbnmF5kWyN+sgzB/dihHJvZmihDGe2pIL/djpf
f/ku/DGmR7Z4omC0E9uH+NiPSeE46PyQrieKUPAo7CQ4U5Q3dUQyjJPuKH404JrS
Q6H9iecQ7NgjUPpjUFgqlqDnIncyBuNw5Cy92GEMLyAJohHYI2g0LJvw4ageWQ3Y
b3HnnwvTg5qMOGXruKsJN4rVMwx9zlMKHgrFUqueg4/+AQCcdjrNr/gkVBk3XofH
qTWR0O8SzfyIiAWN4oeOgQcToQKu/WA0MEVWbabzDT9KhRardkEJmp8kbMP4hS3E
qQZi2/mInQ8FC7GzgOa3rxOStISN2twLEu082TrhBe16ijx0a1VN7Ext3xPUEGM0
DMNlplyE/TI+lNarP460FkylbaJA/nKJVelWFmyC3CA3f00m5fYDXxZTHl8+BPnx
SVi/izSda5zOEHz2yAJq9av/2YxLQogU0rBmWeMUktQPsBAsb/HZL8oxf1zaFu//
m4hYP669k8IOrUZmvY09H75NMtuqjyz7KEa9y5r1aH8NNLrKWhmyBKJeCQJyKvLC
Heyet21GiYMBopPth74F8v8QHBNAWWgQ5BxrwMSq8BZiOfFBz9bROLr+MLTBmvi8
62A9SlJ7DPLWL9JJe1rbZPqPWvDxLQKfPYeYtni6hBJn1BybOD0z7QMd/jPndFlx
8YmK50Js2OzzoOUmfSrEcTr5dBOTMKZ7NGd8r8pWL9qKP/oyAvIYQmWTuKbLrdvB
Y8z/HDyYYs5eTLCaoSNMYK6WsxI74Dt7ktBvreDdilCARlnKn2zZ0gZYeZCxiihR
tlhKi16mvKDnaHfHE3MzRZunpxdpRNnS8WLoLJQujTZyz3BrDotsOKthk7F2nCEp
LOKzYyo8ii2HAQxofDUcsRJM27mN2nMI3tZA4kjg/ZaZjfsmFETPWFLenNT3hEHP
iikE0Pcodaevm/N5EH1iDCiA0ZUbm2lteHJcO5iS3ZXGNlj+++wMfmlYs7jDYkv8
QczWVptaWcBbNtpFnZxi4fuwjAkQP3B1DPKM+sEAJ5t9Ag25S2k8qyftTuZCvwRU
S8rxtlXewyLhZ/7WAFc4KjdRsmoadMxckasyrrOVnsH7UVp9x0Wu2SrupWE7deh9
jBcu/pZhohX4ExNvgu6z5WFZKMQ2IriUCO5mYXN+qPw2jy1KTOKXpaPd3ih+mXUS
9hJGAwrpjbvXC7YpsotJas3UmyU4yZguG7FXS9RDyErw6yqt4f4rYfUqtSKZ1zjw
bdzti+0VK3B8sBiNTFeoZp/aBpAoA9JgGs26qQ0qOVHDC0d5o0czyl5+WQvZ20Ai
+921RwxaNVY1IQNO8pH7RBnM874kekgz9OY+5uXFPVci3cvUHGGzeMCjTF46n9a7
s2GASm7O5ZQkLFKfllJMWTwl7G53WbPHtswqDZi1ci05upuErXll/wLLu+kpDKkN
+ei2JjtuQwzzmj1nJLvGGxTTDlIOKuoarlRC5NbpHZpRnrpHYORvHNOtml4c1UL8
0jgwRA7iKTPiQis6VBmPmyGlewOOwvOgz8/wAaojuNLvq7zyJn+vaLJoyrwnt6S7
R3BSgWfBRXQkjprTsRFflbJufJ06VHhOtXZ+1q4arHVqy51AkMyBrAkPtq3G7A18
GMBqVmfSrRQ5/QppwTdlNCGxgFY6uR75fflk8i/HZDM+53Sjnoa0gJMUjex8Z0cP
VVdsgXDdvbdUxFHRf/mzoLVh9HYA4ogHAQ4KiwmEqJ+gTePjiB5VcQiJb1kihIci
aNBGUzmB2WpXkk8ZSM3XzomS1UFGHDfnYIApjsguE+Uq4SUvMzMWaHZEyJoHIKvF
42a0JDW5Uy4te3I0KPmT5AG2LUWKH5yHJPd7+laIihm2KNO2khViPiUPCuFeuwsL
2QHNhbIMcgtkIBi/WvB+f6YPFxvixnOQYFm5cUkkK4ISJnjqPntqHg1v3k0Hu6yc
sDYgCwnz/QXOeNtqbEAlEBjiGZ4IoG1rSeqlN9qloGJAh+5Ma7sm4g2c0ZYnEH0g
UBQqUMB1lUzuEPoaknBPlRMoW3lUwlb+GfQF1pz7cdPFA+tiEyoAsGStqzlNOuV/
YJ+HV+WsCzsTGnXwn11467+RFiHqmq47KhvdHKgcLO6gDJIblUGRqkDZGujtM84D
YX4PAqv+cx5GwLv2D6k6kHgmFB84KoQbV/ashGeNGg0QGguZ+oqkLViSBSQNAP0W
o0mxi/C5ZtptGkBZb8lz0Idq1SZRVai3O7XQz2HDgVRK/S9EcllwnNGYtbOQay5F
0w3rfg43zXSttZ3kUVJ87XfbDj1wptlQbRvS/e2aYenmrapAtILcHq13vk308hfP
UIsXKdTLpt7/biegAgMWz6V11HTd2AjfrCuLmkYKUbJfE+NPzKjjIznyDP847Zzr
2biGHarEWKDiIs/xh6o85PmxeA9HZ6dC07W3S2wH+CMVO5dmoChFpqvF/cJYQn/Z
cnFj+9jSnxCyyl0UfR3w2+9nhT88bW2AP+PL2SbTfli1aMH4/rvASOaANQdzKr3f
nUpPwRLNQpHKUfXncp5rv6Aa8DT6MNQ2Y3UdqQ8GkBwNcregbHxQ129+RI3ugOt5
w+tJIkH9VutNUijh19Z+f3uHNl5ha0ggSmpWBHHGZe7Y1x4fXk7jlzyqzCbICWUt
dtFpRzQLbtcsTZBSxW8h6CXJ8lVomzMnbZLBYubVSJY5swVUV9Oj1UIx1199ehw4
yN/3KP7uWoeSBUZYYtPu76mTz5E2/rPtWGnwVrfsWWn0o4TFS5+TUjh6cbv7xQVq
8knZ7OU9del/0XOMvK/eQsVmf0Eor+FsI2LSDfWvI18AuCyzJG8ImbDHRtQt2mq3
Udjv1Y+hMSVr3wOdb/6l+9UPNEv+rrKBQF2xBD6EBxlL/t877n4aRxvHxGNQWGXB
Rpj5bnbpgpPTPv6Odv/MYY6AlOsZFkBJHnOR2MN1XgZ3tMGMHRgGXa7h9eCxJIwe
btZ6u8WEN13FM2iBPcGTJ1aZK3vCk5nbQK1yGy4dWTxwSunUsDlreHIsbEE6QOV1
OCM57UMiSjLpMPFVxCdZG+//JKKMklFs5Y5htMh77KuZtxsJuf1htiRLgsuv9T8h
3BWOlxTIlj+OjJ4fpfuT9pkv+Lq3If8oC1R1XAtifgh1KpN596PHWB/eu/zRp+L3
CqLrbJzRjyUi5HEzwvcms08ZZYLpyXP6pCaLfMN/jCrYkxH2ZXPZSL/pW389VYCq
jJjTmn08Ot01f1q08XaqkqIIlQdEZRkb5Jga4tLI+Szr39cTikXs7OpBeIMGOVm+
rzVCqpMy/ITnGUBHY3GtMpVhNlceVR6wO8dQ3AEvUS+XC9aN33vIbFli8pwTnp4J
heZ1BBz4laY4aYbIpijM5Ze9C99zJcXfdkVcittd9lRfq4KbkT7F6dt5ph4dMQNy
5WAiuxCzEMbQ1/q8jRPmwk9IKxOatfywUpm0vUetpXiVkO3SyAI1796AgwKJvXiM
L8mO+pADXYKG3x7LbSeaKiUKUKtpKmS4yvwWxISBkWxc7zsFATdamS5SyOFg9aO1
xV11GLxcXR42/N6UzhMMxkAaC5Hg2pZc+DN/fHElSbt+YaMQhK9NO9+rLTgm7Ypy
7bfs5s6HWFc2sen+G2/doqQgCo+pEpmHhd1vRcMOHGDjW/rqaIdPUA/KMxsCWWJ1
6FixbmwyIIpbWpgcGGsEg9DKrq29asQYn41VfU7Q3zPuYvi9yZWf9vDFeGAnqxda
1WNgr7stzDBObXAH5x99RbQueLi43v8DR3mQ1cZ8py55MIK80ym3IIbMkjAWG1GS
BMk4uDI+A5yb/6uspfXfIf3fCa9Vcp8wR3GuCfPsv0nGDOde/akhJQLQ+XK0pLiP
ZkYH1JCwgDB0jw9qIRvsqBr6NdT8zWt6dFGUhjNJ2wNd5Z3+SnvIGU7tcD2jtMh+
h1VcS2JluncMCSFprX2KjrvnOCJrH5roOnod44AJXJHiBwQM24j5tun+eUnBx8Qt
duDJk/g6ntJKDgtxj4Qv8YTkgH9ZyyQNT4YoJMZDDDJsAqwDEsdl/+mMPkxYmszQ
dnDKC+8uknoXIjZVaxuHg4SVNQVRNJvVJPFw9sr9Mm4yl39RMnpsCykkGnLBj4pd
NtqVCA4JMBJvAiJLthKqqdHrjrWn4eum+MUaG0uiY/6Pssr1hj6tM1LJedK55Ikf
hYPYq8zthBqfnq5GsaL21RcyTxGK7g/4nz9+Dk1B0/iDFEHfbjMWicPorahIpBGB
ExW0OiVss5zq2hisRN+gVurrccyq6w2Fz61C6Az0CRWF5ztQ6K+J8QMBpVwHdArz
y1Np+Xoe/HSeQ6OdHdndFOZdPMgvSjRs9GtPHOJs4CB+UFllEO3Yjq/rh5KRikUV
pCEBd6o+uaG+ykQzcbxIvTncxE1hx4h+BZ48wXoJYm+aWfA7RUTM7qXeAxRtrmiI
gqdu0aKWkWI829IZtTgUvhxNhsn1ONDANSDoXRIOfIkWMtghpiNN3dkK9BNVRhhz
TnxnwYPojs31Lp9d5DRl4oC7/RQ/jvZweYas7Z+l57PrY8H4E7bUxUt9ZdwyYizZ
Mbm+R/Gzo9ctuoRD+MnxPXzmmNJm1jlG89WYCY2O2TIJ27hnG42uyTBNpuXw7aE/
hlJQP3Iz9cJ51CdUAx7TY5pyRU//Wh1mPszeEJ3l/S+RZuLuu/8jjsdchnsRiQ05
zpqM1bBkBFWZm9qXoTNU4f8p14EVQnESj/yrRKFuLrUGQnjoHIwNU6XQRdjjbyZN
13xaTrCqaeDn9Mlq20r5SE0B+3kW++gIaBGTEE1Lk5koY1lckQ928Xi0aa2eV+/w
w6Kkab84F9zSB580a4k1IjuQ9TjyjO4ZIg6AjAlNjXWt/NICK3w+v6cREYr1mbVO
XcJGN+WhbHaMmlj3zAbghNh4Emsc04jS/TDGNdTlvaPG73tgV9MHanZWfG6rPqgx
FV6Gj6scj775pAO1WPeps0IH0ij2Om7EZBKoBXBDKL2S6m4XBMOuZbnOTjTzpRzc
thNo1F7Ej3SK5TqnYiKhIg1+u/vsCPyQxEYIAp45YELeuDT1cJZQM57DMfrszJBg
btJg6NJJ8Vom/0uwvpdbPnNut7l8xAFvBam8c3QXGZmlExKryVs2ISBqLB6OreEb
s/MvNQ62c2xaG7mACBuCI0UjMzwaZo4mMvf5XsDu0/7g/bDNv00qLtB/Zae8+DT8
imYZT6DeFaBjj7kacmExL29aMhcb56iDnNrZTkotPqfmLrsuStrMq3yuVBaHLVal
EGV4ePoEOK72Z6vdpuQRlccMJqjuP2cDPdIvge/tUZCJDMgOdewlXg9aSLscx+tV
dMKcmHsRgPHQF33VMAreyGV95RiBejDohKjCDKcH4xA7gf4ef5t2RhHtxJNvhXsJ
iOZ6+r+rxkVqKJBS6BMzoMeqDmCtv8p0jabB3jyZRQecSb5zT2zZGAl/0fJ8t0TC
qS1sKkFu/8ASW0B+ZNbDJDL0DVAI+3LjomnigHLb/w50ZYW4oHSmwhGZp1jQss8R
qPdLecQmt92wa3USjAecvzA5tJxje246fc7JX4GT+qh9+sSQi6Dw/uqNCg8XNOwX
93dj2/ytk9DtyrveAt53AIJ1co842arS6hWpr6MoyYdGPClMSekA25//SXf/xxjk
rGbEx/1WF1Zvye3TgEpr2KwuwKSykfQYKO9fq2mkPZVqI3OsSMM5L0NDxifCrv2k
YLkAJ1G7qBFRr/BePzIJM2FQeE2Jdj01yXV+eyuZ5Tje5xKh3UV5UIEzw8E8tPiM
8KTOEmKqVIAg5cMoIs+bPnS7ZCTOalCxpN5nbY/OROZlmU9KbZ09RCXY/0xv7X8C
NrorYhtumSvRk+i6WvrHOHP4+e3/Tf7j5Tw9Cuasw7r3q2PK1eCLOjO+mVDs6+KT
R6goJgSSbL8watT90tB4/wHhvDQPaRYCAgc3iYQqJhMIlyiLi+WErZ4xCVmKsQiA
XmBgUskOBfmwEoQr078s1HUzVBVaMLkGSQd3u3OTjWJBRvcsaGqfc2OFzTnN39rV
Mf/AKopmEG2j6lacZ3wlXXwsBcIl+VGfd99OygA2C5mDwnTONURZByByj+bLNdVc
nnKAf0deMBV36HeecAWsVWpIEXJHclArSHC/vxU2IbUgXQ4IwZgr8hwzYiCp4Ewe
+JmCyJNoYsicqueKm94jSGKq7UsvUBBb+HjgCPsmrV/BFnOzG74QQ9cw6B68weu/
Wu0EL53kn0OcnZm+KxAFeE0Ln7H7PgWbm5ukQxoxWegGnxj1aMJXNusSf/Hgf+Cp
VUC/YlimBYNWnAtES8+q1p9NIGWHdi0V9aTxTIqXGrkk7vdxV/chUdEvlroaJH/N
KBXRQE512WsnxnOQ24X2o1H2n0mIRORHbFZ+KbaZzmXKGWst3WQFhMbTXVqAyumX
oyEpTlhEH+a2VrqgaxDHy4x55AfSCTUZQjCHNNeJKDWC4VnWKuKXZJybk/+mMoif
6e0UBQFQ9K0iG1wiLn53Lnnrdow+H5egJGDxUrIte0616SKc6Y0PAXmBBa0AXNVe
3d6soOsLyQWGlIMZqijEpAqWoLBZROLWewuHU/HfK4MpIjQY2l9UK55leyF2k76H
LYO6pVUb6Ko85noesvrs7aZgDC+4I1AtRWzbbkaIxa8sk6ldQtS7PnPMODqSb11L
6xjBPAk4z60LRbgHHmk/FpturMDdgG4k1QdhNtJnF4d29Nh+knkPDcR03MeRLMuF
sQ8VyuiCGJTtvY6P1au8+scsORdlF/Np0fmMQaHremISbL/lBa0pxxc0NKPg+7mz
VclxGsk6pMewpjZJkbR3Dcd99D4VBEZh0id6AoVVpbA3w51Iv1sZkGCcD7m7+RuN
uOLm698uDWAO8EkrvgiIcEcuOwMtImwh2X8TktE4MayIvRc4X7GdPbMOO9BYv3dI
74IXykcq5fMRbIfMOMxqkOSoD4aIpAuuNtO0tKnTOWwiHxZnwWfP4IeYnlsgT1nf
eGGwi1xXg1OMTaVQJJD+M5Ro3AlUhwpeb+g7H9M6W6c193LTMr5idbrSZBMnoh+B
+ozbJNkzyxK13ac+fBrvZL8e5TjDgbVjh/b7Y4omMA9SA9NViM7IHsn8UCfN2Z7M
GQP3D4nBGlxn6BUCmvSOhv6NIGsNM0U4BdaZg9G1iTw4tg8AUb1SHTwdFGqKJ2Tl
NWk0DCtmao5rdnbLPygKQibcePmP0eU/5B1Dr3z3RL6s9+TPTu0ZCPm4l5YQjwMT
8HSxM4IdPla272u0h+qoAX+swkl4Rkqs6qG0F++UklS67Z5ztPnZH7x0YbkQdSW+
cPqOgG2Hae+v4IY0AxJhFqdQUsCBYMYc2vDOCSA+aQlj5Wj0j4V3YKPyr0kc5wZB
+yGL38onag0fDSHd+zhXQwstImcggvWjo9K+gxOGOOl8sLnRe1RFq8QFbt9gK4kO
W3x4mI3kvJ+1rMMZ43tMLTf7WxRLFJMlihGaxjIQFlQORq1VzqFkSQwXylrN/r+/
8ptDeldaX32j/06vjZVOnczPzorAWah8oCrN8iFHW5e8b50UKHXUjYFpC/fCwIzd
mas71+6urXjjTR4ngaV4B9suiUQTP6U2EtXHZRcBy1dgz8qn3M0N1BB/wvx7EInA
JJ3KsL8AHiRvoqehrMjr4HWURi7QfFTnsXpVAC0YnI605KGX6d+wxRoZOPdF5eRP
PUqvbkNwm3X2jnIZug/e0atJylXo9hKpp1rcca9Mjs2hMe6QR+xE52c9Iz1XQAY+
6r+6NtA3qa3FaJGp8yeQvEUmuJQARmXfFRbAStJAs4y9+LM/2ZYrVIZLXIEwQGZQ
x+S9FlorhdDJCwBI+gTZC6nm1JsVgx+ZBqWv7w4KvSstkuMrnuEu5Y66Q7F6uv7y
2Ph+OsIv/Q/b9p6Zlv+/RZWFiiFu4KNmPgFYsbirxOaD0GGx1DGZDAn58bEZpf97
/HUKbbRaCeLZpsXHWPTlLISHyEQdxy+eUituB1l2MOCwv3pOwe4uhHy9B0KbYBIu
uyB3+aF6S7eUXhewpyQF28ksGJopzz8dyaanUg8RiKu+S7hWG09sQ47dYQ+qqQ+D
7StQ1zMXNkAS3VURqfkx529eJs7g9MaOnpjG8uIUESo7PSqsMT1+8EGm/nxOwuej
Fcec7Zy4gXYVSAr7uvrVm8zXkDkoqbCskZt10TkKwaJSiFVA8WSKEcvROkiesuCe
/5PqxogjXNfbdLEctwXZaUxVL7lHCtW58R+JQUr+ATwjo9N9R7urRTAFoyN5GB9C
UsnZ+w2x7YUFn6/OBKXhJeF/m2a/lKXeFnwdCj63hXUslGOgM7nmfNM93uZf8gYV
BJpY6eO23VQcp9GhwQ0dIT5Il5bd1WALuVQYutqGlHx6HwmlU3UlTuwFUhx8V/yn
NZ0RoknDYOuu9FgVJcVox9dx2I6xfrwv/BEkKqAvy97i74GONqHmmYj67G7QQy1j
kzvmIPuWpzWkTNmRXMTp5BR3+/1x8TJC35xeeWlc86nzaZvmi61pwtvFm9kZMtkP
9GFol+rzShyP5TaGVZHTu/ytLnvuvik0VaLM/Ry9ABURSvW5lo0QDp1xlJDVr4un
Auxh9HIlFMPZ+X/VacedDYF0ZPc50s4T8WRdSAyCRM/3+UOE0jqdiIE3OAhQRHYU
vwI4Q6x2WklQnfR4zyeqs43T/ad3qPHEH9XCY4PYDZUred3dOHXI99PjpkBb7zqZ
XvizmaAFKk30xgyGrVnx+wqvF1/dYRrKr2xitkPFvTeYfHA1ShMTUk4y3MPDMfF3
+tN02kUUwclaYaLQ+sGx+nEKq2xfVUKCYG+TcdsIWZ1j4n1KeSmwZzOuxxROTgaw
qrmD3OSo0nx43VIk9kCeIokZ4pzJCpxGzDyLX7UcsKQ9KRSgr/Gltl/48ytE2ItD
08D1IGYAY+Xd4uF8dFjhpsKK7vAB9XRSduyqJi9lpyNq+MYmVorCY8vXAatQJZxx
RzE7g0lTwONyKshqHp4LyrUHLpTj42hw2T2go0pP4J00viFgSbJw5VDzftKrDBLx
qkGm7H1BbAH6pY8NnWW+1iZxLTncHDEGnKdjvZ4ASldC1JVVOK+/VXiqQ8RZcoS8
47XxuJw8DkvvcGllS37SdOEnECxD0oULkY0QM7BhevutmbthO8F6QRj1h8zfAuco
zzfyDdOe/be+/j5pLt7smdiOo2OEinUYo7cdkkbQt0JaAbluZRyxa0VsubcDm4R1
uFcJwCd5pQrjYKtEXwHfxdv2gJnm0ljW7deD+wVAB4tzTlP1XfGXftjvRQJ7qxh0
3VD8vLybVLeXTygpnD0gRAIiOKkeqF3T6gdCinJc9aRAR+juL0q/+GlCfigExbHw
/0F7E+WyJFiLzDlnRije54oZk24HsTWeRA2H/RRcSnJ4NEJaDQRLTpnenHSRCb2e
y9t03qIiMVfU2gWs/0GxIDMZz8WemY0vIbZD/pdI5KmXpcZZBBpqWM8d9PiFmoW6
ya1cB5kopCEKAzD5TLaghP/A9D5PDBmOPj2ZoqexAz2ql/PU7VRBFou+oxCkU/A8
Ygg9cohPjoZfGRcxu7nMJjiPu8tF9X5+QoX6jUoYyGvSapwNyTppa0yCw8fSPZ/x
3TswfqykB7cBUN+vO5qM0NUVyIINVukYTsAiABxRF6NdRyM75lOXThq60oUhQlMl
tQ3TMOSXaioKrQQJMPeeXHVLQ3rGyay/71kKt4gA7AYaDkLo2s7NPfc2O8IWu9nd
cG64MvmQcLRAs8pZD+Ms/lZ0oYKjHuBrC0XXyn3gLRJqRCVjEsXN6bkDXpGEA57s
dRl45Ehxv0a6FGboM0tPAac3HvLCfBX2Dpp1NcaswmDG2lL+1wjrt5myXYjRWqME
m9axdIAk1XPQm96MZ4vBef0M6NcwcE2Rz79E9S4RGAmbCB34lF5hWN2M45li9W65
aOIIVWQw2b+0iwD9pMsuWA6V8hwtTLf0UT18Ej8I3UMHRgiOMI2dpGIPWXX4e5E9
RxnCq/e11KucIPYMCI655ELvkzpSp4OHD/bsgVWPwm8xJ9ifCA93P6X9bAqagkJe
oT9FsvPTRqve5flIj0Q5QuaHM3gJSFkgc8XLZR4Oxlgk7x9YTDbXpz7uu6vPUycs
HWnlqZ2psnEL+OuyGlyWBN7s2kncL7zK8c5TlZl244gx951Wo0cYK+HqtC9CHaWr
xFXaAeFmOOaWYKJjfXAA/7SWTTZp9HpE99AXd0VYryCel8Sd9bub00kMBKsHgRyn
/oT2k4PYCPgudgxDmcHqIXX+I+gjLVq2xOI6DSqVzQaRVNapeBYsPZ8ezb7r1NuL
gTIqhe5Anl06lbTHucrx07tPWMFcXlqX0nQM/napQL1SR44LdISpaaJ/3pSf864t
wtTJvrBNw93+j2F1JyXELG0d9CI/5i4Iptg63GRfVo9Wv9BGYJlp1z5df28Sj3/V
FVo35kmUARUNznlIfL9rYQb/aZ5xgXDHX4DW/47yA5U73MOIuufI0hIqMS+PNFU9
UWZ0Lhlg0xr7uEsZdcDF8C8WFWNm6pVUBBR5M4m2QeOW9DOjlRuXYE/P+3/DxBVR
hUKSp+DnNSIcDOUVRogdYf6MVWjHEW/W5eUZGtNSD6o0YYX/JRmIrvKlyIFl0iPR
FtYR9YjYAZATimeFgxJ+Dr/AUG/e6LskstZmZIRwrldTC0HksJalcQHE38JykBA4
v3JEK79scYKax6lF0Rz6OG5FJia6wDKu3EEYxIgTLnh50OyzaqVbnjyOBC3esyOG
MXeMWTZ6TQLSIM2EPJyDiqTEIjanETwnI+kHJvuM7fbHFoZ8j0EwwHmMA9ycoz2K
GOzdhAIz4In1p04FANfeuMtL+iyiP6dp94hGhhSYJln/mumWvVpIfflRfA0VXg1d
X8bt8GtXZJ2KrWTo4zJi3uxDvYItnaGMHGs8RX5SBWY/yMFtkHQj8ZQZ2wiGcHWZ
wAsHziBFXsEAoHWJZ5sQXYen5QsQNJpP0mEBcpwN8FU/5G+MPZECgT02kYAffkyZ
XzFt1Iu128APw31/HhEyorCHBoSLGB3B1y06UPliXIuhUOBA0fAop7gzGczNP7oH
P0pRQzGj86pbiE6cSaXlaCdWvblcYuZXBNIVN9MuVOpFQLxmG55WliCYfCdBpZ8K
U1d06OXFtkcNVwynwHt5xmE89JAzAlXqgNHplbOMs7Xmtj+8ruS9PrXOzglhQ34Z
lYEZkUOYuSs9hecQaHbBvsmmnM0/96rliNyYOoyx6rd6QfIwShXFCexFc90lKPYS
ov/YvNXSafOUaL8tkrFWqHrIii+vrx9MuafLhK0/T36rPL5KNGrXwbzAmTvTQF73
v7ujBa04CdC9s5C8PF793x++lPEo1S7LxUR0MDq/bvCAzyXgmDs78jFkUuFmCnCY
DjjBGs2fLu1S3B6k8VuNmqQvhD31QSMFP2khJIuIsQa1it3V1l6M3HFRjnhcusiN
VtmzkyCqD/PxCpK51kCFmpLgSmqTdmpPQ+EszmtBIPYxMY2AZM1wp/nBYpCjcFrf
1cTRdPaTJ/rw7HPXw/O9PST1M8Ko3OzCe5GmWd7UW+B6/fEoYAIaRnTJPLMmIBDX
guffTlzdjcRicr81WTU4fG2D+8lypaZwsQvBIdkSQ2KlDDYygjQc0u8lOPZ3yBXC
0Iliocr/plIZsvEcnEweSFeeyNcsToNiuZQ/VdWahVE=
`pragma protect end_protected
