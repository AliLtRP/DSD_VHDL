// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bsf+FpHz1IRCBl1m+Qz5JQ9AhGtFhjMz032czlq8ZN3Vjh6psSoPS+E5mlAHtWNz
wy0koRn83Rnnojqzax9DTBXpwdCm4rh20PMzvzbhnuwXjGTXM8+gTnK7gRm+baIF
KIIhu8rIdacht6SFSIhuWliJuqUC062xo32Ix60zx24=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37840)
KQowJIHBZ1KRDVS6qUeAZltW2TTKcDKJZTpLXajVY0dzCaa6PvzZs83ThW/zWmR8
SGJ1LKOdY/y7NLhv+13ZpC5mbhNZWGO8mT1Z6I2MWg4kcnG0WPc+4QkoQSc/Ukqi
cgvRWg3uFM2paCLh+93Lb3DqVOTTATNK4R4TkW5WxHnV6o8UVbsCw315xSD4gJQa
Dr4lYQ+JyCCl+9f4qjeK5v6P1LGhijipCBo7H0bYlZm1zDLH3JugyhUUvFg3MYqS
D40mxKE0pbyJItRueAufo+EGOqGLRPrQMBYhKG/ZOcYcvjOXY2Jr+9Kgt+YVM99g
Ia42CpEO9wmmx9DnoFSzyjLrR9NSN50q3EEr8p7wWQ77InVyv2OIuaLI03dvsx1O
wUhwfiBbdu+Izg1jgj+1ytWrpaLTezCIcXr43kfFDoRoGt4pJCg8AOJ5TInHh0iq
mI4YTOBRqoLKJWyCo9cySxQOpc/u92ALI/L81nqjDKNwyY++JCsylrLw7ij6/79G
mZ2Q0cyGf8q+92EIfxc5+ICXfGz2b+2iIDseFKTMl1+RWfL5hJyEZ8xD5Ro3WIpL
ICtRmEkajPjCO9lHwwFz+e4RyeAHNBCXTBEMMgX9Qj+/ywpEVEiGFVk6g6xOkZpK
s3Ri+4TZeXvkuv3xoWvYbbwXuCr09+D2nwGaq1nrjQczJNQgJTh171XnMC3XDfda
gErFVIqvYkB9nenDc+92TJhsOxuvLOb7AaSHjUVTTcJzPnCmtuRmMLr8vzrC8lTc
bJ6/QL4xVGEW+9RS/JDej1rxOuh0QjPb8mRI4ZD6GCh7HDfGmYCPLzL6U3w8VxH/
fDsQnJa4YJWbaAGT+8t2HE3Hc75l4Egc8b8MidC/qKBcjFdWSGB42JXie2hUTTqK
VqzjL+MJap2LHzF6+fCTaTSENOPEmBbIIO5NSTVqX4DvsgwxGhPfrXFANpm7hC6o
tlcS5Ds/5T5CNl2PdkqXFCbrdLcj/hnUkSWLdbMR1JDv2VQ/e5JPRAef3QNcIDGb
JlKG4tSaGKtKAaHUVwh/uRaUNmZDChs7xge2AOQjsjLs77rHjISAmNZi9g7DXLPR
D9l9HpsCPa702X3fr87tx5Xw2rAQoQJGUsJz6NKA79Km8/iNpqgf8KP6qNkK8kuA
IbQPyXf/Y4Rj8DuqNgD+aSOnWZ4sCH9oOkse4xYk+IhDVu11Duxidqo2mCPwOlIi
wkU+JSqd7ID6/TsX0+69wqkf3kjQDSAKdo3OQxttfTm+cZGP3PZDxvIUfQS+EjMz
HRljMNzqtS0DNEY6KY8IttKnSfhyvl/3tRbMeIEDOlF94Hm2otdmA5MyIcPtbBVB
sTYgOPSNOtNybRmNcdm4A4UUMHTpIYqJI4J4EEvHpheNUT/jhzblABeGTeU0YVxm
D8lwO5JPAkpI2j7PGY4xnoO/bCnn/P0uBkimCGqaeXhpdoqCptstUKwnLU/zFjPq
9GUkt85Y18wRxO3N/mxm4+Noba5JE3TcRxWYHQh5a9eh1vGeT1L3ZYdfyLK6H4Ke
Bhp8HnrjIRY8H6dqTCvw5Ztk7/ynJNR5kl5oMMr5xT9aiks/fwwR9O1oSdp5xFsI
I/Sgseqy3R9DRLfzvZCPrA7UTzUE0hwmR1z/TUDR0AbGiABzFQxedbwIDYXMWx2j
cNzy2Wj7n+dL2dy4ggy5NooSlwA6CFhxarZiuhCoWRzhUGedZi0MaTWC7tOdwv8x
Vawrgnf4k+2fk8I0j5SAT/Dw3ll7rDqH7QfVPFaLFMNUwVyP8rcEMFXWRy5JDTC7
uwguT6MCnZawuwg1dqxo9rl0PKzQQAdQ84fJ7AodO2wlLXCXgqlIfEC3UBTRSfy2
0aoFpTu9CAEXFcV90tW8MndlKMWIT5KU9gjkVuwOtwqaDBAhjQpgymXhCd81R27D
EKR7oTujHjbka8kY6/Ws73xGJ7qgSyw0yKI5fQ2vvnZhvNo1Slcn70Ewu4eWQ0fa
cMgBCiwHChJZRr2onX3gggFl5VAw3HKquYf2slZWOHIafhxN5qdARluX75eWgj44
fyUG6nOeYSme0iu0O2SBuoSU/zE5VMmcUKPGZZaPwNyHyn0JRppt8NwN/NG6jZp1
tJdTIIudQNUTUHLxV5WoaUUrHOpk4FtriAYUn0qrabkGYJ35EGsJRNF427WDpLi3
ijz2POITSx1sWMMUPWsdbHa881EVn8VrVquhUhFvMX45Ind59kVLCuTgvTbAwE0e
cWmcuvgQhMHTPfzPUdZzxYC5bmMlqTX5+RPA4SuBnNKYtSPnzcuuKlil5WuQX1Rr
Vp0qRRjw7gy+trUY41HQCs99H8MUo5eFjQgt1rwX0uEjiZoBMijSJ5l1qwvBhy1r
+CXaUvBlawNnHC0XHT1/pirBDcl5obDUvx6VnYKMcDAGeTtlsB5p8ch4k5v5GWHH
5/ExI0GG0efwEnB9TL2yxu6pylV3KacSKCaiT6xpqkob9+uJRkBGzHOoFkVJF1Uy
ScU5+mBLTCqkFDDWdeJbT68pOSptMGA1DYJ0aGi5RUIVnDvf8PBztpl2WRpObgzW
TtL4ho+RNH07iOyzpdaQKLgDz9Ex4oABds2YcoJ7MzEN1Tnyb/kFCHy+J393HlUx
DQuuGnZRpZ4HzNE643vY9xAmJ2oaoHTv/PwskzAT5cGGde6InLedLD5Ed+NjrJcW
4pEhF8ap1c2dSixlRGC3EnXn5pYNN0jWSvgHUg2aQqoF8oGgh5OskZWxpSPxxYQJ
LvQzBpiiNzOrEwxHiWWRBteBOyXDdCUuPokJBCyjlqhTlgcjMLSGx3CqVu7/lDss
Cf0QKGYViTIx0eMM8ycqbTPlUZLiv85vLfea/zjDZQHh8kv4vlsKuDQfMlqi5Zxy
fpQwIUo3z9YR/oS9j5Iu9ea78SklyHgTt+6+Oi4CEr9H/e/2//vCS729UdvkcVxr
eSapHeh0vaezKy0J5yxiu2Frt8jgLlvFapdH+qh7fZNilBMA32zi/bBaXJsk7wT/
ToMwfV9VGG4vPGWxSmo2ZiD7DFGUY4fFxB7be4vJsVP4mM8CIpf7y/of4Wq5rsZ5
+8dVCLiBFc/kRPkFWSqdBxTwSdMyoiAbdWmiex/6zlrAoYFgavuimbPMZuTOFdj6
1pJY59xXYuxVGp4L9hljDfIOU7xy7iX6J0GoqYTA3DXhwHm52NJ0JYO+fSqiThZM
pXr/zMKfav7Sr9GpDx0SrftIYC3J4GqW1WcPYcMCJJjnCPKhyhwHRNIaGBw7wGe8
vrwwMYoenT0+Z8AakfUAs8463oH+3QWOhOldxpwkF0TfPWpQAV6JoNqzYWtee2f0
nnKHzT5x+YJOynp3juO99OJhuSW4k4CxGlqDRI8gvl6CG/IDXfAEGeHaLum1D0aL
Yg0aiILSP0mF/EUAYE8FITslmLstw443viB4nJigDk0ziNqIkrODX3dfNuDZMRQN
z5+SHscv2TPySg5Kxx/Nv4qFw+YZEfL82ijn0Iy2UKs+I2MtFl/joJNgQaawyblu
ohDpuek1++qU/LXHlvuT/GRjUGTkT4hENUlrmYnMBJzEeAYPnt7hA635gb6e9qgB
eQFe9/gihxsgDrBDjEkKiYR1wPROO7DaU1cVu4USz9hPmWx8D8bya8Ng3mhIn02P
DlR+d73wjnYgpFSQtCvM5xPHDn2iht0NJmBl44CqK/uKKSQAt3ZQCvWxmL3g21xD
jcQeHSt+IYvyd+rYxMrC+Orr8OYZYIOraI4dZ3j+w15pLveK9/H94rcJuAszxAZH
msCXE3+1znhp04c3LKRa6A7A/B2LH/7mINrVq+m4kRp38N+gEjf6vr2ivcScxKkf
K7PIDE+DdrtBWrO2zZ89ZElyfac2jZvuRGG5Hv3PBO/zzsYaJcozfOWxubxidu4G
wXsadIjpqINVk5sFuJ97oaV9kAT+nLo7V9SkwPFKNglAVjNqrzTHaTFJnoOmJzos
tlbO9Z1ZQUAcLTN3M+3EDm4+k4+VtrxjhiROqC4r3xGXzdAFGKOx1gSbvAQMFBqO
Bwkz+F5u6rY7d5wHr4lXyVsY8HpnmDNi2j2UiHtIblMoVOaj63C8qcXNIdIZqQRJ
JDo/8jqhddT4GsOSxL31NZgrTLitWWWQ0Aw/y//yC8IJAmdk5L7MpwT50dY2hJHW
Y7i4qRaA9NVDyjbStSueUqjCtZJfSKgLOu9s0nLQb1OMB9nIn7rZoxm3RVtuASbI
HpbCOicIbrngTQ+Ib9dXHEw1QZyIHAw1+Cm9wyY3ZhEvwlTiNYVaRD+z9wuUOUjd
dv28JW7aSqSkT9o35Nci40M91kwa7/VANNFIihx81WI9nkmsXb4bdz+08xqf5fNj
w8Xc9qODwbwJptnBZzYgHVHkITaCPjhcPSmx0ddIAeQJR8fO2qsTritSppvFn3Hw
Clyeu/DnFXimbPRv2ezVOiPXTgRPD7fjcS+vSA+Dv8LRFCOnGNsFYCy2dtPKfQMm
XeANy0GdZMnMPQQ1w2LWeWE1IPe3lGbT9yk3en9QdGCpaG4MOqcJ1xMZERndt+eN
kH03c5BTulK4mBxkX34QmhaN3+Zt1gdiZ3FTTTojEWonaay2GBWsumMeE6Em5s+b
9TNMP1WbM2Aok6aKtvKCU1WGh1EAlQU9WykNMoimnPoZvoFHjUnroIG43p1VWH15
e+eJ3I/uKWXbs97a11OJFGP5ahmC5Sgj+AT+FBZxmcufK6QHb+utJJdI2WXFsQWA
7QKQzXuDvEBgxrzolt17Wlms1ojgukSo+pZ3LNgMBJ9BQjc6/4edfTQs8Ir+zyDX
qT6WTHXHb5tTVh7zybSw+nvGPtLsGSfAKwVFWvFjET6oSWlGx60ccbHroBUoDsem
kOARd0/zqwOrgFBb44XVEyNVYX4QhW9PdqAq5lx0weSJNhKVvy2bcQEptcKm8wPM
pQ/74QopzHBMMOSQeyczBV6u5ZhCzZftE/URyBScwJzjBSj13aIX851egm2dUKmn
OhltvXwUnA8Tltivd6DvBYKtlB81QnSSDS5czupcWMFfvPMld7wjwziZuvchCmoQ
TqNSBnSJJxQ40Vi73pxRzOtxjRPObjWk7FjK5EaHtin6buRg/pd70e9+prSV2oYM
JaKHVFkoyQX2K4fu/cZx8leDGvFXvtzkz9stvqIAICX1jU5tshT+u8Nw1V+GIXAw
ZdM/AbX9p2es2BhgZ+SgCxp10XcmCXrr+WajsMSIzC+K+G4F6PkVyrVqejms2tgT
LRfEtTzcQHyZSveFuLnV0iSiX5uTtMlqvNex95Q7RLlIukXBxITpQbdcIo90Toct
Mvfa00bcp5HBz/x4P3JdtNTYTB+QzEFkk/IFEOVJ5Azudt0JlxbUKGSRx4afr3ML
SOU2wz90qyhwQNQbLxBMyap60zgVIG2m7xUoR0BoZ03albO6jvPZn4HQg6ctI4gN
ytJhic8aY1BLqDa/5v0zypQQoq997PcEL2eiTZLhuoXIOjHb1nR3U2yVb7NoNnTp
vmBifAoTaBRdXkyRCFrlTfTeiwVLWTZJYzWKRrWiGdqXc516tpedwB0SLogAw6jZ
w5OWnt0mFWwhYqP/DsYyDgWpNmYwMQS0kKSgMETZM3eYgb6M3xLZByDtDU1Sm547
AZ5l5b0QBNR3o4KjN9KM5j1LY9H9X8BEBCwBQFcx0T0cwW+79tu2/XtWc6P86wnv
pKNL1b6W2BOuVUh7Gz9/ynfU0dlkPQMR6ej7rncBEuRFxll0VAkrGq8hXGnKkpkX
Tc5KYcibcrYJyTvanFAB3n1KOgdO0N2H/5qQXdNwsRrGnbcTnRvu4udwYeImdSVv
RzvOHrg7FHgXn8LT26iFYR/meq+Ycxf2fyAdrBMiaqn3O0lMwOj/N8QxZB3ASH0C
KK1Nw7asU9cS6Gssa63Q7QVic1k0YONcvaxYFeWGXr01Gw8VyY1HgVriHCJoxt4y
h16NaUZ+VMyJAU5qRW76/U0TMEfW8dbH3OUEXOpw0Jc2WXCLagKp2daLDTuVyKaA
XH0AO3VHXVM1TohNyaJc4uVUyb+ShpmBZLlN0BwenRXp7dPVAdoEtD5Pb8JCBqqa
tz/BttvFjcDLrD2sr/SQFI6vpo0Cwsm1ZUpKvsuMIUGQVjHl0w3pUXW70mQ4fTQ7
JAjM1bSJHx+ap3aMBKilUbBabmYQa9EUaXwyP5W64s5SWNXb4BgxbW0s+Kv1aWMQ
Wef9/lr6nQOY2BkZUZiBXsdNVw4WdmrUxB8hVoCqZU1FaA2UwGIuTPlqoXQU8E64
gSdb7jzdHdzXBao8C4GRZljVyk4lLthW6efDKj93NclyedvSCVBuVGjf3yjFrkd8
QHHqagkHwbB2pmjxLx+2ACJUeUdhQMfu971BEci8Y74CZByogLX2yo8vfEb8nKK/
0F3ZktnQvPvdJjdcB+Q9YgMZD8Avx7/dpIK8eNDYzwXBdUtlHUulhZmCCiLXPyHZ
4ltPDBvFYRv6Z/T6Kfu7gcIh8SpFPBLr4dKet5O3UMLifOXu9QJ2RJZVF+tX5G7v
CgDzt9PX193hGZ3IeKMKi1T8bwkv2fu8IZ/c49SNHB7aiRHgmyfJr1lu051XFVPJ
XelC2XciFuy+7h6QEcQ2Gu9l72/S1jr6QE/xkZStYqqOV1OC4IbUKd8E8jEAhHfi
NdS2+gc4PLc69g6t5Dog5DeS8roNA5pJiqDf3jQ4r7HOx3NomB8Hn2o9JLoovr+e
2Zz59eBn8VXoquK3CIvJkr6YMANsoeJOVg0hquyOlww3biDb/yjgGYWG4Bkb3no0
onHeCJEgJOGQoceI1lWLqFfkwzNCrPTUF5jqMVeEvD/jMF1JBJf3TnPX4HiGYs9V
/IBu3rOmQ4AAduE6yfsrJJQ+quIjdoyi+5AZgkl7LHA57abs3jopCFaHoQKksZ/i
Syy7nsY5YgTNepOCCy/DZ5JSAkpS48L1ALglO/2utO7RHYwlWQLpZbKciwwuY2Mq
ilr0+HlRCwRawrYWAMmFk2b26l5SP+EDcVLVit+d2k8QFzKK3n1mi69rt/vw11nO
Ita816YvKlQg49B+UWH6DMuNmghxj9sAWCPJegD2XYpPPnqYUrfkeskWrYsLtt+f
rEL0kh2or5Y1/w7BztaPgCrxoHLxDzi5M4kOaSmGREafJ3PsqWevBIoZ8nk5FzWL
FUmOSM9ZTWjtaUieh67jCZhM3zu52776SggaKAf7ycY6cwE7hMvaHXBCvCKhUycl
Wy+CHXVvYyc71cGcAPzPSlNbCxdNYcRoNvFT4hCDOVIXDANGLf5+JvDtRNUb5cze
WljKuryzyEQJxxiNDm0saXpe12tkypmFXNpmG6GsvBBkGeL7LKHKtEw6H57kpBlm
5F8zQ+j4k7QpVwZWZ1OXEDERg1oxPzoekDATPFa5YMcYtmEfYWbefGhn0zlR11X2
QLGfxlHsM2oe8FQbrgO09tXQ4qlCNbafutUkPsDUEWQlvAxAF31bcai0AsKUw4jE
APaAuQ8TWQs8RyWaIK+YDVWaBeu++bM0ZfMjiISXPPN3UdK5PxtIuTIwKdQ/HGrP
Xa2WrWWIFiTAguR7IsT4Ufhp1qFw+gQkOw0e7FPoMnmU8q+9F9ZBjgNM4kcQHuxy
N7XTMXpzYkpNamuwzv3t9OKTGT8rk3bV2dxWN9FXZ3aLc0pcD3mka9iEMyN1uJua
32+S5ZD+qiCEzizOzhaIOa1v+AIEOg8b/R080oSS/QGg51oDNvkPqXuo67kxvWyU
v3gGVCDmBwYVq6gfN2E9/VFK4lWkW3ibEdh+Y//+O9CQwF6p5tk1jIZB2oyMmmME
Zpn3de/pKbgq6Tf/1hlvuQfKbdrAVKnw/m6gGYceHV1tuGAMStHci7GaRMTVAiHy
yFwn8oeUE90Tsu6Rk8S+aoUo3sUKdp2feD+tS/9y8jp9T+t3RAK3v4u6XUnaP16k
AFMrxzptEy95a/KYxekJSP+/xUzSuT0XiadsW7X1AyOqFyNfai/Gn1EWa6dCf5Nc
A+tnc0sOb/S4WRx78YbSMkdqL6z9llHuZEdxJ+LzGcdib0zWoauh/79xMUiHdZhy
6URgfpa+HpkBUIbULIzzK6R+n5Pyj02QjdhZTFGz9ASnvIg7bkHibbvzjp7hSkIq
gB12rwe8x2xZpfBgJU3zoODjp4f27ReyAtvXcPF7Xf95/hfmXorvgDNeZyGwRt1B
4II/vX8/Fn0Bu0mL8SqhzsJKO0ZY/zUsBOeM6NieuIJSTYrDQKly5LkS4maV2Uoj
NOzdl+0OeeBX6sLoM+AypEOE0BoFQtURwVpDtot4orklk5qslxoWsQOsyhyRyVfV
CcIPCn4Z2cbAs8hZVy5mnJcYu9qY2BHGAgHGrtTgzPz3CEi7CuA0RC9PLchOIBNC
6MVfKnLS8FrcDaEYMFz/UuZIHcwAPktQGhct7b12l8DPGfCuFPd0T99Mu3XonOS9
C4aW3YQWge8eHeNtHzvlD77GnRN1PfN60f7MSFV1cclI2cctYFnyyGNSo4AMiPC9
ApDNhukwFR5slqzVyefPLbepb0bB6JJbXAKDz57ate8KuFy67GnraVDY5jiDk3x5
0SuJfEPLzAX5jpuJojpjfdnb3BG3CGqQCqXu7t2/8ivRWt0yMTmAAIybsJRI5qz1
ySoI3/4UzCSdDAZzarvFvsMMoVUUxrcSpJ1bP5oksfn4hivGo5Pj1s3hEYgBymfi
dxKro7kr4yc5M2yy6mjgsoeN77kdm/owjl4ZkEKiDpFH6rnf3VLzd7odAnuLlNKo
VVwdsEg74WnyCpqcY+aAVAZc/6pbgB4yjM1986gvudq+3MwcW6YC1sZPi2kvsaiS
f2Vm9W9xMIGId/djeLxTYh/V0iBvPu0nwbbUJTT9J8u/r2PfhNL5Vxrbj/jH1dL3
cDUnyMFYjWK8ViC8kYdLxrvT3T+9KJkmCo3D/feaStsEuT+qQ2D6Nye3JMiuw2eb
kSUE0VxOzrNZNyY/WwW9EPIDX1cFIsG4q3V/dxQOCGLPz2Yl5IlrLHnSPcvGQkw+
viT7NGjsTM8Vl0XnhL5WOelgyVIk+4VJFlDpf9Fa+JnbxzPUvVkhzcpHhQFvSVCH
k9aXI5UixGT2HXyo9mXYNwfEtkGWH5pj9JaQEKzeGa22wMJMs2HJPrLN1syWt+OW
AbhpL4jcuK3CE1XcN4RWil3FS4fApiBXFP8DgHeoEm7s+bopJyA5xxRtXc012z6Y
N7Ulh/ju8z/jsKuMDETNXXg1WcilH1EJIly4Go0TFqA3Rj5bbql9QHHBYQP4HMtY
f/7QHpyojVFZ7b3WAwVW1huYsH5/aX6pRXtAPzLIeXlqfCojnfY79pvZMcomAtnu
pGwAdAOut/TKjmEypGYRIuZhM/knU9GkSt2OnzJBhGk3foQOndQCgq5lS7g47hEO
/FxZSj2qreyvcm7gxOiGrHbIdEPdjLbXWb3bRfrBcIzc0pYBIcGk1xYXpfRo1AVZ
6dvWU88pthFcbV1T+EgdSpJU/KMqrIy0lPrLtkBOtG4cCugZFfe0PkF2Dm1cMRRb
KLkDtwumXy78FoF6Pb+dLr9RMMG2R+9SZ4l4YlfENc7X5YX+MSVq6YVeDvqyv3Iq
4w+Kn+8CWDDoC7FvHOyKvf4GYvjLH8T7Da8nwBNa4mAR+ZeTuMiqLl6A8PbRpwGc
bQOizPioODipyQMMamagQBwdjClpWYEY1h2jaRr1PTV3Gngn1glV1Wwb73cfxsTN
17jGEJaVCHnKVTphnxPCOGPa02czxe7mLdWQ9niS2x5YwWBHs5GeWr6t3aOoz4Rw
+mRybZruPMy+arojGTYOstprqWdQYn4TDxA/eVnxxZbNZ+WX/QsVWKGFC7bXb9cM
yJtnM9zgXzwwyTyRDXx3SVuzYmNDKWTzCwL0/JT9xJR3CqJJG6OAdsRMm9OSHcWY
kU18Uqqv9W0UNSTLwgEz+2Qdzd7eN/Xki5l4uBcrTbT2UR5GwlFpeQ0WDKHy7yUV
uHUUnMSCOE8qdlRZLQjYEV33BWUhNDC+XexeBKyqd6/QLb5FPXDvCkTJ0mzIrG4H
WLvi6ONRLV1acYmF7XGK7XNJIBqJzsviTk1Kw+hr8PVKd7O43emo3harAovo2cwM
5lkbPpboCfIsVoHj20FEkkwcrYpnZ80E7ymn0/ZylfrruW3mN9fc/SHu+8qr8j6U
856Z+VARAqhHD8eImlkcPrTqY2yhLqAPI5MJCoJURoTTg4DRygujXgJFU8Up1fw8
wNIOrrvzDdzebNZUPblGLm/B7iCX9S53CjBtvLnxMzJyQ3C988aFmYbRz9MO3L3+
23seHGa9F0MzF1ih+3sUtU1lBTU7EdgzcrDzQScJWR9NmFfbyDbiOlJeqpdYpdWY
z1vtbin9BcGe4EH4L/h2IyqaPE7MuYvB4Z2ut99VNLR4PIhbPdScesNvGHy8pI5d
UfyhNa2TqwqY3U05m2rK4pwy0qsPTj0gBYyxomtliNxnyZhv3g2Ec33lOxVDaRgp
arX6Pi/EQaKySKK7db4xuJ2ppg72+LgbKdzufn74vUHePfiUfK6VaLu3dkuYKdD4
fs8FAdlurqK2QQUwma4M3P9eMwQE/qcigcdgGwFIn58qQ3RxyXPoXzWxpg5E08xD
r9jNvn7QiADHM3X75zTgO5ijRlTPwI+AIW5lLkzNJvmUcgc2NIy0q/+t3WBUIEOY
8nmLhho3XuLOCQIcer6eg6a7r8YbIK/boKrNrn5WO8u8AyfqX5099GXqBygvFaYh
Z0encDpdmLB3/ZW+6ktorMKnzn9pqHNXg4H056paQajJ4fKnYJR9yrlp6gi38hPH
VmOpJkZDgVtUbyVwSvzasqpDCbRFnqwBleMBpj/L4UOY/us6ot0q33QcZ2bklCpq
ImVxEhISMJGK3xQrRMx8bRAOrCSlQYqaXb+uis67niBvbweHWmCt3hoOogBCwFvd
eej954681HbOVCDA3Qdu0aF9iRHX9m0r7+n2NF6I7FUacN2MErowepeWJyZQBJU7
cjgOtaCD2GxEZFsuIZ/m/TBlltYenS7N1b4nIHMpNT8FMe3PmrgIfzajq8qoNooN
vyMnDOcPy57CysJxniQf9ll4kEk1PvqhkOaITHf4CtWo6DymBDAnV/MLydcGn67u
J9R9W11a6XV/OhvkIziVK8D7Fp+Im953AFD07E8WNw9XZrfUg2PCuTdKZLsK2m/k
L75IcFs9lN3RA6izPmJx3cXYMr7r0+CU26JIHcQ5MvpzeB4AhRa22uvxlcsB+NXd
Bt4jn7SydmgynJLvXkI0m77LkwRJ0YF2xBg3qZ1pNO1+BxY81jdKgBD9IQz20Rl2
HTT5rYepy0gsB6CKcLF8kKQy21Wtzr14bLl5eL1AiSTNO7EimB4EO3i2V9kuvtG1
WRyByiS5OjoVTpPzBtL/pSWOMCXY/gwhFrwCzJ6UbHbkQHP1NaAcOSW1mN9uO3mo
9Gj48bUN9v91fY+1/tPE3URWoD+qHGusbgb344x6N3KS11PZr30wst1XLtNdQxCm
D6D0DiECdFewI4yoPiLlEUUSoUgQEXsp00Q77L/tmRlfFKPGI5pjDjOFINa4APDN
yPYcsLaeGxc/ULZWo5qsznww1FurjXW27WsOFwi7lnPWqBQwfOTJFcxIZPgpIjat
Nf3jazrbIIT44kqYmq1NwqbhdN5nUUxrKkj/lm5xlMp12vhFE+4eFEM3596Mxe7u
+moaDr8IQ4tOs5v5cvnCVOZXOIUxdBJyalYcZRyYtv6pRV2IZvGWctaZQYZYTEKr
EyrrVLiyvH1lvMBLoKq4m/aEoeLznXc3tyCoaeafaA2x3Txmq1b3eF6WuEEj3POw
W3QOMaPPhhEQTwEFF+7yZBXn1vb8i4bQmDdzYZ/U2bZcjU1YXo9M8tZKmkdQh2P3
2JYfM9uIVl/3pv1iI7V4WvbIXofD4njE++T9JN2MAyNYuB8Dl79lC5raYKfzXCgA
Xq8MH3x9Mf2zDE8jGUpqcfCiF1z9sr5Ot6lLsIop52BH4s78k+QurE1+yQSDL2Mm
GPQelqZEXiSQUEiliRwujeWY/+dVdjNhAz3cf60zy+CI+upYWSCnjUYYSknmZOnU
pxQHkOARgpNBvkbuyAwjuljISIumz09gTadcQbTa2xSEOp46piLpB0RJCX4pQIFa
SsosADSoIFoTTBEQxVb63/gf+asDejujq45HxfcYHuGwV/d0DfAvIVSHcYDWiQZp
L96EKKqOsV6jtygx4ioDcj/mgOI0EqaliKSqwCW4Zp5CkeqxfQxLrj9SmdZBKgje
GrqwvXOp18jDO4pdoB4mVgT68mq+6fXQAOhgdhILcSx/+Wbp0/Dk4z0CRHJYuvT8
pJxQNMYGzC2+vkLgPf/xzIXQJ7wqJSOpn43K1mNOGw64pVtF4BKKA2iywWwzop91
YgVUcwe5LPcuM/PYVswLppyPiTY8dwcE6Pkj8oo2p/tlsGnrnKDjOugJB92qkuAC
hbNYApKh9PW51oUFkjQU8QnhoMDwsqFUdFpy0APZTSi+vOi460D1da0eTdIlpF8j
jTnPqLLB/uLqlSxiVLtL9PM2NF5KYAdQ76yN/sCkBayXtGcDYe9jAV4hhRjLQfCf
Qby8ViLwon2hbzY+57ajsvgdbbs0OOBGlgNhYRdlP6kARb4dlvvfIsrJnsv6KEna
cVm0QjYpCGzghQWOcVCz2WQffWKgXp5L9NgB4MxKyY/VPurdCFlEBlRR7hyoVW7Y
PktEECgr+s35aIGOjfBYsIJUN4FuqJEe8uqzuVQGZmQ+IJdLpIti8cUN7GFrcqrx
8qZ1jddjhl1JCl/W65Pt6t3Y1+CMknvbAl5AZl357VSspGVGXMIRckeIOs72Bs6/
f5KVcoNaGNIbZ83Z6BHKqqQcsrhZcWDlcHdU22kwcdXWCyxxLTLBbLoQGd7HpSpU
asqeZz4U3Rmm2vRngk4OwB7xKIId3UVVDYxCjq8TpZy/Nw+8VdhAwo5tCfE6YIBC
YqrZ+0bBuh8FqpoATGt/vMQYxGOpVDGly45SAuQoKztA4Mr+WGKWS6PZFyHL9+ep
VKaf4Jn8LJD4xrtvnwvGPfFTJS8k5nG27kz8XZc7901El1oEazmRytRv2l+3XvM4
s0DOsohvrENgCizZ9JSWThCQ59wUDKU4ylymT+qS7Pf8aRBTlNYb+XLcg/wbnCYE
Zyf8TJomwv//wCLu3uM6lm4fRKnzpyP80yOMuDvtepvFCgE8lfvaVxw9VB6rt9xz
iVwStodDwO7NcW75CIrXZWxNAAZJs1fq9Gj36vgev7cOyJT9xoDc1lu5h37VUWWg
lqLZkp2azMvU5MdgzM5R38rD4awV7MA81U0bG2eTKeKT2/9NBLPQeqRdzGBuK0Qo
tot86xBEZmpZhsWitwEnkjXSYj9H2X7D8jvuC9t+LRAUGreo6XkGvgiHyXTgcjUt
4O5VopL0Yj7UU3cFYzd2Z0tY4zyYziv75rUq4r546hCLU1HOhfmsSPM1E2Hnf4uK
f2mV1QVkWRJcLwQZpG1hwQ0b27w3d56YdPbqRRFYeDewxSQdJb0nOQBEi/qDfAt7
F+yGjKlnQUm4FxWF/fPCssZfsf5JBOXVl9RYLTd3nZM7ur4WTeTIQ+Sxap0tlead
LrlCfbit8HZJi3Y2heATpI6LIPveLGM6iQYWsQRJ0NaVLwhghlRvrRsjLV9X4cbG
k6FhP2RuSX2wrzW+aeU51hBFTqhlywSRModEXANLvibYyB4Z06V3SSRrf8QA1EgQ
GqvhyZcFHifUSAMnXzTQvUzQQVEhCk3ABO3UP6256tkydp+9gC6d9hXvWpAnDHx9
ky9gIkY9Ke2zbx6VZrYmZxs50OuBtjp0Hg8ahhZ6yxJxU2D7WoWIgjfMGIPDX9bd
ZWujtFCgznKHa31yNXzY5GTrQnm7jzdvdEo+rOTojAtwfTVDwLlziZZLNu8MO321
zPx6dHmX9NNuFUswo302eC//dx8sMo7bB6Xi+t6kt0ainPzR30dLVk7jTzT1sfxk
092BYmyZhb/A2Ipr3E9L1d6dwXGfXcqDTvNEeOLd74hHZ2DU6RrRgfrPdssTl2gS
DM9ZkDkb6IwaTU0Zb0SVac5hEioRQwPF0Olhbq3sl6bMKego+aa9fHufVyE2+bq3
BBMeQZSAwGz30wPiWqxW3XLmGDaqtDhbQGQYJUNpSTAd/MEuPoWSI320BukndR4w
xkXkTPdaPoTmSK35YBeSfua+gqzWP0ihCn4CNrpusakptNO+x2loQJ7cfLAPTpFM
QYL+aPJOTvjJDsJJU40WvF13U6LreY0GHMdH89a3AYvfYTFrn8JkiTYWTRstU4eY
Q0YQaCm96Bz6YBIY+eqc+oFszKwX6xdTHNXLAwUqlsDOn2WNr0wi4h79pCA450yu
GWsHSUVwz7b/IkJLa9c1SzFzSsaAi2Cm1jUdTfdVPVOP8nWPZ/oUb4dxEV1dXhjF
ykEnCIv0H4kUtLNPg0h2WEMn8NjJQwY9kHxEwUJJQWRQQbPA33Gl1PnCemyPXjJh
ohaVq/5nnKqJ1FxbY+U8YF/3QjUOJ74pp56RyQQESKQz3gdwH4e9Z+C6ze73BVWz
PbLAz08GFfWiRC0q7cQdviZ84DhMk/TQ/yrYkHyWmzqi7wDmUybUBKycpTfY686K
FTrdoSO5fdvOLULdyj9TmqlT/gz5lvI8Uji10zDAYQy0IUnQMhEx98175iGMQcoS
S5XnYmd+CqQSPXUjxtjOhra+eeaOOA0dCvw4JsV/7hUoj0jXVxEz2nEh++Nk2GjI
7Ys0EjnOZfSlRAaleMm1drGbAhvgeEg+QSHQLt5IEHjA0CAmMwyKXLHkV32bbRQk
wac488lj0iBDINzrVhwPltLkS2r768tfSoTxS7rVLkkHRBhPp/6RrMYTPZQrF0t+
8kqRmq2eElYf5yeZmCjJs9TBXc6SkoesSwVPcvKBlqaoa6cO0uFrscBtX/ImUReN
oM7+ehpJN5uufWET3qRMn9eWoKuZJk6tICKNXhB1qb7oXPCcD2XFUyhd4XEqpPuF
q/KkIJH3G3hVNIiUJBU0Q/LxNI+7hzEkdgbFaDLRR0DVYPtxz1m0bI3mwzYmIYVe
yAIDTRVo54Lsz5BMkS8CvwrEdr/ogF6Y+6nwtE0xAdAVbXxC5v0JEOJYsGZ1lbvm
saMOcz658fjJ7KYAMzHt1XYXSCy3imkpSuKV0yrb9v5CUKj7IYS6AsIVbN8DZcAv
eWgM64w/uAuoHe3k9BK4ApM3gih7GftMFtEks0BwZvXLcLSvsY6yaS1zbO1nh/1y
ZEds/TD1GGJJVzjxCAD5voAVOPyKMZHyMa5see7w7v6t+vkajyYsnSW411uem/fV
GS4EQ4y/83BkAJNZmO1YNDuVzQ60tvtGDuSjIQLVoAPMI3HmSWeNV8sdGWYk/Kuz
HelwD+6G8Wq7uqhz6dUmB8gsdo7L6cst2V/5RMR5UdP0ZHB6kg1fzvYLnH8zYVKy
v6XEvZXofpNhtlkKKM2DCjbCcnhE8Lt9NQ+z2ombMDNj150Jr8ZloagLxRIaysrg
VJU6ysAsfIOYsSIUvpFsBVaweBdpkiLu7LlNqEv3ANJ56+dMGSSxNNIm+fiOY0/b
A752bbbAiQsQQXJX3EU84YhpeavlNSyETFC8SWGfCwPJRZDk4F1b748vOvGxs0Ff
m5mlYufhVpFk+eE/YZ+m3LYRiXzA2kNo+VsV7CjlcBbhtphqM+L/qNAOGrLVgESd
uqiOdyGxq+mj/Psf0xUenBIWXlt4HNcOeEF0TVNzPryWw50b0hxQHWMmrNk9ZnBE
ngtcTEtJJnWSuGt3sb04WVXy65nh7N80MeaBhO5nDTt+lKGG80E1uV1+3UiUllkQ
5J5X6q4SiRIZ3fUO4NOFOkAzB4cZ1Q/ljqNHo/Sq4Sc7YA9MreZbNrjismhCCfGP
fnmFQMlBl7+yDOtUhEhJd7rc4sBhiul3AT3eZ05ucR7jCBIMvbsx7pwog84zduD5
YVBrnw1tk3iOxVThFX+O5TJw39bqX+lK2cdqi9aCp7KvGAyCfPUq84OS6h0RbUul
jMPb6glYPr70cKFiBKJH4Ui7Q9Zj1SYu65jwYF1MtaYr+I6+FrNTWA9GfmVDJ0gr
x4tnROZlLen4ptbrt+re4JJk3Y4NLH0PgHGUhMCl2qF7wAbDr/LCrWx0Fo/k1HWi
Jli8WmIPdY4NnTBMbm3keV18c7gJzfdO3UWz81VPAib0rNBDioCOzx0jYWHkvm/1
grwsGENwh3iH/aFp9TXnGhvj5mwMacm4Paj8rHTKhTRQarM/VdZGkvYeeAtcgfFR
u8iw/Ah5C18WEYxDnmm3aUUBevjPdz4qX56I1F5iakWgku+wyUQsIoHemynMXVP9
KyQKtCRPki0uzxUMiofORnILTGqO1Fhc/Q8jsCeTpU/++to60m7zuHFzl5juG6Du
mubNzj/dKiAP29/tfuC5aE6d0CDSxBmYAmEo/0yN4rZlCD3wxlR0We53UhAcQ6oD
CR0b9ZwHouck/pmGYRQW8M6LCTeeRBDOtiaHVmrkTVnttp1xAa06uJw/SndXivRy
NqD8qQ32dGNGcPnqwg+dcXjNLZ2ZaLFWIoBm8UNpT8bSX2u5j+jqKIsQ8Rh/4Bfw
agCfoo+qRQQ+OX0gEUB4AkYL7/0dFpvfo+XnIp8cePHfBLfdi5KzE6TpN6Ey19ra
xHJ6stTHXuSJFx6AsBNYu85RYxVFQtbzUSVfvcOQjHHHJansW0y2OtTOSvVF/HEk
iihg27uZ7EIQKRpG6Spj7FwrjzIhMn9PoSVp/ay1OmD4m2meKdsTi5y4rERdnsGs
MPr2Cfoz7xPZ1YtaXZ4m7FVUAocZFwFCcphmto/Gw4H5k6CnCSb/q34Z3RrqHj2F
RceK2W8fFUncCgsv5sd9xZg+pAZHXoOLM8kgFPocAMF8ymoDa+ZxEkTQraPbQUiM
ggEaNhVzfwHEK9S/CI1YyP3wXn296TURSTBUK566gFK/8k5+e6ivJsG2MHpz/J15
YfgXpkU78Y6UCx25ymn8yUQxW9sKjzKonOn+pDWCkBh2so/Lnb+2bhpuQA62ZiAc
7pzM9EZzyl2S+GgSkxufdxhBIkZfzHUmcP01SuBTNGVDLFCBWBLUl/ep5AogsVuN
R2J0RDJo47akH7iCaoyTAG7s7fiWGbXhJHjTsOtpkTdGBhbB8YByzC8tDTDcz/en
g/R34CLjh6ULyqpSZ00/3LDtJu3YDeY87f43DmM+R5vgpK+dM6qirn67566B4uaJ
OtGxHG4LfqTVVU0FL935UCwLYY1iWmxJkdFnN0Kab2nuX/XIa0il1+kvqR3/KGEL
kH/QN8KYAGUQgdCvPwMBia0AakhFEsE1FQPOtJtDiP7sls0FPXbKsNN9Sg0XNPTr
Bbohl3wGX5AwcA9SYIQboKB5Y+tpn5dz1HkWMXTBZx7PSxbt3rPVotGMwuaz+w59
gMPnyZ9g+dXdb13vf8kLV/oKawSJgUC9TFJOqAC5zhwLC0nJri/k7qrJDxtAUZUF
THMr5CN8iNASDsHC1RcZk+Hx3+5EvQv7fpaSzsXbcu9AyNCXhxTo8fJj9iH3pLDV
FmAjz1Um0Y/zsyZ0VMz+qaLDQXU7Wu2k9ZjGviI+58gZdVLu825voMtu9K+LSYC/
Lzu/fcGSCwPlzGI1p8ZAWnbXtL1Cn3yCNrAqRyKVP311AbHLhDajhPUVQk7mYwFM
XDw9FnZvsrQJrwM0QpKlKZxk3Ltqo2ZGWC8I1EU1rLfVFKF+IUzoDZWYBdgBLxAK
HKgUjw8NKTJcjTFXK0Iv+h+2djv8YWzP2giUbdg0klVhM2wxpzXjQdKQUfmGS6/l
FkKZh/3wf6h2oHZ+2eraBPfOSMhIjivD01aZnyDgsM8JHebc/wpxkkcfjXziA2iQ
spFnTj6K5916wz/vlo/YUNsREfTkWJmFrbxO1Pu/6K/NrU1wAN6NmygW/16TmqH/
ePEcxv5nHZ1tSvcPF2zV4TYrfOWIWEv47EZyPwMh3yZ9D+hUYo8cHKNZKT+vAOjC
mtH3Ub7+kO6M02FXLfcdhCgIUPvAnFv+reN17VeO5hx4qYEBvNwrxj3CMmFNdpyY
CkYcyxPXInUbYvRgZLEsT8LWhRrcsZ7aaLXrvAG0dO8bVlkqtG77etPNFzvy2CCv
OuCWOYdcc38GPgSZUdMHAizvrTqcCygHtfSqPeY0M7z2slhnefJ90Hx2VqB1unzB
fd/MwlpUdczhy0rYz5XxPSh6oLsZQosQLpOlyl+S3jQQI8JSfm5McacmOEFqV1Is
BhMF2QZREZltokjcs9SO8lPm3JdMo8dBjSL+pv0vQOyMPFQ9A9e9COXU9RVA6Xt6
jQ+Wuq6M7nkvUdp7m8vWYdLL3ELVeMrcE6QIR7LzA/cdnW/q93L3ZIER+wJy3bqC
yWQWTek42VvWucslNdhkGTGXHSD4REecMnFnruZbT3fBUDbt3tnvnrn7GnCeZQ2C
qy2NQVm3HkHkQ+atvQAbg3DpMFZsbKfeeMTdYTuvLbAocg+6eeakCOWVslSIMmWh
IYCj+GsGbm7WOlflOpgsIGGMalz7iAMjBZl3srmEWF7sH49DFY6y3O487/VAYPfr
0VUQBZLF0bYnmeiwLj4UAZgK+JrqrAHiNL2OnOpnOIKLxzcA3cr5jPNnF5RNmtwN
/dvX3QDW9A3fu6+hYgz1yd4RsKtJyXRwh47JGWHejVOrhp0uBfve4oN6jQO74g6w
LG4ymvIE/+7bZcTGfUPJtpWN4zkfM2cvQfTSvjahuSyyqGbPWXkk7+hQz24HGVTF
9hcyt4fIFOCC/rgl5Z5DyBTA+XiImhMEdwugnda2dTsrK06eI0y0R8wGEyyfLdkW
fM6gXJYoEmNtiOUGnqkVSAdwBHqZG1NI1bwr+jxTLMDgSaNWaxdHFTaSlM/8aLtQ
AENRSvyaQC8dGqpBaeR/LJVH/gNn9CtQPjYEPg8NGkPCyNNDKbGd3Za4m9ZvgHpx
yHxlevM0aESNrUYujFbYMVyMekIWjHb9subh1NIUlnTGcRDeFXEHE7EyzbjWgy8b
8MZwucjXYhUkyOStITOk2BIyoLymfx80+YDnPrh9pWzAFKTE8/NUadmQrBBXGpMd
+V+K5Aljpw+docKmZi01Fam8I10zV7aRWIKWYl7+HXkBG/O87icPn80SFHzZf64R
f0ksOIDpy0VB1aRtemGefPQR48oGVR4Q/NASC3mkVcIrFDIyGcIkhSVufNY6+32C
ZgjTlLHrzZSIBsYz8NAyEmvnTDEJPOiRxMeEHacNLRUgzf9IB3dOKfy1lno043BT
yiO2HTir+7rIT+VIURaqRN+sRyB96s1RyGx/krNohRZqPko/pq9J7qCwdGd78J12
feUMmr5aJYl7Eq31uJv1aH7lXeZv4+EmbH+06PMDG99N0TmqSMbS7L+OucYdsqo0
hoCmHScaJ5Wn79irqTjKYTG2rd41ATCUjVR3pCkgMbhw+puFH86ApXf2VNTKiiGl
MEUV7EYXQrLb27jSyzCKbAyZ4bzf9l+cV2xauNnO091m+icgZifWNFa3PIBoX3ap
CBF3HfuYo0gH9WSCDrVJyk7TjedzoZpEbkkUaA7fydscfYEjtfRIfAZIFz0rWND+
bP3VW5NUUE0qNX+xSt2/mOSwHKkcfpzMHdERxNC0wzRKzu1jjpJvpPR8n1M3uAQk
TOXyb3aLAK6OAubuzxaNplgeC/CSO/VDP7xZmiE1uE3z0ZtK3ig6IXwJf1YZ9n4d
UD6pe1QNcqPzaozTFQDYp4+L3W/0ZueadtThBELYCJ2MIoMTcvdrjNKPcn0/cBGS
Md2Bmlc9COXGifPrRLaiMkRl8qglzjFkedz1GHBWxaSpDgStGdZ9KE748frOaGoa
NUssGyiAC1XBARP/8IX7RJvi0iJ96j8uM5QnwcNuvzT9ZHukzv+2MzJf1qTD0UeJ
hMPBlh4ljcCNKpGBdX6CuQTkBOW0lfug4wQuf0c9n7r5yWaxrhGGK+hRU7nFjATn
odR52g/1mhS0lDNKJbmTCUu4EJB6wAYg06S1VTHONM71xo0+J5Dqd2SaLZj7qZ2V
VaKruBCFYjOOeDpTnsNN+oFn6qSzpeo9GNsFVjoJeAX6K96ymVo3vPaadNBCyky1
KSPCiQLAxGCPQVJDMESTsP9fXfxaBYxB3puTkiXjSYGD0i6Tord7AUDMURgmXqrW
BhoM4Y397HmJOmStLKm7w+l6+DDfXYQFYLmig6Z1icZVdAcYNeNWaJh9bIwgCLrt
rvNarY8HeEiilft3qqM4RgKusMr1Wqsep4YgwTxXn/Lr3WcS7gU7x8wHhQ07GNt/
KzSfZQI+u8faX3MUQAxSc6IFbgiZwXX0UsZLj5iuZ2VT76cKPgiyViYUKqp/Bk+M
pVSigsVOX6SfzdoZmVLF7spaLHl3dRl5pilwecJzybSdwM1JpJTJsgJJgNGBE+fM
Ifjn2uF4r9M/7LEQiorvWWnVvHkTiRqN3oWQeVKRRIXd7SfDkKW+ciZZ76QQRvmX
fLmcG1dBw9srPTQO79kjUhLrYVlz84gCWT2GEXH+HRTx40tuc23kbi/pLD3S2wLB
2UUxftvutRGhVA9bsqnb2HUMQb9LvoPGXYVKkP8Y9XaLFiD/1wWACSy2Bn9q269v
jxHG0+ZtNshgsfQOvjtXLvb1SAk5rdRo0BlTQdTt4iiugpKUHT57jaUz8jgXNiD2
Eyualwmf30R4/i4Qw+7PMIN0FsHI5IH3x2oIBeub7tg/b3IWv47ELxanDExFZyCO
gSKuX2yyWMKBc22PCHguULUsckyLtdEyKqFfaVuTD8PTIdw6RHpCJE5WPzSDmQSL
TRCHjcOmXz4SPIadAneHXMvDx4OlJ+EJsZABfn5ndtuV1vRO6eGwVl2qKKOidbIB
rikbCSnJ/g4Q1tHzeiNrWollbklyB3ZRvk2WWEnczcoXplSgn6ilwPNzw5iTgVPr
xK/KPI3IBSZUL5NnUh7GphB6yRRPpn3RkekoWxYUs9Jc9g7/cd0P6eNy3sfMyUi0
/a23xGpqZ6gUPkJedl19eXvDAdmiMLoxVbwnYw0HNwihqAowLPwa1JRtHkSdObzH
bA7HIoFemqzplnJ+tIDu8jIw/iCD8+aMMpgwa+AAKIaUuPmweF/9dBdG8T3kVaB8
q3kbFOXijstsWtLZXGBFVXTwRSUtpjSfm1+lcdirmHsx8+hL0/XcPBM+V40B8NbF
AQ7OM6UBnZ45lOySqIEigAzOVqKL6dyc6TH0K5g3/4608pfUdurxcKQLGItH8NnN
FpDtpSBbRJO3UmKmeeums/usJd4m640nv4sI9lUNoaqtGlDFnd29sfXeNenZ4Kmm
ANeA1dbSIRSbVmeSh4pAlGFOMfFnA0Msmn2AeQowpIUYkHmfpfK9vff5suhqDlLq
MKyn0YRRWcMWvQzVXx5K0iV31K4hY2DWx1Yo9ppQlAOOMaoBhBSDstqYDZyjaReg
k+i6DyWc+kbC4v+1314laB9b5SdFEsIcCAS1AObfqaiW6BI5NgKY9yezjJ8NuIf3
xihvX7d6gE6oKyrAmBE7zlswtIpzw5mgUjiZyXkbo1TBGK+R1CAAmHzRnOcVpQHs
cI9u8ZVUX0K6tox94WQk5rW+qoldD90rOZXdGnQJUjVEl6VABKs682CAsnNn5pMo
Ex+NzCLIiDyk0ssf68DpFgqaa8r/+SFd+Gwt4mmuY/CKhWiM6A6NjnaXFXPp3OBu
JlhMt9Q/4j+dY1VQbYHycWogZA7f84hqslcSYg0o14LJgDE2ptQxxQFKNL4wdgq5
7vbU/QixpL8NLSanyVDVwnrH/vrDzyXDmJfULlBJ4uDKxaz1id5Iub0xqMOKnIPA
XC2GYU05geyw9j4NyQ70xbFnC7EYKkXBA2t3fDCD316ZJgsZy/I9V5RhpgtIX0zq
E0NeYd/+u310haHQg/aoq5l1ltBasJfm5HsveMpObmLKZN0BijhkdBfSiFXq7Tjg
NyAs8DOga0VMXwIF9lC2GisgNjYWP5ra0+tS3Lb4uRp9yE3T7GSbX/d0TYsUTZrH
hRBc5YavpvuBogDBGVtVOp7XJV2EGa3vWz05B+YXQTiGJInvaQcwTi5mgQ2pGQD0
MNkO2Abi2Cl42KBilisg48zzFGWQ3AMh5BjEAoUtU8nl3lrj8ibF76PJAMUtuPlS
NhEl4Uhwqaa+sQgUvszd7z5aLbiA+gX2ScZXN0CedjWsN+j/k3GV/Cp2Kbra3YU7
85nkEEKlos1zUqWzHpnI0ffEDD/G++zxgOyMf9/w/ZIICdb3msavyJbp0f2YZmoW
J95EFOZGi+dTSxJc4VXs8yfwBzoEo1UUtOwY/ARFfTJT/gJl3HAUkpg61ytnB/TM
OISTh+kGTmaH/ixPR2d7Kh3AnRZKHs7eON/Zgsez4xWhUmVgZC96jp22XyZgrJmn
ZM9pwvP437uysFPX3Aox7wA5o4LPLe9ZOY4qt0GgAZi0sBHbehWLk82UT0e4r3BH
EcRVIVmxj5t/OOlyesE94oDQtARauL4iPHNf1Zgfip5zp7W7BS17HYT5/SIBT4On
tuRhOYoN9QlfoZLL/rn9AqyQiv9sgCloe5canYdmsmLgdXMEnfufuG+FEw+PS34j
R7OnlrWa9JgNEJwk4D04jwFsP8IS9hhRYudNK70Mcvw75QLB3Kqagxk8TI3NAUxs
GKMacUkAVI01LbfJvy0fPbUo2iwCaiy69XQubJUHNeuyqCe0tR0YY2E/ARwhSMt8
X2EqS3036W8D9zAddmn7LBX2XiQTYMl8q5SnIqHm2Js0U+R7nBCAEPH1TqrGLijl
yGqCtp+Hru7a3YjdQBAwKClIO1dnz4NmypAelS1yxQFsH70UuEFtkeb5OC2vgIy1
oiZ2qldHoGPxjK7ktX8JqYnZGYfr9bATsn2WNWl5qHGbz55E0YL+KtM7VxdryCNe
vI4bd+EsDl920ECY162l2xNjh5Q05/JOQq7i8+Ll2ldNZt5w3Bk2ym302GSUs4T/
4zOK8oS28HZI1ZC8+BjQouSZTpsVYgcRkHKWQhZu4ivzwMrYwaeAM1BBn4QZ1iKG
dPiw7u3VDL+grmJaZI3oVXZsEaKkn0+O2NFoVIzIVD07vhOkbPU9xPrp136T3Fd3
iuacNvfEl0nqk2U4nbvxqCMuTbHTcZvq+KXk1H9o6e7YjFBmB956gEhxo50j4I4+
yYJXMY9rcr53WSJw1u+ENLPsomoO9k3GKO4KCAH4LZuTlscMmZ4k3Bi5xzn5AF73
nA8IGN82cL2GUIaCFi54Ramo4fvpo1LH1WHWXj56zzVcXw+twuTO7Zg+hZ0FNLWl
lxbB3hvr/7tBLnmMZqntLsvn1Glaq9EvbYE0SviI8YQ7W3GrB93A/wDBe0u/7Wji
Gz9WRDLm9qjvc/H+3MIGmQQ6b6CZjHyY/ctFXMdexZhqoFom+zj+6Q4LmtyvurGa
WvljXetbsDxWIZG7tMwZ9eMApbHbQa5yDQVc9ZlQH3el8Cda4y/In9SWQT9q7l23
lsZkMjQXx75Iw0dpqgkZ37dzqTNEDoAlmStr8qQvZlrpjWq0d8/JAAeZnggXUrsp
AJvJVSVDmkYoqQYWdYcmuHcN7EBIDrgGX+TxIdDGFA25o88pVREgDS9Bkf6I8/1Z
4fLzn0SRmvch8hBsP6z3Y8jU1dMLLSpw8lVUESTbdMqqU4cKiFzEYLa+XaLCta43
UWYYjOONvmPhlAJqYRoe0L1JYGJAX/CbmKUtPxlZIoiUfJSMBEnKcJb1j/ZPRE4Q
oIR7NUJ3dIpxmMTDVJ8gqYDgPy5QV6uG80Ur3Lo+qMdBr7o7SkQhVtXRGNevU1+s
sb0wrF6YteQ0ftZmI8ACTRfB9azORTOauK5KKwxUBV65fLZboRM/kiuKiLnz+vuC
JWPvKYrKCgh1cRggZgiwN/CWd3djXBHYv77Tg68HYuFPQTLLRX5a+rgofT/p1EAo
eNxQmRUDS2+guQJVtBC3wZVXqewcQmUcClP28mHtOVv08tgoEbrtyWbl1ml5058k
JW1uI1fJKjkP6WLf3dF/lYprH7CpoS1U1sHPYMHVrYL1wHNx0OVz0vNeb9YeNPeH
Yobe8BdRsFU9NS4avk+V0CJTOyGVwbQ/N1voZMWx3CtB4YF868IlkFRraViaqOG4
O/Jl3pBO+tklutTy569kpVC3YJORKQvoTsDw3u+8b1y84wTuv0qPiCzrSqzOqWuo
PgnPbIZd4uabYsVzo3qnFXsBUwuSDUrNZ/7fIdSnRhVQAeAV8IK/1BlmNKwsUx1x
2yfj/fXw+1cENyXZBS+jhG8w2nRs7e8vGM0MNNtT1s5KZ5Y7DVCe/Sh4rcXaWpjS
7xB4l9rl1VqQWFzC1hhd5pz2JYOCrWRJcL/IsfENeI3dNe/Gip2iEOjIm6fY8chk
8WUXpqyNV6VO5jiE9cgk+j1KezwfXtofen80UJsvmR0EyoLVbFv/Golnmkag3JC5
+gwxHqoRevxNBo1BcjCQP5ibBfBsAjxjlQaryiL58bqcG72Xt6obvkgGwKuk0QRW
YaofgArVajAqM4Wji20a5iLfbykakt+olOe30RBrWdeH1YmuO1rTp52aZFO0SjYv
i6dR1s4t+77h6ZmyF8XtIhQshS5NLx0w2bOZ8tCYKGq6AI85UMvoAQkSqHUvmjbt
6UOdDTK8Oq/HB+uQD4Jf9s9vWaXi1caQq+f3U0CA2+xbwHybqieuciuPEekLQdnt
+dD98a7hvg7ot8xBitnjue4eRQ6zFN92nOeMarYUNy9EdQQsrvJQ3N1ks7wP6hh/
/vBxJ8W6G8NOa0xScc2P5LTCBFQBGISvnYdeQYQEJ6ReuXBGkr/vWzsr5mi4ijfC
Kwv6QYYoN7Q0SMjwVNagANtmiOslezMqMhL4HFP96sQytCzbY8uX1mzmloWAw7bb
MrCzNuYU6oRdzC6RWuik52M3C23pKRyBZXJBFcgPAKAyBxtSfnBxtSHoYSjkBagg
UhnVIf6Qj+lg4OWauyPaP1IfLwnak7say/Z7B7xcLomzgL/QYjKn6bYaughDjMiD
UOdBRCfZMP6Nk7AZ+xcSb4ljXmKMAN0eTFIL0EcZw6dj/VTqa/4Mons/jlJqxko2
KHRIzyYfKnnpQS/uvxHhgtivwgRABAeDxUuu4VZiAshv0+VFzAgjaz9SplWwkUmi
heWyeXfecAP2aakzlKqEtob/AGHBjX0V10MX0t1B66qQxsK9QG6O+8v5sDPZrfX8
mWE5T7TA6FuW+LvNhkbuOYhmQKb3CKaRPxh38vFK2buqSpS2L8qV9Yr7N9sqlW6U
51pEbYJXbnG4RVC3xXojPjfr5wavbfafYoEwKpfiivGA6ijxE+Efu1v4s4CnWj6/
NdTnufOzGGEPHOKv+DRTNQBccXEV9rwd8Um8jGw7XXS81lUbt6EDeM5UoBjxGTb6
goDHfIWFkbOIQ7P0yWX2zCAV5fjKc2RXzFjNFx1vIEFV7CXpk1fKYDbFfhWAx50+
9U4bYgdoe9xM0hWA8UON0H5EjuDiu3UB5wsGoDIuPXZ3tAMzskKA34bPPuXEFgnl
0FXWLptfh7eF2H/JGPXbzXWXW1fB773DkHKNyHds85fmYimSawcv4yMnNNbWnKdU
yRaPLHnWdRDlmxN8uwFbpbzJRmFgGwQxelIgnjVpkOdMMtba8eWJv/S1UVbOi8oP
+8GT6HEPuNYPXNPSakpt/bMo0kwANymNPoSa83oYZkdCrpY4ptyyhBUP6JDfYoun
srJp+v2dDARlidN3GXky38zggSA8lSNsO2o5UgWkVwP+8tP6xqz1kKART4n20mAm
LTiF39VsMWX6kUySiHVDcOsGjWv1S3Eevn+z07WuHEs5kkMX/nZs9o8b1sESxVmp
e31UrQC08LplQSsyLTaOQc5dDaI0ECbJ56VTEhOIYau+HfWnOrCbh1bt+S8n1rP9
1JiR1ifGDQy4EN1if5P2n1t9cW22Mq5ax35ozj8UH48L2v6elRxxrX5EcczhXgmk
4Etn/w+M3M6WG1feYXX7berCVDseG9wfIUSR8j/GCSVcHLocVDblaE5rksnO2yCV
EA1Y05cn+uNLX+fwj+n2sH7efOHd9nPZa7AmAtNLhooOrsrGv2O5wBdGBl+WiFjb
MdHlCH3/N4y2d8VkP6LyRmA6LqwjGKy05GpqV5qTjDFfIHAnek9OmVpqR7dxIpb0
mWcrX9vvV465LcyOr/XKCx1W9ijUQECkzlEqXdQttVm4GT4j6eCCrwM48v3CsNAq
Z30cMQhDP5gk+N6RrhU1J1vndPrm9dh4Z4kQk44q4wC6OAdkk27OirTXsH4B8iJa
pTuiPijVrAG71v6fjRPsgH3syfqCJCsE3D5De6siRIk1msOEN1wTdz3gosThcLFW
hztzRoElBtyZqDVJ41qJ7T5d89c9O/K7TtcF4nc21cPvLOXuvD7F5zfIePHhrPuF
5Z1tqC0ldno2if52uxP6dTl0f+wAhMoRNe0WwqGqrUl8y1TsqVoAvs29I8RD/LwB
KOE46ZQoOnW4wflEikNiIRLfFS04B2ptH5v8Ni/JfjuwQPuETk1J/12BhUy8lzlw
+KftfDS8s2Gh6SqEPV13ei2JdlZfFvzasy4Bj0Lj1rDJLYPhTzTeSKkTWv0nERoD
Gn7RBFX4JCmHRXUC+Hl8koi59oEjuVniVhCL67jdtACOAQBPsCFx/bQtw/RO2mMU
1gr00bDCCAy2IaZBGCSIXKKWOzJBgfsUzIm6ev7z3p7v+3X/uW3Knfzm752DJ+Ux
UkkJrQMygsuy+StrGe4qwHdOMoaUMfIePWcS6Nc7zvwYKGfLPIWCLBDebr4K7W/3
n0cLkReDPoS2VMchr3uXWSCW0pTkgPHr7n/uDLxSJObjSpgsafyjsBSeNPavB2Bb
fyQQ1xCzx8lDcm2Ka45rUNyVm1yRjiFjKEJ+gmf7vSm/UZ+RAfd0sWUxmUsO8hJA
MV9v7UA5hNQivJB+lWc8JCPcKykJ6lSiVvJJofY8XVx1xPVMOpPKX0FRUaKlKjRj
f8/WFENBzq0q0DhgaNRGrOPQp6PX9XYkbgSk7Peri1+4nqT5XlRY7vlgjmU0aJjq
TFP0kR2x/khpTz8bfww4KcnNOlWoVYdgn3tx/6kALvWgxGP7HNlVVIUB8N6bGQWe
R+EN6xFlhoxNbOCwWL7Jl11eswJkCMVg8HRwDsHh4uofDaCs2L1Hp3kegw8L/ZSH
HUvS+/McGwB+i3BmCbGFB+9Zthd7UFuwOi3AweIoztg6ytR4xyVg3Uc8jvshGMMv
zXQgNyiZFtdmSR401eC1OLN0CCm5XaMmc8CRy9eei9Vhv4N0OsKKK6B6JsQzSOHk
xb5WpCOYJBC7N1qeoMmEr3lI+mm903/fKlWlD6jlAHF3J5VYzLZAfPSPDyzRA8lI
f4p7Wjbwpykq33ggRmeMm/tnleo/vohKgBHmnj6oHM8EkYRzHyJ6mVlaQxPipu29
Y90VEvQFcT/8bd4Mr6CmFHwBpHlDabfxrKnIEd3QLj5yHHfTxqiTZHVQd3cPBiig
mWJ/pmOyFuVnFMfO5US/ZXgZWmAlySMEbM+l3KH5YVoPnxbsi5QCd86l5eKLAv/X
RC16m1F4sAgeU5Sa/442coo0wYGAA7+jsy932g2Ady27DOKIfpr9ZlTtL2J++UJL
/C44tLDn5uc/fWWPYMWn8B1/jvNEsBOG5amzwp9F5ldRmZosIuzfiFAqds+5NruX
JhJjYBoB5g+1WpzLkK8HPStNJ80xkgBr/vwQKst82Bz454e4REyrWxf5/AjoBm2P
ni+3QyLe9HmfArBZzArTvMfH9ubUIhhuZTvPZfWav+wg51bAiNzHHe7GVH0TjKw2
OOxL5u+8x5ydkC9BsGvC6XL3+nMpoZl0fiNEsWffwKYHrhTD+4uDh+NpK05dWH7p
2JtHLaWIxD3kMvAaJ5VE2+6vL8LPQxDxgZvJ6llFhjrajyZflz7zPMBWAQiJNGCg
eX8+jJ1DWGlfCtVCUrTjCwxqT9sImAr33gwWBTTo9PSjrouZmpB660dKARVjYOwV
WbQjS6EG47eIH5/mr+iDleZCYc7dBvWULEMmspE8tyb+29NdWmwrRh/Fe4BafkHO
PWMmI0AlvobFDJsUsUEHha24oMiv5CsP2S3Ks9EspLsH+tNosHAANlsX3GxPIZPh
RZKngSbNZkrs+54N95Po5O1HeW2DE5ihqi2hmr+yx77ZUTzfoC23Bhv4KXNYQysa
l5japX1xL3EdMnCiqZ975qsL5imGd3oOByHPxR326YJrMdQnSS/J5FGhwfvGK14G
AQgJGvjO5WjNGKgic6LQCqxBcKRn8R4iGZXdhG+H0j4vL4vCIJLNWV+oigAMHGqy
L3EJA81COhR0Y7YkqWg7Kg1QbOqouqRbW84gL+otdwRWNS+77RgRQkDlKAi4Uab4
6tnPOIeIH9tZ0BtepWg0PLqBlesE/ioI70N2PT2eG5obN+gkN25pdfTkw+TuWl6k
lJW+yE0edv/B0+l2cKogioOIuPl6GwBOZgR4NAhpoocIc7rwv3dqB+bNNyv7lduY
LJdXSavk0TDOf5x0bEAZKaFdxfaCMGag+3OE7Fj2u1nKFNJmoqXUOe+HPMkjq/mw
iL0E148duh4K0MsZB70Oa6fv74NfiQmWiKxqVK0ala5087hLXRK7yMTgrxVnUY9E
tHKiphbkYQVW0T2XjQxm/PGX/yFcBix1X9F57LSdG7jxQThECVgHInLawBT7Ixc8
pQThn8QYCKWjQQgD7TBP/nY1bYnRJdNNqo+Z9xKtviuKsyub8go3VUZ9/OFAPUJe
POsZje9twXLsGcARC0Ik6MxNxUfozBf0/FJpYD9JGALFLNFyQvnYIHBjGhocA2dh
GDXWIN2l5myjxRy1FN+56MPPEUlBCUfn7OE0LSHY6T+vRpjeEM25B2DUzGDRUYLR
8tAXYn3NM35vthuavDQVaFaOyqXCQA53k1KKk2e4nXGdoN2z2nirNiU5vZWh0G30
fc1iHpMBSKFrzyOXeJmXEBj/Fa4528jsajJh3mHstIisjgz7eKC3UkKFgds91WYk
u6mCb/LCK6yLqEWQywEzJNUlq4yJasVt7DBj9u7ZZVTdzbhtC1xBy6knoFpemwz5
xqJh5vXnBHaYx+21qM0V8AvC6eO+SM+9DdTToH8rzO0u8Q4ofQlm4lIoQQ5MKyL4
ME6sJSgDSdP9MEmc5Co5J5OZSsvOuDbNbxlQc7jSnBZUUd0a2JiiNyUzmrKCOvC7
9OP8Ftn3PYnSr0xW1CrBZvvaNV74C74nTJf3HQ4yjTK4ljqjJsOK67q0vHqfxjBS
koKAgIxr+NfHPUbw+USrVUc7dnj5Ko+5pTP7fwiypnqx7wEDA9KLQsbo9C2J3Qgl
bW2NNohaSPcH8viahjxMywxswzBszbRfMmgROHi5ZAo4tJVIXNQT3+2h1UMm9RrS
w+IU0CpFI3FkM9EJ4jzLfYrJKJAi7NQgwnDKOMoBHA5DGxT0EHIjfnbOUE/rZcvV
i9Xlc1RUH7I8C0HShay5cp8mmBCTKC6lSte4O1ZT4tQfQGRh5KVdx9NWLoauEmJa
E/yZyRe0zHRMVwa4b0bMaLiT0U7yA5Uoj8ot5wOGmP5ACIt47vrhDxHSMVRfga0G
PMherYHZ4pEoZA6sDBHZo8Y4Y0AfV0YVultvlIdc9VZMJEaYRvquTftFln1gInTc
vemusn06KLQM8EIfntZhxUZTbIKxs9v0JqkPJfvhJXF1l8oKxDca+tN5v1HvZTDS
OXvcMxj7iPCp89e/De4ImVuY57ISCDLRM7lvG+w0Ho+XlGWBRaLGn2vDmC6tMPl+
G7nFodrYJqkP4porkir+NBGJ6BZkRpn//EKKXx8GwRbAFahpsWz1I6yPgNOgm/dq
5Evm1DjxP6IcWlwZcMCI/wESZ9uikYB27KKX3Vt1aQHU9+rsqU/gcSkIswBPpTpx
gNh0J0YFqKh4JN3qYpPcWlrSLLGray6hEAV88I9LrkARkih082z0zbqru67duQBD
g7SA/gn8y32sWiCS3rxXOslKDQhIwj6ScUVYnIK3SqGe0GNo4hULUF+JBIZVketD
W+sA3xVphucrFN4HdHa2D9iqTgKsLSDf3O0PMvhWRIrf6y+4yEf0Ob9RVZ0+rQDO
C0YnUQbHuPAI0Cu0uIyoviQ+8NvwDI0QrUot5YNpM+Viym7KfQIdoLytol4teP+D
0Tw7sOg8ztG+vGe9tUZBRQmh1cJj0ZZr6sK8/umrrh1y49SuLB/mRmWkN5ErN0D9
RxWKLtJN8niG5GLyQl3oQojWvAkfb2X71VEkwHUS8yfL3jR3W+UtKqQM76TVjL7Y
viN6dXfOg1y6aAFMq9hls31hTSYOFYu7Cljwo99l7MfhuP5T/p/Xuou+tvXYmyxJ
nbQGJD443ruRxARo770ojOB4hLlMy+wto4hSrMXoXWClyZdmX3hbvNrM8Zk3C27k
l63EqwJwu5oQYdW98yg/AlSrfKSjprOTmoecg8i9oMPimqTnT+BiK1gDazlsR692
gBNrlBJHB3ySwzGwgx8OyNIujj/DYYetGr8ZaEBbwml78qB1NA2g9lNVHIipI14z
uhex7k9um0gUbYavFqRzk1CBK8FwAbWgsifjr1A4oq5nB7BgeplIFAtwDzWksUu8
i6CmPdF/POAZfZCrbLcAS14bs3rR2Uurr8fDRdVQ4dT6ukFfdoxjlGXX8m4maflK
1X5TxUdWTfwcssf0jH6oHN+s8K4fLxqZvzeU7uNagHOA8EuYBwzhqnLfVYlxjkHF
L+274KjdyImxKkB5F89LBF8uOTfGVXhXTwJry1LrWJMm6zM4vHR05+ZrzfNw2vPX
EF1ptKUWjt/XYKMKGQz1Z81oDz3d67oBUXbTHwOxmkC25srQgYvObr+8lLPkqDYN
SsKDwEg19MnAlryyUnLf9/tJZ7c8xb5UqKMpRM21McMYFFNNo0JrGSAS//Pqx25l
0pjUw+t4+sJDkc6MuNe73wHJcE29kJwnPh8a29EavuPI7yKJ167mEe5HpZGPjjSr
zWePmh3lybURAeEkqeQrucw6cXEjFDxkHWbQbeGkIANah0u54MfuR9AG2x0wCiLU
HkIVJzKK+TPWZmE/TSLex9NxJhUHlm7QFao/36CvlDavngobwwzHtF/1uLrhahjD
9QokITctkRCcv6WqCfqgeSHrR6i9BX3acVNva11qgAufGqwr3Bfz3+JPCW9j8TLi
50+2Lrn/LjYMSxMpJgl7BkOuoVfpYSAk3mY0ULzQLiunrM3gNZWHqLidjduyL+L5
Ue/pvOhtgn+/Re25axBZCT3ZpKYFngZlTy7FuDBo0rbHZIcQ1uQfOZAZZIco9yII
wbdZ7/ZBKpvYQO+lyPx+1S8765FlUqo4xC4SjZojk0a/hP79jJcrwBlUSP2zyO3M
osAy+1C/RD8Kbld8zGT+c2uosBKXD23SQOFLMDSpgmFGilZkAWzoyooEXfjtEFw5
8iTuWm5LDweLyhRnvUAUcejZikTmsvaXuNHoJwlFeTpR/ss01/RiEh0ieBqROs0c
Kv0cxmBpNGl8RQlSEWWPzgC1DMz98jPcc6VgwvE0r7Qc+7W6gHh0/hVLyc545qi+
MOJAzmQTSqTFEzLZDOD4R+LZQ9vO9Y/LpzlnvXeyrYj90R9w8gacC+pnwI0HuBK+
FRrCitlKjskFESh/8dYhSYv1WyP5jyPtOwg8BVIthi31dMhuBMpSzXAiOIF0HC+M
7w65oOjSFFSBIsfGA+JwFzKPzH5tLFgiKMupb3WYwORMmDF3yvQfQM8YGw45A6p6
nRuD7BgM6YfT5DDeHPT6zQBt1lmBoBJlKjb0Oj8DxwUufUcjJz7vtMVlZ2M17two
1wz/iT3PKoXnJ0CgqicJpTnzMwXuvvxBAvn9/q6GqvHTqLPgZjsS9EZ6rFksSWwo
rIMYaD4QTEf+BdtJq+H7Tih83RF/uuGSc7PMxiUjsU6oqp6Va1YF7hIatrQ6vgD2
2EVfKyuxV+/7fxwa8DANkk0StWar3m0YwISOeyLBzXaztiitPnWASFr4/b091BNl
IQYVSptVs01fpG36qhGXvA+0lliW41N4QCHEV2U6r4ZKxjmq2PV9OhxMqTX9XTql
FVrb2qf8yFEb8mTDH3HurvPFHD7IwA3vei3jVFg6NwFBOhr3Mnka9Zb9GoS2zySK
fK7CcyMb/bPEoVVP3QfHoO16UGJgmBF3Y5AYYZriPQirpbeSip/84MlvHeYfJsGu
0NbZo4XS6cNZfukei6NIzH1+H1Dnu+7yQ3yncSRgt+cV84r1ZiotdVtHlQnUVaqO
SWE4VJpowt3bXueM8kKPmi/lZ1srNhawvoRAK/piTF58T75N7Br/T21QK1xjslm+
PKq32n7i2jrQxQaua/dSbQDM9WdUvHidYdiA9W3H1hkTXyt9KKiMKsND8n3vY68D
IeMDqVXjly0libpMD6EdmCzKix1nB71f0EqRRvuv4V3tm1kZy4ZHzjZT5AyNLTQ7
khVRVjMExi0DvqmyoCK9jzkPBfGMfijz101LWIB5+yNyAFz/uaTEGV23MfLxjvt+
oSPH6N0qA2/M/g9QvM1mmICELlxLr+kQ4buntyymVhMLq0pgv/ciPDfL21SQXY0t
fVf1ivY1O8t0Kkxzy0CKPVjLWLvO/k1ePYKfjqgTqlxFZUr7ViiWLxygzEjrc4hW
8DfsvzGxgWTCWkLn/NQF0SvuM+07NaRMwp/pv0dH5wirKhcrVkywGXuelkZ3Y4uC
lLLqV+BvZAG5ZtYYJcQun7InY7gYGfR9M8ZODefzHv9K16BJdthzOwtl2/Y328f7
rau/UrHcHcm7ZFSQ76Ec29awhlUJEpFwVf1ulgRsBC2qWUzhGCmgeHqk0siDoQKB
1ECz6qJTb8xCjjCCOkPevZuaE3hdt4gXJc01hSoI5m+YAkl+BLp9YdOqtDqN41PZ
MvOb18o+N5ya6msIFVmZ1cQdomHChSKTfmpcXtLqW9tX9OwR/vI/FDMi4GfMPT7O
dwgntnAnZ3NXCPVQ8PVvfOt2Pf1Nyo8BaCEeZS9ou/RZIxxhQHWjznbkpBj3iDBs
1euB4wtf39YsAUo5gVobYzGkzRsd+Fk0SGwhVi1yStPEBrIXZKulmR8XCcgZLz8e
kNp4/kMbRbfRKKXo4UNicZd4UuazSPkbFk27fGpZ2TXIF0l5EAMTYH3IRzvxknCD
lMG5fop0SKKr3PPhj3b+T1B7KEWWzKwz2xJ2SpA+cxQ/Ew5Sd5H6v/BRKO6Zd3Ub
T+3wt4WGrnpE3NK1YiovF/6nGIjiuVndbffJbgNgEF1cOTcDNxAjtwe05MS3Z9g6
BI4vpgv23J+ZrajFW0/RG8EBXgl4NoxIUR/nUmdyUfbSuBEFHbbib68NjGwuo2jQ
/JjOIN1tiDa7RQladv5e/87ZMe4vVkySD+N1avlxchiufxspHH2Lrh7aGtq2UEXP
GW742XA6p9a0WRB/qtO6p0ArAtpqXjFwI9EfOou3CSxGUWIZIJKmJSIAoQ0UFtDo
UdTaDF5S21cBOLoyvnux1rPZaapUjJtN4bPvW7wRA++8by6w5v47f4kXIWd0vvZT
U+Td1kiq8ZYh8D47WkR47gTTDQr/kT1N6IW8UNR3g2jjl0bZ3c/NCvM3+wnO95iV
5l3CHDXUXOBd6/368C7EUy/hc8accAnFZ5YtdUiG7mR9Z695+iFurIDwA62LwL0A
dexXHI/MIG9jPuMOcNmYYCKnKZOBYh87u7qKtH/msHpfFzvF4WC51hnSD8h9Q1ri
x4swxSp+in7xnaHch6EDziNeRscoLNrkZBnvzQp77i0MrbmpzBAUm627HN35aLG2
RpAMdl9wq2ElW9Ksd42biij9qeC5CbIrGQ91EDg2+PjcYXl7E+cOMI6VlJPvBRGJ
5EfXWC72SZpCn+hzgj4Y+6Mbc6xytpPY+L864UcwBiLASznM530WnkjFkaRmQueq
pU0kI4Vt1mYGy3WusUDq4LuuEt3V+4moCfnxtL+RtDhXJRa3jzZxRd6km4JrL7zt
/YosvhInUZoQPwuXyT7o4clqu5vyjNAIOgMSFVPrGCpgfez2nzz2Pd+xMtclL3Su
lcRCaeg/JX0WVRlUjmmTl5PbxfYo+srU2ljzvHfR+uLOyrpiDLBllboCiFVMp+H7
c/nYFZCL4tEgPtbOKAr18+wsn8jo8J5GjINc9QevwKWOTfnl2zb9ve8UOhc9Wb5l
ltYStCM5m0JfJOTOxvOYeu4Sr7s/XERFyRU3T34MF7K0iwDcIOxzzeE2Y8Tch9Yw
Zcp95dQPk90I1KU42gtS6aIna0FG8dWMmn0wdRasGmLL4hFmio4v6tFqkWJt7eE9
VtBcy98nleVTPKoISO0UrNaA0HjBs9qNDQfoH1FjIYLT/IBMGFmc2hhRPqiXWRR3
u1rqPHpjMLeEFqgB1CdbzvtlkyG6JnPjxKDn1Z+VHARus/jwfhyd7ODcHcktwibx
ITUWCkxV0sdEOD2QNz6PrN5sDPA8/fb6P4zbaqdr94Mr8bmaJgkOdaDHQKIpYoEm
CniMjfHnTpKtFep22nUqbQ2G9Ot6ulcOrbuDfbO2mhlD2m2q74tiKUZW358i1TXr
deMt7yiwQWbqRzlZ55Z5C/Udy9BX3FrpZkVpjbuMu07JuRA/OGM0x1Yx9Fw4tFM7
asqy2OMp1sBMwex0W7W9F0ihygDy6lEH4/K0rh7j58Iwsu8tyrL6a5W1VD+k9ovy
iTyGnH84UdxxYsNjXlk+2sa+nH61ShNSC/7qfDBfUm/rf6wnx51kTFG71yvD2jKs
kagrDwky56ZF/h8PMJ3ZzD6NW33SajiKJaG8wl/ct5O4Bep3Y05U805+Q+vE5MOD
cAKt3a+b1wGDzlsHrvwUSeh3sYkPV2GB0KaEpWw9HGM8Vqo5Cw93F0yVH+QIl6zE
/pbNJScc6pRhO3EEWrALhEx/k+7uxWj3YNwd1PRpldQnG7G8AbSHn+sxNPojPyId
mHvYew8tJubITyoebYS9GxUduu0dy9gS+NhY7otPAZfUCk0F4eSLDUW9t8BpdIhi
9mNqwLNcbQautKkwi4ksyk0q4tLf2GFs0oPn/vobXECeScSs86OELKXlALGxxLWA
MC6QWDPLpVf+j7AuurNjISyZIvwNEtRzVDLXetioOR+Y5bc21W7ihZCc09bbImSj
MBzYueu/Z4y8KPM4wQG2SXOEj5etysbdYYWRKX7FOoHLwSKqLjYdl26zEWX7iCX7
OpgVP70Y3i11GZMgwzEspLuWIRcbTJ4myzze2uH8JNfoRNX6esEutX0JN4ubBw9B
F6UQvqsqXb9sC7hqTeSG0LkAEPDRRytVohzbJVD3aMrCQ+ZMpKg5/UkrbSncVYOM
WVV+zRs6wq5t7bT347vUns8+i1XWyPDFyXba5nSDWu6L1B+iYOEgoH00tvZJm60D
V/Q8ShS5oXTj8qjnaN6IV67L+Fqja8s9TUfAm2I5iT9nHWErAHs76rwRma5gey39
HKXzZBeoTojFlx6Hm3+0uSVk/96sAfUlP4tzUd5HhM1krffcjaEpnxK42YjznDVJ
IkbOKWHsH+wiiDq1GKtxDuyPkcGpQ00jhRiNfjxrJ0hnbmYIu5v9IzcBVHWBpXW+
7T8eLcIUiWa6pFhCoVDXlNi2RNl9oILnzj2YRRiaTzl/bjdm68wnsYtONMfU/ct7
vmWGGdoHVG/2VIsCJOyeUSKRXkdlieN9tHrVrbRIv05aqvHx8w4Ia4fvkktWojSq
llTM6uCoHDTHdCwvZmPPcz/2cdts6o5zhs5sHjLvoJobOyCw/N7xdsvFGViig1iW
wkKQvUcM/4FG3K2B07gvbdf5oURT7TB/7fIfDmEz7X5U4GZiomzVF68RBjNAP2JW
qkrOBC7Q5L4gcDD9ELtvwm09g+s9yFh8bVAE0CzDuj+Cmz9Jiw9FquBki/kM6S13
BZuMtrsnTPPLSykAevzMNEECYBKylv76Fiyw2MG7NjDEdRNjeT0vkocKya0L7id7
S6g1esoiSU+0TQM5Q/3d7pX+OrxZo/+6kT3KOAm37rhZEY2/AFQqku4aLa3t/A2R
xUGnsccvb4XkMOHs3s8Khsg6kJlh7er0/VDu/D+u42LhzyViWLiWh2vKx5KXmlFg
7LaimRiTSpM++1y6RbM4bZ0+oI+ipEWFjHgl7EQGTvnzVG2ubggLVQakgpJxk/mx
aLHlijLtS3O+0j4pZDiyAKQZ8UNKKTcq1S2EoixSWVBmFnyDUJKnSSM+GR+l7kWE
MBdd3H2Vwddaa2FLGszzYTbs0aptwPGZWV7pd1bt74xVtyMsUw9T0s4JY5BHNArt
MOq47ARJHILrlidAWZQZys+ObS3TtoYZr0F6jpA+i/iLlpyEM+FYikIxDxiiOwGb
1dr/92KDRQUHEQFUjnsOedxWv+rfQJox86CmXsGi4XZxRtV77vlvoU3kZ8KM3BzB
7xBR1FrVsmdbtfL0mTBbiqevzuLdZc+VzmVQTy53bZL/qOAOW0qAQ/rNh4gJerh+
7xj076EipQoqQobD4kpjYkg1vHkHlcIexMm9DI5/qF1syWA6bvJL8r+QhGt/7jvW
Cna7HlI8bLShmMfT+bEV2XPOVdeIYexvAfFk4UucwngFIbeDi48DvR+MYPin7xMG
XHPARUgNkaQnN2ct7O3JXY7gdpaLVVsfUjsrqdzdHro2JIjH8QTh9jJZvPoANMWX
ych/gW85ctALvXegjkC5XnAU1E43v/ArryA/PLAVlWZydY76bIxq5/Tg+qVRfxgl
SZb9Mc8fgDe554p3xGHWfaIHKH5vPdcIAQ+/wqAr5Ltl8Y9GRumB921T2TeLigs4
brGVGNjSO+EM+u7nxoT0+R57o7EtezNEjNe+wR/vLmlHncQ0fgCF8GS18yK/1ZIi
dPiI80/m8FUh/o1UW1TfexCNT/ZIWlq8IAJzH8ANdguBQFER0uRgk8dK84wyFOcy
x1leEDZGIjeLHrZ2pbQ996uQLpp5f1kDC4u5/KYXRxBKVSBJfoaICQYZOZYj4d+Y
7aYY/rri36fpu2g0D9w18TF1rVcNNfedSuBhql9waxqfpR6fl6EBIRsbylLclpGI
CsLUMnUNQBClpIEAA/MwFnFkWeV7LzrHMlTzHLbz1RysVWTBFKrC+OvJ41mqXDbU
3s+wMrYtNaeubGjmqVpTLycWckOWUMFOI1mMXXeiNAiZPTCKNZxDQAYOZkRNJlXt
L/yba4EkDXwbDRWdZsAMFnx5XcPgS1kG89GuvYPgZjDzlUULp6aqja2GCNQYsOum
zaDeElRG1mK540fW80EQhDL9ypLOP5weHDlO2JZoEBn2V2SlxzPfkXttQ4n9C6im
9LGadcCSmN1I2bskM8xleeISCCtrxgyynHwl98N+FV3lszcEf7fBGmZ4Zps6CQRB
abTVxK0oD/wmcfl/li/whtToRqqozSTc/jOz+88kx8PhKN3m9mo0v2+trroU5JRl
ENId3g8lRKoT8cuDqhO1bnWPJ1ODT4HLXXUEuwUu1qaEkjtSxR1wOYhZvA+LLNZk
g80OO2/SffUtz06kQKYtOZ3s7DeYLR7U4T4m1VPIO3V1XJ1n0oWEO9TxnMJQwIRz
xQ2oJLBYmYnV4OQrg1p5MIOyiPI6FC8moSbvwSA8gvfSMy4RhVuhiH6ybtMnNy2i
HgoGL5zMmuq9IqXOT9bmMNxWlpswZYGHGtbB6ltVhcpt+Y13GdELGvqNmWQnLKto
akb6WjNnf9hkRfi4FMrfhekKaYDPhanknOSc1uO6rZVRDCXX16avLZ7hQI5CeJ7p
ySHmbZsyjF4O7REWxTpE7HAkyV4WM7SFt4Sovfxd/TS8sHtrUbIiDl/rSWHH7+fH
N369SwGb8f9GnfspykT16Ob561QnpQ5iNqLaKsb/z6HWSApaADjy/zj9gwMGhrGr
YT1A+l88orJN/gSKtcnwObMq9Yo+mlPC2NYYk7tgWjXUjGj1f8v6wIYik3QJJfvB
aSy1qH9FEQm6HN6krkNiehoKEkSKHkC20/N0/Uf6TSxNmvzQOwXqCHeQBva1jglM
tSOupUhHOn19hQUQpVgQHBQrTXUxPXoB2BABQDsQE1pOmgE3Z5uvp9LjmOjbS3BE
0VkbdVPXwwYKRYdX0mAtgk5ONz1rsUrympG9So+hgCsMXV7nH6i/bf7p4wW5eLSg
1fu/lCWeHIJE0Oq/wO/huB9TPeyz+wUtDzxqEptNmXG9H2TyVrMCGoqcJehNkRHV
3eq9J76aTW7eu4qlZgSInNUnyV6WMP8PkJPNapDaW0IWEMTNcSMHId4YeQ6wfOFx
P3DsbBHzQ5quob9EpQtkdkeMDIlanDZMSN7O9FQsXYl3PASsHONovsBnpop7AzYM
pdX0NFr3Uh9mcEUiMiNcQK3vf4g8EawPe9QRM2BzHbnqvZAB3LD/yIkruIQLb+1e
PQ4jFPcQiwdGGmdCLqXT/Y3RpIjh3WrpT27bPlIBFqGAe+F9KMykgKHM+3/uBwVw
Zn7iBEX+idfAJ+zEPnuPwVyL8AH7INQWoJ9/rxASJqf8LzLzq0yqpCwNz80+pD9/
YTtIjcIHD/gCstBHfr/E2WIO/kYcsABd1mu2UcTmxZyR4JIiKL2BbHo+aMyqhgEO
UtdP6kK+B3otsiGqWMLjQyvE6onurP3Ma7dhcYIap+ULzRe+miZPOZ39ADOpOr2F
jCnCDnNik8n0FyI1C1sq+MBDC9uCrcQW0TGD5SNXW5qoCRXNcIUUpmk3zCtuTUc+
PtiCRc4h96mRmPZh0r/DGJ71JJ7HrSPCupjV/Bw2D6WY6fC6cQNWGWujK8Rm6kLb
YuFI6XrnbEQR7xxRtrk8MYbNP2l0UJpPzIhosJoI8zh7hK8Z4xOdiRrKrCr+wXKa
K69Q31t0lHKO+F1mdGukSB8pXNEzVrJ4mtUOGCcUygIzNe4oA+20GbwNO3vI50UB
NRK/SQCdfz//N2PXADkA5E+5Zuv3tjT0YVW8H4ne5BTgFrjLRiU+OUfpPlrITwRt
K3+Ypsq9I1F2WPgaawpKYAS4ji+8b6p0bpCw5u1qylmcmy39fgC0sz29ekQoa4Oe
QwBqONA/5Mlu3p09dNTm841MOypA9Ec13jBudpSQJ/SlwOnBFGKvISWq6rSOp6+w
XVga5V+3NG6eDoCmypFcTFT77nqj7SFZm5kMtOCGAzFdepKXk6f5ESCVH45V2JUR
ltPVU3ehP+/vk/dCxfIzdoRdnIbm8GfRyNUpy/5wAelvCMiXbbkBDnGFx7kXyVOJ
IU2kjJNrqYBlhTbt1WQavo8kHg020fBjYJNS4x6lwTkl4+LUNqf7cZzEihszDH48
zTi3hGMQ+rGUYMaSECjjqR9IRVuo2G2G5uCNvxjggi8YRPlME6o6qq/gBSVFvVTx
5bugJP2OlCL3yYX2eAbqnfyqUOAC2XszLxs8iqBMeO95qvCb3je2TGl0QJ99EOX5
OIwgsXCOpPcZJPFrciKv4NAZpuvxqklwT0ezXjv29ehln239sKRnuLMd7Rbjv/hj
ryqwvem4PA2gze2uy8Jz2jya9w5YaOxRU9fcz0L1da28VojPbXGQhgZ1S/E1BYFN
rmBzpnp8baCFZr0OCBAt2A46v3OVFfAB7b9N5U84n1GNY0phjnl3kuSeeIg36z/s
wtounZCSeDoFzPpfuHtGV/gt+Ac2tCc630WTuGMxm6EFesWuY/7OFszJJtdDrhRA
gDv3pvAlx0Tr32bcwyykgCSKND5hwdSn/Q7lmPCy+YTRClDr8o83jSAgLEoji5zs
6147+GisUzoGYvLWccC1MrWcx7Ks10FqPYPjLxeoj3DXJMFgciSSw5ICxUOeng9O
f7hh4e777lbeW9DiQP2DD6FSWmXmVkpwY/Hb9RqUBitbDD2wP2AjmUm54BFnSbA5
vSZ6GlGWHydK5vYcJN2WZcY5j3JpRjkObYMouy6Rp2KrXdw59WyHycy342Gn6zmT
2PQr1cVeZUKJ9yjxR5VhTGMVMaiCQspUZWBLKTvRA778clSEdTvcUHGpW3i0oef5
Nbsyw3PrJ3cYnDOd/mkDcQ2GHIAUpZUqITshbC34diju3pU8hP6RgtyEpLmXJ2et
4RUuVpJQtqiU4TfO+SAZ6+kOoScElIn897xyENo9NoJmI4y72B00YVjQDBT3XvVY
PKlBN/epKFD+RTC97GKzddF82O2TAfnp3g3ItC6y/1lzzWP2Ir03xZbpsB6JNPco
g0DcPp14yy2wDEBR9Ed1nSEys5/Q2eVJozRXgqpHwVHvxW6z3mSE5ge9qmAX6qBz
MmSU21iYRG8AyQVDAxo0MfNsv1aBwF2InhOrD84eqAyki/FrvGvlZyEtJ+ijtDyC
8VtH0B9zHmJp7rdJyB4jMeamQ5y+pPgMQfzM5fIoP9akaIKhawpTA8XgiMDTG3a6
Fz9L0h6nbDDI2LtNTaAhz2EUjvuVZmw5lojCK6jnmwfGlPWfsGqJfsht9pEHBRr9
JwLOe0yRq4ZzOW5GSyepE3eIXEc1ASGyvf3R8Aeud4fkTcvDQbadLDl5gcKrKVvX
hqefW0wan/vXZIahFKNhvOOgWR/XiQaekhrmCU4hRfECciLF5wExs57cYhB9Mq3C
WEN2kkjk1JetsyU0q+QE3rnmrirVz2SS1EHUhg26BFyyGcuWNvSEN5KVX4FDOVUh
E20p1bGVCHlyq7r66SexZ/m3bELnuzYAuwF+ckfI3j4paHY0QzPJTg21WtR8sTgN
fuVqCM2dOtHpAbIndjC585dM/3UQx5018iY85Yu1hTwp0Aaiz6rY+N7iaSj9ic7W
ZJNwXZw4Keo73IOyMnNP1V8q/LMYABV2y+BlQ5gYTS1gK6AE7Nd66RjwKFeUCvya
aFUdEgF9+77OXQOeeBf0Zk9Ajjp1doanK8+G5NU5iBgXHWKi3tf46ZrDR8ParFab
MwL4mNOHEt1dKfh0Ogazl2CXjqbIeqCKYKgD3izBPIgHs+Ys7kUhlvTF5J7kXmic
5R5LttQkCD7CYqaRiXVRdXy5LUs5Jj9qc+l/dfWGpVvr1on2SmueqGeoLI4+DM0w
Q2oMTSywotSocnIX5VGln0PXAjkDbClBxGtE17opCb2EjwGTKwHewU5P/BklyVfB
VGE1knYl4e0LPQaU7g0CC7obT1UfX7Cn4l3RgoA2gKyTsAsbswTda1gxxoJQTt1P
lqQ5tDq+K8IVdleAfDwaeIFDfisNdc+f1v4wiUJenUrtBMdDcCvyx+L6SNkuYYz7
fbcyAD3HXACfd3Q2LTBEY++7fQ4ylmeONKDd/jnFu4NPNILAiI/Lua8JOsc6EAOI
/5doBTtmK6CCUVMJu6KmxX6s9oSH3bIKng9DD9y6qYNLgS2uNmasMgBGdjuVHbRx
sy5SbmswL19poZtTwGvecGa5YWj90QaZtITYKYtEN3Ae7aboDYHfqDv2dmTuhUFl
USk2ig9nfxc+VK19LXHgOM+TODslx6YW3PQi6kCJP92wBnw7HbZh2LGNfoQy6g32
gWrLQZTWfoToIS73EAPX8zaJZMGmb3KJQEcVtZ19zxXLtI0e4wWnMkFT9fZ1CIyv
VvM5Y3cTvBKvTQV3pKn3Ms7dyipIpB/f5K8eiTHwEOHE/fQuMd3BuSQhEQs5q5tZ
7AH2QKhzr9rlLtie5RceVNApIAJQjn4H/ovUsJwonPcWAafiTAhiWlajgoTN947z
zod0icD6oU6tl5hroQiSDAMlJlS99xIoWwRMVZivhhMW3z1jLIxrEIuTUZN3YrsQ
R1L8HgDEKEg5ahbe0VcFpUVOei1emrj2IBik7W2UOeQCkexlu0I7Mi/NhfPGXu08
Q4JjAO1cxWlZTs9D4xpJ1sGln4bu2xwIGKnzmz6kAfnN3o3e8yiwBtQ8HKXqg3X0
BK5CSjOEJvTp11WQgnEda4HVJ4aJWrjzHDkd9KQJ6CFmf9YrAFQzi5ffdC2bloFL
Rlah52gxSAePnH/bDfSAHQ8kvhC/iL4lHC30iH96ilvQZU4GK020WRPFgZXNdry/
JljUejbF9p5fToL0IyichnFEgUH2HX1OH7djovJ/Z7GwrTrgXlCxZ3MNq7olc2V1
waLF+f+NXMj/yRltbOgrJx9C10yuILoq4gODPE+O/KEceDZKzzppI9heNp4ddBgr
d0eUCkiuH4EPCEOZzFXNuX0JK5a6CYM9Rsmy6rxtMgAwWejQjTTXhvbwNDJjCYh4
HYaV93VZw+PnSKYcn0CEohfzFzwM/BTkNX6lg/kEhA2OHRpZxcx4VGkiZFY/i92T
VXglT/avsj+9i/VEfW+V/6BmiTghtq9FR5AEyOprtN4yEmi9S2TsLBABQbocV8xi
HhZlkMRyc3rOgERnJRMWGMKkGXwXIllOtZQKIK+pjEscKkZswxqeqn22DevDU/qY
BDgvVY4kWbhI8z8UvyvcmBg34Mx7VghEt5KkKqeGXLfYpgwHEUYgTsVMWNYOLpqi
T/8E/Dg92Mf6+e6znEdziEr3ZTGkic+X3FeixKFp9OjwOxeTmyW8a/gsMGz4K4qm
mAlrICC4IaayldG+pKUAv0ziHo4i6w24EwYbPuBZDDn7ttuuSlY4X4aJDewIi7Yf
wB3NbWiaWVi4BuoRixbKXMRp+rC96AEh9BewcCzywmjbCFq5Vt7xNsre6FwXa0iE
bNm3aLb78awwilDOkdULR6rsCL4gCix362TRMgM9+RGcBDUYQF7QnS8AmgGalw4p
gq30oZwj+n6jA7NT4A4pYI6uQ8WvQL4iZGbsXoF4Ft350mz8SwCRyDpSaplIF4Jd
re5NccGTaqD6by5wtkUWoyMBx+eyKeyGMAcLnFSkUjjukSp4azz88GOEuNgdYgRO
orqKRmSBpEx9zx20pgeqcTrIF2iTxflsQZkZfaaIj3pCHtA7kgPqc04abJ7kNNRw
7LYTEzOpPWAO8l+IaOlcEL0Q51Q2WEEnImLzyBjC5FpySAtZu8SHCqhWIAhZpyb7
MXQDOlDS3msVgKDSG2m8cvI5PUJ9hZhHRrXNibJ+X8yWJjy/h3fPQCkOwDZf5kxK
obs0hcPEdajLomGjYJUiDiJ7oLW2UEv1PBPnZWDKagVLnQbEzUuqYof/mLhVAuae
Xx3No/48eWBi0D5EYoUWGIW3EWE0I1zNi9GhvdoGKUedV+Oo+3ucVIw6OXZUG2x6
ylvL8FI6+jSTwEKgyLrEKfeim+asMPTjIpmMTsik7+Z7Gj0U3CGfvJgD09abcTab
AcZDuNIR0u3khHF1ug4aj1BjCnfeQcChzrAkkf7yi8ouFgWplxh6Jfg4s/zfLLI+
7TuxEFEbqwWgF7AR0ukzgJqqTUjljKq6tujb9cdb36k+NBxkIjPenFcdM99qMmO4
PVQuFyVFGEt8ghM07HFXBHSRf19K1IqYihF8PnyPFr2UG+jQ3Rc+jkCe0RDiDI6Z
xPRiKijcAEvmmgrVIqaAbGgnayH38HPzUfS9ZYTxb/hMmity4AjPudl6OiM4FGX1
bBPjqRRqXq033ndG2WCvI0WvX+XFbgxTXkeRyVAoGXTJoS13ZVKJ6YJjOZhM95Uk
xvUSYwhEJ2YRkV8+1VDQKRYqjOCTwF2Bo/eeoe0GIF2/Jq3pWuO6pwiPrF2LXA0j
W3zP6FmJBMMBRtvuLWlbxVuI8c/2Bphx56GYiFYVjJVjJ9F+T6PKVUXqHtaCV1Uf
uWKIZ/cDCtY/pnrN/Ycvw0cGGRNUj0mchvt4O3C+X4jTuPuPTNRvGD6t1kDmioes
KR1boOaZruDJ+q1A8LOmJHj/RKFhvCsXfjktCxFs21/qISIV35YIgYIML0k8qVjx
N1D7YSfvpFv+hgMManWkr/lEWaFMJzpeoqpvK1ZX1THr5Km1jTEDvHZBrgzbZXhu
9XvmfK3AK+5WtWDCLOnbcVRy0trY4i2+yztRZTjm9kotF1b+FtWI7V6sxrH0HzaK
HrHIk1pKIyDw/1FogOiTFHBCI2PuVpImx6IrDc8YtROil11dwrn5VylXP8evMjir
ixznm0AGoV9Ak7eWjjtz5GzrcA5pKcWulRxALaqDfDhlXJas4Uc48mOXG37ts5bl
DbHNJN2UCg73ymkV4zcYQ+Jy3551Hy1sARIltiMTZ5BpvN9xOL7fC9xhF5up2YdU
t0L6TLRRsTra5H1UtxE8FZG6j70w1xxcKyuJJebKHZ37tb0R85W8E/kW33nwl3iG
0GQW7jbDiaSm86yN9H3yXcokZ+jrorPJ0jM8GefsBFyByB6jimSkSYNYadx59oaF
SrPXJA+vfYhrkuRv0mXfV1MzT9LPnmehy/nyoc1PyZvxZZC9na+icdKVohb65584
fwjwiKIlrE4YRFrOKzUcDV4l9XbFgIYvMZmmPR3V29CM+iH51KTKggKrCxSeFBLa
HMDgUz7jn0+FBeRGR5qh5bqNEDl/PuGCb2HIarsD8h9hLNgv7zpQNrKwlLypvaVD
Nee5NQUNO5Olagfot7v/7llR6UojYVIj573GAD/Zw12bZT54ckbnnyyXSgAS+lOF
OrOCnOA0vSEINXroMBWS/K5S6CsZ3BARUBYvFw9/5dfMugknRxhpvQKqX3VsxFIr
00kndluwdS/k+aGrDreoJFNSr0zmxnPFY5GX95k4/LIhGGgkvMeurKafmsza+uxB
pixmLIeIBNH+6Vgrf8ylCeR8clQFl1n7VaNkAVcbefl13JJ+Fj0EItc6itaCzCPC
JW2DxU4be1nBNluGkLgRYZbJCmRmfYdjId0Sy3ZsQXGNpeoXwYfpjyLIwkv2HzJV
AcqVatvaClCBKoaD1+mNWZUdrd4NysKwus5l297hSzSp+//kRCrs87+B6D47trDE
c+P1WbL9mGH9uxyW8mAn7OuWrPdT/e73KUJ02FpJpAMerOFzAO+xC/9lbN+JOLXZ
qBd9ssIZzS4UMuu13etCzhiyFrbi327G5VJmFgjjJftIQW+6hLaHvj2nV8b2cjz3
VJWIZd6ySSs7OC9hGOJvncClQFH0gO3Z/hYGBPYTIogo2dI2HjssMMRtZqOaz1ru
QCHGzuIHGMEl9T7RFucxbBzspsXeZFtgUqMdcDPQTJNF0TMWASaxrE4yGi7jrm5y
+IFcmysh6VziUoNYlRPxlj3dfpIp65YJQRaPgAqSp68qMsx6693vIoxKEesKF9qn
l2uDNKUpzUjbOBhRSgG2KFJWk5iTs4Qc11KeYJvegaI7p7I+ogilJhgRUtCPS3u8
J9xHEacj9EfLNPrZY6+82tPdyy952vtGk9+9HufFlppW5gsjCHJEaXjqak/RfVRi
XnRXesonPDFrziMfUXCvF7lvwOBY3R4PvvZJSJtNu9kHV9+sH71nBNhZrMNnfug4
rL2R/tBjXxx2OonP3Inefopx5pkzcXZ6a3KXvsou2OwlUvrYSjoZ3oy6qbyjAZZu
JjrlAH2BttHwnsyQ4IyM4Hb5Ra+g+SIX2xZb2ngp66Nv3Dt6SjRWHqiv7tzDneCs
v7oPx/y0Sh2x3bl3TcsOnfadUKXFCucajM81IBg7ByU49ouZ4woYTGPc08Phpisn
wLoHNc/DA+a+roOodcSus0cDnG1iF4pi1HVX9qWxky2PPnC0qPx+HzFZoG3lvnsD
MI+lYntH3XXZMu6FgQP2QeQU9TAXvXNjk6KHe7Rn7HIoR7UFQAqlzjKaIGQfbOoX
8CF+oLZjndKzSwT1pF4Qu+O9KIQX7d1cbdQ31J2YGIixCQWaeQSOn7Chfi8kBF5E
2aa9o5zwwjrhwV4Cf3KueQqjzNiF9GP9MX4leigDkxLbS3GQPAP/M7uAuH8kj3rd
W2pF3Yb7V5g7jjFWzZiSyVFu6c/KnUQNulC97uVgLLwMuewblHzR7a5IiSJyngdd
x4yg+7olEQBOtmqEKS/Jo9RSc3ytcg2sOsF5GCG2FE/gkBXOnns5OAIxv7XhnOmg
UJPz3xrqIhrMp4uosgdJy0TezWW1d70cMkIWtO4mv9H47qpZF0tMls7s0x+elgyp
vHjzSKCeKLXfekkLUzkFU2ayGizbBB2gA1gCrBj0YDppitizSf36m/aZJxJHxF3h
+qeicfL9/1bs/X/Ogajahs/D75IjSyd1A9Vl5cJg38D2rHFVVbY/qCKX+j7SEfFA
/lqMoWIayoTO4JSHP5I1debAURmmAOWGpLfB2ycBRfhRl0KeChj1bJJ5YUE8pCqq
axUh9W/KG3ebC8fJTJNn3hixhQ55/L+gmxtvvzGpsn2gkWeLzFDm1XopuWNgwAwM
ihdYQ3f4EiphY3i7TywVs3b4FDbEAzM+3MvxS5SBPYEBqzxWZQkCo3qrvZqlavI0
DD4Zmx3o2tpw5MZyA/GSPYVBptM/IJpc78tscvvEm4ELZBMY/l1697pO/WhZsRsF
+rGEXwf/of0zTAJtlIQ0C0r/Q/4/XEf7HWW4gbqUMbC6kkT1/0iJXuT9DwEQEKgy
5HWi2aZEU5XgLwdlpe2O/zMDNCAI/qLoFLdPSUUeeS3YNtSs93r5Q0uWIxHCrxgc
EEtDcU8ZSK0CCA7RcWkbTH43XI1Jgz2tv8kSU/6RX+aDbSp44yG73X3RxcWgkZN1
v4QJbFuqQ5yWzVyTnkYgWHC8QJyjsI5Us+iUhNyDXPOZ+aspb7tQ72RYNawug6gH
KfRaa9q+uVmPwyByLgcfU5bSK5ko8+fgFKt842WXapeR04WWTVDhnZ4r+DBSUrI4
sO4h0LrhMMMhf/2HcHmbgcqt+z6yzjKJ2SWF0vEbzRcamSUJ+1Dk1wMv5qLQWWq1
mbZLCM1KRm5xbtoQ9R27u53Ca30p4a0IAB+aTuS+V1gtIsxtiZiUTcvMfs0KXEHP
E8YxZJAnOJ2SOZTLXnsEjtoPJO9hSrKGI0v5FJtAzljR3k0kZAyfLbkTQ32sfGsU
Xe4lH652J7JY6S2FdcyNST7RZ/H8niP0zeJC6Xf8yL/1Z+LQkMm0WMqmIMhl5/XX
u9hH5eqWkbq8KSqhIGac4/WDjog0ngqsJ/tg1YJOHGQBx+MQ3SLeJ8tl5MnzqAWz
Stgynqe0XE6AShXKzTpcFprzI4DVvGajMRTi6k4IoA8gJBXeWxBKq6Pc4OJ9Zq67
IAbabvOBDeYz5HLtXAewxUs6wReuG5ToF/7S1bRgPyRv6XDaAhB+p8tehxZ+HQF2
jYZNwBg0Ahe777ySn+kIgtOWtvNwp7znsYwrgmpmJeqYquHSdqT4gI23jPMyaIVr
pm/YSUqWJQHIHvtBLSIZmXyMewq1dYKCUY/TDdehWI0ZZB5/WGrPCrkAvpaItGb6
lezqepp3MDEECJ5dztrxtfid6SEKGj6J3T0D9HhNwhOLNZzPgBVTdG2aWboJkGwS
AI368hdUXB66pm/v5wJLNHshfoQsxwd7elm0y4SfgQJsFhyxJ4kSDjUPZPA2dX2A
5Ko2Ny0Q19k+9lb3FOXIvWafpEQFbQm7YrQqjosAImInHTx+iE3dgj5TRyN2vqPU
1FiXZ5qN2HX3Ro3/qITAQSHXCwTGg6wkq/IZ4bbs5L41mgVfzEGvoWEeZbds1/7H
I4uQ3T1oxtAWRpWLVFnGoMAAA2rNLagvHdAPxAoTl4xELNBZwis0/3AmPRHMinw5
NuJQbp5d0D7QSwy8y7hf78Wy1iq+QmPO8yNasAAqq8U63YpXbIOOar01TOwAwcaP
Fl8DADw36wxY+edWDUxtsCbU8kwtTa6VAKjKLGs3RLKmZSazOyjhMwKKAi/ABnjn
LTGh1/6zS53K6KNpnQxT7vHERfQdrGqgrWuuS8NWOFIJkYHe4+7zbkP7X7a7tZsN
A/nZ8t2kD1kFtOaBdgxEEGtJ1Pju/gsmb3M63BXzC6qQ0cwPpCuAAkDjwQqvMC3+
vu062cpQrd3JmK0V8saSD+LUtZuBWXn2uEPJOIvSWSTI4hqm5z0nivC3Qw5g5zJc
CoNIAGodY23Il1DMQv29BXXLDXZVr/FEdQJUQPB7NAISdvXcKfCTcGBL+2GE9J6h
/PKHzPfzzlHAn0CfBu43Vreahl662E+g/km+4wfqdeufjDu/ktLKpSgzaDD0Jh9I
Q3W4H5x8lRRrysg2J3ncCCZAiCGL4hbXcZaivbchyJcG91c8k2nhZnZkS9vEBve0
IirqjhAnPXfZ22hSe2EDAevQsqR3pTXQaTY093RXR1iEMuByzdsNVffTzWW5cz13
69Ey/ZIwxdusu+h/o2COEO7VHKzApL2LmJoT4fr8PCA14aVJdOK0ztOvQzmLBn/x
kk42FuHM6T+b4WiiCUKKSf9Kie0lUJuy3mZW9GNwjoidL6MpwglQizFc9BxZ6TMM
//wjeoN9VT7a9WsYO2BA8rJF9+SxBtq779IY9BgGgJ8thAAIFyOGw2hko8jwoHVy
cBC/iVfNuItKM78Ba6pGZ/8ykbLzGTixs5ppSqShbDsKCosKoG/MEPek4+KgB7sV
fXDVoEJtVHNPdNc7hgBRLfp3W+rLGJveEgO4VZROkvtX0or79RMAVNGXWWBn8hOE
2xZEEBf7wHvglYCp4pmP7pN/+Qu09ukujd/ZXQFyYoyc+EA4CdnpmIT3Ldgj2lJR
z0xiZcZ7ATzrdSMjnKAHn6ESA+tadrkzwgaXXFJvau9bgRy2B2XMaHH5c3lV9PIQ
7DIjoEFo3RRCdc4POxOgv2nI71dRJtUgasy0crxWNtwgyhd2zN/G6CsdfHog/WfX
G12AS5PaBj1IQ2GKYeHptaI4P6l6e5gm11h+1QBvq4VGuMy7pOFLcD8CWqyEr0wH
vFzLd6nH66zP+dsGy/unLXEK1JFWwiYfBoi5Un+wRJUtjxBexJMraeY4Lzn8h3mJ
sYYi05uKVW91MYNUqMb5q6H4FroG/KfdvhXdnqxyBrrzv1n9Vlxt94hGev5Wz1xj
omVtr2XLVC4iVVtYsMsTg74lOkBo5K1SbyWo464bURd5EIdwIKlbB28kmZ3Tg+GJ
vE6G8vaBzW9RAsu2/H2vA9wn1SC6rP5RtUJ/rX8Xi4sA1peJeLMOpcwJG7mqAkHT
H+pqPWKXBAAKcUhEX91s0bEsZpUqBp/TmGB309HzNSqUgdSL5afnR2zbF59Ucrhe
Vd4/y2B0ctl0E1JxhFDz1u86GpWc7NV8604uFh9oqVh0UrGO5evvjz8pOjTKVmya
C0nz3b4M5B0MHK9e38jzDRMbXmzvdFVIpasmliiRwG8aRCBpvHzKINNjJSzCTMxt
Z7AlDWD+dnY1afvX72Y1E7EvUkrff0nOoeAO2HkJ36cKtINQcIkoXMsWyRic3Isa
KHc8wwWcbr9dE1lEc+nQzaPS0iMLKs1xhwXAfS5RdAJySIchw6c3HOkGNCS4O5hl
WNC9kBe3IAZn5P00VMXYW/tQ49tE1lrY3mxk1Unkbv7NzMv6e0TyOzaw3ki2d+KU
4UPgdBwIgl9j73mhiAYVVnUi/x9ctI+uwleZVkYPJu8xiA+iKqFjHHreWtYDYwPj
EkzvtV/Me+Ef9B0AuJyaZd+Rcf0rakgmOerWCvjiEFmFAYSGQpnWJcdls6buNWwB
/qu6ZMn5/VHj34IzjPL4J6nPx/TlAgFkLXHO6vMOoyr3WyzEjaKCuKivCRwd+vOH
pGu4rdoUYOtWS6Ah9lX01pswXANhmqNeuUN5SRFAyKE4Sf/CamvdPlJNBdP19fBD
qZTXw/S81W8cCG/mkHLprQD/D3vWnh0OvCYy3cC7N6Y4sx5oWGdQRdsvGgMnu05E
fIqEkY/AweOZJ5WRfLI292tnlIJsGZuuAMZcmACKD5ovoff+tw+6Uc9BmpIAzc4l
v5xyJgYmQNszL3IREOZWxM5vVGV6kjNXadiU/gU+qleqRX/gIbYeoFJMsourQ7Qe
YcPy/DCZncEiK1BZCYWxxDNgd7q4yR41I6HU3KF2Xq7kThT4U3QOZWnRzwfiwv+h
iSbphbtKwb2oXFn7015tLOHBD7g8J6uzf6dmAAww51MB/ybP3wWekARcVxS1ALZe
0vYERHuqbIakNuXbcPOkzVkmlxVy9Xp2a9/+FhR9n24Rx7j+Ps7kt0WfpT4zwXBF
VbfZ0VatxKIMOr6dlTL/jHF/CiOJs/3mQ6OOGoWYuED6PWwlCwWbStSUqr7T8XvW
7C1L9mK8Gwr9bT2aAitowykSh/Q7GefqAi8WxUeRSYAq3CQzZvVD3ETMaj+JQWTl
T9Jb25wuJsXQIRKGeSvr9lWpZCjvWmkikhc89uCBAUtnT3cem9gnZflDKKgUGwa5
NhoK4uZK8DQ6pwSGVbX6qq0qfKjn+/eYLreYEt6mgg8uAes8j5a6Ld6sHis5yFrp
lx2ZST7NSZ1GJFVuSox7PIJDymB8wkhiSrWAlJZ11UGqw9DQ0VguOrxM3Q+OVGct
eHkyZuCMpuKjBXMnLsmuVQ==
`pragma protect end_protected
