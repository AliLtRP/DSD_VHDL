// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HUcEkBoNLIAiC00rOVofQmmYghLqO/SeFZeZ9PEvFtyFH1s0usUAGcDoPTz2Dwt5
cmhXIoalUha1PhSSkdfgxidNxhXhyPYfa07k512j0TccPdib9E750XSZfB1J3bk2
1fhTKlYqfz66IgbFb70XC574St928pi4wX7M1GglCvs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18768)
BXs/Xx9EWhItBs5UvZZrlyShzBo1ZOByBF0X/hpNi7S889HdRRHBuIasmkfgU9oh
zd+m7YMtsukVLXPTyqHq6dZ36NU5jDSX5PZ+syMc/c9i9MMG0IUI0rHpBH0m3EB4
QYdR+XrP6S21T0NRSwMK+9FF+pJunIoBLGQZ8PQE73MzxkOqfP53aW/wrpY2o6Jo
OeME6aaDAVhYydwnQvuoLLz7C0BYBJpD08SOohQkTwvr/9HIKW+FdEGU6KT7RbbI
kdDt1TX+JgPMOY0bVlU9MjBICJ4Q+x+1SaCWC5sEKrsZEMOVYQYEqIF9PLOXXREJ
k6wv14PJfY9OdmE7+8efrJuf6OZgK7aYswZLAR6xPLhWAGgGmAHQ5wMkExtruEfa
a4tgg65ZeS/8PVPccVo7mk2TH7f+f1bkDDqQqrBceBjpyaALNt755dNvOSt6qidj
V/4j2oDXzerYRv9dtdUCRJTElZYxLXAjLGmYiXkFhvb18VcCWBTfDqznTYDE0+Xc
ugCuctjtgsIdt5OLXucwFKhqxAP/2F0cfz9LT4dU8+AYC6E/6QBgk721x0WUWq/6
HVrIbRWxo6/CPfFtLftqHogv/DuGQPdMN4eMb0CWD/DrszvD7LXFw5whYkX2+siv
3vzzt8PMmVnl8W8FyOyXl/Aih4an/ogBnCE/UaJ/tlY1g2EmITvCnlhYMBo0Mxuh
3nc77iRm86C8kftPwhTKlR1ZCPCKLImtnDtkyHZBVx9UhtVlNAacxWCLPFSxuK9W
6Qk1DzbMx/mgj8hBeLAIZiHJ46sALbF+FnbMl0GomOPTB/MSgFXffWrKn0ZSXrMD
dcPu9rCnLyPEkY9GaNy4Nx8kew7GdkAGN+l2ky9eTu/UaPVbCnb9qdhFEN+libK2
do+OFdzErOZH4QcMYhmu451cwvlfU1mhwz8CR8CJv8ASOAOAGIQn1Lmr+3CcYF9t
iCIpZIkPKYsI/fS/URZX/BfFarJ/66Rl3u/xZSMWjlIM5G8JPAw7/IORgrsfRVQV
YbAWUqRoIw6t2xQFQavJSr1EIpJcVIC3jjgEuqFMxpjT4cYTnZ7dvHpvk7UtEqMT
Ea9y3eQxi4n9/wK/W/LKCsPCjxQD9dT1ECHR3F8F19qTbaJDEt0qiuZiAaWpIveH
DQYo2oN68UQM4hWeJrhvZy3I++DM9KvDtMSWRfkDDRZR1ZU6o09MmQNxh1zlkDBH
1jN3SQym/O3a3mF7JQcd0Y8wbIqD1Cz5270PwKB02VO7CvSNn5ipG5VQ0kU9vQCe
FX1rl35jeTjTmq54n9GsU2mJ2pLdrnqn8nSZpDWIzBnS1fj1K7KUW3tg2AI0JsQ6
Il3n+6Yr/VtEjsYlAFdVaS+WquoGQGFrWMF8vo5Q8PuHj6IlUSeCDyrsSTGSRDQW
k3xf4T5j3O/MNcI6O/kCDffde4X+WIjY0a7uyj6aTbwa8Rvzl03JAVHT2EIS1wju
9XiwJi683A2EJ2mx4dKdl6oCskwL5q+cHXOgxaoklHi0LUEHapD9cmy+SJOEUX3w
7q9LNZ2AZQOwJXPJHHSKIr6c1LAVsch/5BcoWUHJu9Aecao4XcqTMxJpQq2zbuil
+2zcmI/ErBXHMPMpM+TNs4nYeK/QNcoy2smoD49CzNi4N4kUjCJNlJrLhEFz6Uqr
Ef6fWj4CE4sEcsRqde9Bi4UJBEYoTMkgT7Sd8JagDt54tFD7/66G9h0xupN/zdrl
oTWpQ1trRUtOZSEtdpGKohwOUoHk6HpCKk6Y9+BRXS/ac6QFKd091mAoP2xawGXQ
6FcEuTHvG16SLWSXdbc/iAWOCfQizSd29kZ9SwTqQvu2JN9TL/1+nGQy29tMp1LJ
wnRvCIrjmVNJs4qh4wPnFOFZiLwYpbe+qssir1FSSOAw5t+KcwW1cMdh48qHOxgR
XfuR+3Ws7dlojN1QIfS8esgWBTcFscWf2kD6NIiKKq8VewllyMEk96EiAYVJWr8J
WchkNHUErO0AL52bNYT1A1U8vdkqLnErQ3OrBEq1PlujV0wvvMADnPj6k9hTVNx+
u1PvUKzKm0NLkN8x3Ggt2v0NNZkoexgFD0Phu5SLXSqP0V/ahi03j6sxIIP3EEfo
tiy4Dr+6gjv+pXZKB3MB8lApeekIlfCrde+qRMJYYESr72tRmggrbTAVEHqlOs1F
ZRo0O6YPKkVElGw/v9F8+iRzSV3poDNLhDfGNxUk8GLNYci4z6uLOW/BSTxqvVda
ffCzjzvR0JbLaDGYi8uWNsVuIUOs3yAl32to9xCnUtUCEZ1ocDWpjbrB2REYnFPN
tlS6v137nAjY9YVq7V1DwpD4uvFjAUEbyqc9EoJ3cUosJiL/P8LcEhTpsDkDZVkb
85tK4BUYbtQRD3GmFwLYL2Xynh2vvjqvTciVRFMxfYVdFa7tX+QQO59MeLugNmsn
OdM9Tpr7icj6CTa2f8lj5/eoPHxcU7G4LQ9plPqly+w0eljSCKyV1M33pUexBnFl
EJPrlXOlis0wF2gQoqSPTGuvqaroU/+P2vN3ni2pMFwW7SKM4cj8m6i55yPtHfkE
NVv62tXBKeRHzk8qc6pW/7FKu1HQcSMLBCqiSZK4OIW/tifuhzTZgh8hRU2gWooB
ltcRdGBQCqUn7NYKVSf7qkq0c+uvleosWttZWG9u1X2FV9+U6yfTKDwqaiKVx6L7
wUYTEQ7vGE1sGgcRKdrse9Autup+mL7Mq8c47WmufORGKh7Ilk8JKrTVdY79/AiF
pwSTNgoG722jIHzo4whmVPRXDlMlKZtVuW0dl1dOp3/d2T8e96RTrzYFedKb4Nb/
UPJLK3kHhxOmQzUTvmBs4+Cc48GCnZdiKAzDBWB4xLQsCv+OB9MGsydbW5esL9xF
Ef3OegCJu/Z5GLDCYi+S0qu0YKZFryzyY0BcFt2TMOefQvljvmRwcPuhHQXmimpd
jxlMeD62OCzMXdK+uQ+fbw+uKwYjnuOuh0HwXdOW2dadYixSfsLYyQ233U2EL2Vz
ThZhJ8L3F71a+PAYheDld3QefApaT0+0UnGgGVstLvRUl+OS9N4VOomRRPQUs49d
tiG6haYzd7NMTb0CuI+vuat8lnKWHV8OOxYsGwjHXZJN1DCOM/5BlzuTFRI69xOh
v7RewWOKFM9uK7PxpluU4QfxvDRZYMJwBU4GlgI4oCcrHo9G1sDRXShrQUFfq36Z
6U8V7ymkEiZbgjzfIlXtq7VJzQdZEF4t+uWkfuAx2X35KoYsOaNxj2ANT4eguKOL
zVE2UDdHT/f0uRRiwV1lpuV/SOba8ujGIzLVLE4KA0fwlxMLsbsCK5HU509mTuLI
V/A99ePYwRqD6Gwo7SZC2OX2sWXto3GlLuQ9+DLQzYg32NOfVFRIi3D7v+q1TQjz
U0u9er0QxWnj/Gqw/qLyVoWwbgiEU5y67PcvHHuJgvwLFPyor3oG5eDzqrwdMsLy
+ijE6/XErpNMJuoGAWaU3sDF4GBvG/Y/tmQoTR8HiYQpsPy9lGFZSB7qsIDcRe7E
P2xnF39TLPCxNoThRl9HpUDmV96Yaav+i7crUSIFy/DZdRlDe9JdpHpzj86kpPS1
sl6uVSW5Fk3fr/QxE5HyrJ1KNGIlEgODAXsLrTSApNIbRt9GshLwRef2cPIRrBSB
ls1AUDoWBT/30opXc8FUOISPjWiobsPGViaXVsJlNvvH4XM02ODtuje/2xoa1Kcc
816yQso8EUSGxHWYQZeT+ZJ1qjs6h+pFL07y4Qx+H7bZG6tucUCJyWrHy6F9SSc8
vCecN5BfgUAlsnqk2dGfheh6PnolWbrPQR4ryX8layF6XMOJx0rsWPDaQXFwsJ7x
g2sgjW5ChZE/53u5pTzTHW41L3sk+GWHJO01uKUAP3WH7/oj3RQFUH66s1Yl4bGN
KC+NOpVbyQIMZ0mGLqbG8z792Wzixu2tBCelit4WcrpNP0xWEi0pfK8hCA6ybNVi
o07Ky7VV1J6WndP+kLhmSeDFvzLqRLFY8ec6Ox3FOkmaGdSaywdnsjOICBo1C0Kh
H7F9ZMOiq7IyqKQWmFebJQaCPFlWtbd/LbJ1OAW08RBKcCMMrPJ9P9+CKXJmPbje
2geUaHJKTGhUKb6tWOlVmv0QxAkk+XQEKwodieKwt3/KaNq40w4XBdLhVwmtnE/H
u2tAkcen8L1Qhx6zbTCQYsXymkC8VlKkIPk+vLmSsQuZOyQ0g01n8CfTZSFguYIK
rIES8V6uBScK29TGA0bkbH5Nr+XusPKI+n+FccHkxWIGjXe9Pelsad0E2xWx3aq0
K1n/hX4Nw+Zyw5Gxbk40vQCAwPMRsOUMiyFr3ssYTNaibbWHbnCUnOHDnM5NtcMc
QeU5RoEK6nVIs4Z0u3npaQJGdym596SGlDrs9OZI11HhNeby+N0k4cvVrKrKJZPJ
yH2aAQSC8nohjxr+NxqbM6XaQ7E91AbWs7LxPdXoK79EJzJW2z56T2lrZwVw+i+n
8huG+13yV5NmZAS9y7dJerbCvQ7HAL/eWqaJJPWwGqmFrkztV6LOY8RDTEwxFQtT
s+g8fRWQGCKoYzU8QQjhns93fVEz6fwkYdc9WLOBQYknceR02mjMKRxCjplIJubh
KnHCuLihB4F+RlIpMm9NOfDAn1tONCVLAbUJoF0mbAWBsQv3UsrL5uM6J1JQHkLz
dypShv5bnN296nb9XkPu6VsXqyRJvBJsxuegakq1SV3G1cBoYMpJ6Kh+Qn6YaqIr
nwUiGurt9iDbQSP2DTRHeiZKXAS4ULsJOknUm32RIni0yyXjVQKyi7ng3V6MHSEx
m+YuZAn2WIIrZUPX7XLUhANhUPWwtUU3xvPR+3t0pOZeba2STWPVH82r2nxoEEFm
cW3T7ZQ+D382aGYJeqCH/57+iCE5my/7fhgOWl5Wfy23mPavP6kvj30Mp0bB+foD
nwi2sU9pEdPrZcZDpddoBWrlGxFd8oqrD4HROI1B5GJwT8vXoqSqW2wPirVPcpmR
fsDXP/MqZFdy8qrmc3duUm4C8NKSCEthAy8l5bPkiXNGcqKdw4Ioiz5tRmamZCP9
hGM4wXW/V/cXppmjVkRNa0LjonCB+ubeH0DlfJUmwlA6Xtn/hGpnWzePtJVgWBMU
x95hlOctfh2nDqrfpMHd8/MHHASC5cBQI6prHwD+vlpz4h9RemF3SJs8kwf4VEtP
Edr8+obqUdDDQMmJK31c5KlFJB+LVnMHqLQjh1emsZdCVmZVB9QUu4/bth9Kda5p
XoncPxtziagh+YWraVvqHMYlxLT4VgzyaKYuqM9gQRDgDfuNpA6ds7aidtsMcrB1
BjUCja0NfYpjbmpBSaMRX4n83/wqleSZThgpvNjdGAEufGlPM0MAhNva22iv6egv
2onA2GX1BP2kqWW3mRVKkVZxOD+yb1Zjd+aKJGlIQKdR/3c0LQ5rUmD/oDLaF3yG
YETKBQ4BxARq0Jcw1fF3OMFK3S5XEk49X/LF7iPzwce8GNo3ns8ASWrwB67DHw8w
biMKlXenq1RDL0sXgC70v9zNBsRU0+1JHWoLdJp3ahgtNoily3pZXJPEeP4yXSss
ctIZ68uoPtIrDOX//Fb4/q8ix1j59YsQ9JDlmG1Ny9yghw1RXzOdHoCN12pTsJjg
2VDDncndjZ3mtxN0UNzJGY7ptlRyfjI7RRtIbU2aSbIaCZS8je9cD8NxSl1Kta50
eujxue5EzWEYNsQzqfSasiAOtrExFitBN+JrF5XgtJuSQIVQOHhfRshGTk4TGfBJ
xPLdBkylKtXMha3BPKo5jlyojGBMVeetUOg7CUjuKVjok0B22TjYT6XGfgWfdC+n
U/KGokQHhjmPRAedxdoEGFmZ5c0rOo0OXnQPybv0GQ0PXGFVg9YRInmY0ZrsXt1j
exsIiAj4N+OlhefdTpx+RVtysz0A2YB+nJIPdSHwXyRq8xhGK7RXf50skom90rkc
E43WbCIk7IiYjq8FElQB0WAnP2CpJSCZAe+u0uE/+SVvU3ohu8GK8FE4DownhTla
zqwCyBKe0DS2Tj6g3pFM6KbsHwlI5yvAN2f2FtdrDBWBdv+FnxwZV/km4Be4Jwg6
vA8SYASgn+gRJPya9l9eB22CI0R1ObdRB9RJ58uk+cyExutE8wnJBgIWy78ONrGm
vWgPIGV1BfXBm8OwO5e017z26Jms8+LFFOfwZsZX37jQGNCivdk2ss8X43cQkF01
NMiq+w1teqGs21Y3aN7GXcdC6KBLFmyQt+9H0HSIV/oKwEQQUpF0N0tyUsKA9dcY
MwQY0TUEXWRymD9FrIZsnbFLOYoE+CXZrGc9fo/D+sQFKOFLwCo825QPFVURqluf
RNUF/SVqbqvKl/NPa/R73cZI582Nwp/U3eCrmDw24YZ30QpLmdFNfApyKJCxpOXz
0P/HCQVHF6V88K6OCRbXAHDGboNHih9D6U4WsuVhxd15/+z6vN/+TnHz7h5hyaHn
qhgBDOBaJ/DwxwcVULcXpd1rog9BtvxsrZFfb1KedK2e4So+mXBDlevJ+nGjKzui
CXu9e+AKDgfHrcgZoZ5sgLoyWuLQQoX+I6W9gU8miDKcUbtIQJIGophBhRFl48g/
6ZM5jknS4R0tB/t53U10WQathgclw0N0iSCusPFXAdhG3KeXQwAfi/KthGSel658
1LeviSk/PEVKfbuBzkZR7OyCVuLZH8VrKvan+VWLI/56VN27IqyotOC3mQQHo7lw
XQrPSU6vBqRM2/I4urv1MjLtXbe68aasXm/iBrynP6ZcoYlkDvDHhf9JJcEUqafw
TsCMpNQOMiULviu01O2ZEdfE/M85jc6rRmvlRTm45iEZxHE6dn8gasbxX7IqQQfa
UrChme2cjhskbkWZJKFJxRo711lSVxb9Rs2FbgnfyAmIzn/5b7wDKiG9PUKsQwDZ
Ttq7tWcFeUK/16ebXQkjOcLXE8SfkABQoYBJ3hkxB7sf8KVhwaOePK4V4AOgU7ky
6G36UfIMSIy0rl2Ysy0hNQL2VRK3z2pHmql3h1Hz2B+6kce+JtcbUSSQqctGMXwg
eXuzyCdwfp+s7g/Lo8tlsbET/LQPNWOwoq9M0rniFiztNfppwAstL7nkwtNW4r/4
z6Hqc7fhQLZtljRSIbF68gQmEESbR3jPhB06eapsnmk8Q09v8WeS6IpQBp+ihseo
/rgy7R/zd6ZgQak/q4hT0W/mMhcHdCKq+KqoaywJfr8YpZ5pm3JIu2spT3t7vFgQ
fVMDM68WMBMsyEj/J2pEhDiUR3TaF4JtOxJYXou7QQ3An2KrA6bxW9lWC6fZzHy5
r9E5PfXJZ3QYDxdKsi+BHcnBVMUQughZ0Fv/OlJKCBMMIkQpG9J5yRavEGgH8fus
nndC0uru0hRppe2xUmIwGNBVxKF0rMLo1x4SOsAab9SyF7+p8Q9XZaLOmY0HTH2G
PPX0TmnV5Jt1Cy/A2KRupvx88lVSPjJ0yKmhZaQRL2TuVQJyEUG/JMbGLFuQ0rm2
yRC8QJvpy06HCyX7cj29+RwlTDiWoYC3kz9b7oBans5JttiFRN2wDSn8Xtv60ihx
d4qFPR1hOdjjVxzZPFIRm2VhmhSbut6YakHzG+yimlsf+tYFo05khle1igG0GQQs
g2z81KH82QzsBbfx9zwJW5D6SMfyE53auVCqCpEAG5uIAYmioJV9Wn72z/xMQZCq
y/pETnvdO9J6iUKUw7bcyjAxsbFXklwoG5UYgN9q5DCM1ixw9rpTVOsF2z3PatTI
zTf6QptS2CoEI6dVnBtf5sCr2+lWq0X8Qd2InlUAMbro1i7hCCAvtbz83NwMHXNe
CMicn2JVhvEKjm5yG5IdBx8rnoH2b5OHSrByyxr0F7CZQFPJvKNWJ9U3OZ/gO7u2
kSuOKj3bKpQbySlqZZuXMTyQZkqRnzK9uOpA8MdAcKZx1MjBciXUbYmt/qGissru
onbJPw3fbmcYJYwIAvdx8sP9c3KDzXCxmkfz+BtTB7J1ACCvnL+TLoDkd3huYA4G
K9iFlb7mm0QLym8o2ShNiPwLY0jHNFsqAT/h+Ifl4un+5L6u5jWHd9zrGiYoY6Sf
J6s5rbLqe8TPgiHW0ttcR1s0UUXf5jHL9w13ncYd9PxIIf0dQ2t7mIJW5y4cIrfc
/wYyBLIF2OIcIyLSLgMCj4WzMDBDw41rnKaU5SE8fwfeMe9lunlMmC1jh+y9ca5O
88wwfwyp+FYZFqvxkfU/LRGeb0nRXn6JOYarS8mX5yfX93KGMNjJmym5gQqjDQIE
ilAzWVNFSAs8T63+LozxM3U9tmOMHxcZU+D7JDkjGP/ak8mERR3+KYWrqBIo7uR9
fQOHlTqNBad8XM8hwO7+hv3IyEa19EWJWDxUGAMzVoup5AF3ZLkEvnnXu9EuTwCM
Rh4jHtg0aoqSZyzuG+BhiTFl9Vp5WtK8YoWxhOfSXpeSjmW/3ZvaKdeHDQjTNyiT
ejK07uQlmd1gEZkJycLPCgYMH84owPNi74BpiKxOkjNnrXfcf7gabvGoYmubv0mr
kHQSQ10Sw2c515wbdkw1bkTWL7xy3v4ImOlEUZfd8M/tr6Idrk3vJynZho64/0vD
gbc89HhsSbDW9L1ClV6JNlBg1IWHGgvOOvxtC7B77E/0uKjFyR+p1vmyQaEKeQmv
xgej4EXzXx+8cmEfO16ndouxccT84RPtwYbQviofAJCvvmUssciAPtW+FAWEIqjN
AI4fked5Cky12uVO4tTUn6IGonrMHOXGS+61M4Z5kvKmWccjQlCUkIpaH6S5Fy6C
GWALB7ceAsr7DceRBv0uy2EL0wiTrYs6IeR3TaiG5h8AvzjEqpm6xKRgwW9f9kD3
I+3qSu4+QpmxcUImpjr+MPfUbDonLH9LHtSeZErWsfcOaxbS0qnqcOI+YuFgfZ5C
E3vmEGXe5AEtLGKI9ow7wvkv4Ns4e+nfbesXwA/No0t+Ni56NKRICZebiP1y0gE1
0MkrD9ikEFIfsVRYLmsaHSH/regLOJKlLc+kgFlCRUaDZrnLfw77sVTe4OyxOYIy
33UxGipS6zX9AZErhXzZeOkriE9H/k8wDiVCXz0arzekoXOr7LECLgXb+YF5vlIb
83Yfrku6nQAz7hD0b48X2HyzuNpMJhSUWEm8/evo4RCEi4wtTyemEe4Xe4J4F/OO
8o/O9LhV3KeR1PT+LQmsN8LQ5/CLP1cw+FtPVQxQy0la7/NHJTMvqpXOPjM3+LBQ
LFi1glrv81XjjZl8CNVRBPBfNRPEPmRgJiaAS/DM+wVw0Xc2IUdPDcYFuhUxGe6N
+1AglUmw4601gvPodue8reUaq1tuaPUbZNLBvIuP2oF/LswkOw7J6/atJQYbXBmt
6C9sn2BTsRlXgffSz12I4ubgFFGDPNYcbPFd/1bGWHTfp1fc/lVnY27h8Ruj2W9q
XD4Xj3gjyYr5WQAN3c7DbUKX3XZkFtO/odoDJTs7UdJpM+SrkmIMVmuLNH2GOlU1
hwZq3L2MMmWPZps0fSjY/FVv38uoVOkntYO3Zx08jXh4ugxboP/yQGcFFpb89vp3
0jmHKLMBhSpQIaHCd6WN6UAXFig5RqN/UsRRN8bxvdJaWwrc3gyCEZHxVpm3I6iI
nX/mFhDQAvnFeazqEPW+o0nOWvZ0H5oZQFYefM52Q1DUuCW3RsktoJ+9Bpatt5G8
UCX+9oaFvPZXY9d5xuCjtYCowCXQ6iqA5ODwO0hFgkadzyOXHInTdDaFQHg8Il6B
eIMe+LB/1amF9ifyb1v7TRTVqexN6lO9DY0GBk0Xga19cPhvRRKUywnUcvPR42c7
qwcYceivdajBCzqvdoHnlxXMo1L78Zag2Ivm2Czpbw4s4SLWpH/x7f/JztBE46WS
WbqMFKP7T9P0Vi0/QadQm49knjYPG0pIdnYsgBH3Ftc6hJmWhQfyzOXLtakTY+Mv
MN4UbTfzai8JdAUgfVMpdKOTAmSIj5sFFVdvGErq9P5H1R+hbwOf/RpIZ25d/0YU
W3dzPYsIEx77N0BrcfkGLcMHcoCg2RS1v9bVhcQaWXjBl06I8jhAepRfUGidETBy
g2prxngAtm65LWLumzG1tramo0kVzrxlM3Kpp6RJl504oN+6YmGxkwNLMoTG1mJb
YPkocscgkZMN0Dlc4yXIhpSL2+mtwxV5RVy9RqeuTMloS3FoS2a9mQ0aODOgriwh
ug2eo8bknxnMyaedw1kW/tH4KlAq2yhVAFKBxAjzQxLDJRAN1qCEpjbPTuK05Dt4
Z3MS4V5NS8WYHm1TDOOfHTIaQbVHns0Hpq/9wkENGfqG1lr2o4yufnKz8ofdnyvS
9mbkoOoKp/PGNiZgIuZ50usGQBAX+zWxCMxiMWdSg2grXQT3uvJnS3TKKncqkeMN
FeSs5PvNyM3DcnvYiI4VXOaso6OZ4n3P9LA9fxI0buimHSL4udF7DPIRstLmHHXf
WlxzRbzmXoGToPTWx946FGioUVIPhoOQ4HNZ7BUqO3vD6NRINYtbXceBRh5etel1
65lLGsU+/Fyiao/3fKdrx99lbDw2V2LPAUUyS/udQQYP7egJz/rXDTINgos1TEno
RoB+DQNTueff5yNJABgMlq3C4dh5JalkYXB+8c9UfrZLEOc3VIoeLIv9pT0+y5Xm
lYlG56/XTgsPYfEerxTMPdkejguqX/PkGc8+dMaUELbyKuAasnS/2aGTXCttMYnz
mMYhPT7qQncJPJ+omia2Sy7o6TTDRs7gMDkQogwpadqwZ/YHwWWsWRfbiHH2EVN5
b6SUyo1U9CwSwCB6642sUM1UvyM3yO60TX7qFs1fpmKq4i/kzDPWMFU1BdW3heSp
liCZZVD6kU3sX6WlU+3xakP15Tvab4QaQ5Job1wL12X8orBC8ZeY1xJBT09M//z1
nrLBdOPBXalY8WclYXGbsUkjnj7kssZjFzeW/sqJek+7r3scCWGonNIIAk22Iqlb
tOEseV4UDIF5psxfo0QS+eb9kYxUAZUXK/GHL10zdc2aTnFTGqIQqe/iqndM6TCA
BA1GZ2J3N6MZEP4WtPk77WVeczUqqPZ2Ml4BHw8C+d+B/DP0mwGrlY/zAbBaUF/J
H9bgQligFQqm8RiqPlgjlkDX+6l1lF0rDYvK5s76a6sNhqLyUTi9Bfh0ssTCD5FS
ck6GlUaH0mg633jTdnkUjFK2wEU6Zn+qB9taw6CSM0LF0AB6dyzFrv6cJU120h1Q
gPtm9zToIjEL5bDV2bvPJGSepctZLhOEJVAiSlNisQQVA8/3jKt8OAJ2z8j0pfCc
z46U/s7kpfxYXo6iP+2iK07PeY1JrZwR6Pek4ov7XWzPiaEvUmrn5FveywKbqoRo
HJ8UwKoCkPHvWOn546JnqJlHEmaU2St2OLCEQXHOY0yBKG7NXUpiqSfEWhMdlG8y
fFnu1ZkxDxQ+N6L4VO8RyCfLhRv40IZuXj0WN4ni2ZrRz9Aadwkgnw2V98NhECM8
6HoBHMmNwW+52JF6MqTqWI8hIUJ2F8Cn649xKVDR7StFPj0INbwawE2Av0WL4rzo
n5WT3XGO6MzzfLa3+pqFafrZLzssYa/8yi8K47k9YdGWgBRJXxs0zmWzG2EagY48
OFAKZITdA5JDY5gvplLF/4t+5l5sq11IgInvgIG6QuRZ6kx8yHgbCuiMxnqIAUOC
9p7G8eGTS1rBG1BiNIZvBAHdt2DyCVRDT23JlDFnEyuvuKlgx8hESUJGAXOqn2O8
C7I9IrCXmoUDg4LQz7P1AntUwsTzDFU6faAt7wHB5BzHnALkrKCCeyBUsZ7kUbW+
BUe7pDZd8yqk7zZBK4QQq855unN0W2Ox4MARsJ5QvXYPxoXA4nUIsYPB12S9pYlS
emXnpGlR+F2tZuQKrl2TIelHjtScjvaGbl5fK37FpST5sIR2/iw0Qdqcgln0Oy7P
09CTVip4m8Iglw2kdV+bLhaP0LM+KcuTmn1mZCPcFwsoOdpachB676BHjjWPzm/L
ZQTju0VHjlhiS4BmqsuXhH4oxXBQ2H5dmDpMa6fPhritXt9Sc3BJoYGNc6seyJrg
xnGqjrr4FfmfEEJEBTymCwZMY88L3kLcfcb1cjPQeZhjboKVBYOK1J3iAv3y9dOE
8MReHcyXEJiN2z+BkMen5nXa+PtGMxfTF40dqYHT1TQURzOf+xaxt8OXMNPnmu2Y
F0WL/tvzEL8bWv2ThamGgtDhNtYek94QKoxK5P//10dMB1NJTaxaM3FKIRjIJ8f+
KJB6nouUHDsPBXQpRVFdewwimaY2uJyhLj06cyff91L48rN1OdgcwVBWykHzsLz9
D9QXpUmsl91P6Ct6f7ChV4Fvj78MCmi3OlDdOABdPww3XlD/mlvsPo5W1ikugm7c
G6+cT+mcNGvVrX29C0VfLDdtLFzq6s6t7jUYscrK0t91H9/Q6Lg31S0IPLu5yTHL
lChY6O+RIuDhobcOuHx7hLGXkJukSbJdH/wT7DpivrXq5aIZwk9v6wI2FVj+4CqM
lvWSYbIuphHKNwy7s+pfLnPzIsCseFfP4ppK+WdvGJVzaPpDsvHb/riaY+tAMD6s
Ls0bFyD1mOGKpdvPmd30iYrYe9oJEWypXZbLsJcdkMd1NqsfphWmqLkPwSxFfmRl
teicanjxk+M16SNdFOGaXjYvgFCwx6o9Hc+PLrvYJESyQK8M6gdELfg7qaWbF7cM
7MNYUTpcBpRlZafTpnxzqqHT8YOjB1AjRaPjmU+hrPlIkZkltZ91bOUEcpTfJVFb
5mCjYvwmwNVrW4NjIXq/rm6Ky/7AEJOB9TZiMKs3/DUsE3h6Sjq4YJ3s4olPImse
pHij94AhAtUqL3fAR8ebb92O7YeVrjY192TBury3vlUe7RPcSURGiWZWRsjODwZa
+Vu6rh7AoIwFxBkqwUgbU0eV/wOo0aFt/RQzV8UGYcSqN2lSrG4X1bZQH58GDC0n
pzktjY5zwJ8c/AH22qy+Q9koATI+yw6uS/dN4zTQVhHGRTvHgkZuu8QwGPzRZQfF
w29WWHc/QRLdbwK6A3eFULbi+KYOF2v7aycEt2kJ/O71PdB9JzVcJxsOdtE34KSC
edsIwLeOqJJnmu9Zdxp9ENxUDqRrZa4ZesYePndjA/xh2lpj/QSOrgQAcK44X0LR
chScaBl5scqX0M3cwcV+Flk+Sz5q8Lyh7KCs6mGiC6AKfycDS8aZLKoZa/lhC/Ki
AUAZK831nHQakelBY9dMJoqu9GSDiLewCau4CrIchqZEdfJV6kXAKxC4IkbRthPl
rIq4hVR9HOMWAK0ksQt6PAnZyHzwy0RrMIZ3T1o7AnnT/+02w0Pl2KeogTqOuMP9
SzYzVaUWD+25OBMoJBjB0nY+op9nR1ly3bDdLFBIO4U2xpAJklRXt5bswbTd+ID4
EL2ow4g3c4etrHPuCqbT8gKL6WMEeEDKiKrTB70mG5HPKPwx+HLciOezZou5ZhjQ
GSlRAGyc7gWFe3Hvej4cwnymmVmza8xqiWFUQb7g7jSM3qx0VfwgWw7A6UKY7rGY
GL54f1y3S5oj+MvcnRnbMTbeESIrla6ktAmT+7FJGiKgMq8wkoaqJMwp/xMbn08c
0LnIOSZYRbCahGHN8w8cf7R1PBFgcWw3Y5tv42LdYxwAgBun8IPPs+AAqMeDc/g1
ctlnfL6vU0VnzqjU3s4m+YaxXopBxxkjHvOIBMGdl4aER5f8Sccvs2bVj+iu6/OF
6uGcO7N9zATvaFFrFuLdtzDKS1bLwtCTQwDvSkYCmZybbQsy3rQuo8/gljeKnOcV
aUykGLPATrBRgck4YxIX0U1h5eKa0lIOYr3y2f6dmFHYaLP9ty8WIcBy8nLwtpDq
2gq2k4kNBMOZFu8bNVkxGAg0dKdG+MhhUqBgl54W7KwB43IzUeU9XpPFyuB8hYqy
be7k/3r9ma4tWqJfwNcb75p74k/15kcpEJQbeWnCV4OAvBHmKK/T0VHbdqSWi9xA
rhtPkvUYfl6SftCglHQ8hp06KNlaE0zfFYjGUrPawvHYZAZJq6TjBS+DnVEe0OVp
bsTD1m1/ppTv0Znvj2FCrb9uMJ8u1uOW2bUsNpWEqQEL0xkE5uV6xbyKxTDAfFG3
f8ZTb02Xu8+ehVhqDlFkdCTYe3N2RzeGxzH8l7NPxbi6mh9iu9zm9iRFCaKI5ydc
aC4QgZMXKSpDW5cw/gXDBI6BBKNa47yUKYdVl5qXhcDpij+O0oAKvd7f0ZPa+iIB
qS5q48IMKlu3kYZxQB3R7KRMrwFv87Y/q7aVsxs4e4+r/bVmx4ssIo6C4xrirvF6
0anXzDieQadUVKzb9Sc6yV5lcNJzee9pl29FWqV3z1rqGLLaYHnRjA49ph12oeD0
WyTSc7kerFqRwrHNC+B0x3LaTL2GH1hauiNtfdbhYP/2gZiO2eLRyJsckuDiOk0C
nlE8SxrHOkzGD7+G7/MVZgmUGhGQpuBNfv1PpG5BtY1RW07b33k2hZdVDjQ2zrHC
4Fe3lISTfETrAt+KihGchx4DX2CVeyA+O8RXQvnutgD0tPpqFvGdZVE/F0qbpGHh
7iwxgSNGKBsS7VPhySS/eVoTG92W9btl4TAyerU4CD6aZha9l6Dus3XD0sEVUouU
TaoC1jXGF5RB04k8xuVhzgR0/nQXkT50tpolLmN0jW541X7c5Vysn/ImzNZRDnnf
a2nsLKKuUXYY5+miH8VHtc1Vb3rMYWybgDE2yVzdwNR2YWaxE89MioXTLihrJrg+
Yw11YNLvSeyF5vdnJAxef9rVMUkpo3w8aFGaL4IBGovRsnWz9bjEL7nes4juvEQE
ZOl6WzinRS+YtGEmXfDngbghPi762E5GyLWBJi+t3Ke2VywlFDt9oJgp53Azjsr3
fBGz70lLTpqJZeWsAs3b3JlxHf5sqJFr6uMdHzcUlQGDv4FfQ+NhdsH69IMeOg9D
lZDlom1gsSsIwiMVo/9stmrKEt5UQ1Rp5vo2yx0z14jRyOrcjbGmqzQhLpeReQXI
6HCdeeNs1aMSCfC0xltrtyLBQkiP5eEm5iUNVvUkGmiIPpCWlszUR7hPEspdhZFI
vscJhRXn5oBV9OaUQzO9ZXrykfMZupj7wXO6VeH5oxUTxhzqEKIkZJgXyXoWGfub
A/hvvTKG3nPCsskjq2rjgwsRQa8zZ8QkqHrGVwqJw+k3hf9EzyoRSou+dRr5LW68
g7owIpRvaXIAfwDEgI/j0jyQ1prJI6AsYd+8Mqeo8daEq6PmK9Gw04uC1L9Ax3an
Fh/zAfmIg+dlAlg3gyhCUe20/slCb2qhwzfk7B+z1hbP/Y9YY2kDtBtkTXnlvw9b
WRSctQFbGeo8eUcrYGksrMe7C2Pd2834Td0/7pdb8U7TZwYrIAOkw2Mvgj9d7/Py
pD61QQ5boVT05eJgariYcPZUhOyRG6qT/SKosT/1bpTPveG6CEgmaCF6f6W/lHzd
BpjuuTF3oHIcLZNibNU4lqFlMrLlxiVo3/20jvzu2eZnOSFGrWN6Ts+hwuS915FX
M0rHAwhb1aFKsLUDB6K9Acyt2IG6XcLtWnnjBcB+J5TL1ox5Cz2+AKxaGtj6s2k3
69qd8g5m94byv80asXkKMuG3W4mVazCbw7QFznRWWbe9gX6efKGUMikXTFNn4xip
vfuMocUtxmu2UR9FpyNY4Ao/VSGCB/ZZPy68DczshZGcz4xX35Vty6pi27bXc45K
42LqIHGMLX2xnxHpf5t9dJE0BqspzsY0KBoosHtQsR3zEMX8bYRghew/0JIazB5C
K3kqL4HmkkTjJGUUbgFzlRxFnsMYGcpQKRxF2XMQOl26L4nUQkcgujdsk5tQHkyZ
wYsQCCs9leSBaY9A/y+nulxqeZ9kAV2Ul350f2aofkEAhMscbTD1Z9/yFods5Npg
aRwb+wyzKQhI3LRK5muprJZqxgPftk9QWbhjVcyUkrkKxaa+NJbOpMR4oy1qG2C/
MO0erKRKa9cjUYWr5pdvU7UaDVm4cbJkh0AYbq9pV9QYSQKtFkADBcWXrSlQukz6
/hm5mt7n6tHLTvjEVti1AFP4sBnqLI6Rz5sDv6N6KLScWOLlkG4YJeQAfC8U7xVs
5wWnMEchkJsDSqr6CxyI2ynDxfQUaMJTWR8XElJBZeAvjoBbu4pRgjRhHJAZadQy
suitVvIIAL03is1G/aD4k6jI22nZWdeGm46HNWD0PIyeqELn0hi4cQIs1n67vrHX
xDBKSfCrWmsIwDOQAUT8m/ckGh+jwTqwhb7aMg0V1m0wNIXb5XwO4txLNh7NsyFI
wjr1Y09vUgrWdyRaZIATgXLVC45own9w2tEXpOnEobfuSEBrgd11pf/94eO7aBXL
nOE6X4IMn9TR8xXOA9yzHvftpoKGTQeY1STwWnrVzvXTs6votS+13sn9+fe0fYlC
T0lJz3VDtgNFl071KM/6ZHNoqJ5rdBfNfhePXQN9sus1bYmUQj1D1z79gsRJasR/
7i8PbsyVeYbCVEWNcyzuAt+Jyce82cMtQ3Xg12MXtuvvQfAIzYErxJSioe/Ru4Zr
8Oj5XkyQySg4Kdq+3bWHBoXSavFh9ogpvrxjW3i8Nox+EQIYlcoHtu8PXd2jKNWX
XrtvTy84YQywrQFJLhOpcHqusO6C0rnKWr+QjvuIBRYb+GTEdd9SoU7uK4F+Jyfh
Zqz3H2L8dBhU5CDwtK8yUGetGi1Z0GmlD6CaUSfy0SHm90CNts3ffP632tY/hWtU
E/p76N9ekKNTsrP5FI83LR22WVAU7+cfETW/1NJc1npYQx/pzeDKu6unoczBg1vu
i7+/9h8bkPsEJXKnR0lQe0UJ+zLcNunmYMhTMo7zXQ7nS1eag5Ib8BdMMiIWZaug
XGM08nyfYeQSmfKV79B4vrAvSZLa9otwxJI635l4QbhSV/30VSZJ5YXBXaqSP6Ur
056XN+yeOPTh4vbOgYfHJ1qb2wQuB48iUl+G2nW3wQEJ/o9p8dQJrA9/XLTGVZL1
CHKIHlWJ/US3LCPKQgDHgPAOj7Iewb4wrQiM7qUo7+lmhEdiKxQAOVKZW1reOLYy
2UxjmJHzioLI6C/hXSqCWnt3oYhFvmp8U53UmnbnjOhs1Q+8PP8tXcsNUMAvh4qO
9nqmlD2dHWX7UWw6b+cmkNCaUql1Ls2RCCaXpq4iE9aFKgpeVmiTOVz6plkFDuhI
7kFxYxIi6vJovoCpsKaqbwSJzrIFHqmhW58TdOEle6UedUyiy1iyddUh2Vkvwut/
sRNVpgEh8lsZn5tuK2AGd5DmWekGzrn/akphp/jks+guE2C4cPO8y8rebhlKyDYl
5w4ZEFWnGSCdZjd45t7BAXxvLZfpBltKxKUFSCG+hg9lsmKl7yOHKODYNOvOWKjs
ZK75tJDDnCBW9ru2YZpgGnXrAdd0dths92ZdSstDOi0f/CS3v5V3PvRiykxNOLPR
VrUDknBbKt7fXkEwlT0pNR96gWsm/6DDVWpuv2D38pgBEyLHKEB3eNjxVkihw4dE
s26qDV8ir1dsBEd87z840nwOAEyE8hVt8QVl7pJRaEYFS5WS+xTmxAS+N5TyIDCR
C5Y+fw//gKi9SvPHhVJxN/7h/v4tDOriM8NPPC8ceAguscCn2HDxLlGG3UfSzHou
kH9I1ejFf9un/1bPY6LJsOJ6uDfGK3FpbRITxofRh7qRq6OcEcippTMj7QSswQiM
D4gnQgM2Q42Nb2Q5rRlBV29MGTTmiAQsEn3nGYEPlvSJLdEmFsUDqwnvnJMkE18Z
oNQh7XSdi021L9N2Mg0T7QpWcoLilZGg3jlMlUIgNI4Ozpd/wfeBwhwDVe2X7tB3
d35cVlKNle5scsueoFhD4qCLMW6weUYTyeWRnZSw3Mq8BrKBmaauWkirOR2mlrWo
tlAGff2tLuuJ+HX3KX0vWjQs+13fWSgWJM66GV9+jOGrD+m8zBuQoVjFqq3wNFAg
SsTtQEKkz6F4zjFVeMzfbRiS6h7SewilLXW0vQ8I1/FGhJnWKMw2iBwyeUFjnqw6
F1Qr1BunpyKrvNrGDk0nV3kzj+FogLfrDWtSw0Zj4C6ECQ0PztBebHfSriWIEIws
Mrmh858KopKE/gloE1Ugw8xjMps3YGJ7QuCToCDW44gyxgfGnuUODF9J7Bvn8uhd
yhNMdn6u1bkqgRXaefh65cceR3d53Qv5CUL01l+We9mwDf3fs6KrYVfoRkYxMhQc
l58Q9OIaJFjDYHGUpCDyfczgrZn9S3osWMdCCMiEkT906y5KP7diE+t/QRAh2CaV
bWOgKO3/zQ1PHYPnWJwOzqBwNiU8giPPmwlLtgmqEpOZdZcZHg4BGEksBT07kGUv
nCJxSc+K1u3bhG+KH4WP3mSl5nmD/qVfi6EH8+jeoNAgxnRy+diSjvoLVMGL7Ovs
M/26EF7h3uiRB/tDfJwSKriK+enrynFlh+sHkNiKW5E3PNQhIISOShFbMDBLguXY
UV1gX6zVCL1IB7ziSM5U5VPpxOCmxzyS6Cr9bVEaZluWdZ/r2Lk3xjTYRZJ7NHZc
ByfQYzpLW8dGXSpcObglErvtqMvQrtDA5h/uuaR4UaR2KSEERkLeuJmbf7SULMrm
3a5qsB5PwVp1BBNR3TcHTiZNyYAAb2kmKcfkLZJo8s/34Zf5NOnpzjP18SvBvbNW
hiHH8IiRdfg4mjKl4NjjsjuQ0HBt4xfbBxFnqAETQDv8r+TiU2mlBQT3VuPLLpTp
uOES78EhlFxJANNTeJ727cBeiLzpNUKxyDjdzw1PwplJ/RM7es7e73K6Ktn/kT2M
YPR9tqXgRxFt4bI5C37iu576jcI9etZI6AvHzYRl7XQUjgf1GN1QcSgt3kOD8V+N
9O7o/Y1/DrHkDVXJpWN1TankuBAi5aq/yoIrzclrst7uPJADg0ARZS1trZ0gc9ZT
yfgqR17wMr8Gv+yi4gInvWv7ouCtnfEfjBMnD5veZYt5ycO1ldPKrIcQ0CbV64jP
iyCnYXDO8wSgr/rwPVrSG/EhSUii3eZtu6BtNSp0hS+InKVtPyu0O29xb3cIrYJU
lAbRVbB4I3X6n9Rmf+qa3F8E9Qrnpp76IgvcSI9m4fUQ/+erLT80eu00G6NMl7n6
fc1RSMEdeuaPCyUFJo52HYDPNcYh6GuyIql8asg9vn+85lcadoyRKxrO0E9oZq0p
eQUGpn19XTMgnp2USi2gSY2iHn4KQVBt52adljtrvlsghEwAmTtAKB097BWxRSWI
DjuY+G4rbfaqmkAxZ9+vmqDdq7gO4/rnKLjbbI6JIbevj+sigz8Rh18Z90jWYX59
hr+0xKjxWOO06D0Kdx3hHE2cSO9ZrOPMU2F4GgbctdRA31h7G9T6MzwotOCHINBq
pw9IpN7MbaiNUW6jUDFktDM2aJGi4GhFaRF8cCJjCH+y2Pb15SWmbC8oKSa0uKyM
cZNl+9Xh8j9IUEZY6VzEr05dbv209C2QmO3oTWtcJFgVWeaQo5yMKE64FFMyvs/e
utzPXeyByogeggxvHCHcCszxC5RAlUDdTIZdEiCeg3DHIZJR9eWjdsfViSRe5v9J
9mu6ihzBkYdFT5rmJrVngr+ud7OclHi18KpFog+sauGvOFKjV6N0jD1jCLW/Z2hK
hJKnK/rKY1ESrNwi7SOVR04+x0PFBwAosfS3vpxxFctGIeUqFCVSN+sTEWVWB87x
Ufgn24kIrfaxEq7GPcGC3OFdBfnRtPvXpx1+Y2F+haSWemyZwS/eqc4nArTgfMlG
nyPjvbTFUphJFB8SAVXwaGSG4sdetqH+Zr/3+nLwoiJcJXXwuQuP/Fi83AxDQoLo
icjFkmOvGvstF81lgmAqrngKtXs385AL4MxfxJNQH39uK65covVG+k2Y1edm5CJ+
oasU6QOUO+JtPaKvPJvRHaagQ6urp20KFx77rJPTFEIabPm5ii4a8OXJBsPbVqgL
qQmVU6JwW9XBiW6el4HWJKhcKab+J0piY3/XyD9QAPZUUO0SD04akI1LiS+0TMsq
nXtrJ3RLwr5gGeqkOqFGi8+Bm/b89Uo5UI90EV51cJ9LQ+FVHIqp55O/V49KxaOC
UD2Ox2kA8KgXQznLKxPBnyaRXiji9xRSS7gOCiFESKf2QD5W9taBbO9nKMsQpgND
mO4y2hR69XVuIeryDIJCQOciJdBrW3+WuhfSVKjciuNWEDrTJhYUIPgbbxZo+sqX
CDhp0Cl7OAi+cOatWodPpj+Al16c+vFTCXHg7GaBf0dEDukW8dPpC8f7qxUY78MJ
QF5+qvE5FTg9X1NLd/qR9nOZg59ETuDq0G1gTIGMJMTvhiJGjLkYBTXHKw9IOCVU
apwMPchlu6F3cNxE6798XJVjvf4+FSrednBloWiaSBltchPYlXIeeOmVoUA1TLi5
b1ylzYIfwAQL3PC/TG8k5s9ZIj0pwGRMORYoe2IQx44bTv4lwXmAnw+o2RKHwxO6
S5GmCUE4mt/2ygJafW0rwLQNBzCp7pO80kHacKyU3IlKnhntwqqforFy+q0JN02v
4hAoeZqMplsmLwwwfSMnFsMzqPLb4W1cWRUyJ1Uxr4DOy5vc4jpiGn28MomjdcD+
2jMJCYLi5X0wQSlwQx5X8Qas2aLGQKiA88GYKo6rAgVpiGODFj6l5Ri0Tgptszkb
5e14+ekxtoXcyv/giesJrYFVkhrRlPEk2dI1QRXG+8wgeHhmh7KcV8iIru7PgQg1
N/CGHhbOOzIiMUzyrHOgGI899SZr9Yx0cc9KE+3+CYS8NGREuVnBLHWskr1ZltgB
R2DDxGGvQNQlEjvG02fsQuretCdjSjDMYFY3SSF5owqZsjqqb5rhlbIPzDrAAJce
LDbe2syCXGd8Woi9m+85gN8YjMBaDpoWuPUCQFFS/Qa9aNadMebtC4fw7naOZDVT
m21Z+nwKgSsKWMjcNLpEMA29W6+UTdukMtCZW0YTWodxbzPmxjkbwRyHCXk1c4HK
cxBilvQcHzkJHeh+yRO3Ag2em79sIwh6Fu5UIFgTcZ6Md8dkFfGomOprUNCBF5Hr
DUo/w91LcdWJUbDfUHqE9Sni8Muhq7cwxqW9nNuigXuK8pGsYE3HB87CehP725Jl
PiJEKU7Jl3o8vVCiotkuBfaeObKhpZNsJH0lRCVP9gycvgQqD/yMKCCeLXwJreUO
NM8cedVyVPhV+b04bGgDx2+xzFM4Uj+Xl6ogrdiR4jh88gOdcfgdInvJtK64t7me
V5x09PqtvY/8S8m+pZhZ5Se3Jm88M9SzpYZ05H5oGcHl6rSJD87SkGucLDODt4ry
a4T28GuN2ORTz7ui/lKULRLx4FCTuyLVw0Da4YbgB0eBCGe4LEXEcn/D8mX0I6QF
do4nU00Nj3l3pR7uXXWApmGKCRf5j70CH/MTktUYLlCOEd5+dBDt9cO+M2pjs7Ja
f5/WACuqgFuMLAPA8WKZJwdPG336Wvxh+MAb4SEvD/ZTMtm6/Aa7DKs0CBS3dSYd
44NRfR/v9ipDSJS8wQjE+gJ165usU5AepM/U7+GkxXnJe1gTiP7xAATijmRrQ29r
9g6Nzc3jM8l/+7xmqz6eOLD+M6RGhiVdYlhCrqdDlb/z3tgMbUk5iK0949hfdmoo
JINScoY0IrRZx+J70IRVnQsY/jgDoqZpXpxtteL1KcPh3fh+GqwGP2KjabHz5pBJ
j0B74UyjqjzT/cepf1VPL4Bld6sm9zpR/uTVqfHriodJqaNlTUFsSzKrxzC9UfIA
t/CKqVpRAnP1MK8QiLCQYCyWSmCc3hRUNriKsAVDlE++o+hp8rDmnNa3AdHOK1ks
0YuYmNm56ZMgFDsHq2PxyAVjWCqatGA62sXxhgqkwzESBfBWv81kAJ6rJLfGfgXZ
PG1LhSw1VeW6p9wAsd4pIbtn/xyFvTQBIp3gy7x7GdwfUliLIhrqImzNuBmV/631
M6xisVnxaicZm6RHgvN52Q72TTHlWxqTQR7MOeCbFfOzpr3GHAOY87UW5+wY1fNR
JCt1Ch+VuxJ1BDpu7qi8JB9eI4ei+vMNeajaF/y0fIf9ts3IWX0p4JxMn4xGZkRA
LFLz1tbtyPUWhP2HkeDtYI8Bob2yG4hyJO4VG7ba0jMLFXTKfz7TNdqOwILIoULx
ueztsIqclrFKexfS+9kTx6zgnAxmIv7Rld1LASzt+klYYO4icsvH4+g8edCiPVSW
4dOrvnGdxDAmGAlywOnRaKcTpMxhkU+aF7b/jDWB6htRSpBm2IV5IavikTkNNjOa
Q8l77XoAzDTu07AQgv2VdUC2IRyXHnZ2P8xkU37+BZpj8dDLufg5O//0OWzbagdI
NndgCWutPhFbnYTAxGbxEkG0gZadlpWEH1grsXssms9HBuLwaZR+wG+rz+Fo4Xe8
AQ8ME7XcnVskIN54jVhQdt5wmBJ2onPXPV9o8AyeJnlsbrCyU8oTp+q2ltkeEh5v
/8ixx0dG7uz18GV4kBAS+w6rlDeC1DkFaj8rlnHp3SubFrAL29ZRHD4KOy9/Ybkb
k8EBl22qp1l0WQtjemexPYAc2PpjIWXpNMQdWcG0vORE5hAAVnFFVC4Y/F7uv2wK
0GNMy+FO5yJ1qC2IaAYgHud0xu0i6mBjHvsUlmTyMiJ727t1UdmkZWZdJfnHAYYd
RgjXCQ/vG4/qQyQnBajJjxTx9CsfvH5k00IDFDfwBWyKaOoFrBx3+c6lbOACA+cy
eIFKoS8EbvsgapUqJdidsbD4vV3BJuIWOKXr/ni0AZlMv/dPKo3uYDT9qaxp7zpP
h9CuNvz7RvGuebDEI755edjM9jrZD1fweqs0TpgcLytrSCpuk7udGpixNojcXZv6
JuVCtmbkSl0L1BKZ3pRkx9T27b+Ncwr3aydZ0oNqiktEZ5F/fSxM8hzDuqAHHDtX
ubdesh47jKauu7UYPZJNxGMmkzqq0bIADea30qgOLn51dTfdzOeKt3h4Xckj1dgx
GqL8hqAYCDGyy+XRl9MN/JEWzwvLAFuJ+FHeDGB3K1CwU2q924+NXOUBOODXi/R9
VkV5lvqPIeAc/Ids/BonlgRc3zVgTQ5bXBzgQVSU1tDRgtN+I7jMpHxL6eSYvCdC
kUxg6o0d3fI0NEMD0PzcMhcYOBjPn4QPLL9rILzzuUn8T7EUNgJt4svKWj4CqP9l
unmd8G0B6LytazE4t/bRKLImBNBKJqNrFkyTQNXPJSm81N/dqQdN5F/8qTRQr/jd
Xya2dYfP435RxHROonKwfwRU5PgukmwljaWsRz65OOgoZ4NqkyrnuYNmlfiHn6Yj
SjWYPec4aQyBNiJ4XpN/NIzWWJ46D3L/gc/m+Trl5sfuSDgRy4Bhxpvx7+36ElqG
QqzC2bXmbd4cXpPEWMEI7LxY8rZ+Li1x/X8lEEkJGWeiIAeTzSqfsLlUzYmfSyel
VAcs9Q2Krqj93g40apsmkWHaDCf/bzQukV8CgNR/T25tTM8keLzi+icFN/YWk2pB
hlOAMzHZdBH2pIawhyRd+Vy9QqLy34RoiARmQkw/fvCcPPfsanJdsWyScDoAJZGe
YgSt5eLdqrsTggwnAWaeUi+vsvqIae9YaisfoH5NLsEuOaIgvm7UB+S4lcyHXG3q
EG68h6KH4IesvCJnXcfxcDWI5vzaFdrd5QBL1KgGl0qcLd1Lb1WglDjXzaRZdIfF
vcHY8yUU8GtkATslhIsnbCHGc62eVmxOdMrtfLWvQvK30hkXnN5jNB2qEYNa2YRV
YH8sjhZEoc76dH72pV6eO9N6eWpqtuONY93/YcWcNeoLknEaR9EVRjo+A3MTWpsP
+HdMA/OYO97/k/4Ey7kFUzGzjapRCDQvJN7kOqaub0a2vmH9CtOvhCaazmID4LHG
D0C47KEzOCefZGcNAX0WAA8Lr5wbBSTmBk6eCfKzysX29+TFNkQoLnYfjyzaKqsC
a/z4DnHCvNrMNl1DC3xP0TZ/cfjVvOx+rMH7QXgtBxmgKDGXQwluxMDxOjaOmw4U
yjM9nmY3xXN6voZD8RbPS8tiTCrR5ybZiAyjafOaWvqfborg6tr03GtSYUye0Vvd
/IYjA3+clIm+WT6ieLgcXEkVf0WwNtbaJaS4gAwLLMIxppGU/QMRn4+6aFemMgHm
/EAkLpyzw/d2pICa4Kj5xGEOjjdxU6Wft75j0qy5EnNG4LKb7z42VSF7m2aJWTGc
Kai/I7raVaoTXDCxsq4CACIwlbI/gAQVs3KcB5D5+D/EruW/GRVjPQVlL0GRZ1kd
5CFycJflWpSKvo6/W5bI13duhOX8n+Q5jQ03ku7JGf1wkBZQhYsreteJMDhkQrXg
PEccUP/5y9vuNPa2iFJJz9BJU7O9b8/5oXLGkijTNDvF3RjnmcKhAxBikMPrl/p+
kPDFhIMGKlIMSvchdr+qS8vhO8V4HDR4iEQhkyyBd92EaPOKhfUTQ4pFm9W2Z70j
jHx8KPzurKHjhS7QUkZbSftwwV+0dlYlGE5euGtMlWA3O6rRbvw/M3Zy8ZdkG7g+
0IXXZdjFbxVY/u+k26QQFqi5Ei3YINCViqYN4H8Mw9wEC7dEdpHOknIlC0OvTlqv
UY5UFVLFjcrjOcQZllP7ngN43jSY6KAbjTzyonWSg/fjN04YvhPhbd39pWDs0v7O
XoGWRa0OTN+RMAFbuQjG2XIE88awn0qlgE06/DpFHsDVFfbzm5t2TzkDuZ/3edEJ
+lhWvsVHH9u7wAr19PXfuR+WuqOI+MfXJ8BuNQ4HWm9Q7SpA6FYVYOQSlWXHfPG2
hEMwogJde15zvVeca44o2SIVqDVn4SN/20+UtkXrfYLygc1k0v4FNET9hXWmuKCK
1I9R3AN/KkSFB+xbF9cnbP0cbieINOS7718+MyKMPf4MvLRkr9c9HMTWFvgPep+d
JUDBSxLmgIo+aKiv8D+erNCSy5JVHGqscHpL2Oo/OO/3pBpzvHcz6AUlpSJ1bmLZ
+QP7ZRv+K0K7l6BQSHOsmeSRaAaXTJ0P05RVljHirZTxqith/sUgkPqo+BMgo1FT
8WuwImoAIdb+qESD0cFEgwntrLQ09MZTKiT6rNrNfLqrT9by7qedvo/BWXAEPtr6
`pragma protect end_protected
