// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GNywWL8CMkwcsoZ+O+VQh6hdPEqlNxxnUj2s2X6/LDyphNHZh/PNfhdFi/Y4E89F
xJqBcv44zRkdseE+axvHIdW2bDVxc5oPoHHzx9RfLC/QKQProjyLmbbNiMFU1cpV
uvlUo3onFdReJUoijB3y2lj+wDZX7WhLb/a5vtgp3o4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14352)
XE4+YR9MC8z1y5Wc3Lfk63+XYC4kJEoCUc3Q3q4aU5rDcivoH/6GS9zgqZuxiNgM
62MZSlwFsgakNIqT8r87nlfSyGxwoWntfh6QSjRJKNo+Tv6zJd9n7tmoaQO9gafp
IFvFwnEqMbIwzvknFUYrVuGIVeikPChIPP6AJhCTycq4M627q5NHxBAj5S+E6KqM
j+K7Qy1Wsuz9zBkhcyEePOh1P/u7NPvl8MFHAqlnEi0ogFRwXMz58bDUlmIXE+ZQ
7NtB1ZaGDVVsqecwhEGa1lRc0ISVXFIOnTnSGtd4UYd3YRAIUwwVmM9aoX35P7OU
0I5o6R9zv3dQdHC8o7ojrrVK1CDotjN7WhX8Q7CrVzJ+J4Xa5S52dYBIanj8jL9h
1pDBiFTfCpCc18qLj8tdDriivtOAi07snC8ZGg+365phg2OTrfy9m7k/39KC5b3k
Cg5c++oVAlLx40mLT2j0CRnVvTcTVJkCK16g2En4+yHrEpw7Pphwrgof6D1kA3l3
CU+dFRjfb05aZuao3JelG6XOOhoyjp9hVW0GuNQoxd3rT4GcTB3dyTo7Cn22OrwJ
B2Nh3x0YdhNJt3lrOWnaV9ZwV7CTa0He/hwaNmWagJ4J5Xt2UA7/2MSDaoHbSael
bJ8HwLJWbiCelqv2EDJY2b1QeyU31xbrfgU4TS9Mb38eaW2cXWtC1ZSBpvd932bL
h6aKvY6nZzYaJfsxA7DVzyjCbRNboMLw5UChutg1NBMuQSTpGK0GYUkr9K34ox5A
djVnQ9T+i0Er+z+xRUtRGWqTOB7T5WX/FqMWlPP0HNR6dNUuExo58HHTd3H2kn/d
Cq6EkkasCHg9gKfaZ61bJOzJy8KObXyt+732P3j5/HEHsK6M8UgXgATTEyT0jNlB
eppQyRJqTyIWIqA3vCFzmQv/Wi/ygxgvT276+jnepKSaRVAv4ZodHAjz261Jn+A0
O+K3kiyvsmNwbUAHky8qFISf6Q73X6Gf925X3Hycvd1RRgYCUQe7Qb3Mb9mdwOFB
Od94JuYdwPHmD5I/sECLMNSg/6OnWVvuZImMSdzKgaWmGZXCnZb84srSvri22xWi
aF1AOPyH8ETzEq2V0ryyY07vmBTIXUWTspCBSVozESgatpfla/DVnrnLd4QMJHJ5
Yi6LU0Fx8F9MtMt6UNFYy0iC4D07PjoG1zfxl2wx9J1YsSeiL9b4+sDtEiG3cqkX
DxJgFYXlYITDbJeXhiAEfnwj2PILIEk8YGIay8jCsO35W+ePp4bzERQEcV2DURtq
2r6sBvCP6Gnpl5oLyhKPWkx9TeKon3siqvt/GN8XhGB8ujxAI4pFDsVXPf+zm635
hOlHIwMSWnEWpQ5FcMpn8QTDsHiIqK6myj37Y9AejMAcCMveHClTgKtj2XT474l9
dEndiYaNtiRNYohFJkes8vnHdAzSEZciWxn/R3TiKQEMV/f8rvw775ZCW+H2kxTN
dozvCE7OtSDYegi/GzuctellSTYm7FRQJC4gst8M6K8No6tyDf6iZFnYrISOfvl8
Vipoh362SSgxT5iL36Lu8yQX89AXyZtbgs+qq8K7t3xeVwj+FoCONDPjDkwnvrMb
Cn8DejwuGfJUQifSOjW8vJ6/6gMqA827ZVs/tussYeQ6MpNaOMZrN6qr32y+Lag/
AkCUhEkSrB3pnTWKEhKYbGOAqs+U2ZY/R3eKXlqe0xcL67v8unDQPJeuPTlstlrc
OBnfP0mff5m1ZC3AKP6LKSp8Ply/1enZ9+o6Le0A5eUTxOrrAH88g5DM/M/2v929
4VgDzCdIbZeVP2WUdyEqRbi4OdTE8LyWSXjVVDbVQ4CvqtDqIls+kLuJFN8D0g8y
X01dLsOJ4kz/QGCYFhi3w77AfRqks4233A499jdZYC/S4UJlenqOq8Wfqw9aeqew
QHXZrSPwLjkQMNpi1A0ZQg998yEDTjH6iloBhcL1F0OgG8TtyiNlgwHRs5QS9xre
34SJh3VMeciuWRlT5S0Pda7H0OWXpjzz06RS7GR6njEcrRWcpLqyhQ+MRQ0nu393
iVLkxVPcelBBRZGLX8Rk//vOVvvw11kp8/+CfSR+nKtiSAWNN6mNzTJofK+RJXmt
9P6HJ4EWZdRUPJ40eND0MsgYTmq5/1FEtr3F6MNcUxfRxMd4S7U3LVsXVdDAh78E
LUBcGLeozOQ2i9OQ/A9maVcN70tmm8lmWT6bLsjZ35Y48WCeXuvWqevnrKoxpdPu
NibCAVWWEJGSLBr/uIk0DTFEERDK2fLve2XrWNcNybekT26DugM2l+nvXO+TddIk
l/BPGO+wUOJrjmgBG4cISLnrLX/j/hipMYlblqwBZXtQT0z+ygFo70q/+7+Mhus4
szxfczx4C8DCYI6amZL3U8UXSn7iezwa/MfToCOVWRnPfhmqksX5TRB1le2bAJpX
jkf68XWEHIAV5hKcrkYP7MzYnz4eGKhkW/eFo9oNG2SyJsJR5dr8XmuavEuS2hVY
nPkqEAT/bB11oncU8TStNLMp5S2RaTunyvvOD5/ozQpV3MSoCjImvReWwavfZUVB
fD/+Fr6YSebmHebrdbV1uc8MhL37xJW+qVqA7a1SAuZKXlwgfUpq5TjRm74BlXAx
DYL2Xc44yL2rZOJPATuue7LFz6MEtrAoa7uMzjw+N3yIBMu4lnyYrCWqtBDlt4JG
0igoGhMetaHAJzK0T66xKU+zdudb9gBrBsfm9L1qlJpng8MlZ82nsjs0mWurdXNh
BSqQxqBTXdm6+/SjX1zKv12aZNK+QorgxC/XqSxxi4OmHkf30IaTW1oO8tKS7zCk
UzmFEiPTWApUomJUVrXRI+coAqgF7f9sNY83jXbYhiQceLUrxo4M9zNFoLEffdl8
nrBBwvHlZQs6YUXh33l7P+D+oBOaHXyRgi0JJd1Nqg1jGfRJ+FxQ1HrLrRWMcoEb
qeaVeuBMeMi6jakYpJDb7GsxCSoyeLskC2GSrUkKVpF2iZwvWdKRBXNH6WAThoVf
GDqDZD1VC1VzSsr12t3320vDx2HLtuQfp+pzP4qq51YrlBMaQUuCgXuFLs0ecaaq
ZY0SljjjN7CGoQRIwhznLHdcLKNMk4CFhvtJl/TiJc9Ou/+xajaK1TamL6FMcnXc
LFnRpVh3nGcSonZoo+U9ndQDwa5a3c5akX95LIJ9S5OPoC1jetL6CCnrqxWejglT
497+Vud8RF/MVlpiJNpwSM9t7LEJxxfExQu8jqNsgWSEAFWRHp+nu6SjkvQZFHH6
30DxAvWC6GXMAh2moW9MmWU/nLNfdDdaDPtMdQSS1LEHNvovB5yWsS6ttC5pCh+j
08w1Am6MoHbsJm6B6mpwAafoqFt+gYkL2KTTcqx6ztw7rozrSug3IyjbKiUW6hDc
40Y3atT7HVZ7Gop48C6EZURz5PYs15ECZ4nX/LcNgz9JJjx3WhTB0OyVRfRA6iAq
bmM6tnGWFj6UgMGAqI8YILa+qelFihTL4Dj0hrWinHADmM05CKqdLw8uqDvG6ePv
wtyo3xXLAGLhKQ3vKrh5fYkMdTvFiqtrKkpRGWVsMY6qrGEmdEko+dcB5qx9k6it
Bq+IYNasIGvyTJxc0BKPEWbhn51UnYQDPcQnmd0NBPKEIeh896LxffeiKZUbF5ne
z+eSeWcyNELCiQ2TJLhAdieI8uczYpBqTRDkn7VS1Jb4M/vxgNfEYi+R3e9CprNN
HWD9FhEL4p+708gtgkrD4pXxEowSv34EtmnAXx1OE3azzm3Mis4NcqfaxNI3oiBM
5R193mrOEePrxgLGQICGK3ZRtnJijAvq33V3S3O4ZXBkKONZKD3bt1H/ZWL/rDWo
zmEGqn2hRyOoM4PLu5vrNHHHFqOLLKa8vTG7zgOutlX1MrFNTSrUGmP5jMntCnON
+5BZBnS+c4ovEdpLWWExi/JkEBx3cbTd6aL2Y6nVE1aTPot5XSb8zp4zQzQreuFU
YLLZ203KKj+nAZXo+xCsiSfkeQFitCom0JZEHw3A9Ab8IloBfEo7IKMP0gI/QTjp
WdtNaoDyEdsvTN6yUzrPLCqTnNz1RLNVf8DhBStrNae8K/URQUGDhaZakGt0saDk
wqqNrEB9Ffk+cAnjEzKivwxUeYNJbic852KeIoI3E5fDRwLtz+lqs/cSvo/Or39u
aGtjOyYZX8I6wG+d1ZO/millQpJor1C6rPxYE6Q4EYr6q1D8CoUZlzuN8qWEWtl/
VURwFV9exs7cyOpj3e/ceXLM7ovVtufp7IziBXTJP3AgCCOFpowJegCs3LJGdGP5
UhsF1EhgVWaF2fGuDeUOtd7xhGCnHOmvJ7z3fZeYrLXj1dLt/X/ecW/IPbeO/kza
LHrLRE9wvjSjzo5JJ36um0VfPM6d6H+PZ9y6xMdr0w1y74VcDhJwbKVrCOmEyshV
C70CGHVdvC4bgwVbO27GY1Y2XHA3BQpTK013il6U+V4ezsUhZ1OOhp6Fsf9aD/LH
MIcd+W+0H/K0X7StZGWIo9hd/fMrlt7sNHsbRElJOORiE/6Tg8lGUv4z/rdRmBNn
BjO0+Jt3r4AP5z9YTOa7Og/WHMb1CIYZFTPjMkmP5Wp3k0jDFfhKfYCWVkdPelzZ
OSWJGh2xQUXpTW/NTsGmg9uZvXjnypsTNWwQrRai5X+8vmu6hb7ErGopz/NQ0bLS
nAGcQLw10yK/APxafO+iVWzVxMUvIVXiIQ19e+IROWREmCaoLJeoimapKUInWbnW
I8e6u7Bw+iSjcmOQGweDO5aUUwUklRwz8EwOjwaQVR/OrP3Gor6dxV1XU7eF64VS
hHn8hIzRyLlaCnIQTGQ4TtuikjSbiMN9Zuk5gK3UBsCH4dKM2ihdyvVNTeDedT/K
TLzSs1vOk+5ezlIK/wnUzH1i3iz30+0rXX+gPh1Ti20V0eqtfTb7NuwSDJmh+eEI
yuGiZAhkyclL5JMDPZXi4SZCF1wkyhxMd0ECc/7QvsYGt9yVnSx3Hymtq7YEidjT
GQV5JcbtdtysR/xzbE0LwjmtuemojY7Od30h2meLgUvmvQQ9sjmZhes/zNUQnWOR
/2bI2lSn1H5XGRYmUZveLsAEjubOck65nHOjK/cwtKBm2ZnJDu6DM+CFtls8iUQN
u4XwO8aq1y7r8UgZhNHvfVv35AMFz0raBzzc1wFKkjY0hw/285RrpqbjO0JanNRv
0VDsbVlEDyNTCmMwdhv/TuSimMhCCznMvJQyj9i96hwsF0QtcQKPREYQ4c8doOy4
/0FMNN8N8I5KcQ96sUzXQBeL9q2QwlWKonB0cfB+pUQkDAr6lRhU8/ovFs4Uv+5v
+tQXkIYuOfiGYLxtPlV2JuFHWa//XrS5pIey9rRwbe8Pl6+zaTEs/TVomve40sym
We0UzHZixsZZWkTwRYPMQGGJGMKNicYD9zvpGiF6GI4hF8FVJv7mlBvxQ9SY4Shi
ShY/X/ebn//YNmIys7TPbWLwFTVtYZo3z0C0/KDytI/W1j+HusRrwyzcnysxfg5B
kN0tDok8d3IF2rkMcHGLY2Weh8pzYZZwd/pFOLiFYVrW47Yq/+DktoUWInAQOwZM
LjdoWEmL/7LMWnKkCqdHFqWcM8lJUSTQR4N70m1dvkbbNK/cxXLbD5W2gLVWUx8y
iWcVFJbO8XHZdZ87gn+VKaGuM/UKZrz6DG8Bh2Y5rtqNseoUBq/E64S/LAQARInP
YeO7NiD7odPbzXQ1nCvGEG1MxBsxLsuxfie4HoN1/Qb2+eG6qjJc/V7IoScGD4zC
L8sBj9movhKSy/PqcyMrheLiHBCibFOVHVphKXLsXVHwhXE05tKNvPQsAq8z7FQQ
EveuZVH/7qIF6ewTUBw6lH+k2IA2WhFS3jXQcK2p4xRH1AWSTxamKgsJqs5EqlHb
5lmhXwJmh9jWtUtet7Et0tvRf45V2KqqNoHx7zqpyAflcvnWTrlImIvsZ9kbmCFP
H5yhKBIJUfZWKsNadob8DYbe69eyumnT5ouRbyI4QXpfTFhqoOzfPu0oJ4HUBZ42
st4F0cFo4WV8XA2iLaPqa/PCdKyAsJzLc6dshDqFMxm7Z04VWzuFaXWoqfDlaibF
BNts5GolKeHl0bGqx+Ly6iyBcge2k7yeHPFAk6fhOAZ5/m7YcTJwvxKDQAp4NemZ
58JKOx+VbstYSLzFprkgUT1fLKscCJS8092UtPoGKz9T/ZJBZNZQ3t4DK1uD1tbO
vUoLnDXSxVV3393U3/gMX36kpo9HVOBkPmL9Gy9waECyNKaSjRgIHXS7rPBQC9UC
4pq+xXeOiacWAXRraXZjTOjNkrtP8Is6/QC41frg8ZqU4AzoY1Au9POjfNzHvfTl
ZrOJ8hHTDztzfTnQPjytH5Prh7dzTdPMsNw1G8UqowGYI3W+hLUbPSek5Zmkwed+
IpJnGN52U7/aaPYGWk2EBPPtKmkJNwWO+3FPRERE1k4zpisURjRE64d2wPwb/YAH
gx0P4qHjzs0tPvPUuZ5uij8jXcqiCcDVmN/pY9PvnGaVh1dk2bH8b1voBNLXoCPw
EQEbHOm8ufbEpBKujjcqvxOxoqrv/NVpBqxiqyDvQ6AxT2Q5H4MaEeCLk5pcg3Hq
jACcwleCsnFMN+4kLUIwW55o+qEzO2+oqg6HQYFqnhVUXIz5XSQBogzaoKQ7/pgo
PDA7RuKK2XMusIJRbacllAYCCu0rhYH1JtnFvX1smEUY7LBUuKqh6bR38bIX1WGK
mkR2z61aUuUBqnbc0HyAVBXAqlFPYwvBwpyaGNxjupMtMkG+IrsJtA4GWPMur1sb
ROG+f29cc+7SIEDviujCDfwt6kxOo0az6Gkl8EJld+KeDiOaOLITlQ3CV/YQuiTJ
aBnO+10CfQHEhUrcXtNK0eOVRhf1CY6VYEPR6OGpblVrKigXCyB2JfMAxiwgiJTX
fHHRWLNF9FSc2KjEOwLB0KliCugGAx+8Jz+eZ1OX1hTb8bIQzSPEhLIcsUvFfYBe
gIz+6FP9onNIpsIrrNDK0KQ9M7poauLSSqb02wovNh0NZfZQ7wfc0IEsdsRZKqiG
n9AMvnW9eLnKw/yy1heu+zdFeF6ioVol/Q1yf2uzJBi0sCwchuqy16U69x+aq9Ut
oAgKQj2kiWb+vj+390uHQz3LbtP++HLFZweppFWBD04FMQMuwOzUUuuS8w9WwYgX
6c42d+1UGe/tNQSO69fXox+DBZATByHfAUDpbhg6/LnCALPvC/uJr50Y6MnE/E5u
v9/sCwP7SULJyHYBWROtEIDETI+diZScf/1sqNV3ev8RZQ7kTKk58a+BUdMY2dD+
3AZEZ4C3gGdChUJrfBB7Q8FLlX6NoMVXs4hWUcN0wKr0lx0WE0l0SMmEQvxSTuuG
ZZShWUytSRDq+gpcEGR7w4sMenVVAjAE+yvABZFhL/o5D5DEG2x+tadsAY79uDNi
yr2zCqMcDESBV3M//p45CIw75xf8w1tvaoA1U56GPprGerXo9waTx/4WqNfQDxdc
s8/xt3nc4GLJnihAMDLBJ8KAh9O6dT73d3ACQ0GMh3yR+3vwG+sQGB5KGkPg6Gyv
9MXzhuzsMOeM90w+focNZYTfTppZWcFCwsM+C+Wy3POcV/pqzcW2/jwyI7+XGrmg
afyTofTVADguxo+PO3vrn4kBIAX5DT+5VluBCwT8qcGIa7JBcJQO0Gpv/4Ca9IRd
AOq97RuomsCI120Nbh9WF435FjlM+5mfhrrt/in8XJkQYk8Miz71Yi5ADRiOAJ6F
/cDF3EzjpDN5PXkSZwh6HF6LS5wK6ueCNGpLi51qD6qZ+ClRlYwGgGrRRtBTG3lX
dHX49sDTh6AYYBD6y95n94C+BGmNSFxzg/S1a838Yk8huxQ8/FAueXCJE0Tqz4f9
qmiutWH25UmTu4ubtJQEsswkP+pRVU8kOy4PBcfU4yBgA3fkrUFD1mxF89v+QYqr
8XnOeFNNQpCMmGNM6n8tuSAtp3Fx49wfaxcRI/KFU1B24zm3vHUelCpV8OUOTcNt
SVSUJh8GUgT8JJg3hea8AcY7Z7YZOCyaOQGBRTb796vNuvR18AHynWrFStNpxh7C
kfL9fCtSwymsUPqVSYOcrqCy1If2OVedAPoysPdzXDVObXEX/bG2/Kp+NVG+90ZL
QkhTGyuFOvWsDbH4NdAEPJ1fD4X2NWS/9h/KY8D1vM/YGvi/yor4ghU/L79pG1OI
BsWqUI10Y2xQyMRUbxbawRc/OFe2shGxKqlEEsw35FSh7Ee36UtQO3zJ7/aGwEAe
+ZY1u48yWFCBkPY5XjBXIqLOKcFx3tpYc1LfkHsx6aFbQpsx0jrnbEwp+9SkEzZD
olJDQJS3vEQeC2aottI8sE2gddYdYV1Cu+JiWUdUbCdq7wS/5zPaz8n11HNpd4RZ
8sYwSs0kRwfG6kLOw5tne8x4L62ANZ5VL1ZJdmp7E392mwYNP/+D9/XABpJwIC9k
31kq1mXtKVMUwbEkgHfAWa+NGBXrNrM9YxuMdnBjFDmCUXZl/fjfyW86aIPa7ftS
G61pytkL//o+gwZ6MyYxsOJe1R/5jxmHcf3hSwLJT3mbjtkR3PSykVl90NyQdpl5
K3dToKZ5eTlrlV9f+m7oogORKATzptN/PIId9rSFa9dnQfjZOeZwfhmn6M/mqvkr
yEMGde3qhh4f69yYslSccPP3kXJuCFWQLqo31vZeTPnQ7QhigOEGL4Hej9i2npuI
arjCt4htSzjXJ5DzNaSRHUwESV4LoPyGbvDYLrwN2FMyRzqhggBXiDywZz/lQiJH
oIaadUDkB8hHG1E5d6cNQrOWw/ccinwYfouT0FmYXhW5LQzPbrkv/HiQHilg/GzY
4AMrN4Jbz86RFvOUzrTs/yCGTD1qCfP35FmJ/LLXiF3RugdAeRbb8LU0TEewR6ju
C4cflmG1Kyq+tQxVSZhLUeefI0RUn5cvrTE5aUJ+PyeV3jcqclcSZgXi7UUZA3YU
qDhV0HnisdwBbGQ/EfUkOezLAgFE8vVurT2Jy+EXFsWG37OPIAg0NYgCZist1koc
mFuK1j7iUxZSQEub598kx7LuagIo66TYuM+t6ujSt77oBUe1OZV3EY5MxGSX/+FL
bB3LgmqjbObLTI896WV8x9FdU4WpN5HbMvnV7ltEp/8IWU6qdhlndroIdTqFW9hV
x/SRMFDAiJ94OMQBrIqQcJRVqIa3kXPK3NszNEjvJtbiCSt6J/gfwi5CO4Im0jBf
23n2YB7G4RXVxznytbYUe2XPjsZUumvnZT3yceGimcB3rSyPzm2UmWP7Sr4djAXc
Gmdt3tsy0UcdjUeX6Hf6J4hjHm81wHHmofnbiIU0mzs7iudPaZz4QGlgFsBJSlhF
zmNkFGRaOJ4jLmLD/6mKzCtxA6zHSHnCN8Z5m3mPIARRqtsuFWib+YDQZX7JXbne
6nPE1BAXISccAQJM4Dw2Zpl3Ma52hZiV02dL0lH8wUOEM+yNe4NDhKGlHSA7YWUB
v1runoSAzg0Tyxxy9HvHKTtarm5hjDjpC9CP37IDwr9ER9OaZl9c+gztQ8PXeL8k
VcJ787VlwyB43THbv83312aFHkgbdALWQKcrKjaNokrIZ+VaeOwHZMsB14LcODI+
Qf38ckUdQc2C3xZkUfyGEOM17qLUVCIQ5uTkiY8NvlclEslmPrBD3hrFT8j81brk
rjIMzGGxmXHWX7lconNT0JK/1EFzdxjbJDfPqTJQD2yQ5dd+fgs0mtg1Sx7jiMJY
uEk/OoHfkdo4A2HJHMdmqEQa+PMLRFxp2/6KMebY/+FvQCOrEMR0JP2ylcOVcxM8
WEGTdlyRXbxn/GtiE9uP8vwiszw0CBke7KJrndCVZx9ATrJITvF0TDRm+ERGFsTr
0yPU/sQ4orLetTAiao4WA9OQ+3AkzdqaoVSmVtmR/FXeUO39TVWzDHHgW3nmNBDO
R6/YBiIpKztnyOAeDXO6adQpbZP0S5kwAZb3Rrc7u92xG0xNmB8/8AgEErDkheQ7
LLN70q2Rmk6KDDtLHbgNclixbl/ShLlR1AgC3xI4+RWmus2gP0M1fsonYVVxTKen
MnJednPdGf1f+Rl9LfJdhzFFHHDevGbdZBqvAjZvmpcxBOEK/FTNqsKIIgxBThmQ
AwMWNA5yt8cWHpVKKXaWd69KjXnmgqHJ1FbG8JClVNeuEcKq4+BKAyPiLTlsRkjP
90+d86uSChBAqQscTLQYhkTyM/aLlP9XGF9RprInnrMChjK0zzDebbZ4XGxjpvLs
yPeSpAolzYxMrAsKFk15B76xHzCSvK9TktQXIMjsSwl8HNST3oGfqbrWnul39np8
2do74mUO/WQqld0+afRS4JpY58faOlxmHJtV+UPt1kmLccnPsGR1JJPO8LFHzpk9
Lv/r+z8tkmdNWwOoy5Yq8Go4stnEFn5Dpq7ToXoil1Z1D3IpQOINLGM+Lq2fdsJj
BHCKaBJ0KV5zCOnfThin81ZjlIwNycwlg2GSuVdBENo/NAUiKQHopzZQDA7SsbCd
c91PhtB+StUEcLN5w1iyQ8kZlE3aWX8x1QFVqnrTMj6+JRY3+rqq7XTMPnml3Rfk
LkToB1AJ9kv7i4J1/+A77wmVHIszlUIzRf6Wm5T3AJBqia6GRnWG+w8N9jp2mIBO
ntXKtJyCl89TrPgTtu7v4Ok+Du14BByqPU2G0WQlDL/GxwAbLjrK6doPbGtcuMaX
geHUBOF3x5dQNNxHqD5oTo0UuzW6UhDa4S8u8I0Pi6dPoF536gWb67OQ5QdAw0GA
o2oPZTf9O3eq56STPFAzT+PCtST4zVGKhq2Kbqk9Po7fxu4c99n/c/gwAleDyein
0ZIV0vAfCzsRcL+LxAcvFWyz3OJF5wfvW9nJHK/do/OChMlPeYPWs7xEXZc3Wq4W
Gmbp6vUxit6ox9JgAZ/tAw4lkYYWXa8xvOHhf5VCWo72WP7CDYxFsM/a8unmtPEp
tsRmDtq6io5DzeSO6iFvJcEuGB5Idzr4Z/UWLppTgCA0jy3PyoqbknYKMoaEpb2V
Wk4eQblhcnFfY/yGfZGnOPScN7hxyy8t6t2c+NsgxsfcbT4wcL9X8EtrJcH7EdEa
HW1LI+ha4kpassCMCLBjR0ACE1gBT/TMPvtounTYvha/pnkUP2jEHrZrU87gJtjA
djJwnX7NKBOMTtHEB/Je1YZ9xmufoA2Ltj2IlQZ7moN1FprpswL3L7aGivod0apn
uJ+hoYwzffp2yd/PFLKg2jj49SgEN5A0D1uSOVRrEbW2XpIR9sukHKHg13ngA/F/
4vH3KacZnGWz03dMytiEoddo7T2HyWBKx2/m4JW1cx9MLuwBqkNHjoXhcZTFmdnN
mfjEZErH1hdogQp2twYXmnILnfhQIt0omfgvrk8FqRAkmoitOBUOiOGnWHzUmb4+
sLrlSAX5w8LTxNvMovSP7XlyGxJAhidRE5KBsG6QJLLaL9v00amntk+SuLadL58A
TpUFITkZxr3tvvPltCfHEiTt8z+o58UVzcZrm0jKJcTZy65KHs3ozuiAVffVr7ZE
f9J6rs2hEaYS9Bxil6VqCvUFfloFXyDibMeB0J7e1PYOWhgIOlZIN6cusYvVx+9v
NevSeza5OSqMpelre1qSv3dcNSU/Vy0FOepCQr/Z9Uvo7vWQDuYr874yzlhVAckM
1/pYnQndps4eFTBioLcEWlo05wdh8CSowr+ZH32m5temAizQdzAr8VViJzwUm7XZ
nOwv2ydHdEwWx8pdJkrYYJC7L3KmTntBtKGR+A1QVlalPw7UwiGEYyx8VD+plHBh
/CX76WDN+Z9t5dCu+yGs8G7D8zHe0UyY369QBOORtVEHHwW51ktCuMwIuAakJENF
ns1r94p3uectHdPncXQZsAsc3Ul3cZqUFyp99ST5cQ0mjFZmLwBbT9FJuZUQxHCg
AEHGtZVOXesC9GnA+D3lbLwZDV9W4CQIl/HLQ4A+Go2vGcAk7MLKAD5MgS5f8Lhc
bxg6cOTuvzRpYqH8TEULTzRfrP+Uwg7PFK3URyRPrnbDxo3L088gRb2WpM7JKjz3
3BLg+EASRaFWFaqX6M33okESHWwpFxvMvI5TLCxA8Dvhx0KFtE5JV7UmdrNDxl+B
vSacMN1pb51a2FCX6kDYUoHHVZ/k3ahbMm1x3QL8R1LEgeoc/VLW1C9wsMP1dECa
a5BARigE8yXWwodYsmhqjwKMbjEmmodIir+nBuMFzd8UgsEKgYNMkRZBUqbwufm8
LbEvbgOIoEIeUbKNXDGwwU+vx5zKA78ZlW/H+1AclfnId6IfEIck6SDWZ+Hftvho
W6v0+g1yH/f0NPYwPnD3nO9N+1faL+Lemb2PChKXQkGfiAI1zz2bDtOQnqxFY1N7
F3orISw7+h/Af3TUo3uJYgvFfFB5TSL/tMGUsplW3fZAdCEBoGjNbM6l2HBKJzZy
nWjviEsZ/WN0i6j3TvkJiuYNECYdgiaBIczIBSIvsiQEFTfc89Ei79B0gpOBck5P
RBYHU3wHs3Ex/l1lhPLetQOYbOOLX5qoRBDP8j+Tbgd5DymUxQPxt2qTa/xcKsBd
8SNpaGZdPehvgfG2v/edsbRp8zaBp4lZV0CIfR79Y1l+jFEWV+C9eBBYHWAOljYW
9NcXbwgunMEx1xjjfP9vZesp+NH38rbHi7r5RDopraksg2M2pvtKbfp+r1ATXogC
Wpm63uOLDg3PnmHViutFpy5iYb/zxulSsB/XPcZX30UAywBMughTZ5hoHFwxNiFI
Qe9+seZyaCB4UOXC0wDv+l/VcotvUYuXWJvIqKKrhry3y1OPcQuN52QW2YsPb8ca
tXN2V8Q6T4TASbXTIup/QhPwsFnlOZzafohOQTO9gckhe58uJE3TnBK9E42by7Uu
XocroC07QFDgY6Y6OzTYq+Q6M7HWJbYqGWuP9z6tVsWsTZuD1/oxS2xF/vc5sX0l
Y49La3yX1gdHggfSuV/fHy8wpedMlqOdIc2TY3wQE8MVX4tV6A9JfloBXsN6CU5F
mpigj97vvvUKCmgnU3LUj+CPFdIxtbzutMI+1rc07VAfyZLkO1VZZN/3I0snSGKf
BFlO+7V4qLzqh7cW4hjVa7sj9WkRkv1jDsIAwBWfYazLMY6/u+GnVKHwgyE6ALRV
9TITBPrQqqFfdp+wh4/s2tRncxOemLUcB7yWDZt9zajkf+Ix+zeEdzS1cGk3A+0w
0M/p6fFJaPQFJYSfyu1NLLbzKMOOe9Rgelhoml89cequqpUa2NLB+CbJSA91ylfI
sEgSRsrDHNucGUQJV1IW0SWqIbaT1Ep7CIHdbB7Sjb1Tn0b5fjdiwXVRxfnuFz0J
+Ul0JlJ54UQCIqtS0Mr5KJk9ULTLrzpeoP+awfj9Ro/ZadGSVYc0qqHtV46FnPZB
QHKsKtOnZgbTR+2O7l9PTuFT/JeAHRPW+y6yoCyCQGr/4qv0POLmKoTNlH7Dj2VP
Cv8z7l8dYGB0leg0hJ4fAbcxK6deqTrSuTffedH+F0Be4qNqpRELWHJebJrQDTgB
g77rmet0+XzkPC9TRbQj4lmWi14fjWfmiPtjOsa9GeRRY6cy1UXT7z3YZhTBBt0B
91uPxQxvZVuCSpmL9YB5xN2ybe/HdZzuHey68RrnD2od84lcyKRVN2B/sKaWlTKK
hdxMAV3ZFaWtDJQM3hBE0DphF5Nn2IU3PCX7hfgA9cWJyQ+kXmTqT4UYv77M2g1c
xzkEFdCDK61pV5ZFTNAriAbmQj0subk1ASLccF3kvpeyHkfydrsNh65h7Eaw254B
bF6gpX3Yyv7G3Wbv80TvtT6RbD/IGRyseAz2CVUBDzUHUQ3SG4nBK1/zMR8jkjKI
zMtOerQrFfz+xnZIDWqyAf/rfrhYVqGhQb12RbddLJ8NYtXw3wSaqHoTw0w8NYQc
+Q37my6Ixu4GqT8sk66lx2BVWi7O4DfptFgUQu4nvfQsxEl3a4XPk6WJwVJLRVti
8Fr9lYLdR5iGvYx7uSkyRKYw7ll47AriZccEIiI4g2cIAj/tfmBVRRN32s9lXMHL
JHmFUPH+QN+oh8NtYhlbeiC8jVV9G8nDi5KQ31sb5CSvpIXGJ5zO6SIeUCpgS018
R/2SRrwn0Gvh3KYjSBnyg5zaiBkumM/DR3wYuOD8J6q3ThlW5asdgCkxlnapX0sN
dRXIry33BhNjRBHo/OHgYRJrasOGPDIMcgn7Ek5d53BzRgsyD8uvFiWE9WAa9WKw
SjUFJjJM8OUs+P/QE2RyCfvUKzgjEFxvk/3VN9dyDYdMz6bkFB+Zq71hTf4DwvxR
lH3IvSLEM6aY1eBDH3Xyt8EgdnG1bhsEQzmxCU4RvFnjhNen9cvP2H2pBbTWQpdG
yLhWUXUPH358b+H01KbJeakAvvR0qCP/8hdPIa8G/b0wvuQnPK/kf56B2itM6JdV
QZZvk74C1K21zrz+KPlfq12CxP9jzN2VCM+kYmDZW2LE4L4M9TnE+teL709Xx7l6
ZdUHKUwM0+L26BUAimZkzR6Dltal1QNJUQNvEKxizm2XRzCv8Ayhco+BL8S2gqup
FjCOGsV3onEejndgGrceprW03Mo9M1TiPPji6vYHHbolaj9ZHnFdMz3B+eAp8FcS
XfsjVV5IE0ZDkVod37h084PrKPEBgTeoGlOsWInCI7o+o9O2n35tbBjlcyMPd9j2
SiTMAaksvCV4Duiz4USsyBKX9UG1oMiNi55X8eQf2iQcblkc8ZiKMZTTHKS6fdqg
ad8ewpvIqsDtkqvmwQrH/MP+/hC96IdoUZOkVilHNp2VP37/kgZSMwa0LHgypMY6
VCHWHtogFJnk7TQaHrmOXyKI7pLqAmJns9JkzC/Ljy6dvGw54dfFe30hBEgcqNV/
+pgSRwcL5VMH5eDS+yFwZvZLEazC7iWBdehZ99S/In2Pi40mwGS/0jhb3bI5+UyA
+ywyB51pfWPNFgh7zmhrZOTS0V3nTn8FlwjmZIgDChjYDZXrzzr2ASZrEYeh209Y
4Luv96Fcaezequ3/hLoQ4BtJun8UqcmUp3k3/5kpNWgd8Zi5Wple0OYQoIZoS+6T
E0GAHNjSUPL2GxhsPU9PBtlH4lfUcIjgrsiE7ft6kEgMaetmzftuGW1qFVIVozgl
o5kAHfbyJqGEw33Cv+MrhVm5lDPYAm4KzgFdPhYyIV0xhy0ts7fr1cAveE6ANCyL
Xk1SKKWivsmFI8qfFnETLaxLTYcw8+fSYoOLjJLwxvjxAmZZgrXS4qG3pfexXyWa
QtTS+1Ey1EnAkbX+A3ZJw4qtfopyz05Wr7MK/dhol0lANyyy12hBuipjfJYm+e4o
9c6a09cVuaLBv+kVK/hMkpK5PyT6DOWYgbD68EYGA3OU4wMIZTjOasoa1z2XxbCL
G0TA4KrQdvMY5386SmJAlc6gGigPefpJERK15G0Ypa6E+V6g3MF/yWPvYqfFJo07
q84legzGPgoT0zv+proFiBbR1+XovjCTP5ypQV5ZM/Jqv8FU5LUD03bcglx82G2F
TsvH3LsXNy3ImeiMOTfePPg5qHlIRmaZl9K6262L6ENsUSWS4UmCQ9dHjx73OBeR
g5yiGr6/VNVriygCvctqfHCCTiLjIW5/HvaKZ7InrQS6k3VH90PEY7J3vSjzNSZW
d21FlW3mU6YaA5aIaTeNYcDJgKd5352eyxneigEhNe3oV4hVCLJOOrf4IU/uoiHR
77q88MBHWas7LuUJyddCRes6L/7/tCy19R6iyHDxfx6aDvn+cbyglr6NHhe2k4x1
Q9X4OnyaNM1/M34LFXQWRwLVwsMk178tKA7P+JP3gv8aBeQ+izzgvnfiF5/ISZu7
18mMxllPJbXMpwh2goanq6kom3Ix7MLu56dbwy5tWpfZT4iMDz6sLn2qC8CcW1tH
zeVnxR4pbO0sZI3MRlfvpuVNvlVMziKIXv+kWtREUFiBvT1LDt8mwq14PszHh5Ly
1P80s5gWsb2WQHu7flWLFummn7cJUgcDHjnO3ZEdS/xz5/wkNv9T3YgfvQCVpVee
WzyA6YQ9vOw9Ye8oJnqJ8H8ZsdxUnDujGLhoHNeNUg8hCspnU//T/KJjECKJ5lWo
KAQLR+wSVuIcRkdRotEmjT4PxYYXHFQAUm6F6ecPFDyo4S9ZgnQfqmmsx3E9Iot2
JyaMHCjBiLPubTRjY4nSMSY9/sPL9Xc05ZzUsHpLfywPKDivAZOpYwyC+k5WHRDU
5ikZOn9VJshnkq+/aXEUhRRtJK12Ddkd7+vIUwOEeKWoSYg6c4LQdn4AeJya+iMM
lNgGObhKOzJp1Fyu6yMWBDJ6wUK2oe/hu91g7QMkC2SsB8MeGiYFKOxamKIqHth2
idnYys/P/AtWxwZJYIFnvn1OV1gn2mjtBE7Q+9MoZlnk2yr3vBK3c3fwG1J1XkAF
9hGnskKF0EuSjDr4762ToFlFBrAuopY6oZP8pVABNnucdkvmn/8cZESucUuET1uJ
EfzYm3zw/4KCCc3VPrOBrR39SrQBdALGppaZaGtU5LVyuCJhoj1eRug/sr87Rq3Y
3L2cqebzQbXLxGdwWxdT91Rb1FVYqrjGhmGayf7rKGI7EqweyHlhTU7D/wDd1QH8
UKHMQuoMCSRhLdNz2Xx/OwKMqcojp1oELz3ry4Wd+h1b5y1O13FV7/nAYdmkrCdL
LTv6zuMKYBwBrrRfCUlg3eRt+An+vzKKLFqePnV6w4AAGn1rMQRXV2Njeq7GPEUy
Ei9oun+Itny+W+vPFEEfeEVRdp6oD66++TDi5fprMjlnAxPyna75jDqObr0isL8/
ERlMSNr9+cbCC405uwBJumj8ifGX7ABHJUTeblIUsrKpBYO6saJae5IT5FJTNpdz
pwkGgsiTSqKHNjUlQ+mrDWwD6i5wufx87JeLg/DDvh0EsaXK7w+ZKes+5UblzsHc
hfa231AJrToDa2odEJRP+Uq7mdoqqRnB9aRXTl2dBQrlg8a36YdWdpOuBWBmw8jd
DcmGqFr7Fd4xDMHE3W1lBtvFypJ38ltHyd4GD58dLMjazkz+t94D8NL1N+vFG47y
3uTsk3wRscwIbz+HilxYSEgfJ8ddwoVgiyPIjj+LB1mD0xqDtDif1m0evk2wbaj8
TiX+1+/8xG0JRzaWbWz42zbL5i67upVnMpP8ofO/xz7Z/XwjvXtgBjGTIIxNt3iS
Y2GMPUu4qrTYuMWargCZ/s3y7JD2Q0vdFtd+jZN4p2VQVRobTcRfnWNGHpkYN/i9
3kGl71F3WSg3pa/E8FVi4saR2ViPq4g33x4rALd/CTyAtGWxOpoHCFG0b95XMf/B
GHDDUs/CAcTK3Z+wZxwNkZw2OKyWAw7zG41FrZTB9xOO+gEAzTz1zK/x5Cci6EET
D+bPrC4tJhddFgzhSdWqpYCo5xC/b872BMxBod5WtvJhPDwmyByu6EJdxOF83UzZ
aQF/Us017o97b0Drp6Mr5GFV8kMLYHA/urYhHFgmK+SdWj/RHMRxqtY+6F4cZ0oY
afRDGKJkdcNy5Prr1AxUN2FKdw1XrMDj1CquaPP0++3ivbsfB1WmFkzBAzX+0G73
X/youADAVxT/e1SLGGaj4n+PxnoraIr0myOvy7R0R8d6L+7pxXi1SleEcOfwq4bp
qi7IfIhcT0muqbNVGO1bG2rYckZBC32y+NFFwsYEvxlUDTuwgijq+MHEzLdQJNz3
bUohnaYwrqsZez4uIz6tdqEgYVa+WsdTsa7Xifzqy7ieBVQ40yoq8GwTlyhu/gEh
j7YLC2DOTKLrWcecZhdscUXJFJ6HzikzkixN7YxHGQGonqiXI0CIsXojbOSs4k81
uV4VK1m605lxgv6Uhh7FSvpJWlLLzp7UIkDhAeW5Gcqix9UElehdBV+TtpBGdfUf
mWjg0wcDM71IF8V3REgB5ft147+ECMF7rqVSlP/QV5rWxe/X4UqBPfJrYTEhHFet
/nJHGcNtmKDcNWpfhnPJG9S4kzx3Nx8ZvJw412ttRb9fCPo22KD1MDFFy683gzYW
1zRkFRKmNJduz+xN4CVTaKK21D1+pW2tkzXqU9aMCZhedLSavSk5NBaTeIfAx14d
qFwP3EMoAsMbLvJH0X+RViOfqEBR2T3e1cFdhfq4YHI5y2o0xOEHEVK1IRiqwvMx
zdaBLOQW2e6ro1cn49GjULaT0mSxBZ2mpjKUK9BL9CIEAmeATUj03D7GLjwv5Vu0
1BunDLyN/kzeUkfqy6F5payRnn4sGrfTIezbWrwgw3RBBZQ2sv6i0gQz+/7Cmgi0
EhweFJh8Nn1lLsqcXv8TRShxc6/yFjKCdMowEJtUL7VWgdTtlTrimYxEmvA6cEXU
3+daiVUnb/Aslsa3PPBcGX01A6zItxXN8Pn6Ga1Yjeu5L9D6aOcVwSEPSlTUKFL+
G8JoZbXwdiiLljEySdWue2bhzbp8dKIs+e06K7iCr1sKsIf1zPaLXVW5bxCQljso
UlJHZqQ30dNtEnPPH91P+dJpiWJtNzs0O2QY62tPui3jTWzgMqathR4S834uopuz
etZPJCR3QHwIH7Bm9UrtbrO/pfS3rqb5UUEHm8RuJyonUcP45LSThYCCFVvxqtpX
x7Ivg+MPwAkm8QsAaQ5i0zIug2082HpphhOOzL1Mt4Iak6Tz8+uonSh9YMIOk24t
PI885Anz4sT2/Lvaf2/P2ybPdNT+LMb6ji10a4r6xXGAEvqxe2+LqRpgUx5NwAJR
pU1ofXMdnq43dUzgTQSFJuD0h77fNYRSMvhL/L4AmtmbQ0wIsONjtdndyXHk8gOI
6tybcqvILVJoiELbvjCDUquagjJt9ggzl3N2xbF4cRZrYOyAqOhrbINKa8/xwcFB
GNVymTI9hzmbH7Vlzc4lp1IEsF8zQmyZ33AKE8nTjjH/s9tmjPWOSw/gQqnHIFPd
twYkbvN71/FVgj40RtR6lwPTrpxgF4+B6952XKoh4AT6L+eFvsluPb1rkCylQ89N
PhI2+cTVjMYxLAzVmlMvNzmKmNc0nD5JLhyK/44LXELj++KEOkzwPtyEoV+lXcEq
ejrYAKSLvx7sm0/5/1vQ111eYkifrnh7QLnaZ/iAJE3bmIp8AjxzIo+nA7IeZCom
6i1INh3THQHGWVYLFDeYGiCoeWj6nbEu2xZ2+azquL0l5FqKkHZDa2bzfN+RptJE
`pragma protect end_protected
