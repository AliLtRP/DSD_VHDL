// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pGk2KBdMvyzzFxmnz8o8YXjOsS+mwhsyv/UgnxNI/id+ULI61D5oPcsY6fpe/qQ/
fis4R4YXzedib2B7Aah5kqYqQ0b94c2r5PZbSvsJdn5ZAVzkB5BX51S4uTVdnOot
fIIh2OR1P/500wA8jzyqhHsY5KoAbGEbKvT0fvfNfDc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42432)
7gE+GUHVzfBDxPIiGxTArzxMqnZTn2qiuipmo7ofaA0vZBcbhJiGGt7gzraBeS64
eRjm9680hzZgfEWg1IDuSG9kUJ/Tb1/mpfpOjG/klFU/9KasrqImZBYUoWMhjgf2
pxy9lu4RPupSSgsfXEjKT5fG/Sh6SdWklfLICtzjJa34U7laA+7hZdeX/ID3I/mT
Z7AbK5hlvIETcxcPFvpQdPesVQDUeT5oSFyoIZl4jyOf8hEmC2/eZWmsNAwBb9cq
dEurmQU+mokRA/ex7ppcmVJ+ZJ5o5oXLw7MeKTqmB0hNdzTCFbLOSCOn5vbw2/A3
ikIIUx6qfI3wy8s99szi5efflflbJ2DmQ0eyrlhiqNyaxOIsX0L0FWNDKRIqaML+
mW0ODj8klRCP0+z2iA33+3KHAriIjv90DXrNqUDhgsL96HXYABfuGJuRvH8hUWO4
QZ3v08QEaFMgJJCC5FaDaoe65maHDYF73zgT+5rmKAomQhZ8dhADUb60B0hRIVcc
ikhTv+Uz9/pZUQRgnptcaVT9Ngv8CGqn7qi85twVKgJfC2DIdGrl9a4sSZFyKVNN
LGiP5vTlj5mFcD/7TxlWbb8QU2QMqwCCKJwTZcyiXj6BiusJjNg9GYiee12rWHZZ
0GW34SoHXUPThRRyCvpjPK1rlpPKHaSBtk20w2o1pMQSGLM5A0bWMTtgyvKnj0EV
jFckQY73SF9cu1DKDpCfhFoEiTU8U5/WEG8rzEcKvKSnUe/g6ya6T/48xSG2oNWu
Awk8+RC3oWf5xre16hduHfFmLMxhRycr5q0knm0ZkIzMnxNDDlg6Lf0yUaUDBeHt
Wo0i0UBp6xRGzlsW+JOX80KY8jq8X2TLKdHenF2aX7Ml7djz3Rc14mg6pGMpesbE
fEwbjaay+II6NvK49qvZcNmEC7pv8NlAdBqCxVTyQfrv1oWwWhJHTH5BS8Fb2k1b
qjt12K64LxMu95aFp4FagM0h4RoETEKqVmZeQO+vhu5w0qkPZiZPawwHKG3ogGQJ
0+NoFzsuYZe7iy90bTV97ITiOMAjiW4gOxSVO1EhNY4/WC8s1mkmQ2K66iPJJ602
W0Mg7U7kFS/YtYV1DGyotE5TDO/Q4yXw0xLTcn8WIlnhzVnoakU2lIlHarllJ7cP
jijzlEG0lSG/aD6Gbit/I77bw4sq9/c/TyYry7Hm1PgMJCds97HCW5Gv183MRI88
QmtIpixqz8IwFivGkaxnO681sbB/J4sDRN5rt6TNmovi4NmLEzqB4K/4nzgTCyZ+
ZkJmoM9Ay+spZAh5pfBEsB/hr/uUzNuRC5cACrh8sDeqQJ/YPSLNhgvMDD1zzCH0
Rcvts60H4KfqEyEOyucKtd5DpQGF43CP4ItcBxDGcv1V2X1QGa6nhAnsbhcn9OML
jUBYxIfOzg+iuScwZYCQfJ7sGT66bGIRHibYDWjMfaeXl8grtvxWl5kB068SdZUP
zWj6B939wJwA8i8W+b4qxMDQGUl7y8RIClijI5M1amysemJ9ksy29/hG6JofyRAF
vpx08lgHvS8PBYFMAVuv6ugfcWRieLvep1d7qAGWNUEd9qbwSacI+Id0JtEroDcg
pwpGPsbslNk1astHVctcQY0hFx8rvkSXys8d6h7QZ2snBhYMeMOyf4/WpB1xvvxd
dW5214/oby6JPT8nVqaHbGCrgXA1rj4FfpGJO9X2XQpwZ47SafNlYSJlfY9EEhlq
kUouMXY1Snk6kng98IaqesiyVl+9N0kn7bl7Wr8WUTAf+2OhMLxGoQqhZvGGUHGk
ysfuGGHwromlQl6LOUjaTnLtwrcdCVGH5rylyCQ8gJe5TqHSsYAxTwm0rDcKIht8
AZ7inb7BFTL7rMufvSUrj/JO+/RMhuJh5PPigfb9cHWzWpnDA/j8+vRrBaUgNIca
SJhawTwjd/xYvTA9wVsIoqzGbwz15p1qlECJ/iqXZvGRpqEOXC/Hymuiq3BFI7gq
rvVXc3m2Cb7/7g4o851JYf+jGZVkllYCRnswl1vv3xICrBW64LtUkLFqKuv9bzvl
rX1z/ruwTcSQ4/yy4XMnv03V0WkZeA0SU/NOC8UpguCJQFe4ZDdkUwH6INrLyGld
h+atfBlMvuqjkAmdYG6XbF4zfFfkBJN9Grq8bS+lyyoOk3mc41lrjrQbUYqsr0Bc
Qixr8YivMgjcixLqrRIwUcWhBi3VsxkwPEejKnUFBBdLP844tyVJEp84nWfTk4oX
+hO/y1UEWExr6dXzEo1eceL3Y8NvN94j00M31T5C4xgK9A9M8TAfcL3vML21Tcq9
U5AY5zl4R/jPoWri0efkUkiux1xuRgrBCKH9osm79MuEO3OKMqqNBI9k3jd/Z6Jg
dq8siQA1gB/su+33fIBVhPbbyMKqUGxRXSQPo/XFldZmFmGJTm3MUmwDQJCGoF+x
xNbqctv5/9DH7Yju0kOpAYhNEtFBVHq42rXyijLj06nQOWDqjO6xyERzNGv3PF10
Jr6TpsBspnvKM6Wy+9AhlY68Nel0o0N7Rs63D55iRNUfILGE0/igBwDuKmpX/qhU
59yLXfE54QqMqAqxrVEgjmLV571DkkV0ImU8BPidZFeISta1GBlBwBF/U0qavRxo
3Xz2XFuNbAyUanTBWu92VBcegufjEO3kO+E8wfDQYWRW+bb5uePVljoRU5Fl0Pgw
mDSuC16NIxUl5Zgnb7kE93uZ53kyGvFqOPL23nYUosSLGjNQEvPdUPI9HKWXkEVZ
RTFhn0bHIKZu2aFZw4GUodNYOnnbP239ROK61l/jh/8K82QGhGWdNX19YRD+d5Jn
IRzueNCT+Tpuwk3K570q1dLqgvkUsj23gjQ0RfJf8hcth2LbkamYIJNr3kw0CwmV
Nc/8+pYvwNXHSeU9s3iWGOZWhJn9nH20M13S/9NHFE5YgV4OztKRj/vsvGJ0eTw/
VYLUCxPVADZ3IVzetLTIDLjkahcsA7Bu85JqTYOQ8JTAXTy/mz21ci5Utd4qBDGb
e4MvVueUZIcO4S/M8lGqUo8CZ6Ek+MOeN7vdeC/JizOYJ9nTFkv2yFuWFukA+wP9
PHwY33QbDNFGaRbdQy3pEksyEY5at9meGlmH2qhFWDsfPaMho7gS8gF0WP+h60kn
O1gPEKGDRYKh5K3Nmn6Z8AOl3d/Btfxh+9Ih0idRKKNiYdeKG8p40CNIVTxjlmzu
NTFtPulEWxLcoSwKd9zOUauDzN1dWNnuNYPJnpQzZlQNDGBRSRZ3Z6KrLebIqbHI
bN0Jr0tjgkRe/79S99v9UcbYofmmunwpbFHNfQGy8nTPw39tljUGDV1qTLFbKwG+
7DzDZ5SDI1msKup03SsiVERlQ/cKnpfbjuxgQ4M4NEnwE31KlldsLLFNkgnx441M
gL+4uJpxdFjXT3J7qET3hsCt63atfqHnmc+bLS+5egdyLAu32JHeTxIethK7MO5j
RzJh4QRYLTUnbpbVplEO1vcreyEC1SBVslPu5cHGach1gBOIj/0PkVp2MbDNncKf
RLMMkMogbkoAEpglvjUT93MjTwwEfDSdV99L3fEMnEKTop6cS0A2oB7kqzX2G+cm
QHwHSVwXqY3AmQvWLCdWs012SaTJOY1tNbMyD2N0FzXoYASmPiiXXlGxje03hcEf
4cAJpO/tupWUDMhGsPlEhY875llTlz18HWEZpD+z1/1rbxJ/daT2u8cfGFxOs0OV
TbXgw+nF1+lmCjueCpYQQ/LgEQ7Yb+8EvJ2eGQIqeeFpmfQq4cXYtRsk4aHiZnct
udy+h2nKZEWBNZzd0g3GCpuu9dRCuBvqYp2FN9uI6Tb6r6nd7z1XXcPKaIla8gzq
49Q0Z6LJ90zr4mS+TahKlUhAbNqwnNTCTKlt42S8QWkCEgX7TJ/rrrL8O04cRGt3
/r4Y5Qa7Ai2YjMpZQylr3TpiXHbmBW67hBUdjyR/ysmjEsRoXCacQ1XVoG2Rui7X
jBQgHrEsIo7DUDwL+RQ52pwhOkFSuQOXRJn/MGt4eoCAcIWCdhOwbO5KAKR35dy8
OLpurZd9hznkYLNLmR/G2Rok9T8Q2l/LDY4PXpn+lquxyVSZQ83uRTrjn2FWWJ8C
ZG0UY7h63ZE9pjg2lPBTolHjwL6tnJRFga1wmsHaqdJpIz4AgG5OSUawMXQnXm4Q
6Mf8zjqqGDisCCM0U8IXTLoso9SbswssLEEjSFkAGDIPiURHlgiOr1WBkV/Ojgzh
EvZPfmDcFEHW42qSQR8E+rgxNHTjwIyr+EK3z6umkDHsBtok+LniW/fQgIZrXYQe
hhtpRpzA69f6hsfkRZLNGhB3u7nRoLWI10n7h0it8NQ9xTLyGpxfwoiKwUrUx3Ut
O+u9uyTYo5F8zkTM2OT1Oo216AKZlCF7JLhAJIWzt4VSwHiQRC/mhsYEdKc4CJmW
b8g2n8dXagok+kzC9oYQ6Ols+IZ1jL7RZimv2INFri9OcIkNN3W2z0MfPGM6Aa4j
GuNWLwxIAYCRaeRSL2EY0XqQCoYTQnwrQ5VRS4apr5ou4GQGbePIjnxNwskBq/Nm
cc/fqsFgp5Qy9CV0aSMpSF0ZgCPvEPoNmD9RVq9XMYP49JKv9JxIJQnqTZPIwpss
YzNTr/20bhX8r8vVwRb5+FD8WV7rg9ZE1VkFYbIy8Pi3esmJXrVstpkPMurJZSxA
fNUeNBXxSWG5mE/mWR4xwXTKQYVfYoRahX8EiEU3MFlwxcjKcVlp0BZDdkiRWw+O
1EafFeeio4tON4GA52HteQKTCXVHqQVSQNrpflz+cGKvoMiigU9QVn5ubIlwh/rg
cYz4KjhP1FdZ/mlyX8VSJM8gQ2Vl1Ep9hbwRSU2k41sP5ZfYhDEKhmPfbKH+kcFY
JyjV6+B7Ro21yEhJYs3YkuyYnsRcfaUesaLhblwdaE4NXexj7tDtZvHJdc8tmU2g
4fb1KnNQj83BrgEoK6OvIw61Lw6mdtxRIU81w7FnX2uYIzQZcrdIIIawUJoT9LTL
GWZU4U5Pd1+p7hUTr/1B1IrcYhsj3guuQbP83teL2XdmvP3uKwHI9phKVSzx+Vo7
MZP1sgOUoz6up9gz8d8wGtbmtEpTCYOyumEzsQbZdGx+JVDsxqFxjgsf0zJAcpmG
JmswB0fiJKF8HjppYjcdnaB0rn88BGbvUZQJtxoGTdsEiLTnlcaAPe2vHwQMKXBw
k6rZuj0Fz38xsysrCCXwmOITGqcZV0sCaCG1RUuVof1zdT77TDf250NIEK6f9Xyh
8kX+F7x4EmqYBTIRSmK2e+qghbchw9I7v+GGvsBMTPAiXiW5Km5NEV65rC829wru
cjQRK8WUzA2UKQBBqfurgdOD4vZ/wDANNUzXfb8EustBUvf0fCfmzCCoXMyJS5y6
O7MClgCftzIfL2hmniRzpZ1voBJ44uaDnwAyq4EUjEMCOOupgT1tjWcSeBBq4sLB
VRCgPn7POydeBxkUwFKAOyortjzMVsNxaMzzXuI9x4erkWNHcgWbc/U08O1A7wv/
95gSawrRDnPmjbI+GDL/QhuBBhMTaTf94UFHjWO5Kj0hgIquP3HVPZcgRkVnR3xr
23zX2NX/kFbz/3RuwtGQf7Wzdw/nrv+D6J4b8XFhV+RnrcxeU3hfxVpOavhg/N+f
tONhM5jK9YlaUpmkiql3SIAhHXYDydSIONc2tlXHz3ywOQGOoVD4PoUPyTD+CrHi
/8QMvBKEATkS4cyJxwEocpD6iLlrpU9/to9ECV+oYbvKTh2G3A4JJvPNsz6OlN6F
CQsIrPh7s2OWVGoXCH9D4WwJ0fmYG+qR9X11OO5em8Vf1v6Mk4d2pOrL+UlHHQCr
B8OSSpZeY9x+1Es8qE34Du+NyoWjW29TTBYYbkJCtID8xO+TcDXyl+alGv6Sj29i
Dfn6whGxcxJzBZTheE6Pq93NkdWt8wqNTDoNo2Mh/+UTCkivUGMqFm+e89MI9STf
vYWKjr2pm8628zVd5sguy5j+bOPTdW/zCak0NwQPwZRmATy0A74jp/kNF3wpPtQ8
ypeIdoE6uqkokou4gFs3lPh0lPwYtnyMN0QgKQFu2S0KvIKbsWZSgb/vUsca9YZN
+fNXf09pOBLxNs+Brnu6fPzYEdSrFUgmxH3nWuI/wc4BxcAj35NlaDvizh2wqnk7
9itmrY9VCGXwdjYEXy0f8yIvnaXv/XxFeWtdZai0yExeOjmvHerYda6lXdK2e1xZ
J/hfXAxqPj+Ieb/L+7p3QX2T6dbG+8tq5lO9MiVGas/OhP3jsBuhn9FO0Yn5y+Iz
7Hxc2e8vz0wDcHr0vc9wiVc46dBcZ1F5/+HyhXcuBQseisrNwVCa558sjalU1wa9
oe53yTenGMoIwHbv2qMe0XGeZ/GCI0DQWtL0lqtCXp90lqS7/08w0i0Q/1cWeq3d
ERw34EE9qwVFS5ZG4qmG8ItqY00FJkWk7yKFAeZxrIMEsyUSi6YU8J2Z7nr+kv1a
dNT7ouM/r96/Jl4ePMir0VPn3sbUyGNALRUmDeOZiKlQT8/PHK3LdIh4welgxhN8
2NTSXrm2IXwl6JKGKpzMubBVddbSroBdL4twSL4gOnC5IOKz4j2zD/JW3uGXCr5/
A0dXZMhmfJQHR4pvFKuXocBVt6ydqdk8Zr0Cmc2PuNGvvbIrhpeOe+dU3CxPSznw
Y82C9JZKkEUvZqRt1LTZAmPJam8CfzQpZrzPwTJ5DzxKTaljwC7smkf95XUx3V67
CWNfH6YlII4WUWIf1nMOiUwrCrxaz91JdeGiEfqf2xPqL04iIBKRCnp6SrLUpvEr
DLqxyAvPzwYUIW4xDLkvOjG+AsGJefiA4nNFa/dYA0/hXqKU5O7Exhj+kTpAD+mD
m6UinD7NgIWGTUBfOG4pHX5R4Iwuc4d6T/X+BZv6HbsuZ0adGFlJVCGUeK6x2d4u
jMDzJ9+gJGFkGULdhqhIFz3I5hIa8liVhFNvL0+CdcCfbO07zB9QeuYPKttkdd80
B/1RlocNdJUBX4o+VgYlVbJImd+UkaYpXOmdIEqB4Z9NuLSLc9OeXlHIL7D2aGBz
lFAP1p4C0ePEMDNXHvbDSid6GsNCpFOMZ1/oxtzQ9VDR7baDBesSSwD/MgrYKyvM
UDydwkdhPEg8lC09JXNtuUj+S/GeWG1S0wxut4hdyrvv2pJpox3Rng8jLHnYWZZ0
qhogpboK2GGv1qQCiHhzwqyZMjgHaFNEKpfYl70/maw4YEHrlSfifg4V60NH1/+p
pR7IHV6acF987mIOVam//bGk/RYWug4+aXKYrF7m/E0rmxJ/nB3OKGBiKDyKa2WR
1i7n862tZW46U95GG10Oc2iSH5QRCWFGm1tLWXA4KY1ZE4zi1lCKBaKSoDopsmLV
Ft1pXdEWVrFstXqzCu5/0iAPQ0GY4UPpiOO3YrRfM0hpw4xkC2Tsc6sp0P3v7BDn
kTYj3+ef2b4Hcezm0dMCmbiMlrDAGFy7pUKJ+RLIShBKmmFc9rz9dupQSH1J+QOW
qd2Tj4sm+FML0uiODG3MeTOicVsT8SLxxeGujHPVTPWk0u+O6DXfPDs/9zJcqukj
ikqAlerqFXKfXyLDEaiNf75mrAe3gvObVqYarc/HIo4dov5zTsiR4RLs2npHm70J
qAPMDBNgWjmBLk87u5GLNfY49zp8dExbpDDv6RmUwR/GPD0tWjnaBSumTCC2+26s
TiHe2mO90kOoiYUMJPCEHfrHCNTCvCiDWyPIMpx7EPMamuxdMvtE9ELMi3zFwya7
DBjDnwvhKMv/Ga1RoH0pJ/d9g7OGy/A33lRv2lRjpVJ+of1TAyGP9GgrnXkvXfAx
AO16j7HQZ4s4uYpKCpmeXizYMehVVN962NdghsHh2FIJmo3AAV5wJoNAzy1TBBas
ut5JD9oy1VgyfTvlaC4uEg+aEF7VEAs1Xr/Zid+jjK23u+qaEDSZYldgyAdw1ly/
7f8KQFgBPnNK5TBcLHZsuxKbwLczU+p8yG6tEZqF8Mjwjw6YDjbjQ3Jq/qXksTyA
ryb3BbkgcT8tjZPmk5ah+zOfCbqfHaHdCtIIR2yY0gFS8o0XXJ5HUuyhxcWrJlDW
VVcJdAN/fvhkTDs17zl+WaZpAtzaQyF4aka6ze85VXteJ/C1+d0k5pT6jwLwjiAk
fg3XlWR7n5ayYOy5g3WnhRtGrm8Uxu0SwmcZxIpLHrQu0l08j00+LFEnUHUoFMax
uJDXZDtX41LcDBCxj0lTLKiDzCSCuDeAHhBXNj6Yw6nboVjvKiLYYTzSWZt/3aNG
4ssWDgXITaGrKRaoH/I177RJXWtIuubqzSCZ+xxptSkaK+TWoKmTsgTk6iPwtj+h
TXNbyhR4rVj1csh6Q3c3P2Y9PBP1IJZ8KVUfUPFAZki9U4bgeJwapaXZv2X4uqVg
TbqGMN+HgjiujUEPkMMOv3r7F+Zc4uZ9nNbeN8pryjyCuI7c200pg1CZiW7BAehU
0xd5Xh9692yJBNEDUDNAUuIreXhvQJO3uE2XXI+yrzLJA6/ctSBNv67Gk85wAvwL
jOJDDtgiltaTe1QoPRW3f9+otpi8IWfIHTEwFKqKaBz6DzFyMCorAvy4cPEuIeKk
uFjWt6Vav7xP3dpW85BvdqiQ0/Xz99cxivqQhVFmzvCWUOuv9ere06XaqhU6FqUz
5gGGNxLvXDBhs1kyuUkI0IwQbbAXW0Ea2Xakm1/ZnT+6pX8J+pJ9Mir23A3TaXut
vdz2dYnE0lWGB5RR5unkzSTC0bTtILYshH5CHDVlW3zNe4205cDPfauYpDjLrahC
Gs9AFz3Gn/+cmvt+8AoubAKfr+7jAJHTyXwfFjuMUn4wb3x26t24babpEo9xAmWM
W//dv/gfaUYX8+3pmf6qraLzLt+zyY63ggLCHuC83Yj2Zw/PMdCpVOxVn5sJ0vAB
tepxxRN2I/JO6LLMuh3rXm+Q1MR8RAZDY3n4tlFuge6VAZb+AuRkiv93zMUtIQU6
MkbUpHpQGkZIrrarnLKXgUyTmo9OqvRv0cSoVy/CLFyWsH4yqFt6dRpN2pT/uV0M
wKoMC9X4SYFiZC9Qyw1YwTYQyizPUrSghbgEChvoelB4vyCbzBWCO7PP3PABgL3j
+jIj6VDXIVBQdaarynhCDwhRFZLQqniBeXqMCHRu05wtlQI+0GKMxswawXBED/WR
vv+fZjA7uqia5h+okVHHc5wWHGyu3y5SKE+X467v05hhxokCLsq3bmvHCtnemCua
8CItzh+7DAQCbPHz0no9wvvokw5PqpeMdpmDmF/Rd/O63tYYfS4x6Q8njJH+HbLx
60VGbC0nRg0a0gQkOt25Ktsfyls3aITn7ASLinegnN2c22woZ+q9yBkR7fkYFQ5x
Qt11HNlQematI/Vk/lh5RO8pJalAyoKE3j4UAHo3xgMwUhm6Cv93HYj/Hn01MDK5
sJw9r1NGJJwZq3VYfhnwgjEWLD9s+P8kopS/xD72mGexi6OfL1rb7LPxAc6c7mK9
FOrizyrJjWoB6VUC3Q1hTPIeSOZwFH/mk/l9p/zpbasqYbOLIa2vCkl0tTYDJOw+
ehDeRC7kuVhURbXRVlhKnUl16uADC36flwnh3yqMm6wqN07NKps239WNotSV4Npq
2gtVM1GP+6ZLpPW37g05V8y/wsQqYOews6FxvZOHVcgTnWVMOsRUUbueH9yW0loo
v0uRmwAex+mtF15TYlFZY4bBERBDddTJ3IWADBGLqtaAuWabsiCfB3wByEt7d5zL
fv4KqVSaIS14kDvvU4y7+zAkQFNNvC63z0hu8UQigOTfrsTsSKmuqgNlTVfJE0Sa
xYwmX/MjZVCP4QLCCbJmC6R3rnSpIGsnYgKfvmri4pI0mu8mYoXO9x1rnW2Q0gDw
B0bzp4RkDtMz1Qy8rSdXipwrFxOOL3yEyjIEB3rEPQyp/Lb/jNPAb20C02YEKHzZ
UPhnTUQt+L0PLmiekIN8ijXkWscaAEEpZc463mtxsIE0yAe4iay76JZz+aJ7TQpY
HeLSTeuDAY5M25JmVyyagLG4yIOkVbOYRhMm8EpVSVF+SHfXsVH6kSUv7jMJuAkC
ZnYwXYaAaJI3dEUzBQtRkhswYbAvooJWMxPgInKhBehzzpqErQ1cgKKcjmbJBnBK
eAM5qXwtor3DM/2keRT3JYGrVt+Sffqyys0B8Rr0N1IceiIcmoGo5Slaaxbq51LS
fOemJECWTK/OSR5sQFBpJzv2XXLKpm0o+Sbc1rTeVeTCfdOcuIJyugA0xSGALA6F
TwIpkmZQmN+4UrRqiL7EEZuAHjU/CgoWx7+CVMF+jyzAs+e8sgOWnxdrjDTZEXw2
plXZDNn2kZvBU6yysB6bD6NYOfI4sU0FqR+LfC9a1CxofVPo0v+ic/TWp/EpcrpP
b/0t1MXQyW2dKNmttwTGmWjYuqCUwDw5LsZKrTDI0fl+emnC1cf+LiN89NCodYQj
TP5J7FtRS+m8JJhRXrDQr3ydvXEYjJpjW31lCBFoLW2IOkIi+VJEd3sSEKRxlsXo
TqhNWTAnGtph4tQKQ9354vwHrAKXKkI8HZPRkz5hJjEeDhjQWX84N82YVkqlkLbs
HsP1nktjKJVcNZhrOlXrNkUfFQjhQ/HWMYHs2gHDQ9TzKrpZeFV1dgCkBttMqsIe
49Rd4lBAWIG4QOJHHmc/VR9zsx+LmqkO40E2wHKU0Hlsyyjomdcoa/NNFGuDhNk5
BYhcaNL93DOYMP3Y2E7Qd3/y/FU2auC6/k/rLA6nmI6mzHmupxuF2tQVcbv4ZtiS
aBKLmcmaHDLuMYrSv+2Mry1Moxs5vKrxWXHZriL3bR2JNymofiWyPTPmOWOdQC1D
NKq5TP4UjL7/2bk/fzCU0OY9OhjYgGxeqyjUCtHDmgicMDJqTpJ4JGQ28L7w3xdu
crjGmSuttbQbxx0uYb1inoUqWRbX8VJmMOH993lFYvtYxLZS6STWBSL8Mg2PPOPl
hyyvSXsq+B/XOZQCcStyu08bB/yDKvppYXI1YkfxyMIM8S0l6q5uU3bwSkWrtUOZ
SWp6i56Vca8JLRsNplf/vXj69oGoes8fEhNGyy17bO0vZKe4uoQ0PQVseNA0BufY
b9Pu3ElaIClqLpy5CTOWHRSMls8eHSvpuTTRv8J4UQ8M6F3yz6pm/c414DOfr3OI
HTOqsJYigtuR4rAl2TL4hanpayCnEfDGs2hJmBaa8sY9T+wpqJLr7tMLBGc9l5Of
M8fAhHpA8jsgeKLORMWrAYDoFyHvzjyGVCFJqpiHZcLRDkergcMNEqLecIdg9QJi
hPH22+/nV9yzM7i/k+NxgSCI1mrIVFR976bZNZVrMiWqL0mAwxLMlmf2wCfAZqR9
knnfVFObsQL9diY9cTIhSaKBx1j/yLMy/nb7A6kVu9CeCIXmm0EUvJQ/OtuOC+PR
nrX2DvNJbve5Ny5vnLUpPxwBRsl+MA1OZbLiFGG2zPXXjP7LCxGBfPrwZqn5Kms3
6QYx6eOFwx512LaIa8ASmoAaBuo3jsyboS+xQIq6yEHMa1jX8PTjEQ+x1eAa911I
VxI/L8u1Ij+wZqNa67NbxO9QuGTxdWpojC8hrIg9QOrkoTfn3xbT3G2eSdvcdBqO
1zg5ksrtzmyFpCYJSSz+Pj2ZmleaxDQDUWvQOH9RoJvBJk4HTud/oE6TncjqRxx0
WISZJpf5xA+cvN39Uwv4edXpnBM4XtWLgazxs8T5JidU9TzCTMK4fhzxjpBAAtsn
DHaYAIIyG4aEBwc52y1RtZe+GmnPXJaxX656650neYOvn3YCYZ57TTncLrYvS3Oh
p8OdtWtmydrTfoyUmCHJelbrQX6yWIIm9hjhFefMKKB/n74tPOUtk6+qIpDz2h+h
5TcRiZTyPICwk9rrrKrkfNOZKUcJdrwu08eLxxiUDafQuDUzgD2p3jPLKZ8JJ9PC
dvU0rE5ragC6vU+9apsL/6z/+mzdlTj6rK8TC0ZdmYmdQb6nleugb/JUQBaGV9VU
f0JreyZcF2vPZ4No6bCF1My0XVFUyeMkmX2rMAnWqUF1HRZcCzjvS7SWtiDmaZpr
PZwXd3zQHxvtL2l74EXJX0oGp+nyYJJiicPvi7OPpv4GPJ2Biz9/PX/VjYqbpCPp
XBjUltcCJEzBrKn2p8mxlojwSlCrmYLwTNES+ZjH5Nh5alT7gal4BAefwIIPm0VZ
wVfU9DJEQd5HAZg3WinTJzxUvxodp+miRzyPhgPgkVhKjtnj3x3Di6sWoS3ssNmt
2NVbTmunYueHI17OTuHgujBft5v0eKG7OMKmUHa0c3bK1yqqu+TVg/a25AOZ2Bdj
ybyq5ZfgWfTbUOEpREHcS0tDur3sO6AQd+k/S1s2dpXegNgxzr7pj7S7CUh+gOwY
HjEa3tObhn50EkKVDP59r6BCvbivlj63PqqNMXzjw/oL+uGGMfKdUsnxOXbd1LtY
V9KuoQ1sUhuO5hWFeqQUn4NYTejubWwGZSYicXdl33pp/ga1cggPt5Z8GlES8ZvH
m4FkOO1GD1FnB0YOrHd3cwNIbFOM0q9yVtdB9sD4QSHZRJAbjZx+6yeUchafKl7w
ytn4HweSk8FCy0nkxgxb0Zs2N0j5Xz2QVZ32axOnf+ep9fo78Id6YVo9Uy0TkFyu
+hOw+v2IAw4d1F95hs1nXq1lB33dDKXZBRbPtmkYpR79YK5Pi+2EngBj0sayMXen
FmR7zWo7DrEUHIxVILJlh5Nq0yeIzwBt95Cy4tBswEMTo6bFfevqQ+UuEzIyEMq2
On0VCDRNY/ILxr6+9ZOeTcN16IV7BT6R8kjQG8NQf7Pi1KmynnLKQh9nTOll2Pg0
8MSQwT33oQsLvrrgx4Sf26NFtsJmTlkAZZlA3WI5/o8VyQb1SSmxT2jsh31Yd5M1
38o+PIo7AjRRyXrw2E25poe6O7Q5tQwEaBcpnH7LGSquLN/JZ8z2obmDXzcsC8Xv
bLNNUciI2XVA1BVVS1KcykLCFLfd6fxUHJMsocJl5rBNG500ySeq/dAdkWV+n7bP
VWngmSr/2XvcwNPWi+fGZ8uqVY4LeYVXO/u/jzj3xKmeSbmb0x6ZbpH2DWiliUk1
dZ5tV7EK0+Hy+GXpPu3sj7zFjNRVIAG+eWoWRNItoIhRu1r7itS6J/5S93Ag7Zzz
od0PakNs8S8WWqJaZ4OvU7c78JuWBdT0aDy4aGl0CjiPtQ7oUFZU+CZcNO34X1F/
zePiZpPi+1JeHWjRiaHL/caIUMW2gIFbLGk/TTGijW3PYqM7JHDGX5f3s8eDDZUB
NO0rnUBu5vkSkG6s1jMO+Q/2Vw6ykiTjvBWvFc9EjlbO1zd578OvbE63j8vckY83
8wzjC8lbQzdV5uYTwx5lbumAdceXQl2imkFtTwazFgaJJYsqdGEuD3L+GOupILHn
pR/AKPGG0EIK5ZKiZoslnutHy4SSaujEDZ63sKjIobm1vkUdOsMSPN/Fkrtrrpwa
0sqIdwioOeWC9K0f4zWcDR2TGdYgXG2+H4rjPESHdffGiCRkuDFQr7lIjsu93HXc
Eqn+gugnVjbiofEFh564RjPC6nQw07hWcbI1es3wCmh0MO0raOnMOGQprh6bAeWf
IITbSNnDQiXTaYwONn+CqVzcJdU30b+oOQMgYDTd/Yf/eklwhJ3PLarOv1evDhyT
Mm2fNMi1UHN3zbwsb8SgcGs6v2oaUIVLIAr0TX/0DZjNKYldai9herG9W/rlYTTq
cPBo+gFZOiB/TRv0VQq9uZlR1dx2uvFERUBcRhWoGEN6WfpdeGqYKhELhKf08PgF
1hLg80sOtkRlQVGlCH+kraQu8VuFkSZjZe/eZBU3tf1yZrv+qg4qLZVIcgtQXQLv
qoDYbkjp+bBlA2yn55L6b0w1/AiLE1UUXmJeht+SbSfD1RwbK/NCAOpoNPaFBzfe
Cij7bswSPVk6B169NP+OJ0olxbbLVWiiGmZ8xnfwb05/9vuqPh0WnQmQS/+1+clA
Q99VAk6H7b95BfmCuqb0qpDTthwMWNbTIZNj5JsR9NGJWOB8MHgH3hkRGWGSvwMw
iB7ndh3zwnzW58YOsc0z1puzhM501Tcpja5IulLmPpNC6sxSYV3U6OGu+SVVT3sg
h5tlpV9PiisrnjwhRjFlTRZPOh4LhcZBC1JbBE+RQKwndGj5ykNJTfKG7X56lF2a
SeDxWnJj/kQSMhQOf7B88uiIhmMD20fV1psPPmPb4bi1kAfYO0uRcC+Q0xupg5um
zcvoh5VagByVXruY0HkM8DTkfETuVeovulBu3NFdnYJjtPTCBkTfjKOahfnMml3k
UwLTDDdsRa87rEIaFyrIIC8uMQnSd9w2wNoVuLaGHo/zi7DdObC98/a7zt0C5fEs
9tTZt9dRHr1rDtHZ6+Q6LdYugNIP0gir67vD94f1NCs8J4mF61en5C1OkcyK+MFG
dqmKbagGd19uotuexByXwv5QDRVDGsUPUmvq+CPqsZfsmeQSJCCrk7StrUYbZkOu
HNj+8F+n6VzQlbUZVNZu0nCeSOZQikI3qNAosT3U4GA4/HEaKEvKmOu/FNdZfKrT
x4zmOGk0WgzNRNdKi46N+akakfN84WnKFSO2bcJI30rDIa9eFNCEQu4Y3z+y4bdm
TdwaVRfAszdPkZ1ShM88/mjpQHVhQdHAeY0VCew5YTsSssVh6EEh46TetkuH6ue4
9PEyvO5m2dkBtNe0ijngCg5CAKOTgbsm7H9TukZ8y9l00CM4GGQnTGcgn9NqpgwG
2mEXK0drqaqPTH5zjxf3eQB9tbsDjoDDwkqr+50VmytmUm1emE9vIQr3FwIk7djO
t6z4QBaTggitBPB2AWIUyshUFMyl8RiAclmj9O7HzeYeJxAo5i5PHgWljKXKH69C
Cj7qXy/+FkT7NooVIAmE6otGWCiFfe4mNLfu/W6ns55tvxHLXC9EmSIhsxxHg53E
AU38XCEm9AMyOrvrEIgYOKu1E8sqB6eO5fTgCsOw41VjeqnnD5eHyvGHb6z7dQQ2
ugomyQy8DLbs+TDyxftVmftXZLsz3kqzu0fEUSWnjwT+j1KYL4YGJAEy/N09mG90
2QSXCywKju8kXIwD1LNheAbcu0uA6Xxvo+ecDJ5vqA5/lvMBf6USC7m+MwZyP/NK
7yBLgN8Np1pHIrQXFdZgumRUgRNZPlRey88JTTMSMWeUvGVronuu7O3WxnBfVgzP
INOk03ShDTM1eutDkxy8/wUbR7gQ6BNQWFs+nBme3/+XxJiP+jVY/rkzM5d7bgBC
lPcJ2o5Bl/3O5IVPKRk31XQxY4CuUXnjqVOSOhp3npG/gA7RxjWygGrDnN8Q828O
SxMcQCiLDPvwksU5+5D7cJ6P2WfHL52pcxs4qsywGegQnaC7Srsp3IQxxVOKGGNQ
ur7MLLEyOb1n1zfc/JDoIKvtfu8NCTXW41yRlJAWv/WGWA+FNzRkcZ+EwNH/bx9k
aCTOT3jOmja4B5DJDzQlRqCSDWlgcrhwhlNvKQWGjKxkh1ITUH+sXoISL+5VY7mA
v9bu70w9qdqhINaOY/BW4JEp5iohCCmFXXHyxMv4VLQBytQnbZVBZpPnEe99X9eQ
mXd0IVAK4ukD5fa2h+4q0ciQMXI5g/TwxDIyL7Rh6A+t8EbCvWKhYg4DIoskgvow
k6nPzvLIDsLoeAWHVu5tNCM+D5w0U+AlGo/XOq7Wulnbwl30/jaYy7uYBrVMcgRj
r9Eau5HEkIWz6iSyZbS0peYF4XjjwVImYC/qaG/HduOZKEGYLjnZ5sJCI/P7IGSE
WYEvfoNG2jD6Mo0STcaVQjhsAGt442DBkoGyjIUl4halmPFig+Q+Ow0NgvNSeUGm
IiO7DcUJntcYTeAVGXfSO4+T5qzDdG/cgyChwQT6CrdN2JjUMnC8YZfmle9PF3fN
KNqxWg11ReIBl2HdLq4POjT9M/vDRgF3sGxQvOSE2WS8AEiVoL4gNGZz7yqCK/d4
1m5braWD6Ytloxqv3ftsDTQDMdWJXMLEpD/Tz8Ki1rHwxMEqPKEo+qQ1Jljn1bTp
eKJ/iGKHoH3NQIFasBDQMIgzWhcRwXc2ua43q3sFdbOEvE9cYVKpWef1qTpVkE1F
tLbM5TY6AAtMnjzVEC98TuOZ9ewB0tUTw/Rz+eesnLetSMzK7KdxiDXZl4yOMN6x
nlFOO6ulTuK2yYSwRiLlljsQFpboEROeVtcIOXsLVDBbJUDJw8I855BCpEeTFO8f
vLUyiGmBAMgw1TOYTiON4iXm0uBCDIM0HNIofHObnEhvoOXGXnLNjCUBeyxWfLw+
Sov6TMCPYAVeHkDq3YTSwuda+HEUJAxO8zYk9OYA3I5QZqDpQc9s95qFLJYtFD//
i9XjfYxsj+bun1Pa+WlerlW17cSxf4RxD0BWlOyZIGZrWVfgq4CvqRZnt48iXPVw
3Fh7PM/Ps0QJ4Cip/bSSd8gYrONrcbRzSwHFNfPzWz0ZXCj+Yz6C5uSHrmXeS5QV
EFdN8Zl1UOH2nWPUxLxsEbZFV0xAlgWdUP26tq7xwP1GYO5oXgiUXzXq4wF4jJ2Q
KiQoXephQMGzGXTLFb23Znc+2y68TCUnzv8n9tU1vGia4YGQ2upNIgA88B0UfBZN
vkhaWE/6mHT/76A14FAL4g55py231isldYvbahxXSSP6C8TDfV261ikUQXqj2vnA
LlX35v4zNpX/coa0L0li1WMyDFTQBTd7VgHFDSs9jEgYxEzyUq+9BMB7IjL2Q/DK
uNJbrhJ64ZT3GiWKis54+L8wtoGp0GvERvu2tINP8AUbHWL4jJsO9DKmXNKKwmEM
VcfVPxnmm0TMXRrJKEY68oE68LCE6N/g4yvRHvFpPsfJfdLpZAASrKypLA7bY6tS
v6mjgvZyFrizt8U0X2lTOG8zV7yJUInYXR91mLRc6ADXvnPnkEAKGc93DEEw90tR
0dCf6jUeUPWhCxgU0U+ro+1UHNDYWabGCePcDPEnI9K9TGahLEzeZMtHaYM9fNxI
Fk1n6asTevwe9CcYfD9jBgUozp4t7UO5X/atsOrkBUk+yZUampr/xK2zl8qTMizq
LZ+SxgWGsHC+LT1ZgRATCMeOfmtnZ04VdWbZ1ZAZhhvPo3HYzEUHP6f4m1ecnQ0S
pMwrvNjTHaVh6h4c3z54uzmstd4INL53qkuHxPpKS/8vMnt8/pYBuP9kKugK4+da
c753MV4ee2u296at6GNQCrix8xFWj9XIdQqlObc4Q66nrpYHmbzxj0a4HHH+NPgb
XgUw7ZO7sZB0ATvCR5bbUSF6rJEo67oLuZhJ7ugqFOapGIIqg+NAqAAZWPQ9XQx1
M6KXbaYRvAUEsp7u8xTptKNGdCMd7uLALlowdicTxf6qP/yI9isPq+nawK/vNbHr
P2ky0jXmnk8YDvnAO7FzZ+CcOZfUxls3KknLcYD4OUQZ64N4ZDwMKpoH3jeHzSyx
wh1VwIpHaSdXRsGS8MwwA44JjLrkz+eQglFfCWNT/cUOa5fA8EI2Vp4ff8/gqaWO
GBJUozqKPiWSOpaEkNDxLSgMPDntJ4WFlsjc9WU1pgiu4xjQDKLTt1j6wrETqDUN
bfYSrqj9x9a59TVzFikrvj2O+W4l01q1ZYE3uOLv4ax2T+Yv6OQWeE9Uy5LvtyN7
KarhhvEoGE9KGKbqVTnkkBNLbFVd9PZW1J8nZBhdCjaXAnBP6ZWqUARtgPfa+nPQ
slOvaJ5tJ/yTrdqqFosTYY7UUzFte1XJFJzmpbBjJOK0KhvYB43X45gvx9l4yXQM
njGdSE4lF4yZyAQEASyLSCFZFYb5lwwo0as55gjl1MohNXTz0qyv42vxwtREbORZ
BWBQ1OOqOsJViM1Hfpfjn14nPfB8wg+7i5qgtFrgRIvRVR+tU7MFisE6XPSIwB4S
vv+vQk3ix+eMrbBxQ6cXWq3xnVn3c/eiCme1G1EZ3ZfGzE9a2WsnO3i1xcEokX5k
E5zIsz+CrlqjnsTCSXbfTrwkccnxaQlUeWtEFrQVLGTbfIgjmvzx7X4xOUoWd4kx
DgHZ5pgsKWxqZUFt9gX7KdKEo0NS1oy64JdgIZ8vlrKjkfFwzp7bUJ5Y89NE0OWx
51LOfuHYSMfuxIQ8J0aMTdgNGIsnPDX2nTUK8Sb7jltA6kd9WYOoo7orP78vUUki
q3z8rXVMYpbX6IjBTeE1thJBwIecP8zC1iI7JcsQOHlzN3WcFSjyAHpXH67HV18S
N6QIPya9gLYaKkV53JFZOjsF7tbJyVxBwBb75jtaJdP6GhI5sWb7E+Cb5s11VCa9
hAFNkbqbItuUd+kMihfBVmI9JKvVyn/BW0yc6q634F27SfFdHi80n6z0VrbRMwEH
K8pLsbCkcZK5PYjp+4XHnD/t0u+nI6XpJVM2twobxPGWDaWYRjKIL7302S8uCF2U
x16DRxMvKQ3Pmd3c4SFl8Ix47C8/kvG5YnRBSXZgGki9iVpqdTs12WNJ4mwVKylx
9UdS0OZ615sWNh4fZuavw88xoAY4v4Yzj2QbrHGiXQ6NMCl3fw1maNS1o1g8WiDH
+uTplOoGgXx1JIrYLJKSrNLU156BSn9gs30lYahq+skqm9VTYxV/Hs2XR4hpxmSJ
cywYeAdgZFSyZS5PogBzzewu4oO95siOvV1DQu70cJHZ4L09isf5yj9Q0riI0FdT
mGYB3zHLMVuEa/357xI7+VWU93iv3V6Aw2PKnSMFm5Jc962RL6YVRLfTRNCmE5Gw
wFZ0BEhS3Mty3L2X+5nGMjmh7Sa8H4CoyEI5ehn1EIJcaqyHcewjSoYHLAs5vd18
8nsNwQ//njY2f+rjy2QeFopzsU1ELJ9b3zPcmAhuDADIPBTO0xLGVnAw8dz+hlpN
Gtcx0XqSxNtz/YWaJMUF8nKqQgNSX3y1F/ptyUFBZlRoIcHRcsC5MKT4QOdQGFs0
ZagvB6lkDn1C45Avdtaw55dV+myWEPK3cudgGwMeQlJoEBbGzgcwH/Whuyhia17f
F/gWua5e8lm9foOwSe1XlKSU1tDguTUpo7e+HVlkeRDslSTHfGSJesAWpMx7CMH9
Mcmmfimbhc1PIii5yl0zkB1q71152W18q9b2d6pYgLE0efbn7BT8LHVrlnjf60rY
NAcYST3Oamy1VoVJNsVF7LQ5Ak+OFuDotZxIQJ9olZjqmaSsIY57MvOLz6pX5Ktn
IxRoKP4OQmf7KpGMlq6ws6K6jD4Mxdls+9YuZGXvTht/fDkOTxgROJP9u5vpWCfI
4ZutNNZgxA0upBpU3UqL73t1z07tjpax7AwDXMVHrJy/KmXc+8qnZJIZx7DL1aBi
MVoLTwRpMLCGvSTxfkobJqEskDvY7RPSjgrwbIqAO2R8BPlFwUKDSkopel/AJQ/w
FWlo22t/DLbhxC2lkv8IZkQR3NfkflTNDBOCeJPFZqNOboebHbM+89GgZVQWe05s
t1qVeHGy/VIRtswffeMhu154mnSrgI0HRZynVKUumxG1M5gBfPVhMI/I41W040ya
NMZAsauhxhOoHDC6cy2vjfG3XRlyfy53pH3q++w4/4D95YvBWLSEZm2+91geA4rH
7plIe64TSxScm/2OzY1ki+WnpCMrrM7Kj9C1EOFUEhx6R++GdpVmFLqlEFbeFmno
RsA7ZBsxBB6GdzEbPyEuXkUzsZWmWze7NsBgUFOlPgSKOGzI0k1lr4fENHZK4585
iger54d1cgLyS6o0UYyzUIcF7+4RkUXuG0xN4WihA28dxTeJ13PGK0UAxIV+t/oq
VECP10h7zdqs7zo/YxkwEp3jiUZDIIE4i7hVSwwQxzkgdIcVj83clQ4WqiX+bOl+
YvfwCh6FyhOSxpTXqiQ7QTR89gyAPhmUfDiU3+EbMD5pveUG7BSeAjQPXzrsSG64
dXFY+wmo3iLBFl491zsuQ/6Yh/E9WBYtoNyrmsMgE9niFCfL+/mIvr6yri+6vFT+
BGRDjvbQGCR/z7LySefLQRk5JCwsOIaEEcrByxyuaImDI6Jfke8cT1oE5JFvfOgV
FfDrSGNbekgdAcU/rPHmoiq33xIQ3i+mDUfgCXZ/UZONXwubpKANu7ey6+o0mQcE
13Zn9NpGYVDoOCuU2wUVejlwEytPn/qWJT91nMt+hC85yzygNMkCvgcurN9gBH7u
2Sp/opSL+uGFJ4uJE73ASY06NMcCWyJNyLj9bX2hgbDt9jlHmhuOrWVr/bwOQ6ML
Cl42dJp8Rf5InEkemcQmT6eg+XtFnQ0Ub/0YctGvbp0CSC29++xlG6slXqxMkycP
Bvibu3ab4BMXOgK81CxJwuECuCF5tqAXGEDVHBaFRO/0weyyumK88hQxrsGIuhTd
LDV8SfRfhiuGwxStzOqTXCRBlR3lLSvt9cmyUcImyP4vj4Ewf+Eqa1gEnN8JOasu
eby2AMVNiZx+YEk7E94OKhX/vNZh5m/rfLTPKEvQymF0keimdvyMnDjlxvqcFxo9
S/YoAmZWuXcDUbYdy2G3PJqtYUPGeKy7azrnj6kVEk6m1i1+KjrEf8bkhWLgDE7d
kRQ3DyCyRlZoq2513DZSXZvGyZxlazq2i3Nmpc3VSquOHVUwn7yKWxtxn3/wv4Lh
va+dZVhQtGsksoDm3CbWagV39sqP6jaSbLo+KpgDAavWVRkNcphwTAejObVCFyfs
CE0nvo0ROgAjsjaFLKMkzqtDMEpm1jpAAg5XqMK+F/CvAqARpaaA4ZOv3ReuD7Es
Y5vg2bgfU5ofI7c7QlKuKxl4Lmv9aVUE7TpwfcjyHjD+q7Zg5niMmISK/aipPmV0
5aA1eeXllD7VKCF4r2rqQuUhPaaC57FEeTnS3Ry1RlE8ph6weSd1yaYlJn2TBKRG
HXa5PQqS1CkhNUigWodH6POIgdYPLbNH1QOb2rt8c7lDsPEw+H+zcjPVofEkIJtd
ytLmq05vaDPvhCvbc/7BQtDW3LTGSMmpqCkEVGqmpjuAVQ3nZFw7j8IFi/Z/Reus
S+SnAYoIjMy+4iJjjf6nB6zQw7SzpxBO/zkoYQalD4MImGeSYdaBzFKWgIDzBeHl
X53wobJ9hIqEa5hNVI0NiaklscyUcEke9jYRLieQtyBmS+C038+iww3cgtHQPt1U
WEQDyM32qwTMEb8SaIWrYDnw9dVaIiA5i9YzMzQqe59GOeEhLwgcLldjtm0gPYPj
j8K1z/aZn0OpBYAwRGaMN3HVxTf9lslMS9loQv6bamAxJ7DFzmhDd16q7mBfCMO4
rPl3Y2zsLAEeyxRIdnc1fLg+8p09kuxa9dp1W2lGKN14HtWzaUReBK1dAFRq7M4r
VxKfgwlbpHaYPL6XBabREEU45/b8NxKrrrPxf4eYuwTQGgtThxcQJvufUiVacI6A
XT9lq7ZwBGP3FBiqO2BKOdmyCNFuphITW2vylM4S4t5hVDgAKqTQwNdcB9j2hjQc
82lOZm3CGoS+I6c3aRtxJDi0HMwGzAScr6An0w1UIjSUwkpiURKWd3voc1wsY4XU
gzdvsYWvgMJ7DcfNA2DI9718/Nhs+OfXAB5HAE1I+hrF69Sgttoy704VwqatouVR
GV0aKPhudZFaZYSz7D3VNakDjdY8SsOiTh2ZE9CyblmWplhH3aPjRGGR+y+hhR5N
pTQ45OT0Zq4RfSVC5Fu6JVsjdoAux1K0WYEztmVG9FVqwPRaayjOscOLJwYp4Jwm
eO1fHhYf2y6iwn/+u5LOVrPrJGKQV3GvvEqNWKZ1FClMzhb9I+6CL9ljwQU30TPa
/anHtSSQPuUypvozQNy9VlD3WEjZYFAEGOKAdhe5qK0aVnxwbY8Xm0kXrMEUrn/6
T4hWTIPWaC+Z6vgmA99ig/15ROLYsP+mG70LV9scIUy7ORHmbgwtdceilegrL999
puhtFdo5TlfmacgyWZS7Cl400TeNmKs2RA6ifq+8q/m2zkLIxgGQOWb3vWmcuU40
S8ol9q6fmnVSbUxVHjVtIvjeJr2WPemwlVAvkOrsAbN3KP5ZYMdiTfiYvlfbJaj9
NQqZrocgaRuWHZT2Ft32xHvgYEQRPJYY03xTpn5EzFBiMU/wEJBBDPvWqBBAWwkq
Lh4hLLogYf1Yw7v//evTM4NMsX1iltwTCqDL6XwCQ/Xl+9GHVx6TaOY9tnJ5TBVs
0XonLTWJvIywswlTOwvlDznU3dUHZV2O/eFsL4blHGvdS3bIgmTWtjgIQxre1i7n
DMG7Aku26bgT8dqthj7l2kk8a/OXAnetnqrUaJLYEOPdaeeOveI3QcRAH1FFnc4P
hRVq1PSE2cGnhgAyzKKMXMmbObThqfc4nriTHwzf0mz2P7WkJsS6l3blNqn8o6uF
tGxEli3KSaTqkVAK0bd03PFV/4NRVgl1Ii42Bpmz8lLLEKEhdpRPjYhKOWlArt6y
cUqwMxyvMVuCdrxVGQrH1cg+q9I1mFCgR28aX0egjvK8ib79HdpBicY16mHppYgy
xAMH5WqwcguK5gdDII70klS4jpVVv6N72pbSBzsh6/EnNv1rR1hZS5Ct3q+1UND8
oYIaXAJOUgy1Davfd899lMaPbG1pqv3W5niWUhXmee725xUcyj5n3WJwblAhdJGy
94r9WjDq98QriNqtTjKHEtg+fW6/BHHP6nOCLRIpqMHdWqhh+BqwX462K4eqrXJH
+25kiiE+YV+WR1rCtpovqiNFKY7FKxqk80Sx6jkcVtEAunMAhvijV3cZe84j/oM7
KZI80xTlG5cjL731bH1YFuMjJuKRiJzkmjCgv4vzIz8aGrlhLgZP/Bu1ibs1es51
fGyQnlxTY8ew6iC5e9JExbAgykW27i5MrMGCZgzTo3Zfe4tyVX/XP//lU8Tr/h/z
8TknzaIpFqa2khSacyzQ/b3196TpTiJ0EI4oUq9bPYTXYMLW+VBSrrvXdxCR4Ql7
Lg3iRlvseP1KNEF+MjydKdFF6GB9npC3/nwsNoasjn5as2d3u8xh/geLWfN3Mq/P
pcxuOgN47Sa/B149bV1sTkTCr7LtdV6XBCwtqVJB7etjmTVF8iu/IbHPXSwK0e0Z
HiVak48TPm8vNMF4dLLYnS+pX4OGMtH8SEF1OFlyASJDUS2vJQBXRI4ywwhWUBK2
T9Zdwp+paAkpLBxREDAlFT0W//v/RjwCnLEJWjFLUxabfwZDZT/AOGbrpeK+ANZH
2y3cjDxwa5+VgJHHhSpLic13LayIxl1bt0ibsVboP6nzrhrXcvUJPxgzYXhx/c+o
/O5DW5xmmNJEAdsfTL67akjAeN34J+oSdv1NHaWiL04onPTI2FIzMH5yr7l5tQy8
YJ3cqSB8dBMU++p412Fc5QAfmKQb0SMx44lubv2+UWDaAift8TK0pkOSEgRQ0om/
6F7CYLvvMLZpf6Ca073ppj2yZEmoUr3LPJUDMk67j/o3p4yBflg95zSMn/jkf/F0
wAv1+kMRbbXqtRapieXkTNKcgUgkf7Rlx7Yg/STNTJT3cDbDiVgmSGbSjrKX9P/V
QICTsQPwbtxvpPxLhTdWzDFd/zH+FXztVumblXYMoVAEmaZDF3W+1sGD5qKUbok9
EDLti+leRlzdrs3WO6ql+zgU3dc6QPZJJdOvPl7q+bGZa6GYa85iaD4wVBFcY3w9
fko2N3E3KN8tUphnFSGBK27SD5CdTEwyk3Unm7k0+z4nLZopUqd/SHY8pLg2AaN1
OAwqGRBNFx6oMOWjY45RdxsjsiDwtQMysQy/Yf+2a7TiFFfcrkQi3h/lehMtTqWl
PbRSrLywaKPJbIQhOIGdpVHBNNkHu5oKGUiZk2hXj/xiWFe4w/Y27V0l8sdemr2J
zqu8bt5ymrP2+aHqr8K2kxICrVC8F3NMmn+XykpYt8bI646Xuf+A6f37ikdLx4Sf
HpCFEbIyT0i1aAzq2mnPhyAeS79U3ZmtLdzY9mfobrx+vggghY5eFR3+ZYtDzgJ8
aDvs/2eCqU7ZGCdSFDKQwIAbHG+4FkaMPpxJmgRFdZXKKBs5v2e4KoaayGBT7qfR
6X0miIpBTkmqA80o30E9mPN21BiBEu/5xgMY+0XmGfsHlvLMXp+lwBrvy3AiTIoI
PaFIh5sFlhq61RkaRlNMFGt7G4Uv7zlS3L9pxB6Au0VSnKHpZ0mcqmGFFPeZ9Zoj
2vHJQCp3esSxsWOe9mHukCu+EMKIfz3DzLc1MaS1o1kuHihotfOCPcy8WQHV8RAD
KqJfmuiH03fX+TIOtLF2DE+APEtprNxKmZv9divDtJidyx166ENYZVVDMqEtsu+m
UmxmEYIIea3Ce38GcvdzHYyuA+e2OyN2GFdDeJRVxutcyY+ghpwh7DjG1ECP8M2+
hbGpY25HBbNB63x+s5mOAZNSumV2sXp4mDYEmbZ5W7JRXwLn5f3BMGz/1EoSUDRE
zZDJzy3BDk8P6FpdbyrHTWbMBUAh//8qyLYgFiboqp4lvIVbFWY3/mg+qF41mR5P
dGlOG9kSLUm2q+WcMsHjBnPG7EXRvWVsh/dOcxtEcXx4Y4KExmHm/VyF3fcr5tFA
wlqZmLten4w7S5PEzMgQ9aZXUaIWAjrXXhz0fAXudMhVC0Yezas+44+TTUimCTP7
1dHN9VCUd1YTfoKFSWO69RliWStjYSzzVrZyNocuWS+sGTjrsQb/SqmWxHHFKRu2
tmsEjDIDeD6+0BXBbnr1W5WJKL9l+0qSBPXmwGSqZyyGuKBejKTiM1uzlviSkdKn
0giwdQikHw1G3blPp2mci1tt+axD6oclIUlIu/IRT7j4Ey9PCQexyUzlQLHAQYCY
/i+9QhmrNAkJM2Jf8kWQfDD8CNr33w/X+ukPVWlNiXgvy1uUL8H1lWGfkMgCmBs4
jM2kBQlfhcCnqUxNt1dxFBZNcBTyXW74BXm+ovfCwZWqxkCtFGJZYRw42VDGODE1
QMdcMKBup0RsyD4cTWsoRqnDGgWLMsSHL9XJ0l9SEu10zORkbCjYaaQewyLqfsvz
RoCGNBDZUHKuEcSrHrAdhkAcOsS8vSN6ZRaqHm/EPEDTFITn3+Q7S1xeYDz60xz2
4Ucf33n85gelzGfWmXT1pUnAtCixzJhcFWWPL/3QsUfkQhKSRyajUD2VCyg/9/Hp
ZZh+tgVoEXzUv+yx9n7IHoIGneZVrKFxCqQRoCsiP76X2UVgcwo9jZsrZNY1D/yZ
oYypNl9xGQBqKAV0Q/9kXdhujEhcjK8mQaMVZpmdNLJzMzOOQXZoO6pJD0Sbnrl8
jtHp0uGRkqqJv5W1Zv3wLqngD4vdrW8V9PxM55nka4PTMqoFeW4G9FMZucHjM19t
kH1BrGfCR4WDx5dqqMXROS64ZH/OZ82JR/3ITFEfPoNzjH9qMrGlBZhsv0C8sKg1
8N1oZSw8PC0w6C6BFP+Ol68KTTs+rpSMm2IZ69OoEJefXxCmGbXvrzdfhYXjVfr5
Cva4qRpac/B2As0imGnGeWQHIRzOhbGXvKTa1Vbjrr/CGL92PwS28V8DHZacq1nF
dQiuC3ztlwX7G4gC1csQAjU4fLYcCJx37RbEb4nULiLQ7Z3GQA9dNNB4YJvVS16O
GpuhpZj14gAnmarr/91e+ojUAM2063Q2AymLVJd4vlOKbPS6dGZn0X4+clwTe2rS
z3/3X7+ZO3iBcgJR/RrEyqzit1UxDw5BKDVBRcsR4JCGS81wWbx+ZnBORWNnAwi5
lQyl/QUJpNxYwGxo4ncPaTddvn4RRHrpwrrJB82MnteNzkc/grZjRZBud65OGf6q
mf7SG+/9qk6/2os49IuEc+mIxwTc3kQVT3SKdZ147/W0oqs7MSHcZ8LxL5Bp1be8
72I1zGg3ax8jWbffoes+YC2MeL1AQTD0Y1GjkDrO2sbJvLfMDGA2xB2ozwbQR7QL
rkR6krU/2/9ItDQehg7DW/qF/1hlmTeS3TWWS0X5x2ywJ74KtZisnBBEZd+2v4Qu
a8zl87Kn2VwMAQJ/n7M3gpeu3yh1lQuiAf8z+Ol4aOskt0tgRCU/3Ng+sWVDf7e5
rRo36T9KGZ8v4iSDeyauAWXHlRhTX9t2vRplVLzd5Bn4qfXelShoS30rVx3WVJol
w0aPhjG0XzkRC+/Gx4UQC5aWl8JJ7Em3bu+rem1UDWPji//U7I0U25MB3QDxYMYM
OwQe1qqyc+iQLwNbe2GZXEKIOFPIJB7f48Sofm4e5Iu6dUFZn5e8hTZ2OOvBy12e
zyuqsvBQDlPzF5UqWnC75oDpU10o44SQjWO4BIPx2B6+JMqvOBezVaT23VW/Ks2Y
0f0yRtXUZ0wzvjE/cLvwydn8+WDgqVk7UBCjOHjcUBaDE7PkhZ3ja3r7mMcnkpze
RSwSIsn7JHtZEQrIjVFcDa0GwX2Msg3NV7Rs8hYBCESa63+7da3c3xpv3bBpMxON
//OxeetIHB35UeiJTqWkyZCTwJaD2dSLEffvM3GiwltB0xKsJt0xHFRvRak6vP08
W3Vw9udHF5K5z9u+kpkl1rzJEf0cOLsu2tgD6CfC8EWMrb8r4RKZwl6BG2gfUAuz
NFP+BIvthLccV0g7O8qEy53SgqXW7Ki+AXrfOZFYNBFGsBVCWMc931vssTAvjqdP
bjk+jIASaWWmtJgTfnwU9bY5k0jVTS1TaSaar3B2XfYOkTAg3Ndpe0l79cFBqyWR
I6yvqX4jwDpv/VuJY2zW0j00EDaK3RPr2sASE82lQrr1xX0gu2+LabDlnAGO8Hba
iJ9KuCZWpLFHETFxYy6FGHnJtB21DQSpB9zJLuv1fGMe/pTkabZ3TPe+Q4Ibk7Bb
4o0boHWfx2LIyit4Wg81RlZbrRlU99xwOGgdQXslyWk7mcyEy3utzkWU5G6+yFIt
09If4f+WKFJZJRXPUO/9WKqh0utBhszrSIhMwxjVWe8Mpjl1sJYF8fpTdAG3WW3Z
qXr3fxDcbNLz07bKEP+1fqqLR6GZflP1PFwmxgSr+mqOpCmAU3OyC3LREOj0mPjl
d6xQkHdsKF9JiEGNZ5L/iNWUXQgR3fZQOMd8S1O4Do4++QuAyPeMYXQt+zzGiyMZ
p4zQWelwTVbIS2gF8m0JEdtlpZQFjb4l/0p+PPyWjRz7o7SchixAfE+5pbFS7Vpy
qyTU4keUGX3bnGSZi8gcL3axuJtyPLezLmqQGK+nxgXMRot0z+Rs6VaXvZwNwk/n
62RWxOLDVUp8nA+xcX4SoardRWUaVrGsT4gT7FraH3nV5OeCkQAGJcDBzG4VyADq
+gb6BAp35MVQ9XwVtEj+U0QLjV+XwScJQxmwshMHCfyUIKzJkS4gLdVF7o1jNixt
Km564mtG+6lGBi6qbQcH+eIugtcmmZs1vv4bIchcGTMYs8Vc6rZYtmQl3glGgMRD
AOIy7ipmIt+MuMZ/AM2gvhUjGVAT3nTr7FMytnO5GYBzJblXIDODfzfUpiPW+1Rl
dZgqNkU5CneKOwhrUT5+R3gdvGauSEPQAJ7Ip74+AFBXj3ey3tRriliQGyK40ERT
aAW8BzXVZeUEV0TWnLiWdutXjag7RJV9LtVteFSaIatD5ZZzR1MCadFmffl4HXl0
anwqzusLn8Ap0PG+fk5BqWTQezI4yKUwhmDN6ff0QKs4aNghF13zKW6xBoUesVIv
rFsEgJ104Zp3cOEl0X1OifUi+K0mIMz3AfdL+C2ZrfZUu+n+NapmXxn6TvFI44Ux
PWNOG0hmMFAUUS5hyHSbK3wl1OXOaduOQR1jWkW8Xx5b6w546KQ9jpU7kigo+r/g
ryN7UIfRvszxTOkda9IO5Hn8BR4zzlllgNNP2nXpFjqquYClv1FfvgdeIuHAWBdZ
mpfKXUSlDqKs4KdoFqXHd+9v4vHivG5rClCJKdNj2JBKOC7SysmNUi9gdQ0GN5dh
/REfPkkijn/KGikas/Qq+DZIzqm6l4UpvwmaXkik3G+2vBtOQYcaWgWcAiTSINxV
hVe41RkV1ZZAH4bh/9/mJdvWEcjYi6/gBLJilwXmQ2toO1Wx7EPI94y7C/yIAcKA
pb2wKaSyD88E6l9EShUtStdsSYe5Xss8kr/lc1+dM07i208ysAxlbIBuv9EkPFAx
jm7khzxn3veNOfXY8KJzDJiEvkulecBAF0aAglSNiI7tsfh3NooLD5xiSkX7COVX
eCnn8uakbtEmIdIsWYXshUjlaqBGS9RpbuSN/o7WiKp0t+l1YbnC96a3r8scRzMr
tcbG88VOYwH6N2CDaP+AH19Bu6WrLJUvb1123UmtYOVPRbFbCwV0gBDYxUFCfjo4
2EaWihpNGjnaiXldbSH9U8YxdBeffROVK2QgIfNKgOTUaJ8AvRaydFYCsIQerdwF
m+JCkfZ2BY1zt5r2f1BzSglL1yqnWhkHCqeZRCT4JY2gPEDaDe8M1W+hv2yFtF9g
1K0tA+HrjZBdbeGKB61LIdEGwC8EpyLaWU76niERQMNBc9awLzA3J1t+PpfHwQbD
nJYAaTNxWAgSgoPnBQ6t0KukEMQm5iYrdy6dBHqLP1dFsEBtxM18JczbMOAbkeJs
/VbYlN0RZR/DfP3zM3/okIXkrPzT9FqK4geEiEzfciYArXg9bzLwi56MBCD+57ZR
LL5pgVUCPb6rjBIA7z/1UZZRNA/mTLZgNTCP7IoZ4cWZx+GwbKMnzgikPIrlQLvm
Yi3NWcT1WGyUv7FMrm6FSBVCRuhWoVXVvcCxULmdVMSP+Iop5BjjWAt9FnmobAve
9r/6bnXSYVi0wEH3hg11t/eD59pYKeIPCBQKZpQdziknZ8rlH7H99bGUGBdNm9O/
GnWc/eKImc8jbfkZ/QzHYDzz0PXQRVev4TD0CwwwpzydizXvVQEm2TRjAurXfFhy
mjE63yB8fgnlOd4KGm6mMrAAUNQ2Rz7QE3c/2ek6QCSxDQ4GlE2EKr5iIIo1mKyi
u7XCPTpqiXIb50wM6u862YzEfbrUDpHAjN/4WYN1BdLEI/YjgrltrM3MOqT5v9IH
hzV8ddAjZaT3AjS0OvlN8guxwTvvAj0/n+KsKPgimpQWlbZxe7UcF9cw+HBxtrpp
VwZ0S9OlMMs+H1NGDhddhpiuEpQyrHOIfRjW1a9BDaj4ts4Y1+Fri0CK4Sks0adU
JepoUjNR/qvI7qUvO/hBICzeRIzj1rXfOYC57iks7SdD4/yjhC03jEzMsFCSZffr
3maWZubwt8iap9NZjMjfnMGNvOTpqJNFvIPFaGXQyBnhFOxU/0IDg9seOXNlpV3J
F5xnOWLr3vH9X6jN+S5v6YcsEdUN00QJrgvMpj8gUz5rwPdD3gFhsGMw76+jvGbH
GAn91AuqmOqR92F6arOWiV5EqMAy/4nITlTrsaEV/1XwqCa9JqRwpGu8v8AsTVGl
7Ir31DkkRGukdl3q/ofsjUohvqRHRU6aAiQhf9ifGUAqkx07i70uwMJ323pxDzc8
DJNRzHMPuZE4yl/TD/h8tX6kZq5EkAh/r13a9tIlZaxaptqIy5+z63OInk0kn3wY
FUyc6P1AsQgMcqKgMIdOlkLD5sM/YXIa18gKPfH3fhgIc48v2kc6T2JSbrqt5pd3
7gUU1O5nrkeDIbMJ5VPitJEUO/XE02OJ/BppufYF4vwJJp9GKry/u6/1yzb+y2wC
diejddWY3+jXYSJll3PcGy5U2tmHEMsVyQhZ3nKy95fMSE7j/nY5kAbt5Ow9E5Wr
o+jsuhq8I72jCkDza1ru8eztF9EBmTmQio1MyzBI2PV+MTmtFRmBr3affa7FizhM
aoS6BWZZCUdIozetC1921MZU9130LP/hfDDYcLJijq5FnJbZFQF+WEwBMYWmu91g
dCd47YGJxa4L47TJsqBd9QRVEErdQW099eg5cvPBEx5esT6U7L4REv4l1B1uZ2t7
9AboU2LNIVDi9Vi+eSWYSUe9RiKIfkCCAqzn142O1JfgafHxhVVecpispfg429Ah
mJAiKk/1Wx1WlfMjhX8QeGi01tryXGSxZk9CP282wqAad6rJg5U+5r6KudLckgUD
QDzDr8RSHE0IR3gVR1mSVEoIHZ8kNcDZprc9aFOAZ37IybKF9lbXKKQTpiIEoU6n
+uTDN/MqMY0rVvMpd/+tUcqRLJTYCbmnK2TzSuQ32ANqMMsjgH1YNGXNsLwQyIVK
c2Ak9Mgp6W/ZqdtOw63+nL6HiDuxcfuybIxn425jt3X0AsOJGsADQvtYwNs+BGBn
R+tEB0g8g6ROAW2+mFFSM9G8VM1TB5/EBsiia8DPwz47dvoMerOzS1Wlp841ymsn
nhKSAdQEooFZfCJoFiW9e2eCNS+7CIl9UjX0ubLowGNDKdX/pigjgLLDd/43SQDV
qkQfvJdT9STdD2KCnH7NJfMjgHhK0AF0pMwga4fobKXqEmDIyfMQPHhHlrF9z9p9
Peywqgs01wjPGdBQsYd7vO24rP4fefmU6mt/CRM5U2uuqLrdSHdF6qSpLCP87se+
AI1mhrxZbOBMUHVZzt2MF1RPhfljI3tLcWqYKWeZ0p9BX6WcgXT0y1y41f9+qnA2
mz6PvKhhIhjo4uIxyrrLu5IhiwZZIGdY1dpzno1X1MEMfm3KY+LI5wX1PKgMYUA7
3yo465TeQ8arNioTGod1CzKxARnsjlZU5zSpIBGfKQpKM/liHjewYoXQ7pnYMjje
W9olm0o8evAkLKaDQjceJR/uig8QZ8ruWmGmALIN7U9JZ9oNuPkXqUx/FHNHS6gE
f92KB3l0EWAlz//UhIlW5mLjkKvb/zgPeDNAv88+AOIwWcAWTkzBQL7aUQvSrLpl
goa4YklalkPyRfoWD1r/b3vTIr0RZ67sKGoWI075/MeF7mH4JYPvNaq5va7u2qMC
B1QvSA/aLRseLSnzfK8DhIPrKlHXjDxV/p5CXLclGE+AhXTYl6wH4csainelqmsX
aPiLUiVS9iwVcg5Zwmcr3COCwNINipZjmXqryKPC+xqjIMyElvImEEn9/X5Ff7Nw
ocNMTOIheOZiEK+06SHOwXoMJyMrmMBhJb1nm/UpzCD3ViwvyWtPQfiSZup2/vH8
iIxzzBF/Ad6XrTtWrAzpybdkJ21HgG2oxvMxhYyrIg7mRJzXkWU3ubpa9U6gQ855
DkviczYYSrD23DrIWJ7wshgrVMJAjx3I8RiecIy1Lagme+aSkhQpZIMco6rg83fo
gCfBOFLH4eevsNi1CX3D8ofPW5ZbQrt4CyVe4gYnYJKXs3iMtPTVJSUMzGe/SkZn
jP8188/clUbUTmYbia2mILnM91LrZRXiwBeJw+EyU8NZ49Ez+rHafgtW4AS/GNdr
1Rrya7svqxyPYOayHVSR3BElgrP6SP3II6m3wOg7oJqZGKnSQiMNWZZy4mqTa0AU
QQ5PU0pgBSu6Kju+gCrWhMObWJY8l/jguagNrwqxs1AG3tqPnKDuJSwdGYKYZKAB
3X+4zyqwCFYIRze6wZVJb/9K8GEf9UtgmHwvVaPcm5+c+ygHFncVhtKLH0cnfWE1
bdqaYulh6q+EjSP4NUFu1NsPlcq1jCv4VqDunmXlSnYRkZMX4ItENvxJbieqP+HO
jU/71MUStFuNk2g+W25TndgOh5qz6nVg5AqCt89+s5VfDGFwxuwZrQe4b6GNBucI
4lUCsTOKVQRZfrL++o8rhqjWN/ujcWzeNSKVTr/cg14sVyOGTn5WQI7IudnKNBCR
DocBTD9blVPcHB9MCTsJzJmg2rZe87V6utx5bDQ3gsqMUBfqX7DcAaYVCTZEAiqF
6C9wOOQ44afp160WteLUD2IW2hIdF+wQR27PGG68Q2bYVr2E7MRkRLfMeqE6RxI5
ylwVn2IJ2lbOPqFt6xXczo4LvBn1JzNWhNe0A9jFxfDcjQ8eS3YPBevi/XPaoMc9
p3OEqNh/IsQ68BqNQigZfIAdyi4WTIeEVNbJVdtN+iaaEffgGosiYGawtjNE5U4b
v1dnKxO7z1adGBy7o1CMrE7/WDdX2x6CUQCqDIIafRMcKp+hAPck/zF/hvs+KJTg
y7PQwv/HeuyZ1z5ozI2IBhdU2hIv0NVooZvJVT0QAmVStg61mGFx7AQ93TRFFl7q
2z6pmW+XHK/PV8QGb5TA/ec1VIHc+pF58igyFzCyjDYjhxk4SEXC9aakzf5mXb5D
b0G3qxhMN1DBIrFvT8zqR2PCfmS70Cfwzyel/As6WcWp42b1Rl6UPJb0uIqmZE+I
90DEHa0mb5iX1ldwHyWYZ5QQaqkGi88itA5sYYAI63CavIw4ejLaO32TN8dpbs73
ejdyXCZQ1BLmsKBAlholZ4IEhIFIqLldul7kDCwgU02B9XvhFFjeB+2Hj7Ptjzu3
lO7+5ZB8GgARlY8HdVoblK0g33Lr7wEsnFl5g6VTQAHvh1uwiSt3PPFCMl5BlHVu
DAdUaE5JH8s3qP3B5I62PTY61GHGsVHu4RAicLk3wLTE1V10atX59DUHdewLiHBr
yfHMxdrr7Fs7tdKS3xVyT0jNo8nTj6PdgnlW6Co288r+wZprcrHFdnNI1rrf0jh3
WYfxIj/DUKYpnXzTD00h99XDyFu7GhLV8aUGPLL7RCOKyS2x0ZmEs8TyJaJAON4I
lp80NX7UzBZZ6dkQGg5Almss7nfjOnrRRn58RqkTLBNDLaZLVBvofUsFYbGCQdpt
/AhviKxconiO+oIiK4xgS+rnnwN90lY1ph2e2tkd298yTR8hJ26ntOstpOpxv8wA
9dioyPHk1z1izxy5ySK6wMGgWawzEyOLFYIgAtzHdk0yse+4jO7MWpWRajpXyEXd
AOKmQ3qUddrdXABqRsBaHOYmKVmlNKJrVxlM+ZwuzCJdXpq46kkpGrzjAtMqgerX
rrSqtZSt6Oh7OOyXZJFgE8l4Wpx0C+hhoGniX7upGkMJDkspfSy1uiD1rzTfUv7n
y5jgBjNPkQ/N9jY3IaBsCF8fAMkIKj1d8PCB3nNhtQiG6/s/b4OwNFgeXmGs2gk6
fsccNSv0+xMVkfoMiaed22mvBWFVJg7r1nvlG6HU6lwyqDtrHfEXxzB0gGZwZmii
EzbPy9fS7P2FPUpLt/76ctfuq1brj2XL43Kg+so6PR8LE5B8F2tY/HlwYso5s1W4
sktknUYCLL78KQkywP/5JiospakcKRjPoU4qe4yce36Xbn/lOb+RSckhiwelFfSJ
j184Zk9yomKyVORzT+gzWwKBi2s1z+CLu2DUNJhd6NNU2mdk0+B+UncWbuNkJlZ5
eQOC2NtRXZ8fofQUWxowm+K6azTAKf6SFIlo51LizuXMtcoeQfwzi3sR3Ii+5GDn
LUtfPiVG3SE6UnpGG7Eb3I5IUQVi0BgpqYx3Jxoy1QWqTAQxgWXUUenoucxPY8sv
dlcSR5kV9mlnxoljeq4q/7uUVyy1W/qSCRcvDE+YVrHVXa0onrWGoEgknuplafgg
gZsJfjbc4B29PNdyS0sePM5l8fHOv0e795y3XzithTpmHs8oQZzg6BHHhFd9db66
3ZGta1FL6Ap5ZO1cx0PzD9s0Uv4TLT7z9KOb+2oDpayPKKJh4KT/iFigZ4WB0oZM
UNZbJlLvo942EzL7ouXoAiIbMVYoWiSmNC0DQt8qjSPiXz31GvMFzB7BFp0hkh6S
K3VfKNc/L3Af7LsmktWq1dJ/GCbWeYWe4NYr64tjdEeVq7PuZlH/qrS+Npk5LYMF
BkP+OB35+ey2bLKCWdQuQJrZPtKgkeOQIPpuLwtVLmqIN8fldUgvEm1f7MhD1qgB
r7K4H6CiaI3NGATp9IcMcCxnFSWGSRh5MPVGRa/E/VahJphw1NKPhS0CD0r6bP9R
FCZWW/HOPdZYL5M9rfyKzcb0EnjxPrmXJOPSabtwGkpoqlhNOaTTGUprNAyQsqlx
awXlWfVaIVwpyzVnnWYIZ3RwylCYsU7CcbzhR8nK2Ushmw5CKPE2iI7V9ivU9SJf
ZMYHRtNA614a9/t298MaB9At/bo791mWM1E/wV0B/1gRliuqRuQ2wB7hJ25itiWr
N7b4MAhCqiOe4XH7xm+PYLnOKkMXZuOHpLINAGQbJnagtDgpfWFaZsS29UaupoRC
G8frhDYGyxaggy6VbWZjTKO42KdYOZUjb/KJNdi3692LhC8Tj9weqalDMQDVMFMJ
4gMVUeokTkIPxiDCwENJJexFTjAyLYqyNPdPYSyVbu33zvnmgHcFmFmIdzZfDdpU
RZzlgW32hcGikfzBh2qPaW2OdEWu+Had0O0wmDJCKZw5MEnxFrsXK/gflJ9gCudF
Y2XO85Vnb3oTAUyoNW4LOQEtXAdr/j9YNyr9BaWABL6Ekcgq+7pQOotCsxk1xK5N
wCDbfGBasiru5Qwu4wia3/LudRa9IneTnJclwlHoKZRyIL9holLr0FLx+CmiWIQz
3W0/iGHh61oOjE27TL3nYaFPU3BWiHtMNCCfRUW7gp7QuKxOJ3bpTb34m6Mo4WOr
PY4EEoXl2eISysodGpvxz9teMC/xvbKiibMTiyraxsLbDUT/AA9n09lA/94F/Qkv
xHQMXRYuqGe5uDu56jfGWMQ8Egh3QcO0TqKYFLr8PPyIOr3bvifSP0DLTtCSA3YI
my4ROus3M5MgNM/nUZo83Mgc67GiwERtjtxlQj/tos9hNRFCwBp9GiOgtKylyz5G
B0lnw/zqMbRwK+166fmYgWdP5yxyZ/fYxe9I4eOV7aHmMz01VCCtRZwjeRhMBs/6
PJ5zDljxcdyxKMUMOKE1o65VxoEvcTbxdNf0u2qs5/hbPTQRB8T5nAq5Hg9ePhA+
yzye4Z2QOQ4QIJMVmtmqZaVHAZjbc7PyytOo234ilD2Nm0G9ibWRvH6Xxwe1S3pz
tIAF9mY7HF6znYihz+rn/P9uHKnO2Ng+PgzIfJVgDiAlCp0uqPPdXoOtLyXSUmvi
wpvw1SISvwO3vNperbUO1cNXyQ6MSjzCgQyWY1/T8+hH4+t2GUqRYumM8ctC2Ldp
mSXVGGfD1pCOinzprVaaKc+ayMZFvOtwGanR2hvbwNK0yr4ey5q+CjBLFWTps9Ba
CYlGPmvC50pbc2qSpGkrqdEAkjQEy/pFmmmm7jybyGobAg9PuPkdoaosRuC214vA
yf/Fwxz0ZdCU6GMYGxHf/SkmYQV1sY0bO1M4lzNlk4MzVcQ37ItHS+uoE55OoCcn
i0iP0p8+0kvZuE8FemOSJojJkbzpXRnV/liNGiTgix+klq4agTzZlVe7QyLtaRhj
BFABTeHdkiPEyATygfv+eLBIyO9ykofaC7pSADuALP5eZDQR0+6IIvPKEbE6V11F
o9Pp4LFIRyCTJo16x1dZIuOgtr+YDnQ21JNXsDaEcgva1zJhWxu0PsdIos19eqLZ
oEcEIYr8PsXapM9fo9BrhmnJ6nthkqe7aQh5QWU78xjLsTmqpImpeUgnmlPpjov+
WE9YO0j1B5FQJqap0ywhBrn3UHywcw9jnzamhkEKmO/+ZOwfLUtso7cNs6mDMoyv
y/AselzfXIVcOGr1Tp/E1r1/UvYGFdjhZtvESLwErxHTZBjgm1H/jrUut3g5xgiL
f5SLGqG2JRHGFV7pTW2/aiCKyMT+jSoJHgwKu+ueQLKstagQ8buKGyjhf/rkmTt6
qxtGlom8911F2qTkx9KX/HDNupTAd72XO0Y2haa01yHECP7JQoqQnkUptRdw+ObE
tUNg5lq+8MqQWh975wp4nw4KFn5m6waJdSRnWuekH4iM/dECQJZKTWTYrnbS9DRf
5MAdfHpVXGk+Ta4o6t4dc8tkOntU46AekxfmU0Qc/yAQzyYunlpoEUSGhCb/FqXR
0ayNHmkI048fBpkuAhovhTnzOvNLz6gbfNJ+3clzlzOi6amqkhW0ect3laDELBMY
cnrOT4ciSmdmry+dzT21Jc+PsQ4wWHEBztEXrXuc1ED8+S8GFLTfo8UIHhRgfxrO
arcX6pvTpfqV/8PbhKBNz/b9WW8aKoSROD33B5sEqnz8DwZBqEV2/nsthAUonbS3
0Zn3ginRTsoFGNI5cWtPi4Eq0tczJ7WFXtezjD9b9DAEumItDZhIiBPeVAwStmkS
1JgTLxzU3b7PlHmq99LeOp2tYcdSYCMnf60x+xo9FY5H5KQmx97QCG3qXBJUc0ee
Poid4j9uGE5e30yia+W2uhtiMzWV00QfzlXnonRTtBz12S8o1XnOgmerKL1yxsSC
7/jDfLDe9R4oEn/Db0Ss2iTCsA/2SO42Q/aeK1Xj0LqzDTIPG+rxYcBTSy/TVYUA
STuBGkXOYy3ND7jUJi7GBCLmj6FrZLmhKAHY6x47DyvKIK0duYXMdSA+jHKrXX5e
p1chjEA6XMn3uqOr+Q6mQKt36NsPs0ccqk7cvo4tGHxb2uXmcU338EbboC5bX8g2
O+KYTTXukikZ4rwOOSeEl4FLJ+8+6W2c98F5/O6ABNc/iiK/msYNKzDmCtot6+DQ
cha82CFjnT3OexphHe7ktu1hsCWHp4NDpTa+sBDg2m1q7+xav1XjXGkiB5wSuzTE
BV300rSMPabGQtaYvY2KHHMGy02u/20H+bhcgwfFQjU10RBnc+SlYb6tUSuQdo3R
I0cHWuSjNj+O3ju3/BXDv0NEYjTX4dHwLSEBy7spxPDQbBKfzpou2Us9fNJq3d5D
ap444qz2j+Gn2X53+iT1odOn2wvXa1X2LDoD0vnopu3YqfPKpSzPvh6FFis0lnYa
qrSxX8716XiC+Tf3gwmmgJ223NOtV0plvPwaN3tYJtDFtRp/iID4NJNl5ysg2Hwz
C+dQyVoMQnDwV1viA+dG7mnxdexe3Lg88m8Qla3rLQGxiQo9jhDfj7iN+1VMLhsB
JyLk58SlpJzbAWrOkn3RCn43iZRa/sl66HE/AIbRMUd4xQNmmqAuuWxX2D8GXcU0
IFZbOiPaYZUUQw6POzGbNF/HK/iNZ4spy49Tyj9CmqkxCn+SDz3Y1EtO/cLYVEyu
YMEUIiAqFyaiXdPMcL6TknFsq4JunycPOMwIYZbAfVAliyCcXj/SrUnopjiEBHpb
jR8bkzyzoZKYQ6+X6W7TtxideaheFonuQ/pdrCvh4d/OKfhTKDQ3SoU+q/8unQDh
E+KFZF3eBEJDUp9blzKOOT3lY6wxbI0m99fwP2vShsl460FNKm/eMFN124b0liAk
S/fNYN+M+YFSJ5742eCWb/aIlculpDozVOIPqrPhjiSlb7FvP7LcplWjWrdguyzh
zY2IImgnS7HgqhucSym5CJp+vKP5Av1BuntRmgSNuqJQm7Y/v5E6M+/t9aosJCis
ElBUgjSM00TPSbgSYN/P0r5EEIphAOGZnkBaNdY8D4bnf/liUnzdcvano1IVtZsY
5/yGSb4MI2eg+bODW/Jqsjelho0rkbm2ALSR8JyelwXzJQy2iQy7Kfgd8z7YsLwO
ONeAr2ivDkSALDll8NbKS1KmVrEWTUPQhKMt8N8TQmN63TWuvSN2eXnG7mNacn0M
B0BQAUK9FIzI4KyUCaqEvuHL4KcyI7TVqru/36ep1JYFDifY/ccsdXvF0oRooZF1
nnENtbZ2il99yCg9lZrAZsEoCDbORoqinNJEQh14z6s7rrL9Mdcewenvj/Ow7Ka5
jEU7ZvK541ErweI94n7dhoY7E3BxrL3bCgm3J8lxoaHsGsPp2C6aFPd9Z2LhE7fW
SXs5vRFHoaJjg3Jh1SV5yJrX8zzCLHo0OzfrKsDfSt89nkPK2Xu5u4yAJzdgx4GF
E5FYFAlTKmVBZmf2CFpvbjpj11RCOBdOlJTikaYAjIIluJJrkh0SVhBDeL0jwrUv
Q6fo5b0Q+l7y9hh26GEyFBlndfyTzadSHsOuzrmNO4IWDshH42Gm12wZ7SGeJsgM
mllw9fA7x0bg9crttNvoIETUI85QmIcOtZC5MKJxDT68qA3ISSMeLLYDzChlfFCd
PDiaH/1oY2LH3mj86FMSXtD5438/v6Yv4Ef3twJHfKm+FW+el8MRMWqQgp5+Twru
pTVPNia2YOBiqvMEYls7+kjDQxe2Kx2aKI+bkxv57BwseyRYaho8Kpc19I735iD5
vTp+v4OYdHpicyuEVHUui0+Z2opy6/N4cce8b1moGLhDf5BtxPCXlwtULc0tdmIa
8ayN3hwWI4sshQvdX5WaQA3diW6CNH+JREYzm6MuI+ICBVQcA80XYettHYXwZQ75
eWOJXLhH4SHdTw/Y1iRTtj5Q8BeSXPNkLag/tjagrDXgbP+QQrshTanLGblmRvsc
ZuAPG9/POIN4Mbphr5NCb6JYj+j6BG+W7FFktWTkI5srbIRKkNvEQTDaq9qBn1dn
DedVGqvZ3oKDVGdRTE6H6xg2WGsUkXR+beanLwy9ZW56lUe6bYmdHqXQqQ+iyTr8
ab5Ju9nfsJdqAGqYC9b2a/YoF85tVSluE3OpY5qCFUtnsZY2ltoiPYZXxJ5D3PI+
5qyi+rD24QIMi1agS5zPmbAroMIzKUXX5SwI6xBYEqx7giWNuxPeV+z+xnVIJNPC
j25Cv9U/SkOMiLV4NADdxaYY0TUG9pL3SXc57B/ZfrjgfIWFap5Pv8fwI1B05BBK
xF5t3nZ0kfRfNSzUAMY4jMZUSgx4KidKDbwqE1meGwPqXUhK47M1j2yjfAkRTTr7
xXMlbXeAK+6C6J2rzVaCck2y8R9bo8Oo+ljB3nv+L2LEGhNWf8WgzYs5yq/2tL6r
BjBovynxPhTB3vK6mCOVfjNf4KFWO7VR24G65kaIiPkRQcTFvmvtdtEGTwSeiuRc
KqAd2sKs/76YDdnqX9h0QLNko+M9YT5pTAmlWS61P2TwfC2mMxhP3wTCbWNEf29x
7s7+yYjA1Agm1nfkIu+QUGnb6StYnMlL/k4qyZpgUNSWPu+M1zEGubMXh0Kdr83p
IHA4VtWZ4Gm5Oh4qBxnPvotw1pZaDPH1qJEuJnUcLduL9ImtHn1dsmygFDpnDSuE
9wvUOfZHVs3cmz3L4KNT+Kjt3C8APmeQdk260lDcw1rK0Hud5ls/KfuplCGCOYuD
PCmMfIJU58DHttmxYe375iLz+hFHNEajRbCy7xlpcNCjq0gSlpvUmr0V9jTQTKY4
mb1E/w465WHV2YYyP/PuMvdwaRbYll4po6Q0RtfAOfOExEAQAARQ3S2HmeS7j9pI
/zcIV4hXVCiTlpQ6+ZRLzT7PRwKOeCzw7MZZH5sZkvxi6goH+HftOQE55DOzDnIu
h+phJP7LZk9PjeQ/oS6n1E2F1pn9jMaewzVxHZSeWYiBeJ+yiMuvd5R8qID5OmZ3
XYpTcdzukRUMyN2tyuRabm+RqKzfikzWvUelNYUJ06TD3Vj4G3Cq/mXarkQ0tFtt
k1kLhIZwSkoEo68RsVKZaHGWf7i/FWzEalHEWm6ZT/J5i3Hw7Q0m2Igdj+FXFzQS
RondY56dK1VJBwRfg5pkjneTGeip+yX7HLvPhZ+sx7wQygu9n+yMZydQEnTg6m3t
zNRf48Lph+wxfHf9qS0kBAiI5M7F19FSr6GIa0yWdXrgokThA7nkcuEmgjHqukc4
IXrvzKyITGfz0l4N6SAQIRy9ukNY5yzheksP5OThLOZG+pHc7vjlnW5qJyDsOpK9
drK/VqIv23DsiC/5hBsyxT+PraBXAJX8UYYvlqlLYjENLHmbusKhmAE1Mm9TUaYv
RN5SYzF/QgH/LAI6H4xfUG6YxhAVe8mVqGBNiu8hmrpKudnwmhc9mMOnXYRk3cP6
FBqo8N1XeIgpwgmvPPeg40NuBtE7lW4iYGvCNVOeVRcmu7E9Wgwob1e+mWNRgoVr
xZbxPb2XE3cVwT/4eLyB+G1ZR/OJZseAyQ1h/34hmQnNvAtyDuA/dsii/f81ivCO
EyA9YtCcD8bFmcm5cvOEjg0UkwIOYL8LsBYEnZZBr/8EHhkOKYVcNXAgRrK6GY4g
Y3JLxNesVaT5v5WK+HlKr6mmVlTLNomZ5IiP1ATPuqzV0cNkLw6/ccMJBOQnA58Y
6/AOBQnKMx49zp6BJJF4qtIUOWRJN3KfkM7vlaG8BWquMJcmB/l2m34NGiArfOLY
gqictDwhQszHdiE6WAKtoPJhZEZjEmKSL4SoF7WHVfDhFQxn1E9yF+8e9ed4U9Zd
ofSUMN8Zi8T/ZKpN6/5PiKmG5bGDqJL9oCX16O13Swh0VjhK9+eVgZq3G1X3/7pX
oxV23bNWN/17LSIK/NIaouhX3P4sTQ1TviRx8kmw8Jjpr96nbMAu7CXHPltf5Ypf
gzef8GwefJuTTqvsZas271SJaGK4ahdvru19TvzA3vpZgvd2t/Ond0tA2BjREFZg
WtDI/latnZA7H4nMjhCLuDww1guUpYKYfKQJJnmKSU4oNkcv5U8nIILa1NFNkY9L
ks2RTDUoJkjB+G5HKxw+aB4yTk+53IczidrxHZQjj6iWmKw7IWhFzP/LhnEAyxvV
fLAnJ262CkAqVyfi1DxT9Kjxla7pSqDUbT2FB/00TVN+W/7duwitOP/xu3NTGhjl
ZpLuY7VCMr1Qvj8ksBLMoUrRMw/GAqsmmQKeoOl1OToSC0yl9XblMCnK+EDZoqly
zBnDiIQEe4OHiSntw7qeuDKobfb+5sibhgQgbAvP69HEuFv1Cdh/dTTcRFaNeWZa
3vpo12e9zebefuVhzcmL5dq0lKB6pPE5rehT7LupCy3cK26kiORwImKGXPodVX4S
dlY0QRq3msXHjtEnTZh1Ce0pQYUGH5ScmVGW3ue0rGsF22bR9/98XTjyz7gRJc2h
Loxxo9c6tF7xZZpAEUo+ym1nikBzuofpPKrkJKQCpSvDkqSjw2FKUsllZfbnWeW6
aTrcLm2ULkHEwyz9JtCXqMCSk+/QVPSNq8PK8AAZ4lOC4np3GqX/068/KK+qEq8t
UvvaRgCf4YDnuF3gI4b+lzgIY1TPaMBisr+V6ctwwDu7VV9p6Cjy2cVssUGCWC3l
0Qkz1iVPikQHgK68yTcldQiMe+JKkJjoIiNJOPtyB432EDe0jZkWjdkQpZlVGipW
xzq+nplHzeMKSJTXPbLnsyI4t0WqA1csui/UDv/MfE+jped1i4AzOSmDa2CvL8Zc
IrI4pOvyHpNHIs3fOCIM4eBtOI18RHZWKZZjWRhLl7HrYI1GRjaxsR160nQ5y2aL
Mb5H1Wt3xe1G47FWEOs7fQ4XRDwieng9p052+b3m/h5YZgD0DbaSzhkGUTt3eM1+
Mt39uKQ2eyaBLPgyumbhAbMmDKWW1peC63Z0OYgqWQ49sB1gMrVjKRwbUc3vrj17
T8apaIxAK/21zFLoSKWEyAzg4kLsV90IU0eOF7l+vdGIYcbfqTvCEuiAcXB8gf1d
tFHxoMye6rSsOf+pQBM1/4rj/nE1ZOrs2rq1g4RdTiBQFG44H+lT3Z8vSmCzKC0y
IPIWZr2MkRIckC8Jr6ycq3YKcXKmr4MrOjhSRCaI2ObkVvOoRb+j5jVfLiU5ZIPP
eVY2jvGMsBm31A/7dR7HxUqoaMoLAX59rjxAfDJHFrQDyzCOvbZYlNLkeXc8sGcq
FXI2j1L/5E7e3SrI1hbq8adw7YutPFo2Lsm6B9h+QXX/RaC7VXssoumjFU+tPxls
jqEuLG+fdlvEWqs1d1m6+9DzIg/VBXvEiL8kaEV4iBaH7ZmFtQdnSlfHG/0WJ+wx
Aopb/yVRDEHpQ1OuNJ2Vj46jKoRSEUfUOZOyd37C3+/4jQvGGa+R0tEfzPOnncMp
0MnCsZX3FnCssBPKt0r0Xb1oUzexHLykWHcmVDnoLo3/LCMiK5i+nyJqGjpRjHkq
xDcTpeVcgA1VJqW0xo0Aap4YxcAY8HjNTVn6Fq+XMu+Qv7O61QmZjExg+TotF25/
WzHMpVmJKRJZBUxRGfdF7ukKuJfGNbT9IOX7ft3JmrohCEMrMoR2skkx03MHbGn6
jEQRwCnc3jrPLRSkQOpMtbgHznfYYbFWa4bCyop7N/vbyy3dGGT168ZVIo6PiCGY
QH3kVopjoVKZeQDAezmH60cdEZ2BqIKLWDM4DFy3tpLgQvzd2SkJEwdLxgyNLcRr
KS6nZwoxE/8+4xI8+l/BjZpPOAXfamFCt36KOdpIDb8araigrY/Frw0sDgyB5CmI
c3ZM7DD+MaBnN0IT9p1TYF1ovulwbEGrSJbFESmiilY2hPCMNwQWLZFPrpiFrBZZ
WHVbnJ/3wNKqMCDo3yUl7GchW9qpPRgFgoAaJBqXzA372L1kGfRCrT1+zxh3wDSW
VqPht7CFPUz9toZaGGVyTZNXtLsEsZ1Xc/xgB6oq8hsBfnpC7nm71ImwiMMmhRL/
capVt89vuxtrGNl8EM0eQSVCerOeVUWblNHYMYA9WmpzK4GO6z+7DiFZWiVAmptk
ZbJkoGoaFHGoPd46J6ZLQMW/aEOZ9xsl8KY/qKdkrCaHaqRlBFrc7lyQNo7ZCxtD
UrBWsF43d5/u1rcgnSGLwwLm+cauztCwOJSShfkP8KeNSn+8Fo8QjsfcyCDr4nLX
fGHbxU6KJjpKdciJXn/qNoyxlQgajKXqD1ypZ0ttbhLP3w5Y0YNoPAmhE3dZEDJI
Evbf4t5ol94HcXcTkQi9go+fh/YbVSFqCT+6ebGhg7uhXP7P6BtrtjPNrcsgf9Tz
VBZez86Uf3+ptJSXcTW2xFOiiIPovRL35yJ7HMCi7ODE5cX4XQdrd+a4Jj4C4NJ6
oGxn0l8QNOX3iLOcqhnbzCmoilBgWPAIhkR4sOnqJTGOIbRpdaJY5DViTuGWWPL0
Ls5LYId7BKivlP24fDPjKRu5j7z2xdfSN/QNcAJhZtiHQcU1MS4kFN9B7OO8N4Ou
0q7fvmQLkkOIAuVoPWBsDHJSnI9C7IN1//xvkqcZExQkDZquFGc66siQvZwDqa3+
Vh+a/h4FH2aJeH96rPYDOiSXpvrcWdlpqjkpAgOaZgmD17fZvwLGk+gm1CsopMuM
JO6RiPwiJYuKaamjY8HNkYLxymdZkWJSeW3J5M61KqfqxbSzhYp4o86HIFGh0AT/
PDH8OdSTEzJ7ebPkWDDjoDeUoq74anOrk2RMEHWqeMtFSc8L82FBrfwiofTChbTA
yO7L01+Hcoc8U2c+vGLcjjRmurfwJCUU05SPA2y0nmhX6/Pvu871OtDmrmseFV7l
5M0TL23a3U8L13bldqOERcGhjF9rvMYo9IvKrc9untoRL5jvvLxeXyD7lobd4GDa
VFVDWB6m+dp+9wZOyrebpGEaVleKvfY+NQyDgkb/wtuqVGfoDBLfcBv9uBwhlhme
aJWe9LjjYfWtduoJcduVXcMa6/FAsBnkzyrwRe1xL8TDbsLCYCBoSGHecNzeBKdU
r63j+RWGfOGmCQ7xwp2WwWk40/9r7F65U96E+z0eRydbWuJLX/X5+fb4PKQ2uMoj
fgo+rgWepiCJ0wP6KMsPIPbMnLpRmlcOhT3xdBK+59+RwQ+chzvqrZ7er2n2Xdg8
AE5uUcc10fagOHtOmd14rISpPwEaWwEJ1eZB4BeHXCf0WfXGE/QWNPLqXIUq+H3E
kV8hG1X0b+nB78F1j23qz6zPdr4Jaa6JwnV6jmBLWUkeNUcxsKNLiQqGPuEUUMch
UvVuYsFThKWDSmDfVfgMxSqzXmKv26N96fLUbwWxmlyHqMhaTl0MjzCu87HhC4lM
9DXeTQtrRS15yXOY+xq/IY2QKqT336zUg0ldWEhtp6wGVxAQ0qDxh+1Wvqgrm6c5
1QFHMjPNalstHXccoWUzekhdrbIC5CI6AxaUwhXzooUyE2Gbdf8QVA3iIexKoBr0
zYLpVKSJLIRmD3rVyJgDZVocn6gtIY4sm1ikHMP9GF/erDZLydnqLr6Td6fYQz8v
RrxwWc+2vwQmc4tYUCN1C/JjC/1ZIWnIs8Hj7eKxmiZavCWBHe9QZNFPra64w5nG
bLBqcpQLj32onM+gziWUf1N+Q848u2rZ28yluoYBgYLwpNK4PZxnpWTfG8H0D1Af
AA6UBxOhx/OW+dVSQ09cUg3G/w+6X+R0V6z55iRWCQmn3PZEPrJZrHjEKt4auAik
wmh0HJeGfnz61SkOAQZyjROdlJ9mhuACnG4Duhf4Vx/5XjzDfuI1D1CJ3DXa3LcP
vC7ovv9/E8Xd97UspOX+Zu3KB8QNXPHDFr7TIv5/J15+okwTgM582d5FrVwcN1w5
vQIO2smAqzb2I0Hyr8ugIjw4ui96BMjxR07n8D5+Z2Q40fLM7Z5numWTZ/niqVo9
aMO69otEJAIZCtzKDXbZxYS6pYcWDmW8eWs27w4vGn5E+CKxXxoQIcxDipY02zQ+
YBSGJF1SFDFl/Fx2boQWdsvC5ZOAjnbNUBwGbhyN1R5STzEWppK5mL76g3uumZt/
Sy/mYloxl8wn9ZIi2fmp64MbwOWG4/BCW4Kr+0eFetspC/S33RlTcT4XtweP+7cr
5ZCavwsgwB15nlOZeQAD2vvX0IdKmB26d0dNqXMig1X8IaomGzkhuBGrtn0Zlkjw
4v2dMrsg3rhhePxh/BbjWFJS1qptmURya/+Us+5And1aztMLjVV8BCsxrPEun+m8
pep5TM3RlkgmxIZOpONUwLIc9ZHpnITS7VVUctABs0YJqmU9dMnXpf9fg5irVnXE
tLwHXLyQuD3PBVn37Mm1M1ETJTeeKNq4QGjmhzU4ktkdxMDyse/GOgrAUiIXig2N
pcNRCm5K+JdSaoLeXV2YCIvDunb/rwt51wCKGd1tOpLQ/0DGCgjneNyrKJ8iK/6+
5W3HFA9IMpIFuKJsLspaMbwhk3BdTY1Q6nvFZnPQUkVjFR+shWcAJQ/JHrujX+F+
WSedbjmbyADRoAQsM2/EyNUrUPItOWmYl/FMOYoZkIouHX/D5l2hoDfN0LKXhqUH
jf1DXvTkG/1TJ66LbfsNjqYX7ltqELXLzN8nOHRuPXFHXje1CB3wBBuuUZdh1ea1
irOomvhZGmHWlIrjAr8Ssf7jGk45E3o2IZdL2LvNmzSFpUkhG+WMtHFAL/2cnYuQ
19nftQ1r0LCvAXfeBqh9a6y8fei1ZdKm/hY/FCiaM8hOIqqM7EgjvCIYMIJfCaSe
tGPO5JZN/NMELFMVsd8b/ETqoIa4YABAkClAsmvzBxTtKuLpv2dGAxFxQHxVUNI2
5tya2Q4J8S2iNXs4dohggMrY6HDKLfR/mpa2707Jvtgg76PK+rHbr6Qq4ctZ1/79
YKjRaj3hT8B4IHFEAl5IxNOHyvz3TUruPSYrbnL18XzXcykhK2jz4/993CiVyeyU
uk/+bUBamlKGJ8kVoIg5NM/6Uv5MoFhEj2HiDZaiFO0e/6VCJ0zlEYECXN+UHzf8
MXKlDjrwEHcnjVmViQjSb4vniToYzqjvFAZFxv9YSmYxPBE6pJawWgyPxxXfm7bw
6FYtTM5nCW7TpQTQsaHmQ0MM1NbyzEAT6liCvykd1dfvioM5mwJQD0QMisfYakW0
freqZXva+Wx5T7gcjwC1+AZPnT0o9FSEDdX7JjH4sHolXopq7/u4VjM1dhQ1CQxZ
gbNqRJWWxuSwMb9eFJQMR1x2n301bUlX4H3Jd+CgHpGSLR+j9B9sOAEXY0jgnxho
YpH9lHmLwTq20KrTU4VljclV54CaGMdDYHra/4sYO2M3s4GES41AjaxxpT+xM46m
tp/XvQFrxbcV8kVICb4nB74o29SUljjLQvggaKWyLDJEAv993bFV43mJ62Ja+Osh
34ioEJXJrUJckxNeDDQE0FRbzEw5z71RKRcZtlDJgaam/7JPMB2JNS9KzJb1PC67
7Bii55kKolJSKql6w/v5s4Cg1rnpEmU09MUDiQQsimOIpW/Iz6jvUMLixFpSPaS+
CvWDAJNTs609/wXeh2nu/yQLs6T3hGUl+nBYK78Pkt8I3c7hLusVQkUGALRtK6IJ
YAH3oKgY6HxCw3TmsQ/1TegwbgVFe82OIRfbhMsLGwr6N55zipmG1BmJLIyUrunI
4/Luin8z3xNJh/za2yGn3WBiyJBtnWVCgpW3MTyGKpntzqt07gMkPsdEEdYa8jW5
TUaV5psdGmej6/n2n63wj0xFdeiEzh5ZvjA9PEGj1MddHZeA+cxD+loM8xnpdY1+
8Xb7L1RfyLSl3URk02cmcK7sOT8kGU6J3aXWKAzV9HFFVerr22BLnfi1ANc7lVNd
9z1LQcQN6GIZLsDskU/gP4bxtiCYWOTuErj8ZR7sS9PtDfhQiFpLhuloFGi44/HW
lhuWSOGCe3LogEX1C89XSPP82SYQnbfFFaoh/xLD2aPNO3zUUdvDTtyidpDgaXcH
jDyHfENRSGbSjoQ5rt44hbOJD+AKdw5V+hYSHMb0vzJ3n4cWDZ331afxlEgfw2hP
fl7VQcJ7oMfPePc8I+oW/lnageDdjKce0no6v7LzfUcOQvSCNhsTYbaxw0Pad6uZ
1E0/rZLkhIjN6JRN2NyLWJ1bmdpVz19oPsU1Vc5GitY+MoJmKwjwGH1XoHIiKcis
ILG+qxQP+QMhCFaqRwrmxFPd8yDR44lQbu8ISM3wU9Tqspryz8e2jx1ePWjghC+O
/Nv/cBPbltctykbNMf5Kxmv+dcbkuDlyxQ2YNSBwl6PoKDy3WMni4xcD8Icl38fV
K0W82OLGyiViUkm3qDmY/7ZL1+EZ7et2IqUE2yV+dS9BjzmQkNVQv/1+AQWeEZdi
9vUjRnyyliLPKM1JRNb8ci2wnEHAFJIk0vlvNcsvXFjqhArvWsyaJzawG7iKlp4o
OSPpC3VfQ7o5DWReUXNHbDIfStIJEmfG7DKmNbkgkIbyCXnXFeeAwHECkArc7Um6
wByVdkxWJwGD6+mBtbyjNqvm2Wvz81cB0Kc2O9cW/A2RIesFMuYoSHHvlLPDtlIw
/9NbbAcXKKOZR9whllVmpYjocYSZsed7nSWtqBeybg4Rv80bXdiaR1QhG9/93tGp
3pcqqeUynzGQUA9JKINK3We1Bz98cLOqTSBFNe8FCXNaw7dLJPyHMWKI3tCDExtR
hOd2lKCy7PKRHvvPOxGoXrAzjLAR38Ql39NE1mUoqCaPcwaRgSlmCkfOoSOquB/D
Qhr7wABnwvRdJEpx+VAr82NZ/wAiksC5udYXW5y1GS8cpdPvmjx3zJmg/KRQtWWw
33QfTOR3QmE6QFOGOkqblI7UVmq745KkD5iM7IXucvc59TaoyjnW45KY7iPWpWkQ
REgWaKmYyJ9R2/wNl2bJ1+CZzDHqu8o0kqyzk0pbUTsuWR2S6XuwPw3E5LZCppIQ
urMkfA6xinOxJasQhZc0bjMQRrYur5QHmqJErJhmxdtF9CxMu0HkTk7n08AAohEr
EY2FAZ3itfNNvghzjR5hlP6G+0mvHDvqg6AauBHEYRmRD1gLzxpiwdjy6PGSiljT
uc11O+Joue4hdTM+IKjVsYZN35aNdxHuhBiz18BIkugegyBSAHxiOBWXG16CXvCw
lUnPU6J8q6REEyA0LPsFfTvKZ4bSOvgBaqD4ZPbDxM3zrkHKwy3JbkcmjnESiYCy
oOI1LotoJt4SyjK/7jkFO3BDz06HpJt1n3j9Uv/eT7cfoi+EkZiZmEPeOQsZm54O
tUMMjOPFs1PR8+eEeE4bCV9fLdp16rZjiNEdZ88w+4B9hsSxF6Q0YfjPnG+BXG2q
Yo4LHDcgaYtFuelAzqFl+u5fVcurlWwV5A0h2jEk2J5tDSWFVTv2qpMxOcLbnDh1
EHoztpHn32yAGL5K5hJFPBtJMyaFj4vV6cnjxQ9SV21tpvPEIcKyNZTM5RsH9kQk
ajmOwoKL93CvWHp3VTsg07wdiPQRbwMZtAqM0VYReQEifRMJqiHkL5pzE1EGk1Aj
6WkVfOXmm2IuLNTsnc5qWxVBed5GgUzktWmVQTP/WbAe+5Ltn+nMH9G3MUc1FBNZ
3dXjJD+EF3bwWHcGnClHxNH7yxtJJqvpsSxLtxt1auamsvn+imUyG83bwt3kPiiA
g7r61FVYa2DnZ3PhFkV7fENACRMM/fVdLYZo1PXbENFR6HWu4ZoskTjwC+QlAbpL
FnG8nVfm1dKwsgMtacTk3YWLrk3R9RUI1AAI48u7+FbzMMTG9KPmoeQq01+ChVLi
j1vn1TUqyWzwIdDBXSC4TfOJQlkvj+GaChDL22xmBuDPFLgitZCOm22EBe0nLZcQ
0RjhSnlXHm0kLiTkmfP7PZvRiribY7LiO010YFbpdXkA/fHNiYuaWnvPiEp2S1hp
gUtgevRyyr8JHAMfymTVeR72oM/oS5Maf5QyJQdKlmVqCLHc4y8bR3Ri5XBJTClO
oi/azu5vrYORx4QyIH6b9UZWXEKHlqmcCQOk04dtqkV3UjA/EBzGhPxs02ENPTdx
qLtT7TF3F9Gd6UiTK4rJBhTtWQ/w4Cy1uuuG4EXV7jLCZ7j4FRyfLunoS+TC0Fnu
gefH05a9QMBWcR+nxZI8I6hQr+d0iQ74zdP5uGXjvDXlxAKGLDdMTTg3hWLg4I4a
Wg4P49xuLiwC4Pzdt5CFAX/LlNIGCyALxCfZtQFPs/rVipz6KPEAAIuNLBs5iFwJ
EQrKx/Y4HoxLytppFV00IDKpEYCWn9ha74XTTVhOo3GjWFIOUuOE4Xt9dUzY1uiP
sSYlURk0j4r27MCv274dF5KhZT6nI3Lpwsbtxk4yoA9SEhm02sQ5FITIaTOqGd4C
9MZXaefFl8VBKdW5QW/7OCb31R+ypOohVB+o3zzv2UGAO9oNB82luCU+NX9xnxrr
11/MtB04RsHhdoWvfoU5lvIMfdlK1W49LNxStR6d56Z+eaIlkC+qhRIhDrSQ42V2
OeC10p7ReC8Zso7uMkOUhHbj86CSQME279lwWkpWJGgykIgqA81bHl5yEbPoi2V1
Ddli3KfJL6q9fLiSSXvHaT/Azjtw2Z4BDCy7cZZy+VmtVOOFInNqg0tGZclL1nAa
KpQ526Ii690D0ucn46AcgvImws8D97FaGgH5fU3Y0MdgyvOvIeTmpdY7/F2Gq+Br
jIT0jW7B5yokzHmSrVywpMZub0c1eU6OnZUAr5b0x393dA9ay62arpwr0nkUZxaj
VkB5zO6LmNgXtoWnDYmDCKPH7We5QGa/ISmA1UNPptl8IipZFCNmcZ1eMDpo/LkD
ftYVF8F0SAh9FV9nw2kDI4NLzd/U98+ABAQu/TvJ4LOc4HwoOZ3saQ0hZuuuTSKk
Q91viGiF4DwHmNwn2R9ZCOuAjYN4NFItHJg3FKnHx9egftPu+1YuGTmhydibh9wi
vW1ASfLOroIMliiTggT80gzt3O374VHwuCBzR5W8U/E/jQcdJXTgMQV5X4AEWF6C
VAqr0PLCUUcBTJvrwV96CFzmtvy2G6b5KFtJrsiHBI2vBP1rI2TEixn48eEzWrET
wLes29GRf0uj1Ho2qKGEejqtmFHRSGaqICNIFJ5zuTLd7BhG6E0ADkUn6OCsFj0y
zX2ZuESWLeLiUm3uPvJE7LaVoyF5cEHwJPJsCAZEAs78lalPRxn9cWQsfKNfi8uU
DOmWbAhQq9UPNZwQqJnu4g/0w0qdXFM5k1REgALomhqEzOYUOpRiKFaWMNRw/eN2
i3WA81ohDmgG5CxJ/oOjS/rVqwTwIxf6HbkS3H9aWtE4Gg2gMjh6yPnXy85wXD1G
4iGaaWKzokzUzoQNe6GtKwFsWAj696df84lLB0ceSq4torvMCmyibn4cdMnoaVMk
g0Sy405BpKywMHafAzGfYbtyZr38HRoW/IdPu+xoPEVug+ZqDhuN9/YjzHGNN43/
DTFF5nOMAUBaY13/iqnjpsC8ZHgAPf8NqSzZSb2jQ0LvPiMuMS9ylakR1Z2D9GpJ
5TXljEA7zAfud77ZBCwYUp9Qi8j9c8oIgagw8GMjrN/Ni2buRCq+w3mcI0hHq66l
S3Mh9zAUFgMBA05NLNRO1Y8K4IiwmHodWajxV68q8ZC+LuTSHQhUARlpKWUPPkiA
uYoVLSCdiNThZScjhvfWsXufP/qkLeivgUNGtmNUm7ROiPRQoMLEGBVGgzMyGVBo
oEp3QNGf0tu1JMPhaDxlfuwBp1TMLYuuG/FRzUDlqu3oh4kDkThn3wPmDLHyHrVI
jzIBUfY4ohiWGDGiqem52k4pqpP4yfywqvYx8EIqW6vhLTWu+UcVC5INSNpf9MRF
v0Juhul6jFkOgFwhVuIiL/N1IbUfG277jwnShWR4TlcC8rPYTCeQIRKp70bWaOZC
xKz26p1e8aaerzq+cUP64wZ7EDb78KwMs5Rh+GYjZXBtX7sXZ9Z/W19k3Sdpj8Mn
u8fodojpfI/8ZoczmzObWbsswAkEEVI231ZrbcGGst6jg1PH3uxnkRKjDAES5IE7
r5fPf8A2Dmeaank5my5VheHCvnIV0m3gQaMslUezcvHouXgm/NgKXx8se9qXrJrL
p4C5XqaSXnKbkkP/Jrlg8XyL0q3xIJzyLzBDswdOZTjygQqvkT0ob3SAC70XQq49
Y/cny/0z+fxDHM/YbN3OWTgGV47WWbFzVIVaq+r8rCeR7AEOj6nB1P+ypOFfaF8i
sY9DP8wGUu8eAs3a2yauRd8wpfj3+uBl08wSBWLWCuc0uSM1G/xlgrpiKhA5PDGK
Kd0lJaQr339C7ZoTWG1gcdoQEmPTXjOml0g/DUtjJM/H0zdlHXUFdgdgwd1hAqm3
3DvtYiGg9DKc30ey+tG4jJTuQI2ZPtmm0QD1nTa7A0wQPPMPLf3e+nurPSQ633O1
3a7Im57GThjkrTQXZSzZDxUsaQNkbgs+6ocCZwOpf43wbb1KOyVjc6CCRPBge68Z
LkTHjz24BNCQ31b0En2jXtbR1TtTIFPG2wzRHYXJ/uwX7rGA65G9izB3ou1h4F+p
/j/efPFBeZXW3pco+2lDnclzPwbwB5pR4nM1sR9S36HMpIjYBDc9QGwMtmEUbwU0
e0mxv+tIgTfrvAbOlXWcSCV/j1UzX/WCpM/fime+OOeBtVd6RPm80gAUpJuOYToN
hbN8B27wUMMeYX8J0kX4LOM2Cs6gbmXzIlWqI58qEoTWOmnHh2mezPlxs34/eu0i
Nonc1X5JKiKoYVTDotprhD2lB6nYsB7aF8qlzzVxPTwSDhJSgHO7I3Rg10hGWIy8
0jQoJ0ddvLTXaaqbfCCaxJCaVolVHS+Abz60oDR8sXXpk5NQozCGZm58xaF0pr5R
e951ZzlV2kp0cpgrsrbIwhV01/sC7LAIBpE8vquGC/9Xpr5GkgdpPpyNtNn0AHHR
rVPxzp/lVfilfFBIghqa3vbK1/rR5IWfMBJ4XGp2p2svybtBqMF6zjarxx8Alq0q
aeO04CTVlFPaq98x0vjC3y5nFmxzfUf7zHbluX8pb1u8norESS3n4aD+6ZwStSvK
gnvCzex+puYy0ughHrM1IB1u7xJYnUS1SCXVAMt3VTkdybe/vx5zH9NKZLeFmz8Y
Qw1sZ9Sxstf4GmJ73cIiBQZOkDCAvxHsz/M1gHFoXwkTrq/4KwyvOZc/chzPO5/b
IZJj/KUgaowIY0Z+Mr5hbHF8xy2psJrAYYmRkvwYFA2bE/tDpefdYm8JUt47Nj29
M+gUdoWiCz2HLVw8Ozb7dsFC4Z8FWpinLEo3IgIAwXFfT9vEnEEe8+6rcj80krg/
j/FSGmRtt7WJ0q5BxD8rFxBZE1LRNiCU4dXX2cGk9YJ23GPfGklH8IkQ1jyd+tlD
BRFiLhiVh0N1eAIuhf2+bjhbKTw7PwpwKguTqmhrMfPNHDUmvDc4pLZyO7bxcWf6
zPa01kduEvDStQMcrMBeKcJ/HAZ4Qlpo+hAkJteYMakPSooU0nvmzyxG+SQgsJOo
0BpaekVd0uBG8/nhAngQTusFbPdlMSwYFfIU7e+zeazs0i9z1gDQcscpmyYVJmdI
eA2WMSdvmO2UVEyHtAsA28WYva+PFUJGYD1peI7mM0T/EqbZT4Y8kZED21J7g7Cs
HQIYzqGiYvzCj/4Tgh7qsEBEHrmhefeYNiE+FQeWmH6bVvvN7tLy5jKWI4m5LbL4
msKmKZU13P8EmGrNWdfu8XjQnVAytpYqWYED+hujtFIA/QcR8FSxpxI4/f3UH0Cm
T6erVsCL+1Wdk1cxUDnm27hTAXmHDM5G/QePJIr5yodOnG/ekgTlUJC7++Zdaj9G
vNeHCLugRWROL11Vxe8bMltDr/xq9XxReLHEC5JgI+rDZak18gA9iXoUs+piE/gO
TQADgex6hVdQHbjzBJnTBulorLAzpOf44KB2rutVAogRXK5oQQUkXNvmsTqNlemm
YTd23msBgwn7vuc3V9q3dNhEMf22KcyLTrV3kmmTPY0f/q3zCUsv2NbpPBhH+uJT
5Z/d/DQ5d49JxxH0RiaYOpjiTw01PchvKxA/R+rZc8E/HbNEZpmZ/+zQ/GiYxLr8
qky5mWSAv7MybhkAViVGlwAMXHq2wnu/LbXpMaCKMJD5dDjcPzmX2GYQX43J4UCR
7eRWrrOmutZKPxRDIh2OrjEJUgmnjBr4qAG7FTcSF4jyui+iStTp8kIuzxU0CuV1
lUKnQRGQ/Ukw1o/+d8hHYR4VoHC5G/yTFY4vX31g2qVfglcMiObmhfKQ/ndVTOat
GRLII+SHI0K0DSnPxb02UmGL226S3k9g6wW+S0EvqkdKm2jQ/jnszct7v0wFCWgg
yz1jIpGQ/Qs8g72+WjR92aM0F6Xm/V17/Yq/UEVYuwLngYB4cTgOv8cNNNNXhtBM
NpWQJPtU02YSp4WmEhiRZC6uoG8u3Ek4VJuljncyPvZlU3N3o6g9kCh3TsfA1jNF
1AyQyuOOnWkuQKNOonVQRTAAbM1SmgTPGmZQgOh3l6Na5j4907QhGE9OREmVsu6c
vqUW5J/NCqTGXNo+z0JAn0SyQukeBCcV0vKkru7lshxUFX7mbV0phHA5EbSPLp/1
vxygsSShPUzz3RuFQxsvPxTT/QU4MloLlPR5Q3GBsyZZvmRVn6rwHvUCD1gwCwL5
dzECmDc8Vdrc8AFKbMb6YrLsvhxeeIiYnAWbno4w2iOMrk1BlDX1isCrIPuHvCMm
x+jYMRhwWpFqd98pFlEQ6Dv0xgWHSOxsSehI/4dUgsdMMLzw2UEuq6yTmEKmEkDw
3Z9HW+D9FOTsvvhhyhwW23PPa2T/2t2HlEc7Y3Wd171Ood+zcQJanhVZjUtq6iDG
HF+JijiDx/1iY+RugN4OWEERCnLnApBuTfbmMfENfIO1xQRj1oKRzCA1xonRbfGw
s20tUaFPwD65XzITE8fIY73mVnnBPmKr++ShUXPAbYKQiBjcvxRXNMUqRtU91XHI
j7Lk2b18vckha+rez4BLfBq5pcnmUhBiCu8AmiP7MgOsNXO7zb75ajyb6j7rVLs5
of2lBJoxdWLvgG994cXBLFpTSAu+4de1UOeyNsKsF+fQ+EHefFvhTncI95aPlCYs
kgUyLw7l6iap2+56AIUgORh8cVpN2caq9d8xOODZKteieTtOBpDo+StHJgkLOgSG
0TlV9OaVXapWPpGkqYAlL+coqk2bxWPx6QCYgg7fOpS0/T1Z0ZMzHBdZSEDP9XvX
6687k35jwcaSJ5P1ENfbC/6kF/+6/HLsRk32bIby4ub5rWMBwMpbZQtTFYCpFD7p
zO8jK8Zlw8kXZy3DkICq15KV5gFPok9nw3NUGRKcgNbfeqWi3Y6wxhq3ACQPn0jw
C/x+5u6almLAlgxTS6K0ilmIeSM1ptGSf6bv7WTZUtOnLatS/ParoI8qvXfc1pwT
ptKHgtMz8q+wj6IXWOfD/ebkTvDWsVh05L4wbpfhJyEDjLjOXwpJROWgcmkNv6/M
cRO4/SjxajMMwxhGJGlmhjDffwYza0IORcZ3XfeeS1NG9/ZPwVNlOUWxeIMik6u3
1aRJ5d/rzosulTXrddpvxoSdnnwsmZdgP//QZEirkhegwyCNpJVEGYtIjptoYPxv
9Nsg366ZKz5N9SyvT1YqceyitVPuqP4R4yi8y/GnXSQB93tFc5f1rNcoW3nyp2Hk
K+t/dOk8+9pYMBu6yG8tKI/aDjNMWDL5MHQxFCP3xY0AsVTBlVExTs3zjtMGbv4f
7d9vnb2x1xbsD37cSVa0vGWorbbhqcJpi1J3QRx0mbTxUXQrzFp1xDmEkvDlZkp9
YNME/Qcys60WdIHCMSDK9vum/vQfJn4E0aD17L/zs7BbmVbVEA7DCsdUCQZ7Wjgd
jRRbvJLSNC5afLmszULQr/dL2te3r9S3lq2wIpNriAeQQN7eJ4ubYrZ9rwGB3vTO
JNcXyVDEQakisf+eq93B/HR/xfmmsFlenu/S9OBxSre9MJecOmBNozu6BmoyNbid
ez8IwapKJ4ou7tS/hbiQLkKylxaw8FleLVgVwx+m3aAnMuVbxWrBL8cjbty9lw9k
DXLkFPJ1q05GrvNc4MCLGpxK3GjDjufWN6P3rQAolU58+Y4KKdttyN5m47NKHQri
ReLqbX4EZqSWC/2EYcn46kKcXWFmF7BOG9FpFvrCYuc5BsUrGMfvOO0fSaloFB2m
q91UFJVcxTPbmtjwJSe5YZxgkhOhXY5j8pggPh8XvAJbtkyB6Qxp0grOCNGJLjLg
OOiWk+GCaomLN0UwOXuthUwY50++k9jEPdcby7hXJdu83eSnfRDGCLQbQyeKVGDQ
j+6PPwugS7jL0PvVlbrr1eMikzbJk2P8hV8TEvj3d2YRuq/fxFQ7d0/+6tt4NnCa
QTJuAWPOVOIT5KfTN2ixU0TNn+S+0wx71HDfC0ZEgVMzfFAf/KB1T2Be48VLgKbb
1H5lktX6qXbfl4BRTuaYNxknz5w+Nm4oH9m2+rsFxqGKX3N30St5WvrmJelBicPN
1H/0RPiGI+3d9xykfu1LkZx6CrIaxbXC8g1r7za1AHPv7r+efCQstVdhBAOaO2bd
H3UJmMig4l3yFJNN2oc9SUXMz2AYv74ad7vMplxIsiFVOhvyrGiDdaejVS8Sof2D
VpYu6oXFDsKKZhkFPb/LmbvScSEHdyCQXUZDzD/WsJZDY/s2eetrRodbeYAgGJ99
TpZm4tgB1hmtC2LqLwj4R0yr0bdqwtVEuPoBsgQj1BkQ8bopbrwqe3X+E5UVJ+X/
0Sdv/sBJFW97UVfJ0G1z3vefBWxykQKsCgW+IGJZPn5A9VHQ/+bTrjbKUjQMA0NG
ni87ObEAJc2hCIEoiu5iYmNonXxbZJudd/wYSeQ9XvorItBayPO7SEA0DnbCFjNE
7bc6GAx6oaTtOO/f7dlHNHZP4i57bd1OJsDlvtg6KT5fzyuc4sZ+i2KSEWb0uIyj
nP0LE51FLcQGbtBDpZ4Di63tzmhIi+g81FzEz6nrqlePz3VGrBK/FfroI2WBYD1A
TxSrjjXlFfa4ifB2AK589/EP4QTgHffFWBkMlJM7J1eyFADOJdFekXAAYIJ5EEjg
dMZHk5byljAWbViQrI/x1TtS4IPS79FDsDCdYoa56c3xgfx/U4DGkk9cd4wW2X0J
owhc+GqlTaY9X97bbCZ3RDBD2yldqNyYJxUwoBYuWit/PDwFfShbO96xiQf5+VGe
nPgbccGPvMxrBSQEVHvd561wzVNFw1pUWAx2libqIqko6tD0sSXFcB3sS+mEd4kD
ZdvhFhkuyi4M+yw1MAhB2/9v3iVjh9Xh3358l3GKBWYES1jX+qQv4ahXZuxVseoF
WKCusIVofdPQVS4Kjrh4kUmS1/Xz+gqttbLlCrt74UDe9K1+r0006E2rNHCztKze
x9mm7/2esSKdQCjinj79eHSDdi564Rd5fVWw2Jdpn9+Xe44scu4HQzVrWKunaCOV
xaJzDDj3PIT5DkbMF5D18U7ieMbNHM8mRSQgfTHJXoE/5EvpcgspZLtvMrBAZoIZ
ArJoqi7mAu+orHakEiSq9BUlorKEHk6GMqfH2iaJzCcCED65rL9bQmY4R01yM99M
8QAujz8/iRshNDwnFy2Z4aBz5vRctT8cP981nAxukLEYTcl1V03XAPn4+pCDxjNb
xklzVa6VfAcQH3vRbyUUOwCLRsKdE06DoQ5gKeivhyejtd6Zr8qwFX7u1mm2E24C
QVvyEIhg8r+89r69lzS2NMUkz4NLpjQpJlhQhFufAZk7TCKwkgAkLboAqoCkfZCr
Dffuaj1L0Sy/MQQmMNSlb7wSgLo2SO4YgRaxa85QZ7/qPNWlHJnTc35lHcADBIe7
PGHLPae1mzEdEC4XK9gNx6wRD0ETCm9ar98RaMAMgES6XTaaanaQ319seEaDK64u
9XAEvlLQYEsfXPXQfep9vMTJWJFmFhUt3nCf5ReWzR8/fTChUbk2pLv3VO0sL6Rr
gB9Tkpbw+/ltOo/7PfsWK1wTivGQrJBAHrbOMeuX7UHonimDIS1MNhd6/+OPMy56
7SbueObw64ATVXMkX+95Jagt4zE+L9rg0o8mr7aIzubhEtG4DC0VjdUN5zF/nxwP
779zCqCS1Bi+ezM+FQ0+MBAxq89CXNkZ51IrBfN3oDPvqUvoW0Dpc/UvhVoC6PV/
jteW2eGBhoyK+IC55c9jaZtW9jFfTCZkhI4rsDrZwkN0QeCuipcvWYjfEdB2FZvn
X20Z4qH5RPOk3Lz27h4j40+nfaCuYk/p5eL/LhedDD0a2OwTXM2ViCLRJ6See5W+
1+KpggiC6T6Hgi7RGrM/x0eZBZchgoOWHx05uytk6XLVgUFXMSmPbGVxV3zy0y0n
AxTK2Y6cyolcPWJVD7xaFlPo46O2yIXfSUaNVPQH4P0lu4FjzRRnKMHib+kozSSH
iQEjnhHhemSyoW7oTJT0uLurBtH1KFkd0xyQjpa2I14Fdaa36NQSAB2dUMN39Ys9
`pragma protect end_protected
