// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Angc8IrConR4IrDKdxS8ZJP/gGoPKTOmVygvloJgAoYqgsPppfVdxIFGlm2Eo7UC
M/yP6/Og34vULh8JByUpd0tsSI1/+WyAbYrbOUPnr2ZOyRMUFNhrWQkW6VZSc/mJ
cP2GBMwBAheGXg8FURWNLlylHq8XaMsVGipk0WDAHaQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 123952)
w5bNo4AHbnkzyw85Sz8Bmr8K9W6NKZL6uQDfLCbOshfUtPeaLu+0wJHE0Zw2FWDC
km4mwNP3nz+RLmXT6ip15JbP9SBPxBmJEslAMFVsj40WwNCscr/lpGK7dDv3Vriv
NNu+R2VjQyEUS9pbERa1hnAMFai9mCNL4WWr5ZfGaR2mQdvja54/mnJceUW49X9B
y3Qvp1kWEfu3HQi8aOD92PtE4yEQLRzNdOQcQzRdEULYm/ogk29WFbPfgE1jsfck
DPhKnciLgsMgz8qS7y69j0rg0lYt4PmuXP67sXRBDvR4qfY/IDyxeSCNTiJrxM9B
kOAkE6X2fzawwsTNeyLDwp/tQiCQ/OR3j2JHAQIvJIg3Q3QFndJXJ3rBEnuOOttk
Nv0oqGpvGc0A8T41AiwVh8xvleplYj1wq9gVWqnomrHcAPfsLtH/YEcNCplmwfIG
aGBVOerzY/A7yj9D3WnQX5QG9kHzIArEIqSmJV8IbqHK2UXyak7GsolMXsltP+YS
AaJEfMCqoumFHIcJdZVFfJ5OLqDrlpaKOG3gk/2IB9L9HC0ibHTPL5LTdWNQwAPg
jDbf6+mU1OsylW8sSN0pXSsiKe2oCCOnKlK8T47mpCux01zjXUiC+dsKl+qtyyx0
tUVX+XgoqQITV1p+QlmHa25Hc4lfg6Sq7h1u1qUdxPU00jnV09ga/vUiRA7UaRWU
yhmXf/2Ny3Of4OeKKTiDpFfkeFRlLRkLb72ld5P22zoSXQi0ukcZZRJY6zFAh+HE
G6237YKOEPLZ8IRsW4LsPJovYmY98K3+O4/DgHM6X/qU7qQUe7JX+RJ5zjpkvkVp
YWWTqUNZeKz9y9BiXUaPTALPJF26KEF2zl105c9nHJFbR5ixx0d6X1Tm4NANKJff
yj6ePhs9eREvfJq30g2bHPFJas44jXtM6QThJi18w+Uczk9tzbMUIS7gdlf8kpwR
kxo1+5SNfpaX4paiUFZMc5AzITFfWv6wGEnQT87pM8FO5PSw+txIiGuiT4O+or1e
Qpq61GX5TZ9vaW5OLsxalLkwcvCQWC3QJCIFYO45tO56gTlNxkWvK+1ODmtH1LoZ
wvOTZ7iDwiq64pI64c5pCjtYRPaJuxlS1mG6Zr7wK9u4WAVcmC0w4kQWHmudFAca
XjITWD0Fvg6fT0g5AGQy7Uznd3z/+qkVWK3+sP4l3FvuWzlVuA5sLyzZsuau8b+S
4cYnDw5a6dgxdXwUxuhHp/ph1Lx2nu6pVwJJORyqErgJfdq8lyg4PsKT4XRXePdL
HVrkQ59KXnUhX4nbBPqvEqRgZKUD9RdGNgXGFk/I5AlotE3ilHu70luUc+hP8xam
ZETbj6xgN+euU3RmXUwyVJfCL10M8nnAr23m91AneXbw86UTICUJLJmiwc1HzqgY
4uMJGEFrwJW2+vDBYe2d8OZGALGFOlECIpUwEYPAPO3ixVQEfcCK3Y6xTJt4LkMh
zu9EbLdEoVF4z//P8A1sOTuQ38UYaVh6HVNZ9YQSzmjQX/bMDjKNLq2fuJkHJ4sK
r+IJCQTYAKoFc/PlvINwfLO44Y06kBLdlLASkq+YPlvr6CcB4S005j6mzHcSYRuc
NdOzc09FEl501DnE//ZeaMIx+IUKdruyaDgd6Falrpvat4qZ7JcYBVBmnx1KmDmm
cn+0z5ak2Pf+ugA2/Pm7KJfjw3O6UwmQEUkqOtOUyovoQcg0+vTf5kVV95uymM2q
fwBDc4OiE979J3cZk7RVbK4YjSZhEfxcLtwvMP9GlcEPipXVo9EwTSrOS6py9BPB
EM/TJ9W2A6IwkJM3lhB0lwWPNeWabjTMEgoov0YQ61yrWpUyvCI1uumOq2x8+40I
Wy6ENmm26GBO5uc/+qBJBkshE2MfyUvaQkZ2fuISaVtPdiNlxQgfIZbAVL74ECpo
u4WJIy+fC5EzqdK0R1JzKaFGOjcH4aSiEWXfWrbm3XDrPXTUY5f6tCAx5uAsMaNo
D0GZbVhvLN3oQFh3A1zCdcMl9H+L/HMx/IRr3ybdGd7P+hS7YcBvmk2lJSDGf2BZ
4Q6cPoxQc2nYqMU2ZWoTN6mNtmIiSE+sqR75+J3ipcLae9Q2yRiA8qbkvIVXWfDs
1QznWVWiTrxi6uHCGJUgls2zl7Px3Xm1GD7fhbJVtX92EURSBBmS1DbuUv1i7XQC
0/6uHS8VfA7X9BY2UMHMaEKSvl+HDDvhxkDAY55IqW4DMtSslCFRtKu3ENygZKl+
dMyXRaylAV+TNPotqdB4kcbtlsHJq2BEcAnBKzrSULPzDNQe8YwhjXvRfVMkad1n
y1qGuXgj2gnEsL8qSad43X+m9NxgDbObNseR/0im31ZsJKlXTiBNy6YQ/ID4qiID
AS8IBDIdn+UD5FHYmbx+XmmJNofufmkMJfR25F6DZhCO3Qy0XeMluZzqUUlmJwmI
ZOMwuZ3/DPuzm/cojHTHXyoH5lMsBwXSxl5bkFhabKueEhAMHEqOciW25ldExN07
ZnkOD6y6zHpj9N3+De7yZLc5i5fC1bZvqOKPWl916ScWwF18uBJYd22hG4KHkZiI
IVHQnM8ZKm3aM7X4Ux01/pW4g+BBxb5qg0a34NnqAwBosM8hsMdlK/eDo/3OaTvO
ltAK9RRW0Ttk9STz2OqEa2HyASp0N+0fO7AhcNUSd0az9ejLo+Q9osrSAeZZOFm/
/LbkEJwjfiQzTNa2JCe6B41NqnaKTrVQLv3aRdNOr1GYe7sozy85CZoH/77LSvPp
nmXbyTkyq37kgvdoF/G1KW3lpV1Zz+Ch7V2It2FUvnSSx9h1uVR2LoWWMDoNfXAK
XgmN9XA3ex83YHcn+xaSSpSAZ2mfjDs0U5Xp6fYZkRWMRLytuUwBFOen4L3+h61j
Lhh0yGyNsZ0IN0zlm62x4x4a88POwrqLXQkryyuDh3WM43MIcU5Xu1Avcc+ezWSY
CyJwW7ijyF1KmNuCBw7ahYNki0ZE3ssRCPgizTUF0x6wdnXUmzBm1kpgC863DCKH
6MZ86OdbtNYyZbJtx8zbDeYvqhvlhzCctJVElr7cocnFic50Bjv86atixd14nt8c
lsFO/NYBEpja5ea2HmI5Cb6AzZQ0pcHit06ahVNEie76c4M+6ODDAHmclpZzQIKa
GNTo3dPjwbzvmeMRtuJcwy1Gk6Qal2TFBcHCigV6LXBvhdv1UvVYifvvk6l4fVkh
2WnwXQyx8BvddtGc1YoQCBCSmFzxCWkzc0i8nfjyFjvVn/MHv70KGFLmqXIlx66H
O92JjLk7My6yHKYjJ7lFxSa2DDy0S6miOtKej7eEld+B+mcDBnfiHEnyo5C2InQ/
tkAqxREFp3IbJksgDyFWi5JTwr9OtiMjcPQDglhbLIVSrYiyUDc2S1e5XKMEGzP7
urIQkn02UyI5ThOFSiSc/oOTqfgYmR+3WLhoFuB0+YQLbuw80RIpzUDqFgIRyg9+
AYeAHvvMSSiqxofUAZfy44WWi0hDgdY8qhDg8eCikKrG5p4/SU7fKdEgx0SG1e1s
bhwkl4ZBvEt6CFjTGDGrVxr8osHrIjikvKPutEKR/cWkTWj/MpeHj5PbKfRXMU1o
AAD18lYsxZeS2gAG4VjNCUgNUjX6GioLTIk3dd1i3ejVYG5JQuSP0ia03RLjXIW2
is8gmQc/7E5A1X66Jy1/Yze534Oh6YA9FgwcRbLcAvLE1hb02fRwugbdL85DV8AZ
kVOMHH36Ms9rjyXRTKqFrvRlv1RLfH6HVcgpqblLlXQW0uG43jGu02WNuwy7wt/H
l0KRwxFRXsaAz9NdbsQLZ9vGoV2xl5BZNucrZOvmNrtGt0D7+1WdETPMs+6JzKq9
oERmtmU9ic0ESAfHmi3yd6bA2eBXE6zzb/WsUZ1o0fEVVKqx0XI3XHHrq2lAX82/
J3PlVNCTz+MbKhhLX3XtIoPQqeS70U8iFwFD3Rjt4ArEGbSiMh8BqMaOYhydPMsI
HKoO6WDbF5ALiCLznJd5Zjh+CSGpxMZheS72dttZxLfS93aLTOdlki5XNHlP7Ka6
SxoAbsbWfkvjaL65IhTzqtxO4XXTjDT6L2YuSAF2bMKhr2zpS9sP9nzyI4LE75fy
ByIP2CJY1bCjzmMe04xc2sH3SU8hAfSMV4QXawOnDmrpFMvxywEzcOmdhBL7EEiF
PjQdWQEzFOlKM0B4tXZAjx6kql/rVlzGkDrOfjC9jRyokj7Y0D/F13dEBBc99rkc
v0bNLKOkU01Oz0cWJb69J2P1MADFI033uS5z1Hz+bJ2+AxfKsb6IMmNjXzuqga/p
c66al21nJj+3gSUwFHi0BcfV2xhjlbmLsW1uknq9eq/yu8M5dniZRQQ0sjcs9GvZ
K++eyA9A/ZDeR91aKI57Fjoey0VJ9/L0XqiiK2BBIgxGZNFkHbsFsa7QtYwS9bUo
ChNs2n9wvjfMrp1vvaTh7lms6aZzml+iPEpujQeGxjksOxQXwIf8sXsQm8gqCKJD
49DBT7RV3xGSM76Vi6c6F1tnLPY1OwclSWvAb4fVuHk43GaAyvPCaZF4bMzkXq5+
ajsjnMLrQLAScLSrIBOYDzjtLFan+ax9h0MzOq9yEo9hw6rcCbJekJ+bpy0cwn+t
57umhakGmhL/6DpzMfV+WYqen1rxWJudcxuVyHXudcVvkh+Z6u+f+Mi9eXA7Z+sy
wESPddxvO2R24LS9KwySPqfNLgSA+Fa5MU1fLMWnvq8eT3aD9SYtRI5FphLua9Sw
RRav6fGfEY6zUn/Max6lhl6xnl/rjjiv5UMlRZX9f3pHMki1txB54ceHYLKfIocW
XIdYOmNq8kxs/dJVWjtjf3Iv53b5Xmq7swUoNgjUcXb1htu8GcXuYVPsUbkNyvHT
Upr02DxRPpklYoAjuVgxbQqB48RMekxjPfxCZIUvOZHcnnButd4cDARlOPQvET9/
zb45sCHrJqAxwgJE6kIz70wehaYtQ/93OayBnDl13qO0QE+Unp1tUgQhfULsea6n
SAdoSksOHm78ucSVeyA8L1KZ3z4Oj8UAdDSwMvfm8FNUQX53xlsfgf4dMvZIUi1F
7T/JEGOvokZgCKYH6U9IrSBoqjmoFGzUU00b03N5/3MQ82VS+PkQU3gEWCwXtPr2
iuq3mqrrNlb5/RodNnDmLhgv26G4RcWbKl4RHtMfQT1CIcyIHPRbhRHqS1CW2crF
trFFJULoPO0CO4oCwvTb5T+h0T2xYX97Dvm4ArsKqxjXq4Tr7S8gHdZt3GxgSdCx
2JUZWCa835cnYQdbHUORpTxZUpJwfkfKAjEFTKjoQxMOjtT1+zHQCb6PG3IlldiK
WgS8+H3BV66ilZrC9fom+REDFuGCqxH/OKa8q/sKzBUyQ+4c9u50FwzSFh1QMeuG
0lhx/yTHs0/4srHAxLMrcuHDEEhS41/kyGL7vnPb+4Pu1IcKwtrqswyRM5O+Ez+R
Stc+CRfgaaSJg2cBNOHRG2uQlWDqDE1ipBZwunm0DOdRs+ADUXwNJLoaGVXv2x+A
iHyBdgRmjEt7LFNWYvrKP2BwK/Gd1SmgSfuJ5oskyNpprR0RJ9AmnDhODOAXSlW6
v/h0odt32Lz7NWkqrm6IBFRa4xtrNXE4Z0mn78V6jcIqb2OhiJ5xjzZKyyudZK3H
8YDvpKAD0P0akQx0bOJSsKB3hjQSd/TmgNA/Ljx2NNFr0O7mtBRoCLfCszIS9M97
0r3Frc5waNy4LrtK2aD0tN2fAqE65h7F3YZHSsLrjCnmOKYJno23Juh0upn4mkpt
OmaKhE0IKhz3n6T1Y0Dr9hEyq1wO+r4uXxbW3moVSD//F+4Ueo1K1aPV9ayP7xuX
O1EK99guQO0Kh3w+IZ6viEpr7w3Yzsv0Pqg/0sbWlzaFi0cgGU2E/y4M9hhxetG+
SuyuD+xOz/CvrdDC5eYN8hT/4UWhil6AZKqTN7Qx4REH2l7F+PcOVLPAFHDXEOyw
nPVcukbfCp7QlIKFgPswfQOTVOP0mq5YnWy9SyGLlWCAAZbzk4zYfEzRr0gJ6olU
axqhczZxMCWsAUu6V2EVDuwDRKMclLQ4UcNLBPY4z4lMNlMGt2GSb8wPdGunuqaM
ztdegbWvcK4xF6TM41ErglmPCQPgYe37N4qG5xy0uqpz7tC2zcvk4c4+twFJztkz
CQgYXx/BSrkE0XaaykMdbDkJhMAIPEVljIchlt5ZZ8TC2jVxID1Sx6bso/eBmu+t
bOZfYKvHIBjU7MqCPcjLXv0kuwqEMtoqtPE/0lcjQ7Y1Lrqr6xADf879zS+h7Ltn
EvEwHYhJ3yi9C5xm9M4qcPPHkO8xuZgjEV/COzXHO+lSyXvFE4TzEZjvP+/hpkPu
NV0dQmudr3Ywpu/S+OnXfLO+baHvGtqHyncMG9Gbmskhc7xj7OCXvgvxl/Okiw0H
GLnj8oL9kTgJ+d6xeILQrO92q1yBToyqbfgaQFhHCUV8jV+6EStgDBDo5GJU8EJQ
xhs2tTn5e9bvuwF/Ql7WzTHFi47h6o05bROfSyFKp5rd5aFxdNrZO7syF7nwl0G6
3ivSN2PYTC2BZ6hKrv0wOCDT13C1DMsZMDLEMDdR+wWPilko08dDmjwU4HwaLEKT
Fsk1pHYdOkpzx2+WqEKobGZG66mP02L6sYJUzbNN4V/kH1tCbw8XE1M4TCqs6Wlv
WREvVMuRGDS/7ElqpOEifO5+xAOm+y42q8+d9dutOayUb9sIQbTwGY7zA+7jgpIA
308O9XAKqjMRdr4Iv/zLFMNkUanZ7hsW53hCc1Qh2CcULWHIfNAv2OX4WZuW6r++
U8HWW0Z6o3HBRUa44HSmu/UyIesyymwOad+JvPobiWNONivcP+yMf+lDD3l7che8
4ecvwqS1uIQOrwy+WGMubVVzHk2SuEA3FONxQdxQ7i8Z6TH3HX/zz4XHWciZwDTn
491FVZWshS1ygQkuYBLkJ7WQN6G2V2B3R2mqyUaqSimx+a3sNVj/5VxtLCHBV7Tc
JF38tSyW/Z7FVEV7rqd1Hgn3c9Vmze656mAUbL6I6oS8GoRuyrKzs4d4t/Opu8ET
Lse/Ubr7XVcN6roMWg4HqlP94lO/gQHYNASwcLABQxhX0gtTuxd/7ILsII3SHnBS
1ydF2ggtaBonTZ7haWf9F0tlT/NIUK6y8ejka7LOEQ3RkwtT1o3jgchJnQFmT8dp
UVC/h/JtTSfFIM4Ewm6iYjWPg0R4YmgPRPLbtrFVqaTCVAkLzs76K/nanJbAzZu2
mRKAZVK4lPUO+MQTRFwELAeg69PE4cY4g1AuJ6t6P77KWMSPwqY8zmTyxjR4CEmq
uS3dZVDJLTKUooh/z18mzc08Zvrefk2EIlyIL4ElTLmPaXm/TdkKGI+FvLQzQ2To
9sLL3p/+pfZP3K63WgKJEeBTkEYZCZAiV5b/Ww08gmW5rwi+yZejTjXM3jnBuPab
YYt8ozqlIpqi4QTb/UD8yKufyQiU9shEQGiYOTAjfthUg84ix2hnLmzz4iTfAsDF
YmrTiaSsv3HGq4vH+FZX1GbAZ5BQRLpz7DXsDwzVxKgNVAf3zPErzVHHndxghkMk
sahGGYv7vik+TweEMZg325L1Cf9qSl7k/v7Bln4oai/pr07FxirmUH7eoSQyNKf0
NZs5SiVipW1AC65073pentAXYJeSezyod21sV0P4yYz0kubux+htdjHBLkpniKIP
AYTg2nUZh44cMFUfexdcoGOCro/qJyYDuqS0BkzxTjHCI5YOiHV2PTk6y8nnMxug
GTZGQHpv9EdDgqEWgV1iEGJQjGjdGdsPIfY9LbzG37GFETN8P77pUVpcLGHiFYHy
DV9IeRXWlD0Ark5R7l00ii6/Aispzq/IFB/FDmIgnIk5awK08dsW2G6E2Dp6BHM/
VfmSBA7u2S31+i8S7BgSburzTauqCh8pPx/lijlZpE7iAYUskSlKRUg3wGJYYvf2
59dJUsByuEjFB96RvKoQQBQEneLm/ZzR37mc5VWGCSXMxkEQIM0MSS7j5Jx3Sf6K
Pjcro5pey7EJHxgCdAvAgjoCaJinTdVf2wrqK6RqgWGwpk0K27/V1FyJMVbtaser
rhPyvoMz4jh7yhKOBaRpX7MCirq5EjEDmYijA3VS07/57RZSPBoo6CM29AVm6NdQ
tE7YI9codaY3dS4Hzi0uMxU3NgPU9ZqIq5Uhh9vkLg47boJX/WDTNosdp56ZD4ZM
pVQOY/J58JDWOmnOkkpppdyFhQGL2QoubW7pZrwqyJbkM/535Sn5aS/nrH8o67AP
AG2mffMDcCJDXrs8XlPMFJhEvSdwzhneMdqvolHgoCL3R9FBl1zmTjyMjeO04YGp
oJE9MPPrPoU9r2zhO0vBnwxPg+Ih55czeklZ4kQLbzAk7IdeXT4wzOThAemHU/Oc
fQ4vS1b8/dreBR5t5LMExWHptQweu8lq2fqAeS2sfyYUebA+Cf0TiH/Yx3PpDwqt
GPa/SlVl6MYlsO1IGQe4dbEH2/IuwnDR5q8nXNeI9ZGdW4t6icezbAwxFLaLy/om
vqD0VOcFMH2eaxE02/M3s1/6DpH+KpckwGI+MkXUmEJFISEeTpqwttPuaNJGdJmr
N4i3b4GUm85jptRqwZSn8nyUyEuzwTLo82JbZebW+chSy3BYVTI7pSDoRqWyC31P
2boy99mwxhmUMpC0ZUQX+/CZrugDNTTi+9ZJJ1dGsF1XNHT/FEMAMjuWIHIDd3X3
eNz9VGquP2V3BsHvwhz/8NzcbSYPJiqYtEdSY98bXYzaRCpDehlI7vlVMw4DmJjZ
q4iurYPHEfkNadNWR+nAiY1Agss7zMO99l8kL1G11KRzJaDRYs8fP9J6beNHePW9
rylyE+bUGk7GF4o5OFFs3cuWnmf7RHldycifkaghsJ9NF3xJcy3WbgW9oCN6npFF
O4oenFBBYWCVi1VwZlND8JwsAEfLAtKg3WYIicAfUycktSlJquYoxcXKjD25ZtWs
S7BtpE3nOm6Pj7gcPB8bPvhvtDb9t5MHZb6UdIjQNFz5zz3XaDjmfC6bUB4oOEdf
+ZiXPDJc4WfjUw0NWGzp0AP94Jt0UHn0C2DoAL9yDKWqajLHZAM8ZhCSaMLiNTAh
94jWXbb4BRcG/Lv0XruUPneUi4HGlDyzHov6kptsqN8ZlzbYBqTbnRMvjWul93IZ
6wBkSVrJv3JFjzV0+4Y0x9i5AUvRScCoM/oRvkcX4s0nJSapE9At4/00fVpbMWGA
T895+0ZnLpV9vsQ8Slh6JJyP/KNtxD0vYkDasNBz/OAt+K5fL6Yh69y+kqy3UxQZ
ASf7REDACyfHnlR+WS5hFg/j5rtvlVexmwGVyEa+QAL7TpRLcHg2mZn3PUG4pP5R
v1y0Z7iaay4C4ueNKFcTRDI2nojsegj085RfeStOdflDXVK+b2KceEgoan65d6Ny
/Udf6Ipr2tCKaTGTtGova80HozOUFI3Ji24lXkgMoszp/cJFYuoxF982rkVcR/Qt
RxeCHD0UJPt/4ZYfRocW3U4GctVJFQD6W2RgsIg8hMhIMmTJvEv1Bo1LRiNHvla4
2elye7TDj0xeWE0jewCub35+ayxq4MMM1Om9TPmR5SI/cyaNws4Q/tJRxKXQxCMv
GF/MW2eDIQAtZ6913hpLZGMJQmH9T7cB5392AXt5p5gSLFKfbvRPhQx6GNs1gioI
0WurhvoYkwpZwZpw2/5YEKtXRLSNN4WYaI8KQZ+tJHVgP6S4kg2uR4Wfm51M0Nt3
lxj0CGocSaFqct4Wyt2RgNXUlcFenvmHs62WG+D6f8qtCxPWvtRwYDhwsup0rqoX
5dBzU2m8MSxQ2eV3BvPDeFjHe/czcQEvj/MZ0AfbE3uLBK/1SfL2TLs21jx2vqij
2PyvF7SjJQmqISUEdd0y1dvYShlavC2+Ic3bWES6S7UUdC7U6h8MKlAx3iegAW8x
FNVuHrqANkPVe3uI1GNSXoN0pS7rMp7nCco0+hflhgyFz9Zf75SvcL11NTjCm/x2
6FJ7Jv29SVASB2QAoaWTk76ik4ihAd62+djhaNmvAYUkpKuhSdy8DC90iFuBxHxa
paoGMTNxEC69yyDxY/h3lGJjYFEEnqLZfc/YTObPm248i9hUGlFg7CDSTa8oPYJq
Hnm/iuOUyfmwauidM8GUbSTT/Jnu9uWbv3oRa9G4UUWsirkBTE/SmJy/uADGn0Vj
1r9BgD1gLhEVe3phtmXGo6WXef6ZBz1ekLdXqLeABEKmX7SFM6BiC0yCINEawluu
EzMI2SzOEnebS43nlFyU/xFHT2sDgmVhwL+OGvsoAhKBOc6gQTQUuVomcMZb1azC
ATZN4q2ib6NHrgGmWRB+DeTh/XmkThfJAcSPQLnLTBhAicgFJ1bo6zyRUxqP+66j
hMKJn5jBVE9E0GuC3ZT+t/yvTVxuwSCmM8YOA/smb5nEORxUNB5vPZB1xbkMTmfA
ioi2+3oX/bmYrraegoR4sTWxL1n1eRqRLnigF92phVKQGzVvok75gHR2cvD9Y4sD
/OCm/i+K1rzzC6eBKvKM4k1gwRlahwfzGJet/1KLBruWFj4zOVrsUoeg6cn0CJGn
wmqRPxpSBLEVJdBiArXzcd1bgsKpxJLmpWknGbXyBZqagVi3eOjD1Lhzi+wi9S3f
PYe35+Au/S4Y3OwPxMu7cKOGRZw02zvme0zIwBVCCF3G6ckaYZ7k/2SPTLvM6hSE
aaCD76zig9nCU45Rk2xXDZ/dsKmxuN5R26iHA+IlWDKg5yhYiUK7zWNo5HYJwtK7
2UT0FbFlwc/pLz4QXIEPSz2SM0038zBLuqAN6zGpdCmNB+0nhOGpSD26cjpXVQys
7Aq3XBtc1DY3oMNHgceIf3BFJ62NwB6wqAuGRyaacy9daHhWok+G6uv+6l8nLwyS
6JwFLXGZCM4wqIFTw/bpMNm6V4FQBkgiPtVgfFDUGeAoctIa2d9zTSoqPRHnzC5r
cqrej2HYLUrY3UD3a2B8BCOYCkwsFdlAWTveH4tV36j0pzDopqvi6d7+DUiTK0Dq
xxg3ecKOlHUxjvwfvupoca8qUIaNM8RpXBuGH/SBzG5P62ufBft4pLc/2Cj2QHqk
7U/NrlLIrU2dqai1oE8sctCsFM3bS8rMVURzDNzvpDhIkTOdE9+VYhEd+KXlMuxc
ldgFjWv1p5J4ncwIfyRsYVj0MvOhrP3B03aGOTrx9rsOuDcLroY0Ng1q+dCoDTMM
s6MUFxFADYthLJWaAy72iczPyszaH6SzFcjdIAj0SSBcOIX7pZfJmHvSDWartjPx
yJ8ORVkyiNU8zyIG97t32aHpsfCxDqvqy89Sbgu4y9bLkYA9s3k+H7ifvyar/I2F
iXT6kWpuwjRfCpblESRflj/TZoA80SB9o2Hm9bAu4Rmsrm30IbZ3N8lXfW4or3q6
pKFFRVQX3vJznPDCR9EElaRlkjzhgxgEcDxPRMF0l6v8aKg6dQiZjUFqePoZNnuT
MbWkelbIPxbdWLvDIY01ezdyYnKmCG+EuFR/9Xq0d013f8xtx7Mk1bb13MUJLbim
PQ9PrH9fyYz/ULL97E1lh65z+9E8plw4lQ9qCyCZnhfBUgx2FF+WSjHR1QlguFsq
CHE/PEFRVBqyVDUDJWlVwltHPQLDiUN6nHZDyMAo1FsIKFCHP8bY5IlxVEMSuW8d
Yk6epAbmYm3+61rTulF4okWhd8IY/SWi+qT8AW0gqOX4W9qGr3qsbAFfu9jjsB+p
A+PrVn+cc4YEjGQ88/A0SfaT0asgZHEAUJaz1yvwrX+qfWt1dLav4G6UFlxpPOvN
Va+NAbdptOFxl+KGFrZdTGGAZRBKT0B0vzMxZs2dabSuoXIPa+9pDCn6t6A8VMnQ
q+o7gjTid/ZLW4zLLAu+gZD/0wrbJGFjUMRBo067i1+pl5/4IY3DVfR1U9A7eckq
uqLjxVoEBo43E0cDQodGdUCMWaU+IOFIg/BtMUUFNLjYKxluIKWFLmdfq2/u4WZ0
9+d9Rztsa2FokVnBA7h/jrHaLB2YdvH4xKpW7ZQwwEeoMS/jVGmqhQYJh/4Mv4bE
2yXLxhd0bkrDVxcQMEmfhy8Yh1zcujygKdwWRbneKEAtKj2QHjTTdDKDoyrbN10S
AJguBx0ghsxEJeKYjB+zeNIrUsqNlLEtND0lRQ0pWd7AU5uzJI8D5JnwZX7Oza/A
demLjt3flzHAn1OulaYf4dAnBdmG0Hfg3ajClKhGER48Tfwvm1M1Bsx2A7s9P4J3
IHJk2xKN/Gj0gIFxou9HxPWp1scLKArx+zLaHxkkNGnhmQiMnXf/UC2/sRopqJDJ
6RRFRgQrN9BjDS4BDErXFjh5LS1jQZcErgn1W4YqYEmZDXkIvY6c+EH0XDZtLKJ6
yY0GGnZGNIc8MqJ5+Jlki7nc2PxJfJQpTzM7jwnJbmjEj7k+RyGEc8KjI/77PBrU
eDZHFsbGY6Z0jnkUkv9x6Se9ofxNATz4weVfdRKFzd6HRoik5h/sRoV738+GotXt
H8XHpMD/Qij+JGO6yZkXEez4/Ad8TRMznUp6jKbUYpCDnrFRdg0+wB4izgD0R7dW
zA+L2La1c3tpx0ubU+sao0bS5nMcGC/jLhoqESd8UI2QDKoUHeAJf9nwSHdAUPat
as0y99H9odJ1RgfWUQ4Z0/2fyGq0I8aPhJGCbNcl+EoPb/hh22pot05ZmQi44O7E
H5kdojL7EyM8ZBm9r5Ffi4BgDQpnMOmfA8XGeULmwuCTX4OtN0WuE9kl/UO5YA1c
E2jY2NC1Q3IDik9bYTM0e4WQdNiGvpAYHbcXlHzoIdtc3vBio8J8kxIRLQH79pq4
4jHKfPoYt5yxYVjaJpSQTrFtHJxiZQMZwfb1YFkOzWTEtlcYXlvawNGeyKLZzmPi
PmSTZsGDHbGu8Qeja6nUY0uKAfOMxL29RvCqkVWoaIIKGfxtvXThej6WghSQlIrM
0lnGtpahpFP5MCuQrTMgDyAv8AUoAghbiigpU0Lb1HB39mOBYqrkJR/AT8MhhMTE
QlQgPjmEwmwp7Ya6ykiOLfL6SMIuq2W1jfuXsa0fGko7wzVL9ZK0XJa6mYi/tAG6
PQutN7LBEhu8Yhed4zFNwXXlVv+nwvM09Y16KDN5iqMVQemckkeIwfI+d9XhjgCQ
vo4Dfg9pACVG+g9GQlTyVSZDTsX4Ww2I84vnSJd2+cEqUwIgXMD1fZs7CzirF3oy
o/lS3mXgCQPi+0+8cnhszZBuEeYrNBIdmFzVpnv0JkVDqMwyhXIhaGU/MDs76XGQ
Ns+Tvt645sTJZqz2XKPCmQ8Giows1taN0eum/s1yuKe02/SMo04yoDH3mkDx+efC
DFB+uRw8VfXTOT5n/AidpvQwXdnUt4eDvGUf6F2Y+oPyS30Unv8OaUh3zSutLejl
shnGyWuxymp/5ifBeBxWGTA8jDi/wf2oJ3Q2NpQ5uOTb73osgEX9Dbgvlu9tKC/q
eoWd45u4hGG52W5xvSDO8Sx1FIRy5HLGmaOWH3Jgj7bLXSjrcK0AtD0xBJQZM3ND
QGz+GlQkmLUIAPgOZrdArlt4ukJMevE+o2dtZQzuO/dmgClF2FuRaBGPFrumMsni
IuOoSgx7sQMdPIAC2iB4eKMryIIcxrbmYohw1DTyQXzA97SFXKezWWPW7RnidDdM
ESd+w3HedYx6jVf8A8kQm9/Eb9APK66//WwuXEIzyZPLQzvePnNTsAHrsO4vMOur
z4eTy5/iGAUc8DBNgnc6jsPoGVK1TBv397ft+3JKAdpkYbEEXtNc/aDCXt1qEgYE
8l1Wmqut7481lfJCiC9Qiln3Rhwkf5yKDAOZxT299bdIXjfphqDgFypYsFpHN2H8
PPiErq4NqEVsrrZMoSlDb41ttbu8W7+3scJe2htu94AAc6/Y63pbNQ/cO2D1m2ih
zjDaveKUBGO/eEPm6fOfq2vnM127HKe26ONLRjpRuNV3q+bygahwOVZDBvbtu1fW
3XTkqySn148idQQPErf8FXkhAd480t+jBlXkHt1qRgjNIPnTdpspKkEV2VnqFda0
epfnAgYkC2jOGW+MPKWOigd2n7oKTRTLs78V/S2oVECMekUED7Mk14SzkJzQnB88
WH8ukCellgyG/vQCELsgmQkiUGB7NBgUuX5oE/bUgQRwPEbPtslXUcT76sjah+QY
VRGYGA4+Bh/SCiwtm2YmNaWNNX+feeoAiK457i32bjefbhGq0/63+WP8qhAHdBEy
6/JQ+SK83qZxO4VLLfBcfQqUHwk0b1dBhlNSbqaZrnh7XihNuJtAxlf4RLLv5cLx
rMosPOBiF3mGrSUnsu1K+QUXz1H8IC7XfYr1qPpF/NtoLoqP+l4DKbZclti7Kqb5
6lPK0c2TDyYa0YVQD90PDR/HAJ6assrE8kppZhgkTrDiCNQM2SWq4KZIZ42hZeM7
/F9OAvTLCI2NUOH+gv16n47L132W/I+hQz5ADJiy1bRAaUzRlj6337eUp+h5HbQv
znJHwOzn/Mc/zsWT2Xw/ivv3KJw8Vbsy7SbJNJn2DzoZ8McsUdurcZOQc+2LIz4D
a/92a6f3ptw3nmQQO25sRvgbnY07xflLfSSc3ScxQvuH++Yz1QxWXdSdhJaQur89
5SG+ShtolJAKnqc885kNwaQb2ViMxNC7Hv9nnh4i6pGc0+0IW9QP3JG6i6KPPWgd
4zIEVnXpF4bz7HvlaOtA46lbUijp4I1cOf4NOKVC8WvpgVvwI2afhjl9lcie8ssB
stFTnU2H1eI+HfHxVZQMhyZFYh5h2xKqEcVzoHRA7bgwMq4Ubx8Jokgrrn+DsQAy
bdKR+6c+ty174+PMQqsznSaA55ro+a526NS6NZ32x0JQBLphKQVqB+K2BNCJLD69
gyfAhRPvD6wI+ye1Uol/X+Fe8XcLrdrqSshJyTiqYWuWAIuB5hlb+5xHoxGG65UZ
BMMeDLHYiYXCiRCOTQG7gNekpwTdnCdDnIZvqBAXUEwvt9an9i7yx47bfpCHyN1A
I/GAJw64BkP13uqGPV+FV24syZ2EA7TPYR9yeKZGHNJJX0wsZm0vLrqj2YhgPG+Y
iAS7ZAc7YvAptvm9fGQqIOH6LIubQd7A0gcG6h8IzflcP/ZaThSznoX+9vFjDlCc
6m66U8QzDE/OOqgEr/xzPH+TS/mBmZ0YKTtaY0sul5p8yWdkqHtVayJpYD4+Hlo4
HHAmoRfQlOLPbabxalxkcmdzVrfQrjrZzN4nWfk1ayqJJv5dqvgNdVWlx+55CJx5
plRa/V76C7l5eqXrhfwxm662O9cEiidQUTRpaPnQ4Ifo9krxzIR3/WIEQEI+TTnP
8FdFpVVYWQFOE1vUVnB2gzQZeQTcgTpnvwcUd2bN7C9xKk2p8gxkN6rHh5wHR8Ti
6Sdxi5kCrEguvmTljhdWzw9O1Rfb9qOFwymHCkq86PFDq1RavTHmh6DFDQ3loTTx
qFczEDisQuZs6ePitpVqWXnN8Wyo4wzWxOEpFodfxrG0tBMAocwmKsnvWpQL9Z3p
PExuPbzxfIIkwU2rivfAxhEwL/WQl0Z6lzZbCKqayMBeQm9XZfS8JdJlbaUvbzyU
+u5KNZAjv0zv9owlcJgS8QjitsbOYdMs3wdntZQs9U88YMZETTNnnvg11GINt5Az
eoYJANzANfF1IHP2PA/XqkE7irnSrcJQc3y1rL1YW6NJ9OJagjuqcMWIUy3cDRa+
WoYrghxiygB8PWyWI0vBh40wAGRWRV2bykSvbxjdoxCm4/lZjsT/GFmv4/8YDWkH
Zzo/CrMBl/xQCxZQ3LrJ3fp4qxSFMMYKm41huybhDrctTsyBOh6XYY3PaY+qq6Rg
QGJJuEvBrQT1bqKwIssMP04+HuUVZRkZouch2IhB44R5RZIJUE67xto2w+M6wMcl
amgGyIrMxOjUrK9nnJ7r1yFpCtelFLKMPYoDHpLVRX957Sray6WOIIqg16EFOlZa
lfsaOfI7vdldO0gfHkob/5Gym80IxGfr24xEjfIjCLK7Z8DM+jKFH7iFvfQZ5PnY
cRRVULR/t6FCwAPLuK4eWO/5LGklddTT0F2bFAGyAwwN1btMKTAQVUPtVeTAcFya
GdDxp7ndlJBNJjPIAoK6187nJY2uwDAphNLLbsv+bpm0iih7DehUIwFNm1wzr2hQ
6xJOmKTpguBIF4tY87UN3YWRa78z0l/NBgjjLmR7hI+qmxGbOen3bydtCqLEXEr9
4A3RHCdBE1HKSMkh0IVFNs9GiN4ROVlb2EpAhrtmiQ4/RihMNLObXfi13Aw8M0L6
X0WoDNM6cYjE9FdiDgQnMuEGK7q15wI/8UB00dvhzsHGaiIn85VLe1XeSdOWeZ89
/bD0HcCmmU23aKLMGVgZncELzJoE6HGz5K3r72Blk1PXxZ2zBIcGAjWQrrdtB1l+
jEtmugX56zUSCcKW2ulqpX7HI6NBzJ+NRLlHic47/eNVGE5nZJ4d/OJ9b5EEdV1S
jIWemjnTiSsZo9kAsEH+TlbBW4Pb8mNnJgr4yWctXKHv8hZ3ToRn2yarNRCz0FHM
P/hjeGYiV6EoRiQcapQl6uPrUEgy6ANgtBDDBGOV23Uq61zAd1zgl/nUnFGEoO7U
OEXdmTucbCFSlnG769B2FAM8oGx3LR5PAHA3C692lFjBrLP+Pfm2W5YAcPiLjwx0
+QT/z90mgOaajLPtzUpeKkdL9FienL7yxuy+6ETxazBBRQBguLwgQ5ttjWOeDnNG
Mv8o+hYP5bCOr41VGx5Gr2+AHW7bifwY0yMBBNV60/5oTwl8vka2MMRiuVt8x95r
duN8aSxMwWlptrbzrvAkLQIo8IbSIzEjY/s9uQkvAXi6Seuok/Ey2H1PsFVqexWj
iH/kl3lGKxuuf3i4gekxeblV3O5el7QTb1g6aBbWBfHQOZlEVH4+UKYURH7Ut22b
KLfR7UDFTL42IRdqdQhdWgaXWqE/hnt/pCU91y9Qz/GAUDO/ukt2/0acrlKK/1j+
1Hve3mGECHC3nzaapnCYI04BcH+IVhu8wX4VY6RSFcCRVQ1pj/pSLdoClU1EdAf1
cenHjmqEqPDhAfCRKLbJcgW1z+sXwFsjSxHlI1hWnM8ajKVTRF1FfVBShx1N9BuG
DCtqhUengdWxqPeT4duiMU7dv+USLKe9xJhGkZtsKB7TVUZG2Fj5uuJzESIysPzG
v3fjqMt3qOoiRtICA5BuuuZbKQDy+xp+UuliXd2/QqBMPwairFqxbV3hthRuryet
V35vBFIYXms7CjNqPdfiKjyn42pOC5nvRbElN7E31/w6WuTDxgXt7VM+kvCuI080
0/zeELICYSrqfdu76VSbIQH5p+PF4E+OeRq0327SjRb4bhFXd1N1RyINJWtQbW9f
WrcipY9NS7vCTaPhQHHyOE9FD2z39gLC3FLPvTAP5Gk2Bo84msnUbjPJ7N15m97F
xtiNcmw695pfe8cTn2tVEgV2CKz1/W7px8/BMlYSOSbjGVf/Cpm5dg1JPYy1T4I2
qCWqA51w6DqNISjvjsw5XgZq9865iJCQwo4IiIz6M7XGQ5ahnV1lihsBxwhLpA/V
x0ccpr0xERMpBsYorWT5YIHzMThpEzR3m9GZVjeTV2WxknHf7cMUvikXtXrpYPzC
oiE/fEH3Si3hxVRKoAFzojA54EKZw230INXDaOq5IUUEqAW7E2mXBUA6A1h4lyk2
WsYJVQqsFkLYLH0QZcnFKetFqLKrFXGNJ5bowTKLeSlQDPEmMCudpI+hjZ3oaPJI
0LzvRC3DCi5KpMn+AHREYteLhvcb0M7dw9i/D1T28zL/4XK6xnkKjJxp9KdK4q2c
AEOf6GIbLq/udv8Sne6q49B1BjE8oz1odmSJEApA7Y0MYDz3lCHA+81JHM8Cbq2S
SzNi8S1zPgqP0QhDbilfdGahXpvL8TBfORZBPUbQUKzy8fHge1yTYWBDWQEKCmLj
58Rd1ESxbVIhU7xDhOVeOmBibe1f3ixcovcCTgrkyyLbh3XoEG+kqdS0yMTvnGlk
LBU754XhWV93KaFujsS7qGdw3vj93IcfuP8VgcNrvkSQ8NBaITf0nB6N5+v9OOgG
P2YDhOhspj7hYPgIDC0qSlmG3m8H3hOUurK2PiBHyKHJIumjm6ZYPrAMo//kZale
NYpO1JwTAwWLbGYYS9klUsgfwxNjbFo1DWitKtQO5FSWEOXLJThULxjyt9+plu1h
EsjwTTBk2RYqvk5e+Ujf/gojXaMCgCDwk0xIAjoYdw+Qi1M6fOvn2zWOfIEotmrB
1Jmu0LyOMNlKvpD/IIGX6o0EFgCGt0cn/q54fpTesUoiCA3t27uCSDl1r+tj7Djb
YGIi0Lb7SibP6uOojC7otaVfB2kj5aAcqOWPVJcookIKlRdLUofh88Jfia4OUtkD
BjJ9XkPSLRVeRTg/7hHfl/5/gxtiDI95KleoHv6/9fadodQlijamnyfY5n7L5zdk
n5yA8SSRyntmLhBOJmzNDTonxv/OBD1Nzql7sd0xbHZfWCq6+zUupryaUW04yDrX
DdLcWjJ5aYhUzZPTcllgf+eyzJJ8Sp8wWD8Bn8TtIGBciTPiKtR5igD5b3LylxCZ
oiXYbY2C4WjjYcFplLbW6etsOwHHQtY6D3vUXI6c+yi+ZvG/gwaYqb1kEHnscqH1
b/rP6UqbtHNZkslzUxVovoBwCx+ip9Z7/fYdJl+Y8X1of67BDcb8jMTo0SheIm1Q
IuUYgbbeRAo3JkQ03v0CH6WZHboltJlqCfvEriCOrv2X8axJJQbPv0v4y6oVwp81
7pTweEsJR0imswxkGET/y6afZoU+kFtWnbYXqnzEqv0y9OhVVl+GlLPl+H0FDrW2
A7pv1QJAvOqteOLulGPN/WvBPrvx0AoKZJF2QAqGsNXqaHtT24KF/oDhjnJ1u0pk
7/EHAOxqma9J7Z3Q30TeMjvN/e02f4E58HtOQZcGKGXyjX6g7qHvIKfNwEIQ9phB
yzDXN1BEBmD95sqB9xrvTpSMIsRWc3ETHWoi/upon/ueqFbe32mAu1TRFx4p9KPM
oIu6p6OqJug6NpSpFHm7J+bZkQWGHGOy/hUvQ/q8hUF4ylD5QivwHd3QLQhx6wS4
0W9XXBKX2k6QTSMpv8O7VKHLZpDuAQP/cBTwst1atUKKAl2Vvr6OKm8zu+ccu11q
p5/nLrCQwTZb/toHa2tWaPSQUAWiEbC/dIebsBo2Q3h+nDkzubw7ZrzYcQZm8qZz
DKKt7n/EInHJMD23/lP3kN+Wblq599VXWBZqfopt9gL89d1RBjRT8l+sZPyxSIeX
lg6PCAr9BUEC/rJVUSU2vmk0YA5LHWcaNinD7Iv4xB0kgDZI/e8BsQWol+fvDt9T
lAy7Y53KtMAtaVrPMGPIYojGZmdVc7RHDgUXOU2uffahV0ou+zBnC+rYHIA9sGNq
aFr+xxJ3/DLJH5ZvycuFaW5pY9+rEwTiV2WDuIPYb7w++o+uLVmUy6C78yzJnC46
z9bi26Oaw2CJAeMZya+hIrISwUk5DDrMLAllWS/N1vNCNF7Mz9mu34KWJa+UqODa
9Ww6JQh+LQDeAgQGBxD7NzLACBy9c/REfJfBR6KGItUQnBiSunScgJJTbO1NaaA4
kYVaD1eTqISfoHlBlLxOSpdB2HbOf3ZSNNnVen2oVX5QL/26BodDurc0BJJqUW75
HJ8g0hShzQERSzrZxNm3v9vuqlAhzxIZFFUMpXNfaMuQ5M56BkGeP2viDUhND+F4
mtEunhgryt3/Rtpl2bnTB4HnMESNcaCB4ZL4Kk/uoDUn84++EcNlGMjj/2aN2Qto
q+E+1S74et5nIWYWD1t1ZK7XFjxQUhBHXIzfN1cQ1tyIWcx0y1Dq8+1ZGrbElze9
v0dfTXeODVp58Lak+7WnTtSlb5ny6ymo7T+irqSpkdgtUG7F2vWRtKfGCIVraYz8
8zRamdrjMqc5igCA3Gk5vprYStzkpp56K2pFkEsN5DlyQCuXYWgBPUWZy2mm8u+G
o1o/E7XOtTNxrjl0LnUhNaBRaxLhv1J06dEV1wR5cxB0q/Jkq6JJd/CsKMnEpf0F
TDM9YUNuDaqQ9BTkD5afTh6ULYLTTfAqL3rmr4v2nYdwVinkqaAcgEDieH1duUJB
pSZDdj8AWu2SoH5BleXRjcOGmQgnKW96Ylu0Yl/cBvHMnzVKEMx+fIrwGMnA900+
nHyDhLsyijzAVfekSHyVC0zn8EpVhO1c4nKaqz9KCRXR6z1sFkWN/UWZtWp5VxGd
y4x1TuZ49ZMkw+LMRAJ/69ZWhFIMUqaTmX8EhC5hssbNVonr8wXyUh9romZtxRxZ
cJLGnWqF0v0Vnek4fOrnvcrvq63mofpK/2B1C2mMoakGe2+Pcpke+WnGsXsPMnoE
ESeUgcI7z68BLfvfZo3x7U+pvEudrjtMTsvUmkAr9gNrOQ//UP0puBjG4XlVDRiA
8ZaXAUsa7eoj7rLe6GacXLiVvEYXX32E6s+S+nbSFplPmix96lMmii4WAfkmoaNG
rasm7IjCghtkhhQnQYAvaPZ65EPjQVqP/60nL1nvUJAJ+0TwhTmyMrMt92+eH0yf
x73Tk5180VMOIpAtIBCDmfoz5aFIB2UCnoqX+ytmBk+gZ6JgcUzDmlGwK3soFbb/
7WgngXSxh0hczTWB7kjhK5pg9TuG+CCHoraFwY6gv+AAvLLGVPhSsRa2lFAwvL5s
GmmzU6Fmd2XwglKbV//dhMpqijoGIIACbykVR+L00aohJXvNpLzlqG9nWiSDP3i5
U6b2LjtTo9yNxOruTSoLBZR4lMso7BY66LivZGRZbAS4UP8c9K3vL81TeYbNsnXQ
GrMlI5o1FL4RPGxES6C4kbGUGgcDGyctfTyu7vKujCPtjX0XsGoC/I54hE6OfQYO
9hs3S9BwafsH1CypTWSeO448j0DmjxdTn/9BFiTvK2e0rCvHU8pLoBEnOcPCmXYA
lbo6Rs2PS9HN1GOyuDoB4R1UO2CMkHeCs+bORTeSnaJV0dm0YLQauRqOf94qvJnE
I9km9WAXUNtd6ur3T5SlZ/ras+GdWSZFm2FZe8nVXlTQPE4xNNc4bxg/svYxvBQp
IPjNiqyzphuL/0Dz4ldI7yDJELpUXkkBEgU4jGGxMTld+/8Mw8vhtlX5A6+x03c+
ZdlZRuqitge7FEx9+QvnaG6uthXTiSsWVE0SRL9vSZF0UfeotRE7c5/tDQjcZXb1
NPDyT6g+rJZZcFzXE8L110hf6jhccYl4GxS6V2RBhJly3iGp1dEzxHfU/Wqfkwjj
aJR1w4cfAcRnNdTchqtdA6AuK+5D/DGU+8XWrltD/HuIrjVKHofLRNe7mgF9w1qt
s7dRO46bNYWPMwZTO3nC1dFlYguy+tVgiWs03hy1w1Yfgicg2PEotruMpFShmC+E
DKIVFZj7/LihA3KNb43gM6w4YglUepwFMEIGtlG3cMdfE8JSgmRcxkhhEom/wQdO
J1RNIXyslDGQKwTnggaUN9djnSEU7Xe7hhiKBEebeAW+pqdnhVXaxVSAQchBhKIO
jzz11sOi127sRkmemDuUGy6cDUtgUOfkF3nZRGa8qnckqAyWx2KkHhP5FBVSGJ9q
YHVSCSe1oytp7rX2YSw1bdeNKdXG/lp4hrNKRUvyv6jeFIqwTI5HtZxx8EW8mUOc
xYsWheOTlv1W3+rDdgVjBQwZK/g5nauvB1wk7rL+2A/HWjEgyQEoa9xfWDKS6kCc
8N9Ne8lXIBJrt7WDIyZ5OHXvbiFVex7zHMnxX/qWPLg0fV67cyMKhgLapwJcZovJ
KN/lUJhWWKWsUSe64sNfUdTB1MYI7OuxTLok4W4rYdwHTw3OLsLF0gzf3sNcSQFo
vCBMlCEH9kWtCZcOL0YDR05QL20Cc/rHworH2BnyeyA5qvxb3KF6Mt0xcsFb2hqs
N4J/8t3uG6KYanEnndgfvEL50E3UD4t/cgwCvIa4AI+9VzIIzOWHqDAa0D/7nNrT
LdfJyqC9w5XI5oFFUTmfZMqdMEp0XNC6SDHskvw9nc89hmUt8uiOj0583sKZU0Xn
uAhHNozishrq7NvhfizoL6iZwcxKbNbrD6iKipqhEoBkn/rGUDreURS6F+sAXCkT
aCTBXDayKDuYF/QNguYAF74O/Qr1LqGP3qmW1Q3nYufanKqjHt2BHLrwOq/dE9Zl
fxU0Swj5aaIqc26zqr0eE5/Cf9Qbcs37VlL4li1tElx0UGLmlUOvmEuc28P2vhuM
4cvQm8lZHA8BBCAf3YBsz5lWliddXqRDjkNG4tkuLQ0t96BEu7cQ4oXx3ug3U3r9
RgNwrYr5nRib9uafwWcMvZRudF3bNhZsjHEE+4VA7NBFXk5wd0pUh3cdp0JGv9yC
uwXBIoDtRJquS3UiGQNId5w6vE+3OOJ7Vd0/lDVNhqaP9Hctw5JGgBiomqvMm/YX
Yqfw6tS1whZ8JAJCHqdq2wCIRAh34rT7hOzp7KlnT7WPRJ/hInRLGxkbq8U/5QEH
eJSXBoovg6ZnwGEPaKBeH9wVBTgBNPFfE+V6byNRUvsv77TAmjQyJU42YvH2vrKW
RVTkAnSjfmK57fCtouZ50Ze8+zpfFLsdWiYsBM8ZY2kyOhmDDk42pC0PRDU9jiqF
JV+UR1K4gLQI/s7NXaZ6XOOg1aU0rdgR4tBOt8hDocDOJMKcYiQSucCkB6lUAdgR
grplvekWy67xK4TbxHt8dkK6JZ3IR+F2I4uvo2zlCq8LcL7ynNLMIKvEdV7AUqvn
xVZj61zxIMsVdlMqUUOX05ceknVRWRclipK89N34e2S+jLphyi8nXT7nU/g1/KWw
6SjiK1sqKGcCofaIVroM3tSehTbGNmGM6zbD+/ntp+NU0ffG67pcxCvprFRWBuwt
4nzbLPdqzlpOKzhtLvCKSnL/JB2vC5gev+ydLJoU08TgnxR+Bt8g5Pn1srE0yOBs
5VgM4jpsNYCCaP3cSQAUN9mqwEMPhJVM/1pS448+ki+QMkNVQzGFRtLvfYG7K0g4
TT7TsxCfvFJ0mxHoejfMKDV+Uz4nM2YzyZkuqzMGGVchyjiReJO3MpGNTqs+1Jc4
LqPiYYne+g3b/zjuNkQdLK+6r2bIGzVCyW/J/Dz0Fa3YPcGu2yYhPUGlaXsBCaat
gtlsZR7/nMqH+Aoy+88TTSdCpAEDp8LuUb97pXDyEkHu870Q/nsd93oDvBwtPMjf
8zft5f53NK55qPeu4rhzmy45+cQjVZ70Xh3jBbyWReLlOYCc6JzIP3Nx5IodEWUp
TGJr1nMzB+b+hcoQLTwqHjrCxhOD0zXywpvGqcC6pRjxYyEy0fjzTKWSxMRRqMy8
gN+NG2jphGAE+qTHW1d865pTsvrv9Fgh4SZY86Wa852VVnC1poiT9RUDMKu5ojMY
ZpQ03kvsu+6QH8YUwjFK3WVR2m+n3jpwz8NJqyZB4RbRdbl2HnE0CPFeSNdZjDxC
WxobkcrwCrF4dxahVzcpjUHz/NK6HfCG5L98VJFEHKLiQ+xDDPxCWXS9OXX3rshM
xu1GBcZhlklh9HerBK0HeWHlNK9apXouAOByvZ2YCDbrUXKKThUFagL0nUD7xHM+
7fVdzZPrD3OZdL8QZIiqpCPCEwb5XwBnRtGrdacfB7nfRNA8JuiIk5+auTxHErrp
A8u0XIRED/uBQTjTFdlmMfm+L5tZ/TmfeyfQ7Cvf48Yxab7TBt/6B6MqO6LDdzWE
HLnwggYGWgMdFxm9ORVAQoKQnDc3YkYJ/FwRX/sIVbBhGBwLh3T3iEvoGMF6wBQu
/VkMsAdGWeRgW/u+xjeyX/XacF093dDp/WB6iHowqYDazo+lndUdp7sdC2NqvDIh
JIuGHp2rcdrWPQZ2SUxcWJCetcMgxUG7G2QRXN6k5x2D6hI9KxhCqXcugVyzyBlM
q1YfQEaI5YHkJPn0hGwJTEolKRvFee60R5g/mKPI7SElSrK3+D9qCEpMZ9fEFmqa
6ErM6kkVh7LCph4cElC9247o3EAR1Z3BdD5kIcvKa1ZWaUJ48NnliJjzV6xbphxd
bSP0BMLCRGn0ghgXnB3MzgbocpRO4dkqGZjXtJWh8wStLGTtVRcKtrIMUbZugx+A
hMn1QerraOTSyikPTngsuPPafxpqb9FxCyfpHfx5Ke0LA8RhgmRQCuzGNIDPWzDG
zWjkNlDz1/e3bCZTYRnGpck8HmAtACXBcAozdTh6Tc+TqZUzUTJ+KSJwq92rczpN
D6rAPSpKZuov0skfwDwpsIjkJSzomFQ1z+ho5Bvbz4XTPEbsap/uTP+I6rLuSMO7
trHkkwSxBPL0+fmPvIGiCaPJVkaP6/MeSZYi7SSyuasvMlNe8pWDKkLirQbPM1xo
rQdmKHDrnAklGSdGAUYkuojVzDAK5RfJt8ggF0yPOhT3g1+fLHGY/8H9JxrOQEO6
BPxf1pJ+4GFHf0TpJ7dHQ+DxU3qLmGudHdf33xryZejEdVe2qORjg8NZ0la7lXQU
Cu6MumBZs4iYWJjQgttT8iQgrt/zwz7hfHVSP/iWWO3ZdeRqjuovrTowpOyojIAQ
ly/FLk7J8+k+0//T0/HSTEi2AGY6vndydH8ZCkjYWDy86GWrOaUzDx4h+ggeSBEW
s5p8AZue0w2rhcOhslP8efR9gLyYOuQHBY5vBifcwmrQQmceem3lrSkZHnNbhZWN
XUw7PukmZkqPy7hBcQFxlj6F/oOvAjiF6iJgjJI4A78UMiVTO8nPlCVpM3xf6ilk
4xKgWGeSoztReKTICCmtB9r5De9eJBqaOX3pAdFTsQLqlsAkBrogH7LMk6HDI+oM
8ZHNW/9VVLba5SAIznXZHeMgCb8YvZZh+Qc2m+4AW80ZkCKsruy/wfkJBCgRI9ev
EYxIcueumhgyByROOY2Bil4IcGJR9iyv+cHdQ802IypplNQTWUs68y29fZhl1b1b
fBctq2eYr7keUuBULmI/VVHlDEn/KWao2Mfh2XZewLCxjhLQZLFSl+hhyjM1Jp9I
sy5Ks7gwfKmTyHXg50z+rgyQLPUb8Ndikw+6KtGS1eHtQTIsNxHar1iPol4KKrnz
P7ridamfh5pyEfdSlP2f1PUp42F2PIJSE18Th6Mnp8dk9HlngaLF2iKi25cehnd2
t5zFu5zzek044agIcqPHJBLO35uC7hKhHxoooP5phu7WtZXJ0xAi+AzHdGdWtdL3
BeXO/4XXMJX11xsxz7ZFyWL89dFSUojH5i9X7++c2uByMFbKGQ62fx7nnCroN6nT
h27ne+Q3d1BYWiHPfR+lz9SwDVDD9gT1IWnj3miX+hOJg5yFtrZCvjzGKKeDQutC
bEXmWCmDEz6uDwk0ePIZvPG2PfzyBZyZmucP6ePjkL8qQORW5/pmp+Zqp1AxvR46
R9eEwmyQKUiaul2w+h55f+MAOtxW5X1mWz4bo0VXkw5j3ceJqzr55E1JwjqSfvN9
4AxeLnCzDilFAcAS6PzWR5Imw1hRnOvy6dOeknUGB0ay/6emdI5nVTkhr6plMFqR
Lfh6s8j8YY5mWF80VH5jP6u8TZchCtCC9rgzpWT207Uknz/x2EytMVo4vMmupXv9
NP7A8aeujE8ppWqE+lc7e1+vGVK6cqdMoR5DCK49ZnklZYOO8kvs/kJfTymx+c5I
9zq+t3/hdYxX0kLX0+rbx3iRriFs3DtjlS8bjh2qme9Zqd/LDusRoOEpDaMiIJoF
2MAxjjUgP1q84uw8gTnQr0h47PF1aUbOk41J6qWMbebSBmMcNDpdjBAnV7ChzzmL
0bdOCFge2zI56P++6BQiF7A1v4StUdJMJNOlPt1f7PLmXcnPsZxjjtvJmQDrKevQ
UER1wGwsPXczh/SDqKaE0qluA8SPm3158o6TEtK0dcrJSqrOyExqtatET7YbRFoh
WLLEy9dssZPwLtFYCzlUScaB1RPmsnio4bAcDCkOODpHgVHTXh/q0TxDS5VjnMOU
TaOMwwWbiQnE0XbtW7ZgGM1Vd7oq1hItSJZq++MoZ5Xxw4RiSNFDXPMsZzIYhtxq
V19Pri5kp1h8JS94ncWNeTFC0c3rsInLCGUwlh1YwU7FbY6XAOEDx5ffPEuWaNJz
0F29kC2RwT2nsqxM3fzEuVe1IFsSXCZXMOHNzOVuMV9UZCG1Xc4XFr9bvXq/V6ZZ
/FgMR83dUs94Wc06YBDfyMejT3LJ5KjSN/Jqh8pUwLT/AL3MWlftBATtpAw081wO
4+L9m8+/mXIfZvJKNOjtwHHbWLRz4XeeEHAw/eOIvqCPY2yOKcE7jX1b5GYg3PEM
g1cm5eLJEHvQBhdQev8ynACmD6TvET4vT82t2SRlhn5gt7mv9Rn0bBDgq/44PcBl
2yMcbrcjOLj6SRq4S6Gnlspt+VSPgsQMhgDRVXQRdhJdUzY89rlmDW0WJT+HAakc
Mgy6bRIg663InvVYNAE4sjB9kxoJMpXU491p0+aeIbYqVepDByoBfIOK2gSeHHKV
QziSevgDUFyQukGLSJaNQ0fkOXxsnpNxo5Ocj10yXyQN1iqleslwNC9zWOHMJfVr
UcE0Co9UvQaizCONPVflfKaIz0D13ktozMws3XtndbopiOcoKt6ZCa7UUkRDqsGY
1VjH9b4DrljKzgHugEYwLp+BwDWZMSdpYW6uRaU35o3m7QzMFrM0nE16OLhBbFoG
+YqjWsOGCl9OdCgRqqcPui/eaLViOr9nlvhDyAd8OOcele4Ra8siGgQDHx97fvws
ZIXe0P+I0qmRz8h2fSiVp/SkqqmewAg6zbfK6n6Z6vd97Dvk5brITV9CFELtceZr
11Tz+2D9XgQE/L2bT0HbFD7l48VRmmTH4EU5fSdKSC2OszAa6m5eNZ1b1xfAov9r
aK0Rq40awDBRv7TInAKUplqbGSJTUHV6WeIbgmrwCO1z6yjW/IQRG/f+RACoawjc
baCNsRLSCMk2ockRtJf4EkOpCGHpUbZVs7rbOccPX/JQLRSz1krmU4gWD85Z9S/g
OOqpHIcgpCp2onnlMmZfyVUGWYTfwEu6EEW+zJ6UbHV6NINTIggnFG6YhIyrp+KQ
ZbCnZfayR9hMsn7BQCa30tYABBMPjsVeOkgOrG9D1pRYtayPxSAN+nx3rxSjBgkS
glAzj2gUhtKAuHlur9PTeFrojxjWkKez+5NtpjizJ2nKkRoRYkH+1P7POdzgHuKi
gndVp/HG7TnTxswory/IlkBGQYRSivgY+FIRbv9TtyKrlXzXhVOYzMsPYvkyma+Z
Q1X/i/YKQGN6raz+0E+qRXniUuLnp2MJbu7qH0wu6gEubpQSKCLNkMTJATr3cpze
2oRBkKv7fH75dTHQEgulf1PFqZN4IV5IE4N2JMW8d5KJQuMf7QbZ+n95X7eZFCfj
FBCqc2pn5DnBlf6XsqWM+gVzFI9QrSbR33TxopVBPW2vAa+EU7cv0gkK3J2uTHbk
JUccCPEapLYAh7Ijw2TL55FQRHIflXSumTdW/Nm14i7ERs0uPp2T0jE/hXRPjNT8
ySNZ37soEZI7sAWtJUyktJ2izTZZ9bq3sKMnG4B4sbxNhduNjoImmC9f7BRXPEOU
cUXHNe5q+BcBjULPZ3f/0hDoZ099LxifFXZHVWTzrBIHRb6HGbzxn0pMjN9pWp+J
0VTcePQyajTph0gLKH/L4G48OiabLcaiwTiWVAdQzo8cgZHzIrAL3/o20/CXbceD
Wom1X1VFhbCi1tDOweGjWF7ZgYRe4OaL1+RdBzGEHrH5et6qiSMijtfxnlP6uG58
WQEj4H8E4gtqumQIapSg9SFcTkQ1A4tsinl+lxTz+mM+El8/s9xjvLoKLohdTCh/
G/BD3vmdiwVZkxvP4ccY9kV1goLSdvJdxCdTtkxUhvhFlBqNahV8eLmiajieGRNH
RAd6XZ4NHPpOk5ku/Y+FBKMkrDeXDvjtnai0+glmm2ThVgYaXjpBILMBoHoMxk/U
sEsavUEzm0VydOsb5tlUMCNM5KJJlNqbitgrAO8Ftbh3YDLzJIqNvz6BNeTu5Tz7
JTXEd31S0C2TvSxkpM6C66Qh32I5+FLcWyWjzya4ir55t7Euz2FHczwcG6MW2Esk
LyZh23OsWhlw0NerRUIfYQ4z3nN9Fu0i5nQZy+SadpiolCXaDjYYG9NLrBTeh72B
WKEZkz7L89O7i4kEHuxJZAKGdhKxGHx9rjKbRAHMHdGXuI4iwNO3TejEBOo8NIMg
HpZSQFwhzK18Zl9g7IGl2I2mzAY7/88KcQvLSzCfnSu2yVl4voUOw6xLS1ho1pgs
3Ldf4MsTuAEB5H20XQz3MmIR5UPUxFF2ynK/l6pJgTyztywig6jY2MDWaUrlbmQx
8Lxo+38wrv3IFENs1C19WY1yhCORViZPDHlagI41Uh6+7Ivg9NY+Y14IawparEK9
iugv7guP4klGI58pJ22vessHQvWC+b70ULYPfFoxPNIFZRXOHwBCwuHmZVja4iRC
qWL83b/yh7XVjsXmz08ipV73DWVBhbanwgmkXU4BJs9UiDA5DlVWa4TfiDmUdDFL
2x73HcBkc1f0M0HGyv0xRvK1/wz9ayOCx5XYcbLe/hhnhwxY8mxLx3y5NKpHutDR
HUh94WUhL8B1pVM0HtV2T4X2ay8ezXLjflaG1DyQtaSYOPlOXqV7IsgyZkNR8uFe
kQ3NpG6Xr+3Vb+6Fb3N2hSDXpPNhj8vrOmXjuUY+y+lowySuN0EgOk5n0nqOjZsZ
MOIefb8gFCPR9PcVPakJRNdlqJtbpewCD4s6CZudXrghthrLFKrTKbljd8UcvSDs
22CP7BoVMh5fVOb1dpE6PHRVZCwOJhwERn2d8RwRLAVVFDWntoGmsWT/zYsaCxT1
ZRru/rurqpBcfFOcqzFWfSXerK+VDpThfu8x6BDU12x3E98JHYINuYsb75vdlxiP
K/havebRrF7FUPKJ5YIT/b8gXEGECmgVa7mYKJKRF2Jjdf+RrRrtSG+YOr2NUNW3
+ysMV+lRFozOwvUOcSe8fHLIrPSfUP77SVSM46HiNecJVK79GZFDLMC3VIe9D18c
aQTelYYEl9oHhl4sPv9ydP3JPV1TM1//vE9KRfvE7y2GQSu7q5aKtgg8C4m4FfcI
EXCu0rfitbPHRMU3Suc0HGGBtopgn13dnjU1RLBFbQUGens1oLKB/vJhC+ljg77B
LghdaJWodZRAKpU/lIvp6bv877dGFjecpw7qGuRRFP9MAZFFjeMMleXfssiu1yLn
cgxpPF/G/Qvznc07H9cpFrD1cMwgyzz5FUX69vLZvexXXqU3k7cXhvQKMwbfnmnY
r9tSnszkMirAEbbN4VXWycSa0nh4pNmnsCWZqW8mA3/70pMVtWCV4dS2YXxHcNJC
SmNyfp/blNntAtIKpoUgHIMtRJUbNKPvnSuRfnq0MGpAPmEip3Qr/rjBZoJkmazZ
q3RRsefgF+gLkILdTt5IDAnuttVEiUIWAqB+8AtbOFh3OYHYukqvt2VceLpR8Xpp
bSuUy9qJKriXPUFRQsLCx9AQ27fwzc2Lkhry3fwjxhq7WgtinKoafK7U3ZiDnJig
ySaHfPuhHv3ObF7PvixPCVHCw9hhM8LnWymwLKH6LdRId/qlRLYfpdbF5XxrYPt8
YOMukzeDGHZJe2L2g4PLpB713YwP2gkMyJDhy4Vir5nR9SqSxwnPdr8Uq0vrZ6H3
EzB9M6eOoAA0KWaDaebN3ojVv2coRr6dK758Wa/CGKYolaFP2oBguX0FJlpk7rey
o2GjJvrhFXy6TsVx2WkGNEVEz/+FvpKvX+O/Yps1wQZAUdDsOqBd9IGZwnQEoxdT
AjArNCJX2KmpIRuiVBKs1AChifjP7iflAa+6YOppBvCFd/pyWFv2XoiCgrLYeD/y
VRfukJX026vvbhCFe6PYtKZ+Z32G5kIISIfaMkCisTqKe+S4L/Hum9ixR9aGqcnF
jhDUyU+NY2374hM1WGiznwRObl1bwBQRKE08+MOYErxjcet24uTuEgQP6ZnBFcjF
866yPFB/Vu/rcWY9anQMvN4FLVK1LKdYBL9r4avNvIPa04iHfYm5g9brfLsqlgCh
25oaaLpJj4gvYM//dzhqWxsLSl13bvcFPFfoH+v3jFPF3o561QsshEFbJ3ufPWVh
KEOvpzj4l3jgRspz7qjdgOlxvLDqOcUeeQ1w+CD7Evgb0tgGhVydTb4/3Vs7eJ8I
KQL46SrWnpe3z/25/jNk//1itOmloUSLrE3MTufnD2Ew0HD5wuP+hiKiQ+w3+fZQ
Trm80VuhaapUIErkA7puan2AnAomzuITmI36tC1rCQzz4COQL0nPgCiaNGimKh/8
d4mxj1q/MqQCNFKSlyLaXXyVLCYCH8NjSXPzvYlt2JBnS+spPyMSK7oIVxSo5Sjt
mL2H9op2gjpY/BG1DjU7oJoyKAEZ4Sj0YBWyqysw2Sy1UMLxlkDSfIwrOJGDkgt7
sRIje8sUocTYU4HPUKeGg7N+RKVYMFqm7CZ+a9Bg/N7WKX2zJfcXm6EMktVkZms3
GFhjMbehpTsRjq46p4cRdgYqNhP+CSEMmj4XLG0pYtfnyLZVVZKkPp5CAL9Jc/xK
DXhJEERto0DWWZZ9uOooWQ9H3IGVwuk0bUMUuP37QFRV2g1dL3EmYVDTjj6INoBC
WceM3YnAYjDP7gXsFos3XobYGWqaTzP/fab2hdpkMh7NFRzeo/V1bYn2X0DZPhba
uJ3EL9kGNu+JNOli6i+N0XxjDWrCQW9LMfNXSh6/e6H6V8wO5mfuiax+TU8AQuBw
ptAIVu5yKB5U6y4APf3gb7FzgtQ4PDYUE9XMZD+VNHr3YeUJdXcMTNOU/hwnqFmA
S9Ao4dfCXhKEFFQaU8gpoFSWjBCrApSbeVvLW9cXh4nTHdcB5sL4cB3SyYz+HPEg
57VHQ7oGkG/R9pQ3RSU1apxdqns+8lRzATQUi/JyK2Vg9L1qGGpuxQalVAX5949b
vmpLGPBnU64z/ArDwZW+HCCq+LYNiSsfDmeOXLfzWR8SAps6Mtsdn0DQfhk5V1ir
q4CP9T5Bi2tLpRZ//+DzLxdYoI5ArK7tJCv7p/94UFnLnxRARVkcDgCX74VDQ0l0
T9hzYRTqkZs04npBWn4igMkQb2uxz8hIyg04nPNBFfDCZrY8kM7bNG+9b1iHmX5d
AO8PraWYKsC7LwfRUx4NIyXULpdb/2DzvlEfYe37kOS3pj+QDA7EKLZhBZTigSYN
G8IVG3xJ4I/OXd3107fUDsuTd2TxfQhrf4ZylroJA4mrIqgmcA0Qjcpq4UyU15Nu
CxLDvP2ApyQwXxSFqKqAQEge1oVmJ2BgFmEBuN4csVDj0WUK2I7vn5+Jc6HjH6l1
4CxngZmR+7YaT5ATqdE52x+MjUJWVZAWkXUyrnDDuQaGHG3D4wPcCq5G9CggRIhf
ntAL01TfU9slnZVZzb6iVOwQD4UlV9z3yJlL71UmPEN8N12tVvcHWN/1kmFg787w
umo6mNA4bl4Sje5fxtaQHnGZmyAmTOZ1X16B4AU/0rMsqPSEGAcSgz868rBhZm1B
tsSQv7oREq4t0ZDekCtUV4x1WVKOkxj3yONbQcx8C/FuBjbpkJOr1epLnYEoITHv
iJw+QsUydORi76oLJVXzYQEiG9O5EedwsCriP7upe2Qa7WRyI45iHIavCR4G7DD3
AfARp2pUnWWJC4werILTVSAPPOMC9qGgQXjPVEEPkOC620DWu4VG6mSIhB99TlaN
C+a8arwQifpFPEmRdJgtGL0loku7JmjqWzyUSFponnF8byQ4GiLvmksvusNWH4jE
VbeGTdYFXXj14RwX9cdRHUrQeWpfMliTokSgDBvVcrnaAFB/x9B7DWQwcndQnuRj
JmDg0ye9K2u/jPjbrand2lCzAzAlfOZgH6+IYLDb/8yfLN/s+FdFf6mGfD2hS3od
TcHCxbxkbMx19xVcHJpC+BjkQ7nJI5Brle1nNxWIVP/ln2Yn/BZQEWciGE5fyWZy
og9kr0D31kgIS74T5s6uiiTHn2KZh7xAh7OmMGVhZfeuDapg/4cXqF3nPH/UPus8
43vnHEfKZm7Q0huL60TfSyGnM4cx5mYjzYuWC3SsFjjeijVO6xr9/MdeqjFlgTFn
bBU/ptD8lMyKa9+mNFcEGQE4K0Lxo9E6k5ifP2f4592Qrr7RZLFpjBH8g/6pzzTU
+vf8hQbRdDdw9Mm1yzy2QA5C3cqGm6HnrmkhhmXCFNzs7qVaCQ14zl1J+avQsQSU
ShhBQuKq9pPgDeQkgrVFiEAWT8YV2Fcxo0de8kjaDkHOCgCAjjAi0KMQBURiWGdR
QoAe7RxXk6k+brTF3fowYdTq61SRxhetV6YWj8XDV5Cv8FeOJytbkXpZ3Xm2SwJs
QUlQ3HXTRMg0JVZqiAP3D6wZzLNFbtR8Ch+BMnbrJb5hH2EpKM7yqmUEqhsoDbXV
jd1Zojuv+hwbvLjdlYLCHPEcP9HBGMgp+6NVpj6WTX+7NPGdHXQ/Qov3yO0EreUU
pBUqdECCkL4xJZHrj7iw7iyXY0zdf5i7U2Ai/Vu5NWeau1/i3CWrUZfdUj4OIp7e
ITAU0xMzeohHY/cEuE6jy9dhhVSaPgreyHdYfW4kAtbKBZIsRhJTeyMW8+lGz+p1
MXaWvMqVQWyZFIvFnPIVB5yZxogEhzjjJj2RCQMUhrcGAFf2kDqP+r0rqZi8KUPK
HSRr6vsZUpzx3ruyLheQn5El3wUXFLUzzmctgxhN/jcgXubylNl6mafy9PClCpbj
OIe3juvGomH5Slo+kFY5w+Wp6gw9OU4mQ37FI0hlG2JH1vAXAWMZxUyMO/V1RoGo
/yLLcxPJnAlmP4ACl7jud8/N+yJKAzT0IfZZ0H7gtXvkdupYr68qgQYdeLan8j6C
+oZlNAvk33jBDwI4ghXsXl6vz5B7EO92b0E/liXCv4ffR18Qfxv/r8Wku/YCquF4
8WcyYMczkXwmFlMEELbHXuAnwEAfbErZUcFgOLFudpQuhgSESvMXLFi6ZcKNXT1L
KjZcnUDwrKiK8nitJcrIxP5ISlvefMpZD6Fh+tj5GDSHAnMSsVt2QaK+dy1mhAkr
AK+wx66bcTlm9E+ceI1ESg58P1kguBzTpmGCZalbiaj6PqegS/QThtTvsXYjmFgx
gjOPmxkdoZQFZYBCzwtS6NGTUTRf2Xc/gtjO1yPsTxf8zm0B4UFj+XKEq+wnO7Am
jedrnHAE32UjQYujafP1IRtX+qK37gYiDrIzZbYfbKJeA6QLKVmgVnPnbuULkvUi
W7EvIZKEdbnMnaK/oumuE+UtVUL01IuFJz7ko+1AEIBbZvZnvItE2WHFkTv91tHr
jtmEI12eBMnTgwxdjcifuno2Non7/TV7j2Ei8GsH6gdzWz/HY+IiD1UeoUvyYbB4
4yFl4XAA8u3xLi5AlvUPfWThbSQ0gHqGLHIl0we77rs8jo7JWqddNEJtBh2AW4Ur
2yVTY7OQehl4EHIGz2XqXfRBcLFHuh5S+0DeGSdR6Y6FYMUkHJ4Z6kx8vtMYOS4O
lA8emIuosBVlD0ryJD+6tFAzvx7Imn5WbRMYAa3J0syravzBJF1Jt7KR1/JTMnPz
+eqEyXWZmX1tgt9cyjNvEQhJC2mQd0dcNU5VY6rq2Wjy1vRUb/wGv1DdhxMigpI/
pKr+HMDlWrk3x0SBNvWBvainCfDawFB0YRCwFUBZEb4KGQFQsPhPOccvzcmg8aGF
gcPmBrPRNqE84uYea5VkF5y4xHPyVtXhEwTNzOV5+LDLFZvPF8R0mIMgZKnxS+AF
LlZlLLbSnUAscqZyBco4p5iDFYJDPgi92DLceAlN2ekBkMaazmR/Qz22yc52zlfC
K9ysHEuxW54g7TQOKO2BmuDTGGdnSYiA5CbxHs3ch2+nPHKOjv3WBOe+4FQ8Nlbw
X03P0c3PKoCIUlngFJVsEw8j7qqa5tdRAaqrnZ5QZKvi+4CErfKcjdaRjvUlWq3E
nYmg3LaInE+NwFmYg4x5byQ7/usf1jjteEH6K+wMh/3EAL10sN8jneCJebi6s/5d
5quwd2Pz84LVOpBC4cMhr9tmGfzOlSKupQyLXcTr7Y0nmEPv7sYTjmUnb5VMhIff
HRybDc8Mj59aGNixc45HgeyqfpGXSW4D+B0MVrmRfcAAC4YqvE5XG7O5KzEseF6r
WUJeI7iNQVoyQFkafjHXVF49OmEDvc8TNtRcYv0GrSeMPOEcScsv8JCzWcqwXEcU
kZY+j8tyikZgWN0LB90ptLCp7cj+52P6o45qDEeZKWXjvASn4IKx3/k3fb9pggoJ
1A9P5oAr0naS9JSCxe1ek5vb3je3YvnP1Xa/2Q2biqzKsOz8RtJGBcBU1KMZ2QVj
RTDuStM0gVyfWQS+sTzasouIU6SU+lugZMBWXLuWWSFreAZdtvELuVlExchFjtTF
DVWzhJ8pQdLWoUqyXJ9DiuXPSXIkExy74zQo87X6iNxyJw+39Koydx4O4OsBdr2Z
IYU6V1RfQ0T5VhmlNEeWS6EDHzUYLTXFWcl+hJ1ij5wIwY3RAtcogTaTrIcwXyMO
25+URWlk4PLqgq8HZNJ71wicqQ6oPhTArNqeCu6AEEN5479Q1X3o0QeUDCmXnulO
HU4I1BLkCqH5sf55+5lg87OmXjt2CsfLD5sfMFOecXR6i6jOz3h0puaHWlAaXy3k
4AMW2XKAD8a8pcBkK73fnXdMCkkBNyeyJLYqLc3/2mhO4qBvy6vWykBdoDnAvAQP
sbwB9zQgowNqvnQ33L6fSCSdztPJb5pbvJl8Fag3GNaK2N3FUsn6KIAY97ClUJOO
ZwL5m1E+S6EMk/iDpsgYlwBR0NpEcUCvm+8k7v7bD/I4VxeLbcSLXQrTIsN8gs4f
gcQcCrAuZStf5seCXgvgpAjaRFrH1JJSFHTO+NNG/xDUXjnHOrWC3GaX+VPBjRh0
HK/mxjpxkUu/o5PYWlxJNfZoV5GJq9yY/W5V6X+B5HB0Hr0uxOW7uDjD05lor3WW
ycTHUGKqxz+SI4I1S2se/V9kXnUZ8nRQYD0dPFPcuMlXml8Eet2T82jWdfAf9x2u
XNIjJWaRlU/9GO4eNPlXEGjNTjza6nK/nimiX59wXmdl+yZWr+4mnKBPDbf/Xafu
Oe3CNe7w23SzvmQdnrtGSd4+tO4uYWYWAzV8czWbViYfeeSpZPQ/B/onqLIItYHJ
suSV9aOB8ks1J/8beYaHFx1Pb4C+mFDaI3L0WPLpB4fOvm0HcqDYJJIMWXqw7RR8
JqZiNsLm2sqTr3ZGnYLwnUByB38l3gsl/gguzdCf6g3O3nBB5abmPNB8isVJ6fI8
D35Mf+tfdpftyEB1K36JHkH/4Q/8kNRGjT6QwZjI5t0/zumoaAAW6FKMhvQrsm/E
Z/f46wH/MxNs6XadrxTKk26AazrAlKXViegNHfCHrYY/2vy5aAAfHhIKArz/OEpL
gh0Fu9M+yiqf/hkgOO5emdily8ykm7Xb9k5z74cPD6300xDSIL4pD+hoT+fkKmM+
YQd3f9ZlvAQQHPU+99aSUiWPR9mLMGKLpNzyd0QFiEcAYmLMeH9p218iJ5iXv/aD
u4+cCWfG89yZfAqDXTqvnuiHVk3rxZlML7rr0gBGFdO4AA+n+PbXHiEeaXZ8Qw7Q
9bihKEQYajCUopi3wS7dmFofkNnGazvkpMaHobgIUj/8HSk+nEhzMIhpujDqORBq
CofK8c66YdXJG9y5MU4Du1meG+ZiVCasfO88F91WNdcwcAyufr0izvBYXLdfgEkM
aQPLgdAtTlATIqD3OnReK48yMVskig9wFfRfbQxZZGieov1xIeDzGbB7B2h1HWpy
DvFdhSsNtIotGC9A9k7/u2emJYq/UDc26JI3rxE1fwj9rp3uq2uzTxjXB3fLeWIc
dC+CnXpbf5KfUBVVSa8m7DEHpTWV6wn2TqufstHK4WPHTwZYo8h49bmeOMN6ypDw
phQxfT0NWFxrVcw0pf4yfXBcSJ1/YqjdPjyZK9JU6Jl+rx2xFU8Txe8twRmr71pL
8W62ioJoSirlKgVHn4lzYvhxobRZ43K1NSWnHCeAY4YD2slqv3evk/1/aqSWclv3
6+SN+iOYyAoGBWmZPkqyQm9kCFdB5/gJcs0YC0Tl5mntdCRSlfO/n/ds9z2Js5i+
GMuNxUgoyLBvoKnbsQPJndOkLhWzFCgfnURXX8pKOcOlLSvGEdgxkJMO5DFG1kyg
fre8eidFXhOyB7ygk9MkCUO1iFn4grEENfKbdcWor9qb8bBf/HiZ2qLxm8Pt8l5m
VxahuMq+R3oqGlpsrDXUtCPAnkAGGBukRJSsgK/ymlWwfS2N5Kl+1d+qVsD0J1Bq
JmnZ02P/oTOuBkwLV+oa2aaH2DLpkmdmuK9KpqqqEP2e47MSqm10beOo6KzLq/vw
spj+1U2UA22BIl8/dSB5dIFAiaNl9lKk+yj8csrnj21NbTklAVo+nIb3UshMLf86
/GNpgR7lAERTp0AwrIuUtGRyj9JrF8shjoZF/zoRRB1E/K7O/s6T8+XNo2FS6bnS
CgfFhjuCayUnQR9XevGQTaJO97EOwy0nkrR9WXn9+YOL/C+R3zOLpIjtvjrdQmhd
Q5Eu0d/l027VvkyCFQPUOes1zJsOVSUTkPx1Dy7ls/pl0svLcukmV+NR6jKjPDN4
a5j1loTqJCI4TtDCCbvP4Cg6pr/4lXbTkyNatvYaugKQcYaVzgI6xyyWAD1wSour
iWaqw7uGXqUecsXTds8CygXPk3yY1OUBhFDYO3hYNh2yeD/rUdmIx/MxX238TCMN
X06vVp39N0motZEwVL6unyCyTG/LASp6qTarIMTJ5T/wNUKFA/ifS5dLFIM9wFu4
Oep7SKwXdohbQRLLI1fMO8Qi3qs+NOcogvA+0IDc+f/GQ4XY5zWE9JR138Gd/O+N
6WzoXgLoKFXk7u8vapdoiXcX5hVYfgbGOrka+/qB8EKJh7kHSQJhkS/Ofxgolpm3
QXp7PrKVcCtRsesfi6XqtxSv+/Pf+pPDvFvUohLNk1/akmJ1vJcQcTwuJQ9SA2cW
RH9PV+YUzkgt2OagTp4XOmrNe+a8sCPdPChyzOq35I11h1Whw++REDI1OPaA/Int
hyVzx8eoWgnsbxqo0UXT2ceELeQGHSw8mACgzQaDxaU/GV5MuwoJXy10Ec5tKSec
WCg53KvyX3DykYQFkr82ehVYcsD8qRJLEE1uPGE1e7smuwN7pjnD13a0S1MN97l/
DXlLbKqr7KPDhVfgguLDPBnXe/P3F5HZBRR9tRmMsfL/DR9/KTaU3MmKpy53a3hp
b1C6U2wWa8ap+9K8TqOk8NYSJHnVw/pf7zRHUfBY/vv3H031U8A6jaNRkyXUBU+R
8LvOu2dOFSeeFZmN/fNF0Rs3RXcY4fuOQJxdWbNu9zIWH5OxK09ImYah6IXiuoar
zt4o5XPiaE0hXw9+UmQUJANtTqrCs+Jz9Dy8N5Rvuazeu7U831nEZCxPjQS2ghxl
5BmBCI3aCCLdrF/M5yCNiXggg9aLJ/EeyQ1KmR4XNVB2R4ChpmM77CMPq8oLKyT3
wJJCPToheMxzuUp4t+zNvf0xHrn2OwaDUia0M7/WAfBAInYgjMh9VfD51Cy8ZNW4
TiRMvV2Jsc0v1OsWcMLCiarf3hOD6z9ySLxbqw4QHVb9Sp/fNhfv+6r/etpki6tJ
LBM3TTkeKHIL3qWy2iQaMWroah5dRyoKaLIYzczsxHzR+pqrpYd+0Me5DU/LEMK6
xwyA2UbHmqKwWyIzjeCS2/6r7sf+TuMnakbOaZvx3tB6ULCVPlqvY6A+fpW4d/br
oOyZ+ZdJJai9fhKMe0yd6r/GnBMp0DNltqDpQnjzZAVy5iEXGeewTccu1N+p9UPZ
NDoQfmmKOn68Gaw9cvrr4RBDSpamg3RUwU0sIrIHP2Df6ALp7gRg/c4QMbXwE7hy
P6jPYk3uqae0jKXa3qII64/bF7VrwFrfYMM2vohCnTYq/U/+TuPbtcbekQyiT+sg
qthBm4uQ/upAtpGV9thgysIjvZeyuA7tUZ/x1JOpJ7BstRDJhUgcfvm8t+e59BzB
1azVxhu4RFXDvzjhwYmf9Giau4ri+MXcr5m1rLfSlPEwmvgg6oj7IjFh5qqRoPW+
fCwU2bC3u3PehDWIVW65hipHalBKpDG36Vqblj5XhtMLwDDRElGYbF01b4CF6tB2
hmqdjTiiDA+kY5nb5xwUSNK/+hOkWuurKd3QPE1O6KUZUWM1buo2MZtRAu9XCCH/
19mjBHHGsya8vlG+/FPEXz4ntVCHcpDuTggMZALN6/NxVT5ohNevHnmw51IgrvCU
yZ/SYaCDx7Vx0K70CenMMsoShhHvDCQGP+6W2bfSFbUZSdPj540wHdY2toQlEaVJ
wbzDZuYL5ZtI86pe515zqQfMTsEuTUK1e0RsQM6RREBpQGYAsZhj9zE3E4KrLlbA
qSbQxthSTGPIHBmydzBlBuMLB36Bmh1XIg5kApF+kPqFpSsZzYLWEloF3emsTYkt
rBtfe1odx6bwm73+PAtBjE8A5UM9LfovQImVzdcnxv3AnLYF7nGyR5KyJ7RdX3ih
x4IvhRPKikjPme1DNQILM47ung1cFN9NMLx1oJ5rUJtnZVzhPnxD6Fez7SpeKuLt
65IevGl9eOkISLT8TkyDf25RLhQavLRubOeMNSYV6sL3d5of/31H/goyT8XQKsCA
6zkSwXkztrcTne/h/JWBGQSOdYG1ud8YWXt0Ljdc1TUGVZIRiz9W1R15013XSLzv
VaLoo8ymTQt7nksTCWVLQ2yHG3KH5vdJ3QcbVTc10jpr7I20d0ZzE8hDEz5jCUm1
V76XnT7fEP8Pv10Qz+IlO3rMfkWQPi1AMhuu71zfTCw5VP27aGhTJzyDLsBl3zgO
IUOHwe5kEaOjibU/5Srs1KGgrMjoC1MKQcepSAYOJ36+EbzY3r/aMLeOE1uxDoZS
gVQ+cBdjddRdlq8oO4hNnGwcO+nDJRwYg6NURZImnQ2qptvAltDn3xvwSSTwxJLA
OJ8H7gwMo4fHp5w7ZBrEW/evcJclg1emjIAi0r/VU8eTyvXVBvyL0FbHGx8kwHRw
xwy0qR0xidP4Hdt8vdX/m3wOaFv18uVDvorSQ+R7eUfsts2Y8rXYQL6tvKyBWund
W/5OXZ4uZu1t3GAWSjgCJAABpP+86LpgqHncjZIY2K7b/kkCUpAJEKvryJXrH3rc
NB9MiwLkcEoJUr/IsO52dJtYBEYmRrm6cbnqMMXQj3OgZur3DOQeuzVR4zTlQsvv
oCo44ZzhhMS4N5o9Z3HyKJFPCECXs/s7Kc3mbFBbZgfthsnH3E4miwQgTbPrF+bc
mvgZYRvU4vxjPzpzJYvNO8ceSMmsFDsV7YWMV8SHV+8vJIBjXwfulla5IRDH6jRd
eZepCEvu6OdrsUClYvOHllhybNbwtPckAjMPEcFgXRZoYriCIMKtC1nU41YykS6f
fGzRRW9q5p3ICtMgFMuqyfQU7kUAS9nYJOaFQxRMoCqXGFfn5p9DKD7nzZOqNst9
nWFHh7sZLztpQN0dqKsBbKi8WNS6jAcn1Kf/+g0nTCkU1ru58KTgc0NKqUNNvAlC
PgLyxFlMds02+bMBrp8VY4nK2ble5mzui08b9UDLNwVhM/R/vBBJwox1af3Cwrc9
nSfyJ0QAQbpcrRFxeGwfCXp4chhYsoaGX7c8Fqokog/69dEvC47NTG6ItIIez0j7
DJy8tgJKWG5x2X1w8XwDzZgnwSiELzbHFVxO/8xep2zVZOf6BI6rJYmReowlKAYG
GBkVWCceTDA3P9l6dxPAaYW5CiqzyH4c3CcdGff6XzyHb9FwvbtLKDZsYn1SULc9
x7puvXsPiilkIH+yl+Y2Y/YTZ9xAJZz0G2LNMM5vu7ne/TddY31MWEvtqpgCjX48
7hUhAwl8cOLeAowz0HK6MpjPBf7s0kLheRjZOxThOubZhbFUK6ajqFsoHCE9wMSz
aoHuJd/DBO3kJW7nqiLJmeg8Y9sVgkMNWb86eSovwXG30EEzKs5HZzVvaAhw/Ea0
4n/uHNmBZvPnH6+OtkpuH5/lx9fOOIr6qrpCSS+keztM//MFgWm3jh80F5tP4iGs
8Dvm31Lm0Lzi+Oj0YrVqxfWj58BRDzSATqwyN2v5L06YiG97ARS3tEN2/QphrCZY
LiwDc7Jg0Y7dV2OWxqvdt4QhqFyGCioi3iGVWcK8cC3ciiTgGKwOl7O2h7j2Pj4Z
9CYXPoFp92L7zOUXtT/rMlm3ZTMnoUEG9Zmm9snbsmEI3XKnPvFuklK1ijSbHCo3
PHKtLSj0Vnc6GHNtMZ+IkyckHDh82YS5PZrXKHF4WcMSMztsoZz+uqyKe/vhnXas
Y+ROzZXdW6jRZOUEq15hHIGvhn8frtErDSLojm/M019yeAfSRhM9woqtc1Jrgpcu
2bPthb7/Lp3JYVnjLhGhZTGQwwdHZS4NDmQ27gy16U+H3smhju1K3jFjA4ZtDWgG
mA3ZbG+rIjYtmtZDMJyj9TFAN0L+0DiuIX3hmfTe23Dd211PDM6ECMPFScQh6QSB
oreqhr0a6baMIqlOWXkgHscQ35xizrBqvBn3OuHz58pcKe2MPGBZ9t9CRM3Cl3Zu
aHI+MWzJ7mB5N6vLmb+0UrfKhSD5SE1WsKIg5l5WxvnM1ysvALUd2zScLzmKB9Wi
/99RdQzjmi8N+9tnI6L+Hrh4iwpi9HXU4ckc7aNRjOO/VXVbEL99vHio3+v936nD
yWh21GkUawNZUKz3pOqxcqnBZ2Na54btorO7nSVE+GTWSW0l1DcIB8nwIvpWzfo2
GlYEKPZB7SEnV5PBKPU0kxoRRwXWcPCHT7JtvbZvabRzFUUIUBjEpKsHFWaVYWf1
AxRkDHK7TU/22hqNx+2T4Ozs1bz5cRt1Z2rrPQooxLYtDwXFMSGjRGRoyt8kzwUN
mfwurUCUrs0aA9LFH43W0fGz1KTe1XRsbqdiakNeHlsgjPNPMcv0c7gq1RlnWggI
kCrhOFM1W7gblQPQSNQyfy5elBTvRVvydA38fTfFzbfX+YIY2/Zi/AuaciCLX+PK
qrwvnSm4IbvkQcz0QVxkipTMLNLY7z9akWdE2SKrLvRQRyPndbD3JdnjILpWlrTe
jPFlp9/hPovMrO4uAiUJ3Iog5eYpLsEKd67gI044EO1kBjV5kxlsXqxo+HazHulL
YrTf0BaFYyrQzx5lcz7psWma7yvDcNa1TbvzsMTNrKshDWfdSdx0AiDpwqLawhHP
Sqa7cQA2kQoaUBMg83EBew7zIUaz8zDzP9daa/lIowgHOTK62MeM5MPT7L3uEeI4
8Id6bfoRPTa9Q4vnA51OYpaR8BnuXpoWe0sQ8sa56SbGj7igl3MczWESZv5eUCiz
cT3TpvmNxLA1/asj+hpMbmyYv2uqDg41V06gTfnPFiA1TQY6wmxdIFHNadCsRm7a
RDxsPHWs7QDZVY6CydqRWA50P6DoJiuvOc5FidNp5iia89sL9xn5BgBcZVt3Zgd4
0O/+8VV1jt7ZSgoMfpZQaqDXvS5zDQKFGsAjfUEMzLPFKpNl62US7XjUVArxQEdR
sH8LBckZwcLo5HAmPsnNSDyZwhr4k62nAPD5W4ThVTnnSokviMEGsOBd2XPIrr+T
I+Xf10gbvUgAsxCuIJrxEDWOJTN8TQ8P/7bvpxiLGQLYsx16HsgBuK4MIIySClw5
nq440XR0qvn2JIvFrGz9+vg9m6YXTRBCv2RIH1YD5FyJV/mdzgFSoBq9geiMjUJm
V+ooEq6A/HmFk+sMTkOhYQqtjWv91e4k2ILQXSsWxAgHfY7d7xxujyI0lxGqYiXJ
do92XivwH/H0dJY3Cw7xLbBu1xb0tTjoph/6kS/R0Z4gvOO0k9LWAuKnR4m54Y6w
wf6djyaiBBbP5iRxTnfqhChrIJ7wLNQzaBzQ+q6UJeD3Ja0Yhhkze7OfMnY5o7sG
opMXcAKzzrAimadYIa6FVkvn12CTqIzk+tfkJTHEfKyjhJ12IG7y5Rjoy9rlNs+7
yWVMh2lML/eww1G3uUYKhkWbq1qbuck6d7Wzq+ot23Y4FfRSR2i2mq5gcqmcnIjt
wPkwfpTOr0HGc+klvRmeKs/exy5xKvf0ihWiSE7Gar6DEjlYZkqNm8vN48bF8HT4
5P9Aa8IqG/7Ay6Vv5spVk/1z34ixi0LiG+ruB3hK0HQ1VS+G14S7IUeZ2AnJ3YFv
KRhdOo8H02fTmVTck8oVmgifOHOjz7H87cZhR6aWklDEfP/S2kaMl4CDJera7uc6
6jbdvPZrHJeBDMXfJ+SkX5n4YxRlfxIA4hfuoVuA/+5xJBm0me4K8a+jihxETZ6X
AbsLrJ21H7VdCBUR9pkYpAJ5ZvstUo8XrC7JfiPpXrtfheDeEcmu5yEzUyYGucrj
yCvaSl173jmauQZDdqkf959P7ioyRtigEJy1GnYLNmlbOXt/MSQmujglSzS8Ds+H
KuccrUSc4wwxwGDJ46omltvLQX9j7qR6voVcTttrveZeitRKARbGNBRyag4ZeEdw
9Sn8Ph4QhA5mCCN1ysoIonIbUZz6htjZdZ/Kgd6xjXrPS4YfgQdAJbA6S6OkMo8w
uF4/5ZTpyQqb0TSI00DcGKIMzsmRXoj5YRzW5UuPaCoVpjjcZGkybTMNkShYUCdo
uR0w1+UNDbNXzmMBicUhazAMIgf20PCyKS2s1txKpyk7w85wiO4GX54FI9/gwm3V
x8CPRvO10VFc5cBpFkBEI6kbWjdUJGKUsuszkwWLRNNJ7bv+34VRD9sUTJX02wBg
JPzC48bs/nTzT8TUbhrsmJE+5R9RGLePPsDYN32JMELBbyq1bSm44FVGNqujMsfh
E0UsfFw4xSzABsqqCHbUzDUZ4/AVymarS8CgK0UZXRTEv9snu0qphQgoGXaxV+L3
r/tCAOliuYulPuw7iDwSYlwgQ8xix8OaO3ZcuyJsmcTZJvzhROvmuOfQFQnTxmeT
y6kCauCQQRY4mKBOzaJDbW2CIGUbSnDo2EXJzMSNG708zhIiFxS12HDYmnihIkV0
7rwq7LRnmGpCoQv1/zwtBtluZjAP8rUXlMh04P9+pu6WHE6tjVHZy5rmd9KVxEZM
JPztfoEKB311NMnremfU90Hl8Cse479I+lRSFNMUHrBpfiAXRaoLS9kmXf2feaib
4Md0x9aF/IAGj3xO3YOKBZEObQcS1Q8cVG6gXuf+jbsqPzHwU22H66CrIqV1xehl
gf/fhskP3a6C6oKLaijtlC6oTGpQzSJxzvtPNxtFH5suJV4XW4oBYVcLTrds1uWS
vN8ohOwrPNboLOGOzZzk1FL/xrhk9ockqQwtWuoJUAgvHe8fVvglPQG3CKqzcyFU
6CoDezJvt+gVSvZj2XR7KvtRup945BTmNfegEuRMJifp3A8jkNaHXByqQqDivQhR
LQT7nxBWiR5lJqNXvlzdTxswm6AMcWM0bJ3s1+Z/q9eQpS13vxnXpz1QebLlUN8G
nYGc69uEXFFgK+dNOMU0t3aGCiJJkp+lXoDdEaMA/Y5y3wH6oCGIh6knBUcIIHuE
h+8TY5WQv8P0tQu0wAdA6snzmzGMTV+jLx4TMU562p0r10Dpjq98mmatqV9aEQSb
9Mg2GbIRfTnptklOxdVmYeED+eX4NBMHGGdf2JZa/7uwUjUlxczo6IqMMA1qzjkZ
t3SHewK6J9RjrWg9ss0kiTkdnuUGkOjsSPDvpygIO3PpB81u91PLiKwr7StQL86s
xqfNZSnboSOKHWxPiiOQgICx/wdleWu3x/HfSvWfjebv6K6tqc1pRxuNRlrX5Kyv
0PC0KrdZfqgckLbbGbrFtk2TJcBdokVjhYBxYd8EEf/TY0Tvndp3DjnNrQgpnuDG
R8xOXdd39c2MQVyjU/NBlFOUC2fL5mfZBv7IIgC8Wl8kRhpR8fRQzCpRCdGyZyYs
HLLutKBMnlec3PqXbvixRNgPZ1o5zCSveOH2jldfBN55Qnb9U6otpQMpnuXROe/7
pKRQ16J1D3SWzloSI6Dsid0jXO4H2MzTwIpfmP5H4hFq3ETcDLVPbHJjAKKU4bEb
t08DGA0kerc0DnO9Nb5PRnqN2JbXqpHxsbcXE1SX2EJJQbDk/ihu73hYQtz/3KPh
vIv6YCgNTVZW+s24QPSr78gAQkTdn+gOa5jbHhgm9AL2+tKtplhh0sM/9+LUprY1
SIdHfejgKfZoZyC9fe436JQdUKWEtL+5AuQ/oPPbGJBFlS7VJOBEPtYgBZpPfoup
YM+3TEIMb4WDv2mEqXoCkNDYKM42Hze5cY9H9+knvlURrbfKOCw9zcnEZZwhWpBQ
9jyIfHHW4WkT8scxLtW+z5p1A7/HCxvG90n+F6CPqcOvLqgKdEeaJ+86H0Skmg3U
yWBcaDyAlYv24auSdAslXByPPIiO9/I2EBFUGfJM0awvEG/nLVdcR1t+M2gOrZWK
7k+s581oVzLw+rzCD7K/z+qAs1ZihAaxagNzQ+nlp0jZxJjdOhzmIXdzIHRsXhYR
uQKfFkeMGNqQH3wu3EFwCHLJZ4+/c5oIfOdCKMnQHszqDr59A6eXwIz65ChDrnpI
e4eHdEIDL/7sZBd7mk4GFYHNjgY2FjhlefMEW5srhOPQCS03PjsygwS21V7qh84d
sUUGl2+5W2UQ/mitO98SdyErnbcBgYLbVsI+zzuZH7aV3+jYEx5IfOoQf2YJB/0Q
nID66ts+dDn4xB4crb3FdZFJQehKO8y84fxU1gv2KgGgUFXKycRKe3G/E2Zfl1ME
CnfHaGy9FRkgSlsE5126vR/WnLSXn9nf/ZtxWyj6aDW/BdwGRyzlk61u4jcwA19h
6CEkmUfPvPq4bZpRvLDSXkcCeHWvbY2oheY9AhlAPazcKJisD1+2JFPp+06Jz2lP
/B4dLbU01oi0rNKRS6c9l+wyT3X/tvWIJ4AtSk+x4OV9hU8QHHS/lvFYbfpWQDJR
OsjYfRyosOpsI7DoW6C5zuCVjB5wgcJxWcJ/1bibz/Vmp3eVoJG6FEAg0mJQHAbH
zFF3w8b3+OToySEgmlmrsDIqhaIimzKpHUp0Tud4bUJr+DDOZfwa9SRlZlHqRZSq
wpnBmKoBcZ9fj0iDpRAoevZvu6V5RscgOH0I/JDK/JTG4+xALapaY31zi4oT80KG
rVCR0DWydt2cYn7DX1vMjFbOboIFELqvui6naJf+mrmq97jUJ/9je1H+3ymRP12c
dDUmbuvdJqjOLcjeBpou4ci90bHnTMmsk15/XrGlNpnTskmUnrAiCGGZ6L8W/bQB
2Gh0bGmFbDr6sfpvI7uq92dqa8Mw43huiY3iIoJ2UD6VCKC7Ai1+r3lKn0f4WoRs
KpQLHLS4EDUu1xw6cBkgonVM7FxHx8Z8n1VwXCB+SQRHkqn6v1CsYvP3NC2JZYKA
XdrcUS2UlbiQrOP90FYf+WWnxHRxgOnDWPJmxS4aCfJ87qL0v4dYUxWJ/8mJXkxG
+76uv9MgEAJ++ewix4zeuzwnb/kDi/1tHTIn0+cllpOGbUQcTSIrpwel58F4OwPI
l2vQzaJgzHbd4YUcEHlMNRAWyVUpbV/nSZLwvWzBRqsHKfQwPPllR4tRBUH5mKKR
GBQvy9SSnsbKeiePJ9Mc4JX1eRdhSjkNMAHtH7XI18XZupbcM9wcEcpym0YyVIw8
uFXepzey4G0utTekdED15BGFjIdIDKSLmqJBXml3eL3S0/IGMUFnvmsnjYH9mNGV
qJIjzkqwyDxu44jECS6czGcDKU9Mp9E0G5jYZFpF4BozhJ7FEWTlOHxLnw1Ye3gu
zeMaa4FSMQc5X+N5l+9GvNsuTnHS6mXYAT1OU9Ln6At1LlaYitQLxZErK++XLZXv
zIwfjxCQ4iit/WJO358gEJvTgCwgfPpNcJXUtkvDD0zRNskrIlu7XMuPIRScX0mw
y+TAOWIzPWSo9Gguj5bx9WSaXeD+/Djcp5Au5d59uAlm+grCkTuckccs5m276SvW
96KKBN+JxT2NCgCe+NQfxMTuLvEFgw4pkThH6f88ijSCrpx5EROtcaQtUH1az8Nc
kr0+xnlJMV9ZXVcubpW43QE4QCyDNrusrUmb8jZ55mFPG7KuH0L7ELezCZImwDwt
CpPzw/lWGPSNFlyrNvOcXiFWAVPrhIFDADze0cgvz96E1HrrDxvNh/N1wpl8lr7B
0RwzewenObj6DZWqfdngopHIY2kJaaBxQmWgzeM7NxB00p1OEid2peY7T/ReBF80
NZFZaY/7cSEbiUMuHU+d8rpadLMeFtWw0+Nr9Vx6C+CGu4CcVaQlKdyFT/mdEbPF
t5m0Xn9XCgRggPBEki+xnLJvANKfXKV5MJE2NMXBf0M+aXXVLlI5744L1OmaBOL9
1s2vrw3mwLujXo1W94j1j7KwR9KzehowceMJoCd9/RQDQf8zSxfXiPmogBAHSwsW
9LrKnJC6dXjmhDRjdDVntbiVcYlyu1Ik9jf80mcRqSFbB3N4DrjYfCegjOQwCuWy
CzahqaCa6Ukv9EqHnLjCevGVkdOs3poJFyhULKJWiMa1P2K+vP14ho9WNhnxqVWM
+/G/O1ecAqKiHDmkytA1i1OKfrTJ0lW2OY0y9f1HJCfeUArHO0IVj//ImnErjU+f
9ZXzwoDaJUiyxnhjoDnX00PUSbfWVpl9aHxWzWTE8SJxD3juwHmi1SlyX6nyTZA4
4WMRvmnqvJdXcyPCWLJ4vyOnLdt5P8HXfMFy9Crmhgrf4AELJlffAHkRB3fVpYIL
mmIE2uDoFhVzR39eqIEeKY6g19DxRgJm2/K1fzfoTCzMgCYiyhLX4NrYmhV9qdZf
vNDmeJgvVrXH8yjMo5kWM/hJZUVgv9dXQxQVti7R8McsgbcrMS6rg2HWhYwNA1I1
yiNaULJELmy9F+XjX7LjgO68y8RslUlwUDvtnF+AFOntCgCixydqWGnrYZuCzYYV
NgSZ9Mr8kEcuwIUL1/gXXEvosqzou5pP7MwzLpMPWmXSgmt4eF2IukdXywfFK5m2
6a+xICegZ5500KPiIGknwnBCPiN5+qAbhhV5VufhXv2Zs6mulPDFUY6DD1Ore1gv
xUfzTTPWt2mpHpQubspJ9vZI+U9SHvy7r+zsIOTLKyRS3P1Ihf9idc/i8q0GRpFt
PW8cfuTIqYBe+Xs3oQYbntEcpjSittwekIzjJKDEo1z+cXKTY5dZeNdHjn0k9MH0
kzZKqcZfYlRod0v+igju/GD9wKmLY8yWn6tXmmit0o0vvedztxkKsPM+1O3JjMMs
IG17xx+zG+HeB0Fg3zfo2ESa2kdw217jEa7jRoO2oK7gNOI1NJCbRClOGR6FH/7H
bJ5ICoH9eZB79eKfoIKMqLW2Klbp/xCctgYPDvhwgRGpSLigZqlLYHL+LXwG44wu
JmL9ysUusFf+n6DGZ84Uuvy6ixZiFemIwhtgnjQJcfA6ZFoGckbg1blccAzNFSt7
Q54mKv5PCrv8YVwAkhyPlnGM4UltCH4tWlCSwjmE64618S3UBITNCwFYxJCW/BY/
RyvO5daZ/p9OM29bQA31S95DDEJ9v8p9G7tWltfra3/4du81DPum8AZdlbeo7sss
9eXUJBMuwqIIda1jM2KT/8+es2HiazJwsw/YlObSism8CIOgD4p5OMON+ORmqIiF
FCB69yhwNs39qi0zDYAuM/12OaBWUo0tOa1oOpry9tNhgMewBOFhe4P+I1YeHlcb
+2WMixDZcaK++++yjfrRftStRdRUFDG9gJPYNHB6rLAfRF1mjHLx3R0vIn6qXeV5
hfpS0LSw4Glzp5C3npM0pa4c0AyKgHIzg8aft2pELqH6H3xaIBfpDCJlaxiecQ1p
aVx6w5OZdtE0HcVHlpaaKsevhRdvrGlq7gVim04YQ3bkKZsfrVtAGWb6tBfPD5jl
9RkiEDliTleACJeS8lR/C9OxTqO+JY641SEL6dRKE9+meyJRFCmd3PQ2Sn1Aj/eZ
2vLd3ugoRbVC37GEjQG4EQrKruQxECl5xqcoF3KQz3uNENQT8LgFmII148ghA03K
Ix28FUIm/xNocG1Zcu9bn6lYkOFRUDvljBe1f+U6es6exAsxq9h8tcfN5ISg1Sl0
5FETGhsQEhv9WabkQLxZmssQQWcYj9bmOphRIFDHi+9TiFWNobUgMogO3WALs4/M
AMJKIGbAP1N31zLwnK0bITWOYIdr9xbsqKkJy34BHHJlxXq49v4eU8FKNd5MnXnO
QAIo2KcxWahssErXWo/UW4W4dkIusSpwsNu4rTKIKgTWWPWtvKcO7QozCbz2sisq
9w14iiOuUay6EHZ9u9Mn6n6bFCzqGTz/J4OJzB27Kz2qTxS9g5erxH0i9S8nHhkw
d4WsPUNlkaLaX1GlN4jcpeNazH1mx32C5z5NEAHVrmHfLBcmEfNe1GeIOux94OZa
0q80dJIpN1t1054IR5ve818oyIF3Eyyh86qTyTK0rLKraxD16/hLUQPmdcCAIl4h
RsrtuJPCUm6xulbx3DGYnYNc5xgECArcJijA2xbWYjImCq2F2uBqUuJd7etGzPBm
+b16aHVrUDERf5vJu2hG7Y+8R6zVapuSYjSwdMne4tg84nF8NA+cY0njdJwA0NTL
V9YGlwkTpxv1whJt7gsIUYdEiqVq/v53Z+cmcayoFHeTczkp20NXKWU8hAPi4JBw
9kyAVswH99ddd6sW7zxzGmen6CRk84S1cPpKtCuMNwhhY8ths5vVMuwLyewN9sRR
o46Yvm/+8gv8cb6XEpcVJs358jDqZo51aicOwUW9ko12ZHdvhIbFDNoZhPfmpVPu
BjaP5E4rK6xlD/S48KxWHE0lLu1TTa3+ekDcb8HmZQ4mx54i7u3FvcQiHtuq3+/w
b11mBVJcIYd1gYz0FoO76IjAN9NTHqPmnjQEppGxG5xBmamZNeR8uT71TsbzHfHO
y5b1iXpZvzvpbpm1MJYrCtpj7z1cU7o93xWqproTtDZXQBRIRtuR7Rny8tgVS0u7
OEWNGejlCez6RnGJ1XjOFaDhnD6WOS7ctK7KgJncGLkZeKZ36wC7U4/6Ap3qPq+D
FnuH8B2/ElvFVcZKjv5xvaATYPdzJaibM4VOeuYxX2NrbCxZf+zLQznobZZfHggx
j0U1ofbdDJ7+vDdIHGweattwJvOJP3Y9jiIVribN2EERUd9C+6+gUh0yW22cpXsN
XJXZuyQ9HKDHiMQ7dsXkLFRjSp7+bbl4ug+9hnjMNZKkyfX0yY0O+YeiuE50xMfp
KVE/YLmpwxOn8N5BI+6lfa2JxOm18hELFYXAkqJbHPmEVuX+aQOXI3fyBii3bt/i
ThIVX3VG2q0Dj4S6g9B8P5HuG92B3H60lvUokESbPJ5eSyduRqTFStAzq3BiKVda
W2fj+dFWOV/ZhRFHNGzCXl2YO6ucOnnqmAcwh149q7lo1GL9KWsvPa+9JsE34IzY
taxL11gt97/Z8NcLU5r9I2w7Ta+xR9SCt0qArD9i0B0BbGjj0f/pJx/cFzAqtvhj
enyO41SR6wgIuBCem3BnwV/asu+EvIzPacypQHhqtFIkG3qajnLsmYjyh3K79iY8
uHFqY9J5RLRFKlNB5IOd/mD31Wv3hZp+Se+SFO4PwKk/wRds/DNn8p5732ACqJHB
lGZ5HVP14xtNOy9o1I8DqQGM4WM3//IsE2kWmpRFU9F8YLJo+imNHjibNExmDuUF
ZEAu7GVzcIzSp/BEwX2TnX0ze0M0RGXBPaTfiNuSWWymvrVPrSNsZmy51q3i7KUE
bR9Ln2L0IrH5Bv5PQhD4pzlu5YuVGpoplNAewFNKmRRhkRZMWtUOZLujpX3x43jG
KK4yO1Y1AB3LSiBzmg37//AMEBWaqZqUbdM7FkiMVr5X+0ixCZrbPMAW/iyC6ugs
IZCr3BzLI3Ci1nB9lzKYXDieyvLRKrUvpKBlQo4SGQ+tdgSW0QXO7atiR1PiD0HT
+1Ua11uQx81vXx9ad6Q0BO0B9QwxHmUQ+258f/8fF2GINpkJmgYgp0FkuAuTo8he
S+PMOc9xfRgPoWMQ6eLEds/Yg2qkaNkFMS0NZHvUc+mG2sMUqIQq4kdwNrM0zYzi
tvNmjp8N/jm0DDjjSpxvrFvJnSRzRT6eYxBhlwIyzHbMWZ9kzY0kqTK8LmpeEJc9
4y87qxLCxbUJ3gJe/RfyU221r2kCA64vgl/XvGX2afm8Y9xZsFnyoTVgE0oW6OcC
XMYA84RGTyqNvF0BcLnzyDKla3lQi9MVg+hp/cQzRkE/OQpBfMBP2hnKe1/NZ0TS
+J8Z/l5DvykCta+r526NWYifv1dE+pn3hK1aEnQKkovnqge/IeY+p4GFKizpEn+9
fuH7cMOnVqKWnaBcbSryLNzPFm4k+1C86qWyN9izuNhCzHBPKMIll0xoV6V7xDcs
KBkDKJgSrGBpuCv8R1x30VgEvIDNvR+zUPaX7TTm+I/WY5abvDqcn5S5CVszthdb
gD6ujmtTGPHHrZTJpf4NLG8PcZCFDeM5e7EuVRI3RJChneYHMYXvEx36au0xuwRc
SOcxhLIgddTP3ClC3F3zumX1NQEW5R1DXDHmp+gBWeHuVC9xgMpcdvDs/0KvNoPQ
5i9IZhZYOXEJS3dimSfgDmHK+7qCMeEn2Pl0+OYzcVPbenxbLWbIb5MRoJ1ixOpF
q8Q7e9+pe5VZpdHSnuB+zdu3x/n2JVJflahZ2cB3IEG8jXG7tVs7KLdDXipfYkgH
01bPCWTIrfj/t41SbHiXoCcHO8dbC6R/a9yMA5tRBHo6CgckV6d/ruCktPZzecSj
t8Bierbx7rjfVaFFQ/pfL64eOVJCAzRTNF4kr3YqZW05gxalJvlVBSdtjcble7mx
H7pqxjWZ+n/ux9Dpi8xq3ZcH0mneNuS6z4FU+1cm+GD79D50kNxZ9s717M9k/sG6
xrP1ZUTFt8V6uqCHQsViAEQAP8Eo5EjCl91OTr/o8vUR2B40aso8gXKidZ9wjiCL
442AYtjVNTXDgS2zSPivwWI0sNfvysckufcN8xbH4wxMuBxka1i8NQiBDr8CbWYV
1Lbh027BKXFZbeEii6sI7Y3cHg6IDs2MA7sActr5pu7Wzm0zCIDK+Zt8bKDRDZz+
JC3NiLnJa0WA9o+ZY4/b0HEwRAZVyaHamloxnQxZ1cosROrQwg97fb8Fr0DsQRHU
pS/1wn3Qsrg9CWCK5XETdNiPIVGzpxqeGnj6+9lmE86ClfMkt+4bU1Uce6rY92ms
YejnS02+qodtuIi2zdiEbvPu2OcRVgCzVMUjUWE4yskP4GdXETLjWs2Jb/j6ywhO
Z3M/OqGtdWbBL2JoY8hol9zVOi1PxrJ4Wt+Bew6cFQDTMsidWo74aqijXeWBi/jD
LWKYExuFOEIhH4hOYAtMboQ7mQWi68U/5wUWAU0guS0OhmT2LONgNOB37SdRe0UG
2BpWWVNQ1OmYgAwC9CxliZZWs3MPdNlzyHbkmWqgE8mbrx2Wduq8QDQXIc+K5nFd
/QOpVU8lW0K5pRUhOVIcZ9tuvfRi3BaZNHHn0m14AbWazr3YetN42BlU2MDB9hhj
7t0v6Tsw9eiuHosXgxF8PC/ho04/LtO4pWIknYLUBXjM6isG7luG17uEozbwHCuE
5cBfx4b0NK7zHAsmEkDN/EK/GB+vbACyhxoMO7JSuI84Wvl0cwQdwH0Ai9S4dEzr
eV4uT683jICO0J+oKptwa3eFxyZtSehHudprMEMg5xPqvjmZdbXtfEc4j86MsZRA
igRHEa1WimsSgU2rdx8lR0O1saEW0oskyBxz05Jf+cVPDOoc8vawRmmcmj2tdeB2
qRaKZz+6YoNsTNvI0nMii9mIS9Qer6lHpmCF6gCVA3PrS0i4mOYx/lcXZ4Wp41aH
6aScmPE/gOgzM8nkEjudk0fxF1lbRJl0UP1m/4d/h9zmmmDnFDVertsPFcm4XDea
S/yU5I3ojkq3An4N55stYLVZYLTLaVl9xfXo+dOZHBc/U27jIyOEosmxwPlrKj6B
PqYkzwYBDIzmB700lyUCylN0OOW8eNaA0E7fmsbJIkmKHZUm6p/tDJvBAqjKN2Gz
/1x4eFrQBCeobXPKlZdmh6lvX4m3b3WjwK5JMEU8I7wWOkWIuqfNlzq4CM+MNC3A
2AaWsX8Ctkkss8co1IQ4dI5hMpC48gLK2Ya2IpzPha9CtRhftljEWUs7hq5FcEOO
rryAXjOV7cEl6hqeqgtgs/4i+XMIcpGc03ohgVqoHewPZ7UA2eteEJgoirofkqfe
tizT9M53SmY+18ivRUb6meQ0ksYdIPLXxVi287c5HmN5S/4n2R3yn9WQuVmykafM
77fr0aG2jRgBgJcbdDkwQtg4L8EyjhtfH8KMxgDbWFvy1xYUIQzVvuz03YZrBEBh
UPl487FVbKB3qrBiDtdw5rK78pBgUuSQIy4V3Aqj+kc/11E+K4z3krtQCAjZH1Rh
FFuuMJjKn5qATQxgkWCz9pSJjJkwu1k6k7wPidwo+MoAS8QjJCHCrcpSlnRIOguS
eIEA4z1TxOk35byTrUPltVJQfKWrUg+ZZjxiqr9ISuDpeirixKQ2LNb3jMkdXvx5
Vf8OAAnLS7htnF3S1Gi0aV1qvuLOQWLI/vIhRbfFbQJ8o6IJtfdDH7bB3BqG5+B3
GZtqni5mTgWI71qUGfyr5etdX36pSWyHRGxOFbjtDAytRwltTcYv4SSr65CE5hMq
vvPfVLsuXZxvoy1GcFk3/DXxKu/O4XjkqE32KhfYT0FBue+txJtpQuInlariC1Q5
FrajiyFq72UIftaqVl+TDVoQOSezvnF3/9ebj3jtSFyueCOw779k3WhO5TPWkKBn
unYsWsKm2e6P3oOCdzA73l7gEDLhNJY6TmIAk2g7LpmL80ew//DbeN8dwtXKqEQR
9k6kwj5iAzh97N7ahUhZ5tL140gd8F0/0PqaZr+ll80mwRkmxBWlay9JREZBLIpP
UnHXAkPEpMQkRcnCBiTMVpgcUlQo7vc45VCzb60NXQBGXL/LBPdtUeBqTM8DleMn
aLVLJNs7dTm/HuE91E4yIxxzipCvwu7NrI2xdJEO9OW47TJGz9Tm/dzYBd5uoOAQ
py+dKBKlemUq/+PNDpZ0YLcS3g6U/TWmpBqE2J+TvmdTZlJ/xqgCnnz/eqlBCKJb
Md+JmtmCbs5aBCCswLDs3SKupH2xLKFfzshnBi6H9oBTml9iH+HZUQRpVCrTD4kF
NxwekMY3NQn/xk8SK0ggABh12LPML+drYPu82h+Z407wBGraNAZF8lhjDQM+j3X7
iYE+oxhRcAdSd3isUmiMhIizGkQyltdKQmVtCbO9t/QhVMTYrmRerhuTQBDH8Vv9
MW/L8dn2l2nWr2rnZyHCgTeaNMJCjSunxYBpvkUtMpND/aqbD+6uqXpKCHSsd2Yv
BwzN/NWKfBrfz16+IUIwLktfD+BYC2Ev5jUkDJFHQ3EP1ejOTIC+n35gLmoPYhOs
mLmPF7N+1lBJ1TqyG3jNyxyWy6rriNhgePBWKICz0vEAVmUD0hDXh4HI/ewECkA3
UUDqlT8BmtugscIuY/4Hvnrvynx/mY+KSwCowRoIYggxh8c78uJ58PRkreyocj8+
PJQcEcm5kBviZRuMdJ19BpFXfGSJjvVgIj707IkJEvrVWb+SstD8XxHQdgw33VOL
Z23NTuTjfa+GunOHc1Tp9VIzJEpe4vUyVQm11Shmmp5vP/fwuywn5WYM+th8kS4I
7PGvHesWuPmhubz6ZJaGryQSOAn5NR4cULmiB6kPVKkrisEMvUkLUgrIamgGj7DQ
smoLW1Vpx4661ZwZVoToIc7SDXog/Vi96D4liV/t1TBvd4QXQiJgteUQ01AES0Mz
p57WPw50cn9b0xBTPg3fpHHvrEB7WhH5T3bIJ0/i1kdaajIbcbFxv6voyvsoyGP+
xaPZ1DqqnyNHnQeLQliOO/GTkjCsuJsyXixm8WemsfMDXXFtYFAbE5wgjfXLy6cK
y8v7Nse3ZnjOSPtCBXefsf7E/qjFlM1lePS4ITuGBKUicSo2KL7TmcSJe+ueQu69
aZhLHZTANXYwsn/Ap5VNnqIX+w9S/r1j037AONe5a6ivDqvG5ubA/WVTZwJqb/OF
zpKVZ+aVn//f7HcuK1VDDnde3XC+VJ2KmQGpXVhmXlqkdU5XgUEHPrmNzI/qFB5a
hiKggqKvWE6EhrtSPaseXr6wOHJmMifmsDbKB+4srkGdZLhMeNdUC4JtmF8QU4x7
uIg5Blmz6dWt7t9EHanXk6iCtc8J+s2L4iA9Qan5dJFfd/xdJ1uATI19Vy7rt395
GUpD233ThslExa8IRcbA+tI/C4HnHS7WsWpLy3bdQo+zN1WbD0uQMI/ZoYHRo+ir
HZpFDuEbIsNHWGA63dk89HxY4U1XWjAHtdej30JpC9zBJc6uh0ULO9vWksWyq9Cg
hZnMSk8DQoqp81YL9IJIc3pWA965y8NOsMlMkcvJtX6OHhWjMEvzvgoI0CYrgwbK
XpGn+vF/B+kgyuqZkWpDqsuKwCo0IHEwXHk5BfWuuFGOrepWAX9IgbQdfFXH6GzR
hBaml4SgnJ85Pe9r2eI19apU3hpImPXRpVblh2IpovPFyAw76cPuUivfK4EvOQuV
6dgzjn0uGY7KT6/rE7FVnG7L/uv5Y6eNrfF3w6+0kHYj1vhFQ83Z8r8dMxWlJ7vT
paJgcyjg68JxOUNVagVK/Qtm9caz8HinhJbJCwJBZKE4xcGBRArSTrhT4ZKR0hLF
KP/DGz9dBPNZaKYoHye6J38U52Iy0oqjxe5sLpBn39oP3b6vd8VSK4dGp1wVNnCm
biWt/h28eqmSFa9L4JUUrJUt2cIbe8cHeT16uTiqgfhherkKFbQ1Unv6DLA0O7Wh
WJvVnGyS9Vri0P76WODYmy42YDLC0mRmAMQTMT6H6QncDIQaLJ37LByUUAD3Op/+
e5K6hXhqt/IKVWg4C6QCLqFqYcb3gcqizcGChphrFX6q8GWpBlfurpQLb6RAZ4uH
XIJzBcxOgSQ3lnFb3k8oT9amji6jrtRBcAH7DR8lv6a3bFy4bOrnvru9Chbd8OZz
OKWnL1qXjh/9kfIZRCjxG7AQjX49cqcgYiQyphzLq3zlFyHxvZ3L3w6WKrjZQknJ
wNaakwxnD8Khx6M4Yu/jotec91RziJcuQSkYViUcaQqPVT07FC1i7XSgQRjJIUw0
uHqI83i/RoxOy0yAQcDrKVV+uqFaVz+oXUsJSWRSOo86E2t/XlMyO0NyEHuNfjl1
NW/sVDsaToJrA4wQVuWXqeBTqvXJv22J/i5fkNx7rN3+KKOTaFKoLZ3KlAG9DSEm
5e44aaPKF8EITok/iJGn9E75WhZ/RWrqiIKDtbV5Vm3JNkIeTg3BLgeHCnpcUOym
ncBaG0773/vM9hCr7Pde4WpMsY41+IxDzQaoKjagfjd/ip0Ag2Gxv4rwRPvybrkX
+uhVGUkFqDixsSH9I07qmjXGknqZ8DWQdkL2w55uCadOa+entiow3RfxmemN3MZL
hvDEHylX70cp/msdqg0+LxH8zpJrhtiv+5FE4NGJMg/ELzwreXth0BzZVXPlGywu
m6HOPGPlXj4TBhI9nxNVyMz382vyz4XyuV3bVWAjTWY7k8FYQODJHoSPas1vcthK
tn2A40VifXQVAO+e3n1qQjkvR4dyvUdDAk808259VxlPll7MunqtIeCNM/JETshh
5wxp4pClJKhthdCKlvFXkc3ND3Y+bkTO9wUN8ib9Aqqau3+u79cpymCb38jf9YDe
qye5ICd5am5LP14lbLCKzkYFFcJbAIkC9eoPk8okRI/9hhGsVjOZ9qbQv5wvZD0E
UuxIpvusFYRmNqdtmrfSBKZXi+Px0CZiZwWN/pewvdjyzc5kZGkneN57c+iljmy4
foMNwGdcUMYjt9IqX5rJMsCS30NbjUibEEdaK1zWPPYg2CKrLbtqDXW3BJTDY7GG
2Soc/SfpE9gVaUGx8MMvabZo6Sx94lQrmIJn3nbVMmdh6d6TT05lVahos/hK5k48
cd61xCH2sNuvRbipUNu5iGrhL5eYSHunyedJ+mZ/YymJgzYwBIsonayGHv0LOY8Q
0Xtz3Vwf0IDDIKOT2XIRo7k2JtEz32ixDPV/YZkMYwo++Lobc6J1yVIS4VFPwhma
6VfQ4X/hu0R1cZwzBGZm+nfwwvadL531HeUGf4AwQelyFaqrg0W20LyPTX0ZPyZS
Cp1V/Yvj+d0xmOvOYX3IvVc6jefXVAQ17pbVvoruFRytz663VaUhR/77QumwBd79
vUqm3U5TzS8kEypTbJKsXssKPZ63ArVsPR1weQzxM3DZZsOzO6Wq89yZECd7zGGK
rsNGocXcxNdn0nrQfE4NtP+4Xp2ywqnlcd7h3VNq7Ye7gWg/0vwfqOE9870MHNkO
cOsq9zsLNP/oTNU+F8sY/VhZu0jebhYWZp+vm+v7CN5UEgmb0WVjN/qGgEHfJ6ys
7W/mhFbfXxxYsuE9em+JaKn1WzkiQmSpUJmFRHxnSxmoMU9xQOB1RkONk2j0sRLS
JMKgRnsqS3W/OqBY4vkzq4eNzPCUKCSyhqJbbRXLWRX+xjx3wXbGHD4xHlkc6Tr+
sPUUavZAx9pgjI5QPUNuCvRtqg8h2DQJ/ynrPIDc5jth4DcyvkO6EgJ394BEJh2s
/mgF4OYeuY00PfSoO1AdaXa0+EaC0rDvqkNO1HXROL8C1CAu61IriG/njwE7Tjau
oLvtE4IqsNJhqz0GsZhe0TX5hPuEKoUqST85aCRmxmrxtwzlr516/y6HUK1Qg5a4
Cf06ZO/SVcmu9AbuBdR8nGRKugIGd+LQJYrw9Dqa31h8nc3hbY70K+h5FnJwzSAE
wTiaHZO+Z5t06mBRYNPd7f4GuQBkI17s0N9QbgeNowkhPKwNGZPtU8JSCe/iyoL3
yb/cf/2/qnYZ63lYeZOax810RTIvFe3fXdo/Gyl/u3izESvSgkYpGg3ziqVwZlNU
mOmp44eZF5GwaBhkNjjFCkrdXrhqoZNHCmSPPir+mqyqQ17MViJF1MIcB3Rz2guG
oxaB8jFK90rvopcnQsxi+aTqT6GMW7FHL+O80XtiOay4dRsZYl2BlseiRDukOsg/
7RFzDPBU/QiYH3x5OdfcnIN92rTq1rQNB/e0jxtzN05bi1OFwH5/D70FryuARDRo
+fBKtkCO+jpz08QySiFbKZABQ5W6khgwvE8sj718VN2M5U1IB9Pno4yqHshISUCq
Yz5v8bOxuia1iGGqb3K1KF6JR88+DAZtxYNX/zffD/MgXuz9qfhInirbbS2ev3zz
Q48uu0y5m3wnWl21qhrufpTOPudvaNCXeAhG2MJTVeHESg79sIVquiVxVq83GUN7
dlyeol0Feo4+diSqsXuZpzEsj6uxps46LvO7J9R4TJrn7b2FYiy8qK5Tw62JHls0
M8s/8PJUELlBRXrKWzeNISjD8ZJxsyglU/062pWVEzP5rA11jEFodF9vKr7KOWgb
fwMWj+5S7JMGWd7hjpTQNCHIT/mqJQbqHIX3pCCNjncjFtGQtShVLyU7lyslP8/g
hMJ1LhFsTrp9H9XTxfjZDsGa8BGXfB0UIwaAC/w/RvY6Awd4w/mFLN1w/su/LZD7
2pVdJXVcZVgJCDlza44DRvdaq9OBX6Oi6RVos6hsJN4REVp5cHoaod8QpraEIhy7
C2dhgJAZtLcxx6jCSJa8XqlVXY4rCaeEzr/T1Hj7mmCx5XL7UiF+OWAIZNoZ4Px0
PdjTKPbBR50b+SHZAb4uP5J8ZzliyVUuLbR0dLg5GEjZWXJFCgf7BrMPQvxNeZoV
U0/T7/GqKApTjgtqXoZpNs2f5Yi3HHMvp3W2y4l2uFDHnWb/eV0r7vk3fGKe4Pu5
1dDP2SPkZxpXZlOQfixkd4dp/Tf1TDIkA/Alpn8hRWtJ9vlAfgXz8MR6CDdU85/0
/OIk45+9RtnrQbARC6yD4gfLrG8uHeAItismFJMz3kuPW4Ki4xMDBM+9fg0MPlP2
WBzq7sABreSuqlhuG/4fGp+ayJvMvcWINyIWrrpo6+zDQ8g9ZOjWU7tfsFCyqiFL
me0Ov5fPinXbyEU8nlYTIJEu1FbO2P9Ahd+ACOp+S8E4+OtkR/omwR4efXrdE+BB
DlYKQQNf2zZY7OmIQ+V1bMBe9m4EtDm8T030Ahbe0iSqpx8EvAtQfXb0bEGz9tcJ
Q+/nKyheni1mB+8TvQqmkQ0sxML2XnNFbiKmTskA6RbstZdZq2KjAeMwLe1PCOcf
lrW4iZe7qYzND8EHUVv3ZFJYZG0eE1iLYRrMRsXbzd4uc6kIL5JFMXAEt8XTHDt8
T8QwwcSkmglXsTKo6U85oXdXQIQRUEXF75hSGsRBPXBnh24D+ow65h46tcXrY/u+
VwZXjpR6OpK29Qqyabc5kPIT9n5O+jQpN9TKuM3faa6SBoS7nyKB+YJ8rv/go7rg
O1/hg1s4pZbL9l23NrSN3kgBmtIoPHqejOXqaEoNuofei6vZpiAzN9HORTnX0Not
0db3jg9MnPqRqP9BQba7gmmN1nZuwEivERPHpcjl2aQLbA1UbqFT8qSImp36Hyp3
MEWp1Fpiy2R2gtKg8Rs1530Fke+9plWB0Ifuvg0NcZLy9C7RuLmGUmFslE7we4OJ
jQjn1o7adSyaHTkTxcNQmz9LqGNGhJilHV3Umm3Yila8+DxQgGpEBaK1D9zuNvQo
K1XmhG9LtvisI2KXqT/PKGPZaFj2+BHF5Uc7Rgzpb/VwBWcSE8HwwzexQq0quWVU
+j9Qx/fbhyOONvXWYrlT6ikatLhd8AOqXmait6m9ULs3btRziNOXVSWHhm/wlxk3
Bdg82txPkFwZqruRRzgghcVk+6k0aUuqbap9tn5PXEPbhcVQBnn/HvWEIrw9nWfW
o1tS76p4K0ZXM80vsYM9hs4ur5dJqynmfZDr2wBJ6DiVllmyCB5peH2xvLfqahfv
dbhmqHlRxFMzknamUOpfeeewfpADNWHM0+XDFtl+ClRzcIgT0DYkD75S7HVFpxDq
lqvbgvvvzaLuR+72oTHt46S705AlrFuuE7YvFDu3Iq1mIaMPo1OsAli8UbbZA+W4
VjuPerO0sPtabYMoXylw80bh0IyiLOKhQV1SghEDPxxBJx4vdLE4wJtSA2X+2LVs
nkSRpS0TQZ80Qa3HOavYmDFlS0CJ7j6ABXof0SASSnh2wjQEHe9Hk+DQJ7nwtq2d
4KDwXfViI7Zf3HEYf+tAvGMyuCqZJA7F8GSZEqYcL7rjnGtQ1tMzH0uy+WB+QaWI
+Oz5TdR2VCmXs/eikcanqZSrR8Nd9JFipNV1XVDgxRCIMCuxUYcu/3WfGGQ12lRx
jSb1h26UW+oCfIYkCgL4W4d2pdVYwuHgsr1qIOrATPuaCEHnGrLYKmuVV5TDPD3l
icuOloX1B9GcB5pWc3z5rxEqbM6f233oZ/2ha8DljmPjjbrvS3XajCACwe2tcfn1
sdRvegyI0I+ICoaidGbBBesebinzmq4hCfcZZRbO3k1eBaSbb0ZaXDPNi43u6nJp
QATQ8cyg+Dg5rTBSFBDhPZukJu3nMVOVSRSectyEGG9aZU5Ff6IY0U434fyGXmFN
isSMU3VcUKoXKCwsJmoj3szLkRvjDTt4pNKnWzWu06aNHti/edyKUX1++k5blJyj
XSDFb1HomRCqDZPxKE6cisqg0jIDU4hilXGVFypnvKDhErrh+igYQDcdwkDB981g
8Ggj5+pransLD0vr2nH8GaiasnZwp1xJOs5k92kbQxS4gxy86Dh8SpbXHVtpiTtO
hEqcYs6m5Agv3C4eRhffdcQ8iARfwkUXuR38X4jQzLmxNYMQ2k7ckqe2qey9PPIK
zUd7d8KvEKUEkY8s6GyCj9seOYw90EInOjSAXr1G+EIn27aN9YACpis5hScjvfxr
hBElvAV0Hvf7Yo7u9nZGuAeUsq02aeR73aKyw/FEz3LjZ9jcKyTY14h1Kxv976zk
7FNnc+2mnw3Sop8Wk0u9rbrY1ItmSI9GVubuCK8pbluLziyld4UgAG/wvL4qRL81
MlGUJRCNyOf9wDIZ+KjoUr+Ax6WK1hxx5fVwaWXSSXrAxMhmLYUO1ydaX0Xa1iD0
/+I1KUToZoP51h8rOUJSst9IQICzphU9bRVZIVWl03wtATkPjKCROJ4PNaG7Asrp
vNOmpab5PRKYA/CJ2fxtFKCL77IkVAYl96tj74eSrYLXJn5QOQR38VTxxOykp9Va
+I8rDqp2ZMIyVrPd7WK5+8C3CYW2TYY/hhqTXf6iCoQXbP6MdU2H2iG6+nypwZnR
ij2a1rjAZPrLr/ZaJ1NWdsWzOPlLVwjH8cPhWTGmI9q5tNP+UhVFU+9IH4BF+cRT
+lL11P8V2HW4tvVMs5vaU7ulx+hcGp6LsOOXZXeuWBJ/9oM8TfV8SWkWyHIS0T/H
/DPWS44726M5pmS46LHta83qbikkcbQ6782rJaKwaUxUMeCYq3sV1KFWZj0WYKOK
Vb4FG5uqT4J7Le59/T1hfCQrD/aObSPmtAjVC3rgtFz+nvlhu4j45IyNqRPbS56v
lHQZxNUFKnWI1rfMWvv/qxfC2yFe9VFkO/MBLn17IldP5X/4gu1wLdy87mxVLOw7
Kq0pZgbeZuTn3kwLQ2Ss91JsKAqdtDtzYdp+lzs+ebUspoufstelkKrgie+VfORb
hsuOammjyH2JBPvgjduU4D7SjoPFDs2CH6syqSUu2Zgo3Qdc+81u0q2TYyaFhAZy
vz8oFFy3MpbMrsqWd4DUYGvY47Mf5ewiFEecQPIE1mS4HIIkw0vGCX8a8zds1n/J
Oy8u2MoUTOBs+YlUcBkFCa8MzJCCFDz03qdea68EcsmG8+pQn8g46OUHYohUmpTv
Qy3y85is9pZrCtwGsnKtABwgYE8jGf/kIfsccOwNMCJSFxXzFsFuyJI7C3hSW+sI
1MmVwia/lTr8JAPCkxirdxYEdjYa71TJlyDGeZvvkyDvhVgCFhXeqnhVv/W2rgPS
M+MzA4WV4N95NAXbSpxclbFGldHwLbiurZpMgpXCB+8zGvzs6kE/kfHOxt4cWB3H
Tae0O61VzmMweje4fZPebzZRI/mvnY8Ggjw58dV5GhNzv3FzXxp1xDgxHGQ5WNIQ
5oxdg+Vz95if74E+UnvEBIE7pT1G2enCXkJAPGf0lOwcs7b5u6XvuD1bnVbdYuvj
wnkU2dlgvNIQusjANXyQ6mlMNB4JRcdCQYwk2TUB/Vl8E4MLPof9THk/5wtK3Qzj
8fJosEbPV9JxubQckA729wQySIh+qz4dAGQ5tGoxWkwgh7WF/3Wi/BDEG6QHuHfx
BxF53VSpNTE00H5g0Tch/f39qHzucm8arjwHOzUk0xUTZSYcykIbB1qajieHr72H
stvjx43Alm5cay317N7FI3Hag7eA3xC8D8YiTUXv8GuIQX2sAr1MH9gVmH1aOnbY
ph5VWATcVn7ctEbeMHopKBrdluER/uJR2R03ruJTSILkffjx8uIyZjLamzVIfYdF
ZngOSMBNflg/HieDQKQSk70q/DbZ+AjEnxq268wmPj4Zd49DCM+OWh6ejjzRz8ZF
XBMWQpyYxWdlp4ZYey/GwtQBktvQqLwdEDja/+3wMbNCNvn/JVH9N37yTl9Uhx4V
NhOGpQP1qKZ4go/Zi5HCZSIkZRaYoH0yDTpsfsX6N/eK4CdjHIVM2UYXFgtDX36M
hpk8TfccewlmHL1BNg92adZ/WNM71roXDwKq5PmMX499knOZkzIbibtakND0xTga
6bjEhxUcJSqDR1wu+WN4FX5Lk9zdVPFj1K5z/NCTUpKToKP4y9zQTe/4kssFwEX7
m2nA/UrzX+7X14hZR5cSapwHfjvdCrPno/jh3EJC8eAk/XhSnPIG3Zcliwv3usNJ
ByNmaEPVrpaMzhtHnlKQAt6kny3mCLD4fPP9vs7l8tq6f0EQU/ZBZmj8bL7KIM76
wQLsQawvC7lNAdoquwXy2lBgRdQrusc6M5kqEc36y2CJasJ3erWDnh65F42PXAMG
7behY5ZerdLzs2fTwyKuu+zf43uKItN3wZifyqBjxaCp/Zedo3MgfFjPjIBb0V2b
S9P9zpipFwRWa2bIhhk9eYT5A6Btg0i/kUkdJq+pQNbXC0yk89YKrcmgfXVuOPRw
UoOQsu4Jaj8VBucaoiGFAp1c7oLtGL6bSenjgAD/vOkfX2KGCYMB1PswTE45WdDE
1ZN+jJj+kk805Y1lbPSqM3MzDeDcPhbN6SPrALTH4X2KKQDXoGtMk6LCUIQEzBkF
AwcnwP+wza8YRozjhGmQFKyI3vF379c5YC7gqNZhPS7RmpfN9jR2a6My7U82RS84
6RhMKrg8/tzukV9zkt+YAwfbQuwVM0M+wGEcXd95CClqf6Lp7wH7mha6K6IFgl3h
12s1ogPHdfWVIE58M4Aa9ORp5fGjjvMZl9O1Qj29w/aS1jDUEhy/l2AX98WtQi8A
NZ/1TEiEy9nAnQqbWr3mZD1IqUpImj0URQdCJUn0z2iYHFfSarq+m0gO3ZWNzSXK
VvSRPzjQBzGExcHu/lbhK82aHvImRdCDjiftR25ykuOdlY6ieG2FD98lf5SOTCSf
GDesRUf5mu89ld8akK2GShznRkMCzUqCH5MDaDuYAl9dxbZmkwvaLPS2QOV0B02C
9okp+1vOYCA82xAN0/T6DycEqOd5ySXmCQceuFc1RPpaHvD+1EafQj5fbsjp6JcK
F9KkdoUPflhg18jcLNkuA1KGLczYb+QDpOUfV0istV/1C4fxxFz9ztP6hYN64Djn
9tgYe0E+asx8e3JZkQLPyqnRwHO9RX3UXnUJFtyz/gkQpBiE8dvSp3si8B5Lbyp+
e7edKdMsSEFcmGDx8HUFGnaMK6pi0Xh51F8aEQKauuKUy8KQjTd/FBkoyPubnIIx
7r92NzLuIp9cyck41te561yozUd+45QmwszaZLHXzN2LsKOQuMxFgWBxUWx1cJ7c
d8ALAy9Bf7puQ5n4tF6Gdg0WRL4xWAEpP6aUhWbuofu+BcUQlIruCOkjEHBIDTO7
YPL24QejjbJcyYCi/CtEAZvES6X5BEoFXSyJAqa/6jVcryL3jZmtue8bMVwpM0oM
g7YzaOCPyT58zxJ3QjoS1Gjfd86pUzfNg4v9D26r6FmY1fAo7EnzLKSg8SLYZIlP
r69wU8DtxXPvY5suyFl10oi6FOw82MfoeQfl+x1+pQNIPHnghreXhBCvp9ILB33T
s7z+VB4pijK6R61s+0qRlsLLtzXotJpVaTB8UcbATHF7l7n+9G48+br0Zlfcj0I4
L0EW3/Zj4Veg+rhSH101LJqq1w5U+ecDsgF94NvViptNkwzftbFrxY8wPnUk3tG8
4d/50dtIqSJ6TGBPX1LS13imDKMapgKYv8T0GMJfobeJ+lCl5kH6QybjatGccJVJ
+9uKN/lMDJg1I0UIfAkjsKOJqAfvzU++KmmV2zQNp3qZ6wWe9i3iuEsg4hyF2m82
xhR/eF04RHvPqjqptJsR7e7qJjD/1KtIRT2wR1etUpZZ+LGei5DzDh7TlcEdo4+P
PQsHDAkxVZbL3NGxMG8PDTEL5y9VR2Q99WfC07hWXjuhYbhBhrCbP7uAOVc1LSnf
ag8KCrkr/MW1trrdcXMzr5zBP0BUFiMImM9h7alcSH6m8dqaPlIxfoMqpZthEVQr
kqRxb6hCT6bdy0vpxA+YoKz/MPgqS6O6ZRjMe0cXrT2QoYFk1GBMP9TjfRoD/u0J
s2d4Nc02GlzgSbJwsQv2mngCUC2Pr+NN+sfdsKtn8BGaZqb/dksmPDirZK3/+0vj
785F2qbC7bOe9m7Bruv8w9N517Cc+K0L22QDJ/KXAw2+lTX2EyCqt3wIELd3GMWW
FMRLBKkt5t08g5MawPOQUCqr825lMJNTjehRUbTZ0RUulcG4zGiAGl4klYDvnZAR
D1Idouu2OPZoUc1/LVKdr8B2QmZFuFAYOn0fESyt/RGeUId6RQi49J4q6GL3FCYv
rxnC0Vv2kEAaEon9HFeQhiPcgAq0VfGR5gAVi33i4CoYeBKMXzOx2Z4A96ga1EMw
Rx9TGcvGKqw8O52KMANTaeh4ULVWbOws6VDdByc4zWrgamm7OSEvzxNepmA0uHKa
9PnA9XHg286Gq6Alb+WRKvEkmQ8rktQVm62VQnXO8jMNN1hPnGuSrpPI94p3YbrM
pOPXBFMlaGpE0CuDYSUaDe9KGhMFRmV7iJS9cdKyBsHIebsy0BwS6UVpbv2GknOo
QJlmvDZ2Pj2EaEWZBpHlhw6Hg9vuieMjcHDjzYyXAM3xovVDoxd9/mpBt1D41GZj
K9+CVGTQqnK88Se6ndKKphrXfTHRoJa//n5hKkoveAiN24rc8utU4YwJXaL1EiDL
xGKuY4SVRxmhcoFqsy69SJbkmbqCekg2YrLeye7LwsjGfOyi9tNQs0lqFdAu3q6m
gfvSabtDtpaTl8P/NG/CwcutMFsZFwpCRmsLfWnMji2WFAiUl9Ha/ym9Cpl41YyP
XjffN3vSdpftdL3dZIglJCXis087ess8B1CUi9gGLPTCFdMyhPX7akRVpAukWMSd
3FhuIIPFYnco4y8FT7JwhyvMLZILU5xNk3LaMk1RaKTGhpRQG/4l/MPzGd/3vCr0
g2VUomMkb1KJxdeQVLQdMXxieIqktbr8+RqB1VLS4SoyWiGWxtmO3gdrdZtX8ETI
b+mzrOLounhfvlgoCyLBaMGlzj805UezB7wLP4Ag3CTm1TILSAfYrWUISBwiR0VY
yEtGG9WW1JTnkcvhdSmJzgEBQpCEdLp7w1oCCsFBy560gVJscfwS+Nax1CS7WUQ/
tM8xqErk3Jp3rWxM5I+tWnLvpEGqXlTP0q3LW9lxqlvnLYf6ONQI2rRGrezWUchx
YhkMCPzIWl61d697ZAZXrGH39/KxiySUdj/RAyiRa8P9At4EIdJq/WVf7xRkITfZ
F6qQzdCKHU/7rrN6cgAztk+qw0+V8zhoJtByz/GTeBC0DvVGVKa94t+1wVYTNDLJ
I2gB8KfHPtVmLCDxLlu9Pp/uFJyTKsUvso0oou0Feq+vEGpShcAIYed6n7+VV+qy
SxRFu+ItC0WtVd2iIR5pNvxU4NoQ3E7ANLxmw7xa8yMWwV4i3qF3rDN7sfPTS/+K
1o70xVVRJ7xaKFZLOLfbBm9NsK9wmx66dAJaCUw33e8bI8ciL2BrlXy2kSvZYHP8
/ld/YMB81ugKAVTmHswFtPg8CQ8/lcabuzMpcgz0kf17dVU/bcj5KNoS38brfFTk
PtT4TI5SFRvhbyaAoFLMcpVZVfMJe42/YLrYfCgxhJjvOd5P7fUaYiHj/1sL8ToU
qHja0Hq7Zt0PvOdPrZTatkllAf1mz6QCd9qc7KhU6RoQ3ZlYDrPkAblfM1JFf46s
26Ao3Ne6To5fhu4gRqZxQhFczGksKMjPbCW3FT6WFlJbTFcF8JxJdWs366uYIHma
KjyrS53N3K3z1WD9YEJDUjMsT8CXi3Cwyxt9goPgY18IPnouB7UganxcZmOSyUqd
4YGS2KYR7bwiAzcGxX5mo7fkehaR7aeSWY9iedk1dVxe1ybBXiwBQpKSDLijkbT7
8nlQ4HITPWUrsTHBu1nLgRnUcE4bAH0aQkqutNKyLtHMRUTdHwEASSM4CTALQ38X
9esIRyweNlopp+CZS5Bb/ZzUgxds96aTpuAmTi6Z+BNvpPWNbv0nc+gbc+zijJDj
54dQF30yHwyBjMVNpy4qgDZHkvT9rJ0GsMlgk4TtYC1VXL0+cc9o1daweLVtBCjd
i/8I104sMi4BzLYrRccsoh1h3Pmc0bGcxprvOVUqLol23uPL/LBt6XNt67Ah+oJc
WRr2bkUmeuT30fbooHzPf1aPJmSLwbGPlWA2MviCQLWXM69/kztCXL9mebX86xGW
UuQdLOohz/CofYMyE53ROYBet4WtFPlQJRoESzABLyQMddl2DtzsHt6rWKMQVo0l
m0D3yqxkGXRJOwfaAqsveX+5UBxxuMSTiVDlQMJhHkP/2copiyRq/+Z5CpjdP47p
l9niNoxZe1X7DLXUlteXIjrDfL6UjV6NRT7lPX4jgHlpyuM3kAPCgc5ATNlXAs2d
nH8OrkeZ7h7zs7a1al3lfTA4f66fnRNPlVnK8alD5vRTlXpx7TihmdJsxRWa3+bo
BZEKV1Uy0v+tznXu4DCNAIjU0GIXFbKF38uvbZDgLE+1fxpyWOta3VOpikxI6aOb
6ZvPIB8l1hRx9HokowihrnWoPBjkhKxY2IzqeQaynzElIuSlhrwhYvUkPrVDGwmm
AVA2rGVKL3ss5GrfEpM1Ek2+C62W9yWg513v2XPvmitUGvceRwU045bLMXkmFw8n
8nvz6BFqFzrnhXw84yi8Emnh0C83UpD5G0vaU/8bGosqG8Q6ZFDisswAdfVVVq0m
FzkO/M13mKVBCgrnmPhTt2VRtWo9wIoXMEKxE8AZ/AwqBry46tWe/Vu5j/nf82c6
8uw+cUmR+YDKHf0OLA20E0HStMrL5TRDuTqF9LZk8nPeLeILwpx4XnjDKjB/CPah
luZvx9TfVWmXS93QDyArquwQvZSNp6iWrM2DmQ8HKxLxLoIKwEjbcgNjIZ1H5P/x
0EL+yyjngISMxm6A2PuA7+IYzXxZJxc4bhDrNebZcdMe5AaTyc4Px1gixDCmGqTQ
5U07r9R6B7HsYP+F28yIbXiher2st3hVEHxG/dGQa8r7z4diqNQzA+t14X/VlnhT
gciR3GBIuSUC1sBlWZuNrDcZYDrOR0T/u6Nfm3AUXGXCDLqmAAz8l7kibyDUIu3x
4OAYooMKWddb7d8EllM04EOgRkSJTtW5AfyfPK3vvSIqPOkhHj72V/lW+jcH0a1o
45czIn/NPTkQaAAkOKMpg9F168t5hsSYUjqB0tko8khMyvVfvQOynZmbT22yRKku
Liz3hLumOYd+/g8L8OljFgkepfoo+25E4Un0gosEmqx/kgYaNWPjw8BD/JOYOdRp
A3PTfOcxxm1BgHxGerWzghVkom7Jj2OHNCF7wmMJVZVkYqsdAhNdtd4wrR4oHric
L8Hc9/l4/ou5FqLtECJS/317GDzqsBxCVtfgByJYwPLNOgLHhwCiU5DIMrBKWm4D
g+RuKvG1cFChE1J3+ArXnWby1LP4BreYTmLAUTu3OzJbIPY2u45K1Rv/23UjFnS7
Ojk3OY8RhGGbD61jcwzEabuMV11m22wGV1z/GgS84PGDwmVzmdVZo4R65IUkO7qC
qO+mi4/SKfXY7ODhph/jrIbp8KJ+STXrvAYZzJ77vWWy06yw0T9Nnx32ATsYtIzh
etWDdFbSlHYPB6uNdsyICWwD+hV5sQg7dIUfwmvcj8yKG3M5Q7rHqFffuo5ZpSpS
lp2hVYd3hycuZ/Jkbo/CP5QuMHSFQ7S7HJL9BxY+kdjJqFmTeUVRwny6ua2aL4VX
lJxmyhASwCeDQc/28gIRyQ0M03x9IQZxtw/uIZGX2mYq1u1ZnxFWt2O8mhjJ7aet
CSUAxNoRNyiKZwG8YMlUpPEvkVRMDZ4wgqOzwKMgGvs+RAMcq2rQ69JxAYe5Kuo0
DQZ8snyrUtQHY++3UGULsoSzc0dkzkcCDbVTHrRpyg1aS+nRRo44hOTiLZZljHph
ZPKrWcOtXEoqofiwPNJeZVKDVRfPY0+m1qX1pQKX5xvDOz7Mu5cXWUfte9+R+LvM
PJko3BW/qlgrT/lu7gclq0NaSdfjJ3rdfEznZr+7Q+t7K7hq1OLdMzDEFnVcMRCo
+0+4MLFJwP7hB2arDAKzZotz/EY/FlMeZDPZxrYGncX/RNR52peKUOTeOCmrtZFK
FQyjoNtedIt7WNDz0B4OZNCCrC91ODLu8G65C/X1ycQORgho5YDwnqNNw/cYOyZp
4vMmuqsRiC8TqiYfKjCOE8gkH3IfiIXil7voeyA8HuxaWZqeaAozzjehiERZ+RZE
2REojEK/MC9s8wHugN0U17Fs4EHSLs0BwAQbAc85yKTc3vgET/8G8vkACo3gb1q0
TCZRjL+QN3qmq1Dm5yuz5ndBiQK9OpG0w4MqY+8lh+jTTvzWwnqPfyx4H6WobIym
SIvp6fwnILKMh5fV1QH9MCUUfdZb5mXM0fMkiOHTAcv+0mMi8NQLsysHYmUMp2bV
RJlEDi/+WFGgNQ7pwYmGhx1iwHEmMXWTALa/NviShXZFd17fsa4sACExLPl18PMF
XU/kZ0e3DtWP6bxVf81x17QhSBwplqiPdPve9EFk1VLUuFw/CKE+mL2p1tlrY52K
Fc9bm/L/o/0V6NbyyFqsOGuLEag4dy87P3+ZboGqmIYU1CCmHeXhznKjvh1YLs+n
t5IJFEQg64hxexz/xKnoPa3d6wbZteWhrZft20tl5imexu25Yu6MtNg9Uf1mrzCU
srQoakNo4vlOKf0dd5x896O2MsQHHtc0ESr/KzlN1kap2T94TFx8MF73UBWTvZMj
bWa3Hit0Oq2yUlnVVjYoWATXm1mcHTTZY7mXczjzmONlvfuu5m+FIjmKgNUNf/W2
ioMKUFO5pWhmMdv1MchrZTApNmarp5MJUSmvBvjFJB/9ZEdUYdazHODBxKkxa0pa
uELINEILUgd7lSFWvoqUhV6c8zyYpVxiDhTcp9rCfpqhN0DOzjl5hkzXntbZi3y5
2xdSVz9H5WTf7MYDLgo+eiitxi1XJzU3IRG6osp065L9Bnjr0QTcKuu86UuuB1SG
VlXVZfppDxfI4EC8Qsc3ft0Bi2QWPZx6heF/OJ54aZwUzjHL/nkFQFS1Bj5S+f8X
Znee+H/4TFTBYWQiE6kQZqjZoZiZ7xPoNKjFsPgnxawdXGgvjGLEmH2ggSyYJC4L
RtW73/P+g/GGmqUUHrWxAIh2l7ogS3PGOe7CX5DnFRBwHZMQub7RQkfPLsms4fe4
pe9inhyXQcJXtkW3VNN9btG9q3fe2DjxLn4fALssVfDV5bjwHFoNlg/auxUWSwRl
/3keEBEMlI8DZ4wodBGV0YVOrON8QxYIg9KrismqZVEJvsulUsQPguqSled5aGCJ
9L+GT8sap9n5cH7DALsZ+481JmK/pEzxkLlvBXycH+I5Jg6tbef9AHwB3Ju46daY
JfC7FwU8fblYpZxSKXGXM8D38HhOxcloTfmVX6rBekzcFIE3EhAr4tDK7drjdsXA
4Qx2oD6T6xD17TB/2RBmMZ5PqXurQNYFx07Jdqm6SoJ1MzBWph/jQRK3IMQTNKMu
G6Vth/iZFAreBiu3qu/mXEfpuAu8G3uDtSjq0tJLXIpvQCBaBSz3fDrJEjWCre/E
jlYnQrCrTvQd5TvqePE4vDKWPBcGsRlTREjPFbov7hLzsEOe6BETeSOwx1Fp1d52
UzNR4Z0vPam9WQZMNa60J03AW+59cU80a6V+vGFLRquKrDiMcl02sEB4CCu76QF6
4mL6ILNcp9Fo+7pSaWzPUVZED2Oc42jFxccsH6yVVIBcuOT94mDNBKGknJZ++I7t
IUT8DFMYenCwCBgIrrc492eMp+EHfTCm5XtuKc7xNuIrC/tdTm101p4HY+gu9f9g
vwNJUk5/7lIfG/afp1W6UirTZX32SJoIMnxe/sGCH3Bqpupe0Sx4rb9E7g80SxG5
k6ciVS8k+HbHyK89c1ytSddPlm668i7cTon+Qn5+qrfKRK1oW4eOy8WtRUZxE90K
1lTprxi3cK5ySNf/Jmx9F1EZRqh89goxtBYSLgt3c9rlGw33YDW1E5iZKh7r9Lxx
1NwgEnsnICEjY56pR0GnPhTEDdLDOHf/qzOfQ5SC2XbUjiJIJFXpDCfzQH8G+Qh+
horINn/QdGznFj7CZRfxShvTrme6wI9VD+cBnx7ZqwlDPNeXro3FUZFXdQVn82nd
1yEnWMJLnplcIfL5h1OADibTdQiNPvSmzeCZPTOY+mKkLIOcciVTk+wxXoUcSSFk
4i/9mw/xSaPFRfSHqywenrKZHVpbo94O8GDBrfcPgW2Vyv17nf/ZqO+AtlEsH8/D
SmLoFZH84FXWC/mj9Jh/rMZ/CuOJpS9TBtUcs4atniebOJyNdxCc5Sm5IFXFOd2l
nmw7xAdKoc839IuS26XNzFQsAuWO2ZJpf9b7aCRTvU7UrNDqLIUGp+/JMZhJNXYh
KMPSjkjvWiGC8JgZP3Yqkt49jUoxniqvUM1It/lhlrVZ1nIDGqdDn2BH80gD/Otm
h6ivqV4XhL8T3jTPLwIkHDjmsQQJBuQHd4hgb7U9ZvG06OA4r54tIcHXXRJ62Hr/
yOCl6KG4WRDsGkyP5vGxsnZLnGaKLDmZmjt0+f/SInDsPhm+4bS41gQcxVGh+s0u
mdlJj/9r8Vd7auq1vWG7yiJUuY4vCuN9HwP1VvRwkTAOhWzVxXBLiHxiTCplgu1z
A1eAnQsSHPPZNS2QNmJ203yMWjTVkF2Qg9gKT9uoOEnqGftRr+Js5bxYjzDXVdAD
rM80rFf/JvQGUESxfdFE/DGhNxxO9QGOOlK4dvndI4vWGTgnQlScNAO+AUkvQ4Vq
fEZR1QmINglCdm3e3WA8u0eLfZPlQzOtWRo0vHZX3U9Ea1xREs229NpxuI1TOanA
uVYH6yGuLiNsJGmIV70VVD08HW7HpJqEU0PrCvtK+eiuZm9AbFwr4LrK6RbANYfi
sB+rYk6uZ7hQ7Ik7DulpQwJYpvjtkIvTjY1ByglgvTFul9750RgKRYSqH9gkwzwu
Kv+uMWToSrBojuBzm50rVF9P0W91U990ku/804B9E0ENwJy3dtcH2h/8BY6257NN
ilbTe6NGzB2SNzgNKP6fIDZmNF5/jOhWfBllcqgb0ibDPyeSF1gLU2gAevflvn7b
S3U8U7SFCYpyMScdJMIQGNrmc8f46XHF5zUoEAfLRJHnM6SvvfE5wwkSsY4HUKnP
VmPwI2/l+JxfKdqAT0e1+euTRVLoRdQwtiHVnvB39Goa6cXEyzxJfJI3foL1y4Wk
zBpC6Cs4/HQA8ocfiMHoJ/RypLAfkOKA0qC++77pBwsRdVOO5vL1BWacztbJuwgW
Cq/6L7UnP+OgrNYX//Xd52H9zrevkKRYtO1977S7smqmEDmP+7W3qEspv8FbTXrZ
A0BxSA/vvelOaLegC6ehSsaOF4GWYjNa9DzytFw09d4p4xi0Y7fgwAgDhOwgGUmM
WleTXJBxlt1Gv2EBbOOAjmTbmiJ8dtmkBEVtEf9Ow4/QrAPOK2BFpDX9hkoK45dh
FpWR4DjNNjxJFPr1byYlUWkXWHbwLzWEGZBNSgvdCIKaZ+dncsp1eshIc1+npu1H
Z0jCdojlEUQhrfcpkh08MwFuHAeBfxOzvr2FwJgsyvAwvPFFSmhgwSIH4r52sSw4
GN+IxJ+3QhxKoUWc95Kr6OUpB8uU5UI/68TBCL/F6nNyCr92T4pP3OwoguwwnodS
gedQRNtN8BGbLwi1IP7pl14M7dxg/5fCHAQHpRBSISzHXGjZd5ddS8HdzmVADLqt
RiPDArszv1IsVStwLqhhczkTW7LO+jFIcltZvrfyVhqo9FYqtDylyWlEh8bz2xE7
17shkjD9lQjR4yTa7L7anLC3VhTMd77XP4mzvN1VOcpCWJ3zjQl7lSZVsZmrFra8
JwYCngdzVK3lSb+NskJcK0jYBYeBppqlHo0l5z7ATBvPV8bSPcXY0fVNDvfg/L5o
29PPSuD1S18EfWU+jzYr77LOG/7l2OuyRzfxkU7TG95sVLMXDSmwypzP1GyQbyXa
SHLBz7988/Z27teCVQgB/UUuA4rUTJxsz9LHMRL4R+1xAEVBdKWZoQ7aVZ9IXXAF
NaZMraHfzisOx3pFxp6iVqLoAgDGDQcc4ExlmoxJGM+++8SdXCwELFmfVLPIHpm+
UWTUlHd9UeX1PO39774URZNTBPNAjCQ8B08BaS35wRa+h7Cn6oNgf0ky2NUE5O75
zGiVQ3vyg6M1NvTACNZh2oJfY7ayV+CnX+uK/V1SczvzeHEI1cLco/rReDIK3X+g
iFXvn3LOL27sP4KIV4SxJ9EI42DIRW90WNXffF7EV1DCb/qmOJO0EYJrPyYrcXeS
pSqTnl+x9khc7S7R8BZ/xDWkyHngbtvSZ23rI5Zh3NMompQmXXwlzi3U0eLEy0j3
1T8Fsy8LzkOLJHq8el+vd2YbVpdYa8UOiYfn/sa+8KAbVoVZ3v44c/+gv9sDgBNJ
SsSSQYnV7witPVMFc8lKShbm9EqlD7W9DZEoCS6lIP60y5+VPKTDm9+RF32NAlN5
C33RJEj8dy43SJ/62OW63cM0Cm5kMwuu+zF7NTWza49OHUbjVMexancNkUN8jXr3
babw+NOHsvBHdYQOecVPW8/eVqs3jBs6P1M67C1cYW4tX/B4LXJY2ciGTMmwANPc
0DKJ0Lo2p2cM54Dsq3fU8tOHGx2cjQJXe2lzEr9gmSEvmPI+TGJDsJrN/5ThvmPS
ChZKjA6AkAKNljDoyrvIKzgcUJWwHRF7bKpS/Xs7c2MpEAkkXXmIHTvEXZ/6amnx
nY0idKaTb8/VqCgqQ/sbPCvzM3gVR7eYYmkDT09AF/SPjFEcfvdD4ndEhZrDJs6V
bqy+4WEJivTZj/MmdK7ztxVzJLTQP2QLzdnKJDf5+boPvjE4vqZ+rjgq+ZzSW/ON
i5BXPumKApAomlV731yQmhLpZ74NYJe4lGy+WUgeeLh6zL89quVxAQDxglMNk/DT
X3f5fSe/+KvjVdfpGDPiqQ3bYVstasYD6VjURl2NBIBdSjELKiRu6v7uhXvo9eLL
geTPzi0GFl1Of4vAWCC/AxjajaXH7p//4ZRArBrvWDnoUjmBiHYERTaYj/uu2tlv
/QjqpaOaDKsRs3JziNEC7KbUUbN92bO+F/7BsXsggeJ2TnBcKsxoP6gq5+0PiMD4
1358qQ9dtjWR6f+az8u8NWkxmoQSFwif8RONspnAj8oQ6vF592pqtTCZaWub+Nna
l7laft/d2yYYVE2F5Ydt4WQcOcENe+L/9wLPz289oBQyupDxQZCxzUNj9wfikoLg
Qb3Gch56tA0Vv+rfM8aD8eaVdqcvnAAONBHiNe1KhjfYUBfqn7wzLOK7b4KzKaRR
Q5eS/TubY+U4/wZJEL7zSjmP8GIgTfBFnQ3GkPMnoulhZpatM16cHxPwrZZA0yd9
7sZLejlsDZXDUDOEBB6YmdMW/Cakk6Us9ugrA03liqz4nKzCr8d7KLsUhXzJTfxm
yZ9vR9w4mR2/jjYmGlhKBQN/8lYmRdNldNIznJ2bzQe5GjsfJOhMjSoYDKE2DugP
J/jYqDdGfd6qhL9eY+84IyWH01hA4Kpgqr9Gx1Bkhp58e4Z5tBqYNg/S6v4wJQzS
A+qiKhwH5pYTK4+1rkX4tJ3TioPj6VMx5nVsLMb+RDtjms8o6O151pw1t+qdkeTB
Cfl5IC3WgaDP5StrSgg++CSMoKKT48xjG5rhqVZ6CDel9kiKJb8TmnQHRqGpKUr8
CCH6OzJsNQSOMop2Axi03Sw9S4nhn5ORRiSz3CoVQVUTGE3W+2HXWLUGA9Umwl5n
kyOgR8gPf7hQOIc2Tkjs8XzPkMcilRgEak6h9sSFJjlSZYx842NuBFbfQJaXCzPq
odDWYWNh7EL2Ine8VVJ/lcih5umu/Ev1g3xSFPs0SjNBlzMGSGHMKXqLpMqw+/Qf
IhvFugXpkCeLyzDDYhhOP3ourp5URGgYh8r7BRF/MXTDwONGOf7l4AZZ9rCYruA1
U+U8s7i1W4+L/e1LS37ZnwhBXx5bX2GCa0Uo2AmWuj2GQ7+zZhC1cNyEEeXD6VTE
VBD1pl6XmfMVxJl9S8GbyR8/TqV1onLiNMXcXO5RZ15cXUK/EFaXUalI0ZWLzlyZ
kh+aY7Wsn8kSZFUTz07cKq6FEqkiYeSVROYWIjC0xRoYWLSuvfeu3dVS4Q3GQYFV
R1q9YNmVQJgFNtOVmHprJ9gkf270pyz6QGuceXBI/57okWlVWRaCd4fPK7TnXavQ
a2fhYgTiOwdUU2ocfg2QDWxwgNApcIZLmviUCMIWLGvKwnTX2H34ogkNfuGlzYLd
f951yTJ+sN2Pjv5fEp2D7BqTMDlqZaxfUV4bC83vBDYGgFqmERIprgtWgYY06R0b
/rWqqW3AQasX2HOexA1/J1jE96amP0UowDXH6EJBTh/D2FKIOhr+Ji2XDdCRzOC3
feHhLhUyL5D/7hqu7HqV43v8kmmKCMrTMK2/TkE67l3shTxLqCNush4/+6F2Dzdu
JTsXEAirSluVdMw1RudiX+1XyeJn9ZylUhn13KXvPM6lQCRM1Dpv9dLO3Se49m8P
Q27F6HO9LMgfJV5bkebUV9N3+qPZF3YqPaLSudREjXKrpXDTy6YRobiWCtnFKHeo
FdluPDtRiTZV2+6w+jv+jzFMz3KM2qKUHuwZ+NrWn1Nica17CX5xsbuusOmkbUg+
vQml91T2kBSi1wpSmNma7x7OUjXvlXK9tZeaceKSnYY7sxv04RkadeB1yozkxstL
g/GAlcuAzJHbx7BEoHz3ukb4wEpEn+KcH9rufOwK63uRik0XSnC9RWtVRKOZNr7A
CGZx+FAZk25yqDLHo27OHT3v3ZzIJ8I25JwyQkD1sQpXkY03GARxB9/UJCUzSimm
RH1SvOdVgxFVYZfPM+oOTl8xtPRxVx3w1XeTcGq171eUGy+OsXBLIdS2wtgbwloE
1bQjJOIE1ljmeqRPv+QyDDquAK0z1sO0BYRAXK1LAndn5eeIIHmUP5KUWf1VUVmz
tZn/PDf39LlqC9E3N0LZX13HyT7PnDlZfH+BTHEgmplWrAhSBMIAcozvruqAAd0P
3YfChSrrgxIatSt9SSK+MM2OjloyBUTh+/Q8AKpnqCgJdPTg+Lf+gfCBXgerfVcg
+yvTqj1svLlMiDn/cwP3OIkt5uvaJg2IUrgTcROcZr3DbrmT1Tbb4H41ABE0KaBg
nWVi7cSKijjf67ll/R7o8KIAxjMg9vfwZC60Lp/KAO5qgDxuFjSIzBmGoBOntzdw
enYqktqwkkQ8IUQf14za76Mt8PO0DDVTVr5t+k+YLUm7qdRWES71LzV5wRLwQ4WS
i0dCNJdPUUsdExRXcPYqHYdT/dCnWuV7TPMSHfbb0OH3f8bGYp7fdwTwrkRFBhsW
7sqDLEM6eJ4Cx/W3V6kmzyx6QdL+bqrzrxOgFF5KV3nPaQrD9+T6/0CSc9/nc7ce
T8h7/iNRdNRpp9lTnoxz4sR8xlpEYErV2zapDv/q/2tFvtnAlnbgfzUWa1kgp88m
/J0p6AXBtycu1r99P9lnIQwPWT+jI+nnWtX3cyr6QMxlhgaGopapukZogstJoV9P
DoHdNvvzUDWvAEwBg92wSpl0bHLJeKw0cUY5E1o0mkYBO0uQc17RqePhKWMv9uBh
XNOdQ2zs2yX1bwvf+dV0Bw4E2WFB0j1ZiBU5pKdDKhJIiY43zVOHymvzXzELJhZP
5V8jtxQkNPGBE1RJSLV4Ivilf9mdoOCPGJ6nRmuiCTbYNzrhqmUIYZou/EzxCk7Q
hHF6t3ZQIvtQuOki7V844yBKVf4UTTaIk6mZ03c1GpPm/pCRClACgA3v0xFY0NrS
S1Cb5DjDEZoY1+8AYh1hBQ0Y3QkZuMwfLEt3rOzBjQRXJnbwVLvAgOIOtIojxteJ
bslNvMuKhjCNVnCc+srEi7+gxLHtDdPWjtdoRHDnJiBjm+AVhA1iCUB5djBgAK/o
f0wqDNTauuXhEhDrcLRFT+h2rTZQANovwGcBDzTeWjVUT9SDxVuy9urBVLg45Ugp
bqoyw+eNtlBozcnusSAQgesY/mEJ1p2MXT5juXnL1FVNYskqMyKG9doYp1vWBtWn
WN4eDZG5gjegErIelqtQwMjaq8Do+eGd/N7FT2ARMtRydytiERQBhG8IKwoMvLiY
5OQVh9LyU6VWN7W7l2kS/i6GmhHLKCrsZ9z070ubIpU/zMZcu2fN0dn5+F5lzqYz
fF+p+d54ovcglxNqi4IB/WvS1QhOsDodVxWzAC1+K5C4QZztBs4kmWkObJGozdfK
xjYl6klLlzpYSr5QJO9spTXHPENR/fv7XWKy5d60IDwoffASe1QHENVIHajCEOV3
wMXiVqSr4RPr4MEOM8OsihTdO387NnoazYMM1Ay3Z1XKB0sUfQJnhUY0gvTukm6S
GWIBSrBDCkL6PapYjO9fqkcdly6y0iMcdDrHaOZ6Bld2j35dEb6qK50fIfwMIchV
fyFjVrPTK5GMkIFiyYF+4Ux2VI2mNUaBbIX34Ahr50duqr/lmGu8oGpMK8lE9Uix
JWFaTrAXh9+05kYZ9+JTbtbyjnkgBtuJk37YEzUOyFUe5BL4VXqYhA2w3zNSv6T/
V7UMImSbaKO0ucvrJJUXMLW/sRlNiu/cSjMuYDS+sxO2mhCHUrMu/poKq/vQoH9y
zZOlCQxYNZ+YFfdp1D6i2U6EQerMN2XIcls1rjJrW56gxEAVyfcHEU8/33CwecZG
5bN6H2evRSkZNPrGwrUYw4tg5U2Mm5555ngz2VN2+o6u+hub0b6QpHtrb4e9/EId
jWfSMGvU2U/VS0ubmgCvLiF7ep1Vn10zsXS2aHbK6jqQ4yxAUhjCyFUH/m5vwSe7
DKATp1v3Frfo0vUEA5/+WUjbRO3y1y+dCVUCvtlS9Um57UF1rkl1l7l49vokQaZX
l5epcDOCrTwNpE1kYLXjrQij47tCZ3iT6iF050o6fEGHOt41uOOzF2CfZPV4dmiM
EgPZrAC/s8oZOwA+Hh9GV29iwBt0Ide+VKDkQs8Tk2wXaEv/k1iQpIIasczP24pk
hbykJCwZNDTq8WtXyGFWlFD4qkMuYAumJXfOwTehSbhhnSD1ddTwGA74y/PyU/is
tsDsfj+cPCL7/B3SC8E65szWeYwwIJqDB7Fdh5SHnSLjonc0JZxMZ3txIBXfZxJw
c0aS0lnsF9VnugUeV52a8WxsRa/G82+6hIf33EAIbXWcPW4uFDYWrzMso7+EN9uE
koP5/LOTnW9kimELfFFHZq76vja64qEzTDegcUcuuVkAObvoZliYqPHIQQ9sljPr
AqHdkqWKBgXJIToMggjyVggeTLmu4wkvwy7mx+oIjuGRUWOzXGX6O0oo5Yc1jAvz
rjuASqNpbvO/9x0Xx07M3dG0df8SgZXzIBGodVKEolvkzBVOdpsoBfsoSgWTLSyK
EbPB0cKwlFj+9lqaToFkFMrcCq3J4zchPAtA7eGZfhl0fFpW+PVc6pI9cmflfNXb
onX+72rQtkkX7qNiM2a4DGTK4qEcAswy3WnqyGf3hvk0eoWaURaBjAFOtQERdZbb
eIzIIIfK/Eh7tW1E4rCPcNmvnPKh4n22WYor3LcR+xYe94OPSSQgzJhnUNBgcIJe
EldgAl8Bw43UzQK39U/7z1YVdTShV2PiJzuGulW3ec3AnfaAA9i2fHZzu2ueLUUw
bbnSx7TSxvjwmc0sICUJHRt9dR6vHs2gltjTjwv+8adpYWQAYJ83YwKeslYY7fJw
jQ4stX4EO2mJWAUCp2+dmYFP/+FmT71UbZKH+GrNAPLnz/lbmOv+FVyuWklT2RoX
0kPHzXaAnUiubd2uUwyCogfHO8vMkiFbEhTyYRX+LHyJ1k180yZ9MJ1rqZn4LlYm
FzT9pt3JmPtCT12dtNi0eie8kJf+Cnj4XLCI7gjjwn7h4geKmVrPaa+TvCLx+8ud
cVXCKHCm82jtsEaWAOWhDGzGXJ7Ka/WbpEPwGCmiMl61lS4Fbrfzvl6gIE+b6m4h
mAZNTXVIMpSW3gPsgxX+y1N3yo9IvyGZ1d7EvU9UwvO3Vemy9XJqFjlEbFX87+re
XMcJ5sVXgo6ZF2obV4cD6qU+6o1IhCv1dpotoecVJ7j5N5RPDRQkw/RhBGNgnHpL
Yzu1BWI+JVKO42lFH3yf3ZzGyEggK3ul5jOOAU/8oUf22OCPvi1ixRnAzwSGzcFn
2QYT3X7So7qkXHPwR9EiXU/vuUzVQbSULrL8vWqwxUwJ4pKCUfbCGY5xcKCtw0YW
n2R1th6ATZPKZDlCo9cRIAwKNx2UJsQyXc3Jd6aeLdNt9RDb1utgU2KWXgJ0TkW0
KLd+HCjWzRLdXjZEEu5CGwj1Fe/rwboDRQcm/O13IP6ZAc1Y1h26YX7vFYUJUjYg
Bix03XIKx+5FyET8Ou2NUWwuO3C04lqaVuF/RVMNWwXvgZsyacRCcyl9ifIGqrLp
JQ0lWgTqWTWnUN5fNxnNr2wIQ74Kt1OZvc7v5gvK89GJZ9o2ofIQWLiGX8nbCPHb
wp0tC1eWQjFbMTuMZ1oJSdgsRkOvaY3X8lAZduLsWQM0wSX4t1IFUbb+b75t5bYz
dG3w4nbeFM37temCXOshDewD/7bsxskynQC9zcM1nLTSbDghEMjY3f8QkvSu4UI3
ZgMgZeumAmzXBCo3L2WloDR7kp/HnbqzdQm21dNfW9Z84krMZI9lacN9ecNgAwtf
YyMpWEMpqY4Fhtibj2dnyuZiO1+bGHGZ+q7W9XdFAm6twXGHNOis8DD0R807kosj
f/L02yWBlesUZktjVmC5tuzkaxjJTX0Mr3+tSM8cCqmD64OlWrc8GbywHr7Mv+UB
tULqf58j9MtnQVXe3G1ry9qyv8yn72NdSTWaw3709G73i3FurfnVaUf/qs4BEAY+
PZgPH4k0Gc52GKFe4XJPI8F0L6A3fAjeDKKl7XY4CK6bHTmmlGUui6k0pGshBp1f
XvRbF/OvjTUr7k6Q/WcB7y0qnExsTqT7Pz6T/idbDWjXClk2i31lGfdNiyQd6rPZ
g9+gXHBxTd5OrhbO/AFKYgmFk+GH549Z0PNlPSYfktkbdjfWeKIcRua1i29DqwwY
ZyWBfimQ4Webu8puDHZU0c2iPGLTY8RL/ZGot2Rjj/opqIRjG5/0PZchAAoy5e1X
tK/xtkLoMjl8TvYlQW9KNnYlB14L8GHdwEyMWV58lnRXXvS6kcESc8PoNrJVJas0
jnia5UA11qB0TNdKx+cmIZ4Im4mger2gTG8bYkbu/GfwzMgLetbiURyHCdZRH5kw
9eqXENmcSEfQyyDm/l4Gd+/PhC7WdyWgB0EE5bmV4iIguIIhMi2TBR6ZQgBMTZ7j
JSFcuEGMbrzHZuwwU0CrCjvUr++1TByLcY+yFH9vamf7dW8B8B/T5789Hkal45Us
aXu0Y0ORO4eqvy6rmaU+/DjLJ0LZHTDFiMXVZCFxz0cS2tB9r/VeL6BGiVfTNPeb
5Pf5DVLLCT8OQ1MC5yOiRT/i6w4dlMtW9qY73b3MEicI1n03LJIiAT5E1RxH1aFX
Ek1zMQozUw67vqqE+bLbux9/Gu0d6I9SJkLcYbDtDpnmG4EJs/BvZPWIfGY0h5nZ
BmEIEiTh5bIraoNpNNKfvHZy1q0pxFiFO/MDxq2tkx9yIl59cuBfi/t09KGUFw39
UunHXZSB6A9brWwVVjFhflhj700o5/I35ZOwzt398OYNZ3gxlEOjJevm3RrIvAWl
kUqZZdaby+w7LoNn5qZocYgtH79Anmbkuyk+bkfhEDdKhXFG17bxx/C7xzWHcsJ3
0XiJg5QOGuq0rHX2UiulI724R+1w1ZzQHxXIMjNe2Nw/USSwDArtp0sfPN16DKbI
0cWIcINwkkBfF826ZSAwaSYL4YuCPXndgFsqZWlZKyw60US6gskj9/m0BDCRVLB7
4hlguim4ZFk3J6pJd0IRIMsQzmOwtbcD7agIsn7Brz9Ap1z1w4vi3U4HuQTnDqUR
4bvN7k34xHXmVQiAqPYBf7K9uQI+aqyA1igIbBf7a9reY7x8iR4RORgQuEXhDdqB
qRWwO6sQBAigZ8cQcxWN8yLcPQu3iJ9AfRs/JardxYDEQ0uWKIe0UeWtXF7GfZxE
mg1pHXitZv6pLNqFlJCbLxnB0/W3ytCRIK0DUryLnINhNSYqCZUVfNf37ub9Kk/V
qELrT3sVtfEJDd9RSpTNxg8Upptg+D9QvZZmnW7O0ZY+iKQeggyQrW0Yw/47DWHz
YBE7HSbCgGeYXDiw9WWtTYvqZOpB6oiJ76KFEvZHBOM0OBMmU/Tv0qAqL79YxS3B
wFj9UYZRSjrKSB/gQKLuHmC7eyxyRiVdjI+rzmO3O8uvKhvc61GLsx61tVI0Fvr2
X7eqVN23XSZH5gl6KBairc/IqiKIsnJIAahD7pGF9fRQad5B6MSe2GOsiH4n21E9
j4YtLywMHSRNIKXIGaP1HDGxt83U5RlcZy+f/V9w7UKyh0fc2zFQ83uLOb3AvhwP
td7A+dTSbamL2BngEgOq45MkXFTC4iY5AfZi1KCRM0gvHUGWfNx1JKXEIyWMaEmu
W3BhCm5P7uxIJP8SscKmUI6IOj84BGiYrF2bDoIFr24V9V+wLX/zDK9v+tVI4Ysr
xffF3hJiAX16M7ygK1PMM8aHQR7QXbgWpRbeI9K0H0RcSOISIDRqmp59/hKEydaw
FdBx4gHPgbZYOHwMbyPiPWQrKOtGbxN4IdAaKYl2VpwmU7P6Mmx8bTICMdo4qNsN
9nPoPrR9n9tvwo08qtXfDZtq3smwOIoOOw+agRSY0GTzdRSTphNw9XTFLNP8/OAX
M8EAY0gcBI/F4M+erB4NzuX/TqgCK8NbSqx4ytnEQ9Ci8l4rW698v4nEj9L19XxV
JLboVoFD39tebhMdMHihizu+PhVIXsI5V8waWmIdtcoeKfnthkGxg85q3aiuhCpg
PuyWb6Dk2RvWBmHEjzbGWnoZZ6t50tWIfh6KjHqsm/NODUeUdDhTD1nVAT2F3U8E
t/r/tXWoNJRIzEJf4D4crznzxda0vJ3L1g447rEKm66qUcz4oLm5AT/Hhmprr5cM
CaHN53cZSKQIUvPNHwhTW0TEinL3rNeAjQIWktmFCNQWtIW2YqLRsDd9QtFS/5k8
S/Us1hWLdb0oycvkZDDJisdLsfoaEBfs2KSiQYmfQAB46K93/XRcvhL1voXSqHJ4
lfsGxqtg5q6dNQ166g+FvJ5U4GyFYFJ74/lJuI+sWeiFB2yV5Kft7QrwrtkvNPEO
ay2lG0ilPXvUok1Z/aV2ZTjqmG9TmaE8rkC0wxy9vFdsD9bTyP8R7KDKKbglCN8A
H+myjaXuAom7gKo4mKYoz5Ch0reyuNqo5zLL6J5m8nvbNsRXCnNfTPOguLzwhuOl
vFmoNCpzb/VztrVcIMluCSXKgp3K0ieUOBaHpugDr0FhKRIclDlrQeoCzA8LiZOV
QGzribJjiCQAfL3WSctH3ckyM7Q8v0GeXWmbYCGx5B0Tc1wMoVKMw8BrcG36KY5w
hXv5T1quIrwiuaREM6fDoBAmyx5QxvEkb2M1WRZO6rBGD/JFCROC8rpHRnEZJ5EL
KlgDl5M0/0PhMqj39nHClFotTzHGaoae+AQaeCAn/hgYXcfKXjFXroDTsNByBb4c
1wZWafuvkGTI33G3JHQVKNSgLYCKLAUFtZLaM71RMVJ7Ak9RkuXMV8/WMkdS/uC5
TG25qCJ+k18mTaF78iv+qn9ZFxdy+25A+cXtTtu3XXE0Q/fAj78c05g17k7vAOJQ
04cJBx4cWrDg6J+zyCzq3zzj28isuHKN13CmLdEwov/z9i3AotkFgeP0N55LeEvQ
3yF/pxPJyJVVNouQemQocmypqFtRfp8tu4nY/OtIEruBqh8fDNZWUKzvzTewg0xC
3zZM25NjEo17RVlQ1EO1f4xN+jNtxWr5/hv1svn+cXxldrq1Ogp/X0e09Lh9ymop
rNlh5Wp1oEHckvNNMvU6y9kId0I0QimKjditzYPamTUTZiSxZytsXizr3iKGJr+Q
y+8WtUH++6FaBlUWg8sCfC+YJ0N6U/tJXtZKq04pVIGV6sEYKb2UEkvGYWqxA1DZ
/O2/Ca/iTJjdJn7wuctMVlJiwA153u+BHhMEUSe1Xbd01EehJ1+8DUcF+zFMCpmy
pT+Pxunq1JkAFTV8nGejLXladiaUXiDcI/jjNLA+bT/uAvhZSG46M23aQoL9rhYN
aYCetEntg4Fw5wvmulpmef13/kx+uYPVz3yfIOnet/ypZbOCNciygGAacpNO89fb
DpBBhUmN79hTSw0paJnaAfganSLojA64LMCKkgq3Cx7TmnAuRKp+hCn5P+QYxcPL
b2mhGI/LxHrpG0kawnp0iLLBbwzz0msruz1NsnlXZQPPVEtEcIeeu4gAjYGwwroT
REdgG/QyWcVg8nbkieobgGb0N8ZAO5FQaciWxjnoibaHGsnKdxBWlBZon2WC3RpM
GBXTz+snehYB/DTe5UqKmYBsXIjENCWxdQo8UOQ+pi/DJSSS5S+6VxZ/3I4JSt6F
7QuUdAfG8YbahC4PkHvQh4yxr/Lj/qe2PlkF805cQi5v9WYzyCFNb6a6mxFQ/Lqm
3NFPztUEQGaWeuE/CMggYtaWmfq8cStS0hoPeS/AFXOPwgkJY29ojnp/7N17U4v1
0ARF36OKREGxu1d5fG/qWIas2GkEAMKGBjR1pY6Q8M7AaUppvuJ5sDZS6hRKEKg3
BkXYcR5ebFk4+k9K3iSJAsG+6iT52RJFPCIbwR9sXha0qa7Ic6NZojFrG1gbf87V
cn41rKeWW2jh78crlSAMaM+mX5xRYsexmwRekbp3viA7Klt2z+/TxC77tprW/7gU
Znupw5sZd3J2eozK7snJ7CuPrwRzkupUY0lrGjrlR3p9pyWUme+f78NrONj/JBR8
k3DvKR72hz89rs9SknCLfETTj4RNDXVl3nVYN+3PXtXXCD9yxRgPLLlZJtOpAsOv
9s6HtbAV4T4R4Df4JY97tRaVk9szKb09dCOlVpEVPrOMqT65IbwyHWG1MOsdvu59
tfn7BaCNTmfQiiQgTBDx95m0XCRwMt2ccQrV1wSqZf/blg4gP9Dw9JeYUFpXceOn
jhqLbcqqM1aEMuKl8bkhvAOWEhKgU39ASppLSldK/iYroZ1Hk+iSr/R7ufzUM6k9
sBThggisuO6+wH4uurIysW9hmUPj7/d8ozunuPvas5Xk80xB1AaDqjcbUzwEYYCZ
ToSOWNNX1W38tFqHmXg5+iCtZeaaiyvtt+Z3ck0yk48OFl5CYiZkBEWfAULIGiQn
AYWDNirLX5KNY4284LWYpG3yAeFMNeTehTDedzpkqruYoKduEdHo9rvw3n5JrzRa
AqrJzavHjLsmYGHxWJv/IYqnSKnde04yr84gankthh5Hc6qvM0k7mH8yVdGUwiMt
Kc8e2KTkykYM8eGypPf7yRYcm14Qjet0yDFupfsJLGILCTG1ZyNUvaBOYSZAJzfd
hr55/Lg2Kt7Ky5X4iVfMvdIs67qI3JKD8qQP8jGIiM2r1KdZh1H1WoibRl8XwktF
wAyqQw7SctRRHLT4e7GVqNmyWHUjzP/eON+ZANcJPgZHPYPUUnzsyGfmMu+aJFsh
tFmsS4s1O7jfztQYVFGaQNdSsnsRjRFZikmwQ5lGIyXXYW2duBUceSyQDTL0zDBB
JGsvNvDh5EO8F/B8l7FCHhYgPMRWE0gXe8WKK7g/+cXvE2IHx8aFVrHQK+ZR+dho
jHWbJikJQYyhw5/dMXCbdGW0xVGHYtSDZwt0YXk1fZwchfHZzNWO6JSG/Gx372jc
N7Ol6uktkC97h4aIdm42tbv72S4sj4aNIY6y5hV5ytpNp+7EqudI9zk2zh+AnBpX
Ga3/Sdb0EBS9BDtAyWb8zk0hEdbU+t99lXo1BaIst0ZPxdanBNudN6VYWkHVlEtD
jnNJ5x+PYhQI/B3K7HQ0GtFpkT93dp5qs3NiML+u2g2kVVcd9deNWWsiv5cBRPs+
M35okcFzwD8hxM3QQV6Jf6TtVIeeWRZpx00RKH7yg1Hz2/RpnNcL2MWud4nCzf4h
vO2LDN37gbnjyneJZWXN0f1P+7NmkYPitqBm9NKdi+EKlQbVjYHEUEMDmP9Z/HVf
MXyYXpHBIsG3Me617u9iIh40iWqw90Z+XHoh5xGXCpw80jZiFm+m//pW7QnKHGIZ
+ieHZHTKnvtwwlry+a4CAxlqO39IQP3D2SfUAxs6NAjPPisLQJfGHDWZy8xQjnKP
cSh4OWSBZnaoMoTMAR+ACuHe2Sx32tzUVqHiXXYg7HM4qu8JIPXn/IXZF2eEV18K
yBpESQKyNyvz9CX+OCnLq5CSnUXNaTk0QtdfMmmwPskXFMxMrjY8/SXyEYx/ml/k
BMnC5utqw6fdTaD3jnnLbDZXvXlUsyOt4AAetGExyVhUQp9DPgFpbGY0B/TQS95X
ISlTE0HYIfW4F/52UaWNaTWqimMsY43VjaLBsSLd7aSB2TQsb/0Y2tN0zJjSZW/N
TMFHeUKhWnGCjzfz7Qfk1FwXtsP1xcFqBVY5bcWHBcuFNLXQiRBe1qG4Z0pCwytH
TcqgRtyXI9luxZ93+bGIkJ0lvP0ht3eSy0HnMMP5jGbiUrOAp+o5FyQq4PsZsM9L
jM1mcY4IyvJAqsYb9+4p1d72U6N9ac4UrW6cmYsfcnG11ikuIOXr8JxXw+POrWP1
5N4HHw/bdnt8GpwiHievyvVfQtkbSBhcMMGxWFgrNjKwBJsZFwTKfLNzUOU1ZGvA
ljfrK674poMCMcFhKhBVOtz7387TIPgxuvl5qnds5+AAZDi4PtpbgSGffTuh0D2E
FxyOJe0cvwhQaBue5J+GEz/c02fIab9N/9f6N25sWju4TIC8T6UwJTmFaLTte4Dn
hnE3Iama7s6HvKPtX2DtEwzvuAIEyKKnekwTkKXRuOoc7ae4c1ZwCylWtDM6m05V
Ad6jRA6gkqnvvM2HPdyoSzArvSiBna5m0lcoLoc6ikJoaRPEcbI1uX+VKKdRujxf
8OxgZDFqn1ZfFqprVGynFdxvqHy51ZcHFPfeGxs4hKNZtZw1m+ZV4Axx8wIt0Uh3
/X2sgJ6AylqkivpEemJLuHrljS9hGS5rsLpDl/BZyq6aZ8CmaHHdJzno3UJHbwG7
B/FD+uN1ABZ7ZCYxPzRseBzbPQrR00B0LeWrWt7GxZdN3e0uUpwKGaaDz5DDktYS
YpJohPA4ifY0EA9aqfuy08Gfk0HKH+2TlhFlrjJ0huXfOtUc66sJirg00XSEp6uv
D4TL08XxtpJsflu1V4oXElxVTm+EhM+UtyOAVumiog2O+CBamrjgs2kCoC8IiNaR
jrhgtr63zVPr53xw3Mchqwi3YqDI4Yfiw4NN01xoO/xTzbpBZZs9kT+oUgRKfbaw
t6GkVG7SzAtpkBmQon1srjRiScRDSBxKQh03AWwMdbd/zVonFne7xqgJjqUiKm/B
UCiGfadzghqtnpBPYTOMsqe6hRAGz4PSoQAGfmGaNcPQhXA7bC0YqRNGdJ6N+k6D
AzWfD8QZNFSRPeCY6UXiIjQd3XvVVFO5U9e4H/BhAYuxq4lgOhaSz5byP6z061Y1
G+HM7CUQppWZR/dfWAdnsOLUhrwubJGswspvz4ibjSGZsYqFqCnD3izvE/WUKghA
CFpRYzoihtBy+Xgd2EsAjxrNCzYtUKFwaiUxF2T80XYjr35sQHPlxehI6JTrtrn6
f+8YGtcrIGGR5fmKRzBtxkmojalHip1J7A8niCWgGpL6+Sa22bT7RWJWYW5jfQvy
sM8hGsBYKvz2vSqopMqudB4fQJn8Rwx5218WQbY3DLGmdLQk096sp80qjyH98YkA
fUQxMZ3gHx5EopXpLNYUWlgOUl0uuy94RCCJZa8yKzBNTqDo4GhHFXjg8uS7ZAxs
7xWQaQLCworPU9rDG5SZeoCM1ybzM0CRzGKMBT/BBOEEFGsX7Tabp3xZ1piq0aGo
eQq6JQYWkv8iCoIya7azDAnT6HYFOJLOrTiFJe+oczj3YN+qwOqGbDZZcKe0ukz+
WAsKdG40bAN1+dPtEiUGm1gLxpub75z4U+dgnhl9s3eWxw7bG2cSt8P3Z2el419r
SYHSZcjA56OHzD1q/iP0AkjUb+uPea5J9vanXki37rzbGc9jHY+7v6BE1vwq8NcX
Dpk8+aAjprs/1232IEACCHx+ovfIcvDcdcRg99OIHZlOWWs7ujDRfjGGnKbeJEh+
IKCiYOITXd34pDfWpjcQWGgRYnPeSQCZL7bJCjdJKNqcdUtrcrodFyiS8nkQVc4j
ywIIQL7KlJqxC2/1UymAkueEOoh+FFIjjSHS8rV/GqeIwGGJfRq9t/U8ED5emaBI
sCnEm8m1IahhRRqvz0d1HRS9uXaCfRvC2/EekwdX8KqjQOcsoSL9EIgygeyDG92j
qfG7Ju5bGDek8IUQuxq7EozX8lbL5NnT94VuOFGcY76alKQj17ZJ6kqkRn9E37P/
oddeciZxAtiwCZj0/L1pFkob12EViLZHNMM9xN9fFU+wEM+Blr7ue34hnhgt7neo
Mnbo/rlQSlFD8ulEHDQSRo0FUYGZkVI9PnsrfUJxEHi68ZHW4W0EK7DteiEDpqVE
5ahaVpDfoQ3s58pKvwHChg3LvP0XbqJOoQTZoh91dAToO6DM48DVrzT97KrJRwG3
Mbw3d5Qyu7uVhOdmZvcY3gs71i3rqF0+tFiDeNquRK250N+9dBUHTcTIG0Qk1KMB
4ri95wF7rbeyb5crfgpNYsokHyr6Gav5b7McoI2dgW/PY7vzLjRp2c8d68/BCGfg
OmhvbVwnPm2N0WmL5GaaN7rPRioLKABNVyNr6tkMsHRyUwPHMwQALnvAeeXw3Qsw
roHBSf/IH0pJuwv+5u7E2Q12Nmpc3pcXPfTVE1BjxofUMG3yDoKsoK/8GVWS8rFI
QFWIh03xYgpJsfs9geVAQOBQdLBqtLFAGFM9PVpdRYrERZCqeEos0aY24QgSyekI
dBt5NNFJR1IFVECgzycKyr+AkbQIHiYU05l9Hx+l4dEAgWQivFHngkFJrwApzO/g
bowgxnNk4z+/IfpZfPfq3VOriVYek3AzELdsClSA8j77Vd5IUOazc+rOAXBQVjAn
fay2ivZozqfC4NxDl7Ap11h/1MzxDkGNuOOon/SmWxr5tZpoVXJ+fOMjtGtZAE9b
DGa8VYG7IZyLgE5iw3HZsDevBVIU2UvhH2bFrkCNk4RZS1V4+VYr6n0aeOahuHde
P7N3Kd+Gb5Qat7HmbJBNNuNsYPHqhvXZIDwrhruCODcVALD3ctm7yXpwvWVKiEKd
2U7d2BwctkGBVPpS1xyOOafwTyWA3aeEw0A2HBoROnK/jWZvLigxxb5gn5dyVhG2
xegIdSxZzUtuoMRryDnYg0X6n2mNgx0URNZyrsJI0HMITwhMcYUw7zmejTlBqtor
sEyhCeXOS5AceDjVDDGF+TPNdICDvtKyKJ/10CVYpoMhfkVFqOhcen+vkzzriNK0
1vtHxTOxQdR3rwpN9JZRkwoFB/OZX110/GQjEKDDdGuQBUeszqlEmpHO2jB6EJNW
JNH5tZF7Z2ric5GhHp0KJuhQmd/Bg2HCl0A90r+8TlFVEcA6mR6UvPlT0Oj6W7Xf
p25zSZcCTLbcXGSZpEx0+MyGVV9PK7fhV5Wv0XU5q3J5hoa5ZJmRUhoJpwOnzKpn
OuSo0XUctWM2/ELy1uABiE1i+eJFMUFCUA3//wZw8X04JPra1ZILtZGB7nAPuTWh
NAKmQV46MaWYyDc2Pv7N98/yvs3ZE+eYOndVRaI+nXbQwUq3SCEUi9VC1yuNohFJ
bjYLdUM/Ja7AbSDnbEwKDiYQLYaQI1QBtcG0bAQLhpif9ElBOhymVTdIEsMCFxEg
uCvyDQ9E/uoTNE4eIdO39DbX3H6TUe9fQ7JHCrrg5sf39aa2d2zsmGP1WL3/uEmT
/FmniuCAb/jndcdLM5zIyCV6mXXC5c9QsRqWw7/FG9fMOlGP2dPNn6qQBKnRFv7X
iEY5pjPwoKUG9UnmdwZzGPmIE4YG4mnUrOF83al2SDZ7gYH3u73JlieuyDAT9mKm
nohuHAzC5EEB74o7fe7h9MSbQJ1qU7zNAta3KR+Hdr/CY0hb7NQEdpbQL0OJcF22
EMNWZisrHOqvNx4r+BcrNQW4wZ6Z42HYNKNv5TQBwBtyDh2r70DWv7K4CBI0OXWH
2ALUh/lhTh+pV7+Ks26s2gdV+fbB/fNAkV0ZDlHnutK/KcAKREIy5BPK6VTFL9I9
8jFTk4QPQk33mK3ksv/Ga0XWWwkh3OJMTV2xuyj/m21coSF59MxJRvmYb+/TbVs8
DSY3DbKxaXRgBsk3j1DnLMX3eqj5qu4lILgEH3FxfkAZdWKzS0/hRNchlq4QdXT7
2ed1o+aiAJADdnR1V4DppYwyJAT+i2M9DjFmL7/M/Msqxb8PPiGpIyadaRv9A+oy
LZxgn1sNT9u+cC7W+IdJ3ZWrfos63sbfHBvonHYznoAt9W4OTOpFaEXCBmeJpCoj
PkxQARtYAamru/A7aQ8hLkxtXzvEDyzSo4bq552EdIQBYay9vfv7nVRzmlZx5BFJ
srNpr2znzoIBMhmiY7gAG9zKM4dG6Uvzki8DUJX7I+uOqKUJocGtrRIj0ReUOXSL
FtrVBTrTM0S066JTWzozMdt2JCw3K/DGy/Or92kp2ZptuETzcA+AOy5Feij2BT0w
pG9O51lzOsc9FZ5LDrNjeXfrJL6rSGK6suHIMTk8bV2xWWHuSdKSP4wt3piH3ISV
Q9RBxAlMk5zKsODZoDcJAW6TS7KXAPVH7DfFXPtEO+rnjpKiffhsF6YOdYkW1vGV
GKaxXK23WSjC8KRr4VN1HuZ8Emh4wiJH2AvEpSiudu3CuY56SF2B+19C28imFx+X
fezF2C2nVS+UGj+x6UaBDL18Itfs6iRuCDQzDeg7to5XzoGQSetvi30QcVO4dMW7
TNWvbFP7IbKcMjqGo+c9clnSnFZ4EKelNajxTf99xBwZKuS5+bCBMvIKJN7L0PZA
jyzNFFNAnBv3+pIPCt1a1KFSNyvmyRKF/NNGElHcEToFj0mN2JWLvq8IVzvcxwrg
ToPrKUfOIwytgQfbDVzCRBg1EFavEnU09OHH7q72ZQ3PkPNFv2tEIhGn0avc/fLD
tYbkykQhzg6LBvT0TFetpAh+GwE8f32pQP5A+zUMLtpcntN1/JpIToJ4D6IVt9m7
rGAry4wDibEBYKp/V3myRYR++g7rUT3pZ++2+t+3w2pVs5od8qunrhbnWf6nNDFl
Zf1hvm6F0kC1D5gOY7rjdoB1uV9VC/29Nj4ULrIr4FkkGCErDJkZbq20NZDFhe73
Z6wxm0jaRIThVArtMi0Hzh2wXq2vI5aSvhkngUuZzrsQz5pZUjs73cLyTPL1N7hV
xmqrVw33fGjVXG2B4yxFYJa8IKQzOheoGldlWnuSrwkRzXSFPSn3XeRbFppsZ63M
o/PimSlr04yKmeYfNqvq1KOpLj9oQhENrSazA00VcimxDQjGF9l0bSryYYAIWGhP
Yz5Y2r1gR7vCuxsqLFyzjY+n24gRiaMSHHaMpfg5K1Mclh+0xLTKu97q9wPY3MsV
Bo+pCDAsICKQRqTDyzXOja4u4HtswsdlIk3Pv38ER9YyHShG407yT8pAuta7tIxt
xZR0G+CEk23OG/AwC25FvKtsejdIULMpEe89822w9oIkVJQQsyjWM18nW4E2T585
lK18GMP/YgTNbauLzQ8f8pfTQ1jVFMWwi9duiDbUu7x4oRLS0qIkYGK4uLLbmrEs
IcfxmZVBm9aPcYuKFtf2na5RYZ4T7HDPQNze+aanzFv6oSYvawcExcbW8cVtl+IG
vsszw/yhxcbbe462UbH8spI21qDDtlrAM3NbVqBTfJ6t2SFKgpAtj6kw1RKyipYl
Kxy2hqTNwUAfxlOKs5VSnDnmpoaiztei0XhNhxHVQVQPvmbNwHvAY/wPcqqtybEm
a3JxiOxEb1Y0n0zI8Fd+5CzEVd5aLPozYrwlMSkDLehLjKpO3eXKx/bT9g8f0Jhv
z785y7E09iEx1p7Ig9ZOPsUifxFS6We88rKm0skxxfLR8yTHPFnQiXWSGL/r/Vuw
4n5bcoi5+jnL9mq3Cp73uC/+TvF5kDVsdtwfz8AC502gsOWL92DU00C4amoHig81
FqvPtQ9ddH2mjDoNCGc/IoFrLVpRkqya27CIo8KbQzd9zaDVjibIkDuObUgzVL9l
ems4+FInefAgN+bDpcUe0ZiLvy+Qauq4EoP8fNEcPNzg8ErlOROeN6D4qAdt1bjJ
5D3Yzghsl9dNWh24B+Dbkb/SCmNf+Tb92sxIzFdl+oneQNNd4GZR6DIWHBCBXc+X
F7q7KmdyF/szaeDsqQZYGEPXTlho20hA/nLKyTQ2rcu/bDWnUNI8dqNm2ZjTRNfD
l/KnVm+Ewh7JCO8eZaTQw4JWrPa4hExqAwU+bgaLWRvS/M2WMMk87ksta/RCW3Ox
bl2xxsXc/b2syt/ei0pPL1pkeGwTc/Coid3eWJIT+OlwpvSPsTLNKbGgl0K7mUZQ
7es+XO1De/sDAlz+RIiQHqqDOviKtOo8v8LrhWAMnaH4HC3qepotESNHTMuWCCTI
/GyeIzUAQz7OYYbDZszxS5KqcVvFUj+Xp+izT366HXSpubuuw5CSyOH3PcO9EQzE
1geCb6UL9S7CVBDNRn7Fc+3ui13AecaQtGIMECzFejok1W8VhBWBhx8hEELllGkS
rExPr27Uyfd7k4FJT/U/lnsH+cdXHW6HNqBKAH6MDlUBJB37MNiCt5ulBgy9XDpe
ntOG/0gU5uq8ltzz0RwP+cjpuUJVj6SgSNMvyQZrYcnm3cfCnBQVuyT6mh9AOA88
bNcBR/M7M9xAKKFNuy3zRFsgTAXvREfAFcto70HGLKZayICW4e63nFTX5635NPFq
+o49pCE+85AZ4BkxsjN3K6wlrf7vpMcx51HtHvM39cD7Rkz4blr81OA39eN+Wps1
6QCOGziNtxSF7qHhnubqxEysMjMFYN2zk1VjlOaRXDKQquwh7qVGaiTGE+v5u2m4
m8BmTWFskwDkAXaOHv+dGVLGGe1pRuYbFoIX7mM9TyGBAwBbVLvQkxj7cQPqP9xK
API4wVKxOdf8L7FmzY0fxkBkawvpjI7efJk5mYI7438/y9lvotCJFoJRjrQnmkuN
dGpn4VHbIsdPnVKAVcAjysjC5XrxTFjCBGlHNUkVT11obCGVBBGylILHaYXKeG2B
rfPTJ0rCn1TP2CDqow4EG7XJI2YdtM9LgIe8OS2PDR7lusXPb2ZKXx/Y+FCZ+xQL
F68+Sdxu+Hg7e6fd26nBkLy0g2Wp8OvBVL91q8LWPtqIGlxJPxg1Vnjk7Fm/Lom7
my+hyasZXAVPlP9SiRMgIhdrTev544PIOlAnk6mnXUTtSVXqwzi/LiwKCZRjKDoi
qcrhvZJ+w3YCY1PV1i33YUbIh8j7gg6gJW5MHsaF5q1IdMVO/nUvqxoKPGcS4f6r
MqFkCpQb8NYzV+jjRHdmjYycVDlHQR33016wwrbAcM7UZbEnwZzniD/TICw1ZPeZ
DyZH0+oiWlLGYho80NeTdCbSLdiFoRmm85ZmRo4jVFruqmYfjzSCcba1el3BFEeB
jKHgETyQ+8UMX/vlOkL4foW8RlLthS+lAe6exRQVtY0QiAjEOviR+2cVGh7gvX6E
A3v/3xfv7BNQ4NKAK1sG2jIhkwsRYh+lgO3aMhZjCalVx2fs32Z6HcBV6rS6w+ku
Z762VHPGI5H6S9s2ovjI2QN730E2fQCKi7NE2rbWnOR4Ru3x1QSDVgy4EqjoiOR1
xZQiYc5AXN6bbpRalqU20VhaFoqRnSQta7RGTLMglRqa8Ren1CAlun5TZzQG6Pcn
/W8CKcEQCxGlUwmgukN6T2R91CNwytH/bvBqiivr2sZjWUfFx2COVtC/EUIdmpio
jFTc7SvtJU/RoLZBSEuE3C2WWNiZyT8Bz/t0BaK2W48TqnRpkaK6hgqujqzkqEuB
KiDJyJLU+jFvHZUqHQAqlrPxgjyF6Ehvo7k18ivSvuoyUjERttmh8BZnGOgCvqD2
migfa06MVAux5/TGFCkgt/hA5/TMqapRiiljCxccia//HcDfR1cBgbVQaDrXb3Jn
OmcbOSxAGD8+VQccX00NAq1IoMifdUA1g64Gd2QmFMIgU+VlhrzLzujWmu1/KOxG
cMUi8gbRBmwKuWiViSqrwJ8JAo+dqN4nW0z/rHxPdKm3lffF2vitQLA+trOqbUEm
S34xslNoWdlyujbFP4mbzdkFBRND60KbAg7jcGRLbndrAHegY3YUD8YPAsKmxlg9
62tNYBPtl2ayWTY7lC3m2xal5U6hJ6ryu4OnUPS8iDcL8Lkf2jqqIQCp9XrMj2Ct
Rnd/cOOH673f0+g5Wmo5338Vpy5P4vgi7ex06jOeCa4ZoMfPGvO3hBFxx5iAnoDB
qBGHTjdAVMyBQe2lIET+WHzc2P6qGIFNVjo1WIr90xDO9ETpU1aLe+PlU6m037lP
I1u1lQnz6kVnU4qiVQWL9D0FrmRbxllMkni6REysDW8MYvKOGk/AL5NhtLMZsjoI
TnPPnqp7pxovHTrvGUZFRDdvBiRh+Milz/xYZQOSxiOFK7BAut42EzReIwgxWzFf
9TutQewZJezMcYOPemD+J3f1nEyOwWmILNBJjlH5kJavxClZpI6CRVE8AJFMUyJN
6ZwS7bamg+0AYUUNWGDcxWkNztvpz6aabKrfMWgaFf2vxt76M3hwN2hxQhrzJsRR
H/GePpo1xSyg4327xRpCuCaJQbKSB9SLG50kIDdxOrP1/7UQBh8acRJOByXRGDHl
a68oHGw98DoRYt0IsxfYbRog9ReOUcAkjXtgbHnNV2NUZU/VnCHJ00cDQMi8BpkH
jxUxvi4vhGn3mPqwAaN1RFwTJ5w0XB9dI6APhRLnwyYr1X9GYboEOvZWWj/zEmV5
ik6s6E2WZCry+UQNtmGflRBQ8zsNBkA1FjCeUSG/hBIRYgxudWofZq1F6I3OZ/qq
lkI4sPklv45w1J4vwZikC7uZOnWpscAfV2t4mbQz9TC8VsNHdzaCjVq/pEzz3KtI
RIBG+QBWUxblznC8Xc5eaxZdDewJIfgvDBhFlC+XitSuI8Pg8ZCtccdqX5lc56Ad
78MFDENWN3skErNMjkyKZQ05muyKuC9WoA0PDuaRC1X0EaBW2zxH0Uo0FC7WHKiB
a/1k2BXClqgUEX6xJBfhMgazxE1tSE91kv3QnEFTWlZaz0VgVzLlo9Zv05YY1Y/y
P+ix6GzmTjTaKneewvzVDhmM1sNtvpTRCHqtDd9ero+7nkWOmpcCYjtevQXwnij6
rew1MFGcaWuB2GOIZayb3EZZSPbCdXs5g9EIR1vvH4nM+t8ywv3M7UjeiBDcbNcx
ni2B4flB/u4YRDan8bMWYrzewQ2+wi6dcZa+JstpDxdFTbu9pwZdRU5c9P+Ot9TF
QvL0tuJ4PH7QeYVmSlGS+gIrKasLgB/XkthhXwMF7O2pdJVgXg+VqgTiaGoMO5wO
rRxIZ07cm7ALPQ4MBoJ5ZMkwJ/4dy85eLETRIX5Vh6xoawNJiVAApVrWHhbUebB8
ZhlCH/dga/G0hq6XOzWXbTkUdxryzmOqPKcq/FMc+OPDqZS+psi8pLyZF97Mocdc
3FrzEKGuwFDotys72aF3+2PpTqdR5/4jY2Ijaj80shuQxCIpgp8tsr42fOUDGJ3k
x7OvkRDPXALpj9fXgPylcbgt9op1T7naKh16NMEVxB+nZmwawGI4DjOCbBVO49sv
VGe7EcfSimWMsr/7phDRpEskExEAjsAFCvpK6huZpV29Eq7ATvGjl/A+owVdV+iJ
DbMttb68gRBPLRyk0IJX6u5yHkz0upAlL8nhhwDDQk6gT0qRGhDclgd9y3iHk+PL
9JHh3FLButRXMGpAm1BwG3qVjvFBf4rZP2UYF/B3mniGYEPy4ksuGpkcPCFogg4m
NCouUNu623vooBZbHlu0NDL1e859+RH23ts2MQu8BGnhY6fNXqz0zVpjDwDA9ax3
zcKZ+FhQLwO1v6WB4XLWeRTS4ZqEciZ0FkjNvR6elam1zszB69c0/8NEf+ZYCcL7
XL4brv8FFIycDyaife6kNzWzXzkxJzWXzItTlq+Jlcdfqt9SmNTMhjwXAvpwX0At
kwhTXumGrx5xFMaYixztDVHjHq+CXQeyYNpubd08RQqNVTMdLJbbp4coZ2RkwtQW
ThVZC1op84HGaP2qNAuy4rNVyb0DH9TO7FznXQuwOCWtAHONCNJtewj+hks9PT0P
NAIbkx2gjaOviIAkFWrlyL58luKCkHFgM+yZ4X4bx/4Xnl02m6x7qmmJlna4Y4dw
C+HVgb2SdXHumHOnPVtDqdwPcbPrjupViE6e66LNujP4KpmvdbZrpzD/Q4FLLp7B
b46TJS7fJgcRh4H7PcuRUtKmj8wi86I+9iEQrPVpWaeNQRiDe/98DXNgOL2AVmUb
ZPcnaUTMGEW14xON9+gTmoehMH5m10USpLL+MPl7ssnb3v9qxvTxDT5grOWRxQJu
2Cpnr/NGqKEd8PL8xwtqDC/AknwYknV3ue+WRusApkjGZW/t63QgeoKnN4Kqf+0m
CHm06OR23JmwFU1eI7DaxqYEOq8gjPx9G7HLB8MC5tEmDE6XwSh35QquU50skkAG
4MCtQq8Jse8/bZfK6YKwNwbnmYLBHxDAKvLBNTupAmwhC/xnaxDtQlETfJUvXGTh
uPTdllpT9vaTZ5sUdocIQg5Mbp5P8tyC6isKlKT9oLo39HY1+uR07msAfUWHVE1F
ObwIvsm1pCVtyK2nKaqVfGyMtbKK5qbrD5EpPQpLOgVxYMuiOOyUz5zlikjpA32r
UDVsLMisXAN16M8BDvUw3F+bjI58lgkzS1YptXEBWekHk4qUZx83RvEGWh+mV21n
iYNVbiDa7mhGRJNW6LssiCe4FZifzp9G28A9nWCfYYts5k7GnyddvSjJpB2Skobk
8YqRFSYMpHYI1h+LFYo1BitSpSWz3dsfREA0SA7oUSHqeoM6dMpKN5x/ukA5Xzvh
YOedX8tSpoxSLHxzEZo3oJSJx+z3BrLsjnBQIY1XqCpaZ/TED4f5u9WN6qHRjnOg
Yqj8OjBPZa7HvRwrraM0SI49EM5mWq8/qP227xwc7hnqTm7aEPu09r2BXhqLjRlL
GZXBenh2XlSPw7SpndRJtlvkWeMYTtFW90fldEiyXq7S9gAWno6LUzCpeqndKIbM
AFRpMzx76z5s4e7hwldqBpilS5CvTUCLCKVdNcuRFgBqH27wn9BDq8TiPNrcbfld
O6WmiFFjH7bFiE4bNwK5KGJwJVldDNWk7QEoc3+RKfvgBp0yNJaahjKky3KLtqPA
/inD/TwqpSOeD2dHLFhD9JUKhBRftp5S+53ohYDbh7g60nhOpFrQuzucUxNvD24p
vJuSUQFGLusIKKJt17l5/qeZXRJuj0xgcHovXdkm9zKQADvvqgrVrRLyEakUmFXw
p2z88QvwTKK3xk4dSLGUU+i1vCUOljUiNdC0cHVCMhbR9khyTegGGaNdokT8REWm
gVK83am1d85SbNEwbbcF1Foohj1SmKwpXEE4o+8MCGDkb8YJ0K1P33H7eFqb+BVP
bjt2lcyiro82HQyKRLpU4JlBPXZMFjFqLnVv/dZ3TWMwvXha1LgJaLIuy1wRu76M
cI2pViMcNBEMYsJWdoEscxlZqpHJchgfUxxyd3+dN/20kDhslq48lwY5/pDJs+3g
+3+EpekcYQzrJH8MJZ2TKt1mYS22Q5f7gRDSU1PIkYce1OfH0TCDrtoZCId1kIWC
0ozqpZ5pLeIISRKGdyczEwWQhgZ30ubds0jEze1INADe800pG0yCzhG084adcY9u
t/mEYs+XvlxoGMwaR9hUVdDCSvptNsT4a3o8ktdfx9vxIt4uni76pbrcCrwO6RNA
8HJwp2F7pBHVFYyu5Zrc6zMfiz8cz2Qxybud3Ubg0EOwXhfF8ewrVoZdTyaUXpOX
01622y6whveu0g2nt1N2wu+rCqWXLBASRIzRp4UNF/qJJmrnKn0/0grlq7NgncV7
P2qzo1Kqwn+wR+gIJG+4piuBrv1UkztzMXdPgiz8Xq9vi7pxaODlkIqJbZMM61Qw
CIWpPGWKvwxWrvDuRZ78nM855ljL3HqD7aN/1jPa2k0sjd/PFpx0cfudwwwneAnG
ycpKCmHfqE9o7abmtVHYDXaEpGQv7RzL1iPgpvZ6ajmlXKsDSF5Zn/IEFr+iSb9r
8VH+loODlby6nLDGQbezfwAmf8eQ5saJYJEYve1/WFxx7buRSECFOsQGM0OXpmrf
yueiqyNFAcxAA8lz4mvVq2HnxEPpKWroW0ZFZTz1DcW+5+DB4Ga3HbxCGGFGw+2g
N/SIjWl8Em8wEwRGLI0Qr/OVm/vWRdK0qpKCVXvkIJWsG5U7hN4G901MG+A3hsOj
5W1z9wqDaCA2LHk7Mi0aV9lHj/tymhR2S6sq8evo3+7dnuYe+8kaEoGNxha62rWg
PFh9zUX4rB3YI06duaDr2UikNVnsMuoA/jkynblfoDR9ohrVXcCNqocp/pmJTTIg
d0pkHRXtX43f1VUKKKWqQICD/JYSGuRHAjyWpm1fFetizjZ80377rNi0YbBZ/aHr
V7T8tiHWW5vtTQI1gjN16Uxvc3hUvrsab/sZ2wrJIr2wN4DNz5H4/cblEEGgWM/L
lx7A8hCji9JCc6VThE3v9aUFyUlXWu4Nk0pSwAzdlr+fWcxreucZCcHA85Ok/Jgg
rZvkj5xCsUoABPYTbxNXtEGayM/Q1TndK/34lg7YOYpdFzY9DT5nprMoowIWLvLG
2UKLSjPO3sU2PdRoMDTNaRxyJMJtvwRiVnC6RrY1ZhUIDz4Ipy7aLVV27gWfj5ut
a3M95XdS/CqZqy8UuLcOopq7OTURfbOqwLNENknLuZ2+SlCjAvpVFDYGaS/5TvcM
WK1mKBRqKR6FLvILomtdBnPNAqCU8QQrveDjWQJ9qHWzigYR5GG+a+BpAlPYJG88
1FX6s52UMGP2D3wrqAbVh8T+7GPMGfXVpz/T3jYCMYR5cMb586z1dKpwVGfBdv1q
8VoJSKvDTc+F0CD8YI/zaqZYfmBJxEdBpspSogwyS11oEWLfy255/YKs7g8zRJue
PTKLaTsfqcMUGPQQ1GjUmQpXwQAZPswB0bDktNRcgdPfoy/V+8k5hWRJ5J+1JB/7
9q1jRuiqNxBZZwyAfA877U/FDJptQ+5FX+X5q6/ENPgYN6TLI2MbhrXgRG+X/8pb
85KaCTcM5JbFJz/iVHEAEqOv5lSexerri7UnE96osZxQf6UNFC8klMuctUgFy73/
CiG3D5XoIxAa6qwrccefq8w494uJsThOgZsjwCzPHBqywuzjEyvd3oNH+ebVeqaD
uoDlaLBWNVUoTTMBOaNNi6npzbbtpvvxEwrNHrd/A3UgR9eUKXcnaPNvMdj24HLn
krZsXLG9TcyfcVmW+z2VnhWBb7cuTowQEbsGIocz3TBz8URIpZySzO08ZM518/Kz
j2xQYf32snAJJLmFa7L6DXqkceQfPm3ET0HO1wA1b+JpV6nbPNd0wzdls+xzwvqn
rf2DNt6vGWlJ8Z8M9khnVjIYBf6gY5Mnt/D1sNe+b2zsb+o4qj3JxB0hYN8+LSkt
D9abMv4kwvSdDDs4pENHn0PUFj5Ja0a2jTFqkhc1iIX3Jxrbab6iuUiTNaLx9j1o
hLMP3+Hg3cfQacCL9CPedpNpJOXzax/Ds7FB6bz9fdk0CQKPi4uw7tg4S7PICwLC
knfWhCec+g4K7kuFFHHV/5RsJJLmeBezJaeykPTgCCBZJkY+rlWNxBybz7aXrBB7
9uf3mWL9nBG7PVIyXSmcVgyaeMqV/uO1G/Xbim9ezajCOdZ/QLP94xDbboU9681u
1cpJyH5qrTvM7hlFYX7gSHZkxOWOzsabSa1Ak7uNAezxUfl8etCXRaSCOOnGDdYp
Ld7qMRixT7huewyNF8Z43zCxM7QZ2HUXc+xofAOfV4TQUUHH3YyAPOajB3F9xT7H
jUQVFkj8CspeAMlqjhF5AQHRKMwmJ6lZ4v660yz/IXCjNxlHJUiwGogiKFLX0xCI
dVPTEzm8kHwRwIH2jiBJmjRwuDaV29fj+nRSU4BPtVi7SAKeGS13ZQbYKVINYk+o
J9MDNYwL4cA/i7b3R46y0N/ga88Ntw+bRnq75GPO0RiNHFMjsQJRPls6wUWM8gVY
x5ge3hWqS6Kcx0TgC9HWF32pxPwtKKu3BXeBCLD/ZlovXPA+dBLE2sU4gkDYfDhl
X6GcURzuSO6d2Zvx2m1jVGYQ3GkWvLNCpckAqDtS7h0ylZ1eWbmHSGS1uFAnF5nR
WoS3dSJwvU0TkbgePAKCZVvjrRL5eekaihZ/D4Hp7Pe+Ld0HCP1XZ6WXfzQ1TzA0
rgdOd/lblgIWb4xwTb8pV7edZd9obdCLDvqUTo3CXIkcd6YfAigckajGfZ5P38gO
HE4a9bkMiz2tKPHoFnsBnc9G7SxKkIgAuXpgZOkceAPhMKKj6cdgBbkruo6C0NMw
M5bjUmIUjt7hX/fZUEc4kflREN4hPmSl497X3LBh+ytKHjty2Y9pAH9EXU1lvCF8
X5XdfTuHpohoDPzHiXx4bqbg0kck8gnCDSJ8A/PMuC/0H8T1F6W2zp+iCIzLIPR9
YxRIHh65U8EyYGcG7YVP6q93wCGAcwcsRX2nm6molis68wtnJamSqDBJym0mWCeh
gn3W/y9+2Wi5/ZR0U9nf31jD1ZnOSUXusAKQrwAris1OXGxDvdRbEe4+1rLXaRPD
SRNuWm15bSrvGw4QQp1NmvwjIDRIEJFMYTrfvElfc7aqqH02oMgv2s6q95htXIKp
RFADzJqray0Bjlwdya6g/EAuh3rhIiwkEAZl4rfSofq3XyDaKYxriuGI0KFkioZL
0mrGxCX0nJDDzUH7KFrxgrCiJuptKL4hvF917esrsD23z5pzTyhi6/oIne0V3Vec
uubHNSDaD78ana6zZ+h86ihyFVx2IgaCM/NI3eaY2D/2+V3qShcpNCUfRErkWgfj
7UtdIB9oK4jtIE2wAh5uYNw6MiKG7RDSNY8OCB+LVY8lg1ZmCnM5j/i32eC4Q/ke
QSIU5WyNI7X8f3TH2a7boaCB0IL/SQfHzcFPhl8gUZDjXOTCZbbm+UQYN+Ou2Mtc
oYhCVSYuYXsmBKSroNKvQ27UoFkERVDKUTHqKUlyN2fLJyigYTbTRwsZYj+UxAQL
4M13i75/l+7MzoyCV728u6s6D7kqHF9EE+2Abc3oAIULLJ9htbS+jam+b9fo5mgr
iAukkp5QtO8BipmZ5H87HA0A0xB7NgUvGJ8C7PiN6869Wt1cWHsoN22keKUjdSZG
UpUIDp6+CIEx/3/NbwCyk7yHpyLDD4UO0De9GXTl4xu59jZxZuZqRRBLdhFDX+lf
iCt2WFpcomC3bNfsAuN2voO4QAB18z6Woz1RDN6NilsGPcT+jhtNKGFAFUQyJmZl
vaZkP0b0ldgysS3uPPYveFl1Ud9UbtSSsV0tIaGsGZmD7DL4+2W9ZCXK+1R2gFqt
7ugNDXHOEC51JN9KNcXQNLQ8K8XqXhCc2FybKzITc/OVx63cHc1tdJVWQgYRjo0R
rQon4rlsRdFI9XLg+Ylu3kkMR7ZQYtXmfEocneaYhW7MvXhNbGb1ZKPttmfJtVng
AzmJ5z+SJvJAcmM8ew5HukiRD2yTp7eICbhBdysFr3CJqClur3dK13I1EDSl5R6i
LgpSQ5ZDSdfwYfde/IlsvjBXQOZ5ZIZ8xJN3AW8Lkm7PksLvsbEBfm41V4bwPmCm
XsNu6fqL9MzHD6eIgqpEo91gyZnu7kx1AtrH2rEux6iwiGK1DX/P9jQfGeQi+h75
4agNn4Rf9GPJz9Bm9fCHF84JreL2KxeEGIF8XhfAKCynTeQzmFlNeS0Hs3yvhrTb
eJGrLS7iDh4NSSZ/MvWUzAq3wPC7IBeobBfB1jPBMSbZRZzMVFr7uEVb2LYgkC71
oOIMFHCg9QeAVQiWkm/Ljl8cTVDXYpm2DYxyhN7vHgq9MqEHtaZpQb7u9KmBURG0
8S795OmmxpcKmVkCWJ/KeMmO83MOR1BhAz+9iJPoYVJ3UzQgILzQB9wOL2/Nqv6+
tr7dO4WmlqjROv5Ki4LGIR7se121pSyBNKL17IozhJE8yebup7F9NzrRMZMoyv++
aqDEiMi9RC4sh84PeMyf211kmZgHSRievbeJ736ExwjPEi+v7/YuAVL/AQ7DkrTY
4TRqGEDe/PDeJ3gtvzVBE1nKqb1DPRKPDq+hn+oYf5Xy2UAkhODIItu4VQ2zRxw4
Pg9H+SkuWJ8CktsjKaXyf/nN6ns4W9oQeNqQhlx4dfdV4l09gZe3IKpgFfEy4RbY
1g37nK/avy1zoDcppjWZ7kI6C4NauKBXRkQGxs5Q+ncCFwyIOF9AZsWHRqF3/l1c
smRv1wYNqGXmne1Yb8E3dpX0FV0wchLe8TS37NVkTojsoSe16h7GwI0DjHmvETj0
w0XeB3RWOkTzlQsKcFfHL3XKLQ6EZ37uw+3puABbedjr9Co1uKlitUZphUXh4mWc
z5XGBKd3lxvIW9I1uPl6iCAHWVftrEYSv4N6Td8gFeBBTD6fxJkf9PmnlwkP5mzE
R+hIPYqwRvOEmk1J4apV3+nOv9uKmwrwJyEQebtlHshuDSjRaOY4yQ6vPXlnS1et
TrrEYj6XCbHwMxKDR/04hbmu6IGpCWD8A2r9hMflDutsSkCzk4aTX5Vk3BUO+KJt
XvMEoPNp3D47gvi3ysx1jyMWQupI996fT0THV/Bv3uxds1OdQefTGDvvtDCDPnHa
xgD8mDg7ZRHiqE0tOtnVuPvlRQL8NZ3QuZatRgCaGK0I4K6aVYk3KOqxoaRY6iXA
dV/iN3NMoFAUEM4yLJmp72rj50mXubYLxZBnuN85DE0vXVqgyCJty+VgTnJtommg
w8dISf4l+qXpoyYp+++5pEqpe6sV2D1pHIWUGkhV0j95qDhIX7Td4PjDdUlQadTg
inXjY+l5zi2TGrX7kUg547P3sbkjAyQU+uj3aVxU6jKuemB2lCdJR4WvFiYVc9tG
lVTCTjTb5E4sm50oUsccwb83YGy11E2rLIyP5AuS3C3rWSszdjPdQ9PNDVzMpnlx
HRaaiD3In1NDbh31ffWe4AS65dUhzC8DQBjtYJawaVURV0M5MGdXvEGxYhKKXFxp
6xsAuc9ALOjLa9E64gSy1JZVw4JXqa2AURrH0D7E5WiJxJXR/2wLkV1Uj645KpmT
akYtF29l3w144fp8fAdvb6xyqGlgILkwZUS/ZEeailF5/KK9FJ4oInn3gCOMMGDA
vefPheQ+XxBYgv9EXppuvojTH2vFppaUqYTOSBJgb5YL112uBsqjzt840ejTr3cy
Kyqjva/cTbZSZrvtJ9S0MHhJubIJH/+60bP0ldQaC2Qmd/PQTCh8Gv/ezU/FBg1h
B8tdxeZOox8kG7PLUy7zA61EhswEsVr76XNDx38bBxD3S/6ctZ/3cciz/rmjm4rb
SYCinsyj8ZqkFVcycKcy84k0gwf3okQRhk9XJAiYgmyfYZ3FRsc3xgD5SOG2ntIY
nQJO/ygc0Vq6ywWdO+nFTtWXh+r5Kqn2yXh5NFicXlgjV/u766CHFyvt0oKYjZyP
1Wbw6sF/EkEU4mAvDfyx1Kd8jyopUPy9vsx0V4/DBIN83VfghdPDgN0rmVb6g6/S
3+iqSMci9ay5cBvGwvKPmi//4xfMkjprp+rLS46lbD/eguqiZF4zQHOkGZdU5faO
DajjGFsoQMD7Lbvpnv7OCO1Dpw3XtnNA8DYNwblWDxC8XBvyV+8BmN5AOQMvDgwu
30BAOUIS0ma/5DL4iroE49wiNrguq+DF9MVvw469KUQCfqJlI2N/nrm1VKSMMJeP
0/bIXqhU+KVpKs5Kn7onJdtUnlkkIAMvSHl7TTFzncI7RNb33bw6FjYiceYj3RTV
gTW1ns6S++el2UllwKbKi9OjBNgdYb7rorNo78e1WcGP8MjiGEGuhIo6d+N2pg3M
BauVvhrGAtcx8DzKxIuHjzfFKvfq6TY2d7kP99+43Lr9W30idplLyhTOGFlISrv1
u+PK0qP4MvW9sY7Q+3TxDbVzCCEdC9wW76dVdJdxrUqhkCIj4P6Z94P7Fo21ozun
BDuR0ZRUtyzMU6Kwk2onRke1pm5qMCCI2fbeiXrckStvn2T2qy4TindiXp6cuEPO
WNoMCdlTA3PiMmJTxdNZZpDtPZST1Qk/TdpNWIiGfNFIJCXHi7ZB1H9UKuWwcLOT
CYtJeGvmBAWQ5zkZJRMyRrRFT3JyzNTYesnnMDd16TeXNh4IiiT72F+8o6L38gdv
jcmW5mvLkvjFlXRdYQB/CFtq5mmTCdYTOCjPScahjh6Ynf6tCLiJd0DQyqyUyRom
5wQWxdye+0F3AyeSvAdUuzmQ0U/IGHqvhEPIw1fmZfP/cEcay+pYCznMAs0wLW3O
ymr+OiKwo2txTa63l+Dn5J/BXTr0yRPQfAz6FUcfvefVElalZBNjcCSmzIcRrIxT
FZuE7WRK1vxh2LCH4GQlo9BoV2c8R9ajNTulFG1Y3fWhS8Ta6eBOotWsVHzKSaKj
xS1loy9PEoZ0Q79EX5g0fI1BldivmSp8SlDuh2ZeE6SzZdyeZTzKBOiJLvtZyeRF
heER8zf2pzu6PKfjvJseHu7vXdz+Uc8DTGymcslpRzdCoIW+5GbkrQdQFqkABY7S
J1xLRBdpaZBEMo58+KG3IAkkh1FTOEXYl1LEsOXplDiPqImpF3qdvt5zceJpu2sZ
AlfxnjGIC5gvFyZvpTRB/5XXIFpQcKVqEKWGG1EDxZT0RlC8oDfR0sK94HDofPD8
318kpkVhbZHR3SfAh4AlIiAioCEfsHPJrymh43zRcbQZGGgDf+95Jzghj6jx4ibK
VVroQeDts7ciTrTmOW7CTOyM1jew0vM08T4+H0UeibbuewtHpg4PI3VdClrBcOzG
VzB6xVxIC9Uv4RmR1VvarIKGYsFx8xtWmM5ssywxXASE9PQGXAY6Pe0G0Ig5nAVM
JKVaQhctkJX7NNmk/WFXVy+wJnIqfR2fcu9PGzLoTXPPfRhjS3EIZ6MRht8Wzy7s
+Q0/M+fheri2+bw0CAcj+dclNhgYdNr5YwdLsSvv0UARTnQ6iuEYJUbhvn/2VRhy
H6GaaF+j/EWrzDrv6amxxFed+gZxnBAAcLG8V6TXDEWIbTVQqx+TIw5+LtQT9Rnr
whVAzInTsQiN/MlhnHyM1JWVAuZqLE2NcaKgHdOQx9RaE08LX9lznMOaFvqd7yjN
samYOZflD5PK9G58fs+BPUJSTW8sGzgt/bgQDNMGLUYXiGH8dPNoUstF6lcjmdmJ
Jb9O06Dg1AqvxGeqaIGE0dvXTEibgn+4rHXrtIEPThE2yLsFWGc8m6FAGI8YUDPy
jhJTrqqrP74zZkZ8iDC8dyAAFM/S2bt2dB/y10RrmNUZVW/tZep1Sd86maojnY63
oCxmzC6BEyxGqi2UC9FHnoZ/bsWRu5ZjCd4SoMWLL//GfGomRUaXkczz82upfVWb
NlS7JGRaKLoAj/tFIK/hRncA4MDCKan0HjZKJ8JvzPPrfwWsmE6LfTF9r0TlgcB/
XK4UTLifiiPJ9gGIPcfJou8RMpurYygVV3c1gqLhFZH9AiycQC98wxMoCpaXuRAh
3V16hiFkJiPmA88rgRfVwr8igwgBIx5YkqK0byUi4PFX0wHz+trZuEwIyjh69rwO
XMwRlLnoFfN7uUIIfntq2MzsQHzD6tZLKH1IGoKBMObSau2ZVktnHdSfZ0dwU/LG
bsevOmH7E2u/Z+F/dTDHeDixQrfCc82tePbYaIsknb59DoYqW/upaulC/0cwruqo
9LRlsHhu7VmkvenZJdmUnEka/CEsULZuoaI/vOfOElT9TfH5L8BBJKAoWdNZOWf7
Kgt5smmNwsZbFIYiuE8G5SmdxOaxFoiYEKC1+iX9lryUyvjNGNEzKlnYdc7QMcmY
v6f1JIuppBU3xioT2xXttg3B2Eb6cv78gjPGYhRqFG7q9IiWcmrjdSXBjL233xIb
boPv4cBfchVFjZlNbkEANnurQ+3B9WpUpPs8NQHPfku/HGY87pRGB5Vp+hLf5Ly2
rIddjQyzJiek7YGa4Bx5HD2DuUrzPG4uzBhjZ/GsHTooHHb0ADuOIy1WXgv0FBah
BbcT4oiSaeqxA9Ka+G3xzah+zHFFKviFBALaNoVPJzANel9hNqP5oJ2RBiQuo7MM
UNvXQZvVP6KDeR5yM/P9WOTt6fGqz6XFqXLUTmMScuBhal07g1UgB/KSGjItfTFB
RlfNu8ZWO/+gBMM55tkYWB0O9+GHjJOK42qUl2czNWh1XUZQvWfrRSa8D3M0qW8I
S7l9zvsZwCwIDY2OEM3Pgy8kIR3SL+rKHZ67mdElhtBHeUBhKtQKwnpdtB2FtuWk
jUCdVtEoHu6nkVExjfLw5S+L0Ecv4lkROsy6JHFKzZ3dkvbabTcSLFBoqsaxcl0t
m/8VWp2pwvYPJ0CtqOKo0+/QOdvjY3lSkW2lgqB1LxBYyBlWKfRNc3q8y+ICdYbL
hFRY3c9/L2bUVUHOiKZ2opnCFG0cJU1ARhVMpTRrY5iqAAiT5/Pxpma1kEBiYRAR
ZT7wT1Wlkf1Xd/FQbE7bJ9PdPCMJZopky7mFMj0w2RnaVaGST/FuD079xeCukVZ/
4KTjqieVOfTMq3smwSq2VEJECPV5GuWyw5PcT4DdpaLXeovEhgFhA59A71wLqWPg
ntprfzOTGaTfJs9Mgy5MrSjAL2jWszgnvvjtFT6RjSPptZnyheqCwfHgWsEXpuVT
sQvZddIfDU1+7IR6x03yee4FRPN1zKV5ZcsL4K2eDI6xZk/HX+YTS5dUL3HZkFzp
34ZtPZf3yLuR1wEVZPizOVHOiJZSOfra0lBvVkx2t4bxObKbrvhlUfpNmF5er/GB
k4Ml6HlIY+LlTIGfo4tkbFW59w2KlwneRk1uw/SUWEEydttsQ0nM/I0z06gLAa/n
GPiP1614gF37Oarl5MrqHsbQIN3I62FGioySt09sdsZQaDqvkEG2Dm36Xq03Vm8W
Vl2dN7GfrLkTf31G08bJ/AKd3whegSjFvbBpzJYmN/Xn2dRav0gSKb17WlsfFNLA
zL1o3lXg6fcTSGGKRjH2rlYWYEAuprz7CDKF7O6x3MEdWywBPph2WPfqYz+Oapci
sv9x4p7/ifQIPjkI3f+ycMOc9xiBeaYqEX2YW43REJ7nNTAx8+ySQWx1yoc7v9Hv
YTXA7ZKghoWxqJ1+sp8AR0nauBymaHRJ4dlND5MyqlNoX+cLrYLX2BubJMYTohHp
zRcUdBDShCWV44YJZ/jobmXeQvvz0s2QBs+wz/gA6X8oqYM+FX1OTuH/elcZCe0b
KpZIIGfSdRdJfTUyWPi/fDQ4r+hBgp6PG/FGeMYSTAlcjp6sPpcRmtWbqgE3NI9J
C2Jq3mbmvWFxO3g2RA5jBqvXmXSF64fTvHlbsCxqgwJ97xVQMYJAhdta2E5303Cr
VfsmMZ6iT8eic2QM4c1hDpG5tkBVel5mP+j3F4jDwnvT36u+KfeSsOlL4HHV/wjg
p+TJul6f+C5PAkvsIeOhO3RbqJbij+6WMtITUdsghbfmWLCzE+lfq/SCL8XQ0+TE
JH9/gkhFLYqFzDgAGR1sYbbHH70tmPlbPrxjx6B+x0PJKneceNabhDf6RKVGm5AP
AuYE11qbXpYwYzmXv0LEaLjbWynBiYGdM1D7eanpVKkGGFjGPEpSkiUgnATizU+J
02h2/CruTXMsbVv/N6kykpuR0MEuKwYieXE2Nf9NGno7J/N95jL9wqGc8oM4T+rO
grbNcnQ6w5ppk8lfo1EyYSfOiuna+KFVq/ChlacJ48KdmaYnj6WPq2KcwdY75xX1
okdkziVMbnVRBRH3EsgaRUtwM/TyNB3jbVF3lwkRIDJuzJL55A87zdU74WYvA4hw
GnhCr0WZfdMk0pMpXGjGAy51fzdaPEXkqjQAG92PBRu5r2JOkdzZvwilmFle+BZx
25CTY0ujcCQAm7Fc5mFh9ITvlX8h6CSnHTKFpb2PUbAiGtImBu+Q8W60A42h7D7P
+QN3wPqcI3yQlcWEJBnt0ZsUjTgP4hLcIWHGvD/5Rm+TrcTJkHmyXipKkGN0Wtet
o4Lzb8yjjNG2vYD6GxovxEFWgQ/fRYXby61YcYFBaNlZpEtyostnJHO8GqhgvfQM
zEz4KIvApVr8Z1N/KuoQ77P7LP0So2cKboA1Qag2wc/vJ9ZM+9YcO0aq/roEs10T
2yKbqrnOwCtQBh+YNqAVQzVhceqNYiorRHyydpjfW629+K/O5reRwpnEfbgrg7Ri
23KG4vwSKU9RldwsdX2S6Zvg8yWYF0WuOlrhwFYYYhMxK59J9C2wkAz5QJijrm+w
8egaG+y+yAgxIvY45+6uLylScaabCGQmbrbFDyedQpyEwkA4ioplDii8UKVL/fBQ
IbfIR74EJDVb8glBxVMK3TpGXzsW9/jbGdItLAJTj2hu+5QKvAWN7I2OnS9HnztI
eRahs8/Zn5aQXoXddP35tqRArEjBvwaJWioLf+RsV+GyrrYqsbtaXT1WboCCMSvd
2je7zWR0v7BnZYDN0ySEbaux6nplsWVOksDRjbo4KAbnI/vCdxf8lTU3QYEGAHkS
m5ulOIl3D0LG7qJgWvtWw90iW7tCtQvmp/V49JQwnsvPbVDOLr2PtEKFUaZPBCq3
LzgL3Fct8Zqxc9HOrGxY3Nnqtpj9Xjbw3H3CgB3sczZal7LtWI5IgGqacYjDlcLt
nikPeV1jO0ochtN9D852vpC/iC/d0DbPTaembm+dfcjyKbG7awY7DwoiOtseT1SD
IxcPULoFh2g7YYKk3C9VkfZuVUra5G8iGKqByFan4/XzLz/KHdhED1OU8rRcDjkb
tOfuj5KsmKJWmF8VY368gFDKEIh5EIOBQBBkdmdrP1bKPc000eXrA+HEoE2Tl0qr
WLfSe+gwblNslCwZ4nW71g7TgVMoDQWtJNAXsPtRRKdrrjUqx0ynETsS2OXeBPki
ApwGgscfPzSM2Vh/iqVg0GZjW3wHrXNCPu7ymi45h0DXDe3IcQXIwj9wmF17CxY0
PPYqZSncThQ2Hrzeu0pT0vlRc995zJFphEYNU5lhtdVde1J5jX+GcO7snlqbHlSS
p5+hsB/nXkW6Hmd+5ugORn138PlWRF/TOmJbEOGjyJOHMGLSVBrcYrANXdDZDk5r
d59EIJ+2GZ/GmbgTBDS9DU4F2/CCaRPoPQQ6OWI7kYY7g2SPKN/AsdSpAnk4N9zp
3TgeSF+933qWhsKj9mw4nwYXBA0KTT0xZY7PMTwSr+e5p6Qv+NV0TljD4sgfFOFv
YTqsf1kTgzHhh0ahCPnJwxD28DLl8a9rXlbyofkiHlOMjEPzDtqiTducgP8b1RKD
Qbc9BRmrdC90BW6EEEF8OUS7g0aECw8CaJ+ZBfNyfNqAzQ7XsP5+4q/91NRpxREe
IZIZf34OFriTdbpm0OJPuxdwr1FiimtH6N9lcp6jlXkmPfXEbZ8TGaLn1c4R2/Hz
wrslxFyMleUkOHfZDaqI2rl4qpIWytALYjemhW4CBkjZCeWvanAHU+OulasKKhbp
lcxcaiaeMHEOP8eYYip4UWpsfFyxx8/7WWPya0VTkmz0Na3BGZFB9r4CzpT2vBiR
0hBvzhlD9WfyDcnF/ZsqzHB5ESRndaVaEwZfZ2HUZpvjXt8830ztCQuw1m2u2PWq
gVf4N+FRZ6bD5SnQuMZx1vJgBedNdSutnf9ARs3RXdKkTjZswiNIDkkXjuFG3hDk
x7djx0ZKf/GDWZLsNCEu/v/PRZ1Dy3uXt5oN++Mrf8dHYWHYrErcHqQLftvMFPRD
QwupnF23j4p0QAEly2kcED6BWt4sC2du+XL9Xzhs79jvuuWynmCLaaGVbQRdHYlU
FOu/jjZqrbAvkooJTb68X2p30guR8UKVPsw7wH946mMc3VNrSgKTAYj8VTBf5BWA
wi4TaonZY5EmTAp0wLnocuMcLt9EBWubV88kjgBab/MhLEFwKtlejMPE3c0c+WD+
3fQvunMtMTVainRqE6g4VWFvpvgG4swRlsKaJFN83JHGLnCcxknzmEQJLtaGCIfz
g8cuXLB1bGSurvz/V9lGAee597rGBxXeKXBHS0essi3XmtLzNUTppPl+t1DfGdim
lbouwrUaa7Yw1jebLNR0ZmOPuxiDzTBS4CA/9+fm7fX8ZLskTBH7w36BwTxCFBhB
fLN925N3nJOBERcWwBuloq5rtJ5SWJcoWq1kdZ1oZ0Mzc8/Zpm3wvSweabxHWSWD
kE9NqJkmkXGdTFwr16LonDwWtYqEfmhwy9EmnQGfypOZIwJdjhDgm0MdKZNmOgt1
+90b0OKlWCRucVXEhJipNenlYJ47CmNXaewOvm6LqKErnClmYvrs1IOFFOUKDR4P
ApDrA5dkXkJGiVioWTlylR+e4Ix2ioyRweALFVNtfS1jHw1NGdEgRPy0MOh+1xv8
JY8zv61noLzEehdt81jNJgwJAOPDEeCK4ang2wr7hoLrygFvE/jpePhaseEm98kd
BA9/nu6OY/W7DQ9BEcwQ7AipVfWPlj0yBf7s/U4KxhHPJowcFFWRvzYb6OexXNNO
Nm06aJZMxsDw465BN8INcz04GQabzRUML52BGukLlqm5Td420vIU6Z9Vw2v5VklX
xcRC31zy6OWtvt5MSKubKtwWMQXHxvg8ih6Dc7Go+NxdfZXkTn0NfyzBjkwzTx9r
b4IvoYhMwGZ0BdqNVpPXKmEDXsrDpjRUFI+zqAEWcdELmsdil1zddBcATGiRyDuT
MGpc7+zKxz7458FaOD7CyOy9MVix4SiOPlgigKTpj5MpD7V6LL6/mqgtoCv4gw1t
maAlAAVPeCatq3arMmaIdvhgeM4Qv/GHn2liz6Z1gZ86AHmCp0eVENDTk7eLgllE
KrUCSlIYeE86Xf7+PgH8JkVvA9yIBocQQK1S6agzAUqWcrc4ln0XOM/Kqki9cFUv
EgHDz2/+I2lFSmLLob4stN37Nuqc18HflU4K884Zgd2xXQa50qrNh9ZEoXlA/ryK
0gRfDjx3FscQ8iKlXE9Kc8ajhkLVU+f8ayP4dZn0Dr+zYhjo3wLf3KYkiODa8XVV
uhBwUuGD71iMclsmv9Cwh4xXsXloL4Gbiukhx2sHYcrCxceolw8GR58NOST+SVgw
GSaktrAQbjNlxtBV1M0yVCPdviamE7kvBBY3dGyHHf/Xp5JMWfR54AARuSg/47qR
5NCdI6TYu3lqxo4Ga/hxYIM/pBmeYMArP0I0uxNHqypTq18IbpaxBlKwgX0/29K9
UTkoWS/WFx5IVwkEdSRhx/EqQ32gezsfcK4qY1FsXXxT1dAjzuKbh5HKVYcHwFGF
OOK0bJ7/yj50iCpDQpymf7xIBzsW4npwZbUeALGEOYvJrffvR7CkHkYlLskvHxcb
dN0sjiwfDz2QDPXQHglmuN1N9wEOPbg/I3y8FnvyjDvDPTGoMa8vtedDx2VP/Rle
lROCEqbkkLfCbHPCFm/6jiLtyjot2JyQ8O6bF2eZlGit54SMiDDTzsNy7lrcjaxH
cNogUZx7SEIZ7eKhWmJH0/rzqBX8xu+zfjRDcaQamU1OlvMsspuFXoLJ5l3b+amg
xdQqtD08Vwnfbtx55ev01GUIU0LWk6ot3wuHWedAsaS734QoX64VHs57rjchSs74
PVmjebwmXtSjFbJHlrFtffDwieLQGUVVV6jiSjuLXnz7ZWw7FUv/SgyF98EoU2+l
ejzuVySJmxa6WzNKS2Li0PNBuKtvKnFJqpfqeBmDYRlKc4OmItlf5XTJJBjREdQV
pHK90U7trU7yfpl4hSQEOMvdtFOcXEpxT/yekG8JMM8shAjD8PRuROAGdO8HsEkb
B7s9gqu9I9OCWEyOsKtBVqNI3e2q+9Nrda05oiW1Iql28z1NhjwYMPEUpuervj/Y
1OwWtO0BVnUHiG652BpB8JOlmLyPSkJs/L+byN4K1cBPBD2q45RrDrAymcpQIi4T
Gf75Rh2yJYty2PHqdg8F7od419yJgxwR3hZ0M7SHbzCpBEUMKeeZpAtEVq08peyx
PaUwAqslqVDQAfGcUS8Cix5avi2vvMSy7BTmC+Wt/VTWm1mhamDWkvMUaLFB61Rl
VckGrbXuGW/n+kzBgKovwPpyCPx+r4EDONqoIAkDG9/wTelwRfAGPWcvKt0B1v6a
K0VoY8KzLA18C7iDJJ70CPjvOJ6vAliJi6IMFX/JrAOlVAPNURWEnrK5kaVPNc64
wSjsghQ2kpTq+V3PsAgnXzn7f66XdoTD675AhUhr68RqVNrOx6xwCFZ2wRnufUsz
kaBxGSHNF6X6DgCye6Ehv0zwJnm8/At6thTvK4sgJpErT9pzpx7CP5txp+ZCaQkF
csrwcvOlOzFL1nnTkWzsQxjlvIQNTM1kKiAYpGXpG6OXthpkXXUUVQzaFf4wFZOq
r8PIAqQSNFI3fS2blgz70jdK9C0b3FTMMcveszoV6rui9oaDApT1iQ+CQsFOhAl1
PZd/CyGtLF7/guTCT4yErfbt8pR5LtMUuVwyHDpnrduYOZPFrQtPGPdqjNt+iR/H
d/OF00hlXRGS+1WSbCUAVXhgVCveTouIyLiDrWTWjHDd7blFu86hCcwxlM4kr2ol
VQPANToe7a9nsJZDN2Kx2pEY6aw6SUGkj+8R8J+M5u0FvXw+pIuHg3s4D+2iO0cd
fiaxlIDNt/xFzPQECLbyK37PGKvQOVOGzHSdK29Kw4gi1bpaFJIWVSepxPHqL/RH
ABbFrpCQh/T4lEIfT9Fhu61i971GVSTxHb8TdCz7LOd41BMNrvUBXCRnCbljXT5N
pTZeFuKpX7MVozmAWRciRg3NxI61Zw0UQqeD/bnd7cimcRv/TmwI3aBcptuzBAdr
PPDaP4h5jz2y3fKYKvIXDFCbmomAAToJ32oB9izGNVDZq2nlF9ylKbIudkpvsz4D
wnfhOs9K3rbD23B+yEk49SMbVyTI3bYl1xHkCR2sn+EXaZxMPXlYV44RN4A7xfow
I+BDwTIh9xC+UZ90ZlXxJ9YpJceyTeZViYwsFYYL6zrRhuwcqyyMc+1q0wWnY8+p
Vn9ElWXqpL3E52NTdxeuuIPBCpXPAdDk1NOw7hJBCdZvWIBHmQB+6BY+TjrPbXQB
+IZokuE8o/El4EK3g8YWqa+CZCh1zpt8CV46C1BqWCgSQDixCYVsEFrPQhSPboK3
H4CpI7xcLtYkhmS2pTzaFkhp+m4ynRCiNog9CPtGbHEb2zz/0Qj2BgtbZn6HkyBB
wxsZxZ3/thXmEs2UE4nIZ+MxhBUvtTHFnE0CFW4wIpwwSvX2YnAIxhqBn8MOPzOC
0RJCEqqZujtg+CfOHi0HRpI1iSyKnzPZqKZoVgThzDlYZBGxlACoaCi1sHvkAR5c
T4foJlrLfMgAarnmXK7FmdX1OccU3YiI3A0XDnL7+w6+TbD9l8nydJXHOj5Dtsf4
50L/set9UYW3/9MLu1QMszUBdNY78aJas5F2kWzXYtEfSgrWk3P7x2FRjHOhdgAV
Y/9yQyIMU6og/d/k/TUWZ3MMPXp3uLl/x4uvmjt9CwD9EAzHTQ3ESl2JMSpzP9fh
WS9IkZT+4psoSRoH43UoZ5ohoooC5QzfpmDmjG7alDndpxB/IHxszSHrGuuYMEtP
Hm2YbUI/sEv5YbwXYlz2l3tR4UOpx/u4OU0LL0xkYZTt3FYKC+jST609D0+zzxaM
+DY2H0QbBfDyWq/QuZRgzIdwHbR8mljCOJTlZv3yIz+jINXlgKKWc3kb+0JXTaWT
49PXNi0J8r+6JtRt+AOMz7Opeqh8+BVkkhqlJyS+WhjA7i3Wsffh7hFIvYRNXkpt
gnZ0i8aHrLniDolxbJXyKAAChJ3V3m83CSN2oMWvf6GwKP/tvSFLjXHPvOK9EWT7
H9CUl/1c46N5aGWWKCtJ8i4LLrIWQ408aQM7ueBYJARYqCAFSXv1qWm7oxJ+yGbF
Zf+u4VFML1Thr6+ZwyTEMo/3+fagnNGyAtN8ybAK4tuqueC9EaCt3OEQEC/wqhvB
cY8gXUS3qfbfk+yvZSJuA0VGLQwmi56zfLQ1H6pvtagfpR6zKSJa8Lr4c09fYouC
BvwJsYUvwIGOGAGpUIWbkrvT/Hcw2xxjW2iNaL8MUkyX+14/8soXkTQzy19Hqv7U
PG/4pn3T1lt3jLaN0V66uNv3LgzAq/GaRr3sHtg0F3DSY+FGJZmvhqMBeEaYUNaj
1JFZBzICdPwE/w0MepkG3cCQ/qtuz91goP8XYdM3Zv+o0mjnagKMetesGzKAPsrI
Exx6xC8Wc2cMsrKCfdMgt+DNi2bzGAS2hwrVLcyl3T7eB8kFxyXN/Va7l+/S+0xx
3K25903LuDkOKvBqjZXxjM9BsafThNd1SbUa2OXkXuIJvZWQlmp8i28hPzPdPS5i
Ll0kw/j+tBxjvvsqDapCWDsi/DjEcvt33ZYNXpsgRXZZfj6nJR3t1BEliua0xcZ9
lOk3IVP7vzDRvOjz0sCKh89r2IxYi0whfC5BlbZgbOsqutlmQJBx6NqbDoin1SF6
1U4AJW+7v+iK3zHh3McwWEyMyZePtIdhhxr9W6rFx5pxoq/1V+zIMYRO9SdS2qcr
ey/SNGFFYHWxJtAkmbANPAdCNnwmlpYF2Ppt7y8n+VZnziSh84kHW+BRZu1rcxiH
S1SnsZT2O1T+LwvikIzpsLcOFi2geKUMdJ0UVDirdzuEugjI/qaIbn59EiHNhkdX
wlHjXnvDy+gL4W5kFI40Gaqqqis2ElTrsLwwY9sLMR38fEj6GIb6rJbR5zqg2fbF
0LNLLIcbl+hRjXI0u8lJ2d+bKtDEXHVEhhlmvHrj1Jwq5aV8j2jcUiVQySd4fcKK
mN+N7Cezjyw05hd0yxMEcizoFnZteT3nX61lxelhWpoPmS1B6diXdVmIGm/hnrAS
cNW+q0B+E2JjV8tSQ9VK1qDiJcEy9nz4dLvWlJRL4h48Ul7wyWGFNx/vV+//9sRL
Mi9RaZjSX25BvxbeJ5Dw1erQaPui0hssvSgyWdQ+JdUk7rCpjdfniLuFp1wFkuXK
mj9ANLFMbTPFwEzei2tOHfZAkxVGo2QI1x0lfzvX0vsNPA5fq2Eg2OhhqpKxv5nB
gLiTyrs2MYuNvUwlIsNH+0KnQmgkyH0Ss6/4z+0tpXM4DkHgo4hFOsvQLIOov7zf
E2cJKMXZeq6knq/kJ5t4EZr0NJx1nUiOkbtVgDpT+35sEW1uXd0UwTsTT0S91oEN
rHGzO9GienyR7oSV3ac10NgMWlBhwCCUSxgiiQ/ZosXBv6eHFaVU5zzGmjgXF3TB
s8oRlMWD+vMjxJR/a/rbLd2p9q5WLDtMMFo0xO5+jBpfAV92tDovmjufMchVtrhk
gOADJ8oOFQzRTVmTz+6IVvWCbE2zZmVnXUL9JU7YmQ4Aqacy+zLgQCOZa2D+1x+5
dqHIaoebnTMY2WQQpdsvDsVjmk3s4QeNYTVcZFho+jKBDLKLbPaDeDmwHslxMbsT
bNMDbxNacagAioVExvb1YtmsVRwe2kM4gX8LuzBtOpOlcApVADSzg88+cpyAlqzv
3W+s4HCqetuGZynULdBrzt+OmO+2Ra+ssRmn+MVQ7fo8NZ20WfUve0HC8ZVQNv0j
f7P3qrS60sNC6kXsmPbCma3CGDhddspYFmW0OxBwz1XSJ3oCHrggiNoK7HLAA5hM
REJ/m+WLArx6iQXnxrvroHmVOpYTOg44XIWTEBUB0IPD36tNFoHQwilT62OtEHnl
pV10eZXCRs412wmQ85qmTN9HfIqoUlKuswqmk6RFYGdR3nFBnllDo8inaFsLlSnC
HTCUwetRTuzQVYs5a8UQga2vmmb02nCi5pTSuOfQRxp4IijcIYt+PfnwSrYUyC7o
beWJ4u5FB3XTDag3U/3F8LTm2qp/d6MhIzbHpqKbLfW6lQohbUiQ0a5mLh13BMYh
9Id7IGD3pz8h74IoVFAIdF6rgxtXhLz4ojKubYzjvTAeFqC2SdSSq8O29OQHQ/mk
+byk6m3kRZ67B18QZc5Q68pO9UDkRNb/yLCc0vNxB75dPEF0h9kgf6EL/iufpTN/
9h/VGjYNtjeP9rQwT3BFO/DaPZekityWDMyFPlpx4UBIbjRlaBHsFs0IawIz4KLB
mFPAN32pj59tlCqUoWbhIScKFhBu+nwo1xjQKQUTSK4yr1vQEC/RtenySXEv6G5t
wJgc7W/udUOjr9UlbTc/icnUpuPNiXeZ8A5kOz53Fw+1ggq8TJ2UOcGnaSHudZnU
K5a8qoYdDSGqMwE9qRfe1NGP8rLhgUK1APGs35MPx7CH8EH4Rti1NTHMExqYQrnh
2KPZ9Ph+ozwamuD5PX3mwUOT3TCS0QEZrNa3Ju7IXcWEcS4NSNjodVnDtg2oZnR0
YrKFv3DVMyDe+A0GO7AcsVWMixYzBI0+qrDxl0G5FNoxR9S1N8qDiyEelcJ809Ta
7Ge3gnqbGq9jppHLw+yXd7RQ1BE5qZS/v8RL5GJnNapO8XgLT4eBgQg8e4gxBqS0
sSmCRuZVuN/HuXARtTdPiK9s4PviWmO62AYxPcHpNd2ThD91TcDrYEsh/bozpVF0
ENqVgnp97JcOUrlTsfqUHNElEbPQ7TcZZfI3hcc0SIkNmGhW7jYhO+jNtW5eFh79
AvZ2BO35xD0FGeuYYzXFq4fYEOgruDmlbY9Iy6SjwW19vhEZN5kTcmDgWoMuVGIA
kMesko55ZBltos/iTuX9UCzUygMXkjP00TznTLwNz2O/HK0duuQQHSbnnsILloi3
YPrQ64Mmwty8l3ppK7DtmQjR57L2nVYn872iAGhXa2YimZ4MggdY2JYeK+lufavI
a4c5vf4gxCRGwcu5iOsdL5u2okAYjcrtQe+XT1rsB3nD4fyBJzhXh8EUDC/MWn55
f1JzjarBFARzehVL1SMDNxi72I3X3SR39IUPuxaHvd2bQPJ8VdxxNabnw8VvBlls
T5tvUJT9zD39+hL4gfDbzeKmpoCOdEWUfT6MkxzGd8xsID8PbMhh1w/CJQyDTBZG
xd1j+NorCwTc+ikaHYxQDNKSNZKEjpNKO778KQbJHy3QFPEBBkGK5ETB3trtTCfL
H+PaWEi5IPMgvmF5KWcnXLZBBdCOVYYnkypJX78W/NR+QJxhInec1L5fQE6HWKnG
JvZxBq0P+AwMfJR4uedl/X6s9SiXNow9aRWizImm5Up8ZrCCirhR4DBjmfaPrzHo
h29IsrMSsnp1hgrdMoykGHiCHp6yBRnoJk8VeAu8TCX2P8CWFYqvd1IgMMtcmjL3
82y70j2un9VdbVzCe8fUMDe6p5LkEOh7w3uLN5pYSBo4Lsn4kNeac48GC3+jPO56
DAZot4HXmMYE41ROW/CAEh9o/qZF3kMFqZoYv3J77y8dyb+k8+1yeAmVjuIFTW4U
GI7J7Jr0njTCWOg7sw/DxaHjgQzhX78Ndw2TkB2c5kpAdo+F+WjVHujoL8GL70jh
+NbCFHn7KG2Fr1Xh6DMgN2viM6iXSQlR9S0FTaU4zphehMuzQ4O4eIA5QQa9NGUR
wmleLP5oEnAWAMLtXLbh3QZGjfCOEqGdC4jA+3KnGq6o89OC2vv9RgqQRVv9MOw2
6AKpc6p8s8550ByKGWrL/5a+bsgbKzOrkPkE5oLP2ayrUhGNRjpZkoEaSlGczhg4
ZAXxznW9FUAfMYNuwyZaxwUn8XbFwLhdWMmfnGJ9o3KpDSv5hrthUZzBw66ru87E
7kBxPqV+xRO3vSRX8tucn8VriVIwj2MF2nqdDm5ES5SoEZX4f/N943EmSDRhwO73
nWFb+cDOx8i3XykIxJuCx0GywB1wSRT+0HZpkezUD5Nja1H/2oKixrHk3+40vjUo
PwDY1KUrD3ZzMdY9nGQ5vSeqCuZJWSk6p1lKfFxqFuLXi5I6GFWR86MQ8+4SlxL1
eAmJEQ+QJi764uEDI2xFVxD6mEHRxq3hXQj6ZweDQPSn87hMU38+w8+XkTTky23n
1DKNAP9i6tdTYqDFLGRvROuqEUa2WC56PHgr+iu1eQgWGCvSHSfHDv+24IgJi7za
XlFB7YR48UeFCAwLCvXxaiXWnCiWCXoSDAbnitjuLunO7R0heat7s7HhNHht8+5a
Ik5W/a/W7toFlw1JBWJ3HfnBLYbKs3850d7FxI4jjysWdmN754SMbM6y3Tg7xzFn
aL5yKFtHz1Ad0spTJwz1Fi0cERisBT1/cqp9fMljvmUFGwfM3Cfw4sQ4XxxXoJmH
nBXsRQ2AFk2bIoX1tNegrM/ePGsPvMlwDi3O1O3lWhTtuwXo+1/rCvh4PjqTW0d5
/8Yyv2q+9CzxxJ4C8bjAse6f48+Iw2F8efd/7kv2+m58+7SX4dUlt6R7NtSW/mG6
HUB+GRZxOlR4DIgAbgXa6N9JtCQzhRlkABlQ+i8IY7LMWwofbLsnrDj94NtDuWHb
dgQHYUcdNyIOFv2R6t28B8QCRSYvq/nJsAxOzaaIfRjgMi93elixaNGwYpJ5V/4U
15reqwLZKtV1RYt7UnQN+lP+yz7AbrOJHNUtYCPsfmGT3n3ibdW01FztNEdsJUMz
2Q0cJJpYDgckrTt0Zs0JMvIJEBfC7UZvkl6D4X/MpkvdmmZDpbexkc0qlv/CRFBO
VyRfpPjiUtXndizEMulVCT0atU3zlGqmU0vVKsZVBd3FjMXTEIcJwQVWFLCkqtP4
Oum3/9Qorj6xltMXJrEd7MlNlhYH5PgepWYmmQ17bxUKzirq/ELOUKquYEFsHRhL
n41OHZX2tH2F8ADP1ItIpeorPT0JdEytC3Ac3TEOiztBIpolxIN+mtqKUyLmPth6
+6V7AWYNjwDubAHnVcGO+JWzyq9a/vojA4QjEpg8G9t4bYBW1WjFXVbCrv0gV/AL
o6M7TtOvaRIspGxB6AUkANLmLavX5uroUkpERNxjI7w8UpuQ4lVP26lTLHYJKDl+
2yl8um+dmeCsyP0KbGXIbyrlezRHnvJO1ud3gNQq9ddcK0kkFbaEqpv5V1PWPilZ
F5SmwNEJ5nOxU/4SjJ32qvVblqpIr0vj9cVxmEovTE/wZZRX3ajD70nEkbczzk1V
shnDTi6RPBkPLf/kqfV6Jxiy7JqqZZAUVnId+2TzU/nnd9rjiXN2tWCF+52Znt4X
KTLe766AhYkdse2Wtc3OU+bMh5bX3S0lToEMQSeBKNr/FhfrVH4YGr62Ncs/FzwS
qnn0EuBR/EyFp4S+ausi9RR1TKZTjctCTAHBIPTqBnf5ySykkMQpes66iDzZBfFE
YVLQKrPBtgk9oW7vgUuF2iGJez+5vpeyaRQav/RxaPwtXVVIbUBLipc6LDtMOSVW
sma7ekIOrl3WViGEXefIcWTiOpUPpWXiZvkV7qvrh8Rnw7sm+ocPmCS7n9yhpRl9
DLhwVKwfdlFld1Be+JI4pODFgCVHM8okovH/wVMfmXSEwNBigNWiu3IGOiOU6poz
0oqHYrpslIlatzw96aV74Zoa+mxFTAxcx0zA/0XtbYtgS/OpKL/L+e7P2lIa3FG1
hC/OgYu2C3LkRb4HoLS2a2ycjtWp4lxwMpsA1d43NbYHOjPSHiHIS5dxr6Ld/CnS
4cRwYaMEJ2p5PFX6bSkTjnIwQq6VESgbAZ71qXfATkoN2VJaXrFdGkooB6EZxvEp
ws+nu13gDt9l+Oj2jG51HMIzHrTTmRQoH/ifV7bDo28LbKQ2rGuzkBgrs9vMzcdl
U2nWV2eC3KmvmHVZj30TCVdzwiwV3hadB/CScnyRvLWEzkkp3DiKTPrn1H2Yu7mh
GMgmn44mkw4at6T08WJYdnLn6EbZ23fclKvQr0M3Kko2f8uHt0cHNrllopxss7Nz
9zotj81JKrzM1ldXC4adhiN7N+bgdGIJPqUs/g8layrIC15PXL1jOlHBBtkSjRVm
6gkKOZ4xdDKxaxGrfBDGI1Bt7L4SRIV3Ep82O61rLnmlYss4lmb/etLudO1L2EJA
zwsvyYi/XtwcbW+ynd6NzGG6++v7vO4uaTnfLwRc63FSmLkgeez6ZThjVB4jvryl
FGn2Ia4a9Xzn203XnWGmzjhBda/qsbDkgmPRuKXhyhLjypQlFLNQm2Zg4HTWqBLt
woPERyCD5jXJ924SVa7//2wFRt5qmabmTUwh0PoiqzVV1FaWSVPjCxOZ/3gDOCpr
rXh9a4bo7EuzWm/kknIEzQ0tMbdYv9uoTm01IIXbvpt3A20zzAcmOfkzPA2vo1WY
875Zo4hXY+S/nIUKTydjJrPyq2rCwg9ppssm3O5soEVY/qH9XkvMvYcF6wde2EB/
nFkGXY8ROxhz4GJvsfKcLP+ZNjj47MMimwQ2euwMOUAszIVZRjAaUnthu1TQnx9c
4Eh2b12H61iVt1iIHpPImEpRZeIkw9+S+J5Vth+BuW+OXWrxobJ3PflTNG7DWBSx
p5Y3lBvl6L5io3WzTGLjyseW43N5pADJeizCDcalljn39gC63enyf6uBHQ9MSuXS
NwV1eJSxL1Zmcp1r6ug3s0rCTA0X9Qs/W2GqtJ9vD5318+6QEbr/18wEda7mis9c
42RJUp1VpoK2fWsPseTiNt5K6Vr6YF4uREnekw4g7wlBP1f87peRUvwBDUzu2mPj
CUAutY5x/4s0zG32/WmIrAl6Y+AQ4nWysVr8+eyk/ctvMg3kaqXEyqZYwHhQBq5w
e0mx3Ri1/nnfsbNTPoxO9J9Km1ThDs58Uic52DDB3WfwcnOp0pLRoxj51VYzyv3L
vdGHeGm/ZXMnrn0+aYS8FUdEQB5tkb/GOnR9oH4rVELOWC7q1cmssjZQx4BYnDTT
553ExjblB6aZlGG2CA/WvI5XRl+x1reiTQ680nNkL4xPDx5x6UtCexrT9sx+KTIc
ar05ZX8WxUtKIRjs40a9jrE59clYimd6y1Q1lIaN33v5e6miui8annMF+KV+BOv/
bJaMO4I+C9wN8RjvMIMYrpJPGAzD7DLWIZdYSC0MCZ66NrNUvWAH59FstNbFg5T+
fYSARRoJBNMcirwEXf3YVrX6IP5lHhmvv9V+jp2oj8T+eKqJhhF80WDsPa+Cn7/y
F2ETm0QB5GLSDYoEnsnu7iW1Q4fs4tCAATxenX4YXSOHq2vAiMb8jVySPePrP7k/
R+gAlJ2x0aZV3ogqGXUztHxnP1F1pv7oPv2r+uyYWhFruyHhAjBMNy/w6BhJUQB3
YgiGnidmz4ILVKP+xF5uXHvjMJzamhy+7VRHKi1QmP/gbFoUI3FzA13+EYtgx5OO
9YogbR8Fqxf10daPuDWtOxPI9UgvsMjIxF3dHT9r3yco9dGAJVD4yuOmD/zGqz+p
JaRV4x27yvbNDUo+ZhM8A98qE3IrMBRYl/OQd/wQrdcCidfIIdZBULN13goJ1L7+
lfFCUaghtKzqCHdSnGquvRVuwcpjljzFgF2lwxqGnw7TpBGA/PktsopE7xeJ9pJZ
KIrNgQfne/IdxsI54c7zNb0h6jIu5cFOMVZhqJgQ95ZcglDclEDBL5Ph1W4NNj7z
HuddjyusVmEkVqXn7xp8duOJxgJ1B8TXwWUewix0R/ZpRna13dQAUrXMTMbNao98
xV7cUoDwgzYQi+tUbP1KDW/PkkFhNYlglFhmpO+Mi5aDDDMOGxqX/DZFGY8TtmTD
bmV+iQ/pXqNFL2HTnC5eK1T0F285GE6WvceaK/E8k0lOwV+oWcrULXU3yMVuFd78
DqqfD4yJgBZfZvu5bS4IUEf/AfeehQ9BQW70oNDtwKerJ9Gfm9gwosZWmoyuREsJ
IfwvBaUCkkbqxxk4dHxy5aowHFOBAZE4wmaWcPSoRUU75l477zWzh0tnG0oAmkEe
4Wr6+FB59gWaJOMbI31dRbygrbTRrvp+r6bMRBnUQ15HJM17/igyK9W9Fo9coW5D
OyfeVQVZ4ZkNe+B7RKpGm7cyzoX/6ECuKkrGpvic91EmzYV+sCex39fzXKIbfzhl
5TcIzQS7GvmZJk0La37y2nZMZMtT7G29C8awVnZL6dPklYsICjSOhmUdJ0J9IuBb
oZ7wgdNoh0R1YaLxe955ZHfP0eFuQIy8u3c9o3ixdmfEEVI65wlgaAsxZ75i//j0
6Jv0X4jd8FYACGHYtgRyWjey5BCJv69kBOl9gqk9lpdbkPLZ/LNa8KM9FmN3rHHt
344kajPNy2ET9uSNqZULpp96m8dpVoljKGGFHb8FGacEoNYFDurIA9nN+x5L2Q5f
18SKwdho6kppkg1KwTVkvK3HRXBBvQdHCoHeKZhSHD8cCYN0Xw2F1B94qUN9kH1l
UxMbOOIZaPTneka8bsadFZ/uXud9ThqChkkwVwElpHrJDGTRWY6IgziLpw/e8zZQ
mT6XgBfoYECKN+zNpgtzICGMA7WNcztKUY6ix4Exnry47TEZ0lmu+4pmPpa9aYVP
tt671jXn2emybfJdCB6lCITg+VxkS+AsN4w2ov7fnjJF1bhMD0fFo8Oxcxe6BkqK
pOJ6fnbat0/muUf43+TGWDzBDiZU8ph3WSkQ9or0DyG8R53Kxvuy+bDlU0wGLQ4R
laMVV3PHoC9HsFo4F2ZCx0pIHCz8S6ityytACUiN9yXMicT3LWPHPm4URT9I0gMB
ddUEVIpC486RNaw9YGFkOsZFcwzhFYgVPpza5gp9FZQ/xYFHvmcwuHT9uNhPfdmJ
WXAFjz6AodI/ALzlFzXCOStjIszcCWYIU6/709VhiqynAkRnra7lmnEtM1qydBPJ
wD2VmktgCjEqrhUCzpRx4wYlCT74LJbmp9i86Z6+x3EQKKWMH0DHuXZEDZRAZAVi
pzC9BZUYli3/71cz7XxgUxlutf0qyrQfXNtAARyfZA1tEg4jiajsTerqzGd22MWe
7+yRZ6kwlxgF6k70CYRr21xHm3INdugUYpjmhxarDCj0HIzOwAxPMCpbPD8tPRzH
r4gNZ99lJui9VySUAW4HPX3kgPfdhDSbIeD300uOE0kcoau6olYXBuUOJKYAWRv8
qn6Yz6mBgQyp7yci/d+0QpJrficrpEnD4Vyd0reE6HymVJC3HwBwpJW2Z/jiEiD9
I2TyM/zfj6wFplHO5gVR1lxat7phuYr5K2X9txc2dzoq12wxFbk19TE5DeGKob3K
vct8nlovLpBXPyjCG2sNEnV+dBlT8h77cR0WbUeOc/5IJE6Pf2/0AWFim4wPwExi
m4rsDnKOl6M3GXxtR8zisiBMsKC2kFX2lQztPJ+wAYxI2tCKRHfDJQsPpjty/sZR
INEK2BNjwjWooz+TcDHKsyQp5fe8aMYvJdYyrlIWNtBnc8C/cpLp8DTplwRTD2mv
gx7sOEwMaIC47Ofdz7Tl6z07beY8tST/Ct7iFSYhanPy/58UGG/Yks5S6m3JoP9q
SjyzJShsdNCdgEk2Yc+mToIMqNU7RokAxTl3RHGYeT2DfHEVBgYKDjvFp/1jVXSJ
aNZUQTYpsLFtz+8DKTOSx/Es+pqixO2Ukcg5HYT7Ccz2V5X764xRAzrUpyroI1S0
iGC76NE1OdMmr+h4IsnE/CETIO9lBRdyuAea+B6xuKHgCSROAky3Ufrxl7YCP0wW
kadsfcxB/L4CCYr0VKfFRiRUdIWHLF6qKoSnUX7mwn1v2mVmmB5TY7Q5MZ6BWfMk
thFKNSQAHd5XMz2iHrcSumaqSJViWcC1UDuBDDeaXuqncxh30LyQJ/hw8p4sbgkY
HdfrSMjj2uaTkD0OS1VvE2OPeIexoLA9FaeROJYiHMisCCXNqblFTQwhZc3ZtXO1
yXosSUV3H4qUmLUQNeYXPGFKSzAq1I6y3YglnyeD1bOos3zo1bzyEhHCOCwHPAh7
RqN83mdoKQgLWvFdSFLgq0kO8pT745QO9AiabeqruJNdfH81wNKSc2EykcVnOhl9
X/DwhB7y0YV0lAAMNnfi/JyjtokJ5Agrn1yREUT8T2fZLx5XE2pDPyqjaQhPx2A3
jvTdn1RovTqxJv+UGmOo5GKJVl9wTZfsh8oMwjYPJBTc3Ha2vH+zCiiNLbSCWk6t
7n3aopV0dQiH7S2YTugPcloEz4oJEV1YcQRLd1viSPORj5YT7VA9BA0yudSOTSnG
+dpITkPUK9s2zpwBmy+rF5ES1XtbZlTjlUN+NoyFuNnHbi3o+gQdPOMDqgcstHne
9C4t7l2P97M3yp9TcBQ63Afsj60G4/z44pz+NyX8IOOdxAhceRnrJsTd/7u3vSOB
cbc5oTsSyUCsdnK90QwU6YCZmjvxng/s4Iu+6fp0WuUVyLehoyfzkuB7NS7AWFNP
TUpooudDg0wwYbkPI3o0+3yavm1vXesr5vthg7hyVB4m1YcawXdiEkzgqgeUR2h9
jzdoITcEmzq5vBEm38bWzMurN3LCDd7T8S3WsfkB3FdINVv2zVZxM7adon2wW+QV
iN7+Em3rrDnt+ES7dS9jrBHlHYO767kyvWLFdQZCc2yfMx4VWRFDY2Mi84/tyaGU
CE1kqUtxOvkzU8KXbvrlomyOp+hWZ6/H6AZZ78dSRweG1gcT0oyCmqOa0OcysrEc
7yWrna8cynLub+8jxscEPbh9QC3oxOzu0PZZdm+ntxiYedprydpmdi/D9nSrmQPv
DcH4XRdo6mottzB3Z3XJyhYCdZbL+BUl+m2Yw8n0+iss2aN9m8fzvQqfL8+RgZ2h
blBEbfdXUXAf7m2z0cu6sRXcj8X6kBD6KIXEUyjp1fzdy55V0p3NHrmYJwchl69q
mAhYjsURufaSzkeJT6c05ZeQjF81/AetmLJewUWVF6aOFWBf7t/DcqaO9sCS6dgQ
ZpaKsGQEWDENjiYpxUxLnJJ7Y31GGpXGLC/qOD9wqBPKSXvpXmag3OOF47KwOTQP
D56yp3ygAvdhvs+fFd5ySe3k7af8t5Oc5iLdlyyjLo2dFIMcirChkEeR6UW/uZK4
0hcw0VNzWwbN+ViGFlOUpx6uMXzHOrbz2P4sZNTigtjm7senmsb+h3GLa47whoWk
Tto7EDsB3xmBVtxReRuua/QUfQJZAuYC223yxw7Sa3YnJSDIKeH+ay2thNpWExtE
t06tmezB0VSekxw/TsnJhADBvW4GXMpsaC8MqRo7tDUt5cHuqz200FpCoKmgtc9r
wGvspfpxFS4bNUR8RTOR8C0P0KL4gcO7yy2wPlgRime8OHGJDOp5h0QkLj4mPtML
tr7a8ZNjAydQzF7x9OxYfbClbTqUDHKNdgaWg2hSbIRqb1yf/q6OR5OFdUDmRE6N
k7Q6RuLzCCaJHEmHr/4h5km6SWyWAZjVNajbnnHmkGnv5C0HL4/omQbHwvzAY3Qi
TiRE5nNQ0LjQJHSAhsVWhZIguq2GFZOOAo55kVDx3JtKyrcBa/uZizVGPkLEZVwM
6iwTxBhHJ1uBf1mA+aR+iEoVCJ+8S98FtdlyD5AKAUG3TV4XmXzqdmRsCpCoI10X
RzMhy3CHG50hy//Dz64RBBRbfVbz2urEIRldc5rAP1HUQTZyVYSNR9AZVzG7lOIH
JaRqEPCriSuSpS9JsMDEG6qGBb2pcSp03tVAXAEWZIw7kQkdxdB0yEW60Lm++JeF
E85nlKH+vYze1RyB0PIzG/bcdwTdQ0B8yzbwh53OHMDZdPG6LEUaYmSEWNHGmrp7
aVpgXjp1a6MRb6SBVhBCav+ur/ltEA/dpBsR4x8K3+Bo+/QNrrJB6V+dWctdZ6WF
riKbLWFzbpP2idg1akQK3maRssKhLNVJbXgoajffkMlrHisiTKTEQ5w2Hd7R4x2y
sPgePc1tKeQEPo/FAnNH3MnMK10keAaKT2II/kbhVIJmsWb3q3YHQRIFVsQkcG49
v/DpAulEtGeiGhoDLea9zlwuCFQzf8oQthQf0l9DK2cKVvmLUngRwu088eQC6yt3
hyQhzqr/t7AUwcNRFeBDn9i/+n2tNVf1HhZQOtcvTLa5aW47xnZYZ4NclFtgpCAu
Q+iyLbmhus3E2JKLig9yZXqfLRgDVCCOfYhDRQcjzMKujaV24yWq0iUYzF7II/QY
Sqtp/RsC2XUphLys+dR2nAM79jSJkIqa2XwWahSllQGXUmfXwIIC7VIS450BoMi6
sTidmUkvFjndKjcJd3YIkD+6bTR55s4v6G/h2CdlBC5DiH87PbC0mJAl6u9G+tSZ
KOmOAnAHXhDEJYF+nKH2XqkpkIH1alZqX0vhyuhSPbe/SHi/yfIv7CuZzhCEer2a
bb5PVjgaRtwvaWnjG9fAbH1+pMCZ0cKOIxvqYOQLfNtbRbkRYG7h5DNPX9iAVBbd
+YIuKhUO21sShSEiUskrbgMh+qNRneMpRBUd624aJ4Vy/BU9Tq7mT8ZHGAC2D2Y+
SjHxM36UDz9pDLDlIqNewJmP9mkgcreA3G+htHBXw7yePSDjEOTzmrBlHS7o3As4
Dp89k5qICHS0i0kq0i8Io4aNWOx5cPS23HIVwTsiA4dxIfBiNzdRN/Zkfpt7SRvO
6mf/PDM36hO3C4RCbPo9IVxnG0KzVxE8Zhyd1ROdTzqTLFAaPpGVugkg9pqFPT+h
pvrmDBdnoQCOtFaO51f5MxhTwYzE5ZLQ6zw6mdEsXH7lWko/uBczObTxro5LomYU
Agr4p+SsP33EUaSetMS52RMKJcXa4zihzm4lTkr9/dFN/BAHZEnZpCx5lqNqkmDG
Dw2aukNdm69/hjCaXoNgkSuJ9YEtiW6IhteOAh40kMS9DhwfeVXmMqMsL9jF7KRI
RQylvMsLaLbbpxN5x7Bzbk3BpTL6KVE+KaSL/BABDKgGlP9OEP1USTDaZ5EJ+qHA
XSg0s1hQhmylaQHDGfDBMNDdHnRy6GkRMDnaxtpYwI4WnRkNr7r49lIAUmJsrX5P
ftHJLbbrzyydUi1G3ukD0JvLPPThXJfe3ZPOgWPy50kYJ/UuvLwgONWhP7E7F3JF
ni+JpdH1o8k93DqdQpxvU9D9zYfUP77KpaKUwx7qstL1RxNrr1pXSPCQccmMhb6K
DS6w20lwfyxTMMXHVgVObG0xh0NQKrDgluQbeL/aBezqYxw4LFGrWNP5iEmoE6Ct
W+nQscZ3sZc5RCreiF0l7VMfERjSew1CT2csbgDGX7j4u+MHii+zywfu0gJm4Gl4
6BSqvGYZg2CHH4UzjBTmeEJGaJB4OdUuNrEfeOZGnvl30O2SNJUw9yeXaThQzAyi
1gadIi5gLREzHGPUDBfa5Z6J3CeB057JqSFbdLVUnQAxUkna9jnsn0ww+QbPwG9c
6ciwtbRuTD53eIGvd/BCu/mXKegzuam8cGESJDcheq0i9Ti/7SGQaIwKHUadIHPY
2vAAQWwfCTM/mb1Cc5j8Rd5GDnyhS1jWb7aNrq7NFVawOn4M9IMrtQBhae4i9ZPd
LMPQx/nwRGs/N6gXdWQg/5TobgDJiLyqkNJFTnaHJpn8N1pRAMp3jPVXkudyQnOy
hONMGVdB/k6MzkW65qZzqd6hxf15vOJZm+JO+Lnwh+XY1xA3DyG5CRRsdxdaFPPA
uDyHQm3rpNx/u+4VruOREaDjIf62Pm5WtxE4RMaDte9iRuVpcexvwgNcCAK6ViI3
dcJOjNQWCTD8+GC19O51z1HaOKSvXJdqPdNYItA0v97nEPro84D8SVeG01uGwR9l
UpNxSttxTw8qh3N/d4vQFLqq9Sjo3eAF90qyrrZvvSgBPo9SrCbsBFX7+OV/IYLV
AokAzlCP07wMZFMN99eO4YbGrKohkbN09FSssN3RSK8E9MIVNcr5pgM/E17GOSjb
pp4nfcHsnSQAb0lOqyi1c8s7opZPL4wfaUd8nRvPxUeAo6aQ5Xlaja+1T9qkbnrn
P4ydVcjhxLBd4XIlAq72uYPVyUfP+bTmcSVCRpTU6OCBIjTalIGJth5qDAqrWrUc
PPFXduulT454gkAl8Kedt7dHp55tT6EECOxJocGvJvZjdQUxbRm6WtOe1aIuSOw/
uygK7N3m5TypHv3faF0Y1UX2sDS2MXuQ3hlSmk3rtHDMaEiCXVw7yQCBbp7aKoxq
XjdEw2hpLSsGmJH3wPVWx15mK95IEWanNreIKencLDQ7UbTbED1mn/1QrroN0XKk
JPR001NYi+8ORoMfZFnql0vNMQFziy4e5sKGivPs5wiCvvugnI1OFiuhZiqSc0wC
HFFjVebLZrQ1RxzE8D9NJd1lxOJZakMhbSJrjKSo9iKQSDPY1W16wWt0OGqDvgIs
C3QS9oxlobdTr0WzqMImzUMGE4bIPopKaawXsWmHF42aGPb/DQUTwXKr2jygU/C8
+nFbxBvzMES7w/vOeP/Hkp+JF8xq1Be8bJOzJjiT2ej3MiM66j+SYINDvmUiASQu
dS9NR0WVVOcp8j8jOg4K7zsOa+k2GL2JlDhOJOxc+R9C50tpBaPHlAFORkmRA/LJ
lL0+0rI2BkaHNlFa2yqKBVDWwj/SaE3TSeg0NZ3puBu1+qUP3JJ9gxK0tiWnctfJ
5T+ELR5GVbq8/+cFJ4I9XI5FkOcwixvkgbs8+5ZI771kXjtzo/6gsIHe4aXoV/EO
p9V8cf6OcJTmqBLs7iETAN5rr61N0D3jaA2ULIRMc6e5Xp84GEYmeUBXZKSG0QoU
nNegp0gmfuUEMsUz3VShSbSLBkBwd7uYSN5CbhSRqiTsCVYv3o5FuzL8lc3+HAlC
kPYq21Z0FpqbSccERh65UFesZkpub+vFkLSMchEzIz1Ts7DpYZ9mI9wc5zcxIUgn
abhgdLPoWOP6MW7haI544hXwQWr374thPglaBffvcqC9uqWsYO5aZsT3FgmpWB6i
uku8GTv4CPM5NGnxL815QTBIO69XUY4gvCbIuehYWsyAXhuzfyBLqtfplN887bF2
K8467Qk7dp8A2MlTQBtS7VD+tcMYQlQmglNtttZY7bq93s5/Q/i71Ap55DyqQJxY
GY3IxrjSRGLQUf6ljFhyqVYvsKSW/pXvZhQIpINRhq5HfYWq1VOb/Yam3XUhBzLS
M+ZcvHgEZLePgVRu4bsmCDE/qTYNEZ79jBwyDwpWBs3kKpsh2zDXeTS55r5LFjTP
U5Z+sw1luAYbtMD3G2DrkpYPC8fDdYSIrjJy/oNn7pa7JOV1rkF1nRakf0rMnjZe
RsPz66+AfPRpotP23adq14dhcP4eQWwzFSUJS3hioqYyCb8uLDZbjO7ornugXDB5
JmQVUwz3ANqBzyyiTaR8LNKP2Nd2I1hiYBBCHM0q6y5EqmWiNA8Uh7dPQrYyI/nd
VslB9k3L2xjLp7QZ0l38035C75/OnMaQqgRVNzG4lA+LZjy5PumSaLcWaUHEilaA
aZw/t/GRhiJDzRbyJM47xES/98fFW0kreS/cH9zyTFEUmx0gJeHY2VwG7Vu7s+S7
7I6/UI8DJBrnWafUaasnMZG2Gigfrf+eSjpX5PWeOPc3HjXuyafSxraAKEIAXYgv
eknTkQOimH2BkB7oacVxgkOt923RzolLHwkVpkKOuik4/+M1B2sOJ0n80rPorBiY
EgyBDNkE1heESEoxsdTbD4qkXxWwmtpELl0yFjPVSiGtCef2xjODWfA+CSPCWWmM
EFk1SlquHGbU1jb+iP0OPjhq9GD8JFCZsuZQe8lwjfQP++Fvn/j4mcC7DlP/rUO6
aG+MlSq7Hh9kUSzxFcQGZrOiyBCgRMPUtXrRNNO4MGsIMB1D4j8KNGC6q87Zw8rI
g8agxxH8+9xzr5+sY6MQLUImsVjTjRzwhCyzHWeZtJ9hZSphl9TRgBYzTQiKtXGq
lP93TnALpgklJScRTWyYRgvrtvMPOWLv2XS2sQ4WnJ5Hivvjz8vsXrPqxbrzKfrA
N6rr6l9xX0ciVEY+o09VmyAle3f9AetSD+W1fh+anIN3ZnjDU4Y3oG7R95TpLaTh
mI4PA6rbmuwZYTfQLlVhTfLGBvg78TjIwjbi87uuscBWIUorbptbp3v9BgTrQ0/w
yCP/Hv5tm2QZIc3sVXrwWDf1e/Lp3WBntnrhUv5gk8X3iQZl6URQFbDN8YzbkGJO
uyYtNa+uCRrNNXdxRdRol+k14KH4JrxdtGChlWWIvtytJCQn/S8EsRJsY/5o8VkJ
S8QCrfMD2jhtPCOCq1RGXq5hHlcFEVSfPHey69kg6X2RSbwxm6M9J8RvXHV1mIrU
DxMDn467jpWKYOgKF/n6bCy8XSD0CgppjwlCT/O/BRsR9NwhRex6MF4t8hSqkPqc
MqABb3j+ey32+9VGZ7ygOGXQot8y607pIqThq18YuD2Q2TDqMCfJfaAhu1FUWBHr
ZxXRc7b7bLQjhbKn84KYvurEEnyz7fbt4V9c63BzxF3UbUbryiqYDzF/cdbZeN2W
oW4e7CmR64xG47kL3PUg9kG9DteHMpZVJruAGwNtbkv2+V2YXp1ju0XBg7ZnBIuk
tUuxz5ilGBSZPNQM5aZIfPpc92EcVRzJqU/eBhaH/3C6NPyi71n6Dn6JljdqQMBv
n2ASE3v9PQ9NkpajMj7/xpp9afLyUcJluxc4T5+9sPQYdicMHpCa4gCfKW/jpMol
VoC1E9NzYL2UiKXQI2K+Ys24L9C7t34Ksg4woXKw+BVA18UhaSckMSCHvOIbetSC
V6KtlTeox+qWivpWLGO9yB9O3WYCZFS5sFcKPwQOYyV0ZYnuvhk+KmcFLkvoxa1G
g4OfKV4vqVyWGPBGLWZyvYXNKlVMNH4W2U30EkMKCmPSnrZA5gOYhDHiTuT3UQcR
x4otGhOO+2AKPH+UEAwSUnh+4iJ8VifWXmEgMDq2STxkwdvGwx/GhdcW0TpEoiCH
ccSZmBAZqRY8Od4YmG4xqT68bMyg00w0BLJ1xCB4DvsJA4FKj1b9OAxSdBmPqaY5
gSg3vgZV6AsoJFBoJ1oomj8sgnJwHnL1BCgRLGuwnHmb+9WKNl2a4odcfunYKNx/
yrzL/i00tLvlHrjEXyUfo5fCEOjQYLqfih35uxH4tMQtKC0aNEE6oaqflWqB/pvS
rS+eOmXLcUb1bgYlMwMPrdAuZTkPZkSvfY0sD6TnsktsiRMaJ7/HgWp5q5Tl7o7j
06x4KsC3Hu6eTU75wWxjRUxSUKVbLkyVagSsG9WZLF9duc2uHjB1mpI0lSBE3Gt2
8gyOnpiFBSOzcLSwwL8QMt+qtYLxg6EJkEGQAdAdOzG6LVgHklDbZIi8TOvqffXw
Y3sIa5pJkBlyNt+XSvDanYuvFOcUm2mJieSp/lKsWlvC/7oEPxeCO83NKDWFzEWh
8QEP0FugUzMqWsTUxj6SSQ7AAeG+MtL2I0e1wJLrANjJT1sID3zKDBXyvz8gfftW
tzK/DOKiSonHyqm7MSFSSrh8Ys9FMSxoivYdBh1eQZxjAl4m9btUttGXJbcNQC7J
0ekB7Yp7bOYhgN9pGhKxHUDcg6VeLLdtFrlgDJO+EEVk10ZEFXrMJGe/ekgebcEp
QT0rw1jSSroeEUvRhMnwJk6CIBnkHOVCXD3LafrosOXpSVEccceQDHrkSkmUP6hT
2Mbn2J69qq/bxH5YxyYRALkeaKRCJ+ntKiFrX8/FJ9sMFb/NzzYjS39UB6PCv1GN
r6OMbA6EjnpfqNZ9nKjfUUnbazUXF42QLjey2NBueRlSVLnpKT0N0N9b/H2bV3gH
nrICRphButiVWU6AZj3EK0kiUuxQm6l9YARf/K5/PZdnTKZNh5Rj7FrWZ4QeqSDP
vwokF/4/3y5mNfA2cO5WUCwKXT8yO7jDUV/M2dk9En90jIhVIuc2v4yanl9GrCsm
BnV0kW2/SexyTcxEbFFLyWYVQZKc67YZVyL/Teqcsk6rT5B8OuvOpc7yXU/EpdDw
+ch0Cz6QVs9SBvk4YpKH1zj226fY1oLFW0LKGL8Yx3azQxiS+mHDTnJlVruaIoWG
PlMdoGmn1YZdEm/pWjO+486KbBFwmcbd1zvvVN24GHUKR0mmP2ToOXEjiYepf7xp
iIgwEQeqI/sxv/J6LnrzVRv0zVBArU/FHd97WL8KAUPZPRFtFOPxpMIEq+4Y5oX7
lHLTuA+PBbT4akwyAjEZ7x+0onwiIPOp+Ye6dHazI7lpUpxeB1v+V+KNvBnHWhek
8Y4Q9X5VmKpOLxrtlxoU6wYIBRHyyNkyuwLr/uYOkJ3qX/yq43oAscT2df/lcvut
Y0hIR8J1oOiCAHjLlHfZGBe0vw4MUF4cTXWakTVpN3GcEhWFsyBDLGu2MGLFzCm2
5x7LXJQpb4ltbmepjvdJJ2FBSIqSLHXVIBJ0wnJmABA5nzexfnkaUp9F9UDium47
xm1xYTq628xO9R7TX1eCbInDaR5SKT3usDczl1OYs+Vcv30t+SqEN6uCYQWAvYnp
2bCkb3j1q7IPr72Jv/gSzt+qmXf0cFyQ4P3IPpD8kLkQZNKZTwYQQOX9YOw3d//h
9/9kUZ11kAwnyWGhzX80yL/03kkmWednGpF7tSxHqmclBnETl3TeThtvsMhzvaGh
eHYHP9FPPFw6oTynptLT2g7PsjnARkAYzHWKgMj8XeL5Cb8UlB4ojcExk1VrDCCz
+6YLnmtcb5zAtolBBCC2qyi58n/NSG6LFTgRiNNNBcSHwLADBGBeVSdsbv5ZCiHf
wU0nSkK87OCBLqco+NpkYWBhO4uo6DBpguCHL/yuIq809WTw8+dwJiLXubhrFHVA
E17o7uqwakkYhSltMLk2h7g3DX0/kHCrm+z1RiDLPkzGFGXUnp3WcEMrbIClIVhk
eTIY1Sc3bN/DkPZ7/4AhAPK7NpKuKGT7j+owBqSusYlmDDaYwQrxd7ZinWRMbt3S
b7ZC774woBc8aDP1qA+MO3i2WqcLGDwAT3vvyx1x5daNcDq0uDChlWeFXlOM4ge1
VscOeU1jWkviA4L3NIxHkl+nPq6oahpW4TpMdrKYt98spSOpMOZPK5DoQl2ogV3q
dSbHH0231ddmyykfVWrbyukN6IAN0g+878xpdEMhDIYul+6fmprQClJ9WhISR12v
F+kWepMwm5iHh6VhS4d5RfVWZUBn3O1FVMxoShDqu8D9qjd60iJcryb09ybFT8KJ
U+O72Wrnq9TqJHAQo+Et61v+spOeXn5eNcaWFtmRZfx10wghN+ymkjWw5uG0Ft0w
+qKEbEUjR3Ff+ezccxc3fkJK7XlFo8mo2HeN++o7Tm28ZQ0sUd0kVqN9RPRjmElo
VduxKFhpO+dyUCx+Sah7cFEVRJp9Ze6WtbwbsZlQp9ytLAFM4TATg8cjT3pP7NPz
BPMUwxkepXnfPOse0HS+xLgjvgTok2JkAwxWAFQc9tveuVZ4Mt6bEFhYzGSrPSm9
NvpQyBPyvzIiuyp7OHPLSWRq05P7KfrwwdyNWpTNHOve2mHbSY4HHRXKsy4Ennqx
d2BApADnsjMlDoGIa/bqpNUEn9enji6cBNGWRm/JK12O1tu6bGNBsjNzYHsEwGqL
e3NklTpHbw2MjjJ1EYZ84MOkryJaI4jafdC8nbKKv2nqOfI4NNLuQdIvCu4TbnOy
qUh68/QgQEy3V3GSc2qf2/kJC19dVOCHIyIl3rLQv3Xhz/CAyYDfqnsityjSdkTf
HW3nTFi3rnXxG7pVqhxfKLyb17XGsrgihwHnie3N8vED/VwLDL14STzlqheszw8k
S0C1cAWUNXfvTBH8agepJM3Z0A/fLzVWTCqIXC7UHHDRTu2Xn5lbo98gTsVCQIq5
P/TZAHwq5RLITB/mM9mNxn3IGcqcCtMwLuGEXgJK62uEUJN5JwJj8Uh32WPc/BcK
GnPAY4yWgifMrcgHJvzYA5cRJr4WO/lq0hrK6jgvqm6DrpXlkKUQWb8qqvSbJeOx
0of5Df1f4D7UprbNwJhNoL+as/G2sAbMBcoPE4Os89/Zj1If+W7V1S/r3klIXw6i
2GxDdwfdH6/UZA3gIwKklKgLw9iUGj7LOkUgtP4fp0nMdmWMhOyCmZe5TZV0xAHD
rOtyEKRVas6JARK76VR5A0rX6nYtCL8Orp9VEobsRmAtRrMuqYZHB61q2BTLUqFn
DrBKigZO7IoU6tWjgY7ihMmc38NixNRI3tEfaJBKi5I9GzvnpZSYvohQMsGbAa52
5Z0qO51vpXS6oFM7KcQMBdPgE8LOWMaEU8hcpwiCviTKOxM8fX/UeBiu5/8HjxYY
T5rHqa1pp4Vrw2yHW+r1nG7kJGD4pi+faX2WZeMazPXuNhVEyIOx8uohu4yTgmTA
ZvOH7u6u5wfgvQjnHoE9lP/vWjd5EsZcWPtUclSByst0pZYxSLY+UPUyyOu9VPYX
3wTPM+/qVJqm6CI7jSE6KTa26WcJRQYRm7z9l3bEB5j9gqqqAm2Eoxs/mD4Cd/c5
Tk+9xnM6yV8imrXwhl9eVrCgh0sY2a1dAroLPWPhhkCYHvmw6glbC7eOB6QyIIfY
OCG58nJfVGgjekP84Xbb+uhmDqCbw9nw7dSCMixIWnHad0AU65exTH6U1uPWHQhB
ymtcl6Xod1jGZuMs72m6Riqo4APt30IQfvU87GNqigyo8c+lC+KvxgL0q0YOXFc9
ByuDb1Mplz4HsmkfWmhttl9tReyfyXwNK7HhWuV/T5vzpQdgv/G/za2pKFR6wQ+s
JrPnjw5sxcoTc8x12rOiZRMJK3ERh4YFIl+CV3pFy6nJ1YLQWQbb+H1CQoIKSnqk
cP0rcnK1KQB5gyUgRVkC07mD41CXu254viuJZ4wclkMupdfpPSzlmGSfjhUxE3Hx
iRGAWxSn9OSR6R4iihe/LXwYQ6/K6/YFF2oHNYUOuh3lNQCPgRAd0GqCVDQhPgXd
AXHl4ROuyFYYrnkToIP+rj+luEmnPH+8UmGesyC3gbo8F4gX9JI1pkfEmP48zqhW
TcIie9Illj+ixbEhXHQvALUMN07fiOlqSM1wrd2t9JxRzPTP8hLLsvDLzIe4gjYF
HD1ko5R8viugRDLMbPvgfWaum4TGb+6bf8dK+36WGBi5sGzUXY1eEGIP/RShCzPM
EoMcTJXSWE9IkemGS7rOSmdzaKdB4m93lKpz1xTdZsI7iQm6mz+x2W+GFjuPNSzD
1qaYA46sU05llEmqYz4mTDMJ45LpgCyvKUM2gREwIK0wskg0E67LVG8/IyeKoOCo
6Vo7kFT4ayQ2UCxYBW6KVSrMaSSk2j2Hgm9ePVX77qnQAiuYKZZLFWiu2c5X20JN
EuaEP+AGd8UaeQCgzTS/x4x+n5t8/5M3A0Jtei0z+nNvwZ4whpYHxnGHbYyJnmXv
vEtcpp6spiFsHp4ThqH/P2Hy3e5ULbaKR3BSf/mAROKbOXGjebZXKlpmK6FcINHK
2zyFcXdtuybK55tLUw+LhZq5400E/+eUbDfZEPxzrbRMM0tF6UkmeNmEv2X8lktZ
0YVhlhNZjBtnZ+6R3MEU3kqbowut+WXrc3M9FezfEBvCZbwd6jzw1BUcfUwnHmpP
sSImgGxJaUe3dBSJiIXCrCku4EUwBc0JbB7qGTIKH1p0Y3MkmTx4/cLYrS9N84UN
FVDH10rBkV36nG9Zn8fysIEt/lM74QiQxva1ppqZz8oFpRKq0meaf31fkQD9262M
fsmA8d5tJqA2xsUmPxRgIli2UnsyIPgoa6NobYaWBGDTFcFylXDpZNJDNwP8vOkp
xKmT7jlMskM2e+nDHr/ascyesGKhc2CNiQakucKPWwt4rcRAVY2iHZmy5ptMZ5oL
SL1dFJsgniW4uMD6hJC56xFa37LX8smfB77+rCnTuzHIMVAi+qqC5IjYexn/esdG
NGDlSPaFxi/93kgb3z7rIn7ykPVVlSPqiBa03c9BO4dWFc2J/TcoW9mjQ2xYMivL
5ICnTvHD8n1bpWuWjKCR+Q8GIeOquWQk9+IcUUbCVjZCrro7eGqzgN8dB2ZvQb/X
ErMExC8NeG67HNikr/B8ej9kNuURIW2XXSfWkxKnTCmQ53IOiBkipvaSS3JCXBfO
jd3UWBurvwFc62le8RmtJbmkqaUqZSyotuZxOg3Sz72NOo4kPF1HBBTHRDcso1Ln
Wujdr+mu4giIhoEvhibH0yllzDPSazz788V2zkI+Di0A+QhnHtgSj+W+9aodcu2U
HRJrL8w2LKtt7cG7rX5hzZzYrSkLoKiGKecVZanEyyl3tyQigGR9pw5h9o+4CIEd
kXHc5IrEHCt3GBbWuGsuEkP7dAE/DBvsElyA/00t1icGQK8U2+4tlTTdXFe0EVPO
wk/8DorXIsyrr3jpLxwdjs7R2L+Ng1PKpDpnyLSfCbA7ap69wCbtWsP6Xvy8umZ9
XpHgi07U0jp/RNUeeznP/r5V4vTWAdAnDurado976riKZCjIPt6KM3+rN4WAinXg
mZnJ0C+giDr5zQIZS1x8Etr9vaNzLv4Ys8fW7/93WGWWntmEU+oC/MSV+sHwtBb0
0GBVkLCa3MhV4Y93EMFuHkgv3jOD0su8Eva63dX/0bnP8okv6VXhUaBExmWgFdpX
DG7n4o9FX4N0Q1Wc8AKfLFz6QFHktwX6rP4EkfEbqN3pDDAXstAYhheaV2HxyEVP
Pr2iZydaPKdXI80xINUrv58P2MwxE8kCAt7xzfkqt0sLhrpj3R0YkxMxoGw7gaqy
D0BxnKcqLxHTN/rSoiRQZYmuaaBjOH2WbvWfnoxXpbww/ue6Ryhwz+DYRrUI+dak
/lz1F882mjT3QAqHepz5/PySx9Ua+8GguBIyvMmhHFQffLeQMeG1Qmc7JxOFFSIH
/ymdmuWPIUjWl1nr2DJr+v9NA2NcP1LqB1r66BHYgb5/SPn0eZLO6v1eR/5Ecwh8
fquMmQYMFcl5p0X+dxENr4b6PE1ZkiQ5JA/4rWNcyHzJexhIzO21LLxxgVsxpAwK
SI6T1XiYTiz2aKadFElOHEBtJmd0TaRQYMKdgKVnPG2vp3XVLcpkumY87SlTeRIX
6jPvfDih/0z9gV/MLquzqIaSkvsz77NmkzPkrUX/XKJlvdV8iLKLXdJ3YNKy/8SQ
u1UqV1ZNiUv4imwcepZVzi4kGMGqoWo9kXJNNusuqKGHAZmLsV9und1mhN40RYdp
0v27ZJUgcgu97cf7tIaZMKAMIa3oX+/xPBptMhCxzvhS1TrfCDcrVMjpO05Xc0JL
pTr+K4Zh/8A6XYFtkFxuBW0B8YizsGDbaVS6AGGtm1QGHQvUnU/qJivLYSmkYpOr
nHVBX9ESgTHB8B2n+JV/SHyWKZLasWiejr9mkGJ9fvrHmMPZuSMc75va1UGD6ajg
EOAC/hCQUOC0JF08bFq8YKJd7TP/AU3rhBsO9vay2sSjeXoiUU0o2WrKHYj9SOev
bevcWydxknyv/zCvPPcO3PFpgVBS22P+oe1CssBhHnrNlGFRq64lRYEEEFWvllTv
S888bsmMWw5qNbz4Ti6l6JQBLNSQKSl9TZICj3nNbHM5od+0JKPtCj+R+Kxu6MSZ
GmGxzmxttBDeYBo1xq7bT3pUJgRF4uK7M2mJuFKftHuSNE/th+NkKKjY4jF7r428
TCzYR5c2gobW2uVZPljkgsUt+mCrpIMSvubMNBgpKr742kzrNAWCuQRMJGOfWt0Q
CToDNMnz2G10gjvUxtt65HXDAiM3AuqQC8aUEBxwwzjcqQAxnIfiVltYhKcsE7jN
pPaPx+hB3natcVtDetCp1xh3RrcoJWtwbSWUIAHbdsNbWovE26/yi33yIT+LsZCV
RsL7HQxjfQrH0z9zbwAZywyRiQ074ZVNxVEWSQPuShtxszYDjAc/Da6UiacddTfx
odC4mjYHLoaw3Q5+J4tXWsZRy4eMjX9VcLOU7SREOsr0+RrcZZqa4eNxBI6p77xQ
EHI8dqNVSY2MG4R6C2Aw7d1ufiPc9vmvP5OG7OLyQqL0CDkNDQN5m7r1jwAfcTzC
7KxyIR7/djlAF1RDvfM7BrIkAiKMGLgdH6KMxQXuqUwPQgYUNluERmHYtsZir8EN
Rt3kQ1qINfsbW/xTDmz1fRvol0D6nNvSHEfhA3MeTIKIb4TH/+jsS70PUOJRDYgP
Q9srhFAEgKYGPdhJ4uxPgOqAcJ0M6XD+pQkAFKdIbReHQyLDpf/KvdK9DZdzl4my
VicVqFfZyy3hpWQwgul+W4WWfw1gWv3XImSRhv6DJjuqFYMrJ5YOr1S0igVTyTpB
imelY7n1Ljj6L9ch9L5h5qTJXpYqNBmKkP3u1RA4Ee+S4cgBWJ5Ke75uu0rYVsOU
4gyZZt5CbPbS9EyUxK+ilIxK6M7Nfpvoc57A3TynLdWpCWhRi9Pw+0CgjT2bZXj6
Xm78013VMnQ22JXkTZEqLfqtRZtrRj2zOiCOzidiKMM0qwEW6opLGEzRATevfXc7
lLkkLGjlcROigyMqJsfrR7eKk9zZwVQ8lE1YvCm3UG1PRYZLpgux21VMOkN55IJX
uEOzAWE+aXhi0uDMGOPKpQ01NaXQhQ75IzceVBz2tB6c4Vui3WhzFhDPWhYxVYAg
9BJW7Pg2VfWDwOTjNuN+3ESptcyjHfsuT3JcJBPkp2tvtyQUmgqCbxWIw0Bv950R
uHloPITaXU0IaBw4SDPFwIe8tr1zlXZhSlWrab4MLtp/WWMM2pp5I25h1lgFperh
Tm4jCj3iqYa3Q6ZTnf+nN9eG25zdLjmaBbxt9+BucY/Zec7lBniDZnlOqmuKX4Oq
FkePPLxhnloZWBnkziSmsNTErzAMk59yHb16rdi1rPLPOgHsbYUzGp9XfBFST0t3
HVcWoxPIlUfAQ+mNw1r+DZ8xwBFP08tzPZ+3QSXsYZ2erFA6CDWibnAnQNtMopGY
X51WNICNCHUCiF65mgt4n1WsIlSo39i6HLNQM5aK3VybEPXPqwN+Y4DUBIM7gW3C
0NG+ztjxSdl3wbjVOst9EG8iN/67dZBjpRjVNSoJyW1BJNlDcArhupmZ3A8/7iP+
tSc9437VFmZ/ajsgT9/SHy1jf5xwCuDc5ktqS7FlxA6P/t4RxgAcAGXuHv0xB+bK
qZ/EwaQq7xp+HhIZpfqzdsYLAVKEPF18sbe3grjMJLRuD8EONUEWilf1YlIC0mVx
DZ8OTKVp7W0LKVL/BTILVr0QjfyQLmZTjK4FpZfYyhs861ULn18WSNDDBxZ1G17w
slblLK4blMoOshrO6PT9ZC+PzRjUToV74YHqQIuNiFD/OVwZY49vSD1tqhYCRd5Q
9EI2qThv7P3CBVgWgEcyxtJM4/25MuBdZOlKMB5gyxXfIEY2PwpN1Mh6L5igFXq0
NdKOf5UtN7HWj8MvyLqcN3djo1ITvGcrvxvEZ3QBxXNmTWbW/heKaIrre6mN/QeO
xCypVF/PFc1sg2QFdqFDjLKgpuxqp34Qhk6BI1aW0w/j3Ts7AYnObHY/jEBfGHkx
CuLkH6flDshLeX2KeO6I7Cc7sW2pOzgqyFSqzDRz3KIe4mz+ywfog+tBrLaXVOaD
wAFsfQ1iMOMNRavbVqfEVQQ6PsMwxWPCq011CAUFIi3DvkWdXsn3sS5sO92d7JqM
0s7q1BjLJH0OmB8wSHWfJpw7bo2dsnn6WYZ1TfRaTQPvhp4QPCxIovkLEdpGpCYn
dcJmDke+p/Em4f2CG0Ew3oScJRKMxvK8r9xBl+nMnSWHUaJrjts2+J/lX9rJo+aG
X3iSglNRANmnzr7Y1qevA8p+0S2SCIsJ6/D/UG2dAzrVPJh1bbp2emDKNFk+I4z1
xh3ROi37/QYXhycfC507jvBAVQmOuFmUY3t/23zvkkJ/voalfCyzUL+XordGc0Ta
FvIbrnDeph/UyF7vgMDV/oE8ZCA7VTyL3Pb9R+HaOikd6Ur6g9BVlesUBZwYE5rO
WU/sRDrHbU/5yyO1qAR7sKWoultG9Gkni4aiP3TUr0sRSG49ZCGMmxei31VhpwVC
WHJSZwQMiflzjFdplaSs/we4bhKWcaArZWAqeHAG3vAoz0mpKKnQCYydTzfa+YsS
HTlyhshxOtR+4pT7RzlY6d94hYnlJa4PyGZMjklJU3ixOFjmdSUG0XX+Wk7ZfzgY
q2MPUTzBR9pz2qHR8Yqnp5MExKrj/gR0jGycwrJZOzjS1yHFkbu1qmli0IvMgw+M
RO8EjUCPfmvsZFuY2caV5AUC8QVInLbiVv+NE7o3FBgqJkYM9IeDiyTxz1PLRfWn
8ethhcaCfPrbRpjouCfIzj4BahizJr7LAvgsI2erCdPKxJRD1MQuwOR+IKosspXJ
+50Hzyithv8gKVujhZotjLrRqqq7NcrTEr+Gz/k5junZ07E6f0syn2MiikPmZJNo
ldEVGHddhAUcaovqtdeHR7GYNUAGM3mAoT3mMRVcNIf6wgl7YxVYvBtR+tQ9fIYj
aklr6VtGoNQ1m0xuX/u8Otmd+DRiU9+ZJvuwHXvNR8MXOyEYswvrzH4fNJZmFv8c
/Ri8FaIT6N8SZ246wa6K0Abc1M23YUFZgudHkuRAPpybIXAj6tiYKKRy3He+tv+g
CRIP44xi3BSMd3qmrzzTXrUul0+LZSj3uTu+iIPVrqp4776sk/6HIMGbOk89gPQf
2k855JDsZvc942UP8f1PRYVVwQ2PtlLIQaLjV5n9P9Af3Npt7xQR/7OW5kfs4JQV
I6BLIPWvIJdkKXkt4fgf5V8DFNsFgWlk8JrLeCjOrt2SSQm+EJPc4b7FTpeAVqeF
iMObCL5CCk0aMGoO8IhdWreQyYmaf80c7uaozfNZhlork4UUsw03NlryfFhLJNKH
c8A3diFw2++yraVPP4T9wc10hoP7N1rTzD1HHmIyhDFeDSDdG8YKGcttEBCFO5wH
onUhZFO1YSn0WuR3egKzkda+vp5RSqqhxHpiD8PJDtEja7KngjtQCAVhu8jsY1Bv
RVKr/IQWkrJbPkK5KgATEUCUIdyQszDnoMmguZpns0t0XY/3cxkt1FPRlbjT8nSo
WxPg2KgW5QtMBQ0Z5pIffgCXYXOvwNWugzul5kpGEnEI95jcYzVaBN3wdEahhR3r
z8+urHqkCJt7oAcyEWduzyGZcUWmLkEefD1UmG/tIZME3todnvyejezdPwXvTQXr
XUULpCGBvGoMLujrvDIYjYtU7FS/S4JSXFWDUDs93wMh++XuU9SZ95Sio0v2FFq5
aus+kedxhJ65VXVWjgNjz7IEWu0V2YeIGkU1KKOKtkLCz0eF9dL4HXUJiUdtWb3l
EuqyNsbptO3iLTOpVrAqAfBEJlIUjbBz3rX1g6ayvnKeO0icjuWtX7CgY776e0Bm
K9hH7SScg1rRB5/LuIW29X7cep4/VRKqORX6F+IV8ZuAFIzCRac/VheuQR1rHsAH
YrV1EMDYK3pdFpbx4FqslP3MrNWAPhHMDSWXzrqgIlTdbDORicXkYvWk2w4G+jPo
d08tqITBi7dq57nZrWRS1f6ioBeTg7xLpzalTxjUaTg1+HB8n0o+xVr78ZBnNcxf
9qPbeIAm+LEEalbTZebqUNSQ9GoQqEd44+BIOFbdX9QIsdVHjEJUf//cbv+mZyfF
1qzGZ00Kj9KLhUpP0HEBJb2iPvmEENVE6A747ZLmT3sdRO68tcxrHHMJkljD5p55
RlsO4frJNtm/ca2ocJBBhRGu8jXth6RYA86f07BANtEuqbzwHUQEGzzkbndVmrWX
j5tZ5pZ4Z6u7N7IGUhf2JgHR+pXgXrkIERogxpdOWW3bFkKk11+GuNCRLy4EB89F
Y2Hx7+Wuru2zod74DQiqLNv0PlFxx27LFnT42wKEN8CNE2SNiDW8v0zyQ3n6hrW7
ag643qQFU384D/mB2YWGjhTPC2SB/YfZ6TrAipSoIMxsUTnNOl8MHjSw4yTlLYTx
tOxcx4nn2vF7QdmgxcHi/diIfZePeIpb9xK/3wtvnnu+MyNQfexVQDSif+JRV794
V065ZmDVdJoKpdV/h7Z+xM6prijWm2AfgzKcdnQSsyjkDAzw9ud1KqCRqdh8TJCp
CTkEigP3bky/S46kQ1if0QqnGC9TNN4ljTJ3uxRzG8qTvIPf3I1zmXf1lx1EM0zt
HjG/kqFvIMsfkrDy1zR4N1xKB+wBiyDRmrxvHBc3N0m0HloJY3Wu6/nJ/XVM2hbT
oeoXd3hQIJWtg01OLBsPjpLlYgJ9W8MiQ72iId3YkT9pHPatcSUimFvsN9kqE7+K
GCwwudMnzYnySs5tHEX2bzkdl8zSpcoZGbsp5FFdsrqPVGn/Ght8Y9Jcph50ENDB
vOnRL8aZuavoTBMCHUG+Xu3edvtvQfQPq66I4xl9WB1oicL08oneJwZaAkzMldg9
ZhYHzaYeLI+/6TfkBFTBHIeKDiXFkultJllfOHjoQ1s0WxEUFELL7oDIrOHtMQeR
jB0Dhc48rS2AahrL4Tm3mIrSu3zOmg5CxRXGicjhZomPzYnk2mUEuh6ei5w9Nky4
S0fsJxv7LJ3kl8Tk7B9Np9WTdj0fgqkF92J1GnoL0ZO0BjamRyRAAhYqaggrrJif
BKb04Us+OQousppia8q0whov76U0NZP9V9bdVl4iHXZFhSwxZdNoAfIJ/cm+LYLp
Hn/w2F/bJpHlWronpuTCk7Sclcp9BzXgE6/4/thbK/g4CaR4pVc6CqK2Kv/O4BR5
l4z/KFNA2jR3krUE+C2nuuLSFzFxi0cjX5jXdryAR2QyZ48MHFWTDzFaZyfThtDU
2pLlLx9YlGdW/CoFVn/SNxzz01nzkY6LYEeoI+jsUOZ143J8bc8zpjnOYb/G5D7J
92JlJwYx4pY2JzaINHGHfvB2Gcuug8YNu08edFLf/bnBrHxJdW5CbfMwIACFXc60
7u+R6mY8iwUOz1ZRCgXFH9cVlNe5JbXTWXLi96eVSUV3WA5DNfGjuaEa3CCN0VkN
xyrqyiZnuu0NiqvfTEsg8Ww2jfp0TyzUWcLCB1VImTRkhkOc167XEL0OozlbE7/f
FVGp37LHaAFQYSiPtwSN8HznqMux3MdBEkui2zk0VkUxhesp8AgaOoRnP+3/gVnt
WYBZPeZlHMoSDETjNqHUqj5d6cx1YiJNfnZQw3w15dQ3ghGwdGeSC/tINOSTQ1u6
0nF0JtjLR4Y8zg45EU1Qs4eDqHdecMu8Qt70LcYOy5+1mkzUv0H9JOGja2U0BzqH
TXnI3cxI/Io+zFVtGdJZ13Tsc6PqSU5EMs2T+fXMIzW6bo7ikAhVGtj072qh8CzI
oHU4jB3xeDoukBCinb8RHECfb5dC+CxfV+zcLz4vLJRFMlh3r88C+ClpJ0MWYamR
+m9w3bbcWMCqdNX0yowIzO129yMlAftNFZAaMXB2yyODHhvCJ/J8vH87qai+HIpT
0NLzs4j8WWEAjxFLD02MerYe+kKOtMCt+Ykk1OuHYy29esAYGCMSuhMK4hcmzVar
VJqw3jxzHrSCedRiNHP7j8Dxg0Zh+7U6EbRgR+oMuvw0i2vm4e4Jb+zGpb7s8fRA
HMS2a/cOf43HAvDTFiURZSHxOc/uOxcwOL+NsYgXh8Ft6E29IKQP8cJ9jmSv6T0k
iQE8XePv3c56KbO9ddUyJlndmirwsCD2LHqspD1MAL8ELunyjJt5a+FNaopLki43
tNkcGcrIGE4qkF42ezn5SoqqQqhkzl11aikzBTlcZJbmWrOAu4FUitP0C2s4bz8b
EIh/MEzx5FNo7ZsxFzem1+rU13caCfZGKR8B5CpgnlkFINKORJjurd7XwpwIkLzg
jEa8kw5ILJ1H2nO90JNuxuYvaCwo0omF6g+sgSfSgGP4+WXahbRjTYlb9q+vzXy8
oqBIZBO3jKwg+jdnn6p0bHESxbjJ6s+IPhs6SUxTOPfzm1ay+7G2+/EXYTf67OQ/
/ft3q83Z2TZVoN+uumNtPfLgLyI1z2v7cJ6bB2Xp9jP/X5fGgzX27N7h7/vDtcW3
Vpe2ll8tobo73LkgVgIvIJEgD2uqVU2UQu/7Ytw1d9ex9xUR+Y0PgjgDYhBz1bXZ
o9OkzScuUGGSGSn2rZcGMqKfT67k8Gm23ht+CyjFdc6sCvmNOz5hRmZj/g+R1EsG
L/c9X1b2nJDrqpMuKmgKKV2CqcdIJSezBb2BivDThCDto0sElpCfJDqgeafGjG7F
Px1Lp7dcDujdTRTGNMMih4rYbUy53DWTtc2+8JVnGIhitYK40W9L2VLtJ0yCg5FN
ll9mG5MnArTLYoGRHfd7RpTcLPvzOZaCwtoejZsCPd9M87c3EMJfmbYCbBvQVz3O
j2Y3i/K6tjHIkwgb+MaW/W3aHb2jfF4+9wZZSLpABYliZgzjssU8L+bxdXrJJdG4
lOCXYaSn4DuetR8HX4pdHjXK5IC+Ok7ts99PGuKtxYE78B16QpZK20wV9eNsuxi7
3P6koGCCgxvB4kPMWXuVYEFEWbtLBAOntp8h7rlslMz1xYwG6qukVnrQi6R81wZA
DWx5xdn3gH2hjqDIhcEZwSS4HHpCXwcpE9XV1gft7hb3aZGl3tcuLLXKP4+EtzIL
WYaR3wTPbYgu8x+378S4m+qBDkeMFH1vR1qF20q1GJw9ZZVPsCul0uyYN6VLOzac
e/N88QcdUuOr9EvSTGTb1AmEGUSgV3KVHahA5vyyS5Maj/o/rc9KarnfutkluJXc
7CKYT7wOQv6P21hFCLzdWVhmJob0OvPNbEo8FeDByhinJZQ2MwrrluhmDwOVQyh4
mE7IbMQBgOKO34Jd5s8G4pP7HNcws0X72+PUXMxQDBrJXO8aTKX2bTP33vLhiysB
6z+71/0w+ZXLwV4uIQHrP04buE8FICgZxkHkQ3ZTUodPo7qj/FlDDwJ5gP5fNzLN
XiX8JrqopB1gMoHY5MzvsWPw0VuycGEc8IBAvEW0wSfTb65T9Ab9uWW4F5Tx9kLZ
klwIZDSjgQn/oNqEscqz8uE3w5oFMbfy19dgmN942BgGFZmjXjta2W0SW1Udvo3v
foH/iygcGh75j4TKL1B7CkW6jTomDY3oLcW20cbMVA8QD2gl+xKhjLx3nSb5zNwy
+6N0AWRTox1UjnfghIcdLMcy59lJznGNmE25NCSFoNWos+i4hZQFIT6ltw/p6FIg
lFmTTspvEYk/5MDA0n7UK/J4vw9nPl/09yPfuGzk9PhMUOwsaR4G2OIg9vDXceZw
29Mwsa7Tb0fs+7v+oc+QoBbApijMWGeGbbE7jpheztvvxedoGljPQuK05d/CEBJF
25wmcp/QB7tT93T58TCDuLeagIoKgtcNHtkyw9qXEZ7wl6DgmELFpNe12+VqXgaO
MWcXdE3wxYh0bS/akb5KRLG+57KjxZnd4hWMcd9xX7JyJVz/MkAdgS6cKaWjop11
ZEs6g4bEb8+ouSoUg7Ha5at2Vc3r0fVW3tVt8tFCqpgh2+X3ecQAX+I7Z6uJorUv
Ut8W2qJzqUapvyK1t9m5+RHddMeJS9XE16CjcbqVq9uTbJh0sVxbZFdrvH4E4WLX
DXTeyd4xO0yTiFauvCyHKhyH018FUqc+oWABlIzuZtYuv82QGsBSHFtAR9GPUbae
rJB9ik5gpqeEB5WIeaAOtswDfMdTXkICu0IzjrWZhdUn4im8OVQV4OJ9xEfjTODK
yWPlDLz0IKqhpUVF0q3SrsDtvcusJ2OuqsGlNuWeUUUdRMVqKwl2AsMIo2Zop3yG
PwuHMGbB2YzFJ0XBGmoIGRm5hhFzNPKxbU1g6esOVe6BZEEVax0HE2Q5ddZbXEIs
rneq3cZHBcYd0IY7CxXzBzjWsm83QiDI88Ep2Q6EDQYAa9Mc6WSr4ZcG0TBX3ke+
d1y3FO1KHZjYbOQkVSEXnbbpgMWqV/h9e9GOlEAEuwj1+QSflC1YwvX48yyOq1HU
rFlrmj7eANawdgIOkGHSL8eriDvJW+ohCa2UzARQDzXEuAM38+tY6MeAogek78aa
Y6BPfAJ1zrdvdCZSV6HEuHIu2w15k80XtI/lQIGQxH90N8mzB2vuX66iMp3mp1rI
X3KlxCoJUjbyYDICyytfZtlY+SV0lRe6H3qwgUwMA6iiyhVynr9XlelCcLJBME9p
4Fw4/0QI4x5A+W/IQDUGAbdUmKRVAu6zQ3EnhnY3bIsjiYWZUREy/7F3bjWp9I7J
H2caLB0W7R4RKZh4F+GE/KX6kTx9QP5q35fyrCThncrNJ0d2GjQF2EDbiQiKtl7z
Sfos1cmDmWe24fOPW60ymKk5B6CpC1DzMQxWjrO9XQobwqOyK9RMXqg5cynQsU2G
q3VEKwjpOetugBYZp49zIj8qeK0Xa2uXysIg99u0YWwcTfDyF/QMOGjCh16f0fPi
SFRb9Z7z/0igv0OHwfEOmOfZD4wIFUatLhCJiP0h7ReKatAVP0nubDkZWYj8VgqW
+abXoro5WYhhIfFDyfCoi90xno5GJPXA9NymdrBOnRaFNGBcwdnYM/qtF0IDI9F5
DJOD+1c8/Iccy3g743scAWgRzK6KRHIKPse8N7nugmRJOpGY3jm24RAJXjnyjVwJ
nBlaqIQkN8T8VWVV93qE6qjYnAX6dJc/iuc5oKaKgudLlBGavpCJSX5GSnrvEjhw
tYZsrJPoTRpHlf5stdp4MisD0hD4Try0o6EC3ZqaNb75jQawCmzg1yCapRngdVq7
rEc1xKDU17gSZob3P5BMfYuvPB1wYuMZinH3uA+G00Wgqm7p7NCj+H8eENXRdJhf
u49+L3U5Ok1etiUol3ymtT9KsvKuejSDZmULh2/5sdfSHUvLY29SK4kx8WyTRgZi
0NNw6h9KwoulYXFxPxp4IiKRpheSuzvoHCZAmhgX9kxKvMt+SDIopDxz3on/g0mB
vtuIfAbWu9NcT533LQDMECOrOsHpzrfVxCG5XrwqoQSYOA4g1+6ywVqkGWBUWDB8
YEW1lHxmtItMbZGEnq5uj6pquhCDWm0VEKTyGKHjox0IzOFq60kUa0KyhCkkoZ4e
XbJ89xcpyDvESjaFYwAFTQ4TG1MvFh7AMI/Q+zsWofIU6V02RHBQQm8FYx/p/kh7
LXA3uvWOjzzTUmJCk3u9rpOzTBGP9jZXk+F7enzccK23XVenrR3RLXDXzMU9u+x7
vZULyT2jCqjOfMye4Y/0sJdAu+7tKGRsI+I/QPr7tsmAJg2FKnfukXgyXjWLUCt/
KW68FOIDuS27lV0O2KPa8log8c3hEbBDcp/KiB1CzBDOTDcIXD33Nq4CeRC1+tOG
MJr0CBb6FaTjrjBEdEJZE6GeEFvtfoyOmRaSwq9PhJSgdT9DhkOwNpGfiaKkeUJV
iXaCVLD8V2/F2ijPrjEOK9AYMLHFVRt0klH4umQJNU61PxfoziMrAbSFxqq9xoyl
MmdcLFEI+moVi/mcagGLai9d9oeOMRm6aqEYm8g02ebXt6Du/0gGr6X5EXVxp3WD
iGJ7reXq7dvz90ytiroyywPNQ3ODZONzdx9snmsoD+nKwVP4r1AsqATzBU/2074i
aoRAUVY/akPROy8hkKIH4KGze+J78cOxljTRYo8ZK3Typo6qGD7jmpB6yZxrVj5/
09SC1WI4Uz5h8m2mGdROBtKowk+92OBD8P4OSirdcyqC/W8yeJlshHErYBadj0Ko
klhu5GHnOCas/PlVDbNfP6oxpEJUK7DLVd8rvjJVSGgfBgoWDSgOoneX+2zgBjMv
d8lRnq8lk24sLuSUGf62X/5RDuX5yTcocyNaZzXQ+MfwkdrsZgLug/PLwqrTs84K
hyYHimKPIUlwUkeYLaO9ji7uMRRFPbvh56F+XLhQm4oY0ecyrHithIpr4GEO1Q7K
bdLI90xntSHzXGzlHX0dLWpHUO9t2IF33JaJji84kCJlUcSAGYjglU1BhpVJyPw0
ElSM+t/9sO5pfwDhUom0T3ZHoUsL4BILVjH6c/ZoQy4Hg38RZLOGL2LNuqgJ0m60
DPnrWqhCeIszIoIWAtHyRnaiZXE4wWdLotqiNzJ+a8wS6FlD1CYYrDu2u+z6G/Lj
GTe03M1NzHMHE1KaF+ZckvJmTFFeh4u+38xmCvCmGYpD8AdMMx1q3Lp/oQOerXmj
yYt57HrsNlauBHtdqxuiR+4tgERBJRJfyibs4lNkStWOAfM1KUC8k0bpdnWaGVb0
45QyOVbuF53zdm+BhJcm398ZGTFYgifNY9xkxhr2OdcfuEEb/tYP0CINXkKbvuY3
MjcjH204EGw8WB+qlVoY+qrolMPluSsWN+YzOPp+MENjTCOaNAynRGaUsxYyTzTs
HrTfUnFl3Wl+PYPLqPWrsyFn99CEVWo0bTPGUtbSA64SCEfQspKLcR9+rh5b7tQk
axYkrWM6IwYDKTXFt5+Li4A8uyqSHI/+WV6PmZiXIAvBHRkXT6Yu8YVumREZlkeF
wFSgfLM3psGJfGGoI0IfJN/jbtbIaIh30LoRksQlMEn0yV/HmMghGvaZAPyY5mkJ
lj/BYzgNaJjJgeEeLN4Kg3f2banhN32N28RhSpmE/nPisqnqbALRIFu14tIpsQ0q
HESX/ldwRG2BPvj8C+1eDDi75etab9GRc6BOztMTqpMLSW3kjl2TLPaXg36mfNNs
eRLzxE+w4q/C5M0zJ+rAuYGb3y0dOXtBv4C+8UElhIEdgBxpsCbtnfLZknEoHyTe
Y287OknsK5Pje8QhJfm0uJm1jXxZoYmt+3Kg6cFJVI4YFON4ZDrtu4X8WCgwxjUc
893xJLyR85jRS0tvP3EE5QHZHZ64mVsqP1MXF/XUGHBFRyFSEAgmWof/L6nQ2Ug5
BCKxVih0g2hhggvRPJrU0I323d6z9OwNmZdjWcpI16UQSDhhKOV2fGzaFDGnJkkb
uPuWyikykXUP4cyVcuYK/AKyXPiwPROnN4V9zEe3MX67zIT3AeZn3FqUbKaIbxAd
a1IPGlsYub8+HHW+kUkB6VRKY7qKIrjvxEQVA3T2i28Ut1nc8Vx3qUmKPM9UCyvb
aNCw4p/o0Sh2HvsIP1mclxs42F3sYSLNuBth9dtboAwil4/prJd40KnCgrBU2u5F
LVDTpC3wv+gn5Ik9oqJn3pVXQansEqPDUcRb97bfDXMA3gSfwyeGiLFjqVrTiTo4
PtNM/ZWM92IKhj78cw/oDDOKWmXc8iCiG6SPFrS8HouwyM91cHvFnvetXA7n/1AP
qKXEGZudDHoQXrYT50i/xCPGU2/A/gVUbtrCjwOmnd7x3wvfhGOV96rrTPFpwp4K
nb86GIHYw4XvwfyfEul9JeflD0EA1c4v6joJG0CcQMdsp9LFpcajhaq5dTDOJqlb
Gey+ZqyALmjaw/XWyKWm2yhvhsLnoZeS/v+Sdtnz+gvV83Wj2oMpvYOyk6fcz4uL
XtWWxmC9mDzf6LWg1aRhD5cd1gFs86m+6CRVx5AsmZHdtL1iAMepHVN9I6JY+J5z
GLj39UOuSrbCb4L/Un81Jn/197qIEyIty6fPz4XmrQIm/Vc2XPZGGubf90ed8YjH
v29dCclGqUx1NctFD8M+JfVx1WKo8I8e55dMmDEOdXdgDz7xOV5UgjjpJe20Hsbv
unLupKsP9z6js2ht0Z+hlgQ0uSPcJeOIQmZcVmgHzqwDeyVefiEaU6N+1T3iu5M1
rcTKthFsMx5gKdSJ4KfA8seGGmOK0NieKvqxgf3EoP2uaqNckOGZgCeUHNEL6rKq
BgCgWoBACbYC4g/TVvtBHnZbAVU7bC08KjL2/grAXWCD5/6yoscRNZe++byV/bzD
4rLL69htVCB4KGs5RuNT64gbrXWIlrhaFj0skUHQ6iEAoZ365iplU+xQLSs+WeIq
UQWAkt2j4wwYbmg+0ePxZ90NvCDOecPKZC/ouTKdyDMGxBtHuS/9+ssVo8tOnXwL
nZCdFA5Eu7d0OCMWEOFJfHpZTV42YtFQg7YEMYDTEzFfZt/4RxjQ+yPtQes51j6H
Va5HdZabAFWaIf4zYF1TdD6/ftsFu4jFSO51j0ZqKgHBHC33nrvOOU6BAswn3myg
uL69YiCLVGY0L+gQETKngjpSowzEwwR+0Z69Tt02CR6VUWM9/H2CCJxlpOkr5MB3
CykkIFjmiY8WaUuihrLaSu+INya7gPCkcw+e+/xjrm8HM+52fZwddcEQQtnWeyLI
QY/MEgYB1FUU7DUa1fOcSqDR2O677utlun5JIBiOR7XHglLye6gWaU3AOEF6muFy
QuL0ZfPxXTnaFTpGCKzxSmY80BlNctk5xiLmi/G/dLtuNKH7bGdnFc2ghyufkRsk
/8660TgjaPiIGsXYhTOemYustBAS8mLzBwAeQsYiIZtBTeeCSVT1h+/yuRNRs/VQ
f5LF2OSAHKkV81UnzBVS/TVZv3qSLsDfHKnQergz2BUzcAsNJCwXuFvab5iZQUrD
qyXYV4IOISgPubDQRAALVYG5XLINebj7mLc/lHuFw2+FmhNifX2WHlF3FAmobynx
IA0lw0/Abu1O0+oRGMsSVUZ06rlzxAAArjnN4SxXU5HaINGnl2UNaZtIC4rSgxVG
SJZReKjaBNbcy7GumY47Jxi7d+IAHZzYxsnLy/QXQi1UJVAS3bGFc/txb6IkF/16
h5iyeFGkVI64n6enbwxROVyHMSGTt+ihOvRmoLy80N3I8sNqzSNIIMPtmqrEIT0X
Yj/OauAgSZoRDwAV3C9f4snWXqBhmOpHEdlTIAQcisPE2rzDfwBjlAnXE/78Seq1
ZoA7R4PcfvPbHRPmJZtYOvG6K/dRPZyZ202TVyLLzACpI0iUdJ8lFmvOBK7D81bR
vYiGjr5XvaoKS3GbeCSiSbsUb45RZ6Jw2Smua/+lBETTXQ02+lhFUGIAGY2Fze3V
cN8UvkD95NbGGO2nct/dCDnGR+aT6X8ndGr+50jVV6ix8hpv2pS3fImnN4kCAVoi
p+QZM2RdUCS7LBAwHaC1YIb1vX4J/HGwe3NmhxuiEsWvjl5lU3+ecqFu5BsKyybm
5veFb31BH+kog4Mn70eFNp8MELhOWsNvIrMpcfdReG+rDxeE2X91eO4fnYPYDLox
HpLa8lOJbf+rLDs62sVACe0HBd1EZsKwtzh7PF6DGjJeklW+YAIn9jJww5KG+XmP
sEiybh/fTCNWKC7ByDSp0BToW+zOEAx6ZIufDv8/JHK1wA7JMnax1R+k8++k2wH+
hqMLEYTYLZITXx+IY4urJ2E5NFjWLaUGDuWwxj2FQU6qcO/x+gfTdybkTP6/Y44U
rICdzmou/SwaWh2Pirk9sdX6I9zF//mqZajPIMLLAPIjxtwm+Ih66zePNQPqG5oG
2rtFq+Kjlm31VByXeFzr4s5APSBrlaZxw5D/8PE+E3VWqL0vjlYKBTn/C82b/CJd
J+Ms5O840gZxJxtXQxzLmsPwFx/W9L8Ro9kez3PG6+hSURgdK5zk5WTLSrD9H5Fs
bBWfueyXnvvfIb+lpIEjCBvWVLnEKphJ/f8YtCUYNXAmNn0TBTGROr8ukDz9h8e8
0pEUGIZctqEPC4/G1BmIvGhfBO5s7yL1FT+R2GnnNhjRRa5mSLxlqQguNr3ywsAv
3jtlMFk2AbFO7BCF5HV6NsMp4ajYSz0VcU1PYTqr7DKJ/KOdxQ42YjMbR+B+DYla
i6WaOwLo2hd0LGjd2wJli8GQcTKy/C93RiyrmUIgVGLJLY3pWYpzV6yFdSfKV3ut
d83FiP+AhDx0X8Xz5c6dH+k+aDOVgaIMFfKtnvY4E9UKx9kIUvvx3YOARaHZvNxf
yW3+JMfXu9vXZsW9yu3zXlxe7aJcJlskbnp2kll0ZewFFi/iGf14EQByhLHmiSeo
lYVUo8qvQSiEOOd9d/Z/zdJIvdMFCtPvxH9UkYX/JoP4eTbKzF9qkV6+tPi1iMOR
FOH8NTuIFwXXVqn5QvQ0DyQAH8FYWUKfBaxW7M9k322hqEiRPJ/5SEwtKMgvAEEb
TrDwLHZVj4wrV61a/YgDdFMWBq+0fFH7VWE94WRLFthG96oPQ/Bz1Vo9RfrT2IGT
2ykv4mZxn47j+DD+LlisP831xg0GMeGpeL6pYtnzUQvbY654vQ7s8s4gBTKjHTDz
gNplKyHdC9FmLMK4ySz4H5klPqvWgB4c0fE7fHaknJY1Wuj7RNQUYZ45rBadbpDv
DbSp7REtPh2Ygj2EskgmJnG+jtxC+/WKwoTe8SEH/A+Guyrxywl4KwRxu60stmtW
p0/91AdtGanF1OFZtMQJ9S2jwi9LvYdLHBKyhSBWE9i/MfeXT01lACeei2olC8Vu
OmQvbZU+dty4Mf63cYGOT1f4TuP890YXSAzX9ZgRgXF3KOSv2VGFtoTaXAOb75gt
qPTtXFfYwHzqdVFvJ05ecW9HzAgeguzeU7DhWvdMLSg8yDCHTD1EXP8x4YL+UklK
31hxPYyFzeyhL1Crr/cCs1JG8xk1ClUFHKe6XVF7LLnE398DolvWbV6au5GAihN9
LfROefJk1V6d2GPxCcKjNyM+wNCz8hpdFNcJywgzw8w+ftbFnU510fxKmEPr4AIJ
7dI7IMlSION22b4myfPbFmRaWOvFUbBANovECtH5ULEvDzJkrdtBqlpZijX1elmG
z2fkhABTgZ7E7aI75wVH6HtpdPCDAYs8Sd4om0RFlbtOM2AN7lAVa9c6MjYMr59V
Ed2584tdrj0F+kkyK6bSvBD4ngc0HC4bcbP6BgQI3+q417FbBXmjdJW9WdrEPHCW
geQfVsl4SpT4fYwnBo3/ZnvSxldhfV80sDmSSaOrf9SGEZE1u+MC2MiLE2n/gSKq
laVXEbBPcDBeR9KROAtwIjiIEf9ujVrT7Wcnk+hHp96OpL9IwwFims3YUeX4YD4C
wTTxO+NHLSDRlspO4PVKvieEP9/FWEb78TBO5dg98AGm2NveZO/qY5a8EHDmdqMj
8LgIV+gF6cihdS1M55bNP5yEmumD639HqWJPCAzX2OjrN5PijHC1M/AAVHqqXbg3
Aa/fQpXVP7F9tuiFugXvN5zb6U0QxDNaBSiIBiNmKdaluw1MZqgGuKMsNaZJFQ+T
JK5AFy49v21/wla61UaRycq0OWH+laL0hX1Dc3S6D7eJaBAYK74sStAisYdnCyff
FOegxg0KTK9WS4x4jWdO8hiPjbFeul6dYamBbvjcl7PvUWw0Qmuggea4yo9Jv+z0
a2oHN9lMCYspx5Ln53mXGi+RXxBz3ca4FhDT25MxhKjvxAkuNPC2u7cLgvqLXLgs
SXzloSVy67EHCWdgoZDtzeaelxfDv1uYg3qfhA+/kWT4w9xu49JsXQvkCR1gDNTv
BuylozNc6QGB77iY8yuevUwN2KRYYyEIjCO4XZlpc40JlVv/+NFfL5/ab/Eb+sWU
JqDWhVLCCqqxn91gtoFiT2m5pLnyyqV5rKAACjdh/bGEhtZ6hwkHCsVd/XjK4a5e
WVNWTJaF3SY+5fFiGEtAgD2TlI9JaXz1mn9HLHFbkxgdPzeP789AL+EZ59VXassL
uxH2JxnT8/kFLfMn9pxj6616igVZxeW2IgexNa8zKTDh+R28MbfhOTMqflp8/HzG
/O8xHoJjNYksCB5YNPP++XFeitxAGS2VqXXZGBpprdtj1sHm+irz7+2a6WF4DDdn
njVpKQDigrtt48ORu0UrNMF7Ieo59g0jzMq/3flvc6pC/XQey3lNZAcNfixzpami
PcyhQdyI5d6LBx+PSCyfaKsfByvP21RVuGNv6g6XmxTAZ0defwfDURBV7G4Orn03
sVlZdt8g48n+cabr40D9mIXOAMIVkmccXxippZRSFs1BhhAYGv/2ESZcIxrxRX76
1TmgOdEnuEKl/ky8FXTY9ZsfFcLs1D4eGpPDEL746dgzNyzFiF4iJHDByd6H/E5h
cmjFScHHHH0Q8PAHx0GEKZpTGs7F7xKhSk2ENr1zksZSx5XU+5MVtAgyrdueqfua
dHs6eSR/un8KOrQz7QZp7JVR1/C6jik12iilFMYRFSzPP9yfs5FHOXxhAqFjxe/m
XYLleuAUnfqthoTurfrfpjvk8AmnvERh1SIqLJWcAmeH1N7H9XDb4e26sbb+9NXl
J7knGXLhFgmeJXh0+cq0jhid5CEYpXusQVOHDTidIp7nasq72rv2GloQxY2p5kjb
pfH0iFW0pgKPXAJG8hq+Ezf/HhSzPZVlyEv9USd5dGsGt7ykJF4Mm3+lVLBpWnjB
IbVQQ3rP1nWCDJLPYuenTGUo45651CL3Y9gAopz0A7G/LLRwsP4yh31MNsSTyCRd
D7hRyitKSx7GN/iOOBZVjX2OkfF1uHGTCjmfKb3zfCwjRjiquRei1RZj1VDZYE84
1XU1skKQMmz4no7eEAteepuE1aG4DQ6iop8jaL8YyDmGWz4F79PFJXk8NV9mjQNO
BqRzQBLNlh5wHM9hoHhH17uvBi/ixitrSqX2e7JrjAI+39CLXnUOMEp3FJMAJi0x
fS9BO66p1MT3yV5t00bKg+ny93tSu5H5+HG6GEXrVwbGjvv+tVb4w9mBcUvAVe9N
4thJz9KI4c0ufKql5V6V24a+YTgWn2+DJTtBZuWe5ohBPhXOtjVAobqPwIVOAASd
gMlk6KgbhH3R1LeJJOSTymRThL3t2IEXsrZp2/TBjulcwYK0X6mxe6tYAaKiofkG
UDuoYXZiAIaTHTxGoRWh8ojywTFgmR3a6X+rO85/jqlydJQPLQF8/afhdgahUMaW
EwVVhat/MG2zK6cokM9S7pHjmxm89BPZrDreJegHsNVSh7D5/znUyn0jG/nH5p9Y
WeKs0NsVke/59GlOI0HEVgKQU/eR5QC8RfhvjG/S7kkB6QDZKsq0lim9E0XIiu8e
8xL39V3zX7PrsBJF2Pg4k+hYBB2nNMrWhg6TsSRxuxvwakIN+GiCFPg1e5tWbtCW
eMomM7uZlWOOGQBamwHHedqNEuyPfEgIpEcf3QcbWyP8E7p2p/I4qhJGyFcHOydM
UZe3QujhgnHbzteiFLt4tOhh+u8+Tj0cY7QMfuJWdlIl0QcvGwFm3k3bQcsq1MQ/
6UfILannVxXt+9QYn2xJGU9089f93IixVnQRMYlqnFygbnN9OMGTwCnmvbQSFpgp
k4igdVd78k8GhKZtWAdmESDCYDByTVaf6V8hcFiXR3jBh/2CbRdNYCLbNDG510W0
YXLvPTVq+bGMP2RNF8v21Z2xsoKS0GHlm1szT0XC8V3Bspj/vJ9aPln4vh2DdH4E
Cr+c5JD/1xYdFVL+zxbbJVzi36YY2sUp5RG4VNRcqk+k9nG9dK6JQOxjV/wlw0XV
2d2F2FL96tFyl+mzbP3mUV9tr+DFgtJmgKm6WJhaFVUZx+zBzswX2L7LyKOY3uo6
N1aWJfYyMswMG53iIk/ULlUy+9c+cKQRSPWnlZrpBdR/FSz3n2IEsC7XnJaFKngX
Y6Pu3AhXCHm+fnmYfosSNlMBHXtXtN1x290WoDcbuMRZGuu5W+QgqST2SGyni5Ff
qQiNaQtu2mSaQfkfjvkNNMNk8Ft/XTuqm9T0oi2tWQJ7/69oTWrJwLo5pNatUr4M
annufMmrLTdTOCPgoCEZiAStQKb1knSEtNZKzz6OsOKuVwg05aNOFWQRXZh+JseR
/p3NXL6ZvpCddCZePfwsLw499pnY2NgPn7zijyY0fHvhCqw7eVYf96vR8TGgSo5Y
GuvKrDETCIG3+G2lVm8fUyYkKtU/A8vMW7MOt1a6hPqDrilrMHvZFceMTCKRaINW
sOt1LrWQVLgQm2fa/4z7sfdA1KMXDv0qsZs47hykUQMpJSRsRt9NulwXbj+t6bwX
xpVLB7zfHI3LhlvoFdHvMc1KOG2rd+xe2/e3aP7+jw2CzVQppCL5qgmkwZBxoxEX
PbW4D08/VZO/XGdcgn6/CScXrPuHyd64Wl4S+do+CFEpX5aeU9U6t911/hO1nQkS
+Kzr8SuB2xbBR/8enQNJjXtUHzP0eAlxyM3WDwFf1V0H9UvPAjkWZgr1U5fceV6l
GoCsIHv52ddrTL5i0zQVxWAQNTfdPVq3kq9k4FHpS10qe9BD/hwMS5v558UctIee
o1Xg1wDZdk/kstwW3+P8i4yBfJLEs3iK6iR332q6woli3RB1KFb1CCBDjrGBZisc
Cx4M0TTa0UC7mqTun3dBoNMIcN5pH/jDCdFVwV94l+Yn0QxtlI1eIhWoat0r3Is9
vJkDqDdTA0E1ef2T7qIAgc+1b1OQ0bqTCiCPBgMvXw80RHhjgDjSeK6ox9wZXHlv
hnfQ259ujhRkDK+CYkM5w6+SM7eGIaONAJY6dIstfp7w2q37BbXG3RYCi+ADe7tf
2Ff2kfJrZs49DTLhFbiyGv+wV6zCwN6R7ubbH/lh5sza0Z2aeJ3jlIkJAXaXVgnG
kedBRpfFTcy6jYNT6Wv9DXmyK8CCaaAd/ZbTIBG2NCMzG+mH3MtMKwvOniLZiJkq
MdNnkQTLVr8XCgPo1LAhPEf88i7BqtfIed9sZUz40YohCXi1Tzs1cc/KXgDwHCnx
y3xv7iLUKIHTwmxtOlt2Jcpi0XnIP6QSzUOUA2ybOLp0Yqql72CB6C9h3h+RmX0K
HB/ugku8+nrDOowXNblcCAtuVyGRzTOIJD2ieTyQk+kfAg+hWNlKRdrRJ5Lgxb88
pRxcm7ceNLiijVc8Ulw/SQ9iADx/d6Idxc/57hldP9bYK7slpuVftEOg98z0Uv4H
HBZyHv71ZiU+gZO/EwIxggSJTxVSrpztBnRwCBBni+Do9l6sP2G1KBx9yDYM3geP
nEJqHWig8JdRyJKq2eG6aRqr3fqUNmEJ10YWv+FzrIEUN3y0DbTYc+RYF3KHqsIe
jPUADCARvGSA8qOZyqmUB+bQZ2hRMyJznXfd/7i9owxDR9jwGSJ6x5NaO2ggBKxQ
npv1DBjh43JgqOh48yoC+bkSI/cqvJy5NpGLs8H2x8JgponQCf2ygQYX9VuKkAoN
WKorRSkdC+BwJaUng2xRxRDbvRmDa6FgBG5/8XEaOpGT3jbQH4hbSjOhqXGCxfTT
W0T9LUb7j1JM4QrsWPw2vHpWgDsZnOEdfsrWTjTQs9/O2pgLMkJFDHXHn0tKoUaY
oNoLL+9uqeJr3jGikhT285I4Z+BHiADT2/6C+BrhOhXwLkjj1B2h66hX2MV1dVR4
7wN6gsm/AfKZYKni0k/IfYki6eNfIXzSM8fHaS3CGiSVPjIYpkMxy6eImxiWgE11
xhFOsXo77dAAVOIj1PD9sI1c6ZHvcoeodaef0Qdt3aSp1Mcr9+6Op76qzv6Dr8Hm
ZpROrgn1LWozazcsynjuu4fpBrKhgkLlQcX2NZrwwXAu+uew1hS4S/bIksGaPFHS
UUkzogc8FOuST5PI/nhwx8Lzqjt/MeD1E40s/Ymg3MtQuwQLKxJHnkLcaB4a/xHo
e00vk8ERIB7sqwjDp62ZJTX+8FEfkOjTfUSc+BCv7XuqW7X7cHkCjyyB67N1C8Jl
v7D1n9JSS4IJ4E5xuLe7PQSFto4fd9PwIYVRB1hfWXIiv7d84fIwPDCIxn64rV49
mYjecr2W7t+f+1zueGI9mwfj3akpTLFsaV9Cm2uTjTMkpatSy6kNf9HpSYZo2w5T
UzhP30hJVkEbmBP5/nyqzvMWCrMH6crH7GdkxaaQQdIZUNz3yNVU/daVFbBnbUP2
uVi0fbl7vl7dcmAmYFbgZmonn8+M79wfq+rZZBhUngwI6qPKc+GM3aAZZQ084NoS
vt7kv0SH7F+OqH/sop94ZxZUkuYa8q8Ji6KBurPlvQXByyoKPWkycF0268OJWSXK
kY2t2UT3cvMu7ZX4q3PoDlSSnzYoCfsa5Fwet5P6/OAunSv7qm4rcwfevuRVI70n
oR3tBjYjtdQbRSEBkZuDnyhpLRpiZGySA3QIV9Yy05wTuJcEqriZ5JOa73dpHJNb
Ntsy7B9DR8BxESyap7BUeFq34eBTLkjyFUxBB6kf5NrkkUrctED3TYkYHjfQwLpm
1YG/sGqtg0SDaA+ZuQYNj3zm1q2GV83H9FMd+niDotArAC4w7uizdxJdY2Kwc0Zh
841VKb9PeDO3Hib37vpOlVKwrqPHlLzSmDPG8fc+hFLp/WfZ/8lEURLzzjiX35Ie
1N/32qLOtki4T6iNAPCEI1N5GrETrlYKQsOKJzG6hBFKSyBXvRfB1HDz2XaNx4fK
x3HHqmSmvf9STsGeASjbxa5tHmrsesLQcQBNzmELnuWqzR2muhTDvBT8NcwcWfEw
QZO/VD2mVK1N+hAarzmBw1RpeyX5tYF1gcIKTaRUHDIWSEYGNkQ294iZm7JLU/CD
zEfwxVhOvKC7qfM5YpbGlM4kQMe8At3gFfarufQj1luV2SxLHtI4Hsbhtcn/Oyoc
V62m2VIcnMB6cvcTYPQ2pKkr9H3o6Q51dpPlUvyPB4BcZGse3fKNaE5qB+jMb0Fo
no0oAKQSo+sGe+22/5kM4oHLxPz5mslmpvBfckdsb3uNuc4RXXF95yb72oz+72Af
LSkdYKW4wWYvlCMwj7L7vG9Q2KSErfn2MPWrINwYWoB/7eNZf2KHkRCKdCco83AD
mnvX4u2sCeMWIfjd7Pqlisr+vap3szT190DcXXycCEdQATxCzaz/Z5imxVCQSOqU
wd9tP14KULttNa3+en3BCoXcy10xL57YsPoiwh+6I6CVxkBkHcqzacSdCG8bL8Jk
oGAs7q7pAfjMVHWwgC520RKuJMiOs9ApYxwH1vTTCg+My+8tUTW2GNOq452TkcrP
hD+6eBu5g9e4yKydWlKqSFG7lL8XXhBovHAzW5Tz5w4LxgRD3DPxoPidW9lUYOpc
SWTIq8hXcKG1sOkAkqnVJSoPbz0gAc5MJZDrxxms6fGhbnJIZHtqZnay6VCk58aq
ZJldEcfHUJpst9WPbw+p7giaRbwcyzKzSoH77a7cV3kZRo9k4UD03RLx6hfyHu3D
rOu8lpIwZHyO/1tgfi6Bk/C0tF6mrIdRoBx1gHNyCi8Wy32AztTBUjhlbYB8frMY
fw1cBkqpxEsAhEOgv8EsAfCpzmFG0+rDLAVMB1y6aNZUBrxZAEnAMcHOoY2ecVfK
2S8Kshy7thgWIw4zuCQdte6BZ47aXv1ZClbai8nXOpMItA4aAknyUrs3NF7PFiZo
b6WTLmEKB9H/8lcTARn8xTwLHVKTlM7STO28HEVGxBDG7ZNhktPh5/pEth+zd/Uy
UGgbHCLuq9rQ6qwrLnEhN+bhPmwulHYMZj73wPHL7vdNHVU9sOtWpW7EUWm2fLLG
UAb5Nv+PrX0bFzhj/rVOE5/1Puo3t3YoMAGCVelvGh7ysarL9E6tgjj2Y8xi4l3M
KHSkf+6OmmeW2JAAo3TX5uyrQY+68k1dVm5SlmGfP4KkpXg7O0ZAq5lxoqJlpF0a
DFTN6y+4l2NPJyQ0tZsc2DqNJhVV4qnfHcj2M6o3y8GH2IsFRObW8WnSRGF7J9UY
Urfkq4whZtmuQDZBmh+6n2UI93CtSx4ojSav4m+4SWL8a9FUFtZufou09+VhXVQI
+1PE3YXgLQHRC8e/PtlJVSv3c+vx03qWP6zZ0y+bX9eglGTuHvTHhafFuFQ9Idk6
4+PtJ7M16ObXO4+LWyQPL7jLnSimRGhWljcvUXKjjARA1HthhMyQjGSt61dBgpuC
GP7o6kh/PYmSSdH7Rp2KaZd8fEjoSjKgtzbKa7zOFh57oc0dcPCOJOU2LDlKaFml
b35cGWkAC8sdInmRW5bFxWUFcM/tGwCqZ5KgDoTxcxBslukHlQOfoorSQECwPHGW
vokg+M/mM+oPCxsazW4I9pZBaUo5kPSLDlHgb2LSABGZqB6LrUVVWCvyTlQfNpO+
cn14VcAljCkgPv4E15ofDnkXd2/N853Jrp98j5Dx5X3QkSSpK4bgugQ+s+Yz/ojQ
uh9Ls/pqZQfbgh7Ox5ujU5uyfz4+dhE3mPaMmjr1SAs/KTjUsnpfwZLHZFfIFuwn
rjbMY/YBFUG7FbJI2nZPyJgSH3NJFWNTjPwcobB+N7AWMpIQrrwfW73wFtGSu2Ij
hOWjdxOgK742aogrErtRlq65k4D03Ac0gnfq+3o5P13sRGh/YrWW/KkNAf1QyCLS
tDczirr4V8+m+lOJBU5SSw79FUTdxoT9F28OfF8o88Wb2H1F9ojl57IeYbMA+4EF
G6FpE2D3QvAbnro0dSgXGaZWUWCSrEAB2qjdFoyePyVCXl8OyccE7GO+OFudyKCc
EHTsJEy3BgEXw61JRRZoMmn47P0PYbSTjD0oq6HDb34LVQKYx1oxn9PgsHD2UW2+
CfnhNAaSCgenxTOSMmlTO1OqnLQQwq4B+0UR0ubI6uZGLcKAfP2m0JyY5x63zdzC
N1IIa+w/swFOykMWwV1ZgAM3ZiZAvhbpHpjl7sC+StODl4THyy3LxoXjTMa4BqOD
hpYlrDXZchu1pmmbz0oxBIESDcQEEOtRLubfEn0fp1OEueek+m+MHtP9+rd2d8Rp
g5b4iyavvcyHpo8cRiB7xUXnSy92KspWG+7tay3kEJ0MFX8RRP7RZIgtVKKs4+oO
k4wVJNNjlVG/NLp4rPm60o6tng4QiuP857ir+0URNRfVilhKCCUAf8clRYS+Swap
CHR5ol9D5vaOtUWBdawJDtHJt3w2P6W9rBnW0mBVxp1Zimn4VsxNbAXwmfLpQzLx
oQHQZVg0rjtC/iBGEvVhjLwmJQ37kI8B+9MpJiD5ZrbTCg0UhTnOYXbXWzXrd2QE
BQULW86eEzU4fZOjTda3+oWv+CAcdX4vdHMYEoaTJVscYZSHTmqwfeKI6TnIcY2Q
Uw0Z2VFPZPVjDImIsurFRqxUY1/Ft2MEicLPmH9Y7M3AtQf1CjjHOLPXX4+4uwWg
MV/bKPZ6KgZydeo5nov4O8wvF8GLLeUL5yhOIvzr+sslksLTgglrlgSK0cZna515
0tFQaLTmWxLCnrYT7i64TRnN7CJGBoggOd2ZGm5aTO04GtS/rRktl347rgY5xk+w
vomheQS6R1XmxnADcoDEr76evDfraJdDIq15jL5YCAFdQWFEz8XejWwNgRkvTJK6
NSHuGm5NPTcIntdctwj5rGx0JWcIHxJw0U6tJXRoG+umMCwgxtm+l4X8RKUk+Srn
DcnH0XhpQZuCPZIlpEOrfwdAub3Xr9sBd+Nw5wWAtJ1TtW+K+GGLk31bfaAiMXKC
fR1nhxFfZNPAfmRJdjwHd653pKJPs713fFDgZKPT8ZDei/AG/dzzNa3fI3Bc/LTn
AJPI59ca2EqsQO3RFH3Ko8OX2CHoR96bpCACx1x3eY0RGCnd77loPuCjfECdjmFQ
HGaHprk9uWjPIYYEALRUDy5IMUyYAEtz935Y9TNFVb7bV+RGKVeVAvr7BpbMRorI
hR8cqCvn8k7Y3Q/r5k/iL4+FikNRgRmy37Yxeiv96Aj4AcUdk4GsgJlASZCr99Ik
uGoslXKEe90NqFcJTWOkPGinOaxyBU6hK/36xHP5DHvNZpwlrIFGFB2CnGs7nE7y
ThGUsDrFtZjAYzYsYcIRkAGtKOB8FmofLK5xD4aj2nFfxawsRdxxUkrbYiSOo3Bj
urATCkBMcNeBk+7CORYXro+DtSdVj1P9uYWh4AbWyKqiYgHWI/JWl0iIrQuGb1Ut
tDeG3FUWlGf8/C+1HS4Pz4ek6iW+v+BmwlkDLpWttJfPiIi0CgxHq3ULnfGNdZn4
M0jmrXqSR5QdEtyK2q4caeS6Hk9r0EoGhQpTA/Gm9NjCPXTfVuFWAIxu3UO6QpK6
sqyCoytX5pRK5KmUTOJkJ8FfuBbt7NY6RGCnsFNjKHA+eiTLfGowBMjEzox1YRbX
eRkXDSrbsQ6Vr6vJ0Cy9qeSi3c3BbqFTpFa56lX6nytzn6q1pvGfKmFGMmfF6jkw
1EURneXXdbV/M8LlVpsT1deUzeqXEGUUZcKJ0uXc5IVSiiObuaeSSJiCRr7XzHxm
Ycf+ihu1x9Srl0GdrDW8Ina+IhQiftdKEZEQxELg7+QeN072/wQeei0iNj+jh1uP
OAzsqnb6HupbvBNuTAp3nfvVS+0ArBmwGPENkD9Lu5/TARfUSyHfHn8fF2pVsdkt
RlCVprLk4mNsl16FFx+H2J2pY81oucqbnwxwPTCmLMgeJ6p7VEtekEinKqqycKit
ZjERZbHwVeoFy1glzZRUfuscXMujuHlvY9a94EvBrUb4OYYYCl7YB0joAnV1u7cw
fUV2kgWtKKHE+76WKid7yimASACN7ybEgYK0L2usHTTYC2EIw4wtsDnqLC5tl+yH
rb+dmxxUKe4ka5hVobaPDFgj26YwgDshZpZU0SgPyd4krrnQUpfWzbPVNeLm4Rmh
VzBgoQhXUbZK1wD0DaQzbHpb7Sk9RvTwXGqOo2SYAwrjVG72WZfteU+Yu05du5Qn
V5RjpmK+S9lCi5yGpcZbbKcfA0IISpJ7t/CQJ12eXZrmPtMOqGJbTF5Hr8Yx8Zj/
wJJYSnM+RSO6lIKay1b5l02hD8Q2A9tHBA8kzg1ceQ9kuNt5wIAHi1e8XwZ5GNBm
VAXgand6B/eenMXqjk1SFPG6PKteht2UQFqzila3RIXp9c5GDkPaNgfunGnDP1xx
o4KV6MCXoqn39AWJdbHVDn0PrFoUfCcyDltmgjxamdNZZwKpN5UCSk4ef0a9pG4y
SUoB+kEpfWfvTXma+j8PvL4Z16c89Qs+ZmF6OH0IWlIxZ0fI2H7TznGvlgzXBp0d
FlxN0DKyW3OISniHLHPQApZeqp5F/61UjH7sWRdOxvmnLXlXbEAzxNBlPscUGvRw
/cEKhJd36M6kOqV5pDEi/Mhe/S2vgB3q1N2jUG08SGnqeojqLt0GTNzqtwdhXVjy
gj3pZiWHOphm4McqXiGNunXDEgarts43v0btANiGax0MZ0krNbWRRjmiux04wcAP
3el7ZXCzG33CG3GxaVw+EEhlxJrQNYlUQlVqT9MnXh1RwBqZ+R+mzbXlJcZDt4cE
Vsr4l0G3AtXISsms0HiX7qACAhtbzkVLIPP8eUb2cgLdPDkrH82JKmK5prEp6Hmo
K3YY5gX4CMWdic5K4QRG/mKoX10gaORMylOxMTmEl6AQF6pAkCOew5/xUsoiTgXl
fnYc+EWbnJ85KjYAIoDVXhNHC2TOHmbhkcfWfOwSVMf8KMmgOXdQToy9J8q+mI5F
BsEdqvpKo3CuaHWp3FGPE4D3ZG3noeX2hTkWw0F+qnkrL4aEypAgI5mot6Y7gpVN
r2ETMKa4QNTxHTAHxamt69OtrIDKF2ivPyJ2gF1SJhOQ7Zdwc33HZSv8ceO/JbmJ
3ZUt2sw49Ov8g0ecjzWsnc/h1DH7E90+c5NbRmvbO01bXVQw9yAsFUGpYZ/Dlr+s
2wCQ/BxD5Zy5ZoZXosFZb3mZth+COvvCnwStHTKjavC+j15swABGK/jz1weiPJK6
9IrrZde0BCZLbWcJhTcL1IcU6gSsHNg6vMDopUwrcrEuPigNtJnS8r/lHglLaaHg
UIjgEdN++SFk/EMVfjK0GoRnbiqFuIxmWMxTLKHc5DwN+o/D9Ze1Yrg9it4HWTdw
lM3w2m8noxrBfV0QubdO4D7WwMziUv6CssBEgsm5eqZGeyGk3PNfCjQwZ2t9JfFB
sULig8JejMtbQJJdBD0bwBiB41d7DntM+pgAq3+Be7k0nkwuLMywAKZIBt5O6xdi
LNamRI94/jtu6SZLdwUwOVv1TZ6E5DakEZOhKO1CNOEKJoG3a4lJ0aEl9U08Thpf
1IjmZ6vtcbWgzKz5qHOAMp4oDtBkvouCCDZ3eH6bsu/Ij1RaPuPdtylNz3UsMmCV
ale2YToDeVWd/y8n+KIhhoWt5wsI+ZgTHMat+zaVn4vY40Pi98G7hNIBlKQr1+7O
Q+XvXWP0rNdr09FSKvS4xdne/Rli3p5DJB6ahTLWu3zD47Xzkv869moqHJsp7LXq
NyoYWKjLYQrXYZ1Vw3tqROxS0qm4LaFvB7sJEGlgPHTMnVjXVH45wqGwDLwgulu4
okn2qrrD/CjI6DxbKyLc32bWFMzQnRp1pw78TsMySJs3/tnAK/YUWQ1XokB8VT7L
1WpN2zT5H6MmqJWoCq1/sLbEI6mWz/Ywsai8zg879OZaxvJ84jrqeflEmWAEp8vE
stQMiNx1JtiPdEAIx4HcGHtVlOaglZp8de+GmotGILY7/zJylcik+JqcCB7NzPwb
A6aMCAuK0lQLTDsVM/01LZiKVmRVLQwKUR/EoculvxtzYvMYsWnWiw/7PzWp6h5K
0LyxH5QkrysUNUVPkI/64+A24JcHV7L3Y6UPtuU60sTVIatoY8He+dLIKCvJNY/Z
M2xzjRvcX07EJTXdWkxe2CryRaIIuaXuIeVrnoLmiQGSlvCKeALLOfqz7LFNnOP1
kFBQGQhQ4jz86eOa8iR+dXs119LAmNjdPSaPuXhZXTIqcNSLUE4XrSmdU6sb6c1k
enOh6A8jpFykFOtAbQH1QbGbkeYGOfhLw41h/B94vTA/tF7V1v9n0aKES1NAUcoL
ULHke67XGyId4mF+/T4X8teAErkgfUSr3cPLWO43phuV5D65/kixTTq/DHgjJSDm
tJplQ0cqiibrEDcl+1tiK6wfzjd2vBSA+zfiCxtG3xNIVR5KPUD+KIi6G7KcIij1
/nUGYKJIkTydmF/z2DtQWTYqjQsC7HGIXDmR2MF2V2RK9nwOGixz2AJShwAyGNtY
h7PJ/wHvWL1BemnxdarBc8nKcTJ6M0701qIqdqNN6UDpS6dqZ2d9XqMJ6VyZiwr6
IsNjeUFm/GTFmhf/39XCKVayvQAMuOOck0SwhQsgnqVgodb2YqssUXYHNk9aNmQQ
rYi0F7at9gCaDNevma/ccMKI4LNFypMGHZ30pyM2Wzl8RgPbpYKgS7IbqJT28yuU
uvmu0StGVgI9NrKY/rcLrRamw5eFzTOhQZ67ndRpyEDPU+q5Vva0/SUyDYb9mblE
mLYduX+U6rRgUngbibVjCKl658VfgImiH3kuUwvQY/maOFiX63dyybuJ60o8By2t
lH3ncMZmDRxSp64FUbQ04pWjsyMDY0U7+BV4y++CkxqtNDoYZGMWgRoz12f4nu6F
OtZuSFoDFtcqpOwBoFnknZJR73tJF5mIOVDy8Tz12VshHGuTzVLQ3MMQFylkOC3w
srdOM5tnmhaVFQiEM8rLbxiPaHHAi8VXEcT3MUT3ND2BfnKU7GDIFsPZnHNNrxqc
X6D3N3Z5qO1V5S6XVjf7VxRIYpUOZDSI3L2n4h1FUwSmEGvErX6dTWzB+SIkeZzs
KWf74XEgRmlPN445+Du4HMyjmYYHolVwStknu5vOwJj3gIfNdu+0lc0WZje5Ofb8
gIffYQ7SC/5C0xxUO+HuVqaaEf3oV1vbO60X5ivn4U+M0g0M0Cf5d2jPQI/ctpmm
hMWDCLHxWSptJ8Pb3gZkX+UKfXmmaN5ipqtwWWxKXRXig1JhxDwZWXPAaFYHHXIe
qYbd6WbvGzPdEEy0RTEA687uVjqdHAtR9UEPnpQrTJawxkl5moFr7J23MJRjneQl
6zIuBeA3RbbZJZHKXPztkHilkEf2l+GhuyJ94GjB03HzysmRV4sXWLaheAnyVLIX
kvQR7CioAZeYK0NfPbmQAhbon0WQm4is0p2aAEDQYg4ElAQmRMSvo8/f13R39a5v
qkyBtRd3pwU+43MFiF65Z67s1MkK+q32KKvlc3PZcGDlV3WcDKLHF4lkjNgrHezk
w2XP5UjpiUcQ/EUsaiGm08qLlb/ZRNQUVf4y31HliTKhInfq09g+URSHXpacf4mP
gR6Gr531m0qIEAB4tZHtym6J9rUUDVt6Tmoif4QmMeXoapzMTDmsTsJvXkUEMY6G
OlEMWrbluhS4lx+N7pz5UEpECtURiB7Wi9yuV7PvRftqH/8gTMwGmMIyRriLQbEm
6V+ovdiQzyD0FMvZZ5izuq8AuPvIsrI7f1cyjeJPqwqIHpoBmZu1zEJ18zkNAxZD
kcdeodgai6kPkdxrtCxFhTvwdRmotADhr2cp1uMSqqIxAQT/pPahWpzEDtkJoGdu
FmmVo3ASvRFfPMjO8vjgF7tEO7/78M5nepR0CsHqRlr75C9O8K2PQRadxevdrJYL
yxN6d/RKCkDkmsY9eHcSG2AC3te6kze98ZPVZ29a8Q1ALmh22hj2qma+BX+vqX2y
bWI5cNtdCrCvJ3E54mWDX7OzKoqExukmZbsI6weYHyOvE2nbKvHDyC+jQK7Et3am
hme5qd906HkiEW9WqDCvyN8sWj9wGiEg8lAuroWmfziCVp/oFkAhAkDlg6rD5UC7
SpSXNzX/5tNKcUAzSG9mAuaWY6KI7+DOBvpDp2ErCGAGqW6Qd1d71ZXOPGtVBU/K
h3Owxbr204kCSINeZr8OvZYKqWEcM5Q8vp+mbPcl1SzXQPtcUGsS+quSyp+PBwOa
rH56lI8GINLsUj2STKF66Ii1nfU6aAMEvCDNqSf6JB7RPYoy6rOVyaKy7oX6S9kR
cmPUUs8349lji46STJfU1bG4cFtt0vY8gj+G1dLQDnfa5qM+2NrjYwDqBitWtATg
b5Xs4MdN7QXl7/3jzQglqkp4TiCSpTG3e5lfW0/pMhtXc+v+Ft2e3ztv3Z2my+ZS
HtCpqQnF/HKy+fhR7ZE3uVn+QtS3hyiW3rrUZfu360rfvgn+uGi25O99dvapxDEB
TSYCEXDezTVF9uQNsyowcsSERsdDRZU+JfLR/Lzw8yoSZ1RYYtboEOrobs79ogL/
0v0opwW7V/oyVJP8g8UBTW88l/qBiQR7ltr36sMvsU0gnEL/cIBWKvNqUCmgLLrF
3KGmZRDGulUwDZGmE4SryrU6h3Y0S3dVPURuhT7VyYrDZTfgZMjGItb7lKqx5Kro
RQwnDil6uw0hlwMQuovVcPbosBnU1u4ueeRf1IbYsyBjsOb3VO77/3ZTgtrsr9Oo
61Oikdl4cXRp8XM2iDp4CTtd+rq8C8sYdhM5A9ZWLh88K4Hd8tr5dwJHGWs1EfEt
rNJXvwBVLzFnM5i/Ek401WCBH7wlX50AYbOlU7tJOG4SpfyQI/q4IagM21asp4Jw
cathOYq1Art7boDLIDiQCX/32J0RtQNQdJXpSQOuMwphY89HvAwjZP/rAojNvjbA
HSmvYb+0kyQDAatOxx1X/uY9BNSOvLxlGo7b0jOYWDcKTvZ89MhazZWcx2PyFCs9
U9XiXiMqUN+AGzbzaP0PnP5LXaXMLXzz5CchEBHXgRoWM0qqrWZdp1NZeFZYxv+y
LRnkZ4j1k7ylfaQ5LPZ1aH/x6YD5aOiMMV/oLoBEYKY3Elko8ZyHMFhiO+kVcsQU
44IwFNJq42M95rHiZJQiyPXI3g7t+HUWM9oej3KlFo2fN00beBh3dwJrxHv0+MiF
t+RUflxeS116EJeZP6fCYkYPEbsFOmNdczKl1SLLp9WgIIhb3CgN43MLnf+tYtHk
dupC75yBJLIGPaPRWw/7U32qPHFiCnRLvqCRg2VaYtHDeqjqDD1PGejP+UPGjDlf
kZTF/8zrzJwH1JJwAuOQOw==
`pragma protect end_protected
