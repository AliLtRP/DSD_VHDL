// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qq/Txcj2UGCobKo5DJQT92acoHGpBYKdYvtaDSNCyTh0MxDo4ZYEssBdg+esg4rb
0MNWGf3MBjNZ82c6Yw0VLjuRgV2jpTt4ct8e0orHqBxnYnHWwylfYnz5kjRCG1aD
mn9sHQwE4tt9PBS5BpkXArOlBDWSlK9GlIOYLAjSV5A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6416)
UEBixrfRK2lxo4zEek6PkFZHZ16T+Bw256MAmRrwsoLa6d43WLLZR/HxONw6FshX
2c5ZF0Y0lSt4YfxNfX/2L+eIBhQOyWS+PvZHjk0Msq4JAw9pSwb3yjl05TV411lu
7EvD7BcMiILKJv4eLFARZWxvee+RaFVoP/832eRzW33UW0ux4O4y/I0Of1yGCZO0
htfAspfgAhEGttX8RZw6h8gg98vVyWLVwalHGjycHOjXL0Bl6Vnn3i5oAMFSkiXa
8TIvlcgaJqLOmobN6/dOF2eXlVmian2O1NFceVm0JRMxL8mVs3mQ+l+lIvbYY7rm
yB/iqVYVlSPCGEkPYMGHN3IqbdxEdPubEo8cVwp2CkIlnDDB06fcFpNDeFHXK/sG
PchlBcvSdzacyjAQR4dEvgknNHL0eASt3phpwSH8Spp/5tlfom9PPFVVQf7zQR0a
B6RI9SQr+GixFAoN73CWzBT3UQI1rKYQ/IYrwMWR4JijkymPUPF/3L8OKP9Dwyq+
fetjKs/R+KA7kE3aPc0V4FIsNdSaZQxIdz5F55uIh5og2omIC49s+e9j3UxZnKq6
vancHFJzCVPWotcHnkj3WY+atQ6op7XTQ4lbf7gstY0raeF56siykwvwXI0/Jlil
V8PjJ8eF6REeF13hHyF0nUzf0Gx+PVPqGUZw6I7OWjstZwfT6265G/M5a9vkTqeN
lb+s1ekUfKzuX7FaOEb/hDqG/Uc2X6XDgJ0kted/6pqflr0rslb+LpuhRt9mdM3q
H/jKIvjxmM2b3YztttSeC37ibF2LhU/04AXbS9n1xB9nFisc8ffw/jGqV2e8Zclg
o7mn3Sa0q06Kz+DgdblIPFyrFxg2h9mKvYJubcM+BEpD6VZ8KbwjMTcST+TTZtQv
d9wxqaZHyjQ227Y457fZLc7axTTJgXkLzJAR7HfgQWQRon2NuRsjidBf6kUS122H
3owgjyENgRve3oNYEc1ZNVkMhHAaiphK/crP79ClEs9dWfoEWspozoKJRPpG/cpD
zwM3dTuXoLxZsynFUXPVeXBSE7N+h7mZ2asAY3FdXbYi4uc0CXZoWlu37LGU3FBu
U1Cg6Yc32VYY4vQS0HLlpZ3mrPJcBbgnKXnFhz/1dDnWnJVvaDNDt1+sceocLbLv
h3frFvZ9rg6VWXRoXjsiN1Lm5h/6shE2oVHJupdr4kJ8RQ3nIgcoYxt05MqCXxph
pPjBh940r9mD/Ofa2ar/B18TtU0byCay0rzc7ZMLz/2mT8EkxqhAX61HKiPwhIj/
aC9kGpC31AEn71QWFkCKSnqaLv5YKp9VUCqGA4+GTFnQJ3LB4lTNbNj0mdf2daj+
pXLiH/0LOxPi8GErKYfk5NwPd74mUKX75cc2r9x0z7L1in8ZGb28CbYF5hMo5ru/
yyPlrYVLvsqvc3sOK3uqfUMg/2KFjt957caqv4/D903Zne21wkh4iSccVQdsOB4L
FNvLkIo6n7ASYMKmi1B/kFvhC3Kh0ofNp+WN7o/XpiJIDR/dfEKtyNt1PIC5bXbS
UigGoK1dHFJZ6pD5zYwwtk+OfHcrE/+80NaKdgIEcumn0Iw5qzYf2rsjP0spZT8s
x53jox5EmM2Y9wPwWxZ6KVCqouu0mplTz0ctohFa/r292JGi4lT3M5Pnd3THzFzk
8hYe1HD3PsivL+/0rOCx283QWRO+ipwCndE91bYmV8AJC7fpBjg7P/iTkx3qS/jD
91Vk0ZarB6dLRxS+cS82D5RO6XVxEODZYdzpAglDTiMcS+uBC44Pkbbm9/9K+z3Y
GpoRfSyVJP+Sd9HMVnxxofYyVGt8KSXglU8EqKADM7t2liOikj9XV3i/iTeuaSeL
A3KSME6ngTlVOwYqd9IDb3OeG1GNa5BY6BQHHFdojtCwg0ur69+alI2A60UPckiU
1DrOqGTirpSBdLJ8h4QRu1hyAGHyUupco/DeZ+hLkGHDoR3Yv4xuUd0lBKsY3mOI
y+0vJY6G4tvpuFJ9uxkV9c4IkfqPzVWpcRwZWz2qfM8IYI2nTusvYH/I77+Eoh5q
n8GepWGv5gfJCq6NWfoLyz00q80ct5sAbrGCFbNfQVKz4muyvXlj33i9jrCZAVvu
vmFe7zyklOfd/nqvWpfPs+YKnEs6hmrR1nggo7tCA3ZDXNSEzBzJFq0AoWhXPiQf
YxJZKHXN9thAa84thpJIK5EONJ7ZlAq2zc/XTAbdK6zLrudd7rOFoQaP+TTJcx+A
HrNUkc0q+EiUxhWi4FwkQwySEVOkAIi9Qfd7ED0RNGpOQ3owR1xzOynDYLpo63ab
R/7GpKx9TYOmnz69rol3T/bmlqU6RVzcS871TlhhIHT5r1jfZ7yeYnJOLRXdNwGB
5nu7PxurDmrlbpxpc27lhRK28FATTXXesJgztgj7BssZaeHeXABOfes0QtnHS4Ci
6fnoTjoFuPhwANtgp0Rjd84V30Fx3ZusXTqXNnTV/4YRqHyZeuQccpAD2b2ddb+h
H9kr+QXBIv0kScvindkmKhk9PXwhwZ+O0RWzVdz62rI3yvfP9oEXWjTKGdBgFz5l
K9mminJXrkjuWpriPGmgvQWOHVydc8ia5OMFib/sI341OlKaVXhQDfiPeZLzIsdC
aHIf9PeAzMjs90shvodfmWjzM2zdet+tVL2qFjziPVqjNpa8w1FscU7FrBnUjkhs
W55zTILNcsG0U9hv/2RbEJvmiw9Wa0H5Is5VGq68GFIeMULvZySiDzR7gSPxvDra
rFh+8wAtXqiZOdRzrFRycutPVhpDqJfXpydzzznge7y1JC8cU1X0yACT6l/cIYWi
fShVPryh2yKn5RSwn5dQDYsGpWRc0RzuXSeow7C+iguvNtG8ahiJ9iAnijUVKlOW
+OmM0iQdfQ76gaOWavN5NP1Tzy3K3AibDPcOTDsYJr7DlMHYbuFeNx9j+nV9N4qE
mGlVUnhu5BjatDoF49yjqeHP6SLZdtdYy9iXSdiMd15RENB8hVzpmTbwzE45B+kF
aB4PI+woThI6MujprkbFSFgl5JNIFwvU5XdDrqbrOVWE4Lu1gGIwsJE++MYtyb1g
/+37y4WA84qd0Rfej1Qo6cSJG5zNOXYMZ9sdXrW5OWJpqI83vkh5Dg6Ot1T83fZx
X4IZYKvbMZJ0Etom24VvqKbKN7+gbp+T47NozYYxfUU0Ca0X7XArvHZuNss4DLYn
36QzQYlyGyg+lJfa8cJbtXJm2oW+kPScYDwX+DlodgktIK3M6i8HgdGoW2cO6dbB
WoCagaa/i54BJu7e0Bxol4f/EW+m+JLvSo40TegTYkUgwL6nz1PqqZ1vlUrAwwkO
AUtdvO1npVrbV3uloqV/lMwB/rceXFSDkbUht1pxNWvzHPEepOx3X0ACuqJaz0lO
6nuyIZJs2xTrVB65tDwX3HfGsAdm9Jq7pTASccwvdrJp+dUPqPgo4VurWU5tHAQs
kqnOvNLmYOKB9STyrUlOU8u87L0/fJtgziPS48YqsHED1rD5d3vbwiqnIUzO73N3
LAjrK3R2JhI9bOd7mU1fm4Q4bxWkNs0JZD3NmtyWN80E1JSHao82GmTXB0wL76B/
q7hbVpOOvK10ktdoySyUQCX4ZGctLCpBO7lLUNXu3KQCRc6CrDsX47ujJsnxQme2
dwtCSU9ZoR0gOiaykjWI4W3coNJ45ttY5EoddCqmRoscZU+Z55vwucQojh9bgAB4
8l2ZxXF1gmoMbjBgr/IGm1k3OHL4wljt4KksJ93s4ivir2YsLRCBQDFq2LFsuQE2
qzAjjxdXboW4f0R/s/OEZbbmbMZ/TwWDn2/GoC+cYjtQxvPs5A1g9oN3Htuq9TOz
av+cu8xhYdiF8TmykiRNWZFO9ovwK1N/AILpFDcp2zuK0pgSF/RBASjw6JIQmYu/
yaBuRjviowJFsmKKYtBkCNFxEpSGdn6b2oMtalSAtARGLKOcigBajbfkzoAQY6eb
tltTajsnnlQ+V7Vc77vsK8dZ/KsWqBSqYHY5Rv4Uhs3ftgxSo0JSK2y+7X8aJ7Hx
tkHbaph/b9CtKTrRamp2LMIXQEPHD9GsvR7RGT/V8+z2kfM3/WXf2XmTO/Qt7wo5
U+jhbFOso+3jhywRRTF0svlGTZbRyY3nDWPvjrIg9JkSHHwFHrOFXVg8kQ45Zncp
+TGFAO82cbG6l74RBh+uWwgBPIKx6NjShThcDmKv75Prensn1/1WC4EhtvizKVj1
l1M1yptOc95BiQEyUSVuRT04la5J4YJMQIf1icZRWV1dWPoalaKsBuWkAt1qhB8i
MXnDMUgaJIVBMswBBoXwPkXLEPi5m++PzqUpDYA1IFw0pcPQKE9cGCtCqSgHZdtk
wjhIkqgyc+1lWPDz2Ub0OBVdx2DZQzKQls1nIXX44IfPSNYoC4D9FUgKQtdzY+No
9zraZ+CI3keXHi7tE6fdakxGVBDEkkiyouYBcSzhUMtrTF6F+hnRbQvhTLKRaYC2
q5K4SrEm4qBZKfpMxBqsO1yphydAOyP3ELwQj5UxwwTbCl6rkn7mgvshkqb//ePw
h9qn6YNt8NS+82Z6GSroZtg3KWXNE7OJ4s3ahtAdqIaTu7/1S2Hmd6Jfz4/fHkm6
U1RjQlKjsRt5srYOG1KulLH4lYDdja4c6KX28IAT9KE3IBmpQYTmM8k2s6lcevsx
YEPGHcMJdV6Y6dD+kRb4ZtvXVUb1F7Sq+hAoXGMBYJYvjUVMkqFIFeTa4rzOl3FC
FeEBX4zz2ktzVKZHlJ3E5fnfZ6ZfArbHlmaGyJd7ABuE0UzIINEYbWvVvuIoWoaC
VVaYCRvvARIPX2H5YjJ4eHbx1RX8DwnrhAF4GjKtPaGGEBqhfaeyGuU0D4KoMPTJ
RXkXB0KnCgfarLyu80V5dfyXA38g2ZXnbb88QKKjeWR5iEIz7wM9hWHu1LQAvvic
R56RlQWEqq54wFrQMVM/nsk8nfE90eJxcqvvWhT8rcrkKxDH1d3XnaRiF7fXhsfT
cqcuVOkfxyFbyKD84Cay9IpoXgtbdfB8HsK6iavj/GZW5VaRnmI/fzq+W0vf0+II
XRZ/uqjeKUptqlP/pbFtC0sAdcabv/JSUDXf+cobE9BjJne5D7mnk0bv3WhnUs98
vNRrye9nochItlPZ0mAPI0BtDFDcNL1W2wWVQSbmOenRUXkOUY1AEUfXcFsq/vRX
cYNXURA5UIPL9q14YsZ7EU7ZVzJM5RbfaoWP0sok4IJtRE4uZeeEL1npqAlISq3A
IIk7INpt5oO7fexoNZFQ15Pd1ypsu8FCNNmMrfM+dulCHbmvgemx4W5jFe9xTSgU
10zDU4xkZwyIun5F4YeQdKNkBrSALPxwKXJeMgAYmrZs4AwelZvebdqm9niyeq2M
U7IrhN2IP+qCC1YX/KBFuPVftiJ5r+jcflCIP24fG7mfuIFco3KP41je8kManPdf
S5ngJI3kcVlZvK0fr5H+Imqwj1Gsb0a3RU6uY6qwqLk5j8yGzVgqc6z7zaogGru4
CJrYkVyk2AcVQc2oyfIE2eMxLgPAfAt4udpoonslh2Nc6HEYgO4U/6GTXmvs6YpY
6p/cKxwnJVHe4Fs+MMBi0lNfqFvM0Jn4QO58XiWHYd/kygItuKSBmJrj5Z8ZTQmJ
zQs7WutYQpNnuVLHD7cBa5sygx8fpBXzq6yQB7vGuva/OwZ8/pISywqH7WO0HUwM
Be3I9yxhF+gu+KKBh9CiXyLIB4B8Iu0Fv6V+dlknaY+8aoDyXbMqOTAKaPeXJA0+
CpfXyLoqqlIACCFZB8m1G+Co4Ox4VerZRPldkmLeaoJydPNKVDPqarxBi0bb0aRl
iZ87b02t/4w0X1iETiLq5le1+wfOOgxzw0eCImOBMuPyNRFYtPR2k7jfvgAWAE0D
Sy9P3KADJPuGv8wHjKIn6oQzZxfRf7PKDPFNyNaGZ/do8dnN3d3u37n5QGx4xOrx
JBJ2jLyH6Sm+BiOj7UCsE9c/t+uW7jKo6Ris3bGKbQiEvevLXgnCnbk5wukC4yW1
wyDWgnwpLqpCzS1g4QDD6/DTUvoxcQdhBglkqSsMxu/1Elem4/Ild7HQ9+HSj8Gt
eSg6/Vw5HXAWeFpW9jfCq0/FqkCFvyAdF5ORaEzJU7hQpe4lOzJRqdXqm5In24n5
RTabbiuPfnhY8+4UyHIL4aWzT8LDs1bY6282kjc0Nnb89gkZd1EHj7j6Py6KJjEB
nFcyho19hERuja7Q6C5iel1WY2NXlbdvrm0BAiaTUalzU/zKabKNntfFY+kV3U0S
n2RYV8XDcw6kbYjAxcKwOjVrafuNGanQkP/9OsLbkgrGu96Mh/yvCTQMV8Xl43+R
K9uH+rF2wMXx3Wc/tHmZGG1k5WEmgYs+jVAjlrllT/I9abyIo7NBi8rBlNghfbWk
AAs9TAJfCpVv9noch+UYWopj26z9LJ5eqdFhUMJLJEbIFqAx0VJwNJ8c6ruYrGmW
3t+FIHEU1s8eyICB7aBPS3lxzRlnuh9978XgXPHqxf81hNClY1QlygfDd3xkeCAp
5958SSM9AfFUBHuOM9Gw8yRsZ+36iujKU5Z8LqPuaHKqE/D7GQklktLxBY24jnDF
53XgCBJemU/13QsnyAwagzEt1tJ6PhdiScGQWtRX786kzkrm4vT8t3Af5K+UQpyf
RBkyJgKsLVFFT8zNkrg0kaNeAdFya4Deo3PhkEZN+6aFqR8m2VeisBlEd6viHrZa
qJ2Uj3OJ5tPthgpu4shQTEcHz3Tn0nhm9nHOPWgAET2FohPXEragwI+2P2NgPuVK
t1vIx8AHF99uhSxWJje9q5UAZyvhMn3+GDgffUqjQd+4IHmme+O5la49SRAYViD0
z02iaTPwmPV/PKYokj1cbajMkNIBuWBxE8WHWxTOcRWIipJR0+ixJrO4MKajmsto
dDP/Nw1SpPIRMo/vhx01RiiWyoFbH/boUJxSbFz06/Ob+/3iti49glV0x6yTLTmP
MPZkUmHW691K94Y5rJxGwVU+As+8c1YKs9mTjT9BeVbctmYvZJVJFtcJGsFqX5Ti
6FAk5ATYF63KMquq62sYvd///YhoPPFm+ZiYX0Pnnm3hdhGSWp34YLY/z+JAs7eN
G7rvBw7V2IaJlCbmvc3ngK4KD6NpZdLQx+BSA1B+frHH6wS+ea7kXo+wOCzUYcwY
5bUmR69Q9YEQT0uUxkivWA9jWlYEBj8hL5la2rMbiklQA8dl1wbTMTNKL1LfXP9L
tLhw1MR6bxI+WvImn7VMUN3zNkfYO2r/H79yXowgaOGsYLjUnlf+y3LqpwrErP7q
ikwQDIchEYBU3lMdZGqZcwWF0NUCifLTvAWi7V2dGjosQitXbfDxP6zIoZbWsxAy
ewAubrayCwq6DoquZElhmBSzbINtTGxVqdYrxVC4p3IvFqoV0Z0LyvUo3+OvX0Fv
XPAyhYEK7CL+jXyCBiRHa2/l6u/pJCzw/91PFA8bjnyP0nW5jbPw70gP0kFctfno
PD+4Gx+p0Yk2t73GY5/mdt/Jl++1WObHV3QPJ8jiYfB89j4GbS/cckh3gl05oHbC
g8DsNycNf03IXvaRMblfhnoPuv/YzvVty6NfCUxPtyNvezllD+sLRUQz/0iYBaob
qfxntDXiSW//tqaG6G2Wue5TXFs6oSqTisxKmmWj2Gu9kqS6vIF97p+Wk9NK9wNQ
xUIS/AuT7CUUWE8fnoJY0SR5fgg1NyxaJa2OS31NEVjCoOmKxdNJ1GRvgX8rzuXU
j/dVC93lYN1nJQr++nTNGFEtcYvemUXpECpog9unR+Uw/p4c9O3disOFdLPLDndz
HfU0ZhFfU4QA1h04QjCGgErx/AbbLAOl7bVt7fsEVFo+QCMipq9+MnhDbWqSUhsQ
KO8tDbKtZ7tLXiFjaWfzCBXNeS5dj8g8v9lXxaVsjIwhM08ujeWPU+6+Y+TOCRg3
sVqK1o0UKP1++LNnQnHNa0bI1Tr1nz6uQjGtpacxC5KfTpQV7896O/HJpBpAtDHj
9mpdW6HupYvHBn0Owg30toHISrV/2DRJRXtvqRi616hAnbz9pplTuVJo3acplS3r
2wnhqtD+FOoIxljW4Mganaj3Ne3tCpQit5/sPqh4gR35bxuArPkNlsOH7eJyBReu
Gbl4XP19+cNb62VrztHNN7C3YO2Tv1v1iFNu4AFjPTpkzvaYDwYY/I+vTya1lRQM
8GaupUjyVbgZbh/d4bGEmgWYeVzzksLTR6v6IbhxKhj4iWBafg2br65YqXGqxI7Z
NOCY7FZB2zRbzj/BALMOEz94szRT3P9qlbt50+HEOFbuwXJaCsS12fY5AX0DVWe2
ZHtUhsw/OGCbKEY8t3k4qsaK/6zY4Fl3JNgrfCxc5qS70kZ6ukfah2BpWd4S8OT9
N4pkj21LNDw3DPyNn5uQDJQfiaB/WJpI12JfkM4JsLsQCtcKs1xE87xpwu33OCVs
zn99oTbypr186CvBfV0hcHNQ+uBeRDMAWrB6BuXNqsSVUm/aN9N/Sx5aU71PUf+J
r4snyLpJJ+tDxcmJ4qWsF6fnYcjmqonBXKWzOzcIqoI=
`pragma protect end_protected
