// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cMb2GsnsgbQP71+fzkf4/x1v/sY+6gAjCpobwGn6D24RKSvOrS+tUOpx7J2XDvxo
v8Z1sNxvo4UeuXhBbrNkS+HbEDryhyIDrk30fyu8uyfSCoUyjlAGZzz+Ju/5XPoP
3ni1hedkVgW2CqDNZhe+xj+zzU+7ETIz4mW6J5WVdY4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28304)
K9JzmsprMuUxlH59FtHWyI4oaVV28KqpI3qIQedfWVV8tlelntDMcOvBdO9VnrBM
6LcPVi3xs/8Bxw0YydVw4yWNzbKmajGIHO+eTJvtWhAMBXsqLyuW4oSl4wpIf35N
p/oHx2XNvlONCKUK4IfRDDvACcWML7cK7qbmEKJDGKpCCJoYBfHu5Zrcgh1Btco9
9kYUQXFxnfNyXLNV7zhwbDcweMaueV4r/tcXzvIdFPgokS9yV8ar5ZVg8otx5PCZ
mKWmgGRT/noLkPHTz4Cevv5y3z6r0ucONL1QqaXrh4buHFzS1AWywhWtSo7/6tn3
kpCu/5Rq0z5brvWNkDfsDG+qvWI6F2g8CMxzdLp6PHVpKCqQ2GyRW7G8XNcYtpMC
kQ38ck7XtJQ78wxS6pPphi2D8TNuBM/C+6LUg6AUDlDG/FPNdMoSNzbH24w+nXMy
N+JjlnGZh4+l6ojY0e5frbd+rV1rbZNEph4EaTTWXSeggVoFFPYnaUN0q0eXWCeK
tp1Oa17BrR/t7KPNhRRtDQ/2yt8P1+CbHFDHEGiaSzEOsiSjriM6F1z+aV5Did2d
sDr0xk0dNqoP2mpaIWgEeugwK5IVixxg0rFTd3QeAdBDrcHPjGYezhxlJyhLC+/4
n7n1jhG4+YErFTviyI4A9geClUXbv1RtHgaoPFJtZIR+bmzlgkyimevj6jpxlVno
yiSP7n5JkBTBi5seCIaJDfX5DI4RjqEE2bbgqzJuo6pTGamlwlsRhuznlGIvbMcd
Qnx1XYJa0NBpe9N8btovUf+H4u7EBcmbav6sxOtKmi3ysEUe7VER+2Es+N1MA0T/
swiDAuUmEy4/14KD580ZK9gWmVcP8+mKNzUuaOfYY6w8f4lU3dFmpTLhv8EryZUc
WSRDsYVDTJGHhWBLVuymVEUKDbiRzeTadSJovH74pRRA7sT4d7vyxIP2LZeliiWm
T3L3pnXu22dEUoTS9nDXKtPaDqrrnt1SBxbSodYK0sxji5G0q4Abemt225iGQ/EF
kL1a4zDVSjtucQpCsDuNAsk0y93ILqCfAqueVZUXPPcXuwS53zGqOxpWKRa25/gn
IUeSg4ArYAIN+Q7N4mYcfwBCjK3qAchtYoHf9VvDFaylEy22KNbmoBIB97xf/KGX
SPqMjhUcRBlQ0ZV4vc5QrBd5zQ6r9y3f0nlWjKwuk1fLOhYJ+DfRzAURKJtooVCQ
WSvBJmo77cj6MRBbDRH5+LXkq2Va3gOMhNvYizJjui+I19WqpgeMnKfXEjinlZWF
ALY2bpH9bOO7oc4salleducyicI7Dgmijb/4B77sA5q6vyV2grNiJyLH/4YbgBA2
wwEKKwLnneF3vYMD7HO4YB30FvOIhbHXCIAeqkpo4/JVvdepRGRmy/X70QedoC4o
lqEAlXIIl9iVxPuITMwsiCDPZSkNQ4FA+Hr9qE29MkEVdLP1M9VvUQMBlIB0nwaS
jc7gDKLToi6B3HsP6fHX3xwPh7LguVbger86sgwnrus6JkY5CXDyhIkD4g5/LO28
pxtPqW4AY+0feRQGW5a156c+lhQgXn6a/g8JQrQZyOBZPXrNBj75dYJeN3PVvyrk
5XXMAeh0h4mvuqyTZIJlaxsy0TaGsKIbYZ97YrPrm0Y2J+mC3YLo0xqF7T67SrBG
qDKzunpjWlm5PMIOVBYeN8aff75aPi7FLQV1H9iVpQPAeE5V56AAgi/MCuRf8Qp+
pvrHSYoIp36Op0/YC3kSPtC9BnxbVWMw4Nyq2/l2WgOuWjRNDKRGyE9s9Ri77JA8
4SLiJXgHhC9dFqPUFLe2ma/0cArBnCbnPsavoriE+OL7h2m7YWBfwYHkayLmMryR
uN1qL3hvbDvOHRnIOFDPSIU6sm+5IwPvSvDRxLdvdUgDbW3yQWNmr75oBRB0YbOG
UqCFpVrESqLvD1jplVVbiOxTPCf14hq1UQ8VJoAbW/96bapY5qZYOqIm7n26FZIc
dBCNMi1bLFECLg6FqrAC8X1nhdBfeKTauxrJ9gDLHwtLz63CILi5HwsnzzDAoP/2
P4QUjE0Dz/06WFRZursSnwvNmcInvEyKkYaGWyfaHDYdFMLG9P62hkGlwwgl6brh
6/JM+nGbPNBZYQxM/BLmqWSLlarRjCEgxfHkblPab5FLei91iLusKB5pAr88/lFK
zocIMsXC/2vqSR1CTT31j9o/TLEXkVIwAXeztj7hx0jziLYqdfpbyEEpx3VyK+iX
zGARPrkE7te8v+15uK6hsvdxuVAF8nyOku8vRtmYhTup6jIV8oTucrtImMjMkupf
IMxiuELBrWEgTVYvK8L30K9ZFBQj/9ufg0A+eC/au69zOiEp3evg6Yivryenb/C8
BKQFLdONo8oqA94OT/oWAnZf++ZFqWDqgQ4xM9XUicMMaiJPt1RbVyKxexoOWtTK
fVRf1N9Irqt5d/QmzkdtbnQHiY2AOQH2c+zcTWIIoG/T7QiQXvtqXroC7I4bXcOj
heDmYwLsP7Ae5s/HUaw/T1XY+qiajVU1RrHXXvCJY1f6b9dt71evy0nYdf74DQPf
hL4B1ohqo3PmVxn/L9O9Ku6wqi4LqIyAyYTah0Jw/fkKwYQnDWqd8WUNRjtTuk4U
UJo4Rdkc4HdnS6zSZ+gMZiySo0erYZiKEY6r+kUxgPzh3AdtPaK5pxz7ySvX3Dzv
eOoCTk5l2eUtOPacEYGr2weZcOpImhTN3xEee6nbzXL7WGPgw2fzacPH5OG/BYaV
qrDnOGnJhHu7DwCly+j/42etUo2q4X5uczAJDHGIiAEITF0wTBKiqaouoVlqYDtV
Ue86p1TTGOcl5BYAJaQyA09AWe7H7zkeSzONke0rW4lLo96a5IgVBqNaOYVsk+5E
rEjmu+dQj0QBiVErxgjdGydNueysr0JimTTUQT148lEvkkV9dPPV5LoCmXUvYYNs
kIhMll6VmbT58DZ3JqBdplh1wpdGqiQDK87SOkU/iV45JnGAxHHcGpztycYGtvx8
dQAOkMA6czpki1Op1DGczo5zt0OHymFkW3vYH+aX9tZzbiHyyv749sgKz1Fjphul
IPcf7unu+dd2oeNGm+5knq/wigRm7o9p7ZmmwJoXhgY6SnsjzfehKpOujLzMDU9C
P5s7bcQBmihHFyoVMjSYBaHKZ6a/dVT6WYW2zwaEUGCYlpfQ4FS3TfWH95hvdDSS
EuNG5XRF8ZeBUc/Hr4xm/NYNb5aI37KSN4hVmM8w6LyQj2ClkxQzmzMTcgWM15jy
bbQ1OTSy0j8SpZ+abWB34vWmizBCRhd9N2MWE1X+BJG+jF/WseDvvH95C7+bMhyQ
wdlX6G0CUf69cohVrVwxeerzmUD4oez86wQhKvaXqMOpBqHMOlwhD5I969oM+Hqo
dfnH42VnoqQA6J7o0j839TQO0WOUHQpZyEZr0ZC4i0kyAwyCMNF6FZfzZ3KpkAOD
4CH3+bQAbNQYmNlmydhVavreBdXSpVxlyGxgzL3ykugRhTAPkcUjL2gxm6Qv+CJp
tnGUUE9NxPJTGUAfl1onhdNeZ5wL3dABGD2NtP5pPV3YvP5G7SDh9HNDiNAkc3pr
3kvoXCSWiOT85rp399Ai3XSOZpF/vteUilOkYX11MSnm//K0I36EZCmRssUopVL+
Fj/YgGc9BjKhrMG/l6faz8iYjhpBG9Rf+z2SOSfPum7sFwYQHbqGEZFLyQ5zWLj2
H0Z8PDrsYWDXTBjWmcslr4dyggYRDnMAdQXfCRVVFyOvLaWzM+zuEltYkJsGRpx/
QG0aalMCnVfY0/Ck57zvb95XRjh618OU8fFAqKDR/eKCecmYfch04DmQ2qVQ4Ytt
IYoLvDAhAvcKyz5pODGNaLiXkhoh3YZHK2aPPAIhkCSaUKPmn2n0P+4jBxGe0tRJ
TFDrKfxL40NxKVekTlbn6QzaITXGEXzfHzjBe9/mvGx+YaTy5YfmEnmC14tcvFTK
9JNL32PgrwwwiO+JHenOozFRDtuTOdQnk/rYBPY8RMwZaXxt0ErnGIYyFIpF6XmV
IvdC7VK0xmAENKsvl3aRwLYtzg9aVwGTOsOIStzZn8HFGojdS5vKs4gz4LyqJI97
pypTNlk8RCMTVitwRTmvokgFCc3GrpSmbvuCTMLyu3p95X1Aga5f44oxyaKBGBFm
jL0gIa7tl4DkaZfufFDO8kk+LMy5arurhU7O18R3jBWnUnV3b4WYHlZw4T0h7ML1
s3DMC99Eaa9FBMpzsKDfCZsrfTCQ+Nttg2VWI3L85CH+RumZP9zMQNkWi7YfEZAg
v8uDMSkS0v8nBMtydDrggdGrz6kqdpHuRkOeAwXgNAxLtzkLTDNZ+6Ojnob6fLfe
FAb1+oJjK7tCNVg7kWFz8+ksgfPqIhywpCN15AfftOnaVXCFvd55FYQst5maijF5
wAJ9SrHRS8iwX9xGazvq/7YLnWH/BhkxC+mQ1Vz5XghU1JoTA3pWjE59f9BrDVhX
3JIu70ouQ0BQVCR9kYgZOggRBer9kVrvwXLfxHmaeHyC40NyeBXF3i2tCXzMK+jX
9kyNk0LUZbXzxncsLKvPXD7/N3loiR6r2VlqJ7kOX+xGGwnIldYCHc7RNI2vBs7G
CUS7vWsPzkKYjhFDf/a7yEVQnW+CJgKhVZH8CSJi30E92RDb4NYTL2qM61LMxORB
dTJidkBhaj9j7Alxjt/Gp80VtHL35UCD9DMgwDdtZCDPjjVlp3pfBqqKcTdKvnv6
ybZ3j+K7dA0oeiWS91RyCK5tKRAEgKlurdU7mS86PM6MSTdSBVxmxwXkL2Ko0Mx+
NE/iSDeckWZuRKfKFaQNOPnPWK96JL1kbZmS1Y5MH0sGobKSDPfSTc0nMq+a0KgS
qoTxpwpBamCPSpaLmEKwE0RWxi8FVWeMA7xbCoKMLPijjfgIs1xQu2IxGBFwXbEW
sXTzrZVT+57Z7VoBDc9J1bBnu2CPhoaZpWGrOmp4TU2GgJ4ttc/Msy109jkubtZh
HDpilLb4Z3B6hKEPqsk+A6wfr4vXqxvv3kGZNbAQV962Vfp7CzKFLswwSSAkToNt
IxzSuEoZVEkdEHGcWMUrmh7aZcwv8toGTTUag/v/4GYqzjRleX4Cxjs5xvAC1vmz
8B2DKHHaO2fTjOmbnD5Vp8213YJshwkiBdMrOBekcHzKiLDjOFXtcIaqJBCCcdVk
7F7BR/WGZaihv+HQPTg9NGDj4F2w5KqQSC0byKblGt/V4LljzydfSKapasXztEQx
GLZjYK7xiWfCnU9jPlOAFhAI/CnMUaEjSBP+/j8acYxWp8O3hKVy8clnHPbc4X06
H2KIrDy3Ob9kDEn4Z0LM5ZAsLhzFEMmx4D/rbZLauEY5/Ao1R4MApwrX/RSCDItb
Q31KAnTpuw1ULN+3bOT5z2GZ+AekW2Vbo8rn3B6sthBoMwqNrJ9osV3nxgbDDPOy
ZLIw218/cB9ONquVYYEGXxShK9AOalSLCG9qegdDfrI0MsTxtEXFlA23Y8n+YuD3
Msee2rkLFuHaksL/U6im3iEO9zYXfa4pS57NOh3YMj73EsWkP0Uj2OjWaZle0xf/
72lT/TgvvqVQnCAWKv0OXpDVVGLsKON0vH0BhQoR18reUZZYVDAStOeCpoPigFSP
8O380592ti25BK4Q48L31nmaVLlvSUgC8S6fpOLHIBS8qhudgwOXLzA3Zkxwfqh8
vMQ0jlFx+VWbFtioWC75WmTWgxAA/Ed1gsaE9PLpdw8dIn8mC5MPydKuranmHuw4
2VxqBNz6yFBW9gGSjdPRUWUEZvAOVqvDIIqS69pFWAJjwFtsfazdXeqcIdEt11O8
ZziKNcxgQO0BKvFyW27jGLzEi12+caKhbkLmBPceuEMWtP4j0hjzS9kFVq7d6RYO
gz0XhQeqwKD9Bjb8E49+wjG22FKVTp/oCeMsIhp7IYgJ3UKSzdnZEdEhcI9eBq6v
WG8IFamd1wRbOKQwWWRNu04/fWFP19pKrB13D3Dn1waeCIyLho8zUZtepqWPpc7L
bYZA2Ww5xUNvs9QmKq9oou1Ycr7W4oRN+oVO2MUW+jluK59bV1HoMyNWbzkCZSwu
5Giswrod83Jrz1OZrdflzsjSzEvlRf0oPCUEI6qK4aWmx1PRoUmIPBa+45Y8cuoP
hjaylUUtPuFGK8dDAPRofMvjltc+2Na/j3I7qiwM4hLPnGLrwfIxIR8hIhycpnSZ
MMlCgqXI67+URo4FX0AdezFDD8mx9jMLlr/oFW6kIHLqC3E4+hnk+QMdOsSO6AE2
7Wx24jdUzMyY35izN0zX9IF4MAhtLlBQ0ILBuS1JBoAl5I/uW1TS3xgrmiV3ZQZb
hEd+GHEyaUMsP08/9hPDFpXggnjGQhvlY1spvBiAUGHsck5brp+hStGrElgCihyv
7nQ9DVwZcxGIUz7TfF1A5yKAafEredFOdoj6UvkBil0w7rYRJTyGuW7A4ILQm0ge
utfDOWwOWekkYklGX3Nl8Dgt1tC2Umpgc83/H+jxmllD/3mMFx5PA5z29pYoP0oP
+thbf2zXx/x3MfbhGQxmrOEyJZrQrg9LCzRWDXVg/63S8bXEgif+UKMMmWEgIfq2
WyQLZbNDSLwO8E6dANN9Xzjfi5detkX2hch0Cy7ORaXEpEP9Gz9DAaJKaoX7PTSN
f6QTrDyl/fb0ep03HL8b1BhTw4E5x+JEUN67htX3Q7QPg41Bd/JIe2EQmMsXSjwA
rSHwUNTEOQ6JdfKjVRBOEdsrmxvY3pMydN0qP6Q8r9QLotse3YHhMMrugd8DovDs
IZo4+Eip+RU4weFkiK3N5TNrNKnFlrRekCgc4TyO6fs+I4OqrVEN9yvl1HSw8NJS
nCQjEGXO/wF5zM7Wy3vdyoMSNo7iYUy0ANpzkAndqw96b9B+hnPMYBt7E6am2bHl
N88MgTqEIoelWU0sIDFrDyr6Mb/7mWg45DXhkbaJ1mdPtJjXKd5eQ9SlMPzQb801
8FGrYgnv0vR7NcqctamUTbqblg/3flUHU94Lrl9tU4Mpq7PGCIDSCULdznVZIba1
caUJ6jenrBTiJOOtqu+iNIjJUz8aI3eVT2igxJFWf3SCcVL06scSeDBGicmAAhbv
RHXYEAmKmdA9SorZ3rc3oidFGHrKvBQJlIhF6m5g7G/xLNrqfQez9TnH1u0JJ5nW
MX1trHk0aosdmr65F+ja5c0Zv6X95tLgLBuqz3gKPyKc587FIXHgD9rGMVEiZolk
V7GazqumRKAHtRL7FqneQVQCcH4puhrMVjQqGJ0PYdQJyDe3teJ65QpH5+FobjUd
qyLDpsLB6Bw6YKeYS5AK2EVZXorfcXhWUpUpxRkCWlUbAzNn4gjqS1Z3c4S3kL2D
mjcQ6FXQSj1uR5y+PDRFn/x8/2rVMiAiHxplhbCtN3zEFdpEs0J5itIOitVdcqw9
PtQEYnXtrdw1q4sjM+8Of/IO8l0OO7oK/l7Iq2OTDvscZ5QfbtGqcnR9TNyXHQGc
eF/HeqKWv8PFm5PTjywxPQHCbopZqFXKctvdwMB3mmLe1vwSQMKxvuqwABGFBRz4
6coTTpAcNbHDn4k0UBjo4uClBv9jxJa1yCJA3uY6uUoPqxINQS69K+6WbD/z2LhO
rWzx+gvuPK9nTCz8LMIh5Hd/bHuPvfKmTsr+U1VM7sgnuFZObbCoGj5rQiH1vSvB
JBI2awwJcUaPgy/yCuLzmqq7Wvx51yDMo2qt9wNFVP4hGqGbR6EeR7yBFREHA+yP
QVO1IoUcW/YY4e9rjHAc00znDsBvwwBqhV9VTNj5YNTQSkaBTAO+8+HiTMEg6Ble
Kif30ybL/ZEwCInoUxuKRrqrk+OE5+5cHmJZWBP/U8GlAJa7xd68CtmurybiE1vo
Af3cuZxJZZWNRVtySRypCIeTzrwmn9RhXibhYX9b5MyvYthdUDmaSdTC6hbWYA0A
3K/9+/PR5uxMeaxMiJEgCDTLN8ygnfPrmaig1IooL0Qo9hRXGeRsl1dOQPuBj8iv
1pHzOR5w1X6K4W2yKaI8nt/8zmZucJi6ekq5OC/Cag6fEyhhxPbwpy+dvaDiootV
7WeEDOuU1N6qW8X7aFwQ3MLbQaX5WT6Kp8H44dXMKctPRtvbV2kD1lIkQjFBf/Q5
F7ENUUX82uq5GDMTnxm4uS/CKSpp02TOPTN/aB0YVSN9T2mitAfi5arfRMyxKFtQ
yA6YB6+ru4EM7qOhWKpCaarHBDj9GuAZS6/2gGhmIZXhQ5sK8Unm3yATiTsVkkdT
FU/zVCFDpfn+HPc/d2MZKrOgctNpdm1NDEbKRvfbouBWQeZ9D+iBodgsUMxFJUST
1Va519iCSNJ9weydfcd0UeigGz0+YUffqHPDkSIIA0s5M1u+TPM5+RwQHYw1L60O
LybiOPl3ZJ65wMs5ARJgB80CNO1tDoY3VjjVQDbBRVmbV6DqT2VaruUnNphlNPPT
iEIOb8AtjfJ9lUnB00sAjp37SGIWEuXLKXraYux4f/9xE6leyxfXcRaIXyMxqq1y
UNAwf8HDxcitTCnjkCiHEp2fBNP8NuhFr2PgW48CeGcp+jE10BtzUpq1jo6nb0zI
BIO09jPmeEqL9CQ4+BTH3m5/6sFjq+irj97fmUcvOysqMq71Dbrg76gwFmFCUocy
fXEfC65YEjgfgFzUojpH/2QrKT8XTf/MA6aKW3aN3XCPHEzBD4ze5YpdNxqYQDKS
uYFD4eeoYizLErE+PtbEEZwP2HGWsu52evj1j9e10XyVXQ76bfOUSnshNyQL0e0g
z9aalIUG8xaWZjaD+EfEbqp4RXiGM3B0OH/Ygv6VPvLj9oJ/QTecl1Gu6ZIny7to
SN5sXCBAwTj6bYWFj3kNYoKg/73CB7ZCEb1w7uevI9WHM7BqtM726rh94RL0LZdP
qtvhZ+5bpzBgmXcRNYLf837tH5O9Hi1OF3XFtPD6gjJHug0SqJvgOUePnX4TBOL4
lIUbcc6K+aEsDX4gA7jcJxEufXX5yR8698jyvTKeP+8mUxcKsc9zQrIUTxhU8hgX
mTN4q7Aki/VJW1PsRepuAyyE9ZgEX4NA5oa4TZ6RHujCPS1edPkBBfnPuEa6c3Gl
iwyGn5ZfmBNcD12HGctCOwffejwGCy+vP+PtTRhEOmgc4yKdodt5D5RF2k2SZ+6e
Vxp4Ml2jNFGxzuCzK9XDsRhaBaMdGWOmcWWkaiEczLFZNULuTo0mioGKbTl9tK4b
E4ZxRyLlYTHQ0EmDzo+XvgHwoO8RDOn4Klqjva/Dpl4cxLmLetGo6pXhgS7uGYQH
ngfq5pgU5WcvB07hBR+SpXodLkaGFM/1EdDA6V0uW6+mM840GRIt9XfZ5eMt0geG
TTPHt/9YqB5p7aPzqTBPDOrdzayo4EM2hCV7F7RgI7Cm/cfzP4mVmozrBZEwipYX
PNJZLT6yoUiWlhN7JwKR77+WHnRe++yNAE2FtSioHH0pje5lSuA6tsl/cXAkCUxO
aIIe6jkdbKpuJHL5z3rPL1paNnYwbFeRvB4g8D5hMVeODMffDDaR6V7tNyQa8tE8
kDkmGROu4lJf9wKuqsBMWuUScd1zmmu4ODx+c7quUZlq8hCDTjaC8xr7bTqKDDa1
Dr4MIirScBKHpvRsWY3RoI/K7P9jHCuGdjglsDSDOd448kfOkVK8XsMnUYG2R5dB
TfJhQPxDD3lJIfAdb7IElB7Yo4WgEHl1Wqx6gKjL8348vmTWVn46zpAk1qn9lw04
mR5SsdzjSp2SMCCgKZzZ2OAPQa8tcgB/l+MIZXYVgRNh7op4cw9gtxeNfyT9q950
qIwJ7MQ3usOoGJHlpF9U01byVHYs07wCP1zd6T53B0M7A+X7Oew50qH/PlvnjWxr
x1Zu0yTrAGm+mtr8GdSd5fYlAquarnL+WYEEpLcDRfzCPsnmGxxN4leFRxFhc/M6
F3fmYo8JzAeRjtO5JvolK+3U7pkguo4GjpDQL7h6uPBa/VqS0mvpemKQv8xZ0KPM
B1yltaiFg8CmcGRkiUHG4u0apslLcKkdVe0a6P6CVoS9yf0IS9bAKERQoH9ASqNw
bp98GoC0Xr+VK22vTT83Vm+WaC/KvYcVTQFx7U3Atfc4svrJ9868qEQD4QhB6VE1
/CsyVGDb5LROFZI30SeZ//6wbOvTAbnM8D+kCJ95D/146gLUMhpsNM0OetrQ9mlL
lxf9/wwHF+q1OkECXzm4Kb9Xmn9VohFAXaZ2iqiBhswRz+tjPIygBV/RhWsZ9rF8
Fjvl3CxCwcd/exrNidbnH2JxxD1wckqQQkM5q5rlqzk40joDnaoRveytHBLg+2pC
Eutcbdx9KGwuahX752F+ZTz/O70w5ce5tuZ8T8MT20K45ARG/LqV5zbLc+LcQ13p
s/GYFEm4t9+5YSQc1Q8JAhhVfxDF5+Ln5y44q6yqyrfUVFJl6trB4YAcjUQcfWV6
2Ho3Xw6yQejTP+IyWBA5uuraJfallnShDguqJfZoGRKB/3P5n3kaZIS2zy7kCNaP
9w9hYW1Tnqtvx0K7kzSaGJOZ4RL5+GX0Yn4+D1h5mdme63VTV8o3aeddPa+AXBEC
Zq84BxYXS8uafZItYCpgUkTWEaXR1qSqFS9KP+tYUohry88y9Dn4IY/ZpgS2tQVc
7cr920cN9rP9kHx6dAmDiT1mN89pgZztHNS8coeNSWuvJxKyjBp4w7wvrnU93SyH
wq53sulj52WEtiPqcBpC7Wl0bDhYizPgJd6DejbwrIPRJQ7Ex5YhDWns2U1jX37W
nN/m/KVd6xYg7emth+moo02Fl7T/53ZgnmzKUxrCiinZG8leHb+KMG5FPGZDFx3I
vASGjBHGVEnfz0luPv/dtx7e7KwrcW+3vucZInJVIMXTNg/439FUyvj37qDeNVM8
YhmVGs7oAx3DXsaOH5J72Y4KW1m0QxDoD44jIFInApw8YZxIEg9fjVwX2RXDRBXw
4H5aQagovaWJxStoF/kD4/3JAOtGzwT+awxqRQhvXcv+jmRn/xc/9Icws8bISIX/
o8H+Pmk07malba79Ig82romWxDHokP1OTASJqstE3tl4AZpfm6VrAahC+Ci+NDd5
JIMKhTjPfscKFsyIn1OfHnIBRWBMe9eX9QCGmX5/Sd7hC0xI+cTOm8FaxGQnBX1R
DA3BmW3S0UE1RU1dWf0878jvkXL3Z7T83/u9EgcNA4unfOrVv3ha2me8DD2kHwZw
0emtdj5qzH/zDZzKS71sA7RbZR8T5PBm4VzzTcqBjs3IENSCUdX9IJfgX5D3FghZ
Ee5E5olHnISsh2+BOQan9U4wteqfXy/muBg/NshY3oU6y/F2q5ktHy4rdIrYyMJi
CNFtQMIaYBaenWgmUvpDYeJQAncVCuu1lL0zX1wIm+kyJiK7ejyQoTtzLGeffaZZ
6zJlrLwoIUt9iIR2URoRh9RKvl+SODO7qIAUyhxgJuoG53Ex+ZN7hlYMzROzxO8/
ykXQg2Ji4zmQV012c/Vl6M4bFm1EtQsrrg/NnQePUq1kpIFT2XzF2opi1+zYjDn0
0bBwAnDsT/O2m17FuAmofiFXfK/gy5q+mZpTlehijjkQlW6oFAgX1NnWulMcUM/1
T55PW30VtjAkAksJ6LEEneDFfU0W/88d2RD4b+uwfwCESGSvGDWit2yK+hdHWa3n
eht+nVlHW61qX9O4w+IpHOkEnfHtyLNbv1VJXdzbodoKqf13TLNFMOnfIeduhED6
l2Ro4PPDYHmc3KJsXcWG+n2XNWz3JvY+9siSpHTO/HYRqpzrXBFW6WyyloPPC/We
ZY1GeP59nVzcnsbR0L79jjquvKmmYmznIAfl40fYzDv7N6xcGmc3aresAQRk8Ni7
7Ytz/yOe7Lszx+EhADB2TlsPEjC4lVgluMAP6N6+ZwUbt4d6EmXgX/1OlUcT0Kom
QrioFmeSyXBYdIte6KfZsiYfdSBQU6L/GO/WUuthacrdvAn19rxTaBTwaJJaqShW
/g90WHQ4FsUztQlhy5RBySX8/EhDE1lUiUwauMcwv/7FEBTI7Oc+xj2NnWw+9VOT
6xGDPralMO8B8CKF6L6jAGquqB8QqaXROyJ3fDWkYlAl2iWHcNgIo7oh1iwfRcKh
XnR71ul46dONzNI00aiNolzb2tw/0maDfZB6s+HeWyQToMztXgMSV0+mPFq4kWs4
fbGzssnsx372bQTQJRub2XFy8cD+xY99dWAYh/orojnHo+79fMNICfOLTX2vQIwl
kf25DP68ItgAJEmKWWKTIXkWcsq11XpG/C7yvY5kJ13YF6nvam2khTQ26+5HFyPD
BlJWEZHYAZ/92kSCsz6E9v52/5Mm6C0JrLP4lZyQolRRF2J6PcaNX7EX/NPAPbLH
lMR3kO8h2v7mpx9G/xzF/CdRHhL9O4NL03XovwKB8rHrVw5hZU+fUofRqQtmVFnz
aOjnzRr99x85+JNnXJim36GJ6+IZtuaGvl7HZHR8VYU6eBmKl/MaBpNivJENcCxT
Ek8f4rt0CeWd721OgfN8/K3WwBOyaSYLZcAKZPVVkXbp3suVXTRtbZv4/qgzFXx4
okTdv+QyDq3Lf0iUiKbYvCakY7BicRYb8mLZz3blFjf0fsZhmybTg+v+AKmQPzhv
kD34k5zIuCVnAHKbXR9gAqmPY0Gpq6w+7DwgngrOqA0TfnsJmWRFHgzBw3SDlFvy
MVT2qQa7E9p2R7RsoIdZAwyLQc6icf5RPd0xqsl5YDM1SBFsx1mlhgqOrtpCbTvL
bv0NQ9wIi/atdwLlltcG/Ztrl6FhJj0zYYA7AgHsgMgYGuIQoOXXLuUID1jO8cA3
gUtQPP2M4sJzQnejBWxp6U8xPf2brEWiLueMeFrgoxoZ2htkmA1RQTMoFrQQBN2I
hgbuzvxPFrHd3oaJg04+VLqNY9VeRI141FiN23B+PRGMkjJug8AtNeRkUKGVLVVb
ULRAawWOjBpBzMhFEN8ljyzP0qdCMLUl1CwMnN9aUDWe21MeCOK0wp39pqlkM+e0
GzQqG+SzPBVa3YK8JZvq7++30WCwQAooooC5HB2RLyEe3xIfOnvnzRL+s/AT3V9i
hiOoWrIWLCjlYaEIFJetzAsydI8gbB6wRE2brAt7y6BfjuQwUc9CZd3yHO9z0YRJ
sJzwHgYqnb6323NsQWiIRU8+z0VHU/PnyBVIgXmOs6cMXN0998W/E0Dz8XiTwcQR
up6tCPO7CnWwNGUazpWaiTOcFeKFZ4f8AOnIu7Wvp9R5qmN4jLrYi2nzIFoDJ1LE
fB2/sIsEYzQmxNP2CTytt0vK9juM10ONe4Y0z/+A47SJiRkwnmxmFWN7utwB+upZ
96CnEqTg1vtOUDhnR6u+YznLyj8IADzc3xCoGBX4umio2fQi9HXRepjODwqXgaCu
vnGjx4yTx37yCz7gO5RFJ2UVOUlPhhD7XACtK80yeRd1NTWdT5bUiMJhNjKyFP9B
FWYSztnNkX1U0UfxEU1jjNxHVRgmGA29g7qlvRAE3TAg55GDe7yGof/tCpyiwjbE
9VX78AP/AMkAzpNJy460exFeuMkAypHS4kKxTIwzKvhlC0yFJXS50crazkIuNCnP
V/3JhHhizW8Mi2C6DIbFYkCbjNgmSf9D7QbC1QeL0B+Qp2jJuv+u61gANrEsJx/l
vQ6pQO+jBHjByeUj2OD3SUNCHLVx/0OEw1Nlv/Z0mScNBmXp2eWfMnu9zkVCLbAJ
TV0Ga6UNz8gTLLy8+8iuGdOBosG2aI8CfGbjLswKpPkUFQ8J3VC5lZY55bBG7fwG
ng699srImRLi3t51IE+Vp5oE/Tl6LRzLedpyminQ6bCPaGk4duEhUZzT7/jPXgtq
9lENO+0wyCJu3FvuSSdudf1PWVKEDhXlydQEopP2FD/OQOAUiRKCT2YGT3rL22tX
x5vA+0nSOhdb4SMUMxVlsPgitE1PVRqlWIbcaTdGT+wHcbgR10xCZDr/x35nKGKY
QChBsB4pWySoItP9WZ4JLa4vaCxDzCReerxNliOB0PtTZlSxMsy3jAnMbe7zF7Ma
b49Z/2ClfkSG+afPsCZ9yyLETb86TazIl76s25HJFmGCznKOSwKecb0MUN0IimNC
v890oEhmyQ1q5od9NDpNw0V7d4iWslcfR6bPqFzJlBPwRrC/x0W7TJ9ELtN5agEY
erBVH3S1fO9wWC9n7Pa5Ripx8KBncjiBN+EFqkQjLUPR9oOYNpyjPqx6qXV5/X6n
rP5b+DlVgxaWk/ha/eZVWS9Y6D3hMkNdw6oQKnWmxw0ckV/ZNUFUoRiw3hFz+F0g
scSv+BwfCkl2lzVGIrfybW1l8qpduRsonw11kVAlpxEu82JJpgyE7ry1UX88rOHM
OOLLskjyXesLKofoNL88vmHFil7ePOcNQkoPZnttDvTxlJOXq5za2DphI5YoMTz+
dHKiOaUsawrAsHWTUlsouAQnV6OgUnLOEzQL/X/Wgzf3W9NLNrgEKOC59s4nXoqw
jAiHXqrIcPAZjxWDepps8aF7NgT/slnWbocPWn7JQjIgMmzC5aH3Ctgy5FgtHa7R
K/KQaVViAqjqBusqzLJPAXjt2IiTaKkNkaFZFf2FkONUxVmA2KHn7URH7b3fNRCD
m9BqzwwTgbF5CysmnmGb7+AuXOycyzWRLEW3ImLgg1b0MZEzXyK5A/GqaNgLqR4O
bG21B+dxFHoLo7A3cIhBxRaFkx7pgvJcpX35mU0AlgcF1SGjJ29S7MHnqrpZV7MM
ZCtoJpZyJsTHMzDS3NZQiDyau3M9c22A6nUNTWPkv2y+Qx5dzliMy1ObzHUe38dq
A0hF5GxpBz8mPVHOYfW7S48s63A5V4au5PfHZYdoDyyq7VWpT6XE8bxe3sPNcHbc
fumw/vTcfIB8iF1V2kHD9eKQdnUmzeqtTDOJHaioXFaf2mNFX7feh5H9vm3hKs+K
OLAeidIMSot0THDd/KKYkAK0HuAwLMVh4A6IWIcNU0ivNVlrKbjuY1BO+ExFmGjg
tAqXbZ99RMudzUc6+sG05UVP2dwnmOR12KVZHEgqUtFhQef3wIEgucbVcFjaSKaQ
ij21PAgYZ93cyGXmh6tOwaI5cShx7HJ+D4WpeAQiVpCiFGT7kYoSvhK7ULsMIqrq
u5W6pysXrWyhwbDoObO102ZcXWum8Oc3+treXzQs9BZxP3doo73Jxp+EQPAthQRb
md0lk3b21C5p40eiSoNqyyHKXVcq6NsKU9LzYUPLKp7VO+jmzvyWk9hIm0joHaoU
c4hmF5qSmJ/oyEyWBwXrrICh6R7yBGkfUXPLocLKvOeddGHOcGDLBLo5OEiWFLHG
DZhLRvqWjsVyNLqIkn/xGqGm2/qmSuyibIS+JRpMvsPCBWgetM+PwsfyPUwtlLWM
3FVua7OqNoWdFZYvkR8+ZYBeGARVc9PQGjPcMX1JYNe4KWxUTVA97tXKTz9x9hRu
PfILvx2stQ0V2ttRT9EAcF0iipcBWDOPKBtb8x0UMub934XHNZldmoXD/Rvaa3dB
DsR23M4vta56EH+rL0jKxIbsqLxkfIv6VXZlPya3feuH4pPpJa9MO7R52LOfIVP7
TbObzzeUyqyYViaOMv3ZXsxMnLLi24pYRhTZgPfPDEd9a/xvLzXpdbxbgaJCCLLY
o2VPhpfX579V4q2QNdt6Y6IteuAumT6XFyXx253ZaGFk7I6QiGdJ6TC0VA909fkT
mMWJA+H+94ATsRPWh3XOPW/dqaenDDCyQvax/Av1oI8c9wb2S6nT2c7iXZzTtUiF
cPg1k3BttH9CV7aI4ykVuO03b3jbGgQACOg/1HOG+59NSlcVvE33IEfY4+gKGs7M
qKFpivguppJEJIJgRthtjwzVZZxHT5KwrBbGp811sQ+JzzxRmqYKZA8dZzS2/a1M
XDJZJ8GlzuazNx0kzo6q97ph+IQF7zxQm6CSAYhgANaDx6OEtW0QvVpu1VT6apWm
jQD0QqOTylt64wiu64V3ub6sYfDzWK/hdzkP+iHf2Oj9CdfTTiSUQIRM+VxpPjvN
Y2LJgQtB4H5dtyJhNedHCCl5YFkrUqoXbJ2nWVKIJb430sYH5s1wuvkuIRiPbNWi
XQcgzp4GnEXxfT/wWOq3A8ellwO2fzyzwdNywzNSQ4gCKP1mMsxNtGJiqXydTKrO
8h/DunBVjn8+VBy0Hxtf0y+M+l6f13s+oCDVJg66XFzMzgnjc1UfBK7EyjSCU7Xq
T2eOHQXeFMUP9upMD1sIqAOMMkM5pTES+v9Wjt+hrD9fsJq8i14cCK+CsSFhROfd
42CuxnCSz9MDMleYd+DdgXltR0KsitQvm+XNoO8+cvkc0JsZrtbKNcBNa1ObRKPd
/HoJOTGHNVzfK/xfiWD9zxHkzlwtyDJ12PigdRmLhb6ixx6yDm2o2BPCl5IgkgJ1
oP7DEoiK0/O6pJ0YxQwqljRo7zxNZMZnHP9QjmwAj0iYj77giK6CMPw6zCqvSCXT
ul5iVXgssi0CAOAwfTjI00UL5dP7RzQNTPKB3lyl3GeIgQL7/RdUknGPahXV+aFp
31vpwWIKP6rvgkXVsX6M8xZi/Cuq3Idk2JnDG7llpUqzh7QRCBs36nD9pA1wXcmy
rTs8fSRxUa1EPNXNJrw21RCoL7B0EXmNTN0g6gyTmg+cYMwM6BL51bTUChAKsbgQ
7GKfDfCeOMrx14CWuU5uwESKCaK9B4yi8Wfo7CBv0L2KEZiVdKZ/EsbHcCI/sV0i
UGfTVpPztYGcMEIZsXcOXxUVfGSk47H+urgYluovIRXvUY9e1MEuVdg63B4lA00y
GJthynntz0jHQg2jjJHtd5HyZG6TsQVqOwR0M0LcFB5SdZ/yYFJf3eNXVCduB0sj
TsCcqySHdZpkyUr3R2d8jF+PvF9fhmg+82fIiHoIFBR2Fo9L4QQlqGG5N4LLz5lB
+rV48EUHU0fjvydgYqY0eCHNZXrP0AtlrgEV8OjbQOTbLPFcM24Ui5QmbGlB3VGX
zKgyCGQFjoSNILLdTEPo4zgQ9DX5pe00Z5WsphoulOgfJyaNzjwVOijsV1250JY+
GxMEm7ueqzDPL+9MRDlGE8IluMSdlqpKMBQGhUAgKAAgw3DPILt0B25Nj8dKFkyh
kLRCu9DMNCflskXjs/fk83nDT4Ey86Ei5qjJUMM8ITyuzGGJTz5llYlcdRwQ2e7d
Y4Jj0QbE7gPVDUdQHYkPCM378a+kvNfYEZW2wiWmx5CdGl1ZpO5YxHUfJZGl0Nq3
1BIA7qjzfDr/VduWRPWDI8Cqoi0ghYhwtnfqQdOLzqobQKgxMabz37fL5JJsKxcx
u84SnyZWJYJSnSwPP2nwLLOWgMBDowtYTkWzBlzt3xjSCAd+hkLDABP6s+usr7PX
bBlISsiN7HYk+yFDLCuWjfw6U0ehpQiUsh8grr/oYR2iom+6N+EVhtC47vqTu/ne
7I6SZr+vuakG2oTF2qE9lPDhQVkl4yXjfvXRB++Kktdhpy7GcHdzwwHWbN+ZpAVE
CN7pRophypt+q2zfht3QkxSZU9D2gDezZgZvaTqfDVliZyoL31l84qZgyG3xSveE
wzcqHANSuNeLxqNIb2hec6k58wQ3V6VyxbKq7uT1BRGa4LpmGbSOLgSfCe7nR28J
anRsIbCN0LDVc+3W5yKROLnszripDSPDqbuT/VxK3GrNrj1zrDaawHfTVn0ewmZo
AADs8fRUYsXYTaV7/knnmHMHkQV5qrEGqLrEoG3iTker7E3aRbl2FbovhZ0FDIpW
EMab2LoAEi6R4RTg6kb8BTqJnlzNGzVpAYP7852jUXwiByUALgdpdr8VaSE20tBJ
FxW4VkNwWaAl1njGZ5gEUvrDNQerE26JHJEmUKyPG+bSB4cDMLDC3skd1jPbHEjg
iiPm6drakLSVCcMC/mLwaswDNxlpvP55NP22u7wSAnoI2cULft+mLb2zw49FcDr4
kBAz2zNXD83P66ZNpeAeGjAIL6MdT4X5vBvgSp33O6pI4N82G6zf83Yi6ge0sBXE
UblpN5xlMg+XXemk3aBqfFTbqX26o5f3ONzUna6skGwYGHL5gBUDOKuwCEwbOOQY
Mir03yImUefD6i9DX6xvgYkuNjHg9dOvmumE5djrUBwCc57QW9Qbyy/luAXDTfcS
l0wPntOhwgNK58bUP+P3NtucpBPOzAGvAquFatop+0rjgAYpo8QCSsZnW5JYJWpc
j150/DN7uBxV+1OYCav0CjBufoJxmO94LGvOu/enoF7Mv+FQWDYedRO7stgiDrtB
oEmSK6vBhi70bTwu2zjem7njhMvXiLCXmoLLD24CsWYsG7rCjWt2pXBRPBtcSm+T
quAt4w7YelQjSFfAE1IRQl9XD9FX+dAR1yiPp3hq1RFK0twl0Le8Kablrwi59D+c
ArIFsIcQTIMfbsnDg92nBNITPioGn77mrpd5Mys22NWLd5rkxCys3sa0jkL6Ptwa
VkKtzF9B8SVWJulm0N2RO1aIpddeEWypZAyOrENb6Agge5qlK7S/Nys6LCR9KGoP
WXv9PQ7gHgtYHybvIx3wP5QfMDIkVSK2JtaDpNNwD5GYtI/NQ8iI10MT7JAuID8g
rLaAfLlJDLY6RDuTeVWjRST9VZZuduhI1kveCBNfrpI4ZtGf/fEc1LRmzYDxjgV7
AqpJUe3AZKr9pAkbmbGnHIjC/UtKMm3bPcNbe/Tb9OgRvbDnNm9aZ3gybFmpUuCA
RFxqhGMpVw1ZGXcyvg5IWw9/q2vg7s4X8sp6tBaELIcNizIhoELFQdSH+m5FjsE9
r/0tFocTuca+D5jAznCAqLsojvQXHskLmcvjkyPCkG19Pdd1xkjj7xh1HpF0EUow
FB0u/7YrYG2er+c6fRhKQSYnmhM7FMq0PE5j1yVKMay/sUc9w3SureP81BelPKPx
c1J2sg9RNK0rT8nKgNhbIPT7XeM0sVVVsbm64vd1D3tvFxM6pSt0je+UwSzrPN/t
iBbDE3w1eL3eltlizMJkRksxgrDRTFY1fPpLOjj016AzLcKj7C16xY7LXVrSBbgG
eVcBr1h9vhSkKt4n9yVKE9yOnbu5v207xnK1nHTOkUf0Vgvn5XiGUGPTOOuNoWGa
Mi++ubxV93X+31XB2KfP098P9vAOhbjTwwNdcvI848WeT3LkeguFiMqlS1EqKVoS
iQJ6BD8W2noee9dFA1rLolVrcHiURIkLtU++jJ47gNuGpDfp8pCgkXlbPLAybXsr
16IvZnQi6AoNcYJZTD3/yrVIGKaVuXaU6PUcRTsOB8mpkLymeCxBLE3mW8Dvo6mI
sOTmnggEEdXQfeuUCSaZQzJ2NDZ4Az4TnDsZPG52k4PkMEm6p0HCWigo5l5ukzv7
lEgsC7k/h4GR8Tar22P09fIp+TgO+p85orlxFyyJf/9g4Dfxesmrc5lfigChKebi
zwOFnzfvZkuXPgrEV/tQ/j0O6Sj3mTTProcLZzc+Aud0PaaLfy1YasdDFrtyS1h8
PrFEAurvS5Gb+1pmBZR0nYoxor2LUYz7ztpaLxxM27iWJDBkKbbemVdmcgx3Ul/b
JHFQkV0qZCXZVEUjPNrEtvXipMob09q6R+qSivmjck2DOzbIw36ZfCdMB8dIW9/y
pDuru9i3G1h7KT7bAnXFj/6Wtyo7KORqxTNx1D6Zyh5fVXWyBH1NGdPvNMF9oal7
Rrv+0xRygAMxicjXn8pNBKg6BsyXXENPDe1V/qZuqjpGrZ/CjLbrTVCW33YsRIjK
/kw546QVAtCTMwvVjcv2ue5GsFor8xhMAU9xU02D96Rcp+HNy1NXySdU0S05fqxA
EG9zHTSxCcHhQ/Bj1k2NucCz+LcoJ2xBHhfJcwPx8p9e73ddSwEhXXBNgY3WKNQX
kbpfoyU01ifSCW1G/5dUZeKh0QpOr0npUOVMTG+9g5MzmVIolDXL6DVAHgzU6u58
sDiHNcBsNrSR5ISt+r6xGxF57TEoeKVwqgwukX8rZGzvUV06/Oy4O1WcGQcOICCW
6fWlDN9cP60RjRcz0uvm62KIC1IdFH1hz3yrrmT91rJ1nXZj70fdQqQUDnjpGjQy
ea3xtKTFgUzt1/YvNqPuktP9xEQjj8NX4kwEHnuX3lsQrEvmevlHppFSmnQFJIHr
rI5gZu3RAIEpISXPGnXe1QdT/itilMp15i/rBtdAOj2Fo04XSObZgyUlGevqWU5d
GKR6KICVQ39xd6u0pbVl6VcO5X5YmkCf97NP+MR27Ho8sTyRIH9mJaD9+4u7aZqL
YU6hkPx3Kgzrj3oEteDC4sjTV80dNiWbI/1OLzFKNDE1AxW9a3AgH78mVAKE3ncy
a0KZkTLPDyPEhwLw2m0j3C6zJg5PfyCYdfC0jtptGLmrqE2hYIuxTZ+hEdo/T98M
GemtuIJX/yVyhCsNo11QYGn9U9U2bykzvztR+jrbFK2F4I7DheGZxFLdxwsKodYm
Ko82jGXmf/L7K7Z98Mmo11ePDmpWb6bMSSrUmR22ZjB8KIsp7AAWKBvAZUcirXua
DWXv04edVujhD5QxF4vrFVMpTJ0yl3X3f1vzTTcsa/Fysd7yjoR7ooxWEZyLCnCB
O5HAUum2z7iSm0vLimBhJ0WLaBb9qWd8CD+89znAUQyzcOYt+InTt7gk8NQltTpd
Ovu6qdCbnXkID+f72cSqH7dy6HNhnTBPzoom8+LktpXESOeunXzFYPo0rakqdK3y
AHu3A5s71UAm7RO++iJqvxYyITfFmE+EckWnY+8irGx+75AtHPzUnAwV39cRiOfC
PsFodOBy59VyWDt3GUWw41kwCTGe8sFtBUYzsbU3Vp4ssOcdpkvwWnEZtIct0qub
Z1bux58W2qhcGiL3zd+SurinPHXeOT9Z7EJKGzP+IOR49d9t9Q3a99tjEku+Zxtn
55pVaLhrX75P/4C9U9D0GrAoga+ReBLgBh/FmrGm57DbRL7e4zxg+k7SaQLmOSCC
iG1fnp08Ao4bnbhibfP/+4Sw4Mbb8qlsWV65C49VAlJiO2pWr4FVkoiyAvpdeQhl
f0MYVwga1xkF7Neld2r9pzlITPrnK5WTCgzUmTr60zhpB9Xz1y6tbun9x5lttjTT
64kGtp2vmVmmXHRCxGUQjComoNfP/CcR5/bxEql2U+zmBzpgHNTEgqhynV6L/N91
kbukp6Li1jm4792Y1KIzX9/3Nqf/nhnPKHtMQ9V5A8GLew09kvaBgHYneQGJhQAe
Bp8BT/tld626tsW7WnErFkmsD3CB8bftDwTYSNL10iw22Wg/RKqrWqDHiLdNpqU5
wiSOCjGlwow0knSN+AdKohbv8taerzR8LtqQyQYzQHTV9mc/PiJhHoe7XNAA7E+W
YJW/HS2XAyRRIGLVLGoR3u3AQOHjttTBLc8IVSRjC8R7Ap2wmjp2+P9v4Dn7PAmQ
oxkGk5JKR4E1F0M7pO64g4TnaI3PISQVou/znzW71AzRb0G5Ity6lkjxUrZR61bv
uESJlMqQqpnL2y3laxUDSZPOf7CJEL9exvf+aZ4I9o2j3R+W53TVCD1cGDlkgSRt
WMi6s7f/BeXg9+LKPaV3FHGPMksMFINd+CCrM3J1pxAJ84u1FiPpotpmsrDh6VZg
KgKFukvqX4MnkbezeldbOv+mycm7ssrqDFPumjtaePS0vbGNjBkRxMTLW+WMr1Ln
Z+2xu8kwEAe2SAc8AyPf7w4nAHHCv85hLdfo64ljA842FFvi06akXROf0ifYvdf6
mdwk0XWwy8Is4wNnpSinI/39FxurND9SFm48vlymOL7mS12lPsdwAZK0jzUB8q5G
VE3eX4wikWQq1ebom1fGq29gYm01ALq2VQcvpyKq6xJ87kUZ7gaqoqkrum4+e17P
jUChXKKSTgqqLlroLUHh7j/wFDjxMLgR3Eam9oGkTUkWMfSIU/4SXrh096DvzuRy
mW5gtMl3tJnP6sb9Kdpan7lboOMHNEIyCDQX0xZSH/wjTuYIL7edBzgT7TIn0CoJ
wud8s7F6rtT+0gaLttmhVwqgB2M6RvqiCgOB4F24/j07EwwgtXQKHiIRM53sa46S
mAguuhsKU4nt2ADPZcAXeY3GAqkwmT3a2jC+WQCFg7Jf9AlCLtt1jbz7aUDnjOoC
2Hj8WqsFqrEGLiZi9KKw4P1mTd6hG+X1ipUBDEA2PkLSKGz5q1Ov/G+Fy1b4ryqi
0E/dRow7V0d7jIlzO9fasM0D5bfCEBC4gPxgW8zqukmKLGHnMtMXiS3c58mKEfz5
DFlZ06q6LpbxYKLPABzh9j1sS9dcwx8y81Mo1CHRQk9QsxodWmXjtiMW2PUi137h
/sZxLMZptZ3Ag3L4MJUHlbpsonnielhJjxJ5xg2Zt3Six2ihXxK5Dbc4weEk7K/T
QyeZi7rvvnSxDZ2sfqdN9pps3plcI49t/DFsg9CQshVLdFpy3fZVlaBCtOHgKZDG
FWcm75pzm8yQIb4Z6XmMyByKS/83IojgmuPSnGhaWPjKIQq0C8KMUQOVFs0tqd5v
CbQN8noE8QunpzJyYWO/too2gVB863AuL1rf7f0zKDRh8mxakaTZwfGYZeKT1OVp
9KjAU3vTgVKe4QKRKNgs0T/mjG82MLNdk6pMPx0nvJ7nuSjyCdXivPqBZE08rmrF
DwjM7rQr61ERmiet7JoP8oCimpZRFYKdDGwK+s5HEbYrfNOAGryNewK0et8pPCwx
9IGsDKdgbo/lV+cmAtjkskfl/AVi5aH/WxKi73RZvx5StjIrBLTXylCZoaRf8J+i
kNkIlcLodKLMWqX5oso4IJ4+mRPSjZ/pHUAI7wZV0e4pqPVCVtHl6AA9iB4zik/t
gsldy0Y+mD/lV8ejucZ+dLN1YY9VmvSRDdZWux2kn/gkB49r3FcH1OmFpy7Ag9mT
W4kpkwV1h4Y+5P1Cfg/5nMYm6on5/Avl8d+GennegpmoAUimW73qkMIx43UHwScM
0AaAgtNgH2nVSinMEmIbZTzq1u7ax3qxm5upG6FsqcwurLKJE0phSbLtHwJ8BnfO
eGsJa+9T8wm1KzmTffzaEqtRo9reSYVZqgt0j06mTp9GGjjDnWNMCLpxcy1NFo1A
mh2NRciAPReiSIoKeR08MsZ6pWw/9d4irkVa91qxm1c+g5L7Vx+j/Ts6zRLdM49p
vLHg1k4p6C5IMZL+wcgSlmYb31zY2gr6b778corBzKvruDfnaA8nXQVQS4b+doMV
VGTHPUTPeUCYzR62JlWSZ3xHDjYS5EzKIjxzdczxXLqXxhnJQph2yP2jvEQOaRcJ
kVV6BINpE4ts/SB6lHCuJYLNnlNG8KoplrvazcUkCmMqkb0wsGIzjjjefmDS8L31
G2s7A19q9s5paZXJRUv+j2LMWTFfcndyGdOp7UP66XERKcIy8YVSIGJb6et4HTH6
A//Ulv6wRAuxv9dVv6MqIhefTRpiV0Wue+Joq2HP/WhS7qHy8TpHeRNd9bn0UjSA
p7gGPc4O7CZYq7Qt6TiElavxoHPOKTRDQTFngv3sJ8VekR33tWWtpeV8YDXuFYg4
qIV3qQD7YZwVmIVBhe3vZW3LQQYVrcsMiE6W4f2N4X5+Zzw7h5w+vq8F5nqyaoWM
pG7j+J3/PwjcJ+zNSMjkfpz0U3JkBYcIOwu/oAN+pNS4yZMWbGximfkQhho/xzJ7
M9OGbPsIVB46M7ZntjTv2cGAD07v4XYkGW/VxiS017PYpZ79GCbok1M/Ml+lm8++
HXh1Pgp+lhdWJYxO+8CAs02clS39RBF8E2LOsf22eED131V/Lk+L68wgxvH/dU0v
l/uoWE5jkVp8tpRYO+vTZl9bc57F5XjUDarOvcuUXP5Pq9CL8F0oU/GPFT6rGnBT
26n1F2IZ1W+6d5i7K0O4v4iT/p7td1a4a8xd4UqBlYOV7nUKSJJZ/LSS1k11AWDd
ayz5M2MV6fYJdE8Hd/Cg1Z8a08+s6XZZdPsv6XAGs+Y4qIDRYtaO4KJc0goETRS6
bbK5Wp/zUPqRNl0+aBpCnNOk0UjQ4WFovCFFOTxs0Z3T6sOGaz6oSkVx/jXXXyjU
mDqqclLR5/rJdmxmxswpgvwn+GAqD0JNOoGnVM+qP/QVc7LYyR4vSogsnT1PrVhh
FUpbxsS57FoVMCG4E8xvQYB8m0Y/6dKrvZxIaz7GMuwDApxP+zE2CBf+TXrYu2Wc
iXQ1pYjBMVXyAmsmwZVOzVYgn9PtRV7XlCdV1WT3kDEX3Y9hiTf9DoVOzkbLGHh9
KefKV2B8D4m16TL9daaidAsELBJFDb6oea26KqfILg9FbzBS7uqTLDWDsyl2Nvxe
IhDPXJnxvcmjFYoYDuwKRj2wfNktJ5abZjULUgBYaVtzgJ/qRDZT7eY11lpFI3t1
kVCt2hZZhP5MWjZjmgPjEIPYGc6UGnLgB2mEcGWr9C3SduXnaf4UdVTe73H//R+U
OzlCZohVZI7PEU5GZPZJ7TSmcnQ2QVgxlgvgtGdyQ2lqRFiJE5mQUUuHUfxdVVUo
Z16Z52+Yxc8UD5n91bj/7qeHHjI18jHk5L8kNZOOZA0UHro1cyh+Jo8LG0fcpWbX
XElR+BTq7HMWQDSTdzRVHKmU8QXQQdKB4U8UZ7ocLP0LM0Z6oUzyWpil8Hpvadk+
XQ2MZhbgZoxMZVlGA5jqfEyVUSllo0ArwqGh9Bue6x26cEi89sE1PZ0wGJw412W9
Z9Vn3YEk1GaLTg996psHkPiAPAmJ6576OWCjo2qise8sqAthHMwz8SrVj/VAp5XI
q3maHxDPfE9DK3nDJORIOz4AidK7HpYLzn8u1gDzZK6VdoTwnFFIAk9jit3OCrKf
mvzXp/RPeKKV5kPpkjpafIJGmo2cwlZULUUAIEGPB6c/ipRQEhk5bo3JldgjZvjf
rtUipfSnXtnYrg6xIiBwAJHxml6vfJbo2JWhG4nLiiabOev3mRKMshEXCRbexBrA
wddAenyuALp21YyflWyGhVe/dm47Eqi2JO4c9z6jTuJpjf5S96WgYRKVijzzcJU4
Yl5hQ8ULw6rLprWkpfQuBn2yDo4mI01nVBq7sxJeNoZn+OJRh0GZoBL6aQnfE7kH
73d7dY4birZbgdD3GTRRa90CJpCBinTAGq1g9xTZ4byEF5VxLjWql1fBXRK8khEg
/DcXxSM0VnzSwg0HyosTamNSQMZKAERbu9Zb7Pg2Vvpojxjpfl+OQSZEbyUysCSr
zcCfpT2LYskEOj26QC6SruXW8lbOz3ynsdBdNQ5+019z8RYpDYdWTwGfdaR5jAxX
YJg33mFl465S1SaliCdkhLpTlSmfgxkN9nuoJIu4N0VDgba88mwoJmQfZVMZdBLA
rjzJZKo9QaeydDoGCTxME8fW4XRg2BjpP6iQa8eOTE18qW4p765eyK1tnHEMYfZ1
7AmkCGOfs5sRpmKn9rujUYSEvbGH1//rp8sroTWxrto3Res7UtCS4RRlAwdkTbJI
nJynceuxl1pKX6rNCGS0rJm/qQHqabDsz6VpaoCaUJX8a779OG2n8A0SI/ooZ0bm
73EerP3GBkPQ4eGju+gruuMYHvleIKJOACua0t1PXwO2eMw8ZOaybYuLvyGL7Hts
nqMKOC1oVPN6rMHZPUpYQ+up1JtUQO2oSY70uqbAE0/IUA4tDLIMM2uyK9M81T/I
EqXGQleXM/voQxM+gtRYesCdnm/u1HIEj+tS95i+LKvqyML2UpHSHhnfIeZe7HGg
jPvnKg+L/Bj/Cil6yCzOEstCo3VCWgzDClGL95Ioflyaocf5VXgR/ogOHa+VXB8e
754zNS8JwiNyb5Ejx973Wls3qLfuJFVtW52utOnrrHW6MTP9KS+Dt50B1Zb9uM4u
bD4Bjf1H95nuiPvd2OiVb0jMPAh250qXNhoVfeVBxin/xFgkO63ZTT/BaiS7dmZH
BMDsDcKpXJFj2gReBHLZ7Jj/6KrToCKz27ReGVpRfBsEqseO/+7fB/2S5VBTk3vx
AYPheKz5LdBignNA5s2kdIUpkCJJ0ypEnPAv3c/IyaK2z3jDXY2IMAoRu2V3NneJ
HkG7/fRu0f3jTXImlcpindmqyRdk/TUgSJg9rfwKwnwVnmscK1dXHnh3EYM5KQjA
n7OVoYI/fzZQIUaXlJrBJ2aM/6hDajV18F9iL6/CDF0OaPDtQ2lLSpBo4VD6lIGR
2zlTzc+erG/1aRZc1IWEnvSxoH8m+16KmDIjDnlGpS/QEZ65mYZPs2q4dI3EUNqq
CxYI28BeqGjdev6/PbFtmQFpBlH4DeMwT62rPC9AYXGzKnhuCSMr5PUk43q/bJG2
9aduDg1986gWUdZY6a7Uvn46PJicnIkvEZLTW13iCdeBkcCbhuGcgy3QoL89xtd8
kXr3eMzfpo1Ne5u0RiNmM6hZn5M9ydfcgGbmvdxvt5V37VgkDTjek5Dk+ARtIJMo
Mo21MFXRQYRKHR9Issur1gxuk5Ko1r/4z6tWEG2bkG0h6K5vwmZZWJ6isI0eAMVB
mEMAnLSANchp3cpMABjxS1AhRogx5G6q9D6Q4h3NNZjjtaP0GPPngyOB7KlKsA8M
QgKIrsrQhSdcZ26W+qVnqYMAEoC9S2EZ21N00G/E0zx6nxJOTAsJCJ3+CKvVh9pN
iopoPjzxyPFp7e4EtbwZ7Qdahm32cFbay70KUtbTjiVqloxdwLsp6pnCrErllnZf
tdGDHjdyNLaWgPnhdHQuVPFfqbI/iV09DqXS8anCe9XfsCOBPd5wZBOPuaZR92NL
css7tOCSuO9b+ynHS38Pwxca1hRstk8J4d+pKZcdpOF4itxon0Tyee/+H52RLLp2
lMWlYyxWeZV6w+fPe4IX0jT2blO9YFuVt+Z3NSXLeLqxRRoyI+430ZTulWYqBAiQ
P8TW5CfHVWJSdV6oME48FLbi1YAz2lRui3N264mURDLM3Mx2ponV2SSkWXRi3LVE
Wqv4t8Wj3S29rDmQ0Kam71VvffVT1zyEGvUYgl/WY+069cckiTg/tAEfftdm7EUT
aDsMtZfvBlNz/JvXrkiJgCaxtgL2Wcu6tB0LX4itM9DA6s1KYGlRiRDnVKdNgUpP
wyH1B6dTcyZxPxtRMfkn0LjJKHJii0Jf2XvORy2NPoJX9VsQv087if95fCMKQjGn
YrnnAAClNO0u4+PKAR98HJ5znGh2omm4htrBtYW2bXi0Qi8/xzeJ58ABxe2uR3l8
fRiK14NpaDGGhLe6uLNHEbHSh0ZijXBk2sMa1xmOum/AR/cznZyQiUrZfj/RTQ6S
FhTFL8s+dkDwDf11uTLB9+WUU+5kzwHr621DzzY2xxWq/fXdsTtyjPkfK/1mrzG2
btC6ZhdYQRE1N8dMbKi08Luwhpob/Eo6f5u2puV+8i3/mhgVoVa/RQOk1NYtc5wA
r2WEsUM41ERFDjEihmyf+TrWENFkfVIU/G7FTgkfrZvJv9O1R0RYd9dUTBKJC6Za
gmWkXozUV2Wfw3Xmt91CDj8D7FukBZ4l34+pjqBP8Dn47w1X/tp9NyIiIwrocr8m
4iVWekf12GpU7dBOzw9TeicYbJp+KVjOF+nr1vH1vDxf4wzBE5oxS01nzGtfZitP
Wnh8bDxHWzWcHT/JrqRedpqaFPQXdksocd3uuQa1I39fhZfczsZHEyH1avC2rIWY
9YwweklbHcMHLj1gI4p1SFcvF1OJ+ljWF0x21hmHRcIEhlVd1dJJqjKHf5mAISl+
yn3HlujeTVJttiYNyFhj90QkaY0eHct1sgvS0LVmP0HT99ajAfOlRaxH7XwEF5Cu
jUNX6nZTIl2Cf9sjjfg+ZTSGcn6jKlnUO4owy97KQ8FZ/zIDaMkXzdrRY6Q4uj0Q
Tg9Mc86pRrsTHGEHkySEsCWnLX2gpcsKbWb/XuGGDpILDFJF8ZwLq7CN0v0F750i
VIllt55rkMBufOG+H5RaW+Upn0LTOug5U5WmaLP973pDLKVKu1BvxJPqlb79L+np
uhp9R56ZufIZ8T4C8sUsos4pxMeN6lPKxmMmYePpjx6n/AxYcuIpR2MAmjRWhl7u
UWho2H08+OIdC+0vZX4ljt3GTqRG1IRrHR6Tibf841unqBk36w36Vvg1LHzH8sP8
qALIdC0P2mh27CF17X0kojvpZXzRGXUoOsbnv6fpL4hGn4YFd+mc37jcIsXc9tbM
a+yB8vnSC3I8i6YwExHVurpccmK3JaUxEC51r8JY4jdL3/zMT0EmkH8ks0R36sr7
WoqS4nIGfBEBpXz0kZNX6hjBv14H/ydfFsxMC+zpjC/O4DMoukXYKUtyLTeknlCZ
QEwQfTO/ZoNf7uSSQH/zmYVNmR34vjn5JP7wvqgMjH4SNzgTRyuy/79Xi0HVdskw
2Gw6pwOI7K2fiGftW0K0CAzxQ7EkocwBVZLMxlHOGBxxWxDdzztiKe6T0Hy/DauY
bE18JY1/jC4BX0tr0gq/CR+dMDB2Xdj5Ke4fV5TAcCnGRYc7gMJGMyMV3nwEiEEI
nlwJHzeIAqh+MwYzDZR8YoUXcpFwjTCPfCaMV1wacSxv7CZk6joerkATOVEKVJcf
TTnD9HRYyGA3+j+iKu2xS1wYEMONx20uTfyp/nuDtBZ/QijnOQ/pZhfrDDywfDJ3
xtsgDMh2fsJAmos+2FsoSRgEyLAU6FvMJG2n6F7ukCeLl8G2cfzovwbSMsLVmFDT
3y4+6Ue2pT9i3i14W48EH51+i+30KUvwPo35cvHPhEUVL7bdZn9qRoHEZjdCz+qT
x4eFaJ9W1Qig75c27cbX9Z95Yyw2PYZeOdeKf9KcbQWfvdD4E5VumXmaSHKIThgK
fTd3pZudeIWhBlODLcsojGkNZZg8dgn1sI9yTl+Z0mVGp0uEffWKxJljyNtO9TLd
5WPZuyi3hw+94CaPyZMR0tq5oiS//Eis5QpSknLJdKuQTtiUILtC3+d2lT6dKPgf
ZvClWlCUrDsK0I8MP2dSahoy53jlcn+PRUzgSLQT2Nlh3QN4n89eQ+UMX7OU55kT
DX1gzWUKtEEvFePywbq9bMY5gn3g8gqqCQH0kGBBNDmXeoQ2+7nEZWiVYoP6Wq5N
UHgxlAwlIzCQ+rlNJIfYyBDgXbIBUl5wYJfEnKqgIX/ARaE1B/zZ5VGWBWzV7ZOv
pRk4c4GQfE8VYN8+OseG1BvQjQehb57g+s1Q881k9dHFRIZZT32mcHVjA6w0LMb1
/46f6miXHF398qM3+fV56/+onqIv91BXS9f2fVZSL/jHRpXjkTGzdDfUSlRvfV0W
UM5swcbaLYZPDuqlSIOChn7JUiGXQk846C02Jm0xNwGP5qvKlR+nSdI6lRsjrlTT
DZ+uX392DEIMKsYqe/80x/EflmkYBORvG9sXCgs0g9UKtb2ppa71CKX5KgzNMWad
hgiH8IKGikrld0JRgtc1pCwIXUb7CXm8UZEcoVzo9pA7+REuPMLC9FI7m/FBHOWm
G/vXjpcW6H1hPxXFQhUbXUTZwHGOjut8P6g1JCjAdi8sQeTWdxsG1B0j8qxNE+17
bGbKgChbBiuOD+RXfKoMhmbSP3GGxEiOi7bzvtY13vamB7rM/yyvTC74dcnStkyU
gkTdP7amvLRaCAoZ06R4yOWzFYB4Y3zHhPa6sRRdwnEw15M/2u6P0iiSgol5ICvw
Oso1oa5GenHbAv10GBqaX5g9Isi6oM0iJXqShYCnpX3DPleY7kt9DMZ0DWBXZIMh
OozVTNTpNsDL8bxe07JFv07FnWML3xh3rkjFdhXdNMH8jUsaaHsNTFzJ2cNKh/br
HbTXEIo+Kve9UcMoU1vAA4eD/5MkJ0vxPaehoSNtddrL9h0VMniqMgtsZpvYVrD1
EkgJ/WpAHzwBJRPh4CZSXwJuzWWF6es9pD5cbd4hL/WWX9ynK9CygC7Fh2+j2q/s
BydoXsupZZZ3sVKmu+P25+lGlKL6RPrpaNv0mrme3AgBJPM+NyzawOEbpFhrRMNm
0VZnpwN3lLcsTpK9WSoD4mXinEi27ps1mSlyrsfpqXZ41p5MFjt1imbSAwf3HdkC
vd2ca7qMHyoFUVXtkhz233CiD5WT/+D4OeP2+ig/B/RRkXiDnsBBu8swBZ/LD11/
nRPdh4jCmiUEEzc+uFjNoyx94h0QR0dI6/pNKkPDQ5l3y1Jk91p7YVf0y67FYK64
gTk7/gyfB5SnZ6/uT1p7dsEMfCZJ5RDv/IZrpoeEn9oY0oa3px8af19LP+TaQTYn
oyYydV8Vut8KM3YJtMsUt1UDGzuSvCczD+8Jy+alPBD1wZuRkFSVOmoRBoYL8tsZ
gfERWGyvVze+G9olyxQk6w3PJKqS+AYcGHYbF5w9JyE2WEZUKqXSGgFk1Qy27Upd
yFt/Hc+WvBoUWZEXc0HWxK+DsyE9LDVNP/vJIPnvfvHcamyh0vh8ocErrxL+06DW
WC97mfob+jwvVEhQSq5MM22+BHGeQZzYWbFwDkCGpKKQbkAkdId5hHFBnS4VoAJ4
nLLt/F3xGzG1MsTzfHvUl0S24Dr/sbA0dfWJM/QamIzkznNxqHFqoHCVA6wR9to4
qL+OMybrhnS/91GlJKgeT39meiLA2SMXZ2PHlNe1pXrIisV4U3WKkfkilFzBXBvp
QDBXbXMeeIx7f0zmY1dTf93+8VCoGrWhbI1yPZ+SyXmBWde980ii2p+DSBxGySiy
E1fRtrhNrX3UZarXV0JdmoZjXGppal/JQhws3XgMUDYwtNozdqBKTRRuPGCGvpX2
uPghn1tHJ5YOls8VN3fhFqPMiWMkX8tucpmE2W/BMf+o+D7SU9TfC9v/DRnKI0FV
1bkJ4uztCxC+EXpNbQGUEpZzBnoCNBSzr5O+bxKIrImC9TNWEkcFtw44gQRW6J3d
XYJGosS2hM7R6+tgXuKqc1kJ+uXO0EZaI3ENvAIBrsywYGZx50muqhehD5Rdu+IP
w4mLVJV/RR2xnWU0bvT2LIjjXU+L2r1e5JC0SeTjEOP0axL9X8UUVh+p4ehVysyN
TlwRpSzDn7tZUsMfyv0SOnX44r2Pt+nrBwD2RYJWJ1K0/En1vmn3WL2TjllB+eX8
1frRXGdvcVSblw8rEI+5D/2NYnrXcSUfMM1UtdJwFVLlJcxPqmvgiMg/kiyJJFDQ
er80r+AG26JijBcSpdxyJCMB0iZkO37aU5DrUCjYxShM7Hlka8IC581d2lNKH3JU
lkaMp0L7muV8u3KyIeSE//tjYinYM80eyBZe6gfclAUFxy+TVdaXy8YnzPf1Zo89
eEA1LO3UDBa0AkkC7d3UqZMMH/3Liqf1I/n0s+UjwibbKv7rQGhzLokAWz3GnrH9
ftZlcI3XVB90EAF3RnS5FzqE1NqvGkmDQnohQufX0cRgXXdvcYI48xAc5p3yl0nZ
ivq8u9KX/CTTuP8hvaBNBg1Yi5lOZouASGcOvZ0r3qsfGKxfgB2+xlD2JnqBXrhI
pCAdvd4Mi5LcVIyi2OaBcUn+ZqWzOLaa14R3ZGIqSdSIdIy42354wdL+dQSjGHbX
pYLBK4h5uCnlUcr202wTslQzRpk7V2LaXw7GMe8ZtMC4R1m1fX5GaAPYRIt/iqlC
OjJsj3BleFY6M+Sf+RTvF3mTbNSUWPphavoaYshzCWZD/HAHMX2nr2H+zuRZ86jL
AWmiqYtps1xOa5Z/mCCMB/JXYemOc0IwKtc06+gjndsuNQg/ithvwFUVfOGwgscy
MotkWy035ESP1CebqB2xGChi9oO2DjKoIW4gkMBMtW37JfiPU2J+b6uExmHrlnYB
+R5DdwCGIISWFUeCWbugT8R0lWPh8yy5YJuOnajqY+DlZnQJ6e9+zoQJP7d8ZrKZ
eidsU3vfYwa6o+OOL/eVDPk2/19Nyv3WIefD4e9sKTFxrUpOeiJPtD7wfGTPC3lS
1tU5R+hd2o6wGA+H/orbdSBk8Ce8PvtFP3FRIhVJn3ikty27LFfj0rDYk8SA0r3r
kVrxzuXyXBeXUukMDccA7sRCiss1nCyA/OXdzNWUg+m7QJDUrs864ekat3AidMW1
DDRcO17j+khl/JY05LSzVjqFGuhx/9eGnZUcQqCWT931u7VTWci6MgYYSEgcEXr2
NJyROLVFagcnvq8T03//TldiWpUKOm2hzYcn2uJ8xFXv2IU9eRzaw/pYXUiaaH8h
kjZdpeVxsuKXKkzLsWzn9+9InakIeUvPF5qji7khmVzkjzJc1wuYEh/lMQp/n0mf
Fd9JZBAFO+pKI6Ye813JU6SAV2WOOi94UceA6gYLfhVok9xjGv+vYV3D6Gd8cMdB
lQAcDPdK9Ho9ymQsek6mIqi4C+GP5W1sY2gqTJ+coj0JTwa7KAYpS+2gRD60+VSW
XYgDwtVPII6y72vjmFqRhzDee+tlUr6mrFyjE2Wgq0bb0S+pz8uJpeJ+XaDNDLe9
X19f6LolAMPg3sBsFSTo8akwSX3M9Hg2c93dAVwmx7aab2K5jt3oekD6FzeuUB3k
WWcpWCIi9HY2gVYUuBRx2hnZRaJ9j28ouYmDHXba7ts1Py5heNryMhiGKocrZq+6
1NCURYhifxwXLncyYr3BuVYiF8djNARYfOQyKQ0oPYd14pa9xVcYFYBLgjpcKkXt
Z38fudVBK7he7OQZ/nYT0+GjeJ2KJH1cM1fZ6O9AJU501Xw1Y9ZiAQZkjNwTBXYD
ZYq3PBkD1ShSdrj5OZtzGbfUmtY+j3fM1hVZ2sc/ZRdQqE+/O8xsaC3YLXJerM4G
Zq+2xzfUlxAxmLwC4eAbISWSTlRwyf6+Xn6fxAnHvc5LzipH7pq4wgK2v4XL61Mu
NS9WYp9ru215/v4j5RkFoN0mwb6t6KdC1fMIARBW+puDAtsw9MpPVHRrFTDATaSw
2n1tiE/Qbkoh7DP48Nncajw5/P48duxRde78Haety2vlgDBWmWZ2BXPXg0y2poFU
YnN/Pt58lJs+oONXH2Jscb61aabVbIP57Vf2WLzb0gZmortukUp1E2LffQAbQWzV
b+M3zk1d41o3wHQY3LxpCs5M6atQeGY0qYs4lDrjoqKF2+F3hSWcELgXMHrUQn0N
AVtsKkSxf2jVAFaN0UamlU7byc/XSM8eU53uaS5ijf1N2wuctywIzvReZmZWMvWx
fAJ7WEnJ9cPra1Jtartb3OHM6CcNCbafZUg0Gog3d1rEFlxj0ExoQanbNZWwlQ6b
5Q1wdqpWiQZNzFmiWQs7lQ+qSwUe5kEcT+EnMDhXgy347lYEjOAaJ20G1W5fHF6R
RmvKOi/t+JzyKmG7J2xjoID3uLR2wTWSf0y6Ow8P4xFu0RW3EHvoeq2HMyKMHxZO
XbNbBq9mViyQfz/4TXpgKQOiqGYIPsR8Gxi0ig2fX2/NylP4glIv6yL1Da3doa0m
dG9BeFb8Y5UboeTGlTaf7JOQrnZbkYjH8fIu2s66GfFr0Lv4qDBckBmuS2DaZxT0
nuOQaF0ZpirF6OhNaeoom+loc5QkMmsjrui/IIO7PQxVxyCPplWBxz10e0Fgzc7D
kk8IRatpTimHnIySJ+nV5aL2dRmsJrzhD8wBr9DvDL/TFn8NQ6TPVD221+b+GLTH
9DpBoWdKNZLLwaSXkt3MfYDNEMek/bMkSK2HYkgTf5KN8sU0GY17pO88R/etsO9o
jdR7H3qKc7oI09XM1Hkyo/TSXxKdyzlL+modjhu/cOd7zjtl9JMFrh3s5eaS+nIK
LHhDe/5OaPXE6hnf8cESRQ+zCCM4OLwH521A5C8dM9WDLQhEnHqmdDsKbsv1aGkR
PMOEqh67PbFZAGAUZuYQOcRt49Ti0Uqlm+jtwSl2TzzHKREmf7RlG+8k3PUbFa7V
eU2gE6NVMEO3cbCP9M/0JtSPw+Bp/zlfeVrdl8iAyGcFRPRpSEa7CAk1fUVwS7LE
mTJoz4fQsRGLaNvGTYOZEOxm3fdxk1xxrWLbgVpiPgGBib5xAqIytkWVcLBy+EJV
VC8tWlYf0I/f01vLNi2UZSQK/G/cAId44Ff1FtqTO4LY7Ngj7WQiSuWy1t01aLc/
VqtfQw6qZXfeiHiqlKwqp/xxK0MDvk71qCztspFYpAGjLSm8g19mX2AIaBNK9Hlv
vkz3fNDFIjRy123b8M7sZxh/9BpGljNcMfHzn9Ub1QwLiUksyTz830D4uTgssvqN
XD3xZozRbIFE/tY7sF2BBM4w2ahMyXwSnbFieuV+/m77R1MfZRgowtgduJOhMf94
PqMQ5y8Pk1ZeRR5XnTbBbROwxJNGmigoeG0/Z4ZNhg7ykS3rSJ5pr/wg6iLLaBv0
TtQsNgGIEn+oY3J+DsbrPkNSHU4/q8NMpzDMwrMoIIZ6jFaqjZdT7dL38fgzwEMD
wLXHBR34dsO6fOsWS/VzVW9uaZPvG32MK90AFXpuWw1Wr2pIB22sZWtn21bUcYls
zWcISwyz7Wu54oxhleIyWTGDF4WplrNrd7l2lzsRjgvuVjLLJd+n3Ou863XXlDrg
HjO8h6kda+MEFhfwR12uWCKhDZigsDhAhE4/3w5OvZRhFYa6hVBK4G2BlxjKyAJB
h3euno/5MNF0mTmSLT5st05c/XbueflNDSSTSHnPfAf3MPz06P6MLejuOncr/EnW
8MFQxRGraF14Fxz6R8OoQpZFayzL/WWAA/S2hfxi/NOwCpqlRHXJbycCseb1ppL2
gBdJ23z+XKHhn3JiZLBBmGWl7H6jfziRMBDqMJiqF+HHXoMNLdeMOIGAkBUi/lM9
NcB89KygZkKjst47Yl2Plok2cfbaIpgOUMwM6XCoGgVdDmhLJIVk1kGoeqYg9IlJ
1+HalDNDQUEZ+aHKG5nB7DQtCU/B0qM+9T/9+8ySSd+LKPuN3eSIv54eiqZhmXVJ
Y/s5aNfDolbXcyD8omaGmhVVP8W391h+2LgeqJVt7XNPjYEPS8Zmr8uMT15EtzSX
Nyf4GUoEtW9rdpGsvAv2RFumZq4NXYbH7Va8BTn/BgLQMZWZvc36nwqMq5j5GPyG
AodKe7u2v3WaF+P6MhGGqABVCaI2fc+6iqbMD/XZCPsxdkdrFEOZd5K47S8I7scg
erhrLds6ucAZN8/DlS9O/dRgsnt2ytfYrpxaCnPVD9sglXlkOO32w2OBbAcZ/PVI
eU2GbyI5c2Cpuyz4FjslD2KnkAB9bVNz28hDukz3f0/+elNdfMbCPJShDYQ6QX5e
H+7bRT0CDPOPFC4E4ypEN+E34rvrN4zB6K0MJfjeWFvwv/KPYalKxVuaPOv6+tJU
r0wLTsZRLAq8ysKt+1+yQ4/4eGd8XtJZp831p4dKSW51E0dNFWdzYux6mW+FGXgr
+Fe+wyRfglMxjj82wIo2GIL27t/vX0SGZDTanrJmURV4yrNDwIQqfYQgqCszMjHC
WfYX8Ff0qKuKrf7oaFJm0NwXUSYmw/PryWspy1ZqRrU/3p2pnZzx/GVxC3AMv4K5
luMwAfGYzEc1ivlTMTA3PhdtAwx8YRg4f480BvOA2UbnoeYsLYRRQC5pjl9/aDhm
257n4hd+R22niqIuhK6s3A5JBPKEL0Rw6hN/abmPTd5sN72nzymCJmljq8r1Xxfn
/3EeCry2UpwYt0Sxy6j+C8aqOc+It1/1mXUnxDSCNTrgz9gDjWIwNYQYweATYfhq
BsjzJd+THx8xXGj5xYFCDBXEATwTCNbapWrsD5QxKfXF1muXSaPAzjBzHcXpAPWY
AIgRdNnidimI+kp5Bld7vOMcxZjkojCuVao/uju4XQZf4479aDRlIj7Hydxrxuws
ubGC5qY580SC47IHApnLApaYcb4EEmlq75p8kyhCOq1rqkOYzxSSPaR9f9Lk80os
7gKSFgGDgqdeUSEa3XpAcmsuJ+PZJWNnLdWUzIdANPP8O4HJYv3XNZptJe2OPJEM
lCGf3sNIevR1Qe5DE6Ggm36fDDutbEBNotmYSggAA+QikoHwmnn4ygYFio7ZWCx8
wEQa1cvWE1NX/xHluztVkB7jldsDYnVIi8n4JKB9bjFvJtITp6chkmFXo9bGVUih
HrCfP0WpJW/caTT/g3jwKeOvY3zbm6Jib9WsYkhY3XBXnE2DysriXIkrVKyW20+F
e4sNfGPFP8a3vf9RF7iL+W+XMA33Q4KJW2aQ/LWLCrkdPJBJUIdfS1W+bqkabc63
hNT7glewNZqmlqvQbCA4Hepzuletr1Zw5H0kgkAzHkzqk9i9XcSLbqMv2v61YLRm
vHotqN0S0trbznYMvExi822WIR5ycHR4holBmsUO+3I78LUMLbLC79wV7QaX7zu8
JSHqCrC78gLl4LSC80A25l0l+CsAGAdCnpUmCYOdDcvlyfPE/g90tljrrDASFG0i
0NemZLQOha12oIgM67BS7Mygm/fc+5bCaer0YLxJ/m4Y8m3mkc3U2Du70IaahGO+
D7dyxvR7QMvjtdUT0yhNMFEpWzmpMpAzigV93KnJIU3FOmiw1DVpLtSQXzLxLxbK
Wph/J6eim4TrX0C+yMTRwKq6LnrJUqQ4PniYw3Ho2HWs6cEGtNKSZZ1hLk5Me8iH
y56A2lNsC7sElTtdu82Es57ZWB7hYUL7Kp3f8c2Ui2DIomGqKzoHr3E4+E0hiFMp
pZIKPbxOVvF2/ZkXCPWbbVkLH4ZL1uVfDsXHlHcKK2HAhozZa3+dHfnkkMhFUuRj
ZO+mE1cUfq+/jzT2t0uuAe6iH8YzuMdn7bBhiTxkgc/WItodCRoQ5T4FL7SPz7Un
ykg+DID9yOHc9w4qg722ixtGoq7PXwt+1KrbUGARtTvH1YphefZ+Q/35b/KUHgu1
ZZz5i+ywb3zGZT/HRyOrbntRtZVealWEGUGMsqxxJteabqceQLkDJQJF6IZc9SXZ
iulA5DSGQ504JnF5oZxxPuyALMD2OupyVTbllfoAPKeZQaD7L1Jh270YIy5UYRPD
HJNNcP555iPCIo+cf9oPqiOJIEEQstrAaIV+Je1BW8smmsmT/WsGsR0IqSLypPBC
u/7F8x7RH/oc4HpftaBH/9Xty+Dym8s0/fwGG41bX08o33PkV1BT/awdqfForCoX
cMy7BuBUZs4Yawfq8GWTh+zogMi5U9xcBTWkK6rx3/0Flh2gcsU+5BELoHgCa4Iy
/JI6Qr9Rj+94uBQJosQIThKsa6Y9oje765/Jm46RQDMyH6QwdXuUhmXjEoHu2Oyq
s3lyp87gY6/vqGQXC/c8SWxUODZ/A6X3qz8CGal/QxTu6TVtsFQ7ylBVb86KrnMc
VHp0EYO3QHqNwyTwDeDPtRqDYKB9aACkjtBoQ0M2J1H91CPtMe6zYRC3e7Uqh0Jg
iRguM1YRxV5AthAHjyQUHN1xxRGMUPZZqfkJVx5rKaVLE0xUKUgYh8NEdCY/wN6y
vSPWLZ/DyglL/cMGDIceUDPCEhl7RQV8StIimOGX094RsGARbFmZOkvx2Nq6sQ+y
QzviFAp3tEyfUhukeuNdueAj5M1HJndpoLr4EBQkM2PE67xs5oMARpu6msHCbKiu
vv+Rrue5WRXTKmETRIar0fJ9hv15e00XAd0CYIDuCArvtav5U/lKpwH7i3QCJX2N
nwukD6lDO2vi4bphU3VLrGN4YH7hkw6SH2nDMDYJgBfG8I95bTbxVX0eyv77WYrF
KZT1AeFNeyTBGGYYRsyYLZva8oPsY8y16R0G9Ol0TtwZeTMBcwlndEe8z8JrpQ+j
PhhJRPUGX5x03HUzzF6pJ4pObmBHPuqfULS8F7fuoSFa8b7IRaq9a/X57WoArnzn
2SPK+bDSnQREfJdFsCL7VQLd6fcMG9HiYt3auO2bItY5utZ/1/u9gKDkG0FtcsiU
vHyc8Eyb4FvNjBNqYdpNcMunXtT8ACd25FCLN63dygU=
`pragma protect end_protected
