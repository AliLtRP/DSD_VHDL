// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HmuNgIZNcII8AhSUV01teM1OtmJpAxCHjPWG4LnYeMNSO2ckGrWvu/X4UVqC2AC+
jt2KNwcjj6Fwu3el/BWNjhCBXhsmI7kIdPU2oA+xHott1QwZB/8Of/LK+Qbvvbpo
jZLnSqdASssci3PjhMpzQII52DD19bFrKqv3MUsPLL0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3392)
mNqHebeb9FkzuLzF0JV/17B9vViUsFASzK7rGHIBOZH5TlDnXoK2y2tYSr1ajz7k
76oYUysBly4kmL6/MmoUabWsWmw7y/EyYgQudnbGhiu97NrUn7I9W6ivEPecZeu0
BpQJjjM2uUOSm78aFAS9SjjTA/FYRs4voaUvNkQn5rKSEAO8RuTeyPvRP9waME3/
ML42KGU3KWIBDou4WO3AaWaSAuefxiq7zxPGVLD3XhfNS/8VawCfQ8rKB3i8JFX5
UOCkJ2/TEKiKYAAYf1g4EIeNzJh+SHfS+hUSU4YUc4AW5D3dHKR21ZoFR0FoVtn0
jxXwUVRK4hEhrvdgmC6RO0qAvatJkwHPjjrrc2xLLiOTgQoH+vNVKXWMxCJ1ik3W
CWNngNkootoUHVhttOoqVDjAZDhUaNGnFSyMAwPC8YW7ny5W/FDy4ZY/ZZHgzIkh
Zde47z/iLJoKxYL+WrOXslDEyiNwDvOLgDl0Mu8GAq5pQmH14iLFDkWPF9cgZnLb
yPG0E1KPHqwJD9cI/PjxlitTOo6+DuI2AQYhDFMJozr0mcjYj1oUahB85jgwhN8g
ohfmhR0dnEEh2gjDrhpqao6b1B8Y0DIntKpxFbaw3LaDaLLw/8OPPNilrrvl9vFq
gzazLpWzKatkFdbIYJCm7Yjrka/iCETGuBZ2kNFLRojcjd6uxFRSrE8/KxwuP9q6
bGUMZl40wi7whvf1m9hPmr52eya2ShFLwo6bdgmur7Z5XEA8xwEyx6GX+OmnUIP6
6bMnAtTEbPwtGEjaX86LOTX0ooPhBlhcOCl15eUXFVODPeofcuuRsMFtFXFoIBJU
1edZ+nonoeDbOpgEr21j4ro+jIKCIiMDG1X1KVfQyXQB50/zft9gh2Ss8wLDYBf6
uHLe+PvB4lgZK5rBDWj2qyP0ai31IeO4s4HBfxzF3FHtreP6p68CBO8f9lCBobMw
prcYxEF/OkSvbf4bNn/g0T4D1csDpUbCx/UTWEQH4pvGfCd+lPfp0NUb/aATv4JX
Fo5iUsyGQHwnat4x8InI/T86l9RN++RblscFSg9/BbNB+oGxF4yEymITwJ19LAGR
HXltaeBzth1xzD6FH5rDsPsko7BKMhgl5AA9sR7H3PWEzQ8M/fX2v/JcfjBk4ilV
QHQjGZe2hqis5iw00YElF48GKt0M2i728DBkfkegV/1bs0WxkGeHEatewZSmWWqy
aZdMgoUweAEmgm007U5CMemwWdnLuEkn41Fiy1zoroamB4kyXIHmFbYfVH9ZhKcn
e/j0Sv3SXbQhxiTz9dRHtUBraIu3hrCMsafhcsaIu9bT0I5mPsjPP/X1Rreuqzj0
bL4sc0pm5nL1KO0OmpnYjv7gZHcSMJq+xbYYZL0kUO9V+nun8vLC+Q50iXkxDn4+
aV93+4f1QYXkJeQcD9TwVB73i8k+tzoocyuzCmTpMg/svUYhrPKbHd+SLtAU9wLi
ZVr5agUpo6RjrKRRK8QzjVBxDXf6iY/oVpyuCnjcqL6tA3aPH+9Q4haBwVJWPqZ3
FZLI9PIP81cFev37Kvx8QrMh6yB84vdtdPlrOEtEZlEs3uUJAC0soTN3yTipuUbn
CSt1lp/36afehOxcAVDVcNEjG94NXhIUGPCsRE1U3TwkSyv/XlrAf1c1paDZXKKF
Sw1Aed+xBlSJrdW9wJJj0c9YbWvUN/vI7fIHF7cEY0nxTOsjAe/YAGBUaT33LVx1
HWzUARIGipiPfSbuqRjSENuyA3ebGdjm+LmTBZciOF864XCp5NNkaVVxnngdVH4I
O2YqQw0tPbVC1dUNJ8Qceb1CKsFo4r0Bl2Al1t40AuQ+9SfCkZmieSE6Um90Qrmy
ZjTfslFHjNQMibpjinpO3VsuSFuIiykFrFcV/FOMVhCkx/1ThmCQ9jgrYi0IyCum
N25zG7xWwzjx58LTTeV05IilGtvgNPY5ba0bqwzyNdUpvFKuCgLlR52tY2Xq0y77
Wly2+1Ks1wPPfzNhBnpk8JsKsDgvIJag5i6JBf3RzBDwclpSUD7p9LqgEzFRtMmh
exxUQw89+swG/hP5m34iguDvmtERCv710HTwTQQVXppCKpOUDMeDoiKliGqypyDc
kUN/5GZ8G1ObcjIx93eT8+YE5B6JxkEVUh/F4Pv0l7AtkKGfLXwBnfkO8OCji/Md
R7pd40iPguG4B6BL0jL+/L9Yy5/1/tALFCwXMMvZH8LUc3MfUmvZBUCmOQDB9TJe
OiYoZX+HAbARwTWofkD/kRVggodcTO/t/ZRyvxBfHN5NoDQfv+Rg7aNDlpl6VaYp
sOcUi5XQN0fPDVkygqm+6KjO/No4Au1ZTcpbBYAhB6aoQSy8AeqXDN4tbF3K5p/k
KBGBtYVoyN9acz0gqc3g68QtOTSfYZ8eYRcaJmy3d6TnMr9oLvrciLzppzz/4kO5
bOoDasf8iFvyoMwCdWNxQI+VV/BKadEwUZ2ay4D7Qo5Jpjj20kCYIAoFczKJOqII
zliPS56IbrmzYwycYDNEATpzGU8QW5IuWa58RPstsRatSSuKoh9q1rcc3O581DB1
vwXhyylz6UHNGfrCvDydkcvbc3UudsQ1AHmNwg4d07u1vOdj3+cg8AqfS/0jEZIQ
jpwAlVSv7g0ygOXtWlYO4Ojvqcjh1Y6z87Ls9OukwPtxs88uNc7Kdwmr8GJ+AnWC
Aw0yte0cBGO1CbvtCXJIvmgODjbOLJVeVVOpcSwHKG4QDzC7kC2GBciDvTazMH/T
H0ite+TrY2fsRko6Cmw2JgDfvEelx+ZuaWh2aoEziaExQ3Arqm7Ma6x24mWm/JfR
V77ZKGPNJXvjvgo9oZRBS2pff13DFj9XK2PwBqrUhF+K9i2sp3jtAiCvAy3/AF96
4kJJbgF1VpHcWiBCxp57C/i8GSTom1vqMlBHRYHN/q4575LWVpoBRO+UN3VVST1O
mfzcXiKFSHRSrH2pznMqeq9v6yvGTFE2O+jphwITz7UUOch2w8jm+5Yi9zwn7wpi
2vOYoggIO1jwejEEPBQaaorKVgrBC93vWW7e/ELHvkzEPpiUzFcAPLT3Ds2Vxtgd
wTqaunOJNRPf9m/V9gYmQ3xekqL3Vh9eX9RXfdcp+gg59ITfau6JPQwFHLlxjZSn
+ixg1TScQTNBvAl+P7hPZNYpPQPTvbY1LozFhlJK+9yAiBZsLJdpixqDngUCEoXv
BbdRV4NM4lTNMLaNg6FsFJ3Pcdosmcbr+uxztcH4OlfbuIfTLMbk3GeB91/7JJct
2ki73dlUB/BQ0kJ5w8yinCxlcTLG95PArl9vzK/Z0epowUTghTuYj+jLobHGgXyG
gO2hSlmyNH66Et4KwCzoHkVsfe4MW38hlLSMfIppcvkMSrjr+2N8QZao5WmYKi9C
6E7hdFULG0JGrynAdnoIInSOIC15aMmEMnvBAfcbr8B5mG9rHk8lMohkF7IRZn+w
Zv5ALtfLKkPmM7ki2jk8SEdBnz/1MF7eM3spPcGcg9qsyn6gFvUj9KPzZPm90WDI
gAM+n+DTsa6T33nbaaNMx+6X/SvuHAQTs+xYA+104A/CAt9bpxGbWPp6uIXn/Vg1
aiIhjyEsh1GGcyGRz759i4Jzen+s0SWz9K1dMeXea8BWKL1WXU5+7NdMpkqPxFuh
wsdZXKU2gf/J4KcUjZmBHrR7EJi0vubCjJknAnCOq6pZABtYou+GlzOmsiu94XEp
wrFhvXsoyIEkoF3RNhWCku4kh6aYM6l/Kw1eXHo3sqUzrNm7wFRu2APGJ8gehK2K
0+Y271rHE4EPyA85fzEIiz+EBuHu41NXvlfJoGy6kmOu+pO9DxyRiLDO1R2XskNo
nkhbFJlu744Dukyj5u2PoQHRSATTtZnyUhBgSO8DBMAE670z2TSmjY/0/jRFU0Se
pAP0QZa2baM2tzOgd8FQ4VuvA/wxI67ja76llWeSEUh3wRxZWGuGnjRnDNY76rIl
MuaNsF9OphVI9VOhKizfiELKE8aKUx+wvsPdUUDL88x1jFQKlX/f1OdWYssfTy1Y
QXyoBpvP7UA2l5RqTvMcgYuFpRd6IqBqu+FqeCD4KBvjZFN3OYvBE9Pu62ImXw+V
tC/8K7RPJJJU1oqTFk101VGGJukE/O/JqQ5D/fdsZADqptPpIVDDbY/gXMRzxcQV
l8nVYNKjCAJKF2cD8/RShV9W7fe2K7lA6/TbIZs6+fbB/9xP9ACtT+UuuC0H550c
LxB5uwBvFUI8ikxh1daeChrtTMikQLun2ykSooSWJKaon84ZlqA3VwtfWxqz1T2x
Vuhjw15Tb0UzvM2eTXq7Ug6yKUiAxBJJA/S+2mJCRvbX/WvekMHVsMxKdGbE8TQJ
igDtQlsnZBcmxqCS95Izq5o64sXfrckckVc5bAVaSXuCYOjO6xv+tpj1EwOS/+ub
Jmg7WYSYx4vNsKBZ5YefeqNUnhCrJtnRi7nAULNeE4BbdQAnL4h80TvdxGMQ2Jv0
hS6ofhM9aEJVZrOZU9jDwNotUDVVbxFjDlT54cV5+J4=
`pragma protect end_protected
