// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n7D+nMk5lWlLNvNToEgDpIlzkhh0Nj/mNsEDauV7xgfWPwgt5QutQT7d3UC8CweE
E/L1NNC/AcfKhJl2O3Ez1im6KTrbXarr176dbJ3gnJFgtgVLXbWdQrh1Cw2tuxZo
vLusLpvMe17uVwSiZ7UYv2qDkImsBnYwG4w+1xJfwis=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29120)
TubtQPzC5u6zPLBqjWOwK9cnKFyJ2CCd02OqzQC12C+hHQ0z43e3HKxcDZqAAUu6
+eu/ysPBMxkXNJKgbnQm+XA8iiYQZDqQoECjmykBGrFf7rO5aTmXGBCFlytMfzfz
0YqRNeGvz61cD6WRny9UvoNZSMVUXqsSu4vSc/h5WICe94a4tMFGzEKy/geNGv5Y
tUMar6i/QL8QdY2iQh8SRexJZV4m3qes52gVc2E50BoQWGKgJfh0XTMo6zEqPHQ6
X1Iprh44AFEywgc48FrWhxOKBAWmdSvZ7lB+TZGcMwzk89ZJcMFg7t9oM4Ib3fqt
IHf75nMIferVjmJdFBveroB4ARVWL5NNdigVdTY5ZOuofD0d2ZmbZLqHQG21PXbN
t0LtPgbA3KjG/ZLs36rzvN/AYR0tjiTuRKHPTnyjqMDENXFrJ/Ms993RxeUiJgHl
lTybrNf8B9XIi5MD27J8CPC10O2ojOEtB97tunQbrkybZ7cdNk2eAzg8YdKzrbMm
wvIYRTPa4mXD6FgV5763YS/Rv9LYE+U6+mdZJnfS9qihjTs7HSkNzrEP2lUur4kM
CFXgmjE9Ixtv2f43dfuKC+8+avfNo7P01dylXskJ//gHxcJXL72QErtshotXuLFj
on55fBDTHTu4WAFmMP24rMtefBux4nIwLGTC07ZgmiRcHpjxB1sAsRvSqs+Eqy+M
HT91QGpO58mCPblszBCX3utzB8qdJDuFGk9TCdhOJEA4RyReGUlt0xOzWlH8ToRG
bABjlPedJaCT6TUbpcGy8Q3vECiiZXQUP4jjanS8V1cXLAOonfH8r0yUxZa6WnIn
UORYp1O1uxVvj1sWwKOm37Vrb6adk8LXMUQq++o98PZSg7hbw9oZoookZJCwYD+N
gXmBVdz8+A1y0p3/br1OFQTvtvOcCw1bOj/b0gAz8iHJSdlDiSv8C8AHZC9XZNp2
mQZ99lZVVT8ckBtk5mS83C6ZnuKk9qJ7GUYgLvK6EdECNlYE9vTFbGCZkt2GzC/7
WPD1fpiAuGMb1TkD94ujpj7wvg1yQUzBOrfjh6DlYUqVdEBVyDVLcyYH/Hw/11Mk
JqmpJv7uryBDcOjHDOwnfL3P+nudFn/TQjIutDLFYes8Y6H2SGzP02UTBpNr5y95
Qxr35yPa5Z6jMq2SXlg8WJW3XN5sK/QznBGj34mGqzVa2IxaWsQAUVttY4FP5l6X
XzcdHnFd/PG5TLVEhYhZXeXIuzFL0/V8OYZFeVXi1QYP750Vs+uWSXLdZZEB/OCF
81slR5iK4m5wkyIT0QCFwsqviDdCDrjCS/CdfBbjBhRYWoujaKR0C7V0+sNyNIFg
VL/b1nxJLWL84CTprKRhBghDC0TF/yGPr1Ak6TzdqKFdkHeKDb3h5ktVgP2L9UNA
NbZ215ZfTfBth5cr4elN773e8H7uhyNGgmfUbCjLkfjkUI7dGwtmrm3+wFALgT+m
uVkliH5zg27X1k+2xnI4ztY9N+QBX7nz4eifsRUNJVl4WED9wdYK4urhnxSpUZe8
UvwcQfxpcq/4qF7V1MJFKAxb8+nZOqhYhRLFVH11I+v99UdR8oi/mKCOXD2WZE29
hbSKwh8Z25YPv6l5AaImT0163X2n2FW5ovhE52SrbN8dwgwbOmK1oeY6L7jJA5pL
gRKticwUmZwpKnYdSQfVlKUmtMFV4bj4Owjdnqmj1GcRbmtOeCJSdWWNCbLo76Q7
uMJ4SblDRsE/z0Y+0u2iUUdwVk7YYzQBQ/fFQcYy/cckJrlK3ywg/h717j8G0pxl
ZTdsZ7lLNaFlNHoHJgWiRcFkK1PL9NaoRupe95w0ijh4WEq4GB8bEhjCFtxgt7LT
Uq4KYTY0+GPeyBO7cOjtkNMez3E/6By3HX9PKUPe75lI9KhvIMncBqhoByzF/je7
fbl+ebCr7n4WzxANtE456/1LXhd9cfv0ORG3llpmfXhS25nXLZeevoQXCX6BHh8o
4huQFGkkJayJDWiWp/8vtEP7Ip1jH39g/+xOf/0lt+LgT0e5P7p4M7LnB8j3qlSj
PLoO9zgOftx9XvbhCJT9nkYlWKBWsosK7dnMaoHDAX5lX5iL4yJouF7acZGA9bpg
dZCrqzxHZlDcgljJpk00Eg3fJ8GptJtqLRnNLzZ3C3OYGghAd1dfgErIY3hUOhA8
fqYIDsXgBaJjVVy8aoZWKQynH3J4AUjckK8bJGpn932NvXB9qu4oVf7J+MRAP3Gj
f/D9u3/dvidY35F13JSOXy2+AUROahp1qASAJuq3I41QneqFkLO/8bu6ZRW9O9h1
EB/UartX8dR4x82/bmcgc5owNQw0ZtnVmjkmMFDmEYTNvJ6rvVIl5p/TXmw1NpZB
h/4Sg3zHk44wjnqAQfn94RIyImN2PJMg0UpiLj/UCtrq027Gb7UQuqtvMWI1SsnF
lDQazEWVo3C1kybT6Bh1ltNIDScF3VUSs6LMdaSj1vqQabr4y5teFHN9HrrTWaL2
8pZgjIFKURObrzJlmdPVcjHR4acw2qowuK5XTCfqlClZkehlYXEMfKEkw2IzwP/l
exRGk/nF7PsSBFe26KhhWKgtlSuTbaEOZE7AWjh+wZ0mkySt1ksXILoVscdUy+cY
C9fWjyN8w+RrETBbH4k5ubn+veqDR7jeoR3LraeoBJaR6OfzT5M9l3LwW4Ikqg+6
QybrmEu2kMhfmZmbO5honr/ywheK0A6JSSVajMHQdTC/piH0owMFPTrAdxecpoo6
vUJYqzi45Z0/JeQnnDkA/i6+vHcqcCbkaNKHGpAr86GbzH5u/rtnvGOj4lIUBmhp
fTVWYg4Szt9pSiQ5YahAfgz8kTGCgMXEL/d5qVSv7qFpZVclHFNQdnCmCco13V9N
KOzNpO3sKJYlljVORQtVYrXC40GeO1c53p7n/esyjpLUKQ9vmllfkyLC56CtwPbn
dh2MbtkT3gD2KAuXYRHxZekbJ1f7qHkQsctdWdH7YmIGZihsNwFgfTw6BkwQif3+
DcYolMD38YzOHsGOMCplZRRQ47QEemumnqD5k5TmPb5hq6cxgrt+4kwJ1hnuJO8L
84AtR93o8WJ7fLxXmmNhfRqbqpCgDLgY41mpKFEiZnL1WcWd3nYi7wiIJkk7tla0
i2ZLxD8D/I4NyCq+Bj65gZzbV4w7mZwduE8hat7UMwn+3YivEbX6p0hz+BHWs2vO
ZFD6357u0tc8yADIO/DjR5YTJokFNwuOY8+vD8FAelqcmqYmc9EuhMxllJ/kSBX0
Fuc7Bsbgk4QBmRlRhtopU6j5FbFGKbYpFSLs7VNgZDacPVhmxCBiL4GiVVfzXgyQ
slptA1TQ6MC8MlRfgBzNDRJYrQM57gHgY7rAsQkIIx4QUEJ7cfF0iC+RQo9ohWFn
rtLVcQQhwjmCxjBFwvXNbhzzLywRIXhdU9P2D7iCbUTzte07AeLg6nYYUjFX0SoO
l6P6MPvFLqnHY8aWreTVIj7GZURoEsRQ3f0GqMu+SU16PPQq8jPF5aPM6ucoANsV
gL643fy1puP66g06RF09XfBUf+LncQxznU7ATzvdPqJoqXOIOIehzM3Cfjcy9D8s
oDMG7NDOWaKsBFipq0+LOw+/2T7nIlWbsxp6Br1FUirPL/V9s7WbhC+iAM7D26SO
k8LE4Sd3B/LCGD6aQI88w2B2gAr/pSN5tUFNN/gNqE3JumwLmPwOkeMzONASHmlq
zT4PE/rG3VyY2+3Tmj4kn2eXPKr0401MLUYyGlSHIJAJskU2VlPgx8VpW24nxAd/
HSoANjBCKpo2eNf59+vTN9QQUTwcCkOwPGMa0EFehBsl3dc66U/Ph7YYFBeGo8xI
h0HTC62Lz4z5jkMz3GYUqM/CrZAr2joDw5Uox5wkHj4ZO5j09pYN4N/lloP70JEA
ojeiRu9XssFKTLWnhOlUD7COKUAQGzI8osCJl8FCU2dCEgoasxQNpFUQdcNJQKYv
iJ9PV10W1iseyDqR4K4t3tLo2Vvlg/GZjUZx0v4s7VZmQiXc+rjif+0JUnDs7s5P
M/wcFLJobj7/TJI3gZ/flSABtHzXWcz6jyPuuHG3iC0f+r9zAmuAK+AApafb9ZYv
dDnxD4S78RNB0zswqTybbsnJr1dovpyfeJnYdDenhHACNfVo7f6Y4ZItxnV3n0PZ
s21C7iGwympsO/PKfUeWoSlfEBdMqA3vxbhYKdTqZpESJNpT/xKBuz8uGPprmOH7
HXJLxJRlxX+kZGA2MyVEejo9GDiM4Zv1EZgGAD/eeQn8FdQHNF3wMrHe509EyCTA
pN8FilX/cuX92msckRGMLNGgV6fv00SG2s83rNEx/XSACF/renuypnPaYkjQL++z
G9NqYg6yvk2g0tlX+IcpAn7Q3vW8SlG7xlHDTWFFcDVc28w5cjcgydBKmmrgqS+2
//7E/5X6tcqpsJ1YUDFuZxDDXxKX1XCYAZZQ/JeYsLehJM+TZDRqn9U0ZQWORDVd
5Y2vn1Is/fu9O4vpj3bIccvDggwdt1hZIYvMy5v1z0xRtZ+wSdpx1qwFpe2tYuN5
KW4TKWcK4dUZREVUhbWlWBKfwItNpbIOhknqpvzto8VKv32TDciYoDFuu+HCPLQA
Z/EOdh+eVW2M5ZThGGf0L4u+gT6lJpVjcepv7djVR/zRatYgFbu/ocvJhAVTc65P
WerYUrPiZd0G+lWv94hmxnxj4qhgq02BL4WOsIkqTlCk8Ov4Ir68neER7xOFpLWf
UBQRUdei/szX/q91l7N9oJHhG1aAbhhBdgHo2oeN/JmdJlowAD7FXEPgfbqlHsCi
HaXq3CRbrg7yuBEY2tAfrJkx9Fuz/B10AVHgAyajtniUC5U4cl6Ypk1XNZc2t6wB
Ptzm+kjzIFDiD7dw+Io+MRUwaneiDw5vLwo+y6KtS1hyRsf1YxaCLLNS3Qg5q1vG
Pw50/urG5bEjqN1OF+brnCrfA8BWA2mhjuKxbOY+f1CFr+1KbFuzdLxHJP+9pP9Z
NFfMfRtKcGdCLwadqj1mor/P8n13INKSGMsExutYslrw9B4xM1nfIXBhSAdJm1cJ
eb1zabc4WbhO/DKp85U/JcfXssuQd1wWfNi2NAMKgVZRd/+sVUNMGieW9c1MMwIY
UZcvXxyWTxotXB9jD272spxuMIEM/w6iccQVX+wDZvguoCFdgFivM+8p5jbvgpB2
rDxJ1TPBf26trK7MSipQJ3p6B3fWWEsSz4iU0vLStadehe8JR8ENKFpl6BE3d/TB
ZTK9WRqfO63xwi2DKiw7bxhSasy7lHL/oxDvRfmEF8G5QUvuESUVXla08bP/rcmm
6PNwDshIrIHB0vVFBkDh/FXvkAWkI6wzhWSCoyLCtBOjHnuCfSTvs/JTs03qrNuC
CqCcGH6e036qYP70OF2FfTXJIjKpHtYeFa34xZtzP/3vPaiZD1SPhd72vT9gfqnH
lJzECae1w2Op7Zrvn+cF+JGPDoVq0zLmO9xeU5kHYNhLQ4v4VuF9JDh1j3uWR9E9
JRsBxEbYRtiQK2DTF4uEiQ9NQkCKSytDiTmh9ENe7YMt4t3naBYBKAphqRMv1dCX
F2ogrDpZdOkfPvNbiAhNf8EeTo+A82QXTJjn+Xp6ZuC68KT0DLWlwrN1g8KJpAq3
Wae0pz06bmPLQtorSZCV0AKwdzEIxEVLp1PYDe/SAKv+eG8atOWTJyW3B/8fe0Zf
oyDGDJPGUKyaJ0VK6Uvy23DzhW3kzKBX38tOMLMbgPNSoUZg5dKivKy6iUmEjHP5
q+5LydLferfZ9ETGQD0Az/nDEc8bCW01pQEY/+mpxDNhsvQ+B5HhZFM+qVABpY9Q
/4ByQv00IyAuqpgybQvtTgApD8eh/I2Tscjv8NUWPAf03I4pCCwiF8dQcHes5azn
PEMCqozrv6uI4CtPMajMhzNUqRV6y2DbkPV3SMO6+XhQh6dlIHbA2KJnCqi0AWzY
fR6XJnpUjASeYyIgL1yXxpcCS02Xt4p5O08mRqAh6VPX5NgVA6NOQZjSPtpu2eX1
+hgj7tRBCB27Ye5RiVGSpvjWQYFzDedvcJkI/CouHCz/BF+GgjhFarsTitQOtcxl
OBZUJoKoSjZR1l4k+lM9Fh2OP7YHOjcMLgS0ProWdh2JxRMvAA+SFrCbD7j5H741
rGW6PQQLKX6fIoSWOSeHla2OxZxxzoKezPfD4rKpVBMConBKijlF8YwegVhm4Lyr
GhbB/TaeYIOrufz4kkqcU/aqb6Zcq8DU4VQGk3LV1bJUa+ESQMtk7FrN5FUryaAn
0qz7McihVfWscq5hvTm4OyBUM7gR6fU5qeAuGqed4FaEeTrecqVbI3VBmCBs1tth
RQ+8tyLrXDj+ZmeP1SFLpT2jBdFla4P2H5/AGw99qKoZiDUw6Ou4T2Qu907AZRK5
bUNjWY7YlcZj5II9+MgK2s1PRpZxa2zc8A+4kLd6k0DT4y2Y5eLD49U0O9EuMieG
QJC0k9rZ6CJzcXoSY2hQmzIhJbb+IZMFa6KZNbRN0MZ/4s/LSFGAO9osird1G5rC
vRdeQMAgIKjLW4AJn7QZyhDJPV1aoVqXPGJbFkVV7x8vsp+v0ypjiWFFQLGPpnzQ
WSMq7qmlKf/TGB74tdt0N+nbVXg3HY8UiyFs33JzzrIMaXYqsRiiBbomSVP/fBh8
SntGui90YVWSL89juRmrF5BWWDCq6sotNND1OgfG5irDC66iYbuSvtWeEqFBuTT7
pP2+Wv7ZdDhIaBxTK1Jyk8u2szsPgXa25gibhCnt3oOvwAcDcHJNJxSyGcZ+Zk24
ANL4y1xmFi+f7iO4Vuoj+coUl1eBnazhGbBsKNn16WToz6hU6PdqECeetk0lJJ3D
/HLRxCHaG4wCchWvk69uNqa2pRLx5yIwAfhL1497stgZcm9MndmECKN3KDIf3rkt
uYHvUkq6T3W6jOK1XBTqAWLqYLPHbbOcCo6c9s+ZaGK6mdgntRkqVTeUI9PqNXFA
SSsJL4dKbq1Q68TcQtwc0JDoy3FzP7FuXg7IJveahsZFhtQ7e8FoTsttijaQATQZ
WI137lLG44veu7EQlIWs3gqHlrc7xT07+O+K5YDJ1Hfj42XdYFQGQeAUmei9/cjM
3alE4Ntjy+OU39hPT+0EhgMV7+kiRdTgWX+QVe1FBvj/X18NhK1wcWTft4949src
5v+YIcQA3w5rISKs+mOhgfCvXLug1owarpV9OwSAcw/GOc1mGpjJzM1C6RrxVXYD
Lou2exPmA/k3jjwwSQRfXfYVv9UDrAjIrq+IkRRzWvzdoBbsVuAkb0STe1UhBJEm
+Pylirbjc1Z4ODh3NaG1Ivvei8X1SwChE5VoZDFxqsXAUR6FP/blndpPB09bG6ar
8n3aO2K7EenpqyjVNTVG8cfLu7YuFdBETIs2IxQkHtJnyfOn4E/OMFGkFrdNVuI3
hJIOgZLTwUpTiVaT0D02dHkleikJV+jtWEdIV99AKmQu4eWJuVz35VPtyosILBx5
T+9X0sniN8kO4chuRMFT/YQBLdkpvVyypwXbJ/yhSoB1X1u5g6jq4uVqpphsCpKD
fJYpYsmLmiLABNeQ13rEAcB3tqkjW2BA2ZB6hzm/x7U1DwsuUU6TOHVN9KcGZF+z
3Ssh8MyUaHhqJ7NWRwoWne72Yz8h1YrhxHKtRXggraBQbLL7zRqI/Uwf2bQJcHag
XeLk5V0N4bi6J7EzLHACP3+5QHAdmqeS4vgMGpCxi5zxi2DJFG7uS0UwggHZ3sgQ
AWqE+Upc978dzMFbGXJbHPYryuNJNxvbpi4JNDnrQgbKAFUuiXOy+p6cnZHkee8t
8Qid2TsFwo47tI+s0B8NMNOhxI5acp1lxg/rsj9lRYJwSmVSC7Sl9a1Sg/1iw5O0
jMVvDXRnXSSc7eLODyDwQWb1S1+REkh7b6IV9+1sTrWXcm/klnXd5znneJkw0cVF
EAGD/UkPe4dtycL6frjSUoh78ZAn/KvBW1i/Vhm6fSh9M9WSv6fSNh30feMJTlJG
+gP+pUMsLaM8R6k/8CatiaQnf3vJvMRwVexlWJ5ih1W2dyONlsBCN4xkSUv5JkRi
zEzDINWGPmwHxPI2fIcESVWExJhqGMyU4aBhBIRrqq3CrpxMNdw5m7I038okHeC5
ixa7hVBqHgYTzm/VBl3tgfpgRaNLCivtPjCUCskvxm5Lt6UzPy+xfGiOwH9AUiIY
u8Um7aHsBt7MVfWbfEGQYybuWAkQcjmnaK421uqpgor6Z3TaEVnnCG8erTxY37YA
ExdUyPjy36Mkk9ViCjVTBPvsea3GKhwbVW1BIHiRayUMkN+bYbt83DNINiddZMjE
1lxsJpQPhFR8UFipzztH4enJpFPv5K5cOsY44VCurF7OnirT+PCsW6xOv3aNZQcz
OGUWtB76qGtszJerQ3/TcCIVRgmSZgIEYSdh5j1JY8XbLVcClU71q/1eZU+vn/3q
Xp0jQkOKBAchxniOVf7xuNU7BoutxIhUB8H0gaFUIoIbvHe5UZE+6H5ItupUrB4s
9V/Fd7IMZMpolhiREB/snHxG7hnHMnwCsZNDC+Syh07+It2TuAydqqTAO4IX99LF
MbOXIl3RCjj0yazFIzI8fb5O6QUj+mjq2/kEkz28ZIdJgYJVDjGpLLop2B0Y9g6A
pm2BxdtigKSd05MzLlf8w+US0bmRUk1y+HFlw8BRkxB9u8aMxccs1E78OVB53HQt
A4HRMW8ty5nG74p7uD05V0slMt1SE/J6gesKRS3Plq3iYGKbbr2curWlsvh29wkp
SfxegACnADXAOvjoikTcnsHB1FkOEU4ndgypB+oTRIBYdS/Y/00HJ5Ep1B8dVBrv
rcivfMzowg/729DUBXaQB8vgvygqOdptzxhzFHSrPnEOM7lBjQRo0gwbhp1ZJp5b
a0flyCSFcfgIgWic4UD8FdJKrrc1sLsrooJw8VXaxzvE4olm3S71RHaW6cCblRkP
57CgFXTKiK1USf1o4RACvYRPz9AIJ4k4ZQjLdxdvWZBASmWImqFEYo/9bldXuxm0
tTSe5yt9VlB+5D24jnkDH6vd4VgIa2kG/2ehwKM7cvaf0P8kX34Ky1zj6oaQAoG8
mKeQChydSyki4RvNixDOjdj1bkb/gegz2Foa+sOyqUuo+/oce6MERMY/bk8HxMco
dlhUPJLwI4NLEAth0i6+1Ejxn/D5oWxts+A3bpqCclxpBtHIo/78K+pbYIrv86Rv
58eMZ392NoeGoD8yQJMCazg0typgpUZAzKgwNwjedZImTKiX+tGsBlRk8aChfvkE
OTMxlAHRdf40hnPShTm8F6OyJ6KaVhuHzXCyNW3C43fzirMBPHqLruKBmZJFg/05
5+Wqk9aPOVwxRqul/KpA+vxzlIXF4t118ghLqbkHyf0r4Gbb7bF0JuIoQoakKDwk
W6pScs73heYh5U3KzrqALvX9eOTKnXnHTZhM633zvA7b3ki8lI0V4uv69Mgibukm
t8q7ttQBPNmXR74CYo5OLpUH8I0amBDpPyPbIF6UAYav4kha3QNm6IM0kWW+MdwD
uff4XyxrW4Cri7mDDKZsgT+jWz7cruoyzO0SxCcs9W5zIfLJBlF6NhfygtQSzULd
aIzV31vL6OGzjmapHSwa4M2ecU0ww2vQCXszaZynQlXnvV6XQpVS0xN5RE0hM0IE
RjN7JAefEk0tOvTtkZUNTaQoSqm/IMMOe5hk11T3ERrgQalMoSF/gFwORZmy+Gs7
TH7eqO0AFOKLBS1zbARr0ijF54Vvk15KukgGvHFdg/Wq/uh7fC4qs4g4KQGLqYKl
am8KQT1iTR9fbo9Mg14qXwtGEeS3ZX9gbC6Gs/pQ/yrMfn1AfdM7tJ3qNSijSc41
PQ0DG+yCt3TRdoKexRzkgsI/iuNXXYs+K8pTO8l0lDlJookn70+kc0KvIvcqH5KX
9D2aYaOW0a9hTh+xnu6za1aUC9d67iU/GqoUE2kk+pH19vUc6J3fHY5XCUl9LVGp
JqiokDh7XGkQvugUsAfmNCoBtJ7jRDq1YceKzNDDZyu0UvwDnlHT32eSsyyrs+Ep
cwPumRUjeow8Q3P8pZ1lvSwNbrMa0xTX9thFGrFb62834Y/Pv24xufpVfTBFVECq
clXeqpnw/hb13/ooIP1WjkR2LJMozIOGeRU6G2uxeXoMCA7x5yuzEQiWJdhYHdcx
w8F4hh4iLxro4t6hPwI1xR1ay/LATC5xptGN6FB2blRdCom3SEPODhbAe2/B4oOE
menVjKu8F4uWjLQDd1Mc5sQ4JBRdt8HNPa42D9pNNpdOzCsKJ5vOKnqQ17oer879
3ThycNrj4cLE5dsuf2KqXMKbX+IX+NDXD+E8XIB+9wwz0RdUDLCWZ7qbSmDvPy1o
xoWJ2i/6iLEp/dXdLoXQQ+IpdeqP9QYuNcTNRjNjgCudkhgACgm5Y84geyjaVjo8
ABFN3LRjePon1pLJw/6aCPxSPyOtZBxPXTzJntHqs0BN9mLXV7W0wgkAMv/ipMqn
SOECffpCb8a5+uUeXIkCnSqhfQptUx1buR5cwCcA5mnVCO81TUbGpzHr5yOBto3X
30V1Q+3YJl7pCyLgs/KrD8819uG+noivsRihVUNcNhlTyHsUV5pVWrMbw2dlxCHC
t/+TNFPmBUpa3brcZebMh3CLASdUcyR2nosEKqMioSzj/zr7GPrwZkCfIs46ZA3h
aOJrVtowW84pyRF6K0ptl3rh0b7K6XEfTaC2r4/9e6uGgNPtBFLBZYUgLZxz3kIg
Sk66p1iNuiAPNmF6zOyfNdG27/iVqw8rx0NLC6AhZNuJDGKSZebfx1SkYGyuqt1/
U3h36x0PCtZLoYr7txaXgDPFsr8RS77DA6UDsHotfue3xDF4Sllk0gN80/iZOnky
GW3fkQrNw/ZFQrud7AgzgOZEtj/KcMnd3ROXnKFMIsvrrptZHddcrxqSNUG5Ccuo
YHjWhaxOwbY2DRurjOT8PhkIXupfWzjNE6OovEiTtytQg/RVUc06jGZN6ueKJMOo
zRRmrW9YxrtIJWJfsAI1XXZtUz0/kNTWQ3AmBMaG90dU34jWwfPOGLnlpcoOC8tq
zWEHbMPLwWsmHtlu6ZWLnopElAFplzwNvFRhdUqJa3Grb/XJ2F3owW6y1tfLVWw4
jmjSt3uC5Sa1jQKbWzZPQDm8DCaEq+MPqc9bVPyJkxJDqG7TxV9jZGyZ0FlLmAvH
wqhob+OrcddUfDa7MpuCd48lpE+RjlMO0U+3yjQ+BA7vGQrT92Z1hu0YSdLWN4dn
ZMR/j9yI7UwW54c+hTN/DlLRj5Eyms604QcnkQo4EVRPIHA/rGMAlpl4EhgXogr1
jI1PH8T+w+5qnNNhrbhaiFM1+acJySGeelvdcobvLc6NVNZNJYf3pSSjgaR81PwR
m0dSgmbjlzMLLpNlhwI0DuMi7fs/BK/dxZ8cJfV9SsPVRwi6CE7NhpbGotZqQibh
7Zks33wejp5Uph2X3jBmvb85QVUmyQmIFNjXQGanq/xIPXTeaMJp47w2//H/G/3x
C4iOLiqqVmCR1GaWD+sObu4lMsK7y++fjJmqLdqUFJK2SmSVigRoit6BwPyj68SC
J3/bDn/UuRKEluOt6SJBd3YU1pzXkufapOdi1yCjLh7ywhLM+FBIo0o5o01aOxUJ
LHj/K3jRvPNOrhqBXyvb6tKfp3Q8c+7foZDqKviY7nWWIS3NC7+s8fnZsXwGqIt2
PSSuA6HkNjp2UQvJtIzI6P40UPysCiRhOoXpOiOH/XO2dW5erewErKOmbNjY4ENk
FfBRKcAwVUtNuy1CU5p12s89WzHj7lflQuyGQcgnRafeFSOzpuFfjA0dpLTac218
+5LV3NMVZnah7aUhRMYXVBNiQcp35lCQPYPL0EQ4++TAfBLyUme9pBeJ3QSMewJ3
swHnbUvzLMpPvvEVWAxDM02V+z9IO2f+gmL3YKUQIb4UJZZdjgOE3HMPMMTHAZZK
Kh/dvM7mFFqj7E3eZWOIXqx0EmPfjyasUflGROTky5lXJJE5FkzNRLOq+SvgKkq5
83ATL/mP45An/b/YZgkm5ilAgdsPubiMntUjgw5SVqPV0o2z0aT+i6ar6mMIwA9X
HwxalLESRLA6HH2+Pdjy/RLWOHKbgYPMD9Vu+XdXXTfUkKhFFo+h3VCEDQze87hN
wQGAkEnEEAPHfvG+bEJY43sa2f8ohCMR/JMVDdI/bZe+NtROcXHVwkhSpPvCLdHV
7tqoRoBgPA/JwyfSKIN7wQUgEDEMYV/XZIvdJACE6YSXwOwD26C3nw6KBb+ixeb8
/NtGdN6aH4O16ENP3oryYQJIXVm9UrBhm33nICHPgDWy5jmOZ5GrwevX6lwf3JPd
pbhh/Vscq1q92MUBolVCz5Neu03FZE9nwysVTyJzoW3Sr229XYrURXqfy+zfGJlN
cqE6utUT3RvyAJVtTNj6N/nPYa6lljyp85LVbqtkR3VWB+g4oiv55XHHZm8YXmkw
4UbMicMv3tbARTYkFKKH8a3aC5jWIu1bLo1H7IzdqUimJ8qo6wlQhOSfJ+tAtnLV
j0j41FbWhuKvbEadtM76YbbLVivyiLVtMmLw9wuhB4CtnMpkcbxGmKyUnQtrnpGd
OsN5dn2K6seacHU2bmRhYVWPZ9LpbSWiY0QWHlJ11mzLg4Q9Vb484jk27huFxRkz
ozCEiFV7ytQfntGriAb+AUdd4RIIo8nB+6niZa9f/o+fpavV236jpHdVwRzvHDb9
8SwoY9g4hMklCamr0FlpbKYjdIkJR6xjsMLd1Putl4x+9hQIBarm4AVWe9UnTTC0
jqbszvKC1MYgb3JTVgYhWsSo5r+b55RTNXni5bzOIWSRod4AlNoE/ocns/6Y7T2B
CPpj39k3vJaIBihSxkHWbg3mtAHeNjKGKMr1mbYWQJAC7eu5FExXFNrNsa656Fgi
mbFKPnOC7+4kTRhEjlyGYZqEfew2Wx69y3f/Y2An8Z8LTcU/vbSMw9snnXJ9he9C
MsI3EaE/i3kb9XARVNaoxEVClNuE7N9yJ9tar2XanANPcvSXdk8edkncn3f5laqa
wY9IwqqeajiehxTa86jXbxnKvnJudWXd6xipCzDF1xea0Y29kgpAw9D/SbHYlMOF
6sYIupRnAR7j9Cs01qmBS2soMwOZxGeiHWQyQnxiIQLlvwB64hhDBknXRsc2gXE+
HAuo7WYMvUTgTXq+oe77JsZfuhblSBBHmw/zVp/Knoyx1feBNTYTIfqTfsm7EVPG
HOiER9rkVs6zt0JF3PqLqOyO4UxUef5q4No5YhQgY0zFLtTkxc1meNJ1NK2VJOT6
UxheLR8IHLbE9LhKIZcppUOk0rRyPeZoED2kbklwaCzU/7DmOIPs+joQFYCGleI9
yNLWlMDIgHlERsOdeEBC+lDtmeA04Mg1wy05HxzwlOQKjqFJPSx1+UFABV4HSd/z
KB6XnWaIcGOUPvshO3BilFPe+K9I0nKJTWtF/6MSGX75UEFqz8GaxsqcNaoMm/MY
8/dCRxZNnVEG9LG1AogfG+TY3mdVHJutF/R/U+s4wuA0pq7RZPmjJl9T0PfOo4fE
BZeCDsxDHlZdd5fFji+w+A+T/QFCa1DXu2wV2XElulT+GrUSET22g/V2w1hay65D
Z82Zx10D5mvyGhMGD/IkzVlzFRH68qeQguiX1nzENwCRYh4A3GvDXltLJp7eQ1sr
bfhEw06S/1WpJ7OyxVeKp8DjvfD8uWoD8BeOAGqPQ6DGol7SAPck02aT1ZKkr7GV
D6T7yfHhfwkooeNsFdlhAlXQquuOLVMdYkpX41Yw5v1TeYb366Cnho27DHtpaftR
Mm5oS4+V1aFzTaiQAPqqnHaZhAX9/t6Yb8g2i7i0jvN9kZFZdZ3dEVa7g0Tu4igQ
+hqPqt2QteVQIPYfxywjV3TqtUIbI185UgvoCMAZcB52V1vIy2ViTAHt7SDOvfzq
jPLrcTXyHMfwcjyUcfnmPwQTs5eRxRHzDVH/GoE5hihsgALLlYl108JEnqsL7b+S
GgcsHe30KuUimOVehaN1Rx+Iy9NvkKss9cJLuic1Q37j6Tl43QtjyvHs8kbskSFE
et4xaXw+ucb1RS4H9E+bmhMIqQPhKoVrOBNjeq+Qv4sEnLMLoxftDismCcR1hlin
F1IQp9IX0DedtR4JV2c/r6u2ZJPN9bq6bmRbFxVHWQdGRsnAWwI66bjf5B9gjQnr
1+aMas4N/ZgB5sLffMKCVzSbyfQUn3Fg8zyiUYKnTvZRsYUXVfVLopbCglTQk9G6
8L7SOlyM2L5d1+FBJCn/zRFqok0eO2vE4CJz1a+WEWoNRWLXPzv4pGI2MqlOYuKI
erO/ftE3sZXAs02K+Jg4sJA8Qk5ybS3ycomgXafPYFlBvRK7G5BhpP6q/vquAZw7
8bJLy3VjkkiaiMl/R+lbCDJVamjxWdQj30L48SuXJ7wDfkzk8Jo09g/Y81B71M1d
yr58NTMzBjmgdLbGA1YN/PCVdC7ulvVEPSqdyLV6SC50/hcrm3TnYXVUXQMjLKjK
m11ScazcVyAuh/7x4MkTk1fwb6Uqcpz6+RdU1bb6b5kfWcUFoRnojPUXWOAmxWVh
lgFJSaVnmTedebBgbHY0zt+HB+X/FvLHJU3tyyr3bpl4X+7A9UwcLZaMALr7GQnt
tmfyeQ+y/g5v/sqSEsMuNl9CLuHcX6yRu6YjunWtOzoV4sfmdDiomO10eTZGdHRT
/GlamKwYrr0Z7XTfdz1XEYRRwpD1+hSnlHwUVlLSfId6bjyrVigCgzvvGOfM+QYW
s8x/goyFFuTPBKG8/tJLK5cOk0Al7QrMBCoBB4IbuqGo7RtcHjGf57Zkxag4qVxj
hbgnkTfy2InmpGjSr6dvetsjGHMg1fT52ies9DNWLU0eO2AwRcna1byPntr85ISm
Rz3yrLp6hZ/3q/CpQMXqlkBPSg9wOuQNzKnj0nosgOR6dOtXY7+gNhjS3PbP2czN
8NSm/4bV6LAoiDaDNgBkH5Gl3gjqkzj0VzpbZ7I4fBEvv5oApf4UPON2HGCX/fBp
pDRQ7VfGVMOr8fVDg8v3NftlMTBADWiUfkhsc9diK76ZL9TadXvB/wWRx5M4vavw
kXfcCahkT8Pge3+HKNyfzk4Ezq6OgHqL1e/gtN42UBaQKtm5lAIVZUBmqXpluCbB
N+EulhqTv8sfRlAguOo2eGXdwETaxQRqIhUs9/uJkwYTgJHqSr9L8RPdLNMDZrEE
1haCiQQYWigtt4nri6lXZi3LO41hOQ3KQ4FAMbuJdrigI3+q4Yd6xtP3Ggk7Fw1q
oaNCAo0qR2O9nsE+IN1wp5qoNy7AYqSMNMcDT8as0Nxr76O+h8QEH5TyYKywilD9
rLjTXAtrdpOlVHiexH8mxt21/W9RU/+6yrPP78TnoG+p2p6Fvr24hNeUoZansqBa
Wbjl3BD0/q7Z67pOc9oW1mUIR8MuyVEpA9xBkzcyBACr9ofvoEyahkVRDgF1mJXI
WWlVs6Ln/0rIbSV0ljOgX6MInjdAvZxNU2bZrElsyYYPZCamUjIF+NkO3wd28Irb
LdBSFQxoJmbhPwU6fnDIQBb/TMchxHnDeDDaMpo0ifofuSjLumrR3wXg3tHYE0rC
odgXazs2qUj9HRCLkTWACGshmGcefDvi3W3MW6J36v3jzqPGjXPi6mwHDd01CVzg
rraSmL7zKwoARqDlGEbBPeyY/ldg3ugg94xg+n+U7ath/puMzpV+ePNGj6ElXgYn
22zQUJl/WFIhyAFz0xDfYNf8B5N5QnBr9fumqvd3YmoJf9tYSdFQItLZ5q1nw8OS
bCufHdg+OfZb+GS8UdIsFoWe0xFhtFi4StI0TtOdPJqFpjc8NJxqKQ+L+Squy6v8
kAkvHkao3X5e/p9hUnPTQbrYPMQSvXBkXz03BaiPIdwmTMnfoMgZbox6MCZctjZw
8ugYJD5briwNExBiSZFrT0WGccAd/ETqMoDYVjGQ5nStOUB2Ypx8COz/3it7fOZT
nS9IgLAx1vgH5rHdfWU2YFaysqA3CkxYVKrHZENJ20a4RZTA1ewNvzYsKaHVc8ta
C4k5EeLmKy/0+FruO4AG+dV0uKs0ueGVoz+L64vbgI9ESW/NnRDiNRaIX4iuQ1LQ
jJpqACJyrC6TEQjjua2jVHYqVdhCVtszxfXusKoaP6kajRO7QCsR6CpvwZrx9lJl
yAp2ICDz3ktNmP+Yen40a4UPx3igAh+d7GBl03KQCLwL3M5I8HhmlC7R+0/lm6FE
c3U+3aa7SU9IBMD/tprCz0Lazxaa3pCE+japtgEJuPbVJ0gvl451csSNrvR/kcCg
1dpRX+M4VvaBtbf3sH1zOzEEdUOX4+7lz/N9i+RzuzVYWdrB5o1QVTo/CFRHKZj3
6b62ZiOcu4JydgzPt6dL1+DBiZZ10J/xOgWhAMf8MqHWPIUX0c7qtzuAYHMTyDy0
88X2AkoRe/N7PW3d8JeVKRteTVENv5n2JiCcXhaMjEjJFYAPNlTquCwjY0vYISZC
Nx4KDVmx4uaN/aAZna/Vlni2jvZExbmuYxMA7Vy+/ZD2+Kaa7faKLPnk4EqwTO1G
/4T7dNOoC4aGV4jF1VFU7+bvjBxRu9x+ZTrRHeIT1NQt/r/vdVMZPTKf47FNtJXV
GVmAO/wRIuAddHPecg2NXZyk2Nmz4pm/kkdYO4mQvF9AvLW/Krq1IkDVdW2EUrCf
F1sqN5/QnaRFjxNCDZ3v43yXN2jWUvokYoaPvsH35+Tu4l20chHgh5zJqSzwkv7J
WyohePvl6J0/RtJTjSk14cfAcV1Tbk5gkXhYpz8rnPLbQ8auIWyfBnJ/CWVKi7Sb
oXj/SgwN01AJb0iQMNZ1tPR29otpCKFHufz3HApHXf0yKmKShkIHvACtUITmQ5Uh
Rbnz+vX7RZ5nNg43MmG368THBJhyEtrTbtmjTrn5XCGXpBJHWQKADjMAVmb9bYEc
wLprHSZjpU0fwddwuVXZkFXptlvKcdOAgKv+kPcn5rvy2SPKHI3Gg3/fTSLO9MyA
4ruEljouCfTpZuoK0hVLkJoznNUpDT8//6NwEv+RqivvLd+vtLIWv8AK+qXrSlEv
4wntaXcMRKPLQFF71R38OLGPRZkxOPV77THdksKiky2t4s/E25g+7qHo5Gr4m32H
PKK8oPJQRO4su9EvfdFEf9JWhRMcA1H6maIxHhzt04nSRRSCINP2fmVLWa6xf7HL
/MvDO6gGsgsXeR7J+qSbbd6vruedRJbOAZsHyfD4cCqQKb9HPnwIHH2qBItXZkoM
CSQOtFF2dByfokUU3447UfOTxGs37vC3HUeezNIRJEqoUrz1axAfN0X4OqA0gIoe
ifdxi6gyGR0V+CSI62evr8pz19JGh6LyohALzALeknJ2YhXUGpWtlP6ElO+IlXnb
JY2RoA6fWaU5f5IenUIr1OQqskjNrditMBunXONYxqyXUirvEUoqfw6EtLsu+rTe
vKzjyGqcplrUUi2TgwDTlx2szn+RVwPX8mumZwIqBchQ8IpSCm/ggKh7QjvqqMc6
yaRcvW4lc++NntOzeophZnpHrGF6zV01F8E7UVHlv6ZC9wwuSNq0N7tvjUyGD4y3
a6iJW4QyRJ7Rr7AU/ONlBq+YKYhiL5/uyiTZQfj7s0xxoYMyB9Fkalq2oyoY5fyh
7W3Ok3byuluZE4c3Rc5t3b+GJfciO4weoYc9V0pOSN6lSSXuLIEbe4EEUsyDDVDo
iuNCruhzlCpMWziV5yw7CfsAd0QHJLem+i/4KJM5XyjJdM1YpUXoIol9Db5FAa21
+V/3ze4Lw6xQQKseqhJjAM5xcfvO+cSiebazO/VUL7ocnRvK11ASNCl0hch7BLw0
N6Vl+WWMxF/aEakVg8MSDsGF0v4Z+PIH2ub0+pvNte1jRROCVhSzdvAfWvdCVdw1
1/sVypNrRMqPydor6e47sCKfFMSJc67s0itOvJiiRpWlXOeLKMKw7lV0zPQVPSVu
l9Nv96S5yVvFg8PcxEnhueqXjvTeUqpdQJNMC04zsI7ugEv0y+bJFD7Bi1hlXi41
aXFgrgBtpijqNkO4AKNnTanhnG/SJFARQ3hqEB67E8Irfuftv8znYUJ1IzfXb+yy
wXRjUxH/RWN1Rfk25l1UcsPzhqNP1Equ3C2qwilJIt6HI5vGWnCUYdYgLCbuGo+l
8ywi4ebM8GYGfV5wx9gnOmVklaOKRauPyP//XsUyNd9UcmOrBpmTwKM7ktNmgosu
XFHIZe89xbzvL8frGg4QlW9YPI1UXGJPKVkpomxmKBh4E0y+KwR3sJnFSMOEL/CA
irJwxPqqGVSCnxJtBsBpmGvvqjgaChzzVIHL0IenELTB+Xss7gKU48w+jyvsx/d4
br/pIurQoYSuhzB77xmI36xWfK6R3ZqTggKaG1gAkw++c1+8QA00rI3zao1/E/QN
+FnjFrJUvcD9vAAiIEHRUi4qTKB8f5xkfR2Ozy+s/lY71V9ZXw15gUpIaDQ7q5fr
RIBGfC287Cy91WOf2nsKdVYlRf9bMBlHsEl36Jg/3WQaVGLGgzHKM0mRgc8hl2BG
4rf2mX+dFxoh+GlBrIQVpG+n5xVdpycyQp0W3s/mR0oZuXgSsQ0ECRHSThnxvs5n
H6GxQIa5GgfptXib323K9WvZYuXytDic9MnCYE5uTTB9KLkjr9uDqBBX7vvBstfv
EcARgcoo8FpoOPaN1z6zTNfVaeJIlLViAwJA6a25XWLSnyH2xrSLm1aMX0dIHQAS
hdDlQx93yk41aT4hOUgbl3qHqKVTJeeyADy4uWA6Twto8Lzp1H3HqEVNQKi9Gbi4
BxU5QQP1fV9suB6S9jvCZHo57NtxINF5wkC+3eLrDvnCmj1B9x8HB/X0ZUA5VbX3
mqDrfgMr43uZNegmciNGwPINHnD/kVDDzFvn5Ut2xNZOxlBIbnal1t/7jaYU5vqp
RweeziKAlKRi3E6hRbx77WOxHclI3+1U8apvjXx/pYgfe6SLUobDRT42Bj6BG82P
erQPQeTo/dek1rII99xg79/R7Msm0TL6MrReYmygfj9bDERr/Wnhtf7Rx2Xy68Q9
ZDK7F4IO5TmE7KVUj5BtZXG+acf+kj6YyHj8pxXwm6hFeIyvWeR5KcDDEtmjNRZE
mAECQVeKb6U3JHTJKNXrfgzC2yvm6kDR0vB2fc0Iv5msNQCGWqS70/ZjWHjj+Jms
UWR89FFBi7rlGunw7OVjt6A7zzywjmIupnEchH7eTe7jfaEmHzFvX7zK2vAqbY4y
VhdwIhPdJfSDG1iijDl22Y/0aMMIttGA3dTZQI4NbBqctjgCwipXNE4U91+Lr6EB
DnSQYjSY1jPdoIHt9f5k8JZ6cTg79cawhOAqtnmdg87V+Lvobumrt/Bqgx6Uk+68
vZiMQCY7ydU+5tkg6Ct6s6yS4gO0zlGmdYFS7Qa4dw/3qoXlh6pi/TaIkQz8hDRT
AsAodZhO52wlwmAioLuQbMYrMvqFgtre7oILu8eK6qgPVwbfXXJ0LiasbJZ0Fu45
eHOedSe3WZ6QMWPrPFPn8bC3SvI7rV1Thiic/8MorjuKmpHpeiMTd0Mb8HRjLWr5
j64ImmEKjVrSRo7kzFh7B/MVzCrXK1Efdi48ub/9RIwf4YFzn6aXWZNu0i61J//2
Xr7SjJcSFoeVN3WRlkreyvjxfnXp+E7I2ks85u4pXFD9SaKl7QoYc5p9f+8qVKds
DlYjX2MqLyl24sMG3ifZu0f+OyEm6y/2Oskh1WVuRQGOSfOJWv+YluSUcJJ6Xwg0
xb0/AG7Fp0P9jvk3pk3NwQzu5ZF+p+TOuRdTjBYHuAcQvG2m+JGKORoV0vbIMQEQ
/+Xrqe9DLdcaJ96WSkn1PRB1DMdokYAQfWUE8ZqRK4eomiK6yMKxXYaBwmfcWlE3
oJ76LnmGOGrr9KPEpu2zqzqrRChaAFzYgAhYLRExVQZh2oRlzNnyVNxYsFBEgmV1
4SDIjmaogzuDZwZyX8UbQeFhBLC6oHv34XOI6GSC3mqgb2prsjFHJFID+s2IVXwK
+She8rKAPaD5jumPCEKjcPkSuIruounYSoZaZ2pqU8MI+fe5kVIfwoWONUCeh8OZ
4eR/8l9PswEaH/W7FrbnsKuL98AeJ0UwwCO+rflxPNxQrO7YnUSwtGf/7K5FaLxL
S/3ITKSCWCcw95hDeXlPY7laqB6G50Jqk6HFckCSEnnpw9XxGBzKN35KZLTvUEJS
p2m+FvEhbW0cXaKxn+jxlE7itO/5VxSF2TRCk0MCXnpfLgcTIZgwdo/pafemQC+N
LIw5I1289YkOwnL1Xnet/nRq76MgsfE7gCtcoFOtrK8KIWS8NS5lsOB5tpvOvbeU
ugaFx5jcpL/SfCJTj5q7Eu7UDkRl0xXLqB948WjkkAgyVsaSBseq1MtrYnzHOdfM
rVNwnhAe69ue+wW+pj3BPCHdu1BsN9EeABGGlqjnXQqiPLXTz1awgWS4TO8y2pbW
fo8FfNX67C7q4xYZOHsimOV62v4aDfEnMa2AMiBK3hBQVKj0GMyd74fEyCLh9Phx
d3nVZlSIjAnJRsB3FbSUndgaw1o6eG8ebL10exZsffPEOOoJi7c1E+Mf2ST3hgZY
JmM5cKraF0/t72nPKHW/N0nG4UGGVIxQ9VTgg7jK9cWdfh2Kj98O3P/W8zJeF72B
RzX7HLNg4FU8I2bcU9Iyy2Uh2w9XyoKxEK13MPyUc3KM94oLuDya4jkA33YBm28s
8HW6ru7WvRDYRi+KSmbHi5roQ8UdOhhTrJnlIxSqrTHhSy0F75865aD1iP726vlN
tU+YqoOGccdGabpo76EC+Dk9tx6Mo04aJshOr/nl0UTWLJlvZpEEOLN+VYmYZIxX
ek041QfZZt959QvV+qkzQZzm6lCWCdcB8MEoAHiK32mlkob9TVjQ00BvoJHJfVzj
yiK4WWPHPwc7vIYbm/jsL8GK4lltr9ZcOyuyS6dNtbgTcUxcdRwaGCpMutVNX3tJ
8VwrEgpxSI1ZjOceMk2W/UiE4751DKSUFucmb3eG9N4bAy3IC+xZcw8CvhCFxC8C
vpxPmHeG5JRGTWbnjpJi0hsPqndt2kQy/nN64QXrMcNkoE0wKDQm2YvvyxjwbX49
LmZN519d1A4XBYbBY8MMnZVq+YWC8EwOwyh1Fe2UN/NS5WkRUIfCfJ5Ot562cwgm
D2JBFqAYrTBc7mQs4RLJFUHlkSI9aB/0LvnBXReiBQuWMsbKcONlDFfYt0zVr+2K
RBZD9cDqoEw3qdyu/b+oW6EVHyQThRbtC90UKcXiqOn3Adw2e81mjVYoe1uVh/36
LJNEamwuLpLbRX/2T+0OpQCGBc2sIBUnzvHml3CTE5PwEZiBemTATHHNrhLUHwoT
AgWi4qzqF9rttTGSHGIp1G0SD9MG3411zFY4Y1yxa5jvD87w+yA2EkOXglqChAOm
UoY6gZhlRPL5afBWK44fqj/Jamc1EMewgY32j6JsJfIrN7grklwLqSno6MM4hH8t
/sixsS+EnKn56ANW5UQqavAy4WbXOl1zsf/wbUWv3ldjmLxwqzm8KaVHGaQGDD/v
mkKtWZV1xXtlxA1tsxCmomUN5TCBs8Z2os1/xs0Fq/+egNtvtt1O/+Q/0BZ2D/CZ
pwGmRDQWmMbmMOeOSwq+i0V8XDeaoU1hY9VT7PGxVgn4KGKAQA35oCECglqMgy6/
MGm9zmnmhbA2Vlr31hxaP3TlCTKXG2J7/LfctBlewqAmxZumqSdA+PDSWlmCtzYV
ugthl9rHjUElVIs+ZnnNmsn66hk98P7Ts8gbyQAVxGFaFGeq2Nv32WJrWtt3GbUn
QpGnwyMzzkzN/KZoPSE6we39z5AlPzYkyisCBdAwl7vJoKe+L3zYh5itViSsirSc
+xaFzYrVZ6/sPK/Nkvtfk+7m2vX1/lKY7EFBbD2drZqZujgrnC+funcIIInuPHZR
xvEB2Pg4xjbBGdlNmrPeDOU+McbeQ7U7YEYxcUub78kJ8UYUTpTW94TK63FC01p4
IIWHlqusObwNQOaAdsDo0cnCiGsTLmD9GyMaw1BoC6wSi3nb+vW4mU6r6bn/ml9Q
5XQTJ1oyGL9B0eoI0bKV7Db7FOc0HVszAZ56NK1q7ESPQ+EE4SIHqdiBBsxt91c2
0HBZrPZHyn3xooThZbBQtYRWrhkW+Zanu1n22iJc1JT2EP+uZYg3OekNc61W7shk
87nYi6G+LAZXdaToUNEa6pHMSYWdxyTXasWD44CzJvrAASlsDUEy4uKvkTeVDRUE
yotAwRM3pCH0IKQQPym0NlPIAhLSAmvbaAt7vPrTnykJj1/VxLVzqakHQKEjXy+z
t4joh7SjHspqdXugI0qy7qe2v6J7iQA4M8nil1D+pHRjFFBhI6TTjJGeqYVKKGgy
w/pcANT179pilDfJs908V72b2qqLZh0JeZ+OezUWzH2VFP062Ih8iykK71RRCMs2
KLL+WPAf4qlLggfVipY9rBqeQMgY2oTahf6w4kc1WRd/VO7FZkrfOPp9VYsu9Soo
xnlGdOQDGTfzOzwx/xZoBu9khvKifg+Xbpi2Rv6RYGbd4p6jRC+qm+7NpcUF1K5l
GoCcEOPeTi9fIq9Zb9aUpPPttFtol55LMqR47zJ9p+lFLWtl41PDfN4ildAJsXjg
R0+xAonkFSD8qn5mFjfd8DXot+KZCL61d+bod4v58+3F/rzA7dWAQWttrRQ51Z5l
s8NctkhZ7ZVpdGlNoEf9v+kSASKaG3e4yMWlrflNsqGtozJk35hMSMkkUIMQeKrP
bDbfvx2VRB0/sllXW8zq8HbLXz1ZbdU5B/snQjzr9icEVtEQN6N2jQ82DosXlMwD
W73cnK/AFeTgJpYX70ZZQFjoDCnkuc4Gp3YnbfEYiW2T+QouIeo7ef3KV0Ksbq94
qEQ5+ZCjS9UP1wEGMAyxRw7thx0jk91WCzBpnuQMbOt/Pb+qlqUSAW5VVUO+BaVT
cad4ehInD6EACnHFI6OxDYY4LIz51XcI4Byo8oQOGBc4ppxB6OqrBv+j/eoRspyu
SMJpahw4a02v2FOwASD+H9qBQjr86phqsaO2tqOAOKQmUWB8ftYL+T+UDAqcmlJM
1PHmg1u7LTme8mXVatuL0Dvi11/MCHtLg84SoqZIWb0gwZB9AJQTBdiIP6uSRtML
kn4xeKGWsFQwNe7LtK5v6gbFr+JAN9oHkFadose0Txh2IFg3B2rLUdOnQDVSWFuD
tMqjz1IqNJpPFwPzTps7gz6Yp+7C4rfv40nzLMUfrk9p4G2zs5lNvWBo2xQgLp27
uwQMw9WK16qfWpYW6l+251gIBU/IBazeMJWRVb/mmvdVLaK/9KLlvWSg3BsanbKT
dlxLsy/Nr95c08Qe9whqL0HUlORm/goTioQvTX2bYn/AFQ2ysdgWipWsRW9ecZLK
0qz2zhFQVZZNrqV4wvlS4kTxhMm2Dyw7HOZ9/g4D3HuOLC8lz8838rxtaaUXdtT8
aJcUm05DsG5EMLFPToyDyct8dyZtFr+xMoT6uzbOKuAT+xuBrzFQovA/sWaYB03e
TFp97YZCF6hFbnPEaAf0sI00bkypsZ54ip/cfpUOx/iDqsxC3FK2MJ1UBk7L3HjE
AGJRrnCtQ+Wd1fF6iVZXkQwScvVjpT956FcCa/hyAZNiAwS6q0SNBN50HdWZr14W
SUyjBabgM27bnmbTbeGCJuPoaUIatyrH2WW1RzCQ6ZdePkyiGgv3csETSSklE5M6
aagLmZ8DPpGakjH1ghufOR0zrfsIIArERHWGHkV5QzonoMvgU/3tf+hKfoxNhMLt
J9CQl/ullrLQxEpuw/IUtoSXrkyyj5+ckxU+cJhSH3YkaK91hsf0OImocr96TUhG
9ufCOUTHxpICallM3gV1L5e279DEVLmo2xJ548Xtz4txzRa3xMtb4zDJPtY2lBqp
nEuCjQc4hQlOptzl0l4mCjcFlkG7z++irlxx+Uop1phU/Ea6avS9S6zVYwchxvFb
WbT4wefRUw03toO4+DCLOY4NHKCp5tVvVeUTL36ztYvkvZ4L5ipGy782y+JM9flV
8PNzOF8hAxtXPI7esCX+kUTsaDydIGEhHUkKBHJ5PDBL5d40i+hcKypNv8/ZtMmP
Fzr1FiD/ur0CzYGtdT9tNW0GTr+rtkrzIKufMnSsVwP8Zs1c91Y83Z+9WFuw9L2J
KgB3X0hfIGBmeH8LsKyZw7ElNBE702/VRHJkCfsT040WZmV9rrbftVBZNjh4A34r
AmgqZTlkJN+2unQ4kKp55bxx9tTEG1RUvLDhSbT+3ZznZjTbUJEz3HF7OWlKRiCc
ZT0T2imn1/G1u3HW0O5JPilNAehKUMOe6Kn+Oi+aHjgl2JiUhkHpnT7qK8Gv/Tbd
1MfWU9Jotb04EOKrPC9DjXQ0r7K5MYqzJHAZPZXbe6Figqc5q/1Atd/NKafcop5o
if6fSsR+2namAwjwAWigpD2VykYcb5+Q8vXTEvp/l89536DPF2pNBsdCkhkRDUYa
pQps5QqFWtphlcsRR9wMrRanG5567vZZcfhRScnIHRzL4mX4C33T0KjPcH2FLr/V
i7FY61miwL/riDvSJDV+QkX9trDQRJfzEGzd8WNqFR2uLuEyzpt8VyVcxYioktWr
cZcmjbftWW/YxzMi1RBKQpggnXdVSMlWT5TtipIHLtST7AfaYpnDRPOYikrY8PVj
tK/IkQC6dIOoapKdSr+59hKFEOuFxYdw5BSO8FkGLo+LpKznyDpGTnUVhzbOlJCc
VrFFhv8m+vcLsCfIsQZPqiw2tE9VitjDe7AQhjnd09I86udB+FhgcoVIMNbZhifs
7Ky7bo6CUhlgnUV/GD/7qldrd7EkEGV0Fl/nwIMS0RRjwDoa2hzqNQNW98lYWiTC
XyNNt4vwOWNNmKKM/y3fb/BJsbkFbsADw8f0d64A7W7fUjbj7hmOwtk0fpdLPqix
rMwVbVVpiOdv3tpd4FDoeQRx2ERQpjFlrb2DRopCqMXV7SBzWrfzwJWXQWewpi0L
9EGGsZ05y0hXKGWZkbyr9D199AYTcbX+OcmwM+t4p4oDd5ClD1cFPOkjDjgzyAJI
u2qI1D1oABbXn/bJ9Wjg26zhIHAOfBVuJE+f05VJXC9YvXDiicIcVtpSiDKP70kU
59YCrOhLtZV4+J3WaaV8NClyOSjF12lJ2cy1vtbuI8TgMeToQQotlQ8pktyldMMi
Fc8u7lRauvNSJnyZGvuCBKllZUFATzEQpkJNdmhJQtKNY9gWbOKrRIUe/PiGp2mg
UJBMQdXvuffs4hPLhk6NHnYB4mzkt1WbBqZQja8Ee0Kyi4aCCiLrkvnw5MRcYgwU
WNs7HwLBZkuJM3EMkTegPxokGomdcTdsolgAz5yQ/gTDsY97fu3GkdfryDUxQxB5
6z6czOe1dm9Qd47YCnVrGvbP5zJD7Aix2xs2ccPlfy4XKWV8go4EKXCQrtv3B+Xi
DaRdWklL0MioK2wwuC6C17nn4V6L0s8cjPHxVThxBNrl359p/olonJCNaFhsIPlq
7Oi5yaTKEKM1l6Frqx74oGzp7pN24NIXDtPQJDhm3NH9CXKwMV3Wq/rb6kTm/gNS
QWxURO8ZIfLqdIt3SvaMPBHSzsDyUfZF+WEH5qhdwyW56OxhT53Ag05ePOMEMS4v
tHJc/cypb/xNQGNCJ14F6bLA/IuHX/qiIhrdK2jAWYqxxow9C4QXhT5v9jJfRtLl
RfTPFnmRuWck1mrekMYgurFm+Ey/KdQvCMDSghsrO9zqXhCfwDt4avk0rOKE5HTf
5nViqZBVM1KFgCU1n07D4dtdjqdShZ4agSoiReip/bPRMHj74BWBgS8TYFu5U6xG
SI06BbJDOufZfedvIy8YcemIjxJPYGKxfbM33zrLdRnxlmrYOcjmvfZ9BXegkO++
tGpMrYel6axZC5nYbe+6lI3wjMEQi6bNVzZPGfQG9U1vrdFNO6e94ubm6Gv3bA/1
J+Q/Rvjfe1tkFJF6gn8Sp4V4YDin482NK56EGTJ6016ctt8G9Ha78HsqctcI1JhZ
V6USlyP64Z1qHWz92bEAXN8aL96QvX5xNAIbdh3wi48YXXyHdV2yjm+fei7xCNko
JL8mugRmS7WJCgMd93aU6px9TYf1W5sfMFnL78s11I/k57DmqISahAsh2reKnGhX
rwyFhd2hVKGuHQtu4CiHRLwUC820NBPsn7tzsjTalQjDfaiXVqRwgYh/+xYwaVB6
JQLaGC5RcdoXVR4R0tpZWcxbHe4FzJjCezaiHuptgwszT782J4GUqKLCpN3d6ccU
zdTztUpqHZwbnYuk5s4PjVpOp23czyZ4rUL7LZMVzLLvC7WN7S7VM2TGZDNhmx31
AsAT/3z7m/U6hqRj1OkiQ3GMkJ1D/u0HTns5yjzsZm9EHcVLrR1EDz+1vy4Wtacq
QT8nO3rekhH+5j2RMnR4mJ4VdAdDnMJWLEIUVhcaSY7l0qPjQW0chZ7kgH9GVNmi
A5HojGmERvCzweL64gKEJX3EDj2EthAhuyLDo/rqSNY92H8vBpK1TKrhO+a3Sknt
TYOpw9qRVgAg3xoIHY9jXTKHUWs3wvQwBHxJDvR+02njqscRkebLI1zbfIJIiBgQ
dn+/lM8G6iCV0odHoqFTKXKsEA54Ikg005Wc4eNGHioPyQsKtKjLkaJaM79Fhvlg
+NIlWox/EZ8C+Sa+G1/k/yMJ5D2xfFQx9T6k24WvMrPcbFK0gchtrKNQu+lu3Yxs
maPIw5lIy99ErfBxAyFUllTPxV3N/jPJMErLyOh7D3KTSgKXSey0XmB8/EE3DDTx
dYiEIyqnNUsjVb1S/0ZsZjKTHfQqh/kQ58/aExzuTvZhXMcsG7kDs8pYSRJqwgWU
5WRZiOJTiMKWZ38/IX+2EYs5d150XpMvOxKpK5wrUNPD8HxBNJURkuF8GO43uV2K
QfuEfvM18o/DGj5JHIbxyiKppH/byjNi20DC6bvsh4a5EgomBzOO+rQJ+127YQWc
j7ZbaOcPKjZj9TEscfBMX0znm5P+dgImpeKe/MQa7z5OfMDM/8uXmQwzdbSRR0i2
3jIG6zGFmNGez7rnbwQgg+3K1rArDwir41WDgR/AwschD1a/3RV7CQImUyKof1vB
lPpX1qZ717+1gNQzjq2Cu702TyvUagOEUvbqZKYpcLYXMxiKC72U3M7vFcTrk9bY
XdQk/FZKBpfd8EkKvm9CQZj9xDjydBaK5T7px9wqZ/qj11QL7XlW+rHUh5WDlh5b
OE/93tyXqk2lLfYabBHloKdXJhmUEDRa/wVeYZllwMgSYuDLYOa4yuDiuG6XqpNm
IRczIiYu6fEN4jxBU7dIGv4YsD1DEyZZdrnTCXO0f5zdRQr0CB16tb+Sxa3GoO3X
EFYOCI42gFYDA//pPoR2H4uWXZwWb9ZARoofU2FNZiuR+lcipqEC1c9G5qduZ23W
loKjCdI4jprR0rxWZ99WYvmvhuK9wYAVoZCJw4VRr/UlvlazeP7SHMNUXST7+U+M
lp0aCKLA41b/8wQrP9bzQbuRpYlwe3LYVKjC8lHx17+ui3TqZYJybnXnpw7v9LDd
hWm8uqR0//agMDlb33XAHxIlDajSELRGHpfS58QBok+hnc83Lt1AjOuzi/RkCYqJ
e7hfjetMSOXvcKYfvef3ykq1P6qL5O/jkDWO6kHAcY14zx4jKgOdRclqqznLV9Dg
n7J8dSCfDAmtGOYPK//9niEVHgf4H8t8TLcC2GYjzRxyjn1eOAvrYV9x6r0PChYW
biKiwVDDYvBvuH+rMT1UM+6UG5s+DLK4RB+eoVmi0c1xKWMofcswaa1VgeFOz1mb
NbpHJnP4ekgyGk+fVZA5P1z1GeIMx9zsOTJBCG5XSt/B5YEm2iCA2IBCcXurkw6Y
PckqNE6qL7kYRX/YEaXiWuLzs8EKqb/sRAveqk01/9TsJW9eM+TwGunzapKnph/a
niU7v3KA2BanoCNeQOdfAw4liUffvIV6hGSzOTcqTPToz1lLYOoYXmhsURT3BICt
gc5dHm/mQKFVOdvnYWEG4rjNko/X4K43dYIR4guigyEMdYby8cAILE8FOIJbqIx1
iTjPaIS13oGH2vcz4x1MvCfybY0h+qMRjiNwlwlYiCFJZKTuTXpySRW+MC1giBNa
1DAl/GhWM2vZMB9HwYgTi9u/TfTAxuggFrSOVLlxlZTLDyQ1JeN+z2yZehG2WZLD
fBtf+2pFWhMvGGshP1JbOAZnBNu5JtuErS6tuKoxF9Db6vhECDFwueUsddehTvP/
6kN8sQJ6uwP+dHG0m4yX8RDh9pAsKBf/ClT34V974+jLWcnEc+tSvE2iJWpYD/ul
n3Uw5KWqG8ARqc9xtuxFHBs8Rj4s8+Hzx7V+3WuTO9F3iVJnnEli6cwJEBTAydn4
xawRyJ1C8hZeYAp8UyH07TKkQy6UcGaN49DhYdbTFblLeP+KyMJYj97r0Nfh0VZ+
ua9IjoD6puyq2PQVA5IjwjBH/d6j2vUQOc83QJd6OaHom+nZ1s5M6XNGPBDgNbkh
30nomAIzhf49zoY0IbIi4dCJCSIcX3ql+coH0GesUCYwDBNBRnrzkjsT5gAB0jeH
LDvMyCZdIQC/8kYE+XAenoDPpYEnPnOkDKNYNBjt+bvsRqHL3SSrkSQUT4pRwOr4
Ov4Dytp57Xb0Z1YzhM9nViLKLPfdp3l8bu5w/MzJL+ybcscjkW3QEBIsC3sRxVYW
bPJDlTJj7L9vMnl4kCB6FCnO7TNY1VemWElZVa1K8OHeQAIfIzwYa+17pEzCMOCN
Tq10x2fvoMX9CSlt3tW8bHt6NY6ytNVRc0Th2AQKeLgbPZzubBmoAH6AszP5d1DQ
2953kVA5Pjd6oRHcbQTHIKs65I4LaCNlP6CDuJPRQtTRilkS1ATxKB4JZMTEylen
ITj5TluHwoODmPwu6Yu2ODJqvUb6NxQyEQ0/LcvvDwHYCJUcbxTLtUZM+Nw6XOxT
X1lC7AjyeJKfTxdXKsRi7wsUHZyntdaSM7bgfeFHdJiTW8ochleKkLd0uebprDOD
5Bn1Ettyl4NThEiQhWdojSn7kICHc1gMzPrWopgbAWKCTfYFnBelsgpxMwqIW0qd
lGgyOia3KCujWn7jVyy6B2X3VCOkwhHlGoQ0MKPhXQ48vGaiq8+JioVFIZC3Wx5a
lk9DnN0pRoPr/EGJ53B32K6aEdJNxQJojQxW18Dsp+mgPTehlTKec6aTr/JYIbgP
3IH8z2WZ7WNhBql/bJLGG7XiMJeYhuFC6WwlGW+YnK05rPxgvOAOSFvcgPe+ctHc
nVw9wpa6nl4v1gXdBpaywhu8+fdWN1Te7o2l0GFWtDCemnH2JPpKjUEeMX0hTsCL
XOSpxADVjmkEnEGE820rW84PdvP6Ge61FuM6PU4nubjB9Kxl8cIVy1tWJds8ECvX
c7NdncSuGQbepiJ/oUdZ1J2Vrcqys1h9w9QgbSqgB85R8+xbwbxa5JgFJ9lbjRut
rfYhWBfnzVf49xHkimckR3peUp0BByELCezmYdEDyhgY4ivfQTcJ0w0LGz911UCr
0tcOPedVd47UcKeVo1F/x1n3Z6Q0DIcTW0fHrYTgspgwP5in7QMRQ9uBiD4VXjxG
zlszxlQDPLRTxPuOhmoHG5EQN6FhRa9Io3oSSwikdH+7cSGVZN5+sLY3K1ykfLD+
nDCtBIGW4icwNxdp2m5vFm6G7LUpY3mwaLkQ4grB3EA1Mwi+BaKWNp3IdJzfMEZr
dFnWvNX8gJUgmeo2aljSJFSZ2rVpgyM6Q5DnlvnW5WRoCBicbe7Q76ZwboB9A8ry
ou2UhQ8x3QufeckHLnJBtbzKvwfhbPIxjR2QIdg+sr5LvPLWsGs+PvCrtmK+HwWJ
bHs/JDmg2kL4Al5pBQrZLNaWaCDsy9zp3/dmfMNzaxzo2SClNwDx3PAIOqI5M0Pt
L473a1VzN/OxSWB7DJHvkYiirIr4/FXPXHDoV8cqaHIX/L2mhNvJXh+wNAFLT+yl
6xi0l2DPVUfuu+uol8Oi//lvgYF3lr1A4q0BGAJDYb92unjjsCEWKjfeYEtcpfsy
sVmrxlR+f/Qj2ITVWQ/JHormrXNYi0s8R7NR8qadSCUhIfaXFQ86101t+I4FtjOU
tP/Bdb4DkH1C/fGtY2Q5wq/OOvozfEzK5vWAUSATPr8jPLMPwM61v2b4lmHNZuHo
w6M/R1G8TGYS0UBJGxggXyF7M9/6LWLjGeNNwwfWDnrf8r5fPDZ2quMyAkMMn1Fq
mhpC80vPIoDAoMiUYyAKBuEZtDPK/ZR44KJ63Up028UYR6iRFmBpruBSchijLW9T
eQDx1CArHl5kcbQj8AL34SBKmCfwDknW44BbmqgqQ30OU4EzsMx7sXEI2IuOfKV9
ndKPSgX3Nf9Udcm9d+lEb4ihZuJw+5H575qLg2fMjlFIIq70wCeVPbIDGXqoYdWa
GstQGAye6bExVU+8wgFUFd8JbDKdDAhAj42lJu+6NYGlrK2i9UWK0M4HBFZ+8KWq
uBDWJw81W3NyK0bu0T/qoGPK57C6IHopDPcVIgnh00ULgOURrjPUqACd+23qVm1M
qdkRjhJjArrog6koFRmzUsxHdGdRl3d2sDMGh9iuzWq2W7j14awQhhlUKqoCNO0p
C/I4UyH8k71NOiXYx08NNZKoPIkBAWde91TbFPiNOCIRlFH/VfZFqWotTYsqMPQt
Ltkx31e+mZO5RypBk4zolrSAu7aTaHGSXDZEJ93rCj3fesUM50e7s+Warhqjt0U2
KnvT2yYwbOrXg9iW6Hd/mw5qGP+U7hW8L17cVbPHRM+tTYoDX3bQmrBnTxdQpU8I
oKESQMJdrCq7ddS+UCxCmakrEhoZeer40BxfAxo5vphWdKjhxn1+FJ9/z6ybSCQn
s5+1y2R1vf/+tOkvAnRaJ36AWJkF4kwrkcT7dwKm9j56jbON22v2umy1XxUDRHFf
enOZNXG2Icnpvma9h/qpayA+ez+nO5gPZ7GkWzaSza8RpDwtFYl5bdawCiyo8aOG
puWrOY94ZPhnSmnKMDk3xAJuMvphdT9pz/nyzfPVn400GTZ3yRe8w1RADaDcKnY2
BpDUBPwvCvl6JO//b14AqgaqhWbpazmlw1NGUCgxswY4NTs2TpucPC2HbXVJ2G9M
eFlAXtC4114ErNXqrEDtWJDC0GtotcLbDSwf7ZxgCX8cMDOSNmzQjXAJJCe5he/k
/faMAbrJa/cipNm5ejZi9BAWsED2mpaUGVyEEzLhYVGoLmCkjKxFeD+FlCT6Nygo
H15RNlY1AX8esrEG03zJ4moLTC272dWD574h0uMmDpmMiWH/oVVSL6LrFju5Wmec
HFiOgCiJUIcfFeXP8DK1wsIhR29N1JEuhmMhJe9QNMHIv+nZzYUtl+eC7XONn9KM
hBsmpkIvkfuDQcxSsGxKOuopyvqfAESmnbuco7gn0TnOhi3t7quee4F9K049OwR6
9XizBE6UMpKy/hP6MeHI9K+iEnENumDnuE1dv1C6xECMGiUxoPvIcYjIG66tTVwT
7vRlSq9r2W6XlelSXs2RGNOwnYIfd35kNJsG+vmlT91ybPwunSoVrIyPQX1i9Heb
xM1tkXJBfnAaUrCyySqPAE+lJkW4WsaLHfnHvCrlJMhb67bRg6fnhqqvxdYCgfwz
aLon4/Y0KbLLn32Kvemi+6r/tAc18483IHVNPeij0DL3wJOd4FkJB+A2oXh5wJiW
mNnlnJ9HRxNB80I14/6Mia36Kz8WlEChIaz0jHcf0EWXBLIqewy5Ci3+pGdSlcNE
SASYeOxR0wYARcA9qDzpbWVojIpV0bgoukeN7GLD7n9InNvMV642BN9dPYIGC+kY
qK6ZME/Vbe4jtrIpR0E++k/udvGovReXpoGqUtbFZKYGOIksECf/Za+2y2h8hDPX
UmMgy6j6YXuWGqpDc8tFbhtFwngUuu3xWqYlHT0GlFj6CibOMR3dTJSEOMioMc+g
nt7gMoyLCxeiSCkt1Wcut5ztZ9IGYx7NIdE0bZC/BmNEHKZ+p3c21+VINrWfS4cC
P3234Ny5a9sF8hlGL3lBJ3QGs9Piq7QWHUvCz48w09l2NQHlYi3LEy8KUUXi+X3V
gBUECIkHPhqoxNVflWJvd6XFIO7ZLQho5TXHlTl5XkqWguRX0cpD0XYT48lJYZgq
AvHLkwBx3u+1wb3vRpXbRxCu407l/yrqomOwSjS8g1T7gHHGxF4EZDmnb4+dSmNX
HsIk9NQ+xC4TSHHVrjghv54dqy9jhiTlsOi3C2DADpRA4hn9GfcIirZMsqa5lcm5
CPsXa9E+myD6f9aYP3DVj4p3AnUZmQsTbus61QoqW586B1xxgTwZCs6AhRg10OnH
WGr9D9kaiBMBGpMsW7cXuc0XScVTwHuU8c3G4KNEyCyFcnsBtblCRrrf+J2tyZEv
QGHj8O6e8WLDnK+KTo5KmeGYhS2sHtN4310+6byYK7t2C5IdcdlumZO4kIK8tUYz
4nnp0yHOTojoKSIbKNcuP7rOpNxqthhH+GQCNaHf2cjj3FT+Ux22jGfRvKpJ+XZm
2v3BgQyo/TiigUNdjvVQhJnSXBkP7wU8OvvAMZP0kbigiPvNytrF/OxWBughVwrM
erb5Xunhp0aEyqYe03Yo7pGSqPW8iIeF1wns/dlp2Pz5vEQZ/3aCEsckXYCq/Bvb
8/StFYjFbo19lTkeSDoRhp9OgoRM16CfwG28rIy4GKnYksyuBmy9Jvteb7X9gKlG
u5sdTGlHJ5vgdxi6CkIMVBmc92vE8GYOo6SnVMa8hgvEB04ySUXW3uX/OqdIae8Q
jYoxXfV/23C+jKYSkqtDRHk3/uYTGS4uWhgzpd6dUj01JAxDJ5XdK6lbcZZTRUOJ
oi0Puyav/HGMiYPJ6Nrqm2LtrvTqllxli86rjIS1z9e0Bc1gGfEuxNk4/bmWdyB9
jRTiucjZ+jLWhAN1Eg1KR1/oXEXZHBYzcK5MGqBbZWNFUfMIgxNAcql1gLx4Fd3n
Wq9TDlVKbxPBgquT+rT15YFn7sBLYT1pM0GszkDahyuXqVJ0qeLUZ8AQn0un+kaK
xc6lIskDrkDy1ks6bEsOn6eADtCr8TRcdfQyrjupjSuXuFWh/+ys4TQUCSm838ib
pd3SwcvHTI+gv9lA5Ze0qCKwRSESih03j2TlcGpXqJAGtxKi0z/uaorCdMeXoKGu
SeiGOjpd/D+Abr/lkZV20FsrnNhVO+VUgmDdKW+sXc4PsbgrGlux2cGNRpMSTMyZ
upqUEcZ2UcP40XVevJzjrdMo7URhGXxaGL+339T0+DhGomecPbG8an1Yx2KeVmHi
EIy2eTBRMB0OEj0lK+XIHKnbjtrCBPKVBgzUtZajG3XrZc9kvTbfamFb7kzrg+FU
TaOxtFfuzNVT7/qwoXpi3lhhPrxKKaa/8kj4lfvkDZU2eDyFxNp3wa72FrMQzzwk
5qgGtuY0xlrDk9oWYpeHH8j5EpQIkEDFMejNo3ODEhEaa3xHH7xz22z5OXD2NX2r
DITdMB49A0rqKVxIw/tCLY9ODEqBHElPc2cyGAvVuabp1gDs5Vl4ww1SeO6FINnQ
QZw7DdTvGW2XTQHeMkF2pXIwUi8Sfzc2Q+gCtJjemys/glrGQ/UgdHRpMcU14eVD
KyAneN+bUXC3YwAAEFV7xF8OGWR2MtyGHu27NEAJIQBLcuTU6A+z009P/hGwyTT/
JYzZRoanu25xYREkLg7TDQO8+bqDjfd7Smg1BYCuFRa9lbuVjlWfc9+Cn9TsIRSH
LuaiO5it3T58+uxvnjxT94y9WLXh4SGzWOMXl3KiRTRFNk6pwYZ8L+ShR1MNIuG5
83K6WXjuHbfp3Ex3Sx8PajmR73w5nbAXj5Mu1yoHtJDY/a796T64wYh/wTQY+2TW
NoxW/MNdAAgcl6Qn3EFz+IlmhnjgjpM1K4tYPggF8sCR9BXGb7UU1hhluNRGdoA6
MexVRoB2OAwvfvVrqMsZJThhsROmQOqwJWwMYeLY2BMw3AQx5ibz2/wxV2dZyrUO
glWZgop8VfkhIQ6kbwbzUratys3v30l+xIhQZ7d04b3QasrP9Rd7c4r9s/jZq8hj
950okaqS25smNUgjsJ5CfK/IvBC7NiUJxz++Jr9Ft2wqXVUJvWfmXC16jtF+Kzjh
Bnuu+hNu5BofyOv2ZGdRuSN9rrodeXMKuwX9EWIrnzTuIOutBKFX3/dxR8gia8OG
tVvc69nZOJwx+5FRw7Y5zBl4jR/+2+EqXPIqtE3OK32Yuexy1ZfNsRHlSmxF5C39
eQjp/6a+tNTCpq3m5iEtkVpKN+sPzEDsbtaMCKLWfaPo90V5575R9qUw0AGpLi7q
kz0YMHnrs7tOf8b5Kb5qH98KgIoewp0IlJWoFdNUH+4sxmJDIHeEHGPhhXM4dBM2
5/MDBUD6KiVS5JJnNhm3HHtF8vamlCv1bI2IDYaHWdkb1Bhpij2JVQ8khFGhBugY
jnT+ZVTIekNcWBCpt4jYGEBIE+i1PJCVWehppyChdoZlKmXJt/oGFPhDdbzHLa+n
2YBAAlSxcRKS2vwRPC76aacyktfzpetHnjxkkF4BzjJwtWg3MxtoYCn82GVl9jtu
BOg+wocNHMZoLb8BgWAQsw4rWc47oh0fBunfkp8o+0S1uNLdU3LVG7YnHCsJuq+h
yeTPCV+CTI0F7V95HEmKPkHpCOWMbSCog4k4JZ3+O2vSmJuRpQUXJkYDtvk3fAf4
ykW+PtzYHyv6HG5eY9zVUVRs4Tdfe33twz26zyS5Tvf+5UbJtk6SjQyR408/b/Nx
oFJm+J63bAotqByTmrZKUPxzACIWRiEI4kJ/ZbxMFgfQ+mXBYDZXzYrijy1DC13t
JZNJiI1qKc12iq72+970GLHzWJi0+W1v4k0sYtxUmP0iOHMa3R2asZkAHUsHMG4R
nQ5w49IsHqXB9jgsjSHgw8ANP5g9zgdIR7Nf+HvAv8RsaCyYRc3Z8gxLmEIyb9yd
Kjg0QGngRQsWZ87m9tgRxQQaMIVQgiK5ikCaS4OUWiOufsTrrITlwXKge5MnGMeh
J8BvSwrVNSJPw+5qwJ5mG7BDhYHtJD9iXuPj8kxNUMPvewmoGCQyoLOb9dVla1BK
4pQAeUoe0WYNwJjPQcf+AN/dO3435iCMYKn3KngRhB06BcRobv7Pz8p1GH9LJGT7
FFvTB9TyHfZPbRIrg5rbU3g6j0rS9R7vKK1zd6NPvRwy5k7Vp+dK0y/CfMPqgZTt
TJdjBmsIUKZfuXFLq1mZZUAfmeGQEnyr1MDSM6zAIDLdHbKUlNZWIg0IIggKirPc
UUjvmZyBzmNwk+AzOtyrJfK68vdsZO0Rue3NbFstXyg+4VkggswvNC7++7zF9ZiI
Spr94hrMzFG2PcUFQSpEO2qyjXEDusAj1l1FleXIh/Sxsw8Vr9zvLR8kussng43L
VSrwrkokpvrpiTYZB1txRyyV9oM6maCL1dt75tqunXLN2sD6iH/+VKkQ6UVorhIK
F3954lsuavYS5hnlJJsKNnNtGK0la8ei+RRXirR+X3dtI1kwDrrupTl8Ki+3PigL
7Qp9OUxG0PL2B9269BPnMDeUlHgvJUeV0cW4VQL6DjV8spbo3CgB4xw66zcLKlzV
LzuXq/8SmNaGMK9kS3U3EFlAdV7T9BZKlMoosQ7B5Pp3ZJ1EpgpATeWfQaqxPT+8
syR8oDiNNKAeFs+yJoVtJX1u/oXlckytLYno51SQoCs/oA1OJF7cTbzZ/QOQE3/H
S3Wp0ysn+a+a71u7+TOPRI3cP8brylHaPWvgw/u1TjEs28ScruS5Dscns8BgGepC
lmMWSnnShqbbtjuwGF/rxy7O839TTQrTdWFUKOAsFcydtJ3iZ0+i0/EJe3VAal6h
JexT7PqLCYfEqoWWQzogScsxthD3nE42oUM5/cT/fPvSPODaE0/I/8OI4OrMmpSJ
TLyik/bd9GQRZdTgAceHVEg9fNUI6sEs/TAgyfVo0RWGTT5NMVO4jI/reQs6MDZD
8GX26uGyT4sCkeMHEpR7qBtcog4TL2LRrykklHaSidiT1ybHieEl5Eebgceai281
3oUmSGp8wwNCoXhOnLA3D8S3Pp4YHcDDZd7c+Yc6JJyHrmEALR3O0rF2C56xQOds
9joPQZXWdS62++rm3GyojxukkIIL7YiBl63PNjn8mLi23+u2tztUwRGKk2/7vTJQ
DBz3xSZXd+f1HJ5DTKN1Pb7ijPrCJ1zaxiEnrjei/r7HUC+srpKZ8TK0pj2FBHCk
f7mJHBR9BjP62JS8jhKGOXB+Kg/GFnUvvPrd01ocgQbgj0/wd/Ta0l3c2Oif+W5Z
qPbYHeriQ3eOQGeGmtWQdaVVB06pCCRV8PLljdr4Z0FQi/AymV1jHTmO3vqhR/UG
0A+X9ET/JuIEu9AAu8XkUH2dmqcJx9cslofNJ0o9jI4e/29p5/aPU7Xo1Yrb4ty6
JhgmL6WnP1ocbV1yKpWJ8a85R1Wi5Jq2IlVcWoluLLwcdAd87TpAUJxpNEHzRTFn
X+HRgcwkVZwSybxK+WM9xOzb5ux66thFFOR3ZtuuAYeuvNHoGfpkjmnPw9wkGelz
d2hWeDpfA6c3+5OG+2dXn907xdAgZ4AGeVhwRjqd6qT04YgWJOQU9eZTglOFG7wR
ff2ekMZhmQw0opH8KVTejqEUlfVAd6Msiac6g61EXlGe2/AWYlKTSfxR1JlwMi7K
D/94FfdnmxSGKpqjuDvXO5bULypY0ozI4JEC2IkkNSYkKUUqDLNQeYTBpskTINWg
veggt3eGgDXxggV7HM0JcLHEr1mtK9i06qvH9BdJ+9lwovphn7gJkNLl99BG8DtA
qB4iG8olnm2gyR9p49WOizyt5Jle4yCuP4z0wcxP3Up7hlmmD8T/GAy8HuyH+cz8
qtKdKKk+VlPK/jiyeAbKg2n40erZS1zGMBtb3GBTbh78ClZqUZN1hLkXT9rM7Ura
7KxRDF7oEwkHJyvmordQcO8SwJ1195QesKqGEe7IN2QO6+5B9rP2/QzPcAjFFYXr
8f3XGE+gNF5riqoNVhRqFUk4BhLQVn43+1x2KN2bh/zArRRSvW6rsemjIdC1ahOZ
FNtg36ZWYqs5ZdaBXTnfk+0F9dyokH0mjAq1dOXgG1ZEP7z+/RCHDFIlGnUPbx2Z
NWvJtunZC5MU8a+ycaY8FaPW7CQ8xGoD3roNPK1WGVqccfCW02D+t+QPgoYSdx8K
p/TfxS+JFGGwX5Gi1zBEBpop8rYM4FMzLqrOhoHhNClvLkDtMdVFekF67hRu0nRH
o1VLXU++BcWVzH/1azvMQX0I2VuWi9qPAbGaV4/I9DsiXmefiYuqly/fStDOiL9Q
KQ2Rp/TGrxptrp+N5K1rw6rnPPUaUdPlCeacVVYHZDckBZgjJ1DmWMFmGOQzgNfB
WxtWOsyBKtveCeeAuUOt8uvKYMNU1p5hXaI+onrEmUYVNBcUSUaKsznIyvodqKOk
qQ5O6MRBY2/msP4uS5mLtFZKh5tJrD6Lh/fPq+jDloh4YbD65IVcJnVfYSPK7b8l
0r9+DZ+1zmg3nWty110rV1Nj4l+87slINcb4VCzpnHby4ZSzaIuGT3n+5kN/qOCT
+yQwSMPeTEF9D0Yao8r+K9W0HzpBl6zc8s8IHdDYS0vL8ch8H8LRgMndOb8CzHrL
aHSDzDvG+JLc29Xd92EeXjhGo4TDeQyru/cIv54gcezL65W5jNFb4g0GJG+vOKRD
Q65eNo0+ZxT08Yv1T+Qv2C81c0VB+ZZfr1J/ot8xVCMhUaqZ8VYbKM+QiY7Pnlb6
xSdv8zobIyi5djCiQLqJQCJUD4ig7YeSjAgGIgwS7BH3rwjoY46ex7Z3tV6nMIvv
6PnHm/5IpiRn1yRdTkBMzzBTZ3T0uY89R0HRO3xPeIN82z0kPlp/2B+gkpTZBgvM
RLP4K5K+YFZOMg2jkSRtI9qZ3A8aGhnbUs/q4k0+ChFMgG70NbKB3SxYAH5bY9IB
/eqWRjioLDw2yR625AL5+bW0bz5IbqJoLAo4xv52NiJJAFfOoRJjqrdb3UVDeC1V
wDUcfi9WQRSyfXV5UHVaoQmBnhqbHPoDVxk+UQXHhuYR/3SYUxHx9cJBzhOCIm5V
/XdqhVDfpuzJm/VCpTOlkeKRXxRtlVLzZqi3N4h94nuQqgrUlikYafGtLfpEkJ7S
3zQs189KA6ikhtnG11+Ma62hm+ENdujWoiS35MX07BYJhiWQoCcQp/5cnigSdQ3J
jB3YZRRo+8JDFbKCJ8KrOvUBQLtu71EMVbLkMy9pMQtDlJ3G0ee5kWb71GRBWCIp
0CsMER1eWXWw88uaQhMViqM6u+gu/ht2IHLx3fK5YxEbffIZvhysKHHPQanlsN9F
7z9jwua4O5viN324TuLeKOpZp3L6jx6OUmyCvpBpOhC2qe0p5HJ4zwt+jyKKfiwo
Zsmz5fVcQr5VmTMuQvND97XczErzmi3UnokLw6J1WTZCUmGbuBvUPuBbUqK6k1Rn
2mfjJ1aXeRXaido3Qh/GPevx0YCPoePwO7F3cEbxH2c3vBZv2r7aIbNM3cwFRN48
Ql01bCy8U7Rl+s7y0pNxMIl62r7arBnatPse/qK1fz4h9pSbpkif32ej2ESdZgrI
wNik5iDjOZsxN04H+6BL9hJZR/8HtD1MVL4DFRWtw7G21c5Ie/EX+OJOhguVq04S
bxBnHv97n4jYxiGAksgouU0l4/0S9Bi12TMsOWWqJn2l4/bx6Hc6Y3tWA4YDCslo
EnUoj4ziF+LR4/5F571BOZ3/+r2B4bpukD/V7lfYSiA=
`pragma protect end_protected
