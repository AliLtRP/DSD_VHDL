library verilog;
use verilog.vl_types.all;
entity two_vlg_vec_tst is
end two_vlg_vec_tst;
