// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QfFqkxiu3lv/gYfa52EEYInX3anUzZq/N9qmABQ5lcYVgLpk9D0f8p7XtNdaYOYw
7VSzSv7/jITeFGxXsn8dX8hxzwkMyu59re2fqGcMEwoR9rhXalTZUHTlKEE7DJT8
A4JEZ+ElnIL2d6xWM1xbTEYNZ7Bs2MKJZnK4UppktAU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10064)
4BO+O6LQ7JbNrrkVtTwGVEaq/PIBgdemES6ix1G3ukcrypkYdWD7qRBUzTzdoe8v
c/sLZrehSUGH/qLNhEgd7ygOf4Ju6KHrPauVJjIakS8ivRveepQ9Px1gRoIODj02
nHeqQPL0jWyhYT3yB9SL1dhbjPt90zcJoqhU20FkpBpWqXq79MhkPpDPXjoaOj9D
DZu+YFxFmB53WEiD7L/dVw0kk4O+kXr7qBYg4ciNa4ir1HDOsGVP4K49x9Jtr0gi
IBkJ+R5U2U+OItJS6RmEdAc29dHymUavVXROB+PV9JhFPpxj8EQYzdz5x3C1RmTj
nMOoViHQxgFOkxbrsaQwuCFvLW484MBhfHzlp/ujAHDTDpcW+PCDudqDQ6NMrm4S
kHGCcSt2zjdOrdoeuTxjHxKF5ap+ZhO9oImp7qOJYApkUeLV62qJo4NPMnpQZTTv
GTKe84mnnfWrrYH8nZrmuSU8JOthRODwLNvPOpAmMY8uMtMAXHp7K9SQHgdoZa8v
D3yKriFKZnjZp8FcWbek7tjRVwW9Ml6CxVviHpRRZ9g09QSqQNqvuTUBqrMJgfzS
1+22sDJfzwXo34KMUl/BhY6bJncFM+8lzAfV63tZcqeYPjLJr51DO5bZi51HdBkl
WXCGxfiFmPgvilbiyK748MJ5XzHe/VDspgwUdYcV7WjQujm0habwADKamuAvtdez
OarihL1PyJ+6MASc0CKmUy9XLpvVmOrMufTOFP3S/xOOGu5y71UmIUHvChfbetXz
xyqQe1na1Vrv7S1KJTXkr3XAZhiJjnfM9kGG4yeVVwvJ5TB0GBgE/RNCCPelEQc2
yVnbEWbptIjlmfzsFBf/f0xt8R+cdXalunxCpDvMp5M0k3Sxcvnmj3qRtLoUW5sR
jC+DMpubznMJhKoXlRRODPwObOr0m7rC0TwVZUfPHCiTx8cTqVt53/+VEdUvPOJS
+RD6sVK42Af03eiy9i76qY7m6Q5d029whPquKjnFy/Xu+px26nmVLRhXH3mf96P9
bHqydnto6Ivkyh6qDExKriouui62YWHn8qmgrDmddcgtUuuln8cmymHYliuMtDPE
eExzuY0SZHVvYrypLELwXPsT3qV35s2UKyx5qTd7WBYVGnJoHHU1RY9q/uVj8Gu4
Z4yDnIBodRrOaYNgtbw7nSChETax1VRL1RxlppLGriQycbFz8+xcVtY7jt/eDng3
EVogDs4FxJ1TctRrLJD4nhQbju4u5PZY39GzYFqfAkvBMgTUeLWE9Ff8fI6QiPay
MRQD2X7NkIf0PruLlQKh/bDexWXYN11RuZ0OGVb2/M7pVgjdiawpqoXuk1KPques
q6ZQvjj1kPe1zrh6DFLJphO+ud5AsTgqMS8U/CXJ7sFTwy9xJw8IzV+p/b1jaawT
yxYPDMSy4JMJ1UoJ3LC81f6BtbLvRp+8Wcd0MzEezVUw/eXJwO5ogtLnlSzGVHhw
JOF5tDFcOZJgZmYiFErJ02L507ebjHgx/s6fkFTW4nIu8bXToNWID9/V3D8iO1Tc
UebRxEym1qxWjlHhfUxMiZtRxzhI8Ad63pqfphnqN2QZM3PChmCQBvy9ChXl2O+f
A9Olc79pyBDxhaUidHJfiScjq+B0bGLFEmPuzbs5ebbfIkshAa9+KIWOZRduXkkB
rv9CHmrIhIoC9pgNoaF43RfIxjro08RCXjdCa6dY3Dua9fLdnBIAgtfr8k6sab4F
tBLNXUxsI09LMI6k+9e+gLnjVyChA72f9FR275tH4RiKJbMugr4Vkq070AsC2NwD
jjwerufrETJFVQ+IUtmYQtU5Rg4gur31wcRyLbFuEHSv3bKw+aBcbY4vEidjwyfI
vHvnXyHN4JCvSvTCKXY1YgTSnH8cq8RlDGjsT779EkwAq4uboNWKEq42bvwkpWnq
Xs4kdnERUIfwLwh/ZQMyW2tka3tOUQ0OkX1SVtemNCidMCoeqFhkClV8atMJ+e28
UPa5nAZDhy2cPaq1S+4QhEvI5UDBt9u9SGHuQ95nBRC5wnZseVFielSJpT2AZslz
/fpJRU2LVvc+Fd87f2segRO8N3ElEdx4/qKRYwAvX98tX5heFYRQGLA3ghCMTJne
t82Zg/Zt0gHZOj6U4IrQdzqZtJGlAujl50AX42FvDnT6befEofM1BG49+J8s+2CY
+92+aAJgq/HTUj9MrShxcORgP6cnGpAPpqJToPUOxEc1r0qWxwqen/IGJiWl2Ii1
4TAq7mhNBQCJ65c2WF25Bl5U7npKioLvPPhhRtH9k14NbadAmXDp20Y8/6RQl2U1
wL/8JfTy8jqN7lw3Vv3LiLz3TtPOUdchZWonZ9nYigpZV2NrRhKVh1l6upHUtTfl
cz4FyCYOqLJ+UHFw6Mi1awFImXlACd9ip0bIVEXI4tQGJi59FbiPJ7sRHehffmtd
rKarYsYL01eUOPyeuZWgyEXbPg+jhwZQ2ano/L6WRyeafYF0XIVbxH7rnqdgZIMs
hAjE8+Auu0gjCiiNV7LahhCMqEIxx1XlhQraETxJG0ynp06sB5zJYl36IglLfeN1
1+QWZXNU7X2hB4XV0RbshhBtkbBpOHxL8MYMCn8Fpx3gW2v3aF/COSys6ZGd7Gdx
ZBqRrnNC7a4uNhHmbjioB/letZAFXfH9euYGRDkok7EHMwIIxpWq3qZIkiblccvO
JJpce/UH/POsx9kVNc7rJbNnC+3RRssMADB3DykcmnXHOUUqxrrTYk9EWQUmJtO1
BlVVfQReoeqVzgckKmsSHDttIaQMhowILyGc8gmabucOY8yprfa6QWbLWy9zfsh7
cvlfGYcHLtX7Itx/ppXtcB1pb7/mkctjo8lCPUv9CoVBICQ+RBsj794VCwVAaprn
kd/qRJ+ABwSWP+CJS/L3LLFdB+dI41TB/c6GN5Ypv36PSt3LYckHAWIhZB3nWaUz
iDgp1sn7cG4Z4jfxG612VfMgtwd1qsqLKK9n8XCAI2I+0+v9RAaKtNPF5F/bqIv2
M1QnV71OHsxyxiAEfWUgisqvpapK346cSuSj3DyNdpAYEIlbdgzFsNaAAuXMN33u
j7tTXlxNETbrZ0G6+Pse+nIC39mDCqm+nXAbiaJ6xicp1mMr5GCPg6t0A1QCu8HH
2JcQe+W8I+V+B8iaMiV8rIrPBFGasQqOJTGDUfbFIf4F0X4efAWLmShFBuyTthGh
LnxiHlChjNulE8B6j579YNpLQnn17xNwUDmVNJYWxpJsj/c44Pskg7QRyGXF9xAz
dkQObC7y6aPdm6iqxaym8fTrnczfC7KP+8f86Sw3CMOgK/UyQSVQQOVBv2ixvzhe
tz6a1A1haFHPKCUuN6H7RL5WS1RJwjwTbaClWWufsiraMuPiKPY6ntNnv2gyiuLV
IeGaJTc8w4r6KeB4n5JOgtAanNhUt+4otdQCPdctVZxDDbVZGvFf2AFaJ38nqVKP
bmFqNkbmT00u2PkJEUgQM8L/gXnz94AtN9+MztiMZmOvwjV/0E2wMfs8JqFxq8Bq
pYLEgjTT3oCF91Zox8gnDxBzB+WPr5k+i6skTfrzcr3N1L6dejAWSkby+xSJbSqi
zuR/OYmop+77yQ1HJ6keuImQ88D82oms3W3/TZwSIFwS72DusRi/6o/ndIiYh7TK
s7Pc5SixR0W3vlPku8WOlEVsjp3CCDHzUqeXO7f4FpP9OVGWBAMW9SuAGUea09Zw
PRgEXHcaWAgjLfR3OPVDg+HtF6O2IT2Xe35qwZo4x6Nz770DHSboaORkiOSpoSAG
+iVpb8daDp19nL6U+ickCoB/miP/SvUCzOkDvTZr2CjtMVG7UJwitllGJu0wdAxt
Z3UcWDtHjNqkSWggvTDCKN4O94num4LewkXVSfa6BdGl6R4xI5TMp51CW0i10nwg
mE7Su+DlUfA8q33bJcQu5+U+uFkH5D/eKGOG72RNtGQ4DMt/q/27ebA4p861jDi2
K+sjcjV7WdNoSpqwghbmPA6Gz0/CqSB5bf0Fu0+KtnArNT9JwdUSmTpuf9FdvB1x
L3wKBHCcF8/7GANlvPZRl7BoTl0YhacGvKqT25NGG3ASZqEl2YxpS8QZ8om5nk/M
mzmDyXKsOvh+roBBiGqkmtMQ+lX/6ZTxdBwA2oHgB0kURBAsWnjiEYmUf0Vm8Jud
S+sSOTv9xy+JyXnjcotBy+XkDKCVD8xsBwP4AzYX8Kw1uPbrUSymUAPPGaBbv6mf
wHM9O6K929h4lqtNJyHMad6KpwFcuNGwaR6svqbJN+EO2rhX+86wt//Zv+bGTVSw
yKEzbBoNohG2yuaeLYXBl/PbwaFhH2WqqhaRI9Pf/qeQJ1273CJ8CHeRmueaV2t0
2mmuAiPSexETn8JeIQsYg5N20ATaN1sZOQnY8O8wjKycWygBQkOOrt6v1cVSupEX
9wwtcSpMtBkfyJzPk0qqkden1YSEPZmFaNYjaVBDYSHZEqQwG8VWdfnKBM1ma06y
VkZZoqF4IGBD/PaiNzo/GDmFwJAiZb33ty7N2ZrNo0uQ0B1hKFlf6PIIyp2AIFAl
zSM5LxaczAXaYtWhMDFrEAnXdKefkF38kWGlp+xD+8RATSbeF/iusVK8ruRtq9oj
Y3GFSRm81863tKlRgQXdRnqA6ZOqFI387jx4Wpq6YoMfyVRsOhznjuZjJzmlsvW6
rjSe10OF0+g5NH7lsPkNRcc2eWdnh6JhYlxDR0jR3q7uhmBLZrg4saoqe8BCq128
Drt5ay28O9haH5gDAZXoNsz/U26tLUrPFul9nO+5taZGltg0vWsiJUJmUsGTTFFR
Lijey1YzYCTxg+dl8MosIRmqLUPzGxrUY0PNLklpz4jVWgE5OiCGjsBQW3oPlLj1
6fg9W0TuYDls5I+hqmNsa/96lUHMeA6VJIUEFiMhByfWzeuxBDCxEe9gLiLSIHRn
6es3X2R/YJhZmJDl4/owyvatbquZK+TDEKH6WYuz8F+b8Thxb4LLBf4tfcuAJu8b
W2IAgQmF53Po1L4nQiYRc4bol7W/vmH91iIQgOJQSSUNpJAaM4w56zUqnxgmhK5S
SxS6nbO8iV8aLMZ+ne7N/SMlrNnuO4GKFRGHtcYYlpgQJcE5gplR3cUdxnc5hpfF
D8SL3wQE468rxv5cf+pADGOoU+hzDwk+PmGL53HGyBknUVNYXj+sO28sCkh5zygj
i4JETfnj+6/4aQhMJzMHsF1fnI/NoXB/O0sxVRzWL5FVjGtTMAiHC3kIP4FK2bRC
us6s7/7bu7PwKdgyX0LcMFqwIvygxCyD/b6CemNvMuQ8pWBj4zg0X+I1ywtmymQ7
2bd0vIMvggEfeE/2bLEb35tdtqORIdFxtX/dEgJQ4fC5r1Z9fBzkv3rxxX+0u9Ri
9FEs7knE0RAMfYL6Rlnn9pGNp6gMssYwKFdS1iykCdHgR2xYg/xbh1c33iGryA2I
M8LA7REq5Qll9Vnexj+aaUV7lsCWYrtaTtFK9Le429YwpZ+/xFfKAyxHOWkQbMo7
ZFjGaPmhKAk0BuIZ/pucrvELOJywdxCq/4auojjhzpm2Gkywdd+0i5y0Y304ehAX
pOzN882bUrXD10LjIrydpEgquYPU0oymJupG/Wn+UpegTnzb2MqX0cKScHYhQIA1
txizvv0TGADifpY0qHmiZbItkNLv3MWaLEjpOWOeyI83FAgPNosNG9Q3pL76QLPT
pqGqrfxBYS+DLRz33XyYLwHaPbMUaewZDUajF/vpfp9f4jfbw9skO0kJVHLBvZ7L
KlO2HY4p2kBRns6ffXCtl2N9MgmTSpjbmgAIlap4kppQ5m6eYddUjNeJ9poPEymm
0xWbSJM6aFASZLELwyFU4cGWhRQFtVHK1NuQ183ZqJevtyjHUOnWuYas76eLflG4
adtxX/wZX4NTlPW341TwQDIBGZLEKLMpTLDhaHfllBMI541ALPwoMp3Vb7YDB45q
GaqoKal9nBcNQSQ54A8U5cHYw4xU56j8zC+XlHSFXXranK44xP/ywjivYlTeT3br
O89k9CKNvmcD3cNnXTob7Chp2OOyt/XWhHkqO9O9lBoBweVdH4RGhw6C7VuWxaVE
2lVkkLidLRtzr0eQtNugKQJqOwvKNU7IJlwsbVIhUJncBzE8YFjmjUqucHEoF27Q
5jy0n92GY/fuvIB9QxqeV5cukOlUixaA6LqD+UjLKWkYVqNXLOqyuPS8vgAh46sD
GEzmjNDDD2i8eFxXLzgK7rbMFb+w/GdCc69tvgI5EUII+vVgCUug3Q+ur17dndZd
GsoXnRqc555fwXCf9zWM3B4hy2/NMZSzBeZkdjc/RX1yHynJ2e4G0WrXAjheXNcI
+HYZ1BhBaMMi0vWNGZ+rlYWzVQ1w6T8CExTwULiOLwpLpel8eXirWp7YGV6yMESv
4ayJuJKn6MUj2D45Mu40kI0Le9rrPkpdnOi8zUmgsjFW4OLEftLy12dlCbSaab5N
iXH+rI5mQ6rl3l01Ceh/cs6Sx6R0VdIg1LZYv2wRZ/FETqt0Rbu8bDxf5FYhtHI1
0lLmbeYUQ7A5cY9zv+AuCHyQJZlmfYNjtHNKyf0tUPt0I1tIC2p6Lq12EKL0L2Hr
C7CKxVA5+Ntw0AcGdu8k+dTA8qU6yLEXMs+Yfw5A31mrCObNtiK/9GcPADq9+BlE
3xaKkm/25BH9dovzzLfk+AHR/reEHlL4a+YnW5anu3NvVlSx59a+XWb3vZomsG+U
S6ghbavVhSdSjkRbB8eZMjJ6VwpVO6RGYloMbBkpqqPod93w6ZJJbIOkjNmwcKmR
rDHExq24A2wZKmvzJ9ovFY4uSWXHEdrE8GkJHhops/z4A1xcPPa79TlpMGgIiFfy
FM2X2KuRi6n4T6pcF0w/ZT+dHnppV+BR21eISHe8qWXSg9TDw2ziyVzC/EAc6y+x
IP7m6IF9agdFAYh5wa8zjr8UASR01Cvb+tOUzz9kgdrTENgvQIzQA91TX3RiVFaK
ffKl+rCDVMmHufKp9icGRK+0ckArBRH3giIh1kxjq8+JwTEw4CM0vNdWkEl7hN19
bXWbJt5IACJB+Y6Ebi4yeIlSIj/5JsvqWzKyf+oRwMbXLTWNJd5C5epTiOVo7VZU
epb5IJm6Dc3C2KgFRNs8DBT8b0X46wuqSA1y2sPspJOnz6oiLGEVx0wbeCC9/DTG
wiD/kB12oJymwLJ+jgVWUEyF5xTAbai67OfBk9RjXn8REUqsmrya3FoRD/2tQWnG
14CpRzC9wOW3BDK/3BC9I+4bkoel2CrsMZNpHo/jf6DHV4GxeiYplM6oL+O7kjTR
wSuZabRo8Iwuu3eDXGIIBghyfRR+DbPtN5OQjOa5VAOUzUlVfmrz84zqd01hBHMy
GnLtsZZbjSzbjjlzUe4oIY08I79f76odLpSS7ad1QDCaATNgDE813/WTuWYBuI92
zoc2rwONRFa4ih7Sg7SO5HX3WX/bB/61SVKm7hTCyWTru0ZBMpzyy6qumwUHnauZ
3cGtG5/h8xZ0Grfokz79tXUOn9zl0YwC8YEASWpfzaa7wryZ/QF5km5lkdBYeJE0
p+u/iz0ChjKL8KSKWlsvOKUcSFZT8t+PD+Fu34glW1ys1Z2mZIKHD7fxz4wNZU5l
SeGCJAOJN8jPD7G8hJqg/i1FDv4RekiXAKkr1jKvLcL0g4oU5muPZG/J1MC+5t2y
gsGRVM2BVayXIhYbzzRAMsDKEcySGPtECB4SEf/VYZ+NesoQU0yvmZ0QneNe+ElQ
MIIZ/SpLi8c68etdPkIPNGrSKZVCAO73EFkDrA3e9TIL/znsn8VOCBVQ9ZutO9X6
uxnmKNPVqRuzR1EMffUC3o5QSPeP5kdWMjuvH3xpur0NeRNV9VDVnACWBOr1ETGc
Ys1jes7qLG9WMKUWnF+qu+o9snUtjJAa4Lnqy7qbPCf9iwz0kf50wK+yqJLYXG3t
7/F8fOpEwuFytnOHgLUp9HL1V5KRDuLS3Cbht8S7TaFQGA0R7blkzaxQFLzwtz/G
IXKtca1fjeHaE7saSWNgZme+J29QNbUz0yvuDWZK06fMLY0VCZmc8278uTq0BsdU
YykMd/3+FllZrYcC4KzYlz34gpJbZ3j5RRMscEQLf74FfY2Igi9BOMlgRbeIWgLs
d3lV4WJavgii9pThVph80EXCoKeC01Cpup1bqEZxbRiUee6JILZZuiLvFkOb4tXi
UBJGw+FG62KpQzxYxlkeH9foxohInr9wqcSGAB/SfASr88MvKwwHsLcPLB8XzSlM
FJz7OTl5StzFagg2wTdWZ7zSnPgVaVoU0UC1d9Lxn8UX11jqIJ/DwjDZcUVw2DLi
2kJRrjyTiBR4Xl3lGKG7veBy8+ZfjSVjWY1SdC6HCtqvhM50RoLiWi51c7Fbma90
fFIUWCOizbYFdIg+pWgN8yemLgNyU6TbPArV+At7SmGw+w3Ns7uICJGKT2Pj77Ep
fRK9kQChMk6iF9VUXvhvp5dbg6Pe7FFGRoXSdO94yDBAZmA+/6urvlFt91SXgtun
xI4i6sSQBYaUP7LJF22+Qfh6X/vsGUk8PjxkMn0YP674vUtPogiwvXgrLKQ/j8hx
A4336N7IM7A7sjEY47tTEo84D58f7kYw1r43vBtfHqqm1JRtG2sZocTEmGv+Newd
IZg5xrYKRy6vY++wc1ULrhumJ4E79j6vqqM8Pv47jXv5MwoJ/6doTbS7JW1c+2KZ
FvPYJ10U6OQKLjlGGj/qehnwIUx3kqYwVtUqsxIWst35i2fhSOsRCDSPOAMWv3se
hSVQumCdyr896eOHlkPzP0rzlp7whqhJ4hyN2obWkImzieGTuQyNLO1AR8EQ3aK4
olkJ5bA7QVbaMMp1UgCXqK2a3OYbm9p1FZiUT/+HJdo1mqMa/HLyAniGL5K9rIkU
4Kc9PDlDry87z2iX1WvIC8aWHopkte3JSkIT6d489PEm/Ch5+TE4WGTUjv+W+Kag
FlR6hXlrTXmHBagiNH7nf8Fh/Xac5J0HS3n3Kw+QzP7OrgE065Pp7YLchh53+k/G
mF97TvUiKTX8msdWFibSDrc+ybbgjWrUK0Rss0iHFZr6wJr3yL3FplE77p4k0kjh
Eti6nmcdcc/VQxun40n1eKqwJ7uT/fUTqVUEO74UWsrMw8T1zMSkZaDH+5hop4rQ
1rznRL5RxBXjJyo3EJ0XYGnazyjSdy34qrXhSNL+tCPRrmueixT2XlBZ4mmpkwgx
P4E9DlZj6pBDT6fpFQ09MPI/26gZ4udvZJGda8FknnJ9rrsg/dcV4FDn5nKz5uzB
Kk7dSIyMcPEc2CW97muQ3IFE2TRd5g7ndvIX73s6WgwI1jgMmSgN415IFAWTo75b
Sr96mb5TlZWh8XiC4/eGdvhIED0ynIUExEIFPAUr3TSF22TSmoTIkaJdZK7B737A
/wwwYKgYBuWi6pr2KykwVS0k9upf/Vhbh8KDPAYgM6o7eZVTzwJRNJv0xPhoiKhU
9+ZC3L/2eLoz/I2m+pJOS/k5AVbPGEYgvn0OPfSCcB3918oXMs7Nfyk8C0BMPyc2
XvbhD5ymkCvi3EuJr6sEp3b81z5prLzApZAaBVdZKWe6YuTZ93S66PALZneIMoqo
mrMCzNWyHhfIEOWUGA9wBuA2p5X2bXrqmeG7jkr50gLAXoJMKyivn6aPFBePUBgH
7CcZ+P+PzRQ99n1cmNWEEqSp3G6Oh3dz8z0UD8FHYEBNWUj+Jw9H6naUARLJkwDy
GEPK+yDn2JH2WbZOh0c5EKe4R/4zlm43T9+Iub5j5Z7fPFhP8ujAyEWY8DPj/w44
StjuUYolrXA3w3+5gqXwZOxbbQVtw+oyE1d/xN0idQzBuLgsBTYiWhTk8Usdxk3+
HyHT0tkbsDn7E3FKExJTcoeYb5dwx0rEp+CTRUnP6xxVO7UNLmVMaztlvwTi/rVN
f5cRzpoBhC/apZsE+Leqszkw1rORzxRpiedQsKX/QnVvv2MP36JfUc5lYQRrXLg/
hTWHWpYRQukq4OUp3PW2MBPIRtchEDB5zJsUaB3h143xGzuloW8dRfgt7SKpx/Xl
6k/6K0uNuOciUdn5Ohy3k4Mqi0tFu2sYPtD+ABicLy0UEQScFVfTmiB2gvUcYqlZ
MUUef+CvnW+h0LPooWvVYqMXe2faX3MCRMXfOHQSqm/KmN0LyWZTvHVQbTbKfs8o
Obb7fMikx3oiPdo/rXb76rxqmv/5kwsRicGOHD6Li2UJfZtrpmp0+NdXhl9W+Pw5
buV88loQEOHmT2HX75J5RyvTlC/jwfEh/b057Jq8Hv/esU+PKq0YE5ZTueS+gIZd
EH2FqBJTIRhuBD3wX/bfX2G68nLYIf+g0bo8OqdO7Gx1m7MCCG7jYFqJY+lw8Z0o
+nvpfZ79cWB+elHzoorunyA/AvOljdleH+LbrySdFE5sm2erXPTmDLLNkK0kpmXv
N2idq7bsNDv4fTWb2jJ6iDGzHWGQm5ISOjDsIEhfgqg7ggJvoBuNSuVuE+Jlx4dv
S1EqPL92KOtowpbBMRVGUnOFd5KTl1qF7bC+48hyPJeiZ7PdAizrDx0F47CCK6IG
5Pv6ViVDD1ADnOP9Dprtqk1C1Gay+XjBDtArQDj1c2wdrDY8i32Dwx0Kvweb3uwp
Ikkh/7FeFUqQ82WLW8G7jkBAvorBdm5xRGuxLfgtOW+7/YwRWanZQaqYFnhSdGu2
A3qVOguOseB8zlyWcsXp/Aegsn1nGvmpTfru6aEC0qrxFycsi7wsZ7nTvk/GQy18
qRpMBepMFNvjNt65TKPb8SdBgphet32RUyLA3Yqd9zRAzSGkrinrucHmdjE9JgVB
mpLF/tNErwtxYwi0jCnLZINB1eJxNDg+TzAYAzjFHqHe4kQAgJAfTAxzxxdxRP6y
d7ev2WmKDY4KYHljSASKbAkW6diIpB21IWYOjecUnAU6/Z5zg2Ft6bBZ3XPggEjH
6Cy4GEWezR480Q24x+kvL6Tuvf+a7aLVtKQSLPj/l8j5VyB5YfObKzVWnMEUqC3q
BqipgL/wWd6GurhWGvesgnESrsGvd3gYzquIHbpqY5p1fyBid8md8FEqr0X8A6O9
V21LXhPBY3e81Dea97fArQfo9tYLVsqP/r9pcy7c361MI2yrQyuV/Cpvj8ZzWcHd
uk2kkjgVjP4ggAoWTxZfhtttK+sDA/McmzS7fzDE60GAmhc46oDbxnKBDu3deg0K
//ykvqv/AYYGFzzwKSGS64XAYEoZ8g3N4BHEIJZgzsPy3X5SVgAlUlV0Wn90Ss1v
Dt7pWw8MECdKAmN5WgVfms81obMxNvaplN/HTAthIMWBMaDwPiq24ppWispfQMxz
itOSCSm6Xe9tFSRdQIUmK01v2N43sER4YpqvExlRmOQ0bixkCqEUYYgVB4uLypU1
iWi/sBh36vJJt8YCP5ZtXxs6Zvczl6hnmiSa0caDEu1mUXHhJ4zI3SsqL7u5J/q7
0KbQU/SecgQ6249EEmKhBdt840C8S4utV7CZebXN6YGBfLDzgRKj71n9lf5qj/eG
HO3rFU4W4qyWoMzUm2cAmkNHomX1xzV6PEZR6jvYo6GNbjKn7ec6GzQIdfL82QcL
fMRvNchPvmXXE6JaJnJaepNLECnHh1AEgx+p42fgTK/tQpPrdMqO8fZX4QN+/zGM
fSaPwKWESgiJggmaTn/yhM2WzjRki4kgAxiEC/E3a9ZD03Gga8Q5p1yJlvv5eNJK
UKcnjbu0TanLpSrnHqzi12o0J4nyYcxjmHbRC/P89/vDGTD/OvDh61gC0QRH6L2A
xwOgwvBDpxEFC8vD3EtngfBxuKQisq5ue+/dVLzAbujIgB8Y/n/ucnhDuJOIQBHg
TRUCVqQ9BsMZWL/WE+z/jPo9X2dzmCBJ+f5CEeD5RvlwgsA2PZnzrCCVayJskMWF
T1P3fEAVsEUiX7t0Hi6/TbY5UmJvauw8Ur4rzAJr/ubGw2Vel9QbM3I2kVdO00hY
0rTfTp62E66Y7GPntTbh5M3ctSTGYh8zCeQ3q4nKoKMWetx9YHWNnStSwewEt96K
qNBVnGYHbnXmDaz0YSuu5PH9KagbxaZXt8KRGoH0bhyp4p7hr7Vo2WgXLq44KHzZ
GtBIVaXQIf2u0O3Cm9BHLJbUJrbBh3PC4NkflpMMGsTxgyKbwqANpasmLdWiZJW5
YIk+4q1LNhlu7Tr58jJF3u1O4xRx93N1UQvsdFmv5hcqcL6Z2AvGv+ABjUTm6mUv
QiJTTfG7zsRQ4+uDvBa8/htzm1jrWPR+I15tL5iY9nERyLrdgPhALrhDKbGybLnw
JpdWizePiuaqnktPzRkvbwsJt/8g8kR0nFwB5P3D1AHMNaRYgtO7AAw4OGQEyHNd
eBo90zpk1iZsxmQLgaQ92FAkYRICvVUK5zji6fy3fHR8bRPFMKwjFU1xXl8KYtw9
usfppxh/s0lEt5s4Fau/0RnGp/HagLJ3kbNT57Efl0Nml6Y9puQ5QzrwD/vJY3Dc
Hy1kH966Ztxwv5pPorIrR1OpU1HF1zPpKFqzS/pNU2DXoB/LH+m8nmeQ1CPYTTdg
6OEPReDJEJXqXV3/DK+M0/vw+TrK+HreTYN0bVYGKCj2a8Fa9mYV5yRvybtWZsVT
C2L9tO8taikPthaPauebpKjy186EMeMqaXrhZ2M7LG0bgM6USLbejIPMIrDD4nVl
TEG938Y2O0nzH1ClIMfUPSaBbGyRTTWiqJsxps/7LmgQWuULnwCHj/yRZ1o9CVfG
v4GUmpqCOxeo3iKMXLKLRP+WseWpEOrS5M3JyPmBXgtSd3Wc8p5ay92LLNnbTKi+
96b22TUM1LJvwcfgtjcIor2Rk1GCppdwzxXjuVrk5O5J22NBM/uAUBVxTHIT9i0f
BRRunFGekNj3i940xgMxmaWVlC9LYVZuuoVK/ZP+swjVQLaB6R4u7V67QLzYRV6w
YCj6FNubMY/6yErVw/mOew7ZOxPOSkoqkOoHWSCBco/vPJHqQNd+uGVQiSt1TEDz
kJZNZVCVMnwp1svvax5HAbGspgSuuovrccELncQ6RtbU6rhLNoGhyOr3jo7bd+7C
3RrYaJ9ldVqEnQ+eXLQFYAflmhRq8JhspB1d47HiUu3ckBJywcXDh0KIxZ/vFnUr
qkR61unKad2xpNGfnrQ7CbKuadIGpozWlRnfygK+btDe90oI7tDayD1c5qkIkf8u
DHK1xtKdR3joTWKu2tJBTa21UQeH8AKjhOX5rEGUcsFYPo+nvgPErIeAFWmsSMkd
zPYlhY8mCftqCU6OZb60fui2fHx0m1cbEQ24NDRmN0XzUIhjNBWiun+PmMWN0XXI
/1O+aOm69tVDir3IGQiY8sfZRIJsDANxyyCwXl01CKilIZYW0up5IUFwDlvuKDro
PTS1N24Z9BlfgO19v95IwFNepOqEq/WiAQ87ndHYqXg=
`pragma protect end_protected
