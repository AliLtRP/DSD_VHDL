// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oW3g8FLPA6eHtCmx20ZoRwaK8s3JeWKYL0RDZDhszskYkaGnI5bJU9LWFw7Hkyr9
8I/JD1Ixfa/Ve+BzQINRkv+ZIjCxxx8LdBm3uvsdyzYqtdjaxqrkAC6TGjnV/ukp
4UcI0qhy1SiBgqa8Ll2jpiMZay3JtfSVRrKA3k3Eps8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48304)
BtPWtBV//7EZJB5QGlD2t97tus9I92J5wTbbdXlRNIadaLRzq2pfMmuBDN+/vIkz
RcmsG/qVcveCGtrRlvEPGH3vyTWD/qfP988dRWX8u3DYvbnXgbLcOkzTK6URiHcK
qwYHC8F6NGMmf8aNrhWReNA9TAb90BO8fEojHcEOahj4ygt2bHP8hbVuvvV9xRU8
hB+8xY8o7LSN2Z/SmEzJGpZXfYZJ7gJmb7y5JH+wt+eQMFq9yf86BZnRqEMGAyMP
tmy4d+cwBi2mJAQMnLRRr0ZlUVS4LRq96MhUpMHAxO/q5+wS/v/BIeTOYLzhLvgh
dteuA05RC5x6YLcSjHH96yQ63emKdFxer7QFT+mp7GyGIhXXtFnMIWtPHScxBiYU
NLRQc6HEQ1wfRvCsIujDnHXsMP3vISlRJh+1J3O4RKuyTM1C6nA6+u39pNt6AYpT
LNgLB91/J9s7TEKawSrDZECHED8DRDKURJ4p5+zB4dBuLG+bpWcCOqk0TTdDRxJh
u0Jf/sNiYf1ltTCevaMh/jFoyJmYfZpnZVlhECNOw8ltrUbFzdIu0xj8+l5W871/
HPHNA/aD24sSYWV9td1LhJiGaNUrTlWKLjnZ6YOIVFXPjT5WQJqMelufe1nfyOfY
V91XA1mdN0tjDq65x/lT40NsC/wme47Xez+KbPdaxvqm3oHZoB9lW5/ZKL8XD7oE
Z4GCm0zySwiNaYNJYiJZX/kQsQZQ9/FK1kHXDRixzf/SeZIfJ3uCiau+4iV0VGHL
kzTT+cC5nHckRF+0EcIzQ7Rao6JE+YqExkg6M0rO7BIqUInKO/L8DUcx+UQtBzK3
rG0Dun5yQOBHIAYuGwYh9tPvj7HUUOGZciLh+8zptxeVLVZQKKcCMs6EWuWoPyvy
YnsbjHdmF0UJ0m/JSm1U282bTfD6qjWGIt5L5xPkMZbLhJOxvX2Z03+3hy4kI+fc
nEngCOL9IdeW34RTEcUSmKaFSfGLcQttg6Wk2x5iq0vi1374MmU+QuW2hSfR9gPo
POei1P0bBMz/MO0eZCxz5Wfc959w4g94tYQZEuCRaXuH8Ov77lzZUMCfQn0932Cn
e9/YRvIslDcMblpqKXY/N7qAILiowtPsjG+VFXumYR5jueHlivW3EREYbJGzJ2De
nP1y4TWnvSO0mJD5m82IqACrt/dzic3b284XPZkXyG+45pC5rPuXT+L/5Cqy7cPN
XzpcQhurBZDzKcj+pyw26qtHPjgB9vEcF7NA+hevQoCvCcS6yqK2yZZsUxLnidXP
35PJ5rRruf6jqxk1/X7pEHcxe9dBSlqXPMSMvSVGgQpdkT467YAvMErjTqpMbxrT
oGRjUrCocHCK8Xr5FtGvx3cGgtZKDgEovtYstKrTWy67YHEET+9LrRgDYyCx2SIm
AA5ni0lHPJ7/zNaB7ftS/SPcBAPXJ05Fxu0Y5HvjrqQpZmzpC8pEoyxWQc5T3kyp
+Rs3m2LXVwOGp59vabM3Xcphy+cirJqRhPSmC+xMEv3XfXSs6bDREzhdWUNTbHNY
w0E1d1PEt4XUFgvZFmVediCkGZ0Mis7l0gyygvGvJMoyRzEnL7SdhQkFRCof6hx0
wsj4eHooYiYyGTLdrhPP0eZse/gYCnL6vtOvqeOdTHmpJ1vO818HGQlPsanMSeNZ
dUq+IvfMaPIQhA7Ble3kV3gJXCkL6m5x6FMgFyyAXw8D3JH3Bc48VkB0uMTGFK8n
oJOKdIUdq/D7bgckyyl7kiAmvAG44EiOkQzpS8QW6cVMjblH801UWIu1CCBl70+9
qFJ1nbuJPUHrfi33rzVBxMjm6pOKw35gv2hsaUNrtmgySyBvLKokUOWf9gHgUyCe
rhNQ/7ThrYNj7aMo1qGrun6ZDvQ2ZMivFfJeoarmowlaraaTL30liH/03aVLDIY4
3FRDc+aXkwZiSbwmqV6atBi90TL/9V35SC1CSiI/l3zfLiqwaGRq3T54IAtHZHWQ
iYfOBNsLSiL2U2XdqGo/UfoDgtOvHuZ1tarXb7IriMggmRBatMwpcAU6eL/tQbBn
iZ6lWvjzAjEQiOW9WbMtG2B5c/4RFB2037n4UcTic6dSk4SJM+pH9fNeTQaKdXo/
SQuU3pnNuTUeF3cS7FiqQTeeNuoFGdyjsaxh6D3Uafa/ghGfV07Lkx5xdXhmM4wx
24Eg8hc5rixibLpCzkHJ40FfcN+xbKqlkls83qcfkQqu1kst1k1F0DZ7x9zPF4R+
CPVAWnkY+ADn3sYTf2u5VvrQj1xrvnIYhwD+l8srMXFhavOgJbDfAQlVcDGeCWb5
Gg0K1ziN0SP1b0Rw/1jwyTqYuCh0YV2ZrahGGHEzFWE+eRn3gXIkYYCsUwvDkmjW
l7OhQD9eWKFZklau52O7owT9lhSLdGtWMlAhKik5nBkdAp74+crMGDrNYylMuqTk
9h0GEYJ1dQfNnFy18yASqG68Iip8nUpZGyZYNhj2FLJEPcBeKrXQ5uvmKexJsHXd
rtXLFZoi4X9wfgnCFUag+q5sv2677WzE/Y8rPaziNqTVWjnsCrVsBIiU+7OVqRU7
SjnMW3gm82rQqoH7/QY9cdY7K3w71cXK/6aPwYtxwvF9N33Ul5B/zVwtimF8oLhF
f9k6aLsbvRm59jtBl+T+oPT8tDiqDkH4Y/wTAE/y7NT7xAqvFfQ/KEI8QtH4LBwy
TLfrr0qbRP1cId4nYM4iBcXUQcUYwjfn9Xs6J/Vy/zlsXV3nYj9TxzKFxwt9e8xX
Hpz0VKW+To89Vikw1xgF21hTijuX6YfLDiyVOjO2CnJtxRkgVtDSdD26mVuSlEHM
lLDRFHBAH9b+DIyiC7E4PKgG+FunrmKyPxZrp2fD2XlZs8IdD1Lu4QXoYDXgihqK
1BgrAIMwo/WLmUyyEtMOy+HLk7u39EpBDmhttJiFvJBIB6Bi6dPGcy+sfnM80EsP
bgkUE+CaRaX+KUBnDR7Fa6L8BRlmga82QbVdHTYgY0GktJO6ylHUJSHeVSKwrmGa
8Vd4kbnHN9hghIVM4Y+oWAftYXbxHuDhFL+YQX9w6GU+IThkjC/Bb/NDuoU2LO7M
n1dtmt95QHHcqwH///23XBVXKIMuEYISKHTklPSIHm37yzQ+B4RDVUWC/UL6VmR6
ASBLm8gWTOsnrhgOIKELydoF5yqzmbDNQPUoLnCM9dQ+hSZOJEEY9LCUKIjlI24l
cP2VrlMWSoT2LITsuG3fYKRt6ksgRtsX4qJ99VT+el1k8hHpLw+SeTXxeal4lk14
PcF7S9VALDMNzjf//PcrwsnCQoJDAnMhatjNqNhRtKQbQxMVNQK4CRTtgCI2wgta
cRp4vDSxCJCU+D/oSaygwpZeFLVVi+SedQ5OYy/vjC/379sBvCenzsmPDQNaktkt
rrUw8k3a/Ir3LdaB7+NWw9gpo0mCWcs6Kq2K17i4Y5AAwicGZOW+rV3Wux+Grp9e
5iOIALUmlg0pEIuN92Etb9FM4QCFFBNTiDIOWJjPyrJJ44j7Mm9E/LfqptiLC910
1ffwn4hy/bBV+RnSkVyhdPVsMHIZk/FK1SD9CeXKYSjQszYrGzY3wmeDCc9TP7X/
Af/h7Xg2IROFG4zmppjkflNS967VwafoLP6PjNCOH9P65MWEQ70INPEAuisxlhBe
P6aNo++pt7n9S1bxgpW04B3wRI/E2Xmew82CkwWCi1grI0AS9WKz7sBv8yiff2Gw
JCxV3IWz1xDmGe6iQu59KKGupKJL/nf6FVYUwlIyA+YcrGMqM4Gf9T1//lo1x6Ql
G+ZQVNCBi6T2dqXVPObeXZpbE31xNA8PodHupM4u5n+B5us/HKBNdctj/nUk/hsH
EWnHDDV6p0w5MpbssJuD8ApyKfHDMpB0bGOLAemj9w3/E5Y/BLg62lzz1nc0xziG
I1NQDUa6wVCWXiuhVJoxLHkDXF/N9Uy7s5+pCw78VksimG7eMfbDRPoOTG2/YdxB
deTNAoooDgDsh7X/dDYGEArHUZei/9C66xGmH7Vo1eNpBiwT2u7QOyZp4ciEeUrh
CixuXYf84nZ3GN5OfWRbGpPB8QBClSNyWcuHy3B4OkyfLyzrIEVDLoeCdHjdMfkD
LMCMOEH9f/w73TuaWnWK5Q2dpAYj3FV7KaVu5SOlMzHXLNpbBcXRf6NbbuVAWcnI
BtEQ4K4h6QNU+WqKsVncSmL425xxQCCFrnQBebpDf+QsKt2t27qFeGty3bkhoxnL
N7Fnnn8MXv2HVA0cZFYZZ3zV2n3NU12+ZiGVNUN62GJjY5nQZsFOfuBTHi127yPK
zxmq6W2AthIy3sbJNr6KWDfz6m1yOu7KD3n0guyKZnF5Mg6Z2TD1/jLoE1Dz5cKN
x6uveoutY2BIzfLEdY/Dl5aVvbkwor2HBOuJWvcSsgEXRLYKN/WnhbWbUw4Prh/F
rYJt9jt6ksX8rGSUdcAq9LfLHNgan/QMnqGYHg4BixuUR5yKpmeSTBO08Wv24sB9
L6D+WfFVNehjRuE2cf2p0+Qp5aFQjicW6nZbYMj+H8Oql2mGYvJH0C/738q5pMzJ
5D4kX67wwK6tCE8wZNrDWlLd05ZIXdB1f2aityiAnVqtMr82IvJHbIQDB5zUlHeD
hDnrkHgOdg8NYDeIHK+M0URZO+mBtjn2EaY5xz25p/Yuq3KXSzS51exGTyU33/yG
2CXB4zT95e8YSS28r9BhyEpwKIIVagFHXPG0fjoAxiRuoNej8WquRZ9dqMJP8WxX
1eY0j7mXnMUPnCTtDw+qHOSAdDodspCYn/K62Yy6E16AYjw+n5gvg7SBSfVylDkh
o5TsOwsdp4PgyJdi1lyqWt4Y5XeEA36Wi/+NxnhsFJR3Da5tuxRBTMHDOTOZJwU3
hGLkU0W3PFzaFFjIj8Ba5wDOTjXcCJCUJ4+Yb9D7WGKhoLGy9jmfG9W5AIFW4lmL
nvZiB/R7Vc6cJgIrcWf4RjLl59xNayVS/MRQjlO3O0eAvFEInMQIeLAh9twGE25e
D79JS0jPtBE1Qvl82r1lVyO1d8DPjDd5TCSMAXtNcVbyyPrRHiWNX1iz9ox7aq16
84REcIZ4goNGDB7WBC8bM+qEKnZhoypdQB5Rfr7mHkWHQoCBvssNbBrpEPKrIt5i
H72SVXAdHpFYg9nKXCXY+PGXje9FgHZTJUKgls7JJLLEYcN3QR9bv6ke+4lfKPOl
gyGcKLXcxibPEM8k8bh88MeqgJMjG94UL/Mv8zsQcVh+IulocrwoeY10fPSTOqtI
m7tvLYZUBWaR8sdM0s1fVuLc1XW6YqlyHwIihDmZ7I8uupWr3v71VHT08yqmLXaz
9tTIWDpZf/Vq+FUlgj0ic8UVpous8eBo6EHE8DnveNlKweBJdYmpoaAZHy14sfP8
kY167PTRAzkEDWoRjTVvxte2UDix913XWBNEBHxhk/HABs2u8Jjgu1p9SawNPZEX
zn+5OfNVhQ75lm1e/C4h8exoamhNUvWD7oFo6dXuvq050a7F4/fxFbAHz0jxCx06
xNRgdCUl47B4wnzbrUaeTvIakSOyYsKpwYZofqfybljxLcQn5h8+tlP1Qnmf46Ht
FodxsVp5Z03REgj1Opk6ZOGQ5HkgY9FHygSzNIkyS93lDVdJSUcwq0AtX75f05/3
FqXWWGSq0akujznwjcJ3oaCRMusSbUfrNufnJkaDuAuxsyWTSXK9j1k8L6fT4pI+
OY8+/6k9EP5tNwu68AIyXJS8/oXosdCE8NDBxhHHRgpEk4HzuQyNWO4Aj9hNiQHU
2kvcHPJxx3qgba+KZCB3MCKRTG8ezGO7lF6jigkCJc9tXN/KJXjMIssbGJyKWYEF
t6NGBpETd60uMyEsw8fjj1FWGXYoDk3oy0xvB7cQVVAEx9YrXBo1yeB1/1PncApI
HK42YHdegjXloy70uenTBZ7m0JcMw+WpxFQb4A3BIwMrbjZaCUb0Wna/BJbAqGhJ
IpLUvULWeQ7o00Sy0cs42gVajDTpWfD7xscbcAJPNrsHFRjZc1KkzV+eN3dgSScC
94qfWCcSHqV9tH4l3zcH+0MwBxkFq/dvqfUHL9N1vhp1AtZuboooQx5vOX/Gc0E1
6GvK+YyhNJ/GL3fJEVFFBKCU2g+XUdOoo32T4euKbhNJFkFNITm6w4PUKpOJdys+
Zwmg/mlqwyGBIW6xij1Jt15eBieuH0TB2y+R4jtI5Yukbfe6X8xlOpOdZ1g/9Qei
0r0fsl2kOPixxC0bXWzvWKKIGNfihYGCuR/AUtG8tFvJDhgdhTZZiSoxr2z8Ghy9
Jy6sFYAK80A3in1kxEudUSnWOjval+korNwtaEu5er5h6p8/PUt7e69LNrKZqFpI
S+P0YCJJuWTuf+EjAiTwJ2dhuUHxtxNi7oY8kNojr66msKCeccSXh3wZKEO6ekGp
2KBBtV1qA6204ing8k24ks0nHyMWfoT2tHNkLUONw355/RUA7KpdIslMk0tYC1Px
oxwZjSNsGC4jIXS3eeLO8yyMSpBxvCmiDp+XHiGVL04nGFix3nYqAd3oVbP9tizs
atNJ3MXKDF9Ni9PNmI9gNzsSc4P5ghL2FQ7NU1VJHhwiczRaNw+jLvRrFCEZodY6
Vc3q+6jVHuFAEOs+H/n0npij2QhVBmrydeQi2VukRbCNaZTnuopYihZ94s1q8qPQ
CsbqUghiQZLDkZeeYYdO3ctMg0gh7fgCF80ucMkf0Lze2z+bOCl9NVUK+VZ7WvfQ
mFN3rXP/2r0MXmNtGKI9S0xWmnWNAK0etHi+NvMBuXzYsAWfdNLphyAvdV8mJoQe
iAWkI73HbZ6hTG2zL4t1x606ef4Jh0lMJKfmFh35/1Hz/ks0xl1RcRlYHDIqE7Rj
KcueLYFWZCsDLMbCFJdrARpxyV6Waz0Y8kL06k7xexA271owU+YEOm1KYias/+47
aP5lQzpxW14lt6+8FsS2NVgeBuPZGM5jK+W3zYM6kLqeIToG0yiTL5K1sWlF9OLx
9rA9ddQUw16HVsQRLrHsVwE8wsSumlevQL6qVdV0YtvC1syglwMQinyYDjTfRwd9
Q9XEgHhjkNf0k5q3AZImums/efIHoe8BHJzsdmr13Exnck/eIbcch5dfRd1d6ais
kV0r3KaDYKK/9ADG7+eT5iL8NHOuXO1ej++O6Q+pBJs74ZvyCC5P7QikrDA1SBkh
54laH89eS6+wSO8NE4smE8RyqQ/1gx9Uu3AhSHJthNwgZNeTXwxmEou4rGTb4ejk
YFoQkZxEyPJK5A6lFWoWL09/9GBEw2G8N00v+PsPJUO1SlIVeq6h+Th55ATcS2V6
OcRJocD/fAAUF2M1OE05abmHkNVC4rqEICpudfa9mAGDUEOjus3URwL/B4sMp5/H
Hy9iJvHy7HlcF+55Flp0K6m5iHPUXAQJ8wFoYEeNC+QIFjIR6eI7rBwsWrxFfMcO
Rn4piAFDQpCSru2QXs20piYKgEvNGJWqai3lC+FTso/26lU0eypjCgLSnnOIpr8B
r5rkkGHNHFCKV4rdQPKd8amiCJzfs9EBDpXfVuwA7bzeXT23DOGJbereW0unOHd6
cmWx/+ZWJhD64GXV3QZy09c30MUBGUIoB3NonWIlp6UTi6nsO6AxoFF314kdTp7G
n4JTiZipBGsHuD0WHwZf6ZYRDbvwlqqtfZjWleyVNsq2lSs24Mb0fYeEIwwpnIyI
FPS726yxLFu5QfxWIGxVdlw1+8yItedKRjfQYLp05B+bZVpd8bc3ja+pbcP+cWtq
7l8xdkhXo1Uy4DQs4TfJ0zmFRqSLypK0Ot9C/EBLJsnzMWVloEiP0jWnD+wy+SDC
YUvEQfPFsRCQ5cxLVCvzL6sgK3+IX1BnDFFLOxjPt2S5j51RTzEg+GeU/phv0XSw
nDDciCbvliKl+GeSIbAprathYwzRwm8Ovu9w9p16Zkr1HT18i1t+GrayFjZ/h4Gx
l5ihPy4Be+4Rlo0aCXzQJwCtnpo+DeX0i3VQtXdv6KjnioG3hh/OFcpYTyShXk2G
nMzIgVsppn0mHWMwI6kgwh2zb/LYS59j5ykGEP8hXBIHVnCS7PeqmhlxIEZjHy2B
JTJi05Oo/5v65yhmBCO2xHPSprfssgRYNQBj2k7kKZIUOIGzhMdnuiA3DXniBqCl
ueS45KdRLFUYQcq/dgruyIsh8dSH6O+gWpEfrddPJWMGddyoKWZ/lWU7M8qFFf6U
n1dS2y4TwzVZ/sFmRM+h4BVcygyKCyzB3o9acEPdYtMXonGbLzM7D22ebVa66K3q
qduweKRRDpUwAOLUVJE4yX0ayrUIJ14u3YCQxq96deQUxn1049d3IW19Y5kBVYQn
RPfhHORjMxfSu7EeFBcOcMidIhYD0JHa1v+dyg0LxCvpDASHNsaQIyNqJlGA0zug
arLJPuGGlhjSULAnXkZG3P5REKyczbTjB/NDRqkBmhVA8FuBSADjBeLSIK9zEYC/
okoGB1DLBV5VCciIKfNUcixEL4OBbyIr21/L2JLCpoGEeXqpf1IvaJ2JSvpTRiyH
UHs1i3wW5nxHNELdDJIq2U9my3dQr+F+34pZ7NUz6/iQU/FaSAhLkGKT9NTq6+5U
h5s2bcrJKmxzk0tQfjwl5YsJH0mAWs33nQ7BgDQnp9owaaTKHkKHBkZvrXpkCwsn
WkqxZCfHNN6N1vql+SSpD+RxY6sw4/Im/vwxs3x9da4KG7TojG3mV1ZmbT3F1d2g
W5QKQKIOWKer8KFNN2jeG+JQzlf/CMZLjZkCYB6+mz3+CRLJsqbJzNiRefFYZP0o
zFIioVCDBP66haQ4KUYP+XotPf/OZPX+19o9hXbRZ4LaeTrj7HNezZGDitgwMqs8
7q4JvSP5plyC+5H17TUAxWASuyJAo9KPOXtye6+zKIpgYBXaeBhyv7pYxxczc4yj
0+KJxhMKACr52JQO2PibWNWUtko10ZD8R/eSN2OP40NT37u6SZ5mux5ROV0S+W5/
MdA61rPbfuBWO61BDZEuml6ZTLN7SRQSVoeYPQ3yrNlrXYNxRKVvbdUX9c6muYRn
RpKJ0LgxFF6vZNXYhWdtV9AGvHnmMhIxcXMuW8kYUUv0M6hFFAXfVwoATrXd1O0q
J1PPI259K9EwtBIoEk6I6cncEJMDmPPBgKgYXeCqiR7ljZj+J3lnOpF1vt5wUvJm
xWwFks5KpI98V3DFsFfBxTz9FZ+QnPAaV5ExB3jgxz01E2gNF8hDQW7hZ1r0u2Oj
i7dCu4t5AiOpPzgHC/6Qbvtyvie32e+XLWNWG59FSNQCkUySBXQIXPLacSSsunb0
jAll02WgMi8yXezocUVoBefWi9Klioit7BS1V0UL6SW4x6qLyJ33K1TiK0unD4xR
04nmhKqb5vLt4NWCZw23FZt/QNSkucUIvyZH0qNvsiMCVaKPVkHNH3hk1eqnCM/k
MxqqvlMHaCxdOmCb7a4baZoHBomZ99fuYiQh2xu/ugQcjFgEpTdhBfpL0EXxXrvH
BenUd7xlk5mkIH5pXm++ePEr3ahTynB/yWcfRmtyv9xxo4zV0MJsfbv30TznG3L8
LgaAzKFEf0IXDHUxRhGTAbaZHUrcGIgQPTTzkw8KU6EkFUZ3tZXwYYRciwhEEQaa
gPo8iL2P6S+/9y7XDgJP1K/ZjLO98orT/21vGbmNX3V8FtK+sv5EGsZHlCfHL4FO
XtcWEejf5fpC5fsziTNPLLIgcIRNqfMJuBkEJ+YutUxweMrIV3H6jm/tmlQvLRvA
ZLFDSRBP1H0CIpW3tF/cn5pQaV+f9ItDZFfrbgq9qO04q1oYQzEfETQVOWJhytWx
nD7434ilyh8vTdgb+1NypzhcjXitoAXlY5N1SE04TR1/Pl807U1/QS+s3Ga+uoTe
VBxi6lNUaw3OSfCszpV7UnQbKxMkKkGTdUeBXYa9nOlSV+xup4j5XDTuoi6uInAu
KG0fGMJGxwoez1+o17Rlke4Xr9Cch+XpVbNO+IS1HswH0AL2m0ychnqZC3a6VI5k
ElzQ26wghvvYlYXZPpuLWvg3YMQs3pEDjqNqqLT6ncePFc/jYKeKkzgpiGlXef40
+j1HDPJWD3/V6Y72sfslPfhRdgOhP7lRVHMqx5EkyKrlmsiM0ijK7S6QJyvnXyv+
vA+zMKBsAQita7eSEkkZqzGGUF959rwO7Ftnx/sZtGnP6PTa99/fZdpIJSbHSiUG
k8HIvHz6tSpPUjJVvyAsTd0U6P8nomV8epSgXXitLAIXuX+ahTIG2uxXyBrrTS7Z
PDCM61wo68TM8h4k+3wa4xUlemVIH/j+sisjWYm2SfevTmHjfK2KchTe9nkcZ6vM
9XGnV4SsOWcPxLhRsnM3d9yYruQkFGS2/KGnwbwoOSJCP6BKdYSflRsVCxnsE9bH
WmU27R+/W49HBfW8PpCP7BK366cTCMXSausU8HMQwKIE/fOlfYTi+mu4eFDEMKKv
rIKZFQRyC7rM8r9pMN71MWUYZjlvV6OZtrzD4OTeqZE2SRQNhF6xA8CdTAP4ek82
zsF1r64nfLVSn23W34f4L6i1KvXQDj+qTz9doPifPeDzNP0DS0+wgZ5rppdaIsE7
gRm12etpN9J5W2DXti8g0w5GgHoP6AmroXsuhj+xKJMSe9JZXyhyPxqUIgpHdHp7
TrS+dLRjRVDVRS5/D4dIjdB6lXcQx70/AR3JdpvRV5SlS+Wawb67LhrhlRNymRCk
tiLoASs/bV1tghY88HvcY6h+feLp3hfp+VKHOlQLFWoi3qqDIviZA0q20BDHfsb2
RawpTk1OZQXKx/bBhHpxv7Uz0EFCZQIeqrLtyua9oZ5Bv+P0guM/fmj38Nd2/b9T
xmLBSDUQNbbOzi07XOzqWLHEz4lBCTsainsDDOWLE86kOwnStY6OGDLPveSGNmHa
F47/U1LdtQghhDn8+dK3ImThggsxsnFdJJyy89jV707V/MJTiLAJLIg0RdNUIjeF
vybEYaSsP89HQ+UZUIWb9B92hTwsQxin/rUq69e1GpioF63jxUeiQ8C+wzTKJcYG
27xvDJX3nM5yLUJO5lb1wlr0Sbv22V8POHM2IMGPG9lVjf7erNkh9QLFzujHgTQ0
CFkOeTUyUaM6IQo5WH5JAih1DdV6UeGJLjxZm7qq1P4g2DKzoePi9mlH0pgQbYRB
CmrARn7x/iquDVwqtW/LciyXWkigTIg+APaCGdbuyU18qA8BZnA8ujXmvHOcvrWf
BR1P5eLJLwe4mWVk5hWR/evsYR69nH1PWqQ0DrN5vI8FC4AJcDIsgE6hA/nxyAA8
k3EZvTX2nWzYi30mMVacJlcMzXaMKs+9zNzTVcfTBF2qVYFVdua8qQn/uor3KYqR
tBPe4DVVqeHP4my0Dvbgh1pLSQRn1z/EFTsQS8Y33Sji+0fpftcyPR+NT1Ut9r9y
KVPXOXeWw9kfZ/xeBkr6lyjzv+ibaNfdfJGNuhJMPJQwjPYc5E64vwz13mM36BA5
xBO1kjigddWaOl37Vt57DtxPBxM7oiGDiUsxxagELmBvPY8AEF/VIslxXjInd9BS
mWuEMtUOX9/LUIe2yE1STFbXVQ45YLbP1thA2lBBqQdEQ/C7rZ6jIANcO3Yw2mw6
rgbxLLT5HYxy8Ab2T/iNNUzTzWhZM3XbtIIeXi7LIEWXw0OCsWyWJbpN8Fk7Tjnh
BCaYkUHNzV84VBQM9mf9S1c+jQCkqCt2ueP80Ssig/WM5Ga17rNl3aW+htOg7n5p
9Th7ei6pxmMnnaMTtsxLxHD2HydBYYyTG7C+Sw+JzdsHBpUEc31mVYKt1eu1+ysp
OjTWsdWKkrBAsDSpG1P2jCWvDEeE0D9EuMEY2uv/anWJ2TltfZudMJCMWNuL1EzB
n1enJOCJ1pdCcU594W5Gih76JQMITtYo71P3PfZOTprCRmWIwtdS+2PUqQ393M7F
7o1eYLCoQpe2u7vyU8CKU9VxptadI5AbuXkf3lpywzcEzQ/UzElqIndfsuQzkycv
QB2CE78W2kCQHOF3+yMAftpGyaUPVAudXePaduaoVnIuHdx2/62bDZSgL9d8BI+7
F73WzNHBcufqOMHUqe5FJxBZ6EF1W0Qv9w+6h5T2G00FcdOEcJ/jSgRa66e2nccW
sfEYv/T3xgak1iuVLgNX6Y8kP4cW2l9mVgQ5nZjZncgl/TQWxWcXYw5ADt+DEU4D
I+EDNLee/WEKSTTKESoQU1n+3OILe21kix/MdyHNWU+IurMLjRa/TD6/QtABjbfF
ZXiFVuxBTOXQl6qyU666bHdT0vPDUMRCzkTzrh/99NjN2HFMwwKt5yzk4U2ZWo60
XFD3Hpplu+CPK5n7OMgPNA48bvRVQqvHNP5MvIx5dKXwBe3qh7jcMA3QhgT09oq+
lDn2sidnxBN0+3vPH3vvbP6Rb20+1GtmJ0RH/J0uCT+ykM4/h4jk8HW9BgMSrqm9
HOGEckF3mzDMQT3qmeWriLtAGYCHuAuPCymIzdTyeBVb6evqvtopC30XyXwq1LoI
t+bbLKwE7rLDtJN8O6vAEcaeL6ISSz/dxhjGRu2ch/9umywNthhlPQKo94iJAS+3
pwpnE4fmBDJHoAhZ0lRAWKhb2RY1GFngifRf1GY9xME56bhEWjF+Tf47QOorLfZH
FsBwER4d0ONIEsSrYZ4SuZWyn2yZ06q8mDPnUlp53wryJwVNLd8zu/GZ3eXKNcBC
vEtK3mkFgmZyLfzi24PwNyvV7TM/SQT5K6DEzqSVNaz6QEuTCARvJQzLfEXdl1Lu
HVZyGUY4QX7QWNKQcODMlvmfmdwoeSlA75V1WnYSfONLPO6fin5REtnWWH4qclqP
lP5/zYjJyrgDi5lg7c2O92BHvGciXIzoLTKUlg1qB1Saxy8UF4JDE5rSF4KtFzl7
FojpyXEBep5f6mBI5furKCCLZHtQhgUQIoq8zLQF9FX/n/1emvCm3uObDfy3Pmtf
gyxIToF3IjMtbv4MFb1b5TZ58+/3IJ8vdvXRtZh4/GDqK5mTC8++5D6M+jIJirTU
9lNSKHg5TomfZ/86Vw33vnI7xY7B0ApP2nxNhLIPom5vpFB0MKP+k86bPqKjpia4
wvsQh4Z9M6B4gzVnf/173fjGfM6ffXBaw9lKRPhmByOoldIru/8GD2HXjD1NzLLJ
1cY8uWUhMwzMAUuIzgWvQAlFnO6iVahKggNj40WShnhw+oBvIu6+LrJygxlkSyyT
raJCklFaDmAOmznKkWGj0ClkYMmd4g7OpDLo1UMJf5GieeEG+bR+2j/5rBTVAD2o
7NV+bmyhy71qsBAaNHy1cDcyr22O7HQUGzcDPLle+TUn53hBFVkN0biS6ErvF6RJ
fk5/9iMvh6HJsEh8q4Tp0dksBCl7cLkbx4Nzts4g4jDVT/0xlnzJp4U+Uy+AnJDc
t6t48w8732XiW4/H/QpfMIMMF3LqsXI1RpyW727yw1DmnmKmLrn9C/e8XpzP6B2w
jsMyGi1g/rd6lQF/F8vdfIdNJcKPdfvbkT051JpS52LRgv50Y6fJ0S9DFUWyhq81
iZ9nJLNk++n8of5TAkwhsU9cFHItj4kN2wfmVi5MyaeSxJO5HkRxTQ5P7D+59S5e
dHJfQEFDyYOnEjqA43oPGOU8ijJFouxN6OwVSNjtKNbLRWe7rNO04SCrqQbx+Pe6
z7V+GpBVISCBv352q/UDPlSZNFW2Jq19whLhOSbItEVO2wyWFri0JrTYqvKIbjYt
gL6uDzmNz93wkIENVWjaPFxRyXYBB5mBMWYcWSlD/6rxvIzCM5HFHA3p71/skL5e
jAunNSlC3Jaln7rjOG9QV1fgZtjAwxZcfn6ke8bjF/LuDjfBLDLiiKQzhPhdFZqt
yA9AJ3ar56o5DhGwBya0Tn+RXltXApEr2DTOS8SmhNl91NJQx8iwwMo1Bf7EkM4T
W/h2CpHv40gh55wO0Ruf+99DwGFwldOgLk55SuRLbra9CK56hksp0A5yFvV7FSLR
MMW933Sw8VELQv7lObVkXwK7xhO4nniwuJCnMuz7KHbEkbzk80AtcalZExZXtW64
cln1jwEb3k1Jy/lZftB+EHjR2Fqg/A8upNq+SqMFHzvP0OyMETaITJc2GsrUhcOa
nm+k3d9MCD6mxMhmT/rA3Q4Bv98x5AphMyZXWkulCPttrTJ/MGrEcIyrMjli5j9b
09mmj1q7og+jLb+6vft7c+RzRz9BM+l2i57YVCgR3LqCjMpH/cTGsjXUGyb//gba
kAefuN1rlvncJyf+u+D+A00SYPmJoVfCHQsAhRB3QnrVoPrP5tFVkGWpw02GBq/f
J6ehmdmmNMO4HJbGDwBvvms2VUD1Ok08put1u6Smm/4dYbu0ORF4zCs/C2Df1WTO
zMonkRpDAmKJksQSyjOBYGrUKDJy6QJCuMDzYrKK+bE40lMN6SyNZbEosSihkj6u
16k3z7r7473OzC3MU/3brG8oAbMmDkqDBEgvK03w+96hgIgp0ZIbZ9gjebAFqJVW
bUOVWODIre1VFYln85vMLqWtLE51MMV8OdBZfp2VVAc8kQSnvIeVq4lIJtHsfwd9
aAZpAZF0/MIz17xi4UZZxwls/Cuy4LZMsLVNMBPY9SLQkoVA51KOWWCzK/IbsEAc
D7J4Or2sHZJ5cEreGk9DQNub1KY3ojvwwGTGkYKAyJHRxspLbfsg2tZrDuLYKQPr
A1+F0sOi5g/756BqWIWS3tQDIW21PxxeL7hshgQPHw3f6FUtBz6gBqHob+m8qaE2
icLyXyHaG7lj4hEFIJA6TLIf3amn6nUgXyKiLCiixJ/0dGooVsXu/2Cvp9WNS6oA
ijBi5EPtbnpc2p7uZluXeKpfEsSe7uQlsSKpY8t82KJjSqAIlbeJhWFYpgy9iuat
I+TG5A4Cm0CnBoc3+OckPVVOMSxAFTBLR5PIut9Rrsv/jN+JF1qkL4llWZxsHquu
aQ+G9rTQzwoXFDXfj8e74xzwfmERkSr6ChHGfwoOkCQqHR2+luRkJFUzjiJ75slU
crEESz/nWWCvY8PYo/PAls4QrUFvy/xkuCIcxd1bJcxjyYQyI0/DzFlJIPVI6QWd
obRxs31d7y8h9ny0e3HchNZNbD+clVkZO8dRSaUXAbNpfocW8ROhPs81imiF2rGh
6woP8Zn3nb+GBzpEmAN1um77azyK59qTuAYaqrYW49bqZGBFmPwyWoB67WrXm/tW
YUlnVtGj7stiNRGnrLFUWodlbRf7w36+uXvlBp+sMOaZ5i37Z6LFHrF+qasRwSEF
39ltGf+ruIOLbuBkgRKT5jIb6rUWcPwvAMgguELKpHvHM6w8bTwXrzcFCwMe0Iwk
SSrLfzq95+1IUNuH8q33qQ6x203iCwdPsgCUwqJ+woBhyptgsydrBHTJqC5FQUCv
+q54Zta3309aS1DHO8T9LkzpjRH6vu+8KSPFIZM6+d74EA6vbVW1ub2P2GPpfAy3
JO5UYDrvWgk8WjU5W0wawpkA7qIehS3OhnptFbTkQY4lM95okguuSQNDGD7V4DTk
Ct2B9+VPsN2+ijwg6J6dYs2JN9AmFwQkRrwD2BTzG/vQ1UG12MkzkM7MPckXbyOy
LxXSwYMuc1keMMv27cStK0tSGtFonyMEGgZam/C0l4xZfzxEy0CbEc7SGE4d7rAs
YA10A+p/YukHXlwr6M6jOvzpHpJdkPBAHjzvgQ07e2UrB/FeTytj4x9Upz3zmfiL
93YlCMT+3F8/hhxmjeJdjNpa1kIk0BQmS2gMvZkjKaS56bjJJSdY5xZjpjn6rNtb
Vlh8p/+NvbjEi4ZqSppi2I3QbMk66Ned0od40tUBefeLwGfsvlcjycWqfHwyby9W
socbMjQnY0y1M9ipufrxjH4MwaipowulCVl+ClrB1ByLc7HU2M4RUz738R2kG8SP
gkJnSH+xiKZFIjHOGPMfnuDIrzcny4YDzZLd2KUVpgvjGN+QQEX5SFuFF8d95Rjx
rlnXyHPftGKua7HgTyj7U0utOttcBrjB06+hkfEbprsu8Z+jLV3bKyltHdFpZ2NE
Q6YDXg/HcMYrGKSwG8qGGmV8u4bzpVrD/QHYbb7aLB/BZqlPAuBiM/2eU8C2KL4s
jfaDHC0w7iEE+Pxyythr3jUQf31heg25NDg7hQlplbFjJ6XxUUC1EEj4uXP2m/RF
OEDFBSAQk/qsxNBrzFOcastImeI1PiAkccr85wrKLXrxiFv0eF18nD0XOmImy/2B
UzlUHua052CgVnbiUEyD7R6zBFMQZFsdaFVeroKQeSXKagCBHIbscHuTERM2trML
uQiyEmHBPkSFMISPwo/2wqacm0MH1n/uN4/FnuVvMd3JvRJUbcd+UvE+SVzmjiS7
gqHeK/WXFH7D7iQblClYgAYyadZ1vtqki2lr5yqGri/54Q1FpBh+/1GAyoQKYA2B
P43h4lD0bKbl7lhJCXjZALKkwoJo3kofdJHE5eVb9WvJZqxiieD5OuauiMSPOR4D
oY8c4E1W4+mDEQcBaXkRtP5HKwcTnlXIZ5fd5lYvRBNTHLB5HnQF2iN+ry6j5S3f
wmQF+gTsH29aMDlP+DIPItvzXmKl6nyZGfzbngPuCZM9y2FvVD1KshmykL6tcZQj
rcjQTO0x7pQ1b2ZLw0XDxXyUf8WNQXeXWbhKSXDEXIGYjoM6fdzwz5bkiRqsCFG3
0VYc1JsxBsC4Ig5C0CXDg97AF2Ci/HUKE7hD8p9LDagp5Azt9QvHB30RzefEhTrh
XdDx6el6K6Cfy3Kk8L9lfu1YHihLG5y3SBxQycGKZMjCyRK/Hafb2jOpx/I3RGCZ
EJbnYauDfm/FAk8Otq2XLgFl1QI4dyrOpbTEkUSv/YRMMyOGeY6NCMhD6HPnvGeK
I3Hvb7Wm2iqsSlGGbnr+aQLXmkWAp1M2xH/7Hgh9T5WkzpRtQt+jRZLFw00esSd/
UzfO9eygBYEfQNHpQ6qcZXSQ9pref3PzKlpliWqqUkxsSw8mzzJ9XR17FLMhYugj
bLIfkaYoZbw4CdFf7WO7oity5lDCZ7gMMljMli2zmxuJMU3ZygKkdqlCxGkGojR1
2mvUeRdqGUPdJn8+Dkln3d9n2VblCGYGevCnoObPdwlMSH+LhaP4m/zjwfJm1pQ2
4fOEXqt5qdCWGfM7ZUbgh67cVPfcqACe514fUbuRoXU+eUIdEdW8CKdcsX+EWGY+
JkxsUwcWL4o7xlKBm55m/0a/Hb79ku80C4CiTXO9N85TyUtMrit0s4qN1aak4y3d
KFF5p7GVcpRO0pIFoUrox7HacioJ1PUKFjBMzRJHjChUxPHredxXjUR/6RL/b+Yc
TNi08GVaoPJKlC4Zs/WLX2kUEaiHQ74FSrmvQbcMBjN28ceoIYd9NBi4cQsR+2f4
YTWMAj+JrgSwfYmW0jSqD2rwHSOqMUjRVABAeAwZJIzLHZ4HJUMx15METQhqfza7
47qYi+7k3ISMR9KOUn6lhMLmDyobhiRRAcnzujLwnx7wqdKnz29C8DN3kWiUleKs
fEErxOFTtQ6zXm8JUffejk5CleMnhOFOohqspEPzbfL5AFpY2eR4+tv/fp8V/25H
/iWSJH5yj9zU4zDmEARuZ2dZ1OJdTFqwN+/mpSIsAcYnYyTTXKJRmBe6cfi3PVtw
IU3Zj7u3ZlUyjGGkvFR/9xtPaUA7IafuY0td9bAT9Cmq4ZtnEQTnuijg8YZbO2t0
fMGSpeLAv/cBSwHt1g5/k1bKjx1wnBGJQJ+W+SfQAK+sKGn3U2sQIlBsZw4rafx6
S1T+82JT9r94NIeUCSB5taeAcuSF9eCQKKX4jLPou/xhWt46MeOUUpcO5klErQne
buiw2TFhw/dHNPtU1Y054BlW+cSRw6sukedr3m+qooHRVenPFOJGu4I+6Hyl9LgG
88ihsJ2IODg/0jtQA3I4wtZZyLnBAVUnhX/Wd5Ll9vjvmG2pi1sFr5ka4k97pZRU
i+5J9RAqOpHc0g6Uf3QGCPfYjGNMmqU9igwjRG2VMY/BjVZKFbXAsATSCgFRDQTu
owc+nda69PQK4NjSv0aKy8Y9OM4HhIJjE5vb4ht6aT9ycJwcu498smTQf5Cr6iug
dXKaGy7S5zXzA+BA7OOE7+YcQma5k3uH7z4IrKfpeeIjYYD9BZVFIsJ+2poW7bXX
bxuYiUFYnMIve33RwDJPs/SA0c1qdIqkn/FD7amU6fnYsBSa7TT9sFNrtOXmXfC4
PMgbnXXEkFS8SQNSWjWImiDAzDAu23o7wV4iWe2wBGfE3HCe3ma7girJGARtR2Z/
PdKuH6v5gaYxrJggK4Jh/D7HMdUteF/9JuKkibo4MrJZUF6ih3+kXvOCrx7NUEQL
POkk5bT/6dN1t5Ia3LaGYMVvPaPsqPJLUYeecjvPBBVX4/tFfl/mNm0ypqDq9jh2
0WhBuo/07euQdosvKhWwu7wL89riCRQVKjOOyOLUD6ZfzBvp7uuj0Phw5TrqTQSu
8ARJSO80L4Z9Tmixl1ks9RE3r9vJjfrOIFtqApf341+FqNyDA7WnmDySMhgZzRrf
fLqgg5/Gdv+yn6IrF5y1klXWatPenVyQGoPbdjTJVc7eSe+KVoT8hZsMcDvW2Px+
8xxgnbYKrzu3YTj5XQRYz3zLhlN46BoMakrEYA5/X96M5r3PH10jvF9+HkFQKJ6L
UmmZSmlc/XhKP+HAivN8P0sDSTZ02XtJkJWUpfUvVIA9qATy8NgFaMHzmx9jwZit
/3/la58JIk3JlkVlRbHQFsWeKaHaXCkQXalUzA2/YYW9GGUEfHi+LhHv2uPsThqq
SCTNs/+It10SvDkh4aHkNahYYM9uJTOvdtE5Je9HdX7MtCd1EqaCAWSTmQsreW+d
cT6sj9zqdNxB2WY7B3vHYJ8xsVXfgg/YsUb3vtcJ5UsCZjw7jlO3cF8kxlVVObV5
pVNiMBTWqCPzZZ35pQwham6Q5BAY8y8fIxCOh4sPos/CB/mYPnXv2dXwHkZXp/UJ
bI/W4iMeJbmj2KAM80Zlb0JP1lHh6+TICjJk/TknYPKXx0JbtqpW9go9WvbBZS5t
mm/mkQ4Pk/+nHz+FYmHPvQq5OE8GS+nOHxATltAYf/pM5v60sPmBcn2s+LY5VmW4
zjROWaDTU3iHolMs3BBpNQriN6+g/3HO1WOzt58p4st/YlgsZttMUAkeOEyg7DQI
yO94h6ze+IC7zkBrpDqptuL0EoG2BxACOzsLg0btnQE5MAFjcPW089a5VoKmovkK
LaGjCDW0FrazUNO9ZUFTo68TIIHa53RBc4k+SY+yD6X1F9dQCITj5H0+i6dcm7wp
kepCs0BYhzLLLuCOzWtJ6v4PS6f/RRKtiuXpavRhzVM2FaPMdAky8tRDaq2dVcwL
VgMgued0eMGuEX46DG4AsxFihY5lOeXlClpRXuXCSkinL9Z0grGB35Tj5jB5ZGok
t1nfO1f1S/yhE+dRhWSB1230Z88C/xnEr/vOR7CeRq6xX0htAZInJtp3XDv0Gs18
5nG3/Has8NSCfGgFtyo+DMbUy8s+VcmJAy9N5PDRqiIKiOKsG0hZME+va2qjxbwQ
D5o90q9yE92Mwrm2sOoKZjWei6eEHiB++NiL6Sc94bFqPGYq5y4xUWobGXeGT/27
OJpEeY2vgTEfJ9zQECMnTUEN3b1lEIbnzCryG/jPbqUIxnmetjZKZS3FxI1seak0
xfwuyJgFoFkOz+FznzzLTeEMO29h8Osee8RsbX2O9WRxoHk+DG+nr1IC5V8R25JU
wL48xGJbaF5khcY1eNWVm6sDhdcLNhmOhZV2sHonsN74Y9A7sck4sBo0jepxwvnF
oaudd776iz0v/kQTM99Jxa612stEg6tDnLiPgV0gn6/mnwtEbqHf2I7VLpny1lQ1
OZL/lz9D5N7FEC+PlVCSd8O14EtpkokxTB+bQXg2KVRuGnnTgWzENoySiFc2Op8h
XygyeZC27TXseTRSmzsYbfd7l2GLyxCRHamvS0rEbH9KKoDMSvEfqZFo0Z2G1C94
TTCqQcx4aUm9YJn5n+UBGAo/bkJIONS3Ht0v9M8XNSatj3N8ftOLBhr1ic0HHUpo
8UrFXGZ6tBMc0HyG2cBd3s8Qp7dg2nERJGRae5Ej/XZ8zNecdDXjDApj5+slUG7m
3iitbmbF47naIu0STPnZqCHiWn6m6hSG8q5PURp+x5vzRNKzC0fOh0pSMA/pMrmX
oge9gKh1PM2suZpVKoW/Hfa9PPwxyiFqok4EJ2UZWVi4mMPm3J3FKyF5fUiraUiF
xtLg1udLdLuMWBvuOOpwPeh33MjWwkRgFsf+7ZtXpgfsD1eWq1xml7c6Q26jrR37
OWFLD8KuH7xB09JhkPloFioD7tNzGFC/LYiR54Tl+inqcok0nIThfzvRzegUkapy
w8AvhbMgat+EHkoHJR9agdkRvusmpNbTSCDKnS4evXxS0uOEtNBx+GyQ46dDKH5Y
0wSMXZsHKYPzYzWCPaQ0fh7miRpgUdZON3dmA/bzSXMydFpZA5rbzBXGPRppT471
sgGVRhmab8q1mxT9x+7CKUOSj/1Z/B+z2jrCkJ8jySRZGd8HbVoKJUzrf4aTiUE8
XvOaE6kl7+NIf9gcMTKhD39kSfUHN8d5JBjdTufHSvvwiGPG5GLxbcwFbeQsK1uU
prBhTW/5WYK0tlyw74MDMQkwwL6Po90kA1Ux6jvaGQWdnbJN/VypfI8MQyjZ2P4Y
5ZJpRzpBuCCgXVojcO/7W6Hpl54lbjrp4t7oVJ+hY1n8vF4M7ez+0LOG1riLVEDX
ddMvE9oWPTTgLblOzQ5kcRIGLHZ6nxQTapLmyRrTykHqheHndp6v8idVTFiBsaqI
CXsGgEnvocsPRDnGAAmzq1BY3JWmdqxxLBd9kU6LtlNi+YnQSHlRnACWx6aYvuAe
QvZJCojNR92ub0lY5zo67tC8RAWbYw6p5IijpTZS6bchE6NOrXSHAnPw+pqMUSeA
3ezwqEfgBkBos4ZdP3DnQZo4tbVQCnpAJlRSm8atSu0M2sB/1B7E7Xx9j4SnnhoG
VCjrEUcBhGyP/O8vnP2VAXx7xzdoCbkj180y20Lu4QH0zd2jRN0gCbzNA8wxzpcm
ie7gAukTWXcoNSNuDJZoa2Nooi3Qh5Amvqqcfopzv0bmf3t7jco+rof5RFpcGCsy
gTzOFcFpw834oMsHYLWNuKiSZg6Nmtc7KsOBiiEWY4sPjYTUGgWYJUft6c1X9i35
JTj+EP7IYn7Owh2gUTGrMnbUiKHGVpu7c2jgA8PoyLslPrZrer4i2V9vrwZsYXMC
dbD/e10Q7sFtsy5L2gp2wKcFawmn0PhANZip7FXP4XXmYHzNc0dmG5hIllK+ExsL
Y7yiOcc0p90GfgwXVfk79EskUhYWDP2VKMpVCirsmfGbJFrGU15+oQMYDHuaFfw5
UxG4l2ivvoKrx02SV5AZcWPE3r2FLuB1C9xlnYhUKWvikcLuSUqUyU+LCpTR5ThL
5McO8BU9NclhFUMavDIkZaur/ZWpUehBst45tEcg4I0R3qhSE5q/JApuXtpiz9ZD
Gjt0WJAlfsHP9HguhaHceGqYYGmm8j4f1rKEPt23pJgbLFkm4xN4qcJjxe2iy7Ax
yfOIq0YCIxw6W8HPRuTWZivEL3XKl2Lh+UySFfVl1xx8sTObB1RcrHMbYdPmdAo6
jRaAz/VZqaMUD6wYvShB/V337TyJmYbLPMmoWwSlp8esweHF3EafkvVBSttR4sXu
vR56VNfLcQCrzNS/QZEr/IseBGdUY4Co4k2LWOiZK0c36T5m4fIHuB7yDG579LQf
6dYQxUyfIEexFizOQK2M48NkKJuF10GUuCnKZC0bw+OenClH2DIyjdzhD8zFVa3V
8ac9gUnPo1XBcl6acu2KIjIbDucHgOmwAwS6gfK/ncWdi9zKOSpXZ7+h6j7EUPPH
dMTbMNWpDAHguZf0BSu8lpuuh7Qg8tQBTlf44t0oIMtO5C94dsUfCHzkyq+QJgI9
10ftx3hH/FUp989D/HjvgMqLJLL05EeSQYnelD0rNfzHoaWGVutnsNG/usJz117z
F5TSSzOZBAr/qgZNSuWgxf8FRmoM0+cVHVrgeNc7GzFMV/FPAZFSeiDUebtgKOu5
RGvfav81ms4TojVirOD/8k/UVoT0ObQ8tP7f8RPTU1EG5esZF/2xfb6e2u6HduU8
CIzCySZHglk2qK0lMbG+oOPRCOVhKRcPOyyBrX0KIhappmIqaHiK8SRMg/V7kTwE
aaCb89zAQ56k5Kq54PZHpIR1pfUynshDdVFiU1oFv4AUOLmfMtuwFvIH2StGSbyw
Sk4uAA7hNrRZN7XRu19Xci7f6J0rjdBfgemC8UoF8iIqyzqFLB6lNyyHUVBgbkSO
3yioRrXchaLx4lFg3IUjrJnQM2pxLgQ8MPyGqp1GJHAxjCZ8OpAmZK1OHPXaS/1v
uNjjnQkSqeqdV+xHEdBjHWAGs/At298VvKiayfq6KqxYSEn4bNhPsw2QLHkKt7Wz
+AyVd9IPYIFUI+qsM+7RoWCKC1K/3YHhqmhpfkFKxWISyUG2DQyPV8doK63DQMwm
PlGq38tE/zZ9gwex1XSY/DvQI8yogZQQJP5YZtXgOb9Kzb2D/z7gNrpCEALa8YUJ
aLmDfjt9eVgdXQ6VQp45bu0BCSINbe1zDvBSKMCGld3jyxLA1LDi3Lb3Cjds65Qi
cziPha8aFzgGaSarNnrCgoq4xADNXZv6kkcV3ouzCrDqoJIb/X6nwqJMG30nDhmC
xAkCiO+zhrzlgLHwKXkBCcUuZFf/qH4blBY1IEOHrPCeH9dvwpJYguZ7wzf2UZ4J
qI/5ULtFZvynbLItCYgijrWRKRbuWZoGjs8z4i1WIPeO6OMHmfCZ9l/KmiYYBwKK
dMQIV56OzVzwc9a87wcFJg7gz9lVcXgB85xtqlywuT87TzMjZ3btJQckA2yHeU+l
t04HKSdGY4pr6mjaJljCSjFI3sbCcA5sl8YNgVk2XlxgUpwNEHVcUX8/MOFItJlK
lJassTqKVWUp6WzS0J1jcxdzn42L9Ri8Ub8tHeNGhekmv935wljNTLitch8Tn9h+
SmDC65yvn0sy0Tz9btqqhGFtezTi7h9uFYcU1Li5CUohmpRd386k/pNlzr/UHgEU
UFoTq7U5Ijca4VBn53ylp08juPsLK5+CWHdMhhpwPIOKqfKh9BpVMt994HF3Myc2
aKaxdTgPeGhV+StLMDfLG84nfaYwW21LjWUQVq+e7IzYRt3YpVq71Qys2nL43A0a
81rXwqG/R8ng6BIO9/Ir7ww4INKJNHg6W6OoLQjcPTB70YM6TnNcBUzPDlcpAEMj
DSWiUmyqr9JeVj/vk9Li0aBPg+HJ1rlvlHVtcWeoQV5w8GePT9QueMeUxz6zX6K/
EHdkwYyvFvV3O6z0brO2XLAG12seLSOc9Az9QT+c6G9n6FVeZ3McQH1U0xQHNL6Y
4c0Noypmvj4UXMT84/m+7XQkGGNV3h5l+bPSWE++6notHPAy4ARvtw2I6rukc4/H
gMrnzyPzoqzDXeOIPLqrsmza83mEvBq4PcHXdt6gmOdigkL1j2P/QUaiqq3iARgQ
bgacKThdPwCPYNG0q42GHEPVJpHCwZPmOzFM75VU/HXx8XICjwEuGponot9jqWAP
Z8jhudrdqY9kHbeGiI5hWj5rxhYpNDG83Me/8QR/9jC12jaHXC7BQSxF4wnZY51T
WLd3xJTZkJfW2t9juKpXVX8Awuvav+YHbzq1OYhuUlTjv7jFy1YWkU/SC2zr21OH
3QT6wBtot9QBfNUbn7oTGFxAawok88pQp+qQ89L4BgjOErK3hWM60gI5Y3r0MNDp
o+Tblle9e49asWC4FIwvQgHCvZwsbJxR2ZSa/huW4EOY2gYEK5rmPBObzPkBil3x
Bkikn1D/6J+e3n6jaH1zA2WhLfmqWg0/poaq7S9nt8BbMwiZjtquj1YZ8XkmnLs8
odRVP1Q8wWciTUNKOkPpjoeCv6EMer1kCnt/RJfG4S23U+Ij44WioKzd1tTcg1G2
em+7SG4BHsCf8TOcT3iLBC3fuh/KY1tIWagRsox1CwzkYpqHlaBNunxmJajMBwVM
7sao/lx2CKaX0bsQz/U7sjlvl+oo1A/uZMyeH36RgpkdsIU1S1J8TZvAo1Y+hIqz
CexzPC1q5rfNvwQTlKDA90I4VoyATCg/EKUsCS9y2qNGBMiT8qquM0d80FPc4BDb
3XPuyZNqli/K0SvbwXWB/ZvuuK/lEisDD9Ed8lCmoGMiGdGRegM3s8kYcOTO9FQP
L2FMJA5k0prViIxslv6RCpDtus+Yzl3RvKOjZwTHS5vaavHRcnL6hsdRIzT5U/Xn
STBKWtpSKdGDFDokas6MjABZRyF/QZhRixkfcTjynL7BMy3sS34WLWrMyqAfyvtG
wl3khn4yJhD0dF2XnXHrMa/7ESx7qjIH1HkYnfyYF3ZWu3HC1P1zB0T1+jCEW0Z1
CuhbNdd8N2cEIaFHoknv2Plj00NxZFAHwHXNq7pdGvLRogn7pQRqaPawOdTjzklE
TBsEUikifhj86+L4GUOD5UVywy5P7l+myqsbxsFLOzUNh6O/PHBfDZ92kGp2769J
fkpd58PIAo0sApZ8b/c11zjMAZIfqw8Kq2TnqFzroCe7n1eL7mwxgWr+TwHq5Tx4
bSBF+Law1lRynQ9VOo+0CivwbBzoRizp63ipkkchTGLLIoXnJlRcW9+k7M993ML9
Ia6gWKiSKNjYbpA3WVNlxpVA0Ai+Znn9t1xgPF18F5Y05a7iev+YKhrqprHVfQXI
sNZUXzmrVXUawNuOYrny8zUXH3KFkRvf2JZ4vgKpLNWdrHVKy0xvptGE7U+6KfT2
1pDIXcse4Y3HKPAmdKJK7LWOV6dqps3vMVjcD5GkRqiUwX4alGTpDD3SPCRLVXrw
J+eEUroJ6X+l2J28IwYrjL+AabJpbCggi3NmArKFzRqZR2xxIStb8s2tlcrTXftC
/2rPIzvM0zclkUYkFjW5NL7pRJXMHWZvnlsIvVOZMcqLyMWFIR92R+gRJd2vnCqi
HL2dOZYH2YLxXYduK2PzofnpVip19L1AT34zewme8C/7jm1N6qw6V4kEOwpu7Rhq
/6r61IoApmnuzBnAQ4Kc1vMzhsxh0TEwAO4QtvxtYrs8WM/jvMsjEOVXsHcWgXK9
9SUHfxOt9SylZeWqoSgsI534JdqDyllu2lDpmhexX1LsBBgRGUwP1Wz4ApM/1u9j
lUCisH6Ln1cTxTWFdyaMiNEpbCXC7/le3mjmqkK6tQ/dGMlqzNB4JqukiVkEdbdX
AXFllZktK2M4785V0tUu8p23AtDEFSb49v5yHtRP12QIuqzop6oUZ5/thTLJxa2J
7w5tp8+CBH9cA1N09BbRkw+mE+Kjh+2m0HT6TKleuPZwRDM9jBbO2q7XzZkS9fON
Kozlb3rDDz6uJ0a77n2tlpPaTvAhCbEb8a8mYdib4KpYjmyA28vlX8jN6Nx91bGH
Pq9zJ6+hlMmg9G/j94mgnPst1hIH+/GjhGc+uXPcw8Akik0zDYNXUAG5kYsd1Im4
Vm0AzGzQG8seUD76H8qH42nTzAq/XfRoWLe15Y0/ObNxmCp3aUKS64EurIxez6Mq
xGcKDezY6E8isPfzrANQ/DWyiW9iF55AVkrCNj/r5++Vizl7oJ0l2KiaMywcNaOQ
kKRTPd9bpGoJubgRDUpTJYYGpfi8RMl9l2DpWZdv2eMdh042xQAThwZffXW1usPS
HmeWZRET6EdbAUFyAqbh5cIIHyA+ZCJFL3BoTbTMQV2cR2dH2ZoFUBBvl4jE8A9B
yHTfW/tSFvnI8R6X/KilwoCYxFOvAqX008xhJn/Ymiq/ROb8BnDV5ph44BcYSPun
GBqgmX88CjXcivN90/uqfyyBHDgXTqNdZCBIjr+8hSuJ25cv9K4Kh5ykiQB21XIY
p+th1JwHl6ZNtlK4OMzkqfh2qlMvF/6NOKfyhcdjVOPOFQdIUhGB8CPE2k9gOiaM
x3HfeDJ1Zz2V4XUEsey7UQG/tlQN3Iu6blFh/t/fsFmRBl+6tSSP4YZ0+DJzzWrj
jRmgcmc+xiCfyH8IFSe40eWn3BdaJjkcsmWAAjVa6pW/+eD82X+RvRAxT/L2rEtt
A7+y6bHHL6rXPnjqQ9IU335jwDMwyCEDzYNA7ppPQ6tocG7Z519tS4hxZe+mzZG6
UDXDP4T6P0lYc5FBpZnI37LV4ZiUfWoRx90zLG7dWyv7Q84EZRQEaCpf3cFxn01o
lWpEWEVDk4ZVXoPHdIGdfAKlah1yLhdp49Ox9xwMBjWPqsH6F8pyePJm4g/y2bzQ
TsL4pY8docfhzxXfCbdtSfjrH8dgHgykkWHh/T07FbEOHygEYBZ63woJLjqiWWts
jR0XXnvqNpeqXNBTAvNsE6yYHtscMYESrec49W4JRMC0fmwFPIb5tHh6V1QJS0fx
7Tz1vIMTjJ/mLJSxTQQk2vIPPBomZYNoI3CRToKD/RHJ691htYQHwHIa0O33Lrux
PKCvuG0oNY5xOeRfEUF2O66g0PVElafXwcAJIUsKk5H4+Ck4O2UJfIH2u3DozMWI
lNJpOhEBv15xGC1qZFMUAGEpDdlGm20pDtSjlhskXPKUZNPUrhSYKQ+DIzLr0jBB
JY4olNTo0i2Kvn67PZT0Mn5ba8ERRRfD5wQVKmujen2cQ3l1XxzKBC72jvpZFRrh
23ChWTo9J8DeNWeZEZ1d47vko/5WioMykM+antdsM7hn68E5zpoOg3RZWnW1/uKn
NbPLX0Ixi7MdgpNsARe7LeJasJmph/YPz3CmtmLe8WvrYQ6xKlIV40gwJWkleYqw
Ii7vk9WTNI33IpbuEHoBSjeBigiKjmgRbR0C8Ke2SHwLEyEewVFxkAB6ga/8YS5c
WkkqGvD56Lcz2i5h3jzsCoCU2Km0dRpxeBvlXaHLJkBufygkp0+81PF2VlWpbwfy
bPnQk8uh03+QTuDvMkNezPmzQtl4orxOMhh5PSQy5cKE0dhOohaDqPm8oEdfM9sZ
xJjJTXnPJvNUcRMxyl97/MT7m2ELRlCkcyjdtRsmhQa5puFppDFDFWhedXN9TH9D
QPEeF64/CMn2Rp9jB/02GOZ8CiVbUgwCEn/jdJkmAwli+HPzvc7tq/b+CY+BGP8Y
eDPfzNyTzMPLOGnMjtNNGP9/rjHl6J8KkfZG99Xw4+oRRlZhuMWOhQLqQaGcfG3B
BWzN8KZw3uAXl4zVlfvb+sG2L6H+CufBLtiEN3kEGxZrHpcG3t4sU+qkSro+milN
U0SIZMeppvstZtEsRiEKa96QLlj8K4DkTiGtcOl/Nz/Qbnj8Q1NXXYEyExFj6QcV
EJEVlDtQNWaWQMy4dsMWb60QfdqKFRaozhXsNOPtI7thMfnJ6MmGxMXahFPXo32o
IySjHADeMaYC1OBHtu4ISSxl6AJnpCULfLXHjx7QxNaXLmDFli7TfbTv35uSfpRr
7c8Lin56ZapDcCt4NQyfp+QjcIwaAcuqqrGB+cJt7mzHagVobEBgW4ji0V2DftaA
46htwafUfAIyau6TKj0vyOJ33K+TX2d86rAtTE5KrryBpMkoz/skcEKyUN0lrGaf
7BYVnq7TR6URAYyiZTrsj0zaSuyAap08qvBS2tZwuJwl6OoNlTErlzCzC6oc0z6r
DBxF78tPn9u++27Gefgz88D3pS1cx1DVN6MIfNAkjmLXUmwFHp8bW05977OvXI+R
vcy3tB/NnKQNGiwe0bFxw2fFY8i0hEmpRbGZTseFLklayWHqpov0pz6wUpmvx4Z+
B9M7l3rlVnEnHer5ZrLecNn1MxZBPQ4tPcadT0+lcwi5y2CMHM6sY5ioVHElbOek
P0MfTibE1jBDCNrJYVka9/fNgLA4TDXtaDcB9RdYY2U1dbkainHB7l//wntDIIqU
KZEGhbJCj8weGsImT9RLunWaNGwTwHzeUyG6sRaq6GRNv/7RHAi7NxmMS+sIkIMP
WExYL2oC/ZX99/7edBoZVCLQVzclTIY2H6AtBV9UQD11Jl3u2j48G2SunfQr8yDL
RvXDPb2X6dwKTBdFMst5UJrv4z4cdwOky8lgZmI1VomroAdlixdgDzU/OgEijF18
n3IGiGn0CKAqtdpe+pRhX3lwQbACkFcdsQ6vmao0oSLLuiTHfrAViv1iQM1UCMl8
H4dS2+m7pvXpARRHbQD3au1iTv/Ckxvt1vGqi8kGQV9AG9q9sFBhUluEMijA3n/C
0JyXfjem3Zkbll2PTWko8cKJywK+53uoGT6QVu9CKhwl2jQn1S8BTU5x+FnyiG9S
fr1q99OscZJnPjpU2aBcLELiYfNiQv53aTmCDiNGlZxW4SRrsgeS/phlGNbHa0nu
sS32M6wU62tugHW6Vnc3ci4SbnbviijLYMdrGybNXtxMto3kRN7RxPoEd5seaDUq
ukh5safVdlbwZmp3Mj7FShaBtRwa1kA8l835kZU99bFLDoP0PyINN4u+xSWkdJRC
9zdDw1fOrxnq6aEKOScxIS3kyhzuLK+rXavhzEYOSF7WJz9Qo2/CWCHZ/QWiyjxp
3bZBzkYmTuiUl2w1mEz9OBu1UvvL3/IhvfcK1tzXMIZZSzgLattcZfIT2QQHul52
gzZ2II/OhBZoIp6CPmyzrp9F8+pZh2lb6B5caJFOmIWZ8zRYsdZLxn9AM71E41bA
SngLgJXtq+iqtSwqyd07h+m/uBxtn392OEiwp1yJcGIkqMD746iIzq0Fuv2ivzll
cwTAQ3k0LUCPdbJ0W53DP2oS/5z7GSeAji8xHqu8oZOyTdZhpzglbvQNa5kTPvq0
uFC21NGaejLL5mkI7qY+BU4LMJIcuQfcHS1C9LdJOz8V6kZlSqCxXA3TFoCtCrX/
KX0CiMXkg96YyvjWkPJKDiv6gif2/GqCoewJyWopuRNeCLIR1SN4djbjM5aWVx2n
AWZY6Sy5bYmqfxNXYdb3t80z8JF3MBQGTpm2bjkHL3Tw1oQw07RhoNBnyvNvF/Gn
UJ8uWcTGiQyQlRyuPu62DSuPfjPmbtdo6g2laY2PNU0XZDwET0YRWVj0e33maeq/
FStKK8ARuxZKYJCpCVEnxYyAHXCV6phypIEIC5FY0uft8sZwihtBULTxHH+XQuBD
VfJdKaJw/xWVb9n8Nua0inOcVmqZgCWdY3aIQ4H4MAjXlbdInCkM5dZEtRGDb3ym
NaAjqwzJ1sonkPjnyp4c0hniW0zVTEf0gDwVXPFWzZxO3z6bYs4desUjhxXs6BvD
/YSrd2z1CtB/xTJKfZaoi+rLBIKPEyTIxGzalAgZ0sR0QlzZelVRmHT6iv0vCSfQ
PGcpI60ssdJUTdcwTBTgcOLjQMveBppXfwQgEMVFEiQs5C+CN6o2436W1cb9/ZRM
6OFEFmE7VB68rmEiHvsIWuGMgmCuzLb7f1AW1kSXkLPJNcEDxKrAGc5OWo2sF9Ss
cCzSy/GKNX0lhUKEC+0tlMPn/q+0cj5l0nnLBuxQbnMaJ4OA/lJHzU4TOUudmUxY
HxSEQu9nYJ5ZQyjr1R7t1R08yUN4aeLGPEX7uLSOW5zYMgy+1ZiRM+mZJJ+4Mz6t
NFVI7QTaHoIxjDjfBtO0Mr99Pzc5PXF29zh/DZ2WnBCfW+mpzt1lHNiDt2Lx7DEx
IdGdpIXMhL2upOHusne0nep7ZjoMKvVaS3FqA9QiF1GfrXkKG996NC56Sjo3fnCQ
CmMWlv0WvkhpG+AYar1VwFmo+GZ+/8wmEsstAKcYfgJocI1Y9Ns3ikwS0amCVvyJ
ZOO6P8n7jSzD9/Q3x38fr1+yvjCkhs8+HGWd63Oj9OZ6UyjVkyognnVAdMRknn+P
bVZg/mXBrv5IUN4nUlj/G595b8+dfsVhoOicBUljt8TeoyaaIjUq5uZ9+z60lGNP
2RwqUdp+hzeV+RY01uAZ2jFpPAIJWGs0hL0ga82CZkL84H4dp51UFAnL/+n45JKN
P4BPBI6oNGsPH6hjHmk4R3lvs7BUCSqCNwCXVBz31MPi4HOHpotMSb10ZFk/OlLB
+yWrHuKIamY0ytqTDQvJ5FQrni1PaVSu3Zr6PQecP1gGnYMkRQGZpnTeUdPxr46p
G4coIzPzmzrDcJQ9aevmxmu/WerG5n1c2GaGG2JuK9Bj4DNPsn84HAnXp8Lw6d89
ycbp7P9Teoac2gMT5ZidiMq3JxsZ/2YaQv+QwhMUzLEPHugHF5OhIBfW5o2LEPQ1
undaEMUL9kEps+OZvqjWVm9GkaQ244rGKxypQroCH7ootdf2s3VPJPI91COkJZgw
svffBQrwkC2aKko5RlzP8at11qtLDu21pf2adH2kWAGuF9RzBHcLbpG20Uvaj9Lj
qe+dygYlQ4v2qJLysxlqz7m1LcS4icnfDRlC6SLVSTI4QexoqCXYKxukrmRZIJSx
aTLXbciig3doFrq+opciGuMnNeLJmN9WoL95PGzalWeGodFv0Tg2V1liHBjIJuSS
pkqWTVz8cvyrieiF3aEp+7KGTurI4cySICDLLjKwYbZ+8ak3vIyMlsSa/eliAY1a
U6UXFka1zIf3b406v7gdhI29vsT2qkNbKJi4dDMa6+8gasRvcz/XUe9UH2olDg+W
pv0fYJtla+kmgpnLuBsAQyZlA1oqGmpLSHpQVndZPvBNes2T2zKmQ4K9QIAGh6QT
+cbIOKJ9uXt9W9wS05PgsK098LiSAF4cPjw8coKt2HDIXoR08MPk31kFHSXgFdDU
SKv1eeXVeJAnPRP8DNOd2MLCq+brTUghBZrIDJ/ZiwJHNk901CAlqHGQHc+Ci9ga
CWwGfUIzy8ZQwVonwKaH7Uj+WfLWT6QBprLgb6n3bHwF5+4T1+gEQlwcjYhC2PSK
rZCt2XUH9+UI84B2t1Yx1DklA7oDApr61Xb93f3YMcK6SecCSWH9wOit4j4DKRhb
w295HQlDKBAxlfumascS0ZDpr1agIOEz8JyXuSlBWwjRpPiekwUA4e8rGbqbv5h6
kMjAuBM8AqI0QoCrls+Ozz1zs81gs1uUOU4kPHjjishbDy5t1/yjmtl5/wEsu5Wa
9lRFU45WdSadcUu1G0v/CPV9djKlbI2b6H0xGhIWtPwfjUrtwwl24yTZYwCULffW
JJrenQ0wH6556RuYYxJAgRxbYOjMkpJcm9Yhg77JM0UVCFA5nHYM7g3jj/+ogFhO
ykcwtSOKTmQo48dJdlCDrlmr2Lo/LIYRQlB5J5X70rpn7AFqO2SUZieJUKSv8DN3
NrRUx91jabGOqAxZd1v8NgaKQalSqDUoV578Rvfab/GwXV9pvAlNXk7NfJvoe0me
8ND6FvYQGgKqcapqte5zWRuq/uZMp6zw9dW+4IwMv7vvKETcXCRYymMpgJGXrm+j
rTv+a+uIW45sN3h4ifv8AINGYnizs7DHmnnmcFlS0yLtjXNr9cwCZ+TO9GumNgMU
jsAHC4iPhm3cYDABPCGv6pweb5KOu/uiJv+zRdOO6COMrXcwGXlB05r5g7jViOq/
aEd9jg1Msrq5rMDtSwpZUbDfwioXDZ2/UnFVIbHxT6YomKOFmra7PLwINlDTkRa1
brzcoxnIB8s07MY+rxNmeZumayjwkbfjNuFLEGZZORYKvwIerVzqJmtsht9WGRdG
7TfaDubNFiOrIjTqLWlNrrjNrAztc/MoWJUhDUXKyOAIGWLQfSZeOVVBzIgN9Fuc
POFCFmMuyU9mtLCmNt+ByN4i2abKBxQj0sJEgTgQRg2+JphDRHYFKBjhPnscoTeh
jcIWKFzvaf51yvG1wUeBv63jP1JnNt2A3PcMRWDMBJ9ZGt7HPZ2iAF/6uovveLPn
a/EQa9j4IKlurFvRZFWlHkDCawlRNCor6GW+wdwtkOpfpihKNTt2A6RgTT2mp20L
o74wpnAh8T97TpI1K1wSyfpSiUW3O8uduPlIevjOfDWpb901KJ9NiAK2pO1V1nEj
Bi6AeD+QcSMiXc+CUBj6YRSQ1xnEn52EOM8GsxNmgwfshm9sSx8mw1NZs7FSyzD/
PpluUoTrcVlgwR7jRAsQwT69w5eKYQgCHmX9ei5/6Fb6sJsu0Al4F7AcloiZu0z5
kzyItz8o/k36n7bibuGYEd0UaY4XHraRRnbTfBOAEmPlv78ZJ3ORTPKh/Sjb1OE4
4cRTMbITlJC/Cpr/uvh+YYx5hwBFfNYMHyAoUez9+Un8yxIFA6xSopGG7aVRfa8F
J+kCZiTzk/QuHLj1/CS5T8KgHvlw0JNy05ybW6pGH0+dbrVbIjkrTen55xXgqsBt
jM/zbR9RMZobbS8M4QQcudYRjkQ2dyMI9B9D8AOa9IPyAz047rAA4l4nRNTn4qDA
zFjWxizA7ojWfuCndWoKzmnkd7S5PNoaxiiTHHzUPkZAZjNKq0ylCOLqa/N40HSh
+rP5H0J+AJ3vyKgoDZbf9Jbbp3h+iG8rqhIIkGzsSs4ziW55tu2EM2grYgB45p2o
dK08fg8XfW1nhUck1YwqlAdNfjyyj77tVpdNnG4t7iyClX5uf6L+N59iauEug56v
lTIRrVCs+zun9dsSmnzC/dSSi2EYdblT0TJHsx8j9ps4wmYtmV2t8I+QS8k0oFiM
UzIhEtNMl2yBBAOxp0qY/MzUi1YmlidHDCLml8YkTNOM/zJVrzjjeNvMdwTR72IA
kXV3PT2dwiBpb3p0LEP0SyJbw+zx9McLx+gjOnAx2Z3ekBgn3wfz+qCRuVygzwTV
rfnNkgSRU8QH7zfmb1AWTW7Lcru3uPM6zlKA3bBQf7eKIUGR0s7f8NbM2Yx5oRoj
pyZC+bS3ykbVyNG9jHHaYNo2t84CUZMoDnNQV6G+jCOF7YhhEHObRB++toWwKAbb
n4RU6lwDrcTVp1Wecy9FejELOJrb4445m8TsBM1ywn8nwpSTMa5pS1p//o3QD8Vw
5wbnj2qJ3vVyEvt5UYN/Fqk5TK2UIJdy74FVJpWkOPyldnOSzPqDyQ3ufxnuyA83
A0s8PD3dHmxPeiV2VK7igmKo1gfjjcEHDmDWRlWVsIgsbVeQnSkTXAuhtjhaz4mr
7+CnmMMyyYA4XsybP5V4k0kpSTrSuv2s/4+yGn+7PnsWJa5+50I/qJdfostuDraa
9zrB3Pg8Oe6DZpkSh4gJSF/9Jq/fRcQupGNotFRVA6cSOxvwge5AL4sVaAKKHh8w
kzkpdzVu+5TodDB4CmZ+sRNWLjB5ELWaMfIbGcSEY2/c/2V12AC2deNjWbvlWfPO
IWbfd68OAKXpwfVpZXyPMKtZvrFGwsenWnPzcDau9eQcd2pwkvMBHGWJjV+WJWQJ
MdYYueBOyqeJ2Ip0EKwRvxiUZIwdEDCCFDg541V20ErDVY6ZFG0R6PL0wQLWnj22
YzeqMb5H1vnXuZlKrFAOa7uSqOdSOwVdtjmMrg/P+Kd9VNAuH3LgUN4D1kwlfNcx
J7YG7BDnHAWtCboF9wXOebawtT3+uIY81ABXs+HMnjq4MKaTiPiTK1/nuGkgJfKH
96oyu/8TTfDiG2ERcklsZnMa7/WX9qeSoYkuEQ3YdqTlYo3QCTskwEssCzm1as/Y
nmiacbsUsiF/WNi2iounSHapwpvfYoRCrpy9hx7g5V+XdZMaPAe5ZAxDJHB42rvH
Xq5t++0T5sTw9Pxs4tX07ICuea/yu+/UTPGuBFT4xsUGIvqG0dOu1cWqxNu6pPDn
V+wlRqIjWoWjZ+H1GZRvGmDl29Y3ICn9k1pVaN+QRWDPO04b6Gcnj4WSr3sVvDRX
aVCiGwtGgioQI+HGh0KdX+Ljtq+flqZ43bgKnbb1tyedO+74rBRJzDkEmy4sQYWv
4Hui3Gu0P5xmJ+3fNbXHyJcpqX0pOsWst5nBasmp13NoQ9vBinkn2TAditaOYon9
HelbV56LbR/A0kOhfLXjCtGemx/jH/mwERH9xIZss+JX8EfKnd6WCTQ03y5vnm+r
PKPhCyz+7nnySLPlacFHQqNGRig8f0YLFnOHsgtmTqnFryD3p+Sg3jNDAWm8fNsI
OWeeXSIkUqTtrBfmY1EAurpQZImS8jW07GKibq4rygKEBrFMU/DxYFxbvCNxQFSL
owOhlLr5BwuxTjWkI5EQpoIzn0kTpWZhMKgdY8e2kb4q49fc4q/zIeXPFEP6qZ6N
IVPwg38IudJhVdf05mDra+cKRPaECtYVEyTrEk6CiCWuqAQ1CzC4mNJw4Fw+p5xb
uRzQpLZN35R4MxFwmlqKykjDFqotaDte3dIWNwxDbZ3O/71tORAqN9Dn5/rUUcyo
wswEg8NvlsnXj37QWjpo00mLFTKF8TI8WJ1u7QxH2ssuEzQWjqC0c3zFOlH6Ym5N
oTOWzwssK71QssqdJUBWm58tkfsIMkR7g3wKoCRF5mn3ARbFHY6GvjFKIGwruMd/
bdlJRV6xHhGxHUFfhgosVdrvju0aMhUsgiPjHccS/HL37oQTDMAnzOM73cy3CtAC
M+Vt59ZKeRQUtbdMAJ/8xpP7ziwYgDzvDlXQk4HW6kw8z5hv/Q8UUfY4Ra8rcPfB
iW6EtBATzEA41DvlIl73G2GmXlrZcbZZA/wQy2UHUE85ETf5FdvvwMTo5c/CYP6q
Dvmv8GNkSdSc0X7LYmuq5xzeudwc3Ekn0kEcjJfJwJv3sEykUscCWohSjQBVZHzw
5T2FuoFZM1bUrClQ5BMnrPDXWHK4qruYm0bU8BJwR3YqLILjuMOXlEC/rq72grTz
jDjBwqqJ40t1m9hRwR93P0Qw8Fn7WS0IBQjjFxWEfNij9rKwBb29guxY2Tz2DEk/
AUYFLrhobhJOXrjjybr6qxXIDNyRuniVVMlW2epbyBKluzvtkSQJoQuim62iUL51
/dA0GMvzVrwjs0MLhhQG/BCPqs3TsWBsRJ5MdkZg3r0ysxwYaB6n35WqjmfHVCc0
K7HKgqe4wWwy0SxDMsxWHOtPSl1XTqt6pj39KWBd9UB4wbPHIiC7Jpn1+5BJig4R
cVqD580mZ9j+TGOVMMoB150mGMn4T39gLYbrgC6WlNJ0VArYZBJQcWvBqCxkgxGa
3n/wUmLj8yJnG7VkGCVsQlits32J5LmEij2orn8nEjz1P5cVlUkpYULlSIP2UJxF
kMSdF1FU06gr077vfIOx3Xa2lASP3pCzi4FOXcCTfny4a8Pix1pKL577ETaYe0h7
H502HaFBRIzIMsdubF/DFMSsbEKZYdcYh1LmyUYmmHKTMffEQ+lRlrDwfn3/k9s0
O7d3ADyZfVeDDl8q9ypl3PyHTL6KFRbQpEVow+q+2inL0Q5zj7foAR+QEr8mxTJk
HOB1OVBv4vc3D9l16SpEh1b1hyqFK2sk+KemnfC59P5ZnZ3JWoyjp+8iC/ZKWg6o
dxLlj057VO7aI53L7iBejncNVsXvjSrV1sqaRMJthDVFTrAe+1TIUltDNiyrfVwb
2LWHIB0WhdR3lgjecbLe1LE970nWdu8oY5drjPXoI4e8Z5JhZyU2Cp9YyEokW3lp
DDUQ4o4C0xSsyo0nXd0cDtaa5Mfar2MJzAbIRA0ZMkllq0baAgUrHJxYahpsPAmo
DfZsjgRRFOHeJXzBIC+yYV6R/+GBPt7lcdxj2PWUso57N69myHOnUKrHvQ3/wAm0
81LTl9K3iKRGEEMXnh/SXWl9QFyc10GT95uyluY1yEkzpzylJWrn+JFtSYvEAvA4
xDNpoCsSoPeVc4bM1sXMrQ5EwFKsNct+JE96N72gsNmJKNcO4MJLCgrlhyi5wqX0
2dxBn++AG2g8FirqZizFRAGORyth2fC6CENzlPpWCUW3cLSbT0tY8mWTFHHu8n11
hUGQLqN9F/ciyzu+m2Qz2sAVuThXj55Ge1R9AFC/DvB3q6WD8goOnoGxphrgQOni
KSeQRIHybpQxCUfNm4YwuMUNdWev6vuINokM3GzqlS5flm7Wcla6TMHwE0CiN39S
ESUlefbXKoi6QOefeJvJHN4Sk+JHuxbnDOVENdeMXphhpkUYHofZts53zqaIMOQT
SAAXFLJlhEyiqbDEBrG1h1fGWIhkoR7rUwGADktuiJDGdnyeSLQ+yfMKltu2A8Ui
XtvOiA1yikwwSu5dp/4cHmTu5/Y5eLKXzdmmn1VFoj0H1wc3CuMyiam7mpWQAjMo
kvLYCKPz54nYyu4hL3U/kU9riAP2+vZ/7if7eJE0mot7S0uGAsLPyqXKpA4Yz56h
vUo1Ptzr1tffIQwCpaqd1K61cOQVD70fPvnt7rirE4YSCU8CnXk8hJB0EXwzBfUK
krmhHPmHPx0E1bMxNpk4D+nx7+7DRUulhRIgil9IdL1mk3fiYAFvZjQb6Cfcssgj
cohElPhD0Kjvy0qey/oN7CKp2Ittq+4KTnPxFf8jSMl06mD9bp8JLTOHUvdrI4pu
XZ2lbzCx+OUE7br/eIZsXYHjMCwXT9TcYKx6jILsQuYBoBXNhNBfR2/qk4430aF2
E2zy0m3xTAjagsonCKHi0fjuQEW9+jQobcSxJKNBRmVEsZNshDZn4BJ3xaJrp+vM
1G9fGC6MGgv8DVWTYhlLIh7RMoFUz2weQbSxO0smA4V3SvHETMuP+8E8pSqEzHTl
AWO9Zhl805ArIRxntGBR9/hI9+6jpa9OF+hO1nwhR9RnJLb2jCaa0+i91I5fmzJe
BxAPhMX/QrmAj9OOmU5Acl0GIOnMvEVR6kVcmh2tGFteaHPOzr0sdxmxHEHkHVz1
zhWTnPouCn4cbt8htI8sL3Rol0r+SOZwvwu0AHqtjKSu39ECbrmHgHV3lwMZCUo6
j7lQKJoLTa5kSprTXnt3IVQZ4DWvit4B8+3eRKdHswWy4uOu4QKQP9SUBwLdEMeW
tyLlIJHvaOR1r9L+uB10Xo8pCX0Wah09iSvP2dJdgCfegDS8eZP5sxGThOqkCG8z
Q4CANAmb6A6z/Sjo1tXgtJ61ch6ObEzsQC7+cJbS21pfeMpGAxht4STaGD39hSio
10u2ZMiSD7nyfZAqtg960YZitD/5v+/zz3TBks+7oWqj8eOQN1jevYfgNS+8Iqwb
Fuz4Z2tTVGor51GIYbHDQS1BZcBsRUZdsmE3SUuIAgFY1/IbQM6PCqA3+82agXLw
yXTz/l6PyVm2EnH11sjwXX+Fnaa+ix6z0tJ0Aayo0ji9782b1f0biikcRG0YyKxI
CKpGlxDFgolOvI4hX5gcE1npZPmZHHCQSsqm0WjiHQUqa/L8vpXe31Fqpggs28MQ
WO1/EJoPoMTva+oYLI0JHKq/HlX9wDCsKGdoeQcnnVCv4ffPeMdgSLyK/takHttT
by0y2hTxS7KokBxBYWRat6pJbu1Y218ANoIG91lQIcgprADnBLKNbeLtqB5g/DlU
R4a99ARXF4XZXfUp5hhvrsLh2tNkRSKZNYEW6kbW7D64Lqiq8zpjNLJT0A0I1jj/
VD7l2ktL3UkHg5CbGilDUjR63CuFEE3LKyFuXxEiDBDLq+nzZKVYYbPK/Da9XXhO
KeJCys4zqk5B7Qe63Qj5FGXP0m3YSJN/mTXHReRdyry83ybsE58WLRTYHNAfpf1G
nhZ83XpkXsRDIiHzNaQYG4EaaoANul0ec5vL1Goe2QXu3oVotQJC0OqGrMz2yDDi
WApZRVIiB7yXxMtH6KOyoEoBR77ZB5VDZDXMt/QbpC2J+LryMI2RjW0blJPC86Dx
FGRVb7eiZPA6iVGGHZXORlUuFP+lU1AyIudjVedlt8NR1AydEcuiis70LUbU73Ee
bi06x9TlCHR5v6krFWvkwux90o3Q20bW/1sN07zugvpfiPMtIFWGAPp0vf8h3vK1
aRof6NG5etmjYDYlTFLGG0aN9JnFdSPP1go3zYDsXg29/IrKOi393yo4NF1xkuNt
qfLUvSfOqHZY8yuh/RfK73sySdL+Ie07mu/i55zCkVN5WtmO8Foff12BSCK4i+sU
+ArjVCvKCJddial9WGHNYHPSOTXZGuc+P8WFyZADrglXY7I4s8l6ODPmB7VAcPDP
E+dTBltjDL+QFEEK8yIUNO3YcnK7958Bz+zfhJHtkQmc6vXX9wWSUEmryIvFwqTZ
oN9+bunK0Akt7wqCvx74eyYVPYzNxk1Aegd8LUpzzLRkKVGm5mtk1p64bAKA5aTA
wDLUMF+nA16EUI2Xv2y4fr9jZx6QQNRmX5IF+6D1WF1CSa2rmYwyK9v+/BnENLTO
wAx7HaGPilLczV5t8EbZDxeG86XrtuzpCP/qc1MwfhQjeL7XLTHAuvpuCHzSN+q1
UrTwkWdulvFeiguY2Kijqo32O7pKcYe7YYq8TIDcwpc8Q6kSwVy7T6OJr97qCltm
83F295YAgwi8WKYCQfmnkvfwAYzhBuaXKAXtuQey/rTxenkQVCauutd+FAQ5vUhr
fDpciJkMpm3IOyOPhiKomiUU5KKOWbnuVmIkWmiM4unxu2DJkjbcVfjqAf3H/eMK
iWIiUomE6uyOCQ+Jv9Gh0s+NavLWA2zdH+rpSiDH8b/OV5vS36aZ4+5nH/zFta0N
18PgIDFxw/W6SaS+bONhUWBhBIVVRzzbCgLR6pOBtqZl1A/3+4YFotL4hLyq2ajj
QhlhEgCU5t3AlQ2dSOczUH1JumM3xYLbO6BJpJrUT/xr3Jb2pmnj9b+/LY7OUgJH
O1d53EF4gyy/S5YFLmCBoKEZFr32VEaDyQ8Mn998ceMh/H9zyMYUqT/pM/6u+aUq
Ai+q4Z01oBlV4rOPpAU8bZhWBPO5/qi1avtWX3mFI5uizLKqU63ze2Zxdm6H4ysf
bABzvJikcWkLZm03fRkJgFNbDhVBwAPTan0P70Vm59mDH4di7ZysuUJPwFBJK/6f
71rzBg5kSsAQZyenoffL+LYVYYVsm4rY8K8QwUrAchh8A08aHZDKM3ytmIWINQAB
XLz3WCla2PKWhx15j2BllCIPEMGu561lTWJs31YKV5qqhZYEwANFeRVDJa7tG7nh
/hCXnFQEBkpyKxXHMFKVVuYVawdA7muRWbBaTznKABh+aLuZ0JiQMi9t4o9p/P5H
S9nrVE3u79Op1f1YFlcgfqISiyCMj1LjaxTYZq3KujgwPDLGz1A4+Lz8KwMQVWjz
mMd8wD5IoB7F8vAL68FjXhhC67ZCWGkfLFVwclUg16hQOCskhZ12uh0P+67WIZ+S
UsMGHiXDzjblqYMS2ptk3/s89XFyCtlPtiTwMaVJjP+rRdSTj2z2sq079uWStmOh
UeMIlB40GQ1RPeCBr4/o0jtjyAh/LDL53FOTp4PT/7O/fJdQPmJacatrLvgIgliR
dvfkZ0o83+QoRL4w6BplNF+k97MODvkGKwpAnRu0Bu4b3OkH9caKeFTqL6Y+mcL0
GF0m4F3/RedK+YFQZr4jK/OqFecnJITBAeOwG4H3RgTh6WRQZjYT7WYJ4MRgC7Gh
JrjMmPgNbBjgPfrDsvmNy7H+3doNON3xPxtfNQgl8GhEWzSyXwrOYwYFkXJHggXa
PlvJzgDnR3gFH+5lhWTqQ/vVzin5kX5YqgYYo3MExvMKuW6J0Ru46qHP0WXNphIJ
MimHVlEIhOhoNlDcmHlheFwnsxyG5MQfyhrpL/mejRojvRIRN6Fg7sVb+FLPCuSV
nXkX9AXTGXxevZDBI7UOcrV6wXs8UEm7v7kx780+QODISN0DHntmU6LBhtvKi9SC
sCGKpCB3HnQqroQ803qu2hKWmUDU9oncwMmkaNxV5g6sPBAJQH3aei16oh5jzmrF
2AMdKC2qHv43EtgouDyIpiMgZgPrcgO+vpBZSpwN4Q6P67zcK8HsSX8v+8/qEUTH
9po3fFqdGycSOzq1XHh30DGMAl/NXYVTxAliqF/TYWfo32TJl9J6Zwh7Kie4UdTF
I6uSbJOw0EIcJhEtqK7x8HeUAXwPdGK2bpzWdbnsdVuY2ICs5ZZwJnvJ2E5cZ9Zk
HhXaZUJpkzVH+cvBTUWyLHXSEK/QfzKZ84u4zeuAglz8LpdazNKnlrYnx3RiWXVO
rqW/9n1/2BZE/AdV82nqHbZ6tByATZgyY+M5CbAyBcmvWyD7ZvUFgeGtmuzFb7zL
r07RlhAjb+yB8E0bYy/mtnD5y9ketYLF5+XtigrcGuuGIHYaN4EhRhPKzYf1/Q5V
IlTQP7Ou/XFkTn8I2Ln0ca0vy1FCQ8x0L8msBvQRH6tFssoKeHKxDKr8l5m2BI03
nr72tKzI3MsUSF5T4aU5uPdnuzu4OOmE2Fegj5vFzkK63vWWR2fDTli0ERHhsI0h
Vq3o3Rm74h7ZAoCimMI+oyDrnQW2aPWbnOro0Q6HyVmVPVJFGelZacPnQHSpBpyc
8g0QkljLUfUSY1yBpxOtnzUUVN23+fhaCCM2Hs9TQHLkzd+2oW0FXedcsYjRqz/N
WdwM8j6A8vFOJUm6M2qmoLHIeSP4Do6LWgOZ9Q21Zl12oYi4MaOiN4/2RWNvF/im
BK0x85/Wb3vMxyp1R0kNDrl09ubrT6wVdDnOtO/tnbWXAyUr4ZkWdANsgtPCTjo5
/6NNDYtfX/9rg2lHLvPPHrBpo0ufJVv41oepzwrD4ivU/AO/7DHJcNaXELTAtHBK
rrsdVPNR0ug/HCK5ZEe9/Iqa2gOHoeKNx7ppOdFbDAAmxvBWBu4jnV4DaJ/xxJMH
5C6emLZHvD4tlo5Y6KaTQ3l6UUSyIdvssy6h/gBkIviOb5oaIQPlp2m73Zpbpx+7
d99d/DnHRfz+XemBH02InOIxZk9BtkBJjn7xCzsVZCeZ7wUo9X4j3JKtWEUhD/CR
U/46VF2Hs+J3ljGLSrYTPTBCEt0kRhCdi/TVGVou7QD9R+gmMOCCwGDql1djlCVj
+fByXS3FM7dw0iHH5T7Lh7mXD5kD7FCVGlWq8jJzbeHxfuAjnhK/OcRhSEn3Vwdq
Fy+rMpuTfIFEtCoxROjCLA5qEz8iKZTpkgC3jPQq310mZi0KnyCqc524LOxpx46N
hGVGsvVsHCFNoHST7J5lka5Diuna9WNDZJZ5tjZOtPgZ7pIDlFGEhraFX9+I81lF
Luj99+VJHz4HtkzsX2J4Ocna5JLmDa3I7Zo0Peu++8arPqwzoEJV/ngEI9h9Jeqz
oMX/pvx7pWjTRt+BuYD11Rh6GqjAfGkxt4DoDWJxeKUH/i3eM5KgwlSnHwhSTRgv
6FZVEYBRKQcEQhg1F/HpRYHSPPY8X37IhCbWRYRLreY9jt1GzQBW6rLWWXSdG7mu
TgKhCxsskm7ko0tvDlJ21qJCvlMYTIxdFG6pxY5YMLF9pSKjzTbDtLqW3LSg9EpC
cDiY8mjQKYAu8rX2bBCEcvMMqJZvZSy9+tSg7jj78RioXnp4GLuQtmVoh4F8oMDT
bYXH1pTcfAq0+dZx4IUGsxK5jJVMpq3It/r79Idu/CMZxPQsk+4G2JGVyZxs4rXi
2oygd4rf3zN9Vyw75y21HB4FvWqcDEVcsdzOLaWN5hl6NPtlX/OW5sHsfo7YqEhW
k96hATHi4gZB39WgVx1kmNnEfVFPVaIJILN4i9DSMFwJOl0DXvn1M/UkEIdFyjk/
QN1Ehi3+Qdc8GOI5o2dy1nOJ17V5HFAZOLpSd0NIU/s371NVVzliipTpdcL+i8Qa
OBqFrly31BAC/4SvKmtQkaC0JJd48RPNm7fFvqBGAq3ulPvGJ873PBE7jJ4PSqub
kyIy+rEYwFkkt0u55qc2H/WDTuHF2J6VWKvbbSPKocMp0LGCoIh4ZgDdRNQM8C4r
OAXyZQyE9xEG0sUndxs8M3bqEMlARw0IxM5bvO9Cf1oX0BOhoHdohrO7WaGtyyqM
WrO8DiH7uK4Fj0JMXPql2v6iOJtzQacHb36hHQAzH1uL1dIuDKb7P43Zxgg4CT48
guIjNeye1Eh8m2Z847JJrGOMQ9156dXR4C/KARKuvL6RC2Zsqg7A4NorgDqWLr1t
mls5jIbHVyBrn4YILfTh9knZIjgjhDarIz2Iv6QOX8kpXJ7pjGBi7HFsAiPDZug1
+SOV9V3ZfCSyY/4x5dcGnXPkMGBlcvyB9njSwn8ervFzr6m7pqhhuYufXI2zkydk
mFXAb40eVO7jgP4L0eanNOLhb6w/zDvyMABWyhW5jhYN35pJNaSo36CHmDLNXMmo
ucuaW2CfSoCwTQVEJPuXJmpQWFyUpWWL89g3Jj7YTyyHpwg9KAcXSxqdhM3ddB+7
3MsLfjQvmY8H0pRsHofENl4ZAyeEi5m8IBdXIdULZemY0reNqmZFfpHl0NHuuRlu
2AeMlZ02vsftYnhPKWi2P2+21+pSoX5IPyiioAe5EQBFpDOr3I/nrF44LwR+/yhC
6YEhhJeWNcUpeE9yhsTJSaRQMYqYP/f6BayHo8wjEdCaaFZqItFVSK8eoNdNzn48
lkqFP4N6jh1m8hQzoYli3EcB23bQ+R+ha5IxVzMgiwvd63r+VFpMZpBehEd1kDA9
7wZRNfrKj1BLkq1Q2J43QVsnz6rNyQRxutwso8LyeRUWGe2w14Cw3XixXq8CeLCm
eHA7Z39pLN9Igw6RNIMMvJClwec4VXkZ1YA5I+E2UPq7ExP+pMe+vMq2XovEM+Ne
dtcHyAX/sqzMU8ZJLiF3Te5QDBu69lgwb/AO7oRTfBmmRIG7bRpncX0cD9DW4DRU
P1I2bX8azoXFfqwGa3vCIllvX3GbDOPj4lpQ+Gh79435bROaiX0d+BOXLUjY5Rp6
4GpZp0ZJRbPbxteMnNTuU9BdzNWtlRVN9HTIb8I+aHtulrx4327pfmQfnCZrnhIi
+lxotdXLA8n45LzqZfyx/WC0PgULR5hrkiX31sDomJeFU/My0UTCtj9IN0HLYxHZ
zgMkDssDlFGbaZ7G6AYfwZXiQxdVSB2+Qs5M4pPs/KgGqKLCuSQSBT7SsHJEatkV
W9FRU65xdts1ErPqYgOV/1W3D3art44m+uK3S5h4qW4vO7H1zKJS6r8RJGD/VjAb
jnyauT2BoAaaZaC4C1x5TCYzTMKPQWHaTwY9jhCsJVbYn5U+tkaNtuiz51x42AnT
f5ncqNFBziCLaeZQqLA7tD1VjrbNiZTYLju2cSuH9w05yQkWHv59KCJyvP4AUj94
d9lFbxuzB46VuCGNAYCbMss16QfiubHII0EINhljn7b8WDrLVLZAL2IDBZa5kRTK
/jD1gfq8Yn0qzPPh0b5A/GplbL4+jTANUggLRa1k6EvZJxwBdUaRG3tMrjNsgDLU
Nj1hpEEnUBsx2OgUacf/suIFBRT96hLpMykYnSep+3+L5FV2ia25U3mBLyJVVLM6
bcYgKGTGItTD+0zr4dr10D0x8Us9LoVUfYB2rKolVNAUsT5t+fY74BqFd4JAVWIl
DjagoxxLEOwJiFwyMRrIKqXkQqMg37hy+2ibcoMfSb2rY6QpP1IcJE7LGX+RHvq5
bg/pOCNLrHkr51IIX8ePSlE8q2h0M1Qo3f7cUijG4497u0zPdcj6GIMHkX66526O
H4EUc0YAJhZVVqGGI5uXnJKQRawq2d1OTAkNxnezWxUsyx/tchtbEmSzsu9hDN2Q
l1SrRANah1WRS4UZQF4FOi6aNYHLaNMe8CldNcsyFLZC3g7sw6eKy1MB0G7HDBvB
++egGQUKvBbA+j5qtH2r5WlCXmUqRNjgEii7M6xNHIltIeWxz5R3ynnPMXD1W5cd
C/TPY9ZyD3jTyFyNiUiIQZw7OorSgWA3R4bOKbCLaDSOPEqVTSPCHpi25Nw+pA/N
Zl/fKrkJVTGzcey3OfvrIiu0oNljHZCiU08Ok5PZvGRZEBJwfcAD4qMEoreBXer/
cVH/iE5Hqi5myNkgrJ6V7n5Hw4p5rGMxmMboFt1nHF7RiYWC1o/RmIAFTxmpYIzN
6yKn/lOXMPUYvexKKTYbsEj2cjCDis6lEQTZtjiVd0Eehlw+DrDEl1hyagCel5AK
DNGR8xWvWy3FVveR/8FKniJbTZccpHw4Kc29fHjCbd2bjy15iaVmAESNtUcWwSlc
n9t0lYt68JjkNcUlvIb2fISJQTJxX3809fwdzqk4iRfkmX6FQYIH45OMwW+2gF68
sOFM/uHj8ydqIauyTm5vUglilZFH1iTv56xvTkhKwgWBFwDqHcW8XCROqGW0uWhl
riRuQQkybTNnvLRBGrGZCLoNg0YaywvEY+2L6UkkF2G4mZObqqSURKexippVO3c9
tvGzBdamHoYC4m9ZoUZ6Lv9yjUMjnDmA7wjYWvN9uMRsbqHiRM7zkaM2VlwsKdCN
5yfnmEhQlmHYi2/T3XfNVqJXBfyEFb6n3NK5rX819J0Is/aPfwlswnLLM2nYoMqe
fBi/lBug7VaUxls+Rh37ah27vfMlg+uO2Bay3Nz2Rz5uXJv7rjgeAT0zXessk925
tKS7vE8NtpGPtGLGWLyuZS/xHZEWr/Yfp/GMkmaLA3sfXBbdqtoKTRK4RwrX+Rk6
erPGUVbd+/1nGkqDsyRyjaEkAKrewhPxz58IMY37cSrQzjxRlL9p9Uzfr4j4kHg6
ehduAvwo4ZCkI7eH6mnZR3ri2cJ+Tjr0i7qtIbvCxT56pMPRFX80gsljIkJKaOP4
k9246g7W+6N7Gs0P+xk8920nepfpWxKXvD9/53mN9zMxd5tm8DxOiFRXj2jmUjRn
fyDNuWDxyu2mpYHdELocrW66RN7latUrs3kUkO9nIlBG3OQxO983+s9610xw6t1e
0beIVDxs3J12IyBjFLtpFbKQQ1LTn+ikAEKCzvl+o6qSNTo7FKynJSmSclHZ4uLK
nLWutDMGDtQ0JUTPdSQaXhXNyTe5nf1VLJk/H09VSTiKo0K0QfBmK8J+rLdKeJl3
sxWEATrIHRgjNKOqMZAyPqF74wISPOYZ6+xHnHB9VNTYFdXeRL94PXDXXRsgk9qa
MMUI9SYDLvGYvuXU56CRkIb/31xHLQd5aESsiZLPUH/Pdn+/p80HpFOLL6MaUDyy
UIy+YVERu1JU3QNN2RsI0IRw2eq8gRpIeKCGebL1FmENUTd3E1Bz5f9KFwdgGsaM
BN21XYSvAYQQPtNrz1H+lYDQ1eVu8cwiZRcMyhYbB6XzTC8VZQi+IqccjaOGDdBy
mLziTIXns4S5+d0UXNg3D86hwOXcObvKFvLAa8a8O3iT1Q+JtT42w/GkFy6PJDJe
phCCC8ne4tvXcooDB1Qqfra0AGGEkxJJW95ft21YeicB8E0sr+0UIj4th0FoB+uR
hq7RmtZJBVuPlnQfSG02Ry9ANE6GkP3zSS99F3LXog+w+1Ry6zaAJYVR0OJibXHV
4vYvx6H785rq4W5AGOWTmeFJKhAzKiVpPqzXLfTBMnK/qSiDHy0NFiVFyLn0nP64
ok5ttwYubN4Jt/gkKmtq9Elbl/U/hS15u4X7srIcwire86Z/tzilofGm45xOzKo5
ixW9ydziCYHQ7/3WHpLJg0l5VCUXjwFF67F7ORzqXMQPtrRx5mYjAkSU8gbVSHly
P96C7CgvLWQEaghtr2DxmmpJvKIn/rZGS+0Ng7rGW9CiQANrAHwSS5mEUP4aGChv
SQC/5IxRzLxMY8nqMxTAO00zxBTaTmB5y555iLp7prQTwId6j9SM9ldVZLxchxmu
JSWe2LeOHlDddrjOCS9wp1yFXIUt+toDeYb8cpjaWx+Z8CYICZWTjknmBFbO8S2R
zo2Vn5WrBFMaPTIQsYg6Y+Vt3EqRfTpM2PZCZYWf1L1FWkwsAhQhtCwYfxW+O30E
qOYaCbdIRJpKayKdu3XbOcSDHmmOoyJoMl21+zqe2prwIxpC7eNnBJRu+wR52dxp
whGWVpGjTOVzjOBaM7yzALP9ddRb5HVrQhla4DRcq2DINazcRdw+1MF23DIC5DMz
YESoJFSeASnosyjkKUHKqr2qNCu8Fy1Mn4G5aEloNCUSOQ+SEcs9ALlpbF0A1Emk
Dz1waENbAes1GmsoOMCGvlZQewDUI3qTU67ikMWIocsXSa9QYM8dhX/xtAhegogN
fsU0mJYOxPs30VkYAee7mLalb5lOG8l/PsK7LEQlGz3JWH98wPlzWiSCUFFIqn4C
OV5i442zRQSGG0JDr2IgCXAi6WHpLnms4Vg2JCA4rLBoAk+crgRhtThTKe9Mlkky
PV4khBkPHY8qBs6mkPvbupelW7nQ8a+/2cCoNS0VycJ0TGXL/9mhMzQ2AHeQqvAc
CJt0OJFKBuOzOg/KhM7S8ia3rJndiVjo9jTUVqXUb7oOlO9wxBe0/T9XDUmotl5w
YekP6K4Xt0/k69oU0sJ3Ddup6RC6nL2CyAqsmdSzGmL+9WV0wAj8cVbiPdm6iXyx
xIapCbK7RjdOoOOQwlq6b9AteBkQGbjMjGMd2FO3mrsGLBa6//20dspgz78qbvWC
6WzCELqoGaikiMTMHOfCxWA+TtedWb75t70FR6oyAhXM+deyRcHx69MSxpLRt2AJ
fsGH6wJbfjtvg8VAspzdwD2/KDzCOCNCf6Sh8kVjzYtXKn/iaQvvt+AZBg6jinLi
FclTfJGILzld4o+x/xYSnnJa4xaE0nifnfy0bsnuBxcIWUOyMBQ5QldDlNEztr7J
bD0D7YSFujWdVdqRqzF+M5LafTXv6bMc0A1QEOGSj/QAWCMp6rUPzygEe+iDTunR
eW6R1nEMitY2kGVOckjap70LLC2cSLDHzS2fITIHjDO1mbc9pxrUEq9uykwM/dmX
w+Uva03bfuAlYl77+eotqgq/+yPQOfx9nf2GooLUwsVw4/ccu0/JkaMo2V9FXEIz
sd+fvqvKmF2SlMbjVLL7oZZnAUPa/yqNV1LiW6Jd84m6+u8ZkyTKwcAqVERmYsJy
s8CreMYaIGiVIdJ13AA04hw6p1/YoAlybCP+6CclaM6piS//3NtQ6ForTVBm9vhj
h0eXBv00zhy47w442I0uoqi7Z6SpF8M0X2GPUijVM9Q1M/OC7dNZxrqxehWTGBKH
T58MSGKwxberpX9Md5ZQaWd73bs/Ol3HCtIhrp+bGwHVBa/jT2JQkCjgnNHh9hD9
YB8HQ8zLNFUUVe7Mp4tKDvWKIYUYqf6M6QCcoaMt/MAZTsokyJdlxNspXX69FupO
b0nEnH989ARMs3frLRYh6IzlnaGB7DLBNcPQj0KVNzapUQh1hLSvbuXsjOc+tIFP
2Mr6zLGkR0n02Bo1Qxse6CWYvxJHiZV5m1cetmom+B6F8MDblZ6kKvBSUiFcvHS3
XBOkoElua96S8n61otAx01iFjPbEWio0+i6jSLv0uHOcRY6KhPYHSSMfi9sYZ8cK
jTBvstIf9wwdluJDzr/sulXo2YLjpneHQhmxcchla2uwUOAtLckooipBBc7C1Jfm
Ec+iP8rP44vSWdwFNw82QuKTQowDywpHehBPQ3LT+ZzpWR6IqMG8cMFrjH74XvUh
/zJZ7aSJAeS498X2KSQlFy0PxKelCU2ItkSaEdlvA23uJd2vVf9wPi/pKWtf22+O
cCCu3bYabZClcb5hxi5qdgr5tMH/weG/9wawMdN8bz1/DKEnQW3kbExsePaEPVX8
9zB4Cgyw8WPK/kccigvyeHvFKn8O8gq/LrJU8BMHnA+J+Bh3yijZGnLuzKSyOeK2
CTrHQBqlAnB8c8G+wDfm+hZxhc2AQ/p8dn9QU81w0WOx+nsG6+0Vfl/nSY9uMwmu
9408d14Jql5qwKRjvlh8b2/VXzOcbCtcLjm9z5oXxpVmW9mSFtw6yPzkGGiM3561
G6z9EwHUoVyWPG1whHKcnaOeJfXOExv4+TZ0lu5HNfpiVjBQdVtYeikkpoN5ox2k
sfgmRXJ9CnaK/VCeOYpL6RWdsPO3+8iGbVjxrVD0jKSO9AzrVzbntOHatORg6ccq
qhPrphXkKuGm68t+4+rCuvo2UNitaVSNGFSo7k3DJzdlgcEkVv5dKKUaEWO/1jxM
zI9xKHHT9RQWTDyUADxr2FOm6TmruaXeZeKEej9vtSEBMHHiwnqDXuHoij9TH2Jy
Ii2JVqol9PMNVtEli/mHj64NftM8eN9V5E0nZ3HCUbbO1FrG1TvfXv3KqB/Po3Ng
Ct9IHtUlUkZv5KDMipJ43SpgfjhavkUQqNq9QGJ5uGLzL0IQ5LOXrDR/M4YjiiR+
bV3/iT0V2ljV7RKmekU9UctGRe/Ky9xGr5TLehxYdFNBPM68k0VZlsSnC7QkX+eT
dVeknwgXH6bGNZbd+vyh2+VK/vkETXGNH+U99yn4jmXD06/LNty6kZe8NK9OaydG
+h3hy2pgDpY5DP+hIynzvFP09Arp9oYG5mr7UzCzd5nE6V6SpxE4kIkt0aorTtS3
RpPctbkiJIQJ0pP/QtSs9FauTIhcNC3rKySI1e5dvnOoNop0bvfchIrvXtIrRJSC
JB9kTaa9ThlUbXAztO8uUhZ5B3gimWWY4iejNKd7n6p5pJCXuDKVE0d9hbKAwxsN
/S4xffBOoe6bgWtKo1zaQ93SQBt0rxKGVWtGCKxOEkBvtfL7UPrxjqBqY3q6/wZN
vZCr+HxMYOvWSgiBZ4WnWZzOt1GMDXjNHPAyuw82j9fMD+HN8CR5DelDo8zSAmkf
DCZ0WdrC0HYdkY8Uecphxv+Osid5iXlxy2JZde3CfyE8A9RVM6dKSWoan1nbBypB
Q7koYBGS3GmzF0gXMf/dFc9jjaDYZlxd86BU72Rl2P5mcFp45F+4UZ4N8+yEapgE
CKG+TkXnh3efcj22JfSPIOAiNea8f5CwstnmPQoYDFRpgM7t3GtfvK9jTUFYjZOo
XXewmKORiwXCDljSDziUUCwrzjmfFSybnyJ2IDiO9Fvh7Sv5Pir9La2cwOVLNqmJ
rBpSrOOOUNh7H6C2mCImAYLmtNB8Lb5Xb2qqq6kq9Tok1zDQbVpfQ2usUcBk6z0b
Ouls88Qtlf2hNTmvtDuVMHN2Xt3xXCsCU9cZ523+g4pGsadFzcf2QxsrKmyMPy5Y
2iXaX0SDXPIK7nY3Q8qjEB22cPsAD4khfQni5FOVV9IDT1jRcK/ofX/JTqSnB6Jc
fiCBScmXxnxRxGKJw2kDbRoqBFu5dvx7WJIg94m/TCAz7p6DsBGhsLAx5GSs9XC7
pHRKc57ef7+WQYNNTvyEskQ5vc8QvzRaKj/UNH1PEYsrRBNGdqic08yMCe0mWq47
ha+T0NKJGqmoRUc9NurIdJjdboXumkHeTfGWbsB8dWZ0062YSkvMHjLfo4/+Ht1s
Fg/Mc3324lJltPmqkmzwoib3QJOPUr273zg112orqfq/pIbmN7cDb2cnVg5rx8kR
UGyrzxpTXGZhxGJaAkcCqFJd68+rK00lmlNJNM1s84OSkekA8lgwOqDHcEibPmAf
AUIgCopEQ18r2dxkQrtA8c0NdKJj6fxFAxlw6pAfXCfp7elv6ZkQu1QUgEcjgluH
pH2qJF6Qb0DkocoDzvyScit5fuCdZh7cKOBohztuU3hqmbyshB01g5IQF/Z6D35T
IAQDO/vaRLSy7w8P5wbYxAmLJQIgpS0DjX2IZx9BBCvm394Ra7XIgGzPyqc+aoMP
wedd4Z2JFWRD2jMsWQhMsdsqgrBCmVhJJZ0aLnrrz/vfSylwFVe2B5NzKrS79aZi
e/UmvZrlbB7SGyasVSNLBK77c1qFvR8XsXiLFjQ8UCr2O7Jf7xD1x96qB82dYt91
Acb0qBwenaKDBne4HfQlwbcCu68BYShNt6qzoasSfYeTmW7WeOXBwqXQJ9TwTXYj
eMYbhJzCGMEdSqLUgvzI9Ngey5IEcdYdMiAwhjM57RwauCYlO0oM6CUbPOJ5KYlz
d3yD6dCMA2roID/ez2rEqtejo3e0ZiD1BfDlGCyhnFU8Yc4KRSfAp4AR0lT2i2hA
VoncF1fI3nKX27RAXTGAnzLpBNfqHgj9ni8PsZxOeIfS4eZGEek4or0v4tk1RInc
215eIP0RfXUSvkodv2sz+fPi0DiN/R/P0K3huuJwhrdirqskdH+6vrLDXXQ16K3r
Yn2ygQNyysefCBXvo2a6eC+ev29RnQxG8dbGz2DoTiPukYg+sc6oynfW3rQJgp3K
n8q5jaRQ2zS1wp0SFm5v7kmLyOtKFpTjFnypTDKX0tzmKDnI/+xVEqmvE6JugIp8
RekXM1COhA9wRMCu+anE+qxTzB/tCigzkZ/aLLAqAFVZyMXZo9nY7oNIwpc1gPZ/
EqfOZiV2qUJ7n42kFWHcVs9sd/4RBETQefwkPmwF7e271w4/BnxTHazGzeNUNRXB
CGStoXcK0N1RhTB3wFqIzmljFiaV/CIa7/fafqB/L6eOYL0XfESsZ6ilxLXAy8M/
gMmYO1xuYUvV7EdLLSsLOHrl//+20X62w0e4u2jY87qt8SsKuK0ibPH+6106Woy3
dmdQl9ynLVOd0q1rp2hGO2xEl08ZtDCHPIvpl2Szak+/6t1NT0jIC2lpg/llLLgi
h3bmsNgXf4shbpdi/co/ZNYRlzLmbiFxDgophE+tlDANJc1X77/a76SluNkPsfoO
Sgsv4OJKGXmH8Z692so42uGutLiP/sl+y2WGo2uRmk/SNN4CHrGoF70wkB4JVlWs
TkPwlg/B/PsvrmDg9HvKfUm3ExzbfX3d5WTPa6q1lXIJK3laVFVQHUhGAPGSyqu2
bsiXZkFRQUPe4fxnstki3X4eYxlh4E0ve1DfU2ATgLYpm/Qc7MWpVorJXsfA16PM
Ccob0HCdZTlcPkJdySt0XeWylMXL2W6Q8y2E+eO8ZFxjX3KC/rrdrsP3B98WOmXx
xkrNqRmsmnj87yiCIA8C3U0zx+cSuhAjJYqudV4c5HZccoCSss4eSH+xgqvayq5D
oKl25OfU9FbcPLrlUSPwr6zDTLLKDHmOCuacZIQHJMpfKzrEtVW9GF7Jj2WsmqMN
oV5lDnt1pX49A6qLInzTyiSyvAB7vmpg/dbJVjeOCdFjAeGj4m4JJzcYMzFjCdiU
xtJGsuY/riBnMscr/nYaPkrq03tI6fvzb1qAzqICV4xbpc6UNIOO7A0YsmpczBKS
61FpT+5jV1iv6Vwi5+36b0fdo/RKY7fSju1XAsz3EEJAw/Gi5xTYkfLFQf5RPhHM
gVDsusijuSR9DDr4m0r2pXwRD6NWaXGQ/U3OMZDGksag/bwsPhv0Fku80MVO29lm
5uT5zc6rFxJQ5wZjZ+JR52pYwN/1z+QpuWc6UooioqsCr/q9Yq/q/8DsKoONbbLU
UnMM+/Xrvn3fOtYXZK3Gm+9KbtvY5bZz7Yyd+LsS0Vz+aEfcBHEUR0T21gWCfJsQ
ee8ggTnt7WV7FPwhUiyHCiHwVJLrQGY4gcDma9QXzyysQz/yotsFxXeZbI+cE+WE
pK9t0gAOwU2pb8fNCo8LR6UECJObnoCZVPNy83Sr3NmX5cBYlZmetqxJi7UD96wV
4RNcrC8zyRGj/Lgt1po1e0CJ7o1KwrrPMYxzwEk1QPKkSYETplJyoQhhrHNZC4/G
+06vcog04FI87tWU4NWoxuRbYqJVz0vfM8bUDtLlsi0ao/jGa2piA8iAxhBH3mP1
U5c6JzjNRIfpJZrKkV6lczXezKzBmUpeDqSHFv0piIu3sA5ZCOYMxsshs4MOYTt0
4Elf+1zGB8bXTGUpaiedoK022amcpp2RH35HicslTx7fgTJAP5Xku3wY7wBJAA9e
2uvC9GNWPqQUHt5WDuk8r58M/6Feu/y+0TJnYiupO060sY6DXb1DdidyGvCrfv37
0hCMO0sZq+TzatpV9EOxo2CyAjYJ8r7am7qnQkyZfam0ykjV46caPSIzKdyF9xfd
xFfE/tb7jnBkRlQr9/J8HHXcJstpa/NUxEu1YgbRhSCPb+xl0vhntlKaSL0CqE8l
pZZL92bRKZRxTDdVFgMPbVwvou43kYp7ddJJHUmsoq55CevwHf9vbz5DtubZIYh2
hb0l3snRXS9QxE4+fLAjp7rKeqom4mVwuSzZsZXNRvQ5h7KRCHPf3fy37CJdx2mG
RmS4bbbflcdQCT5abcTe5x4l2RANolfHc8GFJjSCLG3h1qdDu/dT2sDMP0BUPOPy
IT6bov8hI8stQthapQUS7CnepdKWd2IhINjUGxOmK6fNxEV81wwcxQOq6Y24Z29t
qF2CmOEOxxPns1TKqpt910jHD4ibZdpY3XPuS/z8Wl/oDHtM5P1D3sWBJYoxBlm9
dQ+g7Yf4j3D/lcLSh51qDK/GDTz6tERhnWoRPms9+s0rZrtwZf+Kgl7/OQ9hOsSa
kYhiRDJNcrdJoEwiuEXZdwXOOgbTq/PWaJjEQTzkqXiFy3NkGcxTj6mRgkopIfsw
COOgXEalnPhslvMxrmuPzPGufrOeFyDp+m9LuoAeQey+yA/RO8Mrb7wuyHVeVxk5
0E3TftEEiKCcXGld0LhGwz9QzKbxpL5158fuE+BfECyZa8jxi07ctjwZeVzV59W8
4ewTXTOvxd6qKALbUtElTl+AkC2Vlbq+jnvKN1A8wkWjhGHOVH6gVl71/a665oka
asqnWDpnIBVrFiBJhMRiJIvJMraPk/W6ooe7tdyggUaS5EPjgmtzAZToLOR6Glwa
XAWq2p5MCU2qeyU5AIUl5zdTrXK03sWTcV/1I5iDo05Ehz6lyqB9dETYqstR7TUA
Y3hTqQ5axKruFnn9m3fJmA13x7a4a8VsRrj+OOxj2lED2V4L1G2W2DVlMycA/H0O
TnnPXRTXu7ugS0pvapx09A8J/MBxZctHJ44gXcxBKAirkuZ1OwLp3YkvbLdQ7YA9
q+eL+/jV3p8EBn9bio3/f1ma/4uALux3IO8AMSG8EVpLVNMJeWH3R0RXBhwmAA1e
s8k/tWAeucnzGHooBwCYsjQMoNUYZ9RrEU0ZqrHGrf7Z9M5JqkEw0oZS5yqfcgDA
O0hk7bmLKndIkqtQA8X1dhjTV95mh+Ra8TUp6e67K+cpnPn5X9lzCxR7MWf7e3od
ZD34V9SUxITkDc2ze8uYe7gtR6j/fFxI2b2/t3jqVNBfMJuWvRKVbftKiclmgPzq
V01He5LBAOWrrboztLlcFW7HOxL6vcOycyShO9NmxiAe5mKmGtTdMxgxbY2RW7R5
5fuu1dXwurNmyj5lydX1qcn0MrLD2nTf5xe7AfJmSpvuZ/WhXSuV389K2eL+oBxM
/Qo+r3gche1k43gqsoP6SfEkchae4O3IqhUs6aCzVOMpk2TpEvo7xhQjfeuVlp1J
r/+ezTDvwBg+hS0FErslSQcJfUOVn8NnM9fgrLf4wUfpBTRsP43rq4rMo44FdOBH
SsBhXVU3HquoM7fm7bHCJlgFTdmVyN4AUBYJwObUwr3HBahKmOUa4Fst7evawmkJ
E+UOJhy8eHEbyXRt4whPzvU3ZlWBubn504N0kkYVGJ93w3VLL/5n/nQqccwwf9Z9
Xat0iBYW1wHFfvoDFiwVIzuZQAMpF4vPpMBIY3iDqRLQqptmDqM0tLFEHSs+x+tu
kqfVXaDqk5ecqJQ/TStx4r0rvwX1ORDgIk5ceIId2rXytC1kcGje2J6VBQ2qXO8+
jx5uEy52I1OoT/8TndWNVBOrfuwLp2fjeEHikmJJWHDVahDSjA25FrOST7psIFeM
hhVOyoQ9GlT6un5txF6Pd6NdMAVNuDinSlon4os3qIDUoh1z9oX1v2aIuIyDAEdw
HKC2olXhxKG9m44A7/DD2uSmnyhI6t1Or0Av3DpO53ygRSo5za71Jzocc6/E/f00
KxmmXvk77sXqktsEy/FL9N0JW+PHGE8xrsyA7Hr0o7tJHAUcLpLOPvCU4nmTfU+c
N1kiSpGasVjpPpemFxjXNrUbeIac2NOd844KzVVd5hTXsYg3YXewSN2MQuDVHuP1
7WmfxvVhzMEq1mGxvLAk4U1w6MYjLfR1to6XXdxfol86fqJrf+RBhavQVvJCJU7g
pcuNGuRUpTlhGBeTlz+Co/Lqx7dTuDuJ19VAjyiE7llBKcy5+CPfQ6RRIdjTCdQ3
DKtHtylktt7umQYhoWdJwJ6HIx6YvH2GhOlRwhYSNFI1PHGLNaUuUVwoVKIChWyp
nFfCHBPLyFcqY5aUZ7oL8DHDZWcsjwuAXm6bpiWkwJ5tRyvCwnKcpN7z6KgmsgDx
PcYhPjPHfp7e8C8na8kbFxR4w2Lis82Io+iabpAiJrUiBa09h5UPH7pRskr65m4N
yosVNbwWpF58hKslVVTb536yR0ySxOqqj4eaRlFShazfgZSpWQU4NBJB9cWBDThv
H/Zl1qEV5HllvLwP04RKViKeoeVeVL6/JANGMrvL3dgdLFY20yVqjUEy7Pczb/vH
40iuAyVySjJ1CkWdqByxZDbJNglMPKPLvU/FZ8+nU1aDSF9Sbt27i4FSEKAVtTPU
kaPLf+5h2u1/NrbbTHzyjT049ArTYuS0wOydgHQLy9dQpagUqc4M9mU71N+IiBry
soOb+J/MdkmBGFSH8A5q9yx9PYR/0OGfocu2cAaPdEvoABZ8toYlWJhe0X3gH37u
g9h51QHYESKYfsFPC1kCUekBWo394rhkKNeil3f33ErWAeEc7UUgXuTeusis+zx0
gBACYGLE5akmKJQVgkJoKNzlFcYWeGOkj3I636pIw4M/Km9opNIU40QprUwhYJpC
Xo2MAjWQWVhPHAJyFWlkpZFEvtTXjU8i3qM1FMHWc576FepISNb8/mUtUOTtMgqE
qldcRU+L5zi0oz1/G4G9/rCl6qzQ2vzU4ehB7TRhdvMwp7jxPxxd9qOPQI4gRIQG
OjV6P/+wgKMCctGbrzHbIcIh5tO+fvTzx+yhF+77LWHi47a264BsO5+ShQ5zHKws
68Za3zrQXo0OBzaWRyJIvvLMNUe9oL+YoEwbMtoy0/4rIoRB7ziYK3FGI1nGDouD
1Y2nG5R4TuJOloCvsOmvLJ1Wye/+FGy5LSrhbmHZuPuKfi5oTvAM8SHA52rQF8b3
6Nn4MDIpSlpDZs+SBCzST+LVLUXniBVm6K1B+opcH3gYuHOyH1xOvHYO80Vu+IWH
Lt36WtFR8uQEx44y/tF3N8koXdOQLQ/OYOxM92/YsVJ8M7F5u+bSdY6RcR9H7DDo
gd3zQmrERzplB1ESBnDT210719L0kuR8uPP/d9Db62e+6JJq12DwpTkALTTYWF/A
GsrD7EYLnYTkFjqW1+u5l4bwRttNYZh4dck8FvxepbPavm54BxA5Ecxv5WyUBb23
TUap+Py36VjlwwZK7wuwjhas88f++lBvvDsYN+3Qw5GUzBgPpRzdRehNd6Ya7+WA
/Vg4NPfTITz/RtG2V9ycIxypKbH2n9+mV8YA1OjEBAiBDaUK0Kv/xcoNLDKwHtrW
BOeGpTST/WlVJVj9RJrmzS9PQo0yI1ImbihHjTBScVQLGrDknMtpn5mwv+GkMptO
rYfXk5riDeGnWRs1MaWll+WssoxdRrjyTCszq5HMpPTr+Zg4P9p1cKZnIgDM2K8x
X88NbgJzG3aCO2B5HUW8OjdWDHuUkikND+e7UhU41XXdDnNT4OGZdBYBH3pvAvH/
B5n8kryaZREw6zKdhH3aJ+Z93m37A+icJ0UKJv8i5FpTo85whS1HOY6j/oSE7bAl
TAswO6q3XeetAN4hFuBVVlgdJgsCrf3h7lrxNQhgRmglA0Q9z9rs9curI5c5la9u
15P1NrGEHImgABdhfG0YPRLRPrLQkgbr6toFYaY0EGGwq6eUFESWTzxfpzMxDXze
7slLJ6p+YLlVOCvF1wSM/XFAj0B29xdUZCBeDYwisO5r+Yv7EQaP3uKuEl16onn2
qO5gp8HKWPgzUuvbNKZ1vAndifOxYIubLkLAOBW/WiRwR94riDUx/EvRIf3j8YZF
ZJCh8KPPCGlYVzrIHUK7e0RH64BVilovYDTjOfVpWOKaUT/7ydFap6orXfdIFazN
B/MWepJd5WT3Z6TzlLD0MdG107dh8rYDYfWdkRFKOLbOqx1xezfiS2scuT5sewrE
NC4viyvo/BetyMeE7e2cgthspqglt+jJaJTCd3VfP1AFjsofkuqGHfmOF7lihrd7
7sd74gGJzML/Cn2d06W1htRIOlLd7qsSVPI5t6X/OvC1IjPfIxRjGS12dCmza/s2
IcfrOda9bh+65vEQ7RcX6C8R3AD9APYo7Hu/c0eUeps9ZvzMNRPFC1h6XJQ4lnbg
Wh7SbYnEYr0W6sSkNR60xI4wLb08P3QSKBThDXOcfgeiwigrZMZDOxdIP/NMLX5A
UKS37NsdH0/DdjnhRkkc+pQ4lK5UiuYChfWKHHtwd0P/kEd7YBCDasreLrk6XYhg
4XqyuatYn30FMq3F9b+gEDRvJK9Eqiqce/yuO6Ay+oYHfZytXLjHY+LoEU9+oLqZ
LLIKOkqZJeJygPvew7vQYyuVGCgYiv7TKf1ieK4T4J8qkdnk4bURSkXVnl3zkHQk
Uv7B2XZg4YphafEYpoJmqmGYQm0JAqrfDPrx4wfdul+1eiOLeeMoPShBqDx9GL2i
9zd+4BaOwA9jmdz5HpRP9IRmawxJgIQBNcpPhBOYWjIuRMV4hNkiUQXh07hRsnyM
Wp7z4MH98p5XMV95s8kvawj8zc2yqA7aZoygR4T75QXwvmUkebzigQxfuE2iJcng
JxyU7lSwYlr9QVHW+DGE5V+uymvN8GG7K2dXl/EDkcxFsSwXr+KSDp7d4r6Et/AM
nMRG1SkWtEfvviaTiELWacbjcr02cbRgbH8awB18H/cLL4XIkHwpd01aJln/p4sK
VZz4XNLspX/7RppIyDKp1lrOJrX7FD0cIrYJdW3P9u28AU8iiJ5ere8yjMSxx5ZH
/9qCtyvtsxUCDrUH3f3wJkLR+WN1v3NJRzlZMKmKGmCKrcYGCNZnjHUTWq1qknhG
iROTDROCC3p5hTy+WgNYN8uel6LjyZ3zvuYWK6v7c8ZTrb6gMEH16FdwSAJtwoty
gkqPZNCgmV8HMdNuZEd1q0DA3+kPyzl9Q88/drtzGvObOMf42nLO2IItN7QySO9T
A5dXIwJ0Vn7lCbThVgt6MtBNGPMaIJFBUifQA5Zu+EzFFkHeJ4l8ue7hufI/18fs
04btztRPlTz+qpjwXtJ9kNfM1pdUxNvTy9BudswXdLE5nbP1FbwgCCpv6UZTFmLr
89K8/M55MTXR1VK+hzFxlF4ptc2ZT4OUmc7r+0vQDDM8iMGv9bsOVuyAum5HigOh
qwrLVoTlcTW2dJ/Z9bIam5GrRZN0oxf6Vnt79XJJx0cs0ZUC6CXTEkuabuWNzDNB
AgFlWwpRA6KArMC1iB0Z6UzeOgiXnkUeHN6/qjW651466nObV+ESc7EunEUj1KCw
xIMyUqM2vg7LZPZMmVBGrSuUHuZKM2cEnftkqL2g7VJy1/U12j5NPjtc3HKIBDgh
3L7yUeMbExTgP3/erCPbDnpU4xI4iXJAA7u45f7zMjwdESYwR6uLT1ePIlOOUcRY
BvD2SgCBOu9Xei5D8O3z4CpRIYO+m0gMHp+ec00LqaZfpV1IP6pR6En+T3q1eMqd
3NvUr0N313vt1ptIHT5yCeIN0dsn1mGJ8RrjkmMKTPwoIopnWjVfmy+QwfwP4KxX
DdeOzowPQTcmQHUQa+x1ssqVxiQchq9FGePho1D9p+ANy9MVui5ZnTMUYnppALmL
++Ye4hzbIyvfVebjlvH9D85qtW3Wf89jxhSwKzMgnUtNwzp53axItpvxN/rM4xn9
pVxZKRsxXwkxkH81OZwLR88Z0CCZfJ4DfgKfIolKY0A3WW7htYQpGvTS/sxJwSH4
P4K6i3igrbRwTNFbD8RSERjIiBNRSASTsQwYvonqn4xYQ35cmLWvaDxkN4qmwpVJ
n4ddScuT5SlAOxpmh7O6MTAqgEBKx84/1ww2dm6MpHwvHVSHBPknIDMnlqKlAKDs
pvCp/NJCpmrqL4rocGEHne56aaCHMgyGJD2XZwvhvCsUX76VrslP2DA6MK5L8ij9
xfYAKCUKj+FZTGReW886qENCyD9qkWSTnzKkBY4kpkHnU11mYPUKwxztbckoDn9T
q7SFZNE5lznlus2dCpb9ZU12XqxQZJJio//vKyRQFFnDPd5xsCPEXmzv2I3VK0b5
gPI7oEqi2aaoxJGSktKvFe/kVTGCZbRAOuNaNl7OhnCG8qpKEHesz/wybWUN3XEO
+z03+zeBeug31bmWtpHLvBt30V+eFLH+7WgFIrXr+j28kCpNU7pTtBzX6L1eoauc
jWQeGDUKzeAH60iX/AnxmvZf2YBqDdxIeY90B5ck6C4vsJaR25Q+6bKXjDinlvGv
6Mm8JJsiIkJHXYse3bhTXkJ9wANkptmfXptKLaS88xhGaBPTjnZWm7X1MEhun7az
KuHlK2ldOF9R9oknfL6gJdB0I/THOBmw6zlptW5WhfvmHj6WhlYqaMm99S8Tx3C2
cP3/2ONAUtFuNSoQQZdmxzd0QLFazTGttgpxtyhuFga+eyab3C9ZTE1jZFmJMJPZ
CLUsaseVnDn6dV9/9qQhkmTP8o47LUx+0gmnwtbynIS+DEY1YsAQ/vgJohW9B4x0
wgLWCwyYvJJX+sQW7At2VC5z4FwgIwxcOwT3qYrn6Ni/l8Nqil94Izjo+S9QR8KN
LVaKIHaUMKm+kc13SaO31bFb1u01vKaKC3so2k+mryK8TemLsPkpocErfY7qZYsP
aIe1zcxeM1NKOqcrBB7JgO/lBxRbP7TYfeDIwMMG7m1cS4/BtWsHI5CXXRnHyhKD
vGVaLKJt+pnRyCAXbvtW+WCxRrET/2wNp6ZgvA5WjDbDWpJvEIIN3ceexBbWAFa4
rzY4+nz68FlkH84dTP7FNQKNQwOH2t6OBM6/AW1otvD68iVvrqFlBQEUWgOuhLMn
xYVsu4yJ8W8MZrHZY8h5Ib5e2vKeyOoRSP7WQvtyrwj+H0FEEAuiYvSBVD6xwlXv
wOHx1fGg2AXFAlLun+kzhRBTSwiu4N3+vqBhF0B9IZKj1YF0HE9FkGrnd6qucIky
+cz6N2ac5nMtUXZe50aCfpLEahbI2GcZAGMkV/mTim5yakR9zxWAZLIwu5NboaAR
/PfO2eYLkf5FtZbNFafaUEmaGGcpWW2U/CWBb+HSB62atg+D28GBQYKlUzoq1+85
uDVUye0cyF+I8NU/9VUPSiNGsjDWimS9ux/fnYYRLF9TUgdaNRA2pBmWQuNX1SZQ
sbNCwN8uYa+VukIVPS2FW2foSH7zefmmcDuC4xIO/qU0vaXJbZf29/eIdrophHw/
sa5BaLPuveC5ekJDLYGbiYb0UDGanM7boYwQ60+2RIhy8UclhXaYWM12RkzYeqZ/
RR8c5yXtw1ilz18g+YZaIRmgyYcdFz76oxU/Sw+6r5QG26Kw3MrJJWLB5WMU7ssq
iEFfFqoTVul+jjU+apXqPArO/1vUMiE7zEZ9ISls5IdgM632aMCWaPvBDAPp2JrN
VhhP20aaVOPyJU2SwgItnnES/QtsDZTg3sBP5vL8qtgFI7dM/bWOUKzr6Eph1ZDH
SzZapfY/4XYx14wo8qzeDlxBatl0WzMi65yLFKQ23mGwz/0k5DHInr3YOCC7bppw
wx3VN1rr3fjCPxC9+xDXbewCHmwuuLrH+U3Cw8tbHN95nvqCRMyx50D1Ikpp0Vhh
XHtYF7bF/yQtAk7hW8Kw1BzyxzfzZjQdMezP9hGr7DknryNmr9sx733vDSszqXIc
g5RuhsmmwHhGbwffCpj8lKDhp6Bdg98vdZvRu0Ly7dpYXOT0KPNtI2N0cBvPray5
xghnW+CUfxSmKnrQpEidgY14QsCirvosVCyj4G5zr9Lcv5bEMuVmoUHH5SnHFXCP
B7TO8nAxMrNo1jhfk+FC0leozwq3KM24PRUX5qfi0IumPQjThoUSVyAFcibJajvF
bdJdq8Isz/8yXgDp6Y9mVZnH/jeg0Oejy94OtSBZL+FtYHVgLAXHv7hu2uFoityq
InEGYftMzUDRbdvinW6aWX1sfXLclHpcQP69MYkDX2NyUbB+CTpUQqfBSagO+CYS
J7a//2aeL8zw2YtwbtWt/FX3gwU8bwmgBrPXauPN72FSCl9EpaoIkEzh3fdiS20d
lP6gV1b+Pm+fJZgtc6dyWPlUJiYAgXiVhEhwj/2H2vXGn3Mef4AjfGivigjwrwoK
1HpiZD7c1wcVLci3dXEjy3wdajysUt+to+GdbfXvRkQB8/JVr9IgS8sHcA9hduTa
GZa5hk8kgfZCmOYk6TE64H3paVXNZ5z4GHsyPrJpb0HW/9n6tcbqYzAME9W07o/3
VNlLMunfAnDlg2jPVY+jdaoz8Qo5sJZ5h/wsHlLo/Im+vwaLaj+/22qd1D7UP9VU
ESpyJ7s9XSV/mBgyoq29Vu9n2/ySy/9L/dzU8Dl2Q08A0WJgybGBcO+mCx1wp3x8
hLgwckOyupwQjta0wlvuPQ8WywBSr26gYn0RvCpfa3Tq9mm/9OAsUbTakPykzW90
AUFlxCDE2H1m2OsJ/x9d51BuXcgSHhN8ujq65DL9J+6tE2RsvXymU8aiTpFDSMKN
+hpw4PNplT9WLNSHex0P8d8UYWJkzMwwBAJ40UFqjerehUZ5BmvdLTHicP77saVj
K/yVYS6+tfpnXL/SPv42qYz3P5+rnF0cdxI9A78SymGqX7Mggt0sJvecw1m1mc3X
MW9smnFIxFq0LBcg4WqDgvG0BDiFpvE9y2LBE/arNtVherBfzRJ4hQvz3NwsPuo7
uyiOePH/FfLezCZP4N82aKpY/PskZZAMUaaCzdm1Ax8qND3w6dpvzCMS6pABQK6z
KkQDzhRX2gFt6dbw/TiZ7ckA4ut7S73rNioTMLjk7xQ+I2DQajsXClkjnyxCZ8sR
h8uEsJc2SThAzwm+3XwGi5Beh6sAl4vLhojuAdCcU4AAlASX4d3S0YgRX/diSWLg
w2XMkEcLGUK3rDjakh+mrGNX7d3s6CwBA+Wj32a19pmffSYdAIpaCV60W9+XoI0u
hDurzMRNww1FAbX6XqMck0ZMhLndA+nJ6HqHETDIge418SHWmbnHnFuqsA96sOTy
rBBAjuC4rDK3Eexy3ZK4A6ax4vMQM1gQdmLPnZqcR4+Z92tLcx/W9nzyfggAjO7u
tHb/Ak+tUFYlRt78A9Cc3GnYDPmnKOQ1qxaxrfWx/wJ4SEWW+H+mEyWQJKw/YlDd
eKEl0+0OuWTmf3mNpizOCgu86aN8LluZ25gCpjJNy5L29xxfg/s/HBKsAcYsX3BR
fDcBNexhs9PRs0skCdVWi+ki6C174jxfpiVgZM25/tx0nLyWHhl4ma5o68XS+gvr
lJNTD1bxx9LeDrCj4Aod/C+COiEiJ8IDyzliDJ29GKesyLRJXCclPBg3pG9rxhYQ
specBlwCUqaFfoFb+Q1PzNYjfqzx66B9OFf3FHGDFNL2rwjbZEzlVDj4WVmpRiTm
7URTl957PN2PvxcZbLHEpWx5kNFEGP5+qo7x4b+DAYbnFe7hCYWblP2UUlwJRQo0
o7dN1R/vNjABHxWDaKCYH3+SH/HgA5KAvq60ffQoAmD+mH7NaQxKbSho9aaxF5xk
T3xPInsIJZp1H+RqedBqBFP+BgBbzKI5mco7gIkSNU9T/ESWt3mc7dB5JDwIfP2e
VuiErgdJuPRMheKIy4qCfVBkZ5jSNQLQ/iPkkLm5zUOmSNFs1xXaJRqEtCwIwVnI
gAx3WlYMf8FIXWY32YRVjFo6EgWipvHSW+xXlR+wV2DYywtfiBmThuir6j3gZH0z
a3lnkYNKz16EevZxdL46kVvhE9KTt4M2cDd68KNLaqGy5bCHbY+SKu5KLnKP3jAQ
qVYorq1nVk1DfoiFnd5WL0Zlx5G7CsiD87NkmjNw39yM8Sxlismikr4oaasev4H8
qIZFXD1y7EygKh5z3E3BIgU+FvYgMVeg+wkoWBc0ox4a0mVa4t2xRrEA/vp3sAFg
OR4Wjy+t8Nn9lb1gW0+jymDQidGYSuR02LKTG/gKy8+WFObl1knCaz4IJcgpTYvp
p+XbnELpvHOS0gt/pvDCh/3Nke7XUyghtBzV4LJGtmGT5OEttOvNkpaakEZq+TPW
78MMBMgk1uZDuo6nYqJJvlhanVCUht3quCdQs14Ug6YNsH81nUaqkYhSuNwsJOOL
DE2EWht/kMPkFj2PT/LlzAzC6XDi2JQlNAWkRWF3Y3ea0CZWwdJ8/W+T3UPQ7hpe
MRP3mkh/1p+hKuyiXNrwJTzfvsLiE9+v3mD9a2g4gTUavKwlXDasVbQ6UsM1+OYW
4xG3GxTP2MrFrp3V0s9P9J7PfBLI/LVLv6Rz06GG+IXioQluzdGpl1q3mWpAfk9T
6zLAtALIZ+qhoT+Fh0VFo+/M3kN8/J0a0OMsTfS93ocSngM/9nciDuqUT46NCVy/
HVUf9CBDF34HL9GBHIO76MVObBiXLUNJUOiTCzuFpVyQkf9/YJ0PHjqf0AFEcHDk
sqcWm2Vuuipzj6v3HFinHPpOK9Q3bfxxpyhWqToyAbE9Df4HDjp1dMgysF0Dvc0e
GKoplwKG3nqNJHy5p2oV0o7ISOyz6RAjxwVlsvKNGFsZWAvVxzHVtA5kS0vKmG/s
r9DMq/bInkXDZfEJeZD/HQeE9rISupcQ1o78vzJB/RMDG/Xn7WniBnmNKR9LtROB
8T23AitxDz7XQqCB3NWJQo8hV0scoa0Op8vRG5/nJra527U8X08d9a41F4M5mrsB
EvS5i5U3gbmVFjEbNKzaeNWAlFocifz4VeC6/W0y+iThOwiN4kj7bzYg+4H5XbS4
EMTooqHVI58Zs8IEhHDqlQZIbsnVgmZb1CUKiyD49cqD8tVzjvDfocZtVPg1FV6x
JXp8XI3lCO88lMN9VlGDWL//BAZWY5jxlJbsALhyuKDpaFTg5cJ7T4NkjW0Irn8D
AH4ziDbgD1hmF2wh9JTDQ0Qe+LAtKM4cttjXdu1rf6Wka38LGB5fXbKHriOXw7hK
NkTh+wULCCURpxaGtQojNL1lYiZR8fDxqShlV1jV1SyW5FdHAxSPDe89bivL2hsy
bE/OSI6gRdDc/xsg0wCtEr2F0pD3I4LoXNPl1IVMcYNfeKTX01KzBdCvUEhB3vNx
GcMX2wBGYqfgV0zJSyorzOpbgELkmMqez6ZE91fRXcn8c2CY/julQ3IFuIk5oKkG
O7DH2KuieVoO3XFI784ZHovMLwH22J+zT3JB/PVmLe+rKPkWt8yV36+6mzBJi20X
t0eksH2PaPikG+nx7PIuk2vxRVkJB6MbwFWCAPC661lsyiDC2YAVAK9ZvSXoDeHh
uNinzArmF8HwZHSLlHpCuyo+hZYGytrNEcD64a+cXZXaO1tWl5BsnMGBXE0QKqNs
zdWcAan2JaBaFE5fbjU+DPuQ+75m/+XgoR9+96vlqYqnvyNT/eQphzA8GyZdh0cC
aAXCSNK6InfyLEEdKxAfgbwM82hfJKwoh1ZgR889rJIPgvQWUiXvEquzgGbWBuW6
uty1TjG5VNP9bLNbfnoFdWVfSXfJ2G+AnLJyTrMM6pZofq1oMqPn+2wZKkEV8BYo
HTGUkH3FX7ehETi7u3BYu1xHaeJntjI45ZWBv1P9OOGyro77Mt64oeAzNsxINjNg
/uXOWHKoam7/st9CZy2KpeX4btjMZCsgMsRA5yK7d6H37WfLdSI0K+ZQW36IiC/7
SVehhgCENPBdLa6b/9D2PZHW9Om/1TkBECTIuX2BOJAjrRsd+KBDGJRFeR6tTbBl
MNvRDYyhb2sPxEWo9+sisf/h6LbDcV743qg5dR6fuIZX4bO1zKVIuogIyzI4i0xR
bccaeufrMeCNXTSaPmb+UsOzv0ME0tsrgCIgKS3dV62ZUtiqzjVXuDbCfrg7oWxh
15eZ+7qHp2jVH5StLpsm91m4cWHqqvGatJr/9df5PchTbpSKZ/2FBWh26zsooZXt
+SC5/r/lT/RMJzJWzJaG7XRkC0U568g2fUAYNi+Myq/ZX3qNYd/hOR3toy6Hy5dR
d1gPXgQkAlBtkMNOaBfRGxTAPP8xEtbE50pS6yooBG+LoqPwRsQf2SxEOmKcfxMq
ymNgs82RhjFC60uupw6Op2kxMtxm5MIb0tmvMYDKlV/KLz5kKR4dhryu5Y4UULEb
Ykwwn3FJUUnsjrCy8r7hT1kT1dcoaowaVDBNcltCNexZYG5Ccf75zUYc0CXiUk4E
qjcgcP3aWJMIkzY4/yNbQugFHTIaqAHPjlVjP0bkn+YcANZiGcrr56NjL/MTOCi+
iROESyzkNWypEqZIAQUwa8SLdtASkACYDWgSNOgBgJq9FiS600TuATQ8/QJQ0aLs
ew3JSLQEayn6KJjFJTHjbp9xz5HIy+gnDkgZ9+/zRT8B7tFISHnJrDvmB94EOQwY
NYt3SBy7YFwVWW5vOv5TqKmkgLCm0mnCduKKAVEtCGZxqQNAhVxZL2QlCte/c34U
//sMEjlBrx2K/GmANBZST8/Ch/RZ/wOa8z1JZ54DCj7p9iJFm12+6E7IKM+9/KPy
KvMMg/A9Oi6tWET+GDuT1hd30fHWZheTaeyQubWrFcyfMmzHxg921J7nAHa5MnU0
AeScoW9GgMWodZ7yvjzjjQ==
`pragma protect end_protected
