// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
HpHdd0eQUfHM3BW02lEGRWXJ2jq+zZLdDjWqeIHUx7gCsFpBI0mKAzJicPE2ITaTjEPH9AyqEnkx
d3Wdg5S17JYECQbU5tqUPsYYTaFW9aDADMTCuJaBMiNmxCUuyMAIK26YY6l4w2UtzbBFHj+Yi70t
nzgXl45i6DEsubUPgK7A68kU/6UtA3BYS2d8R/q1yKBsg37nh/hKwsIVwI6jiLy6O1WOGSHLcL7R
+jg+/XyxcvYhujUSlkor/EGqGiwrdv4U9OqSIBNa32ejkW2WH+1Y+RFU5oc99I8qcP1tR1GupuOF
iMffjSuCPI7WV02YXIMLMhEw8dRH2VpNU+k1TA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
MismpOOaZzaZOhirRhTLank0FXKJ4aqsOWy/7XVT/2wFOoQ+d75bAKzWbqO6oerfLNCgaX2GACHi
RDOqpUCa6Uz+RDU2Ebg13ZpJvsd97i3My3euozluI7ANwGvSIAskqW5R84NTFVo1x+nEW6Ab2oAW
WO2PcmVKNqmAZd2aXI1TSB7WDKo+DQRRIwDf5n4qWnt2TzhenWODc0c+Cw9j4LwodrkWiZ5Eiae8
4OwRuE3FZY0ZSW0Xq/5Mwt/Bdi3JKiSCG5XKlKYThIDmGy7Y4ne1RSPR5ms0hxH+b1RzDGHN7VZp
ZuLjfT7NU3fyDQiiyEdXiJ3/Krvk48mN2LPCATEKD25GclpOclQYWYcn1zWLssIlzDG5gQXA9szU
8G1611KRRudiLX31nn/mijd/WgRoANLCl2I6DN7Bmf33N89PEa6RWQ4DJl5H3C9qBqQJYIjG7LZF
RbiFxrMXiEacXjvL4Mutqy8/YDkqF36Beinnw0+fWr4PPKpwsfaBb8dZFz+u8PsTHLPvvtcIAm9Q
4M5NJhRUcAT1OOlnkDrZTwhA2IkGR2c1LxxYOOkblgcRhIxOoGzfu6Ecqqpk7t9e/cMB2U4QigsI
mGweFBJJCo3Bnq2av3N+moyiDWjSeaDGyHe1X/ymv/fTFcsSiHSlZGLHjt/hWshICzWg3vqNndoa
rFJB5TSvA/JdEsueDTx4ldPn6/SYPKa4yIfLwaueAMzAz/yooND6g2CPFwtmc8zsMe/BTNeAqc92
ts8p0/RU5PJAE/ecyH8IDaa+tp/KEGfvw9vywLZFSOY6SBD5LWPC3jSc6RtA2hWcEOAjj8IiaNTX
cPaSS+rBe40EX0LEumot2hLHxHKgvcK2V7etabXVG68OCciqSgJ3csFng6yaMyz8LuTuStbeHE/t
Cdms002hMr0RlUa79Ar5nsNe8UAUu2ml6S8KLAzuioqIERdIVAQuIJjU94JKoEmqCRu+t7bLuPQ3
bPK7qJt9BObn4wCNAmpi1IPbf9EN5tYtnY4S9UNA30NAnNtFO/rNLX6R3gh4RBfCFQ6CtEbxVz8d
ftYXPK78q7rG9u7r4CbUpMdJkGT4v9oWS3hKISAgek44YuH3db3nNhKpqd3CVML9KDa1XvUsqtdx
GSl6+JqmrjXs3SrvJkKjmc0iK3OcESTEDXyKPdExKsv8a6sWD5lMC/sfiVmL5aMCoGoHAUlYXHlX
7lK6T3vuVimxUe6/QFoKOfASRL5j2B4vi++htL+cOXvGHHzrasYajTEZ5yiBsgP6qFOqdYJydfwF
DIPTqufrasdx4cV6dOoRK8IzfZekKee3qxVqIrT8OXOZyR4tnNHDnAbJ2AwHEMd8O9pwwz4rw1GB
iu2FhFfQTJz7/4ewtfEUXnMCg67y7eiphIJx8q4F+37r0iwN98UxLxII3x9siOzGScaTFtC044lq
hUgRLD3ZfZfawqq+j+ltz6n/T0UmZDapD6LRaZ8J+bQbs79KBJsuj2j2zgGcLSB7o/nNRQqgOfqG
/ZTvmsQqejAgtKQ0fj62lmqoyGR3r10Q0shDGZQOx///GBwv2+URLAz/EmjZ8RDEzTZ0FQ+vqlzk
zmoZtVc3XRIofg6AjqqOTsZeQO+e/fAVkiHVIe22KkPS+BhktRnrlXHTW/BvcYCQ5JjCYKoH0NJ3
42sAwSa2/Xw2khqz6MKGIHz+Ni71oTEroXMsjoUJenwtGzLn9TCdIhDfvD3Vyk+lED/IOIgIf4AU
PTXiw0m31q64pMYN6AAOdwwoEyB1iDw4Hti5dWR8hlpjMhqGc22LqV4TM3UTD2/PqyKhcXCTl5nL
AumO+Ho+ezqaB+hnI2p2tI9YaLV6xslCm7ZkeowsnCgBYUVhfkMlf5wPDZlWof11Uv3zxL8CxCRW
QUyAtrQ3n1poxrMks1bGGUgHXsNPGsHoSjlPj1IQLSjBRQ4HnWnGVjsXqn/z1JWRYZM++LsrNL4g
bhs6bnMtSQLXadNFXDOht+HElyRZK2WCQe/WD0wha1nGcAjqONLgiWzwX9CqTs0ezC0+O8zvBPwx
H5KRiIJstBn/ivyNMJhkW1SAgdyJuEi5uXNiBt/YT2Ou2DEMP/XXW91fNMWqYFkJCgxqcZ+p4Ifz
2VdixYXyB9bV/XCSKZ8u9AxbFV5A6XATAbmXfaBkfvo5HECOkzJDFAKBpSFXDNMh7ssjV0SQ1epe
xmscctwNdp6O7xxWwirvkJWQ7Q5z/VqQgY+W0idW8SK8/1/jlSK7NCAbuRpnFPEXHKHhlsDZbA+P
zbaTNwzkK0jsyULhKIIEAJrz7Rd3JaMPfi7+J1z4V6/VdmUSaDD7NO8L5Lp2DTl/kLMEDIhMtdKe
Twdgu5glI4VTXKbch0IrPYNNP9+wPik4QLw6zrFOKzLFBQV9LlNxzaypPjlEHVig/Men7MZozfun
dHkcBmOW9utV0r4524kZ1gyGn6M0M9f7zAYvSf4CBo/8sTF38sjEq8gto2v3tqjRNrnWPvZbnai2
cvJfCaq3MWMq/C2/A8zQT7P/XytgRC9l6vjvniPYGmwGZW/Fo9TYCpOJtiyrEbpsBOFbpgXz+lk2
qvn6T5c85Sc7Wy29+cE1nS/gh/WYSFGIrjvq6rt0XauQc1d+SB60n/0886zOu1s1TDFW6EiStfpT
ARB1Uu6IHkyn2ELyxzCUZvU3CjyAd1U8kLuACEekpjGNGQVp0R5AI7QqlcBrZk9ZI7jqtTcqgoiG
ZpgolxRUQl73hIlPI1j0eWyvrZKMKsz3eoiqP/3pymwdrtZQF/JVtgZEUxfaPqwG2BBIczIayPKM
TdD/OkNsSDcsDX6Zmt5sOT2zZshDwkl8zI/TTvE/Kgvd/ZjweJKOVb3wQIMOW1W1tdH2MesDukJq
RfKoaqo60Uo70UMHlPvr5WGwOZzjkTl7fSiGmT92NR9S9OJbyKFQvQ0Hep7g/LR9gt5asiW/FAlD
sfAKmH2fHJOvHmLCJiTU5yTbcsFThnYpiq8eRSBdOrcS9gXpt92aiUA/VgxvVVhjjg6/gO3Nwvg4
Q8eTAxaMnx8t7cIYRIyK4E/Ou+xEi0Uk6//ZmhknwwzzeXaKytbUj6YdhEoOSJvx+S48jhH8Qfa2
flXymbcdttPD4c/XqM58u9RXodxWqwsfqYgsg3y66um//MZoiNPxIeLlSTLLwy/z+8jph/3uRLvQ
Ur5GubFS7utMQM7TG+IbU9jWSp5yn8siohb0vP8ngNQc9s71Opjqq51MXAYtpCxFBfoYAU1kYGKx
uCOCASpcU3TUdW4ELW3eremVEvxOtUa2+6cHMXaa109ThPMDXTPLtbYN16SBoqFwPRajOt9AX3F5
Kv57gIFHti97bD010wmuONV7E/rUibZ0CyQiIW20JdSJJLoxrKwPHcjij/uZp3VUBM8PN+pIeg/V
KUqmVFtWBRVx0+ElinIgcuafk7Y6lXft0VF2qbkLfw/EYdPwaa0vkVJ96wLKOgNxKXhLlBsJubjl
1Uz0fG2jhdD1nIjBsu7ATJJ6ak/8Q+eb3X7TgMzmh7HWIa3ioGMIiKPTB8I+7ORNd14WAhxUHfqQ
ZefY81Sa20cX0jRSzIDap3akqDTEXoshuzrOtCW8u+Dja1lUjXpljiBBRq/9T7i4VXZ1lt6Ldy4d
DnyLClcO7PtWAJEAU2upBeiU9Sur0jtRw2KpjxT8/rE+/BxQuDv0I8ut4XpSUrhsJeHak/RvbIIk
NtaWoIdX8P1EIcOjW+ww51KHv3F9jAZfnY0w5STJ3Zz39wpYlL9Zr2ie6TPROM+U9yOEZbXoCG1e
cFNjhpemoijqz7BGn+Rceixc92I6TvBHjdmWSwNVBNY+69wOSszY0cSWvrTRAPsFQqAq+6N3VMIo
EkChKewHWmzEWRrIkpRyjFhCmEP+BHPvt3N5SvMzQyXlHr/D316iNSWrIgnDND+h6OAYJ9DKp0zW
f+aBzFqFDI0snYNFstF+hnkKvFjuwNxp5knFXQEwM0S/WY75pTNP5wHec5tQKb12yAzfcWokUIBA
SL56DLKUBsh2uKcmfHVfwdZja1viu+A5Ld+IhkeY1uTTIXBEBwWd6+pRTsuNmVDfE3bdrdLu0hV5
xvmjPK5sHK5EoS9IuMMZg/CM+FpJRla034+qverhdkMfGizo3ydeNmfTuYLDgVTnECyt8LZ05ndx
Kjb4of9bKI9XBX8nft3wAR9Bss5bOwESnVAvp+R+ekq5SUFe2FsHyQxVwrMz5unbY5MEiiHAnGpv
v47eIAIjq8uOKxxArNIH8G3C2uCZflrkvtMoRlBqjTry/Iz3ZAVgVhZ4qHRO696ZAlz02fVDC3w7
0p7xR+wQpV6fNM/e6WioTmHuHFHd9+cfrFFjvnBBjbNI++KJTVhc0dghW3FpQwHbP4Ho+u9wxVhU
jQcCaNukHSPBEM/8V2Kn+YRmQIxRcLqBVSD4iC2E2z5Ne3S+j/GloiLRPdk0kHSiOSpegPZHE+VA
azG6ManrRkMb+hwRQJ8/GR/9ughWnVqXwLbIlNZV4msPPqo5G/qqc/EAFCH+fv8aDnBh02cjs/iF
gdA0Xm8Ge2svYowOExdu0lKMzrqXmBFGAA80K6MrJNrbQtYGD2ud4SsvBKX9fOrAyW0CAzFw9vj6
NxYQQR59ibvsy1O55vY65kDGAhksAJHZfH7DOJyz7A8W+lP0QS0/4umrmVX5jKe5BQI1xqm+b16B
X6e91xdrHjhr4wLZ8rTxoVtWa9qAgbOzQCo9tEXpfkQgOtzqeWiFdlWUdtYRHCNuDy2bhkyZGh1a
hjWT0N1Q5LBDX76p4epVtdX+GaNwV+nCjxjwyD8ZeD0rssC4MQmCmRjrEkecdWm7eQpq+N/UZnXP
R3gBQThWUbggUl6w04idQzrnUnjOoLMceReFk0BLUiWthO6GxWYkvVNJcGJzuu6+eC1OSmLx6qgF
5ht3mhBfw6E1ylYHPlOZbMqMt+O8WKWRUC96DKBVACLqy+UZk9QAEvTFko1tdr7xIQ+6XNNrWyzi
+q9ZRKrxFmIL4SrE2Y2HoocKHrFPjiqQvsT89F/fl+oYuJxtxlw+npLHr8rBrs6LkAyVF5ztG/ZB
/gLWGT27WFOjidGsXrGKn/N33s95ZWNAtm7+wBaEJCAJ51c4FqpdvGWU2DdxMhNj3JEQ1oVVcVYe
u4Gup40Cp0ZFzEwd5d1aaJsFw8+Sr1AehopTJeCHZiwzHEEzgKycCiD2cSJjpTjsv+ZsbY3BV7x7
NbtT/bPHYs8Ls7VBjlXNm9HPxJFuqUVxQxwdRKfEe3TcIC5OKcyUqn342XAAduiOWsvrF8OzVmj0
u+0lcgoldJff/Akl9UVYCpfZDjB4h5LqP27uMoOGUOIFTz/ST5SdQbU+utc5MBBPTgHfp0RhvRmi
qRU2rW/uganFQK137bwhOO/RVpRi2AbADFnmKPN2FAT7svzglD2nB2iyTFQZKDoJZ+U0Mi5K0/ut
d9ICg+RWyXmIPZ7SJk8Ucq63lv2PpBTJvdznuwK0HN3BVQJR0Cmj0Hx9ZxTPvcovoemuqCztHEAw
cq73xEei46bQ5xSVMkqd1jv2/XUBqJIwCscbXuF3DTpYreJaQs0cD3m12dgt09a7+PaVYb++vK8l
SP6/Stks/lV0yA2i0FeGafJhmwcrzOavJ+RyZMXjl28FgSOZRJcXtIlY+JUSlcl7KG+d2Q44gVts
iWRts7QWnp25Ztp2fW7tRUnx0irap9Q6Qiv9viGwxixELwAUg2kn4fSX/ng9s1gtJ7wRcCl5oVum
Umwuqf3ilVM5u6xjkhrR4IQqjVLdlTaSPWFSJyMRhgnrsDtNKbTmwp+cFWkTC8D2ARA+PaU48lep
UqxK0cJq4FyBJHFKeAHlwNDfoMpLNcHcPXn7941GstA03IRDd2GXDMqjda6wG7gUseneMqCloWyD
kLYimrenQIbmhHHPo1tmXX9QTpWopuo6bPfnYsOARwpFObgaKAzb8sGQt6cq/ulx6RWUPi96VxbA
QQ+4ush2HPk99IeLAzo3eUBtT5dRucMIAYGij0T1GnkOw7JAz76KVFY9SvQhlgSOjuTaFbDtFtMf
reIZ/6Lb4Ul7c4rWqEMqM8GPwQmow/7uQKX8E7XI6E11ZTaF5KIglBHQxnVL7YOWBPp9X7P+AeJe
H9Cue+9TWvGWWgFU9fte9a5V35C7zITOfQL2+pCpwJpvN6CBdypOngzIb3tOjmuU4TmVIBjlZyz6
U06coGpLrqdC06rJ0iyrBu1AJ8DPmIZk5s0CF+Lk652DEWYjdZbQsuTEk9F+1rwEvWZH4hlMKAt2
LLEKoRcwSZhISzTIj9gCpKfKyzK5bpJKj1qoWZQPOZsM1dwZLQ2JZD4I1Bgi7qX0pXocarQCCLp5
WQvQLxQROMZhZJwg3ohNNq9RkiF6yCmrK2h/OgFF1yY+ZDTqzdxnFLA4iPbYOc6jb6gUCw9DI0T0
DMs2+SR53RfGzdOFYZUxMjfdtwpQHaDy2Kkn75XbihzE0PQgBp5BW4QjDLS8hUYbtdBwOSV+Mx1L
1zHFX1FlhZLIs/AH4ru8lT+YUxCOg3qWOBiF1ODYppK2Hfe2FjoP4xJxjSdrGDT9W0Zrw9H7Bap7
g5uhv2xpatsleHn1+5rKMfa0uqyyhGbDs+Ya48vETGn7XMESuLdBNW8ovQ76jH3a+UMZSwp/vHmd
KLfueIr3lskAZtHzSqq3iVa6Xn5z1ABL6NhF73u2ElydFJsyj2n3MWhz79T1PGA5FyaD7q0MPwAY
hu6tpXfXHpQ6mmSFjOl5884PqNN7whuEl4HA2FDJDhtLQATW2GdUf1QxBcrqQYX0AD+Y8pOSMTJE
1aj0b/1p5NweZQIYvBCMLDKou5oIP7kHxbHlqFPgUV7Pl5IsPsIP52w6s0J1gCLc2uz4pSSuNBPY
0XghBCJWu0yJ1Fm929o376gnnB43l/+Emnno4AimoJkpn2P9Joezwbadjj7fzbcG/zRxscwYcRPU
CyNDIHn+Jt3wS5IzsY0V5o1lgJ0Gb9UwM93VoWLHzJVRUmaLv/yL5XHw4gSrhQzul8caeyb4T38u
pNvXNtwh4KUyquUfdpx2pJfOUWo1Qf9V9UP+7OBidN4gvn73dXYGOAGu1k2JkNxMV9MH77A1LFlH
2GJYjrqX2WCRJqnyhm3EebxceQq27DVjuVZj0hu/gp0VwX9Zo293UOlCoh8w3hwBeTQ6RT0OrQXW
th3uUhjg8ocovIKW7Rj/CHkmfboPDlxP9sPVD0X4DQT+fzCfq6MTp2swsuoPuzlLYXq+aWFT9zM9
Cwfq5qHsoJsBFzr5nVdSQZbTrmryAwz6Eaw0SbibBl0rtMGffsBFS6OICU3PbY0B+frLnCL0EjNC
ue5O7EuZGsX7bPM+rH9sI1XaVPXcJXqme3bREUGLbP2ieiWRHTYsp6y+1HrXXT4qBr9Xf2on/zlk
+AS4DVYFveXHMTIw0zMa8gHBl7Kmyri2M99wc+kho3NP0Pj/7d1WyJ1CG4c+AFP9l48CPghx//VF
welplr48YvqO9Mp8ny7o/Gs5NhSLIUUzSZrDycahefJ94RRwcURfvBuNdkM2Mx4qnHi+NZ2qIka7
p8EX7HFywNTYEFJ6MJv+g5wsnr7PP0A4tznILhcUgVHLDv20fuqlXnCoEn+GnAxXrj3RxnaBY08O
eHACB/bzoGem4BIsB1Htopne+BOYHcCkOiRegumeW123eeneyv5e+xlkc3Xk6EQeO75VnTFwrEap
uEE6GGfbCCVpo/QnUnvSOwV/EIH9vlA4Wd19EzXixUMS1MD0OeuTvjMWVNmEgUZkjdeAHdWfdSuo
12dg+84Ej5emyqgHxqpPJFI37C8TTXkWFZPAe9yM68TXCjG6wOOh7holBOVNGhJmcKu5Ev5UNCkd
hru23MEmW8cUKZY5RGAlD/HAX+uVSzoqEtIlPhGYSYEA8Ra/JAlVxg03VT/uzJ+fXoJVdNMM9Nvu
BaD/zcQ0WNGVxLq84ZyLpfljqY4yy32QBJNCUgKytawld7Eh7RsJjXP+qvZP3j7Dxcfj9HBkiHoz
dFEzS37DSa0LbgYKhbe08SbD1hHgOvscf8nPEvZyIeWJfe22UCdizFHlvZToHVJNVdZbXWBpPSSu
vTUQZjPtZ+PcinzgGTWJbHiAjh6uxcodd5NxwC/nbSeA03WuxwoMm3vu51ziyIY/wvKEXonR3TYh
GR7MshY6wfSRqDBuqVyRBaXAQ2mCQ8FVVRRA9QnOmTnGJRH69C4dBS6vasXsQK6jBP0QGmkk+Uh3
Fd9TRh9JKSYQLDgH7rNo+1xCV4v/SHNYd6HMZbucT4wrYXRfp0FMfOSCyvDaCTi7QAKyk2F2yv7v
ZokCBU5p2BzIP9Cv9V0bQyAdnql2IUDPoxx5rYCDcYbCFWqkSG4LAcpypwBvc49aLqB7OujSK3Tt
sCPBmncmfxrZmxkNBFDXCemgWdza/NE5ZRnQj2kV0RMlqyGDkT3AnrNqXxExYmUIQVzZqExtIz3J
8BdH33Qx4Dwt+YokwqqZTsFHDLqRAEQj1lv91kkwukCPDTI31rtHb50sx3wumMZIPZc5ZZrdclS/
9sup+7LS6+oYMamqJXt0L9SY4uSbMcUtJ0SFf2cpmKnIdWyrIJYf3L6VCTMYLfq1/evYu2pIULDK
zQAHCqiKp0N4Xx3nUUQp9lHeBN8H+/uMzz7b/vRkg1LcbRmkudqBdXUbHSjPtA0ClvJ19r7tIwzD
9h8o45VTXPoebbEHmMpMfcvz1VcXyJ8kjhEBAcy+ZpWBN75Euvnpso4RbJkNxHyJPfBW6LP6bxvE
VCIm0iyZnWrAZ3BdaWlbIc07sPh87bxCvw7M7kiqnnRNRN6DT4BVl3/4eKmvzu8L5pVYxZ6GX+in
OVkNFi7NfUGSe8sqnmBS8qxcHQ1WdXoH6MDSusjcZzzfPuJ4FHkuSodCDzqv4P8B2D8c9sc+FNC7
sxF1R8ow1RjUWMO2FSLPXAgjybrV3lf8t9/9zOG6WD9gv7MG+PcxZXW1yvNS9gIg049Ua57jLD/J
Pt56Y2FBFHfJHF247GcXW6FcooXPjDpfM7Wch1k2AEuik5HCl0Lzlq75XVqfnX1STbH222M3ii0k
7uK9WsTgxjnq9hxvli6qJgZf1DpqWQsnMf+dwCPC1YCJQAjRazN5X7m82FjnXQusD15D94OPDekY
8nVfbCaABW9PKRErshVvWtNrawZD881qtJIMrSL1dBcQrTEUsdHLMro8fZ3hnZ8l1KcK4dFLGaKn
ezIrYDXq+K3FoNUU8xXpCCPm7fOjCET7sAJH1SKUc8usknCdAYhfBLLhOtsyUOSVkq6Gzxbptu31
1XRHdm8MMBN7BylDkfDbdEIxJd1xBgBWPqWX8fyOsQdRVcNq22smnAZI2n5zC2gtG1tjpOEVy91c
hzy0sJat+zIDTZAhxxIeCPtyfALz7EFfWNVJaZY7/FCTovTXVofmzGYdblP08QVoZrJiH6zjYzJE
v7bJBIzuGOwo9ssxERQwLov35jO45gqqjvjxTMB27MSYz3NJNZm4VL1c/Mr237v8YhYWRrHhdZNL
W7+GBDEM7/OH1//iMgvpZD+g0XpyeRnDX/fc8X3+i63xGjhpkuCA5QItXAk4rePN6RYcs2qjZGwG
YCsNzwrW/zvF314h6dDPp5a87/e+JQcS2NeDHJi7ikyb2kJtdD0w9wRZ/3yyPDzuSLppcSZ/70YQ
OVBc2SNcKrxNBtDK/gghpMuEG8GiPcjLDs9LsDe+7+LU1mZyDbegBPZKwXHZiC5htWMAX0e2eEHD
+La3tP0IHlW3sYj3RDZYAmQzT0d5oPMz5QAV59kTXaCG+21RQJtDAxZDlgSsLxJZxM6SYrGbYx2h
4a6vtk7HDp1/TpZWmKU/kC9p55dWk4Fo1bkW/lTaUGXLtWU7AgsA3cftUT1GGE7nztgTtxSm9BK4
5Qer2B/LdIPmvqMhG8KhMECQhfVgCHNNc074hsHh9OboxjAILdxAQ2J6YxKoHzYDxi99zanmaTIg
XDhb2XuwsDgwxVVwWWCMjbySMHZoA9GQqeG7vPJ6nID+XLLH2Zt7WHze1raUs+NIhLiluR3Tnt/S
ra4PdaAdyMIBaKDr5nqIuOsu6k5HadPtueL7A3WPTvy5BRzHNobQFKhtjZ8BdHD2Jet2zXoEI0OJ
M7qRzooXeFoMja87IdT+cnW+uhO6+lDQpreLeV5LzlT/ieuxlC2BEFtz1cPfyBkuMvv1RMtLtlnI
kzUTUhbpJdD2VMFMLxlfbH4+0bNlvASzgrqif0i7c5LmKsCZ8CEDXLwKFlbgJuzz8QZjw4xg74MQ
T5bntEkEwMyU7R7POFQRhPNd8s6PSZm9IZ6cno5RiytaKrxGpNPDlRGs69wDjksjCqfy7MlYgHHR
juICUJ2w6MSawup+BSOKpeyqI9n8fGujpWojGf+mAnchTMI/ZnEXcVlmGVtK0pqz2+EGeMIHhAko
4dcOoIL3qSEJYkoYyHX+Prv2XkqWdI4eOYl0NOpGLOs2I/isSqRTU7SZU/qTk9EHIPV6TpuB6urg
40famRV9w3Zbd1HALl1XNa+z2vhYTW4oxHcdnYdYfGf3oGNbzxijvHr5OTTkTfAf7WKe90QhMyUi
+QWVlawPqP5xtehPNKI6zWf66JjfJWAnGlpn3vBZYeqr6Fyk+TagRS7diJX9k2PTej0R2B0hZ5NP
Tw75UEwRhBM70UrExqUgGUtAntEcXdCxCwDdIcRsoZxyQOMw/rCmrgu++cjOEipN5r7sh4/KpDlC
dQAKUA+8dq20QIeK+wIrwpaJJjKhnvGpBSiZJTPrmX3ZtbMyDk4RtI7ZZXz/FkijPk249Bjzjsi2
Azt32RsJGa40jKISwcckioL8SysDywybN1tYttWqkM1/trybiV+2SX0NJ23w0+f8WzvrQ8kEH9b6
xPevg6PzEzoQfu5ds+DMGb9L5ztHp0RgFT3b29asQrXlrMCay3/NEgozZ6TNXEIDwiZ5UxSgA4jp
8+nH0UrRQksaryogkCkHYwNW1EsIiP7lS0IU8bMKPEExs6G3zU6Cgu2UCoJuFBKJVBoWaNjq2Qr5
WQvpNqkifSbDpUdTn2kAn7PGX2b6+fufuXcRRGIa7vDH+QpqVzJsdFcwxDTJK4kJv9EEjxRH+WKP
Ykb4WjndDvBc+FTxsmdVn/de+31jhXUsR6l4dH+KOvpgxIO7z8Lu+l941YMnshMaqCrZOd6FxRfo
n1lnQbvtyYXl4w2w7THQTBtYoGmKB/1d9tbxNyXSuc3G0mFGZcGxBQHYLdZxIuHC6JjAF/6ZYxkv
cjjH1IVsqrqCu2Po4Q7+pjaPdigqr4yyah+gHaBdAJ9XDOgUx++LDG8hwqQ7hLC/9wzklo8NasFo
Drlk9kqozkp0fdcxuOYpCoSDipbAertaB/gGIho+aFRqdNav814GmzDpSATMN3yLG6SZMHk8ca8t
xVSwf8tDLX5ccP3D4zjaqQo2y0SlXax3sSU7NRZCpojiBdHDeG2QDyqmI+o8Jte/P1d/QhKqdj9W
G41r62HniWnvJHHFxKC7yxbhTyV4J3l9Y5e/VZhbi9wN92hhm8i7kRe0eIBXh506Cf9YsVP9CcwR
9vqfgi59erKyrWwDbWppHM9GURNS2OW/YtZaRDhgEqt8it8VMRloYWMCpdtfRo0LyJy7wgWH3FpO
ar4gogbEf425qlOXhYJmDCjMchep3lKf72neQUclJHgsRYetXjKibt2OfgpWk30cgMk1PB2vJ2hc
SqdDemFYF7ad6rGKWxo3cauo5qwjui3O3UNE04jz8S7ripNMrVWSS+JUQe8OMJ6PeA2w0V6RCpDM
Du/U33VXePce6dWPe9Ojs3f6858RA2UYjtKP6g8xdapzp91mNXUH6olhoV7A0O8udjgt8PlJpGyH
VCOCYTPRW8d0U7VtKCtIJClwV5EVw5SGlMb2NVH8KULKooi8KTWvZg4YRd6LZUX7nIt7a6KHmfUp
AasASvuyoOiDEGoDsa7Zkqn4qqPvyXb0zfZ8pig4EFDadqAAPTqBITPYVycfrO2UfROuN635/VBS
cdcVVkWqpn4eZtS43axDOgm6903NT80xpEmfY2rZO5fHJsonNTQKj5fc3bdpHsuJ/+lDiUEoCNVr
XZbY35aS5DCcQWuNA3XVM+XJOSpMubqQuEd92zZnySYntVWsVIefVyZcS76g2WXMwucI35+KmHbJ
k+Vo/dmbclZklumG/6ENF+MaJCjzW4tb57zcrStSM1QaHHcCVnDXB8Yt3o7swBB9d/abT585jDF3
meHdDMnJ4YqOt9Txa1R4EXRK6pK+/rNF4CNIF2h/KiCq8UCqiKLk6j2Dy68NTQ/gFnEbJh961F6C
FXo8+fqU94x+L7iOaAqpdErGrT26FpqnzVwcTEDiaOzKwdTZZ32JkMiTRGeslHgn9lmce/LCyP40
zR2wRL2k+SNImirlLJMGmEnasYqfbAbsEymappIXZMD7t8UK9JEjhqo9Wi8PIDjXL38rXS0obXOp
qLKDAFgcrnxROVK+W0EqV2TNinOl9fAtjyH2vY7TB+wRDAXXY+pmNdH8N4D72eY6u+AAtvajGrAK
s3hVmGMwW/ufUobgWvzADi9JGvNh8ITinT0u1g3JPoYElsUpJcGpprvz2owWzpZ9PPttM5T3po4F
kwhqCz1YDYDSSguw2nt1HR+8q7XkCfdhBvSzrXg3HdKakJIV96X0SLbH59jwZI3DaYZk/F5mVLUD
d+XLhtIrGqPF5mbdgv6Z8o266/XQP5v33K/IpKzjUAxRNAxiTHytq11NPuefFSmJtPlUzSLs65jU
CuuAh7cTNGZoEwuMEqz/mrZ5SkmE4EL/pwSfttN/rfz4GGQsp4fxw2Ekq2AgBmMBfgI10LDpF+Wa
7tR2xuWz4QJI3zvKUgGOEPJ39vf06fb1B/5+9zBccxz7JYY3C+Y1yDWUeJsWgTMHi6kI72Fx8ufs
ROd66Cr6lA79Q5S4+VVG6PVKRyv0nxy9ndqkKYxeX4KYtahjI73TYMew13dimA5Ik++EZVAdYgHx
Y525jcAfK/lkATO2RgbQ6+KI/Fxs0HfM62AvIZSrEmMotYcE2E32WAVCuumKbXmLEcR50abuDKau
HxnZ1I4bqoIH16swDKAwthxExu/x2yg4iCpzWQxlRep77SVW8JOslsgu8uiSd2UwM/L/BGfdC3Nl
HvihAjOTKn9TRKf6S7JvsfTMFoTXCWvSDZAElbbRVOx0kQ1sjfRK4KU+SZFGBIsrZj0AM4Xaj+fe
jqczcY6+W9PVuyIyHZUnS66aU1zAAEABlNmGQpkEF6t9W4OBdvtEzKFcs1wNQO8a8a3zgJJ2OuGF
OdR9LwC2W2jdC6PZrckHH1MQg4OdXZ83JFw16itPPib9dpa0WA6czL5gjwgJWj+lgO9sZoxvtgCi
0OLtnDF2+vV/hXTMk4cQ+LTGUPdy0J6VXm/Cb/0C++/UhqzFdfOzrAj2edCqVTK8krdkmnthPq2b
xhLyL7suW9k1TXu4KQzfHTISWWDiKGuaWs8IBlyqR1qMfVV5VTvSA0njhzbOYhHWBCOSzFWn1J1l
gFjRWicZG4WujXk9HPsF/3myXwK+7bbpxhq7SbOrV4XnTBqYgFX/K4B/bouNof6xVn8c4eAPwPj3
whnocWCpAFSMfqlAq57+u9ze5xcwwC7qgf2YswZMz9BNYqgbw/r/+BnOX+SahBLD/f45f8DLrrsW
AMANrnmrbdx9wM8BPLVX9cVjKP3IzccMT1u6jZSk47VdCwyzNlg/+PyaKBa6ywZYnATuLiZeiGCc
B1aG4gd1zSMCRIw1CbXEAhFIJtBPdHNsrHR0QWpGqrOJa/vSbttzZpKW2BtGnnN/iskbqtJ2nfOz
LUSsEDH6WOXulD1o30c4YlGVJzdkG2yWyLScUH/wKkgd3IMBQHwdR8A9FichHulZT5k6WZdwSpnP
RjvCjR72NR30URY12gdqvLdvm8hguMoXzH9YJe9zplugZep48zdFMHPcSPy3AA5pmAwWGjV83yPC
7332RHuKOIwkBM6PTHQ7q9DfYqiRWlV77oUCfojAn2LmKMFzBn/+SycJ1zFQu7DM4XptlRdMswSD
XEvzCJfkyI6lHrP6WCzugyNc2u6b2Z65qDHCiB15KerZ30GtRMEHziKKxoM3UuY8pf6gBLhuTX4r
hOThcgAqXoImhEcgjCtw/Pp/aTrq9OP8KK0y/1MLG7nDGRm5Mc64eQzzM16gGA67B7t1hfTXS987
GLYekpqEL2uAN+BP0J9b8my4seSxJcuV7WqLNbrmHo6g8ZLgP/C5yXhxFjtVP8OZ2lwAYbMU4/Xt
vQECkfV0wI6ljt6L+2i/GmQssjiquFSp6oqLlNdBh4p1hd3OxaMo1k5TDe896LKuMHpa0NFL6sLz
tku0yVcihXhBzo9ftWV7THElax0l5r2c4/hh9y3gWc0yZxpXDdNV5LeiOtvORNfDZIUbft+pb0Lq
zZJKVNIrfVGraU4yJ0fxLpU74RtSh6dxLUS3nHp0BeQR2WabZkat4+6nbA0F6754tCzkYdWzkNLQ
kaqjpOvq2nFeYyhhu0xBnHR1SQWkGxjpFS/U+5WyMbzDFjfQb6Zrrd80oWvyAD1s5R1Db1AQSl8W
sFxsnP0UdTbbzVKQtVsqq+al/UAbSXep8+yAij5OF7c3D14jLFQLPBRPv1x0n9oVBZq6mPL2DkEe
hbSMeaT2myxq3miLDZEX6i4DhXRlcwLuu5hjx+sHc/8+lH9mkbzxzsT2Ec3KmjVfRrFRrsJm/I0f
Mg1m15qSBid9FZ3S0/vmYdLKKKN9nvwANsh7XxX9b7gyikWD5z6BJ60aIqmO1wzCP5snOR1VF9mJ
ajzl+Td+FoC2YY9ttFt1gUgZFiHdbyX7AYWl8VwxVtNiPOnB7NxztbBV6D/gThkkX9eLTHuNkOkG
SFz1CQsx3MNYuYgDFIcqFa0/BTfZ91+RinC0aitQCHOTSMFah8Vs8Ht+M+RZIL6QjtDqJuCiSTmf
QyDsGdE48SY6Yhac2zfi8tec5jOdRWJaeC8P/zO3SavYD02eLq2mE8EbkEky6vwZdCNElXN2BxUN
9JedmpC4vzeaL8QMj0H/eqf235fGHtV4zEbcB0fH502L8VTO8NLTz+kxDLIiTE9i8AlYQkAbbli5
1NXfj2UfiwgpAg8TMR3uyOL14MrBBXH3fg5NXJidnI/bCQe1OBQ/rxWaYkuJidEUft1tzNulkw3p
kVI276GSCdA04NRVF+ZQcfAQFhwrpefIMrGGUXuTNySxYWne1vXycRrrQBBWEze/Wcl7i/xemo6j
zN7wRDRr9oppwYoIkICaR4hYJXQLDdabTsJoNZRhxbzTa/lcH6bLThGpsZ/i3f6g45tmqDUBhQIS
F/0d7tEs/N+KNkE3mx9LkiSMpubrjLM6qKOhXHAL7NwF8SCuKiFbrK/hJF6cdKWtr6og4sAW4c68
9++jtudHZEsxkPzZ1RdTF20fmUUI1B0RRTPXsVWZvMhOdchbIocEbYqkU+DdxrHxNsHChoOVx2wG
xApCgZMsN2+a9TtDEvdnkktdM8L37WfbHuTsQLlAKbC4huoOydSPL02+/pOG8b0uu3a7MUoPBAtp
bcu5FqjaRSJHp7Nqu3ipr1y7OkodgA5lNouCkwUSDddTHDnE3ztVW6KUcYkwqVrQR43snbNBIZUi
JFc7wRqbl3GsSe/JzZZmgfWXm9LXzzzTOXEy9nn6PDfu4hROQ9cqOLWpvRuLoYSSadb8YlhfRspA
mbiNKEd9UBrYo3ECM61bSg9+0YI2UwkCP+BRydX+K0AUhQzqzkOfODV8gkl0QlleJkXwV/0c/aoK
zUpEIJnB5yhzksgAZ94bjMnpzVv3MSErsXWd43mQ6ADc1XA6Vjt/+vj/o9XDKlpUDWu6gq7j2DLH
DSkZLxydGNmOrmeyMeYB7dJLM582kBd741dbam+AGey3D4PCjU+FE888JqbTN9aDKq7Wdokv7A05
mV313cic1WjKoue6TbPDuuhPkBO6UTSuAPOlQSWY80Lr3ljZtkfy+WhglQBjNIYoPh4pbg9SpdXb
RT8ng35il08MrBGr+FFonqQWCtXdO2nVZDVurIp63656cVFXnoVYSGhowwoJFB/KLdOBw5++Gidg
c7D0UIIH40sx90mXHJw9NgS4wCoEdeWldhB10q7TYp9vLawMO2ZdSQpzRrPMTR2RlMkuSKzde8bs
B5/YIdwHIHVBt/NMFuzTSPgYzDAP8fQucnia9L0tuGhpmH3/gfbqXwtbRc3hhgN3EcagBKHODT4F
LToZUy7KeMpQHc8Fs0zyT/4+bivLBdghS50Fn4v6RaDzL7vds7W9LFug7h1RTkFIE56OOXFNMJOK
MXAsCrpC73TiCgKGxdFkskPqrKSYJox7GdGYuo0S6O0PYF4kz87LY+lmMMFRrp0hMUYEqXa6Wqyq
E7kUEoZlw/dZpGNd1gtFkJvsAQ1tyyttu9OaULmOB17ikv9BbLUbdvkDk6nvBFlku274cPQgGsIk
Da7bBLSwCPtj/pS3B/mX4FGKicLmPxmV2V5ohvzGzPCbbh3MOxa8CSmiMDL7lnqIoZRC2YYFQuLL
hJHuPnhFS3YCcm+ueTeRzFmUApODeKQSkPZFojb41RwWeWh0WMPF8km6QPMCKFpKnH3fJl7+U3we
fAbZdmvbW/n6HjcvOSyvcAKsMvsbguyiiCehURR6Z9jEtEeA3RcOX1enTiTaISyiGtprqxMBS1r3
w5z3zQA46DBfq3Sdtc/2DKSfaLyGSKX51hG36EvPNOOc0U4tONsuFQT+ciAmPlcVwN77kHYnBgRk
oeDEymTzAs6BnP8NtkJPnJ95qJn4GNvsvWjwyK9VfO7azV6xJQyxOVOUpz4g+7FqNaopY+CecWnd
hc03Sna36DK4D+hsPbnf7Vi6MuKyaEsD6hKDPx4R8rwGKbOWId5sDNN54dwZWMMAWL/fhNlwgCwe
z7LbVkTEBlO37b+l0Dt/bH7OFroNKykCi84t7yEqvXmCM30QO/ut7Wila0FM0rjlxuM6yde05eop
npeM4weq0Vqc8oz5RnCS+ojVT7l/RuXeakKnwrl8AZmO8mrJX6KcqCvOtITF6V3WfKt4QlUDeLBy
cyL4HpXhzSxv+B60h6FNRdm+ZHZT/1ixinvE9tCm0qpUQB+M9btbtF+gK38+9JuffyC5swXVREHr
9gFAFh4W8CQbrqBD1TeMoc1kEj+CVzEiu9fsgTKAVOSsNaiVAw7lmtucSuSdj8CSFU9BSZYar9kN
5nv727lIJkJ6niAzj29GKK9F8tqxQIldHFYH/T/ZXP/V5j6zISPGsTB2t0gyr4RgWeAtwJUOssTH
j5lR0i1xN9/miG07asvem657Uitd92D9tL6XLt8C4QAGOnaTCcODDuQODONg/VQhraNyg+raTimS
Zr5QaQ7n3MJV+tT69J5lL1PVyeEHtkJhXJAs5GxnpUPaSkM0qrW806QJ7sk7HrIdm+15x3DVukZd
n6hKe2yxouWjU0+ly1YJ5MlITT+YrQX/Zzk48GZ1C/jS7GFzaLoeEq7YWDTvM+XkzbtNA+ZjkVjy
wyXfw6hdVP7R57h5mwKzDkL7j+CC5VVhSGCUpQEGItqhis0+Uhk3LypGjdWKIPqHPcZvP08erpEI
JC+zklOgjQrks8yh7SNQxMNZrxOLJOeP92NI1m0m3NvboRwLOYzx+izYRgX0gaxZFJYTlrDInOqQ
qj9qSAetaBz843WE1XpOfaHEKEKCxsmLN8Ptd/FqETKHHjd7ETmAQiq8ABlFcMWP6FjOI1PnrL9F
h6ea47O3y9gffRpyZXizdBUW6lh3eZ9oYIDeG5lKNfgKr/hQFKAh1UnLND/vhLH3s+fWSfge7PdJ
5knjoTeBRhjBT6qJ9TY62+3a+gPErPHWhEH/H0cXYLqs1xHavsTzJ+BkZqq9zgE/LCJUsjHNzZBZ
v83tGkDK9/YhGHlv3g97qN/6LrwVuXh+s21ov1rNwFTUTcFk4yAxFW4pN6kyva7s1Vz1dI4KHHg0
m5RKHTPL07YN+LyCJvk8zlvWS6Yg8PLXzrVeeC9fdY9tM4C/0XkMqOZRsATJf8dsCjNsvYkCrnq+
WiXGy9uX//EWyxuHhSBrpE/VoqQbvjK3aFh2WEmUTOUAhfnF1lp0tgixH0/+4NMf4EwrIUqnYnD7
DeE6KBGnhc0hdQWxE1QKS2crLF84kwDuvwHlvu83NBonXUIGy3jPB0F4I7jV6JjL6PLn4eu3xRgE
nRLeiJKFCQHOgeo0PGtwyLKK6cYWy+RhJEzlBqzW1akCaDlsbPo6qZujO6e2z9pE6xq7eGeE5XUe
z59xRgZhKwrOAPD/fdGVH//wSidB56UPeO6PrOFrfjC5kFjtXBe6sdoyeq+eZYgyJZHonYyv7roe
qTaeFIWEzTBOzDjmy0c/kJdP18ticEAz55YAQgLsQj4BmXorfBcy+JME0g2XUBJyNiFpn0slStWC
uqdHyO0yA6KGzvGOvjHsZsYwVAupVl/lbuL/8TSimszl83GzIhodbZRra0qx2GSLxsUmZCNKuCMa
/89tXpfua+eome0eycbtuE4yTWSXuaH2XuQKOTW4QhEU/j8BC72q72xcy5+G1PuGqvKooFQ747BP
MOta1LMIf+kdUgVir3YkPUMhfjmIst7gfj44qEDytMbqqi2CAIc7ELhz6BiNe48eID4etmixptEb
gzPdptE4IwF6b2T/6aGz/R6spVa4/+gzCaXD9CNnLC5XflmgJlYmJEE+S1Y77qC6faHwsnZfp2q6
N30igP90jlc5l0BTXypbac0zDqRVr7NUbBonb/AFAjn1jU0Vq081j+TDMo9+R+2+A7+5vLYcVaf1
GCX2OfrEc5Jd8B9w3L9bChMrnSjmC2D3KKvpvQ3XWR2/2Z50r8OBYYFwfeVt/bjZqSLKT1708FRl
P+EqDayluAolW1S7xSw3r8dei/NbLjheCt286uZZp6N+YYXPGtMF2jo2ERpov768RA8m1QMXf5pw
g2b7ultLU8WTkU2XkaMjeA29hoBV8/S4FpxOqRgq6Wn6bFUPmZP3evN/8Vg6KuMTQwBrI4IYV4f+
0Y+tdOk2gI4qVPlgciaSKUiTKjqK7tW/ccQNwIYB/M1F7Lg0BbGIt++mMCAnx9Wlk0o4pbYHTwI9
QfBlt2jCXhAyG+mgK9DXZeYflvVAVIZyN//BCiZzGbWhW/xtTDFKjFLX0hQxlHjB7M3S79VyA+14
bttl27SQ/+gvaLp5avfStQrXy2Qpnv/rTExp5BZJXzvjoeHT9G4/olBDz/MxCFOJ0VlcEy2NFWBD
ABcuQHwqAaifnkz7EETOu12wejyMhB8osQUaqumhVdKJ/+K7Nq7rB6u4vzHTKAKqHcn6jh2t9QyJ
w6DJjBOcfd/pZC03ZIMAhPbtZjrrkqRq3w7mE9DmV2VWLYQZ/QtdqGwOsYFFDgacG8I6GGonBjGi
7eE1RgI3oY0I4B4epJuVBzDWAPagXu9QFOR84gtfYrI8ysEZTE0fBlM0qnSDGYaaMYFVaBFEJpE8
sHPjmtct7PdLv2RGa7mhnR75okNeL04JkjUg+v48RGn5YR516BjaT0cz6yI0ozTlFAtZYiEnIXNB
QyjYgBtnBSawEuP418jDl1MwdodgBAAOV0G9Q1qayZaylDkPB9jgyDyCFwPxkk5TA8vD16GLYqse
qXDAhuk3TXmWAZSPQnOsyFDUE+ytlnKNNgWdw7wVqT61fYGfoZuMYUuO+BOEPPGQECmoBtWlx91+
CgWDaqZamVtyXT9yWN9Mgw52bg==
`pragma protect end_protected
