// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Im2zHxZj+weL4ZaQO2vqar7Km/ySJEcWIyI4wz0LrgrGlg/UlJsgVAhiIHOz/yzK
JxbOYpLcdj/UfsuyUqKN8aNbqxkh0ji1IZHZgZyCypeamAdD9v98r0jhfiI/TLX1
8P7Y9seYn8iLJfFdUT6Xvf4LfVs55NDjfBELt49jP6A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8432)
bUw1AFzlitVLVOaqDeL7Jxvb9xAEt85/XeVmOtQgKa3gqr2SF6knNiu5OfruuLpq
4wgZMQgrwVAvHtbtJCiP4dPw6lmXem0whs2Z+MVyv0Ceoi3Ybj1lJywXSVWA1qNl
aJC7kY7gnYnnPkzmwJNEXMnHYEMQX/LFle94JVPb6ulznjmQgaA24D/SiKOA81H+
+C/8wE+MphPK3i0ZalUNaa7C/jNYpfRdlnZ3MLY7ClnhTMWSBs3kHs9ybjsg+1pD
ElG3333NbNRLdvNFG228KsXUV22MPz1hfdKdxRp1fpTXX12BUnqb2bx+k7ARfXtJ
zGblTAtWrC36W8Z6GxNLNQQ2QKicadEGrseCWDHa8LyA3JncqMMRuLHcd/3oYVTP
xFAG2dfDuFpmGwDhe9abwkdaf7xgCwgrftrUtwc7Ue/muxtuI/F2934Qvh9HelHa
BBFK6sdzjoJad+YTTNzIuKmkqZAtTcizQHB9d24pQcmsvOKxWZ+JjYnnK9xsqS+K
NLR5pqvz7NEbnJ8mio91+6kopnzwGqnp++rQjWtEcpNrXaRhxcXbwe8CfAEDaUTP
8hR4Kyj/pOyYichWj5JZD2d8BlYXrpXqrTHwHby+bT1kEjZlMHvvtzdY8rlWyhST
kytPAuOjrOgmndpJEk1DjjkPwIVJhIagjHW6qKOtCAbBkfAyh03efT7z3uF5CfUU
U+pO6Z4S2hyBhm49OywFC2Ff58HYlTtmi2PXpExhypNLwjylfW131Z2tvFIBRYIc
B3AC5v63+8xRqSaGsvzsGr06HHJSlMCLVp39AZC5JKThQd7rdJhObWC4C7MCEgha
2OzH4b7FyOo/ziaGJPLB9Q/4CJO2tPEAK+huPhwxKpilBhvv2s6T+RpBRDAqtJGd
Dqt/N0Qiyb0R6sabyrol1scrSgkRzctxtZzdHvnhm10QCF7VmjKoPJTiyhYKsf63
8GM+e1XThXG1rkiUl3VRNEispB/H9JpFuyb5ivr/O0io1pofxS8NVfbCpyMyyBqS
eFHiDP1F1tZwrz4xjk/n78+4XXd/6ch/TJYiLbKIWH+yQc6ZkNfTPfzLkXDiKX+Y
IlceYgL0pt4mcclVavozHwPD9rEh62F1egB6fUk3rR53rnw2yBqtaQB/y8wL1C+J
GeHwVDD1pcswqU/MJDrwIT3p9Gz4KilcZAsYPV8XN2V479kUorrsV/+YF0rhU93S
OZ6evL9pEdPeyBc+ODZaSLmrE8lIG9xF9AGCOAhCWpFZ9fB8mGyaPHqncr1ugJ1P
F0b5T1D1+YIESpAzredSmpEY20fKb7LsHFUdfEKdm3/OfyYU6pzVngcYV6c0cT20
bfaZnS1DBpHsdOsISGkJjglwKwBfqFgwWA3TywEPr9JPlD43bYO3KnqTTo2LIFKg
24yDGYpndISQU+t8KKknLp8+n1KMxHi7Y3wV+9oxGxSSXDHuzbsO5m4ejk8y7E4b
x3uBEEF7Ff3IFv3s9xu/Z99GEbeGVdQXXHCVr1gNLATo1AuDX7TTwIKIGR4pz1Iq
6hHqsgd63DGpypvaDSzVz4M9fxYycKGNNTama2bdwAoLD6evnSap1cBg+fkqmmVJ
gmLuIdj22vsTph8XNq8pBYXw4mfYXEpSBUdbKCsFFvVYPcHciD1jItM8fWyzoS9R
w9JdV9MyUv1MAcolF3kSXn8ncNTxpK+Bke9tED3B3cugUusJzZBWFnydRXaFAQzZ
JuJYY0tNVIkU8kRR9Ia8MTn3f4islwBwSUArPSYTL6PCtnoYlkeew3faWjImOrsW
0OsWW7YIto6+ETu8pVt+AiFYGzLUFxgdjn/BzIMYSVHsuCVjR99/ee7CTA7ioZpi
oCudUwkLKRtMKrffHZFaEJn9+zoabBPLxeD6qAgauL562QVgUxjlnEWGPMVO+gjc
LU2nWzIr6JQnZ+BbjWi2AZ+YNeBCqiWoK+/2N30IhMzjqJupvfzb9Y7GOxhjeVCY
hRXM/HpHFSLZLgrMoa7h991LZJAgGcgE4iWt5l42mwXPCUixJ7UyDmGej95Mdv0t
em/IGjHirrsezY8X3/g3oZY+4SyX3Sn12cL6E8wtZrMLpDEnwcGxEtK4ZL/2hz2N
U4EVNfHRDGJwMY1ER4wOxuDRiR8IBhrh2CuCAp8dxkkrRaT4Xn+sikAzTlZIB0it
dKYs3w43k/4OTdxiusHCPttDyIYgyq427iA+nzPM5VZYYOuSI2Yw6UkzP+xE44PC
vD+LgDcMCa28/vswB1Nl6Bz+1SgvANw8n4IymQKsaEXPDj5o0NdE/Cnu7Z2EY20B
zdpPEUPUU55LjclibInX1rroEX6VTEtyQjWxfGwWytG2gjwy5mWcaRYX35Q4FK6f
BwnFWk1SGMlImHUkB66ZtCARmf2Lz6w/AkLm5A1ASTM7qKyQza7JiBojF750HI1j
a7/GOfhgI/iTCBOrVNcyaRJShLkHY8sQjDYQTglYrR7cSjvLQ5M4oQvn1qqRBWWl
EM971yk172yiuMg0LDLq0uXooK/WjFVoegwVRiQPS5Fpy78b9opRB+blsUhREuub
k8pEaC1C7+N6AmqCzyto2EjnePAKX8aGx3DUC2JGWtnas+esLRumlJGF2VB5GT+C
tiahYohb8yNG0jTxpNeuLyoxaMcnIuYkV0wyKwvRR4oKfITuvctAG7tJ4m6QZ0O3
Wcu+z6w3hdPW+x0+Vs87fFzmOSksWXeHgcYZ2RrP3JdiZ483OOxmn1dvpuzVFtD+
GDt8pgtvzcOg+9YsxGThZHEVFQNiSbNshExr8NmCPve3czb0FPWhuCcGBjweYQhK
XYhabZIm+dCx/zlvgm6de9fNQ/FYWDwQTHiFjvKW/5mYxJsSTOH6tR9fec0I/9gx
p6egcjUUj6bwPgBBCQjaw+3YhM6Ljq/HH2sx31OIwhWcICxfCoukOizasUAeKwAC
1Kx0Nc0oudyU4nTmSoP9HntAeRI6Mgk6PJQ9BqcG1Lq//YpWJCLMWPlWx667xTAW
e52gbtKPjC2dFtUhxmTo1MCJonSj1oMC7NMPLxNa6KzQ4IWW2w8zoOfo2ckBTmKM
pBW/p3vm9QeYMZv4lU0bymhtfsS7BI6fu2NjFgLd2W8bvagW84ukSw3uyS/ryqe2
hP1MfFzOF+mtqWta8p50UP24sLVV2EFKGhCvTvtOyOpeUeRuIAaHCl0+xEqzJP5y
Bh/wuD9eOQsX0sn5JmBWRFCyRWny5YYwDOwvWFn7EnbvoQlYkZtUux5MBDvJpp5X
kwob8LHpS7sPO5FBxyFbwGbzZTzfTAxXQgsRlMqQOEW3467Qx9FwxIyZfrU01LE/
I9NwyggoxP8b74sngakJi/qgyDXG5iuQsVe1atJFQxJ+rRI41FakrmshB7aINERK
va8rd1aRQPIEBJOmd0f36gclvo2OiNZLl27cy3aw+cHmwZCmV869ybrsr67NyayI
LaBL0/L72QZfmNp16e2rqhsKfR1B5luZi2rVuGiJiGqYQg1xYgnk0XCVFx00iz9D
QbTdlyJFnYoKWsMNFbLB7naZhxXHC7yEvknh2iKWwnIKBdBi53u1/XZ0UHfkznbj
JP+17bADXLEU+f6zh9j22Z1QLOUb3/EiQ5H3D08202UMn5F7g2mzsSe1jA6+8IMh
oTQlAsgC8AmevigFMjfRjgTVyn5ztCMaKRncVCaqYXOiUYqlGMQK3S9Db8jriVMw
mty2QQEnOx2HQ64d8B3i/wLjhDsUwzEZOnqjtzu+XsfiTWiRX/+58+bPA0Dxc459
LFETLyhsPkuAUOUyPzyI8cXg8lXI4YPS5X5OQzQN9e4V7foA8mzC83ZJ/vCy894l
jlYXYKBxuVSkwlOCFjtN/mGdTQPEsmA/dNbvQdJ7naAAhmpnJPTiGt7OwZd9LuFi
4xskV+tlciq7Zdrwq8AeAAjRGsx1WijzYhm+e/hc00AVX56mc6VtNfGV8uY8XLJY
croDPVJ9ZCX7ME0T+PrJEjmlH9iZHUvfiutEy0RTB+kVNu1py51WeSzt6BzLjoP/
UOd4cZ0On9ObgmbetEwkWsSOl5VhEiX2WNhWvoSvEZIXO9dnF/rrgoNpTxYjIhAG
H0qe7kHFAN/q3Qw/tvSARDUGPsyo7hUAbSOBT+rNxLtnd+gmOdy/q9uBjz+acMGs
B2Xgcl+e8X6J/mwSOO96cXM3+ARoMrtOh90/M+nIOTA2z67NoVw08lRoPEvTRp6Q
H/KCsqq/peYQMohdoewGiWw4L4CzHo0bi6Av92mYK2sYOSXPoUJpDCySg0x8dLvE
WZ9MwFPNC3oylIcG1QSkC0k3EGhcPcUOItouizRHboAlIZFOMr9B2jH+S6zCXAP1
eGFsqlogn99velF1kM0VeFpnl0kllm+ewH6ksRGInnHZfmaE++sdQaGUh3cEe3bL
EVTkHkTXkeC3e3K4b188/wTO3dvK8IN41T3KPHSh+DzEVD5P0mmdzRgACJlV5lBx
cx3mHqHZ1DWYh7FD1viXAtha/JeVC53pzECzwg0DMsh1iXP0yHuki9eE/BD2VunZ
wI8Ij7l1x471KB97HmkbsvPqfc+mod26WSgrIf6su+c//4oQ+hSofI3IMkRQp8/2
z4nFHJigUgbuQhjZUR7LUskDjEKhorbsSMYRvw500KSHMXBnz8U8bmVF71pH1v92
ML4q36KBSijHcqp/044/GRc+iwfSzhfafAlJ3+O39Lo7DURp7tx8xz28ncEaQZWT
nfL026DM8Gd2yTZ2tex+IGVfqHs3zLQqpsDFDcLhg0uo4F88BRrgkbiuPrr4/syP
HyN1pCldQ+NvJAu4/4C8fHTbjwslL/ZJ59K+d8jLttAw7QXEwqOpDWNTsLxMzjXU
v2rH+SKz7Wn2nFDv0AcX/tcu7JCxHfy5REHDX6jPazx3DswzPVjv2I0xuvxQX2MK
7+3ouMKOpGwSmGL2nBn/bLmdavVXJ9il6Lj6I9O1ecLOZplOOsstXLt8Z1+KZKjF
CBjcUHM+7aZfCODxFfpigfpI+3a4vf4I30Zj1yEjMr9LMpWE/Dg59RWxOUPH8seZ
OfbhWNnIXGN4tUAuajhS810mffnXnRKIq7ushpvHEIA0WE9e8EoxQvsvL/No1HP7
1KpLTf8yGFnhdeDKA5jexF073Eh01r55oILR2pKHhqn3cPtOnloh4VLArZ6m7nDn
ZvnHXWyvtvdGfa++BcQxfDJUK8onGhevExRYcawaVq1fvi+4Tv11ysmO5zYSax91
Cpl47X+TdQ4WE94daUr3RTbRROhz6OT4lm2Vm5VnOgEHE5qAuN1Z+OfGBgP8ycPP
3OVSH8dA9cqgx9kDgng3HpxkmKWYXp65BQ2wXQCLzd3yjClwg53hBN9f+xHTKuHy
iAYTdOs3Vj15ReDfMOTk7ZXl/iaxtJuvKdaRHi+Lt7OuhtUEWQiLIeYnMUpQ4G59
yu/50xneCoQ1PsyHtWp0xqQxuR2h+nXN5v6JG95Wvr2Ewd41H7lBULeuFZXX4hA6
w2ghffaiPSBwDwFx2fU76qwDjYcRd4xD8m94/5ewmDYRP1fGyothp8uHoZojK38b
fqhpp5JKMeGo8PjJGKigIXOTmsgdZzrlecQ9Cw1OKRC5E8kICRR88b0oEWHLtjDG
JNwiWOJRQZ/xT5pOdAGzVDOhjAG2IlL7SLy1bAX4+JS4pVvEWOF5h3ht1WXfb26X
hOW4/vGK9bm+iGFjLhIji6Yac2LYw9Im7YnUxc9XTAdiZvHsqv8uOmKlaAizmyvg
YW9iQphn8t8iePjiroEgf5BV36VtF8DIVavMqOTJETLC/IGcaSAqzhJdbFQUqsUd
6gutmXLmrH3gfKy3lcLoo8SVNgKYuxnY++0Uvn11sAPZoBdwOyV6dwJH8MMJ0q4H
kP4zlrmfVwfHuG83zP7aEw7QyJs4chV6fenuko4jR7Q+K1Q7AhVfyc/6v7Gdrwk7
x9TDeIlR7Dj6fHs7DEiPM8t5EKGlDVWvbm0Fe1Fb44Tlk+Z6JuXh6xqBQ12dJj7/
kjbWew7N1zinz0uJV4t9xuNCqtXkucF05CJDKtAgAGtGsjp29A+Coy6bpHgXwWip
bV3DxyZoN1zE+Cs6OADCqp67m00PPIA4otCKvhDMbdBhD3hfAuUqYHbD6+qkruX6
WDCkkIrAgALv6+gbtBrrziM7+zaEkyH/JE9qwqCZB0k+UTnfvtuzxotKOv4PObhc
QyDJL4G4VjPK5XuXiiYW/Ubqmjo0nXx/Yd/xCdLQoXvgKmh5ERQguiZe9Y/WKOSk
9Qx2tPymah50BeFilJknoEf8ktTuKHago2OG/gOP00n5NbqW76miA+f4cuVBqdiH
ahz4aBQmR7GjMOx5+qlbWKMnV3f3mQz+KH8vvNDWwXKyLVwcihMTYkn0C15a1rFR
gts8Ddkvu1TDiW7oEhrIdQ4itkiT0LdEiyhXmmnmdOdYIe57m39wpbbWyFR6wu4d
pxG3RcRSzmwEPCycFXocBx5DZ4+6+9rQbrODu2f5EqLMtuNsbU7LgnKu6WPJhzzi
FrLjMWA/bwQYvM/i5H/ZYVQI1WTt1ERkqv/8Xc/JpLrFKEmvEvJlA1YYTJYfYiAO
CuKwNc3y9LUdI2VfiA5U4XJblsME+p5gipIHquPQPBGhsWbp19rGasj7ipYznZEH
vadxO9g+rrJFWuvwjk2yjFrSBh00VfSY9MdvOZ7FwceoXn/IHakLgcjtxYvhSv9E
A3qMRqQKGshv0IWkIqAJO2ZuCPrwPnRpvmSsAAeCylGgBc4c1WuanwfCEAOcWAO3
NZNkXpK0KuYQLE6XhB9Toy16OJCalV+Eu0vb4N0Onu4LFgoO/kC9WBLZWTGSn5id
mNE/WsIaOS4JdqH4hCvsTXGe1Y6r5eh4mxklx6M3c1V9QqHKtjvKUX7nSAh7i2zt
FaPVYiu06UmNimB8dx3I7eu0W+L5bEIRunRFSFoI7jDLaVr+NjZYwNjm1Jywdroj
cK4F60pxqJYgPz+7bJEczB9Dm8P9SQBtDF8T7550jc83ecwdTmJABGds3l1ZiosD
FhEOJ/f7D+fbBRo1+M1fSnQbIlWjxZjeVgIsMQvnZ8kiFV1u6fvKOAgr8MsHvGS1
UA8YS+I2eaE3R+rqPuVUEHHTSLRQe8ATYxIDhLtKthx8NcrQMBFfm9NTVEwSLyVD
l8ZzdcISbtyx9Mr9AjruDZHwCEQTt6tcgBfaBL1onZsbRWKZ3g6L95MGKBXX+1p6
VBzc679hmDdJXJApVL1+rwL3gpCebwM6AG2wY4BpXKw0KvDTx7leBbxIJw6/Vw5E
7z90GylM8W9ODKrkDi6r6HZLH9HqbLQ55pCBxhKnx8vZoC2sPs8edt0EM6hrJIvY
qw/NceNH6gN0115cSQnWAnYSBww/uwBPilna9ZrAsBOZ+aL+hAlLhQaWoWulLz29
xBcACDqWmoDZhRhBAeSRa2T9vP9fPQAbRGL72B9jyAbx/B63UGHOkB14ZpNEklJ7
3XbxH57gtZhaNdXqMoixKW1Z+V1Pf15jj5vpY422g7me5tbYjRmnAGa8nu9/2gaz
mZxBGWAa7nDNvnyenpoRXjKa1IUsamXW4kB5MX4HP5gnxxKI6VP0VtyQXMw8P1yw
UinDnPYMcvWPI7bt++lGzAcTpHP7UiGQtnbRjGqVN59zj9P3DFZNtQQX18lmnZK1
3CStmCXGKsp2jqwVlKIlX654dyef9tsMpEfFXkcq9LJkjaMW8btTC5HX5galL1q5
+puXw0tCqKApZBMJkV7XUbdtRcC/w4nEvEYJ8KGaWHes0+cB+JNYD3Q6g2jEpzHs
ye8pZhKXh4L8Yoyzhl8O1g0wQNjxgF1zQrCcvCC8h8DCgUAwiCghdyOEwOV9UcWB
1YnlqgXRjMD8cb5MikMAbCftYDa28NZTTRmW49VydWNBOM2eI/T2682OcEQy0yBl
S2ltAPp8RB+N3CQnSxvomriwj+80o3yHyuXmc2Y5BgIy/hzjHIElmbNmZMI3ElMv
pbnbxIK4bA4Jt3USA3R/u+EBe9FlmkrHo75/oigF9KP/qawNyM0WzTn+EY7ZQrAP
5Z7AG+Xj1pv+BaZIwdMA/226qrJqLk37aQqVxuYBH0FJipvL5vlLl5URF1NY9oCh
qCdy1xVSqOJKDwW/U/fjZ/Ib4y2QpGTl+IluEaLJwGFXDhC27bNzNM+oScqIOKYO
7CzGlL0pb4oGcP5kdrKJqxV1YJam/KYy80pG16u2uK8N37oADb8R1qgIM+EI0Hjf
7Po8uXXcSFu8JiCxdTtGsqQ/MOryWUupVzn3fv/MckgaW9LfzamnKCcFwqx1Xq0A
YAm7bWUoEc2s3/U1eXfYRkPUDZCtjGOPpKZlZ0dHmIuPk2EUtKNXhaYfiWdzvMG1
m0NeWUGIG06X7fkfRoJV+vt8RfqV4JByLr2d9e/eirtfYyBqRxdT5Y3HH1hDqOno
AvxTOxMqaKNfASbkdrzR/038pCW/0M0P9DkU7lbsZvUxwOOWvbKqxyzz9Ffo93TD
jPY8NnkP+zoXXitOQ/N4LTefjxJ+Y7kC3RDQbB7dnSHBPunUt+uze8yRov3bjGPv
VrduIDqhKX9T+qEGHn0l7tZxG9gSYHvyK8NEMHbiPAuxjgWUSd4aDrx8/k5Sgt3+
raJ31dN0UDfbXKWsqya5D3cQ82HOxjY1clSneckY0IQh0wHDsALoJT+uCQfgWrX1
wXS2yArj3betVN++we1yF+10lTmneLjTpRMtLF7SQnGfLEiYhU6E2sNI91aJvmNz
qpmKII/p49APyneDNyHvN6fs9Ehx5qv1Yr9FOk8b9MLCTWny/sAffuhFmp7o1q76
DZ7JXfKmVY4qhaV5EEe3mCalEsMo1jOQhd887OfqQgT/Gt5GecxFlnl/MCkwm/XW
RX2Pf1LqMzJEkdED8SY4AJ2FfPjvis4/8e18qB7RWAwn7m6FIKH5q1Jdd+ksKu8X
sv3iro8cayJqH5Bc1zuU8n3R5zhMvFwak/QRQkTqPsNNE/M6hO2T7DDVT04X3f9Z
IVlh0J0cCfmdLHmUpmBbfWj/aZM3BqGFI0Mw5IUN4K5L4Lwm8g1RrJ2ZYcI0jYFW
CrdRPJxc9bS3EqYdcfnHK7tJ52cHO/9mLi8UnsSzcbXyLXIXCgE7puo1FLWRI0mL
/PcbVtGEddd/HFnAp+hjiyG0YVIOoE1XyQrs1s9hdJy7CPwCE+Q62i1YnOviIM1U
hxXwBtBGj50Q1CJligh7MDFa+Tk5fhReQsoki6Tv7Pika7JDNaz+H+VW3iJwOHns
uhSJ1G6tb0ULjpwei6pOuQBK7ZfFbyd1GwwTd5uh6OyRXsmR3rvw/1lkmQImhbWk
qPv85doGDtTp88j/TJLJzpzBFjPf6d25GnYFIkie0gg4zBzkWMoynTitKjiD/J9p
CkLJSjsxDX0Lri0pxlPLbvPDC8jbIhA7r1uiSPA8uLyFSwTfdspaHH/75CQLNKqd
ld5m9GTrGp1O0Ofh95KRgo5r+Xlii/ltDdzpX+1hdXiFNxMq/ybMK/T8eE6BM3J+
GbvG4AqCZud8hKY8iCkvggMrVa9Fm7+WsY8Hc5zfhQuln3VQG5j5HpuzSB4hozVe
COOXjN7ZXq2iCGDWvCoItht/5SlsOpT/tROQMPqrsK720eTPNhE7qP+UvE8UxDdH
WNxicxttGOoTkp8QGqRqSkkRQS5i7W1hr3SJ8HMiImpYXIi5gq7AxP8P/IReufTD
NLqpnxGWxs1COrc56guP8dg7GxI3EnH0kkTnhPRMh4uEqK4END2bO9MbW5ajk8W1
XA2Y703bepMN4Eq2ZcN3K5e/vPBq9wVzXFgYLjKaHx5DNo4TMGj+C48MAAvnd3D9
TE7giQFLPolc4Au6KwcuFO8OfiMwV8o5H1DyjzKhapkJ/VaAJoUAQ4vLEnQtheMD
mbRQ5zeymA/lBdWdAqgfQsYyn+AdQqNHhNfhsG3Mzqt+sy14zQZrRdlWMgmznNVF
F0aLpWdGGcF6lUfHgfRqOmnUtWKcqgf5fTIFqPNx3z0Y6C+GqqwteRRURTCqLOvH
Iq/dsV6US5O2tBqEowwjuRwuGlwQuqBKrOi65aMlE4XwjfsDG3AJehkzjWJPwQOx
hFjoqt54T2qX/7aM5oeWJWKDRMugd6Rxxqw+vgFCLMXKfQn+DHim13LTaCLkuSL6
ZmHtrFDHixJR6WZr4JePNE53CVmVqG8B3Vz/JJM6RrBCTHm4kjIu+gZrlxvnb80Q
oxbkyY8PMKN7k94fE0zPbbZvzVF10Ahs6gTkNqweJfNMwCJ7Mkw8ATqOtPKT0jSF
QY+y4VG8zn3jY8ug0M1o12BaJiHu4d3U1UIh8HTxl+YScACsFRP3bHq41AgsbV3x
Axeu+piYQFTElnMdsLNCJWKW01zIY0BZEAhURMEJqb7aEc8cgO9fiCbtWoThIQO0
92dz/tVoSSiH8Con4SkGovc/L7G8gdsQuaA2Y+n6mnjEC8ZAjnFmgN72Z0nUPTQs
EKd2GvrsGjJqnxzWHjlndl2UBC6EZAbipEQVIkHW4A49bgYNpqwNGaJVFxPe+Umr
jtgYPS+q9Erzr7VHxxGR/pXjpOJaHgtsUddlffzf+noD8PEp/ly0aPdv8/i/CIjV
vRCDQ2/LDesvTdhgF1h7iMqgZhQGkXwhGioiVpar7+Z4aeUpo60/0WfY9T7FgO2f
SeFKAQn5nqCeUN/mPfKTy8Uj6rwO9CKXC1oVAfVeEUTqbh6tGHVaWz6zXq3L4cAq
+5glk7l1lkol6/VJCdqJigGCw87UAbpID5/z1yYPjY24O7CpcxLdhRct7snTjtAq
/uRirKrLxkp5XCPEbbzzPGsLlOOgrym1vxDfQVXad2UlfZzGue526/KF1chDtUJL
mVAebxCosBLDc0FEzS2Jxvn/AxrDw8zFHpA/jAUVOyJCsgN/hKg+8bGGfzHGFYA3
AuV7AWIsfj3SK8h3NWFxzuugl7RG/0n0si6sSd4thlJnTghT3/164EgYQpLcfPHp
89CuOhw0MxbuVeMid3IEyoh4Xnte7F/6ufVLk6W0DzYscXRBEYe9aqlQmgxEsK6k
Kykaip50rvKxhhfUntR/Z5XVh7/Dxng8vyaY+q6CH3jfZe/qw0EHz/OAW5YKxoF2
TNt5E7Tvgi9SFdCN3Nq6PBzLaPfQnuA25Nfa39DWPCBlh6SwPoCL2J3ztqLu9dlk
OuylYbAHeC2yc129H/znM+OpyQvk4DzxeWSOV+FWR9M=
`pragma protect end_protected
