// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gLLx+BW1T73TdvV6TpSEY60ojzGr+miMdt9HTEh3zLPy4/HGVxlAw6SbjrndKYa/
u179d27uNmh4Y3ArAbvpG/ikPKtgKGUQLk5FPEbtgV6XSftM6LoVviXv1/YVOXD2
S+Chjl7YhUNb8UWp5QVTot1QPnoPAlUCxSczLlEUhdE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23120)
emlovjdsCuzCM6gcF3sF72SCfBdQdtBvm97+jPBR2sbR0G2lVRhBhBFaa4DI4G1D
4xisBf1n/pqe8wklRnpXZaAs6/LWIpn7qwWiy10TJ0/oyiYtnzuwwgHwbR1/npOB
QCdbRpmMhqCSfhd/rgMBE9Zf0ZDVnvl+10pAzbpcJT+lbEiys6DC4o3fejLjy4kT
VyjOfryNE3ARLilEz5I9RIyaxFEx6Sb7agVctIPLHtTEPaOCgunUOXAaTaS+YoSE
UsQwka+NFJGYFRPM1eTQNQbQBJ0MBDVfO0XyQe3WcB17TjLZObbogIUW3y7E8N6/
6MxJ7J+ZTC7YNQCYm1eH2UcoJJ+Dj30sHptoBv4BhL3nM+Vse6FPtqSnXulSluiP
CCIg+kfTSnx8aakG4R01CkMl3wth1guKYVquKmo0xiyG29uMzVTGkvXIOl+eN4gH
X5HIMyFSAvfOuRdDRfo/J7rx33gz+JPQ+A2eU3sWifR8oxmprGSqt/wIOTTLm+bb
Z4GUszrW93eny2ydWYLaAJk/ChJEVxKVZhMWp0wdKs4BpIVhV2NwGlZKiiJ9rJBU
j92qKl5NodDXZPQ9cnidlw+u0uOD9+JPbwBLs8uVNm1llZUwBLGhQu4LSS8BGLKN
t6xHI8WyQXMsA6UTTfOFKJ639xljrf7EmhxZl4xHUlIqO9GNd6VKaiTVqOsbv7zV
CIix8B2VBJRO1Lb4HUT9W/eDp0yNCESREg98SHudbuHDtiqAtLmHEAdHoAJokAuy
0H4PcK8ZO3LAckIzZiS5NXTpGUQ6HKcCEPxqvBwHrYbfzwkGC+kwKC8Sdo38PQav
Y3iWLyhW4wD925OfbccbG6T7xIl8Ka7YOgd/XXg1a+DGOSPh6uAa21n2ibx/fWG5
XMBdWOtKR2GYNTdN0vMzqS/9xOzdczjQz19oa1rx6UcssKSBMaWGMK9GQP1Uhr4Z
mwNwu3Jlo/qkZhSexcMSh+SxoBtdGknJhszBlqn/EHtkl+R939fPH15kvA54aNLy
mjF5rdwS2CzNZ77JB1QNzu3sAHqBP1V7jc2iosaFQpMzLJh/ZBIbw9btJvZjh3EO
gnJnYfgfd3e8yRUHCKsuz7Z1eAjJtINh4NB7vjkIhssICO/OcK5UHvoO+eU/U3LI
A7AZwbux60o+Ea3uKwKFO6/oUHytihfLSPsaLdmOZR6cQH0oceYdISvsr18RtHvo
3K3f2wxPudwpcOa+TKQeNsbZMT2nHWMh1ak0cBbjnBcrjzcj61LIYiWEnn/sF1g9
ojgWOsyTqtqu4nlYHNV7Nhfdjy7rtvM1yfOD1zldpmqyHOnw8xo21tLgSlhGNlaR
qD7TCHpiq7PucvkGJTwmZVSzPO4z+PaEkowYOeFAugFJHIaRmgKBkTbB6jrlhQ9G
U7yiOG00mHeS2Ek4UdIO7J2+ER49cn32/X84DXNqqVIIOH1YKoLO6dgemu+AzhVr
P9iRpqW6LIenHMPxApd8d/JH7R2SyDU5wDbctW9+DYjgv8SfQkNidAoAj6tgUuaq
OugcIJutXN+TOSIoG/5OTB76Ggc11RjzbsqsiKGVS8Z42eUNytBiIHQE6T4nccPQ
xwZuugZinszZgoQtP2xkmZsOIMUaPJFLCT80zYHfM/M8wVkQCdVXpXavmnohHxow
8ydTC8Z1jkw4xqIciEORAWPEQgKO0YEj+tDmaiuxfUEO3DECqEEjMU5NPMMxHJHC
AWI+IqBzBS2Gh7UKZOHrApUT+vF8Rb8np4oiSDTJ6V7hQdagRZb/T8zy5tYILMZJ
AmnqNyRNFM3H7pwyfq2u0LtvN1eCv7baaTTUTOZ5dWxmcsYEpv1oYDNuBwmk1539
ybmPt1zEOhyaIj8+ynm5D+6YZm7UT7kNys//33QLpdOT0EZ6+YC7fId0dcAEULF3
pI9f9R+QIR6N2LEsMge7VWKrJMybm9r9COQ4e1vuHul7AB+I2MQfMQwRktZfVEkH
lete1TAeJbW2SdCTjror24PX8xbCcdB+7ANjJVEA9eEqXedMJ3gTc3gjqKh7GdWe
P9ggrrvtMPr8VcOC1tNKlOkjOvCh9B3BdKD5EcnlLCYhNrfKAMOgRKdHea4XzPml
tMOQ0luWI6IphCVGvmtI4VQ9iGBwunmPObaR0c96RCwJ72GUc/wNxRF7QRGnij+o
SdspJl7szrvDLAp1QHgOaVbWgw+0np3wOk2v+QHXuvF5Zuc5j6sFnGhBE4XyS0Y1
kyPiTRMDrdtefQ8DLrPTQxSicif+gTWLhTG6xzvcyrEsRuyeWFjCGWXm4G23LNIY
CGeNU0mQdx09uuIHbIZ0H8/NsCBmrVhUEBYutUbY4EvDLQuU+I0JAKFWPAQyibUF
S4TzgU+Dox58Y9tCTrCTCywrjNFkKopyi1aDV3WdSbWpCwq7rwMJFBGIKou/KZdX
rk+nM2cA4sCSFisxa64Qf/J9J06mjH78aI922/f4eGRwP3n8tRRuG3rMzhkanv6L
Z76cARDLN1wTgG0Lht6ExbZVjFUgZMrTg/kKmfekL1cirObzCRIS/snWM01SwdMj
Ndwo68tP9yIxKwFROFgGawuzWHygr+zF/TG6B4GWliPP89LUnnop16SRTu5u2Mu8
VAQcfAdpsqhaAS66Hq8JvO9PNIcl2nn93hExZISLKKfGOb9DCRUjudP+aZzSq/Pk
OC2Z66vqWBlb0h4ipkfioNiLXQ3UEpOiUaEYmCu/8NVmzkie4jbJYgUE+7Xim+PI
UYO1AXm5/Pe77nVixKKGeuCI3Hh7vVgq0hya4E55LQK3qI/4Wl6XnUYA9kA0palV
reURwLTDg4G7rtnjKHn3tqW4hj7TahH+qmENwgfuxSndYPxA0Ga0TTHZgSyq1tN+
77mr9gI0uZNvvZGuAnSpYWWVv71DLO++jm4nkciOb87WgMB5zlSjbiX29XqAeUhO
PngteXk5W7v+eIBiSjx9NbfMvSRZQL3YAhfa4H9oM1QmMSXUOBqJldhFTbx9AlVC
LZ5fXmdgel+TguI4ADEZEk2N4v0CkewnrDDwaoQOFh61vzMZbVFjdCA0Cab39MwU
S+/VM9J5ikmqJhVfKs92XpS0Q+NWYOVtBJrmshdQX+HSMB8wb75yTpS+UTK7kauz
agpQhq2rO1zxDqHv5fidWK3kWdo2oC6EfbRcWli6XdpPp0HumqTnCs+MSLxqjB6O
O64kMOd3iIWWRK2TASJOW54LQNU/T6WlKE4TWfaBsAhSVAAFFmHl25+vJcIaeIqB
WlMTUa5UWOnCxGtbC3bekI7T9OzL5GE3MA9+7art6PsuSLuteq4y/VntXvMWCGHS
iaJIyNHRWVq8xsVn+ow2PwLUw9MeMZz2uI3/9943j851qBv6cZbb7MfrL9O/l65c
yDBfH2D2zZZ29x7FUepgLNS5qGm7YASvRT9qVhLQJG6XNS9PlegqGvwPk3lL0uXb
LTwZEmVEmBI48x/xzISsUGWjKDsQ+NSqI02846WC40e4LNXYdUN+pccEVbVsL4y7
fGxDIlU8gwcUFwNb8mBtdIZjnVg+xw61A4e37XRcCEEnr7uHvUezlfyUf4jL7Ae0
RcKNSt4/OrtQKT2bJ25b/2xytGwL44430IgvQIPk8GU2XuQxfzKiPFZ0fVE8ITHP
m46Ocai83wolsCfQm9joc507+dfKWxY70R4ym1XBPynQ6LZCabjgr8viwgT8p+KV
X7iYXDns5U76M3kZTiAGTcUzVCTVDLH+YDR1jfcW84GqueBo+vJc5iYfpbywJeR9
ChTaVof5js/tHWkYEQUIEeT0/3V0Nr8AaVEWU6PQ8LDOvJmmuIFNCEZqJrg8i0IF
PI6KGAyoP7Ti86zpWeV7PGIFNQc/3fZrevfzFYtOFyq1hur18kX8Nif7CTQFXY83
Mbl62gt4sN5/HUUxC4Bli/lipUXERO27ee+3UKpB3zSlcF8w5TcmAthpcO9UGgP8
x4gc4/yjGZmemuemdsn+PuAz2/b8s4e54WW0MSveK4+RhuEbBSTHQuAxlq5BvLzL
B0Ma0qKtn8wBG7aNYpHHALtUo/5tAgepoQJcFM5iTS2AxILZYHFTmR5DKW/maQgR
OFjtLUqIUNKueE3Vh8kzFDT8L11/zhOEhE6rPrygWXn+/iNsSWcRW2IP1s1Zewiu
aX3ox11pZkZz1BP/INwYhx3kVQdbjZdOaGM5YS09TtAul7hEUDySRh05AI2JAjPL
BCqSrOCuDfCLffB27xv6E//qNLR1x3ulNlPJeHkMfcAReONNjqVdJKglAHOPZj+s
C02+omJT+BCqXvt/2tmumbx5llPsnqbTtH9sY67W3nSjZzDLEHTJB367ZbCxtd1z
gE3c0YtEo/60mXwAjbUYql7Lr1mlGRHtbXMhbZheMH0woXlzaVFzL0UdImALAjNE
i4NoSg5gCXE3T2vXUI0EUATzinuPOqnpgQwK35GLEL4B/ZOlCT8Ss+vWrqtKaeo6
0pfKx6EdV9T8ecSvmjiCnCksdiqgqWY6N+xuzjjwB6RdTVdHkt/rhIGAKl2SdIBn
4KJpaKT966eRLkjC8XHn45TW8xQZ3EpWyfyWQ4gakKppkoqOl4q59+71xmUg+wlO
HePuGKhvkuCIPJSgfPiXfqYDTbnn9G0XIiH7oPhQwDZtFVJ/VCo8tMaGLEXWks87
Tu0Vu7C0BSwer2RXKoiYYBp1CKYlcxbJ1tQItDQuPDCLK+Lvoqd0tqJYRO0780Ho
DX/B+FetqNLFaCgLiFiG+Bfbwm1YccPazLUnaMwNIvWMfDmUxuUb6YqyfiqFy1H2
gSiboG2P6wAWsG7U4TZwildw+1VeMKFfErOsWl1gcwh3JlTVLnDXfWweqoWJlgy5
z4DRu+yhZvqllQHT1urfjHNld4tmIbTk7D7OwqKSkNmfDZuXeh14uMNoE7EGCCr7
YtcD1qub1vcQS6A0o6gXfm2i4GjZc6/tKKubXasALzIkSlM9RJDp3+BB4Ok0A8f9
ZR4oS8IgNxdsd+vT+K5lmJ8IuL+p/QObmknwLx2ktdKul1FTZYsjRvmh82z36AhO
88YOYvjYd38w5gwaX1arh6iLgMw8RORl5eZOuj4skdptHfbDLT20Pr4F4H+RzII9
NhIwvcs92Vme6WZaQZKc7Bo2qFEFbQ1dge52jfGdsLeSU53m307VHnTOtbibGFdh
u9ftxK9DQHzMqhiQ3uOusEcVvN87qluaAGr9zUB5FTlvQa4HOzYmXDcuacIhre/e
+YasSTbFhQgMdhaKGmPR/tmgIDHFR7Iw232m3Vg8ZyMJyazBfxHHi2qMSI6XIDiV
/8Rhq85855h3MBZD1QoPJS/1GeEauFr7Rx3CRFsI3+6EMhS3SGftYVNfd6Nbp66C
rGIL4ohopO9uEFbCb+SThrH9UeyImvD9CClbJdAEUgnHx+/4GLTglEBINvipdh96
UYQ4F38BjKPk+XjAEEtYYOn76MP9+tVFMwh5s9U2yFoVuUmOEnU2L5X2aocNIiKa
/hQMQd3Aszw2iGcZNGfFlQ+NiA6utiXvIdJ9xtezg+d4Wi3SRQCnxb5GNlRE5t9g
TyD1OSFwa0KuRSxcd7+5Fm6NTBGm5Dv3owwVBZzS5pepP7b/tW+DzF9ETFQ03Wqp
dY67KqOFAmOqB4nB6qK+aWPuD2rKaMxl9nDhpovh7FT58f0sIrK7DHXQ6tQefBzX
WL6Op/QvT9jATZJVditF53ZwKJdD5TUSsilP+GZEoXATW3d60M3D0W58joQJEh1v
UOyy1dzNzWjj2VHAgnlIGSXaFKmHtr/9mtN9e3ShXgkbOLx9a0YEk78Np5w4gMjx
MEuZYQbyblDlSw5dAKkqFy1+lvbqd64P42v3m6xilGOnCrE+WaDshqpb1ZIGzPHa
c0cN/Yah+m3F356qHAvwOnfJPdHOuv2t70I5PwJA2w76ugCQYFiakjxAOppKr1Np
zD+poxRtHHnhbUyOyJlQfoU4CoiO47m2aDNqskNG+9r5NsN/nezMyBgwsYijh15B
5JWvWF8SNc2PpRwP0Z1B9QCZq1sBiL+U8ihfSs9RQk5a0nZq5Mm6riC9UFs6gXpu
Fn8G+0G9oeiPUK6+JVMbsDnrojIz4wnlzuI2FcShmCS9ne4Sh7hAieA6y+UQiRAt
SzWEvwlYFblj/6t2tsgNzKJTxZERW1ueTGFV/JbVKGPXVRYFOn9YnmHZmXSw8kuu
vmtUp2dcxAmjbfF4nTgLJTWXlFEn1a9GR7r+4Vl/k7uFfD2+RPneMMUongw2OBES
FQovanDOcjz18y63qocPMDNivB5XzXMY2OethWdqbm+dfh/ZpiY7BqOR3a+ankG2
LEYdZHs7WOUf3FpniLl4Xzuwr8ziD/huN2RCg7efT3JqQJLNoTTd8xlQpUEVOLVZ
tIIrK7nxYSSu3MACCyxDraXfqAp8WgCzSFKWbm79QEhPzo8EMewg4Sg86eSmg9EV
NXjCalRfm9UGD1khNorVHsUUpJLxK7GXk4ymm1We4RW4+aLiR0N4DNMyepNWysE1
2yZd4XrAwgFD9vnSQNLKgtUwd2kZCnVS1wABw3k/GE5lfvuJk+gFoLBPJV8hBFvq
QAnRZAhJLgSu3VkSYSxXOnbS2RQFIj4Nj1GuTPHXgG1cJV1sBrPX3C/Auiv6ROiM
HunbCHqTh0rxxYsNMpuXqWNV5nu5UFQEdgcbmenbCDhrExuBAz5GlxLlX+L9i6YF
ZkNIuVCQgqqpoPd7xqA7WeGy6ihOjLO0fiJ3zR5/6+c5XGPmkNYFae4jlqmJNf9U
X9CCgQDKiZMvVU4p5TWTK8AkGltwEGNgNgaZrX5dGalnwtc8nKM7MqJ/3jTg9gbC
+3VOpbQ1gbaB+hHhrHgKdn1KmvDb1um6oEetC+Q4Goktsf8YzMgdJIXQ7QtWaMCJ
OolJkJHcuGYKEy+LyXalnW40j03xWEeG2GOxa3Q9iszE1mkX0PVZPeMwH3w3a4Nl
YstX3GF7b8P5YTS4Etu0kNVo6Lom/afkrdVYFX5ThvaNBNzr2g+rwOZ2elbQvB85
H+I9hTipCgZ4lIKGvmk7OzMprVYrXuKROHw5gBemI9hSs/sS5h2qs95RJOC9S/QK
1cPGLPjQ3BP6mWnKrrmWwFVDlBiAIfDzFoEemjKDJN00bGjB23kjdaPLuYnrRziu
psTnuz8LIR6KtO7+uDa7CIZqL09QCWVIwhLbl23yLNwkZjNG+bQtQs8LcpB0q3UI
y0X7RTgUaJ9bbeaix/N/D42P+jhmOM0wg3mqqSMaXIE0UuQNReOcMRlcVevOV/VZ
a3KAAxOO1QyCfzVrVcxKeY0q6+jhCd8/SMqloYzUXLCQczs8A5adHBj5MnLvpYXY
WhK5q6h6GcC3bX9SZ0BIToPBEwxJinqmoTAxBF8Rg9xDLeO5Jofy2r6HBE93mSwO
Kf3pGoIzt/l9j1/ZcrMDzRdcqAMey74rCn/PlxHRsnh+F1wEKDE7c5HsH3JA5CoB
NfFg8g4EwgKwMdpPIfeoAjWZZzduOa+6h+yb6I+Bs+9lJsPiroZ2YIJkl8MNsCcL
ZHxJnIwuHeE9mxxd1/s+yYnVO1xcPYvyzcU94JdD5+nv1V66dCniKEWmaZDDDiZZ
a5LQ/lWDrOLxHJDTP+uHSRemo+X6OpFSDapOleKKVWIW1viBN4DqFGshX52O0zPd
3ZG0i4CFVl1tmbSvHMcHpQW9BlZ3PdbvsUsA3kpv/AvjhbUEjSENSi42x5WbQt2I
fBY33lYppjvw+JLV2owzpqSNZtoh5ojOo1bEh/ax8u0SiYFgUDzu3KV+r0l2PKQ+
5A8FeB6X7pDkEb5FG6KYhtXZQtrOoDm3DLgAWj6gOsLEx2AZafYqCcjPZ52ZSrRi
oQd9ePAnOY7sZSEtEETdzTPxXcli85S2o+QTZ/Q8d+gkzabtV5PG7dqhOGEeR0LI
+KQ1nIgnR+8z4CIVF8zICVy48Avm+TtASK26oNre3ir4R5B71zNgoRxfEYTkjxFN
tXnazWyaBDNt+ItW/H3dxphQuXaNxeJtrO+kpHW5Y4aKWU9lns4x0LxlNh9QmLaV
HpW8GqQ8G+QP+K1/x63Rco3Dj+ihm7fX2rEdG0RlcjRFWmYdzHB1gPrk4DD+zscD
Iei2qby7tnwBhh1KzDqVXLaXbnVf+EnIO1Sf+t4wJciZjbJ1o8pliOntFVt3zPpG
gUvPNW+yFj25yh13r4pVUUIPfIEQpbSwRK3UVMb2cwGbNlpcecOIBUFT1YjHL+vS
L38rsfgoZyzSINzqBywAYVAydPThnoCIU1NwI0ARR6x8wBIZ0qZWOLm7AZOKk3nj
vU7zx8Qm6tsikodCFpM3SOUAswJy4jaVcoNgBBgMlv+gnssPFPOpcAqQJREXlZaM
AnJrNOpP9khkIxx8nyLo0UFEiUg1XGg/DvM1d0V0vg3/XhZ7rRKSVJz2AZLKDl+d
b3Si7YiuMhDMQPcUFQhgH2FSK9uLytywRcKUm2E9AmYct4EtCbUhnQ3g+2jhRqE9
1dKCJw6zAuNW+LHuORNgJLZvuV1LpjtukqHPQ6qZAGWPK/R6mcK5te0mENZv0NFB
EjwITHiNP0OYo8wO4CEdC+mVfhIzyPd1DAmBOUg4hsB0lhSM2hVLG6B3WRjFrYl5
4oCL5GyH2sH0i4yDJnv0n/ozlZAFknld0XwUb+z5Uu3MZYD2rXXAcdSTZC/0WUcp
RW6QfKYt3WusUW8ALq6D3DYAWuk8VaOYs1nSYD46TIes/+YLS8KrjMN1tDfLnh2s
STzGdthJh1RqsIM+EZovBJ4kARqbdkJlb0yt8RekI/me1iA/h4/DxbOyqrcb+CdW
RVMkIoMTqrdjRdpmErrNToD5VPIC1P3qN+5mNR4bRGTSp0h01BBQhAmHZ5Bit1Bo
3teDgQ7dla5NySt8dxdJIU9/yu9URukjuXylpqEcZB3iQ6wNuu3MPNFX2kvIwVJ7
C/9ioAe2X7eVvvrqIcCKeKnT24s/HltzIe94D0PlVtpqBrkDtpo+ZlTl3HEviJol
r8OQEq0M1wEW1jOgluyHohD6Djz7h4SmlGN2R2agvBfKaqWDOozslLjGDVDFAixL
u634arvY4Z29nr/eP+CCJF2M2dOPSJVEZ0kZEKi6EEXBagyDfYAw9cyDDb7ANDHI
33eYAlxKU/lNQXHNDohnE/tLs6iHv1FPZoYn7rxlyS8m7xpmQmg4q/PaNopdfcDe
Ooi3gsITDB46O8gVDqb3m2E76Z0+LSmfhdAYMhLOzeCLgtOMNcghPLpKlhSJL//n
rhGbvOgp0AsblmItgS0J7UJAP+n6NgkP4CaRKl9kNr1hlkJ5jhwL6atX7tODr37v
zYbzJDqnfFYwvn1gE4nERZYyiXdwNRj9AchSi70DZUmxSNEcBmQVnGIvURbXeIwc
EZ8JuzTINwz49o48h4BW+Nu/hboISefIuL7qow3NDvSVoqPh3RXOOQf3M1NclCZJ
60sL36GiLuD0HQBHE+YsIg0sK6JRk16w2bnVQypsRTuZQOy7RqZrLlfZKNMzNVbN
rfwsHF80wvcZbSV3Ybz4fO8uIdB1Bpbx2fMhp+jghe8l1rpEy266A3t/XXdA9WMY
ASWIIU3rmWFOnfcGMBSiUvQtgAOX5ZJRIJ+2Lx6RV6bR8h1fpy1kbuWjECP3bJhh
+sACcmM5GH70R4IF8xfV9utfO5+vyoK+NztRoE+5pqj6xCIlkKFQG4iRCbk2FRgQ
nJAs+ITEOHYseKIgkXj6hrfhyGAOgczPc6eSXbzrsKSL/5+YWceciAPovlDdhXJm
IKtJncALv+B1QlYROrOLXdlbMTTKq4JC6BS1x+op7QdnaUunKcYCqBWnnC4zQzx9
w7ARYUI3NlNEWbsd1mj1fobnbcBB70qsi0RGfh9L8azI7UlBpIlkXCMstPg3T9b6
yjBDGbdmXAWdeL7JAdH17etLgzxgEi2QkbHze/Lv7gVqx8wTRSoTtWq+tlICGFO1
dKqbhQFQwvUi2bmjLZHS/z6orHJe2ntYEvC8SVY6v3uibLYizOitvVlfmpKvBnQJ
VJ4fS1f4VCfb4a1K34Kuh0fRtQy7TmHY2TBW67D9BmD9j3KdIsz/MzAEDota5+C/
6jXW0PwiP8BDT+db0hlaVOuB30r2qCZfGoqjP9KAHoPZt3++DaLeRyEPMWPeQjPI
sUQtvtpeen/JEdV22LGnk2QmS5pfg+CRU1BS2/r2/5vjcLkaojuo9qzjQEj372Zp
ZBnhCY/PboUuDNufOmNrqNNiMtqwicatu9nfoQffhiSgrK88lB73Lox8MoOVi582
ls4vMrqJIaBBUyk/dXlXRjeUDHHVEkUn2uCs9pXaNihiD+zlwF4fplbGxC+s3eAS
s2piNw1Mf9p/HGBiXB38PQRJ+aYhbzm0KUlOCFS6l5AedL2zEWh68VUynG4SVIbK
D+JLbUvgsmK39T3ByWRtFOFY17Gz/zi4RTpp3m28uAsg4xqxFOoiGSqqhbiGioCj
2MS23Hi2s90nYnmFgq4EEibWdAZ3r/W0RlGAr+s9451uxuzPRbDcKftMIp+rI482
ZtN4ALKDM0MAcnyrp4v5Eb3qgGbXar1sZZjen6rHaE/TAbgVB1zhVuAQeaFydyFm
xAxZlYFB3pMr66oFL+X2JiOQ/fErA/Jo75wLhmLOBu9uVuUR14dRX7vzt4awetKP
CdGdbNWBx7UjuW33csfDpYxjDpTNbDGxApCinS8F0OPY3dGCo1IeuYcJhF07RuWe
zRyjSLua4HjmN/kpbMerKVDzjGGjHlKyLHfjBE28X6azTOLhZKAsxhVTH584JrW/
twNiWazRlwzAnh7iPMZ5KVVtHj7y1AuVGca0/P5sa/iZsdOhoaITuyB014R3ziqS
1E9msTCBtsZq4fjUz3hAUOHbL5MfU5uQeLhQi4M111antWxQ+5eVxdcYOtM5reW9
JM+ZWFTCzcq64ctoTZwXLiaLV7O50vnfcxifNE5hRe+BPSzQCesd+7jhfaGoQbM9
Kxvt/bzgKtltmGF9jsQSwl7wHIaXGe0PsKVrBExycFlT8Lq/msNaSNGyXjZPvoqW
QzQjgDGGsGAfFxKYIav2RE9kHdNm0Zf7iRPdzJXfoBVHzbi8d8J1W/KIucuLbmmA
aoq9t0oe8bTZsblpl8esQqCJyfTbiOQXHlGTjcNVjTKCXrEGQs/1kNwmiagBpMuI
3xBVt8UM1oPe1OKdn9UpHZzD0452JokKfvJp9d38OR+1geNIDnFE860cApGPPW+i
ZyZuXfudCdgxZjZA5+OiyTUfX2wHnAeh6jpGzgVp1dtaSQ9BgC4xNeT4wAwHq7nz
uxu6Cq30wdGMkh/NXrkWxAnZtG+ja4S2W35720KXcqQIVbpOk2BKvyiWmMgAapah
kTsUWP7Be6CJICYTQ6PCapqrB9Q9Fq7zFhHaqAJvVeuX4pmcENoddODE9QVL8P2p
lBbpoQmZ2Tu5QIzy4ApZ3aPwGuX6MIloPD4jovqA1TjPurERWWa0aJCBpTabKq2K
oXPbttlvDvlBvEMYSPurbox79EoFg6Yhb+HrUeDwcLqcLf5LAlS1jwUXX+IyqeQ1
wB7pJML84aKkMSeFwLedHxai+5nzG8J/alldQl2jeu/NHX2EwJovkYD0GNsm4Vln
xn3oXjw3L81fQevy4GLEMZ0d31dO8h0dTZMgpqGpAMybtVmyI54/ppAyL92vmBZS
0T8bVjl56ez7cCWzxsG2wlx8bjQirA6dvpVEJKLqSmbO0bmiavpt8G/FKpBkiS1c
TPJn+JvGHSZQ1C8hFIBTe7KUFkiZE8Dr6VNALI2/atCjHHn+OfeTVr2FGfomiVQI
dILPfTDqb3sJKKAK29OOACEjWsr9snxJLnL+nqckOwo+j6Fsy+Cr+fF5qCkUnUkM
Ey6CauMZqRLISey+K7r5qI0ioYYCxgw/k58Z27W1J9SoOF25wwRAKCk4kghZecTf
TZ0wDUpkMqyeFW5XVKT7vWdevVEKy16z2bDBT+GhBzGxB7+VqXlzPYfK6oWuI/pO
v4aZOq8IHUhag5fqL/gozAfzt4o45pjWSgMow/r6gI4ey5h9AlGALSt2t1lkaTzr
qeRSCVtmnGn1cV6R9ebgMuGfTnRsngTPFk7Bf32mz8er9iofzhIZxDmYK8IxKzPr
ooY8ly2UZjTDpn+d104IjBYHLA2RN7uLyZwqrlkmh69P3b7qPp4G80HUil6Q3In6
+HtbekpoFTvAjwN/rz5Am78oAYig1Gm7igPKYx+PWaO4m27InuX1l/Ks0SUz71ZD
kq1ffLYzM5sSBtduTQeCuxV3VZGU5FO5LUv72EXCWKVvOscs+3kwQKnTttgRS5IC
WLQgK5AOaYj7t1f0WQnKftv1ASc3bZZ1CxdBIm2f6HhVszw34b6DNmo0NZfVQCvF
ffva00Jbb3IgYUGSR5mVXXZ9Dm7fp48ni+wOXQmkz5c9pvyo//MBAWJdWDCJWt04
e3o55PQmITSDVBHUGWUY6ru4WSyux0+J4FFh09lmKFsKrra7roFEgJwmjmiT7wd/
+6QABnEw5ahBueKGAvAMTAXef3ROfud6+1FSiPe8EAWpBTEzEJs327fLSE+T1BtE
2dPEeO9ahcKMRB36klPnvaH8BbyKFyyQ+6JkZl1gR0Z5QWIutLnWq4X5x1x+jEeW
jkqMFF96JKGecQcQJZJ4POPRJPkVaA5k+UFGDObRwaC8klmLnG/NkSE8Hgi753vE
paAfleXUcwMh4Qbobn7PoI1Ts7DrLcmJs5amN83qJ5HrJUwyn7lQKWYVbAlW1eRG
E+fMM+0s0tfhpAwRSKMWmoVtTZhJnD0GsLttzCcjhOBL854tScm5NkN7P0itxLII
8Aa9cdGK5wv3uh9hSAWL5If3BdfatSEle5LbMtu+KV0/EhcpTQU/zyrW/bzvsYJU
F7Qi50SRBOBTnKj1rjko5+KlxTGBG1KKuf7jQ0+nYFw6kVTOhZZFV+t9/a/UyVF6
foY5T8SKvE39Gf5evfa0Y7WuqqYC62yE2g7sNbzT35F0SGpMSTrFsngTpJH8dXOW
98AVd5uH+V3BCta51R2/hWj68lt/RV5lyH8OcuESOdYyzxBM+sFsae0zUl3v5SLR
HBEwNOF37N/nKwmRGzHeQ/Iy5Uw18YA7X9nyqrOdTz1sZmB3IvCB09TWl8nbvCr0
DNxwLl+9Izo+NXSGwI66CYCm2d2eUzlL/FOJp31GD9vQzGT+CD9aqWYXl9k7E3LI
b9T0FwZKf6248lSATgbzYtZ/BzTGxBOj8qlA8QC70C6iUStRgiqYy121OYwPw0pY
jcQeA3rDvqePSI0x8zcV2I9hGSxWe8AGS/9QuQ1x/7X0gaqI9sY23Z5PVa0KlBba
qPq914CouB7deJTm+uKeYxmal/foxJeU0snkhxzy1WhXcZ5jShgNbgf+GpOJ+oQc
V8XCGKTRKky0fScPSQE/xo9qCYNFFzv7nVGojKGp7L0qHk9ZZGegOlSaJvhJhK/e
u5aGsjN49zn/0hYhKYRy16ZC/f1UdhSa+5WBsbVUROF0U86XcMRIgTBUZsSqECVR
JviEZnQ52Vikgl9Xagl9NixtpNHHWtJaw7nWOz+EtkomXtT/7Ir7GuSje6cxvYf6
bj2tzjDabsOLYn22LmJjuBzDJUDcT9xskWN6KekbidZTjHB6eIxVS6dksbAwm5u0
Qtt3VtRZWz/ONQJvp4Lkl59zK+YRxQD4atIq14TI+JSITVawe2h8XkeHJ69zmnBI
z5zvrI4cfbrZWJuE4PC9lgNhKHi4uu/ySdmZ9O4dWmU8fzNToIoQwu3/SewOZIar
00FmYP3ikgwUwCZgWdCvACMLDSRtL9WSEv6wr17EFDYTuLsdJWcjc0i1jhEqr5vY
d61XVxt7qBNuR76uEfUrejl38DDdFqJhWgT9CGAQEaQBsPWYfGHa56tgfWbXLcrN
Rco9rCYlxr3gBwqT6ZJ2pnm7ylsk2XAhGL/6mvFpFxmOfJv33Nrnmynp9/xOxCQ6
y+17jqyhBH3qy7plUzD/yhxFX40R8JJD2WZT/RUGO4MyO+LHwk5rYTloz1sVDdGr
X5fjKhcvULU+0/uIanCubqUFakUZTUXyzCt0SNBhx20NYjh37ztK34i88064d14D
4NgvgC4Vn8A/42DzYcUcvRMSn20XZn3GeCE1Mstz0NTL3W5I1IkQV8SR1yhYWIvg
q5lzteVvtvzOnYvE67Bgj9NoZHgvLx0IRRPDDhdsEAoXVtqXGSy7k95Smzoi9gmU
WXfDnlK/+NiO66yZpMFJcE2GXGORH3qbeGVFXHMq/Rv0iT/JZFInjZRcH4ZLOwtA
BNxJQNLO7m7FBX1eK769e9xsMzedSY15q1me06t3nCnI36E0517HfMDbx3wG2Myy
pBz9kT6huhBfTdhZiki1whfTfxy1m/hZq6G5wFh17ahwXqyW9s70gpeFq7OnW/JB
dD5Qwt3qXiJtmPfZxphGB7AQZ78o+XrMEQr3B0O7Cd2eFwrQ/PKRVopeQ4iNH0iN
QWf/qNGQhTAEYbdK+GVhgfclpwxaeCi+BzoHK6gqETD5NpPKvMDDSvAhS/zR4t4c
GUZULsvQ7FyLOO6OdFgft+Y8ZLx5ThsGvZpxHxf1Qr5uM1f/ujvZ+BYvjSGI35YV
4Bi6Np2Lwml2yRiYsbeYWVzZ/sxVOeZ52+bLOM5JkyUR1vi1+R/6g5Z55Iy+VwNP
2QO4o3yeG9e4MSnVq86Q9UQFJK05wf4Wg4DK+PvWXjhvQf7J/4tdCpwM7OJd4snH
DWyszOlX3FFt2ZB0P/kWoMG7ssK927XfdTbDeN/rUFd+kgi4nFmWGj8l7Qee3orI
Fv3bwB7r3YB2STKROcNS5rz/V6seLGrViEYmOk/f7yWWJs68s8hbMxJH5l+IFW/F
/wRxYJ4dWBMtVZBBz9LMCxmwago63pXWHQV8Yz4/bxdemAR9pyctBpFLk3M1jtaJ
KdCLtIAK5hN/r3qwRbeKPg4ZarLefb2BntkKng9GnbhxOZLD4Xiiwmq2qCHbeFfA
/8H2wuXbj9gn5mnWQdhLKFoh1BQL6i9IyqIaipO/385Pn3YF/Lre2AA9HKTRd7BV
4xkyl1gH4PtreClMIglXsS8Xnb5unhxWFSlVfbk6bGHMzSYnhNN9+GdwuYAXxKAM
hweNsFE4HpyAaoqQzy5LrQFsIw9j2TWLrw9oWegOWqXJeDhDCFYOywjzqSsmY7mu
V6UzV9a6lC5JLCE5J2/ld3WwYJDhK6XM4nmG2/OyplrsxN89PVSq3iWEEv1cEDK4
Uzhtff+VfjdNVGgdJgZrlQf/4sRRI00sbOMBmpg5v46keSCodcfUJRU5Rh/OWjeK
X/EheD/j6imG5Unv/psdggaiNGFRDZI7NSolsrM++/3EEsl92TMZ1FdDJJAfOR5v
7Q18sOcDe4wvpLdsQDibtnUkUIm19H6PqBf+aVbVtD9Mb0o3gZk3bCoPnJRRkVbn
xfZU0xfPv59eVwLhi2tAIkCnLsJoyjbu2mbKcAaMJLAj9/yOnfpdmnLiAP99LGKN
HepGJs0gcQ+uxNghpq9EGp0vjQCioI4nqyNnpeFUAvPFOS3NmkK3WppyKLJmdLV3
vZx8dph8vQXUUY6Cmd17JUVf0ze773x9kOgGzTYZE5R1Em54B5gKnaHQSMOSrQj8
sP2x2kzkJDJzBnU4Jr1nQUZnb7tVgYnNxLrTOfHopJvUPr2jJ0WfCeSaBzl4LyTw
AYblQk4PYKf/GuDH6fkO1xSqZOvbMtBueI7GeRL0v+w5ecOcXtxRhm/N5FqMyE6D
lquvprnO06G8d/eKXoLOJM7uJVdVVPsSFfEb5PXHr0hzRuKrKaJ6q2gnEXi9wyEB
ujy5d14JWVV6xOfuEl0Bn+Bq+4zfPz4kvailUQLc9JTHtDO/0odo064jBGaQbx3E
ZvGzKNARiAMuuhFqUzylRofkUA9i093KImpmN0aD3HT2vUsAiax8j7KTdGe49Gdg
VG/h9p440FGBTa/TceRv3yybXSjYYRTxDv3HH044Hfi1+2qXYVNgXaetFgkW8ucQ
3KoWMXCuWnfNSWg8Ao48Ypwss0tFFeMmvPv2tja6Bxwt0fStrn1VRkGa/pYWztEe
lwht3FnISdAZYQahlTHMcaF+tx2L35IFrPAFPxVyUEaIqr/ZFk0X3Zh6py9w5YPD
U5/mLgJ6/jq9sf2EhI68IAf4wtanp9GGFbSqw2GYASq1bRbcob7GDtcvrJoI3o+b
ZfQPDvHEZ7CMCcESo3O87ZPqX0I/U8EaUsXx4aJJkF/UJCduQ+cnXIrTOZwtkLwl
C/2JOvfWWSX0o3/BrVMQdIh1qbNx4VsjwdqpSSaRbKo9f1l4eI0rnhdRbhvyTUBI
XcLYw924NA0jpfVOSYVm8sIqmeR7TLRc2csw8PHztbSGc7iSHGyOvvNEI1LaGEDd
/HwT+0CU+DffEbHqlmB8uh3w9p8SuP+pf0NyRkGlyk9m7hle076Y2eJZJ+1OfyZL
I88E1f0NbRr+nvRvIw2HIkwonnuGCVfxDCegF0fsi4MvyV7uHTzWDmHiqmHeuMez
wIqs0SUk4PWfnTbaKOl7L6gq1xj/FdRdrLlE+rKkhJ4MVCJkr+QbNqd/q7OFmorF
74ugzxtdGrGsNIVXoYNtCpaTh+/b/vlqTG9WD1aknlTl/p/7MJ7XVRhLapER9fzT
ifvQ856+YODBdofugmBzROFfDPSLwCmV8EphV60+Pfege5dOu/ZMmFRZcwgPyXYm
Ws6UgwTbQ7U8wHlQLJZ631oRxZSyFc8gwlv/fhWNcKFzwxwcqr0VAgw7FrXzh+Bf
UDyMlU5mrcrDK07I92YoJcf3Ks8dtjrkH5bh9I1SOD6TCEmID9s6k8op0PvUz7NI
Tm9CyUffRlzt5vY6QR2mwW15szaLTaYyt/UbrgCCoG0DEuBkSarnb93AnWTvh5aE
t7jDZEMzPw1LRoUjtDh5zTmFEnGxIMl42t36giHKuBveLRB5WdzlPQPkILmTya1K
wqcH9I85x2U77/6CKmFX2+n4fahMgocGlPnrhZMIXuyANEZyawhwE3xvf2iIPsGk
Xo1Xf1K+vg3VnqM85wWy0G8lh0UsDSdUmif+bSanMnupx3gZ0Ylsx2SCoxwQ78nJ
k/TOA8vt7+lhqd6/3MZTnMgUnxBCA3SM1PkjnYzCnrT8mRKhE/gRoHx9QYYpZQrG
sLO4lLOvs/RQVKQGrhfooU20bgK5mWoHkv2+CRMkpIeuDkXCDlHlytX1ZeT66UKe
fUQ/NOiBIjfnsets+DbVh1/lRMLmHNczvaLlmxwgSCkUln0oKTYkTIu7uj1HCUrX
zvKAGFRYcNFFqlQ+OYIX+asnB1VeQK/xAUPp2oESZBlpaKq7ZJ5K1OkosLSSWfyU
nK6DLZDBGhP/1wfYeIALTXOVa9sm9X2Ip05MJ3md2NfFd7rfNGl17y91TBK7FY4i
j1fQ4r76fTpofssMyJvVpvQUrbMdUgjpRwvQlDY92gt1to1Sw8Yg8ot43yWpLUjW
+bZ2HA9rFZImZAPxV4usnHLkqcGeCKmngaHh1ggP4PLAYExyINfRCeqWudt0kG1t
t0+DpbmUIjn6T508YNrJOH5OREzA1O3lOoL8b1ymY8WhQinVBwiG8HkQaneg90Pn
IWT9AGQQ37fXHmySqChp3ENQcRV2u+oW/RYeYnrHTlBqH4jm0JDQh9NSANCvvcfp
MwhO9nfNJUf0L9lp4pgY2SjHEcIPO3mUTf8941PB+CPqIDne6xZMnqz6wh9JlCts
O7lEuSVruiCzbt21aBZIHAEGXb9sXRVZ3q5WNuFgBxE8jMmXsY2isQx/TQRBh6m3
lVOOKNl/8t0vxvB3tIuzbeECP+HcVO/m885m5S1LtiXjxcaISB6uF/O+V+eDAzhZ
aQEDQU4mSngqS9D/BvKjiUn2//JcqONbnjxI3f56uvKYQuJ6zbpY7I5+GxAE6rYM
m0fV4uEuBKDv+jVIjtTha9OulobJFlB9s6EwWXxlqNsLxaQEyP7vIwtGlHFhFial
aEwvRJNupwtkDOXm7kpu6mNTbBmLr6WTEW2zTYiZbG2fgRG8Cqrm477A1L2PKTQg
cv10wA0+S+tn5AzZ5DLYiAcCJTpBCQAp3KxTF1l5DVR3qVZUBtvkqw9Gcr+OW34V
xfDAohq76I0ooOp2muGCbzyWbB+7b3ZhX+tDkIF5vO4+e5TTWOkFtSM8f2ACLQcv
UAj4wJJyxqlFX210KBKX0nKczvp/5ekycRTENGZTNvMba8QnEMnOIhfmtDe35hEo
HVc7IpXc0qTUChlC1BxcSw+dKFxULgFKsHF/u8ktYnGJWpMRS8ptwprgyIXSckHG
L5BtCKQPPtYiJS6H8KLjdSU2ytHIyLt6kEOEqoWhm8U20TMYL6z5ehwfXX8z2nvC
8+ybRBQqbuT2/PXzEQq11kmUezQsFWjItSnCwqx1ZQxl10KzpHjKwA0O9EtbhLZN
O6OqO+coYJNk7kNBGpEOBHu2snbM6nqOmqSI50qjXRlKL28VwvfGTV7TZ1ILrHfv
yt/2RLcQ1X4jQODi5Db1U4/eZSWIwx58EoeCGUoPQLKVeR/3tisC7g2AfBgXjWy8
egpUOLJaPiOJvzwcnwyXC8g4meUq+KzztrWeuOqkmVRQlTAVGVpEWA3ZWOEB8DpV
VxPEs2gJJ6QEz5WXz+93B2HkwlzSQ8zofUVM0cEAhltIAys2zyo/fpCGARWoaW9n
f3lmK1T3d8aV+0AGYmLRKyg02CS8psvwhPKm7ROlm0eLFL5aS1Raes1iWE3ZR5zX
aBAo7OBcAAaJ01/byPeTFjdfM6k6SeZ4xAA4oMCSbnaT1O5JDu7YobawglYBpyd9
RxwRXXqPY8LzSJCQeGPDi0UcLurtasvYDxmiU/ZOb5dyiSXt+O5JqgOPvzoJGI5D
bMFouwa14Yt/Ksvc8uRjUacSLTdwEsnjOex83gWXXSFwFxlpStTRNO/gjjifCLfM
D18QB/cRsOFT01AGKGmHUJYqarIklXhs74DXbfjtiec+g3rQcER1xkusQcgpLt3S
ZjZYd/KXfwmBZXl8eLBePut8FLpxqyyCR6ss2ehxG01b/uLSZGQUPQTp/Qs8rfeE
Hz65yT8/tPcPv7K/fY4ANXyuwTOZdnMWLeoqbcF7lZERUvBa2/lF9h2h20GhJSFO
5Q0Tf1oMnIlMm3KigOUVwS0yToeQg0VYDBr137U27fJ7UuWcpKp3bTcGwu/uT8jp
owlTkI/x+/35qtQx/J7PwYxnIjDnNZx3HdRynbiBSVp4ANedkdnWA4NIMf5CmKqa
haXh/tgAbHWf+rb2Ft9lzKwQJyGlCzhcYkEF4FYa4O2p+zQzhl9jLMYkuNeAtHI7
EfOMxIAdN9e26q8j2N2g8yguHkii5/2qU0pjaNdXXCoHQjhIcUozfa3EhZle719M
qUX7wbEFgON42vvV3hRyVqfQkF3SVo9KRcew9jALInhEehI1FuUNtxqRE4Q0zQRU
iDyTFbkivwDYor+88zOZfE5U0qgLWUfEtCeynwrjavNafUh3crbTPGrvgSgoAyro
A2FoLMdsfeSmmeRYk1OFQeu7MPD9hkmCb46zdiaZmt1T7zvg/mhqonq3wA6ycDa+
wcuTE7DFxzCuJf1KJ3fpezfXhi2Zph9Ory0Akd9meqQAdbuU+L3Tvz71oINDcX2/
Cg8RzMMDu/aLYtCddai5g2PlP5rRnDlagR3/ViWEqihzl4w6Vg/GERu7k3phNoTT
DCaYgHUI2Tzn89PzthehhSmGCxGcF4yyZOSYbUt8Nz7MDSVgdZWlmqRMt0qYUjqK
3nCMRvwlbRZJCL/jYXrN276UaeB8Sd/y9lyZJOzSke9OazNAu/5KIOyWnRyEhOhr
cXW4uusPJ6PnmcQiOMZOkRoXFxUj8iKpNVuDhRPNj1289QfG8viYeD6q7sQNJvP8
sI6ltBqMLW0ORXnO+AZYLOZEbxKtBQvZXYBW0Cc8A1kTGYZft6Rd7EgXZu9MX3HH
crglq/nT8O3fIjvd1WBJztaJXgigvuTJlOj88UaqusEOOH8Uj7/BsebZf299Ocgh
UZOrXF2ab4CtGU8XvzxkttCu7Ws3s+ixp28dX+mSXfC27SYHS9Z6t7BFE2i30F4q
WSs0fANpytS4FwJoCU0UpLAVW4IGE44D894iymb4LRSUhwTcI0+KhxHLnXwC2p5f
VzeS8itu84aNM0y2UGhH+rhU/PXb72IddlxRNvZPetijlCx6dLCaqzvrGku1tiu+
Uy0Fb96wgSeJKJo1D5luy4nzI536/8YcMRz/N1iMBHTjxVb0Q2VpKxb/QSwgODI0
0eHBZFiq+rh/rB8RX1huuon2oJ5pazS/KBOxrMOdzy13MHnXCojEdF3blYw7l3vA
dpiT2SlfveksQQN8TxUehgm2V8sC/c6+i4Okw83PoI1JbYTPlT6gKMpnmRW7tx+w
0Ywm0PKDjkICZaoksF49RlSGJV9trWK/R04b2HgCHK8H4uCp6T6kVMkYrO1vNk9V
nm3qAHLxnftY2owXR//jkLb3TI7xdyjR2o90LixWKGlCmaxGqgPtatARGlo6Inq2
pJsLxP67p77j1DzPwyxtDUWUGyQUl+Pvza8sOGaHcC0JxNYrcHF1+cZG6rzKU9R+
q4eUkj3gfFdrEqyLp+rakkJ6Z5SpqbpHUcX5vKcXKmh2lZaJs5U4TXXIlbxXC3m+
bBhoPrxo6kM05uOMGjmRYqtAUA8z1/2/iAbZu9vIbFfyYe6YvuRcBZIHXzp01VuN
Y5amIsgBVTuEB5bQUxVul3r8mmGmGHoPD4WOQkr7Ct3kbZOzNrNS2sNZ1329IsV1
tZdWVRgZ8iOS5RbNfw1pjz61GqfrUQSFJdLFpKL+qRZXaS1QuXr2mTOBC4XzcPHi
XQ1FHXmLgX09IXA+yp++NzpjeeBTDKTkRXqdm2sJ50NuavXIFmzJJL9YoSTTJ9CL
zZfPtoELJfJ4N//y3bPkb5+HNaeiOUxBpD3zThM6DI1HD4eiZLwRxomQZv7qBx6b
SSfYldNgdphf5FymxzMH6eBtveZSCmSNs3Y72f8fIThKVEc+2YdDLy3EYOF3+vqf
8j5D7/aGXb6yaeVaxly43zWLN3pizZHGJywLAUFlMg7LGTDjQIbETvq6f5oSdaGM
dG2ySQKnLqLfHNuwfUXLPSAxDfJmAF+9XkLbKtgxUoTB+L3E0Crks6X4sBIsdnwE
6UmZAcUqhuRH99y0Z5Fssjy4i6atOtaAePKCAh16gAJJnlLcLOzvAxbsuzJXlqnI
RIxiTof5PCkOZy6LIav7VFKMH27JbViWgyuNnKwpcnvvW+v3m/0QijUG1ikkOQ55
FGELr8jFuGFRBtC7OTEc3DDA2RVzUhU1SqFLt6dZRF+y4xeYE/bukEEmgjWB2jOJ
NhJifGLck7MPOPKrCI9VEgosQuWMG5u+zPOSFOJC+JZ/t3VUN/7zMeAgRN5gvVqF
T1U0yb5aWnfcW7gf6R6NEJVI4Pobd4TuqhSuZfdklKuJy0O/GazTqMel5cTB87gV
3zvZpuJ2ZN7DOFPz3ruSTGxcWpedr2NAIQNIE4J2LI+4qxsxn997ybryGgavhrcq
pSezqxBsYZ//hIcnMrAxO6xsQ6tuFXqux8/YzoRRDuo42C+cgSfyAY0Ox6Qhl/do
fjPwCLcdzwfLTTbwvJ3QATlt4S7WXFUNjEVo53TTd/AOb8XMs+RjGsGDd5IQPG2f
FcAg50wlrHSh4PWmk5JqsTxw0cWf041tvHSGrjTMo+/kjOF2SIGtSC1Dg5ZSsFjl
MwEHS+j8WXeHu4byKDKyyjzrOuYwL+FOlplKkt8nlaBK48uOHs+lzadGayewwKEo
tPU3JRSBS+fnyga2xDLYvKKzndVCL0YGgy//nS5JGIDXa6QKWFJDfnCCHIpRI29X
9I38bwkkUleyIbOdqvBU+gvD4p2/XSlMP8LVgWBB5Kc0UrihvkY268L3mcu/kFki
VKevBpfkRB4hY5YFlywPXIq2iErQS0eQzkzoVhDQnRPG9Y9yNaf3zxKcl11s4PUs
YihTgJ4MuhCHLbkPOzAJRyelhzZ+ZlyYyG0aMFQxLrjjqI+TFQnxD3/f6ozozHER
E/GAuCYKmRlLPp9DAYmclDpr1TB29PgxDielIcO3x6BIYROAKhoabf6sKPidc650
8wKA0HD698p8FxhJWg4xPFAchn6gPeCpKqrwtRSl8gz0bSV2WgRXZF8cpz6+aoYk
Wb5s43ahAgxP8oVKt6Eal97PZNlYDxfiOZad1n8DGeu+41xzDQ5qzST1t/QuOAQD
DTJ7PGd/1JzRILwJBZQcf5F8ZL9Z6Iec11z41WyxUh9aXzD8IVZYw2FwEvvSw++D
ECOXXFtZSIgDHOMDgHkjhiBckYzA7bvEmsP3VTcykhAh7Gdq/dSJ5jFn8BB7DNkE
/qLOAUywZm8GIHzLzD6LGuR5MszuL0jqHu9UPkBqDyshqKnmTqobpwJGcGvculKK
xiB2A0KUEQS0uAM1rh+Kuk0AhOUbFnpnYBf996kI/N9NXWs23BzN6/ilHZWDRLYR
WHC1Zn+iwB1q7lxA8chFH+8NvkVU0ApgVxMxmqYkrn+AkNr+HceAw7tCORM5lOpi
Sw1Eyqdnty4Hpsg9CvfgV+zyiOh2Cd8ORI/Z5iCeroWmygiIWr4LxQvne82bsdkV
yygGOIbjFG9828YkKw9oqKps9mTvzAMx1nDwkCUWVtTDBczYhlZNtjwvC8y0CSd9
OUHdI90dI4Z55WtJ3399G+s4WWfiixBDlHR5qTUsA18RWyV0pGKAxTfu8yZvne/r
dij8Q+DHPxqkvCjxcDr78c3Y0d9bAaV6HH/3cMBoxUdJflKvu9v6QSMTdhocMddn
fCS/kLriU7AY4T0qHAd1srAGXI1Qtmpu15KY8KVsJJ7PCYZD/G1XQHihr5TeyH34
r5UefqT1t2i9LTvVXz6TbiJEtC00vxeF6YUEvKGOohdh+eVbiqhaT6bNaTAWBm8e
mf8U+xrnj3m1BxxSCWKGQEX4gwLFdzeR0MaU/g1UcxviuFfnfEUif4vT0co3uhFW
y+i0pOhmzY58opQJGTOBgtpLvx/mCQR7/eNz0ogMDQ351uOhVpdFkDv0+nw9q1Rh
xC+YneB+iDtjYZ5xbZpXrmtnTD7e6moLvcQH59w5cVxAk831hnRjUTljaML19vdK
2Y449DnS1xzHkboENH3P3y39Tz73zXpL4MMtWcOGUJJcZKs3rB+wMct2+NeekW0u
73pFC6JGl53Zvg8pHgkTUoNv45tuoNwiNSJ+fIRS7NF2w78lt3+HxkyI8trgwF44
z6peVMnscbs96bj3Om0MX9HNKXjbmJb4WcXmsgmKl0TZyRdDU0alXb18HPxWKCii
Epe8qeJQh43R4XSDX1z5hGbss+bXNWu78O1hLpGFHkHmhJt4KJQu2Sbt5TiDl6pA
4sa1YtPShLcEfuqe0FJxM/78yp0Yam/BY4mmPmN9pYmx/Xq9XLTrk6fuBL6Qx3Qq
HQPL5iX3Pz3gNARW+eph8K2wTJuSnXj+ia2ffVsuCT8uDHJC92iNOnJxIrPhGG3m
S1L9XqRh4roZ7Cn6GkaHDqafV3VwoxZU5HUiYqYoDO8J8ujoARld7aVLoD6pQfWZ
DY18gkmuzf4RpnP7vtcAtVGtYl939nCyIp2uWlWKc8aUFFKMEovIJzKE8nPaPF45
1BYqdv/UyM5lCE8JkOiFmyoJ+wR2lfz1KULN7AiJeWCRb0OOu9vj6wuuspgOVNNq
bz1njs2dXZgLaupCeNMXqLqe/neGmfUGWBNITZTjXMUp/riOggci1hcj1jMhhKY8
gpPk6e1vFZV9o7EFBivyYcI9IK3Uqu+fPyoLUTJEdGhIPXyHoOH1ydXSOLBvO+/z
dLHMxJhBxOtyrFR39ngWNLboMlD7G36shzJH2D+mlEJTObh9WgHhI0GcKY2XQ01R
oY23Nz1qzHNXGRqYMzgS+wr+p0e4nayM3NyIbe4g0mnZmUM9kPWZ+QUML3aNlE+a
P3x2yTdrrDd4an5yzRuLTOSZiy4efH4bbZ7rJk7mMFwFYg2tsrAJIP1FjN1vSySR
/bG8Pct/ZwxLcvQPHHBU3TyBug2zpGwUw9luucJeW1c8BXAmgH3yA2vshwqDawTX
VGU21p0wzsimKwZDeBFyuHIIy2UDLzTGeYhggPx4M3v1n/kib9SPqbPeT0PKGkD1
mqHQYAHb5StSUpOcENYv5+kQTtlnsJFRBmt/EjXTwdWQE9o/ahkwPGtfj3OBDy9l
yF66IX9KCRrSQCvt95h3QLrmeEdTPac5OwtiWIZwiNn5AXRsh9pm7pBVC2+0PMkA
eXKHBALViVFTNKMva2L+QdMrurCBJm3l57D/MTNONd9K4XieLPktPw7yR5BdtA2i
kbCEagkYQpi4haN31jxgNemk1xEDzKqS3yyv/BBW4Pathk2dAZRDIl8IZf3kGBul
vNB6mnblqvdR46B5VzmC/2TuvgwzrneE772MuoRwiN6c7apQBPmE1yXeiv1k6Z2Y
roJ/UwfeE1icGKcXiJecjNciFUMQFJ4ahh3kwxhV1oXUmm4yLKse8N9lc74czQio
9D7Xg4tP79WFzG02kYampCfO+tkPI5okcNwMgUD7vK2JN3v2fePONkUSmxvPq2pF
bKetwHCHCmHT7toMMhhf7AsABioZDMUlOkSxnCYt+YIpWL6Q4Qms2a6pcBvDYnoQ
0Qg3kq7BKWJGp6g9jAFwNHSX9qNqp/xYhStW3AYKxHl3tuBGpcJCRns0N5uPlmd1
8q6tqTLaoTiTb4QYdBFMWtzxFp/oGToY7okEthbpfRnjooSXwwUOJVarAc1wyLl1
D9VUHRL/Bct8z437eXcLvETj5XJ5kJ9rAOvUfjb8qax1k228qFCuT0Fh6fH2ozmY
L6kXQ/DEqSWkq3BJvzftcpBtCf8B0Gq2EErMzx0JsGWleRmS7nqTJhC2mILvR4t6
p4Z5YH2E3s6c/DClPv3sIsuTLa6EeZ/fSVLkLDhjZCuT61n3/n9hIZxws5mZsI/W
mNJgjKK5ATqKMw8jQYcQccWajsT3ahK9i9SJNgtnSi69Ybo/UfQxAj8O5TGHcosE
VJq+PTqSVxfczAyHM7NycXkCL7NPSF8yisfdhmrKeRfS5jQaW48WSjZDa5GkuyXj
uWR09eLG5kwJrFfwu2GI8bim2CingPvm/CMnESPD7sp4ekYfPrx0tBDRFIQ0RQvj
2G3xNGhxhWZ5yKIGQMBr7iru8R3UlskbYQBhkSpZ0dOqF2lqFzKBkwAeocO7es97
/TzafHOopq/OirQujix6pCcdKA43USwuxhwMfCBLNNllPQxtetEC0BUzoe+6VMlf
o7DZt4kDMMDeFQOTrcGc85yFrDQ05bp4O6MGWLxTGTmTW8gbUGVgPZNJaFV7nH0P
NWvOf9Am5N52peRyjg6e8ijIUIyMNW/ugHbzlNDuOg8hBWn+Gq1mhtd5Z5Vjf1SR
IDaiyNc/nCXHD8M1BL26mv777w0ZXGiyiRzzSQxZDTHoDrpr4gighHa37tLpb2iu
14tJExSj+au/4XfvGfkTjyE/RSVJATeoY3vRGv8o4xRk9o3yTxFoPnweikFJC6vz
EhQwD176bsN3ZnTdbgJQ75PSagjnS2lwWZcJb+ROOXkrgbBv+Uk9bfzeDqk3nA5K
pfUc8e3myFG0vhg09YNgV3MlLTeYqstbu1wZHgMGoPAEeiuG/zBgzIZPJ5L6ivH/
zu4/4qNVQWcim+hAaewaBWoHLt0gzfh/nxCNJldbFlIKNO9iu9B6jmLR+whjXe9M
p30qsvyMUJHlWbs/vC2GGFJmTGwunIiRwPFPnRZwJzXj1kBpcLvBTeKeoriz0SXI
tlyzJCx2Wy+FkHl76dGnnkJvOH1k2/YrigvMgtsWlSDdnQpPwA6PoolA2aKZSd8I
rfm9PmM2WE45faa312HY534BNTMnIaC+rnD3/1/08F/iMSB5G6DZ7336MpBUxjlp
HTvRtj/hDrZ6S4qg3LO7EgUwlNrEv7slOXutwsK2lLYsl80Bx/wdUc3EYQFb+tQ0
WqzSb9BvD3jK3n1o+XPEcLvRlEEyqeb/3uOY3JXTaqB3PlBH7FpC9Y1smOedfO3L
hqBfkKXmhdIL2LyfTav3T7dG/lbbICNww6Z9ba91a4rjvZGcdSr/hS0+OUrQW31e
WfzgXIgHLEPBibGrfO4Zjs0aTitj19uevwTXd5BYNdmIXzkIKhYQtHWRJ7DhEIUj
IYWnOrofN0sfk1J7sHlonzuRqmSU5s6/JFwMUILFnRdQPBPvWiNWFRnkf/1rQS4h
NrrNTU+CIQsywJEZ49T8rZvCwFbdLeHPuK1pmZVA4dQL1eccdTidyUaemOfIfHsY
zg7D3F0N9bkL5VtoZw8M1rqORP8ua16XevqbcQWyzlWAcPLQsA/7NV+4/dIhqKT2
9ms4v8xIasJxyT+1FXwSiHHoRhJpFcmzyPE/fzcthCxOg8G5OdL6xcN6viKR3VGK
2ZJSMgdVC4NrUGiA72GR5WKPxJ1FX+s7mDX2xaiKzvpzWLSPfQMq4ljct1isJu+3
slpSZGCMSQxTcoU3AW5M76StVdg5d85sP5DDtETapQTVn5fwNT6aU5KEqK52qlqm
p4mVSUxO0G175318NasiQC+gwuAlAQYS5+T95BWRYbwgyp89fvq2di+BQKwgAH8+
Hn0TuOk3tM11UsVF/7rtPO8xqwRh0OEanNOKgI6BCSnPfn5gpSttCyuj8DhHI0QD
XU/4VB5Kpd8t+u/zQHJq4yZwqxpLHY4HmUFO7tmfohTm4CH6YDJGXx7UUJilNrRu
D7hjufunW6mvAG4CjUMKxExqyF7b1UjhXUZhvJuIwcTRkYeSN/+TYZ32bkoyMNCV
KMQiY0srZgWOf/9ZFYuMGkGXicURsffhthrfoLbmFZ0n/gOk8wp9ymn6Op4wA4Xt
8JU4ymeU63t6C4PIo0zIrAbZ0+gXhrw7Sxeq/46x+5wSBsKTu9oVynlWfwN7++Lz
VL+DIMy8mwISnlNJmKouR8aosvXj5a/drrsjSbiUDOVx0Cqlz+dxTxM60Q5HVLrY
v4v+P3azd26gLGyPLjQls9vulKX/laiKMEXi5Ffwt8NRnJVITLs4gsMKVbBi83N8
Pj5Y7d9SKCjnS7OV+IHhAafBZyGrta284xTl7RVpOwk39eLzzloPGJMYLrEB66yr
7Uu0Y1nDrv3YEVAxmdKYywtTiMAlcxQx7wmgO1kptG83erfRP/HSGjO03q7NTNrR
uR66/Y2ovAp07TrYp58JwOCoMvkw/jNmrkFOhL7HQ9X/6FDu8IZwu3sWjjDfQoLD
VjTPXKosi6Ud/I+V5ClWi5TiHH9DCeuIL9wRFlu/dq51BZRZ9u7Slv58IUxL0JYP
zyPQgGXgTdk+kdOS01qUfFAgoEIcSj1KsTLhA8gZmI87BW6VkjVqZMj6oSTMO1Sc
0nvWV3wjEhh885HsM99UyOBiJvuD0mmHcWOK/TfBnCVAFl/WmYk/R+dPxoe194kL
ZpOzVP9eVNc2X72bK4MErRAZ1aigkMI92nO1VpzNhHY6sNVi5g/8MBGCHBO+8RuP
8+6xjvph1A2KrFA9abc7zqUSEqvYC9IkmUGjWqj3a3V3vr2qpJBp1K7b1HOV1r49
2l3kU+feUd7lv06hO9iIKrTdtWipfRY+1W8wURQ9QZVsBQX47Z+L3toOMg1rl+yP
ZTDekr+VXnAUnv+OFnc3Ohu83Zz/zh7W3dXI8bDev3Wt4om8ngvrvdtXITLb4UQQ
6JtjljRyGWsMcsLgm5d4gTmf2m95oO99pkHC8ZGIcoTznSRmsY2U5yVlnN6FzIcv
QyfM8+sE8EbbA+nz5y05KndsctH256GucppJf6MyklwudUnMsA+7GQxFC/E79Il3
mTct0VpJafV9mB+wluynj5+ktBpZXPk4xqge5eVAqVrB/Qpop7lfGPBS6MtTt1rK
ajsCoST1G3u9stGCI0Lp8f+bv5oFb+sPXx1YIk78ZZ2d+IsMxlZ1ba5Cwmp5R1EZ
AyaZcQXnCiMdPiOuZBtpQeCI8ZxXxB2/IPd3IG+FD9WMZegge/39eIy+HiCNuEkR
Ux5GHQmwka5+QxM7pBLmbAOM1SBRFuiaM/q6Ku24gOX4sAe/vYlEdSYW391Q25Rf
qMbRWyz2xg0lhiWgew5ipHuVP5G28q78PyOEU24Ou/ha/n58czwbVcGUBcyISkEa
Q7EDrJTXWUUJslzMVt1/qlyOfV+YF9pNAt1hQLGKRUOd+jtfYMnXjyo/SdgSA7JG
oidJgw9SaJeCxgHmsOBkFoXN9aeq2h+Bk9epXjNuXtRAlZ7KDGtndXL65aAjratA
WUHM5BLMIpRwaDZBfTJTzRXWBVzXc32N9TYG64N4FikZLScOHuh2edrNcqRggdbu
Vf7lGC0P+Oy/Ay6/lSvxjIopPi3Y49xcCLJD19IRIUfN0/eujYrpYD1/mEhZOBkE
Gm+TGFaClwaemhmofWaltpf26NRLaEZ3qKifNHYA3JeVyJ/3JLGOe3pQ3JMZicdQ
9C55u2W4HuUZTtLJBxpv7Z13AMctUWOANR2Px0VxQrDPmWBjhE6JejaLipXXydtS
Ox9vodRrGfEfrLCQ8SAnj3epeBeqKggYFW838dme/6czJ2Q0kU6JUZyfoE7GrNoX
pxZpCytj0c64QkGmD5+eO4uEjbmNHKdzqcQ6ghUxRBKuJgJGsbdHeAZ0us6KSCCR
hsCIXVn2xf2i11OsffVQ44hKdqZNCyfsntspngSODM2JoavXXMc1mPlzXXMxm3aQ
AdZ69+FNH+T93We4nZlNaTU2apc0b2mBtXY0kNla3NSSOlTs53Y9sSJO5lnRPWGA
juXz67VUoZdmvWmXixqFhvR+b/ulcZ3WX5dGMz4hwIEzDpjwE/3OC6D7YKVPoS5p
PdxxOzsh1Ki+MuUJxkeHLcfgbiH2vFuHwd1PktgB5TnsHR9ybwNs3+dqHRsGJm3D
CPqOZS7lsbbMUns17/56UiHq0Kyj6D1S8Pt1xEZeBXdI7ON7sw1UpCNefhItBOSs
x9FFyXzrQ58pDgAhybjQmPW4FhpBDPYpE8d29bbHJlPVprdWPb/fDcEj9HnId9OD
BiOQakz2wP9VeDQU2iKhmAm7aHbLb7ABhxuOXaLFco/xW0CUUB6J+g7Bh2LVqlSr
R7k5C1YBDzgkg0gsDQiQupyTtYXN2sw/GS6nIT8U3P2o+NTeYwZ5ED3spI7DLeXp
TlvAjmlx7gXd5qpljUSHeUZ8jJVfuhTrhREeJkqzHt2bPvsnp6lo/tzYsgcGQnxK
hQB4lDTDyBa8wATO6SNz4Zp+IVT04B6ry06mnPRwv5lGGH+m328mDNV9zxc71x6M
oqWdYVL0yfi2Ym6For8DgvWGmYYeCVBblN93z53rlfAPBj3HHnb0y0PUsrD5uy7v
7I8g4Ebtomu0MuEJHNDEhVl5XudzVvegzacleqk2yB/ahQDIdQmbI0Gjfxs+soia
cGVR99L7+dARo1kzc6CcDh4nD1RsgfXMDQfvrvg1xbBuHZYsq/dBkc0HVkpvTmlG
rYuwdvWS+49aez3VUKh8VbRSDdkZiw5/R7J1rlBsgcNnDry4sLhQ8NqKvwp7SQ8c
4DDdp2JPBOKaBOjcR24p9HJZkBbDmeqsYKFLNr8ysk3K066zN8QiLPXo13ULLIgt
6/DxUfDbolBE0OTWHkOHrNtjH0NuOwyW8mIDYr04qGBC3q6oAJu5ymC964KYb6zU
PxNFECwWBYg04NOfGY2UgEIyU+5f0g+xY6ZhTmPz4SeyWsYPISmKOHdVKIAPqxVZ
UyxyTSKqZgrvX+nqGEiqGmKGPRmh6GcYhydt1Il5ky4WyV6716MYa9l0P4ie+MzA
Yllp22VHYz7hNFtAcaIMxuN4ZZZukKFxLrRX3m4GJOCe67Y6ymze0VuuJdqMpitk
nFJBbYcHOYj2p3k3BRxQYw0j1b16/moPQGNP23QFtggVgKtbihQjIXGrxVX6Rny4
SR4QdnxkYXtb2CmxnBiumIKkpLPC2a6ERCk32p+JgEOmU8psPkBG6PtUAJHWlVgD
zo9PGIjUTPPoU5cGQRqMvHxqWx5bc9N4lQmJiv0rBw2nBUlmyctAfZ99/Z/bWnjy
I3UkLysqfBgXdTopMD9C02ZY8Zk/dpUOhFme1q5kY5IfAGMRzuEjMFu4CMWba4cz
LAB58vxuJaDUvmshH4nEAEEU7dpmwBckfhVVSSMA0iZ/ctQ1sU6fKUED5o1JQMHq
lyJt1QjvA/YjOu5B8pJpo7q64+qaGhFxpSb9TzAbOKaS1Q4pL0UKXWcMRDbh4Abf
wbs0dJqKw1lI025/nVkMcmX3PHeJYLbN6IHV/hd8iWnahRjfxQhGtyXErSp7n+he
VNB8LyjG/xTTRc++IVp+TPY4t26AZPrIpg9PLem/OaOKFnJ9PFNlFeHwfHoILat8
siNuOYBq0kQmQqBz+UmxTkZae5JJxU7TAfBYeDG3Ul0szkjx401jfm3Nyl+hq9io
ZR8ZPPH0cxLT8Vi5MizlKE2w5SAmlEwKFEFrotNmxNlQmJxySAsZ8SMZsXfpkccA
3FoiagKBER93niNlcn2G+jgBNPh6cDbfMEy69sgq3etq/iyjuc1jmdvngXDCHXVv
dNZ3g0Pa5siUWKl/RHHrUit0r3K/tnGmhegIXnNPsZKt26Xe4DCoXtCxo4aSXWk1
vho4dizl5Jw75hcgKO0B9/t6898yTGImbimS7xBwiJg=
`pragma protect end_protected
