// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TNUTdJ1OBKF/IYrWQjpxf1N7gaRgANknt2vi5D3k0K6Dqg6h3qE2Gj30F52xrDi4
B6MPSZZcyGu+fTol7mwz9bS9cypYbBCWoeQE6fCWSmCnALW3uBvQglG7IxULgJgh
FOLJ5gz4VNurAQx37mCsg/IF0QlRPczo0Qj4AnXDEIc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26080)
49zdyrlUJXoLtpxz3kvOM5eZyk3SOVBw+KqqBxpcXJ5yTZLMFaMKAJTZHTqAExu3
IE4vgh5UHA/icTt2yintL89ob8deKh09/4YSQqrKa8I2+YrPoSpfeCPQjBmUJbeB
yOyANOw+33Y/AHhqYWWQ+l+I1E15J+Wf59BhHSOBGzMMLArQ8uXoJY1dV8r6/yBe
NbPCvzRHAdQ8hXz1h+S7VzH0LBOP88A1eg1HTDVZWkgH56rKgv/S/R0f0higAkAk
BUl1qDLjRtpCek4Jj5ly/C9vwlC68HUlJJM/GX351E9U9RF8+Jn942d5+AR9fgVS
tW/uHzzYDRyzrCm2NzNPBwyNRY+J+2hzkNzvggn7P8xRvf4bHAkbGnLa3vy6BONm
4eKDIcd1LTrMseYB5QI+CqfBhwjfBPADsUkDd7q2RiKVyleIOM2XLHWeRWiQsH5c
vyNljOAFcE3h3j0SbBu3YhrlEIoDPU6Ubnet4ne43twS+VVsdMCzo/dpPcG+WFjX
pkmrFfotyBg4diHxcmW0Toj4zAHsoHyeyoLw66kLfnl13bxgQ48o8VADFOD9gxYZ
gURRUcgztHC7lpKQagYuE721U8u+HvnWgEN2It70cMRZJf0ymt95e14X24QsGCjU
z5rH5/i5e8TSV0T49wmd1edh1EDuF9FY8qEFwnXymjPCi0Drx5FMNp5PxB1uJYty
EXrxmjzVJfG9OS/5yKuDZE2IKom6qS15CG/9ndMDDSQ7i4n6VtllLCUXNmYQsFi4
4Ru/CIMb9q0NqD3L+pKIzL7mlTqqoeqLCpHfFeG+ozjaPxT2KbenoDKnaI82nqGR
hdPXhh/RjE4fb7yx56UUofBhghzpIFUaKQ45RocXIFwZzfTUibu0eYGrYyZ1fS5X
dZQ8V3Kw6LAXxee5AkCWOkBIuop45L1LjFwdKYeB9AnLMCU2smkYKPRP1azvIA7s
8D3FujSGmF/Yd9ELxme0CE3SfVsKRSUGOMoaigRFan4QjRgkpWUv/ng7hH64eUUw
Ppy/E89Ikm1r0gTkhELP2eeO2R8ep4YYGeDVsg1TfgvR/H8bZUDpcAK+Qe+rt7qD
73NdCV+nZExyjhsP8DVTJDFihgJVlS0w+sKcx0fjXv5mTH5dw2Heho4CiHx3DPW3
ypz5+Xp/ACHvUhWCZqUMn7lA7TqbO6Id+LJeDt3bchqG9ZbjKGM5Rd4cpdEYgB93
X7TVssA1WZ3IL9TiowrBZ9RyQz4xZf/VT+f3zHNfONv8sfEKTtnHv08KiK9x/WpB
nLPX0o9lzyTpjljUup+HLDSFWVwlx+XxWlzc8EHCFJf2eaOE96f9fz9aKq2NuV9G
ZSVl+SMxdc2eWW6GzOfWJuMyYxWmghDwGK9JmG6rZnHyRWDA28iOwY9ULJxgMHpO
bRgnFpt8Lc7tXLBxzTjbU1GuXGdz5LKaxSUlxF5eoytbcikpjt0VWVLl5YqZf9Vs
SjJsWoGXVqABt6gjE/CkvGdkQc7ypJeabe93jEtfj69HASku2TGtcMRSL/wCE/J+
0wer9zgkX0FdkRA8S3hTuJ6aD5f4gTyzKQVj4F7n/6g+LFnoW1DTOPALK5OtBY/E
mYwANA/BbxMTgxo6v/k1EjvdJB4kIzB3gvwwA2aN8EDgjRF9ABWH/ntRGf9fF/98
/JoJcrOkMgQZuw3GfE//k3aX8jFksSnfDpA3eGjsondEzNzQTJPwCt91AVoSUgR6
HTdVrWL3NkRBP8AdT29Xri3X/Xfwh0Q8QN9psea301Qarzcn3Y/8/w7yd6Tjgdbj
bx/VtVAXVOE224rKxGl0jLPLXVEXZChurFwj4/veP2pu+lySQbRnCls5rKfwQMJm
9QvAxhFY/6sSc4ejPJLFA3cpd48s/D9OaRO29KpqwqFpICEZJodrxdduq2HRXgXy
VcvCq1hDjoghYhgkzCmjN7QqLzC0mDbU3He6Rx8xaB9UE6Rm5ff3ECwZUA3JQXSm
YmpS4WcbpQ5KBIEYNNTYHtjNO/n1fD6p6BFTC6y36orMbnEuFpKO/CMPZB6FjmU2
YJGbx+ouEwXcRNCfHm13NwyX88bICDPraaxgqUvCADdFjEjceCtr3q4QJYnO+JKq
bjWcsxdekCebBN1fBysRsHOiBul6nKKmikfRI0IHtyzWfwrUc0wl5x39+D6UMsHY
LczPaor0lXGZMoL5GkXIEnYKTGv9ET1l0sy64IdXAMIuxT1dcjR8DO40P/xcD3Yf
HiCbpRwNdx0xPClUbVO5tndm30+VVtcMQalHGVDSjhXd25Plzd3jZCiPKOqW3C/8
g5rtsPx2dhov8EN7MXPtxB5ifIA0cbl6F/rV31w7yqStdD1olm898epOlIYjiaTi
zxgGBiNlhu3/3icn1wikxCHMjV+vULw0mJACsQU8t8zBnTT10KBzBWduA+/zbycF
UDA55FdzNB0wXJYjxfP7RdgRb2rTJ2gncgB2xQ5WXRmefp7OyG3ulXl/xCMWU/fJ
mjALKp57MshTNUYkwJjfwW72k/nhmjWZXlH4c97W+aMxpfUipEckwC56lej1KDYY
W+JV1AXvd5Syg5tG39CYQsVFc22YrKwclO+lZNOFDMNfW0Y6wxv0QUbERzM2gwn+
zhw/juzgpI+5+reKB7IiwTf5PEFIBzbr7pFHrAC1aPbsdkZroHW+jbOiMCqcsOd8
cI6UDiMFI6Ts4eVF3X9KKX6MfF7ydWd7JYTm1G/r438KXa3CR/o9AUVcWoeuLZzy
RjETXAlC6IejObjXWl1pAWyE1tDCL9c+Cf/EHXLAt8tK7IY5Sk/iubRtnKJRH4RN
8ILkb698Y05MGxJ5g/NyEQ5Sy4hvbaSjXV6HyIwP3L2liv2BABj+qmRQPZB+0AN+
/uKebfNeKIS/l3BhVgHWAFt2Jhd4J7Ek7OC3egg1P5lKtSx1hStQrGE04mhGnEzZ
LLwfqju4N2iXgELAgwZ/PJBCS51GGjfKBU7XvNVJtiWbhSKzmVxuEMXm9GDJhSC2
jF7MiI7TWhFKalFC1NR/M0hEgSW5AYkL/XwowULb7V9HfBLzM2bfv+39nYk0KnCh
AsJ+y75gQ65VdAGnMRW6t8KG05ZBDy5zndWGwJa2vUvmoCX7TG64EyRCDszWwxID
i76/nPlTeCDyZgu1HLSW7jTNqkdAgft+oydGtDSbPcLe8CPXAgGEq3H6hsonkczp
erzT50eJxoH8r8CbxNjRNJx3m3g74jGiaxcADcKrFz68hyKU3CNr6Dk6FDPQ5yME
LJdqpjULi5M2ALxM2x0x+ETnB2vKtfOkTZiFy2JgJC2oW3WcqN7P501e0SddgZX0
gVdRMPMGPRnDE3BiM3BP9DmmfS4Cvfw2eVugFmkF8IsAiCgm6EojEtxcAM7ZKr8a
kCRsgxIMkfJuI/gyRkDfiE9dyaPYRyDVM2FCYzYRgFA4GocShdaP86z8RTCPgB0o
dvXpSkqidLn1TGE5W0jIWE2LsGWQmwA6KrdDRrUViUx53CUpTFDFF7raXd9ODtGh
L8D0kVBsZWxEMqJk2DZvXjIMmLetBmd8COMEqZYdYttyvzgzx/UdlF/Jt7lTXXGn
T9h5fLlmiwmoYF63ftb21jjomRqHlwcQ4AhQ2nbkj1NtfGvPxjc+zIlOI9ao4Pcz
1zqhbzI3Xh1P4TgvMOZC/HLk0f4kTnL3qXM5xisRWSdigoDO/9l5ny9ASmzWzMpQ
7VadzOzbu65Vd3u7wvNKC4tUwWzltBJrHst76zSfBrJekhGOWoz0giXf4SWydBAv
mbb3YoyNZlkQf8z6vt2s+v419pDg80K9JI1jaUc6klC/PTIKAJq4Y5ysWSUwzwhb
UFerPw2zyslYZRjvt0R+Lwz778ER1rruBICQ2Mw1nSyplKT1mycvJbn+nu16xloV
TX3P9oEP/MM67DD9AO6tqOlLP+2a394q+nC2Fwf7AaiZTgteg6QGr3+qSlZHHxAP
BIHW4eKUf44sNeboWTAUYJ88v0qfYuvPR6VJi7lJ9IIMnnLUgSWxUwHMwbfcn5JC
hIY0xyLNIEJysUMHdVgfjroWbBZSJ5Gt8YdzyYcJv0kvF9RELJA7Zhba0Rqpjmzu
cczEiXGSiUXKRL6+DBKk3Noz+18QyhqZUvtQ/SD5d+X6deqbaLTU00d+i3Iw96Si
9gj0Xe53vNOGbd3uiqWhWmEkVQ8RRggXceZ6vb7iA2BockjXRPF0M0iYyqsQ+FW0
QvYLbnVpApCOFcVMGyhWo3hxleanuBjl2aWxTmkdBuz9t8flSpTKpDSgPVGvUolP
EuSQTcDtKV1ZAfhsb/2GwVErJN7y4kGxBgIrYuhUtjeU/AlaoSVrUc81C9jV7sLQ
QHpAdlGVEJ+zlIyJJ6twbPODzHEAMKxYqidbMGhmDUZJ4wkqqWQwiXh79iqLYRuW
XcrtnHVVeq7IjzY8p8KAOTKnX+037MBmoNFY8WrDRLQHWktKo/3hogBJoxbVfITL
fHriwxNaPi3N3DBNp+p+KJ/BZHrfv5z1K23kpNoWOJ95oyf91OGyjgVgTZ/bIECb
TeUmTlONCHmotGzbOGnZ/OUENjQMrm/UBCg/PzRgCryf30BVlS84WkVeTYiNtBIp
xnOMMRoXtUoCU5f0MTPFUwtsN9jPPv7xdshkHJjPESFyZ16s2OwClcqTZl1cx6Iv
fFGLlvySCkRaE1xOz2P942t6JLbegS/M11EnpeQmqBAktsXXnYMFJyeLnqkTbe5Z
ilOT0VlX04A+sMdHBkTQWZtf+pQ50lxIBOvo59MaqIVwgL574cpYpRA+ILCSyKVk
oFQIcVJ03suEtmeHqf2I9nkmNxU35gfgsdFkjJYkr88Ul9aWt75BO8kOAph9pYS5
a3R2cCwd7CwHI3R+dpRSC8U6kFT2Yqs3iwrzYk0kF5dCIQUBdoL90JUsLd4yYpP9
AFOC0KpxBIOBdSq5HyZ2mjolDHwb4ZiP1CMQw9FAPNXXIAUXp5//w0eqbaGKLrjc
YY7q8kOA/keVkM5HApZt0NbnR4yewK9fOMgrWkZopVEiQy6BOvGQ8+gUbmA67BGu
68fAto8h+GCattY4YstFfkZ7mnNlRcV4t6q1RjPm3uRFV1W8d06/SuMbV2YeL/RZ
6SKIOOxsko5eiJEOFXZWVKFDMb2R4nK4Yt2c85S2ROK9LWtoRy/0S1faadVPyiVq
WRFWK0VqSmSbAdzLF93fkk3SP7C7z8/Cg9tsUa6ZZBx9g5PZs/iPaXfQ/hHnXi1b
QL8/H66TFtVQ6xQnLJz/OqSfvpn95p2T9SQN2pLvPPp7dSZJgbieH9CDvGzjIuMg
BYfDBP+oXrwQqEfyIfWPi5CPYJXGTxNn4bLjfgsC/ADrgEX31w5kZ7miKrg0vCon
pNAXY48cYU0iqb2G43mws9toFMKb5isNru0M11W1J8Ec3+Pb3QgBpvL7yjblm9qq
/i1gCmxjml1P+7AgJTQ0ndM3DdzMrA+XVJCK4E7XpvL7iAFVKJ/2qmSSbr7fANYX
qPzxBcAUEY1Bge36sqr1BRjHPXL6jNXJPtW4MXqhPJSY6ZynCp1wVL1RNilFhhuH
M8aQpNNDISAhEx+S0RmLftpkzANYSOSlXbVJ3MVDekqiOG4Q4vUUtM0WFXMmkjhj
Rff+iLVe3hzg7F+/8ZqfQ9nsW7GosjrdLFdujKWJfSX0fiSVQMSeoS6fhCYqO0Yd
La+4T6oMuv4vuQTaUsjlMetLZz7R99my3pbkpzgqz1yYULg9kVzQ60TPsz1oyO0F
3jU6Tt3KIMXrtU28AVW+Ga0At8i0XXy/QkGiOXRrbHOwtUceyEJvcO5lVNnBus/y
GGo72hhh9eNvjfpLlIo8Hv4ycoqtUCGRDVuaw//dGn/3PfA1bfmAc8DOSNRuc6w8
32mxT3btx/lGqx4YNQGrwIV58HAhr+BtisV13mYqUHSOGAZPGJzEfsymg2zvT9nW
irOB3o2qQN+DfhzgoVwHLIZL/8Rp8isORyp6Lnk+5vZhF37g+8S95R9I80McLqAO
op6CzOnkHXggYkTFdp0BtBiGVWI5ZzHvspZxn2jG34jr3fYClbl4zW67n89TIDbb
+DTpHPW+pZOGdVC3nZmfwFIEzCspcGswlzOBnirJG5kwcrMhwOXbYFZC+9mpGR89
CJVsG7b/bD4Ah82P+fk6/sewJffM1mYAHCs2O0lyh6xFIAPkOnXI2KZ9XEFXMVAB
VWpaU1kEbLBEAcz4YC7R5bo/j/zzZQjiaL9YyUvTxsuV9GcSC0rkVihdwDZDW1n+
gRl2jx8KU+mf2nTcb4EJFrEmStQZQdRMlJk73wPM2yd8VeKExzuPaXl4Ooh820V+
DgakF6SqJjq+42Gerxpz6D3EgQpCszlXRGHV+UxY2ALuazbz2OyTeBq3wClXiIW3
97WzgN9KB7G2E3wiYgwqFPxk63Idxsp0czs2YaJKBmOO8MD5XLBQiBm5GBKaF/+U
SpQWmVIb+dlgZ2mHKUg0dSeCj5x5IL/VarV2x/zoo4f5aQGpFZbJhzLtze00m3BN
TFyQNaidSmlvxeZKMho5KiRoHXCocc+RZ5MRzw3D5NE8Vm/3w8ZexVMStqV34FGq
QYQL326BJurG6BrQAasiWeM5QCvSSSUdIbvzsC9DUycE4f+NIRXQgqfMtHkRwvC+
MXABvt4JRVBNy86IBQ2FOdO0wYs9Xr/fgobKJ6JAulaS0yiBHHuUvUPfxoTQ8HdR
XlPE/2iG+wdtq6dRU7q0IZzTZ1GHdcOJcUPuenKcRGyoFpp0w0N+wjp+IsijKP9W
zKRt+t7MDMDFQ5KT9KTN6d4joEG4NOOcBE7dzKm/6f+1OcfLbG+b173AOgjtg3T9
I9J3pIFzuan8mkt/XH1zyP3itu35ERe0kgm1mgLflmRrS+Ez2Tz2oHC06h0zr5Ko
1Vvp4oqmqSdMjDLEIlZKZPrZVa7s4xkm5qAYFTef3gDvudp6x5i5xoeznYJqm9yw
R1QxtZNcPX8axj3C8tJxuZ3wpx8h3YaOAjTL5W+264zcOgOURQS67SJf0QvcB698
D+JYOjLP7FYmMkuE1652nLGkZMWI6muam/fNP9zXk/JTrsS22s5U6ekyvVkN8sak
bBkd4nWYDCLYM0VQPsuHy+RB7x1fuaj6WOLw+VWssVF1QtFPzI3xiZvaL6e7s3jn
CtKxPuTe3lP91YHOiTJA1IJmxF0cFWYMD7kSMTgdacfqsgU6dwF6JVRw/mQ9158v
KlM4oE9gDU/1aZjXHdXU/E8e6twmcUPJIRT8ynpwizDQvoncTUJpqMfN339ljcTs
Wt9NnCPt2GQSR4mmSmpcttoQRflJOxKYYjnfziOizhRTqDHG2cEhm+jc68gReB55
Zq589EIeNuOe+biphXnMKWDDCstpyPnknCB6w0XH5fcEXhNCgnk4PMjgEqpR8jzN
/UfngRD9pImaDkDq0RnEr9Z0SGtEDpz1xwhKPs0tZOJGaOltYHlULpN/YyFkds9Z
XSNGjgOmEDArcDscsYeIKrAVodpQAMonaCVKBGH4LiSDVVjYr94xOUiOOrLQl74t
yGz8zo66OIHhlITdtiWRns5QPKYrBFl1KzbBpjh1bjEnuMT0/APolODEjczdRYx/
M4cUxBR2OYWRkqb+0nRQvAl7YjrIg88pTdZQTLe5VsVizuoKTBVaGofptRdsrTvf
UnhZF2QHoc91+g3b18/pO498GLomR60L/m2b0YruIsEY4UUtMrYchgSnslgfA41J
yXwWXrtETK37El7o+6ia7jm0yDypwKTKFJ7nEg1w+9QymPsPRhjjOtrKs5sKRT9C
9zFL8bfjQ6AdAFILqyQBabS7L0C2Qif4TRWDaIdTe+wlCbkHiGwEyEptiQ//cfdv
p1/TPykiky0ZTFRuz1swQ2p88Gf5oJYV55tWcIaKJHdzJaS8BS/nNxrNfPJmXOXx
ClqLyAN/Q8BeR3nvH+NlF2t91vu5VZPG/GZFnH12IcUR+brwFIRNYh/FsElko1CR
L+cWFbklASKCg2QOSj4X1SkIRNL8V/K9etWwoY51yGo5RbRdgN4Pwrz/7OQWpT+y
/x2noF+cPFbUQWsENH3hwrYqLvUrlxpyHm/D9DPFquloJu3BGlJGjpu9L1QAvM2e
98hlEqY5IhXwdPtuITdFvbS53f23ZaKRinUOPXOzRe6D3P3mAbXb3Li7H/+IQki3
Tjh4AzsiNqa0k4Ay20gIyDhpsVSJb99N1/x6EHLAjDEdjZnFiTPOdu2NcCPMZHOH
WY5mhq19JVqq/pKPREK2GwJ91195fZcyMo2eAaj7t17Bf+GsQ+iwWL372QQK9S5a
/flaBldG3ihX1cJXhjbnYoUvLykYoOKPXDkC1sXwVHDFMz08jMZQIBASMjK1rFhh
KzULGdb8mFM0gheV00eOJ3HxqVJFtZU7b3VMPEiJxbhimbGv4Z8JahflIIo6KInZ
NBkl4hKGBcL1CEYX+Thin/+LagOxn/luZ7o1FYdncaL1G2h/zbt9/I13XXV5PN/g
VK4/s3dML05GO6upY0VLAi39Pma21rKpj3L0QljVhpwU6z2ml5ZC8xbpMp601miT
3eYKAYeE/3yrNBfW+s+yuPRVgDodD8+s6FEDnMgNyt/sa2gVYSHxfHVTW51rm9oC
5z7xSouua/cCFoCp/yjFC/AQqrs+AD0QmdDnTqqzYY7fJrMfLdzZfYHFPXxHHNpD
JcYCtNUNA6zYBGZll3F2vcYyymCJiH0f9uPol0OxLfATugqUDowRmTw+N3qJJkUb
4eCyAKKI907A6TUPiuevnl8Q8fjqJHuj9bYccWFDkuHwuqS3abg219tikzVB41LF
UlemUb8uL1n5F3vebDFXOUwAnvJj8ee0S1KEAug4JUPD6JK0jcatfyJsOYHIOSN7
J2GLSVk+Lmb2iUufT0ZxheZwU1pks1PjYfU9vbisO2JBWcavhWEmGqJa9bG/xvaw
wb6fPDSsv66haWXynW7TkKfB25nWcIiN5edrilluFkW/zOYp6oa4ImqUZTnYKono
KSYRHGZ1fRnfWWVcmsGv9O2fblMZ9qcwb9x8/5stEqAJ+A1/VbRSTx59eTlZztR5
rc9vRKj4+dDCtXGVUXUsvelGai9m1jI3+MVPcfeEveYDvCo1zg42/nIL1D0gSY9b
LtUajjNO9g35G2Fcvi4mZ+nJHbzlEvv20WMFQSGp+28UTnkGZhLTuonydKlmLNPY
msrgD2AV+ZUpWzdRTD5kD7pu/zdoKbbSIp63EsoiSDOjNuLEzYET22tMMG9vexYl
05Nf/Wy2L2cFCRhPhPIvCNVMrDqyVlg4hvTjAeg4xGdGJkntOeKeoKAn7qgk/Mpt
JgG0LFj2cAcCiPdgQW1BpS50h++qEVzeZ6EkhSuJ8DRG/uXFd8srA1eMknF6l7l9
4xy4fWenuHe2lEgUUZhuav1N3ooCR355LgFiYbntpnwpaeAlknTiZFuaabhkVMAf
aTT2p/a1p+UQz7V4eu6WMTQO2DUgMFpHjTwPViwS6aMTtYbnTi5pm/fvUZEy5+0I
JGgZjz9b1WXraBbw8tkrnuPPM1ABnEk8SvuAUgDba9J0MIVi+JD33YciGDzpeNzc
HO27xuRhb22OwPGYX4dCXuf5HNimcjNq7QoQX/KbK7dUcR++bwuAD/h8AQS1e9dV
G+r+TuED3g3t4KgOVLPRGKtmb8wRJFhG91mCe2oKribj6e0ETSrcIv3tVVz6tVEM
7++AnWwc4uwuAhikJZFZS5eiUf3uYwl9kXA4GZW9hdRJYbFJXsbtJ+IXhRA/mRGi
fhxshMYX60V+8Z90Iy7fPvNAFwhnE6GEwmkOn2LCL9aI/LMlQFbrJWODZlnLZ88s
41TPpbaTxULCPNvIy6E1fS8dWAZCqak6if3JAQFJPcT5cC/kUK+8Q73DKutWktKi
SnZI2L/+VdB0k+hGsZqAg+YCLPmXNqHVvY3i/D2GjKbC/6gq7s036HmxDI4XPvpO
TlwxXpBUdZkLluiAIyyUx2MJDTc8YOFEEA9J48HSPTiP2TMbTAPZLdO/58cHdjhu
exVkbgcLU0BbtzCrwuIGNM9R+xrZKpkd5cEnf2a/VmvJiQqZbxynJtr15Yu9VdXp
5HfOcJuTTvslsVEsF/1Uy0ESZ9IGlDg/NDDlxLiPFribfiT7mlpc63eDz3NnYFPW
CmlazmBFJ16GyebvTlVUcdPNyDb7hw9sa0jSP5EXqVDljIBUqavtax737amd+rdW
lwsvhY8SMPDr71nMqh3mIzlgi11SLvPOUiDRjbSz1IAGU9E1XKd93k6XpvIGTpiN
3VXcC0mo7L5jICLd17kb+HuQTSwBCeNYiidJMiiY6xGaFA6F8U/Dta6TxsdZccWf
UhCJpYlV6G7LVDxYVHKw/kLjfXYhTkGRZSZ/e6Y2idgUL+4g0YQc5Zds3tE2wvCB
/RPOePnOewWg6fioK1pOVAOB5RtWVYb/CMJbJ9htNRhC3nTCBYGNpwKjfMVdDOkC
9CM7kRTudmxJAuLBk/6TD4lUIVXcAGT5vvlqFvEoSHaRSHkIq98spKcGfusEvNz5
R/BPjg34vlZ0x8dlM58jpd4c+WfPJ5kfYzdtg6h7oGTyUx012+1aVSQ9i7svf/d/
+UggGoNNAksKt3U3w1y/9VYes87ie2LhgvECNje9+05RtTcO/RSYtgAkCZQ9zqQZ
C1+a7fc4HNL01J79jN8ofSgWH+WuhUFgtdn2d8nnvbJsd3H2Af/9OcKSCHVDQ2aZ
PqqDXQOE8mChR8tx5/+89Tj55x/nrK0wnH0FIhQUzbNS8wzKrnVVGYabV7YHetIs
69rH90MWSiW3ZYc0eHcYLrYq/FZa7RGI5O2wjK9VOzyvws++lKYZvrQJQg2JSaPj
EHPG6iDw8FHcm3fRu8mUkIKsFneZxenyNB/xUlLaWtzpIDiK+d4jUQ5alXBMk6xy
xqDfQVOL6+lDryrSPF2vYcbK3YTgrNQ4dup3IM3Vxw8yBJ/AfpuPYxjlGFw/NNDT
liVWNRqQS074P3/VVAWkwEdBiUZUiXHaAdeMhLnRHoCyj+uMMms4uGLQAzUm/wXS
njL0BvOquvpGYb0NDjlRNwDhZ06N4BQaoC+FImc53fOk7yJEuDxH1iiewlG7qoSW
mP6yXXCxzYiap2cSDrqVYOHhvLjFHC1BlhksLsGQakxf37Y3cEAmiJ+hF8lw8qS+
p1uAp19KTSyJeWj6VWGpeliWUQEnBH4bABtt2nZRQ8AAuBzXqOw62MVgFQba055p
Ezg+hF22CsKJCWptmbXLHy6WC9eOMlBhHpfnJd3BsSZnMGrT3Yq+iR5alI/2FrGr
0c66M4wyxXshXLYbVLwDQPDAvzAEuTDQQRyW9xXcgJ/gUEgObNtyO2ekAb/nZj1h
w8vVVGS19YUyBjta9hUhJk+b8l05LIhuDm8J6WrZDVg4fqunlfBuZFVOHYde09kX
MfN2utBokGChZgeONGWZcrsetJYKAD1OkTsbOf8tqoGqgkQNCMv8v1LJtsximU38
ubRVEj4lOQUpEIL3hppQB9kdlGCxMYKTN4ur6gtzgme0vWJSGRsslN2ndCc1ui2c
QAcDZLWyBIStRQMVICe2mrN8507Fco9jowtl7l2Ey29EA5joOuJx4+nzbm+em83l
s+ewp/zCu8K4F15o/B8zaidVkM4vcjElObeHi3l4DHFqI88/ZoWIdAqTZFGoaPJV
Ecrb8T4N90Qi29on3rI5Ayj5DGYD4eKneW4xFGXOkYGta+1kjIY1HMsazURW4SSR
nFDi4jWzrPHGZjDxBr+PPfIz+OQv+Y8lEiOhCuYzvRzRW3VhXt+N90NTeweDK1oj
5I4eo+rwhJS4XZxOBfGOv7xcSju0gkgB0Da8OJkpT02ev6PWJV5+002ljcDBAFFU
zSzHr8qa5OqK5XMLlWWJtuW/WSrjVtr7H1VxTT+T4zY+o95EBj2RrocP2H8snxwh
bbXXtbfrfAo0Mzhb00IhumON6QmyqI1YYEedIDHosc4poXBTNeFh1VAI/JfWd6Zm
IIDWYSm4qtpcyCXUVAiMVvYf4tSHk8/Nvk+I9T+3Au5QP91yWh/2K2O6cOpGejEC
wLXM25HtKPHHz3G8xtacrUVUIbPW5hwqRiZXF+CbKghB7vTjMMTmrBkL832Dunev
lj4C9+HNxXrZy9I3fa1lZ3rR+a0B7Zy8hH6aLNXSil8l+vdgtGFXdTzVKT+LNkue
LsFAw8U3JtksB2gSiLxPnpLCFOk6QDwZzzYdQSpRpMm+z24ODKMc+xjI/SGY4Oe+
KViDCXz58gfGO3qWj/czvrHyF4HYlKwEgxheOEEwk2GN2Ay+5XLMTMtGUpdBAa2j
VnKNVcpl8m8TVoW9UEUJH81qKOL8zXgmFPOi+4U/20b3CImrb8rd/TEfi8+CcW7j
HwJo42aCJhmY/SCT68k/QrpxsHkA8nCKSSFnIwvCmEEDnVmSOKalRVXPRr7mIMzd
RhsLOt6CuJ47ipWmz6m/6/I0TwFA6hn/WKFoJVCvnBNIYnv02Fa9n4K1lEdKT+Mj
eXcpudPLSCNYQOTzzb5zaEtJTQKw6kR7BLbfIHC1S1GrHUTeS8fCXsjtPCEGPp14
TiMOZnJOZzYCdzd2NFQjieFpDn+x/UIxMLJlIUtJx+8FBphowLEvqSjfqL54Cfs/
cK7uoMNXiwCWZ4uWLYYyZ2vTH8vVOX6+XLw4fqTMQm8py+WFLXPj7P6EsuYxC8gA
AvlyLO1h2yPieeB/6v/YuR9RUSxMK2rGQYmQs/0Hfirm143ssGrf38H5k3Iq7AZz
Syuib+TKzfuWIxg5h/LAWp0flb2jUL88b2QHdtJd+rD4QNk1BDrDKU4VMYpikOW6
S7M0rliXwlGWCpNSXxIXdcllmNCb+0S4rdbLYiPVnwl+hAYcI8sgJJOi4NGLg9OL
GSMzH3Dfq4hRORZZELHdPy+GqwzpmQQWniQbHDs2JBv7s0ylRgDAzJolR2wPANB7
cjIVNxriQR2/AWOnl/brjfljEGeQO9+/B/itKbnBN+r0PY/BdAlZuphoVhtGSHli
VL4OtiwndxZTjC1fCpeLPj6u9jpIvsSxKxInIRAMaiwj16L2nP5fSbQFME8AyhHl
g49M2dRm1nqNBqmAuOz+M3yxOwCFcgeihWMYorhnzchKV+cHxNvTQgB8cPFJ1AUl
A+Pb8zkMVDs9V/lQRql4uHWhkTswILpgZ7zclAbfSnfe8go+JZz4PEBzQxc4Fmam
u8D96l313fC8PsGgfjxYkkmc3Ta0s68PgRZ262t+NHskO5hzPS1GaXa7xOXQvfuJ
ACZ5k87TpSUP0ovwn2dQbdYiqip/GZUUYgxnboD7aNcWdnSNyIJnR5KuJnx/XvUx
NrDf7CM7RSEykNZcS5uoeiJTkmK34pqlCFd2tWJTeBYe4BMT+ILljHOXvdjL2ga2
d7oEgLJ2PVIdNBY7OMrCxY7CjIPKP0TnYwnzJi005fBywtgffYVhfTWx4XUnU20+
ywmF0T3n81VgHDUkKw8Doo61jbENF9hC4479UyZD0sJvEESt0y6XI88ggmKihDrO
4M+PEJoN6fLbETyA3/KR4y37kXjyCMa2n0hXeKodo03+ucRy0QdWIul+yWQyUwFk
XPdKdfHgsBhV+KI7XtNTmWM30pKkQwV8YvFR8PjqHCBgiUjBAST/tHdC3DVUBY23
prsrEUGs3OdjVIAoV6QYs9FeYcPNf0OV77e6pPjzG/meXdHfLpfCm6EulJeXKYtG
lHWpvZrnOEFtmEbFSw7gtnbWGSzdE7BpuGVbbwSFAdwMpmg9kleU+qauD6Wrp9xh
j2F2GtP98f+DZ7u4eKExM+Uoq+R4GNa+LxtMtq1baWte64hmUh82gKzbY0GveVDl
QMc4mT1G23k5vNntYe23kvuN7oXk2OlYxYoimdq3LcQxKG3hV+R47f57U335epso
f1KWmkoXHoe+PTAgX676s5ePNtjFg108rWGTDUx7RqTnmHg5zVlTdRe/Z03G7owT
uKfXN4xFU71KaBEHe5fzZv07ykpOroZxtcn0ehBIyl66ZD7vSZ83rs/3Fboz8b0J
l+K4waeUllFy7etrd6pLG8cXrJvQu6EGuv48k4pXdjvW50pQPTOWPshguOb8o1FB
6d35pQDYWqNwBVLTGqyrxOiFL6S92u0pUnDnsseUQ8jXR+TiH2NgT7/cdjdB9MKS
eMSa4wx09GF+XYTSMPz4lQS5refzuKqZoXcjeVtRQralLMap9njk+vlRjVu05yoP
1AccHWNCmV1EFpEL5JJJ8KtzDdLgWNpRkibim+sKYmc0gGRbv7N1OFWpCb5ieEVV
fkft4wJY5i/zNYbSUoOT4Zt8+mR1zyQpdu3b6QBOU4jjl/XjZXUzmYVLn2B8+mOp
HpbajDgagZT+KCn4lKc2i1hYrQAddeNxJL3aF8VS2u2zPy6AE6DURB9ytMFMtQ06
3Lr3PfCMjDqn/ZuKTjg3jn0Tk1gcMPPibmWcTOhOnCRYmYZLVVSEHZQQYoZQqa9S
AW89Nnfnk3fAt9RvQbDBDAKS/xRaH9NeMeTM5dgX7ci3t6EnT6aYa5wQcHh42Jv+
OFI/D9qdCrvNZk4TrncyFexv6uZK4tw3XiqZtla25zsvMsG94uXGsXC+2o1XFcuR
U79+Ji2wubA6EZ4K893Eob30nuBVDUtbdrXd2/Rn7Zd3xs/S8eiLY8MjNT0HtsbH
0RCF/QB1VEfte2PAEObDaEtgPnpa6DeVA2zV67CsaeiRwKqaSwzrySIDuz3H6nQU
i2BOCv4hovljTzO6W+sI32TSw9Twh7TBhlxAt6jivnfjC6TCrUhyc/SVepDlnLav
SzNyA23Ivq/JhjEZeyIJAAHLFozccNCXjfQAdv8MjzEZWPfn56UiV6WkRvR10rhz
GbhQdTxdB1xrAhL0q3GoO2hn+z2AhTzUSLMQACEiaz2VgcfqoGoi2NX2yqgkzYjf
fkR+OYe0LC1WPVDiWVRY1L5ytdugqMa3efMYaM4vM6WsoPS/uPcBYTKyboLpjYm/
/YDei5ojIF+c2DATxrSQr9noNpDMJqOHuMTIoOkYDOt8kgam0+GeR43X/nlLDJ7l
deonIt3DNWJPA2XyRQxDprzMjf8l/o1ZuYVIMHZfgkx+XrLRMdQscB1FhvIhJQIw
0chmFUVZ6Lgjx/d1QOXgPeSezifdz4KKaQjOLo0m3weOaMJaGJEzuF08uGvNU2MB
jpYoAs5a1mcidlXUdsxYic2TP6bcV5AuhvN94nVbSVGBk3VvJp+3gBvQUvekhJpu
0EPjwyXChIznSzvVvH193WWBItHSTx3Z3DZ53zq9qXX07z1JzY9FB0iKpl0Rcefm
AqjHjH0FmhPLTjn9wK0Of+VM3drEU1gsbw8D8YzZvASQJ+hKhQ5pTc+IArm6oyTZ
X4VczbBSX4LWqBqln6uI5I+QWwPDyXC29DjkCkF8RX18cUSKgzFNp9tqP2lHbXlF
YcbcqTIeNsLSVZlPvTksPSlJxTsfxBBQW/NqvKCeA3bIH0PwOXsqGzUOogfID0MH
Uc/Evw2B6rydF02h+t8oHXUMT0RZRGB1/BiOCh3fPjHOWhMEj+6GCoNKg2sWCBZ5
gOHQnqFCJotCtJk/XMf6YJj7DwDzs8rxfCHni/u31f+9WQ7VENJ05+AZUO/2oKy/
5qVByzgLC0ik9jq61odh354zuH+xXvUmajfDTDPUvoyW2RHegy9cPAzpvZxWAzNc
ZzRbvgfg9XvDXwh8L4IrNZFulQGkxFoIeNrZtFRLKBbd8A+EzcIrNGLU1ntdJdL4
AuioP8epePURVRaMP9b/lJOvSFHy5EwClAg2AXWxlREC6dz4dUxYbzTxpbYlFFUJ
6b+ND6VCpZfNB+vfxvj3BTaHeXPFLS85Cu5hiL3OGHq1n4d+wYed+CfJiMrf2y2Y
H123HJY2M3JoyTbI0QYJ5ItOjePvJ1xksnmZsLwjBnIEaOKO/Hp5qqxKzoJC4Q32
DsqcYKNWqe4sZU+1eDVH1GF2RfSgf1K7vKNFnyBN2ebzyovvAqSe33PA0VXA+R3R
JoiDZjqdacSIh4VUmh6aS8nlPfLbPZZVd9wYNWaoonoL6n4pnoR/ThPzH+qYZY95
MtPpNe1cSDBdQJpKA3mdJgipII/1VPxyGKQCfuVZoVaxDx1il3VuRMTNrFN9MFwk
Q5iBjXNgLewJJlWcft67SoxR4nq8e0/z7xC3dtg6Iu9Sc+EMGbozdgRQp7lf0Wse
v6bVL+eZ20px+tPpofml6tgavoQNEHUdvUTqnjzuAXrGssh2pxNNK1GDp8xUBzqC
TCP4f0YhoSggOAG6plsjiF7P9QSSU7lbqC7Cy5mCocSWisvAhm37vYHUoUm90uB9
DYwbz6qC8WCYRrKjh+fc6LqBNKWg+9VX2XBpu0sov2cA+MowL7LfiuiLz+fm7RNG
gx8EprZH5gKvKEqedGl/ireQGHVbvcMgb6wcEXfFeP2GyhAkLhAXYum2zPscHCeF
VXT8CVU+6Dkoc8JJjBS/ms04CkX6LiSFm16S+7e3DFEdd0tULoKKCn/8jreQ2XNk
DBDLwGikvQBHlvy5/+cSP1Nmna2p+WZS5po2l1vLsmh0mxcgVYsulgIx5Kw8fYkJ
5dlfHARNlzNtsFLbwP4x+Hl3lpf37VKMsH6Y26CpHXlfzpc3d/ILLz/6T+JVl1tE
bw5fPYqo2hoNxvs5C6jzI7ZnU5dNJUh+MoHK4Eg+vN21VWgYv5LlOMdzy1qSXHq2
UOiUwCaQOvin6F7/XepfpseJVOPoMuk8n4NWeZFgiZqWh/GJ+sd3bA/5c6RnyBId
bbfYFlbD4QRUjubNae9fRkQWkhu3SPojUr3+QxxIRxKDX2Y2KTT0hyOvi05rMlw8
5ntxMGQ5n53BXVRN2vRvqpXSVOxAELM6grxgUpntKpM2lHcIkon/4xdUQtkHPAcz
4+gqBdDmzybkxxpjvUvnTFL6VLD96F1LhwfdaFd3HUOIxM/0b/IGT4h68jQrQqwL
emOiKCdIxdMYCa5qzOPgwoFBjZ8kF1X3aVb342UJDbh++9EtdGAOU/WnUEoBPfSL
z8f/4mYFQ+gTiF70SXE1CwUkGITBxAGoH3FOK8AV7b3MvQ+Jq0BHr1ihZEudd4Tz
10AR6lH9plFZ3JHmveDn695p8VKV9Boq8IgJAMF1AMMnHtqpTbLWmSd3rSiLmpz1
IZorx/7qRB/75jtBG1aaVXj1fD6Bpa6kVHgrd4u/+kufHgaGIPJzkoV+SmZ0KTUp
i7s7sPuziAaukN4y8AfVPZwFJIUkHKudiQPCNlKzVnjyr1eZtEYlHZzYJ5KkCW5P
S8XSdGXt7UJRs1tEXovMQy0uU6KNFdD+srbGf4xJ+ekcDqs5Z+sdls1pq4CNIhnJ
w/Wo0a6pc14mvb/74CE7/gYJKpYd7IJsmbg+xZgFRLtcRvG9iqug+Ig1WoQhebfJ
zg1iFtWWjURwEV964xjlZj8FOt6xC3YJOFJ1i0lTpI6iUmXVWIeJZBN0l89aUhbU
jVabCdsIrku6SErHwma0soln0p5+P/+NYQ1grr/StGxjqXDLoD13b105PBqlzDKG
/rRCs14lDtiB+O8V4PqXpBoyrTN65cF3a2rxQJBEpdMUjADg9lqyoiqw0z8RZ1rN
HAJUBkof/VqmLmvAGkvUQLD2NEbZMa8L1rUWzmvuyS0W4UxsqUFcw9ZKXApYRf7U
2IIV7PXMO0NTXS81oAvyUOvwkHM9N+fYB+EXganTmvg9e2ISNpbzqAqCtzeRgZeZ
JV/cnwQDXq+5lVWP8hjZjVDKvb+aFxHmVR271CUSTfyiqJ2EBEbUTeSOghTPbuJw
KXd9oVi4V0FNvTUEUCzwG1a1O5PPq3tew4Vmv5sIMG0uOXEC3movPbkrbrsQEFtn
uXTNUR1F5rii0yT+hFandVpmUHqH7hHbAqdd+ZSIAYWe8BUKEZJpd8ydFdP8Fakw
HS/Mc2InnG7D4swlvfRXYVybudYqZ3bNOppIdT5Axnq1SzfzI7soahHuxTjGYaQ3
yJgCpQQqvY3Xe6GvsIbuz/CKJqI3ZD8xqlJSPdvfJWH8Ip57IOId1ytDmcHtSiC9
HCFJGL17fdFDJxZV0S7au3Ebe6ksUJFBOGdkjmmJApiykF0g634tvZ7YAtuEppZF
8z5JsUganPxR3LQJnloFSZa9b7LuTOFLH1oZPbqJmMBe8QCNmkKW+PfRWMYDSOaK
UzpEBXttk+KOgW8AUDVVrb1AKly3iWup3PrJCbLHgGL8YG4kqXO5kDjMWbUSE88d
ZjR1Eeu1M1qQ2/itmewx6gH4x9hVhUiH221xAqiV29rzPWhSM55OiVsZ1gfvdpuD
0iYJxtinAr7y/q4mENG60RKOY/8urPCJm5Y+vpATkPrh4BIJX+apGrsQZ38/FSP+
R3vqkFbydCHH1fEUv61t3dwkAKX0ygd5uH1Xq4t6cOjHm4/0plhdD0QVIsVO6SjC
kXM+NDzlZURQMiAXJomsVPTmLUXjbQBT/IOB15uubmp3mqw0RXDjyq0zvhfZttjB
SSr5PfWnSfHXh3BgoJe4Q3xRCl+dwzd3nVqCMb349t87buIAhQDSL0TYFPZaAbmJ
4qpd4Js5u3tqLTZrUM5Eyfc70PDpfWpuHnV2HIdk3atFTpUOp+w31WJ6LdQDyabT
L4FJ9IXcEHBvCSOU9Q5GjrIEL54hZcydtQjZoCD4XNAfFENkLEjYOlbFh1HEgKlK
ysZPtUuvHfFU1Z8NunXwZ/XX+wY3Fs+QIwMf+wT41Ht0ffugZjyr92v1Wg9Fnu8R
RxCp/h3UrD94ksJ6snXTAuxGlJi5ToNAE4y/dFbqMmI/sBeBu2VEAvAJhhHd5pKo
Zl3Wc2wyeR6Y8WXGJ4eMMy0tf54eT6Q/k1DGpKqKHpenrJ9La1vfijoKNMPO5lKS
cqIymDLVQOk9AFJS+z+HuaMQXMLjP1mzez/h67X+9ovDdVwz4C9bdlvG/dXTiORt
1IwSEs57553UJPprnF+W7FQ62+Z1J8zucDee7zPbe3Peqg/+qxlnwrVvLnQUqlNq
yyK7yR4vh5h7zpDG4jcouFGZ6rJtusBMGNxZDnJWg0dSKHve4cSFxlz0Y+WJpjz6
jSMr8VE2FOMD6QYl7REcjyloLZjcqIJ4tWizrpLElPYDwLnKuDsocwP13e8H8UI6
Tj7pkIIItLs6zLsffxifi5Hk3jzYvHkmUv5Mu11andi3/1KcwBPyog4s4ds+Rziq
BaJVGGLPA3JvApHKMazi9P/QIoTh1rBqnOUuUReGrWT2sxuz53oijsUYB1F4fqgY
KcJr7er5NhLLNowIEpOCkzXvX6Jwseyci3OpZcQGxJdhxmGxGd5zlUFaIGPIO4+n
48TMNezB9n3uIuFIe3p0zJzbCTRFbT+xkjkgZrk6K7TSTu4xHh1ROnxy/uVG6BIA
FR2J8oe3yGB+xNx0YoZ/NAEYmoL9ZXxsSy1YAvsM9JBWf0PMSY4aCiqrNklecRxt
rlmbS27d1ImzVyfNDP8pItROlFwrJgZz5Y3odFGHI/Ii1fPCFSfMdgvq5yhPFPdC
thmiwC1GTOE79zRLk4U0WGKujAEgBzm7NC+KNXgGYIoWdjsRJuNEVRxYjOpLo7Fr
zaiUC5ZqXVCaDzNt1pSYTiNiDGfU01JSPv8m4HeFTiuALWCS6vG2drDWAiV6hJLN
Mx7rXUnkUDGK9M7HcTEgQ7CtdIYP1b7pBo6zuldrnVF/HyUDnFM6qGpfqLpKR1uf
YUfnYp666qZ3nVx83zF/x08F4GU1tAHhUXWg7Ps32biHHbJbzgUWzWX5v05Q0lEq
PRUxIbC8wVdSDXQtkJtIkYdPsJ2ZkqYyG8UX3K6ZXNrh+wV4DVNJWKJwcmdY12G5
aHn1Nnav22n58axigzaPG47TEUqJoEg0cANJls5u4+1RBMHeWsPJj3MUspN4xK/g
bvjcDhvCOHoiVgZF11Slql5zNoZgf8CQ/cFqdsN62qzKrNs0kbnLrkgtVP9CAOtl
itHxL+6oOXTOkBI0HwaLX8R+xNIE8HjtADKyMB4ZZHDYT9oYzVq7YgWYB2SB8jOR
bXq3Fqx5K1h6jG0NrEBD70Ov1Q4sVlhiiNq1o2X362yBSIQJcIvNoDU5sNwNIt37
nqZWYnqwGS/t7xb4GQnzaLr6CargdoT4EYGfUPR/60cKhxZ4Sv3Frp2JzUxBIXTc
WnWd1cW605UmwUysVsoJKjEaMfOghe791dQ0fe0J4jzgEEZB2s3BzaLpC7OU5ZmQ
v1woQC0miNqHoUcb5foDJ1OhwrZXG92KeLfzoU38u9aBs9srpTAlwUoNzH3GDWRF
Tr7u00PfIwXfBhwy7vPktIF/+Bodj98td4ZyHEz1qVXwunKDBkOPcb4+YyCcQF3s
Ru5o63UUTKX1b4cg1+YSprPo7Vdq2j1Q3sjmgTmc8iQPpHqT5LVkS/FE4Wv0Bt5k
lVQ2n4gHVuKj/wq56xXtr+dfgQJR20KhED3g2QMEWQNzwV+w9Sx6UKu50Vx/tK41
8AJUK9Xy+F2Va01b3g1CKUxwPfjdJtkU6F9oAef+twFa/ufTL9XTWiEPz01TdShR
yQ6bP96kc69312xGJAsH16j51lDADvEzVtnFYQUXvcg27Tv72MnL9yIWLd6Y41PK
hMZW/ptcfUy6+zWKI5AKvo6XN78YSOBJkY8QaiBvXZHxfLjmb8d2TCXCyIqc6hxd
D0VzI34BxkkVgX7GTecfGxUUGq3Frv1EXR+5pu0eaHiA5JdgiDsx+36vWD6npH8B
/v52Xi7PFLU+pbhLAPjXpyfUNn7rBhi3GTUNaVDmMPW4pAildmd1uKV7nrBF9/Mz
Mc5V0RKk79qFNw2hu5ETpvnR4YVQBBPNFD1U4UFrK2JsN5VbU2VfnA8G5L1qhrNM
z2soo4hf+HqEdq95MmscdVf3DDfNIWu/Lvv1Aa78r6jWmHkBu4Lp/f004KnPDdZD
EhZKq0T5nGLwBtBHaHT4e+6r4zNO6bh0m1/DCa0Y4nJmp3uZeDRDOibzCNQ9W088
hH7mYdG7+b7md8A3xRa7NSMEI8Ua/KdjbQTu43+byVNDqPUbrSi1NKt1/BvW5ybG
pt/jMO3mV9shCcxD/z1KiCVnpOAghwH9rPaWhAFsbzRufNv4cFYXmh+R7/8amgVP
0+Y5/BWwABKNQ7zBxS1PNGwUFHYD10KaXGwwI2d6ZfuFOH/fX3P7qp9YzI/V+FYD
TMLtjRa0e6FBHd7dwtbtggdRByJhDCyZk728zjNJC/VzGu8063FAmVBhZmJYWm80
UUxRyu8U/uO2cgQhOQEQft/d4nDBRL72dfgKJERwwMMsGPSzyR3MdGA1bd3VsYWk
mBDrCLQSad67DVCdqh00Mh7pEXe8jdoJxkWDJo3m/ArFcmnBSo9xSWQ39HJEP8xZ
7fP10qlY+g0bFEYlTV9wHgR9SmBscF86MfKIYq5XHGNTvjyhXik8jtIaengurr7c
VpE9sz4Jwj3lFUgW4Z62X6sRuPwSg+kgFFvxU++bDs+m6DDiqjk099MPRSn+e9XF
YiHnC8RT9AweG7Ff7v5D61gsH1NusEolJ88vcCHTqkKV5XfSMCh8y0n68GggjG/1
Hl05ijlETPfd7Izz3VLCbTziCLfzmDOwTWZF9v/MakLAoEAkuAZvMEcR1FYkE3ka
cR6Cx3jZoQ5vNdxmowO7G17aGNO2JAUC+BilXRgpNJhIICqdrVl6wgiVM5HY14Z6
OmDTB4B07ABSxZyxLhD58lWZxzY1XvTOcHh8dLTLcdJSfqHuNr3X+D9OMZgGJL7J
XOThQTFWHQSSWd8gc11a96jn8bBmgEJtkDNnxzBn+D/SMuSlRSuwGEdgQaPWSMwD
4FYistJR0kl8zUYXs1+OwDG2tf5exKMqwiwNkGgWC4/WASr8RDdkxpTqxbgrVvm/
u1sjXJxWyTET6hDPJSGOQJpS8wIIxGZOepDGlTAZDb6NmxoE4plZA9LG5MxakdBV
/gt8Bfy0Em5YK9Qryzrtd/8CoAsGx7DZhWgPKEgmlBTdBw0vP6GyqsgQsuL349C6
dKMKBK/8nhn1jUav8dcV+xaLnRwC4QG0Bb9SKxv8aR+VoDrC8UMZ0hZoceGsm68r
DYAR5oJeLmJFEpCW+bWekbTmH2wAMmKl28AP2aO2pMTqAeVDCuRqazBikT32fq+N
NA1K8BaKtD++caqMtIw1k8f+7GhHMgMPz2UYegA5N9Su9aiJJWC3A0tg9q+n0vvW
lH9a4SGNz4mI2hvfdtzSLcfZCzAzIuFrTUgPsf8mk/a0VLQ4hBU3wCC160haspmI
IjydQi+rr5QVgIUj6eyX84YSi1dtaqsHajsBIoAOI86CpgmLF3oSFNkzAw+ugXzz
V6qcYHshgJTcGunwoqjzdKHL1AS1XUheZYANMF5GOAoZSEplji7n9l2ntLPYw4bR
8FpzgVLv1yHFb657HeXh1iQ9V7ZQ6CkqqAFElp8a/LdjlXARgklM1X9IPw2TaVpB
U3VSY8puSllfMQJFHMm9pl/++SpdIXXl5Sf86RdU6Fb4eBLV0u8gVTKB+qKigIty
PfmnRO47D2Fddz497Ak5n0kvd9Zxwaa/lm8v4dFttmI+S8caIDX+e89bmx83c5lU
rmWgQt3JlrYDmnrzpIBl0/J2omeGtcGq0JEbAyP/y/kMsb4cvHX/PxOeiecIzDXU
Pn/SEcJ8Kv9jW23+ilCo0tvJ3phIQAY/ZIPD0FoZ0TeO+C6XB15Auw7IZoUVqhqq
WQsxVgy7WudD9m/zkXoj/NcudrShMk7Rs5Mae1o+HahlZ58sZSxw287t+eVZDaZj
DS64/oenhqCWFk5Yk+LTSFFNPOMN3+IAHJWJ+RiBbjxLIyt++rqxATtn/cCRmwBq
tmzPrEwoDhY2A8b7lOKCgTFym7kjw/mjfQQLrZHApO/brt87Q/u+VlnJSHTtCtOD
aEroObreN0twGooNOf1kW5SH2D5SswtdYMmBBb4ewwMXBZFAg/fGw5Gz3xfuV357
0ZC3HsXWLD2wlEOnCWBNdISkyIGCamVZzKEq4Uz3Xqv9co7VVZX7muYBTQqujmin
9GxWUlZ7nSPAaVNfsL1xewKH/UFDzou+t/yItNLvgYVcj4pIBJNzLDZUq0JMDFug
xHkIb/P8o/0T+M1nt1grl0UX54qeozN38+WH0vL77TMpDEJzxHUH76O4WsLvdMHZ
YF3lI5qOTK9xZ/dyjAnhd3WnpjimEwYHGFMhkl6xhRwAtnDapb0wsIgFuo9a/v+n
iBaREz087nZhY+tlB8LB+TAgRgjuMi4m9s/1zIpGxviYny32XgOr8kXABuoDgKSA
VqG+OVvkZr2Y2TJyIwT7qVM9ZpWLRiKJp3aQj4yPJkpODfWWIHFbV0T+GFs+FEMg
8oowe6raS6gTntZgLa6Xy9W+6zCIRi7z20Jpr6wOovfEReqIh3Fl0MERXcfP0FKv
T4LoZECAOvHEF2wYFJCFmrx6OYunADNwaeKusUqrS/k2F3Fc2GZO0jtyNKMQhpwm
p3fdoM3zATai6PJf2NAta29cZybRIu2ZEXTLZYQlv2m5T8ddC9I1zE/0SINRabvw
/s+noObWBB7fYBRJugunqY/7jsGpfMpVe5gdIH9Rpli7wR9hTd8oKRvnczIap0JN
wICMteiU2GXqrkj9vjb48JlbuRs++0UxZo7KdI0GGWYjDTNJUMJfks32/mW3n/II
YB6KEcBr5sZ8Smjmwv9EVuB0JSjqnlZr+AkPSMNXvjr2HN4XMNe5hFzYTRUbPjWN
7n3yEcZL+xMNV4oBqe5U9JXcRAFkjpho6EM7/yHqUO71jlaF9wcBIbPwGdqx73Wt
4554JfLxFCnlvj5zorPCKuwOfCms6XfClD2mswLX0w9CBZll0HWNgb4AxYW1zujP
mq8i3O06BCWwj3SWbgnqYbkBblGE0SpKZI3obgP2TkYKukxvmNXQzOBasB78HuY0
VBHaAOB5nb2NJ28AveMxSM3J+nZ8SCirY5Yw7lewyq3NN8Q5iSgKA5H6Mvdb+IQC
Sk0JEuzwuqOD9b4Ac4WLZ5dbCpFy/grMiSTRSxJfgyDrOF+Nnt17vw34Ji83NI2v
BeRC2FrmH25UCRa7XIvkwRz1YUQv0sf128qRSJkZpP5OnKehSgal/hP36b1lsKFY
leYcXDp4nc5lhwY2DvkC/ehGIxIGCO1R1CgyO9MQ9wz6/tMjLVktXFmvmhqIEt1f
dn3svUAo7PfwCNK87t/Uelt5CX2AN/MmOj06MLHYL/kLOE57gNspgqplqbH98oyr
H4sx8I9hLA7W2HS7upehyQOTylymPfB9srpI1rgPk5s95/uEqbStW2YLNh0+gOU6
uLOy5frnyVULZ62iQNcYB2g60JQ8iQdBDsfjK2hlJlvyHKJiYM4HsUFOiploDvY/
np70cNC04xEfXlcXP0vV53r9qpkPLbTO5FEnE/EwMEmPXt0pyns7HVXQ72zWqS8N
qZ3WkCmHIMbiQpDWb2W5kd++Gfe88O7wARK3+BLR2ZPtN9K92UbTRZJ1Uuk4rYrQ
hNu1PkkcUmvquhUgBh3VBSxbf7EEHo4dW94u82XDCyHEGsHzrP/ZhoS6JQnWpvW9
ON0JtP24D79+9x7vvKN5MOg/ooAuQfzbZAgm/Bd6aNXtUhHk5YV3bAgAbWvOZCbi
bVjqXhDjTY4LcxyxcIOPEjeN5NznXDT/dXj3LUjrMqevIreXZbJZNq46Ea+3E31A
/GGa2PHwFhFm2fvmf11I4mkCRUw+GNLLkBEJLFECDnnFgGtpT7iQACrhZvL0Qa8j
rc2iVbb1Wgb8mCkLuulCkjBflVSTlr3PEjnKQpsndfSQnjoLfp8TzamKcbBFG13m
yyUrykkhmPKNaS46IwJXjy3hPrRU2c4gaDEObA+jBsJWSdVJ77g37bfQ+NgTTRQR
hMBH41kyE6io51PGOV6pkyOhbtgrEI5Hj43szMdVBhfoDn0Yebpbkvj+dlj6ScZz
w1wPpXaWcxe8jzwv12k5/Z8MmgXxrx7RfcMJ0G8VRnxUfI9wDpBhTXtfOv1icSeL
heoEOOmX4FQqG2qesibc1fRrbBiXOwRVuzsaD2ovM2V3BNkqSkqvtQtBPbYXEn35
oiJBTYxm+L4PdTi4l+w4DxqM1IxXGscP0yFKL/EvMYqI73J1WJpAUoicCwX9dn+1
4MA1WKbUDAg5V6sM18Lfk65Ox+qdwO1aer7711t0twvZS+7QkhzLcSdzL1OJ0Udl
/gGWX+kzr3CxDnWuXGIPm1QqD7zbpzuMn8iu+LCKudYZthUHXkrsaeM7dXupI8kq
B43IB2G894b6oWHx1cgVseuCS2tsEzDjke3b6Sk5hLvbu7LRIRvmsCldrNnNYoXp
/yfhkvEBIBA27sJmuDbH2Ukl/i9IccG0IhuU1WEK4nPb2xRdNsJaR1Vq7bml2nY0
VAyBNv7gJuTDpHrt2rdRiasvOUNaaVGrSNLOWdE1v006O2dz96Cb57KB6I+4Spad
Eo4slzUtevaanrE04b72EJT/M4Hj7mPnnCG8ABoX+4pDpIMl+wlxdrHt/FlQ0uJr
xr9LREyjpcXYddSJlSQY0tkNC5hA9eM3E/krzV9/AmPY+bLJgJLCDq3u55tJjQBG
Pg8kTe9GDvb/KVFR3KAALm7GQuB2m+8yIV3+CpyjE12Cx3OOkv8cc4lYplas1KRo
wIO06YJNvk7ysaEYQh3cLgG6NdpyttEZxL6SO13yuhzS+qJ/Jn74Zmp9NUwq5cSd
dTWUfz6EeXqfJ13JjR7NQ2gWzLokc+C9kPh5DjHCp7cLfdTiz1zPHt1U0BFzVBI9
wElTERDzocn3jYo3F/rOOKzioa3b0+I3iC9bb+j8QaAFd5iTozrkQ+kKhfg7vZeQ
dqaJSdXTD/mA1U1ATQbzuYiXYL6IRH1PLZO/ipo6eaYHyTgRClxQHoQ1dw/87QFB
jcMpdcfTP92ZEa3VWQ52PITle1CfIzACLs+2rvcVyZjmlt9/MvJdYbw7LEYIQfU8
UQDzpcmECgy+J2+2nU/5f/oWyJrNvB4U51BDX86NYdCd8Mid6cw8nLAG7RAJJiPy
vps4sHp0jV7ZSGIheXBBUNG0Mr284b7QN2pguUH1Hr7mBn0lJhrJA9K3WRuBNLw6
4ZBa/OzbeQQ1wg4O4rDXjwScQOQuj5gLJ6oehQm1XNmN82HC0eGOs9ctNalYdMx6
CeNoFiUx6LqV4DLdDbcgcIbh1rmyWWbGDL3rBQofJ8zAD+i+7RMWtY9eJ6EhBKTS
m1ncfxPSDovD4UiSLLbmbagNHVSwN5fllI+425UYWxw3POLslAq0YwxQf+3xLzbo
j8TX9EihFLV0wApGCWke2Xt1qSXwQTszaxpGY8zAzhGrjdENR5y2NeZ/MJKg4sKm
otcj4C2ZshRyzy6eCE+1Y+CyKjowhfs7ukuEyiDFoyrlFTuUgwnevOMUSzOsXUMQ
AAWw9mRzj/uQZuQ4toaGEdpt1QaR3hfxapvix+0L/kTYSoc7vdQY8QrHMXkQNoj3
h5wncS6NKGg41pwgyeukalWQ+vmkgidNUurZbyJCtOO/psmm3VYAijIZ93G/mppn
O+G/q1aDICDhOK18k2phUW5znCZKjbz/3XHnhEvwhwM1yKp6UcANEonEVCKkMQIK
w/vT6LmfziI7xSyDJF7jsSqX19HHXhHcnY+I8ERMp0J6UF23VHWPgOEqdZ68ooK1
uUGWDU0e62esjXFeh8+femQV9/85F+xt84omXoQ9C71Sgk6bGiPVqPqXnFBpBrQL
v8rHAYstwg6WngLe9BkQ0/QaNWYRzRkT+iheqN8S6ox/8OszH8LiFUkMxZo6xjXq
APf0UvmUsBBnxGDSvgSROcYQtQgwzVej4PFv7tjGSVeRlFCFid34+N/ytd+XdX97
z0o3vy//VEpXJ1OGumetC6d7/aeRz6OIiK2Osq5c3AyQ5xM+RDzT2JKuHzlJ/gSk
zIn5owBM3DWzRb+HMWlu2RhzA2Wy7/72X34EoTjhGsTuaaS0y4qXj0/GUlgLCLL8
LXUzdFB0z46Hc1JE2MU0Zlf5m2vO01ur4GP57OU5+KTUe6KvzNsLXOBS+wF/2wFE
ivgCFvPRb1BqEVc215gGIPvEOAKPdF0Q+aHJpJgjpvwagJQUCm7VC/MJgOmimg3q
b4O7pYgPTP3KIIiGq3i346uOVl2Jzu3TCn0NIQdgw8G9nzq1rXRTpTXAX5/SNVNV
a3b10LhNU32MBH1XO0K//H4SXchII/D1dwHqdeby3ekBGzOqKsWoshJUUNOVbwuv
Dym/KP/ODk7cfSPBp2Bi12ZFdv2r5PovAzG/wY7IQth1Pe3coftEQ1QLbVkPheE4
oD/cZLcog1J4FZexrp7rgFjAINlgCcREQsB6fOCfcOw3vyudtY3WafevTqyazAn6
gHK50X52OKfSZlrToUAmUbKeaFneb+Kj5LRtwgQWYrHK0sq5EGUTR3RLOJbyzakx
3hs80Vpoq9O2YWu8o1p6zqyjfcc5Iiv4thmQwE4uzabHBXOwZhwKfZz05HnkJQLs
jCqlxIYXtynWoveW8dTicWXPemw/wNxrvkix4TwXI7hxwfqXssHKNa+XJTaAEUW7
V0iNc43EU3nSOmsxxP480X32YbJawpCEfqVlL0QiyeRPLv4PCMu/fSaNe7HJQfhj
elGPSw1Ls0q/IVZ6VVobWtlg5b2gLYgNikH2A2ppGFm3we06hKg16GbbPBF1vlDS
hD3tA7yIZuvEzoOoMxeMICkw19k4Q0GVusoBoKkSrNO3sLNWmj7ZutD0hZbD2rSM
GQcTohGmeRJO6UrLLRc6FcaNMRr4lWNr+DhmUxqypbWAcZ6h1k3j2rKACdKWdS7j
HKhWhqrgvfT56XJel9rKngJtKLOLxwovCoTzPFmDcPUlVGPr237sSxVQEeyY/AaM
drHFn0ritaFJdjcxKrpgIF2PE143SLC2IgOhD10G8aMqBozZ/uIlKQmzlp3Uhj2o
SLb8EzcyYeK9t+uW+PzsHEYqnC/jQCNRxBwVjUyi6RLVSlGg89vMSkKrr6In3Y9e
knpf2DV+8MpCb6iW/W9TXIkje+A2gi9G3sK5dvNSGVh1RAH8Q2/9gMm6TdCH8isb
FJVaiLuggKDnTXOAosjt/Pfj9r5XwXlKp7wbkjz/r+uSstjEqdevE862NsLNNuTp
JZR+B+apQeSYUlDoIxlgC805mj+h1kfdpHj8VygVcPF+kVErU6iTo9kkmJnUxDru
xNhQ2UNB+ceIO8pje7nQHPrJt32s/N6RSDx/BNUGxfM4UmueUERzq40uo+EkT13z
bEbYb+oe0gv2zDp55FyMEcx/o/4hng12+4MoMisz/b6UFt0ACws0XELIfGil5WOh
o86842Tsptb2CBBwNDX9BiKAIvSUTBxQtV0v1qrqKkV0DeraPhlLui1PB+hizaxV
nVaVVqfr8mumAaPcFdkFWEd7MZtkz8GcZGYuvzRzBBUP01BA2F7jwgUi8lFc+h4R
/PPiQksDo/vQkUaYQWXTFkf1CVEUx5K/i+8DwiVi7OHTiQP+f+WJHmh1qLHXDQ65
KL+Y1eAR09M44yrtsAsO9P5Cqh93N3z5DCGZNKOyDjeO6/NI/8rKNJxxpnhMxorC
OilCYN33xNbZ7ULORbq1URXOat0iztH5TRjdDFzACuq2QM9ne9vPQub5zH3gdYyF
+tZu3Fy3y+5IYVUm+ueOH9TaqdCwJkXEi+YqRZcwqigLfX4GEBz7kNJImyk+7GjQ
t/cb9lW6hLVcy6lFYD87FlesLQgzUfFCMm+RM/JWrQFUilj5fvHINSyvFcmijuRV
YAG+6DNxKq3No6EHZahHQBYh2CAdmZL7PT6zHWIQaOfHx2qS7k00SXyIKeXfM6e5
Vcyj+B5AhFODRXdW4TGfjoIS0M6XxLbWz1eE+wj/ZPqN83XfOYDbZ15v8+crWObE
aMbFFwVCOVzwpVlpVhMm06PLAC0+KY7/TVSRy0IQhy48QdnhUA4JRaOnZmBz5kff
AuqSGkH1cvgHoYKmmAiJCzC7h6BK/kvm6AgOiP+r1+LbGFySzEgKOZ3bVB/rfbU1
uJ8AV6rWUcnKp0f4+PF/d9FYuS6mYLtEDrE0HpCBWKNmijmfNxWNFgmJbaQE8+LA
hSuMEfUaZrX7qgEtWKWspYRvsgdVCYqvFeo5EMRCabun6uc/qyKFcgz+qrm7sb2C
JpWp4DgGy2r0h9L0UZWjmlvW7AhWPmkFF1yprttH3j3xBzmZs2uDCKxw9huGI4QE
05SZmqk+Qx/XqQ9U90jMlxKUaVEPTNemUpItdSdKEwvDsTC7pnMGh1dnln7PEFvP
1/QjXWrKXWQwgRxu02xdPLz5aCu8RH5fgZ+N1+g1oX2zJvc74/nw6HYwDgcmjuZl
QmMBaICbRLEOBRlb3/X3idzjJx7ZwjjqLg0jEA33w9Lw2K53VJaf1BpJs/d8eBwM
D/FhWKNuSFVth2k0QSbQo1KiUfGLXeJzTw6nws1oDcNjIkjpwxOlNBgVB47vC+7d
6ChUeBfJ0tbzXkECbWj0NPk5R7szz/3C256CKQKLoO3Z/jmLhd52dWkcRo3JPneP
9MX6ZwlweYnXRjN48+mIFKa/ljZcAGz74WO0jtKrGSH7Cn9UZZvHY8zpQwJUsnJ6
FYLM/xYlGxMNHdXfQDpYehO045Sr6aBba8mZAvqIrBu61t8Nme6OYrGQBibtACII
HeXhLnrj9hC4uQdGzSrM24t77m/OPJz4C7blpH60/y8/d7KxiFf74yC1buEIOBzf
YPgvwtHLkzdHmNAA1J2AtV9c07SMlgV8eog2TWMNxwtW8zvu8TErLTyuJ0CPb6a8
PGrNvmSQiAl5A4jI55YcLKmu5OQkFFfsgZ1ovwbgMA09ybDcSmFcFVClJ6Oed3u/
DTPeSoeyrhy17hexFSVcgJ4qCXXS0J0ptKGqvGGouX0NQwU/Pv7SaWcO/dqrrSIZ
4frdN0uPQzsxsEuqEWjRjHZAxkpPXbtm+f67C7s8weiyFciUZTuyM7nDpL6+FDQO
oBmTh7QmvqnvYWX0kINibsNK/UVtCTUbz9lsQdaDsuj6itQyLMo18bjZmFmqLMv0
cGUkHYGO+JGlxp/r0tZueaf5eiRTVy0wm/FZ1e41bGIWSYU0YehLsSXZpJA4ft3N
sm0aFY4qRKzU4I7iN0jAyiCEKLdKVUsxwxXlEinTAy0uWryVrt2KlJfMEAWsFQaA
Z8YgOKsjqauzkV+b15qLh7KsFb4FabFBjPNyaIUMWOjqk9UYJwSX1HiA1eY0R2Kz
Fewlju8IK2OqBaKnkXQRQh7CVbPdW2yarBSM/koDcyrItWwgmC1sTud1/daPlVaw
gT1kw0Za1pDEhukd/8EmeD+cJ4peGHp/cURUaKqO/3QYRlGXgQmNoNjPP360pyJn
A4jKZNyVp80iGsxo3zAbbzE+6GA57mpk3Ry1AloIy11mrWHS8JWuOnhP2urclq1Y
z0PS0W6twVxlWPPwZAzGpsQw+oR31MsN1Xo5yt6V/+MFh9iRDWJY5dUXQBRTfhCl
F+GS0GlxIbydy54OCJrFdOex1e3v35G9kP5iMPzukcmyLXH0CPRFRvi0RzLkEfj0
Rnzxq2vgEIcmNikfJH1YHs+d6JnoKmz/TtQhQihfeC7+oIx2BIVu5pIiPdY5XzmV
AzZvFTlBHGRwJN8XeU/2u4K6qsson7rOnb5x9Vx1AJvgnJlYNAhUbxv0W592L4qn
rSuMYznR3QBTsRaym59IoV+9SORIMvwPshQfUvuhEt5Gp1Vvtzy7rRVphZ/twtek
CEL7MNiIQx91w77Bwic8VdfbkNaYiwxhYDG3+hMhlB77QFBlViiFjfFdtDDFTw2t
wPabaNJ6lzuVpWLcmVdve+MdcFuK3VSSOyeJucb/oySUmweJt7MKzbUe2jtPxCxM
vHo0bLmAg+ErJ4ykraaoRaxAJQPhzL8JPYo36klkLoYHk8Rs/cvaWiHtmqJOBCFu
DIprUiJvpyH4KGOk+BVJ+sht6M4xqW1dWJnS8IqVdbfGDlofsP1XjN1coltrWpEp
rfhtZiG9YMJgfa1QhYXQbYNwRgv864RRlzUI8a7LvXXoL7XMoAXUkE+ated+DyG3
mKTAlXpU5lXG4x5DwvE4ajNCI78Q6zZxX1z3uuHf45k8LsnJdRO1srmLRTarou3+
acawI5WW4k+tN48tRPfQg8D84k2L39T6zp06qU7/IDk/loUYMwW/txe88i3LmJSJ
NyLwqhPugiia/rjkKrmFaGVUAChSC1N2LCQB/+oSNXhJA9ANfp3kqSyQ1xRTCyEn
P53hFsMLDlFfx87uREEefgkdAWHqzYun0VRd8CJg4J3EwpKNwbsyxLKYe7lGoz0k
snh/nruiH2wlFMyxA+z+Krl9qNoJsP4Z5K9yYr+2Zwj4YXDlmrXKCwgKvCv99Aqi
SvJJBhCRn9ci9NBo1Fz0bF+uSSni6zI3ubpAmWJUYtYLV+c03F7JxlukYQ2K+AON
OvXPollspDhhdRa8ep0NjARWsUn67vbQKO89dO2OTUcIZseVjAjTuy5fgeI5Z2d0
g+yTbDsrNN8WiprkqwaKD29GJryi43PCMh4PzC4eVCkAkvrUsDc8gUA8bMp+3Aq1
eU1BNNveHlBqB1Up8tNY3UXHGtsFT0i8e7lJ3c849Th/oP2HOXUbK41sQANJO4ZL
T6Gw4k38/kvCsE6XFqSuO304GRVfZpc4t/eyxnGUkkQBTEIZu8K8lMNwA7KFkt7t
USfW1G+thonlJ+2pIiKCHfMDcmHb3jSUeXPAvLtOdp6MSRbZhym46umrJZ7ckfOw
4pSkcRqBBN80oHje7quBuCOSBXWdj565JFn57nFZ94fgk1d5DroflQDZZQAgSYnT
oqU9uPZOUwKoFp12H5gRHIrbRoBZxMunOOamUWInsJ9pKrXdl+AUNtwVBAGKwVSq
xjGE5P/qAG4HA8z7FHsjBWwfSeaQ0oQoKFmyB6DLxnFrMzCIFoLOPmwiSQVuPhkZ
tUyRMnzR4A08aa/6KnrXnPpHky5SlSY8mTz13idasvOMUW+wK2NAkuHIiHAjdj+3
rUfs+xqLlNomqJGgZ+75vwH27YNRMKTi2Enc++CYCTR7bb2Ygb5zr7o98PMYhIGH
u4vNX0QaqZZqgzjm8IL7B29LxzYXwr6KXooFRUuDNHVLctwv9zuxYnA3JHFBIYPE
b9zllmR1Ej7cV1Puohbz6h8AtDd0oNCLWOBzeOCvpPigMXX7466OyLtqxcbfqQYw
zWHeTKyjvw9BPGszB2c5hzklF7g+P00cQZDx+MJFkFqU3iI1DEWNFLbGRC0XojJe
oPnPkZp0C9N2p2+SbyXzq3cG94cQB/ZxxV8g5xYWLNoaHuDLtuHyD0BpPd79xd4w
hn24+MGtCC3K156WY9doAcOy5Dx1nKupKfcO7xuLZTM1q6pbfX6wCz9lH9vIWHue
sL0hc5AhPdPNwTnsjm0tUIGZ+7G95TOirA0jOHEMJCdfLwA/J2UmdQs7P9SO/YnM
2BCAJqtSJTThSXZ0fFORf7/xvnZoBshkJFz8OKwNszMQJUNw1JmIhz4fr13RwPry
C29mBgaAj2HCgANW90ZoGsQPTjY3sYZkIKRy5emMzyrsmy/hl7KekpzaNe5ioCFU
8/qTp7zaPr75MJ69BNHOuDKMpIc0w4fB+wB7PcshzupLeOMlIg/SwKFefWzlR05b
5xhMVgc5IjWkwJnLLDtOCkkRSqwWChnRrwTsg469o3urVMpUsyl0BXsSR2ajNVGQ
QmAh9goqMEUwtpvzAweKMEZnxKwpRp6BJN8QoFO4Pux5LmzznxncUoRW39+inu5d
AL8pUaGEt4sjn3dLH/EASuoW+oizvNRtqug3oXAZa3f+KY4r2hN9joPq5iRUj2Hj
yopGXSfBhHt2M0y79P7nioytu5doXkTEI6x4zOULtElRM3lRDRcpyUloUJDd030T
Zl5cjKmWIx3ZiQDUngRAPAw0FwenNxKsTKqOAdaHPsJKXwv1TWGzWBuP1MrV4d8X
M9qWxvXlLYXLaodRYX0q+Add2z6any643y6BSU7584uAKGr7oukKeeeBAwDK23az
NtmLA0FBtQx5LKTuxixH+SGuC50vk4Xvn2bcCU2kCJCku9xLT/SRrNflLNxP/R1m
7LuzR1VfmddzlqBXz5pwFxBxu4vyPaii/9sIQclaf8F+WVAiWN+vTtrIUGwG2p3W
xzbbomHgZcW4HyRrcvY+5L0QKlUjf0gh9CddcRM75pxMEhN8B7/NSOEK5vgCXh3P
bgY6Qw9qkI4+mJN3i0wOOsIm4bgpi4lZu0Bphp7tk6Qt24ECoV/OrtFTnegY2iCS
wXLuulSvwc5aSs4RzH+1vjvB8cyiBKRBNY2nte0m/mC/ytwOAAwJq0eTrLTcsGxc
9ZSVxqien0x2heWW3qYe3nH+g0aXVSMff3LtYW4Khy1/dqlhgL8SOl0pGAU8HfVt
Mzzta7f6bvPmtlPa6ESqtXXowJEK5oKWQeQX8DLU1p0PM5HwIOjyS1QZebSp6Ob5
43DebtunNCT2wdZW2sOHz+7RvLottd+59ZPxmFGWn/k3O0kcqh9zAou5afrtsIxB
5HqkPU7VQ3dUu1w9Az3M5HG2R33F//poIqJfgkqELfslqdFRFhf8s5Mj7XFBjY2D
cNiJuBtfu53qnFJGDz3keBhF6cqIyKQ8SFEeXz7ca9xZpnh4qgG+TzL58B64mI6H
6/TPIFjdsjXgzfv63PkXdeHsTAEwx7e5VhSE3El8tbqgZ+BPGInwS+/w4OQYY72U
exRLhwEkwQnNuOdXkPOp60Eiwocr4uiSxDeN0LYMhl+O0Kef+CtDNt77i/SPBjz9
TtHPcuSvaoOcukvjD9Vuk2cud/4TN6uqq0nL8JWkwdRsSlj7j/HLa0jon9DVhmNr
0NG0Wa8JmDlWCrizfhVHMY37uY9bMhvWvWXV8CP7s+ezv66veZ6YXuR64ganC/F6
tRzJacvVtJnu8ad6/wGDnEWf5zyjlx67/TJ/hqFH8rcDbdWFLuZA6QRxvGTM78jk
/5gsTPMmiNRwpzkYBkMWvWmQ8uV1+TROCqpJqmjpIhiZ8a79s5TjAfIBp1UANCd4
rwxOI5Jk0IfwNRqcgZ7UxFXV2kyy5HoLM+FwtqwmdmxAgTWp/bfdliFOo5z1PK/F
o9KlCRQ6Bv2o/gO4dEGRkIxarozXUbXVJHcnLVFonpnlP9PCjs2yYk3pGJSgpDPs
uSY50BoXCVk2bgPxCqJwi8ZjfQfeSjTQFBxZOq+EBCPiNlfdSErZhvzsyfbHIg46
/NujDn84z1YxSPfjdqDHVl75ffoXYRmxVByLJqPQ70t1Yncw1sEkfjAndh4wKGja
cYcrhR2Gtj8Pmz27J6zv/O/v4fMjIsgDHZrDs8Y/B686KOPlp+XNg8szqlKEdLNr
IhBREWR/BD46MJgpZyp+oHmrRBgC9rP7YocOmx7Nj+i5SIh+NYboD9Yl2ThONc3R
60AhGdA4/d+5YFZAYpGwuClewhNF0pAhKXuL+UNaDlq4ZTYYLtwocwiX2hDB2suL
nNGnk0a7K8QFguAH0yVg17jgxb+PvI3/hhbIaoCU6XGWmaxPr1LXFPOra0aKUMJk
k0LZEhvPkDNHApGCFjXHJPTiDqelVnZ0IX1uURiInCBZw8ZQvxCRlei57cG05vcX
u0JHwZcreaXC00hSuWUZ8A==
`pragma protect end_protected
