// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
i8U39rPySjPCbEoteArKGzKRz5VmkYW+v0n+Dwyz/GQ/gsA08HKvoayw05LT93x5JP1GtDKlJ2Jj
4V/VZO/hynqmPJrmzO5BKIlnmuKu6Sxk4xm87Zo+TxuIFDHmu7xO7iPGCJwfKJ6ZvA0FdDAtKlLq
BqjlIOH4v0mLhzoVL7xGb+7UOa0c+Ei0qCiBuFF2xHsDNWdQdfg8/FMxlcz87o/Hi1LmJQ52WUoI
SLVm4ZOcz10EWusInRcYIiP2vDN8Tk53odarq1t7MQlpraATfruYux/QizsekRbh6QY4UJ9qkRuL
2AN6330FcLPOkomy+ul/uAs7wOSr/GszSIEW/g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Yxp/DI4BOY831aAiQ8QVqwxad22QXb9vhL9291uctyjvI++HVf8ErxV3FCCOkCD6vpwTIBZ25fYY
b3mC6hB45lzzgdXwftPYMZIoqUqbri2/1WzOhaAormLagNogzotjSqQUF22wYVEPu5D0u3vK2rAh
dmR8D1e7i61ksjMFZczlOqHiMik+zRmgxYfoRBUe87nAEfGB6BzBSgWOvpw3ymqYMjyXbA+CUxDu
8cmzhSP+uJG9MfIBgqnRSWM0OLFB8EM6H1W+7HfFOfjpigne1YKS+hKFY8DBj2K7JPb5+26qtgeQ
TLOsGHyo0JvFXNRb8lMORqrIB5sj/vqawceftfmRw+5fTWQtyMQY0RDkz9Y710evV626PuE4fQqD
AP+LBGq7nECrbrtW14nd5ivjo3Fy032FFbD2f+rFamNd3RAHmeaaE2+htpqC8AVyAaXs/gTLDgDv
5L1jUcA8y27nllWssVmP5YtXKhUq1hsyIWXdIwS51Zvtt247EiMPZfI9+XO16QvpH135H4U+6dar
Eobl2lrkPui9zV9xqC6HEOk1o+C/03LTX05B/j29HCjALQVHka2mSuAAtwGGj0pp001vagkmWAKx
qJmGSaOIucAXjkyDINdMljMNFtG74nQZewKISDs/lAGAzqVzUYd/t7N1qyE/lL6a7+dnmrCVwcBx
nwqr4bLjwgIP6n6iZFFHOSSHYpq7ffWk3erStztHd+owE/N7HC0fx25XUEXA5oeO2QWZg/+SfUab
IIaEjTv5Pd6+a4TRoRC7tgl1/LrJdisK17cl1+4yYbGo+rAzOQUpaNlzQ1QZd0stEqHPlEBiT7pI
9sVWd+IPih8HVYC3CGzmn4Hf+2dQ/sy9zIAJLIlBD+l7blDnRfa5Z93nv6XqQqvuXxMN/t4xDnAi
0Wf5aiEFz15N51conNJkvsBBmWGHkljdsXsQXXpf91fbGaP0feY381bxzT1dUw28mRi5MU1snmPW
TK65O5VWd1MgJ6Ks1MV0EQuTsbnoHg8miWcQSvqBP9NUVI6GzX+Kc9e5JM7fNe6Y+zuD4x2iOhal
2XOTXT37DOBTyxBd4zdFsZ7VEaQ21Qyj5voGRjRZrC9bcYwH1gU5oRH6x4Z1fAicThPeUPhI7v/M
rRPmEi9s4vQ0vdIyYej+PODAEMRUknWCpRGW0uKvdEQB2sStTqr0aJKC8MhsBrAa2Lgvx5x1yEPj
/zfwEROmPyXPdy74NrA3xRfKanb0cA/nKJ2KjCast6qJ15KPf/+XqfwZ/hmH+l5Tz+q+23mx3T6N
TwpmhZwBrq3YaDJ0KlJnbuaLnAfMI+CLO38/ktG8v8nYBR0/IJnnSCD1vZ1B/yz6QxxZKRsMc7bx
HS6CKyQVuNeZw6hb7HsXzQogp+3Wo6JoCM1aDcfOG0GmFSl9zghXKtJtV/Oi7UwcnihGGq4iE4a3
IewdfqOgESsKZKhuTM1Z1hHqbJm4OAzy82qLp39x97leu7fWkHuwiWmfsCPcFNq7ofDrz5LzWKsl
594KvosG+41OzmTOaWMCD+xPy/Qz7LpdikOwnb0q1Pt443hiqdqjs1jcL7RgmdYB/cDhx6+3VRrb
DdgwIkMWKjSfmJQwHkYhkYhl3xXMkbQLiCQ3GAVKd4UneB165oFtlJdq1NcFciooIjQ/fSQE1cNS
SPn4eEKFk0xugQjQatkEI1Ix4uVDKc9DE9fb91gLsVmLTebKyURTclpYLeq3wu1FkMtEjjJ+ACuk
0QskZN57/ZSFT9lJJc7sxbRJhIR8IL3pAjIo1xvMKVnLN5PAMeXVtDTtWFaKlcKPeG8ueOS7vkDO
qTeNfsMtIr0XN5opEY8+KlIEuJs3kgvVs8F3828Sr6qto5+IylMd2hiz/pr0b/EkilPSE5qTXg+9
UhTnbfMr9eb4IOnjLdmJRtxRt1Bv7KZVXFVu8AvCUn5n7Os6678YWlxd2YjPfFY3Thfq16p82egd
hrbMEI3pQbkj/uw4Ou/TPi38A2VcN69M1AH3FGLWkPyZPXZq6xuJvNtlKbuINjouBQkqI2BH+SP1
vky2r0apPOTbXDlJco1C/qvNkRHGlT/Wn3R6eoW1a/3UcN6mh9HhXPXe1grdtqQjZulmOBH5JewO
yBtaJz64ZYCffpsrKbqaHn7qTtVlQp5JZ/1GrIXF54SZJPeiXYDjk4bxfKsqVE0JXqtKvkfL8k1r
qoLdK65cni0OA906kpG3jT9i8h3YYn+2kH98hjznZRDVv/Zsvwqv8jiatH5aQFgSNS50PlH4jxYH
MQ9sd50sBtaPnNA8C8m6SsWj4E8qRSvSmd5HgddqiydqK7uGHlmVuyJdmsikBdyTAWJ3K9wkiQ1l
7HSUrU6UdIxl8Vtid1JYXewUe5R90CjTRfEXmE0kY+rspO0nOptBNIi1YP3tBTkR1gCJ2bdQZNDU
nPkAmPJwAlLcTBgl2ezDIc7sEq39Py2iZG1/G54U2m00Eg2Q/ZsJ+OzhNS83EK7FHE1NGK0E28/2
rhFCnzgO89etlLCDY66G26guBvnOKrjiQyK2fKfc1ZT1Azv4hHSW40BEG2aty7WA+v7E/QLdnlLZ
Q2xoQOu1AshQrY8dLVhR6TSEST0d1W65Dp2tLxGR2pVJJvq9Ct0zrgBdn+0Xa8mST3XiNP6IHv0A
d7A6GFkHEAideYpz/uj3D/AIf3U1j40PNAjOr5euO+8ONQJeGRtpxpSVkhdxaN9yL25RdVVYS6oe
9NFaVexo/kM9y3oQN0XxM5xQuD9jq1NxHm488EAU97atDz9Td/A7bAQG+3Ig5N8BqBJh4OrHYA80
YHnSThcl2yBq+JzB4QotA28SYvByVlxYiE3ggjMS0DOBJ/mAydmIfQtYcg1GtGOab3b4a0g8woxW
WTH84nEUXL4+eQZ11bR/jL1jKQww3p7BTYoVoHtLbvyvsAC/CUtyvf0/KG194g4YsycyUb+7jmwC
kZLkQW4jTVmvge6N3td0fmOECJLpf5+Lyo7tOQW/epOiNU52cb3S029SN+3orgsyUFxy/MUu7uS4
F7lTQ5BEedHRD8AoDzrNumcS2bWDM7kPvwhWElGuGASA5Jj8kkoO0kdounCG79+9vSDGNIlhieO1
CqokaSmSG8CIqdQRu7MrQ/raje+wSvVaR4KE1NXdVaSh/F+ZaMYy2VpKgolq8zAdmRg8TMYtmC+W
2EQmrueUordJFSB7zuWs+s3y5Ezbn+IuhiRLu/K4+0m0lW8ycf9G8zkWufCD/zF4tWDg4uBk05Pp
Pl3fScQ9OrZhzFvsVO1Ajlko9L0aH0PvcCcQ6NrJXPFW/Jjjtq5zcMDY+Vgn9SfpdwOcOnrXPika
TFXYCnslViu4VVHBjKZXgsAg/EYi/KEAgHIfTx9z1CHvohAsNfPgFvxCVP6jM0qLSDEOCt1lx1iZ
abemHMEcjcT7lky92W/ZQ/GtxgUUomZVWnHPFMqRw3j+GxpLVtNNA0UtYIBcBsxPpnh/xTX9OfbN
aFk8ZOn1zGdnYjDA75B+sVd3OCvrjCwoVjaG3nf4eI/MPywU4Ek+dUTDYpAN6SHRksCp11StHFGu
+I+MO/d3h+QzKXnKMyfKjDN35bTudIpoCiuCyZTK+t/Gdq7GRys8n5NZWwxfAuA4KAbdSj8zclTL
ElSclLx38zeMxSEgiEawZEzH20CpwzYn71Wz5uoOePbLtUQOa4/rCa566OyYD2ug1sMJYrxHE0kn
rsmPRh9nZiurHJnAF7cGSUWpZW+DRynRCwvbqIMeOwNNHxpPwL9GdzGRYPb/QevrlA/oyeMdIlJs
ABXy9klcS8CXQhh9rvI0YPklmE+gDSU+Zs3gEYaUiA1y7Tp/vWKN+dsV8RPOOLdbwyyxovlOzcsx
ARfDpy09E1eY7bpLBgy6Hjh1OCkTCHM9IVUvDwfeIoEw5jsNFAq7XFZsZzr/g80hksKw5ZVdMlWk
BlUi+JxNJb+FCqHireZAoKtGob4JGe5QHruvwYiza7PTq6BYFGKTmRIfpxhJQcCp5GfYEdW9evCn
vA4oEWcqLLMPXZ7qYfWXt3FzydZKYGYSSX6emki516esTrbvDkIN6VoPrVVVEhoyIu45eUNl7UJk
whW2EpH4fN08ntoJvFy+0BJn3HEjjaHLWt1Z3FkEieUnDnHjT4N+cRuSwqMYh0b0Ref1V6iU4xuu
dnPWv6x5/3apPG4ipoxVxgeXwnF6KnS0tIfgXgrZXSL1qrjdBxjadYV9A0vDOC6mGQSKY+e4/OCn
/xcrj7WVbLwdgPj2RvEPf9Pe6d5CT2LfFwn4Df3quQGr8R5tA9LyOcSpSUBfBvA54da5Eo42iuA9
3NRTLHU1JAL3k2nK2oODxRwBVhomocS0ALwn7gyKAHylM+Hk0RGyK7kNi7TgrNprJomYAejOz42o
ZaXx2o7X6YUBG7uxXZf9M2Jfnhj8WpJYh4xRfdyMrpRJjSBEWojBLiqsl6l5LrykQzX/4lTY3ypf
2V9bfQXWJhfDPYM3EQXyS6kQ+jKf4kwraC3GTr5kHRAjSkzjK7sXFQ2hsc+HdTMHlCUFPCLJ97cK
uxlhtCdnQkKJhmaj4V6zT6tANCPJ8ew0WPGnQtOVTjS9GdgGr83aLjY2DkATImDTWcGy91i0li7j
rc/Hs7JeH56PuTvMtMEu/lgU31AxRljGIIWFzxLcbar0+ZH1m6ydW5ZLi90kScqf2u5JF1spdKrS
kjGUHzQVq1/np6u+05j0fV+O7XHOQvv6dZ1qkZmk7hyMg9qcyI7EPcVk3Hp9hsHM/pdFwdskvh6p
wW4GNa0UL5/o5B1Q0nuKLcIiKkD9+4AoKnGHixSQ1x8JB61At0tKL7S+KH0twfiKjs/6GXaJcZcX
MxYLkABAAvmDyU3fRKy/VLR7YfhFWheP/jp1RUSagYOcaSGR9vvewACTuhEzI9u1AkaOS6cM4fXQ
qMaVEAEgrgwcQ6BTZTuHERU4OacjbCNeZNqzyn8NUvLELZPAg94g3iFqNEzj9ccLFauH+sFY2ZYV
4j2I5hjUvTLzvBmhptC7Z5k9dn2GMCLDDGaeiQZCtOPYynR9iYcKoh70DcyVssMmLpmMdG4lWHHM
bk+MG0t9+bSACM2MN5fUrfgjt1Ft7kz9FM5Xb1OYQmQIm43bxQduENDg4mV3dk5FsBk5fpaGXrZE
nw5357zARyDZVbqNcQCu+/C16j5Sz2Lctojo6phdrL1lt7VJhFmvyRD8u2UTpqTxz2v+zQRnh7ai
Q506E6IvxdVttlR1hzNIbsaQ6ZeAwmbeeTvN7a5qB/cqn6Rk3OXFr4XWcuV/FCc/fz8xjIsXbJj4
G6gxLcnNWtQUBBJoUlO5lFGOPCMXSG7BDORfhWATH9/wGxBV4zdhI+P8lCpe5LA6frWsNG9eOwyF
j0/GVl/e77GBWe0gPxEwMGSgVdxobRauxt0BWEirDSafnQzw0DGT1kQ8Sjk3kmGTBoRuNTd5HGSt
yeEKUoImAww3KEiuNnxJL5MNWpU0yMu+tDFLx2JHxvAKRT/HTm1T/EETi2emMgAzI0vgDWYSatcE
a3Xlfp4Y3bZ+lvBZYoZRY4P7MJI4xLaQxfN0WQ5oAdJvCxncEYA3s5Zp0Ik0jTcK0/Q/i+V4UX1/
cKu1VY+9lPRivD6i3dfhqckhUCK3mneiH+2M+8YLLZIPpjoOcKei6hs04yR4xEfCNL5N9+fhALXm
QG38fIbsxg66RgmKr4cMi/Z4MeSb8DY9AD85D2c+S7QMd6ZYMndpcjdVypbF/uEGPd4ooGiUIEYB
sRd23U5KzL7idYMaFUO5t/0Cclfv0JjR6I75LfBLVQdiw7FLFRoiL6dz2X/BXtd/UOVM5MZdT3P4
qrkDnJgKHfojvY4PDtjyDSvIcyegxOHzVh2Vi/1VgJWm5BkiJlykiPpW5yY8i2NvDDPduBKoJaQk
vpWkyINoU08+WFWAdjMKq/FHKhM1jR14izz4ojG8TcdKNsrStVuAa+qRWYtpkjSv2//+m9x8sZsO
VsM3NNaAA+bGmd34XEL6jiOKd659WL0YHFFEZUxl39ujTX3Amj9XZIxJACXsa1LTqe6Z0SaqpNmy
5ptnErBFwvXvb4gfXKjY7YM0upawWJsJCZqYYC1CT99Dtt+CbnhSLrox/0TM3UkmHtlu8x4Uexx1
yvapYxLylJJOj0YaTNFUWUCpeFGhx/A2xArjrur4hev0uBUspqDovVfopGCqr+UqZMmeseBDIPWj
NsSCay1v4KabhN7E1KtmU7tBGXsv8/x3720geRXx3Ra2XhiDtv/D2kE8BjAcAR5syvRqypsN4hZc
gwMhmA9Kk1xjNbumOi/0spPjQCZnSSDCOkKSMd0DMKVPhICJ28geACohyS8+/rfC4tJnXZgcrazC
tplXwCT523aYmGaG6/S3lSxmGD7x49etKOqCvQT9EXpalBYjZnlh/+WmCb084w9uj4KD4xqMHWc4
NraNaYbl7EGxJVFJZBUizkUfLgHRpxs1acCrWpzzFpwVj4NfN+op1vI92R55OaZrVli1Vp/I4Wnp
HjA5t5wMLG4qHu8XMW3JYXcbIdz1Y1Ez0z60zWhkderNSPfdpcaBOyzSoJRnbXt7xxTh4VMaosch
t8uvG0DebJ+VYaQ0MdxpepHzoDc0xnzW0M71IpY++meiZjviyP2+cVul9vOnFXmPNta0td3BVo5y
iC6s8bf44gqHBao+H8sXvLBv3yxgQRdF+SrYRDH9k90tVVyfgO5BQ7MiiKUEutlu6gW7vJkKw5RW
FbJ6ql1QDdThGLsdopOaFpcAjfYG4zRFsNrQgpGHxr4YyF2HnjFfkVd0fIRKtq9EU3hznFgZ2j7e
ejJeNioxhP4p9O+2JUusFTQZ5ZXK1cHD8jdvrUsZvBFQkdi01qbGbp6n4Cu/0AFAtgBdWqagb1fm
BKGTZtxwXeX2Swtoe/SkuktxEtXrDp6pwn2iLr7UBnQ0FFvHQ2PHayWaJyg3dUTp2QM6sryBifvu
qTaUclW9PvEB1Hx0F+uO8jdRRmW9NyAeTDc8idU7ylu+fTep1nsbLsE2D9RoxW3n76l07VhMfCZU
UhJqCHOviJPzjl+kT7I3qHoyMmz2fUj2AKxznucD58xiPN+g3RIDwmp4pAdw2UWjVMnh3koKpUmM
eNJJjaR88KUSwmfhdO9Vee0JeiF01USj1plVVlQLctAGvSiU7RUeEjrOkVqLakxZSXsqVtibk2cE
CpFuUGRoEQf9t1QGQh+LC72H+yuQikdLI/v3FJbeG77jw6rMV6O0iIuj1eqhEZe+25DujF2WX1Ar
faEnMZNnGSnf9O1HWiZYpmendgoKsGXCCJbY/YeKEUNbFXzUHDSn06zo219bprsu43RZuaZMwqvc
Nk4dxWatiZgVwgvlZMJaMLKXpxYYp3RhZkh/NNcGJHnQDVLv52NJ+mMJWGtNZMJijGyzqevtp9UP
m9pGbzbTZSiX2Vqwam9ARHCJUN0kMh2rmHIpZe10DWhck0MoM/fX+LKqkRva4NpVrw+0UCVJYO75
LZJRdtfaVtqcQC5IsKQJTt56pY2McK/kkFXtSUh50/NlBYnqgBUAqYhUQwDwpgGsyjmnCtF89BuG
fHNAuxhwAcSGSVNcyghof/vj5HD0h1oiSwkYG6k2pQUL3rUFH13LlutsIDLsJ2XPoO8EFgFVYkNW
sbUq/uZmo+bfZB9BKr4NJyqt9OapkA4wuSUVd+mgqiDas5rFGWBt9VVX4cCi4SPcK/ILAUA6/CuU
UzzWT9YnvRordw0ZBsKZ2FnC4ZLju6M7lfpaihrjs1u4rs+uOvGheig5CHGB+y+H4uTyiRCetBn1
feRAdZHKQ+1SrP7dmZ6z5sJGTbDmFa0jWMWqJ3W/Mdf4xnjoHTcJepL2ZMw1xQq6i9R8FA/JvMvZ
B2bFhG8nBkXjHmig1bMe+BSlvx3dpCcbOTtVYM6EpB322P85dhRFh87B3piXVdhiQ643gNExyF2X
z7fi1p30b9mLGfp5ws+OZfjjwI7XF5jsonwVctszJQzMDnY91euKTlir+rOfTltuxFmIWG2s237b
mY/OvvCHY3PqWlWGIhZun3E7qNnkfdWV3vx6QPdRbug6/iYnZcSSqFQzvNwfjobpW656+fbwtn/n
eYekoQAt8pfisJ24LoxkcVYx63yE2D4OtwoFYLTXOd9hYLL64jsjn+PQ8JZViSSoBrb51z3/U8/+
UzxWX73pMczWPHzexb6x+AiZLbHxWMOcVdQ8Yi0N8YtpBufuhWRU/xqGS5A5XESHjksyLcFZyC+P
RJIThACAa2yJ4TBXmXUElykGWSb3UqaLML+50bzNvfrxNvkZoTAeRY5fbr5O/VzOmTnlbh6SAbdn
42B1avwhBvoJZXpww30juu7CX9vLritADjATgiTET4J1CsaKZAtr9HgUvusdoDHPmRLDS2blZq33
XB9TkLfGloVQKmutOPsucveJrKt8xpMhplv58bk47uWMemZOX5RbxWOECy6GedMeQv85TyjBlq0J
9KkC6eb3zxGvPM4ONSWoFsZdXvwS9oRkY0kiLrgFJSbixFocCEg6f8/sdEdwd2IaUfCifHEXkUtF
C+vksb3pr2WEclyvGRUlksc9fX4HxYRD2jAvIEk4RqsPIAWJYfP6f7ufIkvZGbpXKjDSyfx5XMt0
SvtmK80TbLdxMkrsoTkuDIX2DDn0a7Jp02p5Csca6pj1toohSpPgQfeyM3lKXGCKwfFe7BJhyCvI
zUsOeWjSTys36W8CYjBpvRAevT57/QjQjnY6wxM9vVGkWUmIFo84oEdcMNBkowUnVwQFDYFopi6X
wSXKyiy6uGZ9Pqrq6Ng3NE4Aa8a/m1FG253VfU3UysbmkJm0vzatC4lGz0Nr4xaRgmGEqB6FLuLx
vn6simb+RGL3eW0Yw/xdTvbHEHTaybgXpB2xM3xrDF/+A2HURzJ8FWj/9Gkz0OdPpHyPAYYciUR0
YyHewD8VnIvPjM/FcWtqiqwxe2ruW7v1WeDtvcxyDjLLotUjPlFn/Sqeg/KXYsoHwAWOxhTttMEh
LcLtZm+OTSh4y+MzUR33dpuxlIeR5XUVBtF/Ez3AhoyvDRXc4BLNDPo4mc4sWkEXl7ji1UQl0yOZ
D1M2QxV1EJ9jsnyBTDIZeahxHd8YrTyLxag5ghDf51ruUdI5m93JoN8aWH7ZNC16dQ2TGiG6VbmQ
4Cvh1zJLnOxiL7Nyb/6whquRKxUcOSn05ggaibvsqY0IVeuFhK9PG9fo66ZbdkXo+zRVFYtl4m1p
KK27EjCFxOrgUdGsKncDJqexfMjIka6eVgG6Pvv2N2qnSAmhW86ASgxvvnC4oNZ+JiRfMK0gam+H
B7H2KJRKCk6044/FDmas8WScarI0TfmVrpYlenWL3sL1Lr1My3rBHpx6CZkUfGTNwfux4pDgVuyP
2HrK8IxnWzPQPPxGFgYjY4YGwhle+SeE9HOWw4i/gmJQhxYml/FfbQ5y1LZjaxVIOtWW+H4q7iuQ
DCIqD4mxA43tvH7hZk1gALDYkSL3q8QVSlWrewaQ4lKygIzX8rw//4wDwZNLjbHk+bTN1VTNkqjy
bUnDO504TP2zufP5kYSGHjDhflzF6Lt0SwnjNz4KRKum10JyHSBsL136sWTlwyHicavPoWesu3mf
HKWbRMX3M/WQtFTcb3bOCetCCCTwXK0eSztfsgr3vIh5eTdMhpCkc+QfCWdb5I2AsZwSzOdS9MC9
xDoe0K7ar36wwo0wAjpz1awD8RPghh5kXLg+NwLioovOSZNwsJXXDzhrE1x0hORFBCOnBa5e5T9I
gXHhbovOClW9YW1jIHXjfxmXhNAj95YKCJcDXmKRnrR1gVNbdOPX2Y1E7kg6MuAgF9mLlaGbZ0/R
bemx5i1WTPD1DO5mHiV7fQy0A5p9iPjSa8v4zR16M5XhasuINBDwo8q2VUJHdMCe9dUxlfH8JDOc
f2o7PzIMPibyiZnzfNvltKuCO0qTal/Faub7uiJu1JHZ79WdpEVzWiBfmpsLZSxcszmPram9UbAg
A/DOuamp+tTy8DgJmHjy7c+CZTxiwt6qvVNmQoksTlRxhvVyP/0U4nO26fPqcrkaVNVMj/7DV69f
kZdbjGhnsiP+zE5ODa1xchsT+BMxBUON79BilHlZCJp1qTgs9gABDjr7wXMKy9cokQRw1jnv6AKf
Y+5iP7TZGIvz7aPrx8sChsUaGoVxFoegQN0VGyukIGE9XQUmZetVfu9o0gndanDwq1nIalEF/HVc
bSdiaOoqrE9nOsPDa0T9d6aBmuGetrwAT5JMsyaH78HK7s5mweO/u0LdgWXx86+R66sorzJsABy6
LOQ9HfkzZ4Wgxt3bu21KrDmbn/9p9ugXpjiCFHwndS9JCAtbldqe1R4rLlxV84iyBf7HFqiPYR6r
XS2qzgjGc6uInNmirZQM2/vfHPyBe0cJlobeOyJ3AwYaITwVQ1Gipvu63xnO1AVcOuctX2Uax/gB
fSdxpcOVbe9dloluAot7oVzwcxjDI8K0f5K1d84Q/LTjBn2TbT1274aR+kOGEKGuPBCb/FUbJJIK
2ell2bKN6E6+T9AEV43KlNQb/80aPrL4nw1oqiW55DD1/rmF3Ks/6IGjB54ZCOyrVvMd92+5iIP4
JoOCSkq0e2ESS8O7NDADxM1ilqlFZtrHWAEowxbJJNAQJviehQe/sujRaPRGWw9dyXBbM2dvWA6H
DB7T01DIsCgYIVyD/lonWuI//X7N2XugcH4NPR7TFQugjzQMtVrE7gXUuMICnlR9bnZY9p2l5+HF
FwmcHtBCjjwgKzqTnEB5h+zQU3Non7lnMfQsi++On1APCGnUBqkrXjikpYfqwVUFX6l77+MA3wbE
nNaDmMuoWp7YMkcIw7jMoSNVjp2mOOrTt2Pead+NrdT0freN1ZkLLTDn7r+6n1pJOOn9tnTBXrWJ
xrdNSLDGLSKJu/O44o7Z3GhPOMjubotjPszHQnfeAXk/okADZZ1Wulv9/F49sl0vybQ+REsAczUq
+cGTj3Ot2xKuGyiAeNS+3Fl7OMF5S6zpplChuD8IrI0la6u2ZWKr9Amh7Hgda+MwyM673LCluIId
jsBKLq0EgbHs05BvEX3Ck774E6AZxMlwekSbEcHfgtCTgI41QjdVsbIxPVZYv0edZFXyk5ChKfHn
Q0BI8RbIAVU90F6dc7KWTvDIDQSad3/R3koFTw6LzprTAax2hmcOjx9WppTgfyWTDG+uxA107au4
D1xZiq2l/abI1v8UF7AZiEwaGlWFdgpdAjwUWgoqPEMLL6GDejY2YnGYh8wwEhvGzUTEysy3qonw
pmhQfc6VQ2m3t2BIej/nJQxSa7bePTBHfFQIlZg0JDx8lOfq+wUtO7Fo+JZIG5R3Dbq9E0dq7xCX
hcM5/S0xgc2/xghEnxCISDzJmW8XWoAv4ZVctY7LaUrd7PuZfRYU+NwVxmJUqZNwYMuxa9wm62x7
LshqYEUfUGG7rEm1tX6y8Mipxtowur/MmjGhBhGid0/uk0oDqEbDbDDYo0tlv1grqS5+b3hlX0De
CGTPJGuwAXVKuo9E/WQnKpfilFDs2pvm5TX3xo1YS+PZHu6SOtGfJK5lOu6VdaxY2Oj2GHFU/9El
j7OcDoqFYV2yiqXU02+VLkgNBJOwfZBEjg53XjmliSWYMDUIhBAFj0f3asRzBee650fdPc1TSsEE
ghg7nTb8I1IM2hRN+YEPC07fOVzy79ROaWD9k0DK/PVsgFsjkM1xDiSeft+o/kTgIx3FcD8lDT+E
4IqOF9asaLv4+tQZJJngX3cuRvHiD+JHWxlKiR6T6eEQxYKkZus0bXFPBgsM054JHN0Ssi57D0fA
yEXhoOpCW+Q3KPIeqErdqym6giHxozAhFr0tvJXWqaEWrmvh+hBJcKA/cAb+wBj29mkXcN+sWeMc
g0+QrPnwopLpNKhiDDZVFpbdyZ9gNMrmdRGyczm4csnyvoFFkn1/zNFgpzocfZ6/YaAfiE1yG5iC
CIC5DkEGbhk+6Xe5GAjPbnDsSQrehRkxjDsnBqeRH0z+b0x8fX6PfXZnqhl8xNnPQj1I64npOETc
GVWEQlVgySP1rfy/gq/DYSQ0hBvzUgYmMAN6h/Fj2qoVCpnX7GMA+O7d++eTIsZFyZL+PeeTjbX0
4QxZt7zrbnmS1ofuth54H9xn0BEJ3jwnzGgvxqoXTqUvO6clfQLojQdHDJmzjxNDBELMR9GUA2sQ
pZpJ3yj8dDajrI1ZlpX4FJQynJCDCIFvgg5alJJGC/bzerqjnIz10bnP0aCXLoSigM/IGgtT+um+
in3OTBcYjqwM2WJa7f0XAa/swTrPmcj/LKP2f4G8Pw5rSkgeK6sLgEXLufh4v3tOFSgMRaugXNYJ
c9YqA60eE7hg7l5Pdlf4dy2vXl00Lcxf1e7ov0qtgevYdivbvjXyUAfRAS4FVzpe/6CsN3rqhpqQ
ISS8/i2jEAUVaR8+o1qCskIOcX86qHdIlj4MIONxUjVE9ktfLo7r9Q0uHAhZVDu+lqxEAJdYYf7M
PKLyzu2O4L/KGElZbG4lVPnMS0dY1pHZzh5h9346MbuWPANxXKNBZytwLzAqUZOYEY7K5EAY/MBH
J3BaHZQmDOrnRXKh62OA4oqnXMZQTqjCQ2R2urzn7dZ59wiAMNY5bQsUuAxZLnybOtJImUDoD2Pu
+x5fQJLnPjYcTgjx2DpVTRCjVcSrFKXcjA83fmqlKoBrZAELbMHoUaEncw5p0kCpMTYM0miyiMuX
7xWfH7LdClL7vdHgXHl/YM52K0BfyjUNsc26AiyjwDMay8OpgFQuv9keKoEMc26Y9lLxisrYgi9O
9GiXHjGv2tRoyFV4gANJ8RTXa2ABaumzh1X6QwNkhflc+4yrOwFmWbQY8jTzmGQPZQYMbRh388a5
qwqseVBCiGHrhLcSa/wXGcrbDhs39IkbNIVTopDcpJeFC6Z+vYChzHIEbF/SiOV/+J3epzss1l/k
wodeePxK0o5IiJM/SKvnGing3XzGzxmrJxjRBcifO4YxcE+uJzSuOaldN7M3X/SzRUuEO/4v7Uym
CvXTE01YMU7/issqHVPQ97V7/UQATfWyYS4yA5PqrKLNnTCf6a7SMDkrt8O1PQy4jPeaDMVUXlp9
Ry8HSsjMnX8UNIxBW9aoQsECAQGLdoNAaL+zQl/PBAWwuxF1460RfH/QTscbg4Imahy+b7YR+wcb
TOq6n01rzHF6TtCAcLGbfNChUXI8vB2jRTXstLxxEEWYIiZB21wUTATPmsks74vF+9S8iktWYIBl
5wCWJQoZ5Pmk8ULZLextqDCb4YMlvuPJiYIIHYCQ5HSW8/kmNT9dG+g7U5hvEto8sW2Sn9FmRPvt
aKgpwCXifTgdJKwIDvKwNZuEp2WGXOw0ZPhc710Zles4rh27ZuKp1yewHVET/eYidZqauNx/U6EW
uo0EpOQcTed1UreJHrtushCnJJ4F9HBDhg8UKy4zY6CLpVBDil01T23xAobpXP5hfozb7ux9OnnT
Eubd1JI6EquyRCojQCP9kjALo1tNNqhGLGI7qM5NO/VP1VpTt1iSthzbL2179eQVKIM4XQepDtMY
5vJIWIS9v0OcVbVl+J8qJwiHgyzN3v4ibpSlwke+USD8LHZe6OeuYm1x5NuN1i3xHk6AZfpqV0Qf
oypqpsmbYsd27Rly9cHMuSX1KUVpeLP2+HBCOVpTuenRi8SsDniS0Y9YPz6zjp6J9gtrHrnVNqYY
RE9hP0ltKTtNLCbF3+F90yYK784r0jvRKMHfOfTsCnZeBd6GWqJ6OilzPTQyhfzjPEvGP14GI8Fp
VcwtS+HOATwtcg88cx4/tFQDkZGJFa6R6SJbn+2LzNwVoFGjRL78nJ2BmNFnuS/bckLKmEBUD8EY
yZEHoCujRPUQZTb9AgTTKo/HL8ARueXFcrkEJOGIPW6LITIrEBdwGgI2WguzzFYDFkiJs08LR23+
eiLNj99hLsPXsN/YBkkulqnSR+dvn5yH2N/GgO9vbEyHUhy6dfVe8o4b1JFlpft2fM/6HbrXWGz5
hW4jeDGSXtgj3msnvStdBOxvnY+xZ3ojMy/vkwjrhoEOccUGYsyzEpQm6RtBznuJMBhHyOEl6Azm
rUw4OM9dWY4Ysn2RLCg65Xtd45SV7xeFFp05byyyPPDlfj9s8zN45TAlEKgYvz0TnPcs/RaUYhBC
SBv9JgDmAjU++UqhZlZd8BZTdexrgmdscz3oZXnbWj2YyNNhlR3RaIChfhHnfN7EfNsHtrQ1j2Yh
+tdzdyYFjFbwA0Ax2uaCbCkB3r8rPwDncQ8KXcnSXE2jzVIOl2aMSmeLp5ZbjWaAx8XVZUT9x7rR
rb9LGls+KNmsJtACqfpxQMqQ8uRl/jX0VTwW2ceeDVhVpJhgI9Ty8FcF3ehVG68lKstjejG71VNb
8+b6lq+GziBCLVGXY0oRcucxvYjv2/RxuBuEPWw4hkIVh+IGaFiyCezZFYIukDJALf6J41YAAnTn
P2CLL8MZP2kfV7HwWFGm7UrAlICQnxJwCxu+rwV2ZzWUKbmVRTUv3rMenPZFw9sBs4KU48AxTj5G
BS0l7sxJBj2JeZsXOZZtwBkiXmW9VKP2wPSQQ5FeCTlUqxaxWAeCR55BfXQdN9MtchHiTwRtFkkX
IzKAsLuNtJBpw07neu3uoLFCVWQQWX3HBgGwlkVive4BxL4rkOoGruJkWji6C5AWTWPabkJDAliq
VAsSa4x/8oLnJ7CYPP6jkVEBUlH3GzHNcSvTxDQW687JwTLYbkMEO9ZrbJ+x2NyJ1K/TLLevYeDP
9xM52eadcwM6WlqKSeLDORhZeSAFYQaUfD2CSrhOQtk1QpQMsDSj55tzLC//5Ya/DJSqAz0bTqHu
JROJ4eK4JaOeSWcqNTUE+tADsisZ842O2I/elI5mzm7lOdv1fR1Y460TF/RGHZqZWpKPUFFHlnla
JJXUZYVvuKoZVUBc+GpA49/u0yN5gTOLIyhyHX4LCaFsDa4VL7+xg2FvvHVNDGSJER9o5UhouMgI
O6O/0RWtsD9gqrvahlihBFWKb22Y0ngVALpx1dYqYXBCvs3GyWWDOdtSTGqH9BTlS07ypFucy0Uh
Le1u+tgYJKvs0T8dgGyhMqGK/evFMSBFMnyDZ3GLjOm0ZnX4wTX7HHfRgHUCioyoG9SiekLp2lva
B0VUxVnuWo+bVlhXccqvfxGcsX3YfXZThXN/lNvgOj0NdO8YGl2qdwv2GMc5Sqs+NSF+l/ckQERS
s4/1yX9IMh1t8nw/U50u7TUC2r1ctUGDTUv9VMoNXr/2EsXevAuRj3tOvclVRMwOx+2Lv+aw0sQr
ka3CaW+IqwuUqsYNVwXVOa7ok2rv8HoRjukzde1VmkenAfpg364gT/3GHeOTrpThdpxExiP45aIW
h1/z/CUUZ/7L9ehKK+N7XnJpbgbA16oyKqEY7ENA+NR+O5g5dosffMyiWLp4kiUfr4qzhGHoRjLh
7Dg9ntnfAV5xbvc1Nt5as9TGOCckR8NS1jvh3gNxGYelELXzdMDACEvtT2lA0h3oirAzOiEsedNc
O9QaaNh3MeEC4pnJxF1YGJ3kcrS3/FRy//oNxq2ojcKMutZPWRQjsdqTLzyuxo9ZtsvzUHcGvQh2
jCGwBy/dTuvti+azOgF5t3PPawZ88s+pPLIb1g5kG6xO2Vn5K2AIwA9LsY4SFRA1RpgmcMud5XPU
raULyFl4Hogvl1iAbofNRMJHI0B5c7k8piWhsVtJH20ZSc0p/j0nEIQjdPjClLD4Aa+cMqSQjC7V
d2S5GA566r2Bs5TzjF8l5wmymPI6hIgQ8vZbpy32TCtjJNqYw+pGz1xLW7wKsejpF0CgmhshLo9W
aS33nOjKHLEf9oWHGt2xXRpa2GmWjK/0WVQ+rWdHzlNsTvbMt3u28+T4pbYHlQy5qS4uOcGXBfon
e4uhfVk+tcQadQlaBbA5D16i1lrqFyB2D9mAxC2WNvFwH7x/oBDNBMowaD6T6KCc2P46U71bP/l8
Ga7icC3I0hflMqZrE354Dx3br1NJQR/trYKQUm/u2yNErZbrj3YHAPfWC7SrtUL9DL25Yz1e1uRO
PGx1J1+PJcCnTIZgIL9WgBZ3qMggklbIHO6U5gZ0pWWGaqAZLKYyZ07k1xGGk8hssbURZBrxe6Y8
SajJewUnJhp0jjsGTFC9BgxLzztHbcaKDozQN1tKDJ/4mCXa6OmvsJGFKF4URI0ajX7OeUODvvno
j9ZK7ez0YgXF+uY+UZDOy4r0d+A0Bnn3Jb3cp8Zakh34QwIRlIAd1UEd/G5pKuEbZRjWBUJBd0zk
lfJerAuIbBc5EkcsJ7rjS9/ktuaosMLXrYxGttBoAr2b1LkI6gnsN9/HXZdIwSedtKVYwiZFrSXG
I9d7gneUmPWyLfzEacdOyq0fyOQuACrvF6b4mwzEDmx3aT5eBDeR3zIyc65Z+L/D20NxSzcYiVMQ
XCHvq64OtygTGXQQEI26nDZ7ReNGg0xbKEQzvhOL5MwWL2EBMBrL9rthK7cHgUK0xrAROH0EwG/k
JKdl4LNjQ/KjDt7CpqyDT63Ye/O9SFcmimNrsVQJDSOWR8agrv1hKifEA/hZUSDIxVUdGEzykMj2
Jl7K66AgcyzqxrPKMEmb7UjDh92O3DPCcITodcM0xoPJ8CDPGIi7thp3hvDaB8EMtPYOvbUvjCOd
gsvXDTPqGaxkV3Sz2IjJXzvgHgOXi0RZjUk0HlxN8EUNsAgkpXawVS/49F5AS/iDiJUnRGVnfSzi
EMcJJ7CEQ6cDa6AAmyDq7nyq03zAgDHGCG5FsbzzoxJbsSZ/t9NdloPucY9OZke30Mo7X1f2YUW6
1LupLv2AhtjJNj8edJN0E506a53Y8s+KGTzn+IOJSgr0fPLf4voQDEPYckGZMsQ/6bYGpMNPM/x7
jek1Trwzn7gbGjgfjpm+7V+ZtCNWfXI+1gGGVUmdxGQWRHpMJXtEUKmssRjscDWlwCI7eQ1EXE/B
7Zh+3Ab0/w+bN/053Or48CWcpIvvMkpEqBXuSn3d7a/Dp9P+W9n9mvZdE4GAfT6A28bgbO4BPjQD
gjRASJ1MhmhtZ82Kuuz0MBKB3yWrwayZt0Si7ZO0ya+6FlhSn9MEzNe1u7t2H7ao5tELTUpbn6NP
8/pUyco5/eJAf7qJmVMy5JKBXJ+yPQU88vzIbaw8IbB94FlO1vXCFHnVXBw+tr6Q/2tLiZWy69HP
9/+6V9g/HcddMpu3l/uNt659OyDG5jEHuFEWMNbe2vaoplvVmqzabQeeSCnIZbfDX8Bk7VkmEF3F
v/rgr1EWPTrj0zZDPkADtgugm6m/s7rYZ1y6TvEH7O5qI9vB6IdThw6aRqmLhfKVKbFk9u+nu96Z
W1nebRRf8QrJcKruemQZnB8HCB9w2WEs1ArL2o8j8ZOKQ17Ydc0pLnNkmA0lLsqQ+4kzdgTEIBRa
jy6Kcgemq8tfB1zXc+FnSep6PNACZcG5arQn6FB2hxbU8OsfdwbBSxmu4uSMXGMQ4Tb4IkVkkh3R
tSrvjOSs5Uo+Qwzd1ERcsbjc/l42huKmNJ8o1JSX1M/QkMaxMz2/hsj8gT4RGpFHBVxIkjJ1nYwy
sbtBAUB2pBemupHHHHerOWtLYLbWvsz2d+4a/qyJCVPjxJEiJyexS9cVhHS/lDGMEeai38ycraWv
llrLxZYfw9qN1rqjUQ+DzuiEz2xP9CaEU8w+6fwaSY4XKBEvvn4gubA1AbJpMLkXYaaof4ysDa1O
sNbPTXcbkyoYoaH4pweYA5cDmDHkmgsc5/xoFRYfdfNYZvZ4e6aQ+KNUbS6yeKfXduj7NvOFEhCP
YtHGvvH2lRCsDjCcPiL1siU+EnpEmdGX6V7Hdi38kQ4Y7FR+l3uUVdzsb9K0tOMykBuzmXHzXso8
6d71dtBeSh0l10UtImtCw6jhmScOx+th6w/J5xk39WbWEAG2A8OzfPQGQEv1p+WHHBWzV2EOTC83
FeoVWq6adMEC3EPffIG70mf4sO7uNHAKRacSge/rMj7uA3RUgsxmUSzt9rp0BFlz/JFX3GArVOpj
hpl35/Wtm1qNOIo/RvsMcvupvzOCed1v/kDYt77wI0cfR2S7YONHKAINxZjCh7wy7bY/HYlLfRxO
XgWTZ/yyj5pJ5QcjjRqUrCLucvFPsS/JLMyYusroWmGJz8ePF+HulTfryZEHN3e8D6de/UV30pVk
rREWFUzzKcbTQ3Sx6ShH9mFKoj99+Ak2K8dn/IiWBqP9bnxGD1gBYizGwMhfE8cmUT+EAl3xOfjl
HRyM3SlsubkpDHWlL1lNPl1EwHz7HZLxcgwL0zYSzJIDTPYYp3ocRQU01rJd6EG8QfQQDLubwJiU
aTIh1iUC6aeQtkOp5iMbEmPi45WJ6+ijDglTEKnVhL08cG7l7pD0fkmh2G2fXClo0L42p64gVRAX
vFr6XX6Y3Pzf6BecDnEgd73TfcNmxJ6OTM44XruhuY7YDy0LtLXbZ5g/XW350L+VJNHHpdON1MRu
oLX3nSSfm1w2IH4DtenoDIYifLuXsn+ofceFsr9jT4TG1KIfQ8XwOyaQqIx4xWusoR3/7OR3sQqH
ckPsl177TANnT0UCRg9Bjmz1FGg9FJSX2gs3cqUCocaM8rcGt6HUc1Mj92F4TZdBERTWcWTVd0EG
cN0b29dj0jZuDk7MQCH/pcFsyrw1/q19MJtBv4+xjhT7PdSGKjUYVWz8+58TE1EIKHtCcBhBc/Ub
9+ZOh8U4PlcK2yEeaxbrek5tSViDeBeGPafF9XtJxQVXeCFLFW81E2TXRIEsK4OZ1Nya6fyNp/j6
JBkku5kFU+LaWgDqkaAuD17VU0fnxLC7lj//HDLQ22sZAvVkAMiMgB2mQTDysGnLAGYAiuvB2RCq
7abAqir/67goPO9d20r0FCPCL78BEkqBhdYf/JvIVw6P5Cdw+0EBQtxbvBLcTv8zyVx5QZO9jLF1
xsCrXym6MKoZ5vWmoiEA7y0KahKtkltOw/y3wD/VlSvOfnPr7vPpbHIhSqd91yql1QthE8elNCcQ
y64ehn5UNihY4qotLLd3l1Y/4MLYOt7j74lkrsDT+Mci2MT+0xiQ4yr+5RUwPc4tTQ0cnh1SFBLg
iHLWD2N9UWqnFmS2yDRQ5v1hJN1zQPMDTLqfyE/20LuPK89ALyCz7R6lstGD/+7vJb1ZWLeRD91p
EWjq0ewIfhYmONcbYovxMtAKgiSXaVnWh68KnZHeF/XiMryKN/UcXOih9n/AfXvtv0V0GBLw1mBL
0+zuxUyXUClJG9rp9PSOJ7DII+J/nUcXvSS8Q+pRig51PmkM79n+ihk6O+TOJzNenJy+AjqMySN3
S69mYU1QleHKkju/HfEOTySrUNOBqHnKBIPzNC4GuWfZ5cFcTsHVy4Jr4xZNbwUxkUODQJKOZHll
86pjQsrNjvkParZ4Dco4bV8kBdKovRfgcNW6VziacDtGhzeWOuwYh/UHoXCnJnEj6+LvoCA2hgZA
A47LbKOQCJSmlSFkrW/RURgqBhRLAi3bk3cLcRP2TxWpOQO34uxAZMF1J353f1bl90RKnLx2MP9q
DipjrhK/x8QYq3L30J7U5KFauEu/EfiVDbV/ttENVqsglDVZKA2HCcQOSkW4UTp2c1xl4X13cENN
3d6WrVZN3HesNKszzvxftw11JpxEsKoP7s581UIvUlWEIV0P5EVQnhBmqmUcderBwaLPSP1K2C2K
5u4nypyWxljci65tc5t7gcCISwnX65YiuLeKgJ4u+/RK2129jvuu37eDMcia8UfGOzeTWgEx9TNf
yXkaz0ANrsQCVEP2LRKzBsX5q3dBWqacbz1NpnRdaqedZ0tWHig4saXREVjI/nDw8y359gmUySF8
QkaSZe0hw55i4unz9udb6CLdeWbEvdNO8vnShNU3FuesnOtOb32WlXRU5OA81Mq6Jm6WnvW37TAV
qcZFYRfXPZNbiCzbvJqc64pEiZFAQlAAvchVouCqwTQjiYUYApU4cpcrpi8Nec0k/AGgyL4kK5Wv
kKZJVnzr6sJhENYGJqj7T+gG/4e5J7QBHjvhw2E+/H/8/D0iEqHUsiI6hjU+kfEyymJTa0tVHYeF
vyrxhHqJoXuZgStX3MFdA5+5awqtPb7ePr5gSthyhkNGx2Dh+znGCByA+vVjDXzPeA3MqcjBeaue
gXbrWioK/0gGe6MfxrwUYuj2N/nePDhrzTgwWl428877XsAxy1UoeStrYDltKk1BJWRaSpqgX9Ys
MkmrwQ0WRL3WjnO05XmyyIo3+4p0TfT7grCn+mKf166mLTkUyeAvEcJ2N7f64uEOdJDkHRBijcrw
A4v7DKy3MwDMV09J2Tf9zFU4ADgmHzIKI3X3geWtfeV2rI51OPdxIMykMo0dvPN0q0v+Vr+ml/UM
lmcpch+H6IjHOxWRTgCiZ3SCIG1EPRd1Y57f29EMBZTN2VjucSqlFFggHn9FAarVLljWsckRjHU+
30pL6CfB5ziKXqFPLzXrgzF9F+USsD/A2tuVo54sep+TDpObZI2WDqgoJOu67kxX9uYeadt6QFBy
iE0BN/g9Mij7j59ZKIQiZVDUEUdtBL1kwb7/YXAwcdq2tosZiemzrECKL0vxh6QKyJcbhu1FUFM5
YTDvVBfh4WNA1M/cZUL9YUl7dbED8DD/xbtNaHaxZqwk0SIdkXq73X/hPGYTwu8rPkrHVczISpCX
U4XO7g9UwAZav1gipSDAKjHYWdasJmC7F1tyvyY5hLk95N1/E+LhLs8JYOPTYk22sC+J7jnnLiKB
klehJBZ9Ll5bmh27lQ9A/Ewr6qzZOYI5fqE88RqlA9vSEmfSXa3S0CqN99VsIar56gOCs1LDiJIb
wWeiIculM8ZYLuZai8CBmfwMaL4c1AdLGTMsnTZUOlVDkTufMlHoP7AWDFM1fxpW8UYOYoAW4LFH
GRCYv6gcgPrmKg5xu3bJoUTW7e1+k55QAyFltsXLYSaN4RYwPqYCmYVaWPaxLJvQYLPFeDgt/UtM
xMim8KW75D/4BYV3Y2AKF7FVOO1hcs1+bDBKE+DZn0kkz4f0DS1muqa1NazxospYvetKilPPtRRu
X8DeSR3c2jYISBn/VgYPXY6waA83RErBGMdVk/yIYKcxkh2ik+K6xFcqXo6sgwceJpY2M2YGVbly
O0/HNYsJLK9e8/hVtIjYUeb5rATmonkMQLZaxattLA4zc/94PcHemRD2bjFzI9PJx4p3EdBn7jOJ
TvqtRemwXJMXleeU0+0s6YtUiN4jZhWMBp3ZTMZJFL9MJQxw2T//OIuy0xf81WyXZSZ2/YDcp/P+
VWACwmEosnzzkAnolKSjjrdXCLHXueGgrGQ3rewRb5j+eCZvd+r/C9q7mPGbJqWUDuGgLZyIWXS/
E6WeJCzhmb8GabTLlRFxctMP2YHZW9PhUXBuQZGZx+cRS3Tu5gUqYWiXN/wWPA8ROEt3xcrMHwxp
/NRHIpqYFREXuzHTB51oJBIkOKTUTqD1CKAllLxETLTun3cn3Fp0xGXDRWsXvZS/ZBUsHdJo7FqO
N7CPwHWrtivR5g2mgGw1gVK3ygQ+iYwsrv9qInQXJEyyHkaX8JcYdc1+EDo4AYTl4EFxL0LNB6g5
VjznoBX0hv1aO32h6P87PHfY2xX8Ok9d8YonYdwUxKsyD4RCgeinmOVz+0CPtwB4npY4r3YqKmTW
1W8H4NOTeVURPb/vFaSsso0J0Db1cX8mKPXVtMddKs+Y9vcSq+eh4fbTym4lcmXget26BE8TeSLJ
V2Uh2h5LnT+fOzXtAT7t4ADzC8+5TaKRT6oQ6SYtavgpfxgInvHpk2OIYPrDWOjTBw9sQDBXT6S4
m12odbOtxxyqO2fLsSDIwyORVwFNGGiQOR6x8nc4U2SEWc8g5pwZs6tBfqUVGsD0hOkAAbiHRx2p
2hPdksePCm7HBABYfRIWCkRt0/HvDzijAkKOaIqfsMQWa35ciBrIF0395Qdw9ZKt8kfucGhe8hOi
9ggD4WQOInDWfAPCp4mDcDvs/mBiJy44rOArphnca1ZFhYpaoLrvMZI6OrjqZ3Xeu3hAZekte6CQ
1+lKrO73rrZ6MipnQ5W0aKLdwtymP35NZufb4myxzhHe75W2cNWtFQ52gkBpurbcpJHVtmVeH0GS
w4nL1cQLf3WhCJdwKj5ELt6DKGFeS/0nmcnCPXkWSbNhCKYqUevHpnpcMHRYiKUB3oMZrK6GKdj/
6Squj62yKS5wPCBY/MgsQERLFRafwbt+BTBJC/LkeFskLfwI31iz92Vt47FGhfTbl34CGty0/WFh
z+V+RbfPUXbNjI7IS/k/kxMoWlYBay84N4AXfFpuN4lGHYOogyryXsy/GvVnULmHrIg0JgCtW4qv
oh+/9xDmbLgmU/dGM/UGlNRgnLmTxfESLq2XnfD26yiS6X2WJJUcPTvwLn7gKr/+Mt1rCeO9LZxO
pqlzBWai8T3vIsF7hjy35ue1D1p0B9z2KRgR3KWxj4NEzURab6KbyRI00zLAOhxuXzz5YmMaq3s=
`pragma protect end_protected
