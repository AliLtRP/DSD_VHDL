// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U/eXMq0aqaVn1mUHqYIkEFWa4rYhSHUTb/nF5pv1cyKlOg96Tehh/A7bbFUhtso9
iZ3WI3edE4L8Z6uJRjEAbV1f19Fddc6ZH8op2/4rtnBAbOC1zKmW9C0x/mbLx1o7
1ue2Ro/D3c3ia4Cd4KmLkeLLoa6j5xzalXg2i4Y3oaQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5136)
LwKV9dTt+cu9IPoJQsG5ZFgOMsa3a7723MVo45rVSM5q8xwJCsuWa2SdngvlrIkh
zHgxWn+mLCcO4HAVfBjRKMkNSQe3x6pmZp15aEfIPO2OMB6gsJVaE4kieI7PYAzs
IrGnbUhKJgfrjVWN8gURPkfgVWmJlf4uQ1wKTQhAAJ30s0dJFTPo23HWhRow0n41
NKdUZwaKxca90WONKeQ+abvB1O8fZyGFbGFXQCmjlWDNigDwCX+XTKTT2qJloiuo
7hS2t6a6nv+W8MPLQEa+kNFY1Oz5nulntEbufI6pN1egmM/fWQ52eQ0nxFdZjlrp
fw6s859DN9Vv+fKZhOri5Cgk3tWDCM76k6MPd/R7HPE13hCG0Z0NyRtZiMuhhF4H
FmNUNGul8NL1qr/eZ3g8FpA2DLO8QZNSm33u17062JHT4lvukB8MZ+xdrIYtAjrx
pe7o5ZmS+NtdCZHiL4XnosIImFgQ/Zo5gRYbPOCKFsvqz6jODwDtSHuCfihiiwVj
iEEKMSNeO/t9NeGleM1BVoUtBU/ihlrIaDfGT+0IruyYPtZF5k0mcv6tVefyt5qj
qFkxl/1KjJtdShEfMadDI6BmallCSvp/9FUqnd69icumXaktOfZQx/C61ecKUxfd
qWfcxVXMsX4WeLkM3mtZ3DD0RG7DK5kMlZq5AcAH6g/OWFbhHxoDw9G/X4ZxtKJy
0KQzETcNXbiLZ/zoMzFEtd/STd2Ph4fDI9yhuS9pmJQXd4DZ29q4w0L6nIuGfvWp
mYpIfzI1bPE/FiAa1Pn+EeZZ0z5an+fCzwqUjj3L33zKKeBzeyYi9HRoqcYQOsb8
oMyJwd8C5jvN/3GyDPFdUKoU+Ix2e9dUOsCn4BXZwKOo/3pqCZRMwkd8FDYkhU+O
BevUTogRjBLDs5gEiwNJHpZsUEtNK2jwJQ3mAM845bdDs+Dgf0IfmVIYCzAghYVK
6EqJLjJu93YJw4cl0QUv/cn7aAlaT11KzvLfgkqY11PZyUGEj90JryKA66qBDspY
uu9sP06J4SLW1jl+OzWEvYaesrMmflONq72+giuEKM1oDcW/F7lKXdg5Km+BVcRc
WJbU2bIkYK5VuTFa4j9yr8dVhWIxt9M3igzyKYzboi4GSGIUmMpKN+GxJp8ItPAD
ENMlcQExWUdXjV/0aNd+lLOQjyCoe0WO9rXVxbqDrk84OVIdkckQMpj3EFIN80V2
j71p4q9ck4cPjjDiWikBWbGfa3FrW4JfPGXvXiGL/1tPEJmOOGaTpewkj65v16Sc
aPoeTAKCGdp1STc9YEDi+7Km1Lyfx+KJktpjcjc63eWk6S5ZewgBTsq07CCyd4XV
33vWR/NETUQG0tI2PnLa4J0jChAl/Ef8T0LcvotW5rAaGFBK7tQMArM1MVhY37ig
E5MrfhE+naOAqfkmr7+Omm07q6x6JK9lA5wMz9ThIHDImVMCZQE7gXyVsTVaC1qz
ULhu7dd3mLIW4BAvN7/mf7Co7yzeJQeH4xur49x6rXP6bRvR13SLx0f3cKvg/arl
EGnBPb9awKJJZBsgKcz+ffZzmt+qd94zObk1YyHMWUGdUIEaa5hisMmRo5uqIvdV
cTqmVJb2lNRvzRhzJnbinkRzQ3lDiHivnk08EGfa5un8JuGXVqNNxKELiZTtyTmt
KAvd0P4muboKV+E6T6B69Rp4VLz5r7rDj0xDjTJXb2mYzCaPF/Z/pTG+xUJvV1L/
hKWRmPPabTySqBHP9Uxb+BasTKKddYyYMGPdm7DBN8dFWSzfUhhluBhsoaNhIKRQ
YO7LiAaLtxslQCQLhxKAJr49KLoXcoZ7Uf8WJ6yi2+Xg7inDKgCIUXP8OGHeb4Fw
fXnFYpFDw/4Ya47JSxqzGGjIZGOaQeDtCtZ+HR8MYelQBJGQXUt9IwuoJksNT6ta
AKh0ng2GgxtfBw3OCU8Zph5Xba6dEjrtrt7YRBhsHRcZ+yXlExlrtWFpHKNoZ9qk
+ga8otc2jkm2sTpRVarOtYeX6wK+kI1dRiF+VT5e0guCNI49GZR59qLvbXSvAZDW
Vow1iNp9vHGSAT327Dmc6opIFZkVB15LwLiErjTVjmp2vHOf1kHTzSXsIe18m8kB
3U5g11LwDWfitW0/lINGVfqA9yR1Mb+y5rI/XrPldc0tMHm9c/QzQIaZNRLG3FrN
dCBPeL4xZADMcVr8OJWBwvmdpl7mo1mJhANVVjNa5m4XyXF8/wox3PjkOEbvZzuE
mYLHVK66+9oBk8ee7BPNaSKVrNIqfhgSMGRKntFCHPGzYzz8Ee5qv80yMQ2mjE3C
UulA/H8n14fs9XZ/v51xgk65tpPRMgh/jm3MzLDo74KibQSP8Vcc1KLcLecUZhqj
8QWq8PgMjh+fsCJ4z6jN3tOV4MELaghs+uerAlfZDqeNJIP7QneWL+zpQKyF0dqv
4L5pLIX5XKDBP4TOv8/GEbrXAJjQG/pbXnUW8TA550xI0i7DGlYmJqPpDy82SyEo
8JZpABMmO5phY82EIGvvHRZDeffI4gPSqwGBO39hamkHgfE5idec0hKx3Gz5M8VT
COg/RwcKG9KFpvD0T6Oef3Ubby+a7SYiezhzzruCFVHr27Hge7KGyT3wGln4CtrF
xTfJM2RW8rH59qkpQEBu/mGipjMl1iQ/UAnRcxrwP4/AUgZH9JUU5H131nFKCT1K
gMD26PqX4nwaw5F0xBtXMmBhv0JTuA2Ori1MTbkbeNaZPU1UnhKK+uyvwB0Uiogy
pO6053Yi2C+1A+a8EmxqUifOVr2NzARyUghykieh056sfBbV5AcWRQ4sq4q+eJQH
NWBsceTX+sIJTHgbBRWXhvxy5q+ldgNPp6WiQFn72cWSYW4d+9aXFcLxsIbE4zJX
5XoVHir9VVE0MKDSRfQoez7kdgy4SmSKQBQNPxpEUaculyaMrI7SrWh1A3T/FenZ
u6/myUZPU6Y9ALjfIkxRE/Fk6EQOsZANhh5rgPN2guo85MnUb48nBL0yQgKcT9mg
XG/rODhgFPDUFNhKJhOB6De37ezP3snYz0c9piiNd5xwNSDZ19OAz5vBcNucxIwr
WoE+kk8prVnpjmj86C+Glb7mQcCarx8WPNKNVR5Bqc+puCGFP5ni0cfAtBc8hO/s
FcUCRcA6GhXPesEEe/o/fh3DVSd80eNe9HXNHmY4gU0+ZEt+LodseNg74kzULH6q
VWm0pBI531lmBJL8sglUmKJw8Zjs0rpkwd20tGyDOEFvGvkmCZd7oI9D0ELzgiY2
TN/1ZWLq83q9eHs2kTytICiLza66dD/U7taV0nv21U9zDVlBKgWKwbYDA1FUaNkQ
Q8VUW11kjinAWs6xgh9cIXV+lX96iKdmMATA9TU5H7lgoteLxezpi2tz9qVpNmWL
/bcOgIm7ey9mvbnbwU7HwGkSlo23WWXpC+lKZRYOJsCv33OkQ5SgoNwAgc7G16cU
plLrE/W7yYIKebziRDqV66cGgyqSCk7+MEciOdZOkcu0Q1jzORIADHV9rrYVC6gq
1TE05yWEqHc7a2rxDbm9+5DyXJHkXkjI8GvrUcVZvL03IajQfdOUDloe3ZR8LcCg
9z1HNcK1LajO8iGtdswVOCLlTZKm1QI5lTsnGk+AEorDqamsiH1n4OlRi+rQzm0y
WWOkfBk1gSZcMPIMOnsDzhT9uI6Hre42b0fVRbyY7ZtUWJ4fmzPxQVhK8snG4R29
Ru6of1guieRk9kYfH2mcOuDkPP9Gk7vcg/lMZCF/U9QuuT1UAxywmuyK0FWayf90
PO32RFcPY0T+8/b8HR8rRdakUbBPw/hmsWFQy6M3yyyS+577Dc3FLq2PaaOdwoR/
WCELAv2NgXM/AbmZOTOTtoNYFLMYAF4O2uKmxKqPU0FI+rhtzusa1eiLZsFOT9tg
E1qWroROVTb/3JHgYhxbKPdzguVR5BdXzrPd3jK2ovFdciN47B2m7C/l9dzolL4c
OgPkn5jBupG84qev98fFUllbnErq4amp+Ad23sHbpHIhQtcXYZjGXI+qXAJoMwCi
a+z0ekV4dOeI8XhKb37E3QsCF+PhJQZq//y2BGdu2EbFEYAb0JzeR0l1y+XR3bcp
8Q5CX0kTk64HCwv80JeJ0pz7bpQZZCNu1OPRmLyR1vIxCDAtH50WhnMnjn6zk+8R
qd3Pwv1vgTGdLKneiT1v+YhNIIs8Yh1tJu2GgM36pxmlbaEH4DH1YIk9fQ07gQXJ
zcto9cZnTWrdg/tdCwNkeQc2LtcEpOtGE8MOlhxwrx2yBL135LIg/F6RmI8vvNNl
DrC6xC62fUrUsOopipSAxDNy7P/PeMH6s4nBA1OMNZkQSgFPRP7LdIKY/NMZ30hp
+atVZgXcX6LusvS8gJRJ6duhL7JQFY/LMfUH5ozQb9uhkULQ0dmsMzo9FvsKGfkm
tOIsUPDXrfiiYUrhuSLMkCl8U6bHLkC7KtOuyvG9ZWYHCT6q+uipAhQ0iv50aqlF
PE4bC4mji3kJlqIM3p0tK59xn4G/vhu+f1KkyafleDaf3s2xGN1yvaEbcUvypkc4
3OOnNZAImS9ulGr+vluk7N/iB96YgAy2FxPE/qo9tVitsjoqfIsD0t0dAMODqun4
1wl8MFC+yVtZbWztB/IfoaVsTj2FPKzC7PhL9GDh4/RiBIuYT4Rqlbm25wxgetcS
G2JrBj58xxIfGYzdEPj5f6v+qJDkyrdr3/n1pU4QrgfKqw7MZF8o020ujkhwObpa
XlIb3NHqLpwHoLqY3npOeN3R8OOXK5bGm3xv8vIyahDfe8XUYzIOLHC4hEVIaTh5
9iflN8o/WRKcQq4R6maOAhZQUS1N3IFGeC5pJ7aqe5B5W3sv/N1edh7E/toTeihd
9RW/aXpcrfehObsvp6PnzpQHWMq9vujKVsmv+dtLFun6OemgPaMczAu6y5c3jI25
v7DqlqvBEbYOu7f6KPTi1gTmHYxpWJK6BouRqwLxN+NkWROpkHaH4y2L3CaQZoDJ
CoC2Rst9tqEXhSPZU6TCX2/kUyusDZ/mKubhHTLQROGP4aJLzdS5kBF7qZNDCzLO
8IiE2aQavXDG7G9ZErHptCic/5fsi6wF6Z+LOnapme1ZNv6hRmrs8E9OXWrSpIPP
4dv6Ecl0wPrKPu4pGr1wh8ZWAe9tHJhZBlZ55L2nMOMcH+bbAcTOnuNyfNcA5Tu0
gpMOvEZz1zbtl4ReQjN7/Ou+tzw93Vu/mQBdswo8Gmp/F5dWtOSaeZBYM7R8UGdZ
jytuzROR4q3mJbBezNJ8X73lZ1YWsGTyJQtIyHj1z65Zvm79gghgCeEH1AuzZReo
znuMNum4/Zm9rW30dhut4bRePN9qp+FHG6tDsNkYVjRt9EFZDYo9U74IzGEqvuU/
ECX1BhSFgxjEEyXDa+WTIavA2gzR+y2NP+sN+SjVcdaa/2ODXSyZwCFWjY2cksdu
n3S2bkXF9Toz68tOM5Tgoy3QRFdPVqSoSnTPn2x1Ue4IOfV6DYLIXvaFGwTPPRLc
0HJu0jhTDVOxwGX4uCa0IL/nvTf+8vtyElEnlO0s8CPEeUQs3JmycCW5VM7YPhqn
CZg6wWnQ4s5Np9kLpGQz560336gW0c8mxoliXZbvUWYudXBDQQ+vw+DalgSL/Ur+
5l7yPRmfEDXC7B8kiqLxJUBr5oYNi4nHmrV5TqxxBr3MdWE/HGqfz8RlKwbcbEPM
GSwaAnPBpdTUo6GZVh/t61BSut7HXc76niUXE10qZpWb4EiCilUtVKiziuhWRciE
e4FYp4bepT+L6SVy7hHNBSD87wLUkKm0NA5b7Wx0fociY1Cd7cOPNs8spjTtf9xj
+taMeDv3KwEYgZAoN58cnJLZyqSoTT/u0FHY4XKgFzpTSszwbLXW/k0/q0QfeNUF
7IRJbvi2uyWoTRsEJM1YCdMoN1OjtMggmEUCQn3eCEXLV5bAxN2vPHiHd3sDaZzA
oop2VKMi6vLfCN6CS1GHAFh1JjDi09Z12S8GPkEGit3RrTRKDNgZ4mi2y96gZdsM
6CaYHVH25yFDzaz9AfwJxxYbU6XloUv8qogwmsHB3gJB5KNyIPcwY2iNhPzqxneh
OiI2vxV0ghAayq8u0D6HVvkRZZ1zJhAmVDBigLz6S0SAASzRC2P6aaS/ObHVFEaR
5jxNTKXV0CEfO0ZI0DnW49+Vme8DWT7cLnM3aLQ47KV0aUmb5KcfpCIxgVTWlX8M
lI/ODUi2pCM8RxYMnQ9rUbm1VCGmyVBLJddYv1Wr/QzxWAQnFb5NUr0QkH6fopQO
/RV4AUsIVBVLSIfsNbelZOZKGqUTpRxgQr2HQP9tJ5cRBUuFDvI/Z2ngm4zQMmcK
91PB5PV6olMZz2TZsR1Jen3b9uM3RybBIFfdf2Eg/WjyzDIPsCl/1NqBOMencMTP
3OqQcFKaXsdJI/xlAN9f302idWt23eS3P/qOoydQc6rc9ik2jNfW5iJX10TsbWdD
xSocm4TWcfjqM9KgkHaikSQ9hEF+XpmpWostzODp3pKD/FK89elMH4mAll5OaVsa
mFD2f/vw7MZ/i3ecB0WiFjgvT9nHqoLCxMmlVFDdC8O8UJw39LBYDRVgvo881D3T
tZOSr+5tCFI5+sWBYNakCtE0Gtwc8XRCbc4bNm+89qxn/ExszgmUPKwgk5VzMWdE
eRssBey4OgCqO0MsWBSmY7HubQTQP+mX3QeYsNsbsmDt8Kim1mmbo8KAi51nnueh
pdBz4KlRh12M4MLwQtB1OD0TYHopCHiouk/SpWYaPtM+eyXkBDq1H+ay5Mieo8e9
+ZvA2C1GjSycqb2gARQF2yjFnmyZTA+Dufj7glCaypmGr1i+lKRfy18HTwJosM3m
`pragma protect end_protected
