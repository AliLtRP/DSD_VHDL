// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DtluKUYvIq8IC867Os/P+WUmmw+8HgO8ret8YUQLe1EAwGXMIHRhFFb6AcU4hAu/
MGO1Tl59w9yOvUFTPcIR97aUaoasgngL3lZQ8kyLkuMztv0D7i3Ta6p/kUSxSHr8
5xywSkLAVIwLl8O1YCI50POcf7k21l7JyscksNS7fQ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8064)
C1uQ1FEV/oLIhGsDem0DvOuqjTx/Eu0GOaR1INnpWQ2SNT+eXMTaR8LyQI0xiNUF
AiCmSCvpm1MkM1wKaETVdniBvfZqNe3D0Fjj0CRN4YU5XD958A5GrXs6+1ERxCCI
UQfZas0Uqf+MJFCcgzAGyWIbk+ZVqkm/m70/PXMdHN4sWd+0BFn1A+H1qXc7UC1b
mNc0sJgrlXWsfsoZC3Iqi9MaNgAzsUpQ3e/GmVi6Ah13Leeh1J5TwLLpd/TmYvYl
WJvrpjCGlQ+fWuvXqi8icctd/VQkUSwhH73oYR/uWsjde6p7UggB00RJ4zne7D7P
LNqkmjk4Uy9jWOJDur1pIbhpuROeHZrlWgSAGKa9NtYmcAU71OgKPKFrMs7XY9bc
+OLxS1U2dQ7dlcKS0Rq8DrQ49xpDRBun8CbKBcnD6TpZ/fX1oyWJnKQbfLJ4Fizx
4krlM3EMACr9l/K223G5fsHjEGHue2/9q/vo7cccSUib3uV2r8Sub4gUTWy8p3R7
TDFny+0JNAA9JpdF2fWnAcRM7yjwObkNmapqURmeF6+FdcbrOP1vRu/3BzIHtFpC
bWHG2fFddPAtZH/8nllgPpsSB8dbHVru3u3XdRrSfiC1VHEmPs6YQCRZuJON0B8n
XY1A5W+0M0Mf8A0zhQKyypsp27GKe+R4GTsvJXpnVs+fALbwdKh5uDzl++XAjooj
A7c0eI40qYXcxaSa4O11Z/1JEg1jfNTbQxw1VNWvpGQksE52jCP4SVFlKF+pYi7q
YA/Ey2psZiH5eHTi+OpkDOnJEtbXDj0KrghVb9G9O/SI5PZy5yMqJdFa+RfbjaJk
Va+cD1diN3s51R3AOno9qQ6fZr7AUd4nDiA7HPXL15x4sQBo5yeDKaeviH342b8C
UygVDjHN0DBIzAiGHltmJfTofIbDH3VUascurQzb9C+hNkudehYU9SdJGmQzmPF6
ky/8YWADvMbqihDyUIR8S5arIF2I3pVapPVkjRTtbJp+XMK4EZuQROWe335rNfQU
AK/nG95JoSgIy9buE0RZYQRJS9XtHeuKU1yX5MIjgOcsfmdei9hKgtL0w8yKikQV
27xxFUZbRcqhNCZL1dX7kjMevdTxKu76jKTFhprC6kq0H+7lLwjV5gT4xx3bJMe2
ODLm1gAJKo3VEyNm/puFILtUwximqGdzUp40WYhHtp3Mi9mPslOyedLwk4BUhCT/
lL71Nw8f53SEZis18GOTtTCnE2IRb+LD5z0elsGm/uVrHIw5dDiDr6Y90EmeTQ7c
sdtEqzP4A+ubt88cePo0h0HPqT9rdCRO0D6bifi1Uc4gNa8vdbhQziKhuaoRjeoN
yBPFtWN++TfYq6D49XEZjfxHnkOtNMOR6QFCGx++DkV1YY7gVVFWg6eoivpKgK6t
J/3i17qllE7xLqV1DoQqfquFTYhV8u9oT74g8M+acZUBpXOcLhjoq5zBfU5iFEMr
gRdGKXrtAp8SgRmxllghmjRhUf5IVxlGATqRFnrgyRS83Fz2qi2Jx8sRsp/cwLkD
q5CqQ6w6ZhEl42jIFg4En8Pqz4LI/7KPN1qBIENImL3+4m3C5aKkjZ9irjYBa/Dm
rYJWwIDsUwln/ozWi/goxke/l1hD7YGEMV6dtXFHcAz6HoX7xL1QGIhh9uyTr5g2
j7JgKuvr00IE+C2zqihKIvH9uvxZmGuu+5+wCpCZ+K73P3XdWOm3DrPZyf28AoLY
dgG23BbmOL58kKSgt+7zkUcSBzC3fBAVKKSueqrlR1VCVeoNM1FYbIUUcwNnzIW5
94taKibjVBE286Pgv1A/17+81c1sTmr5wbd0mYXOuIslCB2jUnH82VwYae4Kri7m
Z/9pbMGal9qnSbOO5wQLcyCNYWuTXwYMgznPW/SxriNss/v4rdSsaBojxuOKRqlm
8cbsgAx4wtHFXCkuKYnv8pvRUoDE5GuaXTttr1gXsCYqJJ3g8ir+Tfbfu9Gspg+l
gQev7Mqr8NmwmWca1Q/UEiG6b7DubcJlPw05WEuVgSTB789TD95KJDO/wf4IKOCe
FvGjuVXKq29cB/soAWWG3/cL/lyB1wgA7Xsp3Jf7EvybfEvK8myTFe0o8PN0Z+Yf
lFWmzpWlsrBeqmIWkXqskabnFJIrEbWkwt9ytKO5g+8WuL7+9ru8/684A8buO3yP
f4vnwLUTpYzA9KuLYzjCZrcLFUlNxfckz73kkij+/I2CLJc06dB3QPxxQdw1cBtj
N/6XeYtbmHffZvjQyWrhLc5cjU2kJx/DSB6ncCBqmyDCjLWlpg+RIKi4fROCHYoV
Pqdrn186/VeWwnNj2eitx1sK9rGqgrDz4cNYp0wUMTlSf/+Ajntugl5Dl0kEo/p9
LRQ5YUAStPNEw+HA37qOyN1n3F8RIMLm2ac1G8g7O6ADvrE1M1THbJ0Icbhho4xY
uBxEfjHAXr80bam8Ak0SmZ9pdvq5rv2BsS6oyP/tTow7XcX+/2fRhluOCWZsf0+b
dT8gvARa3hGUJWE60TZ5qwjDoUngsOm7prOUCIt1c4qW6Rh/ejrf1jt3EJuKX/Eq
QynmClKQDAN+ad+4Kbn+O7cCAtQ0iSFSKnJmGbTxDSDDoDEvlaQ4OVCSltI0DV5D
iNkp6bJE2KiSSlcvXbwK2hpk91DdWIHUqcNbCfaBakL5iBWEdRSucHXS1D0asEad
h+3z3yWnne5aqG7iK5IZeCipSGIhlSOXunZM6dgCfbpWO2v3AQ4ro1vFmxpapskn
+umKl9pn8mpbSpTU6KWZr99tPjtoGArVOm3qqZS/EYebmE5f80GqUfA687deIVLe
RnjvmUAVb54BnzA+UjodHUTYLQait6jWo2HzewYsZUkIAQ/laTslpEk9cQ/LmEsp
BeqjXNLQXINzS7E3ufedFVgpq6paMbA36/Cv0TErAL7TCEHaBQXyheks3sY5zKGp
dKGqEd5c3ARMXszxBMI8mNv8TOis+iR85rRrWqpoosqabmMwg5gdi1ykpIgriI3C
+3l5yizETsq5QHwpHJgnxqlHykCKcZNWD3XESRrS7EQnaeGTW58GZmL+ipJgDHFh
L+uyxAla2TeW5rCJvD048oN2ES1cSgX0PR0LkFSqNGjqUaylQoByrC7cdhxLBq2y
XbHyGqMSCKldjVM6tLIQMhM0DPWPYboB1Oc6u0vC1al4xUNFI6hpw1t3cWM0FL71
8wwnQUeWwQrGcNhW6ZPDP+4tjxbFUbteBSxzVeHcvul+1vC8SXKxUSg6/2ci6YhT
RvybVEDp7iTyvvIV7qHh7L7jZQSFsT5j7UpHkwWJRI25FoA/hlbjV+mOWv8bYTiK
du2LRaMsIOZFX5nerfXRSs74Fz4oqdxhklfdQOv6sQRafIsKupdESi+ST2PY0FrC
9It93F5Vw+mMICtqDmCkyesHc4DML9i4etpYROYrRACJR3QxmeFeWgbQvHdzM3GB
zGQoHcvZd1zxjlY59vHC1ae+LzF00bmNpnPq+dr3J75hXDNNATz7gQqolqLIT/fz
lY/vqN/0knfxZzVXxxwjsAeNWoByKvGuCWRyo0OovX5h0EVHJd3uTLEHMK2ZlPAb
P901AJU4hllxOJgg77CQrhhkcXmzWYqaamScfNJ4MvQhws0bSSeH1KZmk3wr9tw8
3Zrb+k5xiHwa9LACulKZGqhD1xWldQaLWzbzOfbVVaVAlxvxpTJN219gNb7o1Ldx
R4Bip3xT6SbCtHy8DJF430iAAIehKy8iuLbe7STAOrOf6SIwvtPWS4MnY4aEpwCy
vlqubBYShBlse6rzBauMVyO3wzhyyQOxrs6j9EWQDN/ct/AgHESUUiStQpucZdMp
Rumk8XdQ7bJ52o0d8vcL5zKKcr3674SYXSHNom7khgxe7gly3Sh+gozTmrDVYM6I
VtTFexEOLumR5nA5JPB+5noA5rh5WSue+Sf1ceyzx5fj4OcI26Lh/ZYBA3hPDxT5
8K6HkZsiLSiASUrby+gKcDiiHNR0MpjQ1wlkweKsOABYQ5aSM1MRj4vxrvoDHowA
oyWTRHqY65waZeqDDyhfvo6p8TTLw2jCFolYwS7o5L7cuh9XaqvzmfvgJZEjNEat
t3O5e6f5mmubCwhQi+30xK8CYHF2+PxDP5fnARpbZR1ezD/TKYlLlk5k5dYTQ5+C
u5mNHPTZSKHECxmZ7eiXmUIA19Jtp0kMchfcffRI2lCO4s/hLFFxSKYGv5YpNnoW
PuTenBDrLf90xnf0mvV/a0ZePNU6qaM7TDQKbgxIDTVNpiwqE8RY1CgFFfuoHRJe
2CEqpQPuYOC1Yn7VyopVsQAZ6yP/LJ0f7Itu0W+cxEqYUfTdA14ldKl3NMmY2UHX
mEjZZePWo4CymlIQn5hJ7HqsST+WPCD6nN0ddMHpuG+InDkxjdYbJsF+TEzF9XJX
ajy4X2QZCEM3nqekyq9RIkyOSVkzvjerineuc/UJgW/ZqFGY8PasylsgPxsTdTU5
JIVSCCTQd0hEExonSdC+57dgX/s6QHFFpRmLsA8NLRWbe1ImZD5qvxXndU8KWcpB
wiJzbrG+Q9Qq0hiFbTl8Cl88gw3I+5keSGyqmZ3hWN2wnW+rzLpWvY+fZPDnXD2J
8efIbm7VmW4fDwtdg0q202KO+Hw3/gfk5FBMxZOtwhGaheVw32zgLMqnZcckHEAT
j4wz0UCQZXXe+wPur7o7KzdoRRi5AGFOhuQAeKDintG1SXQdopRhhjf+dA3GUB3l
JrG162dHMCJ+2LGzq25OZ1+E62NiCXbLVDDnfXrnTE9pk0FnBu5loKQYHYvNj1AK
+717lonCu4hDQ+oH5uvaMX2RegZsLqLdvP63PUUTjF1srD/1MKAkEwWB8z4umpBI
yDcyL9uq9cm0COM5Bt7dsFw8xRmjNOxEvzVoLUMroyQrnFnfaTh7x9ppWb6c+aGn
+3Q/SiWbwoxxcPvhyxwaNtTOkEidKtbqLbM6t6Av8llh8DNwrhhmfyLDRVjXvZmW
+nG9ehnGn5xtmpdaedJnS7OxojKHq6YVBcGgL7t6R0kajBJyQs4ZUQ+l/CQkMt+r
zDRnUIf4BeTZ628c80Z+qWkepfEYA1w+fcM6W4nmjsYZo2MtZCVqEUN+LPrm4CG+
n1E7rMG2/WZp0Mud5pXPLQYfMb836gfvctA67CKkzs02zss9MiuH0KUguiocGqEo
zv1DMi7uNww9lH8RYzXoC6+BJTxXkBLOIUKW9qtf5gZT+LjjUvoCe+9PDu1KLa+m
QH+DAuUMg4DlOQKQWNTfDnY6ynAH6tRTwn384YMXPQHQjiilD29ShHf39qgV8cai
N/6oFtCdmMz8eJEqDN34yLVOtXXnkN/VSE/kV0MEAd1MsCpVN7MWjTkOPd4yq3Xp
O2DsGqIzyl4HuyAOEHT2P48SfMKmO5y9AbQKcfzWnsqy/YJWCRK5m9J873yXWg8Q
yQ9ssWWkXnbDh7hi0YoERaU3b6+1I1zO/FRKXShx8wAphi8XxlqlwQ8EUrlqmby0
1k2tF1/wQUDZrT5brIj1wwpqQnWQR7NtBa7wvqaBy4MDzS80sFMTNTx3cDSfjaL0
lVTfJz7BdpUqlRgxiCHgbYxKpOQ8Zf6Qbu6/8v/CetbuiiJlxww6yelmP1rFIr3g
55x5hLlchLeJGl0jvsbfjnaOj3/28jsyMHxzt64r5GhtcQVIhTzdXcrLrqQBiKSY
LQL5Q7YSSu+YE1w0+WXSdmKVTKvAokeeeUQ3WzqM4n6MAUxCf9pYXlSoNOHC0GJP
y35UiflWy1iCHOnfhhfrO0iPRvy0jUYIWnF18F5myJQoZ9cR9ZHbK730Hsoe3Vaf
y13cJPF5/0llm/KWq4YUbKjtfsXsP5ZNCwjhwA+7Xs5BftVoY0Sn6SD65bDmhwuK
kN+YjasUmSfSj1GzJmSQiQSanbfrP5/kMT7yYduf4CHwgbFLlCZJpSIPpJDuigF8
WZLaNSa+d/k24op8uo5R3yPrhRE45qKnAwFnee4Jm/YXQQpES2rozCA4xpYVXRqu
Q7kAtUvHwKNLtzGxmRCNHfpPCLnhoMUofHR/Uf2pkRXTl+KS+58tas+Wc8gXfc/e
cabURsJiH745dla+WF1plaF/qxNF5a5IiRKMLBdHil6a1hjh/EkEJF0RvYhUYl/t
L7ohrwyXxvSvSibO3PhHpevMQE5KISlOMxXBelDOjQHGtIu8KKk5YGvT222O8UcC
GRDa10LJPp5StAgk6maf+87BuuNLFXI6DSA92UVNKwMyWQwf3/Ks2h9+/W8uqIeP
aceQ1rExOIBOFiRtgK+nhYVuQCp9yoNRvFbl4hpT9o42TluOwQmwpvlna22U3OrJ
DADgdu8nMf/1yAHwDbrCrYCEtIFIEhSyIPEGOxSPobbul5bH/avnGvBnrCVMLsre
33rKY3KhjkobPqxoiIIf7i00zK2oY9tKwDq6TEL4PW72iIS3KPwNkcvpMCa+PKxw
2cfxg2JVTcOIkJj3bfasrQtSW9rPPb3ShM5BGAB5DRZ4vh95zBo51p3rxmQY9ivG
vXd+K799tdxyohhQ4ayG/BXHQ6yT+XCHCCEqLZoUmN8Dul9yIbc7qbUc+MVIBHoR
ynNN+2YnAlK4kO2g7cpkYMEFVERYmuugN29rmQc9ttpOErBtGMwF8nNKcohDxz2P
uOFk8VwewqlYwVI5or76B+00f2QBIJIkwaqpMousQjOxjtMFE6KQjHaiKmCZZd8y
wElNudb7TENFHsKzTJ9IBrWKYB+fubEIlCIbkSfjBPFVRe5QRtIdPahtrN9PDuqa
fjlaWp56dHS9yDu3BNc5aSTXjFF/XmEFX+Sbwq7z55oA4xBsUR8MDM+bQO5z4uVk
Gy/jqUWb42Yupj/hor9focOJtmAEe9iKMUp/8nchiR4DODeijuFUhh5GsOjcjHT2
pX5fh9eVB4BLi1q3L4qzZLL8I5vYcxATvwx6VHsLpLmjHwZApN78un2Lz8WZz1PR
nwwa1yaFBqhYvUtTHyB7NOhsv8S5UQ69ZSo8fdp9DDgSED7mL2imLuf4Ptf+nTh5
Y2ZFchhgb97yaE+eUDpW0GzaOrcl829tyKxb2bM2SSUg0WJNWuNs5LmrTlskub5C
lz3sp9We/yun1U07JWjWNjVvz6XhrUSwaGpQyu4ddZukk7euIilxh8SIMbf3MFhj
tOgJLo0ErbOUaHNGfoGwkOONat1rJByIwwn/Ub7Bx4kMWMPRDGc1YGfdi/bdrMha
mXsz6uApcdJh7Kl+Vn24ApD42dmmvc4v0dHrIAvZDsWKyDEM3DBlPf3GnwrveM4w
OHCawe8hZmX4ntTkvFUNaq5pgTxBXYotX3Qv/sAlhvCqkoKhDWzGIJVIi75mawQO
cDmmkIKLaRMC4oS6LYXV8FAKUaCeXIj4Eb+I6PsOqw1enyoFVEMtJOo4Wj3Ja2Jq
W3FVjRsin/hu1Z/57S0v8rnljxoZBkiE4Sp48RRhqKb/a5KfWn8R54HTqOJ2DvCU
IjNH/sSd/4evnyMT/AXqIePLbbUpG0EokxYyTlAdH6XkoDSC9GkMTJu5H/FGmh8+
UmpHBaiwQQBQABNOILBiSMnpExPg8x8D+E0pr5LV0NEhDIQalZ9mncnmMsBQStLR
pPDcxs4CQKgi5/8fXLagPS+hb4GVuQnResEAywOUCdWGCyP7Bsx2JjQ7nRJsUChm
EVePHhviANHJto+LXDRd5+XPzPlmEeUZ6QbLuhXHrdZQOR/Lj0lhP0uYg/R5XOWE
T0Q7qTNEB1WjTfil7eTk/lfJ6MKOh9wmHvK2wDXHEA6Tu8bFgTmvvMcW9bY/2BiU
AtKIbzpImT/Q803+e7L/xkbICNt57dklRSKCfrWE93DUhwubfpUbG7jSsr1VQ/rX
ZEj1sPKJkBMZkFRYtZc82x1ejT44sKJ1rD3ZlK2pIKaviglqJRkEAOtHm1aOPBPO
EqwoauLEqe9HRxscM91GBjuc0RheZx3JnkOIAYnxJ5qchuER0JSyqMD10j0xM08p
Gh75ZLyhrxULuJ4jZilZcRfrs9X7WpdlROSzLs1nypP2JPD3tnk8f3SW8u9tcklC
ThV2rdleeviFJc0Xa7LyCvpzqUVh+KDBWu0ilKNWxX4ACH4+vOtBWQESQSpARnqI
VfaEcHca9r/geF6az61CX9CrM82hfX9EpmAeBPlekzNOX8IGuZwihlgwPMZodJFe
BSSN7EsZo0iN979cSJUN487aBcdbOL2l3a4Yo8bWeJt2zNiUVWmE6zzd7baDOO+k
iRMHJ3PwJmh+eJom4Mi/cPdSvG59WQXaXhRkC5i++5+wncdiuoME9Ffmx6e9ebOr
yzxbQozzyBmBw2SxP5HD+Mt/pO+1s+/L9ovhe+xih8QKA+fKiyc9ZbS7bvY3ych3
6BNAo/pjWFv4p54YG8XtMno4Y6Sl3v8Jj/YM9+nOGLdqLT2Oilf5CuW+J+qT+JXD
oarvWmzTLjv/ji5heBKuGgk+zOXDocYmbZ/ZNM+bDZrmyFjRD6Ejst0GztvUf2Gy
no3fZsAj5WxAt77mTbf/rSqnyy5oAoCtFiY0doTS5w8W2nJb9rcm+Vr5MXvAug7D
0mkw83p56dzyFHk0xJviVatwmn8B/LF60CJABmdnxcFzHYxXoNtDKudndSukHd7R
2TqFcw7K4/J4QegocY1a/Q1JqEaQ6H42Y6pvcJ9uoq30jWfOuDc2tOIeI2PLOPBY
GJSH2Iv8zfNnc0HR+mBMFgIhllOG3lwUXfxGcGbmre2NpUcSDQ1e6WWoKq5wGMBt
FkzVRmy4eyKKK/YXmJQ3p7j7oYNRSCtYkviTMJgJXfaEIN6NI9nZRzN3FAb2oxL9
jvr1XNp+y/ilprzWglgRc2augDFS8D0FtJ3STmwaPNrUB48Y78KCxyFgE/lQEwB1
HIzFq2vU+D35isVhVGwO2g+qgkuavjKcubawu3LsegnOnz7sh+d9VGlymhBpX3PE
uphla76gP4ZfmT6MwLK3l32/t/nhtSFSkb9S8HQ9BK/5NLNoSoQ0arR/n8KwezTZ
bsDXV5W4b9wTX7U6UtiIFjV2UHL43OGMTrXiicxzoJ5mzzr/M+MRNWBqN9Dvy9xW
+c/3f9t6xgKeJ+urZhuccUwJ93RecV6VCxRc1LQJBfG1d21O+38gJXIZZj8qK2RW
I8Mmah85TZcoy/C5noSyC4NoOxmsI7n7xjjMOySDHnFS2lmiwQv/VD97/P8YSt3R
HWj7SxnusPXatIM62lBA6dKZICk7+mTVv6va2ucH1sTFrwIE5jqlXsMvD2vZLf/G
n3Fj/ZDu8fWPQrgbDRGIqsccas21P68mBydpEfSWgZDynkoyiRpKtxxItMvBnwE3
SXgSYDqejy1xX+IN8z4F3qnrzo/5lZPPmH0zJgZKvUi1UjYayrzfoBeQrHwJ6UQV
uNeqLcpByZiDenVPMoXh+HrFVB3jWHrZ247Imqp0tUMyDdpmhYRM2MEzE5gcLuGo
avfGOHc16/C2t0yB8DgFETPlAYp+2G5WUTJGmVMbHgk+XQHDN63qBT7Hh1+zx1Ks
AvubD9ZZE9WXlzIKGwTqBL6gKY50y/IOA9BsK4AWx1xsWqGZ5xK8QBBVg0JQx4p6
49icS7F7XUkQxBZQJt0JNj2YZO4sMR9w85JA1RhmQCIEnruDlDqsfiUGLLk7H91s
Vlzb5hqYyqs5U0xDOWvOeblyQGKyFul8ZwhhzyOtgjRI2Sjd+IYNgdNcfG3ncS7b
GRUjkERBzzlDtDDTCBEP9TbvrjPhousTebnem6Cxg1IAmvYqFqmWh8LjMg0jGKwm
3Q3rutzcP4sGpDFe+o1+fNu6Ycx9AmWmiOLkKx/vowfhL7BZuQRQiNxjmaifqq6v
N1h3Ux/xmsMdWlShdg5unyFJAKl3z+RnFa2v29/Rm0MOI2wzpRkrp93kqj2uq46p
NHedRilkDmvR6gL3XBcyaOl5GSncWFHatdUL9X1BXVWO+Czo0Q4bbOv3EnQ4mAqe
GpDagD2l2seP6Ewl15sED5uwtVWBa9XkKEfnI226EZ3H4fTxIYHlyjz+FIkEYwv6
kG43kRKkbCVIBX2YpYs1ZbnEiFee4ZLUwd8TYoxMroILOMDjiIRxm51qImat1ylJ
p37Qla4f+eHqSk1O93a9XzYO2nt4FTe2BXpmas60BRhRuLnTWHAlc9op+4ShCsnA
Dcgo3cRQ7IYP107uWZU62WNtWadS3WrPgzxI9XebfbcfFPSaiB94mJgag1J+YyY7
QZE4/jP4/KYQlz7cH/nyHgh3AfnnL9WvknWTphK6Uo/urwKi80OV0hEgOtPfKf9m
OGAADAO4cB3lP6Uo88SxIW3TX5tq14JX/wTmYTrrFXjtmKnFiv+VLjfZvGbdTYu+
SJAVOYQxBB+ZxdHNUiIEwfXoDdJSc9kwLaiNkoIXbQssfXO5xe6F/ZlJT01tUDpD
bxSKlO5YRZJPeMTnHmXYMyAKzEVIpoR0QKQtfdQMEOQzE8XPmrT+5fsff71qs3Rc
mpVJWcvsT1m37P/jKNGWuDfTdUXgEpTWjmXCygQHSgIxkGt3eX/o3tiNzgp/Bt5f
InqS3tM4utof2+uiaYrxk2YrbzqYp8Xer/Wmc0KtZIz30chLuwnulTlnOTFcTMYg
7usgkEG4pnINbykOl8aTTKT1NSH5qFiUd3Xis7POifsUFN8K92DqOohU9l5fU+EF
U72ccqHI+YEB0bUBJp2z3dEYY7fC/8x8Fl/k9GYwS+0ZC2nyEJhNOcXGngEo1UiL
`pragma protect end_protected
