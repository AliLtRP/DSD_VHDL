// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
FxDHrP0oS8IOdCa8LIN2EQwshcFLePwEMUpfAmj9nOxW1KbC6k2x15Sh7WNp+ItxgEj+ZdkHQDIb
hu0cKl4HDT4wLa0Y83QRvWE6Mfeo+jSDk738kWp7ij38CpAUyxvbUBaT6JUQMYM8S+tD7LhM+E9S
49M3Mz5mKaazElh4OOHFKGcwNQNQ/1NZHiiEF37SPbU/jbYR9wnONYGfquY6HJdeD3AXt8GFI4GV
OPWJnZV6QXeDLRfWLxT3AizJb/PstxBKmHo5/jbwrDU02B3U0qhe9ACP8MwAllkkkDT0z/qmHJOH
vW2ZIAZM5e925fYep/yX+XmJ0MVIwcoMjTdbNg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
mTsZTeLBgVCaV1z0TvWYtiTwyqJS9K2dansjnN2jgx+xIAKV+C3o4bQ6RPByb1OTeN60oC7GkE8Y
WcWU2UnGNoqAwK7EAKWEw5AvNBL3bBzQBoQqlnLZZLeOlJCWHoTLz2AZEHdsetxXizTm0fb+BYzT
EqNG8noi2R+J57CJpL3FTbeGQDbs7LbmgXfYIigx6kXfG0Abg0KGWOvyM0xoobAb4an2zdTEV+1L
xw0PM+C4T0r8A0S8dhbyIr3402BzGMYmr74dDH1zGZrWqGU2UUvRFIaR5NNYfFXODc7Y+fTBZkdW
g1bsGQS7McqCkPbczE2jwrmo/cbqN7n6bBSRRnyHJ56UxFOLr+/9QFdiznKtnoFZHz/7VrkC3tiv
Al2xHzh1IwURncTOEF7lnJR6dQM1uT89pyuQQzVpQ13ARk5sWuFAez8nplMWwv3X77l+e3z+mwm3
g7fVANHdE+GlI/NCvT36c6nEl9+lAUS9S3tBzYhZRibYHiFux88QgJ7o/KumUcf0jenhVFPi6UKR
pY+u6Pl47N1QqtPxKNOeBhDleAep8Wnl7TBn7Hop3ik3LEBzj8xva7UEaEf/KT7ZYbvTcn0Caszw
E4fA8Z76p4dgkDL5W3C+A3LLW2r5Zp23DEYRSlL+x6BkY67XrLi8oZEmHmaMOvX5VhaYBj+34/0K
5d/SrNLJ1FeDN0QYB2AWwb8JIe0KgTvqMag0BteuIdbXY/ICblpP8vozgfVE7PJiyzzUmJb7XXUp
hq6ooAYiAoCXrKzhHQ4jEwQvbreLTx0CsrLzzDQkD9dTxJsfdgjbCJVEv7qGt16UuYaYm93k/VG+
0NzuTC7MbJBfrYjFo4TFs7zeDlY5NdNSf0ibqi9EoLd66hd/fBsO8Fl+/ZvAIkFZtH5UDlPC4X1k
3B83mJ4qJhZC0qWI3Qcoqnwt87Nbw9FZE64vuIBqkVitKebt5M0X3x+XJdb+HXYGmxFlQHaslCma
JS0tQ9GMLJn9d0H6Q8A8kMasBxW2jlTAdEgZUBySd90r56F9rO1bSVMRMGvvJ64Gpd8zlyumbC3u
aEN6UdOCSpZLAFGRbPFTm0GT2jtKBANxma3UKPNSSH9p21PfgBi/evM28j7U69uLhaH0PM2zgj/l
d/4KTttr+h4l46SKLa5RBu5oHX+s5fCeaeS2OmgDSkynJh+97EeYemfXHHVMs3aOJ2abrwwVVu2o
ba398QAIa6a0rxzcLTKWBYquvIIbozJVFXaa4ckX88FKbcohm7QlbUPoPqaFcyRrzFYKPdnD9glv
QLykOkBBvDWHmCXANma8l9/Pxt7epx8YR7i4s3iOdokdaf5wBH310Ztd+vsia2Bk/Bv1eDe6iZL9
AeWeqGTS0iPYw9i+swtxviBSKmFv6Vb5GKsQILQyvbBHvEXSbihVic6C+AeJ3tLmYqkm7qZ9CIBx
empNA8DvIWnThm1Ri3kIYKFzexnpf4uMFM/uWo8s9Grc4u2hLCzSKVLmyf4yVEtVNc00OZGpWX51
NhRCzPg9of2acDZtqYxQIjUT0xz77aV57TBVyatzkeRionnPeyDYRhjnB/LGG4LaF060+Vhu57sD
X6c2Orp/zTuZpR1SyLjFsQYeP9tvap23IP7pysghtCQ8VkXYQyrX+UsHejSgj7UpJHD1e96/5Qm9
HxDURsuVhD+XOdHSQOdZhU3FKQDngRKWsCmOQq3CxEmxtQY8JWhLK2TzlyVcsHcg5KVBz/Jwygl9
IXM+1ci+EoGhU2WnhFrj/bg/6aPmGGLhnRHESNUNugbRltqZL17CWmEyUps1CqbXhtMB2yN1QnRd
ArbrglJr0M03S3BQa6IZdT36DjvUXGqj1BPh0FvKkDJNEZZIwZMw63pCBx2YDJLR9H0yP7maahD/
xxHzJZRy69qblD6Hw/DFvUpkyOLuy/Ev6vs+O/UgWq7MTEsuwNu4PZJ3IBWxIMUEwRA9/32SagGW
oAvSg2yUl0d0mIIMnK0c8Kud6DmSla4VSACUPdL+YPUMa5ByZhUjAuS59Ipq1jwjIpqd7dTzGeqx
ZJWpVKdKagxkF7xHd+RJBbkg9PiLVAyQiMIbYVb0yIwItQN0n2KtF9wH2ff8Aa0pWykZlwnZCFqD
ALLB9Ui43QS+s+U/2OqnbXPifcDGC8nkMh+cbCseJjUSyCIOLzAUIqnqTdbPawtaCJ5Z/hEC1jZk
CWcchav7mKbMddV7Df1j38w/OT9Ad2v10+505j7+1fgRE8wCTSsVdQc+diQLQVbadDSyBmeB5ehi
umqAsH0DEsZCFLN1TSWzKHmTBr6mXeH60YU1QbN9NGMmQfk3WfbGs5WSwf6KV81Rl+DW780hNJmj
Y9p0/cGdfC1uX7TroxnELvgRrPIM9US+PqGo/xZQXeTfzdgnBEMfOoParJJAeodAYrAr+yNworXo
mcYrymdYga3bfXDxjRiplctYoPsqNMLOP5p6SitVFBwKpuG596PZJe+hhzC1h3k35fHDbKNs8+JN
FiFggeoWuNQqqYkfQI4CZToZfZLUpuD3mNK7k6Mdsw0kT69uRWeNC0MNsZ59NG71CPlxINWAUNZq
gT106fJ56rUAew00v9aH8IxPB/nJP+V85W2G7DXta1JrNgwzPtxy0UAa6VxhpmEXQjU1JFLBsUQB
z8LlpTBQLw3YbRrZVJw4e1+KEt4jPjC5ueeey7djKkR0ScX7HMMMJMTKwvfDI22jlUu946JHz5wh
j2fAqxVaaBo/3hp7dK6P6XKYu4wacvxsSuglEPc3Q56+k+6RrVLg32NseTj5V615RVNj4i15tZ7T
+Ls4GPT8Odux169wj0EfDQZUUuwOr0odApad9+UCqam75wO8FVxclr4elRxYYYLP7/MqNqI58TO0
JUNc3Lo6n04TA1YMyvcl15VYdMWatEZozru85VtWtmI+lk7Pb5sBjvE7MYb7mSJfl7vA4MBwpExO
UvK0JyZK4xnhL28IZs0lqlmfuXhe/FeLlAQ9z59ey0y8FrXFzYBdlyFtPq9lM4xbUjFBJBGWCV7z
V4NCB80rBw5ooqI3xOwxQ3Jegz4skzqv3CqeGNtEsYWujw2kfgOKCO+xNOO4eTwIBm68VAjoL9d/
7isUz9WDibYf7kBwFN4I9SH2qskm1UQUpVC6yE30OFhZXgdqZX8oK5v4F4f/Jaz13y9F3A0apL7M
jSIaz1hIO5NxizjgzZmgLTSsUrAjFrF6xSuH0rRurAGdPiHfNxpe5TrQZH3bYuxL9zE4R20ThcFS
MnED7hVqEhfzBr/Eh+tSPF8eSnaJcWmeBMc1H4P3LwFjGl6oDIL8pdIaU8MHvdiu/tb04ScMnhtB
klASr3UK0rlaz0Pu3uiUZaHjFhKGWBjhes5F9W6YUFaN8USr/z/AjT33AcveBrz1h8ipV6HrW9vI
Zo1xAOqls20kH8oKWCw50SRahAYmk+aUVtwgxSuYxUffuLKS2uoOuS91b5bwF1313rXB1Cge9Iuf
YzLadBgsAjzV3AIz9BjoqvjU3YxEv/+LmJGAy+HdV+z2/UzpFC7rzXzcKd4xV7NU9eZL1lcmKVXa
7T2x8LnZThKBKYOBLBJyD5YTtJnqroTvTCpIfxINxo1ud+82PmbsWAD1uKm/ENxCaMw5Oqz7CZnA
vOpCsNQqj4lNEntdT4uKi7C0AZrmRUh+vB8vS45upt/TTtN0XMPoCcnGwOH3WlkDO+CHXq8PPRec
L5+O0K+ihFtMV5S0R0bWyvQ6OJ7udIgpPacRhY9pDo8gqx9rkA+8j/9wicT11UDf1O16T63p2Pdc
cdphpXC5f8tZ8grofcql23x3GrRvOvyBw9rVKOZey6plbpnQuuOtfFE6NDEEn2AnUy1KH5ZcVe+G
PJu/6qjgDhjfbYbLTWe83rjJ6dtN3TwVn67zUH0PkxoHw33wNIoiasipN7r5QlL1ZL8YSz65lTLj
c0nQphd4bQ9pTQbvRE+B4BfrEC3LPmBjFwwQQ63SsAsACnUwrADYYBc7vFtEW/nXPm32ttMdbQO4
mEThJjalYXk1rnEvL/K1dxb0oyW8Aa2/oqMK+rIa3Nnm1y2F6PJiG39pUJksvCcYTwM9s6IGaqay
mp6YPP3y9oeHm8WJ7Vq8T14lYzEe8imZhvpsFPJOVQu+j42J6Xdsyy3vM1WwinV8/J4sjvv4/2jm
6fd4h9DGPe6SeL3odUYlWHwzvdYQEXQm42sBo9Mk+fAF044oyUnBY0tDY+nSVKvlJ8FakR1Obr/k
Vh1sQXxyosKKxcFk56q6qbDA1T06/DicNfcyB1URnUp8dK5iZMaQQlSI3kddnUxwwqF93Upu3DHX
f2sLhMDHe2bV1FSAZ5NjpgC0nce6ukltGPyTtUySIaSRgjGK60lHh5vgtwYSezqd/5gCFQeqbu/l
v9nxe93ZWdng4x43DD4I68nyYZpSi4a4S6czohxfJzQVPQ68cmgPuZu9NIxk+6xa/ZAGURLgR0ah
A2RvEPCpNK46nN4Kueow4WZ8WKhrs+YqiUkfAJxNvpa0wqFX826vDCquz4QenNJv2QHJt6UfHmJi
ed5/oW1722DfL+f4OJKQUI3Ui6ImTOZ2iRxhdVUNqhNiM7CbsYnSLhg84diubDMN7VYVp8NhDZEG
0j+Uq1QMEVeso62l2RFV9R4/QRHtJv2m44DVaMfO4b9yelWcrljwb4JsLMv0CkV6Cw2vWKkqFj8k
bzC+kpfXu6R7cWC+RaXWtWlv0YMf4eThS3FGTv3DRVKhvkcHYiTbrtVO0omkGw/xcHb6/aik95T9
y4bbatjKyyvbbNy0RDj+2Cq4i1y+4bv6xBD7b07pifWwKqtcBJeFFSfLP39d2/hi9VVXwbEdAmsh
1V4HOLTMZS4dl2DzucW1SBPuOGZVtPMjOJAL5zD/bHQ/4GhMoUCXPUCMdyiV8b+sTvkNVieerEau
e3sczctbsHQlmv5NU6tvVF6l332nBsifXi2c70g1OUtK8qIaHP1yOIFPA9ZBEyy7IagohbwTJkKZ
oZ/IJz4J746nONCGq0sUZifK3BUnruYWhdaU8Aheyk21EZQfV+tLRCg6X5RoMNNRzwoYjOEVCv46
FYQ0HYAouG2QMiTyIAexewqsuQBtQI/zssdhPQ6cqO5ztjeh+b4bfY41rzB7OZl7VxyOamTcv4q6
8PxOQGc/4oy4HUPT/tgNxrTkpfL3HGMXj7E/WYVFtwVOgytAgJw21fzXpqfbE8lmy5NQAGn4TBNe
QFI4Jpt78BGO6/MhzvlFxQ3/nnfLuBIdGxohfd0wEhUY6BqZ/aGdOtA7FRAAxnQ0FsD+TPBAP81l
Zl1nzm5LodNzWt82DvdEaWFO8eO93yOO+A7iJgNjPxzQPgwqnnhxBrRvyKZhbW3oLT+DZMR3leof
TqvyhS/cGddlcZfUMqUBonx96nAbWua4bQBhDRQ2lGA8EtG1W2G6Agth3XO4mdBXcB3sM0h9mKuO
dKHOdj5v3ZcUDypzvIYvB+L0q9/KPSRt4vHhcH0b4CCxR2cQQh7i1ASkvoWHR1Bh/Jz9U+WsqX8T
ehXCPqzVClFD+I0HW8ZLXbnASzlOepznFbFGTlmUYCGuWWrgLnLwQ7QZpNf/MMTefV8k5sLNKtcR
070FTSE96HHLQjhEYLl+hDdxh/DMe8r6992L5uuJnghtY74T9M3tcfj0twV0vcemeBb3ABuAURqK
uC6ke25FHfobkHuDQJluMsXgLgilqLVTHP8HlUHWxtu//jTffp9a8/nRSWJM9LUN5pF5p2pnE4jp
WhpCaX9OPLl4IWXgPnx9ye93JWNLqHlKreDz0Ppxgm9W51N5VYJoQi2z2jLjjHI6zvmTgJvaAEYe
iOcZ3Oqpzjc54D6GXhqSB80FMD4NbpRnWafr+byQXzeHo7R+0c1IOVK01aQDOfJ4O7DtoSQrHBUZ
zbdGjZ3N0DeYHHfSYnkk7tcQAS9YzVEUpdNVVZ5WOQlKGAzurQD/4LU0Z37QBrPT2zAUbkUJn0/V
KQd1xACVXzBPKggrPFMFPUzLyFRmqFn/zPu8nfRJZCW4RQ7ot7kfMLxBzk7dfjZii1HrFaOXXNeV
2sYM8QokSqgfNm0g6OSyYDc8pSUqRNb6LH0ZHM/xz1l3RkS2SVP6FRrTpKXqHpJVmWInfI6NwipI
IWOQBEQXpd3w6q+5XdJAbm6i5Vy7BVtEg3JSuE2G99El6mdRVGkzk39W5dPvnxkn9dqC4SgvdjlG
ORPzRs2HvJ9n1ajy//zi+sVaDMZHAqSOkD0Nf/RQsfmq0XoLgDHZtArWKaq1wI3ZzMG6hQSeTsR0
oYaeM3Gcb8jM7cklNNbs2PccqXNw7o88cPFvsgCBLOhBS0khdyQv6l1r3p8NLr4UTlP9MT305E8+
QR6gOnI9EVPs53Zjb1vQ8ZRUvEonC66TAbOYzjMFQJ9eqt/mIIDHPj5PExBCryPMe5Tie+KFvaag
9PFacZBKMqjlU/mvqoRdalIcUuauGLQzfpBBCOqvW2FsyHuE3SJrha4DZaTMiS17/pbbFugOHnhK
ebHh2q4ZQgJ3SW1alADvMoIc7TfJnlpb1I5YF+7LH8M7ESluDzO0rO69PjHyLv5/j7CWCf65A+e8
SNm7npZ4rGuSAPJmDubf8jquaFChhN0dzYjVZvR5HmgFh2Zvcb83Xe8E/XfOurgNI5182SoU+q7c
2iUX3WUGCUZHn04g3IyybaC9xepUH6GodnASggxQvrMshQ/27/asxrIfE8yZnAndOXQFor0+AKu/
wBXvirsIZPvv+l/0K6ahDZWzB/vN4AE/OeUxKI9U4i2zI3s8MKJX6hZ7rnpadrSYl8WfCVmKF4oT
CrMA5bIIke69hkxazYG3yMTKbSysWgR0OI6G9w1L1DXSZkMSayRMGRpj5nzwt16aeKMduKM6ZtOm
ccEnXMgQ6Y3I2r1b2eSKujdwX4wQ8UzFY0xJPHKNm3gG++VhL51qVMs9mJO3wmt8Hl7smoIFyekB
/X+gkDlNGwRBCK4HIGG8Kr3jQu9h3nRJgGdpu5Wfe4puTi5MMZBfOF/kTr/Pl+ZhHWW93vCnp11x
UbL3/l9nzOQHSozi1wD32ghm/AGoeJP8kYNkAAsANw8D1qtUDeWcRav1taK0G87WhyBQI2QxfE52
QvCcwGWf5nnRE9Kycnfz14M2RjEMffttN8FHitqJy3oN4HPogUajDGGrIKo02AuoOCkYMQ0BCh3t
h3GMyvNk8e7HWSsKShuE+NVVAxuDXD8Is0e8cfKTlon7S7hoTkA8urgi8LF3w39ELC01lM8raPnH
2caggWEQQaZnWjnmXI7DCGRw6jcjzBGJryaTdgvXB/1ldH/P5+EbM3uJ8kKGQAkr0TJmR8ABlc+V
RAgzrmntIG/CSIQd70kHb15Rktep0RyNF41JUVvCtg0bin+QYjwz7eKpaV7fJaIfDykz46nERExf
ISywaRCy3U/oy7h2JJC6k2WIsW9FNne6NhikWwTvCFPnIKVKpr6d8sgnQq1UtVF0GwRnLRWLst/F
mMAVQd0p8WSlLYQomCDPSh56XDhJFdiaBfFTwojZ2Qn50VbI4cnYGphWttanONNpAv5SGJnol1Uz
wK0OoBggybOG62FdTo9DuqGpQpsnjDOnCMpQjZ7qKes/67bWE5nBba3FI9mlvKTL+eUTl11I8syO
egF4rJ89ln+jg7kNHVT/PsJES85i4Crp6059ELGLEEMozKOuqCWQtxXa+gYG+IfNXa6Se5rIKMJ1
SSSuzd6Q2FllnF+iX9kqLRjVPH0GyBdoM0rrUavk3LYWbg11n5N03c/nz0VJOjU6CGFwG4Kkj3Tg
NlZCQ7LsCccHbO0WsorprgTvl9eItKbMg7s5cNGtP/AY2m6pHuFBy1kemRrR2i9ndJ2TWSqHmNzI
TJ+V/1MLDR9bUGLhoMzDUgJYsFMhpaNOScw2fvtptJWil8kvNhc/fnnj2JQnawBtL/yZToMYFb15
yAYwCWoNvMExGxg0dcG/q/PqJY6QBfBtvBJBulVkfSThEWmYynEfAECm05XFkwHCN/cGtbWbLsAr
dZ08e4kcqA3jCGUQ8Y5cRE+b52nO6IgpnzgllHEM4qGOkgl7q9MnAqfVn+wKOI4ENWZ7JwSY+gIq
TF3XjmT5krromWz8IEX2l0f/aUAJHKqHqk+LOaBekdvwf0Q5XIOYWuqB957A/w2uJguYGsft8d7W
kMJ/RQpYPiZJZhzr7p9fCQJrvuZCIPEAD2IOaV/vIW8FU7+kUQhomFJKcfqbTlGQP4vJtZt5h7g4
uEw3H/ZNzd3K6JXlSOb7KOfWf0Z87BsJxiGoFjXHw3m8khX5VGAEUOnagxuDJVMpQ3hO7zSCiIeZ
qI6s3yHj7kb6y8+Hi2QUtnd5nmcl6Ijzm/5L8cV9CGHcPhUI6qIN58eqenxW7h+kfNZsV1aK7iGF
yrLFsBD7t/INJChoqp0BR/fOYiEyqzhNVNobIgwlYESDvLVoO5nMoqYi7dbDIEITHt02HEb4UWYQ
1kjHgD1dDU9EXeyNpVedHrt5+1YRkCteHwH0wEKj2GWZCuvCRw8G8ToUBbhedd1H5BOcNZlQ7gZd
hOif0EsmZ+M8kRUfknZvZCNvCRdPeodMfllXsCjJ9MG+LfB/szJdK5bAoFTvl+79Cp+4Q+X5lM/y
G3g9eM7afQh47Oa7QW8sZkVKw/taONZ1yf0AtNQdqSHlxZP5zS408OD8fa4bJmwD4FjqgVms9TDX
caHvaVKApzKx1hiPeGVxMvuP/zoWcXA8mC2u6ba/KpAq7xQDQK3xhvbUjpWEglHIprHcGRLSKWvz
KJVfzPdPHVe0IYcVr+G5a22dtmsao4HJ6bfeKJ+W/CbZG5aAxW5RHTRTOWSg98SZfPnd3NAOg2Ag
nmgFuY3aNsN2bjD3FnAOe0ebIKBeIIIJv9TfVI6MhPjtzh6ffPxhNAGXnYTrb1gkYNidj2E5JcE2
2QmtB3BSPHL9ukbV3V+wVfVv0Cq7VrSC/JBCf+LFsFqn/8LQhmVwDKoZq+wP+w8j9gLukHFWZh3y
EjR7fMe377nJF68ZgZJmgMSB1z2HcqGoFDZhTkkA70y9/zAPZ/lu9aLQXF4ytcIqGr2oVTW8OnLn
hzagx5geat+esLM8eJeWUCMxRwVYb1XOV0Y6psOunUYMMFZsc9w2I293tJeJ2MlayrLgpnq/mPtR
9A9Zs197nAXObq5FFUUfGAZtpZTrymzTTU8iihSYqkLk/lIy/5AXNP2UvPhEHcu+INtnaOEHbw2R
pybFOSRt9SZ9C8Mi459VL1yQuXAugILChun6Pg/U6VMSTBKG61rGdoA4X+DxdTwCVKZgAozbebGa
J/K7kogr0WqTr4zqWpuFkN1BwXo2ZwTpiQf+n81dz/t9ckyqCO3NlFPRtDufPC1UXHq6Rd4zKgMS
S5k++zx7NtA0cDkbFKY9zonVK1q/pWdJGhLmzJmSjH4hGwRHB0hmK3jlnhkjEXJjXV715QNVviXs
KcoQvQPlnppQr7ixfu/cWO5uREXmP68DGuAg3JL4M2WC5htzJAY86hClDWedgNgCJfJpSQO2kpw4
o1DR/P5YsB/5c044OBV7yduSVnl0FRD6ra4SLI+dSUX9AEmj2npxNSF8fV/Vd7C2kSL56X1FuZe/
bBumw4GhDK75C0RuYZQo61n1/lbz1KBb7AwIZhCCON1MF+B3RcEsIx7+2TkRLQDB9nY6hWSQ7RLz
m1Whp4KwM7PZciq2xtJZUXEbN1spqVL3uquj1lnIJUy7Hvl0dvg3AcP81UluHMt9mOb3CCSjovJb
rBN7tJRlhLJnSqq+tkRUGZMnT//sbjc8Nqv8CjZshamVcP4YQ/1CLtpeTHZjnukc/dtqDvtm0XlJ
/d/fh9NdQeR9+8omk78XJrr5AS6W8MCpMyZWTgrzfzIrcUMxwAsVQgLZlnGMT3a7hnoGm4yTUW2B
kHvHvv7FkCwVRoIj40uhOfRDZKWWV7Z+gPO/q4sZ5vzFIKBaE7Wc/lef9Gs/Uy81n/6G82Z3e8G2
j0ySEWnUDX8XrPkaikY4RXF//nMzn95fonA+coZSJLl2A8jxV2I6NHR719tGBla1/M4ZoVQN6TM8
edBzTESoS7e99On2Yxp2PX8WYdhDq1bfdB5mz9lv3bJtMdcGy2ccZzaIxM+plHuZ5leXFLxUr+Eu
UyKgGVwLR85ERjN1lAuPMzrCRgSLnKL354skX2KvP1uvL5rC0RjKaZ8Vm6tdEWOFvWEZ2Syw9hKn
P9kM1US7jmwSxwQw3+vq/LV5q0Nwu/ryJupKNPKQWoa4bWXFWMd/mCsZNPnVq6A94MX03c2uY0ji
VK9fhJjLEb3AamsPHwkePhdRZQKj0kUAnq/fZjdoQjxSkZgnQdk9yjiQtkiqIv39Gwd3CyIMaDq7
2ebYq/RSMhU4G7aZaPhCQLRnCVc3Hw/2tpLswrBHNXgz1QKoqPU2ox+CEFY8hAQ4mskxN1wLwIZo
GjFIY8FhiNZ2r588tdMLksAeMoqjtZvsAUlCjD8u2wCy7JC87EudJmBvNJCPHAeocuzxap7BjHaL
KcBJC23j6W9QTnUIwpD9z6yfuHeQS2SWf+MxZpq8no7BNhskYTfBEFrbCpPKNKF+TzjHObauliaw
aLY/zsS7iilk2qV555E8TOQKF64pynNbA4d1NEge7c4L8c1yXQfPIhWy0ANSbSKBK2R57U06mEsC
jGKt3K0P3+cM1H5AuL8hMXE1GYSJgJN5Tc7eR3fB10izNXuepnBT8f9MxCp/xVzx9aKH2eli5RL1
Qr3IKL8x5bUttdUYvCkJIFNUmNvqiV5UTV+g4kp7tRmsi2RHlt8QMWqDqVq810AD+/uJUaTNWL7Q
IIrvsLiur1q+qXslbZ47rfQBQ1MGKw86jGd8f1b/jJAY6TkAiG97kAG+hvU+QgQrPeMAQT5d9X/Q
OUqccibRMXZ1q7+91G53DsgK4RoaFerETIcx2QEMFKlR/Nr97Wcd3Ql9nOcv4uhRDyfguSSCsqtT
jUVAmS9AnGEqPq9N+7vQ9OamPEIl3yO2147dtfqEuL3yHt5sf1oYaZacBbsnxeX2sdqRx66Jo0I7
MeOuiOhrQ448oZwBgtEbDb2JLq1L1o/UQ4dEa2X9CONVkENJxss36kagiCQZ2HCfFn0hwTdX1p2w
oVw4GeM+FKvafFFO2hfmk9f6a7b1npRbAfNLq3DICF5tXf6PctNwBy4ACnKAWSCXyFNDqa6O3bQq
AKetkx7ipJnHo+wPwrSCUG5flD2f9nSnGQ3AYfkz+oDnZwZ+3Yv6pGZroI2Sm3MHcfRZ2Exk+vGZ
iN3D4PUcCJ5EQRL0mf3DbmVGpBCiDOkzQBwsGNiyOkc1Huv0wU6MZrpsfs26BO6OiTeYA47s4Cin
f+5gBaoWChpQCoIpJf3TafYwsyOCLxAf+xmIT2YtzrMW91FnyDC/LlYuA+jnKN08iwcLga4kNFwX
UwgFSEK5b2KnEfg0il7PFDqRkB4CD32Csz9V1xVwJolbGtTIIBxnn5v3O4GsplUp3EQQAC3h0/Vz
4JDSZJyUGJ4SUVZhUEthgiANy5vDT5OypqbyjTkG+QYcoXcag+D0okTDiv5morF7K/CkSMaNJbS7
0soB9U6aCd0o0o6Goi/YEqps6gyyVimjB/yDGqdigEQzMo3rT79iEAAK8YC2tr43geSNdWOHO0tA
dE2MuLEebb1Abj6qX1mSULH3OnrdNSWAX2rWdYMbZRMhuQxlxfPyg+Md7/ov8j4ZH0vCAyIRhx2B
MaWI9kP8RIlTer3iuiCdWupd03WXCtbIA6WmfvhV0jAI4akb5NEcx74/yMtAk6Lpbi3mLP5/ib61
4HUZll2vQzvQLxedUytuumw5l7f+NFc32BesYNRjhkQgEFn936SlE4XtxPijx3OBMRVn/VVTWwSh
47iXvK6gDqzoJAZoTxDTovkILe1Z5hPV9YbMrBS+nf7+c0iHh6E0VDY3Z3ByErYRPk0bPZTWS0YW
Um2TYCqzO0bLNBTU082UL2SxcTzQEdqzspoUJRk51LsX/IfFNa3r19K0AePNnW0ldbQ=
`pragma protect end_protected
