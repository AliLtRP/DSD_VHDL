// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rwytvv1XIrboGvEMCKwPJfIQp6b6Oqlf3cDqp/DStM1v+6/MWscQYd1BpA+r1CnS
SydrdfHJBMzpySUPs2O5hf69Sw9LCwpD8yGdixfA49nWP20fY///ai5GiR8n8bYh
PFwirUBmYYepq9pVHlJLHABLX85o8aoVYS6ncG4tidA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23248)
R6+5/AW4JlEQ1i9dbbP4xw1UAaX7e4RABgmhH0KNrte0EOKJdrw+2/nYlauT1IPm
c04vTMd8jC1luJ6dnbtM6WAgJtIGiByY42u0id1kPM9dHUQr6n30e73pt76Nde9R
4HLKo0iKZGWVQbs/PMDCEHObBsWpVRzTZ0a2ws6JdVcP9nxmUSJkEz11U697NvGz
NVrehQIr0deRAHmAPIiFIuy2xrH7TGKMP6WPrkPZf7EHdkgqdfXRMuaoFjyhtyxP
TAoONi8Li39Nk+b8SPht7jAsOfeiUhy1J8MGjfOHCAtrFJfr3Y+Dlh6xQmPsZqnF
rsUVR/1vgAGCfRB2c+0xO1VBl9Jr4ri5iwp/E4L5f5nPjFJxfMIdhClzMMfzNfUW
sOyCgi2y3gHQBxS1oK5AZnU2f5a88/2j3mMXDdPuKWvdbRGbL52ByEy+6itFoCQn
Rhr4JF16VW3/UHZRZ8jGMKKmheDjcQ4ZcrIPp2rLnsWGI6ndjUTObqA+7DpikNcO
yvDj912VAJXf7S8Qd8gmAbTQzMp53u/sCFEXpJQJI4dH5mZA/bD2Fe0WCdfI/Gih
jmuvbB3M+uaCEriyqHH6FsFM2ZjdjVrelATE/UhZMX+VqIXygUqiDowfNLD3vKsv
Icac2el09rRxSVRaJ8XZ6nU+44fVIWOgfUh947e7FDohCx3Dh+gEI5kBYXGsF+Ga
OVMZ0htzVMPz9MGVSX9vHV76ohwNEZROkCcSwQ+WYLTkmYG/49Y2xqIA4mPfncL5
xjU7XFwIAO5RgiMYV3PZ6+M57QwqUCRVA+BGvx2KuX1LF4YPX72+5LCq4XUE4kgS
e/lJpsc0KS71igzAu74a/2H27is9cyHm/axOGHct9TZdJhxA+kt89/H4G/4XSv2u
Vfxn6TfaDzq4KwzSROhUyh8pMN2i797yrvB3Bn4xYjUm4v9AvPMwBcN25DcsmQjs
a06U5ZPKNL2AK+yF6sBNOaBGBcQ3dLd0BNphGKQ6NtENI76iba5u0ugAh91sV8dc
trFKQGv/vV1nYm5mhgp4vmMXu7SYmuadLnMvIn8J4AUf+3SIDWLef/x9/lloX6/V
R7zwaHNrnLuyJoujhjX/tuJ0djdC1jJoQ0ZMpaLZaMdaRkAjiX03cAW+K9NjNA+y
lDXwjBTqh4ZKJqqExDQumfC9rtw6VR24J4mWUUG8vQ2lIEMBZxU4nEOqs4lPYZy7
7vecu8Q7yQbQ6KR0QloXnr7rQyuTSv+R7eC7qFIP3okSvE6MUkbvSqWClZbZn7QH
Ncmf0KG6JJ9mrZhTE45Ivfmh1u75hsH2ZZ0TWozSCj+uMsyCPlTNpUp3YKxRro2x
RyvgmS1EYLAWAYzaJbnXcKj+ljvC2qfAUtERXk1tsIhwAGgS69rkCSl8FU6dxbBh
sNy3O/UX5pd85OTlzk9IpuWtcoxnEWaaPGVROVCFJwc53JUpCVGZc2gtiEXvpuc7
M7zazUKBX88yxkyAW35H+rXHOiKPWxGcxX4t8iETLIgjf9l45QKIthj/zwHIQ5FC
PDFhXuKqFClVdLZmIbfjKpNbpNC1D/naHCsCbEm1cFFkh1amJnfAoYEdWPqXRH2t
zXA10K2QjKT/Umj5QfNjnDKomhCxQGWBxXdjJXkZ7jA/veuNnAwr3IhSEBRvYftV
GdVbx6ECpk9PQ3gva1lRCoszrZXcL+sN1RmLtrgZ/RqbvkSXd4xaUfVqTN5jzgSV
gHSiJ7zSqpg/fyI2+6oZxSMYyZWBdc3nBZHQ8SAh2q5UY+cRvE73/4HmLN9mJWsh
nuQwwF58uamB7MAia88uhP560jGxTpZAj/ce8cukCJRrCq8H7BtenQhdCg3eBdnR
4FuU2e3m1/gKi3EGRG8tkOVsVrSMfn5/hWvlG+9R910I2DEjYpRPED5pzh7O14tV
7YLFBv6UzywgnNb9BoWrhHXyt0V7DNBP1z5zv4g8wFXwkr6Af5L9cQ1nV1pUssZL
aL72z5CZjCBEk6aSLbGetS62FPM81dpvUSOfXEZSt4OiC2Fk1jeDAE19yNdFtJm7
sMFthTat4QRpBmDzw7a5bM3viVSVtTkg0uG+mVL95X3YsXFbzmYnANuIpxwAghgE
O62ORuChUFDeX82kZm8AyOsDScyML2quyzVS/IKzYTc+Wq5YQ4TcoD0mfGSUrHQp
2YpR8GWo9F2vA4cxFDhZp3vr96zsyTL6RrATs0gIUELFcREeTLQ2L0y+2feCBOjp
MEibZaxedVMx0aQP7UsTbb1EZpNVECks/K/Trix5CLDGaS0WFjcOj6/9+FjEyT8S
xYUmlxQqNbBi8FpfrgdE6jrHBFZo2K0yzbzsbf+wla6U4WY7AGJbOUdIZ53U8LBJ
gAT2B6uzxC2tVAmSyGr8YTYHA4/FVvy2EydU/0YWQP7r6L2Z0+HUAZKegGKYDz2R
RTFAkeLfDrBfNuOFt/TcPF2U8W2PPHYYS+50aVYYQNLPU+bRbf/wGxS5s4ZKWzy9
MGlbxkeUsc2dNm+EF+9tJ+Qjwa2j7jHYEAk6JjnZZXn2Nie945+2IJxjCOpbpUOa
vjhuW4xL6/erWb9q2syBvgEhNBzRQq//Vt4Z3faf8AB7kI96eKW7NewnDCTccZSs
eY8fRQvNDmzg7Q/IPr3QEOsAFyGMZASlxKyy4IUXujr3MMZQJFoKXG/MUYSqxAr7
Lnt7ope4Fc7vKW4jukB8mAX3eHrf1b1eFl7YYKjWYdw55RrX/KXPzI4GUMgLP3Q5
g20EQI0tikzA8erYJfyuvJH7F+yv0VS83bNC0KjQVgMkLLA8bzW5Jri8v+HpjwZ+
EzDkre+MbHrJRWbAZI6Zjb5efBCzXCaG6LnPdfYu5+v+YOFx1iC6IDgp06IyjgoS
ihKPY25cfi0PV+mChQG+uYEI7jjNCNluNDLQLGpfXWDg/T2BI3Zyjco+sx/rYFwr
Wtd2tM6cZbpus91YP7kJqbRD58cmmqIVy9Ldk4HAGqIS23GYxs0NvFw5VRyErXBH
XVSRGhqtX86zg8ZPetbJY2d7zlii9SS2DpkeBuNzhsTfZLN0TqtqeiNruTjQQaRR
6vClWZu1KvNtXoLPEgvc9hGgQs1Xi4H7EYIicbVyaH8KOAkP4hOyJusUc+mm7cfm
aDESRd06xmD5uEZ6aZtsKyRdjms8SAoOb+9af9ECCYRsI7fiMMWHClc8SIW4XBa/
Ku5ee2Ll6MW9qmOJb37625pEP2mNsJ5zF3EN5RUFtibz/wE366858RfNtQdLtsnC
ZAJb7WR5gayPB5snpQ8fYWu2+UV1O45fyztHcYHSafA5w35+IyV9EcKvJCUUvUIm
hLfhrXfz2RYTcI48uS+2Mn8NG2FyTr0bp8uSMAQvRCD+9D+oE+EjZ6spiPePpvLw
60yi+IlYAHYsPq6B1hQXFQ9EG5vdLZqnlcpu+2V973FHl4pzcfSWI1vs42iZYNtE
2I633vAEDMe+2kPfztXMDAWX2MxSDBAxiWtJNW7EaH9z83UTlnQ6KWFNQ21dXcI8
bGeLN6h9w1IQYxhU5/VRID31ELktSoavNPQLgg2MMe8+RWMhA5P2Quv9sCNk1kRU
T259s2TJlyxlUjvsWLhEuqT0kxHQVABD8g3o7gT0/NDK/+/3bQ7UhOpFB5Tes5/I
f83/c4mvmsPvX16AD3CRAYmZiVgmZ4e/fkVXVVMz5kBgQ/fHWXZ2TndILBHwQhQ6
9pVxg4NTAceAKg0ib8r7KRY0Gxl9lQk1TMTzAwkzQMhzevNjuCa1qqycZCYixcMP
BJY/qI23JMV3SCCAV3Rs/PUQthfSwRW7ZkDdhdn0kh8z3E2sCo1oI3Ab0Pv+fmre
DcyH79OQ9G3zfvLq/H+Duw4dbNblx2KvVn9S9PnzdK2I1v6Fq0pbpcJnsbdiTvTM
E7LZW9hOpo4K+mm1aTh8ZUYvVm22yEPWNckH3SWnV66sw3TGQ5Jcn3FaAFkloYZW
mIV2kcsMQhFm8+0gJJ/ZFVrWAwMDr7DTI7dMj5ndK2vfls74Q21sZ16aqKNw23nW
JvevRg6uFOlZJvhdzutZZlJ+tJHYFho+t9FdvJl35NLra5W+pdATwU0bhu5Jf5Rl
1bcSL5b2I2XGydG/gFMtXo4X8arLRo2Ry7g4FVAIhQf8zEz2iLtN2S4J6HcC2y8s
7lxE0oUZ2hOkbhqmp61q1CYfWcFLLT9vJLDm/Sh9KWx+BdkOsWVof2Mqd2yCU/9Q
1pW2sInepq/Hy0LJPYChJwpqQrh3GvlJ66CX3rwNiZCbzRsIvZN/lSUwq8Oy9YcN
wGreVE607aiV/oC9KfgzGWOHnct2InPiM91unBFdnyEnaybvrpWcCp1xdqCyq2CG
XcqiOZmzxUa7Im/iTwo0R52nSRM9gnKFsc87r5BSrIUWnQ5nikbBGezzFbDyV4Df
Mmwa5cK3zFq1VQ1GDqT73MBkc9VEUJZmEBPzOYxkJvJ48wgyQsBRBLoeC4z17rg/
7E1lwc1fXtrxs571qzI+kHVljZpA/1ye1zatP1xIdfnqUJYrY1xji1eU/X7gOhcv
BaqK2oARpcJVFMe1pW66XSb+cQZpDJBpz7eKp1OHHsoYY5MfaWHDs7PJOK7zTF7o
F/abHSJleXbyfBw4ouxLu9YuJQeh2exaVRbQ3/FiEqBzQ/BpFMzOZlpQm7UGnnbd
z/f2xK0iPEP9+hoXWXZHsfBC1j9+csw+fpGRvlTeoz3QH1Zl0DfD37F+0R1F14L9
vTeAPOC5ZN/kkgLNlEzWFiI5K1/9xXYxsCNAc/LFF7sXgA6JO8QRpzFCXGBiVP5E
JcObzDV5PBGYn++GP6Z2Wo4qaZlAW7m8BlANZEqkTTO9UAjO9b9z4UCtRyEZaEn4
TZnSfdUB78Pn+W1i0j0TrfwQ1Ungz4bfPGrLALnRmNvD039S8hlpBVPY3y71lY0b
Vd89d1J6dMY4oxkIYIeyYImc1kX9/jwH0RMtlLjlqHNTMi8sUx9Uw7XUM9zL6vxL
BHoDkzCE6uKuRxDJ9GfQoRwmOQBCQPKA/jO7EDVEEzKIIJ999QfhcNVEnocn6gcL
pmcn48fW9wIIpnNxtMtZv0LvqGjjRgaPPIgnmMQhOsyM/snLSDHPo6mePeAKu2Ao
mSwZjZGKbUfz4G5ToaB7xfaOGVcOpi/7jcBAG91NEs3j2aUEJW5L43rglhZ1l8oG
3FSt4v4CM7G6iA7w0uUdC4FwnAfRoRvIfmuVkdMmXWLgWZigQ1VgyVccjKWP7Xy1
/X9IGOlzhUMQpPfPFTAVd8bQsOeKCLfNEProW5tvlSTXa7We+q7+2FffaP6QEF0m
5Kkyj3gCvc6dTKkK2ruuv81ZDv4eAv9blccP4/hoPKI+VuRlQEZ0cxlgN1rKmx3b
3BMzvPjZqKzSZbzQKdd+Wt0mAiKbfXW91sirVPWLdv+ySo/ym9wQtR38FilLLK9F
h+JxbCzksvNYa56XPoX4+pSbP8F5XemYsNWsfFKppSTVNa2iYLnwi4BIMok1QP/N
g3jAl8at/XYBZAV5Ir2pI/kRnHZiBaUZe/KVzayiLW4yiQh73Ykwgao20N0BKy3B
APOecdUWF5wTSz5xcqt5t+CNOGleJauq1H6VTMKRVR+0i3Q3mJ36/lvJLElSaA8E
VaUhAIMtpzybRMLwUGZmL2L3h1cBGrjYwai2pkvZqJjC7TpMtwKO1KZT6bqjQEx+
L/ZyE971q6E00bRAok0h/CMZY/BTAmb7IR2AAeA45sIU/8+xe8dR+rQ9ciSmboOI
RKY8rRisf3o4EuP/JGsohgF4i8y46+sPEWJZM5wEH+ZZr0NF6+fQJuaUh9d3nJqG
ZR6D0MOZwL0ITn3lQvT+075GRAwz988Z88AxePTUWowe+AsW+Ktk26QWtQSRk6Ja
5cGb83PwrppqfIEC7VOakawlWQC6NOOceGfmAOuogpdwK1zdz0opYQ1AcAac+zSM
ibAsu5OaMXkPfuKnu4SHL8UB21gQEU6nl+IhOYvXyhkFlVfvOAbmZUM7l1RK5F7R
hzEwEzRXmPSl/Sr0bCXy1sFLsVTWtfNcd/f5A+nmWFgqYfODMyvWtsFS0rjGXVYS
68w6p519Dlqt/y+3k81B2KcmiWV8Mm+yAzbQ3V1d3phsLxHwP6PWANOw2zV2Stlm
vZjFgL9XI47D2/ln0Xyf1HU/gb/qdo8Sc1mW3ZCQJ8fqN6qTSJlmiAPYK+Z7h+Mb
aWsm2wl6qw68ylpUHmzK4lkk36QHE5R/Lj8psnvvVd9976pZ805XNXwd9KBQlIUN
hVrA7LIsWK9c6WTRwK3RHdC2+2pFSjgmcbgJ4W6x9vOTCr6VEsfVP4Qxxy49GYZZ
Q8QnH75JWDJOmajaLOMeX1yknEM156K7fl04tdWSrXY+zIDE1AD3pjLZI0TVGWRe
et6CkmHODUZ4bMKjaCqU00zu86N7ofqunS5yMikYrN2vQk6CfhnCQJFfFb4s+ZyK
HcIE34KzidoDY4Y0XA3Nc+12vESkbPTydyvSsbUdcjpUxsjmUJgujHtw7hnlZG++
VOa3ceAXAEZ1Yjac6xIVlC8jend120JjKC8edSQwaU0pjiJ7PTJf9KZlRTH4Xx1g
2qXrzjDKa6HtEVF+5lojoxoNjB4WP6SchWzVrr0NpebV4qTvrxXOIIb7oqAFXhBh
WLvi7pcPbSaCFHmyQUlsHV6KZYJYVbTq7qmgSV63izHtRULG1EW4DHAdMtDSVUdY
1PQOHQcaYSUhhlD+VL22zHkygzejh8u5RvAkNezh8t709OfTdKKak/kwdL6v1HGx
4ZsDbmdzdaGWxxkk3YFIacZCrF5fSaX6jlwnYtRkkqD4GHMYKPqbVSq0toIAG2ZI
+x1wndfGzXeX0IrgzWtqFf3BMbQJPuar5y09Yf6ggrYv9i27vX8PV2IsGSjzx4ok
Dk1HXXEr0/m6jc3p/hcQA9A6LkQ46Qhy3ncldxq2A9USdby3P2x2T+7PmQW+7p7m
SHWrFSmGyk2Dr5olLLw6gvtFOdHoDP2IqPsMoooOk3Pm6ikHtrNU7jMi1N6h0DOx
D7rC3caqk4+MS1VTgR8Wr7YvcfxpxSldd5xEnIU4/lMivTWhWKsIaRiSc0p8ZvNv
gJSmXxbs1encmVFuTrdeh1FX3lqPRKmIMXeqi2p2hP1wk7tcZoWR/DEJZCqCeSDQ
kJzjmuzLUI8akEThsrtlqdRRDAa/soXMakYKroMY6H5/dbY96RYVb60C2sqnZl3H
sgCI86vlX+TqDpjdEGlUHD7xj2q3CGHF1b8ZOZC1YoDxTAkX9TZel33mGMXpNwbP
yF92WOzd8izzAybo5N9l7z92f0VMy5cnCAMUmZV079XHg3VMzvkT0hOuAAt9isY2
QtipAZc5K2uyDbLP2EWn7tVgr97NuoSepVKzYCOq2kVVeMgOsTY8+C/nHXp8tCHD
60R4GRH+GCNoZ/th9f/cqz3UL9FTvVAexljJC8AvZ5ZbayhwwismgWVfwGhaArTE
GXhkn1xnQT9gwrvRFpPXdCo6LMTbML36Mv4TXTEPVt41T+7NLOla0pjZLGBS4ByW
HfFb4qSnotkT5zRdOrIDSqUNUEAXBizds7Ls5SiySLH7NWOyMtymSNoqWFsHduUA
vZslI14UaYGrq/Ehmt5o8LB7ORQwwMi41A/szvAj3zjZeWCMhgy3m0kxNH6UUNKs
3iZ/RpckOBwRKYj0UFmUG4C6Gje4cMRe6br1Uo7IeQWDC/a7Znxm8pkhCAl7xhp9
k/PTF7ywOHMAaiE++zGIUdmByivepje645cUGbp88307lB7U5VafQmlCLNjsiEbG
bg1pE/qlsjt3a+SWALC3ccUJRwKP67TVCSwhks870Utw6SUkXFaptcRdsX52QtyY
iE24SA4FupXn1/As4uUL9X1xjjiZ4MBRzIlJzydXCa9WIQYspp9sf9MAozLFPrxb
LUDyxlyh145WDLrBuSYdQkQus8fmKT08UAmI/uXvEMMjaolN8FLp1feXYQ231aHI
XNQmi+rjXdKmfH6/OYty+st8I0Poe+E8jfHlW3ioqzz78B7vNtOBNK9oS7op8DgB
qjcOqnzglLx1Z+3vteHLqIkfE+hnTFM/dhLvzGadBWfjIHf/GfbuvRO25KipEUP5
WxMuTqBxUPz9rhlu+E8BC6kb38gaDRC2XzKR7MNg9hWWSp/shbzk5ruTT5r9V1zF
qfCiRUMCyVimMClmmJeHjlhyirAx9hJWoaiirzwb5hGxVma8zycyStb33MO/O7Oj
mXcSp9GugUZ8XFk8hLtGVlK0G5N5LnALsvrWReig2v2buXxqd2F3+/i7kLoupdSZ
BDVwsL2fajdcou4lrAOZdL1NAwN2nq13CC7sl0bpebukZUoRnO/zV2uAoXkKwu+t
M8BPlQnf1wNGOw0WnBJFzCaUv1+B2Dz82S1odUwpfS7s0+hYso0uMo3BMMMfL1VU
9671I+DV8GXVcjlI2QKEIPSTti/hiROOexTJBKg185+kSFDn1Ww/ZyimYEVHnrmj
CbuAGHpXuQXJIvp1bEn+iAKrkOZEhbCuxMgd0cv2UlOHZ3NwUTjyV/pPTpkbaheF
7r6DsMe3PMuDbsYTnNLORSGzCpidThzFGRZdmN6+LOnOsvqj5o5+lxU4KXmPlxcm
quMxllZ3chu31ifj/dXjEdDBD1663dk4tFjBU4ah+k1S41EUrodg8xySgqU6cFDE
BdIk5WvanG+s8hRjYGWYaRJvGJ1AgxQtJpEaBgwGZW0ADNWzvf0Hb+ByiITthBcd
TKL7tzh8MIu4fO3IqIl6fTkgiDmubayoluNgi6AA80mQoEossq4X97yQ9NHnvW2V
1KKsFANa/3mlxy2W35Zz+UyJ/iSLrHJoKK0jW8VfyXM4QxsHfOf72RJaexp2QhmK
K78BI/gngZM8t0vq8SwHCg/jv9K9zCioZtEE+xQ820oiQO3fci3rbWSGyDfVr512
ViJVb42kgbNKBo0cmFpFcHtjQ5oc2t89ztsOkTxc1Crnx3DEpGhQ1OXM6iI7YIYx
NI2XRjKlH7TlVXiX58bxbWTjVTW0/Dc1GH5OUAO0OfG7kO6t4PA3ABoy71tk7Lef
Yraye6ss1v9xyEQBrkOe1qmGPtOwacXD0LrDXalKw0tjLU8QVSsV3yQAMv9veXz4
be+b5eJAeWO7gyt6i5QZGbkgGqBwKcuXv8GMiSBMzNqvE59biR8ofGAWlVMUBZZb
IAfKrSqxwAW6pEPv7PVCUuk3dMiY1HHSi694mfBBtdOCkxjUjGClvyQtnKazzF5R
1vNrmeSw7OQt5x8+OdpOtnyIbpC65eaNt4aU+i7XlitYXHfMTMdyc5clF/28ca8S
LvrIJJO7+zqGiS8UbOeDSW6nZVK7aF6ce7xVnbDmjWk2zOZLha65Z7Z1DJr8f7ET
dv8D9Lk3xhwDVunt7G3PGfgvGU5t6gZLmkIpF3pUvIOz8GBBkK8NV+hIQmsXlsIU
Sw1P0uQCt6hkW5WEXQjfub3gcX4nXnEESDb6sT5OAzCJX2mZ6YGCSs2p2D3zDJLE
JQKgWGA5w6mLx0mgI+oVBiPs+uvTS6OpxdUUh7fYVfOc8qXP0w5KD40EFJLTvjdz
S8x/DasiSGAgTEzpS2InnVhOciVyxQ8ybtqV0kNn5hll89O6oDnCeGQ6mJ1Mssa9
aGrcRJlr9KL9iqZcMx/uXzsG5zoKP6JFHhxhEJZRraL9mFOz+Z4W5rfBUrUCfWOl
CqT0yKcptJBp1cVah8Qlsy00v6BWatkSzvR8JyiSEqk06sCpEiMMzqNPZ4DvF3mA
ZLT42P0Or7TB918VhXSd8rxAJZmHIwp0J+Kexj9IgTsCfp2wdQtwWqCZloPcwgTR
bcrV3gjmKqEbh5KHLsVoelE78E7UPVdTViHJinBSky6ZeGqSUCyYd9XOW/zxH76F
AyTBW+6V1ljrJCownSxT218f8T1oqbm3PXoeamCbHTSpVTeexAvUUFVeTgiKeKkT
BLO7HTML2j7OG7NKtkrf+8a9CeMPRb7oR1CgTJ2FoCJT2tnnnnEGo/GMhysjW41r
NG/TXO1stesxm8fmURbTXhs0xNVG8ArBNpiMpNVcZSU77SqViJS+Vhs8SgU6pCJY
nK57pCm6OfjJxfeOzj7ryDETDZfbrV4Ia2poz4f3J5My3/Z7O8SVsqDQRhl4II/5
vvrh+tZRxwAx2RwZ9W81gTyjGWTSOS4FAbj4wOMu412+FJUwoJJhRCdlYjbZ0uaA
IX7hvLQADWamq1YI2ymGbinAKB9tBkodWAD5xpp8xRI6L+TG4L1pBIORZfX8V3uB
4nc1awwzUwIyJd6w6Wagrj+lBS9wss2CVesuhsXQDZxpUJGUEQPaulz02w6cUKAq
FmF3SRnHbHH+EKR4je0bNoYLkRbl37Kh/HbjAoZ3OT0CEXfAe8e1u8IouE5CzBl8
4Mxt+4kQWsBjVrVTAmgXjcfe6swfmeIpMIOYlmbAgYkoZJy9eC6XaJeLccCkcER6
+7iKNVaIWdJ192w1L8MT5zpbQVz/4uOGiZeu2GSirK51DGYb9p0uWi3TS92Bn+jp
GBwsA7LojBeCjJOjDZlR3YJYyXCve7LXr/ktVKEw10S48FASGbf3kQ1UbFULula7
3xE/fIQQHVjMk4HIm0JDw4p1zjQjfeV16jUYYlxPOvk/gC9r6lZcs5qOAo2vMmVs
jKaQOCg/W2+Ps8KyMhqS4T7jLKK+pOgwIWEV79kTEsacbtf6HfGQeP77JaTr7rds
2+cTbePFdjXy58VHBR/dNZL0SQZwjLTyGqR7Hu/LpOipk2B7ju060O7ZRc4T7Xc8
hw2Zz/eW4LHMq2+y3SLgO8pcwcCL1K+xpNnCoGXrevwrILDXGPgaNwafpu7dgbgK
hDR3cDv6L/dEIFX0Zgj9gA/uv6Ko+D5rkCwEG7hHskkdTrtor1NClG9sXE0i2Fli
mYCJuHTylEbD/a/ov7Yo8XyiSb8SQzChcFie/xuBM2NXCLiakIcK1V+TFZZkOxae
klBU5g16XxNH1U5/NHzebWsi/KSGamsfPGErBcDpKiyxMKdY+dJbfD7jrBG1yW87
ImSeDJQLI9vxP97lfVdMQGGQgGTUzuqWDyO4MLiggzST+Mmoe9lyitOM7Z9ynDNp
A1lxP4JOpRjR9mLZ2mipiLZLOdhfBPC7b82URySueAUn7qtjjDNoNYBSm+IojbsN
UJh8j2eX15RjLPzjgm/dhwM2PCVP6M6SC9yOIuFBwhL4RmkGXxThMpJBllHce1rh
t7qtlNz6H5DkKjZKYkwS1sZZtnm+lwhrN8f/wLdtQAROgMe1fWs2m92Wk4kb2i+2
nuEhoVJpX/XCLLTuv9E9yNmYZd0zD5Z8I5M0+olysWVX7YIz8ycMOAWOZbPujU8e
LPlDe/BvghXujIVKGmXx4G43dXWF5jIwRbU+RQQ+uDAbs74PDSsgYt6oMzkA+J5a
8AEUtVBjWCZUBpoaWhDujDmiSv9wQs7KacKrp94HMwln/vmxZ2f1kKSdr1iqCO9O
JyPz/tiOiSpTjT1QrOWCEcdW0Rf3JlP88tQHhUujdtiM5iuOOqYd0bpCUixY8A/9
pusyDmUGTOOmb3keXe5otPijogPgvMLftXGQNL/b75fw91sx9sgSdkgNHQuF9Qpk
jphZdzzKiFcCN23LzhmuY1aRyYymQvaFXtN5iK3VS0USOAbfZiWG8+DjWFyBC3/Y
eJYMv+OZVURKVzWzUEMtqP2SWRAEm7U5gAR2+fC9OcPKZUlLMZ0CwT8m1Azs8ikM
jSJY6vHgF0XAMo0RGSXHiHYhbg3//GQVyOmpawM/JPZ7xVEE3iYgc1nZXNxni8uQ
itY8XyZBDHe1OU73f/uizm12EHYrlvgDqdQ9j+M/Aw2nVNzjZXRsuORv/1gfg+qG
R0yZ3CmqTj8484bQroNrGpzoqnvu/s14tJ19V7yVX+kl1vQz92H/3Fxz8YKxZfDC
U+HFFeNMoS0+SWVk0ffKbw4WrP7YhgPQcMutlcK+HlOhdlCw3Vaar1v9TonkRHU5
jOtz209rSeScvBF0G9lqfBe0aB0DgURaGUKuMJRNNgwO+w/C3ea40l51Pmtn9l0x
8N/Ep4FAEi6N4DIZ8Wz5R58CDT87ZyDtUmVvHn5beUbq0GY7aalRl8O7rCIkVS7L
foOWhN61W+X2wiFS5rWq8G1g+1iyQyXRV1uFg/TyTyDAzf1HFbvHHD6LHKlpPn5B
nrcXz70XL50vQBTeqsrhXXfqVo0xIa77k1aR5tR/HcqRl2XtCKQh+ktFPRLOwEYz
djMbSrYMu4ZfVIyT1gCS6WQ5zHSnF5xNZ+xlLCdMT4gabhjIUYEcWLDzgNGVHjyx
ZN3c/44Pe9vg+k4u1jcexWABiQwcXlE7FoTUncT+QQx2FMZWVoVOJiPR4UMP63nP
AkQoSngePkE2i4bBqWESPWFg1NvOR6Qq8IvSCXfP1CjZWVpePJhkYfbiV7r7oJKP
aijc3J0eNy0kxx5dNIFuFobY84no98Af4L2Cfem3Avgh5Pv9fa2Weg06dsMeDRRh
OrzRwaRAM3PQzqsqpdr7yWTYn2nWcuR8/pS7Wb+JSqHZ/iEt73xO+gLWCAxam2nK
BImbEvHlWduyt/LvCgrXrp+4iazMzOBLCscYVFABoomRutXiZdE4y4O3R9ns0KIE
5FOkY5s66ZzLv/CHN/UKCQ2O5R5UCGjNYh0x8XOLItDJoRjWJvEKGuimdzYZ01NA
fX/DO13/zohMbKNL+YZcK5Wa91DxOn80DmrT43iMsXIk5DCOXCOPUdasVY2R4zE3
J7phfWvFkOxm+4k1H+1EAqKF8tXgObSVJfIRgPlLYKi0D8KXoO0h1M90FIhrva7+
XLxR3aq9lJ9orUAWe+PzzXOfIPSZr2LQMhGU5JTTXpxEbCPEw6F+wtKoWyqL6rsY
soLuz62IpXK7R2895kahtxQGr3p7VyHv6v2j1XCggy/GPkxiZfVz+vK2elvndbWD
tGgHN0xCOM7KuOil3bZZgSXgXtNo2JXGVkPEu9diMUNryZ3fep9QZtitQiXOeADO
Sx8JhHdLzAxQskHUow/v+u8LC4fXHJR5oJjqu7MBhjUV7hPuwUYlWetLDcgfmhl8
U8vUgr7Bv+1uKL91wP+o3q6/Do/g+9bmBB2mf0WGgkRjUqIPe/jLWZ4kNBiAvGhl
cP25P8d9uvxbrlxAuW458tn8a7xkOCge7rGHsAXwrNi6qKFeQVjggSuiz93jlc/o
jjDjvKAENisn9qeBcRxlUh/8LxdmaCrxRF5BC9BI+V1ey3T7Lu/aIYhewrky2I0T
ybfS2pbMPdxcu4y/MoEx/cPS06HhBqpyeLQ9W0eZFnR8jP3aqj1LVsfY/emBqn3f
GB02OsHbfpGBPJlQi7HYGqGvqAzNMfuBzG3lWlQpjLgT/qGwSdsKz02wbecA27xZ
fTYgKgmSfFJytOMmzFxwbDnfBOscXLRgErIvipZDrtSeOgQosAg2Gr4Xh6LECfWI
KASg5w1V1w7t1VZHC6PT5v8aMv4CQNLxQzfZ5KELP3dCbeSmqbSjY4gpRMcc+C4L
fEw44BCGwV3qYx1ITGoj3ol8+XTuCd5lfuLcEN1NrbVZ26Q6oI0bzWYc52v7NoiO
Oj3DL2/R0+t624p2armtLXjnrqanf8bXYNGQLtfSQSrLf1fh9NKi+6OCw8ocx1cY
Zor8yIDCJvIXRA7Hc7One9inzqLr1D/JfabVSv3+hd6VcaGFGhLtYq/B4FwzARfS
YsMhsM+E1VnrqNB9NGljVY1QySJuP3A9phPp4ot9GOOt0pOUBdLhQ0EQjG7ITo+q
XpAWjmqWs6u3i+AOWbl0q6aRthMb4yShUeFhrmKzimqaU1R2QC0NZMKPyiMuU23R
ak1W0B/zKCvUt5shiOghpzRjfNnvw/pDLTgOhk7pIe5glIRRabTtbxoiaxIJQIp2
5eLFmQovvoephCdWIPKRM5f53WXOczYUkD0sTxP903rnJr92k5zio7mDacdCrB5h
6qjRBOkXjwdC9+nhshL8MhDIy6/w4cLsGZJQHHzffSMZTPsQ3Ez1c3if7z19cPmh
79UpQ6nFJvcqpYbINAaR+keHYaom8T4cU8071g6HvCvdrpkTB94UbtkwOapToiwH
olMHKYiqHWx4ANNtdD4jZ9Aqf2Evh8N6Uqp6Se9Y94nBhrR3554hfxDI9fPrg+EV
wIWChPqkcV4Gwuwth/GlsUJmdmDqOMxeDWhi15zyyTUZYd37FGbTyS9I/xdHKDqC
eUDA5d0aTGDzQNOS9SCvINpntjXU9eLt1BgHOr565DtE9uBRRLz//k//AFEwOSf1
B6bnJld5tkHkGSC0AHjRBqXyHSOhnmHn+6heekZMWU6FiEFdtCMDdSe0/FSeqqpI
EXfVnPkXNjtoZ5fOeypGspBgcT06FHL3e8BKU22E8eiZVopbyvAZGMA7u1TrY8KK
kd2VFBE6cPrzyPVSBQDXGut8ykOLjafxlf74iUf/5lCltFJfswo5UqsvnMEJ0ms3
7DoD96W4WStSV6p00KoRBy8k3u7ozxexvSDEof436IpztO6B6mLBFTDfZ+7km1ND
cMNQ8G+s0wG7Qsv2KBWrfCdXeWN0NKXpjIZVR/lJdpp7MdbA7dYTfysLVkapWrkq
6/Hc6Emt2GsL5WquQY7yJ5xieZ3g1771x1txg22VEA63Te6d6sNpNQ2CunOKe3Pk
FyFVSRhlWTX0o9aRdrskIlUDkKn6csPAqHgEw1bSA170gMftQGogIeAUerCXrT+i
qfZbsDZ9By3lfQR5fJpCIS6Q7ZZZ5JrsLuVzWDAMfXQJQ+2rjLso/ulR0eQTFM6G
h2gKBLr9hrFIhBwxST5XXY5/p/Fnfn3zLqzIwdILcOdyNQ3yX2Yhjtu/C0qJh2Q6
sYWS3phOFczF7RGTDpa9mZrNsHr6cA8DDo3/GLp2hF5GWU3r71YJ6u2rlARJe4ey
21YpqJW7l0oe7PvVZCql3pFVl2Gq/flOfZh95P2Dba+CTqY0CqOV8KMx2IKfuSaQ
eybhhqsrPKkLoeZnEYZEV7X6o9TESIIEvhoLpiRQ1i2mEoHemKkizVzpQar51sJ+
YeUuMsChpQ/vIyLMSBrxHS+thJjE6aEBts4cElPE2UkmlyYInS3/5L5IjNneXUvn
eKusAgr6f6c9nWgOrtm9r6D74TZeZOgzLEojkO2dMvzDTfXUPpeK2QKNn5faGFhX
gnFpdfCW2NqsCenzr71tAgk1/h06nc/EGIGuEqP+WJdfLwpX4Rk1Bd6dYlIFZLqS
PCE+zacT6EVOZcr4LBz9CZnD+7oiC8nmlFK76aJib8fokleAJfAasYUZFOMWCuKc
Ym9CeXpFxR5WnKhlCdr41d424rp41yBcsDkiLMpTa/3RwIuGw+PRO+Bu0LD1GP+H
Vd5248f68N5Noo3+S2VfcVm7b0FJ7vb7VDqdJfF1ax3NXojZa+7e1XVT4ONNsurp
je7xS5VxYdLGMNfkJSwnn7jB1imRiuYUgIRiBVTl6JCCWz0I9Wqr+8hwnY5LJWxl
89Cgz7D96xBwF11gWSd1IU7ABy0MePAVpTDgfSx7r+IrBBBR/U71/l4XMIGdhEtZ
jSw5Zzdji7rDfqq6ov+6T3jQMMofIc5BrGQspN3Tm5st8i1gvMey1LbmlC7winhM
TfEiKUTeToPgjlOLHIp7oxi6YFNTntO27eyTuS9rNeb4tuAAeW7o0s05FfZIx2/x
NU3l+lxluXXQmLCay70Z8EMshpsq6d+HmrTotfyVb+NjUe8aE38HNIY20iX9BpKf
VxcdRE0NYu4VAqZddzIuPjOU1MHsfpBembQSkeLN9dEo0AvsTB2EqUxYxB2vGRyZ
em29hQ4hQoWAqDerEUCwSefzMCnnC3BSizvCXHaS57B3uLmqSZv7oDAMNjtIWXdy
YIzcRoMSHk3F75CILdVV7TYik8yTozMXAxlXmv9kOdInZPBHnknVazf6txCeRiUI
AcWNiShFpQ7y58sJGeagRdmHjzyliAz+H2CfEA00MJU0yZ1FmZX+NBzFfVIwPVGQ
KeH0ygpEAh2Tsh8SgcwhH4S+PUaa0kQb4tYbMtndWyJhl1KU1CYMTsEFGjDCeMT8
t45QaHX2vw7PbHdaUEJRH7Fshr2qDufpGRmikXUv9Kzit38spZQwUxSrZVxdYTK2
1E0N5eoF4HH4bEv8zF1z0rEPz+SVWnI3ttZrqAuxItxP7QoajpY3g8TE/j08MVJT
MEp/gRaBCmS7Y+u4P0+Q5v+8Cx9YqQgrxWNMZT2q/iUPSAELajY1rnw1gUsVpwsf
RYpahV7L0/MT26cDgK80FdHFHLCLI5zJhR0PJb/y6jVK+H9OEYuMCc3zwI/KOZeO
sC25WZ1FZHPcKaOIzlWXIuWUMgWTM45EPm3IlCkGB7p0SVe+wP9cSQOKnEU1lGHy
HNvwrZach4rF97gtoD0s4NehEEHa2eu3iZQaBYUzjcHGv5gOTsYR6j6+LGdfqxwM
gf6nVxMKj1evX9odc4QV1UH0fJ3XNn3vg0PzWXtIeNH35iPVsLTZa/sDD7k0+q1Y
VxOC7kRYGb4b6vo96DBqmHULEAh3zJ+femLYDlai2zBouo8ODs5r96lwulvEjlGt
Nm+MPWKbnmEwmOWTgiBN7JBKWlhHEnxPer2QKitRiPv7QaSCft2wGblIrwq88Auh
1vrCD2MFBuJChCHTDaL/4InkS5umyzZYhR+dMzNOhw0v7IkcXbouTrjmpDFqbjJU
Z0wl5BFogu44jPhtA7wJORKVBZ+NTVr6U/OyQfNVJJ7y7FBECSVsJdEfhZcNAbpV
bOAsveaZR5TqfPuNX2noTX5K33SfrAw0z/SR14cCxGbCC8NBR61VxYOKGmkkicEO
SjodzD05SJ4G+bIFL5qD4BJGS0Y8Udc3m/FWOJXhHtJHJ+1AThj/uKzEZfeovWLq
+/ichfDJba7tE5eKMqYo4NG2qhKRD14buBDMV2eBRTiEfGY5x36Cp8goNYmbFgkd
v0i8xFIREroJ6aVcf0HGt4FSAwL8qd4KTAfz8n+tX07Qne7TUd8/87tT3F99VWX9
ELzVT425OEJb9875TVU1mJyLwjeR1xnn3axTiW76GBgN9CECf7xH8BBvoUMpHsJ0
Wfa4e29eqyxDuFgITOC1ON5ykqYEMlB6y1JPevXGn/vsr7CMyYM15f3KMCgZ6atH
qywPXat02LBFZDp3tun+yztzZznWig3S582t6WwgoaYVlTJF0KfJ0XqYhDBmYcNi
FvIl2jEiU5p08a2QCzsa8uA0Tj0R+DcprWzAdy05b/m550NZar5TMYIhiUH++SJx
2m3Ua4VPxuj3FD+WkcWkG4MiAC9snvCr/4hgoAUugCB8qJoF8ZKajvx3/P5M/0TZ
wLo3KBzSJIMq5PPQXAC6uotSntI4bOvIV/AuVxCrBHZriumON7E6ERTf8ezwPVfX
+pFl+mrSBE5G1WjZHtoI+YJOHT7KDGLpROLwzt2vi6UG9U67ucJ0j0LKmb1mFWq7
EAkB8UlA95RgRffyMmPtWmWLSEcEoGTggyAoWjI423S1U+g7KsVAH9gWZfj2i8p5
D95kNpcBXxk4pIlbQ9JFrfniE5RbnCSZHITTqfyPvJrJo7Wndyj+iYAt46nHjvwF
Iu7wCp2nugufwIJykdGUOovgXuFwfkRIOSQ3kl2AD2qGlZh3/dk9pZwi+FVX/P2N
jexzBQfwi2U/lUPT/P3YVcOjfgQ05xwChJIiahACqoa8f9wSdCOyDQO/5dPuPiUr
+z7lq3lrTkHBft5nztzM/t0Ck6YtBqHrmwmACTMdcO1kRXufnEUvIgiDFMsg60bX
tQz+3HgMKNnqk1ILzQHGaiS3AxoPAV5hp44AYp1MAiVpWG4XzktanqF/46xofD1F
AjaN5vZJBd6EcA2JOO8GC3Qr27qZpnnsSj5BoIagjD4TsnGr1jb/31EaWTp50QAV
V+T+xJyOqdy2lI3a4nKKByJ/p5CMf46DLsij6pVRgB5DPLvx53kzsUDxI6a9i3bN
BKlhRl+jsyTgNXgQtkbhmJ5Ilgi/BV2K+LNq6StcFgwACx6pl9/NycOAc2YVT3qU
K2oe4C8MZZj71t9eSSuoUWjNqanOjNpHtfx9Fj1TJXsxynSB4owp7cwbqGuz0kml
Yjp78HniLdvIwU/aJnNrDiuDte+uAKSVvj+NFrd2u4/UFCv7IE+jZ/rGIOHX6q/9
uEtK4e7CNjiXvMuxihEIQwCYWcM1JO9md1Nb8BRCTtiSK+HrCp4pgU50HwbCtX31
RLqPuka8bjs60bKcfo+Zs07uzsrY3SLYVy3skXE4dxSp8SSvOBP5f6yvhEXV5YVC
v+WJWiVPoAROpZbUvYA520L9RK0HpSiCAD+z5WtVVBPGeFqS8dHO/1SxWgaVmlfB
fZwxJsF7pqkd3mnsynEmZqhhc7KkSIgDmIndSdbuTbZxjJ+0n1AJe6rFk1dSt3OD
lOL1MZbbKNzS1FMLf7LQy1KAW2LHDP+l1dtvrwnb7+8j8oKFdVoGHnNFlUIV48Sg
nNWYqSy4cCit0CPu2bEk2A6KKDvItt053H9O6MaRf2vVqbIgWvXTW7H3xbolDTJW
F1ki69ND1Y07TQLKiSiDTFC1FBQ4FdTRKih3gfd7eVGCKEORph5C1FJ90mToU5Oq
n5KnoFd4J6FPjoS/dvlV8oAvB+UE1Kcej7zQG72cbPY5mHlRL779BE6sKFEgj88R
woALNuReUcBvFdl5Qx+dwj1IVVNEvkDRBNNgTnKS+sitR3UYQh0AX3MxTR42CD+3
PUWsY4gYczjOCx1Lel8Ped52rju/o6MwEomm5NKbxqbShUM4ihfcBYcoJjPKNtWS
bZg7NUKYeLLmI7Yyt7zYFewseP55taQnkK1/oORViKvWN6QVeET04jVDC9+Gwrx5
6q9z4Fsf70RaYzXndMNfTdMxKp2bter6tfC3gARB8pwYK3R3OYcxIeE0yJ2VqyDn
VSm6jA5UDH+LYnfJuvdyK/fstHSSNdnAHD/yuoKj/bCwNbyM3AhE2e7Uz+Jysu+U
l1S5gdYkWHAK6lDNoRopQwK+hhXeK3IYIz9kA1sUPVqAf2lEqszd67CpmMjl24nY
Hb1uC7IcNlC71Nyi/lSzPO3pyiMx5fXTRHZcsJIJJXZqPK9db1PIy0LzbV7ojGSu
a6VFY4s+8etiuzNsMNoN49IuJ5ixmODnubsJM6RmnMQ2dcHzEbc+dL44I+dB4UBX
IXJN939yBhAaGrpC4ZOLPQbNwujQ4A26tcja+TvcMb5EdHu/x/g+HA2WB282HiZd
psFvYn+bEY2HXW6dZlXYvVpNqHeSe1ZzPD+IU/GNzjJCx+mIgxwC5MRSQ6yIkeNJ
jrcmm79b1VWqBqtLLIaa9LGcmrjqZetcRK0IwISAtSF1zn/zQXe/t/2J96UCO3bc
pFZZYUA747qScoBGBdd4aFU1KMfeE4LSqkQe0PtI3uFe6m0owWjkcoqhFUqE8S14
am0NJqytEALBTLP53VfK1E+X37e3Nh71d/sx6/fAOk1lBjd0YEYWlBImpo7OJ5yB
BfdRsV9MalnfPTgmF6QLRZPTi2NFHHoUcJH5Y1iTnMKBx9K1iiN+yUa7HZFlxhYo
9bK64j1TLCOpqtLsZ2eHttfUc2nlcZDHGZPSrdflevCqolVDA+ZsG7lAMn8T7PEp
O9nYNlF4ik69iaQZGIR0ayOqQLjF2gR41Soy3qd/5KW6nFlFtzcILxPuMwrFSIXv
9/wYP0uq4qyZw12CI0uVR83rNnM0da+4wvyLFrwgVRmhFH+J7a55bU17gCz69tiQ
hy8NZaeJ9aPCaRGa2Ib9smj0Rj3fZp7UO05ukDvb3zDi165YV77lGCkw/aziJc1M
qqkjLkTN++D3a/7W/NwRm9mdwU0WunCJ5mXt/2npQ4yDnoyBE0UWfEn2Jba5FAl1
PkHPtipj0yZeCeMWqj+IscyyN9Oxpw9P16b/fx47r70kyLQIxFapL50JYpS2UYa/
br/4mL6BlE51YcCnPbkZdEMjDbERekwxO/LesqpkJ9ea5HMlLBqyZlmFwnsHasJ9
qSIS4JbIL/zYW3cEQIdzsqHFZaw7A7yICKqcKV39d1vZGfagWtWlCna6kwR9Ywb5
+WJtZRKuY8X1PBEoYFI4YOMO7IFcsbnuw/a5rEpYQS1SbfnLoY4BmhOdpYFCZ8AL
inSmTy0RpxnMjsl1p/nlmNX8Gx9lALaQrMwsKvuwkUFU6bNsY6gdWmMNOiygDP9h
bLpyuDlFM/NoKE00dQWiCJCmXTPcGfExBvmJI+d4Rnk7TdCWgI0vvQ+J5fcCLbq1
qYdj5g/+wsBeXtpOisU7xLtYbIKilHFHGhqExsZslS9P9ke0GjPgcUIES7SAy7lU
pBM5y+iLBJ7JPK7/4VIHBWVlwyTEO4j3hSBq4l6nK0izYYHv5OC8h+5pj5rqx74G
MsxSrKPxYa05vbbGc6xYMqk79LikdexRqFgxysa+k6D9utbXDqERkxWPvXCZssP0
gKXztrLQefbkhV0QKKmsCym3GInwy8FM4/Yoe1BvBDrUsQ55o70pyHseOrygCXjt
8jf9PccUGvH9XvdTigcb9MHVnz+V1e0ImZhmRyBdgzdDPiAcKq+o8L79+td7NRUo
iwdXpP6c6cLM6fGzpARhRASKqoM9HgS1drZobc/jN+sxLk0Dw1FoI25O90yzXuFo
sYMh5eVSKHNR5Qc6gmaTdMyk4Ns9rKU2zhFM1NLl8CC3YDKhelwxwJFAtclTksXe
HLcmWkcf4wk2h1+CzC730onHZlbHmFkKXx8UT+FH8FTu26vglwuT2mG5g/YQdRxH
3VBHeTmdZZm7zmkb5aO5GLeDrz7JdC7dt8ppl3nmddsdEEpXqke396qGmSNvbzBw
eCOJ7D0Yjqhpij/9DO1uaJRZ5SgB4W12bM8ooc4MCHtGAst2hwNBxeUiuuA/hnB+
9JFqLJLvpYG1DGsQYxYJkeZXhB1/v/4jOSCCwf9BFdBikZxoInW9/Gb19+m5APby
zZ+jxwdRhuBnMhxCRi9+1cY1sigfditEwcnxta9N/iVsRyALNCelmbGNTpHgFrRH
tLX4AIWvSOyGWr+3C8LPvedKQlBgTPt54GA/WWP/um42Oy+Wf/6gouEDjPjMhBvA
cjrK89cOchDeFRK0k3tU/8YKVQc4x9V/d6+IsQwZ3gB52ciOiWQJ9sOSqonZiRoM
GCnx5y5MwVJu9B/ubLvnHHHjsuRdvEnPT88Qn3Xf6NqyUQMlkv4nujUi3jS3M4g4
7AAkQR5DSVXD7Uh8JFVKTOKWJ0LH1uARRBJrrG3KcB+ZIjFMl7aqu7y1va5sYmn1
9Om2Eqj2WhxsIXXzcOOVHxaZ9hJhwO24paZpsMIT903yKksA9ZEPbkkncJai5gPD
X7yVDxpUixe/bC+QXbMZDgyLAVRax+U43SeAGI3GPsLhJ6jmQIZ/He2rDCbfaV0a
6qk9gvABntVRcKwwpVYNEb+RIuI6sfoFDsTdJOV4Y5pCnw9HqZpQNbNouAs8C0mK
rQNNlSb13o/wiPKa3IFvC5+G+r0eQGDFiyNOIao8dUSCks0t+DOZrqUVIfLMxOch
QU9Hdresw3rB2uSAqADpF4eRRo51Di7gUHWWWLepjdVY/2GPcCs/UxwqDKuFu4Fx
a2AxtbVN8sfM7tmzzyKJvwJ9YpCD9FWQ1YjWjqzePvMmBHNldrwT1aw6ieXp8pKY
Ua1uh+L1STZziFfffoGFjNvNFlK5HSJyvrGkVy87ZITV4BXmGvm+iApobQzLDYBk
wuFJRkZXAbTa+n8RbK3es3yS1Hg3QnjUlWHI34v2+o2p2Hnb4fzkxvfXI10g7SQt
jngSSTKSOkpN6lWXIWMPB/uejJMER+9N156mYJr8yTKNEadXQvNEmv2dt0+dS4Ng
IqcYpDA2rZw6mXQGPyOzvNGOyTwp+1rMdgQMj7Q8JwuVAMHyDp0WBA8vNrR6mFzm
cbIiv7JzdPQEF6gv4EZ40fWlfSM2qbNcR2GThIf5SiB60MKHZHMCxf8dPFgL4+fS
nw4uTb5e4TjKHcVL2+wBRysFwJfzUvT6wDfsmNu5/ULoXalsHDP24R4uo5BgBQ4O
Ufzzd2ugLnT2RnbkOpWaMTtP/eKlhr8cJy6Z18ZepHLoyBdq6ODGhLJpwVRwM7gr
Nm9PehT+GSXK8e1ASRYOwbtWWtJ2YIiwcFEKTj8z50l4Y+g7Ml9Q3sXZporL0Zfe
fa4D00iYDok2I2T+qIEFVC6jSbxqV6DCMe2nSjK2jlSwYlkFhuR9UA5e7J5E7rGD
ZiPblrxQCT4EPMmxfzA5bPtcvHhBeI6IPGFzMB17He9EMErMZaeQ3XecBBbpnKbf
8QJVQyJf6Udyg/vi+UbTsx8LGBQPQBFt7Dv4dFOxWeEf1udQbtLDmr27CAUpOgvg
GQl+sp95Sgs0RYT+Z83QrMG8Rh/7DTqxXP+ByOplFM1cjHhnclIidGu/3pjygGyG
1psX8c5yBqj7elvvJJABrtywA3f7erUKh/TBj/DbsEUPhdcYX7bd64da+9Qh193K
hwl/mg7OEm/jH2l69ouPGCcDf5Y2AScWd2z5oB8W7r9Vv9eElpGNXBeUQQKpP4yT
54rOYk98mtJNe9M3gzwEi6WssQPQsLraz9IlHPAzTJ1Z0DU7IZDjAVSgopW7RKDO
fJ7CHsYeqrI6MNvZg92JnyAc7Wh4VpJDAJDnYXNkaK0XJZplcMbxQZBhlE34qSVG
57U7enKLq+q+GiOVLJoP8E/Wxhhvqpy8eJadlCbZsnX9KXI+hwmCk7B/Z0sFU/mK
h4P4qUXVJts4hBAl5lOabIGdh0Vp40hDlwy3KxU010b8ibGw4yHZq2/q3IIkGJUk
YuLiF6R1lfeIc77vKOlvoTv0DyRpRzdJdR2eXZ1iNu23SP1qP5pR2ur91gCmGROs
E5xAUgjZlRv/bMu2+w7GBZC3nvQE6yO3mQPgwyNvz580SuhU5lSGFHT8eaL47HFn
JcVyDmLnWCEA+OmoTB+2Dinim5v+/vQGesktKefHBez0xJjIrMyatu07GsKu67fq
P+xgLi2hgN9C/+U3Msb/osNdwjeVfmXKaVChJErixu3rm14v0xlf2HaN4UYKDY7y
48wteoxbWNLZ1+k0JRXJYZdzAsIx3/azcMMW341alrQKVjWXVzwferxu5CLOkeeu
4hcxlMZlf0vQOs/A2P4RXDuTAdcn7p7togAAPBkHtKrQmyztO4Ul2Evfy+iYh4G6
dMyvFDTCeJ3jh0Y45Ty7fBZaVxXdurzfupdK9dmLeb4diX1wH3iDX5KJGXJ6uWgN
WEgtJLgBfkX4bmIuSXreW+c/3wwOEfIgqujAeSFp+GUA0Qd7hOgaAIh7yUUA8DVV
U3UstcjleJSq+tfizHIZfXQUCZr5taWcMGmTTIErRpy4K707nnjCK/FVE9Dtq5IE
xferVzNqMyscTEysiF/Arv2gBDW+bHUYlNQpVVQcTaTZ+xepnz+rpJunwAUS4RUz
lbOwsksqjnM03oDqL+eCrgFolb/fJmAtYOR5qZ4bLwjL5NdPD53cCYTJzd97D6rT
SNBEkG6FT2fkbWAJ5IcR7i3js4DAOJueO6coe9pm/ox3YxkTgwOjrZ5BLMfWNVYB
wPds05dGCXpbbCJFIk3C0OjgtgE6Cd/JORsKV9Ecq68m8qxi953zG4Aq/9u0kRji
WKAJQFqDkChlHW163j0MrcrnSaaWuhzVNxhDVjrLPKnLFnjjrRFipW1rxGhQG6cR
600JQoQMg7jLCLyp4j85MyIgEm7HKtwJ7l+ObGrkM6uifdkOolCe+CNEuFM89Bjy
uY4f8YxwpGoFQMWWfI5VCYBKEHX2h/gOPbBqycTVFOit5/uM5sRL0lbAk/RiR8zZ
c+t641ZDeRvkzD/6Q/7nRUzzB473ar5UydA3odtMyVusMZrvAGT+2GgEo+ga8UFV
Vj9rwrVc5l97RUk00BinHn0SMj8ITUsZ2v6scmBkExUOcSmb5Yv4PyUVvabRwW3K
28bddPGwoioBq/uoj6psywp3tMJqxBMdozNMOfLyEZaCIOsKaSrhoA9otJvrjWbA
n2OpEcSlooIEIt+3XV9JP4Tn6vhzL/PaX5eytTW2+RfYbrmHOcaLXEy6u3nJga3L
yIsLuWqe+cTgmMZf0DzCTCU3TrSUiwIdUy16lJDTLuOmBBrKLCPyKOTfUid4a5xm
e87PHHRRWT+RA9pSESTLUm4hBrJlEMVlicGoVeYiR98Cyn6baDhwXiiKIQyhyFzP
9ItMe6EbsGGtopBGtktDZMmk00jF0TdwrJuG6Kci92uNYhGqp/xpMxYR0bdnOdxt
dvMS2HbYh/aLl1LA0jV8Ckt9R0XPeCx651KJ0kYHXPgH77pMGwweNvo84+eY/w0O
YVkN2xp1dXDOuj+9KRqnYuLAeW5K3ZB25GjJ2u7HLeUOpbhRZOdyuEi76tDT0jc3
+vYKAFuSJaiUsHV1ALyslD0zMQoqiYxGLUChX9kWWYDnYdDck69MkAs41ZytI1CU
mmhjsSkrFZ3LGGKaWGMHXunC5XLAVDi1m7/ydZtJ6ZueahsnQsEr0aD0uzsmaGh8
v3LX7CsEcerseNlu9k5sUMICI/VIGH/GIDVctSvTF9je9AzJ70d/7zS+tm9Zl+Nk
UhxkS9JLCbi/KaGFB9XqlOCqfjUsxePWRlAWJwLxDTuCKaPQG/Au9VZM1maAKa3I
B0iuQwe6a45itCuA1ycl7Woqfme2Zm4jv/S8I8Ej8rMnSMXrl8HnUgKhIDD/TBmx
2q5mHKrce7GaENdhZKsSVkxtHCniHaO+l+3e0XnvP2DMFnBDRm/mTzs0Ixhg0RRZ
gBwag6eIAbUHJnx1MFeV3oUWHW9TMAGtBZCrHz96QNzRgsT6ikBp0buOiiX/8s07
P3+gCZGN7kQbfRZhkGviibB0ZH5wjgOs3C4EdPR2oy36Mo5pwVCXzF5lJLsigvEz
OrI1dob3c8o2txEVOhxrVRhbo22NoNPLZBBj0CpZKrrQIpLAJ25QwZKphtGykqTR
4O6rREQBYxJPz3B7gTRgqVjIcRV1RTEw/gb1yo5cIF7tkqznTOjMYYNNsr0MfULx
zG87hRXia26Nitmit3Nn4+QmZTi8TWo9DR5pbpiKV9OpcX5GyvEOAh7KU1ufaUKT
hbbosljR2QTL3BbQrGhUKfdeZsIbrJ1Dff3O8cukPkEBACpYFgYuuQPvlm+Znci2
PfeYGl+4SFGazMkbRi7bnc9+WdBEUHOytq7UFhaKPznO2nE2M6m4TFMYOGhyz4hW
iYHsOoskuf3adnrj+rB9NTAbpajk0LuFg9Pz1FmasUBslTEpxU6we8CO/JyRDGjb
O56FkJvqxNhqHAjGOrqi4q8fBvna9e9qNSBvECY8P6xxD3fiKraANa2/pKjmJwUT
rzS6Y5dkGERDKDlvcsVaeW+f8iKXyCc3OLsoBeMt4RLU6qlCzUTR+jb0462r8jlv
TyfjN3Jno/oKQeFwcEHO69P6rD2PxNpZBrsP+L0TIEVAbcjRM1mUV7mft2wZH0nj
x3l7ioysK7gqATGbwJPZXNsL0m/KM7M2TFYjb6NhP8qDTnJiw58mSBSeQGt0K1lc
mg+JTVXfnq47PLLiK+89rMuq5sktxoxGMfUXC0u+24F2htiKsKiteFeSODiJEQm4
fLAiWoAf/f+paDADheGaF9OA6HIN3C+n85PiOp1sArq2baZON61rZHnDE/Rx/0Iz
v+F10UQrzxFdTuRFHxJ7ZkPuMjUlgEsF7dMG4Zc4CG9Ofp33Mdkq4ZOcryvEz+Zj
35ZkxVTOtXFgCiSytKyyERg1O3L3Q/HxxeHML0Op0CHBAEc1chqc4PGnZ+Bv+ZWW
GhWcLzhHaACu2oNXd+Lnz3a2VUKLWGN0ziDQ74T9HuC+nVY+Cal4jf+wZAEV5rAi
mZnr2SEQS5g/hcLBBcyKcs+n/MdnHrFO4QWOBxGmyL5zEvDYdk4MjwfNuNziEuXN
qsHwc7YcGJixlBtqdsHGBGCQ/dxdcVV6V01LBJdUoVhm0iipp4JWVNXDJyoHrnXV
mMK8FoZSkb1J49iOEU6umtTM+/299vpSMOkTD3AfP7lkE6UJF2flzARui11ciHa8
8U8pe46983MIEW225TR4YozRwq0hgrVcd4+Pkp/s6VTHXvzC0R+KUthlVDIXW44g
mdBa60v6f9J5NRpj65E5EBaB5g4j/V4SInzYDFl0AawT3hgQqeaaixf4X49N83Ng
nKmER9F5OhxS2D9LGUkimT60pWI27Ko1CArAzUd5HrOzaIrkUjlXrqI/P+EifvnA
GroqrmNMpJK2bkfYpcQkyVu6thC/MNKimBarafDy8wVNWG4n0BjbgafzhpBVIfcW
uF2s5rhBmdKX1295QmgAQ1ivPePUUabLzwAjZiSW+YsD6jNOy6vBuHGEivwLxkW1
qGDGi8hzZPi2I5z3b7lewr+0hZd+oJa9y350dODAezeHlCXYgfdMRHl5oUCzQhY+
jZbmlbaP8vFM4+eTFyI49M91d3YnN1vG3Kktct7iMyNLYDmVxFXqrVfHsHzNvNub
ZJYPfVNSpOSGGHTVHP+YU8JksDKDfPZM4q4dqnXi2MTvELLhKR7e/nMWhB8qhANR
CWskpX6POslw7bivmMOun5u7BhIpup/L0cgjhS7seJ5rYXBl6171TwuRZmE7D+GS
g0b+e4v5ydaL4+hh8H1QVNy0N/moCNYWLnDCRgh3UlJZJAcCG21Wm5hUH7j8U5qs
yJG/hR/Y/Vwa838eLSJkqwlIT/XLu/z1NexeDsxuNFaO4nIvBEfwHLPzH4jo53Yj
wlC72M4opJZ3BdmgE05b1r/7daT7ZbxI2pxsaW5Euur7MlCSIVHszMG26BguYAaf
Qya65AQeoe7A+fQ5cYYvGx4CL6OelOkPiGgnGdurU006M3HTnLQzsfGCULx+E7Dh
ss/qa4SfQLgwCOSvM8j2d++b8GhcmVK9NKjp14nmnRFOZHO3MgRowzUN364bIzb5
cOo5zlyBOszmYUA0eE02wbx/GKULpvL763KlSIMNFhcvwTVMQkOq/D49VFKmHbOw
sW4YTlbe56viH8Sw9wu4z29P0eIbPABk+sHGhomnOQX9NvIM1JF3L7hW6gOYMbBt
cqTYyg6mK3S7GPchrt5LpyP5FSHFJsBacEWeiwP4PMW5q5EhJvUtZtV0oc/RIfsz
xPW75jMpViMbHgYj7/u/StECPyjhVt/HItCnujpxhbhsAWu56+ka0+ZTGWtO3NPn
jWIYY0KYdoRi52qr8/OadH3qU0QVo24ja+VFPTa7SklXcARyHMlCVtr0jsSj5dGs
UQ5Lb1wsQ+cbm+hxIsUPosIjDCofAI6df2SpV5sfN6VeFBsiQKwgb1a+S7rRmmsh
RByl7Px9JpfSfeUqOY6zudriTUbRF6SgPCBR8VwkowyvMcPx31JRcJ5cpLpKcen5
zCjwqCL3P12vpI/eXjQHJrC0u0xiDxBBC4tUNi23j6V/kizvG/6XElr6D2Nd3CwF
i/ryusBz8Gxtm3kz67k+q9Bx5Dt6Dr2YEzAZLVPvpxFFSrmlC7mcXAVeIXRKvW5H
uOO7kZJ5SiZlRdT1xQkJVK6m7D8oZvG6O6Id0OQviDwrmQqqZjYKhQqxlTc8v6xc
0tmv6/aeBGSxXHO8xx1BT7fmCqiUBUbf2r5Av9gwpxOI8z7jiNI9VwY+RCvia7Ms
ovJVwa1JXJnoBFxugP22mlEl5/8s6J0ea8CKQGYzHJlgkOz2/Y6z9frx+YC5jdVf
xLS2xjTTnXiR/wCivElJphdV/1hqgaI6NTwZbI6gs85lrFR58RTV+lKis8Jjaccr
K5sd5q/B5oR7dFSeVBsquDY9roGdQQEtrraNFJcIUjSE6h18cZXpFHeEUTfmCs2+
92W2XP13oF096f7OHs7wdqCsJPmk1b8OhGpeYGF4C+dILLqRVH86XrKgpFYgytYQ
k8KDmqe3vj40QdpNoYpmb5uP+lI0+ia6MUxX30Snp68mCJzOG5BHJs7jcO5LpLe0
on7pmfwAaHEgtJJD6/FMon6PubfEyJJxwTZzDJXUlgyiHZHbgyaKu4K30oCdEwnx
56DefH4BIDTV52q+YlZbXCii8VvcZAHWcjd1USJRj7hsFLH3nSD4TECJzDh31IAN
JtCcnLs8RwB73rnIbD+dNCno40MLsOUXsxTGjP0Iqtx4KUCb8k2u86jo5JzH9iNI
JW2CGquA+wAkZyAhSPLCfiJVAnlw0ZTPsYoRFF8RRZnSMrNygDHTwGhlUZmNzovf
a5B1nDO1m8KVTSMjtMHxb3w6/4QLr48jUdtlS0ULb2OnqJAQrOE7Ieen5a0cu90c
j+3MrWWN4zDw2Uc7oteZkTMZLW/c2GgCwzc+ZqoutOfditMhnHS8xUwgZzXrvfn8
ZosxRVflU0+FVRFni3PZILueenDMUqa8Dl/qkEbgeLVnAl4UnzM+9qh+pyNASR+c
kxD6kHmYSat6pyS624OBtA+CH7RNaDetX6e1Kzj45NA0Qp+N/nLH9/PSLCgy/4q5
uEs4VgDpO4NR8QQDIybyx2J6eBl3crHnAzCeaB4Kc5u8VSYHpOCo+3ae8KGB6F4/
URyaMuNgHfYmJP1P9DUACPr4eQG9lYKMcma9g0PjEOGVIBsGdKLSHbbWBYkBFMGV
+e++tvQJSg6SVsq0Oo1fSvn60H4WSp5Tb2cPHYinoSZjOqKD5qT54S21Kyxv+ovC
GF2j0cgN96JLcxB3x9RoeIGkLXPNm+SgKqKLHAHvArEIWuBYk7a+lNKgzNGhsZ/O
X3sI6pyc3NQVsgWzMqefJXJ0M60vv0VeTeBBxFo95nF8SiZIvLjBSnUg9mtv2em+
dyLQnTECQv+wCAUBKXLOddXN97U8IaH968Bsa5OQg1asHMsb7t+3m+wvEDs6IR5g
/QIa70SnxDqxxXxXnCrHJZInCxLina10fswUGowdT8u3U2CPJnelc6LQ+lBiWyI+
d5PPMUWTT03YPClPIkAgaweT1p3j/OQD0VxOIUMP/Qs1y1+4hzFmIX9kpBRc7iZG
xRYTv+peyJTkxjxBxgvY03o35xxIpT95g+hrnWLHxuw04PYCduyuJrUled3jFsM/
C5p/1SalVj25dG15nqnSa/VB/6Z9LnoQwkxi/vBBuzm0NvpFqZLE9abUwjJc/bNP
aeMbqhriuM1z4qau7sfA6i/nRgSgAozXosL5WK4irSHIIBXVjkZJQf+gPpHXl6M7
vOqANWD1zUlnN+kzyw7DGpXUuubzUDLxrO12i6U3wBUPRJodXQJxS8eBwKUgn+a9
no1jIcjiYP+GeOcj8a6WFdlkGgHcb9+n5D6TY+850ZHqMRxyuvaRzPrRQRcVrbvg
9mbskmXw2sTccLwtyh9fTsUVhRfoSMP2EB4cUUSzah3EIGoamSM1uM4Hyi8XaFh9
2rloLQVlE7GaQ6snv4fJ8tnD09P/DYh14ZqhYmmsbEeotq5Un0qucbPyanVrroms
H0IKHzzsZ2mIWqi+OUL+XIAcglidrkCIWSlbLcPwVr3Qk0LPHaY1sQ30xgw1ssWC
XNu+pBYufncRJeoTffqGk2g/RIOBwLpGYKHA5WPZZufH2o1xazfzBRTKnbtYKEva
1eAeGMZzIysYr6N3MrvtMVV7kusRVXmO3rvgYmQsLIJyZMhlHkfnfB4mzzIVhtTA
Hf01raukB7lc8o8qOeRDCcSACP8y7dSiBS3/hH5HB75Mwt2YP0eFdV3R14qlUhqD
LV1YEF0OfnfFro70f/n/MQTlqHN/ij7q/smMp2OfoFpudbYocqAuM0r4gsBZq9Hf
S/eGf979eYGNJNAduGBYBrzshUWiQsfGkZWWnCOWA0cj/mH1R1PsWcM7DZR/E8Vk
xkVimVBAcZZrkD6zpmTfG/COMf/e7aiEAM9Fst0mzzuds2OzngFe8d46+soOBV2L
NwgJWEG8d21/n7lIflg84xTKz9bAQgaX2gJAFd928FT7uyu+k7V3N2AcXuquJS51
am6wbWq3RjAWbWO8hD4v5IkORewbmsv8rG2UZroLz2XYOBgACNdSK3z1QImmTUKR
H4Ub27wg8c6sucKsYP1ae2jPU4OfYt8nFSoZf7Kf/YmnYMN1FGdRY82vU3vScD0g
kPhGmPHPR4FF1qJB2Anr9VEXW/rvdRFsf3ASCgHZ704PE83rnSugXbylC8bhImJP
bJ5LjEQ0K7OPS+xazAS012i2jpRwBFLQ8bT2RBoCF/2RT6y6ENM3Ym8TE63G4ZbD
V46CJ23Bl9VAhhbXf92E54Ap6TDAtSPWOwYPpNLOwdVp4k6IB7bjPUa3U5xBeie3
ahC0zHdfJXGobjUguVp8VNXIc1qx9Ly9Zr7R6lp1DwaCoJRmuTRDSXbOuAiuKlPF
szn/6ZIZqgYExso5kcmB4pV9Vsw6MVmbKwjD6HKlVBiPs+QggBTetJ5nBRPFFaxV
zAzdnAS3pwhwyIoj72JjcFMhzaFTcax1SfrWcYWLuSkgtQ9kSGuQaMekmPod5xcL
TlI5VlpNusUZv8I+YRseX9KrEmYJUe3ZlMueSfsG8OGaXjm1GWkpRlHqA5RSZU5Q
J16PxgNS907VGGszBEzQLmIqODaA2oVcdVJYIoovDCk2QuO7WLW5fHFm7wy7dkLG
eeTPcPjU8yFAlaCLqYb270BYTxMSfZQrd7l4bsxJN9xUd80uPlQ6VeHiMG9Bx9q9
FOooSgzCC/93vHQ/e3n9MoqBksvePe98JG5kbdUIG6cvlio+R0Pox1WOlf8UD4Dt
fzJQv1wx+fXViinzYeFvW2JWcXPeV+edH6lAgTuRTIehA9MThFNx9Z3fNenZsEUW
/DbFWPGnQTyBceu+sOwwRjwDYVl4Zwc2nQZZzucpsty1HW9BRa8H/omaqGyIKayI
UOJpjMicAsDy5ivksfAOxQ==
`pragma protect end_protected
