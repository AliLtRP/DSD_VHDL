// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FezjPvJXW4Lpa3yBHriiKomIrIz/dX1nJaa2fFRu+5WhAfdi/HATex8Hue5UWTTA
5q8vHE+um4l82vsPA4v+cZQx7GxEgrew0zFip2MlSmUWoSXQ4oQ2IfzGNzNs9K0q
NtTTcst1mJlvFwx8hEYt5zOGOMVtqtUUjSFud6fyIAE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24688)
C+BEStKKawNJgJtBkjOUvf9kRKu1w91NnFbxix904D89s0r9LGBAJ2TtCBsbad2w
Lh0VsmVsbeIA4Lx0Och9nX3/nCVvfQ7c18bPqdhSzk1xFMib/bByRWVi+8eAtz+Y
UiC/fAvT4zyKsfppQouwom/cU2YLXZ0XP5TBHGkSvEsua8Yd72iYAatTnxVM+3j2
52v5EPZOAOEtWh4tfm7hDzO4tMwh7vj3lRKTEIGh+XJYvLVWlTFjcCD1Pv+QBYeO
B098Bs/v0BsmsOA7fDClaPMn2z0Q2KaEbktTmfK6TtlD1PhKdCUGdtDNDas32dO7
cSlLQ9WsGbGHxoJgVEQhuVxXIKWDU2anXpWBzPVGhMffXs0dGr470IDOZpH6pOc8
efNcWJ4bYK2BPtRsMSwvHX5GiiE4zzOnOCpOwoydYdBLhGxecVrKaFzTT6aqWIcs
nzKg6oKOZYnlFOnY78OcdJS7GueD5aWe9YhCCe07axAIdKrMpyoDnhMgiD6WVXGQ
m1cKDRQsQ+Zz5iasu3WXw5FsBfk0KS+vJ8DIs0hBU2ux7j/eAdTYZ+qsVBAhHr/J
Nw4iohQyU3f90B0KayFkV8VVmU3xk/7GbJ+jukis9mlrCK/YK9tzZEmq/i+rAvbw
pADnmlaimFgdlFFgONDcsWMbuNSn6/ZjQJODAtkj/dLb8mLZf7O9XiPTei5WK7dz
VzNpaRl5ZayNoXur7g0VwtMG9aMwvi7GvwfL8ZY2JUXYuFae9nKY1Zcyl7Kzf5xO
IE1R+9NM8KIgdMjNMW5LFxfZbiR4e6fqcnmUZzbyzXxBx/ZtgK3qhIX7CHYbOGaf
cTPE0c3jD1uknW5kD9+zTYIMMUrArjsO6Yyf8wQVMFTw1de4MhvEJA6n3ubKbEHh
X/D/af1UBB/JyriDPY1GoaA7dF1V44SnRa+hFcYFWitscWLTAjc20d1uW2xKlCEt
+FbTIxZIyBO9BR5pCibsnq5SBQ39h6LZBeV0xmv1SE5mJ3H0c6+TWz7PKkrPQ6bg
WX6S0n298thOzL1OMHKQpPeym4UKueXjK3y6Rw5oghc3k1hQOGn5dscKo25Lz4Lo
5SK026n7B/klhjcRX7FsPGP5yb3OXVJ980o1bV/nGp+qWM2OHSI/YdwX6tzJ7GI7
MG9juJ5wlqBYsDe4B0npHdJpoHslpRfFup1v9D8CCIEN3juJVnCAIKN407WN46jU
LP1WR7Om1ollemkAmK9IdhcajwCav1CfkJygMzZedi6hzgcDZY3HmE+ISRiImY/b
XHTic31VnWG/BQ6y8qM4QSuBugYQu0+Z2Y1w14+8rngvFxwC/VirugUThujz37v2
epHqSdf3io9TXjZDvyo0HISah0npUPrLT52/XerQbiHV5Yiz0nYWxZ0PF0Ts1nW+
YmXHvUkwWcjdoQ1EK134fqXtp7/Y1pZUfs9RzedCk6LNr43YaIA/6R1SCMe9H/I4
T9qhgPl6sqMpmYKFFQTBCJw94WW/DXmwacauuxW+9cJ7o9Fn7HkLM1BFS8nOTQnq
yW6beVvhr6/KO97nG0NhdVFAT+RiTT4mF61D/9e6spalcP3ASfJ84UoxvtCEszuN
fe5YFqfId2VSncJMty9PL5clfJOGUQPkvYtPhmwsa33GQKe6cJbnqlQLib0FHO4p
KIDFXY9kNfGNdDPU/jBtF9bCq0yaKEA6JsyEFQelMogJ7ECxkqsSy8ePwkB7Aftc
OxaaFQ/Q0e6buSykIPHnFwQpT//nbjzOVvRLdn/yBmcDLXerjcl8Ii5lidPHLAJE
o90hw/+K3+iOfaQZtu4VhwVg9B73oyQYW0JMQTYCXHIiJRwTvFBItvcT9Yj6eTjN
HnfpDe8jMIW6V0shVftVkT+rKamyba86oOnBgN7BZy/yEDf3G2kQa97vtghD236f
MQceAlwsDwOi/vuW8PUs5YPFPnxC2YNv9JPy68QjBfeR7F/rSO8IsEP6sWzg3HJC
cggs5Kd1k159lyd5WfGGIF5wOAyaTY02yk+R1xZTJwa4ORuf5HMOnVnXm5fqhoqk
N6HnA/aL98M/hihFbOmDMUA97GYR3PdHvBMA1fY1RwYJMLD2M21nzHpOrY29ELwS
qFoJvi2kL7LQEbUNf6bdia7bffvgMjGJKyijFVJd44Tj+cw8byUNq0YMnJltgK7x
9Ox/CkO/TGjdDTn0gXA0BH+lJ1MSDOyawoez9J5dSkk3KBUbFosNsIK23MCvnxUM
jauL+387Omgv5p7/Bnzw/TbdnX7IsLzsre1JLXgiiD+inZzzxrlFYQU780CCrKw+
+99UZ6hS6AHbdQ/vTeS/F2FUVxS+zy8+a9XQ73B4mLk9RDsqGj4Aw9ftwYBIwe20
wBJEcB3ok63CIqGyx+Y6EirOcLrkXxhjsE+v5wW1UG46GHR6pX9FsWYCbpp+NCb3
ezDwnQ+5evSpOo/6v8nXJwdzOQyCkIyt9D5LmOzZ6SUD28wy+0BiZLDeVD8/eHLl
aF1f4a8OwvQwfjIvTXnmz730cDRfIpJhcir3obTlYDet8djaoE97t1llPfsuIOhm
Yq66TLqPYvfQEdI6c8clrHktbZmC6hXvaigjl8c7jBfsNMmhrCFPe3QPXLAnOMv8
+L/muZZZylQdExN0HCGJgdS/AqB+M4FZT7eFPDrJejmrVlCzUP86bmAQFDq5yg5p
X7O2hrm9bsfU7txfq00S6xHVoBA0Y75G038vB4WIdC1Jp+OwTvsqLe+GLL3fGzu+
HS2VYyQt+j1K5Mz7DQ8+4BU/dfSt5j1X9P9JmWnI4DHUw16v0XeWpur42gMBVaS2
hSQU5vvsadETepbV0JNytIS/x3gGoD6iOSQUxHRkK8dkVhx8kQHCsgVMaG8C9YBu
msEke5p+qBLR7DrE7OfcLMM3oz5TpZOmXfnRER/HnsBtVyCRNsWr7TyCbh+M4Uo3
NzoGT5wbY+8Hh3rUuXHh9HGdd7ThNqi4kpsR0aZJzYGS4jBMgxgLQl9xJLJUZPpb
MsXwBsS924r/PViOKpftoN7zTkQg11y3ma8pSj5eNm4X4HNBGzCmUb/0QNdWciD4
uxLvEbGb8fngYWrcNXs7vpKFP5akDi6vKa/rIVjpPGTuvspSRFe8cZVif11vD0MB
56DOm89LRXQHiCuZvUQLGfyT3E14emGPSw2Hcl7Gz/hKRJCTOKEJNgR4ODioXdNH
2+QASyD1PNKG4gU81V2ikOUZAQYK2xON1S/KNkbOIBTRpOpFQYOSrkgbq2TC+uXS
c3SiOJdxo6DjCPEiJhuHcl4fKZGtW3dIoJ7+HbaOQs3FxeKpJ88ecOQQIAwdi/44
rEsqW/p24z4wPCrihTAvK7UdITJSz1fPR1FZ/PdFKKfVwpDJG7CtZcUhOcgbljeE
sNSpGSVs5UjKUNWaIrt+vUnkdUZ9K+rXjiOmX6u+zg2AYODZCXXZmdBK4yEWdQZe
ToEl5lwfUzjrRM6HNaa1bV1eDRVQ4esD5WMF9GuLzOYwbwjJiH/cNe8IDP3492z9
uyOCEuhfhvArPiCqrWl0RwPiooxb6vdU8bWnrpoNG4OBfYvyxvWpS+Ynsyc3v0w7
3gGDhB3K8RmhP8xytKhfgwNPxiLIwoeZIvR/2K1+BcLTz8XKGsbsvpA4ndtdVOh1
km5AGG0UuDwYF8AKh41/4W87AlTrW8Gs5NcnoNbMs3P2evPHrA+3sKAiWvmZGP6D
1jbbFOIVJV1SaFlGAIB5KfAg0PUUHwQQQAHbcj+fgMGHCRLKmxjrAnnhg0Al+jHN
gE5tAVjFpx1dEbFXwPpVRbqfHu6PRIWfizDax1meeefi0LIZwIxaJr594Y10AW9G
nbzM4fric/nE2FYWi0hM02an5xtLaCRrKrbqc///Gxb6WLwRdc53UaDHk59TCgrT
Tafj+Isk3KbLuPRZTflH+NlfiZkZ32Fmj69FyUwGPJ9VqPecokHyoCsnZtaLxwVe
TBloFNv+40Zvb8RwExnWCglunMsB4dvf/zZeqeC4e73PiMPNJ3bP+iWZWEh9sATU
en+eBN8YWKKQpD9qPx/U6XJL2Mz71MuHIwu/iWo1d8fkVKqryoeJwWxwu/llgA4r
Gd6GGVOiS7etSTF5me5n36VNL4CE81LT5Gz1osBJB0oRikqNm4/BCggc1DlFEP46
LtqFcNXjGhkEDWt7916+Js9pyoViDeOBnfxv8+yxlT47uaXHObdSaM450OxN9qtf
06yYLDdx7tKT0v3+OSo2wWxxOk9hoabXoy239MBfGAHHTe5J/cePSDlX1nnzrv28
I5ti4sckszxe0dHR7BwGcRo28oXrU5+64cjTFIfa9R3+nHHdT+apHCTlqUKsy1vU
zC+q4CHXCOWZVrHoeDJeTBD2DFuJx+k5MOXOoT7QhxBqGNs3JB5zCTXK8qwcc6+d
LZYoMQVGY4HZNmQwUjKxxPfeB1Mx7cDiHzJce1uI8nUhFzVtEdc2mglugtDWhFv8
vP1O8Pp9ldUKP4ozHfyTFFIvnpm0T4PyiR1zMTLw1yFib7iPmZDtD2DOXcEi+7HU
cFHufW6y97K8+xET87vbbTcSx+RPZ1Ks7mvvFvLvEozY7qlHd4MJTHqClKsjCweP
0xx2u4cHHIeGpIVcFVAe12r+6WXwZzdvccO8DzOnonsBqG5or63J8e98qsBpWCyV
97jRhO/LY1P8boXkOJbMlM47HSTOeAzKR7fGytV/9SzA1n7IenDHJNK4kPQO2BQ1
kLEwQvTPXNBJZMPDM9yApitALoUenbTcP3ql6itgqbIRrWhyI7J3eTKWu4qxFfs/
eZ7VadHI10YA5vD1JBrgy9u9xOIN+p5twmQcsBgmAP9uViEA6oY3sOYYOp4mbMXU
fUiUnGjrgxpf6P+IQD6jNBVXkcvTNUhI02CAiowcyt2WGM+LmzNWWLURhKHL7X93
dtcCIxFWiM+l96WlTxEnt5jGIS4CYjCT5JBKm/AmFuiz5jwSsw1y4WdIsFEzI9uJ
oDzgGuH4t6YlN5TQo9fGjH+8MTX/PnDP9JHyBe1GkcF/0C/GJzEFW0bA7Qmv6n1P
nkX+69I1/PbdqeBsSQChNzbfmvk7GcRrM7CWT6aS10nH0eE9FLNDq9LL0Cv7cop3
6xLz9UvkrcsabKO/ZgxzDDAeqKGAE08ZbGHV0VN7mqHP4EnvxgGUk+jzGQaQDnfO
m+i8lmot8TZvik3dKncuBNyOvEgNx9jeAzG0argV/PNyyiJM9XuhiqTg+jWJ4hLt
oZ+TJf3+i1l7Xavpr/lbkRxRwSUbkqFtvTrO65zYE486n+XSyEa1dnZA/ybr1XVt
5w/I21DokkyK2VBdpEEKGHgq3KIW9pfPSr+5kZ6t2NIuqta/E62OhtVNG2TvOOXr
VQXvJrmsOoDlujBG8VRR4zrqAXhZjX9eDo0QjlNAMiCpF/JjghzojURSbv6sAuMa
3j2KQFtT+NgMcdiQas6GieUATt1PMBGw/b/dTKZDT+0QN7j7Ry/UIRSdkn3XTiOC
cYKlsWxOZpKJjAGNKVjD773pTBBsUpHMwiELUxQSKfUbXXUjU5FkIXL71Fs0YGhV
/f9GtzcFm72+36+INmlcFQ5uZkSnqrvILj3Mz/d//iQ0PtUZgD/jFbY1u9NEbC5D
lciRkuqLCmqUiwm8kajQ1oVQb3hvk6fHFx+jY7y07vcFE7PERi705crDJJ8AcptA
BkICawDObfKSFhLRB5LWJfWCCd1xnsJ1dcdQjjWnkgZzgu/W/VxPKXusIXrMopB1
lZjzctknK4kLqjvGvZOLoEyV1+I8caWfn0jhq3QylcgZZDqJQfTqfwsn9GaDLTtF
WgKKgyfLMxZRz8HWwaUuMaXOTcDbXJuAgi96Y6lsCAAhe6IFTOdI2jlTrgJKYhtf
ZeTnQZX8vlgSlRamjHYJBR4T06Yr1ZPA8tKUFt0s368Lc4iDwc07Qpz39d2BWSmJ
s5nYGWW2MClsmnTggsWQ2j9e2RRG/Q5vQeroyW4iaHcoHbnBnZ2py2sfnOCpW8lI
1HOphX0QsTW0NTXGQsxl2puqG3dN3LIUvv1zAUfXMRlXTgAAa/KljVLqMCmOIhbe
NGvyLteVN4d+y9W4wLAeayC6Mxl7K9pQwE4Qg75Dze8qIF7CMlEubCYnGlefKBA1
+2gAtA9AeyQDmLIIC0MXZugnUbei7mFUW59eE7mtQSu/dP4Jp+mbcUCZbK6/vWOx
PyOncn2OIKUVvXGkQsWgolGviATj8+y2ExxqYdbic+JkTjRZc2w8zWwTvKDuKt9E
Bwxks8RktY09rwOfiQfCTokTaBO1aNxaXyls7K9jnu1t8BjuOV1JdyThPrfs0B3O
1+vITtEyUJVa5OQ1OFl37otPXeOFS0mWn/7uSELTlxuGxuVl/kIoTf0kiKq520pb
tBTRUkoSrVNOtCTAI/w+3D2B3/I4N9Eh7coT8nz7WS3PMQkruAl4hIDq0XlEUvIG
MoYCBCtrpSFrVI6oqQQHFuxZXecyFxEQmvcYDdQI8MTu6HJXAUtL5fnTlGX5MYIk
qorOGzJe327paCi00a+028GqLF7IDicUYGL+RZqdL2R3c6h4g6EbgjljafPZL9uS
kkS6Exqn3+6V3cmfqJhlUOUW4pKy59c4jP7CrdUGJB7VQvBBm/3ijEDC2pT2ccf/
oU/tCEBP3ZXZb3S1sTdQVj40p1CFFqLLgdUJxfGcpRHb4WBU4ywZk/ZQvg03tcTa
kzQStOTjZdT/rXQX9++0OjfvK+JVCULBFmFYUHjTEwVtzSWpJtBcC3rt8cx5+yeM
3Cfh5tDzeBgKHTpzWEhOWn1iMTi9Gf6r+YCRVlBRN7borrxtN1BRsoKwPYZEXh3q
nmue1GXrs0kn/7R7wUeJabt0WRKbzUgHp5WoAoHeLnnE5r2vDVOT6IeLEwQCfSoL
SU7sk/aZg4USO8noFpBOSTM5FzuU7CWvBsJZt+hzLzICACkeuWVBlBeFNL+wkoNg
q0v9UP00P1zajHlk7aj6jVP1VVK9QqFeSBAnRV3kLwl3Ikk7USxPFkmtS6KIqGq/
RhuExHOqPRiqTlRHUBiJw78k2ZrTOzbIDoHmUmOIA3HGTjLNsMAIoqlyIQuhVuJ7
83yWw946ZojoZbhylF/rzalYRp2jUGnpLaLosnaJ4dyLlJBO/FVeHIrxa2BZJd9y
oQviQUVk4Vxm/V8DQBdAW+7SyMZar82ELi01k1KMo2ED65EoBpDhVJu61hRrVRU6
AlxuUxdIYRc1qRJiMtKwVKDdybnCCiyiNrXnQzufeWiE8AiTu+advvMm18X9xwVQ
3HVN/9oQc2z1bzg7HOaqtsZJYRpMN9YgiSJNWNBp/dKAilRTELGT3ppeusLwe+r8
XMw2yJt+X/NgAY6kGNLHpbIhsvSY7kQOG7auHK7zn4PccuViLr8Tje6s8LQJNVht
JqErB0DhLgnz+tR4n0+EES7mHcyyVGwTcdP/8mq2Z3HAj2B34MIk4zZqomY6dipo
fbwmwtEtC3FdNpZLFpuujy7Ys/YAXzY3R0lYjHE49V+HV/BWzrvCkR0WGejAyNAR
Av/cob/ZPxVsS2KTZZMpKk2MXWQd9MxPG+zKN0ZMGLa0vs/+E3Je3Sk37sM5vEes
7WUnTQUWXV51V8CGRLOtTuD6/Z4iIpBq/hl49D8TuCI6ioAYF7yg7ph70pbsL+fn
zV6/OgYEH5l+Vdsg+V2T6OE1DDEP89aDxxFcChl48yLKvCsTdjUGQi/TCfMRmJMy
RJ9DZhOd/1VOgHwF1Sr7BD95yTYIpuujcJipvm+iI+7tNO8et0GsZX4/OF7E1FfS
/AnSKXnflxJxyzPyh2HTM8/Bzaxwy4q4C9vpTAr/iHz+4JoCof1WLgexRHaxXfmQ
VhmvZosYx06jBAcONC5F2gbFfIqZoqoVCZDMM0pO5R2wtZN/0ehu8E+xaN45ix0b
GieyE7ZGBzykQc8PE8sAkg53Zfy52goLrNNj6d8+mH/F455bjX/l6wuRo159hL9V
kmc24PmxgzKpsFxRJB0cuyI3BaORTKGrNpyYIjICBYAgI11wkPztXFX8eVvp0xVD
eZBsEkcG9JIF8Kd9tzCM1D3jDf69DfKLTzCYS8YgicskeEMER0i68qcjTN+9XCZ/
jweMfJUfJEjnHvYvUsa1lRQWHpgRhD7OrGq+9o5soL6n2XWbUQJAUZOp9pzIdDSG
kBG0JlpPlVI/jTuUHeFziYS9RbI1kTwiFenjclO8Qc806tdb163SdkNqmO/b4Yzw
283usv3TO/j/PGTlBFMPgrMu750XXrG21JEMRakqJmlY2ODveYbO9KiXDY/JFj7m
ZlQd3yuBv136CKeyuavdAaieg7EEz/Ltx8mfS9fQ3HzO6VgchajAu0MtJ1nfV2+i
Z32u5EWhUgegYpw9R4aHIIEYhPSsZO1cK2T9/jAGg8EXFKZeCz37OeT/4nmvOcu2
iCdJp57UZbm1cL75ABgpgwY3YgNr+hKnstXZp0ZVRJfmJiTpKdBjYcVnpptqbpoq
ov/3jxq8UbSZWTe56DM84amTEohIQ+6KtSYkzHze3hS1KLkjfTiRBGcmAQi1J56Q
gLmSy/zUfvRS60C+3CYWodCQQR3yRW+ggLUDzP2rT1/K4sBCepzIaqKyKjEh0wau
dHbktJ0o+hJS7Q4Wsr/WoNv/7SOXI04C82mgri4Q8U52Bjm+Egrpsoe1h9HwAgc8
XKl6Qr5VHrp5ajPnIcThP7gdr9KeDtZTNmPxoC2q2kfjEQ6Yu0s17g0HjZwkk0SV
iM48nbKSAlhyoRa45zlHZ9swJev5QoNRGZAwfwQjsYw4WJY1+Q5wIlbEQ9Ila03H
JfJlmvaKD2QPl7xiREsgo9ZjW3qRoI4yDtd7RB2zkd6iczdOVEEMaa7YjHU359NG
bY/37ruvMU3o/SQwI55A9i5FLxdtuRDTaU1cLOj9FSacqHl0qR2bpbzo9afTRR+Q
isP+S7c/oCq22Qi4shtZBMqdNPOKfooaSx01bnaY6omZzsF21Q85mPH88FvE+oG4
LBqoKIjnHNUyVI07fyrOl5SMCXKGdKPXTOQeP/J5XTxdze9pX/3jZ/24tAmGZIrr
v1690vF/xj4qYcgh/Qsg8BMFFiwWGDfi0VMDsOONSEkI13NhUqIa+NA5R0kkCvS2
sZcKQVm/olcaA8D6upgp5pOkDTBeOOQmQrDNWgGkUzWL5pzp7maNtupAxSqThyop
lbkphN9tC+NBVhJrfl+rY6IeIREaKW2To+ASa31z/cO9z3AdHC+5WI39YtKvsMxV
RzrWEklt8PWSFDPfWJOppBKgQ7WuOmSb9ZzgM9NrHYVcR5Kkq+Gv64P/KbVcJFJa
SDyR1VHDH0uIVDRSRwvY4isuqWGqwQjnjeYBIuhMaJG5IEpD1XJUf2MFYCDIi51s
qY1NnyEaJkFEUOmqktd41KIonMmQW1C5oRxZsklF8SseNMit1MhPpMrCa5FfAGTN
SNAXCU48VLi7kKMJ0j+EmT0LYbu4mVtwJb2Kay/WMRHhIg4BRy6o7D6n85l5txyz
5rHIrGn0O39xbdNZuQIx9rSRE5ltqZxQ3O3BLt+X/bFSsFx6gNQsaDRDrrGPZlF8
DKNiH2aFhehtmqKW6doIebM0ITWFmp9Y3BPAqAmt9YVR/zOLxkFK6F0EyNjCdggh
UVFCebPwRtlzSQ5Rit23tM25HRZV79LThosE7kO72l6b3dcbGorpvl/g7ab8Xfr4
tULE2+RYg1AGb2bZdWVMDxWC1MKdBSIgQkIu5uLmnt4Nt0tKhlXMV+jkcVgts+le
o/DjM2hncGOJs4Iik5/ZtIApDcCHBKkVNmq2rJbUEdZXMNSqWbz3kXBCjh7lUUYS
HLfrecbtY7q2MEbT/5QCm4DCzbANovj7PjUHaRjz26yiBSGSPouACVXskYpxuEGF
5LFnKzyBPM9xT1nU9GJv+QA9QiWPON8/GF6C8moSd2byA2JpLrzQho8A7zvyu2IZ
H6goFQrnMWTItEiZdYJezuPECTtrcFKCgXaTv0yTk77OpbLRvHSZkH62j6Bpvrba
uFxdUCfaLNSYw5850erAn60fjPzmiJPEOKpTc5BNi/ZBl+MxWA2xjMkwBIK313Q1
lMPj95FBl2du/ksC+thKLdaCLzRznbe8lF5s83TzOVtiuoe/o3ZkNSPStzVciddt
mRVoNEcYfK63GXZWWONIMu+p+FoiuTbGe3nKnwlDAlqbCJHraCMpn5CGgKJNxv7a
CGEFvVuAI/0LME8sxdjQcPrBAMN6zqMRR+YQTxbGI5FMThYOXC5EjP6kU1ZjRMTH
YE3z1NWUnGrCj9dpeMEfH+JoTU5cO6EscUpBP3qw/wFRT9x8RkMdZHTBsvKLXsm2
W8F9bnv4QUcnh3iVIuSIQJldWR6pker9QUcirf5zihmaRL4+9m6KYl+yyU7hlyon
lOapcHputH5J6vSL1OA1erZhWTuhoBwo4zsOCQZjLBSYJ8ABm1qgn0nDPI45ZsSp
jBVvggH7BAW2KDx3ouNYfPYhmIqF+AIqJKIQycdTu8zOyav0inrg9ADf8gC257gN
PJEqWo+J0kQX8WfQsP+8cg0jIePeMf1kO5S7osreXJvDmuRLs+7b6ykCXp6a7dbm
m9yczTK/XBwHr74StXzvvd9O2z+LB8iLDGBKZG+dN8mGi36Izd9uleKM6RT4jvOt
3f3C/kcDa6jOe+BfU3sVJuOSeqFOsZRE/KB8M7SbVMjV2Fu1rBWHT4EzNoQhD6U+
dEfuFnYpgJyIOhSckB+0D65Pjo/jX6YOwdOSaLeq5kxWSggz7dz9i2eN8U53EL8R
ZaePoqe+4mLXFacZ5SpFVZlEO+TduM+4LFDHYC3eEnhDlSSaRTp5+J0Kkrp2ptrf
3yFNPtJmcxwmATvJhiOvLI/NdMYb452+9Za5QMr1i2mHT6QCFDyOMgHyOaeCYPoS
wFDeJYUP/nxH3z14G6JJPAteZfWmOAz+QNOUywTXcOXnlBC7A1aY76zsjjA43uJ3
9fCwGbIhUO5D2MFsQEzMlAihJlLZ0BSH80Y+LXysrVUOopW5GAGX7PFvL8igV97t
B6sV1zR5VMgweKonIgWLF8n0eFSCb95KX+0mb1mBv85GctyL5xB48RH/zWefqXUU
ZUbLdO7jJoX80YkojFYw99bsVdmDoyap9cUmJAHdNSJG0yth3n/iby4R1K3Mm+8V
9Lqbiq8hUE2PeTO7Eb8DW7YlFaI/JfVTxg9KoCPgdH5uasqpbxCL7ln8qeO/toKK
z+rDATrQHuV0M+UwmdLAg7CYQjJbV80qwBhXqQxivdjq24QpgzZlLz1cHGoUKO3f
frixgVtIES8eOQkI5ftYC+BFYCShmESdBE/zfkv0MDAxeopTn9eOxViPjwktrZm0
cVAgD9+ddExCRkRF1FUL7IxM9jSsPBaAjJtMLOVb5y/Brt5NBmKwvvsfM40N1YMN
w/R9Be2KCrd1ET0wDUxY0Qo1EG7r1hodfDHQUAG6dzZHUBP9LNkHLNeuNgsD0VxE
MA2uwHIl4dLVwStuDGOEmFeZ6vsrqxHj1zbVElbT8xN7VK431FHgJ5cmrDW5ZgCw
gOruCr8LJfLdhP/bOgecBharUtkLxYdCUqf1o29Vy0/6i8xUiCVYOJxrTsQKiL7R
8MO28wJcX8StB6JlGEFH+bQq5JLIIoW61/h+A9reGTCTeYlKcRG2Y4uqbmJt7KtH
zo1ZyIFNGJXeB2g5QzZfj7Ymn9SUG1byWyXcbJ9nydZ27LsHq+lPtv/tHBpT+gc/
NEShocyNo3qQSDPPt0pF3ANV4Qnt0WRICtvAu7Fz9sRADyuTZ0+8XnHBhC1m+v9B
i+r80qx/zfudVUR+02MCxikkD/k9LxkFIJyLvYygI9hlVWcvnb23+kR5CB6mL7zQ
+9Q83rOyO4Hi3lgf1Vf0I1fw+4grTsBPwqomY/F0aoh/WN0a5slJ1MsSWGG7T+Nw
J7mTJg9CPfFRExTR2C93sQwVtf8dhsSCVYcd4yJixHFGLRiDNbjEIwiw3NX9WSW3
J7jMBUpUsKmw65MSbX/VTC44qNFD74qUribOprZNi9tVLJp9tpeF7sZmfoPU1r+s
9n6JdHWkE7IilpQLchKuU7OgIsWXOD+4UzXRShAnNouykGg1G1o/e+sg1iRjEOJz
8a5HvquxMrlh+Iq6VkuYTV+3RY8MU8Pme+DOkJ/Ktai41cq1TPTasusXALlraAPT
DHTTbJmrVUjjioKrlVgRL2LYWIa7DZyV4gCxshTc0A9fqpTMOYcM6OC5NnMPGFyP
ho9+6U6Z3xS1ktxbO+Q/T8MX2SREnnlnBX1+SOh8i8v9h45wbsABKjmzNQSoVGTr
JdTTxGviNpBM7l+eNF7XAtj+lwYYjVNLO3qWK5nz0gkekTlJ7drIVsjUeaRBSpzQ
FdWi2Y/UeWdgGqsEF6VIMO5AoPzND5NLGCdS5RWqpGi0z/AGBfobi7CbRM+CDpVF
VOh4cDZUcvMDexqFZCDNCb8t6/VkiEqAVXhL4PXE9ObXqijbhdICC9RYJZIJfhAE
imYKhCCq8q9RLQsiTe0PDu46Ft1tXQUoPkLIBlQkYMgXkSvLBV+Gi4BIBy1JCeUe
0Cw4fCWx/n8aQMmQ0RInTdZs8jYsFpLV0mRgfZ9TSiRMMlhqHkURPkyGJPoYBmDo
6kIFX0vYZgXtTpATgK+yXEleDN64COmaxAgLVGLLGD2K6MsEmqjF6SdGVDNa6kAN
nflto5Aw9n1mT8dNQstwtc5fYu9prHd29eb32I9xNnBZ0Mw1uKIiqoe3LyXFtX0w
CBLHfD/JekewAn1RtePXwTVYvRP9yd9C2OPRcyuT6I23YpqAat4OMuLHFhjmSnSH
mFaSkkUYkBYwsvkkypOLMTqyOIHs7a7WJ03gHy42abQbcWwoU8EpdldUbuSZLgMa
079abhMgMLRtMFKn0Qh4SGSCEBhaZfx6mAZn+6U2/naQHdExrtNb0wWxbGHfb908
SeEqgSwtDzHGwmC2j+3fDYs1mgJpi4dLe0pumGHm3caS5Vjh7SblGBqGMIevOS0G
gOCRhiRu1xkAB/VG5vZK2W8Y7ix09HBLeOTGe3ueORSoYwQEF6TmhNFnEj16m4jd
DRqch9LT/YxweHoYD/wErew4QafXw74Q2qfrEpizRDeQCgL636J57BQzsIAxgiVe
tEUxf/bz3Exz9hTkemeq6Myz3Oo2GUDllxHI6hKzlB475j1eoohAk/xGQTBuOG20
HADDkSI4wUv+HT9lj9fjivm0DSsvgw6sU4LHDvPQWj10RmT961nlPegTkbz2qHxR
Cio68VVaBOymxhyxCLEH40G3SVSOfIAVUjiK3QiN5GAFC+rOA1OP92marQSBFrCZ
AA3UUPKzWUv5fxA7eIijzJsi7feUFMmz+dWSmZCbHltWCIdcZUH021Mwy3ZpxlKN
g7EqIrQ1CfRsUEKDg9nTDyKPHQ+XdQYTbRYjFW+JzJZ+JUVBQjgXDT5eDNIkdZF9
BKcLhvjZZJW/0joG68LOB5GXGkOjSbetkptAzppOh6e7wyx2ohrFCsknrYrc5fte
JWQGMe6hMlRupMMAtD9yiTXkkzg+H6dfGs8ph4xQeaZ9NTh2b1IMKxdhBTNlAzLF
CYeuUK/miOWdaaIQk1ESWn9gz6N1fQU6XuI4x/ZqpAQeSCvsxXFxgj5/6bmJcTMl
gjf+XQkJPBBSZOtMU+xofliyx8rfqC8xLnDW86Sn2uvh52AUnrojifgtHBfUKaWU
ejgduL8oC1VuFLaeJ5fgeBSTdxl/ArbTB/phJO27vYh+4E0LqhoZvRd/i29ixbzL
0abB58sYJ9M8CJEY4l5FnJfakBGgGWOQEhprIhaYRnjEVmYwTCXqiiorZ48AgN4I
PL4CySe1QxFAmF5nC8O66ZP2Ysbc1t+Xpr30d3E2iQ37k36IirtZhvsn5Mvfe3tO
d0BZPM5MVIeQNBAVoJZrofmvD8f4jEOKsLMvEvzXRidNlKDz/FIEPZy+1WMp5RGM
uhKWHbmS8f0tBP/b5BxbqZlOVsYIYgcIv5CXiMNxpbStYFvoXN6jDINyDHfYXFNZ
Gs6QmTgZPxus/CITw9xNh4vMgsT8Cy1+Dr7aGzZQqLs+X0X+FHMNCb21I16BuRUK
fEWcM1as8csKMqMja1ZEGHwtRgqsi3zDgxTZug9Rn2wQrJbuV5w7K5on84JIEM0S
fYk2H7BtytxzGc1Amcn7N0l5NzCRclRUMi8lEJftAOME1nwuKjLVf6rjVw3+gJVS
SiwHjWDgTXArFtl0+4y9umvEcu+EdLRQNzI39JX3fqI8nMjJYYJ1543hIQEpJefg
/kOvMJvRmTfFoHUVXhsRbae/nWpHX69ulGrAQyQlyhPObxEQ0QSNBUcR60ZQEfHW
Km3RLZH44Yca4O8sD9B4PkaORMlgJ3CjofFuoRSSrXGmImfp7iy9nPfsDTAXzNYO
+xW3h94FL716WK9sCvkMEuPWyfKwGRLmkBusFXhD5Et4pxW9dMJ+khudrSYq/Bh0
N8ZCmpjJhm80U6JT+3Qu0naCJHrbqR8u3z6jk4b6tysPYe1uwgrlKWoAmcXxNLxX
qOLZqnDVYEH9OOqM2q/eT7p/jzNlVKl0jOVXwVmZd8rZ+8TDEzLKyn1qQnrfKCT3
5B07BHW20rNYyzcKJ2IU33VfY4CTdQz7kU1Kho09P9DHYZPrzF6c3xVEz2lzOxIO
9fgp9XqE1DwSM86qwGk2OVSDE14GDRs1GDrDG0ANlvO5Nt4XgB4tuMmVi8K8w8Vl
FRUJglsnjUeR2OPwUW/4NwtrF0OTaqn6Ubcg4lxSViIJJr6ffoRlXPXFL1VdUFoq
z5WgX5ur4Zxg3QqvOjtZB+tebl7cVHQoG64e86PKA8lzoBNS5Q4tys80b927d+WT
KKTygslc5K3HbXU7F15cmS2VzEkfHzN9WqHR1jnLGG+E58sLS1xaroZn2/ksYsAN
rYy4SYnb76mMCZy2v0DzK5aoxC+RuXjkfmHRocAOyXMq5di/boa9K+kjhCtD+aXV
pQFHEyOeYszGjmMIpAUX0EPHCX0i8wxb+s6PL1DHtasM4qu2rG9bM9tJINW+uHwb
6Ljyspu/2MIdE/NLJCd8cfQ/UOwqehboBfIAsBa8SZr8Jq+XAgYH6uK3Q2d4nvjq
oT/4pJOFXnu6B8DWABspmd/HdTmdpVKMAQJm3m/WS6BkOMuIN6Nf7s0m2uhTJPLy
r6JKxO9owgHKfyjQNNGlnKscD3NDzpNXVsiXYArWKPlKVeVCGIb08w74e4zLZWrq
XljuUjRgXEYPD6/zN+hnneevemxKuMl4eemvu34/pqRFQ+CQdq4jm/F3Hzbw/Z68
LqMVKUsgvF8wiGGBElbZ4SnJi1VFck+ATFW7RnxGZDEHIRCsSpnk0IZClRDcQyA1
NrStW4H7XkBXF2x4QnUVUgKhwzk4JaYo2cnrwctO/z2cXEWLIeDQV4eUrlDoGkLK
rftVtz9sBC5uDuJkcmh0OW70Xy0vcZybF+S53C5cSBDkJs1Q8CQNj3UP8BnXx33C
Pq6h6xMZWcxvPMBEJ4KUZPEpRgrmwEZ9nSm9Y+tMrbDtMnE7yYw39Q2ZVApYlGZ9
moNtIkWyjCHpCBqqtPibQEMh54Wk3chvXbUFP11KWSQnMJhIdv5ax53KDkb8gpMF
EfW2W1LMCoSqlG4DeXzhl9uH6sh6Yx1AhA2tNjIokVPW67NSo/syZxNjzGZfgLVA
75w/0Hf2mZq+RK9wFJqF34Jru1bIs6jAYDofFardcwXhCFw029rTeN6u5gb5fxqb
YpuiBxIrhqO/qeLDtCTmqr2FvWhB0r2LC0vzGrHuVereStu2NyEWbHfQK0DvotPs
csD6RO1oa3LatSsGbTGGhsqryst7BvruiuAWH3KzDnodDnzz5SpFUwebtxnPcBe1
gaQMDW03Hs+bt38VYnkNosqo235G2As5WHWZqODk8MtY/0bVs9ho06JNSEjBLjwJ
CxRezBEdhmMxfNVs6p+RydrCTdsZM1WpW1y87wuGWUWcqkfE+diQ8FjI5zdf/0N/
d1N4DMIbRn7C9qv3kZFcJpgUnfuA2OH1H+q3lAhbqux/YZjx5ZsNClVnV1ecLHij
iFVRPZQXMfA5o9OKQTMKJsXZ1wHszf1ggOYXYtmcM1pXz0sNmcpxR71+q8uWoqkA
AUG8k9MyNT5xn2vnTBrLCYczLrNqo3noj/B838h/T3+REhX6tqu/EWL0eM8YhzbW
5OQLE9jyq14Fjs7ww5PXzmlNydE2H70mkiXiAon/jm5njiYCa1gW5DXySnrD/RSO
rBzWQz2CfsyFU6WY3T8bJiG486Qj6PA4901dyVylEsKkLbegORhrv9U8bvgzNTPN
w0R9vlY84iq0dh8HvcpKvttEWFdvKgE7bcSSuE493XKXNAWjqKmspf5IEZDmYJ5J
SgNTekH+aUX4BsjvVNJq34IlDkZAZ/kB9SGg/k28SjTXvJxQaMzOOwFaJ1RsfZxf
I9PM5P29oon2uo5Cn1Tb0yGhEf76uT+I1ljr4lKevrbSga/YN1oEr/W2A37ZEGFO
W9GI9WL7xrCI4wJdYx1EPU+vF87VLmE2EQ9GJtBRJmDiN8kBfmi2vwBKvYIyClWr
suWXozDeNF3+FkKtEw1bzzjxuHgPVYlmiAVJTvT6gkR+l3Sz94vDqtMeuCv0EqzX
ZdTo3KEvWtpj7J2NkFQQThyGT/CMONVeJRQKkwbNn/tMeln9YrBBEJaB96qwkbH4
UwHU/mONVN0RZ8LCYDmybWTMQYq942Pwq6YAj4s7zVMFu0jGi1OpXsZ5+sxfVgDJ
Qk8TYJBVB6VzKb7xYF8qRr5InzFSFdsN6IMEf60i0207dItl/0NAJ45tQTqzSZ4t
ZhdzWgtMN9KEXnlcd8GmWeJYMVbZwvl/V0uUm0lbY0XlKa8kn7tHIIb8jkRsZghI
tRErJVDnJwj6mYKzxtg2XV6GLX7ivK64CeRf3MzJEVhewgnNYBIxWiyvblMmN/XO
OrJWpRaYzm/CSCsh+UXqphZFcE6n0b/qQ5tgnPn8I3GlXkIUenEwVwo/q0kJQPLP
xIgkc3RbzjTfbuCx1bI1+u2iZwhHiJxIOozzLJ4q44NuPVIJqsI1H+uN2eKgVW3+
I6ofa+9634tna8ZEls5t9XVNM96T3o5y64xJo3J7jmR32Iot41NhKhs3WpjuA6t9
zslS11NX1vKyFZQgobfaTNSlplGUAN6hr6zaiC+IapSfXUDblk/5lGA42IWMkRW3
ikiSHxYxDefD8x5YKY7m2B2WRlG1PyLFys5Gend4mZPqivvKDtcEnRabEQvrZNCG
qWnfk9s3zz1mbZNGANxgeRqwH+mksJMaTaoI/YG5tAlGXMoW7sSsVhVZUBo0Ib/r
2ENJ6UmxJ1EGu0sd7aYZQ0J6kMarW+gCgji36OVAcperidthxXLgd/awS+Wjkao4
1FxWtqY9LOE/UcXTtV1MtzEM2zY2hqEUW5gebpf1sAekoy5Km74rCoUeVLzR/ZPe
tfDSwoKBwTezo2wuY2lbBgbvNuG7IAhBT9GdPUfkeoL+kkzDeT9QPDIW+LZPbXNj
uCYgkVNQEEjUXgRiOyq3tjJHvlsCXhTnx8TBABjm9tDlQPoYUfA25OVkGzmF/wsK
venJqhh9CnW2NS15ElB/S3aSY2c4yrd+y4R9IdG8Y2r9zyJb6dYU0tbQivTxRVi7
cf08FLGiGUSHx6km8PO7nJobUCiTrKxfg99onF5rc6IXF552iuIeSsZTbpl8R4qk
iWYVkJkV8W8pnuOwrtJeFt6cktfmHB1X6gbtPm9iQqxaAzTt8bkAPC1igIjm6pKB
MaZLm7KzkTgrDLVWI8sFkQB+JI//DxH9GpkHIDM35vVKiKN0lXO1SZNQEgKZd4bc
LEgxawNoZ5S4m3rL/rVMMycfyxLd4toSubmQcOqfNtIdt0KvOk+jnneMMFLKAFWS
/BK/63Ri3MqsAnyM/1aVwg4KfI/btwgZqAP7+XwVhYV7g4XXL9MIN7UJgU8pGGyF
uH37gOUQM+Jgb/Gl7B+9qTzHyqzXWzkD9wVTGSPgZafyBGksngM5oA2zl4q4Dpgl
/NEdLllDKW8yEKyzjN9c7nzadCk6xr5Q8bDfAd8nv3SuH9oZcDaKVwihDJDC7vSE
E74IVSkEn4kf47vuY4gySquGKjakGMPygZ9tDzRLMKxYdeGYORyuW+1mbMg6n6R9
VObmyYClOyBZDocl6MOjnM9oCtzGr0wb+J3HskauGcz0Dh3nDIv3JA8O8s2k0XZz
2kKeafkgXWqDvbHT8xC98MwrV3kcST/Q266Bt9D879ok90NLOokR7xanRr+pCKt7
j3sCAKSWui4BtBxsK8AgQ8pREmTHmjFIUJum84MtbJPmL3bdwWgddKmdlFdVY+f8
cqJTgyBxw4iBIIv6HqpRTweAxVWDOQ1up6muxebltFXbICCj/SGezAuSIWebINU9
KYexLRMwoTldF4EX4pDCn5RK5YCvsnBJiA47Yep1Bm/oy/AVWSiMDNs5BzLDGupQ
LAqPyBjV1aTljgDpE/FJIYHL+a8e6emn3Mg6nsDhbGQre/k5fQS5IK30TBAI5Haj
whje3zcAQTzpYmJXGQYqxge6uFdA93hccB/HnVO/zwa7guSr5cqY98rJo920c0BY
sI7UbZsKpuNFAHX7FMGMgJbAtxnseGxPHwejJrqSBnLB4Ymgbn2SfuRXFpAS6sI0
v4yjqz0zxDRLc3awc7wvYCUHZigE3hwzmWAvC7k+JCIYl26fI6NuxhtLE2AJWR3F
XB6heOW7TVeBUxY5pnNAt8cnKV4axXOIPqkWGfIuqJG8p92i96+MukKFnDLKe26v
WequpRccXQmE/x9pwY9YiOET+R8PscsO0wCG2ur1DwJ0IwVTD9D6aApNKHsPLkxM
7/MYoDLyO+rYsF6xiTM/vbp9sCpULCHzza/Uw38dDFjCvnYwdzSsLjlgpXevnW9b
WFtVnFTMpJcnjOgEDRRtTsj9Ndolfm9D59lpivoo+/KtuM4fodxnIL8UpMD+xor9
cYqW8/8lgOdV/4L+J3YJsHaeGonAPvat9yk/yA6LHqukD368oV0CA0XT3a4l8xqV
A1Yymjv/dZcPJYzFm7bmFGCwSx512nhJm64nlqbq7fG8ZtvjY9LweNDPa05UyKIr
C3T/WKmDAR/rLqb9w/vQalooqUb2/fgOEpjeyEYXlE+lSZKY6qZ6P1CdjmqNqyVq
m9I0KZQ/DXdu2eDKMARA56n6U8DmOZO6btrDjw/BkeHxZPX4k4+kB6O6eGKo+omn
qrS2HiXaGZHLEC+LM/IJ3MwgAyMrjG8lEduB046DrkckyzDNwyMrpt/6WctGXHEp
W3aGUdS5JS7F7zxhNWmP7EM6N/0dtfcFEf1dGKlOLp5cw0DgewgC2qh9c/ILSTCX
9iGUzCx4Z/KLk/V/A3wJ+ELYHeXewov7zzJy4yPzQ7SCeisQwtUclJHLj0VXT2/f
sXOUe2oCrmuGMt20VKLt7olkzBx2FD3KjSsn7TVVPii9WWj+DwAcBLnht+ZxAS73
O8v9eM+FhXDscb7XgEqjrIfWkUC2sIfnAtYscVjiF94UOYzKJxxQ1eWX3DxAEVfP
v3nPZGtatKmduw3Lajdf5sfA6MB0huyCbWstwLdnleKnsxIJ3KyhhrIXztlcduQE
yeEx2/Nzjd9DqQdaH2TE511n1IxiE9VN9LXR5MlUNw7jfplPizQ6trAOjMSBlI0X
K4MrNqSiZJdQND16zl6O8hEtRPZuf6PNDLjHsv8Z0NgYL+2grhI+SI4rayy8a/Ws
9cWABw0vcbzqGRrzgs+nPENxmuGX37aJQ/Bo0f9HV+UzxGo+1yXzmMTuMuBqtWEr
jC8HJ1pYrjgoGo6wEGcSjGDykXRp9l1xCrgVRhkjsgPRsrjWdMY+BYZxeYzw43iK
g1xfqwWG4TjHHjYtsY/UvcY2XledOH9s3HTVQM80ub4UWljqcUCLPydI35t2cY4c
IFWOnEACvX5DMkvV+8olxZHFD/pUHnpBMM6NY8NKl11g+NXRX5Od2ZMFyfVIbeCX
59BqGSdgFuh/uIHYYOOYqgNKOA9NzSsb4+oa6ZrBdj9vPa3mM5x6V/tQRRArf73l
BVdLZFaa0FUXGq186YebBP7l5eATIWRXEjD8mEguXDcUzW83bITHx7V3dSl9NPT3
rS1GBDjMUWIdahI977enAfOeeHBDVqlA6RWex01ql8ct+TpW6a1ibTo0bzfAiQ9O
xRtzYntQ9J1Yszc0WCL2w3LEt25DlZ/81QoXW2mAn8a9+1nTCUNn9Wyg/ReewBtK
BUqXx6jRjZFvPiPV+wW5/3+v9AMgGrudntKUdssfxkMwRA0O/ny0MeP7y+5UXepi
bJuUA73eVub6RwYlEqdcKAQSKQVsuOiBYOemw2B4XAuFGjbiuok0fUnlJGgC7Psm
QaV7jEWsr3Rfr1ziPLyS57JvK/TXIGV/2I1KNMUifCm1L84oT3320e6bsUyQo8Np
6YorooM+JALJxHprm1hNb+SRoibaZ92R7u/s0vntI0baxm1NV20dLrKZQp+S6zkJ
J+i39OhAxwLDsrXgzOTV2CSraWvG5onC5PG/lcFRe51XN3bFHrjpuSAPURh9kRrA
E+obiBDl7TqbSwZx4TnZU+pZA3TZFQPVofgu/0dVs3nWh5XVoR0EbFMdJKWA2qxT
/jBR8K/Ptpk6pgv5sq2V//QXF8cUENvIkdXY/1unHl33ngiOnnDmu7EC5LMoJoDg
TpLVvkRPSnd+A6RKSUj3VvIOTFybXAa+nlyNHhp05U7Q8qWj0rfVCvNhxZoMWDDJ
rnTbV+ki0MlIc+Ds9S+quCsuBXxRRnPre6GzegmkDuJ3id/pkkRFAjYWtT1sOv8i
kLNTaNRe7J+50CWJ6QfY5bn5xWFAKjREqHPYQFTTF9cll7h6UrYPwV692NfXlfGf
WcMZ95i6/sEr1kvgG7B6bwXIHV29tBApa8jjf4jMd1yhS1zAj2w/nNo90607Qmuf
bR06C9jAXywLxnFAU8VU9FQAdbmdXD8wJqw7PcPUzcnyffEbaVBs/mTT0WnlWp20
58HNVuW9WKf0g/sE9D1vvE0rMEEntoqa5Rus1VXay93PKYvhybgb9n4OyN0yuxvB
sXT8lqBhWb0F4ByIJ9tmmmZJA8DVEARYJAQH2MpL2WdThUQpc3RFjqxY9MQlUM6a
FguOBRgZ7D32OOZbYYoN/1QH2P21eNsHWbHyOfxT89nStknyd4KPI66ZumxnTgAN
4CIPlz3HG1svmo4wTf2iNc79n0g0fWNbtyDwacKGHmidIHWs50JO2IcfnriYWpMT
gZ7Gi3+Dtc6AB22wERN9ychV/EmOD/Hxt48FgcUhQOJrdK9uLQbM0cQOIt2O6bpl
pbRb6VskMr5HRuVt13ZvIupoDj770lBOSkKp8TaaE6XJZvO1ZJolKMPujcMOVmAr
DCV0e6jOpRnCBYHNe9xF//AgYameJxCVQ5WQiePe24O4so/ybAhUEa9i6yNgqTnd
r5SwkDUPZoLR9uoK1PEBAv+Opn1ZT4oI9Oi5p4OMtwmjTzAdBChQ+TOON6LelcM8
buIX9xTS4sdv1vKc3NRW8ZETKTtdauJkLClgG6VdOZkHTsJXKf/pNPgvUQfuxPoP
dJUD+CHbuyXe1GzoYLndZEab4YfjR9Zl1dBkULMf86hV1bJpEjc0elpumZCDsppY
sQ8nYEubEAQLyHIYbQz+jb3a2+sdSCiu8I1DBWMHWzOkZGBYPiDOW9NP1gsbOgZF
SatQwK1lGihZge9BAxD7TYqottCnLfU/jBo3gM88j7hhFFFbaYq9+lWvUbO1d+BA
OT3s+BGzVBYRqHqYtfwlpbSN26rFN5BjfnyPxRDy016zUa6DNWLatf4fX/FlD4HF
AKyiWc+egWVGhMQyxEEHtRuDI7lzw7T4eraBVNEWLBw9vUQZ06q5YnSVZeliLC0a
ecjMJaMzumYnfRmKeDOq4zfCEZpbyvXArTFwhlTW52id/AiXXm/QZ3ud6NC2jICp
+QOSr1+19E8tQCpdUb7ED6DtRGl/tBGeG6Jq7BuOrHw4h1uQDl+rdS6gcqmkv1oH
pbBrzTHa3+jT6p21oI78GIffrKLYRJFiEti9MUXnXVYcR0a6d7M6vT7C/FbGtF18
CTBbfpJPHkFzXI5brep2GAgt6U4phqLOL6NJcJqQzHqPNss2ZG87r3br/ngXEPB7
Y9/ouXVYufEIkTgSc6cn0tkRETw0BikojoekDl5JloZ/z/UYanff6nXhsihS7tgv
XUCzVdXbx91YBCvcotTKNMgsNW67McxtWQOYm7ANxD0AHNXdX2iDlw/8mlSoHp46
isL7dQwlvxShMlDk1thgbWozbEG3GsGBwhXwgG4dm8dNYWKlJGayveLuK8/mrQ98
/GQZNawvvoeel0tZzMbfKZxsDytnIysoyfTbA012I4qtFujfwBxQy6Efar6i/ldP
Y4wCEI0INFH+qWak+ebFbbmuotgZAwrbArIQq/OZcsJW//pwgi8wFfuC6SXQ65CQ
OiDo3gLqaepPYWapaV3Ki9EGNcjJBy1VchIUD68LUW4KPIIexjpqCVm1/j8WLDAs
BykHxKi3zGZ1I02VGoDZaQNqcIQj4J9V1UffOKRwHwF1Uls5ooDh6KNsUThiv8mY
nK26rWPPhaSMuZ771c7fOO0uhXQQa2WOqdwLmwfaOV45XdAkntWDL/Bol/QakPuV
bn3Ej3deR5CsMfQMNXSeNTmIKh0F000gXXK5tgLaZejHnthuEWGvDBzzlC3by+Dz
qIfkKioKl+acUBaW7JpB3gZLqHOjvf4TXd0sUj2k0QKkCSqIGAJuwsk9taIh/icN
tmla1xeNbrR1sywtsXawQ5bT9QeCH6RTpU0DZ2b/++a93+qyF5G0mYplDZWIVbqX
CCUcV7JAO6TWRbn04we89EfBmsLodT+41KHKYViWW9iHvKFBjVPX6FLJyFp2JcHJ
VZSF8j6gIk4i3p0pQGQje+Hl1iboUU+psd6ybWO/+oYvmxDwhUcjC0x9Ec+cVp44
bvKG9x9GvTL2vrBqZCcKMhOpm8/arOq3fgihHvNouundP2vVCOxW+A7HCQDNXCeH
oLw8zrk2cptaoDlA15G+eLQ8xF0dXnWkmC6zC7dx4oiL8CmtH2A+ks+ThzH4nNAD
bcXuhj+5XTQ+hWnVSrd4tG7tsZFAVawxLvHuC7e19nM/+FJwIxtUFyt/p+DwG3DK
uLjn9bLFJzM/8RpWSwg1UEU2SGWhldI4yAisTaKvS8edGK9lGl55JA20gyZ4SmTa
ZnKRQTGeS6HpQxZlti9XD2DdM3H3T4ZqqZmNyc7+heyjrJ8k0+4e0u/SDlf1gft6
1sCIQQZ1j2mUo74HshNvxJKm4At7cPdkeG8vveR806TUVTrzDBo615yw0IeOozcX
Vh9CIcEt8PiVBqTZxl/qUdXoEAyRbNIIKOVibIJlYS61uGIKx3Pq3+Al5T4IUn4K
fzBPoR7p9k8dJdta37r7E3d6yUXyiIhhHTZAsmK01VJXXdVP5Q+L1HnjAOBkzaug
tspmzfd90n4DMccD3p/QkcVImQLDAK/PBPJobT/iCoZUsHv/kJQ2qIESRh4Dslzk
YFo8qkYk3chxO6cSTTx4p8zTe0JBm5IVuVWaYqp6IqslsyWxKCPumxOAA+El11uR
DCgtsv9f16JcKZUrPen0LwHqXIHX6/cTq0vPvZWziYlGtF7ONkYu+wymfYeSaxSl
7o/J1TsOndIdoTkFEnQlMYaojRoRQ9y8cK2vB4Fcpace0fDlqOJnxPu+aBtAJ4uM
aHeFnCS8WL1Vm7WvOiP6x6gA+5Xt2YLuat7mNIR70EIuJmEQUyK9wdH7AN9mrK+G
JgYyfDgeXop/ZYb7IPFaxJYzpqzqNFWJVI3htqODOzMbHp8+ZVnoWb4eBlfd+iWT
6h6I/8rYrrd4/RkrtMIV4R4GP0tPCiTNc00Z//HaDtmADBTAPx8tdWL+0tSf1u5E
S9lksDfrxCW5SAwr4DTkDYCxZOKfwTaeLQcKSz3h9Kinxp3GBvDcr83ozJJF9JlT
5Msv0u0XZgPri/CRZXTnwtnWi4F4RJK9kHh8snGrgC+BehcAaq+t/ljuWzredfnj
8VW2wxvuHA/Z2eK0WN2FrW8r2FvlrndaEXnjAs11R4Mojvaof2qGFh8wro8FldQz
jR5I1WCkMdWyxlgBrpcFQlJ6Trf3SGQns/qNLQ4rfq6jgLd3kzEHuaKp9TSmHqux
6VFk5dqPYMs1xPh7avu3eNBDtX5qoe0iExom38w7cbZKHlARkiFmwJ2K4ugb2O8x
wGMYy46o0pND88jWhi2DR12DQtcEfOXmTwj68EtBGkow9Vaj1Lwz2/jPIFCyw4Zz
ltpRYYHoxT5Pp4XM7znkz1cTpjV+uClEeRpeyVAWUbUKAlgm7f+88Z9TZXoZiqdY
TxCv1ubSPqhPW5caMhPTlmY6YRMT5uD8ZpSEQn60lxZNpeg/OtfxlUSPIKRPJmHc
9+CnYEzFFKiTOsE4JqwET+sUxsPgCp2LDCL4uNcMGsEdPgfVwC25l4a6d3QYKtce
rV9pG7Rdnlmqm2L+6dtPPA2TiGRI9FFm+nuwNcg9XbUEvhrELHDE0tNcriwQxUpe
MSn2pbMhfNVbRhnEwmNINS3b4VA28Y9MkuuSdCJux0/Gkjg1aFV1sW3swghLdAkz
e2tx3aqJM5F2CO56qX44SulQGz08Q4xQPovnv42qcexjPpFETClrmEO4bDr4ntYS
7aINJKDomdQLT5XCWDOIkJm8sCStMVWsLsG9O+6J0Zp8t5xuzDqcjtBt4fPUhF9R
L+zytI+/ilhm3Pz2MUEtVvFP5ECFp3N8HnAYLAToTkIcMk+R9H9OOr4a/kCMJeQN
rSF4K5MCEh716y6bt4DPmjghp6pIBRnXI95zZzD7KrMrKpSQXhk1qtwU5UmVpO6y
+5r9Ojq/1T6A83o788sDvYLEWbgFUgdc3wjQhddbX125ZfhKLkPeguKzwZt6c7zv
2BrHvvPF6DFeb1dVHL1QVgivbgelRGW9/wJher95qc301e5W6VbAuAx10t6jmRDl
OQJLGs9D6fAhWEz2VOXBDVVW24FtDK1mxC6s9Kb0L0AfldBFUzIyG8b+ysQmQj1q
zB6414EM8LbWqUuYacYbuyhVjM4mIGRp6Ye4kcz+y/kcVg79p6nQ3WyDazHYeX5Z
71lsRQ2hyRzyBEpx82wh/q32kzKsOEQAMdxCnnmWd5bI3qmK7RwLFaM+xfwWOoUb
10290bTGw8olmkTsDE5Lt4YZfWV2mjawLvlIEmZHVbwWE72ByKAJKTvSIEspJMfl
gMbEHo+EHX/+x4M1GeZMMJh6w5gG750RQyFxDggn2pJhW6Wwp4HlDv5ApKtdbbsS
2KCDNDn8DCEqve2TpgJd1pTwg7dCDN6p7FkFbEu/idh8za5wSZfrwbtIhnYoqnWR
Y9VKu18dtZraJD1CbMxh1rX2/gyz2nfs0h5SZKq31jTy/i41V9sHvcfu/hkxn7Q2
hQFNLQOXjehbb3B8P5ir/NWgozgBmEAtf+lobjQRbuXBq5GcZNzKW5KHKA3Zlr/P
xHz85GGVUxPi+fUFRDtsu4GKu3uHeDDwO1n4kFshn2UAAK+vqlR4ebKy/w6pz4M5
keWWP0nISnEok53XMNNiNsG/j/2CftSeabtgdVV4HUJA6qQeDKpTAm/ACyu7Gp/l
MZscn49hEa3iaUIyPnVV1MkOvvHgvuS7tSYVQtPYwnur8Xb4ZaCVZ/Ax3IbyPt1H
dOVwn+cc1W5aYJ+QVQ50y9p4z8DvctRq25Zo9+1DIIe2FQctw/qTJ5p+CM0VvD7a
y3aOY79HER9sg8cuAqj+dfrzmHgl+9GsqtDoRHVRYw9+Fup62eivlKR8nH4ADjbz
i075DYxqqTawZBpXdmL0m5EEr8p2nqV78f9pEG3VNZUnrdHqHN6ISsf8MC5N1S2t
JIbWgbQQgpUGI5CH4/1XUcAdPC6oQEnoVYymDMB4U19N28/rCbvkPB9E5Kb9GWKl
7x0QSgH25rjKzisQxIhQIIv3GfauxV9kno+rzUYywgnsGExuYBNDmfjCF0rCjR7w
AS8PQLj1IXJlSXiY0GfAbJTimxmJ5wfsuloNV1U1xLaW68s6G72IxhRLTkxYh9NS
JVLTvdABomA6J8awkGFuuA4VkOnd/OZdIkjdxmUVx5VW9nRbE9b//V62biUu8XDf
8V4lOGp0GTjzNJM92f5Xbj4Ps24b0BmmfNn19ns6hpYFAi+IasJN72dDblFi/bg6
ReuuToljLV6OQMCtqumz2KF5sH1BVbHO8uC7CEgIQ8EXV009Wkl/tV+b8axypD10
GMU0zJDPjg6ICvPMnIEng33Be3RGHicCwDiYoHIDYmNBj6QjtsuZcVLDAx9E4yLA
FYs98Gya3ULu8qpgqS+YRSdwAzF3nK7wKOIxZxWWqnLgSUJEjfSClvV1cI71x5jH
Uohvtib26qsIYjNBSP8BnQVQQXTw5VAZQBrUiL0GYpfr65Bcu0X54+QShCAB++7d
rbQcPTNnXyRiFoR2NkJ2zOtZv/MUi5SmhXU6gfUAoEhCzBq6JSxf6cMSly4M8kYc
aSurux4/3/rLdjchhpNrZy+1oyGgWYOybeFFOy7QHjaDFN7IEElZY9SPCi8g2ORY
/oFCuaZ7FtNl4Dds3jtQOHaD8F4XH2cPijaW41cMjo8kwJ973aJhZ3nasXUBDILX
qegTVqdBbb/Nj/Pt/Xrx+WWIx4SLVybkdUqGZxBX/7eb96SGsVBpc7v5Z0QDqSuU
Qxq9zyKG3jwmai/54d4NVMLGEy/Zl82Nb8J7kPytkvV3Kspsji4r6zaW+1veUL/j
TL32fmrTTq+mCuYesvN32/gSxG9rae8OG5zJXQoqxJSibCh3PZ9AdWlx2+ImF4E4
yW1dqE4sLPaFiHZnCBO5U7h2LcjTbRNgi8WXtIIe8F6t/PqIRGCh07HkcZO8FZ/Q
5l2CM57sqDiRNYd/H7zDzm9sbvoWXFidclXV382xCZp204HXZvuYOEBnSlZG36Mi
UE3z30j9O+UwDgvH+e9QvfwjxDlQ1WHiXcda+DDigiBg4i0c1sRzBTiRYskgmAmb
nYFMkfOGkuctMdYtSX4MWx/68X/x1ku8QmfcRrzPG6R/VpJ0mh5m6ZUpRiADLOB+
5VwsAQcMMowVTS46QcXgybstug6qD7yrE2Js3FJcZ/LodfypV/cETlcrC7OvQCGg
/yv+uswZFay41sEDBbIUUrmabcswzWZLKighU4QFhGl9YYDwSJIeO5vmh7FAyzA1
EYz6Xxlz3Up28S5pSyT6ibW7RurhNfyRP0Lehq0djYPxrngOPy3aa9QWa69HN1Qq
qNU6rpyRn87yk3ksGfQJz6Yr+XATwKsJE/xfqSkAn+UKO+EGhZ1Lu60g4XpuAf5T
vKvP6vJp/r0H7jZnR3JVdx3ufLsr7KaBQLZ1oh03BZUgXgyXen8bcg0KiBtvv+7u
SAAOP33MmU7Y5+/Alo+hUU6dxXT3tVb8xFhUIG6PTrVxidhAEJ6+jReioYL5elku
ZOJUEBH7KWdpeS1Pp5B4wQcfs2R+uI9B9/mAbXI5ZddtPYllVtylteWDNJVNYoNE
vLW/+J0j9U2IA6GrlKdGajFRa7Zha8h7L1rxO2La5Dx6jAv5cI5aRbIu72+BKacx
WNnmVKN5/2wIDbrgfpjHbpmIR96MzHXpW/pESoUoHJrvp96DO4xWvRLDRCzeurt8
oPoqZMOO2lRv61d0tYtiNxEAW+I7yru0oozNRd68dYAAtz+1njf+5jjVsOR11GEm
RkvBhvp32hh7qXAjYuvBTh9EscMOJb6A2jv8p6yt5fakgjLp+LQWIAvCeOX5Gvyc
IfPVacGTOhZxG14PG5bmz0gkarvdomVyppzX/DiGoR/jdYiPQAKWTScDLm1L2aSV
cgT16teE7lf+kjc33dDFTpXfixWGbE50kIGtQV0G841JUQB0lDN0IJzQaeL/2S8L
sUWA81u1VS/VI1Ni/WHhtCYaMMc5r1zoA+ef+DTSsKkQgunnqXINvCmqI+Iwzm6w
xmbPxgE0Rl2T+dLXJ+kmMew8KVMi1ssgVq5O1Pl3pUBtx4oHlQHQkHrukZGiqgDI
SZIHfxg8SikA1/NNXwuiI05+hzU2pLaya1NwoqGTF1iQFmW55r9vqYSpcnNhV9Zm
7Y6IqhTMibaKI7vzbn4Vna/b/y+CjRNtpEqsvUyo0/At+NwOrZWQfXJsc6gXXA7K
MzdLu8mXlJMa82rgMsP55IOgYFvl/9MtGGOvK1C8uunB4sNMuYqGG0ihUDfDWhpl
2zoyF+Df/zhMVD+RsMOCAFm2DtjCZVTDsSAu6is+5+MPC8k8ahTrWi07oRQ8BU3h
Ja6zLW6DzxyJuYSPTfAkSQhEbEhHS8STBy9tMTb4h3LcjBYJ/lZsNwut12Cf/LQG
x/Q7Vdz8BeSZuiCZnvb4JR4r7ngCIeYy5lr3P+h/uu29ExS9g15FouhcCkrgvc5d
aF2LenTg9wAT2mpF9SdOz3RVySR/F8qeeBZlOBUxePyC4++7mcfqk2TmRYrlBA/T
ycOKHPmC83URsF56gG6Sj3Rv9fI1v3DKSAI0spp51nGTtlkgQ4IQy2PXN1GNNv3+
nWooRGRuldgi3vcNl0yOrWUz8hcrHie2ltNg83w3CgS6pDvTDjnfFWA/7ULVj79h
z1LvKfvU4qxUR5XkCSi+dJ0El0kJ78v9nS+oruI+z0TtVpfh80Tz7rvdOm2jB4kz
KSleGShGRHhJ3CjWinnNpGrGzbGonFnj+sjayT2zT6/tEYwRPuV3saozC8G2Obpm
tvJoiIIcjI7ag2XNuQYnroBvnkN64qlQ40epqwH3KX5w0Ar5gmVESxwwIO6wejav
PzMwx7IvBb3mY8uD97mBXGZ7EcdCWREMUApD7rXnkg4rM9tMJy5jZ3RE1eud5YGc
mLdbDPIs+fhHzubH+esAhK6z4oScRPii7YjMO2x3q5oqMPoKIqtyXpH7L0K6TbXe
WUDR1axX0Fd5UgxmRWwXVVsVm4mxVpev2S80g1Nr/fprrl3f55+nIntNTDfWqXlC
zSJR/XMlHzHr7s33vv7QhArkJGDVEnFlhrArhoKD09xKCznP7vsJHiVPwBfEYwb+
OAQ5xydyXXeQNsfbEZGYqdNjvvtQpCBKxHF08/i8w9Ey0vJraes3OFa9R59d50FT
HKRQwRzx+zfCMsjWFjWvDIYqXvG9gC0nG5LQTr4skFMJ7eBkLrnYcOI1iFLOB20s
gm7vMnFDWCJzABnXHP9P92/FQpEI+XY2yx7X4axe+QhVa5MhwTw9oQfPNLGCkXXN
CisI23Zln3oqVcArJDaZj5PvWAZlviHx+1gm9x00ULDqxfjL/KjaOr6cYToqwprz
wvAd6XvRktlPrtGh4wM9en8Ubm1UiuAXc4fTSmbEmRnBuDgnDkLstouu5Ip1WFSm
5Oy0ziFn6fLWIfiDyyMbkoQRV1VJgj51rvDarZd5CGrivwX+ELoYk1KBsoBtHWGH
nyEz/kxHgR8GtxPrsbe7rJHVqghHHVL3DNwKraS1EmQa3WDfnXg0Hcw/DNkqKzqv
sPBRGw7XdeHqReW5Hn4v/Rf5KTyVRx2LhEBcB12JpSUMMlChWz41VO2Ib5iPz6ZS
NvOvZgsiJFg+uDqJdNxgfDcXenVYBGco/Hv/PBNMgNQGpHKHCXX3YXHSth8OkiGf
nBc5WLq3eBg7Qa/f29B3pHLJ8/tWNXdDnCNMCPH1TkpEQUSLzKpjdcahLXJ/eR/K
KEm5XkUHgOVizO4wVbWGQui0qqOuUXX7QwhcKl/BW+EjaDVQ8eLZeiltfgKXU13n
7ooP1qGfJd0AcUzPkm9h5czx2m74KfenrMZB59BkGmLAsMK4/nopZxPoLRQT6TwY
BGXM2XNz61f2At25iN3o7SXeOEzSBubtBHC/WIKdipkYo5GT2UqNcTZTwmYVNXel
ElUlfpusMOsf/zIbD8iWqzQXnrx+st1YBNA4/ue15RAISZA8nusbuVsSNkO1Y/VP
BOVq22xO+KqNeuEnT1suTKrc38s/oYWyj7LXqD2ywKFVYWttsX7SdiMGOGvUD0MX
/WTeXJIYerkZkq3iG53qnVON+dtIWOx12Y08hoM2GlBePitTc/70e62G5YRsdPT3
53vlwx2PogsdCgGufMWMEBL4G9Og5w1Ca1ZrCoLk9t64vT/GlcBbq4rUHvIDKp6F
7jhV5HYdhlzL84fhljA42tV6pWmWahrhWoiddrgqOWdRHRVzAzOdSVIzkM1kfX28
RL/l32suT1h+o6X2nsHYA4iCONGsdhez0GY0B6iFf6Bxj5ghyNE64CtTMeqORsL+
NZ3M8hnPqMLgnvih2G8cieRHBudIjwCDYPiS5IIJC50PmrJG+FUfnWP4SRI3TwM5
E2uuRN45PQrbSR1LnkyOohErznb/uKO010fpcB+gtXQRRM9ezw+GjAYCtB1qt+mB
3cIBxF5dgqpux+f4qYLtDzWcbTZjgIkDajYFr3x4mXESqtL9HqBa+GH4Bf8EhglU
nwH4TOulK+xTevbDZLOSvZvCanuwtiL7ahTHNcF4/kd+5yliP8WsVH8+8hdlfr60
ZnoJvS+d6tC/olf6qe5J08ufn7+kW5DGTKrj39eI9Ifu7QoM6CwMv6sqqA6Ilw6f
/saoxJFvtGvRZDRAx8VzeoIJgCyefZv4ZnZK7jEfKgqem2QI+HuR8tBjnWORSAa7
elLHX7Qefdo4t1QX72HW6tYVcX3TV6lAGEWvIN6p1KCcfSWEY5Of+O4sOF8s2W8T
UtdXid1P/oxqnOf9jokB3QvSW++HtRh8rRQVf2HYTRDWKmRBtO1EhZCkiFBTyLwS
oqgEe+WRNZtt856kXc89l4yDTZLf1qYSUyddVug/+d7Gh+hsvoQkN7UhugcCrnBc
dNMJlj5OT3pF+qOyjWvk5zQJMGVUdQ1mnJDyB5007zCc/Oqzuo+0Ga1y0WZc7HdO
0Mr0fiLPe8vU8VK0JqJEliAxxIHtZVSE3FyqL8J4A1DRW9bMn1Ngnc4wCXMzq/7/
aUj0CqmmkgnjJ0y+06LXxBVO/hxALkYmuYHK3l5rzxy6OfpS7Wew8WT96mpxleNS
u4f7VEt9xRbNhkY5jF+BgSBMJbE223tvkJzlqV71LXYh9attSLLKd7BQr9HeGIkl
g4mnSNVGaCA0hp4UIFbTgpSNwuscDI4B6xlXJjxEjuqzgvao0ZfLsVH2rlXyvDqg
HzpOvQGO2rPEOS2qDOj+GXAVvKB2yj/8clpDKOZ4JKFiJ+1Q6KRbU3sB8OCbsd0u
QgqJHiiQGr40AhINBQ2Q0DYhci1xld3h/EkY5Si3zeojtkWtIE9uSc+GOx48poFn
clutm+8LlB3Z8aePGS5Wx+HBGXJQuxlzVyzij7Jx/kboK+dhQOuJD0uyeS0qBoV3
UUkIEIiJcirvAH8xyU29HWkHrb8Fr3S6fcfIZnfl87zawV6+10kIel3KdwT3JNz3
zBXG5VPOKiKTA6vUr6Xth//9cWsv3OKGcd3gtbVrnBk4ar4JLg1ccFHPq5QLqimd
uc8ba1Q0dt7/WjpxkxmTrsz/E54K9o6IG377CfmtY0ZnwWhqReEfTTRmuOW9yzLd
mPNWGkqfdC5Y3+TM9IWtLcCjTvzoS29guAzc1J0MhhBf/HPPG45YA+4Ny4ltSsk3
d4fIMTxMYjbtWLAmpJ34p+wSU/QHh8a+5orGclSiykxsQf9SkZXvHZBwPOcnxGeI
vJEi0xokqaxLzAvu4LtErcWeVzkgmwfnr2Y1mholtD3S5ya/4i+94KgNOamtGyog
mK/HnNYqhcNspXHG0xY69azrnryG1wkGBKjHbcHNAkfFKteVrmjtuMsvTt76ZIko
FN1/6PpwPjeoDjha/MTB35eli4xhhOEBuE3tXYCV/yxDJFt0jel1Mfbkoh2Hercf
IztbHo+ErzG8FSRXakKIqaSQtT5d0DHkau/pwEXfo86gHUfJ9i8bUD+OY7VEYrJw
lBY5paL6GsnQm3gQ1yS87y/0T6NXSgRL6W/sk58BTxxMkPYEAA3Jgsxf086hGhRP
tlTgNUwzYKjRmgMd8sAM9sk9kg1+PkAsxBOHgG9VWH1CGtGPl+Az6G2SqbUXu4fJ
J7Ip4VTR2qEnkfzQ+1b5pA2l7rwXB4JwpA83jvwb5OmFMFwTcjQifuSVYsm7+eyv
DlB+sf+qWDMhrpsDkFhXP9u/XyXkhYSzhDM0TFocruIC1PtmhQ1GK+fI6FeHThlm
XgkV3GYMQdanBI9/P8SkkRhlfp8w8evDBhL4ihgKXN5bUlD0h00UeJRcb4qgyBod
sLXgPTSoZXDXhd1sx3bJ5Yl+EYRCgTqraGnNusUudysgo2lErnji+Ul1ssKazbp5
KdKQP07epR0SDhEZjiIqGH92hmIvr7TtfBGfa9f96uJBeCLfVdSSJqtewT/n+rAf
3gIE6UlngiGQjUcRIio3TVsNqewV+0rCE/v/AjcGSoevqE06xANI80iJX9MEGhac
uCTaBTX1Jr+Jod9VMm703+tEjNjvgMwuwGPoyUppNciXzL1O+tOIofrz6am/tywq
MfU2qM31804GqYEeoHt68YtKt01II49w18CfUuKb90y8RnopgNwNmgoTCSLWJqdc
9fOMMfyVBBf/QGcNHnyrGMRCvmoZVkCjk7teaL1a9X1x7NLGXD6uqIvFEe5WF0qH
HU9SDCuyUcvKY+lUywsdnRHxvp+cvSA5qgLVodW4pNZ3DVcKMn15RbGQhuhhPvcY
Atv0KTXDMm3gzLE1Mwk57w==
`pragma protect end_protected
