// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M0XyIHpPvtta1wXaBw0KyAzDqINsFa6Sn6vCHLKua6VF5G3+Gxptc3hHiFsIOUY+
wQHTiRpm1ZGj2eKceD8fl3OOqxWT2MZT3Gw04z28NT6/nekbtAxLGmnBLhjlik7c
s13x53VADKW+MaxmmLrXU9poqq94+OIDIh+3fOGmaxo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15952)
v8yQ/ge6ehWslTOnP0HZY+VHIqzjHSe9mPPRZWv1crUAIrAAi4E2iVp6dhFWE99q
mBrtMIJ8Lk5k+hOpXprUfv85JiSpKSncq5pHF2Qgm+EFzBCaG5gYzwLTdkaD6zGc
uxT1ULroIVGpkzWamrJFJpsJqQCU9ihSWnWGlS1aWR4qrt4n6lopFg9/2AJgaaNt
lRAimjl6Hom+uO6D8YY00uZLdNOjqn6j+EQQZn/imScsmjHM4ArhyTEhT5SeDXvK
M2PNd6MVXIyJjdTmMmFWiN5RjIYwWEwID03KnlyGMhS0LCALZB5EAQIoM3fjTqQb
tZH1wl2xsfIyCqJG/A3tpzWkj0JyfY2aTkwaldOr5klcwXlc5f5pxWpRCda5lCls
qsC9pv4qGxLTNmSaizcawXT2Igipg9FVWImCLhdrOkQBve6N3MmaBXqMl2QIqgR8
9jJoQiAVEm1eTiAjC/oxJpOq5MDxgFtTpVPraCb23VnAelG83VDxUF8z2GR1Htax
zaqxAmmQ9mYZDABqyzTbsK88B/oHOb8woOwstw02+bSAp/4yhxNg8b+xYA0BSevi
lMUP6mFzvZwKHd/aTo/cAXh65h+Bo9BTMVY/flTlNhSX2uOT/YEgT3s0uxTf/5JU
E3iTSXGzCP4QsEGcIRN0B+9bBLZAdDAG9o4QQY2NjUoGTh4kL/hUfYhDY91I7Zpl
zqo7s3n2O9CoBJqYIKi0f9cCAUxHueID9HbPMwNsSh8GNWZErTiTZkORzBqtYhMv
btVxcY9KWSCbPiI6gj6a5Mucj9t6BJOPUjmxW3enIz/rHaSyA8IHnYnyGAOkJZWf
VDAeKMfwBL4WeQjJeDlsFgTAlLKM2TxzWmlfOTUaieUsglaXdXErwpk0ylATyWfK
MSzNcnhazPFPvxqGeKdSmaRSYFIDeoTwUGW2O1ZiN8DmVhU2UsqAWjlZSLb4R240
vwru29ddN6CNyttkmAQKYJRgpg3Z/kJVq2N/bEWnqGZFruBGAXlp3VK6h/0MPOcJ
0VzBrW18YZSKBH6dm4xSr4a1E1gz5/i/k7O8fAnET8TT4sFYKcm5X0eEwIQFQkPF
2RfsvtGSW5VBpiGhtaMPo9N3uXZW+mNiwEAwayxM2bx7s5wtHxD3D1NbtxMqJOEf
dXtyQVloCeRY1RX/7W/WifaXjwTLvFLj3/mqiD4twRfU+rqytWs1mij4ORtYQ4r+
2QOhJ2AUYw0o3rk86rOVnOEqFBi8GotKtqmZNTPfQdXhY8Eqxihh1gIv8FRkA2Vl
baxXaRpaSjvM/yc577h2IQpNbl3DaOdC1WTBtSwog7n+sjvkjCtYHNpWG41Fv8hG
sk/1DF2rrdmeoimLowI3croaumSaHc70IKykHUO6HXTgGLVfza9vD8KCrdLIUj+2
rTMNf/5Rlp6ydHiDPY/V+2mwvnsNXSEmKs/VMXOBkZFs2Gmy9QB3Z8SoRwKoddTP
n6ztwQzCW+LoRFobMZ3YxWCeD9h+o+IgAKWp8L5WZnjaN2WHSXvNgMqhZgqGC7mn
sNwZG86+6VsbSk6UrHZ+HbmgKhWUh5n+nGhNsxGk02fL7JaBSuAz0l2lSclYhhsb
63PSJ/XKwK19h+YHCze1agXaCGoLintgLhOH/99dE3Mi/Um+PcoDvReBzpYTtl/u
KeRImjUXGCplw43WLF6/zV4qxs3NCTZXcM2vmbdOU+DAYmawg2kvf9fz3KFLeeNf
CP+15lL6PpbmwXjgIkrww2WcID5471x/A/ME5q/Q9I8L+0ui+BJkSLxgbABEVwen
qZDOKpJOm9pBccIdcBsiN3Wfg0UjLmZMCsPUCnVr5/my8Cnqg1u3GCPrApoqK2W9
IfX7fpmQ4Hp02+QnuOJMNZQXwavj11OAdDpA3XoRI4EiBmJCjkmw3PXuQ4SY/ibO
h3uElANuSCSWhTPmgTYu5VGLfvxa2XUXSD5xbZYffO/nHlChqd9PfHMKD3BKlTTo
Cc4+ceg2SFuaFeBiwG0Df+qx4JzIKklpWML1ZBF/1J4LLTOv7hs6tm3bXEX6UnYO
qszoMcADJtiQRyYv0lab6DlHoCso3ffS3//2W/Uao+L+e9k42cQwG+L/AR8zi+80
Ww15x7hpQ7pFKDEFnVx1BNhx/ZhKUuBpBv1tlZrxxDX8wm+zkRgNd0NY6ask/5xq
vajJ2YHz6l0xhgtu1D2cpkxQghbnzsTAD38ys51cNIIMe/SVHjdlZhMzMI5wuVnO
i/Cg51lsrJHxBPCkguFoIaeV6GuTyiQoNcult7K9/a2YUM4HKh4KEANq8fvo6FvP
iTAMuXtmy6O6/SI4cRWCWPpEsexszLudHFU6Q9qU4KQSoQR6GcVX9CQc6UsxdNi/
H7RyuOft1cCT5/wzPRtHs7n6j98D9QCI7tEVQpLSTxW8eBalhI1mKO7LPsPkpR4x
x/il8wB7Ja0PK7k4iN/6jevmCX9jzz3/RqjDgBC6hi1WLPeOctmCweNw+YUO7ryc
drJSOq3UMspgcIGJBR+eW66Hp5HZTy7ZAHrNO61CJBHZDD3Sdw/kophaFpwQ6sjH
SmwaVVFASpyqx3uC/mHhzQUaI6o/TvlCAKcY8olkQcGb/jgtv3mFBYPApxaszEj6
5AxHBprT57/xrYAVxmmB3P9cpwDRoizZBuAncn2UIdmAVI9tGDtZLtRJeteCb4MQ
ypppzev9Bupqpn9bsqnC2OSxkl/gZLLcvigR/biXsLC9mCXfaXpL2WbuBGNg50tZ
6/xVeS2Qih6lSEKGBuS+hlSicVNQs7UJQp38UuVyDZk9PvWT0L6kPLugE/OD6JrD
v31rnHOSDUCe4jgXbNrqtVcWIZI+PDVRs1lllomLZMgrRzQciONwCBnm/ANArk3A
iJcGOj72SOjq1gkrLC36/CMyY3V0B9x0nBPLC6l5uU0V3599ZSp0W62uZojgo8Mf
5NS1pBaOlwJMZxTGfiJbPzNzMH9IHx3N8L/BysLywc+NwAEyvb2HJBtTJL3gAOHj
wxtNyXPWz2/neMRXcL2S/jrY3MkQwqFcrHfyyh99UiJQjkaPkU294JFCJ3SK4k/m
C32naWkNqI7e6M1LZMHpDDiBNv4lwuv6Qr99Pi0n0zMJVJcl+uhI+wu9EnYYyq+4
xzoDzPIOXBfEkYyiIaem5AuGzFdytFECEZ8gWkPM1SrmYogEYo9z3rG+bjYwuoCC
N7TbQQdx821M77Zoo/BGtSSXb+aQDOPUwsgob6nWDBT/+qtU/+V+QEOIdq4zoktH
+6iTiveLhh1F0g5PwOClMl+0RdZvTFFGTqFw6oYGmgL4d26lp4MuI7dtrDxUi/NT
85p4RLlGzfg3FPtzWFSm4RcUpcLB6/kCfHJR01gLjIQxDNMtvGSTRkJj0BJT+mDe
8v0K90y0I9U+xoCtHOinQqA+6QwW6BqJuK3IN2xZZyaa7QGkXi2b0SHvY3ufL1gO
IoFctJDUaH4sz4cncyFMYZas+YD0n5/8BU/G7PXW0dwESpi7yjty7XhLOBo6jtTE
ePa8DdDtGdHg6sTekS8EYcsoGU0WsnNAMsYmpNjC2REih/nq4E6NuY8OL/ELjPOi
DKC8Z/T9Z6niJDp4yT1jQ5eiznRMV9H9pE4p1gP51OpahTQFW1gM+q5dh4WAVMZH
KFeCMQFCdHAegsglKaBghEFs7sF3uBnEnyWtB91uzit20ZOq5Lw1AAQAmiIDM8Ka
eKt2J+qidU6N4OOsDIVIGa+0RS4p76pB+d6anO544zaEqQ8XgRbJDncRMBWuNMh0
hIEhI/gMPbID9qDXSKkO30qL40UvePVXtcM8D6IgA5wU5t3gu5dvh+Eylz0kCQ+D
gCZiOl+aNyysZf7KINBBj9bcUeTSL6f+e5OuTRzEeaabk66+5EreWHhM0CBdO6fU
38QDYnSyILqjNPpMILPG1rptuC8nNx+xMQFWoJS7q7J4Bjwcm1gN9vVqaZqtk7Ha
fxj2nlJJuCc/kchJHJnI/eFHlqBmOQSmEfni/M14BjLRUbptuIVDTAdXeEk0P0Tf
+LtgTt6f/KkzEgiQzy0qM3k/m0H7F6k2FdRP2AKTVi8vpKz6hFUB/sdE4J46fhkP
STua8dWoAwOdPMHmTnsKXEe/5we8uVr8Lsfq8kuHc2uX08lrG7b3vbo7uqkl+ZBk
sSek/r+RUQcCJeaKr3KyghPYugoz/afQLxVwK5Uv7WAiPJXlwhxWXumN1d5mBLqf
24ttR1nnZiAvB7GB8SGyi97Po4r3QXdeEB/MDP7YvFmnYm+5rk/yy47Z9mngXhSC
1PXCgWls97NtUIWJ36+nWaXOklpdcL32gFpW5M1qslGgMO0D5FBf99LQifQpR3J8
HcV/afarX4BW0g++VqkNN52zG4ZXKW2ZCStsQI7ilQfIlcPfjaDr+753Jx8hAZri
SnkGicnX0Kv9yaR8lLpE3XGT/5LhMGRpIvl3bZL042beyJUGGAzyQgw5uwrOkb/9
JsKONiromR1vALWrXecmkbqKDO3Fv+KO85JwXbpZtA20v5lLiMzg+KFrLwP5n0ah
/JMgfgtRiH2w5ba5OvdzkAn2JlMQDJrupLNdyRVPLUDi20AFggRv4ds9GW75Vb4h
J6WOaCl27p85/GmbvuXRKVkn0GXNJQPFq9xUVwx4madarfDCOmIzeeF6cCa9OgnY
fDMXp0KkBBE65+ysC9ktWgrRb1XQYehdeBiU/vXU56RQOncl7mCNEJDG/g4Mt2w5
wDXPQazCDcfnrNrdl+50+4gE4iBLtL29cGZ6cuRKcTXxo1CKSFdPFCXACp768ga7
iTdrrThHWNFCamfVLKkkwU5Hs5u7jFNFizUrIKTx3kZpmegbqJ6agH8ORyHAY0Oa
oinFus+l903fSOEY59jzkJXMjLwK7eJff1AmULUdX4wQmL8I4wpVheNBd9jT5miH
NymJXOSxfOoiCYMRdIh95TkAJJnmros3Rco1o1ENzqO+2FTgTvip8rJYNv6lQZPi
Vgvfya9dVagg4DNRskjrPa5N4cqeVArk5AZCvq7L0eLvSYnsY/TwmL9yQq2+DUrh
FqRT2UgFLR+XLY/fNaPHMs/dikZmhuxUFob/IHstg1eqhcNGGOAuV33jfdkbKPKX
W3Qe+4Wf974XVZpi1kzjkvvBKiWh2mPGluK9QZhFK98CWe5eAOtuI48WJZG4b9m8
I4EPUYDyDWrB5v168r7QHRbGDK8djpepy2Un98VFkM9OGwsLELzWlSX+UX6HCMFr
skbVKWhAnd69Y4Yg0FwiJu1RfuJCgWoW6iV/bPWvXWT/caO9LP+QyiD/+98FEs2b
js9TKB4MaQGDyuW+CR8WpfQVT2D56RkgAk/QWRvudQHNqUa9emffqPFnNWgEbyWi
8p4YyqK0ESrRqX4tQGL1gAdVKssZIheEkuCsEL6zLoDlS0hph0UactmGGU/9AbN7
aYNmNs6LO56nsuyc6TnYmn1dYo3Iq7co1rsg0YjQDYzVk964ig/4q3wEcvsjQ8/F
8vU4APYqp6NdfbBvhqMO5iu0uiA3/Cgx5lX4etIrZ5obGIAmC+zMpTzAPyhuQqr0
Z1UgR9ayeSDabMzoC1xoLNpAJ/h6lo6/WNVgmU8jxwPXsd3lA3iYyEW3Q5TaLcq2
yZAuuWOa9i5+pezx0MdsesFk077i336qxshbL38bjQSEBNKLf970g5fQOl00qR5J
PE2eaw7xvDumuhWhUmPuf1DbANMa824bxqnmM5Pm8NBkM+Q8rvxH3g87G7gpE/tq
V8jxg9yd1XrqeOjdBlHjcsbgOdrq73UDS8mID2UFHsVnuvVR9WJj7xeRz+yKBZSP
pYfciY0V5/5ioUttCRubH31hrjtzrTiMiLeFVgedHMP2INC8DBQbDKIAhGUVmt7X
8hpGz21Slt/16ZpjqdK6PN6kRBcNOfPcqx1MUbMPzUdT35cnk68yfkogRNS5dogB
AXNZGpXu69E+p0XyjupzoZAlyhQjf4wEkE5GFtOG73+hITBdBZibPnQ/c6E3Fsvg
9SVW+U9upa3eefKbE+jTYcyhvZqhkF/HQVGQRvDFGwv6njVqgz7mVMkpkfNUnJ8z
KJutUjgOWDai8ZyB/40LFsWvwvqAb9D+lIXHt0BHSFxnnQDmChVgH5FkNKx1s/yi
In+7i8aTOz1MZNbpJi/N7/yUkfmE1GYvZcpuC5ZiL3/OcfVzkSWXYcbBpg+YIXA7
nTX6WZDCw4XqAnindG/lICC96qnIwgt7gGhaekdOxNr0nq5TVHwTTBBWCx4zHi/l
0ZraKU7nVwns2fh4z9KdmfgYyB1oq0c+DQy8Vg2NpVFuApFU34h7K217A172vVL9
lYMV1Dyzncva5dVthDtBsPzMNuo0XItmsYfFSH/aPU8PqE6duWrcnukNyrQWALwK
NF/QPn1lVP5Z36aI/BRvAfChYud1yBdfz2m7gNORy5QMmd8QFeUaU/qCIX/wdGwO
rsVkb9OSvaTkVypxJ+BboKNtX7zYuOTh1sqaNE5l6G+8FpTpX8bv1tGEkWqiAvh2
2vbbLIyWUvYpkQ5dx/QzTQhH6Owlo6umaBmUeZJ20NEfk4jCwEvkVBvlxkP2Y8XG
XTIKFyystoHMjs6yVVxdLF1o2yzRcq0Mvy/A4HSateJDyxXYYT0gHOFwcgKenG/n
mdXcV40BPr4Sh69SWl+dX/AvsO/uHF24myZ+75pb8s5eSdlnZ0ONBvuOD3lAijEl
JM8kLTmHUm0b/r2QAb3s+qgdgALGS221genT3FO59GuLl9SIsIerSi7t97H7AuW9
QLy9O9wYlkJFG7wXaMzZ5mm/CFnXJibqV9VVDoBO0kGh7UFEfJkbOCi/GAV6iYhS
GtuetjBzRPgETAzAUD9Gtl5xV6tez/aKR9uEMNBQKGOgsIaI5Bwsr7sMbSFo3MN0
Kz2QuLo10sNo0KvzHtymfyPq1wpkqlCw0NT7UiuLRxte2BulII6h5CUiODUN7Fbi
LSonsmxo1qQaxIkLRjvLu3yWsGp6loWWppM80G9f+tZjqVX+idm6J9Mu7r4jWyZ4
nm/qSyYqJV7JYo5BJt37guuKaWVY88rrbGn5jJjLIGeFzS5vvAwwn8ST+murTnYy
qq3tmNi+hTj40WPcvAuAnTfRmNOF7QL5BwDngq75r9nyfzgTZhR/L9UZX3+mUag9
XO+34FudvWtO07375/pcTp+QQolRAe7uHfXpQooKxvZMB4WjyydjNOKul00Zxuu+
Uu9xweUrSuaoY9yNytObMyb0OXJR6od0+cEVtG9tGbjQiWy38Wt/uwmsOe54ZDg3
IJVBx3/RFn+lQy06Pr3u5DG1h4pOwbnmi+sk1zM7orXbeGUHD7ILeIswYdS7ekpC
GoomTkxnAZ93D0KE6DpbrcaWJjJ41qn1uIDPBMDIPZsIEmuvef9sOpFqhMFXcKTI
4BB7aYH3ibpUPtKkXhKa3GR1/JQtf/BilJM6WdyIdz6cSrVdywwuZLq/3SaT0eAo
z5eOCLZVRYCyezK58x48Dr7L8lyUYdfuHbz4gxsxpxuqJzUO6Me83CKeciVn8ocb
5QFaoiuBRChnOiaF6vjSHTj46yCbtGilliUZu27ro7Hpsi9uswplsnxLnW9HuI+3
2J5BnzMX0L6SZ2CCzc23Y08ug6gkn6ciMQ4f4jJac/QC7vYsC7IEA/SFCqFUfzK+
vQjhV8UyVHVmRMERiiarcHip39SL8gPcCDysJ0iM4ggU9irpU7mDJD23wDU3L+RH
uA9RprSwc42SWJMx7n7w7OViqVt3yrQOizZ3RkdE9RILNfTcNoZ32n4TPy0MaUIq
7fkmGrHozUNOpIBpLS5YFOSimUsyZmAEqMNtCE5fm7n1bBNIto9NPuyD2ApGXlPh
0cyPt4Z/n8UtiiMXdKMQEWF7cXYR1iDINjNg1ks7MzQ9BUI+UrOKz9q5QHzDVrpY
J6kkKedLn86afu6iUkFtKb22ByJnM27VI4pEncjbjqJpwNszPWYRACx2ohBQb6Pe
7AfZtEHBlbgyav/ZmVIIQjmrRJ3J/WQh4UssxyP8O6Bub6yyEXtMyumWaPz5fblc
WKVI2lr7zbfnqzltmAZGK+8BBxLu8JGQ6bv80B2vBfUOJD1hkQkV9PpjA6b0/waM
Yr68fterxiCzrCC7IxDFh6Uu0KkutMqI5wyX4xazRN2xGjowVHQRMYfEkJhbNAnu
joQ1gAgMT8C5F4RMkY9LpauJy0F8NMAccp8tH/aQ3DEQC0ks/NAj2P10C+aXb5yK
fOXXlH+fi96SoPcvmP6VAmaflCxTWPiOP/k6o2/CdqhYyH71myIlveD0vsf+4YQw
D651/PKs8a6RA3XOj/E80b8ihGigbJHl3wx/nZB0TVcw+jCq8AkkXRrMOkSuAjqx
y6l4YOcOUOpApWNVFVOjfcg+NdQ/xOU4ni7k9Ys7C60Cj7ySoKP8UHXdYgymB2GC
qokoAHnVQgfg7t1scf1cuGl9OlpH1Izah/Gfyv8AI3x/zgCAGcbkx1QJGcNxmdDC
mjGTxWJrJ8Iy7D+1fzGA5CU9q/NpjayA4Kfe7sELadbzh9F8B8YuyOjSz15pLZjm
+m+pfloG6/QB87yaErMwpkhZ5IUYaPyCvPoTTRo86PGSxtNWNXVACMYoVZCpstHa
B3rlqtKtT40j2DsvfirBzo839Z2BeMu30r/6+ziYSgKUyS7byr1G60P63FDn0o+j
egWqai6IBzke8I8VYNENx50YF0N5aQVFb59O6cYlQlvZ7R8dWktQmNpVk30vIegU
8u9ASeUFrA+cSFUNHqc3EnCjSXxiM8JEgZUTi2VFVZt327WXLYczw8Dag3bwuW5m
6m6w2vpV6MblYJHAnlGNA9Ml2dIwZrc5G0Zvg4vOzJR5SEHe9vOtdeZRfwIsQsGg
GlDFQvgIaY4kNCpoDbL4t4QShOEqySiNCCBR1SwxixApEN8B0S/+rHPvTeg7UGc9
B4+RZWaiTcfKtjhx1g3gS/gwFCLz9rs/jt0MzpHLPx9cCJ3YjYXY8KUctOjjcu/q
jQ4MzEKOcTTEymJKQDp7Z/mGvR63N8vR+OFHtayiJxLW2vsFapD4UQqgzHbMeD76
ByIU6WK79C4RtXN7ULAPY4A8jHHhOZSqSTs/lo2S9VKHai0Hqvai9cqMc1kuAwo3
m2JX7BtyGhfWMwolWEM5tbNAG2sJzKxqAdLy8rQOQSNNSPPZfmH6M7kAGzhukwHl
VvbWveGyr4KIcLW6akGLbe8GMiM3bplBEg9g9ISbC7JzaUhG4MXwwng5H1R5pwrI
1mvsB/6WryfKV6yt8CvvEUldzd3IqWFQDemOIsUESEMVz9AAMXMEPdXq/x8JYrcd
EoEdfCBsjml4Aapz4ufFRiEcImIvBnx6KQljzl4l35YTQ7J/NoqwPptj/TjEaEK2
P8ZHseeN7UBewBfpURnhwChLL1ebZWHM76WmuNEChMQ/cmprAHPMg5exS1XLZ08X
uTeLTkpWTfQFduhVWX6OO+HWxpUFhSqo/GGmRb+my0534wlesohRUWiPF46XD2DQ
4Rrl7hqr8LsMLka02gONIEtv4Qdf2U69OuZhKss4AygoTHp/6bBJSEVzYovOWSFF
Fh0ha0P7JwSMyhrC3Mdc2EebgBnOdThdV9XJgOo8k2laKx/ty351q+TQ4kfj+GeO
MkqUe+cguJEQ89EXsly4w6e6OQ95/APUzvj8d5OfffHVTHvPtv78FvVi+NSRNJ4x
MIAU1g0BOGoHjTNffguEfdVpVbXnIvtktd7INbYfOCL/oYYQgm53mbsFqjk2Tv+Q
sm3D5NqJchdCyduc7xGOjQUzByDMhMg2YjQTVXtEGVZzYckOWyJENbE5YIhh/rjd
lDrk7Vjka01NzIDozidzOHJf6xmYkgvSl9r1tvcQy68h8YDdw2ZaMtvvxq4mBzsr
HL8733qv+6zCmJelNx7oo+8gBecO7/w7f7s5+koU4eXRl3mJBBia6ZkUVg+MRWYX
KVqfOGnw+OWTIo5oJvbH1FNxgME4azvW//CLrdINcfUAsFmBgOGhTEsZHfpdj/aD
NmnPICzSQAosV1pS55/I/d8+/h7XTmc6bFAPEn1AYkoBja7Nms5YIbr5l37W+rNQ
hVppjxUALXIaf47y7FYvtnjRy/1rjRHAGP+eEHiP5YogcqOgVOIjbtwSoX83Np1U
MB4h35yQcblQyrT/yWuopLQA+0ZAX6ut5IFbRa5c+ogMiYwbtLXmCByXcwez4742
Ipm+76RD6pLDnhb7LZMX6ggBSZHMRWimJVi0ZQ62xz5F+9tjshhydbcOYiWPf0Co
jks23HNXccGnXIGtc48RWrOcYqgNszgByIB9xRxm6HVALU5d5Q+GbjNcgNzRE6U/
cQq2UXTo/D2aRm3iC2UVGZOgDVZlGajapCo3lzZHgazndrytfDDRKEE/83zWEYkW
AnV+EXA0ZEIG9I2HEnCTZeHblrDZVcKa6DhTJYe+OQ5K9A/zEIxszVMX4x64vI/c
al5FXPury/KXF2eK7c8ROw6m9DCS/JkuAkwxonRsM23Xiymf+1G4DgTs8zarO2Ka
cItcmyJHiEIlk5jimNM1no9Xok6HXrxzcF9xV94w3E9BfsX/ZpOQXo4BkSl3OE+f
uIO45MH/3y6Zb7VtPvmxnCoXvrjeLTNM+XaHnXSpTUYMkjAKSbA2mT89TyIHqafg
vnh0G0cVwX8pxLctX8xk8677Z46kU+2IcSgTEmK2o+pVWWIFiQDIfuGmw5ZOoFd5
owHzPvxK7OH9Y8LCHTGz2vbCvCg8FvDr+9M2D2SoPVFjz6wWQdyMuIrdgSOD9+Rr
Ur8ZhXArPRxUJq9b9z20xqnOnIFZt0ZqSOkTHO94xAYdRycDeIjaP75aP+l0Dp9p
6znP4ag/v/efRaJq8ohJP+YzapzAfcOerFlJmg0K8fkaMh8enlEoGH1tcUyVT5MI
6HwrSwxTUE129FjmobjcZqjR8UBaNG3lAkpLuEW0hHpCTTCILBRKGaN8Qr4J0qiB
mPnb6K/l35haHiY//9f3EtRrAEllFbQKcAxQNL7tJOtp8Q7y1WfiFOmA7uMEGHOF
HD70NHaPRrLfnkDbjuEDhoopEftff7xD6m8BHLzs/YBwtbpOWj7yxzfdkzHrj9f1
Wtjgi/Oc02x14YFIS8TWfnSSfKNXp+5ubnw+cJwf5MMnmFng2kM7fVaJ07DKzOoG
U+9qoC/VHPYvWct4Jcu9IXVnb49LZGLkkRyLF8hcbkgskLjVsr59iS+ozbFmBvLb
AWPptxGkqMpeHjC0KpnchCeNVNireaFtqUhKSFRYPAVIRx8NYRweN5PuoBcwCGEf
O9w6+R87d6PqEFULBwwY8VeXMuXYWBwiwl71bRufSIaupM0Ot6HCSFhR+1nnq7pP
ePpW4pNhPgolDWvswT4w5fEtGvIEj3n/VO1KyUshZCIJUxv5lCCYlv0AAxtT9y2W
KWRGwGN06SuCT5rzx6W7W9ZMpejeuf0G75IWMlLjiC9bzRJlLe+MOK6N3xDKOwpv
ZhyfIvrqDtwwj2mGHtVMG623Z+ck6EzeAFxpXa0PQ8rrJIzfucCjESzZqd0zunlA
y/bogHX62AyxNNY0rwvrg76oUveWgDCnyLmFGoNgqDTxtiWfzWaAVKYEUIEjYu+0
ju8ixvLYB89pjVrTXddVTZBwH9S+eXpA3YMgNTLEjr1wzsh5TXh3zMBBXuPM7ByP
TB4Pxm5iBUrWrUaj3lWWU1qjoHUzy95kSk7DsA5eJz67S/RI28ngcUJsotS9XySi
zvn/nhMq0fup6T7EDzOk4TZf13FzwIFssyOsca6pghAOh2fIVg952dswQfawaSSl
ruQJLx0/68x7BVWJOkxVkIF/lhjN/ihu4ZFIb7ePH2GlpPlBJL5i7SE2MjdIiOLt
HgBgJZMwKe+exe0AhoNwgLJ02xl4mrCGmYshYBAaFMmLHIXILktjz0T+r3iu6iUQ
rZzj0D4HM21PDSZhHgdjrBieLkhxXBKT1tX4u/2MUWAvP2yAOz5cvqybp8WLZ3zG
jVY9Mfv2FMwEnPZzYsgmFgVYhUpI17XNpFtFatSN7jXzJdBahBlaURR6Q9/ZcaIb
u5fucDcQsGT5oDY4Gz7l09gA0OiNEkqFhgjFYtCiiMSUAbDyXYPdtBKJ2EOe/5X/
YBqFg2t4Y8NZhqMdb/oOW5t9jhDkTST7hTakH3vQ5xvQleAek0ON2HqfCNClWBzw
sDNllhLPDQcTkAx6j8wBzP/m5xHGectwnlBcccYu/FYVUP1hqzYhBCettMqG8kGz
r36B5PeXuYOOj/Ep9QarI1jQ5RbTVO59y0lOJTWAlVEZQ2rJmwB0ZqTN1oHofn3b
MX/9FKQ4yZRRP2Ned96WxkZvt5sFSqAnccKvxqkWN82eJAkNnQiGMeC70KEbOHp0
KXfpr8tZQdsXIH9REsV/g41+O/33UhfYJ0KsY5PctM3ohXpKSvTxF1q8+EZImRvB
O4jwBhTHZTCjPfp5oXsH1wh+zg00j348dVJk35L0KnDcTzb4MqrW/dsmF7UPlSn+
M5n40z3dx17dkyFfnYzcGEYk8R2DyZlt04zvy/cLVqFnA/iWyUvg2GFXKOjtNsOG
XZyw1wgyWJsPedQUlO2umWRjeCuwkufbOU7ZmLLCCPlyqbKV5hIijdakMTTXlVPO
Tb+cP5I9rfFmTAwcfyFlPpPqIMLyBWGM8+koTcn1AaCwqnE/V6T+VsWjd+baMPu1
0YhE2C0PrAN9dB7+1iVMCnv+N5C5QEQfwOMv9dK7m27NgB3jxqTnVHKvH5l7oBY7
XtD3/vDb+uxRJcziDSX+OmbOU3o0IRy0TeAc7SMDsd9FC6pbi/TzraaGF0sJBTcZ
tcUhkoMReU7s5twV/VOeGm3L2IN02ufzobF0MI4kV/CJVYVnTUyjwtEUsY+JVR9N
Kfho9W9pk3LhVObfcERJ23LOb2rxMActY+a9p1seTUXdavb3cIYhaYLnYgUJov0C
fvNf6/tH5161mhj3rF6+rEJm19VjxwwIxRqEUiF5Xy1rXSZX5wnPy3iSLr6Y45QL
v3dtmW1tqMW0SCWRPiCsgxCM0WbiOh6Yg0HaYQzRwTiH/7Ce1edk0iQvpt0LheuH
yA2k+zhaWVDbiBmcErdWumdhktKgYWL+DRAosmSQXhpWwK/BODFe1SFej7X/bwy4
zReUMQ3NFVmqLFyh2PoYBwvCbnsOydZ6VqSGDOGctBM2toekqc/b54/MivPLW6wS
e5HsAJMadz8iKSWKLqS9Evos3pNWhgLv1s3KKmeW0SSrptfKxR0JxgtSEvtqjgDO
8NtLrkgmUgoa2HJUA6YwJODbOlngwCwTlN0pPaR9mvwUUVqzm+vI6q1LIsflmudT
KjQnt1te12e/OlYxSWuC8WZr73s779VGUJ9xT8uh5qfl6j6y36Ho/zzQa30QoosI
AiJ9K7UTzHy1Eyc10h2of0uusPT/BLg54pyNeCMZGEP7MINsKzM7uNrsq5laCX1f
GtqUv9sUYmPWxaLufO9FguigFrOLn39NbgDAfcBK/4MRwwyZ/01pCas8mHchu+X5
DQ+N6aYqOrUi8w1SNMGEUpCuFLIta03RNzz5CSa0jZDFjkt0r+3hnT37FcEsxiSy
fhx4SlPD1Wyc7BeXgvZlsY2QtbkgD89XygHBfzLOto3IWF6n4ZtPCbAdtPHXyrmZ
a8QvIDXCEiAOvefMmsVgModH4Jvk3dUoZKrtuemQNA/0ma3Hx2SbX50ilGUIErFI
LCI0+b1RRNlo1ZvBweje8zwPjJegIEt5WZB1QH7BFlhWRdh8yYBwQcIbE2vSoikm
Eh/8DJtMSrOYcbr/zeILrDqkf5bzuVQUWGPFItZDMZ25Zl5bmULNKThz5nEQ44u4
mMeVAUGsYpBq+CAbah4IG0kr3Qy37ehT8+B8h5hBMGKPMiqBJgD9VlrTZ/JvRKDj
dYoxBlRa2qQeXjI2CXn/W5tqPkKJ1xf2tzm6xL4+LpMSxdh9fSqgLvDIUytTyIZR
QuJ213yG9lYWPU2kEtznoCMPRTtPMOQ9hR9KbenK8iPMZVOcZ9wEWJ1aIKqVsMMv
oLfAYXbNsncibCORqXZo67aXYVfiKS3W80Cw2iUdrUCDSanVrYtf0s2RgwQ4BKhK
XX5tnV6P2unZGdhvaqpE6xFWBfyglXt9b06UoBdQ1BXU54r+mOcTuKwsOX3SolfI
DRAn3VvmfLq39g5c9ZYp6c2eVGOcIoAMc7t11fAgcyAylpx3dauLN3gn80rcWHR4
6RYxzFItVAOyVI4di9CMYNBW40DUaPykqO9wETyIi9JR7qk1AiPqVP2Fa83S7ab7
3pK8ZfmpeIXGany3NvDIQGX42Pn+2QMlbIbxI/9APM0DiOCe/O4/a89rVAoMyr5O
aSUYdZMLMg133CkcJ4rXecU+Vwxpu6DVEf71tDMKOkMycTyptOc+nwvVPaRMe3wF
ZH96GEe13JbeI6YJpPYMaxiyL+uRd/4Iv99IMXNw4eXJALCvDuoOWc6vAqleNruM
M2jYqnvpuW5tJ37zSFazWZg/CI6cs32355KqCdjm/pp7yJStlRPfRXOS07p2GOSm
xI/wjtQfLBj86zFpjnvRU4aFQOepxCvlkoGlM1I9FEwQEVbRU+auCxdW8Ma171nx
6GmH+zWXdhbZywk8Z2pPxLaPXcXQ3b332FK3TpeTiYVOxOJwuPi/nU2i3NIeCnjN
RLPIMBjrBiX9YMoro6hgWwt/olvMBe4jvxqOpu0SmHnsNMHPwnOlZYUDqoxQDm/d
LSSGcKq7XfqrS8GM2pVQJx4DcHgM/BbnRN/+K5zaFX3BRyko189bCMPVAYp7B8jb
oGYW+xIsOH30G6uyUPkAOxRC5N0rNWq6NhtKj/7ykm1S5nOJ0x9EZ6gk8otWZDcL
fwLliHC6XikWfftNq4q8eM0AuFVfnmbU5PI0tAzlFUd8NB20ry3e4EosGRIOj5iX
NqIcI7CzYXLPuqocXyy8YM27ZKe9NtFFcv7eGxT1Tt8pYXAxJSFnmk0J90bEH977
Cdw9DCMSGGSifN6WLRNsR/MyGQn6xAkHZ8SzAdycsQiMliTRcdGgQXxhOZvhifE4
kp0W9cschNVpGoL3CPUPuZTp/aASbhIpEpwGU3EWe/PLXdwV3rcApinCWKmnvRgq
T62PQ9qry5keC2GiTcEKHV0syztNcPIFfh9SsVsqlc9PftCHqENedmZsJFnJ6cZO
WSndYzPgekgZhNx7gt+9ea7M5m1W8cRRel22UallqRED7+XkMP6HKidmMElUq/tl
uFoOBLQ3CwficXqQ/0eJllPyXAAafvuyOX/C316tnE5hHKsFfsLcWAJXBLX9hEQH
KsvfTfOYFl5YtFZjzV3G7d1RFau34U8dd93CPJTLpXL8kw8ukMRPkNZ5miFg3HG+
WheGaFyDUArZkNziCILfynxykTtZOoZtg3tZh9vjTCiLGAHG5pkUrd9nZ+8pkULm
P3PcxwyAc7/+WwzpL2veEOYa3bsNaTsuCPZCSbnQldDt5yKNnMo+fSQTXa58upb4
gaLasLSkd1R8547YiqkSdDmJvDELw5b2Ogs0MyVD0a425FUFGtw0LAaJGqRboTS+
BVRlMQ5aVekfrDv0khe68jxJYP3uQvCabYUM5Zs4lyAEUd8aV+tLEoAI5O2mkxAx
hj2OkMSQiSUARz+WPHULOmnfaJHBWyQOC+dUO4F66qzXFL0GSOhvRVmljBsCnZRK
cmsPozxTLY/S9D4QVvrjVL63Zw6fQh34MtGIOW/MWxMjo4if4pq+bbCZdQdGKSDW
/p+AMIirI0i4g406KqXjYKyQhlwTQBU3scvrEW2wGDa+3nowMRbBjv6H4xp+Ns3a
5jLaOQ1eko8Iad6U0x43CxnQ0Km7I6LggSFXLpjxzX/TNyn3uLGk8sIRbw+lPRKk
tUKtKMCVsv4F2fWdN261D55Zj8Jv9Vr4MGaivrvHQk640xsaNIYIj/PPpjmwb+W4
Ai9KTXlxhVaoTi8gJ5QvqdDQb7p43tGcvQU2BCX3pLNDMkbK94cVBXiGDmkuGANG
KnnDaGdm6UM2pgS83cRlm/gnJuVKpYaFmyPP/cDhWL6S56bCTcAwlZJirAG5t0yW
sX4xbK3OGSwLGdeh9tSP2EAKUWxUY8bDWPQGiIINFUtM0W2ItAwDYI3Qc+9snWGw
CyaNJD5cBln6FRRY4OdvHp0TeSrH6c1kXEcPZQFAzNuEr8RL9Ce6r/785kSbrFi0
T+Jl+WZJE5dS51AzvGOgfDCGzPEoIlS9njHpN02vKXxHbvUWsCdjv2kkFrZiDIV8
TQxwbylyvuqB6mzHAebkcJ+FLu/ApLKyQ3d5s3CwKxWoTRwc1F0SEHp1pINjEUk5
zxKlPD0u80MNTCTtEulZyPW8ijujNIiYyfaL2PncRy05zyOQbH9NChUhI9mx7PqN
ULfx4TeS2+DDKMtCmzqydFCN10Caf7wPtenSR6farzaPpOOFIaQ6cgm3rHTrW5+9
cwtwPzTSwfqgczrltAxvNIo2YuACh9nbGEvV5T+Az/vO3TWEgUcOhFUBDk+HTJNQ
2lzqRv6xXk+YmQhrg1vX6wFfMzDfVv5bqDDtopNZCQoOYsSnO47O5l7MOIjdJApS
o2tT4G0azlV3nIiT+fBszoO9xXmbBzreD7STLGP7GKh/od1Hu88oOx5AOF92CXxA
qZuUaMpK5s9oYj0wogkncpXCypJA8FJalA2cF/K+v+EvtsySBjWKawxF69FReXQp
paDh4FJ3/RETji23PX2WRvEGYIYdmBiTmVPWzHES0wf8L0WOIp91OUD2sPAliyP9
n2CKo/R0/rvryDqwtAVlv+bpCr003BvbFdsgmVbAuOwugCKTjNjHgrG5yfgL+Ww9
IpbmlDqq9m43ZZkSw4eVwZLWH++9/KgxkUEDe1rQxUO66BXDllGWyHYj6X+Pau+K
k5If0wuXL69/XBuZvJuotkwsuCvQ5M9MqZfy5aWWQv+F58nhcAIDuhEURc+j7sQ2
lO1SxmPOZe94Lbn45AWXF3zaQ4Ie+c070fjdryyR5LE/+ouf+X9WjbBNdrXSC/Zq
nC4kZ8ghp9+/EUQ4R0OMWEObUPgVC4xwDfE4i1Z+NVlzQfEt3wSKddcm0gPGD8DB
Tw//VciHmbogBQF8VmtbKsmy7ASfqASsP8XrGTta+vx1FqbyWvQg5bq9sSOTmZD3
meRAs5LdamlyCAvSoKMW0gi3Ya7jwW5fJ1tfqL2JhQfseuDr860aqh4pFSc5jfeA
BoJKz9WMzvCDAAD2JMGfKGwzc7m2bM2DQYOgkZgsFSCIIk+AA2KMCUr8iymhNpQv
xvOnvSR3N5/yU+EP8IBfzxuOajx4Z/4xmxcGuGBidLPWX5rOTKDBgA6Tk3E0moQs
eKs/bksdW4iyKKNTxQrHStKO9bFBTlOctQ3R+NvQP8qls1zIgS8l23dCSI4z/SbR
bSN7fdDbc5d7Cv3CzNfRU7Hw4kYapFiYk8Jo2tIs1U6CSRswKUSGeJkPJyBycCYE
HMz/NOMCUbuh0MewlLlcuO3qNVPTWiaBJi6mE6JCNVdyMfx+I2IyyIIb61oAFsPy
UJAlK9MRYUEMktg9Z9wzbeNA8ES9YY9CQXwnIWWMQgN6bmRyaGlBq0vHcZF7EmJC
CbEOv3hj8md6n32Sj1SDrW/vBGfbzjSpeT4Y3DMxMcyKRae+GJwagpNdRGS53G1v
ANbIwX9Df9OJRCRDZkB9f2ZcSB0uCI4XFrKWPonZv0Z8lc2bcRRQ/5uae4zNlvCH
ADF1/EsUrzXUFQpLpAezjalEjQX2end9lZmiZWhgYm9UDyP8Ln/sChXVdYs4Fzgl
XpdzemYnfeqpbMRqqT2M9cO58sF2yaico01RZLzL7uAkPY3w5vJhvFDIZ3F5Ifle
ebW/RpfkQ8i7D20hKujhcPmYS7ZjFImjF9Y2Sb+0RH6Rj4oaWKp7OU0Laxz97297
MDpHjxQH8JqeTWH2pw2RrIblqGFklYi4IWJBPlhPxB7NEScu9GRHPG3SgUx5pKQl
sYFspL3ErCMxTv/1J0RRmfkYYEm15SJV21x/Qh+hcNCAkSvFIdD9kZ/1tLd/h9vI
okhGFYmdWmkx6nxQ4mL7+/iUne5cj7bSePbZsWhh9tHRExbXJs4daV3UTz80S+Bo
iTnGx5xh8rCYP6fp+x0xMDbugaPewxwA2b++kSWPMd+IH/b5ytkXUQMfo0ApsPkB
jcdftawepN3xDeEZCcx7VVg0h7arnr7A+2qhawhy6uG9pOYJCEedKET+edzRMAG4
kqpGD465UENfJ6GaveeQVUcO5/f826GZGXhXbLg3RA5VHVgFWGqXYpdgRvsiOru/
UjpwOA0aTQKAyOlpVRTFHlI0LhKRn5KhetXuXmAX7coKnNo1F/3+aulrCHzIktrT
G3Zkj6goMZ3G4aZOIKD2ZHX6sSQiYbp7iE2dPkr4GFu7iCrpwjf1aKEKHdGKLQPJ
9sNvmX1rSvGQ/siN5wzr+Us/xT/NF35WoQ54qCTk9AMC6ni/x4sn5EOIYZ/tnfMu
4QjB5ZkJvEtCYCa0Vci/eIINmWdYwNnTTpZ/4L6mSRa8tuSRkSyHDIEzhVdTZNIx
XAoS8p/4Dl7pBjf8OPKdsYUrGogyj1GWDVpzH/b99VP7bWr0Wk285stH4X3G5Uz3
ljN1qN3LrFCRi87j7JjhwY9fcetNwU7EpcQyeksyerDcLcKZgueCrIMyef4T/qz/
I+T2Tnx+S/JQoT9QEzEW3lUw6gRrFhamVGPLuZKAa4PEPn02JLWkcrm3ELp+6T2B
j2IPcfPQcYf/VF382obnFtu/d5ll3rchdA3RnMqoZ49mketIfhm80rgw5QNNllI5
kwG+qZRh9SRtYmx4dIH2ZqrqUStYAcWJwcbuzMu3LF0PCB0OKeG5W1MG73t6RcZ4
0IUH9PdJbuzcpdxZngJJV6gsMgJg9631XNnY8PIDKo8DbXBmoPtJAacsanVhvtck
lijhokm+rmwaC5Jlgh3VFppJX1Ko5gUwbcHUqkvWN7lejlU6lCUbNYKsl7YEOiIG
uyTxtm9txlg+SIiLYnkCghJIceuOgFZj7wlXd4jhh+X1TMDwqrerwGWlis885oxM
6M49LTNAAUX/3E6a00nWuqu/Q4fL8zVEFvRt0a6bSAdfo0mECS/3n2bQqGA7ra/n
aVgp17xjL7OxOyZGrIzevAFm3CAmHaao7Nh9YuPhqfUDS10hGaWNTPAmBICdK159
viph4229yEKSuXPjN241cMQWHlqvJxNjvNaV46Sd8R3JuFeh9uy6DEDmRsHoUWJd
HaRusF1nDcuryFWm6MHeEgOF2p1Ut1umyhph3hjmG60Uz78+AEuehCkjmylup+cD
I57mVVD4vSt/J7noOBx1RRaKZjoNOeeOKVtB1lHAWq/gjsf0fRrCdcy3qaQCU8NB
Kyyh9uCtpkSyc7PkIuNyFYDybQmpTxF3HUacMl4IeSI4UfA4f4LoNtakqptIH0CA
z77oTJSeoONQmieK10XmsyNoKCuYoeB9uiX9LrFJOyAWKwRvUQUybEUmSLZ246lt
JCUeebx/UQZpH3rxf92kQ5/MjlmQvFQF06wQNy+HyY+FxkYEHNnu8QEIJQeAcao4
muPhLKiUUjbrlnXcwR9NnKTj6yZeWa5Xi+zhnDScziDf91WC+MM6iMeQ6RFWkWFe
YurjOZ52v3DI5spO/jnlnX6TWmh7rNJaPr7aB9RlkJj6fSTeb929XoJjYcIRr16N
3eVGXoG1/YIotGgBAzXAqljYdopNQREq9Eu+uXoo2c96os33HflvHhVq1RXP9r5I
EKDOsFkfdAbusfrc+6DRysrjAJX1jMnDqvPp7hOuYrqiv8HJ0HJU49UtnO91I28B
pWu2US7gNLeYj5AlbD4baotvxFat4LzEmDgzzbs73SqSXJY1K9FvJor03Y9v1gRk
ZLgzV7QVuZ+JWNkHAoFlksK7PpDu8rIUDkZpsYVcFBmXJhWRzhyQxyW4K73k8wUU
joncj0Ecm14MF3xYjpZW3Nfh11IkkTxQ7t1+nh+xjOzaSaJ6OWue1rb0v+xLWC0h
7F0ctnx4kgO/d7OAIMBPkggeiIJ5vbZN4V1ziku1EpaK+kD4gMmY9R8+AVj+k+ei
2Ya/js22gRP6y4HzlMd6qI/w6ko2YtioRIwPZ2NPdvSxTf9Cl0lfZ/eqmWkOB2uE
k2XziFZHpNMM2OrgCq4XcckVvc5vXTPjfQ/NSGa6IT7aN7hjwT/pu7GbJK2PC7so
6nxfpL/4y1wXukmSxeSOmWBEmEWpCgsLXvvOtJ0beZHqXSO58L7JlmdU1pXJ6c08
LnrkHmYCgg6O/GhqP2gOWycpySS1nKdvhw1hZ8qsSXxFMg/e4M9J7XOI25qRhG6B
FuC0Or+0N9iMXXQ+3mxl5fGR7il8Es6lZsSka9F2uSUXDYvnYnrBFyA2SAbGbg6c
W/vG9iUwYOasPvaGsChR5PnxtFfz9NU+/bE/jmy0LDa8i9e0hVnAlvQrPZJYPWck
23QD2z5Vtgu/pFmMzC6/ZlLvLqzZ+V/EX7ovMdUR3B8ibAt40Ev0BasrEwbZIBg0
rULwdE8b45REXnMwlWr7LZqnu6MWhcTsKfsAdTlbpEAuASA/9Ef1p/Hu23rE5u68
vNEt/NMB8zUS95+OYAWtOS4ZCKbKBaqBSdm9N9HXY+NeGbi7kx9i2zbWmL+SSGO1
mtXXyIPGkrLTjZ7kRCYogldMCzy09qF77iZM5tC+fh5p5zOGtqYClJtI7lVLL7jm
tM8ZlStpppzQMnJv7b3YJvesDnxJLHAnZsioppp3YuOI2DHyfvBNpj/gvMQyeOgQ
mvzP70ESryz5b5TD3/oYHTFDpr/ZLcB1D05CDgzbgIObg0Tc0R49oWsi2+Yy2UE6
hi2vvnYzqxbgxF0s3K88/yCVa5M8j6LnkyJep1aWR+4aSzj37+PNWu13+K59aWIR
3toB+Ju2plLUxrFkTFoJJ9JoIF1TO+UtU/2NUT27F3wYaPNKNca1Laux0hQL77kW
NK2HELYCnMbztAq+iR1UPq0heM0AYU7+e9pvgARvJI+ci8qLSzaRXX2+bs1Dr4lw
EDqHy1TMRW2xXGTaiwH0rrd4qKE9kVA19qTXoEV3zR0UYWM6FxqEVWh+HALrzQMv
QIRJt7gE5v3BR9pOl22tlj6Sw98E5IQ1Gb6SznwjpIUHqKR00tOcPtjwTykLcJle
RD4ye/lRL92twmxoXMaVTA==
`pragma protect end_protected
