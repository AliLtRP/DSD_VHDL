// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
WuajJprBqnBMwLkUMnILKRRKW9Q/zxc7I305EdXTqxLQmP+3/+XavJS1Cyu9c42zvGCOLHuas7HL
CSsjPPvlsf0HAuBk9JoFZaoNLo2anIDdeuUDmkDuIpYMbNgAWjt7VPK6o+JFTwJdxbs5IyVh3nlx
6BdwiwvXkdBDW9yD1cpCD/KtlontDQX5ZBrwRu8N+nDsAeVMKmq4nZwcNAHQQ6tU82+ihd1CCaSx
QUGdnyMGSNJcV0vrsTO8zNRxUyaHer8crUAaOuOak2G2X0oEuqTivdgPCtZPxCRQxnbF8egF7pij
LnhCz8hYvH3f14KksZNEwfGFMOP8gWWX2iSzhQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
nyMqbwbQU3tFjdt1W81gur3iIcQsdoPhP+qVFoS9V2gafY+0W5Uq32z5lQn6WhxaExbNNnpAUcQ/
PDNY424m/4u0tZnZtHbwbOe4VUP3TnuvqlJyDliW3Voi0MAerDuR6WGbCc4p8sMKOW+muhfSnXCJ
X1smI5/1gMCGMy1hktvWmr9e+XxQj+AZ4kKMaTGTbF3O9CwEs+vb3gjIW9J4sw4I+zmZvmRNVHEe
N/hAw0zyItjk6RIALklxhw1PtANDsGR7Hxg3ElNjQhew9yDMPswzqds2QNPI6+UmLNae82S7SU05
lGwP0qfv3QN6buO3MGeMdZkQakVzGQMeqWsj4vhFUJUC55Bf3Ou5uIkubIhBB9e1+bm60jAOQfBA
kRM81U770sE35l7oXlK4ZEBJG96irh8Z9nbIpU8oitP23rmrjiKAfvrphzHvXr57eP4AXykcp6H4
qhmtujd5aEBkIR78XpVQ+WqtlzAUDh8WoKYW9eGZJDveVWGt4bEBRCexbNOCARILK6wWi1WYdvU8
Exqy2Vy0prvnYdC/t8Jp9YC+Nyf+i1RokQSuur5a5HT/47YofQEzAYmZNIR0ZckMAgtSRvdfcEDI
NdcV0SeWKIFhTnx/l5/2E/NCcfohWrCQC2VcdgJDaQNI2JWq8c7CSZUTy2xqxnHabOI8j2dNDgs8
vKr7uVHOLdUNRV+KQndWYQDS5rs0sljHWltrRND3LV9fGNfnhufzQ0iqnovIqKlK8Rl93Fev5/ni
zELJHFweHjDWcRyRA2Qk6xUnxM9AGDCmHT2v1cG99PjGYmzp0HiJepaIXfZRIOSVEW7KK3yx4T6b
U2rWJ6iwpguvVbu9V4hZZmu8Ugr9LnFm7rYzHFiwTq4TfEr8eWiuGgmMmX6WnYZzLWXVQJxeWYNx
UwSp2JGn88Qc4NUXuce3Jmerdf4ZJb+m6MQhY439t2kB6qdp9LDEFWy2d4V40Dv35y7hIBI2XwuF
3MODAEbB38TRH3D5otNG1h3RHFckcXt+glEJQBPW1eOXMmsYjCRihh8aR1OtspUplKD8fGFstH0I
j6h3b5QTbGUNuCA4Yrtx49C07DkUFTO+eP9ECWNaPrK52nPoP5k9haQYHLqfOj0HNdswwOfJpAqL
TegoffwGjtBfVAnHCO2MqegZWGRRlq8qEl9mspEbkB+zvV/z5NrqoL7EFSHJTjcjv4oFZcUJF3Qf
9Id24yxcqpGUTUY6Bxi7V3ff/oPzL8KBbsU/it0nWkH0yZ9tR1xaI8jIqBtyp1OTreVU0SRvJBb+
7ebFFfyU8Wst1XsUYnQ6maA8Rtfl1jxSyWHNHx+b7corFDr0LFeDl9iSyaytRY6dZtGCd8L0hwRX
cXdZnzqJB3gFnxmN51ZjjIIKytym7kEarpKHf4qsWHJwql0qWaFbirbQhEGdvgq8JerB4D6HL/RO
gLppR8JaF76z+UQxPxnvEpOkNdKuAgkCiuZHSu2dEZsyNYtdaGx96kHPO73az6UkUMZ6cXBH5IKv
+xpPSqYxNcsRkrF0upgMwnKeQK3X5dG2DogufAFu0xEetoYNz/Hbff8xHPpxVQFk+Adc2QiWvJ6p
gVr9eAix84y2L2SeqVqHFd9BUXD7as2q10rJInUpj/UePM4q5SffArXooH+z6vR3bIsN5XUlH04Z
z/PUXCgyD/CNjUmr2o1iLipeSfvVzClfLmVKFeHFgQAXo+Tol3XG78QLBJTa/Rg8MPKhh6jb64Bl
WvvmEeonTMkmoDs9IuBwm5AMvnQk+XI/7wC1Xj/Dh7rXO1yYnQ4DuucZ+0lfQsNgUW9eoNIViV+K
kqpnU2+QjRBPVNJi4N6AKGAijxU0J5n9Gp153sWHq5+HP1o1Xkfkf3e8xdNmjqL3XpKC7kyQOOw0
wn/8Svwfz/Fyj7LDTPfcG2eyql+/89DMLm3Zvo16nT8DPe4ktq+QFrn1HFgJr4CM2yb09Mlq5MEl
iDjVQL9stiW6x8QE+U1ESveIy2E7K3mm0+Nnw+OugP//4qIudxYK8TMcScsT+Mzi+LvBfCpxFzs7
dDmlw7DVUAfne3I1ee3sQGSolwTxAZj4FwyLtzmKFw4u3d19HWtrW3cDMdpJtiMsq4qQi9kxbvna
ASHlDnUnEch2htSufqypTc2SAi2saFQ9F1PHECO/4zXqTYMlYn/VTWXWheZeYtc6h7nvZuHArL/S
C6Mxso5Z8vmkF8ZQDX4cx7wVYBYFDfbpIb9okfh2qdKvcptzb2ptWWfyKjCU5pddn4p4oITKJ/cO
zRgw8AZiu9QnpHievdcBTZvqAgWvTjSjwjOUmd69IlLyJWfK7fMzGR3x7LA1XJbnDt4IXYGA/Nzi
rLIxInbJTUqmc7taenmzNfY2npHZgx5tLOblNffy6tODWKzkuIq9QoRmcAVJyfI0fQnRki6gGeWK
ZhE+gxY/o2zmlRDKIivZX4lWX+cacin9VKDBQfqu1bwPCpJqufYIqvWT3MDtXiNqLovG1/zlw65E
buoDYqEPAN0isAYEUO+1BhPm9Bb1SodfZxSJy/Z05FK3bsdUUUGTXZ7pNw1RbL7L69xxjpABrBAo
upXUR2ClRBO6AGmAvfNpxT1w8AoK5vWYtxhZMvP0g7LQW9HNd9LbcHdDp1yqQLmqousRNQuHteFT
mDPgasqiS8cwOR4y5tkAgba3VvLqRyQSQ4EphqIk1ADKLSiLhwYxLIIQiDYuD6v7oZFWJFjnFXdF
FlVKW/KLTAWe87B2JH5K3pivQ8MKX5KhCO9ZZCrqQCL4/KXFek86AYvbXBkA+o7na5rAzaqTLXTw
DkMInsVCQoEA7jqZYscx15J8CtgaD1gP7nMjDy2WgM95FwbsO+aoVBNGTDHzXX2Oz7IV09MW/JcS
4qGmmNF6AopeHIe+hN8oPgd/cl0BsvdBRzB0Sd3qtHp/71F1M9G5iCFuwXMMm4N0c/0VZga3axc1
hb0DiR7+4BX5FWgdb/HNEYzT4eKwCJYYQFUgwsYcmNNCpJSB3aGXej2FWOYKtZtE71RFBq+R1emv
XDWJZUbfgQH6sQNv05yj8DSYV5fO9efKk9ujr2KQ2116Yrg2cJuamIS1IVXmAlxsNfR84Bp6puDY
LA/CEY/GoZp8jXHM/Nqyy3kcpsTQnvK2IUrvAJtxs6dQ3iHk4vPOgONpVo7oGwyBDV18+poJYZxB
HZbPnZnjTxrzF54Vy/o39Yla9SN1uS3FZt0+g60r7wvtPL+2UPInUQ+nsCQjjwaaUS/F5Shpk6Xo
zi5KreyX+1v1OWS+Y0cxIlgjqzzJXS2aNDd9hMBWkDwM1bfUTsdkx11+AKvc0qz0fTr38tK8lLjQ
xzU5iodssxz3Br1ooufE+tU9izyjVzs5Siyw/DbFxa7ALXwPLxS0DpSnbCqb2OJhP44tKVhCGs8t
oR66vsWDYdNQXrihL5GLojWHX5dy9F4L1zm/O+YnTymMOpOXMhhsdBjSme9+ZYrlavqR8QMkYP1g
ewDWVprLRD6VHf3xKdIlLnFrZ36upjE9XkxI2P5WZrebL3cwFokiXFdb1THpQjVmEaYGFB0KSXCK
fm1B4jl3ixQjGFaJGlGppEz4XGMjNMngb2+EWQznTNeCsXd+E7BUeXWfy0wHVHspbl0S+qtxZOH+
Bc9vlSoI0mKv1zwwtqCFtC1DgaZ9k73aITmLr//SN1HCEPn/H3XVtRF10yTJAl1B5qoMZl9z9SU2
ACUwdY/dVla2odEolPbE62NbklF1RqUFU5J9lzu+E8z8sngnFuM/dHZFZKlQvIRi4HVYNGPyZSHG
EzOiXASap0QoJXl2sb8+K6Br2cpbSXHOSSZXb3rLlaSSCgZ2aO+y2Ev7OTh8ahBCotYzL7K0eo2Y
ZpT8DdvLKo1h3I5qXRYTsHJCNc3HmsZwSF+tSfQidP7IduoJlwb2A62NkMFEroxH0m0cJeW/mB55
SlxhT2yB8W7gVnK1yR9q/v70KJ/JsOMbsgwF95jJ1Ae9fhKb7r4ZKGEHMc1IVAahLKIAFj6jBbmD
jGaVXd/tae7JuSZFKogIYPy8Jkthzo1HKFVCHGDQ5Yg/VqGt7tB63u7msVx0uDPqbbv6dDZLHa+j
5+rQO6sW/RNV27UBI/t8aPakmxbTvg2XoCJUh93umU6Ak8uPXNdBj7ZG1iENR3NYHnhh/I46G7iU
QG6qjgGXvdaenMCo5FtldWBZdxkxkxPeaMO0ecF+fMeHNA+EUgc1aJINgcc8vmECg6ZZA8IivuZJ
UWM9Ui3iv4s+A38X6aZ3BCXHBK8ITLt5vGbP3xak5y/DLNr3Ti3ZEXlV7V1coBtKLiF+ZCai5gT5
SMCaIgleQmkp26j64LJIs55BbKvP0jSjqEvap9PgTbcbc4ATZYlGdQI/1wcCZ2Xmyg8H10WZ54Sl
wMEnUddaDbQzQjQiMaoYhe7SVCuvCqLUO8UIP0/nG9SyctPMEB4uSstKABddk3QwvFmihrOjLBR2
dnfv2QnicJRxDecT6WJeSV9TTYneC+iq5s74Oxq595V6WnPFbpWob3BB3vJ62jeRSsES7pwe/swp
qCbx4W6rObs3Y8oLQdtZGbufNODnABirVw+06MNs0acnHoXugZ30hM/HsGDIzv5aN7PQIFbNerJp
J1L6b6IglIrEtDI4QbLPJ3oljuRV8RNGKa0qQeSoUBHQS0jsAEeHfukl72fjGTGc7GWdJEWnWZAy
ODKrDPS6e2RosLV13pQCd2KQW91Iq4tQfr+yA2snvRX0BUuOv2gr/i1QPdzkpyeUl8KXPvygVhp3
pqByFWk3aMx8+WTqMJSlMENgHWy9/eeOXdH4jFDVTrL2EXs7sSud2m+zn3SzDPmqeDFxdGvKHcug
mIMCFw7g00apWKmffnobI9iKuixUmNY7G0UmJ4lIh25porIz7E4P8VJvbifBkUgPYxaHwrDWBebD
ohwhUP3ZF3JvCB0U1tkHRSEqHjN8ClytSg51Ym5JHT/uWE30yaXU2IH3y8S4Hw0WJTBAt6k/CLtn
p5JzPmvZaWc6bg1s1Ohm/U2QicHkAtjsCqG7+WiWwlNibZmFHMxqK0mo4Rq4FtuXHj5NcRhB9Zdn
+DXKXGNqHRo2d6JwiyMSVI804Sz9q10Hlm72TrXJgqrU90NucbwxhmaV5mcXv7spxFQfyiRf8XYZ
P6VwOZl583PmEWFX6xnfUud7O4TrrBRBGaI2+R3YonptL8HSEg5fxI40o7HfJLtn/DVs7/1MrSlr
rNxnRI6ifaEe1fa3vM8RS/4tAg+VCYLly8cXf6MXvkXqwZNN+nkCueiG6p2l9nzjLwd3t62qB7FG
Nc6rDMS8sXRt10mKGv1OELGmh5NPBp9ZrVcvUVxZ/PN9QNkgL4SB37KWqRMWD5yWiGF+1qJnoCFR
BUm7G3o0oj1RlSU9+juZ0iXxS2xRiv/X5i4F9LonP8fE2R6/ooHNvnwrKyftsaxvVgv9EEfPlZLa
4KHiWbM8ImX/u2ODZIPwydZgVzNH00uLlZEFKPGmK+F4wfNpY5xwMuBQsqTKNb9TVDjf+W05Rei3
mxa1XSbyUkZvQRthdcHLGFomXORR8+c1rwG42x8Z5G8dg3HrioqK8/wYNDyKWtKR3f5sAvK5lNIA
Dcb2kxN5NZ3Gq33lLqK6Jpv0ypxyI/7uyEkbB0QYw7z6/VL+wP1KELbBGPRkewBFJSo+5QpPhmPp
0zYsv2JKMCv3PfknYM2h2GZcca8+FArL0dHjNYAf6gYji4x1qydHEAwe9b9chKkeCLAchMtFtgAx
hs4cBDrd4N0x1XpTkD6E4jNKjsblP4klLi9rhynAA1cXJFgmBU85kCOMAETbUpS06P/VyXlaKN8J
gfuMo4nC4MJXYts4rdVWIIfa5PtZ/iO7Yu9mCnfWDsBk/0vcuVSx2gvNtIvavCEvA6gU4pou46kz
Q2Jh1G/P4V0iQjkLyuweVUp5ekkVVReg6plVLpWSA16Ag0JDvhFDIVZUiJy4udPNtvzFytzrizVi
x061MtOTJmxR7Sdz53rX6eCyN285FVcFigy+CV4DmFiu0nojRteMzMl5noht1NYTsmj8sxz4tZUw
tiqoIiTufr9cR1TTQ7rtGXzo7CxeFAaaiX6n5CRY+MkVFUWuyxC6FllSHOvmk2V+V1FzEaZn8fIW
pufcSZP84lO6Uc6PYK2N2gUMz2UwuJYh2gpjD/yegWbXccqEvc8Lam9VYJDP1swuaA/kKldKcXMb
xauk1kq+yLj0GnOa5nJNzTp0pSFGsNzTXs4PD+I8/E33EUwoQR2K6bkGT4adE2L8DIrdHkUSWNu9
sUzP2ErUA26IVPdXNZT+8V6rxR/9DCvWDOwuxPou1mYPsGD8Ii0YR9U3oQlV/nRnNfg5ZpoVRunn
vVagDe/JZ5k4hkFG47Xmw/DGeIG8WTkaauvSaSELXtEwSBn9/Cv4qD04FfN8kcWNE8LHpdyPXuph
KYfoQBu8TxdCpPUGUx6zFS2N0KSyJDyy9fa7AAz1QxVkL1bRqBqvjPGDjTrwLEz5UADu/0R1yD8J
7ls2gp+S3MVI2TJfuDEt0p08js8QE4hszjBZDyZjbUY+/5cscan/gJnM4IldKzf9LU4fWE88nt5D
y8SSQs5j0Z7Vj49Ocl3nsXh+8AaiaabF2VmfkwQnI5Mq39duWP6vN53LJS6L+CP9PddLOQGrmjc5
V6jYLyg5r/kC+3pbF4hJCwVB2Ji//Bdx+P9N9oNhO47plGTZIyq6iIw1kNpIgC5cYwfVqlIKTMfv
oStm57nHlZCqp1oEpUYYrJ2v4qp2WN0f67rQ9HMkZA7eq6atkAFGodhe97RQILI1da6qKnL9FBZr
xIhampcLhjUZJ19THxsqpydF4eXQfR0U245sjvAFhMH9HIjQB7AdVAZrLJy49D5/2xxMork4xOLb
dDoSa14j1yjIDB752oFjbEWCUmIYC2jWcH6AhEy9/01afslUZ+KMxzVt6cqp+oeZMaN9JXyWMo7g
BEXXXo9eSIacGMPFsrY4aenJjj4ClTcpjftBQTS0bJNnU1nMzd6Oqf2vjMeLMQStt3/FA8NTfKWT
/urkXm5Wb21QP5tb+oiBGoeyfCkzqIRz4dDtJnR7EpsgDKzxu9my//LjEnYwolawduy4SE5Q25pk
ViH8ppFJnNMia9xyp0WCWBrHt3tT88awq4zuszmnfqfIytUIJnqhIR+OATdVvlTShxA91cAEUrPR
6zOP+oOG8q5/ks7rM2BKFDW5AuFKyn15oW4Ji0tYQeTd8GifqoNjQJDpj9VhjDUPgRr46s02pSoh
bm5L2gPrp3e8VZEpbym/IfOHcXqPZrXKsoQnClVY0hpygJAWNpWSqm6uFWrbaT33fJhWznld7M0B
RBJTsJVhQNEMfbWn7T3GsEZUAli9wWA4Ah2qLxJZRYXvztutLrnIExnmWhx+lx/mi5ZpbDy8chYO
Eq4A7i95ULIo5CZStBNxviki+R3aniHkv/on5NmChltGxhYMuokFsg/KR8FvbVtnq6hTqGXvSBPY
3/nQZaWbqtTZuY/50vIZ7xWKerTaXFbF1/JW6conXx7pRETdZhknvxhrSggJV3QeiSzfOLAZMy8K
wN6c+INGjM8+HRs/a6xiY4mh6SXhXxnsau9MSEmamxGb+5zHPlRGDu9X6mZc5mS4O3An4OGqTODG
N8VrdukXzAKzoho0SPPV/9QUU2EUYRvjhAtGo99pjOBbH/Sqo77Weaq+CCY+xulxp9ruExy5p/OA
RNcoEqaL6HWMCE4P0H5BDt1NUgiFfNIbFd9JiDac+WDyztU959IY0zIYA69T0f1mjvHTlzd6AfTh
maRdaXvyrRf3TOmQ25Dpm4lPdLC6Sphbxvy28BHnG4oZM2kjxGRtOKbLyBDRBrapEN4l7D5IRsFX
EJO1FbwGza4i0PVGx+jwMBObv7DT7+WXUpjbjg3XsQ9WHjN01dX7x8J1IVBIryzZiXK4BV8XuJXe
uZCny/mlUJ4Ie32G/tTV86P0ZxV2p1YukaMntcpPWLO0AGHeKWnTNRkk4oUt8MUo1LlcrDtlUB4a
5+RnxLA0LzgwFAJzc/UUBVFfnd4vaSPTDLyKBHZPZ0xbWsZ0NvGPBx37c3WAEP6qAyRj1qyEkx22
aGAdFpmZfaC2MFHHuQKYouPihaS2y+AvdBzq+KNO1Ti3lGyvPHBKEiInf7qi44H2+s6kfmBGvkpV
hsao8re7+SCNzn4bp5/4e5LItRAKVDtaX051CSGQb/5SzjR8Ye2VBRDPreOfmxO5N9MxHnpm1Vtp
4cTWuJNUU6NmYi7uCkrO5EFaDqajkvRW2M6w90meyIodR7wXvFQPjl0Yf7hKFcUWI9gRyolHovdd
ZNqWFaoWeOtLxE1szeTUtD9LXj+1jhaFZ96gsUYJvPK19+qSvG70yT2tsa43xCpZHyQKnkEbOb9y
jQcSe/RdMNo2+9gE9RhbjUTbfXwplxdfNCFj5/F506V7z6frr5U0uJgd1k9C9GPnCB8wGwWwrqvo
2l1HHhYqTzBcdwA7PHZQsSend8KnTkvLIZhhfkRVmf6J1+2mD+QXRRB9wcFB6GrwIOpxGqr7e3ME
o3ADGbev9fKbK1qzihU2Xe3E84RLft7sqtFK1MP3LEgK9OeDxMOPcKn0y5lNgGSWbfS+WaYxYunx
hnt11Njt6A/pSbxJhPQWfpe6i3Ul64gGRmp4ja4lliUMV1t6GTTBVTnCLJDP7thrtf4yUAuOgnyo
PqW0LYVqjODDatNmWQZABmy3x9lLvb/DIZNeVGBtklDsXFnKUP75kyzBrNIL/P4qcWrss5rvNh0K
RXKTelG6ybAOUNYPENixGaFCt0sGcUkcQwVfgmLHNHLxqRwcFgDHN7ZcZK5yqYkKZdugjrl61ivR
K3X8BxBF0pn78Rr4YzJB4bVd9sNGYuO2QA15364gMimqJWhnmCDB/cKfFwghYh9/xGsjGWU9Hk0L
tutYJREuiYkj5am+a9SHi25l/WANwqF94MQWblvFWDa/INpWBJy8dgMPlgNb3yJIX7UhpZu4uG1K
gooIqde+2s20ocdxjQFlF9/CKC6PCeKY6l5Y/gZ3FFoV64GoSY81CD2lJRL9OAAI624WChTYvWOm
u5OSiP6J7M3FVOj94ypJheZMVK41SSYOqoa0odT/pifK+v0IzDbBkQpDQEPIbZrGyajx3tOTHUjv
S1F2JAPkP+5mA6exS8hXL5Y1CCvvKOkgaKiwi/77aMlAtD6Qpakr3pUIBLOUPWAp24oVZTwsnJcy
FkwKOb13o3rFePGGDTnWqKW08E4j9fkehem+3C8ycLGUyl4I9Qro9JMzA27EMQ5lSFNFmzPYbKTP
wn/aqxXG8XIKLfJ/1Gr5GSuIJWkoTeEL6isjI0fLQAdU4P/dVGavrZ+WLIFYVYiLxY60uxWk5dNK
Es9khCf3X6QmClK0yXDGeOHZ4zZJLzMvk4CgnZRFYyfyfK0zk7Jcohd+YQ4DALHTtpjntCHEj7+6
o11s6qXh0Uuh2u5CmK1/A6bkMhh26zuWK19TYxvtiOOwpMVwWx1FajIq8XqKNAYlx0IiVcPhWIZW
KqRksTl/wHwBDSpfRUsBEyzw3gu2hRbLB2pCvZeAOlJyRrSNRVLwETFuSNZIbiM/SGgQ7FfGyVr0
I7e66x5iH1ICq46KyLcAnahfXkHZ0m6rtO6BzI39UlwUhR+URGOLXoiLnEti4pfIEtmLz3/RGEVm
ogcQgNWLIfxhNYUwEHEOXJqG1Pv34zSCx/WGJ4KVpsRrL7GKL2Kmj5uGaFf11M7BM5b5kUjF/Cno
vXJI+5JMxsPy2HQE751C7WsEXJIF+XgzjKcNhunsIWPMRhPTAZ1KrWJc/y1NK8fDYAsR1g/jtj3J
8fiBPxylK+OA4NjM2MwLYnT/VmI5SpuHv3ugLUisPJmd9CjpgtR4CSqJevD5tsFIPCpfYj5Szl6g
O/csVeKbY3x8vljJwlIYRBBbxfgankCfyPXhdnCOKjggvimqfYryg5yOiRxI5nHKMKBFvt0+Uebd
kFFry1WW1kdYO8Grq+attnsHzc5KOo6cNtVKEXZd6MVvps3lHhF8TJpLQphZhpPe3lk9W4a4wpBk
PSyLHmHCUPWTDrLMjpoLq3H/g7bMCodA8g6s3ZdKqHgUmsZ3ihP18+A4g0VWrZG6SG+Mqd+0h3w+
1A8SdSQj3GQxtWyWRPceqdFm7CGVpW27FKgYj4NLsgkIX1qrwh57nzFrdTiE1rPN+kz66YPqhYcq
y6jsoytnRqHrg7qY/e+l3SgTbEcuX8z+gRzwBrsCmoWgf4a4iHzQ5b3tthKTaytXCCpSvOvH9/bO
awJECYcPIOHmyFlR9vJfDVFE4mB33Wr3+WDu4XcJhnkbuIz/gq775qMCviFe5xQRZE8KjKC0P+/r
7b+AQCOxIetuIFzbOdRH9A8/FTTeOgwSIPh0JRHPEHFDk5TXGzw70kWACQmq4X2MeAgS4IJc35rQ
fQWrfiy+yL+XAXPWuMBL1Sa+tdmPcMV9GFoYmZ+nP+OSnRWr8HkiXPi6RrEsed0ovge/hzNXz6eV
P0wTx1+EgI9no1qVXgEGzcINnrGbc9JA85m3nbzck/SzrzdwlZowO9YqmIMjyAATY0m+GL4c35vG
gcXLtJLkEEzWuwQsg6U0Fn6/C3j5UKV91efvCXQA+/uX2QIyOGecpWHilvDo2G9ayoUmOhQrqDVw
Qlu6uYUYW4rfLeqLBXs9En6NsO2NtkIFLtwPldOBP6Er0G90fhGvHOguN1BgYVRWAZobL/519xAO
Qg6y5/1GQFs7gtF/XHZpFtOWEtX1siD9vj/cBBXWorjAGlKjgL0CSkeQXVtpjqzRPkbK7fbczLZD
wi40egB/5EPGdmQiC9RT3uh+vwrIdlSNc/d5PNWUPa1JH63vtKrCBTmgWcFkxWJ1XBv2ibg6Ulff
3w5+2KB+I9GTWUPZC8lEQv7MqjLLJxV1QUgBpFcI3NYpz//jytCU+gnQIC8T5EY0aNaLuOdb0ZTE
tV/FV32Azdr+3V6Jjlk6aVrHimY17iH681jlQeiPGykWNkVR+lT6mxW8/56iSprPnAdR1htRoTb7
QcjiH6+4/x8i5ZURAqJYa+CtsEXoXIUF2Pksbyoqu8UDSQ3E0983XjwDDwlTu8MsVSvNXzktCjxv
wupUaAgSTt5Oag9iVty03ENhkoSkfp3SkPTeTTXyKpl/KmnxtLUWocc8sdGgenUsz4NZYCdfekqi
gOq91BxB2KBUCPx57FrNDNR+6Q4uRgrzDDJ4VAr1evoKQVK5UXcXv/CwgxciPzvsjSP/MKiEa6kl
9/sM5cNI+AcjilWpyRj6gUo3pxbdkspgqCbjCMQ/S/EzqNv1cw7H9j53AOClST+aEBstRJmiMIKw
rPfTuQeOiW/VaK3cnR7Prj6s2SgiD61l9g0AvpiSMMiviuc2tUGikCWj0WCd8vTczRIvavRM73Z4
VediNzsL0kUlhILcJvgjnq2PvRrHVgK3RDzR36IaVsg8dtdYXQk11R7anHkKuxvCl3TlPfLhqsFS
8A+gZPxzFQ1lkV1rV6wTWBx9uX39+je/FoLUQmHmu8mzSOWkMvcUIoPj6lfSqw8x8TUE/LuTQjk7
Nu0gHJcidnlg5+G53JumTTlkJR/GzqRVAPqOfwuuJZVdVjPY6cCd+WX073FZhNmel9Ttx2hv4sTd
z1QbMAzKlBR1RvTqTkRv8a6vhODn1guJmdIK5fI2//tB76C7bGu+8fDhYlF/zJjxcO7dnu2/fEt6
00LkYAgz86bEqmXjZJjKAm6MremLATMOShrIe1XJQIC+OJVI7uqyiT8BLehtDxhZD2/+IquB+Dey
EiD3imyzkktOZNsKcWrqVyyd09xNkRiOEQyMALIanubw5vZwvNEc+LZYesh7craY4dxcaJ3Iifin
mpoqTiAN4Ep0VW6RiynAKrOJLZBIQ8F3Rj3qILNh9RJRMR34eNT5hitdGoxfY0LJPGTZbN+9A8ye
R7KpgtWAYTAYZFYs2tFp1D5xhwBUlw55Dfy/k4Ih73xl6UKjvi/alZDMhpz8wYEKmxExq//1mEpU
/HM7Dh72Cq9BCS3xlK1Jzbe2zeXvzhRgOdEfrJ3MKYizSC4Ll7VZ5/5fNdnsLhVg7js73QuQaKzu
vy4TDLsTzGXDbavfJfIEX88cqkohqhW4mIrFEh6lnaQ2x69fSjqM8X6TvZXnH6TXZqkh//SwtOsa
p1h6K83u3BOlKAbC+At8TquIbKmpfHGfEilsZ4iyPxTILQwhi/Lva97NlkehF1uyIG0yY61pGkeV
n82X0OmEfqOP6knKLHp41dBRR6uj8rrRvqLHiKuhWsLeK02PT0mrBikUKkgcV6+Xhe7xd0j3EfIX
3pUpHZvVe0kMkNI9yeIZ4xA7IXRDEl6lFB7Nd3m+LLwLmg3ZrPns1pTucw4DbgdEZf41Vm43FoOm
Swk6kXOOlrZN8mmu8T0PFoD/LJWFnE0bHiRnUZekLewxNRMyfbqOUHktW/EJlJqFpMSX0wy052eV
N5DT+iG8Egfm+aBHNfngmvtkvjSXI/NQU2o1z2lFuyRBW/+AExyZ/7U/7RRYgr5sLgOJ99qrUmC7
t0zTr6E03fbsAYuvtcBwZSb2Q+BtIxChblJDAQjCWuPtroMs/YjnqawDPQDa3pkPgvjiQhh5MoLU
IofC2QcTgpGR+qNcq71hIAci48kJuge9Omus7HEQTGltqPiYnfE/Bg7FpHMf3qFOPoYBWnzpR8/e
JWPqG9FzQrCGFiEs8KGqkYpzhARYpkDxrTM8D+xZmgEtEdiYZTmvYpg9+KqcHmVkd0A21mjk5HVc
n+TVAXw3p0X1gai7C3icz1O4GX21pdtl0cAlkGrdE1iqspTwGlvj+gHpeJvJuLjs5hvCMPK5L4qG
hkKal2LoeMQMmg/nyRo1LTexuufYfzG5WTaPYcaxn+9l2Wq/rCd/ySHWGeu9J6uZk8g0YS2sJecQ
QvPsZFG8GYzGKDDeRH1hbgVvO8xgif/IV8BEgQKK/t1ZCxaXdaXzHaXFu/xIU4sX0PLbkSrg+QMK
PsJlLVPgRzHbTBgQhIG+2Rw023wOelcyj+bQ2tp1Gwr0IJoOX9CZBE2KTTFfxdr7AS/lAwKsxLzY
R8ZxpWx1WYSH05gXKD491T8rw0f2oOJFV/3LXPihlZKqD7hXv2Yz9L02ai6Z8NHIH5wXn+E6xwg+
vZm63l4ckbEqIzyKbWI78CWQb96fb+H0Ea/LN2pFJJcXZR+v67o40vSgJdqeOdKBtn5pE1t4qPqT
wCat2d+qlg5OpqR/upVK/P1K/L8dG31EdcdhkxfrWDe8q48U8nazxyL7gm11b4nEwVQ8ABewbQKo
ZPMyMEmTwBDCqTxg7fQvN4HENk4USfMmdvReyQoGDx7oqjmNdIy+S9mkHs53LvfeM1RqjYPjyMPd
rIz7bpMZoHAu1OfNHKKXQTmKeFE8Z3Iv+zmdS2dFTGaR/4BfZ2HSy85aGk9AmVwN6GeFybINdrX7
DfX94WyBggZ00jcIuB28j6WrHpIBm478suGXsckK9cTpUVJUlm+CDR6Om+Pat/GdG75asemCgqaE
A1zJguhYRq542FTUtZ9QzqcIyw66eaOQ7Wq+FWb7kD72hEy4V/v0yDsr2VbdJ+mIbwJXcNBNXzh4
HTjGdlr07FmQZTaa2kEakwacmKpA5OrrC4lfGbTDnJ0wxzbKnDFR0H64JAhTJ5l0gPrlwQnpjjI3
cvQetMJ8wpYI1Uew8kDMxYvdyA1yQ8bLBZHGl1IjPJZj71rweOXaxarBaxEL5LusOjMfVPtQRG6I
Yx1QeaMuMqRG1g8exDtnvANGCHQCxYLSPKpt8tFM+zkeTvF4tBqHULKhosBCoyxILw4f96qaOONZ
8GSiJHDLaiw1NbLPo+VKslCM/BjerGpUn1DRE7CjF5qZrJYnh2/8nyl71/nZPiHATOeDA5u0chBj
v7jgOYhqk3klFGVHRE3J+j6XyWiTqcOGOVX855s8VZ8R4Ij8HcGuajbDMJ3mIUQXomVx73M5XFjR
AX0ELtZiQAQ9kNUt5GwJ0pTDnvMGDWt+6dj74JzJdsCtJVaycev9PQxkvToK6J48YL1H1IEYm9v9
Ki3BX46Sb3OXr5BYzfxZLiarZZq+45QIDbaeLDhT+iHwUaEDJQrLFT/0sC4qBEexzSzERIZdgwLc
XDPKuQJbMAYKhX+MvkbBixN5i6+1iLrSZt+Y3wXd9C9hEZQRydHgtQot/HObE1U6zXRD/LaWoDLV
PG66h/XsFTwzYbGCba4eHnaWWPEhv9eU9UDFNlpl3HE/G297e6SkQqNcBHTbCT39pu24g3iBPQAB
Cz2jjnq9f0Ir4thSf8OoOvGtmo9ORF47jV2n1RuFzdGFDt1i/C2v342qUzhrWLYbr0c2WJDGFLiD
/3jSgfkfuBQgsonLpNJ+6kHYrrRLYWglWF/dAl3fuNYk6UgbOOGhYUqpON0EJaqz1srOO0HWGUGg
bngnczvlDVXQFcl2vhDXMlwiAUpSM42ljUCdUN7YCrha9ImcKVvsvrVj3BN90Mp23/lXUmzMX7U1
Q+3IVSEmUX0sdaFU1w1FFkezm0LvdjQl0VZfh7vtvxVzn5hIY2Wk2ptzm7OG0xQ4th3PPBxUhDyB
F6XQL7xgqk/TvBW4zsQ4vVUJcyjcSQCzyeRtWSw/1JjGg5PhHWoxv2OBZwXbp3i1L8Lhw83g9ez4
RmrpE+kClGORGadACiFUfeTvJfZjyyuVfBTF9G9WehrtULehh31eBfIkuct7dfO1Avgr4MaIDiJr
+MQn+tjNlBDVGqCBylQNNwoFI8hO6zZ3zb4T47IXgO5V1/ubNtokAw6hZAa5lQF4vJ25TzNai++S
z+4gASnhiI0x6lCPC2muogphm9cbwkCzzMjJ6EaM7wnO60bs4ACMaxFQI+8bt9vYs3Vn3MvfWzZI
agzaYXSH9LkdyOqtNNF4MUlyccmx7RBNSW4Jx9XrYt5wWvhs/OU6NHG0+wLJEEw4h8iYtpYIKX09
AziDqH5Gw9ntURz7yPA+msZ1RErSaIf26JtQCPMYJe1+ekiK9dmC5tS3G7D+XQZfoDeLvqzU2yqs
pHMXIvM0gJ3fWYxLgg272FZSvo2gnRPjnwxQCciRYNZdQJL1oQI5XUR5PM7SfmY5k5OcImdsi6EB
gRDujOFuvzXCzlshNuPn6U5c+fuya6YGe+j2hGymiNPfeQ2WN0/NWsnL3Kjeydcw1w0qcmkisYxH
nHSNXRt0vUE+cq/Cd2i6s+ObaDwTK9udQ8bkSApqxYEKr9wj0fKc6LqPkDV7sN8hqjZnbpge1v0A
CKAYrfmhGmBqOTyVBSUPA5ZMWrrOtfQWiC+PG0wNx2abUuEJkdFGzHHMGGrO0SbaMWq84b65Tvqz
iy65kpXLrKfI84j8kiyucPosvWYVhgVlmHgBqoaD3knr4/fbWsppN920ZFpfm+xrFq8Sn78ZBFw9
DtuEWQD4buwZkgPJt3v/KDC8WJ4mNxaw5nveGiVxNDzo0Wg3+Kcs0DDOawsbct8ifnN4lzRznRgB
EISk7Vve/h8NmlWKhLmHAUvWhh5w5qcLITE3HCwTZMuVoL6VGQz/ftAS7sSV6s2fU4bw9SAwujw5
2f3G/W7I9QpPXsSkFQD4QONP1ssOKobI3wVhCm2ldjfqqpHTYW3LLqRUghVT4YJicx7bcytnLBPl
1sOvSEHTvRWT+OoUgDp5iC8+04vW1KUMR156TRckyXfd35HZar2vs2Fx/02SpSyxE68pJWcceE3x
TKCBH7dRq+JOJiG/Pnqledg9ku96RjKHTInxkwQbPPDIn6wrMPqP6rzvx7moxVDgzknWFoGKnAnd
Vf/fPMWs/jxSSrYjh8yJ/RsEDwIAqbiZwaygF2ktNTq+FFPeNpDg5rXI0zEMEu31K1X3Vd0ua592
HG4dEM2hipfKOy7HZq12NmxV8cpMDBd3ieB+wGw1BuYiY97HQdsPvLqt89YiLQDzHsyWuC/kMgHJ
l1zw68VRfDhu+dtiWgDxHwgnttQD1aN21t8vqGUG8MDZ0H96lLkpqDaVSndiUK/ZXys2zqvnYmKm
73+MBWMJLW7+m+GQRJDa8vcJG21qslq46kyb9HyK4q1n9MwDKcZ2GJiFthhzNEubHNd2yi6r5Ezl
3pO+7WdKTCAf7KXLKvTdUoTGo0qfyZwSUvXs3nXzcLMHfef7lKF7McsFpD1uGS529n5ZUKrPs7qi
2nMbmMha6JRFcUJO+HnTFuh0/q0P65rJyhYYd0xGp+8E3LAR6f4bVoyqCixChMZVNdOP0NWHS9X1
XTlp930j8LRzIZIbqbjvr8LWEG33yFKDSWQV/Qv6BR3zPPzsngaT9ViJIZnVxMz8HOFXKIfh7Oo1
LBjZFqI9eIEfjo1/B584hpa7hXVWUq3WCmCZjERnbpquHVpCx7Gu1VJaVWx2wcq5ZBpV3LycmM1A
i973CvQb24gcw5JG6znVtqYZdn3tgHqDbZ6HwvrZ65tFSJEzyaGQj5iLe5+oEiaxICf3xeOz0gU/
qgQLMYQ4u790+M8FBCAEEsM6QK7DMyPw6gFKiPZJV3z1eoUByNWyno/sJrKgON5ZtE0G8WhQA0hQ
vBYaJzL13TRwPX5PK1HXj+Kz64Wr4LhHOLm+6BqwYAjWaCSyCe810haERqtZ+OqVsxbzTiKC6Wzg
boNnRbv+W40UXYW+wu/PWdJcRW4AmGtRpfJtBxKtBWdD+5J5btC9PcFWQOfOnfQwf9dpJcoiCIya
iRS//fjeu/GDGLooQO53j0zhIckd0ad8rmUjIENPs78yJf8uuUoupbSKvSozVgiAB6a1xYVnM7P6
a9/nvdRoUaGfpLSKckQlm5Vea3d+w2WhERnuDDIMMAep5/OqRUkmSKef55olYS1JL/x4yzLvihfU
kSRtSp9ysquOhhNV1cXfwI/r7d3v91K4qji+afyPue24Vuv8i1x9pnRKeDnIYlAmxxKMPq8Tbiyg
4DyPzNP0VdfI8M0Hq6wBVEkQlgPqUlrZ2h3yMxR5hcHe3VLGZwV1Y2z4UHPfTlK6wm06S0bvmNba
qS5V1AgtpWf2zLAns8oSIy1iyAMMcmusgmWM21pRPwRWRguyRumLlHEkzQjN5rlOW/wyI5LhfX3J
La7UDWEsYC7jL2Ju5talaELJui/j/2M4T5ogQOagCU5u3P58nkd8gb5V/HyV6w3jC0fkZ54p/8zv
oYDkieExtU586k/fwXv5iyrYlds8BQQssAZscVoU7YYTaKyghuFytOIHjsnnubvDtwNM+cb8+kuT
xYkIdOD7kXuepqijuAJOGE64omJZKsYy4fKE4DKaD/iMfp1zt478Ao1l9J7o0wTbk0abK7bcRyzw
moKo3iTsQjJ7XDq+L6fki6+eEfMwIOZ8/dVWZ30r2Sdmo+570VCCSFX3bFRKH7S7dMXDcDnFBeZe
ciLi/N57hDQ3QLPVTYZ592cRndZ92dEJYVpNWclrJeIFhNPbXx5f080rp/uujMCVNuQXypWug1D/
ZLxxbKlXrvuxXxMzIOXJedybA6n6gSzldkqR9/pCxuq7iGBdntZBIuLP/IVnKhQ+twsiBDOfzhdU
HwfrWdZpwtP4VqqHxocB4VhOB8SBAh+eDhLaLNqgrfygokpTl+e9qgZCfb5lS/FIjtRECiVTdzIv
o5lT9c/S/gMKv7KCS7824pe46oneJJlHTOdx5GLYmkVEhr9G9A5Nyb7o4/OPDFG94ZyYcBC6ONRr
BP/hRjUXJVaY6xZQ/CpNWGaHbL7DG04vrYIYKDWBjD/Yn69cflDi2sX1Rhf1etTYvWJec4Ae/hJt
Qlom49PaDMC35W0dutbkD9kp4F6TxI142hZFxjqDR1KxkusoBToin+hsTC4PnvwTm0ny2uzBRa6Z
2PvYIzuROcts30lB0h0cL8ShLFLR0rSMbbgLwPVzyJqBYpLySJpWb6JRGhWSY6r54K+/iIF4l11y
NiYlNn3YasRI835l8g5mvaL6RY5tzh459B2hqD2GLAT4he5ZLcOak3J76kijP/WtCPBUvkgeiNum
YvAAmHmMZPPN2id4D7q9fkeMnW9xcksHvc9SCWDEnW7ZyBZuJnyN2keBSpYlkMV/C+w0mu2Qd8LQ
tK9oV5KK/zoevBbvfYc4uQs0GJzSjzpK68vutqabQZVVQVSrSpmO0vk3JDiNuhGCdH3fWH6SdMaF
qFLhgUyy2Lun5BrnAn1rJWPF9eaPCsSimzbYLg2jzQLQXNpxQe8K2fWfPqkq/9aig8iO32415UO0
K3MQ9D7Fx0LjGb6yTwbShWObdQl12eTK5PzeAyzh83Td1dVtIB6duUV/6TpeeZoJ94DQ/pFkBQEZ
2dSm5TGSPS/N++Mso71I7zuuAg7FMzuwa6RUXK+3gMgpqQ0zl2QDZvEp11hiFAZ81YaILJLFiezI
BgXLbLxnXBhQr6xnDFWu+ZDIJmYMa4/XGJ1/SObh3G9ATpSC13I+dqOZJnJstXyB2GDNvbx7+HgN
hlatoMsfGm++ph+6u65fCqvJ7j4/+Q+JPq4FM/dLhlUl22l07LYjs6cz7C4XN/yjXhX9HF+FFWL9
RSjGdNI0onmidZn1LGhCl8ayZXTsYqhaFaCndfkMf4Z2FL+CQFNoPEsK5F9M0ES+4PiGSe5k7SFh
cpxIJUslGFcFhPMtwJteVnEq2v+KkdlvFZcZU3xhHnp9Fx3R5RXey9ytFVpkZkjuWXdRJlof7K8R
F6JGAOy0H6M+tI9L0+srgKj8dTzJWqFZAzCgzbZWbEK4yHQMcGtMGI30lUrosunV3fvkw8jY9Q9G
R7TMSQKET0VMl6KVsEBfQOVuuYM6Oqo122YToWHtjVpq93sM9TSUVXIW/z4JJaztsEAPRjWEA81c
Xcx0x7wI6O77vH88+ePvipYGV4NIZMzgiv+1t3Z4x2lk/hpv4/naqr7a7Ox06xZhvjAXEtwF71tr
l2uiWlByQBgUgDBmMV/5PVNXN6Vn5jtR6CUhMRpzF3qMP8p7cn4/3sugvrO63THN6cSlBdnKJAGp
9EWgluHyiHu6d6TwZOJ5ixslh5v8O5yHuaxJUez/gNZKpMYYXGYbujNIXz/2FTd96ucAqFVwSryK
maN/4zYY3AeFqSc9VuO3CsFhBvin+3HCPtnm7jMywpJM/yfx5RUf8BtkYg6yBjZ2KTU664jsJaSq
CPhVblE+bEdJJTY/zOAGIf6Gi6uge59qkInyMOVBdo5XvzTrZ5V3MBDwPlycI6T9SBKaSYt5MAth
KVsDxo56Y/BBNxLGuD4dQNcSM84wymF8fT+fyEKIDJ3o44dHAm1ODhEd0+E59ELrsC80h6KD472G
z9xw7wz5G3Ek+yhhCKIqi7KFPIL0I1hg3Uu1/EoJe5YmNY3pLqfEooU9m5XoIK9ejGAgxYr/GMra
TXxOBZ48QLr5r72X3r6ZKUyxme54SrqFHmAofX0ZYHG/oNJyRAfrGyWQIUNqc2Kk9q7J1ppHv+Ax
2OwPMKGzSRfeA7Oc2FZljrYlnK+mI1KNMuvSjGKuzybkQJ9qweRa8sHa9lCCrmAdwpUPMEtQpUX1
TS1rj79QVG+bM616MFhIvsQgF50HfHxn29A5GNL+hSIDLZHhI5kCYChB0wO0rgslPGWX0eL7oBvK
jMZKYBtEaDcIoFtJiSom/jQiXRx/gC5SlPTjoe3UK+618XYCA+TVTzac9KRfS/U/kQBaMjTAz7Gk
yLympXeIW+1Wx2+malZ4Ai0wjZDIRoWQfOav2D7lt6euoq5Too7s6sYVx8jXMQnbCigkSbJ3TT1A
zl7I/Ynojws3fJTQAsTOZMOt/rP8bLni5c4ozRC4ClU+b7piErOY6OHKMFmjXnR0nLEO8w0/nmMo
eWEsCIfE7h0TUsmYQ7T2vClEH8zFR939qyepCe7HP3X9EFK5HrqysJScls0JymFD6mkpqRCGjFEf
6QL5RwXJLynsWZqd6fLv4GaSGPBwCOocGeLIPkSdNFx5ZM1xZbWjpS43Vaz6qC1SdDbG7upyBhc1
ic/HfdhkRD+8MFHe4b3mr4gi0kNzjnI9DsyzyC259iC/JjtecuLfmrp80U0wjrzHmNUMGQ9IHRno
w//qHK1oV7sGroyu3nf1wEZPGyxaLg+ExfK+9M3aEKgDKAusSUGpnDglkFKIQJPPWr6qAliU409+
6x+uqsoZ8pRkXtOmjvJs0FVzvHwk3lnAZFPPmeV74aEtpEN4n9en6Bb8w5zOYMJASl8Z55ylTKcY
wFaFRryUPydMi1RuELwSxkLHekflnnXlwVeA4czmK/SO2jFwtXLhhGLni4cyQ6TqAoF1KuDqc2X7
E/SAliSGu3cB60bovVEac7+od5uYTM4iCMUTCWpHMSX8RmDsS0mUE+G8cV03x1FHW0yLyYE8eqDS
Hq+O9ddunk957wh3TCFDi/7T6LrkmOp4F7XjfztihCqmYHDhD8k2oxe8EJauprsHprLFjzAtrp7h
UnXDz6g0DO+4cMzqGm/G8tqV8ZS0C3thwX4oLMs6na1C9LNZpmuYNNj6HeKFOhCkRQW5qHwjdzoj
JWEeZQsIb38yZbOlG5Zp2S/m8MuPT8nem3glB+2OMkLIQ1K4TV5tYTbJZRkUGhX5VWffU0ELIXHU
exvaIjfNSKiqkBI2DlaPJX/iQXNjRm7KYonJmbVS8FZ9ST0t9Rd+9777pQbGoN66N50vO+le2MHX
GF2pY1W9CpPY49QE3xJvF7N/vr/C+4pOYqEp/ysBxCaEKvcZIVNCz+b8i07+jz5eZZzsJlYQvuWm
c5wK0UU27XPShSVBDvfX6AVyfdHXbT+KivAWLFCaQTlXA+QFUBMhtZU8/m2y3gKv+ukS//y1tNxm
PNYi5Sb5Cz9Lpl7v6TLq8rhVDcycWBwRbHRScoPUmq1F3uHOKVbbRssw03fAsax+HwAfKxI8BdrD
MMmusG/XoihD0cv0ZcOfuwHIs8frv6M6BqXXiP1R9ORGXWD+Lc4QfUsZbMSaSlk8sPPIwYJ5WNGl
KkUQwa/IRWSBAky1rmI1t7KXm8V+uBcpBuOhdDNOeLUUDQasc3yyh7uSrNtj8X1KURS+lecdEseS
iBe3O/T9nkAvWHuawLRT5VjpWxSc6C/qmfz4TzqSTXPcfFfIZLYYEEFnnOxWpGk/JosKsbpgcIUW
X90XTM5h/677XvwcayN0VhSDeMUExs7/KsRvCWpsuagaA0FtBQ5kx02elTPRsT7SchsZn8yx2wGZ
9gUqcQmxUFDxiJCYvVrvGgz2PX2Q+bs1Rxmi9Ekrffcw3AZRjfTF4t23hCHVActZ4rP37BwfYP/u
P+60ntn1Z48oGu+QlozER1ZW7aZlEP2/QTlMMaCD1M8cZ8IkKrVBousq5iaQH93vtecJBOU0xoP1
2dJty88OGgDaPdsuYkkvN8M52Xrba5yEueOTCNNITyGhQlZt3KvqzYS9NEI6qVc//hNkESTqAfG2
cXqx/vFEbt1qeIVclNAggcNSIOVErxj6k7F7P9IB1IQTeV/gS9F2AYNvzD+1Wwi9xV25Np22F5tu
nn4INBug1duVBBCa25NeE+DDzvYyZaH2dPv+JCOfkZrDRWx1m/KuhKp3WfScGznGWm87BEkPFn4N
8j4D9d7Wal9OS54WQyTH/QTmge1Upj+uG9dAl5nTgO2FG220uwEq2KlTWkHao8+2ORs4sGsq3bQ+
BCaa7ZQl926ZZT3smGpAIwX7U2JN5efQH3ec/v5V6MxxZ8tO4Jm5xMxmCjMNFe0U8ix4Qnhgocni
eSFJMDJ23mZdDfH6zZJ/tJbNEkG6NPTPXvxHBtaziM/YmiWF2sToBrxA6eoOBoWDkPytheNVPOvM
2L+qRoSeul3uV3+jQ0yzSl8Ojmy4Kj4vImBi5lwNTPZ9x9dVJTqRixcdrpuaTJLAORAgbAnhDBfN
/tCMysK3gggsjpFWdX0RVKlrRNXhzeiGWZYtej73H5bSmZ26gWZLEnQvts3ZZlPRd7A1dmDpxHzW
EozJZm7wtEgnuBnfc2Lwchzf2SM67kQhvb+K7FrY84AnfMhxXhP2xfFlIKqrq7A8b3lLNifnl4SM
We5KJXQrXFyui4yA/euXAH2Eeofj7XaMNYP5TpuhQYHti+JHkTnkYPFA8xBPygxPjRZxuQxEXKYG
b3Kf5K+M91AsbTufafAlzRy/ZPNxdWOEvTtNm74cZnBw5QYoFRGU7Q6QNiTqdV+SlTP4N6XpExX9
h5MHPXcSkzJgmOqmlDnGi8GquvpVJ96aNqRL5WTSJHrgh+00QQdb5V7xxKM5q1areIzqPw+l6fGQ
SbljXaKP7J4RU+l3OPGKDbW2zDr7r37UR7BB6iXURRlPVvRJdVpDBR5vRkqDzDkH+U7SjwWEhwzT
MvXvuxQaRtMQ9Fabc1NWXT0OXtesp+GXmOyVT87oyrk5Xz+quX12JKrltKbzpgGpiNU/+lCz00Ul
q4/aTnvVxfhzPyICbK2qqHfDiBye2E99a41KrrgcxExX/4cFDLFs3vtnPzo7TpG4EXcDnz3x0vO4
GqDst6qGo5myfZ61o6rxZZ2Wi1t9dxUOL+6CSFxOPzHXwzsBF+1j75/KOE4RF9s0lYWZmjTHL/hc
5vJZAFMcpCVLG63RymGzZJ/4SsVHXlY0accwvp88Az+Phi55hHZ0TBFBjuxqE4kBR27w0Ec2iA/p
dKyFFspxWm0w/wVLSHUHjB+xR/sr7mdeue+wim97AGflF2CD0oyMQCZAlo85x4/f7OnQ6wHUikel
cRplh9P4n34CsQVwbox3gsWlXjGFQT6xxP1JbV6y1pEZLBNX1x/V+GqWNwRhxgxK620sy8lQusDK
U688Q4lGFZdT4UWDD3TxeGJKFre3EGLjZ9JUFUyX+C+qmpZtuDYGqwZpBQzdeTjal/NxrlPiTmQP
qgVKKogt3ASNIYGjt52sPE9Kfhbx9OAXY1+1COqCaKGTdVs9YJMObRwJn2WUFwFwOkx1NVkhtNHM
neUjFW71VUF4OYILfmslKuiZMiryfGzRY+/mgaR7UoMYXj+Jzu1OaVb9HExXZvpQIWVIfSOIzYnv
KmH2d383AfpobiNDoP7MTzYM4I+xR/ZttbBhQNF0lHFGEoC7AgsidXxxW/KihyKVX2tjVhN/OmPS
JBNnXKsk5KxbcqGkxpe6r1I8HXGAhFbWkf8Ihfns65beE016sGnCPLw2MBXcRce1IFG6CM69S9pf
ygEpWwEqXnn0xfE4KUXXRA96Hjm56gPc+Ybd61WfGb0vZ7zwUj68Uthuk8/VIOPy2hj8QJqF6CEs
bmVcQU53bfvcR08QXYMHaUVijKYTb6MiXQkq24jGlvao70k+mOEz1h9SiBcLeFSYgLNDL7g/kHwl
fNnU1MWZI4X07aDDlcKJZXHUQtskw6+ocNOx3gjBGc8nQbT5rB956xV/DWGmAvdLguI2TOIdFDD9
S18PR7TdaNNIqNMgoyffDNSz98VgolkNrs++uAxD/Ukd9K+lzXxNJZhPHtyCFVXvPreAzhr5tLlr
p7AGs89KUblmhXb5gap/M9NbGfd382UydYZN1GFCFrmv17S+vFWzQQ6ueGqNMQkbUXleYRnDBqV9
TvkzP9fVAVpnba2U5RvCS3Ks6wxtO7PrQrc6rlQwPprVAgSBuRcFGUk15Wg+FPrEM0sPjrvvv0p7
D25VH3h7UZughJ2bErR3yZaJemZK9e2OQoF0Az2QsMBO9VST4C76P84Ngt/EOhaHtUQE/TUG6YxP
Nps7ICwBxqeeb3EOjxG2umrwrwCo42JLeTFwFd6korylMx2wnnla3i4PpVD19HznO2woABjwQbZZ
pd8F++jG/6/gc6g06P24CS17n4Un0A7RuI/HIxEPM+cDu5zj6rgE1rSRshmNBJszojHBHfhqowSl
r/K0qpjkJgqmCdqNaBIiJJrO70luUk8YngrRXjs5xObYyLznPDmAJnxaTHMpbw1sfbN3LOi2aEe/
o1fTJWZDgqpYaGV30PmHlRIz2iql53aht8H70nP1dNxnpGH4tXSTC2cBlL+zIdgw/+u7a+rUZ3I6
ADKIp8HuntWHbdpztLdfULEcPAvPxNG0rozKZmudLGkku1d3heaBNiPz+wbWoi/+iykiWC3ILS3P
0sngkRDVCPcw0I54AFSOxNc6KPGb7AIxwhkzmOyub/6QIIk/WMuaM/bnyB+BEameIjGXUU98gNzV
Msrh07kG7CoDmygB45hHuKs4qKwJS4mSp18QcgEbYGBhZnTP4vXu/Bz+PeYgP7VggemT/q1S4T2n
a6E+2fK7bvP2tBUl9lJLTIuZWRO7ZOQCO9DYmrj/Zzz0uhPWusYYfu0OUSe8DpGX87VHbOUt683i
MEtYTrMypve/f0ICVZNyOjvdL2xoYKAK2DIHbnbSaK50zoCK7VcD7m562jJYD2hb51XPoV+M8MSG
YinSSKtwH68zHp1Mjx0U+o5/skWNgfM5z076FvXDjm3nZE0zBDfPB3T+XI8eWr9oPdBvw1DWM6ts
XnrUXG3BIJgIEcSoJMhWLgkI2ehnyg03YaYmqK8X0NojgCkaq1mVVi4Vwp17jIov96UH1C6Al/wB
mM/PskG7bF2E3xKS6REq+/68ljoazaNkAFT/99T8BHKvUe6uTNpihOrdqFc7fUwh2W4dj5gNmblR
GDbwjcA1IzP247/VCrkvuwIN8I6TNs9sz22QTkGxTBZY3ua1INQXdqxzPogIVqaDjXcjGLFhYQpA
fyltiBC/pxyFqzA42ZreB1tZ3cgFAHbHXLijRXqBwPHvY15DQyS4dLYodvGicsz4CPf+rTM0cHVY
iwYEhnvLjvtvFbAGGWgdDNLr2VFr+OpFhxov686EaaXsu71EyVPtTzd+ryYMrK96p4E1fZ3gkqUA
5SgK4oOYrTMCEe35Wx3OmfjmNMFGajRit0s/FAwdsB619wXVmBoIpqopfFDfLVGkEIvIzOchbR6V
LK8GiLzvtDgyOfzkuKvX99RNV5jyCfcxHm0zhL4G+LYNtKFF4pLc5fiylrGnkB4QSOM+l31rCoC6
MMeEYtIXru3+2UrVTsRaADbo76+SHI1c/NI4xacr7vqiQ95W9a/n0KFO6Ap6QRGHToG+EkTFjfFI
gGh3RV3J5WfLGNrM+pnaLX2yyFPh71qeCRwto0h3X/CmeF+k9cj8I1SoZO+6ZNl9IP9Bv2DAU9qa
LvgVKTuD9svlPi4IZ8qOiF1IfwpwM6WmFy5lMhyla6KjPby2unG287cqmdujivIKJhyP2Uu91z72
kzXV0RSny9mV+7TA2CoUUqqBbyHWUEB4vEORwvmFJ7I6BUxk/o1Jcz4MF36dIuq2ZSdEsNR5CqEO
jTpEhU34DvY5gJzBeohZjZpU7eGYtqt5Qsp2YGJvR2VwVARmW0Wl9UzdkssWRWO/usU+I+FQPwBh
7HmlAemvGDEsFlJXoETVejke89+A0bQy2PDTDwTwASijknL1RrkdFQ9cIagiX9FMn7Tw9z3s1y5X
mb6GVbjfGkHlCknUu/lqQeA4P+UWj8GeMpSx7g1dvKEQhM6pBq88A5VDzdN3BhNHSTEQiKd0PtMm
HbFtUPB2z/ltmCqxpq3YfUUoCgYUq/szRu39Lbb3vx02Peay6ksojoXrG9osqQlWESFfuzROSZt6
OH3gCekgu8ivaAke9m52LIz/e+bK7tqZ4ydlkXHNsdajmzsxmTsWvbzinKChqBd8VZCAwWX3RCSr
GLGHhGf5sF7WYFva0TVD3kSCne0mh23EJnNbSXapngG+nGE8bkpA4faKnWqsOk55cKamtdGZUj/j
rIN1X1TAk+VhxLc2baWhq+sxjMzO38PJ7QaR/M0dvZeP4YlJNzNMtij1Ll43jEmQAF/bZWdvlqr8
oBF/shBMtJVG+3RpAiyeE+FYnkW1l31QkGne2TC9iYvP5bNuEglXgWUqizb1vakmvAu6KWCjb/cj
S+kzdH3k6O41ufRUPS2ak6dRFzahoZq7LsFonkGK3Lq2Z4cmf/oal02/uXaqiScIbUaRXjocGcye
+1NSDQ1MeFa+ulL9ofQhWmizkCmjfNsuXFgYN9wwg0yY6IBOoNl1qZDhwP1wQYn3TQGxK+4dkIgi
N1P9cxQO+N1wrJ4t8LrNsz3EQ99FZ8LyXJnEXiDXW3IeAer54pwcH3pvNCQAjXV29IBo9bh1sxT1
ZnkFZqLKf1lXuAWNagb2kU/qw8+lzJ7QNd8od2oBH6TBCnmPifQMgPGuppZw40VnY/fAnvBlp8J2
vcBUQw3EWQBBH8cardew7qoKaA6l9MfAYuWAYuAZ8XT+/lloIft1h+7tMXxYwOvKTZV8zKbuS8Qa
tec8msYwt+UEyHnO53El/y4V2x+mnrOJiJAHiPT73XkRiQkCFqaJh8L4NU0jqPgxvCeG5J+o2a4l
1tCCQr81jlhB+ttYaICE5zvcf08SfBn0OrI83Q0o5DSqQxoVldyfvykPqnfevgREKko4diYV/TlZ
gbhdoqd5YJ7EdZKRFMYQfBjUpn4DCSaEILJQSXz2rQkD7fKm8HFttM9ABqVsDvQD6UDvDU/uZp2V
SVPyA1zuKd1BQLdAZ2K/d+o/Yt6Xx/80BEvMTGtQEm8yuKVI007TdDeMkZ0uY4J+6FpHUoCXRgtn
1mO4uagmG6ix2UceCy7pW5Ta9rIJ8OO4o4otAdOADWJYGS7xthW6AiK8fmUoP7TPsZ1sYj7Ob5hD
KC9xnmRvvZvPF8/353PQmw6uVNywbLnoJcLY5J6EflDACznADG2SJ5yIJiemIaEZGabn+N1wZvFS
aBjOXV2Tp4U7Er4hQ9CTnH8eYvaZv/mmNKcON1jced8EMm4gDyokKAHNwCqvN3Qh49DRg2LZTgty
UFqu17bwtCrx1WOOL65tomYQ+RPdgmRY8oiD02AQa1tc28LrttQkXHMl0Jpn91xHLOkjOSpbGId1
/9crs9F1fG8SNYtJYUa1C5ivt9tsj4otpy8JeAY218KRfxsyioEM/FKB3Z+DNMpfSESGf0wzt6IZ
nRqNGjSSd4UIIP0epVHR/f604z+kHCHqXTq+/EziQvaab/niEIzowOVsD+eF/BEVmak4uDveVzX+
SxPXZmSr3ZTlax1/SFbW3bFTLRXwEkO4+rfeCQNA9ZGved/ek7u75KC54TjMDaUTzw6iFZGU0tM5
9A7BH/MJKOK6UUeYu3VoFVHr/a59vmMov22klxbGIB5WGZvEtsj0b2MC8jRUIrePi5c8BSjGmSzB
wFv4u7m5DXhDctvRKo7B8TN/2ubaHoGUrovUkerNjxJLpdfCCFFOmy/JkMQo7E+zKB6p2lXByU9f
b2uG0iKwfpwoVbHO39NzD9ynq0pjnd1wHKURgSdfS5WHKbQ8VuvW+zEWNpnFohaFi/A2UduR/piQ
Eadhkd/Wp9X3X5Kte70wz4yho+CxRBvmNZzB4nhX2KfgpIODXpaiBmtobmWqFKWvH2UdbfE+lulv
z7963NnvdQiM5Y5stNFgiVhiZze6rCbcn+hkq27ev7W7LQ9VRhIr302AeXL9FqKkNF3HnUpEpTK4
/AbkVKmp5At3fEYwDqnQgvImRK35MVwDz5Y8alcp43QvTh6lhMcQoNYbq68zldNEqZW3FddIajVK
1ztYsQhoYgYNDjLNh4v3jcPWC5DYgBY3AUsqPMfNURqTcQd4i20AP57H8nlRdGFEFnroT6lNz6IO
C8yx3cJOSzZaw/8AMlNtrrK7yd+Cs9TLDWG341sL7cBSOLdRzCDRvITpr375FPidqon1xpI4PeU8
fYJlfnsiCYeBX+pG8V1jryzeiPOae4gyR3991BDET0VI00JpFhofNgLHT1V2lKMKyCWCjvxqPfKs
kntYUFnXkLWMv4mjtJVzRftvCyXfLZijIgS9ySePocMC254DPkSoxlUrRorQj8fSQ2ZqZcCPSFMu
EhnyADpg4dGJJfuMjE8tYKrgjPX3CPaXDYYP01L8/cwSFbLaeMCkIaFOf3Vn6fdPNOwJslOQpoLB
0VIi3Ww9XNx2pOGwRu/UvNA31xMPQEkmOqMc+7OHud5YaTf4twwSAFCr6LZfbMkFIq4fHfaEgcUO
njUQTsLRMbX4swRVA4s8zA+4quuM2Ccejd2UoiqR9gH+TNYSQRjxMmA82mhtB6tD0NaNJEgF4SDS
9koeL0fdlauDUR3vGSvsuCHTtItcngVod+Ab/n/248qvO1j6NXVc8XznyZB9SHsomVYbbiiSEhV+
pihryClcxpDtVChGPVLsJyazFNDRb1fPLH5ttPFxe1bwmeEEfX7Ot1x2ZiNFaA/jaqrlQCM/IdP+
ikte/1IxJQqfqf2T6A+aS2KNS4pkLvXJx6JNXo+kAtn3Cvj7VQgFzODs6432nkfFbtpjfKuhoNNi
2JJqDL1qwEHyg0NsBHWzBFUYGZZdCFFcq7vTam6iv30s2U2wWfwzVLQOWoX7eIa7MYAgj5qCB862
jccEYi0wJBnGs9BXhwRjQKbngZArg+J1R56omrMnxRumhpzCGIm5Ac3U7TG+o+iVXV9mUf2Tu0zY
RiHlGnpA5U/phe0N2klbM0P8yt4gITi08JZBYZ2IjRn5rZZq4a0koky0kGFDbUQFF8JOId1WwluE
M3bmVj4p0MSqTjKR6OZHT/Yp5YgVakaUZX24CJlTpzIdn2OHuLP9Jfilm1FQKLToVHDe7DV7VEGZ
i1572upk5/BkLz61xzuUp98PvQ1tTA+Y2kBYoUG/WdAXiSmjXI2NiwwhxvmIXXKua5vNssAqx9ps
SAaXkooYKe57IgdRPM6tAXjXYGnj/aLWNnpwWB6prLEBmEjOP2YJluKNSs7YGual2EYU1wkZUZ5q
TPdT4Y/2jwepaVVAEEkvDByMku6Cw8tzQbV/jjxYo7sNgG6VvHXX9U2YlcdTWMrO37mGTomzedg0
YDdTDnj8y9NxjkxAusVJVXoo28XzS6wvCqpgR7TJa+7MLQ8B9auzZ+HowLHhFALMGfKoLVlC6+Dn
Rx85gefyA4hYyafuU5FJ1MlL1dBovH2gVGwGf06ZytWTldeiGwfJJUUG2oAPsDIF1nC+/QbSQXeK
ulUmWIWgCnq7MfglnafLmf7phqQ6B4Ra6k6jsgr/4QcSlyDuK4dU4Wti6oBiycYnn/zH75l1om22
6t6/EurHzJXHzZKZm5xO39nIMhUrJYL/x2EzdiNVgLDb7tee6qTWfOyEd2jYXdJtZDYU7GxNWiNz
MUujxq8vJ8z8prQY79qPJStN5jgxXFTDLI2krOkawgeaZAzE4X/C3mVpgloakHEBVZ2YyMXrA5uI
DG1hZ86QZxSG6224R+Gjc1niIyxHZWHdakmsSOqWNp+ZAuW5MlDSfsnYYtnCh0UlgblI7fUsRdku
sjbZgbd1sjNrITPBXmjzzFm3++/A45fT+8++o1SCHUJ/FdjG3ZFaHctBadVcvbCQ4u2J5ywer76J
AmGLELUpUbWrtcYlcxb8DXHCzlQOHiZNjVciSGUTI+LBfz+6XXYhzdxzdDOlk/J5q+1KB5jtgAl0
mfAufmFbRlBpCW8+kyYUEi6whFC916LKgx7kXsBdpQvl3k8goW+TTnaZX1n0U23Qvy1jVtYfZw3W
CbC3visaweFwIuaQicA4DabAdp9nHqcEITzEfZ76WfcLYFWs7Q0vT785vr0sDXIHvUbUZpa3KWND
9MfSdGxlRmmRsxZTaTAlhbzAIxiYKvoWitpHr44bh1vvatFCqydoWMneUH46lMBUfCzpYjNFylr2
etctGm3riFw6EBRShgEJgJ0l6KLl4uXSXcRnXet0ugCGkiVoHrIZmljmgJmCw+bf0hk1pTkqaG62
n6gjgERPYWC1gC1BAg+RqifJJeF5fGPlKMi7kA7+WxX0Q8AndiQZoWQnZb+n9jrK9GStO1bnRH4X
qB2V/ROL+POodeYdjXkMMT1czhl3Tc/AFPw4TGXRPN5ubdjCW1LYkywaMrUYuD2cNp/PZ2rUDM9W
0XaUoCySca0//ujIkBXBpmBHKvu3ePZFWM72Wg8PVOKNuqbZfWF8L6YaNnXB09py/wSNP+RW9vtn
CFDHR3I5RjXmCxmYTZ6ienAdZ3IRNdnNvdXU+RozcznJ38o6aLWX8c6DpZHKLrv66vQfBw7zORKU
ZaZTjCJzKI1l1lgfdpwa4h2hxnjqR5STKl+shVLF7e0W3BlGSqHFLfuqdeuVQBY/8Wez1CUtwJhN
Gqkph3/Z6JgJoFfZ2T1Fx0DalUTF0AokrVtwt07t+OCaIvP15aMmh6i+uyW9kY7eupAlbak9vj9p
oNMF7ck5u4TutEhTGz4+F7CZwjupskTu9S67xawLCZrynGuWC5oAB7dUF5abSIGE9HH2MFwtPkxD
YmsKucQeRkZzJentCvNhYUJz2QUYq6Fl3uaNtSPtpkOqpVsILiLFBA0WYtUTy8jK7WVXGHA8zIrK
K1lAt3/ZPWGVfyHkApx4FNOeCUZSwRuiLn+pKvkFh3mY4wLhC4+5UTy6mhU58p1vZFTgCjbjZg1v
XjwuP/4Ri2JhYqGRys9fajjWm1AajiFyK5EVx7SHTTu9EFaLDwQzAp0R/BWiLfbd1vmvR5Y8zRPv
2UPsVZcZ3V63H9o6YNUmGDz1mKchNWv33Nhd0tZUI6IhoumN1XV4IdPWz+FBFybhGNkfYJzrp6Hi
uRTQ6PXwaIquowcuoRiJH/7GH/vxHhXWilFCx24tfsYKXnlm5pJ+MmVBENGfkiDirIwIFXfTIB0J
Br9So9FoqeEH2ApKbdgAPhKEMylUE9wH/Gy+qLjxGFj4VwdB662EOfUK32HMoA2Ba5nBX9/Aid4j
xqAuxV0x2+HFe+BI8yTYUQVxDiUY66eD4YBfS632pOSlyiA1sP+BieXBjeu9q0X6u9Ag2iINR3yz
GolU/IsfdBEmr06NKjOTj6Nprl3SClEEAWRlMS1t4VPp9ouxL0YeOq/FvCCPXViQJr85xdSv9vDo
aiP08C4pRspaQv3V57VgvC3NeEsJMcyoseI2yMHSDKJPunoFCSqDq4xEgR2LFUFTxnSgWNP4Qx+x
MwJz72PXLuEchIMiIO8u6rmwbYn/5zm6CmfI6icb7I1D0DHbG/CPThme+CaJxTTHXfy44YHQ2PJ7
C/Snt6V/mYMUeFpZ66MPr8H68ONqDRvAB3mNZs0VRYAV13ZrYDVfCssjCdau+SAHWbgk5bS6jJ7t
iDH/eW6DGJRqRKN18cdClKtD2iJWI4jDytxTA8IZhCg7XF/PK6SOmY5NLmWBFwwBriohw9K/7reU
th/XvgbixY/kmocd+3AaWN0hSmxefUKABkMzze0s/xY0jhYTxOr8L7lkPgZYlg74iyODVvDBc5Sg
UXj4mA8ujypUHCIzHLn0otjsV8QP6EcniTSjRwqHw1Dmgdm/Rvdg71kAaO2xnLVQ+rbnCPYcE+4H
uBZlJJbtWQGUoj75l0dGLV0jn//hjrXd0//qRJI3EBPbrCsXMEibj9TvJfiv+PdfLK1OGE38WdHf
riPlR4wV20+8fT8ZscM+YPbjqIeCXm6FJXWFCoQzJI5IzcF376OWwzEaGXbaD8di49UwryRMfFvI
Y/KXKelsix0nHzUhf612k90IqGxg/8yZLeooefB39htez026LbzVaAdG41MkBxKoPIbx43UdGzR3
vWa9ozUds/5IYWpJXBkasQyYKwLy5J8WBo9onJk0uBVvyPqoTUI0BnuQcbyUe1cLES/ztpKw3h/f
tpjYz7Pqn0B9jF/vk7JT3Zj2gnTIKQE0EgU4XhZYdfZFyzHhRddTz8GjlLxo70jtF4ggcAx9sFo+
XnILrUz9hFxuRBbl1EZQfHr3oaWd8SteaRiC2KNmfmQ3iNe9bUudeEd3ADPOqH8Y9koRp8I/4ENy
pNoYik2YuOWG1+/mcsrhm4ddI4m2AtkY+yGd68IMbLvkQSiDWeZq98eaGq3Dp0NXC9EtSRZO7Gdg
ItzuYpswkoibB3UceNiJdQt5CypyK+P6Gr2ss3D0H1PDE5AS8PmjqXEXnhgcvc8NPY9n5Y8FaEhs
4ZnjHSamIcFixGVowLbI5N+FrjrerKhn3NbIf2d9X7YI5zbwV0wlozx+e7L2rg9vo4U7en7WtXjf
7wfVRd9AC03/fki0W90FEgrAkD+3NZ2WSv83XaTiqGZOkEZp5X+EkdV053ILm3hY4sVMAL/pQJpe
c0U9UrrhVnM9+ETxv5ND3o13qeN1B8aTjc+duOY9HNP6pTbXiCE+qrvLDXz6kC+4JWWS+yTCGdEB
lXE/I1knhsKW9XBIXa/iMawhe1Zd/HHI7ySmWi5y+NLr4r0bpDs5XDgEt6Vz8jD0nviZEdnL/2n0
VgHeL2KDihOWq65ljaXNJ3h9J1DY+CbMPOOV/7TxZYQ/lBZXz/nVrySDlGZ4v11TlwzvYr4STJMP
SOqi5CzDK8/LkD0bV02LaTNCvh/C8Z39qCi5E+D9i1fojkkuLf0+IrjEfvfWzfi3g4kEwh+vrXOD
sJT8K14ozKhbLuBE+uf4w7/Z2NDmLRC1aD58Z2QGwY74ghUzKEfNetXDIfZC+c3+M5NtgIAlIGmw
dsDYGtkL+7iD1fK5T3ww2NO/EMzPHPgx6W42NYbG07UsFIFlrCjaBo+ZgMN7y7m4raP3rebJfJB9
X9AFzK2DIlTB2eJ3oTulmX7Tw0OErHuPRpobWGibQYWRLtxRgdxLACeSIIgFuWfFdMdd+yRttPRt
buY0aLONR8KDkCLOPJxOe5r/qxl4mi4bYUyIt0QjiyIOy4/aXsVVpePLLofHbOWAvfZhL4fEvGDD
wqDyujfnI6zHFltzZb/L76LicrBJ/LrhD6Wabqy7vdEK2nW+3HMTVZXgZ7QLP+4Wz5EAW+Durx8Q
xUaokZ88lVcpF+RArozoF8aOon2/BBPz+ZQ/WoYpTw9CywPjzebMWzGawEpLDN24SpDoPqctn9db
03EhVmEzKNkI42M5xKN3IABSkFcc/vL73oftbabXQeLuZlx5f2NY9bFK0zJoFJhlFUnKmjau7aWl
KbtL0Ij8ECsFgSIQYG5Soh2R+x1Q2Lhs0+dJDdrTSYAGarHEZsXvlpUVrsgp9iupjV3tCRJuf9bg
FXcu6zvvAGDJJ/RCCDVEd1kdFkgBpMuxaP1FoX8Z920Qrl4lrdsewAb8Hq3BLLYtfdEN7z/5CCFT
JnPscHH0sh8yuywor+bv2PxuBxTUVHI4aDmCFP26LDFNtWGMNhqcSwcAdTumDCnhS/kOlMVS8z0Q
PEsJ6RUqs4ipH+naS0rIlhsMF0m9XopEpfTvaGeSHczk4fMsfgxgFRz71MIzFpwxNpM7vHyGWXl+
zaNPwLtNYJGp+DlU1JMpnp2ikCWeJxs+EiZJoVrKzo7WTfif7nHsvMzOXfWalBotebrj5cy6vZ7X
dUTHZM/qVNTrnpAGKCJmOzLZAfehgl8A3ZHJNgNYxlLFNULKOLMZdDI4KIhCFfH3kTAqTeYhKhX8
4G8CrN6X7k7rxWh8v2XaXP2WT0w6U0ON8ENDfl8VUlBnGchdx1CDlpaJRdofQcFvjmwFTjU80emo
qeSFfLTaK9xTEk3v5ThA2GAoozaCVheM6MBIr07eU9bQtPGHKWfyw+oJ6xUznRRowBAiQF9q86jH
XQiKISZDeTQHY6ap1P3r5jmARJvGQ678KjrcJU1oiwEk34IL/hm5ytqr55cJXu4YN7n3k3MLODRD
fpcPrf8mi5ac7Eyfizg+kJAPzTmTrE1U2xOk8FjZzir/4m+pUMIA/wsk/F7wXdG5Sf1TNZSSZQxS
sOVJxLKccWPSjfIlJVXdt9eNv/HCU7RjjUqecg6calSLWoiZQejqURz325+HXJvL9RT2+R4LO1m6
G5NZlvTbnpv9QCc+V4gMG9ajx+TppvahUEvVrr3M/jMeChB6AEmH3IXzKbYWh1HfJ1nTpi70nuUl
zH+0fOBFsJ1/hVOpDKJ0hngzBg8+oH2o4/xasYh1uy4YzA7LHSQPfvAFnTKw07F+bJhrFImMZmTN
c2tb74ArZIELAWXlk+kVgvEPCEpHe9Hv/JIPF3VRrSKPKmoz+851epTDGOdRGIE3Cz9kPuFNC6D5
WjU/Xob4+QbJt35hC4aY+WMtnTXRuDfXrP8BPB1fa7goWs8o/GrbQfG/feTFrpTr5nvnFHv84qTl
ce+UQIaq/NzFI8aQl5HGoYOyr/YMIqtB65ta/rOGaBw+PjVPD+jV03s5edA4f0X7TuwqDbCLggoZ
AGAIZR8=
`pragma protect end_protected
