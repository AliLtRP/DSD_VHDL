// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YPIsCs7mRRD5vrftc4rptiaKdLmuUOVPCaFLwhhpCRTqvU+QRFbJxl8TqwgHanqH
ahHvXKlPxMXYEXfhLNhav1zxjovgs6yIuPDUCk3Xdh9kQLbJ2DARP7pj0X8xBCLP
dcpE4/wfUacP79vPXWbjGP/E30OniISD+7asveQ08Mc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17776)
9Mzs/DBqnH/7OBbsieIyCUw9ERCxnfk6ITwSSHf7ZuOY03pSSPWpnz7zJ8+mKf/T
FGena56PVEHzjgEdGltn4tLJ99XjOr0aK9IONYgqMa1/diAw5xBNLlhOpiZ0HKqt
PIKy4R/BdrWL0h6QI/UzaDY3ah6pHomlJQSdjdzs3TVenuvVyQR6b9ZqAnIvK2/P
wjFGJJ0tGabGQAzLKKe8JefF3fL8eItr/vOPqvffrN9zsMGS8uQ2IEdsPfmm2opU
ynIVn10MfZ6xM7mWIQ4w9xe5g5lVF5OPDdnx0WsQ0VnVwU4WOUcQ+J/r5YJsZEVw
A0XhYDD3Zmxx1TASxOQ+wLVHTSDqAqnTQ3FAddkbfIwSABsfM0tM1obvxvUsMKsV
Q9Aitm9cT/20pYmej0ajkA+dXiZcGCebnFDz+LK+ecd/CWn0SDh+i4pTsDjUZ+u+
zM7ZwQCTOQfyTqdjgCasuBixuUz6wiBYTMA25XxUhsMNbtwqEpfaspUMrIm2NIty
PHAU/LdK5qYed2t47dH2k0e3jYjA8rsX7b4/KUW4QBLzJuYvt7BrQvyJEozW+T4N
+SpfGyIIOLIkzfW9Z4RoAiVA71j75gmVr1Uo4WJN0nfSqGQPW7xlPtI/zopmLbeN
bn6A26ArqICK5djSK6gVhT1q1419YgizGejiGeZ7qh0+kV7QbRPxZ8OSxd9j1BvW
zqH2Zy1WQPidzYSGQJc7iXpPIfFgIXk/RpEbUxfHkc9kIe5nxiaCM259EnrCeFyF
Os9bLHRqdixXG4aZ0Qb3367OfgHZt6Tj+eivHo81C7m/qTiuA+qA+MYHR3xP1icF
NYnlJwHsjJSue6QxMqCMkuO94K6qLm0VUqBb0qudFBVzAMGrXLPOBBMNFRdGvQcv
6GCEutpfyfWFKCBNOsPG7vXB81lZh/oALCE0LgUnAAt48wbnfW6C/8UiPhq2fkLG
bgLEKQ/MWt/bx2sJM+paYD9LWYe//VEqrB3CehhSpPSVweNfoXiBg5JCGU9Xy4Hu
1IpDUHl4s628mlLU3YdVywx3pT6G8OnRoF9H3aPKp9kzPPieUXz/+pwmcpPTdAMg
tnbV3x6rAhGb+he6qArJBdaxlBf80BhmQ1XImmLdw0wxF8jAJllLBeVKLA+jxCfx
oyYPcJaX1/w5UefmLkeLjTH1GcwA+bJ7sMZsy7a01ju4EIKgTK/LlCEc6i5/pc4G
3zkkeaVtjtAyf35gVy4/myNtscnA18/9BfCLc2agDGKd6j1JQfbKRqAIiHrkPPow
pw8UjGaNI8LID+DjMp2TaUPxDxxTAXf1KPzks9a/ByMlGcPJHmA8QfQ6hC1HwLBL
xWD0PgGqgYXVIqYCvM/bGrMXpuAfJwfJjk3/VRdnP0k2yr58YnKRS0/4p53K/oV1
5cuk6XdixhaCBp1ibD4zfSQsmdTVAXjwJ7MbXSATRbPYbQkmBEtWLi6B8j43frmP
1KuhAnhMGJu0hyeu3e1n3+pc2RdwLsDUIY5kFVtcr0dRxCrkllw/3E6XyH3MrUIh
0iXd1NgZ8qEAJ37OU5gkhmnuyLeDLScN1VzT6iM3KWtuG4wom9vDYR2DwRw7HUI6
sWVLryV6mqV3CHwmRUQfu4z1sNwLNNP+rAL0ji0W0s2UYcCT7Vf721xouz98jzh/
UHrXiBSBGxuhVuVoxzIHUML2tx8dbgNIhrGn0+peX5ANYQ3GhNw7UwE5Y+1pm78j
cE3zFcZMYPia1cHfyw8J0H4KVXwBGmxgKtAielfcCVeQhAfeeouWNBqQeMMS+jCV
ZFNiUrR9lVUxhcv48F9PCZG8wJiHvTdKLFIQyA/vPHyoO5ghp8UY+SI9q/wvcNsj
Begps4DB7Qw0qbjpdB3jb2njZ60kHVAPSf3XDxYLcIc9h8JZES93SpwgVEQ4lOJN
pZ6ITti6uf8zndb5YNp5ZE8osLlkpjEUC4JExaFUIpQvYPynaL6bnBeu0abYTysE
gB2h5FYP2InoPf5oKBi7HRVKy7i25LEX0AmMp0XSY9snnIT96nWD+pQhO4MYZ222
EvjEaKboFxf6mVzM0tcVXOWYyAcG9Iexkjr04+SkZjh8ogJ+4Y/RbScZt8vYTw0Z
J8/ChHJQnAgPA0iwR3ep2CqF2quYKC0vxcTIO5RZ6ayixErCEIDM6hTdJ4z5KZiF
kRJ5OM70hZ1xD2WOUzYjf8Nadv7XnwfowmrfCt+ElzNW8frM7y2vUCzBRmT2Unkk
hf09eMWDIC1Xu9Vr8JR//TDBfrqoJeAzTVxlFo8kQwz9DZMHoPlqb+q0m83yPryh
3KZp8yHu87UHBTTnv7ZQo/V88330uwJ2ZWvd5i1z7Z1kpgET/8RAcPERfNXT9nEx
uHvNbKoapg3j8MB3KOAmvMUBqO1eknUihTM6jxrQk18HG2cuXJiWthFdBkvPNEuk
9854Dvvf/duy8PbscajniB/xjdyHPhQIfz9b/dF1fWnTPC3+fDGX28HnUygulp7i
J8fuYHKsPZcBT4C5k+QU2iq75QpozL460q71pV6n3LCzukevvtj9Qn2CfCMQDtQ6
d5bL+IgBmJ+nMeeA/pqrXtCXw3Xo2goa0nvm1xvKMPkRIrH8k0aGBRku5V5DEJeQ
5slQEdp6WvmeAQ1OQ6troyUVWs4zGQ02I2CCLmIZncoycotZ+RixZba1cFSuPWhQ
ejaa9ZvJoOyrWy2kD7puV+aN8U6ti5CaU5hw9RnIjxqwAjTiMM2yoJ4KhJX9CtzC
AD8RdqqSiNXbNe2DF8A4w2m6jmItEA/I1WVLd/cKO9fc9g4EsOFViyKcbEUh6Bgq
ZrozGPRwRckoFacoAHAqGm4tfD7MFW4RgpbFkDTHsYGWj1YbJFan4/Rg1cfs2WQJ
qIemTGmBb+icmrOnVHR1wtttLeo4ZMsQd2UKEq5VRAuRzPkSJeog9v433wVvovBi
qqkBIzgUs7A81Xx3eOnqFnANMBJ7uXNz33RXJt+I4IFafyu8C/d82D9f+AjK/OIk
W+DLjKCzh0mdnMnvvCPfZQF/FTWlDe1eaTKwdvS2g5h3sHf7o2JTi+DOogiwWd/s
AXskk9zZAsWTYJ/Rw8ikCFWV4+dZXnrKHUyrgCiBJsjjIkDhVZfMlsElQMB21Dt5
2LPd0tN+gMmgYoqTmliZxbaO11LP37+lW7BppR6/QtOqcGdd7ArP91IKLZdDkcXR
gCg3ZFgd6Ro9THqx4ziu6iz/eULwqB4d1RiYsoNf8oIcbNOlbfhPqi8N/NwBYlaA
zZqj4rH/rT61KVfrWCIjwFL94wTCCvyxsPmdlO0UNvY4XJlm0lC65681+VoU/A+z
TPY1QjkwiD2mZ/uZ1te9Qy0Zx7ueipnZ1LPP5Q7gnwWtMee57UuP4yDgOzluYuOx
DavxEzQdRyHJrUDljIJFmrplIU8iBEZpjZMIXoSMBH5LJo05uOKw9K49lzJw9yRH
sMRlt+aXJoc4QKO2BL1pUO4gSQUsWqi2b2Rs2iEkHZ+Fh34GoNbSTn8u/QgOAq6+
NNKv7H8PSXIUSG3wvosmQu6TpYDmb4jJGj61AzXuHg81YvoxCsh+OMNS5j+TtUqz
63+nl1IS6dQkiUQJ8vGwv+tGyZQSDfetc+d3dudUK7A0wwjg/RgoQYpeIUS2a0ML
5QCF0Fu8DerqNBRhh9Wm3IufrpOqoqvf7PIEYL1SLlfdLIRh0E8Z2tqgqcbP0a1t
ngWz846HRDk6ZKE6mkYrJhOcdaYRO87zOnOq44vBi9/vZMih1jKaMBQHoIH0r3dC
+rU7ag/Wco9WbKidSWnIB75pgFWcjEcUMoUttvf1eCbCNCMtEuY8jU6651DReYeI
Bh7eF7H5pMDniGAHKl5FE7qaDo07dmcCNJ/1YY7F4byyo30zcvSWVqRas3YWYLuI
ZkoBmrcxr0OhLm3esf7L2NqmcgGqgW+KPLNLLVzUvHH5xHxk2BDzWt7OEO7na1bE
89vhJEWgTobTINPQ4kr5acA43cSU45/IEpK4vYqRfKTiRIwY9mXnpECbazXwmOIj
M13XZgOcZp8rLDS9OIcvGVrO4lpWq+kGJw5WQ/8mGYr4pp74BvaTw745dB5eKVl9
/fW9/EHK+986BH14mdTceG4bHjVg8yAV/1ALGYtPcR9koiqE8rLG0sH6ve+srQSr
IaTs6T1IzhwuNuJvyQCBj7OvjxCx57P25+vSLcrcXsBDx1KhcJJAE5XUVzRm5FLA
SH0BGJFb0Yn8IKmmw0PSZ24vBgB4dw0z2JhFqp77WcIeBoR2mlG/bLn175TMvMjY
RHKTQJPGrSiiBkV/CjaT8+li3bdH0fafg1ZKvU3HXD5vuSf2cZTzCcMv6hmqqYoI
D8ncw7+UC8T/jTK3wThXzadjGM9APNwSGTz4lQOfFYtbsABk4ix+H77aGIYrSxNE
gYM9Sq/tAdpLrb6A3kNQ/mJXOQJNp/nI2j8LyvCrGyvmCX/PAHQtW35dbiEwYq9f
mANTB2eYf7dkyN+trGNDrEicVFn3vv1j1MTRkclP/w8bVK1GNOggjJFMEgTCMsdi
LnMJSHEvgkEZUudVvXosVJESdcuzhSC8ew3b2VVPVdCHtBGFSfzfEv9jtJYMKMlP
wVqEDflBFtC48mUEMA15Ojj4DfxF/Yj5f4cUNomgkgJQCAfiVC9D1Lks3GtuFFI3
RTKvXtz6q5qihnmXtNjztiaTLsgXgt9aD+ZrpgC74shg+RFO73I7eu1Jz9+4wAH0
oRvp6IcivEQ5nWgs4xFFY+uEF5BiqvU8VciieDoiGNfywVPETVo/K3SxpLlrBDJg
5ohRp7uu4LJrzhyzFzlDz0XUudBv5D30ea4QriwLSxCQG8eqC1L0BXuAbo6Ip0s/
atzwdpGICSHu5264pr1jlUwDnjETug0QQSwzL+7CmjCev/bt/OJf8+RjjHgpUAa3
BCfSpR76Bbd8seWJLelqWCPSYkYgJLoHzEAot/zX4SMxC9StpD2Tt6y2/Ylak3ir
CDX78v8SZS6XuRi1WuDrDB/sLYaF6/Thhub8L+RFVWr4Rb8cWz1Afg6Zrtoz9rce
A+FBP+GIYbAmNP31WlWNrWup+dL7nixVGJ2T3/AEP0i0El9UlPeqF0oToFxNtVgU
ZGpblUkztcWWlhhk6DSkgMNUmHF4DXx9Hb41X4Scc9TOs/q8JtxOfbDilDhE3/ix
dOFrOwJP5pAILhzI5m0DaCkZrGoWYQkGxm4AUA4mKZSZoDksz5jJ7RVakiGgllVJ
dN+jzGWtwPu/zFFGiPGhbfWX54KI4Qmou7FdCqLhbHAjPcAdX4g+4iwTcJRRn6fr
CVTpGx0gYmeMGwT/Xj9SO+jGRPXiZhJLRI2imT5rI16qAO/qpPT2e9Dalr6kI1vu
6HJlhrqpP8MbuLMa4vrTsZuLnec6NMjofzwH1xiK5RhBx+qc9q55ulqyVm7Fdd2z
Ya1BroFZaEFvhGqHu/VmZGH7Vj2ZiCx3tkdMyts+Pq4+KABUm9pLTaTDLzFP67f9
RDyG+jtebKWYXO15Ss4vwGGCJuK0oWMyKaeLBo84gepbhS30pTSGC1/QVmlQrKzP
HFGlY6pFGeiGzZln2wzz1SLGRdeC5SHphOUIlVfq7XFPb498c5+pO3yYR1g25dcb
ECYyaMKv8ntEK5ChYspJl87utX6cTZI5KGoZXuUKnucKfTIqcA9rY2oqElP+/8Q0
/7r1DlE/kGY59DwY2eiEHBu/5VmEE8ewH503vDruPx+Yl3o4VS9DZJr/sbWGoNIO
YJ/ScXPfgzY3bzPBEH0I74ZSPEmoaWFj2jNzoDgJmf5LyEBN7dW+/uLuwx6ypPo8
5ptLiAm70w8/SWDiutjnj0+5lmqnPfPzyp/drdpn9SGtNzMKy3xnsj/8agFqkuIO
GDHMdkEmdH5vsuyqiygLi9VwXJvGN+vkJXyRdewyZbl1xUno/La67/Pmhfwi+S7Z
pP7bipMpFX0sVcJuqER8vCl9tSAcaNhLJn1ywDqDtl+PTNk07BtQqnX8zhwXyeC2
T6YsBDIc6uUKYsa3dAKMKlR4b0ZW9W1CbZTxx25wcvlszDxrsPF5ecQraVf8b9yT
csVbGkhUp1MObKBgtsDSAZwNy3Gq3SMDwpnu6NDire82R+kjPqBgyo1w0qYnp/T1
UNBDqYxSN4kKNlmJiMiR8n1Vi1XoQpgCnTT/XQjLAhG8Gfy+H6Nzo8eXq68XlCHY
LGpRHCOyPRxNiN03KAhHQdbeX3hCfxNkKO/R6VKIgad7aZMjFXW++jRPfFK5+QdM
CTz2bOyM/VgaSXT+JoYPieGZnk3DUKeHLxBVF4Z+f/wuM19qIMS0wndqy5+MmOyq
Z5q03zSQsJ9UUC//rMILgBezuXCsTfkD0pRvFdiCgKD2dKeCmzWc5uHA2+tMsfzi
+iwmkuuxeXG6zlx47pzmv81w+3qe9TbOxahStTXcgaWXGEeJbkBaYKDdfxGvKM08
uHopaXWZK4lgFsM6cgmdkfhGatn3FUcvpGCzKbQsK8YHat9VvMhQQuv1UbVi7S8U
fb8TkhtLevg81CM046dkfLw+Y3UdBLIys3bRpRgP87k9pmWOECPT32bBW8bHoL+y
alUS5DQfepEW4qenY7MWzbfSSibsJkzOeY0892DQXvWUjCdCVvOs36kBLXTCHHzt
20IcV7AQCqj4Ud8q0ddsGLc8rmwNwI5TyeGTJBbYhThMllg7e0koHifzDJYCHk6N
av0Hrmn9chOKVxDc8THFXWCa61F4EBv/udYHu44rwoTm1+g5OevqPLvGS8TJpvMP
AwP+3R9DdDXrifqLlQV89Dkr1fvHYfTOVEn8q0NjSwksItgZcsMTNs16IWrIfZ3T
mtcuZG+C3M7AG8/Q8KxyfrMEukUaAwxa9elN06FPRB1ZLo1qLl3pOepynQFltL68
7tC9ipic1WsHkxInh021wJJqqch21DOIVan2aO/ffG6kRhJS+ITpd8CRUEKXl9uS
l79JXIwkwaDtTxDG0ZMRBagdsLZG93D3SYkqn70J/vg6vm8U/z3mUG6AcAf8pb1y
AvTVC0DM6vfJBdBmfcYZYEAFzDShgTdfbVhI0V/0VjelSoerfd0qntAjAurFsHWg
J1KqCSI6OLQQyEyGbUwNwzS8ZBo8dFUEKMBWc9IPbno4C6MMTg6s9XrqHWJbrKY6
WZuqislW6o5h+BXS2qiEUr0XXPSXENbjuvVuizqrt32z8M1thLXYeTxXg00s9Jcz
ZDLPOY8g5xLIi2HbJoeBvppjB/q4lK2Zziblf5SbXWQvSybaBX/YRZiBkPff4iDb
Y2Ed/YQNDhdPKyoFCZ1+4E1oxRraCMup79cS/bTg2XRKi2LfTWHVk4RSzV5WPvWK
wOpQTrb7FPzYui0cKLQ5sCDv7q9BG7vwaqAXSfc56m38s6oMZseztZeSCXH88Nd0
i2k8k3ZlTpbcLfUZLsTzAf/QX6vRVpvnDy9L27pRGfHQImQkW3iHOIyZbYIZcp9L
b7su35YvPSeQEHayfonD2zWV3tXwxv4wzSQELmYftvdjLHKaTnLx6kkZTk6jHkO8
hzlXoPuqiDJ4XT9kWMJH/79IdVLpq1OicMcqndf6NBnvtsTIiMZwWIiSqj2hJzYp
trQYsjZPFf9s0eCzPmNvO3BGFGIkTTi3j3bxMVddp/DffdcJOWuDq9ByCHEnGNaE
ueWtCsIkb7cNLSbqGw35KrNOHvaFdIYPImxjfwi58qPNZgHyMJ8FfgjjdQxhuLr9
3MMdPs2qSOhXf3ZGf/c/bDh9dOL9TD97Pp5Gd+OTIie3a0doC0zEf09gud8zatRU
76n84M2J+2WhoXEjHzFh7QaV3t+5J337bhWIXPDWpUzdE8W7A3qPtyBRdpeeg0hq
1TJF/JbMAX2LLB4zlbX5HbE78yoG8FajRA1ajwzkRcLHFZAkBM33hrFobBNhpWlT
a5rjTxT49CAq2EttI3ELDzdcvWhzVLMxDNZdNUsArtbPjo1T4qMHSiCfSzObD5oa
Dwb8HULQ7lqY3MB3UJz0WW0YrWnNxeE8iVh0bGBq1HMVu8mloz1BAe6Ij93L+FnN
ihOtSTgaSDAP355nyplwAVytyntQBsjXHRx7lUVPAf0pmcHRI6oA/Gs7dIgWoaRh
r25br2hcjHxdOR0xZMZ5S8gBn1kRPVWiLSzYD7uj0eTovDu3VJ1T4BlHaVZvJo+c
UEez7lgGVQwhUIlDLMEZd59kZW/OL1d5MGxJWDVEDdMdMWcy9BhIFEGQTktFs+mK
l3DAij/uun5td1L+/xkjYZkE0clKga0gTZRb4kNB4Nciyn7wffsHZoXGqRLzX+mh
DVJTNfSyqbG2lgjbE37iR+/v9WPDjyuZZG30bKWxovrEkO57Kh0KSqqQSya9q373
zWapWtBvdVxfJE4oWAp7iV/D3xGdz2mnnVc9IaNreNOqWQR7BiS2qvFW+EHtZw1g
7LT7G2r9T/2WcTGCCmQ29R3VKJkq8ziVsr5/3hcR0KgDCtv0vhqWFLWlaGFHkM/z
kcVxEuD5GFhkqjx/epcqB6EYL5iaNgiPvwOrZ/Und4yRM71cRANAdfIKNkJH5qrD
9WDO6Crxp2b7Y3EJgcsqkCbIUIwxI73hc9IzZj1E+j817Ps8N/qzk5JFnbhjx+oY
0Y7lbqKNW1Kfg2po+jfRGBK92/yQ2+hf1kegm4sSl88a1Lww6svqQKsqnLVnAIkQ
OYcUAh9vZIYkpaJi1y8kBPXEnqLxh1t9GECuNYqua6RAvGOsPbhzRql9rPc7kDMh
TO2zLI8gF83IVgO5gUjVDBGJLH2BJnNtknLux3/WvxEctqXo/baYJOj5YkpMsDSn
ae42/qG/J0Lz2LCGoKla5iomJc1buHdD4JQRW1BoYqBDbSuvp+sXA6ekESbPwaG6
E2w1nSmL7gszZ987BDMR48HhGjQ5wDSrrXbvL9PU4HadwxyOpenKde4T8NSIk98i
aYQ535sgyCBZqDiO3G4te1l7UsNWo025gT8pPw2bhJ97QbwKoj3KueU1uXCsbTcF
VJFGfRtw1oOe/KbUweVFYjatZHs+Y3ICi+A6cOUpMF3THc30Mdhz5DYjVfrBneHi
xELC0tUSlqqcAJmqgzHFTK9jc3gtPXHm0fE7vtQ8yptMUdb6R7SLy17W5mceaCWP
3wUGmuCAu/WCIsS6BxYGO2zhoV7p31nAvlHp8z0q6CMYOyHN7skrfWpjbMWtBE/E
17d9ag3GPMqOaLLLNsAJLjMK4j/EebKW9WUW9WxUD5W5OSpWU/ZLatvyfXIutO3Q
73ZJN9iuRWjib9OLssB5VSQ3oECbNg+RQqeffw1F82h6HegaBUbhSlPg7zLr0iwW
7oRtPt/M0uKj+uKAOMfUcxmJX1UU05qtrPBDY+V2bIQrArkYNo/+pK0NrznqvMpl
XFzZ08tK9/OO75291PIlzSeu4sC8J5IYM+oNLhPIlhWJddRR4npHM2Vhv9ThObtu
k8ZJzsNCBbd49SKF0oCHvW5UJrZT/RK5zOjRBgk0/W+4eyE/Qmln4xmJvfDqEjwI
f1ouMzoSvBhBBcs0W1vuR3eqE5r1ftbWh6iZ2vUCY1T+H94Zf+DB7xrHFh2ziOF5
tQn3MyKOnUy8WJzLxa4Ey2O2AfnhvhUo1Wx5KTbc5VI0Zols6BJI3eux4wQ2yT+w
tTgPoQBQqvysBrKiKTA8f51vnqqJKx3bTJXgJaRgYffjr1pInwWsUmaxhtQynyxl
lUuahBuah5UeW3Dwm4q0BH8MgIVVOXig129WOaUs43NY92jMgaF6RusDfKLgPoks
C21CIk+YPUKVfqBNycEsFgblHvrpWmBBlziTmvE0EhO9oGk3GSlb/kDWPYKwiyp4
T/9vNiF0niBuThWt/qkQ7z2VD0ngh9bHoi4XpmEcBTQpbX+tMlDXRZSRE51aeAYp
piy8A9kSg/h+chs4E66LwVBBFeP+GLcVRvcUFsqSu8LFosD1h8WHcAnyGs/HJ46p
597wecjHRlmYkCOVb0hMVA3UCvF5dMECLItPxoWFrznRO7A+d0HaVu2j7eCJnGdk
QygptttrAAMc5OryjHO+EI3RxQojwsf9jzR4rgENHO3hqIzLkWSBRoGUWDM6iSei
OIkjF5NzwWKRetKvH5zJ/R7kxG+K1sKizEwon+Ru2hGrVqFclgsKoaPnE3+Dau+r
bGK+nca+GMTDhTNk7XMaUKR/KZsk6plXGADt1m1X1HT2TQopvtBywWNXBExZX8wI
cbagK2J4V3EWIAJSRljHm82yHfpKGWRgsHVez9RVBv/WdD+8b39n66GO74NmYsxA
MwXdL4wKGdbXBUyKT2q1lzqLN+EUDr8IrlXP95udyDvFGZ5LTNI6D1dlZ8u0/pkx
iyhhlkvqb6oMcbQr6hJTdzIg9SFZYWxG1+oBWTM+jWRO4GagBOLa2FYyWLyZfkMz
pM+n/x7cXDVU/n8WEZ1HJ7NadmspmADUSrdYQmOrnd/MztkhmAgTyt1FMxW8nVLD
qsXBYyJEB96q0qTNRv4zCFc9ZpW8UAUySZv2MKDkF0sd8xn80rpEVjEtNpM64UEM
Jg+rXB5pJGBQL+OysXrZk9Fw6mKVGLmFyIdZTV8f4fzPB3sUX1q3L7mN9nBCR8mL
BJFABbv2ckCwEb7cya5duCe9VUoKJkweEC7MHhfVX73YJHdnrm5sQi/o1HeYPIfk
/Uo2ZvUY53xE3G+mjMV0ca1Gq5Ah3yAkg2Ve3u23yg9nG+2lyY9mX3fpNpEezPtt
JsSRCzw3xeZJZE0uPR+t5U6epJZSj9tLLo/kIzvQecdliTcBAQy8xugKj0KGUJBA
0MtzaB3o37ns9eOkaROrauFRSad7uLzVfFTOy7iIskH9KypBV2tc0vMrcWKqigKT
g7SXN+51gwjgAPe2rcqnr5GYeW0640X0eKUKiRvxvBc8DEf0ouT2otUHefZfXGCq
5drJxPDEx0IdZHXN0ZAq7/joQ04jkZ0CoixY2cHwgNT/la/RxhsHWRK8/9zndKWG
Rq9M5LaLiM9jz7khX3YHRzyfWESIoYRxvamQp9FnBcZY1ut9/liQMtBTDZq6Smkx
lG+BqtHXvjtQfgzIZnPJq6V01pPnh4rN9Z/sY+SoFFXoK7ZRuEi0JK/NzaEATegI
M1wQ80e0rPh0oWldY4AloiwsZ3J5uQ4k01MIpw0olQ2Qy/XqnsBASzfjk3Y+Ha1D
v/1rB89CI35qO/aA0Ey49uWnuf+4GCFgeguMz88QBxvW2sEzszJj24hJLdWp7hNW
nUajGvZ748M+/J2sI/LqDlVnO7fLJetsqHm4yFTeTcxBVN93YtzHwRxGLEEVJ5uF
0SzTYqukIhuJnMD+5pFOs+xJDMnXNF7qoQWSoE9Q+YnC4ixQbyiVbr2RKWke9zP6
cm5ZPl5AN0p3e/TwROQj/ab7+Yi/Bs7z1f72hYFks6KPCEhXpkIPmUXDVMCiCjrx
C8+blOeW2fKq7W6WE9YnYqibGzUTRFSpM21QSVF6wVhfCQ7ywrEO5SlD0KjBkZG4
1z4yDH5pBzaQ+4QTAp3v2KL1vyH/AG+gAPgey1SsO+dioSkSLIGXq/JvQvRqOhTp
+4ngMkPGvd7F6Z/NTe5fG7uGsm1zVSsRCDAGPlFPCSIyqejb8hoEjQ96rBPUyDso
YYsQINcnGV6a4s/OK1TSlc/W6wEyXSRTenapIdLHCNLjNNLMekOyrmJqxMdIROYz
H2i8uCNUZGx3DVL/sdDHX2y2cDfhb+O51nrCOQjNbCti8j3eF1Ju3O4viTSj8fSg
7prsgzx9ApJei6xk9vaMR+qKTP5BvlFKip8V3+ZrzC3A0UdMbopcPeoe2XQaAbTr
fv407V/gIQ3KdAbwa7BLVm4X09/+LPu8Nd0Sgri+7qJx2amckECU1e1n2XS74Sfv
i8agdjRloZM2U75Zq6shUg50ZjHWabOQml243cFzx078BdeW2rgjtvnF6uwI2aqD
iUtnP/enAlcnP5ml9L+Ha7qDvE5ovTkoqwmxccSiHXg2eFLEWOy0fBpGxgQoZnMb
ub5QTxTJEvmrkHEHrta7rYCBc9bpgBd+Jd+sSjqie1ZvGQiYl+aimSWaE/z4JxVq
k2xsbtRc735s26eSFkCKcN0ekPurOibdqNeRd2/UNSRajzH0VlwkogI6R4Wkz68K
QAnRLWRVdLD77AVT01HyyP+TigPAkcyyrjqMMFi+EZcberOKkAO9S4dlFl+9r8t6
bdQf4r4eUbBWFY3ZGwZ8ei8GtoK+2PrCGNXzbEqT5Q/e/OzxmspLnzycgkqvh+ZJ
QbwQ9GRHDXgSs4qVmrAT+GbeimBy4tVCEtkyM+5SMPC7IDxXtN8rIJe4hhcrNKbB
0TLkVQY9B/Nv5ITPY/fXY7+RLO+gOd8u5vxP+xMFjuxKGQnRcmT+92WxgH8RbIzJ
Qh+pVmNZV7Ytjvpft36hRS3svELTHQCvdi09fQtTb8PV7Dybp+SKa5srqlyVYB0U
v6fqSZg1ROVyB+sZrBJ3xgX4cvhV4FUEoQ0pBNwhi6ZwocV45T6h7Zznjrzip5Rh
sPKXokDFSHF649wSmy94V8/HV4WLw39GUuPbdjLfP3UA3SQw/js2+Ro7AfuVID/6
OrNP1O+Yt8ybPioiZiLu4CbRv/6uOfjLdXuk51ywCQE6GshmKyNdWcFrEarmaXXY
aplilyRegyuoSRID1nb39xYgQEN8Asb1UY2EXgfHlRhb9SQKUR+lrfEe3OCHfpei
0x96JLVKNl4eHRber2LJHmEZuR9IYwui6FucFLqkmuxeExth9r+hgoyhaPOzKMrN
AXqJCVkvqT/J1FmeqSeCibfQs0YVpQEqWuiWzr30ZktB52l44KuopGG75KGj84Jc
iI5J04aLPFJbz9nvyjUJC49voMJdvqztG7YGhVdn7dKlOMhd3Rb4mAr0kR8duq4A
vzePAHNbOJ2mvslWirUQMPayNBI3EyFnpsxMwzLWgMVvBrULE76zctdPFKZf64rs
8UlFWQ6dSSSu6F7J004rLxsTnA6MKL3EueH0jAUG+k6vxGBbdiWUP2EphbcZea5R
qqwZ0NfQyRJVTaRGcKZY8cHC1X9KWk86LHePasQEZeZSq2+eS1PVdmUGu6l1S2I4
eUtJaSfhRWBzJZcB7W6oQ6NjueRy41mDwhGfc26ay03urk14RSdLQL9qeGEHSm4S
yG4NPivytLWJu1B0o23n/CFmEXPwUrkRB+pGCiEJOLSSTTlyi/HOZnA+jcMpbCq3
WbOxoy2hpR/rIVYjE9XY1zT9KdDwSJfGFF437vNIAdtuH0zBdJLoiJC/n0Rb3+E+
2PgOCEbPnncRVAwdgm/MZqqvKLdIPSKARwRJLLzIsHdl7W6xLRHg01XbwrvKDP1B
+BEljDJNqXhTGiFp22rBJWBZnxQFe5HdOPTFUX5aWUTgIWesyIZ9ldQM4Qs29h0J
PhnqYnuVTuuaqdwn7XSElhFl7BkF6ItYkxc2omsmZyWC00QTCiXKsPDs9kWSv0yW
tGf22BE/ymoFYdxv5nyHF7lCYEXR1sHKo3naE1Y4Uj+vSB0axQosXamF7fhAz8DB
zgkANA5hlECOqHkGAOCglFgQG9aVCFHqJEmbpTseopLHSW2W7pFRoSgcUes7T3dt
9NjbZcUSzCIPbU04x4eJFGv6E/WOl1b2ebVhAB7Ovx2/y4b19XXXB6hCeXKqSIwQ
i/Q0YJfhU6HMfv8C9Oq+XYPJg9/RjUsfOaiDHHsnnmnrhAj0B1nAVlhc2JTLMcuA
bxw+WFhmhPldLSxkWPvc8r4n4uqvNHtoMkj6wwWoxtnMXNDYwezy8mnCbc+CPxSj
i3WBjiAJ5HPU5FinMapFbXsdYpB8weyvNhjgSzexsKaNBjspe4Q05DI/1+c0GyzE
VINqZ9wr7zEwzjhrj9UdlW1Bo0DFg3k1IvhcRcK0q+q2C7HihVFgCemWc4zDFz/m
TvaLkrEXbOJPmiO0mSg65TibJN4fXUFld+/PUXCXut9NyXdz+Lhwh9355SPpHZEv
5pS2YsDgdAZjreHKdVapqJ/am+ys66qrzKoAYxxcr2WK7erf+gSof+U+StWp84E8
HFiP4AzIobdQUYgn7GvhSwrV/+dpgcZEg5RqsSnVkmhsuDBXhk6XROj44YxSwVoc
Di2CNg6nudvAX80MvHfdAQkMMYiqd4OPVtDz1hYocibAxa73Xc0oJ9Fayu6Pn1C3
kxl/kH1QHwLWPbuESXbak2c64TlzcAhBaGNh/EG7yJk4IpKABdswaY65ZPIhmmLv
rWFMIIl61op+HK7kE6eEGA48Dj54GqQQ/QGHxzG83u1/93KZkqjnhs0s52qe9UUm
+GpKJHg0ZPq92Q1R3x5yysh9HEuLy4qBxu26ZL5DeifFHHJquhttqv8Br45Zm8Iw
C/rrKq3shF9hlMoStyln8HzQ3LoiiIYYBt09yQa5DIDzykU99o5tKeCWwmlufeIO
BeG5D/1r5OOLc1RjiNAU0XVgVDJY0LS4ULGzCukpqGup60+uiBGcC/XW4hqDve8R
/n/Jl3RNOmbqZSsjih2C1wQ7ZgW1CgGLIMBcqDybnAF1O7pLcLA5j/Dm1NFjHYr2
4kj+JRLkc7pzMBY06O42qSxym5wpCMkwS8KNfwB+K8hRCTqUBKo240NIQsvle/zM
yOtHGNErRx9Q9cFCNNXhnDJsYv/asDc2SH/pXZbcdPPhjS5sj9IqecLBV+hrG/l0
ZQgn3gi6X2Z1UmjF+LorkkIYaXSrGXE0eVCxSDjmSO8zjeTatXnldeDkbXRyB6kt
n0N9824d6amQxCfz37wu+C5oCmSwszNktJ8GKgonpd4AjIRO88hnAHwXAo2M9zOz
5Oax2lgyLaZ+/CaK5YFMkBYIW6eC+b25iqTFKtX5ujRwUtwlZ+Q+nyU+2qJQp9X9
oNWEz3dwGjbOU9QSajMzNI8LHMG+5nnK8tIDtIbWABM+H0TJ7nkFyP80OoHzEMJh
ucF7U2bEz+GHlsEEC7yHwWOcYD6Tw953fFEk7LhRxFd+bQ090uFwwOhK0/hQ3iWU
wU7n6ZBYsaO+d2q2BAlmD2LxE4Y3WlS7kf8Wcmo0calbNIJiYP73hgq4AIxnxWST
PUQf5gkBXnlK5VeJ2HM8oniNbqwDOhhKyAVeIzqEkxIIRc+wEs3oTn1Z005kC0B1
XcX37bp71TnBfRajjU3auiLpWvdZWPT+7dE4n/ZpyvCkP/VV4eOO1AoxFwrsa5wo
1mp5cAMQfA58+wKJ39trf3TbMeEEG3DZosLjLAy06f8d3URgINYOgF51e5dNij9O
u+iQusukvbNNH/2vJqr7UcCB61DMLI7B2R1wnsNtheSJYY/yoxao8McGKFfGzGLK
YIOP+zhcjc4BcOoI9g7UzgL2YEAO/mYlfUxVVTcA55TMrc+9FJSFTQr4TEuY6Ayy
rSs+P8K+AOH9/BEPeQOdlCAS9Bx6vfVVfV8OKefNS6v52Hih5sCGkqSPgrxJ0k/Z
/Y3N0mP+CnICwCRFFR06T8EpTUJPpnFiIQOGI4ZO2As6f/gAd1THw1vigVdIk1yZ
Vu0d6IQcoBjSbi4rg/w9BYjZGS8JYKyBKfGtSlC62zWnLPxPnuvLFuFb6PrIyIqH
DLKlZta5eJpBkVCsX4rm5UsyUWAlxw3Dp5d+0JpbgIapUEoljvyoLcC6bhst7CLr
toEbGVIHsRXB/OxAnSe1fSAHmg0TQJdLg+ibcfDIUWqDbExfcykgTNlYioavFViI
y326jlLuCApVeENqcgA/NkLJeCf35HAN3Jx8T+dovKxvfR/gYzNsnAsDRX1kr99L
sIv2BaTyhjugSWMA7XBBQL6YWMx15gxQo3uNMKuS/LnN8eYtH5AQnQ0YgUS42BRS
Jgc8rNgT7vS5vTEIPmQVwtn2HrAMP95MWj8oEbtGVVC4ODlkt9EiUoxXSzc9vDFt
Z4JPGyX1DL6ZXUrtLjTHCIGbEjAy3mK/Wq5bWUwbUL13f0srWbgVh8DUNAG6m1CJ
3vnVwGPefVtx0w9qgGixU6XE8Z+ADbUzfEtt+iMSUrXNhiIarICte4VVp0NR9vow
KyknQls9ihKQCXfY6nhaSpOZSkDtcT1UNRI28Pe7a0ZQJf9kcfFrVSCtAG+5SakY
tPEVWdrB+933vjvHcQLkzUz8khv5yG3zumphftCMgTStJp6GSX7m+HYseHRcSX2/
h+j4iVsaSmkFtqjDId9Xsom5+v/pJrLiRGEUcT+akoz9+FNfvbBse+Wp0HVnxz0v
5wxjUcOoPMtfjo0jwr71DLfYLgholmGws/kSgRYlj+t26VfAOKCwsQawnLM26Vb2
iZ/YlAzrUnLuKBAAiXUiDlQ6VYFIlZ5bb4LfEoTK12XNoX+Ihd98ORMRNB2GLzP2
L6DuqPitL/qCBr9Naz4KBHCwHOyJg54amtnyFjzriW+LqRLR5/OQsYP7q6XjN8Pf
9bOeTGpWc2eWZwd82hcqyrhi2O8lE5riy348WwUotvKyWWH3r9KXHHIXbAtb5b4/
40NhHBcmCDj29KA9UaeFUJTFOR7c/PzZQNhPziyi9VQid3B06jZYZSTEsIBXSE+a
XeGO5bsxWVzw8ZkoGcCMh5JvAFJByQ2jnXmH7lOlvEfH+vlznaUdkIGvW049TVh1
buwbDyKsVn4MDPsImuSz1CGmjeVRILUf3IH6fqbH7/4kLznnr4WMqJdM4ZcBwtls
Q07OMinl5eTH8bsiCUilrbivOl9K10a66pSPjN/m36BwSvfMYI3PgJBj6v4m2W9P
oLTGN4K3Dr3/zYw034KEuj0OYGmqKKEBRz4XE6WPL60/5yGWIw/JaS5oASLy1pFy
HODgsEOXzTWm7+THO6qSJyaY2CnOzT+IIfA4o+i7EyzuHR+cRsxtlXAN+pkiMerH
J9MTLA6wSUvJgJxCQjxwm5K+O3c82SQKLAypD0qH3LVPmwGu/BwK9sIbhs8Sv7mT
8QxTOBEiEA2ig2XHvHlsaX/aUjpr0hqb8vtgzgVyYpkfVl6iZTW30FOcQCa8dODX
VVfsievWtswgxZA9L0BNobtkDeWYvK9FMFr2kE67ddf4jEIOl1CigvzMUP4fh/K4
04ovyNCfhtTVNmgbixoSkOlMZTheXc+9tGb49IZnxe+WY5I0ImeTcclpNX94dutf
3BqPvPYBPmxS4FnHqeYjOLhi+tMsZsHXEjtnArCNUsSwu4ioJBWx1OzalZD43pr5
pDq9PNypd+ZVdkeup/1+dACnm6b/jda0xgiIYmmzFN+CuaNQwaKK8/AEUhogmxT5
i+PKCEiSO2xkX0IOwnlG5detNnjeth97QArtLJlWuqhPY1Ke4utWa915OjdBxogr
WlBwyST49Xbu8K28JA6CAx3Oeb/VR9SkFbla/+K/XgPwN2Uuv32jUAgdJPX2d2ot
jN704lw1kHCbHxHLWHaVqSz7/VpLmdbsaKejOa5ylaPqH8uiiPJoPrQv0bxe6Pxl
eSpPf8ZpYua5qSJQAtCmDqEB/u+8FK12VfjLJajFsfxR9i3Klfwq2zUayQ6krviM
Y0tCg5yU9hgvF7+JzLGCxSHjaa8Hg7NfAdXVCRNwRdBR8viPiRFcgAhGWVNEC+bY
lswzhApr9qygXNmGAWeTiLCTfgPnoTysVQG/vllh/u5XoyM4FhdOkWd/St4g72AG
/7NoLetulYToIpkcXsGIdu1NYr22e6HIgRLWqNb9kVqQL5DI1hVdAHfRyVllped/
rZiiREJILG8EeZkTt5OdKmbjFaLBsSYguQXFgLVGfh3QCIZ33/nAcMwDDimdj8w3
sBmYmXBKvJrLNHcrhvhRTERsAVZx3e6uOOTNzjny1sDRH7eSI99ntkIPkd2o+gu7
7Y4dMEBgOH+hTTzJOrzAV7QaJfZdP3AwInYo2xmsYPRzHks2WAEzlQmknxaT22tc
531Gnd583kRyhMgxRcF6pyrOl9Yjsge5cqYZAMStIAMeJtI9R7j+bze85lLY9Otw
748b4t+BxIFzxVRH5O7jbxp5jPibNwUfh/VOaVLs97BtYlmvxk69RJh8x7HIpg5Z
X29+8UvuBNCX4+J7TW63GpNVi/QvunN0y4mx9d/MtKYqahnK/wPRu5ShM4OWbRO0
bblV+z5rUYTdstNLpVm36Ms5b7+VILwhcplNaDTA1qKGc/aZjBNuirgHIu5FrG9t
u5lXak33N/MzolCA4IBvI7bV63L/G9jCTxcZHRUjA+5YM49/2Pqy8oEyLcs9dmJP
vstdTJJR0YwC5l3tsHfZLvusfgbwOMO+OIZzLQQ5ZTB0fRaz+WnODjkjK5d3nN7e
9VYSCUJ+GJb3+lhv+rGeKGMn8CuHwgdKpzwKts150Dj+pJC1dPg5YA85ByMs1TUW
IBleMoUvKqAnKvJCVi4FO9VP2jkt2ByHFyDwBxe1Oa4OHxAki8WvX3F13mfzZ2at
Bk09QWwofX0aVDp3s/m12Tw9rnF9peG2LnhC7FVVylTB0B/1VhA2KnMhhFAyDVZJ
6E/J7GDI9Nngxok5vWokYIPzobKeTGC8JSfZ5PSQmRS5oGY1RnGO0eQBoSxpvlre
+eG41xcxJ5SoZ/Akcziz0siy8TFfmxGkm7CJQXjRnD68r6lBHqTvMFPCj7fsoZDi
QCmyjors+Mj7w08QvdsbuRnbKTilZh/Bd7MndTHvKEBqCTJC48M4VJ1AGucpVsty
3SJLbKqTR5GmN/IvIT+hgh80Yhf7e34lrEYwW6Lv0sk054OWcJA9imip28KIUPBt
9ZlARrXKXjM3cSNptMKzrM5DdsbUgzszDeIxssQBOsCxT2hift1cDeWrRvrDDdV6
2PipWSxMx0DPlIJJ1nSv6s3FUBmRhaXBh0xc3lEdAroM5oW+ggC3wCQYAlMkRxfU
VZJKLuV1wlOV2/zu5ZMo5ASTEaZRxFHtMrp+bmvEp5UebN+bBPjHLbdyI7f9HejX
8QN3pfwGslc2cZ2P6r5I6m4IZ0SBexT2sJSqHK/kcazptHPyW6Hno9+/Od0pZa9O
So0W+6htQcmktRxT0tPzMRwJWqbwFkDWOYG/ivn/1TML9lNX5MDpnd+TX0A8WAUA
/eQvoRO7HbgjWT3HmaCKx7Ay1KdfZF76ZfhTMoqaET3xeshDA1xXg61xOU0NlF+L
3TjyV3mHKKzl1nsTNmocq+gpqT8b/lnk6hWaHk62iao9PhSL1jbWToqmxH35Pli1
N59XR0JrjkhCLcVBags63QgLDEvl4p3LZkAnahpIGlhjPdEZBnt2dUYqglrT3/Lh
vJ9WYmC4mwq8kWi+bV+njMtrxBx9cu2n+915VGdlQ9xuevju311OvL2zVYm+X1cN
BlNRJZWIjqRNnG9p4Ur1BB13BdW3FHIou6pfGp3gKTic2aM0C1mNFjKq6/U5wzo0
0XEyCSXFBswUPLqaEEb/SZ0hUIl6MkAj99hLlVDvtfhTeJWoGMiEoR5LVIPwFFDj
1ya0/1lHSXZ4xxlTRl4niJLfrjfBt3iPo2LLAl3FYaXpImJBA2XD+C9ocD875QcL
dMhJfGJ6ne7HVoC6Cl8s6Qcjv+wj+gGtS41gNalxXIIl6OLZaWRh9qwKn0FM3j/9
fKmFzMG4rLqhWgp0LPjsNF5vHOLkZvxJCVZELAgt6bCSAopACgFyYDmqRtcH7MWz
CAruCF2E94qc7w+f+ZOd+GUIz1A8SjfGv3l3iPgZjDBOBQlZ1ZiHmzR7qzeCTC2P
Y0ZSQYz3JH61VvT5w2VqGPJbieIFF/D80Z7WA3+WFgO0Cc1wuZCy/d6msxAJ/Om1
myPpaWgppa8Gyg6AvqusizzVPyR7flBYOBn/YryHjbKIYCqUMnU8+0f1lUzuOfzU
/knao53OWe4wjN32PCcTNKSaMYK9p43FxPSXLunbQbKr6ZlP6txoagKWHAvc5EHp
qztCo/CG6DGl9I2c/Xhwv+yN67LTHYxVXF0yJkRHBqkaWyxniQX/+eEhzBIiw+9E
5anOCNJBm/m7ZXbv9Ueg1C3eTAbVohDl69YZMM3EA/2n/kR9QMap9vuwZWiTirMB
JAvbYBHVUDo7Df8Jt9bmBJl7fvU61PxuIONoymXZhg3uO1XPslNFZJ/0ymW3ZaBT
jf0gX2rA4d/5nXgQj4rGLkRochFyS1CzYTb5Rb4cRBTZTI43M0lIWIuF6HUki5UL
8CjkjxJv+AHoHA9WCizvWo2M2grDDd5qjSz43ns3ihzrFX/X3+ye+wZJWW/slxos
B8aEeFgHN8mqZNdyC9SiMnUJSQgczTU09hsThVXmtkyvy0u19FU4fm6O4M32yYfH
7HVCJE8037nP0c0w/RrSgzc+qz1KbY8+PNQ9KgpH+K5rPTlqdACIE1FrJ975/e5u
/uQGN2Gx7o42Kfbqcj62aDNLOA6KE3Mmo4PMJUHu/SBSosq2FT0WIJ2+ZlhKvLFp
73UMrJm4uOjdoid5Rv6DQlMj9syIv8WbkLJodWtq29aEeBsggHmyjl3mT1IkYdEN
lbwL8q4HDAEY+78BKYi5Jx3oUrXCcr6gYa3NnDz/O2XsTY91YdmEXSiC5ugIM/yX
zySK7fRGhnIdVS2FPmlVCu0NbIWMVT0X6bA3MMwPNUtDSXhD0albv+rkUVHHIx+o
KNHYr4HKV+9si4pJhu+/OPsVjLa2Cc0DLUzmiBahGRHvNn9OQEDFOOVs/F5fg/S3
VzgQgg9PaEPCFRKJIm+B7E+1vvdLDBJYTh+pBkczXFgxu2JxX38B2tnY/C9UXuyZ
o7RYAguPhVfYC7wTBnXEUtuY4aJmMGNytsDdEqz6sle8RVt8d6zDfV/niky+fGei
/WZ5MXMLpneP32/9Xa3in7NHe1Z8L0Abum/VnPyfo55+R5umrcp8S5c3dt2E/LmN
XSj2w2P6ySVmOBayO4Jw28IiNnag0K3W2n7naT4xf/vGL8qqm3W3c5L2uBA74jv1
BKbfKVxK/S1DrMc3boJ74nh/AmwQhX5I05V9HhvfDMtlU9DhA/Ly0qgyRllDUzMC
Zc1WjeJStKqtVeidG74BeMFN9tXjby0uWNyvFP8rBo7ES8q2z56Kw84sYNN1KUpu
Fvpr7/QxdBjOxq6hotoXmXR3qnbkAG4M/wc9pgPhgU9lxSS1A4ZZyTbvGyosj7qI
xqdfLQvOPh6bwFTXy9q/rKQbRVLWDn3zFEwMhYonQpNK/j2+o5DWF4EMykLEtdzk
U5UvtPljTsDwzp2C70E315O+jK/v5x+DyR0nqU00s2DHBspj1Awsc/MGYh5Vlm08
8X+j2VhAS55UTL+A3USwG7dmWGM/u0TAXuMGfoTfuEiJ/Rx8Z8JstnCysVX+1wVp
J51KIwkmLV5OlqB13wb8wiml7BaA4yBz5sn3D+zo5/BDb5IHNuAsyjzJifpWeye4
oTw0VNveWYch8cb/HR5SIpt1fa9BcJr4JajJzqsKgRVf3W9oI75uwEFKK1+kqXLM
z4KzwM9HEDAhF1YGaKL6jiC3+olVjhBmkgHI1qhFMMGF7a5cRPWBUcC+LGDZoUbQ
h91oxePuJbwNBozCkOPMTVbZP2K0ZXnnC4zuDaaj2Z96arvhIVsxGMl/YSXyI8VR
UvJaxctFWpzpIsBkxKwjwTImHZY2MT0bBKSCxwb3hz554nPE6LNJiZbEo+06wwS6
KhZIpPAORVDtOjZbnvvkmZTKZ6yX+EvBO1C+lbTLiwSggjUBIWKGtd0Ev0pRg/Me
VRKpht9qSgqM5Q7Dm998/BNLlfHL3AU77GX4B/NtWykkGWnvkCaIUlsUYDZGvZDh
iMt35x/Jt45TBfuw6a9PU/QxqBYzcW1ZX5aKNjtBVshN8JniIzQ+N39nZeKDmMkT
1FBL5Y3tQfEXJnNI0kpIlhIXE1mesDvxc+WDXB2IPo5jnm3KooTFCeLUzPJYTHRn
rqgvhF/A8V2eD4v9gSzjL1O+3uQxTpcNA99YeJB71Z+r/UsYEUtdkkES4Ew/TXQV
+qwrpZ7mEYEu6B53nspn+7BKpzIxNqQ21k7tgzAkNKdNmifacWRSisagfJ5qVUSD
KB+rGO5QBfZ1Wk7Opns7YUEX0P+57KpOaXeCQaCkTBuq0gYE7LMXfqjqKwd6YliZ
yRWv7+0UEOowmlXx5kNiV+vTvJ39mqKFTBMhKVdjnOmzOoZLBnigQXzVhbmHPN8C
93EhXDPW1ZdHEOmFTghpXKbeZoCr4FYeiLuXQgHRzflIYGdbjqz8dSjGicMhiW8Z
krvBBnDScohsGQM5AnBAmqSSX5c0sflKnpneb0wuWZjlu8jRR1UB1xlyBSWhSvUG
SrHDTXSc5cOHtKcka46lG6SPslu+pabisDb8OO2+AiNVT0HCcsAPKyAqKZ3uUflj
a3tQh9TnY43HNHDNYrPlUKYWFPzia7aPVMLNvO/eBJ3VAz3ylxRYEVy5t0o8xHV2
w/+OrpGhYRciCgO8zn3XuwCQBUkQL7GjNdLDROufV6KPUTvBdW28HV3FDN+qshPR
yrCMg/RGuPe/zy5J4JZZr9Okik81sYguoLJFwkmXiO0ynOzRu5fTTx0NDMyOghjU
z25J9LohiPrf0azYO8Un4SOoFSFginH61dfqE5dWzangNI1XKvGEjdv6oatFN1c7
dRPIl5EFsjRfrniMR9PuSr2tYvgqD+ObAkq+5SNd4zOqsYYtnQ2j49iQzRO83+7+
qu2anqya4Z0/5rXKhmWoIaPi2AhzAAFodNbRXJWB4CesxCNW8F48Xdlsm4FiFWAR
Fz0fo0e1xz8GT4qMUluTsnxvbtzhzkM0C01RbW7N1a3KSsJUAe1OkKyVWFweOI/A
7u8y1kMlPVKqMwNtVoDJEGCxE7HT9AfT6GE6PJSnFEpNgtWgeROajj56hpdF/T56
CIo/LIf5UDvM2/+uLUf1kch4fRmXPfFbJRfLsIgXAfHJzoH57+diZvhXwM9oCvb1
B6/HF0vVVUe31DjSLWNUCkAtXLz91A/J9RLf9+QtI96pyUeLy0EI+qvOb/FpSIo5
aEqr6u/p3/4isKMFHx9VJn2cquLouMgROye7430tq4DcsRviAPRscirKgJAX1ChW
e+MxTC3CBIenffW8Mr/UAKAEhUR6TvSjtT1JKRaoHNX+csdAZhVNEr64yr6Tlq7P
bxcaysrYKZ6FEb/qDiicscFMirkw6zi0bl6A516Vg2u9sHdAEnzNhK0jpS9R6hMB
SCx1DyM6EVnoPjfikSK70i1nm02SdARqTRh8JeVrpEVGk+aL8/GdfCymhqSMzM6i
KlXIbATOYcEd0TBTzEEq58Q291+1dQL+zI/qH7AtmCHAWrhxg0wif67kx69R9MR/
z+4tfr2WQQh6IZgMPlBjPikanCVDHRo17P2uLCPWt3OgL6G993wGNiau0PVmiNTd
PT0jXYIBEQFk28aSULDtAGw391dJDhFYq3xdqcD3T///yfozd/ebPgXygLj2hbxl
T6NCjczmV3Z0PUXX8GjB2ZnFp3tZjQGYdkgZzN7qlt+yIQQyl4EonMdezGTQL7we
wI+yZ0QaU1fKAmivYSxoDI/MHrTC3Il4MQ61Ch0LDjkMM/dTOtPrH0Q6vmR0KEoX
c/VTpYxuIEqTlKDS6uuBfql3XC2bbh41meLNIfnSvfE0IwI31GVS/SsXX43DkdJ1
xt0LtGA3YmjS/H4B87/SWAeTr7F/eaiCijQmK/HzaoUIbaTC1NEuJBQ73u+bVNx6
CfFNwDGisyggNK/jT+YqaQ==
`pragma protect end_protected
