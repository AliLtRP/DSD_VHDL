// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:53 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gG/L0Pf9vlnbMzfNEZIqgEBgwqTbcvp+C1p2wd8T9Hry3OrcxBWsUkrltGi1AnyE
TKjinHCMiR0toAv4yNHQkl/afNQ0fneQ7TU2PNPmLHqLYXMbKNzMyYmwvdjuep1C
Zu8XFejXwL4DCP/ibxTQ3Y8hI+MkUcn9i+07PZBBFgM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14000)
yjlqIf3VYAgwbCvjCeTCAmpZTX7VQV/M8xSI5H6E8FgDXOJSHCiozxdVUA5hTDUE
RS/l2qIbBtYBqcKkKCmApddR2bel2XFeGu+Ve7M/t59uUdxh7ptyQJRiiWsBnjWZ
i3TlZqTpvd9kneqYRqIv4ihgflFMpb1aLB2KA3pC0ERzihzcLAIUuZUQhm2iyTNh
dLqvbTijatGPIspy3C+9sKHIWqGxNJgFlc+gUYqqpDZFFzSUz1ISnpwsQfzygrEN
XxjV0gjeCbDIPC63FyagFoyW32Se0mxSwVdfe2pSfCCdSU73uf5AYfH0zJ2FM1zT
0QeYrbLwZK3gUfySbBWI9wl2vjqU9xcclevsupLR5DFmUsHs2igg+C1lHr6cxP2x
+Tp0WYxAyoGgwyAf5wkaRm57IshuKBqo0QGFlLQN9s/X3SQKoetSQbITkAZkkJE/
Ym9W+2hVtySwuc2b0htpUuq956wbU0jF3lAG8irrUhZK3EkY4mI8fmCfldC8M9+4
2R9o5eqbnPa0NBhdkj2RKz/OU1Pr7FGA2OrMtMEhMAMVhSgsE5W6TaOiAI/0AcFp
rgAx0vA1Q/km7bEBtrTVxixvKV0p2/kFEhrj9o2tasRFw8jpTvT0kAE01lzAmKVy
Xv9u1Syy1m2795OhbC3wOjWBIXrUDxGScBd1of5J5konlLqEh+cNO6+XPFAPRE8U
n0luElMuo6PSKNM+y18TpKfjdJvdgBEdIwcz5qw0fu7kNlaS0t2Dwh5EcDq05h4N
QJhBLuaiD6jnAeE68ggQmtkrGPH1VcM5ne/ct/1KrGM7f0ftVSwOSXQFK5DF6R8g
KV2fqvJp8AZmHV27vtcfUvW2xCYB8dd6IOG4dvttdFe9RiYPq/u7FlMQskMohFuN
z2Ehhz2NiIay/n6gV3RGmE6lPADY+9CuxwwEUeM3Yz3hyWLhpjHtokwb3WM+MnHV
ypgtwVtNTs4+Me4fIm3NnDMzCK1f5yNH6RexR8bPA4OZEnJhZzswfa5CtWBdfgCu
b9YSOVed/N77LFPoFZvwFz6mwvt0gFg3naU1azyxD0ktwgTKeNw0XmAWExNdNbWo
EgeTJosQKtjrJVNFIcvpbct2El7eEDVTYZm8e85EKl8oSQMce9E9lkBl1rUS7ts5
rMJVow+jUZaLbpn4N8O9kvQwOSYkwnC5LelH4wWRTfmynRbIRHhZSMaqyIhMVRYa
k5MjK+he/uyN3vg5CiYcAWqrflu4/LCSxRdfhA1fw980xI46/MIHddKLe8wDppYG
5iiqPnkUarnC4TAgYUWlNi7WjtM4FWofEIDk2a2j68oLDnEJeY6G9DBP/MZAWZqi
cC+6jMIEAGJXT8tCje9s54E/ghBocuNv/rhfxbZM2qj19fYUdK7PuSLRuQLhrHNh
er4DeO6dt9+gVg28SGSLuW/mArNi07SnPcojguxWc+9RkCYg4Xaybzx39kvQVmDF
D79PPF3yeMT66Ehi+YWk5EY/PSzGGNlGG6B0908GEVZzW6LN6bs/hHd+IGl8FZj+
dk9h7f4N+menVDk7nMBiRqtxwKdJrUSn//R8VgBcnS35S2rrqli21pId8xMV+KKJ
gmzQ8NPFgU5qXhTwjcyXRiTKj7ibSBGmBgOVd4Ct1/BXZFK8Hm2KAxG+pgqrYAzU
POZsN7IRBbhxNiY2ZxhaPiFxDO9gVy4v0n7f96IUSbSRUqZQYvP9l/O6NAe4bKRI
d5UROTKq/EpoltsMhO4uWBX33LfQ+TStlf7+hZVskFPIgaBhIkYkb+IIo3obZCO0
jfn1PnzyDUFb3bvPRIKJ9lahzFbtqr6H88bNtawiQDqL7LDqCNQhQBdSLAezNIyB
f0faJxPsCcUPhgRZQ7A/PcZXgYM0q5XB/jZiihzhZv8f31pXx4ZQu37eM8oDUyEv
r+1miDNMjYgJB3mDfQErKWehmbJXJbtdKTFuwXUmyDuSet4anfvv6wAN3Pq/zcwd
KrfGyHbCIVvGVQQmELbS4rYIDcjRQuxMjr9dg87ZI5mI794xv8Lgw5+428ehw0Ux
ihaIR5EKswX4uxsTjl+rX2EhHuJ7nsdx991vOGkKBdPv2rvaQIh/ByL7uHDZkSJv
qtdz63j1aefXmUKGaF5Mz3dmM4M7cipc6vfGyxLRIP/gw7xR+rAgDByXEYpGNF0j
dMSVXYaFtmwUpEVRjSLr1EfZmalSh9FFMHbYSL+3stmsLiyUFpEHG6GkzpN6HxnR
dFJ2SArCCKqnq2dQ8SwTxZxB3nfMfv2atK4Ccdp2lUJhlQ6/KnCNb2HmDcopIjCT
Bg7063eh3MfDq2QR9jegpEzElLwJ2ZkJp0cuuglaU//hlDKT6wFBECru26R2W7xh
YK1rz5h9pgMltizKQCXRir7yDypilWITzvns/tLKRzPVDh8LZaz3CdUWC+nQ5777
Okibcy0Izt2WllEhdPNDmf7ODsh+BQJvruf7uETfyoxo8T61oQf9PARHzGr+HorD
GFfXxg4fwAK3f5Jgm32FB440hwtArGiojV8TsnD0dedHJXiq/NY4aNaaaaITFGdq
bqsGmyU4wtlgl24b0XAhfGoqUtAET4r/kKLb4zP44e+pY5eMJdJkWT4/jUF+0rwA
npyl2j4GGGDgh8MfpGTAtqD1zQmcmJspjcW5Fhn0KNSrdfnpIgthMjHA3aSI1V2M
+mDabGwbrbP/tXOcsP/A6/3VPlTGugou8dE69s402oSbvP471sNsr4vjuNWD9H1v
71d07do2Z/BX48yVQ9AaNbahG/xdhjzv9/3ftKzCsu1WEAAoB4k7xWy28P7AYoIm
ID46S68ElfgGIeBlOSb91FkdU0XmXCXe3sh5rDlSX6sp5e2cZ9sCFYowPkHszdWt
dwfOCTLQzU9B4sE6SI81FL6TEvy3HAqn/9oSjqWX4VnCrbTj+Tq1Xi6/9HRzAqy1
2IdF1qezzq+5LGQB0X9hmZ1VHeg+J2fQxgD7AbDX8fZO+AbjKsxwcxB4xmJa5GZW
EZKzg7PLUIhv5AtvE/RjOkzYh8Z+nl4fQ1OMcrUjY+vv2qWLk770Yzf4fWxtwNxA
N2yCxojiMIb0UAL4H31DMCu2EvLKiD18c5sVaP6jdm4gA2s5MY/vPn6ss63NQPac
3h10BfdUBmcjTL+4Td9pLYK7GaWQDmuce0gIVMhkFItcbhvSgtwHfiW/aBOQqThb
TisIPrrSjMjxZH0FsE7BfhdfhI+E7RzPhXEolC6nNhhoKkPapI6PkLFtoMtpgYKk
HTQX/s7EVPnwQ9+NBkpSUC4nAewvKgqFo2Z6E2HSx+t/8JJOt3gA6AFo/iu5kA07
OpnlqvkzMX6TrJXQAnKPj0e8G13namNXw7i7EzQa5oYlHSPp6zeR4wCmzUE47Jrr
jEdn8DUeULPF+sCPmWg7V4MCvv+5ETTLiSRyBXbMTHtBWw5CQkS10UiV94t5QI7v
b0jagvBQZabZ4nZ6IBsa2Mflf5gFAeksT21wUJjVKGHBobUw5vsed2f/C1D3urC3
pu05Gd7jO2xCtFqpqn/n/eSEvxQQJCZWXJNSSIrZDTBq87NsUT0SSmGdT//P7i/d
yEf6pkbxBzclq7DzpmWSx3bkS7eur1EVdxKYAziOxEJINOWne0PTjc+6GkN+ROLd
1fJkwN3+hKtlr3OYA31n/TR8uC1NmDQJ+fQFEM8wQPXnV9A56cWSZ5HriIPfN307
Tu0R+OkNDI7pdM7vzbLv2AdsVxbKRVKzzq2+8lNd5ZrD1uiYmqcfGtr8qcJoaDCo
cvBRnkyDTlvXOfIiyUugD9/BfA4doDP5UzvnfJ8DIOApAAAIrtgZhMyVtF34/zX4
0l01+tY/LWlqP0SHH0snO8HtMkMLSNpKTAGTMtlFAjrgJCGRT27JjuJxMrUYa83F
YSWZB2A+xtNigElwIwJgV3E5oT+7vN/BViRuYtBwNmIJWhfqLdQV3taUQNsbRuzN
1kFCZUw3iEUS+caO2lJ4qn5yZva4/pJTvUz54fVrg4OewMOg9fn9mm4grIwPevjG
dKNBSxdQN0VodsjR/29N/qOL6epFFLT4nhbpYI0YXBKxhqYrvUhF+BVIjN73Zql9
XxM0tHElYyYpD+0McBTSw+R6k0If15NAWEXu34duOQBBOIqG5qAEyZh3vMQqfBFO
3pQRtgczhEmrENc/vD2p6PGDPttGn072UBsaYkT9HOTgeltFnecj456pIVNeThVD
to7J6EUxBF1jrIaQzZNvIqzvn/3H/FklamdQZ8IvLB08EVasHXiL1rSnuO0tietq
qwvpM9aibVt8myvc6RmiUMM9/sjY6WzWsWGkQKub37pTj7uSRIaO9AaXwknpKz+R
O4XIp9wMTfHKhh2RR0pM/YZTIwpCNWVfAoBWQxAeT/NbAjo28VTciwGjOKVCchXA
KuqPZX0oH5cWx0n0mlRMbSBqDCT3er4NgB7LJXFLGy9oejvpkqBixx4jfN4aZpr2
3h5wyq56BrnhdXTr+lcHfSShmJInBZk76kKGGmfgL3e/E8SOlAG5GmZ0u+d1kU6O
6rUiSnhu//Pm7zZOlKS/lGw0OVauZI5kIVkf5N54jVHEoCTKaBO7aNXV8i405P/j
K4ZFJNFz70DNeDrqURKAKEmuy+e2pKZXJf/FfHVaXsLkOMsqDvbE1zJN4aGPcfUR
ylTRi3DJrno2vr6bQIsIgg+ZV1qFsYs13n3sqT0J6QkaMd8Al+URDnXwnAes9YZN
j04Y5QZeAkRXUlH302OMOuLqQFQPeXHkDjJReOhQc/nzCzXoUklukvfxkBUha3Ww
nnuVoYqvBIRhB0uzLTTtk0xvZ2KX74diIFPd0doXBPXrXjm9Qq5Hnb/vuro7YEuW
JdVOKqwEuniWAiDwFYCa92kqI+S+YCHF4CighnRNEy7ghHgAmamN07gKgNiEVcQ9
uNPx7IfwRg0RqZ3hX6oOqyRF3VP5tLzG5axRp92AQeLxBv1ti3cWRfx/LvDrc2AU
OgWrcGj6MvBKI+LS+O/tH3qsq7OsetZSALUXeHJwaTitkyKBsgci8r20uvvcORMD
GiOcXEDo5QiyeGq39nNhPTacOQXLoEcSQr2Y+jmSoCEAf/jfA59Qey87yAjrBUsv
IxDmqfkwLELE0W+bmrb1TwgPt2m2T3zztHdRHYenBtGpWoxPfbrq069DBDxNoh0O
TEzFvHn23t/cAD5joT/yx7ehbFnEQjWXAIEjyDbqRGOzmSrpDe/gZMKcEulntECp
xgJNAw4xU/g7AlrgcVnEZQ2Fdrcd7RJXqTk5nrJRjYjBUa2I3fYKtGfXs31tuM9s
X6V8pB9cIYXnsJxqtffPauvQY7/H7o0qBRyLIPSWJ/MsH1wepfID8DtUKICHWDMV
J6NqeTEpncpWdzxUJ/QINEloMka6eHs9WSTn4cFIWU1M3pbXe5kkpvxsWukDXGMc
5COZvphFpux7gOCmiJfkA4aFf0G0VVBCz9f3Fm8We08qyRriBHx7xPPv0Xl7+kTl
sk604Gca9TBxsSZlLKaJrZ+ubBuBYk1k5N6tilBy7i6QEV+xr3Zp9cDnJCL+uWGK
lJnlj/gm5x6JYpFthS4XHAv8Hu81RFDILXUFIsWn6LmjlxC0ZumHFmKLgPwUgwoe
5Vt9xT0GQTMmHJR66VuSon7OpumDpggIJ1g3n3QLFqfORUAfO7UtwTE89xdAs1Y2
Uyt9OAWLW2Pk1NZuF/sM7xxvMmhDc9knMqzPGEv+MCNw07TJ37Rz6YX2SuTubAn/
BppLLY2/tKdsthxY6zS5cewnl51/+JdHMCX+WiTAet95MqhWljda4FyS4MbOoocj
JjtghizvrFYvaH/yDlICXszIJd207gL35isvaQ2OPQy+U0478Sbp3Pvfo73Kk7Pn
AB8u9xlXK4keeENys3IiyZm07Wt/X7ms0vz1LBbFPyYQm5hzRLXLBTMiS4Q2fwf2
NsL16G9f5L/KS0Iwwh/DbSVBSGjq80h6JO4KPTy52Y2WyBArXmhdyLQIXjEXgdQe
Mkh4ZzF50FukQPxv5uQFZejg1Dx8JWPprLqsLyV+BpdsI5KVlqUW6KUUIpKntBod
SUaQBxR880tqwyD95nZHcWzHOSv0ylPaftNwUCjSRQi1TMI8JzMOwx8T46W1JA0z
uXoQn+RWR+lEcTMXfABST1+0hJGEKUrYxNlrKvNmV8xW4Clkogb+Fs0uw8LX8Msg
lF2OJSEDcrXXIMwdUBalpN8POtTiBMrqMlNmFSbdcrVr34cTJUoYfkAoEDEFhFVW
c8NlKV/dq12oiN5wrtWAiy0H7OqoK68Om6mGKBfgNAzqN+AmCTJQrf976jkzd5PY
Wum/1hKIAjfnJOC5s3GtFrwVEdiRarYvX2qbWDjAuqgxjd04LZFn4CZrz/msx52O
4SyCP/ktcPleZfXxa4oKBonq3VbbIniyqxq40xJFP7UoMs9uRz/MxmOlMZji9hV2
WWY/FC0IX9heiMGMFS9UegrWchw+L86XdCJ8zzddpNywsrr8OHwhcACUStpxSeUe
sFgSKD84fqxBZZsZQD/PvFzkUOk9+i0SWXtwM8LQJwrmWLICTl7LyoT7iwlfNnEV
M4V1NuiPJr4zg5W7C2w1+xnyJCLbj6A2W/bPmFIFg4tBMLTZny7DLiu/ssxcXc/t
eHeG8BE5z2YVKaQ+xzxuq2oNJzuHXazmkiJnqXln96flG0swreTjb/kvtqnD+evO
iEwkhOyrMDS79MxoqkiNiydPrwyfnRfTUsXTWlBBiGCgA5nPD1LZT8U4pre2/dmd
Kuit6vSsUUm5iLWuFH1LM/oyQ1B4XyuMf2RE9W/7noa2FbJf85gT4Eedov+5tmUH
JAiUJNYjv1mdYeJuypkPntT53P7YGfmyHh5pWa95EgwxjUWd9i9cgTPzQ77iYRjM
i5btiv7EHhRHItqZOQpue7f4je7lm53ZD3gJuVEf+IX55VvYJRg+HgjH28oT1R3r
WjrlCvH4wFxFiJo5Cf1N0dEHh6c+82F6MpGaspna6kxCnK1ChhYBmWn91Ynvs2mY
y7JUl6VACM0uDFPTNOAOHmWJwq8b0HRnnNLhlJDwb9hwoP+zots9vdMjYLr7xfT5
zrsd0Fk+bOkleCPD/2LS5srO/MYHnv12K+iW5Cg1KAqNzOe6Siw7eWbkoPBEQpN+
KQkCfCd7J3ds83z3YLOWbXQTuIxlX0abuwvjqhY0J+xDsaS3ud6FX+y0oAHPCeG/
I6MDtYjuFOMYQlUfy3jE00tWDvsntsIOodierdaxgrfayT+5RQZo77TdTyKxPjFX
h8fq/SYl6Az+NcaDdX+42hVXm5kXKLVEVu3ik0MSjAWRhSLJbUrNLcklgacUvcii
/aOoTODy3PqdaVD96A0oyhW+lh11/EDGbBbHYcPuv96J52cx+f8U/vsFLzkhrVfd
v29vtnH4iyHzwKIJKpNYrxboyycXAPtG3aMsaMv/AGstL/TcQ6O4VnSneRlsaR7V
rme5Yka48FGGjFWkTYnuVYX4GpWA34TEs/loFxzf4P5walaFjFmwbiJdvWwDQWbz
HiKGjmCjx9JaOENzMZscMPUGwn9wufSFgKL9xMpPa5lutMsL4g1GyCdkxsVGL+Vw
xLy3Uf+VPSLbvJz+uRdL47LtnZ+IaN3oo97TWZ4HsmFI4MHkB3/DhX8pZ0hoTkfM
Xg1jeLr9N4uPVbkimv0Eg7j/XZO4Xpbg7xvSINncvIBejUq63EHNaSVC/KiwuZ43
A5ENhqPB5dDa5bj9AwjQrghMFmUWhQotQc2LUDzhK8fhQUYfcYglwLUVfJFAW3Fw
Q9Mzqob/LfWRf6qwxV4HYrdV99kdKebJg1K08C5Mv2oCKtgkqtX9A9m7KNO0Rz2G
x8c0Kr1Zk0QYgZ+zQO/nyTBrVWzCQYmQODXqn6894hnbLHyoL9ruxEELUlZNGM83
bIBdbvwSZ0u8qzAF9+BO8lgAMd+Ej/W9YISwIKIMHnoS3Vozt4l9Qtw5oxRorcvN
bQOz8NRtH/+qaxR/J0sKJqB1vyt3NngJYJmvu+5pT8pCIPPyVzWELJbdbTmWqOhX
y5QXE86sKbA6y+BEogcAZzY3lx2xLu2o0H2lzoFp3UWQO2wgwjpVMsoF+ETUHqad
RanAboThqHg2TBOKBxhXXfLbY/qjBi/h5otiLtmBU0vZS+4CwJ3+1WkxF8rh9pEO
r7hQzurIaoGOcX8c0wuZCptIHNmJFekY14PODnuUEIWbuWdpEIrRRTCf2KXFICie
mlVNoQRCs/StCTVv3qqPVHnfRJd3v4WI9/L9vMc/0aVzdX0+LshcRzfMw5kzv2K3
QQ39UW6JMof75xrWrZFz9ifF795mt1ehB/GfKHCF39WNR27BBZUo3tVCDiV1YHVX
MgJkT1VBLwPz4NX3pRJ6EmTyNX4KoIQ/oSGaTNaR7POcQ6eKyx+4TleUBOZ16qMy
uhS5L3N7zZTcRLRaLON/1VjDyvEpK1jHf4F4Ja9FKYX7zO9itNM0qP2YApDA75vn
eBgJFtm0F1jsfl2K53+29jN8PiVhyprmSE7Bqm6nP3aDyLx+Rm6WoKYzci4doYLK
ubRtz/+OtfJGmdOJVUvWKTz43Xp7q1iIIxztGi71JmW4c9c+H3Ktz+Qd51SUuNl1
rJYnw/XLLPJCKJMWa14bMYrm2zaaKrrhYW/+UnMiWs5q/R1hDqTZ4jm+c+8U5IC0
bwL0D7/HgXBnT/S8VsdA14yss2jLlUsQNTaRBKCT+HFmJwenbqEkzsQw4lR7zNw9
x9oO3y0wKuCtPu1mQPk2LTjwCPC1JOrPrWtWK9VPjGPJbD2DyvjGY3JGiUAp+a83
VaWfscH2ATio9mRjdtiBliWpMT+71WSxNU5xDItM4iLXoSgHLAZiQLE+pJCYukq7
eQiuUIFGtAYNHigS0yJrBpt9ULbJNqCljzr8n8h0RomzmbsjYZ/Iv9yKj5oRXT+O
wxg9Yxc8PDBnWPnv5DuVDSw6+F4ZosiD5Rq73nxuCU5I2z/faBfZAaGNGxaSqTjC
QezZ/Ros5latgd1kXEwFZ//k10zz5W5yQQrmcbD81VX0TGIvQ/ubhF8OSfUoCrg+
SdL7M+c9vJD77Lixli+JN2i728y9rZF4MJSZe6Z+HiyrCou6YlSQOM8/WTbwuhqX
81RS/nZ8jJSemwGwo4CaaRtPFjyO+bFteRkVTtRSDS6u8ZsfFcIo82S5+KQIlt/J
OJC0ehSNOOM3EAp/wmF9O+NgnnHqg3fLcPoiea1GvQcRg/7y2SKfapgiSc/Af4BJ
UdGuzqLWiNlZYSB8EgjmqVuJHYBY6o9XwApK3DMpxwqTYeeZZH2P0KS6ui1Lwlbz
7KsIhIAPTr7LmbcaZlQaynkl3jyYQVZC8uiTXSXTQRBdg2D+SN/UUoxXaUuXaqDe
pqwVEvcew3IeNTRx4lC0vXq9JRVKEOPoekH87foyjEGbbdTPkY6ajQxdgEbAjCUE
OqlS6Lmbf0xV/ZKiKX69S8UWy4zC88E8IfdoG9XgJeGo/0v2MEBIwY+fmr69bhAZ
1erhpYoila6Nm1vSRGCCcoBsWVar29PbZ8TSNrrKTIwbVs7A4CF1N335bjNtHfLu
d1+ry0Vh1LuQWVi1ukmVcyf0eXnckM2ymbVjzVKxitLMfxXL361J69Nb/WNg/d+j
5Jy5qvwTmuj1VAssshSb7033HYqLL2CSGJB3EpaFim0ovtw21ye1qHgpc5QVUlw0
giLuGGRtyef4Gqs+p9EAh+4//l/WpN7qzP/LgWdkjwHowPzuZeE1r24sVllo3WVX
0XkpgnVzphWtJ5Taxuz4Z2FGllGK41t9bLye62aDOOoLOXyXgA3SuaqxerjkqbR+
upWxcN08DYAfb6D2Ch4EXnvhOYNwxiN8FunVwLpB/ohV1w76BZeF3WrvU1jH6DDK
K1oieqeVBDKu3CS5zdAM6b+D40WppgXruGh28XpjgbyPmCMKU18NEzNZkaKNJi+8
gml6sC12BlH6cyjj6JzwZCSTxKvNVH4vbP1cOuI4eUfbarR9Xo2sLlFBVccAEvR/
nGJA1Hy5btKoXlJg9TICrYt8T2W9+leoUcl5nL6T7XOsjRzQLbjzJIZs4XbXeVTg
r7fE3bCnR03L+xxsvr5F2dhypalrKoraBYH5qYZ6DhACXhw6g36uLEyifR/MqEnh
xufxqUQgYxJKQuZ5jSnkcQX//xaydUp80kA+whClkQhQBVtFEqvKR/WiDdOFVbwJ
7KEUmY+j45nXSKONA+XTHjjo/qaLtZvfrm7q6vPa0COHFee4DQ7+fkc/R5Abdck+
7oldxRUA0FM3iO7oL4mLH5rhA34BaM8xjHqkT58Rh1SyRtkKGR0c52SE84TydmV/
ORwnBSXQk9QwEWvKsuLZClHW5n9R2EqnAeOnUqrvRY/WfMPLRu5Pp20GQDPE0tXn
QxWpy4Q9h7j+reXRHyDwbqQg80aUgzfQOC7oQVZZeET3l8bPLpwZh5fMWkwgkady
5NSAb8palSYT90fHi7Z69BJi86PFqVz2/Y6YWmRTqpv5ngpgiwveAoxThiGTmqin
vpEsUyp90+Yz0LxGqo0Dd6r4dxwK+S118zWWqkQiinmTry22g5/pwZwDMLwfNPfq
yYuwRFoYSdchRQ0ixVlzJ+kJo5toAKDTI21ok7khGiiNq4mLbbAkjOdGCI0DEENW
UQVZmPverJQ/GMOAQY+NedpfcRBtwwzcf1yZnO7ibfmi9Tllwx848oWCy1ezu4Ra
qD33tYmoRwX/gZJAN+B3hVMZnGHh9e4+LOtkHesmhK5//4nJ5gjw/zulnOTQkgd1
/aPiE0SLR8h+/lFp5Mec2IQunLSxkV8DNfAIwC0b2SgPHZQotOPqg28NQM1scdas
sfp6kakV0vSCOF+W0hmo8kwVXzuf5H0NX4Kfmm/BxreQS7P16uvwMw7PzV+icdvE
uiJiMm9uGSO8CQQ63sikNulXtGOjN1Gd2bnDCqhgA3DVNLwmWuaaKA82diK8rlGS
pnYrLakLq7KZPINHGZ9On1uhbbIyajs1lwbW8zlSaygsoQSfFuSOVxDxBAbKYOyQ
2b4stPrtxFduR1G1lvIS0IzOuTo4f+KrpFOZsd3VdATc9hGQKb6fWU9bRvFYCMOM
ETYfW0S92q7QQvu/Vfn0GWewAuX7d2pvUWH5kE/kiUmlqVqjXnCK/Xxfcrs33VOz
9nYV2BwDE0Jj6+6c45tKXqjeMSH/KEZ771aIe6wXuqq2YISPFplhOM97+0iJ9Z3Z
3P93jiGG5Pyk5Wz4fIrh4jMHMhqNewrir665dfYhcXQSUl5dLUYhy2H75+h8OFvv
RB/EBB9F5SIqPfEK/wCfrZBwVm+fvVnhiJRtemjR3Mkk0HC7pMxuWAJty/BqqShh
4vNk1gjGLf2CdgoOqLyqLc8vkCg9uD8Pf2fB8pXCy+tRfpA2Guea932fFy9rK+K9
Dk9w5+/BND7XyR9mJ7++eXlYckszDxZDvnvJJzei5vUQojYkt/JV/dKARkNg7jtQ
nzpykEPfrKb7pZgoU4Dj8Y7qaC4AE5brszVdPIhvz6Uot/hMGzxX1oXTI75y6NAi
yUgq5TcRzDGwPc9fWl/25xm3HAcnils3PWw8Ge9QIUWrD706xBtfDpNqzAcwLdyg
VEEal7RAeD/mjfmaRQ+Zkggs9Lhv7CVqwqxkNoxNseJBpjGKnhBnEjnRvJNP0rZ5
VN7v7vZBgTsujnjrXHeubobFNkdNmD2xYIooP0SZ68g206ZOM36P2vTHYpb43jaM
mnSxJu5NaPNeKZNG+ZlED9VScwurJI4YzyECwIJ/VJDdR3mMdBDGbBb1DOv+c9Dr
aHuOSf+WEDstWItbdjJ9fZYAkPQ8fa8g46O0i4uBzMc+cOZ4uVlVWUCuyezKp9Ys
aX1/QDDJwWUq1XWQKmXu0FJspdYLL1yJ+PYHLGhKrLd89iy7AlHkvs6NXXGcTiRa
fG0S4PZMlmF97peSIz5sUJYut3rsLmSD2WpwVyotQHYE3b/XyhKHbjuSFbAZyJhc
jIKRnvNLTE3RIOkAJXBwDTP2sdZrgBR54mKKUElivsQFki94VSVMMSE2Db9OFr0F
5b9mCibtwaJSER8YYd/lNb2xGLRbte6EVm9kjYp6RGZjP54hm2uWdVdsI5f07Rlx
h6xZ3sq0IZNo9tIV79CdyRS/2xGRhwoSfxbJmM9pami7kXYt70LpJ/sK45ryXxvj
MIjcLCG0b9Bf3EjQ3u8DqOnmLFTqOum0ZKVRmbD4PBdzLGgjxkyZvJPYjfeD3ywS
p/WpJbqOCrL0y3AFsoLwaJs9YORso9THpOVE3HsEN9e1wPj/ojCvj7qABw+Taqio
sXzrUZKFU8GtjpUxrZ9F17ucRF1WjW4dLYkrLSG+wXOv5KygGyehp+nA+YoLkJu+
dCof2leoXXwxAvHyKSlnwKNdu2Te+hmjTy/VwhdxDzLzXXxeBLLRlHNnIxRxflb3
QgrHLwHDsyOCsyd8jYr9Gn2xpJ85dK1QXRydK4Wph/K2FJNGVW4QoPJ1gX+KE71N
le6h6QNKUoGSSKMAhD2TZMwqxpbl5o/Dpsu+9PTZMiAVHiomhbsIvVooCNu4wKrP
7mS7hpdGvUcy+ThwExprYW7GvhNEn8r3T+gk0HM2wL9QEgXiRoutFjPPX9c30k/5
KEhXDGAbGg3YD2shpmeACHy4pc/sGOAfD6HdiyJ6kAteCEOkaF4C2iMLHsI7a/Qh
QcruTQwnYATrfUiJJWEFETli/h0qCfj901oGfWNWFwHKM3bTzdE2wxPHXsCys9te
dgvJg5DQc5W39gvDanLG/aP0GrZ0WFidbXX+cLCTSBFwCj2ggwFqCSwCqbyuQXmp
KPEhRFt9s0BPWbSydEk4tpJVhKovzsYi75hXfUnbr59DNEidl5Ex3SIKIqnXPjb1
eo4HlqIJ5g4IWmm+0k9EymjyOJ9ijZAZRF/h6MtuQ4IE66kKOlq13NlKXAi4nwtD
FG3bo36/DJe5j6WVg3SL96XA3JrBXQqPHH9Qvzo4uOxAUES/NWQaCjshfQO7ylxS
LwkisShJ7tbwJNGjyL9RmZVspyhxlH34lD9VJrOLtqLevjI/eoxyIBrkRecM3+Rk
OTVwpc7R7NranAjXS9thQmDX1Yl0AC2kA39LrmyUZstKtg/zFPCeCZlWxgsE/VJx
vs2RnELQ8iMNiHiheqRGDI5dCHUtvEuY/oMj4S02TnSoaRajCYi1Jd/mfNVgQXSS
QHmT0Z2O/qivwmvw3kO+IXx8C0BRqbo9tC/eeebo/CeWWAi9t1XlGJY3lSTmLPip
aPVBzraDeVe8FaRG5nz3iQa5vbGQqHx0k14CrDtt3sTkZSEVXZEqnjqnbXApHi3A
qQeelYR6qsLDwH1vljEJdW9+XFPsG1FWrHwF0K/1MFhqdApqNV3o4MxztIt2rsPE
L1XRcIIkcgJlajUI2O2cnEmkbTJJVF+zeDDSctXAubYu9WGXlXccyGyD2hCIYBoD
Njjl/ADFZP7lg6us9QBmTTTBA2uAC+sNpku43vvajQ37YjGCMdt3V5ZAV1Qm6mY9
TWqkXYvVyyuiqy6isd6/LOfyftjg3vUCUV1f8yVukbmG8rl+lvUjFSPoTq3BpKUe
3Yiv1T26VWEtRESnCRGlJHLkfQMp3bI533RWanwJqeD9mgX44tFrhsmXLKeKto3D
gBxgTmbEbxQKp4yR6ZDDsM4xiLSnJTF0JzlifNg9tY5iEZVIBnTgOwr1m1en2e+m
i/hWGq0FmX9S2Na4tCDLu+JW1w9+WWIUYAiQV97zNWz7MTxZKfCBxafWxDvt6/Xc
apwGHgKpNA+nN+Kta5c7Lja9xwobAFj3WjImjDSOdZyeiYO6GHMIOCh7OxNcfKBH
1UWaRMCTm/2m2uGHEMGHN0dhyce+aS4w9Waq9xwjNUMlV1moMF73BdF1pTG+d/K8
jcbEK4psBu+rG/ZlbAqgwMtUS3coXpkfMgIJQuqfB9bxh1ii36frPexN91gJVKKA
VF1sokqrkFOjF29iG1rtFptBQaCkQOGWzjbaXsEnyxmAKMpCl6bXePmQsmD6IjQf
uWAepTCulUcZ9sWY77/25ojNHjeZkcNweziLqRpmF5aDYdS9C6xNwZk3+kcIoVH9
be8asXu2nzVD9rwGePt6mjI/gmBPp2rB6/My07Mfge91e/xOZnycf4JFPeBxzvNO
52O3yy+zCdmDPcmPFKYw7KmrJgFrHVdnWXA8DzzTPR8MtT0LymRFsWRru5a6goup
0E8kjwZYUN2YOBwqqMfrOtwu1/VxxAWySCBLDNfxJ6ZNMCvx58xhKm7eQpy5nblJ
2QDjcN8Jfu0P/YBXF2Jz19YcjO/OyA7nC6INkDykqOHK/IlU4mjXAg51B/q3+902
iepI4Srj77Wq30hCdKHUKy6QkiqCl2Dos8L0ozHgYOlQeQe09Ymk9imsxnh64l5u
bPYnHMH+oXQjks9bxK/yqstUALYhGOtxOuUtDCTyK0o6NZrI+pB9rzHMkRFW5Cwb
zmyxitLJHVKdkl+RE2vg+JZ48pmkKBDLZCg75DLIO+AliM7lZ4bPjxXSteCR/wFn
OV44872lOZ9lO5UofdDs+TS4laj42DCgWrnh8Nb+EP6EW8BfS4dhrIEY9FSdvzjW
vivhyt6gNOg2T1J4tXgXpTuU52LlrlNW3GQ1X+IlmI9+fAE5yIAgSDcIPNDwTvVf
v0RvNCjEGrF9RgsJnUm0/KIk4agilXEKV0rQXs+7HscSw6MMsTBoaIPqT+n7itLj
bjwmxCF134N3zZ7VIpmBJEgu6H57ngc2NbKRuGz8uoMgs/JnZ3xnokQ7bK1DiekS
BxrTC4sxWv3cJD49WrpLZOsa5dDUYswdzb/QehdGjQbtTasY7yYFrXq0cVHuopur
/eUdnXvfBlMRhWO6EagNsH+og8SgTMkdUMQi34JKrnNXYHxOnCzTJdPah31UZ0u7
JmivOoRkKOzBVYvjlTkat4o1+yfM8jawd6JIq9m6FQbSrfNpMQzundnneJRBkw5U
JkcaeWVrMnK5FPNhnZVCTX810o2OL5DXLqoBsA7AoRVpabLvPQwmPO9+sXzKuEDr
7SsY0/E5uGIRUbqURtrA0CyKte5DwQGOuRgr5ew3jQv7P8miaW5rx55ZeRcnhFUe
BqldqGlZOQBL5t2UaMcENldp5pgcElHryy/bFf7N/B6HcIsyL4w9jgBu6BEvY9U+
NO3PNEOvgdSHUMbhlRqb8Bfp1NewOj7ypMOvZBgZtTSraKJTbwF/mzK6vGBTKGXp
69Zn28teewtLzsxveV/ItrY250BjYGgqS7IYDaVVvjND8FS2t/+RYG9KVeyw893E
wHhm93jcmPefwmrfPIXfREl/7AZw2XdKZL4QoGQRmOnZ7Q5wPG/4SkLFG78W5kIn
8aNC6vHTfu8oTx0nVN+//IFXy3+I9aI1mKrAaRU3SNOVsuVEUWWwkQn4xJnitfGe
xKfj6UyO2d/MnSr8MrfU/lUUGjF20XjuZUogb+NAP1U79f2FrFwXfostIRVG9bw7
JquPHt/0+/J7bROVIvmwzJeAuGG+sErW2IOFHAIE/uzTOJ0Uu4H8MEKFBxgGEixq
yg2Ghfr8f8ImZ7N6lnd3aVgq7ziNKFSIEbKTskxl3ZcjVDq8FbO++k9Hdk9I73E2
TReGpGikofHXj34odzMNYCVXVnV6fmQ+DZcwc6g4RD4DZnnJAn1o6tX0VUD1iXzO
Aih1KQ/Vi4xdXP4P8/nujaWJ0eFvNkWFGwzAucDVoETqcmU2UhB7JyqEaaR/dFvs
NfKFVZ4/21U3N5jxkrCIXx9LB+WDJZ5FQPkOuW6AJQbxO0+oCGfMDB/IKkMZZM2Y
5+YXKxx5fOkdlfMH/H+5CDjlWugSrvo0UAVn6uc2352Mvkwz0LSvifmF4vA9y3Za
iHMopVBuKrVeePKmeu7tuc/8EH1ajzrhiWD1PV4SvYRb2F89kYU0IR40N4lmszvp
dRZbDKDJG5iZMa5kOvWJrYtf0PZJGbIowHQcFy0hF2JZTcdjKTBlri5WsWbPuz6u
tFQD2ttSKcuWzTo2SA6kp7+qZT/D1BtJC9iSz0m8UVD2dsilBlQUwbbrr4nlIQL5
2UaW3gBtPV4PFibBtV6ng4GxsxDUlEwFiZGjKvCmQvTXY6pUcPeStcO80UU8KaHX
T7IcGi0O5nmheWDetnHuRVBzr6Mx9FDiKAKleK4J0uGndZ6PRBvmxGqwsHz0TLsM
ej4+dOJzg0h2pQJ6D9jLry89i3Ut+U1/Lmeyx0Kg0AF9nRsXHUI66SNivJxKAb5A
guPkgY79WTPYbc42vCni2WKfV5JlTxaeUaadlTqHpPv8cJkEx7VKDVoYNHsSRtu5
aNqEGJVIYhcCTUqiQ4gMLSmv0O8orXD2qcEWd9BBZCKEGTMYY3jF0LR2drYZu/4d
jcNmsSJXBDsnjFEe8g63SlwWzFZrw1bokgNLQimi4ev163sMGI+tWr+WD2RAAei8
Eqg6LJ44MOVGTLO0SVAY40PcArSVgpHVGOHxBBnEiY6WKhY0hULopMnypfjcUjx3
f5KhzBxsorIWtn2YiYBlSApV8OegMMKznI3MN7hKHIMtxGdT1wn8qmsgSnwM+gB/
P7Sp5yhnIYKdei+ZERy5eIzy535CJhvCxkdswIYnV7JjWxWOGmGu+bSC37hiJjXa
6MmBGQzslrks1j9VeHzso1wFYv0v1UGGwNI1/35rAAuxQghZaja5tjA4lbpOsB7k
5Dj1uC7p7Mp3fGKKkxRjgoMMoagrGhGw/65WecpAtqDwqr8F3z7TqqP5HqYFbcLH
37dL4wmIiKmousxPzCejQc7Mkscr6Ceyzbd4/DzCttGa86qkvVBfe5PoCu53vWMw
17lWGHI2xLoq+OC/c9I8E5qKaNPlTUwwkOF1EEvj2PNiwkdnJsPXmeg7liQp+e1K
U+P0imajCTC8sIDFA55d4IZUiD3pYineKfv7ZH57606C8SrlsbUEKKBLg/WNxP8A
iYdV24cN3tPCeGenqCRMOom0SIgSyiN5xqGJaI0vnbCmty63s9WAv6m0fcGmxmN6
Qc+TabzRv9j3P+Go75HEDEqolw7a5+2TW4K9RO83RcAkvYZAma6ye3Tznp2sdS4h
Jq4HcLSFNS+gkiZ0C8/Qo2VK7qyL+XWOTm4B0fk5UP7WV58S4KJvmJQt4Oru3qNk
Rxr/T8JF7+c3Dae8gnqnHg/w76BCEt28mjwEFXVLelDnYm4zvrl57Gkq1fOwaI3a
8LT3UL6vBd/cuU7elXMP2gSRg2tq+H4dxnqC8htIEhcifvGTs8fu0C8RCt+M/HDx
VU1SRNnbTfeWh+IxIRrM1Za266x+O7XTbtT/0I9VbulVKNUmYXQRj/8Fy66lhytB
9b6YbVshCns/3WdmpmtcFwg5Ab9vz4yKZ0FLwUSfXPt9cIGs+NU7BkE079GfbzPF
qpilk/dKAk/R72tKyOf8s/h5hjI1vCk6R3bu27Kvi0nz2Jj2S9DZVAbMvaxgy044
UFbLgtawsIeaNmtVuG6WmY4NC9pY0Fnk0HzVIgMd4kE4OyMhfOu5kl6Bpuf08gvS
lRxjEtg78PQQeSwCAbzTgZ6cvN9FFqxIRJVD8Tg9mbJBYNC9YQNCQ8H2JijV4V2T
HHRFX1JikSwHn9PyOCS0TWwbmgdfRp+5GgmNT9xtiQbU7w1QJhML/NOWDMfdTmmH
nadmA0qCT589SZL6HfenrpKfnYTKRw5rXMQCOfoypb34NlM3sO89IvKCGKAwRKt7
dbnXnpuv5PcPEm8QKKgOjXavVlgLCE+xPBgL/15xZpzmrJh9vQteS/ygVojaUYz5
JtGbu9ABhybpRkzwNbktG/UjolwoP7ifhc7oO8pIs5I2L8oLJ8slefoZe+fzwtq3
meR1iqmnovanhFW8NbdMxu9Z80usri3l2dYRf7sMW7GfYxTJqNsTc70OUJt0OPS5
j7Sv5h3RfntDHUysvOVlBlI6sLfIJmkiOhBr0Q1pSOqXSYoP/6Yh0q830AJaDJM/
wkUKoKjOs9LO/2acpb5XqcaPXPAcZSGwBjmR2r6LaeAFzI2vks/qoSnDvqMm0Z/r
Ie749QI2Pxcj0wx8jKlusds8lFmbJFm5G43EDLs7jAg7FRDwCaYJqJ0QLtPly2rO
9Lf3oVho9hlmdd+HkF9ANbfvHKe7eKKdxGZsYd1iU2/BuRHL0xq/kDvfO2XwBD+F
5ao8Nay5zUxRbxNF4lUxmoq5dGHafUhz+dfxTZ8+2sVJDhL5yFwNNW6HInC1+t4P
xWO730twFyI1lKeNVdJ8hKwQypy6MLnK0fLyrpmNxm1fb32JdZXdgImvFiJ7JtaA
B1CnAqrP+GTCKaUwbFqJ8rEf5wTA6UNc8p8PJnn2xPgcNIEEgJqCA+mzWIUXjHct
xVyirdH8Hqis5QH+eNNUw8pSB2ivbL+ac033X20HCgwJI6v1uR+97xyn8+ydXRs7
HyqmHWmZltbEYFvXZYMRQg6Pu7wnSP1dv9bbQjnRR+5+Pg1AZA/dAQAmdIL7g7rz
aSzdDW5RZPQno57NTCgZ4YbSls8KPA0mer+3uGdIDLk1E1Ugz2oPlXFTEzg4GpkJ
YEG/cveVekILJ7t4JofLfZ9fv1RoENrA+qHrkk11C+A=
`pragma protect end_protected
