// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MWiRNdCvCmhANFFcpG66N/yYRH1/64Rn1Gk69ZWxlG/6o0eI16q6rUDH48l3pwBY
SJPU5laIuFkZNtJ/Ypd0nHc8cmhrDLB1hiUdDm+uxd9p8xZ44yXhL86NLLahunbq
fU0dmCleiiGG9LsrtmJqZmt8x5xFVkTvkS8Wt2DekWQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19264)
1PuTxpL2fUboCz74ht0gC837tU7a13L52jBn/GdSUFoUXK4Suakjbm23edYjupYp
BRz9Zc2yyGB3Ij9fMz35irqVAYI0oyMc/f1K6X1eOru4YYLGDkSnkLwVL1gZDRfJ
WPZadNH+L6VQe6XEc6bHSbTo2DdR/cXWmGmS+GynYcZvorFQ2PuA5muk2uD9yOF1
8gF2pxlPP1e4WAC6HocjrMCLW1KmQV0vJe5Q+iZ6bQ6g6MZkHYHr4jocJdE92o2r
Zn1iLvVkw+0UrA+5cT2mNJCTUT+yhTSwLKsm+EvxzA2XAVfPwnajRyduyTUPKRSc
qsc8vatM40HioJtnUSusaalROADXmdYruYEkny0h6H7wSKIirKQNeYjMLGoAVTBn
+Nv7Tsy0NeaRXRafTuiw46Br8Gon0PiyNVslq0YVxU11fJKGdIkNKUYHwFhNKYLX
sHujBQG4tWcX1ojuvnV4JuFCiSXjzAOdRWmmApFwhkNfn7spWmukEaLUion/A9mn
c2k3/qpBbxjLjERJyenBQSJDEKYG+Xv7wfKHIrvwZLpc3Ts2Q+FwXn+0Jzg+h9D+
i5XvJVlWM6YQLz/sgWFJEJqODp8dbSWgipOLSsLaYdXOEY1Khi3w/v2E7TcQrnPP
COWvKtFWlvO8P+URqX0rQZKeBPoG0NtyvTOuWbArmCZTASQIcxCyWfx1JlOab5Au
5hQgP8gryZJnqpoatAzQofrxfv3ItDJD4sRhNMuuFkit33fFBvaq87ZF5cJ/1tsJ
WY6CsM2avyZTRIlZEGAZI93jeR2HDFeGLJIi9c+4oniZQV/CSrG9jAE5DDMfbSoV
man5zWpyz9ehuVd55pCRWtzHfdTKJjNwjWWqzgJtgcXHrycEEWiZh8kbsE8OPYYB
vYh+sqMiQiQWcNqDYQcljgR5Id6nfLYsiU4YHRSHlCbsl7Dd/lpK7kjGmn5xZr1g
dBJbTSNglkWnTKftnWsbFKeqaI3pfjFylmItXgHDOX1QTrxvxwGlOjAyDVC3Dv3K
KX0jDTnhhbto1FOOoTE9jjUEmU3nm30uGH3BI4/C+/TCFgayqY9CJiT/hbeDJe/o
EIlE/Ajipq7Qz6Kqs+dN/QVnLy+9spVfGTXowoAhjvRcdrGgP8A8vbPrR78nySZn
2UGb69uC7qYq41aUuhTqOaoLEjK+MWb9HiY+GqWjFMOcKkl4l4IuLhlGtmGJuzQR
2SL1DKhNHuMzdA2jgFJam5/j5P03IvIJD+swtyD5IHzPOkhPNde8RS2uXLESO2z1
mgLeu+VUXWZZFfKwAiLZEWx/mMe4biR1lYsiWb9Gji7ceGoBQiVJ63BOC3GdoSHH
5rfXJEJkn2swzZHcW+ax93bV4KQisHhJoS8R7KWH0lHIlouDKT9rPjV85XyHXfnU
PpRRZFQeibhXkKrtMpw2dlqmHkYtnHZARoy2iZebICSLxZMq5hilWMT8RDic3l0P
FOQivu3sXEX3/HbK19L9Oj5PctWDzO6K7MCIYhd0UQ7LIe3i68tBYfsB1/hLK9Q/
+JqIzwK0+v6KBQiVGqmNm+6HTPt+VVP/WVLqjeJVRug/TtlF9UMNbO+wib7yl290
eMHbJrjNug2XYpZbdgzOX1Ma9K9Td9+Y9khHOa34B7epit3iLBPTbwVkLTXrpP6t
bAbRQggEV7FnW8+8EU74Z8OlatPK03ALHkTfv1maSM+pX9ESFwfcbRp/1o+GrOGm
j11LLMgQ6ZxDKsJGrijpjG92Pv+9A/poNX+ZexJsct/vIrOTy9wDRBFf5jgWw33o
FX47Uw1X0pJz3dcPNYtlQiTXXt1Cq08Tx61LpbOIf8oxoWqTD8mSt//HetWC4EyL
ULCSWdZok48U1w5SbFpnKHp3tTDC9mrBz8G0CVQpeI1g3MNrm2kkouxTRsLrm3t7
3zxOmQCsV9ZrysmYBslAusnzdM7jRZKHay97YOiLdR8pEjDtjUPJXt5FhcTlH6ma
nHVCGr6ckdsGDs4KCpZOsbnVXkJ8NOqzkiyuqr98GUyKvHou8OIHVnvT3tfUvR9S
Ec4a7lAUgaEHawEJfjrZCKozPX1BqPFr96BKA1yDaoKBZoCFkvmG4uXC5/jEYdwo
OVrRYowjF2RFqI0PoJhFnDJuGgNxsI+twhmJIOHB+LktgVoM+emQ6WxhZ5jcit2t
/eOHJbtItbAPEBkHJNBpRSqrqNKPm8TinjrdOpapYkg7wIGBGBwUREmMubTAW3Po
DngQshd8eOIyupP32ikRUfooFa+lIBVpOTAb7hC7MR50q/M5yiXkKzQSKfax7kYl
IhKZFmZU4sU70SIkF2Ytv2c9ZYqmmbRFOu1LkblnMmedAl0BuFoxndriQTeL9wv9
VzD6gAE779e8v6++leMArI4m9u2zD6h9hDf+dlZ3ipDg9q9/WbNTmeou/1NSrFFt
tb2+xS4oWjn1su2pkoXWWxo6plD7U9K3sKmBSx8rqJ/E1TGgKwQy1I3S3en7gYou
duwN7aFfE7gSOT1cySyuvXtevBiow8KfatCSFK2P0eELyIjJAyiObVdqrJTgnMPT
Oie0qk2WlmIbOv5F3Fm2mXeaxMJHE5MLSFMHSHrsM04iGio0uepgkh8NMabtKMMO
OuBMSuRtKh01AzeAGP/YP9o9kM+PepMbTy6lM4jx1E/Km0VMq3uwspkcdt2DY7Cu
MFo+tKi4z/aW5jauc9PaRblr6ftHYlyhauoU9NpMXrXY8NaZuhS2j92r//MgGXH8
mh3VbWDZlWgLRdBPlmDk/ibiDjpScKy3ChAOlwx/3vD66wk5hpT/FI51cBEKTLJm
TUrUeCCuTaQtyZhAAq+0Aw6sn6cm9O/Kf9eb519qgpf59tUN2Mnlvp+lVYm8OV2u
Wsb0UZXPHSk+JTxCQnyj5+EjKiHKdezxk42KjibIev/eF+syrA4wCOsK9IfKAsoW
YdOujOL0dr6tkkVwx6X4UL1D3K18v2U55Plp1WXKI1i+MAPGkWjv9wx9xxx35y/R
u+vGK9dr1vofKOcHNd9TUSEBWL6Pa7LCF6KsHaT89Jzf1BvVuJlzNWu3k47KDPE4
6HJvMlrb7bpvW//NMAAwmCQh5pHZk44B72mlITnA2rT+0FKzbxBpkbSNBeRgcbB5
wdSC4W5tM0duuGELvnTgCi4nHc3iL652MxpxE62KI2diyEePb+a/E1eBDVpSYisI
NeLHoPc6lq9ZY/PitnWxHqmbJOEyvOr1+eZn5zMheQKtqoQyTS9ktuyYdTn3Nlpk
Bh17dhyO0KfuDG6O4q215+HAvr0A1kY4hDZcUhP4NUHtuvBqXhFKVDcfzLCtgc8z
t8bL2M2on3sHUEP/JhxOduh2lp2uzQSZm25vsZRNetorSxuFVaVv0CXGlaF7A0mC
sGig6MaXSiFcbK9r8qof5bEaI4WNswxKiqS3O3I/iOpgeVbZ6CLMW2Jt7v2q0qE9
oJO+DwiPzAfiAxpniMNMHwquoBaH8vesf5ygYc8OXfmtnmZOVy2rVscbBuSYZ8ro
ES6tJvJmG0DXIQPTL2ANWsAfx5/X/D14TVuKRi+lylmBSD7Fs9yXd5rwxLWgelvI
+fMhQG/maMWclsnKBoB3Kg/G6KhukGFXvCbkYbMtGwc473JcGsrpcHQ52YrS/665
LGE7p/EQqEJ1xQY3a/sKvdFwFaBO+5nPFpgGmZQBw8I78pDuiPkDG4H5lDDQJGqj
9w+8JGSMO1qsmkWdBmAwvfTe2el9JSvhhIX6iSnQWLv5r/krHvtwGetCmI+MKo2w
vX3/b6VtS2JJqox+kYri5jB8KAyaNvKSWev69SKMSH0QSCDbgn3SNoPF0081JHTT
kLZ9aVBWgWEt8LbS36xxb+rn/3eoV0/cSXp/w2UB8XVPt35HkRpyZJs5RwXfWjpy
8+avX9WQmpdY8PKKo8T5BMJL/uc+/NhXPiLIOr89H7TuqEVZxQfEwamqD6AnZr8+
pD6iPuGrb2eMafvIIgCvK+p5Af31wdrvU+s4vPz08r21GZq3IsI5JPkcPOLqU8JC
1TneH0kJsuyi9XcrNN58HdvQOG0euDauRhGW5gb0J9k9j1GBiqNnfy8cSoG7ryQu
APontIk1u9lUJ/7XCdw4s8jEKymEuSFyn4DVkNiF5Mu+3VZJkfyBTo0GrWyRJyne
60F+1VEDcVuPvNVJsC5cIzjPaBT807kIEY8y5Wn+8axXxWCm8/VPvgMv/cIns7HE
1HIYTQ2evG2ozQcnciwXJVUsrFIZVSMAdfi5d6KMkl/pXudrCvb9V0n9PxkchHSi
NlCyWLi1rKTVxUvJjtevWumQL+tSwDJovrSLqWYEcdaVflvN1iVkJhHnotpiR2Zx
tfY9mjexgXsijTisygh+AAH52GadgSLEWSUmDJ7y3/82MjKRzC482I9WBq7O2XfD
YkhgqM9iL+AwWw0PJEnOWDSyLP/MEyv9ZmHZUMZTPVF1MQkRhSoxuR52MMhSwaZZ
ywvG/la0kGw/7B78YucZ1Kp38176x9jn1XTMNbYwEduLWrJ6hHp1gZFLjlailWWs
+OsI8ZnZQ9NzPjtTxIBzh/neIZrK/nvCCofUomyGAxQiU6dzE4vPP84C9awUfKit
Fw1c9xZIW168Dz24ZMrtVcVObmBngY14VOimp1qt4Sy9d8LUtlslN2kfP/TmD3Cc
IJPhslztig0YVVyimabgA6SD8g3QlyYG1WBH/8iqZNl8BegRnaMhFfwl+Bcztq8A
49cEFmipRyRbDX2tzINZB7g71KwZQDOjSmo5HWxe9EvDlG67g2NuH08ogxQUyLT7
Wi9MYUIiIo0MZUhp+4g0SHomEpffAmi+thDOH1Rn3BOJ4rP8EUaLrV63UvyhpECC
Vm7eDM+spYBNmGJ6WCbv5Z5t0+xijO1JBOvnj62YYvJ1ZMzQdLkI43dMZXGrmQUA
xvbZbZxWx66KPbYDmSHT+8v8kpxTeJM2AY68wVxpJRrRhXh1emF8dXUm3++ECyF5
PeGRjlWuGU15c+1SjhvFfOwHMLZBW7ymsuMSx6YHAAuToy5ZYoY+qDIhOPE6fWB+
QbjZZpBIoWD8bFAycl45hq6rXNso2q8mfqWDL8TTYrVUNDcTeJlYidSmMaX+cd5h
K0715yt+DFqcpBcPeBn4OfU+YwRbVEC/Vj1eraPGhGDRNi99/xVkJMjHmBK8eTJJ
+6WDmRcuc+nNNcYcev0i2+VxJBL+lcKVs7emg/xE76hlrDctn14GakaBxTie81a3
TNXHJTxHFq9yr+3HvLyfGq0u3KePyK5aAPzVppZcoJKUW2vgIoxBGt+oBgZLQhiT
Xxw8jbFkqO8aFSrYb7VWXM9CsnhotBvYRf1Y663a6dMtxHK7Eeg8ucrUmHrFToBT
2k19ZmT73PVEYYtpfEINHuNadDpAI2EPoUw2T/IDc/7Cbm8PuwCZoV+oeYH6Hejq
fK7b/OSMGk4mmjW0H27Jpv3txhqVTmjEu8wxCFCzH5wTmXD1MEf9Ey2Gml8nL4mN
ixW0v0TABMU7p0FvhWslWDdcQR9FlQXccugcaINIMNt9MNvW5mOL1rOXX0FLFvBA
cDLJbS+F1Pem4mlqRGgI5pK3/1Ve98u7NBtw74XefARcUBF5qRVBIYmdyYg5xP9M
NsfWUYtKcr8TupzbJOxLzwa903m2qsbIbXZPWo1bZ/RF6gKDz0+U8LNtvTUoeHND
frH8aYyTg8KP++j7XUK/XeqbLhGu1cTDT+Po4AwHtTetMxfdCgI82sspEFYgirGU
PRgyzvhRSK+W9BNmw2qoGfDEASjVMJBE/2gXoOXx9/41KjeAagjkatIdLwCmE+QD
X6+mbne1WJyVS9thZ9Wrcwz7g4XMF9uaKwoXea8tO6xOMIpdqauFgRhYFLNS/exD
5+CWSLDIso5xd5m+wYrWLoLby9pSWhzsWWR4R4G2EEqsUrrm+h4WmyEu8dfxtBn8
01Akn/AK6Oqh6lwcVGW9RIzLSai4zQoJSFXlFZYR05p0SBmYDjSxeCOWaMrB7KQF
og67so8Mmwk5icY9WDKMqIpk6sdX0/Kq5cw3TxRvoAE3vw768os7ygxjKNGbEepl
XBrQ4C10iGMZiJrBDn8mnAMXkUDa79SILUu+xJzaoH2gWhq4VFPBPZR9W4hE5+ba
GAC6hLJQz56FhcbEfUdrZ3vKTojVZE9dWo0pCwxKlaSA/u6Mj1vGpIdd4Otgm/cr
8I2KUyXf5KWY2P7HbwpmadcQ+lu/30/8H5vxBZPAG81fit8McaJeUlMwMAahEpZc
HuynAXwH2MJV561DwsoYZN2u8Cg+7o7nuyrx7ox+nV5PwuC8RgXYKDYlyN5HDNKE
fen4YEmGZeztJux0wtAOWP8ORxNGduHjXO9vfWvhnjUmSeNLf2PCQSc8Na0Fl3Ai
PC2eduCJYVkV2/e7byxwTjhD9GyqNYNA7k7ZUKE1P1rcSdcRzojQA98aDDyC6uxw
OBgcQmVEKNEk+LgKmUa2shXK5w77lJZ4mrXoSq+rFahzOG6Njpu8f6KkU0fn0ltT
86OQNoeNTZe+eO16zDZpg/Rn9mEyh8pGLO3cHQ1Pn0v9Jr1Gmy+nksfy7oSj8CLr
494KvvqXpaNznXTXGoU4o+gfcpnEXRl67PxwlzMLPVsdesDAwGlLToxwnQUDalEw
8f/sXEaN0u0ie5i0bEkZApc/6AlTJMHRQQLHanBH07LkTzfOHvObOhTNhcBjk7wZ
zlKOoALPF99f7F90XRXqj97H3YwOxuMmhcv+YZa7gFNriIZM/2f8U2qIo4U8EePe
y0cZZqcpPFGCyahrUwM4TcaK7VpzsaYYjQmL4MsrUJ4o1zzQ16uxoi4u6oVZuw3p
JFh3OllfpgYShY3wZbaB+sR/PXabsnQc5lzc0I89vbx6o/qREbwg0wMplEhzOjhp
X+3CQ8CbmTPOXrwLlm/R/tGnsB1qlzSKXvPQV5YpB9Xs7Jn21PWjHqOBSl9OFYkb
HpqmuLO7M0CSmfZXTj5AemK7s4dCtY59W5DyQBdc5wFEMGhQSsw+teKHZpK60m7H
u1Uy03+qSDR9RaH+1t6R7nxemH52aXzCr/98RSUQcw41jmT5KEynwkoYAHHZmvmQ
apIHNSbuo8w7nRKhpCf1e8fXe5Xtv6T4TSugawgqMSWNOPfVjzcCaHvtRFQ3q5tz
X9yDhlCfkoxfMkFn5u/3oio3GdKWPJfvXyMDqO/BKbI0avT2L5/0epgd0WEMqRt/
I1ujTgS+lWzFj3lcd7KqgQZQ2fwZQ+lFcuwbcDlPSjERg7JxhVZGWR4gLT3g2NEg
GUA6jmOsWw0KnN7vCgP1QjDayfxCzQaDVuVNd8DgDINsqGELwCRM1auX4EoJVatj
DaGPlb/hEGVhlRkzI35a4UzTM2m+ObGkMxQpYI0KlfsJkzNRutc89gP692pea+Ls
lsLpESPg3r4s4jhFMz857El2UoQzonA6z4kisuDYSLiZDFoOZb5ZvhNhQYT5eHvD
EmLsHefOX61/EWUd1K9twzRxRqX1IiR0A6opWUpUbKRbfAWmnmJlxcyh3wJ7cSka
sQYJVQlGRgsKecywcJIM7Hf2QBQYp4A+1KJ9PF6pt70u1V2YwUCtBwbECYuI2iJc
zKg/vzpAJ8ebKFs/g9229J7qed3VHcPI3RxzYu1Cw27tbTZzWUUEK5YSeNsLEOPY
v29j9w48gmzanS0xsEf5KxlFvezEl6TwxaoIs+F4SPY1wMOabqE7rrkeKNqpJQXQ
KsfuwZPKSYj9Y5catearQgF/NjBct6/23NC8DRhZVaoF6yMU5a5fZAxbp9CDpZ6K
rGqwGqYfs2jwCOBPeilPVjRQa9AxUukHP/nk7oSTfJ++P00BKwfMora/x3vrJqT6
mw+pIhsuTpKP9Ef8JHeTlLZys2p9edX3cHNwCddIkT4seNEqCu06QqURhv4BKKvO
7RE+tNnNH2s6dc9RD++uCWYB2TJwq5gyc2GTvktUZd6muVlezettDs7ZcfwLTPcM
cePHukrFJtoCkG8pBAjcw9f+h+AIHzJltXvOzSN91rCD6ZIvbDoY4eiuiJUrxX7v
vmJusZ0AQfN0jMvJcOCLxmeeRO4HXv6ps7xNsz/YmBEpQA3beULUqFVhpwHhHwZ0
d4HpAgcMeXxFVfnw47rOgqknrk14Vq/LXpoHM0A5BbYVwdknhnFpkKerHKDZE3E8
3LS1to51FA27kzgXK8ooIaWqoC7m31iL/XGL+BONHASFXZDWLwSYNsNPdUNTWnWZ
euJDI7Cl+7QEYVehqCYkUOXOdf7dMrKnroWKube2GmnZiRJ3ZM6z6D76PqPtj5Ne
H2Mi2DnxEt0+96MS6gqtw0EQn5BX2gPv2wuWJTHMaXMlvYTVJ/LoHWtPv7pho2sh
nQaO+xQOdaW/Hb6kLfUegRnDrupM50oNDHW4X8acxCgrsiziknwgjZ7ZVHDfNpmu
/3SKM5jlRQs+Cvdp0NImfr7k8AgA6ZR4a8PXv8eIyWdQThk6nFSKcZDe5OJB1nea
Hp7w0q45bs/XyI8g7yNZTQ8uEUixlHLQ9lTm1GwrPg6A2zDUeP4r0pElYip2PTAr
Ou67cRt8g5p/m54XiyWNMDKRq2NhOoE5yeghxWhCFhnoBrvSf5lQxTEcYWmfMBpF
K9t+mwtmi6DcUuoFTycIoR2Ue3R9CGZ3YQBk2T4Q3UDC8g4jV/O24dXMXvDbOBWN
hnzRvMuGD/O/vbeLvoJJ3vDScs2Adh2JMynCLpunJWdwu1NIf1Bmpga7AtH9A/re
RIjXIeqdeHaAPPUaN4Jrq/xJGhQjDh58PlXMbXLd04KQrHGQ/5wzYM1hHS6ulm0v
Cn7wDQn7+jZsrLwEhNhYhDWS4yfWVSbRulFf+k06NB+rumDcqJ8nA8a3Clq1BMxq
LWnITcxJsIYvjeZSpB6Pb0NsiTn+36XzS+wmladPzEK3xWXiqKX67YFQjXDaCfto
/68y7AvrH0LX0JaLOnYUKdjellR0DHEaa8WFv3K0nmki2O2eVPcRA6QUqMqfITTN
oSiHj8pAxNHKwRi4ulPEO1AnSPNBolRt91HvfJnP8N0EpPjmQuE4H1YzFzld5dUi
t08X5GtoOqTa5aIx5aIS1DNIKIWeDHUi1KzpBasOCEwH180paEpB0kXJjFLh4K+Y
7K20eG9BJ92drIY+KfEAvZj+Kf+5r07w1qTv41jgcgOoVTtdlRM/oOgt79+2ceSK
ZjAlMF0F11YWqQRiiu8ao28+VJnxuXxMr6nFgVLpWbEOywFtdvKxjGwzEjKLm24X
o1YkKejkRQHN/bBw+KxFIvJ5u3OZH/lbs0VWNeZXnSxLOG82uj1I5P8rALTLIy65
52+m7XpRAL/kPuYbesPF03ZgQ9BdRVYg3AHI1eZ/JdDjGI/H3Usofr9ydpAIA7CE
QM2Y1BuD1kKRTgb3oFcS0p1tFcUjsiD4RerOYpHKbtbeyf9/Qed6k5NT7XpqZ7bG
+aBuPa9H1gMfnuzjaO3ZaS0TtuKh0yzq8XW6T3iIMxF9gwlOLsjk3pY7iokKh4jt
2xJYsBbiBi84IGOr7QKu29jl4UhiXoGHOY0ab+kDrA2Kz+/vvQegOk6qva1vNDuV
r/x6pjKRcRRsRBo8beL6i3X2dr6v4HSXC19H/0H3O1OtENjOLzcAYvni9efqG3or
LQKxr9fczHttT3LcAgGq16sCLCg76ds9jllqOMmMWZPqEFwyCqV+DJRXK8puFWe0
51FlGwcGjYuZ6ATFcwnx4iCvwPTpLmVaOLMSPJdqZNYRRuh6OjM7YJsBnJh149XX
amEyoDoJ461Nu0Hu8dGmk+oUU7JVmUnlNTxdX0ROhLJsugZbKANcYF6Uqd/H0G8s
fVsd7DNFLpIuDvxi7hbjtb+YSt/eTqkOLW/UsDCf47XF9n2R1q1CqqrDrCL8e2Lw
sn4fTFfFc7UJ03VxSoAQBt+5kNoV7nPw6ieyjkPXnRvtKIZwW3qe8lMrTRATwwOM
zOS9DYmi6G+4Mqe42sdlSIScNq0XpgqLqCYSMLT/hqn/ruZTnslNt6VBPGWojd3Z
DBZHtnGunGFx+aCitAIwXr97tCBltyaK9QC0kCWGC5vlDv7lVDaUQahZR2NQUvh0
SaMWteRiUoO0Pwgt0NcJMIjMjgn9xtpLhWYOqYjnL3+P45Q5NctNknQCDnR9Ctis
mkOPOL5PauOFAKn24UkNWufnGvkW6SBAdbgX+SqwDymtmI6lyoWq7ZJraxI8Wr1B
Ik8rwUfwzwkQm76XmJ0DSQJpP1rF6eWm8In8b2aqe9cG8Tz3GBRXT58skg0Gkp6y
yoovJu+3o4Gio0qNAzZWwZ3sHuqQMWR4TBX6W7oPLkzY85pfY/YcZm38XwFUkC8z
bNcIGd2DOEzMZJJ1EAk50zrRcyRki1GgaegPXNbCNyMAwhpF9is3YYXzWUMu3U0w
KElV70d+WKKUA1eoPcZa2VVxWlANr0wjAQKJeVINss8f8PyEiPKx7hV8wsKFDWsx
+fozzMwqaSU3QLKL9z74Ra0q9GDqaFPCLDTH+x2QAppJRpXHGxkZmyiuwWnA7Jqw
lBFJzTH9Js3On0hP25nnx/LgZBMKuRh2QEM2umVQehAFdf0kA9/sBGlgjoZu90ea
YvUb/ReA7Q49IrGym8JbABW98ooC4JfuRTKyT6KiNOehNCPX4rgM2fx2ra2vBGSO
rAN/7RBDoQAfi+FxZx6bGRcuaz/QwBHo45iX5vIwd9pq/+dcsj8/d5yWPwdGRVvT
s+u2KyRES02Jlzf+c0P8ZTabe3G0/vD9z7VJlURvQ2xo4072cogba3iwP2DV5HRP
1HzBxwDUo8JKPOGWJUKVFDlcl23WAeLOI3hbAAdq9VhGfqf4rzeczDZRrVyINHnr
wxN+UmFLJAcdEYRFcdii1Oite00Sqr+xrT5T2Bkn3bLt7hU+OJekD2dP/XgmCpVi
RSoqo7iTVJyewAu0Ya3qnEMyB+gHYQ2rg+VPiEhkKdEfEV5vOPiYc/KFFR1CokzU
dyB7QIqrf3Us0LWo5K8/yRmx6gBLWYn/rc8bF6gR7IQntW6fRe89l34OLAJh5vFE
NV4AaCx71dzWIKMtowbSQ5MDZ8F0P8gDWevqUj7RjhB1FgDE7kZTTepp7uA6SdU0
aCwWYfwhBgEPZ3nJOnQljBaAJ+thaSDkm/bVLgurSla6bgtWex7ed8Pe5ZBhOUDg
5s/2iJ5T0KSqptV4Cr6LP25jmYkGCwpum4kEVp5mN8qJTL4Xb6Mc38AkJ5NJPSrB
xhkpZS2vinEEjmyyNaTgDa5FwVxstbLKCFvsynB30zD5GrXQDSRQtf4Ri+K/WNPL
Wt8LKhaUAp5yg4kl6ud/edhe9mmoxyVy98XYV/xqV/A6ZLjUPR3c1NqbkuInSuu8
QG/dWHYD8Nk53hjoSwn+MfgrbC/dngZdGdMK/KRWOaQ32AuoarPRQdcu1etPFclw
hYdRy6kupTx9Uw1beG/ajeBCWdl8syUHRq1PiYYWaxsc5Ala/BJNVAgDafsDCC6C
V01aazfHGtqHAfDrBxxo7MndhDB02Odutg+IwyvkQCpCfqa0SrpxXqKLg+diuUzg
eZb3QgF5pkyYTsV098OI6C8zR+mfDJntdEXx2gqmn+LRTBcE6FptDAajCWiz6RHx
afC69awS8v8LJ+z/n4iJYPc75VoAdEAZhQWu7KB1V58zaawRKWVj06Mf6RDQ0zNN
/jixc47GUAGWad4ho+Aom9ehsZq51Ej0bEfrlAr61zHzhdQeQRWJV9ToLG1WGXfO
LegPTFTDLs0OIF8tZ/AUjbzL7yeGF+0Nife6+x/6GjVtuoWANbbtdEKeD950Ot7B
ZosEJp2Ln23IqFRpNIiw+JwOAzOVLMdTj7OoQG8ImzpyUdUqdvXaKbcXu/nz9II0
iglUaUatHBI46wyHQV5XXz+sl0jyxf5GvX0aNYY47bi7kcv4Mo9ic9JzMITLAROz
ldM3eWaqgCxIlvBr8+UZ9FAHM0l+3+juuPPR2pQrp9GdgXfxrpY08g3BbPIDK1ea
nRoVb2KsiSgXbqzvfkVxDuvnGVjGqSAUdNsdsr1OkJsJHDoJP+XmBh1fgMkc4BLq
tDkKKJx+A6MbGn8IuA7CyLHlxBqPwGscjFT+W5fKpCRfyCZj2AH0DqkKNQ4m4j5U
fCmpth0H8gOw9ZKjbQoekeObnuiFqH/T3kJh6Lyxccq1po4wcimTteAOT3qCl57Y
RZsjlepMbAgFECYcnLlidu2mczqSmG2LYL/Rpzh+vZ+nPLgG4+MHH2dnq6UjXOfN
shsifuIF3F4sxAPgrIiRQf6NAwhXo/8n7MOZ04ZyIcUzi4QKQ5LIP7rQ6clbpFTT
x5MjUyH6eB8Gd0zDOHBFomfL4ysuS+lzO/5nlLpQHqsND03R380Mj9GrvVfo7A7U
I/FxKcwFDuqaHc4+XrvdbiAeRWWw+emJXFVGZlcZtzl+SYscgGLVSBsyAI757k+B
Yg0Jfso1wMfxt9yfCncCUOQJF8BDHhHoKUCPVKugiYSZJVgifOTvsBflC54c5Kad
GmBqmReULt9PTJnOO5sqM2Yy0IkEgw1YUIa2Fm/AjFt0OHjv4v8DKtIUwhHPu+3V
Rn2zY2StOtRkV1FOBAuMVrqxRdaWgTtFfmE0Nrtzq630EpCYQMItbyoA2PUFU2cy
E6TaWcG3m3BzkmmGV2nAM4GUEo+vK+4qLOqBK6/AQTqrUw/nfi+aWRJ0mWywLpVE
uqUoJDyLc+s+IbQcO+U392C90V+0EFjB3WqbdjGxYdUhZe/YVeF5ZxJFHfNYKn78
Ro8yroaaKeKdm2rHWdySKKZRB9c62tlLNqLZq28q3BhgaiSMypibHP1mwyg2dfrK
bnhQ+pTzd+JzrxhjrinApJq8k9ZzKwdjjDjPv9S9mUs1jX1HNh2u5fxTUmcO6tYk
Vh3SkPs0kL28wpRA1hdZb/eNiy5aV3Pa0ms/1cCMfn5jk/NZ/cNJ/68HDg47XdaA
9Ewy1QBT/VEoK3AjePXyaUmAi/Tflx2UfcFBivkaeheDGMCIGsQlnp/YHW9pIwW/
Hb4AdAsyxeo6Raklxa03E25vkptt9y9T5AlXn+i0YGr542C2pzf5ucovakbkvdrc
14CJMS5/mh3lmMN8k48i9pHVlWqHrgmYmVCGQbDmYbusOxjmo/Q9ICLdEY7iyxow
sje7w5eGvR6RrXbqLr729c3lRqjueFUx4ENfRBz+fI+AVRTqT++uIMWPfL5B1jZM
hGvcXhvapROkMNONKN7j2g/26B2fVD566MeEUkjZ0ArMM6g21OezEL2RCBC+LFG0
XoGS9t+AtYhTs0CeNlSgMY6Nb+tmNmsSw5UJz6NK3Piz9O/z7PqL+sfwBNv2ujzk
czyuu7AG+l7fj81cCnnRKCOOmu36yWh5EyKh5IEO/GTkDIyQ+dX7Y5HNSNHn5w0h
lExmxuYtZ92riM6HifrV79ZjDZd4Rk+guePvQX3rbJk6jd38cL+XtU68aclVcUJO
ssZssi2S1oSl/pj8HDhYeFoSRd2/Vcbvd+9BqtJvU3tx3HLPWXlUPkFSgHqdebH+
0eXDPLcwb3tc4G0GNB9RUWha7C0e46cYa7U2D7HEPAt+EVf4RpZqkcjV/NfD8+NJ
/S43gK3wr1nb5UY77NTufPHr6yZpUBQBY515S6SM2rB6NQ5iYk3dq+uZ1ilpsIlL
TGA+9mwhTe/ZX96fPRpXSxCbnVsdykHDDaSkT1r2fHpSv+SDAanorL5EUnk6w1wq
UEYPMtdXbsVBYRyrmucJQz+Sjw/3oEyuehFwOWMVSN2EIv2B5m4D0xMrsZi+t03D
GHUf4CpKNnZ3oxdNBWMCZ+bxjr7rMvt0SiaRPuS+3/t6VV1XrM9S2gsgc38i3D6w
fi1ehmVYMrgRQWa7c/mbAJgFWQVaoGzsw4Y8ZZ54C4zjtHitKH3pLY4zpPuKkHLa
8KZPxp2CRj2L90SujhKPc/bjEb5LiN+bwyJ40qm8LZgRPkgLtLiOUvnutXAc07p2
fXtJgLn9O+324HilKgsShaYtoOcGNdKIj18eN1KSNwJ0+WB3KT6cR1nQ8Oyd6dQC
7ZTjZTYX4xKUM7bZOY9Q5r6QuCCnkejNd7hWtDkxvLQjqp/IEG+zV1IqgHzYxC6c
zMwRP66Wwv4JMUcoD82gPeLDjT7LxOxueChlu89fNcD11Pt3kR0h+b7bzbgeIWhC
5n9WwCu+b/cK2D1im74nQBuNEks6SjAJDN6z1E+EkxvuRzqeReLzySdXbncwxz9p
rzS6DNsIV8RHUDHncllkYi6F7ZRS0limwwztCFOr4BXWjxIkjyQQCRAwxIiGpZPF
Exr/5R6oXEeneFxYh339Ozra5zO6WPnTdWmICfLUXdKITzvFGWoURPhzBTJIh6cD
tL4CEuOjF4zbs4tvnjF8Qq4jrEf0n/HHNG8ZOax7bfrr8M8lTwMi0DEE5oTY1WW/
0PXsXneXPLi1+EotNCFV7G2mz3/KEmQUWjN/B1k1mpxx2XfPjotQqq/Q6sGwC3sE
0gWW8ywkU1MkcQy9RNa/xi8u5d5APnkdlbP+xxpglja4MJEn+MyusEjl6C5Elt+7
5hO6uzCyBVgCQrvIuU76WwjMqqNAh21KnwFQV+1DvoD0nMzwnF+ltRBieOckoMwp
uMkJ9+VAnmqIACQ8lKSmljQs7LV6IRZXyRMA/DQKc9mZTfDIX8oP0ws/zqNgqXWN
r13CgdngEC+tVtKqcHN2jzt6B87JJfMDqh50kS3hVv+HxAjK8lMPyROE19D94Ip4
b9pU1lO17RVHZ1nTpLws4FLLUnP4X9spD9slUklwXHsW9fsYGTMefnVcp9JpKJnm
DO3ZXP4/E2TidYnERKWvtheqm3q40e/OUqy/AmHj3u/jLTpQgAWiwASm/SI7HBvW
yRK8KdssaSAoEKLDw4a8SFFtPpUWr/WGhh31BNjYzpfcEE4bS8DQED2uNs/YuROJ
A2Xdd5MLrdSBpGhRpzYpttzP9XrZBB7mwIxhkJ++SaCTINnIE6XmTqvQWruLxTCR
93jIcT3JCAGFumtSuecQn2pcgWHbIhX6vbTADvzQobgIJBq7Uho92WnArgijQOz8
650zj/neGtyCMjMyOdfmy0ZE2UYtFm0AkDhBmkAFRWYlz7z0cD6o/On9Cx7RmI3M
5jjszerKyWPQQaRfwuVtHKqmUdhlbJCu8YYm9PV04B2oJ9Qyw7Wd7/nFuhk/oRbn
Py41AZiZSMVt1QqeGz6qOmzYLEb7BTkcnRixlc4rhwIFU85u+b18aZhvAY3mTksy
uhsz6w3AcGpSnaKIaoUCybYS6NrXhiMNS3XcWYp7skq1Dcj9ONIEXlWBFnLcs6R3
+WL17qlSVy40qDd6b3JrPq8Gs3CKUjUlyKesAL9mCaa/c5knb6httc8cPvzA9Qow
O1bWK3ArLYRTkkng4+IItP6wjF1DE8CrxD5AqXjX/weSUkrQElEBd7IokuGD0mag
17NagXXxioUYe+m6qxl2NrmhYKTzZC3VVF+TeJZ49BxNnnJe9DdiuuYAcAVIE68g
AIAxbGFG8Eh3ieCoalveAzfntagozQBsnrhnb4bthHER08XSHu1wKfRneQHe9tIS
q5zcxgSKuDxEtE9PXKpZTsxdDtbJz6FcXVD3RMatKKyhtf6RIw0khqYU8ycQRKS1
Z32r6sG2/3WhUOWJZYLxbOqyI8rY+a+QPaQHRfwqdUe5ydgZxSwPW+DlQb1VmRbO
kz5JCTphxMaU/FrJR+f9+VK1sf5IsfrE5nVN03Ph1wnXFwaV1Z3BCyRA7hGOabOv
aSEzlcXeSYDOz+yvUABeV9opbGlsaTICSj/PzciZuhoX+HxRxSVC/8OIK5UZWb87
XwR3ArRARdX/Kjk9JZjmDfWE3fy/K8yf47L7UXd7+raaK60p1pM6G9lCFPLkoYV5
y//LCEeISPZn0S+gsdQ/2wAx+uiRjDXlo/qeMhUh6r0JEvwetnAn1jvIG+zgel8l
aB0T1TzsHJ/fy4n20pWVLKl4mBcnOc5dwHKzAXhfwAQxeL7X20cUumZefeacKCAu
flmQyU8RlUjobTgkaOpHCf5IzRhpCWthE/b+G292e6EOx+UE+nLXsW4R93XapXu+
W6gqOqbKPYQHOFoftxIlnB0jsbKSaUzwqByEFLbUpmN+YuGKZMZfkZ9P/csONLj3
j8/IscZbQL8z/p+ibPSAk2S2SqVGKAUQDV58VjdzAoctzMO1gG0wNJMgJWJy3dNX
iojEEe1R3FSm7LGoM2JqqdirLWoUM+a1/pF/i+CltNv62aA9WR034ZWyMfqD41ed
bku5ahsPnigjItcoYw3oLF9CPxWFYOky5gaFBV0dHcaxBzBQP5WJG07Gpf0FQa1r
F8k43WeXOoKD6guU/L4Deu1/bcZI250Ptf97E4b/A4M9MTZS2bxHB56QUnVmxL5l
8MrvSb1tqi9rXeY9m/Xn132xLA338V+x1rcKZ8lvr/A5BVUoJDOpWXzjbgQm4LNT
ibRQqDYHv4c2eHsweBXG3DekYjJad0kUGRSma46KE7OoMqRjQFTRM0lwrM5P2NWd
7tAlqCqNotS+GCKQ6XFhUWyUGoHAh0FvdNuW93OzlGLxutNIEnOGoXrZmSfSJXSQ
Y88WhvZBS7mwu8prgo0ih1csQ9iG4QYysBw4+8YPcdCNJi7TuKb8H/w5AOtL/qO5
a0kn3gUVewDGEWnCslkxs5gUIBT88oSlGYjiciVt5/mXW+7YffJTUgn2Spc86JeI
zbezBR9o89SkMFEBtyCDoJzZ7OJ8ErnV90B+WvHjA4jagJd6T9CQKk43GEujmRJR
pw2DIMSr7R2OCDqXP5Ux4oMlVO8/RtzW+5Yz+umZP9wVTBQ1hEW0OKRG4fNxkxUo
AxH/wpjWOOyugTOUGcRniqk/nLf9duxBloTijjeWeBga7kNU4l2UNS/RnTpD3g0r
vg2moXoNRRmSdK1JOICa3DQF6TxNTUpmNabHtuvqk1FPT3Xw9Alv1arXTTRwSerl
TQCwu9HnLpeG6ju2uFcdZ4U9kECyF+knHxeX0UaIv/OqAJXB3i3IPwsyOQ9TyALq
MMes3if8kqDb6IOGFf++9/TrlG3GL9d+nQs/3zK4/D8TuPb53EuX51FN2wiYwfns
JKZ1eMDgoyd1ufIS8RrfgmmTWOksZb7+ha483bkpfKqzpANuozA0qFV6f86pq/G7
a9LtBBdo6GnWTVxvrEu3bveaRbz08uUEadwTS2Hi6CziFq3mwB/D+KjzOi43Aj8Z
grTa4WSvr6X+5Je9v2OqyiT2VygdeA2wRgYFClaHI4iWYDmdaVEqkUfXR/dEx0Vi
wQQsmNs/jU7hJz2FS1q/FizvZOdZVYhyKUredxOhzn1PWVHjlSng3/kSmw7PFqc2
D+gc5FsIraKLwm/VP/QKUEQQengtuarmcC/NFnl/rnDFrxSPC5cDdHekTlBZuups
DAmxOuxZR0YuvyfsYzmhIiozwbFdsLxIXH9aF5E7GxCl//89pZRUeaY5myyApORE
L00nkSeH49s9Io1mEOasT/K28Rgzdlm7ebqD7L6rtxGv0snvTmijGi8mxYAGH4aG
Xuwi+Vo0z4HkkppTX2KDEAlqcuC0Mk2CwOY9U8GAsqejHYKrWeSY7aHAeKTMv9Mb
bCcGk9KcV7gTGZg2oJqqipsT+k44K5Sc7oZjX//EmtflDMlRzPtj4BRpJrLBep/h
klFpzC7E+dPsuYeUANQY0I2QzUuH4GvVjXMKLdVYPYxRxYWI09wrIa4U+kpCE1tZ
4cZxChIO+DLbtgqLOHTWPZbuTnUdf0xOWJwk5NbrFUHc+lEwwRbzuisEeyNXno9j
CsV1XlRCwcz2GQFGQssExBG19V3/V3jOxnOu5GbbRKDYqFOZ1C2nIxjQPcqFSisQ
VJMkb9nR3jsMEuuRTgOsU+Y0mRbFc3h9dX1HVVRD+tdhmSpvl1+Z8gy1kjIP09BV
tJPeYY2Yex75gABRhvpCA6x1gSiWcD4YDmqTz7cTrw25LSeJHAk/BzzD0eKViZpI
DehVfLdr9PMLVtWaNCh6wceQ7pHycawi0lwhf66SOKl9vF615m2Ugq01XdnciR+E
QG1/DtuyvQsEf3bMCDCtF+MhkhUqjgbbXWlUSxZzNMF85KVJkf+HvDSwYE0ivxtg
fn33ilIk49jmQdbirt/6cOfygDiqen+KO2CRcXjZbtynzqyzQxDFFwxFoCXF/tIv
UlYP/26vNd5JXBdQtrf/anJ8w0HrXoIft/NZT++ABA+/K6lg10fWxfrbO6crgZMe
c9fKg5gZyAHYthJU71gzpBotq4gkUu+5rCd8grdk+PQwhoDln7kxzAmALHb6Q/+7
6tI9v9zJ2+sypFNxgyPmx8MwordPDoOEWoM70GrBfR9thlHpwmSO7cwgpUAA0lcX
7CoqEjNPJqGtvvfSXxV6ezOteZTzig/9Gf/9cBKokYTzqp+NmBIhZVVRm+HV3Mvu
TdgpSYwTN0U54WQmrP84xg1H+q4O89N3T6KoogGJcrImjdBhRlIypQrkGGPyXmES
JHGp4icdvharF0s89wWeLa24rdl5DVJATKV/gPAdVs2to4hUkWlOSpkzzx9XsBT8
Huhk0YQZJNYICxQWvFcmDUtuIWUZ9WQ7xXa/+zmvBWW8KB4tq+wampJJYSUjzHv4
NmrqY1XpADoGY9cgUimYWED1xEgUiY94SnFvIi6llUTVAcqFVyuAC5SHpMUwmYxB
41pIyJ75I85m+JxzGAEqBv2NJ84TbZTADshfIqiUZpuGMHogNgV22MLtmBcLRMLy
GmcbgizAa1jTTerHveyG+276M4lg33hUhRGCzYCo3dGhmBhw6WrZXNR/LppR1VNb
WfyxdoXk2zL/R1RHxky5EaST/IBNu8zjnILVVpdA2/53mv3W+05BTglv/MCR1TV4
1cksHHOZsWrdFyDdlXvtqhXgyKJtTnHCnAyy//omfURj5qEcJ8P+ZreiQNgFLdpt
fGL6/OBE15Kc2rDzkP8+0IdRzHF8sQ9g+UDjxoAUqI+nRGBbMl731sYOwUWWQhy7
xe2xOCZXNrUmLTYpNJ5ZEab/0+RY/3XmyOZ6Ff1Y/4HSCoYFLmbUDt2Go9/c3Uav
le3X78D4WFwkwwDJBunIW8QlJuP1ygUr+NtKTWLG4WlDHVhn3Z60BqRf303mXs9e
Je0pWvR1SY5+N2QBvuzo9hNEV5/d2H/UThgK7MTjhqh/3lryxo+NJFPSNe9q+4wV
hhYM1/klrGtwhWPszxqJ/0Xl3urj5t2/sPkQ5DROSsdohpYjuS1nnbH0CKhYwVUB
iYOLp7hwLGqEIJD5iV1D5nK+fK9lWnK71HIpnZQ2M1+TS1JcIzdSx7ZVZN91Zm15
maAtZKJhBUQl2/apuTzApNMsGAyiz4J4GPmqm+R3dzsM1+Gin/PLzc0qXzF8qvdh
NXFYqRiBmo8n2NWR1E2L/dp5R0cQkxUXY/zor5UYdeYQEPWMw5S6c9L/EP8ghUpE
abhtMqa3Ou487LqhRvakRh/QofE6Am5YAURFULU9dn3mSeVY2Hna51BpATAZenAH
0Ui4396Kl8PqAebIu/zTl7AYH/5BADEHGxdSYN9o4kUVAtTp4P18LT4tC70ZhOT/
gAz4RY7GFDxMhgVv3vbkLgiQzf0HODO2kLW6e4WhX4d0doKJEwip/tk70HGT6oSi
8Wksq+Qt2slNcT/uvU4m0YYMtTUtzG3qfA5rb1gb06LlDEGKY4ZVEl3iDtxBnww6
pkkPo+JpAZRlepcjjkps7G/rR8LqAbeJLlzyieisymJeRRzRt09msg8FBGe/WztM
QAzk1OPSCXjzcWNCfCR1gDyOzKpbK3bngi5E4fVc4FdMhiYaGXNoQUXIsmuE6w0E
E7DxjhaoKGSa/y15RRfvocX9kLKmH8MTddjjV0zuV7SN3P9G8s7tAjvLIdlQZKKs
Byy2PIjxbZQHkbHBeUBzJV/PHfIBejnunTeET5wrjCshTREX++jOEWPQ5iWULtSi
UvT/FCIV/BxZtmamgQdkzPIUQYcYZAiUXIdSpoMP9pGgSPfGSTOwLRA19PM1IptM
a7l9g21YaV+p1ZTipkBrXKvO+/x1aTHQX7Jt47dn/TvICxZGQRPbaY/VhAHkvM8E
dNMzmxOhVRKbBwNhmJxytvDWZUonMu4GhesXPWV2oSmVxjmgozPVkjFAybMa/DMj
+fns/55rGFU9JLIqUqI1ta5o4UKE3tVKTVWkcZY3SU9+zOH85BtnNThsLvwvYhc9
BHuV3IpxS4RDks9aAkS930bH54uIQltafNpS2DWPnupsiM+LijY0hqxED8jX/lta
PgdvYeHLgbCV8e+tLz8voyr1SOuzKJOF8nLLx4hjwY+GCFc226XIRsbgtzYitlXU
lEaw+YtC+UMsKdjeMzVhZE62Mt4Dt6QD7XSPL4kb0mqGEEKdTtRcQL53wH7Q1PPm
BAXlQq/wCVSIBXJXMrMRA7bLmTgkjyvMBhLVuGqoyCufD2kb+lB82/ghXyBOYGW1
+4Gq+UtmQHtb7cHc88Bi4HZwI/C83CTKBcTGFH/9MC7zJOG6ib+/ySNyA0Hgc/9j
ptLGqYB5bA9e89vzvCMGeERi4lAxG9R4sAbu4pQllUxzLJLjGlLyv0P9weOVGNqV
6cv/Z8Gp/0KyInBikgUOkOTh5SOqXt3GZuwLiR0fPHCdJNDf21PE3i8R9+luJaET
HMdWMbOzuUYi93ZJ0mZvN+vjzz8NjwJ7VBtaOOFRhQRiR2SLWG+rBHHp8vGMH2VF
C+uFvw1jAwZN1JaT9KjQQFJYcZOQZp9G4MNIk3jHPxTJWUooSM60/PDMryU7MeYT
U7FoBIc1Wz/1y4sodRVOhmsXT+kKoyTjT+WAvTzhObnzOTGJ+ZPmuoZOU1cTY5z8
fpx74RuAsT0j1qXpv1Hr8xeyhJGWXhhYSfCpKAuC5+fOlhd+q6pGTrBH0D0aFfN9
QfFd12HHxFGqJv3kkMpM3YleQI2WwEiZs8jp4b4uNTbUhDGjCFdRbdp31d7PMJyq
rOZ7yyv2TLtBTQB2qSHpC/XEIUn3P1a1yoq7k1RKFJgY7aNYAPSYt2TMjiT0n0Cf
egOYM7s8tnY+uIbFlJ6fsL7+05jkYTD23SV5ZxS49wJpmqFlmVwiEStMjGM2bZbk
hETkZ6gFfZ8jEf3Vk0BSvgvgo/xhv/cuxh00k5+qFrlfIfFjsRWCG4i6RGrUduBw
C2qMQ+f0R/RPWbI6sjtQpijbOsH7aqhV5AUgUFLJB7+SMkoS4/9zp+JZ5gZrDxGD
jhGgrGWEZs27s/Esw+VBAx0Mf8L38LAdcnWUlDDnl6ivSPr4lYKirGToCpunwH0e
GrJsS6Z+7pIcx02qDdH1ivmy8lvGupfbIB29vLvvJD6DxuaFWo8Q2n0X9+l916dq
+hi/CC3Jms1wo8YJyNJ3/JSRdgzds3XjzbZZ5qMd+okM+GpaEXVoQAL8M9Cdgu0R
BvH8uAaOXqlw/knxAo3FZxIG4Lk/7Pa5CNjGlOKB1J5DaHKqqTA48o2UFOszZYq9
2MRs52icr+dD7ZAZw7QaxD4QPTiHKnn5CI7i7VulHglTAQUfn3i4y00CvFY1gLh+
bNV3Eow3LZLqkWzKTufyMqVTrIrZ6kTPRpX1mu+r0/W7HjflnAI9Oef+YW6U/nsh
JiBo9GEdZxno49kAiCfBPN1Cdq6Xy1cWdX0A2JES0hG+n+J16EsxHvZeX/8S4jXO
2P2OvtAfM59uGMennL9lRm3YOxrc+/p7am9WDfNuKpGjnH/P933Q+pbQT1xMsNNG
Ued87JRVH3GMCXc9ERT3bwMZFdcAv6pgNL5n5/je79ciKgXX1L6auSxTBWkJpFHL
RU2qvHm3QX0v3lr8R4mOyX2fv4NpfJv8c+m7Uubf4yqhty0Xj9A5iY7/DhIAwgOl
5SzErDlOjPcSLSLIUbnu/1uqZ8ZDY0MsL3S5WKDCVNq0vYdMr7CFrfCQOqwTzHii
21FDKN01TYR+kszLoYvMX3/6bjBBv3XUkqgonh0gnxvkuYT/lj4cGfbGLUOuvDDJ
7I5pMnBjdD41LdL+K0kAdERXXhCPvvrkjL+RNscQaqDOU86dM7OCyIgr3TZd6qbQ
KPDQigflYbRPVjvnHKY4GOdb9PbLP3045TZwjmfVh7BgYP6/JnuzsTWNQ0WiLEe4
d37jWuzK0cQyuBnNOHHvZQMeVirmyVPCHM3NDSKL+M66RyEudtDMeKmi4BBV1sNl
DvK3CYAbOfErglUEVndIYzdbBO6B5Ma1Xw7PkjvFyK2/HRayJ0Z6gbfd1GooMFwn
Mjuh9PY0Q4qsqXAJyMWk7PGnQ/97NZq/Lglw5sVfICXBAtYKK4mN78aWpm/E3uE9
3p/yvVtPl7nyBOUINBAa0Fp4uyERXiK/a9/AqpLcVspZWWxPR+TzdlPEBguFlaPD
hvw4yDPIb539dHSWLW1MI6SJxJnakFNL2BnEEdkvI7l27Ww7fiYEEbc5ZZwFkOn0
WXEsbN3PSkaBdjvcyW08nBUXPwoFV8fb7XpqA8Xjcz9calb1cA1H8Ib740pRGZJ/
uQp6spA14CLPgkwZhYA9i50B0Nte2yopEBBvS62gTkykKzZEubJcVfSt+YL5IVrB
lrQg4vKFHOngStg+JjGkjytmMLOzpVUPgrEj85uKMgcm8X+EffaC+2pJuaG/zlB7
kFlKaASsjj3qMPS3P12E9ekis7kqEQ/pxq1XFRqhrFMVMUaeyqbbAjIutGicBJ//
839q/+AP8GngLBAHI1rtMfzc2bJvegkRMhcJOXRMNqOaWXaMqtwoMkhHvOyvRdkd
d9NFKN9Y6pYZFdrW+DVG12ZJmYd2bP72wlwVk4UK03NiQaZ55Oo+yZljuuVX4rP0
HNMdA2B1KjmmlLd5NqCjx3Aty6E9GXvPOJ8PgwFibv0YXvvfFaBprLSON1vfTGDc
lhdSLHMVZ0PNiaTenk8B9ZtSp7X8AcvUqoh7LpHlQhOiR+psH4MbcHbPwb2InbH1
mpdZ/WGlz4PAPvzMJsEjTqXXwUiQeGhie/rdj/wY3SXZPdoU18DH5RXQ1yNWpXUJ
WR9cqstY5xqkCmBOniWXvEfHlqSTmo4cfF62FrmfytptxSWhr+tbC8tXmaxIF8W3
rwR4yp6ZHQgXUMr0Y36viMlVuH2jQgbJQiGwtb47pC403xhvYQbhluHLTW/5N2z+
aHq4kTetRiCG9er0XZLSlVbdFyvDi8LAP5IKT0+alHQ6xVDMzyNkg2RVzx5b8ntT
6WtnW02kWyxjkD/GxapImuXfGXYQr/LGxAclMg1VGZ1/Iks98+pjHeeGKA5v45gh
jcRBmQuwSO0zhnEk9HttZB9H+RwSi6BU+OKBTKjPKld0wDXGKuOnFNChBff8YBTq
fJtXymBHpv8y1Y8xdo5IMmEnphKYRFJjU+GZi1kzEM5LpDtVlZE03tjt4wDEezng
SsYesm++H8ZmBXKzpS0lusmMQWJSMEwHyHqQNRpIQ/+EBC3xtHMIxS2a9dxgwUPb
6dMuMEqleqTA0H1RBNr9EY4MNoEzOms9zycrdx3Cm8LWGFA2DOWlZfQb1KcuCnOD
38gY3+4DwnhOPgR41ehGC5rJEbcL5ERPEbFT6wADUipf7+OKWL2RjnCiltxfr8oO
X5ED9yJ2g9Y/OjF08GW/kkNbp1Perdtsvrt5r40+gsrkbCP1osyCLvO1vX9SGtDT
gfUY/JRpMz2zXrIedy3Wa9OlIkZrhT/K83NNi2hRcIxJqL+p1H0WB4wz5nPTxTFp
d+CslpVsuGaI28kdR0R1kb+Cx8AcNWVUGJXV8ITpe0gHVsQaIAUS84kt0GuAxVmb
T9b/ufROHr2CwqCddVrfrpfUO9yH84kUxLVG7v0xX24A0+zJcXk64KeYJ5Y/gEz1
oeZu8nbEfilO2sJdyc2QVbJF/xknAIf+NRUIvTr/f+hGnbz7gxpgVB58XIiuyawC
hsFjDcnfZPb5zo0xafg8PhPvNHFZ5kLEQRHyjwlB3uutceKTtOvf+MCk8FEi2WL6
tf6jgK9JrT3zMTafOXHw3X1iIYFJpIiegtFxyUHHh/np0IYd0oEVb8XYTKju1as5
C9VfRJTQZOaYjCSBgaN98EVg6nh1ZL8VY466oe1MuQtpBeHHkE/mfCTwbvD0bH8p
oAHk2uku5Qu9bIGI0rFrH4nWIVKFbi0IAZE73KELjEpen/ZShTXSPYva7uVI55uA
dUMTTg0qHg096FAZnVmqcl41NWvmrm+rggdeIgf8e6GGzjkR0XeJAyoV0+mcgMuw
uQZoqGOaky+aC8RfGoPMJzRQq/b8IU8onlUYJ8t9D/NyrzANwh5lUMGEXk07+ukM
fCnf1vD4YcwB8GD3PPaoPdnlKb8r2B4P+FYV+2EPPVoGHsXgsUT1Jp2c5Dr18l2o
tNkR1wefgwsm4vwgqRtuEqsNlau1spXRYCw4Y4tJXeykXGCq8sTOWuRCX0aWE1Ue
N7Pf6xE6qDBmDvkWf21WcIhDT0tIPEtSsOV7nAjQixj5ymRX/LmiGFoDZ3Z8fIoZ
tYx/BKyFgZhTw9XESQ6LHNIw7WO8T/HQ6OzR81cdE7y1uZwSP7qYymaZ+qjsdQcS
dUdQ8LeDWDzGS9Va399O8jZ5OZ/QJh6tQ2J8nqMf6RXV4fM82eJ6sf+4D4sXaq4Y
E/1cpbOwMr01bG4AqOtZMFIpgchECF+OPIuPgenfQsXX8Qk0RSp19vQTJw2ORlPn
UjCUuLdBaprkH43r0FyXlGjNGKBIMSY551T/IadH74iOC0MSQOpY7tNPPOMK692s
afBF5uc3OJ3tHoeMl3OFNC7AyHuY0tuEBrRratGj3gxch0Yosl4vnyseQQkLxqsk
hMenAWirlYjpZZoJfPNEtQ79OYXwkFlBi9+oQ07K88Af9DLaESRyMwtHdHK+niV2
tZUU6Ngr21w1GELZj8vS3SBMU0GKVNv+ihZbmLfIxDuqbisg3cUqfxoV4dXxkMhi
DbzDHeWNKYSt/dBK+HcrQzLJW04MlC4dKpjbYbAdPne+wOOunLS7AKTDiLmVSrkI
AeUaDEN2pJcPjTGhnuD4x8pOIOA+14fslWJG1JqdDOdGC+iOTQxPNylNdqQ/rf0q
tRGtc9wzVrSbPolsx1OwHC24aVdfzwAoaSMlnGqswNLlw1Z735cb38t0PF0ZBbjt
m7SVtXnJV4XjK+v5A3ZW9qLebhwmqy7+ziw8bnUwZpCPfYphVI23brtus+LN2alF
zo3NkN9XlECPBWaTxP/zEIelw4nzdIaaS1ECaUg1PT3L4Abx7mJGdSXmqFnXJ0L6
D1ecE6meLar515ZDkXIu7UmCa8b2Yp114HaZ+eFNAR8WxqeVOJmr7jnJYDr7CBV/
CAa3hCwb6F8QOxtokaYqNBeUP8M3yZn4lB5/ecCDEHJ2V1on7ROT0K7sORGZIPz0
FEgr10t4JTqr9DXL/2M0hj7TyAzIpCpu5xnI8QJXnwuc5bY/94kFohOiBJN9oEUK
+nJSmi/84a7cn84sQkPqrVgyqPgtfNykuekJp/sDqho5zJiiiwgyUiyrCh4KTIIV
oxROPaRulmq1XCe3NStriVeMDLsV/0kDShLlxQqP5VvniW6vVFfF8DVKbguoN4XB
+PR7npmMuoCdoiW1KZ+uDw==
`pragma protect end_protected
