// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z8ooq47MgAR7ydXNMEp9ocmdQYKj6/J332jTVBUFKKi8kAQTjjPaRqLGDaslo9Ew
b7lqf7aqQ6cfXIwjV2R6l4Clhc0ojAeRyJh7W19ihnMGDTu+hP1FYjvZFmYhYe9b
oVcdsnUFvD/D9qlq3xha/WtcHgu8NJAh0GLHJ0lJBqs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35328)
zpK05k3p4HCvWwNV9flc+7T2Axs96JgHTebt2H8SlMzditzkxkKWKlsaHEjaBHU8
uB76bBILr91chadiE+hCG1xcOSdTUggvi+ql52WAmwKEBsbVDHEnHFfgHs1qDSXc
LomLDOMYuYFVEwswxykiw1GgsJojnpYebyQOCsv68im0BQT1nOncjb7jDI1FV3vi
oedH+kh6W+N4gI7M5TqBbQWXpPKvKgqwdo5RHFTY8eZhbrHsLvavww7AH9UkE6jG
WJbncwdCAbIGV5VwJzX7JkdU1b82brJfgMxkHAhLeJFdVzxfeTyzMhhAlONES5Gq
KGPgpYNlK9yvacNV6iQIkdKvFglBCrvT2OVXR+P9ZPvblspPcN++s7bHuIxZjoMd
O+7wbsA4L85p9uEe/+kcV7o7KzrNA8bVgQBdjDpO4AQgGcet64d/e/4zNdCvvPmq
0HdPzcKfFOgRonLKP1ewJ48G9Ptacm7oLG8eKh5LzRcll/tWoi4a6ck/vsjORO0z
i7Z7Iol81TgfLO6YdfX8DsrlZTDaSsG0+Yii8dqpSYqCZIazHSiJVx9TXafTIM0Q
8A0b3uSUO5OSRZM/27tfO52z/3Rb2BaMo55+YXoswiVQgknQryklEEDZyC+xfwjo
ikd/zcXpm1VSGVkPQQxylEvG7FaQ9i+0GNsRYSEs/z9ff3FLEl3p3zIJDQorXZM+
ZL1dQM+a2lVkUUHXPjoGWolG+bLuKtf5b4sQcPW3NI5FczBY/cewGyUQrE+Lv85a
xUinw9Tv1dVz2q/nc2YPULB3FC3B+zxetnms/34rSbCPemT5c6p/+L35gTZXCKJn
z379jJnJroVt6++yHQvmp3cl8wC5vf8PsrxF6VQQ1Wlm2fPSZfpLgiCUCFTOs7L/
eTGDVSMyO02OOcvRlIdsEB9feF8AoPw0duxqoLuxODdRyr/LTGYgnPFbzjh+PucK
httpoV/yUiAi/l082ExyRpQ92kWWCMo9POUDB+YXN4VdpYxm/4QIJQCsrhXgnz8u
pPRUWIgwhL/e4+UyHTbzPIJ85SZZF71M23bgT7Ig5KUcVlwrGSZV3F3eCYGz2xfb
oY7fVKwI/SkKu5+G106a+Nj/sJNAe9CvUUg9p4iPTWAlYpKq8dwkv089yCBYISWr
XV6vtDzV3vB+aFpQ16ataVk5uT/LeSskLLq+hjlpVZQXwvHRK2hzKn82psoOTXCc
ypRWoOOVPcWlh0Tb+c7Aqu7wP+0+8uP4UthNxYsvZiiWqijY5mZtaS+Dy1LOpYd5
TDE/6qV/kP8RATrxp0MfEao6rz4p5aAXzlb1rBBceYliqSlv/9U04R9ALlDwr0tG
Q+HDYi767ubI0AnmKL/JlUjPyH21F4eigNPhjoVHUvLQ+vYpwdozujR86OmPdGad
BOL+B7IU6R2fOO+qrxm4JBOSyRZbA7psETxCMTZW8twnb1fZlV+wC9RK9ZFwOMzy
u88cfDu+dbsGvBtpVrt9Tk2b7hmsFNKotAFSr+SNt+4fuqOkqTQG+ZnzT6KPkJ4W
Ez/rfvW+lbhSJH1hIjXABIQnuQTCx5hWJub5OdQYAby64aEZK2qrDFThIiZUI4sS
8EcgDqU/fh33/cvfBJ4HUIYlXAnJW+oL9RTrTB4eW87YRk8RPU/Rq9jVDdV3PI7T
r+XjScWu/XSJ1Nxq55LUW9Yrqtfo3Wz1Yo2jVDTbpxkWCmgoOwtG4BrMjJiE+fI9
F/BQzScdnCrHiAmcWlBAuWUi7ofDj29yf7a09vOq+QsjnhJtOOvcEAWwfBCZWSqX
79CJ1c8HWikuKmdL5LqZO1bEoEbbDieOB/JTKPpQBI8oAR28ztLV8ij5yu9wVFNP
S3/DQqSunFoRcEnR23kcNSoNJh3ajbAiTFSHFmJM8QoNJSt/CbO9B60DwSvyV6j1
OYqox2Tx+7u0at1ZbaK/rnO2a/qS8M1mvnhWbyQk7vYZIouL4USQJsxRgr+UvJyb
ZEEakNOy7KD/nnuqYLQtODfVe9qTSABVB6GYLYD9rGUBSgY/yzXV0TYk22BqAPv9
KiSzLMU84XCZJy69z3kIYQYSZUKSX5RnOIAWJ2qfYzQmblFgo6RlH/yxl4FIkAkv
gxDQKEeu6JTnmNfehLd3GdjUIKXVuO4XHjhJmcS5MDiFhWnGsGNr4vw029BURi3P
zpo98b69vK7wUYCWRn2MsRu4s1AR11Z3lkDgyrHjtVwtNLg2T7fhbK08UmIlk/qv
ZzdiSODfxfOPqN6HxgXn+1hFRvTINGEaCOhWIqwUAQyHY6Jdr7QK15oiP0qGE1LL
XEqhZnx91E8KOUaZHkaa00srWeew8LDFIR1JwpZszB4bDR5GK8XyK0+dx4CM2qy1
mnoBT34UK4lbS+kKJUdWUDpHIvUmqMnJGU/DC1f5OkkTyx3xTjU3L/OOo4sCOChP
5mdbTw8vyNUkaaXngQbpdXJ/LALeBVnPKitSaC7nqjPCnvwCrq+9hz5h1yQG1hMI
n3XZG/C48Pvv3nvxJYCcnXk2lLK4H/BZPIkQBxQzI128UTXPdtJpZP9f9JQ3/Kfo
dNAI8VqNn5+iy9GIGcCehTDsZdCeVVTxmYzEaaPIlyq3ZZfrzfAIG1Jh+lABsVrO
JjdlYX2UtycvXWbzP4sre6RprAqw/OvyVu3DDLlrtik6Wu/HI3umFG+kF1l69mz4
QB5ibmfkL4mOLq1lQyJ2WZNZyLNuvYZRrKK2nyg1+o73Bg5M1zzfNIlxxTmg6q/g
37ChbvOty0pusjx8aX0Rt89pWsKqSmRYXf2n0XAeUT9/MhEs/ZN90DD7y5U41e6V
gE+OYXwQ2tbp+qrT6ygNKmVcsB/1sY9NBIIcLdJV1mLWmEOxDSIJ1EjUInUj/Nts
GHNWtUR+gmnSTThSlKd0T0Ii2Syu+jkXdLbJcZZu24Dy7PuCq0o6rF6I5T6xV6fl
ft50ZtS6GVj5WPhRxmlrCvAFdR3CA/Lyk88iwXxnxWH48tWNdoOdU6yz4GNZZUDa
QAc5eoyudKxSISt6R485v9/PJDpKTmwtBlmAHZscF+YZkgvwP9ZMJcRWrTPg+Jc3
KUrvhJMh30pw2qQea4xDNn+yRablIxxcKt2jnde0uIsS9Ipn9KvsUgLk4tnQJCah
szyAzs4FoG0e8kNP422z10xCOrqQYcKHDAdkz0rchGBt1i/+7x/GNENgKy9y9i48
AarrOy/cNE7b5VOeAXgw71JQRPiINpzqbiISiwJ20dhFR2or2NAk6xNYxO+AoIsZ
za0qwqkEVgEZa9UU1iRFYvFqSU7Gar5kvt6buSW1s1qq52lKDzs+sDXsasdbSz63
MosTiiHKthgXf7FW7WgkAHdW+7LK3EUAYHSnItH2uialipA29gtcpaJgMGd+XXCC
5VVGREnvyuTDF4UV2vyaRGttBOMEzLgvICsy1C3WGwmktddFNG9FE9MYwusDMsjv
9mLlJNO+TW5aBFY4QorNNSIAvd00B6w2GNreXr8KHY2nWTMydM+M8vEOmk/XbQLR
fmGrXkmA1UxnppxvYLbMexkCcaNRYSADYnVvyphzVwpkWnS+zWdRyH2XIEpVifyR
/UY4U1Byr+d0diXdHzxmPsUfxbbd9FVaU51bLpLgUFWD7P/tmXjtnVz+7t9Q8Cxs
2vLOwUvrX9KTqSgm0IQDICF5a9vBzxBBnAHsO5VBBN6+Pyo1EGmVutyXhegawinj
1DNdVoTW15upYa19Cd4V3I2oZuMpryEJ8vXhx/e1aJRO3v5+wUmt/Y2j2Bq9Dww6
8MtC4Hfyc5++roPtp9rdrH5IBMCvq0MonUZGQOWGQaXe0eMJkHe4acLKwI/EjQiO
avPhLKVtEkvypQxI8tXYIUFTnZPa773h2OZCF9bZPqGN05otGAte0MJDZwU6ofxs
BfSGMMYGrD5CEMcDdxdJJiKUoBSlr1kHkvVTj68EofrUk8nmlP8s4eWI2xV7NkQr
U0ZtidZiveL4RXG/NybMCsJlduA40qSCgk3Q4BggualmRszEKjQ+X8PuFmY8oQyX
yX0NS6+vMyMhaZjhFbfuKdnZ4Gz/XGFCDnqMKV39pf/9zYiPBizFFInuz0h8OHG2
nPE1qetHUDetuVokuIqP1Ovmhw48K82qw8rF5XWUmHb0uoqgBR0IWeAhtgSs5cdf
88YhNDs2Zi6jL+Bkp2716Ljtq22V4toF3deBwbhIQvZ4SKF0gs00QT+ejW7WL9Tb
OVWPaaMhmrvaPYKqmj+cA3pH4S73Y51YUjmMCmwwy2ozpRovP0IZlZsKDFiU58yD
dAjvo0qEq1mbQoZ4+2Rqwz31XKP2X2zR5J9MTbwsJcsz9pTv30WlEpzJ6gxV/Nqg
N+9S5+Xd7S/JUdfUe3hRSnK03Kpw9jaG32Ghz0RF6YHPC9DtVonTQFtbFyskBEwt
UqkG3M9aCR+f1YsBDB4I8va8BV4qHAP65eKQFdg/hiwvuEiz/nxG4vWEuxEZhYm3
71r9aHKxL6ilV19IjOBUSZZL16KIQD+gPW8Wtq/ocCECueqFxEyN3dz3R60N4mAI
yObcPK7StCzjo1+ssRMJ0en5/NRXlLR5IJ49Tye9slyBED+dBbZZegOWvuVVAaQC
1Zqjb/U9u+BXp1pMZdz4Vbvf6k7//QGn0VXbCq513iBJcLz9GQatS661HGApBIGY
UpjrLsOEbSr6qxSSi3HAL+Fot8V/0lhmYSsd1+lYaSOSfGRS8umio7PTZT4CzYYy
BtRpAzviND7uHgOcpe+GNVWVLYdl7+iDKLR7GzYQ5Iesl7loePfgXMaLCH4Y6vWc
eIeuRbdyJLmTms1yT1FleJ3rfli+wN4Vcmet9z1ABDYDeYVmdE+hN7c2dsL5mb59
5gYB8u9CVcSv+4AElATdqSUBHBfHbg6mrgKK9J6P2ItciWDL1zIX7TDVeMnySsUx
XrzUcz4lvlRVpkG6WlmykQNn5LFxsP7Yum4mSFJ7WpBm/9/CT+42w7iXCgVZVMGW
oDcFyUK7VojcQVp0RYUxnvj5gHAR1w+Th+Bj3XN89jgvCAXKiEKn361rTR/h3eZY
rVsOhz7ZLgID14vtNTowtWfAHt5Ceo6OZaxZ1dS8rFJcKzfg34JBeebUf6wlEWYn
1ULy67Lz7MLjJ+cCe7IQz7J6oVEtspATkZYbYKRx+3dq1149/NR56dTs24xqwipO
U5EWVzJkU+Gi5qUSGAFX8fS6O/DQU1BmNlwOW8tFDMLDN6oVB24Xs2ZZ5zy+aVCC
TXVHmwq1i5S6rdfCo6OyH5bpdgRCPgwSgOwr2F1X7E8WqNqmOqtMU90dn38cYam4
dtLzqjJvClJdrMxYHse3vnILS6ktpJ342kQJ19Xgyod0aKUZQ3/32SylByw9X3O8
Bitolwya/2MyjA5QcULUNBewye04vGQh5LvILQbIxvoFLZHbt/GzkevOu8JojAS5
iaqXCUHPfFM8tfNR/vAH58kz3SDTEb/E9aHB6xz0KFgstcuiBP2OEDL4f/c7Pnb6
NpNSVbjOjB6Csap+YidZCQdM/6gUYFKX05w0+6Qc7k6AAZpIGDukV6PeWYMVuNcp
l+9tCb3er6OQmERtMZxj22p1C48/tCpNX9bIG9QGoF9CTQE9wiMQDdgGkNfEwW5x
2U419FMlSPotSOReYM7iWuaTThW4b0+o9yLQgKWiWDJ6t0fpkAlmpSvZa2pI1PCi
sHk3QQp8KdqMM1fA4auXgJnzLQuPYxqDxIunZFWS1Atd4p1kWc50aBgWmAnIX/81
j/h5pF0lFyTdLr36Mw01LWzeHAWtEVk88SY2BkGOqxrMbtQzKoB2eMiKTfk4n1AP
uHkqzZ8rvuQgXPToS/LdsmjsniKnYZnDotYwiumFqzahbRhE6c0I6BH/+f9CVwB3
naUZAr4tYRyf92NFHNOQBD2J9IJqPi4wD46pB9vSwRLRYVpMVW3Oezqpa0op0m53
xHsjTyjXUutXGN3n17FFLKtaTVW2MiGexIxNgVSCq6TgcL/tXm1viBPE7yp0FEHM
FrrOn25pLYxIrnfOVmmh7anD70sATPznvlwYqaR+/t2K/jGQjrx4RVHKNGPPE0mY
bv3vDFPhYmTfUg26+GNSHz8TK+DVRsp+mHlsDnQBK62TbYjJW3AcnczSRL2DdG2S
C1bB8jJRyOsyk3s4EpJv+wEfLUfTH0MWeMflh1g1Nba4J9fDvD20kITHu5X9WpWB
y9p9JMxVE4dCaw7Adfuahye4WoGN9ULUNCOIE90YcMsUjHAQ4MoTAuSOwnafCo1+
pzdv0tvfrHR4S7H0Leh4kHpBSeMH8OliDt+0G0XjLfMiaiDx+cLQ1ktcryIhxfmc
kE2yaQ27nIyoIWiNRuScg0Ec0myXiuEgH1DYNbVNB4PiFCirmeXqP5J3UMgKhV1E
9JNRGoPkJf/W6NcLXz1TyIC7MdemUE6KVUE6LlSv7cHpOcu/j6FB2lqRrjcCbLuE
biyOsL3D8fRorINlg5JsYHD9A/hNp03GON/+B81c85BcRzrsy6sqJgNr+sSZUI+E
toDGoBd7Ikw3PPIAP2x3hvpihZs5Fg2jG28nGcdpAR0HfzTRc7jamPAXaDUm6zeD
U65U5+nH/xkHgj6MmLbcuLInHVVG8uiM5MPJA9aaK3bvaWOTmWTtyuGh0OF3s56j
SuuUTL4kHBE348mG8IqTNkMA5hajVKYdFn+RX7tVf7VBegC+ESV5SQV9z2Tu1OX9
logFLYe10oyELLAewVNhY/8aLfEHCUtiTGHVm2GrfDZCE8hKYl6QDCfGiPIZ7urv
0N8Z5++yQjxe2c703Z4HyqvEzLbXe1Q+5Rgd5G+xstkM80wTRinyHIY0J6BVOvxZ
JeCZu8ALzoxfakY6Q/aDyEh1dNfTsJyJa9tDqFulMC6XKSAKEHJOY9I8vOLxEeDw
dpdu2CpYkFT+jbTAjRWLMc8whqQFno1uxG917Z/XYsmz5/o8C8Jxq8R4OZN8kX3U
M6+4/+twSC83H0txBV5US0ai4FOGuMDw9Dodp+Ed/9uVrb3FvLWr6ut7HFnq/+8t
YTmi1DT4QnKjWhWTMOUoiX15LO+VbtKV8xphs3ZQxdSNWhhxMF+BjP0dB8LZX81m
wWIZ+Qc+rS6pafyg1t7pI5AgelzT7yRGkiKYZQ+3AeLacx9SJNmUTk4Xu/HnINrL
x00PcfSmBAMy5FFoyUbDyVAT+RVMylDQ0SF43/MYPm0m5eN6mea6AzyzCJdddqDh
cm5MVEe3seqFQFsSHQwfXR8SV4T8buSCmSGTeZYmbw2sWCHN55YrOJyow7bpLeZK
M6HLwTf2gjylGJEpCCgk3YXoUEaXOyG4HNpapkcZXlz+XtzHQ6yBhrK2LK1mIU3E
WoeWvRvYhIge560b0iLWC9PKL99KhJSmP8KS8o+f4EbThoEsYH73izoApI7h6Tzs
py+DxLlKQ1npOtlBTQHEm5dbCrv6090+SSWQxAyf1xAL5+kVpYyz2YSeG8H2PR5C
CxgJBy5wbesmzebauQ8njRqgna9E01KDEEgohn1y039WvfyxJDqKttz9+eMUOAP/
eIGqvAGt7wbJm/qx2y8Hjx5KciN9Lv1SqgacEmyWiArbRQ0eYd4xQaJ8cUx88sVQ
4Mgb2DzJVpprexgldyWO5yXT7m3cZanxNvoaUtgEnHVY0xyDHm+3XiB0dhKvc0ZC
4CWq9LokjF8CIvO9F/HMsK0umlyTcgeSzgwwZrXVvhGC9UWxLaBr2Xmzhyp54f56
q2gxXeo7xkW/cDjP963NuDfla4eEIo5g0/E/bqWdCl8c9FVEhw3UXaRFQS0dzSmY
E/9NE46UTwVu4BVvaoEPDDSwDQHXks8l1SLZogKvcPigJOPQJ0VdHjgXUDpKezZW
mOdxD9voU2SgbY+KEATp0MbDJMqAw3EHjtW6ksYdD0B8WWR8h7byHPLZBJZMDjXh
ihBpa9Orlvraka/tA0mj/52qog0TSrBeQFZ0/5S4qK6qcCfPASzn3WVzpYb7T4Jn
QvUZrJuTK2AHQoRL1M9zhQJ2ysr/WeILzkpL3sUcY3uo/4Gs/t1r6hIjJAe3dNoW
JZTIlUGOMoD/2JrUvobzbWg4S5HeSLmrWM20eJHOpjesezDbbKGijki1/yl1C468
MHlQQHYmQ7SUic5f+7bkElWMhwMQjrAWZXfNqQD6qj1o49NX7rc8ojAwWXOP/fRA
KNL5+apWJj/6OAfHd5vU6xGck6TpQCQsgGPdj4xaVsw2E1gBx9nPv23GIgwGVwrX
RCOTcbg8eqyLJq0cvuGrBu2GnUeript5KZxwdfXHQgoS55t7+jEpuW5KIGJg2r1m
KttJYq/wyVaW3nWff40jv/Bu6UaewjGvzcsr4JRUiHgBegsZiP2Ipl0peBf5ebFh
6WI5h6H8kiXkooUs4wqmpscBNNxJ99gX/Q0+FdKG1B1sgVYeXrLH8ZKl0LjBeekd
PNXrhIO3siN0uMpXK8oMLqHMIBMQRM1DBJ+eGweDyQg1viFO9SfIeVlj/brJZb/n
PVtBjCRxP9ac6UJbeW8yGuBCV6F1AkOC5sEll1/HUO7vNaq7yP8GE2xtQXeVw/Qm
5zDIeNqx62lR7ZKVR3fBB+GTq1d9mXC9p9pZ95hLZqzzHpLbf+fT1D+vMpK+1GUo
oSrAU985HgFNeIzOoBJKzsOWbMw3sb5JUo+mDN+vRWShNdVuhOfCH9AZMmYnINcY
AQHWZdXoglJ1CvnCvvA13GsKeGD7BEyTvi2QQAdiAbXaTVqW4cI32DhvPAIzh5oV
EvTohhc6S/Xelx6+EiK7+mOlUC2pw5/NuR/ZdTQe42LJvtmozEWBFASimAMi6Dfb
DzaUBJJde/Mx7E2oppKtfbppOcUzOlEOXc9Z+UNIHaeRDDVIqs7Ho23+Li9g8j3+
7kNx958cUrTosb3hxechFdiLYr6XoytLkn9z4CFYJmR6fVtMiHGtQavXRy8gxBq/
+TAz0tyEoDwwywCdSRjkQhvM/KqTCF8iN3Kxhrac7Xb1YbVLwky7csDbHP3ah5IZ
QAe1lEOigFYa5OurFZpWaZP4dzxNNeX0R7szkFymd8w1bDIfpg9p9GBUh2mC94hj
rFjb84ugJYvx0VPk6qDR3XCKMnEvshCvD0Xkmp5yC/N3gGi9YP5CUYsbdYMikSMx
+LDLfeXYpznFNaNqJGP/GTceZcyhUim2x/wL9ukV+ZCNI0hznvwo2kX1PTN5M+Fv
hH5+a4cS59y3IPoHDIU7cd0zXnuejFfjeqM7p2RCb9eaksJSpY9Q13RWzc/v2CtL
D7QXXt01YL2U2PyWWX2vKkAlZ+pujUamMAUFTg+95RDRkM6Xu78hEzSm2y/guFng
ycDzROT8LwrN2uGVA3jyPB+iD9Pvo60hUHjFBHWgLmujJwBzU16FdZPuZ06Lm70t
1GfRaxJbJt9UHPtGx+6wypAv/kcpX9Y4OCK0r2jnFNxV3m8A4ZfBB7n6r3hwyoyu
yuBYBaO/9VQYaMBpYwlfnwyM2sSpQkDu945ao/rQmJvYdWs1wbvv3Rh3s2o6XwhP
p2RMyTubLrPLfFZrb8z4eOrVM6+m0HESUquJ6liutD7xU+JRFcQGlbOTQP3N8Wih
mwiBXImCrO8RV378tEC1kVrk6gw9zLVKSZ8VV44TDytrzw4kRmXYIpdmJtkPAwpV
k3uWY8DBy8Zm8E7Vya2KjPZUR1VAKyaoAlMIwsLnnglJqcGopRHJC3Nj+WSC4rWi
cUj7KOA7USbe7gzsYst4bfUNKRIquVJ1e6ikKAeIj1CmWFt9sWzMSgLAiB6kzkVV
D3yGEfNs4xPF94drKgwrC9vy3y25ThVIQ5KptHtsh4fnu58rgR2GVJ7p1zmTSlUU
KtKMS/RnjjQx57caGj662iQ6T3lMB+ZLqMnTgps1rYO08PhTzYVwYn44GA1XmV8U
nuT7Nk5bngKpeXYAXbf0mVvPDUJQmM9kc04lm1q9W+Xo90oPVpGbHDWS7rOt+qxc
BIjNz5IV7Er+aSp64errxUaxAuGdRMu+itsgT2N+B+t2S7Z/oywabaE8HDXkz1GI
ioPFySzdvGO5S9TEtOoIwhb1xF0Vp7GrHvsnxr26llfKtlxIndrftlXiY4/ImUsg
WPN9cTE6H+wGxGat3enwdKfT8x976ztH9YXhe2tqGCpNehJ9p/MuWQrPplg5VdsM
t6G3yDgyiE9+uAzr/cJNIqKVhoC400N4ExhdIp3a8aOlOapzkFYNdzSqB1fPVTRN
CIZ5tPDRTgVeiDPrFqk7b/yePHuXrS0Bqf37lU8jdWyOi+4/Hw+xdAoi+zxwcfS4
CTlReNLvqjs86ll5AqRAIOBGKwpo8Pfc9eduJELVWvg3LfxmgCUuDVM85nAXG/Do
h7yCGI+hVf1UIu5JU3R+mTHKNXG4YjMFyk3XuY5B+uPFBNxmQOCTVIWHszQFHngl
4HPr3j4s+csi9aOs88fFo6G9+0nMvfIFipc31VL26KAW2YzNhvcS9yLcbbAFewK9
xHuqvgQ3eHXfrBkJYVtAlcUgCSyu6jdInxAb6vKSAPiDDG0IGkMfr5Si9hSeyFLV
yWvP8skfdPbyAuG3yMmZ6HK0uN1dMRktMXOnwJBtdHaAo34QwqiGYP2J1brEXkfZ
/WYPzi80x5lK5RmGzGMGWo+HXmnuqHp3trquxXvNWgShsBMtNENCimFUO3fjnKWS
BWVEeGczvimBw1MrAJy2n3SQRG0PMRJxAhqPi29QGVZrsD4vfCCEenQ1onm+5V3m
Jh+kr9XiDqXMz2EPIXh3oMiv2jUPR8bx25nJF8jAlaCTmUsQ32ydQeH7ixP849KT
7IGKyepVtP1SEUkVem9HQsMTW7OzWuUxY32K2wSYudHKj124k8XibLVTeKqBGtFo
WyS23I7VYnmzNZeYG/xoXqVb2o//hmFOJj9j3p2uOBUb+/D8Nnok/frbo+/VoKtK
lVl0I2r1p0CnTlAfkwGWRkpA1+tzkIre5apsvwfQqaqysaJeVe6z4kxd+XOBB54m
AqVyHxMv0nuohbVGj6lJC1aBXrdIijGGW+b4jewtamoRFQUsNFwodcoXYvQrVx7r
8tCjPQjzeFZK75lZioZYC1291cs+8dn4jR3OK37kSEH5qZOhG1XLSPYGQsQmJJei
RzYfvAyDpuWfr3Y5R/I3oaoEd5I7xIuJEaDWeUTrXLCTeuMPTF3hizYwVxliMh3P
uIUy3sriPOccwHEKalRLPeiGHOy+XAjJ6Vb8GcJDmjKLLvZiJxR03Hv/bmmBgguM
1p8mJdUWRot6F7av08i/7wPdg0aYMfe3r1Y5v5/wBZHe6/V0CiXJ5hCfX8NiScR9
b8fgMTye8fqh8Xm4Z2N4kzFeBwoIbEPhy2HOogcKqwWECI959JVQa3p3cEkg/zXZ
L8l7D7YAZdiRD+WrrK2Ea1K0JUrhg9mq1ljqqUcuVxxf7CjCF0ZGnzCX7Mwz4w2s
i5ox7zehgdYtQ+KDFkiZxAi30sIOTXpi09h/hXCnKCzy/Lq2sh+dXqgAacoeklX9
vmw26qQdWTg7pTk080NKkxtzax79qBEXrB/esO7qmS6wp6pU0pShYvm3zD0rRVuY
ryRsLpYzxe/KfOhMDgr2H25NcOb0rmWBuDHh0H89HhzH7Wt33a+xh/TqAJZfbm/5
WS501tbZfLC+GzUfKpQMHIzMiUCIQYHwJP/fP1O9km4TPzjouAsUHxv0AeMZ0kK3
+krV1431MpVIWPu7YO7xKdansfEKDjTgzPwvjxJimaV4FP6cJq8NWNEG6chqUx4x
9R/aykqSQ+57Khrisv1ifsZ0gj/PkaTe0JBhoO6yC+mAPESMMjWLszg3lGE1VDYw
vG5FUQyzAr8qyzYg8ruPMU25mGW9dFJzy7xLXMq7N1Nl08yvxESCDcfsNgEsDpr1
iUvYvZIloBVPvn9NtKMWeGoGKitf6KTXBQR5+RLbMTYpl6zSraQE0wPNb6a1cD+W
p3SN+BqvkS1RgvvgfIQ5zRTatjbfTKFvr2o4fMDcZk42VJtmPWNklI2Tbr+2HWxe
L+aXjSEN7MNagUV6qUyPR2z5j7kM5QIFBzXuK/s69sjdClC8oOTIDoVV2VONmBAc
oyV1LWvDQMcOd6WCN5ydbvwg9xZXktPefzNUqaAzYbGoXxTaR1926UJxf3NnS1jJ
w+qBKbl/aYctyGJ6zRc5mWeSaAsDphW7wzLKr6CTPG76nspWDi4Bn6aecPtwNHnR
5XQ1qo1nZR8ZkgCN1qYDX2gz/umuVN69u/Ub2/PvZ2b/9mZLHhdrkRc7/FbNlZ9k
kO9YLOVlDfZ4bd9ozG62Cv61YiGt83dZWtr59C+V9uF0DScVIMN83GNu2lFzWJV5
M0H/Y0IvArZj9QjAe5QSNv2pSKtJKmi0O1SsZSGZM2ZfnOxdJmby1vbGjn6h+hHr
7SzzxlJKVLRqQ50B2SkSnZpD+qzAauPAjAugHWShMP5k8Cqv3Eu389QJ6Y+n6zyR
LbC6OIMQ0TTOT/IS8OWADRXgj3lrHsNrfpiwt5T3kBDrDQE5nd4F32/mXVKGIkPL
3wQXxQ4DEpMmnLEYAKJR4aPS6iaZJbSGpg51//Vp5Kb1AAsuZPl5Y1bRGYahb6/F
4A/aBrJO810XtD6Dczvygv3J6j18vIym7FR/3WJQVJZ4IwG8WJij3C8h4X+kKBFq
QFLKr+avFDm7sA1z5Cvlr4I4HIEZ7VqlzTi/Htk4o9w1WHOPpCxbOPCld3mwyF9z
V8QMZvShqvtpK5LfmS014gWYbEjp7NA5VLahdaVASbdo6dFJOuhpp5ALn7Bb6mOV
NL3JXmzwcoyoh6g++ccBk1AGhqtNJNGGoIswIMiF4wEDvPjkQTaC1FBkm4ohQtjZ
TXk9J3yiGZbgPBwtsJozMj7zpDEdjevouBpZlk0lyPbH4NcoqqvYlrH3gPyvPpvV
2rsBw6h9VEhXA8LGFzMkmKqNYLz2JmYRG/KHA0ZfAnFl10mI+bZTjerSjB+Wwn0/
Prs0oW1WwQmbmGp5vknUW07K/zomAHT1npSCJvKUe/HspTMdm6tPY7T9oSrGEZx3
XEZnjIH6Eg0QVWtWjO+46k66Gd0lrr+7yMQFwaTsNnznZy9uQWRtXR4fwR8ZKPU4
ZJAwosdMPToBopMt9CXahUs8XtDPseJctpYWX5b36NT5SZcRdW1sIAFAv/2+fJ2/
Ze1mhg/vAuFisRojNZPNfnzPngPPZ2Y07HKLc1eq/eZLQdglS0u+7Q5wHQImK5kN
7uImKYRIFOO6mNvTbHKIZdLGPsNZhb5clttEd0+tR4ik6WxKJpNq4Ds2tDR6HQLj
vGhyI9VmSJ355sWBNNx0GF15gb2ifalbMxDBWfjScsAF3tbLi0YTu2EHEU9D2gL5
gbUtsMoYb3HCMm46ZvheJrImbUwBMZBIi/qtMCstbyeDyYcLCENBBwoc3KWHNZHn
W7ujkFj7PTrZNqklaOHqLw1FFDeGiDeP8bYEAKz4tzdD8ubV2H5v1F6iJnGVDqmt
QKb7kGRGOD5iRu8TxuylSBKNEXwZPuu8EziPED8VZR2mjoUtNksisgv5qoNaJ6gp
rghkEN9SpzykHPYMgqzj0EBBikDiPJfN7GuoAsuQcYEpL1EEKTmBFPZuDXTGA5y2
IgJah/XyCUZc4ZXQt/iLfP8Vvlz1kONd+utgnDUPsxO0aKWirGUnTX0K7V4QJiiT
FiGCsUl6sG4Qubkd1v+5LqNHhJTs3/QEa7Gy1F87rB0pE5ADTAFdw9VA5gvGBsDJ
izVXDqUTiD2HPMvc0idRJx3seOswRdqq2SLpF/cgSQIkP1ZUF257RjejRpVgepAY
go9qas/gdoRZUIqg+BXMylaF/LfpbeSkQ/4ENqKHUUN7ieXG+YbZrjdsLqRmB3Ms
3w9L122f98SYwcHjxZTA30WJttctXiWcOJlEmi7+w1c7a+gPYbrX811dcYeFojdB
/ZSohqP3ncMsSUGr2lQk4VoQHkJEPPfP7ONa5LDg1pLKhM0FB1I4LKcmgyHuAmqS
ie/eTU4hFxe/HRWnEKcoM4VpX/HBq6QzBGoJYZY0sQxtav0LkEL/XJKoARWuaXZE
2WKmQLybkr9mjXmivzIEopYQg/xzlp6RW9uGkH0WN//zXzcMT0xAuN2URQpbupPV
n+dqKEoptTTojW/OaAYC3NUeRHgPJcZNiptEoIY+UBnGX6x7v7VyvdYbQTAUI9SF
L7Xi/pj2PC3jx/Vq/i0ZQdXh+klpWAmWe2y8NTjxgrGqETpFLqzE09eKRSHzQh2Y
kGDOC3Qy2LxeLquiUPJyQVSvlUNd5xAk/UEugks3rIY7e2c1dBvkZp9YpDUVm0qe
HXMxRuuTGKWjq+1AIlSkRJA7aoFL5gOa97/Bu1oIYInpFKXCrNcqaLH11UAQXnKr
WBTVXEPjEhedKKMbtWYuaWDLLh6voOJzlMFM0SX2epDYZDKfNXaWwzFIe9cYoUzr
k12SIODlLJopoG4zBoVGwf/ZYxhtegL8uHBSmxpD2NS14SCmH6IUWCxgnwumMFna
jK3xu7V17SDMzAPyw3mmxS7Q/y2qguPhQd3ugYh+vhmPobtdMU7qy6zdt8kfgxn+
8jJycAxpxCl2yyteCDRsJKKOsCQSuPQnzFU+TY3jHemlRI9YWL4VXXPfiRJ9sI39
zpyulj45ZbiAtEOaHJjcrmz72iwu2iSyKux35Mjdsr+utA6xndQJQPs+wDaFOjOW
5aQQrFtuqAZ/jI9/lmdVrD3ABsWaVARjrBsg4Zr/3Rrqtd2T9pHwlcGHuJAfyn6k
BTnQRxkR/6huCoaoxrUQafBMnplGvV7+5S4MtEF3X0UbskVcxe6YFSf8VVVD0N70
BfAXcxs6Ijq1lG2QEFljBdEsXok1h6hLU/T7jUqYAK2DN71nLnovWC0KI6bGkQS0
YMGf4n/SZHcabPWyLur4L5IGUrRjARruwC+7Q65M+IsBaWFHkUga4JC50ZVJ02MV
7HFxqKBrikXEW7myebwL74XstocW69iRYjfuv3+wGRJwR+flhSonC0eFl1L4kwcH
ELQ5Y3HKb1tQVnLJRbzaJD2nbdyFXx37KzJK7wmCa6/pMDLFxLT7gbaxxQyyg+Tr
7mgzIc4WOotkyuwJ+lWY1Y1N4J8OpqHNthn2mWVZ9sq54tXZ1p29d/hfmv14HTq1
3utY9nmbU+H8JsZ1CE9b1HjZkkDsrUlC+jJrlpYySPImruK3iw2q2s0I69RuQt2Z
cTTn7jzDxxPncAkoIlpLKgZejnRwr0wzReZu5Q//FSGShLGZnzyzE02pQ/buJn2L
1ZC3Tu+c2mdqI21F3spEHT6NrP4DFHiheSss4uoFEiSiQwH025ixHiAD7kX0E1zi
Ml1LMPP5cP1A0Owcl/+PUY5bBNcR0htJJ9vqUdNYSZvye6O9xiPGRcJjQq8qAyXw
ZU1h0eB8VjvdzPnKviOGKxdnVAm5VrI/7lNGYyaTs9YUOT8Hke13pkRM+nDdaBFS
tBwHxLsPAdhiYv7mdj5qNE45+n7tWCbfSetiUGjzfXFlhcq1uN7bpdEO+93q4F2q
JBQMnP92enSMG3SE3DZafIdrFooPWrzCEBsVFnUsNKSwrJ6kNjQi5/CSVdGIm6rG
etDIf2tn+lL0XferhSJKMsTcmRJpJSc3i7QZhUYpeNLS8GRL6AobkC63Q+8Hh5yY
abvyOSXcTN+vmng3RPDlrUjhL2EPHjHgOriDev9ACSRBTuDKGES3St/DuosC6GPO
bftHlDZVmlP6nTPaVNZ/RlpCBckWTVup/oYutJWaLve5fb6uuKpK/ePwEOpf3id1
goVnUucudBF2zKVshvyN33lSFju1VEFohabRg8J191BO2csK8wzekwoQwRp0anDt
3/DtLiTDKAMtaomujWVJyZ12MGTgrKSbACj9FUMyeR266wV11809+ONqoE+XQ9rs
S956R3hYhmv31d4OqzohkronPEZEzYuvVbLZKx6Fz4rbK5CNy7Gt4wtZXxWI1xCS
AJ9QYA92uSpjUhYi56vKs74WtisiE8L8XyzLP91T0UXqte/I0ieY8W7qEgJ/vBaE
U8JxUm+Wa27i9bLmQ0JiMHSQYh/9mg5BfoVPrXtZldHVcxlAzPi2G79VTPPQwLNH
T2J82oLa5NUu47IgZJLlxDh1a/teI++peFqGo7qu2YGo3V0PfCIxEEpLX/IIk905
MG1b81A2hpOIT8b9rVUdIsAZchQrSW4FWUCMNjJL1CMtz7lwwi2vEz7UHhZRfiO6
Az7cerFUFnJipgAh1OjUeVVN1KUzPV1L+sSaB83TS7Dfzge+r3hlHqdZ/9okfyuC
V41EO6CrgK/ActsQM1STIEvvIx8Nx3/+EUUNlYnaGamw8XiXqgc3q4PSsTcXPuzO
8iskOoHd1a1uCtxz/BnQgVlVhT+NA+JbkaVjt7/kiZcFwt+zTyagxib4i8phmW9g
mw3SPGLr/KS9BE7/O8fSTWIrLObcmf3Et1jhx/UMEH2uPEmaCvgp2pd81smXyh6S
vs1wqq90qsV9LD3Td64g27d4hONDbOxRoozUhcCLMAfcZNl+E2xmYHXISCqx5L2D
PMPS2Tx57FiJwrALaotDCG+bO5KVfJXR8qHTQORalx83rnC2uZfI734dQnKlDnUh
VEsJD7HwAifHfzGeFg1dCOYGfpPbfrhMk3xeJoIZ/0P7CoeKb6FsxwgfaIclZ2xb
ukzlAveUgvG7CNildAHnEKecrLbvNLFAD840qx1yYBobE1kopSrsLld+gb01+7Im
gCeLGa0sAVfiZPS6r6ktt7tLAXgn1IK3yMOR+kUFD/RdY1MWv3X5llH0+OqUuwJi
oVF43X2N/10hYQRdG08mA4VkP01hETjBkzH/T9Tz/ofIHPZcbdMZg8YqiplgzJuo
4ZoOmIOKqwYQWPD3MmSZrByJn0KpAQdVyO+xSdD/R9EoOWhDi6PxJ6IfxK2Rp8YF
36icfB27KqZ5sHIC+ZjiHwnhi1TrUSI4hjlVeP3jDnVpsGeZL27/daXEamRbxJhA
p2qY5LzSHLMxDuLfK9CSbDpcSLsdtIahILbJ5lEMD6MG633/4YAMW+6ZEYEX59Fk
JB95T4EHUZ80mJXIKNQuXQFR+WfelUKHMTZvw7ZpmNRNujvwhpxw7wTnDRe1Ws/x
zBaJvFFU1HuYaXlzc+8hrdVa5Rr/LQEYBVUNH8/GA2pEvay3pHvxXCsDvg9NyNuV
YM1WWR+aoUdBl7uoWAihD2jpNMUaPZJMroFGFE46d1CrXdl28fMRazMS9GMmXwtY
bjktEtmwVw0n1mTH99CXfZed0EoccxfT2Pk8Kk+9luq2H01GZT7fpi5Zm68DmM2m
3o2Y+Q9wpE216f+u5SFpJfzu0CmpEmr8XDAITQFvpdT/WLnnFnFkxez657IW/ZKJ
lEPZ9VL728cPShtBrERH4AlGOVvArotCFXEp2LMyVii0F9zfzLolJvd4HcibcGj+
UkY0SqCKBF8Tov3t4RtICLQMgnzrjYX0+ecKuXvyA3vTt5nmOwoywdFFKm/6BmIB
mppqwsWdhr75jnJznbf5FZ2ULZtUIRGJED52VGUFMuv9p60z3/l2iyq+81+BcRl/
uCEIrHlzDzNq9WPHq6WIxmtUt2KXy9nyflkDPhnituXpaxmK1/W+jt/HkYa0IwCi
IIXoGJ5it7Ob+PltocRUbGQ0K4NLTepIhChiUJl59h3IuQQaF8Q/IlFcV5Ombqn3
PvE4nxy7uxuGnqDopk0g9XXYT3U8I9NP4WR3VA5thUH8YXvjReZBWld2dytbjhzC
6JxCH674WK7GSEL+kQ8bcaeuFGnWPcp3myi/Vwml1n+cqwwaT39vOZUnRkZspIdC
H+mcYCNgBBYnkpVI7EFtc/Ks5qZDk4cCdMBhr/g1SBXgDKNpMvUoVwE60QkgZBRx
nvG2C+FBVK5UxildWBxE1gyyIOPq+ylS4hTS8qc0KXZKBvIbtAbeFW7BI693iM6M
CjPwoGwRfzEhvl+eoBQ/UyrRgelqHfalVkHUy8+ghWj7goDpfHe7rtPy7Tq2g2M5
ISexQwav80ZlSm6it1Bk3aJ2zYwTSr5PJtnI8DM/v0gO8xtcQZF/OG5AOO0HoBhL
vhLuwTdPmkLlJSF6OKhM25K2RG1yheCPCBz9ohb6RzBg5Lwc+SdsdW1NyA67K1KQ
1oEdl2I/siDbgw1neis0CRdXvG2CTvhAECXzfgeQTFZn/ttczHEygkuOG9ukCyEp
4hwBrp2MsHkjEUBATPE3YuxB7/dgYz3cyBMcw0SgTL+zIRqYFnKDCnL7XUdQ3EJg
oz2AmYzLuF09zlCavZbh0E9ON8RiJxzprx+NiragF0SMc4IFhE1ZXT08HkALjwLo
++a3Qnbsfurkp3KGjF0udO6JKBqLRw4T2f3RxxSodW7WZymTs1V0SeCCxtTzpP19
dLwbqi94Tu6obJsaRLoASpG2uFbUhZ248nrkzUPQMpRitF/TSu4d0lvrh0JS3vrt
M6y/1Gtk2psZ8TFMgJnSqT6/pNQdHU00GXEBA0GuZ6Wkbr4cy6vvsJVM0oe6kikD
cUZOeb9lSfIFYpvqNL82OnEbB9J9dyJrB85dLYyoqOXJ4hENxR7LRKII6u/Cc5Cy
/da1toJ0i69aXn7JUT0P+iInEZZEkaLCB9IAeuUBFeAeTntt3kDVDOEVrpWNXIC2
i9DaNL4txfs8XLj++OCrTjgJqDa+orb4iut3NioILBuK5q7tLQXgmPmbQPUgkvq0
CDAldBDAZOHDfPzu92cJ+NdViRjtzUNgz8TZQ1g/qfpa2WyiiYv2C3YtUZLGj9HH
O8us7heAZxQAqG+q5gjkRhvNKdUoN7B/6ah7N7wEZms6KwQVaZ0QCPWX/ufbHCB4
ozaC0L/kQM8X4gnjZPTS7EgbxmXdDO3oW9bspNN6N6x4drmpV/GbQ29zpEhVeFXh
h+fXxXEXKC4GrZq3ERYecFLRzWWD5dWfXiwzWmfwJB59Z7yxpkKwLPuoa/hKu814
Nu8PJOInVl5FrJNQk+sKRj/sD66UO772jerW45leUQ7fnmOIrx5peYQS+9bwE3Pl
qcPCRLP1Gt997e+YXQW1LerIl1wCxxZA9Hl7ZRnN9RmPLvkGq1nfuEPpCnAcJyrw
zpeaPWtI002dE8MWE3keoW7Uegvs57s4uSgcTlQWRwPBdVCkNBSd6kMrh8zsII5c
mNdmn8m7ovEHRaM1Ib1FmyjWyHVFQiR2raUHOExLuvV+RjbQOT24g2RtsNXBRPrs
DjxXNfQnFGlX1HIDTEQMNTipZMlaisWgDpvUtGqdkPBl6OSPhspIFqBvGiaf7OCV
upvJovFxgdg5Y0rhIvCa1Wj5KP5O476HNqw6KQYUwqNdg7jPxrjKBF4/DMJ/7T5T
v56xk7V3Yb5iqn21/+6GCd7EDvBjZ33dUK3M6fLD89hhw9Xdghd+CIFHUlIbcMiA
60CXu8nkjgdYpzSlPXPHY+jP+JKqnHH/SqcXk9TQbOth2AUCqsWcMwZrBaWsI6M1
AtbQi0weVYptdJSINNo6zHsv2VUIY70MhdFnDPZUXbVDKMJeC6GjYMSbSFtLOEpR
OQViSdOrmg8XSFPhjnYh3XjwDG77b053dpiSqdMQZ+V2iHX7jenzEQJrx5Ixggj9
VvnpCJpc+hP6OBSLIj+2ux9TBMPbhdzn2BVbaKyWosAF1uBOqzwey8MTNe0ATsp8
a69Jk7U4XVz+1xq5G6iaWburJOyZSta18lrnvisoFHQrBzJR/3cnWO/ye4g8MlGJ
pRNQCWwAx9fsEBW25PXARcqzU5qDjqtvsKE91dS7+LfDJM7A6BW57Z4aBv9Tsehv
HZiEG8SvGsiY9zLghRgGo7/I4KFRowcFGy5pOP7YBy406XFRBhLn6dj6xNE4HJOk
AGP+P0iX2TjPib/6FtciUMYA1fhTrTSo2cujNmm5+5lsmiIhNsUYou1DrSWrjMvH
SYD3I/d7Wto2FOwiVIOwAjjzaTerx6fgAN751WUEGS2TDvcbz+0qiV3CpGMA0fvx
fOnzFzHPEnG1W1Fc+P8+bCpL2WnmtayTCfGivPtspp3mpMQiv3rSmIJMEwmAGH03
FHH9YLQlrZIWkcmThCu9wrE4dQc3c4jJLAkcdI22kRQN9cMkMU+TNm6b2LZYrM5F
UyIAK04IhbbugAX2L8uS7e5B2A8XKluJGjrHVQJT+uoVmDA24/MLTfSbYCAtsYha
3zQh9Ysn1FciQxpNEBplqjy9MzG9HhLK/eO1FOr7+66d1zKJzcq75Xt8+bQq6d78
Z5hDx9NoCtgycQh9KscFHml3riPYFKY+5duHQb5gIBNdWXkcmp5iMB3hZ3Q9Q4uP
vrB+Y0kkQkMRS3Zq+CZKU5anUeb7nQ5FfNmnUtgzGQFpr/5F2P+bYbn+XNk9PpVL
dQ2WFCRICreUHlqZB9bBaKwo6FxsRUP00/wB4WShohH5fz4rJ0wiy1qonxMzgRlR
GmS8npfnU5F6fOsxS8hSoejjR1ces0wrDpVIrQsB62Su2HxRzWABG1jUyCohT5ys
aWSmtgtMP5gx0y4p5MCmLrm1WY7gvghZxUGYTmh0BqCeVBBc1p0BOt9EMiPgLeNN
vlBkImSJIJUeBVDlRcGniL2qPIBMsBGqa1s+pPq6Vt32v5WF4ijZdFm3jmJRXznk
kbDvDLTaj1h9hF9BxycpYWSif0trmXZwr3h9Hv2FlNnYHNgc51pwDRFVbKQIp/XC
JD5IMhaWD9M9NOzN+lE2zUN+KexnCuBtestSaU73cxtB3Aix1DMeOL+DUVLgFPKK
qCMlFQMQ5FLY9oIAYwh9GD3SOfbYrMcEzf4Qr+qsFsSSTOxtvX2sWOP6bmdBC+4i
hL/bJDdu0mSlxsrxgqYS8y9QB0LMixC8yceWI7TeuoLqzLy8etwxoNRThP8KhdX7
77iVgNOIVuCVcs5TZWeWKP1pmHSTWLVy23RP6jMckvnWfN3rD1BckyDYr9dABuzc
4AICVyxvLzEpFxe15p/MfqiaUYc1O8542Kjuz5HtIGdybEaKQkEiJXSMjRK7XKsH
tebvbCatKw/XeNdvqJfXeyb/K0qenAJNBertfaCFgor2UbxhwkUPOj9pj4ZgcjtQ
QgOidRbTQwGgYCCweXbvSBeUUq14zToRGtLje27L4QYyrK8jn0pzukfVZCjjceSV
pm7QkS2Z0oBMM8MpN6JgQb/IzdfJnjJmCw5/grPpHNoBx+WqoTl7vKjV4nFX5yzl
iGxbk5oBmgsHIhuh9YNb9IAMEspYnxZqKDKndJekRWGAR/r40tWUbjz0Kd8lQAZv
RfuOiW0Ad8sBjshixlu7gSB+ERKcnxh6zjETWpSkpm/kmYxP5J24FDG2OudLPi4A
ZLJ1F3MSeQKs8huviPrHh/j6z2fSxdIdeb9T7RNwLEIgETX4LyYA9dA4JBEZ5Aqn
xLW2kylCOKyCOGmc9rRS2VXOKh+7Y+pC+vnBvq20uyNWIPHDzPlyNqJXAHBDxXtO
/8J7ulh8V1fAt5x2XEgnY2auGZLu7ovQxeq7ZdMQhQKKtSGNMfP5xTgtB7yGYq3E
1QtI0gPGlvYzsCkm1z+sxzTl9mUiz1ENlULBMujqzVvlK0FloM8mZU3Z2B41H0fw
Hx9R0sol9RaBuxJt20P+ngFwvuGCiwZf1GA1YJvf5Lue/1FEg4QcvZ+njcH+1t5e
ntJvgT2isPQUUPfU2putyjMx/luB/C1I2muaOm62Cd70S8/0mPq/rAUGnQqVf3zc
WgWSb4VJJ+s6EKIYctbUnnrR30UNkrGQ5XoGlaur+k4Dz1D/+c3NIkSIaKYXHOUR
k6+OVByoROR85QhS3XHw5lf8ebwze3Sqz0chqx01iwuVdmkgaw65pm1piAA/W8Rc
1rRNyqzZOp377pB61rluMP3yd9fooZk3InyDLCVkcihuugy7fLKS0B7slmNzkRxn
pweswmfISnRbocphxuZB/0LWXSWRwS9ag6pK/g7gwses1FNdhWy2VlB9WzkHLrGR
Am9pyJKa4jRFd7EgfW3ujcnO90ITBiEh9DDs+JigbRyjhZy8nMLm5oxjZWDItM+T
stjc3UCgc11NS2OIUF3dgUjHSk9N4Px7fVgPTUDibrvQBQvD4udWfxT0G04kK9qH
Nrmo5TByfzkCoxFUQ3ShWImagn/IOMXpv61jStexmpgmraR7tcI4+Ppr9RsyTOKU
RLURxRwpHpHa3GuJV3trPEvoXtc2jCONlTgi0eFRTd85zy8LBH9jfhZD+jZIU52s
3WAQhTbSHGsG9N/arJo2DbOfxjQKlhJlGlqCzQtTkRHiEsn5535bvjhkkMasti7e
wR0CLkDV6L++sp0F44U105M6ti0EVdhg0ZfwOkKMZNQQ9rZGsEB81tHBbILRgfJo
iwsLm95FQ6ldLN0uC3tcnfD/KIKTfFSU4wLrunDvcmKdYvz4PJiU0euHEq0GHcMz
3PAZY8AkneZBpIrMA5kdf5VGJVQe2KP8Sexi3TJ9Ejlv0/Dfp+t6/yy/n61dyl1y
syI+pIFd0iFXlZDo/XC9fCntAYGmR0ocLDZE4fDe2DaXtWHrIVFCiP6FostyJLba
G8i+EIajiti+CySdpSuyeRHhC4qhJElkR1EC1tXhkik7n7JJhVwhHfX0mwyMUnZ4
sjtgpnZHc6i/s/e+HFsXfiMXm3b85kbHbgZ16pgPo8MAWj01CUIcaouUfyosvRPV
5yDhHOHy75tKu1h/3bgRBNqSPszlsFGpBQJBonY0mHomCz7JOqxOCb2XeXSpVuXo
z6o39wrnoxtPVKxl5VR/DC14xf9WLIE4GnLZdGoOuGsqZw6IHNl0Ap/fx5ThTxZI
MqPOrOe8LHnN2QQhaaJHgAJaPyIUlQEslEro6kSXwWnw/GPrgCrZqRJq4xlmOjJn
nnKGAK/jPGwR1rxMklkawPqx/9cCwnugQKC3Fx2n0qL+nPpmxpoEQS/n5fFyAvSI
Rwc4jokDgvEwteRMsl2DyptbD0p24H+EvnFShAPxd/B/COLKYgJJpWY/3M0jsKyr
j9pxpoF6gU0kl5MqpuotJ+rZ2Wy+KILOxC69Y027dvgzQr85bwTXNCxa2EmddX2Q
h5fnhGkuPezON/DojcmSJ8lEmdsh3rcv9zL9VmumV2tmD4nr6pgAH6BbLCkeoioo
4q+MXz1qqJpsf7dH531Qv57bR9QdpNajV9LmuHOtApJwi7jCmKy+fnzuu8W9p5Bj
jcw8QzCWr6fklP2p3389qxJJVt7AHNxMSNG6ZfbiLf4tJdVw4c9pkBbpR+L+HGv4
jt99qYoIn5tsUSBwIwE/5CI6MCdTWyuSFZw//vCImc0ZlkYNqFNSCOiO08+35T8O
WN274HVIglPEEmoX27bdJLAEdUDvYE4qrk2JHVFkTD2D9QP4JAqiirZhTJykumeY
XMvLME61/Fok0K3Ldobbe9aS4yxNnEA3D3xyi8uvEqcYJcVCgI0QbXdrSE/P6kfF
IwsKlPbffslsvw1Wwa4qW1v1ioIU6asxUpzlR2Y+QawE+3z8N1/sBIFJ7aB6Y+0D
at26SIhaZRSQj/uEGt+qzSq+wSoLH9AmSiVWNSJprMKTpIQDqslg2lTHudSPiu7H
RdRqDv00V4Wx2njbgsKCJQ4WKIzK+74myeyX8rsi8dYfx+uMRgGtjr0HjHredfiy
mEfZJ77NDukmi0tDa1hJ/uVxIA9BWWc3fS8f2mY8HZvrKWdkGIFaUaJ0DqxtttpN
HQru4DflNHUJ0fWM+20vSg4x87ZZa0JCrqNWmkjDUefOCGNPtWFbyYpnpZyFWUpZ
m3l3uklM3jV0mwm/I4TN2IOkXNNtOnEYVaQeKf5FIBtiIGgI5PWblO93FfnGL5Bv
IFRd6bQ0pf5q+f1E3t8kVgquMg2Xgfm45o4yQEbv31VxXxwJDcJp6CB+fprZw6Zk
4OHOueeQDhXwt9o3xgwZe/cUnm0mzV7h7mW2glOl+OgOCU7PMcEr+n/hiocOavYR
lZMaxbTZJf1CPgxEwW2ASTvfLNEIX/FxJaWSZTmkwIrRXxd9yKUyJvXQHGiA31cI
rKVncvSmr/BXmOT0qR0JOrIr7IQiLykpYpBMZAiyHtGZHIuSpfYA8PzjKn4ZT7aV
iR9jl8tEWCcETfUeXhuqyTPts1NaJGiMC5/GoxAiP+CDHUcSEMMXE51hqNJwaTeK
AS9bjiynhiXNZbF2H5aXKsE9WVtL9Zbl9r4ZZQ/dIyRc4hD7uikOo23V2TVKF+fY
WUAxaOg0BJepwmF3e05Ev73MIs4MJgTD1PbqtuwFxAIB1P8f5SZMPoicjbN6eOzm
94c52WBvnhaL2dv8ZVDJ6av/2L8Vt1vTkSq9ByQKZ6hQZ43Vn5aaZ0C63GjnpWxm
K4Uf1Fexd0t3fGP5oD2MWRiU77fn7MrtO/9LF6QW17ikbn151aNSYoDncTDgrhFf
N2ZbgMQBxRPdaZmP/Ke6siCmM9tb7iWG02NV4x7DV2Wc9lLwLWDfE14HmMjOpcTf
AZAu6CHgQkusKQXcRFVNvUQJYIgmRe1ScIGjVjNbT+2cowqcuFPZ1SY6Aq5TAyFO
iu4cgvylvViqcBxSgYBvaVqkm3cbzxsdVZb10N0v7aW48/FzlqoGwP7TxumC9GQD
8QPuUVFDttxvzXeNClOB7/PqAvaOlryo+C2RPcsW8eKGRNEh1DTTesrA8+EGpJNM
oJufYGGLqkCfQgxpHBHEAR8zMGZ3J0F4F82+hP9/6vtEYXevYVdwG6Nb73AaYaOF
u1uWTK3c3R4xlv5N8DZpCRREAf72kbM71fWYDBxLEcE+/BTyzwyywf4DYScM/+AL
wM30KrLcAaN5gIvsrIjf2EBDQxQmmMsduVmp/XOQmUv2Wkj2/M3cWMVC73RZJkGX
fLQkxQTLUGaR/Tknv6y5u3C1n9GR3f9bWM2oPHBq3PTHQYTchCD/LAcTPX4f4AXX
OD9mvBQWbfsKKSOWmDm0HjyE72ij8q1RDlxfoTdEwQTzWTAbKsDHi+YNAT5qHeMO
j4afPKEq4amtTU9n+S7krwwBshn/uWWdia/fe+5f19rtySaMTx96sxw65WmAU5cC
bq7L/npWkFcHUqep/yNaXqf5e8y9ymM5aKFfvR02XpSdR3K6G2/uIeVy7XOVhb59
gZfU877hMiPYU60L60C25NMJoNHoIulfP0d3fycZUpZTD+Z0Ws1mLo+U3UdtY1z1
QsbeLZ2yV1kc8f8yXKMnkTvAmMlQFGxSQmsEfNQ73UXm3ivPADUCSMgqCsKkFp4d
HjhtrzEaVsYnUyBeXuQccP3dCyn0nLoFlLLx7KV28oDLgQk3LKrwnO2Yx0aI5d8Z
C/3Gxc5/VQeS5MEF14chfQg+FUYQz2Vj28YPqcF2Sf1imrkLujZfN6zijqFFc8V7
mjHpAeWJ8oJaQOZfdOmhwlrVjmzr2mVDfqczx9P+kj0Axy/TDlNOC5UmXAtbR8XN
irgjmcR1zLDpK3CR7yZwaal3GzlDYlOjPTmjhXXDiTw+LVTdpiz2gdEPZl5XlASl
bVrWuYog+3qY8S2thHx+uW+f6vzqa0ykE8WHUqJTWEm5TtNx+OsRhAU3XeJvDctS
56I5TdEkeEf7MGS1SK/Lj0AM/TBPL3m9yFjHD4t2+0c0ItJVJif92L7JrEaW1vFc
DRv1pm9UT2vV8osk9TNUsbkMjY/RgQfyXZF1fm5LbNOUGo/HAysbM5BqBHP3hGgt
MaqGQj/V8rpUlQJ9Pz6eNHZtabCGv8qdKN6xaHKtwoW+EPP5k6HN1J5ztBvXrf0q
RErG+oo53JD1f0kKbcQ+B5zq9wjdMi9fQKuJpndGhAWkGNzZsAlX/6usVHqQvVcv
i7ej7SHvD+2clf8CZrMNBkg0UDmqUa5iUR5udcHM4V3Yyxa4DdINgnAN3AF+gi/c
+q1vblLRdL2PvbESwykqHKk30JNRB3n83cyTGHUrF3zfpt3L3MVG/aIWQT3Lh0ZR
fHUctnvuPlzZVVGPrqFlgBMDxfsxi21WiyKYs9jIB1z4Hh8aEZPzvvyxqOcEmlpn
eFPhTLZEDPesJirMJeIsm2gLTqDfOLJzJVW12sNyXgV6EMaLNMNado66AOVrDNKD
ndHr0VHA+hd79ZVq64cEZ7EQkq+krDg6A56wUiB2BAq8J3ZATlBR55fRNaEFgisN
4b4eXph19MHgN4mb7/B9Z6h1cScM/Hn20dcdKspkHjMv5GU7/iXFgtozB3UkTVl7
3xXzrOFM4rpOBenFTnkjiaDTSSefn89ByrLS5zDCsnPkwFHcoxcF56CpQJMkBwYZ
7qxKfijFwnJVXJbxbrUuMTjJdNjTfMvxnaI6QoKSESgl0pNABHOXgT0OHG4ZHyLu
EfwycLGwT3o8+g6YRsI7ofs32iBShli+siC3yaF/D0WJcF9HJrofT6G7KfSZ616j
NMJEi9rZHHG9f5UYTekGZxJDF77aK7WlYgWc0NBwHBEWbOA2ouvkPPVfSDSZymiq
iQCIeLpmK78xFc1MTPdJdFX6oPmqzrunjdv3+qiWM0A3F4CcCvmytg+6Qkv8SIZ1
82koKvRSQ196pC+GxlYgT1FQNJwfVVUFnk935xrftsK81baXUh/TDNGA7HBb05mk
ZyUr7sV51qkZehnVJs5j0gIPMHPLxQzvwr2NGrCcUY2gLJ4J4UPM7tHszzLYYPdw
Sp5qN177yOujlRXDin7aUxGHZQzjUoQi26VtwUjNwn4Fl5vpT6rJKHLsiSscR6mw
woRsnQ7k9LN+gWoSPyBkWx851DQTBLMUb+DThKBYEhBbjXVedKr1mHiWqjhwfysr
JGULJOEfqMoIbYIFf0JY2UgRBFEK1ia0umXtcw5w3ug2ZKoLT5b2JeEGSPm4tFzF
WBCKMmyRv1AaKS1+9bGLPG4oZxaiYwCc0ciItA5qYnqinxc0yf7eIyuNPXPgKTCv
twg4vbUMfM9ki0JRWnANnrpEFergdpGEjh18K6LNbvCVl2rKFzHPdXEXEDtanI0j
qlc+/rM7Xy4vBmy2+eyrmCBZig2erj8uW3y1voIn5u6/O6q10cNUHxze1O4f+ih7
1GpjKJBoF6PWXrW4n8I7D+hBIVQyrSclpbjYkYhvZJR+H46ep/blJ/fS6B+3QrS9
rJO+75a1jirOQlN+yV3gKnlRibNfX/tgWKRsvs0imn2ksgl4GM0bDqT3Ovm9WzQn
eJVw/CGBH7Y8qXsHbNJUNdVVW0NorBFIAnu4LcR/YvEqX46DGwv+dQVU2NXvZ/vN
QFPTD++Dzjuvotm7QqV/mC6F/CPSuWgrD7XNuJfI1qu170HuX5Rfgw5s/i8w5yn7
6cirFTDzn72inPBnzbNN4wN6eXexOmw4x0QMp7tzkwF1s+rgHMcbbN3rHeoOvCQM
8/rnLhsTQDx6jLcz2V+i4PJqeE/BQpS+lY/AMl5fzgXKRkL2vMnbiicadgT3gXi3
NN8bbD44a6ac3IGZZxEdyxAzX1vIJX9K5fFFjbkkcROnGonJYImM1vsNpAk/GJU4
P++IsKxu9tMxiU9r4gifn5L71hd/tEmo9s6K1ui+ymc+t50Y5fpfEbSi86KrDJXT
ljPD/gI4nFcADebhME+69OVvB4j2is6L6VFXOtF2BuFtubtr+j3igTLr5D0V8CJj
G+lMMxXi8jvRMaTurk9QqwIstCbPGbMx92hwr1yTPeyNmq9lfcQk9R8ff5JwjMb8
707MOpjfHnrgnB2VEo2Extt+ulMShYJzMG6Fa19mDtYAK7/YcOnWjRr/e8+bPvjJ
dQG2pfrLrUFkjZGl8l3Io7U1wkAJ5FqjQRq1dkYcK2K5XUFmZaujv5CNH1oUNS12
LPijOcZGK+w0jGD1/G/0jmCEXSN0AbK7gzOmAlLBmDJz275fH6J+YttviLQUD5Wh
826XVL2bNcnaZFgrUqE2eqLgJpU1LxSrJldnHV0NJanH57S4QaMHOCKz8n9MmrhW
wz2Lj4D+vTvPG/OIojtbR+T0djqGRC17dvBKVrPEfA5B0xWPEz0s9bWobkJN9Ckc
LMcq+PBroUVQiPtaPuEDvXX11+2TF6bcnG14Fhk504duayV274ba+SJmPOpGqTm8
XnytTVQWHGmtyIs9IqBH8H0f7+cODeSRqCddcQ7XaM3JFOJuHaMnu/MKaBmuuxGd
pZBgSuEIXJy2iQ7z51xh/wumTHqyVikWH8RnkqQrL6sBNy+cW4ZkOq/z6J9fuzq6
uJ0bIXlqPOdr4/DTyqUVc08J+EsMR2QCFb/98GppXfVaAbvsJtKUy8eEAv/NJZ/c
M+FQ73Owr3C6LfBRdaPRQfVl9vq5RwwXQr8NtMxcNHkX72v5+BIoY89yNY1H8HXH
HI5ktE2IiGNE0UH3Yga/JJS7ENH7Q6iu3zzoYjkzQIsVQeYFMb2TU52TArthPca/
hH7NilQSVE/RfWJ3i/H9muBoc+Jjko8jSabVND8rCwFNXjc2GK9ivSiCyCWa7frz
TKYi0B3ZKXeCMSkkoSOmsRc9srFrKj/VZ6cPp87HfpZt1RLY9PsVvc0b7CFUbbYQ
1RYA3varFkdK+TWg8muNkgLF0J7pkwIlLzs5hQCdq4OZCG2TSUf2RiXFSp9azcNO
Y6QXx6OBizjt5F2ARMJdyZ6tTAGLUyx6jbBU+tRM1qGF77MkVuyZuz9iionEKzjN
zpgdCfkhRWhEKh8tQmTb08UObymQDZ1ceA4N1DFTCxCB0lwh51arzOkbGnQeeC9F
y/GTo7vtFWOcO6pzo14pHKEN93YgaqkjqIPzOQJ6XZhHTcM4CroqtbUotfYquPs9
hOXRTd3W2VTIWU+wC9M/116j/SU9iGAsY1iU/gYhpeaUUddDiv7U6wnM5kLnB89z
/ecnT6Jdlism5X8dRwS117OPYEZipqhae1Gv81KzJMZ1Vyf+MZcfCrxi+1vMBwjR
uyJqb0P+dty5989arlBiuvPFsQOGKLlhTVCqy17MzveJlvsnRncOqcbLDnGEjgbF
xp25Q+HClxyd6M8g3mHZMLSqo6jwTvu10JKNZRsv1H+DbloGtCe1s7RZKwKQDBMr
SLsQ5h3eImAJmh8uwhk8nxUXYbnarpmzBze3vMVODRpxwrajaxIMcncY4YzytWsf
B6DCmSRKENfpBNzvdpCKVoOYY2sQT5ZzpDCl/T70OMkOL+ardqo6Tb2BbmL5l2ws
1panGN8+99TrNZnCX5ZAP97cYzTADKVnmhznnE0mLDNvpI6y7OxfuawPafFHPYDV
VJ6Nj8GPEt004RzwKXpHxvpRyjJZD9zDMUBXMJTohYrX4xi01vFMfKviqXlp+wRm
WKLMAdmj4hso7bzW20dY4X9Z9tCmIVlguUvwsDaOJwlYnpkqTDcs8BjREZ6gEw5c
+Vk5yBHfuHCPRcRP/T3vcr3uKGSrwnVYjUHv6DXuvNi80yk5XOTSJ4y2a0i6ZuDt
T0JdrT09TskE+2mzCm/XlGPRBm/AthyM4qXrHTeFG8PbpmtTD7Cs/EzjEjqDGwCg
JgGt4evd1dxflT8/2OWPe6oc8xJnwB81nENe41QT3JTEZNnpIlD643OYxJqUaRUI
unByLjpUguxfv0lv6VIj4zlx5sMMa4XeMmm/VkteHRuHf1BM0qMIa7COB0znhAOm
8Eq6MaTA7sPrcPiWjTbGJVddFJ+TpMzirq1Pzp/RC+aXFKqLD0koKDJOIzR65q7g
hfLzDHajPmcHQnmyB1pb9M0ogR+yWZdaf97DWiinvL3NdHebBeCudX1E0kzXvduX
XqH9tbikpIjbaetXAchhmwz0KGsnUxe438vCcRJmcqGKVBmvdy/pyBIqLkBxByxx
GKKNnwp2nF8kImydCuX++mooyg+y/1mI/0zxazLUJsvnk/lVKa9IXV5lGS4F0nao
sG6l9rzHm4ZXVHPAxLXcrcxwehIH4kldlVscrLzEIcgBgXGbRRE5c1dETNDVgNKP
syVYwezFd4BmznhSOqw2a2Jy2TJQwxovqwZuEI5V/PAiFKT1nUniSFSMgXsHMtVr
hmHgGuV1eqE5l7O5wvHEbO7Ihwy3cKs5dSP/27ta5ClfxHgh68dVFxxQ+oU0Qv4x
grKVWZBNglZYPc2yI1I4YB4+dr5uCh1F1pFaZ4A0hPO5BeX4FuDQ8P/+Qpd26yND
o9CQfBN2VN91rNO5GAo8h7lRzsBc8xJpb4/N6+KNBa4vGOK7Ho5cp92ztHok8YSZ
FOJdIoJ1RDq6PTIhFP+4TGzE7kUYVMFFaoNqNHwDdqhvhkhJ+/BpZVfIosITrRR2
O1asHY5LpDChg9iwvqJOEhWL2k995vgM2DkvCZcqn2Ma3Ew5J7eyyrbHCT0/AItD
O6UkHu85nCoc8PkogY8wk3AhG1vzNeeF3T/YWNGESTCusLvtAZr0uINo3jdjCxaB
8YP5yhNmHHmvbmXB692y0bPzetPTlchr6qlDCoIAgyLlPyaEmgcXwcTWx4O5CLWe
YAKG7rYdVatoYF5ZlSrTi6RbQ+l5C8ur6aWDwqn3blu1WdCUSSgEyTJUcYcSsQn5
7yEOot3zOPcpJK3XFZRDOswJLtHPF3KdjYFBtTqHteShplai7p14j8XW9OTZinzJ
cx8WIwIAIlsMCXZs+PtS9BO998Q416yWf7QXwSnp1ZDiP2gahOB5a5HK0DhElrXa
iCGbMTk9oBGMIRxfLPkf/DFmh4lge6RkB9l7krhBemGYL7goadMn8CLjrLNa+WeH
ekR0ukoD8Vk6QM1sGA82oUUMNND7yKS+hUpIccDF9YOkRinR1cfVsyUrYpg7FX6r
uAxZAeyfIliM5gjEA6QL9mbCi4JWiRJMStphVB92iQAtrEYBZ80Q61s+rnWYSIbS
2chmtWqCOWDD+qd0oQGwJSIc9hPpR8VQEk4ItIn8cspVZcT4+7iVSdZqkbLCRWWl
Le1GoYMVJ3IW/+QkSkTZaE4K7bkCDityRkvUlEeASnNnZWCOYS0Mhj5BZuGwkP2l
YbSBjt4uPKRFFs0O/nZKvcyAPw2ljvbE8XlU8ENMyL4NCPw9DZYHSLrtSKDtIQdU
h6FWgao3Y9Oey5RtEVlkThpd8woxx4akf1aygsBEZZoIYTMm8iKtpSmLb21V+HJT
snMNA9HPx/MfNagrmZvP/yHfoZcLCdW/H112HGimRLUK2ea0nqTv3IoiFMSNFL22
mSqPw6tt4BVY6o2fTkJRUlaoZPxG+ETkQTQvaNBb/f2epQsg8UMtMO5udtg3zaRy
JOS8tHar2r6u+4eJnYNWHLmKqYNW9O/yxbs8agj/jr9AIDgVi9Jm9kIjzGcXbTeR
4bTvHHlfTjXuaecPbQgFE+dsxw9ryGjTGDOkitZhamBqNM1wvAfNeuMJCgI53/Ma
CLFXniuvzTDD8AUJf2og1efyKfme1kK7VowIRY7brnMCt9/axK+yJo8GmhZlfjmC
VDNOxpYAGF8hLfuiDBOQteRuibje2VkUXiteNRwmK1RVeoHNOz15ScBC+xlVuO8e
NvXNf3oqrQOf75jkupxnIkGPsM7Vapn9zyIdWAONiiPew+D4BVD9tTU5NJ9ruXlx
s7Ex6GGvQA4ROByArCmliuW6FmK+p6dKnTTqLzUUdDFcAry5WBXn2akpkzV6+l8H
NjQIhPG8LrSXx2JJDbbKE9UlsqUXzFjG3goUBPb7aQW20/tCGcduwXxDhz5g0Y26
8Xitk1Cb01t0JL4ElYcWrSxgkvZzywvWVnN3lK0A6h+8UZBsUDa9Is5MZVmLs5SY
PRK/xNltiXvsx00hCEaFmXXqM/yyiZwhB1/JG7RSSz+mgCVmFfEAksZ1apeE6ct3
LG/q/LIqlwrjpJw3LqIoT9OhdCM2Nnmu4hjhLx1vvkPMwAvmdDqn4oWpA+X3Ftbc
daOXGF91PNuABMRK3NB3pPkCBe+hdbAzoyj0JT1+FIlKCo1sjz13JtusLtCyboWb
EEf96fcwEvEzs0CaNOPGgeQ8Pf5DDf+WVVIKp4CYAHYPslcewxAYxulznxpTxv3t
yv6OXEyt4wiJowFhVt5B5NAgjkR0928h9MUa7F3PMn/SNW59wfJoh3292Xc7Y5TS
dvowBFwNmxeodRtGi84h7mIHcUN8ExGgr8ybNbUI8LTJ76NPf2jp1kIOOmWpQlGe
B/bGg5r9TzfvIZ/bGElBdSyIMy3eHSUlGS7O+K9VTVhA8wYfYhIYezCzrZJnzlNU
daPIN7myepExt1iyTLVcwGwoYlHRYKSxvTHpDWyD0Zi1WEKVxKTVqZdVuGv9EfZU
TSV9iYnSwdH569POMZRbqRGlgFQlllXuuY+kntF1VsEAQkJYwxyV3lI0X4jJeLse
PbmXYq6domUvt4qQ1o5Lj9elKZaa7YR7Nk4zepQXkhryKzmqfB7ruiAcvj02FhUL
wn25xy2W28b+kHqvKR+lIqDBehyGf+38fr/jpCqdlNYFdNmQLytrs+puFYMuR+dD
ssGmZ0k+tiu9oA63oIHnEclHBgJ6puHrkPmEIXu3nvQfTYb8q+JlG6acFXs9f96G
/uUWlyoCS4y0/CXnzfSl3c/cmqhpRnOJgBg8/0/InpTVhyYC7zGgVnXsjoeDUqwQ
EBAiAk3s+dlky7fAlwXxdDLgHAt12fy/hRPdjh2hxvVA3hGs/71SpQf9PU4UZ0ox
341r1/oBmpbw4KFJft9FecbqQftHAbn5t6tzElaDoF0ufICLdOI0JIGadZu0tNIj
W3lz2URFNM22feV+Q0CdX/zeLHZ00T9Roe0ehEISJGCY/icqltyGZ7z55upRgjF7
siMqCxFiGvJmPB4dyp6Q8ZhHZiKIq95KGpkFJBWdcijfX4zSfrUOir9sFsq6n+Fy
5CjivF4IyjqKsMMhW1/2BcL+B0Mal92Hnzvy2rE82l+qFyLRy4wgtV07mbZSszzN
xfDGq9ulN84c71UybfRD6J4Ug2C5zWb2H8BKfJndxOVC3EooCsDuv19xqogL6QYk
BKUh24DcQ5HZbOiCeuq1OXsMiYISHSAdYbac7j1vsmb8AaBq2IUmEViBTapbs/M7
6o2m8gmPWidyFvuLcBGY6WkvW4Hz4SPMpyfsR4C9Ki9CSoiWhaVSWs2M5qWatguk
CLL42K2le/BSPIHJLJYV7KoE3C4jWpb66xj9ifSgSMbcvuQxIIbXTnQhKQNzWdFP
gLewutp2wTk/UJ21u1pF+hTJ9XH/reEfTjTYwhAfDJWV18qOJuTS29ltZrpveYX/
wPDt06j2mcvb0P39RTTawNlzD0rRgOqHteDvc1h/OOfN10bQxhLgk85mNAfC6es6
HYzNN6Oo5cbGDfN2G5H0jh+CpcUEA4eTQXCwjxoEML4dvcbD6f4q7gnkNaiodr1D
jqnFUV2qWD6Rwtiac3LyGwrOOZerAODPDC/vFgmyLjZu3cXMipqvhujH+fS/Xb8c
toX7fM6xgWfAtmxCb0/fS0Jsn0zDGsSqQEFfOOOo2TZsC2U7sd6lpL9XakVPij+j
XJFlm5DYOq28NKZAb+eFQqmGj7sPjATtPYx5q0QuFRK17RWdvph3X4TWwzVY4hZw
xjfqIZGvjLlE/acegby++vQyDuYk8YPKn3XC5SMgurj6T4NFvjLjIXROHbRGVSFg
pDUAjVFffBKpFKCQHJJ6Vjb7jZB6HmaKxH/TRSQr7ATpn0wWk6Td9w4EFsbbMFaV
gv1QW24TiuWjn34u4gRaQNuwiU/NEAiZxY0c4KSh7h5cRoedY7T2vj5mwD1/4eyV
YZCS3UhKy0qqjnob30u+ZRl4tvDrPyZyBE0Mtt12Re3cte89JucB+9tyinbVs3/n
7gGgZ5au00/h2/DhywvRo+R18Tu3vwmP1yoZjDXE9YNozYV55W0YtjG0lF+Y/5rv
zbhlYI6h0ZXf5mlJ3tsGenGO0IOCwHJAFyO3TZ3AoPoAUOakkh/amMJ3iHmjphfX
Mnz2iI5Ic90lSuYfF8/BwCOQeff+mre5daqGwXBwNfKw27wizRyKzytIk86WwTJO
jKX7I2FyU09hJoSky1sYqJjvBHmVWCGzViDB+tIlZDd2NDExcTu1S1VcrlVHcXYS
OSs9nzgN67PqMX4Z+bzcw9BjrTzPi6G0nAZMsBMKNM9OBEgsSpuC10moqbzyKc5b
J+tQk766CyhPM3ARId0tlTXYGOzIkA/Ung4gQ3PtDQdWgCMCFM3hiLHQerNmqawe
euAfncO9i/4P9y35h3zI+aisClLDsKEUWPcuT300zQSZWx9r7TW/suDmQ0EHoo7e
nnjpFQxM0aEEG1u0NQY1pXHiL4jA459tP0NRhqizn59aFRdqq7LL3tcrAjETf27F
oyrnx/bnuFK31hJzWSX7yZg/+s5JSsONfg/nJM7kYjIhEmGFrjJEM5sDw4AmKNM5
fWzUY1pkT3SBGL5FD4BC0qEfnsKOxGPAo476LuHZoQLYTc0zRn+EUk+TtuZAP6sC
L+sIuvloMCG5mDg/0PPoGmMKXBJeWFTThg2lBuCbtL28O2dQH8Ab//YnS9xejtPA
8luJrsoP4pEbmDAQPJdb5VdA06yNA7aq/8B8KzrAp5ZAK6zol8NucEDeoXjTQQ2o
jyWVeaa8KH2nYvleHmrtHWmYoRicKXYKTdWrU1fsJ9L09FmI6X4YcvMJacTkR2zA
4vmDTj10Dl+id3rHYEwWRz7EfJhFQibLdAYjxWL60Vg8aonOcXaU+/o6S5yVe7ZW
wiHMOQwxoLMUExYHHq/5VP6Hj0+uzsagSf5b+JY6n4CiPgP0vW0coxu0lpnLhVM2
geMEhh7M2O0aEqaN4tz9FxYCX6AoBRE4N7T9YeRQje8a4iYo+tWkmtMpViDwOQsb
jVHisULWgn7rSfJE4HLhgLj27i7iJ0z9q7utKq3XlTpR0u6pjTzm+awqTkfGNmfP
S61YHQ+ik9jpdIlp1nIfuRsouQpU4Ma2tGpgsmxQLxiVTk3+HdNorC+TLgDB2948
7vlAI2sCGtmkgQ9Y4rpXbG5wUcLLo0/lHUj0xz8FfB6ZqCn09b8/+ZwU2SJiXiHz
/AfDwIR4DTM9/c4Y/ytN9GVCm5O/7wW8qiiGdSRDzY0m7eNHTSw3I61EvJDGTuI/
/Duc7W4hK7dg3O/x7mtn16okW8TUJFkuVmkKfrBFgLXT01xQohZV7ynHnGryoo55
KA0PpTmbWjH9wink1Bd+XCwrSTNAif8Xs59T0bFzPS5amYRQ+Wf4OSQ4H4iFvpR3
8tr1rBbJ6PS4nsVtvB41jYUiAW0CeE75APmAs+OlmDcWVJbi+m5b7acs5JKqP12S
EMt4YfdaFsIBAe8Nqih9JY3hMZPua1KqGicl88YqerdSg4uPAJOxdVfIHNql4x9v
7jx6mIs7vcNGvZe1ecC7PzEf+rTQApbqAZ0q1l5Z/zG+gOzQ1zftcl9LdoMOf5JY
m16VWwUjbDuiTQdMnLaz+NirY9K86TiobjeHUW6XEb4pY/jNctq18cEmHtBbeHKm
5k59dOawVdthP2tzDuyunTiXOfzpzJbnHVawVmJLkEME6Zd3VQTm3cjvlCecLe7f
oaGOdzek6qKq+TlLW+os77hSERD+7R+Fb6KkNbs+L5fJ3geTuabAPpM06lSkyb+3
Zh3bcKv5z7SIEQf/huwPus/UVe8ctyUxK3sB3SZ4CSVA0ynkRSovD5JhoC/p4MS8
Xv/EXTLy+0rdOqWMaEEvaXOoPAjkfGw9GGwuxnaRiqfNVYwThyPXC8Tmy8hQC04a
TuLvehsTmluRdOfPlF71ZwTvn0GM9FaVISkKOVSOSikdjaTgBgrzWtSiwMHoWO8O
uTyuTGCiWtA+fm4Lr3XdHDApp6rJdbvaJR5QzI9UqHDKHY81lcSTJsMc0zC4ppWN
B4rE/SRmc2gi2V37BqsttoWEI9rj0+sBjFMCCTctyKpXAOAIYAm3yninOlNeULdG
CulTN5yPaN2bXy5mXreTl/fE5WayKaRrGdgK/2EXsHwKhPVu/t9wrlrPdWtQobei
TZ0dxRxrPPkh+RUtDDjYAVo1Bhn/D1PbZEWTS3yHntJA2QD6pMcUbnYHn/jEzNC3
/ofUKgbDK2vFlPf/L6AoyEbjUY7+uFmiEuT4X+6YtvgEqV9Zf10vwoK6tyMaT2Co
UYP1r8Tn049pOC1jHAqtSPNkM/W06FkMKnYwR3KV4CgSqHIjdie7btfMM0cRY8Mm
ZMr37lkIGK4lXfdxgqw4JPMQdLCGNmSXwVRcrL+5VmqpQqrFqM0cjDVtjet7FwKt
SqVQTdipUnfPebzkriKpRSxcbmQwJ4IlaerzD5L2RE9Lw8mGwh7/jKQpIjE6Sl/n
vNuEMGNxn62/A8ppiGY5p6a/DpD/MY5Rjw/wDNn7ik7whQEFVgno2UJZoGFp8MSu
cWs/3NbKBNcDiQk8yqEenpACQXqPhva4W6A0tneSeXLsIiOv6eDhHfis4jZGgssM
3ggRksqGFJobjbRbBvi5yamJRkeWCkWtKCNX5WE3BZulctrf9PS8ktwT8ur83sfd
ILmLMjXUANZ8LSN/aoSWJLHBtlj30Nd0RHpjJaJaWLKqOukkBX4obErOWQNAxr3b
WZYIplMfxPJflIwcwSyQFzgEZLKCJwOxpqjut+903sZLWGJaoKmXTY7ramJ23Hgw
c6lTo9/v4W1JWMMh78JaHEJpH34yOX63gTI9UXq1e0G7eLI9lk0K/2z/VKx7mqlR
onkDLkz5GJVeHPG/8ze5fH0gS0sdis83htQe5Dfou3hcLlR64GL0PtQ+Jxoj/xSF
s6jaCbqhEN1JKsdJBmVQheNAHZJgJTzbDgDuVY1Fs6hvJY1iUxUzRQB7tricuRnI
xmf23DO69BNs1iUbaEvx0aLFXSXuojm1ME71O0d2wopF/Xuiej40JdWTNGe6Hcgj
R0+RGd+mODugYpBAZd+sr+sPQTrJL8YibKJcsqSSlyuOdZqdd20SM+byoqeTGCg1
y2h72AOlcek/LGI6SenMBCTrRCBX5rjh7+max8R8wWXDDELvCxcGCvV4/jiV/YGn
aHbZkJbJY8SZ9XTzBeqLvYjj1zul1wmn3QYv63/DQz4NO0mGV0j53cvW1ay/yI7X
EB/luj7Sjk3/ca/6k+exTwJoFJ+9gh0P1rtJfWQVpwyBv3wZr+hmfRjd8XP0CDED
V4Ki4cRh77kX4Yj2Av1uQ6Rf0H3MYsiE82WYB6J9UpTfqZ7X21uUdRnX1SHf1eMD
T1MHBvMzFBXqNV3JkN7FQEV4dE9wgSodC9O6Np39dVrfmiboa8g8Z1fF9fj19Jz6
Z18q7+uxPXuxFI5Gx/w8vocFzrbk7LzYlkOC3Mr/0be3YeoKK0G6aLwDgNt6CcLE
zPc2t4QFA6OAjrP71lEU6KYsAbc3HsZeb9D7V2yZ39Sv6VK9lPqnxYE0pF3zxWzf
H/jiYtaaUYEKbiMzjtGVFSpobtUZwsI6q3KIa8s2N9wcJi7irfB/bqy2AGpqYLt/
G+697m7+jPseQ6/0r4AzDbMebUeKT0mSxO1pdHEjv14lfedW1sA6mp7H97qA1RIs
hGQwTJ6mrwssc5NdYccSlcxO1sKNa54hJvQ7/T5eNLwaVH9pp33RKLgEkWaPPhWZ
I3JwOxUeLxyOgC3PACVBrs8NbPYWlQ1Wu/tZfktLHRVheeBp6xGXbS0ulP5H6fF7
FjUMnPfVLF/iRfob97rAJitSd9cSsLc5lV/7hqzo/qbOnApwM1+AsikPykTzYpUX
iQLcwB56+gvU0gczoAj6/G2d+/Ghs4mATAGv5rVWgdPkkZxqnvOR8awzauG+QrY7
2D+N2PS6FKDST1Vc6GERSmiciakR4GVSMN2kpwYPaEtjIRW5vq3NB+BBu5hqyNYY
mYApWecVg7SKu3aAbAZRxoSHre3S0cJCRSMvq6VboFcz8KrxZQBP0gbbDeCDgpwR
486AhmlDvBkFTTwNCy4hCbrtB7xXalYh+85NB7P6RjrkFpKMmRqsOsTb3imNO3to
6WtQqSdC6Eaxq9Y+GnNkHoAOYd99oXzN8Ymzdw620UbX6E/vkrtuYKUceXPzPP/I
CnhZDOh5UBxZalmLsqOxerZ0EytTE7ymdGG99t9ZG8GmEUmJm3gAqY7+Bp5ZM5eR
PEAZFLpPsA9Z6p/xb0EHgPDHq6NAiRxLc+o0o0OXuIGWqy6R1+ZlcPJpijC59AbC
y0KuqEOf6qwSHTW7FeprPGa6DsWG7XqffKyV/OrMHHGpExrvAYNs5INHXuPEGC38
2nUaVD57HIm+zB/AgjXYbA2GGlCmHUT7/dRjACYUt+f6/pQ/oSo8PmrDmmt+E2ph
PBid+2BjM9HpPRmzVUXlqIHfGZ5NrPAIY5nabeV9tPlBp30q3+aWro92PWNaJuzc
HzySoCXUbnBRZe/c+STudqi0GgNzlalFvFkEdtqD797J4x4thITR63/aIDrzFKbK
/T6Ohyv64kovqWuTQb9os9Y9FibPa4PNE/cSkRZfDQN8afgFUqtD2Zs3ptxM8nVk
XTa91Cv2DxDQB4U2LG0YZ9xHS4fF7JYvUnqMRBcY0Wk610N5IPwX/1oeuyWEVr3Y
YSmELWecWd/FP5pEKq5tzC2PscZQh2aphYNoVDKoE21njZCw++4Y3DFQGrf72tCv
+lnWbOXx8GxoJnZbdkho4vjKm7geXPBM6ny7sBoko+0rDn2ACoZXltPoq7Qpb+TW
YYDYo4wjDDmIkAuultK0KPrZeBF0Jlxl0kqbvuwDEEPJVn01XfbBybB0x555KiHm
AlEHQY9iehsM+G1LxL1LvS7ANe2lnMLc0M8OCmIwd7Kd7kdeOebdurnXxU5xcoHn
Fbclf5l9PvSLMCid1Ox8wWZ4YSzCqfq3BixYBzgKYQmoDO3QA/dSLCpZCBrPepgM
2r9MSb3uFuY7fsZrErcJh7pJvkawteT1/la/Odcm4gavKj0qICn/7p36r53sKwsb
oSe1O87eqWdgGf9ovKRG82zbHs9laiDdJ2WFYPGons6Jyy4AfBKnc+o1Zp5ExRg5
v9Tnux38eiXM6XSyhEfrhQPAPXl82pr6sEKY0N21p2x4rm+cD5RCYZdVTGUGcih6
LyPbag+vWMy7TNayE9igadj1WBnnRXxOZ0tlgp3D1h89P2eDHC/8VZ3yvz7ooC6S
hraXXWyI48Iz1pY0aWLJp3hHfCZ20F5Qnq08J0N/rKFm3toHthZbpPI1vTygou1J
S7udsly4JDPRSM/q1J64h1CeQr6RGWWGLK7/LA4deQfV3qUP2+s17dVqA9pEzvFw
dkDkjMkvTKqr5J8i9HgW0/JdE0JQeo5yquLvBeAbXrsnhz59AK0k8Z8DOvD5bzDH
2Gv5wZftrGLzsmmANLTzzfJbhykx6F+eSrDqFOAxSoqDqLMnWTWIzJiiFsElvQ72
JWZNpSBb5/dsOYB6k54IFS3yxEXR6sNZN0VazJ0Wopudeh35pqpXy6cyFsKLrEJU
kNw863bF5vvhczInDPYoZCGe/PLRey1sO6+nm8CyfFIrzx2iWFwXx5Y8SVnydWb7
w/KUmpfBsJGXRCDyTVqVUisJp3kjtASd3adDC+lcmEj1IiRk1Uv8TmE2yP1UTqfv
Y+g1zS3l0JgyOs4VTgQVS+57CWZG5aCPnvWwRKVSeWoo1hR667ClU5uJVwOjE/C0
mgNm3qpBvBN0c1Ckpjg7j/LtCgZlsO4PBaCuFmr8vwz/KFXaY9HAiNQM1wA3A2Pd
CnWmeI7wDAAp1kkxK/TJs9SIKvQU+++09UpTroHLwYgMgzdfFyLTzMdiBfXTe6/t
HeVyx3tK6+J5OIbyhR4zViMqpvSwTW9GCIRdn/G9SBco51JBpzAM6IN5moUOWKiL
TSzk7cqdqQU1/oXvt1k6BOjk55PhfUUfOC9dE2uE/Ki5J6hphhwYhu2RwUiSHtuC
tKWFLegoCx30kB6u7MMOgDycKyw+SY4EGptOKeTvVns9VZyC+m7VpwkYg8vXhgCZ
Xfpx6JEmz1O3JK/VdGejNj0RdBi4gdDrcGvyp7YiMhgDoZvDi12ER0LCN6AVelDA
KvbUaZiQlOqfDw92Ds7YqmVdao7p7CTwR+b/9EWJVHH81l4GgvUBUed2Yk7s7m2O
l31zluHT3a+HZ/CZPAQIexw0yMOXxm8G47kEfGD2ctY+h1oCBzVKungzLhyDtrHX
5H16RbOmYDAh24F45XopKTXLHLLjSMpKjgCqnXl1uOh0G3DpNFqrUAE7uwgqVh3C
W47x7S+8Bt7bbJ1VBfuCra+Uos1QwLHpNwydNMPwIIpk0o0e5zMHx64+Hm6uAvg7
es+BOscCIC+OX4ikgWlWi0yqVGbDwlzFk537KamOoExu5pTxFKieoXkFwVIs8pJR
w4Gh5bwnZ88KBXcmYudID6DsGi9NTCj3UlO4l0axDP5TA3xEQ8rMLTJpQ6VWCsBA
4gv6IUnYj6jiqLQBa+at12/0bTKOPwFbGUwpiboSsI+A9YbwjE6VbeOdTedCQ+sk
w7o1fjnTbpniedh36POWFR/VY+n5JPbTQx4l0nMbzp7CamPy2WFHzkEpaQJ/lK0d
fELSw4IbPHojtjpaIJi3uz1qtyQEkcw9TVNOtAfFhyXoZsWVFP5ES3cuQfWIFuMQ
Xiod/I6FpmEcQ5K28nXmQDcws66ea61uY7Bvl//TM2ffGhiSlZ0y+AR5QF0UUcjT
Q2gVjjTL3p4zkKEbV3QBUCZa5RanYZdLoCQL5hyf3ZXxrQtdi4NzLf2OR5/8Giyd
wJTRhA4Y6GVK+12zWb1mwvl9sfI490lZ5BeUAvSzN9b3ItRMNvr92O8oyGUMgMWm
Y+58muOuMOD/XIc9OfCN6IMYs3dCFoNnULCdiYqqlk22VQRO27J3+/Ls68W1g6hj
2CVYDjnbSGlKQjp/7Eq9ioIwCjWvLZS7710R1sapLonVFm4j743hG9Vton4RD0os
NH5Kw06DgzH3KuD0Jqurb2GxgtGBTN+lHLpbu7nlzLTWCg1LcZ3Ul4rC1VojOmyT
ry8FpCtqZ5whf1FD5+ipPUhjBOp7MumLN2NFRgAq1N5461iJUbP6Z6OH90JOO1J6
qcPOhENwnI8dHPI0iSp8bj4D0ZUKiadBp80avHpdF0/OkpmaxjgOv1kua68u8my+
TkG7TzHpCLHNPL+3q0LD5rtjyOGYUTvmPlif8/ObIt4C+XnJWCEXzil/F6Rql6Ec
GtRfj4PwjcCILIW7la7RRMHZmJ/HbdG/jgq8kZLE9QHd3rMmJmh4YJGv1KCoUGPk
BrX5AgF6WdLpGv7rJC13ivEL0Q4w9b6OUjIPWp5Ie25fOzSvCXg1Fl83fWwweed8
svYe4Cb3LOAtE+YFBj+QgKqSKhlQVyziY0unWuPp5JiUArnjApTjq32nNYjhb3e7
3yA+VOhfIhdiG5qWMc1JkCwH6dozdz2X0f+3wPwqHai8NY6tWY8G0JD8r6aV6yQS
60/quaxMNJ9qn0qZaKuVWEUuJoa7xtmwb3IdSxPTxcLz6GmuXdjm+zPAaL7Q0qqn
yjpPrmqktoElrgGt9aHm/qGgCa9uS6YhuWPBPR9k/Uy9seZdcvme5MzoqpBLVFSE
1s9yYjqpoFJYRvMyNg/3AO4PZM+mtS+zMdhosr6UAXA19GyJMjB12h44bHfFS5zi
HWKqaNqddcAGHGVktft9gJCMbI+7weGHtf8RBb6vkeSGP8SaBuj9UGBQDgkKLMeo
7L52zIi7BaEZDcZQltwurWNGGYuHuYsjguY5nfxTmOXYBmH1hncRkGCkxB8WYLK9
sBeH0QadkRkuky+N6KY28qA9wQWB5WCBdo3ZXquNv/KUqzfNE5XD1Ch96w9GRlF5
gcG3KzPz1cfzwi6A0bgRKkQgY8ksqyZhfL8/Qu4pqiVIc65XMQs1wLUExGjFNRGP
15Pe3tOXgTv4pekPsp/L+Lo7gXFjGYQQkaSwjIS8HseBg3e2AqZSf0+UsTQ5lWkS
3wCOiCokVJMwhWrQIYGF1rpJetnziukTWqO1mlA3iyvkErnh4owY/IEz0YQyWMgS
8aKavxYoeF1xKiAtFKaX8xhGqP2OC2VPuK8keKhenxi4xPqNtZh+EcHzeZyliOHG
WeOhidefHpqFztHPpJ2mpE0y++rJIF8TQoxMWiaoO0lTTglYvDLsDEpNL7pto5EI
lB+kKgYwBuX77ZNBhq4SagQ9j/FYW0R0s/XYxh7QdQCjK1VvWJctIPyukFGHKS6G
7z5nVLrXPOWfSZON1wttqMdTXt0XfFfjG4xhmUZsWdPwAcbt65nn0AVA4BWwmFia
rgkfLa6hi4rzmMPGmvDucM7nN87OnPNxlVi3jPjLRcornU0Cn8QsRDzgwAb/CbQC
nTSVugiS91D4tapSSytttYXUUnKwTOwf40d7OaXFLzYRj/lJUB+py+VGUfxZHKgY
CBZq0h70UOOZBdOT8MZ3NeQ6UUYSWX7GGKfZOneZZViyE3FTUEXR4DusZXh3b83H
VdCH59HEETnGJm29Kz5j0hnPC8zhpKfJSIFXApDykI6TkBwmgY6JLVNtr9vSg2Km
crBa6c4ZRpZGGJR6VZQKj6T98uBJcjoxO969sXlYT5XKtR28fqnsGdoIwvON9h9X
pTzpQ2ordruOy5VfexrBy+BkDmHqZbwuHlcp/d2aaQ4Vkxz8GdrK3LNTv30XF+4w
jw5eTmGupwEkmg3r6WcdVPL2t3hlEQQb+C+8HYGBxxfImnk4bnUEVJVZqkynC9Jh
SUcnFp9LQ1Y8NGOawcAAez5yMAJ71fizNq5/YnEY490HJIZn4C2dQt7mV7ov1nXs
np/RQCLwFm9+31Z7RAYySwkwE16Y9IslfugH2J0+J83z1G01pVVl3BhZ5mItNu4e
b194g3mQcYPhTXer4zbKFkJBK20tvdtUt0p2RuNr3FpZlhDLkiKfT+RmSFmLI1yx
zbEqgYApV4FL6S0AwMdAxtU0gRHYmjhSE6UINIcS4mn9MsBeJokUHcs2VwVVnXW3
vTFHd1T4PZD+JA45lpr2p15eQFkvjVnkL2i0quhNafDehpv0Fl5JAlzUJUdDeO/v
HBwi79oZvIIWMN9lwOuo4shMAmqANKU05zW22647RezVMvy0EWgk+wmf/70zmDoV
qsI8OREbBfyD7ra+gt8JS4AisY6zzut370g1BVUNR+Dc0/e6GG2HU15EG7QJDbsx
AUMPj0o/NblfWJCW8zkgFG3wFCyxIYGvptxzqgau85tv5+08Atdmq1zw/SsE1n3K
XXiYCF5c7FRQ8pX4U4JNacgBeeqMPt0u2q5u7hQXH5owVxzqEVZPNMSrepSU3tzW
FF3vPBsINJmyxkoiVEloWMi1ty3aoPyOrLLUWxlS1CIIPchE/J0AKBKE3HwLOP3z
U0KGx+DwVjF53FSGnDBjmCfrpBuUgVQaLPYEyhqyooXCZLWxtCKNkgXzisw+CJsv
mKEXTx5ZEM+rcifnBPYnJyWvjF/E3LREuLi1ww+EuI0RLleNoMkgwdnefWRnoSq9
8w4Y/CtndKYwg1QpFaCyQ8Kfut4mdFcU1kH60+NNkru3PCvZ7bmvaL4j0ADTIpWb
wa5swdO3/rPZ/mDm4yMl95SL1qaM6PvwvAfEF027Zmj89iq89P2I95dAhoQQWU3z
KHR3HQkPVrVZvkSw0kz31tC7+uoE9zjiZlQi9yHLFep9vAZRUwbfi/R16Ou/uao6
AN4TQKOR+ox3Yqe3bOkUcxpOvOqOZseypdyRkVZrLvEuoQxFd45p0XtJ6hfBkEgp
Z3Z4WASz2a4U0fmRmEaxMXyvDY5OKBIqggvsUQQsDG0S5H+Sw3gsaI104ECiceUJ
PGNE6H0DZslfdWN31SXEfKo8pbOWtPCCBRZ/3wCVbfQsDZS36R3WoqmzWwa4tHeL
S92SsLSZaeg2RJV4V3KltnzSgRqK/8ru6wqQzw2mIdDrMlrndpuzRTQZQJaN5jS3
jfBfUnYED+H9xSzf6IHRoyjZLWGleUUDwEVOpRSOBPPWrLEsfK/HzvOeRIpr8z2c
RASO5Kr75QIRB01wd13bnVYjAPciO+bI8xIdUZfFkllGllcK+1ZwZjhIJNRJ0ScU
mksT6433Tw9RkxgwPhtw7WHdt5yFvcnx/isU6EWMkE1W+3kh/j9wdOfaqkdvgjXT
T88OQfPY0kdU80mDNVfm8wHJP7OUvMURL5qhQZZLfzz1nMRUzC9BdIDpzNAubTdx
iFg+siX48pZnedG5XF8VK/lFBPZOIZIU8C2oSGefXtfEiJzF3F8LZ+hSrERjFLqF
OibiLg7bCPkYDAe/X4ZidDSElHd3DO/fDxfZnS/7PPklCO0z+Vps9C8XS2aPDBqK
R/PPqkqghEfcVSReDOkwQlwW3eyrinThtP3PSTeC0C/ogXB3P0rZutyjEBQ2eRVE
pU2klLVFJz8x6qydA3PAloz3AOXUyhpsUgZGVxA9RgKBwIGOClvHRdhgniFjKRb+
ZIgpYWhytqiV0nfI6e7frusy/MOzSnppqrquKs9BYgtpuuWkqQyV7/ZBOP5Ar6l8
JhpOxT/PrnYpjUsjVsB2aq4+xmSRkOkGOkBpakvJ0tLpQj07zfj3uoc7qYRI/tHa
uWQcqcKs5hRPvPmpKmu3Mc6qQJ2gMwOtZnT9cNfcAL0KSeMBRgaZIlZSy+kyc/Et
BgNzY8BSnymZmXhUMtJY+l3mTpe5pTLw3Tl66ep2qzTb2L22MPuZn9ycYou8PcgL
j47tTK70hOa2S7CbvKCJLkAJJA5ia5CXx98t47jvxCsAbi8aB6bD5wmM7O6Lr1Xp
LiJTXj9A+XIcHaeDwc+OTa7dvF5zCc8Pzq+uP0UsKWrX6mcN3AXtFwMJyDbHu4iv
0dTt/MOo+seB7xcGD9eOyACdAi2mVfecicSLsbE2yqueATsbH0h5zjJu2i/Ml8ei
ule5HrsX1uXzLePq9u6OmnfL0oiWwOIjnDBlLHkaFSP5lxprstdjMmqIF6QN8vAP
mvxyvWqOGRJs/oGgUUQirEbP1zuMIdhtACEvbNkNtgroFFAzLmtxqTBZhdfXdFcd
we+8AZK0YgQRBK8OUlmJen7F2/pmATbQrq6F5ozH6kLalq1szCLiweNSX9PFsOuI
wfmyJogN+QF3sWVU9bzLWRVXq0LmCw/nsConR41ILxwkj6MaQZwUkupPP07vRmXb
6WeV7xOjiqFHpaBxKSyd3pyWagwUvndYUAzl53SiWnJuh86o6CcZYJOapUFHjLd1
Dmmzyr9+johDW1eyXmeM7f+vXgnmqlcHiaYg8pO+lhFuD428LQimSgExSy1zbs9z
J42T/G6HVeBNM8TOqdz3DE+kT8Cr0ur6Qs9yZDSjO2QAPJtHHOUe1ABHoO8GI8ew
uAVSGs/uH8n22NE2zOHWYhdf4bTR5Mw3akBLs3SAYsPu0VXjT2q29ATs6X+HGdZO
rs3eBAUXG+WdyQhTvnv+2gMctDtf9oBjimIls2pjm3xgPVKM0gnWVQTNWlXq2cV9
PvidEtJP7dFHdBlpo1xxOU7VpYHuSKa0k4Rm+dw30XcH8wAXMv9WEsv+nBGeidAg
Abimi+sA5EEA6sceNfXWHIgqYyZYn/D/l4WDyAp6uKHwM2DrUkAk0TrL0lt7KR2x
boPDrx8f8lcqum0y91KIiNppsR2m1ZALhBHXvpdYOFLW/NW4CNlSRFBCE9kBTp98
F2adlZcqRTOjYEkEZjkC+IuI/ZwoCRcLUdQT3iXFvk7LaDDGP/E5c1nW7+oBzMg6
HeBy9DeHTZ3fEuOQTlLzoQZHZerW/saAmzUISpJRNt2s5lvdW6gQOimLOVZla//v
C6G284+FeWq8Ev89IBcQt3zAKBfOpuIE8tzD+7C1UzTInh7rp9KG+iyM2LDP7SD/
qtg2Pooec2z0rb8/jHWnXCUjbX16ju2sai73EMpqwdR/VAjsyfy+6dcpP4jpOIPw
PU2Aca+hM6iM8HLnglZ5NL2dezgPD68qShDFH1OR8BKghUwmM7xdT80o5unnq+U1
ChW9vnGZkoD7qWuIcBWWiMhftOKyp+q/vx3GbPbCi9C8vdCL3/B1IEABbMtrVTw1
HWZnAdcgzMzQL3RTCm1uUetLa4MCBOecD3BXYhHuIcbreUvRI53zKu26/9njkLaC
xpxztuF0nnY9E1uamoU1Z/ztZ9aFHrw22Z5ZVrdwcifRT23QbpnjY8KKXAqfv1Fj
jXOtzpX7lQYfNJfHUMarL1BnJ9oQ3FR7qY7GKuhv3n11JmhULXBvSUyNhbMVvWbN
WjRMVutSeKnDHe51jUQ22WKJKkw0ly3hcexxLXaYLENW9fcBWU6jMmakRxmmzeDu
08B82tagsi0a+//buzwG+rdInMfxLyQQjaYITEYAlm1XGG17uwXaqeVdE9ww/fd5
s75sGPaAzC6OO0xeUKKiBG+LuZHZHF0ZKbo1yuue0DNCTmioxC8li7zjH1z9MjHi
s0v8QzrTcxfkWMXs4Jq2ODrKo+ld2KqRodFgiTWfCt+tqLgnk3eUp/fqKwk3cmYC
2AF7XMJFuhPAGVnBRXWlomgV28NzTEhJGs7IOS5XBUOLWHvtl+9gOIef/l+yR6ft
OVzTd03D5lucP16btjTO1HS/RH4xMGn3Ehi03xX7e9wEbJlpLBgPiBErGRMqR3D+
EvD3lhqlzxLO2+tWRj2sIikYFgVk0uz7hzuqS4+fHC3BYmFmIWkqYWBFN19vEFmp
4mUPGDpquDghmUqMRr/m5Ef6b3enyozmsitiDbv5nCfQd1GQ0F2TZ0MGlhCUcp36
fbYg3a6k4zME1Ub8OlV7CYiuD0tf1/JpeFjSErUHqC7qUeOKr6VD+ppVe5QEFvXI
ciwZ6ag/MNwduo7tq6M4X+JnY/9shVIUjQEJVVqGvb/z0Tzb68f9n/bFLc2uU1vd
Vyh8O0K9JYlyytUKFQ5kNDVL3X9M4OjC1P7owBH1+RP5FXs/cUu7zI6Hw7GFMeRO
C1m4j7AEOHeeYPFSamX+mHJSDkgQgXD26bHztp4FW0RgfzZqu/W58nU+zbslQ38p
+b0DbgYfZtg7lI555kJRI75mS20Z/qMXfFwkhOUhV7K7Qj3z+54+1zb7RCAxhWM9
YI8RGNLcN/j6Ln9KI6b9Yk7BgU1ZoRMQO94y8yeE7EcG7cyhrzs2iKph1ngRr89Y
`pragma protect end_protected
