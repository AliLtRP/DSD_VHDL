// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X4T9IuyCQL3soXSL6z3thoA91hjES4iZG0j/DQPEsZ5jIoYdubzUdtaqSLlW1bwx
QZjDCm3h1MC7neVV1SW/DwFxBBK87jsFG5IehT/9llvY2q9lxKmbAH9cfvxXvEn9
SW4gdRUY0VIMqbW72ravH1AbUxNsN+rjj66mmDgdycQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32304)
sZuvx4ExZL+Hukd7/0Sq0UBBVnVJuMPWv0BXspIz6csdY8uBmMgrgqwTXp7vmOQq
dLG6OMu96RnngnsHMKjPGHv+4p2en/a2+JYdiWXP4f4qlvag2WCNTQDlPsEv763E
ZqUt2MnNMAmZBAwHUyCFA7BM6OqmfSx6aCG3PdyPb8RGS7J8U9zUJomdLkOQiYvd
om33b250nHpmXT94o8YSseIiRbIgDslfyu0ceidqus9YzB5aQnz2sd2hbIKoeVt+
Ff8Ru794uxPLYHyHgG6WNBqHpYCYOtAx0omBVbbMuSTGecdOAog6n9idpu5It2jg
oDg7FFtnNlJHY5Q0+zlCVxSN+cLufxoyElE4Mt3HrDf1o1e6CVRojLpYhfMIEtll
jVv7MpfY5Wuk0SJR/5UgzD+gyuqHlmpwxwFLNCcL+0jMxQsj0+O+5Q2//AEfCdD1
LMoMTQegYK5n6EEXgEYB13pps9TLGhl8Bw4c73G3YR13bPkaSzHNTz/osgC7Dt/d
6n4YIno1SX/qbT6O3/+Q/wHwTlH4SY1pifvNwTNFGPtY4i1W7ZWZUVEcGhxe0PFB
NrFuH9f3ZydppXJanU3HnmwnlX4ym3Vbf+LyKWp7f3HremXyaQK04mb/cla0eIAx
k7u7mYssOG2Go1BLdsxikozbewG3120F+9/QwXivbN4E2QsSEfavBF6l/jkkRGxL
CfQCjvpW4WKTjieoVVQlWjulLUvi+L5iLDtifsNFg20lb+eEzVOKu4X/e/L3nv2F
01KkXDNLQ/djeNE6S90HrXSlT9Kk7BsJe5Zp7ACmFCQN+W1n7RkthYllIqOT1M2N
L+n1hyW0dnubUkPTGqjRV+S9PLp8g/Bax43y7NEsQI7mfKoBFDvSpHetrKReMZVN
nu2GEZn020s4WG0NRtruSQt5EtHeJhuYKUDTl7YKlrxSdXXmY87o6x59kkL9YpIH
kmbMf6LmOjWssbgy69QJOTY5YrWfd5Gpkfv7hEQjUc0l4QRplBvuJj+vVAiaeaHT
j0RrlXcHArQKe8Y20k+ae6Qx5kjbSCYHBspbdsAafrWEOZFjKejun5SnN52IY59T
XIb3Xda5zp9WR/rZrGNV27TarEvqJERjdiXQb0JH+hr20B1XSMHpxeY8Pnq1Uo1i
kcvlw/75txaHhPk5apNwkPM2CWYCoGcL+qqcRCtTndWb6bCkYbsIETL4Fg8a4uSK
yfJcz6Utc8rXk3oT8EQTbQsV0tIrR5/qyZdxvA9gNf7C8whWWAVH9IIQu9rGjuX0
pGI8zBlApafIMJQwyMwdUFbF/3irfKBw0TFX3QtB2HoHKLGdsE6hjVBAiNkuOJ1p
M0BO0ez98G9K6dFpdDGAO365y1kGDZkvkpfUspSFy0yajuzIhy7RH4GB+lj2ij/f
kGBKSlwIXa7KZ8PS7arNbfKglZkGbxro7UcgPJ2kITzwNnKn4HjP/EhN3/q5+J5Y
0ER5QuSe4TKbRLCAOK4prQZael5ua8MiNpMktd3oe+rB3k8lgZjizYU11VuuvSMh
V5wbwKGjAtFr4KHeoBt2zVBtXntkxQel/U6bPNrrQC2+R5Rh24iyWzsP3XDW6mrO
5VWldotJeXYt0PB7ROTvlPR9dlQ6fxviVq7I4Z8eLSWK4eQ8VbaM49AJQwrgr0NQ
9ihVCOyTx37NVCakvPcDhga1tv2Hxo8WgLXWKol+GOmERzSsbJ+0+GU9qOWW11xR
9GzUaWyofYDJ2S36y1oDUxiKGf3y0kAiR6lWh73vyjIo2ETrXQ33h+hIloIn5n3a
+eE7EZHa4hGDAg0AHFxXO/LhPBAjdB3FqyG6RELwxVps+2aWZdxBQ9QQCi9+y9fg
ruQYDjOLmFtClLRtcRAV8IjeXja1PLoUkh/7zBe7t7t9NXTUDhpxKU4VQ+WEKVnB
ATxWXQulw7RYaWg8xTxO1+io8fBCbIiNpp5vwLmZ5uxNQJZvEPDoxSZqJ8Cwn9+4
wvrWfIHL/0w7SYpq522zL8KK6FOTgX1qrTDL7DiiEuvXEYmqAN5qzg+rgFxf4FCb
1jDD9IPTeG8IYoieFY8TMEG3UeAiMjj5YI7kh6D7CM4yj70HxCQ7TmLf71R6dqRz
q+BMeIYXf0QgUkhRe0H60iGWqcx2MHwDqVc8M8Qmgf+JSPxZqWyOAaw7caovEPQW
sCpG2G6/wB1Nw+zWxlTrUIZkphf6ZCryPTj8v0JoePYJ+jJg7s/XvYzmZgMDysvx
0RQi99ph6H7ECbNdtZ4idSvpi4wgW5cvfmkaM/5b1iWbvuyhK/56JXENzACbZ7/q
GMAkw5pUg3I6kH9qwJ03Hsakg64FLmnEybl+zoRynTUbHM8J3IpPAx6ju7nG/71N
rZKV4Yh78TobLa2ovaAVCNKZFPF2dwTzVcoUQsQLsZinoHdVlGB9pRx5HgXN50vB
WOiao3vCRJFUQ01Hk5iA0YphdiXOie4EaarBgUW0lCM39NAh50kkpP9RZacSTYzA
oYjRMtImAuQ9QX4df/ZRKpuwv8IEMS88/V0KBZY05JnDhwWHtiOeDaSz+tApWffW
/+ao1RGoJ4YGnR2iU9TI6mRJgJV6x/XJn+KOhYKLOifEGWOY08p+WzIwiYjgNfP/
13Em6l63eZIKkkwLr1WkvS8U2Qlx+s8gMd5Cu3n2Z6ZQO2LspP++sn+CYpDp7Y8V
rBMZFxoW/+8Pco1XXeKTOyXPtPYhWYWXLZ5pIE5boaBrPxQ8NB40hYYzMSqCJRAw
0CxBRDj2d4OTt8uFb1t+3qvYBYu+cfp2HJcwJr3zld7iqLR2ukIkQa+mGPWzsjin
30em1kLgjviK99sJR65aoScu+cCmsH0IgvbFb8zy6fUoOfY/UDVKrna+ccANkfzi
5yIedZzQ/ldddmm+/0OteBb02ovm73BRbpVeKfGQgROpfu/HPItBEiYCjHO9M+Uu
zyMZF3Rl33O/g9v09r0x5XSN33icbisCJmWexstBflsOt2rbYG3PqMjgXME02W3o
g/OrbAyahk1c891xgJZI81yYsfvbgTulctjeFQCZCXEKlw/+IdYIDRDFtoU/5AdI
RMffnedJjtMRlVAeZMYpESiWwEbcKPzCL0tpMYh0hJmEWzBYlUmXiBnhjwjsikx2
WP82JyL8lBNtlkgxgN5eHsjc0R/blTH56Mzqwe5+UX0cQNy4SdWwXbaIsAlFGVe4
Z6+sH6nZQ94VCcDW4eaRH3qnUwLqQIphc/rLhahrZSviQcYO+/eeKFgkiXImv/5+
vl8UeylZ+LY1vbOGUR/mt1t4VFxC73BLQOPLzIpOdd4k6jox+WxX0SM0XSj3VzHo
QLVH8lLkPAAyLxG2MuElR+SOwRR6O2tTkBg3nWIEuLxQFllkxXURV/JompqEPkMv
qmIZoQwjuCIo6Qz0N0PJCiXuJNnvQ86mcphdZHhWJGNY61HDrpEM+s68lmufzc2D
g9WnRSU7d/MBHNubSaWpUhDm/arDexnkm0s2uQQWX0mWl7h4hdTUx5ZBZ56fG9st
GIJrFcZxsWdyUWHgZPQhXsPeSukQ4G8mUg7XMGnz1Jebd6WpLTbM47VFOHTRYUZK
MiBHIAJNE6aUzQuEEnJSUbb1c2d3qGXe9S/XrtvfA5yjV8fqSH+iKcbz54uL4pKF
yEKtov+jJYOl/84SS1QEgjUScHBcc1atwURQDUM0Lk2025OETOVsUTx4ew1Zvvhe
+a5yPS6w5/XXaqFMf86Ix/DG7tu1Ddy4MkwI9sGJR+4bMuCn+GDtYFIPADGQ0UIC
BeOnEOjaBBlFbA390lprMfttkdGrXinjzKMBpFSeTX+7MBhjnxfSxWGm3F3MXuwb
+g0Tb5ZGdqaLmBLnfltYE7SwygkK3F6zX9RtBm3pcUilH1NtkpzSKH0rV/PTM5dZ
t/dp2p2dtz1hPmdw/KFGEz00JMzwqfoqkbvux19ClcwaBKD8pZxKgEHT4veypf9p
s9bWpT/0dRF3XIV4e7F1mG1REdbH3RMEd4p1OTeIB/NrnJEWNRxzcNeeB0CijtQE
bfpuEhl1qQeK3e3NwaSe1CCP+FMphJlsIbPljQipcsg4qsMXptDGTq7Ls5mPdzwq
rm0026ocSnpjDg4JFm4HK5Bz4dAPGzyXyum8jwoHRetjyYKBjyzJfoc2pcK3Le9B
BhvqNmhYUOXXWzR1DBVQyfuUnPMTIHi3/AcJ4xdPqG9+DoEGO0NHa1iO8r/SNTYj
A1xG/l2I3wx/BLtwAy7eyEECOA04+mRZ30gp7eur0ZOv79iQ8Z+81781kl0vx/ys
UhmHqR2LJtHlFXdEF0tm+cxfxOGzXQ7M1mGL4i/UucR1pxhRsH98raZYiLb/mRsl
BcHw+YML5tXOalvqTalJW7/EGNxoc/fBuIZRYdlgo3W1MLgINGFLeWD8pXi6FfFN
9PUAB/bEKX2Vyb1+YzA5iCh2WaGbzem2zDjmYj7VjJOYo7KVlpFBRCa6v2NQ15m8
jyQRgyqx3GpHidWVUPjXEO94mIsySHWsTfP7rk71FLfcIBTsCaWPCd+e9CzuLzTI
np0B/UFoKjV8cBV7BFlO29dl2/mJUd49h+gCJDZcXrJJ/+6f4al05DH7Dip4IcUh
+YqJ/lvvEvrVanoKiZ5v2gSzv7F4bhSwoHwgQ12CpO1lYo4RYHtERY1V4xhHPSDw
yzpx75VdFz+Sf7ARztV8P8Ehn5ukq2UkUVjkZKp7KjY6pDqbAIzfVx2yYN7kqMpk
YvAOLZ3lgVdCM/Z5jyYmRQ34p4LbDr20iNX+uA/RrxNq2AtX11OTnLjgRh8xCODQ
CwC1SvhEWM5GS5p5K6f4YI0ftIrm0+JdkXPRBI9R+pW54cUnyOgrh8vDBwI5c/Jy
ib09qUhpp7HukJ+lHbAqIu1XMuhWslkmUBouBlnV6NsJnzz6s6wfbZyqfAyUEtCE
7WsEu6D2Fz4OQtV5XuglVUahLqP882maUrnhzVVmQM/nP6aMsWaGgI8+Tau4rDDJ
Xoqd/g8rcWU1eIzQUvQlPDVhL58Jrh38oeB9QfrkY4I8A28DI2/ofLMdl739vdqR
zAW42C96NKFDIYMSxll8CjngcLCTb95uNRXzhs1iOcT3o3vlwzTs88iqrfW6dOQA
iORQmgH0HVxwjZ0rRxeEdcNpVjDlduJpyPzC2nADUTa3RRkImiVYCgea418K/eKp
4HUvhpMXPVTo2XAjiuYUmVoPZGDo/un2UCIBKC1a65rfpp0VnXu3RViZeiwzmE+m
SHdxRmTb2+GpN5jFpEwPMHl9Hz8AlF/X9CLKkrvwq0+peEHWGGftUgUg6aAVPDjn
ZBAk7s2KNBfHD1yZBk45MgyWywIkH4C3yrLGmMajr8PqTkhEBhjuVnqa5HrqRrvJ
wcf5xMs9udoSO8M8XNre/dK9UF6kqdw2vtGI9KQ/go3tXP6bDJFJE3PJPW0wxdXs
RfeCA63MhimI0VhHu4+RdIUOMpf77bviUrd4ga+VZGeDBsNY50gtxlA3Qcda54L3
ZGGregzuIejDrxtbby8BPNVpBLLUGsjOdjFUEz2PdMJ+OEBlByu99SJOVjy4ecsm
3aZ9jZQb2QEeurv872TKuyremXpGIdqy2SdtllpQOIQBlaxU3I2JtSceJLt+7jaq
BWEo0xGu3IyclDJan0LFgser/Y0hhMI7TJmgEre5MZHAeFq/TlLyerLqWyR3hsiU
Pj+EWC6K2JLOoKQe5qKodgVe94ooA5HKTdGlHp7BozzmhRnPsdQmPBZ+8Bs1IaRa
M7PZ7FsPyWoyQIuteGxF6B57RFtLUH8gd7ErADbjpNv0Xy9sYw3nYtMUjFnd9v1p
8ph2WOn6vnfOfd+241ChgCt82dGV4Sc2W9xbNLwHc01BtnAhkj4xiqPc46voljej
i0ObHOa9rGYtZB2YX7ucXgdz/Zr16v9Ny2R6A1rYWVyQZP3+mh0GhkwHpiGFanth
dpYGFwXvNxomz3rRzduKzMd385CPhkjvK6IXU9Yt+M6M6Wia5K6MAQ25c1EjwTUO
Ttz3fNen/ps+vTcQYmgcyeBVwF4ulR7wO2XUok2P+qt1vcJwAQd6E+Zx3Y31RJFw
oq66gpm25vwuEpmlTp/jYRXsBIBWQ6tMcMY7qdohC3AXdTBbOt/sLE7EVEMEhzCk
dhNtK8ujhpOI4eICSjF+G5l/K4HCph9mbi6h963l8nn8wIx7KjXWqgUIYtxjHu37
TLSVGlgJ67vzNggtTe7Z+c61Vt5FrBF1zD2ohQK3ZTYPkWlaxkvtaTIV5NYV3Sz2
LKswaJ+E1CYHKkhF9QWpPYiQOm3WiY+rlf47IJc14MNE+O0rR7WfgCxtsPugcvpk
x1dux6vRf12xq//KhZDnQzScfi2bntl2vqS0PQXNMXQXYuFute9qG/E4aszma3UI
rsBvk3/7Pg9mjt41WE91KxEhIasuWBGA0Yc+lB7GQMeBUdmHux74TlH2ooJXz3FI
JHD2WXB4JbMeBoI5/aLd7qwThiLbZuLxkAqDOKA9gDmrZlggLllW2MRBtQAtLn88
pfZrwSBBsbAfOP+LjrSf2iAQSnWFef88zevQ2sVsYYuyy5q42L83xiBkAn1gxZcS
t8Q9JXrlgxH/VEwSMCHqCw8Du4Nxi3yeO60Wo1LklZMTIRnyai0T4jZQk7fkTThi
MBvphVunFu8yp5mxeQgx7WDC5XidDIcsiJVj8AepPgfgnZW+VtuvHpfxv6JwDY8s
KqfGMeFL2HI3PyYtz630ret/aQ4avbY9kU2GQbaDRQjZfmAi8GiuFM/IssbP7Mmr
gt5SrXfJyHuWVsZO0EbcIPUzZqLVrG8uYC3guFfEe9oHVKw05P/YpT1C9T1U2W5z
OgFzxHSygmgceS063hheJlDpXoCx+HWWpqsT/YOWeC/UPO1jLGhpZIhc+0iY2iYn
k51WhFl+2plpuKLOIjwSUZCzJgcO83T5d8lXNdHa5WyMKLKzTlKKR5/CliQ39JFk
yd/Fr0bGPG2VOE+du9uwmnDwa2sHKEaB1hu3kr/u4MQ9vaWzHHEpL7PejR0RLAc1
Yzw16p0Zc6FtL7D5Q6yg85e4zekfNXdLIIfwdhxa1t16r8OWWQkBuzwEtfIr2ns7
ZPcUVrrsAbaAvx8M0R5cBsouzhUQQBphGjCT+O60TfA2+nzrlthEvxhiYBYTOH/2
m4iaYaEFL083nalJMlO/tDnbYKNklgjaNiPelPAYyrRTq9b5/96Ya5qktxJWzrXT
ikhS+y61FmxhQrC/PHpqtylV6K/+os6Xokz4j2l6PDl/oLEAi8hqqvdW0/RM/NWR
GxFiXp54tgZGHGM/V97jCB4jZExkWopk0bTKEfnT6gK2nWkA1WSOtyDQsLslTaNb
OzXlDpXZPYAaMIiD/4hsPzoGELADJlCj71DVW5jCvqEd2YFh+VMd383WKxSwo0J0
BEm8YbFj2rJSNHnTpTFXGZMv5mitwAkIrsJ9+R8WhvVOXCSGJcVOsFAEI/7JnmxP
sKR3txdxsHv+KGFftb36XRTsINixnzoXJPXoQxi6px+NmVsO9zaJo5mM7ulSPGns
cPGEeXqa4q3OJMscDN6jLWJ+Jdo1Gh2btXmk7jTbynrkg6FqBozfszyvJv0tQ9w3
3okKFlb9ZL1K+xZzxXQGlSwAHUj5TcFqCRChscf98MY9fK1elbeAskGbJ159Z6dn
JRp8CqdV+wRaHm4u71f25rfRh8ChtPb8e3+1iNyUByf4AWRVbfut5g7t97pE21rI
cdNoNH+enWUk/UFThTDg2ZbEhmFOmCzMDs0l20CeFqFBcYIe6AaI/ll8DlkYe3mR
jEimP+OVpayvhCk/HKSWThQvhXzI+GlIK6vOI9xQIEDKIPSlkLZ7K4i3m2VEOaey
jw6/dLwYdWKow+f3TFEaP5I5gwwAqIkPLuoKr/tRqvCXtTMw0QqhF/9usT9ES3R7
mzbIjiT0ZICSrGxAomr+TPp72f56SaukTJVvDqvvqDUOUMHZDZ/gc4s3dk7Y1TIE
xcqspk9xxpFJQkaEtNxxh+lUM8T5BVoZnR1UwafiRYwfnbRrkDEpDUB6ahDfz+Qi
+II7H/VMG/RORNTOM5M+ElE2/MqXJ0iG4q5E5Hn8L21v2TjWyrcM9NUDJUoPd3aD
CndQacUEN/LosovZQxJwaJODOF+gtzPEhjDwVfiY51StOc0mnmKo0h+27SMIFw8M
xQpDpwtWVRbyuj8w7aIr6dWlfeQwV+USyO1mJhqQvqoB48XgfXpnE/ItmG1gUj6X
a3t6XaQJN8zcDhZQpYbqaWOdA1+PZa2MRkAM/NMa2MEQmYkNqUrfGHeQaPTF8vw7
jbQ/C8SRYqCRrNzD1YTYekUXqIjFcWCkuvVPlVUeO/DE+ztBv9FSrqaoapHwae0N
iw+MsFrjm5YXiOZ0D01Qy66vJiykEiZuwp1YOI3qpN0ezDjUrCVR/3z//JZ9fdwm
UuTM3/7ScZS+/xwNRGObF/6Mwh630hZDVuMY1eLKpTZsj/TFrP1NaaQ8gCKkQfJ9
78cFbxehzKEL/MPudg0IQCtyDfdm5Z3ZyaOAjlDXinqU61AIBqX4BsVcCO1iCi/M
4lNtJEnpvVsFFN/SCTupk787hZPo/HBv8A1aIsKI6mP7uL2Jud0tAwSDaxxuCAlM
72ZhDGMCMG/Z0T2qNh3eXwtHKmz6DrZZm9652BxgfIOcDHH8TJVkjRxF7yzeeyjn
N97y7ZW0FxvbMo23nqpzuzLjOnPc+X5xQlRIzie6I25EItZeIofOlcFt27snfsu0
+T+FY7gWrvl2xlenAfSf+5qmJWVDNA5GtEtp9kBntH795Km2L2xK8Q+xCOMRrzp5
RXW/7R5eBjRRoWUM8EM4Hzgu1o/8sojEdvqaAf3WZGGpEFcZH+OebRF4Z1bm720h
qQP9IcR2Ln2geGhygEN0DcsIAyy4rd+bazTCQym6PqxYPctq6G6EUb6C9Dvvi6H+
N6dEaryeR+Tsw+6Zkjh+yS+i7RnHMc+YJcKiAzg508EE2croNoKE/nygDfniAmC5
J7+zTPMZjoMzjW5q24mfewLA/YTLp8HNtv0AnhtAytpztR4TbMTnt0hs0E6TdZt3
mEX8n+PZjvRgpaIh0Sg6mSlKxD/Mpld58zLPInFSJ2QfmDwj1FftzcQQ7nVCCZpn
1P4mxCwMur/fxOeqa+M5uC8lJPWpszTSiaW0Ts4VmCUI4f7ILasQUS/44JN6i4PN
qk7yNPgOV0wqUzzYTSL6lasDpXJV3VWyn5FOiXjMQTa4Mf9UMArQ8xZAR7iggdRE
GaGXqRBkK8+tuX2fk2u6uLxwhNhbPI4PmcyoTbycHATUsd+l2zCn7FMkK0MZtCsY
HdneC5bpVJFlQ7DyaC//ZVENvEGEW3sZL4zjXNE/C3CEcCfZUDpMVCf3Qe0l9xlz
ynJzL20WyRkiEQHFkSn77LbfSVvTVPH2udyAIuz7Fmp+2RnfR87MZxJHKpEKngE0
20X8sL2URAOxITsJFCkvstFGfMnI6aUKCsRC2qVjKd9nVbTE5JbjywWYiPRpmX3M
1K3NDwRo8vZc1mMMLnUM15rFZT31NLlPeQXiC2aBQarxv8DpfL8rPCzfBJsJ1CYH
LqWOBk9sluGFA30AehL9obb2suUjIdxGnZ7f53nMIq2+4LTRBuqhseRotZ6ua1BY
gl8IQp9kE9Vvz9AEvl0qq6aAmJA1dzuWDLgHE0j0dW35wWKAFtnsfCPLMypV+M+j
Cj56bFP0TyFQTSECuIEiLBJKd/sPO6V57hSqemlFPX3f/MBb7PEOvngS+g9SxQEr
dS1cUoipFiqcwV4QQbpVjLvBVDWDSwlwVWQkVzCyYfA3PXn02UXb1qobHpPIc/4B
7t0iyJX4AXUrYlptZ3Ke8pIm8h1ZhC5R097jIAdFYOxPkSlKvwpv119mPIZZ7n3b
xlo/Y8J0tzCk4PsXy+P5RV0a899T9Hu5Er1PFfLIeGaJ2N/v6Wm6+L3xbA3kRYbP
q6+2I0MvWbB+3b2auis2785b1NgIGTyrixsba/24syAZvVCGrILERtst9ajyS08v
FhcrwMPZbfDIc6Ml/0ge6dCQj6SLeo2GhFlsHi/xD5R+bwI+DmOFanvYDzKciZsS
+wcbxUoA8wxO9/DivHIIbFBKwoWgJmDm4WumnWtElrKHydj0df3f5n6pOTeu9mNz
qR8dAMV/ZWy8+QCRc7gQ1CdJppKtdYlMA+Jt/lqNi1W8n09V5qca3MdxWg4vcXLN
Xne+Nq7bJ/tBSx16bu7pRqYiumLppVxn6hgJ1DJmYxY5MHqg5xEr+8HNrXlG5uvT
j2lbbG0m5Gxjk6y4KXr492Kub+wwos3LgXMfpiV001EWG0ExlPqkO1wdL8JQ11er
k22h1fMrENq7O9+An6M3LxeeeJrcSLaubiLVcnGk118MHZiu+kJ7Lmo3FYhBjOUv
DuYW6k2ROSoR/qKoT4B/XNkYRs3z4v1TUGsibaHJOGRA9x9Zv5cftsDlXUWiPm4i
jwAo7sIKtTEcS5MWADGL+C4UVhAA++H36N0OTHLDjqRv25XO3hsJllQC8+5YLJaB
KSo0+Y8S5qe31/iZb6vv7dsJHJyYPxDpir+opDx8WvAgX2OXLl5sSjUoY7ZR7Cbe
vQnBDigf7Rk/8ptZEY0Jea94U7v0sg6sPgkV+5rNsVScVIAGk2WPTqDJPSXnFyVv
0Xyr++AvIkCT2SxQtFIrP45yty0X3gNkhwo8Y0OYvmbust5uzX+uAvvIXTo/f2Gk
jjjXCK94JnbcOW1VlJ1qERmFZyfK57tBnOSCp3Dvgji1shBeS7OLwd/i7wnOquwF
HZ3NZE/2ngZ8qlqzhcoIZiC/Zn2rzBTOpQjeFaFWtT7mwjZHjBC7IZDdmEftU6ow
GSL3zHI53aTrTGs70yRVozj1ja168IPGRpMWrdIz5LkSrRB9ot1ukbZK+lhIxpMq
wjJ64Jr1Ni8YsiTsZTuHU/Ngz3JBUSHv9R0fe1FsV8CINj0W6/3X5NvGoa/OOAYz
1eVRJSKsICBFbsgLh+8dlh0Tn2onJ2xe6tAUG6rCKAhs13bezbTGJYGummGYatST
Gi/wuRrhmNuLhLAXpRmTBoM+U4lHpxxOl3ej9LCD/ajDE3JzIl2Ene/fCF05tvV9
yAiaJ2jP8DkMRLuEgg7yVXx8EBApM5EmeUW7T293FJmsrqLWWoVitkUGctCW0UDL
UovZ0fldr1a5YaT9BCMpzYQeSSBgJUpQUitDZbqbvlRjNOP/Eebgv5cCPdNhGcfA
XbiyWVo7i9TaJfL+8Ci26yWrEIrqdwuBDsDal/BVfH2DOLQIyFmpoXtEWjgz3ik5
Cu2Sw54w6I4oyiJ5LABUhu6fxL8N9F6ClqehvXez4M86XGgQGiSAE056RDtskAeh
ODRsEUIhURcuIo+eKmAlT//BbDgj6Flnj5I0KcyY7zIS9qMKPGetDVmkmZ1EgU/S
KW72zkTm/k49SQst5X7Ci5jy0yeBjmqsP/yyVovYX1e9N74+YdbsrggjNmLY2uVw
k/6gN49a//jama3pDo8nkb7qBQDwke7Fgg5hwX6tpAVSQQieQfO7dB9d7pZ4ZcHO
eOKsPUBTLIKJ1UXQU0ho9XhAWkuiHDE7HRMCEDUvQRVgD9qFVGIA3i/baKkAs2te
H3pewSanXoAhbWbOLfIAyCBb5WUEVPrvhWzZqrMNDDqCG7W+VoFVUAhLfL9JPrwR
RR7TRk/96RqtJ+IZD1DZ5jWz1kHU1FzBSF21DNbW1gOAmRaYiWya1WNhUbA6xzaN
NnmaIEE/iwj4IZwUCnYMvPEUw4UbhH+O0x5LBR+1fIN8xhTTyc/xEWPwIkiClkO2
4yBoi4ggQ5nV33KevKEOWLwmJrrP3WzMnXoRhtcl/2x4ofZuNuaXUbWh6cNpwfgC
AuB3ZPxhJujoPExYniM1Mf249e+1oUMtXbVyG637fBEwjlCaN/LQp80foJz3xxQG
okjwQr5Q2ZkyBGOCAf+LWhDU712Fdxnhd1+IDZKM7L5vKS5fSRbPlV09OtORdJ6j
NEC7mCi7gP+MmUbZ9kVWVN+3bNaoqptb1H1BOPAR0buL9XJNZwgYkB7fj3KZtjqe
+zmV2eKuE04JIFKAoHb3N0WBMPLbbKBkvDDbMOhJAvsPT9KNO6BHFYCCQvLt+U7C
bsx3KlkCJ7e1S0yChqhY6Z8HzNbBW3gyOfAAqEmHQ6OF/0fQk5RdTvVnlYIwjAOL
2XLXO3jGi1ln6fQKjpriZHJ0H0fg9cvuGO4+Znf3H+FlOrsfdd2XJZWZGBJ/enON
7hauJec0N1uxkqRUjULr6DcZPatPgRG0Xu1kxMM/WS0imZ6iZ+W4I0oGE5qDc+Oh
gzMoWD/mKW1sE62S9ikgkc9HmvTU19um6yzGoGZjMiARtMvmsQm65FGa8mj4rIOt
LTwpdGRB4BvUA2j/sdeLcSbcMYafI1BEEpVLwkKaSwaE95WfvNgOVD+tM4LFiqu4
DIFhP8wLVa/rRTgaUycp9EWEx5vBRv6E8A+dP8kvmJKgm3MARDAVmVCJ2LTf8Joa
8UbQxQgXln3odmCjIoaT7zVnodsV7xsZ4tVDzIIziYiAW19F83QdM9kKLjBC+NWb
k5U7UIq/ApkO5IUqRz7jc1bmXw8U0FX5iCNM68wjiE5o+wv8Rn9Wz3DqKyUQpsC7
uAzzmipTt6EOLUu9YKDrefE12yT+eGnmPT0AYiMcbqclAAT8IplX0WDYXUtzTxpg
u4846GsEhXlU4aZk8QzQCBj9XKpBvczosg7EsVK2W7UcKwqIuNeB9zlZAgXW9KdE
3lSwQlWWNE98160E/k81qA/72ZksF3PcRpXuWtCF4qhRaxoS2+AiP3fpg7GfHx1S
KDm2xaTBSXT5CFnETz3xDNodJJApwr68KMHkic2Juvoy/fDxmkUItkUg/0GCW+5p
jHXtvqybmXg8hhbj9rLqzRLAQReZpTDJp2a/XCRRyedkyLEVoxV3YBD0u4XGcbJQ
HSMAA2nOuvFViWBdalQ3bdVe67P/AFDovfLb+TG3WbPDWjQdms13G8zlkmKoVrci
TnrOYRR4PrnzPqTHzJAxdv58hsNDaxkZCyLJwggBbrjroYYux9+uw7eLJUpK10qf
Rzr7MBvrmzSb5GoaQNX/icX7pkQuC63BFZXQasQsO2h5qYcDI7W6B+cneRfkWF43
8sEVFFxTtRcU8/eUMJjpCzyUqUwJWhCLGisOqqm5E1NlnLtDfmyyDPWmUemxHg8I
1H0+KbZ+2pqCSfHYpIIZ0WWaSdUijHANA+mgBaIzYkeJ1D3c/wn+MempF/fsVCFv
OmyWtUKxbztmr1jlZOsD9p6R1NtlBTB8sabkzsARzGDSZOJ36T0vzav4JaanRCT8
dk5q1OLiwxcloA4nWYZBgCf6ZSqls67+wZqht2xwMY/sL9KHPCk4P7Kt3DIzzTU8
SSBLsG8pfHX3vKcrzNpU1Nf61q8FGaC2+HFrbDoeSjMjBaivoLExltYhH5wQ9cy2
mxVgqNemV337gEPLZ24X4bCCsY22cX9zcTI7VPssJgPb9Jyx+Of7oig1pr60e3Do
GOX/SchhLqcbBjGi9oH8u4bFHS62Dlhwu284GqTqgN0GNxx0ZRgScnzWanrA5vcY
0GQOs6nUD54GlHVmpGnGFAcjXuJpR9HEgiU8qurrV/ab9z4K1SkrtgSmJbdRfA+B
aG2WFpnMWF46U5eA2CUFdlALVdk7nGgphquT791B0OXwOxrWxJx1NMV1sgTpB36x
aNhjuami4uHnv+YkfrtMzA0jKLyxepAA0GJBiBjx94JuI2K971yIHChdqLo6JEq7
QAsFdmimYHNwGVhC9fZ21Xd/lrh8H09A92icKKLSNJRA2PLA0qOnNll9w31DUp/J
YHc3jRJQYEhwLgVZWrCxTw6bpOioUbmg1lXNGcPwt84iu3QyUnGL6PbS2lbyDaOT
cXajBjexREZdVxla6wGDkCu7D1ia3g4cvsnghf09lQtBe/DKSzApDxbAKyS5UVBI
6gkWuIkpJIbguKBiE6pg0/MyAZS8IlKTQrsHc5l3LtlmvcOFEzrtNJzze0gh9i1E
0bEfaffLq0hVWa0aAe+jYjQV/Ai0Vguzq+InNeRKCN6uygystdIfVhzQi+iNTR92
/zB/tsoV6R909Kr7cKMQjIXYhybHZCIZ07gvrACvNGIN6VyOXavAsIbebmXSfuYU
ce/uaqylKmSnBMs4/wgbWc9XlC1fKGuNIGtQtFlUYiZGl9Y3ViWlByYpjZGnPAIw
5WVzvwkBK0cwcxFhKKGkc7pfrV2VVdbdxXCMDNb90Uvq9Ni5ec4eVK+o1YKlMczh
Ypu4K/PkN7aZ/+n3M8gCSB3DBTyb/zqfhLfkPz/hdxJu64oNemejmHmsgkzprnd3
IB3j4RtTsNtN4H/2ctEXrq2mU14z6tn4a5ZlhuI/CFVQViSho/H7FgERu4ROX54f
D1sulbXut3UIzUfcrDjXqHMcgrS9GubZT2UCOQGa168b/XWXFFWWYHCpGnWGFksv
rY/xGy4IySxsn88s2ILdbZ90N6ixnOEp3AA12UihGHNwXvEakRudSfUuVqP6AdPL
L4H5WhXEzK8RriA4FibkSZoQCiqTbTS6QXfPKj3kCus4o7YUveupeAFGEmFmLfTz
tVfZQo1z0aWULCRwHD62XQBBCkADOjqIzSpz+3YOD2PAhPdhj8x+KMKWd71asPAo
DnMrefbdwpQfUu1G5lyP50LzJjaf57ugaoGFSCWvmTSR5NX2uKSIeWX6ToigvgS+
9TvuxNixJNUs8X6palldVRUsgS3zTmeOWvgtSIVb1uJeSK0j1HIMBJJIoN6HzTcr
afL4PbQ5Bw5UQ+p1GJChOqCAT1UAuLmclewuchbB4wyqggaJBeJlOej9wGjMFt+w
BzkMQ9SbMHyKg4MMxgq6EEt1xf2wvacyOp7kvJ8i3lGF+TzmYOutrX6aWO79cTid
SskCaL3t58GfuZXfSG9XgotuxXY7xWVnZG+i9nWOfu8ah7p+Hka07MNQVC0B+Og7
paMB2lXA4GzZ7S2QxtC76TEeY4CPEjOptXb9/ALBuVTcXjRxgSk+Y6MF+7vOc+nt
M7WxPG6JBbs0/EqQ8fuelNMQT2XqLDNxzLglSjiLAGKzgfsVSuJNa762tOKbRJ3A
MypHfzaC6+0Psd8mVIvz6N6CcqjSrZUEaZmSc/P22UZMXSoUagj6gHoQLxS/ub+c
yezvwllns4zkrm6DB5EIMtfsnjbcjTGaQpCt7PQV8l+wv5SjalXRKVBtMW9YedpG
YnrI7X8L3wEgG7zcGRFU8MgDCwj0zROoyGivWgg8hMQrH9bfgFIC7HI9MLtylxTy
QZk0+o4jg871TigawbJQLS8vyLP6D6jMFBVJVA/J1AAJIgs36mjYm10OM9c5TVuu
18HHl6HSAwYxv8sPlyXkFrqhCSKR75lJYs4a/++UQv0bb9CDy4AjP/1Ocpt5y9Qo
moykehaZL+SJ2Yehn+ARBtqpe3MNuQZUAZMQ4yvDLsD9BWkYj0zvbSLMIltd8Bf5
9ve9CN3MgARyzLAl0zIe5ljhgpMZzbqfOz2TFcpmtIwlxQGXG4HynCB5lEu5UJCV
1N1WZ+O6HOyIk0CobvpAcc41Vxwk2ZJAbYwdgNxZhEc9JohaQ8ZwIYU0GwAcIdzD
jvgH6x7I/R1XPQHfpFPmTSsVprEN35Y1pLyCkoPUFG2YMiX/RBDUPIIiY5d/hv5T
KVoU1J/y98VpoOl9bH9g6LNaX8jEgZ++7Z8x0e/NgoGdds3s8S8byJ3C0eZPKZk0
9gtrkY0l6I+REFQPXADc1Q6DKP2tz+L8WPULWaH1tTPrtQA+UCfrs8KU8S8wrCAr
kPaWgdZG/U9pRdMU7lM0DHVNzWpRpy10BV/O6U23bhx2d9qgsDayeSfGWT29xe70
jZYK4Y2AOlc0ELjU2HwQO4NCc1N5GIX4gmXHK2msZNax0T0dWj8VCRa7FneUCJxI
ZYbkSAfHS+peo5pd7p2szcMQqBsF86ZrFN5ZE8zQD4H+VhOS41EIkXOvBCEqF3IZ
5Y1qrsAOmShTqyzj9WQGJIVRtKPqC2+O1cjchP0V//ptw66uZ+5wABuzpGJhEDsk
53uES5g/2BOgijupe7wR8neSeZ95ZXBJF1ZkJbDR+Ncsi5Hzs0oUIII5G1COHnFp
0bAPUdYNHdomlqZlrYKO0C0mNh7L5DL5IvA5zXxr0bYTfUT+jmga5eusq10Vpc2X
DHvDKpMIKV6i//UT53xWPLM2YjKXmaYa7rrd12VCgnL32U1C8uoGErUhTERd5TW3
se/PR5HFrD87JKNVmQYymZN88ZiKbFMnyxu2rJtNdMGgeuLK0xuTil4aQEPlFtG2
oO4jOTWQGmFKbI5LbmpYK1IipXtWEmYNcp1+bgn0m2vTvlhBR8vVlLweiVCrj1rR
5M15xU77hRP83CihLhBmXOJsPQd6WeJSl+5ATwVy6E+VdDUWL1WbUWR+KYJuyGtb
DHwG1NdpLEt7yNTOuVOeMox9hBlJwD5zE267+17Xmvtc/2MqKqwX4H7zwXi86NG5
Cx+adkdn0M3hZVednRsqm5aWhJJiKOhB+JLvc13YWQfmDAErqFFPFpnxVgBNpgJu
j2s6dlsZS7/IF+nkqVHbX9ohg8n4b91mVV3wxbQyCVLjKdNAn8pdFPfrjhfyrmwE
Txc6LahYqTbHZuBy7VihQJNB5SVjL3Nk+tAmqbYVF2ecVtugoweCatPnwf/zYbHe
HfxYcDi2iMaEI2bScnPlWZmxJ8VysmpF8NrjWUGhfCLSUCMIsP+MqFLXQd3gCHvd
VQtkSMr4ZFXlygfkvgsa9Ok0iIt3KNCU7rSfDDs7YLzKUWwRtz0jVRp4zDcLghSl
ueMpe7aTq5pJh2ou7zx7kw81q02SsuKJdCuRL6mORBxMj5n2RSyG2v3WupgwKp1s
/VRVnRMpyae/flDiVPLAQQo6MZyK4HGXCIcxF5JrDUzC4lpC8V589sMqSJ3+v/CP
IgB52JfNxrMfQAS1tP6NopDAZ2sf7kse87ejPhAPfVaalgbgJ0lKnZS1o/3quaGs
VFmgt1tZ8thMH5/qojb/vRrMNwgN7n+vvX3TtZhzanAY9Mpwp3GlLYBjVOlc3RAX
oNercwJNO8PMWXfJzdpjl7hTFowCOILK2HY2rAzdYL+p1aa9h8KFcVJzTN1ilHf9
2ialXeB8YbYPmNQ/9mBQPvSAF2WOS1Qfxhf9dYD6kIh0GTNh1Tb+Mi2hAndZKhyG
AvW+nmCLm/UUeMULI7btfXBl0Xnkz+h10DlxYVZiTnVGEoTbf++gLL5/auQZ4oJT
MSfzVKwkKpWvbgqEYaoW6msQuhdMxOetIxH/zoBwdIGzeahCoyjEiCwMN7GXlyqn
B7UrLmfUo1lSdaicIazqBlPhJ+YFgvsjRe3g5reo4b7DwaRD2DSGSL3UddzT5mhA
MRDpf9wlLRfv3/7z/MYHn+aQP+cuemZ4R7unPeZ8UoaSqsHcHzvwdSZuXWas2ivB
SR0Ft5eYm/W80B79FL2FeAHnPy3wjbkYG5n6oj2HGZKnEdA573DDE2e6IfK+x+Oh
8DPViMeCM8rOKPDSUEqK5Er7bcT694QLfWkjUGNEDVqSXNxSutUf+NLU57Bipgfc
Romnrtd0mvMTjaguX6iEhE9Zp9K0IveuvKGXyBfIoM/dJlsVi3HZ50R5TvO5LpGa
UZO6QQg1F+uuZafg3rULzVNpsZWPeerKk6wOtyCp1X+DpoOyYXqVG8UUx6rHLVoS
IZ9/jdwLkFRtxA68cNeWUXRujOeQhkigg7aC5Znz6sm0tbFw1SYZSxplH8EIMkLD
68QWVDUwmGQG+BGSVbmpF2o/FtHUvWhEeD3gbKR5V9BGk3LcqBZAxhgJKK0PRlY9
CWMeWRcCUo7614a2zmwrGJb+mhDTTt++SdNAD3ugJhbof0Zaxy9KZlwlFlMoNfna
muA5yJKkAjnO/JsToWUOuAcm7AySsirbWQiqiv6SZ0hxtqw74vLQeDEwDEvTYqGX
2KRjEIbAlh96usJ0t5skxrQYnj7+ksZsiHlRcN254t+PqbvDOw8YRyKs5yqWJm0F
NnYSBbAW6YVlxaJhlBaLqUc76Fmhao0wItiELEKLCpuMPy4r1skULO0gY04e9mcY
/q6WsegEM59K4F3jKegiZoI5fj6Sub/iaqV3XOBiViS46PbxxOQ9cBY2avgX2ymo
b74BVyQatKtRZ2ycsxvkO+FVtbFDlKM5K7slkTAiCFwJ+WgF5sOEPHMWY8JxENgw
Oo5RwbYn5T6enfOaVpmBYNzzh1UGMWmXR7XW1wTs4RmtdB6FwdSroB2m01JPS8Cp
Bl/DMiJJpY88fPCd1RBThuWtOHhGEVuzKZ7TKv+mHf21fZJRo7oeRHYK++foJ8hp
YbTUqVeJwEsbBb//er2hcjcopINIdI6GwC2jh66/HomEcIGWNtXffhkqIrokeSEu
yxiUdI/UTDSGwgvJPUisA8ekgVQxklK8sVkc942BYRKMp19iWpmXL1tI2hZh9BSz
pnhRWNBm6zeMdTIP5perIkOKDjleQh1DNXeHskzw6SIQ16wENOfMeKxpnDT1A/fU
+qpXD4eAa8XKReRO3+aPbsa+QfmFQ9EXblxm40kkig2cjiAAUrCqpRUFfuF5MFzV
oIlDb8C8nyIkS8uC/1vA5UuY/dJGodUqRU0R+zzbAS4aeCmO2WP7/m3anetqkp6j
9n3GvZHbZhsSFHAdqf5LVOBLmpBWSg9woCeVuobFL1BdRiMIIxMMZSbhw68VKkFy
DoqcHjcKuOU4kBog02oChIZTqREovJEy/NBUWPI4f6aZXScxvHftRXDqu7AZ24k4
d+yqP7qNRgB/3J+eN4PnhkQF5NdDPtLk3lF+4Y8eTXIJsDyZh3I8v+ZFZk3CQPf0
6lgZPQ8czCZk/v1S5NpZ3+C+vGh6oTkjebl9CupHTEo1qc7KqsOaaFB8enUQZydi
keCrMIQDEEM/DyALH6Eh5Ousw8Vm1nXCEZ6yhFX0SgsejA0nbWCRQnUAL+COEo64
NwZYodG/NwJ7C59dNwOL3kfHo3zU/ZXmNFsyazGYQH8MKpXfa1f/Bb7WWD3kBTL/
AoroESoRFbMok2NPr4hvhc18xkKLRxWXjcOyboQYEa9F5P+rNxH9Aeuf2KKm9Zg0
vbyzud8gqzDVG4J2muy41mMiJdRrEXTczMHHCARyDVoy3/ys7bg9oCzfXdg4P9ff
VpjfflXcEBn14wYvZHLDWUv7I674AQjvahNz8wM3BGJMVfR4vFSSRizMHaR55XO0
dnX2mupRy2/AtXcilPhb0SvdL2tfvFSJgA/Tdcf+81jx8qfdJpNHPAl4R0A2w+F3
C84FiEH5Du4dpK7aeEYQ5fR/32cqOT+TN2VZIr+v8wsW42Ax+uiG17nw1a/ReY8k
C79VndBQ0i4FuoN+Ea8iu63JKQMf20nBF2w+I7RDmihJrj94HDw/ZNNLic6Or7pl
tnXsf/RbsEWn2YtGAqo/y1BdUz3tHOz5j8W9ZPZWspTJlfgFmBEDVsATKdsPCowH
RA7brZSvsWq5y61tm57ivd3p/J/0Co63U1iH91b64G9RVo2fmSvjsycKvWqyWUqp
hFmYc4tUisF9+e8W+ppzWMJ8t4MSSvEzerweLFiXt0ULz73r72HGug9Pvo+l2RPy
iCeyn2xC9ip6h8nNk/ntf9EZ/FLmwC2pQ40EPuzeBLkXlvwWDeNuwwhj49oxLdYP
4SoGY7/r85bzq58GTCrWxONwMr13VqWXRbHNLBCbztxt5mZWT4pjOvBZGbTfrYig
p024OF7j1Wwi1T9lFGsKndjUj0VJpxM4V5cUfhu4TZXUmGCt8bNTIinEjtFRMzhE
9JCdLPVFyhnfX6HbSd3oVjI3BwRq91+CPTC6Ba/pd0KVz+Co/03RnRVDuwYcapds
JLI0kYKJzjgDVVvEeEqDDz+xfiTv8cFvM8+YDlePRik6xJ+BY5BRag1N0Qb50y9Q
0psLRaPtXv6kZ6yU36lgpnuB6+3BGnOCcnEj+ACcuo0nzZSzaBvOIcH+2NAY6h7A
DsY0gFUk/4/hz+4cE0sl0EZz5vHnlauxxaKlCa2ArtD1Qcpn23RFJ/MCCPM0IQxr
7+eaqFo5XjxvkM9IyxV/cIR6ELO7doUfbB3hMuhZ9HMQTME7UaYVzQ6kXz+ANlVk
SAyoDzVvyoTA7t11hVnXB3E9dbiwjgmCoo4FJHy6m+n6QEXcHjVyd7kyomfrK6uo
qYv61g3xzzYajnQMEexpFeeexIboPfeVlcmW1Zf5i01TXZNWPJd519iQhsuV4x88
CGt/FtAWjAEyexXEbTXd/mjMW0dkJeXD0O2gBb0sW8pySgICClj4nDbVSXD8OpLA
0OfTLg9zIQK/hyenxfrYqym2ZsjL7i2/OOZppUo2H17REYVBoYYfKZf3bRCBkwih
pccoS43RtXDqwIDe5yU0gFQWOKcU4XCE9mcs6u6aWlS8OxC2vuWQrXH22HZX4tRv
Id0eLTX28cfMfOW2qFRmRpgpRsRJwMI/zDNJRl3lE0JaB4W56u47hOn+G4GoORcV
bcxk3qsqFTgteKPlSfyzvHfyJLvRogfBbtQCy4TadnKyGA4YNtv4fURDRGPpf8+/
YK45oqCIN4RZb38YxGt89ykw2zNhwNMkWGRL9pfAmt7HUD0fq66SEcrXS7IhG7dp
wwZMyUOK91Yd2qvd5TFNCBPIqDSQZb3TtUbGG/q8nncntsrwEpkexqFRgVDiEaMV
cXr6pZBAMRcg3BnqFlT2KhKgiZPwE8xV4A2TfbkZ77M7wkC67c1mlGGxRqRzUPpd
Pz4TKCLe3WiTRqY/Lh5gtmyQ2Nm0e9anls2mxJJxp6sMARKsPAZqRGeUoSDRQSKF
+IcD3ymAIXvy105oC3lDD2odAUpkPNaVqQsX6rzSTJqH4A/2xltlK1rF3VVyrhUR
E7Tw9VHwpF45qABYH/udF2syvs3vmKl3fG/vgqfo3aRttMPnfwvbF73cpv+pr3s8
2urXQGuSI8ZWkLRoqcQ80qqpgrs98zgE5q+bdaQ06WBVgjcBP3iQNPJ3CHnjCRYg
1AbuFliWUfeqJ6ab+iMsWVNgF/a10qfIwPi4lXYBxJ59WK2kq1Ttxh5zGztFiDMm
UWuAnWrb9BqCfQtSti3Q93scORLj3s6hYsPSjpLNRAvYdh9Grq5lCOUJ3pR47ebH
3TXb70s5M+Z4FD9cSDpDUbFg8EJ0xJoM5zq7LXxWxD5vzZHDGc2y4jM6iBNhvB5j
atlU9dIWx5qPXQy1ZXXpzsxmS1Abj+AzX1gwrt6FX8fMM9AQZQEotW9PIpzO3XY6
RYhdzr4B9jRm8Hhxa+D/QXk9N3eYLSv+EIYqnDQSVqmm/OU/ElQIDwt0LHs/gbyW
6BwyAIx9xE7brbtXWXevEsVf+8BptIEb9GlADBW65zyB4oMEubyTKedglF1ENbip
6e7c5auByi/7CiBel82Jg4syqW/w5a63Ar3KNHF9RHYFmG8P0ozC0+4Lbwo5Db7U
OCjBPWvL/+ygiJ9c7ROQsFJSYle+RZAWy9bu5JGpjTegp5fUBliSbsSwjK0V3uTc
7dyeA4tk3NoTaekIVwzrdIHz2fWMqo+gV6E06Ul/DQI68Gw5TQvaXxMCSaPV/vCJ
ve2/5C5s2GjAgH4vPtmwOsjm4YdJx4IL0Zxi1fErUEM1TzxEO1snfIYeKuBLSG5z
EJFpBS6L3dO2QG2u+WK9TPVPD1/di9R4GkTxenH3Xmwqz39Rv01ukfsD6cDcoR7T
vpnB7lIFwLLH5Qgp7UYAGdFaKpixqmu64JIbTVFLihONGTnBdIrs66TyuSRKIXp1
Vnx4gdGWVyJowyJcCtyB6MAetr+vNES3BRiDdwL7Ez0wyGhWIu2Nwf0J7LYhwaZT
QdOOTHrnEdZOgczAqYHANYeZl4LGifnkcjWG87K1QR/2whmxMLSXa0Jm+Gb0Zyhp
0ObRoT0N8yuWfF7kFrcDzXfYILcjvFn1ZyEUNFaoiJyWrF0/A4EBU5fy42UAIT6j
oUiQYxC9ukX8SBAYZhHEqfhJ3MsvFyhPzDTG+uv9VvdaTCWL5u7W7zJo8+huMgUH
QtwiIJwi3rL53RqFf++yyKx4CGTqOdK+T76gai4zxHX8gFO95eG0zP+f92fxzn0e
MgKBRepH95NGqzjqYQN/XIV/YDE+0bt3P8X+w00EwdbSlgmF+KJTvvS98v0GQw52
SBW4f/bVMfNohvmA8kxtNi8pS8BlQSEjHcvvVgyXHMd0b/JrV6/66JKSzQxD1Gyu
lEcDNjf+hsXW5jV28qG5v5cbXnft6m3SSWRAH/GYUq1YBE+Fnk2RW/KbuS96VBYT
KN7zyYK+ZwNSWeorMbr+x64giTNDcyyJSNi+t6AEf0oTSPrOUmowDxB8FuKfDf7P
UDvNQVMPyJ9if+YHzEHgLccw9/UVpPLJ5JwjJyaVcKO1vo53lkIra+EscCF9gsX/
bfj0UszV352aLjbUUO7/h+vg3TPKR8LJrH0vwW5fo5sEK25suObDA+Hfw4reynV4
017x72K6K7ezLGp7ucXmFH3j1ouAM7K9uJuZGST63nnX4WZXUCa0rhoGMB5LiiY5
CqOmQroNauddcUSHA7QjAo1s22TGHyVdj3wEjWj1VEy2qoRZZcS0L+Tryz2KDC1j
uCVD2wccjHHwY7op8e0JCExm/Vv/l0h3G2UkqBnIzkgDU2AjjlMqbPUCw4kz0j6V
KQqm6kWRbPvAZdIwQu+QYhDyBIytmvjYXR03rRTTTiCg0Tzs7tavgwi+dw8NG8yN
5QIflIHETQA0q+j8c4Zhb2dJshHcXw5n3O4CeZGIm42JyBQcCYGM1e0pzestHbhV
N/joSyMXL6FWjje7xYqL7Lwh5M0BwUic+kDKqfr8W5hJpWLU0CVnNLQnJpP3dQ1M
9w1gWex2EU7C4pTgSYgAUBy6PwBgDoHuRNW8HGf1G62zKMkgxmVoEGgvQBCkebZ1
QztCu8empyGH4dCTkytVcW90HzHxVxFG5owspJVJm2U7ZYiyrCgQ+e3SPPInuBM1
t+RSsbKZc/35XKY3pEJ00w6efYbs4d8RZy7g6b6iPkit+cbp2TuDbqFNPH/4HP9W
sA41SccI5zkWNR/4ej40bEfqG2+QUddCt/wkH9lqGJ1MYm4wuEFoPv5rD8mhSIv9
bE8tfFLDeV3JL2TsonTkkKwcnn9ZTpFikUPT1ylBrFg1Hye0i0RnWOL4ZrcMTMyo
N995D+11LSZNwRjBBba+nWFFW45lewOeHrQyAaqkbgnt9OuWf3octsDQP6Y/9yRo
GcrfQx1hEXHMYdZHekyN1shA0+abVbODv05g8ndHEAK1uG7Nf6ntsEIfc6Gq08R9
VqLjT/2C7msaRy4RBno5F/vERLXWvlIB+HOipIieBd0Hy9C/zqGb9L0pjvCMc7/F
wRPGozBFzSMLvrfrhjjLtEglESpRoiKfXa8IQVH6RR/HrWMt/q5fXwAlKzjnzBFI
RgDFW5VQZ8c138Yh1lsfW/xXILFAVDL7Hm+MOLbR8y+Z2qzRbQKhNbBicQvclMYl
xnDssYw/FSGz7jLz0fNq/f6ZqzAEon6PgATbGOCSLbLTKbnqJHhRkZoWdghGIIIE
t0lbTI7+r99F22+n09kmVuVuzLUYPi5b06RldCslB5WgaY9FIK7UBj6S+CNyRMIW
pfGhgg2TqTRH7slchMwnAmdZZbB+NjWOB2h4fRcut/e+v3gdKvHqzvJmCHhuHh/1
h1HM3+FS/VelObEkL13d9cRSoEg3QXXr4wuCOGgpnJP9wQksjI5/cZx9gfzE9jDw
QcctybHO9sgwz00uPqSUNUDQE0/ipuznnWHEq/XKl4SmJwUG/WzWGOfSCkID+GPu
UXZdFp4DSPLHrb/oti2kvMV/zvcsPHGBYamSw/OmpUlxDp8vw5XtSdVENydh4CRw
nQGIoY9AGMUyKdjMkhMM5227Ea6qvbDaqm8vqJ/VSnrNrMa5H9YALGlYG1R5B20z
WwcREyzDWT2a+mRdppsv4IRz5kNpGuxlslJVwTdxmJBA7p9FKP9z0kI63RJfKaK0
UzqIlxSkI7fdoGuJ3/pzDl0Hhfw/CbpukDDBcYuOcOksLNno7ECF9231hU2uhht0
d4TzNZpcd3nw3sY5wZC+Y+nMQR5ZqE4fRyMawX3jz5QcjcLMCG09NleJpGuyNoCw
rwq7hDdnimSOYdck+SX63kVTyjE5PWfSAGUrTBrhG62kUDMnmzLUo0C/2oThcvV0
S/ImicsAGqK4tf5eGSDLs8GDiKg6kpycKuBpYvRjZRLRacsvCFaTrx6NcnHIRZdj
qPfp3X2CduRPZHl583iX/dDHQkXaqr0qK5IVJTzBcw+MPweZeXjmtMGenBfj9ZAX
7iYq9SOOvWTeBGpaGnsDrqRDxIe3KK41mOFWc5TCTup/RTsCVLn7I4sK0TLK7YA3
lSsBkxHjABTZOTMSve2vCMfNp4PIavGO7VESDP0UBkU1UVncosJdTLfUrNFKupOM
dPJ5d04Uun1498TCsV+HW78xagQz4fQbEIOVl478toU/7IGIImCYOvf9KiTEPbs+
S40j78J2qtqxEczJU8GUcZkj8cfeWIOOKwps7BNjmM9fDsNXomn4GxDW1o5aNuf6
pn7pZeDxvfkbU0RMomZGaskb9vKSsPZgwEv15HPXImBSctKtbYlxa5MgltRy4O4r
UR+8bDKH3W3hW6gs2jBo2PQc3lWqldzSckhrdXtT8elah9gUlWA84C1k9RfSrRJk
4INC/lwJhpYkbkLl5GFPkDxj+GI/ZPGSzwwB7sdNZvuO1KpC5I6//HXKs7XDvgo2
h8xmf+9cagWe69Oc/WIsvoM0XY2iFz2JmF9Oe8Ircylp6GkrMKwOMSRPBjPXh8Qg
qZI94JKAjjTIXmLnb67fjo9tP074zWw/OogdTYSCDk6jDAZUbEYEUWYZZOqa7ga7
7bhGHyf3gOfkVn+8Iq7cnxNkW5WSMeMuud5HjeHywnsZfFoQx6DwtEaLXgHRss/V
ikyd9E37t1ooDl52y9d0xQTbc+QJTyd/8RSt5+ZiE/z931VGo3sFvJTVyaByCMOz
HpAeRzbZeY4DosZdmIK83Ae3js6z+noHp/hvE55RVUwGU/VZs6F3Elz+WA+0/O9l
zDrobOOM+UEsRLB2SuPQh6Yo1yuXmu2AFcnWcgerlZiAUEjsEoOZ/vEgh/2WGWvH
HIgt5Mdtz0CAETj5R/nNQfPOAhKtfbWjbDF/+8CQ1bKtz6iMzmvl3zVp6E+G+AJa
QuUf+FgcowyDabwHXOZBVYnB9+PBiD+hulhrHrNeFNjZ+GWz6BK5Gwe4GALnWEyX
VwTolGXiuS9BT+S5+f39ClpeLr7iqDUTAr1SM5aVuFPoIwtWHyOG3udEb94+h+cR
BN6aM/A/TxsS4BkxnRs86xiALpGCRmFpjRAwXX97EQCKDKdGvItmDj3KoYoMfnEX
0wGzl179YIWwW8sMH9wyMR3KsaIOHelqHwfVgzHjUbVSltroEQQGPBQVrLH9eaRU
a3A+I9u6vMYqMdWdmRDY3trCGdlLo5XkCcHiDXDMaSypRxbWoyHJ2qCNT21lZQtt
tXJS72tCvO+WY9nFWH6oNk65bfpc/TRQGmnVwH5NQ3sI8OYOfXUNShRtzP6jqDkc
e0FkisTswu9DLc/HwNAaCqj2zTUC+1nn/Q7oTtV5lMijU+xHDL4wSRv44uyOl33Z
tR8+lyL1ue9eVv9yilYW6vVP5+XJxUuJ/icWKekWTnE+RaEiuA7ZFU498LWjSok+
MNB+hTUH40pNcw/zzDsH0Xd52oXbjNqqVEyfPNy+8zOR611SIzPhhzRRNjMb+PqL
zxWR1q9kCCjoh4zVw8y0IRpOBGOo8zADkXxEK3PmkA4wb8f8ipTcm8ir8aBXPyRU
gq7VBOQwKpaWsJ0h/pjqd+Wcptk2egdVBrqyNCvRthwbKCeXBFo+UKeTrXYPc/q5
ChhFNzVTfYQOVRI6nSnGFLQ65E9pbvSc9coJhlQVt2mI+EmgoLVkzxdrmYtH7SUA
0qA1PY3ciKFTwtzlp65CSUzqjUPRPYuIWiSRr6LkT6KqiS11A+YtQzGggYKbtj1m
N6+2etaY/6fQX/BY9yOSzUlokMYarmL+Aaz0SZb3Uv4G0YCuScJUQ47vD8waxHOj
T0nKQAitd97eZP+i8I5disY/pCh1r61HQci8ssyj/BCWLDG1kgrPtNu/KQKRzVa8
DwKwwkPsn8Y7ufalZ7zEFIVuDYF3mGHHMUMgMD8xsjHvhZLCi+j8iir0DKuVFboF
cRVlrvO5LcO0P6ICEVE5bgPZmZkjOGUMj9r+Ji0v+kV1FR3TBC0Fws7kN+K+cdS8
n4+64XfBfbCWkpAGfZwllbk4Uy7xt5d+qpCZqrggpH7EJDkruuUDhslT/QI9cCNC
RjGzeez912E+5ic14g6eXaUBkQT16XIibvU3bgwL9Crp+6rGbyQqPiMcj3BvBLLQ
vV2HZtiUMHEETkLlvzZrEC41jx0g6M+SDS5Fs3/TbgPm+KmmzF//Zs77ctcqHODr
C9Q9kQ9Jg8nDMQq0qlV4KkPXvgx85dcYcHMnkmARNxdhvmInix/BEY1i7JDmpehU
w7MsACYvZjNzPon6JWpInL62LkgBFNNCnFu0LzEi3uHqO2aya5ZxE1zpxE+bxfde
zQQ6PtsOf9WsCR+uC32TNG75El1FTu72bkDlUou+zdd6+SuIk/OzwESzq3SCfaFv
0o19QDjq8H8j856yejefsxKW4ocDcmDFA0D0erFD8W3UqFk4zg1v7tJ59yOSpXwA
0wlPnBiUoNh3WnFECeHzwxrAKUCpO0+GLPu35JWmnF3WrK6BMPj0kPqfOx1pERps
3nO8qVBirgyBahw8swfRmYsSdado9CMP4RH8IDITEgo+y5E1aqJWgXs31A/ws25F
pXylHB4BmMjgdTr9lTRXZ3tKF9rsqxdW8ioMA9ncqvnE/W+Dm/6EHpHRdQ79z8s9
1E2MGjiPX4ZcZja3Z48zcPyxz739i3iacZBqH51Z36gbYGFNtM5Mq5crYIDx9RKB
BMVkCHs3jC0xxMW9jqYFhb+sT47SC22kniEReltR7O7bjgJEyzaSM5N07qKKo3FY
B5Wn223AheC8qfg4NJyb4CluZzgWu+19b1TYXoOMAG+hf2BAlQ78gKjq7Zp0YtNu
tn0sjFqIBdzcPUcnLzn/8q5u9ZBqbSHHJBueHtameOcohnmCJsZXHuQZAr7HnPn/
O/+PGsNUXrzU19Dndb1cGnFhwVUz9FQv4RN/Y8XpYc3yAIZmxfWn2F6qiU8lZvOU
bW1ZJISgDP97mW7O57EqSgqMifExHcW0EkiAZbj5xtYKph8PYFPTRTmskQpbRUw8
zxoooRhKqka1vbS7YKJkPaXvaZnvVrIARpEcV8KztrGkAmzZgr0v/s1/Z2jqfpuT
WRmJzAF0rQ8QKSxJyT1apsRxTgVcyAL++8vsrKo5/nphxXpjKwkCT7ctTGcQ3FVh
4dD5lnVLzwS0KJPG/Q+Jn2rWOTGeweUUFIKHdG8jErgbseNuqhYcIgUWCOe8cIZX
z0wmcC0dj343z+A8oCkXjc0M7WGNxbtXu/hH0N8gMCkxw/DhjxMMD9LIUm5vvobb
ivWaSbPWddtDHk2CTICDY7rY4jTF0VJ1JavG14x/btv+LttI1mGjeyCZSy6WaTum
62u+mKAmTu9OmBSL1mMJkiXCRU0RHJN5G/BxdOS6kBuWremi9o9qH16iIjGTXPy8
YPSVGWs+Nj45jrx1p1qWFKrvr8IOVzFq/jDROqXIWS4qhUUPgAyG8YkS7E/oBZHX
VcgRLL2vQxZyoOWimneJG2nN+kpdN1/kMaeirFzzwistHcCAQYK18mO3pnLQ8FYA
dASfF+sd5EzFDZYHgC4UWWQ4SZ37JUS1iFouEWpbf2zma2qiw3GNBAxCFxc/e6Ig
cpp0iC1DF1xHdz8lK1ZNoWUVV1UT/LOsOPxYsPjFigAev81i/yaRacbi+y+1nz0q
ecG4n//IhK8a//LyTl7wfx1U1gI32xMfrW8APHDGLcoMCQVp14AHsNrGcmVhnKe7
ztPFY1h9CDc4LmMD9J0woit0GsUjN8Dqxgm+bCQNqTQuTn2lNgBCadtTjX0tZszv
8e1mMWyfNqLPO3FzPgAVz3C+TRxc7Bc3ruLHxeNq2ocCR690xLZdPvqLdkGYka0I
GhKYzPca2GFu+v3bAAPKQemyMLgA9quBTM/1WuX3BUZaS4+uSFNGxwAQ6Kw91a3A
6TlThCzpXaYJD/K82ZQIm4ctF0dmzUsx7SXOA1M+WQ10lohmonZeerOrdq5SvvgA
3vmxI5pJO5TzN7nPqCmoSaMkO1wz+9T5V6fW6NHcbQJEiRWgkgr1SMautY0DH96X
9IoVa7kgqX2HlZypcp+eDsrW/noDD72Pi3nyB9rpbt3OoErYJW7ar3qIT8blx/9U
Y8QDusMpDyTIsn7GJMb0j0AfebqolKXxAry7uVoCrGKaFEv4tZ4hDcCXmNqEHThq
OjUzd4/4vquGGzTXFCEUi3Vm9whBGZrxJpasYq59egM496Fxo/IaBkdTSaV1hikL
biNsqKhNvtoETHzdotBUFzgtYxs78uckV33sW3viuit+FzUHMZ00gDoq3xwAwkBk
Ffz+cozo+e0If2+xO6L5TfhvrbfPql2lLf07sRWZSlxPXNa+2YpulBq0MfcpEURa
Yrn7zW+lNrDCElPwzHs4dmVilToAFbqNOeWXKRSAzySNyg2Ue0BCLZyl60pCi5hZ
GN2Ni8LfaqJdCPJ0eqSla1xOWyQ5/hz64yXHi5erWth2VgxjqCPcfPD4xTG5ZXDT
TbV2uO9smTU5L7PRF2czMV0aqhuf9hxvZOuio25LmtwMS8THBw+tPRdVR3qBontJ
E9zVsHVwdmJ7Il5H8MPdH8Il/r9LOZAzIsZqjQ8U8kGNZX5c902DCMwlKD5CsGEO
FX6iEbkfdWwpTf2PVe1Xe44xrRLIHdOnB2FPKbKNCMlgiyaMTPhJAzspfgodkwrL
u5fOoUYA37fOLzEFLK9LH45QU2RICvI2bclgsWjSISBdfpwZQKkYT7W0P7HyBKtT
IQsiiik2Zao976x3NjjvQXj6kzAgrwMemxnarfcJtMIOkKnVDuVMqg0z/tKlQekv
2+As4NfJLcQ5ZjwYqZ5IKHu5Qj7BuanGj8a5XMyRFqpqdau5BzZk2RpqXlnqM22v
4iGGII1Ssr6B0GQsgVP7sYimmxkRqwJCtOQ/IarqgCCnvGg/JJ0W6fPzV2OfcRhR
engxFPg1RAmn+1ttvaNf42gEnpl8EqPa97IhksCxGvKGF8xy9AdBNAOqBEFc0KZe
ZWiUB+M1IIyN39qBqDD26QYsphvWgxYzEX8xPNibck+UG2rSUxVjJl3HoX5OC47v
sSz4Rvnx4mocDh+kQoL93xUQ5J451KD9xqA4yPup9cO6iBkXRp9y8yfsdd686PIN
7QhrLw1xe63dUgJ84yHuSoqM9boo+QfkVOeO1F3rH/PN6Pi7AqPYIehUu5VAZinb
8rWXgCcqRznjI46XHSPYGTJpKDueFYHy/Bzq4qXzNO5iVGU4tZjIbf8UWK0uar8a
qDTaK3Uhd67L1xDUN4c0pgVx1v/PzYgTyj0ROxVemKO+3nmTfv+sTMMxm+qxWivq
NFqQWTJpChiedjhus6X1Ph/oFi2yFKNa6QSB+56YNXLHtsf/p+Oiu2l/1ugxFY6K
l812LjDUHZvhnqYXChy7kVIuh/VZJSTGN3iOTyAwKGvHixa93FoS3le+Dza89tVo
tdQxCJyoUlF+MtiBO6XEMgmxuntu67/6GLdLS8SDSzj/3Ife8REjTFEFkGsqUkRy
z0tS/Ie1n1V5WkyOfiwhOZvyiBJDRK+x7ae/LzpI+zglMoDgNg31bOZ+VY5IulJs
49ltA+UGJd01L9mGc+6CAVBgZFR9/a5SrjI3tbTu9vvx0iRiLIIjgi1stYUvCuUr
K8A6o6HTF4WkPuTUw7QBzG1d0L8iRdQD34P0Ui+Vq0J/Kwp63AuIb491WDiZm0TB
XLuCEInxU7Cuztii2CO/QfxOlh+G+Ll1KNy5Abfkdk97kUXSIH12nltYLP454Sff
wqqaMy4v6UAgF9MmaPIKav0nhg9pzHoOXdwc8PiyWGUX/Z1qRFztSTecuwNR+lDG
4VnnOXilird2NR8EUp14BYiXRd/4f6JX+Xj6qhuWBcG0jb5DUdR+hMMppKTKBHSu
9Nwv2RRDDZLOzxGHQF/5A2qZdv/5c8H1AAKVBun8wV/LNXmtbG33VyfZLB82e9Qo
+hRRIIL6Ps6lRZWj1p5j/BqzDnqh0r8WytYWZ7zPukH9Eedh2SON/OgeqmGpPfJw
jobIQ44wdERUsB4oYZT3w5nCwJby63hCEVJTN8fVsvqUl7/Bxh9Lq9KrD01/bo2d
sb8aXf/xDwmF8d/6jx2T3SHU++NkJNHbXo2mCeLrtayKcIMsR5LfajFK3cdQhZPi
LPBgpwlf/sPzCROdwtGlEWh+BKiT0glHi27vckpYmmpXaJmY8i6vowXAJylWaxW2
F9+LOiiekK4BDIMvs6LNCMXwJWW1bDlZgbUHJ6RkcHX/qRX4UlO4YY6ik8FxCgDo
H1NIerfJg3ut+vqVIjlQmy2UjxfvdcNv9bMli9CIEzRGHK3/MU28SZ1jjp8LM7Xm
lXWgFhXTo5cf1NaNshuV4xAVrERa7Sy8wZGN+wMwH2CHowLEtDZDU98a5qioGC1i
seXxyIEzI/JDWUrZNe3BLRPgPdzDl7HHPVUPXMhZMtocvtc708pngolUwKuo8QO7
J+qB+rKR2AXeGpWpDn/ekynGvuGknm8k2Y3nS+tEpSI/AFn9f9ad8ImMZIZAU9AD
++mV8Xu6Drgi541udlX9d2fkF3+Yc+qVztPNr8d0pVurrQS6jdpmMegneSfxYYU/
aIsLiivBLipjEjbXl805ujop5fk8ZKRc7TU6fORdglsD93G6o59/rjgGFquAzGw5
latnkMFVtsnoLh0VnCSu4+NARLdf9Ww5sUgZqfWxCK3ZJ/boWJNqQosvyaNfMcvQ
Kp7mZkAOUNRTH20JVlbYOPi6tw0swBWEIBPJLCKGgbLD/3rYhJejfNXeqiWPDpmO
Xk/Kk4UwE58GMX8nq0vkqVuPNGz431vp3f/dWq23spfPco3rSl0B4GCv0VmPCE6v
nJvsT4ZRPDhFq7A3wiFv6WJa8igCIF+G6/RVKZ3grctaJ3FENwb3qqyAl5tvtSj3
2ljWhGfMD19yyK0d5g0v5/rGnNuVBVc46WrNehhg2LuhZrYYP0PFHZ7Zm+Yvbbs4
CBzSowGT9frq79gSUHjSij/XmwDTSIcqZ3q98KbQcJiepeKFtg+j+Z72lY5dIJdL
KIZQYQtfpNr2QEbDYC7Q/HqMIbA0OO5iz/OglIHIC2G+LoAHx30MuGdGkW8XrYJk
7YDXXxbL+SHhGXZ5KmoFsjvEYUpxTNj1jrs4nSv/mbv7dXkuR3ayvH1+g1DIi0h1
pNF9dRQ8fOMvhMFK7lTx6GPzD3MPsVShTfAgaAtZUv/vDiIlMPDFUgfrQtQ06D6w
MOaUwbsZD/CKtboC2hpCEsi6jGjXiYSeJj7LZxBl90Sr9LTKmv3/e6n5HUTDjrvE
wP95zHYAdZEM4dyb3xTsgqxXFWTvnlK1FMUPgLM1eZm+25oWL+JkVbQyqCAtg4mi
Py6kdLsdVj+ykS3pf7piNc3SHPWoZ54nhiZo2SUcJHFraQ7wfz36Qqd6Mp4REmfe
SenxYt92Be833OSrhN1nGjcS18/vS77IM7hz15Oi0uX8Ka8A9RpChfCiJDcig9c6
8X7y4S4Hk4LVbxCmEPqn0fhR4qmE2yuG5ILh1JsDH3OnCSzz5xt2kRAgQjJNePcc
sCDCVsVG1HfEKREAcSFKWbGZigsmF/qcYAETIYrutpOYUDMbDSkKEApcUvN7akcR
03Qajf6C8SF0WNWZZQm1jGfv4BJiI8REUwiiXLOzgehCOniemOWwpeyR9R/F6hwU
BmRREqpEQ6roQrz89vlMUrNcQHHFFFuWBvV7Fs/wkU4PReIeDTh2zPQAo43on+m7
WHFQbAexnkZSKX+OQnct/8h4vZoL3QbvKdGYtX5UhWFeeVyEFCA4d0QANuFwemHs
Ses8TFa5AaJ1aSvK3Tmlmama2O53LhtIGLOZDOdjRSLlQKwAUgRMTNRMr7OQcpF9
AR4TdZEFCV4nDKmW/JsE4ere3EJSNbJFrNK4hD2sY++fEgITl+kvsX5aBV63IpBo
VFHVcboIv4gfOaxe1bVTovTtCjJRpQm4IuRY+UTHWHJ8ivYAk8XFxuPhPTTlY91f
xbhR7qsr2VSZYAa5kP4Rb314sv81h/4mwU0Bc14lwbWfsK0RlwsiVlM0GXfkgGfl
w0fzb6Uve8u0gxHpTb8FQv3woMFgscE0J7BiSkHdZxD/w7kAOurtESH876e/Mt0P
QKtErIywCiL5XiLMPevz2fZ71Qbuxjmfat7RyZAnoHAHQvrtFtQdWgM0qC61xxvR
FHMQNwgSZBze4cVAMSJ2kK/xvDlAe5gFe49OaVlBLADBhCiUWGl8v1N/HzPGSa5H
dpLkT6QEKqd8Jc/RJLtlBv4Jcj/2R/yulV6bZEEwdFEFiomyKRV/vNWyXX48XqWX
DwsZEprxsdvOPKcg/JjjKf3sZ3V7NqHXBsJ9ipstnetR1zPYqxX6NSDT4G4IqT7A
XCy6KiIUB3LKQECTg52gOfrCLNii0TjU0QdHLtm27/w3fYillFi4j7po04mUw/u8
FDquER9duitTIR+tkG4L8Ft4Y4BsHPjDSz/4TbzErB0dcu7eBpSwZidCIgez/Vju
Oa15dOxo6aNDUGxEPWhYIu34WjNPhwHENFzb1huPn2tGwT/dbv8HYnT7h3VzjgX7
ug4kOkLjsiq+03cbFOmXP/rpRQlKyZPCFzWEU0R5/DTOqEz2dujqSMabXdAXH5lU
tJxJ8CNcsHM0tyBHodpURgiiwqokWt3Ffq1snIwRflMJK2qEnu3jDv/bvYAJztV9
hdQtUkuVUMYhGOG1agSpCfkoYY4hmBvjrAQlldDAoSMXSIF6DrOO/sepCLJPWWOb
EiN0AwMsudDgq1BOzO3xqY3wt6sHtwmPzn4NWa56859vrI8YUallTW8vKWknyiiA
1/mLJWf9rVe7ERTBvrpRIx7YoxcV70eeJDLcgmhL7QwOqoVDhYIeBAK5eM1jg5P9
Xaia+tITo46IBE0dvXUthQnTtbjIhD6I7kVfYd5EiiWPT5BTcxG1ps8FaydMkIp2
zS/vmZhqA8+G6x59ZmkKKHa1UOgfgenczssGBC+fMBQAetlqiYlwTyjEzfNYryQM
dTVxYX2hRv/8GnMH1svXpWDmsV3jy5v6Kbm1vtznhNfIZoQqneVS5fGlECLc3vey
DDUMKl4qRh8X39oRrmbJ2dUatwGjREZWs3is6SUvOcHrL5WD74yN/bgyoE07pJOI
Ml3Z4zefBc6gIuY0w2fWrr3xMBqIty17ZrAsaWJbQpDgBq/yFqbcccLe+xoiIC8x
vCWl08OdRg6ybJyammI0e0UFN9MObrzioyhdXWkaS8bmiDsOmEE7+jMt6iDaFZIL
MJ5CtSbdY/7oW3J1zGpGmRAKocmb/cHMwBcxGX4VnSuJO4OppI0Z0fg3URhJPoK2
Qhik/foXaLWK1vW2UckQyWwzVKJBwA1QCHDUXbWFKMNkSI+yZuOhYsw7j5jIhTTa
dtW15/9pF5dXuZ3zHZxM2yLPnOhQv3HyTgpYzWgrFgBBGcb0B6QbpXi3tRwqwott
AO9/CKuLU8NoR6lUGR8zmmYVpR/kV6RIhLEuC2IO4ezOY+NbmAwg41Ikt7nMJjvL
K8khesxhnT6JOqB80tMkADbFS19+o5FDCzB4o8noYbxk+iDYfOHKBDkP4ZsjxHmM
7U0055MoUbNmwv9bTCCqu11nO1bIpugQtqfznf5WRvDr294z4wMgf2FC+Kinwz8F
D+uKHRBxA1l9n18Nmm4dJxBeKU9vRQdIoEKEOAzpLBgPRUbsrYxsOdVv5FUMRcA2
D7K3CZwe5SKq8o9NP1zy8D/GAc3b3LnrnFSqNC2584pzO4/H6R5tMoseMU6/4ppi
gVVwi5wCLnK6K/HsVV36Vt5HywsDLlMadAB3YQoX3VyhN6/2cCNOj5VTidHtpmZ7
sv7DsdQ4ltPs8KbRmboHl7Q8m+mIB74P7gGl/2m5hM2oZ7s2WcDOkKLkGBkxT8cz
bA6xG+lNajrjTDAfbgwwg764iHRLYJVh7QXYTqw2owPaTAVPR0PUuMuvr+Bk+8vV
PysammuSfc8wJsQfUncC9YVRgbYCO8CxZn/PVyX6OpZIjkQ6CtJ5lHEM6Ije9vAq
/97tH7Rh6oAz8NDIahtGH9JcM2PnXvFSpwLTcr8UGdtkShoIGx3A/iGbXcDIV9qY
wGZ2JmO/HR5jtXtoTiOHPsgITGD1s+blCA41/VKS6jo7cCNshYJr5LQGYfdjeFYh
7aR7cwCursu0URelDzwnovSOX4nsRZDElZ/Z9fFa6+JRWAg5g0PfamSc3OIrOV4H
JVbSf4Iomsd0Hwj3TcLchHwpZqlO5IZlBYoaqYQ6wvQa5A5PnrIxSOOycRuv16ST
89Nn8CPy4SfJf4uwaNe8hQG3wFyjlSxoYGcMAHTT8TRNNPdaopefhYwRn+4MX5DD
YWkcOk/LZtqXLG2Qx3d3e/tOdfKoS8oa/IgUBcWOl5V7bXJNYBoOs1VLRBxsw9d+
yrjjmXJLkJ8EXDb57tYlgG6z5IhCuxQ3x6sTWDUhc8ghK1ko3rzY5ZtGTG/jZAeQ
gqlK/ik8e0XTDjv3iUQK3P7darUVkDgJoW8xcUx8AbJiG4tcsnKwDSpiqHXg8qqA
VrA7nIlZGY9quheKay3YVPgoH4BeWmDzlDRbM1Uy+fJDCYlrPgthsV2Vrfh1x4vM
Lp5AVJd9OEGAFo5FxCrm3eUxet4fhbohXkeI+LYD4QUK2FPGFPSLI9Nto/IGELcx
kJ7SwZWFR0awvf+3DaGBIxT+jp6ZXdeiLcc3tDSW1eJjIrY/YtJUY6dzYOExKvr+
hoGVqwaTKpImYabEHzZT0rVw+l3a55z9PnU+qeqMgEhc/Hsv2wd2CBGxS01OwB5M
s3GKtTDRVAU+FGD2E4aybIXxH72tWy/pxT+XIVa0Z0MlGlStGdJWCcitsSwPqEXJ
RhQ6ZWZFgQIEzAx9l3XJbnGQboU32gjqjZyZsE32OcAWvceEDpiNl8LpKgfivUm7
OQTejvHlaM1ROFHA/EFx6Yvu5M5Y9OvOxqUfSJCGywkuZfjCiyCrgDWJ9aQ/NLKK
sRMrAlt5qHGEL0xpsXDtEl8EV+H7PdVlMQ0y7xqRcEKVtqbPWANzTmJk0qnCbF7p
WMMwJfOlAhBG8Y01ugRfJ8PDA05RaD45BFjDwC5UCxjfYuLFQylROz9kEMp7cEnp
BCKOMojGxeUWvPox7fqI+VqxT1BLYWBbYc7lGTfx631QPuZODjjkErkELuvy4yAV
SllPDNzDmP4WZMhEPmwlo5x84V/+LhTPeA4jwTe34vMBwd1qSi3uwDnyYyj7u+6s
jC2mIJGYtFQWMP4uaHuMHai1uIsAxlXCsHuYfHIuWumVnOtVgVmXiMT4HmV6lC8x
1NNZ/xr9ZcFjz+3fx9ReD/HCID90fuHLsS8CaNVwxqiQbVIwlzOdXB68IVXXRKeZ
eltLBmAae5aSE99vCDRizESjPB9n9YaTz/40JNSWZrRgzfzCSG9l2tjJNogb5ngU
hEaAsYoU0tlj/7pTY1ITZrYOOrNmA1KAiDJnfDaHI3y986xJYgsRbDppmIKVSDg7
B8CqKAeYZMx5HjPgYNyJ3/jWjjxwsmCf07STOZIkY7CyN6mTlWYO3geZQ/HTr9yy
7duYM7M/mYOkIzeRyokOlDzJck8C72z9er/pTyoLdDNGfxBpWFBfEke29nE00ez0
r9PyZcN+d0mnMaUtZjhOKttb6ngeTY8J5ionKV80TwA+ePQoxAaNOQNRZGcvPzTk
ZJEYuk/EVAiGbChPxqDeaWr34jKXTYXP2gxTrROvrSqpi0xUawDeMqEbSgs5K/nl
xVF0fqQirTol/1fjVp1iXYxiw7tbXpKKMgrIKczU5S9M7PjMT7Zq/1J61BoI8AcN
XyyxcZx4lJ9ydbSpfdTrCEjhlENn5WL0hlEH39WreVFbQtUmPGsoTxOA2wAZtp0L
D/RrjayBxeKJ+qJnl1EsmfxZ5bqqTP4Ot4izXe1UKpGA7hCVAvZkyOI8GuC5Bdgu
9FVN8T8OIdn8S5rdy4nzD46TcIH5+Wzk6jv9CjQHhOQT1qDBdAFgnslhf59UxxXw
2StroGgqsCLtD20Z0uLrodFnZ/H4Qmcpyla5eapwUdf7tcteszSLwC+e52T2SM1o
ESNMpt5xw0MX6Z15VZoETmH/iGD1PJ2k4mJeO3XsY4yeMfECrcjJUCse5q4SVBB5
3e0KbIVuGdEMaxMnrcTknHd8siW/7qBsfrmRKSkqsgaXgKSkfFz4ktiBfk/yVic6
pq9GV8X8VTmCMiuhdYsXZMXWdH5a/xZFyKgxWqoMGHHuAuUBbv+bPOUFIftOgq3i
xL7XojGbwLQ/Bp6J5U0xLpj6Z0dYu+ibKsqlSt1JGWL0zHT5b1TwMSdEtsZDS6sA
y1/97aQpMtUEe0wn6Egt5Eito5uWKx7GAveYXeJCVNlIaH0cMvICmWbg0zycBSNC
AK/rnDCtXK5KRKLaNQuss1blacs53GTBzf4pQ6n/xLnaoKraKK6cIkRiIgAO67G2
6+pNogQBbnPzfDluXatpEBoV7SvZxchjj8k730yXkbeelL/Ftr7zCAWCGFo+PI6+
tJ1aXRW++yFB2r+yYK55io0JWUdVEknY0Z24b8Sd/Y/mnZHa571WeKqtVmlEivBa
3MZl2MhIiK/8b8lJDA/1eH+Krjtkoe3uIBehW3SLh007PNC4uzNpTmuIRCbh1zoC
pPOjsKAn28QvqfKHyJJlW97IsVN5niVP37x0ixIJaV1iTNUgXhER+AxFk75Gr8Qd
v+5T9obCj8K8aAM7cCmIT2TllmEcKIfuaaLtPiVxbsA9ie7khr2WKGZTjW4QlBts
Ak42C8/VjKu+MNfelwbEYtUZ0+N10KdEk3VMrBl/F4EXONfdXe/tqOGFsTQ782Pd
han0hctQlADxTwgXM3mdWh+diF+cc9mjevtw5dYKrX2EfW8ZH25i84jstZV5fDMX
h/OsRuwJhECODeEsKf4+Y9yvFIUx63/JBpCdWKuM/bcwMjxEroHMDplMbSzIbXny
H6utbtqVPf64Y0XBsNy7maHWiIvy6ne/iN/9ILypfZMRYsjvDhcE1oaUQc6xVKIq
x+TO5vU+VWzYMOgS0Do07+FxO2iq0YGGq403X3YZjMMsT4WSayAMNrlPX0WjIPE7
K3/ALkZ7FeAEIsA9b1+cD5YlODl5MRGog2PWIqTMCxTIOcH7lgSbXPRNsICsAhmH
jX8RnXvxkW17HdZ/m7WGs1fPjIbSvPmA29z2wNfhVD59NCrUSE6Qqsf/B2eYnOdJ
otIJe05E6MCKGKx3KDbMCPOr7JQw+uMiw2zz/UI6zmQfv4ImfQqQJfhBKTEmZX9F
2wpjImhRLlt5da3v6armfhx+XFVjUYiiX2bsBynu/mcyPSW/jRXC7m6jZLSWGG9q
wvJdUPDNxwmeE+PTzyIVzDuOIoU62xaCuSYrlKamLeN3S1iUmlheZbpQvqfoqEL7
hMVLTgNnnOxPBVibhqnd88zMBKSIaVm/KitVXa62GMVXwdAnTXrbAEVFhiynoR7G
LYAjXWuOxdO+p5wrZeN6UuGSk7TTA5zlxx0xA7DUZM7bCmrMpWiPnuJWCr4R4XFx
mF549/gtCTAToNRETCdhdf5YqKQA0Z7QguykPS1SSoDQJDjYBKjNYzBgpD6KTdB1
TTc8xFy/SS+7+UK8FdoLEPCU4lYgs3aJ5rDQON8n4hGEtvORLvFPdpvg96mmdhCQ
9BU0/2ISsQvAa3w8xv5ADG9Q1um2Plu8LW3Rv42D5/ph0fTkORgAzhsLMZF1Pfzt
04M/5sjCSqflNJMD20qClYY9i+BTlPxAWjbwK3y/c6IZ9+F7bAXttI129/u2MJo5
nyriWC/wezAbHBQVX0sQRUv4WtiIfZbgBEWcBgmNYyNqE6Ix0pz/4Klc1N14Oqw5
2cLdyqXf/OCcscUKxBNpgaIr4irOaEYwvAyxZF306ci60uVLFTWguPwec51XvjqS
6Yg0fDDMK0L6GRNQtrF2oAZfSF2f1Msz+6t6f+YTNaTxVJaRp5S2+VlaBCos6v7P
0PmBNc9gz4YCW1jr02k3KsmdPceyoZslCQ1hW63iHaS1kyFeqQ0Jv/UNeqn2QSaB
rgvVsPxMenIjkH6U77aSsbCDU2mXUC9QXAZ7rg5RAZkZJ1BsTurYJ2igIKFoq9H0
GYkK4wWnKBIgZAguPwl0cAVbocdh9orK5k8hyBGAOfJwXO+CgeDK/pPvvKTYtPOG
o8ZvjUDDheeH2lePQzK1b8eEky17TPa3w6L5KDQwscemaIldaxQ4+4KBiVzFwFtP
TYrsuymqqaEyDzQOljI+xJMewaTFBSobkAjKgzAcCgU7LKNt88tZcDs3YKbrCO1I
hSGW2hHVyESJJ2CHULEk5wdzFL6KgYGQKQ9r1/+VhqnYY0is6M/GLpEsUKj145ai
cb1I1TNYxFo+skHDnkytyILeFUbR0S0JhLeAithiWUYvoQYyf4qKlzba3QG7ec9E
xEt4yJTQVPfSNQhyUvqT61NdmiwnybWoMCW+YoVkFGrUOAQ+eGrMBdl5WmjGNRev
OzTXmCAFYJ4C+ZCUgEMGnkVxkBLkKIzGiDwN/LfBwBPhe4kbOeR7JpgjzYcdAMWe
MhQ9r19uh+vh359Rox7HemtB+0MmBAJJqzbgBub2FzCElhT8MIQb1AD0ccpssN0A
QyJ6+hNoTUBnzNWeSn3dybeYulfPbZWRgPPREEhNLwMb8N/80B5v/WGMd3Nx5oZp
tylNoTH2MeEdSmA123EaYpp3v78GIVAz4dZgJ9enYiSnxgU131dV7al0BJmJNGuw
Na5veLC6FZM+8181Z4IQK4XbkfwPc/3MH1616ULWpthsLEEAe7fN+ar7af9MYx2v
qiEILYLiGsLitcWblti/t2MOEEZIdMotFz06dwTA4OZghitLJd8fSwbdgGK4+Rm2
Zl0/uNn0VJy+7xj1JubKpbnpm74eOOp+3Oahi0MU3v+2udZCMpjRLdw1JxcZngt8
O3BxB2U9avWvfkRG43etbQRoR0jC1ddrv+KJZ7Wo0wQbmBzzrSxyZfJiY3SbfwYQ
cberUJEztwf8mtK0Z2Y93xBq5UcM7DjxzZ2XcEM4z6fGvSxbXQuUjznxJucv65UK
ybgBCmo6yBuVJgD5tbpnznpjn8Vi0EAPw9BjbtQAg4ej2UA9bPbLk+QlhnsZauUH
8SfwEDCEkv0r3HpTpt5yeunoapmE0/tcuVQj/T9D4zI2aQbPawpr0jS7D+36d1yG
XQ1l7kAEu4KIUfs+YEX7Qpvg/5CBSr1mA2/0yobuVh9ZvWfo1lul+lIWMncTjRcf
f5Pq8jjfmE0KqwRn59HZd3OWRWAsz+0FgZHBwd1+jFtmsbpxs512p6XByatXp+MT
hTlZh5G1IXKWDFY345v+/r3tUVDI1StmB80o9KKzJxH/DSK04ZfwHlr+qQbzh6LD
/L/iHHRYrA/mlbbfkQ9OqkIfv4Ku4Vs9JH9y9OyEpKsIwmvXrT9xT7IGTBtDQYrJ
7k2cpPHGA3IWwIkUiTAdjIjiP3iUeLLvQNan04weWKEboHasEE9HoHMKBXQrTBjp
skziHIRPTxs0AtoXDLKFfci9pL6L7r/7rYR7xHQHWzexBJ64fGH9zs/RQwadN/ns
Uk6AXQINWb+jIjvt6mNckPD3yTI8qdg483fzFTUdDWy+b+Kbmy0PYXAKSFAK/3uz
mfK82BrY9JeLOnek6FD55tKYVeTAZTvBvMwHCPus50J4/zd+ND7upkQuSqtaTizU
/Q54x1MWMf6Ex4yfMmyoCGvakPE+rdlKKC+ut8zsvVMjPxXm/N9lEwYziUbnIv0v
PbZuVkU1VltsWVILwTWipxc50JdpXtXY7nqaVNsu0K2dh/P90MjcBIOXThQ2r02i
8/bmgCQL4oxphoS/1O/0nDLOVXoO/8xjBpR+78EZuBOh4T+pP4kIl5gPtVIPAG7P
47b/5wxaCFVNoEebX+5X1S9LRk9hOEKOr+NXa0yrPKruvWNXCuuPvlVK+H/eIpGE
L8t81QM2z0ugSOdsvM54lQd9NdeQa3KB/KRmgcLFDyuom7FqnKxaFzOAlSeb8SwE
IS10E33X6I+IU6hB5QZMYwHQh7W3xaCD3D5tk3pSmNLTAFlbYbj6rI1FKwRlfmpy
vhM7XTqlQEmP469UXOxv+zebawDHeVULfvvpqY+SKiAqXDzRFnIchtRVCva1l5uv
6YzEVofNUIraGUPHp1bWGFnAAW1X6YjHS2g3i3Er2L4xbvt/Yxwi1gvxw6iXZWAv
HCd+Nzv6TvpsyGkkcUnoMUbUbS375ruKei+agWenqN4DsiTkXflIsvQGWFtzgLte
h2A+WTOn5sPkCznXsaAa70qoSpLRenK129sxLdXIZuXKsXpWmchdpNyEQI2kx0SF
FzoGJniwP07vkrWezGhUkc6TS33cROsEiZI3frelU/nnOFEi56/2HSCrkaK1pjsd
FOIqBxk1/ivI/E+RaiANrvcnNBKxo3cXRSbvE2xdfNetOYkhGS+jusKYYqpo22/Q
jqEbOsm4SWvaG7lL6lTf1xmvDm2E53jexHFHnrp4bQki4dRnJzljQJ/IW2Sw+LGR
7MWGKfKnrTVJcTFCEDHLLxnbJhyi1grZ6i7RabvFgkWi8+t60jEy9no4aiYIhalf
OREfnr0ARyXC7NGIr+6yksbzBRHOlaadtTA5fxb8+/3XdF8Y0yXEVZXWsI2DBikt
m/I0NB5s6/PONO7dE/hj2abB6uh6vCnIHmaI6tZlg3IjNJ4iTeOoLFKPG7AcWiqp
Wf8GR6G+vR6t5QISIufbr0WWaGzl3WBw5+KZKadIR+bHozKypM0rGKrA8z3dscGV
h0HDexSLASXjUWrzVB/n1HW/in6r3NtK2ttBjKrK7pYXXM5x9lF4+Wj1fQ4HM3RG
wwdtGmSLwE9ZPCIFRDaLVbx6kE3O7DnhDc4viUdobd4yCSiRFdxGUCK04N84uzAC
kSWKzFaybZohAhdPJHn1iSNRrk8skSnUynikOc1P/LPkmv7xpoMa3TF/8zQqSkcr
RqPzoLBqvO/gpBcGqVoq4HFXOglMIE6Chr0g94uTdbKHaJrHJobB2flvykRmH1BH
w9mQMBWu0iaaVrhbynLAD1ljgQ+o55XfLRmvDOKO0eA0Wg1gtxX8VRh3TEpwYFf+
FAC7MtXh+ujs9pnqTzzf8o2zwP+PN6VH/xLc0qUfTDvXkfjqn2ijUqMx5ib/ykxR
e/Hvu76+AM+55b2EGcvj8aEWWPEfcN1Svn+fQSskUh2gvlAjKeu6We8kK+qwr//l
NKrOKpoTzITsy5p1MmcY20jcEIT63ioCeaX4tIGgBB0+U/2LdZsPXPQSd+Wk/rXK
cgvdBSwtZLP9ebnm8zCrbXsH1IDZK1gEnLeh+3WpdUFJtIUo4CNOvWw/lWNGvXif
TDnI7PlfWmmLkwC+88ZlMUAKTjry6kv5ChgjrIpbLa4Vq0dAR96dwwdE0X1hs/v8
kusonsIIVUTh7KmXVXX92jmMJIv9ynaap7pq5aJe3lhidl3+a348vHf4wTxPEJX7
4sLxUdeoDDc7NLnIgqlW5X30yOdQYyH37IFG9Yu623SKzyJcw9Ik9uPaJ7cIQOmW
EVZ4Bew9dRX9V6TwQzZywpOVEGcJAxih3Q+tCg4tYIcv8gygS4mXabzFet3JFShx
hs8sJtYgKE6PfmSGZVKF82NVWN6CuxzIBNT7FHzrUCj4XmQArFZzd1HZDdMd49IM
w9h0BrZzmX6vsNZB1HoTqJxUcQdYT1Q+y9xpXVl4oPH/AHHoVShInq6CMQO2Uc92
lj3kpZMhAark3uBkIQ7yHDYVCLaYx2NhoXuM4x7J5eiEQXBO1JwQ55vxWjEsI8as
lND0NzzGo++OOxpUPjzQOOsO8edrYmL3hkLxv70cq4QnyEoe/bL6h6Je4SPRUgRy
rW5dWMugxkJ9SCPlHhpQmt+ezHzsGvV9HLyHYG3ABFfL1EyNYg69fTFD7GqTB1df
d/1Q1ERDXajUMtkHLL6C1Ge5zAdl9f6TUhvO0dh9+CLm9FmynbWPpea+asykU4c+
/zYMVCX0SXOKVhJA4vEtHxGfVvp4pqVyA+vXT1rmWCZ16Ru0drw1xav9qzkNTJQD
e+O+FKHIEyY+AtIcePE4LzJlCweqh9bLsau7YtGY+qx7ypc2/B8YsFBr7NgIMJnO
EQYtmoy4IClFiw9v27Kk5MiF+xWM2Mcqc21reGcEib7PMPjSLPKUnSOTuLzd4UO0
61pHH55tzaULgWvuCF1cPobywZcVThd+ECk3tfa0j/PVzPj/AjVlvxps65xxD7H+
emkwcYqLE01wUuWsO2uv8HyBA1zz74KhqtTubvMuwwnn93i6lEV/jgoIv1pUVJYv
t64tykkgSfSKKvzMTQ2u3shDIiST6RWlALT2EFhCq+Zyfz+sdP7Iv/3jk6ojhkKA
qxEIJsK4E7UrdLF4Ssr/ii8zy3rrDGIlOB6eV5ZH7H9pz6wqQoKmYnlRUWpFXrWC
/jYumWEMheE/3tQBBUyQiRoswZVlAvtp1IdmDxyhzpm58IOseo41DT20Y+jHRqdA
TSexOpPOqCiMKW0pIw9EBk3Uz+X++GiOu0onJmKAml1haLHxiXmvhAmuu7LI9Bgd
`pragma protect end_protected
