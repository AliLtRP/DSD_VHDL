// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mF0uO8o/JuXt6imH1za/afH83ninzpGdQBLE/niKpYdsXVQI3AbVC4RXd3v86qLf
LT8RaLLnHGLpOM5/t+pmJUAmy5BpNi1c7QSWos1C5Wu1Dh4NaQ9G+SdM3gsCPwFx
9gZxkCfCvRJOhJ2xUALmjpvaIe8qRB91yxZYPT9ASQY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14336)
V4u6X7TQdkSW3jraRIx0ZDQAYIq7l5TBabZpzjQoyNCBKgD6QJ7AGTVKtRME478P
kb0S2zw3zZuXtQQf2dGpdElF5Zx97glvLj8Bqyib883gYO/949aj677vNXli+oU1
wCz7GfeLKRJM1KN3D7M+dIjbSzHCNGR8LkSDLsBT0gGf+lmwbRLqtI/aSyLGK7Th
U9iEzw6DF4Y4qeo6YdvePNcJAW1+pnTL1SD6RyIMBJvw02uxsMf1eN23zScQ1Ho6
CRZwxf+PvMVUN2TnG7PdccdMGPiQFLViB4MMt89jfvdCGry2onWfBgFFfYo3iYc4
YNVcIMlzfCszkCqFkO06MykILklRETW4gEUrRfpjWPRGqRkoolbVPXFRjD6u78Ph
qEvuQ0oZ7UrIml1FI4GQXPkIdmZ28ZxRyayPSzH5BcwwHNVrWF2I6NaBJHX8Ch5V
1pR/AbmZs20z/wTCb7GTCPf5hqcJDjOAb7l2flIc7PeyiZ7/ssdsv8rCEeuoLp7Z
NK55EJXzSOTKfxhxC7YeXSIYtDO5/JV+AHGDJpMkk1eVOFJ2wwXFGHLZtkl0YLrh
LMPmpOdx3Y7eFgVj8qf6p84vjGXVkVCxrjanSnnJzsweXialChDOIG+xEI45jOjR
rmZGc0Bcw7W9iXsIXMpWOBbXGqTyQuOPuk7u8hmAODGVU68ftWy2RR8DRw4ICg9G
R30tFrsWLLBXmtu0+uDUyvYjTWQaUkVa6tZuG50INj2wQ1RqlZlyNWlUgMHXWb6H
BaMCe2d/ydHouCWaf8KKF7ozk5xxfbJ/hGiv5Ghi3QlKqb6uu7sWgUcFrIzmptku
vByisLA0v0QNpnsErvMSf21KEO4QE7/4vIh9rZEOh1ErCMyVfM4o09OuJN1HaYb7
pBkICaJtiv5yWOByGg8v8neI8kD3A/3CFlqniUmB31b4G37yXMWq4VvGNZ8lxzqZ
8DZze1pFoDQZqDRrVwMpTXYMCnxgf6TkqHFEuWiTuU+TevwLQ9tFpeqx+cL6mlBL
oktdaACobAQUjJ/yJgL3g++8ylk7i5Y6wVKcANM0g2Y1vJ2/YIntpYMSgVA4u96L
RZViT8zfnx7rn0wf+fpiFeFfSSZU+WklO+M5i5eFzisDczOfCijymf8KU8UB4Iu8
06uV2bFqsZj0oY/cwoEU9Pa6WpG7c6vnCs80WGDJjSt8tbtPFebbksTbcKcvpMAC
rVOhqQpGadOCfOhMywLNF1yQypp1o1y4ucz7qxp42cVtfuG93kqrG45m2XN9+yhe
QanCmQ4cX/r7+75HQPtMf1zzpvb9MkVxIs1wLCsMgQD6vclL9ELBpDc6O6Iinbc7
Ngp4lHpp+i8XOV8uOtkjIkSFmdWj3y/1heJTh7MoBQtC1KGtQLxxkMjei4Z8/W5N
AsVP0p7od97vP92wyVPWpjXBm64jt+0Edwa3ViyJVViLCrwqnhpisZlSuu//Vtq9
9KBvlTSQP7oQE0FB3j1I5J1AG3z+oR5Lve4DRQueWWE1SGveyu+R35jrK0sHHCJW
CoG93gLezHc0bY8j20q8wE2qtdtFvMXO6d/IkqoBQNpzQqXwHRXHZakgCRqWlB/p
hMSqhQ9JhNZmh2CtPBQ0ZMgyaMl907H/XAlz7IQIlkAbzSPmebW9FZCPw8hjZMVw
uRlbiQv2g/jfrpdxr+DQB47PuA8iwCwHXZ/Ga7gDUeqW9vc7EJlkF19lj3uO4U55
8wnJkmbRDWwvQyzZSTjPWRM5BQ40ZAwYUPIz0fSnet9d0pwnLXo0dDTvVGrAdVDx
kT7AkGbucZritj3R4fM8BTBIcR4KoBLwTITQe0EYGkvHAruHzVynEtmpcAcAaBxT
dtU0ygtLFXBygC5GGvxJvU1MdAXra2Le/MtV/J7hY4KdJ1zIYYfqcrgxjS4FAk0d
m+TOvuLoKrC/j27/cklvWXdNbqxmJl4AkWcPPWtMedLMwwTqnhFA6hVkd+sB3mfB
B4twtR86JyxZN486iF7W56WM03osXmJKHkw/hKxTvy7i+SVvS8bdKsjZkuAycN90
q18/n3O4Q6hdtHTtWW4npjjvy30YqBCH9f8PI6BUDBejla597mWounxT9R/A12Xu
Uhr94N184rIir9uxuuGCjlOE5OaqxbbQXCKUVerO8p6WyQQpzXu6jpKw9Pujb4a9
VBP+e5vCiLxD37X3GZCOqamJPel8hefyBTJmmWu2/eZa6JWCzp/U+FdoFlAndlb+
BpJWNXymckRMOJeSrVf610CrP6N0u+aweMc6HjdzaNsn+0qSRyp/oCDj4YzBDIRb
mwCxaKkctOmdKpvOEbfEB0WftsZ6Qa/X5eGHGTeh7e0U43mNJEMh4xIFIx2R2CDI
DQHc9/RlgC32JvLXDjL1qVTxiRyYqjWetAw9d14nbfwQvkzuN+f0daTrW8KtxcMe
OuuEp32w0jEygYGfnrNKWHfdXNhr43TOW2bLjY5kgN41JQp5YNZXGM9KiaxZRuEu
9twnFgqW4yy2fxJiwW84ExTB+tUtgRrCocig2M0Oirmv+EUcW8SsBhIsnnk+fLyH
zkmPj9hwj4kFLrQHB9mmvRTvKw2usrf07Gy9IewPf/b2WZr2IeQYJW4mk2TYW1Sl
U3xXgcl2M1Ii23aw7uZdW6KcnZgC8Y4Gu1N5rcjzdwH1UgBWYJzHmcVHUyJnaAgh
nsvrygijq5k7w78V8UbHAYXQsq/jIL5qPLo5wy6MXu/+sOE/yHqorUKH8TX76fBq
ltBsvXEYeqWpLKdd4eMWidmsLKrAs+BIM97s6GvagSHCquYx5G2Gi9CFSsgL4mVw
i1pi5NpfOUmBMcXh99Vrktu4N3zr5jpXf65tysONn3ReP6CtGOQOHV1m/g58TlT+
VUtWkoMmHddd8thUT0mNsNQaouYGllNdpZCJIkzPSzRB1zntESBk7glZvy1NFnHo
e8mWi7G9OVwFWuAxfaAJbpbw4wL5RE+9Uh6OQzoUKfXc6+EzS0A5ThhF61x0aCPT
7JjZn/TTReSYsZYKtS3lv7Io7h/ENprs28+VnkFBtfRWJiyNEBFCir3pIOJw80BK
6GSJc8UiDzoJRjgyLaRkkO49yPkXi6aiV9fFT5gazLHua9KxVmYWdLaV35ZL0VaI
hvBEj1CNuEApUqAMIFveYYLsQazXEpfPnt8ybVL9bkI1OcM4J57bfwBBEQaq5U6E
N2FmqHhDmtkrWLwD3X84B7pwcY7cG2LCYSIjt0STnhoT96ox6v5Yhuwt43UYB2d9
dFKSptpKSCaMg8cce3g8GzaQE/xIvu9us8dOihrW64zIewDHxlJlg6C44fm9EuuH
8lBauY0Ymc6EC+pp/kd0CQojJYYVk2koc41+xdqlSo1HhyFJIFQWIkVnGhGPWRhZ
CHcWQ2IhBbt7oRIPgYnwPFHxOngETx4KyR4hFVtuIlKYzJpKuRExMWrN7ReaFQvm
99OL8zfwPpA9xU9smzUA36XgSkutjD8Lb1i1swQPc5/lyOhWkR3iKcA1HdoK28+3
InH++GkQQRXoe0kxwawRcSKcriuja0XngOcIIVD+ETWsDofIAbjMtylIUyNfQAqp
voiJ3YqUsOr4EL7Eu0M2Xz5Ddyg+nnQjgyDu65I5zBKxYhMsCgLzEn+SiKLaYAWP
6C8fQwAuMHzxKNZadx3BeBgJFaKJBIp0SnrkKPip9kKOeL5OVLRykk8xcGQE+bcD
do+MFNCsGtv9cZnMEFDTb1EsZnZ5ejhRk6GL+ZQehdtRWfCEq3AM8ZeQDgbub/u5
RxtkELtKRUzj/f8hdqhNRL7Hx+2GvskZKoa12eio3/uGrK+C5mez1ZyNdT/r3ijS
6Z5goCXPwh6R1h7SiRVaxkD1EuNDzQMeh3FBptJBOxXtJTTkISzU5JksJtLGfX1F
q/rXOD2HmgeijCuGSm8xBVYKrobPrHbP2SwSe7gDV6CvRxHKm4noYaSTqd7PiYSg
YW6rn0SYv+yH/PvWWAyDcl0sEB3I+VyMt5XzLrowHzqouCdv680HpiT2x8mkLfWB
GEXiLXUu+rQksw6n+A9sI679WuD1kUJnXMTv+BqB/q3nvxsbhaxDTpaE3Pv0dBE1
et/9F9xMEauDxf732o1R1lRfQsXKuVwy3lWLom5OHSoYCSdfOs8lAUUpUzPiWcuC
8wynwCya5Q4W+rG7xd0eiRGsVG56Ke/IlMM1+Hb1E80aPyrq3/YApEyAIUca0UlZ
+cDKnUEyNQgucFngy9IwHkHEDLiYs9iAqKAm++4Yn3gV6aLHX6N0GU+hUtn2Uumf
P/X3uPxlVWoNx1Uy53ASePviX3WFc22qTHCBCJPdzZq3KHih2riPZEbOPqRgz4yD
GhK3WFGJ7LQ/sssKZDaUbzfpE72Nv4Xz70g4pFsco+TE06SeBT8lkWYGwgYlw7eL
UwUWc6F0+J1P2nUVwfFWTHNyoo1HMSHU7B3wb0+R/nz0Ygo+pDzhAFjst4tzQdPX
khZ9KO1VEyznk2vf3zjSRwygqR6baADpri3ivGg7jOE8HBoRI1x/AL615cOExzKo
MsHiTbboxCRRYBfd54GlYcj+jGdlyWQXYmMYRBsGOpCNhbraOrMzI+4oacIz0puW
JT9OUhbFAvzGsDhg8Th3HUP5xm11VIFMqxc7vqIhaDeGZlpUFuy8REyOXfIJNT/x
JPUnG9rF4UE+LvkmEp+d9cKYn5EJDv7vcM2lrzI685H9LpMjutPMI7mUQKYhj4Py
Xg+W6dwoAsH1abF7PZz5XVF/OOTbL+67w/6u1CzvA5tzcZ1wm7Wyjw9goQUTqyDE
E3HScp0NeWfkYxCbaAlYeITAJf9c/nb4r+6xRxCVU7oSpPWPWcwgJXsRamfVMMHG
6YMRXOpEzpRe7i8BTmzJsDvrwi9nm5ytbHzA97N4wUkOzs6Z2YA6j88s6Lm2F0D4
t+1dWC+pzj7frqEYDrvoCdQvTLpjZLtIZQn0F+hV90XL+ixyDD+461NetWWLF6th
752OMqmksYBPZ4KJ/uvzqukOrOL9vagV//macGNqem0SPum1HvRS4KWnV+E17GhU
H2PCDBaFFxbpBa1h5NNJQnNE5UpCEa/58JrM2qhlagKhr0eRyjl9RTI1UN1eTXwO
ef4X1d0FF3/9Gh2SNWD+CrBuEtuYDLyJJGe8yAaB/g+qcgB+E3fZ0JvEjr+d6Jx0
Wkr5yq4b8OE0G8yPKjbA5zDMpTxtAEn3gqMrlDmPsxkeO7/RbzrRYcTYibL4EXZk
iia6F1qg359f1ySxA6VXknpjHk6c/p+eY6MqkUtK3iLtuWduUr5mRmfjOLwxxmIO
eSWuz6UIi9Gu+mnK6rE+VemfTx4iMMceGbPWQkpoYVBz7oreVxpOCDL7ehgDYFRT
PzSie6Yzcs1RNYf6td2p2EoiHUKx5lipa8/ZQ1237oQn9ukddiyEbdbASSs0e2+O
2gOdzkjW8H6XOo9xeACaBeBw7YcQ9fNecS5fSarPXWBkYQDXuovWJKZLvdNEEggm
aZiHxuyP8wLFomOmgAw01ynIYEOKBSTByNbexDAAqSoDI5yrO+k7lzQhF48oZi9u
2GX2/MZX/3D/Z9PRBSexcjuTvmp6/2B83ZfPhp6U/QLLGsH65cMNA9yHCG1KSqAn
tbIPtyaJMdNBjBQG2sffQiDvSTEzvVYPiRXgrLPiOkVItDu4HlsYs3AITD0vjMZ1
vJ/3JxUQvxFixE0z273gd9jYInxdxPaEukqstS5qpM0kgYj0TYE4nKQNXyWRw0cQ
9/25w8jqGAh5Jj+8Cc0/Fxq+iTphqDynjYvYB4gZIZSRbrVHfM5AP9+zOxgiSNVt
fLBecC5xtl2QMdCsLSCmv/jmg8sfryi7jygK6s8NVLTa9M9uAPZr3TQI7Pr3rjJL
HAPZtS76TqY7auuZyhfLPqGHR3FS/q5bGGPCfPWqJX8jLQ89f9IRRV8tsdKn/LeM
Vt7bJiascBzYgDzUEMWAytvKyy52KobUArz4xdUQDGTNTwlxfkOlhtDVPbq3DmA7
ZwYZqQONHjwNrI1S5uTN903M1/u52b2utLuvzGxcuujDSJL/6Sny5n+SFPaH+Bhl
Qxmcudx6Sbb+uxae6hhk9ZelShJGsaL5g51z1ZvKFodhWSgUFaDITKXXkNvxd9/u
W4R2M9/sBZRpG94ogz8kP+w6NYGptnFCvJrXLYnwMmn+JcmcBeLpFAewZwM97sGt
rKYtGL/AVB8AEQ8jC1F7gepZwMzbYEcX0KTUIlgFkZIIN8dVXr0dReK/bGCsVKDu
PPxepBM9JnXttDtvVx4ap0M0IeV0/Axd/FqGE3lqkqexo16HzkTGLDBmF8TIco6V
DN1DJQmgkZHuafWyt9Ic1q8A6l+ZjmGZRGDQ6Ngizc/YQ1N7j7pkhqP35PCMTyHY
MGllfRmGM7ZS2sWFObkRooKp71cMKy23aMhalK+T6hTc2WVXrK6t42OE+QCGy/Dc
1JWzoEJ+eARMxd9FsLZIgN2EVWo4PxIgMTmfV5PNnkk9XxGtWT8l/h4+/uaGoLMR
753WFhk1DhdXIhCbJNeaVXDyrHwD31BwcjygDwTDWSRx6IvRwxqLFjqQnOKLCfmH
hKWPpq0bK/Idt71VSn+KrtU9ZqzD/Qw+9lGekaRPQkqqOP9Dwzz63rRqJG9ytw+Q
pbFpGkluaCUv3o9o6LsnPE6AFF6LM2jinHFKK1cgK5YIBUo7ncZG4qFsb3ikX+Ws
H8abgIGIhYuhxkeYlM+PrQiIDn1KSdGXLKXPydVecM6m2iiePbyuNH0ktZ0aUpj/
2Mm+XNY3fIw7/dB3btU1uUR9JKX2pfRVP5RMrpxRUK+8TlsriV41SSS6t/4BMTd0
SmwqzV+v57NPcCVJApiaEYdg4h10UZnK8qNk0gqFsnOwQHvsLdLu5QEGQYaKDh2u
lZEAijs3GRFsDglP0nD8aivjqtTuynIg3+KRF7fsr29cmr1vbDYNZb26PLlxxjBt
NrxTcjfPMpmtOFDC39pO4zgarGyX05LNyDDNduUtujV2/LZJVF33IqjPzbF0rhUR
4pb5GsFl+RYmcEOHOo9A+YJHVCoLXsR+p1E7mjQEddSxwKBGgaANIhzkPdPk4aE3
8kdXMg0eXMDNiy7EFZwVACRKZx/xNw6C0vEplUwgz/nXdf29aXUAL4JKrS/cDYXU
KlgqMAnYzFVnl6yCVa30ROb2qn1jX+wiBQ7z5COfsoToMKPU/b49mW7ByrIvPP8f
GpPylaTOCG3X14j/BQddX6SAbVJiWa22gVZApRAxrr6Y0+RCB0GTZFdnFq8acUER
PcuxErTlUESI7JI4v4fdZ3N4AKYtCjmIBessop7rgNE9XnKLuMrx1yJZb0Q+jqy4
uy0pes3NB16lsVHqjYq6Qms0Igg63mZOM1tOcxcrkTlq8BmH68AcSt79HpPFbIqy
AkoQb3O8t4M7IjorKH8WHoySQzZ3IrOXSxSQHvUN8ZDIVN+Cr/IWrVUoG5RLyEPs
1hjcldVoY2Xw4xcWGA3yuEQoz+5r6StHTuyUp/wGVHqLP2oGAS0NzrLw9pGTHDNY
t2YGAMovzT4hV9fC57jSiW4YjKM2byfltV+RsV3bOQqNZ5jvhaG9Nsmpeqg47R9I
RMhDVSkkcWX1uD4KvERJpOqfGlF55QNpljS5d5u/9hQLD7IZRK+x0StPyciHtVDv
/S+jP8V81kvJHXgdtqELkGoJzZXQO3vSAdQR4jsFONwgrAE2TSwibm7Gx1w2I8pC
wjgV913bNnlFOPamRxOWpOrQCym9PbTPxYO/OQ+a9LulUntfudyRkjpHE1Bng2yX
6ghJ9Lz0OIvcwDzqQKOBDzm0+G/Nlc9EKxBONU7hYD9R7OT45BBH/rekaGW4B7xN
6xVMpBv9GO9ZsMFpCFnlhqgdvLzdfg2lTfbh3Z6tGFbeDTsa9IyD4biihhl00WXa
1gwkLywRLiPw248B3LQX0xFLW7FJD/gzd9Cj18LdGeWMwa+11c3Y0ZYdgcr1uMgB
7gnWLsdNNE2hPxQrtyMlibNpwZW7dZPlL/mEkfC+heqho3r/WNAzp2qkScFzvlk0
GMtv2g0ZOC14662TkP977hcBWtnU6h6xSeEYoJTZRIA6V86HHgwFBYy0abYwUEpI
+tuIrg2sBt+/RXB8axmJezQnwDi/VePbPe+09s312kNr6KHuShpo0yN7xrZkcDiK
uodpE4dXIVUScCZFMRtjuynpSwDB+LEP6vD1UBwslKN5eEI6ydVYdMkiowC6Ecth
AgcPd3tm5A+os3+E5/HSBpr7WWAcsm/dKWUMMVL6fvQiZFlsSyC0l8ZyjXaEC2lv
OtUE09ptOzo/4oR49MhWikI71P5JM3GJzo+YKYM5Pfrox5mmq6N7ZBtrFssbicV6
NnKmWx2EXyK6DJrM8JM7wyEirCY0mmkMCIpje3vFRcU7FcioFaR3ic+pyG9OWDsM
QXfC3JhIIWCHuM0eS58jLBNQYB50XMk5RbcP6IYnTBi+hKY/JMLm10J5jPyb/tOT
sTDARzV98iN9rZb0oBOQViQmF+HoPD3AjG5a2K8MJBf3NAwbQF3WCHbXmo0Ji7Yh
NAw+YmV78Uz7aQ59bhp3TcGvvuv7Kkf1J1C/v9Ewc6Bm+8BWhLjdRnRoD/g6ejAL
cidLHbnXipd446Ch7rbnoZ67FDdMrI8ZJemuNJQOTL1lB/iYWlNuKR3Hptm06rcf
kX2ycCLqfxucDhOt9TQavE+8lOHLv1JSSAEqnAsyU4/jieVT9fmiHXS/sIyywBbV
H+uR8y/S6kUm3EPEvaosKvts4y8jqvuowTgrMU57yCPXOA89wMGRnY4LQQOX7bjR
aH7LYcYT6SvjJmu5yjGcoxIMQkwb4CJnH4YwSmvFv4HtqYGYsekGT7zTCNljVHPD
ivM2PScdHf9dr3Ih2NNiJi0b2MS/DqG1A5o3LFajYSfAm3vL8dhdqpnUzzvM/hpL
cUy970U4VfrkYOJVjXLa/2G92c5EOGot4BacyCKPNizTKA3PotBv6TUEAvuvvC7d
Z12mqmzT7h0o+KUik2ssIs+uAFmYYZKm5ouekdAaPVax/l97Zl6njluQkjvZJnYQ
kD0uUP2ZZvvdxHoMQnYPq4qNJduw3h/vK5CfV4fmn+QOBAMBlAdVnklMyYwhDAdg
lNZcZ21PGzQqHJziWxHmDtUdxyo9PfNdasFAfHME7HzO8HFICI35c4nJaDmsEzHX
UKcCQDzDw7Q8E2RhgY7c85WEqo81UkWPv0l3DyhbSozDleRZhHg31bHc0UGXKsYQ
2dKxSJ7CqeWjVOH7AVme6v+mK0LBkyJrroAqmM3h72k0PU6tSvdL5uhtRTkTVVCX
U8FAJC0ooOHsuUGv8fQsVtjBebevMgrResJzrGNwIXcr4rp2JQnjtIGINzhpJMBo
ApKaokEqmRGQpA0Ho8Tqckr4zvvanwEob9xUlnwfU13UzE0t+P87EZeBYU98qPfy
XS68jBKtNKoPpqQzH6R3Ffdf6isQWpJ57soU36iV8p8J/Y+ujl1Ui3vZfYV7VKIq
Af8NMVm1qJbVUuyUOi7vNq52dMUrfxGrRJ1giXAlr3m7koMbPVUq4kJ23THlIfS6
YNc0eYU9Z67IZUcHecs0Ct8Si+ZaT8MQStg2dY+10Rh6oz6jq/rUgDQfg2UMHbmw
Pl9wh9hyUj3mn5Vn64nL449X5fPSZP2e3mtGcAVaqtl4ff5UfxPasxGgotsLJlWZ
cOaSvM/7poK+2aWOPt0BmWrKbUCRnsMNLt/ARSjV2MA7/MGP3g8sAJe4aNCmQQZb
Qv5awkFYLa6QHJXy32iQPwBNjOhyA5uqtwso98FInSMSLiOdakbu2ibhsLTUflCu
DAb9PL/rAlXJCQNjaXsEYgORL0R8XSHryPoYudKr8Bo8jksE6neetkjMSrYoM40w
VdYXjrze73G2Rs+AbLpN41k5Uurt1mRC/kXeobftFV04nB1lQgACV67TfROBSNb3
pBSK2azgjex33eNUc+LdnkEkplBh5QT5j3QSgxu80GVsxS/0PP/usqH6BdhKvP6F
iHgxijwIYBA46pdoNk9O2E3qTUK25PR+MancIz9svH6LSvx+EZb0nTgtooqNI3D3
QutCFanb/XSfD+FfZ62y3CKRQ6xz+vuAJ8hPj1QKdqjLh79+AP+JXLgTXVRT7GV/
GMexnMuX1xRdxCc8AD1wTxaT8HHM1ZS7RQ6HasxosYq/5CvTY/ELEgKKRxFcINlf
UzyR4RtRBREXiI6RwkEotOVQYVCgDJbfncfBaH10p+CTfd/AtOxFpu5qo0Yi9v0A
OL73uohAO/MTWol7qRLp9P2V9iD4ReriefMxemct0BsK6C+60c94jPJMHR0z7ZDu
b/eAxmCcUk2WwVyeZEH+mTiTZAMK8RnaSD3y/K4Dcs6AMzFR+2mjHkStSOW3VFm8
vWs7Np3wVj0s1yH7tVW/oMBb6IoUkDllaidljHA/wHaodzPGO2lOiFWPTvCydvmn
qpyviLMquTv2XmMJCToVl/099+B/2fV5K1RpA7XMwLayZGMntJjjerRVmgR3QC02
oPBylkSqmkIAjKLDxSuVn9H7hu6Yqx9uPnPFMoRm8nqj92c2ZKJ3aHTukfd2EMK8
b+Jd2EJdayjX7e2yxxWec2ifhStnbKLI1LUZ7qiAp04fVtImpB9dujGZ3nd2zeQr
Ge1Tp0FgUVOhL0sPLgkOiC5A5DLKH5sX+DwQIyn+NZRWXqKbnT4IFGaIxXqsoTHb
9KiJWHsjq24XOyaqDEoYGlUevVmYfHlRTE3UiWaa6sgZJFk0H9SU+34GO+lI3RZd
Q6lOsAnXYnyihbwLMHtyMi+0BwNDP4USPsdP130MvU5/+QTwUC+XWmu9gUMgxFDw
ASHgT8lAQFnmegEifkEtic1hrx0ukz7KUX61WI/lscgP+rxCK2DxetMVZ27t75YB
OzgBAxrMIPrT45NX/DRKNfoCbl67kNiGd+Krg0ZqM7DqoD60k1sBF4wUedaW8Cio
w4NOh4hA/IB+GN0AJauje31grbT484n/HSKtGVjTnDFxyQpo86IcL6OwaZGHRhZg
ItrEEt4anQ3Xr0mKI2Xn9t8xKgI2AMMJVfEqB9eF5kRnpAJOaV6GUeCUxuqb28WL
mcsfLEMvKLgVKrkNGQxUj2gLCnAsHKaJ/6uQrunTvMVyqbwFMsiRZ2ZyKBj0Os/L
a8OSOQS+CyN2FeDhUg4oDNq3yyIqmhDNknzUBMQfH6rubNvCxPoqjV9HcNctqUzK
hcuwUIZq2YJM5Uc0x27IYguys8WyXSS9zX+mPgSVH4j9X5p8+NM82JXPALapDBoJ
HFi3vObcYEmf0pO5V6Gm48isWTEXs+wSMi5ncp6bwNovKvd6P0UYe+KCLIamClsk
pQplmxVvMVDmrKvZVgWFN7/AdikJSKc1ox6oZYIhcHJvfl8oJ/NdbyFFLOAM/URW
1ypRuw0QZ17g3SO59zixPZjVt1gttVkkerqzzFXuDBUaA60jd2nGreHb2N4fa4fE
hLDY5IXPAxVDzfAErl0ebUG+eamwMObtRXPWho/ZdCXBAWp8Y4LWrT/swYjL0Hz+
crDBMPHKv0oqVPpcHf2QSikfgKklhd2BkZPLAC9uE4iBKcls7jamtEgCN675hU4X
eJfiHQTTL6nMZnCJctVsK1w079M/kkk91XVdygbeeCmgCIX2QSKqDq5SBGQaCPAy
f6LTL2ngCG9wa3+jBj/xviy1snOPGAqKgqUyDSmJ/+kNEvUzGUyGnyQ0qr5CdlMP
hrMrKgEMlHNFbXnMG6MXPCv86eYUlZFHhQdo6/k/PsVQ2+JnI9xwCFUUMzjAFf4B
RiNMTMUULFjuFGJ+KFdO0GeCXFAXI4Aw93W8zEYeowd0ymkzY7XISXowO8L0KlfM
xd/XRlWX1dotltd0MEzbXS5NGGFIfSzI1DXo5UlV0b/gh2B7wUS5KiL1T3mZZnNh
KygZAmFKAbH88xZUSwmvDwkz3njX9YMcjkAyRsOJxMIKUN0TO/mL/1YAngDq2PnM
aizYro3jXGbSm+tPnZAnTGHCykxuLlrMgJy+Qx8045UDn/uKdR8jtx9qxOh7OVTh
oEKyZF9UTqyL8wY/dsEjFg79r2fy31INlHzsGgv5AapvhOVqQCyW/5u5c66tngqV
9LxPwHreYJdsjAsZvJUH2EfPSQH4tq8WijIVwdShb313sUpX96uSr/Cs5Lka9joF
4VFU8KTWCnSmXOpDXRxiNklbza62h4IhI84DnqUQxWcNxQ4n0G0JeoorMc1kxOBi
F2YikZM7oPoHy7TMqWfA3rB8LHR8YDmgcTXos8AS9mvw3OfaqgJsW0JBJhj3Esm/
htqSyKIwg+11qGjpu9USCze0MkJntjcoOcjNY/V8LMy1p0mpivEQeOjRoiZ8CrE/
v34ij4McXocBneleYlzCk7FH14MlbdDJAxvk/gZKw+5tJqSw/HUTqEeTG06fy/J9
ELpuCtVs9PunG734bewQXMSS+9ojBEx0A7AA9qrcILCZMaRyXKxiio/rWGrlpMWs
R7wnuAgb/kpkmJttD7FhB48adykc0P5MbVaTcRmfhN/iOSoi7ynagOAfygaBK0hX
QddRaGkBfd33o66H4mQZhbMCBaZpSXG0sH9QEhcvh72iQcNEnuFBn5FCKWXWfELq
IRbzMXjkhR78pDsctcdzV7eHtWO25KWdi4wvsyk3qgrHODC2fsD/3Bjfe/vNm1E3
HMsGNb4Pkgg5E4Vovvm8otLQLfwqNx4wX0b1NKBHV9gCDNaB5/GMQBQoqwhytN/f
bpSYAQU6K4Q2YjRv6XnU6W58opwKxcwprMv8h8pBZxjdhhIU1IUXlzOzfH9/CtL8
kunwcvkhdTFokmdt6o0bsGFGGZwe85uiy7UP6iYQ5owFePIFi+PWiTgoMeufwNgz
hBVD9UU3slaYh+WTlQBGgmxCAn7RCgJxgnbdLyu4VHOL9F64YmfKRpHqzpnx2LyV
shNJxFEDZyZUDaIzyYZs91rVmno8lYtSMSl2J7CMuvbuqI7CVX8G7mT9QWjTzWkm
WkgM3eI7Ub0FgZGcB78FBWKT5ukHc7icXc8p71Qjv84cORz3IaTKZYNZCZtkligd
8uUbOUETjYXRbm6Ku84+Hfs3TnxuAwqPGSJkp6SILn2hqEDLrfEOt1Ya0EteGhUt
lkPGYorvAssjwtB3gERljXCGS3BTUtDdi+DWQh6Vt9fpIqXfGkRUpVln+w3+bm3O
hJMrOlpA54WPUgSOiokClRVsho2RfQKWtb0NvOQXAgyiAjMZBsUvEPHPdr5g4NM8
nyOk35boVGBsQWhLhHWMmX8rxXfudfjkSaqUIr04q0mls7YxrBBaMEXv1ljDqqpQ
E+oHwBYKM5Qd34w23zxu7egUCcygeB060iuC72WsPCDqFtZ9Jnq0Rs5t47FV/ngo
6Rnk8b1I/7ADiKZRezhAjxHZ8WwG5anTFPZhQeyzH+g3jCrMNOG3AgAcfcpwlmZV
pwDWQ3kD0+XnpM/cL4UqeHynzRqpHqSeEoUegGAbIVQlsr2wTtdsX36E4z28RiHi
G3+h2I7gVQ3uiXDIGPux6FiTnmSkGhZukvAA2YVpVbab1l10F/4WXAQTj+G+d92r
gt0RT27SZe/1RPonad9ufNgHW+r0P2jo0CtVdB7oj6Ce554Lg5moIleglCma+JJ7
y74Ei200X705yosdQdRtk7YqtFIdIIK0FipZsm9s2GkdJLVU7VJ409LdCDp6f/rl
/xt2crkerlskn2fABKe4EhdukSH3UDU8pBdxo6yMOA2Soku19/9OZ+dusxm2joSW
OuFIjMSL9aqHE5wWTzYK7atEIC3NEVrejlUlCUoHFCdYKgnXQfhCrBKbQ6MZpydT
kwF4KhlIv7hLQ8b8pGmBSijPxjvdSpbDeH9Wjf7nQFazb8ES6DIDRXJa1ao4I/Y1
14y9NVMjImzVosX7ga2ifi8ifjzO4sWSGP65ukP0M7H0rsZFOhZtwqqsxlxChLW6
UUlaBakWO88Hk8BTGkCCTlzGo7gFJDMezKFbj0y+SXyzaHTzY+kU5UZGj7A/EGzb
rNBENbFKcMY3EvJCG1dSHOOZ7WeYAeHoX6JOcoAqypHdFuCD+KKczMvIuiTfVAN8
/q65a1jnD674EM/oN1KQhscI4k39yiV2zbPlVtJs9CVreNeYPbg+Hqsjk/GciYe1
9NnX/KeBl1BnCsuBn027jLyU/V0sELw4cTsWEVLapPkYzaqcJFe3T4xL+//ZewqP
w7LWbuX0+Y33Joo7KqWI3y2iy+Pf4GPcGEDI+EtNBqXH0D8DSskyOuK9kvSuArjy
DjVS0eIQQ9gPHMSFkLIaamWvGCODUmxdYdgOhSvpU7+QHoJBs2n4sOesNK+l+jQj
nc0mAe+SmuJaWmgtVYbmfvW69f6WriTWGKptFZ+YgOLjqg10nPsigBbwrNVElG5D
GINYdYWOQXwNt0k4TD/uuJB1GqOfE8+MDGH1D+Dp0G9L1yX3WMPCcBsyzhiHMMkt
aAMoahLL7TCNdKKz6RHZEMbZeMN+T0PQvibddkbDBRExFsewGv8QRJc4Tolexn4b
jKkBXc6qErLXsXn+lOYO8u5mZa2yukuVIrQeGKXTuk3pU3+avzUSECLK0rUIiVkL
GDEoLLvLq5BX7erRzY1P1WvRLifbPgzxvWEMxJ8d+JlaQPCVNimV7cRv2l9QYoXp
U1n9mhdGk3ZlzVZDSkTdy/IoP8VoM1ta06yY3qCcwc3n9jg/OCeCX5Rom23kZCVw
EiTnuK6jw4MSQqCYP7k6vTMHGO2vCwaGcTDyKF3emYqNfZHxnM/4QoUxirMNIgqH
WkKpvXMjRC8aqaXe9oLVbn08SesaY4dUnsyHbwiSjTIUETupLavDizLLBnJhMKda
lmI4yPXRZZOn96qzCLR4AVRhDW3mOfq8rP2v/VQum5yUjMWfL+8HxWaVnx2nS9gk
VcBtbi0ktIo3Trp5/Czec7vFVJEuv44sG2Tb9KgrX+bpceT+TRAfPnZyyeLpTJqR
WevHjNOyR3f6yS7tXVeYnb4T+3bxKvNDw4vwWRKErOxSS2iwMJZn51NzlGA1pu4/
stCDZACpn5ZsWRYbnw7QA8NKodfpwEn2OyPlfdDcMI/0tALP/7PUOtkPLqNtcfTw
Kuv5epOcFqwbgbg+qUpn9A0iQ+BBxqCo4L4hLZZbOcK670129r1TWIfQtCO9imp0
8pVAAv21kfpJM/pohDWirxcL4Z00PVpcVlr6v/dJjMcsCV3HdIoOg0D8tWDkQgEi
+k+CoLIrtPfhXEk6/TwIsDcLBtZ7kz41ucpD2+JOlK3Pywi/fJRWg/d0FghzQ2Ii
Tvfjmo8SDrwEVfo7Ns+d4q5ECyH4o+nOZUDwoeCISxaXacMahzYo3gTlawKDE/td
SH9x5FCqxJuEP+PN826ig0awCWJh40iMG5UQNLZ1yDvOcuqqeubIGr9ZRxWQya+g
Pw0hExlQZ461wdlxZ3bH/JNm51Ij5JJUdRkDt6XUIRC6p8o7mYr1glOR5j54Da2l
6xzMpT26CuWgdt1p05mTdcsrUg5Kge9nGA0zD7V+T06eCn+xDx2wCphBhkOSJy/8
q980v3/zA3ggClMf7nbqhp2+1PPsC1IkOUfr91X9NZHhkFHrPLGWSTL3Dics1Owg
8ymryb+seQ0TOc/A3RucMk2RH+cEomcYwcRmlRSpiKBMNCJ/d9pr3i+A7GZQZ41g
Krxw5uHralRC8BjK6F0v5SIbKsH3GpUu7Or/8CwL2oBUZ0GDGUgvP7p96TLbK7Bs
sOpzohAPiwI7+E6SQ11ykUOR4+5Ro+HDGDLyxq7Kk+Q9+JV9qQCfYzFkWv3TwbvV
50IY0hRn1EnA0jesXHmolS/P9e3kt+QK+wbO+DV6lGWBKcs51aK0qyoO1nX9oC6C
AHwrtyUOZ4IgSzgDVvXuIYceWQSvdlh3/2LT75T+t8yq0S93H3UfLuz/z5lv9eTU
zOZaz7tBI0GTNVJgvklm3upGd/RdznCahz9RRy1/UjdjAiCyUkX7SftATGLVbfGI
vBVC/CwcaVFm1NZkJVQIUOkGEST6W6+JFFRcCKDg5YMGJXmaW2Wj+q6L4BGNBMgm
HImODf3IPAzYZjC/DbEVkCqsSYB6e5lEgqnoLa2CMTvJUZ5GLIiJEG6iB6J56g8o
3vnHPy41fIzbIIqJ/ZTwyFHRChBv1Y0cRu+aOZ6zv3hxUB7s3ifIrdhhHD6hZ+rG
IvtBTYBASK9Y0X6mEPy3uujoIRihvwjIKFWY25vXHiO4g0SZXIhszzqbFTu1l83K
macXJLEkuTalyq6epCHSD/wGyb17iaQGo8DFO2pyfk0ZZk4iOtMY83yzYZter4g3
iDSdI16/gOLySbyb++5EdU2WJVjr7qbEmsAO03UedFhZPgvOO3nGMBDfgcevGTFA
l2tqUy4SzZsM2vLBqy38Mbp1qf4JkDx2Tv9CrIFhVLIrtC6IsLogqsnf0HlQ5O7E
aGNhNc7QZz3/gM/ZXyPe/cxwl1l5Dt5HObfe1DUPTQctBXTwRBFnGOwxA0DUN0cP
MAQXWCjdgSsRMu8wNWWPde6NSVPRXfArWooAeUdK2pe60H8xmxBnNymeKW6JBOQ3
PO2P2W2Mtz20wQv3HV1f++mmhAP+YQ3VfxhHrg+8NmZhE9WCImeVJirYvIk5y2JO
20tXypS/qrEaTQCEaGEihEE8F/3LRAdK7eMmN1+/uF72KU0p1zcV0IUJiNthHZm/
TDKgwUEIccata5mtqS3EWAopVpupI+2Y0YQA/NCzhswcIxaLamAeVAV2FSKFjwyx
THxJoqtna+QZJTMFfa4+e3rfDsodzSdpXNSQuAYCDuqe9H0ag+nhQ+7WmytoA4Ja
tUROphRnPk3yyX6ojgJ8qTW+RL5pxIK6R7qX5jlcaO3X3LyASiAd2jiJEHZyQiT/
NCP69BnTkQGrjvc5q/ksU3iqwGLDm2Pz6Vt8fBfTbsvXqv7vi3AJajVmZ2k4jBMp
moUJuHiKQ64wzYEMKpOxFCncPKKnVW3XC1/5h/kDHokYQHNEqdzrCEt10Pglj20h
BKbyTx9Mj7qcdtIqzoFElSDixXINozmKtuV2Pht/anjRuXN9LcCDCjt5JyofuOKH
yU8284afuFbUs3sGxLag+bmdC5e505CwxAmhF3r9IyctxwUOQYUDa5XsEuBLtRxD
azqpnz2I+dBqkcpq0UPoEJExxxbkuIsg/l3XhkLbtlWpD8qt9K+h6tWQp5hoTXPd
9/9v22LqT2+nlk8pFwa+n1MSDUmog1GzJmRz+WlwxfDnVjn/ftCX+Htvua4obVPv
I++CStN4kKiXLuCdRY0oof8NkrTQqK8+8z0VFd2Fi4tiyDJZJR9BHxXYVPaxA+DH
kRFhZaBkaAhWFLmNl0CpZOFgse5JZ7h8J3wOCXMQJleYs+MafnSCThicEfEqRxEN
JzHB32yMaLKd/l2VMPXiYGcT5pmK/LRawKHaJ57FhzO/9AiayuWHaS4QtrM12sTK
x7/LQ1PgJR4PQEfGWlZi/zb9PtVx7sWiYx20/6dn3JqXm9XYow4jy1aYlkXrLQdo
4YDkLbR74TokYAztlIqPGqWMkY3kemnmwT/YwLv+80q+5sAymQkr7CXDHDm+FSwv
2bKa6zfIO4donrXuS/tQc1fMnVG5o8h1C+4dDvW+IIiby/C0cEdrd3X29pbIuK4v
hnvih9E3z60hgAV7KjelKJtehjS4XXR6BeQhwrqGvD32SWS+ueCyeFmOyBVquY8r
2eFl9a3edoAg9uTWkRdmCbXmXHUBLgAZNvsMvSHsCmxWkkoKpUPBym11KfQIriJb
JvPHuvnwyvglQE/5DTa+aiMPbak0dILYlV0+Y7t/AhQQ+8Y/pb06thF2GvEeB+Jt
p7BStBLmpUiLlfuxxteF02B8y/zhSX85VkX/FQE5w3/0MttPHDEiLnfS7MeZQYbT
wixE4cfV2CtuDIqy0vh0YzHtEl9IkcX4heYQ65uFjxmRxGe6SuU1xoGUEGqO4kSY
t2IGfCjyMnAE9nrrn7YLittF+IdKlecnYcDBTDanSqKX27894KAjHaq19ID0avf3
gx5TaRYTb47MS1LR23wFncd3OCv7762kBOvUNeEe2GeRKIgD3hH+FDNtXDXNiZCg
l6oBQXHvMXqlHrgrBcrzecPhCPzFoJexPFIUX58IN/ldmILBXYWxqT74sMpbcZdW
pjnad061ZEKnJp3L79CAiMqSNHkHt9Jtef7vRX3JHC+4IjH4BMwLo6aVhTMdhJi9
q/RtSSTdHvMyTbAhbQWyTwDbLdpoKm/9ilnpCsLv760SH+E9HzxDTwofPPnzZQ1l
Zlq1Zz3MB8gSp/nbWSNQ/MjebBN/HpFJsTKQMqLuwmvVf5PSkON1wtAwMKiSp5mn
9isNYJLakOnawfeHqxPiiyG4+Pe2z/4RSs56xW77WAu4OKeA/X+Owi25/7SDhAqh
I2aip12l4ZnUp53fg/qnTgoK8fa/pWko36DkPaQA8lKEPxdvAMTpYoOJ3ZXvHklZ
nKPDpBgNidzmkkVF1DR3+jncumuUT78A642KUsNc1/odspqDC8MQeX1BUUIoJHRm
nEhEGeAzcXZ2eikX0ynCPc7Ib70xZkJ/nqOkhOkDmUupCvZ9cTWJDZWATlJ3esM1
7VONhQNL+mA1BjfvZqSihUr2YIrxzjIxRC31hSMP5YpTjQDfBfmjgbDO381n6VI8
r5JUl6ckljB17ZQsrtqYMB34sBjR+eO8j7qsCbxqe17fHtISJhfGJneSgRSYvEXC
XXJx8QljR/VVL4ODV+dgPxeqUPpRPwgstoLbeTCXO0GrVWJVwCD9BDcdjLtYjUfy
UDickdwWN5ysFATYNRxg2YAyb+2ZD+w6F2Zt7KDpNvTdVol93dipbGaaY7nlLJPm
mvVOXqwh9ephvFSNRHLx55q+XlAgK1FCCc9wX5+B+DtiW4RjXUcPnvj+/yTxtSyc
Hmy3Rc1qk9ch1TmGnJVPMTe60zQU/KpcrDv35cnN8gGUH5fF0zsTPDQ2jq9/SkHH
NV38iZ0pm8rPevPIw5nKFs5u069HvNj9B149Tbqam6o=
`pragma protect end_protected
