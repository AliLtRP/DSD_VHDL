// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HWS+PAs6Wr+wq+PbO+yckY/po8RcWyMWyucelw+tgPcURLmLEPDYp7C4F+3fmXeN
JUYka59shwYzoCWP9W1DjlLFvWoLjFM0m4ELaIBT3VsCxHe45Qa6QxEMVVo5Z0X8
MeMbsLqw+XjxJSC2CUtiZLt+iEtwvGtnD7I5vHeoEHc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11616)
OZx7Wa36XYVoFNBLfe6dvsEEyljmbVWBs+nRpfTqemR9wB4RYmvalaS4gFl0DTrJ
rG6j3maeTT4PXAIS3ffLZG3sIw/oEXnCCoblffRa+IW3cf5eSmKRW4B/eL2dMjmp
JzHfDK2profUEEPaFnpQiP7AIMFIB3ymrS7Zi8NWGxET1Fvv7hfMW04q4KgD8lPj
IcmePqjMRaL3Bm5t+DwaQ0h9Y1VuUibYOB6KEHfot84v2qSPM9a+wQuJD4PGhd3C
i+xQ6YBuHKIdSnq6Q8ndr8e5mNIre3pa3eoVXovQRBUfqjbQqr4kJyn2kVsEkVbh
EEIUdZGaPEU1z1GUGoOYeBQS59bUDuV1CG5XM/1G437KylYJov+HjC1HcSwU6b2M
fOXLqy1gcmbcI+vDJK3GMKM1mSVNROwMK9uHzW7IkMJ4Oax+mfnm0gr4Q9vl7c4s
fZPVzuRKIKXtygE/VEvnQ1v5GkQWGmryMBC9JGMbaJ9cnKtT5aGv9/4sH3oEHkND
GyeLmyP/J29mdhx3lKJgCDdgJWa0FmUDvXRTbHRG4Ih6vyV05+yXI1XCcF+rfv+q
EJ4VCL0bHzpnsOs3qhz0a0xCJ/WhMWj6EymfSEOTdUz+RcSCTXrvSo/0a3g4KRIu
xDqIx4M2VRhUaNVmoiZGgsppZqWfZktiGDoR7/M1uWBPonnnmeB+/Hmh7MFESJSe
cLeh9up7gJmEbfg38yf4IT0UnH5YeopaAxul7sxTi8JYjX/MyLZG8EsT9ryfTLW7
LoM/3Zk8JRAk/qlksGsLBlygRoK5fBJ0QttJCDvoB65JNTPszQo3De8BSUdKZrLF
vX/LkiAN6tg3ZDyGsT+z4YMC3GvcX6b1vB8ZKEJikpWQgGrzDKLVycmMWKkegRYz
FCd1jUS69orrt6JcuKJlT8XuXPsc+4nN5ImchF+LuJeFS5WJZYoOWA3Da1P6wGvE
2UUBTkfJ0aqFSKCawh/N88+4s8VJIiWKbLMBxzNmQmdZfI4fk/1SgiBEDliYiLrH
F1tB+l9a+PCTKkz90xMQOjIMGsgSVCXgqVAJ6eMsfZmkVtcPUOdFtjjhISvqKaZ4
RdpxJ24h4Jnf313zw4MsbkxSnldEd2vd1CE9c0tuFlNGQbsiA5TgnKjduR/C6xZF
9XWi4HcGBzj0lpAyRSf+saWKjemBXXK3+Iwe9OHD7sk3yNc3mwsF5wr/ATELJyMy
Egm8aktYDDKn7CdvGsZd8exwHAI1RAdVlZUj6AqY/JFWyFsm4hoHt8RSj9Bu6HAP
2//oQgzuApV8o5Rp4DxXW7ry07oT2wLxYhSEL2/UGS+NYTXtbS4hbd5mZy24a1bZ
Uj+H03oYU03q2wMF0JZ29AsdTxjmN5UbBDNwZHofHzMFeHo+ypjJRmu2kjIfPlWt
sSM0nhdfL5MCebcmQjyaVtmWtae1oECkKOpyrI8ZvcHJ93tsFUUBSUrwz1nYpV/J
u0PR8E+gdxpi0U95T7ggg+bq1fnGLuPgOa/8Q9pXMsNT9X7rbXQ4e8+yaLd8NYEd
9yl1g8NSmEmBsMN24r2z7d5JWqAVIYb73yDCC+FXHvya3ao/GXjh6gZpdQliKVn2
Gj/Q3WARP41mKAVOpH5kHp8gPMB6hK19oWAx486bSSMu0mdD0Suz6ubI5iXcz0dt
VAAiWuKP3S9l0UyMZUc2B0Uw28Nv2+4TtNiFxtaIpRIbv8ouCkFiW+64i9PrZCUU
37IFifVR0Ft1wf4DcrYE/eDJvHVZE7GgaCQB/o7iOu8sk51ljDLhxORNIBxAueAF
mbxIiNXPjkQAchGVKqfG+MYHuJmG1vt76Bp7ATDHE27B8ua5af8X+B0hi+mC/Urb
Q8sm4SvL8KihxG3p/FT5yYj0dsEHn7I4NgTaVXyXnhMFUYoQZ2/HzeDJJZ66vbu5
uVZ1FcCn3AxRHrXzE6BkS61eUbG3l0dxebZEogcA3t8VgHtAong/kSzYjTQ7SMzH
Lg0xh6P1i+C7qiSoup2RQWwih4QIAKiXChYwkrO3cHesvKG+4eWhIMCBNOd1H25r
AuJXvZt2TZVhPT0tMM2m+zhvw5ZWXeFHysbUT43DiPXCnoxoGlsaYlEG/fxMcj1e
iBPILe9hAmiJk4FgtQB2fMaGaA8A1SqbY4BLUsymX3FhgGsDhZT4/j7v99SFAc6/
rHBbyyCYQ+aR/gON0t1iG8i0QNYIKCbZ/JuCMZ5oeHvWqO4wftymykfHmxPaz6Dq
ITyEgIOVwxW/zCyDm2JCMWs0RsUQPih9L50cvgJ4KUp3lw6IUGtGkTwSKSl634l1
dvDQaWEcl7R+cbpcWal6xSGMyofFULh2oIJnn/Pf5M0lnebNA/ErksRbd1HE985Z
le+SXMRwD9TcJB5QW+A3gTP8xg8BYO0lwGHqZjDlIpeMtNjxrIhIOKqToIK+qaiz
xjnGavLeZTv3rsb5awYn9VMw5yaUQ5jONMbJ/89nxKh63iYRXjeLpgtUArSFzvLW
jeo3ne7ojW1TnEXV/0aeGCD7IhRJz3Di5p2JoygEr2RHDraHULM3QiSQaxXJjwAH
WxDjEIKs2XsIZQK3CJ2N+keqUefZ6ZGbrOzg/i9t15WufTfjszRX/Imv0etEPP5g
sP4Lslih1XlOMXktzA21rJLE4LHE320lKfx2NNFi5bct5Q0HWNU3s9XTyNO0HMtA
FO93Cab94TdMHcwM9e3AnDL+vLGyidMHsboWT857uJhoOH2N1vIWJ0rFMnuqk4Zg
rcTLrW60463NWaClzp70GZhMtTKZqLEu5V7b1YON9B7yhASvJpjs+F9OQdQwF6th
IVswXB8zO/MWNg1tDtLj6YN1VpfE88KMr+0o7eLRF1K6IOEPPb2+BK1btWiqTlia
6hxsnt7saF2tIcWbkMVVxRJIsya6mYEKlPjzwKi3Sz8Zxp/v4wksJejFvnGiwEC4
ISqthq/yKrDBiOnaAjdaiceZ8t8OiIm/1iJAJDsv9Y1In2r0oHZCt24cIt1mMEJU
Ja60oQghOB6qddeqqwShXFGkeuYQFtNkd+CtPlaWQ8T79xdmcLmI+kPgVWiT7qWA
4SfR51FgEdFtr1Z7ZdXi2kTbzhUv/kzXa/NNmRu30yqS2LA2lR/JMhalr5WVWC87
IQIYrf7VdfR8ANwLbSBbLgQ9OZ9Puf9Jos6h5V9mev9PuyJVV7S4ggepcvuBG65K
tcv9OvDFlK4opzigJ+hxGkGyJ2ylMYS5rVf3Yyhs3LKbJ+yWF2ZHuBIDh7WF3Jzu
lIz/QFTRiXkQ16axStZVbK47v/cGjd2v7Y69Lr/1UqUjYogWi9UfdqCha1AMmfVM
5Xnuw7al8KtZ6zARviAw2s6p5Xu4PrQGnIFubGGwrRG8mgo6FN92mJovTH5hkMFv
menyyPv5l+HK93B0T27N5oBNXyDT6tmlUVKzdq6JKgm77dY5flK/0szoTMnzBncZ
6Kjv0a5cTEQvicdR1ye2PA4pNUED/EaR6vPkjsR6pG9ydj8gTG+ESw6vJzTWYaLm
SqtSs8pT6weuSSxuWEXTD37mK9zFicICJYLzHCj90VH1DUd3Hvu6jzL6B6l/6Eou
V9yIQTy5zJEY5GwZoNHkYlsgXn12ngjpvy6uhF+DJuyXVjBrp6CRboQo3hVpo16W
HpozkNg4dHEpnAiUifGVmBU8LAxIj+5UvYB/O2dAIO2bs7S+AuQwL+SrTJJQ0e3L
MnfFoKpF8POqcsLl9a+MI/8jL+60Vuh7bKZUXVgng7ypP5yIQwhUTzZXs5xgriy4
qZyODzfqLfjMA4FHaJ77462xb8eJRSCYESsA263MDgGseVFoq+2zBrZlsJDc4kP6
V5Hl1rS2Vh0aJ4f95Cl+kp4W+kkB3vwTzGK/PKSV43MYalSayZHH3ElctSiQPra1
68+US1br1aNRRnfw0NmPf+HFz+Q36hoE+YUKIPjPpd3myBIiAs+CAk5HxCicdSNF
FIwwDRTm+jLTHfN1ujVudP9F0pjWf37NRwHimN81Mn99R2FAy+fEvFXqWru7Eogw
yBnU+MPWKVMwkP5FeZIcSibn7qWGJEpk3euGjNP8avN9PBoZD/WlBM9L38GqDacv
vuwzKaDRhwKrP8ZcUTg/ssVsx2rTaxGcbEwLXXr4z5WJ6k5RUlxQbqK7TniktczR
BxsEA0c1AwTZKTQ77Mx9YV89anmAEecruJ0yGfohlZEyPwqnoK8tomGidGxRxW9l
SyMKnsXucGeHg+/FNECaP65vE4PbHx1ufRRGvGZShA4KGSaXu8tqbL+BiOiB+0O/
jrKyJVAn2TuAr+2nnM+i/eBtbQI/ghFzNm7Td21Pk8aDg6MUkIBQpJDOyryEiDP2
iGmwsQ4H38tgPLKIS2u7V+cvr5MKx+BsM9zgQ6bg11xHj++SDT5guqKXmMHUqzTp
hyYA6PfIWX/nBXoJjjwLKwIGfo8hc/1wPoODE5LHowmm1VwhkIGug3cAMqbmbECO
sDEwMN6XnRjh5NN5DtZ3lrxo+wNGJ3r4O+R4GKmwyW44cewoBginU8WqK7L8+Ovo
2zrbbjkw7R3Jzsasaot9G1ecTgOB4GBJwg3Y5D3b3LvYOprJYxRwCU23wrdlowtN
4rfVWwF9aF892O8nsuz9d6NJW9a/4iIqlA1cFu3STCe0H2kbDptoP05s+oAxS2Hy
EdUhydpqBO0k00zW0x3H9sg1TRGwqYhvtC716c26Bmo1i8Wxfeezj23TXvoSAyN8
gjlUymD9fseOdRUDCRM7dH6VJcXUUH8uTrHaiFHgRxR2Q1ChMmcOnSzW9BVynedn
gVicfeToikPwrH6VgeQBKGPbf1wCkG6G7UwaQNFnhxVvzsUaHhSZR34hKQt+h7U7
xZpVpp7MO042fp9tZTKplYfz8DCjfjbXVmEYwch9gcyEEpQqEQZzOdjZuMshodYA
bBO388jjkog6OQVL1bUSXfMB6bwxB7bJQonRBjblHV+hIJCN3SHWwbblTh0pKSYc
8yG7WbB+Uc/iS2L10zK2TOyrLe1/EeJQ5raHngcHEC6DcMyxBupBMClPqWeBdqQB
QSglcXO0kTyqfYlmZXnDUn06t4IKhv12RLrNwmkQFqZtkqTL1Deeb2RAcj5uT4VO
EqGh63AYdyDl0sNy+S4r3f4UhhSjPkIeWJtRdfBH8U05gj9FWkBdlr4SHMDhY8NP
lEQ1S9LUOP0zHabsEF3RB8enyGvau8CFAMVGtC31L3iGZliMgihxeq9Zg4HMhtkW
NbbyBM2Qlfx0crkNjUeoiHrvxoHYbFFzjbBeUZbVWd3os/8nB1h3CXKcvc+RtLDu
pXHYmHRCwa1dE8TXzR3zmqkC2DHraXtHVBnbqxH90lmzNYMGfZS66gHhlJhjN4eW
YakLxz99jgly+DvV2qzbY2X0sGzXPE1CxooGv5GKVye2PGvvJD0fQJ26XuRBxaz4
GFMrhad3BXOGeYDgkUEmA0Aaod4I1F48DRPGOeXUc3J8ogWG26rWaTAS/yf7x11b
2PH3RVgFS8xiHDfo5ZmLududDWUaVXxBnlUf3iBNCEn6hKW1VixxZWB0PJfrZHuL
kD9835Ikz+9hwr2SN1kOIOIBzZU7WLwhDwOwyGvqcizXhB0TBOoZE4ZB+XlS0ccx
6hTsoQcnWKEROu/WwCeddj56sWJb+mBY6TOL8Em7GrGMfIwyup16v+PQUZsUS7RZ
IL/azULYEWm9zHxQsVrF1VN24o76awk8h2Dk61bGHkR0mfoWzWziFWBV3/GyDlQS
yg8BVigNf2Nh1LumyIyuZ+nMyPYTZ9nZy8F3YY7HsXqaZd0MaGpNpiYDZS0fNHdn
/vJQ1tCQQG98f8zFcKUWq3mvDEUpDllHCU0/usBgLUUY/3rWRYVNYnIX0xMU7czG
ATrDRnUa1vHgY9OzgU1LsAFj1Adm3y5HB2fvs2uDzoqxmipEpfUe37L9VUC/aFIV
WsmzBHvewSRgXHCExNyh6y61MR/Ybsnuk3iNdEvwq4IvACwj8y6IdK2Lybtn/BXB
dE5RekqvxN8hJZd/MWD9Nk+PbHNLB7+Nk6ScjTvz7UrBVubJLynHr0Gs6Rp2P3St
BxiBiWRyaDJHh47FytacPvXOvlDfNlufFce+sPOZLqFdWsSmWJlQqITpleTTY0PI
eSi3Y0nckf3Cm6UMRYnGuIM1hHuYG+1BrNwj4v7hys7oHMRCR7imRSpTsRsjNvP2
y0p5aiV8yk7wYkZ+MQcDm8xPsQPxKoSHgNfPvQtHJDvNeRorvAniaDEXOy/0B4z1
Vczbw+ymu1S0uDKFwF6CN3CnekHu8SlwLOMPyvNOWNl3GQvx2ppxHGtX9bg3ExXK
Mfs9JF33SzBP2G1enWJ6KZrW4+T8MsMwN3XzqtaqARpMToI7STPVjs5zwzeIk33t
be6vl2/tcq307lGlLlpDFW7LtXeeMDiFB0u/uOLfQJCvGb3653ZbDfC+MivtIrlZ
JrIiaRhnk2ETKXLGbICJdUpEqNIa754jHz0ccMINJY2tOvHL+3ZvBI36TKUomyT5
bAIzgtY+lI9d/A8dCN9157pFRuWhTCDxUsRcOo0ERfCSeE+H7A2qzo5kM+16sWU+
epCXa66mhxHbSFhIcpuA7XHTpOlDiX10EWZhThkQiNbqn6SiVe96F/GPgRDWkk8+
QGWhQRwXsSff2kzzYwAwcSPnGtM3lBLsFdoUVkk75vrQLPLfiImJ8Xna3k/iJzIR
WBYknTcYV+Xs8nuLK6eVJClsaHDVFt9isEI8GM8/z7TNoj51mLuW3qep7e70sscv
shI6DDaULVfSPK1SKfYuols6GusezlN6oiVSKCGL1MtZnLHE74+ih+zlWyt3BYzx
m+0wDN+boAMJXnpjzQZx0X1Ic2qxaXSfehoacOK1EcUZV6LKaz68c9GFcnxD9IyB
r+8lD1i4joT/KDJhgkSFDhF+3On6RPtD2KOH91AZmReHLgDJHaeHEiU7h0MimN5J
LYz8rBbbLGbT48hyQ7TSEIpuycvTE2SJzJqvNCLiWElfdchTPULF/a2DxfRRCdHQ
sYUwBnS/pCtD2n0BFNdfQEssAN/hRZrFxPjlBe/n4yGQDFj8xcz3BSkU25wKQ6NM
/b7bT7wiQ5vCZpt4S5hgUlxTJ9zdg4X340SXMBd+5d0jVum+IYubTtrzY36u9WXX
IJu/BLzzfOBWcK/MijzZulPQ/dr5kKioqKI95z+Bhr1kcu7319l+fj0Mz9/+hkWk
JAy8p6u8d8vNLOKpYi/c4MczfuJzSH5u/O8nrVSAK1xd3syD+rm4DIZvrB2voMZL
2s6aU/1sidqjIDMVwzdPauUNhR5znlBrvQtLQ/AtX2UuwkwUL6stmvSPbMkfrARF
3Pfh6d17RA05QGdhIkXfuF9sTShRZ9FfH88MhTHTTUnHcaibK7qHLsZKDFuRN6zO
mKQm/yK9PqNYw76dD+YFmSq1y7HPwoBWDxFhLXwh65H2QyT21q2U16jNARpotjrx
i9A+5KzULZYslQDRoTgfklCYWId8UrahgZw+kH4tmISnQPrTF7LXtrEKQW41idec
Kze6WeoZJx8Zvph35ro/iqdIdeLNf/Yec84GIszqAp6VJmHHH1KoSbqPDDGdb2wT
2M5sGsw2C1b5I5GwbIACWJ4reSG/5/kjSXJAkBgS7YwQjrUAFJWhK2Nu/vhRVj3Q
Wtm0zC5BvVp61rshgTqk4f2RuauqE8uAPlNUHdGyTgUxEx845uNY2nJxLLVVqszd
m/fO5tF7AyjPyHsQjkpZOro9ZFp0drO51CWevw46bFNhq+iy3/MicS0Qy29+72hR
N1lN3DTI/1VmRzNb0N75EOYg1DFb/Uc0eaMzFEszFCDWrHt84yLGv7UIMvUTXSv9
Xe87MU102iOzBKrrZ8lepSSywo+lyM8nc6FSE2VoUnwX3O7cYAx96D/XFTthbD/l
SrOityeLDYN2YnUZ5N3N/7u/xgRdxJ4f/GVvlRe3slbRvTSFqljuaiNO1c/IjHXg
rwzFKUoj6A1baILUQWDYBrRqL+Q/EbtU+hthNqbV9uliJBWkaDE/DqaasPZ5WAxS
SEBbn67tNwHnN0BS3eukIzr2kv3Z5kfPta1EH+0Pf/XiJxHxsof47WQEBv+0b/st
ZXNWD898j/OlTFH5wCJ/Ab3oEn86XxjdqxpmvvQiKajpXqk0+8pCMkzjB85Ol4Y0
5xpcObnIDJJ7xu+veFCHgURZDgxXvNJNKXGCc5Kyu9poy0wl+ydpMwUrdhyQsO/L
TC/rnvC2nosmJF2lEQn42Rt1o9n3TZ5B9uDvuRqntAznrfLtjm3tAfghT7CxlM6j
CqggNDmfRj9REbLy4NiWP7b3xZCpmT1FitR0asLmD/Z+9E3gVoQT/psZzDVlNtez
pUbK8pa9EyN/jDHsd8ulvIPr+UJxhkKT7+bvLqcU/cEO21nwzDLnuYPKimtSrTqR
qtkshV0NaAFJUFeEwaARq6qZvbZH6ox0it8y14l9EQI0bz+amYjTqCcJXxMX3IUI
DQCt8TsJQaQvzsuG5ynKDtiCK89xFqn7eum4RuFOJ7VlTlbIxMFBD81qNQpXhzkV
e4gqVErwAMd8cD5KnUcZEkgIbJQlXBHZ0O2TEeJ89G8mY2e15o1mFtfOwHnCaz3w
pPX5I+RBEdvQums65g30B0SFOCIKNnZq3BpDcl4zGpTnfCF6fv7kiYpWwMUjezJY
88F95ERHitxPzMzsBwBGL/dRa+0LLrb8D5w2XJXtZKjt7rV/NK6WHMztPFbqwFIG
Xn6HfXHO8hBo4uPqC827oaHhOl83+Xlg0GQ83vS645s8JQsPX/kBwmnUyPubZsO3
/CXxdXgQOZk5YdH1PKm3IL/yKdgf5eT2w3Iec+hduQVNBgdnznWHb8qoeoHWzfWO
CCFM1unEiMNZSzNhBqyH//nRm3o0N7bhQHCWjFKIC39elp3Ic2K1yWQM/ksCU0J9
mhsITvCXbu+BOQiEE1/JzGkNBBZzZ8vLBRbnI+W4W3CgL/XOCNPECx+ImsX4S0ta
j3sEdAepw02GND2TYWUTICllNDkuD3dLWAJgIY0QYK/u7+GsTlHjJyN4ZpAv8Goh
eDgOoy72VqLCatXnca6ftMEtaX76bN9Yo7MMLquQ1EfNQOX2gOq7PtekaA5ji18m
hppO152YfXZLBUSjjisSb3sxmIivYBwOA9AHuAKHT7v9z2oo61MgKSr4yVxDvEPl
dWH1KrqeQ+nBRsZEklWkM/rQgLwf9QdXm6bIV+98puXcmTPCGl8U9b13HInJSpYE
C2iF0uWqU7HI1dZnBGRfxKyjY/cZlhHS4LbqnXuNVU9FAelZBwHnvCU9jcucGD96
FaJIGX5O7Jq+odbxazfIMFequI3MqPCIHMY4TjPLMmhwoOo5F63Jd4yxxYduiSn3
QPrsDXuTnA1ixNcIBffJFCGujjkvvMJz0KQTEua4045GQW6H7grQxL79JTcnuaEd
XECSL08eT/by7I3SFfvCeni/550nehjJXHpGK6bV+rRNmkVTar2naM1RM7lbHBkT
VTTAdjXsLqCa504JndZsnttfmFiLJpBIdha/bJTWOR2U41egBUWScW11eipIK/xv
lOZSPKwV/hswfhbba0XRkvlqpzedTs35SqNQUUW8a0XzhgtdKHKg8zeiKVDJbIwj
o+eu5roygNZa4GH1CMomZyI9uHZ29GT+DfeozYKHiyE5U1/RIQVsbA1Xknrx3UdM
pFqOYHg1nyrHWl/IpLrWXuyFyDU2xwiDMO86w5T4a50/eeiuXoqJBY1cVkvCGqJc
sATwsI/JBM2cIaTM8zFaPUDo8JQHoh1i/mC/d2vIVCHajCISpvPbha8rhJJDUZkl
qaLxkFllP/TbmvjNaQZw3LMAFx03THhOFC5/irnkCpUNHG0z9nGPqOBGg9lyc+Ld
PA4kQZq1pTDAogT7R9d7thw57HOByQ3Ug5If+gz/WAgxJBsGsnBJp4o/T5QwMwL3
MgzJHX05S73liSIBdMIvHI5OSrjb9ygvuih7pPA9+AWSy/CDazSxgl5TJZ24a4FD
yEMpUnhFO5CcoIcbiIaZYxedzL155vG6sxcUS6iJTG6p67GQPgQoqstvxQ5tmgSU
XgboDQgy2lInZ0m+rzzJF/JHls9NTzZWCsBZe4qwwrRwn3QjwQcngM4nTbrenaXb
gJa/B8idPfhJN4cUy02xGmMPnk/S/lgR8l8R7UX/E8h3O92ec61b+shCD6mJQP2P
CYx6196xBbf+yO97+6+4WNFt1W35MHjAm+CLwuOU47yy2Bb0h5/D4eq8I2ZOr/Fu
1l5pWvcKL1YcpB7tyePl3zlfz0W0vllJ+YSxPXCSbO6Iot6UvjBBepY19551abLH
6nxcfdGWZVhyK5v435JVvFAS354z5pBtjj5qm5+b3maSMG7TNk7Ba1S4Si3mKze5
Gk2U4+bFrsIhvaSWi9+xDjWG0PVbR82KCUpP3Dp/rRsgxoZHHS8xCi+Zi8nie1La
uRV6N9SPQkV7KRSCXzg1wDqFcyq/vouwUK+mwKPfZemgT2pvUor5cxN5xURpPgF4
yRnmv80P3NrC2UGrPrHtFCZ7ELm2jJ8Vb0jmMERedCnALNKcV5ifTTIR3xFXTw2E
TvLKVRUZsZziozeT8Jit+j6SzGcQBJvQuQ7MIlfLvqPVtZ+VjmM95FdYJ6wcQ6h2
AgWKn2dy4AgTXtu2Ij9FV1QjMy/HrOtYeEjXavDnt/99fFo5V+zFBTtwYwZjb42A
ZV1BFjvvi+XXqxZ5AnGWTe3rK/izAxW4wS4QJO4Qyv8OGib11T7/mC9gRqvD+4W3
xvill35yodSHSHZNJ5dcyBUkOFiQmdhw253TfJp+xFtWlOCXhrZ9C6Z2NJ8lI5jV
PeIXwPBjiJTvRPriJ53Gc+61SehpKvjZ2Fs/6itRI479qmvwL/VKAPzUpPiEHz27
hnr8J96whuafwCeKrdEpQ34PENOtbHkZZS3JOJK/8UnRi6NYeO2JzsSeYmJEKq+E
0Ddxmp5+3/yUoOaRxa1WMjafMWWiGC7BOjL6JBrGuQpNa6hfi8zW3Ar4lGIY5iVl
f6E9UKddd1DDJVDloWuSl3yHwzpfOpV4FqAyrAYwFkGuppdZIadOs+UcfsT2RoZE
W5NSjkGqPU9w4pFDbMjY0sX93SbC3MhvbVuRqWatB2g3ELC14Ft9dC2hB1ZJo1ez
dm1J2006/jlbY5s6AlxzAE85MW0Uer+4lV4XrkSq8ZDQddWBxqDH/NaU9yixx/AB
ShVJipRuOFgi1XiQ97cZsbv2zIaJGVMBcWqjSS58+bEF7yYfnCrQYgcJH+Zz0oxp
zW0K/M85sBPaXlm3z63/Pko6Cag+L5OXrZHgr5uRfdomZH+ilaM+ajopSzRqjihA
S7+XfFZQAx2vFvA+Fwc/oJeYDfZO9vO5G54o+2cOEOg6RxZ6YuJlq0PcmJi95qBu
gqCq+OZNSBQoCOt0pBcPYNcBnr90uSaIfZKazoU5Lvdxo+2xRPKTdMvTHezsJz32
y3t+s8SvwLBld4uU+PhCOaf0v5wdQPoloXmDzF7Q5ScgukWu6l3xu5oZGty/ggJz
3lkxj4wccmPPWbzEVzw6H+oyklm1XqimG+lvFCcDd7X/m14H7HT2lHXAQrZoACF9
h4DCOCphzLLerUXv8Wj42hK5jWN5Q3qEEZF+0pUQk5RebScGr2x6FWBVoCc3bG91
9yTsygRmdh5UjNiM1Kp5YUFmvhl0uvQrMcMwRtonqX5eHGMQT6HdrI17CG2Wmhkc
GhGjCMzCXRuSFIzB87utIl6C3Ce636mouUd2Fvj4zBOHsh+Uv/3P1+x6aKp8VjsM
ODWsT1qGmWu2e4buapPtHDGSVzXbGIGmGE1/QoGCHhQFpMK+mj7+IxzG6OKlS/8Z
digQdRTWA+BdmBJbrOIKCPcYCtRwSmH5UxDTyfztS+unZdiXEwH9O9A8cB8xgOSx
eAKN4JyGiJmO2pXS18U9s1X5KaeJrEq5oSYuUhYWxr1ji4j44Np+xq1g2J2o+Iva
ko4xOZpJ2rj8xfzP8PnAr8cf/701crU74CQe4WCnS/KRV3/+x3BhIIrEDD9PSBbZ
atIOrdN2n7h/MaB2Z2z7PAQOkBwsXsNYeOB/uIzRI+L8Cl6pVtJFPv87D0yhkVPq
+2K4Z+y46+6XyvhY3C1GGn3+dwUhlnKqWt/7Kn3iznOTQr904AdbmaNW3+dAM6Cc
NmNO6sGCSc2kFkcA7H2doBpV7OaJ9pOfEEImSnHdjNE4W2I7AlC+yZKRXdHxMQlo
VtZqqSS0AHJYZr/aga91le4wXIg3vzAdVXwVVBdE0T6NmklZ9ZL75ZwE1VNn4qp9
2CWqWwtUFUkhHi68oyLsS6KQ99LQBTptAKVFrQyL/WV3KBZGujU2bfuidHESn2R2
qWJsW9AHATaCwdqXJcUXht2Hdnb3NtGY543edT2y5rkkGJKplLE9GaoHLlWsaWmF
NEdHqZ9z/whGzF/9+iFJ13uiok3xXQypIVetOAQ+CsW6r6QSor2NW1e0d07G/Hph
5d6c7ii2fwj1/OXSasV0n65uE8F9/6CH81t/W3Ua+TDrr7qiYvJ28HZtK4fkc4gJ
XRh61HP9y22KuxcPNGpZpf2oLDe+VnO2Dnno5jMpapqhlYZSdL9a9xiJVDcikHRv
EzfcmzrKN1o6y3NNRirBI6I+YmCxk8i4iibyj3wRBuwO53KYOoVdIuKsNkVyfWbs
fuM8dV1o3r3p6vIH8Dg8CjpKRdkCxMiQZdt4o1NbfyWSuyX5Pi/8XdRSC6KeCFft
zPMrSYLh7b0nPRLbJl1uSrEvF/L1q8z56B/frtQuuvmHKwq+t0Ju6E3g8x53KQzh
qNGdvdSDQmaFmgzGLUk+3HrJfkjSy361arFHOlrf/08Dt677e/0VEnWUxdaFHW7a
1OKktsQ7sLn1o3bwL5roTUMPWMdnEfj06xUc3v2JAoxtRHcPnBH9meg0yWvadvuY
ILl7Q1kD1fm6BFsG/HN6fBChGf7Qboj49LkGjGYBZn+ENc90BgUDE7hVlkXpzIEp
rnaNK7gT8sA6erCUZnVsCzgHiEjhLsHfMKX7lzeuUITOLhlU/LVbmdG7izW/W5I4
TCB7ONc3ASMgieEB4yd6lAsEQJuznXuUBAA/phXyh3TMXVXVtU3P5Fh6Xjj7gkEM
E0Xu1gVKF7akU/nSH8BG4nwH32Ss+FO8lt9JhR8bLem4TbJi3EYcLvkhEOp0hn6h
gNwySBBdnCWuOrmfgtEsdEUCx6QAkmFmWKUG7OCq28fTCM2EuctSEo1+lOdt4Bm8
pGMw8QAKp6RWeo54AFFr532mahGKjliBXKeo3UqxivD4cD+dgUsBDy3/yMJS6K03
vxw/2/H+6ceFJW/PKPFQdXeCdPE/kpSdNRFBr5+X7dtlXphp50xgjanW4VYUWBwk
8Pwvvjl8kDkW2e9y6xtSE+Ji5muIT8RYypitucug9cUSKy3UglJH4vd1/s0dynT+
U5IxEQiW2tSE/+CkAnFevrxFkB3OwfVcKCbEgVXxlc6wM0GQNr0MHCxFfYezKfF3
NVGqgbnxbM2FjQf1ignEsjftSy1vzsMwvidPmNzVaIgm5xlA0+lugE3R6lofKNco
vJt2blUrhG9/Kh8HGlbVXpYdFzSOKAnUt7yGNzHey4pW4ygS3l4ZzwGLVAflWllU
1ePBoAB+qqs+U08pKmZ3gG0gV9bNYBj6OQXzxkg3yLAldMfSUJUgEhDhilHm5jsm
g199LEaDHR/KcGkNVe1BTH8xIWussIg7tTKfWqPHxmt523bh6fdVd1XH5N/wqMTr
dUKFH+K9Unf/fvT1iqZLH5LyO6wml85DJPExEJbLknzfnyIZqNMBC4r3eLexJM/M
Sn1l3CtJ/Do5mKqsNmNQgZDNbg5qVsiD0OTMnGY53yoAuPLrN0dxc/+brltjphPw
vaZCB3ce9IRIZ4RGcgTvTIXH0VtGMZjpVrr67F1SL0EyscxUMgIzoCte6pnlEYgW
SqCEKbmQPxJrMe0CzALjaVA3bh5mSAmb0hN77QoNEmwkoMwMEqC/KqzWJzHDnU1P
UkcT1UWSEAXilLhhd5PHHvTLspjhd25SUHIsRB2Y3xu+XJcamHZsBl7AOrWKYhvc
E8EUkbWTix+eXLMs7HybHtn6Gxuki8b1YB89Trl2Lx8Stv+JGjxw2lxRGw0FbOQQ
yuRe29XMakN+17xKN2L3wbYTZq2hm7VwO5ap08er0eam+NNV3f5iJ1S6jvxJ1joE
a8YC7G/QmNEKutWwKg33sycNEOpyCgnSNDpwDzvz+gsoGY8ehdDXoOarc4Ze6oBM
JWfE0XW7XEcCnJDVqFNAyyse7yUStEd813HQ6QwmwGHqL+Ey008dai30stLIsjje
QWNITLJfhROvB5Z2ipeYUQcXAq5U7zDVXpNfBtjzrASAoA8lMrxImIqo6fevqbhc
tVkuYxWxRcPSr85SjNB6Lmz/x4Iko0r2mpo3F1NQYnA1vkbRuspk+E5HKjLOvwhz
wmEKVV8YazpgddIfISTWckUNMV69P9rlaHGOEFWP/FEYq4Xjl6axKOFjGFr08jV2
7dBehxmXybS7534wSNw/9J0mZjQLngzUh/w+wIs27ZAAlLmz2FelvBDDqp38gSiz
YnU9jnGCd+BNEw4P9UNb065iRrGVk/MwrNJMNxb++A6FH0e0RhkiIU9EKw4D9rff
1B8Sc/Z1OecUr0slV62x9vuRM1ERnaXg1oT7OdnloSVlRMEGD9TtDwEAngfmcRTH
4chTHnnZa82r5CteMOHItOo7ilfVLkLp+L4vAIPze2AMSqCrGV4FQsNuo7qpvDCb
Fhqjg9YvzwZEs2B/seQhA9LCqoT4bCIIV7Z8Fi7ZyS2PHJtKCmsZpfcHm943vHIn
sCux6YlQBB8EBl+GkrjpjrN9oZnf46goIIpj/Yr7LzLoaFuNs9NMF5Ek6izJrkV6
QuO5r4Ddux9vgeEt4MIHD04rPzF7QmmPBdpeK9fL8qhIFcxtY+Udtc/4yYfgmw+9
DV7hZRewMn9mJcaD3MHB9l1O5hh6XHn6umtAcVTAcgbBt3MDcHxDsBxZ2TPClTkz
XLl4HJs4Q+A0DyMkJoOE7PClPJzZJN6AZzBDCEeTkBQ13ULq6OacsQKz/gdRSgTf
1+z51etjxnKZ6gQf5b9w7W9fgmeoirB7JlrQ4PvsIcCVeWN6INsbIEOiDtXHjrME
FG9DjleSsW27lIBbVqI3OV0uReuGRMyT0RoVbdtLYGzLDDOVqafhX7WNAB9QmA3y
b7ku62X8pcpRPFaJUjFy1vzyvFnYA1CjSu3IHjKS7nbk8w7UcuLfTfi83KDN2zxx
cRj0wc+mNasbhZ9t//kXszz69QePnyQm6BjF++kYaRCO89JBMe5ohOnynjwtPZSR
RK9UZ4TTPhmn6BeZPY1s7WSFpSVZRPMS3cuROygqE/Wml8xrAu2mBWQefozA+aEc
`pragma protect end_protected
