// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dMz+sz6m8P4xmLS4dE3AOFtE+c0W482OMelYo0YcDnGj3NzCykVn0VpRYJAtYCYF
uucyaFo2K2An9UdtZxTfNPHzwsMH86YaE5aP108KhoboGKZEvKMKShaCeLzOHNIK
k6FqBby3LErlK0nFi3mabt1zDXHe30i0evGnoninK2E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7472)
a7d9wEU68hdXjWH+gSBNRzZY25q9i1bFI2fCk/9Lmas4d6VB3gYFTCfOw2BkKyv6
SETlkggY0tIwhUv03TnyKy45jXw725IcEnZErsx/Ba/qxVH+351wOCuTVMiFIJkN
8VTWi8NUzhBBUYFQf9CtSsPck7PDh6gKCbVMfrJVGL0nNyWpvTsdFIea4+tnQ9c5
3uIgptpolpBbxrgYwDYf9r+eUr0a553iHJQljvK6PFcGANRc6c3GyjPi+BG5q0ww
rm9hEvJAyXD39xnRyAO/PJXVMPyMYT1RoMo+d+jZN+YDm7QQMhnMUFn/d9jdN6/2
1c3kSWcDmAJRiRQSJFhHe2epwZk7ckNNrInR/udG11tFGaFCuPkjyLsFtrb1s3Bj
PbcZemJfldx3jFME9EZRxLHXd/Q+k28HLeN8ZI0fAGVrXQyW+0UMzXiCMOFwkrX6
zBiZ3M+f52MbYWNtQP3Rhn/LYPKYwLAtZvLCVvnLfbI8lEqCRP2ETvMRrowbsgpC
mAC6m0hAwhOcr8Hzqh56pnzFrcAfCe8wFbM4+4EdI88rdGIBfwzCA2MmSFVag+Kv
aPv7vsq0v6ZEjbCi3bO0sirWeGkHyYwn8ql69+WhzrhIcnl06MIy74426bqR+EpX
LMZeHv7cvhAAvkUTa97rFtdJ9FRYf60m07KzbcG9Fd69RNffz+pF3lX26XB5KutX
TFBiT9erJ4QFho5NCMRSdbviGSe/+yn5ZSd8sz2+07djmtPmbF0QnXMQ9IRbKo0K
6UeVKkC4dImwToWyNS3f+YPVWh7mEbfifS/F81xjKMDNzBhoRY708gO4/Osltwyg
ARfoUuuf/rA5En9KcSaM3Pyl0pTNRZ17r0r7qfteZ44hdo7GlK1Tbw4Lh1Cb05U3
vHHipnR1Vkh1opxakK05INQ7ysVKVd5ODYJd7v/t30VzARYf9lYuNWFuhRk3PPw9
AdO3mpETCfE038IdUsG+6mT6ac4Dh+ByE1Fc0LlXVB66hovlgmKXjGXQ0K+xAnxs
eluMzUqrMijoZ10d1LACvOL9A0CsYuCavERrMef+P5Zftb6g+uXorMsJ768n5ECo
3xZiwBbZExySHj/zH5cwwV0k7MG6OHFivPGkooiq+TPT7kWh4yGFGdgyGlTnQQ5A
oKQcI6gB4ClOuKSmV4T1oR2+n/yFdc9glDhP9cRmU3JkuXlNTXuBhvdqGqzFBhNV
MRBQBASXKSIqy4vZMkSmsAKrGZGVjKVNHah5TrODdHryhecEscq69axvUM5qDo2k
3HclU6L/t6/BxRod2QeYpmPRbh8Q+ksDdQYrHDw3WtJxWI/E1c4/gLgflp9OdSPW
0a35LJLN1mdc6r7rZ5KhdKBYJorS3BiAIBzMZ16OfpFFeDwv/RuPea/FTCMv3n9r
yKUbvQJHJH8o6O9mIrgwFl9mMKzckDAmYY/e2ebx+lGXDShuQ8PH9vn8GDBxMb+0
gZwh3HjSEIvHYMqrp1V1Lu7lc/B1IBxwduC9hCce51uEizTUdY6bqawXWx23hXz5
srUordZpyErAnX2Vy2sBxys1HoFY73tTHVu4vAa2HT/TeeV6ff3Ag5i+SVjsEvaJ
JzHGLN7HIOZHUGaavwGfR5dYuzTDhch64tKSutkxS6MSieVsa23t13n7FGUGF2YS
Xgoi2B5O7xQnxgkTF2oPwrwy4x7d9zHu5d+mutOpckqufj8aUNfOZHhhJ/IlJACI
V5OtAX/dIFr59XTsuxz1+hlcPn8x1jik3k/c1zg7Lv5P4zBAgBe2x1uNPABIzmZH
bq8anH172pvUyNfZQmxh94kHt+tsyGyBRBKmijVp230omt5nJFuphThmBib75j/8
L7dTlWhjdBQaP7/y8kDpw6ypEEcqL3iFEVSv1aF3ppOyxY1r234JbCO/C4GBJcNu
DPHOEpMOkLWlaU9/vGA7p7YYvEpfBWETrHX0uM5RzvoxR6i5OVDikRw+vTqQLtki
xvSs1FN771ILuTxxi3T2hzLLpY+iriYFlsKlPJ7eXjaE6FU9w5MdN6CguRbhQ+be
cCoHWlsnHjtIkKRWIhekKQiERxktsiqo9d307KnZuo3/bfCcI5zmHlq2dPyNn/9G
ScPPZwciFIhwGS+lm5Vicx8TjDGIgfKCg9o6EP3LeM/DIa8IdKNv9ho3I4b01GQY
DhtJlhjkn4fFJMho5HMKzpuJLciZqWcF1mSaN1GbkgfQAqhRasuOw3Lrf/cW1zq9
VXVTKKjPyKYwML74/k0Qg21DR8c5aogTGYLmHmgfhmf+l5kogUwWyNRT87LQ4Ozt
+8t/rqt2AaZe/DazWVmpSF4HjMoU915eNG2HNBNn5rAbTM9BVvu/jXzEzZIdKMaj
WqPTjcFHWlmQczj51hTF9cNkLA1r/b6tWKG6USTklNF479cS0W0O7qIzvb2XlbzZ
L/a2xBUzqFHdIn6NaAXwzEXkd4ArOrfmJjCxLRkCKfrE/sewrAg42RAsQV+HZiYA
YnizgnBneww4eppwSVM/gWPM+ePlkd9FlG8xyJY+f6zSUP5nOVbHimJcqTY07ruV
dw3u45+Qxn6fTohsf6phW53i/QV7BX3nT+JqO38sPujRkAez6NElJi/TNqgF4+sL
oMNTmAvhhudqcnCa1v0Vw4K+ozZhS8/tE3d+dUcywL9E9Gc3PjboD1y4+zs9cIx1
9BTWl9XLHOYwsi3em0PuyHuz4Yu0W3iuxoWrS2NutOdLHm0WLJh/QelghzWoiZbd
c6du+x6d85kAZr5pogCPrzWd/q5Ncc6BxFM/bDwh6smgXaQyhw10mGOEGzvKAYIJ
NrtNEm2a3MSrN6+EmxFBc/M0K7IBs9Wdo1Xm4EJ8aj5MHamTdDrsLJ4jratTyxcc
J/htRJ2L99f70B/g0UhHsYAUOPqGxcTXvtlSVIgSDG9xe0/z2tcA3Jc2xPQcatVN
EKLPFxf9S7l/f2Z+JU+xQ6IlY8rDpDgu9gbTb5Jm8YmIsvFRYHJbZY4wSw8izCaL
AF1BphHzGRGjDuJsyKo/nSSNd+EITIpH3+H+yk2eFwlFO/T8lg9p04nY754VmaLp
R+UVlL1STF2LczttUj3qaJPtnYrfmSQ/5vdaW8nsZAekRnoSQ0rRFxfu0XuRM0Cw
Vxze/ytQ5z8NlmC/miqPYh+rihcb/EDpZulWJ+Jdkr9L0NOosZy0ypavIG74U876
4Ou5oeZFVY6eNw8Nxhv8CL/N3kJLw5184F5d7RoZId6fDX4D7GriTtuSFX/+zNR0
5zKx04A6Do6Z7zSmPdA0jVQGH6tpO64LCwdrHYGbXJnIN6QKFRh7y5M0qOQzHyDw
T3uebmqg1dGz1iELIIDJkPjLQf1iofIJDc3OqJkApwYwiMoLq1P5EWXsRAFPEOPx
hPFa1EbFGPh1Gyg9c8CFIM0q/G6ww3P2CnTaKaG12IlyR+acxo4UOzV7HqfbBqNo
PJbqKAKUNpD5gI6ugT/wPZF5GlHZGqiwEuAXWBUY6uzbbJ2QJEC2pJRu6EBdo+7r
pgtX8Yc0ZG2UT5IMSbMRzAUO4eXRRQAJJWrmOPgBa/PqkM/lIG9avtKLNcnnyNBS
6K+WmbBXX9uPxgE8MFOFnvUMUYHfiPhFbAFBw/idwa6oCP0QaI2aZi6uDhKBXHn1
SdRyPAD9BkoWbTpyRNvEPM8TiwyhB4S2RdGT/Vk7GVKvU61AKr1vb6ZP+xFrH//V
LJWlyotYgKw9i9+byk/rzveaZ1y2zZop0yAOOE3UcBSfOiVXsp5XWIUeG+oJZSJn
ulRjFzFsHmPcnYNYEEYcgetHU1OmWtU8xCJ6XI7Yb3vzG/+ENZJAWwH9lxIS5RAp
wHSEtk6jjIkptm0qh8xOJXjEDq4iRk0bnTbvJv3K2dIqYPEXoVPTNZeusUkY0otT
w5/iu1OEeH29dip9R0EZ/vD3n1gSLaJK0Rz30bnVjD9BUuSM5huyr8Qx2wfsbp+k
EOyfM2amp614J2aE3ITgLsv78CuYtaOpRsqaBcdUKcq5W0PjXoGImM4YYqX23uDK
O3ATwhY3EhgkbKhWLzeKUBc7YiCrPIdDqyoGWSyxr3B47fFUxIdNb1iwVlGdlZ9P
5vaecxpdFhJQ9/6ppGVGVi6GNryqyCekj4gUvdzqd3WNvujo70QTKs0+koKr10Y0
67ZpIYKimwIiXEaefmrFhfiIuZdDubE5AIt1kDgy/1BLc5ptZ0+FePbYEhXIQvIB
w06zN41qcDHuEl6lZh6Kmm0ZD8Eej5PhOIToaZyQq8K44mURq2KFXUtdt3Oy97sY
t/kDSNuBT9WHHCfDGcPAC88q0KMoFF2W8YjfL7nODI2qzjSTK4c8uMxedp6nl2pA
lNWt1+96OUkMWLxqO1K8Dt+OwktrRYRt4HUkJm+ABs9z8SZbOOmmt430uVg5L4/V
bwYh34ipq78CXcvo0VGf5cc7TQ+7MY5ES+dWzHmp5lFuREAgOrahmqJFvKBslK5B
AbDFcob11HyB8/V5XySWCR4I3XPmiQpN1iJaIJHoAT8wRJ4F1ED8TJdVXlJ2bVA+
bN08e2qZTS5Vnh0YFkuIthqO5soneL8rVvfSfpZUaiUKpTcL6RniOMkA5kyh3cqJ
TXIGpIZfR/lx2hFHWjWiidh8yUR0AYSDrm6egUT7p8iwda1wIFGx65QvoHo7Qveu
1CpDbTVyEPU0ZPFvt+by/Gm+xCoaeyT4VtF7oxY9HHJAdPcnJ+Yc+DkJgB6QJ7rO
qLJeIYm+9gPjUCK3BGLld72ZO9KsG0nkkZkUIu7Kmdo1zv4hOIlt8hpo6pW0RFT+
iT7cWNiqFvEmjWHlFac36/Q9mEsKkIPGStYnPyURadnP6l/brbdXSpB3UlGs3Jps
i09zWbzcjWMgLeAvJY63v3b6zcIiFTl2qTJLORMwSlsA2GCpMhKCPo0xe7yq0QUG
5ip3t+VbjdgSMwI0oTY4shUzWgduTmFeDdMy5e5G46anGsfIy+gQPPCVs8rdm9go
ZIx65RuQ+b4S47KvYVSa19Uqj4EO5Bxhc/H95U3gWkO3IIl6pb0nPCdXkeGtvqC3
PIFz9IxHswf+q5bySoHJv1XHf2XgPiGABjf4leYygilQQRUaaF12NUz2xtYrwApm
eF6jeEO74CFarXrnT5qmOr514sgBqjbfRTkMIIg6sf0JHkLXDrk1MGHpShKI7FgK
7DTpNZ9W1Oc3exA3go6J4niIk7gN9yJJAEFGLhjI878oyt4uWb50ULPE0UgVBna7
moZFymgFn07m1vGtjuTO84hoXYmrFRd67ZSpq+OYBvMYK7OTh05RaI0xjK8N3zD6
gqjpb5Ynk4IUTVT8JwH0oI8dszyMsIZfjfj/HNdu9bYml42BhF8Qa19WA8eioph+
hCe+YeU5M6G/xR2H0/VVogM8jUcj9IHeJCAN/2R5gro1FPbTr0JUnRLLYpr2UqHa
YAkoDYDSx90xDIs825JPw6ly0Fq2h3iLa+PnhDPzBR5cMoQ+IBFbavhCqAeqTI/B
zOlDpM5mXon/xX0btIoCBCjUhVN40/Ny3lMcWU33gveiXXNuMboMlBrQNhz2L3LB
rS3+HzfPOzML94O/kRtBIk1ysmTsz7qN0J3EqRPdOlEvgHDUkyFNfXJClcJmHV9F
rq6iwf+ApUqfE0JTMLdsJJ08q+KnaKxi4XZkNvpi4X+MBcBIArsaKxwEHkD3T09/
xRHvyOmbTHXx8qHRabcGmqtK07Iq8rQSkdm3aV2nAv6CXNdbeiWkIyMOJ8YCCJJE
9Rw//FzIr3ehHksRqG/57pxjj5YtIBgT+WaxBDSOmLKAmv5ed9xOSUkxGxwv5PlO
RsAfJMg+YcCJY/lyfVQHJXN/MavuSGqO/VNHYSJYh5fzdwepDd1fqsq8APCoji0v
fiekkjkWQrvvFR7b8wWVngclHrYCP3FWqax/qPcyWANn05LHw5p4nDTvC5CGpPUz
FRWbG35ddW4kKC3OWlpFiiH/zpf+tT4B5Sp7sxnXeAc8GjG4iOsEUNmilr/+FZVD
tbyDwS18gT2ts2gD2Gx2gD+lI4EgN94ePRyV89fgO8v6KE86ajp0ecDLWnv2qxWb
a2DXCqvqone40cdbQF8rm69jQ3CWIuYXfnKN9/FjgnUCpntLUsqzE9jexFTKNXSa
Y8hVAYpF/SNhr2x0SP22io6nqOYgeUyzk8WdYBQXq2bu/p5PDP9yXj0r68twN2/p
Ws6jrZ4h1MDP621UQElqRaP3PRW4VDG96yEuCWvwXkboY+BApGRIG5asO9LC5iU+
dCYwjIgE0emOvrM1uUhaNdc25zbB9r7pNoU6DI/6AfYJM+ba0TDB9Dt/X97k+TSS
QNVzqngxsQIjMStq89d+ed/8VYc6xw+2+zoVN/ptCq1oiC+P7xuQvM1O3d+TRFpD
GkPGZIUTGqlivtBz3/+2FzR7eL4O8Ff5GZugEwPVn+aWvaNeYhgkQfOf4T7pCkaF
bdfJtLRVzOnSa2ReLVOcRQcb9rrRlsdQjY12SlEkvsHKk8587Jmw4wpiX3M8JGaV
7wQk5iiyHNKkdHvpHkkGfhK+lU2emR3Ailu5PTUN+9xS/D3buvrVDf9aXdFNrExs
uwx27jLy6eosmpKdlFws4PfZ/5TUX6gbytYaFHgeTRM8L8t/x6iOxncPC6lyelxU
DYLpfIlScjsR/+uwt1NW5cvMERA5es4Zg0ph7994mCxMkifJrhDTlqrygl7MUfgE
JedraQlXmOqhWO6ZVDU8WBr+71zvvw5jToDPAiJrdcJxs3PROJXcuiqfJR2BPZfs
vivn3RuxilpcvkoXqJLTgxovbw2XXnnymO9hL6RHp5Y4Ce9vgqAjJ50OQtziEqN3
QBrT2d11s2RPuJAURlja/GuYvCi7ebIQxADhNTmtwnaGpP05wmjryiGVB+ZdkGQo
y2n+mvzZ29QKQgs6EtfMXIVm5YGW64vf0Xv1R9kaVex7VlXHdf9xlRAxDzlXBnDn
18mmfy8OPKKW2MHVC/k8cqWCIS7gMoUNlpkxzayisa90epDby04bhrF+KseofmtC
QXhCy/CLtXOtm210lkElmhKsNSDwpgOJZLT3cwojVC8Bb4GlSDdDgXeXFSGnscGA
zfpkFXSQQOALmAtv0gPYTndTpjiKCnyxUsL7yl2Ydd/bRBgb/pL0F7hey3RV0tcf
MXFP4fs/UDrDIT7jq/w6U/VHbMn0olJCU1O+eY9P6LsZ5NmzkS++/U8iSqDAfRN0
gpk/ckliT2Sgp3HwX4rT5D2j5J8Wl1bKCrB51SWvb7+ShZxOIOJ4YhW9V/D6MOw0
2WEmSNqWtO8y44ZBunlBOHWk2zLzrpiXx96sXp/6bd/bUtQU58Pyo8hnLbGfLeVi
qbnF/M/nnnp1Myda/BFUkNUpaR8A2kdRqKD6jzqJs/jH/lASc3ebl6W8XvB7BW9K
szExtJhCvAweqj2USdy3BdYiQZ7T79p2B8TEiwI9RD0nubpiOFnZbGcGMFgcocLg
yz8G8xL+rOUNIR3q44YmBlwEvgIsrKXBUa0SV5gdrMmueol9jC/iESozN/eUg6eG
2fElj3mzJqYc5Nli/65fTigWJ+MjNUE20JgtEdxH+rf/A8vL8uhlURj6AQDDztAx
KaK3e5zdN3Re7vurzhBIHIxw2AKIcBZK9ZW9AW+96Ugmyuv1c8FMqTyduhb5Eehq
9L7P4Z0+EiNtkV7vLhswGqrv0IJpki8ATZG+UjbRYmoowSHaT/xf+PGRFROvKXm4
SbwNTwPSjaWGZjplnOqlTTvZXWxiG9FK4ZWX9VSEWh3SeFju/mwN7f35Dg8dX30L
HG0U/MTFLLY2UlY6ar+QxSLH4PzgvZH1/v7UvHfwgLTAVnI8PQySvUGKkU41FjVV
BCab7/AMq6dqrjrMDglaLdoXA9Qx40z+7aVgiBfoCL+Zp9Z3ifXF2LOu9PYG+gNw
Cm76I1qrBfrocAt/dBmpgDo87lglcQ1Pu4L8t+6rP+E8SCuaaiqtYXcsvBq6CgOO
y21N+5gzOzNLuly6nGlHWKAAJjUiIrsLqjC8qiZuBID1RoEUPMgC0gMKu3Q+r89Q
UFIzZjKW9+j5+jEK8PHjzWEcFARiJ/x0VGK5fawi5CmWZ13mFL0ushxoE5qo4qSs
btS+3f3rxWrWVbW9vueaHC6Xz0x2KIuk8VZIj22fMN4fpXoV3o1eQMDl6DGigXD3
RH1ZdevJrKSwo09JKY8HnBQr9Xlh6GRuTCf6yMhGWOPpWWfRODiw0SG+vhV0yXoM
Pb76/Je6fO2P2buGLva1H1KUIduJgV7Nm/k7Ejqxad2kXS+mOlr3JP9WoJQQCqpK
a7daLjJKDn1UV1Mb8pzfVoyC6EGwMmFO0QGRw30UO/AiWS2UsZ/48zW7+jZaV3yY
74PPE6Ut4bXmCJcv8nMkipMAWuPZ6l4Sp8YDZTD29qY7jArlSxKuiYWRO0wtDHb3
TpWB/F7cNkYAnguLv1vYuIgLOr+wC8QzEF5WISJFke1sLynrH587+3H533p0my/F
teDm7rBqSLBX2SjM5r2d3ps4irDhpZkXmgve9BVToUEaQLUWwVyvn4HwNtq8tL1A
TbeUSmn2LKiWiMhfpi7gmDAPYbU6juGjMlDep+gghF8we8VYmlnNBbcRB+fIs+Dq
8cIK+bOGwwL/lc4B1w3HrH4G/m7jJcPW522VeSbSm1XMMSQO/MkXNr9bL7kHxOtG
ywJxQ/jjFvlS4AQ3pkTV9LxIxFGFykocLt7YHmFmOAjaeN9CXwd2ZuJD+5J39N7c
1U8XlsIjmyqIOy5oZfqoQB5L7iagi1zwBq3R/s3ddudkAzfKRjsBbwb9wSvtbviY
p0dZNcT86wwlIp4rInd8ElxPi2UTHVk3LQBomg52Ydq8Qi1DIU1mfX1H+hCP6gPH
t7Ws9yvOE8G5iUJSyUspTFw05MSV42dqBNlCbIAwFDQrM8+ZXHljgc95duYrxp3v
JRgk2jlYSMgC+cCCXLojD2ogbMQJR4zpAMtEoxni9GmJFA88ppfF0bGJ8au6LbB0
nKDDZ+/cTBDnZFii1mibPsHBk08O68I2gtnCAAdffD12j9M/myHwZyaG0f3T15aV
gvCG1nCdSqwuzL7m5RoM+bMwpanIYhWNWDqztbfYlQZsW6F+q5UwUNTSMndsDMpS
ODidZ1fDf96G3uBdLd9gphU1pcKOdBeIkfm+hf9f/Sz560WYReS3oqAqnBB1QVaJ
0wlKIDyZZpY14eLd0sfaACepVYO+cJqZAVM3L0rLCGzhlZTTfj5i2SQy43Fr5Wri
tY/pyiR/p/gCwKmryCQ/OOtFV5ggo9W7wawhQulpAGXaEfOqy95V0GDDaJsP6Qb0
KrpecTK9QA3f956CKrrIXXNYneBDaGheX5Go674rXnbO2ndhbfMXsQXKqysCt2Ui
1MMWc3adx5x3LdjzsCRIHfiHTszTNkFHBgL0EnTlCD4Ln2j/H7zG/RzmOvs21dd3
DlRaoReShqHkR41LQzAfhk9/1s1yJIRkZBhtQuPc0xenosTL4nJsfEnMW2h4U6Zf
5dyhByXfapDM0Uty8tDsBIDkDWMEuPrVGIu+VUC9TWyMkca9ffG9LqHSDX4ELUh4
CIT797BKaiTLJGUHJ4nT9MQuYBBbe3Cq3RthqTfo0IvKmdkB7NcQQfhU6D0MMGCF
LeNW01UkYWu6bkmJrSshyo91oa291DOOkteWk3fpRGWg+2vJiGiZEEcAcWQyVuFA
yNtSoPocPwWkehaYowlAb6IG8mXnjkWsm4R1ZxA+HeAgnk4BgQ9iH2/Cv3BonfDZ
HkzAMu6nkNIs2QhJd1JKWGNi9b19LcOPBS1uZFNgZvH29+6jObewtSL/x82sF/Hh
oh8sbcOAVUtW0n4srHxJRhmtRSgKRFRMTFsoDzUQUxceBPBaSEPzhJz0GF6pFRwQ
WC2jwjKa42k6BduHHkb1lqLBytlG0L79hvlYSn3ILIE=
`pragma protect end_protected
