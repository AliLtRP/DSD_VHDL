// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LtyEdQgE+YYXVNljpjpgE7nhAwOYQx63a38apwRuBDi+ATnEP102DmnipCcTH6m7
6WJSP7OYb4lYRaMRBqksPCa2LMilhNNNMoDfUFyQP7uzRCb69zTuUvH2p92zZn9y
fOn56WFwKk7vqQuqETftyRAxPfC5GaEtoOzHVfL9Sds=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9344)
bJSLBBeLuJ/p0PB/NrDaSENLK6b9nfDUZ/JZzKsKbE/JpW+ycIs25jvPPFGZddvY
or1x416wwW2CHZPkrB1Ivcw1OZfOpUc2Z80Kwe1rPelehYXjQtHbhPfUVtxF1U7c
FdPwKyvC5xA6Th1hEEvDtQ2fWDAln6N5bJDPkUj7frywh/7xtwIvPCM700gJG5Ci
TsgCfH3v+2bQOOFjNBv7u+VHFxc0m+9EA61oILn1DZgpsO3yKJmUEZhjMnUZ8fCn
ANwZHpsnU07gx8CGMJz2sb6uzPFqq5BVvgZIysRQE+bQl3TOfD1qm6TmbG/prEyb
+vM7rheQv7D4t04LuXclsPQzT/WXH4L7N0S20ceNMXEKGuqrNFOPkhiGdPkje1/o
4d+XrECM0ZT/0tLvqAnKNhtJKqpB5YgW67poB5U7MT58UOzv0zaEhgqg8Sz6TzFL
AUWjnrg7d8+k0YTlxN6XDV+i7v5W9aDCKdDJ1EwffR4RJD8dgXJFT9q6GhdpGC78
6P2LbEdcmfuoL7lrooN9Zrgo8ORqumUECna3P+1oCsCEEPy8cdkvbZRFRroyTYbk
CVf4sU/yIsTAKafKnsKTMBaYTtkcXU7JlmM529HJjfffI9tm3w6FqhRlGaIJW15v
rMTs8er4f2t9Wemu4BAR6VeD6YJXRojUGmksijh0CgtdLXwzF6HaK5+vLKMrw477
nPX7sGwHT1buJ8LJl/NppvS0HZlebwlA8hFhkeKN6wRFoYGKuhUAxILlOW4gVMme
hVVTbvajcb2NSvkpVWDOCHk5KbwVEyCwgUfjj/BACmxu4nw5r3JiUyv5J31DVEOU
RnPMlXn54hYq0uLkETqAsfiEBbU4E0RS+uaz5cb3btZGW6s7pIGaZb52NHQB1czF
SkP1tLG6PpfihwrZrhUjmYh6Qz2/e5d8YoJqlQnBf/hPDzuLR+SUhF2jYuYCRJ46
uidJX4bxPGl3mVIAnwvp9D0rk2zfmnwrOsEjs+4ilpoq1Oly9qCp8yni0Jd/T0Y8
XuzMLUmf66B+mtg/rSLpUvsjUkYrOGMw4/9KVwxpwSHCfeOHAOxx1cgWrEUuVtaX
QJluCs+HNn4vdKQIErff6TFMRxcmKwTCzB/A7UkNgzVazglTmOgi6OVg13d/qD8L
IMzvJ9PQmCeZSuvym+ZXpa4wNL2gsT3mqv3uopnSJ0rbkSAFMSx3RlR1oRfsK24V
9WLR51ShGSphi4ihDiDKRG2jG3c5t2zvOzJasdH4ctfF8SRm3wO5dn7MehjUK+e7
TmzTrMcSPdfaO7IIE10pT1myiHXQG0omkcINaY2pgXiwPlUBf2+jCqo8k1e2DRpS
wAQBdlp6Bws9Fy9wSbqQzoFh3K5rzkVMio5xz31Sl/2cocRdwIK1Yc2MSAu+Uh/n
LECTr5d0UCuve913K/VYfKpqncalxAa4EkWtuJ09+20Q5Nb2Vz5vOw9v628uFS3o
HLk12t3XX8Sv2s92FH/OLSkRtrXj8TLtdjXauiyGLrhbzaQY6KB6y257KSQ7UtzG
fPHiyjCfI7DtnZtW2b+qI8niZFtph/7WoEPZX2ttP5erIPZ2rtNOnZPUbssedNNO
d/JO0Ki20ISQCSuFpdSZEMDNog0bTa7v4c9nwacojgMNJu5RzLMNEoRXGtgNrJjq
ul/VhRhCi/V9xQNuTgHEZCoou9hH04guqvQxI+lSgD9ld9NWk4/UsrC+b2I052A1
R6p6TzjoP4tRd5sn8aXdtG3WSh0ItxUxi1LYflk4Nejm1GISdveLzzVOOEgXgVW1
vEVQBE6s/kwxDbk10rsvkbPNVgb80nVw1FNJQl01EQmAq7S0UzAwg+F0wlAs1ZlC
/TXCb3Mel6f6jYfvYSiAdMCPsizJQW974PNr4KVbuaDGCEQW3Vi6DgqQ4AfJhb5N
3SV/cPmKpiMbbiCRrLAWeNIBeuqECr+8GXpGjWGrlJ/ocU9Qg0gOh9DDv/xudOJX
PJ1SuUW+ZMkj0GUIzpAha4d+J+BkIay9uLWX3RddOcQ16o+AyyOAlq1SDmaAHLeE
o7+TWbyBobT6AQqU7jszK7cLTra/R+8jlAnlECaLKLTTLP9Xs5BffnObiH11ntYG
gFE8rSnP8XsWB90V/D/yW2D1bio84JurGgNCpxvrhkTfylLO2H3Sn9g+b8qz7e/o
9lv10WvUFkdEPhZWyuJslHMKjCkICPhxw8cm9DgNcteJS1bY3lsG3JSTTjHlThtK
89C9BDXpCw7ke3RqT8CjjnCteQ5QPl7ZyflrrsalIFHfxufBbLf0Zli0nXq9ktb9
aT7/EZ/Fj5gJ0CXkql99SMx/P/8Th+0seybL46wWhxvFJkPy4CqZNhVPNcyEQXcQ
XNcZK+E2BbZ2NUEvSCpqTcpfTpMriy//8AflkD2ANIxnwXg9mIDBICUb0ceAdmeP
wMxu2Q7C/vltbZiDb5+2EB9knqcqtXW0SCyMwPgAqFAcbh53LYi4eHwRZod3XGJw
xAkc5AVbV8ReoXKPmcSmWqJ9rAwpmUgiSFxOp1SNJbXBxDrFLs4/3uRo/zwTFD21
vXD5ACQe5t5FXVrNF99zUSoch6W65YFvHfBR1HsNjb1rQcY1Itw2nZolc9YUTxK6
0uiZ1tSVKkNt4YDn4ED81tx0dZHrdqu/W1/Pl6fFHk+stwDAC5lE6GrbgVZ7FL82
8QjpAc+lFVhEguLUspMXr83SFS/A+KCHzSjw5lT4dONcq08QEtVQJhkF3YEw4y1P
hgvK8J59R/kLj7AhdRJpEOi5GyH7UNSYjuBOjYxBcwwbTS01NZaDL9b5Ze7KEVq8
V6RYrSNtD25qJKTDGB5NYiAGtqQeyacN6XjWI9nMmqiexZtT+QF5BQ/B2D/bxNWj
uOa8BGsuMQAmRZ6UnAvzipmmuP/Re0xZPbssiy2xsamMT+ako004SHrhUP5gqR1i
Z9Yi5b+bX+SK/6eFAiN7y1Fl+OZDiHOJkdZVE1Ma4gSbB4fc2WIwS/iU4GRAQPgy
Ej6pVod/HB2O5HPQX6RTrqHazxdto1XFC70qi07YSR6ZzUEYsZtbSmVgXG+0vmCp
v3ZxR6shZwfsQE3MS6+Kb+4sLWl/5t1sf2jM77Wdb4K7ePlO7B5UEBJzYokSjxIw
M7g8lUWHekC4BcbU73lrtjGOdXbSzFivtb85qKQrdYnqEtR0cySIcehHY7vHYMht
rT4Ke4G3WeDP2XP0iEp7VXTz4jSKExPEnReUiqEou3rLW2HjC73AKbaC2d3qLaPO
FG29ZYIgJJCPpjVGaTXZYo03CvIMbO561Ive5ENocOtyZvNdGbb5loFwiwXDjQVj
xkjLPGdz38LlIBCcxZMOd3Mxv9h8VobrKymn7XgV0EtuME4wcDI9ac30zoGcJuWj
IbjZWHNechuo4xX7LywXX8q/hLMm/9M87agQ7y/O8BCgMYrEGBkrGvZVXlww9oip
1EbPYtSoti6GdCpOKEX6UJacgLYaWb9UVhNU34khtEgr0eycfXpNASBDH9YfLNRg
DTbcDg6nGKsIM1wdfBx80QA98MhLNTmIuukprtfVVsOXAwEuwFq9EMVHUoWpCcGX
D7+Iv7kpFshFSl2B9GeSyUNb+dUCCWj+CcNx8Q7w8IEzIuvUtRddcwwBOKI1oyAO
OJEsVP8eu3DfBdCRPzFmbbb2BhSdj4zKga62ZWXeDmL80THqLQrOErepjPGwQ3QX
Km0gg11plchwBwu3hRUdAk6m6+yUSaccqoZrEBYBy7qEL9he2wJNF8wXjFqnBIU3
ZA8qy4Jz7p6FFhYxVGPUFMLPNLrQwAeHyKuVLh/jbYkN5yoJIgsE64cmmPef4pSv
kATAfZUR2YOsR3+8ppIk1l5Xz8+mzmEmJLGAHqyJumCyYDu/wy02MYQYOjkN1TEp
hPmpH+2AMuRE/pEKIaEcrB/88VMUPB/awwAnh5StQVfu8A5ggUbnAaUL7iP9Msqk
JTsYLzTA70hRAMXgqVA2fEI9Y4rutquNI5G5FZ2hK80ezSzyZN8z4Td1Ehpd1spz
VU/U7A8SVt/ybxitjbk6F5OUGU7MksifK0M4jSNnkb2nPQYBNHBEaWSK608pd7zl
xnnltQEprovuE6wjDckTDamscsRtchV9TOGf/Bsxypj8SlOMPM2pp1IsjSug+D7F
08GNuvjDwuXtd5ZDgq3OJmgfsOpyvI7yS4UY16kBnG7NgxqbqvhgsSYRutfkRtRp
1Liy8oKJOKavI8HRdmpZKKUObb+SSN14BiqlXV4bhbQk9cxcny9m3sHuGbl3NBZw
vPS0WtsuSNa5EZWzcbg9O1SlUk0ci8StPctm5cVV7OwqgN7AP7r6Cs58m2cbK6sf
DCZsnCowcaIi26+q1LKeHzCfjx49ztrXcJ+Cgxwhjixop0NRwIMw59QHPPfeKQWi
nXhiyZiBRYQ/d6/okvoRKiEwP7XqSh+lGBY8+H58CVBjSZHUtt+SWhTHxVxeb2j1
ZH8FmVNlW8dnXVKJGhSglZj02KUKB85k3yexbu+JMwk/3luP758sAYRx62OUNK+4
+dxvKHJrQW0fM7x5fMruytlvBt2dEyg3ln0TPGCvJaAFDeVPPu3OhTpx4IxB/6bn
jf4ipD/6j+5fLAVNoVJrXE879OyBtqy/BITjdy0v1hVQ7EoUQOlTc4aVwKNgF8I1
y4c1zQg+TodZMbKsr94vaVj5mBaAvGJ7+MWclXXseqJu66tkkJzYKgVq01cwZkV0
CRuVnsE7D+0vP5ig8h3u5SlBAs20tVmxLj7kMDnvskscT/lkpkg2DeU0BYDNqs2m
l8UvKi3aLlrNRCjH0Cp8Dg0jASMs3JRwTiCZARDCx+IxYhpq6PtsH+kb+0WOuV0C
fLAahUSy8HnfqXu42kwzeeiF298Yw9qUzGDo9tZoqhTc+CL5hbDIxE9b+FGaZmei
d+FWPLjw70f/nnq1qSYCZ5POO2wXCXxPvlpnSmSpQXXDkFJe4B3sEBfhDov6Ul1L
iCw4Ll+AhCT4y4VGA6O10KcxN/D5Jy27OHg2xTgEWDYlWgXl0Gei3PiXXxPCjdvn
5iW09/rBBWmq3/OTS7HtbbxAFKdptWNzKQRsap0BPYBg8t3uw3iMrpwD04isSsMx
rFrfTVdSjKvECrIouKdFEPGEESqcN2DiCowzPYjnH8mbScp2+sKgk61JRqakGt/R
6hAyzUeoccFZNyUUUgIjNxu84cNqrh2c3tPEQb/WCF5GM4UcIKRj5UAFbtrFoeRa
I/PezECtBFQAfE+LdOnZ9HU9Pnk4bu8isbG81w4W4eKbODNKCMss/ncehrl4doso
sQoUPD5iBYkGms94rCQ/3Oly77JxqNIa/Y9nTzYo1Z4uha6YGvxODjHRYBIfjxvz
o0T0fgj8mJ+QF4PPg9WspTutoJnwDniizgBx2QVBvPVo0Ml6rhOUueynTsN7BGt8
jfxmJYp8RdVDPXNAjqZT6x/QRGzCouc8hA5QoMSP4OiYjo4Zl6KvQTlD4kVGjhE5
oYNZL3IXYClRVeYqiXQN0Rn5UlelJaymMa6Q2w4t7B3+3JChv9UTpY5ogTdwssfd
pnI8NBbSSrxNFBMU3qqk3w1NJel3EVD62IBBzsG46u20Axuqv1Nsmdx4w/uzwaLf
+tCgNjhbbf28rkfu3D46Bs9d4tK2ydRycPRYAxVb3ohS6TGtciidM7k36hyfosBv
lOsv4fZTalRUZdlh8dbewa9uE6lts3ZqpFDfaz9HrPQnKWL4bxBYcJWHSbvyc89l
FKlg1Q2lDLVOLllr5YxwtE63RYxP0MRCeLFwHK8rNotvg9r2cDUTAyY0hu/2Agw+
WAZZGsL76IDeCx3kemNv52bik61mvp9vKft1Ovg2lS6QKqgauc7l1nZL+OwRH+a3
BpMjSmwIWQso39S1U9RDcCOvuSeML7N8XDC7STUOUoNt0tU7ILR7ypZamvZlgwuW
/uo+ZGX07QDjm1aKaX847fvmNNRhXV+McobcXctF6qxfZ5X7vHrDDfCedEjs1FsY
4IOWLVLfrIRCxs+ENHL+DBo5v6dEglDHc8SjTquSqyXRfS+2JNQryXiMRjkq3xOu
Vumeq8M8NZDCj4e4DTUqd3uhYd3bvfzipigljNbW5a0Y7TV7EiZobfAJLHv7XoI7
EyuAOWoYxRlxyE2Se/ddC80F1fdQj470ZUNmP+dDvdOo9+uOmzCLqLtJi4L0QsX5
uUJq1cx1XDyucXLaFRBD1NbY2FA3tBMw23iZZXWjc5STAmgQMg7sjfvBi2nxpZFu
O+i/5XKvBhxeB8nkJ+kBhNYCfVqydgiAtSD1/pUxVuxF+c+VftDJwQHrIaAjx1fk
fAkg6UeAppzxnwCte2RGGEC7q5DcJbBORnUAFFf1EhEyT9zW2yVfrBkYx7k5AhIn
RBmPCX2n4NWy4kGaGRwNSLk2r+fEW6ogwhyBQbzKXE7ixIdhqEhLmiGM3DkDYPud
kWpePtfndxA3hCkxuJIOWZFP7yRaaphNKrmKuW7BphkxzS9alWd1ag28MHE9WBsf
LVlIQS+dkxDLORTtFUyCj/GWTudoWUtghpEnTFjE5qlRwXSvjeMco9/1NQ1nYvNr
MAx1kdVG1jUPuue1bQd0/NH89uDKYThbzLc9/gHF979pGj00NHZCJJFEZt+T91Cy
dWuK2myFz++ejnt6OpvP64Tp0rGY5RWSRq8IWFDwIfbvGGCD9QHE/lPxHbn1iu4I
zfbXqn9KdYioM7OXB1YB5uTjVU1pd1ksi+ktwHAJiwY8/WVzkJzc6DR+C+ogWHFc
DZy9ZOO1y+9G96fS+W8OjG4bPMZjl0pE1l9bgf8i/OrOYvA3YKJP2f48r6BmQ1ae
d2/zPn3jxAefiCdZ8xcXDfcNi0M6Gjp8ESbY1DRPTt7ZdqmEBfpJPibDjVY0BT/R
7WQdDafvFk5VN7iXGf5KHO+0nQu6FGReJOoodu1pjnBTcacZucHsi4/AklzEoZco
ehbIGExSVoPab4uI0G7H9Tu//bd0P+quIJl7R5oMbSkOrc1LB+ZvuwXW6ti7iDer
3vCIK0AO4AmmwmBpq6pObcB5LbFXlb7MFMBCyCWWy9sHIWfKVRwB0Xp4HNnbTDIy
ZOubSBjo7/LPXX/5Zz/wB7Wn24MHk/dODyz+1n7kUur1VI6Nm3PRtB01f2t/LuD1
K2ysw83tSk202KhMm3PuKBppNeZ+clV//OE2geFBu0t/+xeCONJYsabrrrqstGVs
8/J/aQe8hltJ60dJ698FyRO9XeY5yE+qgd1SsiZEiQYShGJW6Dkcez1QezRHJRd2
sq2hhErhXvfF0Awvec+rJWrvRbN4NRON6YGc1667IxbqzBtvhsZyiYvlJsI4m01S
WXuri3Uxz1WCggaXcIm2BsVUgpLnUw9PjXKavhxJJ1VGvs0o9uF5OmEM32J9Ekb1
fCS1glt5a81npwb7oixZ3RDNORuzE2JzMrFM0zHTVC7n8rlW6889i4yORdRsPKkL
jDsg8y+6WbetMLjEAMlees+Y+MNAA/sBVnQfQYAkf+Ii1oML1g/n2pnc2bUjdgT0
uJnB+rzFSGBN+I2xTmfhG0xcmrlQVw3jav19VqiRYOm3cU9jc+Ev9mX23kkC8z7k
YiSZTaIj8Jn6DvhVHAVgQl5dZQ+yOAGz4WWiZrSITacALhwvkEUwp32xPex8I3IN
P58Rc/43GPPLZdZkJ7RC0SZYOCNfwjav5HMPrYDOGc8FMMhmEbwPwdmq4uYJYxcl
bf/Xy+M1KfHmUGkXpyeTA+M/xyOf1qtLMnL3+aA1pLzDphDWPO4ZeQ8XSdRjwnn2
ImNlLF5IsHHRyF7dr1TsQ4mjkyfo5Xr5geV8F4Lij/cjD7WUavT8hqKiV/BW8R8w
svZnwXjWhKpE4Kzp16XmZ6oFso93DBGwHH9/j4TEZgX87G8whTAzcPhy+jUtOr5p
pf07cQ5DSsEXzRMOGyjggnFC7y0SmJy+oVSyOvzeOZmIKlqqOnx9zTbkK2ZMwtCu
p1ZCCF48S7UzNaEaQtaLqI4JiKxubxb2erWeLlXrtz2a67ZWit4ZCszmxx3gj7Rl
bomxUeNly8k59EsTlvvRKTgi8QN3CMSP3zDjTSRzhIpFhm8f+CA4YrOpZuxc5QyR
+vpV80eereagVFAODpWD+DZKJVKCdSpli5sU5fYWvYXVR84/GpGxf4E3XXxzKqnf
4S4xHVMiQYcFoqaRnXvCWzXvdgpuvUt0768Qvqov/8+vOJ6I43Iev1uYkpun8TIq
X0gD0JpNevmiL2l8/bM+16zqDQb+RjDHLA4hnG4v4XNOH/C+gTK91oGCIQjgpMY+
gKFRFV3sSRTB5OwpJwZ4Gd9mVvQiibVzVl9MyERSGts4yJlq++duaqIDEkdXaakB
FyrQFDtLPZxeu55bNVvrUJW+G/4Jq03dHM8ztIWUmiLf1puucmrB5pKaT6OD/i8q
WArcv8ueHsFCfp6/A2uHFR9D1Gocy8iY/m1uXeLWD/GTlJdR8aUtvbYyWMBLlCxN
Lg+wJYZEk4G4RhkqBmwqKhhkNB9u3CuJ3a34d+srSMVOOoegWds48Sxoe+Ovd5n1
xHoZovCDTvmcIbGkQoMREi4TRNyOXazxP85SpB24JPSUr+7dEwD2XqSfgHocj3UV
yZCcdezsvzw72M/t3yztxcrKLmnh5404lbHYhvCXqH0hFs3vSYIZv1aM40q0KG24
VLb4MC9n0Z5kf4OWmL2gop4//jUQzoHKXIj/0HK1jrxTfBYaqdAYYF2e1hFdbXqb
tPtRQk+yh26vTyY1xUQTmG43fCJyPu9dJz/8Mq2sJRughz/WvI2K33p0ye/vs9ys
67u9sEkq8uRqawWqtJGLokowJbQka+GPzZFVHJQtuKUkG/ToFvFtNsgWLzzczLTs
4qFvHErLviewMDQeqY5F+kRqn+irZuMwieh2x0JKm6HPHQiDXxjVC4W3B47An1cK
DRIHV+BxG9LQgndaVgA16uycE/ULJaKBDuEU9MJE0iWcU+DdUen02xXvDw7zL5Cx
FaavOYVQXBf6MhoLc+dZzvskm1Jw7vrjwN10zQLUQEZBnShP+57s7ihnwxUIxALl
JXPiE5hxqkM6jh1ipXh7s4j8bPIq14W/0m56CEU01/rqXPkNIHJqxTHVjXQbBjU/
5apuHYkAqLRlCpHxbYMI8QajYNQOwXsZ+LqOn2XHq/9vCNC+K8GYjtFwxVao5WNZ
Gxma07XcZDwz1di+7KR9xMSJkazByaQ47kvThMb+23q9EcJy52NjwsRxavd4M5sx
/wD1IOQLsk9Obr4MdLXu981JQOhWClbMTBCpC+wJDFfQiYKGgiWcuPWdAdu8uFlA
YclN8CgVHyk6uHpwq3QteUM9jXrw86BJHQneXXRaOCIaXsbceYV3emS3HO+k7j3n
4VNxt6sIROL0hLschAAY0G5ixuJrL42z91Pt/47wWcITPlRTnF39uLInt5Zr2pYg
+ZHPnMaDu3YVy2xngHJ/aiGor9sZU+WctuCGTSdMouuW0ftDbi5MLBbnZORMtjE1
CWBfpZfj/a0i1W6zHHxNP2X6nZG4F3MOnANjfuzkcKPcxDPFxVFFoC0HQ3P0qk+J
IFNwVnP4iXKJnR68IgHQ4eQMkxZUynH6ElzOaroMhZh6XR4//iqtP6Bt96lD61RM
wRndji5bzYYPAhdIrW0YUA1kJqOQkuNm9//b/Ee5VtwzB9R3fGINTaABwuBUhoKU
hy+PdkMnXkLD7/ywzZCQFB24XOMjpvxtSIqugCG8urATaqHN969Y8osJ5KuYZHXD
y+DIS1Bf1Q7bx5dkJTOTLMhDHgB1+v08pXXXJLXXGhEj++y6kIaEq57NPtz4K6tg
WZMcf5UmitVH9lRFAGFN039nc1CJQ/+lgSuhvSkzu5I1SgUVvZU+vdGxamj+Op/O
FZAzEAvPl7pVW3TblRJki8aaFeZe2yy8T6Xx4w161mxl2ZFRerSzhbeEBYX7G0wn
q+iUcfCwfXghT0D77EFrefRj8sqnERZnR8rtwuT9pTDPt9mVyvzyjNCm/XPD4YeA
UF7WNG+EoDG0148ferKqZUpjEkDXw6211oycrxvHcZeMHTIgxQGyWdMkqrkRVhIx
knj5+x//eGWnQk/p7VCkfMVMkZj1duQOk5IJc+yjlm5qtW8J2Szx99pHPt/YnxJh
/6S+9Ia7GxU5JMYrW3ti+UKF4TxALbQTmIRf5qSB+VEpVN/01tmyPo4uH/y9Juf8
ArKYgdz67nB2NzRuY6Ouz4XFmKBjbhNoCIu6zomEUNAqgugzb9aLZ+JbZ9MPJXma
BGKoboMjfSYiOM7k7CbVddzkXU6+2VX9M3bP/dRkojVXfY3AwJxwNaz1dkwwhXtB
K6ei3URjtgl6ErQlh5IzKuLFViIgLzhoOVCxp2DA4ILTFbzG9wx0UFIilgKGlOkt
dxZxCbrmTBomlEfgsd4H35uHVEPfUdvdsFRWjs3QKJLE5oFqe29Pi09RyBfH9ooh
kFkGlNwBB2i2Zifshnm+kKfhJOFB4t4VC+bITnCS+vnySbn2hoFTTRJCeOI5jC4K
911KK0W1tMJuz3KdEaThbqVM9ARWkaS2b4kXhcPNpM8+Rc+lAzn17vrDRHMMZ9NE
rrhMmHMBeFmWwsPNVnGmWzG5O8j6ET13QkRDWodea/7oSbRLzxa1p50lAB2QcTFz
lJiGhB1+yf1kr1QADJpxW4lpNICNNXHT0FVbi5UA9nXcLXeKIzsy7Qxnl+vY0yXN
fH77DfA7PJSNRSGVELxy4TQTMX3fycNHOVt86jofaXJgkTyT0xiM5TOza9WxQmkz
zKL5Wc+JAdHM7UOBZ/zMdZko8hI8HV2QwEg/nGvV3cAh4+tFVs/5oXki7wgl9o47
00rGnobGyh78koD//gsb33oSSC1lgsytMBlZEERbgBstFPgP9GpurBtZ0XV2Mhre
K+Yppyee6tQy+YPeQNXYt5mOZCqUYxOx4C588hQAa7O+4igdw+czr9q0N5xh194c
ybPYOddhoD3AFeJ54iv5ZTj47cgJ6ZAA1rhsggHgIA2LtRbE1a0jFgsItJIydrbs
ZVtX5P/smvbEVWtKmtnoF2YG/hh8A6FuWxppBjl7Yasv31R9DROb5O1Sgp5OL93l
V9dPSnWhZ6/H+eVtlQroSMjloinS0I24CH28m+tKoLXRsho7nyymeh3KMOFtGTPC
YUpRgirG+O0sVnLY07XlmoYRD3dTbxyZ0g4mrltIlK9Pi+e93zRl+ldsPy47Fp7/
9h2RIUms/eu6ukqOfSgJ2y/t4sR8iMv7nuSoP+x0aToCzeQwfbWVpgMyef8H/6jj
MDW/S+RuyOHkU9Sjo3yy2pTnKtHm18ElrtxAGVHt1SZAwLGVBjJL669nnpchL571
Nnu2RuOTpuy2mR3BRLEGc5ezaqXKihZTthGT+Y/9Hg/9uhVpDWweuwQUssoguitq
90yraKxSVDPtP8vViTyTyN9BuUDjwO1UbnPdT8DRKNafEV+Mt7d9G2oU3dMywYXI
wGDwlyzTHotJhjCg56pPkYuzqn0TxkKWIZFBtZ6NaKFTx/927A9fmTXnFRsR637Q
blFLXokOZTqhOGLBwt88BkZQyxJll0OmHAdy+1nrNLRsHLv/ZKX9YgMSGw1DjDnG
qvRYrzAI2/z0Ipa1imtV5+WJCAI6PQQob8IDqsuOd9te4xiZeoz/8WfRBGdtX9Cv
Rv1+fVS85JKkv3M884H8QrLN62tx2K+KJ+yF1BQBwHM0yGm8sDsABdhuY696lyDt
0LTMQvw4dO+aCDMeim+I6APh4ldSzy0e4RHajXjqIj2XWgN7m5nWxEkOEWrTBvym
mLwDSeYlgcW6epnKEN+N/E8Xu56eqwWYZMUqnVfHFGPlMazqddAKERu/7cNrlSKt
UG6Jv954GelqqzebOULcTX/l3wy+r70u6kxD1XR4zK8ruSoZiw88aibhsjaDGa8t
aWQ+lp+zVq0PWOifOVuhlRx9o7+1GmNmeDiGbxPa70PbRFLub/ZyPrBpCFb9AntT
gidzU+cNYeRV+27dyfy5TRqUe/S9QhtyMd+xlnVSzMhLct1hnG0jWHlbkAkvrTno
2VE5RCmN3stcWeUoErdYilHdViehzYGiMv4zg8SXv11CAhs0F6dohOCGUJ911rUe
sXC3NpxOq5DsNgQ2G1d5TdGgF3hHKVF6PkcSxEFCWUjgfUoiyN2hRLDukQQatQEB
6iPtAplYKDGTj8TWiaULpkH1xpyrzC+Nu67fcX0XS4xZIUBnSbYWew7LeVTzGJoB
86JG8shFTpwAZpsE4sum4aVJ3/QZQyGkFP4VyxeKPk+BSqx0Us46jOyP1z1AmYPt
ViFIRjZd13t5Si80DCMpkS5sz8E+85jTVdQJnzSV4JkYk/0L7BXQ1Jo8+3I9b5x1
qmjNVspbXz6zShjxOh4+ONuwp1ycxUY8aUNHwdlPs7k=
`pragma protect end_protected
