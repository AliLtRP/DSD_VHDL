// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jKHzdj8z8atKLLKyBu8Of8QJVHzIefWYxKhBAEi+ytT7VboJGlllRfd3TJowZMFC
tZiQzGdRpstkdqN1VJmqw8wOrAsXhxD+O9ccf38qS4iYgT4DVY3Zdv9ntygpEv3w
HXKj/+u5NsrAFwYf8QrIiqNFt6pz13Um/Pps9E5K8Ak=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 39248)
D44K76HraRI0pP74oxyWFWvN25YrciOaWSwJunnVEdDMkXPqlwc8XsJI1+EfSUM8
z8Zb1ymyQwcNaEph/BplvMJTywvo7AGg4Fl97dziwIIjygt224poAyU5P+F+W1gL
CvlDfEW0B5xqubZDrPcBT17WDf+qYYXhrMj8gfNgWDFhfmIsA5zqma/IwjW/pp0D
zUBbt9FMp61ZBH+O8c7GiOGd78nAYU7r+7UULVCeVrKEh8QaMTTXqx9bAcU+cL60
MIpqZfoTdIKaClouGWwFm1h3TWkCIFlqto4Ow+Qvi1iRUpwie7tYjB1v4Ee+D6Vo
BzmOUltqdhm6lAUbIzvh40QJ+6TUrs5xyvWJUvZ2+qqyR+cudkTT6MaJyCGAL5NZ
58cxmGWLO6qJObgbpehsBoQTKMZF5kzqyAxuZXklISrM+6j3V7jrEM97ZFjS76Kr
hpQVLXotduH9ULeyGba3BzHy+N1THP/LLq5t0OJbD2n4vNl0H3XC+KYOf7EV7wAV
AHhQDsiwA/TRKunH72b1bZ7edYpJwuWyz61GcX81qL14LtMWHDCB56lPdvFngyIx
uV/iKgW+XaYBgP0dC8stDbPoKEwQ4Pu2WxtnfnTmOFx7/Dw9AkRYX2BZCLEKcKr+
NIm7dmw7XrruaB8yV5MU3Xx4vMqLwGR6oWl8ny4y9fvVGKis+IlMdHwjM6AcoRAE
Qz6YK+LMoms6/19Mvugt8geCfjUDe+hCTLHyKRlv35HbOfGfFnoMyyEYSF/XRNCx
SWuY3TLBYCBWNUckfCty4InEobMfezfLrb9Zw+tiM+CCN+BA9DzeXEsH0JgJvPSm
qQ/m2GDN5XBI+zaMPbL8/x77Qg+e5ZSmnNr2HxObjpPHb9RdOZNIINBNFNKeLSYh
bB/7L3BJC4C1lGnchyAIMwajFaw8K1Qv+DQ40A3jYo8Y/XNqES7Wb/kehuK3iZ0D
/y1m3Jc3pvL95SG20f3TRzGET7RdNQes7BlocqqGwunc96y6/ozP72n2mtRZ0v6W
EFDvh2d1V5arcHxi+5vJ0GmZUhjPBxv9Jq4U1EOhMu6gitfeXmtzkvnANCyh0IMA
qJizf+x+VwSoywjgU/jKkY3xyXl1IUnOQb4eGkycw8NhpSVbWr8KmopZ+3BREFSX
377usU48kO2/AdMUJ80ilFu9xJOSXWH8yl8LdNeiuWbaKxCMQHgmQeixaBCidi+j
bd9jMdnJI5oo7iQxPgjmLbqPzScJKTrvarahftX8Tji7uUAC6KOwAeqBL30sOWxb
Pw9GYL3QTDkduL1uOByiafSN8CkfVfHnqdKk3VHSG3N+96raiELRYXnrrtYQYVm8
RfO7KsMvLNf12qiIpdew6OHiq7wcQJKnG8g5qImKto7L4+HmNtnlQ0ZuhxTh5sr+
I00C1rigyetdXpmsl3Q3h36Gd02Xy1kyrCnsU/H/wHKU7jgUMBTYJn2GBkUF9kwN
9YSCtTM6tAmoK7e8FZcUDE2KcSnn7VTWDVI156ZnsmQ320YMoWBN9e/eVpsQLXxN
ItnqEMdOq23sQR4QNkKfEUgmgXO+HYq5H8/wsrDVb/Nd6TeA4z7+NEFBUo3Pcxwh
E9qJBlJIjUuN7AED9l/bXyp41DL5alKW1bgdw4YqzYtnH7BeP+hVfqtdOmMpdL4J
qVdKDm1RmQelk/H0yehDoBfR5JV5HA9x4LmO4rTJ/ZrbLkK9p4x7BzfEYpiMGpiv
ZLehqCTjR2BClkgLTTVb1vnbBoMchilBC3f+g84tXqO1eiap3ICsLgmSiYvINryr
8xxO25s3B1jJDI/sJq+DjPgGhG8iLfx5pzzZuaPXQCkAAGP/YhqzQdcuqHEsmVBf
H0PPztPWjDh0210a1gD/hqpq7K/TRGIz6rtUdlxdE8JOi++tuJrwLS4UXErn8fng
rP52HvyzRm4mA6tWumod1aP95puLTEII6U1GD/B2jdDJq8k5+HYWjhmDCUdbBf1u
hVIL77TnvghHaG7adQl27Mn9+ksZySbUeMys0aXHq79UxpSYTQ7imfh2k9bl/WB6
/mmdPuQ8fhLHkGan8GY0yrz18oek/kFaO3X/pwtP3So6RMwnGMVV304/tJB6XTwu
3zqFoxalYmmqLAF8uYG3luGJGJewXMrxf9ExB8lCXT8SA1l3dvHyRLWu0ThMaclQ
GVO2yoa0zb/o9wsdxK0V+xLAZswOVn2GBlgDBNsuxOAYagrb9deHl13xdSBcV0+5
42sOLL1wWpsv6/HmGU9OOs5KzGchqk8AmgcCfivphzWZPZ/UqGEoROrjS69a/VoN
ISUhC1rev8G7s/TIRvsEcm5kEt5dCMzEQme4C1hkOgTG8rvGf7g7zE5bEvL9lEew
4YqQCDlQJ+2zYHTzIFs0E3oeJYtYRgzikj7gAz6y4Ac7VIee1z2j7HnAjaF+l7ce
f8jveKhp+cC8zH7ovUhFTBRbcgGUtv6wxoFnsh+0eDTsFxnyXG8XWOGYWMC14VSE
GDH84P/vlYsVpMcP+9kIq1Le11ysNzes+J1bOcZ2sAEDeLCHh+PQIecHlBKDsm/V
ynvsYyZ9/s+LsLq/XjaCC88Gi33oPkEFZ71LfsfWAh3DZjMr4pXYDp2WXSjKZ45g
Yk5js52edaf/JRpBZUAffjThQO5HhcwCfNog/vVnpybjq6I/p5aL3KtxkfW5vud8
u3GmNZZrZQOvjMinUPJx+XBaP6Uo1V0ijgVHBdeg7J6zptIX+Va59y2iqPhpB31q
dqdN3WVq6O4Ud4TfrEFu5NhnXc/wLBIpR0jZ+J401K5KSxd1CGVKpHOtBdwIjbd5
74ftk0iyrpogZuPHiF3qkIlzPdDFu/o+/s064vcESCwk1AAI5IkKZ+iJL/2kd63a
9c1gf+pY9Sn4/vA65jl0SYnXB+CIIb+Go1JHuIOHxvtHobnOW6XHPw8CxkdGXKok
hsGzCrQ+phGi9qCdK6AJno5fihAAGqUtuGXQtb2fi5by5Mu+KiB0OViRftjPOw1k
xLkKHsNAJ8XLzaMrkyskJXRBU6cSsJnOlgI3yjzb2TH8Dk0f9ntnYpMeWt9t1pjX
/qWMPaUK1jvcuxr1aJiyRayUJgDmqBD5JQpwsmZM0bdE0rVI8q7IxdLzs/wMpidS
ImtgSwN5h7yxcm0Pj7sYUDiwXK4hh1wNXfv01M49CAVTYQa8J+cwZ3BwiSFS3S9j
eazLo7QH3Tog1iF2QlMCidM1YKg7vVOu30F1XKVn3uaI+s1a6akwEfZ08rMjANfH
fXfwMG2FWbbEICmueNPB6ORC4PY0q8BhTDgBI5b/HU3nsGk9blj4UOh9LdmPkkLT
4JRmDoyMmUiGRXj3spOS8y3KL4Dostl/pKbBVIPLf4pzzA2NS3L77NcEP/FMJmOL
b3TeN5xeyoa8CEPAVXAKYaTDdNC8oCnsJvrkEY99tUp8gOZadbGg11F3cQLbCXEV
jFVzve4MLm1DLQLTivEESNdenMeeOjDyQ5fKmU+PTWAmER+a/iDt3EaDm/a0dNUa
6B/po4zzYCTOMBCfqSwP0Jcb/6Or+p7y0UGshZgNV0eVsfy/guC7bQyFEJW5o9NA
5eArHT4Qkxgwsd8Mfikmhb53vBTXSDydH31SA6r2lw6lPiBVNdBFmPzQ7QgrhzJ6
JMZovf4xBlo3zMYVMh9jgXRCtweuFZDLyV0mT++D5as3GF0azJQlqR2bDzcxEKS8
S+D4uc6mT7D8a9p2ztV1+l/8nWGqSAZ366juQW7DyHbO27yEnOLama92by1FINhs
p7Ngz36am5xz0wQUtbgs48M8vexvcsFdEC++uNH+XPbsntNaBNaTiGGH0CtghCOM
W3+RAmytiFOOQs6i2Or1uWBpeS+bZjsRPUPid8b2k/nNpfyCA174DEgfGo+K9iqK
IleIqk4kPrWxO0zY2UKR+khJ2lk6CEZ54KHp6nzaU5zIR4cnRUyz+B94Jl6T6M3F
8qtlyfwr39ZOvULRJ0X3+b710lG/LFk8zecgSzdt3E0c7Ao5L/8cyPrzH1EOoO4Z
kVs7/Svjr51iuXvqslNGazwfbeyrNSKzBGraNHiIjFRlsOiWQLteWfzAChvtXmlQ
uIXjvWUkToLk+/qH/vUGurzpUQnRj06cENv51Y4PSVi68KGMtfmJvTa8oPxpYiUB
sQ4bcrxZ+5/3hJLmwbo6496DpPgvVcTGcLqT8rUvnNvwqWuOKMvC6yFFVG6glfVW
bvWNmH9mR4VRg9eV8Eh8ZgCcavzAoYLW2mW6KKPuyXIg426iO/KE/R/kGQQcXqno
izICPTUDEb/nUogjTYvnsaG9qlrs4kBdJamMPu/7Es+KrT8yc3IVWn/Hqn3KWf1s
nMw1S1EpPHsIt1eByvDnAeiOCq4nismxa550+Ao9gP/9Y52VY55wwGgzpUr0wYES
8u/lwcWxU6fUI5o0DJqvSUXBw+Ybhxg/C9yNxTo1JeUdRKesW+kYVdLRpLyErnZO
KU0TneNgYrtIykgYsyhWRRYLVtxqpDhFn9WqyfUH73CwEibVnXV+LzNbSbzFF2kr
fOTzmnjfNxnSqwCyuQUiZ7IkofEnrJugUcFx3AYYuuGKuzoVDWZLii/kFyfaietF
w/bss/hd2g0maLc2RhpnQKIfQrYoNFleJVl1oKxPhcFjT/eAudaDQvCq5E+/JMo1
SAgzq+CKoeSDgQCf1IFIFlynEM9gtkppbLRjGtI1XyIoJ3NWdhjPucHKaz0WwkhA
AOvQV+wE4d4jucUNNxQfDbQlWd6CIK2hnFBRs27ZS60tRoXhQaS4JLVRRkpnV787
o//upUHaWFrDsstvluJhP95AYX9g6+9ylVbkGC8KDiFS5suRJa4cMEachehXzuov
7M7ZaDh4lTHXCRs/XsXQP8tNN5tc3ynQfgpJa59Jk2OBziiwcgvCKeu66PAxU7V/
LfZNnWgHxGsw1vaHMWauuDqKXLK7+ShIBGJlCvSRRue0oAShFIDj3AZYf0RThLDo
/vYZi1hm847D4E4ASlWaoKarqqtJ/gt3bMJCLDBsAWqrF8Wr+24XVcBElIChx20f
PEfeH+iWZNf6p3WoKgW1O0JV427aDPNWYl0v606LO0lYG/PkwRci5ZKD+z6laOb3
fV6chToV3xyG5HKBU0tyZTVzIzefB8SF+yHEeK9eRuMVnnRC1JhFNmHim47Y9Pw5
CPduFRWXHRGtxfLmIFf/wgWSbbs1LMOuZc0OSNvhXWh+seZfysfAhYEouMa6u7P6
uUXeJPe6KCspkwTXdkTXH+FwNFcO1Q8dSMg4EhUSijk8Frzs2DtQHrHiJotSSedP
piLxOJELqbjC5E3D0RanUDBc0UJW9llGQM9V5c1M85vd7IIHXTxX3BGnz1kQY17k
1JWsemd8fvtKQ4BHG4zc8/GcQdGthLminwppSjjlhdOwTtA0/bHCQsHjbBBVGqpi
QslT1ncCT55ztoo3uM/MdsnoSevKfq74yFwsqCQssFa/soW4eqBmY1v0swRIaKhn
w5FuBwENzHOMyriNX5b+xXtWKjhnS5IyXwDhvdVbJDr85gxyUlSliC7exTdqIrd9
LsIAvyjEKL+BLyulktvtUhmwEB3kSGIYFUoeT+5Qm1CMDsRxpPNxO2Vd8WnY6Ymc
DYgbwz/c85XEqAzyAX8+185QS3i9gqg9I8RQPCZAyC2PyDeFnpcl0K8ejIfvRB9L
yFMccFyZ1q/l29nUC9VY0uk0pn+2mV6WFIrIa9oW0vTRb+rqXd0mPEX9XJFbF05B
NsFl0h19Wnj372w51tyrwRYJ4fBDWupYANHOGDHf3BZkS7/zzrox5fg/kZ/BZr75
72UEvhqIjMKm8Yslq5aNW/xWF55IDZMXVahtRUpWxAYBObEpi+uRIYTO5F7EdV+1
gU8Xb3IObyMnCrPszvuC0pMEg7ROSIswxhzScjdXRsEuoIJki+kciTfZtCG1F7nI
H+SrVppGtI+Yjg/G7tFPBZJBectZQciTAkE7rCHYUntnQSplLcKU7VxNLDMB8rqk
Is504+c7OsVmTD0UBFihAniZ7IaqHI0xMY7X1xfhUZR1VOyc4zLR62vTIO/gqdiA
iFJKDFYhAxjQ4NhMduPZy8WmnXKjBfc70wfuXqem3/gMo8toEzyLNU1OQHHBr8hc
IZzJXAo0WTsx3RRNGDjDXqt2X3jJPlZDNxsg2IDYQAaHYPnNqiymgBEiN/X624gC
f1UICaAb5vdp9vxwV611+6PoZTEGPnI4tqDbgAtNdzsISvPqHcPFYPlI1VFu7lpP
2OMW1A8nvrdKPHaFu1iV4Nk1OLdJ8vK7VIQc5gcCFvQBVUjuJO1qLiQxJAk+gVf6
mTHJG2w1HaOBYdkKAz3moo918OKPX85/YC+m06RGsfCN6CDkxklNWylqbNAcKitc
EgSN3PlxUHD0jVDVC8f7cDUW7dxcPOPq8l9sE0/AQ8P0k310h5WKQXJi0htCf9MU
GK8cyr99lbTfPwemp3WScDEuE9pyWEuAX9FcfcLfBY5CsZt5KRZL9MA/qMuHlq0x
mcEXrlgf1t+psfK+IpwI6MotgMW0Fdzimiq/GHdLn0K3yO0KJv+5rYtEtTZ2mbQl
Yk+aToyD2KcojuiHBNUkHhTEH6Velu7OPJ5Y0QYi5aZBQljSGyB9lw2fZP8JWfn9
xjahCDoljOCNkFESJkCZCQWuxdAKe91xwS0Pl7cZv5RvELH3tP3yeImWdb1Gd3oB
xA9qvBAVwCI5hlYxRLxtT+UnL/yl83+AdZMXq6PSMhZHxRyY0JPUEtPOTTt7KHZ9
rhp4zQXTXcCuleNrBlaonySJ9uknj+l3rtFwQae7bjkquan0t+6dTcqfWnYfmi0+
5bP7bCJQbutpmYJy49cNqZXMgYTQH+xRiRJxyA5UHiIavcuCYRnQFCgd/qeaPMl+
mG/k18AcaTfDgxF5scfraCzuGaPoXbDxum+GjU1+ya89/4C49XnOvtNTnAmRB6Us
44RD5KB9hxV+IFMczTM85xKn73j+cYMYQEppU/ujIkIekyCB3hc0NaPxPEaN0cXX
Mx0dS4jtJlhPXBHOVZf3CKpy0iclX8YLoV/RN/j8qLL8MGwQwm4ZgRHc1aL3gA9f
D/+K9/TkjON1uPd9oOJJyCe9CJrEnuWPEgTX2iarzQC5bYKiN64Xbop9Sn7Oc6DX
N0su5ah8wbDKJFpLJPIU7FWW/QSE0S4XAF0bKin337IOq6tD8hMG7Ev3j//fexAL
EQNwh9fqHstwsdrK9IcafZJgZLb8lksrIGJXhSBUQFHWJtrViw762nKDM1G0xfGX
kuhHOJ4U4Jertk6rODXvUWw560ETLZGunrXuajb7FKTwdf3lv303NXlPGY3CzVRc
iO+NPMJJkRFkN2KfkFfyBBT35fFOYsSsNnp17puJitOjnhUvPHAnMhVRfotDP4+x
QN7jXQUXDyGNEvZZgsYItpY4CWBUOpFEKZOZkdThGuB2yCuLW67xYrqqP5nmp7FB
fYV8vJQrn9krXMIJHhX64XBqayy6mprJUg725IUdVCivn00rJVg0/IALM6O0vaLb
R0NdJ23BqxO0FzKedPF3VZcdl6vmn0hozs8GzEqqrJ/kxA/HQnVTRd23oP0onngo
WaRfKD4zRR7Lm4Vfyg4UuXf8A/vFT2s2zIA7nCBcZxXpjEaZEw33FnGZwSIW+WWm
GrbQp9QpB8ix8W98oT5f5hxypFvZsTAfqmtKTev1auwb+Sef4gIOXi8SQoHx0anP
OwaNYW2iSzmsEKBitclQQcoM6ByGRhsOHKHGSYiJMZkaPck2pGkwdBVdMnsRuJ5v
hxDyQ8sL1WuXxCWIOJdZZWOjZWckzd0anFVJjvbN0kX0AjTst/nRDTkEhcdmIegx
9aXhUXBR6llKVR8ofiWXe6bOFyjAlgcRfpgsBn58GOOSSW4YzNzfZT6sP5sFGMS+
CjNplrSQaEL5OU9gJsIGmMWmGYf9RMtbp10MENGIfdSr5mvf9NqBlh3JhIsxvdci
jBwAnvCvt9vwsEN1a+c0rfCZZgqsZsKjEOKpOMvCN6hgIVDaSNqCB7eBbSH8Oq70
e6vGUH0Hg6vGC3/hLsRvtuqpr2ZCL2Jw6sKkV1xiV2mz5XT+WUR7hOm+oDJUyCTC
TuPxqJPDS0WDns0jb4D9g6fuDmtoL0hM+W984y0Lt4X1Zz8oHvDKJc8F2Qn49iB/
t1qRM8eWZRNz8BB9s2K/f7fEAhGJPrn21RpRrXFjQEBJqQHC3tSDC3gmRSfUdNL9
61/+bphGqKTV2YiG4s6MpJc7VrT2knRn8uICTRa9e39cB1gNfpJqVBe6659pXIfX
huulOOsl8TW5v0xNPEI10nxxGNVfaRN7CL2T85CvrIbEkRG9r5BcCz0AmQeyUsJj
Rr4tBolUd/AKxBvOi4HjbB6iwXHte4kWLKftfGjbog6+/VW6i0QJHBemUzyO0OVq
iTYsxAeB4wRBeQqTAxpw8CcdW0ZfdRQjy9nDvBMJBaaJFqr7niyOUfU1/+y7IPw2
gd/+jQo8wGCsFzGJTa9wNKHBgjAXhmJZns/QnZwVP7arp9i/UGm6f5rpSnF5J3lE
2KmwtJL9pYtTewIoZgvCk6NKEazRQKqKRURk8qCRfOa0vh3q7g2Q0c+xnQMfGRuj
xCOt12CxTFCh6WJUAdBKiqvKMsJRPwHvo5w9HDrTLFw4nQq0j6uB2T7J0LqiwDZj
5P5PIrRVxtkfv09/4MCNqCYmO6XZGUkjMw8sj1nrtW8as84rTe0ruCKTThV8WPkH
e5rE7fpZwuRWNMOvge38BrBTBN33eCu2Xr0RL2GP2vkN4d1Ir/6Yoi9bcPRPs3t4
2mA+ApVY6duBvtcOgRrVYmNGoW6itp4+rs/wOKLZSooj2zhFYhTEyFg3+8ubo6Cr
mE1HToZhQjmnXCAZ8Mltws+yw6iNBj0UablGjEy9nks6zkH2M7V1sgUysohACOQp
2CYQ/SxAhqYFOZjUmImcj2LwXJ9haRQ1nozg3M2ab2a9UoKEtGqn6kmQRI6g6/ef
826+jv1f22WWrYXyyT0rj/x9IbEoMDzAd7Uf3Y9UyXwYe/MnLmA+0xFq0qz8Wrz3
w5iz/WHUb0j0h1YrWqXOFBbxjKScSEx3wLpH//xLJU5fbnWoHrhBVCFmGWS/VB89
CxTTGZo3YiJ8zSBiakH9RxoUIGWwIfoPZROLfCmD5LKbx0GYogaV/hAbrXgtUyn2
AeHxs0i3eP6RR1OVc1FoY2TEpCj5B4OLpIqRthJJXzobHsA9NJNkBa270/ZxzX24
YOkNS+pflaySX35nIV1+heo9BvZhzYHL7vlKBVjZaGItqf97JAJ9s8QDN/0yQ0ki
hYYxntxfYeSVh3r0EwBHM0XS2nJXVx4VLd+QVxhs8hNKm4DUPz7FciWOVZQ/6g9M
P79IcvORk+V8teEzIIghjNmg4CkTPh5y70adI1SyJHWoHT3S6esZM+8P+0GcIjaK
3ki5TOKTNTvQijLqLTftexzkLc0wGGEGKzg2q8WTKB6uWstKGZU05nqj75q8GNEJ
UiMhAt0rjF4HngmoqxoqJnfrp3Co0haZWMScMMzuk9JPYlNfJh62fidOZBg+SflB
phXpXcJmXx8ehouQyQ0JyC5n2l44Zxq3CdTmM4D5PmB73XobYjQuKMj2yvyKcY9c
lsisTIyETQWkXOybJc4CwO6xsGi19tMkTRtVq4ZtlKJT4QdQo1klEIHyv6/IRtyU
d017lZD2d34Xx553aHJrKeOX5Oily5P12FI5F6iBFfXiHQeh43GzkpXCloVdFvQ1
LrHizmi0W47z0QQ28yrIEtyEcvxMNaOj+fILWcHsWfklDl5o0DjMxpu5mE4aIf7X
iGoK8W26Ezlnbm2EW4JSin11VGKSklKA1m5qtz5CU96w8I36d3xXKy0faBLFKvRa
McDUSmQCVPYqwnxkrJ7Q47QpNK5mcRL7gHQL6ekcFtd4M9OX3Gft2hegflqHlDZT
pdnbpammTRgBJmU6oFn7274Bp3eOhj/CVhDKqiKyo8Ouuz+Rm4DxdiQwk9tnMYkO
S2va3VSoTQBzW6g7AMIkw3QzLMuGVb0Wr4gH+/adGchGT8VRc5/GNK5O2pZ2jRR0
yzzeryfo6PbE8kPrq+nvaqaOa+KpGSYzGRGLdCl+0AppMJzd2C+Ju+XsNWuuhPnR
MWdQ7fi+Pt9xV9qam4Xpt7NozDyoU1cepNpXoFRzIeiNrBLi6QFDLCTmTnE/cbuh
Zb0nV1NcG1gQj3CIUaT0ACMODN/i19SPEIe4vT71Vjv0vu9QpBrQaqAADHkIxh2+
aNdNOZ48eiVDsa483O/NoKkkGvJ/ap6RtkK183DGgy3PEN0/OakPatr72/z0mGTQ
HTHFh4Cr0C8+TcrvFXYXILluwPJRrqqEXuak8I3gAu9W7lB1YQXpVRe53qzHINf6
wZbte7wqFx5vErZ4goSQC6cPi7qeRP0MQAXX34RXSPoVKb7OR2dQ0hkg1OISaRv/
RBfqyouu5Lp1dNj46Ixl2/ju0PfM9128xN37mkmQ1HXP1+RuvCpfNsMtyI24KuXJ
JO8FVijEZ6Ekm1cJMWIyUInLUljDV3OutNcMtKZF1vThcikh8AAnyuR07BrHf81W
BoDxz/YcvJRimKG2DixdJ0qyecfdSgZbw7aYLJFnaUHa/QwIprjEjWKOLNdvnru/
1l2hYDRw1x6aqOTDLe6DHUG0RUWqaibZz6rDqC8j6DplZEufRN6iXgJ55onmK4WP
oKn/ukV4CmOe+4IbB3tNBliuvkvPDmKFjD49J3jnI7C40iaLVsDwO+E+bnZUy4Ag
sHS4I8fH4lYjlLOaWGwdAc7NfUm2IqqBN8LRu7pdnf+fl/LFmp8L5+lcDwJ4RdY4
a3QtHIv85FJvzdo/+3qtu5AZh0v1CAczI19FZ6rwTDVshG3SR7/q9EgUOlRvRTY9
8IZeXAjO8q1HrrO34LPP4cuG2z0LZ6212AMHTrlxU273TBjW4uS8GiPrdwEk+lfl
miMkiyk9+cKHSmbsRPbAsIGe+y0jkauTS2Iz8qrWz6yPj6sYd5CC5BrvvQ61ZOtw
xeNBkMYVhONwpmIi9tDtHFiVcXCBh2BN88GrDuan4moThL9Rh/or7bmKxGCtUFpj
h2VVOTuvbuHHVZ+JGqdz6D07UiYPb76NzkNmwqjHXyLFS+fdSOd9NVEWVwL3OgmC
ilOkY8BeibhNjHR+kHzaGWfEqqbokK5DaGsaBjQv0c7c1xzUoKdUJ2I1Ci3YGBhV
K1CKLLgmGB4qQDQKVRyBUXLgeW8uN1QoVhVM6+7orOxzT9pvKPQYyCJ5TBhA3Mak
hy1E3L6sVCdSth8mf3vmOOBzh3AcYWnMUPpXwPN22MZF5DZzhFOzTPfVOqku+18Z
JWjytJ7nRfotLaZnaIBcHLiaxZydi1L24SCiWwPE0HpJXyzBtK7HGuX1ZJPS1kjb
9GQBxlY15t6udm5jghKJ8E17chNuVbb7tcq45n1adeAWULujZBDbJkbizw1A5Fd0
XUxfMBJDhx9LUJQDPcbH8dZgA2+zoXQj9GBMkvDceydkrmtieGmS9VpN+BrwFGjw
c16aA8N5ynkg8HUv+p0TR3X0YIo00DdDvj2psIF7OanbHXp2gJ2KadM3f0sKYnKn
0GXfZptfOWuOSFUBfOpIsT4J6VR2WblWLF2VoAxVmxGxw6f2HEcT3CDDD+mNbCwh
i8YMh1jcDKDEW4eb5mLgBS8QEh/PvSjgxmjD9nFS7eyEMuWroMEy/6rw/1QuRW1X
KWj0XGS3CUJYq3dYWFCfiAEbvf9gt0Uk7QPcRM3Uq3y3youht08M8rsvBprG3VOH
IR8QG11sBbYJ50MwIRZbzZwRPlfrVOx0x6NjGETuWTo3s9Zxxh8OdsVIQGnA+sXu
3f46Bo/0GPKWmESjwm1spQCfvJO3/3HECBJEECp+4WZWKXhq1JSohOS+8q7qNrHt
iLNn1mzRep0If/Bt767znKfD45XBGenKt66nIhwNX3NWPtcNMer/cLkO7mkg0+5J
qBpsyob8IVC1SXJymYRUlmZnwGDuk31CBV4jzFVy8cF5gw/oBzqccBD32ZTdYlm4
pjDKvlJKo+oX2R7KzKHY12+b4AnAq4S5kGSHhwHL7+MMfDWzpEMBywREhPdILnU1
RpPgPQAWAOPSvXKtJYy4eAgoJMYYzcsisL3I/X7FVubsErscnQuKDlo1/X+xPqtp
hEx5dsplPl0G3Tzpqa8ALxmD3thg4DBGwg0WbjAiCmrhZy2ImcJXejDv8yow03k1
bpsT5kYJIAAO68YubdXSsSlghTVp14Wnd6eupdsl9NvQKz7QIxakCLA/6k9pLViw
HBjouPbzy3tTN2bS7pvRNXUApjGLWKeId4izzum4wJtO19BmFuJ9KhYwzWrf7ttJ
7lIrFyeeXC9qcgM+GE+BfWG+11IwRAhXlm6/jK/me/y6ZpPRVfoxLKLFdPkPHfM8
kaLto5AkaNEfXVWJcxCkiktJwBvEHmBPPINP76vetoUBnO0D5s5xfzSLPJFam23F
6C7zfeip+oyKkDDfXVsQnofFW7o49GwH1V4e0TPpT7RLWs5R8RRo30mnD/SEjUbx
VgKcCp9Yd0ZpG/uGzlvzlRbwUVZ3SnwrZWPG8oGgiIuWQcOTCPM/Tf31CxFlfszC
4xWLCE7wVb4wDvOxx9ZwxrYV3ce9GnEQzKAWOPmUL1Ozwa/+VzvOnp/jUD2jxiqr
EwzQMivR0758GLLmEmPWxNb+vJXFtlwOrT22KZ1pVjcpb2i9cTvpC78e64n8mILe
IIlHGTDQGFnvwhhYYp3AK5s4uHtdEkSVCNijZprxQr92hVz0KhagZNTWSEItBnyU
DUfvmzuGjK3EWm2dztraypDpImqlauFYT6XA7Ia/h61CgZQjoPNSeiZFpbFfDFjl
bvnL2qDnzSywDiqwDuJn0mSyMZFLwDLQLQYQRqDao/Fdkl970UX8McASM+z3QxHC
1xhEJ5DCKUV0XOr3i+7yFaJChBaOTWqQXigQp3LrgelKnPtK7078leL1Uykf/imW
h6YLyvXTU5rpECecU9fCD2nVX7mW3/mxCMzhpB6i858YrRG0JKYMG35BbfP5sBBC
0MbOnj9mDb8Ahk0GrqFupRv59m23dTdillDshjHwwfDdDRD2/t90u/rvkf2wGgEe
qdWRm1e7Rdopedmt7QFbIX19efkdywB4IHmRN31Qt165+qZl4CXSzKvk9kP6FlJ0
gR0a19dEhzraPLNQ27jFzbc+WXic7g5iQ2k1HAfjnLloo6or6ye619z4OlRVrKLn
jEkAorTgqXJ/C+QzYw3zq2zogx5+KMHDxOqyl1whjfTTtWqvBudNrFZgBJ5CGVPZ
Sp78dUN4E8WuuIyo+tS47BN6cJhzyEzMS+2+9ABfkDvh2DHzS7ZpP0Vqr35Rep4U
P9eW5kgJS1CC5Cmy5IanBALUFBI9LMsDdj/eOQ2F2DziuFJbIjKYfaUGQDd6rNQB
EAI6QkUCAxnRCV6RwsVla64NtauQfSww9SB05yxa2zRQjmT+QoHiRkpOou8tleoQ
evwfiK0JoAsiclhUHDBR/me/qK4WW5SAE5A1rnMZzknKVbhw0XrWtvyCm2z38QpN
/E7jjiQRLqo1nHrrWfjtR7w0UhDds+GY71s0OgRXvD4KElediZOVeQMAEyWO0eOm
GUZfKv152oBapOYkViV+jStuNQXqAJrdtYEYGS+tbPApKxGCmnhxUBBAU3yFcGaR
9qN/C/ZkaGpxlf50zXrqmut5nX8MdvB8RNI8MOBXpt0jnKk8O7CTuAJrNL6awcxL
zTLX6DYINKi85jG/wktyKktf0ELRDbSPGkNha1WQrPB74ArZBIfRlYLzAsoEka6i
gOsK5gQaTaJi4ZKbsY1AMJzF6JM75iyZ3yGp7sCEm9SnZZ6nf4m1io1q0jJuzQ0k
8089GZOoBMFrha/RgIsAIbY7nH+9JiVwdH+2FdOceWtNjaKqsxdRr9UIepuxLaGg
MNdCwhueOBtgwEan77q2NPxgAROVsMubz7y5RhqzVEn6TnZdxAhk+R/383RY/CH7
dgLXe6NUrRHjrkpeQ9UPKH3glO+gK7HCiSgnNo/uS5y2+1oCx0NgpC9lR2q/UMQV
4gewYIpltxkdvNz9NAM8meryt9GyNYei0lPwbfH66uv2D1JDgUBflKNLQTkTap8d
w3etrdqwv5mha/aErEXZvxWUbI+Zijw0H9C5mTEJcYQZ3GHxJhq5EjC6hsNi7qaa
jLCtMfCTiDtdL6IqxG+rVTF/NRyYA4Y2l/2wCa3RKbSin6tfVRQTxLArrjoFKD+F
dH0Mj/ssC9fibA+wT3pcK9lRxZ0/FtvLEC7We6aYC7T/N0FYeme/vZBgnPUYifMl
8MccJUeE/7RMnbRtVtLZ7DHl3fx0vteynb1MBWXvQzkJ/9kWjgUEH4kA8gkw+pf1
efYuLSfaTAKw2BtcVoaS7DlnyLYEqSan1QerbfabvhRE661tPVW+aZFEsvTsLLm9
eyHj0DMIjbPCFleCILHInm/0HC+VBQZ2oCbJ4j6UBOQfzRCoa5OgPwKe5iTATUau
ksF3VYU43UnNKc7Lu1w4NONueNb2OBPonyM+VhOjFgUCHMld7SqtsfRT6uHYWX4Q
zitl6wQykeoAcONqFC9a0iCt8kl/QGIOCKbVD1Ucq6h7GqapXJn2ynQORcYHk3Iz
/LudDaPehCLw2jeYkFQmswERG7mW1Gon4UxsbotlJVGjdJfUIBO4xMr46KjvAreG
f6JyP7W/8HxihAAvIYulBn/FuG/csYFqRq+XrMcghYnLfy/kwSGMKBK0vSWQHWCV
aIFCiZORMCo6r3PqjvuurLYLKHVDkFg9+jz4DL1efBPbpyy0bqLAAHut/V/dRTPw
46M1c/rtV2F0lU+y2Kgwp8FcRwLNvy3IhsvUfTE9rjDi5noxgQQE+LZ07S/3STn7
6fTVLRYTFIja9qgdJatoFWVV1SphrRjNKDRZpLupbISOFu6mDp+Guy1g3NqVzIbF
urCCv4o0uQm3CJD3scqv4bTd0XTjkqY5zAg0Utl4IJt5gbFD7YgxwQdXuEwQuhen
P91bR5fifwAWwcVo2bFTlaeyhuV0GuD2kAP8IIbWeO3mn9F3Ehyc+BVnsdP4WHvK
PO0v5zjE0ovUp8fRf6dHU2fiSgs45o0CPBxdmGBwzmlnnsKB3eT3naMY0e9DI5LS
OiHa3ZsQcy40K1XFIFXzpoq+oewaiXMZb2gtFh1Jp9f6OiUCNeWDZJ53+UiN24l6
C10EWIFA+l+Af9Dakg/q6HxcnsHmoleZZOY7+GRGJL8ZjeV2TEZOZ+OVNHKQqYUU
3hUzSt/vYA27+pvIypUpsBStfd43VMhHclXHHdabVgs7DyGTXP0DiXj4CoNxjtbs
4f9oyYLv0bNnP7GHjj3yNB79Q+Ylye8zH6mlKjpSGQLTGKr3TXnDXATUBz1B6Qnu
nOJvyc2iJDydginBfmkTTG7Kvh6cgoQaJybLgBaoyOn+SoFbpPJcfSTVcNrYv4nU
aFH1+E8ujzuv79mc2N+w1VS+FusKm4K5pVsyV0dRQ3LAyNzGnHTfHDlLpRZiK27A
uzECgBSuC9ugmf0zDESj44QgPB4DNdq45md4Y3rh/YPKl4o9uoe+SfUrDCOhr2Sj
aXmqLFJ5t+r0v7K1848JE+ZhsAYoOruXwXj7RBDH83f1YCnYMq4J5PFTkGn/XnY2
e/+4XcJxEBEPmfEzkNjBZeS5H2GI8Rkj4D2xAMppKvd0QUeFuRzo7gOMFEKiWyUX
RXoUJII7uyQnuGope8Vibzycp8vDD0eLIfZFlgIs/HaiDqs3eUte5mVIcAA2QBxV
M9GUG7SzIamIs8ZT743PxC5Cu72u8jXgB8HYTVrsZ2nZPuQk+uN81Hqz2y9gtRyy
V1A2o/dyH7SMNS8/fLQvmGuwuYiE85rG7ho7wsNV0KBbSwHzxknPZfIys6PWUW3j
70An3hKY3IeQy0ZuHe4n0UHEoAxsZV64l5oioMlkxD7dhQ9uXNhzLIyAdqh1YTGu
mPfBVToUoRpTGpZDx7xueNUK7MTup0FjPxZanNhEez4ltl9rvMauBG6NYTolmqYq
foJk9oD9UcyxvUqeXxcHn8eNlriRCKth7KVct6syVZo8agtdQO83kS2hSTBnBWp3
ioraqqAGfT5qnNgG6Z9cWQHGkrKWFpqiwETehxE0UaZTu7Tbnvi5JIQih8+XXQyn
685cznlOW6LI7ryN4mEt2vsok+vHg4Cz88K9r/kRRD/l9A9cehN94IclTZOZdnLa
t3PAiNYW6kr23nT1Pzj/3d6L5WRxPrRdWKIrQKJHahzRr1Lc/eH+VF3yTrp1T9SQ
uxPyChTzQLgnY8OFIXdBDEel0YDULadm+lcQIaVIQ8h+gnYE1WoHZHflfZdDXN0D
MCOllGwj/nsd39sXugRy++/plfNNbMV7OAo0n5f3YO7BEvdSCGmVA8rBKexG5vm7
GhskGUU0t1F6Fjzdrbveugv0p4O0EukfSHCat+VDkURBtjlIzVqVdc2wLt6jacdy
8FyKFAlZ8mTr/OaJoKeNJY5DBG9wjnN67BZzM0ixDVjCqOX6rmcbHAyDhV7T+uzn
yPZc8lVlmjGbcIwrkI3l5WL4XpOuiohy9vUuhsWDvzdVhWTphie9YB6ZR7vAUgrd
6Yvtn0GDKrba5hsx4aJJ6FY/tsn8n+b6Wld09w0Dj+wKmfSc50eVT8DJV0FpuPUa
FSN6YxmHgDNzyLZffMu25tBVEoWUw1HRwZLhbVHS3icGXkk3pUgzmI4bB2RB0fDe
MQqFa7jimrhiBeLTNqkvyTzQZ5/mbWfQx0u4WcZ+uAbRQrRm4otGP/7H4sNcTIeQ
XGIPa8LMIdopc83FxDdCqiNUrOFaroP9947aT6yfGN8+wOpGskvA+CqjGNuQWaUe
tRacqdQzqdFrkSiifyabfF4D99/phooDFbTz+qu5xVK3QeomwolRFtnQ+VfVTm/5
nPynTSmiMMgypNs0ZlMBIImK+nmE2ZBWG6M7bvxi2hK+iJhaeuNOv9FOyvcixT1M
kUpX8bHvVb47yH9pf9Rezz72TMVQ4ngyCze1ITO6NNEJa2FzIT+4iZsFdXn8uQ4w
sz5uaGhHSjddHcDc8/6p9ECh0yTfLxPsIKjRfV9yn4jTbI8o6QAVzVx3R3Vq4u23
phN7IrL096d8rvb95u/vN/pH7pFi85tSbY+nLKbx9idKklVGhdyngAgxro7k3yPS
yMo51HWOrxMEm/ZWXiscJp2GoJujECoK80mu8vQpTQJMkZ+766AH8TJcI/9q0jI3
BXsKe2Q/hUoA8/fI/gd+q2kT5AW+xfWYdZwq1FoerIrkWcQ9kbjVUJQj4vfH8rwy
8uXtoY/HZOAbToUiYkBWY0b6bBN0A3C0L8G0ZZLwJQHAyyqPfrqUt2ABgK5T+sYE
C5pYW5GtN1GiRopkKdSZiLKgdvGONgASt9aKFO6Fvkn0QCmHUQdahh7nVHAdqyKo
bT0+MzHIed1gnObDBBEgRTwRUXjYyB+uUQ8emgTFpeDE5qomUjX41u3zUDKjvE2k
vzJVjUhZLwId5Celwt56tiPYe5dLhyCtYEtkpPvUtcdeV2UqVOJPCb7iDBaYvgON
r/8e2hH2tzPDR1QvoLcTJrI7wfNIt+NhYpQACMn1bdmg+5q9k8XtHMLq22Hh+ek9
yXrmAM6L2TBjkvjbhzCpb7Rz8F9698TV98uIDjp7DrdpVt1K2nzNrskpzLBt071t
lDYHbfh1Fx+QRNI97LcezyDGxIhWSrnbZz9UiVPzVdb7IEp/VAqjqyvo4egKWv7+
jgGCF2bwb5B/dufmWSONtCc0BGGtrtLPGY5/z0t74IRbdg7h7lASJkXoC78R5HGQ
5pvqfcR3KwXwjTR+yZPp5f8wRwG3MJ8t0fnAjjsHgk3uwsbQU+eaa+93SQQIG1l5
A938a64Zex0azTLAGFMq0pYs0IOCYF/N6KlQkGdAGHT1sUSoUVlTBBy5lkmdnYB9
ivP3pLQxEM66ctKIyhseoFCDwVE3c5OKO1JhmUHExwiknRajAYeC0JXmimQdiJYp
YNJ5ugZh5LjZ8dsESUMazdOZVcll8SnvzjpexgjkHKQvy7fQFq2sdvJF+DIs7sFu
WgzXjDMLe3a2xEcIgKn+Wy7/FZTaGaot4vcCY+aa9uLR2s0+juHGsSvgnwoX0Z/l
yv4GlW6H39phpIZ7zaAxMYgVcrMK3dmuvce9gubgu5/a8a3Hu2ezihGBaFrsR+P5
JL7eYAz2gtir7kla6qYlXefP0noK8nYuM0V9W/RpNuUnd1RkWALymi5WLXcdKEk8
n2Img7xWxyj62oh+8y+4qN9s0tDnneh8RtRgwOykq3g++3eGKRN7OnX6Cr2HuLAL
/L3vGIDAMOx6s7ur+xOfoFxSJj9iUJXFbkDhtEeZYlQQCKUj7FTN3egKGpApmCf6
84SHvqOnjGDZxZ/rBUSKdeaJMRXYTV1ad9TTBM8XK2wMuiZ/UmYunwqCHvbVGA0M
IIYJn/+xJSeef+DXBpi+vW4kCk9e8t80dIdPr0rsX+6WmCBMrO5JXOkmubySmoxB
78OPJgWqEztRphzrQ66PVdyrDx42HiJc8UIw1mhBoYMqJylOUMOPjE8NctwGqFgw
yYCHV+v4YMr4DhJE50Vw9zKN+3tsQcJjZFpCvkGxFhp7AKuEtKCdtJZNCv6lBFEG
4vdzvWtzpMrKX1Ymj8Dl+wGoGD6dY+SsKW3EDdObYXYVFQZ0lMFVn/c7PVF0tMiW
Lj92gO+ms6E7X5qnSw7jY597ZKbRL3+LSBYx3mEjgyWoAkksIvj0JslIgFG8zGYk
6HrigdvVk2ZWmfoMidq7q79BwfINSl69RDZ83OGm7Ev3s5Ue4OmtW/zpTS3sK0qk
DiUbHcQ1P0FvhAKMQ39ZrdZtCXDQaS9Fn4eOawD77ataXZCrP1bCtaoHm3boJGVU
AsEWbJmDn5LzWBYRx66wQlv7HnX2EBZV1DnyRNLYitB9rU9iip7WkTSzZqOXI0Xc
zUDYAFIi+oEujeHFBxA67C4wOQwZezElHpH2Wm22+8MUdZcjWr1E6SplkvUfafNZ
HXQ31aOflxvOd0TynNWylSq0rNOREF+W1sBYVHzAq/i0lnMUJvPF/QcY17aYfwfc
yBuNd/XQe4ILI1voS69Kc0GJNoXXvf1By6icu/bvJyRWWBBfclGfTnyiBx0iT08o
FN8GlccBgCGc9q/TUbXU74XzRtpDFcihO+gqw4I6pX6LL0ETaZHum1qEne9fMXkD
6RGP8idGXkj7SgNAVSEHUbSe1f4M5kUjU9W06fNR6Dem9BbqazpVEGmraSqQIf/4
aZHy3PS01KrzzKa1cnmRkDIP0EGzCaS197Yg3CY8kku8LOmSSFzVNuT6tEP8O5Cw
pXdgLvSsIIT/8OIXLEbH4KsxTg9cwx/ngrUopVU56kIvXietSK8z5QBFgPTcGGxe
8XQX96Fdsw14JrVHehED+AaegtCHHzRY4vqza0yh2m0UYMN03yWoBm61bLqgk7v1
B6EyB3/4104W06gmAOWPBiV+qjbKXvFPKlDrJ1HtSCJHfqqsvxZyeXiLEabXleaj
C0m/LDqjhXIxK9Esp0i5ClyWiifuiAUGLhPK3d30McWk62Ya0eGj3wVMHh/HeK8j
HIEiZEI1duWR+ftpfQQQw1PUujhd2AEPCTGe0UQdZng0erQwq89s4zCwB7k6dsVS
x4xQ9pyZqkJprBOjRHjkfd3PKAf3D4YBe+fGtR+uPP0+7yEhLyBmFv1jBE9xmApW
0vU+3gyLfoOvy3uUjUvCUku4aW5qJoiHhDgBiSe41dDbIbeLp+TaiT091J2v3yPc
aG7/x7KIU6OyBQJRsCOteFuAAe4sJ/QRxcZM0UHagizF2wByT1pzZXk5zHaanUUj
P+xETqs+HM4TRSB3o0YmcnbE/OCTEoJN2D0iaOAC847A97DGwvK0PjLrpu4LVOVL
bJerifEBA2K/bEyJN7h/I/otY42bev+I66PoSlKyyt0mXj1V7+Ef5mKWGAXb2tKe
dkotXjcNqPC0eP8f4Qbw975ngYi2Ky3RhPSGLyE/L3HNJmTQoVp62SyD+WJBejFx
sUMt/mLWy4bpV/8DZmZQfIs3KIrQzBkcAiL3WAdvB994zCePmRzu7wUmGgGAq+92
kQsaYN62j3c5QVQuWkZzyGy0k1ObprtDErbH1bwMhdrU3myMLrJzaGR4/kIY4uVl
hSvAFjUVGPot8RJccsNkQn4YLbgs6/l3Q9TvcZ+NjzWPP2IN9WvGwF65RPzO38LW
teDzMp57M3peq39BcK8ykQRGh5xKdj/zFpnntAugM6ZvpBu/C64B6aBWyll5Wy9E
DzVGI4baohOWkGnsq89Z3hbuGEXrf1tVXl2X7NC3hIzhgoxL9MFVdbsa3OvSdC6W
cf0rNaREKZE4NYoNKmIEGhw9RRPRdIETIMl4kxlnUW+7fjb7/tiUsDUjGh2H8AF4
5v9jSWdIUAqS0putODjciVIYvLwIbybQzU/b7gsmw3G/v1I4FsW0wSnlEkDU9/HB
gJhiaFm5FxoWcxZjbWhKt0ofdjZrFKexFssESAM8H5QhNUrDcCWwuWbDbLC5h9m7
IuNtsk/oEpeZEdXRSUoMcWTpESOSKuO50LYY2IsocelpQk85JukA3DQVSVjLFh0d
yPXLY1l1MmvxXyPdBv6yLKcKHk/PPuxGpvesubaodz7iKLMqjbwvxnDu/gHxaHG+
wQwBbiupSDOfQDYVUSgz9W54azhQXUP4cW96IPR1SOLRuIRMtUWXdYg+iVt+qp52
2/24KGpXsFw/pJKCE+bHsqCOlqAFhB1UQsqKsiV8hpE2/N2EBWYqyJVSqACdXsQF
5rh7odRuCEAtJbtZf2B/M78NSCsIGAeQQoyDUJU2b4HcLK7KroeaQ8gyi8/F8+xT
qP+8EDLrUW83XsP5ibyX7pEgbHkKZl2gn98ayA/GlAMtViqEG/ifYY6vA7mkoKQR
eqQJ/pNjDF0QT/cNzFJmPyvoRgQjmaMq/HowbaKMT3eOVoujZ220x6LBPVjH3Qtr
u4G3RDlRohRVfdxn5hf7SDhlLTkOFbbY6CKb4JiuiymoICUpqsBOl9oSlsjkxl11
NkJDr4YRHXE18uzXYr/w2xiSOXrb8bAoa8tckzAPVLLfs9OjoX7NAV5VDse/H6Zm
yUVG9BmZHlH2wdr13xwkmFH1dS2+uA6oqMLO37T3Tq2KATyWAGsDx9Pdyh6Q5oJ4
h694nMan7j1zq471pP9vREqtpHKOZVuPD9SXHV3J8RToaM6Ux/i8KpA/ZvO7Yx7F
Hb/AgveEJFfoDeOKH9iwfLXY62qUqiXWz8EI0R2WzfoxP4+lS2IAILiNBfNl5A8u
8TT8b/h0Ks49v/+pxph/u2Dr5a3My9gCYtNMKFia6Xs4Y13fuds7HVNV5CNpwMDt
IL5EqZQ91F3KOohL1TCmA+umSIR1R9EbZZz5zaymCsakiVJJodlK2Giiag7NK649
rEiEkj/r4DbYrA9qQ7Otx/ayHhP0yfmGVnBXJoMxjUnrp/MV/aAGR1JthRxJ5DUg
brBHGCOyfL6E1d8lYr+txpw6/mHXCV3BWy6YVT9QPf61ldWuhftOF0t6S4cWS5uM
RggZUzjuHfkpekdiLArTPENYEQCjl+6SlAzvwN+HHpeW2Vc0igkGbpe6iaw2pdTe
2bSlZnJ1pNWkFrH4+mzek19d2NslS5dAG3IjwFjS5WIIpffiPIKyGMkCmzXEMPVU
UrdovJ62nWW3zba2vvr/oqIBt0v3smsPuCHZeIuYGBckZHb8kSPOZ83El01Nn4+4
LMkkygynfADT/WDvX+YWU+JrdCiDygs9LCVSkODwwzSTc7SqjVAbtBzUXd1MLn2D
gurIExdknL3ee26tYtud7CKsV5hpZzCswhk//JJxsDsODXIZZ6th71XbP0KRryZ9
w8m8MgQHee40J0CEhd6Gvz76ou9dFT9gbgm0H0hAkvBZngH8/mzRsbKcGgrf2j7L
MFtsTBgrMoiBfdcXwuhdM7GnNCoHdUGz1dxDFSEpsR+twwSOit8i/T8UqDfh7kYA
GpydSt5zPTfAEDQAcba75E9hAu5o1r7t8Z2lUQdsr35WozDbKTNM8OqnaTkEwp8m
L5hwGqhMwOypGKiXF8gJqCFN8gBgZ6EM6bNPVoU1qk8j5p23tHkUcPU/LchPES8z
88Ee3xo/KB2V8k6JPA4cmrrAdJcm7hrI+NSSqW6Cu+NWqlAmb991ucaJW91oFB88
kBouye5FK95dtqErKZRzxfOzYq/PSsWrAf+oAkG23E/uDHSCHyAFaiYVRjhl0xQe
bLYWA6UHrUYrIb6ySxDZMbcRO0rcerKVjE3tee8DzX9l6eFECQDMJLOarXWaMl3+
Vk295M03P028PTUij/dAZz9275Rt/MRqRMXgcmnI63PQTGBbSgiSvWMaIdeTHUcb
oawMwOLK21Uf5Vohdft1542hXC0/S+zHA1GfUl5AztjUfarN66k5oyqJoc5JscAH
iA6LrjpnbTmmwKEBCGDea885pEZEMV6tIo8XdcYNxC88dkEF3wo2PVAcsqpLzz6m
DpwRnndfEQGbcOktCFNS9mlEJt4PcFRJSmIMbxipKew8j4TP6sMRYm/wjF52Ts7y
J0DnZKgfNAplpqcckWX9Qu/hBDucoVxuV1Z+WyBA7v27lRLE19y1L/n9CUan9lkO
yrcbgSGRi6YuSo1xAPjRwA0ypPdSN+gPxhLysepApUfe02RH9hGWgsDaDotawpfO
vfuzrfyqS0+Ul/DGQVQw+VfjdUFHMy1nIClpuKlnMONvD5+3kyPmCKvWDWtraw6x
yx9UEKE6BDIUA3GBWt/f+6dJgPuxJs+sIom3iULx0prx68aZxObxLkCyEJep06ho
+f34AinjFNvqjq+SYWHbrkPH1B1jjCsKiHQjxTiET6I5bFhsYBuvERoGGKyMUvvI
iXZHo+ZR8fhtqh+i8nKz7NNTBo+4J4NSQBnKyF+3sXCIPJ44Xsdt9pxLlaRNUMQz
9ckIbwscLwgQgx8SELppE43Xhao/8d116d1jXv866HJzit76CDh0FbO/zSaS15LG
ZDUqiCldM6J+iR02CQYQdnBRjRhp1UQqak0ez0/ypxQBk45Z4E7bIHOESxMrc6Ea
W1djnTub1Z4YdgPxZU5fs8ysaKBfZiEGGI3qUCyzQibX9KEeU5hd2Oqf+U5gcJHt
3mo0HWjWpJCmaMqkHJAbQLEBL7bNSLRBAuzhv0F9+FmG/6kFBP/sS+CHFNAhdbkX
u6dcpaiZbwCd2GFGY0TbDvADhkvPLIEp4aMUajwNc6BTpcQvnmcDbcRNK2nLZXHP
gw1YA/fRGtcOoPqKJOxvE0w+P3tD5V9Ceo33Jw0lqxz93Q/h5Bcm5PljI+prdhaD
D2ftwONyJxLsKth4XoPJ2bUITp038bP0sVtJPFRoDyi3rVo+L9JSPQpLViUP93/l
jjuiEloPZwWNYj0g3JlmVyKUdQmTsKnnv04whGoQNKatcvfKkQyxMHuMnb+QoZ0L
4KGRyNp7nA5rWBYZ1PDnw3dMcbclX2hfdL9+MdAtP/LmSyFnSW3Qq7izQTodTekQ
zXJfRQbIBaO1jBLS86l0iJzVBqowiLpQeC9JMHwzSZw7Ybv1b6GpWVLRXWDfqSrX
/vFrAre4XgulU+zk7sl5WrlY2zuBHTilQ3szxKqth4Sk+VLYJWMH8mlb3Ic3+WCc
txEt4Tvge8iTzKynKgvWmvSHSSlaSp0BGTdnQQOySvmkSe15jgV+RF2ffhztcST5
EPdSVFFQ6ET5nNjXbLXcoXgESOjc7TQRe/jtgXRq9PYqL5Cgp+08jLLqroRUq1D1
OJlBddoMD0LD8GEi8LrE+u9yP1iFAEaToYbYGKD2Aesc2yXoX9JaSuH4NIZL8wRL
YykCqpHZl9vm41EY4DKWZba7aRU0o0QlUp6JVbmJtLv56Fxgpuys1t+eecuBmWMM
xozzV7t9dDTmMBvpE1LiA31KMuGO/BVd1Q5FkjPKK1lvNdLIHrYjMMoYHGDlI5Qc
cARL0NeWrFS1OlX4IEIDG19o9f1iVF3DIJ2z+Wej35bsEBp168JEv0OgafMfFj7g
0v4HjtT5rtUhXGbeOPj3lUz+FCn9D4rg29ZV+p1O3eSfJBuMLcK+che2Mhr2cMhn
z/fjIF0B6zpEibhU/1vbR9E2tboLmt43vBVs1hzPwpWzCpxNb4JKNYZ/RN3V9iwH
qQoa0smY3+i8gPgyYX0u1kpilHhMhC4ar98bY9/FzKNTsLYMCBJpFfwb9fbZ9eos
jXWRiTdeEUWIBV2SARg4IXQ6WraqkPvDYkJMY8hZPNPOTVfzUhbWjjlbXJoROOYl
B3My0m1/7pomLjaN8zEYWq+NjXwOjij4vIdyH8s7LgM28SOc4nrQhylmwgbxrZ8f
FENc3j3PVjzH1yW9DPo+mlgmV//nWUMDDIqNefOk5Yc63AnWb7eVIu88XW8aj9Dy
v7lCO0Og9agtzRftYdhcFlFV+Y2pmnO37fZfdmlclEwy8ZLPgopM4LiMLVaNz839
Gt4flarFTO3Ap5Ssy0TB3B4Z91jMsI31jUL/aRnZhfJ0UxHavo99l38syhX6OhNN
8wR4WJnCip89hXhW34Y2wmfEGA8tesbS+4Q0EN6Qv9dqlmB2ea7VmveyVmmV7LMq
RelIoFzaYcTZGvYFJXCEf7a19xuMCR5FlyjxwyDJg8YJBO+fwZeGD2Mkjm6pNRsF
CjI04TTdS9IbB5RnbfmV5PsOy+NRWKlRGkcnZ2m58bNI1VrXFXNK5nLyXDtT68R+
FT1KeCQgZOgN3DP22BN2KGAooxd4t4kfSfqiZPv3A7hTKUVEaHrxZV4aGorB/SsH
jI+pG006Wn2UFbSI7B9MUkc2jrm85n+SUHVymRiF0+KWofQUcEHbjHbZImCqw1Qm
IHMZNGWJh1PjPxtvevJC9TWbtbw67446l9geWPInrabIJg3kOtMpr9NHX2GpCONV
tiwHOXY+yA6kw3+gJxbC/QPOfbYZ2m5eX5dNjFn2G7Mcrm/VAoMj6AEv+61waEWg
MLwj+hHkNDLpGEFlQpWrXNz19H9FDTgGphLARKAjPyuZExEDb7oq4WCsBgvzqd+U
k1mTS/riVBzXMzL6Sjt8/+tWHVSJZ7OB6/IZQMlVKux8XKzRSUzBZ89EK2XqsWiK
2hqp2BrDIZ5jbhdcFINEp6RvlGJVl99UJwOw7GOAQRODELXjPKVo6aZyxaO77uga
t9RKCoMGdHWMBNZPJrlqwJPmBkybZzSSQmY/fzagxhdYxf1pl+RnMh592stdltWw
eNAIUiJZYJ+7D25gDcLmzarm/JUxGL7GXBenCqfffHYbm5PZdYLtIJ38zLVym/D/
gjDa5kAWDkoP/Yeaz94ZAtoCuAyb/0iycpqlwr25keaLfQ+IHmiajKV2zMYrPcIT
JNLTwXE5KyJ+juby1ACuNrcvHWVLvpZ6PD9LNhOPIs4ynHePXfl1A5+D8wT2XImh
TKEmViD0IjR9EYkMawYL8y5e/UZqI15gB/UCQmPKG5/ERb/aYw9wvz9ZC/GJ2AVz
kmKf5CeY0mkQB11LraMjtQLmrcNCfWb7+/QBYh/Nz2ejmj05b5Y3DKvEqe13E1YW
pD42/osLL+Dxu4tFmBEWG3IemYhhEYumhpZH0SzeA39mEs3dUh3OC9dap3ra8pgv
ZBWhZHLVgZHin4j9wiC1xq1vGIdNYns5EE1OBFV3qSMtRVuAAgZJq9Ta0ZMqXfFe
YpIt6tbR3wtnvQILzviCAt5QrvWouYrXw5DPixKSv6L1cf0iBTWE6TTUt3/CLyvO
em3l7UTKs7EOO4jdpiyMgXe5vCkS7WhqEjXmjgcTw9l1Km+TQsJZpL5/+mnxlJ06
EttN4klyRTbhffo+AmcU5yPpoU563AKiSMrxpDiAHGtQyxh529mXTqwj3BCecl9d
pSBzQGubZEv1YynXRRs6b6vGpsWIxUS4uRRJJujVynRvwiLxQDLBNSCpxWeJ8YDn
G3a5Da4igfed4Ou0TUEjT5CWUtaGd3D4DQSbOLXhn4Jtr+cgo0tLbJ5CpyncOV/1
aVouOaGqSPScKAQRvu6HyqJneKXq57b+stdnJ5Rz87Ye/7VhgAOclD3zptmtnE0R
0rl2w/8vzIm6++UXotizNn9AUQmqXvQhRaUECaNRaDVWIuV3oGLNgrWywMH4WeRG
nXcnPDEb6x5uGYIUgV0nQ/8BUpuJq7m1xgy0rEbtbhgkui8OvtaLRaBoOuk5edTt
2vQRvhEE0UrSm2z70cKGWcF6o4vl1TJIlLk4TmeDKsGrV0isoPUvtyFx/mW9jIMB
P0J36lzpQTAtuoplW2WbmkiaDS01GKG3eY4Q3HIVo/1SbrVnHbaujwyiqfzcyK3n
Iu0ndILqjAW6cIbRHOEMa5WmKAsL43q54S4YoqNGbV3weFppHo8mnYbGl+g0LH6O
tOjw/iLPFZlmmZhWf5CWQX2COMFKLnInQvvREWJADEESuGcs1xLjyuKuVQTn4fcB
ZjMzNPSBEZmWNg3cGoTYdQIli/apu/5jeelhLzWqWJ7RTl0uaLxgk9m/uWAgh+Ly
CYXalMIyEKSntJcMQ7Gv6dqfwb2q2C6iXTVL3jLZTRWn4SnvmobcG908cgwXEcu9
tEBVKKjs1TsDtmD99ghCgVk5EOebjr1QJhXdWURJA4PjOvPtnjt4AsbtS+nMXI4w
+3Col5KO00h/MIQqEmp+KHlT4t/aOecCWD8d+K0/Z902W8NdUgYiRlP8EJ43iKbw
CMClqmlFLwwverAgA25zX/MoEtOqnk5of2i9biNMviX63vQouMkBpu7FFQR3ajuM
cRe4x+L+D2G8MbTs2WTtGto/tr05NG3hGc+SZm4VNKn7GnNs14OHp/h3ThUerB4s
TrUXXViEd2CoiGO1015XPmDkGtUfCiNvCy0MbX9dO7S+nOu95rlMIeZn2kZkLCO5
C7nFnvN40Om1MkM2IaAJkZlxp2jR2/cszESAunASdgIQOKNx0cjWDWuqg32AvH/0
R54Fosp9MAJAbkmTxRRABez39RJAT33Ap9bFYKjkNnt8r4PIoDHDNt6vA0gkFQYb
4P7mNku7A6IR6MZAWq5fdVGnuaqiG+W5n1TkHGhPkkbaXhuJzm0RCQKXOoX7uVCc
14+yJRPe1TCwq/9SS7XtLBAdQELoW5WSSpSP2muTGANUWjdTX9xJiXIrDy3YqkKB
F890mxufGaZ/icQrdOjGzhZRDB+RwEp71jrw9FrQSMUlA+Sh4c9d2EWM8sn5Q1Z3
IRAjHqkMc6YHvt9Nn61ROJh5xZEDUCGSt8qqcSPBLKwZYs4jT/7cOzL3yCmvvrsh
PB0YKRlhTVl3vDERLYn8FZrSKLCyKRPxKDsn8tW+3n9cgKmzWSe1zVgeGBNsZTOD
qrzJBBJDWI9iXqSoAntfsvHVU3aiq787UM9YCudT1pUcf/bFdAHL1u9GSWJlZsNJ
hxIimmNBI4a6A764m6fk2KL16HHGZHFBxysjM6hUJdlg+VtAuOPkG628WkoQUs/G
CAq9Wp/d+coY6wZT+0DVTok/urt4hJv9k0NGLU9yYZoD/6NAaJKTHddRHNMySMD5
Kx5yBhCIWEEDPeximX1t3wjy0/7PmtaAQHfkTqD9UtpS1I3Qlr7YYw9opgBu3oFH
L/4SPSYGvKBACogVfHkMzj1kB/4dm7K9Vbv04hhy5WzGW62Ctf9Ht7WcDuKLt3L8
/JcnJl7k7VbV2AcXMj9+StSLjjpdRqEZapMVTGI7gwiBAE1pW336adJ0NrcH5wtx
fKAzeZ4aZIuSYffOPA+hu55hKy5Dum3BkeqAZhWw7TPYnZLbZ1S4JjEVsu/SGrXF
lRUXApR79HsZH+hARtxv3mdtNXwdOJZO7oQqzlhQjcHBo/3wHE9SS6ExXJxNuxR6
yTjIWjeEtP1zK9DjXjKICBXr1rOogBlfFHAn3wBJpxjBy9xtEzOjTmrpntfqKAst
r9CUOROkXScBtmujOlQVEDCaZ0DQ11NDrn3FoPylwpZnCkzf4xovfekmff7IuzhC
AO60FMaqrVCOCplAQLjrVhxeaDveMpm9aiD6xiqaBABrYpFGTHXVQuz0qAfbl94t
NZ6u0GflmDNpc8oXhCIWtIIUXwBbDQ14HhW/bGNwJROooo4agPR10Ew2TO/GdYFA
NxFZJVIxlg81JrJepVF94+QWlYpn9B60oLRM1UPpyTiBJ5bh4B7VUIwzi6Y//fRn
tfltSv5mtfQd72Klh8FgouoVQmM3mYiK5uTUwlLi+AkncQ42WeHdgQOF/W1+EIX7
ib867n7CXPeiWFyhZRfD4mTLUrcFN8Z7paPINoFLG4mEJ7ldS8o+v+ubodkp1AQw
+gdfulBWkhCBUCwDRPzuSyJi5yrOPpuWK3px43USgqjhsfLd+jYAIPIe0ZqN14Ja
Ai6REyCrq4MbKDnokuvGafswG3a8p7i4oSxmGcJcJSnVAEg0vq9D9ch75IWGkipu
B2bZt65gcjJaYYctLwjwqkolJw9pXoiAAfpCacB63JcBViNS1jQ1bxuWXdYpvqY7
o0MtCX3VlQTiC8hMQ89za1JD1YaR3Vkp0w++HnywsT+emcqpLVmzhMxU9iF5XcBk
WjkhA6psiS7x3TIDCKAH8vSIWt2NE6HzglDqY6xOxRb9dUL1NfPGMYJsdupYQl2D
NmD6DAaZgom6gp5dvrC1fFFOY3A/cE28fb6WH55+F5+4b9p8r3Fn5VFJlSmNfTS5
m06lZTL0TlVE6LCqJXaFTbnk5JMB+NQYTxYhrZoSmZxjeqouK8gW6Ci1Eml74Xs0
Yue8nNQ49g0158/k4rxrASlpcQzUucfBn47DhBmY3y1xox+QkDB13prnQtIo44WI
ytpmNfO/C7tnz63wujsLjPSU+r0fHgX+4B/FgnZviAx92TntEceKRjHFbHHrfxMd
ZPPP295E+dMQXcnuZwCBVfECTVdMPLN4RrjxvRr0JxWYb3C31lD2+qyejGGMdrTE
l6l3JWr7sX4Q9zrQB3hwgvOEwhgFajbO0jerF9ZVzsgUF0dwAF3Ud184rbjb5CKT
FpbuRD77SjEyXDR2zf7xNYSoyvSTQww7D5WvGRlCQxxPCsskOA/b8ikGRj13gwBq
Eh+7g6XDICagxdIi2nfNphTh6ehyFYjNONTCW6gqAY0YT8awTOOX0FOCk1S308dx
K1Ky2rlVIDX1iUnlDOjc7fDzh6KQzK2qX5GINVIwYmEcXc6jKobHT3UL7Z83YkvV
T+T8WMb+7091R4hwU0GjNkEL5qD+ooPhV5oDRYEuwZApBTOjT4e9yjBH0eN/29lR
k+W2soRqjOedNCgC/Vf95hJOfp+VcmhGNR3lCJ8Ky4F7QvzBhQv6QFOp7A9bOoX1
GsNIx6oPsKNjSlS69vx0LdOI8QkGJAp45kWuiPSepm/lvHVvunKBE8MxmAczhL7b
l2NuQqyMDFOFgQtSW54naymAyy/artc56s+9k7dOxVNcpT/StDtaxYfJmwLECVPv
LchcLbr7zpNPMKGl9MLEqWFwBsljx9LhklCGuEmvVQCHjzgHf2byUIZXPag21W0L
xchXLGJc9SpeJ8lOZG3HpOFWXogEXwKq9Rrf2Ovqt/zBF3ng1giOxb33enJgqFYo
7E1xYKW0iFSfxqVvJfzu5Dj7ugP2/sQTtXCirIYG+6JKiMBPV/7Ha3o1Tr+LQ4aT
qfmJB7Qj4B6xwrDJlEjesSROKoNO2gHKQoeVCyjpamdNepABYKT92GZBms17OZbt
M6SRxVxC0a7HtgurjqKzJsRUpgsm465TuxjSYr1UH8cAqCNmbN/1Yq2NmRoufvWw
nNbMG14lPQ4bE2SfOp9huqtAIcifMYWMC0C47QshnDOhGskG/KbQ2QEiU+czfsBL
gUrQySGIXnmPDaZax4mBiDIsOor5l9xMDJDL2g/HsjNNngOQtDy8Vt8OvFYMwRJR
TaNGCmX25D2DtwU6cOZvKOmw6wf0i2tuuK6U24O099YKeXN3yko9gyccR+u+6LeT
xtt91bsHCSdzbTWVwoyQVki/geaFdqWu70QZ5E3OIqo+XxE3WeFnuCOCf+lfoXIu
lQKXBn3qqx2kS31wD8OaotZVet5/jkFvCZnqq7RD2aOHqzBEfRsZt7CLhfxHG13S
xCKOxLpZJGoarrinUTGV379HpzzBYTsFTTdTHtdwdknqQFuiQOKWck7rZjM01upx
hLMqt9guOTKD+nwptvm1H8nrk9vQeiF+Pv3xzq47ilqyMTN17gwdRUxXPYcm0t/4
b16uv6Sd2V2pzJqtWKAXVm0Osj3ZH6rFc9KwmW0UNgX+PxVuswRMhl9dySECIxfK
IGEIsdPrQol4ob2CQXtMK6V2+Jh23gSd1fAFgCpi5TabfimoxcL7U3Cq9UFdzPJI
U8wyz8kpb/5lAqvZY5xRhwq1TzsdIwAyG5Vzu6ibetN0ongm6pIHXtZOcw8w2PDj
IMBbxx1+nPZGT+oW/+cH0TO5ywtiox/EeX/bvwbzBVcQNKJERWaym2oJpuYozYlm
+7BjYba0eh/ycY4n6acA4Ll9w/h2SVxLe9/1samUzxsv+KT49U0JA6I41f0fA2V6
PUmyjAIireLjg9rW4RH43SSBrluX+dRJWxXHQP3A+m9IMQJgpK3L6waPYkqjqqTR
/ERJaw1GEYBz4hI743k2tAaedlJ9AX1ehMKyWFxQ2xW8FaenDchtvhR9QAU9GugK
DA7Mvi8vUJEkD4Lwh7FWxURTgwmO87w+5Lxj/wA5P1+DU2XdZXNkjUexfBGipRgt
QLTD2cNjYtEzPl+adnzIePClInZIuqC/1zXNxgR5pDNk1XADI0AN2k0gZZGcUkjF
XKYvU3p2GpaVzmhcXxLope1WYe0js1s8gjlkHkdjQU++200WLU9Pq2J7TIthRddc
8ffU5oAuVDtDXQaCnjWw6zVveJ2H/Zz7a7lSErd8/fK5pT9jLNZZpOcCiiJjaTLR
WTIiXWOBiTvArdJGf/G9+9nNakWAv+qYck8UQUSvgG9AHwifnFLg94WkecfSYdOC
O1bgnO93lhPRuaRAFCM7OZR0KHPImsLjiKK/uc7SQ+Cyq5h6J9XeizQr1ZqJyzN3
aOP6d9lc1K+8ju/f3wDwKDRD6R/lstO8qV8jPf2b8NcURj/6MgBOQyZtkdFY4F4z
RZMRsWlPzXoHux888mwQlQu1fYbp4MOnJHQuxL3CSPYHyb8uJsnA+AnE1IFms400
GbaVyJgABTBL3gkcXc3k7B92Oc0HIZJiXrMYoGp23NkhBOo1epi+mv/xDpwzMPPk
xb3+1Sx2aoWcVW4kf8MWzdiXggJiQfMjadcVzmPkTexS3n1IvkrifWdhhceE7wUk
wnhOsTpCSZuWgPixg5QuKFzV5K9qzD8lPoJflvYtnvywbVrIEeGQQMHXypRXk4XI
5r8Uylo7vXU6JsCtZGSaOWJjTx/qrNWIgm4C8B+s8CZb8zZbrKVR1ICyWG0o1xS8
cmj3LADJTJXpZeS2nis65VgMEXco0g8k+s1+mHNadwd4/FY/nAaxSGhlguSewL2J
nZrPXSbNrLEhn1hvCR17R+HqQlbNOt3hMh0AmbXA/TgDuUdz/d49b0o4ZLI9dLBq
6svaVY/AP0Lb7BNqDkjpSbaQIJf87mYZliue1m0kgED2nTAXMngaai+DyIFnF/bS
QxIPFvjyrUf6Bmw8ikOp0BhEPcWWCUkNVJAde8SprUWg/XlpFWMQF5xxOkOB6FjR
bTL5/HHp+df7yIDm/oKFnx+nGK5KMpcO2psZppxmiVT0I+sGhcciOuM9DJ98a+1R
hJdBTGL6S1AbrM9OyiQ13s6dQ9t5Xrrt09DglWVy+IhPNMxqn3WykGTy3hIYD5fY
R2ppGvk3cgjwfO4ek/XnGFloe72GcyFH/gktSj+CwBsKFTBWEvbntFST1yD2lM6J
iyIrc8KD3VttBrYd86X+Wa05wI89aWCNR9hLtxY1u07LWsxMBd1TTq1fnWm3k1ng
FSGJ/FWv3EqXJnGoPOJp+8gFFV6WCrlnv1PmwxaLgSyhCcTos8TBcErju+5XMm4Y
dpuvxNbsKkJjJCKwg0vnnoy7rRqK5EfFwwBNnM1iBO9YAZc81b3PoGOFgjERhlQ9
HxRAmeac2MXnpBNnLpeDnG1yaHQcke9kk/yt5JHtwlFkBH1GXztVXa+kQra2Im6G
4az9CqjuTuNcc0FerT0TvDEb8xioONrHWmHBRgqw3+sq8qAvE2OJc+ZE8U3kNw7V
5glRBguGirI5yeTtOll/evEIkhzIW+Kh2LRrLciNAVq2qed8pGkB6e/g5YQQZh4x
C/oyLE3VQAW3d+6kOpOOOqXx1bCKeiWRbpRrXM7Rea9cLQT2AEKIsjfxwgZZaAfS
K3H9jRJiAJ//MBJRrXZxNYf43nyK/qlB0Y7BhgVVC4tosEbzbnud9r0i4/YO14uG
Q/yuQb6ZCpzGgF5QsnUN3wp3rsGMae7TcIGdupIPOrki+dE/8+AtWIcM8lwHXdUS
qRpzILwVa8zAYT6NLrYUIAy1yFfthEpag0qKUxq0pmV4UOhLebGUOEKaHxjIqMII
yt7H3FplYt9eNZP9fzwQSq3T5bSL9OMi9UvQ6OyZTMmaW2BfECvCgoksxWq/IYke
Md7EejBQzY9pqyfRIlvYkx6b/TXzyeNMzTcDTZC9jO1ImmOcXanbmUIkUqXPOfJT
rGwWG7JXiL92+RQZte6Vxe6FYnaXNJ6xCT70hyAHMj9KecABichxRjJoDtV0lbYo
h4qkrfhbuuPHIwjg2euUNUit5s4j6jkozml37Pcb30TLdyxnLYGK24rXEcL44spR
gSdaCdyrDeOiW2lj0cO7Gq4xcn0oyG4RAD+yWNI1tYdpwq7RZCnJ3A/gRsSGcTGE
G1/9KacFoxBr77+rBpmrcEruk9FLKQJhB9rkaAgl+o8kXfFcjL5vTvwYMYecnoJW
ecN/VNHtjqGURYulYTtBYasp6ptXLxyFx8NPfSYW39OAINM0PpVK3guagVWl3Otj
o8p8An+OJvtYUUazebWxkSvwxp4kpl9SaJIoJjzacyhBRw9YiK75fkr4aBCkFuzt
NiZTfG+zS3rMLPghyl9Dwrfk5RM6jRi5zFR8SMcIE8F5iz+nF0UzXPpflIsQizBq
R5nSRjgJnzeS77x+t1asGuZRT62fjuExcPrVjJ1QqZm0pOuPmdVGO5D+sq9gyELK
Qbw/h0R1jACtcuWn08o2fDnCF6DF2nGCH4tog+hvXsJPCa4+ljqUdi9zLLxGnW2I
Dox9taDjJU1jIF9IYlwM3Ilb7Zw3/qrQWjkUWBa5KY60Wwv6E2O/E75P7rAtYptC
ohST5K0qSNN6tMA6HvJfpBayvk7p8eQNPJaDRzrpIaFHbyFTJvP/vcQr5fRuY6z+
X/aVCiu38e/kcTckjMgnKk5errMo4WNVrIflA4C8855rCgzpBZ5j6h4vAOP+G8s6
d8f6yTh+OIM99KdzSLGNYK5tR+mpm+nJdCmkuXhcay0zY8uNVRGJjTEyZfm6Cyfu
tPH7r9OprQ0wGPTbDsDGbGV4xM2AMHJk9MDN8T1rboRb63aqT5VBSW07avspmf4A
pfcqqzDIkhj1N0Kq4ies4cz0asROuxPJVDS4QCVglr84MLmiYJWkxpxViniYOf+f
eIFn2UkzMeXAa9QQ01bAqD8LhD3y/mm+KnGPZEuJqvsoafuF29pgYmKErh2554e3
N7xU8TSiPTqgdWuGPxye9b4hYQffV4AGRBd4lIFjHWw0qRNAaq+Dc6FN/RgIOy5w
gk9Ua6TUeH2QQWA2DHSEDxe9pk1MKSEfBgYt4YisMgGoVkVdfA9LkmgsP3Xdvf5G
jiJSQGAnoX2K+9yWIYEWysI2sE7VLb2aOW9XoySqSCBAO4wzO/mFS+LWjRYQEX7w
/A3O2AcNZAaPtBqW2By5DJ+S+yBI0d2ByER611bLhA9hMxRzpk5oWjZfK0dLx2LB
5/SAnJPqy+SMM1jGtYvo7SwV1LNLaH+HTd6ez/HXrWTRxAJpgoXHEknWxJ5jsyJU
hBqz95ccjy97Sywns8N5z11Sf5TAkzyiai33VVPOdC8qQGWC5/ji2TZL5oQH+KCo
iAjZ4p9QOa/tp4I71UksvwRC8NqVCZ6EnSdw4CyCRK88WpCVVkpp3uf3lsNe2t0c
eQYgPWcy7QIYfdNHgXkqZYW5sKtwtc74F3p7+SK6UQVxcwavBphTvkqUeS9OTaG8
T6kJLguTAATBlU30+3PwO+sXffJaxb+R1rEPmOw6F+AjJF1YxU0yDismSKOgX6d+
6tHK9nhImKzK4yM17vxbqnF5cdUOJgJc01SZ41zdpMPGJ3AKA5L/AspOc6A8dLMB
VD1qij1Ek6mMzydTyZki33pHRWUUWTffsT8Mffz6nfJEbeheeoHRIkn0cIPMAI7K
kDZNG/HViWnm/7g11fOUyC56qop9WWwIfGdpRj6RoNrEE1UMxvS9QQqIuQsxepcu
jKJA19A2GiU31CpEcFymjxlD1j6gQr9B06ACkph5bCcWcuQ5yC/6zUI32g4GMj4C
5GCOi9xt1Fn5/x7HhCUjuqeJ5i3jJ8TzLbXhwHyfef0yZDRd4gemQndr+dhtxs4e
KwSLwiKU5g2pT/gPgrE+vKDOw2VzSgLNrz7s5fDI09OUoYuQ0AQiIIw7N2z3BNoJ
BINT1QcRZfJh1je+tlp8/F6Q9SJHhZx3witNeWAY3x58De3p9cb/8D7zWtst5vU9
A2e7z8XKGFzbJLIZ9+PoXuOM3GGNwAXcbtcq2hbkscPc8kC2A8kDaweCURzVDsGp
LpZdhZ7Fgfcy31LSO2vitD/s3f0WGOd8rClOCcq9Xe3XAzyMIVICI5l8SLoDleru
w5CsG5/3pBlqg3//MN745r7BDUQ0iUDhRW9CoIxqaMvralaIz6Rpc8DrV26JeygX
2sM3YVxJuqyCejgAsBQZNNhk6h79Vpevty6AS9EWJl423zVN5YK+cxaS3J3+yft3
2rsNlspM+LfvsypFY4vCu7Sr/yLubUxyPb+JerJNBjo5ZIRH7PMHbr9bM8tLqOpN
SItFgwnMiQApX+WeNpxDJIbgqMU8u8Cd+4XdBUE+xFrf/Tt5V3Nn15/SQdLAii/V
t/FwRnR5tZSywcMKCtwBuspxatHqvn3fd9uugg0hsu9TG35vkajSMpoVSvzrVTUo
rp4B1pgE1F/L+x3ZxC7z5LTj6CtVCkbwhIwthZPrOagn4LaDVIgjjTNxiB69poEE
WJ0aBslwzAe+aWgAYiwY9HtRiCQx7hucy6/rzTpX97LGOwjotJajOndECZb3XEFS
u1VBZo7FRkoliAW4/woEynstrZZqroOdngOt6uzhbtwFCHWpxIUg6kmS1R9HyRrr
iIeSJuwK1sdc1mjAY0uytaTif/boR4vli7uVtFW+rLJOx9bCqTaOgWOtm7JuySJ1
wzJRu2BkNYyL04d6WW2dmkcOuuvHfdpl5rNfaL4j5xnPUqgqY3Rtj15l7vy/REFz
OHfzf10Vcu4AYWn6rR4eNm0IPE2iIqOQv3cMB1J0G2ZvM9tQKv66YOSrcChGQALl
BrzwsJ21oHzElg6sNdI8DI01DpYz9yvzdoKShOha+NFpHvNujPPRw2A0O7xhsHmt
/+nA80WyKUuwed+CUcXH+tHWL4D4LNl+pga36hnX2BZg8Gd3XuLJTq3/RHbVQKrA
w5P2kozQ3Jleqga+zT28z6Ks3xTaqFFYTBmZBL1axD41fv/2f4jwT1IAlAZ5HOJ4
v6MHOWMqLgDi4hYlSVBOnYZhl6rxuFsga4OLGNiM9XOXt6Bozc2Y5JO3v2o22SBy
LDJ6tb+6ooPmgy43YOrJLoZpojhQoGQM0Nst3/uj/mCpKX37NM8k2DcLq9BLL+kn
XWoeMdXLRIvzNirghobm0e3+Et51Rh8TfzGWFajmnXrdXrviJb1F/Twu+kYQT2SC
KA1FNDjfEc+ZpeGjIpuHATq5pwK/pkOTF1V4R3OEJ9U0EcWW/3d4OarT6qfG4mQw
ynzN53DCQIt7O070sNpUYDjXUuRwCQFaLsPSzq/Z8iBBOCfAuHfrYMD9SiJzIWbw
6KhZt1FYeJ2CougK/L9a+Q1Er8gCc+eY/pF/UjX3vG0GVEKHMNIjoncLBSnLBI40
/chnXJmQtEztW0xXO8SzTy5nHExhw+VjsDBV2ImN2RCIfwH5ZW5hHIiuJPQthD8P
r+4v2rPDcaw2K1/UOYxtr8AM0JiI3CXmLmiVSs6R5z3wTB0tWOAcXlJMuMmWt27r
AttoR8B1qyx17TQIMja+2QFQvK9lm1m4EZ+CDiinz7tw/t38CeUn0gfTwIs7r5aY
gkpKZVT1l/Zbkeg09I5Y2AX/UKcq7t2d65uZX/DPQu9EQOknykCkJjv8IKonrU2d
sDIaVLiLS9SLDQJAUS079VdYJLJ70zMdQCbhWXDNiwz9o2UKfsgw/J9FqEIJWtpI
ih9GMrwlTp9OQ7/oqOpkIYmv79V5f7j1+pR/t0IvYaQSWYCE+X/9tWoaNN2+wXml
0fAwVd6VvHQD066JMShntnZi55auYFkwGQ+3dMZOXikRG8wZ1CnbSkiXe2yhGHwq
EbdXMJELkXg/MVzh1pqS0qSzTrIhPPWvk3s9I4GSv0bedEy6ZEpKDxas+0Qq9rXf
RlrW7hOOda/DrgAxBprnRj2jhT7LCYz3d+DmgKQKW/qxqq7x4g/gFOaGJ6klBNCh
iS9cZ6iw7STYmykpmK/9pppRcfQWFaoZAtbbnRaBaWqk/beRI/F4v/Y02uJ2e6Kw
59gUOD5PB2nLnjkKyREbLSyfDM87z9fhfqjfaUC5lvIaV/GsjLbuxiZ04h0OOtqJ
ouFsW+39+leWGKmzoeYDglFils56VmjvhGyvrd4ZaGr7iz5/7HZWu3HlLoErzxpz
koqukhnIwRl02c/Y5dNXvEP5O+V9xyPGJ+KhkfP5rd+WyuC7wJASIIBjuCHER2KP
BJD0/lURKmNHvAoHZNjURKVP7sz4q5nMRTzE8wFpZZXR7APF4mPzalLZq3WUgQds
lEEEv5MLa3bjRSwBaF9MijSIrYMPuUhKF1XuHzjL6ICJzD2gZDWpmbI6RIbDdUN/
LhDielXMwOFPH6+VM0BZl/CNjCMutWgm11+JpMX6TLPNhie0yGiFJ/sTlhTDK8Uk
ec6X+UFp00uMctefbNgEw748APQaZ1Mw1YT68+cnbjR3/jvcFC8vjgw056Bwk0U0
99+8RMKHRBdXLCbYgMzHIeo2A8KPeS9DwcbHCzCLkSSFGG0oAJkIodrx88vnfKbN
31tHREIuVYOwqfmSJsZ//GPsniwXuG+fQ93zNj7tYiVGArfnYY/8w2B7tMNoT2li
CvgcuJ8j3zdgntSXrOZGaPJa1Jmhv1tfH/bvGnfsJwVaCqcyR7difalHu95LA+Zg
eTH91o9IkpZkenVkW33LrCvwvMnsT2Cia5eZc00aShTViCrZHLIKCfCbMdWBH8cZ
SEuQlKaCWCmC8Xox7AsFs7WwTxPu3uHhozGn6TX6WgirI1bKlOMQfYjiWuKMnFkX
uEuYHj/qXUsUKGpo27KG++Nt5ra22Bs4NGd8rK8FIoCPj3Lfd5l5Vfa9uSTmCQ/i
ANJJt+9nWR31ERqi87fiXH0NUY3XVPE1OVzdZyp6X1rj3UyYLfQ6IpGjcPmcBl0U
Eiud77rwMzccmcK+ffiZNDUUXVRgUcdRElj3THdkCg50mrfNqXy3MOenQNU6LWi2
tHQeks4rnotdzlSx+jgyltqmfP/RVB27KgC1Y2CEupHmFC5a8VDmCyXwhLeWZGwk
sXbfLRpZCNe+GkEsmRC9JRGT9WcAtpxxTalWYfKubcx8Qrn5GkWYwWGtCkmAbFmp
7t1nne+YzSVXXL8dzVBwUh0PeLrLHqkPWFiXX2MFg5FOiqfxxy8+I99jQ8OkzAKe
AJuDbsTc4tTvjFfj0WBD6hhFoiOSQ3hHWtjal0HvQrrfItps94GJCpiI1aeivFMi
RiRdMSOAQSgmqJCuFxYlMV7GDBsZ0Yj019ZjdUN+WwY1Joxr1YJ8TReaI/JOo+9w
aUPrGiup8CQ6e3jb8XTs/4e7hDSYYo7OJu0VsECWETtT+lE0Pr8p2ts+r+alNbIs
/nwARvlJFjc/X4PexakrBzvnv6ONModLaRepzLsQdBr36iQtYmmNpZwSHhPGzB4y
f2YZ51APamaLr1vDKRB09CJbUvWu7DVb8nzsRLytzT7s7tf+zqUqlL815qNFAEx5
Us8/IL71gWMve/JvciDHjXk15BlbuTSIipV3BpUdsQGRZ4vTDFum5dD20oVohNHR
3TUa09EGIFPgbh3fxpW2ucI+gwAmTA21EI5nyLonHR8/UpnsB4IcsroyHdgdlyBp
c+s4pW3aKmzcdDzVq5vCHrGlk9ifTClNlKCvWET7a71rVy9F5UMlm4hVPqUPOEu1
nce0/8qxvAyfRVbYH3VuuU2pX+abO6Mzp7uAdYEzumjrBvxDYQI8zkKRuQIJb9Kn
zLrL1aThLgJtTVPraDl52ZnWnXzmE5vW40Kg2/uS1qLE+JrRmwp28aIpJ7kUSOs1
PpgKSHAHxwT0VweV60ze+bvz5/rTb6fuQByTo9FxUAbWXSMKmY0gYi4BQMfwyghJ
HT5PEKZD8TBOKMx5TVuL7dGZCeFQUuB9GwxEm5HKaZiJea1BOkJVM6M+cp3hS2Kt
vB665YW2TqY/BIwUVZYYzWSl5kyk8KSMEJcz7l8Msa5ogTmLm7XJeedGT/KW1kYf
HK174A23O24v68yCI5tuvBdq1/tujFdsB1mgFimNsTL5kSMhoau0aGm9FmgOpQTk
1N9WmRa0DrCTGB0v7vEubIcCrw/hMsBpfeXoexnIhAhq5KzesNOZPli2D98BrlW9
6sPmiLgZ7jKz8Uvv25WTyzs44FpfmxuIEeofHhUbBKrFy99nthN/c91doFswpJQl
7W9DTGw3QOVGUhYK3z56fS2PNGF/hoBGVOGBSNKGqb2RwTFoh2P2Yqx3FWWhJ36O
jXmAfCcwKdy+QZmfxK/VWZUahxO5T77FY8Hse9nmocNuYLVyom8d2Bpd7j3iWPdh
1rZFbQ/Y00P1QBYSY5KhQomAobQ1rg2oyEVL81j+oCF1kqYayJDzQ+EnTITa/p66
ij5eSN3z6d/pv2aucn398ltsdwlNyzqsPVxROoZum1MJaJFVm+WV9hvJn0eOyPfA
SP4ScLFvdw73jfWTKF8KADFi79PJAiomThKI62gVCpCDcBxAahR+Rdjot7eU14/y
9pBb+x0UQWtHXq8CMfKvZ/pTUW6PeJ+Vi4dP03gBlYszYMPF9xfTYTW2+tuV3JdK
79cAD7/ZNnFtPo99RLnIe88m/K3+oDhGU+H+2Nbf7pY2NtMDmjEIXCWSJ4bgzol/
TRfseyYIlTtyyTu+1YboHxS/TI1McDTXiTv/AgDSzKVaclMLyrsw9LHOdR9Ezu8H
Re+dYOIQKRS085q1XMo+KhiKKTaxNL3sdUtwHlzb62Lczm4zsRNrJqIyHJHkn9hm
gOcHI0oFvuPEXgfnWpukCxf2fE+ASVr8TI5jHYRbBHeNSYq/p7ZbYen+ylGFlwR+
a6FLNGiAce7wjzE4b14SJ4EmGhpcKQVXt7rmArbVdpe6I+ygB0cTpJiSDqWh2A28
nKTurR4OIsU1Pe5r3szILqWN4qajPTwfKoU+kBkgJ+GKWJLh0/geGX6vgIIJmaHF
/fvC9QPiNgwVZU6B9563bJ9XzRnCQBoqnATb1DbQ4vi21Yi5H90zcEaZd5JHkAa4
HQcVHOQkZx9himF81Tp/ZgTrRcnN6c9pM6A9fNIN7/j7semFNc1g5ztBvBVjigz3
ntXoqL5r5YrvWnIcnY65KLimmRwbCrm3ChDLFCl0g6tQUDvZKN6b2WaS4T2yGbKA
yY5TCS4LGmnrspkqgo+poAiZJfe9GAl6O/T42yoEUfavMM3ocPKxpYZWWwUo25uL
kDiJ1qtNxjFzhSUJSa7dV3G8p5Lxf7QlOgsPZ9fi/8DU1rbRZbYSCLlG1EfUQ3G7
PdaVuYw3QS3Oh+KFLP3YZTM3UA7edcFtKYDYxpmOAjdqn0smc0LuB0EnCICvrHx0
m1qyGWtWOUHRhfPvxwcAVXJ5YBew1x5rRDUDAyc7LC6BmO7OEBYxvVEIucAjJloF
aZAyY/zMoV5GpyzWc4lHZeKhMImLZ+3vaz6jQSpLcx1ll6xSmDuLt613k9UMMP9P
py3J37mgWzEKV1KnvDER91K8RmLPC/rEXGo51bJafuOWe9qZjf8JwG8t7xhWZOKF
TZrCZYteMWhT+0YYfsMI2TYItkMqxi+DTicnIqq5w+oS3tn+LHU4XwQawSvt0YSE
CqBZbYy2lF2v80w125a5F9YldCX/I1oy1YV/MbX9F44ARbwJaOX3g9u1q6aXldza
7+6DNcfQzVZrEr17/hQg1/KNXCFXOob3DEwNfVza9x0w3MqGe3GdLkk12I0Um3jb
Gy0qkNXfNFf/7tNUnt0DGJvdIv6efHQBOkUqn8rGkkW8J7Y0zyqP1EMlBd11Wgbu
v54z05zRnJGs8KNsUeQnBGGKGOA5VFmKUysONRZSPh41miLdGA1O82bQMMhhoQ45
k2TmUPWZXp37T8xF2tQ2CAnEFbQnRD7zdHWnfLJWWKCExbTKvy4as3sdpwW+zEj4
JyKY17qMo3jwvla+pxMW9/nsEPr7CjqND4wCA7Qls5Ta0s1VG1nh3lew7ZHn0hGA
Wa95bUa9zRYRHAfAEaUsS2/+VI03ZwQZRMC6k4WrS41/jTWsOEwYoKVRRYUtEuzW
Wua59PJidOvfkUd+Ru90/zPgSRixso5cdOD73pWcK8TbE9yMeovpmr0T6jPdJOgI
GSBeDYcJkFPSoLn7qZEq8qcKDUl/xtiz8UB6lOVGQd/+ANiBTuydturSSGz/qj95
lMIbGZKen4jz0osrLL6tlf+HLNYx0/fDW1sHSNuebRGGSuGTQxioyeAfdb43feZ5
rK4bG29G8thwPj7Z5VB+o2KsLfXihBHBshYX/niEamUHnviMxxNOb4S9L2rrcq4a
F4Rm0Dxv0sVschGe38LgMJ2twPiF3Fw3772QpeAGwFK717VmWk5rxUIKXwbokd8Z
1Jc2+QHCGBS76HU3usCa84+g1l34T8VqkUXScJJApT24QSGBYyQruDx7wKh/CPGy
nC6zBLUz6EhzgwjuPqYJlZcqe4d8j4KdzCvn9f5x3WidEBU/oIMRpx/Koixhzlv6
eFKv2kNbGGvbjxt3Xntumzxms/ftewhREqFya4VeIPT/hHjflFbzUAkPON8eDNpM
oT0QfXvmEHEmfpdtTIrmxUPG1YMc6OuAZp6ng+X4nGWDznI+LSKv5lRqLlTKZjRw
TmKaLkmWPyAlBAyBeJ2/Pk3zys3LZS5uLIJSeB8GpAMJcYzoRdNmLsOMA31Fc0Sw
a1cGPjTbqacUMLRKr3xi8KgX6FpbtGfCUgfkKN9Ufggr4IlpDFkrcUR/XA0jNj+Z
hLw2vaa0CdU3By1zkB6KM7P8Y4TgW23yMmxNs9eiJuBg2YQoLmnwfOGZ3wImwOtX
kWsHQMDhvTwOxXuPiMrHHXNxrFUUjv5wiy1fJN44LIbu9Qg3PJnWimSreg4E5ccR
7kAwhkfTHVa/ilBk99iwkfcNAAghvzqIG6MRNVheN0VOqhn7W6tes3UegqsPyjit
Ln2jBnUxGd4ecmm48TKbVst90hmnRmE07eQgtrQXvGraANP4o+RMPIZBb2/4Pg8Y
YROhKdRpkmmfy7aydmenpiMmnoWS+DoHQiaPpt4pV9npLxxvN78U8lPCkS2B9HoP
gxEgeY6ggAcZKch2BWxaiaQJRsF5MeS/m/3N5iOEvL7tXURAILQNCvkZkGDAnmf4
tAnGC07PhLOyhr7M2vbxq3N57n9zmEExmyVChfhrtHnvJavRJmaY/2ITQfhrZE7a
rx+J9uT3WJcTcn6Nr7x+P9nveNiUCTJvvkKBfenwxXuNgk264ytSriNgjZ7+1upv
/pp84KhvuaimwrL6tGQCKDhKTRGDxnuVZV1xGdujOJqb4t2cyY0pSBssQtbHaN1b
zqtDtnbFLKgqIacjWagM5EaOYGFC94veBVeLXgLfkYwmtJQfnzKBwTawmTzedYx0
pSEd2vsjm2RHHNvnKupQ4j5FnRAteWbbV71x0BnJU2eTsXjEejNtdlNYV2m9h+La
Za5JhwNjk+cM5lncmkmU1pCMgxTXyibJO3t9GiQsjHYsvcEsljSeN2ljcwLCAzmX
3X4Pn6QVT9EuOBhxf4tVRVJHibjvb0O3vuzV83/otaAXfAM5T3WoDUtxst05sKRu
9eKX8KIa2+cGa1TvFkStB5TxjfBP6p98u7W+LHruynRwinnaW2OoACcBI2cNfDwn
T4JIvcktGPvxOOWxCL0v+H0hhkM1WevM23dkSd456Nic58iwryZxRjsAHfbCuuD2
Pbk4MadjSrWDc8e7aXDM89EyfbRuN0Re7KkuKYTyAP3/SQUjfv5kZi1WzcdvyURJ
cS972ZjJTX5M5UIzCdf5Hlz741+ZULIvAXRSwir/riSmi8kT3nSNP3E/OCarWBbh
nkbjvWSOp0kAqtB3hxpFSzEH0CvBxMpo+zBhi89qg6IyHiLnYJRGPnfceGeiboF8
DZoj6ROShuwxoVZ4kY4I4jW1VzpA40ubtpd5EIlKVpQeYH+abudwKyJlgIKvEMMM
PUh1XxxlZqbJ08ivp3lDBLRLdF3OZ7eVkYDrf9t+uKzcqVjD7vJFSxofh3e8PUmL
s35YFXn7fdL1Nz+vDGG25lAcwhZPbOpfhUb2qBZJpq8R84rHZYroppSVFS5ni4tz
U8+WgAIE0qlwfB1gff/yuHebndPPtW4SuW26GWP0dVbjrdv+KDFdAse9FOEWGpY7
yAPE/MTGXB7kU+WZxb9U+Av7BdmPQBwwwjFA8U0EiQYbP2qCTFL3kyVKNtqoCkJd
6XZi3BZv+cbqyleq050zAwGA+eqJ8g2P7bsAfXxOJTyRUaIysTBipaiGBXMHZvYG
laQQeAPw5aZa+CXgjB3Sb7raeoYBIRb0SkIgEzv7m3opIuo9fQNkb5xbz30gQLYB
1OLrFfT1SQM/RNjOvZOAzKFPuvd676DR+TYJgPQurzp6550j43FQe3GRgtnpmXTY
ErMasCxh//aNNAqcBDHT/EwP0bZonc+homHV6u6uSDtHW2Mw7rAvVoK9FQLa1SYm
QWBgJLONWsFMFS/qah0rmEJcZQV9UHdpVK/LFXYU0jsGtv2e/RzBDQASI+C6IciL
7K33QXXwXMVQaQQiT+L87dFAUPh5D9Ku621sXTfvmoRBdeGJS01sQYbJEErRC1N2
Mv/fp9L+ILiSAnWuVmktzKW+tG1rTwHgJ9mm6AVxLiUnUVSqXoczCHw4N9dF3xdP
M7DxcekQKlpIdwm32DY/U6IdpicfENmgC/NX3Ss0Np3BeuDxp1QCp49kaCz8TSi9
EeB6cPzvKutZHC7WUOtxsfKNG2fbZux5Y85MZlJbq2A4ukvBk2cSFFr7vjZgR5Qq
CmNGUwEp9dcXU1r/uD1veHb7umYYhww1AsHWGbl/aVL5rbl2Gp7fiwau6NYIalgf
ReSDqZy0wR+tMawKO+BsRvA7HXPSvOybF6UUmZc4hyvUnxMjryRHHjTujiaQfwVG
dDJYTvPaPiqQP9AZ9CA5Im2telpwBAm49j72ndKp6V2bzsxIVphsxZAC8G13G4FX
keTXSfIPRkGc1G03yegoHH+1pSdSVs59ZUO6ed+rz6LlHyHLFHd5SZVKAIn4k+8/
9YuVLHOCm+C66+Vf/GBzp2P/tQC6p+PSYXLYs8Y5h1Hzw0rQRXRKsAValA3d1BXN
4MD8dlMzSixPoN55EPRCKRi2azx5K8mhWuHIe0lcQJWNCSoej1WfAyZcg0UheDu6
RJcOvhIjsVrNx+a5oF/apgGgzhM1EVr3V5eF6RkwqsHnew+U1kkfJhiMfInygdvL
9+lhye7S7WXtqr7YavEFElNfOSrCH5UcSqd806D/jhv8qnxpfYgCok4KoEdOmZ/e
qjji/ls6aujGAEGFdu8HDhn2Do9uQtTrmfDvp0Ae9qZjlOEs5DF2sX5HCvKbpyAn
ckAf0udCApv2n/POM4Ls6U/qnmoyHZPiVo8jvLroH1+ZaaIJatK/CydYwCfEAFu5
utT1InDafiop2FliL7CIy1VZZ2vY+ut99FbK7so/Og+cKVkWg5m1HPDJWcTPDME6
6A6Y9Lr7bngWESROpreG3Y/C60GA07EHdzEdpp6MFWYLM4jO5KZKh5FMMBsyFI6x
za7SNakMIbkyT5t1gKfrQ+FqpAUIrtax2eJIUWTwD7gS30SoTWTNOR1wQlSZ4PTE
iA1JtI2yaAVjyilCmcSzD6dOMBDHp4oxJGUCaAPp+Ee9Gkx083YwezaeEiCKXx83
+/M7L9g+Hw/HRiErfmmU0EGylnaRS61q2rIZKuKyp4UWXCPyyx98jYiJY8K0jbfw
RrcZUIEp08gPZNxipg6DgBNFNGeUQDD1Gu1HtQPs87uEToCFUEBp0GPh6UxDygKN
2a3IzM7VDbw6Fkvq1RtF9mpEt6TEwX/JcsxSYqBNPd4q93CB3abm4Uoq1i2OuTE2
Eynaq2Osc9B+qkMa8xQNgZtCtwCD643uW2GVWErn7X4rPND5ACPnWerNLqYIZEiB
n5K1BBWbBfd8baMJyUGTDJ7NvEuKCm29VUgn9pCjg0PeMZ8sH9KocW6BwY8hFCUo
2avmaLsNE4cFn091BiP3ev3MxZ+M7W15yXfjWftG6T6W0C24XvhxNJBhyCmZKPbq
FtAc2Vdv7JjsBLV7/lOOxk/a1sXltxVdTeLRcftFlIvJnfRtEK7HBUkNvAeW2Qj8
ZAZIhRqL1rcluIsJ/k0ciIsD/fEBrIX+OQUOEW37jk+vWvAwJugBxA4jUQdRiyHR
HKJtnIBO1vEJ0FtogP+PQqs4T+twotDvV5iAQXRjRlEWKZRablphXsprdkBd14qU
fa/jxAhOmgY6G7sW4WdDtVseCKeY2z0CPFE3mKDM8NGuNg1MWGqQHwnZRAM01nlJ
k3Y2rAPLvuvtkEzJQdeRkMc4/pvprEdZ+HPaPTh0DC5DhqReXDweKOXRW+ePJ+MT
2Ahx1e+7578Zc7vRqyW+sisLc6LspFLrxUbnP9parRGpuXWlFlb94zWojEW6HkUE
vG9bO0wVpFO+pUNKvJK6YMHPIL++WoWPIkCvgED4pWgVtQ3rpN2TwAWWn1/NF2NQ
gysLeMOiPLnce2lMzjn+lxYJszIbQDZhcO2N9Eb1p4XBpcSvtI3E2Y3IYaBHsv41
4YwZ5txREmrYwRpQK2lFDL1U+2pMorC6mbXP7UY6mae6P+4uf/0wPcFdPZtED8Ot
k+4iYlt8UFwLBbd+L/RAvPJZC7F/7SFGH6EzZELP1N0kVKCyon/Pite/BhJMdLlH
zFPNUVX7yfUaSKblPhW9wnCdrT5QE/t2hS+t4dvV0ApPysYuX0xV0frUNXBtBeXR
YyfIfTqNsPwAN9x3NffEcxsm9iieWDgRQH7BcCINB+XSWpoLwLa5QkOU179BBU7w
Mi9YoebxWEkZzGGcBgYouEIRHenAU4q2Ew6nkU2AVJNLZJiblQLYt9g6OSBA7+o6
5meC/zfpkN5EaZcTc5aIUO6d2PqVCTJ8LsX3kINFcZwRxHYeaiHcz7ZBKeRU/LTf
8IPOTNe/vIAtuCsbSJFZlmYfIc/KNL4UnR551pxdimfbdpyiScggH8vPoqvB1IEy
YBGwn9F/TgZQZEUx7Q2IaIAo+MkhJ51Un1yMREGAbPMGmf5F7jhB17M/5EN6RZFy
5x353qPGCbGpQUsn3VcbgFfMI4D+gwgTB3Jqsc2hiC4+9BL33JqWckpl8aMbJ3Vo
1CGqQMwjEG794Ou0aTTN+9v5md54BWaJv7AjRiz2/WGKz2xmom6XCxKOIZA7lWMH
Rv5sTSsojQy9XOtMnyahDTGbU0EzKeZHgazsgK+D8A7CqvU6514uUGrpMXywKF5A
60L8CXuPhGuV2gSjLodLpgOePCB/mB4gS5BDQ/jzwibT8uwqD5CkV9IxqjStrEBP
siFCHm16p74xM7WL2D34MfaWiRlKf6nwnblosrSruFdiZP7daYWv0EikW6PfkEmh
0kcDcstSNAsmjIPiuabLZWeP9y9uY8nUjW6qznD4XNAhDLC+UJGiYO0tt5dd76NA
c4WH8I/9yot26rMwTmPdKLszVvPvVYDAFCdxsBDrRr9FGLgngBUt5KgdDIEHq0UH
2wgq5kmHNRbdowzROM6aKQpOdMEGX3/oohLTxjH9nzfQCa5FJGI+RMljU0p5AH97
V8Q22Y/2pUkNpUuqOmWd8rNcAw0sjAqXmlPrlZE4m9La8/wplElGNVP8wg2OfWrT
r6GNb/xfDVGbatumcIwv4RZweSQjvGN5Nu+dzPygwpZUTcG2Z7S81z0QR8RHNb1X
I6AUSPxAyORWZObhTuECMryMFzQJuI/jmo3yMc4oCwaZrfZX9D96LYc03qph+atB
YmMDb2P+8dJP2kYXIN/JOmB3OKCbEnRnOyVBhCj/TwdbXCEnYPfb4uDWvJ+pe848
sL9WanSIj3XC2ZclkH+LLoCch/b4Iu3mX5ZenBHrcWskW3x3N5gzc9rT3aT4jKcW
pGIT/uVF7vQiKpvEoPDFgFCbrdmmGPrTXzmIxh3M1aOUwn1PqI2XutcKWlFKTc54
b8QBHIRlztXCRNMqcLEXV8eUKNpjHhXfuaqzN1qQsrB0ib9CdlYQm125tdYKBMBD
RFUA8Kdj9Pr+dHLtHXe+9vvm7kFzKGddXNGkt7wYc1nyieI7VnOU4pX+ZZcaUHQL
qoCPVFN2j56ZafURCHxBEydUWUf0snX/6WkqZV9Yfza65wlY2W1ee8CdVACiRloz
DFWcOsDvdZXT2MNdzBuHn9AHfFB1V7L+y986In86tzdEJ48Gf9eQ2wSeHIl2ETAZ
UjxxCwuGifFzmEAN/kJhkujpqII7Mdw8KKV0rYMJ5S9mtKfUHHgNC0Asdr6fV3Lu
m9uCMtxGMdJIycq03pPdaa3FUsaBzrcjp5TItXLBeRY8BRsoDQJsGPg3PKdIysRP
RK9k4LY+9KTRW+BuL9rn7XSU3lP9u5PJhI08EoHhdCJOoiwHQd2LeIg9QAsRBjpK
t50L9vc3LbyVxu9Erj5oT4Bode3VFFi6K/pIknFYOsObQO0buzEFvQUzeNusm3n8
MzxmUAe8SL7KWeWVM/vbOfeJ7jc5HHeJHmHM3eznP7RGbz9gwCCt7Dud+J7aMLWn
vN/1CqD0n+DXyG43O7vp+mES7VPKnijhwBumiqME2hUW8ysh/md65acybeNGUeBy
QQoiXtHJ+DsWH5y+NsoPUQ9YjaRi2IvkmdnUh/jk1hfvp1OHkDshBlzwRVM4vk+v
V8Th+kYdcxHJp3jZSHqXzSVUWgD59EX/hmUGCwZNjS1ZtkgTNQqFP4HzlnCAjBi4
JJNUQmJm5IEcrValr0n/sqHqu37xtsCjVcdCQyT4wo1EmqavO98iAhcY/zvFK7XE
56j16yPYkgX7g8t/dAcRzWaSj7XFcaQI4XYWKi/tGShXq8xcpCZhtJRaLcoB1tZD
2I31kcitfPyM6pnMuEBKinso1gyNq9FM2frq/XcvglmzKL7q+rxe2mbIXBugvXK0
NbjKXPlOgrblj5iXryInSqAt4e0tkwVrw3nuUN7ISRaER4GeAkdnIFYqteDv32Rj
X0gmOZtVSiKjSuYT2q0NBgaebF3apg8DPFPr++BS50DzC/6tsttAg3ApLOe10D07
j3/TB69JlOQlgsfN3KImy0bCmQLvLA7Yu0IUEJjfsYpePE8KV3co0s6zDV51xN4o
QLePlWOTUY8fN7tigJ+dxhPR5UIJbVTOmwoZREHxSY+oHasju9PmFRAIGF637DxJ
HhlwyWdjnZgH4ocb/riTJQWkK/DYENv1lDCso4xTnd1Guhg+jDoWW+3UazadVjBt
MxGlA6Y8GrCDROvjeYxi28/VSUYE/DAsMIjmDbN3WtPjh2T/86PuCVlJOEP6bwxQ
ty6tQeBIpfopwij6B9NxSrUmakoNQhgogyF/xSTVzd6lieQVr2oFzdFSQijT01gm
NpDxcU6Bf9ylim7bZen+4hzAyR97wbbejy7wp89VHIBZqRV+cBntXpKC3hJz4A98
A6t9f2RTg0Rdd/wGazMPBAaqBDlNKDymMFS0VTMOaIQpDOD5FJQFC1O9MNq+xyFe
rURiuYl9O6g2ZmV9XHYaQ7i704pALxosq5S81VETIpw8rOZqit1KhsQUDAS1ole8
CIcbacWuhPL3al5GlAosFgv4sJdKKrN6THk1v3aKP0BGAREfIqsp44YuBF/YtUbP
NGyEUSkLDRmL5AR8WOUZAoKz3wO7u8qKXKWYGw4zrKDcx2ap+rGjkvDJg+ZhXD7b
Z9jlpf1cp3XfH5dbh7XvMzkUbgTis14GpX6jt6ckNbemQBHumeRk118JlUjWBCXn
O5lVbK92Seo9nHtQ0JVRqg2LN9+khNlYEx9sFQhVea67QqL+UgurHP1EkXU0KoBJ
JIAc8Tsxz4KH3NDzwxAZS6g8MqGHIc3/BWsi4sJRLjWRHD+a/4wLyQvdtvBZ1RMg
mFAAWphtQkytpaAlq8nsDXk13M8iWRtaPPc6wUC7vQpOOw5+oH0jXcClTYY1yDCU
mX49+BZK69Rl3POB/jh+ffvt14q/TPtIFExYps8geEfW/aQHeAFKABd+LuTRuhL1
UXJcMjdbl03mIGMLdWqUQ1kCytlHITe6b0LT6MgDS69NqcA1Zr0nncShO/B71ofa
Oic/u91PY5onM8dMGnubFflsipQ8/SGWX/GHbLDFLJHP44vcCYfVvG8+MZ55ntIu
9y3CJf9aOklKcdtg83ZECfv/uSRGy9lMygK3VjnRy34qb3T7YMWncc5X8iemzp5w
pRCeX5ysT4opdfZRWoy13NFjjceJ/XEbN3cFzdpHNRu+PwUbnIbbwfQ7PfNe0glr
v1NhSr7ocUWnil4+vIo4y8Rt24+gHYpvz7zsKD8YIJHHZcLZUvWkzu0sx6L5F/dM
F77dH1Xd+FmtqCuzmytiM1nBr4KE9RiJMsd6DIa5Ij7yvZHhP92Ss2iL/g0+Sfgv
uvsNtmDx+TWNf729/DkGzIiP53T6bY3BuhCkQ1RDbquV3H9MslhZ863CD0VIYN7o
2CC08/HfI2A9b+ycpcvjWWcZusTATueqRrHkzUDfH4QOyyfRjPwSiyjNtcbnW0gQ
WNUOAT9yQMbGvZxH76Spjjdmm/v46eOIdy1YnmBgwz5TeDLRNPdgur/wLZw4Sbo5
FqY0gtwAPIbRRlr6//SkyYIzkaxAhopKm8i4OKPG6KavIEfjJ8yiUnmhJM13Bz9k
AB1uxNSRJaTzsF9rEEgGCJZhxgsbH/XKwG4uIa1cylalJ7HymHA2FWovp2TFJ23p
WoPs1bkzHEYeA+kY0S/Kgeb6MpUXOaw+Rh7QMyAsPGdLmBExTNduWLFwIGnb1RHE
5wAVtkilkYPXdbNw8SaENQ/jq0oyHQ1y8m8gkqMmTB6DJUKNOEib8U0n9plQRtR4
4kZJ/x6TC/mn6+S76yW1RMHHtxJuPpMdeysO5cUcCBpdqHNlEwrXoJrvkPcYOF23
gYdZUtDyX6TGPVYbbvQhEOPCa0dOCbMvrw+lpE+u0BMGA7gBMTRf1GJL5Ph6N0KH
EYZbCCjMT3hCd6pworEZLcpnTa8i/nfMhvpWwqi27psCYA2fP9Tca83bWzQ5dNWp
iHuF2pCKZmZk1YOCGKAXFBMxTsIBD+yHZ2Za6dQIHetm6pTT6tCvEoi3NY/ZR7mf
5dakBls2ZSif733QfN9Y3yO0WwpCB2iB8CTUytRJzxTYLmSpK2VdYOF+I38SU+L4
zm0G13DDbeFU74y8Z2D/O4IMoNoDJKLDqdmj1aMMOtYNphm6Qsv6LWXcAv6oeDmQ
ikqGtSfFMWy0/hnNRhPfnov91NL/Wrc/jGeOnYBKO4D6jzxPK8Lfo2tPGCfVmavY
FLxDehUgzL9eYYN7LzY62uFDrNQ7zVV81VawqYHXhSSjVXsGId63ld7oY8DY6YOK
yMLJx+QY6L8CpHHxjPHQYapr/Py4nsjStbmkpVbB88s7EUUYiFOlYdd5kba+0vJZ
KHdedC9TW+2gYDMnamSjqHqS+EsXpbIEIniyVKELyS3huvPwpKAu/LPgK7rz8sBT
jRxXIJqSs9nhChE9QV8r5iwpLfw7hVVd4+cxHeH9wXcA22wHObc1U0U7GN/Utg1q
Iba/NJAQRAlnN/lv4iv6+GMYu+gR6Df7PgqAxEcku80lqSeTGGLVttIsxQcX11uH
lpKyldV/JHXiaYX7aBsVJQNJg4hnTeyxn15+46SnCeEORhxIvQdZDP5qaYKIsOw0
8/K5jqR1M7SRSkqqSnO/4pUrtABxnuVUkCfB669j5Gdymu5y2PIBM2oTop/b7NmH
yKXTmphPwptKY5t0O7bJgHpYqX17HqHz5IqCvmo7SqLdX9B8e4J+z9Sq/gWj13M4
90AF7trC14KmEW8gchVWz51wXAwLtdb1ExtM6Tysmbq8DdB7x4VRdnOiEyBLvto/
qM7j+6Zb3RofyZP94b4s0y8u6n72BdFUXda7J724DezZwPuJwKWlffuPhocyOARK
z1Ru9F9Sq/2LmqYe/VXDbpaCT4vzOERoYwI/SM7X/UjWzjMFPiXQVIulwLGzdrL/
H4OflOrLgXk1EEMwG4l2lAvLZIS8lhGEfIfwcf42ns8WfLb/ELAGX1xu2GR96mvH
VpPY2brkihGX2z48jq9OFlyZ1lBXY6jr1jrBMK5diKolgn5x2/xBTgG6gLf+xjms
SbNmBUBxQZ3AXd6SXyZxbNS+mebvovn194SsR+/semHUJkqjQqqxHeLVhWb4nUeT
KLwjgP+CNCu1qsDHBQA+DIEv48yxFn5t8G64krk9KAFk3Tv+8TKZDymc/pZzVQ0V
0BYzV/bTfbuRrKWJETbCpjdoQipMtfyRe/6LVok/Sk+oVkceUkMGitpcrtWtEe1v
g0ZfCNVC+VjWXyQSyOQOu9uINEcwdo1kIIOD4e0fXN6AV+r821dCY+utYPqnuk59
bZoihb3QPec2O5Jj3/qzmKGSJEqPyLdH/hfDLN+p01EHjKo/lemaoZry9hqzFITM
i1N1woh0gF1uxhOIPV7BV+lM5uiozaRXUceI6cVYuKdQ8eRK/No9Cln6XZGOaC1G
yID5mYXpamfir0VI0oA5qsAtTPJO0oHZj5NpnADgIKVHqMC9sFWAKv2CQJ3KXirp
ub8Db7B8rGazJl8YENoEXeDA6ZvEx6i2gloyXYqqE6nKEtEbFrOHdQ/LjmgcrJGY
UJ/UEUxzL93kgaEZ+eiPJWmA+2XYbi5mP0LeAlnjbRPpLpS9ZQ+8PhJRY915NBOq
WQwDdUxxvCCUTMU1IQfe8sQYZe+oAHTAKxPdS+Nb5seFhXysF94VkY38Rr6Z7lIW
HPOAe3+u5Rd1qyUj8Kr8evvtU6nFYGXYidbrAHAuIriqxZyM2m1IAFla5823FCrt
pNN/s2g44h5PAbvc/rrwyOc7zdqf/ctzMUWnmOCJXoHsFCi8Dsh7AK7buDDGkNrl
5dCRyCVfKUE+iWgJva03Qo6FfZ98gW5fmn8wLxrpr6OrXVssKhZF80O9PI/MVKXh
zBgoTTigHYQI9ClgrhGfL6y+ynI5GUDJ0eh+k1dj/qPNUeFz6FHWTNowZq0ioPXp
SIo4mohrfhbSNsc82OcxW1WUKnqeVAhHWNNFo1Y3dgdhqnPGmkHBp6kgeeTGmeQc
IJoRjBP67n0vs6LuYTjxYsgpOBj/YPgFGAqsupysVuYylTj2hZgbWb0AAGYP4nEq
OH+yW/PiU0TZ2VWlkcWZQMpVooXeemUCbD29KGgJhU3s85Lye7rs5OLuQschkfZI
fZ1JypzSivxxHCHq1aEcw9Agq3KmKdN8j9VQEbw8tDk6dvv5RZ4u6ZkuOVRlQfBi
fWWLH+fV7xb+HfEoKtWvAetj4dPbsGOehC7fHEVO5D8xi0eIPL9avNjRvSGZI7aC
1e22ih/7ZumbcokzJuhk0U4mxofMBHJwJZkfxkSg6Og=
`pragma protect end_protected
