// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UX1N/dNfhxETlr+KkijPsrzlB4uIKwcB1QUYvhNfI4/Ytuiy8iuYQp5gFSeTMwsU
V6Qdh6CoNgpCMyz2sPVM2rQQtJs5BGU+ZAgCz031VPPT7uF2/1TNA4/8wiIWM5XU
M+rgsCPC44ATmI+fSLOc2LpF3esLy85DejkpMHwxudw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26816)
285AV72bUpKu02nQdNV9Dr/eQejQIjdCuizOFbZvpbabD4/iR41FTlTc8WXqlb4O
IM4EH64GB5ikKaL91vOaxRJjufDaNPmBmlUld8YvlsWCFwih0MmOh32rN792yo5y
v5KnruJhT+MX1nGRbOagmzQvS0V8mHpFgc3OJ/owbTxdulViy1VQUxMFMrd79Iyd
IbzpDfjAw2eXe6ShlQ5XcnBOhM1D6EPJXMQrg4kAqenHS03Ea1bW/tiDhmJTzBaA
6pMOcIMvd5ciTHm7Bw2gRH+z0Gf/ob6geY6pXlbeZdZg2ja/xzKXP+MHnspp6oFS
ODHYqDKCJjuPgch3/9/OWVCu7QzQBZG8O8rutd0ViKn3FNeX5+yx5nNJueYQFkIp
F4rjKzTqRd3ziMVadN5CSS852zyoMM/FW+9M9bJJz3W5PidVs788LFUZyqveR+WD
36h8ntbrGwt/97FiSMDGF7A69By98RruagccE8+tbvMP96i5kHNa5v7QixhgZ+Fi
0315c1L1Vt9/Mdc7zmlWL2aVgMD3+UDxYvmhqnJ8Rk4W/fxfx6lJ5FgY59shtUx1
HTLgkelx+dVmgcIrbMy8+PisvYwDARtC1EAB/Xnra898RKKT0LsjnJPQjG5BfnoN
j6S8DGpjHm8W/39Zux2DrNt5hTf9MMB+emO1+zsslJmLCXR9e7FAt0RX29p80tr2
WAVPd7Z94jqWYClEA3jz1tmV1Yf7A5d6pExNsFgz1ASyt9VihqXmUowTY3Q/bohY
PgGNdVgeuxCnNyadwWHwqOwo1c3cGNpq9+DsvVbTFpFK+uiffLYeqgk+XbkisT7h
ipvsoY5u4+XFlgQDb5WPfwuJaGNbDhP06rXn3hZmBoGxoBu1xFy8EYoZjzwAMfov
ZyjjNWMMEpZ86dHjBCXD8YlkcIstFOV6n0tnvKZrpGUHjl7v21BdydHZA/RSCZ5P
PG2P/vkhatLJiI8ASuAuEtAUQE2GkE7Y8IKHIo9gJv41SlZMybg+aZ8dxiARX3Ie
o++y3IqrYNGuaF9cxxyyMB/93qORi3W3zf+zpkKdouZU0rYoS4sahuG3MaSFhKi0
anVJfuw5Q+ML9lBhS71WngJkFXCzJj/timaPnAz2b8b3IpVJ93C4VCbVGwBqNsdE
0v14q7ZPP257OozBycLbYPbGBajj/FSjgIgiWupoN3g5EiP9jSMztpXTncB2jAfG
/Wvd+90RB/P8yPQRsi4iM97Fb4p3i9nqjsTh3hwJPRSl6AA9UaKUE8DpmoorRtDQ
iiek65+7Y4H0RPVdS/IPxwpEUQACOMuzzX8UQz0In8b6gj/N3as/CSTXv67vDG47
xojP9VDmi+164vlu+EoOCL82b6GOcYr6OdkyMORrdD7/blBoftnpZFi8KDxwv8wk
u8AOsgX42JEdkgSqk1FWY4uhJQIXr1dq2qay7cnCBxH5REFvr306e27J3UtqelBT
WF83FAtN5H7nfIAkM44/wDYePlZHppxT7NhPiTvgP8w6kh2FmKXgMRgSS4lXDPrz
clbmPRwbRctgquLnQsisP0c0hWKQwBS7e0o4wk49eY1Q7iUYgjcm/qrMDoJwVCU7
KgMHpoUQ3wmD8R+J9CWDjizylU/vbYqA/nQZ+Rw3fgBeHOdAPq45LsTuIPeHN0jo
l9rrGcdVl2s4gfAyOwU3doxRsxMcWgWLOKSYjwxZziBR9stD6Z4zFr3KBO7//JZ5
lfOSDxlVuVUNGNtuisPf4w2zevS9f1ob1C+qbSNXNEZ5NeOQTiY8b1Teb87jgyiB
GP+jQLS8dpD4Em0OUH+i7yjWdJ2tNc938Q2iqhPWbEosyDhV/TJWfkSo0beAbmAL
OpEhf/in/XxdSQXRqwyYuMTShfvsM2invhLQv/ygaWxNUanQxFUuE3WUmQlm0cBx
Oi6vTtoK0NOab+1HyulKfS+NDp8xFxqi0QHcBGKPe6Y4WHa561QGv8Tt591rA2lQ
iW2OYz0jYROu///D2VwkuBsTjX7S3M91EUhR7RWzbfwrBjZWjQ7mlY8RHj3YwCrW
XP5m92u1wNzSmqiMi3yK+5CFRyRFW/ulf9UdbZzq1ST/ksMJSQlG1oCqPNsF9e+S
od4FCN1xJEZWt0N6yoB5KN0IKgTCOYbo5CF/G1OPqJyFym9pUl53TO2n1F5TYCJ/
oZolOMd5fhdH0eRbsYlhzW7MP973eeSDifSKsj28+0KG77N8wBDwgyd1licv1UBw
FZd2FoT6lG7Mzl1exkiJflNWV2C0Kx+6aRUMAwCUFF6pclgocPp8AgK6u4ez+q2c
4lfYjIIB08HrcvcKRKTZRb39ko69BN/NQpV3NPVXMUfk5KIm6yCsNfWJ9TjHPd1l
L6RR60I2CAOf43HYpPx9UjmUT668+HpKmvvnGac3/MdPiY+bYC/RZAQJxItV6rh9
1qwaMof4vjzWYrrYSBAXkwx8U3ZMRPErMdvtA7Mc8yuIMr0FUnNSO3972gjntcdu
YwQKobw6IyLpSufiy2DVVNy4L67JrihaOAk4hgMKDsCVXSEYuRZoyqdBXharKeMe
u+TGTZtJxkpdKwqoxrA8YmO1E9jWD30XeySo3qyG5V4ewuZByh4PAyUvzhppYO1B
nbIreunUigSJQeUDdFmRztw7GXhBru3GeHAe3IT+3Mwr8DbzWCbJi4j9v+UwqT98
ohpao4RqI6eqKn636UBtg93/hOKOcpV4rzszOZFgsqjPzXjiy6EPgc0LdHMLE+am
bnNvXIyMMJLwM7ymVEaOw5s0vwli1TOlBGlxdp2vStS4Bs+e/JNG1Zrewy1+8LqT
H8s5G321cEuCIA8CPIris/dUlpiIplreQFSWhAOfvNRA6YrrLl4m8uDa90BKVh2v
Z/mmoN3l7toyrM/THyjTDYlJW0b+3sFvly9UEE19JeqfztRsNx3ecCok1Qa+lKm4
Q+7yU2VNDfSHpQCCuTk3jYCw/XAEHVco2LnPEjIb5mEDMSvQaImB8UgQczwvzMb8
WOmwJqKGwY+ANgFyvMe2DZNssSCfKDWknZF3pEk9MJM9+mb0ou+2whYwi4Eu/QSc
ndfVhTdnQ27FzUOvP/qBygiymrfNK6TkVzY5x4xMcRWrkI0AUHUjYM49z2t49FW9
BqCOfj0CRpGmnQBsZ7tV1f4MtVpIrf2hN1x/IjNBONxL1c7qO79pgGXs4owiECY9
tr6wP74ua90V7XKbA5wOQOcgTJ34+1gpO7fijJyRb3FgxcaPvOTTnF1q0NNEbcW2
u2ZnBucXhsBZyWfZZUQYpxrq4uNk+E2O5RI3NOzhSghn+VLQsueMkcJjNGhKRB5K
cyPHNjkZxMo+au41LtCnSa9UqgWI6X52FBhP7IuR/SUh1i+X/HsXAHogWfCcSOW2
u6OV7YyvRVQ7Pn2PNtQUbBb2Pw5y6P7wblLhpKScp4aXN3xMiYSj570xO0W0Fq2M
fg7aE1u5rRrAsknZUj7+5kzUSuBmFhgN7ah4o8PzR9Ff252qDecOa6/6OtxOB1rn
gi64fS47jkwP8wHkrrH+Gfo3qBSx+1icpfwnU74Pl83FFDnZ/7QV6+zRs+vRF/vF
DnRQJgFZNgU717P/NMAcG97VS8SRwLaoNUbT3CYX6tNklz5yTTtVd8CJXlQkH3Bo
cm7+sgYnwq3ail4ebv5HEkuEX3RfAsm0LzmXYvd1J/EJ1nzK/vuBsaydqyPqSkCu
meUEJtPUeU2L7oaoplERzulVkZ+6m/nFg/xIp0+I8I2opbHMPWOdbQXa60iPZN0/
GVfm2Nwrrny3FCJWoke/9d12mNcroU9N7YRws2XbZw/rSmsXLJzHBuAWJkBWGhCU
sa5jQfEvr5BlvzyPc21ewIainvGYirzjb+1GKkeSDsP59y9CmBaVS8NFKGhIkPbU
sx99HBREuYzWNrR0bBnqgLJFMZOwU7TLpJpVnRkxRg+OJS05f5VYhBJjRe6P1kLa
zcI+2w80zpeI8geSbdbYyg4yDOzWGtl3TRNQ97tIf6H8dcMXebSrQbHqPkvxZOlp
5I/Cy4Y10NCF4Q10s2Ea91MXQGU4cXyZgu7JP2ZItVFAt0o/VFY9HOLzR2exDkbz
Ms1qsMHCKTIx12mCxpV1uQ1ZUh3/OypxTJmJj8LNeIwK2sqf+qURHQndWzufrq71
hT8AMDeoj2KtCZjqEH/JKCncYzXfISc0eCdxqW8924jEI7J6Xq1hP89Tc6mVMT2i
ZGJzn1FZekodyUpAC46Xp3UWk41JCibj57cT85Zil4jgqlse12X72GqGqixhrRT1
LYevJMjrs6K+BkNBnwJbUWY9QsEgVVlFs7I6O/gY7P00fqwkW51VZ7nDCOXcUtWH
LhBP6PNfyXYezt4F8cxzlAPdbutDRDAhwBdJ2NfImZU04kJ9IyrF5IH2Ad8C5qfV
LmJbw8ciw0xTMcX0oRP5+l+fowA/HMeZtDz71hQqNORCPHWnc0yMpeiplyFVZ2xM
3w5Dqidj9lPYhZhDzJUvIkp8r6YAXdPTJbFJ3qMVC1nUAPGMELyzcVel14b+YOhY
WwvE05Hind9dXZdCAzZnogiet3sb4bEroR7kpZX7mHur5Vlr/QVufZbrCrojmk8j
NC4/Sq7g/fRN1uTkLCV9cZJBx6pYjPEc7d4odHv/mG6loC3bXMZWvQu3eQY1KAY8
ZyM2Mj27mpn3baKjNlg4Kc1kDB2sZPhStzi5f8mAgfZ1wzNhAo9puMLHSpr6Rdkx
4rP6VmNuY9U53vB0IR6D1dNWsqSXsImzBoo/SiXQNnBaWF14V4KH8u08A9e5Jj9a
nBwObQXAH50xOwgPgh+X+ahSaL8mrjhQijsIEPJdx1Z2rlWzWO7lHkf7eec0EeXo
iBCZSPLX0lbqLYgzrk4ZoSIhSoXOtNkMFIeyDK3LPRglSCbUFQh5W4nqaE9nXRE3
wx8Lj0DtLLHL4nSS11yd/TaoS9HYn9lSDAmEHz25wouE2BtjYPEjsH0qvq3/gedn
/GPRmbLYCZe28VJrUmlnqn3+wNNs2aeSzu5OFut0grYPCHpzEhv7qa1UFF8Id2Ef
kxDKazhzetA0+RhbrElr825F2x58Bm6bCiix+KHQWTeVJ6xIUjM8klAeLPr5E6hv
gWllcM6OlohsUOPWEWL66U6zjEIJOK7FyYJ7rac4t7nXTxjsD6iGOFtbI4UuCJaZ
xma9QNTRcTHwlxuRJ9Nn8gzEuruFTHTOp2Icszccf903qKcgLWB1lD8Kw1WgwPDZ
zRACL7TqjS2vWoarvCh9OsVGfNpR69Si/c5FdVDo2BKkCmPwqhIlJtBekLrc9eH0
ij8XXAdmoQb6znlH/f3SmpC8w94+BamHDlt3IqwThILLi3EDbtzhTqU0Gzl6+WEs
Ee74Hrxh4JYapdi/YJ815NsWqsrP3Md0PyGZGPNEkmusH/kUu2krHG5E2haM/ABs
3oK18UGIfLZZMPcdkDliodDEctLRjYh7C5JaPlkdvCgh9REjamS/9PQEPUcF5RZu
Y0rGjh6lyErUP+k0pOnAP72WDJNR0t8tjPcHXCD5mm+ituI3ANb9g9BdbTZncO61
3V1cDXdurj1m3cdu9W3u9gTQDxecVT63mkSNmDYa/Z2mVDl5SRafrkVgd2ZOcCQV
SUQWVXvfKLcldQWT8bu7BOddInyEwS1fvCEwlVJMIXKVFOl6QZVDQykNHWoM2p4x
m2eRJuX0y0ZLI3ppHpS0lGPVPWSNxJ1baqus1cKJkVYPtzzPGia/JIo+H/0/N28L
U+J2Mxvx1uKIH6/rbm5lTC/KWfmlfZhwmiHS+C3qojWG0/4IKDU6He2mbaG4X2Jx
oPPyK0Kg24fk5N+uaPsqsR43JZC8MktfrJkfE1Fw4xHlfUMLTnMLDFyYgRzdWoLw
YJcM9NBurXOEi/yki2+dUUsKwlovqPeQuO7WrT7h+1f+5kQHtllrvm8uR15zcYjd
KsmsGjSlvOCzwBAEy8xuN6/PbaMYLAYpUTmyfimaqXrn0THqco22wDJQugZev+7I
uB0UMfZUHqx6Yiln7cYnZ5kxx7ofPMzKqZA+Eddt2kafROJ9osvdpwE/EHrKaxmn
Nrb9v4Nv9yOrscuL0qRQmdpYt/qWbTD6uQrU22mxSvMOpEGEIxu/jFJ803EZNS0Y
fVbQnz9tOqYYIIV6+fRx+Oq7laVza36noL4k5msJq/ptZELTb7RaUIm6WFUX7svg
CON4p/WeHQ7dvoYhwrP6zi8U1DWdKDxaY1JA3KiNEFy07TX6yACYTKEXdmpXwNnq
3nvauDTUh05CasBUHx7lHv5vzHEO2akpWyFIGhDvRLyz8hGIZtugA6qlDL6oBNzs
ogpTQ1ZqKoFkne4cOnNAZ7YBip50NPoAJ9WxYT35e8+Yuc7j4JJORJ5XgAqkscHs
m6XWddM5vfqCtoZ6cCB6yx61jI0i1BdLVovjytjVNaMMEHDDKoiZHfoKSHXqJ2Fy
cq8wttrqx2buzosUe2X5gx2mWz2xH3j51lHYk6CEx7hst3652aVRRa2hGFAED/fF
CkJuWjJMgi8xDeKvaiol2t+bmeQqeYDkJoTn+x4UaokgrliTSDrBBspHuQyBPuRk
I16ZlXbAAgL6aBPMobvy2t/wYP944wSfRf5ejrXKFs/fymvskxTRhqX/H1FyXJ+O
wgEYXfZd4R550YRMstISdELdz8c5TSoF+kKO5hOdpsv2LroSkkTY0IPFtrELgQTY
31H10TYrfzxTLnw1yHP743cFdIUFRItBux/UT5KNk5Jj93Z5/DSNEwujmRTQatSb
vAIk7dEk3QC9f0LjrTANwq/W0rN6z8ommnm0kkK5h+qibnd+xMwFVz3rvYYDy52i
6zc6iITRz0hDMGmk058cimRLvRDn1+rRU5ylrNB8amaqoBLAopjKkfb5Lnzg4j+7
Ush19nbuDhA9FUIH+rVuZ9Nbb6xzaCLHgANYESYke1zm+ZSiXqkpTt0M2ZVf0RP2
H1tqg/dFOBUWbeOLfqbeIKXA51hXkwKgn0ySiHSBV3QftxGMFwmVH89bJ6oViRwO
Xh2E2ciMbKWlCs9pdsR0rVmKU6/wGd62Sv12wrKrCIXCAKj1XQH0vA73h9OTtTcK
BZS/V+djNxxV0SFG1qn1XqkMKfbkkJKtc2JOzjN1vUigWNtW0l8cDcNjaUhKODL6
Py0bXve2KRoGZOzeX4zbsust4XLK0MMf1K5nU4LCQ0QJ1oTv5/3UWLMidlhkbXux
SXN3pEPxgHmoGNbSlLELWIJtSQkJnMPTe0rVI5UJpZa75Gp+WLYHArIoxkD/i4/A
cRyTW/8NkukvvdZoe2jALhnPX30gfyA/vXad1vlG9MUn1k4Wdh4xSK7qIOUEkYug
72s4pbK8bv8hOLREPVuXDyeIYkbcGG2ZyINYCdjVG6SC1h8wQRnZtpodOrHb5e3x
48hCf1/k+eUmBi4vbyEertFBKGqXEP/afNw26w67HkEu2zNmxgyCrq+M3Y8B5Ouf
vfTdIMzvAZHBMjOoujiRGX21mhsN8fLfDq8JXyJ+NWoMjaO7RiamLmH2PoJPnCx+
EUXqXConAiZWdSXEztxTqB6oKwh4/4IH1/bvsn11bQQgGCZT6QU9wduXuM4ee7F/
7pLbThIckljKQpQYe6x1+xebzFP6mD/rTGSUPRtO2Bi2KljMRjQzA7i5xBwUZk2n
iGIvde1DhzgVB0Zh+GJq1y1muiiMwiU2s/dPuty1i3ytjSR5qfo+RkRRmH0tKdOw
cpTluUUJMvgWt9HFGs0Ikj3dlgWRMI6QLIFDLgE04B0t+mECUW0I0JOYgHfqShuV
B4erv8sDXAJrd7bvkKsbQOFme+L6NfYk0PoECfloM0OMUvLtcuQsSuxSpOA70Cgl
T94rVsBgc9wA0pZahvGPL+vQ9oOsyYoh/dD/XgeSFR5KVZE6LYPEq5ZmgfwoN4QS
F9NOeeuL0wf1GCX5TneJ+jEMlADIKT3YxtKB0R93mvF6/CjP8lBP9Xkn7jbiL4kN
s4M7BHG+wJH8iCCtcMOMkRu0ejt2YuazwabWt0VgIISM8pqoPxBmQSucBi2ltD84
XgzUlOxSWQ12oE6aY4/VX2Z01qwggI2qxtBQss1n6ZL4h1LtdtpgEgztIqrn7w9+
ViszilPsFQHTt8oP1YKSq+pzL4I7/t2U/nnU7sd8kEwCkGrVJvm2dCtMrOGe5fzM
Vzb9O7arRu+iMJiEqm3NJt0WOVZPG0StSTEX0sfBUUfFcxuYnQmX3SyADVXoU18Y
pM/x01oSx79+PkBV55A0VirdF+pQPTO876Do8gKa9yjJevBX9un79GlxinrVnctc
JGJ8fyS2WSfn4T9lyUtLEpdDykdmETZWeYPgeTNrNJ5VVgun5AseKa1DXDX8tVqf
VIkmPgvQrGhoin4zHwQb34K3WncRQNrt+jrC4vqa69ukLGbtm3fsuPfweuyYP8/i
ufhbN1tniBbEI87fX6nNgLtXl4A2/tq9YWD042V7weG8SLTaZccxGMA3anz0QqfI
U7jue4oDy80HwoWbj4YfNV+Ia9Sb43rs4U7c146Teuz4PJ9uPWsO9sf151I2CEVH
66EYjaNBgymhWx30tKacmql3QtRyw363DVKGyxQTHWTdJsFnJ7Qd9wqLY8ILCBBS
VpJaOz2mbBbjAMOqle0dCYrzo9VobWTIu66ixhNRbY3HjUGJrPhey3PlzUQ1v2AT
3mmhsjyzLkedxT8qFJS1B5VWexFuoQADtUD7f1JFL/Ls+UT89wCmj2/EDQPOHNLd
seTfIZ7b7ZpoQNf7jD7wfLcBGCubW8MToM5P+eyGJQc1dJnE8lbtXCa6vD6ro95M
pBZs4QoYYOysk41BOjMF2wxxZQATbc1kddvTZq44K8IslEL58Xr0JXqVUfKS76oP
W1udGuzRXl3ulXNfMmaSjLAdpVT/YrSJ2GidsZRhV6WXkxPeeVMN/dF1XjgAnRac
NJXLFRjOgXghT0kY+R/1YhAzLg9sxH987CN7Y1MWenkCljTC81YX6s3zXM3MIb4u
ErDPFL6cXtCHJWydocWRFCbZq0H78Qm7DYr6SH98v+eYdmXwatPY9gdWPSCJO9gK
J4Wx0NnK8wG/WNxRBddTHr/65V/zbSYso7vg2KCtMq7JWMNdFUcnpOflbxCIxcoC
oXmXUxdSQuSAkR19SLhHFj7aguFrUn+MOlbIonKr/Ba4zPc9K4josowAPto/zPJ3
dDk38nCp9byJ2XkOzCXhSDee/dFq1RZXSRHdcHBwLHL3XamN2+gI8KlhNRBqb8P0
HLuh1d24TktX0B151ui2iWE15ccY3z2cTafD7IpbGpBy3FYSW1in3k3gDMda/VYE
CyHnAxDD1N05IAEm4LtA9XFfCQX1ouWPBMj7YJ2FC9dTmrk6a3tWUuIKQ02UKGRn
mw52KocS35pD961HWNZOVlW+fxwivxEQGXtozJHnJWTDhLuqqmkC/oXpnpO0eaVU
kykVDKBKA549kTHbsr+ruxzSqyx1RLSXjSF94YinW7sBxrGSFPfMsTy0neX4g3gG
MuFsY1nRMoEKesHenC5GkGdNIi1hxcPclY1gUh4o7mr/b4UmZ9j7JcSfLjwOhlQi
BbmNb4KGTaw/cQAN8gWHfWOqdJgjx/kGmhcVldYnlV0kM0CuBh0NRult6ZmfOf5C
SXml+CUbX53R/+cmTG0FZnjcKP0k1SztglpYK+dsKvEvFiVJ+HO48VmnH0oJJbjc
TlxBLoZsb2WsDMxfbx0UUfhzVELkxHniTfTKQtnLDo/2dNcgNn+K460U/MlT1lC2
7POi8S9SJoWzPDzRAmzIwm5ynCP+tHLUloGjj8QKF7rmnmWCsZady+soEYs6ynTY
3n5cQh33hdXDp7L2OqTL8U+27Tg6hMb8q6s/3+feZxlHbIO3scBqEkjKPbDuYSdJ
XHsRKsKT66yhCmMJmUrBZYUve2CFeqTXTHZz+nIRoqjQ7/LlHl9rF+Ne2e01qec8
MY0efo9q23nkxwlZ8TAgllMgAS/4i2sRNa7foJDtybJgBnYlGFpJ2FgYPTg3o4Hc
rzgPD1aO3Ahjp310TsPJ7ev+iD/d0+psZvqq3chiuz6xnbbdP+f+UHhuQLXXXNXi
6fS633dDC+lA5sKXNZ+fJRhbtZjPqdJPo4Orcu4jVCwKVzCaCuj1a3+gx7I1aFiz
8/+4pR0zcNvIoiSVvEIBdhAR20vi8Kra1feO/4QH/Gl34USiAxIzfUgXWKzRsHWu
VhwmIDdPbXZGnZcgIamfMVKLyE/nVS2GRERVL7u1GIkAAnYV9HG6OPd9B0TTbG3q
LmwAAkGHYMI0QrzCsIUJ61QF2Oc5K8C1kJfFZ982qyVLV7FJ6feFI4oraNLDZa9I
anHYBGeEpc095L8sq6AFOlM5l6qCKKAYNzvIU2SUQbdAF4LqVdm/fyp7V//CUMmk
LuRQsUcJ7HiWlAQecvnqNbF+Ws/fwZwKVn4SP9854YIhAFQpq/fbGLrjDB8aXkS4
w9vFQX/GmI4viYZ+LDqPoYduGZ1K7hoTgPRM5jcyXypVato0OCjxbkH8hqhubyoi
nIGKxmGUnktpJvuMfcCsd9OdD6GHgIOaZIrjlvcSYlpL3hBdnnTNLCkCcdL2hck/
RoIxo7dRsLTIQ4NqThF9f0s3/t2T95opNUR/VH/GnJL1vmNFQRtpsL/m6Qy4GKkB
1OJSkkGktkIpU8/AElZe8tIAxHltmPwEFWgXhRaNXJlQblyqlHZ3fD0/TP/SK1Ui
MwMtxXwQMMMl65BqSXE5lttvHQuNt+9b41woo4L1T9B1WB8+swzVCn5bsloI/PVz
iL9nXaX73+htmCDF3u9m94AjY78SdZt5QC/OtjHA4U2UtAAXIAcjDGDKOLPn2+Ku
clb/DTw3FNwPCpB1mi4ob3XgejpKHKrJkRFhSLvkTDIVN6hkIoMBji9NRaU2u8Z5
UN52+lYVnMp6MABzT/B0atWfE9G9Z33M9T38WQ3h2U4EI/xtVdGVWWkRunYV28NT
rl6P8MphYeF92Y01jKtxnsy2PyYwgJ2xiixRsiexueVR4SWnOptOpTjb9RLkjUD7
ei8Hoiy9Gr9iSRFH+jCX6bl4s5AeBpg/rj7S8KyZHA42n+7sNPXwoYLJoQaVL2Pt
Rze8QRHpmCLJs3ovFDFw+70+avnZpidjd0nzOekkMNN73Uk09eumYvIcJjCyQeKn
8K4EZFND58JYJk3bONdbX2mqi+d6u6a7zhnG/ptfVH1pR4Ymj+u8DAjKfyfLjSbt
BOrf7q6bxW4nSpNVvt46KTARQ1gVnUTQXnIJoVxUTpL2q3rXWZPBFku6uPHfMF/k
hF7rDqJq3pzj2ciu+1J+RQ7GAHLKlEbDiy/m/KJrwU5WwobYqeYlrQdm3xmZr0G4
pCcVTr62xRmxJBL1f6ZdaCohw5CySNG7LohqP3if7QhJyDYot0V6VRbRTYUK4MU9
4rMpL0uUogZ7fsRhhwBveKA4D1VuSCNGNCuApWLmq00oPLQMHIhIX7UJc4T3hqbj
iEZFTJgqZQxXvqR/nE3blln/eOj9GNSy08runxUlvWcJghPrJ+/9WekG7BTZ3KRF
AM5gFGBMehWklI9fTIEsPZjJJuz5zw39s94FuFCipu1mxF9uDzwAT51c/SwtBue5
c/4UXSmeS2ntRZCFVWq2I73Dfgp40sFoN70NW8ZUiQpT/bPlOz5+MTa0Zby1pHer
fcgRcIvuyGN8TNybKsHGbx6dZiHyh9fsndO93ZDOPUh4Yxp1ndfxUtwLfxxRJNZ3
hUbMejlLaJSyQSdF3MyH19pjR45aHReogbBvMdnmW+C5rgRjbJFy3e9ueh847vcJ
ELh7+c4A6q4lBkAk3sRReorkRkehectVqIravAqAs8SsMrbLLOU/DfcNh5d7jq7+
QTaryxMQ3ay+fRIno9MKU7t25xp+iCQTCwudhDzQLZho0hd7DMbCFoqd8+cUNd94
6GvqqjlY8v1EwlSSx7w5pk5BbyECMcKDKpNvX7Uam8J14vGmp05kX3U8gUBacmja
gUJnXgP/YUdmm+LNc69sWN4CWOK86uDNHZAS6fplQXtiJpbX1kF3rVbde/MxYY+5
OKQX5FoQ60uwrgW4Hdu+A/pL0Y/od2muQSIL7zgr4Y3T7DtsNTwZbLW0V4KZR8GI
y0BjB1gWjBP6loTQ5XVgOJ9DWfv8i4NXKJ5aowCwBNHGc3S809BzUzwc5M5Qr4tX
JgsHBdPhraCH5lTA+WZOBLnBGOIWYJowVK4bcCGkBKCaewsc0lxe2UXF+9DwVKiA
sglmIan2p7poM365bUTDmXoyMxQRkcuYZt3eas7I7x0HWJ7VD/XKJdbt7cMLIGEn
bhamhQGjn42TgnziXvlXG4f2xHLxyTaGM9V7cKaNM1kOg3DFVd5YTRIw6wFuln/9
vYR/uTSrOnzs3Ep6ASxc0AAQfvst0QLrjP2wI+lI6ACuFvAWTR3GCn+z/bnQG3mg
Fr621aw6YfROqVZsgmycY5LGaJiWJuwfSm61S3O681s+qACNhG5JLZCFbC/rLfJz
s2H6BimUate/X5UuGdzGLoVUeftkxcuobGje+HXlJgCqxwmG0jCXVmDxzW9gAP4k
Wbe/QQmyRVwWHJv8nBzDubt8qdx6LByhQ5wSV0rWM6sUK8rn2Lk3f8A9kLxhDRdn
jogV8dFTSjEzDPeu+9Fm1arab0bzBZTzqtm8diy4xoHJnxdxHP6oXprzd1oWITeC
NhKEdMkBn9nMXEDpgHsT+iPUNuQSvv0rAH9Dr1XZ2ptdaEj96dQ6F9Y5z2hau9cY
CaQe227UO5T6o+8S6Z5CAiiLKHXPvTRtWvX3ploG+1jPNw6q0ayuqAwihLFO7e7z
Hk5sqKxRvTxrdWqMEWIITY5ZpIqeqFWmfr73b3qLcLpd1VCGP1GQzVFPKHxpPZ9B
xKg4783n6k38ehI3EO5yFT+pZKRTSGbqFVwPdAUUfk+h7JtuqOh6DAiGJ9qv0v0a
Qqe25GTLiKhVHyC0zZ4Q8ZAZfIlyR6gzCahtB4iwIF0t3GGxHQCtVgc+k80NPmub
AaU/GsUpnnhDrXu+tS5i08D+NUymuREFh4KfW0TQXBSLto2mR+m4LzalvPFwralv
N1ynwI0Afdbtt+6kbi3o+Y2hYqWKhvZ1YmtXMfAt7h32hh5u4MxDlo2acY5AzmOA
3ae6q10cajNNyz+PQ/rM/zaSZWr0BygMt7KDTgLI0QRYZsaeXbTj8pyGyASuBsc0
pSu4Y9BvzTFI/2o6Hw9RS2oPWdWh6CNzvkcLLcdJrBR41C8wiyZmNhR0ayRgFL6G
wOG9P/rJ5eBIWRC3RRqpOYdlUU0uAzh3N0lsMFSnXBBTC96tj1ALtX2vrVD5PikW
LoQNx1D21VrVtVTwgUiY6f9pTz3FFHrkUAVFIPdN/k1ER3CsWFi5+fufqU1dKQFL
FY2AddSk3HSHPFQlGeDt57Hueo3dLzVbqYmCpfF3l4P4ohahJXHUTyJFtLAISDeu
YkS62CgPU0I0pDSHmJHMg1qIEwIrSCJ4RS4iUlAASRfXMatDE9fY+xyg1WRQ7p2I
oB9LXksXxrxxK7BRlF9JViKCSKd7zxLoYXAY9pGTJkV96TvbvfQNxjmQUcFLiXUK
B77qhZZ7jQqMLLxF5P96lLOKprniD+lPFtLq0vL02K1nJdH2Pjsfh3nujP02oXev
4QLUoBeKePFtMGf4qUmLby6CmI3PnE1N7JgYTs4ue1dfBTVYQs6Uko+BCIe9vMZP
7a27HqnByVautptzTWhh1Ar+K4Bwj/xirAeQNa58nPwTjF2EF3CS7qJ6kXVMXdbn
uNG4Fs4Q4iRkQdYJyKOC1M7vGFauZqN92LQpknMQR068dCSlKYch+wWz1r0KLIlL
ycH/o8zMBq5k7xTQ+WnpBtAuMZlkARr5DevHFcp4bgOy4bkEEtYk7+1PF+2dU1XW
FnL5aH8hsmDkNoL6n6AParFsMvPtAejQLv9XlN63Slx5DICFM+X8XeQFvzulcRHn
yMw+WLp7CAJzcehIYQDAQ7NQ2A20QyZA4mTpGVFz7bC37KLXvhji09cCNrwXr64Y
VKZ2IRdnNJzHLdnj8AybMgMGanDTDusnRK4DP2HCF2atg29EI/opk3c1avEHHA36
FWYiSUEfSU/WHEXy/hzhvOzufVvGBq8tWz5QVQYN3UBJu1bcoktHhm36mLfXzAZp
FVmyjBIsnYZb3sn2goA/6pZCax74S75ft6wKZFJL4godLzSrseH9c0kTOjohBxaS
6qxEPJHecbgcvUq7kfogNZBwWJhp96unduZ6DWjd8Aj8W0iHFitUuHTXmdKy5lAt
1U1te//8LKWpCjSltvcqRyUvFY3KCiENsB38ErXlLOV872wVPqWAi+dYbniQpbv+
Sm+hjEGS58Tgx/RdBsrH4+4mkrKXhZGpJVMGuJt2H4Om5LSLH4CxVGKmsDybhwvd
9FGNH8E9zKWE30j59TZzNgXk+PeOaNz6e4jPO3B80pvewsnvUL5ZbwYT2nV4POTg
VTy0IS3Ndx2cex61l/yJPiZz11tb2yxsLPbuFcF9MK3KcmYRbvHH0AruZXJkGusC
t9D00QW/LzkFBzvuNoa1NjOEMHcbh8JTi5ctZE4oUlHxhL+mZ7s/mGijGfEl+Ftl
ry/LwJPuY1W9xwPQMjHC685YoC8Us2Qc6iZ9M1L9TkmctWjwtKZ8IepC9L85DT2/
LP7NEDaDVawl1FYY8N9f/bfbJGwttcmfCd0m88rLyz3ZsfY1Fo1khHvYmNoeCS5X
Crgp2cE5kr4h6tt4lodO+1coIgJNcNoxLIX2ae4Y0m+zY50uPe9cxjesdiaDuLcD
LQEoNvi1Y6qFK0NckNjQRxHtzKpWpdzoBGLJRLsZsW//fjn0dLawQsTb8CEAtnnr
2x8SYDQvgZpDWUUKAAFBnfEnX0sHibGCJnjuAhytwoDuVa/7MiukyV1afeXVnSbX
H9zOfga0SXWLd0RG6tker/eOU3gTn6hTY1MzYXI7/lyG4v+NiewQkFHo63F3rSb1
ge7soIqjoeA76QIbj3h0I3ZyoYlT0ijY1SqHpsBc9stMT6503v7k7FH67yGs3dcj
dTip28BnI6cxBGN45N8NVYyl7jxN+xGhzz/8u9wCYVJN++fIVQcLAoUqjX0lL7eP
lpNzIe1tyGAIa7dsp9lMQ+BeEpHBDNQWYSarEEJviX6UeNHPXDgRD9TX5UFLInSE
coFEKa0iR2ARY0KaSKrFUkPcFMtK7r0rGfxzAP/9DIOFOVPASo0gL7bUM7WpuxuD
IcklAexTQcwygR7RnoI5kW0jNRu/huLm/9AOJq0j9VVK54XPE136VV7jEgiauRgJ
f1p9X7+s41+ncLJX+L8pUhc4ocSUpZMykSITHeRAh7Juhe7Cgnz4U5cTZC5UYFAj
q0m6fbZi3euhAIh1f1YKJleDIxmvwdRio2Fhl/UpXUiJGUHHPX7NO0cKjPHSbzbB
p160L1ukm/iMORkRkWVCHCw+Q9NE1VWBsiMvEoLSLlGtQ+P8T47jTuTYP3Soxmlb
RhR2MlN8tYPDZievmdm0rKWGBm2HjWZPi/gJWx19Jwsjtl69wowLwOGh+LOS2vt/
2uB13yflcLnu91529cxPbUKBkqNqlPu0/jApVLEs/dt2vaYm75PBOHSGEwQt+Mji
hVEPgsWOJK8nXlVKujrVW/jsCUB3/Pm04MEDY01T9PM/vzoVB6IKI/NgsfaSWYIZ
1+3Bf4R/FbaY/gT/7gqYVLIyC5VxWBXTMC4wCUR2drvh6bZ2dMOlGT4bfqJguTDi
kEg1lQEyGeGL0eOpsFIaytBscu0lniqjt/0UAGVTlLzmDmuUdYTo0dSNeGz9LqgK
5koSbHoo5NpYmyPupher8qZkKKBKYKLptRBkXGLMjBrJGxONfxUSWyhvmXRCJK/v
1PrmDgJq2gM38ZG2jtIeMMLkEf7kfxBM0WM0kXVcK8PW+OM3bdsbD0OC1Wndz3z4
4TzT6Qb3ABUYjKE2aXz7C1TTlRwtLYZU4mZlXj/q31UnmwNjqwlfsRFDVXVyMK+R
csnTqEvJ+jXpDpv+CMfwRAxzuNqBqyIGWChu9MwlFaN7+QkrvSFJ3OM8MtCzvci2
Cfisu3QZYoPCehwRdzV4VckGGCjK9k01Rq9KDuzThub1UOBDfb7zWCedkUp5rzdm
aypS0Q+R5WDUE+ICvYCnL/l3cRv4ScOmaRqXREs7G2wx8UIvq6yOYzsKt3ONWo1j
LWBeTwAZOZcnWaNWMxLVOi8a//oD+z24G8/8gS/v94dIeWCrrp0zm1QJI+PNhAr8
ysbRcGVJLG6OcxKj93J/zvlhWcVvp8UTGRFiSzsr8BSkQxKYp3rR+Bb5dcrj5USm
kZ3qDQg1rTEjpZo8WLaQiEDTO8R+27igGoCJwh/+Fu6dc/+zZuLE2J54NdRQY/4a
kedSQFRZk6mQoFaIuEJqFxcYziptLDD/vEMvCoJK8WU7yD+SANMV6XDRM6Cf0/x2
6CrOQ5d5vNCi/AFvBHLPhon9M71cIXzMW3Cnr+YWQKM/1W90Pi4oUoEv5q33GasP
tX1zJJmloUM6ulD2dPjhasvHQ62DMD1hWNSfVT7THYC0JI26d4SgA2jfN+bzw1ij
Jv0D69jshSmQyzjgRxC9j5k66dxHAlvVcHmneN4O+hgY7KRp6Rurw+8zvZK7IjbX
di7M8n5igKpA+h9tat7tHpcN/WZOP6dXP2bOuOY/Rf8Fe35Y4FvZa3NcAHYnhZV+
vcdPflO2KgAMsaY2YqThE1fUKX46NXoa4dTmlmwoDazn7c3KvXJ8pjHnuPR8hzHe
FtfEjj8RfeQZn1aYw4EJw3u6657/WtpQWOLZhAfklOZerX/BZOZUvRAT9gBgJGDK
x0Heb9rJqmalItzBirilGHGeoeCY3hPMpbnZk7YkyL1PkVIzDdN+QO3YOcbPd2ZP
0cOqvH7QXyvvLGxLlDR6RTRviarTGNqIvJ+rQuLlKt72LxiwH2ghzCBm4ybPPchT
oa9gEryc7ajJoP/qV4WGo8po2Z3A3iA4/YUYYUj+7FKyUMswRl8JTq6uInMDM9xV
eVRh4Gs600VFjYU9WxxH4t21y7ymUBklOmJ9+7J0iW4SlxKaUxAd+zI72aGyHTb0
sF6680eRQGZVgRflYOFFo8y6d6HkMcmf1FW9+ZYkTdQ9I84WjTUJHRGCWegKufBg
YvcSsQQBQ89mWXmcdIO3Rgb6eRLAS/3Z//6xDg8JwMvRnIcHsHiKwX0BVtvGnfVh
qHc+7czgbDAsOZj7f1YWHLx8dBuSTz+xNVPdkLfxdzyJqH3JqOTHQOhqzR7qqows
WhMT0yfPXvId5vdms3Yxv2MBpHM8hzC8QxRwJepAW/xTSeQewIH83f9wuINYyCiH
sjdB8smSWpm5G0WI5/prHITFeiN3ImJbWgIUnGlqZtoZNkcbe1oOxBfoZWQc5+AA
GoVAj26UNsdLGxdSWb5PHMry3GWwIx1eYJrFfAogLxyK9Mu7KtAuKrL/cxoxdtQr
NUTC9bRnH1M9ha+e2rre/ObODKwuyy6nJTurN7usJ3NeyeNhefxfsUN7e7UEKh5I
mN7eXIZ/YJ0C0PJV/sKdbdYtNcUzD/G8AqUPZ1ovJXWJczirPbEkmluv8Vti3YsC
qNNBMowZ/oZakWktgjGVfUrfCjWZfr+VLIxdRcH6clbvphmejizSblC7b6WJsLgI
Pdsw7nUl50MSCv8venexWFOAaKDAO0MyoL5Wad9yx5cAK4vYQuZvW7c1T3h008eO
9n0DJjMxnVWRoGj26BPjra4sMxicPcMukOmbRgayd7N1g89Z1o3kPualornySDOA
he2yCk6gd593HypPdV/UDuk+ZQLiUIE9yOlTRXvuKvmJXdBP7phLQ4q81Ed44QDi
YqjFRF4c5otXfLqBjCxj5LJatHAeSAGl6shEKg4AVqsnPpO9/2g3LW7CqqENAp4p
PWZUoQ/VCz32OUeyEtRnO54wJm9SqbCNT/LhGsOvyV58fQVIR3ssBqHHyMBiLs6u
gD8aMu+MK3IZmO5trNi15iiy4rQenIQaIeOk/T9vW/7PH2IGIyU8oZzGSNwxYvc5
KXGL0Z2164h9d2tgvq7eUTJFDm5pbsa9u7syslCtu0LkKvk9uKG3Dm/AbVcxzJal
RLldpufjHtlfyZ9HZCUad+ogqonfMuvwEnt17X67B3uAre0DOJ1V8NxZ9X8qAPpq
vLIS6x4F1rx/4+9Ze5A3SkKH6vpBS2Of3YUSQunM+skKECyimScXEngkKhYVw5dK
ACVy7NLBeecwOisndVPfmvbCP+dUmRszozHK7CeeLofY84BQZV9kRqY+g9VtSl02
1JW5/ldzEeGgs5j/enlazpQxSx4BIMDfKyznudrRtETqeGcBmynHvmSI4arK+1FM
Ps8pUOgNMwLKsiezd4vQEERVzq/uoziACf912C/qGVnjY4wAtJx9xUftmSLxCcRt
0YVdd+RWH+7GaeuxCRyKCcsrXp+2u50DT7UtRCLxzsXhHNSoTJ3ZDpds2N2TQawj
+LZ5Da46ZJJ8RhP0LNRMn4K557EeEnMrApVTsA+HXx30a0t9x+XedQVTyUjn/gIB
yYuaLlqco2NIM2x8CKCzNQ1EIR6/3YssEb2lM28Bzub+nI5WfUhdAvs3tyRd0yJm
6RdJ+LrgEmsAzsRvZ46r5p661DjEnCDJtESuXahly42Z/yYebOKzau1yfQcPsw7Y
selTSb3HwzKOaBo/WnLvlQkYpWEBBPofU4SdYxz5+CkMEVGp9Udxwd+E2fY2fs6D
LvTJmgrbJxZ2R82SpiQuTgIVPXjvcA9y7u1olf+RkebqY/IGDCMkC0vf3iqb936F
S6Hsv6DQoUZFkfbuW2G9fQZ9acgg+xlkFRey1GZSwWP8vKyTvdPD5VQMH+5rsQlf
8gg5fKbeWOvu57g+zyVS3UqREcjdL1yv18E8VqxHP2Bt7OCVBl+ZpqiitxNuX1YM
EQS8+KEFq9+G8o7SxGwUZ8x1ITsouSCVwsqJwbZWIfmLu1EoNPRXk5qiLw7gphZV
pK03LFtdm5ylFxWrkz1TEhjHu/5C/NpBUMLXdsGiMl6V/6Za6ODqKF1F8G10VgHt
XDfpAkpJKvLTO1nBu8BI76+AwNqpznRfBOd3WsnhwRWQRJKq1P2Sa0sxVux81ikE
rQjuiaIl+SfObC/BXByrOfezgXhbieYOuXu1OJ9wYJYbjxOTbbCI6I9ANldczn19
kog2Y6+pd5TvAEex6X/qyFYwaFtsKUH7+1Uih/yBb2rCHN1wxbfHQorK6KhRnLIL
+wblqNX36upOp3kWP7IUxxI4EeQwoZRFZJI/dmpl8xYKpkpZXRnA9lE50DkFpd1t
oNTdFxhc5PnrzlJZLH/cwdtscmuj1YIXoF6uhY3sLSpEfSwfUFXZaGVTgimxX8/P
K8wUUKOYs3GmpbwHS4hZ8A2+cQ/tGlRPX3FSqvIr+hSaa4NZ3YF89QO8H4bNE/hy
i1hSfQb+7UHBl4kjGpdVo8s91uDpf0tu/YWRRBkEhR6sZN1I+GUE/pQ5oVCT907N
FYMs5FXMZo58offAk0qdLA0d/IbbkzhsMF7Blpg8fcGTVgH+eDcNofPtYMpjpj+6
pmO1ts5f6GPktnOZkb+QOv2/pApH7Lvodvf1halgOGHj/o0zAjWImcxIS7SmuLnr
3Q86kFTEPEgHfdNuiPWd4ZW3zYNvXv3EyG5jtVcFGxrMLw9F9B+0TgrbrUMYCF2P
USwHeukGOgYmUW94C0vN8MZFHgzPfxfXpdfZ9PyOAmWR/i5fLfNHbcjYsSkez3Ar
PPmj88pJ13kTg/PfSkcBy8ONl6PPG07hmWIdjtS0lLBQrK8n3eJSuw2F6FDzcAd8
0dAHWqCyqbh4i1UatemPBmC/lGxqgemCY7VXKpvjMsoEnBC4JWDXE4ATtyOuw2lN
9P5zgvK3WNyrp3wOB/krIEM/afQXz9YWK4UO3NWTZ6qcexK7J8HFBQCvjXSTvzCj
81tn2pIZIwUSrDXmuenuU90oghepl3fxswflfBBd+zxJoeU5c5ON27qR7ZbC9t7z
Rx0HQEyu1OpbjSGs4E1Om2QGrYQhYoQR2Eeu75QskefSVIanioMOagMwQjiVhsgI
T7LeGQlYFL3CY3Aeo/A6ayiCJKBjYiTOh04ks1H1tvaO1mFu3mXoSID2HzSrkwPx
uLICcudHkm9vvTBN3/cWMoaFd0WvP/OLNT3+OZR54BBAvgnaCxY4DG/Q3ffIcYzM
saoYrM4IuUnAWSysSgWmzdZMpLRSIEAdkUW/zo4k2WzErC3aZNADO3NCJcYhPzHP
JVWU1n52HELUJL/Qec6DDDdOP/GpSeIKoI/UdOnWB1YqpHEpZWixNc0L5tRMYiLL
vjTRuA0XA5rvswdOsvgpmpMPuLLbape1UKHUj7UzysLCJRkGbilF0jyfbH7u+4kM
tl+0+/S7ymjnAwCLOXTqnG2cPhIBUOlmYcuouJnhaJnYfyFoJqCDTAlHsEdGZKqP
8FgrlEVF2Wd4VfRdORwL0D93/012TdrGWV4MO4OdpIWbbDukVa6hWVbnAYpAQqDc
6n19DkBoRRD0KuWfAWQSvLZZm+oJXjigwmEQEDx1C5TGO/QCAQ6xWD9QePyeuJLi
QgnO6HpjAjTXSNzYb4L1b9IlCfFXP/OAIYttvndgY8IzwIPOMmskMxkuTxFgmtzI
Bu7KuoPlzJ5TGzP8ixqy/buSIuk2nZUzjAckPzikscKRjmOgSRS31LtWWpmQIE/L
7C44SJrK/b5RlRNPZtn+hwTgitBiWDU77SbY/HHLpCbGZRswU7YDdk/uz9Xzc66i
9bLpY/O6VmNvny0M2OVTGkkUhMhLJ4eKYHV8dHVUBRqtdWOHtbngEIfpvmxfVsMn
UE+dPCw7kQJAuLk/IDWqDXJ6KWyR5dfh5fe+oLdC5EbQM0yihUr1DOQ+c03FZG88
KBXVre0GcAZC6kl17TJls7GvTYQveJcM1hxU1pdBw+wIgEF7F9kGpKMc+HTBzFbM
7QAHSIFlA+OFThSgDBpdSTce6ua5nn5f9S1Fq29y9jphbpCyffwr7UrYPE6u5D0o
p5DCh4OYjSph9u1M3GWJjZB/irLWWQtkeGZGgSu7/LjixW7q+rVyAecvsrzRkXj9
lF4LcPbvpGVCa93SPKAW0xRHGZB2FQuDn6K8lDMJnFva16Ok1IFf80P9EPzujwoG
HFVuek6gC+ZIPc/HQl52Rwv5u6KM16zdbdRwMRMjkHFEJ9S7lM6WR1z+uX4H+v8m
OvgxfbxvKASM2bmfJP4LHyOo885aZn1bVxWgoKvnrpTZ/7ANBW9CVdKfg4MQ7BHg
ObX9sYfspZ2mxZdH+3ywRn15g6a2SPthdY/qHSWSwFuBwAwzcQtGa189Bnir5Ns1
NfZxS0ybs2l6BMsh8QlqJxOLKw9uCdhXabrXVBhNMDl/7ezaGHlVf8Kjhsh8GTuN
NMqxLuMzg3g1Qx7IZmBcRc66AFnursCDPDawM4sXbPr3HqBkg/FVuRi0zcAnskpG
fBWrTnZvdgKG7zgumZGZ6xQXTRMekhcZwD7I15jC2ReWbW/A7IMZ+PcyU86B160l
Hboa+N++Sd+RjiwpNAiZ9SApoKaBwoR0kMr441UbUc0Av0ckg656MhsUSiSKLBM+
U4YMdQ1gyKCv7l+F4LjLATEoIUufS3aYAEJJXhpovPQqDPS/xwCiVi3wqpKaTuok
1M167Kmnvly0nJwJ29qxLpa53tnFx9prUfF45yfoSGa83Tpysiz4ZcVj9cMK9IcI
x17uHGI/phmwisYi2jD72UbdlTfS1vOKrCcbkRMK3iV0oiljV3kNJFBjPasbRwCk
m2c+rnKE8g5/bdPQfbQ0r300vrL/7bhvOxsoOutf583U8VfO041/089eGvcx2adc
1KpdvFuVMsg0D9gwsBlO0sAfq5KwbMYI9gfCi9Z/vtvBqyqpXj9al05f5MkL1uRS
0xvH5zHvst85qmR4es+VHIyL+Oh4FgpkCjtichku53Cu8DnkD5cS34Bafxde6LAU
JXiaZ+YZdKKQu+PScj6+E6fYv4etGaRkXEIUSfWeJtD7IiNhfQZqMaerFdIvwqvK
wTS3KU+OZ/n+WFx49RvH3cTZG4u/s+2BDlHa8mwMivxLoe237+mxnaj3olQtdZWY
P6e8CKHGYQ6JD4DBgU0AwMr/Z5/Ds3s2/8UhINVFF3jmLKXqm/cZyy1taDLA3RJx
U8BaJ+c2Twc+XU5IM5lSoyBGgDLDXLOcux9YOJo0J8G5zw4B/jLbKkZqf51FVe8i
u+Q5ZtxFbLlI6KwPqNZngPE1aHdusjxfBaYYFZg/150JevMqFI+M5wWUyOnDPdw1
WZ0uXVXJh7gehI/KMzCSNIrNT+lPRWRWwhoynfeRj5JaVMNMPsIN6IokdLaplcAJ
c4M/gVAfMX8xLGlGbGceoSD9MoMVRkxeHbVed6MnjHZt6w2/NEGvAT4dioaCBySx
MB/nsx0R0pK2uOODahRHAMmLc3RNRH+E6xZ5dGGy0sq7easdvYaTH6nLUhSAv8k9
3Wg4Qy5SYZwpaFXarCpuKY8OTm6183j1c0WAti8ae/WSBH2pnrwV2Y0nfvQUWxz2
jZeeGb6RIKjeCBa/VgIPuIFjoUcVRlRDsmMa2GQgVjvUIyQPvkBXmzw2zIH7D4pG
uV075o3CsYN/JpF7wW6dIEaUdhlpsnx/V9R0Fxwyv5L+ibEcyTQgNthnDSJ0ZlE2
inWaIe+RmkWcOp88a+Pk8pdA63KsaDtUlSsueiw6glhpWJ+mfdExKJG+zCxBTQfe
gA5rWT2fx4RSiHmwVqdq8HoA0J6nUTB//eSBJqe+9b3V1C4jI7zKffV7uiBMJ9Nv
pkm8VLnIxSf3GVeU8J1ECzuWMMNP4TzcrwtKOgmsiM5y3wyvOBBOZQUyKG67wpHi
TDFASTCuPzOS43OsXww88UbCbcrBjpPVmRS4rhRCaY+3TARBWewSjk2S9VsO5D+5
03WCITgI6JwYS+N3FyP6hZaK53fppnvSYiyvTbldc8xoExo5JiTct38NWZ7y6WHA
9Jmz831dgubyXujyaRKJX/SOiQ0CLcw5Z/KDg+gLlJFdpDrKE0yZeNvXQ5tlG+c/
WcpfWBaD+XhBAm5UyzuFBjp6K0xTeRNLvIzQhklQFfTlOmU8nhwf+TIyT8sXhW9z
UOR3uVdGYj3k2hWaMv3IXpAEcU7cLDi9DPOoH8YaWCOmGLXjkZ6fM9yYMB4WuBTT
42LBPg6BJGtXFfkZF4nMnGIgcyW6n2ck0hIyjEGF0MR7eHcZRvfFCwOcoFV5JKFE
4whbV3x3v+Ytn9Jw2+qm3ry/5L20csOAFcQBK///64SSOpxXxWQbh+ByCuGWuY5g
uz9f1qnlfUNlk2N+37/xfJfXifvakh65suyMyD3qtIh5sjToX4Y9pigb2IL3ZrDk
tCPfkUkb+qunz/JY29l22+DHspMYZovCq96vAXFjGycLgsH8LwklOZqx0vg/9+E8
+AVO/jsmMJ/7b9Eh1+5TulgEOLE1CpWvVbAFHacudMRd2D4M7fNknr4E0etLB5a3
XkOC6i44vVzbPaDTTU+0BeHGKcQii0qvomnEhiUOR0bbt7yo4hmvLKzymxAPwVxH
AOX2Mgb2BRafU+n5QIKB+w7kGkqp2j85+V2v78qgXD9FP2iQgJUyb+CSoTHeeaqU
AJMvoGbR0z1P8R1QU50+0w2ZfvrtTaCaNT0Y1r8WzrOlZUla8dVc5RIN3I2vaNK1
ORHvpg+8b03JWzuiNLS6Hj36fTk6HF5wsJDt6dsE5n959A+CeoXGqMhXXzYgH2Y9
cA4BFBsrKtVB7T82YhGc4zQL/oKCJ/4u3LRGXeezDIoflcfL6U5+iZ1oOV4hkqcQ
ugo8BIPqY1pUrylf6gTpdSAyqxRXw2hHpwH4Wseq70Md5W9minyKZaEKyNVuoEFY
8YdPoftdMWXT2/PMEk+lsGTIMO2fui/r6Ihkjb1Ndtg9brSfEuc8LA04OQAuJ78o
To5XPMRx5Ap02pSGRhOUyTKjMarTMZ8GavYS0laO2zEVOVsEoCd9MZFUZZDrJcf+
OI2glPgMciyunk7hr+uLRF2enQckNW2+ytOWD+CjqvGXKU+913h87+oF7ugiB6ks
vKtlUzUR3VhqUWhKPuNpdCql1vsIbhLjNQkyx3rbGxMXDMXVN4oijJ2ZW+o9/z6/
HN+Gso76cpt6Ugrtj6/oO8fycAR2UXN0K9XWMN4g19Gs5Rfp1zHWHkJ14nwW4+qR
Z8tAz8kfWb5CVcC9r34dlbKQRMQp8MI77TYV18Oo33/tyCS64qmkdIt38ZImQtV2
DoWvH7kXF1weF4fuFD356v8qfeZsTqcytWFmtqqOP/NG4ObEAe2ROCMhwXUVwwI2
q5AalHga9sOXeKhkfPM6Y7I/R5reAT5/0adHTRPWgwdS/jRdqDOJ1WsznW+M1wq+
HUMTPyIOtTn7L1EYkVjkzwM8eoIXnlQzAgECXeaniW4QCYc9zIzSMtG2XXTGM0jz
uJ5J6l716kgYdNP8FBHgDIcJRElz4ART9G+Xye0k0qPJw+wBm6P1AIfCL3kDxJeR
m+VFvcKlavzodmB944izNRBXRagnse4WJM8pdl37w+SV9FVhvLqNXYLcFFIIFEIj
aTXfjAivTUTQbV0aLOvsJbhGQMKZWmW8UkCrxZRguppb7DLKD5UrRbUMMGEQ6ZZK
vnq6qyNy1CARNXT/E52QwjqCK7lxPwj9/WLImjk26SAoAeuscaBe6t0fbyme+o5d
K54V1Terw+ClLMWvSPDZD61mUMQ54YpoXH51XnE2hPAOGjUHdgVxPVSkepCyk3xf
LDPEnddLoeh8mf4f3VDXM1KeeITuqWNwwnsHpHFw3JQYpZtB7AjX8u/Pmqqs56/H
147EJNOvcysga7sZXlGJQ6C1Z5hfRcmc3roQf89csEg4h7bClds5Ig2hNvq1AvMc
a074axkDlSeoGq56nbZ37PfMobUcpW66fUzjbSllrraYKnWHSmwyR/ehAGVaIROA
oQcMGxd6a95JvJ4FNZPZ05YjZW4QgAaEMC6+GA9++3ZkJ7+AvK+ZrwdZipFHu1XF
tLNvFOEZIxzvKdMn8boE/6K+6mJdGs0GVA1qn1gM81GY6uMhud+rAHeaoat1h7LG
wS2qDsjSIIavsbZv+jH3ZSL0W41uZLdbfoe6WK0gEQLzP07gmSildrnEDGbHCgBs
5aOH6iIk4AT8FGvTgPk+YIIgcVmbN/lIN6eFMY3U0BxwUDbMqclr34DHOyFbz7R1
V8ikZxxZs3JfUnmP6VQY+dic7OimI1NVraQJzeWKDfL9EQJcCnZg8fuofU1sxGfP
uCwBRKnilMomvgFk1TCA5Q4XuR5EBQXbSzV9K0tc4acd+yFGPyAW1+Udf5bkYAB/
4UGoedZyX126oIIperwvFOTiEzuCYKhvnKf83sAXdOGnA5UFr4GhSbh86xMPXk3P
9EPztDkQuH4+l0un47JaZEyYB4noCAZen5nBnsEApInh9OY3uXBHh5B2Xjd08fZk
PDajK+tN3lCsejn02hgt5Q54xE2YnvDpwIJfph3zOI16c5zIMdy3yDRRrhxkLv39
+CkMT7L83DsFXAc1XbmneKI4/zaHlguJThkDsnBLUGT6jCeh0p3FihrdYYP2lj9y
l0PT0RkkjaUh91+Yi11Cm3JFXWvnTg9+vY8hQOqT6wGVcq1JcCoXb3rm1L35BJ9v
xy/MQ/jqZ5bF7mm1MTCo+a0milY+Bd2h+ELFgSUvypE0UAvtyoEwD0XZUQamWhG/
PDhg+pq7WdyZEJ6ckYhP+oe2hyhTAkJIt6jFRfW7H9/tEMqO4I+Hg7Vz9uFiZ++T
WCSZBZZnLaptwBNn0C8v2SPWOo2+O/24jOJoP63zxVKUOZWW7Y1t1i16fv3PJFrs
34f9H/SbWLZYToEBTmfkEf2s3zteGWALVtwhvow4coCcMUeWu3A4S0JdVl9oY1CD
51FK77eqUFdfN9ZcJzGUtDWmlB2tq/6HLJ9UUzKBBBjjC1xkIQizW0N6oNVXlkGq
YfS4hHtjJZVSpNtHT8Pmah63nW0gvoNwOri5UPu7J7Z9669gB/O4Gpxwn+Ciivvv
dZkhanuO5N+0b+qNkyL6016tHZmjz1x3Q9tgVjXYI7zla78e3h+dBMKJSTNmCrwV
U5b2zczVgZ+JbVv6am5BY29cpbUPE7IgRZF/vv9M1+QHfThizZPXkuuJKgV64UIf
zxgRDpfEHJ+hlwvv8t4qNy0IKjLl4XiEXbW+fRX9HDh0QfCHpDggIQmoKg1mfHKf
+mxzszmk02FOp+664soOpi4LIJr/CvBxtir8KCJ+5enLAD48sAZP0wPFbi3qHlhB
AC/Y6+Bh3d8sw3nj5WBaKGwulsgYUI2XAXOIsiX8iRNq3yl9HnkJ/PXtgWSYB93g
zCY0SzzDVrKH1agFBgSI6aaleuBmVopfWjwXGCvS+uJOTmNO9fcJzXR8q+n2Ur5I
OxUaQXZ96g3El7rGU+rR73L+q3kQv/fEGlaJlgR00HpceY7bwYA7pR37TtIYU5cU
IPjOp5iv/Wvi67jwZLH9ydY2Pw3EP9sKCjtdT5YpEnu6040pjCQATg3BXPb5InoL
C3NVAwrlp/Uc3Z8vtrcrqRPHMDxwM8pPVS8n4vKbQbTQlP2ngY70wH6h3WQ/kMQk
Mist0ETxvv5la2OqbS3jH3IxhVk31Vz8zvGH8KSSJunaOrodmVF5BLiGrO5SLN4x
WOmjfz740QvsajHyjR7pOLbhL1zeRd7ImU/8pNwK4XC+xhkhJNFIundZIXCCszIP
uvBdGiNeZ0VK3GNHVGUNkel5A/TyZLlEI7/FTF5pZQYa6pVoqaHEWOOIgMaAZca0
omgR5sbflxtE2N2zdZBNzH4pq49b+XIRv1+A59NFnGiBKV3MUiWcq4O1eOWxI/7v
fCJfM7HyDLmQh9GsAIi1w64Y7rAiq9qYMmj4BzzEDOCWA5ixfrw2OmEuvN7IKM/s
PI+SRyUYSSxwctDagSOINVjKCqmSKPyhdMFxLM6K7LxTlizxApS22NI9XsvTymBw
/5bRjxhXDAkxD6gUON1zexb2poTyEfEWV1crmnvPk8brfq+/H0nLJztwNDG7ocpH
PKUqxRYHLHhAwpIIBRVjyrfg2pfoxioObKOqfSW2B6BLs0qxl/TIxP9eMvTn20uf
iAEaijlU5yBoB5iPcT4NoGJQeLPeZmknPR0JqTQUB+KVNvI1QKwgmrx65C7Xe+m+
8e7za3NVbikA/eP/urStCleAk/hk5CC850Sxe0M7yC0A0F2TdSnSLLheUMhKyDII
eWQsY58mWWELxX2pxCAkUFuRsqdIIVniBMRyq0JsR3sHXXIyJCXGKnL3O8htY8j2
QOaIBD+Fj2/TWpI5JeTIb6A4PR6TrnxGIaDFFm/txmDVQO0bzhGOYwnBY5njtKZW
fCDQuNwW+thvIc+oosb4VkcWkRwaIbPdHMT9jsT4HKk3JphDyuJ90BvarrebllTa
e21TL97WJHK9Y0WsBRuRKiATmYjzGNqwUonR8r3VjaRGnc/kRkIJCGuGR5Q5/o3F
AbWdCAYXstoUqO2EMY+D0KmKsgDIgzEg9rwZk//tG1YQvdY5B6edW/74ZRLcIEEq
vjxcWP30eToxf76qd5C4DOfrVWgbOmHwHwXVdpONTYW5Witmqe7QfDEESDHy0Bbz
brwMpKb94UwfLe1Ioy6/m9PY3E55BIqEvhe3q1Cl73R6fio6175YxFcv6kS7YAua
37HENEozj3a4dFhH3cDS6Qq1Z/iWcCKp6r0b3ciO2JS8fUqZqhHgLN3Izl/O1zv/
mAHLNBAuuWE6lMB/EJGDhyZ4m8ZrXgTkx11hbIM+otNM3MAehHAv10ujwagBr+zW
iAUQwx1PCfwHrTPu8O82mQh5o3Ol/bkylMaBGCgspSXxUaXGP3/IxUnHA4WlhncQ
HBDzRKcFafNud6FPlVo5iOJmXLGBhN3kCg9/gzCzJavPzLj3pcsUWhDZDVdwO/n6
e3vtTR8BIob0S88osNiRe9EFWe6iwSKltdLpDJuI1x4iocWZJ9VpCm5kZrQdbqIk
ZaXTMrUZVBffLk66TmETnFYLoZsgeQrbh9kpuxFMHSFvXYr2pVwZbWRfdAkusMLf
6RKiN4JdM1HrakcpN3DuMssF64dHPidJ9Fi8vnc9MCi2HHQ4nDCO4iexsvEvGvjr
6AVBKrrBjqS1g9es2LN/hI4dx8H8IAZvUY5tOnGLeeHjkRvKmIvtRDe1YV79+XPv
jnLolZ+21cNmpHzi/BGD/8fBM06HYvIK/syxEcXVmrKG4MCg3s4krVDkteZa+dhY
XhTs8kWB84erYVJ6DMLvLrFK+fSizdTXl577+y5B1npvCxX7hEzF84q3D8aIZMtQ
20Q0T9cUgABjfx39Nt+tPjrDmsRjB4FhvNyZZ63ZGWarIHiY0vONvSX2HFhBX650
jlpf3Ixy8ESzyoQBKaQ5P/H5p7pcvvbQs2FLrG3lWwQfMjGj7FeGYaPwVXgLUm5W
jI5tEWRluGsmoXiD5lLxvs9G19No1PcyTmIMiWM4PJk+ZJ3G7UzHcJ43J/VN5hKJ
8rRxtGviFaQ28kIPWFjLkErkfxrglSrBj6eZpw5+tuCOULWhTmlfsv55pcloEBMt
vatue371H5kIEZj/S/DwyWjDLBCWA86ZkJBOkErn9F4OZsdEDzMh29WvkmcDefsj
sRdQ4qEE+GrwKwICMNeUcf9j3cUWz5igs0j9St3TIHpAbAU+Y0YamitV9jJ4e4b+
iMSEm/CYQj7n41KPQvUNU62HPXNji7QaoHnAbJ1XmcIpb73i1y9Z+hMq/L5cJfFg
Ju00jLziJdgBw+CcRcslHwoQMHHQDNb1ctigKcncaJXaeOjF7lwaoxd34iU+qw1t
iLgXOBDceynFiPCueueap7GYikdxZWUvxvl6mQMlc0MRAoMn7RD/yecv6y3XlWCo
k1vxfevmK4+Re6zqs8ucut0VABJl0abOzubiSeIRL5AzpANIKrlz7GJCDbWdkHku
kC00Ky9G4VkAE6ou9GNePtieu+CoCBW2D3dy37QdhqjDBSjZjp1AsHiPWCXUOF4B
+OSACxYv2vVRkM4ImKqTAUJFL29Pg0CpzS/+0xvq28u+Vf5hpwnkH1GardQx3ZLg
/eH/MZy3+pnSKzeNTqxR06vDishG0flhjZJPxhFpadkfL8k8NPMVhoM7zGkc56OZ
GTZiFKbkqz1nDrKSraocDMbhQle821YSK0om0qQE3T8zhZlkw6zTToTptcKAySKY
G8vnOp/Gtmv6EcaEQYLOdYfPyFHek7UWIK1umSiv5XpTPpusJs82bbOLBwwyJ73j
q6tLQBQO7W1i3M6LKMDO/lkj5jGSZZ/Nzr999o1Ol31v2Ihrr/NqhPjakvvlgnL2
5IEUU5qUjm783oDmX20Cm/JFVNLP1lmqMIiHo7AKY+ERL7Y751Y1GBRiVpaBKa52
mbkIUp48FNAusvNoD+cJcwjJVlzFYJ83VPV6QttYP3LSdvgZzlcSqP0zLFR7NggA
EwYcDJ/sXDtsPrjFiPcAstLAnFvMtoXazHvvExws3x+dF1FEkWx1cN5U5VKMmRbf
Z0zkmpEI0YEJcZyVsAzzGIcIp5ocnGzxcYi0of5Ao7euAjFB4lUXOOQWjnHt72LD
ZL1BSUMYeYMrHtY9YPkLGxDIFAauU/4SrvIpREv5U5L5wLsRqmIz3a+qwNMfAAjl
sDOvVuhs5Wq0hXTbHc3kajXEwtYSDUkVThqBdsqmqGbtaEy5nLilX0T+RquHpV3k
VhEMpCJzMnyyX4TbdcImg5q0/M8n4Hmd8xWzC/KqLQU0ugoGJ3CLSQQyVGhORAKM
3Kop+E4Li0fmLC0UglYapZvLheFKwe5zDPyJEwK/WYp97KV2cRThxNZetJYvI+SC
vzLe0Z3KXtj+eqpy891SchOzGfUavk/2TJDdXfMipxUqZfENsCIzJE+LChMwzODq
oQJXNkQAspXAVph3kVg5adY7Dxf79lBhCLvw2hyx2k8cxnnol2qxZngjdB/Pu08+
kmzypiaJ+XT0y6mFRDkqCu2Dp7RPlWzdZhBZwf3QMhQLDy0NlSUGYX1UBvEBHUxa
E0mhSNkYKt4Zw+a+O0fMAGMTzYZE42FPPz2nO/27Vk0+a8EndS8VN5GUi+aivlXq
s7hlTSixhmTRr46ZI7w5htMppGlpIdElUnbVJ/kdrJ9nxzJL7pQ/iEJGj9LW3i1v
tG7TTb0H9baE8aly+DZX611IGaAEVzgwuBGYsCFrF4SFRdRz4EH8X8IcGhUHTLUA
bYpzZnPi4rgPd/t3DeNlZvfBfg2D+TzrEVsT+1KRhafrI+rngEGnxAUsZYOeYXkx
TfOL6b/cYdY7mT8wsWkBwrjJs+mpVVdwFi5NrFe9KVCa6myFpsrKrvTE/4p7/4Jy
Mq/1HgAgD7dA4JNA3WJIdyWB8VFrkTWntA//QA+GOa1Xm/xQFXZn8oe8cFoNCzke
KcRaVA3bryZO/rmXZqM2bZXTvCh/YFA6h/m2/pppqgEChBqFokh4ssndppG2ssDm
AXI8MTVIrfjQjG1TwWepYFukem8P/gL/33y0Lthb51zJ6eTY9n6GVwfraFhz3G7W
XqbFnBgcZNm8zUtECFSp7m8bDxYE5xb5nPzJZ+slDyvc+lN3cT5mE9Ut9UumZuKj
KJotdBbsL3y6xaVLyEj4g84XwZk5ISVMraoMwiuXIWuH6UoEyOJXmWogjBT79m3H
Y0qUc5SaFk5hcL8o0WR5qER2XVnN7l5/i4sFH+m75Uw+7IjgdSXDfkEMrIydX/7F
LYznjuZhggCUew8mCQ34v4mJca7E3cQjUQHeATvGWXOzbUZJU7o7ch/PHn5L970g
OL5QuGvI3Sw9rqR9/Zd2c7EWPeOblvO5Tv/vqKhlkY+Y6uuTUhgnnYSu9w/+/WsM
T1e4LNiN5QXTD3MDHVhwKNR/wy5QXDWLKcm4MK3oVcPHVD7aq4H0FGLkOoDFZP0Z
q2kU3By+ZyqxcQBo0xm4wZAvwY8oCeV5Q/12JXfbfebBgot9gen0iF6bReVoU8je
Zhiv6Q87RKMZBEzPlvo6FhoPy0p4J1nPM+49i4DWfMTm0v6ZnVLKTZXuheqd7m3q
03S1wKqLIBMPuCQaEGvHm8wbHCD2K4Zp3TaZfoBUC9tKBmcwcEkQaodYCSXWBnGO
PHKRIYnqbDASCncofgPyBgP9c0PffVZIebEF7RqQ55p4RMRZCo0Im5Rp+nCft/fb
R5IdC5FWR4iFt5N2k9+zXmaDBHEQ1NE8ErtPTgy2hGk9ZzO+I4rAzolj3uxaYYiR
/UZhtCTPilJZBF/GkSoya+7DKVmmu/In2uLi6f0HQUv5QyUVLXNUsmaU4bV1CEE5
gLGOBqJJ2cckazkE6jis5N3jttkBQyiyr8Y3BaIOXZYNFhgofKKD2OM33bIOUsHv
Isp8EErU8LDHLYKqSETrEsmjylmwXwfwkss66E6FhFQq0KuYE8Uy/AdBSPff+SFO
uer5GyvgrJH5klbxiMhRi5t0nPCMx99BEbLZ1GsgBtV+sfGugeMAamMZjXmRexKq
+adUdjmDYUY9WXNGORTE4WPsaMQMUuAoE/ladXQpzAZbmaC9Kva/k6UiTC1k6piD
rMgO4uECwwwS7Cz5OR7AEgUiDtBbklCLoKnhIN6b602GAaIbIaCQikMrpWtODKa6
5LWT6v2a4ORTJthoy+UrvqA5CX0NRIoc3hrDaEMjE8ohTMO+t7+t1Y8OYXrzjsjX
QkX0pqGs6/JNgIpWeXHCqCBaPFfKWX5HjbFEcv3OGD8niJ40+gtAeUWnzlVyqFAs
7Cy9rnEncdIiTToNq6FbdJJ5dxTrCwT0zEoRdTH9RFb/13EosHifeqNKONlJWOiA
rSPhDrvt496nJde/yZD7acrmNrQFlqbrHwdZ8pOoxpVN8ldMkOGjR4lWCxSv8v3u
65opfroVs6gBrkIc2hmOrZQ7eY73AlBMhi6pnSDD4qTD6NUksRGkasLR/EF+HbO8
wANb825/vT3H0/euhcZnORUxJTBcHi8n7S1wDdNe7xnbhKLwl3TEYKHEjEjiXJ1d
yvE2k3pPALw5JjA/1xnu8tvb1bdvDex80iEz9m+9xfmf6pVu43U2ihML/OLampFg
ps1cfsZHPrz7z2L9Em9FbTFLYoQ276QkCx/IIvqu8l2lrENcib7zVKpG3QZWSkcp
uobG7pH9mWN+diUo1fEf/0CXfWWwj6pRNDR/ChTOT717jiGYcM+Iftp5bfdHYXLs
tEJJ8c0ameA0xbbc8F+g4J69QfIXGjAYi0OH+0W7L9/cDeqW/lvVi0fklJabt74w
+Q9nVOm9qfFwTpFJxDKdLq7Tg7vloHGRDwrED5bWPRvti560knUUOXIfsbB1OySf
4iZbd8IjGZP4T0dQwGcA4xKg3vcmV10e+lPH6hQrFRUa1diJT7C4xh6NbPaputWd
0CQLq/3IXw97W8H7BhhduY1bLjteca3J7lqYKkgYl4Xg9rDs7HYdq2P+svTb1mSk
U2eu8lbomge8v4DpvjFrAZsIMzSwaQLNwjuzBJ/+OaluNagHhyUUtNFX2cCjKW0B
i3RkMcblomqxgFhE3V2NCUfnizl5WpAzd2jqxx+cbuePRY39JU5j2ohwCc8iZv0C
x2nd5VsvT3TmpDKg2P+KY38Ft/HYWgWhUxQla1WsMAQdj3kF1HRsAgJyMvIbhJb0
CmYrLY5km2/zgHsQJJPjH+NMB0DTaauiH0z+YLUatKGjOGTxg1eq451HwsUgv79s
NRh5f+nYFT8mTXXZzrAYsH7VFlfx661Z1E6V1e+SfGr0CAIBf7Wcm9ZuJZxK/BMr
G0BkJdsgAI2HaaYKWm+n8gUrm2kNx9lmUI4WpIuNv1FzMzHp9btWQwESgjilArEE
7a0e5GQbXo/PWbfmtDgGffi4JlcGxuLwzEvQszzcsQohd+Qa9V2xfpemPYP6zhG3
DRy9te4+tbPL2bMflU+j70t4X0GPKQWPNAzsj6Ox5MaK41+MVqYrz1xqu8vbzO2A
pLJl0JHdW2j3czqN8UZ9+Z/fhxBFzAPRANUQ6qSi7rynfJUVKrexy2qj2XgLGxlg
QlwvGxS0FGBmoi/TLsc8u6F50Mq7NPpLwLR4r1HzCGqVv5504Ji6Di8/eNGAAuVC
GnjUrBz91JL9BCdaay26p7Rq77f9VSLg+LTwwXUm5+wfhW2DCb4AS9zVN0g9pqEC
L/f2LhoCHd5nnKom++defsXAFGBqUMQcfAz3sZA2IK4DTZC95rUscEQowY0lyQqB
Rcy62RwQ38TKo/hTlIFvcfqxfk7RKTJcv60D9oWzDObQnRcKYlH6kWBqzni/a68n
IEBadZ3xd+W7D2YXlUtxDJD44839hToeX5wIoOeGOloAjflWgn0ZRfxXx/siHBtS
eWd+hqnEwRty1Ph6MMqzB/0saM6oktNgJqaBjDDcbQr8jq18ZkiBmFWPRDcfIgFv
I510YJyXzz17H/MM11cjc/fr3vSbkPS2axZtBYxHcJCAMEH9NHnznqNqr/6izsNA
EYeAoQl1Tm2SyQMejAFaRhwP4VnuP99PtQ/xSCDRCnsuDfPNAE/jDX/RTCpFUMes
APHrYxsRxeTUpiK8biy4Krsfn0mkNfLLMTLQxDU/qgW1rFV7giu/eQmP+hn99dhg
fwxrZ9eWAa2LYYRK2kIThBQjG/zWgp7mypNwzVevCdVlWK/8Tzh325x+/xw8HvAA
+luKlGHSZCbafDRI+L2ZrKHEM+HZkTt6avw1h7Hc6GxNvLThPfpMCXSoDsENCyTn
9bFxTSVDJ0XOPSD3M93qeQjm0lSZZVWoDJ62uTTMAUTDWRYZ0MiP0D6EQj6AQ5do
zeS+egTo15SHqYhVSB/0l9Q/f2OJSYty+R9Hf74BR5zhlOqwuppTBIv8LBsEJ24c
FHtCTCgNZYlUgKGhaobUhOniEWSHSWgkuphZ92DyHcfqbr6rK6Wa5ooV0MVwwkH5
iCPp8D6rdVt3gaptOUxFRLQ/ZUk7UIx+JWigakbvFlp3bX77eBfg/7M/1I20Jc/r
9lLWaGLeEEU4u+uGK7vAbiZLhXzTlLuwbRD0V5gxoqGEidS7XxVlbwCfg/yfbg4G
cxE0oD39oWOgTxFD2K0GK2k+gONytX+qbOS6j+ohDEzQKYILEXZIiLpjyFVsgjn5
SVKV9qFm9TN3KrmrgcQFMsWAeU6Hi4aFtg6NAjQ80mhSQLkXCsB0R/misUOciWkC
3otMD7DwrZOvGTjzOqPBC6wILv6limHgOvaxR7MVoI+NydX/+DTtyzldBSc0e33o
NSUT2PP/5Fz3Sh9BC21m1FDXcGpzVExf+bjWLwy1jtad/5MXgxJ+VuBobmREl2PM
/NjbnLhtS/3pT4E832QFL4esBRmZn18ZRGB/SdYfExL8d5AvdideM50mtDLGTiHf
jhZu794dy7j4Z2p7Dfqx2RP9HzIO60lDgUor46If2nzlA5XgV41N87PmAUlQiGO5
65cIsdkxlib4NaCZsb2Pxm95zmV6jYyIbJyyWV/BmkFZ6OTP0yES64bsXXdjWJKW
jDFf780OblGDGN+R/3p+h275BKqvVSbTvuNx/SV+7McvNHxgH0NHJtUn+tYLmr3e
I3fvE1By5Um5iWVMAc1XX028UOPCXwoOUr3xmYhp3LNmuaNOgEuwX9FJgarDAPym
9LfLv5U+WGd5cwsPrPjEb/E10PrYX8QyiZczQbIixwl5o5jo4MWbCj/s1x9RWlXb
p7uWBENwc1fG/c/7S8kc+xl+CwcnRk9IfNMyrciQqFZtH655sd0dqgdSWTi5JdoT
z13+5qlZZUZ2cj+dEK49ZpzCIlriud9u1zsbgIDk/hICYiiPSHIdrDUyvNKhUbyb
Pe87upWv3KKQszUsvB/WmYNTuK9K6+ls53zfgS2lUhZhZ0/pJXTzArC/e/L3Oy0k
YhcfcsElwKeNA+Ev/nZocXkAVvj2xPlH0TPeNgsWJ3HFwpUYq5A2Yyhzqn/AutCx
TNsFFrT033FvfrNrxPD9gP+T3RZttvXSYAlUiVs7fxR33gSpFyzK4MS296UQ5HVC
HOcxVBNAzozRp93AehtoT4523o9kyOJWpMzAv0nqTJspMw9qIlIZPCeOWvWVwQMl
OTpnh/tQwMsBIETGqce1yLQoJuRIuvmN9nwDu5Orz3s2YXPx1jXe2HcGfj9gaB0d
1oVCpX7tl1TRHnNxno/38oqmVair0nLmd3IxsyCqu+F9RsRq0rjGQikxIwcso5QC
ZGcDLe4H5L4wPLO4AD8uIHIVr5J+9kkJ/FWA/ZkNLdwjXQM2f3JXTzAqA9AsFPC/
bty8Peg2Qn9bCJQ/wEcYi+CnwLsmuFt21CfvA3eT9oRcsm/LGc+VFtrI3+51gIOR
d3TkS1bG/KakPfUz6E9sNwSSvvg3nYIN4QkdQg7ftQiuItygjIe8Dgrk4vquVHVZ
07GS7vvC9rWCWe3PeRyelyjs6KITMwjotOukNnWMZVJugl6q+wp3XCyUySKTlnCk
4a9xFCNAscXhEJX9CZEr/q+JjbELXOSf9rKwCF0/WvtZffDVYQ0JB8pUUDHaXb1F
E/EC1FujB/kCH+t4L7N1rCJYu2S2pgE1qYIrn+YjmlU=
`pragma protect end_protected
