// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XMVK2kAFI4T4AMW/kS8cJFFvYXffHa7e6oS5ok90kCtbXXL2YjLhI0YZdLWb8p6/
G+f8xi2mkM/Xcq66sIDD7yvJjrgV0oYRJ1cMoFJnL1OYxwWwQFASslHFKsLuw1XR
9wH+0nTndLoK0FsGMpPDgpZZc7hEWsWdU45bjmgTnkI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7472)
/DuWF7FzW8YPcEcFnKfpyrRkSLBQIZ7qgldYJ1ymUEntLg6156SFlLJqNLqRkWYl
7HrKkmyKokUiF4WKMx8tcqLLgXS5p5i38zuxNVzKyTtTKmw0xiWUVeK69gDZ1pXR
ETM5aw0U3zkDL4ZpHPlhY10ZloHXe0mwODEf1S8769hTJlxq78HP2E7YymrDECzM
17E84tuYNabCBGB5uTQ7AX6rygWkDaJ/1HNggD4Xi3oAeoi4IEoCThb+PGORoe6a
mQZgov2pI+cim35gWEekbcFPgeqBmWngLOnLQPRt7lkhe9Oje1vno9VqCBjd86Bb
tICwiW8ZzxiqzGQ4trHHSe1uRds19QvsLuLHFm3QHNBokPwKKlrbwSEyYm/W+u1z
lTwdP36SoiCXns3i46E36J9MaBBmc+6TFX3Y0siNVuRkFCtEk3HWb/H3stIiZsAY
u182CSglnowPFCdXapmynsPt0v6u7Yz1U8cihInBhkAwrdO0wUVohxLaR1rqEXP6
sxvAti3DXj9tspSzRlMvWuvfvdlYLjfdtZRDxhqsTneVousCHAhQzhlNfBDD6AiY
dPMz9u4IiHbbk0YVsBbNPLgnB+BaFupfDuGAUiZNZ0yjP4PBJ/5vo+p5EHJMzmcx
PGeVQ0tX4uc4OdTOVe3/LOWhVwB8vxC/5FO5JxCJuAj6LUku8Pgw5611IWagXDmk
kZN1N3GuxP9m85AWL18QlNke+K8BDro9sfclqdjzjgyzj00Q5rwHF5J/4uu0sVLy
HqS0OBaRDs5w9LxY5hCwGQeCiirQFvzNe5cc90mjkyLV6JcC8AEglDHktpMsvSUo
Uu+pD8lTTkVPeV0t1iBaEEAmkYRqOwO3uRZW8ywU+e44QsYqb1SxCldgFAOhX4N1
jrBTSOlIIU/SULmf8scYLpbFO1XnHUIbh15jgHEfuauskVe4ypgyXaOKHqOOwIDn
q77bcLB0XY9gVvFW2uCHNTxhi3KvV4GrBuetECWDsOQzKcBMXj4ISs6Nx7dl1nrs
OyQCln+qpWfvD7UsVi/yXzqh0KGsrpJqAGYuXN+SernsVG7kpO6XeW5bA18L7rYr
typXVin224mA+vJOy6MdWI1NS/szTwLkYx1Z85UzOUlnaIQJ/gVKcfR3WAx9QtpB
9rjMxy3H5SaylgF7959FG4mjW48V+2Aa5rxs1dSO3WU93IqpTI+flCsrCvK1XNdQ
k2wzhAs8WbaBEz8gz7l85JrF5ey/sN8M1jX5UkMvRc1vw+u2S66PYDrGvLeGmYzW
cUjP3jRQv8Nf8n5ZRm5aiKNlF0KLzWusN/+B6gmQM7uSoehD+Q37ciiCAxFmrB+S
hLgyM0LYeeUG33AwT0Bfl+pcPlPEkh8xXqdY0Q5lCKiqePn1p9irxJh9ftcqsKaz
/InXmDrbPqHJmdVqNHkUeDxU/Jt6pxFEFYoRJZBzD3mQALsKZ4ZMzcrb1q5Tq4qd
h+dVDoJ3TVmj40bYr/5Tu7vrspUzXxQj4zfIa8zbzIjnb2lYaSxSYjYepnwVu29N
KbstW7+6cr6ViaB+AgL2e31q20STIdKIMUDCIxk/64+RccwworZqkP+EqHETXY5K
ULX9FJaeZ2XxvQhJpWa2k6t6ZOlm193UZCP86KQw38en0WL1bO9MKXLhA5oSqCyf
11Bpqwy9+m+Vim1S7Ms2234jQ6LDwy5Q5TWf7wknPgk1+qXrVS4jWpMoigEpHtKV
H5AhOsGK1WxPJs4JcslZ2cO++/tzIckwy5NB6oTIqTp8NBWElKH2fZx/jq/VpMkp
eBZhoGxt4BcRXYoTEbuWFG8h4XcutkK1rQIR2U2HadWgXBQZ1jZ2TGZ0eYOX9PLJ
+of2kffKEV8mdz1fS8bDTGTbUA8Ff17EoOktnjxymFcZNPuVccPEvg8c9OaezmQE
C1GqtZo5on93hVFihxKU3xEI4ZaxtSYQGSBRAfwh+3kGLfnzTAHQbrJ2Y6KpmDhZ
3bXAZLdjzrdHZvkSyl8LdxAcHPcvCGh3ivJ6ovtlQUoDKy78tGFb3johD1qOmPZt
N9jaRS0hK7toin8QG5H/rfEv4uSK5qmDqVny2HVPuo4kPSpHB/+bzfqdOIARh0gH
HUBNyKq2VGvudFoqGQFeVg0FJhcjpXmv/GL66AR502lZDJKDgMvVRRAdMc1imq8t
dgnR3vEU2+7K4eFm9c8Y1/y8llPr46AZf2jWczQKbCFtjGP+3XVWLKGt154FZQr8
C11jmMKFkNbxoF6qP1RRlqKwSs3eMow/nquXC94HH7kIRuq5cQhPLUioH3Xit6kM
MIOCDh8T5+Chky0+AoGAvUl9c3aBDEOjtjf7CVdB6aLCVr3h3a2WEwS99iIutom/
TB4tgms4aTHtI2ZIz9mCpWKtF4NAoS79zwO8k6NZkHPOzSgye6VAWU3OFV6mGj0v
7nOkNwxku5jH4V6t812KGoBSQzlTQUE7/N1LIg3XcorzgqhvqcUxtWwohEHKlNdl
uOhCIs1XbiCoi/0LSWaOOsi5o+eqBtA72T3L2AuP7EusrEQBZDoLxh9U6s7olg3z
hFW5lfuwh/VCo2e5TvFHJ/izEQ9dCbTPYLK8ovw/RDBVQbYFmQ9WmO9P8YdI0PKV
igs1vhX9X88Ic1t+jY58Lp4Nf7lahV2GppAfD3zmpsvEwehNQOWF+KwGu7YY3cRi
q5TQOtN0mikAGmbsBQ1klYIfqgJndE1QGPZ/jAo9f3zRkB78HSUQ9aWfDZKzQYHu
8rQ3E7iGwOIvfHoDttNnM9VV55ChN2wwifMKNFIxHs8gEsZOPYe/403HLelRI9pR
FMUXkuH9/DAQ1cT4OL2n/UY/tX78o5ChvFwdqBO/A11kV1WQkAp5k4yePu+a2MlQ
WhMUDkasB6p8eZblhVhIg3TJV2KlOaFWsFWZtNXlSHTk96ZRemkJhreyNG1FpLTh
lewS8AzWy8ZzjgECHOplcaGmmPpp5g7D248VlTtf8udGfmuU8zVw9x57CgmKAz0U
kGlzm19n+RQ5hDXBE1wQNo7hloVbZZHsrEKAcQGnob331hcPuGJVuStvj81IrfQP
w1S93nPel2r7/8kgUg0lyu/QM1uNLGAOOrUwMS/SGuFMsKyTqWVK5djOUTlQHLLu
n0DCflHZ7/YEx4LoR24+rkLcasD12Kj90XhYqWbmGz+gQbzSi8/AJiOTEU/QXytN
yZJBoP8Ls0SxYFCVf4gfi9JeOxw02LGOFAIDa25b91FpYkcfOhndni4sbIf4nHfa
uNfg8LZfSQquBb5py1p92lhiBoNkj1LgmXPLZZDZ6VIuWP9fd2oA0gWLlUuDvsv4
3h1s/DC/2xuurEijl3QSqEmDxYPBFXjFJQpznvnC2kttjmribwh9cLkJA3y+9rlL
CerN1cmG6H8LvVIZRtTNpfkcphgXixaN3N/RYVrM8C53Oq3wkiGgOHt/4+BYL6wm
sQDHJKfXik8ncUDOeDBNy6UUUtyApLaP405jki33BvAAQj2OqIH6Te3HOjWWCYpo
H8wA2zmKfpwCib8iqu2VzjftneKZOZTtESJnoNYtbUIsdKkqO+tSrriXR6q8wL9r
0V0gViaaaHa88/Gr/8wUPwwzgmiJUHMPbFgz3kz1LBoVnvk+6LGVnQJva1u5gKc/
XrciXGPQEOlijDcUQpXhNx6ukjkBgOBenzr/OFAs9wbkhsfzmI1zxaicH1G7ci+s
u13bIccrn7re6cOXaRfrglvLmclHRw/6DREyt+ouMTTO8+h8UBLjl+UReH/nM4N+
PjVZZdlHMEXRk8gJ/xPWSLVuGGv3KtKjOlBiPojLLNuUjnVu4RFGjYkJnZM327Qk
JdPBWL+qzD6XAkNm37TC0usSHMuB9fzQmydYbNJrwzb4Cyoev9t3kSpaGi1burnx
vvCsi6AE6/sWFMLDtATfs4Grz2rLI54zPCvQrIQ/s8l9cy7PEGoSnmXFY7GVxMfs
PPjQb9qBZi3OvtTSQXTOyfRhwFpaEvA1jBwlKD0fhm6angpurRR7CBDzD4y1eWOL
t8livcTG1YYh4VmSrBGH6RkxZ+B/M3q2qSLZ7ovxZCGSYLhRBfXmynAozvTglDZl
nFsWu7vACgFS7FCZGG25288QuZvrE2Xb1wqappMgT6fcaJgqLNc3z5HRY2SU1nMb
SpPAywrc7GDAY8gW102bXF/417WzdcLZy7IhDG5qA4WVdTTra6fbRBUqlo4rIoyV
24m4X6EhsSHum/5ilmIe52hbKqdJB/DrFGB6DQjsnNhMA9RBimIdo1uwEkH89sXH
lx7cORpHb0VIFBRkkUtmLhM67uMAxXFB13JvG8cNOKb9Wp071m6sA9wMXGkAdiuH
G9TeRsb9EqPQ3rUxzEsOpUutWc6EYJ8l2h4JwSEVzb3VY4k8MO4Szju0uW3DVfx0
7MczWKPeiJkcQ6Whg/r7QUVIGIXEsg0yfA1IeZbvThcqrDNyoGATFH19Y5wyCLzS
4y/t//u6q2b8kJMVlwOsGiY+PKcFWxJlDFAiBrqaz33zzS51Y6292WrkO7XQ1/ON
TjEzD+E8TIbQ6ri7P11jB/9nZKK9ZkK1y3vdVeNHnvGRuMSDN9jfZx1CJF17kpgH
ONWCrPcTVqVAEYBwxFpfxGJ94tkZrn7+JE+cahcCChYGHTRfs/CUkmBbi8+ZKLib
MjuArSZY0wteaDPdv/4nA2AqIIqBSL0inBrLfCWxhqCZsfmKRuBc19iRzcE5IM34
eAfRFuCB6oz6M7jOHsSVwOemy35crpketrNaSzqm6/MlYv9GI0vzAhT1U9ZbqcY/
n/W0gZ3rWfi1oZDusch0icfV/TGb9u1o5dQSMaJj8C9DU96ERzSLYLHZwFdumDGC
UDFNKPoS4LuhNVLLNUTwYft2aJ4oyaB5vtsT1rlLa12+P+mnR6vQMk4mg6k6ItI9
rUNEuMwI8j/Kpx4IXuD5r+UuFGEHbJGfZEZTd4O79yqmQJXxeF0i1rkKFIZjdnz7
y4KE0rG7oWB7/oTPII57BhnWpzAIsbBGAcFdleI4XEFk5dt5M2B4049DcvcuQD5g
ZGKelZg7XvsECFWnKPlDeplWxcXmrNq4ufG60TnmFV6s1vufPsWCu5/Kl8cfu6Ez
9B+hIH/Rd8kj+kgIqFCjs5XTaPvKvVOhJ8JWpRXNONW6XaNAVhK/O/ZJOxzEfaMO
mRLsC6F2dObapSIqGmsX70GpglR+r1ZbMeVuIthd+b8mrummpkIt1xnORFBOUjYI
CumtC4JprsX+8Zg1OoFJUt4Oy7Hqe898m9xLkc0vtOcFlXk9UKbT3ZD60+s6qdGH
FmTB+bPSv7MHigJuSRee4pT6+h3raWwi7ygT91fZgndy5RBp6IzagQeZ0HO1sIRu
CyLg5d5VERteMP8/Dzi4eCbcD3snEd7hTrv61wAxEmQPOs7jN8lmpCktlqOOWvwy
oZ1uPBoesGaVWN8EIoZaQcJp7x/F27qZK7NRr/UZY7tKZFSFPNbbFoHx4DJwuSxR
Wzo8uxh0fa9ZBOqkxpWMo/D4xJ4Ghx9haJWTXmNYBFDVLE/ru+NrGaZA1OG+r8M3
xrRNOmZIkJM69SvZQ3ff+aAOZF5/xv6frm9Mb+cVfxJ2qty+6649cQBDxZaOQOT3
grq3LuKN2zTnfmix9ITtiwQ/QnAe4bHwFZk/FvHaBJQfuDomdqi+MPMW2iwWijsM
AoJ2ObSOQsCywx2ltTF9poiwomOHhRAJtHjs82uBUqS/CNEGLDCS7uDwxGhwRayl
w5jEWRexb922ErgSkNfJOClXYA2zLWWD4OX8A4T3DiwQv9ZYniPVLQ/fBGznPhu1
dmjmZ8XuaJRA6KBNud3JLohco/QZe4asKXaL4pZb4otwaD0Jv9IRkoNBkbXhzHxC
SjwdckWVbhp5bkodyFzu38Z7Pg/OqHpUaLDNCs4G12ohgGwKgp6KuRK/iqgnV83S
Bh2O1i2z0Z5zZFItTRZWY41KbqMR7KYwDg4MoTbRSgDjaxZCEeRsCLA/0R5XZpon
0hAQdNFISxnn/LDIGd60XIvgp1o+qea2VqgjHdLFQdZmoYIorylB8iy/WDVIzS+X
uX3kL5nrOHxa09YZHrkGYNRmy1PFf7aBYfeYyHsV6ANQTrR03JeA25b0EtWln7wb
xFtlFYam++sBUCO5tmgpGa4dz2Os8d/AYwvP6CyJQK2foxonNF9nsgDpSKTTpGq5
YAE9apLDB8YYdicAI211WvrFmOFQP47GXvBOm14lcRZuj9f/Nqg/FTVG8Z9HqwsD
J6odh6hPJDMBazlnqSox8GlVHV/wUD9A0g7qYkGsEqIzQXbXBdmZrt75TOqa0v6p
CTvdYyO6CdbPO+59ycU6V43HEIax7W+RV/+BTqCWGJBBTm/APsvZ1iqRFvp0/FMc
e5PYdBrNvhIcrNYx8SN62XxSELpJaCyIkCnSY3uUBvdTJf4WPz1Zpz493MbREuRr
6p2fm/vrcREkxVLa28qJphejbRF+imN0N8YS6MxDqoAZK3Z8teeyvvvK55wi0qU7
yCCDnXAqxzpb1Y9/j41zNUW/V8jFtZOp57b/W8MjPihoHcMbLJzxN2zrr2rv3wRm
pSiHmef3Sn7X7mL0SkTV/CU/nGQ2f0o7vQltfvvBLNHunNChNiToIRhFg5tLL1ag
9U/H2rF+oL8yRw0fTsBHeX1PTPbjRTSFEkxq9WO/9Td1lmfMrc0+DCqQBr9KZfNY
7P0ArFD9NulpDxRIt78wavZhFdf1PRTVijBsBQ3Z1w6+Id0bOnemNO6AP9EpDozy
E8CAW0QxIkkQ2RVumTuHIkA85glTJ+E+C1ScNX9REG3X/h4Y705gEs2Imp1CqkPZ
4FSHyTJh+xNWuj5ZKFcak08xETRDheV2E8CFYTX2sh6/QDnKGvqMlKFeVQBNlSqL
QxRySctsTvkz9VugWdZ7diryX5+SJZkVwAD6sSGMc6aQWBlc37OGHSjIhM91sBm9
i/tzi7+waVuLqYittK26DFpyL5hQO2X0rsRcggeveB9Tz94QtjAi4A43s8EEdX8I
VRoyut05hyEgZtqYY5WA6TcfhXlI7e+ng+ySUqG6I5VRmoAG2WTA4bDzugzyV7fK
wtdDybN25dSL+z95q6ImyoMsbdNrkeFDWZ+1pBHNHbtNkGiCUgDQnWr+SvVe8Orw
TEXntFK4ZUGXziGMw2cSW81XtIze7YFuJfP+z7Fama5r/NpxhYTlpv46fYy52vmt
t6ZNVYfLXGVrcVLWlRgegsgniXrNh0TubUENWj8TGxyxwtk6Cn8QPqued/TGKsUJ
PltuZ+1lSddK1OPmy2Ndwodo2jdY/oE0hBMG4/yWVkehrPAnFqOv1/B3f+sWUiOY
LsfvQYCS0zvtHUdNkYExu+yIY2pwxAF0SR0ZdNlQJWlvXZKO5uwt24h0XBXeowyb
hTkDCcA70tmaf1f4kVEOe0+iGMLNpoj6TvtJT4d1n5Nfj2fs6Bj++xqiip/ClQUA
9lQ8yXjFsYcfcdc+4oPaWlZLxJugry9Ll8hDrUswnH0W/pdS6F5zHL7PXTlTUDL7
mwUf7xN3B9WTvxTjvp6v0+aSLRkKr3wOJPLS4657SciYpcbMm47WzzoepWAnWYZi
1gZEiVbRIBArKtGmD4VMQ4RsDHantJ2s8ppfqhd/QLovn1VsfRhRjsW3fmQuWujO
n5rGQkIvTCMxmblvoLGZLiE9E/9IlZBrGOX67Y8n8euZOz+0w179zreFf2UJOwHV
HNSRqL5TOOpL4Y9kT91wMDHzXUfq8rDAhSUxmyzqSylg2bN/V6EdV0U3/qetPt3R
RSqRfRbU/fhmx+WAo1l9aaZp2oo9TBV4Fx1uV9fDmSKstU2N6VTKL2hZlOPN9E7J
tSp2MWlqU1ux0aEvmbT7Yh+QYFvQBGkwsnTPhAfTuGhaJIKuuCSMdI1hrulvp923
9++eWEcXI1sdOixohM8/DvkqVx2Gom6N8AFZzEJQprXzYHrQSoDh+fA52Uas9bYU
9yr6P0/El9jspjKyDS4iv67BHWALE+NyXsxF3H3HbzlYPpJt/5MTve4GrtNmOzTr
WFHnqSPpuFYI4r5ninWHiX7PHkre2/KwfWohHcQKA4Ha1Z6ehzsoLd1MtBxG38v/
x0wgdjs9I0Db0GRm5jS7UAaIvcpjKbUHHF3bD2olUEbfP2KYZXd0yiYq1jCqIG2V
x9OgcHXeHVhhbBol520BgXLVg0uQhm+G2Sxe0kn4EGe8eMSIMEUsUhFKpfdYi0WB
0q9whzUfm4yQQpas5QiIZ33yXVmmx6E8+VpRQHgkeuC2pJyIAiB7qcdolQW87NDu
flBk/urX3KS3rGKFfLyln6kW2vbn9EAxQvzJej7Jc8f560sF97ypniJsPupbyYTB
4JBApqIkEYmhNYvOagAVguh2vnw1fBlKpl0OkP1c8SGVlvhnrhaUTQHRd/A1ExD2
9ulVkc2KNdCgnM+bKh9BAPtqr28fjIW1npa6u/S/dujR4DVwZRaoy28wFzoHPPdq
sFwULSkIPVm0uaF8xli7ty7NHCMazrAFJ4KDrCYMvCRz2G+hqh7YXDF/S/NZv8E9
9gTw3YUF6MjuYyETMnqf4+OM6wUELhMunxzpc5gi18jU6Ek7WXTbV07meOyVNAq9
YZ5g80l+9YOamRb5ax/qaZ42w4Ck3ZBwpn9LA5QudrHQp98ysNnUSNlUa/zr2I2v
zSWB84xuBk1p/h72Ofo5J3B42xIR8DJ7wVSkODzyq5vOnVK/tuHa0J+eno/aOnWR
CfxLVDs3zL61ebeTfJP94mLWUf5F+epEaCeDhV1Br/B0LMYLmMGOZ5VonXtMo+fA
DVoJq16wkTJfHW2afOTpjcQxZZtb73Avs1D3gASYA/iroRwafN6tCF/fWSmQ9yXo
tCMMY+/vZMdC7qwAls2iZ2EluPjTgPV4NE6Rlhifbh1IHeS6/ARkuZgZ6D2Ciu1P
d0x3FFV1WQtqdDVsfPMSgirua7LvqBFIaaFENMJq3F9Zsz6Tg2J8q3cu/7bvSUN8
6+FiF/wG43h53xeDOHShRAVikteK4qowd/e5maxFZKOi6XGykpe3OU/uWam9NaGB
GKXjjdYESanoGaKCUffVCrLS8ruLhNgc90VOOH0RzJ4UPHJxZKW3hRMEETVAw/Jy
R/+8NOTOleStHYtK7LPU14EvP70DWAlgH+e0u9ksLcN/NbXc6kP9FC1CGs2eYcC7
/E0xbMbM36ms6LzxpOr5P1vVuCXdyu+ThXjRYGlZCDykOzTOSAVIDFDRyz5fjIYd
IJ4eAZ1ebquDHameqkBKigezvAzghwW2Lv7AYxZBDuZ9NkMM/eAe5bAUGwkdhJi0
Tk8K++5eiMKO7XXN9X7USDVs2mEDxQcW3PGEYkahYrN++xvx/GPDck9+lz59DH4F
2X1iWiTFOOla1ICLqemmmiIs61ssgScGMjk+s/SpPVwBYEpqGJVTnSlAj1y0ekkJ
85MmC7MK07uCyekR/9RR9PFg/fvN5DJkBS/pRagkrc4l/MTO5wPI6A8MhLQ4tzTk
74kuHsna2+iqlU1O/itVCfOEKtKxfoF5CvbUW4UmdUpYW4Lgcf5NBMnD4zB1VnTb
Th/tV4pfxaVadwdxXwcfbtygsk47SZmf1JiUCNnnjkzYoXQau6PG+oPiE1a/XOeQ
SKbDYcjMH052/WEqtoKV8nNVpy36FjwaIeOF7T3IlEbi329kDHY0UFhSoYRZFtvR
Q+JLTUFqxfh59X07QdsaNmSiB9kBNkoH1Gf9HJLL2t3KI+3Q0Y4vgFHgA6Zn93Ui
6A1UW6Pc/GfQfxexX17+JyYHbOt+MiiDHe+1GTrgdkihvlX4+t/YGDOqJh6VrSGi
vzvw5YdZDUU6NuZYnoJHyVKJWa5tJZI+CaTGeIBRUTkEtU7Sl08CBZOLR7idrTbf
Cw5fkOnfARwT4Vc+egHY0EGMlYLcYXlgmrZJNPlvzFo=
`pragma protect end_protected
