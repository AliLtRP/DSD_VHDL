// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
anyQ35UT78lZTe8InYTTeCun1Ka4wcx/OQJvpEeIJ6DwEJfw6kT1E9wgB9qFxBRi
09CNXNPdpQDDEU3lJwDJo4CpK9roGcChku7QoCs/gIBqVclZyZqEZnTSDMlICEpV
pZYE43+eaHyNMFdyiWWKIz5t1nQK5VvepRESSYnap0s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5552)
zPVl7nO0R7MGwulPHgS4mbZaCrexwO0HI3QLH10FxpOCtkPGDQBV+sQBBRy2kXWo
kKTycHprIgFfKO4WfE4OUZXrpAwI8l6y6ppLJp6n0qsK5XMSGSUZT7SIlYgnrLqD
6YhgSGCP99mIzeYK4+QNayk2qlUMuRquGONCUvM1QCELo8fHoT34yLQ2ljldYnCO
cm29/hnnjqNjXEG21ssg99l8u4awTEzeiI09/J0A3IU7ysKbQwNd74vZs269i5It
+E1359KestEeDxoTsqW1yYmZYlryjpaAcMzRRJf+FYnPnFJHCDm7wfICP0PpKGn4
Xi6Xx4XvHMRkXqZjpRgUj3BnGObz2+MUAYT4x0yrcv0WnR99LQZyArMQNHcviaoF
7O/O1PGdalAqDk1mx4lvARU1nCJSjfhEkU39Gr/ntHygMy2E8eZp1c2yUbj34J4Q
5jXN0gkoxLkXtZnubXA+smZvRaeN0VITlMay4eCyky3NQNrWPhlYP7DaXSTPM2QC
vMkPtZ60zde3B8/kbLmHSgNCkcHf0MWVytTi7nb+u/B/iQHJQjRC1KtYSiyy0qQ/
n86bI9rogNCOTI3CsiBwSihI7LQO6jlJT7Qx4SptXcDNBFb60O7zh0koRbxduA+K
5ky14vkWJ4wjBy23TB9FEv24rKa+2Twmo9ERom0PSm+rgM/cHCMACTLSy0z+ir7z
jt/Bf5qitWGA8YA9kfcj0/XP7VDmWjZiaUOXJyKrMPBvQdM3onTGm2YE+Uf5kmcj
xpo/6wOLwRaG0w9jTlWM6vCVQiOy1yAVvMqpHD/1euYNg19qXjyYAOFI3+ZHOWE4
fMV2RpwXELQxUU34rTP76UmyRrfRscvIizykSmh+tWIws8JxCJwPqXb0NtO5/avY
jcZNivs1Zssfb8Vkj7qer1xGIi24XSbxY2J+z3n/U+eMfugkX6FOnJbLBjspCFh7
DRQnCxv+uldVmqcM82PhDQzJjTVi8vovSLWXwrWTugzDDWJFYPI4Fb4LcBKvWEPn
DlpnpHSWFwluFBR5ZEm9+jz8dIiLX+MsSiKxKDFDlE3QV2Ff6LkWr8uOUrW5RK/P
sQ5jVwji5hnB+x0B0bnRQKRFEj6s9GcC5Ujki3n+tIzkKTRWZqD95yi9ge2enbCZ
KfJwyV6vKqz3cwAwQ3ADiOzGQQ87r/n0UwJQQRqW0GGBTw/gL/AAbeASe310m9Bs
7gRT4G+ahtmRijc4qwW7lVZz98lHyDxsuCcpIr55aHIppHhZW4XLvpjoFjIrRWyT
EVxccoSpqi4b8m3VbYJXm8rpgm5Jvl4cYxZo3VDgGbEVZB6lUBWRheYokH9bES2N
dPzCd4EWs0iNne7fS8/L9A/3Duc6RqwpRCQG53Ywjg+MfwyBN8/35fFc8E4/1EMH
Yl60aKxL9zi/X642vcPw1orNWmMhhGJRaOQj7rQhg6wXHbi8M2OeCdlqmd+oqv6w
5viHVDI1Is3LO5ek5j4wTUN3Ysw9a4ZIhfpzVOfWdGZMj+DhGTyZlpzyU9jySVB3
niUeHsrT+zIFQbN62802+8mz/+I3FMUUx7hLObcCBfmV3lHxEHZGquvE4FBO98Rm
+OeZtySC9VyKSXWaKaGgpvf/zs+PNrZ3ULVDYIhIkd/QOjE7L0zWg8mWWLiWiNqW
Fv+IfSAO8Di+qwwL8DVfmHXmo8E97p3mbNM7OUegFolO1XciURxQeXTVNZCLMGjy
y7tG2t45ARC9E6DjxVq/HxHjFhQwQWxVoXN8nkNnJfMmWgge7qxVghKJc8PiLH+p
jrlCfUZzlmLUBgb+kF3MRennuy5c6OF/gRA+Z/6eLTIOAHMSQdHRhxypArf5BaLo
lJ0lcuoMCwIh8/KXe8qgkxpJ6Qk34wAkjBEvHGM2I8nBbK3nVq2fboQpMOHXwo3/
7xJU0tck9WsB8c7Aayyg5I/vFPvG/utsHzSK+xr00Hw6mNcYino43hlk5hIFdit7
ZQhSZMNIVefPZXArx2w1dQZiyv4y/7sNxZt07hb6alKMv5KOVh7pe7OuyXqWYZ2T
Vr1/piyX9v9NGD8as/7BvVvD2W5C8KrnAmAC3ydaYve2UVOpFJwfl8d41TztQCYz
3yAw36ufo61NItrx1fx2We47DZXSYhSFW6Bg1ulrapr+xWPBUR9skVD2ntaiE0Jh
AH+ZohUi8fGit1oQB7+Sqs2BXRcm+0H75hxFjtn/WD7MQ5xyFWYWEfAHI99trnzK
/9vTKDI98ovmQ92mVQXYL8nlydefzSKSwMqikIC7TVKBAYUMZPiGJGqK1vTbMvwF
XsNUETPTZw8U+GShpVHki2AAHIcfoqltm+lKX7NdhmGSGZZG4brRL/A7/ufhu8zw
SnHfC8oCgmOlcdvLw5zDcdbEJuF1P7LNRqRt+TBgTsay0FmDovasCimWDBz/mm26
yNIbset16RVy8LwB5INwfZftp7djU+mByg5lkKs7DX1Hn4JHKcRNdCmmgHb9gmEg
hMGDZlYAmUWSUMgQIJ2iEO6RnGIIzpowmgL5mJ6jWVsZHKwByJONc0QxgWGAx7Np
hhgQ9IffMmN/t1ZEDMA+1/SCNj5c2l+/GPWr5l+dlauQAzNAfqRlXCvdccMe3nz6
i27WT+7YGO+lqYuErp11FC5eV2LL51JtFbFvPdH/kQLt1Bl1hU8Mxme6nKwyJlQE
4O0nJK1H1uwezUMgc0VsE6f3XSrIet+cl/4opzRMhxTDO8r2m61y0H//xV68qo+u
FDAknIl0AD0ziO1SV7D1SeLWd6F7ysxbQCq6UXNv8jhU3FcpKz97e/EFYCoZjOLx
pxwU3HxTfjXcegOT33TarEo6FAzgYpv1W7L2E4XB/PyyyrovOO+84jn7ffbT0UVf
Du52VotAsK5GyVOQ0opH0AdgtJRUIuluDufVQg6NTq29ow95+XFYNYClJ7Nsp5jd
Ehv/gZ07oHdNmn5iIw5YvHZuoa+7ewRLE93MwenH/U4tfJ04U7PhDx6gvg2b3a/w
OjF7rrw0sjN/8aVH6seznZWVBJuUsnC208fRJzkH/E6oTw6ShSJpG5JYrYZmE4OU
kUhWY9g/l1wsBf0XembZBEqCOqCgcO6w8G4v5OkurAJ3RedVznqmtsvVYombo+ck
qzuwoPmjcopTwq/WiTBFbjchwZng7Oe6iKMufGCboOJR61aWvRDMUBHlLqea9k0H
wIpLhU8n7MlV8++HEaqGwjhMqPAHyxIuNFyTOWTj9tLFmcwJnXopqjQi6XRxqYCX
FF5jz9pN0wzBqziNeV5ggI0FFkx7IX3HmzVYeiXs6hzvma122DF9ACuJED+jDQQN
xStB4HtPCNfh/Qy+DzmmTYCBRraAiaYugQzPKiC1JpRJoZsk7mkpMEX9QCjIhReh
cIx69+H8YV7pxQYrHD3CTh7Wqk8QG4iexzsm9ZvIAhSGT+Yw2wctBsTQiRSkUngS
qKvtJXgOw7q2wAuc04U0uS0ejhNE1hRd2vzZzGoNm+A4hFeoDrFnWRga8QjfsWDF
nTpejdWmOL6texCRIcs2tPsGGaAN6cv/4m8ufPMDtCmwuxqL8fYkMyH55fGqzdtA
sIJRWixifMKKIEU+5v5oLwHT/sq/st5ugSK4HEbM0/xmB8H5CYKmLdFd+Wx9RdGz
hKYewuA+tkxSTKBMRdqaUAPPbgDGqsOCMRs/odL3PmTzT8noM/Ch7eYEkl2lXKVq
bAmqPVzp08gR+3s4qzjEb/9K/dAfF2BJU4G1VHBBrNWrTu+zzxssyrLh8wvzaTBS
WUfnNaDBbqryQmFMfJ4ZzuezUsDdZfwrmW3Q0STfXtyMWdYClwsnD8094Mzf/PqA
gtq04OlyQ3rg33c0e8gH1gGzX7H7rW9RyvQO8bBgUnOSo73FLVMY0PP72eRanseJ
E4FCQ+3mlcnGIJjXnkjc3qr27T9FzB3pHkonLAPbsyW9SLJ+wyJAAZIdeajAkgBY
BN4WCkqMjsPW46gJIBA+t7YOFw5QMFKiIYDFrY9TEI1mngi0I84jQXHfXoa8BNWq
QVM9IsiuTW50tCHUXo7jy1vu/MNQMHITbhPfJ5XEAj/EtISaWy15bcqp4/8rG6wX
to5uP0nxTCUfBqMNwHUKlna5dUw7IXQkDyx0pOzk6cajHFxDpMCu0tP2igHIqSF5
teUAV6bsChZIgM+sQXOJ59cZkFcijrr9d7F7EIHkz/k77B5Ae+4HrY0EA5bMbJvZ
vS270xsucrmcCrtt1zki6RIzUgQ3PTHkdjplScchSUf79liVqOBKXjiCiupABfyW
p6mswOV2Ra5jfUk1JCZNtQdp3H3iUhFnB5PMIS2KbxdGx5L9cvzjqZ/xotn+Cqmf
3GXCxRdcDWqDPjhygzMvEDZeqGG/kVoY+clfSful5elneLVVZdjvCdYl6bD/aT/Y
VfqWaRTQHGtHGLOkngLjFuB9NTzjbiRcUtXiuCbF6awpH2OahzTHXJzbnvTs08kB
GGqSQPpiESko7j+Y59Ozy6A7Wp+hMMBPZQbisnIFLfgsdvT6k5q89Lg01WLjxhy3
Yj12N5livIHC3SNeRkaGWb84tubxbhIG8QgmcJ8esHhOv6B/He0tDXKBArtVX1Jc
DlHOGJq7wk3LQ8/K7kPZwD/NVUnbYQunph5jBosjrTMiY/G8sRotNQPAOw1IgOt7
x6m94gM0pTH4UisdooS3GSYHyIyrayEZKqnD5SOxDgpFeOIlXwmCmiNHmn8TMOBR
YfX+Mcpo9scfuSIdnWOpVkk73BhODo96JpK6zi9Wn2mnyLXJDsveddEPLMR6by5a
TK5RB6WQVFqknsphPGZ03KTTBDTUBUay/holP4QnNp/I2MCvNbakKa247dWk5zlq
g940gYGQLAo/1pS9jOyinB5Ma7S7Z4bBEYLS5msHRLuctoQqTHhoTNzJZ2/BvV9Y
Oh8BDfnFiIwgEoDH2qu/H6qmIA7m9Mz3S19E+TjHgD2DuLAxdvcYigUF+Ax0PWGE
lNplwrroX4lT9F2EtmBAJMgePk7C0ren1123aSxR6gQlkqbEyRrIssCl96+o8ert
J70HezbVNU0meBQe0fate4RwZuoJHIqF5djCEdxBAYsQVvDxtL80mlCDVttJEOal
4LPcQkUqxDdFfpvGmNAgzGyuwSrObTF8lQ5ZOQhkKrGbYLuVwDU5VgyOOzvJEFrV
gaWlrgg7/IETZANpLYCNgb8huzjfssa8kxR2lQqUh5/xaxAl9IaNL1OZJBBHO0xJ
9tHXrqH0Wpid3xUdog9ambQPXni7kll0psz46d1CHCvksznNPjwCBm/oOmDHBlNL
RUwAJCiNdC/+Ttm/8DYILj0igW+Eup+1aVtmiOKWoNia1m3CzWa9IWGOufk8lT6C
dJNGxHEP9jg5HBfJo1vbEbEW9TNoJsdfXPropCYeQM8MkIUvEuG8H4Ew38iBccrk
2hGlMasFL4l+YRSsGP1pEbfWvvjKj5s5rnSROrCugpUGXUx627xCL+BqRKi6AUGp
12fdHVlx9byKzCYRbWwCdsgkhOxhyJnZjjxcJ8R2dTrglBMFh2jko16+sqkkzjcB
ZZJ1UoYRMOQbgI8tAPWBjRnEinPhHGD90KS2+EW0+AvfZuZuDbcTqlnvQtyJRRJt
/5Xt8xcGFMiUP+81yzTdtTBQlf5kPn8EyXW/9XrRKKa1cGN7M9gMYTf4tLyt+HaO
rxt+cRXuVbmWYBFaAKLuyyphE1T3ArmFcCCL06+htwUNveKIcahkcBvkLQ5HqENX
RXeb9cINuoIP8JZm9ZiTgIhPUQ26KdlooRWgMkv+qFAMCSZ9JsC+f/xPG3jOUp5E
7AszmhD2jsYft4P9xCHS02PU3ud5t/lfgq7PNMzkjdK8zlee4RZ52SUbTZfb8M+P
l196SVuWVlg0RDboojK3aQBxbWAo0H0P+RDREHa1FFOQmIeWtRjr1DPi1e7dlsj/
w95HJMPJutzhb5iPqJAyvyXovZPZLCSxVkTu0hw2i1QJnlDY4sMVjMWaLXkxNY2J
FB7Al70ZVCmWms7hHP8l1qif/F9Ft6QEyYsG+qh0T2hQtXPhOEQqNAgvIVMRensP
5elrAz9Gn5f9nI4a5eZUwvwetXdWAWqYbyLlcE/kZsYPdqJ83yenAMg9AvzELcKT
LIC2wo2d0+YxrFz5F3DSSe3oz/kFyqJ9HeUb6yOkAaC1Jli1PRKv7ooMUWwsZ0mu
2GLnraVJAN2Dtc/vup0KpPlP4kUTY9FSF+93KNlCO8JnZJHNokxQ1xJUZeehNVt0
e+J6kvTAQEN63Coajr1oq68+LQnKs/BH8twFssE9OZLMT5l6LdzP8IOHUZGCNYdf
8NJXhVQwS0f1JvOJD05aVzzoR80Eec7GxWnwSH/j0sodBodYQaxaFi62SdAhgMBj
ydF3/pP8V2qOsHTFfA8yqJZW6yNIcBZpgMOVmsJz6XY1LUXLg5yZ/pNQ3CWNY02g
Kg7WK32BXGy1lBhxUdtHBTGIWyFuCeqmXf1xBpwf+cq12HPTOw117/vI4cJy8ZJQ
YhRIn9NGbufQpSDk7WzCBn7fAM6sY5jaF+HpeJFFfMBmYTlCCZsPccT+Y1WlNn2B
t8jIE7z/QjPeOu8BXFbCejjrnX+Ndgfc17U41U2wuBdK92izLUh+Bhrmm6SrsHkV
JizAcXjblSd6pim4axfG3c8DoZFIj8Qr1UTQa6IbD4NC9+1B4NhoKTnLuyh+uWXs
7ZvxCDNdZx+1CfJYjSk7nOKvvUh35LwA/qVwBGK7hbsVz7zsCFf+BxxXX3TvVebs
Xz8dXXaAVk+OYQTreXi7ReCX4YXaqpd7SvLA4faNNVewO4+nai1TcsYCHf4uUZEr
WQK5ZkETTOXfySlPf7yeFxT89209Tzpnrn3hDFMWtl5jAIeB+xXZ50yj8wk5tsmo
pM0p8ZiARb9JaGLeEwVAk/O2C+xN6vhkdt/VaK26MCIgNiF2xSKfQPwzNtqUu27Q
92Bsb+n4ZBHSrDjC++qcYhC03XOfKITPzhnWg6x7nkmsqWIEgf6+tqXQ6I474Gzt
cQJJ4XwE/IlayiXEeJmB7RFtiRzEJyS20pa8UIjtBIfAYKkgVnkqoxrf7OAl9PR1
GzJJ7+saXmrqdWbEGGVOMFcaVhGT6Wg3/HxsPSSvWj65I3eJMT39y0LMs5QAzyZ6
X3YJt4NikKiGnMvcne+5EQy70hE4bb7SveP79dEMTsD460ZLlUOYAq9ZnpDpIGUx
bfWQe7hlcKKBa155RT6pVMjdzOWnKQPrU2iTDnLQr3wHXAAuF0ilxAPGzYC0aaKY
dw/mnLXHd8pnMfbEhUtOcZ44mXPRUWy+ZAhkAciqAVJWdrXYdjGSSGF3s7tOPnpb
djTrTBFxNMyfvNZZxlRm1BVAdBRlJ02OIG7H7MLE5/I=
`pragma protect end_protected
