// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ADWqhpSevEF9qeUc6k/xiAcDwXSd/5YD8oyYIqGmnGP3roIs+ugNy4n3vz+3W97P0GS+3M3zIKjQ
uuExuLR6sCX4meJxBbGoeSil7j9fVm9qC+zqIm4cwKgIgE0JqHGdgAnHOp/8Zv2oYkbFCcOCfEbZ
pGWJiof+vlLl8ODKmrs4kXM7K1CSxh7/TgSoSemJ9ZkNr5H6NVz+7DmgeR5w5MKJEw4J3X4v+kC5
hUL93Uok187qquze7tUVvbdmUqRaeyjuAC7tArzwC4aBDHAHKYADgNCl/4LIQKTi6MGkVxRpO86B
2pLCyIaq7bNtclE2hf9UZOX99d1tkXhOj4hCVw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
/RtPZWKoeurxlOEF5LydIj4p3Sjnds+sz9APvoX/EGJOB0Ey9UuBzeklR1M5pmWR2pkAWNf++tie
5Es/DuzdjgZxNNVYVg0jgRCZ8buVK3PqZfNABB93UXV1vIA7XNH7ogSgOXtIbQEYDNMoxZ/1OjnI
uyXsm6SyjXun7+FuoVwcby2s/vmLDdSlXm88ggLWbeUfXiW5Z8vI10czZQER0/KpX42eb0R3TTu5
0NAiiit8e176YW/RCpZlr0q5ql+kglYVDCSniU3ZkmXIcT0g1UH7h0o1kYNktasR676I/f7goy2c
08R7PytPyGzyqnsGz3dV+INcG9y/DtBuTyJXsTB7CGUQmVPOYXTMSoDRoydqozi3AvVH1RhF/CBq
3RsaaII2HucTZC+h9EjIm+dckLci0+WJOe7v6c6VlvaFmo/n9UnnnFSHBBMABfh5pq/nZw0pJ73O
BAvBIEth0HJFWaK1IU3AyCHRTHqexYMukztfY5Gs4gvUf1716vfHVyStPwgwF1IVAwK4fXgG1f8Y
BrPJuk1mxh37c+1RrWfXvpahg0Eu88P6KWEcx4YnlTo3pQoM6WdI0rzApRbYFVqKR2EDBj5rNDdx
D1p9tBJ93nbpnX+m6UB+8TSKVN2KSIgpnhEGX7ZSyiexVSO5GmHRfNoW5wEsNjMLy1tJPSdYuioy
xNatFaGnKQurXg24ukT3/cbG9zrbseJiwV9htrjprKZkyD+mgta1IPwaJmZZ5rRgdsZtCuzaYHWn
uQsJ16K3qChV7eiadk1uFjXr4afj9Z89bcQ/bK0lwdu3pA1auEjzIH70FFeAamys5aPwdMsi4Yu3
9GW61L4djDOHWssw3dZQMGBRO81hfcCRsJ6RaIQXVwiN2jtmrALbeGaFBRzeTQLei+Adt1iDojna
lSnU0/9mt9caAcC8iIKOgwxr4lx6ZXWg+/Nh/XFQkMx+52Y796ZXFWUP3ERecU08I6d0COfA3ERW
nzjBMgk3qKRfBdmtMINOXihs/iuePVVsE2+13PUA4fVeN1mBG55P4LJ5dMp/2mt3veSPau+BdB1d
y0LqcGAaNvfaDrN/xgVCb7nBUl03pGCpsTYPFpD66YjXOaSbhJpEClKHMybUODBWGNnuTfV3HF43
fPfn3ppQMpXunjYYgfEN+i3icDdlzJf3fNqsRUKYuf8O4LQKiwG2c28C+Lx0FG/nReM34ux5c2k6
StRplK18qH/GwrLoMecueQOdK561dMY0xR3BM4LYzB07QcztGsrjjN6ja6xIt8aGsBrAENqCaSET
Vpr2VLBn2c1qMifzIJiBogp9WNNEov+ZUCfOZcH3FvgRNWJF/8QE5LnoScv5oe/5fObdWAyxN2z7
een1NAfeS2fmvYjvQYgU1B30NYxrYwIUTbugfSIuiTH1sOs9POvaA9D/CnHy3t0Rw5oYIFGcthrV
+jluFGk+2LCRgrJRqScYwVE2Knehx/H/34nfJYqQQ96wYrNoBpHp2oX46go0cRgqT1dn2qSRSK2C
/S+T8PjYipwkLJhiCm2ELCDnIbwhxigQgUQoPVlzrPwE749ZJfFVrAeVEzouW+bfSGl/2Z8gwNTf
y0H3ELbBD16vuLHvBJN+tdVnjMiSN3sHC1b0M80meYSsIRHmq3LK9rp6SC7s0f5O4txgGsaqYrXZ
Jdu0OdD3O7ahwJL4fN7SHX3VFGij4H1euqrbm10MvEo55whlh1X4QsZMVZ3l6fiWwZ8Uif+kfvEW
nchODlO9x7241NVv3pjEhVvsRWPoE9n6wH5CbtdVL8eQGMfMF2+zAfdyBsUq6ew5satoXmory/Wy
OAD5Brox8r4KkkY5grc36RJuRyhhvTFYLbQKkoh8DdP33vKtM57nDs0fbEWcB0dTY33gjEaGN0Kw
vpE+8ZpXhtofVGO8CX1fK6JBdv7NmSEeZavmMgxibrpumTjVHLPaAgWUPZtfT0AcKUkP9rrddgxx
MBKXlB7ahvhZjuO9eXbQA/YJYh8Sxc7cRsTtwMyAMDjQn+KYkNk832cenNSWEgo/I8DS1XiwKFiA
R2Oi7izhRbJpdH/BCkJdD1wJm5hvjzSWueevml9a5AjS1fy5C1H7j0Y8UaIujra/nYa618HSI/2+
KSov7lJOKrorVrZgSGZv4gyMx+9deF7Geo6yDuwhfgYl70S1hQNsNHTAKv0lh6iTVuzn67mNzXSJ
sUHYP+pvWsaEkQW5z79hZmM0n/cKzE4RvIxUelOKWeNKFc0XupNa1CVWkQaBwRJTNiB2iDpbX2Al
YVIBbrkeiCJ2pnWtm+gaZqG3stXeL7An/uiClXscNd6T+H8P/rASZ4/gvz7BAk5RTr4Tl2jOZIKA
LqNQORqpv6gSCHvYOSEH3XUsRGNKABT+DTZvMlsIOf6sNJv77/v5hGEn7NTyU/fLwJNVwliqumlO
0bqhXNWqnf5YEOblpHP5B+bMlpQEZmRd/Mj7U9XHLjh1gUaSw9oxnkOy9W7bP+gg3sjqtn+oZCv3
H9Ba/qhokI8efK820Btzdx1Y74gJ4SXomDbdnoZ6YbG5cWRHv4pp1HAIBSK/Ue7Aj1UFpKJ+geNY
j8FfefGi3WoNC/bskbJaDdAOuDTovQaiuEBVatC+6ABS7wpDsZFmpNtTaaDFLaff1BGsKghwNGo7
f6nHc+VXouqOR/u2ldIXF+gflExlYMejDJQm0Q1DfvcdNyrBkgQCzmFivHdv1wObPnZpwTc+v2Hx
/gStQrN3Tj1eKErBDxVKE78EjSYx2ihbITmZWg/GlNOYPy7vpgqL5P9VTnMNG+1EMWvKVPNGg12M
LWdmbXRz2UYhffdZvY9IXXIO0bq4OJBd5uGd+7pwi7B23nXFyKksiizNpsup4TaQxFZWG5MC1MGB
h0bQ5sYletDKlVWRaLDkKN148Rb1816OkcoI6lSYxrtcYCvJh3gJ7NFl90Zs1pYIqbVEjhOwqvKe
xokt9p/6HLV0DGnuhn4IqW9YFYaGA5Z5ONONeIJ8dCHBMNUGsC7ncAaC/VdYvFPLtPb6cau6Vzf3
8//DhTy7P5+seaUN6n9xigN89r9h/7TftzXEcv+ShU3UxfGb5SHy4F8Utm+0AbW9YFv0t7iBJV0+
S4+hmHav7Nl3nUUmyLgF390L50REpJ0BVvXAiXYMWhFSmMbW6lKi3AmYjDoSaOIpMcduSTPufNt/
aB24+JRhXsJWDU2QKhVVhFU/vfXnD1JnaNZS2a79oUo5KNh4Z5id1Wx0KrpNzSEaJee7ap0IZfiw
ZooLjOjrkhrrQYgszS3/b6eMxwkUjKr1zDpsI4eI2X4aumXVn6RP02jvv7USKtpZ4HRgWCDBEFXl
ZqFe8dZPiyN7VkAAvWptECggQ9C5+SNmVSuQ3FRIfgj2K5uLc4fhZ4oU5bpFvV3lN0prVpEQe2vW
hkZPdtxQCGBRryyRpCQ6jfo0kQLxjLFeAK+2wLfIP/sEH6t5EEqYIgI7LuhjDN8kCaAJDdudLQUD
b/uDzIfG/IEJE4G7Lo1mYbLqiqt5Zm2lXK7+4TDiEJPscMR23jSX2suX97/9techEdXheU70Ln2t
7PlTnHHQhoo/5ifmHR9+vQu4RO+rOjYTfhN0r+IRBzjkqoSH0GfXU9vnQ/5gpo3gfrYT7AoXNtdh
t8i0+Du0+rTbRwcGZzdnIIb0367ayg1AADv76Dja890UA6oEmYSrl2aggUXeQ0AftOOdLPiClhia
uIuD3aNfHCa55l2ZpRnpiGF7gROupDqxez8FlAq54+mVVyFJvauhY/a0E//nilX/U5XcT4v53Yon
bZmftn0+sJvdn1lWCQKGvp9WeWAY45zVqaqwzLWdJqF6UgrlIgnpG+nN9+Ki6CoiCLy9POANXgGy
OpKJS9v8gLPSpvjWMfNVcp8zAAGNVC9xJcPGvOCQ80y72FUXdyz2F/bXrVSk9u7cPLycLatZ2jSW
rcOsTp/gENqXzTRYBBjVX2AcQACj5kpmGvEVjvadqmJ9MpNijxxmEuiffMIl3MQDBHUqeiHpK1qu
c3FxZVAE9cGEchg4Kfg/hDlNclZaSt6N5r25hWth+4jt+TE+Pwky1jKFD3E5BRoAT5dKlX96g3NS
nNKg4O5nrCf+goSuM2zMycdgrkA1cn/UsGCHmqG8GT6ZMKczAjOm6nIDcv+rajGADWTDV/vkISki
y72EDQ0rYUTjiutsmX/D4qWEAd0KtvkgSF0eWjR6fZ1KnhquXGuipkyRV5ZBOabtCJ/jAQKSUwdr
Dgskvgn+vk4pbeL6a6erotjoiM7BMefHzaKyqAK1u9jfrsJspsTIdV9s7gonRfoBv+HLhtCKEkTj
h3B1xHIijQpeJI8Cu4OVqZ8+37puqfrclJUhfRqhXyMmchXSi83XUej2q05X+AAF7nbEco0I1T6D
wMBIE2sl41H6DwTa1qCfTvbZ5h74ZbfYFmQ9YIPsw5a8GRH+b8Xw6XXqqLSbLwghmNScwb44pi7F
GTp4aw8m/jBJB/ywyJfiILbhrP9ywEhGUJbW2xTwP2vWGoBlzZXWCHJHqNo60Bx02+QhjqHauCsK
yFxlB1K2OwJlK6hCIlfbL+Xc2cxK7jrnSDFKgKegLv6IY00+8uCt2IzxA8xsUiKIDf9pTkGw0QKk
zekywc1sc3BiWNprcEWtjCiLfUCTvYVu6XqSdT5rjMiMDZMIie5++eSG+dI7ojAkI4IF8JcAVeQI
6bBeSc/86exlcCZVJoB8BOlS/Y6ZHxfHO5k7fuu0/iufGYnNUImYcX9gwxvtppAZ2o6rpAcTe9b+
bTpI3jEIaHL/VANDq0rbOFR9+5WuIR0RcBY2u7yDQw2//SqtvdZFvxfZTRW6ZQea145gx5pgnq0M
6WTOK+m1dUcRWEOwGO+hh7cJGI0mytPKTGhGB7F3Oezs0YON15XbAHchKMpRr6wZE/yK0YjeTxn4
5hO38JFzClwm/Px/ub6XO5ynp/jvJ0Oy1jOnmzUoGgsUqCcRyvpN8KO7QMzjUu3qEb6A/wOfwImo
FXnnk1vlYYYcxwTCs5rT5fK1368C7obdj04KyfQDZcb9fA9pNH6a67cOEomuNlx1e1sFQxxUC7kD
ddGxyBNKgkp+uTVhiaCLrhWI41toI8CfkJ0PJ0SePXA0g/pWlcsg0olmX1ziNpF6jCh+exxqhvqH
UowdWfoEOo4h5wemNRg098VsAbe+8rV/9eN+h5agoxfXE5Uigc0UgU9E0Gg/Uj+fJ0tV/th9cNxV
dMKh6/ZdwGehz8EPP8wYy2Ll0gMrwMul2zssIAAmEKTyEafnuvUdCnTAN98jc3GiNwGejDLU4TAt
PkUwM+K6heU0vUsFP4Qi1S+kpJiGbjuJVV4DMyTCJ+EIhAtGEZ/b2YpTBLJPxGiOYpQ/jL77Tgo9
fBFDkZWKWjmk2LOygAFammjw1i+8VCy2SHBvM+3XykkCIRTVgWHn53894edzLO9391T9YbC/m1ZC
193jot3CEV4aEiRbXwAw6KrzERkF749cXlCjh3ncrE/qdoEFFLvPyXQe9OvmfKyhxbkXbzKFy6eQ
BE7hMKccTqDXsjPcGSO1OlJbtWdd/F5ZHym3vfdJUDkp8EIatpZzEskhtKZY/bM3o531fiGSpO2k
w8osQk+mKNWqhf+UOE6fhNOIg9Tjht14UI0fGYpp4mcVfBi8uf2HlqM2fxDjlVm9GKEvBczvW6pk
yqJgKJegL0oCefp+ug+CZeQVGmEPex4Jblm30TbhCBE9FYG2j5mVrk4V5Xb6gTekKHsSTIk9A8JC
g72j/zZagtv4XQEqhYEN6qasrdjPsTMbUlV7W75bnXmeSwJAVDD8tY0iA3Hlx4EssLk3PFOFdWIn
eQM0THqdyuJuQZUgWdvgN1sWYkkLmARl3sjsY7Jx+J+/DFv/MMyaq++w8esE1z8mZRlOWp0C3k/J
N9bmHH16QYCUhfwEvIRzzTqZBJlSTdPiOGET/mQKeRX2hkpX8nvd/N7qd5gcTwlSqoPACq+lhDqY
aVWIL8jHmh7t+5+04kl/bqTLYWTIzDteJTaiPvqpH7xm4M5ymo5KXdVUUPJQ5/cKlRnoYwBvVLRm
Hgke57w4oOtjJo1+AIeuddlTBD+GKc19KjLQm+BY4cU0F+q5a2Mrb+0GSyDcMe4n8HL0i8x46WHy
SPnapMN/Yo2xYewl28HYB5tn5TYmmTHG7YyDKnPyq96DGxTakg9dzKg3EZAk4XGjXQxBKEh4KULT
IUanfXyBbEpdyp4LJzNdZIGhwuJYW7C+skuZ8WCH68Z2IXSYVkBRowf2Fvfb9jEH2DYS2RQazx4V
K3TOVQ9+wdryxSDv+a7TxNRDqxzvZDxKbOM0FaAtckabcAffZARVkyrTgdHHEgToY6Hp8PG+P3/O
+FgLX+XSqza550FWDys30kJKv25g133sYmdfVFgyCp869zuirnsEEvFxolQxrlD88fy7crGcdVd7
b0Ts2md3i8b/QyAbquFFrzk0rnHfAaaP1J9IZXuaZyYhgMYwsLF6hfOpp72QWwujexXMFWFw/+Gn
6WeyHeK3MkfrBhwdSEb4Iek93l1jAoZcnafoxJxloOWdXH860jCYifa0c0cxfWy4LmFYQMHiajmB
yVbTVqWf70YfaIlT9c/qBEkw9x4QEQcxfV7ofrWuCpHKiv90O6vjKYdOktU7YEkNs4Ly/2J5hTlX
ee0WqIvmbtBTgpY80Mwo+OCSGwuX5yOe/BivXNC2EXirhM+Aah0BtqUCjR8bphtarWE8dsATIy2u
xBovDU/s8k8rF8iK62Ry63CiQ+w/XKLMsTawPuLbzTLVC1YuCDaKoxeK3lhvGP+JXgAQeeizNBHA
0V4LpVja67OvbSMy7vhOzqTMVuqcLbjvg5iIyAVsMmNUlJEBcr3Xbk72vqMO7oCg4aIGxOvsBOB2
JtZcbiD0NgO4k7fpy/pzSFKE/eGemQjaiFAb0k/IzprZx/nctqhh3r8YFNIVuvgi2FzcLmsF9Ryw
w8CZXzQkjqBw8n6gr8/tCr1FAs5YHZdHTOxcsIq+Kox8sdupLywWljMZi98UQHapM9WGhsw9zBZu
tWehBRlhY6ufX78n4He10BmZg3mzG+ngnqnmsbq4bWRGdFUvPTpRhq/UIiqNMF+MP3hwpcQFkfp3
nZ0sdEV8o3ErtA13K24qV7WJ/rhD8Guu/1pjCXMzhKV09slWQAb4/bIzdtqKB5fND1x4Tkj516g1
YZgPRTGhyE4SUOBPKe71YSWsPVfMBXCBU+uPCguKzUJa94595mKBqxsv5smA3KMt6vbI31oFxOF5
dQ3iOZ/+8s9iDWLmXSCmKuvWty1yP41AzJShp5tPBdVD7j1FXiNCQjBaqv3dhz8bj7XnFfpq+Itz
7+68Mg8XpOmx3utkjTjL6A5ZGnVHFj9cGBRNwZ8ObFbx0aQOklSMFKbf3Ni34Cj/wbGOSCARBanx
RQJfgZpZraWFAgsWmMYF3evcz6KyHFIP0jt49OlBnbQcwsiEe9u2zlJca+5/sMVHPn9SVnQOGwBW
8CR/bpbVIq432AeY5dzdtpxYoR5plKl67eS293xXQ1MBPwSjxM9ZX9IsQSpTYVP5XNbBYUNidYD7
N+jFQ4DQJJEpSVxTJ7J6lB55Fg9Fb3GXM95BB0MsN4xsTX2JOyzVLz7tmxT7G+h0gy/T7zwc+DcM
v2HBm0wReU79eA/hG+r+opkb9qX3mK3QBbJlqI482GO4vKShlYhOiWflVyHNBHH9v4RqthQMLT/Y
qUetU807JyG11ryHZFFFLd2bgNJsZ3NyiGT67tUBmtQ+b4vdCE3z+/VbZrpLoV+vDSAPU40dK7Ra
VIZhF1skps/9vbS26NsnO4sQdsPHFY1jWHuhTlBc1r9HUN3nzoY3JO5fyvR59a8mhItPdqilYB62
VoDSPWVzhgJj/icUWQSzZ2BeJjKnSG2zVrx9PlSUHb8e1qs5XZLlztJ9wLJblgisUF6Mv/qOzmkU
RNUGWz8V+nfCytwdsdX7C2DMGpjmapDinCsQiOgk4NAnyqrtREnUgKdsZ3BTwutphb4q+wE0x9rG
vy9MYtG2P+JPV28BaOQwhW8bigbGunHixRMh/hORoUiescxqhrfB0OtR49uA6dNw8+KC6Zf3qpHZ
FBrCg0nrlA32nKcYf/FB380VeHW3DxSkjKZy03THkqw7FNsLIK5YlYun886nm6EbdC45O+NL3+W7
RCJpDuOTNyO++s1sgfVt93UsGnvpVHSly7XyWnipnO0XMkU9nbbWh6eQw91LW/DvWZfOnFLkNLdv
2lWiowVohPbYb5B7nl2yvKIURkObwcVn9DEs1k+U/17+KHAUBkx5bRK1ht0mGI+/T/v8XY55bPrU
DS9g53PnnMjM+6sU/gsrLMMB39Cbaw0fNI7G5ubkkvCydxY9l/68bNB1f0mnrT9XCo0peaxFENBy
1gXmZ3+3gX0tlqNDvcT3wb613EqqRIyQnmyhbRw7nTlv5Fms8PJT3vnmLYvR+veiom/hvxqgxB7a
tn8ELWS8eYFdjFVYrnnrU9QZLBVVACn/BOIGg6OUiw+9AotZFhO4sM+/9OU6YloGOZhMV8DEASE3
qk0gBdrOwvDxcqrb6wzDbfmYMnBmS/+NPeFtiB96M719WkCVtl6TR/p6556lge5Xq4z3sOUmUrxt
DKnZWelvyi4mhI/2C+/y90q5R8dyz96S1aSuwwobQWtu3VwOf9o1EqpSNEO9MXoCGzmomkzrMFgQ
V5FFbqz5VgJAWHohC32sNZ0ccHA45kUQJWMWf1Q+if/U/C6XMxMrAN1TCwgHCf7Vd+It/XS+5Rch
39x4wHlmpPmZaVevrqRRTUF5vXVwD0SmJ8SIMaKkP0ZdjJxcD+hCjOFEDJuhT1IdVOqfCclFIuGF
r3mY99GC8I3MhIszjvQKLf9qGlcqI7FIr5ef+COkGlcArSoVFQDFgP0tUZo+C1/410ygaiy7i327
QNgUfQdD0+XZjys0dEVYR+fcAiWhAY6g4mJ7EeIp3bPqBA0kNcIE7wZvh8FbdQSku8T7p1tr7oWV
JfdLv7/xadrMh2pgGIqtwgK9CxpmaZOZgkQ0Sa1QJXjkhYuLjDIbUuVwN6tn1EpjnIv08jUkIyYC
Ww/dVR+srhvn48oLlkGM9IQqPFOwbJhFXuFZXxjiZL0a1DQNeh97krWXjfECvv2Xv9M23Cc4oOex
+4A2u2/AGGPtsdru5LW4YxGoCyIFONj8emouYuvEpPqj4Dah45BV/ijOO0kyvMnjDVYADO8cckD6
jOhHMcxr+gsrg+TCrs+J/bbDmPzzL5z6NniU/qpRaggUU9cmxAoVPHYjojXc6pEd9di90erGxQ6l
NlWhEysB5nwfDofMUR8hAujScNefjaV9i+E/zupe5ON5+HbpI63cBnWzUmqqbBeqULfb5sRvxTQj
eqW71cgiGuVu+QeB1VN+D5fAVMiYXqfTX6pQw3KRDVTLuEW1rMnXYgJpwxhNkWO/8dAHDM8f7viT
GDOVXeViv3N1uHEkGU+gHhDwdK1rEzltPIVF+Av/NMGSnvUCz5pHHrlonNFgtgRMpUKIPNjaOL8Z
IT0W5EWoCsHreHO99asY64tLZDKcqDJyKsU5b7M9qFWfEcDKGIEU0GWh7AzYyEPmFpL2ieFplErl
s8M4ReH04aiOqNdq2k5VfcSlm4KD5QR/EOM0JG0rx2Se3iV+9W4TZdd8+tioq2G9zrrC3J7jreLZ
PWwCh6Y/lFE1Attl5nkYkL5j1NLhkBgKLYlkJ2riM/DNktZBa1JL7wUWS72rQpgKacXNMKh7VCnc
9fdOKhfw/kRBMrryK8VVRb+dqnFn2QupOW7S6S4tPX3OGkuBrLhsSt3473+GRJMw2eJk6/14tuC+
WrPUBY0/enX+CNZTrItYBED6vWtukC+XBufiPciPpP0JEYk4rbC2nVOqdxb2bmNJIXIUzhazMMuV
wjWtWhBIySOy4R3yl9BC61dvUneR+tKAijQ/oMZJJxkPOrcAkaz6a+AGasjo4XWj5mjccx0BcX1V
AWZ9tBZ5NwHwIgQVgfqk6C9WOf+oaJFIAniObEkXzVg6h3o1U1AePRRJqW87B66Nhznf7lhALoFJ
Lx1jwv2lmJ7g+8w4a9DqLoqvAwKfaK31gUev9xsef03qojgn1UFqR0pml96/2cQl0/5PoiuXc5X0
vx+dUddAAehu3f18+uranWGBL26B7ZVq/bMiTlaqUzi6ymbxCRxcJuRwMjgBcj8Jf1yYirHv1OfQ
0KCuqWrFdJJzavL5J6BpDVNco8Dus2DDfTPYOTBz839oNpbeMkrbaOvTPnP253niyBRmktYFfoCm
LNcnC2UsZv1oHQ4mamEWqe0HtpHMi+N+beaaKWT/UZwiguzWpqlQ+w1FqnFA9wVIOEYMQ+Y2Uh7s
HFQ3e4q39qw4PNS2KVCV8zK+l8vPC5rUR/iKnVpfLUSDLwhd17n1YjU+0dNDEaNKWvxo2UASK2aN
aQwWqzOMLEc4w7XAbYBgxRJ2vFxhkLke7rF8Qjggl4OMGWxG0cOsy+4SiXUkG4uvH3f25jIn8KO+
KunXTs2ulebhxE2KUzLxP324k1pFgUb4bOEbdbNlsWRguqU9n2xLb7vhLzjS2+NgYG4XmJGIY0hU
kI44lGKBV4pHIUpGeYItSDJ9gygccdtDnQza9K9W7N+DxCpUtqpm0j2kQFdg1UUSBkOX6et1Zs9g
Qte7hmpdwLfmcyevbP14FXoZyCCwawq9CgbEbfMCwE55HL1R9zC2ee6g2xyMOTb1xxNsVuUMGBdx
3bGi+m5bThoVB5pgBbNBiXY9HnKyal5quE2KaDJq5j72H98SJoGWeDdQlvdICIlmFCjtcTiRLZd3
SQKJ3un0O86BnpsHFBdyrL/zn/4UwQJVLdpKpHljFdpdrXe5AgTXk24oN0ckJ90+WcVOfIyIKwdn
PSAXraXI9/TpSu7WG/jnAnt9UIA1zwX+Cj4mUBSzboOoXhSAmK0hwAwgTbIIPy77i83jTQ1CCsUm
s7GBY4v4lRUaJ72NjxtlWbTSPXgeiWXsbGiGsJEW2Zj2PRruwAWh4Qicn8XXX8isRYXo9cNsXyrX
mBYWKwlDuBcVZBt3f/uPY3qZe403Flwf19DLj1prb2zEm+ng7FRM+f9w7wgPhwKmrnnPYpa2cIDO
pv0LM1u8Q9cKPumbErlh3BAs51Zljchxr8z9dTW7iFdBItqBxOa0Wf1VVjQreHutYcClFFMM+I95
Gw3A3zZ1OB20lrAA90zLdf7Rl1gWV4xaJLNr4Qqow2XBbmbazeNpmWPmTsazlrxUFLWAejrC71Xr
bGT2CwYhhhzS6ZL+pEH4386u2P0e0PFsv77emIs+rgb1W0SHVUemcKifXjGWjG3Td/5oboejK2E3
qv+CAjvtsShY3TFywi4g8m1odyYQJofx0zWDSKxWPlcF/0+cdJ32dDPrpNIc2YUuVq3YFO7EvaGa
5+329VgA8+/UYNIyiQxpZCoD3o5KeyMJbnwXtMiTgQK6KcjpwB/6GGCcVRp7A0ZbRv2sOSJsU0Ok
ukdssPDzcH1RsaypGMj0e3LTlWjRvDhSG5kqlnxCEPX74wKJxMDQcA2q20HUY3gSMPi2Q8bwL6sy
wbTqYx2cM7ax9pdvWcmq+sv673URGh7zNPpEV6egp9JuBiOGpeh20YdEO7h2PXD3/fpe5oSiOE6F
YGOgQb/ZKZ2DoLzyxkMW6bYDRvMDSIZGA89UTN1pU/hyo9vevepVu4OOmUsqydCY00g63k0ufyb5
P8G0kBgJc4RlnVfhSmmArCUXnX/P2Pr5xiuCeAcKx36e+y3GKrkAuLFjObh2QXbuoYjHxkgQo78E
fqHPvwWFZvhODox2LuELntyW7agpbKWP3s+QPWr2zwnvxIfTHks9CBZDQ21MsKTUoWhlgwWrh2RQ
CCHlCiaCAESiIOsZ7dMhTcJfdaCe9xM2zv+2M1qGbFkAWpHsaVveSEutqaDDrfb/YDvxiYYn88kw
sqtoG0vDhubcTcKqU6UexT96qCCu5M+OkArkTj6EW7B4mlcbQzjTw3WD5g8RAj8Zf8AZJjeYdNGV
OVHSH17+Dt3iPtA29GE4iMqBe7B5bYnAsM52SVaHXvydTgdRklg4/qmYRS5iq0/Yw0fH8PwWD6S8
wromXHr8a5B+/PaH5PEyzStyVhVWDws3CyagZeghOY3GMhwsweSX/1xxgKUxdb4bx3AloCxGTEIz
tpmzvw2dD9KYqR+wfuC+GqtbboHNChT5qeWuJNPS4/89IC9LMj2mLneZN3QAcSt8J5HvTHI1oZml
TRl01PZNQQQUuTUwUashrXw2L3aTalkUGx6rdQt/mxK5hYQ8aYL1pMk3YAbpINXuWgwE03golfIp
Hq+IB2G3K/xByvpjYfJV6aJcnZjRGZDG/ydpzf1s0omES4d5N51SP/xrKBBQOegxoyzVC7Mln3mp
o9Qm6135kwkxTpMGT70vN6B1l059murYXGNfYFENFVFIN30xApyzQHE8hRg04f5GMQU8QaiPfeNO
QmsC8cnOW5/ckstOiRKPuerfxIXdko6WK2+gVu3iN/Iyxu95s+U7Ch1S8BHtIdv07vPH7g2ucdRU
dSTkKZYcjye1LB9qYmowp+71ifP+69cWNAQ/1tLbJ0reEhXywPfN6EWxPVOKFviufPHHJoSmxS70
we9i1vd4iFBmeXulWRZfvclGZRBi5vHWhKIb7XToXpyq4ffHPnIphFZQosU3pKL9BC4wyeMMqsQx
edGnYobhVEflbLCRoIYcAbVsWnNO6ApG/cci62KPQ8YIKrq8bS3i+imAmkhqpgQ0zDERGmaJEoYh
DttLp5JNnxdem1j3oA1c17F8HaBnTkOdUxpKcQuZO2AKvAp6XysgUQ9Uzw749R4UV/zghtBhrkm9
1XdV8+fE162OtMR7kLiDCkAyKOzgB+7MVHVGx6IymUT5h1LPpJnW+JPDc4jfpuGiF7khdUhdycvJ
pJO8bq0ip9IXxIE5GnwryFx+rW+MJfJxHO6/HuMS5P4vkEtPbdLzYGwveA5DKVcQK/F+0DCrAZHl
nBpjChujP5E0JgluyrlTZIwlfHxpygX6W927IflnzWWgCux6WZYSmZNGlWh6wqVRRDwl+erbQpFZ
pcx8J2QOIe+TNsnP3Bsg2j1f8qKZ3VNSW7pQ8qOFQdbvFxKM/IAbJCaBb5ihxkvjkAL3ZOyO+2v+
Mcg5Vm0KqAcwh7FobhoYwAZCcrls88LubtNA6R0xXTkeGhj8w1Je2RTHAcnX77ALnXBxhKAGlveX
u8NhgcgQxhbmaFib1jBe3k4sVnEfp1Wy4DSym0clcBO5Q+7aHAOABBiIxZn22jYbZL8i7Xbxf5ty
jWo9uc9wYO0n64S+ipQtFYpAmfqjLWNOEbjy2adloM/1iPKKzGFNtdrlqvq82uc+05GuGUC0AwBg
tHs2LTVJhY2qauGeZTM7yetvhz+eWSTzTs41osPnCwrgXidDOYEmJaX6U55VzCuYPRywUee0od4I
lojsd9ISVrw8MFo20UEh1Pqw8La2sOgOQi7UVdrnUEoiF+KTMx/mOe2gmIzDO5SjQwkW6wS7s9sm
c0GePcyPe8T6Mwq12ujqx175vL2+X5qO57s7P+3oaiHkTiVRPTzkxGMOOE4hn60B2Y+wRX4ZVJmc
DP6xtQEoGlghGPzfFMXEh8tJNDi0gh79EeMF3DsfY5aDQgVHomGa/fyF97psxXori7XbYvFZmzTW
wo2ZOf99nlutUf0j5VRNhopJwhtrAT7/C4uIB+zIUlhrRAcEuG8056WNBseofOHL9GGsh0EPkPIV
5f4tC9zV39m46y+KKYg0AI9LrPfKtXMLWpXuztjh2pxPq3ldieU1l4TybYxLGLX3G5mbF3a48itN
gdY8Xc/f0EchDEqbkBZImFRuvD2pfuUr2M3uRUM0hduqbZxzS0yk12H6gf3XqLXD3Ru9xBlZ/Weh
FXP4UC7Mb/voJC8qMaR3Hdc+uiHZ430QN3c8hjZlCakH5vMcX9bCgDEm5Uzhbs1ZmHx2dIbdTVz3
CfXoncAA2xbZu+YqWMPsZQEtrxQ2tDpQPOde1/O8IBKeD5US2xssm2HgkHtSY6xB0Unpm27xSWcx
/PeoA4TDZfELcOyHUg9pnzEKkNt6VH57kcwkSLPTVLMeVOX7YyPqtMibJZxOO1oGkzpPFBRA+X8h
Iv0FBKDR3vzTH4E82bh0Yqkc4uReQWZMAsHtUaFtu3zDNo2gc0UpeYSkTNkozOwvTbY9X0AbuyWF
q950liaomaeisXwyXEOy8fh/ZopKCnsJ+tk6MBvYNipv8UhubTc3RWeCTQmwo4uMaEtSTswnUmCP
UMhjxVmMBzD5LaGa5Ss6gUkL9W3HPKmN01g2wH1BIWVor3Ur7E7IPIIG3T+8BNfLwoaux5QBDFGG
keG+H6hMJ/TQOS2kGizBVoesAIwOB1MSbJThW1b4XOj4RnYp/VCunfIoob2hXvorrOTaOQAp3fkw
nUAPsg1oIgfyDMWnfFUemx+OmSns33vVo/mzq7fojipZf8G4ZKFVQZLDYWQNXNBW116wqF80UH5v
FbMrpYtldgTynoxjd4ImT2y59Sef74xWxz8x4O9xljC8gJIizruIYN9Fi9CTpilnz7zYsG6BE9y9
oxnQXSn+lX8Qqoq4wNS6+TB/1C+j1sx/K11GpE1CV1WGpMlFJDste/OPlc2SVqaA8uLL/WjcvJsv
f09PYC+4tnj3WB+4oYOMTt2GZ1IGmvmf+fOjwt/y9PbQGEBPDcGx+5iwAW0E+Beb4JE1vdsxZbgl
LWNnQis/oxALzRC0wNGe1vqDRJE+1crZjbuHh/A/F0VuUDM8/LE32AEB+DmgsYAp1xeXXPGbdtAD
tjrsovH36fLyE3TmqPnW3OLg3jUs9t6BNm6HxRS5XgE0vSAYY1VFtCyACVlFziGE3wcNW/0lq0kn
3cWXqoIj/GNv2DthO8QL5MRWcIFjRk3nxc8vZc0Ej751ZaLEmeMSNlEOOj8pt3r9TOtxUtJCicin
SXIKWBz+Pxv3E/nE0G3BXBsEfvMwaME1l+vLX+OcfvZ6TUZK8ulKjuP+f0XERbOCFjD4qFvBPCnD
qAMl6TKuIXh+Q8OstmepZaVms/GvcHAdd+I6faS5NlZQdSZgmRqX9GyGUf4J0H/j2CAbJ39ROZX0
vpDMQwR9/1pP+61A2HL0IdxMB31iawDhMvTpvdEK/lVsQy/Ti/LZ9cnZ+UMjRp8oz0Xj5ACvkJIB
cmDfiQEgozLqATQ9wlJauCW5E7pHQz+qBGpGtHfRBJGdEAGS6o2sSmh5F8cTVas/+Y0AJ6bPslAF
GokyyJI2/b1xu43EJuk64rD0NEUk5M+Nvk/2ASpUt3YRuJMM5+vFLSw5jsLbAp70F3eX8cYoVJs7
lbfCWDZPlmkQvHoK02VVyTsLkqBeVfBifKbyX0dS/9L6NzS51K/GdVL6NIxOT0dwMKwhXDrXJCpA
6VdbDY2i99YfcGxoPrG02hvgh7zVbIikXP97hO/VAlTLg5erCgHiYJA3HTw39BqiA0cUwF8/BaJt
uzZ9mUq3yANx9YE+t9CzCZu50c2b/xfC8qLtSN6KnT5qzMDf8Lwz9mEWmNKgBB9otPpBUk1rAKWH
Zdv53Q6sEciMjgDEUcYOBNAYl3yFTbeNVBx3sRoQ8L0Hx5u+KhIZ99y/Q69v5+cReoUl/UBvKuyQ
S42jMmyIxUSOPpA0OSbVqXy93CLyqGO2HiPHj9SZLTlSp/SfS01YpnmCTo3GUrC+5V76wqUgtFla
TnQ1rT1R6PeWR21LyNHQOUtSvM73cok2tbE2H26FfjN/Gvd1+fPEK6iEDq3dSiHAETLNJAsn6ue2
Nb8lqZImJvnAV8vy1EWErqKxueydSZxpqkFoYmmP91ph9IUIDjIj7fYiJlhMtpNzXSvq8GNttyvW
eoWhOytWvXVBNbQQdV4M/qsFV/gCgE4KOmwp+dp6TlE8hOadhxFpvRb7dMwrO8dYTg/X7Vbx40T/
K5JsGMVRnL2/pf2tfHG9TBSXP/02sUjV1FUIrGRJHE/p5IsBFxn+mwEKEmN6Huu1wQ04CqThBe8a
xJzrhu0CQC+wgObGcabW4vzH/I2xHgKbvs9dU+dIPR2+z5mjfDTnb7K9Yb2trGQs7ddtsKiREPPm
8mkrJ6ZX5bGt/DBR8kTVc4bjmhLilpJrsqHo39aDgrFg4naP3XLXiZ9uFcavxOyN/U+FEi7JZ1df
zKIv31ie6kIGGg7fGWw+FWZWl4bYgzfJ2ubFhfSp185hdRWZX7rULvmE5jOdD3aQVgWk8iQ/TdjE
XEyPhfK5ThmjmvX8JeYdEmomtIDFm93sy/uUalRIEyRhkqMYL+Zf4exTtkfiVlx0h8lQoPJGQzXv
A5FaC4YqrktupIYvQcwMNzDLJv/SojRCrSYTZjagw1tqVGtf3YZU0QtbJTthcIjQnPv97yGvm7vs
hHDsucZDoHokHQQkw7JWXn626bWbUEO0MVxhdfzWTAFlTPSMcB46YhGlGScz0v0i2YATc/ZYvWUD
uqCrLRcWP78UUuFFrURTYt5KL8lme6aMz23FkJ9zLV1Eh+tpA+tXqj2zxQLrGhJHm0m6Tl3gE3D5
62I/5xkAmomsrhq6ws/qn3Rll2lA7am6fzxwoFKwK2DHJ+A+2FK8xoRSY+LpBHy6v/KPL07etRF5
KhhZtxbgDRle3+05p8WHoxcuAM0e0QFz/S8jjsD413zXb3qV5Kgf+QrefVUcf/dfteERMs3Ii5cq
uqEhXp4rVmQuv4IfeK/gG/Dh8SIzkNni8znDe52Cs/9cL6dlpojbTf6iF+iv9lrP99ZYZ42rPOlk
bs6UTJnqTnnHrJcZ2lLsO4oXWAM304O4cmLqAkMgDOa1iEDTce4DG8rQWY1kgyoG11SIMVjzQ7nE
aGdnF8sxbfaXioBau6nqiUcDgn/E+r0QOOKYAANpNpbE1LD5crH8NPMRbcZ3Zj17P9Sde2wONAGE
LdrMOMGEfdsdC23/90chYJl0AhyMF3ZxkvhWwTRhDO/lbpPfPBVBW7kXUrhX4496qrH3Ed21McZx
65KnCi2SEqkFJKaSdwHyef3obEXHG1g4CydcnnjN/4oD1f9CeKGhsfODIyde0PF/QFzBsCHd3IwQ
zp8x/ilvCshmV6dQy8fnJIitcwfEF92JjVCiS87A6w5SNq04z2JMvwVxUpEZlAP75EiUrWRrokXk
5foyV1IhDpGsRz4eHmGRKBOhDc+ZPQxJ5Q8ObqfMOrAWUAzYfYOuCGQNmeSrtd485J6r4ruJD5te
AVC2BuJ18tEKi3FSnaEIteLHKltoatlbs3loDuX75jMebSh4uEFzBtsnpVGZ0MPMP8W3IprXk8dR
k9vb7R57++HYR7WVFf+xZ8tGelmSEWDzrkezpYwsQjbEXfCbSa3PlepmmhtbW0K5o9aNNGGvID1x
C4xZka+yg+h7CdCdvb2L8eQWwpYZ2tVnu7V4bY8HGPF1zntSABknmluyeLRmlsjXceksQ5XPJCGp
zkarRZ/Z2wrXGmjoerwQJ+mp0d1FMPq/62uBaiVYSFo41zXxntkpRdgN7ZEYm6ej8JP1ttMCgHnE
ReKze1ANVpg=
`pragma protect end_protected
