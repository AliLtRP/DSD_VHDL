// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PXghcTQJ3c4szUhXD06DEiCHsOcI/ZoWu8hH3F6+bREjyr0RHMZJ97zUyUpMePpt
UTa/1IqOOeppJnFkeab81DU/kTxLmbzQsdsaAOzkXXZdhn2YNNsyi/hEca4/jJF4
8V87GV30S3kqJPKzfSwaH0cMAMy7TkWHeeRjSqKk/3o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10704)
Xuuimo4iPzJ6wbJHo8Z92iN052iLqahUaT26xl3+nIBPT/DrJFYB7kSTAvJk6qVI
xcYBVCRCm7oz78mKV8Y2K+/PPVU6hlnVcjd969JiMU5FuMbJYL0JfORf2+JZd+ff
44zmiSuNHAYnB7hcL4gHeL72xmFJ8XGWZKHEkTT6u+NwNcVdosnyLwViwV2cq5Jq
h5VQBX/gaxnvfKfDRnHsp/MiJ3ccJFdZaD/hnvWYW+R1LQX7qSHoFuk1SzKR1rU/
mrXOZVP5cQLKTDRzK0Au5kzYoX614toGnGDQpKs20QAOi6YtZe8yQG+rstPFDBxf
nhiivW4pXhKahODdt7NkDflUrRwDvLPcYHpI+OiNqbglDxIPiopUOHS5Pz8h38pw
16blfOU6eHP6S1wzsohM5SSQLBL0djtXbUDrgBUYlgYNRHTsvrkDMhVuJaIHFCNX
+TCu+8Z0mUsYomunp+iRAWOBcpl3jzKnArR1k2TOB1j5tryb9X2cCB4qTOQdDt29
JQ9bV1++sYR4PpZVtEKRuECQcMslqm/WAYIuO6SLV9RHtzz5Uu+nzQopbaMXZjcZ
ICaJevXpFAJJCs50q6WRPLK7f71biJRHkWPv30LTXf/UG37RZevne0FW47u+7nXt
5PT6F/VKKW92nvK7Be9omx78UVyacPhEFDodMTph5OW4hcBDJ3x+PerufBnn8AQd
gXOgliEgIyn60NCH7aHVS9MwTtGTT2YjGz+tluH1P6JKCCxaaXH/viQs4KoErIUj
fBPgWCSrS60Io16lKwsKM4ld4WzaOonvZz7sauR6j2EfV08vaYFa4czQZugRItqn
DJEzzOj/tm5xqfRCo+qnqRRT1AAWy1bwaqZ+ATN/tZtr4g7W0RRJ/VzNu7wUTSQC
mAApEhExiCpXWI3uxHO9bc5Iqj7q/8XCQkcFRZCSvs8envz9EUj+ehRFqJAtO/NZ
wkDuMQiV6gLI6WNuY26rFtEySeKpYtKizhG02aXYPmSUEIuTEVO8IU1i+SeI1HJB
exPtjMDL3gavfc2BE4HaxldMw6gd8LCGXurhAgge8H/9SaeAE0336KvCDXEjqbHS
Gyt2MpmrEdlyHw+Cho5C5vzdloJ9hzMYoiYcVBw7neae5f3kYh58sHEYS36yQvhe
C072N3iZ7cToGhN4DVrmcDvEM8O2MMy6mpac6kl1aOJ1ZkZYpqggSjMhiOmWNkEm
SOYakg+DolAJzcHgQzdCyrsDhsbPSL1pJpU6cbtUDYkbr/xVURjavFDNP7qDQ+V/
RJ47k5XkF9iMHiCVBi+sDNlDUc0uOKIGfcKN+Z+shTTlvj4bVzj5lkdYTrJGElXk
rueWThWziD3P4/XxINLPqK0nBPrLFUklpn/AQL9a8Vzr2EdjS7l1p8ZDmJzJ9U8Z
mTlhyEXXWH4QjCQte3jYhjiNeCbWfyVWPftZRCs/7qFCI6iL6ANk/szU6+U2CyPy
qIx2M1aewO/cM3ae19RKfIL1dEAPdneA4ZtzkloH8sE3/8isdE/swZtdF3nN80zM
BfW4HPGX7tIWSDsa57NKg3xmqZ7RfQWI43uM6ZQmdeuOAIapfODMyaESemo9STFj
tj0t0nDpQfk6sFfDDQyU9clsyht4UsMgXYyB3PODY6oDXB/tMLtWgQmTJhwws9oh
qhOb+gHdVyBgussFPTR+RGDOhrRN/Yua4qC9PChVVedb+n+vdsjVWKxVuGFFqHbW
gmLUwzmJqFhd5xK7rVw6g4N7ZenrHRTu89O3HAYj+mg6Q8vbVvbcYIkNEQaOqSEi
DMQoX0dhdLeWkwkZfOyE4G0qp9MXr2do2G2RiRBYc26QWEvrDQt63Pt3H4NK1kdH
mBvwKAktLOTr4GdI9dMJra25A73DqdTBMVtCpqOLYf0izbYRoO3ZRW+I/Q9sjpMp
dCtaL1tCRCMHVn/ymkcksvXn7YVzE3b9RgDRAxQ0wuqxo4z/IEo/09eP+NOAQK/N
v3qMSw9pmPftQ/9EXFCVLsG4DlknllzWWYeg0WJLVrCwTA572hLpae8hf9nVaRuQ
rBv0+xU8yrqiv0+LhIpahFNubx03XRrvYnnTLZpjXUs09d4Iu4HSOwk+X8qOCrYZ
vfhozO821R7hRgm6icY9pU6nhAOEfNbkutF3jfo4w0qx04Pqw/ftK15X6HKV0+wE
9g/N7ahpn3d+EVWEzirp9dLgImpSP6mjitV0RRhVJYeUrq5fqSo9M1XxO+/IWL6D
9rzgGWpURWCWp4ueeEsb5Q3eSXqh2YvWvZOCD0k9AXA3+8WC1hXW6GHsA2HTy9ox
mZaW+Gh8Gl+AQTUX0WByCUIv0Z2Dz56u3ci4LmCCeP9+DiVLi/7hRGveSmFJ/7q0
9026vHVwEpv+f4NKVMwtOIHHDP0uWbuGU6RBJPT4dD/jJPuTA/N/JJibEXbGRCVJ
1fSq/QnypKF53UOpeJ174Ppy7Trb9gYIQCXFYGhLxS/M/PviU1/baj+9tAnDmqNf
mnJWVPF/l4Oo6JkoA7A8JZJOkRiRlbMeEoBlj5hyYIWm6OvlZX3bNTiIg2DPcBIy
GjG3amf3J2LzMVC+1U+dTfVhSMWrzrKGsPe7ukL77FyLI8te61wTMtO258puN2Gm
kzQpg4AEx8iIr0xub8+CfR7UCAh5JV+0HpM+ENTGXQreTFDH0y5I4ULnagjZYsKa
nE+XuPUB5Duz3sTIMJoiYxLZxOwzc/u6ExnkiSXtRlJvR84p16ULlwS7XUiYGfMq
MSaglsx6OP7XghcjQcFK3q5sBZPltARvVEmtMyQ+WXN4OE0XfGzptovIXAkbwSLK
vWvCU7hF2SbVozpSFznpIzvIlG7+Diyfe7q/gjO8bJaT32OXNrv8JEtgjvZN2A/E
Z9+ci7fNobS1B/Epc861AG5YrDQWXL2tIeybrt1ndt1XBRUPM9Na5gvjeaWAEKJW
SYswhLH3htRNpgEw/CO8oT28I3jw/idD93jeCPLYFUwAvmd6EbBQ5iGgcHJLn4uh
um90324MOfOk+0IorBC1C3fy5Z8k0zwc/7u5BJkj3LGft7hHbHdgAEiRmShw/dhf
y5x6AjZ0jJoLOPW9kSbmt9jUafrLWCL7JFYQYlypAJfFARFdG/2aZktlEgJ5sqPt
DXjhpL6w5REAHr8uTU/F0lfw7tj9uD5BIub038JVlLmk4vl6Yit8cpT7ZSvAGIZz
QcgX5+zeFkt2oxSGh11+fh8vM8wgTc9OHhAMYUNstmPFoY5khA5348k7ny9P+ZBF
JpkyPLYkGSXyK1SUGtf0kZIYrSksORFjb5EeZGBeVabP6g1jfzy9TB2W6xRsBDhU
CqlxIU+KKs/PdYsfBUieQGi0PoLrFer2iwOiVB9xyUpo+Ur8k6k2rQVB+HyFyODv
bQb4y6Ni8sd/Oo9lJJRRoQCJ5iCb/JnBQeOMrAR4gyd3LdLQzvWWp86keLf+Liy0
f0JlBsua6drAj/eAYT7kfVR9iNWoxXh25UigFjcFYNgLmAUEYltyshQ7cofx332E
BTBHGD3JGKP/7I6F98EXf1uA9B7hxOO4H5bR5D1Zaqnuo04XVvMutCrvdUw20dIh
PRf+ZiBukkoFvcbptiS1t3oVRRZKKKYQdzwQ5Tsz5SJ6S4WbMNdr/CwRcLcyzi32
AFc+9VzJBdmamPui9KxjDN+n2Hw7Tw+tAZgjXuONsIjI56ZPp787JUjhYGrWBBVH
T8mBnxp0+Wz8VCtJFynD0vrMnCBSeA6c/o4sKlSY9owqGkLIEaFSDl+v8nmGrhLa
Jbv8pjfPS2l23lztK1tsddSNV8qPLcbCU4kz3m/26zpzpol1otaqLUNjbFl1F+2V
M34yq9NZt5i7v7Q7pe17svoLNAa5NJpFyBN21Hp3Y4qu1eSw/MHJ/29FOqVbs5zE
7axzVItzNTwBpk8eP/YWXjIMntJ07zDAtDIl4Ble0RF2geUomIwRdBCaUw9aWRaQ
HBvSP1DgxX6HmPakZtEub2gGJTnHbDomfqGyG+oQP5SlUHfMEEJLxU9koNtlpgBC
gguTcCUh5A7lFSBdyOTjJXHq+WvtV2Fwp77xu57NbgPuJWsOtFfmhytEGpPBl81L
eV42UlyVmlcbEYy68oktwHF1TWn8tWOky91K60GTZ3J1l2ov93/7YxTlC0hTDNGi
cGzri/vn+FXLnu7l4+hyX9/dvvEf01QkfNlgU2v2M+1X8dVT0yQBkSLMeY1PmU2H
7JzidfE1pcLqsUThTIHaWlDZcq7oedV/lFsztQQIXhp6Kh+XNoq/UXzRzFQuXPtY
E2doIkUXmVMEGmiXcvFL2afkG96knS2YgGo/9sajOCUY54sgyrZyksXvaR4/cJci
dKW9mTPMl7qA3+t3JQfuccHfUjV4DGPkMIJrJ3S6MnRffNQjYHlKYMcV6PL0VksN
9PpFeVjSGfhqJ5ciasVb+obHa2j6x0xJm1DiZpdwX8O8dbfwxS1FUHsMEf/OMr1s
sa5GIUlHfaEkZ2/XRdDwa5x2Mcl39jC+c/TfX+O6erQNKnjXr/aeTBb/07Kvt/gt
22IEy0wf6B+6mmmFenIdzASARSrR3JFOskynWms+fwhi2FOl7kYapKotxgxxwU/I
Va03ukH8NPhW1iNolL+xX+DVcJzO0QBOsGd2JWJ1wOUyds6WSINEffUFKRl+vnyJ
vWEPjPmxSoYSyqQuPhpUFCtlOIRSTwbNYa5+dpQvGZoAIcaRAMdQGkTJWPPjaVmw
e25/zeGV5kd7RS/JdMD26g+2OeXO252ffD5+q37tOYfQyA8M7DaM/H2InP0/Su/d
ieN/HeNf0USf5B+WSDW7b786OKIWc+GD4E34zzuBYqbdnXs016diAc8v+eyCILfV
Mu0d/03algfbMxIWmhCaT8JKSiO9PO3vJ4tXeu4B8ArIQfpGBCxJpa+w0i31BW8z
3e2pgSGqJjxQD+2Hqm9LTzTqPJWwCV+7ack0z1a/efejFI2a5LBw9y7I2KvsGqjm
+flHyth28J7nWq1ev4yUMs0PsncRkZMEH57d6uwB3ZNrSDHfG4jCWbBJsxd6LL4S
yLAkpd6T/wvgG5VjAXt22LpkhH7Z2oHfvo6/jDbqZiefME/oJ/wzAQeyvWEVrovU
lzla6PQ+4qxPDNFUtRSW9LpghkRRtXsaK8PU3aW+W4I6quGluQjY5x9MBmtxcRvb
cmNOZWh7RW+9lFLaOnvLwhAC+wn9fl9n/JJdkDWEMNSNvWpKnQbuR/98xBith5Fr
nV8mD2AyEzJ3e16KVta0oDavxDU9SxvLkUPlymKj1BPe64nGSzjhvbF78eCL3htl
/9C1qMg1OX6/0aQBuUuf5m6kddJY1pc6gdVfhbDx6d3ZCAFvBuIyp2z/K+Z8WsqZ
pGGJgrMuFYFOg/lrbG71l1IrV6JKVV6nrzKU8pTrrSBNLR/f7Za/CP+tuNaqi4lb
mbIrZrgCpKYyBQ0cpaQePCNcZtrT0XbfEmwAwaZ/0JmD4mMY4l2IN6K70As6BbqD
rkJVZQT8iAG1FIPBqvtIWt95pgtonUVYIBakQsyhCGD2SayDdTnkvwdjKlQ1CFIK
fgs5t81oGbGbCpImaZzIOCK0jNJDKNNG0NiAlhqQFa6xyojJAeGxH/7AZ4rx26Nl
gJ2/70DJNxgrBJcQ2tu1tzQdSlZ1fgXQP98YES1WOCsLd7rTfW3GH7iIVU4q/LRM
Ep6sx7rUz0YHwjZZQoIKJYHEVNPABoClLS1I5Cf7sZJtLugHNsVzYTUTdTR/weW7
jhoDL3JI/BEeJ8wb2KRfkex5lEBxFMUgR9MthYk5lE9PBo75THiY0Xn7S1TJcH2n
HQCyeT5duKRoqKOEiTKbv0g9l2PUYCupCcHk/HLRvf6xLzSv4mruhlOlE0QB670z
7MvfJxdIxv1NYec+eBSykAAN3ujVMjiHxa1UBdlvqFoGzEUmhEjZl2YfBzZXjNmZ
pDckH5mYOJ47Marg5EkVOF5tBwM7jkUjBY160IUxrswzPab7xeQCe1VFPEymhJU6
Vx1gAozy1Hs8UFqKlJUKIuTwC7T20WDATgzMxG2qMwUu3TkqQzYsZjZ7l6c43nne
7LJcr6lssC0rHexMCcbOdOmt/DNlkknh6Cte7ZxXQPhkihY9t8dkNxtSauZ2Xwsd
aAtC10ic62bpkrAFbKJ9Uh/XnZSndljjaFUB+CE5pDNx82iHBA8v3H3GHVy44PDG
rxC/VYvoTERa8TaDGJHT/fOl2pqeMSTYspZjw9G8n39kgtGsH4yvcO8a64Gpry8W
6BRb01D0FTmXDJY77LZe8FwcBJPlhoGtgnZJXa06MIAr17pUZltN0T2QUzyMim/c
x0VUGpLBfrebxl7N53Dg1knaKdtoD3CNHrkqyihVLhfc/Gwn0mItMg2IwHEwTjZP
cNxvXQ0w847nPg94puQds8o4hhOlI4qqWXAZcMhPEAtSRiNh5JTakWAMg3XABBkI
mBUjNy2r+7iWsND0fdmSepvfByfJEgVXPxmJETbJ5CTetv5CMyTVHV11rNIbI8SF
X9gJEVwsy/9pvkt6g6PsJ5Z5aw1ptWmZFqxZdDwOX2oZHOlqVf/hkypZZTQ6PAq+
JVwAOUNCXDG6wcn0/Cc8kmsGx5NUTzENpmKE6RPzh7x3oXbcFjZtCRycA0nrnqko
sFrL0by4lCf4avvoZFZwbusJ6pHA0ybICV6WeHVsZTg+HsKDzNpzDu2h+oRqO6i3
YceeG5A07NYW4EqDtKZEXP1bF14cIR/2RbPpIEMdeHzcMcqntphVOQ5nPS+VtDac
3dnJlGL1B/VYD1qqvlrqI+NEetd8Z1Xw1FwY1YnoACm2WbQwO3O5n3MgDbg3Ykvi
K5/gYrZjHZtZRBXJgp7kw5G4QhVtyo0FQFYWPIwitPhoyjqNccc5gyRQG2q8lO9G
biofiCUVBZODFA50Jg9RL7EJl19MEtrVYB7WC6OdepcId5eg6Kmxmhn5+KhGi2BA
zt8OlXTawn3Qo5yJ8l9COt69zZzJdvJLa9Rm7KbuL0FEfwAvbZICLEJXYKiePn+d
vCYhZTHAAjQWo4PiM8tRPcX6ezwtwkE7bPYXDZq47a1d1gWs5p/RudlgaWh45JPg
rV4G6UoaWKflL7pw1U42WboBPNr///co6xpERHFggtnHFsMBjL72yTf8wrI8VHB2
sHKKigblu+u3Gv5q+G2/dZO2heufV5he5wuuZuEsnqRo2ycBWRwqCbn9PHo9lLhk
dxfpogMcerY1anpafyxVl53Pj/mI6KIangu6W/9nGtRHcNsoAXf1aj6xoe+eWu6j
twdlyza/dwG03VDWuIgaz76bUU+0zbn+4w91OBi/33fPOwP7L0W5MmADKP/+5XDC
d4w5w1HIk9kPtRBR2Zcv6AnpQdmP3e0sivWaDHc6ukqK5dVSsdWxhBTUXGKk5jZ3
W7PV8LmOnbnTwQqaQwQcFPvWDkQOSm9+++qp9a84yUDxpVG9ZYkFtgJjg+BAPyRY
Lt7zb+pRnu8refW1EG9p+DUgD4cXPtFtrekl7Az2dzNwGEvNKrHriOCO6cWFrln0
FkO+UG2VV3X2F4JqyVy4Se3Hbdxwc0L8zlRaDDgFamtew8gGwVUVxPiacU/EFPu1
znwQMZZj8WeN1acVLMocVXpkhhSAo08jZxnNLDxcmC5sETHowwMLwMTHr1VcwKQL
a63m+OYHlIdJ2D1DYHWqrKxm4YcjaVTL2uIN2i57W15rVXySQSMiZ1q2qkWSB/86
uolWoO69Is8H3amcZXx6rof/q/7VxfaACn0g6tUb8ZiUzU33grdzAxcClTBfT1B/
S8IruW7tuL8p0lxI4G1eSdU6vuAbWutnarJ5AqnbGaxPZuHu4Kq78qNo2ywP8Sp+
k73/T235ZtrKQBZhV3dU1UGoX2fRRU1CS/9tvaMwvOjDE8oSmW4Fgu1/axPhkQ1n
aFR+O+6TZBEaLIkEs17VptP1pwIUpLveDCyLXNeKn3kejSIrwdfH7VAjE3Hm+Yjc
FpcnTIusp7SHd2bm0SNiciWEbPmS8AfXTnpxr6Q6f1+8tLvtXlzJNlAwE1nmbNkN
APkCKfINMQt6opPlFKJwTV3Et04SlyOw6YOC8uKBZO9UdcjII35oUvWHtsJJSv78
BRMmXcRoWX8PfN5+3WPgLJzE2Ga/PDvbDB1/UDjHkA4JuutW+ZtAYfwSBVDB5wtQ
6EpacBOHR2QtKWA2p0EDOT4WzdrMgNdBokHGunMhJUxRMoitNKIq8fSq0rPGVtR7
Ft1owx05QYa5wdv1ecFvL7qVS+4eSxYWtIt+G0ENyDe88inBllaEfjUCKN+afBqg
N66FYua/ZldCNofy9TFQBvm6G0eQn6li99+l7d9X2E8ekz7Y4/45r5ViqYTsRrYj
8syT9TSX5Lh5HmgsDoxprwYTile/L87qg+ZCTftXOit5pQYuPfxdTMJc96tahpUJ
cWYinZyd9sch+YSrpIu5t6P66EubfmNjLa5hwPTyReKKNKl0TfhT7+oGznyIsG3o
rPmE05XivTk241NXWYtilRk5t5np19xaNKoLiA+XqAuHw3jF3i2BAE2ir5vFZnll
9KMhPqBtsze7PMR0pLg1gbhN6U3k3L9nd2zlX5D3YoBqO3TT56vCby/wMPmfzkbO
vxGIA0Qh9FjJMruQ1t+tX1/fSaonJ+acIub0dF2SjZGGbxrIEzOrCEGTGdo3LscD
Uw0YH+X42cwAKR8ESDSgnmEFpT4bhnpK26bOQtM+uuy+zresiI+PYgzNSWyeDpam
tPNwzJy7rfcKLg+6/FK0orLoCirbdFziBTgF4d9MDTLoUzsvjKWKAjBbmK/dRLc4
V1LyFnvEykwnXfCan7zobEZAqz5/3YTJEsvZeqyuNaGX4TMY2p01LUXbDquPH83f
qG5GBzMwflWcqeqBmEJIw+eXrs+0xgYmkjUK7ZqvgwerTlOFE9DwDXliVUSg/Ndg
7qMQJVAxR8++es48srt4//MUT4SPbV/er6M0y57IbKPII+1q6Jkwj0hmabZC7WIj
MTcWFmTkwxDx6kaY06eoF/R8v6b8V/XhDo+DOJoOHgO5nvtRwp594fuEp72dWw5j
3d/vckkjt/E9Ap9nwU+trBC/aafZ1eolmkgGc0TLnanGR2Q3DVWqzmj4W7NnKyRA
GJ+J40s/WkO2LaiPURjnoCsc9gX281dIECByIJqtd9vv5dXQkf3kDIda9VXuvos3
3LfAz/74DlrvhGEPcnFIDh46zAtdwsbo2ooBjHmwDrSi70EtdOeHwn4UW01Jaw3h
/ZKNQ8TuKiLjoJTaQIVJvQ+7/uckMpPvmx8zElIF62CVwI16ZE6tpluu/UcaW3hy
n2HkkSSsCzJXPqSN8FnSKQVCuOYkUmpqffdDHZuu+wVEkrkA1dOrVlvzMFFYcrrM
ykmvvIze7eBHdBCA2TIrbFFFyouOA7JXY5jFVWNnkgLMpaBL+Skz3Bdljc+sp/VS
MoCeLmDc5PPEfILpjAJDtGOWV7BQQgNnnjyGStiXVczSLSJTFkRYX6PNxo8+zI3p
hzPMIhKY4AcXUr/zaRA8tmCEBpOYT3vwAOMUX73cQ9F6WuLW6BBAn3O9qJfe2X+2
56d9GUlvHEcOsf+KiE6b9JAmn8cWng05tt5VUV9M6mnnSgH7FdfA/Hc1gYU7+TKk
hHb7XdxRnB6eZgzAnE3LRVMa1hJbFQZrBdPGIm1+j79yICf5QSaEYA43wp3wAlXW
ZUERjQL6O1TDgS3eEFuv0bxLFGkS38HQG9eLg4vedYwK6DNvYG40sFN6g2eeHhTt
HtnmId6s2plrqFU91ub3t1FQLclKmS4yNrK7pgIEQ8/tTi/z97FChm1YnAl3/RGl
aqN/K4CMdAQrhmenuRlP7P7hI09hBAsSeHXrRIM/jsPgymDtwnGpnzCAPeZM7mhr
jOiNBRT7dceGA9A72nRaFFYU+z3G0TNEPUKOZefvyiC33wU/hCCdrw6nlk9sXJqc
EtweOJaupE5qaMpg5H27ho7RnzOUrbCjEhzr3sXO2nmN9/CAhZicy593kPcBcLoz
ITlXZSTrgTi8uPLKJJCKGYUj0bxf/8vSE/1ZtEMOS35hXp+VsGeLUlEpwXyzyw5F
WVrIK0SYuVrNzNj52PZ8okVcIDffctKuj5it2ybpdyLvnmEYAapHOMvtKCgGS2HQ
Pcy8V1xwLEJQhJAS+Bc+b0ubX0z4vK/rd681hglyvw4c7tbTJ5I4PQGqR9VTySPC
34+eAlh5adSz50kc2T7jU8p7Lnq3RyBPd43ZsqmGC8cs1WXWJ5gJRswW492jfAzR
r3R+bQawXV/MJ/1xg+NBdw9rH2MdHJkJApyXKBnmUSTvsyv/F4KTLlbFCdwEFvX2
fXP7cFmkfdCZMX6r+kvwPS2pDZA0PGt7ngoVTUUX6h4qHIFes1p72HFczNMeg8Tt
jTz6iDK7Oc9kAWH1bXwNYhQvmL+2TmHdYLmqEEbpqyCOi54NKjlCJhYQ0NV0Cix8
NRqSKRB7TGiA6GLtq/kKaQQdAvOYsNbsU/0rZByWMzSoQYFfbjvKdGbS5Tddmk+B
Faw2Vaw2rc3a9iNZUu90j7cgqFQQLzqVRezg7/Mg7zee5neSV6iXt9/KkGkgokU9
2j6zOlHABU2WC9PhtuX3C+ICkLotcsZETN1u1DCty3PTPSE9qJ5NQ0/vc1q3osoA
lI55MsRCR8V/V3oawC6IX8zs7qgZsCBwo5JfQwxJb3IvZwWy9AV9qEWruOeBC2mr
XPM4F1Bu65sTWfW34RqeVXBOlBx5S+XA8mx1QSswyP6tKMMgaQFhIUIubieqg+Px
/JSgsiZT29ocQmIsg0+8HN+XFznxiDpfGmgSFT7ABAJ0E2qq6L3tyg6ZclW/ekCH
lxp6ta43nvGq0HnS6zsJ4DPTy3vwauyItJOQ8kl6ZM+Y3l3r8LosWmHai16ttH0V
9ZNZoT+FbV0T+zi8lgMu3YZ68wbwn/HhRCMh9ttnjw6ZHmWaDEihEjwbNjvbso/c
zUBjN2Fvra4QB/wJYmQt34/R7NIGD38xa4hddBCQtV+sV0edEKp1nSKuyOYiuKUV
xir5kH18iWMYgU4MrWF4SaSD4CWVL3jk3RidFTO6UTw61sj6KK1a1PGDa4gd1Qh3
DBBDm4ynItmQaMCvSxns3Spf5IBqG/2yAH2AhbzjmsZbu0jOlkdnKkV54edtdFwO
O3ORClC5OF/LqUOAlyk+YSvUwWUZY4ycSdYb7zzMNZnFyM8zFxH7D4S4d/fqlHfb
AJUBQblQV7qCIK6IIM6qeA0FfeMTPmCxuoQS0WkqCBfOwjyMAj/GSdvgk/UjGf89
i5ldLFC4OtxbOOLagOns1f6PUCJr6wGSyxRTRvK8+Mdo2nvBgU77IqDE7zk9ZlhH
Hk+byLCjcatGYxWpDINc4LIVe2LN1dR+XvtAZSQr6ZdY+SbHvecX7tIE2omJo5ak
Wj/ANNyS+XN2nCmcH9u9SQCOiIvOzdRd1sJlMEz7+uJmVNahRE1f3mYyPn8JirB8
E+oQA/WuHJWzFWBgQfl66YJfRNAIf/odqz8aHJ5wYn0PhxypfTN0qjz/3RzBL7lc
KkhTEXpwIcRSFs+L3qfwZdTBCrcd33D1cg6Mtrs5Td/wxdrg2WM/i395gnA3D2SY
XjpJ4jZrFHn4QliVOg9MyYhbuesPjuslsmzd35nJqh74y63o53JHUL5POCIng2cj
XAGorOhTYluAR3rKUie2WRjo5tJ/SVCpwkJ5SSoiygOllHmtdze2N6ERK7x1X9+2
aVDH/zYXeU/1BEYpiOVnlHvWkiSGXjacE254VWpCanJJwhF+apcnZxzakxs+B6jC
zJb4beKUaUwcShaayuCUFJKaqKvqhenAr9dHGLrifRr6afnXJfJ9inhDIhBwj/k9
QWJ9oJ1BXccfYMU2vKTpHlsdY4cIPqCzTFWZwJrCETaDdYk30o0P+TWc0LFRGu5B
R1xF/eSClSRfTWuqcxmuZjMzoCYihZlf6lU2Aakbha/Jgh6gGKIe2gvYBq2O1iRz
JqI75aVunA+50tjsb1ro0sYcXQPa2FXFRrgGJ0qEflRJJmyT95LSqzu7dZJHE8X2
cBF1HaSi4yynIIJDP8Dcj0FJZFni9HqdoV5KbwMY+8glYVOZa2Huluua7/EKKp52
LdwUQDZx/s6A+34Wvx5aCfSffCR+bEoRju4/hETwqKOHW50UIDa9M6B3W6PiP0+c
Qc9Ms3JkBFmLdRte6vn5YzH0PfhQ24sm0hKJvzFn3iSY+zvVNEmIeYVi9jkdvYoP
eNJm+1n60a/8bVupKh2pCUo5zjvz1NS7EyAdKHHmLoM/YRLYoAKGQrzJkFMre1TT
fvo1HVFzCCLCmUj39BnQQSykCS9mq4OCAdLoVBRk5tYUMEv9XHVH5KeAl+3UH1py
Y2NwRTeXMox/q5uvEy3M9kShpsPb2e3UZ33HKUDy55BQeBKYhwNVTqdbb4YQzxJh
iZbr63+tIaZrrbI5OHc8aJzxl6XxdmNtEFFvesJxjMRzcfGZF5j9b3vEyTcPKipv
uuoqbQNkj9b8+40rYUrITgJVj15OLuXh/7fNZqcF7CvM8Gsyq4BHLo6XZQAE4CPa
4/6XAXhXGdC+YsCZiYvIpT69cqt1wbYwHXWKUGqSMP3I7prPLLklZvJ5c6hMSob5
ikn86EDzx0ve9j2E9xK1cDtV/OU7EriQRV3qbOs7isj5yjWbNf2BTS766KqjE99T
tb5/OeRaEcqlFdp/xcRAskEqHY2+y023jiSi8j5y/ye4KcdQUd8hiej/RN/Ltvn+
eeHqmAhuja7Pt8fsw7MrH3STRFVa/7MNgtmR28Eh1aBVFFBch1io/ISnjZfDg9sG
KJKchuYZ3KiQmSMnQJX5WegCUDZ7+WdrM2yxHueWb8epXFHkwQQq6z/Sz4p5ZxNn
qoHWGo7sJ+XkmNesPyht66ROoFC3AzGBWHEI92zrpZjNEMWm1sIGlJi5J8qw9USD
0iCy6ejFR1JkVKdxgXdaP0ze1Jf4QWHVhTvSVwbIfkrosi9wv5gMmsnLq8M5ftJI
xyoiSqHKBP8uOGwTHtdQKswF8iRxbA9S40OIRYA9+VqkpXAblSjQPQcWkP5PDMoh
3JHn6q0WqLZbphU8ce6gxHML8/CIXnjyL4fR253iyLrnL6he5BINFQVY/doARlUZ
903rTVxoriyQ+MSQo47Xz08Y1wONRJlEQCzAy64NfCj49cRv0FwCn4QGBHnWKLP0
XupELPLUrvv30uhp5akbPCt7lkUkx5PQeEgqUMr05yBW3x7B7xYwxNmproyihQHv
QBU81CH5OYswtreOhx/G4Ec8iB6rRDcgZyAImswp6dsTXO4j6FtC3Xab2wiN4Sfe
1XHjz9hXe5wQPae/lMWXqw+kvdA3VaWd4S8mRoXurCWuizgY2hN2AvFXOYhesePp
I9y0jdSKlVJ5oqXDJ02yDRLle0mOlRWxC6TznQ7+zl+CAtyGiDpGyz/UOe55faGE
wI4QEoc1lTmQg/EZSp0dfv55oEqfvRZ18deo0BhV7LgkKUEAnPARL5H5HAqss4TK
1Rj59w/6V2Wa+/GgC61XJDrShwBp646yLxcddC0zquvR0VVjYIpZ3JeaZAfJBicy
IqP834gdwRKuqONXgvOiwrkbJ2OoMxvdOuijrTWQsgeUYFMOy32Y4K9FVLBGR9bM
0xyPYwKfA+yKRezXKcolxH1q6FXJeXMYg0OCa2r+4PLTcISDprz2sd7TJ4zkrcVM
dqw/w4zuWANqapp8gy8iN0ZtgC8AoHcf6BX39cUdUDqhap/g6b/7vZYiFLVHZzzO
czmWPEVenjjqbbvIwNXSNdhiqXmsto/a4KFKFHB8WfnFuwhGTFiUUPd5lL3KibOP
uf0PsMTTHMdxJidju+7thqXtIMiu/slhessM6bC367CTdSQp+qIzDP65bLKgoqcc
/A6EuoSVvQ/jU/8uv/wQ02bxCIGq4nNLbO+siizGTvAzBle/CzYsf4pQKyYH1hy5
RvmAvdL9FFC8FBdTnsbZ2Xy6DYmUuPBUKGXE1KILTxnWlq9dZR1eqALX9vHlqepP
pagsHbWA28QhE7Jdm1weeSYlzuEl0cXJOwa1lRBBiwc1llLfZLW7KNDyLJzSUjeC
k6hLqpfleFEXIThhW5IWW9PYf8DTmjA3orggKWzuSNel1rDeHrQOT+435bGZO5Db
S3JD/OSfqIPv6Hd3ppUbFqgwAT22NR53NguHgPkVV1RIxAQ5RCB6DxKw1GQiFMLG
`pragma protect end_protected
