// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:53 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gPrmj8qTH/+xCGzIMYS+FwJZLdKq+Tax1mEXq+K66aBD//DKYLme54hRMciXxVGO
aWJD8FbYXIqZ3UEDMcDAz0OuQrr7euizYNxKKw18Mw3zsRDNW21jc2Qst1JuVyLK
NRaolReBkkmFkspyfT/0v6estkMsORIrQmoOIOsiR2c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20144)
TitM6h7kz/p7eW122CO9BFREO6JO9PVZuxyb+HIxbObVCk65S8q44bFn1JxyN+c1
3vI00C8EOR+pgkNvDWe1+JO1KjvIIs89cb9Vt1inFM0zYp/pLrbzw1QxJ+KCNZ9l
ivPHNX7wspYf0fZ/FotQPAN508qSls2VlV4ey1l0aiTMu2v05mM9LeWsbZI1Uc4S
Lpfqng+9+539Pm/3kLW1yn/40EJ+Ba3s2zgHzq8D+LlNZtrG7NLRdvmqlmN9SohN
xtaLtKZV6LWrBPBBLc94MzXEUIGvW6qgrL0BTlV5jLxlgutdtFmJD2eZsT9RnI0p
f1bug53IluhVpsM1dgibzXxxXHNhwOXVBZdAutGbab3FUKn0sjEtpqTQKTT9pcpJ
CIGxJr8Z4yX3BNG9NsYTVX/BBbZJYR3KZ1XLu60b4bj0wPEIuyw7D5l7cvU0lU48
sWr4BeS/5+cJO5gTEv0V87o89tPrhcSt3kFJOoUeJu0AdgGpEafVlbeKDLAlLRia
okXoLUrYkvJrbzLSutx2RHdJxzL4s0pmj/MK4oq9/eZfRA3uakDBkQHAlz8DQn0T
E6fAiy/KWCc1Bq0vGl7CzoacjPFV6YyAICen0nTjxTrGL/pvfuniMPNKZlUtLHQg
DhABf8UAtxvfaRgVWLv5O8CkoMj2jT6YKEmMUqAVE9Ni0YriBoCLh7EIbp/UlWun
x7ru6nfzcV+cWP5r3P+F5WSAlgJzaG5e2w/eLfO1681M3xKWI35dOZ2W50GVv5GZ
6Uq2m3uZ1YQxW0QQct8rdzhsZZFUnkwCgzto5usNLbIlmP0Yq/KTVbgcl7JrtOU9
3qaVJIu+KwGWjQh5XTUWQD9fu24+jRDO+ayPMJtq/nKHtKHQnXDt4UKkKqkhmdRk
1bfj3HAyojjiv1qcM/HWDDDnaVu2hTXg+rHXSwEawrrci3LGrnw8qJ4dO9ftyCDh
HVDL/eyHTLLhK4ZSDvCjlu8+5KoSq5Qc7UNk9R1A8SAWqZ7EvOm7GBwAj1edYIm8
pn7WP0OFdTNVk3mjVIqlngpsuyJ7+oPlD7kywQu8lLn5nb4Lqnz/jTBh8BgTmyLk
Eh/09X51wxZao+54/tTfrwFCr8+E0eB5zSclRof8MDCleYYcnPm1cqN9ys2wFJHC
id7kbsgMrE3SLnE/qL4snJhraMjGZ6+rTptl6FDEGMd/pTbehv3CvM6gU9a+ubD2
/KB/bVOWQnqnaJsqs90E4q+J+D5ZdomU8A2j/pX6Pib2ndc3a5IHWWPpfvbFxQ+3
grU4IgnKNjTVx16P7NUbNCHKiDC9JWhhv5GTKowV3bcAsQch9j+eBWYba//N5Esd
z6xuVswwdiRHftc/o7HQ2tSNqS0k67AJqwC0cuX7UUwvzcN63F69mkv+oCq27ZBw
vGAVsWmXBCxlf64RdpeWdJaFl6oUIayZqt7IVBioAL2FIXDtt4phxjJUw9gwSfXr
b4wSKPXqRTyFSYdKn/0Wf8kMgZ1+XLAeTVVPer1gFaaFvofoS/utouwAgllf7WJa
yMT/Zd/9qR08Q3NSREQS/Yk+pKkrY5+EcZF4WoFABrochKvju/nKWN7kuirnMu3R
dS2VyNT1xZZVadgxulKpxHVYFoXrvdxYqqEbDrP8jhidPjPoWbROJ9KC4kjVcXpy
2YVbmBME6ea0NwQxGuylZEkhk/W3WPOPyUze8ZaH7HE7zMJdu6YC9Pyz9ZbtJx7a
5pibfvWaHerPYGD1cWbmEP0RWUM5ZT8f8qm8BP9SpYE+nKu6jDxSGopE2wTEofPO
ZyHIPaYWjFzqAr6yuBWKfhRymqxZNa9TUGqOTfQzRgdnxpHUBqg6llndn0qSZHg8
5ckWnHSA2Fr8DslT3l1fESz/dNPvdXdcAPX3tk5G2lb0IjfTYTvnJDuIBmK/+fz2
N4iB11VUYnprUtY/CFviT4i0gW39wNKZRZMBFgt320As7tllIUC0v9uQCbawgxzY
7IGoKCdp3t5P0jABsCNGdyeGvBibMIj7JWhNhzjFs9Vsld+7APvlFK5xrvaSd56o
p1+svLCmWuv5j15JpA951ah+q2HRNBlD875SNF2dq/C27rmeuruCGbCaC7pFlicL
HMMz2+iZL79AVzfUFtV4IKBEHWO5poizMzdRm+pQ4ra/whba2pjza0ElQUXe5zCx
Rjw1O6kNEMlmWjeF+sosmJZdieqIpIxgb3lKScEUMYGPF8MqbrBtl0uVsOHB246i
MSd6cnP4ng9RKB40ACPG6yWjEESKziMvPbZArUjH/pqh4rfV99mPLmE5ungF49xc
/uBTMgyDjTfhKtNx4jP4IX5jWtkN9pfEnR1mVGTji6HvE9RUYFffcZKcar0C3v/d
pSLm9c+3CR68Qqbx09fEEJdJR+Z3JqtNO4XNSI8CgOcClr6WC2lGiQ9hZqpI95+T
NWTwvnS6eGJs/gEfzK/tXyHd77Dg8VV3nZ0TyypgKfu0MhLZm/gzcL5nnZZpwde1
nRG4JBSm3VALsAissCoHqrIH6TJ5mLR1ANJuhIOWT5DY5dFwIoDz2lMkBnlICzTw
Wdh+DAFnv7fb6HoYaWC2/yWRVFzWcQ04Dm/XSeUKu4lXFHA4mAlb/iMO6exhdHUU
dVOk6ztzomI3ff7nmLsdFfyvTmapjyxAOBh4/XYIHMrQJ2NC04OtR3lFXOZAHzh8
sr4kql3nkMvIQ2LBLW5rE51st7jXRA3xqYy2JwMzKd+LpeknfwCW78Q/Yl5r9+Sr
t8CnqStcszJEP3QJl2rXnfuvr3LNMLQ3rX9kCjcE03/aQo6//+ico/cElCAZwgWd
vPGF18JqSIoIi8PlCawL7rhDCuqmLoWHbOBHyU1RBgjD8kgWOTeacrWk7w+BdlCK
DJNLX9K0hjwVaUl+6cUWOs0z6F/PWPEeEUjqDDfVx3EJsiHZfAn2c2MXoFf+9ZD0
/m47ZdAXM+gg69SKRtEulo/SXmjYtxuYnKaPihtmZjd/+ajetdwL6ZHt6Zc3yi1r
9sqFLHMzgs+mP0KcMAl7GCQhYrHKmRvuVXvHIZPLmpdtfzEp3N+8+yzrGWCMan2v
6yQ1xgRgPkVdomNPtqgU4vBFo3vOSzx/KLZGkeL1kolYMVnMdiJkcjR+s6ml/TAu
WOCNOF/YUT1mvqP5/gOcB0ii+DkhSddpr3J+mxtJDwRgeOlOnLuxoUTkOiR62DEO
0w2ItYD9E2e0WVj50NIt1dy9UVbsATqzI0k9WOTvTYPZJO8VGGjEoeSxIowqEpQi
TESVeycsHTny3dwTC5nXiGLJHcPg7LUJSBszMIxoCB87IIu16zQ+Bx2fDgDaL3oj
KX98Zgn6jlgjRyfpj47KpHUPzg7jf4HaDuiNb9soVfXoiFEWgI7im/64biJARq5j
CsTTHrXRdPjrVEmfx9YGMLTBUYjx5BwtUIPUlGzikQJ8Db4DcxkcqiIJ/nMhFW64
NBx6vC1Ppbm7Mko5ja+vRB2jOTbJAEJM9xlbxvLUA/7MKpSyWQrf6yjIOq2dqPWW
UNTpgwWxJ10HfvHhdRD0R60E3h5aYB90E/+TmlJvB0rXil6BlO/ThM565/iU15RB
amJoeYKXNaTqPUlDOqRw/UdYP12hBMaBGTnTepYPyxdDh0s0+wKxXZpMfp7gNFu+
rBLnSZxIkkt6JjevdL/B+N5ZtpnkYnzio+qARezDDs13uu1mBQQYeSO7lsl+EXhb
4w3x37RktVvkr2V7nhb7TANaC6bV9WCcusxLvY6q2twQCTibFKd3UyIOCv3qHwmR
XqYZ7jfnnmBwFlb2wUqpf5hQws7jrlzcv5IB7yTKFEaJWiatOuZcqq7Xl5EBR0pi
C+JpZ6HQY/oqL2rbfwmjK8JwAPzusRSheSB9/5/DIZPDzeBflP54nEMomQf0bNcS
cfoQJ4xCX/zRmuf6NLJP4DAtI2h84hKh27S8KPN0IsdMW7x/Rj2rX2EMqBltwpCq
Iu41+5Z7YRJWtErOGLu8p5YsmpegQApywZWqW0D3nH3iT9KmHZM7KGfYm/BNFTns
08436eOyN3KcgOmAAc/FxG37M3/1AGeM1E4INI2zmr1cVLYYcy5/bfSSTcVngDuB
eBblQZNlq9TWqJ56txIoYDVNleLK+zvcKWMe8TNP6mMunvWv54taEqYCKWlUmjhl
0eyXQvWoU+Cdt4HKSpf+NJVJRKGPdxRtKfYCVV4pAz/ihWeQTClLN450NWVMvamY
B4HOV6cs5++3+NP3fOGx4NLlxl1pF+PSR+8SLKR8K+x2Rrm340ROlGp2TVt6rL+r
uFjhLbno4kL5iOwpqyaXplY1atNIsnz+F3mwCpU+1DwvWEJFK4Zzmg+ntS03W0od
iMl2jHikS3C1Pgh/dmjAdFvwY7TZ+O9qpKDd7B4n0GxJW45stxRNmoYxB5OWqj28
5Z05QhI9pl0AeOZDEspOhsMaDMIfksudfAGBl5JVDvxFADyx9BFm9VYvaSScfiWb
gp0gEJwYxeJisI4kOFMlDxcs2hCxfjN4eXM0Bb8FbY4G9bsn/cL0cNvS5yiGPYqf
nn6hI5kzRzZCMJIFTSamSq/K4gIgiI1FlxmMaucNeayvsYZfi89oDnjmCzEiHeDX
+l/kxIAeYdsxDLGYQgJWAO2t5gnGE6HV2H+uvlic9/73aJrRnAt2R6qkP9MAr1VC
59w7M3ILLJhFiGAtZNvwEiFgCWz2A/Lnzu0ag5QDpka3kgrp6lqExqEopwAuSvEX
EhKKQJRjdYt7gJFrCVPXM7qq38VOBoXDd+w28TGN1JUfOIjBt5mqTjEM1Xa1TqSF
v+vp+p/QJXeKFPo0ipT5tp2moNigYfIHbxZj+NTV5keumsV4yB4UlAkL9/BYcURQ
9W6GXMJwyYvqBj+pFkTDanthkhUxys9pBk2llTfGFpPKvIEpx3TOsgCLPAhRUhea
w/DdWL/HYCGgPYdJ7Du/uZ4qquKFVSibL6oWawh0bKD8KlnQ+m6c5hn/fERUg6D+
Yu5euKm4D5YUoVJadTQC/eYxEP3c+9nAsmpFv7i/9CkNQVi4oiKzlUdAnLOCef78
+fWvsAUECt7ODIEWiXIBCggZH/q2vBC5IFBBMbqa9vQjCc/GurvhtEwOJYkqspzj
/dZido6mPaMtzHGBr1vrgBFdBaCfa58GC8gG6btCOuM3SZ+LbkPXREaNh9vt6Hvb
gW0bQwkgZGQkG6UL9Yo6DwxbQLYcGVf98vhF8X/N6IMO49JMKJ1li5j2vwTari1s
EYW6IL2N0HbmTQXeGR4Ug2eVpQ8HsQ2d6jPOAEt/jPlGHDnJxST4Zd06p0+tDqF5
X0vJNlxmWaqD6dDXivksDTRj2yElnamM5kht6k4nEl7ej3aGKWHEWfwEqnA36tLC
lb6dXrJNJf6ciLTcdAYsIMswm2t/UdSJ2N7wApL4f+h6XGcTkHzJ3V7qS8mAbZad
n2fsUVztMTAauoyuel1kDiQIqZcTcDs2yWRapZkRK8kkqTP9cMX0zTa1kXV4nH++
PZ2T/+HooQyoubFK1X6F02bMnmhOKIjHFSaX497dQ1mBY6YKJOGj/1uH5onFW6qe
lHEIwg09wkfWeVEePLgbqo427hex88PGCzHr21bnHoiu/Ho6F2A+d0cbrRe+C4na
7H7gkm6/Wb8WUi+91VikgM8IxoUpNuYseQRK5G4EfLJezpGKO9NmgRTX0SCjrRWK
+h1yXlsAOtJunLEESWfkGlftPHy2Jca+CpBd4PseAwM+JjIzEjCRAjajmiKhQ/I4
361xu1nEnPkIkpsrINPLPMjYUqgAfndgHnsNbIj8eLegSu3QF9MnU4iuvitkBtTR
RKW+tjdfLQ6D/bpgkqq73i8RJV86ZumWvp05B+JiXwsp3duiB02zN2FHVnAWocGc
EyQB9pfSVewrqp5hX4kI1LUYaGEJTgAFeH4z1u1JbzfBC44Lzyx6RxonZ0ehRQfB
6lhHqT+FQlysJUTwKFu2FfkYqnzgi0+NCn1XI3jCAZH/E0GVigC+1l08jXpQqzO4
8vQqOAheuPjcjdqIXMzuFtfOUsZmGn8i6Oq4qnDRB8yLuFMAPVc8FfxI+mbo5rVq
A4FbAGhhHMQH+gCuNcPB4B6udPseMOCnUfITfoGW2HSq/+qOzuG/HUN0h87TU80p
3+KCLRQGmRT6ee675rX8XjqSNS6Q2/5kjxJr3B5OqcB2IKaiWj0ygaOREdCyBQ1T
xfxc4fuAmyuYyMVXixqrBVC4KAaQlOtaqsUtSvEXeSM06svszsq6Z6lVQpS5QtMs
kiZBnM+HG4nPUEXcCbKqHL3LPOsnGM36v+zJyE3b+Pn9mf2j/MQ5dS0WrwjBcBX4
hqkMC2iA/j5qX+VVI0t5Y/sUtmbGxD52YeJ2euVMrKd7S4wbYZREoSGeDshg8j8l
C9IRyJEWVIugyC4iQJACXBoqoi3MkXOsaRepJm+zezEfT0IJbG3iTwGoma/if8FB
+PZJStnEFMBxUyi18mlw3gtm3w7URWA3j6LhxZoki3KHcpHEOxwnQTGdhd4lqX2h
IxAUweTO07njtk+e1mq8k5Fscb0aVu0pXRZJp4iT6rVWRUOJR4RUOyFHg+j64dfu
dQykmGqNo++PD8q27y4WUwtrROinVfprdHWq11hz/HVlXPXrU5twCsGmhZEGPrAd
LFmtuhm0wXyuiJ8SIsoK0CmtffcrxlNp/kRGRw6sQMnBfGE2rsClMaqaAIgkYq8O
ACDT4aQJenQCCe8fG6NL9meBKf0BSIzNrvfQUiuhr3hGZKzdRCov7jATwUf+frD+
XGMRLqZvBLajgVBxjYQrA2p5Oz+qqeI1+0kKZKGzTSc/ipq4ME1LspZHAT3gMETG
tDLx4c47Tfwur3H4mfIKXN91H16MqJMloSWEFK5LSDziO6v/KTpJtmLfzq8gVl9u
NtK0UGWEi4UdEUUWjXcSFln8BWUovNn2KWSks+GPrE17QWfkLnB8nOR3rnVF2uga
0IwGyykBiQo9gII41/OsY6GiQjqWjQvBo6IoGGTCyYrSZEu55ZCyp1hu8L2b9ouW
N7hRBDQ2CkCU5L0l2lDKVOh1Z6QCSNDo0Sai9kTnzRZJnvUGxLdzlA3Y6fq5W83L
IAf1Qugja5CXVlPjsJIpbKBDrKGgzG307jcXtWf81hSVvnLL1GD2myNANbjgAGx2
PptGuALQrr+X8D4D37fH3ccSsCmmTaje7vbG/4DwN/lf27sFt+IrO0FL2lGLmmo3
a90fMTqxc0Igzg66Y01au6uSvUCTYKpXEifsdfAlqXfD1b9RMyKxqYips4MIglIq
j5x1qjSCwlYOMHM+YMgkB0XEmxT1gaSa0OsFJcKZehM3j6hi0mUt2mOFm8bebfMO
yS6W4s9CUz7K81PEiDGcMFbUOpFrRMqesuWUh7APWwEpHzyYASif79dbWPc9+oTc
qKSNIw893R39TzjYg27RYAO09fz2Go7A4RayOvrEtcWjkvLeOUs40kcWfvik2lO3
KD4vqCpXhSz26heYXBoj2N0M5mukYpr1XvrnRkVFw5Et1sFNhdH9br39VY82T3JO
cKYsRpdKwAyS9JP5TSGC8PNx9zO/KoPY64WuUBkCdvNJdT1E13gR1tcTSOKzzvtg
qJMoNcxxLrzO0f61PQ2bas0hNmebUFyawTnWk8IdW4cR7sZe+b8KQZ/aQfJGOqTF
gTn9POsN4/h9q7DR2+NWMn9FwHMMK0uifRscjbbCqjYKVe0IuhfyER+qDOzBngzI
6YrHkxO5//o6mutmeiBSWwHoEmKUGqZvn08EjvNmG0H+Xc9BPHh/hxUP9EuKN63M
yCxncNQnf5A93q4rPXbQlt1RyCzFvWq/wgbbQ3QlZ/HTjSxRZnjFe1bOsMvyvaLf
EzRJfEVbtZoHQYyrdzI8jgHikQbMnR5HIKEAELyURmiEH/8EPypwFx11LIa4+8eP
U0bqHULTk0Hq8BQG6DjcrPoHMLXwVOyrS4Ryg54e2hc6/grrvvfSc86+XA5CWOc5
ZxmGjnWG6zF5K71bGsCSamEkZAvlyXyFsBLWFNwICsvBF6GAKLleN7Fxis1uAOB3
ThvN960LjeyZjubiXGhJj67WKVxAf6/Fr0/fQulQ9b2I2eCi80w7Wh370gqtQyp7
calAG7QUhrd/Dj+J/obxtTweaCvjvFRMnftoGjT6LbTSb3oSHExRhtBGxnEGR8kq
EhFiz0Dy361PvgBI1C6XyZaL0gJXKpinnHTBjG6lzi6IRSdVweCAigWyezaQZS45
IUsjno++PO+P81DudpatNUneO9zW+n5CCInpJj825x6mGV+HA9py3SuU264IEfUj
amn3+cI84dQcF8aQtCf0cSndTBpb6kOka3YnjRYXnWD3NTLzYziNBoL+qORRr0gs
x3JVmPxPeC9qRyhByAo8e5F5ZKuMIDFcH0bH3VUgUfxmPp4MLvz9dWOTtZIusUIg
dw4EMULahEOlQs4AsIC3djo/6kL+9jlB4USxknHNygyjCylMM05emAdsgYOtjuKW
8wM4W+Ex2fnrhnbi0VBJ/mQZJweC2Jk7M+5eC7Eaulr4vhRB10uPm8O5tef+gZYi
iII14nLuum2QuggvwOAKHqlQ2BMEe+4mQ+7ghX9aI1qvLHivnWNuPA6XE6O95VYd
wKApuikyzyXaMnDBOPo4NFKxgZwHkk3X03mI83isoKBxOGdE8SOsXQWmbMYuZ8fy
mwoirgYlzStWVK3wfrZmXCGwxOtXV7CrExbL6LNmq8WGJJNQRvTvbEsv8/X4lUGK
AY6ZVSg/prIaP5XWsOoyHFn5yOM5JBPEGlF/Q3OR/2nnGNniaYo+igauGYsDckHM
IAFt2KUuamTOVPjU6H6jTOSYQgylpHgfSbCXXManx9a7+Yi9O15iYVnGHcYH58/J
pU/chN4utyZmlSlzlEjaBBnPr8PYBKHrLoqI5rVBqzMpdWd96lDQHVo3WjkFbafj
QlAfytkX08b/faVkjWqkOgcBbivBaD14gxe+GM5RVoQ6GkHmXrV0uGbjlq8f0dDy
1/01hFjQ9x5QmbgCZqekqcqWBPL9dnUV3tOST8FEA7xmj/UVm7/H1V8mdU+Qmh/D
ynvgeAZRpdosDYMOGoMT6hNYpsKTRF9mrpffkaVXfGET5W206+/NPZR050Ym4e7j
Mu7jVNlMjnf5F1ltlYRs02kHUVE7Em8typxZz/fx5IciN62LsObqURXkz5KkK8jk
5oEHUg9AvDIBqHkqxAhX6uVZV7KiHG2dXKMGku8nxDd9fsGSqmyG2hyAYHoO4qA5
DeXtOAOWN+eAuxIbNno40Nb6+jeB9cvW7ihXDezOL1lUZBpFMtNa6+L4+OG/yvKS
bb8kkAzvS7X/vM2j1Wam50RXqMynfVYhWkq4qmYgaJx2Rj9ihZiMyknIA7a2NaDH
gUINJdrmbkcPcmZhVD6kxVlaOodiqZuSZUNqodyGoAREPlYN7DtHzW/EbwMBmcun
EWbrpfzvXi7ttop/3udZVSC3fZtpq7b4Pao9jNMS4K/m0EOwfqqV+BxkOdfbf//n
sUBPewPP8rFvJBKYy2/qyH8miyCJhRxJuInwnlD7m4gQQ7XC10P7GDs26HIaR9hT
B8P0t3HQOSDTCUAAVNYaqAxjSxAMAXXMpoPlQJVkaysrxt4nQ1MR+hYIBzA3t2g3
dRxHdwMU8PXHzhLyKjDH2wf/s564IyZzXi8vfNFnV0FHwa/2cAGLM5rIg9ZuqSzt
R4INGX2vttvcg7Ekb5FFDm23sUDHv3u6oQSUnikiIWkxHPwa7wyluZ90sqpN0CjV
m42CL+Yng8CBsG9DJsDucqXUCurojKEauoXHl1qRuG7LHlLDofEUd5SQGU7ewMTV
BEEU+D1vV6H7g+vEwSLiFWpRod+P6NRSfFwKxVm1OFBgTcXcr1+e+JKNWv8AsbB1
x0FOF5ISs4TM+ZQC9LFgia+QVMasIN/Nih2K3BHnFFgj2JiykkjmuiDzPityZmaW
PSsoisuYqiFeJ/Jx6RRPi1I4P7kK4TFNYTMCmRq5OudB9Zutj1I1clhELHqClDVS
ceYY6YxZIS9iK5jGTKLLqZs0hhzHF3rUigTj0leJQyubT+za388mmGpOG6O/7mCM
iOHw7Eg5yopmlT4rN8+5ZI6ST4K4hRha7bRLYvX0CogdNy6K6izal8ioSpB9df1Y
3ZDwnIdv7+48Y8R57zkSFp6KG8Kgm0AX+dL/sj9I5WSdhgYlGaH6azVYmQIoAtsA
nKWTsijTmxfqAi5lnf2NUQVyqXZNyu37PD24289x/Tj4bwKfov0c8THIXaK5cJv8
jyAnBSwfRdF4Aq4lyYz9lG5p4iBhp1eIktB030JxkuoDExE/51Ly1AromgwvS4m5
5dzrGrCQLRlF8ijWzuZHbmLGchzFjQ3Dwm6md+mu2PhDgzS6Z1UXorG+qhx4LdL8
qRoh1QGJ1MOA3a1gfhYQZpNbuUMK8gBImF9NHyStFSfYkB8m/YltZ0Z2ndF9cYXX
69DrFfVE0bmTqP3WeE8Rm2xIELSFTBKkiz5olXiOi0P/IMB7WZhTozq2KBkDPsf1
WR/p3fEq8YCwL/ccYoUY9eAE/8LIIUYv49TKiMI6glQWssLhn6GTtFjXZHoPmXON
x1mUofC+vQ8DFq0lWgaD4yF/NKO/WI0hMVoPw4DBBzStYOZww54Erl2YuRWs5YVY
WiTn1Zsq1DGRX2aTnSgWsVvyj10+HnfPkJzZz0ALVCfgbm1200wTvg/zo6qgowvP
MGl6P/fHg/gTJh+WNl3WMUkuGwkCBoMDQEQ4QqDDzWsrkunYlPNjvYw9g3R3FSzy
5OSH6yCPcx3Iqyo862tNaydHhaSznyTLF46DpqxFR0YwBm/lzk2lJKJ/vd//AxNH
fk7tnhQ+YGJ9t6EuO40GNJtmItTVnfzKWxZxZ6esYfxIY3QNL2T5jUAUWDzSrcaW
piiT3GSM3zkJU4sJAYJpisVMXhQP4rE44eVGDYfnoIf0yqHQQz8jxW5y8dBI+xzw
Oa8pftylD0llvReaDQHnZhmV9aR61VbuY+q+bFESdWq2hvw5iL5P822w/iOo7FIJ
Ngisjjy/2duEW1Hdpn2sgwKAVP02Yto9U62HOyHAx8HOnO7EHXxjBSpWLFVT1AwH
EtzRFvF6S5Fwe5+lcrP2YzLtzY3nXPJr7TghazBZKF57dKpf1ogLdrDnAUK2F8FQ
cVI7wMAPegAbfD2ODh2yRwL78t2e6aw00jEMgg2cngqR0CLDhj2HdyFjkJVV2r3D
dcjGuL4709KkuHg+yGc52ulScSbTsJ5022KEUqFbepqcQqfpI/GryhAktwf8GFvM
Cby4UB9zBAnds8flq4d4LFisXUmrByvThWmvTdYz42WKVftd3KwkLUEO6mG6fENn
kCnZYHhBfnxFmbAmER77QP5VTu+Jz6AVXiRESIjkpV6tRr+w16rhlx02OHwa8rfl
wCPzsG+RnAGwGDc8BaoiSL/yGGLWLAe8VqOMCQsih2Bx6DBUK41kL9J1GMHQqnIg
It+mvsawvqZNWI7K+oKvlGkEC9JxE5UIOMSxkcV71kyCNqOGvNaYm3CG1ORUz8eo
6cG71paIr7/fsWnqxYdQb6MPtr+BnWZttI/CToElWWW+18Wyte7vHcAUXlXA1v6p
L5EULvGoFRm6YufjLW67PnPdED4Ld/fUVCXlvSj7q9WkeyGnMwtNfnV0SjEGRIDi
icxQ4AJ9dnJybYQM3myfKpkFmKb9iBkVHXEQ68Cthg8cBdI3z7FXt5LJjv6vfNeP
qy2eH+t81j+M+w5b1GzBvCqorUNzFzI7poxvOxQm6bHUUWrbWDz5TI5ip2cuZBwm
eIUE6AS2AQ8ymI9fbnmAMEj09sgxNZvubLH+H7KKPvUc1ZY2N4JWt54ouCCfwFV0
/c1JUJAgOoaUCUadW6ipLZLWdYgwdKSLET0GKXB4/nng1jkl1d4QqMHLCSBq8IW6
NMtKHHTigMjdvM5p8JtZRv3/9o5maNeJJfXV663YOHEn4XxioPck4MyTbfMsLU5i
t7Bg4lXVsiwHsT+pj+Vtlu1wJtetMIdVT8leDIgQ22Jf6PCrMHs8465Qb2xDtuVK
5JK8Z5RYs250WH5sVqvQ1lhvwVHHR7I2UcJKPzY2YXo6ORuD6t2S5kSbgiKljh0A
3pR9xqx0H+Fd28Lyd18VqZWYaqCuz5E9LDv1AnnRd4zDmWkUnGIFdwqOPn6DCS2a
BEoceFVU6cYwAN09zRJ/drcXQlXX0JPdf6nW8VEA9I88Eiq/RspnQ/Ortoxy8QY1
HIoE5H7ZtV7X5MOpS5zVlXmjuVhH4ouZevmTSuEEtzd1HbFOTtnfbUW/cNhZN0Cz
A/Uwxx8mvjpBenOGIpMaPdO19+NN+LTRVJigSVoeP1t24abjTC2tSJA/2X9o+EH8
WvLgeuwvcSF0ATTO3tUch2Gra3ITx00B3xZEICGtVhSnwIiov3V1w5qW3sD2bCsq
bgV6FE/9Lf3u4yvyqhK+9M4E/rFNAOEcmuqzw1dx1kKgezhm3W82fb3EwUCpj4Nk
fYCAYcVXmjWuNqAu+GVS492+JQ0866jP/QXDjjgF8Mw381rg/9pCwCC/o/4DOa7Y
w4SvBOcxkckEjHWgBTV/rKYwZtz7tZEzWU63CnvE81qF3dF+l5guNVMdUeUKi2M8
fVtNcx9JtORJkXQ5Ow86vmn9yS/n44UKSY+aZSSYKj5/wlTEQ10dz4CayNpyYlOa
4qTBShSf4km4frAFrAPiZt+5LfNovoeLGga5TPoygvSvdgI/Qaswyn3nEJK//IhI
TZUHDeKiYCTH37oo7rG6yHfp3Y8zP5RnHF/jbN2lSr0jztRcTBmsF1G3cPARdQx5
b5CwuNgE8C9g+8Yx8mClPcyAsnSXI07Uk06HcAOux3co7BPgIZpzwtaEOxV3SxZd
YNp6ojCE78mREAoqN25AYnO1yWmigXe9y7acQNr+Q5EqSgK23LV9+umD4/G5Wtkl
WkBwuIZmS5OHhke2XDoObLz8b5KYrjina8/lasitSpwfY4pv07Ujcmp+cYhIVRLe
3w8J7qialSGyeBKCb4SsPCye13iiY+0s1SGXADtiLeAzaUjm8Hx1i2x4NR/FYs/9
sqNh7vGu7pZWS/ipbXmFVS6xZeiqjfk2htRpFvI1wOK4uMCgeh2G/Ssym5NJavne
wJpJYBIxxc7fU5pGfarOHnhyUszqZz5nG65xzBPH7nagX4aixbSjRuMcLuWKMArU
uWfWaPQQi9kz1hsS2udjpqU19xfk1/FzOsobbpJ6VRokpgVqqZdzjBdEOE88ms4q
DjE1EoTbjichHydo74TQg14VCM33VeyzgJiaecPDLjC74KYUzpSL1n7MFYIgCdSZ
XaBxTNm5NpYN+9W/5YliWGwXpqFrycxvmIlVmlmU4t3iPK4xAVwiQcGwz3aMIDSO
EONVAZhUCqtdpP7MOqZdJWT7pmFNZJdCG9Clu0Pmp7Uj3nFjZrrZgGvAr2QhH+NI
1qUNicCziZtF8Gbo4c2haQEijiexZvTD67+lLiYrwPtDBfNF65ltdFzKYQnS7OIU
wqSNGSiIxBvJe/pdn4x7zWR6/4db9uGqB1TNnhZyEg2SB7YMc6qezib2YIriv8ZO
SqiwBtu2ysVDMI3QymYEAL7dncNVsTJwCSx+QdFIKINDsnnS4+Ted2tV1eczyCQA
rQrk3MX14ajQkxWLxKeIo7v/PNx7tDMZhVzKuKDRCIKqEdr9Jynh3cbS3kwpe+kr
u2XHCQgiiSTqIQztlEUXvexX79ug8W/nqbozCLE9Wtr29rqPUD/UjE2hIXbTR+ie
c5tgLCtDQdscp0C9nnsctJSWeD+PCd/oh0pQfD1aW3g1jaNH8OINNdW4G4kIh+AC
JcD4E8aoPzT3dt/jPx1wYdjuTpkF6qVhzqguKKMlK39vlDgCKfSHXVgFfqCaX1iV
T2bnEkUptle9sm4EKrB1FWedxJmE38QnUzo8iXbLFhFwfVenDM4O/Y0e6j851KsK
kNtprpIDSTKT+s9TOiNDxhelvn4URs3MiFZBOVYn/wYoVIkW8oqqPWXYpn+MvfiI
7XQmbR2PzA3/lfZebjGqIzdp+/jXofCvzNP8setPj1aKrXGFrNyKGQ6B5jLQn/2+
d0fnfnL+Dwk2pJ64/+xEexnYAHO3P2X/Uirp7HGb2nxSICycgOkq1yrbvFzgCZ2M
00/0pjF6N8QzfcEM2R0XniV8o0iIdOjayZiU/GeFlGrGOa310JOsBCDOfavEK0BB
wn4ICdh2XMYd9Esokr7+l7IXLhzPkXVy4Im049WBaq7oaUzOyQ/FRDz8+V+yYMMK
EXEu0bEMNZgxcRi3OCe5ui6gOpahsv9cMRg4HYizqIgxryiYktinnhYhLcEzU9tJ
ZPT9iRdrpE2Q12gUwYSBgUc8EJBbyImyLf1qu4VKMiNt4rFWKPfaUJ97JQJh20oS
qVkNrdqE9rjYCQLoDnQXLwnXHNsziOJ75e3gCwKfFxpOjF72qzfRHmZrNmwNBscE
9f44v0AEen0zuW1Dikh0STLdJ65r/szFzS5RlghP2GkmZvYfwz+QO7RNmcEuM2Gf
q2PD7uIp/Yy2MaL9FjdKHknFVooWPfcb1yLBEpexy2elHIwLELPWNN0jK7bd6NPT
syeewAute0bz9mUVmOlRIkx/yHlURCw8E8kA1+jnGeTiOA0XtGjtxk0wYXxBZAEU
R8iwDARTH17n8GiuX7WWVFz6TYSaYxgomqnm8RKP+zItlUMoHCADO1EOVl/pRhWe
Fhd/e9yzvcuqs2syiYo0GG6iutaKHjTMSjSi/6ZZniprsZPd2UQH2/+CQzyTlVWz
GCEii1zRdH+zm7iA3NUU+k16Q3/jllG7d1Btb8tz1BdTSfYKqZ3FmVI35oJ2e0bq
NQZ68F7GaHBJ/d4UkT/YNzwo7gKLfvhFxA+tWzJzp4yw/xzZ2Gg8xUq4UlBktCO3
1BShiWZat0CRKSbUjpRuPwCunbEggYKXbHBjxGh7QMz0aWIZpjKTaxl/gXcMzqMk
WFqmw9ZEA26edJ9aohShKRPDkqW6SojkpwHaIGP4v+4SgxWLlVYikLrFbE9d1GMU
tIc6GA061uff9p5c/Oblgw48ZhAO5O9vw7RtIx3jgoshRXjkLsS1YuFlfN8bOdDL
CoxZozR/JUDLNB3/sojFCJRqDKJ5S1luszx00SYPxr1Anwwv1X5VcI6pnlHHK3BU
PNszcN8a2pTF9BUxGPb/4nFN56NijPLG2dEAUIjThWLC2F6FCnGuDNi4qpAvbrIM
lKw6HkH2fXil+hEyHNgexwBnBFgxaSKFSBVjR6CXHRP6vtxByvxsSBPSfPV8C0h3
SiHMLFSrgdC903Q2QhcP0oX8XsyLMx3vl8zwXbP08wBAD8JC9OwB/OGrg/aPseny
wfi+TCu7eirapTgI7AqOVspTFGRhGYtGLLtrSslAaQRbK143aBCyAciHM5gPzGbW
kIf+04YrKZJN6U86iBFn4QJnwAHDDxrfo6uNwUxbdR3WZ8ZzDqdPys4GDOZx9HvJ
RQwP4nMS1aQcUC6MXsYA/V+MSfCCC+g4uvZOCuEfCLnBTL8z+42W0ybcQbt6pL8u
8amfTPGJLVYZJMu9Y3l/a22OH9lom4oN5TeRnma37Oe5tQpdNSshBMnZSR0gezEC
STv58oLldPMdgO9oYzoQv5me7S8kXzWNAWK8M31SAkgBD0bNBGAj1dMsAnXIBB6u
vBWiWQaHg99mpP1yFDlb7QB3FUz+SHRfnKZkf4K7/qfgPW8NQO97RmsRT5gWnB3k
J5RwfnmDP08+5iqLahkgHqNWwN6g1jSPqT+BOH8lZg6LwuyGqz65uye+zg9SbYur
uHAAuHsU7nOsgnlzmFQBUo6oOqHPn3bgBet1tb7yCbWY+5KKs5I4QEfRxpYTQE8i
eaxZeBA8+F5Gc+nziIU8y/5zow2A4ZgTarkLnHDsdJbWb1pLDnc4+n2wf2QkSujL
E9PnzDFBrKzTEZGr+68lWQwTOVbeAn36YTrTpT/KnKaPPFeOuCGe6x44PapCnyvu
H/FTntYsQpuiwj6B5O+FvsDlJbGl4GsEQdIRQJra/6Ja9cTQx4di2gS/3S4fcgzw
boZ1NcWxbj5XCDezLNScS8QQeHzqEhRYXlrnmgkW/zPaUpXJMNEJZhy/IYWsAE9O
zn/Cqs405iiP15Z7FZ3Yq6jVRKg+xc/pshfH7U3gA3aEMuwk7TSaytyxBa3Bkg/1
0KwBRe1n49a3znhGHqWj98Qk5d1IY2Y6Zynlh2X4Lyv16QypLuIXPaRLPOTQ9V8y
4BEggzK5hBWakgl46O7KWEA4tz+AhacThyIvtb+RBKAZ6j4NeqzZN3OYwszeBz4P
KZ7IkpRxMFhxCBIHLVTmJObJrSOxkue+WlOD1YP2XmanCo8owJtiXoNmnDIy/F7K
gyN31ULBMpycRyprphGs06tQbGOx3qfsC2Tbhb/lK9p3vFhcJZ+D5dElLC4f3qaQ
FstrU5pB7FCptcw7lPMBS8EkOKnyy2yqUWjrB15ICIQyK1dp31qofJYKM8VsvOJv
IrdOTvk9hG6ZCi8ho3uH8mRnqfBkjoV3A6tlkDSbejAkRWB9P9yS9cTGm7uk81xw
PuhQlaPJ4497zkKiuiH2YwT5J7ZcuJkKmO3AEbJavhBjJXE++qi/7j4Aa0IM/rMQ
uvRj1Ti7P4TX3nP3b/ttbR6x96xPygGHNWwkS1Yw93AiF+er+fvIozkk30r7wdM+
0tsHYXpLGgTW8GpTR0my8SV471i1DyCojb+++eXnBKwB5/CbJBeCCuAJ7/D7lYO3
aVKCCACzjIo6MVGVvSL+XyY3jIdV9I/aCqIh+EWVRh8ydn3qaDonHL0qoll+0lzn
J9QoQ/9wcGTLDI+IGEFeI7FdNsvPLDZYnouok/nUEeGXx1TQx927rAbZynPMdHBU
bGJEmgN94JxKchs0Yp58911GExgpi824r/YP4TcbY2Q9e4kqNaClmJr5A6NhfJtU
nMZ3u0DHePHV/8gAagzPTCl+zR5p8XZ0GDd83YBkORMWSHbhhNldyxQgygyaOWty
0k4IoCrgyZ/GaB3X2XuEFJB5TjXf3uWNSULWVIJwft/wLB38RuzoA0imDa6yGu3h
92npwNTpsjfSQw3frS7jMfCz1ewTnSvP+KK+GPn2Sj74avDMhlWkiq0PIkudvBeP
hTg+iBZMoE1Q/WRRBDqyyioiUi9/KOZnzuQOoHBjzimVrXwfBg4YPAtcLmN3UQ4r
WjtRtkd2tEXFV8rjegHwDiWIJI7p2DJ5L4ijbJO4LpqBb3j4LvOEQqGTx/xArx4q
1DgQzjkxy1+zkWxGNfVCW8T+eOavnH5hEFHruiC6EwbSt2jmlKWkxB2JdKFSNJur
x5OOB0dtBxaJaCmNA/wfSED3Y14jFWhPfK43pPttwux7V3HAtJxcMu7QMTRfDMZn
ctJmidkE+PUarFTNCPfyenxQoOdnIXzaXaddopqoDYHscr3tUB/KpSx1xDHXQyr4
blRX+67ttMB5+LkDdIWtxU00k3RcLlfa0i0OzzlPRyfS5UxU4R7os7/m+TxjjM0O
ic0evyim0Da/HoQp/vvf4UZA3urtqUMIv4vE/yISh0R1y0OsSSSAQ8FLuO2mJSFU
uzdFgqTugBj6ixBMzeBFko0HISIgsOnQ2sVBqAT6FswPyDmYv5hr5h0mvCNwu0zt
+V1PVjtK4lxtMLC4HBLA0tZOMvEE8U8KpvlkkNZHRqkl8+A1uUS9WuryI2748hQv
y4Csh3v5IM3CB2ByzJ283APdhC7ONNaqJGn4l1H13xxjZ/qPPTn1QeCUQkXfUZRf
H5gb2w7LFshqiKZK/Zqg7MqhfZUmfQpKUlbFZn2Bn6CHTAwFZPQ4BulXxAhhHbLw
Fo80AxFqFm+euO/j3nUifNubQCgxrC+uu6PRVCKPvicXkd0Ln5cQ93R8PPCJ5CJs
T7Np4uZt80qWJZpYtlJj3CdgthFiKPmuXt1NSaZy1wCqb1POn5tylugi6u5WAmX4
PO68bVr7aFBCRCqJczFfcCyztP+6oEZZACsjxvChzebNRuMzfd1DW7SY/K2pLhUv
FkDMts7in3NF3u7wXWDkp16l9x7VAAtzQCOmiU20bwxoymgzbQ/aAdeBgNNUm4lg
gR7EzeGkwjHC3EbKQFK9wo6cVgoZTyWkYzkMNA7q5wF157V3NrTmwBIBXsyAIAPp
1qVZb0DP4xmwOhlcmIeMWFW+hMmxd4M+cu/wEYFYCREQXMgKwxRJWnUOdA2X0Y6o
Gyx9pfUnAUvraaM6crRqPnLfLtYYjJ13vi+8jjrN6B82oxyZTRpFJAevkD3h7pL/
s/zyvTbVx93b4bo5I/O5DdtFp2EM3TZlhenyvavTxmBn4mQNUzOWHjFzN2H/FBhX
whSsDe6QH7JrStpP4oMXety9nbqFFnasZv0oo9BgQxyW/CbN99Kh56WVeprmwbGu
MaUyU/vOjAZ2UGk0Yrbdgv2tY3tTWp8/KnZ65c9RJrVUlJaue/JqcI/ahKoTNCpL
zXfTChJFeblNYYTbdXDplSwAvSFUFGG51PxV38WSY29T38i0JPgHbHa6JyjTw34m
EpS3Zk9m60r5pRfui9F+iq3K6Rs1Byj/+Iecgl2XfDrxSiA0Tfc3ElsX+rTDq/ER
meXobeJCGHhIrij0y5OaRhk4HMBZ62IYRLMIMvOZ0nu+khx8wty1GrWAlCdJwfqf
OLrrfF10AMhZszULwNVrtmUhuC/M0IJ0weLC+VdTbl6jrgT6XiAkgHiDKnFCSUzO
Yw8Slm8yQ3ffaZmzZN2diP9xSx76gQ2kSF6Pm1OCD2msO2CMh0KYfj1i6ym+P7Rq
HaDsPnlZIxPl1L2xHF7nLdFOWJTMYeBpvWps53qgfd4bPj12iNm07HKbDbIcS0FI
ahTfFRp0JL0jL7WsUyb2H8LP6JbsnSlsLMnTgq7EFMFHyLmhtt988o5iqvDkNJ7i
97iO1C4gftSyHm+LqizrNs7OgE7f9f6XRcneoEPdAOb9iwaxGyveIBlAVcLF2L85
d5gEc86euTClSIDVVW0S/ao/KNQB8xm7sVOCi/Sas/jLkSv0t7cD63LegyLY1fdM
0V+uolQ7I39CEcv718PwqwPyc6jCr2IniDIuUni+sko9Nue4eLJBBRd1KFny+c+Y
kbWDFw1SpHIuyKFjhLs1e1gv8zpFvjAyZRph6PoUo0zJJb2DOzHlqG8RPlSGjKOo
tCAXBFtOyENC2B61dTsrvZwXPGQQwf5Zv9Cwszv8e0NscXpFBFMJClwqFs6r2NI0
GCFEinXStrlREGt34iXz9tpbdlo6wliW76SWLEaSpOi+2n3pEAuZNv838aMGsXfX
X/NJJDky8OvCfFPPyv0LzZQqKCXv6e22sZh/mEmG5RvgHs/joHSDxShhiNP3R3XV
NZ331Yl8+kVv6iH/qfp7kxmxecOFcw2YJiAy04Olr6XVaHmgwf9JIecWkBjajFzj
4tFfCU1A0bCUhzBh8dgkQ06SctMm5ZqNTDfC/DMlVyYaBY7iTJLfF1p1B8wJ/CX5
QnQtVv2tEZuxYZm/sBCtuT51TPaKHiD7MEbuExcYTBQjsLNG4ixXuoIeMopWZnd2
dFd2VuTaAz+hkFcuxYYzboLcxq2+8YiirE1REC81duJbcbzMBwYMFGF2iMAfvZ5M
PPq+HTJKeqcAGAIHRJuXT6SDdWBauPk3wZITaNwf+uBnSwhhrnBIQwI2nkSClh3J
nIGUSElHF7L3NySfhD/xvgdQ148xJBrzvLUV2jSZtN7TxVSPnfJ/UnczxC6otcq9
Wt5MEkQl8Mn/2b9GCPwb0+snRTxcgHmnHpUQj5sg+ErtrMrX4gEmCd5Ob5UL6jml
kpshcTS0p24tPh5xX2083KtraZi5EvPJd8gllRuFDOqZQ+hc910HnBJJ/SCdD9hX
KvTlXljV8lDzXbQCtl7WfZXJUgZeP2J+N5wBzMcVJfTbsgnnEU/vLthIb8UhoR1/
nwQOBgc0THNje0puXzzZksGvVlZF9d8rr9pGKRRJvpaYHF8RXSLTOcyefndCPfYa
vBvcWuMhD5Ttj7w55gp0L3bsxyUJ3IbkTsRZXfBioL/KHfOC2zUhEHdr55lhffn6
97hBEVeyuG0ogR9sV0LV2qUsSKfYB9D+bD9K/fQmA/KDESt8z598R9EGvX4I3sQ6
xwAsoBESk1emLPptN83TOwi3e9+uNiS8ztTtt1ej9075wyj+h0sFw1Bo8HCBAiGk
NlbzUxSRiIMnsyBoFbPQ24q3+u3/S+68RFtoCjuD350cSHS5AIiz/7y74Q1ZlfTK
nCzGwpJKHRG11kXb0LQ6ILfkAi0GczG2PMy/VBRGGPPGa0MTU0UB2fW9Ct+SUAYA
N+7LKtMkJYjSS14fmtoKissUsqBmhSyyq18u05rnvNkUi13zd7fvdXn96gAJiCU6
u9ks1PrbAelxlTTjRkqCqjTDcILxzijl9rUdt+YWqYbniF+Pz9gzpmX3qlxrUOvB
ywNdOTE0ONKzJBAz4g0wwDnvxkX9RHuT0638TmyI3dQIqUG2kiHCSt/HKseS4+f3
1YmN2z3nTaT5SJxMMkGWkNMwAS0ddds+9unYTgQFqW0FjF/W13tLU8folpb2JUKJ
rMGuMwNK0Kp/q2gzTY1hmvPV+LrLyGXqKlS3H0l7sZToDuqOAJTBYa29twecO/bO
T8+itBRRHCKjmyKJR2T7MD3Hittav2QX1x9ByvCLOwdo0kf6irW/bwKMXZ85iKav
CDEnc4nueDLUBHqhuEfZLlXTscu6KvPTqrRCj2tOAeo2Vb6xsZ7vqsNO+JjtyFrW
0vZuHJMuprzN8RKPTVvnC1irSUBQsd4wgvctno0gAXocYsj7OGDyVz6QuYK6IWrT
UIicUcH0lF+M5SutlXBQQQgIrNDB0eZeIyYWm1A7+hTxdfrn13Z9QWT9R28Wdti4
9mgbDhSgcMDYE39ejNiQn1nsNMYEbAAmMQ4WWfQBv6ZlokVKHoyNQq4DNkzQT1YZ
/xRabkINb3lh+JZYwpAdeyWZyDEpG/fj/b8D+hcJtlHcKGxRnSrjJwOFWcL0NeZq
t8mALujv9bEjE/49ihK9p6F5EDpZp6+BDA/2L7FpHIM/HotdctwBs/3hLV5i9Mn7
fRUzNapmE6UebWQV74XDQznSnDV04lj+Z+to9DwHZyAsJnOumoSOpbabp42PAFtc
ue4r1X4HupzSc7ArgpsCNJ+vC+Lf/ry2Bi4BLVDOW8OZLGEJJg3cBB12F1LlwCv/
7T4QNIr6k6wLmNkbGt8s4knjNlmM8SaHlAOXdYAirjql53gwe0zCERqtZOyNZu+S
0FpAsNcupA8+huq0iHJXLsbVhC/eQjo/1VCHdK7c3up+SmrtqQ0SAfdKr4ZugqEV
l0P1JNHcqi8+jxg3RlvLW1K3pyJdrFo0IvdtaGYqNL4s0GmKirZh29K95B5xIKn0
Hxx4Em/LVNothgQ/mV8lEC46gxAq0fV3P0Vjg7xOx9mLSFx+YrTJE7kNngRS97iS
nhAOiiN3gPQR1KHeFRESPksaIAWiPBara7CNI6OYrY69D6n+d6vrzfORyzRymxNh
8I76mFFqEvaq+dIebWdrMWtzZodMxwh364pUlrd8wwL5ZAJeMm5T1g4m4MXlNvdd
3MiC72VvTPH593G5DpZKzPsJ2QpMxajr1ORNZ5OxSFbSs6uFYlHRXGl97VJSEQ0v
6kTd594QyPqMgTltBxESjTzMtx6qHiMv9M7VQlYPaGFnVwNjsR/B2XMfaj6gYel8
bG7LMhwOsEI+TJNtlVKiHJBiicn+OScrt0QA4fI5K462dvRULPUzon3GQXyJnoLV
oqdGSUhGGRZH8KhXqhzG7SiH8qOd5SIoscciAA0/1KguG/+7oyF9e33EvtSx+ReP
D40Kze023eCOkg7qe07JJbX16l2m2frsMyoycuUiM4wQDexjLUlOw3SrOD3CNqSP
XNT5u5gRTE6kEgs2g04oJFCpPloD+yUpGoU5ymf/hrN/Q2FDluUIMWIPHgXeSlw2
bOifVxcDeL0Aut3Spwk4iIQEnc/Fu4aUZEGnswioL4lcbGM/LvAt/qRVWIYNQTy2
Twz+Dikqm6sA4RBRsp4jAtgmGYibLE/5piS8wEMUxvtk1oC4wcMFhAxlX0WDjU39
k2bWor8atUpXYa7TolO2D3AJjb5nQmaJMFfglJu8Za1Sz8PgPZUUl7y/HBrEINOj
ha026+kLDXJYDo8K0hTsgKpfbO88ujCPKJ9tdp2YAddF9DBowI44NdNeF0PXrRQ8
OKtE/00LV1r1i1G+jzfSbYUNcTxYG9PUhexd5YEsr9kwyjGxDKvtnA8gubHz+SZB
2HAoA68jiiYyQRWbWA41by9fJUB8CIW73c9aKk6vslICUVkVcNTMYB430imbBAT7
zW2A0FagbPQ+Zr9x9WRdGVtdZpBRZPaFGVtxqFCysihKP8mByFlzvCy8jxLAvOoi
jDNBM+COGGw85F253E5xy3C58dCUq2XuJqihXig2+Dp3v3+xZvx+ENcMcvppLrLW
6lEnz/61JLOLwgkwWg36uOqucULuYYKZCwu7unF7DwTlVDZr5q6PjOIoiFIBueQ3
WVCSiT/n68LsgcwsTX16NOBgkWIr1YiX5/dd7SAAThgd0ja2lKWe11dUNq3QIRCp
leCw5rzDWYX0eF2BTDiLjFnMeVtBxo2LYdCkPZzelAhIYkDA+o1Dppon+6yf8eSv
+6dls62hjqp0hvVhwdzQP1mDIG2s6hwAz7gDY8o6mNM8ZEWBuSOJ6NjaB+ZaXXOR
RP2acnRZWNIeRkuZbHLuIFCjNvooGlkys5dFuPKKoYd56ZkFHnu0QMVBMzX7H8Hh
FXfGOofvv8kBKK8ybCs/49Cgxq1wRUPxowlLfB52DkA1He+ZR/WDOt4h/ZJ1f2sq
UQTUyLcoeeXAO8DqcygDOjTNzJZBeuuoWDJMw8qD+RJ0UnuH93d6Yq0StvKqusfM
+3GKhAgrrqfIb1j3ipcyvRWG8R0AQ068R1Fx+ycx4UZsF/s8rleB9/zJJaH//LHv
r3/gfr0Mzyoa3DavABxD4l1rXt9JGyJ95cDOLmJs6O958emFXKC1RG2o89Wp9OQy
/1UaM0L5EAQVGRXZwBWfN7hoEC7COHyJN/lEKG31VcX3Jlw2nXW0BgPPquBDDKG0
SHStYVb1nH5p4KZf1GDuMsFBcsz+l4WOYp9US878KZfhNMqwyEGnlcl8L/qyCR1v
LOiPSdvSywwCqd333nzw0xqUU3v8Fr3qh/K/1aVPGaYoP6WNQwU8NHJko25HnTqz
wbFWjC6UhMg2JomAaQTo6oO3vSaV+iny2lEheJNmMpGV3SVRZwFGg1zC2l1Mbvua
0C9k0cY6dm+DuZ5yCVnq2PhPemusIcBkpzM5FuP6f8if8BAHHW2ZbDsguoRX/xHf
WzJul8RRP3ur9zmeu3wyElQTyha0QwpV336HZaed7GCeS2CU8ECxNjAsPWDFXaMh
Xj7rN9aEzjrlFVPMvVMnNNSqaIZ8gkYgJqQzcvmxi2tMVoq7YvseJ/wEUeHFq1KY
A/ftjP4Avb4LKMou8xE8wN3vpH8Qeelswkb3D58KenqAgavX6/+ADEQkapb4zQpc
YDtQqDHnFZx8iMh/kJxMryFnkQRtf+c9b2bmbz34z96ZUbCPaiv9EzMA0x8vCsmc
ET3HdblZBpZizTuXChNmUuvMhRAUYlku7rz8Bf2rmR6vg5VwhHQpkzU/95eFQaEo
xR2BGSXDIoSZyVmpr/bsKRh3VRTBKRPe68Qzy+aoRBR3xtyDH8i6jK+sJvss/5DE
zLRWZja59Bx03iJsfbxy8lCUiunG8/WfzzzUSVwqXyVcmiqTv9/w7gMmQUGpx7h7
J4INTt2YH8AjRtwDw13giNqMPSfLY0vTOhYS1cL4Vr9IUTWAeZkoYJwvYtr9d41R
6UCqjSUYNp8xJkdIe+twFZFoAP5GeooRghh7kfD17ZwUPVAF3wwqGLHns1fP66kE
s1obqXV833dPeeFLiB5NGdT7KVdfG6t8qhrqkCJ3WTqYGFVROoMru8iKdvQwsRvO
k8wDjfJgMnHKsXI0gI2+auDPR7WG+H6hZEh49yD908C0ZyT/oAAY7rtWjyYNOHLd
DrFjlscMyr8YmaA7ODZgi5OXBk6Cya8wQ7y6JX0sbuxofhjFwMiWiOt188HFoyKQ
XCqP9w3p1qLMieHiFuflTwZmzOdSKPOE6PNTbrKUlvSR4n+oGoOeY/xsIYHfAsuG
xpGC1Z0IA+Z8sGj0RCdgbJQgGDJD7JQSEpekI3h4zcHULQ/CPGODi9/NSlfV5taA
NL8NkjchPCcsGzyJluG1r7LEW/0f9aqJBxkwesNQtxZKgtGzyq4RD4ccJNXVhiNB
7+2i8ZpGm2L60ndxGRsx0BBjWRDrLZDxTbSXOFIYoQDtPZ/1N2Ktial/P8Z88G/D
61Flsk7qGZ64kiXymqaRY9LGu1pUAdgIJMDqRQ2iVTkuQpI+GXDF67Mk3SdgE9Yf
IL6RD1iQVoBEEpF7rfc2EWeQMjlkYoeCsJLJWTDxJ9l9iRT5LIl+OL9S3vZrowGV
MWwyhjkJO0ZwFvQdyd0p55QjejlpxsYKk+R7YwoI3w7F3ewo1b6BRfZWGWwE5q0y
vkE7RNQD6JFX6rte+1oWcIJVVrcqAqXWuab3bPqsauKireDkRZxlZQrQxGuysTvd
RLTc0SbDrerSevogU0F/gW1wKBDIFft0MbMLI1Z+VFWtJC5TxkOB/gQnSFh1XGcX
0wos9EJPrVryrxf9oeRvM2F2eNabcJFuRJVJjCOMvGWJpBTRcXaWFNCVjofLfkEE
tqUAL8K3wDRsPbc1MZQYx6cSDtRncW94OJY+OjxIFZAF7SinUFthap8HuG4cQjmC
q9HSdJhdxZGiu9oIZZcq2RmdzjTm2JkO61owq0KEGYRDlxzdA1k64NFMLlc83z7W
9Ihwmg7PzlggLYRDmeklWsrj4b7V9LTjVGg4yGLzlkcOdO87RFVcr1LsWEEL40fG
tw80yYLGSvdxE1iqwxn+xbBN4HyE1//at8oscggnW+KojXdQZJyrLZRQs5XRdyG4
gD/6kJb2t/mH4r4rXJFdW/wwRRhnXgiVwRw0+ayBs5P+Ni7UaIzmllyrKDkWuAVE
1enpQdEHKnw/QXbMyg2gmsnI97gJSO2aEQcXypPV/26aKZO0cx6HaGJZAr1jh5XE
EQNtbq4ESA4mJhThwHmneMvkqmQNodVQrD4nIuwZcFXxIXW4zQtxFHw58hv+f6Q3
CjwD0aR/7N+g+a0RF4Jhm1PPc5U6Xt42eg09X6zztdTPFD88j1MkyjNd+HnPNHmW
EEgu46/XI4g28ArNiihvwOj2phUT8Jso2rKKt40fxV9YT0gpJsifons71yG/Dgxb
2NpVLKxWM/ogrGoU8DjF1Yy1yDbBiB6T5AeZPnwtTA4PocEtybxUZnAUO9AJYdnK
SBXB/fy5jakCZGxqfWdyr6dizapX61G2qktc8LSxbF06+gVKCFHtOK7Szs2UqRKP
xvV4eD0tF5nd+ArXsdUrzds1zPToDm8gWak2EL6nLTSG7Kvsbp0ysrtpYo8G5dnj
Q4GFvWO3b2FNnY/vWWm21b0FU1sPdpN6BTePgezV4hP9SAIGqGRKT42Pk0lpw9fD
Awfpt6TqLiY93+sok+ze6LDaQrdkGxMLljIA13aN9q8M7wfBrbvYUoPcyS+A5sgj
gk9tXvpaskEO+oS770BMBwidTc757+Esj1mN301MpMQo4wOShP+By9wXi0aVBbZN
U/Vsj42OFsnO820s0KSWnagg7jPxt/jGo4oh298RXs4aKoVFNRikU/+FNFBgqFFZ
t/4ygHXtmDMy8+VnHZAQQjnOFnR26s7vaNs6cb858fxkJ+9y8C2MG/K+4V+PXCob
wSiUsgVM/LaGgUXQk4k4PAZ9U/IhV2hswtEIdUHuhtEpjLbLZgFu/pFew6Jtyvma
AZkoHsPHomj9YC17ObPDXutZ74cgrBHEihjcb64KiUAL/6p7bEfyNhR7SR+uX7bA
m8eV0gF+JMjh1WWm/Vfcad3Et4/s2+Kl6KSXtKSOp8DJm4LONU9lg1Oa1/JLIRIh
KthnFTh1tIsHt1K0GFjC/H8+T/Wc8ft/WVTnwLfbPhvE4PE6xikCDSB2f6P13ZeB
y+M7Fu5x8TOvAEJvXycsJ3iFU+4idQ3VbPtaj6A/2bYG7GYemeGwJB/5NuZJWa/y
eLl1cgwQGyO4DcqTTPE1CtzOKtjWN7MgSvhR6ex4GxdvDlyKcMakUANaRso+qqY9
1rkAbHC52s7Zz1ThZW6jb34sEfhlu99YjUhf7Wvc3HCsBs3dnP3MJdzwPRg2/7g7
nfWv5g8nmtGJu4v7uJRSZOjuZ8laPNfNpv6eaXcc++eZ9rqt8QbjQuJDhYPg2bV4
BHteBiM7ZsRwLDItXhtExv7+jdD9CFtQymLP8k+PqXLG3iPtrvkfU2oKqhrG+dH8
0QeqqqoOLv64K8CvwdXQGcFY27mjsn4BBHTP9/kgJN3IZWVHQVpiee08BKZa2ipH
rE9qdTrBlzSxJ1lXLqm7PkBBpmoCHyi7Wvcm9lh/N9q/atdLyPVu+J5t5TZEyGyB
+eUrdQuBhlJjjiMjYS9fEJzovtruXA7evMKOZnKUvWhWkFepgjonzp+5/Fxn9IMz
O5SMkvYq4iVxI+X+CCBxCQfplCxPuPfH1uim25XoRaoVyKp/r+cpkcHEu8ZT+Xb0
TplPSyUcHJ/FGPmNXeqZIpBldqy1tzFNcJICbuzzR+E=
`pragma protect end_protected
