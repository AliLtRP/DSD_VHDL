// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AbCyCk4KsNZWhzNORmQ+zTShUp+QgbT88RskfIR6+L2uGriIK569I6ioXNoska4J
6S3l0vODnafKME3MKX5b7F5Oph2C5gJFQdGGlzTcDWRLU12BbgGASuimBzKUypKL
ap5piFRKMwwTyjGHBlAsqG1LrZnj3f6z7ZmTwmhbwDY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62144)
ndM85/O9KY7yrfSh1On51NfKyx/AFzZjIxZlyh3Ywj38PrrBy8PU0khp1OQfrIIs
cVWl7CMBJO+cN4OsJENd45UmbXup7JbGfoRkvupdVrBEbNPR4sQAP8ozUyKsmUMp
vIt8y7IChtySdlTObykDwxEElwmx0Ix7kmf/th/OrFXcG3ct0fiGu5rjkpuN9GkU
KhXuAbYi8KZItJZn43TSgoIcXIEbsUErCz0RoCCdOoN+RcyKvysaMjFStzQZRmd3
JpCuxWy+1cbu9tfk5m8bCbZkzJNIeODNgCBWghqIUlpFmPugDDqcwqU8OXa5s3iU
nr/gfapZhihydM1zXxXM1UScLxvcgGE2kdXqJofM86BFtHacR8JHqQ6MGEkKksJ9
SAxmEwtoWXC1/u+boMTq1LnpklYMMroQtPbNogsbk4nsWmwrXPCkZopGFZdjkiOS
arYl/gzKwwZQe0IODVvolAUmmi3SBCWti5mtTM3/E/nzhh7f/1/lwF69v4TYkFmb
3GfXEFLRciqNHzj+cXuat5yc4UUZoEPTO/8de6+MAq322aYk3Vwu5X0ZwmjVdlCr
/Za3n0N2GWMFtVOno2jTx3YvT+xx1t4Ssaz3ueiMz1T66AsuPkayXzNXw98MKrw3
UAn9xjRfOe3QwJHlYbRE/VJczqQRSC63y1ebtbAcwQKGkzP8tt9etJpiqpXyTBKT
fQqwmbbDEUACKX+USLP19pDCDUL6pKzY6n1mYTd7ClFgZj+6Ij1O54aD9x/wgYHC
cNSPyrO4FKV8rlwQIlXs2aJWB6TYLjCs3TMviflb4SR0K7rLAwE2zOHsKzxQhcQI
TGc0j4H9gPLBNPwpiXnso1ChkJMeJd5T7ho1jC/B73LkZH4zP/ss4NZlGm0CokJ2
DXXKpOXbRQmVlloAF+vVtwAJpyJzYs7JLr32H+VXg5h1QZ9Lhjs4Mngi6RmPeXyY
Pk035XTaWTkXL24vKLqHq2QQetBAAl7KpOqGN7B5sr6r/hKx09XviBC7KeBOgV0x
KBGZe+G/UUcFY5d3RefoFmG9ErkMn3MVigz+A8WwLdlKqOix3gbDDKO8NIgK31Wb
ZpVEWa2TOlL3R9mvdScVG64RfwBdhhCki7G4BJ7qCImxl47ba5bq3emom125Gd1i
i3wpPyciqBVnfWh8j8BXIjcR43PeYmaNGb5IVuZQ38VoxW3G3E7IkG9hFGzp8On0
7+p5yX2QBTMLvpDfj4UrMSSlwbW82GM7rPGYTDlp9sVQlfZbDXl6vEdD6BfmZf/e
+JX+zSAc+MlJ3T0Ssb776JOaBXoNfaDNtMpghVvzD/ojqbnnmJK6BXWAKheYoZH/
efXnhf3RkHesYvi4Yog3KzlPiP1HfAlIeC1MnOPvqKnJKI/7TG/Vwaq9W7Huraxr
7/0elfITEFWu0uSU8ey4c4wkRg+1zcJ/AdOufebXB7JCtpbnkJYYWQqBMuHX4Agy
O1dzbRtfzNAN6ty/dQfYCcPu4K2EC5m3QSnHAiIf54qrnMuI/qEYYw1fnR+8aWNW
LSyubtaIYoiDgeXW4WJA3kmVm1zcoGFWwiJmPk6SIwIf4N46fKH5BUPLbK0Y+mcE
zrDIhGjLluppTWJgtvHmadrvoQTUGmbVkrcyVezJLvtLhQo45g0p4UQpMlwEg4Zf
dG2irEdpNvxIEb2E9/ZP3AmrlbgW43bJxLp9wq39Fj0M6Sb/JHHV/K7Anisk8Pke
A6V6QFXwOhQj/4pUULfJeJxec+ZH3fjOzv2YuFaiOmGuuywibqWSGCKEqacaOoAp
QBq1gI/wnZuJketsiitDaf/03kgUntcg1NFjIfzlq0iJnJB2s9xuKXQ+joPjXbU/
oBl+V8oF4DqoRMCFYMa52rtZLbw8xb+rMI4QKglKD36S/3w/P4oS/AgdFBgrV4l6
0chrHqJS9OUruZ1Kjvfy2d1XChCy+2yGdkuJhX4nXHL5ND31WmcEMVZ2enOB3q5c
wKi3ry8sO4cZZJWZZnQWbzR6sjpQ4RxAiWBKQqlWxBR8E7WQ6Hx/YPx7A5oUwLYr
t6ortzvBKZjgk+mWUnvulQeMZhy5+KdwLKZT4ex7SZUVe3jDzZaQJILC7szjl2B3
J+dV/6jLSVSKfpPvGe2y4c2N+UVC2pw4PQJNMTHxJ0YGoUx9LP0kYHDIgbwL+HOr
gCmYRuw+AphF+4042b85G1PgtOqjTJ2rU1IIA1fCaoJmcFK0M0smuNlLkiw3eLh0
nfmXJbnIcqDeFOGC6Fst5Lblk1Ic+W9JgKIhcVB12NTwInttaw4x7oTuVrVNvvkz
Podv4+T85ePIrZOQSW9ILQXUA6aheC+1xKTI1FUgesctwuL+nZVEnrBjveQeJJeo
7EUF+VtOqt9eu1qljDSeSZaQUjZIvrdKg4ZjuBie9chKXfj6arcuTKJU7CUIoxqL
SVHfyVaEfbxsN24aQt9JR7DN6HxHIOFIDo8JFmQdeeWTapJuwIAZ+lHcobGGW91l
w+jIWHHj8fQFg+dvvNvtNGp+HlH17fMDjECaWtU12uKaxIZrxuAnroJYiKnuyrH5
JPwHoEM/bqb8urVkhmdv/FmXNgOaalQjEZzAhtrzhcgY8yoKILRrgCLHJlgaVDEv
WRHCNUEXIyp+/+Ws+9owFFTg20Oof/R1TTuXnku/YtJddAOVQ+rxd7NyhOlbQcb0
VTwYlCtCQMQWPf/rkL8cMz1pq1MI15zhoxPmTu4S7Dt5c4Vi6pA1yCimZfjjm6uw
lFM+iO129L2kWt9XH8wq2nZdqsxPWS7jX+5ARsKllR54Y+5JuLHTi5rPlJdEBJBP
1aWkdEZRMGPFtR5MCo8smowwH2TZ8hl95fYhYUinkXioTu2F+ojrVlFtsWgeG17d
TeZlW53/GO+UfBUbfKQ5Dm0uYkp6pgzKZtvYpVOj7hJ9pgKPQEFcKcHS5idDU31t
11OqpjaWDbu35KyHEoYq/fdRU4B+grVx61uxRpPpQ1VMEjLiaf3/ijXN1azs1KFW
aRpe027z24e0FDEaoB+2GkPcaCXI39aMxv6p02SKTu1i4AcoGrhwMHkVku7fdQNw
KpMv+r4lhEpqtpCQ1EPmqxRobfbOnk1KNqhgGty9bXvzdB63dyyevjZO38q+g7O5
2JB6IR5bbCcymsqXv5G03GlE8hPc1MdKKJUjNUrSQMFjwNPz9FxGGCKum3weVJ7q
GF9sb9vbGIQOe8Bo2xfvzNG3QEc8jOgW9MqZOHcQ4nM/wPE+yrmh6U0KT+wWTkm1
kolSJa/quKJvNtWaT3rsDA/kSl3lmB+n+P2ToCyyTUMOUuUpZTpKTfTuQCm/CrMH
CgqC+MSuqZ8TDs1EykivXyKsK593cEzcdWNEOpUvq5hbUP/3nqNT6CjEbhQFd1aW
32xQwjCW1a4ndZ+T9geKC2rD+4GbJQT8vFkrz6HYnDToerOTBPgtiFogJJD0VCTD
TMI3YQG2tmIGQC7Yu28orW4SFjRx63DvL/BJ18gGGK23ZWZcMxujxBb9rGtNY2+X
dlzo47IhPtepU1aNQmkiAc+60ZwGYS9Ld3WpuyBzINrioJNaXLYA7DOCmDAw489Y
Ud5IqHYy0aBBhZE0IOacZlD2PVukWS78iKyAuNTfLwekLrKwR23pBhb6i0QhGY+B
FqW1J7dLS4XRQtZ80br3lKkKEcPMurA9uhCDIyd+HpIj4tSUiKa23/bPU1gs5DUH
NerJ7SLv8czWhIoA4L7SFcBitZ+y9f8Tz+mMTONzgzNC3i2jCZrh6nLZZcl48En2
NwvR1t86QJN8mVv5v0i9OLOgpjSEH6/goeyqwKElPVrwNhogE2RFknIJlxzRyQ0f
l8B53CrBfWt12V4+hhrwT2krB/VlRf779RNx1b5g3PHw+6u2VAk04PEgHr9gukqW
jKyWnoEm8pHTwU0tZ+M80towdC55aysL4jGEuC7d5YrM+DnurYE8MBMQeN+lSQCG
9X4+3+QYbQL+2xdbBRzVOXYh869d46UIPiAV6bHCA5rfBfCCDO7H8pu4yw+0sxKX
l/ZRLlwLjOGB7fVJE5IYLxePKYVXHWqpYOZLb2/blR7JC6UeIvmW0k4oj7B9V+AC
8JnUBBxBs7P4jW2rlXhwY4gY5eNUeMaLis6gwp9P1TzByMUxLj08Ud7q2C9A6T3Q
S29zLeXXZ0tM05J4CyMN/SYSUc/TKKbfmXMhet7piOkqHg00IzlUxcRo3Ii7X8de
PyotApdvYLfo/nejpfublMciqC6syUN/Zvi7FmHcBr94JSNWZXmzwcDrLOqx/tLJ
+Y4xmsVqTOVA3dLt7sZP6zDHpMfMzVkdWUoiN/Us2c0TBLOkY7zfMrn36r8aUuO7
YCF1vzaPTPhOF8i+y5rHYwrToah+NNFOmZhlY60FNctvvvlRbdR39Z0i6tLcSAxD
z+R4bswtGOOIYsrJzGfBbaSjqmpptJEQJP59wluUZM9Zxc78hI7Ohqv+0z6tSvZ0
5mkMxo1NK9XgKIXdxtWXqE+YY++mpsMwydyxAHMSqDtixOxBuHufHHJts7evrnSm
w2iL64D1RPijxeqL9rEKBrbtoBgWC6qW3ePIUYBdNirN1lRTcsRU3N3GOPADMH7F
DH0aegre/EGrEjZjMMqn1hEZeTQCYqk4sLEhskxJxtCPf4rPJE3GOSBSgpWzub0w
akoZVh2ZsPRNKu0d4QJjeUCMWzcmmK/oE1cgkbq5VxaFndhJDxlLm9L5jLjQ78fO
cB+bbh1btEpwOGt9sVmTIbQEkyC+wS1ZXOEFBv39Nbpfca+rvVC+ezOxP/RuAest
gu5jZ/i5Ui3oAienFcXPGVtPfg+Nv/zzZlNa+MujCSx3+Vl0Ig+WuMmVaHZMMcIO
cfJd8EQwrVF+Yv5+bz5Kr762Q8mH5+soXyQIHaT+O4lhPAE6C37kmUrn1cVlPQwU
YckvTik3HMOWQYjItjwW94bVlH/STkRi7s3DXEVHwXhTDLrRyVobfHZAzi70vgJg
lGzJ8K5VbQLMWfZ7xAJRHdJfrQqGaMh5l/OlqKdBXBdn4gi5xMOxm1cMmlTPclp5
nvIgc1KRs9W+C8IwYjXrZJmzx4GWrzvor/MKt5LIZj8FYKAfU7D4C67mVtusPDeZ
hUcqs2xQLq53/SOONUMCcuPPxoVi5nVO5xcuo/o+HoRWhmY7qx8+WID6LO/jPf1u
8hHEMKczALsZzxQFVsBLqGYgjhpV8z2ZnQfauX+Kt1KnPNTp/CKcp8qiFdBYENX/
NjbheUXMb0Xt8aBqklUcPcquOohU7dN/giRDkYxz/qF+Ep45Je1fQcJAb7Nt2ooI
+SC67c5TLoIQzoiWymSgxzZ++ttniE8nuEWHo9ePDLgduBAw0UeDIYpWSviXEQyV
ekRF0fU8S0HUWQdSU9LtOtJWwu20hnN0ATs5XlUjxKQPPn2tIJhseQv33L1rD8Wc
AWxK30Oa2tR/Ejxs6HmHGXdul8OeefKLrQsw1NAv4+NjOc1pB2TUnzCpYXsRKZnr
0ZtnhTrQ/PPx9Tb9bhh54EzmazoWR0KcpDjuM/nMpJHE2rt3s5r9k5K0DLQp2Vlp
74spu/058pMAfyXBefTTdMkLYU/N1nKBVlErV0kwlEuXO3pmz+6VEY6lEd/DCRiL
9R0FpGj13Mi0JT2V7xSSTD7jcG1rCkoz30FMNO8keGDwfry77hz25FAzqqnUj1gD
l4HevklxedsZFiRZhQ8ThTXAoQEamO0ZC4heidn3kyqvFztnINFb3zKmrFcUkTjT
TpOgE1NpnPPNmCYpcer1IdFwlniwlnY5kGNF1+REGOFWLiU1T6tGagEb65bjZQBa
z8xfVrQBdyUeur0YkkM3ycJwrZYhXho9nABozLEwyixH3pejTRtv4/eLfFFSus6f
CQ6Xx1j4gHAHJcatCPk+PSn2q6C8C0X5OqBUz9eMaFzS7vqI7B7XGpMbteYZh6At
COws1X5F/JD8BZFf45narFaGKdluGVE5dsAmidfcRn0G37oVH9GkPwD25RtVA0aR
WxLYvnCJl3gYAXOQFRMJiEADHMW6oeGkhHWh+j/NTNSz3x02nkhACZG4vY8I4e5m
AgXvGgGkejh4tuuZV+An1VP/9Rq3e0ky7HS8FEZ7ecTu5Rv2kpL7IsuZA9f5Ujc5
Um1cqZdpHNSuT1LGsOuGe7KgUOfq2lk738vb0YIFnNoCX/A1ZMCbd/Zzs3AbStc3
iS/kgiCLHUp41aKM+7oPVk4kecSb3h0GZhpBMrTEyoIw7N02LysQizJxeVCxU2af
N13ScX57cc2AelD/XE0kXN13tsDmf4n5XVqLGUuDtUwwFmDns/HY7fsFR4SYf7qJ
db8EGw2B0FGD7N+xBeW+DjFt1lxePZXuDVQRbV/YzjWdFEsI7vCO32DQRzUbjAnV
04qYbaF+P1Xve+ejtIejQAs8W3md2vRf5BkVog8ggAB0Qw0cnf/Mw9KLrG+NPG6h
bJM0rJOkS8WeqD9jmsJChIXHOJQUaskhCKKZ+ffGafTAGMYUFjMr01AcajBfpjO9
oXUQdlXuYs3qR8rlsoWjm5Pzf068hfDQlWOkUDrCM+jfOrpPS2XmyxdOWm0ACgxU
xuPJym1T0JpHwUPm5OEfwqik02vcH85i8nhHH3XcRrVVi4rAKhmERuz0vLtk0yYN
ne87ZCf4jCDYmybBqXHan4iiaf4ss1fbGy9BIBvFsounAdQfRexV3M6SC0yW6wuy
ZaZFbUkCDeEST6q159U0BaCc2XZNvDfhsbQwym1s7e2Apo+f+hsUk4i1I/XZ3xGB
hgUshX1Vvs50SJsRRqjsFJ8OCRwanRrMCVZF6BGwjU2WFER3uii0h0w5T1tTuSeJ
8c2Iavnk/Zf/aqirO0H0T6Lu6xOatpxxMBxirvVK6wVwZQYG4ccTCr5CcjghfdA7
lXmD4cQSDgP4LP3ORVx0iZtNr5tpqfMb+I+DcnjxcwlN7IrTNXmzm8uhtck4GMcF
/gcgXimERKokHW7OAzM1GT8fg9Ar4fQQudfOyIi4eWH5wnFnN/gWrq/5T4+dhwcN
TYaCj25C4N1nB8B2qQ0/26uXn8XwogKlrjqr67GMTOFpy22iXmsPNvoXStCIKorj
ey5OW/OBgcOzYT1yGHH5HsfOBXjwpGoSPydQacp+lu25mCLKUJVx53Gxe3Dnt+Dl
eRdB9xJ1iGBv32KitpJbIrMqJNyp7opMcen+x9xmRGSAex4p5FgvMxQUI35sjQkj
tEGOt8xgLhZ81/AAKx0CWhtURPW8HFAr4CJkxE9d8Gbv7cNAG/CJ/YFS4qejgaEB
5TWw/oIk1TDHeVRNdERjl+kPZDnNeAdn2c4cP7vLlWXkcCXtkfgCW5SJKFhi7g/R
KEjrw2KV5osfkngxSzV8+kJmXi8FNQ9ifI3Ao1YFTmplMpidOtcIdJW+H8oG8+3k
ZROVjFVXyvwW+qOaPhJD7l2wzR0GxVigLCplSHpI5XurFuZ3Y/m3SsX+Ehn6fjdi
ZM666njvEL19yvDFy5rcgGYs/nXcvejz1nM30wWExYeW/FbptElkrhRlnWT7zFbq
xWE43yecKoBTQDvr33wkeVLux4to+NtOXxgQJ+zrGhwb2c8p0Hef6KQQ17sxJ3MF
czEPDs79BFP7HLwZoCEm/hFM0fl9gB6ajDGvbrE3sOidOfVyV84O1bU4zJEISan1
HD9bswkQXHRgTJ9t2XmFpkw83ROKMPtgKQb2OR45ZkwGKsubKce+sxPA1pnWiAr/
rhyLtdTr2Hcas43KzF2/DR/qyFG+2N7Tx37tl5Qk963OchJ9jYC3J1zw8toxancE
pTehNFFWDR7rXa8HzGyEzYSHb/kc2ZSvAZWw6f83scPbAwg9pP15OyDv/uNdULFA
znw5uwRyGgSdkz9x0jgyQgtSm652StxIgPOdGgTrCFX4nIuc42wQpWJJOUzhd8SH
vqivPd7jkbbzufzK5oj1MGeFKfy+PhN23LOKOPbvi2LRXMB65AR/vkqMhTrzXwtn
3gPGf0ptg8nxM/vazEfD1pqjRleISuxvLeepGZy1364GMWZ2nyaywbEMExoElWkX
1zuHdr8NbVa2d1CHWzigF4bk0ULeZhQnAPNLWWR2fZRQGjXSdzYMTJZznVXaIrdX
n8NHKqy0L49AmAZzmSJrUvn4+7vVvUQcVJXTPmgN1M1j0l/eRemmApyX1o+cLWex
s9fcMPZDjMJFFstOdn4JQ+O1CvQwmccj8r4M//LQ0FtlwrJo+7KSCZ0V0yKEPZRv
Ld3G7/E0aKwh3qj7mWefEukd88Q5Q6FocTBoNLe7UaLpU1bn3vsue1a/5pxtrudq
RloKp2M1J1ClmqKmZFPQHsvHjpbEMMQ+kHJMpVdpy6MLmVh3iyMQwwEzOwTWZS19
L8xYfjUIW5jUFiQaHwW0jN6vk+UcrK444EDfpjY1j6ZWRq8Tk7vwQVKu+H1QqnAC
uDnMRcU2yBKbpnKCH1KGipjZipf0Bv+5sCiChXPCCbffEpfhAk/fVSCJ6NSrWuQj
bes6B+1PQgpqKWX2Kmol1Yvtbu++3W6qgdjohSwcpARxqfXsHuMcPLQn+48eTSss
ZpbJ7LFRe74JUbcxN6R9+zZC0jIE724Io4YDDW8cFvTnl8w37GFkeO3UTOKSpvg7
OguoalnKuE2qDDru8iQgNyDyJycIdOli+dMzBVqo5/C8SASDthOwOtx2Wlf2JwtS
QE1wuM2lldeZReHhKUKJbBn4FXpusH82OOjw1E+Zha5G5LA/ZaCYHWRllj0DzAz2
oZUu3S3udgEXiDKM03bE+yXanjw8+mi2A5FXRb5GrWZwqAFRHkyOmQjfPySgjmK5
yLil+ZiA7qWCLz7r5XctTUtvtFk0L1qIZ/F9ByRN6JtEuXoZaY+Q4eyLODQ9Ytxc
J0ozQYauqAtrw8jSvXhbHwHgQHBLNIf5mO1L5kWgmmhs19F35A3G7T52QdnAUigp
kP6VazOvJPr6bJConIVQwofjv14Ne3FFYSA4PKSTUMDWjjJFInxt27nSBqMyhu1s
5ApWd1O/mFPMKrs2tei8lFWn4/Ft0MwykbwEclFNDVBeVCUJ9UlPNiHjyFMHk4/k
aDqwWxtvOrMNkWCUgvtrXjjdlN5pFiWmSng//SfDXHT+tg6HkkC2zlruE/tMU69b
+e/IzYSYsVQsQAEdRcuCa+jfKrb/TbHnqOkdenRDx1FM65hZivDWOIWpdHmWZHDt
wU4FyL0v+YfCjd+vwsyUmco4Lw96vEMmp1CpYmKyAro98D4uCgO2Nzq4miUYbWJE
rxEIkGTV2RImoCTk4u8lzlkWtCNvC+EfmYCvvDDIBZYhswl5MerTLgABWYYCcvvQ
8CwT1T9XqcAuFtM2wxo4dz+or1f7kH3anCjMQw3qaZj9a+qRKVBKzFXA17yyoTeS
9MTO8JVQ/D9vxnJnx7sKR/qVnSFdikctCEkOCK4jt4u/nwhFnI98osemFO82lp9q
CjVdXigCWI8bgJLPLyOO2cZ5/qZ6E+BYoM4JTZd3ao0ZyJUGtbNZEU/S+lJ2FDvx
PGi9xqW5pwrsvB9LKYF5ugIKGGFHSgtGGlyu28slPwMMPWkX5fK5yp1HqtrbqErh
vflNuDihQOXftIJZUqmds09s6XL2Cxs1NZKnend9aUKttmRI7dvxRcyRgtnbiyCY
71GGOVXB+s5gpxkp33m+WWxYTT+eYhBt/be/sPbspDnERk/dYavhUbj+YestvOrT
g60zEBLGoONB2aDAW0jmCUjH9bKtLrrREEm9ZvkgPssEsUC4wBW2quQvtaeRm1YC
qJKd1O8d+IwXSoTN1y+2OIsgJ+uCZddA+YM4sjDGAppCS3q+Y44wT9sCE/K5lNIH
5jIyVtigBXJYTRMVPRega7lnIJkfxPK5Z/wdSUEHA3rx1Mcct3RU+C3U3Cqj6X7o
tNDWe0jeTX1zLcMbC5pDxVEuLIMGE1cOz9K+YUCOLDYe62oE7mqp/SWJ04c2CQCB
sWCQ/AHTPqswP7aX4AUIAQIXTpHGV6bB7S4hU8Vd69hTMpJnXnoW0FSflhnVjHkz
aZLEK0SM6e4srA+9crjLo7opeXMQBjZvlO5ZCpf4iQ7q6iS7zVRpjFOXxiqowm9x
dELX3Y8pPhv5j2YHQp/9i8TkeqpR3gfet8ZQv4QXixEiVgV1cvoz4O8vpF/xOG52
B8HShNvlLgc8wggD6rE6fJYRV26TJytbDpAOlKyrCgzh4c+J9Kskjw+YT1R0uGsZ
UCmI75K0MvNGKDtH82rtqwkpzKSG7PAgMrNYVLuGHREaXH4vPY6cRH5Qfe3tkyP2
/P5AWtUzK9tSF2VsHuHVLu5gQPAnE/UI9U0Jlugb15tTz8wUN2ku3hLv53uF1PrW
+tbhY5fe0ZxluOCDyfi3hWZrcjJ2mvoRxAX5afd9D3ndDsKSqJbE25ABRi5QU53g
INE71yIq1m7wI6jkAKQ7sorpgDsLmF+A26kIJ30cEQx7ajzROyvmqFwC0RXnZoue
oWoFYqNaPT/4gdpMplBGR+zlhQOXU6DkUy5JvDt9qcNFlHYHaSSeOTN1IJy2kDRh
oRSixfDHSsXxCCCxIQyuCWdId6i9uMmIGySipCRsHU6YUwuOLoVA3iCpjVow4IbI
oHpOdUb7lt4Gw5FSUZO/nsa3q/fU+3bTIUcO/5hmkO62t1qVZZzmuj60urngFqvi
5WIjKmWSm7jm6s8KjJ4yqKBuqBsfGJbkbMrkkpdWrmECCcTMZwwPSjrD0KYM9kK1
T83/1t14bcjW0LLl7Lk5KJt3tlXyk57q1JkmJSXwPvZsDicFwhl7Ar18ZQSIGSsB
Vn9/sF+yNgcHv3G03F8jhmCZL/7YtJMNvFJVUXVLmtlwpxqOaler1e7+Tfi6HRAW
AHgfl56V+XIEVy7LjIKsWi4q1A9R5wePL9AUDCTnrpdLUUFbGxM6dQViHgC2vUMl
b0sgJrcs37PsNoP16AhAqWdYcahhb04VBHXFy4Tuw9kFfoiTgPXfPBVEKRkDSv8q
2fJ2rIIJ9V5ryAcsf71qh2h1VqSipviWM/z7U/fEHbtzi+fIBwS+AH/cNt/MxSLm
AA4VR3klovUkMFfmcWvwAjudmPL0D1EdUi4JSeyMv8qH+EctphyjOBHcFZ+D+if5
TfhAT5huzwSJyj0T0B8HcVTV4XBcs8mosWE3s7wM1OB1CFPsROVeEn2w+QayMGAp
2a48y/k0UqyPQm33RhEI1n+SmegruttdN2oF2MFdfCtL6zF8HlUo9dsv/Eopx/C8
13i5DHo+WSaGqDD0mRH0yiqT0tR26LflJGruVca6URYpGZdvALCyqmX+ViIbIRmN
aqE+P7v/nm6XxiQe79JimmRpBVq1Z5bqvdhCf9BdtKWuLT6xU7giyBrJ1sH5A70H
8j746u0AwKnd8xS4J7XK4P2p+oyfzdPjAlP6a+o8ogv8Zsrgk2DLgj4nruDOYGGy
2VuDQTbhQz9EjDCOt/8QtR6681dxuiZi7ehn2J369YzZYiTVnQND+sjgd+oCyifn
KTMYU5OPQGNCn6+lXv0pwOQZhiEWcb82Y1EGOc2Pb6Jm0VQAqc30S0VoFZtcizpJ
wMTsSuwcIzk1lXo/wgEU3RrWtTwdBfZHnQ+Twbu/qVkohFdAxZPSAn9pGLw8EHro
lTs9JNkqP1q7nsSCwDzveCLKrpg++4YjcoagTYs5DZpMA4EuuYMl/3G1P2SjNXTA
xdL+Ey3TVLXS9Rskj5tNjO7t6gDNp/EFh/J8+3l7ypI5To/jjcm39IGweP9r8t9m
/nmRuTD8/mRJOSFwSBLzzfQfnx3Kh0Hou10PCeTQOvGxCQSMfw78JiY3+rIPbTHR
EOHKNYJ85B8iCdUeAjDBoAfsb+Vra+sGWjw4UMGVu+foZk2BqyMzgPi1VSqoA2IZ
eAZZKVuDiN0ZqSMz96gGc7dUjIJWgzyi0R0fxV61imAbwO0uu+X1EO9UwB2pNrE0
9R3eJ/5WaagDJRTg4t7h9aol/wCzl5pvpv2jt+qTsRBr2Rv799ZHZkosvAfC28ex
+Aj7JR8njsNMcLybZpFVfUVYjy/RyIiy7V59JEGbm2AN3JyYiyTiymAqyL2L5qM/
NXU4TFjfHGxoDNOFoJ+uKNeouOSB1tWDvrYphgvddk8tfF4UHtzikKtrOxu76iyI
r5LGtuzA8reQ6chDx5g/IMxaLeeFFViFX1N1cHM7LxAiRHlHVWokSAPkC7Gbpi31
B08JD3RWtihUj+h9t8mHvVNW+Hdn3BCat/ZY5MZC4gRsHIdCcAoHGAAmZAmDYLA+
wxC5H5XlGGhXQpkUd1AfrGyfQlJXAJkL+//uq7U+Ymxz++6W1It5eP/s8suJjfwt
KYFXZe7vNnyQ6j33Phpe4h7XIUDI6y0v1mrk2fTmXNiuEdYwIbpEMhbZRKpelofP
d0yEmuPbbt5n7/8M2GSuU9hgIbi1PBXHvE26KQcJpzklG96Kh/GPOVeqI0cj9uyj
R/HltS7R/BZlDzd2Fxv4Ivam1PTbkN4MfB7ddTcU3Fe3EhPu+f061ZekEm1mOGEd
0P5JgfYX0S8ZQ5kQWRT1wQ8MuDA6+OKg9Hn8dVe1xNwDz/bBgncz+vNqZBybH7Zq
N4HGwskKOsE49m0E/1mstIF2UlAEbve1dkPG6uxNcHQHOATjOvQMe5t/rjlF+6ly
MKKy5OZ0WiTuhrMm8yDPyBgccZD8422akWeyPDCAJkhCkE/Rd1h6EyBy2ERFDu8v
gB5UPTNJlKBXIRmFVfNdNu67cpxQmClC86IqcE6+jWU3vWpKDNLf65HZQPN3r5M6
/0VEKwW8O6xc9jztLYUOBlBth1L5UhKmNnerSvavzN7HmiqbPrwNqsAg7Tqz7Yew
I3Ec7KAtMDfau9wf31/OtTtcjlDN2JoUm5VNeaiChutGKDOvta84SXSN8zKYNtH4
1O42xkekkKNIGdRztStmUIYC4xBgX3FfUx/QYKMES3Au73mKWbVD/eNZLGpHMYe2
hy4xADom5JVahTl0SqNz2JeY88PvtmL4q202QFT1GdxO64lZIcyRCVkwlTdKA1kx
z6MkRabtin5QL9SFjWk7ugKHajJafbebFWPdOqidYiQTA5vuu4vXh08pXz+BIy75
tF9hoDhxV92wtkGnmZ5XFaNu5ek3k2auD85gBFp0SEHI+DhbwgNkl7xEN3CHUXMb
sgsk+xeXcBvOLApUBqRNjrl5VpiyqhgUHkfS/eMQWwJGOBqKaFkcm4WWnPA9TpX6
b2kBHFzDPaJit+6UPwF0oW79ji8dVQJX91fQzooGFvlQc6ONwJv2wSV/FBkMB8ni
xyH282OCP80w3VmS2HMhg1pWaI/WY+ktZRK1ebnnYaS2mM9dLUQd8FdyoL9trk5m
kEwJmDa2QwaAnipUpn+hdKdw+6/mUVmdGsOuYG8ngtAz1eCd0HX2xy/P3JFLE40w
DGw8w8xHGaAr69ca6RUkAkS1oTnYwG1AhZMtw4W1TiD6Kqfl1+omDIUnCbDD/RWh
hTDnMZQNqL0nmlFq1rfnCoXrRRq4hogTubNO4QVY0tEckoQHzE7kai1mG+ZXKNbx
8fzFbyHy8Txth0o3qDYJm5uLduYYAoUGxKW58rUIOdseBWtrMN+LXC21J5se3DGB
PG1J5nK8F71koEuZlJay015Nvl8XIum3dalf7v9eEHT5l72c7VeyH2CWGFY0IOq9
FNfMbgK1aup9ZcvqE+d0QyX3JKxH6wHr5PGUS6d+im88DlLcV3s/gs0Hfv0/Cke5
HhSGI3N76F+xM3GZZscITIKeYnkSFlk+3NYwiYC0x0doddmIs6uPI5Rky9yzJdYd
pvKVx21p4DlwrGb3dw4yCa+aI4Xp0SX0/2R2hKpl02J8KiBBwWJNjsjJxEOWiAbi
e0Ob620hJexRJmxhHYugiIN8b5vA560mkrGH9lyzJWO6lV2uCRIpaCimJN5djcG6
/ujdzICcZOX8VQlBQkQ8Zf22EeITo99HCfWm91p6apbE6aujJtqfV+Osd34S7oqg
7YlPmqn1XAn+RW7Y6+jdrwflYPC/QF9VZYnYC5EeE3wsr+pJWes20dtYVC4PX3au
qGt1RBlVTMPYCP8hAVJZQ6NElcctUaXm/F35CYOPvLnBV6qauNtI3/D8EUFRBrGN
zIXwVfo8+b6KDnJG8T6tcbaSD1Ravtp4TzGmU2j8qKGqiT/UcFf7NA9wPq2/QEi2
Ygzt0ukfr89thcJBGqYDqHmcFtVvPnZ0zhPdxI9h4DyAfPW0WnxejUJRGgaMS5mb
VqIHTySqpabqIO3gRTW3kt0CqhLojhDRSGjWklkmPpnPz1QdujpDULatk/5iPv7+
A13GlBLbU1lwPCryvHYu/SnyVZq4o4ctj6ifJTjRtBT4lbnOsJwMOE6xIymxS1Ol
70dmx6dBK+ZZ6Y9at1NxFY+rpAgVgdC6ALkinnNRrIgs4NoFGUfvK4ATmqZyy380
vDTH1/lUj6qpa/rh00Yjm3QuB0y98Im/irdEpBXnA0H2ph2+3YSgrmJlUAK+Fjcr
Ru4vqflHZtoqmsAKjQ5eunecO+xsheydQSPbMSvfglNxqD1b716gk3X0NxAjV9zD
8yvSWtXYJIx/k/khVexCOhN9M81/rPeqx55LaMgM33URXolhtnMCdupjy6PKuFIQ
RW55nWnYTVIErzXQBOSNAyihECJthHff2RoHYHsdyyoUoJXOSadWAHkMfGKkcC5d
GIwoaOD/weTIUyb/cGjScV/N321bGrV7CXnmZejPhykNqwFB/ph81aehEcqjmyzn
99S7Z0puGVla6N1S8X8lJfsDAkAXbBaRDYwpgzC3zdNadOLnLkRsYOvwYubcbsRE
UgFOSHYqqod/iAvpgJ33kNDku8nDquWtXrnm7BvQZltFYjvHm6kl0S4FnH1erYTl
fkKypMOxyDH5DsYFtat8cJsQLt02mZI3001lsV97U/yX643MZDvvcduY+peeK5Y+
8GVwXKJtmm2bzdZTOLx7E+tGM/jLN9zUfYFY1RzNhP6X7B2MJXXcX/omy5RGlY01
dWE1dyYe8COfXF6ruODDm54+hTjukz0D+lcvycbNoXkP1huVvBAmDMosTk1CD9tu
rFXwV2yB8f4hrKUTzcTeq1cp94ToeGrjDRVkB2ZqNmTkTl/UXNqav7z7kyciM3gG
sBFL2y7mGGoyQx7X4pOcI2NIkvU75+NC16INxjo/0/h8moh0miIit6vUN+KzFpoj
2tTToMho9zyYLW//YqURUy8ZM1qN57EAroadHiaHa4Sa7f6YhMjcuS8x1zqK2dB9
YJbPqO5meteuJJOIISVBPlVxQ0fOP8uk1Q2KJKU/fkBg22CdcTtpqgbVir38Dtkq
5Pbo1eB58LueYdwuaIjCQXnk7XpW76JTOXhMcKhtE+e6pNvuRni7+jDjwjbyOVUG
Lcc7Ku8/3jSwug/eiId/BCG6MCpAhhPmiSutPR3GkAeySLtaBJnw1aCI2xYNWBjo
QDp3VvmfbiEnv6X5ZM9aG1wF2BO1rNR11vzZfIjXRyBNh+IArFi9wF3yq3+6tHB2
dDsmKxVtd1ncBYnpSfsUOtGToH2QrZaoXPjaaw5C0EyjJAG78p4n311IpyWDOa9P
RUtxeHllipU6bTdzf3wug1C2kvHYtjiNQncPBHgm6s0AUUtMYaqGMybmFnmQ+TBv
Pw8SN6rI0eCH2RC5xWabotN/uJlHTzr/cWekNEyvstkM6ci301orQqGrapzp+iJp
Y+sKS/J0vsQY09Hu0Z5CP2i9ZhUA9XcM6mffIrlk280qwNqD9nbxKPOBW5gW5jCX
pY2XrCict4IFSSuHg2ToLdeuXhVvj8lLG0bauWo/eHZYhkTdSUYRQj921ZuH0RbK
GcQ8UYTKNRFXNqT6lhF9vdZaGNrK6eN1waIz0eZr5fkBKQt8ln7gMsynTEtva8yB
UO1EAWJnyKPQdli9aSIFquxSkvfKuwjeIRhv1TnCWRTG5SwDZ/Sbtm7IA7rWrXET
yd/mLAieho7Yeas4VUna4HVdWFSnjgw7eN1/KGqoXD22Hjx1zBMLWSPCc+o7FEwY
2TLIJ3N2bmRyr7s39g0BJ0pegNcMDCqmCgFPdByfAkklqIKzwmUXTcvjylEQ9kJK
355EtQ0sl8ZGZoVC9oW6TFFgmhwrn3Nfm9V93SfMs2BaKnyOk+yUvqEzrOxZibU7
oK6HykUFddOd/xFQtOK9ivhSErxKa3TR+S/klqhh9QvNM9jIpwKBTmdoOSg5mbe5
bUmkQeTq9qxZksYKzGrQcA2ep7V+TmfuCEpgteu9s30RyrEQKJs/P0UP7B/upsnD
yc6lpbdKRbsOTqh7tRIIT0nLM2KqCFbckCv58i7vQcx/Jl/0qzjCd64VjeFFS8mj
KqhmZyRQIcvBpzWOnkATSacpscwfvnYJ1Lrbv5h4XlL3DWiXZ7sizfENOGVo9bOx
49hH5qaestgFOY68C86HxgD53JpQFDNj6NWl7Qz75AK/akQRHG+lsRxcACXIh11a
nY6k0WcX+I13WYny3174Qmu+vhmwp3knb+qSGCm+paddqXzOZko7tERjlYOwRk9N
uMp8/ddx87M5atEulX6TQvxE1xXgUCGJ2KKCmBEgG8SsgcTL5OeSbEOq6dUCoHiH
wWJdOlooHUCLFZpeQKLbx6yBX0sEFZS27/zjpxDd6pq1KdFKZhOX8PsKmYWK6eE7
PJABPvzOs5aEdYHMLZoA11xoa6FsAfh0IKmR4rvA+plo1eD+V02dTz9ABLPAyTj7
rTrGSEpwustEj2hWmMf1lkD2jKK0Dgi6txcKXAnCo1rMg3LIjzTr8Hu4vOKyFA90
UhKADWbi9HRGG80afrtDz8m49YDNPKR8uIiePz16ex0ojSJJ56teVRpoPgEYxVhE
k9DoYv9FX7RGHJknLzhwz8PhkQEOZ+HwlfGwepqQqRk/1f/PdvS6ZT0U3Li5qOtK
hk/cen+pwkXs4xRxuRb7kPt3vntzdy0mY4YCH9/cZziaVIWF0kPtzDfmthLsjY9q
CbSWYKWJ00SEPVrAdp7e2Xa01hXAUI5W/JFSECGlbzZO+ovnllrMikm5+p6oPi84
7zbbVCaHhEuPzJ7SSZuScSoim2EWkO4YkmmvL84ls+m1A+fut36WtzYcRrFmKCAH
nusw/pMnXJIVM4I5HF4VuQKf+W1gKgYbDgPaXcqSZtsfZrFXmaArK8nBMAyhAhxF
6+SW+JlzVpOknymIf3/jgo8oOzBpjbbbHnQClzX1M+FfDrRkmy4ZS+sDtTgZWkuf
QSrP1RFxBwUi4sXsppAizj0l3DrwNEA7Teg/iP4lW3TsgLHD91UEFtL00Dc80wen
NUxb6JuEC5rebUCQngk/N7JSFQIsLziBXD1RFtyCzP5UkIPj1pVwbCvJOJ0GX75u
mVUOX07Cnv5bTeAx0T1edfAKCilXX7fKB60z9R/4EEDF61PtlRKKuEWMT87r9oh+
Wzl2qHP5w1PyGF4A2gn4/kaoyDJ8cBsnrTozOcsZ1zOIl9fqq5K6Lx8jqJss1MEs
rPccbFpokkcG5O9Ym7t0Bt75Oh+2hhMu3BtIxT8cn1nOGl9cBap1nQAyvhAlMHJU
kCnyPK7drTDb/xjWyb1g5oi1O0p2NJz3zZjN7uSR/4dHjLfrQeKOGPJ5ZUN9Z+Zo
zJEZBcGBR53tA9hPXmATNreipCTTQf5aCv+0SvNlcLJ3X0wrWHpzK7ozuWrY8XP1
KwW1zsl6iZfTEzucXMdFm3hUKe+HN8wezFDd3YDhe8RfEqxJMeL/RSDTeoeT/Qdk
zeG9Z7UrZbD7U/DG1h6aQlVTx1dtT0uhicwXqiTAh/x6q6qkMC6aMEMLx/v43T6Y
nAlGgfJdraSZrMwdmbeb16+C3eNPc6hQDsPUOnKOpYIuf/jjZjPNi/kkNUdWrYxd
c960YsNWo8fOgBursjvFacc0/q+jRP7X7aOnOnk6OBdxYpZaoiZLcGPvvGpMOcb+
Czi/IJ2wl1LONSqwXyfijnfaZ9Ek75VCgNzpVpZyDW+MMja6ZhJQN/WbeRykJbla
FPnHkkhsifeWejL3jX+fgSXD4/j80yQsgNZkHVPB0YJZyzli8EsSk6U9JaUORUcH
ykU6tZch/bcmu5Yr3mIaDARxNfXIN2uzBvmS1xTBeoxVJ1bbbBNXMlxbgfD1ElH2
AR6UgNQ1bx3ijURVir9YBBCHliL8NOOmOJlVBIstVTXnDLOOCjmaxtcRHQf7Lj8C
DO24XPlT0lB842mCKJHam97fWiDSo3dlyxComWvTKgmkc0hacWxke9XhnRuzQhvZ
JvtL+5DVP46ej172nVXomyRviPz20yb3rBm/1ZnAkO/rCGPXmhKSGUwY9ZFLal1n
kzYbnFLdMeXizx5QyvAg923QYW9UaNRQgP+97A/HKu6BouVyYzwcfJFnpjEMNI4t
zl2R5KjJe4xY88+M3sSSg357a3O8mVlKd4+8UAXWMC9VHuxng6V49UyKZnZ31dts
BOnP9VOE31gaa7DSfNYjkX1gnJU/milgpt6vxGo0MD8cnsq1X4LFGS4TjRT2n/9A
jInPq88Wa8riFJfnQZh5GwyhdPwUBsHklwThA+jX5BwySV18JvXB3WiSWXDGNs/5
uzwuZFJwq50Ka4dvGPvJ4lq4unrPnSvXWQN1KpI44FqD3nd5gAuuJFhv+oNCGNFs
kMQ0f+uV+nZoUPE1oWvB2PbPNbseJZTNR/HJgwV5EE18xqi50KoRzDTq4yu2CosM
lhVi4kCoe1rW1b72XwqrnI/fZQKhYbwiZBX1VE+dpW6RheDujEX3f2PqiFKRfABQ
WLZuiPMTgik893MRrrrYRuH3KFyzNiva6J3REDcpFQukJPxa2f+rwEkcDWE3gccS
+W2AJS0NuPXp0GGLxKKNebs9yIBBeDrUK7pJ3hsindYV8MzJQkVq5UbkebDcOp2Y
rKdF1/Tqv/oz/HD7sMC4Py2FOIXYOIOKXbbPaug0AizLDw/1MtPrFG1p2+C/uv5n
/bYiVwsrtkqSmQXQHR8RHgunehcqbUvlsUfFmfjOJIGcLQjE1qrCkFKFksNJCJZb
LgMGZ5xPq+Z0Y4LkTEWyERjrKOuHahWbLdIKk13fRerj8hDbBFiaQeNXz6HymaaI
uzOX5WDbTWxmTf9DEPLg6BYF8ot7Suku0GIelHtGB8huIj7hlRpJHCw+4S4Pl+yA
1OADrAJMsn2G1LnNN8XEyQw51FEAWBf4RzpGzfXccXMP0ktGhVNJH7sRMZaFOBam
d2J0tGwj2hQCj+27IAVycYghjtZE9uWpf7ngJdonYZDixmfnlXMumnbu/FXV9qXB
knE0tCSiyRsbFv1nzNHmg7f5Celd6/PBzV1FE5E/U0Y+bq15/m0zyoANQ7q8OyJz
wpZvVeE/OaK0LuUFrd3BGlQpkx8pOr7NjolWKOqSTHUILMXBh4FZuDdcl5oyIRfH
nG/DTWNauNf+LD8yCgRoKxoUBhMdViwiQMD/l42YBSuV/CzBvNFXp91WlI2Mfx8Z
wbdTKszYT2O5GxxnabmijHi4BenzM3Oq064e7lrGxVxhxkVOQ78J64S2X0pYpOUi
w8QNCGXNUb+c/zNfrp9xRVZqv2IkMJ1Na6aMY50K32MMySPxhBsZZ0iECyJCwhkM
Cgk/o02CIX3gYiW1opMEr8Aoh9BSnkA6HEGsWGvQBiyMquc6BuYwoYRHQJfisVUV
j5RxgaN/up1Y64IfZcF8nKdmIYxD5yE4fEBwIGwN3LT5iE54EdWNYQI+Wn9aVHWI
VJ75/+IdQPQgidfyRhF7V/b8ae/ArbvlE80znLcnRxn/xPn0tIv1v2F0R/RcUv+z
GUOyBEwWBjD7jmJMj0YsUre9uSR1kbP7Ju0+vzoj+RSDem+lXe96yCGdjltO92V5
N8qadm102P1TzlUHx14LnCwk6F8Cp+cIw+zRpMFqX+TanQS4HXZNCYFkxePZuFh7
DgggHfX3HmQMvgCXfJB/+rgo5jxOWZnhpjbXhZHuhqCuPxD6UB3JseqX4W4KVxXJ
ureTP44izQOIz+f3CXZB1obR/L4R2KUWFldQzSYQ1NMJ77wcdlr6yHwi9NYS7M/o
9lmT29A+Yl6/dZztZ7XbfTS8pGDYqNRuWpSTSUWDkR4vYBlB8XAAztuciL9ZlDNv
6Bt3EFIpIBRYjyG/Kavj0Vi+JgHDmwApFB/hp/EvXBGzpZtXJthJXNZsrUFhIJ4c
u8zddfhn2uC04JmMLC/FXMwrVfHbmpFbuvGOczrsDfy5tGOK66IgCoSSTOXtMqUW
06I7xZDMl+yF+6Zo6uxVKYETqRSVURyyCjrawVfzNV88ufIwifQJBfBlyzoyesXY
v4KsY5HHLE1Vrfo0hwYzwna2UWfoK06dUvLtnmNTgoq0Fvcb4Dx5Tia+cOe7Ietq
ZZTOHOZ23Azt1FCwB8Ywk/x+CCKCbmBsVANHpUBvN6+oZmhQaT3qOyyfXRQr9MMv
4PANv1CteOTm2VLekl4ud/NlsiOUMGcAHQjYIaCiHhcOxhpSNofQqTn7LYa+e68l
RZPhDOY4wUMqsLZK2AsJjdoLzht2yg8+1VCWHAidKgp/zx8diAUlxHzM5A4YzmBx
rveb3gfiYhbRNoG6QTJJx/KGGLqMQN4P4CmfSHhbTDW6/VJGh6YnP/7cfyc226QC
zbBxm1JV6HdQQiiIk34ui5yxF3tlpLpMtFWb+nBlakljxxqX3KXcuBTvb4Ki2GZH
ahPvwiJq68aN2wFvhYkICtPgWRKGfwhqFqgD1mkPnx+G0ZiPiKJ11n/mHe92HMC5
Wk7GGSaBDLDXgkNpv1AygH5yotkt9x4PmYL1lMGKnaNjkRceF1oNc5av4IjXyBPS
xKuWKM+9zXJTdAAIijhOKMa7yV6/HU8EX6MxesZdqhlWchILHPBXjdHLsXQ8uMoP
GS+WkhoP3gnxNCVhcem0NiuNJi2MUUW+rVglmj5lOFZqH9NRyaawzhdV0Qd9jYCZ
BM0nVAsVx89VuyTJGmGcbRQ6vdv6LfyemqLgWEqC//o5bVdqB0v7UsGm/tzBLvAA
0b4+x0xXj3/ocqk9j6dMjttUbFQ+PAVgJSu784m2kE/6vgh7U26lOxiaip6vmrDL
Wsl5khPl9ef8BF+bCNpZodLc78NS+FGKDBAGMwybRnOmc9XnnND1Vup8YUnhHRC+
h59pIvpl1sjNnENyLB7EBOg8vnpJudN1NLua7xUP/cdIGWga6rw9aDtieUTEOL5i
nMJs8WuTDwvf8AhpdS9EMTAZSgYiz1CY0tmn+UATniERWQRuiGBiN808YMGNZxii
9A40ujf968LoN92DRiZ4UBhEV2NUc3GmD0Ldv+fOASZFi3+p+VhijXFwBQJRg87h
4rB+OU4bypR5FQFCiU0c5o1likuHY/5BGDVfyReFH/jpr2sRVUh9oNuZ4rbG2luz
SGihFaI8QaOtBkjfU629+9PepS1pOqOBQjY3bUS8+FIXyt8dMRXCmxUqAiMxlPj8
hYP+RmnE22h0/9p+plHZ0WcHhk7OG04vM53EmiIoHoEqTkWkRbR7D97C1liAViWL
6Mqosmzo+vVtaliUrlV+zk9SGI5FQeW9BqiFWFAd2bmOjT+ONfOTsLl/m+FnuwV1
JWk4oPu1KjWiB4EDy873uCRNPLcPaqJc7Cw1Lt9Rz3aB/SrEl7ACekQ0dZyCPMIF
t3R1ImgVKOA0LeXcSSnE7bi8OCwA5E5puhYtBNuMp+rIHpBto09likhRiY+AcNVA
OLmskJ13wqskih9/R9zdUUnE05eAhBUd1Bur8iaAT4JwOjfbsIL02wu73Bddy2vN
y6FtBXOv+VvWiEizqvX4URAeqBR5eCkxvDD+hmXhFmk7unk/KafcWvax1FFnnkQP
1XGMz4xgqnrpVoCD9T6Sg0Mk7Gh8oGNPElIQE2R/zYo5kjocqnkOHXenyC5MI3P3
xGOiJ37BUOsmARZ/dNb//xNiVYpoMCfW1mB09ZFwx8NnZqG/DPvLNl3CSg3z49Jf
IUFDwyxzd0aI4UpQ2QKwphy/gY67w4ibTlLW3qDFeS69nOyuWDAQoFRfMcpaiWWO
yQpHb39CxdggPjfM4Ko+m99q/BwVbv0z753WJmQ/AhO0j4qSAz2YyI90AOFyDa3V
ZzuTXOFUjvg8WpJ3euetvtZXxWYqF5vVdzB10aqGJcZdnpU3q0pjrmO/6YJPliiS
HfJPbc8qnawZIMJ9r+ZRuYWlXcnLJVoXKLPL12xaD9C+iIdYlMoHz+a57cwvuGTB
EeMAQsALkV61BJhW7WTyDkdo1Z/Rv6Imu4ninImTKGwygayI9fJI1EXwV5C1d71B
cL/jbnK4bOryqlwQIGlse0ONVkW3wm+mmBnO5VZBnlpENXeq9BOiD6eGgMjkJHFY
TKg3avs0nSomQzIT3c9gqB8+aMx77xMWEs/M83D7SorKMm7JHefU0Di9ObRsKB0D
7un10F6dDb0BaD8Mllyu1rvF7XygcxVSJH7Hn0aZuRcGaW+L+yq2b0C/PNeAMNmL
k1UrZP7syGJR/qnPUhPEYJn98gu7GxjSOC3dSUzmvzGF7n5MvB7g43klYZMYF0RK
q/TEwERL7/EffAMMvxWkH3iseud4xM/yx2+UYxC4aHOt0bQmEQI9IDJJFMxjEI4g
x+TWvTZk2nRmP07FtV6fjAQG+RcNpaUeBuFdYoJ5CC4GqATdoquwFNL4uFpM93sR
oqYeO2F0HuWfdj3Am6QyGUQ13jZRJJ1evET9B7r5ckAYF9IY4AnH78eWlYeq93DO
ZHOaRgG8OO7o4dthnbQZUS4Duf9GjhjyV2D+yTA61mjqOFqzW0Qcrzm4G+bSUMg5
Frqrs0jCgLaSPbSTfwdarRg+8dzd6ZqzWsHhPLzgLcpCbadhsHLOVxBR8X1xWF0y
zVbAfOv9UgbjBaQSjVgVJMmsZUsuAf9zj97+eAxLI+7kB2vVX0pWag5gspPBBAz1
Az+zaiEnHPBEn9diXa2vsI6SmboOXSlFubahSH/9mGSI5seEobZr7JvDXzZJVNDb
fkzipBKQCXOX0sA+Yg6DS3Td+hl/K5ctA7qzyr96PE/38l6AdOGQPvb0NJORJRpJ
LsViudblMDzvVdwHHgP9I8erVdZucEPjk8nLa1wtMcE9Jd2HwjhMY5V/LA3RkTLN
zOnsazKGU8gCggIVFUuxf+YLEBlD6xcDubeOsDNGsw6qmdFbxhGGqFHDGjkzKbbm
VeaTTloWgEXIDAfQ/5dxfv0yjjgmxteiYc3NSEotuBaE+VPx3Zj2Zc68eL3SmzRg
xm2rEGaXcDzr8YF+ftQ5uGUGA7SZOl5RtdwlJcDLlj42/4vwKrQSQr5MUM7J+ckw
ypkvzM/NBwBoBeJ0BpE2zymTMGlAseeOTPi/ubH7Toik0Vfru8gGZaENLKqn/ndy
mI2+sfoxSQHgoFPzCVMlwIMargrAYZNIuFM0xNxtHZ6MAQf0s99n0o9PgZSm2Pq8
N8VqsSD8zpPf+Niv1noNO3mHRxAYSu8HJeFz2wB9imTaiPkMfj1QfE+i+aSW7+Y0
DSpmhUkhVWmPi8aHn31aQsnogj32n6O1Vo2goLy76hdExHa6MQQvECbjohfk9jUn
pNH2BPg9TYmCn0QIjIiqcnm1+f2Ow4k3oCwHa7JWu0WD4esFgCW5FU2s8FdQzuNl
L6o8iIRH2+iUEjO/h04Y1jvyN9ot+ZCUH6oabp9YnGBXVyBUFIJMTg09Y7KucKOm
XP8m7hD+flcH75qOeP6N4Q7jVsgZbbdqDjJiOuer7XaDuum+Inj4j77hmRwtV20h
SwRNwALwaIOK9p/rxhh2T3UfA1GUVwXrZEwLVNDWbJPKgv5AjApUCt1eW5NzkUnf
nhnlVdPmyn/EPm/qeU/8kLSBMxRXIq9jr33cZJVEF8PDbG0r1zwnrrlnFZucNFP0
O8RDIKugEGQDfFA29QWm8q0OR0mH4z1Mp7LguVs1jIlEl/icTYJG5gezGHtaI6Tp
frNPrn/VvYsderLwb5YxxfFJbI4gtZvUG4bGlmuvxpKbYcOvzCwPFjukdBLClMmd
p+na4Qjw0pXQNThOrZ5s7X821YKCDLaPRqlfEEXHYFrrAq7pM53chqmQXsaeomwi
HVtzXcYxLKjbhGF1eoveLkkdsK9tEoUXlhDxO+9uZbtXedq8ajjpl23sd5aXfupO
aDewmH1mVsGcVKbVQtY1psyH7fiF54sigTIGdLAaY9tZAlAnWqJK7nKeRez0XV/I
NksNHOpJvAs/CWwgt0Pv3TdaI4CCSW+hKur6uP599JqjXxmxRjpf8m4BPdaDcbqA
CAgi/pD/xdC0M86VdW6xFJBT+PXNrvCJuKjTBR/QeCpVgNbx7NSowbRjC+ygs/3v
OsowOX1h99lSrmzJVxwb/bzMXFbEt9Oznbgr11ZlV+4zqNroeagwFYrwPLoP2SVw
XIcZhEVfyB4Tj6X2y9ypOxopmWuL4j7Ka8CcznIiopko8e8sZjt3wDxVmN75ssr+
OPM60w7n6C2Ybiy2AgHNiVq35vFdvWZTArfpI40rm6gAzfmTARiK2KSimWlAhr5s
xuKk9Sg1NwyL6TmKNmdF4glHt5AVrXTuKPHE9zIAb//cNESjDE0RCd5KDJwMX2iA
52ZJXC9A6aCQ6jtGQJpeK9xYLzvHQtAt5wggbmP5QpP0bD/wMDgGWhd6j1dhoo8W
7ZGmwqVOSVxC9g1LsU7CU8TgfZkFv+i8mSTvrFYXHnr9vC1Pqr871YSDIjc/qUlq
gALucST9e92uWxQKYA4szBNgeLCSv6v8V3DyIColZ+9SV6oAPIfPZpcFjrGQJbXg
PGzl7K3BObfACZPyFlBlx5Hb1J54EdWjmf2jQzGEwTw1u0bX4GIBDXX8wDB6KaXy
yPD4g/6QDNfi/DQf73p9Ax1TTQe/5cktpa9n7pgt3BDiq+FZlcz4a58R8f55+XEA
ofqUxH9iw53ovLJNpGsuFZQh3dDKXDAsBWWOtHBHQz9X6uxR6YZNaHf++W+esbvm
D9LmYrIe8OYvEJHOIeF0mbW7qE3YaavP6ZyE58JMsIZH2YdYWCQpmGO3AcgzUZ4c
gEt3Nl5vDMnQfYJqIeal/SKt8/p3+DC9itiLtxqgO8GfbIh4Ua8QZJPEOpHhPogB
nrbO6bn2fQyiALlcDn3z7cPAUUwexG53POzDcgqa7lf/pG1MZyCr6VOfkecXvXyy
t3fYW8AiHEzVupQzRTcUrROKl1lzDiEfL3nPny96D9wmuvWh4aKO2cHgBVFbU31C
2E3HL3ImvM/xM5pPdHu7aU0mRHXivuyHcXj1eItAprvZNKg0j9lVBAppbtBkWLcR
MwGgepoI+vPHS9UpOYzvBRirOax2Mf5NWGiOSmB3a68vzJPN0oU0wDTh+pNqlhF9
hPCX5irs+aGd6cH2+6HR9j7MvmmHb/ZWEiU45lP4xA5zQe86GSJaJ9jEYZYbWfrz
8JYU9hK7cTFUbq8rvdYUupcyG3jqcXwAz+c5KLiCDn1LD2juSvgZ8P1LsYaa+ed+
K3JZNzS6l2cZerVQ3aubVajE3T7mNu9cjC+bDkBv/zbLAyodAX8q1ebGqcnh5xC5
p/wLdvfhD4850CdSoZzu9WJVQiWpFROdO0iwdVm/56Ua36iDFXswX0q0KvefGsQY
4UnqzQTS5hf3Lu5gioRtY8NCF/veOoBhv8kCsr6aoU8MrsrnfZnn/XTA3n2DbSV3
Z5ihDGsqWHkl7sjuHOxp6orjGOUl8/hkAMRuBAe9bqXp0KJNMZNix7+da9k50ojx
fFLdyygw1t8iL8KlZrt6FWxjBazJJ36oZDRpBRnVF5bI+Pn2Bs8kINttClGyKmbA
KoG7m8MO/dNB5RjS0qOgx/8S6Vl1b13PeiokfNiRyMseDSLPwvwutb58ACym2zk2
apQdDnB6/uJW5ioFf+e6MwEix3pA0rL3nGLFbofamxWKfJr1U56F4JSfwvrceqtb
G3Wasg3Ixe+l10W38r9oZBnExBmJ5st/SIQExHTgIkOzVrh5gC3sl+ZU0DRw2mPf
W/k7joNAZhZIAjp+T8p3Rci5qBqfOWFNygCNlyKhIDX/w2pC2Sq4oZnuhDDRxmlQ
A33ueRPErvbWorii3MKe+q2JdXskIDI56/AQB1BL0dn8owvqFkdxNZRLO5dcJu5l
89CKhwKA+9tzIVMJEOSdin1jE430q0shCpsflie/5iJCSQ10Vmk5EbA4PnVxo69h
Fjsuhy12exfwchKCa+uHsUscHFaMuzKLkrTGl9h+FmDYVs9UOL7iiW0jl+cJ9Qgz
ks8K8TvtmxlxCUAqrVROExRmbWzyJj5XSt/f1Nhf/0UYox7zYHbNrIRLIGvnWpBv
C6xRPkVtt2De72VXS40PUSLHs4Lfn4ymjbpIW7HX+mgI0TgzXm1xpqtmE57y24HP
qIUaeDolCMDDF2jmFdRxfhYuUtpNqmHnH48AmsNHg8B++TbE59mN6mc4wzR5iq8R
Tk/h43g3NgiHeW8dXQeOJfmwXgKvZv6l9jUtNMncpQm7a1KSf5f0xxZ4El496Z3x
jo3wjetuHjyal9oPVuHI6qzz+liWvd0uFCTVibfAx2ns8rLghMuFrAscpCqZmAUV
LOI8wK0hTJwGrnny47290/PzNW0hT0GSkvYJeO4Jd5O9IDPETSDE3MU3Yp6JDGWU
UqxNsWw0hHYIMNL+HwYOPJHqlafQs7RfbVqScOh+BCAIwG7GgiarDNUwx1RQiSKU
rHHMm3aT3lHe4FlGqxlUka7boCeF3x5XKWSV4KWkF0zJgOuuglFqPyxEQgrBKkvH
GXIn3cz0xE+JuSa5VcqICKDYTXtVB5yENZzaWOJGDLqZ8+Gb+fywRs4OTLtE1MB6
h9A+/UDjVRwWfVzM/xzZs2WF7Ih+aS4HknziXvO4TD5bO5roFswNhDFAUILCw1uw
pl4CkpBq7kLC6hX/2HxnIjj8bfmgPRhcRnjwzKgKnF0jAQ6POUnLjmCQp180JBOS
HTnDksY3hMi1DfTCRKqngiL+2E9rT/sKgcoyPxBFtDTlSvTBYtiRgbmi+R8v54gk
MxYZGNoRrJNGh5+nQexwnabgjwQPHzaGash2iY7APFlv92EvxxC3xTsWahVr58bs
mpUtGi4bdfsmhEW7hTe4k9AIrVKxSaHWYivMbswvewEGv1CMM98eJ5lfeofaCGYb
Zbl76G1xcrTVds+n5hgyRVRLHG/hr8+l69hHLB7zVwmV8J5BU9J7DoRoo6zTWEgN
dhcSaSXz9e59BL4lyiHmm9z87wjslJJgLOzXmt0rLknb0M58871KSZ5rEYlr3mYZ
a9wZyT4H1Q2NFaLz0ozjwBghsZ1bGX06t06Gd0NlJjkWF9rhGR4f3I7Dbru3BESj
+vz8tHSBoC0xvIA/sBBCpa8bDulKnemRwKtpORXELvaEra90XvBC+htGlKUtNH8p
f4YJc/CVdWhrrdaDkHIQEbnJpMZHUjfRIqwdYhjJCYc0CA79Rmsi0XePT5oIN5Mu
/KLRAD0aFde7JAZ3jmfoiQRaWggqx2T+KSFHkSn8s1Pv3FuowsZDtXA3rADuscGR
U/8bNiKUSGv7Bwg2YXnX3lSI8KcSo7w2KbYLspYYNvKoyGeIuRUFSBH9lfws/8vC
UxnDwFG1C7pkAGOknbdl1PpgnYK/4hast/3MK80TS7+e3NJrbdg1nTvkuBTr04MR
HAGxPC3tt3QtdDiuIDWxS/s6vooW6AmhvnDYEymE5XncuqnjW4PFziI2/sBoJm+3
UQtYbO7Sle+qRsdX63Y1DWC9QIugn2SnzzYBFKo0iOKWasheLmTIHgGqgQvh8G9d
GHuwNwNpz+RfZTzjcbmXt/NPpK1Qzt3ZnqO6jCBF3//xjAmFIe9ivG8l3MaL0Lyq
ACO9ss8D5fk2rkfBKfrPio9r8yUuww8wgIq4rmr+T14XhQUg/WZO9UTgExqQC9fO
yYxwgSi2m4XfvQZNYKMnTP2idhKlgevZ+77BJ+tGDPKiPBCzTs96AFjy2c/hUQvC
OpnZ7KdCuRAYKaJTqkVfCjAxuzE3paycFlCAFpTj3bpRGGI6N3ofesiEWUdRZt4S
FthDWgOx9OGtOcLZCpyR7kEDhxBgYt9JUacsZIGPEUSAOmrYDvVhb6TN5j02nxvI
dQtXoQx7hciiFjsgcdy66I8hh7OMgwg0+2kk9Nkm8/wspRoJEQmQPJkFyqQA0/AB
O1unEy6Wfb5ziZmEl6tH6HqNJsKjVlb4gek1qF9+rN4By79yxqRqNvNygBnlmWoB
vqaRV3KOieSXOVz2BFIjv/wnkYu5hhdYpk8bhBX4Im9LMRjSNR+hJthHS/smCqPB
zA/IBxIE2LBFTONqfvzFOxVowZI8xSDHsQFKwYtUpRae283hLImjb7gpgPo7j+i8
8svNRvTCGHkjmKCOJDN0h1MI/bavFYH7HjieKrP3NQsTnVoDwMrZRspDKPHq3nhA
8asct5+ofVMtmy6OkQcowBb8jDZBnTo6AJXAbkDr+D25p8A1YJqFjvbFIKnu14Kj
2bM9HT5tbSJI+9z3TeTKRYHqr6ZHnksOA9zOIIgA9TgBeaI3tOt36vpmNu1/6DRQ
KKLgq2QUK0zZLNExWbFtTFv3ZMgOEz3ifrMgsOO1/Z8MFYCkFZCamrY5ennEJ46l
XYhB3q0lys0ftSPpDe9oyRu6OLqpYBtyZgyKgAZj8v7eUqL6CIpJfnkcnuRpkaJo
BJi+k5EuDxEobbHH3w6nu7eIE+4SLwsRG/nMIAAeoI1oI/LOWRJ0Lc1QUu9f7b3F
LDy/90ZNTkvIyVLJqaC0Db4cJwnSXMfT5tiwcTpP3xwMkq+yM6jNvT8bmS2TYAv/
+kcd3xDOH8o860K1onM00HOovpMg6nLFronmjHls7w7lU5DoMpo3DXVvMgSPPfGf
XH5ld/E15CmXA7BXmEIv5/YyLs8KKxExmFoIlGIvUOONuNEPdDQySyoCAqj4Wh1t
ziWgqFyiuG1kWqGIKRL2Xkor2tUUZKwmfTyEv2fi/MdJvpDXgzvWBRKN2GAKoDn7
tI3rtZ47RkBwMESottHdnWQSYt6s7XEj9aioqw5cjdaiprzmocB9SxEeVloaqOB1
qv2HYTJTkKVfXe9LUMWHU8NOmcpAYuNRUp2r1WwzhndBoF8UccNvJW2v4WCzqUvA
Vd0UEHsGqzfityKmvhCsKfqmPyDnD9xv1o50/8FAejD/IuQkiUVnYJ05UBmvtlPo
CQLBq3jC6KYfJG9WmAfF5fVEdc8Km84o7lhIglPaAGe9RnKaGxnfzLxtV0mzW/Rm
K06qqjIJUYsL0HErrdgYlHZ+Tb+LwCZP43hnj7IikbPe7z1e5+mK8FrVcMyUxiuW
9eVAdQSiINOcFyLumZ3A+5J05Np0/7s0xLdy8t7iQm/WrAA02+fbJX33COGNt7mv
6rVp00lE7glag5pBJwZAFpcaS0JvLY5QrkhDq+upCLetkPrL1E01ys/lcKZrUhQl
lmrXizVc07Rrl04kuqXMw/R23S+3FRriytZDy2R8IK8gesmTlrqAB7t60zYdvtP+
9Fc85r4zwdE0COF4vs2L7Jk1062aIYIEI4dyof6MzSsPYAKT+ISyaxInLV/HH/45
ooEQR9uYGtJS/3cGuFhcGhW3/VfuGh1dM4+0t6wDRqmhkpNeLQIq3ecXAKdzUql7
8onFXTlGVKbcPCEliz1fktGTuM7VcvKgwMpL6Uj2GJ5GDn593/FFt+F7c8AMhTan
+7h3znVWyIKmL8XLUEHatejdWiNudkVox40YxmDP1bjihwNFGsDKVHM3dGWEqA9+
XCS0bbrV0YZS4a08pENuf9cQDNoi9T2+Sfmgbjb66wMMZ7vg99x3M+JSJmysB+jH
vxVUlVgVtrnYKMyHsf61HhLndB6/TCf7hM2PocV7Q5+jdYmzHdM41QjKrniMAARv
ZMJiD08lJX2zkugRFL65+pq8c0k3cDJaXooNjFsBg/phR/WNIaAi0KVmNhlZZ8B3
4mDnY2AIcItw/dA+pXcGODgTTf9jGEEv9StYJOr8+ADo1VkmB6tbSE5lcDV6dc2z
WLlQBl84WgHWNR06UnoI84n6YXegJ1QlD/2OhjSJ+8lfO+uZexp03K3BBu+rKlQb
Hzd1rywem+hfxnpvOGg7/8oPlT9oxToaxaXcqJZ7LJqStAmGrMxfTBuspyQyHfBK
uFU+pInN9tWdz+PClUhmIB8ZunMg92cC+djz6AvwxWj8ykOJv5LbiAfhXKsAjqgO
WW8JPv5E2EOC4EO1AWaEo7v1iMuKAzzQE3JD5vQzvn5AZV/W0R7BV6ZqcLCvUNk3
YBdaNvZ68t0wzDekA2tkkPwVNoSp5iJPPnXzatEfBL6FHXiCAVWQ06FTv2GDFFW7
njZ/gTHsXCj18IQExxdcPAmCPjlhUh5RaUfWK/aMhjoAZayPYz4MRqJBGHqpEW0Y
uILc7UQNe0SJne1yaK/mFPQ36TeWVS8bisNZKaGaCC4pLo9/xmcZQLkg9xJX+mM9
e3mpwSX82zR9fq/pJXyGAWguJ+tmXGHJDRj0lgsLF6imre5IRt/kK2TEiF4ZXbQM
I+NALXMP+jX6arpDfVi/WXP5XIGa37wtH4cYvEJdCyImaNnvBQzJWNzrye30JLt6
zSSHtC6AvMChS3D9KLEH1e88O2CTLhsd+U/zeEsez7Z0ioSQKI4P+FLr0kqn+dov
X3bTpty+ZqnsGTEoygukbi0wBi30zAnQ05yCeoc0Z/H9gu7tGeEZcnBUdHwZmDPP
V6u8ajHO5BqVnybVGHORot75yUPmMnPNZwXRXriiAEU6Cwft4UQ85Vbb4rGp0xyC
I1Pt4CnwVNsU1YjJjTQQZ/aG+8KT4vvS+yXBdM2fTSGjtOJUISlMcMHm1+GQCmtd
FLGq90ZWH9phJccdKW+f25pD24sFlLXV/hZJCInZmtQfKO+p+KuA/y4a9BEc3ssi
6BRs2BRYtSZBEWUTzKv9qME+ZOFnSt/+t0ByX3mwXD2PHeEEMRh0uK2PuD0sZRse
DSnVuxq05iCwboykFe0SoiXRI1SmXti4wVgNRcaWuOhTVinERzWCwKRWoBhVGTB2
gDKD6hr49JBH98Mc+RO281vMyiLC3Z9Ys3IPCNoxsuFYoYekNV+PMS22mpDFLTvj
MS0mj2an9BkLD5CuWDHuNRwSeH8IEYtXFFMpQXXaKNYfMoUW9yWkqntdK1l//WaC
oIe05f93svfoQw2ywBPDRHO/RfHHQh8qky8J3jfgd7nhDhqlprRwVRJ2KPs214BV
MB4dA5JoRIMtgYAJdYwhxfOZaMgZHb4vX6dL69Mld4DjyzEwSYp9u/+AG5/OzyOK
XTHf1nUdxTlc5qNM/cu1QHHwSlidA4FYs1FeUU6pmW5eTTODFQHSVt22gPFrYOfZ
qt9U19kyvIVMpkavy3C5CyJmh0WigsYkEufVfiMvgemYgbzTNsybaCF/mw44qIQP
hAtmsihSWNfq7uKRzWdPURNQmqnZEWwA0NgJDoYfCi1CWFxrmHQs4Szrnet8yQs4
7QvavPh/De32U56+sCUiQ98VYGsDlNPjw+dKtcpupHrv7V3edwjS9P1VISsof1P9
7/9MBu1nPY30jlyWeRvIj4bnv5nomzceEL+SG0SZrGg2FVs2QmoDj9shc9KqF/GR
5rtkHFYBEwHxHazkN2Ck/+KADvRbT2UOaLwR4WKsQXU5Ej86piu8O1PXYkGbO970
9CuOUo6kZ2umuc5viePZkufJ0hz3LuTa3LzqBBBjWaQYhJOXBajkYXs+foIm4NEd
cvG5JpMN8jnb+sKETJVdo3XdN8ZJPHPcs9+4d9YEV9Y1kaxkv09DIHh8N7JSJdzs
Ncfu3ucajk+qWav2VN0ZUy52+0VTTmUvmd7DtGIC2U37U2Z1FmgjPHpAQVqCcwJ4
zWYu/aeX7TXmY7F1ITYL6TXPhzr1FaVqBL3+Dor7rWOMfo348JSGlZZp/5j8YwgA
nSRgSVGe2hMdWShebs692jnQ1QJmCnD5Uc/B9Q+rmY+aebq6yHHx5Meb1fvNCwHX
ZSYKzO82rdd+IkwTe2JSa87CCuvdI9BZnviJ46Vs0ab7GRb8EgxzHNxRBOBzl2+D
1Y6vp6Ka0/0DOLymjPL3xrlSP3YwdN1qWXOR0TBdSIt5fQxqNWOvYdEstZgNVUjb
VDaM36Ajbu+ySMFZLsPhNTuiXqXdrPqWv23t/MpsRl1DxEPOmS0r7q7QRSO83BmU
68e9OQ1Wlu2k3pZhomdXM+yZHqkyKeOqBDsjug09L4PUuX5oEgRfPLOd8oNENWyD
kSMCrrGs1nxrmwvaffQxCYTXLD1vx3ke+gdDZ/8tk0rHwqlZWYNs7KutUrloapR5
NC+mkm/56Rl/kNQ03rkmtqeOwNbKlHrv1uiP9oR/Lt/0+OVOaOvyUZqFLu0YGxfj
r1lvvn62rmfTbdv/0irHDSLlVAkjd2hbLPwrNC3+SThLPBamiH9+w1OpD+x2e1IK
vbvxVuz5sC0yYC2gZfa11xLwlIlo1FE4SwZbA8pXoDVbr7hRnrrMMK1otqiT/bGz
n2cP+l8i57DyBnl1cs51MPAkJHT34axtweeSuVxjvV/9ntCZIr/U5iD7zLR0AI8t
NYymuODdKCafDQRcKIdp5Z3/b9ae2JeLdvjP4btp5dqCkL0UKT2Wpk6pv7k5JEbg
MWXgNEaLS3JdfQzDDJ+jcoQKUQt5euUvwmzxqONaV6Yt/gU3MdjeVNv30+fAeN+1
0Gi8OAUkPDGyqKQ3mfruesAO1tGDtH8nSFl1O128a/gELYWhGujTu+RHVnVRRE+A
n39VaEnT5qcNVXj/H0kjOgNrVy3zDy1cPWqM1cYwkxA/34aYuC1BZPgvs+uE9FQ2
WRCtMYDnYwk6bod4GzDUepE9Gu+vQOb4dB0npp8zylP9ornYV+pnFepvYPbhQyzs
gYyWXUQJHo517/LAS9VkN+KmW557C5xWAutrMCpB+939ZtYo/9og9ilj7qBU8TKD
w++RzFiJz65T+myCoLOSCCyn67NoYOjkOvH6eVInMyEp5Oha9z7SIhgj+/2TSwuW
ig3vIFrR49cCha7sJY+FE1Ekat2V5Y86g0c/762HJtHEuitD7PkOUl8znEyi0kl4
ZCe4gm805UGwppL7jK29Gmh8QyIIMMR27y2ZuDoWAyIj6NoQvF+BLSRmTU3Zh6XE
5mlMmtbD9qovhGHWkvsJBaJyoBjBdYYmt2HEXC+0mIkc0SnUoE41q9dTzEdyuR7O
VJoEwANnvwEDq51gFLmAgYRn+Q7rC3vL6TwGi0pSTXAGN6iIp+/Tcg2eOu0gnhLm
I6ZpZY+pfPghhcn55lpAfGPU/oi1KdprZu+7w0/xt8e9g3qdYJNMPJMpRD26JxRv
XTiY9wGejHMVPvZjN6TBxUp2NSfb4JTJbCR0SaJmre9bN6ZHRcfwL7NaksG/6so2
X2yB3Afln8rfZHufgBfUP2lg9pAFtLqhBi9EZiQ5q/uodQNCmTcIvYoERuIEUf/5
aXxEksr2BD7f9f5QML0Wxf11yVcEaw5fujyEPEli+b7Kc0+FdDyJuhHgf4x+5sL6
c6B4QbR5Sl72DCIhK4OQAbz9CDe431zcrr5tOgfM/IIzgZMC0KQo6MDB+SmXqHCp
Pi4sFe013E/I5nvFJofBvBv7VkS0iSDVIiKumluloiFf2Sr/wj3vNZ84NPPI67Ii
CahAYJcciZghrqYhXbK7oZZRrvntE0dgi/VYym/yycJ2qsWTSh/3oA+JPqCSDd7V
IdGJyZdk4k/1M7WEitfN8zCOw0KhqmYxgH8Tuq9qkZZnsF4LN+gMziJ2Ts2xrUOM
qbsN+jus7kiIjtZKtpcUlusFac9YCmZLNB5NpxrTeUqMGCIWrwybEf93dDATBTGF
Ga2/PxaQOzZgtEw1WTWZz6bj/DswgRR41Q0S8q6xGUWdygkZ5eofcg8WOJLKP+Q3
+0I46KeqNFUEPFFl4pikM3CAYc0l21Es7pwVn5Z6d77Eji0n9DBO6dknIShb0icE
ceBPqRgN5w2VfQlHEbj8jRuuTrfQdmwJfwoHburPeX+eoUtVxvtI1cEJJN2xOYRh
8enNuZTKKW9Q0vKDxFEYCUjfikpuoH7M2l2HqdVGTsiQDxxpEuZSnwnCksb6ZSHE
oI6Gmi9DjlKSr9iG76XRRGJ/ZwezbNbydWGRBsX7DrMq8WAGpoZeSN5KHufJrf5W
StKWAWr0tj8xdCVdkB6pm+6PmrTKIiOByPUxcnr33YS8Cvov1ETBsWXZenTMC3qN
GlWlTchWHLSOL9RfeDkJG/gLdp6F0vhCI7hvaL32mtOStzeFr+YUVLil+MknR41U
dXsTy5+bTMLpOAfrtK8KJjjfKeNwIvT5z8pKfWDjGhYDVQBfDjU3OJYTaw98wj4y
Hf+T7ZgSxUj2n3+FFUh0rF+TPYc09USZUR7kF+Ii/pZ3oWe12dkjer7YBJLL81QX
ZoCKK6prDWlCZZrSiqGDFdghRHGc2yMoXH8qUiRVfck1RyPNTe4rFQpZRjo+VSnY
5483zTB3EOeSQeRLmV0ucRviFEukr7PHI/IKXFR+pjCAUkpZqebRnq1gFurYYvd1
EIsET6muqCg/iCEGEBir11hsiA2FlyRt8oi1sr99tn18FOOt2H0ei6t3QWHaflMC
3Yv4fuVtNDn29q2lvOOcmvnooOS1HtHWhGjrRkx/gZyymTo48bjiVuALxjzW25B9
k+XcWP76bpYDRa9R2JSR8048RX1h6H0mfy9Sebg1/oCl2FI7ASz+65IlNc+OMQa8
OnZ16fOT9z15hAydHYIX+1MMxD0Hep3wMvgDGn+zqnYWfl0XJG1Yf53a+PDFbZjZ
ThZ+2cKcEPd3RmxyYWoKQe7nwnZEZH38JfF2mkYNivSTTnRfXipOUr/Z/SpRsfKp
agRb9X9R+htTLEiN/XXgDV7phUAST7y9+GDnZ4eVSV6wnfrFd8VvtyKSbnV0Oyig
gm1oCw2l0np8eUSR/vjsA5vO2tEImIvmgAhOzkKidEOYciGBD2hmYVgPSCup5R9b
pgUYsIxXStRS27A6oH5NevPOeHPsRu5OAj/Ppz4vUcNicourRDgU8rsAp8B0rpKz
6oTHHidmS/L3S326U9zVTYJcAk/SzOynHqoc8kGjVo/2emsXRTYTuCA95pvpac88
xbzWyLwJrFuTEi3eeX3eruQ5hiYiAifMwV4VZ6E4ABDxH9Yj9mPgxKi2hCQvlqV8
O02RyBjX9PVgqfbLg05Iwk3SWgUGkXabOWs0lIKxQPPBO9/B1Cdk4JMH+OuLcPXR
S+GrMOUnIVSeI9gyYyXb7EiFpxTWjUnHeKKin4EHqqaWG9d9z6vvr+n9yWcoHrLw
Y/zV4aikJcDDlVryiDlavnHcGzCefoLmoG0qgf1ZjADorQ0pYzSU9rH8dOxxRTrM
M5UT/jAgvNZIkGaXYZaQy8cpaMhMwmmBIwmo9Ync1G7WYXjl5EWLjDWywkVfRZF4
ioYFjIxiPY4meEyHxD7tch/PDJvBtnlEVugJBZNjqpfAItj7GbrSMeiinyiucruL
yGwhUnuRZzUSkwQIrCCA5wjJtX7IlJuPZC5teFF1w5Pe/olHKEq8HF1X8vNn8n4P
vMdnRM7iItGe3lpz7rIRO22f6+7EaS1pz7H0MnXr39eCdDPDM9CGpcxvtsAYmTxT
H82xEIh2i8czNNkbyERICBHMRP2TXkYGTNVT/ipPqwtkhR2F/ksyymLF91V/6EiR
0CPCVsQoE1eFhW+hBP1So7t3VLcJgto9wPtEONlj3/7RhdanYS0KvncwCyRF32w8
jvqlyhTR/4+S+SRVY5GfXkxI1wkt52MGh8mTgNU3d4R7W4E0G8I2jiZpiACMGdDk
dSJJAhkk8v1xZy6KAjC08GU6zDla6wJMLMnEmU5N5GJ0Qa0c+3CHm/fBYdTUEQFv
XbFVIA5jJnYIQodKtjpb5+4c0yySrUDiGQmtpdMa0v+Cgmh88atR2cfXESiLcyKi
MoQpnN7C2RkRaTZa0aDxQKQB9IkJil5uZnJIdpyzv7OTdv0XzXF5QusR23m9TTwV
ZFwGM+YbusvVocMckud1X4AhB/fKY33uLuUdoI273fosy7YIiCS+WlzFu3l5a22U
EoKTcaNXdhwcFmeon86JVHsN10Ac0F14pcH/l8iXENx06zfbVprzgKOWMFaJfN0a
GcBn3a1DeZee8rGyy6kXji/QGJlnoxKXCCOuM28CB707zNFNg2HOgdpLKj0yZvOE
QTfvRhA9QdK0FYXnfX9Z31aGnOgtPLsC/REmOiKaSkR6H7PshKEq17e5CIYesDsh
qmes8Px/B9gJ2ParELV6L+lY/qTGeyMo4tXgfUZLnSxPFSNdiUWow8z4934IpTWQ
wfsUcOjkA/o30Q9bVBtSrRR6bDois2eOa9D9E/7CvBV0IQYdOGPegZ1dIl44nHI2
1MM8tqt/VGduuWbH+nGEiF2cNICzrXbO5H+gA531N43to2AEVkec2U2ySsEUmfiD
inpflkDa+B2GmmI8MpABwfsfVEvVmhH8oIVRODvHF8FvU7vNiTHNuMukTeFZisII
Bqwg1iw41NV2AMHWFAknqRZxvUAmJzCn+ZH3HvBPcjwyQlJopSz611iJr3t2+L9A
kimilg/v5DIyJcrszfTnLUH5yhxhffORhi1gEvRqQPo32fcf056ZHVsxf9tFPufH
+aDSYPwOtahJHvYfNUqABi1UPv2ww7JBvYTZoTm+N5qbo6wU4GPKITJr5Yqt9nqw
P0B/SI3XHCpc7SgB8HPHRjB/7JAAfzHUPAeRLArIUCf0XoBdtvaE4xZfg2x/5xfo
7rDWfagjoeNHOHltepBBndn/dtCpsXKMb08QxcNeJq8aIQ12n0QifFPGuuKvZylk
GXJTwHb7WKXrENl3jWSfnSC4vyXnVoXwUrbNHGsfpTorWe62Yt0kHg1oK9dk+xxE
7U5W2HTR3F9EagKUv6YLLJ8mDTmrzknk4kZD/ljDxG5zBZnFmK0gdCL5CXi6aPlt
cx7dxiRgH+IW9t+ONAnUatkOAEP60vKQGKlOcxaG5WkcpmFfH27xHjdi5bMT9zvP
jQweyW4eIaqyRRNrgi3ASFZTSR0PTcZWAsLE1RfV6fyPe6ZYf2RQ8zjrm4SeGdhe
E/fj6UdePj0vcaYhdAXzbVF/+UDHNniPEpu770CjwWwK4ZYiFn1GlYMEn4kGQUhD
/beGZjw/ekvuNeRnx+BiUmhukeh3Sjbtk5nx9qvDWL5QNGdve/uk54zlnI2+g+9f
oPx2MU8JCIHT4zL7VTogcgVVj12qtfOvhDtaZZgubdBLLzqaWokZC1NcbveSzQGf
BJf93EIBh9B/Noy/SNpHiRxOc6aTSs3yaTXawQtG07GwI0OninZzipeByrLjlO53
PxuTtIGACNHaRjfIqGZcCSMuA9+EBosTWkzEbzEfNy0ZpenfxSbJ7qiuMOukiDKM
jwXYnQyYSW2zoxKfoicQlWeF7EhS2BeCfHcyB57VNhz/T5s4SGcxP89ubsBGgqnE
2daFp05BTgdXclRdxuOjY2XqA6aRF2+CUT2Cl+GlUeMM6r+CmrQvS4JjD86aDaPd
7vR8s4kYHwjSCbwlWFYfQt7ZLoOH3G6iLzesHSp6lIj9BSttclVJTzjpImvxFuUP
HiE6OtVCO5bf9Fkn7XkAg+rEdPEQMe9/dEeXmaw0T+U+tZ7bBkeeCSw+lKbfxsvF
MuZbtoGZyMw2Z62u0qebqKaN3B0IhCwYN9aJyqB8iwmKaveg9nDe2i7ucWd3Bhdd
ZZ57nJW3RGfLKoIZPmzOxq53C77DXlmOn0LZFcM6RwnGAspctEFUIAlNJQgtS3XP
BQeDbIYcNd0Y7o7ujjDK3B3Ix/GwUTkIrn6bM9LvRSWO583JNfi9HAqWrrDaRPkw
qs6C0iLz184VP13Xaa0sE9dNFCJXTBfg0Zp6zNVQpOTirpqtbnt1oFgQYFzPfQan
D4qhF1Cwk7/sHCA1JqhMOwv+hV8S/hreLePi7yDQoPWyYaoYmwDrlvk7YNgFQZNa
yrv1kBa+Qc3PZ3VzLMcq+dArl/yAFDDfv1weeEYHliBe7sOvUyVtcca4W3KFD1EN
0vKgoySJQmTsW1revbFch7WydG6oT41fYJEHdSciL6IIX5eMnMq0CqIRMnXmsyNi
KapTVhDRUPL/J+G0/lOYfkfTK5WfZBqbac5Il2zBXRAnzajvu/yRj8erHMElAJAM
uKMFB/qsA26aAz+aT3CtMxD71b8De9mIOut+pPDh/M9dK2gVRK9+PNx+jAFOLikN
wgfuaMZZRcHELEtENO5guAlvNgJkgZOVa93Ds+g2SK0NEzXrpo85NaqxE1Fbqxnj
LGatDsr0l+IyTLdKBKpesqx79r9LL2z7A8SatfB6c417EnP2NKO8wk1AWIFqzFIx
niWMIRYhGmI7uGhWr53x4j12sy8u6w7xW8/mIyr+4NY6wltc0IfS+JcdbUCvQvzp
qWIhKyXL7TVcKQVHrLLTSJR3Dbs0g1ZMa3ooYmg5qdTwaC3u/7zjExQFDjOM1cD0
RwCzW14To57UsAOQbzHcg736dUTRu6SSjeBis6t0QnXttnJFptoVLVG5khyltcGV
nz9N7QkSksPR09+FZ+uPMXoVDzrBN3Wxand6ED2X/ennjcY0ZGa99lRU+BEAtNlt
OokB6AbDXSqeC6jKtQ14laFuesWxcOuEGmmA/Q8oNOvC0BHEBQIH4+o/x66tKLUE
8LKt2X2FyJmoO7Gy/g6AtBe0J5tNVSiobh6l+SQh3dS1NtlS71322NFCM58JeZ4v
/NRQ38RET906/Sb/1bxgrIPOJsUFD8NlK9m/cGXVlhYnhh8q4T3CrrDsngQ/ofYO
O+MGWCKAYqKM0bBXoGVqV054eA/BM5LKuWicv4q+e60gcmF6nkRvlFEGfYLZ/PGV
VVbPpw37/+p49RpA0o1MZdkAVdr/tX46Ukn2GvvN2eaXRL9NbRDfR2T1tvE3qUwo
PqF6J7XMzYe62Lvol/tVPKXiOCgD5y1VE1nxWjumvrYcuUYTQIXmUEQwVMV4koRt
s0wpyvTm0QPK78PENy4zGAoN6W6++k5ndXzmdPm3iUn31XLnMz2zB3kj3zeEgVgc
5IiV/vXmTm9cRme/0R9Voyj7DZC40HPDt9C4iM/i9PW7mc2RbN4qgVqPH3rXFfif
2VjTJjeVAIZfsR1wVIWkcHLeIsSQxjTeELDa6dSIy9o7Q1SOIXpgt/UukhQP02PK
PR7zERSIc1ZXw0NbbGKONHq7E+9PLBFiAZjs/1sxGFXpzPRb/EQPa6Y+kUXHQ4PX
XgbYkDzmlcZ6G76pNWPFWcWZpWgo4xR8Iqs2Q/0oh2SXHSWNEcDE3BVIRwE3ZWhc
Gr1lKuin9D1ym2vrZHN1p0s5KmMjFeXmh5hsCmkmRhYy7Ys84UtSCK8e4l9sv69Q
1HCii2QGtA09crUcWj+O8s3IuNy+pnyf019QivvXIzG4FW29K0rJAFDkk5sBrfOz
xvfpYMwdXEB8K5r5bx9l9of6hT9GMYHcS2cV++fe4000MO/K9uz3MFrFmE9IysoG
tRa7nqbT1pIgUcTnmEwW0XTABouN8Sb86Q+HmJHyUKf5CPCVvXwfDtK6lZWkiE7x
GLFxkTmfUlhhwwVThSpqoLYec0gS7g5NVR2HksJisMk0fkH6YHmV2ZfLFxE2ZU92
1COGwlReOlYk4CzUATEdxZxmELm/GVoTmELTeHh+zRewAZCBOSy76PHRcGXYwCyx
ADL6B2n0B98E+BWEsqQxN4FFsbSUEV2MmUNA6GscJDphN+d/yg8TUhAW1c4zmhIh
tI8tmR/A0tpRV9zvVtZSZ/r3qECreqv6b6KodARZH/mBR2GvjLodNnlZ1lfZBN/l
P2RHLglAfgPnEAWfoLooUlWRbMU4X0PnmXJb37m692iUa7kAtWKgVIThbXTMZAEH
8DMoHqZeOlHFCg/XTZLwDkC7cZ0U5sDeJt++Cbva+GgXeD1VY3YuZ4dRqCc47qdy
sXgLNbNN6bLp3HKJB1wr8rok6DPGpkWZxkOo1KN4++m2uIw8vsozHfdwIPhCMDro
eLL2LbxkWNm6zVglOiqO8wTinFYKNXxMjLD2f/Q7+zaXvyLhXlZ7NdKEYTjNW+TZ
TvaeKRw/0sp+rPkEMNge5uvxRAh4r3bG/8JEeD1dfeSi0z0rr5s/nc4sA8Q8anFl
fzuNz96Gu4RZmSYUEwzwQm6LWuYeGCsbKnkEPFGvo1/ueg9o/K0iPFrrIvdNx4ST
DaU5glzXBMOeTCyIoMVFB0+No8cIrCmG29scDmQ2ao8cKGfc7Cr7Ri2qTGKrc3M/
ahajNfTZeczbrTIH6kNzZ+jha7k+QiW9N8I2uFeXwwbbXEsC4wyxkZoTjJRgdTev
7ufyUPT9YFp/2lIQXSCQTt2b3ni+YnuYM8pNsRRZ6sqpxyaCyxglAdD2KTI0P1U0
zhDmq7FekEZou1KTWkOKz56dg7B1421jlGAUMLPkPA3RNPly7BJ5Q97z+PxrACpB
bydVBzdMPAydWJn+Aupcm7OoGufmZDcu7KSwl/wPF0ozoN3ddN3dS6NNBdC2ZjLh
EypaL7TPyJz4+pmBpSG+KCqtA5fpJDUAs54NKUAloCPDsplKocCKkdx7wb57FZIq
DEkTPlAehEXRkpqMs93Jw9QnnvMBqckyN+EG7/Wkd0+r+qDUX7XYN9AzI4uPZMC3
UPwp3SjpsPoUkM7taANrHNBOmmSk/uaq0xsvJBFPWby9Aq7oyijFx7RaEzZq2iTe
kotwaOizcJhQd/riW276x4YQ/opPPUwu5Mg5e1dUJvX4FjzgV99gW+DQ46XCadQp
HbL4FjgLmGTclWzP0KJ2QLTm32enVaidHbTDcEi4AdDvkaDKsfQXgp7XUrAhgxGI
QDzdKXk9gyd8aTDV/PjeJ3/i+S13VfX7MakePPJf06yES+nAAmfMSALRV08yxgR5
+icT0rm68TRAyDIvGREWHH/lnsDnf+Grq1G9HgJBCL4asXlrRnh9LGkDXU4OimzT
GcbsFMFjtGU1GdGG7JSz3ceD7G6udukrjidFl273Zmj6rO1FaLK7vskN8O4wlp17
CIjLDJ91hLJJS9NlucnxZduaY8smO2TPQRo5ZKXdcFSraNavxTbewj3knn0QVwRE
sRy3l3eTddxwgTPHIOApj1mwZU+vmVESDSsj3iuNDtf11BknHWUyYo7l+TVHF5A/
aZhh2A4b5dZKHJjkTcY6pZ0WfyJjwiAMEnxaSQecZ0sfPM4CjA4U9Iz66yzjYOGB
x5SYA3yWJcqtNPyaFVAEHUSLEXP0Tx0fHMpkzVcQrxlI+Nq5vGI6zDuMBusv+s5X
9hnrKk2jhTWRLrlX8sbDhnZTdDc7fuAKVN3hSmgVs1gS/7aQuIbQ24sfSjIAnRRs
I9tuSGWnLf2Mhlp8VsG/eQ3DK/dE2/YmQ2XVjiTSS36YDVwcsNZ0q87VJMx8xzsy
DgWwU/sP4jde6envfoifxao+G5nAwwEeV9cpH1CcVmTW4cCKVOg+S3vyIZpjpM1r
phurE+mOD/PFHeqoEZEpqARtVi3zKB8h7pFUvehTtyXwSmGpmCLVmaNCXcSY0EDH
tLMxn01Puia1tHGAsxBUTppcnnXQXG1j1FwFhMsf3gsOcayjk6va4jDpCJg/KHLj
vNs+KtpiQPq0vl6Ld6qgaL2FRvUJ2GvHb8IksKeH8J1SIPFT1I+ebQLX4dIwvq2A
2WV4AONeQE/8TvO3GiSN7fL0clXgUgqxDoSfbuUAebJnksPQyGs27V67DTZYelY2
WVaYLKdQN8gHtN8xYKd7IFUcb3z4o/JalpASi31ZaSANaL5ChiTu2ZpzeeoBGEp9
8/Uz5K3Mx8nq9z3NYjEo+e4nhk3GN8MApBYJutRMMfnTiOzAgVAmtO3wOszVyyWV
rEj9095Nb4jPeWZSqZ/45wAixwpYlPJhi3XDOhwGjGJkYX1vx01OQvOqHTotfMy8
jVI9qC54VqGATcho+50JsConVGbN4VkeuggvUMV7BarhRAuosn3UkU3rkC4gXG7A
of7ThXoDS5h8VnEMB8lARcjPnqPEB7/yJfolYOmp2g6wOs/VYMdizAoN5akXsnZn
m+ZaljwrEzUF05hRlLN5Bap/2kCyv+CYTW5WQW/FY26evQZKs2LC1TBqahgprp/+
O9Md4IItCc6Sq7RB7uOKLgeTm5oaaA9Y1EBnB1Pif8gefTJ9T0uLmXdDKGjxj3e1
tW3AgwTR80YHv+XaTDANVTE2yH/tlbPDi3BGecgWCl7Ve85HaxfHROqqI2zKb3eQ
wP4WvcBZJCptK1oPo2TAPbUMxm9P3CNE9Eva/m8TgqTr/3lbSAvTeb9rkFYWfh94
O4YYq0Ly85XA0+AMj4PU6FLUp3lItQW33XDCoUBItARj6q0Qn9JHe5G72htQ1FVb
Kb+wBr/G4v1Z3OmmhKVYk6mLsOI1u7EdomhR0GplM6gbq534s/Ug0UOIY/5A/XBa
EipnTYXxIoUaumD9yo2FrBnDQHV2lgkk/T4yovX96B98q1xYbaHxKU17qIsSyOg5
T6sCHaqO6l/RIf+J+iOqilJwgzFDOa4oEEDPtt2kjAVSsrRS8D4SNrVn59ML9RDw
h4Dad8Gd9trsl7OzG9wGVSNZLjB5ryL39kJJrcQs/0SIX1MPpUp6cnbZPZ7c7i3L
cZuwhsRgZ2ahgqtbFJJ1rAbVFeF8FeLf09NeczR/+so/W4utngVCWCV0eap6hxo7
nf32HRPv7Z6IsPOMDfKG0lJT29Xer1O251fuejPfO6d+0fl+Sx9NQDn7s52hFSqX
ljbcU3x6Je/ltT6KlEPpbgWppCRLId78c6jMziexc7Z2cck/jCzNjQr9BjSLnVSn
oupyAORcXu7SIR96Eo0yuKxUWbD3zrDOilJIbXlExK9yL0tP/Pq1vv40WgsWveHo
JUVhLlsMf9zrw/cZTrdaw1uRS7HGynwTAeAL/99OnCEB7LHo7p1GQkhvcnAdn7me
oKALvHf5xJX1whQk2mjkVdFGQs8PLiwDUBT8dZCrgihXok5f/mBJ+13tpYdfrrs5
GjQdhVAd8duxjK8x9lsxZFqiSQmfR9xfp69VnQTu1EKOBUyySx/h0zFmk/iT6hsl
bp/4xxwSne2oduyiInIgHu8iu+72PI7KnjbGJ1pT8Wrb2Tov10QOpy6LGkNz2HpU
N9u5yemaTY7K/XivKMvGXnoRq9DnunozRYNsm0oCWkrfRyLk2LQb+GjiLaM9IZpo
qa9cklwbVkHmgEyowNtQgX7chXN83kLBTwYeZt13L6op/pJenLFNI74kc57qx+i9
tDOgHMhzSkIQelexWuAQWpeC9FbMW9C0mfnrpSXVjnhcOo0PAjJ2niQYlL1InbX3
H8h7Jagbe5WhIiQxnkDiEmmNxLl2JTZqPQR9YKgTdg/MsNekwfjA9++T1voY/GgM
z1TWQGMKwTdgy65uCnyQi56I8TLakUy6x2qrvUKCNh0PK6/uvfYMEgdX+MK3K3Zd
2YQ4bx9k3gPo7GOL3kQDTtaPcY0mN+poTHSHsHyCafH8ROwilqchZxIfpzuPOVyx
JuP2QYZcElJn3zRfz6CE6jXdPQ3S5oENocagiItrQmv2RE1Tx6YkUkVdCiliiMlT
x8VE+FN1JkyHCYpfXldRJ2FVSTxw9tqhesgkwtzEXeEV6Pth9pm7pKKow2nf0fEr
MzU5s2M/KrgCOZcDs01yOw6qIsm/J87XD1zYYIcGpKp5R1eYuxO1PFYleIGOJMID
ioHVJOGoFKgMd/UFqrJ24Bxn+h9SFeLAIOB2UZLGDr9rv85JWt1OGDNa8K4a5aqp
iwDe/oJzMz6hpeGNmLJY/bg32R32Ku092TEusF38uFvsmhnzIkCueII8AISIF74k
Iy8IdlZg7ERpZyihKg/8RtMW+1rbG61E6M+NQaIqFxf+E8v9owRfFCt4GpRdVtGw
wlRrrz+lOFqKcgkKrp1rJ6HjHXL2hQHxcTqbzuGGI59YvnhaxW8PErKcCcaJYFsq
bVdgpw7XGtH25X15ogMkIjJwD8DQbCF3FHsURCI0vSB/XmgXzUpM3bWYR+21jjgM
qBMtfhZyzPwZfGNBV042/1a3NFSHqTilBooOpAFGojSwrrtVvr0D/k1leb19y/rR
t49gl3+gYeN6RXS9p/8B1fj0rvplOw/WdynrIvMZo07LHL6zg/xmaqXKQ3PeWYA6
iCIYrQCt7sZBQAmyX4Hid81krroj+4kOA096RtyeyLUlFFG2mk3c5muK2rVzAWJ8
dH7ZvbWXZpOU/prxeyFb8IetShi5IP4B7oYQUvqVwRz4Ic0E87HzHFAVYBncxUf/
PZDlsb5RakWK4/ZUD64VFAyUje9k83bGJM+CakezUKKALLSTbB/WkbxD15W5eTYI
5WHPWRSDd+p89hsmpS9tCUTizhvjZg+XYcLzTyqVki8s3NRqpMnBQhjCqfWEwfQf
JPfGTp+j7Vvk5TMfXT0SN0z7TNLGtVRxvfQ2xXd3AfgpSILJX5wI4SdA0GyFvcuc
lt80xAh87uqC69e6Ds2zReK52szsTiScuYfvE4lV8W1rnhAFM2Jq38EjAObwlh7p
fFBRysdA5hI7YpH59Pwwad+V84NzsxjnX7Tog+bUEUYl7usFFEvnXayv49On5UuW
e7QzlPV6Fd7Dm0WpYBCQl/Ilzw17372HR1O6Q3ux8glchAu788mMUpaLucSJe5IU
N/9wTzC0VczmvszXX2u6VSq7N8Vz/1wRl/MQ6+DCQ55sO3xs9icpR2C6/vtpgyK3
sGrLVL4h3SoKoi9k3a87ERvSBrk1a+e6NPbPcYyUH16IOv1bp0jegx+XClftuM3r
yqOVgAR8IuNpLcHcZjNLEBv2Wg+Of2vT23pX8yT+JFKeyHqaeDxTcoK8fsvDCkTv
gIMBWfJPX2/v8tJ1Ph9ZZ0cPXdzdhjvLiHrj4a0Yb8OA+zJ8OcqUis1Fs0lcWghF
OCzC4fON/XifKCxQo1cC1Ec1U1nPaSDFJpAbQUfZhOvByenzK9w1p4JpqqEcTkKX
Mnn6oOkeg4aWWKmCzmIj5GTJq+VjYzrq+j7Y/I8wYNu3xNd5iDfGMcIcplJn/5p/
mZm57r5fh1u4Dfm20B9EouPIXmxtJZCC0cyojDdfeKGqogp74UCDMw5X/olCYQls
lkkUL3RFGuT981S74GcgKXprpCoYGhFvMNCmsreYqIQ8MsHc2xojaQFeLxQ9jVOj
zC2Cx2nZjOiF4gSnB8Fj/Xwuznwdi6k37+tpZkHRwIghVV7GCNUOcQ6l7JaxlhcT
PAHDQGDGbVI4j02iva7eBqh9/ke8ZDaFKAqY8xUJsF4LUHG1uTErovZfJRo9VZbX
U2YllpjeFGuJ8+PDHM8ExN82fd9ELzm4/yT4PiIwqTPFvcLl/HR3kWXmlQ9Cb14T
bCrNSp+1VcD0NTpF0Q5S6KBgDjZbGGY5S5ajR9DNP3Rb/d/ax3Kmm2T1mRQi//9j
k32vPMKetC1VRFHExJqlb5C78f68pcgs8o3JdiUAaICjrZENPICDWq2K558uCF7H
lXeCBUGYnkg2McMx5bg0DnaZnES7TGus6K9viHTHdZuBN2hwfBHP0QdoFxO9pDNi
VQdOBStJBUbPWFdDQg6tmwFoNxFmPuhp8wfdZ1v9WRq6tL6Rdlr1MCxFZQCg8C0O
emSWEr9J9rvOgzHV1BHoGjAnR9GTIU1MfF0c32GYi7xhwq627Vpl0K4yKPz22Qkv
Is/9HKE7FTNtULsvMhzB2tjs10OsMEDHzYMz9sxC0y0yJ28GNziFnBohghTRHz/l
j6jUQ+x9CfB9MKUJLY/aB9+wdAEJGTVYf1044d+ipVodSJxwyEgbODmnbEcvB1/i
L4a79nrimc0yYTxVLRUtAjYQI2Pex2KX5IczZgnWIEC3nQjrUhVUhYAeD0iZvkrO
cqHI2UAAIkTUkUfm6M9O8mjwuEuMxmGqP4UcdH7FB9XBZ38EucukV/i2M/be1d+u
+0oEjr4P7DL0Kj8pUv0IsLUX1buxhTxlZtJ0dd8Bhwxa0r2CE/CSAhqzscnAGgWq
rTYOvAhcrWqKBvbkcQm1Y8APVKfsGwMA2y98No7F2YxmGfrbF0qPLM0vYDQJmgr1
UACIy+I0tFRuW3hSJYUIM8++X1Ye8YhjHJHD78RiHKpe1vEUNW6E0tsC3dkV4KTA
Ayb+rpQs1Gf1/ohhgchv2frbwBnyuVD6T+6PPF71fASzjZibjBdIoXW5o68sIP36
2rM35S5gBK8kA8z+JBig1I7gZ9jtG8H9DC6dpG2VTi3tAlWg9NJUHssjsmg6zOSm
LL21LH6gzBIqckmE/zYCLZ/MvxltE2HL1XZPsI+u01OPZNpgciKsQq251PsV+K0+
FhgNfQEsHfyQF+43gHKhOtpU9gclDxVjiovEWcXOTcJKK7BXMUyUup7lLVBiU1i5
kTb/YwHhRra3uoQHfYExEjuf8ICeHhHKgdf70ZrmAU4MPeLG/jqVHCUVJ9W9+ZNQ
GHO/Er6YWggDqnrxmOukF8sTxZwdo4fN7sN+DlfwjM1+ZxZTDZAlk8833MheXtgj
0otDm48N1/G/8Kz4kAXJXENemDC5ATbTK776IELN/1nhnTNmT7T3g8H1JX4gpxXq
kmBp+8mDqWuwxLJ3VYSLFjnEdi/GRl8g+isNstvTYiUOS1pe+tvQLt9O/3yTVVBo
4Lar1hjXBIveKA7JdOabReALbmfq3Et3t1HIfMOBkd7lcDs0y+aaHKxXgSto2NXT
UVGdaA5+Nvow2U5kivIy/nK0a+Zd+QXpCGYBasRXejR+EFQbMfaUky/8ZZd/tqKg
knkXkBTNw8LI2FUnbRZjQJltv0Vhxr0ljb4ixhIFB+Sdpfdgxl5+jRKgq9c36c5h
RXhoDXykTW8J5A5UiCXOvP7TpwgNOsBAiHuer30p/ocGifuDCLflQoCB6fXIAMBE
qNS1X7E57HfksBXrbC2FoKUrVS4f0FzFaeSuhtnySiAgpGsXKtWym4akPhmbEInY
zSDhbEohvPVK6V0Ar5RpRLNREdt1Yj/YyGfjvwjtuB8svvmlZTTQUfYH+nOL1KdN
s4iurr3eUFREEKPASEaAir9q3UeScHeRqVH3RK1qDVkvyvCy2NG+R5Ppi+DI1m6E
t7zB2n1Juk/+XB9YdAsGgkG/6hl5PbtN5FWO2H78JR+SvAa5tG95iJ8NOEdbhG+i
huBTq5EmOlj+bWrQeqd3A44+O1SvZIbNJg1mj5nomYpym9htQJ6sP6tTKrWlO1gI
X9GBRvBbPEFAMYAq0SgRmptGtzsIbdPtUTer3gCzWECnM7ubEZ7tjLHKpoxCrEDi
jA4DnNe9N0LEybJf2+r5YKa5Wc2rrt6b9oCTX/wgGkpSgDs1o9oC3ewMun7LHt0k
0353SoCNpYZCll8iqEm9agnGmS1JXmQ2j0++h+7YZU58E7ZHbmL/7W8vJv6WF2K4
ai9c0rmVzuZXJ52R8kv85Igj2MWog6krCFEeFSku9eqmygiIm0DFIIwKq0M0QR5v
DjL9EHp6kNL38ivMsWucJZ4/j9M8qrZdyiiD+TpOa4dLyWNwrmUj288ecQYhOTyD
bOkEirdqAEQRIbxsITkVhdzm2o2GyvjvryiitycEUpeqfT83GDFP3h1JbFqUcsVn
3ggEyCndox1+11ZyinB2qYkSgwHsNgs+Z4MY8yGy2M/aZuwP1T618CWF8bsz7uIb
P3lR3ksfvwNolj9VQezsZbCsQX8hSVWNqFCNi7btbuYneg74xTvOtCu8RMVlDm7Y
LdwZsghAuHXRiQVkGiciSSA6icvOlVZDYfMIUHXQhsPhqByGVuiBPQ5//igVDfqF
q9548boFExoCX8Em8DdqdEzhJ8ilBpfES2rwyPL2HhYZVFzUf5cQJwNsw5RvOSls
NWp2HpNW63uAqhTUVbjqfDSgKqPb7avc8L9F9roFZdrVkXybT9HnpVwTtyCbhUpX
BNOgr8D/1Igrv9OrkjANkXS6AZRD1sUTgu0dfudTKh9LcQnXEimA0X57fw5zXROr
/lUS9shXYgPBA9agXDcS6THRvXdMFakGIvGysjoNe8kZD5AQ2mVZZT61Zyxx8GCr
dRGk8VAeOD6eZvFBulRc+YU6L/ARMFIDKfjQVmZuPwjeVDDFFiYVRHjRI7ZTQhaJ
0DY4Bn/DfjkylHY7N0AP1upjiQAZOISHR/8YTVWNe4gruITwEd5EVJdy3HBGYbC/
gU5/0Xb3HXIF1pWWlsVSaVIlqdwW+7t1IQPAYEIYDmiqAzG7ZVSAU8JBOEGWU7mZ
VO0wkToZ10gQGTVQHJ+IyXt+Civ3+6V7/PhVG6Wk03SHPuJbOX2BGecgtgUw0KN5
4N0pQNDr8OVrFFKbh6RVU0aInMfia5MfuhBFQrTM+ya9+fYouZvM+TdTwMGpeUsA
Qv0BmrRQa94UGCw8eqvjKuk6SPI0IIyqY6ISe1pSfpdXUsMj6jaFt5ClTxshPpRb
eylEPSR8MEvj5PJ+EBS6GmaDtqe9Q9CDMB3Lg0+s0y9hOsQk1JuG4weo6Es2IUp2
f5euC7FsxCgHVT4OJqSw//AoWyxBqpoESVtur1rLHWi24Tuc9eSDuD+60amisCli
TTz/AT8VO++5rzb3xsgZiVjMDs6J8x8shUIjJ35by8QNuIMvlq/oj1+NqG+czb2b
FzvXYQ2lRzyIqS71cu9Xo+obiMccXTBZFNJB0JpfI+dcxGxjT3lt3pT1u8ULMIEn
u0iTAkN4pqWZWLUdP4NWyHCrP7sdEeEoQ8MHu+FYnSpsrJ+sBXIwwyLBPwbw0B2r
yn4w7a/5Mgpl1OQU+4MJE6GTzH0IR6p6yI5OmzZ+ug8CI7gnugqm9Oc9pZJ8Vsgy
Uf+GxvfXq6Nc+41495TxNQaHl9qJmb7kSWCqVzu0qgbZjOFyw8TMYZjMS4vfycl8
jMY6ctijsAp42x++kMqhe++0QQm45D/UQ47YUNKnNZ84/UhvXAVCdhH8blcT9UxM
p0wfYnKv/8kP5tS9ZMdS6ndNrJtmayR2DjsF/+CUXKffA+UeoKXu7Cgma7ni1hy5
uBUoI5BUEAsXqY4vrjdqJqtPIWaZgNdIfCLT0drLShYBeFQga3z1aEjibeEUYNZS
yYhkF0KeK4y2PCrgEBFq37pgWB5XoA/2PLMxdKHO0uLvGUOFgo/WceWu5ADnuxlM
Y85fmcB3omtmtNqjJvcw7cPwQw6Di37ss0phA8bcWNiCY27GkDTBG2n7N2Lsrl2K
VYt333Lw9fuiFu4v4oTbRJviG8LGgAxdWG+LHsNmhHd2AQx3Q4+/ANF5+TZA4UVM
mQ4ssB6I07HmXpdr6R8AJZquP0fvNcKrnzosKr7kPvFFSLpC1KstxBsL7Viyawe5
LAL3mhSWy+Y0A15DT3J+J9Zy5Uk1MPGTBO5ksUlIRjHnUH54DvjiugflTX5wy+10
SXGm2MrkCKCa9tbYjrgROChdHNPRyL52ChARbREf008bFWA2zLLES44SfeTkKVFx
a3TS6z4UjeqczIgh5HU+rX4Xjwbk4dmS9niS8Pk056if57TkFw1dminDbc7lh3PB
yuNcRjSm8AHRSxO9TQiVTUpFy6dmdeUT5RjP2c3IQvgyQ038MmKFA9P4MLu6FFtc
bX4V5rPDBpK2JxgQvcFqGEIncQsAPJOgxEPcFRnlZCgYuA/lgIYVkdTCuVTt3hRP
tiLQUEE+JwSlfbZj5fGOUWv/W10lHzPomNTY+xj1blG3cwGmzsNyWbJ25kzNBjya
5qB6CoMXOetuBtX/+BPcIEX7H0PLRpHx0G6uXFFI6aEWyorJT6vi86+NSer3fnaf
CUSVjyvI73V0XePxmonFtu2YKjtouHhqOa9bptYhw5S0NJGCI83Zr815JUOOBa55
bv1PrEu+DkQEeZazUUFPDtbTBkesbBEWWYWwTFO+AxrVBBXjwrGyo2wnvX9mJkyS
wTMsq2VyCkkVIL9ZQLdZvZVPLj7P+BvPpWsHd8zcyi/48ShmuY4tpcpjSYpRaGQK
K+z/oSVRy2+0+WLJQjE/hw73zGDXkPRejHAqWLlk6pebiSmgZ7+MAbCDiX7d61O0
+4HK4egfnSC2z1DsHXBPwsXUYPbYDLuJGRYEdQCf39COdR5udanURoxQsumxCFDH
tEHaU0waNlxyAWmH+qEAhYZ4z0ikgDZ0Pv3fcS5wFz+jeVvYn76KRgLlEbhictMF
+5p+IV6GHHVkhNRlr/YBj+3xabI6VHgfEdG9cMlnRsos7R1vYcQWtW5TveHgB1O3
WuOX0ZHfnDCZAHGRN1IDHlywnvenmMwrDrjmuyFxpuRocG2ssWSDHZZIM26nMwBk
dif0Paw+5ok2sIFwjxnrKhZBUd30KjjhYoEiI42gHory/QyRN7e2eMzvAy4zlBXH
BfNR/GZKRucOYWicaeihOLB4CVe9v5zBdR9zhMXWrJD4jkY5ytm9w0pYJeSwMT+X
Hn2pNQpl1oh77APPBqziOi2+59bFEh6FvlbrgFUFj/LOt1OOUssMfRQUNyrejcXb
XVKThHWmCeSP93Uw7pIJrWEmd8WIRU9DA4QXu2G1rKnNRKx6PFtbQbW7zMj89V7C
5dDZcMjaGJWqiRW+g2xOLnp5CLlWXAKmg/qgMFa35P6w3uK8LMNzYkc3iNkWlaP3
PnRuHMP6WjBayTlM8yVJ6/+79YkPVLy87ALln5WTPc31p0HmoTy3lt5CEx35Nsfc
vg1nzOGH9+A8vh8YCU0jd0z6hiTG4EipCU3qnSfyV5SjzhcGIIdVQ8yTDUfuFIak
bFMkdDSgMdoaBDKTuVYGRFRXDb1KckV5MVFuIS3hhXvltp0fmzJANRxzdUU0kXzz
zPhHYhcE1nm+pPrHsqjjLxi0XO/qMGOYfGvG9w1/X9s6+DSRVE6w59+xcUzH2L6r
8YOn2oasmbxtvBgjMIpH/KpYGikOcDRs2Yy7/3sBZ1AQK4AM6ybCFG0qN+D58Kmm
ZUNdJhuGVbBkW+6/NnK5zFHO/+FS2CAfPzWbSIo1Pu5lrPNKY3kd5WjVbXTM0Nnq
ZUaMo0CUf2K0+7fXAzuQ2I4hLP53TsXdIJLMhuI3rLo6+5XDiJEd0lpQsGa88c3I
95HX03KIMXQrP3RxbTjAWM5EOX9kHB73yRfn7hsvFUmHbC2CYYWLknjWP2vM/Gad
w6VoFZayq8Oho3APdcNnqgVvLarY+zTvPL1pmaL+GJRaBghUXbyHkiw/dg6tm3uk
XGc5uD3dyLpaLQKm7v+RE44D4UZB69RxucReRBIYBcMvWhYZCvaTjuXd32sSLRoK
L/x8OHHAce1ITJiXXDf3oSbo7ytnsD3Aw6OJH3WhMg3munKxS+1bNhuGmY4gytU0
y3PtRSkdiOZblQMa2Ol10/RudJPY7PgqIlV1IjMYezmIHrKWSkqssa1iXRu4vJJZ
WvP03q/TKOAk/89hURqqXswB5FhH/YC0iitKj5nG62YrMIYJuFxBf5hnQt/wR3/X
Ujd37BSH1WFbJWWpEZu3lIoIooytLX/51sJstH/hCuIRdHYtxj4OJwyPCO6itFVW
v28TF7yvLxQBj+6BxiveJyJ0tXG2ysakiFTFa3klQbD9MbVwpFUUsA/QWIl7FD7b
okXokZHC2y3DIMuZmAwWESOvEDo89+PuLnIuTh4tMW9VoDn6svkT/vpCnuHUAvc8
yal/wBT1n68y/H964i0dBKYC+F6Yvzn2w5ToPTod1O7UeJ0/k8VbBE/l3SUBV3Oj
z7fsUUctUv2I5pxWW44m1i1c4cmcjONZDYWtxZKLuR7Iu2JnagJp8brbDVfzvQnG
aT46TH9t5mcnGaa92InMSI+T3yTvNaF9qO6KfSqIF5pZ9lantCGEe6HwqMF2Je2H
D5aniW4nE/pae4IHDX5veBmHiqX3UaP4YtM7aG6qCJTWcbFHutrYzu3fBuiBrcPF
lk85qPp24W4H6iqa+WusEIw5v8uVXBkfkFQGqVWmCcMGk7hMjwZF5+mqPpHqy11M
N4SWPr2DJfJp/sxXLXdqPq1iEH9eXF2RSzZRAwAAKxLCK+MIc+4UbcyinBSLG9Uc
rVtZSuLj0ib57mWBkSlerX+VgGLJksrYjHpecyLjf+fyKmeAUGmtYz9+v87D5BOj
NXUlsouGw4xarhcuofIFBAxqTISZfXrdC4dXt0CyK0VgPGNJ1bugKewAD23VG0hv
GC8UYcG8ii7X8qK7A5lMK6veTSVhEo+NQDXTzVELgcWKH4j/oMg0+B7czFXuXSKS
OelkkPZ7bhI0gvIxnx0xpNnJnfqZmKZzM4vxHo5cUZkx/r2iNgHKNUW36RFmYzgE
vqsvSAn6IMhW35mgpC4uXlsqRWTrUygKoVl+k+Y1U/etuevhCwWt/gXXCcslZil1
Np/WieQs0muClsPJcbWeQpl8QOTUGt9KSo1hRJibfWVAtrm0YvPBto5Nzw/WF3ux
JMytKrUn5r9A7DxpZY5rAtBBRvqcZa24zEoX6INo2b107JYhsvzzxmMarBiVJEBB
He+zT1OIE9wBH+44TepLBCy+J8lKMeiMYFL1p8CYybmKYZoyqPMX5n4bLxs3ccr1
dj+bQW4S5cB8lCx765IDvCseBKRkLeTuYA5dx33QgYGDGS7Wr5ph+tc7U0psEL9E
qaVH1QWcrZpBAxognA9uyVPEDPUo/VctNoviJQlX/uYCD2g9ON5Apcwc7kiGcTe3
5Kix4if3BCCmQcH/BaYy14PT2Aew36wJbNolgaSE273x52F9fR4f7yrQLFstYIsU
erqiXWGPbByl9yULMdKJiXmrZsAOwUI0wdG5LRwxwAOT5twR0BCYreu5d91hW9nA
wjNxTfn5DEdAjqIn5sT8w0yr3ohoYKEJ2i4fe59INrhaQL20qx5Ehcu1Ao+NZRCy
njgnRUU6d0lFliPNj5PMY11A6HHOTZI3jvodrwEeCUm4EcJSo+INXbEme5wOipUG
HmjKdWpjk5cl4aQ8TpgOQzlBkIOVGL15s4+ZCAUw5Q1gvSePSokyteub1bdh/ENa
yfRwXrZvxYnAHv9tTHZOdKUOf9xcxviy1r8fprLkkA1G6MZk80q11zu9OtlhvbHL
LNUm/guvFe57/4kQwCp+aRsb31PGOna7hGmVlkPwDXOmFdxhLcYhTG6Yp7F83GqR
hY8o6Qu26GzqeMWqJJusaTbNsi2Bw1l32kE8cLi3eRzlvPCPVc61CPcx5dcRHaxQ
kNQ2q8Rdc76DHi/+Rk9L0P36pPl9+azyKgP9BlRo0I0GagvQ1TCDZEmn+83XBoUP
v/CXZ6O4GQ45WVTmUHIX0tnJ21PSZ+SkugOlfiDug6I22oHmPMOQgq65HO7i5iiM
Gxel6xZ3qJyb17r3okYH9cVbebeSVZNggThe1pDMi3RbvLAjoDkpwWxVijMKOrF5
gFHjSG+ZIQa+IWRxLCDUxjOSks5jxEk7R+XJEkPiD6h/uJy135mzCP2YsDTwT1o4
cxj9kUR/bsSe6aj9ewEYKhWsyUnmJGnt1BD5jwsU3c84tz+Yq9M9YgEUXP42KKf8
4wLX1dVUkDQnLA51XL62Qe1QdNJ3tXMaODEuaVD/bZpsntx7f/QDPGfULVVlrgnb
eg0rPf3HLHb2T/qy4yT7+HVFGdR9em9fDbqZl64M1heRd29XYrM4m5xVhqUP5k4g
nfQu8FIDxFtAiZYq4rzgcs6b3X4Ll456fXlkWXX2XxtyuG20d1kayX2PtdUeUI/K
XuCD7aFp8Gr3EA/7WTQSuiWuTAVB52XlWM0FM5/G6CWxRvqSgV+fmavAxPowhBNR
V5y2CMESKY0AjeNhyXitF1fiazxRihcOnUJj+b6CkqpcSGAr6q6BlwtGx//0eiCY
ALr0IPOBANGynbuPoIaDCHf1IOqryhIwTU+Dauh1IPSGw8xCdk5U8OQDlqFxoSIn
7GtP647iP1WEZahMTyb5Dvnf6Mgxtp16JajZx3xIJlBvlR8Ptw1ac5gWy25SovG4
7UpIvK1KKD9x/33TIG5QLa2sgbUOy55kuKOB787zPJdcRRtaOoMFZxQ0dcIaPson
ZhpdUDJbmzgoYv3eQzLmFNDH1XKvu6U6+F//bKNU4d3vzifrNBcjES+V+681aiAC
mGcW2PNQk6JgKPcZsCXfw0YDyS9d9S7zttH2oRDe8XoiTIYCn+37SDr+kc+WZYpO
f2jwnwMwaqW2xHU5O4O0+yLs7LXTUp8D9Yb/tOlQRAkBx2vcQneJNZwiQ5xPDyy7
BHJ+0798yt59QMuByt4Mt4XmkaErvQiHueoDQt9RpckhFwGyxqBc/OFNNa7kZ8ZU
nuEXmPBUqKIKKWF8mn9lQbUe5h+g7Fm1KS14jIrAnJq4benlT5Rc9JDwZoF0gH9i
Dcy++MM5PA1yj2W1Dn6SSo8R3b7oW2gg2wmYMhBBPq0zu3ZAVZLl15HSyOy3VkXT
yP/jYUWny5Yk+78VAjphBiXf9B/XDrHL0q0VlURm5I6wCHDcraGuN3JETwatp+W6
8L/YZ/7y1lUWBxaQZRcVSICZmS8JCozED+0rHf2X08FyPsBzVrO4gDJlHks1rDkF
x509upI/ilOjKILxgJMyNsnEg6NIQYPjJwNR2yRLplzO5q1GJH4mU6HqulCLJnrn
QlC1Rke/+eUTh7UcKLNGqHeHACeaqEnv0Tvi6jjnbz/kN7dG3q5qNO3EkBTg9BgV
N/84ZPaTmHJZ+4Z2jPWNpgJQeJ0DW4R60t16sQqpJ+YSh4UVauT3oEedzBVYrMdW
1g9GQmW+XgAU39hBYisvE/llrEwQsJl1DJOUIACO6TDGI2maXbBvsjexDxioMuOl
DbV4vHb2s1+QkFGfG0ZJDmo8sQ0dbVfICZQZedhcjT8Clf+7nSiJOL5x8cu2mOWp
9FN0B4zHCulHfl0dwVy4q3H3wIbKnRg6vn6W+uOSsVu7xXHKppfvCW8qnk5k7dhI
GqTY95xzHr8//jWSLvctAbr17lN1TxJEVaP/4AiPo7FcoK2I88TvdLUvAW6o/R1r
yOcZFYg7CirE65MGneJPAvDggvPZeUJJ15W9VccjuY79AU1dQ7VdpNJjGLnYag8M
Jp0BP40SKCxvbFqJRbYJRHjTMgKHGwKalJgjDNqB0K1CSzbFNm9XXigWbAMSoQAr
t2UBUdGKOq2rrNsIuUuDF8YtImm85rxkD1xQaZA/Cdj+IaoBtvzeKMK9jH4nTz1y
VjV2LjPHs33wRcA8PE+j/ZS7RCRVeDhkzra2gHQhFV/lSulP5HjCw8L7rAlg01OE
z60vyA87KDJvXOo40KXGSNbA+S34TOD0qD5AzsJIbsa1O4GykkHqSBtQ8MzmZypS
9oX5DEshSjXMI3SRyh2+uifXBOchmA74rwKFXPyaDKtxSSQ4uUBn7K20EZMMdF2a
DPi/94iUb7+b+W0ZaycoBY9VL2oAy5dZ2ii5stAEJUg6mhCYKi6mEXKhFIMlKKa6
E+TED9YgMzoZUaIPnjdMkVgg9vTc/Wq9p/mooqgg6lVVwzKcT4awj0qYHItsDgx8
uiXmFYwNjtlZwwo0JVYfaxKnOKYLpc/EUZDc5Yajtc8/H3W5H5UWE5hGS0AVvF1w
u44wdvN2sSZrBML+1Egytl+vTozLxNGKBA/XxNhNZJLor1Bi1jLeyEN/D8mlYut7
Z2s99ZPjAy11DymjBqr7ajaDJUP92n240oByA6u5vS9jLFOYt/vJ+hKFrt65h3T0
EFbP43FW43+FLJzvBuudhFZ91D1q2yoEibW1cWbDNMYzhwyyUF/IQ4m+UeMjiDE2
jfaqchXZ0yBtg9g52n95Wj0w7aIjZfZBrP6sNXBrTKvcEafcXS2oNxTHxePZ8JQy
ySWkzlJKbAsfTisBmlw85K6TsYYk6dLLNod/kHAWTfAwpymHjKwAC0zSgV9/LAuR
HxHTt97QmzK5Pr9EFoahJFyXPP1jSfGr5BXvuk6X33L7rO7KXvcCC0lCbw21X37k
bNjFY7lkFHKLlHX2kEmeM1hGXM8afJKHz/u1CVtDriVEMBhbBsOnoMdmGA/XYgMU
GU0JvNHlMMdObNUhSI8A9w1hmvXIyqtQaIHfbxWgezWag43PcdV1kF3BC+xAG2eS
9Uke+TtAubV82B8JHBBUURPnyFoUyPcnBq8qGTunKWD7K9FRQjADeK/6bdqycOG1
UXa4xNCvk0+nq3oYsMn2IwDjALwX5m77vqDiCloPS3dKCC8HuBIjAm1Hibd4o+xn
kTAgAcYh97SusZJVlGSB5R1OaNBuMyWmFYAhfqto4t9WQE+VOg5+qwX8ds9wjNYk
56hOLckO9oV8MFi4Ra5rRNY0qAd5asaTCXlto7V9k+VTCaBnyCJUInzgM9uYwMEn
NHXdTtepdPN7l2AYMJOF99hA5/j9M2NnZvq6qPMoSMIWbK3J5sgRbG+et11UMkRr
flYt8Kml5qoijpT2MSZ6koKquypS872OnJUy5jFcRjb0IMbvNflLsf9Cdj/iryO1
gxqnm+B1NAEZEt9RLdfagtLh83z3kcv9rPLbx+/QZqvHpsQRApxpBRFQl7lywFTP
tcwmGTLsa/6HEWvljalzi2PAF5SB/OFuWR/N/nA3Q9WLt0PCl1ckdBx9YB+hJdpq
m1gkvkGaIR/oqdI7oYJ1pWZ/Q5pjmeNVRjs2KF6BzGonf5TvkOuakWIXpIp1vwzJ
q2Ai6VR7AYWlLtZv3l6Unk2/awIAdNIs6VcgDhPBlcQdrqDmkoenP7ZwrjS+qm1e
v6rEwMvvSMutAeUxhTvcXgxUqkHTGvDcF1Rr75CRnNL3EJZYAUGf84dV5BkqGvmS
UH8m0SwjgdkJpf/nsoqk+FWWaH9p9cpTnVBrP9uCFmagriOlJ9YUCSX4gVez477P
ORRoYPnb2NCdSQ6HLhpT7POswpK/xwC5px2WzJmbHW5TqRIRtFwNrBeHpDtIIpud
fQBOvxyOy2z9o0RrMDNyfXM+P4xP6EqCEi2qGCptEpTOQWDA0t7V75LU0k/FDebB
Fblnj2zQ+9dBDo2o+2VeFTI66KNHL5iSf5BiE2jR7A/nhqKjli5TCTdIo4Jcn+yD
FjHQSYtBlBiS+ufcZNK9nJIboswPlXow884aloJhtL4TI+H/ZkWw4wCr81VWLBK5
oRN2m3cgwkif8D20IZJ25HRrOWPyMEzdThK+wFBMLrUk+pZWHard3XO0afAYSyxb
ff+kL8ULauyOnHmZxIH5dHX2Md5QTvn5nTIsmUStHTbeieR6fWaClj/0owczaPkA
m2vuN+KP1GbyyvA6z2z8bGbJz7IlFYUexqVv3yV0XjRd0XGGfteG9nep0xzU8/Px
oS20laanKcf1/iPR7zTDSSDw7z4Dc4EHmdNaj0VstWUkearoR+SUmvpgqJAck0Zq
yBI6bsd0sUmM/flkDYl++ulXFIvQFgSOrwQGdFUzuPgYH/3wletOp9pTO9wAqIDs
GBaJ7cZMqaBGW3PNrYkGNw+YcuQizMdDGjerXHMtxGcuItxxNlpAlFQPm4utNvC3
j/UlBK9QTjhEx/22+E4Xunf/h904OGbYLkkzhsOUu/eLwJms/xhAlbOC5o5FodeR
dJtK2OzI3xIDFbok6jrPTj66M+uwjmfDtcG5GDzGyKYjqLcTFjKyIh/VMQXsb89G
Ifn52rf9T4rtEK82ge8apPLepbcI5xMzKSjnWgxDI5Q8Ee+QqH2ruIzSWEbdzXNY
vPI4yiYTAfmpB0+25MT+avtXkehNRF+USJx5P/mLdFKiwmsM/dpik7ZIDqs7Z8mN
gCpPGaO+8vOxhHgYoLmtW499WM/lwOFWqenZL0+3PHflBb1JvgnotoChvedyZovU
9ZJALA9z9yQdAcZsgg/bHQFXwxOMBapwEyhhL6nQZ/YXC+/hRYxkZY2t7Hu6+Rcj
trFiHrKonBRSj7BnAXziH6XK3WjcGcw5aVS3FlRztiXdgo42jont2x5zJDAxWcXN
NZWsqroGhOrDxPZh7yjNKzhK6SSe0v9asEMSD4nY4DMHdWgQ+ZE745eK/mqHRsm5
FqTX5Hg6YgjM1bhIqIgK5Ejrwpsp78AjCfExRkTDtfTKcT75uBg7LLK9UstPWNu0
hh3e/wP0Cf/Om+stsR5SlQxwpvatQHCzxUTWMpj5zSR3iHtIRL8Dt3+jNeL/ZcHF
SLBRTJM3A5XSyEAj5itA3/nkCuaeSTKsHOSwFdMFBIJDsZK6r+j7ohFah5GLMQn5
mXHFXhLKqaM9GEC5Rpsu72ODN6ajASiiDqIfO1uTz/L11Tllv8J7WGxl5HSGOIy6
VlwhjQBT1Ecw+2pk5bQklKZQ2NyQ1kGQ3AO3G+ELPPcnTwTGr0VKd3lm3dpWz8F/
r+AANfP9vMArJ/qkGwz2cE70BdJDtQGmPsTlCk+XtQTW8hOXvr1WCcSLt0JT4J1Y
nf4c7MsfKIERA/bgCeqGR75//PLSi/9H4il3OHgg9wYe7PzllTsCjKVm0H2yVS3c
R4TeSagl46xf52ju5gh3H4LGrkKR/uBtLwkauzemqqi00fNNLR9tPKPPCANPKHNh
15FpAxWWjgQ2qcYDQTDnVd1fUrY6T8/ltM+rR/Pl0WPKmGE4trQMgCBPzfFBlydR
WMYY4HnKN74eCrX/E3BEW1RnWg7nTuv8HACg35yI3mdMq2OiKhOBsjVLi/iI6Udb
S856OEGk+VZAQOf6lQS8iFEBRsVGuSBc5xaqXuSDMLAZoaea4bm9XE+dDjWy48W+
JDu/+/pIyf2sKFVSjlRB7vk/m14cW0vWxYnw3ZnMJe8WudHXmgjjCiD60tEj+V5B
W66mwQOIhNfvzZMQVPEW9+OmLuQEggcBdcwZE3eo3akIS+enRbaA+89Tm7YTg9Td
qRwemj3FTarwYd0aabCU1c8201UyLnFYwfxZ2UJoiE9H6k4Xvv5PA/jtFMApHPTx
T+FtQpySO9K9bMD1IvrFGiyGGyvnVNLsqmmK3qKX/sKN6dULFvrZEIn7FSGu0aK3
X+rTc6M6wQMHXuKU4MEF3qgb8esgzKGuqhOt0wXgFrSeioBOb2yRwSAy0MfUg6lq
PxrCHxsvi9b2PU0bWmsmtUfPi8am6a/FLwN6XWc3MQxS+n07CSEDJGor27l+is9b
Jtx0xNR2YWqGgwMRUL9fxjBfQ+Rnp/knDtgkqxNC/xHYTn4UnGz9oPmQSjrDbsPE
+XZfsT1JpXwdGqW/u1HWeF5FYaYPxTteZGO6cOn9jv8QDXzsFE7L+J41FnSA01Eh
4b47bi+cpjieEHfvtHJ5Mu8ubYi2mIPxICroTleJn5+BDek1x3uzXXk0LC5SrVlx
F64ln6TS0UWxqFQQy6d3+/ZNbgkW7jw9WxUW3lFNXvu6fgddaTpd++UhNpBZuQmR
NVo76RmNmoMEfZEaBkg31Dn0uyEP7FHqHzhenXGXLg60gLuQg/z84cyi5WNVyCfg
DKDefuVN9rMZX5hhQfFEhWfV7NC42pNbkNz31M7mLLgq1niYrvwxqRhBs5NpBTKE
eBp4bo4e0YVZU67gnf9wU9TN7d8bR4pON3+/CcgV0+CRwI/13C9R/nHQa96rsz6m
hJFgejrcg3op8VuGZxhBrgCi5V57eYZlZeJe6TXheT1d+TzK2+J2WUyUq1iJEYNe
YkDpfud9OUfPybwjTLaGI9yMafQmDr9sz6rHPycvvWosFYz3je+b251Xv+LSKmZo
em5gp+hKctaJuLoEO2srAW7aP3s5gUoj706HliSpUDA0UAkImrkOjL1MEL2eqI0K
p0Bb/fO50bM+M91gG3nD1Ywv8FBI9k62pkJuoJNWSy/dGICVSdI4AJW6DOJohjKh
WsF3kc42IKT1FjBIUk89dC47Cv5wTIgcCQEnp0ChF+j9IzN60pygUXvnsWzUatN2
rwM0opotDmPo6zMbSkahx/Igllw52bsquEqsIrMas/NYdRL8JsD+s0+EgrFSE8Z0
vO/aEDqTpoTG8i8Mnj+a8XPeIc17LyU+9duamLlpSPN0HTjNlTfMjP7AwjMBndmN
pebpg+ogVl3ZD2wAXbYdE2bgupfgsJsV6Zzt40/1kFumczSLwUlBRG7JCJtztT2p
o2ohyF5EobTlOd7k3AqjYiZhoXS3v4i3PfiskRG3ZQaMTjyNlM8qXxTnB29lKF6f
mml4gYxCyce77T68Y7AyCUCkA5ba7wYWPUNFrp5ZsCOjh0h8JAsTj8p8YJMHAeGe
noovExKm8PrdZnuwqVAqvqA+HCBu5qSJ/tLtM83a1bW7p7Fzf2g5b4lBCNmtjNe/
8tIp3YZ/INLDe7J2jrl769hrIR7B0RVdmnSUQJonTA4ZVMY1u0YbkJGULfNRz6lL
90aBSmJgOUoLOCQ8718Q0NN5uF94E3lX0X1vryhSTTU/bnNqnM4xbF5s+WPF+5lM
tk/nng9rd4mT/bBYUpRLrQQkKlP3RmbmW176s+NMQyLzQReRM3XYJm8mFRZ6dieM
mhBz/iKXfQSpc/nNvZvFifBeVwXXzRLt50ICkIKRoh/D0/dKSCGCqdDX14uNIYrG
u0WhUMaAkshTvAEEFvb96kQYaBL6rNwsVzWsdv4Yg0ePPOwAbGD4aVU4EnkxrGP0
gs0d0lmB6sncCpl56bvbZyz/D+Gk4ZZVeqsV25BCykV3o6uKYCJvUopvYxvCPq+/
Ed3z4HR+dvjjZjxWQrI+bKoAHSWrKqf20VIQKQs7WIPEIXIL+maDtlO7JxEVY/6a
UmREZcoEWn/tvln+wQN9Baf2pOWgoFl+6au8lSU7IkPA4KMUyGmEq4lNULYuN5z0
XzzlwSYgfnGnY6qFKQgfKNAaP4aNNEt8khsMcF9XWwHsNFOXGf5MUPyOpWp3NBP4
PS1OtqhWfXd1nGNRPJ0yN+ulZAV+bYYludVeGarXA7r5dRSs62DQhDZztmK5X+Uq
kG21llgbJrl3syOMADH7u1VVADI4ZyS7LHAqEV1r++4vk63JVVRX4mFoFrrwvdkA
WPV6R+3nQ/Mh3aAnCRojRY0fQKmEudCMujA/4CnQVNjI1w0UPRG+YvFKY4EMmX3H
mrHmkWANmmlDNyGnsFc2cYsfD1qeYsH7qWF5LnTE0/2pBCDWy5PJrJ/jGxif5eUa
W99DiZ5BR2JhAL3fHP+I1anskt+91ikg3A+L+oZyq8V5qy6jB1kZtyggsPc/sMni
yKsR4EecTmuASULQo/bqnKk6HNidnGPgiLgevTT/tqNs59IgMPNrav1HRmB+ORw5
/PaFB0z98JzqHP+KXh52jhzg9wbnu7nImaAO/FRMJHV6rl8IBoM8Vzf1TJ3ZBMd/
17euvAndmZiCgJfrysIkW5oVs1b0YOcNgc6hi8CxZvsED6fl576mOmTnp79sYbP0
9oxzhRofv5KsHJ6tvhjWV1pkr2ShIuAQP++KqxB4SQ33UpT4+adGfXJB5jx7xN9s
Uaz8uBNqLv7EYKAezxwQsoscpfZzwYTJK0+1W5/BAFcGe6o4aYiMkOyyhcnLDnt9
hxjQerTdsaOyrTAmVoZfs5VAi76V1JC1AjLe5j7KA8RTlcTZ4HLMR7BTfQKTUKmW
SsZExS9gR5446oElGLKA5j3Yg3VbMDCYHoMzj68qZ2TckjbfwpdpFA8j6Txuryom
LKntybeXtL5BNMNoOwyi6Pdj9EiH6nrQWOVHvIxT5NoNteAtFL1vJQOj0wBEvSi+
vlhfuK4n2VmpPkALjUqoYHsskAj0UtHfe8tUovLZ+IyFqGx1Chhf1MRpAOsUnuuz
M++HoTxoeO0rqb1CGra7uKFrj7KthcM3wq4Rx/8PDqobnnl3cG0sSHWB06CP0egh
TXWEm0wAdwOAPLd7zfzZJELhKEJFpV9dbf54bKXQPvdehnkJ0HTO+RtPehu/JBAB
t9cPHG9UfuBakhBFRAUJHxbBTnRWd7TFcEeOIXY0UW51FBr3MdmZeUZEDu4J3b/m
P0mg523cuqqFXr7PtAy1S9Lolx9JOhtCLotAFm3hZWDWq63FUAoqgR959NOhwWX9
gk8xQ5IdnelSsIrC5bXsGkL4GKkTl2s56MIn/L34ane9MhZM5jIV/gXh1BIX9C8r
LCX/txeH443RykcTb806wRZg8o2Qo3+3tqGUc6r+zU0CgiodLNRAkJmv7o0JyYOH
vwltb8igmjXHS001fMm+HG9uGKp8jO0jwCw6qlPB1w52YKETK+Z1Y/cpFryQdA09
hn+z5xv1NB8MyBbSlEVcg9VpDrTw547nyjtL602FExf6nqUh7ser5mXZJCLHXtiA
VdmEHy6DcZIOb0ai1pSPi8qVdhQs1g5Jyhtxenihwy8PCX3J/41wc2JEkyHXqYKm
W3p0p1HlXiBZG9GO5ktPoihQrjNiypoctJCRV2cn76Vy4IDcSdzM714EeEyr/EQ+
27v7LSgPprc1nNikbmjjSxMr2gv4/5pl4jzEZt4UOs3qdw63yiCxU9DMNPY2Xxan
oW39WbG+IpqWEefsaP3s2zJLG7rnjV/vi+Rtt+la0x4x1jq0LmHIY50B0HEeDWbM
m2x0y1aDGYe0eDLNDFXrfS237EetM8C4uywpKUH4QrZDWxxnYtq2yyVZjypjoDoX
xMLNo4ABF8mFjdcNM11fV5vgT1crs7IeVmogiDxBFccY+HT9KC9boi6VlKYg2OYW
F/7xIH1H+LQktxz9i9qKN9OcknTfniJMq5WOM1XfU+ZFF5xibPzuGCSMu4uEi3xX
pLxP9LYsOHhAgk3RL/ZRdwbV5ifnD8aTsllZfZLpw8Jytc2GX4fA4DB6YbQAcT/k
PbDjNYy8SaLwrU3lBV9R1e2+QnlZ4O4LhgR3f0K6tmLgXNg+DXF6ZGR1OEHBhk6o
5vCDZWYYv0zPtxC4RqphcxbibUiv+27nqP2mmekYRmMlbMO3/0/JBk8MCr338K46
EXu1xInRy4W52kPzlr2hwSlSTvtPzAkttO2NjhUbb8F6tv+SmEptQXCC1jxv/8LO
SOuM3ia/oyQL6qx0wfF5LQkkmZMHjnQbMflbR3i7EuRh1MG763ffWvLb2RhspfPy
yRObu6y5GStJwMlPM4qOxO2DY+Rn1mPEkPSqBJMgtpN6so3Fm+HxpbJl5u++jSv7
ryCyXND6TDVZxr/zdh9YXd3WO/gWZxPm9aDMBeutFmuIvg7zE78gf0Q8L98Znpy7
K1IRlH/pZ6p6wjy4MYy5kogShMai15s1wETZPA8ccY1AJj3OeN2Lhcy90S/BfGsz
FIkX/ub8k8DkONmQVetqAvv29uYc+uTOIWmWlYzu8QnZJyPPKtT6EGE9IlKspnwa
3KJ3YTK3aXRj8VNcfRMVc2mFhBRR71jgx4LRH42wYWUST/SUeITj3MAI2ZeXB5h0
UmcewqRDxURV6jxtX3RMXbiW+WY21eMomruLiIdyHiqwAbgP5fsDYDKFNxhohrBt
ulyTYtgYeCF0K1//bfscl/v/JH9CrhZvR8jLM3VXYdFUbTaN4UDuEBboEA1e7UAg
Qxhpft9EI9wjQugpnGNoZCEMraKpJfswRHkaiLfFGf+A29IqNI0prphCiq/WqFjS
GuTU2VThJG//Dfn1ZcRl0JjBtMmHmqtQvlEys1xlVJWiA+pBHF+iM54eR29eJwpw
Mgo4/o0Tp+hAr7HKkGLSvAwd0WnLuRjAdLWJFa8qnx0kULrZtT2jxWRf7ZIkG2T1
g/Y5v0IQnhgk7W8pYGSEs9hGJ3aKLR/HqfU5Xv3jJTuWjEUTN7RC0UQRNj215rnM
tbkSKn+3e4/tVBwqswtkH8AfNWiqYVPSoDamTmX6aIHrddz0sesEkMMO7RAlpuuW
Yh01VxUMRabiUJkOj11Ox+RZbMQ+472ggEBTCoAgFtDeII6Z2AeBvrHEqx4yAJpL
d9rZag2MuRcEKRZshpIHCGtVwyNp5DTukRz/vwe64G6Kj99VhDQi0OLbWBlORANA
tiYnIB606AHpNFvG1SnDJecc6y3Ujm8h0fblluSWLGiQMosYHsAk+NsqUfJBk2XZ
y1JFlDZjh5REWgmGCe8IcDmzPFxmOY9S7iiiBABNpCA3FznjfsuLPImaXhu2e9qU
/f/sCMAoR95tQK7s1oVCTBy0sLCUP5FbjLfjmIVGyHLmCAUvxEZi+MA44HBt7W6p
pEycu4v5eR5zX3uiNVET0Zn21F+IzWYsPBPZGWdmdtQ57MmBDZ7BvaPdQGPu0WTY
jelR6nu1Pjp7rQFNzmNyVKS1HCod8VnC+/tT7mZeysaEpkKSHezpUO/gCKssqnH2
ZntAZFfuz+vENoqz5Kn8xyv5AYEt/svRxvnG2MNCVQ8nlcSLzBVzibDqmVGOMhUu
SxWK0m86bEZ4mhwNOE7KpVn0bZkoT4XI2gVyQE1DvlVk6XGYK52+5MxIcCitJMCO
MVXcOAFEMHJ2F+p5RcjI8Zbtg9/vkAmPeoTinCd3F16N9UlKjmSJlWPRYP/KWIVd
xP8T+Pb6gW9UtaCbp0zKGSW9qCE62or8CqYW5vyIQWwv1MAPo9t6w2t4peLVt05S
YOfakVSpvGEjzTVmk0yqe7cTyj/QvudSFVs6dEdp2OtR6LZXJyqGh6hFrSaLx5qB
nT3q/0YWcVs9jF3mSpgMiiElTzf9UZ7gNYfKmtvUnX1qx5HjkbE4GzV6YWHGDbLb
Am6BuRd84/mdnnsNycZiNPJQzumo1naqlzJ0GW8N5pZoOl1oGj4MCS24x+r1ftTw
O7al8EF+xXhEQFnSMVg0GF6Umhr9EPj7BtLmDPUPz5hrcAHxQsrqGc+0XrQ9gsoz
MAz5em8nD1kmunytMTzghon4CbNnE3P4ld/04L7FnhqOJXqQ8+bgxEYl/HyWwQiW
HxV/Xh7s4j+O74l/aHCp+FZhf0f5bsNhuGe0Vz1AkPWJEAuoj5EGR5rMuxXSquXU
56L9dVy+mTy67fCHji5rp7vrdmM24zvqvedwjxa6/MWOuNlzQyM/nz1HDMYu/gaS
ZmHHc2Zhl6DsoVApPR5pjn9eDrWVBkR0kTUyvjij01PfxbiQ1+9Hxks9O3zivGpl
TgkKaXXej4M4OoVFGfrY90EtPlXc92KwWo6w404L1SY07ieuFTOuTgpura8mlzs4
8XE5Gix1+ecxURAHVphDqgD9vryewM1+emBfv4GVJjnhORJmATOlsogW7HUGN+E6
BkZXfCR0kFU6oP3HveJMOFm67qAs41kRnLkYRR8Db5E7GRDTp9mro4P/ez+JQ4n9
c7cISWGUJ1HvC9gEm45LligUCuoSJqKQWrrdoMUSVgNYmpmJlEIdSNlSnMYyVBE9
l2lH7fmvL35dV/kzqYzM21nq5KO5fJXz667xU7o4ZoANLYVkQfnFOW4yMv/EUp7n
Gz95EITefZu8ulKIUuVM4aspfwlkeO5CG8NAD139QZKnUODPrtAQtXu7H0oK6h7b
Rp0+qAUhmCNzu1qf6DAdzd51P/8q0pPOgCVX72OFa/X7sPgsKLUHS8jdwhXuvRgS
4KBRPVWg7bHtEdQitHC41ac+DMUfV7D37o+NalZYww/Mxh4HB6rij9wCLVWgo0EQ
PliQeoYbJa8a3dSZxrWcuMVnTdnNbk4Lnb+FtMhq+bwxydg5cZCUpvfpFNay/o8h
xoD6ALhs+gr8VeZw3/p3merzIzBbaHItqp+BXeEVVkPQClnB/jxe8//unOb2CE3W
WymY5BHLu0AkzHOYlDtrDMwwgsU/NORFMhClCvyuoXw/qRdPBcvZ/y0nUb1cJLyF
02K/X2lBDid9HoD6pnZhGS50H81H3r2ns7EfdFg36g+RiUaDmGni8Ypx2lTl2p40
HF4/RSaj6K/OlqoXZ4QVuQUtSpBrWiWR/TyS6yFSjnimjcUFWNyTiQVvZbSjwb/I
Wxme4jFiOY6HzoI7VWtKWtVX00T9833uf38jpmJiMVZTLoE01ru7BPskIb5b/3Zc
MOb2VMwPCRhAUfb46ZJxsVQQllgIQf1DTr+iU0qxdpx3s0RRowkK8JcKxqp3wy1m
iNpM821Kus5VZ6jMq6sxcj4x+84YdqOqbFsAksRj+o7IWaOmFuzXq8JFTEYkPqgb
nagIM2ueKcZ1eX07thTc/LoWbZQNOF9JW6jBIQyo8dKekjx00n3AWixaOimeklWZ
aRHbb8aL68exoJTfdPCkcmgZY/5PYZLTJaDjJJeF88R9YROc9ghEpG+M0mavUeGD
uO0uyflUfseiXy6Xai9sNU6gvzwkH7q62JVKRuAEZ3frsSgSD+edYBffI5qpI20k
+ztsntxvTo8ziPnMvnUeLT6er9swKZ9kqVA5G5fnAe8+k5Q/ALKz48xkKjKVP621
WVzVee0jpOclhpJdWEni4qJ+9Ej1e6Rk6rWdWnG5Zc3FIAmhkHWzcOPuq3e+35xf
U3NqYGKJ3oxnQ3Q9B6dZVAUHLp4PpUKNifQhpBcsmhi7V7W2cTcCzIpKl/2KjXtZ
7+JDHOm2L83LiIPhP7iVrwtMlblGXGpXbUKU5e6jP1nF2SfrRMZKAm5zp31z3i71
XzVeumyTx7tGIjrHlbazlnJwd+KgeNOLBMIk3cuMWzwo7gV2B2isqwagbqblf/N/
P7GffzICtxlmfYqB7//L5Wjlx2D0C5mM4j9wfcUqt8K8N9qbtcvYoWHDPhqSRM+u
Gsg3Ay284vKkoFdwXzYSKlZ9fELrWd42PGuBzvdl4pTVPruKe/FJL9Z+RJFrPR5c
3jXrRUZBdSZVumGfwleEaw89e3F1FS0/P3b/QdRO5g0Kc79sZkJnLBrY06URQF6B
e+6fDoeCBkFFFkTPY6mbI3dofM/fShE7/XxnYArR945RGpDQmLIqn0gVBRo8qXXh
Y2Zyio5EUq53bTs7talSYUU8BRpwRuMTSMhPfZhF2thS2NSbWX98Ypg/sZD0Pj/D
uHH1GMCaXrKCKDby2unBHBVXKx9FQxD37CVqIG6g6reMxwoQ4j2F1PfBoABXoLgi
/RaUKpUUI6u8sGebodNBwiXXx8nzrlIUNW9qnKOZv/zOeEuzWqkV7uQqfZIucmTL
xtBV5ILcRBkrzQ23UN6cErZ4dAf3Sq6REjCQdhOYwJ8fEA9AQ2RG1IGawI4KTYsy
WwI9iqximQ51wE5DmgcjaSpP2jpK8hjUNYxvXOkUOe5li0nXfEA8lTMrIaMXdxt8
8dEsGEGbYt3G6Q95KmJcGOpFw13WSCvDcKpvvJ9wbWqmsQ6YbH67oASFMFJW4NN1
dEWP6AKQoSZn+LDnuFGMaI/b843mQJ2MRiqtD9u57JpwxrSXSVYXoN/oQeSHmchF
NNwynDGW83M6RBDyrNqdZM/W142CpnQ+KAx0v3Y77xdXwgH/rB+8N9EOwVZ5r/N0
M+rkhoKZFHA3HrZhpBCkt6FubyCb9wbv0Cfq+08yzg2Er7rs0dzWDOb3pE2Loohu
QllGH40T6VFxOGo+kWTNS72XIZ4k0+0RSn6eOnEg2InORWhmaSnYzcnuptMdniCB
u6Sjyue04ty1+U3eo7aFQJuq2ZpTXGiUWzfHsV7AoG26vgKj2Kz5UelfciB8ZEsl
+6oFIoZmLANUzUpnKCt90F+azqgKNFJEFRQscKKvfAPtiKI/QzaK7W2mi7UdDtnU
D6fMwFXXeDhFdQJ8akcPBYjWqj7JidAhiwvsMi3YfA6y+oSrFeS/q/UmNEFTDRan
4sI+/v0dlRWboBDz+7mKH4Odp9u1xSy7kLVb0EJ+HHVNsgHLawWn2oPxNkDQSn7e
pQTTbGDIONCa2vGwonBP5vfA/2qPpB+uzJcLUpcKLxulnLAljVI1jqQBwTaug1Kl
K/R1AtBBDUTp+6p531mytlpnltrZ8oPZ/9k0Jz6l6uhjDJaHzRHv+vsCHnq4fy9J
fAnxS5xiAozNg1YB5MChS9BTy1vf6bVxgXkArKomfXVvflLRDRbrzhj4fxSe2PNN
/SWJND/wm8raz08CxP10J4vfZKTXB7RA8nv2Z5A46iAeOaOCUWZYICUcjSs+Qe/o
NeziqUDAFtD+ViuOTLDBoMw1l6OvqbOlDD/EXXJtBf8hpsXP1x2J/xAaMQLkWVbz
JsoObsowhwF1OO2Pvx4/cFqmssOEXtzmx4ahnN12TzDjIJcIdzIoYqxAgO8Sz4BM
JMHsHP5qx2AmPnfbCbL24G+rDK54aq9jf2+Svs8ULSjC6pCiYW1+av3jubX546R+
BILrA1m02DbO5rEFrJZEDBi5bMr/sLG1wk/QgvgLuhEVO/f/Kua/uMCe5hA93/1W
HZm3RpVx2zR8ujgpE8PQeArtMnfQkWCGMO0XHTleDwcS2x8cifaejhspmqawm+AJ
bGYCtNWbdZwF3+FVBHPiEyrN9sKR6HPO4UXleAXUHVGUR74tOJAKEKc8o2UpK67S
xADWKO+xSbJJ7Wi+I6XxGjzi6vFHCV5A8FRjHNEZhwAiCBsUfN6drXrRE6YrAk1v
SvTTOMVl/5Op12AysQUqdvK3JbrZc2LBLqXLHumOUI0TGvLcxnEOrSCI8FdxgyKn
lr+1V8yNUBPc4zjy+mVP6PBb5oTfHPpAtM3KIJWq7JcBsjoUzrviIKjkN9zB/CUd
rk+qnELMF2mMBH2lNYYyHrClE0+K4AbvBxTX+CGwds89DunmactCQsOtq2fqs0z3
p1fmd/bWXWS9NUWPqyVPlKo5mXA5G/9VwdgSUFtree3HMPrtpy8Y/ebh8qr2loc7
zcRf7RE2HomRWDXXvhP5xxxW8iik9Ygc4filJeq+5Dd5NYtBmNWQj/yHkpDim8u+
cYsktJChP6lcf4cJqFtDYvX9+y/+GQYPxTjhQ1Yubd+wvwD6QWuFJwxPneD+WD2H
KCAsVPzLTFc/Y6ACbKltW/NUrVhRzjHMqGL+ruetk1uMbNXOR6tsaDo+mgZvKFoP
8h4de4/PXhJ8EkG+WKbunZZVqK1uOcZINJ7iAyJwUM6ba/0TzXgz/DKvcbVw1dYA
FJLBAU/4a8aiKRVFVLDOYr5XGmZPebCvbzgWZ5txc5dR08jyEoRNdpjZGRJLwYGM
0dPjr0EmFOSvoChXNQCfhi1Rdtq6uK7qgqbXg6zM8C5nHsP916hhg0O4XQuC80w+
avekmEAIX5i4/E2nZqO4ODxSVtcKYe3N85TPhA6oE8k0FXGb3PU2duXRLNArB2rG
INrBiGOEhPVpfsGfAG/lt6zvRRFhwxXExifd7+bbSKtI0JT/LiMQTnujkMc0D3Hg
m57vSFgJO9R2f0Fq0gfGIxfSsoqTSpYJ7/3mrBuxEYfkFQUqCnSRIhw1dmtjyteI
wXVig+qIwAzpmH5555lmXICw2DcD4DqemGXLwU7o4GC5ue2iXQXw+KxmapbMMAg0
ZhXy1J2jdnFvU1rejKPVPejxa2+rk6IK05guWTcZTwMGu7Ait5Q/jLkdCG24GpwF
YC5M7FRoBJfEYeXacP1KKGlIAcxT3v6aEQITQRttu8f38GGZdZ0eDIX5wzIF6U9s
MSWjQfbuR7+hTNzgVwBDUngOfZmIQLk52mmh7/O+/e+vJALlk4ld1dxedZhnhI9/
9cQKb2vtJ+6uxYwyOQ8bnw/R1OM/S/JgTSDYyucBq09M3Yn8CxVzk3Eq8//h7HKN
CDPFeRUUxiFJ9T5yTu4wviom+g8VbOJL9J7NOmYkmMVwFxN2InUm+mETrmPRWsS2
QrWRkHSYkstYGcb7B/+CPEovLCvWRELU6rcuQBq1AHFgTtec7w4rzSetRc2nHI+a
U+oNgG2jkEYBdm0RIo84VEpJFafvKJch22NUavfPuuL/HxnNd68nVc7aGOHjaa8n
WmcQMLYdziX3f4BgKC93pb00zJ4cEMsEUFQm/d8rKFqPh/S3IvLwUi5JAyIE7xME
ElQg7RsCzP0o7QuTHTFr18pj5OBuQEgQX8tuWFjRTIbG8KEUTN/++Tv3pT+uE+6Q
QcNpOc+mHK4cyBfRX4figGM3N0QwtOGvHiWS9EIbtpEUFjDlVgvUYVjprekZWQky
BG+XUoQ0Ftzz5TsoInOpOk3acvx2xfU5rSRyd2szmJXCaTb/vCuvAtW1OPLAd298
I5fWUEFiIdc1Oq2vdAGv1Foxewj3x4O8kGkkL/B5gVO0x9FYrR0wOJ8JVqbIQfE6
PwUaCqigQQdynlc+U04dg1sR7ZCaSk/PeR87DZ5FjZXNIl98paQVQPGpNuAv84Yn
ehbi+b+N3c7PLHoWfl7sm7iAgpFn0dxX0kCflnk93Ostwr41DOOYH63ZWOyjVB3G
qS90IQu89brYHl0J966ZV+SFmBO1Y4XjuVu+LFria17O6Ay4DmLUNUUNtwY3XIcu
7514TM2Xolbh7RjhW4uR0AJ4vI7D+2kWeFw7Bbcd3fBzI7npt0h3bUSENmoknH9b
QWU+sISPMJYkRNcgI3ugtZbOqM0Bb2PYsMPQo1tkN91pyc28VhPrB58vehBMefDO
kbdWTARZ/cItuoEccXk80D3zHAZKfEjiO0GM4URFlA6Atll1dmHLTN9kV4N18CQN
zH+4YAMQuSeoaaozaflygL0CYfDW38yii2oxchxm/WEWuxnC4ZdVQL5B1C0OnI5U
fdjnrvtHA8qhjjBhTOrAifgVcsCb7wlWKCkBhi6WQq5ab6BKSMM3zZIiUHoveVBW
xB7yYDBbFmHRMNfk96lHAFkpUikSCm79Mq1yc9G2WPa2jtZmAyyp2qHVfenZa8bv
J7Vb3sfyi3/jKRJGn/aoiDs2+A9MBHYBJfdTGWn6AAYZQ9xGL6n5NbwEFKDTWVIv
O83Ncgh09uSRRp6EYCpqDKy0HrzwSCsQgTkMMzPUweSEmopQg0nxtmmAer3tLAFA
lpQxsOVvQtD5gDqu8/aV4zJYeZXbD3vvqhbUChEveTlsBGAk3Nyx08C+phRHyRAq
SDGSdbq5UYNpozu805LBk96ILajErXe1IG5x7NSF9VKtvZIzMdlw5SSfAQPUu6oe
R8GQyBIy3RoAE+dCw3tcrOvyNOy07m5XVgkHb6PTQ4W8wcPt/ONrvi0d6STj2N50
zvquxOF7rp35rDux0D2TWwYZ9sG83vHo1J0NxHBFh+knexp9kAya7t354L5ULt6N
V/bofoo+2gTL+bDx1BSDMscRrn3WghwvTZvHnv8lO4hpSWpctoacYvSRMI9htptQ
Obzcwq1s9P+Ekc/gDRWd9Jqc76aQ3rasGG7SXMXUzsz6Hh+nhp8gcS5vI8QG86up
kvfDMSXNRyDEfIJdOZAfkOyNbungPe2pgAct2GlLB5tCm34q4voSHniU3HUhUIow
8QnJ3J1Q/c7BNndIJ32+laTpXKDszsgAnvhYl5Vr5Eik09lMRXbwpmE4KuAhxyoY
jlInuljSDBJvEPbSHj3gh+C+2fT6O1tD5G68qRpNJZLXaZ51JKwrGxpM6rL8QgD8
OumQFFnWQfMunsa9ZGuswhr7y6SuXu/a97Ws/nr0V5hqB0Ae7wyW2nbG8JqQVQ7s
bGMt5RvPCiG3ktsUrfsN/bjQ7C3wEhNyB9oE6UPDtFB3vUDJZqybIAvCUY8sMtr8
3lxQtdRF1V/Jc0SkkV1hIa1Cb23Dm80wEz51b2t+jEQh7FfGUONkWsDwEaAtYnL6
u3JBZv4q4f081nGDW0LfOhfisTVxeQ/8NOjIM9ggbqYRJQDBjCW4f/VOfWbc6stW
c63KYaR5AawEZBu2T9HE84yCVGtSKo2bekcnG4OqQstVxe/8pJ1pfG996bxcn4Oe
b7j/y4qNFks9YcJ4IAT3NsIxa4sQDMy/Sh6XgrE2+vVfY7raKlU99V8I7eqPQ4ul
FypKkr6Jk0m16OjCySdlodbEqJijSjBlp/DjfVmOufTtt2/ByJvjxvLRdrKRpjxE
R1d14CabhAuXg27IaHwQHpGMSuxbDhjURR+NkBTNXXfUfNLCiz+9yfETWr0zFGVt
fdZC68Le4JflsFnuxGVevBIKMIB3QgWmY9Vuj2SmZIac+f4apiZ+rqrjrgtEndT5
fknMb8KrNj+vtSkUFsvJulyLjlDHysl1nKNb5Hu/kCKc81o6i9LqwcU5Bo8cgfh3
+9Vy1ab9q6omRxN9UI1Q7l8/TAfsYzyaxdHAZfX8f2QmsvHn/l9QDXpfOEOJQqUC
ROU+ie52UUZGrJi0okgxlV34XX66q2oyBISS0xHD2OgrY06vvg3li8/CUYd1Ud0h
vN98D97oG9XCGbKo/iv4Q678IMSXw7iFBIHdAiZAq4MyoMoxGpmNKS07CgiLYV4K
jvrHv+0MbxVRX956qorqY28MMU6e3DU/Ydem5kHMyUTvHyBqS/GhMFGSe9Gs1eVc
jLG1j5LYwZ2+PQqZ/+rJY4GfH9mEgETMxnaDWYQH0yTZVFc8SdxNE7Yuzvxt1xWD
vQRGvaS099tZP1EHRXKR3WxtMxdQJtHRcOUKVsP4E5R5WS1ic5jSbXb36cFwhW2T
mBsL1Bs5yQeJsOHfO83BCxNo+FUWYw+XQo7DgI/aCxpN9AWYAjUp5HOtmiK1E9WC
03DO9ycXbaezaGByoOW1L4bJit4bdDgLDU2Zrhj8W0hHJnDxrXbBp+haICNW+HjG
lXf0/oOc6quOiJsv6zGL0mLmRSN+68ZjKYoTdrwbyUg6ZOHD9Ek6GXvzVQ4HlQM/
B0Ns7NlOImVXyXdjUTAc4nwabXrQB+x5qJcN50+YIF4kdpdCIVWI2YWzrLZwk/Bm
LuDzEK0MjGGld0VKnXzd2IJEtmpQQMZ8/R1K6y5m4RX6fQAMCStJSpKBpMG7xrTa
6l9ktixNSxYqR3AeCaUeTAcNKqDfP28yVTdnx43Ok0bdmhAX05Je9hWudu/VTQ4C
smOBHIlg3fe01m1QuQLVp7LvbWuIYXEN7H8cSHxwbYdug2G1t8PVNEfg9QtTOc6H
J6j1VjxLFWIlDLPO78N7YW7bHu2PfN8/4Q7DPxejWuFy9ODKfCgU4iCANAcjYhjq
huyctdfsbm3989svzkThXWAiFVqXbN0TD+lnMh6CdLmC//hevqqomI7vIpcZP9/4
JGVbUVO4vGk1kUhql0xs4vlFuNpCuND6i4c9UIGYSWoOZgSBt93m8LPR/pRIHHzL
p26q9VRWCyh7xDOhEr+ZPCx7fAmVKUxKUd3DnT026uCTk5OJxj5IYfsgIsvxndt8
LzG139C0vNu9Btvl+raKvW0hIwSVGdaYDWK771E+tBQwfYqGmZ04MtHhONXXi989
xZUGPk3CFhl4FtwlPCFHk3nxBJkznTr2bAwzOpPJ6p5Me9rK3lK8kdwWk9I3x+HD
8qKmASpTrad/E+hhgj65ZEz6+0UO6DSDFcOHfclyNAqlwJ2Sum1wV+2VkxAVcFxr
efK9b4qhU2Iv1LdcYZMk75BR7N8tUNo+Y81LQN5e6M3OSxIEX6PlibDYZhVnv3G3
n4HKKWkyLV25e1jRmIWrjL6Y/XII359AbM1j+8Gk0CjzsOL9Tv3kNPQgexfO7gOu
zW+s3mE0sk8kaj4YiGEIv3ShcGdjfpq0v/EYroRI7+BjbqCHRehInYPQSMqdO+SC
V/5ff3P883zBxuvcBF5oO+BZtNPMxn9XUSWt678FpC10a0sy0suard6MDw+kVIg/
OTItjlvEhaiGccDihiNdq/m4DjbOZxUgHpW/Q5TlY50ifGSFdFu6BfXtKzOj2n0y
rnrC0NeF+Wuan/MM4jXDwKEYY+K83lmgBYzf0uEgQkIdjuOBd44HWGXSqBpY74wh
2qbwmIZqpLV40x44TBtKG5Onz3LFuPmX0dgm6L5HHXPwQkMyhSXsBOtQJE29c3vp
Q80cvt5lYX0zJhD+KNYbD2C+yl+vy6OyY8XMG/c6AEyX6WgAQdNcVMqd2EQ7Kvs5
kKsFAqpg0COsTv0rq49pAz1OuKHgnRbL63+vsF25PxTEINqf98nQzvQqPKj04y4W
BomSMDQwAUY+1y4eDG4Jvc862VBY+Q11E71NiaxNxQkofnfUQr4+FAiAXh/1atAB
Dg0AqB5DXQMdlBrFAsdADZmv00va2hq7aR1c9U7fqmBzVfvFGZ8MhMBdkJi+Rs8V
NkwNZAeRrO6UaMzTYgUjLP3falISNfnC6eoSkqk11DzUM/sWXucq8Z7d7HTjFqTn
xmCu0ZryMTHJAoFHq+oYSE8nCdgbxxG+fUoSTy/nlKzO27vuAWB6usQnzz89hbJz
cmNVda8fUe9iAJ/oRXCsw24XBDFPjOXNcdFoEzB8YW1K0yqm8s3ry4hVILXktFAK
M6ZYKyyldP+nNCm768rlJvy+n7p3B2DHNWzsFO6vgD076ud1TNbMbqLXuw0q5nej
hxRgzMey+LPBPf4p+agYFaK738sHB+eVIv4gcfgIuVWF30n1eBqvtNuDTmmIT/Je
f4jWBDPz2k815q4FfsN0+KEoR3TzieAl774xREoX4juqMUY24+eT4lctDZoeWwqf
9PCTi+mIRIP26IXiZAf56AjXlwdZhn4lZp+zLmfTL8241G9SSKjj1x7nH17LIHDQ
u1HUhZ0i1MLDxMuCeCKJRep8KoWNcOodfeknzzZFb+TOfpx8vkxc4jUXRYObzPg6
Tc4Ue1dpttzErjgIWD1oAYGHoN1uElsXpYPZQjC56oRdQiWxtMomoI3S0sIfNAKX
yzJD+HlGbOfSL/xa/NE++fbHVOc/4wnA9NtOV9T4saYITyw/5ZJ4msi1JTeuLhxn
GrTZXyku80t24g/yt6j5EC8iBRDqma+De30V6BGWPXi2goz/jRpZkqfzAiolEM3l
Uv+ew9yCawiZRnAeKzIKBH9qdH15EvxL/9y4H/fv7bflhTXgjmqnuiHjbDc7pTQ3
Me0rY5v1FEQypXK8aFivx7gbLUF6SC+rEzk9yDStTnb3XTr3RWFD6Xhu9sAjANOK
Pms0ZNs1RyStZ7JLlIwYuM3eK3FUQ7eeJGgv2Q4mY8quCBrMv0mVXLg7qHMgigtT
nYmXNWlngJeh8Cw4cMlf69PetccMMgPZWm7Hg7hKEtJqXabyMDstm/UHA8IVWGbe
/n2nHprDyFrrG76EugoBzL6scwqZO1gvcluoGhvIGcegJt1udPShKrhhlYAPCMnL
z76eS6chholAWZeUu3Gg20llbNxtaXvse+3u1myWK/79Seh+EHriEwidnD7H/Jzl
U0zN0rhcMV2WBiX0K1Tv7rcMAdhuN8UV5J8HMPpmbCwyNSSmupeVjtnjr+U5bKLa
6l+EVfqXs0S4Olp29X6/Vp5nNIzy86vnozzvNRVvld6ai2ndF6F8Tk2Vt0/d+CZP
uFxx91FLKggQMqEfmQi4RGIUdE1sMyASTALR1zzxDPRqxVh4bIKZyG3teaK/cWz1
fRDQc6UWaw/kbmVGPXVDywRcm09innZC3+vIM4zQ4Uaru9LEYVrKCighy9T0wCFo
VvurXZGmdGC4ypsXQJYbi3tL8yQlcyjccKFknVQ2c7rI4RTokQaply6MSKrKMc2v
h8k59gPGLzUFo0f1ud3e7OhbFTtJoUwAkFGCJ89qXMk4uzplzEklG3cjC8wVlN9h
joHDDdAuFVz5HV1XCN1WfgXFUSgz+qFjeKSMxNjjlkJa3Zc6c6NbJv5RcgoQmOS5
3IFK6lHpZ60bvtqaAqP1Hpj0liMkMtr62zFU6OsMxnnilH7SFGcizU+Gw1KVSGJK
IaKZzAQ/k8DruUpppx5QdqCjKREdDewzCKrjf08VJmRNxWphRES4rH4Rbr3O1A6Z
BtWp2lV2efH/bnDZ21kMGmEKrdoF9O534uoWi2w+8wQmE7Jwhch91tZfR5T6RdQ/
UGuQqS69ieBSSOcmU/o9g/iw4FeT9JPvwolcOHFyNgBNHmJ3JfgowAFczuqbtpRd
oyHiJCPEXN0S98OwMQqsQnBZlKOS8WfE+XFKnLeC0iUFfQFTdQd5Xc4Y8A4S5kP1
4hT2YLXlhOdHno95GQmcEt3WRLFnCuLLmtlD5Hv1VOJ0i/VUkFS5Qx3B5knQOpOj
kgS5OL/6HeTrwbNz+PVaLLPp24k6+BuDgtNv91V+AJg4btUNFUCZrhp06dd+YSEg
ws3NP9Q7vKVErx05oea830dgZFJe/i1bSBO/sMFyjxR5gxpLOVOUQJn18UHoTrsz
DJ8SimJZ2iQxbF2R8XXCunzWu3ZFXNgNk/yQBrF6vGhpdIiyDeR89kPJJAZrNzT+
aVaqTrar1YAA/Ar4e467cujoFS1dvgOdwt3zQ+pvI0OYBmwvLUFu9J42hBXk4awH
ysNpsPl1a1GB0eOy7gV7tB6PNEXaLLdk+oIwImGQjPwR7X8Gl5XOWWbdV3qtkGJi
jVYbB8YpvWMtB54x+rnrsaXhBCaBaZ2l7KbitT4N52x036MoHjFNVxpxdm0StdVQ
TbLKC071Jdw8uT41Bs9p3e2oHiukW8R4zr0aegJe6aksmuyidif1ohgy05x4W2ck
4nAzxe4q+V6jApTlivlP8e1Gs5vLUAKINrw4lGviXWYtR6e1/w/G0c7dn9BlA3JG
cQqeZK7hFarMNF9lO5ojqAVJHZmdxQoEuMGRYbEjaxr4NaMj6AN5xmiXOE02Iofh
qDQHEdevtdiMuaiEKkDsEaNK7ISZpBW6BAUqwP71pvtSw0OQw31Ovl4CMV2//wQt
1BfT2uhVMESJYD4C+Odx11GUoBZJOHSVcgTF6gEovC6LQ8d6eyP7j3Jl1VQGqMCm
kDY08rkjtTxEkNFvRzF1rpf0nQMGy068QkPXjg/1Ug52m4DATDR85bAhBkku+2fe
weBY7Rxd+Qp6/534VYpCEDg6526godmmQ9bSS4ETyLByvgWZ616IyZrgfJHqLkY4
X+zSl5dncWZxtOPVb+5CEiqYTxU0Ka2iNReEhJQBVbO6HabNKNkDz95W/Jm9X7bg
rfXUjSdEIS+MZSKzqFJfTbaLxQoyyjHrkqwxhZn5uGm0fU//V4RqB+9gUQbJ5t75
hyov/k3ezJGk/grfhNUF4Y2/C5k/GbF645CN2Uyv01iZ8+73VI2etsVk0Ph3IuCZ
w4fUvGfxFygBQzWRwCe98bN1xpLr/VkHG0xDnsfuOxSXb9GJ66BrYkYs4SX0plSt
vLT4Ud9Azv9xtDiwWepRC8+Rlne1ZgCYZo3pxgOYCDxUUa2ssuQIjvaACcbNn2uB
4VsPbVLLZwSt/TeGoP12YXZNp+CQmRKLl+QwoQcw0qcy2bUCjHLrtmQon6tqmycT
JUFXrBfAwlgzFKL430/xsQBjBery4oOdNZjriev80RSax4LlVr3MG3vTvxyJnEXY
jtVO2lqOh68NXC1CVnp+7qwSd8iWxJvECzp962H+HViMQH9Q3vu284YLM29I7riB
WabWK/7jBdiep3hs13CndCMAwKnJd4ThRi7NKYVcTge0EGhEs453pH0PipgfYH9i
K8m9UAfdHFIs9XGDI5hghnEkpq6nobjUWQF3TLCoNKjVbTmC+9TH5SQDnRty2lX/
nyHdcr6OFZpFbwckSBz8A7u+r6kUFmoUGIkhuyWIRQ3DmreAjPyuUwavn0aa9/8a
57r+0koUfMnEd+obDTBEXil3db1VzbYVIDrH+GXhzzY62VmpYrjqxx8RshKOY5Oo
FnsxYlCP1Tt8UjAL4gBr9ENu2ZWpSoy5Vu5MoZfHBdvbwpIHMMlcQMi2kmtAXZlY
IJdkCwj+GUispqi6wIPHkp2tnlR0+lrOEWi2kHthUtzNIUrOvcoR+Ieohurk6g9K
sUghWShmDhnrGi168OJu7P5RCG0gaBEb2i3nHhCoa9BEy+otS74ycJH+sMBt0XPS
Zxi93Tw/oIlPSjAfSDsfU1YxPaxhZVGTRlvNYkHGcROvv8QTUgqY5/+xUzPTEMOW
bSosRqGC0BS+XP34K4EymZs32P/Ziyi5pRr/FrLffvvPXMgiVDhPwaaX7n0CXFVu
E/2+wEYheTArDZVdpetZQI+JP6fdzcOeceQuYxq7rri0mzgFvRAv3w+RCe1sMwCr
CtYgQY9WW7DUEC52Lt/swYSmeQeFna6XbdL6orncLxdFvaZoZoMb+G16cigKlGCR
uqpFDcfgYpsy+pKRvsGH56bgbilLVE0JlZ5hP8J8ZDp8Pa2kfN2MGAIR+yv2ocj5
feM69GoMV5i4GcKnHa0O8DP2ZuLfB8TEREsHkKdPaZk4WJItsN9waRxNc3Mt2fnR
TvQp+bHnbgMG67SofOJe7avE55Sa3Y1noF0sA4CHNIVJp1n+h/ChgDpCrt26KPG3
ZX/cotMspTgeOKfqUpoISyT/Wc78SQgvDd3QzmVxmdh+UszksWrQ8Tc6x2vgJM3x
kkHM7XMhZ+plZu3UmfoknPzg6pmVvifTxi3xdy8F0b3rdJzYogztTZzZ2vnuj4ek
Yzwgi1XsdQ6QbOswisZA+y3MVUtDKjm0LyqJGcsSOBP4zjNn6RA6glt4Oqr3zB+Q
ewu0nuthtIRm4vJ0B/R/0tukFlA0hpHacJRlV004wK2/us2fRMBSWnLlwkKWdvUl
h9BjA5oqgwEfKpDZHIoRGCo8ZqUNVDFBgdmkHG3llo/UodTFMvO62NByHK5d56XQ
DoeC8Lkk94p9wNS20gRUXX/PMv/F6z8ejsZMvArZLLARFxyXNmwqQLsfMTiQx0jg
EZ5RH4acLs6io1IF6SPEWgH4ncUSJODnc0sygEVpGR+VtXVpX3x+M1WOk0/CVfjz
AHPLubBLixWkSzYy7/zyDAJebwXR5PPtPuHdwHudAUb7ujVFxCn6CZiXTtkbGq4R
OquVGc0cmoQCkIQKSeTtGenp2IKDa+s7Vb2LciVPnQqwNAH+xrKm1fJXVKYT5wmO
+yPoRjND/ded85034lgZ9O2FpGtShp6hvI3DGDu+NuU445nt4MsgQhttYC8OUr6M
DKeN1l4aXhqPL1lcQbrF1tI3F5UL5zKve3Uhu4Aa7bZF8q8LhFZxS53eHRqckFAO
P/qVW8N1bT2LDhnquBu5pg5lO6rVqnyB3oOpjbBGNCIEftZK50kGJjODUESzNwG0
vjBnchUIC5s1NvFLZf5/qe/Nk+By4bUUkwvwBL5ZSLgZ7UahTwDllpDvsCGwi6WT
gyuC94Z4Q3nMdNhir4xu2Vy0+Tcqv/6UXeE/YYoXAQecro1BSlyQq83uEN7hkOzk
Y6TgB7YyQV4feDo2cDpNhiajwE3vCGC+OTtE0UQu5yMLYyYy6wPqcipQrwAOfDDc
LK/fdUCMZyTJhc2WwmjKfA/JKLs2ofjadM+JRxrb6GVsdRMO4SRJDJUVoAvDrAwJ
1bsHJbADzDDTHSTvplVWa5o9PnW2ZRbMD5MwE/UTtUV1iu9Wly8OG3EFd+iOu3nS
6IbtFmhOJTnhvQiYroUMoKj5LXIVY2Cos56hmnrQKFxBxDdnz9Jv1hfncadZhywf
quMtliAXbiT1vIp8whFc3ndoximjOVcFdhuVFWV0Yumc3Cw0PBwUum/N5bSsHbiy
JACku5o9QUX8s7bzOJaWXJCFrPLtLC/eIkTNUvkCqFaV67whC3D5x/FjnQlmCSgg
A3MsS9rzd+KWzBqS+Mh7+rKgAQu1ct6lwuIsQqoXAWvsQvpjjbdGv+dlUaTlazf1
qN20XDM4NMax0U86ovi/3K7s3aELRl2znOpF+vvD9Tulh1P4O/qb35Tt6BhgubVj
xKisxYuyFMRW3B/V3lGn0S6qZZUj12BShy7Afo608yxfodGbISmj39YG01jezjwx
vMgtF2lR/sJXmlKa2N6rcs/xsfdTtxzTLtGqipWY7C/gVW3SizfY5yD7zAlSf76l
qD7eTxIwu8AKT+yrrOgWxyix8QidZ3MAMFI8pIl3gtKnoIwrsWylT4Zdd26oLxQr
WCpXk+pRz5aRR2+Qr7b7LuxQN8P8WaI3gpIHg3y7RnU2KVAgNL7q1f+wyTD8MY5P
ixTtEas4geEIIDbSD3NiGdYh5GgSrBqQu6L+ogFG6NhpUN127qaJwqnhc37SGkG1
PPl0t9OCS4ZN9iqMzPxeByAnmj4qNS9Lp1DMmmgGaW4vbf9OfsWpLmMzjaMmnLBS
zdmGx4lznC/tnhQi7i+wVGwIur439R2KQma0evxTI+Fpcnr7hR6zqdSQQFq7aVb3
vhZuq8jPcS4j3+hPaCEmScpeUn0CfwhP6P0QF7YEsSoJT9cmRozqGJ0fOqow3VDK
XVexkgGrAK/mjDmwmbWpkboXts8SH+OEBs0yqC0VuBqkXIkl12U1wz6r54xDOg8W
4bHsZo160qlXFA8TyB73MsAMgOj0GnHCr3UxFWG/tA9HXBzkNg7ZYGU/Pwp1UXY8
vbpSUaqVyKuWBy6ev2rnT2DlkoHGGGG/uBLeGRcO7gSg4fA2LIZzkMmrbOq23FPS
G0Dmma0xWn2Ll1qesWIzJHJAR5qLAjOp8o2aphEAbLZUTb8KJ1HogwTSzUEkg9Z5
Yf7ZC2HQvygenjvr/mk/kvaVdqJ4G9qcfMHOzKBy7QIFBFysBYMymbKpmiDU0kmV
ffMqkoOGi4pNkiWjUDaMvEBzCmFTS0Hg3zCV9fiEK73k4c4cM2yW7teWv5Hnv/5r
7PotORjzCEbA3BSdti/Pa7UvPtLvxDNqS8g9uEtqE7hzB4CwxOAWuu5covJeCAeI
6Kcr1TBEpKKtGZMCuFHISucJM4Y2m3eCOqS1yUQH0rj3dh+A/ndpLo3aKGS76kH5
h9FQXlFJzvD6ngfI8j0y0KLOzkVHlf4shW3ETDz/QPQXFTc/9hUZ+B6d5sTS40jO
v/Q7Ck50OfdSlFQNpom3q1dqgwnO85VxXvPRViCEm44b7tgltBWT+iKOnO6n9i6L
piEmc/1s2AvpjgdbjmT4BYWmlt2ftHEtpQ1eGiYQFVwCvoFtAUvCMdmD6di4nmvu
YboWyxMiKvbLc6aK8K8lsPjhzpRitlmw/6ahBMeR9GDpfJr3YBCzonLRS/D0fv40
UwFz8k/QlziObFKaRr0h4yRxBjSsunpdXl238FYQ6P2YtxAJA9IvAQAEUX5EV5gR
IHQOWwl0YCPlH8uVBLqqblJ6LBSeUJU4hcCRj/D0laNbaq+L5rwHIenyuErkmfnW
VXMrTJ86wNnNHHhsxyfCbVkkRbALYVi7MJcTB7Tp1CXvFN0DaRpcqzcSCwuzTNj4
43tHldWGCoa4VI0iC1+nhliL/LDkyIYoaLmGWWm1sKil5OtCemEJM+G5F3g12wto
j47xL8HMZVkVgVkXvHsl/YNPoYP7HAhOOM4wEpBTL4BMx2y1M/PWqH/dThdOzh+2
9ehYdyPFMk4Z/a3Ee/A2drAvBuUalgcQ9uOObPzPJ6RuKM5NOznmSwMaGmQlm/n5
4S4ifWmzJZyJcgQ1YlKIqrJKNGoScB+twygt81LYDKrCkdXtKuVIGuxosiWF+xva
sBApQVDrUCaeBxsyfKSUUfMknjnyRk0gmOB3BYD9LPhNSc9JgK63GZ85UmqxFrJN
DG4yweCzj808frSWXLKJJcL2W/WQODe40ffNVRfV5DqxW0hOwWBhNiW54Opq8m9c
qAKV0TrgF/ze+rOtygNVjWUmM5+mMLRuUn7pqD+sm1eFldfPJkuazsXcuU2EbJnu
1bzrKS4m8X4+SzvLP2YbXi6zuzfXoLu3IKcgwlkL6x+ABWpL/0HloN0vHbge+nR3
g+op6MaLfB2+xLXPJ74a9A15w2jnbuuRAnGi99YCqZmGU4D5ZdwezuUPRPbK3zv7
slAXyYNZOyGA9Xl0uyTVbc85WsyodowJxVQt3QYgiPeI4tHIAhGolhsNsmdhPph7
36h+TYNMZ18zp1K+/NwUOTiZk2xeaKZ8zsHSFeP3VTR4SdKt7z/bJ79eFztLtGZo
cQwzkxb4IgUKfDhTf6mDpL0TQGkByDlwxh9emlBOR9NStUof9o3k/1yoTJ3nJxk5
mDxrt9BEqqfzbEpAsTO0Md5FtFyFEnAaHdDc5vcHPV48msday39jBJw3T06LA6Em
OmLdjIPoFoqukCplAD0J3oiDCCT3Fy7r26rNnePhrQ2yMirihrGcEw/5d7NE2f/k
csdMyBFv8qPjbd4AufPvPyi4ksROYmel4QZ+wQeg+t95TxlExLI0be7hCjI1iwpt
SVb7RzHc/QViXntsQmmS9x+PzYtmdIzur02pHso+TKlSV3pquqfv868VlNXJYCj5
Zo+aslhq8Zw2pIC8xsWFuu/IT+JhhG76GOsY7Te46ewp+JMpCxcBF9++6Ptz050u
nxLRXGuzwbIPFp4Iar9yNbnMOs3e7gOfAGX5FAAgnvFwZt7OWqZokQrj0jIEfekv
rP28jnJlrTw24UOOg4qP4GVcYpdG+Jd9671kTFYAdK2K4sJXnFjecOUnc2GyYG1H
AaPf8BqX6h4H+xE4QAh5v2p5rUTNEl+O4AZ9qYHF1o5vQpzAtdyGhAKdhk4PqeqE
cI4TVVXDIlFpy66piKOHwGg08Zw8tgMPr7remZXsVdGJANg9ieI3wzQtAUYkKLsx
T+QRjlkmhNjU7+6hIiS7ANE9TtxhtbpVeeVKL8XXhrbKUXHmSnIqCiE3yBSv3Myq
09QEuQt6EORrSr60QTrJSzZGnNj3Ut5J1Lj7S0q97rRwqKvYGsle6zbDLncj0/NF
PHRcrv4Z8TOUwvnUZEPqXNB/xuz+0amMGGYO6T/QCUkYA0UBMAoKHxgfBTomXsCh
QrcQb8mU7UtENHdodj/ALrrpIM117EIJKe1NcvjZ5OeV8D9OoonrQP5pIqkPZo5f
ZbtruPsh6NKjBtnuXYHvAXUYaiLrb6xGIz1wVN1KT2BJT69Z1lghj4Z4CXnP9yiL
qwop1ibqk9OBG1tVeHMbWu4+PBRhP7jung/l0no6VmfhM3i1CSBAH3QlFrf5CLm4
BvVAPQegeuCKh2//rPackN3LLouqGSD2OFcYEbYy/oE=
`pragma protect end_protected
