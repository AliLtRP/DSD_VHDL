// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cb1SCgnoogM9KT73SI8vw0/E5ULun/4bgQjYN4GqHf5FnYjgq/1uW5mDiC85AGr7
vp5vZi17yYwyqW+yTkr3lctEXb/+8l/dehNetz8RqHM0THufZE0KE79JvT+SF0Qz
lIhdKazbpOtKMDtr3wnnde3DoYRgXvwOIFFo9T9JwXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32944)
wvSeyGQwgnWm22Y495V1hBIPkCkzQm3lsBfDSm/ogHJqCUP7sggOoskjdx/pdQg7
ZyzodAhGuXkWF3/PAcBgvB3rW6vr8FJe7BQfSRepkUDRl7wmkHgfAdqW+3vefjfJ
ldEaBCntxYIlg41xgjLnG+yl5IngM8kvtQBPbo6GZJOIXUQ00JxWlfqk+met9wPf
iQGr1UBENU1RyvJQvKhnXK0rSFw5AhvH9U+Bt5CjD2Wx99hOy9hu4ihX2s2s+LzM
udlQBdMVzLsPrjppxXlLvBvUB5hyqWJiu4xUZfoI+dYBfD5n8JjIpWpsEqSZTHI3
h0CYi6O6J4uYIIK4u879ZJy2nStfasuzAik4oyNTPZuGaTAGU9Yh8Gi9TLqGnXXp
t7uzt816/gI2YcVTQVelsyMXrB+NPWNClR1PEqHV3DjF+TZ7PALHOLhrPW3RQRsH
3KvkZ1UPsMtoyYF8+lGv7gYBbBXeH6JrzD/yJb/FMNI0oAYbp9q44Tx8Nwe2IwDL
iQhwA/t+jIs7/Gw7w3lqmwtW5Sx4jr2f95vGu8B6V/9D6se0aEyP6AFh1O/kEzR8
Z2GRMZ5CIXXYSiyNgAsn1tBe9PBAGVnhPMk7UJMDd8GgfcLXNmt0y5IT3DeGZ9om
oV4wke35X9r3/BcZoKdto0ErMRwbq2/s2wKxrAH9QWTtnsZ8nUfXG8fdQq7e3F5h
KdB3NTuJuklj3sicy0SQcXfQVaefaq1kkQcL8i3e4umODvOOKZEHCU64ek78MOzn
VxpGWwS25hsDDAQDzRoEAjx/Tbtp02TWuPjFSAoozL+Y3keF1MjxlO5gNwkzUtHZ
7+4eI+M9jdwAot3shtdT41WqWGf6fjmG03nlVpk1cujcWas7idHlXshb8AaFjlFE
SMqFvpLm40zY/8N4BAQIQyRF/2TBiMxtyesYItWMm2kKeTvXqUSlW2e8po4P4X/r
/ri3r+rvbIWa18+BRWrayhooKk59YtiLj5X3Yp9RhmCc3edJiBHmQbE5Flqco8LW
xlAxxwsbNemrEIomjYnoXn4smkpF3Z4gurYQMvRih+x1Ax/WttDBExhJGXcPy4+7
FCebshMfdH3gTmMsnE6P5J6qGJ8AakvTeshPhUtvUCmtaM+BcsmKdZI6c9e08OLQ
ssQXIF8F36/K9mU28fgJ10OAYAspTpBoAcU2W3oF3iqS/phGnRlGgxV1lW3yJuLk
pfGgCdCUV/x1cxn4aL4CL4ZqakH6JZwQtaFrMSVpBdearg7/Eo6ndKgEUEKrRQvK
/EX7KuBDUdFNda3ty4+sUgTfNc7J/VgML4ioDU7jgN/CrYuBVEhTMGY9k3ZdkMfN
CLXMVMqymc3quTRGAQul7gH3cF761slGweO0c61ssw8+mfmvDHRdi3zX+vtGvAQy
HRwxUJilmdvZswXsAi0xpJV06lrTLafp3wuc3JqHRQdKYIaVzloo1AJjG1G6Lqn5
JVKx1ODsfvieCDzYZn+vbyQ+Avw42tg9A7OLbL0EzGuEeRg38fJqtBeG6ccqvt36
KlvxA1NWiwKzCrmrK1Muk8NwFaG9hmhpYPNq/OIKeUZGlwm9+aQGhU56Ioy+miQU
O+sI1Xahivh3cXAo46IGgsVi4BKJaBVPbNHFJWcf6Ni8mhwvRm4n4RzsmKg2Mo+i
llEdQ5xTo9rgc87XrtlExbcc8WTVgKWqFSgTJzwlePqkoCP3Giv2dB7hfGsHJFRo
/YFsVqtQ5U2FDVpRhXE6lzxAlRVpG0exfXxlk7tZi8And6W0eSYLMRKJ/KXQc4Y9
gWQ+ryt4RJjnO+m2/EhmE8w7Q0lZqLKtlTTphPMp+77LDAgbX/oiAC4lFG9MnYOc
fndgO9tazsspWSx7zfNb8lZp153+Pb3EVhtwnZfFpdvPImElD/kGCT+wEyH5Licu
nRLpH5MoKdo049g8trWPFu0dabQytESqWqMikMsIHVfIB4ZxWv1poea0PvU1gB6y
yECWz3W5+UikRgJRZdT6J+U5TWi1h5CnmgnZ9GGLjapDYSK+AVYge49wbN7xc2SV
y4NCJgfcpj35YWb2XDe1LyLGL7KT5GpESPuXqOQg3FYst1FZRMx/KxeSaFB6gwiG
yRKH60JXGFXwNiO3ox9UbEQbVseAr5DGiWY7nRvz72UyYoAgvmgarlA2FBzgzJ8n
1kxhDgIpY0g4IlelwMUKmzCRUfUahn6XHcPHL8RdJqHVwIJlRnhIu0bdNvsElebm
NgMLgDS0OFw1NJYwIm5qLJ3VJ6/38XOlECiqs8ODjKbZg7tl7w9kAMFXfCAFVAsZ
I/atw4lrQmsBeU1YAPAhxQ2dfxlCde1lyEuvk+vUaz2WFf/hVOh9nzV81lwswx5B
DmljW2/4aD2Aoc+Tx7XcoWOSRNm+4zObufnQ5wN6xN90UF3UCt78mkWZqgaiGWst
mFgwo8cXWNkc/oAGJrBE8f+lnbRG+NITzfknzxYwZvhg91N/AgrC75Ycv216a1s4
TC2oG1rkTCCoZx+cMPId/cbhJhiewMIT5WrLwn7mC8KmrHhKLxoyHpUybbmrWDRd
IkjoAKjCz906VD6QgSVCSQfwsBrSdo3FeMSuuf1feFHiCPE2cVSa6CwAH6NNjkqQ
mtDPaAF5Znn7oS4/6eMDWaB/UunPb1u6YO1Wma9jQ5WHqJ7SPhSZ2yqrnGXAk934
aQiFxwtRkrDk4DSzWq7i0fvnqBSzkZpLmbCTVMUtBOTbI3XjMTE7wGIzLnc5hXDe
6WjJ4ts4VmfEAKUvLnKevlsEs/rOtOytJt6C82BUx2P0CLhznNqvRsslkIXlRemp
xzqNtY0jcb78EKQff0GyYPDgfoOPKYVchaC9cJs2b9auw2UFeCpAuwuqUlY8RYl/
f8yNh6VAFHX0oqKcslbAd+y4rBT+ZaqlAyKzDE0uVtlwBG8RJqZ/IjFkCd4yzyrF
mhXd+1H9YI4XwPip9HE/pSgiAwGpwU+dIo02cfPQeIdQZYp+jFcwWvTNGK4cGKOI
nLTs0FwMZgIQesgJUHbbFQdLLmyX4eJGScrEokkSRChr/JDLwwW8YZdfIWqC5jM4
8mfGJ9CbHcDxV9U1PrhMIm/Ehc1fKC4xzp1MLYJhOdlpDljEeIevQ08QeL3GJjP6
BXm48NZV9NH6PciWA6aeJOhfqE3Qek3iaKgJXhvuXtTom2nDjYQJOyBYnzR1B7Hg
Jcv+SrEzymOaJnLqqBMzQc0wLKCWbU62Z0SS2a8zF0dsS5GrZWKkrvDpjNWAufEG
8rsn9BgJYckJntFVa1lTHTbH3bGl2u9HiimvlPMOko2av/euhYkOlzDTfmuiHMUp
f6COmVJfLXdZbF/5cpUzk6urxCoTuqvUs7pXqI385XSCDQQRSfZxwMGv/t31iLN7
rzZMoh4QFOFT29Z447sPBA9lornSiskf9NOzQDuJLtq1zslG7gtPJdFCJ18+1Qem
SsTtXT3mP5dTeApG45Isjhksum/9DsKP/4KpN6WJQAFNZz2yMtlmacUd7BA8CMiT
FU648/tfZ2uRQTzUYZRIWQDG6UUnnXCQHYdULplP8Mztu/9jbNEA9c2kE825gWZ4
h8+O3gYKKZ09KZpH0vQa2230DXmeqZkU+adA0p2OQsd0PALDo0hfb860Ob03GQDW
MxgcL5tcGUQgctBlRPfpvXqzhIUS+zuJ11Omrlseq5AaOpTO7e3g888GvSoM2VYe
S4McS5CWBpDqlSScTSCFQtyrKPa5cHpFqANINITw0pm/aMbvUR/1uCvGtq9oH4dK
10+jS2satUlUo8g0Vt+/pjIgez5DdiukQcFXKySBVKiHPMd4Er6J5Fr0Bn+urSHz
8w0E6Gy7QL7o99Tp3YbzINIeHDIn4/r0ORdGa68d+XLjgS3VJY9Ia6L/WhrVZTZi
j6R7PHfCh8u4fXo0+E5qvKwpsQA7eChjIxtWmSg08B5KAQ/jPItLAg9p0nvkTisU
SHLJmUxQ91mfGiQmTYG1gIvScGJq+UUQ+IqmNCY3vl6AmopzJR8m91T9QD41LVT2
SRsEOu7FpMLjGjs1tyNdACmtht2QrQdnRTmqYGxPDjtitfEHXn8Ut+MRxgJu1weB
nkrl/NRUqHpGDDF8HO+D9KZtFEk1E+IfR0/VsB/cDYfeTg/livwE+R7Yf1jjgsdM
fV0ePyZtdPYADH+DZONQ8y4TtQCaVTlZTZ4OR/H4E/jNt0g0jan1EUdWQ0K124U1
3LnQEY8Ct8bJh5eL1pKPDupQwoaDYMhSsTD+ukKv4B22pwqeJByn4b8m0suQugM/
eY06WFvjXb/YMY+MT/Dr5k9fxe22RcpPz0dqPkrA2UXihCc/kzZPjG+8NqHKRba7
0Q2qE7SAEWZmJm0mz05JqjczCp01M4M+CKanL/wkpiSLNfGYpQ2mRYQncODf6KoB
CQf1JDJ9MLdUIsjP/wUy0hZ3iYlzNkxulxxuqSM9kZtNhXDUaNVlZWy5Me0XTCDl
koEfJErDM7BT52TNHyn+LvymEIU2fE2aMrzwdtKeQI2+o/tPzhzz+AcyDlygw8Ds
XiXwtVRdvZZ6xctR6jKpgtzuWVnpDp8PYt+vImsaNofO2vjkfA/JHd6y4Mgmmfrh
6XtdS5uwKluhKANXfEeEnMXnPm81P6lctm35sRgMzZ0c03Ktm2+BwyewnoeKhrG7
Rg2V2C34In84y8/Q+/aCIRV+LiiA7FvT/u8QblG+ped2/Q40lnlBHDts9PcAbwT0
slghnZFrN4LgpGitEwoHC5VaRWaH9tC9e8sdm2LNx4luc0wgCux6p9Ra11X0lsWN
SfOW6wBi11nOm/2Uvgx916dx75U5okUULkyX5miOzxA9OwCH5DXaEY+MHB9wT6zI
VTy11rZ0UV3tFZZP1WJxjzHtWaBRECCB9HLX2/tqt3+eDC1bCNH2UKGHOm5SxjSe
O8hL7o4Pc4Farbhgo77Wc5TSDfMBRFVwxM6lYfgze/rDaaYkYHZRF+jMUfOzIJnS
cfD63M9GFuLOX0G9DsHUEyWbxbOmAO0ubkiuLPjf8f3vDSnoPGMgtfokSwcdXkAb
h7OddIbC3BLBL+0aYLTNpB14CQUoeCSzhcyg++cUrwLxkkizcvD8KA/7EN2/euKS
P0NfRcTiHYN5hO5EP5Fi3RzKxTcG79kFf3bAQur4oGXRL5FjHPXj+RSaFZ4vk2kE
VhcnDWirWpmhj3582TYeNySL62khi66j8BxjieUkSBKNbYObZp81ceqZ7N6qs7jq
5mo72czbJ8IVLpkEaA5s6dqEhLt6wy289oNI242FVHpL2yP2wpyi1aPRVg9zzqRc
aDJBaoadRvfFWANqUsaS1nXZrQUjiFRckgganm0DVANwq3P4JZ4DYEyyXGtSDoM3
oF40280Ac/4UAXYlpIdr/mL8PhENxRD9P8Zw/mV7w2Ol1wNz0KE6GbdguWuV5GqS
nGLatFiA2J2y0DPMlL+PN+ciJvs+ae4tjBvS9af5maay4H52FcVixiM90N3WMGc1
z9BO1MF2EdekBKyQiGfwmdhEOEVKyyWqgAjyjPbsrMsNqQHoDBnCi/kbXWFzIcJ0
SZuwZYFzcha27JToGGDB2E+HlZsikJ+CVDqc6wnuezwrdPIlB+GEAc8iKqiEP9dz
FDdrvwTCwV67FRMGcQkXiXF109I496S3sCI8CCKJIn7n5riIi2NqUtENpwJrxAH2
BuCwo64FVQxQYTreGWmTrjjhZZshvTKc3xqgKj1cfQ9lw8UjXCzFidVA+vI48K9Q
9qnp66+3RCXzrkMIOASGfpOmKHtmN7EZdrS1T8n6OEQPozKdnXL3iCT96Q2NGTZg
zb/E/zA4q6M1ZoIyK+f3OYznMt2K/0I7Stoez39sZmjTN7O+hV0mM0CYpd7Exom+
5TJp97WCDghn/pa+E1QtZ99Zmf04DxCn7xk46TKBjZZzpbqpeDeuR6XPr020TgE/
SVN6UbXdSXKZIPj8vasqpEgaY5CytyNbSE5xr+EoqHLtAPnVnllHgS0sr5uRnUCj
AArZn+WVNvDJ4wwOflsRAOdnHE9p4WCrZKrbkti0K3MCgp7xk3aTuEsuVn9RkLOS
hDNsmpyk2V3xRmTRf7ScTilncihvf6eED7knqDzVTwoT8h5elNbA6oabuq6kCDxm
tsSsnfUZuMUe1XEB7ovnwmAHWtCESVo81gf+QIqEPjPRO7n4tlT85EssZVDngXMY
q6MlAom6Gg9HPzhWLAO7a+dy5Rk58ayU6kroX+kuGsTeIbHsd9f5NTVM5VzDeg/t
LuI18LFRh2EFhOrQ8iLRo4HW1T9JiXp+T4JE0VVp+arCtx3JmRGlD3zps+WL11aL
5eHglnnqfUgy/3wAxobNSY1vnMqeOEmO/614ufeAsgRkccveZnHiNd4TPKFbfpB2
jLoK+d3+wkZxGMKbWAat2H1r5T3V5KPuSsgsmCOPN4B/yUPmfkrQg/woFqrpDGWA
LbKYYZk1/VvJMfYYIXiMh9su0Eote/ae7QA1gJrTwUm6CXZXVpc7dM5DJ0cm41Os
N5gOhXk1Y9eciZHZKQJnUZT9FKhWHnPtNn2Oq0sMyQMeKh1FohZ+tjLXfqjVctUG
SQ3WCR58CmtAn9uq2JnclOI22+6XuYpSnY3c6/6Eqwnw5yax2JNydxnwE2JgG4p5
mMaFCJ4CwhDU5Eiao3TM8ASCe04lACy0Dbly4qIMIC7T5dSlzUYrlu8bye95E1Ep
QIUhF8+7VZJ0hyjYmxG8n6WkLyEQPnM92PWqu5dkzUOVrOBumdJehU/X69gV09lo
nEdbm3g3YY6tWa2HgUwk8Hw4IBshi9xp65qlp3xvdKmAQhTB2A1mFT6I2ATgW0ze
y5IeLmTkB3XilG3d57exDbKc7CFU53L0QOM1aTGlZAnvdUnO619/rP6vjHO2PqD2
iubvDxwiPlc4Ja7tyCvsD9YI+GHiSmgQ932NmGv9t+vObnmKD9pIZa/KbE6y9qL7
Kcc8sGIgWTDdx2IM3ZLHss+vgdxql4nWUYEKJKrFXkhTu9DguMf2Bmzt7sHlIs5U
Rn6I/zXD2ddAosQNr0bCZhH72/VENxIY5dYcOwf7vDHGLjRZWY1iidGf9XvXL05H
HgTIYRtqj3faKd6qJ100Vg8uHdVkTO5b5v5zOcwuxt2VOKBkwMSm2HH5iUi4yUFV
xBRgVFa/plQ/AXFjv7Df8R79T3BzoGFJN55M71rvNZrU05SHPiZy1vebDlJulkXX
p6UPWLY3EtI9WQzQzQRkg7sH/CJuvBoVdJ21xy1BVmpp1jr5eHLQhBy8fjYCOzO4
3UdEdOqQtTFmBfpH7jQ1y0FjDPh6DrJbuh67oeVS8LJIeZpwgr1osdtITt0Zsspg
pvZocD9xHI3k9hl40goNwp3Xc37jnHadaPSEBwJwrmKuQeDb0BS4l1TqR8YNQ6t0
CrH0MvAbPIvTrxRkO/DmjkEXtfnjz1oUEtqIXICoc87s3SgmgwgbnkglWwpwD0Gr
Iel3KdRs0esAU0JJfMJPCJv2Ge6IB1zYU8dZeLnLrkaLhwEl7fjXq2hADHK5HfRd
r90zI5nZ+g5NwvfdFZ71yiLHl4fPuNCdReHZFtrXcqk/2Ypi7mXhFU+8WBlmOR/5
dPfYWL33/vwKopp5wb2ieJ8WiEvWFkBcfS8nN6KbfGiDKYAZSkIAmZek0oIgemL7
2f2a7b6oBvKGQJjl0YDcN0agprpnIVy6go9o4CyY0RZ6afw+I3thkMY9p3FjpgHl
8auCHkUx+MLg2gP9W0qdF/VCeOJSqkIL3obRop/yYHxexkKvWxSn4j9+/Fh8W68U
WL14EnoI2BfCC/vnJ70FycEeSQDM3nkzO0wmNp4VSlw2iDM4F7DQnieFQDRvaG7k
sAtYMOGvmzcHMxsksw8qctl/7pTka8xbEoOYRv5vfH5LQK9bu2/UKtMNA0bW3adq
WbRdx5eRIqsUCz4MYl2DQ3sh2YIl6PRLwu+j/2M6H0jJek2CVpZwHYUTUM6LcEhd
WIN1sb+0eHL2mu08n50MiLUUggjZGJoWfMI875zat3okYVlRCJkgNr49QZ3nNZGX
skr7UIHRmLUOJjt+vfAgFjaJtHobfn0WKsnQy1mkVidvEnaFeyn0l7Tzd/npfYbQ
xeWonH6sz+WNOb+vj3eQ0jHtZ6VJoU8nvkfhuIT+FKfIHt3qnGqVHFVc2pJ0X4eO
9YQIyWFw+Q5afQm9ichMQxkN86KqbNNcEan2sajN74AHLP9U8tzoHUtC6niQnj78
NCmtsXcQYN2H2+ywGpZlXSRlXZkqM4MlaOnHISMusAzOGiW9OPZpO7Sv+E0VKLaw
Lv0jkyK57pwS2CnVirznzu4yizImshBiqtmfLAXz46YE2QTDZN41tgWFg9jjPmCs
NsiWFaOPzXYgYEtzx8WZUARHmy5T5qoAgPMKYS7o39O9R7uwWphX05QfQUPRzcbF
Fw7veWLXBybP/g3zwnXf02SnLAYDVbHfDAHbEh77lRf9qO4hU9x7MuHncLbfStcN
4GrKKhu+/1p5XUGG0ifDeWqHT21UNCs0ERqPdRED2P//60EIJJndZbkEVsYYH/Ac
ENehQD+cLhePONuplvUQKuBqNwk7BUXAc7u6U7vu6OnBkLXn9H+JGYRQiYjEw48d
bhCpvxQD67+Xs9DT+u8mskJFT3QUOIo1gDiolxwx0enDb3jMMCCsD7LhgHgO1DQw
dhk7NpEWCSIAkonAM/+ldwIJgeH9oGx3nlemSEWpoJAnZrTbQM7hDC5nr+LwN2kk
UtVUFb2wTUH74GMay8HTxvY/Me+AzuFexLV5qcoRJkYTyYEFk/0lmwiZnCzy/6cv
ZTo+zr+JzQGc7wBdEIf95iQTFP5mZUuHi7KGHz7JqTGaN9M1UKwZhwSe3BizEpJs
gw3vNrZ7HrLwATv5OzJvE3NcKv9odrgg24Cni2QRW7d0GM8k78cnSEyiRFUUY1JK
zAMV9I9NG7+8D+9qTdeob/btvI8JN1miGVb1ZGGj8nGAbk9+Ls/qC6MioY8OYv/b
guGqagHHURf5xI69J4LEs8n3ISV5lAyH7mz6Q2wm5PSDHyMjuhmoI2hf+KhcLv+E
8Ytl9vDWo7MjvC845YBIHsr9FWsHlvGHDd04u7ii4qIxX+tpKXsNvIcMzjkNzXu7
byjhMZgyTXuVWx3mNkMmea54YCiRD5J0qzEJ1QdbiVA7IrXfFqVjc0OWPK8srxuW
qrM2JzYJa8gLDfP/dke03ItsK2APCR23jOmf0LVjQJGBuqnbxDd3SFKYjwseJ9Dz
VCb+cF48d9Q3N9AhOYxtsIz5E0jIQk5T2ajZte4yL2G0bWj9e7EUR+4bAS4hwRlJ
rYjideDzqohj4F114lefNETYPQar6uMqo9ix23hRGbbKzdllUyvwin9MlPIB9sXz
PFZb9ci0Ixp9CkoedjICbd05fuyAiNbFEJgwcvJ37JrDWcEjhBZ37lGRl1whl8yw
jfoEd6Jv6KYmCkudCJc+BSt5kCSAa8V4PwZLNICkhMG9NNFb7vUruE4twUKT2p3O
aorKuom2yCcXQeQXp6Ht6pEfnjPEewbDZJSkUPZYlgIkjBpk9K1YeFSYNjAzBrbK
AE46ai7wAmrtNEw0rBrB9NGfSHuAfHkIzyYqyf74VGXViENgWQ7UFKqathSQwUS/
cX6vrcgLipxoYxCjEOm1z5ZsZyv/dEVmDFG3+8h2oADaKwmlrWt5hU5U5GBWeLvB
H0kQ9qD02FaQD9NnBRIDQ76ozhn2oMV1UpdDJIawr4bJS9j5A+5npLO7pRH6HdI4
pIGaUM55yQbK/S4sH/qg6lLzPu3VYlaNSVTbdaJp92bJx5kJfOKtHLIiUWA3wgmH
8iPRHwKfprUOFeF/sigSueJGj6GOpXOWJhIwLECjr/jQ8euBQR2V9fta+qtZ1Sn4
3c2weId9makEuIuS4aYSfhmCgRVgAJoAO5K79YKmihWqkj0j6yMbpDp1za0KY4gk
Xm8AlGLErNQyzuf2ufLPm16VEsgEy0p2OHNWSdUBGfdQ4tTLs2jvStjGNjPNg5iv
cFJi4wcvex4o9jzZZlYtXpcJpiiJrf1nafRIHPnKaEr3eKV3Gl/Cb7e55822d90e
FR6HRqcSHF63qlKPCRMrb91e/T4mUlQc7WtbXTP+0kKkIwDvNuzaQ4XV7Eb7xZAQ
oEHjYz96SLbugEOUO3AHXE/G65DnQzirVb16g2qKMzb0uh3SV4fZPCyo/MEQnvMM
L7Cb673gLSPRosZZVeV6gVAD1u1d1WoTWnkTcqYsWxDT7CFnFLmpZDMtPBiz0F0d
G26cPTAtwgcsmM0n1m9igpBpj4KMjX/DpP8YYfgYUOcAbHIsELtdXn+GPeYLeGh8
nEW5HovhTYpklVFjv43jpXs9OLJzMt3ubfS5M+0DBpyKO9g4nWXThSlm2n5cBrhX
utPS2plyAvijoKcHbeZcFhV8OxzxaStyXF2j3uMSxkVS3wDspRS9wCpeMrscV+H4
+NLz6m3oPy6+sNyHNg2ZY933ajGsXEPACIjzuAF44tmJaKoqDTvalF64DmOjZkgw
NkHlU1sZrhszBjbDq+KIPWjvWw1E6cwfrsNgM7GDZVHDLruqwimrMLnY11zl/CP7
cRllJ1Ita+JLqo53aHpbZZNJ6a7HQ0e2hIr31138IyT52CiqsV/+IOrEexqtLG0s
PsbWc+L/CA91a8G9PrU6+vU32TCLXQNeyTgOYUu4QfNcSXZi5XDGsFMjfmEdCOPu
rlvCh6UH4hKyRCBUckD8pvq8NNyZsi5ft35miOzcv6hsFCoGkSwr0j77zA5xMCTn
CwEx5vGhRkeoiMu+hEZ6ckIL8ce+WI6crwbf6X2dmDbOIp5sCrtBSyoicIIJTyml
dJMU5+UjIYCBNxeLmss9Ji9t5CwGPB+PmDcAtue7xGWG5mPA51K0NXLxCXteIQph
+pcLgnKUseJPbkp5AznDtGBPd3lqQ07HpQmSFNRYlMAh7xMAjcFSTAtyGIeuSx5j
hOIWVTP11H8beNJYS4Ogiy7XDa3V3rcrBZaURSjdddG1JXnR16ARIEgkIa30nlsh
bIhu0n/fW1rvNitSrPVMkguBCUuUS5vMDfAWbJCdLrXhwl7Ssu9j1zx7UTqGDowy
q7erNcZK7nTyexnRyA0T03z38fr9Gysr910h3hFTn7h31eiOfOpjQZO1dzM81Rsb
pg11wWJZJdQsk7GFWYcjPb5sIf9tbRR51b4uwB2m7Qh+1F0l0WgJwTHyqUGfWd5c
heGhkOrgWZCFqNwAALVMP9ZQ06+s+coYjWUU98sefzzC+D7zVTrwmcTA3BUfxwDA
jSRRhsr4fql86ig/wz2eb/UA+Is9qIhi4A6ZLaHxz1PkaeEgvTdpGuduevEERHwq
lgh9EqOcBRAoi2gk7VdOFmLMyYlumjGg+LVMl8S7VUtaeM932nDRXz8ix9HrFqnv
D9OKIUVTZCzp5M89rgOlzn4wr4au+lV06uXRiOcvUq2WrHrZSUuVhd06NREyuv6/
44MWUVWqir12ArxceSxihdjGg0+EGAHoBKA10goKl7nVDikOmHw0TcNj1AzA1z+e
R56ndOmcZ2pq+EmvM9pA5KfUywXajXDB+7XVfao+txqtbmuaROrkTAnPRrX6xnPe
3DD31NKQKYU2wRVYViLCeIsOqdhlCj0d5XGicoIom4Ww4//f0e9a59wGSTS9e6p2
z5ohhtS8xGoELopvkTfRtLLi2EvRO1g9PDxEZRSrMJmKhi4ET4CM7/aZkW/C6Khz
zNetOuk+VdXD6yIT++60pO4SlUmM5eWUwkNtMsM1eFsZ/pCKNGDY8hyxOXNv2Jcz
hnaVADzgt98BDAC51xg+wAoLOtOMhK2eZAtmitExKBQxw1PaI9NVKwiyogrXVgTg
XtKNagG8Xr6RW8iqGUWdIP7pYTysQXwQ3BpXvnGr6pFuowWFJN8Ljjd0JH6jqQCw
1aZORpB0GMbgmQgclK3nnTxQPIezURj/fhzDyJ3C6oiaPO9rpxfe+cp1u8Qnlsy3
2aJETY+cKR7ihY1n2n8XlcRyzHffBkrKphHIo53GK4B51ZGKIJU4jNSD5y+o3Up8
0WMWdkXq0JkRNwLJuVSi9ahw3AzT9rw7PyJ1WO/+cH8lGVNOEQIjQpbePWl3biy2
a1t/NZ+H9ACLvrzvVxhWHmp49mtCO83zKNOhPb3tV7rqIrgMXu3aOi1zfWWVXdfn
RJd2O3bEEgeH+CEWSoeQVArQruzD0DCmRBSAhOHjVh+J7WapAEAlOsLESH6ADJMI
b34/q630Jz8EuJUnMLzxLLMLTdRJzHAGawXLR1yocE2IXx/oK4m9u3UM9GKrsrRA
3NECL7NYcTaS2+u578Slnkblor5AU7fmZiMy+jKoC2SPYCfJRoxEC8QYsNkeS2yh
3cYBmOFfQvapcs6Byu0bzM7HoBhYbeqV6RwVrNIF/VITsPFQu6z+4sTka3kULYrh
5pRBo+9AZ5ioLLTxFgj9qqepmbT26aiZbC161DBQBju5pkO0PMhR2shZfAxv4w1H
aWQZiGUBKW9V3zQp5gKqJN688dqP+aRJiv0WdqdJbFacs35ZsptqOKz75w2nvN1q
MTN4VYQ0GabFGz/Sv7EdVM3ZDfTWNhbJO3lpXmwxxDyZOrdxSlkWBuoL5hf5RMV9
zeaFQXLIY/M604VW+KPzqrkKNSazI/quHNSynmEWIGZwEJ7hKhQbiWBtWZ2kg0Gu
GIjCcRkZAO8ibxG58Mp3q8ozOwl8FOaq69moKgjs1j8t9yoBKEr2krQKutbdsOts
IqCsUnVYRbHjmjVshDl+vLEVeg+OGDfxQG2ZYxE6AIJTeTlMF1pmT9UdP4V+h11u
fEwdYyddOluVQGSXVmKa5IXghg91pdmsgvijSvsEsIgfmqtGJaUXwJt3dKLfS53+
CW6DmG9cCXrLVirOhklaKuzKVw7EYxLRj70MnnRVs6Aq4uSQkB19nAuBJXn0E+NZ
GpSIpsHry2EGT8w1PIsRqsXgNMLhWW0FMD/ygwliTKFl3SCy7T4J4gu1E64Sn0S7
35h75jdRNgDp5+Fnx9cijQJlqrrmgcD0xDcvlKncEV2U66P4OoXtfEwl0uFyqxW+
Fu8OIeCQIcobH1KsDBig8AXkdM0oasI+cdkDmx62YJrhbkIbAt7zYBwX9/rb/s4g
nrMXgkJz63pN9C94ab/LZEN8hzK1HaCuLZmtB90e4p/zNyiOtPJLj9aF9EE+hGMU
q1N46UZiBFggDnM9ZK+0tDHBmN9DcMfiNZJezUe+0aoaxBHd6ws2P/IetTLQ64MJ
qQrZjb8lN0PHlZ0OtSzHR0Sp1FHKDfwI1wD3Am44XX8fF/kCccW045jK94teIXYa
pPyIJRLVpt4CP1Yo2sDhLssYHSRHuLzIomIvUkiN+EJ2Cv615l5QcLEIhorMftnY
VwHW2X3hJbBMatdSiNVtg115SIboDAZeRdIQhDLhTn7esFhyMra9tK064Hr7Nb13
/5DEnNdtkCXnPr2oK483NYedesjegEGBRtL5WZgJHmRj61bOJZwcQ191+CGtMQoL
0SGRaU/P4gBWhbZggbaFl7Y5l+/aTv+1+t5TcIE2X/33ASv8IJgOdPdjUXpx/8S2
5jylxwgq5jozNVyptogbHgHQSP60jw9aMHVp87AXaY7Wl5OLWa6go+EHiI+PlUAm
n6H2dWP1KDcUT5l1vFQeaMjT5IhhljH6VIHW0GTSdsn5SZZZbMCFK4dcKd4jAfoq
hOZ+4v80mWEJc/VBZvLdfNvcg11MuOLl1BMEx0xWrQmd+onr+y6XI7VyZDe4c6lK
eO0d7uOuAYQAGM5zzCt3pVhGWmIbFOuBogMgcQK9Ffa3D/1JeuUwVsJzxwj+YPFK
dZAqh3gRXcNF5VqUffF46gi66fNEDiXNJOA6J5HiN0d9yT73lFPIwga2hhdB+8vr
NbknmRg5bK9360OSXrpuh0JO4UQgTnIS6S0Adjgcak4lMfGcxoswb5RrE/5akizU
DrrXznluXvwQZcaC4C49jL7YqwpcmXRNx+mDLS1eF4c/fzg9h+dr36J+oEFOJntq
0GL2IcH5ToqXUjj012DMXeKlJQiGrrsmDjGTEgMJh9C326VgOQDDbGvYz+/oLmN0
R+CmiumG7WuDTyu+NvzXJt09UcGrdKrAdOOq6Iy3hmlLHeMtES7lExyGaGNV/jhn
A7TS7owj5DmOktq559/7eXfIobKG5S+U4hUCq4T1JH6AosIMdAfA3BP5pgDkxU69
xYL3WZwemR5k0VCEFnXDgGHW4JBvtxxdkYNmgPMXEeg9bzDmEwXfcePFXNBPM2Fw
pdnsbfwBH8ZGXgJO3K2F8jAJnmI4JKdFqwywApdhWtYsINW6k76y3MXNOPzJyDoV
HS0tuZLCVUPXElgOOT8+lwfZ+czxTMmdm9JXSvvnIfnVlavhBSDcD/pQZnfB+sKf
kLLk2dWHtyho2nZp9wk7vLr+SPKPRujFlDDq0sSJFz5xohQp/orfK5KY/mOlh8dD
7Se0kUOcG+07UMhH1HmrPZe6woq1Ad/m1zyrPUl4R5BXItSCQdMfdqYvnp7TP/0i
XpZWOFse9To6OM08CL3U+eb6slBpwCoDwl2UMnud9yJt0GhP6e4+RKtG9HaT1vyT
GQWtAk4cFJGxVzWG9F662eBahTlEH7CXfoJ+9hBCCPWXX9sagqc2qKb6A7lrU0bn
96b1BeTzzsBjTowRw6EuMGpGdqDoAKNBZCmTLBHPdeG4O4eSBV+SKZiW8fvomokL
N61Lq0/8jUTu8/OPg51GLeQarMVR+lBD5JIIIn9hA/Q4osFJfcxaSlbVFtr54sW4
YQeRhsvB6E843zdjPN6GMieYC0KXhk+tDbwMq2rdMtLtFk5tzSAg7BMbX+k8l6ON
pkbIpnilBrEP/9GS0zc3RSYOqr+tL2MbjLUOOxhGfc3bvK2pJz8EB8vqaHa4/mkd
tfMhMKEkxHnZYUEKLZufDmbeWl+vcp/jeb3NlCaxtCr6w6XKjK+8TbAdlcqrz1cD
Y8ZCh06PxhoMztUI/JsNG7zGaDDip84xy0D6H/7CzBNII3p0x0WHjdSLFKJpWOdf
Mhfd3W49a1UsPC4yCZfnnj0SmpVLLBzpuQH3AkFyS8ObvzUWfnM8HGCNT/ocZAXW
lQGTZ/ZbSu7CxSrjn6eMoPxeeBLPBEagGjELW0kb14ZtkwRDg3cTO2D3/kflnRWI
FiscOpm6+CyT6kDG1f9tvVHfYYuELECVze71WXmtOkXegCpdNLdp/+SLuJZcrq7Q
AnDwzSk1hLjn4WLMAk18N0oKeVHsK8AKvTOhn1YJbqC76s+FMVn5gFOeDPux3tZK
V0WGknN2VCjDOL7HkfVcIScHDaKGbVx3ph04wPLL/r4RfPhY84dzru31HcWUtBf0
b8BYWDaduIeuNeus+e9cSS2PJ0nRUiihYxyyRSmRGkpYR1W2CNHF6E+xqAmlVA0M
mXDkFGWILr8UiRPl7RVDdbSehLbmVomzmZGoYRXxhdtOxI48Gtz07HEtdfL4eHEd
EVCvXctFO0znecfBSUaTOaBxPGrxkudAgLEvUw1F+ouvWTTwGvO2y6F8uGoLDJEu
na/Ctd+LQkJNtQIMP1r3PnW9QdxHjc2ePdoLoT16BV9zsVQpGPBn5fy4D+jVrPW1
iOVqYMI2AOpmP1fWfoyvoYCvXdLj5AibdEcwqnzB0EHnKDUdV9+zHXHAWeoQVQbf
HfpEOyLVatr+T4mKH6UiTRnnt40Q4SHa7ylOU0n9OwqW8IiTIVCHbf26YZs8lx3l
Ga1RGpBbgYsrw/LTBQMv4hvqHeGZeq0ejQ99AYY3KwTwGJBM+5e7dQiDrI9GQmEG
kWGjCc0kwK3ou108Yu4vQL+gifAROMCreRoYRtxDBUer4M0XHoIfQjwO8CfooYiL
idWIqXDvlM35HKT2TRoGmWafevr+BxLDi3vRdo3qr5ZfzGCJ5LGz/rhDK75GU2Tj
vkZXnjDBkZnpT3yHqYnQNxyQ0E1gSgu7AMl1I/qfgVPFZG7JcXqXf2YSesgdiFx8
i8c9rXdhQprCGUQNjKjFOKQKSxH0NLkL8trDNiGAZFXI8dCa4xGHEeFhmhu/Pi+G
EdFgdFT8cydrjJtbnlg/AGt9/BCtpy4KBwOtMAcXPtpRB4BXR/yX0ocizzyPskNJ
gRP3e3sH3mQdnXFJMwCxpOExNY/reDQqXNbzt070ZvqOV+XLzrooHWBpUe4igOY1
w3d3rNBXSPfx3TIXq5shykP/OgzwQd+xSmLQWHPGOSak7qTffptq3D2HqEpqc0IT
bWaMXiWOlApug1aC6TAl4QRBD059UUNWe57Njk97RPLD19sRSMh+6SrDbAe/WPhN
634DdH6MvCK2eWPlqAjVx89AhgvZ7CC4Zhcku+i8n4pU8JyuxvqD4tgOACv7nxyF
MOfIkNjNBNLsJlPYmKQ3WRg3u/CDhHf3wTY2uOBeXxk5j4HBMFqxflpKtS27zPpk
mwOUZ40kSQwCNzChBRBHHXiJXcAo68oqbGPhhIQWBVCkTBhRJ3xKKju41ZMkezIP
VHWsz5HWJgUul/frMlb2dRc2Rgfy45v5f7/MmAToNTaufiv/LtcEdXipw1TvjhbN
1bqm68fZZA3Y7zcDulG55XJAfMZlqU4frx9yupTIQNlOljGGp8uUlF6kwgMM3UwY
ogB/UIx6/W3dqGCQ9y5JTO2gTHjLTgCtunYx9Z8Zk4R+fCy+SWhwNwU8pygV57Y1
ibgTQ6MIR5jh7t1oxxAm6x/na4+Rbt9AW5G5BbPb9EcdoG4GMfaC7JpBnp7rDg4M
aXEV8clTsFdiJHWLjf4eQP4b8orR0wRgJ24QZL71vWSVNl4aU2MtgYWCpbZUhUR0
kPNxUIPOWlIzm0PxiavhAdyFD7K6zsvgspfUzhLC4RzMqU0Y2EzElmf0YmP5bbdB
JoKmVGZQMEg5yMnWsJPQfHMfMeqURy36BiMiTDQ9Nl2q+hK0KFxeirpllIyu7Ooo
1zeWSObAO/9LCw/zrQ9ce/ubvssXczYDZJUBkTu06WVSLKgxT1w6E6mENxLf6vlX
XyCRGhmSrXsQTqnV7d2Ur1qSuZN3u8WLf7LmXjvNnXzEC7mRtLfxQYjmnSslVFcd
UkIfaT9stUMH5c+UqO/lIYW/3dUa4VGKvnFXWcrYjTbzNubNEROyinx/Q2w8BFaE
agnrrk4mOuy0B/++enhXMsdEkXRXaKSY7BzmOoqpbshty8fnZbnEbPybTGMiADnL
E7wxa/ZqX+HfDHOnemKyl/Q74UBwpE3XCcA8dW8UmGz9NR3bo5V2uoBibtgXz6Yh
fDEvi6Ydy/Y8v0GqQ1Ir/VBffHYHhIgO6H4Qaj1T7HYq0BD34eGMSbDfHR99kz0t
H857fD6Brr7esmlhj8E9U9jIQcdPXAKWLO1Pyfq7Xp87lG9gCkan+oy3Pzzovn7n
ki3jtejcY2bwnyQnAMdzHOKtiiouxkNJ6pkURsqrQixN4l1NWGg43p6MRrZIb6Pu
iAm8C+mbfnujdZ8FTjhbQ6rhGWQzR3BZjH5WwcDDbWr191dxZbr2D6MAJ64jMWIO
ke13hsD6nHtAVI/T3q6HUvZtyJaIlYiX4P9YXIA8s9UbnbfUl1Ymck8lFYQNb02G
8dD6pfWKL38GDFgDV3pgLAps7Uqiea4vKW13xVg+BDK+/AxvVO/mtAcaRS3qdr0r
v6Ags4FBIWYxfqswjlGzAMF1kvgmRIsg1FwLUOCOd2xjfWAxy2NJ6a6ILDVFjR+f
aauZtkd+vhlKvgP2u7y2VEG6Gu5ec9LBJjuzPle8u3zqINxSIMwD9WnuGP+vVTkd
BPtJwLqFAqQJi07RQGRgVGFPcbMgzpvobvtHDz94cy6xa+6GLk0wu2c86wrfHfgP
zvdgU93fyjZzO/KUqsPXxu5ei0a9tZKz3enNB1CSGfnQKX+gNwI/k+QoV2oZ38x9
MrEdJxDk4l11B1OrUSwTFS+LYE9LwQxD542Q1Sn1SWmjq/efEZewh/fdMOYsPmma
jQSnY+JyJJ9xwdaj7hA0VY4o3YHEmUaUv9KrY06BqCkXWYqtLm0jvaoBiESeT8md
EXk9YQjFLb5s34pwkkCCXZyaa7rzGzl20Ew6MrVfs3WzCidtX7AtnVv1MTzh1pvs
XpKhzM0eEDfN2zXwHUa9QCmOQYpDHfB3aVJtA6vsENPhu5XI2EKY3yaJd7GmmroD
L4OZX8EucxeI2V7amMCMl+7RkEHE+e+imzsMTlv9WL5SUcV3u2TLvztLvR4+FPW/
qF9V4A4rlaqSjQyXkNSOItHb22xIwJ5BWu96C2Kee17lciLsN4RKThQCIYdykcN4
VF77VDvvb8P9s6brHRpK0AJR4/Ho+RqgGYEo2YFCaZ9EesmW7o0qCUK9N1VdIsLB
ooHxVa9XlVTCojfhClZXF8/ZbnlNTM+telwMqpIk+UIeZEcaU02Qr0m67udy3E1R
pv9MkTAPVzXmcNvT42+RxMIYe248bHFLKe+qmsv+EzkFykQyYQcTybi+2XMx06qt
+ySYpPjDcEH7oTB44A2Ws5okxN2N6h0KTi+zafPJlzSaoT1oylIdBqX1fdCA3uwT
MLnOY21iB8MFu9FlRJOCJ8Nge1v/yHxrBNdVQX30Ykf7+j5xrFaELcwYdohD8JEk
NlhQ/1EttWc11uJDwxvbCm6uN28pBX1xr0T29vRNYL+nEnZKRBngWAMgMrsExgwT
VR+uDdZqI1oaB/Z8oRVCQvTGSEcCKNYnccgPbyj0pHiAQOfOJewZB1nKFLlyY4bn
w4Uzt1ZTsLgxFYdAkQdHHM6fIkzqMQ7BinmZsdXoJs+TqmF9wd3lEVwweAzuFFtd
a9HOiOVIqYIxHRXM7K4ZBlQ6TfvRZ+jyNQOtJxWjWifQtypBRUOcP7UDXC6oDN3A
mAEyOT0xC24QDd9xJYAwedD7LC1Q0JWh1UxXlabH3L/Gd0viYd0E3sPqyG6WuUsz
BYtAUvKe200XTk1eNxBgu96jYQlywcB/IOeSQDs8qP7g77WPYnb1sRpIRdy3tcoW
90X1G96lT7AJJYD03UKzc7ueAd4+2/AOx9b4wCQf/61cmmpo043FVAX21ygevLxS
EALqdlQomHCmOHuuZGUhQbMn1A3q4ht2D5Uf3nc2q/MmjGHBoh6e7n5ifY78CjD2
0A2cWufDqLrqZLF9Oh2El5vxlD60fT7cC1hMSD4J7Qf8pRDHS0i1Wu3a96naN2mA
/lVrnfoVOQnsDeR/6+CXnWt9rOCTWOXq3CkKdh+kg0kLXNXbKQIaoRLtr8Yd68vK
PnHqySGJFIhT5Nfd6dcQO/bhWCIucC2U0nMnIP5ARDYy/w3aOE5HcK6FDjoplwy8
JuX+K3VZH/o25JgEOIz1Oh5FYZEk4iTYUiV/sGRn/mcw1JqYRjWVFEw9INr3yAZu
cYsOBPfnpdS1pxe336/17lvuySVx3kiIPN0My0HUNwVn+3hdARsh/b+k4rSC4VpQ
25mLzzXhYOmENEwTLiTdUmRengtTfZp65I5DwHyMa1x16gfZvwPTIgHYmSbAZTiT
k35t1lGsR1cMVwNSLSXHBNERChGlrjqs1BXngPgQL2i/+blQh9/9aAtx22uDeJvH
Loyihrb8GOIhAUu4kig8TPFfLyNW6fwnI7P4RGmZtRI/zzyANxH79MTMa6zjTD0H
zItERrkoqpr3aLHBfS3bbWLGTfM8l1AfT0R9Vu1YvyzUCrqs9T93M1RQDYE/qld8
AhONDZfXjECT3pjiqwgYx8jbm5XPZiwp6PvyzP/dvwo6H/4+pS5veKNorTobHwh6
gHzCQMPUUw+JutGyamzDqZXEhEaDljjoVcxSZsdVBBuHIkEhkPUqtGdhVd3lajP+
wqdac0UkyDkPpmI7IyXZrefHwk6RreEnmHnGTQjpnXzbZASyk7M3tp7k4YysYihA
WemT4sKt2IaImDR0oMyYXWDAAAg9R/G0mHzaCjthfm9Guepj+qL3C8lRqrn8VzV8
1ELLT6MsujJkgxl/hqTpcujrfiRJFxBxpqRTJ8HaFQPm9wA9DI0WAprY26LzpEMj
HeYJIZeGVtWMKfxivoe5wzPF7UI03WO+dYH2YrhclpVhslriuoO8E5Hvu9wTswI0
LAI/TICXx+e41HUTgCS0+HS9/prhL/MnW4nhtPJZsr/u7UTml9n97AeZDF3te9UP
ju4cI3pcTkbhewW/7d6sktYa+oNGLg20OmlFac/K9l1W6wHjjmVTJJxXrAE3zXO5
3lWZlmvuqTDZzsqrVc4lc1DIhQ0IdOm5wl3KtCvl9KF6s3XPwEcyeZyqGU3NjpDY
b1ICXfQZUg6yFgTv0t50vFXWNxupTG0hVOrZrpZhihsD8LDWX/6+MQRLWvhAiaaE
tnV+NXLyF9WOiuWxy2eNOSmOukIud0z3Y+8kPVqr0nbURKucRG9XkLvw2VUzzk2b
D6YunEQEQBoQxrxrHYDI/ao1eoHssHijANGlY/A0/kb93fMrs4ggYa7AYwsHOYyD
VuJ2hrfflMTICyWCo5uTMtWCvI8hLa7uzwCWfh3Jcm+zfXfDz3M5eC5z7EUCCm4Y
Of97yH6JNqNrZMtK7YVm3pnfKYVr/IPSCw/zqRyVZ4Y+9aOAgaEcAwqdvhDdDxNh
wx0xrmMFWpBntVTX8uU6girAE8xpTyxbQbU8aQMJmysA6J5/5BBsRSWt4iRFlyWW
1DPQIjUSvkbjAvo2UFb1UsBJur/ROtFfw3cGfrDAsNVa8Peny1rPcB2THgMhQ5BY
AjjDV8V4YEJJ8OosYNRR3F71klHVJ5RcoQOFyj78olge7gh3sfy4g34DHavARk56
1wU27N7xD192FU3SUVAlLOInDl6XRcIxcV/eVzl/kqkYy/yH5Q6Mzf2wf+iqf7l5
HIyFrt0EMO9sVtn+opOrNPb/j/aARE3nWo0Shi+WifVcjHPdDLNsZ6f9BlgnergL
A31vZPUVBS2RxdHqO1WgNEWNlMVCqO+xzfQut5P2nRNWPYhsV9dZt9k93MZyi6GE
G1GNM9u7v+rCRn79k+rRAgL6LYwcOsjJcC9laRQ9y/xB8CgM0/quE94DkiXXgYPN
/l/Uq8XxlkWdhAE8Hbt03CveC69ymeyXN5Cj9lBk92HVLN1yafHNVlsU+C7wfCzA
eV1inwWUYmhgZavsyXyHqd2T2H/PXwQXdeNXWIQyVHNOsuGOqGeDjef3TmuggTIH
9ufzt2z3Q8YkOrrM6u2nnjkPf+bXj3RmXnpVOufjoqBv5Xnv37A1CRVcwPgANg7D
2h6JaJGAEJxpEPC8bqp7dHqoYVou1unqJxFTa6jAlc0QtHuZ+9xIg02pAzsGu3eD
lioB9qQvKEUaiI1gl/4dwMgufNSExhKHkgsXUncQgVYOg02Vr8S8wfYlCqcf4f55
rIFwl0csED7VYePsaUrbl0AjgQM32lDn4yomxKOA9sQinCOnNd2WKfdYmbxiTlHR
JKxrGKzmL1GOn8tni7265OLxpHoFvXOiGUVqx/c9nN7JdzS3/1kZr56r53ZX6UwD
UBU+WFLKX+USAYoiSt01Qqs7XjLFq6Zd9dfTBQEIcl1bnqliF+3WywLK1gtJBPJJ
7TbsUCf7IRjGqNBbTeDXosiyeUjSP32GOONH5VtYoJc1gPrRQ/DhBduoVz+/H47M
yiaxKOzBZKfH59VY8pn3nE0BTCfa8NpYwsfsY+t8vtUnBCyeXZfk0iJ/xCp+wy8Z
Y+hm1zV05vwOZHHPdsJG4S7n//R8vkUkoDjEtNSCvyYwHBfe5z9XooYT6tGKDx/n
zypBrP9U1ij+eIDSktJZQnaDaWrqj5EQ0m+29CUqhhkfH3IMGS5iPrHIRBvqDbcl
qdzKt05NnaHFd2UVD9ZMthO11Y20Xi5WdqtJsEkUikX3rNTxqVxr0nxzSnf/wMOw
K6/bFyXgYiaa7fV9CcivPSmq168QDsg2BszyjXnhJHp/VYff4GBYTHZ729l7meuN
ds6mJ8M1KuNUOuOeOAdFv8n0ueCz4G+Q3j5u4oe7apIsPbh4U1j+OEh3B6KkiT36
kczJrrOJsRkXiFTkA646RatKhuN/MYZu3R33iKfPdqHkG0jSRFh4qjAP74EHrk1h
Tf4s1iNysVuzkZL3r+ql8/9tQL/fUoOBaJd/cz4Jy2jeGuudx75AVnLs5jUPsGjs
DeAv+75krcsgYpkDLRIu07Ll04epUKg/mL9COVT4y86+1CzOnkDOVK05fG1VmrVa
9lMrN6m/P8LKqGsZC+6bPNZ/hoXJilaJoRO9nhO6MnNe2DwjSPElqw4l26Nh59t5
aqfIMTFxASQjIlM6Bu1trGBnt7dMpZrTh5fZKCDK93OOXkMz92UKL4xcf1Dv89VX
l8VaUT+dpXqaG1rPAynxCLQr9fJAbXRbJ364bo5AxIRFPUv2GkHYzhR1FO+064JV
sxxS9/hCnjPPZiGYKHnPlxoIj0zSn1NrRMG6fZE9gWeGbPtYqQE2Z3AZLAa7jVRt
wX8qMMDngpIdRwh+rMSMzt9R515Cd9cOEhv7pC8tKwSppiTjWYHd2QH3WuADe6h9
LZMPwjpliecBEa7FIb5RrEk5pflDXnJsQ+zv6dWmbiH1rhB9GNPVS0JdBfS2SKcS
GDuyX120UbreNze5tzGxzfIf80xJy+9elffK04D13AiI43cSoBC21aJqUHRo64Hf
kkGIVd9b/aA5+GkxVifVrZXJbE1XoS1u+g1cq8lX47b9QgQ3RA82KmuEFX23JrXg
GpjKtFSLJ0AXvWncTVujdwV6qdDyLfW1X7E7Nj6QNpydjiz3+z6TjDPVHGdSfik6
rhwO6M2bop725b939My+xkMXF7hIeSkE+1GsXeJ7HbDT1Amu8TMUStcJuJFOSkN9
cPHJK1x8myNQxERHsLgCPyoHRzBbQ8CejJPhO+9VyfIi1kQzok/dINgUBBfh/k0E
Wxq0scecHui7zIAWUu/1Z7w4dJvp+PVNC3Wv7KCbk3D2zDa50KCVnFZzKcMqjdhM
GDBSAFqvM1zC3uP03sOFGMnPhdS8lj9kIPLLgxb1XOVYOHvjgyroZoOlRbL+s25U
80L6nI162D0Ii716DqYSbdeAWouR6DGe6/V0pOWu2GIFKt77Rzw9yP3ddwc+ldX4
ut6Lllb8HWGm91CBLO9h1CjVV2gVZ+utVuPws4jyPxFQJIC8PYPv8bgYg4+417tA
fYlwysnqmFz6Ix8yr9cnof9aE2QqtF6MhdQ5m0jQ19xfNp0LbObLf+x3z6xOYhJP
1ydreMVTPP5xmO/Qezt41Ejw6sdMIw9gzU509LqEg/Og2Kn6xsXgQRvkesDnftM+
wHC74AwjhuVnjrrUwLfGacNgJlKaT9yMJmLDwFpPFMC+cI5nDaAMxU3SPVeggh01
893mIIzKA9UzN+hyeFMHlpONzwlq8lY2W6bRYTpr805marsRqSTE+Ru6ejYkRBwf
D/rlxWrb6FEYSvO6iQPFVnZnWcUjsfXyTe0359B/RBq6XkyFM0ukLw+iF5rCtoue
4UN4dMq8Y4FwZyPgGSv7mNionMwiUpp7UtznG+a7oRZK2jizzsmazy3CPXJlwUfy
0KZXrcO1ttFwwRrw0h4sKl2fY4GIuPMxq449n8276tE1xZKfZiOQgnEl5xnyPehT
MB8TXJ8Xjbz9jjrOUUeTPa9IHWA5FBKXSBAXujyVsMuP4ePqaxiL7erc+Gq1BIqA
qVK76+q5N49YPzX4elHqRV14MPkVzQ5vtHJ7cSbH/OrONMOG67GxjZqTWWohyQzZ
Hl+sWUXLzCIYw80js/t8GKYwY8qIiWyVr9C6LT5Q6xG3sYt+AQcUfUP1QkVR6a33
pxx4tE52Ng9L0q99IyN1gwPv0msp7sVvvkJI/XOGV0X9dfzXG0iqu2oPV8KWieHf
qHiDDuvAzLtm67xlYyCbWrcqIr8NfIfS2j3H7+fKSgcX2Ka71LvDqtRuPX8XHmkT
6B0sYKnbmoauT8qtlPOP0t/tN/NSNovtKcXdFGCIzcHMo5+gvNvG70mtPWNvr5zE
EZ9iO1BFRghCaodpzF2az5VCywvGAUBglMHL6CmoUCT0j6O1IuMGrsAiKZ1/zZvH
vM6cTyLPXE4lJJpfjh+Gkf5jVehX9mT/dBEcfKXiZT768oH5Hi7kLMYhdRFzvc08
2+p4G836lzJp/pxdyigR2xGgOro8gx5OzR/y6lXad5QpheeyviuQu67pN04AgDiY
/+LHb9MP2L+DF/KumMC8LWhsen3Si9KXADBluLjBtDunGVH7cdDtgvkvwJzNqOTH
wyu2WQMP4sfpWm7PGlLEvpLSIMsIJEtwKZNQmz90I+slSFoqmzwgY/sSehx0/N4T
aJcIeZh+rAAlIz0UJB8di7MtFK+I5+6kQFkKtR5Dr4hUbTfEuhk3RC6sm7oBH3mF
Rci2e3wlbRESwKGQVRlX2WZ7fEpl7iKOMKxLoa6PnAwoMg/DAi15xtqfxyYOJvyw
FfB+dhu81av8zbmxDM3DDqugy0mrv+lVS3uK1zMe+v94RIjAJeNuzSAwY1K+xsxM
GqGwqNStSK/1rDCbZZu1E0ekDBYcLv8VZWberRaEz2zKOvOhb8QCTZdUzx+Ttr+v
eDDTwmLJcp1GryAKT1keWp9JstcBiJVhPR5MFGjZOuKUZr3dcyFbU/q8WbyEYc1S
/dEZhEoj9esCOs0kj24D8V6QsqXFOCTqOOClJOBHuW/X08YkEPZm4dRUSO8hQPf7
2Mg7lErpJRd/ufVHl8jdA7hIRbvYf3Bvya1w4XmluXVuhj7UPzr2Kc6RBrwt5TJE
GeJJYPsLyZHo0Gej+8ytMsDnmbycovljI/M8rkCV+2n3X6MeWq0h45+91lodqTZO
sL2SDsT6E7BRytMOU/6tb2VlWDwPGaqi9sSZyr6DKtdBsNEdNAH/d+i+sGkvgYdM
Ze8/fSIUCtwFFnFTsMvYCYNK/JcYwn29gjXngvCHv7jRn/PRrAHPrgjKrRwOjvS2
MKCqNuj/taz7Zv0JIM24ACI4Oe5eD3C7H/eIZRsrXzB2bvZitwqPMUTwtk69C4sz
BnxDEZjCCI2Ciq5kVyRGmtjgcGLd6PT3O62Ad/Rsh6OYD0wxWKvZEP64e1s4LWjz
d7ZpZDguVNHg4mp7UE3E0fneLlSEXqDGzjuLbtCZC/qe1IS5ate4gwtPmWa8lRD9
SBqSs0AYVrpIghnfcDP009opO/hg+xwGiTbQEjg/2crAfu4awhmMGwk+xnQPmYqB
2IfWvGABbd9jN5rh1P2gOz2PkUGQrLtFlv8MaPT4j6Eo0bSHnrbY1neuz3Xr3Fd5
mZ7WHAQG3Yt2fXiCGvRKA0d/qkLO0+ZZHlPUfBXM1fqHw4E7LWoCfkFchOiEOgoy
w3iasX1E4kZf8p8nIO58XnfGcIGtd3nB7FYqEfem+qC7FzueyZ09KkoDP8vB1xW2
V3X7Qp4+fw/5acCnSZZmU+SNJidFUcrwL0dvEZCkSGV8Saw18nw2zGmlu0m8ub6p
sWaJtiPCNEpFFGZ6d6yTiNTFtzPKB0cCD0YLivXJXphZr4XTssJoPMCbc7elf1pK
pgH0UCI0H25pRcww4VI9E8v2kMWIMmItzVNLhn2xN0LBWS1ppEhaJJ4FH50g8Pl1
2P9bmFmKIBsIz6+cNadVKkeNTeJdo0NrNuq8Fia32vuwifdf7vpdEAE6HPXevWsE
ieC1DTdaYmTPobJ3cw69IR5ilRwRk7jk9jF9MKsuOcOyFgvfqw1EKDo9cYRSRc7k
zrggSn6WM36ufVlpFQF8KtZEHUuYnpb6lX3b7shZcZEuyILNhMZhV1wbiqhmP6z8
suQ14jfUhbo/LMEUS7aL7N5zWlJKXYEWKNzio5quMlAGgePanYY4MzseXxCxSKzY
+NC+zyfNNGYuXf3dZmZuieDMmAgvujrvF1GuirA+qghkOeK6MKKOm68k09yUyItu
dhtfo3GNlADj5dZPr/T85243SZuVv+/ekPOkIzLJvOTyqN/GDPYbsve378QbhbUz
9lKU1B1jjclydOU86KaGa4VALs98ldzK8k1GEP+mqxiDIhebOCu4CJvxlAh+XyHE
IuV8PJOTW7OTfEYI9j8mKKP6YnPTGkn7s4hkd7yk3epD1d5PS4GmQPnMumij6y7L
99qJE2AhvP7yIvwywIDkx02OneH5OdrO4Y6y2KKkUBktJFfKJUIkxd/Wty59zeCJ
W5SJ6B1RLB3WGyMj+GfncTo9Jcd3eXiIoN00O8cIytSVdmLC4/4UPiwHDgMVWGO6
Yoom9TlBAAlWEfwX8KY6afTON8bqt+LATW77RHUfPeMs0wPGAR3fF2mms2cnjPZR
Jqv1bwzaA/v1H+/QIdhB/yEwW6f8NjjsQpu2I6aNzyIhXpTvZOn4hyvgDTcW8Pdu
WCt1TKp1z9Tn/SgXoe+dvmZVqNPfGKX9iXuHbs7vu5nYMQ86yUD3XQr28ExTrw65
n1lhZkAcPWXJbw8LuVOiwkRVMM99+aNXyUQf+YusBM5utTIAHNpb2HqDgNO3h2Ss
Hsr+BpniPik0wjEw1BXR8puKvi6N/4ecgGRL/6XuqldocRW7ddP35hBHBwvJ9nwv
fHSTFXvRuPJJrUzBhgGGAtsFZwII7l/JZBgkq0YDeXybHnRxFahkAfeaytU5nXOA
X7wwgi99vkM5T//qkqne/PbSoFLkTc523mxZGAbG4PmExfMT7hMuGfyTgIWOFszM
LTJGtbjBhP6dbmSj8uBW9w9wxc3J05CnT13X/s5HIuDUoVJhOfqw/xx12bECAeIe
ehB06ZHQZmijFfXb+XRyqfXvBsnzzXXGvrm8Zv/NPprpT+8lneR6WiDgCOUZTThx
E3POdZzf+Ph8Z1zfjNNObZzEX0C/hgfrX0C6Bytmyz1zSb48lqwbkKPpe3ME0N7u
nXB4Mrm9WxsG1cHVgesqXFWxk5y222bp07t56oWNLfW50cmy8yVPD/e+viKqjmHP
BZM6NC+mxLdLOryKIqSB7qtwzAbQY6mHhYCfM76n8kcUZx1E4I0xETWS4jE5+Vz/
IFr8MjCLufe5/TnazALvd0n6Qnh3A3Mr3OEekYxKDpioHr4fFxgGpBwQbBMHjOlk
UUurwyL8HC0EzfMBGb0pU/1FW/cEoj5WzZchZ+FDiklIOFbW9CET8a32veRGRVJr
5NR5tUEkv9FvmmaDyRHcd1ZA9MaE9An9bwyRcrOgoZs905XQ/eRWoMHGKpdTDf0m
wiqolkeRmLsfLBvlxwEGOMuuPM1lYAKo2wodcDup3qQTNQZRYlnBCK1hti5h6PjS
knn/p9jer60S+ZujVNOiXPkdnH8nFLZPUzXNQqILPCbDWoh/j4ipe0tdvznMpdvD
0A93czFqE7fhVwCIvQy3tfoYjjEBq2gR7gXGqROnAEwZouUP/PoozR2F1MzzxRSN
NKaQ3ESK8X081Gjq3McLi0J5lRPgv7XHKf9ggrZYmUtYN2e3+HyyGCyNw+g4jLR6
K6otrfB1iIWaH5KltEWNUiDbLcNCpMfHe1bg6Gx+TgFWDG1mzLqJxgW1x9MYROUY
5Q0bqMDSRAhu0SwS19/5jxkxRkX4eWtjMqNo5q54tMZJ21khubK7fWQ40Lr9Mo+P
ru/MIh6JSPl4c4S3k3T3wp4mLt3bqZs1E7QToijMNPO1xRzcD7d9jEhZzYiQAzH2
UxZRwELD+t8dsjGDPY0OddcJyVs8w83ma1GHnDiAcOgwFZhvkv5TTfDL5Ksy5AF+
KjYF9kuv0Y5f+lOCUSnxzpo3kjaOmfDzYaw15HT/xM5MuRjYvhGiQ0smXq6Ftk6b
q/QauU86mgtBo51PrQy0z/lUhYtflG+Stu8O3a3ZfZZ5oydSyMEXvVueaPOItNGh
dqVXl20DjiK6LTMw9FmU2Q7Z24Oc9IgM720QM4PjgR/84QBK/V++18KavWCfwsui
blrf/3MRixrZwMHS6Oj1QxjO7vN01LmZK+kYgfjkpTtBfXQqNWKZlA5URpG32aV6
UAKbj/OBSCCZZGeNKKN0pnx8SBzs0ctAjZy0JZ7Hbup+eqILzjsGLNyPgSMsIe+S
+CHxa0a8dRbRR57essD9FTpubR+1usGpTDZ5Vl/9PofagsB3Ez55BWOs2717bQ36
bcgKXnWtLwVNlE5wDg4JodX+JumDkq9sfIMMFOJCHPwScMJle822OQL/wvk+ADzn
TW2/tAs7/ifWZudH1hFPxYsj8hWFYGM6a7Ofv8z9osm6itBr4ggJ7xT3qWWn5lOI
t1aER3Muz+PmT9IFfiMIQwnIMuqFJkfk95w1cXmVE8EVH0wwEl8tOOvhVJgyOXcu
Mgo0sw2ozdPy4eFE16uTmQkErwc8FFmbX37YziP2iHCLQA42Dvx3kEdx/OQUcBjQ
KZF8Yo75oFR1UbOaY3gBG6FhE4uYCc32K8QVHwdlcF8jX9fmOofditS4owLf/ELW
Hv+oprJpzIWuhSXSTfGurURSWcUbj/8aeriWmUKBvhK/HUdDAo8+Dcb8HA15MHgA
NGKNX2FR2I7KNKnXGvCsoIHgGLNxNnLVntyeeDccMB70oV0AWF0sgxtKThkG4mak
zwpNlUNg9FicB3MFU2i76WzMokCFy9kGlCMz5xMXOkbYmcQlcz6NNAj4iQzccuu4
I6XLo3czL3xXrPyACs7rxsF3Z46mUzPfdDBE7j3R3R2wfZZmB2E/mFYQiOIow2fh
72KXw+Qk7gTDBBOSNGXyht2z/t5ki2goYzPxORHF9VMU9Pha7sQzi9Rz2C20iLO0
Ozs3CI45N2mTRGLeHRkT7+8t71qm5wUoXGN7LWozJfoquajdB+sOO3RBWNi4omLM
Hy25vR37xQhyAo/DBh3cAOJb7tt2hLr0P3WsacZG2A8pPlqLiTmnDCI9hCdHnUhR
L997Z77MmkiWqv4M60MzeFje1XT1CTeBoqtrZoXQZ7mPlUtoOIMgmmZMtdgV9+nE
12HNc0bpvUDxwQKWh0SHngo4T5TaqMePlMqpGVEg3hTt8aWF1OBdujBFbbDAO6o8
TblKcSD8uMUUZLwmHIZ0lWPJ6UvXGWZFR7354Bs8gOtBCWtV2Hohs7o2nHU3WkcW
ji5EMXhrw/tqQVRSzu45dWZG4MWGe5kbZvGw81ZXYDPTb+es/lu9bkJgIRm1oCgL
SBOuy891CSRdZbh1W9hDIMdyHI5BDTrqcQOZGPWy4lQgsMHHNhvU9o/f+eUqLr15
PFW4dKFYfimyE/aFTyILLAcxgKrDEK9DB55vry5LmHexGfkeBaxfourcLegOBkfz
biHUPlorq+QaIFK0a7nz5M6V5WLla5n2ERsrRGmltwBM38E+krMQsOIaScRB2Zln
Paj0PEg6cWODFygV2nc8THFJUBgUWp3vBfJSfiVdA90aZJ11kv6F6NPPKvGoyQoi
Jw37iCj5ZoAkvM3zNy9reF66zf3PjkpxtHpTA/hsQqn2Jcsl5igI3q7ycZf9ZThX
v2M2/zpiYk0Sj8rjf8BrOrYE5CRLRqiH7kGj4/RCnrj6tefMphZSnDouG3fjjakn
v+7pKs8J8YP2V8ywlnlm0wTq8xLZ1l5yHC+wsgGWdYQKkcgBTTkB1JF55YdfYQBT
FBC/QYsLqcKkU9drs4DW4NS205HcfDIKPqHN3s4gj6T11NmB6xRKwJsgz2BrIjnN
A5q/yS0MdcPsK6VwnGzooeo/w/81VVHcalmLFTYOCVral3QvkXcvM1XoTY0PPN1R
wYoYwmOnz41MvIUruPh1Pn8yP8RTU48UgMnBQ9el44mM4UBH/9ylRGZ3nradDYdW
30t3F0sPHmeEHAKJk5IRYngTw2E/5SFTJNeCHmINOVcXyspYkus5YbrXIZgy+3Ai
V15iNmxL9LBYxQbHPFDp+WkkLIBaV3BuXN8/deAMI2GKP1SCQ7IPY4DUDIzVzmwA
dlS/zGeGTRun+xMo+XWLBnXhs85VOsSSoex7s1XbrAX5X+YkPzeWAs/B6cxettD0
eaHYIkW6ojkwmGw7wKAi1V6nV46s7uhdsMKdwZmLBWXcdwnvR7tIY+oHbq3jcaR0
9uWVxf6DD7itb5vAjg9f+F9/4PacZh3i+/UuEadCy8isbXNz1BMhvbOhIEr2BrBt
Oxv7IhXRDJpyuhCAydCNVF7bEvbRPN9eKjTtE7prYi7rJZsY4HBuItDD/i57G6KI
aKo1lkZmSB4xRIxPw9qAklloJ+iSAORdLaijkHVVcDvLaV2uazQ81UkDkxmkuxvj
JcoNgmu64dILhPhEuTGMVvZGTXs2Zfc0zkU4BXdFWiiiN4GAE25Wd6nFyG/StfQh
L6fTOD9z2hpawqY9OiBDgDiwNYaa0AMuTxjmleLXInFAE3s2xH4YteMW4f4OmQcB
3ndDjcFrtJNSS83svP7a/6cFqZjbqwiVzc8JFoT7N0Vwc4i0cwycBi5t4az7Y1g+
DzJ3soai2SHm6P9tGmwr54RfBXjZZu99wxz7FUK3MuwqNegbhyw+HHH2+5NnYToq
4WtGv9QrAqw7TO+3tW5CvFc5dA1Cc1DuWhsMFFy3pZfBjUdoHuiQfAM11p+XfRCt
hyfR/1oJM1I95RBO0hDM62B462qwhLUwVDU7kWNA5dQ51kEFIWp41w92Yzc+1fPA
QwRC1SDc14OabaePFOY0HnN9+ApjB3Q9rpVMCVDfLishz6trM7gIKlDq6zT1596t
JXgCiJipwrc8Xj0+HFpjj3kESaUa/Kl6Eqfc3rQUGrKvf4FW63mtHo3hxYZWsU5f
dp2zg83A7HHMyIg3GdU5x2CzXnn1v53maezw0u4Ee/QRY/z4aMoT9DlxCvIG/46L
loTUU5sHuAriqW/Qwjo/aBNhgcXSY3XeKoBPvfeOCeGtvf4JOMLdDU9U34qVnV52
WXZvQXbd19dfN8of7NbtaFbLCpJCb4N/DVamKkgjAOxQYd83c7PUE10C4y75xDTF
KILJXf4kxvtRkJBZnR9NxZRFtASXfycIdvHpqNKIFlNN0/mVV2EyHG7q38Ihm1xl
7AEpd8x3MIYj7p5CWpUkV8fB0RpCZOZ6juRV7E29c6urQpMy6zpkGvRWKi+EEgxV
s0n/EBz6WAj4Eykj6GFL8pC++IR865bEl+hdHv3WH9vLDKUBabrRjsHM0lKQndQ3
pmwH4SWyV3sCQ8/AzosGAMJy/voRYfd0rDvcIXf2MAJJ9T++Yob9ehLBIptc3LFv
xqlD6O5omoJbUf5a8L4GlW3Y4Np6at+vicOQ5+KeefxO09ImhLneavLrvcILmyqF
SbV13RadNvXrlBVNi3tj99cQMG9bIO+2hl1YdDWUtErC0xJ7peWW/4CpntaaqQfb
9uNkbQ16NlAMQ+lMHM/wsHnbmhxAfpa1fqrG1zShUxZ7CFfFLbdOWSUrqjxAwhtC
BTIxlt0K+ByuhylYPRpcK1mB91H3Nc8YVSkxwpSMdTMfeaDPZ7UjVeOcpJMWRo9r
hpy1mPxtLMERPxX1+JyQ7MnzCySjACDksMUnkdzsPJYEtDZMTUBJDfT/u2euqKdR
SrrmBdIisOOidbNDIjoul0PUv07psqmiie17nRo/HopHPeP4iyiGBLSed/gqTEDm
0E8rm8OeHaqVhLm8QumJWGjFlFm9yYWEKGF08xkigz5QLDaKA7Mp1J01XQ76FxCN
GiaLLbuDLEp6TqiH12P1zB4FPw8Q0LWLL4mE7KlKYLvvJS5T5adLqTlwB+l2kYrQ
Q0WQyxnGIE5L1GgbPwCJvYT2wsrvQxW2k+TXu1/nAP/fqhfRjCS77YZhQY76FiOT
yCrHtSlxLKESE5b4/MR5iX6jsNa+bhik1LAMpJEzfc/MkUABuSG1aCk3J+EDCAxL
T7yGF7b9uj8ZRbdQqrNSiJT61VfMeV1ZvzgqjWnjc+VO3aZV7UdPEvqsBK12acif
C/UNnAsfnizZPiF0En7XqMU/chf+/hqx9A3kxDWqjVBA1Er+TTyHR7gUkIqriy9K
YXVWnMjSHlgynRVxTgC7x04Sd4MqjOu5VH3gf/argcl7sjqW06nYVs2H7ktykCyM
GeoiA7lZ1QAq51fvENJ7Fg86xYjk+KcTSFMSEdwTadL1378cGh0WJ1mtWGrFxLym
lgf5Edl4p4OWpnVQ2lxmktgiuIzXtXdTpgK7+f8M0DmnH4bJRRg9CloyheFuhrbM
SS6XgldjoHOQwn/0czSC//jieB9XNjIpRV6e7QmPGXFzpkE+0nxgERfF99S64yWZ
crZkRbJ+bUqVMkuR35r43YSU6G8a9BfjkK2zs/zX+X4oQ/RhqJ8UoLIRpd8kXbQ+
iH+ci/PNxh7ASfoCKcSR2YZ87RFL9Hk3BYIBRPRHmlv3jKRAFO+NWFtpNWU0Uw21
qNQk8//EUfMIWn3lzWMjvSkxKb4BqhfpPL06J8HKh8ihsH/xzCR0oTQdXfyi96Ty
LJj3JkQPFlk+Wih0CHKoeMhGxX2In5VUpD5QS7nyEM8atAPeyfgUuBcyFU0KeT4p
VSiZZOdbjaQVhY84FENVUrblDWRlRu3fqcdf376pnmz7+/kLHyq5yHJlS6AlJax3
MDkl9qbQIX6GOfG439rz6L9NlYJRMuRvqcBy2JgsKzFNwbojLdEBI3Y4yP1tMLf2
Jz1h7sdGYyRYf2Pv7HVD+bnVj4bkjcuIE6tuMBfpXSBJinRXqFfMIu+dfXw7tFA9
mlNLkK7fhARGAQsoDF44qzcGQ+0ruDXv5tk6tDNVLH5gPR8dPremmPyVDRFfq/wq
chLWnyOLS8KsDfcx/HPDqWCRvVRW4kaXkImHc80Q70xo08FyL7sEfPJxeUpVyTkz
xjNIlhkWQGTV0jizcCu7wq21Y8qeJ5Kpq15OW0Hs4IxCTQSY1bj1rbphdFf0IYo7
EeBs04tsB8qgYlFaeeCZDRob80IpxJomRpdLjr/MiVf3Ye28G529iGEk2e4hkpxQ
l7ky7CTMAZ273spEzgvMQOUC56j3T8F99FrbWO1GtDalGZaZi84q0n65pvMX11j2
IRkUqK8t6b+BXPoZSbbRoWG1NuJr0U6IsD90oDRNs6e6S3jf8SpmroUL3JUpxr4h
ol9ftYhW1jVdRnadHSq3mxIyRpMfWkft6vQiJzMcAHdS177z5RmDsmjQUumw861x
xsS9gcMsoMeHy3kjx3uAllneOJkL4mZv+5AkDFuz40+NUJpXSpaIevSg1kSxhlV+
bj+r2YDMGBqbDqGZLm3gCMb4WHyjKg5P6m+aGdVEmZwSHGyuLi/k8X8nJYAlbP0d
bjsNF1WNTQnIgyYyKuZNnRuPiIY4Gg+Unund70C1hSGlMx7CNSSbt+9k1hbzTnTs
bWACJ/7A6+ce1q3iWsROmRULTZc9z2hkiscMEGCfX/DKVLgw8W4N9S8z/eaQ4AJb
IATBNRKrrjW0Zcg1Uom2bfaSBiHrnwXU5hn4/cTOXwUuK/DZIuocCiN4eRS7vx6A
1UlFIoav/s/FlVOVjDNCrhTFSsXZl7M1YH2cZ7nbRuSkQSCxIbnLAoxtHqi94AT8
bFBzRhHNVQfO7ay1OYbA+H6lcX9nkdHl5QEzjPY/cCSVZX9zvh9HFdcYgRLkOFFm
XqipMK5fiMa/IeUR29syBcSiDR9n/W0hdoIFA91IWBQfYAnsF+yv9odhPjJ/n/pL
3iY8M/6FIxkt5TLsQQKQrwrtMW8eDVnOkMVNYWCP2OhHVuhZc2pJ4ij8Kk1Ro1Kv
Y4x1cV/UjkuBGQkvHGuKW2mZ88g/OJXqP8W7muYT0ukp9IV52BDqQ8td+61jFUqt
iU7RLxuCxB+GecMbBfWfKS/oY5zgJNtkW1hDeyQU1zsYRTOQ1JCZ+jDOvL8DTaVI
EMAeD4rAQKDNd+Odu3AHZaTS5a4ba83u4QM6C0BBbX4If15TNSfC59FaKVygubHq
/0FWu1ot6Cm3lqxoaPze0qHYT4Gv9wkcKVY3vEymgCf0RFL5o9RQH+8LN+MlICnn
1szuoPfTgnYP5Hx03mVWPO5IedSr3pJvpHaT1FmzktgQTebpBe4Ga0rG6Y0KetHC
s6Jf1lpqPfyw+tlazWafrkdj9aQ6rbQrjPhml4R9JKriPDc8Rwp6tKsdnqrAJzx+
o86hv1x3EiZ6Yv7mdSzN5lNTs/1+G70W3L7Yeh1ZNh6NKVSZeqdEowP9aTvocgOi
6rQxlek9/M0ruCqtmke2QP5raOZB3GiR7fTzAyEadd+0ccCrlW754P6YF2jyFqG2
R2SxAMB8Q41ushHaoIcrV3g9myb0UDg5P63I7kxN4bqCSCWR0OJZXYTsm++1qV1E
v14c4jAk8HVhzb7rpS9OJsbur8qWnJivAtTxqLO7O2MDfha9gMgbYXaXBjBwYXO/
4Tkv8KIZv9QORy0YuwpA6ZNpe9mNV5A/8UGDXHl1CCHZC7WR7Afb+H0RWUPSwOIj
0ryPWzuSq78ax9dAT7KoG1UFzfv8g/YNjhYtVwTDHvs3SIds089o0AofGfs0gh18
g4DIbPJCqhkGz0yPhkReBWofdDebOEli2tOLK+QePtqTNOkWja+KeYOxJm26BSV7
tgrlufIFp9p0TmloKnSaamp5GWz37KTF+bkyUZJL9IlaEAYLCTuLaJ+OBfCwihEG
/DDEuX+APsoFmotJr0SbH2+6CGzXep/45yAg+y1ZFSevgCM/ZJGJiKy8cjX//spK
nuQ94GohFMsuRyEj6HZuimH85ahQQwARyLtzTmEk+1I7t+opcmVsBmEtL4fbbJzs
piyzFvaUqEGaLxH+Xpsd0c4JtMAoIAr+CyLNVIdJUw0+8lBo98lrQjeC5/pC2wZU
fitS0cSGbSZ4mxiggRbJxCbo5BAqKGDMoA+/Que2j/fxE0LDJ6vdgIiTKnLB9IAK
EDJqRyjitZrcYQU1HFP7rSds/Q5ScfkwohoGpQYCfNYWoi2xU6a9FdeLG0ckxqRi
iUslrxFBiIldf9i9ESq6zccbYvy4rEGr5CILpqXzFzV1bVZoOHXoKxc3dhE6hkry
iEHaZR5JBXHoLEozu0Nk0hv/x8kWRiX00eotH0a/iG5GI0qcXLKyWqA4Z2mTS/4c
C6XP0XESAtM51YK0Jj3JJkO07DrZJ4w2mKO5HAczbgY/Jwnnr/hz4PWyyLXL1vTa
EGzfBLE3rWYTZI98yvNXFA6hM7yZ4jV/eBzfxkaIm4+SQIC3T9BrrpqBOldG0Rgr
NJ8NvSISIKjNjOUDIRV0RMk3LRBjhB7avVV6LtL6Vctpl6e9iWyiDdD4+GVgOq4u
TII0kdeFIQ0RBneFyBuNCxpV/xqxP3BxLRm6BbHso4Oche7ya/gHAeCDqUR+Q3PL
hdzE0mk9k/EwVg1pCWdM9io0HefkujPPpNTHJb7/D+98g6N7mv1jnTeP0GGlU71F
goBrx58eaYiWehawl7m4tesvhPcSxrNZGBKgJs+3xhrYYhZRa+2hFv+3d7IMmYIk
TKsx5cV1H+c+AlFBfWBsu91OeR8ZSGXkMHClhCnEuzA7h6Z7G6TiOjCK4pgVzw+s
YBbOnT86zW0+HDrDCOWC6vr3EL6AsuSlW/pr00oRYonM7dkifoCnfpFB/Dsciist
qYZdv3Oa34uHXwcHRbvoyUNvLuu9RuBeNlPSaYMmmxFqPw95fXJ1zHdNxJc4H6hN
7WzZnaqwIcDOa3HXU4RKu/O+lqnJ6FH0+yY/by5wJD8y/HlEyS9Ekwp5H3LPIXoN
BxJV9c9AJKeCkgYQb8dYqqvOpEynOYLJeckGKGHIsnSaq+v/xbSNxuE9W8mRkFLJ
l+ufb921/wm8LtjaW+Dmjo12CQGLW7fEvMzPpKeK4wV90gimgVtv0Q/NkyalPouM
I/jx320hdU2o+KzEok+4B7chkdj9VH1DhOWoM4b2k8e0hB84b5Sez6cXLWadBygR
NVT7qx0eMNtE2gkW6a93lnNF5E8j2/Basw3ztK5e2lKZxgrFAD7mVMCdVYSnDgXE
/4X9LwBT+umSPCt8h16xz9nWcPVSYLZkZpn3ijK14b+abM4yCQhcWhvH43wb1sRo
wTWxodv+Ip7t4pBXU0GRV88bSjuEfIp5N6MVBGu7XR+MyCWPoCzowDCQzqq2lJJB
37ZfhLVtBgTLxzCJLt/s4R4aoXuTh6CLh5gC3fx9XHaiSBT01mNgpiRoBza2CP7Y
aogwxdZcsmhtUKtZVeopdNGb205Gfo0gcUwi4oMQc+qFAl93dYQXta6go32JCFdK
+PnuV3504R1wRJSeqE7jzS7OP9XcwhINMzI1AYsIpWbg9EqhQS0sCD2MqB34bt46
UCPdiBYJxv+ib20ZRejhwp6EHyEUCcTy5X7TAYiyKVZd5HIi2M21uJU6NJJlcAXB
tjmoN5iZpegSGsseE8qtzr+kwh3YYepF2T3oG2qv0UakOgnbACfEBesRcQ4+pCwg
btChyPOgcOMYNvpWofQSlyYRlNHR1w5SdgVYqgOE0ySfnOnuyLho5vaKYgBUg92h
T6gXGATIPLyVe+qAjdVW0sAlE/44ouSI8H4+b0SWFCGaimFIoopk/jmGQonCGY6I
jdhZ7Ri3b3UoRU1Cg+Wt8RH9jJ/NkY4hAMWw0JeG6fuxhVlwjt78bCxmac1fHNLx
/VsSY5h1JEOYZYzcGa3gfFNKgR8T/GUYBSnMCt6xck2xgBSFC0edDSlfDbPxRG5a
ktluTzeD8Gdh84JFm77c0cxkPk7hBZG0z+VpoDknQD3DUc9wDym0Rco5AV1y1Fpb
oPJhimT25PNl2q7b/5ClykI9hSXHj1l90FcuB3xpCzYorobuElf2A6WbZE/YC1/D
AbCEyLru//rNcj2X1TAkMMAh+TUUIYxphZLWwX6K172Cnlw23gtAhAFSxo1/QAZb
ow2b4rjaJ0aw/PiREUb+QFydzVum0qrvdKhtJDANuv/xo3ID8foqxxieFWuh8alx
k0C6MmxU4/bCsascB+RXZkwcad/WPqZ+w4j7Pqu0LflwTPdh+ZyJxIZBi2fthMP3
WsCYLkes9XOfhbcC5ICsDY0wSB56ihdtx5s1KBzxXHzztuFqPIG3IYvXT+kZKRAG
RWtExllkc8RhJ34eziVyfEnJWiInI5PoV+V8zcvBurWvrk8EfnbP91u6Pi/y6z/Z
nwR6xOm8LQKGag9Y/cjKgjA5c62Z+4uwJkRdavAEg0JqZA5Dt5y1bdZVN4pFMfTE
ZQv+xlzK8IHZRYFfo2xOknefiJbbnrXbRJZjylfqxo1jqxjyAiqx8W+3pQRkASWH
73CVmCC0fZgQZ1C6FhCQjzSHHR0zuBPQCPZKjxQ/1IefYhLjGHRYU1i4S2P8mSg1
2STa+T9444NtbAyKtcD75f7+LrQXI40ncpukOiFR6MX3TEkIn9Lymp4aKFGButmt
0d7Yf2orb/HE3kUsSx9vGIM82fMDfxx1xpvQ8F+i4TCbYs2OBVZ0/B1xzECTcst2
wpQJ/y+qjqjmO9NvKDx6jaWZWOdcb+AoHZ4+kLCmIOtYlF1ZoRLs7z4vyOu8LDbW
YJkf7lZv4Vt3GAfFrwzTScljhzp2XXJZTfT7f4vZcboTQKLoIXRdlNCauE466dwp
XodMYRjRkOTVFgihzIUOOxw6inwdnIhIiXWYmf1ynsDMQ+5HfdrvI8WjfkiYIKq5
bD/Tc4KhiodbrR08PNNoqBs1CejYhzdlInCo5tnci6CCISyyZaAs92la9XL+mdTd
HNS7tLQqiPcSN4d+Y3wCT7SdJ7U2Vzgdvx8loqvS4CSwYSW4uKphfqQAkYwOaeLl
VVAlerovCk530rCSYgTqzZ/C4LZ2TZ7qzP83/TgkU6oXbaUR4yMElz9zwdvnmWrI
Thk1oOHo5mGQ7bqSOJsHTzv6OGkCPkQghzBtvHL3JDhyNxpgAEe4jHlcvvGte9vh
xjfzvo3srVAiU1LtTwnEurYyw/nesiJQY31ZjEXUTZPEkaXHd4SCkbnhh0s1lvg4
SDDYyleEqbPtlpK4XEKBPTuccjELkjGENJA06KewMC+0c1OaTua0bCzBmmQrMTDf
/0qkxyJ+Jgbpg2FkWodFAFYkwdHjWqzvykfwWekb51YvtwJIn5L6XKR0TnMeWRlI
1T4V5uOwBaeTY+a6MUzU/nXPw7Xb4a6Sa6gMY94sgmoCpnhV5iXchbrKhFXLn9fg
Jf8oEcCyX9UNCwTx1gUOrL7VyU7eQgVAn7BlwEXFCu4Uy0xwWqTNZWTADz1DoNU3
pNqHwnP4EVjwgk8qsM+Yd6leZkfwuhC9TqTVgqv8vleQSBElyOP8GB+dYPyn4QcO
WBIjv7bmDnc79ty3b7sjV2IwHM4j2yRNtEzIgCsEP+9HwmmoAD6ed9qiObxNXwlY
BiPklHRgIYjsC9aUYk0m3/bO0pXAniX34+ibD5W8UEowIii70finlM4O0Wqe3kre
ePyMsQhCFNYCJBgVOzRayf2ugTLEV5RJ89I0y4WQP4UnxEPHMlAKmT0RvoM2JqJ/
LeTAXzdLZFJ/3Co3KPKjSYb+N0x9lHqpDjZRUFQ/NzybxgdomM1Dkti4iiaLDEwR
0ggz+2DODdJeviV584ZfqVe8r3XOObliC6Gpd1w9rn0hkdmJaJS9Awcx4mTeXyml
hIcShKAedIwyMSB4wUg7DxPAK9mqRFtSydwD2r1eGtzZFHw1/NR8s+wLKvvI9RUq
e/QT0GewIaY3n88P+ma7jCyEJ3bFS3UNsUXXiuhWzkVY3qcmyt5vQNJVYQ6YxDob
FWyNtVP0OlmSyv/qlWvSs2SswTzw0lypBlTIXbxGUvW06XADLz3zPf5icJCKJSxL
b+7TorpFFTZwqi+z3RCpwy94EP9XqYGpuUl9fKicxyQM4VFHSU1Su9lHOaAl0CML
7VRa7BwU9Yy8P+pjbTDqQ/lsx90xd9wPurduaUHn0y+zYh5Q58cqXGlZp4kDZipd
H3ElWeUQvCMqnCthuhgRYuV+TAQmeohwlucDdc9f0KUS7LfgJneBP38D85Ysj+KY
i1LCWNyxxkgscGw7bXUNuiUYJO2kZ2Y3Z23mF0b6mPq+ILzTVITd/Ca5ekOFByil
UnDmUYtlsZ4qRiou+Rux3LQqZjuZz5M0lghn6ovcVf/JpjgkkcxcifTYGuupAcfw
bw50iLS3eYKZhhfaRHryaePFVjfV69UzbtJpGsLg1UJWVa2V0IJEA8tKSFWa15KP
fUdq5izuyHJbun5E0kzDSFALtONaIKp4bPx9mFIVEj9zgO4nEXaOSrn5yzV+lQvp
zBPkYSL0EUHZFl6kD+aW+aYHgeUr4hjZtD5FpimX9qYA2BPINnST0jHk/JwdEI6g
NUnle7X5AZAumb9AY703mD7w5n2mojMqUj5Iz83ygF0t2FHK+qN5tHxOXgchjaVI
SIN3rYPkwx2aGJVZJdOErpejwMohHEUjqnuUZpcvBqZ6uQ0Ju3E/5ITSclHFNTj0
gc71heAJyk/O4HrRn/216bPCRAMTr27aCGKRizxuhXvMKVBvoUEREUPDLdKgSZ5C
5X5dKxoQt9CsbDw1OWYmrekPsS5Shd540m1ZDjdPUiQ6HYnXBgeqNCArA65wKM8k
SdqZQCGUti/5WXpeOOSw/WXVpyO2v+cDjjuWVYKvGG136wjapPv3CVwRbosEWipX
OQIuCs4K87V+ZxTM/1Gs8EAoh+0lwto3vDQ/2uE2tOjddbAU3VwHxCPEymQtjvK2
nWv50aL0xHZwU6G1M4LfnM4OpMmlhF0QvVKCf616gPu2DRFDqf2RcPPXDMx5SC7e
4KplHwlB7nEGvuT0FYKeu7BNoqgALIOS/ovX12A6mpURYcaNC5IJ7JjOep8OI1yw
0W34e/IOfdTJH/yLtCclvAWsPyaGK/AXBWT1yAs33OfDmBZSuafRF6pRJunfalk+
S39+RSWUySVBmcjV5p7YrDP36/GXz9JgL0vDBMd5GkHZAUm1RPEaQ5moGQgh824I
rrEs46K2Afvv+QXGcxQL2SpWSIpFTepy9abw6rtaBh6awwtx677DYekjG76l1B4m
EtSY5JTmiFusy1z4OzZA9chDcrxHSgNUi0z1OyHbgZfuQzdofAE7Wx3buXGCEsno
w2fpqi9hiEZhrAmMwlJOQlpsTcPRX4HJMKSyixzhbvnfWJkhiRX4hk3axcLDC2Oi
j/+5uNDAzZNuH/uqb8maZ0rEUo6OcnaaU8YbU6ltQfw26/hKt2/Sl8D8Lb300xmj
9/ItRRwg0nSVKY78jaSqvOwK6jINfpXKJcaqIPMO9Hdc2pHUK6iU37TZLeAG5vUD
HoRWvYkSKwFbVIzmwpk1eHmXKpAeng1WQRTnYfI0vFc93a1ewoMM+ileGF0TVsoE
LcJk8grccsT+uN+qwiLdSlKJwoQ1VSus0QgVSr7jZ4NBa82ErTWN6GAOi4WbCnGs
djo1XKtchxpKpSvBWeKLXBjoHEIk2qy2LkRgkMOuBZ0F/f1g1u4GGPh6QPP9mDh0
kVYu5oxW4UU4S64Ca30gJNdaDe/ux9pk4hQXqEkPgZ2B7KXlg51aAvQQWQOwkXy6
h9Ayiba+A1x1MKg/kN6/4X75WaES8XHFeEFDKvmCmb899Cu+KQn8a628hMp84Ps6
GlJ/xLDkCDjPgbHMmZLnrpMXI9aLrcBgWWOawYoylulDWA/VruJmmkYgEPeYuOI8
r/2pyKZEbXw67DlAuVyDJzTQ+qijmq0bbUGot7x/jFpHCGh32PIr+Dpyow1enuyB
3DogQrosQJhjI7sNm+cQ5qcyi5tJVlMb2J7bOWatiT1JBM4zY761aubqXB5/3AXG
pj2F7mvU1siDwf6GWkzmXLhqo4BAEP/KKVQWUkc+WjfnlPu7Upgj/b4o9Dmh94OR
gIrIGoOMgRubpR9QBfp+7ad58BBvW8f/HZ81iBVTFIpBwOkwFoW7FN7bSKcC2SFO
0o6YyHy5J73nN6mNl0SPoQ6zSPKZ/wuupg6CW0ccBepA+gCc3y3O8YOLvSvcW3Ce
73VxPVkY4u6qkkuxjGVZYfzjBJndP21rS+WcDJS7IVHrlg0cvdfVl4/sxq+BaJKF
tScXuKBS7ri74BvDiOEFREyn+C5Qd7WxLf2Zb3JgmdmjEdi3aOxB6CoU64oSsf4A
1j6A/sJ13JNZTKuwUg1QZozOI/N8CGxvyBiultRHZK3KgJkAlk2wUkpK/T7ZeCQl
DpjAh6/IasxT0i3z+HQOFRUbCRSMPX4Uhad/6Zvui1MtWtQ1mLZqgegRTw3hcEr0
0a4CsknNpfd3HcexBuLSDXp1/GVLzmf2LqWe5/wrsfIpojxCIQbyBbFZ2fwBXJpA
vXOL0J65Cy6uHVYVzIALaf+Cz0DGSW5tmMiDlQW6oc1ZMy1u8WYwaGx1f3odO+XT
KlN3D8eO/5h3iJ0hMLjmCqDdP6HDKRZnw25swKDbgnHGQhKx+kVKgzp28xH0PAee
5XdMXj2mz5iw8ysSLEq8hDgjZg2jy9lPXWKRDmn/vz9qtJBgJunsGvDO7D+d93sf
DytY5LQ+lL8pL5nEe3m/mK+QQ5ND5/M94iRHSebtGBgNi6npdq0XsmgSEUZYcK6E
46SpoigAy5N2sKEmKpWwG0o1DIJWfM5snaxOJmGlaRrSif+vL0lXPNCBe5hCaPLG
7VrMYTF9j0IuJCxGdjoLXEAVkREZSInuAhrvr7mlVrr8CeYdbsPIj5mCkmy4cbgO
UdR00LUSs2LrcjP738q1xpfRnBivdrNcs+JL5Pic3hpMTIiz1Sofi9mqZhWQnmiC
iuV6vKRE/iuVopFwVbTTr2W8IQwUXilEtLF7wTrzS1kM5bO5/GG5FOI7PdZukhPK
48it+PByn9XQaBGZLWNo+nzcFjaMKE8xSlcD+bmfdwR+kyatpbHUbcSFl8iErDT2
BhWhUT0ViEqukjh+J1AJhVixFDmGes7hFaf8YjY25sRhcjp9AL8MfTIOoAbeZXZq
JnfeZ2xmqy//MWcIDBjxeBBICODJAmkGT4o5LDnGMNSHSGcW4doQuQjH0w3ctodl
QM+SAvYnlYN5/gSaGkoBcv5yAzHzpLxpTpovMh0QCI16tdcE97Y0l7dZoI5xobN+
vc4CmcDlpIEcN40g3nUKX2v69ou+o/xLfYqOeGMQt7V75uhXMHVQ3PGdS09dHSd2
DYVfltowbEqrarKGTbS6h9BPnBwHSInmUSfMiwcMHxxA8rsDJAWyTbfTNeOGJWqc
mJ1YEGHDWQzRVEeNj/Rf826aLobPmqDzz9OcaVdoI1REJysQz4ZO91UWQNlaB+Sw
s/boFHuIG3JYITO1IpZrjIY3+Po/l6888TSzJGxDl0oHh8KZZ1XweLq3cdipY6WS
g+VP7t48Q5m4sLl+nVozlBV3PL3KXOONZMKljkZvqO1PNyfI8rFuHHlc82Lry1Qq
Mltwx9W6dp5UZHwXJtsszSDwDWHibhniRP0db+njoPd7ljrilxyYTGdfH246N2BN
Vim7TUMASzqcI4RbdtxX7DERB21OlKt4mvyZQd424HgP4b31J3GLlaZoaUA996LJ
cGobZ8dxdOLQpI7+ZfKzjtkr4aaJ0f4j8XrHDMpequf9av/iQmzSl2KOldoIwbvh
Cw9XXodJVl1Mg0j+G+VSuxwZGpSQd7y77rtCNMtnS/EVn324UGsPaNxCGEZfBxq3
nNtZS8v5nG2c0xeeXgpI9VMK2rnaR/Kz8MGtfeFYVfIiiBsGmuPxts3cneO68TD1
P8BWFVw7gTP1LJ7TWh5iAxtj2jn57a20XKb2PXaBzi0cHxXNijxQs9/8aTcZca04
1vBi+lz/oyEITR1MJ9O2crCc/HDw9zS7xdBi/8Z5V8W5zCJVR5TxZnZPPAAZjy/V
bhseu+2JRNYioMft/OjGlmQFJKKIBkWr8quP4PzIl8GGZtqVGF+gGqGLUSn7SRyV
Bp2GKdGcOHYfYdBHGRSVsF+TwgNmU9WIAyIWAVMrMiYUoGzAr5DJA3XmwBKcFn8K
ihjQBokh10ZdnZzra9idO8ONnS4olioO+gmfseXyJKv1wiIwe4PAWr5Vi4rsntpT
SJCwyL+lAcgclWe7XElsSeoUvJ30njMO47bIChzjpKpyKPqqc1UN8DeC7bJ/jTM5
k2vUczM+DdGe7FcaAGWYcKmyBM9vEjDNPDEKjHqOdNUL4dVAvd7IrWMJVqbP6Hhz
SPCO2ggH5gbXgIWx4oIQw2rfS7dHsPenIsD3j46Cj9mlv/G3hJ+JzyPAggdc1WQr
6K/ur8OZMKYLb8rq/ScdZgZobHtGAohnr85Yb22V4/i+5u1dkyW4AwgiD+rXcqcK
ff+SyQWnXh+yjMS/ZYjRj5SUawKenQOIUR3GcBKpz8sU0ljT6/P1l8+BscZxKzKU
ROJ6bCWYGS0E0lVFSZVgiA8T3oAMAnLKeLxzhhyeEEe2zhlBGRnMB7X04bxyOOH9
fdwitNKWUETNusVoOkcR/ZYcxLpwgpaEUSaYOUSl5znNs09MM2x27WEVW37LEYae
L8Ymir13f7igdZyj11qhf9pDRHrnH63/C2lPQvoLZ5LPKFk4rD1n4e1XL1hkxtKU
sBWNCueLNI1+Aw8njyE49frT+BMa4HqFn2n8e4YnYuLSt7+0f+BgG0JXPn3el71I
fwDcqZ63hlZjQ4nngkIpDxuJS0E5FPznQrQUMhmQyB42twVa20WKR/b1ciN7pDDu
AA6BjxMP2DWIl8OMhG1qssqwK+pjUFmLAD7G/abJwL37yJMoM8qREJG+ExrBH5+P
px3Y3BArEfjVg9BE/F7xMY6MEl+YyTyqvoj/ldOsukV5n6toP2Y5Jud5II1+uuEY
/uPUdglE291bC4uKH2YsIKEdyqgBzdewlyb6tFGO6TL133697QAdKZ6SM2PHL7hp
iyUwEaeGUL6XWoqUHtO55aaO8C8v7w0qg+2OnfQiMgeXwb06XgHB3Arnild0Z6Rz
4yDAxUwENQ7X7ab/Msypug==
`pragma protect end_protected
