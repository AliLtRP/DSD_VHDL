// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dxpJQql+schZjXXmZeGKj8HwbvoQhZozX5QWJIzxIY+xy/p/1YBMHAsTBGCJNfqW
kGzZArs9eUGwu258ZapmYBfIkvJbw/6LXR/+WXT87WoY+l6PC8aoI19zfRAqDE/h
ZhDT/EzvQUU2JVKp53h4sQ70lksZux+j7LDp/fRnHYY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5744)
Fsp3unOrN5KG1WGGMQ1bFqVumzBPksW9fSd6scQzw6iroVdgJGjBOKsc4gOZScMr
Z7WrdWoOPIp9jAHO7+93ylIgqdefvJ2q5std389wlBlqToHomwe/T+BgUwJKIyHf
eA+COYvixWiLTHojgBp8DQNFf/TZoOPQ+mdeDyB/wlFnPXAI2K+yrdzkXvz1HOSj
NFkUORDWE5zGVQO0wcXY9IC4rKilpI39YbeEefT7WhcJ4TSzz3J5kJLl1rVweL+/
W2wtSRgbP6R7arKbJWibwOaqF9Dn1RM7uL9TfyUJXjqat9flCXHxiMX5iB3mGT1R
0Jo8xQQybBqezZhJ5HApDhZQnQxU1/Ra346yeE6UxhPWEWIR4+2qqoFf1/egW9hZ
Y94kna6SGGsvKiI1ZPD9URucGeBJguVtewg0q9ReVPda5l08y3EOIx3njT8bmzZO
7oIoNpC4MLW/bfVGxDx/c0MdvWs5lzFKMHZeyjzFCcKFPry5A+u+d2EIOBHcmVOj
kq2ywhDtniqdxIdPdSMnodX+/iAy+nT+ROzZJ8aTeEapmtiixQHpJ3qhTUfo1Tn3
cyJzIb83gTWiGoupLrMGhrNMJVFD/DGvmnm1DclEbFD3SnHGv0CtvUkQUnX8wZnf
RNbygD75KDoW4mU3nmRxf5WP2PnjgJ6O3Q2HNRM7u9jNp65Wgf6YtDAdKluKViLU
yvTu8nWuY6Zo1ZNl4TT4SSiLYs1On2KBD9GdFA6kl3j33UoYpeSSkpdRIsJhcwzc
lQD3gPZN1uGD6NZSBcgCDZvelpkgEtT9oq/WPTECr0ov4Be7LUyPZAogrJ41UySv
IoaQvkeTwdh0wJabY6MAVc8jCvu2418k7NPOqhh31Un9T5xAOnqgIrzf64pIX0Jd
nEZPtgWyhvsPJpKRVTD7ApGKZGquRuoczfbQ66WYhx49tf6v6KGzyBEgXVTzw2F5
jnW1DSu0AeRhtQYTaoedCSf9q4fqU02f11PcC1PGgK8Uct2O+pg4+fkrrqkvHJWq
CRRCAQL98RuDZX4EgkOP5OzjhZOtGowrCXcUTfnWxftiyqC5YU+4IW0pqOWXMIfO
cJInT7WMIzoU2/NMxXDW3k/9kg0Xgf1OMWbvts6Bv39UlMhutuIZilVbQLLPYahu
2YbsZLDM8pc8s2kxd9fjaNbTVGN4FHJllM3ipLsJZF16KZVcPJHvMG2o7YxJKzJi
xj0w90btc3QZJoTSS2b2n40GAENPCGv3PgWtkX7Omni1P+FlZVLYSLhpMNwPptMf
TSCKmva+TfIYjk18Zwu52DCDLN2Io4jGd0MUS920CInsm9fSy1Z2bxVMPX7nc0V3
+RjF29A371p7TXFcd+HGSLc9UmB9geQ55gJgGkk70Fh1GxHuuM4J6hddSemc6yL0
W+j9WaTvyo4XkRpLLId/EwZc7Kyd2klz8O8X1+W8RQimlcwUCjMYIgezZV04C47I
wdXA8IDwmoB+FHIpWRhyClUP0+OPbosd/PxqKV9Lwl6FkgY7lmH00hGCMxdAGPCw
VA9e3MgJrAsCoAPh64hHGzHEMKEKlwVENY9rX7+HbrOcIXXYQIbHOIRk8r+jMBhK
lISrilWFLd5ce/Ai8j99DItEPsyUJHCcRzNnJAJyfcs1WPYI5osnyLJWGfqaypog
dI6jDV+ogtrH6UWy9crTWV3MuTxGMaiO4MoOxmlvbrDsqY8TviprnL0Y0iEPG6eM
OflS99bYt6sWgO8n3Dffw7MxaLMoes4fgOtoAl/hQo8FDnjaurcggD/2em4C2YXl
piKSXnid3cd2Ww9RUotaA9Fc0MDs/K771sBCirGMg2dO+xWkCrxAVj9kMYsVQjCY
uOUUvt+NzOXuEr6iIPt0iWB0lma/fX0m2I2ekzFKeapFBV4IDxrRdKCxi0Fg0rEY
4N7NYofyzKVRpErRRHZmbqZO4QGNQ9J+9twk8rHaQDCyX+1HKULjkhm/nYcTD6fc
JpXuMnuGOxH2s+jJBuA4BPcY2Hu5k0YAC6tS6e4IQK0vByw0JmjaPtCloJQESx78
dAyhl0RKfD+7aYafaDYI1P5V1dFk+NB9oNAbZqYp3A+Zl0zmYhfbmHjXXGzJIL3y
hDp476NT2Hd+u5zAZzApiB3TvgXzC/wyAaOWLCJLs4/PoIJOZ7f1WanzxZsUegIV
ElfrS06qNqR/5+kjkCP2+3TXrP371/OyZnnIaBss0LncPchmWdLwgouxaOaaopov
jSaWKiTUFkt0fK+kidUFSLeRikRI+9RFArwKVLJMnZZY9FE2OaRXfu9ZobTZ5tSj
dmdn4/e2vKtQ0eEVdkSCi5xubdv/yFLPn1SmY8dR61GVyEueWOvTzUgiI1Y7vlTq
aj/eCTGFfTqsZ8PYmTbbyQQAFLe5yoEuukDCVpRBf2jMxLPbIveQMPVsYto3XIEu
Tm+6zYPNhWpBx73QUzM9h2v6xXvDjdB/uISp+XoJXfAk1oBBY3p//f51D6Ktyyns
MBwU8IsoaIpJAJhOfWawbwuKow0OUVAC9qtMQzaTZiENpJJCdV0pMz3QrcjwK1eW
DJZhNr915wd1c+koFD5rxIg+shgBl2KpiBDhE3CjwHcXFyr6giEm1T+v1E0pbiEg
O0cwKKWgIS6WtuzkzXiDd/dMVe991rjCIsMFBhIB6WBABbE8MyAygRMkg6d0WfGw
kuRCi2bIVWey9M6zqRTn6jm73HbKfeLgqAifzvikvJR4Fp56XOiN3ULYQ2da9u0k
nz4GzvtvhR9yXawzKTOM0pQuSQi8G0cP+qS+y2+uCJzYwZr/Vway9tBNxzNcOwrt
4iUCKqa17mvA/57VYARb5yCzIjqFnsppB0Clj2wyFpiQJcAmh+zU2/PAh5K9n+Wi
aazMchtCkTKSQvZl4xIXNOtrqQfDgj/cIKfDCTh4ckRcKhODVejhTeo6MnB6kOoo
IiI00rieXwB8Ivs3CK1RfD/RuL9Ur0q/g+De3XflNdWrmYau5ke+baVqJRwxqOa0
KLsHa1htt7cFQ2lvWIB/oOrv8FLKNhYz9za1ITqojZLfm+hrnhuPJ5LzC5JLq6Q5
LH0hkwaS2JURB26qad7DwyL6mS9CpeFAewSiAZan9a70+bAd5qhOuIPuG7VzaTtq
7B29su0IQlJ9LdzhYKungIy51KNFSXRuESIDwqCir2QrRAeVOFzJ6Xa5RDEztvWH
Qnr5Rb0UNyHkiEf2+0sQVS/yFLdT74/A4wUpPGoVMOX6u3xQAPjU6djQ3WAAK4IV
Q5DyaBAbdx+T++g7bIu6Rb8nJfz2GkQSsvy5TMD0rLqfyD+4QuSQBB3ssVfrmc8X
d/fhpyUy5Fd4wZqRFQy8zPxAtV/HRG9N4RidkKpVYhuntBimToFQ50B3XLM99PQS
qMIpxbqpjWTrS7diD4l3StZXapvg5DYg1d4ALrAgcx7UWKgHy6hME8WNoGevbFlK
jsF43QTG1u021nHn4ZhQnyyHReNX+pvv5QxWQc7jlRwAKTMilhB7Aj+XMYb8gY3b
bU5XRTMxl1iluhhJYTEIra7EFpdswEGha3sCGNAy8EM0Xk9/GIk980Bp+PLbdbCD
SIYDNkDR+2YyP6tGI2vF8CJDSY5qQj5MiSVnKejis0dK+zeeJGjdbccIwQ+aGcXH
0X/aPluoHPlFCwo5lA0QNz+XoI1HtG0rvpBtF5ctEsW93qyr8HecyZLIFLm54o04
HA6JUrDz0I2ckCz3ZyRNMPhbYXL1fEu3FW5fdFB3b/xz6GxmD+A5AedBUsWkDnRe
pvSrNXhbEqGIS22Qc4s0EjJMS+1x1FfOxkN8HhHl1rCz+ONzNZLUTVYI6Ikid47B
hrJEIXnpja92ytVjUKu5yo1qiz+jBCyqYIdSnqVc4J39z/K09UcBZXzau/y2+J1s
XiBwIFGg/u/MCmHC7jggG/Ao7A7ox1dUl+z0PEn5dYsJgkr7TdjrvgmMINVyn0J3
QGWhHYyVgOt7oE0zD2eEiHsVHP5MVIseeYg/waVVLjcz3aNqGKQ8gPxf59BJhsFI
XE2lgiHDM+Pl234b005IY22i7t7vlUepulQt/H1VzRQBBKdCIP3m5WRaaM0GJkRz
u27Yi5jBsyrKNUzGURaxf0qsC2/jSVgd4E8kbMi2vVIIjVHwPZ2x76pf3x2qPX3U
ZZod+MHFJ87haEmgj07nYxks82nqmQgxgo9V+AznSHaKFI/UwkZaAe0IBbOIaRMK
OrRdI4ikrIbNYr6Q2tk6S1gFHzsYn3BQJXpmqfJrjaN7/YfE2NmjsNW2h4Golg8u
7KzzKGvmF/Cd2fV7N+LfDiTZy2uoXNbYb5kHEBnd4/kG7IgTq76gJDHo+e1VGc3u
gANEf9kLDU1FYucjuXLClAMd8CskfMVRt5YeWIFCXxdRLZO2aacWsSUdJGXh3Ns5
euGew9qfLrV+ssTQ4Tu4YNq3v1/YxCVcjsS1CSERZijj/aGExfvVAkT40Z6x0/SN
ikY3tqa+OPdjgEYThm2b9aB77oCccnvgqbnT9kcSuodSYDdzOQFJcWBPQF60+hGA
rdTfbxXFCY0efINt+J06tjT0hCIvehhrJMLQ7S6m57IxFZGQtg+FSEKweMP23Fwp
3lgATmIBeiXk8fSKQPKvnn3RV4JC/xwrgSN/NuQ5Tp7BZuCbiLZiWX9Ov8R/3xrI
o+KrqYySl4lcFNHco583cUA2mSuCq8EIeje0csbkmcpIRIKlNdb/PCC5TuzLX7RT
0REKg7AOd+LlRcHGxH78iOimuZQAUzZ73i07XvjsXuQcYmgR5m4h/2aoRa4vzOPt
/6ZsbRMCRbsr8aUXMBTna9epWoRTcU5tHToSriYmh5IV6DiMllKZ0kgNFPToRffs
MY6iRfVMTJLq1k4bRVhUQIOyXGv1Cc2dcLxJsgqoezFTSp1LPELYXFhIVftwB5yt
X5qx0ag4J+nCBoPhst0qdVVdTWOS/+xSS4gS0hZeCYGUd5RUbcYf3LYbMIdL/MBg
60Tf125Q+9hxERTQcb3XaW2/86T4ZSY9tnJi8/5ek8r1Qq3bH8Akb0IId3nBJB16
uEZOzZCaLETLTRWpSCETng1/BymEWlARhnQJVYsCVlsfdu38RLSOxZzuEKtelE2e
v6p/awEj1kNoq//aNcMmZX0AdKeTBIlweU1qw6gIwIXQJML/+rxwmucjnvouslQU
+yWBv+MzM/QSh9it4lfX8BI1C+FvGC9gXuS5hGfSvcSsBzAoGd6owY7UcW11adzH
rV+u51+Zc1tDaU4bKXr2N/PISvl6JhPYXpnUax0Xxf5EYsphq8QttAMVk0iD7HtH
TqzXvV9Q8je+rIw6zfHyVRYjYnOnla44pDuv46V5NYDW07mpZIkzF3YvSx4nedxW
Zo3ejKLbiPzyiSnZOVV6wFpiQpPjeGB9HKS2ISdQATl4qDTb3iHm61XhugtIr+UW
vRjfVKisMbT2O5it89OTq11VGKu+VmWQtZ058Lh6NPyWMZRR5EK5FLupO2ToLaug
d8ftzW2d5vVsnm9Dv38H7VoQyeIJ7fK33C1WqWV39gPtyIXwjFunG3h/M2HiEGTA
3ZInplvEWPwHSUNL79hRpHniSEtmRf6OqJjNPsaIHuTsNIEREwfKEz/JP4Ii6Zu5
Woy5w8yQOkPAYFNAbP3NeGcUMnZni6jDX2JrLQY6SScWarCc83Vn43YTDLQY41+H
6yMNo6NhlcRZnhlipcAxGwmjgCmVCsUry4Zi6EwOfZZuw2JEnibqIrzK1T8wz0Ok
AN59G7YqaSxW6X2V3SVkmgF9r+LJsPJprPoMxPL/qIAA3J9xOMQ6LB3N9jfc8NxU
/ufKYJOFZJz2NV9DX3KunT82d5MgjCQvN8zmJyc4xW6ZmNteE8HNy6Cp0MJe6+6Y
MFSJw7Hob+kETmvdUKT+r3lzhEIAPmRCm8JpSqnxMbT98iVL9ncs7cBfhKb3hUBO
hRnm+t/kenhjLkwhgPpmbaCHWYZKux60WJZotdX2iauzfwJ4k3CtY7FKhMiX16m+
sNyaHJXLZITYEL+y7jd/996qhtW+ZwvXtU+PHAolScIMDAahPT5g0lSdQboYtIuS
SEc6uJugYWj59GrOnBg7UpWOqNghupEqpGmP2VqIIPpB7DWyw/heE4juCR22xchp
Vk7RKaXG+ZC4dWsBHthuN/Nj39lB30nIKEUq1l5zOXg6Pv0jAIxu2p2BX9/mdR1f
JvOg03u8iOzR6JluRvGihb5U7A/exbPRrucgzQxa9eC45V0u7VwCQ8y6G6HA9htB
8KSSXdwy11SVx9bFkW6HGHLrOsY7c357a+x4ZX3VbG8CYCrj61bFb0uuN8w/7PZh
5JaO1HzlQZST/IUXRowFZZeF4Z1QBoGePKa79d8uENRg+WwIzipMjaYmhpCHq+OT
I/LQ2hyBLc0hKjEv7W/PF6sXDTit6YkjLzM6eJT1nfSrZ7+KiiAJozoMzxkHnNxc
lVyUcP3peA41K67ARgkberYuTcgHXoClYa1AkEkn2Ziwf6P9tJBg0HdLk2PLC81T
8iZfBPaIxT94QwqkVe/6yZdikJB650h3+oLJ0jzjtdtqsftNPBgQ/UivXk35wSye
W0avFTHVOIJPoHlwGtE4VLr+GQGL5zVwJ4le3QzH26FD4Pr3u+2jWvMWe2F3G5PI
2bF5U8QYe93HFG4uY3tLCAXqRHAq+n4FrcOKoIU6UmficjUKS8HR37ontiHOVka1
DLqTglHFFzWk6vf+cNEyateOqjPpm5A3WQnwcz8NfT4bZmcqlLJEj8np1ERnbSEA
s4tsVrYVEtlChfRO6DjRSlf9xbg9U+fcPKqP7m3pzqeCVtzR2D74x7uO5RZDALe5
RwESlbgA6v5p0eSUTM2C/6KzwuvGuN0efmx5QGc9JwRZN2sHs7t/Gou3feAaD4kB
67aux3NJeZpMLsLEtPlGYoL/FXjOfh2ci4OGewiHs8k8lbLF8Vfct57tQGf4hmeD
orsCBVhBK7WeLJQ7WDZB9PFOhgpmY1LQSXlsjWWsWT7t+XCi6DY24t86/ZqRlpfE
vUXeYaYhqyNZCcegfd99eqAFSd28WIlkCj3lLnxYvwS5hBb4IOJyLBculj3Dv3vj
cLpRA7hktac5LfJya+CsvPCfNWnNy0OGsyNHAHmbx5PZQae/WS+dYqWBzlhW+yr1
P+nzp/N+9+UsBOLjVT356TsPQCl2NQZ1VGLtMaJYnC5lfwjHAecITf7k23JCENw2
MoB2kn7sa/R/54WJLLfIfzHQnG2t1egYC+w7qp3GezS6ssm+bGpiKMo4IpWAdBGJ
NXMhjZCGPWwXchrTYrKDXpfMq/An4gvhP9xklyxkRqtBQPi2Re3ldzxLd6rPf2tm
+VPyCR1J/pqnmJnkHprwiaS0c20xVrtgMXIOHPJOXCsiI4Ra4CpXxr6cMPIAl3s9
YFdmvK7RBfrZZMb5+A0+kY/2LnTNTqZeOwD8STcbmU6WBrdo7Rf+uLsiIH2H0vSb
/hecrWEn+W+RUV5svuEXIubCdeT6NrfW6Etu0R64NNiuNkt0GgVHFvW6ymroD/Bu
+lPKIhJNvmuNjWrP6hlRO87C0yjoqq99vGuiKkFDAWjuQJs4mftHVkEWEyBvNRbu
keGJ748hmXT5nBu6ul3qSRytm7Mymmbf1F2UyM/K7z0=
`pragma protect end_protected
