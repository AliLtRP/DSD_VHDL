// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hequaHqKzbYDKAfDddzqnvvuPTRRxf0vgjCgfLDU6/xYhqWviDi6A+1Gxci7Yc7j
EJf7UF5VLwd7PK9xWlWVezj/eRmRxpe0fJgkWr4asUtbOpccLgNc6Rz3JEIRSpI/
c+8hEcio1lKoPbrJu7mDghwgDCxgjwQA+2Bm5t+5oFM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45200)
eJn2wo5iZ3q/zR5oNl5SqYlehFljjdcu35LT+bPecSOnchgjIDVELM3vrP+tirTD
xkpRMl1TEFZMFZV/61s2cKRP/nTG7GxtmzLMwcQ0MCw1Tk0nwkHqbKcyVF47yKLT
0JaxUKTtFlWNWWkr4clKwaZRozl0gGWJz8oMa2ssuaeZK84giERqoLIgsYFleZr2
zN+8F9t91/eJyjC1WgASfiqu4+88VwqzMMSARxPcNu4lx5rV1MW8fqDDt5GKH6Se
JBLe5lQRcmsJiGVTXaEQVXAAd0ci95aoyzsRDLSj+NEUVSwvqXqSMfwinfRgcgtp
PCGItfIBg4GLiRPPJz3gjQhtarQxf1xyhiuS+l5h80Cksz6TrS3oIIiN94Ujpma6
802p1dKbu3UU13dLQ9+x1PChZvrxaJqaWC79uueG+SClwfrGOULeTr++CGPhvbvm
el+Ir7tQ9TBjvwGWlYqMNLvJBUUxdks8Q+9G2xUA+E0UNTIlOMzieCeHGpk6snw1
5mVH2/agj3n7lVJMS45k3jBKpgZyTsPyKr/xq0Eb1FwSqEmWc1GbK6cs1Atu5k4Q
LW1+aEbBEVpDE8GKtr6r/r4fxEbtKTSEcU/HKvae1sz05mNk8TslNC50UYsbdtPw
LUwF2lvcdD7CU0y7kKncHah8Ouf4cMJHDC3WjjBK2R0CMqnKWGMmxg82J9nDPtI/
4xcobgUZKNQtXuwhOtMZKwc36iHD9F9yIJ9B9q83+BM2fmDFDSPiGm1Ifo06DOyA
Sq/694kK+XfxPRzxI1n789KO9UCa+keL3zm668sgVQ1cA/QkSTXlWMxy+nIoenAn
CM/h8whLmrKgvpZ4Pi2KVHrXQg3H/li+q+hDwB7DziyKot3hFXbhcARNK+6pSdv+
U/EOjWs3uiV8Ma9UdOD5KehyBCIBKTYlBWDHnXj0p46DM9ZQi9wuEgRUIZ1PeO/u
8MpFf/eHZ0WEq4S6pgGgvug8HzI6BiGwR8/eXvAPr3qD0MqcSCzqSgLzME7vcOs+
HWKVHs4PZV1AYvIHD+q3zzBry/rQUC3Z+PCzmpNyQ4SisSin/9jj1FuCAUkqGvsK
7XzZK+7Cq/rd85bScQzFR1PRffKBGtBM60vVP31EyTqZW+pg/RjoY2OezQL82i6l
GF0DAsR85W52amHaQJ0y2/tNCtyLkehCCJsPgZn20ii4JKiAn3yvWHALaRzXntE/
vrpWX9/57y1ED4DgUaEXYqZi3QP1grNTXXpJXLBvA/M+69kM4DO1oBxhcismSq9Q
Kxx4e4Ow5MXCEbGteIFVqQ9+26wwvt0SD3fwvqOM4sXNO7gaXtZzXBX6FxC9Ye8J
R1ktx+wvBb3//hSjc3ZtO/sadSDtYVvuaKZGGtOZeunNvD1mtRsRIVvIvnnymhNt
fvCXgbv/nvCM7l4MPK+zrr5BO6ihfdNG7Tp4Esy7VfI8iQslsF+JW0/WL11ymI5O
kSaW18nL9muKaU0/KR0pm9moYYZPnDiCdTPcWSixx9g5ISUwF3U0p90SyGNYalea
EP4VxBwJhkiBm7wXT9HuE8RxmsC1iTjQYBh3xRUHZDkTxIy0Wl/c71EDY8FADMiu
H0tORQSNLrHg3nuVPK86gC77I5XNXjG1xRjojGFjXLjITjpqokVOjia9tUNNpsXF
ZtzMODN5mcq8HZzWYiAMiYg/Rm/WYs+dUEofysj2vSM4qTAHVnNNyofCK2n/3n1g
pkuaFfXYGAhmGcJz/YrMKjj58JOjaWf0uSZuUdhDQRAJrL7BfYSL0Yn8CjR1nYYR
vi/0OAFT7kDALGesfO+OwDWGW/SsD9dlW0dF+zJm0ezsYKbuK3Uzde44W1k1UxGj
O2Sw+EgbdnMGTWudbVVcVoOPX4KfZQCcwBU3QnYe5gRoeu3WUqLIVFa/sKOt25z4
Ezx1oII09L3mmGIYFujQAT8OLuSuxyTwMO8sDaMxWlcttBzRNkdh1evOt0miP/3C
V2WMcqA2uetEIc5i7FHGoOSSR7ZpqTxBOwkJLQHWK+IFD4w7Mu7BYlkZDSE3wZyr
QbHQXhiKvljWfWUBhmSXe73FfdCInS+xLdu7/RG5JbjifH/92RLOdguakppGip/0
dvtc9dbQk220oJtrme1XdNi7mc8i1720SVVAYkWarw0Z92yYRFvRrQtKNxipLnKw
G7LC6OiQzlA10sAFpeSVi3iiA7/D6gNEV/Up3AEc4snjQzfiGtTXHPFGTDV5B4Po
dZebflAFbSILM+ubSm+l4ppedN0wXmDFfvJwFsTWNJpsJKAY8usT/p2fQLFw02FJ
vHdZtBoJtvB7NtC6VzmXFWQ1pNHZcYQS4LChZYIUU1+GGM/zKCu6UiT7eIWU1rUm
NNob8ksP3lrTITht+dFMvXiz+uB2N+LOEEe4SVnGkOrmL9syh47iB1v/bthwD/4X
iSrlNaJY9qsGy8AjPot39iEJ/04N6gqDYfMDZLAg6Os0dV1nIG9c3ipleYWxxYQw
DS4a42rU5f5jwjDFcScIwtnVq5xWmp5zwWgOq4BYJcuDIfNwKyaGfqosR7fnibgx
J2cQ0Jstg9OU0cj3bac2HG7xouPBS5fx55+qIXx0Om8HVf0HS8zTkBpoI3wFagoy
PNkWRBsE8rSG3ukuD3313JU/sxUIcAHk1EvhqOZo7AICoZ/pU/R7X90lJCnaeYfg
xlDyuAHSo9g04fJWgD7xvZdvUtWYXxVNOeiZ6BlhIxc7tx5OQ5mnE0ETREQj+MTZ
Gt+73GMGSik5T9XkBoGjHjkBXUNkAqsbz+yjD6/EC6ZAkCWVrDJ2QFdeKj2gY1p3
pNus0KTxa3ZIJIQOxe3yV6T02+2doyJveTWo1zEbqZuKayPb5UK3rXwrv8vEEdPi
ArWXZwYdn9eFLA3XOvqdDdTyt2yLAcShSFZVH/aqruvXYQWSGusUf46FdA41YBTK
HZOwXlGaE9MU90ij0705uE2oJ+ZXTY2LYfEzr48PX4dF+qQiDr7m/wN6Ua0MDDK+
JytOe0JhPRdMBPVxq2M5PXEUn9WbR2hEGIDNUEzdll6uUTUl/xD9W0m00Fs0Jjd6
KkaEMjInXEP42hquoF+sw5ARTi9gdrM4h/yv3jJ3zYiHdK/SDaCjEU1lEF0tPccK
ZjD5esxm4e4ioBwKbmsS3/KUduQEzkGFfhatOQfjIWzqum7elx8QUZkVVdaJGEH7
DR3hTJLvqh8mA04PIdhNgaXHqg8ZHsQzzuTdCxNFVF1M0DcEcKdvKpr1VmDo4i8q
k20PPKlkLbSdvoPCbe/0Vc2ZyXnFHq2r11AEuDV6/I4yU9RmzHFsqJS4qb1AH46k
eke0cTdYxtciyuz/gat3Yy9ZxhII88POpja/h/q6NGLiHn3ZKtPVi6d5lYTo7DcN
I9kVJl+ImHvenDsCYyQBrTQSqkDEczAYP0OBSDZggx6qzuYDHJrRTQee5F52ciqI
HHxA4BfnjRSE/DAx5pUIg9PCXN+qYjdG+eoOnjuwLqsSEBjlO5owizFfAx2WF/lb
TbXa1p9W6Rb5ziFGiDX/2psWXeUH8dE9souoqLzh5uCldF2wgx2uR2/DFGJxH5Jm
vQGOCjWDspKbwj4QHY1fuEsLv5tIRt9EZwZMQ/s3Nb3NgDiRopPLSE8f83pBwMRU
2745lSYeF1CG6AaZMCm2m2tUbJFWvqqqkv/mPhQJIRZlECxrCGVmNFWlz0ZoAqH1
KocIxsXYhoaJk98MBY5K1HN1/rJtnoG5ul7YiC91DvsvfQxh5cah12ArdGS59EIE
Xst/7LiIqopACgSOd01ARP4++4Xrl+esehjPmFmTYejOjJCmqyM83NBKevHHq6hO
duMpH4xJQs/qA2z/KVDbFoRuLIuoYqf3lyp/gmEbrn0JSJXivBLyD9Im9kF1kvVb
E9sjvkAQ3fdEvSMsYd/pXalic7xvnF67l54DiE8PR0dVOgiGN/GOmqCjRaZPw5Si
SOw1oln54v0GftgxtOrnzPXN5niAtvtp/VPtkfIPqdGJN+NZzIlQMDvPLraV1s57
Un+pkUL/sAiJv5ZiwiEznYUBBN7WtnEL3vJCZa7GN4uufM8fQaahmdQUQb9ySq3M
WzIX1o/1n8jQ9+oNV/1LHIN8rZh1m2M19+beQ7Y5TexdERe3wKPC/kc7KZ8eqU/l
B8cxHCV5uU94Bj54MGHpxn6bf6qqjG2E+rxA6H+Yv+XwSL+5tShbk8m8ONgQTGD2
fS2tnyZSXHZusCl9iY9pROXCZEkHS9cKVddznoFpdwIaZRjvoJzNm0+05zYX6Vz6
mpCGjW7DHyvMarhUih3EXGHWc3mq9fr+j2+iO+mlI8X4eVWclzgxWXihJO8hO0KB
SQH18hRjP/E0ism8e2tcMdkvm8lfhEHkCe/BMu/mnsIZzWol31Q27kjfb5zUb2n4
PW6EmtcB9RFW+pwx4pcKLY1GLo0bgJ4Gbiurf4PR9rqct3FXu4a1Z9pQCH33I53R
pd5MPp36viH6rdC84pp4dLEeSeosXfPDd6WnrJZHOlL32CCpshUAI+ObX2wlnx7P
j6ZSgqcUZ6AK0n11Q1WywU+r80pgb1CBCpqk6tsfzVTZxpfjYCuVh4BV7sHmsaoL
HGxbPsu3bG8EHA+R9XEx1FlyNFhdBke/R5h2eNZFNdIQGGx/YqCAqGvujW9mdbiw
ReOyltqRMpfiUrIBD70RC1IurW1Lu+eFMJyPmmnRcMWrrHyUtKuKF5GoT1SLwaj0
FmKfjFFR6G7PU7Tyks8gdSaoGNQAXEYWd4tC3yEVeGJJZKD2WeAB0pqqQBYxPoCs
sbvrPWZXjyYn+sdqs8B9Bv12xPTQzGKFuhVjQCsAilT/ldXjg0wVcFeCgEEN6j6p
cuTbBeeI4m2W/ctjEyh0sapNi+Gosx2KPBiPm0We6iud19zLEX613BVW0AflEjQu
5vVNHScYGpTTnv42Y+7Toyk4ipGaIkK9jT5Q73rPVj5SOIzlt5gHPiARLcTLyiEf
d88zqpa/5BcmFSnh+eyl3575Y29M6NKfCULbtee/Yy0ikV3qYnYdrb8ZBi2I6s51
fBd9/anU9eBkMukpAdHIrfwXHcWJSl9fqm6LOfueT3x8Dqu3UdmGYw4I0bKJHZ/i
xDnMC0kt3yfddNcNzfjjJytZD2U1Gtl2zivXx6ELUjckY4KZj9Di4DO9hSZKuocl
8MFPnaRIBJz+1ERpPzlrBPw8RFeHl1QhSiips73FfCqnKV6jvZBvQdMlN4RMl01+
IJHLHIPE+OKPmzathAytE0ECzy1lOiaJ771BTl0ICE0pSgFgma1fcFyUxphSsnFO
3yjA3RZBQqcZR+6Lg3/boMKfNv1jw65zm7aLybSM2r1SFZoHaPSEIfpwlg2iVI6Z
D31+ZLttv5yhaYorNWiyDMizVTS6deZP4pok7lOvKDMn98h8nzUJi5e0gxRvpFYP
b5AufI+G1u5tUgtiK6NOZ2CvXPNNw+a51a01WDEyrvYFkrn0iw41c3IeOKYda1fc
z35mR/cIKph7u/nlpE6Ny6Sdl+Gj3YN6waPzthLWf+eC/6o+erB5IXLIEtmFfDNG
qGyLpLeCwPzjhkfW+4bE/6F5LXIo6NmyAJEtqQGfpTFw3qY9tYKC35d9Xq5MQ18N
HoaDzt2AdwHLSmQs/IoeAHsLUKEyaBHoh2cWMO0qNpYIgrcG0a8Ge8+130RpiTvK
wO59ZZPWZ0CJY67r4yxskW8vLZ4oLitUWjb2mN5di0enRUn6mOENa6YNGyn90Sze
KVZ94xKOIYiXZEpvEAxu5QXF45sgYkqNFbfPjGVlrUUBa23KAz9A9XF8nRHEH1pK
zKFOW6jJGSUR59Hq101SndWGYOTtSXGFXyLlw6GzKHQBM4zX2B5TsMdGNZ9/YZRD
G/VvlOXMX2vQ/pwSJWky+GAwZpZFVWolKMact7MHa3fHgIS/NSGr7vpeDNEV44v8
KoZrjSV8eMZHH7P14HYRn9ODKQupDtFlkXQser1a+i+byQ26BdrDr7BYKhePtiVA
sutXfBty6D1F0SlAsindr7khk3V3czBOnN7OhRLvC61davDUb3p/510UUUfJUDAk
HVT5ufm1tqt5z4Pi7Shuz5WMiWSlcsiBJS/afd8d86/UeI+9mhJ4cn2dokZstx8T
bSZzgvESngpswS6AJiwtTFggSBSMninMkVNE0YP57F8qkIvL+s3l4qLqxFrFz0jM
PW8pLpkhc4YVsRQOdX8MF6ariDBpf7zVlwmKN/Zko+fY6oIx+vSGC74Uybcu4EZY
GmIEmPJPxSX8S5M1DyXzhIMuJ7sKNgtGBu6n45bWQUvRcxyh1Ks2c1fhPfCR26TX
l6IfFQht7gg0ThPP6Y97kT7oQlHzBo94u+0d3xX/LlYaEC1rjyKjgQFgIQPp7YVy
VdBG6A85aUi14maZ9XJndD711CCqfAfWyvAV7Red4B0kZmPrkU2E+7Ag68xqZBRV
xxAIj5J4tkjMK8rRx4E88gftOrPZP+D02UKj5GC3xJemjYjEk9iXQfy1NcCHmDsK
aUZRNd1S1Nc5JPT0uSPfJBDZFAKDCOwZqdkcK8SA5oue3ZnCyCPs4eTgikfTvS8w
lOnICNKFQSZ6wkm32/K2nz/MOipT653kj00tmj2nvtXZMMQHEf/V9hAY1SxDTt3d
zlmfV6WSRZnEUt909pjZyXEEgS2MgSaw0pywI2UDPuv2pTHAGWPsH0iQU1cmy4Hw
2C6y+MZnLoj+PlQ/1YRAjDZdeanIXWmfD31meN4dC0Nt9MjrcYXZGZ5KZQ4Jrf5v
miTWW1gXTNCgEXDm763i8lHS7UmL3LSGeJckYRBoYVgD5IouqwUDYrdhASSGH+aX
MY6ybEIiaS8TEb79Z4oT+VF/PjOq9oSTY0xzJPoE6bmNGkNTnQZrUQZDeFCuPo8Q
uhU/dVYUvKb4JHjg4wUjXkVoilNo16E/ba2+afNe5y96NdFfCPXOXFP6RkV0Up1S
46eqQbCDG01TtK67TgqzKED7DqfFcSi2OEXES78AasLeVpU5JcUrJ2kPlAgOtSql
ZLC+tC1RY3ariE3XhtvPCXhb8OXCsY2Hu//lbX3YNRdmwWJFpJT8ugW3GjRpUqYs
YC2W9Asg/ND1qxT5vx/bkFYSjOmO7Z5xIXmwP8KrrWk3QmnvuN7ZN4oxz02j7DSM
0ENYQk3AQPxZZ85VwpQRXQPSJYibpyFbJZl3fKTWIyMBWfUyC2z+UYvp6DpXFLsr
siFN9ctRX0JoA/DBEwOIeLr5OnM6tKS9z/h1DkhgqkwXn2CAugMI0UugQ4vqHYqY
Jl0Axbm8rMWpxwMGx5ZxtMRrQcoVHdTglm5CNBdrOoefLG/IBOcfWBqK4S0vVOIR
YRZHb0TiPBUd7wtQNgQxWynYL4cDsdF355ZFZcQXfwP183hmaqsbF8E60C0NhMjK
msc/nhsjGQ10pvxFlv7fvi/hpZQKpxHM/WDJvjSEq695KqNdJBYQWCfFUI5OauJ6
YZGjUCrGj34z5TLS4Mc2yM2E4ncHgLWZVqAxfuf8bu18mmeDi1B7CutvgaEfR8qY
Q1gdFfcsESEA7hEgJNX2KeFgobGyAEjfVyXXkesojsq6xe3f8tpHbBUxxq2Fsoo0
56wh078ub/vRITnFyQB0kHf7RZHnymeYoqfOBbBOSRpCoAihooo0UBvsVo4Y6/BX
HmDAUmgHMUp66m+HxgRCySuwO78ObgzWWfkLqIH3VNHp43fY0BOiouvFtk8U1JTc
6kDMYjJM6CaVMxlfNkjq1Ea1x5IIYgUQzxzKg+QeFSH3DOKGivoViJfU9NMEYgw6
Ac2LdgREkNeujBDfd0NBJdRaWkw+FXBTNpZZTdP8JN9sTiAr6g5qGUr9+fKo2KCB
IZuoNtMzoqsser0GL9eJu42C8l82baAbBwicIyYi8lXDh8q4LLv6xnJYXVkz5qyy
cYfhSlaH40hf2CuocDpWL62cmhNk/YSGmRhTrPwS9dU52BludAnSUe8eWl+CRYwH
y8cdjNblAi/ynIU7fkOIJckO0DKK6WkZSNfWnikDewh3SmbRp1Ez4/fa6evRCz5k
8RVND6oRneWBeqobftiVfMGMtAg4fFPvtIOj9DBgTVRkBbuajeSwkd5gKii2nC0x
0m4UJ3aA5LYsloRdHlEeXIYvleGxodrGlcG6ptl54bYMN3Rev9D2f36uVjt3iF2S
6kEQRjedP7CdO/riakdjffhiMpk4oxXfbPbjAp4Xjl0unnPir7qNaPwfhEuVHb+y
RUGEjOdIselU0MId0c7KWkzVTXbIJfB/g8/zEIH5gbpKx3pPu/mRU1PFbmMHYRs8
8TUnMLzMYGiE7AZHFN4jdG2A/3cnyTmglJvx1lH/MvmNPznrKD0eQE+mj/QNsUTI
rnJW9ECv1o4Nz5SUnanUVP+WdTJAz5jZUURZ65r5416pb6FDGnnwfh/Ej9RpepOW
JXqvkojVd8LBObdvlOzY7W51ApNSa5I+HUZrueffDEDN1CsaY6URBk1oDfx62dvT
dn+JXfnzLLk9AdCFSERMDKyI0AWuUlcDYEboIq80unonFCnnj/w5jXKo5g3w+ziR
wZVGsylJgSHgZZQ+c+ERppn0DoCTzCJ71c/GC1PLrV3EcUodSNkd26/evd4IVTLl
kLd/OJCugdMDL1PJNg/z3WTzBbO7HGCmCRhu5V+q2WFBR3QHv+NUH8W1812D4kKn
nQoNXWZNJb8YfrA64dZe2hdv9ZKcw1CZA36A1L/T0GSkQQa30Rd03iLWM0jAbtxM
CfAmoZcNNO262r8WUjB1n+hrw8Kl79lO0V26C8bVs3ZKyBR1m/DSj0auLq58Xhcd
Wx+c6Bi0AD8dcr2qb9YYhjVYF2f1UlVLApLR9XgOESg6v47M4xAHqxEFyxrtUekZ
diiptBlsbBoTSWlzkY5YhdPseH8wueZBqcSRq7qXqzmzZnSCX1xdSJK9j700MKLh
HyzTmw8FUzmDeWcO3NxCZKaXqGSfimLyA2nh60gbv97Y0ES7TtdEct8VGq/OivkM
9pj/VwMVJn2K7dXGrLN4u14ruNWOi0HdlPlM6X+oDA6T+kAKIDEreKwXl9HKszaE
YMbzXfdXBxgVyO1LZJKmFRjDgKYQmanglHKfwGqMmX7kUzLINOI4wA8BqVQrZjST
Qw1vCaAlZEd7iImKL3kWF7IndETsXVwPiaMEoebpfVdcawUT7MWtKT6oirjLKPeB
4G8aeAhJ3/2JRJbyO3SGME50NjdoZGUXamfj9zdEg7qnloeEDCd9uMekyWM0Ni3Z
0sBPT6dQUPUPFDgYfsDyjvhl2mjxOrd250+fBhuNQp0+pTDws9ElaD3+nrlNy8M3
E94uCaCPLa9n2yZ9mS9LYCSwVxd1a36uEA4oNVZ8tP3VIzaQrtIk6kNtXMwgPaQw
acva/OKU3r3mqf9Mj+598Fwv/GxWK4fMPrT8+FJ67wogtHUviqIpX9DgIaB6oS/g
e4k6BvJDjhF52fTIYVpJeCA61lf+r4ieqrVwXKhaq1P1wJrVZ4JwJpXt5BzoXr9l
h+sR+E8fLdXV7JcMGSd0N1yh9bt2JD4bsxJ8i0vj7jeVT/0+nC3/Boa4tu4LxZ+Q
2Zfa14ZDSFtBmuNWkUE1ddbw/+CHq6Emco3ZymcLu9RwDBesYbaIVQp6eHvPBquh
CcIW48vMMpY4OCwqbmYvzP6CcAdqL+0/R/q1hE+drFAENSC0+54UIflTmAmmbBpS
MYpfPgCcx4ny8toKmVHfjbQjjxLwUpgYPNh0xfxdZEeqFKdh2ci/P6D73R7FNlPD
CGcGVNjKgL7qF/gIJoIbTivKfPWfMazEboSAJCPHHU+IQo1qgV54UAmwS94aEHO4
shXmFb8B0Fmdv+jRv5gwWuqtaTmew58KAiMkOaf5/RThbRnAwqnSEs2zE/uACOXc
8WdhIBGrZr0M+o+fqsNPxu16k6zBh1dCRvXxf5RM1VGGXq6hbVJvyWZXLePgS7yu
iiyQ2cKLovYafPmcXZtMfo9cMQmGYNwPev0LVL3hgH8vBRptZpgRXiUP5Yqku7D7
V8kSsfGWvsmmuedyzmrAa/5aS67v52trQy/a3x1uYquzDiDdVaaswOIKDiHROJxj
OxMNZPiYiXLUD39bxpbmfAix9SbNfs0Aa1tzpj0dHNno35Xqiz3T47GJZG/HZyGf
clbfH6QzBKk5Qgk0fIVBaEKL2nxhiE5CRw/s8GmSugjsMQeuPHEFq7pyF1YCA432
80+Zjqb6bfVxKDupvcBcRq1jS3JAmB0QVRyN2r9UaW2bfOBjMdoYJMNhGb4zYeLt
REk5y4OAVRbrUzli71n2bBAlZZObiOjAaN9dl9nfY/SfjKyrXenHENVjoA5N7HMg
+Nm0oIxGhM/FLREWK5xZytU7Qxi/i9zOK7KxLnCkxf8xQzcn6cXWx3NSlmC8K30R
BkEicU4pO5a2wAneilPMQsuJb6JIU4WWKWZ7wVcPtcL6DM2BDPhlR1T8Thc9D33A
L7QgllIJvzGksO84FfB3HRZeFKlKbANtPL1wQHzYqjSno8N0Fsh4mQBzlAp3ik1Q
ZWjdzhFO1Oo4OAG9Dh0WHfbrV0uumRncsWiUWCInsMKVq66/yz7pf//ynHJI9P6a
ogz1kWIGzjv7m5osHmhhPmrAtj/VVfkcbwkCjdrtgy+weNpLUG2NjaiH8+RFw149
MaUMa2gKmE46zmh5EW+pzdDz1qg4B1US6xLN4oaYiAs7ZqPgb9FlqER99b1s6REz
1lUy3RjsIeXRKOBXbVg7t4cn4gxDmxSyJf9eiWDWhoQbpvmZjQVsLcp98SNRR2zZ
zTmoCTPzOo9sMPcWZZobZ3Pgy4/z1qu/TuBIMb8RgnU/orhGmLF5CmaFI/a6jzjF
kUszEPVMUD6NjH5uO0GP153B0eYuo6+iqPKZJlurxO2zKQ5YlcrafRUFeGn0h8YR
FlDPDAgnm4+NsiFmXq91MLnDN6A79Sktf4y2+Joea9NGVi1g+lG47EKlGdSf9+Tf
9rlbzIIsgaFCfS877TfLRUiJF8wyCkIFOBq3vlEEgVtJkHJUJKreJBY0ArTazyM5
M9xZrX5YeaGgpUGqYDE08b7Ww5Vn4S3ccyEiIYrk8CwSBIXs8Ba5bAvN81hhUOE4
BYK4kpcz2/GDlD8h92dRVIPNj5hpAio8M9Ay6k6W6oRuntiV4nLOdu6aFbynxss5
2B1y8Vr6y3yfDBom7hCoDUGqCw/sYBL6+zz1y6JdNJkUTcNa46cBQMKlZoHKw1qy
C0Ne2Tnf//VUTOp0DtQXPzL1kJi4RejBsIC30w0mfmcdkXPp1SEUIJw5L6y3NU7Q
ZSkwohhhvKUOE8zXjgxhqPR5FWBoouDV+6AnTaoUZCyx7M5KkmY9bZGukT8jHoSC
PbOfArWhAUx4QYi7L/o9tSo3n+HkpOR6zuARG2ZqQDOEQuyPZUNH7iKbMuakAPV5
CWFcQk16AYv+6yhtr7fZGg11IcmI2jpShesPshBsViL9kw/wlZN6kTC+gJFDYtiO
YATcxhDLoZZIlalweGdxp4yK34oRwLRtXwQPIQOJ6L0WWtXc7CkpRK+HJUTRv3AJ
FzQfC55v/R6EfPJE/ASA4EwAm/PvtiQjKN/WVdshMha7iFlWsnHH6Zwwg1BoLsVC
VhFLs5j9Y0vcHBerDZoM+WB+FTWSxVDqaHRb2+Wu+OxwWBfopvp12eFqROHWkHCn
oxXe3CA4fA2oPdneaNJyFWL645KS+EPy+btxE/tmaOITMqxFmktTlHCB5PD73pyK
u4kplPLXS0t8mls4wK92Pmn6B0gWq8yyQa5uVCgs0cPINbxp2574/3envcyyeaDk
3TRFJOIgjj3yQzLRD6DdfVwh2JZFgt1YPoPrnqqdGD588TiZsKEFK0VWoMzeTHM3
PaU2Ep1Hs6sjzgMoSpcXSCYXdF+QmbJ+psH3XoE4H1CsG4F7grvqyql/ZaQ5EEvd
2KxnIqrxsZOQOg9B37DeQsCeQJ2hS1+8PhYwxxUZblQ8kUQ2ggdDyIp6EVIF8o9+
P8NOWpoqjMXvy0j8+r2UDkkJJqcmplMh55twj0fiD20/4d7YjUPpclSFWefua5Qw
tv0tkDyh0ia8d3763gwAE/k+0idaSFU+B4lpxj8hbPRJLaxPAOPWadLqsyg9QcGi
ruw0NitZ3/tN6hjy1yM3rJivSaX+NJgNaQepaquqGfvNkPUAdmmLxs7FqMabun0P
3/csm076AW4ZfFL3YVXH/stNzDq+tcT9NkP8FVTXTwsRLvghRQn0XJ6rxQNoF3Bx
V7kEyjd982EYeuahyP1gPR47unLzvXV3u3jofPk6M8YIKANLeqC03AmNgNGoBXQA
PeuQ+5NM3q4m0dz8TUowHZmgFFMVbh+2iiVQGUGBrPsPGvHRnpHI5bW+bNgwWDaf
tbluyS/lhDpYupAkuyN+KdJY8UjeKU2gzuoptbiJgVc2d7nk4R5UmZSzvq4df0bM
TjCn9e+wXXX53b1DTEcRXF5GLrhTKcJpNMrUvoHZHl+nHK7XhyEmjs+iCrZ5DsfC
lBdqZKrVu1rsj5275IzIRrkraQyy3A7Fdyave/yKqdhFWf9HfxQrvVNMtpzH6lYC
EZP/S1oKPzVE9fnSKVQAYKvVmFSmNiOPhFMkF/+IRjNRwCq5nt5KHYdQxEiU97m0
wdOu+K6hMbE7NLIKl+BgWP6rUEj/K3YsYjBlT+zdt2I6UAJbMcIx0hVbJvbziSzS
r8FWGIw+I3/4p92K8ZaQnM5JfvUb/ndxIY17D83x5dNEsLj6TE7wBi+shzdmgUsP
To870yAK5AsTugojgkpOWwQCGW3GR2yL9uGOt48ZMCcShqLRP6vCXB591TUtch8w
RRpwmNkWxxOEYFh/ClGTOK/YbC+89n8h84VKTuoELcvgnJ0FjVJjKIttC7aSEUm2
idfKHkDWwThaWou+bpkW1NLBIptol3EFqlq2DGyahc885Hp8CjJ3gyoyZmiwjIH3
OtHx7H58QGDzNgDpWLafnCY4xiCuMfhafsPTvS8hB1HZp9B/wBDCyzxdZNTCz09Y
3tTZJqnsiTQRVC/8WOPl5Si2AqQoGoUdz04dMDkAJjxginj+T97tuqZ4grvGR7nW
cN8secPGVNyt7k96KaPTtNrCKe8mZOLG7CH5gmw/vebB7fV4Vhbu/93VwoSiXQJa
T5MqCPxyI3Uyti9EZVePeSpB6/L3I7v1zz2EliaUQLhTpXmXIlXEiVKDyNrR8UZU
++w95fJMc+7jQhYo/m+rlYAYRPbYNAjzdwZfnhU7/l9nKmXdaF59facV6qpM5C3t
4t35Id3UBcmVBJSlO6MBMzbYHVfmeTsWZ69o/0B8mOTthss1ezDI20Ij0tT9ZQMe
mzWWL9divI6vEJWpOUI3KF0JsGcKOzhS0qyeTDeCLpPPh7s9JeQzUGWTGTFhl4Db
q7Wfdtuj3CMWbKVm9xz9JsCbbPwrYFD53ntD4CV8fZTmDNFnFr7Hudo2+SF0F4lo
MGwxnB+e7Kf9bWvVHtA/mh1caO3/UMUS73AZR7aEJkSFtuVo+YoEIX0W+2pS/y+H
6WMbQ4ww0QsWBUmfBK7Y5l/eLM72u4mtaijhLNqAqFeuwmikDX7P+yutsrwpvxhx
fbh7zyz08mF4RFwyJn+5be4f9AKEJvPSPhi14ZukuDjvzeZ9CUMq+1QgR13wELNi
lotVOxvzWQVTrz906nC3vCDAYoLxJZl+YU04UrRUcK0p59bUxRw+QlOs2RlDuqyo
b5/v39klAVQewXQ12dr3u3HMiYoPXJvrJGnJeA0XygfWwUHKbmPXQCdLm8fKq2Pa
KAII2+jPBU29Hb6fPOh7KLj5ci4MD8z5FAci2SKgjIQnNwPzxoxhH4JB0r/fQ9H2
YLOMrb5BWv9VCPUIu7UlWoPzz/T6ASXzpW96mCgT923qRXviaYtWdF9huoaoXlqN
3QVhiGWSYevu70hJjuIpqUV5eRl+X35hwij1xz/aaXuhaV04Uw/3MaSKXSGzwyl8
Dki1olRlbBlDxkmDHoS3VlnWq+Z3wJC4M72qrVERjoaagRbe6ULmT2oMcFcoLnel
kVJXS7oZCD63mVqb7V5vQWSFC4DCM8ANRjLT+rzDP9ZhwxA1zL6KxkXFWfVxg9W8
VPoJtTUdZX79LsqI7db6I1h+/MKCQJHGDgosyBgwf/C+WJ5MCYuzwQlbVjLQv4Xg
zrba4Z1fkYfn94mUvKRmFpIaqXCv6CMBVSXezOkcDW8ARHVAU7eSu52bCdIG3KNM
HFBhT5Gfud4vjrEHsylnqbmEQJuKdKfxr+ZAvQo4jNmuRTifbUrr6nBc7kN7EQN1
4wUNH4HBkV7Ytk0uogXsllFnjBJxkSTYI/H7mocqw1+ObvX1UZ4JcMqaZTcpes6P
fPHwd2oep/hy5xRaKc3MN+rWFJlj8S1O11OoTg6iecJKAtLhTDMZwQc5fZeQmHEq
MyPhCTVpvKbnvPKZSGbsZd9bpRlSnO9rU6AUA/lhP77MzgU11lUCHr6K7ZeEZoTb
0y7t2NS4e3Gv+tu0DtWdAEyqd9pgOBpQZ+5MWzecV5YOvzXmAVwyalSpbIf5e7Kl
bi5uzmh6gw7U0QUVU76p60lNO44kwWJtHRFJqhGXDE0HiCFUJuV7fzQLP9ALyP8M
fWM6OOCNmJuFxnMW/jTCFHk++HK58RGwc/B5v8akAX67r1xlBS1clmSiN2AQoiVl
vFnOOpJi55PFoU25pRduKhBe3ub7X/176uHF9WYFxGDyEsPWdkYSMbz57i22p6Xd
bgeYk6sseYPq24hsKDKV9qdjqJzpYC4BtF5SKdNs5eHtQ04HdCR/kFCix9QFVuEl
1Ghh2IhntRLbhT54F2JPIyrYqiqRPZeLr5fmtglFOLR3gBitZ592hMkAkndBq9mf
T3AdgxCgRxzv9kaOkYH3Qt6A1HlZaWnB2jPIrLFd3t9OPqPjP490iihCaOEw5fkI
pPSRCi66T3zcdiIKs9IHxk0S3pOYVR9icmWp+ATvwiqGeKg1IN4ZVrHIHniVTokB
bur84eLcZ6AgvtGGPHvp5PU3Om5l394RKLIbTCPrWzf5qsxSfKGNdescaTac2LOX
ZFVXFPpMokpPnspQgp9fH9FT3QUiiz/kg1Eb23DR/9DOvX7vi72esZs3SxPCg8GN
EqMZ03yXX+Vi6ELc2kcw4TtwMuJmma0E+FGU+JBjElR2VUt6JCltbX7VXi+gnTi4
rQCQ6VzCecgv8epydq4O8nrOTe7nifM6Jhqh/V+xHB5TBsEJoNIR/0etVr5GEOEg
ApW3zc7nwyrnIpjm2gSoyOEPCoHugGtx/JCtV1UQNGg62vzLSODONG5BNJCvHfRv
gDFUl1k+Nz6D/qcq0zXp/aRqzdhES9EpniUnXhNleKEULMsX6BnHM7FhR1sWBxpc
6/2XQ9uUm1nNCOhqpsYrytqBpDYNz97tcANNlvWghSK7CGB8ClIjG41VTL+6XW2I
rOkOjZIwSEF1WViyBfuyDUk1+zlqepqFEgIu1F1EvK2IvtvXUqpbQGE0xpKMy5pk
Ye+CqUvdt2jit+TMTSjlN1HoWHoSDlsioj4W/MR00LRWkrmIQJXXCmTSYnnTWnbL
VBNbR/KWGL31Q4h+mddYhh+Bv7vaNMKVGXCE7xsg6yIJuyZzH8CQ3luUFL3ZaQlw
QrMz3NZ61zXBPLgSSWJmAPxX0V69t5czh3abS+oKZeXFXeCRmK4b8LGACONjUCVH
TIhYTblSWEXswKoZhrtqoRLT0MmUuzCzQ8pQhjhc/Pg1VpHj+iayPjXDAh7DTVt5
BVpPfKk9C3PEL44H9sixOXvTpz7EPaDaBwmUEyq/Spf0Zqmq3s6OzFW5I9FrbxiF
HlAHnymnNxuOyL5137l8dHH4mdprNUvJ/UbxjuspxOAQ7eq+5CTzIE3iey5z9Qwf
TSsDIxnbVFnc6HycCq8/uuNKmq5tTiHOazqFqviuy96HqmRX6j8uw73SJjXUj4u5
W1311aC5nCRVB2BtERQDqeXg5LQ/56UnX8JPfDsKdHZSb23qqorD0KHavCPYMj3Q
9mtSsL3GiFjj3gVntplsgk2NNkGuqcVDN5yF13tfw/OsLcl9L7ody0RFdLSyDhFb
5caaCTXezOA9YFoalCQ4HY+aOJM6E254DA/82SXRdpXNvEo/EcVDpX9BqjJRgjx2
4hVZL6jDydlddoxAwK89ThG0HGi/a9FqsAtFUajSlaKDq49ZNlMxxprCm87MrrLX
d/XFi9jqelss5YN4V8dk5RD3QrOSsoeNsB2LokyElmMVtAMHJQbglfQ3FjPL/dau
xG/gvLCt7+SQGgD+rUDP++h3pr2z3U6geGDPVWOZMK2yLXvyWM0iqNxp1rDJ8KbP
i/BHYjNXvGQlcNCK08bbOm7bCqj3neI+viIcubqC20pZvsU35f+MPmd+FpJ5UEov
Y0AhEH8w4Plh7D8i+1zQC4+mhAyXrvTMKFbCukSn4O4ikBxQiljG/vVwtXf3+a+/
b78fHW5jQ9nqJ2yQj9UUpya4vmaSfPUR3KX4O/P+SOHep+VIT3fJAhZoJE7Kkpd+
4A2sEHMECO6Ntr20pgQ3qNehhEm1U1EbM34vp33wf8QRqADskMQp8VnW5L21S8o8
RT4aGS4Yc5d4LBcECP0W217dGclZadk3BqmoGMiCfGS/Uv69UrZ850XramGdsrUQ
e45ZRo6k6VEJdpWUMet9A7seO0fk2gSu0y2BjsHo85u4e5hxWmxz9Wan6LqozsOz
1R2TPXn8ZRGy3KHNHN/60aflTacH1TmOEUM5JtWaHIWDhuLtY0/uXvVx0+igrAYT
4Lkk0dCyIGXNCZ9nMufTcIvvsHo8+tkjSVWpIXH8snLx+fXzkk9xvkNloGybjqKn
z3+4ZAfeqMhSz/sYo7/Um87+ZiYs4RlOyUmie6zfoDjqyDSHSwtvnRD69MM6MZ2K
DMUBk7lLdS+XmQQ2Rf8CRdZ/hUXKo834MJrw8Oa2LmqHHxdiqPIw9P/59JWHZGgm
EI6+98GQ70+S8WmiKrLSaYUi52vA2nBMor9oQElTIlzLkOS287U1RLvW/q53ZFj8
o/YjuogHybA5iyd/78p+1MCdDz+r3YGDAw61dIejPfun4y+goQOPtqt65rPHKUx6
ssSild5CZ46W4zSqyGmOgWATWXhz+wCJN+fWbq74J4IQUq9r2Ksi3bHh38TtBM1a
Z8nyLgB/8P/3T7HsRRWU7zfA7hMYbEO57zfhbbPByfEBnmZcCdGB9qe/mreMJXDt
QNUCkOyGkF2zvnSXM//dtWvyLyDXOlI5VewW0pR0ERqxFZOMJEeOmnzl1cW/Jphy
R6rjerqS4tiWvsNsFxawkG0RfITAlZgNQ9bb7PC+JPaDMYyLD79t/7fJSzW1DAy/
LEo51AZOlvqbmOFU97EY2k2qLWus03UmtSE/15OxfJYMZ1JmypMJUzEZN3oROu0k
5T4HQhf0Nit6hgmQsJpQR/h8+ypK0LTutowLdFf6gpJRz9bfQHBi9sHOs1z/Y0XP
6UxDL8rkKBN8vUIC4h5N4X4V3MCyHo1R5NDQmI2PEc8rBZ8HEE2wXntCOixMS7Ok
GeCl7TUeaKfxI0a4OXOdVt0gAODRq4+L0rast6KFfnls0jUL8AnqEmHUzaY+/gkD
kOhTLSE+Pfp3DYsV8iCkg7e4154EWwvHeTZ2gglhCIi1wJHERy96Bfpa24oxweZP
ZS6d4p5AqfBv6GHNaFfjTcelZ96ZFcpMHcGG4kaXXojEDN3yrkxIrghXE4wn731Y
BaqsvnC3Gt4I3A36D4gv0n3Kz6GO9HXw8qN9y9FRAe0a7rsXi1d1Nro9UB5J/fMp
rqXAnBU2V4uJVIEbDUDpdhq+sXxZo22zNxfCqx5UhhV3GjhwFsdm5wRxpPIN8fTD
8Aj3rPmPAaox8Q8zjrgx2WbTHCxnmC1J6DHNe9pv4ap+Bror1wtDHZfhfLXheie3
QaI8HzDOq/4C4brWLo4cl7hPZxhcUNq23QtxMXdaYcEj9VKH6IIa4+6aSAvRjWGH
TZnUmfdtnzhhxK3KGhwCmBHpAMJJ8Dbyr2RKYRibq5s//tsS0HerS/X3CdaBWmMT
usKiSDLCkQCWsxc9/zM5uavh+EPiMpHvEIp3iiblYwgSy5Za8LT6Y5zM/560XnO7
FjSmR15PNGqdRjOdS0cOR3kuCR0IqyvT/Tz1+DcyfP2thOoSA35aoVGUpHjZ8cKd
AqULnWWDZ9AAkYtOuxsy23bTcbTBpPQnnUVFQMD3Wj2TQBb4zjnFt/eLo/c8wa/j
PvUG1jrML+OkkcUuWlAOTdlmi5jYYTNcqmAXvJSeaP9z6kmm1YUinNqgYiIRcLNy
R/SNP6ihCzVGjwZfBZq79N9vJUOKnQ02ZQV2pDAyPiplVD6vmy5VVDUblUUiIbfB
APw8eL6tFaW1Ji6gm9VFRgbCte1kVdpiHatA7uprJmZZLYXMJhxHtMHd6VBxN7II
byd9MQ6P8CHt+ryjs+N/WqVhKFMQRtJ+85k4ZhWbbyhXWUc8sQXwqxvX4NaiZelB
bFhMu17gYkRdcPzZs/mDIfQu8eOMfD9TQEVxC9/oNgiH/5YpHMsptXF1a/A2t0hg
ZEkgwJ2ModudBe6XWTtuSNPX5daRZ9Q97njZxf6r17KTOAiUzI8uX7Te7NyzWSLl
Xx3+Kg5wECXfmZPSdFw/0JNCsBgFkX4EfzQi0pjSBiIR46lkmcoK3+/2e1jtjfNf
UoiJdZ2EaXLFrf9IDdaHk/wLSJC6pHb4x4p9QEqKs5gI7TbjIWt5LrqZ70IlGz/L
FtnHgFvc0lv2RXh/tMbGiBgbVhqlVplD9CGB5yXC2e+NbWky2We4b1uIAybRFCKb
MJlbrShwXXCLAmW8JFjoiz0z5wGGLtcxN3A7+RH8qJ8FJr8JDsvT709ZUV48SrfI
omJyvO75oFpw/BlMtdaNOUYGyZwCLzJaFdTw/2bNLWlasvKKvtKZ9zST6PAS7CGp
MeRzKVc+xf+mpTkg/gxk9M5j5rxOA+sZ/Llc/VDXEq1k//eWbCGy+0aS4OXmkhoM
os1UAllw9HjR6rH+2NgoSES3LFCNtnxdhRO6xb3jghNBb3SaOG58bXgI8u0Wz3cY
SnHZJK3UbUb13pd1RbL/+gvIk9p/uJ0y0CkQPLGBwE5XdcQ/R+OhvZ5TEnuxt+r4
gKRs7MWCA+1PrHXd/EzkgfqK3FxSGBYTSkx/2yNmpwUUYTTn5K7htDWI9yNAYUfr
98dU+fN+uy4lQndoPDAkXCphAQsoEKqOx2T3DtSgB3ojP0M9GE5E0ts3cIsjxpJF
zF6mYdg8YTqX5tBO+AGCiu43K9xL+/AuRJc8l0A7B88brUNccSiFdStwTOSTWTem
A99xLoLi9Um4Bo9J9OJxy2JxAGSwJf0iy5frIIARJDSh1VRxyBho3Ru+W/+tkutf
BWf2uQ2/6JZaBy2fYl3+GaZJZw7UMjJoLEoRXCjMdz9WErbpjDaMRKreACijDcVn
5jZ3wtVOx5WSaLhUchabHhkZsgz1/vdc/XrPkppWCzEoIs7UesmKw0Y1jeQmTQou
jMrecFISsI4WjAlidJCLHkN/DLAMdGrrm2w9dAKwE95sRhiKR9z7rYhzYLGYxZNl
tgTqgzRNrQtyAiUlds6Gvl7SF4vh8UVvimty5swFMe7LahWc+Nm4fhigTy/ZTbKo
AZxQskGCzv/Fyws4ZM+yGneXWatv5+opfMXWsOCu4QueJrnfUwWb0xnswMouH51v
mCgX0/i/YDMvF6+G6wWxD/WVQ6rHO9OrfSkEozJqCpZMuuY3pwLtrjFdq7wXibi4
XYPfcSQ+A+w44VJoNjheqNHT2MON7nott1/ksmnc64gwrNwbnn5vaJMXUfQLUOWJ
PWPLh6cAE4r5hIlLMk4FCioRpUZwXBcJWCMf/Nn3D+A/PgJHAutSxrkWRn7Pkd7J
O0TLp2Dtz8ItdfGh9VCUeiuDB/lBALFvgliGL+L1o2PnPhUh33au8XNS3nuvTYn0
VDbtaKAiOK0BztrZteoEiQJGU4oKjeFzc2/ctmlCGABOEmHZQMD0sFwEl7W/K34F
bV+JifyWqSbLGPL8CvAMoA5R4X4Ssv9RnUkToHI8YI7NUwYTYtrlggYpyvjoq5TM
IA0RTct0g2ZZBUzQ4EqgTBpEJRnZ99k3ZSKHabAwTJRAO9YZB2AAVWffD2MPxFqs
hTqRDySfEPLS4kLlv6czlUPWwTy2WP6s0RJIUQt2dmke+I2PzHFwScCBKBav++gR
T3nfNPPgiphqy9w+I3nTXSDR3zEO2Ak279F8msrQ2/2uJRq1rTtl9Hc9qR1GgAF7
0s0yaVPEbGTwUkxf/5uQygsZEQ1AjlAaTUXXMdCgUau/eWOQaZ9dd6QhfcuIwvWd
oA+vRtaN+1E7sukQl4erJneU0J9k45HVhlJjcdwgHE8aJzQsAne6Bu5ZIzY00MXU
3MURYcc98I7JXRCLoQxrcv0I7sbfGFa8QBjpmEWFS+m5W2xMMYGNRn+YTjyCP7WZ
KD5WT5uhcXM0lFwfP4z2CEcs2Xoh+NfsIvkWT2xbAx4CmRg+I99CkItGfASnnrKf
KL9EjBykcfd3gJJCG7uS9YWoc/Hf5RkwHRDdxsjoSsopY2vAN3b6yoEpV4ZfFMYs
1yUi06IHElg8GOBttSgr05gCjwdwbQws+oTQXAb6f9zb9RMurcaVWAvviiItoqqR
+icEg3+eI6M29Ix5Z7p7s5+ATnmBJfEIKTiK3ir7bSuozFlPZmRJKRpPwi0xuomX
8a/H1E+Bmeh1MF9ijX1vfCjCbCJU38PI6dJO3CVKlA6lJt2CZID7+UB5+SFPmxNu
gKmWi4BO1d60F/4e/SX+fUPPvaSQLQ7VUi/0phMEhauLlFeYbj++6Ye1g/ORyOPG
moUdtYMHDd+pq7RyxjcqeeqoVDnJfX4V+WA0ZB5ElC1dd//802480bgfnZ4QDguS
adPqLZuXKZGR3vDIIMBH5+/kGyofAG+aTafSCPNSm9sR/0hX5pJyOgEdxpNnR64j
VDxwn7wBQznpFa+GH9j+100slxyMHgvbnaQQnOzsW0wegPlr8NCOO2HswTbB0DNo
vXiw8n40MspSJMddlNMBJSwk4ycBfbpjABHwHMeD0xZH3hw7s4TaDobLRwUikDK0
Din0GjLqp5rBoDn6hZjoWa8NAZI1B7LInLS9PIFRtrc67+09FKWJhUnt/3BcJT/s
xUw72XI73qlLftTxrsQfLw97TrgjVuPgb8llLQjW99TJzvJZ88mnp3KntRN7fyl3
hCaQONunS7v3Wi1Pz6K0tmYleyTKp4qoodBYi5SJfp/wcgnIEK6FIV/lRm6FZnV4
Pzd75YBFgVaXrShByqqIIFslyYpeQDEpkuWYb8Ovy3qYYxJyvAQ7n1Wr7l6WMZGe
QXlmeB80VP+hykveF/LUQhs6k69/HRYp2xB2mxzyg0k4EMzmjbBmc84u3fJZIvpP
jufZ10v+Dy+nAnquIhr/MQrlbODeJdrOSRMWU3OEoid19+KdlMsviIDbdqZt1XdQ
Q7ytDlGEeSaTEqmDHpadCpXqZoP56sIU/ZnE4kBVY9g+rpS1EI5JtmfWEs3rx/3n
SGxcLd08+zUP6RohIuLnlI/xb58RQYX8ltPq30RFd4nAkJ7yUrDpZDIBPSRnUi9A
gOgDk7rooUShZdBETmqu3uF9wYgaR2DS+MNtzjjOpv5ZmGsFNeEMz6o92TErJjd8
vczgbb0RNJ6R6UsQzcZiz/2kUgmCM2pmbznHZK58pvQQL96S7qTa4MrdS7rGBnqY
xX7c3mxSd5ajg8JESQrANCoPx52hHgiDzQfn5E1NVKwq4e3UGuftUPDrEtYnc5MO
F73nIiQp/axhrn0WMd8C9fukdBbkVWt0tTYAe+9IhxXKNboVK9Wu9ApIauMO6t+X
8h4F0o9O+i9XKL6RvXe8c0W05XjnioHcxg++Ii9S7zvI+hlqyND6FF7oCkkwCaP5
G0BR2PPqvMLL16Okc7/Wx76COY2wZRb58/QU2arjRoQ3TnExgC3wVI0+Ev00RY/8
cSdngvVIjD89OrlgT18yflEJdi24wULHdkolcpGbrMmI4Cgar7urQ8tMNUZyGRw4
+/l/OPagEHJYhfTi27lMbjEkWearprD+60F7avJdVkp6GlbT135YkwYrUubNIpG0
JoeMvnpB6nFPdHKV3PiT483YlDlIywzjB2YIRUKJSaqC+j0isocGvSN5gc/AgCw2
KxCLPKjhU83TzTGJ+rStAPY6rf5fF+L9WsJdvAmCwhIZPH0O3AE2kFgC5/oBUHNM
uhVR6+XK3hEX/JU6jRjVBA8sUplChKi5oGRJLTta3iLkAx3w9odl8jAXmtV/Qurh
RqCfiFenjABG8O1xRkosa1SHJ15b8xoxdFrb5HFIo7EtYBH0N4aPhGfNEYO/vj/J
kao9t0Za5Im/FQIqvgVNDiuHOzmz+3xUFr1FB2Nsrbb7pfCmKyL+LGi4MhI/bAZ5
JjCDn8lnIerbFuDXYZGqFbN7VABjoLMZGW6FxNE18+5BrhYKESiRKn4jsZ/YOA09
bpy9x6wL48oCDv5QfFWtwWtFV6Aw24TNQvbDBziPiV0Br+aqjSAcovXUt8zqBfvK
jhLKWm39OSMQwwakjkDSA3N/3PpqxlgQRyEPiLQE8AyX+JA6ngAkGmUc51+VUsu2
79sX7DdlSfz5QrqPeNcAYuPvqb6cQ/X4Go4ekEa0WM++qrZx+27fMWpb1wOZWlHP
+mv8+BNy1/IM131MTBBjEtSOW+7H6FtzrkDCfv02X5MMHdy2ND4qf7IYIxW2tgdm
2+NemFiv8oCETN8DgECoATxAhIAkWJDq+gfOR0f5yZx2p3h9RiVa7iNCB5/g8ECP
ELavcgwK5Tq1BfdsvS4/b7dBa1DOMLbP8j4FiDs1gLC2AH/9Svsr865+jXqcs8EF
uV4rrFRzlrkozFjkyVLLjQpp+NnciP20wLnujkPAygv2FkS5FtCQouj7M6ie5ezP
BlMb8gaWoFlCQuN4KcM9WF0yMpsvUfM1fpgelWEAwWRG/8DH16qKdtStDzctujC3
iW0jpGmKHg08NKqLsxP+k9DEfkvEFnyA0yRKegJbQCx7m2lGdgXhKhOByBKe3rCJ
AMXuofhE76cfYtA0PW24l4x2k6FIeOVB1d2rC2gD1e6l03ScPRxWBD7enp3URJcm
9PSeXlC0OL2pew0Kmc+fhZtjxiguUVaHlt590vMvNAQWOJYTLFkmfHmXEOdnuEeH
Vs3iUVy03Y3b2v+UNQXz353rtBFxVY+H8nUDwEb7ZI8d4SwCJeVc8O8vYQ9h4cAc
hbdipWm3dd1nQGl4MWrFlfNxLA1xgBMOAhU4zHMD1vuRuO+gVCNKrUj2bR1TnFNq
p4YsXdLOoKaiNHASGvair6y02FeJQvY3nMYD9LjbUhNDMMSODgQckb1zJwf7+bRI
hpmN7XjFOovYOfMPynvWaeAa/rlhTesv7alrFwoBlAWob/FQcRrIGMg3t/iptEFA
EUOk9bsiE0R6l4HvhxmQC0ty0hHkBNcEixFaHyj0tlb+juWv6rWqgL4BhNNOsSdQ
DYGiE579NXFv6oWNGIiPO4eJ6b1N+JziBYPuVMFcvcjQSLLkNeetYuwp3dC5mmny
LeiwjfI5T12nPXCLhABWJ7PZTGjskfL/f9EbOUfF5HpRdcFaZuAZsniyfy/yeMHp
18QeKyp+x1DUNHZdmtanWIaT6F9CuI096a2kI60d/UqzAew66J41Y+5PQ0y0MlEU
28YJfpbWV1SLl/D26k1EcMtgQM/wEGvCgEsESnJQf8aBuovWx1BOwPzKE2ki8kCs
+x+1yW3vXrFlValku7OuLMr53LREKw8UnS17HbpBxT99A2DdSS5f5UAgtf1m9uxq
B/jbxG41kJ2DtsGcbkrE8jcJa8wHHRSt8FGbW42BmGLGQVUdgSrJSQqXZwhbBUVV
1ZSJ8c5xEjhxQP9aM83l2zfj3uHukUOe7P225+OfzFi5/8d9yXU8vt+DuTSeH9eW
8eMtvQAHbWoKk3fRvnrJ4qk9jnSuvcaRBrobuz+Hu3895ku6vN7Kdhfhho7U2adJ
BaF9VSCjt5Csj08kJDaIvNFchSxQ+nL5wv9rMzySWmrQoWnE/DlCP+A0uHM4znAW
eO0knE/eWK3vdE/oIaGX8/BhDIW68koEMaz6cq03DeD/AjGzbLFQhzH4CJ9pthjY
F+74ykGu1uLg6zoqAdnlAOxZ4AsbTdFAZBn1raw9YxQ8D5D1unlUbEUrqcf8ocpi
kaV47hsfiScvPoMlPW0ZoNgNbZU5J2w8dHtDTYvElQiMe7R5I3+8BFsOnokUcf5e
KIIbaQfFwNiEquNwBWNPp9RnRWS5NCJHCrIbe4BCTQJsFQBVsSqTzO93QaiGy/Vz
9bS0WTOa7boVuY4Rh7vXMLd1QFlGBYG2pV5egz68VQ2RKxMbtFLuECJwHAXg21hm
dqba5aWl+ISL5wMFtXR6ud2dL6sE9aQFj5LiwZcg7xVieeaTOdp9JXpbNthLtrZb
/TU4pgbUM7f049W+kswQkZRXv51oKByqeiHB0KRsVa/sUXA8g8P47oYwN8ut0/vc
97l90+XrEImG61gTWjnNm11vD/POoGeEVDx+JdiAbj5E1Y33lH327vKPam29jCoc
UKvaZ0XzIxU9f4XYKWzsLM8AbmmyMSyeAGgHDO+sSmorWvBDKk+CfVK76fsI+fZY
OKY9LkgQVKR3xJNKKTjub7CYfwx3B/K052QKz+dNy5RSInw984fzqo+x/aQmIzeu
BBEMPamSeC8mGhOIZcd8GpfCFW4g5OWzW6ELj49ZUOr5tyyi7Emnt6E+ObWFe5Dm
kB8BHXQNgObr76zLAhz/HwEJkOqagimdXcaxR3HWv2YGlPfBlgKaqpjNrN87uz5c
vm58fqOHLt7eFgFYvH/bmK+A9eFccD6778k5Of4/ZodjXw8wKlyCnn7eRD9pPGB6
NCFS9QnWr4I6/917lnh4/hhC9Soi0n5i062IUPkvjDWgZc+JDVBVXhmtGd/P3r3G
Y+kNacMd/sY8vikglS5ZXNVxK71Lwwnp0gBuimQbSwoVokcI1nD/J4BGh9jIMstX
4i1x/EvsHXi0OfrDcZQmcd7bmC9Dyf+MAdaZMH1e7smRnsGrzr5OmXbIeCLr81/x
A/kxwQ3LMwFN5L6KcCaeZb0AN6eq2rY4Ni3gzgZlX+/1D1kpzuB5rSUZ0uXVM3eE
6rbBcrr6tIlNZMoGbOnKxi9R7alqKag+EigC03Gd9+OaCSrLuGIxdwpKK5Ujp/qy
TtXFsNuNq2lxgyxIpuFJB+b7UE7GbiVV/cffEuIIjgyE1JZQeChhFCkONMvYWApb
taHUox3557haoyLGbzNHxlessPgGyCwz23HzVmCNYr+vyAdeSm+1cgoIYdKkrHA4
CMl/Tv+2uaBXza624mBFMjhSvwrS5a2f2gNkepPNxEo8zp1qEO9pAKRGx8XKtHvw
eEcXbXgc2l8nY+w3ydUU9/Rfv6hI8ABaYFF0O3/O5NtPpZcc1wEMZkNJkStJonE1
hrc/c5GUeaTJPlC+Si5iBu3CV5VxcCP36LmoiWX1P8wo0ucEjpT1QUFSLZmPBsNl
5n+xVOjgg1lQgyoAu3BOcMPrGG8wHIn9RNC5Jxz+AwX3Yn78NnyER0SPCKYdAj7q
xYyehhdJfXOmuhhXbeP5LeHgErh6Z4NrXMptJUeAdy6Ba+sbWVe5c2TL6LK+qWIB
NF5bXY6Fc1Mf4ewcmCtGWQLuASE1JZQD1UVUHx2uKTCOMgo+wu1qyKOqfvENVbdN
lBPYilft7R/yO3ifWQGNroE/k2O8oc8kz7EXvJ0cw3fILulCkhxsYFMFvmhFzM1t
SydDc6JQN29nu396Z4wVjXcgn52Y0zNbEpUXPkXXx3YhGpqnFw3zuuZC8je3Pvbt
hBKFRMAMJOxvfH4AhgfsuG/LUEmLkompW43ViYvAqGvDBVJjU50zoKY35t4XyOF3
3VWLw+XmEwwUw3/8IXxymfgy+zlfzSGM6tVYo08TUDisDhqGX8j/CYdLOTDryo4K
+JiewEvVhr3mSuwwcUWJYMBn2GjUSABGG7Wmt8NwFNV/tgdLe8N8EiwVw6IyGXkC
MjAjFdwe3bfuGu56Th/LsFZVssbaNRJBQhFU4r86icP54AlmW8DfrUQwB/pVCHC5
OSGOeHO0ldGCGPcit20cqer5N2JBqEXu9qrex6vGa7M+NFi7scCvl7p4KbPTxDRK
jdhCxbrp0aLv07t+xd8OF0eJlRB6qyKIX1glQXYGOdDbKtJU9HcNbQu69yKqTYrw
HQoH2BEM/A7abuiR7pB+1kp16vQcZ9Rj1Luvw15hajbd84dg73fDC879kyC1j/q9
GPNTo5EmPPjQTUE+7kFPbzUQ4zguqU7t6h0reVLqJex1/BctUYdbNXDbdLW8plR7
FUsr/q51HeSFl1RBeQ4HXBB5TSalTZRHgph9xEWsAx5E9al4j78VP1ZpOv3Pgvxc
CSDhSIEDtcD5zTM8JsJKzNdHMusxZbftK1RJNcSZy7HfQeHJj2MUSm4yjFdrI+8+
0ie4BDxpgsmDwQ3V2G/7B+4rpi6UMTnfsnQHi9U5hGe87NPolOulTy2/JCV3dVow
vbYyDs11o7PQ1/tH8PTdvX6jCuG8YzWq4qSbOxxGSA3DyLI6KW7Y1kbLH6wdn63m
mgzMiTgqDbjtJ2aAZl/mJJD2J43u+/ZDiTwe38960yNcSuWUd+LXHTibpkrKQeRY
yEl8emUi+O6XzR+oca91S4ThOgcE4VFswbUZtrrXnQ6mDmH3uEtUK5+hqcB3H13n
3y3w3FH4Dk+tO0Qcz+ZtPLZtbif/c/nqGOsw3sQoC2koCZPOPYZ04o24dmxVGwsA
LUFXulO0JwmQsj3GfzljGxY0oOJVmePyR5tFTR09oCgg/PQuLvK0XcYy3vr6wW2N
zZQyB/dnSAF+mwFO+VdpmNvEdNBwMMXkL1BbY/uUl0QISLoJiIlq4RXsIu9yusrj
MB5Gmzep4nNafqPC0epqcUAk6BLdOllby+S5ucxvQa4rZVq2ACobjrr2J4Gt1h/F
kSiuivX2kciNVwd76oVUMoOa0Hll4FTv7TjLktbaMM7sC/Ga34xpaZsHFFsaI8hv
DiUrt/fw2lS4dwulouawhnPmDHhoZp0IouoOTCEs2J2l7If92wB+JQZONW56leA2
AGW3/vlHUyKbZDxlR6EFht1qRGO5JW8p2Cj5wkI/082HR6xAwdtwCNb1GUAya3Se
ml4ySUWavwCJ00tDAG68ejMF80WiwmupaTuu6STPVVDlT3KOixoHailpvMtdB5qE
SxfyHTa89F4dho2HqTsQ9+GpzkCLItc+Ps2RjrG17eFEZ1anjOtRI+PDv4yC83UH
KT+OAh7dOocG4BdbmLhaI/aG9292QADozwVE0DkTxquPUCnpgs7/inPDNhUvnYx6
8VWywkII6S6HvpePBJtmaYhO8epJzJ8xzUx4kwnbZCc76DbcwDrHL0ih1pF5iI4P
wiMepCg8aJtHLhmYo21YsSDeco5mR+yH+8hZHzAAsrezrjdNL5Z9NZFS4vret4tU
5IaimGjS7PETnfYyIoUKV5qcQQIyhZrPZqGTfxWCFtpEtmihPzMsCz4Kn9PmvYus
+F5/WwLg0/gCIJ4p2l1H9bC927DTv4TKpAb3EUwhAB52hnYZbRwvrIzLMwLcoo45
t3iMoGKkOcx4KaWBF7xSvlV98x2tPtwr9SDNbjynk9czx8T4opa70jJ0w45Pb0pq
HcdcOupDFl58LOL0IOzDE39xOXoLSqwgWvEIulb0QDiR4TnW4nAu970tN3j1nkKJ
0FJ5R0P/lESvTGv4UjnS4uLBep84vtPbowQdYD0CgzUttD0IyN+Z1LIJOSjomxrM
Gx65qm4inevuRlPeR4iHsQQMmaIgUi4lHpXdZyNYTUDtkW/yJW16Q6p7LDy7Oh1e
jeDO2sKCZPmjoOSOSuD8B6ZTwVhXomioZp20DcRMMO7dGuFJM3Q51OSKoH48hipp
LHnjDjTqyBK1SKw5nSxWC628Ylke6OfCVy6eiyOvIB60sXyD5tfTdfbco2BsIXTx
y/9pWbv3ocOi5K/iMBZR0AMKPZt2sVNWfo3MBXSwKvJnBC4+aJoanC/+jMmnL/kM
OMfsSSt+z67hP30D1gyL4ADruchjloD8ii6A5lhE1xneStIXkNOJ6v/M1g0p9txf
lTugQtpf90jUb9oxkkwMxXz35GpFMfKCPUYGXJ9Nv6zf6Qjxlus2HEwJOXA59HGd
DLNznmuq6N0Morgc9PggBccHKloB/ghp2rERKcvC8ovzR4OJvV9m5UXTATmCuAdl
IhrMBehTQBzYOJW6uIA4B/c6vjoqsc28+vGYubt6qQ6BDZIHgPtBzzirLY3UTbGY
6zhi9OinWVLXNMjvYZAZLlsR9CFLv1VOLzkDjMVcCMu2yg/hWiHZXPmis2k2ClWG
9fPjZlIfJLKvS243WAHyRJv5el+81PcFv/6SV/VYbU8/ZeRkRpuwc10VrVFhJKPG
Bc6vrMBb2h6c1bTFl4Bt/OTq40hKKj1Y7dIyvPg/rhqWYU1qy7NLdvJ/WmnCCGPr
19sIXXzMTDDCf4WS+HPQF1ZkVY+zqN1LzvkKv7iElWEvn8FXFo0zByv3e2dVCEO2
2O0IS7P0PcH3BZUExtYQJozYrMqDBZnXUW3m3hGnPZ9bDVIfJWpMQVTWEwGCbCf1
d6dK9eq/5sPnze4f4rLbjRJH4uNki1F8BjRcbF2Bv+2CXPXflk6n2Rr7Z/+3EKcL
1gtaNkJunGlGyTj+N/lLIOaiYcChkPLhdycqhnCGmsu/QHhiO/VKgsCdrHp95dii
6KgOASlr7qa4sRAXOyEYj9In5wmGzGzwrQRQcz9r4HpFL6qn4xr+0kPCI9lu1p8l
YdZw7p9GsEQ5aaSHEZYeKRHH2mrXKDxwopDZjDFWaM6uJtXMSvBAL5pOtAsPhwkx
F/IuqebDpB3AYxBMzUj1tHdNypRASUAcQG+Rq4P6FVhUrJ3T4MXYzzGD9H/Ul+9u
kzV4llGGhq8rkOkz1U+K9CxLZccY6sSunzf2BC5jJODu5klBF6xKs3u3z8bL6k7w
dNy1FC3lUnLaox6B//IEcAixTJAOg7ug6I/L5RKmsVp13aJmvNXoFRbjiDPxOcfO
tdrwBDwcyehKeRaSsdvkbt9EjqlBskAqR7uP8s5e4GsS+uT3BKgLJUP/JIZGGmTu
t1jkrgMLf+jXUnNvbqGQvA8HLkCRRbXRbm2WTEG/IuGdNfSE4X4d2dyC1NdVDBFE
5fgtkQmkEHoW7LqOB7h3g8e/Bxt9MfgERKuucH04xs5gXbzggKXgBOLEy+yRHaom
uLrzQF10lCyy6jwtBJbVF7fJTESsFsW9HpNQ+0dUrmIFF72jANSoRqsJg94KARXk
+3Oq+8iweBfL8Tr16Hg8Q1Zo7zsn5pN/1df7zyrbcnvrEqPkTN5RFqH/znh0srIt
x875w7RoeWxt3SXyIVLVx9hsFyWhKkS7R5nLl1X/I2SmpI6PvBeqAylm57b2+nzq
3JkzpUretj8xbX+1N23nAAXCZiMzBlPUMrDBciQUXEBG+3y6JmOicpEPl5EanlTg
/Dc1kKnwFiu7SQahLPIWW55WIPII/91k1slXI48OUoNfOLeGgAChaK9mXk71MIBC
3sNjqiZ8YY0LdnwPJSV52k7q65TY6+E5UhG8wuPtgsOa236Ypi8oeAbLNj7BsUYK
Vw/UBDCScnYlNv9oxzL7PtR3z+w94E27DLh0rSwfqz+OavMw1XEbLaFGcWa552Iu
MJPYh07u+ohU9FsphBlXh7ZbEGZ15DZT0h9qnC3wFlY8mvEMR15I28hEuDqDY+7n
qtNCg+w/6ZzNXyS8p0ua6/VMJg0BwSrYqsAzpFhdSCFeMbe4sMiJ0l8T2yuNn4iv
m1yQaas7Hc44j3dZx5Mi5LhVbAAylv0dH65PXa0Bd7gY767sN7VjLtTld17lmiEa
WbzPt/EhcIRBPYTnyw3RLwM+7GfhWAeD4D65nszUg8/BoEOX4o5aC6haXkLsTTql
KVnxSz4FnEXvx6BslU0vLUVPByxxtCzCReysfRCufKxQYZjZxcapVqiOgGjOlmM7
6dizAeYd6V7G+VGLdEX2VxmMPB2P+A/8mzUqc96gpAACxm/In0q4jQxhXxmSGoW7
6HCbCCIKzBRFByohZxNsa3hkO4FIpFXORLjMMvVNz/ac5gx6R7Otvn8aBLAav1Y2
8hdymP5B9fJl6kT4WlrrQBW0xQimkWWb3UEoJDAvrYvuu3aGwwGs1LC0uZlVSSRP
lg9Zn8UAM6ZuvxNlqzJSJPC3famhVhRJsRK1x25bmZIMTEp1B2hJP9RQbsokfA6E
WvCmG2yQgD4G9igWaJoed4uCmnIKj3scCc1o+9N24xHZ9wWawVkRydzdlc2tZvbO
Iq1GGfEyqZhM/ZrPqIZ6e9/mX5zF1lDskgwi0e+VCA1QqPZmSPYBXtBa22bCoyqd
FZhBfp1SrMzXSYQxC8MFKAy7nNd8s2GnWKyHvFsVkAMMu3xn+yJ0xgItlH/0i1V7
0lM47i5Nul0Xr0ixiGwPBOIiXEcOyPMR7Isy76mY+rb2x65yEi1S+M+vkZg4HkTw
RdsXIXPyWLJhOOjrRcGgLMjylgFn3rX3xIQxlCYZzedHjufD0uBWsgtgz3tnnEpP
7dRhK6uiuUj8Aw0tUUEsbXhP6WRkXEWtGue4Bf/Ft+CPH9QqlXqpApmg4Pswzm7t
0nWbQ011CJRCMunUlsntMQxJLT8zg/fh6MMvEce7ZTcOgfWFr+2LwNX2SWvu28kw
nBVX7zFckyMKVVw7DijbHDe04E9fB1R3wkkDENr3ezDWrB4OrLoF1/m3vskCBMbD
pY19rgTrWlYG4LIGcaJg7GHOgUPHLS5Nbnq1gIMDqjy55hu8ZoqKwjGMaNEZOf2k
EjiO0kRR1dXz++CIgbmt8gbVtzr5ruBHjebPhkJ0UWtvKKMkPqbALMm0aNdRYLd7
NUBmkhE1CEmX66EsmZ/Bd5Q2mvhAVU7+NHdqdhHkobbt8GHpZPyQdJJtNN3Ub7VL
JlyyiXOeGJOI2P6S0jXK+dZuOFGW4dIwgYr4wp5K3pVgdDe52Mk+QNzTmqOEJlAJ
qvuDL/Zf9ut4qTEAA+vAGNQdk7h74zjdC21Fa30BavBQ1Wr+2krubgMy9ua5TQkq
HCR5SbVKSFgX6J0A2lhVCGR6szacj/6gtX5lHI7xKt8XzLl3dfRjkkd6Z/1BYxA4
eH8gkXT9jC7QayNCzUL+DYKwIKVtGtAgB30+OE7uJWBkOuVS4Vl3aerhW7JENTa8
4rhsnhxb/AnMFbHQAaIN90IpW9vqT5HEDSJii91+DRpfrKu1SX3zLdIckDeiKoEp
dJ5LWSXmPqhhQoXLVqzwtOVUtKWwe2hnwdN17VQBHopMQv2e6bBw8bHm5NeuHprn
aB7OYIwJp85a+ckM1ZceDziPg2AqfLAjsrxz8Kc6yg+Stp+YKTXH8sxJ/ZYBSZtu
eVDZn4N8gWWIbNAsuQRkbH0/uYKjxn4yxagQofSCyuJYdQUP5QXoGrpgqf/DOZm8
KOrvrg/Ent1WXg/ixGuZbiF24K7XhCL6LCKuH5fb09n47UJtbw5mKh+rO+CsuQeG
JnNUt6YNAGovY2V3BgPPJEXhz6FS2wUx0Y2j8wSg2caA6n99HITSt4HDlEmD36sz
Jd2gf+SRl0jmjmKQhbzrUbzefZ9goU9ZYJfXABH7dAk7F40znCIF2OhPK3bu8apJ
hmUB8k7qLkouMFgjMXspnNEcX8bIl/JoIpPxgii/JPWou11/NNJfNmsxdgWgPnfx
bQ5noD0+agKCFAkQfuZ4JtJZ0i/u8m7XPzoMzN1O/ZvFz+ISpSJbdi/jlRRjKeNP
FZkXbXRfn8+RgFYxgxPEKCY/K413F4wk4oR3SpZD/MryZEXScZrfbHM7dnHGULSe
LxGXnWarRn3dqxoy3KkHOHB827O4T42dkGzAA+HvSr4x4HrtluLFu9nLrvOJTdn3
MWORJ9lstkGKglX19ivMo5gJkOZnmq7Rk0lNJXrkLPyxn3uSlJ6y0vav4a1qIHBr
8LuLqIwa0icyvXTQXCr5cwpmnxUttL+o/zMmawD7mlyGG2/SRJUadvezw2UIxMnz
JrFGL5RkBFjsgGa3aIqs3zQZoUZxljG3eLgzhvEvL88KwxbP4AxYe3Y2WnS+N9Hw
sXwtTeQb8hKZmdEz8AmA3kEozmblNX1NIV6/MAQaIpUy090iS3b5ozutqAlSiGx/
J6LvnV0cDpzcNd+WSMmZFEtEZJXc2tAbVutJaLa9mma3sj2GsWx9b/vR3P5Rp/8B
7BH29zAFhRWkZ37j3WuqOldZF3t/ENntfvtmh22T5lJxy7wIiabf+TGf9uqz6qrv
cid8OcRx2n1ywyU5pwGRrsV2i1Rhf+Duom+R7PJEv7vuM0TrFPHiMO0oao8e6dX5
bZETBP8RsxFrkjcjGlyoXWWIX1lH4A+G0EckV1jmbFiuUg4XlwjxmoQSfuVs8/b4
OGneGiz4GOGlGYpDtNwfNNbzWiJ1oHxAkrgDkiII7mIFr8ITW5AIkkuokRnqGk86
cryjdGoQhzVJDPyvJP4oHlmEKbJibLsGOMo3A9ZvM9d4KrSI2m5yNO+jwva619wT
3w8jd7A1tpyCNnDbAr3JA6G4yKsMGgaTvaDDWcRxJkdcfGJnVj219See7lhD+/K9
xF5g9bjPjLUBpP36f9/AnTEUvsIXNa+2imdrBfQc46WKtMusYYXUcyo5pqPncsXy
9NPmP6qtnh3vSL4waQ5MirrrcHqz3yf1A5AZEG3+Z0WZqf4TcihFOe7U8jZiVLdf
H4S7TRFsu8AtxCVDFspZeobgh+m4ofM8Z0aTRugh5wbhwczwXjuAKqtzv0n5nJr+
FwJOoMawUjjnc2RRt2e1py/LtyV9Wm4a2zLnPpamAr4y7PIIcvUBeUzrPcKKH/3q
KrjPRXUbi/s3IK8agxAqVqDmTHTblFv9/D4caN2ubhUGkb3/SaWNC+eD9O2I40U2
EVCqQfdtTSDWc9NIRUQAAzPyHLJr9gT7MD/RbGlUohXGEWhBYnZ2VuprWnRZIIKe
1cAALKK91hxNFzsms7Rg8O/c9pHdV5ZwmWM9zRAgK5hgGkEVOV6YI4IbVwyBq+HY
AcgzEcJOBatkOb5hkXgV2ldslpRj+dwkJPR0+zyekPgjvxb/qIQW+JbIxXDnrPex
2POtc7En6ci1UiBy0MN39fsHJCJlwMx2S4LPlkdn6tpu5sC9JMYBmWyhTDH0PcYp
EMV7Om87rDOEX+mWJTnbr6lWGqafrqpOVMheHEFIWA8OOCnNzdQaujwrkayhVYE6
pbigKutArIKFa3NRqF4udoimM6PeVdZ1PU4Qd5/LYQaZfwwOtewJVUvx9yZT7hwQ
fyJnLlI58To/qjHO26LCE5GBO5G4Ue+yk2egt870UpZUzTgrAGVRiJyOvxWr+4ZN
/kEaeIi0I61Z9PrPu//Wjs2NQ59J04cmXP5CXk4hM3RA/QmHyfYs7HKYUcegJPXm
TGyrTAsP3pfx2++yzyUO/Tvn7NBYfCN1eOPSKOWFFL1RtefOn4ehyPz1WIL4pp07
yUjo5BRv6lJwlXLo1UYkl0D8yq0KJ7a15LsKMxrZJ0V7z8wcD8OpGqf6M9sSyFCV
0faEqsyNzlKXPUmbzkKJ8pNyoDTWdcaVmbrZrLCMhGO4y+fw9J9v8uaEmWQYtxrt
ErOmlmNBLpYnu2c6obF5RBOIQjbE+CGQD+maZ4Ro29gTpgh7w2YUNxj7ew6IT2aY
6tWK5euG0alTLHAXkY8wVgNOXevxtjCh9loAlRoFtcgzveKve4lLiMUNFdq1fei5
RjHIVpoY13GR1F6iOOF3YvKu8LEOcKpYmiJRUi1kSN4EfZ/ETkqzTQmDCcnbBFG/
s9M1FXInRnB85bYkwwmUEziiPmKm9nIRDHIgrsxQPJvuhxt6J9ahGbPLENl6ojX6
J/3zdKoc9GjPSjh4WdEAzOULWaMKQiD2JCj7KnNKqEpsG3CSp7X8oOh7+KYen81W
ceOy2+djZwufYLgkgLU0YCnjMIKwqIwFUsqCIW+KcaPJydZVnkrrPgVmURNBSa79
/dj6Z2WF5Lp9TYrtTivhngbk851BvNWh1rSTh58teVSX6igTyVDJ3eJ7kG7GQOqp
WXRDGmIpZonk74Cb74NUzvw9ILw3wKTVjhLCDQ10NsPcEkvgpUITAEOMxi8AZtuQ
HkiCI5imKHlo27dKpYzCvMQEg4eKO2mwEM7yOGjhx6m6a75sRPz7KFuroZH7+E8x
09CRcuNv/DKvtrThp8VYR2jkw4q15KoV3uMtNrQNjr/p15IaQxFN1jNbFeFT4OID
Mgf7loMVfmkkGch5ZykHsx45C/odiQP5x1y10nxEXvYGkRlmCuVLzlMgBHu1NdM1
7IEI1FZLwk0AR2AZslyGF2es5J/MYKsz8kRSTJ7dnXL6UHhhDVP5AhLkR829nFha
bnTL/ezSykfb08B/RqwB/mLD6MrRil1MgmFB9EBYANXtP3misOO3GJ6XhBbQFdj5
a8gXcwtx+0p66Sg2hh5D0qYfsXfH0MixEjiUpN1cEQxkzECu+RZyBd6iaeVRFv/o
uGZD08Xjs1m4SRUwUm9izCM3QUGAccJNdr+pvE6Y+Plkw1KdIK8O76ULT48hq2kj
cSkrvve90sureDEBJwU71wBIppEvh091vUxEvd7aUcwolrYfTxeh1CQVbjfP47u9
PHr8HdcoCQjqtmtk3T5SxpcKAnZ+W3t1iaKkztQHTqmRA02qfGcdkrgBXJty5FV0
BSMO0VDbI+6IG3oocghcGKgpJEl+Q6G0YjkevUE7Pe+jJYDOkZ+Lr5FmG+m9rkHX
pByGznyleuDtfROIYN7z/XOXY0uocMjw+cW5KhouJdMaZ/s9hQ9FUevB4mxvqMBy
C5kxoduH7bsTaaMrjbLDZfXq/OSndJkZN1yjRKUGXybRy2BEUPwcvGsQkmRH2BLO
QvGQWF8OVa54rnF6pBkX/e6nJXw6FwOE7VFtesiED1SXwiXnff7iZ6cS1yHykJbU
gkPin8iV9jgkcSlnK3nmn9kcAe8UA/Z5WVKKmlCk+vdK3T2fd7FUH90SVnvVYNZH
sfA3cF7Q4baSGQ1FrkpEu53AjLHs38blS/uNeI1G+Wz7Vm7Hvdlpo6+GfAwMlr9m
eiaBXJu1cJJlnf+gnJgmXvdWLAZW3Mks8eLh2A/qV27vNyNhmAP1nMz0SRXxjhZG
CFDKmyiCw71OkIQ1ET9Lx2Lk20Pobn95PWzj+NkGbZwNYz8t8mS19vDqHiBaUSC/
COcAMBYHlsmZn5wzqYRdwVKpHApF6W4Wen+ENbeuNae9ZwiwAn7z2otBPPqR6vXR
8jMsXThQO04vKyoNFY2FYg5OaK3f1OvDcpJ7T5D5HdIIRV7O7j8b0OeR1uU9QKtP
6R8oxHql5TPsL1bKWv0FuEfnBoSabJSqT7Z/0+h4E86o1mCrT2ve5JHxfGY0V3LC
YE3jY/jNIZ1FVCRc/yOZKAGg28cCit/gXXPFDeTTdb7KqJjQNXL4n0hd7iGsHI/+
JyxyC81kfhvGS/xLlClvSFStD9YQfUf/4qYT0HTSSzQGgPkgk/LAzsfI8+MswBF9
fnl1dXT2/JR31hzIfxLvEQMAS3EBTRScibHIhmQBxcTQQ7OCwiED6zNUJYViup1f
QhAv+VLQ5i+6MsaMclOS8AL+MadWrRss/bRgRsfbdRCPIFzDOv8CJh/Ntxdwdw3F
t7HwXcdKfgeZdZ4Brh2AquvAoB49cEmq8ajuYNGCPVv+Cvx23hVdvP8NIRLd+eJM
0dl2+oC+sgXSPm0QEnPCoKFSmAm1OGiWBcpPqwtGekX1RAfjidNTkM0elIRRZ5gf
Vgj9xPqtPu1mekDfXJKp0k9RQ6nB3JdjfpbjUPL1GUNFthbY1NFQryEH0mlOFkbs
IomkJWXnzYPIis/7GYetp8aY8Z4HrPOsPqx8FInSYoq27desqOoWeZulASocz8FQ
ktwvKBz9vagQVzvK7hnUZiO1QPfvXVq9iMx/+h1yEcdLiSiRrKlisQMMphAPhiyM
gsqInKlBHLpYVi7Ng5dfXENd+np0rUEfDmj07RMRa/JsOttsF3Km3uqFUGR+3TZj
LOzRUoQ6sFdCKyNUT6xMiEI1z9DBTHGKMM1sh1AQBamD357XFcaOpquB8HINOF2e
R0u5aA9aW1FWYaCZHbiwLKn+TsbEOlTtywoKTuaFRRNmazxzeCMf4RjWqHtFywEl
EV1m66XcDoqx+Dq92mG2645dcBiHuvgH/NAiRLlyf+Dns41PsE/Ub/4UR5dDdyoh
cUbjsexVBUQcxGnwtYCTDS4lJDeFS3I6tYqbouuMjsf7Uk1ukgkOIg9vjf/ZAqtQ
b7UmVi5kN8ILJYJB7lzUUuajLYxdW78+R4iCq4pTUQ3QmrGddtVrBsi+28hBty1L
xD8i7g3BqmKR9Rm6mltPiKioFO+qXtmx2Lmo5h87EuVa7wsCXfypt/UcIJOKe3ZK
pg+u+cYLLD6Cl9dsiE6lD6tOWDPl+DMIFbrXgBftv9kgcyM6CNA9huC2hUsPss7d
yrnEHiGV9vxrLUAmE66y7rqWsbhY+nXFGPCY/iRxK4u9aQ53QB5jnYgJIH9eriHm
mLCbCyRAI8JStiUuIwDwUmkVysiIEBdyVpjGvhgwgFUPJEgIHQ2pB8nv+ZWrc9w8
QbYq3NbCVhZmqNuTU0+GqCTvMOMMTcGAncuHWDkwsAzsVsLS+GiHfZ0FOobsCN4L
bYHIz7BxQ0d2YkduX28eboyXY+i28/hQz0XlKQBHe5jfzLEbSyp7KtdEk/iAL1qV
pQuSXxDwcD/0N+xgbn00rmYrVsbNQHTEguM7nn3Z7OijdriG2f20sohKsiZgrobl
cmk3lNF3/AMRQgTMlvKBE5BEEGiycxTVaUaA3J5jzrxmg8tuCiWiZlw1HlsvZ+1e
JUDHY8S8uTey7kKNRiGpBzPOYSuwQ5QxVulZv/5g/XIBcDSdx0DM4EHdQF24p88R
hysNOf7VxN/v2YhHMg48jCA5nUoeDZxTYSlZtmi7lz10apoJnGz30772mLyWyfPG
+L7x/hpKwE3XJc2TczfZLZvlfQeAI7NtLV5PIbJFiYWaowHnXoZe5O/Mg7RwmC/u
5Y1/gViI/0Yl2xhXh42vdKO2SBo/KrdjfN2SGP/5L8VG992TCUR28TSLW9NrocsD
JxqBlvr9lBpJ4eHApy6ejyo5jq9t+UL5AOj27zGdCR91UUuBDQdT40SAOUf+r8NF
/A7dgxWHHjNQBgsNgCA5GCJcdkUFJhca818mBNXDlLI2UCRlES93pCD1h/H/nsnK
bJ/Qf2H69N9m+1ocIvJirL42DQ9xyLsEE6eR4v8xBN28muehwDRc+sd8C4ESvCuM
91QScFhvRbL7EEe3J1hzxukQ0xd/DXdy2Y7bQnPPzxpKej9laG5zGlK1dxUbw2bJ
nTbo5KKWmn346VCBnPwcLsEhcKj0hioAArjifrKD3NLNxd5XBxlTnfRunBJzjyHd
Cp4ygzkyoi+f/72lWHkDTFHfR4csgdnCHabKHg47wDW31Y+QGkevuY+QWFMehQoI
+UG+LrtPI1qm9YJWtgAaY12dNP0h1xjdVxxpv5jEPjmQz5CcIALicZZXk8LbkT5w
afAqxZlJ52ajbM5EirYAIp3+R1R3RJfp7+x6Sh5XUezpuBYpUa5kwdErz3QXxLPu
lTmGuGkkYEltMacjLpyhR0W/Ba2vFQO42mCgnJj8zys7TZJ65iCFcpGbcLXQ2w4C
P4fCYNdkBShWIz6WFuzR9RWStKLLPgW1BJz3LSTbNj7v/xl0nSJtxFaWMoBLfNOq
wvQOVOGxJXE9AILVS2Nj9YWagtR7J1EMZwTCBAUmUB9cmGxwsPz7CZm0bJJUWQ1e
LXy/dpmXMx49JaAciQ0ZFoH8qGBh9TM5JOiwME4A/noNuMRvlYI3RFyLc3RXcygH
OwAuTIj3VWOuYCn1wJntP7tCn/N8dNSJWrollHZ+jPzJifXkRC27Ynl8iDV4i9/9
ZSo++rfRgmE87+aw9ZNjyinXFPJko1VTTEuRP6vVEGwfe4shzShKbY9QgS9u6Qfw
iNBjixKXq3UD7hA50XCSIMDcmdjHPGL+iZF1vlTxTrMyHrbl/NHZT1um8Iu2HQSB
1yollLtG0cdvPiQ5RrdThW0XhcENWGZkoMiDk7u3ZycwBaJc6zSJ3qmwivD8lb4D
Kg7yAlCLMVgodq3xgGo9SkPfUd4Weiz8LGi1vLT8p2Rz5ZOYV8P7Gv5kkwj7p3N5
qEfE2AfMMhvy0bS4lQaqeVIa/O1TxnkcolqGa4fyhrhhLzhPENo9gR4G+tThh++r
BDm8+Kv5tdlDCP+DsfxlgV0s2Q4ontQbiBpA1hq5jLkjGajLKaKUUXhQgR+rF5f0
6uLwy4TkxRjFMR5r7e9wXpi3Jo3KtPnCUMZQh9BEViICALccnB4Txmc2qpm+ATlq
OZ4XOv6u7BhrTCRcCd+TNOJBa6ssb76J6Dy+Mj6MrkoYzKom6CURrSa2PufoMpRR
68x4ulPGQYwZ7tmabd8NqChF0it93bMYHzNrlEde0qm0jTxYAVupq0KjhJ4whaZr
MAhD/umzbRwBrL8jH268dZfyv1uGGXOfsZQoOpIfEPtn9xtSwrmDLb51IUGMvLlk
mNXBIl3dx7wbPlTpzKP3K+WE6Ozig0DTD2DSHGHcFmNoG4tqMKQPg3TCJWVbPs6k
fem+Kvc7x+aroPwVT4P7yapep0HoPmzbZCT6sp255HA1Ac+vqOuelUCxE68+8q/u
qxRatUMsHjzU4F4579w7b6OwzDb+LVfgq5rarEfdzem8F4r/7SVXH3+Ig4N1paqR
HnkGmTaUq0+XSyn8bODB/r0ErOeALUFWkXBREtrTB1kjHFfsm4JtOC2aAzX2sSHi
neYjSiO3gwzKPm2oO9IrdQvoZ8NogMvGw6hZ3dACr48XkJRwTUMgK0J3KgcPDqBC
tTvDSy1RQEzS7scrMoWF1fYTRFSvyS3ASs1WA2/utgxHe71DGdoQgLhapWi1Qz2d
AhRY8x4tm5jLxCuVzuxP+lmdIz73A3bYsmolYQhj6KdSd7Vxp26eXDnu+o8FaKxK
jDhgqofh6E9kMaDvRctkL/LD6oZprOYw9aVoFUfE+rxUu3aKRVNDUUhumQfQgUAC
0RiWq26fKXKHQSrpU4cnLIlsaApl8H5xUPfcGZFl37i6VVBt6NMXhbQy3cBWEjA9
glyakzL2vYopZhy94YQ3JM4wzkSHq+libTAYN6G8yAJFu/hZzEuqwT2AEYOHF+4O
dxZK897UBTcDhq+dJbCoYc9inSQq3/FVunAqPQOv93xq2eBJf2zGJNm6/e27gmgM
Ettp1UmQOp3kFbBGfmClAG8yYcg4UAdaQcel26vinh+MOfy4sU4dixdrd+kuxtK4
s+KUnWf3erH+yLsBzHpmKWEq1m0w+cG0Tc4Zjz//cfzvdD0h7hIkzLXcmuYowHcV
2xwNOnUgUyHwM06MJ5XABtD6qocs5RlGj95uezgeMi7BjZJzava8Qw9CjtdOaq4Q
9DhNiqJJ9cCRwrAKJu75exieFLKewn34YuowogLAaqgbBPtBlKfiE/RCw+HBbzh6
/Qs6wbJVFVofTQEdajqtyfSmpBRm4JPVJZkNdTb0hHCuNYboMsG+wxx+Ngb0kD/E
rIfNdFqBoIoVtCCCJcA4deLtUPFRfv00fJDFRW2cHYBXZSjC8jvR3YJkpWCapYbP
dGHypF/xqh8lLTa7dSinFm80oUt5jUtpBWXkufWGO6rHgkuMrG5C5sOZojSl6Gag
kTfO1T4WGLH0wwogvOv4NjHd+RsdPrdKYF9pCsoY/fnO/omh5p72H/lk/mQtRKXs
GhbFEtdZCAPKRQRC6kIRGDSAcyuri7fHmA8pZwCaVwX9SpIsm62o6VVoxMogiJmO
f/fRM8TjdlCm4TPKlWZE5jp1tz6md4VEPdlh/NnmH9+7vVmfv0ome5999ticclLB
0gUMk+N29as+iByKDDfbu3zEGS0kv9ruBCRLiZaZZBvwD2FgfTdWivwcVh8p9Zb7
vMjCYFoEiG/Pde96iHd6wkD01gclsKsh4chWCYIdloI5hEEW1RMMNpw8BePn/0e3
tIq/PjxPh+ZwC0zYoNiXuvOQG9fz7pFGD7m6yzi6nHe3DanbuMHhF2jXkTznsOoM
2iL4G58T0F8t3shAKJAdb8+HIeSVNqK8zXm6gwUtfaBBnQNEYAtjPdJxT/n9Ck3+
tGzv/wsJx+Lyxb+urHoqPmfXkgNcegxPSwRowLZkaeS6K46pCSjtK5IoHzcKixdN
ZXHHaWmd8F1Y8jz9xZWe3ZCu435NEcbPBaob93lMA3EKcEUqg1T+8/b+7I9HP9m4
q3nfLKE1nEZtjDVEUhHUypS7z7MnROjnr/drgqZyYio0qEarQrQDDXf7aG+wllrM
VkFZL0QGcIwCR2lpnhJb00RoTJ/t669szhh2cExXkrwyq5yslAy7XPpJ8eOhmi94
8MKOsYBB12tMcHwf9Tf0nOuTP9o/BgmaboAir7x1Vepoi9U/JKPxDu7ljQut7AMg
4WRdV03ebnYDoemcyXP7rZ6kglVsilHpCN8EcLq6o69LR8HKQJKxtGX3ryZRgmWn
B9rPAD/+Lu6YvwO9gJO8dPlkwdXAy3EKcpSTsa2xNXmd92RMtGvY3jO2h/AxB9eX
TyDRblQ89ij/aRm1oZCdc6WSf6AR0O5rCdq5VDogwuz2HBedkkwAXiN3R5PLXZpb
6LDVHio9rRY/1D/qsL6Irc/Ree7i77vGoFc6Etp40TwW3bQMDZ9+3gXpcekfjQID
FmwrtIZ9vz1ZWi/WKQV8ooUgpxUe+xAAWKiXStVI7aC/TbN+/0ltY9InK8TUU22I
arrvs7sh0SGtQAw5VdggvAvPi3uptx1iylCkHSLITOhToj7a7bKFSVrA0T6SQzc2
wNvWIXUJaqCacY8A88B/3eFc0FAVneR2WrhMj52kOeNLiuhElHrGPkUIiPeR+bnD
9dKeNc+aAC+Oyf/1YJYLtci0GemcXkHQ/+u+O74EZIegqrIjFqVACxbcBPWeQSLa
5mojbNF4Pn63YqB7idajq3yTgCTOJJErR8bg/j1n90+zx78ScpUfO3Aqff7MKC0L
5HTIcq+myMjV5GijTtjYEVCJMoiL3JxymlUpbL8UvFRhfd4vkoduuXnUi/LftdMe
9ghTt3qDNkoQxBm4rmmaAFVWLmX0mC52MMz4Z7fu2hDI3XWX5Tr+k2OB2mj9L0lM
FQt623oU9Fz0Gj8ZrZ0lD9obLDOA6HfYyE0cq3Xw3oynnHgidx1PNIbestVp9LE1
qYB4GXoywel1qHm/ObmIH/cHAxtKSE9cISSLk6BXIvHVF9q8Dz9CtyvIYFzEZDT1
VD7i4SwpigJilCxLp9YKgmaFujYNJcvPnAXwBGCXg9k3YV1nVu6KI+sLIEAX7fRa
D1Ri64Sr/K2Xr9HhvBxF9luZqtbA7XmgzTvXoZ9EBCjMcbEsmuNt2V33t9VP188Q
n+Vv7BMbMmVFtA1eq1fQomBaM1lBmX7+cKHaJTMBeT6dDP4I1by8KITA8lG1BbRt
UwwGQRIlktJB1tsoS1AoWqh8NbVsAucGyRdz56SBzTc3BR0V1qLDehTF48DmSTrC
N1TpVC5CHXbwc4JF+Xemxa57UEZ6uwXDEP433ZkG+JX5lx12e9jFqJl7GIwr2wtB
fjBeOYAlzCNVF56t6GT21uhQWoEedJ6Ia55uRbjCqvOJIPFJS5lgVHNg4oA8sW8j
rTKFU1qnZxVCn1aY72aBMrs42E6F9WMd6DX114zHVeqs7onKnqoMl8njO/IsNPgV
lOo2hwRpe4wHEzdqBgeRt+2atsRF0TGC1uoARYOWv9zCK6ZpYINB7AB4HF84PFPA
VLL5t+1Y2a4IBEcnnVtIFDycO/eoSO88zbc9pwfYSNEE8ipBA33s10r5wjd8d4sv
TaAWbQcfA/4wRmuxDqNwtbWzM6j/2LQwlYx1U6EVIpq5W6rgyKkPwiwmN7OyunNO
y/f2sOhHrtEPoizGx2nmiw7+5aG5lwDO/Bv9DNqJtUj+7f9ht0z9mzciOv9Pk0tN
UX+VIS4m8d4iziQpmqOO+EdzEsgstOMdkh2YmjY+MqJ1a9oGUbM7J1IohuVRO81t
5er1SgwItsLEfDisyl291HHpdgZgiQbz601AAKOBaaOlyrevhub0hwBkA8yT+1ds
lg2DCtQoewh0vpdPIg+zYDfEOEZowhvPutUUF/bYvz3H+eyJboF2SFqk7mt4Elr/
COnQW59g8HRzpl3dXafirBk/bhP1wHdbw3sUw/LqIWJ9roxlBCKUmVaRTu3yNScA
EMkgdPeCliED4aI91b4mlCuqoE+BJ5Iu0PG0weAeHpJ4okUIsT9uYAKczOQ/hoI3
k6WJWFk4tcdPFTF7ojOC4t6pgwVN/JxhrXC9CkHK9kylfgfOcRXkywKK2oxTo3K8
sZIpB9w7goKGTCAQ0xJpmiW9i69Dzk1bjsX+SuTicMYvmGlyOMtcOowXi8UwQMm+
rD5UmVOX2OIS5XCF5kVvy70ycmptmmrgJU9C2Rfr0piBfAmSXLI2pm67Hpu83xsr
XfP2MdCJ6L09AKerfXnPFdKLRXzLjRcbH1YYGSC9XDJZR5Yq1v5AtoEeUqRuzwls
wPOAeZWIor3NTWiQyjAnmyvKZnTNksCi80IttpYuKEURJYkG8An0KmczrG7eIEEo
JIoyFsFjGS5TfjxBIIWC1volyFi93GrSMopw9ZrZSHlT4w/IEgQ+C3UqASahnRaL
3BqBN+YO/IaXjnMKsUunK9kNS5ahT9vYnJLwpaGY4WNhS6ztONuX4w6FRbt2YWOy
PtsmSTIGXitpRaKN0VjU6kh/4MNDq8SLvmeGov8KblTDwuOOulEnDr0MaWE8NPnX
lvCgRF2j7nHaZ+GH8+PCYoMgZTqnMxYYFlGBfLoPEmCmX22gCoVJQtXyq/wTv79S
t3g7jP+Vru6xlO9yWHWsLakR9KWTxm0XMpa4YtaZA0q+Q0xw7QeNGfqtodGDbWIA
4gC9ZWdjPDaDwSFeC1ZVZNg5F/T65wnnR09VNit9fEMOFKXQSkWT8th/hneuZ1Ft
O1H9fNpWoHz0ji9ga2U/YhvIgH7iuSNPOI+5BP6Tq+ArkiFVn2VX1/9xRjPSvb8d
LJJ7pJUzatPxoyvFlkjaoSyK0suTDiZjiqflAZAri3yNYlmFk3iRK4/wpN7+b06W
rNuM4x/m1lncJaLBUEi8ZrDcJEHVe4CC6VgCmVCq5zr+PrcZiCD6HVAdq6pr2RNb
dKGtE9xKnOKah3bkGk0PtW78y+YfRgiTM4D+bFPPsEUJkTQ5qHmNrqYf7llHBumY
orwj6T49N9WLWn4DTqNKTU2qqoEYMA13ZVvqRvZXrlg2ubOfKiw3wY82gWnQu+X2
pK9JoDhgYzaUrHBn3/g6fcNjHUB7ByfVm3zml2O5rHSYjtozuq9k6L/a/K+jao2w
ZD7Z3TyavrR4zUaGa0c9v0RerGMOqzamXFTJzdwJzhuztUHD8l7lRBgi+Lb8M1I6
QOZN7QRoHxcHnN6wB8qa4inT7UxRmIu0wgHoEKucGBQAB5fgT/OBXh/kNKdqbhlr
AdtJeLoBmZN30RMGSyMt3gfln0sq7bu3m6wNelEURjXE6C6AeHQSOEqcIUdUHNY3
Sb0OVx1zLrcPaBQ9epoXOG8iOT8IQMM2Y4k+8LK1+Fjscb2SoabCaZeV1ZS1qJTE
krGJ9+o6l6olmf0jflrU5eM2sfiYT97DuPTxD0m3i+9q88jwYN6T+e9VqeqXT6bE
MGSGAbKVFr0uAbqk3FEbnLgcpnYwr37ZLDr45r9wuL2ia6qQOZsbLEESdEGqfqHd
6DnjJTHOVC0+VHFoFj2ceuuRIjcs239Yd+xnjy3uZWS5lxy4c55MQVzpi//Dg4uu
WyaNIKz7268XBB8wMRdSmtmh8uW/qc/PskBHFQa3UgmLdHTN3+yoiv276PFeLHu0
zywArk6npKq1uPnEjXnnxA6ML4aiC71adf+CQOiLgB8WnI1ebk2A79BzTUwdDxMd
FurjO8AR3rRgxzWS0ta6VjE8F3mmaRTh+qtfWD3PKKEhZKomcmRbYsBbBQooARuS
Dn1xoz4olotWodrb8hWgBr/EjV4kxpOS0SXxx4UWTFoNouBp1CSVzVc9pOA8jUZ/
04bz6dpaLhYdSlOSRE6VlIO0asOhCgPNmgjw3jWPzbju9k30L1Xb486mSS1TcGDZ
M3Du+gvdOGrijepm4TkMCjTl5iAcDERvY1LxCNazYrdM2siMHDoBgPhwWyWjXwGE
PVxjl/zGhfaaWLIdoT5Eb/DRtfuAdIqqlJsEBa1s9Lk4QQahBMQA4RX26O7vL/Sw
A1/I9S7xutR/QF8YDKaqHA7dc4gQ8EaMouxXes2W5XHKva1S4L0pj5guzbAz1kOc
Ykyh4uefCu76ReDRY6v04j+lOOfmAJ7qjlSrHGHATbtFelfrmdJOIwgV5TJSlFYa
qUQsnzrkRioobe+VVynNjJ736I99KQh1mKQA2uggwLkhnu6u2wY8V2yIjv+vtjN8
tDDYnZCooLkA33iU6olszQBGzc6JyK6k0OElUCB+FdtC+nZUQWWfJWQlpL+Bt03q
q7ciGFSraUhz/QC1bD2HRvSkOw9kiAfjIrVnVlub3OhvJfOuDbGrnVQSgD9eySjg
aDqibXrYLG7r7Ax0OFACEH5YXfsYxGCvcfDPsiKtlWbYJK7GmhkJkuqDcOR6k8Ka
mpgCw/Ub7kPUCfh1Kk1t1d5UiKf05FMBu/aiRtr1stNp7FHEzvKmflHdv1a7fPS0
DAaF3SgTMfGIQiLokxL7OXmWbUxAsqQBuETCv/YWaSwXUZrs78QURQGu5Gyi+TN9
QY66RzF6aqWtmShEojkb6vdhgdYRaevsDyxh0BuWHi90VYTZe2i/qEUmqzFE1sCp
/YroAAa2RD7fF4spZu205KFheO4hP3v68eFE2kB/oM57rxQSd7viAgdwIqAKmN9O
criJ5YEJa0IqXAFlumGznVpCPMBeluUHzNDmLhTwiK0XLD0pBQpdrITB7F1joGJz
w18WQXB5eQBziOWce3C613QMehhHHJT+uLbXjsYIdu7mQGZmnSd3Ff3PByE+/sc6
qx59DHFvNP96yng/LN+rBQoJDxd3CG8vqsaTNYfND3A9AIMCQufomEaMHCMKIBNE
6YtsOd1W/seLcwXsThx+t0JN1knaHY3wmlJb6wTZZnB/M1U7ycWAAFk5cTBvbXWz
IcI2RuyEmReozFNBry0AYJ+X88XdVS3gmesOfYj0qhCxvg1VtTKqY4/cRkZHXxP3
k/SxjkKazAA0vnyohI6c+igNCNhW186OGGvLtZrVtcqozjxwStOThCF47MzZK2cL
mjL7CznXSHbY0Gv7t3zE26mSFJEIMD0rmQPitcRFKs583SEMX9R3C7RZe5hDZo9t
dkEZL+s7EhkePcIF2OcpNPrl+iH+X8VoJCD0G+2/MGE950zl/mMfUHbxBBv7QE+Z
Rxvb6jd5AlvRy9L+yvB0phT8wlIrMH+wJ14gmNSrBVGMgjNclLxOyYxLwYDV92Yb
2An+UdwYP7oNVhfLEa2j/VOJ9ge8F7iqa2Dgjn9HQ9/+zYUGLNEtBrobQQT1WuuS
4qiyUqdXIJjMRN9HvAtanIqrSWKOAuQHhSDtMNYkbqmeV2ic1pMfPP9L0favZeXu
/zE40yF+YJCZTF+3STy4OPxHBYZvW4oSHuFuBH7PtzVVo0FcM4xYuUxoE+rjd/Xr
vaJd/su9kwyvzvGjbDYaO01hS3h5hTAH7XYoPcb+tB9vz46j1G3C5+T2Huixw/rJ
2Q2ww7o13rHAWkv4BiV+FtDuOshI7kFbdB+0gKUbJWtyezPaKxQ80GyTYkXIHZFS
T15emACkc2VGVQKgww1RejvmbVvdgQ4UZsCYjpFViPJ30qV8booMspo7bTbk9yxR
M1+Sua9KGpbA7U/Vtyj036HIsszz/m4UUxiagZGrz8tcgiivvp8NQqZc5rjVjmka
uVYVF1maKlzc9EHBaw9YvvLZ6PuLMIuQs494lZdV9IPfwSV7LBErv1mzii1drk9b
t8OMRIkhKRPFQFBrwNdYCD3wlijv4QYePPezbcnKiPGOBGgmJAdnYh2+9SGSPFY5
3izXyMgt/v9TVLcbQGjCHD9ckQCm1JQ0GULgtpB5k6MYfFhmaTgr5nK1WOz5scbD
QkL2E/5eCaHUThvOFcYzwWyUgZZ9wDpFoiHvBgtqi/02NHe60Wj7Kbz/T0MqByCn
P0mWPf16HhqYq6NZlu6C0IdrBeoXsV+dUAZT/F8ym12kOmjjOWCJkRBpi+AUAqk3
K20VxBmaTVxqG3uKICw0kkQ0jy5eQcvPak1GMMFWhCGm0q1oVnEeaHwO4MucXBmB
10knkuO3as4sckTcKhrg5ExiMsYUThjyKIB+T0QH5B35gHMIkLjgMcV09yY3LCt7
zwf5sQ2s8xCyrUQtq7GhfQkImYa9IoyCwN4JNCaOjWpxrvnfXU1EXTmbvRY7ysva
SQqpgED9UmiFFjb6Zas+QYjc17w8F5UmGKJvu6W1B6en1Rr3S3WfxcjRm0VOboEP
7oHqFssQrhid0yWGcTeX3/rAtmcdULGsnBP27Wxn007dyeCba8ua+jDBnS+JIw+w
0etIDqJLsIa12U+qxQ5AK0hkhplU4VrEhUeYOgQitzzMExPTXdvRTHJ0MvHOUWpD
iqCRpkvbATzw/9WgFQ2K7doGVBlhx/lIUuDK0C27K5a3W2vPwzR6/Cj4OpdW3PHf
Kcx6IOUbLhIdA5gssI/Lkn1o4p3TjPsGFeiwzxglHJzT4PxlnritpQpzUmaqfvuJ
8WRdcJiV4b4OlHuBEZRkWITKZy3718nz+XhK1UWGGrMgENbJ4eb1D0GSfd9w/zHL
io2PeMhy0ISsXMk4olnRSNSmS4YUopE2mMylCtXYMgGW0gL7rT+TiYja15isI5Yz
yGpmqy8aAdEsdR1jtuhN/yzQ/iOzAkipoYSLiXmy+RF0wsoliZG//S7/a0VMgmw5
lUko3GA07dHDxEYNczR8KYoqMsHnU6pqc0kT0UTd/K10ysVCUY8vPIsOIhXVBhny
QoXRQF406fo9yJRpkXY47b555IyUrt8Y8tjz4SrIrLTXFSwEXPM7LCX+Q+sB9XbV
E9jW6sktulwNma749Z1HjWktR/cnTcpne4PvNWt4Zk8ZqRjV5VTWx//6dpMIO0s8
xIMIfY77QoaumAqqDu1Te+6tDAsqYIE2PXKEpCfjZww9KyVilz1pMbsmW13BrEHL
fydvqANweC153dh4ZvXOrllPZ7I27flksqF5DDk6jUIGEqhKHqvLHq4DagCBZ3+4
IGsJFsQpVW0KSTBdKVA4tdfKmyWxkTEUCBFhHOi256XKOpHUrbVUNkqLJIXADYWc
/4g8Mzoi7x95RyKOydsNUQy89mxZf/7fs9lZgCuSD7BFvDAdOMtB/kv8LCYdTgfE
GmUjb7+krhv8YY2V3RhDcjKtP/y2FJMgE+TE9I/IOsaES3gN/Q0eGNMzSq/ALSYG
3VA8Lkv/xMoN/PkUJ+3pATUvU2owoH/SrgROpRYPqpZw9zTZp28fR/i42g800lzD
4gTES65gDGa3NyiXCZiynIZlSAiMB6gBdPk1hTMyno/gt2Urx105IH9J7THwZlJS
AMLZYjkehR0eYHN7OKvlyhAmT6/91fu3BdQqVzWxYb5iECocZ43hN2mZhcmfKVxH
A0RjCN+nxrnq6cjVdWq6jNCswaQZDl5h2QWaTrMSSy3S3EAupW/Y4+5R1vkkz/jH
kBtMuViVIC+nWDRQHzSZm/yiMLWR6KvAdS3oW7dVyVqBJ4C5whmzlQXa/oVxmHiZ
9MIR5+pxzthrCQbp/CW/7mRRQV48dgZVZodLk9y6K8wUN/KKH7lCTrLvFE0m7dfE
mFKfSl32c5ZMwnjmp/AnECY2lEMFqgu2uk35losy1/a0C3sCy2EN5QlRK3avbHXZ
xHLojSZlMY5uY/WNzmfkgvUXja2XrGMyf1f4a7qW1Iab8Al8lsRDSCmLN842UQyf
ckJU0vCgPofgfOxtTuBnZH2u007pUYHhRpr5AkoPJbZnauKiXeu/TI1oHEq41R6i
QPkpRQ22KuCst7evAgAJpqJtwAoRikJDNAd3Db6CgUtnxzewe6gJxF81VbLdQbb8
GJ42OAVZoZqgcuZTANpV0MzZsGhOieyeg1CKsEQvTH72Cclxh6NRYI+pT5RX0jKL
pUNZmKF9y1DT+8XZx/P/KqjcC1Frxb5Dx0DyX6QrpWVsyybjyy9dKKxPNERlRzP/
O9UDfE7d6dU2hRZ94N1X14AdYOrO5IEIO9jjvppKP73cRim9+aivZJ4Oos6SlWBm
bOzZHyiISvLeL/QiDfAs14elPp/h/7alfLAEn54oRCiv/S/BXZCruLDRb1OPZZD5
pILU2jNrOuDdD2fM8r9MOQU4Rm6vTqGf2PW7ZUpa9czyEFnGjMDv1v2SWEBmXag3
IRbfvsPhrFNKsivH9J5v+K1LDoogcWaMswN9fP9YNJ2c13HrWPlgY9vnZ0gi9E3G
fzcRwCbS3x6AxioSAgVU3UtW1/E3QCc05685+zD7Y06lrrNoXeLzO0hrBHqpf7f2
1hh6yQ64g5fULmoek5RVtUx9aGsN6VIOXupUWKVobbtz9OTNJaqrQ0Hyr2jr66y1
ydo0cZ0LXAdHu4QADDqbU/m0E5vEFqRprzGu8GVXNIuxx5EUvT7vpVNrtQyqBDKj
wuN6WG4tJ5hM5xLESOY1D6hIpv7Cw9c45suHIbObZdx/z0a4PH+C+jpRx7qwH0s9
UOUbigYeMS/IJbH6LYRYCtWIsoBwBCnJYaztNg1SXcSVvdF9OfWgOBIL3FKELPgt
ZYzXv7X9hAfhSQQK473xsOqURKzzY08Wx5rHzRkuiovIEAKcXOeeXeTGwqAy4Jne
ummBponO8F8dnzHv1NCF6hhtKPTF+oXZaiRWLVwF8orf5AwlZG9kgxkl8lAjYbz4
1fB2HnFa5Ie2N08J3bIJcNOQgrhJyWjd9Q9Q4pstppWSHOSaQvhD7vc22bSzHwP3
mnO9yqXBKTTEaSp3POmub33QhY3EI2DRwMKDZoqjCvkzvixEsh9b+9l+OCklJdvg
YwIm4sCf9u3Pe1CqbePS9kAoarJwaS+rwf//DzpazvqhJARDh6/0BYXrBf1xcwmR
QcoPDwrv24P5hu9xHjd7ebObOumXAvBBNnQLt3bTCRID7thkyKLnHo23Oy+5fhR1
UMNzux5QGbRHbIcDYDC9UCFfsCrEA000pKqukf9kjwA/vank1Se+0GAPFm6xa6Li
FTm0ll7s+U/GVjsYph/wEY9e5UaNqZb4dD0ht4R+HyaFq2A8QKzRsOv8R7Qvi6yR
9a1lWVHAvnIIM0Vap1jbtV2PEga0QyUuvF1oK8kFz+pPUEsQoCm6iyJqPlxOtJTv
Dcr2kzedkhr4QsVlRaAX2WqvlmYiwL141bVf1HP8WuaUNEQ+9tONoYxYyS09+hOX
2pYT6z1NwrBOVPJ/1BEU1Eo7aL+CoUnPV9sT7xpVApS1y7lE5ePEGZQ8M8jhuKHh
4sVrYddYfC71zToVyBTWVRVcxtWBf54jQ6cytpUXK9CaMNK7wmNmJsU/hJOvi3GC
JMe2dkFrHlToJ0Z1KtZyEh84tieKbkSVQ7VIt5UuQ1+WAutDK+cQti3zZjSqI4rM
I6G6snqkwnfT91FARTzOzhg/JKqNSffeVFR13KOpnzHh0uThcA+/7GbpVvDP1O/X
BUxZRMGrtEpt63hca/9HpGi6XJMfOUPjM/ib+2gvUvkgk+ecfnGsmGe65KPHJjC1
eMbVupdL16aPbGJqd70y8iiz+l3TbbblbyknMiy66k/nJ4RQbfj6GJawQwTct31Y
/aDgKL2a9ULKG3CaRSzziMWDBWg8ECG4pYF4nku3qlEKU2cl5NdTbY9GsX62O+4L
rDmyX2YCIOpFpFlGSZw4qA579QGhbJSHcjK+ZLmjdA/xQPcO1a+OOppTf1Mt21iC
fp5pGHXzJHjeeXtoKpsEOUJfntbm7UYZb7ZpBpOQcz5HugIGIi2SQJMc2zD2+lJ6
tbqceEMitT3TVuUm9hXK+lRfs6UnERHwWwl6aC/1ygjqqyE5Iuii8Z4GYPiiuv6y
JoRiSh4QoMGchHnBaSk9Pwujn9teq9+zktqy9bfPktP61Jmoyhr4MvtLX422Y3Ut
+M2UUFdVVgEcpnNMg1Dhy0T58hjdGOTYz+WnQpbYzdCHrdhCozny1yKUa0tfy1mU
oBTOnRDIF+H0UJZkG6tI2+mr/gSCnZasKuMOiDxIxLU8jinYKYJ78o82CbkTe8qH
9QGZ+E14Mz9y9foz0bO0SNg29A78l7nPofUu+w428Gia4+ipfCTfmtvqTjG2RBmb
v+sFPnvNw0BCJSjdzaIisvQltGF7oe1874BNJEjAmxSNAmGDAMrYOu9QwjZSCDpF
OmeLDhLIW34MpXkpO+vnZkriS0jAwzRnCNS0g01JA85TtzR03MF4PioZeMV9SXek
/+NRtPJva2xgufhEhDcRh+KmLn3JQr0DEv5aB1Oxk16qc5LDblKLJskqz6pqFcbq
RBrA++nIaKGgAJLd0o6HJ+/zYRVN8+OtHYCb4cG9+IvjRCa8C5cyYfiykuI6+rV+
Y4eTt/8+oJsZfdpNPKYa2yg8uG5tUa74Aaym8giPhhp9Fl4I66gnCH2NdXZxoSlz
bvovPc5DjZ38WnI8wJ51tPe6XK1hTPGFtZJh15EB1+7mD/cXCXIf5Cw7RTv7SVz8
6mdjIQWGKRgZnm7/0JJ0+kniWyUVDZwzz/gSEYEEBlPng0zTAG8OHVLnS+2kSqr4
+01SHaxTN9CZKL4wZeWPSiUlxtS1wkAnM8ydrPi4NZ2JAopVzOXI5ZVl1K6bSmfk
xpiU6KE+ch7QIVuEVWNo2gof834cyb33di4WOI1HUHl204moen7wPiGRP33BV8Zk
E5dY/woVBu04YXKxyibrmzidOF/FOj+DMiQY6qnQLR4UBdGQZKH7SwuUB6KmUze8
oDozN3dxGW47AAM6cQaWf8vmCh8BjwVHg9EmIzqOvJCFWn66pL+d1UpXiOEElwqf
u7d5k9fpvzNk9rYvYycBULTII9Sjn05MNLHEM0lnC0CovyXvsHf66dssjXcNVkY+
656QZcr50tEdTctP9b5vrgCAWBNhS2GCACi4Enabq+zuxWwRuScKACIGHpX3hgMm
YygNzy96qG+d8bshCpyM7pDFhZsH51CBvizwt4rMx3voGarORT3fTdNMqInT0ggw
1Lk51Vut/mzMMdn56O/T7cAScXVUOuh1sdxh5WaW5s/bp30vmyPXhn6VH21p293c
kN5H20kYbqjyKtb34zxP4ECCDJQDb0N1oRQYbChmWrgNgXoKpShLMf2W5eCD5xb2
P9G9jBPMtU14IQbY1LbKrSsFtTNkzGPMyztJbGUtsMj24ZwsR2o8PuYPlPP1Fz9/
AECWvPLxXruqoJS5Ff8F9xad/Ioq6prrE0P+CgyVO+5ufq2ZOoXduPd3j8gQo5Ox
kOrLE9V/6WXZxedTnP9geCz+P1zKryq9thfxrHyHBvNT4x5tq/HHxtKG+hCb5ZpE
9lwfDKHbOD9nqJSskQOAPRaT2v5inkgKhTH2E7jrjOhMSCbeMI6BV0l2SN03ArEc
v7XEPxdJyAS/TosiwFxy+JGoURGWlBpZ7rVYWP7n1UMAQd9aK/1NAFJRcH4mzG38
ot6gkyAlPaYXvAL+NHF22VhXD4Gl205uDmRVqjRaGQpvXGVl65pxnnFXqlgHQYHm
E7s6Se7PmTfTx17v+FR3Yg5DFyPsGZxZ85uQrd1RrgLDm+gX9ZVnqPt10dawqwqd
XcVu5HV1RG64zESNzZ4Cal1bsP1BIg7e1so1NNbQqqm1110zvuo+TMpvVUWXSwI7
SuFw+pJ/2tJqV9dOZTJDSiyNAqh4mgzIz62MHF04jeBBKfrj+ij4PKNSFY7njTB7
Kk5hLzK4/vsPFvFVOoch2a0cTrLYPbylDkTfaRWyRyld3EhENBKhl65Q8/Nw/+sb
SgL/Iww4pzjXdVwvZHyWXNr5cYAq6bh5K2PWaL4744Rsw73KIo4kQ/3Aup+v13Wc
A++Ezrpvl7d+wGuSV9ic53vHMWQf2Q5PBUceRmewT6RCDMQzUr+FEHp23xKPxuiP
Mw9J9D0I1q+dHSPKQKIImFIJ28AtwnE+pO8X12OpVT8TFOFiVC+2Yv9ISNJWs7t7
oWZQHV6hvDQCzBkNalEl8V+wpgm9wkX0j7UdRi6LhZ52qV28O/B7eUIxOkWiBEM7
lh8lLUMuK+nK0DP3kevzjVRxZA/FQK7J9jyoJjuV7aNJweHANPKv+bU/ZlCprEIw
Y1oL+/u5Pn2tIFjwL8q94GdFcIUsIjK62hlCYMTtJv+8t5R1WKjj5Ngvq1WjaFoQ
RdNoRj3n/h42SfRfUmFLt0wuY2zapCPcXpZ441VAS2UL6jVZ58eLbTk71g4ek7Wt
+8MfLXhUyh+cuMvwQiMo2dFkxXQ8JnvMqLnoUVwm/3KB8RMNswIAVCxtMx1iL5xx
21JkWI+DM9mavXuMSniPW7tShQbkUfnPFyb+AtYpcbGz8BB7eC/zjXUXNyq62Jjy
MPelLev8PvIogfrw1WavzOHafn4EMx+wDBfHGueMdfiECIPc0At3rkjQY736aW7U
mMROt3xvqef6EnJbbRJMp1fNkiz99nbZLvxmgqbR6Ob5VgPbMMrsCZYPWkou4On+
BAclXgFjTmtCx18I1c7j9F/3vOuLIhsjLg3KQ6EfPjS0HG61Q79wsiUeDoJwHeP9
OSD4SXAhzUx3Woxymc1v9DL3byEbV+inm/A5UA5SKZkghvIlZh7bgqotgQrLTU2s
Iq/bFrxs5TpU2VrpJChZ6JC4Zb5gqITfRR6n97+QhrtDskTWqQa8Rfr/n6/UW4Ok
dhf6FiDa2XtxbZ8ghN0NDtUqhDOhWXAdMFFBhXki4AJK8j7jtUuNrz1805cqffu6
v1nb5Q3kp6ko4YIfcIL2fXAXHLdjB1Kbcmx/Ve3BkunYmQCL+eqrd6frMWyDnizn
V3doi6phBDka41a11RvNyMLZU6PuFrXqvuTY3hWzWWKoidFiM17Yjl8X9W2UFPvW
FvXCXk5go70k+M9WF/aDrTPloAQMIzVkV46zsvYtSOGYpHRcn0wFH9kJbrXnZFB2
Ht1iv9a0t1ABU5vzgExf4WWPaDm9tbpYEa8P6kyUXENyA62J3WFqwV34lzrwpcvC
63tnUygBwHc18QNjwYtxC4sEF38wBAFiJT5hjGwxSH2iyUs0SClVz61j0QAW/Nkr
m40Xn1NAz57adfiHmWCSmORsNS6i3g14zpfm4NUfuaerGVwTqbq+Cuc8n++eRnSv
D8Y9xWccS89RCdJBsMZjkGupN2F62RS1lSK2b8m8wCtDAEWPgqDwGoz7uEKd3Odn
d4m4DJ4zs6u2dlHjj6DGGuMLuPOyH3G9VGNp/azwhwHCNaBIzvT+0766mPuU55YQ
/m1xXrn+R1AWvNASM5n49qTq7bf7iCuMI0IGtgvwnB+MLgubeQJG1W90YP7+bHjg
qBX08W8tSjTmG6P54+CljLO+TamQYA2Ad+Od5npHOIvy5Knh56V0DA0f8je1pAZb
DtQxQ9NJ35CTQLthlkWt4eBzT4ISEAph6YIQ7TkLHWX6krlPVx+MVDcRaWYoPG6D
pJxi61np06lxuu0v4d7ka6suBzGQVPk1Tmgg1QTX2Jag1JAeSf9QNOU7K5+rOJ7F
3d9sZX+6fA/5bUuKexMTW/p2TVBpqVtZH1VGQCT5i/gLfQ5s3bCo2CZOwd/onvic
Q98HwLID7NjdTAJzkAXBKbgzeHjJHr3nmCSIAieynzquLL/SfQ+yh+k/UBvEtsUm
023dgmDc3P/Fyn6uy/QvVqYbJyNLhxPuzaXxcENJ2nhe6xCFYouQuiuyfq90AYUM
hFauhmsUnVWTrfl7BLTlN1FMfWhnckTzAAuuYm0qn2uaU7IYoPO5lIv0XX7S1BZz
eY1r/WmEnq368OzGpsjTVowjxJSSYohYCGY3ON+gRqmCCEPqtF4up8Mtv0SsBILR
GDwEhB3L+jcIUi1nQyV82Pqjq/wWlnk5v7ddNK42eyoWj1wdQUhZ/vhTVs0O7JRd
j/xjy3GatldXTJrzH3ROWpkvYLtiTAhjLDwcvt7w8iDNbKXOZUdGnHWrLdkod41z
3VjhbrFFT3/yDvkqWsr2VJrXLjv9I7w3hggWhwE1rIQ2S/D+gJ9A+oYDrCezAZJL
H5W6C7t7f6sSzGiFLywh2S4fJ0F5ajCvO+IvlcioLS2oIqW9oXaPRU5TLxDkdHfr
W06L96QHlxx2GrPNY6LqChpWjp+Ge7sXowL0+cGI9AqFHb+TjBBoFdN5OcpftSd4
nItBQzXd12hRj9ZLuWCjxM8nt/43d2tIkCfECiMtfo0kmAdbFXmYDWdP9HsyfkG+
4rLRSquQRJKrrRkGdVoPtr54RqYeLjod80U02vikmQDmFLQCoiBsnCaYLPfgnE1p
1rPsEEV9orLMMy2D1Sm0wHQC3FETkI9X6eir/tc+v8ScJyV7bSq/qcH8sWndpzc7
9om0roUMNIr5zg7//NxDD3Yk3dhaASDBLcg6Sa394DYXFZQSNuOU80hWr+yuVn3M
RBU0nMxcOO8QBn7FAjZe8ILt1RpsYCg3y9NM7Elgl/9xBD6YTRXzsxN6szJqZqbO
bsDPiE3aoxl3XPamdnk5D4LUESvXwklICGqMIk+7KTm9fN4zyAnSbgFZwWxUUaHg
JVEYR2AOKOxnCFzuM0LH0Kzw8zFnlU6oQ2Hd1w3sIUoxx1WAJPshdZfoo9l9ecOD
GIx50LSYWYmz7C9YRgUBuZWBy0l2rbC7cKuMME3vkmHPiCk8GNV7/h7wYnJSbrj9
wAeIZvALlRfNrugvt+mFkQgRbw1qEN/fDPgYjY9VIBnFzeAPfV/UjhMC3OPCyCHG
gh1MUbg8YL5UDSEwne9UGj4b2bJbHDFhrRGXtRjPzJ3dBuDmnLIXf29iWRTaLhNv
il+ybetsNVmA1BRUMmLUFUQ5dAICmAdThX8K7daCuzku9M6F+aS2s0Ncs9ZgQzYR
DqmwkLfOza9lAYQXYows7tkR4Vx8A1Vvyy4rOrbZwMHeSCUvnXuvYLSV95KO4irL
z7Y+16hTGAzxWsx4TgAsRKHg9c3O/spXdyhFMRwEQHO9PH9Ttq4PiEqpuZgx3Vk5
KEWAle0gN0Gm4+azH+FX4F1SvOb/pNKy+mMTOWJBMsrxdlqf+OXPoYXA/JinB8q0
wAd2lhlnLS/LC+hiMqcb/GU6uumV530QZYCqAOt7JRqR1M+0Z4jPZzH2ACjZii+5
0tjjoBmjdfyxZn5CRsDAtQbS4V8R+uwt04TiPyDZwe/NMDxoqqpnLK748wUn/LY+
RTjdWp0Sd7PkDkmjHlx0w2YM49/wimhIhclxjnzkDdzpHdC9DgLnqczB8i+EOeck
IpmH5bL3vHdP5dJZz1wo8Y1wi1ci6E9/Qa3GRUi+lCS441xJC4QF3EPAwnnjHPTb
3saGc+QWUKJ3+lpesnb4XE3a927GaK4YAbMUBk9pgi5r46g8GBvfYtle7pU/WAf8
qToFfmcaLWtazmAMUt9pZamJTC3hOJHYn39hY90nvNJTM9iTNvRkpYI59WArBTNi
jXaHa+LeMcS3hAMtUuEB6AKZMbbuV6jFtVSy6CK1Zmm6mUTsDRAUx2NDs3RuE9FX
lQCYkmoSqQQCO/y3qZU8u+VWxPMMdQB6gIfqJa6ESAglEqN4HRVqaaR4etUAtYjA
EhMDF+Y/5j7jduYOw+p4YiKXMVFUaOAkxYReBhZARVw5C6wp9b7lDJcIKF7I7Zp+
qxSntDN3NKH1Cc3l1UD+RMCZMQ2yL4Pp7NGTsB/A6bAgP2UG1yWxsPT65LaGhBz/
AsTIlTKrE+zRcWtIpLI+il10j79n3pRZYiE0mjVs+5xB6q8SszR6ZHEEDmD6yOlk
jNniq5qw46NtZEKa/EjrM5fjONdS1yHxewR5iEcbC7o9KAWHrydoLriRnHugcb1t
x7zX8b6hhXmjsghJ85LlkqIyJt5pEZHt5QfbC5LL4P3hpQeoR+aJPWsXPdkTEoCR
r5ZmQVV8yIcfVsEVJT2932z/OsehP+GWbnuHpKjNaQ+mmyzyAcSCydCf8SnOxgHb
CaH45MEVL1QIdoO4VhHk3qnwbsgfFvv00Z/pfqXABeKJg4Lx44WCjPO23Z1c9JqY
qx6iii3z1NRuC+tGHpOQ3w3sIWstNCpO/Uox7D8xZIXAUEd3oq6ZW2smQ35zyHxt
vmFE3BeSTf840W6LUEs/Vtse+dEHAYVsv0zJqQSFi2BL5z3PEi9drZ7t4klckjA/
g39fcsyq3LdmjfPzBFHYIvkFIg9IN7n7KHQjbIypUalRnpPSYELQgibTjRyc2Wzn
Cg7AVraSE0+2FXa79Ax8aCsEfoQ/nCJNqw4nyZNiobib3QlUWApJybuTYf89V8iZ
+bBbrcnTMegQypZEk/66BE19l7xR0bUQQQ9cUN3lU7LnzEbNL6oWdD66hnMW50QB
ZVhShLeNh4IU6RKkQafBdFzqEZXf6X+LigR6iYF++gG9Njpsv3/qnqTusX6fbh4t
8pA8t6w+zcFMKpV48ap3cPnJnvq5qqGYTi0wTir1rOTdoh3SBshWGCchgPy4PKcd
Dz5F1nH1S+y5STG9+q4jDjpxHXuebuTYbM16GydafMlaO54fcbXI3x11cHJnKNgL
ONkXLD94f8BJLBueKJmGRQjZimRpc7lE+BIgABVSkbMzN/vjO9MfdiI3P7Ja+V0v
ny0K3G5Wp+wNZEDBO/tpOJNupRnGtMFQ31UhbOHoTXnlXundh0BPcoC+JAw3rfUw
vd0Ni+3WmFzdpf8Z3pdm5pWMzFPctNLfoIwf/2RJp4WidRRqRNDRJRgbdtOakMUN
NL7p3SfapUtl5+U8moFTqZxWAz9d2vSmEQ/8uJosiKnNa+VyaGYLnYibxrmeDZKK
1fNVKuoaBw8dXYGa8RS8FxK2UaZbScJ40bgP6b7Wo7oJCobKnda7Wgl8+JtmaSaY
KWOJu0lvVBOU16CUzg1g4vkUsXpHw0mgi/49GA33DWFLyIidunPKoFfgWE2AXV2V
xqCRJJYqZtclRwa8JzuHjQySsrJ0zk0SCVujZ5eVH+6qMTZshBoMTfC+viXPAhG+
wc/V69IcJAUVqQCRMj1FqGZ4qvmrpGPAHLSUedtLKr123a0wQpbd8eP/3CfgY8I5
9zQeaMEWvMZo4RVFo056FA5S9J+wEBoOgZXBbdGwjuJitW5EavXCmTkJNg0Ldd9G
4TgsIoxBBE9T3e1aaeA50Q3Rrqw97iemB9o4Ibtsu5wf026tIDsrPZ2IQcFmvTz8
Q8J4UFyu+QFIqlJabrywKsTSAbK/Jg6J7c70zwZcH42vshyMJ7CXEe0iP+eV6fQx
y3ZK+7kVc3j1YnWFKvFXOA+PM84tgbpYc8syAe521qs+tY59EVx4smZKmGHFliw8
DFD7dTzRmGAzTjX13g3xAhcix+7uRiHP+Su+jX63ndbzOTH8w0rJuopkI6m38vyq
nb+tVd6vFbhXK53lSJfdWYLfOw+Svuoit/pNv6o8MgEFN2KPO480w5msTrdXkDZj
iEOWhp4l7rHUOH0GWWq2DqO2baHklUaUOZWRBl+3/UwbqSUKwOLiUajF6tO0ui8j
Pgun99/UDKUSWGt3Brg0AvztAsFf8KcXey71HJVu5BChWtt+76kluAbVJd2QFUj+
LY3oYx4vlWDgxc9aJtMq4r8HW8QGF1LCjHsGCsbO/erLoOHUM2iIrB1BO+tWcnEB
7GXFk0NmVp886l6jKjM3K+CwN7ZMY0xxS9x0xmyQHVKI6M/iOyJA/tMpZ9d782L+
YMHIOkN3/bWpsuD8I61bIFYAhJEOfLgdmJOeYpQl8y8h1V+gkxTsGJ7FcvyohkSm
ynjmzWK1glo5hnSLIK7bpDytw3v82pVmS8i1UxGh5fmEGEspCOpMci/ZMZeCe5Xr
u/M6NTRfBZS3O8OefypI6037ojvq029ZoZfw1YWxSHpwOybi1HdcHjJqIxiEIyhC
U/zw2ItuQH+KLt1jwxVGhv5XW78rLVTes6cw+8wdP2ImVid1jQpNCBsGUfOHrYsa
MA7TxER3zj4r7J9nomf5WE1qHnpyXSNWEyZgsA9HTPPXCA5kVwvWm4fOo69JmVJb
NUO86bKsTv3pvIb0GcylOtaARiZ7Q5bfpaQlZ9Y1iZxvAK1YZeybscu42+JpDh5c
3Fl3rkO5j5LIKlfljojcrw1NOCdfzUpSLWQ/ZPL4w0lXm6sLB4P9YYqlkE9v3PZG
hskOMny42OIIqQVAHgb6eOKmAzgEzLhtFIBBFpdijnQMz1tH2Sz/l8C7i6GeP5FX
DINtiYSUZtSziua+xr4g9fB2OTjbBsgn9plCoLUOawfXadH3V/MCpQzgW8EQ9RZw
BOe0FykDs+/OzsFk8QIiLHAWPKprpi7WkeBaASiyQquZdAzChQetDIfzuB+lgnFL
mfTs8lYITbDxdUEAc8V4q4DbsiPQNJHdVd23on48krU7/v5XcDdoVVPEA42tVqk3
kl2c8D0ehCjoHY1Q/g4c7TBFJRHv4OtVo7x7eu2xblDeHq5+sNW1UxnJ3+VS0HRq
bdEcGHv3maJlJT3sCfENzw6qJd4rTV0dpAZPBczY9YGbRmFDNK+gZgXSKX+BkcBi
05bHQsnvqcshyX6uWhV4UV5tge//uTL0WrasUhziAK4TK48OMeo4SzZ18mW1ve1X
8p3sTXkvvWZCO/jYoJ3KKVSbyf2fTl0CaWb8EVu2ncBZZlGSoY6etyOSCxlT/itr
7Qk9bRxZP+Z9fruV5Oz94yeebX2iytV+lPiCn7LQN5XbkQ9B1CCVjDZ86X+Zmvtn
0l+iEet2MQqGllu7jQabq3Nh0NJu+07GTPNsGvRAg5IqY/y55t0IVRHxw/gGgRkR
EP3WaWxR7rV+GWtnSIZmd90Oa/WTqklWlDIgub0CF5xo2XKevR77svMitr+CBhmM
5kil5xbEIFj0gI81rOZxyaTUSEg0mVxIH07Qnbb8gJLXBnaghc6cuQMYw/kdY9kg
fU9ze6fmsHi9glKemnBqLfmyFOtTA6lxMvieQekev3Cq6LgbrVXGktHzZFF3ZuLD
ZUU9x68LdYn/zlGuUB1USX/eNbvHTcc4Vvs8Wt19ichdoa0HLmrcs7q7/8KMiIcf
q9mDXpdwuvFytcXbOkVc0+oVKqdWrxl7WUlrvkEKhm9Pmf4jtPpdtqZ5BcTXUOPi
ha87H34Qsn2ZPJ/HNI+loPHSgEjtJP9fB+m82+D+0Npz0PlLtj+8NHw+Bx+9BW4U
O5PDSzolwZSDkHQmf+CnEnNMvC16jpJcrLSTE70Q8OvvR0ytWEBOTHSf5isSmGrS
+AnpNqSj6bFxe12WRIjruffY7APJC0yrFXgymn6rXbxk2jdcb4NI0jdq2qd0dgg3
e01tNCrLTbiss8T6KQ5C7mfveoZS6RFNpPEKRdbsBQtoF+RQSDAgvAcEFIR6xN1X
kRYd8t1Tfe7ICwJ4qEh33Q8tI8OsKXsIMxc+S1f+blfaZDdF9loDhlIxLqCH6lI1
Sa2+gBTvQmEcHqJ17KOts6Gpr035iLFjoqxCl+8VWC5aOv+YIkVhcc+i6ezWezdC
XkwYbZkN7oCr87bg+swCsvMoChejKcRFI+7hIqJFqZanfvr/PG1kBG0UNZ0zPzh0
yA19Ekz81UIqBjAlwUL8SKUuZ/NrVONS526pFSHNNLzpQEkmySDBwiBlg75Uvkwg
ligRi+KTw61CEw1Ki4KEfkDXxMWGef4jRjiJ1fuMFFvTwNRLfV+E8Qby2GyPSOQm
Zns7dWGuZbrklty1D/37FHf7rIeRX0dWQbiowpFtnYs=
`pragma protect end_protected
