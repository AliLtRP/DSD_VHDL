// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qp5EYce40bSnu/H++y8iRkSi0+v9wNUpYo6iSLHwnWTzg0DloYiHUEAENlW4B4zC
0rbEaBDy5BHVIlyiW8UmM4pNVmbFY7CUqDvnMYPOQpzcin+enDYOwCV/LpB9wuQM
ef+W2QUFYGgpjz6Fb+nn05WRseGlZwn/vpbNGrkorNc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5952)
0hqYnclhnBofdbnzU7yUwRh+Wxt6bGJtM20MOAjKVlw41MecAnPSat5BMFahbRvm
wflOUcJKpGSCex7dsSecFZVKMPutVHo6gfqkoS1VA0iv/z1ECld7PtrJUF25TPL/
PVOROd5+EgXlZ3zYxUsgO1X0X13bcOyrSdGY40LNmLrkndzkaxozFsk2Ee8ntagm
oNjyWuSGt7YXBFgxCbhYtkFhv4S5LevQe0LLfJrmNg6IcPTF/3K+MpF+hdNsucgv
kx8fnaWoGULtSxQlPGmvpuFeVvCm1LEfsra505urIab/4Gu56QIlfPOEe09OrWwG
/jGakUKu7Z4ZFU5OKodCQCJgTdC2NfHDiEmwn5dT/aR6M/d77ZqJYHqDirptBPQ4
jGF7H0YO+MCmoulOCeBR4WKD3C5f6GFSlM4BD8SmoR5KcvsHuW5EALefbJ7gAb4b
fdSeQu/gIaxh1Vg2SIfsnvm9nSxDUTTiCxozgt8wqtJ52j0q304tEqWbmw7ELgS0
qafSp07X4XcPxkyWOPlQqExmevgBeoG+YiVP8EMIsgyPGOS4gXpx1wZmzSkHH0Q6
W7fqZLAPR3WIyIL6TZb0jBvFQkwnkGnjR4yqfwzuFnQw0Nhtecyud9vwNdsTnPqT
45Xm2LSXg/cG/hQ75xrUP97i2eOpCMUQdVPZzRe08tbGfDjJL0ntvCk7oyMNNW7z
MQO3Rngo02fZBXo29tlhsbkvWmphehN9pTMIZX11y3CLIEVfjwcFnmm+rJ5mJGXh
KC3/ozhyby/Kf3LMQIwsaGBZ3HCzEOCJEwyWpt3Dc8bcoU2hRjYUwvRYiZrVN5EV
ZXSfMwbd6ksUek5f1XEAs5ipIsSMzFb8fj1uk5At46y3w9mNTsTZL+8839ONv6di
l40R9nf+CoU7qDTL4Eacs/lm91eMbSLzDhZl3JI49ruDqixYpLymm0R4X7zoccP/
NWTYZfK3ZV9O2hBB21qQnUZslBJIw/JaTYSQr8ZeBx1j2aFAy5j+Rr6fqDVHbp1M
AxQXrgsoMv6R9Toye9L9jWsc17C7tP+pnDBN4txtPn38oGguQ53AeuBoGt1XmX3a
PPqgrN76cSJeeySI2bhrE22MuQ3LIjQXfBgljB7K88NaS/hNtnjVvNisP8pmtbxU
MWyF1qtHUe9X1fUotxyRst1MbpfTWlKohyGq0Uh3fwyHVXy6JBqAvwyup97XlORA
/rJV72ec2mkyY5wV3zNYX01LJspkk341L+/HO9McBj5spO0sNXDHVHH3e9jnMMiG
29mFSRmzZpb3l2ELUxQlvB87eP8ipeCJRtqfIyuZ3qHSB88HgH3/YNXT548ReJXk
4U0R7y7b2R9zyko0WforQOCKInniEx2kAV16KiUgFa8sBXLppGdS3hMOmNinimcb
CsDaQUaMPUFzHhrUnW0emdzHydHvxUO0VtZZdoKfI9povrmDfzysLDjw6JdYF+0p
XZ9CBbsMQXWbIuzMLRdcUx7yEdKIW7MLGCphlMoZE3XkD5+Z6VGxtB0pOUOC2ill
BAXsKNI5qf0gJpGWerVm5gPPFUnWkquGcZ9IicCO5kfMjO9eDjDrrEuEnX97+hi7
iPXuYDyci4ItN2z5yjhGfJjPiUrMmV7CHddf6u5WlaDOcAZzrhJlATQEiVjbZ+Jc
zWsC8hS2HKDY10Jve4W/KmpexfUDv4j0AZmBiG74JWnze5XJP7z9u/vjYTozGgNe
Qd2gnpzXvn+tqL/48RTSswZu7a4ShtFC9LaJ5gmgTR2YGMz8LSje0yYXKXn+mXyR
RaOK73JGDr8fqNB2XKroktuEIBTKPHreKI18zlb1lrS/sMza/29IvWYy71jk7Nxv
KDCdfjuYs6ymgQDHVLOIqJ5MvoLXs8TVW9xXM28ccibVAXYXCokuAhKs58pjLEsw
XvVry/uL/zHsP5zjNGz9MnFu4VqByalPwKeBCR9sCHIX1/CmSs9vp/OjgYyha6Wn
HoI8j/qa5kw0cSo1R2QgbOHSiys4s18BvZJexdkyruYd/drvvMOsk0Hl3EHi/D5b
/4Nia6wip4VrIR27+LNg6cAVRCuw4vaiXxvM7zRzvU65EjRJNyUTKoU7SK5Ei72G
AEVuCbiygg5poBPv0ViJYmfM5JmR5eclhKOL9/HVFYpJFRPm2yetOLOYAg3HwIz3
B+kpwhPOYWNPu3enevcGDhCJ26qremFAITRRN7+5Ykf+ShjIqrBSBSP58scZzwvO
lJRGULsZ+AybWf7FVgtjvEFPjC9y6GXNCFzEtkuBQ2atQo22tEHviKRTkl1dCbPu
IT4QKBgl7JRrKk5e/JuzRcA97RRZ2wgn4Bgc2FlJ1WYzIdWdNnLm5K2dfzlexuk9
PxUNpT6m6m8Grp3Sv2DNMSAtoVe2N5Jzza7oulJLNF1qsN/v1ppcnxlEi5mVSTl6
2cnENNup/k5xMxywOaRrQWa/dh/G48CGd7vgwL6lHR4b71OGKl52g1hnzS3gOIvv
n2YEFsoUXE6xLJp/nryM8oHNg4dS9vZfMBJqIbfrRYPgOpgh110BQfyCUKUX5rzG
yWehuDeVSvw3dsE2YxG5BcqFq63X2rOLQMuUMtoxMb2sT496XnHA86hDVsvzxpUV
DZsQHEq0qy1fNnKqJEXplu9AQJ5op2o3cobTyEKRCk1GVXd8z5HtR/6w3WK/5/89
GEkPFRj1ISJ3z5N1O6kYkvx0maMVmG+p+0Ko717c0eLSN8JrQj6p0cMRc68AEcM9
UwSfYJXELdD4SHl173DS8sWJpgF9svWUoRN//c+gIb1fSGnIbvJxOe8+l7Dab09w
kOpX03W3iwdZOFHx4ASNIKE6W0Ac73Yx4jv7PUrC+JwDGC44svT707bx5Z5uPDZ1
vSHlluVFnRj8bPwwewjsvWka2dxRZsTvkWuKzR/i2D3g6G/ACFyspH6TD+mepdJV
3PY0lSNVAFmq+rDA0Z+R113nroSoPX/3//wT8RjjRo6XjZdC4FAAwvrUSzJibQTz
LRsWdDhKYJOzh+kKIxbLqHyQBdY9+LmlIM+c87WFvHazHZCkgiR5cOKIxoKhJE5N
+iSx98MYGERGY1rXFM5HUUnTdXZgQjYT8jF1u+7IRm6Z9vBCG2/OFxQFIgMbwU40
+ZoP4yCE0Ybg5LHN5fGNiOPE+q7xyywFt8QD0E9Pn4ZnYtuwkER/qNQ1IFGb/Hxi
nLMv3oRUA5nEUVw+a35gnbmSLo7LzIrTKXVINnKmzLTj6DclCDswg5xUtOcQZJ1n
qGi8uThC+a1vwGJoBcWathgd2pGstqd+lHzl2ClF39FftW6egu4JQhm4xDt6IRWF
zsPIwZtUwvTp3s8htc/PY73NCucu30E8JMjMEoQ/P78JpOEFOmEUN+41kN8CiA1H
Zqos+u9mqsHJT77K1FnaduOfBTvSTx53iqIyfkldLwlcaTRFbD25GdO2/BwIozkk
x8UNIDg0wZSPsXWB9QXaQiMlkUg89Kk+5UvTR5rPDscjxxrDoWA9ZY/Vnjy4VlTA
FymMA+U2IvFMxSkhmphYRUW3k3vEH/0zX7dwa0JySX4NPvjZCUDAfonm9L9OBs/5
pTHSfx0xCOoOgRi41OuItIaA/2scwFjNeKHvxpYXPOhHGYiUOK4SeDni4Y7Fpxs+
Hnu323jKLtli3QYM2BRMTQIXa7sBYVfKwJrotXk58GYRYQF0JHLL5GF/YTENne2k
3uNu87UTdylNjROAGTO71t47Q0Krgsy7iNMnW8z/LJHPaKHDlyDLXDR9Ik2/1iQR
aYJfxVvIH4I5GypBFCALgHorLCQxoJMXbZkCKTtXArRHxK2FBSMq+OktSVeKZjsR
8Du+T2YMB3+J9Wh2hlq55IYvqkCyVSkuRpkrCM4rMGs8YkTYVq6dF2Ig1FeixZQf
pLgtSDhhjN9vwrWGLFj8Q1TyHj4HMadz2Nr34KPBKwm8r8s+TMYxEO2sJ+Gw0Mta
Cn4Wd1VXjN2oXRXeuNVALqe32NZrIxcBzAmiXtCRoD1ro7N6p7AL5YxjY1ZXeODB
NG28i/3dRaUmpHEj0lwByKkrC9R/kvUiI6qVKEQaUY+6c47ZRnjuON4JkkqmQyzO
1mQHsZfENimdIe8JmGkEdJWMEN3k1JPV03RKeZiAgOF0kCnr884Plbl0+5Cvsuca
u+PTquKkoTFUgrUzlJehXxrzB0dcnaI1y8ScB2gUgRezVR3QwsVLukDvzB0gOl8+
DaNXm/z8wzn9x51NxRCSFAxj4pjqgO6vNBHEgYiCDI0RHDe18RsCRRwakNQCGJvL
1zX9s0W/gkx5v6SxpZtGKjNF58D/rPtDMurHqNY6Y1wQr/MEdIF2dmQGmQ3dsMA3
+Bo3Jk+ZfIyp/yZivknmaMuMIgiju81Sj5LqdnbHvld39XtZbjn1kOyrV6/rXbF/
NEzMXTF82tYlll0i6gtd0cTK887/o+hCPwdxWcKCsQqjXZ9fhbZg5rSGYA2fC21N
Sbkhd0oHlqpPLs7ja/GbNwxecE3lLdgpehlScgBkq60Lt+/zdyAPHeUwBjlanATj
XTdTvK2+Worf0tk7tq/Uoc+Xt8AS30TpUmo3nzOrJ3/x31mkbakLiIOxk15FXniG
eA8PN0ue6RpCJmAm/+tSPjag/lnu/sSQWWUNT2lzMJzSrexdeVgFjWmtaxgZZwLO
ajFU3jtUzsOtV0MAslfN6BrsbEIydp7L33c++a0sj6UG2KzO+0HcLsP4EnnA/KFd
ZKFP8KRgnPF20/b84+w7Td8jZ6SN5aq7Qj3AbTvRBpFLDpBWF4Au3f72gMN63PXs
BfD817wB84lwqcEHMZc/n+o8pIoaBsg0C7EmbRh+aqD41EW83nN2V6Pa5b7kMixF
bjts6zJ+JaCC9m6VmmM6OzxgDLoart1R/ysmV+5bwaZzAwOojsacXtSSqSdsZl4p
jhxgRZjQbnXrE38bGuibsAYosVUn0qUcd+bbLGKwrss2IJUydXpVSRwMC/95MTvT
ZrM3lX4Avkw7GiLG3IAHv+bw8JLRMJ5O3AmGfLmRz7pJwZBKzgQvwAZoWE17Jid/
3zDwTjLFyPHoTq52HywGj0o5cwkvPIr7ekHWaPFfHfsw/0FIkAgNSl3CUpqr8bl6
hWyeSc/kSwjuQ7L/SFMu31/VHsHJZC60htAu8ye0RkLs/6xr7b2bjJAIsDiw2cvT
MHYlhgKqPw4hi6eLS97lBgnN+6F6cktmSZm+vgLH1tTMGwbOEq8aJTY4rpmUgXOh
B7rpUfWDA+3NezgeW4D9FBse0roAv9Szf9uo2JafGp5lzkAjqDK+LYKYPOXmGqz8
tp8qejw5R1V1ltWe+P6tL89CyqQXNgk5Tiqx4D4XmSVPSOX+m95blzc205Jb906t
B5GoF+gnxH3drmPQCo1UNQpmvyqa2QJfUgw6u88V1vlHr3HYnliMTjuwTX0HC8J6
iU8Ka0c0KBrz70V5076nyf66nRSfPjrx5RS+bdibWuHjYg/Bx1z6iL5AJa2ODdTw
8jt1Wmkx9qmjSFRPcRcw2BdMqLgDHfOvGSViLtjV3CTHHbS7yhK/irFPZfuDlErQ
otfdXFhpD4leALs5zB+VgtPfdIrliXA1nu9bcmmd/Virxh+Fr+2hrxmdOY7b3ZIQ
qmb6hA/lxmH3rSPk0GMmAS0MjEIkJdCzyVA8AahmV6yGjV6eZndErveTVlnZOtCr
YpY392UQ/IFr0euCl5/K5FjYGQiSKH59ipSX+bkHzWZ/TObT9zKefkQHY7nmkEVk
ofIjm/UdZY6LU7Ul7oxDMZwrksfrU3WYWYrhw9W6+o+qu1JTfmLqA8s59X9EKhTJ
peSsX1JVzsOGkDLJQyg7GDyMYeVQaI/VO+wpgfF5WraDNNKYD1XhyZzH8DP/Dt9O
kWW3t+6mtOwncnHKmzclIn8S99ocWv21E7muo4gxaL3tZhtcQ6IqMxLEZbNvyxCv
imxB3wF55JpyVvNX9A7wl4vTKmA1q/czN1fTw7DyKbKC4qSFweM6YcWIbxUWkiVK
2BQgpZtNopfJQdTsEf8vwwMzGxVVQCk+SgDhtfXAblZhLtDuGq6uP+LbwLVDxzKJ
0RbXVkn0AvCoTPkgqokH0vraPrRqysSNR9fNyjGUK7OMoO0i7oKHS8/6X/y8trw4
4fxTWib4Iz40BZXIIqFtbBztCNw/8+LvcehakiVhEndfTjFzYY08jt6xC5heJPJ2
ArSVSLlSb6FE2hzO2XDjjOzOgGsXZZiUmrJrecwG2rYldgYw0dGd7VRA3VEZ8QfL
/V7rioL3RIpCgNjC1Cczb2okg/shWZQucrhx82kTenJ49gzDdk9CNem1Ud92iJz6
EiEdnW2f3FVDVVKE2ARRq6bLbDMqm+LwC89cQlsclo0dnoWgeZozLqGS3kT76/D4
QnJFN/H/L1jol2a7dwuYvfFf7GXRxNhR0tfYYj6+LlE50vFt9gMz4+XRJRts62AH
kZVwEtkg8FDbFKfS2sPifJseiMB4KJkxgSJg3hF8fuKSI3mRwhwDNn5ny7lIijdU
WFL8OHyL6XdHo0+bq0wyjFnkJ0vB2LnT2OFiXfUEsSLRqvGnCCysUL8GT/HzZ6zT
Pq7h1lazAVP7c+qxGrM6ds6KTfg0bbXaWK9CkpC/SF9JU5vKbdOs06ecxsVBbQtT
nhUjH/gKruxYs0ozMsgZZWmoBZIXDM9cwqv8dxodQ3+oT1auVzaMTLDnMp5/EkzE
ngzsR3eLkR642jYhasvFjibp7Mq2W18x6N+SOieyN7qxAA386/bX7Xr30MqwWgw+
MOGJN0QXEuNplpU5RvOSn/9Hth9GGLuoKt8zrDqe31M1Fxv/myfXOPwBus37LNHq
fDw37GfGO4hx9swLyr9wac/L6CxG1OJUTBG2dUAvzYbSt2jsYMMVPAjt8UFM5nyU
AG/8BMPu9RWd1FSxcmWC/+Z243q38ma09MN13tsRIE6nT+I4Ie1QWRk9LEm5eRU4
kJkMlbG96DzYXm27NaE1R5pW79yuV3/vZwsjkA1zqaFCVqs/ZEmNubIL8R95dJGj
HxoHogVVG8L7I6wQyxsuTxoNisCj0537z/OZbUgOzoS/qG/wpnE1z7SXyzWIxp7/
Mg7UUvrvtCOZ2hGZz8fbR5fWjYfTpLb/BWJmGYHbQkg7MpJ1YTIcQGXDyO5wgDnv
PCXbeRO+v+UyGRkU+O5sjspf60FSx0Pw+3RRk4QTTEEeBGF0vc+dVtAn4QflugWx
69dbDHphdO4Q1igK4G2gN+kwY6uAX6ZqJLrvi9cRRU8q6y2lFRP/VRskbsQHBt6d
vKu6OLWFqADdlIcmuJ4lM/os7PVyyZycHng8dU80MRnxiW2YoxNtKHf+Q++im2cA
exj0KE2MAubXMzv4C0HwyFI4PGY4Ld1rQOvm4zhKUON7Qbv2ES7xJyd5yXDknSbV
h2EATGp/eBTc763GpGkq8qoYMyNHFWm7sQHJdYr0j3/lwgfYJV29zuylhk2lupXU
Wp41PQACHdMPmdtsHrtbM+W2WRl+1kQSiQsFoCl8Mh0rI50fBDYnSkhwYlBWwlZ8
tjAkDwZnAWQ5+YObQhM1qn1iu/faG0mHxmAxxW6ratxjNrSVN5frkxKot/XyAmkJ
CfJxM++j4Qe9FZkun1/kI4yNHQlEjhBTltXbQGXyJHnXNxBd82Q1o/MBLJRl6iuA
rTFD1LWbsmJ3QmrWfveto8CaZEzqtQQ2OSm+dPsZ9aO5GMdhd40PzfLeXablQMek
L3RW0qRsdGKa9gC4cMesrosUcSOky1I7QESKOVhwAx8jqvM1/wwG9NvBpHFt7O0r
6ZLiAxdo4CnDs/s0/T8pUx50XkOQj6PMlaMH1dveVoHdO2p8DQ7QIwQOyGVRSbA/
DOTHm44QO7JNWaVKh2WY0iwkDEaFGnEwuFVctWfYowRj1G1QTacRqFqmNcVyCkQb
`pragma protect end_protected
