// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k2Mn97KylNEqxygoY5x9MeofNsffuPFftw+ZZBzI8yb1Gu+6AkjgFj5hWTBbQ0OO
obcO3fM8qzXesSeDrguka0lNzNFolgm7ptz9MToN2GSxrtrXhvQUXsvdakyb3vWK
wvlsvMLlShVJdQ9462hvzphR3pdGF0mg498P+p420as=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11600)
n2LWu/kaqH0IWxsnrfVRWy+Z/3PZqv9QU8ohetXCS/zO145sBFcxCaH5VUgBE0dQ
Yql1cz76eOvUOQtopD8C50EXmFgaD8VcibKVgQDkPFaGh6ZbsQ44zvECPdUzIx1a
QB3L0PEVGpnt8ILUrBDwyy3nPsrB9z793elbWyc0QDC8WA3DWAw0iiB6L3a0pAs8
MODBA2T2+DfnN+K8klwI1lX3orGZvdJ32SlM0pzdHod9hnuL8fET0y47qCsL9i7f
9ayEDDN9wUxFu0gP26ztnHsMfRhmPYE81W/FFu79aH8O9z+XgubYlDSZeIgqoYXn
+tTW/Zi5EI437/mwCSFn0cLTsRjLvEH8QNbEEGVTCBYzNNNcAoByoujt/3bz6z6O
kvXHko/Gy0OOJ1IqxkJZohkDapUyRQg6YiNXJVUnxct6Zw9agooYKzkcnr4p4PB3
b/vFwXMDFi7ZUsvDO0ZpRBLzeZ0jyronBKFWpLU1Wl30tgANBKsmpclxkJSlYVGP
vv1hA/k9vTynETK+gJH/V88TO0rdiA5GivIT1FTxTq+gyZaRbo1AMK7gFU7pv8vD
qNRhin7amyq/26NpkbpN8EO+L1U3AsEPtbXP5WZP7Prej4pRO9K2ng4H1CKGEkEW
vmbBRaij2V3LhSx308dEYJ7iLlxnm9aoF0L/wp87J4UwnUXhFzjLnVU6K8UqcD9x
3H0zq+2k/XHdsM62rhzdBe1lk9XLWjX9SHdtsHb4DAWUmK9kcAeKXv2pYfJnUXlS
BCG0Cnrwp5MUWWXwY4DaYOqIeyex9CUsFDSAp8ovCfZOqem93maJL5y9Rthmn+V1
h2BjCuOu8H5bBQr0pxuLgCBSiVvV5M/cn1+i4dsuexW2yFAmBTxBVpYEMyu+xjtc
b+xwtCbDuDUwRu5XoTd0GJNlWWI+VoXm5st7Yidbn4leANljBJRoVWaiwlGyWe3N
zK0QMCivwLQTA/iqwzN84jIJIq8/ANMwfmveJOIrqwgHHcDI2znOTYJm7BrDYbwj
eCKZ4/x6yliywKwvc4i0boDiJHKjJSW0ZF1wQL3sl9z7kO4EtXJNt6tfKMX9uQwf
0pJ5pCsI1lNH3D7zviFGtmC2gkDS87J+oYDEkv485S1W9P4hL0ip1rOeABAtyBeX
JDxKUKlEQgcLtd7uXg9EErc4+M7878UMYhtB/5rRVbxbkFZpyb53q4j23GtqqCDa
vraKB5oVbu7AbflQopW6gAy8IJhQxNU/IHpvWHtSpPzPZHEGLat6JTodQ48F5o0o
wUqd/ezljD2TNUVBX64pv3IjAacrW/ZMvhTiMI/q33lHsHrzfH3yCSagAJtdgpBT
csORauK/klwJdiWs8dYhwyO/OPPTpM+xy3Y+JfTj9VloOL5HceunsoJ0otHQnd5F
4XIMUsismbFL9Svms0d9sXGjHcuc77pHRx0U1AhyOm2asHyNzV0F8GeiVx/hu6OZ
xvkGbvn13r3LKTdAf3bHpbmNe2o/fbdKG0JB7mtoe6AkTIgTiwqSVY2dnLhxUYo8
1LwXEsEYlN/Y4lM6ITLGvJMyHlzGCcJwSW0ZAXTV6yo7c9GREs5ueMWA6sLZ9Tcl
562CN4SXs6K1NsBqWlpJUW8K0eANV+YFkt4nDEHFPHYji4UFzogcPis0zZkao3nU
2r2Z05LaZoer19bMgjZkLa7VreuOtYjuldPKYl++8+zOzi9lRy2Ctx7RmfVDcl84
2JcLDR7rbFnA1POqB228Yfp4F1Zjxbcfwrll5ZQAF3Cppyt0NOv+WRpsXtJfkXnn
OCrVZeyrs+vkloSJkarJ/Rolv4EZj6JpTG62PrRBYOM4D3ZfTiX1T+gUJjJ76Iw8
XagfrwSPI8JzVKWVh2TGNYenkuE156dzTHz0V+Aw88l65SUFp6kqpT9CESas3oUL
VC4LBw9uhGEqEM54l6UWa2RvlQFuFpUrQ8goYI+Ri8QJVuDU04CxEuQ99am/9hLG
ByNLxrwWyWzcaUKRgBbK7zTOexhR+nQWpPIcg/2/CA6gbuUqfncdEL2WeFUU1TL8
2GzPBPn2gNy3cf3ICVedvHZDh0ubBL+i8Y3oGOU/k2QNfB4trmGDZIcJY6HvG/94
ipcWs6HabMHqmZHBJaUV6rGkTzioStDqFeih8Uu7DKvlzp0O910g/B4uJ5evGiah
kkuPgRqtIvNxnKFuOshQSPoyRs0Lk8Sdh+QuCv/I+qAzMU9T2+/oGvCJsdikEX2u
3mfG4Lcw24mafmyAIxc+ssNLYtjVrstpSUotUjz4eHlELjqmGZlA4igdWIg49sVb
Syqx8hzUDNSexa3z5oHtBQlsRg961uhC13oM25EV7JuvLpVZdrWZvZ9GNIYKrdoe
Gjns1k0KuSPyou7U/1OnOZ7NgP8MN+RGJGKhLjaJKjGL9wDVWB0MKX5gQ9EEpfiN
U9BkBq1mFQ9D3H0+rwfZB72jFDD2eKA9K+jBNU5ddHN5uBhSAM1kI/n4c6kiZizH
s1ANL/IKgaI4P9KNzVsIDO8q7rlT5RK0DdmuyMHvXv4R2S2Mxd5m5quskLhUA7t1
7I5AH5RjZhfeHSI3yhjK5zKfptmMiDiENcKnKC4q5C8U/qFv5cVo4Nnm6Nf/8Mj4
ncRxRGnMV0RG3h6i+13KbLQYCJ60wa063lZHwkE/NlEdxTjwCiQ/jfqKVCEOSqfm
GP2KsuVmsYCEo2VQTjYkMqEzSahwtmf7COzxwzI3VEK4rb5Qv82VjdKxbDqXO0Uu
SimeiP1+G1Q6dftCowzVtCIYnHnM5zyhbq6ynbV3CD9FF6E4DyvMXzvAVdpAjuf2
CZcgJ5zcd+GFh919b8BBqX511Hgf0QhRqt8nolgEgHze62HI5Kqd7q4Tw/ax1UpD
ibzbC+/8IONmEFse5DvG5OhX40XqjstJk7ELxRoYjSMNHQucX7XJ4+hgNn57h5zX
6n652ACXw9/R6EdAATcCTdMXoFSNbMLbRTo2otGsIvs+sdeYL8s+yEeGzkil3BIE
XdFXHKO0/dUr0HlWD2AL51oNOHGl+xzt09bs3Hm3OTI8OvJCo5sW8MGA6w4ibDmI
CpSXalGSagAeIvtHLzH8rRcdEP6dVqAE0SL1NHXtLLaPJ20lOSmy2XLT4ppoSRJL
8eQ8dicNrJVtEr/vWXvhl8ZvlrSsg5hRCQzQQOjkhuon8s8zC+pNtktlg0nWZ6Cr
yjCxpxuLexNUalfCiglvKGwjGSMxsqwQWatNSU+dmrfQlBRMDjwe5V1+sE+Um0Pv
AsWHZRoqxDV7nfZV7PWrQ9iQAFE7pvCnuhjQzH6wnbBILHKW47H9i7fd4O8XG7ZM
T5zN18Lf+b7Y7fMtlfIq4AUDAGOyK7Om3XMy/e8RlXVm2a3YtSsWujsv4oeHeOuR
MH/8jR1zavW3M34igvXq9x/enedwfysOYs6g3AE5pKQvhOochc41aNND4FCnkhIQ
HVvPnWKKdm3ya5oU3Q3xPW/Fdy6/Ea3AdZgzO3bDYKaP5HAubF4bVRfycv7OCHib
btrjt6PG//F8ao324kEELw/4LvivG4rahU0MpO1Fry4X8rcTL43oOAdM2nu6Jgjo
nst6JjCT2xxSqV0obZkiY85okJ/R8oKF/m24o/umznYvExi2XzHOleIwDV5qyFXJ
9slUTtORfl2/8JgKw60DLk0sXvZ0Wld7OFvuygQerXp0lI/xFxGsU2wSRpsRnLiz
WtbJ3kmbaJtElne/f/v0iSKNY+rzxDnRoi8toO1MUyVVTf1L11iS7goP8aPRgwa/
IV6V5Fr3Ts40Xk0afm4o3jzhEO+4JuM83i6aG7vk9TCXXhnxl4lBmy/XExv1u6cx
F2qsEec5Dl48p1/5LiT9MuKbZEseJn+L2FHoLgU+MyWXCpU6AS/Mg1I8/LPySe6u
j/ImaWsrJ21mespHWDcShC5kvnBgrdY1SPVqutzIqT8zLfQG3MwLIo39XFZz+yWa
3x+QC2E8nTSUmd9uRX93mjMOEfxPH3y+UapkVsOrxgRvoYvFSAT2mK2Nsc177jtv
+ul20KG2l6J/tZyKWNTfZ3oKF736nNc92/dDk7eozTz+DM866VM53vH9umZZfVLx
nuApDtMin1eS+jekxmOz/GBDiCbBOB2ie0np/1W8R1kkKgCiA+FkiCvddhsXJMtK
sCMUB8hSJkfk7cp2oQ4/Q9Pa0py56dFkGIgkd/SsGfow3iFkBjz0sK371VjoMPdQ
TjJN7YHPKnqUnjbtzpsyfqP2e+dUtUsvoZzoMgCMDNhlBNX/oId4rgHGndde6R/Z
6grFfjNIqOsQ5v/mBx6uoZqo2iOJj8MsDRFHz0Qn9j+ZhQyF82dtY4xftikqgQHk
T/1SBaeosvHb5ynoQRSA3Wc+ps9CWV2H6gKbKV+LN2pSauOSSPSoO62+DktFERAH
hO60StVxG3nJSDeAqR3NGfXnxoJhlrdtcx4NYMuy2qCtx5pCN172/Pz2YkkPivg2
mpqJngJCdQp9BOmtJcZrvsJv786/HkgS49DduhgEh3NWJ7l9Hn5Hh7db79rmSk5l
2k9HoorA/FUtFm3oL8LEbAAQ+wWX5wPjKVgDTUKOErd7NxlwtthTq27T3+Q/gjvy
+3MvhTh3NKaKtScNi2o7ExP4iVxzZRU+XQzlA1m2sIc6WEvtVUBrY90KjTuiHb2W
xA+JBEy4e5MJsk4Ln6OyWIt9/mR/r8gSBzkXCJhp7zqIvLpegr0lpvtbFN6dk7yo
3JHpN/Y5sKzhz76wZCVDnykxy9kqxm6iIQXPqg6uG60ryTOedZTgtieS0bYpiaGw
3faB5T1WhpOoW8K/86oJcu+xsM3d6eP7WQKx9slf7HRcYrENTYxoJwQRdx4WETaR
APBnPDnh4RIDDF+x2/kTx3iBMmg8kU1BSlCoj3hmM57Cgl6kQ77QdOGtowPoKiOA
nZrwVOf0ePmCcC4CGq8Xo3urgl7dGDrpMwz5mKUl4poLFxsLC7EWoCIg/mjsRqJI
KA/vfyeYBQp8DtfYqhhGo73v1JXiupEM8Z6w0hXZDWtKZBUepYiqcIQzADyjIyiy
3NFN0+lEtcl7MMOllyOzc+p2jd72zuq3XMxCoOKK1JfEydnYhFekmHqXDk1Sa80e
zpWu0q8h0fLpSB5xs4//VW7dtlAzgo7qbo4CzPLx9a+2N8TA1+VQym+noV5yO06V
H0LqJjg7rP+Rjxi3QWL1cCboRMAES2D4VyHG/q1jEG0oTpavQfdqQHguD88ZgLR+
0l0vpLiKeMMXWkFUnUSH7tkexxLvNCUxH0IzacfSYTYs3dKt75nfVB0f0K2t0t0e
EWIGYSsoiLyohCMX23STJSwakjqGCAfO4pJC5dKHWTTbeAuto1bidinyjy1S4bB3
BHaQ4ejLZQVpXNpg4gzVMxQx1AliBLX18ezkpGIxdsYS99KITTNyg1uilFA6g6w2
p+lJTUx1vT00ko3OzOeIoL1Qy3kJK/KFQw9EDUKBkdbRmuxO2mqjaOFlyxjn0CNG
FKAAJe2n2p3BNpNAnEL7aMIov4b7LajvDya3oFsca/jP7NZyUfgxPo5p6RjGm2UM
NYusO/A3mpYI+HxAKtenlqQwMaQrNYGiIwK4J+6w8rR4ddwXUVDDCxyHYw9C9AxN
8ZhLEyZ5PF+N3pPoiLypL2Oxq1ZM9fENyNizI0TKb1wxLr4ZbI5DbHlyeeb8w9mO
HxHC06dFoZ0S8RMz1Cmz8Qx9LwD8Vw5wG695CZd9fImZsjmCfuVvt6O6zDKeFQc+
yAvJ2AyGYzWuUlehCnAG5TCy5tKo+DzOAYaSxAJzo4ElsGvzSfrbYWW8t0OW6Pml
m2Q9Cw+8eK2P/lT55DeUBWOFKbUhAUFWLIsxUj6AsHKEdbPiTIIYBNTkr0YhlMKW
9Yy97TkkfwtRK2PMFiPKL8YebDEjHKT9/lTlHd613FZDgRCdaUxQJIrHikTlqw/K
FfWkz/RCE7Mhzb6wLgyPQgTLfjOW/fPxjnXj1yeeHHnoOcKUNPo8I7rGZ4Rj/BGe
GKvRPXS3eUuMAGPQuKNAJQ8sthzC1sWB9VcU4F70vvvTHZGSQ4QdkS5HN2nTr8BL
GudjAj2JLdpFjJagc/hTAm/u10SKjmw0mm+MBJv0FES7qel/0QJ8eFHZ00+dgSyG
asUEIaPt5T0wH1VD+RKXiePrnNpu1NaChe5CoWIMP+no88187fE5lnNZc1R6ZOSg
e9Fb4cf0Xo3J6QrDChKe4Pfe4qY78HFkb7t1+vvmUv2lFXWTBfnCwWi37NsTUGSS
d7OUYMCHUL3vAJ1bvf5RpuQh7d6USLUt9Sj/VHIP0oIplzPCiyGqv3OSmWU3biof
nNE322slOzRSA3IvRPiYZXgIpH20nEyL8cIteB2PV12nOnfSC7ZlkHQcOsp/xPQu
rUuh1IlHcmLcMpExeefgCsmLKBPlXczwLlW4770M+0xqUJ/GjE8YBCwSsmFoIuXA
LbbRHmbPB4c0fKToBBfShu9KYmDKMGlVivEbA7gnY5431DAX2fZqFInU5NdUod/U
gHdMBjs0EZQu9N2WmjgUBCTIIqtxQ9ju2rTQJeeiVGqQ/KeirO4c/zNOSwUtTJLn
vdJtE7vwAeIEAK7MMZ0XhQK9BThcnhkVkf7h02YzX39haQNr70pL5FeO+Moekipe
f+l+aBE3e6ISUXmj30V4oGvxt06KzVLyb58IPD7cW13y37FXr+ZR/AOuZfSYM4v9
sqNyvTpnDzDjqKsGpT/oPTp0Mr/UvC+iv/Bg3xPGGquA3Q5DPBHuRQ+8jbfx8ktm
bHq3quTislfLhpFLu0nZrpU6Lb0wBwkfDHjaw3vb/dtOB5jeFVlkpTNLPfQT2UqX
Jbxo7JYzVTMijL9b+BCocGg9dWt7HQAd7N1+Bkb9ipB3YNUCOI/1S1nU+CDbnJw3
a8XcsLA5ks8IGL1JHc5+rD0vygh9VmXEmLuUXVJyc6zaRRMdCxOWQWgrqH4PLGjw
oksRQjd1H6kR8pLxi4tO5WR8T7yiQAModQweac6WwqlfWCNPUTuNw7jcrvc3n0t6
cIsUofrHlm8KFMB6zVvSrQsoeYq6GVYK/CYX2sShMuEq820aOfKoGwaGWEK18Eal
ULf4mMBp5AmMp4Nv3V6vqUj95kRFmUJNcwAStRbjuC7SY0WEai5353TT5F+s4qTq
XyXZo/g1FbxoP+PzUNawo7sfz6cMGkjqnrepxs9VcvWqR3pGysB/eTkdwRZ3Nh0W
iXSIkj7B5+uwxUd9JMGyve2a4gwZzF0Q9vvKpFLPqTwLZgrtoT7MpbvahKu0lKli
oNFdjIFLi1FAltErcCPVOpkB2NjILHGJRPICdBcASd7FvM9P0Sa/Qm2OMjdy1D9q
B/Y+gmzZ+BGwSWEIUbjf0xD9gCM0H5ZnU6hyosa5vKzTG8tjNXfJ/Huuq0W/Gb1F
H0R+qaqewexeManekj7+HtI4yXb1Byf9AlG4ksDLXpmk6ah76WAqzUk3lLBEZRy0
Vp4TX+l4I+QE7IKZhPbwBj40p9GI7oYqkuy50EVBV5QOCl/VZpRs8o5Vue1k1O40
3JR5c9ZfYdtimAkNRmS5j3Jzwt/6+SHK+KZn8kSzt0AIXzAn3nGllLs17HsA2vBI
NW3PFuaiKL0Ob0+G+6m21jcHaW8M2KnUquZb3a+bgjTH/9pt7XlcGrMLqrR2HRBw
EbM24GMZI6NA4GrOznu3BQWwwQlN7/Vqj5JSajhnit1UMK0LFjffo+9UpBDjzAUR
YCb1f7AxXWJ85xXHmRjXu+U8iNOkmVUupz/BFiIw1swoxpqE2oXi7Jexll5Ri+R8
+03lyvQt/awW1CtE56sjG0AFlYfpjrvEVzCY8Qgndz+MBTh/eAabJ3VrYTJYVsZ4
Sjph/jCk30CIF5vpgmqP6rHeEZKAo8NdijRNsRmZf23Lw5CJGJbvgnjWnC9BLkjy
3FMNeTz0ZNuTdbR7IMkDZQYsZGJrFqL9scFPVsFS8MBlIsYMUiJcZc9t5lVDxU96
e8nq7DyyW+OEV0FfefdAiyKUmT14qUvhHcTyciwQVVfpnQRKwn2TGrtHkU8wayGp
Z04sjplBTo5H0kqqRHoht7vdyu+VaGEaacClyHIAwgsZ0Vodxgff5kZtItDGIXgQ
nU+5iv0KT5vnMYKybHEovkjimuv5oH0pUxwpahLD/KduD8PCFEi8fhg+w6VNc4Nd
HvoY+RxXE+ls+67LCB/AFDMkJO9BMd3hCfhTw/0YYnWyBER5DGUULoQsyDt4yJJy
54Hj+/NrUelheccqaFw+wUmGjK7axJbx//voLCOMiXvQ9M1pg/0EWTIClRMvEEP6
ErKX0l3NyxbHEG9pEUgSrgFGBafwujkEbS6B5PxT4Nt5rd90dswnMz86PK360+Mo
1RBRa25T+Gh9oKDQJptYaqtmZeMR9GB3dHcaNEAefmy47pN7hqQeHGlIoQFDETlr
pttTo+WLEnYRWh2AwK979k3JbTNXCANNv3/jGzqvW1g4w+CZ83Go+6R+wa/D/zGd
DUG7ShQtKc31ZRTYU+VMwgGQjw+I0ZBvWM6Bi08E5Cd1K9XvnvJuRAchmZ1AhDgE
tH/Wb4VLuBmDjb6U9tHQ9GmcNKyGO/CcmzDWBUcdWiyzbpBWUXt83dPusLpZMhnk
PiQAcUllNTOQtxXy+OeBkvR9ef/BiLheG1+ycM4W1iIUxu4USHXTXu/MB4AIKLyf
AtaC5Brbznvq8whrh2IgiMKGlB6Y9mdvebIuZGXcC7Cr9/LTw/OpMWkd7JK+f8wS
bYJMdLZ2OiAdPHCpz74QKHZ+zSsk9aZQHbr5z/JPyLr03kIutSkzaKRVgCtLHa1S
+QTnEUdhpFB19EbaoDmj/Lf1oUNBgW1Slv5kpc/6DFQZPr+RqjC7/HJ/MlqX8s5f
g9b6TSINlKLihy5QH3LsDzKLjQSfxlpoCyKWDBomiMe2kGxiSykkka27fbHrEdN2
hXdE5paa/ebR7+SNFKShLX9lylOBtzMFHDoTQE+ONDEgMLs/XALyRn0yg03LHskP
Uh61Q6PkapqqS+hv098nJ5Dp3XKMUV50f7XkQYVGeXf0+HKbMzViqU/kiAkTkfS4
pZIzkixE+g3leWodizUTgQYct+Np5sR8YsKCX6a3llSUmQMx8V4LR7uGoy/mAOmh
zdAxpv2p0HUDYC4e3CinQWhXxlG9DyqBYOq1gfnhUFGGPIiEMWJhrApc5urMWFh1
GPjiROoWsypnfqEPxGimtEBYOfeQj4i9fJkkae1g+2DJ6LmgKqa16NUxsYXRwVyl
/fJIxrtuO0E4dpDMDy3MSx/t5LnueI4BGoXtUQNFXs1EUGf2s06rAwXi/63zXbSB
Tmz5jrIx3HVbA5oVsC4B7tCyyytm0gY6BQquGv+g0V5HQnHRdYlp3DoHTS3MxdbB
IhkK5Eo519MCMlUIYHfyWOa+v7EjYQHYMfXR5OYQcZx8rU9Iivl61A75ZfVoYeDD
RdtLm3CblpbKx9y8vYLtJYaYhOG2nphX/oMuoQ6f2kme2oaYwoT+R/7tiDQywL3f
lEzqyThUcTgpFUyXS89w2wr1MP3/6eJcCW7WQh89sHgJaGkcdm9vOzDvY8vCD67D
/mLkHMvI55bA7yEoBunRWO4AQJZCWmmKJzxlxxZEnqDhT0suZl4GW0/oyIyXuUM1
Yffk8OdTcQstBjZbb+eSrtDGQmGKGBNU5mwf8ykn5aFDM3X1DmShR3r0ZznwXHi1
eV/0NYN0dua1zCZabHY7zjC9ehOlHX/AIijb0sYGKtK5ivoDNP3exxiu+RiKC4zf
ZWFoJwWAcLxQxjntT/v6meu0EQWWcQVS/1Sp5pqcwqSfe6OtBWrB9Le8tUg7G5zl
36BVSg5SgMSE7hVQZfwpydwS/KwbWWgFWVG1GDkwlndW1umV6qHSUosuwzZZ6uZA
ryQi/YbQyelqOAxXtRqrmsbZahb9mJAJRHyyFH+YOnJ1lLyUL2bCRkZ9khd+yvGw
sMzpQ4lEiWL03AwtLRmhiwrgMFj9wg6E6QlDAMexXwgh44tnY6C6aaTedQsBGfSC
8O0d2QJjv7irH50kpxiEb7xJAXCB+KkwuFEgXL7gLwrOpWmck+Aeq/aBFaX2j3Fn
uuACZjzxHFs25oVHj2vcz4jO07Nzz7UbpE22qY1nJIg1m2wCWcPSoK2h0P3CUvQX
2Wzo9BCXLRYdu8WnSZ8FQGD8c1ebXXK6ErUuCpk/ZWUAzgbf17V8JL48scC/ovUI
I/1Yv54lO7AneZ7v4MzB9p5PYcPy7l0vAh8kUA72Baqn2tHTBvkMSmoymqPorqRH
eLgX5jLwxuzGV5mKEpn/1FIj5HWI8YshQ0svRyR4HN0rzwifDNbs0Uq5e95Dnf/Z
1I59j5UOfq5z8EIPp44tGMawQnAAtVXNtMQEKsXEuq1CThfz5tQlQVhVRaByS6g2
wp421Eac7frUKOk4WS2D2eXv5Wz4ebAXXP7icxGcnSdYS6/HJMPU65Lq1p2h0BDT
mKAAGhrapTm6aSmtRTSPZuu5KHeA0L9aPjuj2e0UcoWz6WG+Ld9QNae2SFrxcfaY
rL+xHqiag4Xc82Puc0QOhf4ObPUPXQ6wIm0VnAjUjbYmG+Y0aZS/hSpqZfe+j0jk
nKDCA/xvrVQfSz6Js1lF01ODifZdig6PyLbcO3OXXp/cgqHgqVYjcvjVYKiXVMGE
g9WiahY7aJr5pkCbwBmgWvTyN6SUAB8/8ZCCYcXoPKXeP6/+GInrg4Pz78OLKIH5
lo3jGN9OKh+eFrnv8T1PF/7tPRwzGR6YpCbX+AH56fObU0OLH22iJy/iUY7VM42A
bt9hYTB3N6FYZTVvTz66/qSeTS5LDWO/CuePmXeCY+ubODv0CXrn1igeedHVhHoN
Fi9etI0PwY4/MJaLPqnKa4exmyh00gTbLf7qEcRgwLZZlSHZqc4zM2SC/sjwOgn9
zQe2yI16lmcmXz4n97spJvyDEzGqaOrbXSpq/QvcVT8QceBE6qtER6LRugRIEPhq
UXntLme9DWCC3DbayH+ssuBpxwaTFm4d0SQQienTl2PSSksNi1N0wWgbQzrs+wIS
nElmQdqqaxkT4VuKBB7DY0VXKkDTDB1rOZX7LOYoO2nMmy9ipe4sBgySTMmgPAqZ
Y9LVjY5iO8nx2NlPtGD5bkinRBvmDZAQtXre5cxKL9mwYmElebEIqAHGORbI7vhR
hgTa+/H4KbzyA1kCwzyjxxUAoHRKEx5YMd+S6RX64Czt8DviBMtLlG2ZuWZSx33Y
t/JQNagtWS0xFX2JIQJ8zOhVvQ/Tdl+UxXtjhrjkKG/91JTSf3DJzsS1Xh1fNUY2
92cEaeA/TliJTHwFwKM1f+ZkrBmXhS6g6BC+jOkFFR/uLhUqXTgZhKyQ1mgMHoyk
VIn96UeN5U0htt8GpWklMeqlaXKGhYmdssyvxiyVO99GYbFF96QhY1fDrPxUmttV
Uyn0zwhtXEO30xM9vtSyV/LTk30chfv6nB73YPfyKfE4GsWNpbdxwyvLcb2HcTEN
BrNpGRSZ0Gw8nhGTjPipuD3wlxp6IAYh5WHbReMsa9YF4DDceM0XbE52ZmYNz/v3
Oiv6zMZeOkBcIG6ezPWU1ShRNcwmijPhcv68eXJXZa9qD9XWThGSzLC4BiMS1URy
HgmBUZDGUtZhTzR45Nk41ESFyNeTMzJVeh1TsCcw/HzbevDQkK4QxREtmppikr1/
FAzaAP6d+jXTwcLaiy52BIUS7Hu0d/clUs1OEpTtI0NAAMvbaY2UKekFRbyEFqpb
dw8RKtnNJS8NM57y0P8VO+Xhoa06dw7nLZFuekB2SHyW1sIANIR8Y+z3yZxaegtY
JQogpLWd3wmAf7b5G1WsrFO+nm/ceXq9ftK5GBb76L141EIKbGaTt6S1DNntSyxz
JDuMjx0wJPbId4HL2l3ovpmPe4ZhH/SmlFF89+QyDEPEv0TE5X8iFky7U8FQSFkd
6Hcf0GFqGtJfOryYcbx3F7hhWxWYmErjUKCUvbuHSgs2SPx/0epyZtKkQgVbaF4t
cm3u2ZW9oI0r5yVMbtEruVBU2+VLtWnt215SFuVML5bKb69ads9K27yWOJLKca2b
LJwRm9h+GFZ8ZEobfWVe8Xu1Nku9gCEWhNuN08BV7n3SmMeJzKpyEiehlcjS/+dY
ms/HroBpmMLoIDqA7cvm3skgbHCskzRnWz9Fe+xr5LoNQzZIYq/sS1zvGNQX08eg
LJhdLpdHmiO2dLdBF0PoC8tjG7FF8W2NkIh5x+3n86h9rM1Af99JU0DxNZl2UlTt
i+njC6VqtGTUJdldq5EW7HlQxJoe89hjUz6F/wSP7nFC6B4TE3CPqs7XFn8E+Y9b
CNLAdFzko+Qx+7Y8X59WTLW+otaOwAJ8corAemY9K5JbM1X6Pb6h4BXNMg01D9gt
Au2xEDoTxWgKVlLE2dkyjoQ5TUMQDcexyHIzZ/dqA6TcXE09D165z+WnTmzeXJlW
Kxe+joUgoDtuNgadhFBo4rgn78sowcws92oqjt0qSBFj5kmM+4Q8hhmye28L/EHn
hvl0vtv62PKSIRaoi8v5pNFucafnLf8Q7Z/e+TaW+Bmfo8U/Ng+kY0SPoFNoWrMg
B4f0mFK9BK/5HEYoAsZsVZqrDOBu8bsQz4nMUr5CtPGeO3ftTRDeGfYSIpm8eC7v
MxSdYHLnyyST+wd7Ua8t4dvnkVnzGR3ksZMDUSXMSTka/7O8Cerx2aNKQxrk8ID9
Y4M4Nb51Ha96Ukla+J97GAR9/OKPzoDAkc/5ra2jr1t+mMA3aI3gUUZvKHjLL9/E
Ex0u7gESL9gVQQcklzyOi/V95xTBLaPdC/90PmWlEyxYod5xYke4PaCpzqhnoSo/
X6G7sf57Q4ryDiDC9q53M8qzpNelW4gUJxfNUMx2HjBhlIjKmCIE+UN3vEI/a+xl
ZC8RDP4eO2yv9y49AymDzMhcx1eCaiE/FAIDSpchKswYecsv2y/VNjLUsOWJNSmu
XW5gBSbFka1CkJqEBpiez/vP5xI8AvDVDr7CFHnNozCIbheA/zFksAQ8GZA4Sn4E
D1EGC9SDVAyLz7ZiEEeRYfNETIPBbog72tyfDg6B3dTrCZYCXBa6H5pY6eeDfZlT
ec8lbUmdizSx22c7McmlJlroKrehtaKJQj+wMP0ScDh4Nt/UCtgYwEiX2qXCoY53
HeboxzpLFNvau2XLbTCe6AAIqBru4FDKq3IFR50/Ln1cLrIFqalmr2lWjXs0QwRD
XinFfRPNSKndrhBgPzYrsPo5UE1qbmySgcqnBYojBJfAF6cPiRocla+qu+EqyJvt
oiIU6fs+sZyPwl8KJC1C2Z+q5cgkdzulT3L9w5iUMjFyQixLV+BEjo3o8QixauZZ
nSALwtsTIOj7HqWwHfDDGpzKee/oOQ7i4wbG5zA5SuHovUqsqXuvysKu//YBMd+J
SNM/grZr/+a8UcSZdqJHV4VSPvl9KMOWgZ+8NDLe5nPwIjcY2BWy9gE/ercrIIU+
nTPxijMc+falIGUfDdvdNMzlxfqGRGYM1GSZRVKvykZV8JIgXt1p45+d2LB625ZA
24OSX3cBAHV4hDI63HeVZO+GFs5cljx4+YkqDY/P64RVACSCmXsAv+uoZ9ftd0jM
iI8T30hgE2w5KjqNHgwrpoaBALFQKRKYoxqnAfNroD41EIa6vpK7caqHmtgxpiPl
s3G/9LWMWYu70q4lK3HbPrG1yTHP0d/NhI+hKEw4+MluuhRDAPJez8CLXKjdECNU
2xXsrIOKo//uh8FwoOhWtIF5osWA62ngkfjeHZKPWdZMjdr+aZ9V7FVjNrAWB1h1
m2Sfrrdbq6L96zSzLxbtqV6nrJT7aYR2HRnA+aeCB5SgkvAybXffIksR3DJclY78
zt28MziWnPEKjKQjODMbTXcDYgocH8lyGQ+Qf5/sMYYR93lO6jJIEk3cDtkH6T4L
SmOBTqe5GJXSGWTX3CXykW8O/t/Gts8xdT4W7qm+4QQQCGjSSyZP88UiOAjSNWhy
VFYcPH/LNMHRw0UbFrMJf9IOb+y+SY1jWU1rB01A/HYHqz/1ReuPwNKpLlf82+YK
+g0e+AG71fGsVpTJ4TwzUF+m7SU49LRhgSE/FxJuCkucHdX3phkJagr8pEQmqkNb
A2r1QNWnjzcO7LC5G8M/SebWmIBGn+zObCRQdZYFo1ProVP7hYDbgmNOoxOvdw0X
b3HqZOnGO7Q9V0CAFanAq8io5ZbDgWIBf/gh6LEQxoMcE4n1HKctl46mhzSUlNpk
I/5ffIo4EHvKhJkH1pjVhCuMse8ap8krqv8KRTHu3zREuoief52HvNs9JZJRX5Li
8GxL6ffH9JElORzdooxBgqbsrYDPnn/1ZEAqWwraWZ4HSqnEzEaFzM7/QIo9/+3G
wcJ4BBEJ9NwGyugN543JIdnwoZNYD64dAeO9o0BMmioLPapbr7qzqrOsKkDwl7WW
AbFB1uCW7vUolMovv3mLMC8SQ3CusNHZZcuEOZMYN23oZmq9EG0G1gmCqendLius
hBTtbsZXQ55rCwMmgNpVLLEAMjaKyNvOuBVUFWWRR13whceiFlIBjP5YCvcXHOml
egvNGBwFvxO3SWpSG1FvGT8b1Iukq0d8XLHdlk/Yd1rnZY/OElsBoDnWuxBhRU52
hyPmS2tXUW4MkTJmWQv3vN+gIdjyqNaEtABN1Umw/aRxVH4SH08smN5YH1m1yN7Z
JntfloVXmfYbtn6FzSFE7zM48ovC3K8gFPucdyfvm3+qTGuW/MtBpdWa00vygdGT
eeujGI4eRgJuboGNwbtcC3jhn+wVcqI917czB7qLRh7V/ZpdrSXWFMTOVDAtYJlN
eGaV5uctY1CGLZbaq6HlxBjHixWh6k3jKMqJ8I92mc+v4jBvir/bDXaim5Y4336O
4zBJpndSrDWL8/hSuZIVbMMCK4ZFK+lYez8faRTSsDr/pv3FENi0rHsn8AWXDzGq
QaxXSUtxg9ZAt4+f9iQXi7pN5i+vk7wVUL9aMf77V8/zrEx9LIwOxESAp+vb5fPw
bz3tC5X0x/2Ct0jW6hBA0QY+1/kw2cgMogvkH8NTg7I0VGKbZfpeH6uyBgsoGss4
6F9Krn8/JiTibqCW12QmWFWEfHrYlCazAPkxwR69JYQk//pNJqPx9eJ+KZlWBbg0
UE4Lm9oKkw6fMluR9VYfTv50Y7gGbxbgz+5QUgstzou4UOhFZeEAIiPZCbuUZfl4
Tbd1Im/m9stjK7YjZKxOF/NvJri7n1QhTnaA556+3ytDsgF6g7YZM8YUjGwp1B39
lSlXVcJrB8gaeAp7xwNv7Zpwd0+f3DudixCMYpqQKhJviTY3MMxxqoP6r8FLbFCT
HsdNoThC5ihvOO2KgKNvzrC4lLh+8ylUJsI1mhothQ1Tku7KLKoKENVCPlYNpmot
Zo5Pry5OYiqcSwdb15Z9hN4FAhh6whlfAy663s0cUPY=
`pragma protect end_protected
