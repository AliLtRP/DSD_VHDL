// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h1TKUHG/i0ZHDM+2plgtA+nsDrYpKqFL/Lro0fZrQ3QfOMCUOA951QQM9YQ92QdX
53A/4Temmfho94r23U+4VS5kPPK4gj6LvJZ7nsYJa48T9ApPIsHIpE4ezGiiZ765
XchOn9YeW/3IUYZVM/XOAL0U+mONLYrInFwEecH+5JE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7424)
Zk6BuiNK8H4H7uvSKCu8Mi74COz1SfNTu3hcd1FftzLaQBxrCeGWLKHfPktRJcBn
zOspjKoQZ3q3J3uKbY/RbQJdT0BJUHikkK79q9txlkFtMmp2Gsjc8sCFFAT5HV6j
i/7QZuFz2MxQK1b+h4w79Kd7dcgpM+m7WKStIOtLsHcMJkeSfWnOHSRVgSKBfRiL
47gvtSVbzRrbfqjTmQkBUJZ+G+YIMsgm9SmyH/lNMLRZzag4MLbBYu9JGPwqcXqt
fMK4mvUAr8k7dfKwm8X6ZDzooE78cn0IdYbeUDo5d/XfmeQhCSLMzmIJDUgbSGfw
MqMK8JcJbHllwNK3qflvATKWsUufmqCONG1Alic8fm+EYFRKx4Rhk/OgFq9Qhe60
RSaQ04bNvb22M1PBxuEddyS8fjHQ2KkNkOJ/xajLrrj9duJ+zVpgI+Lgpu/LSeQp
pmCKZdfvspFDEqvEZBrAd/OIyGsPdfb19scyEHTIlRSdL/T5wgYzV8paPzei84P+
bdknGaOOyWdlVrPiL9QdmzM3nIk95PbKA9QQoskiNo1JnowYbpNqwe3QYY3dkklg
0VpVYNn5RG+fjhcEZWWd+2eT9IphOyL0ssTZwbtCF0PNAvudVQ2UBu/JePVX/bWB
9PaQH4+eQJRxs7/QqkPOJOAo71XnFpWSW4D/PCHLhhY2lsfZs8rgRA0n3USHGxVL
uFSGVZjb8zDYSJH1kua4QVc8w5luEWX9UL1cylQa8xipyRFu5jvltaV8HdBo0u9/
20PkXPqQ/8kNuKjre0SuleFI5YR5ma3qRqsfA0yx8+0ibpT100OC0IXvyU7yDYL7
H8p2RWhhXLHqiCSx0WlLcsrtOgpXczQuJDdWl0nr6WX4AqZLQqlr9Rae5ntNIsw2
b+spqFdUsE2mPoSkl2p8yIB+tW9rpmZUwIDK2V/h8IJzVTi5LUkTBfvvqc1aESQw
a0MBGuNMmbPw/1Rc/9DQmHSMHPXpp5ScYGpojupksg47J/PLmjSUxBCSXr9xSUYN
O3GJlywabesW/WvnnR00uAN2TZw0lkrPVaRdT10mkbMV0efmtHDAiX2cmBiI4kAA
RrP3d5YUqGkAaRP6lOh80Our+udQ3cy5UO4AIDzHYcK1Nb9rweeTMSNJqGPwx+xe
K1IeuceoQfttAyJkDLoiCWiuJ9QyLSbzM59dCTHP2PBStPfpomjf7KX51PclMknf
5cnOFQpT5CvR21/oRjnqTR8hPwtXoHoSOFU4QwANW9rt035oOpPpFU19A9Byvwiz
9mFyWkaqbdIhSH0H0olSJO/ctGFkshEYzBGq3CugeMr5u8PjH8DGQcNDzZy8vD52
LHS7e75ESntOV8nw1GKl5J260TGjGqthTkK7IScPrHL7omwp+/haTOsX1sswLjDb
U0yOVtVidJz+G3P6WYmIQ2paFFnghbq0goV1gsCEu8gxhOeMlWvCHUItoMWhOEdd
BamwTWoPJ6lp1Y0SAxn5PTU0klP8VrcwcsV5XOfYWodGwmFUJRzaBRxuSFb6dMi4
u2jcwxnxxNftFEqOf0wXdUb/hT+vC4Knm7buTF+ZoihtKJBywcLcxkYoCTWCadQ3
2W0cmyWGPCr4cN+NNqywPuzNJQSEdBve8ugYjfOl6iywAIHDSmXIUY5zVf5VPfLP
QvjO8JCjrM1qP1+2TKYo7pI7lqFaLZMGUTNXm1B4lZZSwAxNhoJsKgYYJi2/Kcwe
DyU525pVb0c+AK4Y3xTCimG85OFkq8DfBZb+fDOQ2QfApqln9cIn99k4+ugPIOlS
RmnA/mE0jsTP9uJyMcHM1l2W3SZtNHSHZvbGMEBjL3uKN+TQHvAToxkZdyCngVpg
KsYscU3KAIQldZY92UpAw9gDrQZ8Ud5PKZ9W99tKas93mWvqS4JFvn7KMO8ReIjy
43hBlyBsUifuoCwWNQlCERAjyxVfkC3WfCRAQByMJwKg1grWsmKUQCZ2ii4VbM48
q201ir6PNoTGJia4yGkRXV1a6YJPwhf73rRqY6UEEOS4nG7Iwju7igIXe0u+U2vx
GNxxV7Oa2TXpXM4cU3dMf5/RfWdYvcRdFu4jSX/XVaUa3nYfuIe5BhWwXqekk5zm
ryg42FHRp2Kpe+W0FwOaoaC6sCvNjOciaIMeDiVuaiJ4R/71RAgBcUr3rv1pCnyu
5tj43j49noNemoEz3cK6FQgIpdrqQuOxnNesgQw/eDPScZyHJoY3MVP4aEosha8T
mIhho57RrcEmY0HiOTjP+LeAL9UlqdO2bUNSqd6qDwirAqO8bWmy+4KFGhSOXNN5
vE+nRw7dGkKmUpVaJeij8+6FGmmL7NPAPC4OfJO0t3iLPfJrtEhL4T+WkVWY/VjK
KRmEmf68ePKK7t5fKPIDbzRmJ7g9gsU0ynvXVaNFTGAyFd28VdJFgziOdp4Ng3q3
U/5tNwcCha63D9Tq19h4GWgPGoEhytfzJqhSLUAANyKr9iAfQ9RFl2FsQucn6cRo
1bM8c9fqPknQ0EwUCVfS8SV3B6T+VRB2dFGP/ZVdobDdx36IKX2xPpQV/F1+wGZq
AFVS7d69vDfrz2Q6viZpjuFSqjFhI2ypMbCfGKvu76DT23RTFPCwwr4iV9ZGUbUx
0345L6q2jdoAWb5BDahYTjg8EbzLfkUi9fYGmaJvYVy2D5qOZszmEUkDJPP98QJ2
kyH22l+vXavXc6jmRGNZSlbvuBBuyJX2xXrzoeDOBrMW26pCcEx2MVPiBx1SrpQt
wrIdz7L8GdseFQWmzsMA/tdOX41bLdK36HcXdI4lQ3aUY3rCoThd5xGq3ZOPcDyU
OYoZinpt2ev+uFchfL3STflYrNUxpbRr4PRplxxdrTbnk45mkxoTxGi/2R+ZpQOP
cc4JTz5n6c5qfGHEaBhp5aw2F7PAFDTyVTs5D5XSpN3YuF5++SUyJ+0FyWEKhNEx
dVAGgn0R8hsIglw0ToBEWTwKv6P75Y00HHJbTGizg+H2F6TEKt5y01IzfbCDQjvx
Ro6ubxFz4OA/fvSalD/tGukswjZ5dNUNoDHSzquvUVMDuRv2bnDQSGpDnI4jZQy4
WQsPyP+7iKrdf960I8V5VoCH5cSk3fu8qqchckWt++a4cM2rWKk0+ygeN0db+2uI
tcGfaMawOYH6tlbdTyz4KPwdZMbjBgBtSBajmh4GSTkELyMzOd32646By6MN/qFA
D08S+Wc+FYvVBkQH6Q0y+q2D1KsPl67/oQ9fhKEbZz04IQ8I3mWB+8ksXkX1AJKa
pDg0tOz5AtV8QvSJ3lmaqERLHbHDcgNBLSPe0ai7Cw9kfoSrPSnbIYx8AOXm8I0z
GGfgdGOYPqfYJaF126WzRV4pGEVXzW8hw+yspdaA0S0SFHj8/uS07qfTbyLFXQaP
ssB926sZIwB+iUA7otUSAuoqMSYEwzxCMX7MwUocYeVgqtSJ/tw5QsFKNDI/uY2U
5/jiMLLQEcwi9XmXiXNeowZHsigkL1sb5eHU4jRH8GhuUhJp/RFjgcS9sflF6/Fp
PjFP4AzN3iXNv3L3JnbNFR/Sc+vCaDnrHhj4kjR7HZbxURvQdtrCuv1H9OXUPKem
H/7J+cOuFiWvL7oz008opKQLAHj4d7CPRrS2qBx7imtNjMfkc0cVNavcgrPpbkBx
zwN8RuunsJ43Zhm3ixJcTbe8rhnudq4huqN3PCucae9lt5+B1J1dcQjXKhbPiGMl
NISaVQ35w/xgxss05hM18R+GcLz0E/xvX3Vjl0EEz/VFOAtjG9GdzseJPDJqarCy
P7BOeJUC0HEHmrhh77+bqF1T0ADTF3NX/WqGip/tpE2Y6QE0Io1jzAZm1LmtoHZv
NLXrOqXqqGgm7JLTpa0ZTzm2f9tS5pmbohK/wYmw4PAqwSq7082f9+TG+l2St7Ih
qLLJDK5aNzum8xFT0u+o+e7hvSI4zQyfJo3Q+RGO8jkd+7uClQRNEdhbfaxIqdoC
6xtKiOP+2dxH1ENT91kKNjGURVXHpjmavJsJPw4cHxhIelBN56c25qL7JKkGGuMf
+9/Y/pvk4j/VUAhif6lLLnZoq2aMF0h2bNnGX06wfHsh29M+lWYH61+QjToxX+JA
GNhDr0Ncyojy3HLAai6OV2b6V8iP0QJ0EuYkLZQyJRfIyzH/CzS2mBKh0hutj9T3
Rg9CVILVrwZCVLNSvk764HFltWM4HCbzkS/xfQ16CbjC3mGt3LmcJ58O1iRiDbk/
YcVBvgfeGMNlVi2ARm3epUsUYiJxn4pOd3MI474T1nR3NdRlgQ7sDFFZzdhu455J
HjUKa2JpYGMqkj7PsBdh0nBpP9k3OYDs7FZ3DoD4uHJvRl3N45MTGQAQHTouOujC
GtLFJlIPgT7WlNvPZeB/DBBtApr47RNAzq4AxyNaeu6VPjwUUTRHKqEGQcAXLB3k
HRbqg8o7OTecuq9sUCCOxh6iSR/UvgkALbqbwHI9C9KSVUgIbdrTpSQRvF5Eq0C9
rT+GtF/xXXzIb4kOBxfLvVDNzP8hOuJW0diwWGmwrHqc53CwcieL1y00pkXXhsaq
nQqwCV0Ar2eQKrYqe6gOuBpCYG8llygSyPnX7WNsARnZYCylElR+2gcAZB+jtb9j
Crw+Stq7vvgCanoA4RNkAcxlm5CM6jBhz/jgtrSpggDquUXtdtB0CiW9L+hxUWJK
I/CHHm1olfY8J4J+MJUFzXypXqZc/s9C6lPsSRWn3LunByuIzKG/U2u3GYUGWW17
uBR5PBVJOcnVmmaZI88rqnT99S9N9AHm2/gyqg95JgBGQ2L4rzuL6o0Jl6qVs1zV
Dkg+qHnggxVfBcc3ve0Jt7/VHiQF8AaEwmfWRu8efD11HjIaoesO0Zy460cNgSM0
3XUjSt+Uhnc5roWvKfD+ZlN0es/hvA7qJfl99fOUNe3luuLPwPzDQdmdNbFwMZLz
w33t6QdIGAvTiVkFpF0dnJC45nrQOg+eQd2TCxtkxRtTt/QvAOSKtOewMHZujDXW
RowqhIW7mS5hOciEptY8mLI3nc98sz9j71SK1d8b5wfE7KBj9YGUytRZBkkGQZhF
4nu32vEgno34huo+o1Qj9CLPuhjJZzWSoOtgHtpXw27RDubSf02Ch+eMxnEVJ3pI
RZ+2LPw3XBSIF9UGa9Kzefz57pFQdFEBvZnvTAghFGM5MTvEPQXI46ZAP7EdxwGc
SctSLgXeuAhu8IPfzWKsOc7V7BqzLCAyE0LgaE9JjsJBYO60bLr8ujXLrXCIWXp+
GU+RMpjHjlTj3snk275Up36jw8jvlJlh2FzaMQ6A1leKOt/IXt+y8w7qE5oBGlaO
oudY65nBWgViq0nzvEoRl5BylA0PNqOtbQUCdCqPHnB+aB2qTXtHgeB+0lMvtRmG
EfJC0TN3zRrZ5PVi1oHSS2o6ds4VTZ8j3nxXo/D81Kk39atdkqMeeRruSuPONt9P
zQysoPLWnpwjUjaTyawlWbHkBnsvhwE7+tk8KuBqNaItAv2Uc4tm2joUp1gsz7Sz
xvs0HSsXIFAgFcqusUdWotlEE7vLVEc4eQsA4PxoXXWOQnjRrfq6sldFAHoO2T9U
9voRs4BnoCYn4VNr+YKuDUpeiTexTO6Rlb584axEsz/fIpzDsH/SXMwkCPMTObwT
hNTzclyg5uFmKBQsDRMFnSQIiJGN2Need+vTzg1CKNYRfCL3IidBumfrmL3xA7FG
v+CryIRD/wTxP0dK6RyyhNRDLWd3OugKJlzm+q0w3HYJfbt5Dsgy1HbWV7fxgUTc
s4PfPwOW0TbenStPBdPe15hqzOm2fBj/B5im5peZlThl1mcR0eE2+DjGz+eucol8
za0E9mf7iGFQEOQApaPm0L3ZKHug+g580lm9XgD9dNLvAAtHW2vdxvYuaUJry0b7
/7IyLZAw6lUyyyjSOCKDNePkpXBSzBpCfuppwYf6Sd3h0Z2B27WXTHNC//JNppXE
A6bMzeN2kPswLGum3xuCbsnDeEK3NpfOXrpv9A6Iafz/ThH6/ClbzYWDb9Pfr+yA
Myzz6gmCCstvGPqBqxgncT7NSXcA0Y0oy5RmYOTWM1mUFQdMWnttvYpakuDlCp7Z
6ThNTZBq3W4DSnnfHthi4j7mU0baNfSNgsMy+SFcMfU/qm21nwtfoGsNBGnNI5xU
fAWgLSVhtIwIYnZsYhTwX3ILP+usqR6gsyzxFX3VG2IWdjjJO8UDONgagfOSeypS
iOhqySq5E4wyKJE/CY14RZA1O/pQjGiXVkjK9i6Kp30S/xDULsN51wo5Q9PylpPD
87pktfdKgli/rd0J4kBzbLft6i/dUMW8VjDPBfRP087kZR0yWRNp104Czz4Ik4hD
j29QWUzCocWX79oigiflA06VXnzrk/SmbCkWdNzVOUhhLzsOaD9lu+gHaA0iZL6E
cAON0WTKJgFjIyc8N8ziMr6tM8KtbEY/Re225yO7zsTIR+Yo0arprrX5kngmdIck
jDsUITbR60zn9NH7z1uC62PW3kf9gh75nwexQ8RfdolnWpAkwA1CnDHRVOlEeomD
dVa+FonanNyidQ3kMrZeW7zppx7wDyNIIhHdWKxXsplzximepk1Xh0LW1z9bt8yC
731Yzdaw3aucpXIyO2bACz8n0fa9ZhalMRupkNQD5bkzaETlnsgwV+p1dCtViD0B
rSPu2MuNRwvwyN8uDDnJfG/C10/zFfIJ96l+Xx0GNIjfP7i3T+SzXUbnAF5rVgsK
mnpRhI5SJ37jSDJr3+bKr8te4kMfumSwA92FDpGbGIy4MyRYjBIU8gENpY0HAqW3
mRgsKZkJlYFNhRH3jqOEFOOpj1V/hQPPS9nl4vLsyjJnbQGVs9vxlPk1loneSJGM
Eg72q4vrYXIbTA8OYXPUl/qdc09qAkKxCol7QxUQPt0Cb4TDATCrr3yf2E1Bq+1t
pU/UgZZ3Wq7Lx/TQSagIM6VOMGM5pivhtzuWoB6c+RS/Kou4BJHPnQAG//QolHWy
NRwGycF0aa04UNMLytyAjrZxuv36ns1MbTBvBSgy6oxF9qY8UDYJfHwIyEb9zxZ2
s3Y+7jQc4cbHn/q6Sziy6iW/kjDwdIER12orDd1lyDDKNQLcL6FmVeIe/VcgDNQX
gTME3h+8Pbmaf5Vie+8N1KY+7O9SD6S0LDz6QY1aBR7NSB6cNi0eA4WtbzRQygFl
gMDybtXDVWSxhbbNMVdtwx0cK67eEM/ZV0IcARs/O+TtoP2vX134Y2Q/IccJdslK
vkaGKiLY4qGW2S+aiVeULraNgp6hqSqP6daOQWF1hNrgsYIrfgGX4g3+vHSuGYQs
hdIzFJWishOssaKjG/uFv20iDMHG8LN4pw0m+tHrHMvkBFjMP/Qvzagfeo6f5j65
O37K+ZdfJ2iC5MFStDRlYQSzlG7FFKLs1sANXmnq4mcZGjAX33vpl1+GEHGd8CyI
WEEpAtmh85JrAh8rsDicJbztgku3PjhHL838DrSH333E7c1uAuIuOyL6gCkw+5HZ
7U7PVUDBu0bPCBn1AZX+YVyyAweMibkOzfZoAJCMkket1FbS9Uj7hNwON29WwqrJ
NSsEkI94aAhQaK6syVqawnLa/z3miA1otaC28KKkYWpUwveEBX/lprhp5WaMKzgb
MLXZfIl2d7vLOyBgU0G3aLEAhUU8DDLtcd6ncLzWZgQXtIeM47l9TGYGSkhnGYVL
Ikxbx0Fyt0GkIeExIpDizHJRdal/iohvtHveQ5kbf8n0N1arhq6xCcbmiJxGQbzt
xx5kCKv5vEJkAgnvE8umlrzAV3SeS/QfqJ/6HtezwWx7Q2eNC8RZ/tvSbbhsVt/b
WA/g8RZPSwSFdw2MTTrtvK5ebx4Er+I0cp8dUlCT9B48VqO5VG+qk0OMWkeGnA1V
H4bw0iarxx9cFSVxq+UqXqUaXCDO3qljZGKZ5Pn8xhcZBh2U8F1QkVDPtyMHxHtD
NcMBFt56xZvqYfoFHJLKEA69julLMzzfvNBaIR4SUt05EfOK/EMfXaSptFx1dbNk
O3S+RhTAAoJp7WF0NOe+EQJoqOEgPt7UQK5wDdI+ko9Q1XugtSFTa0dVnNs8enur
voWj5TFfo/oBAiHGQpbVOcBjHauqByfWE+ibEnOyr0DZHF5IiG8Cc+4birH2g+Pc
T49F5SiwPOqHu8qCJN65dgTfml4qty8LwQrQXVhVNc6ysfTnkUghctMG+rZ/KfHo
LxGNRkBYB968n2ESFlszSq+bQhq8BXTRxa3cQ76EeWA9hPOg1gOQeaNrTan9nAiI
W/QWgV4suze7ZAd5qBdRaRmoAf5EHjk7t4jdcn793mWByJQWOT6JUK+cZlE16ZcQ
DGuziJ7hCeGfJM9lWYBDx5tUJ+n3T3gGMCqANRiX2j1gujVTCHW5Qfb3svESRaGl
b49dDu2T7qxAnGuCZMttgs3FimNkPwdoRM/SpiEYakWOkEn7+KqyvXwDo5ZDgtSx
YdGtHmbK+H54N31WTTUYrcBYRFtXo+2wwfbZdwOM8l6He4Zk9TGXESGqEvR5r/p1
48rOvno5cL0+noNp+C8ja4Ae5Aq4hn4A4WTunyoAgAG3omKKDefkh3TBopBQ5sUy
Oyy6DsRNmgAgl0msHZYzbZBP6YRgJBliMsRw10EE4pV/Ca7vF6Wf2UMg3ex99q7M
na/ltHn7k1s0Yx80hLQ5AW7HrI34BbvksYp5E4XC/PSkCzVNn+wuji/K4DwJHoV9
QgTiVG0QWyr2uX0wYhi6lXKQ//ahgVf19PBTlGW7nLv0LFmOc7RldiS/6KMpTjco
KLs1WiuF19bQhgMc1nCzTbGzTKX5l+JFyikSuHhLi3TL55TNI3V2zaYWCwuK0QkP
sQEjmH1NbpgxRYyZxKH5jhtfvJGe84uxaziJV+q1e6lBtuPVUV3qG2afrmEMoMVt
YR89oPrmAucrpvH09PZyk9H3oV36T1dNntwyCLfAvT7au6baFP/rngzjQ5FdC4D9
lDManOejh4DqTIVY89PWd5IPXYbGGFX4intlrv/lgblEjpAq+q4xijpsw7LrpRCu
WxPvap0wOMU8uXSxhu9qxuPhjDpDXG3XfgrdIDRY+eW1pme3gMN0MVLVl6pOay3u
If2WMPFW8coenj8Dze8NiyNt9LoKVVB1/OF8KDjtRgJ0QDbhg0rK3I6UvJjF6lWh
YSslI8Jhb5MKPQqZ860yeRZ9d0EsFyQRmjKNm2+F1/YHM8l2NGNauN8rwTqRbj4V
4OM/OZny8w9SzvUhxx1+OM5+ZUbRiw2lZ8NWviZMr2Ic6GZdWd6F1mPAPKDBQ2F4
2jQRv8JS9s5PD1tZld/CJ68I02t6mFvXEjRHAusZGD//cgw411iAin3EfFR57AfX
qrAwIO7v2bQHljiEecvH2cczKOGnVevkcZRo0iXpP4HM6LWt25QCmKrFM72N6TEN
eNjvUeNTYDwK1La4W4pCfVkH1jH+JbCrncIkLZPg0ZRFiUtoHqex8eN7eAhNfGQl
xP/rlhN3vqMQ32JIIJDtjk7aEmm5jJxEb4zm0M8GmvitV7MRyxboXdAEQatwVZ/G
TRB/Xw/gAShsurLuYgZeAqe1wd4xXmzzlL8rVzOKobI4/JcvkN+gc8GYYkK5qPgO
nlGjez1GOhBOUHqvPFXVLdVZk2RS2pcsR59ViZJqzmaS/GO/mUTt/XWPXkQFjd2n
bE1E5dfJ3QQh35ZP7PbtCbaHtCU4ZIiVhkubWdOLMpSC8kBMRQWEPOzVRLyOL1qS
Zt2fhUv8VaxgY8+rGH9Hy5fcX4KtGzNq+zvv056Y9ZEaybQOORS45Khinz79BL3r
OJbVhJXO2CZV3MjHJ5RmXTJl6zxCV0sBZ751i/zKW8s8HvVRCPq7uKE7St4poGWV
vUJc0y7wQE6D5I4IMWbdkSD0HGZqTYdpkkbb6vcE6wA=
`pragma protect end_protected
