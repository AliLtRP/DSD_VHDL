// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kHbcZZ86dNOmNM/Os8j4sjDE3b8YXorMLgAicG+KEy+86Uz+YWifaqESmBgytY4j
ahSyN/MLV8ZrLYGjcbEeUGXxw+9T7l52T9k+OuL0AvU7rbOPacKu9RL5PyN2fP0j
JhMJAcaXy3iunLhe4ngzEb6ToVRjMn4MyoEcbsOZ6qY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25152)
TPZqzrAo9TeFplQTPiEDyMLXHwihGnfPXGI9f2xUwYHU0yqfYql3LcCskdoNIHFi
Lf0+gt7Fcvp7MwvkMjzO/7C6KG20DsdlUwfZNxfmy4t0F+niPGOzwmPAskEHzEBx
qKttHMr7zdhzXqPZO9DtrtVEj1S5d/MbRt25JVceYzlRA2/mnSkvd1FvjbH0eRfB
ftT9bf3XuLfBRSChsZpsJiotH2FG6f75XxLe5pNk02IjFeuj3MMWo9H51hkkw4Sd
A36djzQKy5EXMTI6k9IBII5AZ1VISStM2funIfVr88P67Vq2zIkbWWJPTf2o9xtd
hHiAPoa1drINoDzvkhnJhmk36LeRlBe2/al/Jr6V0e2hGZaUzVVQCBJnCJs9AdIh
JbbIb3qmOHXacseWuaRMPPtYvctENvbptvWpwzkGB5Kg35fjF66vfZ+Get6EMRQ8
o2EUUyh/yuLZSv43Rm/dXWNDovUXNnbPhNzvFULHX/NTeK6iXgsE1QY+csmickdM
52GdMvdPaSeD77qFuKX+dL/u5o0ucXXbqdXd2Fgk2KgCfk4Epr7S1LIfcnADKvWm
dMQpEwFHvIbBjmaG+b6nDkNKVLh35MmaRtnL3dX+u4rReauV4/IZmpiN7RrVmPfS
VCLF1biVOwMWCzfAF8WlcnuG+QpmPlMvDjAd/CAfGzljn4fRkBsS7kb6GPo1TQd4
Prm+yaC6WgZsyj12IpMJkxy0rjW62oxqrkZ/OK551j/wgXzi4KAk0A45358W7fR5
QuOEmANongMePQq8tGlVNlZD6gVtcCC6sNqEx2XkwJdJ8BPNOgF/9sfbljOnAx/e
4cR3HXLItBkjtrdqLFU4DWhxUMFqwDk7OpSbbZWuBy5TnRTC9E+AAEhmu+Mppgjh
SeFjOsufFRcxzwUqQk7hQCaANQi/0dBA+ZUS1aafMxY7rUcENJV3ROkzuZe8fSXC
AQgSwqJ+S+Vy3Skljz5I4Ehb3rCFYlOvqo26L72DYzf+zAIe+l28L6aXUUWCBKEF
RhVx8tpd8hkJz56MqE4whUdiMPqKbKaKYX94ojaodJ4G+T49aKsBfjMm4WIRPchw
BAcJKKvwAIFdSdwqIJsIvVuj3TSiaxUK4Q9DZt8vZTVanU1VuThClnPJub6yENDh
16EVoogr1NnJLDxfcrsz0onf4G2RO+1EbvoyqWFuZ/SNbMoPhyWdi/H/u+StvRaz
Tdn5RueT+A6OtFr0DdufrPse5ToPSU68n5lW+BYiWKvJHof+e/HVocDP/PvMi3Kn
99PkGOcblpTStHY9VtDf18oE0NwkSrqTgrKBEl2m1th4Beg9irZ2infPZCXfyvog
fZD6H5mOH44HuMoiOpnODlYg+a+qS/DGqjrHtsg5LOCLZeKSgnMUtxuIwQVV813w
fzDdjKaQRxB9Z6ZG2iziCpBXSWvOZtEmX5k2g/8+5bR/A0crYd1/gQjNuArFbJfZ
VYXYcSq72Gz7ux4rH+R1MQNO555XXg9+/0jI0687L+SzjNtURs2nYaTJ9Z+YIVpR
4bDeFjfSwuSEv3VNbJrpR+ASEY5umEUL2y6HfG91JkcvPSuabsN1bEOy/rLwfXYf
s0OQcIbtt6wyQMSzT3/AA5k1YXCoiraujb4Jn25/F3B657dB3hVUAceBRCVBKaiU
/fzxyAIBP58XpmQ2jMxAyJ4YCK8WeZxfxQIWIkb+GArcrRIc7N2q91vTsILau+Ek
OMHe5r3J+Xewhsj2iFy7RqsezGk7sGP+GqG0pf93wo1SUV/0jfuaaPUOufBGw9a+
YBL4jrvlsUBFZK/n11J5XG9bC7K86C//LfiuRoA99tfUFEpEp5bZfUIDnj2jSLYe
0aSTcDuddV0hGpSBa3sRAK3Z1nrfw0QmW3AzpgqFXvDMEWPN00p7+PDot/kdPl1i
YQt7whd+VJqpyNw6NVW4G+d5oDRKqE3ce45+tn4YKY5IYxVBbd4FL771A3+LwLNG
Ctpm7+2MJS4+Qfpk1sSfz/cp7ShFSMsh3J2bRd9uX3qWHZhnajJ8viadb004qaQR
O+TJP4ezvGaMHyKZjo+QI+6kPU3rIe3YfOPhk1Fkan7Y7q4GdUrytv8mt91FZgOq
be7r54zOcQhP6qa0rw187Ywhj8k+VfEoi3OJwZM7RvBsJJSquoK4b52r1aB7v8Q6
cVgRBNcpHwFHZl79wnnuH2064DdX5vTk0vREED4AlKZ8h+apOyFqY+kXq4pOeu5l
STLRd/LFCQIebBOb7fqWLWXPp/RgaPhEMSGRPujewXsIuCnjeH9VQj6LFS1eqGfq
9zXqfq4uTbOARwWT7SmYivpz4XK7EO0QVSKZ6ykcbedKz3p+l0PHM0tXLCaqos5G
OV9WXwah+Vn8bFG0TPxKPJU6mTwn2Y/32uJUEbNFYlzWQhLiem8Nk7hMniCvPh/f
oWZIgrlokyiZGyjw6yKdhnk629nxackFrV5GA3Aw1S2UxuZf9iDPcZNrWZD12QZs
+dfg/cx2rFW8IE5tXmnokV1D8pIxMIaZNAvoxcpGkkvVmeGhMj6Qw2XLT62tMlju
wYF5w1QPlskpH8Hgk4delJrTrpGYhuh7yWB+Yjr3dgc8pIhdSh4Q/WEMyzY1+4vv
wgPPP/ptBGbLmRMxBDwLJxmxTwoXVudUyRCDpGfUBsBCy6NN9CLLbvOI1ObpHG6c
xyuwOkksN5MwrZYsfLqfvC5BHquDlRcWOD3f6cvWuugvFw9duzpqc0psWA7SGpzR
8slkodEy0Q8VOoJTEiv925lXH9GTG+CaobRV/ZdhG38DXcVJJUbBQ1IrrfEBD7Ga
plGRIJ6ABwxnIYxrqfW1f7tf8ABHjb/qBOoKJOoRSSJ2RZhO5hGMeccpJSwT8Fqs
NGmJyAjcVFeNpdOWIukdpq1OUFgmkpRV91n0ILW4p0Gofk8l6GOzivetHdsgUyfL
NbZsrpMWmow0Rhg1nyFhS7W2yBY3WceWpTyTVxpw0jadjbSQ/SsRG9XbyMhhXNDH
lpSlc5aV5x/FKMZnhFg4IxpE6+lg3K3u4EOW0FOaUhOMrKqSMfnQcv26EpKY7GwO
tczpBcqzgz8FAliGBNz/sEDxw1b+xAl6iSvD5Vbk33z7Sb8g3aIomBxX0ijgXEV5
DB8vWx2sY5doHUkUO5Ksw0qkJpYuGTlEt9F1gAgXkKKNl8+jHPx4ORlPRRsubxyQ
9bfSUdintrqhy1JXc/PMSvYS4iMLbXSF51y3gnPeydkzoGuW6kDQg+4NC0138MMw
/V0W+Nk/+gFESJQUmcQThuzKr9D9Kv88MX64Ft7UUsI4+gU1KPwowkFOyTCCHlge
ASWHtl6werLE59Ic6oTchjd08FPH6vr28f9wap0gcc6CN7Sj7LvHosAb7RI8ykam
ik4BUQPfL+OtmXAepZfObGKcnVG1QmfPhTG52fjHLmHBUW3062KO7bQ3PJBeKDDa
fZkhZps2FdbRaYIIzk8B5vrG5hbu1BeTIkzOOLpI1he6clzLrJquMjyELiPjaxEk
y1pq/KSASAEjGADCWJtAP/Q6DZgSujHdDZdjIrVfmolvfyzHeuemhfYGdFBvj79M
a9MA70sBjTHG+nuslNA1zSOhTB2/UoJ+jQ3niK5IV7v916fMkutm3qLoB9x6KA6s
bTzh4bfTEnJf/Cx0PUbJmmMVkmhcirezqebWpJyuVexKyil53Hs0OZKlCwsgKokT
7So8fnFpczRF2L82n4s7GBNkzVN7gnxdxCTFV2IYYdYPTynO48Ve0TZJhYT/v5C1
P3qRK9ArBDPlhVCx6FdpIVg1MvuKoYt39F9kW91bCVW2a28T5bLW/z31X3PKqauB
7abJPd1L0dKehuRj6SdG5HBmos9wf1mUUtjyJCxKbcFfR1hX2MCpvFgdPciYKYmx
zqG5sFc8axGejNB8Lrp5tsKz7Zffd4RMEw9sEhbmZ9BMjmWZs10ZMELy2SNqGpNs
syvJxyhr3T4qS4B/awYZ/m41fjHYpQ0zLE8cIUEKilemyazrXj7Gbu6M1W1eEICN
hDEg7gizlQs5DSboeJFl47iUmJtfigynAFJ01iYK00K2z6Z/32fJMSOKgNsg17qI
+UWoSfC/5yBvwD508G5B2ocCs+9oqYHm9ZxOPX7nLoAqorJURFIWLmqj6PfRcWQf
1ZQCXIRe38exue/UQq5rzOfwg3UAxgEQDKEPesKaNKIssw6J8/4dRYofSiRNG2bo
AiBxXtekHUmUyrBVtDnI/gCWjX9JD2fp8yMIwfHU07bXsWXupXRRsUCgVTLLEC/R
u+138Vmu8k7W4owZXt6SM8+LE+vsgRtn2S/wr09ZmoonZNAgKTZA8Ju3+UjcvIVk
TUlma5ijjWyf4kQ//hGIL/8ZbJGzot0OmqrLDc3bZNTsoAoXqz1ePvplRL56IWE8
gam51HH/ExkmV8DnV3qLyZyEkbCEfna7O9x3bfjlR6Nj1SZ56y8mWUSiEsJM9Mz3
TmHu0CggkMc4D5jZHgrDzqTxUrzujN31/iTZaqCqXlvku+spmmHzXZJFZxbvoG2N
S/di9NwiH3BYi0Y0wnND2iu9wMF9EtfEC/l/Ccx2+6NZu3kKYANydovyX+08WqfC
qkmgqCPRI2wcYXz282fc3dV3p7c3KWulIAx/ijrWdf0GqZT2fWXzzo/2Ip5pOXrz
eizseLZix7MI/a/hXgcPG2CkhmT3eO1++yVH/CnoirfwgD/QPVehKmO9kbMyrSGG
fpLA85DW3WqtaTuRiEYajkTZgHSQlKd2i8gd5MnbMOCWPqdcggeOw1g1S/vst85l
mhPowo280JIeCddpvPkYfBas4g27qKm/BaakX4M9iGPBZJqkfCMfceid8DyiW1yN
25RoqRG+GqPnd4fbpp3bqQyz/ioeOCFBKdWuZoiRP8aaGjSyEhghMtSxQBDbmLMR
UMZy/hyJdG4AgLxaSULoHldLhhozJdlJfMDl3TS+qHOP6xsTCZWxXLX1efesGTbj
NTqUJI/H9XorqTJ1ANHTN/DCWpmAn4LH/EPlDljxH5nc9+Y5iwpxjqOJMOxSjg2u
CjS1KKsNM+6C3/xd31NzFjfcAV/EAz3xB6AKYlw5oJE+r5J0j4PhYReXTbIU7bh9
4opFcbq39iXs9FQoNBkc6pLBcu3fb694iXmPvqxsnPzm4VtUMnfNQ+EiCVAn9e+m
q24QH320FhTUA2RWeIukYKZzoIZH3/K+D03lbDClVS7eff2XRKB2SYRL1YNu1bHn
86cheIjeoIC12H9H2QsD5+TjEyXajUBEFDzmtfoRKqXwQEM4EFzPTOJmyM13mmaU
dKXPSjnu8To7YxYdy7o95SRlrNLzYWnaKEZm90unRTV+XTJOFBkSm4gfsEr6rA/Q
ztUjp3JZoMb5RiHBoO5AUuokHdLrjNnvi0WwcMfmooAI5HMeYb7X2owYAE4lwgkc
yjbRKaDy1eGrgqr+Y1CC5gqaMsTGQ0Nkye1LHXW/olnF5YMLIVY+F3gRPM+dlAPc
lE/uL9E5n+g8pRbAOGdD424rDM0uPGqiX9xtrOc7RXRwaKTfxhqrv9tSTALY3Zxp
ZHHlrx8+oVYgJoEkV7iyMGrNEK1X1Q86D0ePJCTavpVCNyBJk+LrNnLXZrola+ww
q8v6i2uD7gABb9/9arrYnPN7GvpuClFvf5zy18KuW4EENmZ5UKxswQnCbr4SGZg3
lM3hfJGt1p8UUnwlUSDvqyQQnW+jMkUyIbXMuzBBL7rSFQuFcM96YccT1yuuTGRm
AmH0cw8/mIqCs+bdm8CoOExL87+liQ8AvIeRQ0nip221P5KJKkAe7koRE/2K9xjc
p1/R27Xsdxg/5e+yisgz3u7OeN8pQigYboOOQ83SCrxyNiGW7ASfhulJz5iRo8g4
4IsemHs+ld9KtOKmL4TLSjOMYjWFncvPJHTYejq94DvtGHqw8z9UPif8eVFGMZxn
N8Nj3E1cKMDvildZuxpHBUlLM1csb9SUlOWdBqYhjP/1zxYxdO85JlkUrkPAAD4L
HQe1Xz3OSOxvLHXePSLH8/IJpPZuU/T2ur14Zy8Jwr9dLU652UZvCw28k8IK8KXZ
QHmIbCoBxoqqgdX0fIFGJPwkseUt42tju3lqXZ13PhFU2/s0V1/hetiVIHTEg/Q1
MzNLxPkr/GC31eBrwutVrYLEmM2CZD2xq2SD1r41O0TWM8KK3Ud4OMUREYVaMSFw
ONLfP457Oi1A567quDhlk2KplO1m2NzjRpmRLxYhAAr7iAybBD4yGt0aOGaOFOAC
bAvvKkq464rt6gfgOl7rnCVP76P/u+CJLfSRtYlOG/KhISYgCll4mKFwUXvWEP9n
Av28vqcZe8+WVV7zO2XLnslnQk1cYQrjc/x5jxqop749ZJaIoy9Oe1uxAMxAkBox
TyFIAexM+goi7I1pPxa0RsY6Oj00ntcVYSjPX274844YpUlKSnnpktwdPlvK002p
JDXUeYr3VLMlMDxtznDLgQj5NxbNqOCgnfYYjey+DXI24w4Q4liQIImR9lcvoxMH
MvSvfzwGSkvP3qG8NDlUHrcb5zanGCtTzOWTU7nV9JiunToZ7cGXqkcT1ERcvCbs
N6CKbbpBouyr87V98aZ/CB6sbpfIJry0dIZ4wlNc/5jSYjlKUCLARJSSgKDvMAd4
+Gh9YalDuBX5jdOBkyQSHKOByTmytDpwrX5ifYZ6IhViFGCJ0cHLtSHruDrWbJWY
3KUAGzkYZ/Kyfu3RqExpm0l/W2O79f/pMbDOANQy/gJAqZOikT0eCa+xg/JBtCXQ
zsAqcQaGDfYmRCmd3fwMIdxIMirQ7SdI4+UZIjfj5yO1O+EvdHjrInbn7PP84v1R
GQTOf9R6BK/+Ibmu4Z0dJjgCFXMRHC6L2jTjmVIY5vHJm6IQa66/xDbASjDD1l41
99HipbI7EqxRICRZ1N6f/9oGTtqxBag+aVhI2mKPl9OEcNugV4ZzWls89hmM8rEY
YNCCff8v4faVt287wwOWD4uMvYNSQQLA2drE4heQkitoa8fcX2nZIqJ8ruc5wzjq
iwj3iEKUoqGcIx2TBnIxYlzjfy2G/gWrPS8TnhmTEjlEiGfoTgCxJXWBi5GGCHVE
r1ZJSe7Id2mFx6iotm9yjE0KY3CJ8mz6VP3Z+Z5K7Tqtm/cSu2dfRMHXM0P3aY7Z
bUzW2t5VsB3khs/V0qhWHqN6KCw1JtHWtXRipA1TnUO6A8rIy8+GwfYQsaB16wx+
vh6R6HQKXVLif1TspHLDwOBmcggrnRoqpWgONXKD3FTnxZr7TEycRiU6RgTx49Hv
2idX0+EO8xz6x/l+ciWwP2FIQHXVHf4paWt6IP6mq9V20MeG3C81ZctrbUgXEwRQ
D0WFDGLGUJQ0jUiNVMoflsCsmC7cTbMk17f00dnsZ2Gfke8hsi/uw1Aw/Q+g2Yrv
oTZtO47sekDitaxVbWH1EA5P+zf7J/Gl5pN9iPsWJ8x3iAMc0i+4H9OI9r9wd+Qb
RGVEpCKRHKUa3kmSC53Xfr8QFCvz5sdmuBMkss0CkhH9lWArQxWvMVOWjevWr4m1
+b8bMIOiiGUXX2nt6LSWcVVLABu08jV/DfvPgS/9/p7bLfYK/XU768TM0ccehbX0
FYFYT2UJvveY8TlW1fdR6w2+bvdzSimwxg4k0yLQoMAQ8UF525vFhw0uVvP8qbA3
Z7R0jv06ArRJym5ipxfz5ONkaqv462nm0rrVuQ5A72OTXQ24exMcA4TiZ36Kyxu8
zwHyeFMxVXeDWvqnmZ0UvDjgu+r1916+EW1+VQa2CRDNTp7EtL3tBDA6Z0xH1ZEa
OF9Nn8J3wsFEjDp1wixxRMvj7VvbgxHp4uRcubJR8s++fElhouOKFx6hdgvxjBm5
AwKNE6iMVII6PFl85gpZDCJ/znoyacRujdcYT1NL679D5xEd12pRn+cFQVqZkZ4F
lQ8ninDb4jsutzvhSjV65fWxhxqnh1JzBjuboxPAqdtUEYAknMtU2kb0Hf6kiKft
SflZsv6PzA5iw2J7jGWAIoJTeE5OR0OO43U6OkPLFPMzXgLkA2Vc4Sr/5s2r2fvO
XYJVOpmI8gIt+ccC5x6YqgmQw2CAqZ62ON/i33ks0BSa1gwtT74EPOUQThtUu0wv
v0PKnJnpYD80EO7sGlfaI8xBN35liDYveZDnysc6Y+MtyP7FhYEH8hyjaZPcaKIR
LpdZm3WHaweoMHfvNIPeVoTxwIMMGT7+xFKpTmFm84xEvI7+LJUFSrHTrRD15Lle
rKlYQMkqng/B/jYXVVDJqDF8qq2jxGBFFy0v+xSkffJ3n4zPBs5vcwTLNcDlS35J
G4/NOSuaauW0+dj9dpby07oPVIjKzFIGlyVC015DXzw8qG7fADiHrVUi2afWfPPK
dzgbb2Za+jRuOJFg2KNXsqaIfmlcb2fmUwppUvwEVM165Cchf5KdzQQNG9rbvlQX
sIL5F0LHttKodfC8T1y7KCQPtFlsltasny/TLiuFkDtlfO0UXgqnVqT8oLphuuzD
9yOHKf1w9QFMTyvYSsj6E980thS2ECsNwjg2nbRVmzd8TAo+J+rFEcq4SZAtgkyL
f2MaxqvQwHGj88/PhNON888FpaPCSmmoBC/34/bMedGrIlo4Js2zjoZe8atLnKXn
fOAy23s5rbBTZUWNiwnOePDOXDoyCLnNGfgyBBwCJQZCigm3sXZEBQPvkDDQVWAd
aC8SjjZhKcVgV8QEIv2KyfJl3//Jig8wi39Da/gyhRSP9soj8x1/Lx6dsgwYtRXP
zM8r10jeb0S5LOaWEj2NZGQLiL2fJeLdi4PBliFJQwZi9T1McZO6VM51v6L4iZVu
wz+561b/WsqLCQDt4k2Kpx//0AV9Sk2nG+mUXLFi9rntTbxppw+cweEfPPxhPaGD
IcYwygv/tSu6jm7FQRunzemOsSPDKgS6wWmeWSLXErd8jLfthZneZGDC25cl0YWu
8Jl0mjB3a20skkLkjQOlUys+u31KU8tnUgSVJCAdZ5EHIk7933/bOswuxltZ9UiV
I2INTRqHFXfSCOSH6pDO1gEsRduJu68gXf/bDOtGRbK2IXsXLqZZwNoD4TV1DCIn
0ELeHbCjE2rw6lWZMgHeqB3bIY4rxHcJdsMrqMbxhbOvLTlhZkRQTV84H2v6izTK
2XWxvTRj9Cb5WulPbbOafNLgR4MnuRJEiSdz8YPXHfaHMrOpJEOlzyIoKyWysq0E
Wv8vhvGY30qyr928r4BjxP0vdJdXVW41x3aeyS/gjmY3IKkVDdlUolSa2ZbX81Ao
ci0+Rk505AEarCasKacFHIdTUviKuTvJ1bwLIFqEGoJZqDnweZietTulOAp+4HN7
87MDRpm/xSMqGQ1NTk3y/yl0EAhXgJFVHPPWRQ7kg4P/W4gkWbJMtmkFm9fofJzA
Am3A3op8pKvyOSQRBvWNEjKUI72xFoPfHqMFSKS0wzuSjA5kA4x3qbqgDdL/aQdk
IQ8yilE4dOsy32BzydGkw7/e6w903KQs4zPf1Sjt3CcjXS3uQURqYE+DR/QydKYw
0Q85n0kKeFn/AAeYpGkZXWqNddPOLyQAop/kJvPgvgQpaADBE0XOvx7LUqviC9oO
ZofEF2+eu4Zr+5xWAT83U2y8Yty54GKkA00K0AziWDPIg8rE1tJYwo5b9mwwPw+q
LK8n8er8ZZnaoZEHyTtB+ua+GaBJxX2BlgWwwSxBcAo1shu0wz6orQsftaAnFxTA
LQjKwCZYMsInEbQOQ3pfqlfLzoNUwou19GNRxKqrQYdSHAPbdQjhmvaM+2KljfMS
B80o3EZ/in8+SmTt1yaHxvpy5l1FeP4jZ5EdtfkvifM2b4UhrFq2aFBCzpDwe6r7
g0e3W00Swxu8gd6Souvh3nq7qc2ysRuqIjvZq+f22m4zvM729t050C6NiWwuZdpZ
GdJam0430HltAFocgGL+Z6QiallBJS9U9Xxk30JSTK75aH/aWQU8/YS+UYMuV0ge
Wv/a9QBO76UIFDVif3Jl0kl16uVc/FkSwhcHzRvDrX/mddA2QY583tYNY6gDWdFi
w7YySF79ybtmmck54mH5EpSo9GY66vK5SkoOVf9lLf8SdYVPGvpCCYINncfNUHNL
S1jdvdH9W9nahkTIfX5ve/tQmf+x71Q+0Ntk7wdsVqvjk8u7zOEF15AcM7Tc04Ac
NCgfrfD4p6R3CGTQVXkkay7kuMvVzFtldis35h8frNCeWpNdRQDsb3H0KQtrmphk
kaK8p9fwED2VvqlY9ZaN+kl9JNaXbWgZWdtwvr27CvZrk4DpIpSzd+kLn2Qg5ymD
8k1KWTqx4XfVZfGyW25QqSQMET8M0/oPSZIYzW2p9ZPs3I0t/BSAuosc8CHKxRQF
/Tl1ALPkO/hV/VGC9t1Ey/Q5t88id1Y9THFehdr4NekSJDvhSIXlu6NpjH8zC7Tm
/9p+lTS2P/BKwoLYnQ2uz5uDFWmAR/ESpP8+LQyTTY/gukxLYjUN3PAeP0suTAah
7huHhTkSyBei5ueOrGKc9l4NpmMWyZ1uDmUjqQ+wpkaAz6QpneaNKHx29dv1KVUO
zJpv5vwNuCbRSH156HtFqHkbvZace7geOcRAilTQ0j7Jo/fj+9hvCja0chBqjn5H
RpaWl3zH62NYb6ZdZDIH63Isc/kWbE5cSIwvrRVfakQDjugNdR3OftAkVROwzDaL
WlCSxFl+szwwplImlvoLQLvIk45SfwVVfWlr9Dxv57F9OHZgJODEUbX+aJyIKPYN
sZvKg70z6WAmAofcEX+bdvglregPfcGHNGLjLDozFpE4UyzcuG4jJnxLrKC8K71J
EEUmiDhwNDRGmfrcauZ/RyI6FW/5q/fredPVaDJvgYmHZNaawjQQEHbK81iRqrz+
Adqqq/gIiyBBnYYkO4u6Z0m4ZTdTX6ucBByDKXHzOfDLsjGNdYtqbzDYn8sHsHd/
i8CeMrDS+lPO+SU0eWlWzmM+DqfPmSJeMuQ8cXatc5QoVtC3avUmqRmnG6ZjPrgq
IxUQj7qszbqL71xG2FNaVYaC35zre1F/25oHglr/Vm0zPXDTuvku1U9+oDijJCQp
qBaqFe3EGae5Sl6kRr0WZcwy8IfgyjJR9M1d/i6SQob2K6yOI2rnoyhgStSzpxt7
S/xHTe3qZdBb4E7ktrNPM3a3gu6a/oEvlPVw5YjBTY1ILdJi+dYEOSgEXR1ySw7V
HxY4MFSUcCTbf/4YStjog9K/tP3O0P3z4ab2LXBftjBq4rBN5bVKftCSItA+8wzh
CAgA3f7yjUdaubCNP/zsqjuDxheT+0i6BEo3EmYk0bziQ2YPBDsE33546MoQwYAe
N/6lhOTwjKA/ryjVKy7Ftkm/SWfmAfkGrzX7hKmHgIEoz84iR6+A50h34w/Nuj5E
GQjrQJlUZIK6xuPm8AYSQc+iZNi9bu+TlwRTAFs/VdULyhdjolOPb82S3sttVuPV
hDYxqnP07UR9t3apU59mGnLCOtiDk2UiKjfDGCTbsdY6DSpMAMhQdMJKt6NeSv70
s8dN8LyDeB0VT3gCQVWq8xKhfv361fnTgTJs2fvljZxClA5wewNjbDaRLgeylDON
oiQozeOM/s8+9CwuRVH9fcWKrtju5CqCN7vorSerV+bQxwJGoSm5RPr/fc0yRPH+
/GRI3l4flfKVLCkBgTx6mEv0XcbE5uu+I8VqqUFXwIHWZwC7hVQM6ifLxhZhMnfh
wp97hrKi6wZePh2B8z426Zuw4twUtUK7qYWqlRn01SFpBAF0R2LCJJrOaKeFw9u5
UQsLP0bejfkUkdvfmpOLuU2Ey8l2ZDDDpch6b7v7ahT6CEfqK3fiNeqVvSXpJytn
T2wMahf0mkFBbalzu+GgvafxWILtKpXdNLYMYTPOgtAs21WWL6ZaSNo1ehtVm+bZ
2gOJK5ctrk1hpZ7p7Ers4zAIuPLfyATMfvgFD+Y9UaNz6Nn0WBM3m4YDLxJdGIB/
bEAZTdDDj3M4h+CdNmdKBRfkWcTPL+4vT2KasSza30H4WAHbR0koA+GJluwwMGFO
VSQF/Hdc/fxsrnibpr+az0kXHbrZbXJys+ANDvAbPUAXpOsBmtcSMEcE/rEu+3wK
mvrXotympXmtgCHLD5syf2FfAV8Khj1jB3dtna5I3d1ONi/laswhKEdzJC3O/L3F
A/AWDRpKm9dRsp4E8u9EFxjAa/2wqCF5RQL97cs/qGy8LGOCu+XLXGeOXp1tuBFt
kwWHx6hGQa+d50DDwvfxnRcG5nJaDquAU8C0DA4dunN8Nk32bIhHYuIarB9pnd+I
UqwNg3NupD+IpQqMDZdcLa7aREuKwBnBbm7ZAbDraYSwa/N/f5b6jEWtEg1pOkLc
41+IKlhPJzxYGclthUTwxUXMZKbMsSU70Vk4srV7GHkOu6FQ2KdDXlGMMaINXuJ+
/VhH14oc7sD9CZj06toM/yCui0RKFkz+iHp/yX133psM9KVhZ0M2ODXpaJuWqQFg
2nywzblnoHn9DB3RUFIvBYl2lT1dQg9NIeNzl6Icr8ih6K59j+ri1ca3d/pBCv8r
0PWRiicsKpcEGFZG5wCBJIUPhJfLZZEYC1VWEGP6xvxGd0/XhlG90Cx/AR//KZEy
YlI1qfb5AIN2K7STy78IgIj7Wbjjk+2Yetfp/EMbeF0IkbTTnvX11IFz/EVHBatf
mk8NRvl4RKJ0k4ARIeKXfso0LuTHi03v9GaW/kYudBDXO9UfLPPgJ1OJE4e1KHCO
WI/yXgcNuABZuukZn89ppUj9wYs3/HWDn1Bc8+WiTiLEy29PAvi4226NkmP1xku7
H7nFwus4gao0ZHUoRFNS7jzOC0CgIjg0Q8Y3pyCKAxvg5ZBC/V6KbgXIyi1ZAaN7
jL2k8CYYy1s4FJBL3s1Gthkp5/OYCD/T2JXuRUelIaN/et5wj/hmmf3NwwOF2fvx
NjfCI7eQLkVz/RDRsskVvET+zZJvHdiWHewfnVJtN9R8Me+uMwV+IeJurthXyXYI
bvQOjpzGgOARFoVWPfjSiG6ztWkmVFYp77onNVVHaibnjS+iqHdpFbAkdeH6rF1T
6tu63oEbQ1yVMF4jzmyrQaGkERzh5mLK0A0YIgSvwzRKxtjT7pjjJ9w6ZxIFeSZ2
k73YzVWb8lGcZs6FDLoBBvjt9i/rMGin69IcA5dWZP6Z8hS9gWxb3R6vg+oxYZ7I
alap7TCKol2JXQymDpXoM0XhabDmPfjSM5rytChnuxZhuBLlKrArFvfBp7+bOVQV
uenXzispPDIyI4nc2PCQ95D0evWAdCfmtQnYKK2+V+nYp+GIoi4CaXo8/3FHn6Js
9aaGIEStLLqks8/kmhnIn34XRkCdiyROjtHr8j+Zt4rm58uezIEhbwpu3He3vyme
w3L9/eMHDALD6ANUzDUrfAnULWI2gsDF9/ujLSz+t8qDdm1RfO3Xes42oCjApQ15
VrjcKwg/GfJdtvofErfXBy9NENEiUdhJhjqH/k73Pyg5lTV/Ddh58PJZC2z8NZbF
ACSZ1T1g6Uhfb/qbveGaZsLuaK4Ql46+jfaFwiFFNjlAuJa55HCeUW2ROzhPT2l4
FdyqJqTkngykIiAmMxKKekL+Q8KW7mqRPw9LtCNvcf/TqHB6Xi0fXFdXavB2TCJq
RE95MKV/3uQRPvfUn/gsO5lpqfE3mtmV466x4hQqJA7qn4jUOM1rAbLwI5h9fCwM
n5Cukc4tV76eur2BH2geto9FNZNvUXP/Lrc2iIkxmBT34mdhhWMe4mWfAj2ttu89
bIUz7hS5M0I2z3G8v8zQ6MwUPzHrssa0X9OCOj3dDKLX3sSvYoJaXxw15KUqwCJV
ZSpnSw0j7Vq3Z5WMCh4Rwnv+cMd6VMnuwq3QZ+g7oxcbB0V174CNbjrRTszQBed/
dDMx5U7uDf4fyWh/DD5Ik5TUD+gt3Z7rZE59jEUgcpGQQwfH25NaRReYK0ypsw2J
liqv1FIlLE/0/QzFRH0UlVo5YjihegYFY3VKwU8JI7t5xRvGRNeOMrpb1U2p/+Rs
d91vGsgIlZUe0TDzbneCNPc0vKWz8RLYqmk82OYhM5dA+8Q/Hoz79a09dM8QflGb
jjRbZAw6Cnef0lVJL3lF/c5yKoZCf1c8pXqftVneQDT6dkWQgqZ+ubgiT9PC2www
S6UWscBwLsouMqqATcErqg9AHjIY2TKhq883zQUKeof640JExaKRP7kAbUQS7kEg
RoTq9yOxGMM9kWF3gAmDhJK8RddtFXZ07sqGpGWKUXfeagVfXWBl9zy7d0OEj+0d
v985Ay0SPz0O4JsnXDG6bUApkSMiC+v30I3xWBsNPA+b8Hip3sm++j14xe50QHE9
WGtLQ35KAvj5fK0ZYaB8ENI5AZcgwz0G/doZNTPpKsRIWe/LG9gyUK/IGE8A0+S/
UrfQTIInID6g/rTFRMZkk9a89n2WjTNl2GPYdnnm2Gz3LgWzqg+0vpcyyBMVjmwE
0Y6Edx0HMBQuF5oUXquCrm+OlhAHmX0Lcj7CL45VE28n/vhAiD4blnKFztpEc6ZL
VIzH/9Nto39A3m77LNFMVcMYRHzE3s0auYQZH+8y2cY6WgtbGvPxSs40UzL1ADOc
C8tj0IrRVMf14Mj7/wXI7/ifzlBK66cnsAe6NIWF+0MHNnZh1R2eiGZBjqxsXBsK
xL1vAA3Kf14OD/OKMj4M1Y5roIt4GFmIKmWLQ5xow28TXEwPtzOYBJO1aRVYwgrU
cObfFlqpjuuU5cv+KIfhYhkT8yVc/c7jhJ2qbHWHN+h39iNcIHDfoHiGlt8uHUuf
nJsbglnKzjmrbemXi7ep0Oz1CJz6CyqlkgX+yIihDOBTEkdloErJzMp549vYZKCZ
n4DDEkUwDvqtJ+51/4Skn3a7AjA1MkXVUS8xbNoe2SfxLJr9dUodQD3HRJ7oX/uV
kK0KJs0+FtNlpCN0nIiYKyACzOt2BL50ERN4o/S5AtvERXbJ7gOVLmYNlgCHst0g
2a3X7AASDR7UmUl9Kfz+sGKpJXwEwoB/hBQTLT6MpPy5A9n+FVSG0K+hZfU72Rd9
1uEcrmR5IXMjuKQlwAq4NQnlibPWcvGvp5RM1r0nHrWCkYD1muCJefTPzSIHrfka
iaVtHF2oauU2VmBw3oZfu9M7j6/hr/sIzaYVPJPtep8s/8z8QvOLGWYwg5GV5O7a
YcSAJknVW8hEAv4OJpBKVfGx8CURZLkEKVMxRPLkuH7yO0kQ7SVvhmBTwjb+OZXm
PJHLNeyK8z0MHNwacO62fq+N5Iy8vMZ/D4gwct7TczYrEnJotyYxS7Q6TrEWjF4H
0TvtQsIslcErf943IJXPg47f9um2ms/hLZjCKEvedxyyDlO59ydsWtoWhCdCyyNv
UaaFQap/WSnrxjoI5syez4jeKvW8YGXbw77KF3U1O2bnRtdNCZPJewal6d1919vS
O+mQhZVe2SD8m9VaTLr/trCh8MJVt7RlUeN2ktOXiECmN7sEsTIb9RLqhoynBOSR
7RoS8xR+gwK/dQTSZosqyeeRcHnB3zHsJPpByI8ODqcXOu/Xz2/aDX7r5oGHdc3Y
SaxbOZas+uG9JJ+NpCcx5tnRsirdBokvgrTUG8jeSHzB4wriWwoe8f4PodTTZVH2
mPjY7kJeX9OoY5Oph58YNBcS+C6hdwYVs0cQZ5xGf/2jS7zV+mH8FWvsQYjejvMf
LV4vmpPdf/gR5s66ab7ydRz5N5Y/T9lkOMxxO4jHqTfEgYYWAMuGnqXYbtzT6dbO
fnK85BwRoQKjeiQAOJ6uLyVEvIPVuje90DIB159ehkmAr5SXGnc0tl8b8ivId/14
fsPbU4+UafAwRyjORE1zCOowucLHYMJILJrpUJRBckMLe6niINPOTOdABKTzjlnW
WlEtW0/5PiYgnXliQDhc3djt+Rr4NIMGDj/iquv7vQ8LZedodBIHmSfLM6OFq2Zh
CUSJjtPiX7swFhMtwJZ6cJv52TNGgmGjO38k3nTEehrJ/n9zyvg2xluSifDn/eYo
ztlSyAGVXX8FHFwo9pvEujRwIk8cGuBuujtstM0Bf7MIxTMWGmkuARuIwEikWFKU
Mo0sCLie91bGntYUWcJGy8xbyJ5VTlYi4nw8LCpi08lsWQLfSCODNALc4XZK7a6N
dbW02lPOdRQNA4XSioq9jEUNawy70iCLw0EmhXOrr+O9xSMaxzGYg8UGaAB0Kiaz
nwnn7Dj3FBlC19qFKSm3OcTlvomdosKXq71V345rDu+Yt1DL0zDfivvpufRF0pZV
I5jLdNij030toq1NC4fZIGdjP93JmIX7NPGbrrqql6vYEsYnLSAAs2+DAJubCOif
kvLkxT+MPFpZy5gXqSy6w/Ws6se/AhD/iR+8UmsDJiKTVpfPTIC0MomsdQS2C+mQ
yuFxUv2JHQ1c0DyU+ryK9WoH1/jMTY7v3hQ49USADDl7uhjk8IK9bzijSbjni7oJ
PgCWLA7YWKRWJVte1Bh9GTV8QAcdhOvfI7bydxINp3cl6CZ/NjtU3JCTR9TaGNf/
EYdua0+Oz/b6Mv3KajsmtitygLItQJP/7Wx8uzGBcE0ONb3MqBACjeg/3ZQsJUB5
uqimKoqMpZB0J6+GB/e5WXlaBwQ4+/CwYh5nMG56IN0JqZ1crtZmqXKiAJjv//Yv
ZXEF+x/swjACm6O2UvgZkNEZyIDvCBuZBhQbLou0zz8yjKF1Ha9iAv+5c6D5kz8i
/6q5w/EdXq1tumifBbTihjMWYoV7G9V7zfYo5XEhArc3whQ9zGcvTz/Y0QVmKfzA
6092qEgBPE/bH7me7ei5LiHGsZQsbJncidy/DCkUIZzzVSHi7FiJC/QELeVCYLe1
31cnQpGY+s2O0LC6j4CVvs+HFHa7JUAfOze68NFDkUCKmDKmHJG9ZDy3RJ78UxCb
DF6h6qOF/K1MgG5sz3ZpPzLGyIBJ4b3jf5+KlAVV+dtpuFowqMzKoTt0fNefPYkJ
cREHZSZg7l79oTXa0ueA8sKKBTFE5CkJg3c5Pxw1qsI2L2RR6491KTQF6l1jqol6
629PX+PmPR3ezUqkkpQNjuDl+Q13vxkRUHIH1g3TKamW3diISeBVmpR+8lyJOzqu
f9EwAL+2STU4ZAfPrUKxNA/sJG5oKRwxcjpBvaz7xXG3wwssBl4nDppdNP3Un4du
gAdPg29dMKcHmodnyLRzaF5cK8afWVuBiBibys8UILeCM8++n3XwlCfXtxWb/Fnj
HpbPIR55r8gd7xYGn3MUJYo8xyRIlqGmNcoA5Q/2zqMkmERdlI+VDvzrBhc3LGYA
SQVydJKX54bHJeHHFlda7+SycPji4QUt8B2jmb1u793vYuKuri11czmsKoKzdsQQ
NqqDLjNOkxkuWzR3+fdPXAC4f21Im6l805C1yVppr+z2zsCs40VUGyks4hzcMuws
7OyFTfTQ2tERtvoHk+CsHRB4BcfabLR+WX+EoxzhjXp91qUtGYI/2MA3udFVe+88
W4TSXYaWU/SFlDESppjkJlPB9ARKteiyn8AciFgavMTRT++3pwje6+Dw1bPl8k7Z
dFBpYzzESp1V9oIbQDi+veDJmGoFgOHBlhiChYtyh6IgkgcyhRnossQRuKfoJM+t
fRf2gj3h9OHGKqhN3QDQqBhY5Ufiwid2DEcqTLg1ZsFm5pRH1B95NiZHIBsLOt8R
u3yv/PAQ2A9KHa/oGEBcmvvGkDIZU7CeQvCUU6kG7RGWtUWcb7Nt1ETiavofF3HV
hdE5O+SnPYN6hj57cFryqsIQzwirUnk7R1oQMjQKMMbunk013Wj5cZrILTJUtrKm
9374nYq/iQbbSRL9v81RsaO/VPKGtxSqA0qAGzkHJ8zmp4E5uhR7srnHhIyZ7jPb
WWEmjdMz0to7gOamG1C7NKuIMZlyWcdbQawIqqkW7Hi4x4zjwh/VueM9BGMfiu0a
WbyG/7i7d12ZiwMBnvEG215PTs6OO+H6Rk70K4Qc/wFqBA2cJdKvzcE01WthZvK/
JaDEqWGfbddGhXGjOMr5/8E9kQOS9nS3Eu9t/Vkh/iQ0E3M+lklcuSvLD3ziUDVy
7PTvJTit9iEal75XQKKSfm3exzbIWXDDOupsI8v8aSLl5h/Zi9FrmSCYY1kG/Pvw
fehqo7zEDTMzLoi51B/zgALPloQqAlnc3VSFWIyw0UfbsOp0L0OE8Wn3REsNeJJw
T8CrB382voaiTSoqlp/8r4pWyUnLfjwTWpTcc78uugW/8/CkAT6i9OBeFfjKohUC
gFhW92aHFNyeFmUov1dcbj5ciXjTibqtuAvdihDcaLvPrU/Ecy2mP5tu4eUA6eK8
nMcPstS82li5iTLFxBQkjmRrizc1WqBo9yAQ448opXdMRtJvtEG95RiFZ+6LHrCG
QJSSVdtZWmCuHM6bDklgA/DZ1efJwopvxcTAOhHdqQGdPQJGjwrlYeK9tzvmZ35O
bwrxcYYbz8+NmKAetAgbdR3E2mrFV+utlbh/ircLt/vd0jFwsj9tkiuRXtAXWzMh
AHMEHli4uCJ3mMI2c40VnLd/2oFlEmVcx0d1/NQTgh54W6gAhFRFTPLp445p8T5M
4LWBUa+M/0lwE6AJAdEaRVcyXN3db+G1RkLzaxrhSwEbHw3Lti+m9d7qnwDCCVvx
oEgUar0yGvwSqgl05Ie24CGhNhVcYoezbtx2xMx82R8HQ1Ee+gCKAIZsq/EYCcrK
TH1F6gy9TgVI+1Uw2aq3e+lxo6nfSSioEZEGqQRW3VM4ybtwPbREnge3c1yXj2GW
Co+DpODXfObsWgagebl9Bers6K6bYc3h5d+4RPnDTu28eeGDqXdi+rSEdFkcthC7
WoUw5tgiSPY0cidPpesCRZ3aVAU7fdyVWP0XhRew5NIZnjbQznL1vfjhXvfq0W2T
D8LPI/6urdD93IN01O+bMcLsMOz4B+/QxfilxeRjxcG4dN+s6o0VEeB70Y5Kj/qg
lhxPG5fcVj6G4KRbJMOX4Bf58EPS1SsglMxmo0a3coXvc5GKCwGBy4+mbLuqercG
hlmctNm1bKGaFU7q/lJEoLNKiver9E+iMVJaSDm+d3pWFmd3/7mgyHNyvtbfcfxv
9zfQqv7sBVtF3/G/5v/neM5lsEH5G4NTMVb98Z/dKmUaNV6uWtc6OMA7MV1Vy0Z/
YLmCdWIB1163YKHSy4YMVNuh92XKdHBSoxMTUMj0spoFKvwN98n9K4fUeULKUBj5
BKSa6iHtFG4s85Q7erTmZdxiWh18G99p1TXYSaohmTFqai1idnt2RM/mPE7thw+I
UjGWwmJrTZVJ4Kc3m3cSMkANikvrtCtG2mnlZEsOfvIdhlLpAPQ4saDhCzuHagLU
6h+4ZYtBSmKCcoJiCdX1IHzSmBRSJ4oscJM9UOibn+7aKoHMNHAqzh1oquVTqsK7
4OFbQ4q7fgbYqYxnkbTj3EwVw7vKb7KDKjsZV54OdbmLGlQ08U68qwrTrIq5tppF
kmygFLUquNAQwJ6+Xk4Xd+2O0oGVi6gf1Vl7nuVg9bi7thJb7YZymQIIcXrraWG8
RLjWV+47HnUZxilvXNkyF9jAjkrM0BH2yYPIPbgDFSStkS2XltdIOKYz3mmz+6IP
G4F6Zs/SAv19txn3xjb+s+SVH7HjKbxanhCP8YJ5NWF69Hq0ENWr2ajCf8rh9ofR
Q0/v/IpEAayZJb8fl9aq3kag6dxS1/EYbOX4XF6CsNjBaxP77okSu1R/UgkGBkHo
Yu0pIjtLkpC0Z9NMzc7PPFD3UHTWHY+mjJ9z/W7X4MnHv1e1uXhqHABrEEsiQbcV
+BcQ9BOHChoaYvf14+BUOvW8snGjOYzx+uYZvgwD0QFFC8JDDnDx+TN6fj1/k4dj
YT4o5eRGqp+yn0YJVBhnuTRXjZEL851sjX/leZx0NgfyXAQS7XXvDES0tMGXTP7s
yQwlq9x/o0FaW1f9GnCnwGUOFgVyULfv+ZdcQ8979EVqNYeeXXPYMcs9E9JNQ24N
wR1x7woVjvKR/BzeaaYCmIIiJvrXM2OpQZYCuhobod1Istgd0wd5ALuYf+1Zn9Qr
o1Kp3late4WanqFRf4ATX4WxAdhjHRXQ1cK9xSlSN/0kbOVQGymbMUDjzEpM+GRd
rGPFZC1m020bxL6lbPIZ7P4BTpDi6xv8qnQHGUN/LqLttuNkHzBuxrV6u+2tg+Jd
09Rh3yFjZ8mSXft7FfF4IyEtL4QTxDpt8vBM/CTfp6mcpcorAcaw9g0ysQ6JnJTd
MwfPhMZXAVDdoQzHprbS4ZmdaRzzNGA6ny+NTav5rYd76bB2FavARSrYXz66A5R1
sZsbCWFMLUdOwg9lBTzdYJ94/gietUFVf6TAJxE8VjVk1xTomPizQ1LPHYT9bAe4
12p3hxNjNgGtpsXgqVaaZTWvS7qQ1Y9v8JVHQA4+AQ5VJWgjEHY0f/dP4OJ8e/dI
Arm6F5x/P3WNcigOYTCrmZlK6bq2CGbGUvwy9omG2PpswWdYGTi2pGfRrlzMP7ZE
96EfM7mLgiRXT1dXHXBOeZT2hMB4KHQEgqA0wbAD86DekgFzLIO6dOwtzFCGUb8h
FbamOHOXqzzeupMKXD70SlfU7yhuk02a24gjarOfudbVKvugF8lsc3rVDC0QTuPr
Kk6ZH77DavEmRHVSU1WKe/ekyIsWmG2o71RT7ugLJHM7mdTMXXWPCxvqp9kJFTkC
QHs8sdCHDlE8Qgoqlb8KdFyEXbcWIyUF2PQfqegVJ2SpXoyShbwxG9MDWrrJuc//
/0yIJASI/BdbERQfxwr0al+Q8sW7MkAImy4x+md5XsBMSg+rDt+pr+wUpTGr/IHH
XLL0yxUC535qacIQbdPJ11gDyO5LT1QbmQIIAD+KnHvbTc2axmOnBZZmrXwygvi5
Nxuhnhd6KcNnhObLIFYEGveF4UQQQo+byUjP0ZHZc9HLxXUPdE2CpyXq3O5Azx02
/u6/07jYW/oqULbDK8FIMH6ctBMgh+ouG2ZI+0qOnoN3QQ3iSgwaj3TPGsjfV+NB
mzCPTdyBbI8tXV+qNlGGDFeINpo8bFGpYyDwzTUMrVmkoAHRSNCajUTtgBz/Z1VF
W8hOdnJAtxGoy+FX/4c8keRk/QD4kc084PiJucQpTmuTyx1BjmjOOPOan6nPmmXM
S2lxNHEZBDC2Gp+l23CJuBxHEchYNNwHagdHjP942+D2DMsDhzeRHcXMM5Pbg67E
G/nwMgpLiTBrGVTWN3DnBHxwAXU4xVg9GZNcn/oZgOFJt5eDp6zTs3uyfYhZB2dA
DhB9SJ+73m+FqtyPF9nSyi2ji8IHSR4bWhjW786i2lYzYFHTtZLwH5MTdnl7uvt2
1B119yAHU5JN8apZTL/QRW4CQPhT1ILI9nL1wHEj5oxZ4C5Qi28xLbdBCH8Exkze
3QGfZfq1SG7j8HP7LnqJp7A8tYkAC3khtgoxFh2UJanJk43mKTM0/BmgZmlS1xJb
d2gcgumOrahFR6Tm338CT0FTqGNlv9Fnz9Ahykl5fSWqRdKmC7lXCwebq/ArmxYL
XWNt6v6bUWLig2oN4Ma9FOhhdeTZ3kvMd0a0U/wu9dcu9ZoyzapR9HAN1RQnhxeb
/9htR8jy/ND2n20394e8zBuI+Um55wYmhQqgHID8F7cDfmxjI3i6peiwTf+tX635
bAKIavDisk00KHayPo5ppp2eGnvsG4+MrdUOOZgqrJFP5/XoMUJL//fm0vFKJgFl
YYq+6ATcAx7+dV8BuVGCO2geP7TLFaRTVd3RQtHfYlH+qw2P378B2m6Fg7Mb/aja
9geohg1YWEq1L9Zzezo54dOyqT7YGFiiHMQbV9aCV09t/uCYgR1u+EhNE4od7xEZ
UCxKoZOyGeWounRb09Ip/wiHi5q0a82mqAipuR2JkLJeyaUGWGiu4BkBUk8X060C
cLoCGvc3gGGBAJBXGXCr+9sc3/NZO+ISeiUC832vhgWaMCWg7ZOCuQbPMWD63v2E
+N+i+0tTdwma6hT26a9YHQXQwtYtqHPrR+d4jmkUgjGwhKa5Q4URFxp133dkYo6E
/tpGQqf+jwiuLGDtf4aEtDqVn2axvw65UqQ3njWiAcTzN59cTotlRTUssq9gQ6ZK
gy798S+Ui/G9CYmSSZgMtpn//qSr3SFVpDOtxYk8lRb6uMSpOe+UY4h/f0af6wl7
uQZPa4a4DjQXP64L6D+0kA0oX0x32CFT+rLOIWd41moy+aRBxCRBqsqSl+FofV8p
8EF/0pB2ET8UdH7UV2s29IKMj/1U92CEvOF3nJD9hiZkMWBW0tBhIt1zQMwNxnW3
cK2gd2cAP4u1LJ04Z2+GYfvyGwJVjrt5Vnotu2mn9/kdB1bTFeYx9O2OjJYhGQOA
Y8C/1C9aA3xkEbjCMX/LGTxOfstKvL7ylwtRzbUCoIvrUV2IoRWLn2tGWxUegPNG
IjJqFas93vizIojlXinavpWqhSD7m/G2SYmHTp/lT+SPrSgJA7ShSV53Ly2M3uST
MndO5f1mxM3o5FYClUVS0BefZYa+/xe4mg/UL5YM56p2Y15JkiTkQQChjIwA//1z
486AauLCI1bfUn/L1damIXdl62yDVqbmQ2chLAi/zhsj4F7LHCEMnB+SMwe1jwYo
bdMM9PpRkDeeYPMmjJ7d/Jr5TTYW6BZr9DBMCghDYrdwKj6RpkT/bcTgtQwykYKA
Ox0wvdOjOmOLVuVy3IT2fQw1pGY/atcqROE9M1uNag17BK1j/noiVcyYsAteQ7Sl
KwJqB/lPHVazdg6d5QLqlSGcWiuE/coZQ8ZuOotRUuxg27lL3V1V2rWjl2lLxyhr
Du0u6YEDJCHlr2XwT0CQb9dMH/axXmZL9HBYuysAaqe/1jyINKRF5xW3f5p8hlsB
AvNsDSGtgUs/Cm9QKLAusHH7j1QYqqyT5G2lpMiJEyClcHHemJqif5srYpNES2l2
InRwU0qS4wyU5cAUlCUqhJK422eKDpTUBoTa3TsLRWDnEQ1TeMrBQyWCHr5ekpOQ
tiBRqiGLRnP7hXQKGe2QMRpUnHeLo5dV5FPyKqbUu0bJkvNz34d+kvfAEnar01FD
H4JhfZknpN2DuZo9pQvgrKN6WAa/isp3dGiODRJSiOUq5KF76TWPNdx2vn1+Bvko
t82Q25usXEZq3Gk+f4ak0cax5CaCK6SDhirx2Wy1S+K/ej7OxlqLZoS/zCXFQ1cN
cCL3MoIIYRt9vKTm7UQ1DBHpwcqCWxuGIN3Bh5dDZHLWUMhk5IR7mMeiqlj+K+Yv
x2Dzk+G+8prAxZHG2DJqZW+zbY9PdSCMNS+FBTJVs0OJ+Td24RpLIPzfYQh+qyqu
c7wGunBDz2Hn0aLSfvcJ4LCOyifStFGnAxbjHhD4uaR0h1lQGXNtcJpvr7VTHQY5
hxKLgdtORROT4aKgTxlvb49ExEjvoHRqNsqv12stD9OASRW4PsJfY2Oo11R4a8oP
Xo+ag4TDVJ2HLX9kYE/4DC/skekPy5vfoh36j1oSCT90Ej00MJPs5hhEX4oeTzPg
r5QriQ48maQ33kcXLTcQEd/DdMC4SmiJ/tkxkDws5dOXFvaqQhSgsz/j/Nuhk2pw
gAcmci4xhzpbqb5iwoDN7EjenTKl3nMUFg3ZmmnPtSMpo+91BX0rFfGs/VAPSV/M
jydE3QrmrnGI98rQew5CxG2GxYb1M+Nh5x6WH+xk+BaVJgYAYaNGCyu+ktMF5aN1
+iy7pPeMN8GBTzbN1ygjGVNSrRLyWZFg56Oe6u2ok6jwElbLdOJTae98p9V7uV9D
tC8E5GOKec26ar1bcX3pL+mTszZPRMymybYI0gqEJrDFHro3lgcu6+3U//EjkJnI
sBn3LITBXeDzDdWGePLHAeaZ2TNSGSHr+QskoHPfVMZOPvVuh3svfDcFaVRb2Q6E
sm/yRr9h0dnAELtPBVVtRPmvuh/B5/8Z6GUvzrXlCfHLapQMZbR59+00TgmgePRG
yrzpiiQSogg6AAfhSploL5hMWbroSRqEY43oErXnh5+3PdThU6LfEkXmqA9JiN62
zennpA9H1gcDcXkTGGUk/01JdXKsuX8AemixvyLO2yU/459N6nsjyzEqmsdfvh+R
njXRQ1ZQBBGHIZJNRc5G5V0CEGyNKYwLAphIYY2Gl/Q6WR1wu8Cm0rxWTfwQB7RC
7KSQJUs8Qc1tGsyAnOfTNA30aT8O+fuc2NgKBu3lAcFoeIJzm3wmjk7O/2Oj+8E0
TTlJnl3w1kTjGCVUzN3FzzSrWsl1b8xjxBnNFbRlQ1lBBJ8aglxOhNpeLOWgGQKb
5U0yQQflK3h6B6x9OnKp+8BRGT5/qiV8vEDWa50Jt0vCR9d5+S1G0vHPk26oIaeQ
uTJvfyyAYCxrORqqsSqnESYqqQqhbuWBhVLq+tmiPuBaloV8RSkaA2Lvb5InimOZ
5Cbf+0IxcsTWs3FDXvzEufgWj0wK8Z+Hj7oHeqgNt5Ol+xbqZUcwZ70l2btypA9a
a3Pp/izYP2kTGncQ7xCJ2lR5kw5G37zUYItxt2VFBhcvxwIXjuSm/cuaV4VS6J2L
YCmktmxkZje3iumnftzdK0PJ/+eOseR48mb+MPD0MslCQqdAVpH9btbDsNzEzkKv
v7GsolPns4hxQZBq09igBZ0Z8zjctpqq4qNEswfQ2oR7QMlRxGMaRnYhUPVZPq9X
kZYXLAER9RmC6GMHHPMbCcIgN/CNdrSRVao6dloZdiJI75rjRAoNouyQ4D1HaFxx
6t6ubK0Ywune6I3NVvyruGOk8bRLfqQUkIjWktbFR1XCTB1J6/CvMzCFwTTq0q9W
wH8CragvwQQYFLIoSUHn/fJY786FEMNfm3uyzjSNI+AD/QZSWNWJpjgKIN4xnP6P
S7dNFRnMZ6GIXUd06KiQG6SpHGJZuF+vWwN7gxdIKbcvvbSRKTkwgMFhBtdbvghV
VdvqWfI8CqfPNMqFNiQ55HLhLpP+BlxE4rTZPeUd78TpQxontSgAV3CPRROqI3QC
/dVwTMEdHxns+M+j15ECh5gwrpNnqnuwslVA5TqZik8tIj2W/OacL/SM8YhQd+sB
cL3Q9x8VbMOiSIgserBKOAkMoFPJ7SORjsHhmzJc7MFl2pni+6DxvOe6dxIw0awU
wNnHqNypLuXea3yQepGUicmMmXvMOC0WJrfrVshU+NendDjXvF+uMcd2JNBlsXc7
RAsYT0xECDQM1J4wnb8zP0YDxeh0JhpgdJILLyiyz7olmkY5mKL5yJK/kYBAoHQb
s/hUuylU9jeUsG3MDgHvrMyxIWRUQFAO4RTRTNuDVXHkwvOSLN+scL71YDoSHZ4J
Qe4PjL9EZic7TZGOiO9j2FhgvOZGEb1xlXgixD4Ulz8vduIvRVfIX90LygoIPGHY
VAVtc2fqjlT2lU1Z5yRyj1pDqGg0Vh4uG4T71G9/KdxumU/ynZa+OFMKATU3K75O
Oql45zJRtKYfgTi/liSPPXZ/k89Jft/bm09qjI3WAFnJI/teSOVyyWKvKhuimNgR
WZRwUBPgC+XROVBJdcEt6dT2gADD4ajCpbNzZpqdbmaFHXUso6d7kV9PxwWgJa14
J5SE2+p9GmdSNQDFaTIXiU7xvNTjsKHeJJ2RIkcKxIjk4kiDVgud+6UE1bgpZw0q
xijSXI7J+jnWUO51qHm9K6sBPL/BwyEIxIQNRvNZszBPu3sRJGgC3TqEglx7NQ2J
27pXXqgHUKpmwWtZbahrYd9b5UfRROZr/Gly9acPr7pQcXJx8+G/2ueiHOIZcjmC
Zoqoy60FHyc7lHwWFbUwOuwu6htV6KGcMoACFs+xxrsAQQlLhgdtGXNPRDlbXSdS
YgGzR9zN04AfwjlYBbXmqFr5oyZ0mTp6haDRWqgX/25Smj3buC6fzIr7h8InSf2p
zDl8A6ia+03keaITSWzrbDCUidLPmsRvvEHOx2mdB8lxvzQCxFRtvZ0PwWYgDNu8
kEgh7uxI3x6d4D6TjTPbPo51bQKfioEBcUrw+Q2/ZXtKirU5U94fRhpHv8nTA3eC
zAlTAV1m19ycdqPy6i3RbqlUgv0Vs7sD4y3rdu9awxm42NJ0S+iFUs1WqbJO0LXq
UOf36L0yFACVOH6lNgTHWsY7hA3S6n764Q19li5sv0/1rPrMWq+vOhVT49x5PQ4c
yU8E5q8bS1Gu6tiCEatxiP9ObzEq9+naYrKD+xzjvkBJ14rUDvk9doAnH5EhxrQ2
zXYxfTn5DXXJV80r1oBRwrzlQQtRFP43PC0zCS20ihAawsJFLC36bU319R7Ze+Hj
5kxyHmy93aegyo7xYKFcANi0+JalhjjRkgghgEmhFEpkZpVOQsEklQnCsjSkBKsQ
EPeZ9nccSz8u9LuduladA16RcJZBw1cUqv4ri6KwbB+hhHyipJeHutECTkdN8uYN
qd8EFwnm66xycpCfwVOJFq74zzrGSxxHqtvpqQipHJSqcSoL1ZtsVHAS8m+VAMrn
1ei/j/LzUQBhWKaeVX2zz0v0zWIg9VM7tLhgoOuC1uGU8kGYPeNXSCDkUgQUOo69
iu6HdGIAmde8wygoKOssO6eyr1tfTmzWVedY087RVf3FrlMccv8xzCnZQdNmqg9J
75fWwCb5j9vj6rv1UWTeMhb+s3V4f2A5cX+uz/V+uMjThl+g9PgPyyfZ9nNPrcNo
MtNbfBO3BX0w/uSYFy4FlbQWXVcWoAg+d4SL0vSkfA0embKV5ctaogHant5jVr7S
KkcQxHv98+izjauyzVRn+zrHnHcTkg/YHncQW0CpE7/akoSoKcyrWMpfBetFeAs2
mbKjH2LANIu8lKT+/B2J/bym1C+CocE4FsQRmR4dILjhLSxieUnriC1R/WNKBh5v
aqlAl+LcrnHVLr0worCkddMmmJrWLaXEnAkWLuKol5Ez94bLy0DzmLoI3E5PXBLz
fmvuGnwuSfXW3VGzfaCUW2VpfVz1utsZDbCGB5YjElb1jgXTPoZlmA6AMVRe5gDQ
PNj9P5yi6Boh6zSxIq3R0GK+qnm8n5o58zoWWVIEC/xxnmEWfisVIlT2027IVXc7
+ZY7vyoIVjURDExYQVTKtYqepNb5xSIABn3nWBGrO8gbgixowhsyIgEz16YRT42u
Dqm67K1rsNfd950c/NbEHnXnz6tHEXXGIS0xlSBPXumlxds+m3wGh7uOQ+vIfxp3
uGKu8a/2lJf90nhHdoYox4PHrLdHum1LDsFECP/yuNVNNT+8tZVnuXh0FAqqq0Vg
NIPWGjs7zOaDOX4mZRjmiJFK6PVaP5PCyNYQOZcVALzYPFJIKRdWq/Rs0aLYt5eD
73j/pKYfqjKRsSXdKUtt8t0eHUEKvQL8jHjlSGE3mSF8y/BQsFr4X3P1VRilf+CI
avivLqKm/FDsLowZMhq0cZVl0BmnKXwnLrOs+YtETxZPIc5vbW+YpQ+Uywyja3Ec
JnonhCpjpMMAHoGTxSjZBKJ5vcYT1z98GY23TiOKIA4dLxN8qFUlbJggWvtwVmfm
ATkHHujmhT2q8m4Ms7baVYGgdHcXsdj9p9xUdA4FvbcsF2NTuZUZodDm8mLlJieh
dmQmIW2Rp8Q+PeTpxGm70zVrt4xi99M6D+fe0wrkMky8G056wxB+6B5jNSl2Rupr
0lxuZnNi6eXuo5/k7STcbbTxjFuxKQEzu9jUkF1JRg25h2hXlr83JL6DMmRaWuEO
fQ3n4eCx8zybnz5VwjBTUnW/aLURieqnyXo7IbgZiIXX/isKIr3RpLJR35DC/c0N
OPZXL5JaMyEkV5ptxGw0x/M+93ch3aQiKKxb5SKHwGPLhAIRjSfT7aDO8gWSfgC8
vRmFyZiyo5q1f1Q6bMzfgj0wg9LkuU+7aLHLccFFWQHqX4KTYRzO0CASwhL79X4v
1NZFt7Uk8V3lkxo01/iORl8bDkNGSCDfMwt9O30kbNCcDLNE9EzlKF/eOtvrtQD1
fEaLCzJ7uOTdmEc/FRMT23H/RuZTmhgq/SPujLQHsbkqibPvVKrDhfWZ1GksNtQb
vWmPi6dG+Sj93teDvGpC5nXhcRd+R07pOUd8+MOQ908CfcSqxDZK4reQPoy5qXLT
YCOhzKIGtfgmBDde6MPTSoRD05y0dXwnJdvseK1OsWDCjNT2r/nCUg/Y+BL4pTJ3
Q2nKsIQJL+COmxTUdVxHU+wAPQdLsPeKzutZKi9sj702feG+NKidYQjsYeRb5B4U
ZrvSpL7R1o/xmkX0MzK2c/W58CEw3eIxVJG7rM1ZRqqpo+ws8C1Xtu/LlharEOnV
0uGEqgAPBW8AXFRraOY+Zn4D8lsRi7VEUNlkClPh8PbWDbkaGjSbx0quikjeAYZ9
2KZMgJIEfMYT/ciZq1BykE8GA/evUTlsYZ0LnmosVOgih9UnBQjyo/TOTv1RfVQM
fomcSxnSVNaRMvTRq++6oYu03GJTvVxLGIEtl7TCIMQEx5AvzqRd8iMGui1nJ75n
kPEGmFvuDsNL6irEObvAKMhUfJvTh9MZ3nUmZbMo04nknVB34KRKidMcIprrGae4
cP0Dg1Q6X+/Fip2TOb8trq40OZ487rdN+DS2r1ijPtYZdfBbE7kOyrZ+pm6oIHam
tCCaIgFvqS8WrRMVvz920umz91lz1t6i47B3APBRlGwkq2FTL0juuj2i/7sN8z98
6bTWi2pShT/jzof02r5GN7qerc2RbTxNwK2BdBx9urdEby+PKxEuxpjM7h1wExsX
kgdkGHNW17OzeBkLTdLoaXEMtlIBbJOm4xisFJSRCmkpZu875oclvVSOS7c5pyB4
XbhgTsGtASjfFe5h+UnRA+NABTpRL5WZK95INe6/EupdXZV7/xwG66fE645sv21H
AJyBBZKcay3A55dSRqa9SijSQ9oWI2RGfyFmNv5CfbhkWT1NPmCEwHR418Ie/Vxn
F3iFxXZmBUa65VsF4/waY/UB7SqF/oOv7bTXOzZmS1ixe1XbXd+aWbx+YqMW320I
d55bXzln3wHJbG8qNBdGUFQPruY2VuoZLXD/Pjqte4boAG0h0dgh9bR9DCYH3ptl
TcEfHFJAdEQ4dCRYQunbDRfeD+GWVzNQjeCWYuSc42m/PV3t/A6EZ+b9i6x9p8IM
tX8rS99JYzohtJnkA+PEMfcKGFn/ZcHvweUVsqWPc/SzqPZx9fdHj0LczeSMkMPb
GqPFcyvwZ7NZOjefpwQDZChGhDZhUrSw3L6koErydYHt/2a4cz7y53ODe1YqYTxC
Ai9Fim4RkTyc8Xk4q7lb9Siqf2DA4zS3s1oFQMRriZzw+dzhYZcIJjr3R/BvSmUv
ROVzIvR0vbSbKjD2vYUZPFaVIT8gp+pHDrCHTo3I1fSLx4QBU0uUOxpv/U7Gq0to
r/tLaNjMUPYNW9ni4av8/w/HBisl6EO+ZxWvnhfUoZkw/loOXAsy3wrjDiYJ7XCg
SCESOU4huPTH8kHCoBktonVbbHMVhrYWW12HrAWZJnYuHHZtNvm5RqMpt/KRvldH
oowHQa24g5ZHR61avJp+TxRa9TqSp4qs9GmxCBu8Z+MOJfm91UxCxTCj+7UZRp88
bB9v+cN3C49zmj/EVW66zvRTO07rS0BBWTaKdiVsrA0vaUwx3WS3LFm5fBeJJ0MR
ah55AwsA+5m68H4QnJXbabDtnpVJYUuqqPZwncxw7OkLXa2QFAXi3xSLdehxHRQC
fvke1rpI3IO1ebJCN9XesSEh6r9fnGdjp412yW3+cOGUXuEJ3N3V4skU3gsttzV9
Y3gi0h4BpqJUQ/hHIlQIZsWzwUNL3CtEN4GRtyodvOKllsR5lg+cIrJddQMcCuAh
4lBNbZY1SYQvZVnFCplT2F0VFHlWrF+lV54WvduPrDEs6WEywQUv7ZnK+vA0xCBL
vLUM1GlkraABMYHMYk9utk+kW1fVvm1PEXEmSq/g4/xOiQxNqmnvLHFKfc9C1AYc
ClNnq4tPnaZY6AS/rGB7JVbCvzcOjccK2PNYVLzxJFxH1C4T3qqXIK0UyRxN0T23
0Vt28M7MHMNaj82ctwL7eL5sowP5x38OsYFGZeBgwE2pep57ER4S95ZO54ntyfDb
Yl1V/ITsHPE6R6p6zWTB3CgdbwyUUHHu7ZbmB3PrzdvyWzCoFrtHYs1a2reOxv/h
22cAi1WGO8K0wiHICLhkj4Ut/xe4uCZ8hLU6OBwOTgxWcP7kkMshrbthA0rE2/RQ
IUptl/M4l1OR76oOI1pPE/E3NfVnrYWpgI9H1ankPMvowwr9iVqdUnW3ywVzGgch
mOTOb0obTSuS9GOQdc8w1qd4XWOQ7Ap0gmDj+DC8vwPwLDc1tFXDrpx9/S5xYB7f
/Miwo0AxjD3vD86kN6D+0hfv20JeM5pc4O+aheB4LrjmHq54Opl8r/I8ii+OsMnx
BQzmvui4L5UQ4Zz9htgvy6e2vINsJCDKoGZbN0mFbeZpgeC1cby0zEI2SolEIJDQ
BPwFGBqkLBSVhVZqtiMs7sq6IKyE0MvwRg7uZ86BgiCxyRKMp58K+aGallOEzkIv
h8bUM+OwdVJWUznlcidwRg9dlJ86GoPccppe6fyEPszaB9W/edMIe4IZzWCbFjE/
ilwc6bjhxDwAIEBmQ9ksUD82efLDJPri2fyaWMn+ARkdFAJYbFiqmZRxu9xKMozs
o+jCml9ulYQprye8UeLnRC29DJP+57vp7NeIzbTG8yaXeKT+YcQXJdtBd17IFbLX
RMwINYh1kGV+z28jLGNciTT6wSKStoamn8+oMJfsOivj4/PhrkmAthcLnXVs+lbU
1L6bYVEhV2i+MzDne2eqUwcynzOnuhoZwFFpD4SyTkNhRKLi+DIujgJFUvM29UE4
Oucw3EJmFy0DehVP8rnuJCpPeGryewUyvlP8hpBmU9fzbgowM7zKb5VSoW4fQiHE
N/uQd6rnyTW5ViOrGnEsmk+cE6Fn9Tyz7Z/eq8P5lclgG86GBcRo1p0yFixSZbNE
PkxOm4hVQWcdUq6nRXDc64bnOkTvuixX5F/k8yKM3GILgUDztDF846WvivN3+fGb
W/zCnEk6BfmTT5ipfy1wkmqN7F6R/c+RnwOQaBG0sOhw3aWm5UQz8PcthlAmcL/R
v2gyTrA7wILxX+FpPXIG2ThZq5aA+6MXp40aed1M1t22cYBYVk8kCvTQ2X7zccmW
qnB3KWcBbfrLOfik7cO9PwxHA45Y8tzYCz1f5v52PB/vHdDyfnX9jkNu3L8RZJJS
pkHzHaZ4iE+x55uyyWk4OkLjT+HTayamL/9l6wpkYlOnIoRQxEcwpQJhHwWPt/jy
RJnInBmzFTe9lwjHXOf342Dfq5q/tSHuYYzwZ4iBGIJLXHzO61EaPEMJACH0AmXe
BrfV0JoWZYGfSvt7lNFaqI1TKoJGLlbNCntsGOE4ZG5Otzt91n9Mx9Xnctn++tyg
FXDiQLu3xDJVlscrhoBd6PrstGktYLfv4fkgzZKBulbeAc4kR1nD/mR7WoRWplYB
QuKi9uwOaXdMG9KgR/mM3nVA3mE4NDc6X543H6JTl1A0A4ImhyBcV7DdrbsiFNBj
M7GjqRDPp0j8em5D7iH3Phx1RGsjxcy/O5b38vQ3Gd+k6rdqGlSUv7mlLrFI+y15
GqVPuYVZgieO+ux3Ho1sBrVrMlkpj2JfDb8yJhCMICQzOqtOFkZFFu3i2UOhprQg
esd8n5E0hYa6nMvsysGEa8gq0l39g+ML8ticdCf63da4OSYyJ49dJpmgiWFfALJC
Sp6UR299GdZGNY3dImg1Fk3WXe53m6yTogA3Ogf3qA8fntDp37kXcRSUB4Jm+hq7
MPM47RkFqnsVYcFk2gcynKvfPzwngbvocRtckq36ij5+9GeNMbDSCd/4CSah7MeY
FkK460ClwQJz0z/vic9wb2D9w/A4Z5lYIsEMOQRIuL1eYowUeJngkAtbSfUSwmcY
vVUjU3vcRAWlAhUSEA3CtJAfyer0cAs354jHeqr066vFRsXt2MLo1GPhgve10/5N
phl+Yjl5z1Ne0QtRDYLwtk7gXdigywIraCUSaB+1sPDhrPtIwxvbYhn2V5hmAcSx
U6F7Wq3WP1hObGCE2lwFpDYfB+pBFPDtPd5u0QUAX4y7a8RMxZS2n4MM0dFpA5qX
s93xpyeUdz6NHqqQ/MVpUTM7vSlmRScaLaCnn7HyPa9RAA/rNfLLIKKlyEHDgxD3
h/AgnR8nbfjTWFqSjOBIrGJbQob7n4BwKHdx0Mp04eYb3GCGw76lop2MSPfuR4z2
dMdabC9VeXuDoRj5ccKkAsKMtmc/sMsdfUPYifMEjiPsttzv276y+yLKNT9UK+Nt
O4R4eWcoJM0AdVD+RvmOa0iAec6F/9J2wvtuFgDFhf+W8uJiMHvImTjw63QBu+hb
Dn+3w37EYLzM0SBNNIe9LVRJizcMCTbbGIlsDvERcJ1rQTADyAeOBrIqx0AFR1Xq
ENFvwAu7qvPrfMRAcSw0fYuUCnUgUL3ljhVibVoPnTZy2bH9DUfWewXDVR5izK4s
Xtr/H7BMiZrILNdnTmW1XEWwkYvSGwibKGYGOHHn8XUmdumpCeaekdHIr7yVsu2N
QkFtHdF97uyDjKRBjHYh1B9DvyC9U7enGW+/q/xEdMMlJRsrBGZ9Med5MRlPYcyf
Tr/4QrGLqeHUrKLVpNBcOsUhxYBdmRKkwfwXOphqUi4cWdgbzXr/nXSX7RwJ9Sv2
ImZlx3hgyK2AHLvqAt86vI8UjJVck2Ja8yvn6/lj9QLUJQhw9uapZK3FtMASuGZo
s3z5orQIRJG7x/N8nmlZ+PC81bO1BtLDZKbn7/KymXzP/3jpNE07gtpVsfnC7j/U
HG/3ud91ry4O1DHeoxk9ASm08vryfQOl+NS1mPKuhmhzvnmM4d5T3qd7sNEnZvFQ
X8ukpoKTwrBD5VWW5tiUkjIuiFM2IXfTS2PWc+nl+HGBqvpbSpDKHO1ND1baw0DR
/4twLfHki7J8HZ5hnNwF8pUCkCpOPAbXDsXg5zX62N38kwr63Yo41SnjYVwKDFNW
1xRZ/bvjFr/Y9CxyVXviyqD5CsAtdj2mfy4nfwGvbqRt0KB/1va3khU5gtqgPJux
sYpmpabvD+WvjtOSJaOmUD25h3EOH1on/QTQooYOCYBPhmL3SUMStR1KekbMl3wh
2UwLYGpEb/6PFKqQXrTYCc01seiiakQPwH3dtK3KvIwXE3tk8qWojFzB8XbviwPw
1Y+d3yjoa9GsJsR8wlWVEPo8bJFrPPa3zg986oDD5g0a9CezqZ74jOvmBYtm0u4y
2T2Jney14Jw9YBKbEako2JgMqQSeg5LSIRWIHwhCAY5jNJY9Yepb9XNceN+WlTqF
O3UqI3B/7Oi4UVg41WbAcDLk5eDz2sqfRqajG9C2u2pt1R9ZLu6V7bmkVxA+jNbz
ZyUxl98BTDMCc2bktZSEGu+1u53oYIyPYZPMqt47kAWBqyydiDwPCsEmZLS8X+SW
4ikH5BjfeJGsPAPFTUYiOfmN4NhFmw/29qx1O4/oomUzXnvpVGc4BE5Yp3Mnlnvt
dn8xW/Rcza1HPwSc0wdij/NeNGy/zSfXE9Y4IwA5TA0v2pO7jhBX+XcP7e/s9UN7
`pragma protect end_protected
