// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IhyCPGUuCvCCF7ADPc7LQ7K3HiGBxhmmyG9Qt+bbDzxTpQ38Fjw4oNcMdeKS0Wxy
dj5gH8uE1bEXAfrs1dmjoJkXf7jJDkvB3sRf1de9qzjtfSWQhlrkOv15hcyZfhY8
396i3SIgQDp650b9RhGw1c2uRTXeYqYm7gxgd1P+oCU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4992)
ZItohJOiXFrxje9H58mrN+hJFXQoyZJxAozGJZT7V0cUKv52KqAsGxHMmy0J1q0d
YLTy7v0WtqnwUCdhHxSz4lwwpgYMD4tB7fUsQE+SOtAVKrwH2j89HQ7u9ms+yPwu
xd/6Zwh8KFBpoHyaVrTSBV/3QwY+zkgzKS04fC1Nfkh6s9ML1xyAmsQTrMqoH+E/
n1xwwtKA6am11mpVL8FXQG908Z+uzbmgUkuajbiN34JvjtGbNZdjhRq978QARxhL
QR4SdiLi02WAMN/WEpPGCHve+xiywhdbeeMLI41i4ixHGW7FcKKW+1i/AvRLMBuY
weDVzpPXqawUfXX2n8MVRXbfNXt8usyG5kU39Vj9calr1mZcG+4VoAi177/YIvc0
Ur1WmX9pS2OsVcYrZLJvM9JgdYq2wsRn+vkJiGyefmLkfcCvLc/hk7BMqqX9rxfg
TNX82gkHcQc1kR2urcAfZw4tqWEct+7GX5H/Il2G0tXyVZmxWSezq3nSHCZFPaUM
XH5f9pj4ew6R6LPF9+vgbkWYM+4TwRtRSa7kJ2GFBI7yK4vjnolHtst0vXv6yeA0
t9Eq5Px7rikNBQH+J51gyrR39FP7EzyyOooT7DNdA0Y040nPxuWizCwsx+HvqQVi
PhJofIVCjwVkksc+5cLYoq8ibsXr1ID0JM+DFvQt1hPDd+d4f3Jkd3nBNKkQlHY9
6REK7DUgMqefkc8yDcKRVzM024OfehoDclioNVKjROhmYyd4Fzbqnq8BdEGIYL9M
CWWvEEugOaYnkWMP0Vl4AZxGyynaDniDZubnaBE80vPeQuuIEcxBkm705UNJOfkx
KVbZIqebE06eADaL+ajozLGNWb7wjTZA/scMWWqK8wRM7hvRoTXO9Fe+WiXdcuyL
u1vBmo0UCN64QtBZ/00tRn4Vidlaw15hAUk6VRNCRT+6BIaTNJIpAZRAa6zmohqR
s+9uNLRZiS+qsTVV3eQOjTBG+Vs0snKhhV7TbXmsiG61gWEL2S4Fv3QxGdtHpRaO
6VGXYXqdeoGFjGvaV3pON2/5gbiKdzpszio0/WcatLv459lxsP6o0ahtrZVQoNhx
IHZwxtK1GTvm6HLvXKdBy4C86ozNryK0WueV49s6vTNylarX+9sQaolQdbbRp7bq
ujFG6UbQY+YKEdwnaJZtp+ipq25fnAmiwY3fqsX+9btx+0GbBF0AWXZvKq9ghLqM
47KjfR0MxtvT2e360Yxj3pTxVLYEZCEPOYx1tMe0HEMiGzmHeMykFXb+lpPgVbso
nm/Uhg2YUzHZbSXTrDjO98wIG/hlPxH7jWpPbVY7+D/GmHmtb8ksiMEZzj15LNSA
wcA/NjkShXUi+ZU9+VakPwMUM6ZO845m3Str0Ig63RF5dKL3IKrX5nts8eOqV9Zm
OPnFY7fhx4Sg/EyCDujjDXiwK68F1Nbz9draDZ6ZBwuYz0/vKuIiDoVrATJLUnhY
fkUbdIzVr+bluClKdHa59/330rw0/mMVqC00uFpeozYD0aitv7Uen0qD1WLPXy3A
WWvtVvFD2N3g/VHM0KoIWCt/sFbh6jclWmvJSEby/q/+5KdhviCfkDvRFueHBLd1
2RU9XmLXJ/QFxg98bLleX21aVs/X7/A6AzTCcFbgnRHIwccXYOIsmxcfDvy96Ohy
fFj+KAk/nBoJynnovPR70O4cmH4dFfOWN3TZ+kiOr5fp9JNJELkJZB9A0bx0y21m
CdecZLEdZcwc1xORcX/jYi5mIXXfy9AD3SU3YV8usslD1L7v0LbdA3nR42qNato/
zf/sa1upobzZVHAbgGwPLQVn/eT4hDhPcUAQ26qUwWu48OxDsBL49m2KBYUlh4XG
KLJr6fAKw5qgS04JRm1memqbYPXGPq3DEQbUwzlV51yx7Wkv4dZkWX+BaD27txoU
ynB6laBFcZ9wYAwVfL1MeX1eabTFFv82B7KU2790O+iyPdL7jDCfJNFDArS2ktAQ
zjHNikKRyftpLri5n/zfyZ+1F1NB2auGgj7imuxn4oVPjB54Hxrq3vua1fkaCRrQ
admpVc1qULHo3IMaGS9UPoeIrJD0D7c2+Smg0x442NbQklPUm9smkAWcqaY22DqF
8QEkRWIoBm6Kbffogl6gFd95CMlG67ZXyzvo7ZQCRoU9/7Rd2KmYfq+zND1QNV8Y
xMeZhKsO9iVe9tvZ/4Y/lKKMtuRY1r4syYmXOrG1Or98A/z5knuUDrnHukIfTA6X
9RBvt2oRTo2uMkt0qcv1D+OEQY2APqKiN4q9tsRg510P3oZ6Hs/suYIpX1M+4SPT
Trj9oc2uhN5ja0ERjMlfq9KGrIQvmPpYi8dvNFPh5sLRt7kEhdCDFimEOov/b0OW
CDN6VLVh/2lEI5vSClTA87Fv09J0tBYEhCh0yuz20LoToZzcxsIwNhs1RCTL+Abs
jEUamEsGjMDw0MCqHOgFcMzpxYMujgNR02c6hOpDZT17pwBdvg/swrQWs9uRzDUe
kJ+k7uYafmVw2m1KGZSKH1sSBWKuLT9KtlhEWsQLzDPCTNtzSmWYW4NXfNjRZevT
euQ2LRxZPnbC6LHRjGyeyi8RzzRfUJg5WjoUDdUeagYKr4QdJet+WIAkrl0yI+Zj
PsOmPs+PUIwbezVuZ+M4TsIuGPuacxzfIclyjhvo99yYQCQ23NOnkinOSdhTWCGL
yASxp3rXBsjCnKCL6MPJ60WndkW4DIJVNOCZ2XpAFCe6CLddyLpjTipRg1g9NKCo
atNppnkoKTHNlMEKuU9z9T9da4gfDIM1DOnpwN/VpucyYuMDSwghuOoXUC+6zKlM
V7asyXvb/bt0JYiowmnIHbh4S420YMEjV1qIKFrV+GhgChrGxu8uRSc8X8LwBHDZ
q0cE80vQypz9Ow93b3tihsRvPt+QV4kvnoARqAKcNTMtlwuJJZvuzjO8VCWoHg07
0cyjivk/uRlwLmIhROWCpsAzh/gHp9F0J03OlGo21Vc4RUsb/fmj+Tc/o5d/zdDT
7G5fh8MFWl3yjJvEDYnuRxV5B5vyol84N8sckT9gSUgGgDx0ijxBrJMf89+zcJg+
3C8rQb81sm6JA+AGmY+56DQOiNMGhdeEiT8mzNwDiiZnP9jiYBmbxmvBp0sIfXA2
M6SqGQ/Tnigu52mspQw9SVEX9niUylm+K3Kz/WkrwJjcKAudP37F1/wRPTjOX2q0
gdVn0b9ZwJXpD3wR4r3tDe3vdHQmnDRe6GKzo1hibTMEyj51qzZx8hvCZqOe6WhF
GpaQYeQ1MAxHSzQ75aACTbaSGS0hdzXXT3sbXAGBOWFp5h9s3/pYsoXhrZ9TblIm
38QiuAXfCVuotLDGMJwZ0nfKxL0WtyIi88PLBaGPvGoimuukStFsrbelwBmIR/Sl
/KtKfZyuXWpHiSFrvaZ62nmDQ5Imq9jtTH4PaYW5fvhV/RAr8w6vYQ9ZciYwE61y
SH3VB4MnDV76HXGp5CIkapmuafx743Myj0DMCc1oE3oVp/YO27LLKlaQ4i+L7EbK
V6h+YBq3ACVuOIIv+OALJgCwwU5ltjrXYc7gydJYaeOVRm/CJ6MPXxBc/O62wsIO
jN/gOB0gw7xtAvmew3chps7z8Tnsoh69fhD8evMFxEoiA5fIroTXRcT1adUONpyM
89pW3YYHBr7YWG61L0+tD1mCts3NCpt4igd9pmR9IiJuPRTdqAbYnKMrkz08z0RJ
6rH6f0Ez8fwfcQpGIjXs6+If4wZzygmh+Ggr71ZezAykbBouWlb1mrT4WeW4sUmo
Tsoox6V+PPQghiC58XHCbaB2h7co6KkTbR9iYralrtCw07jANjbg+Ct1ccJnAfvP
/azmvLi5zQMbpkVMJGNzEDHhctIDjmD9WDbZHlYuw4usIflXF9Wr61ohuL8aRe6v
rq/VJf6Fkkn4vD/vBSvSf3AnrDKHOoyhbYHzbUzrvPqbKUgj0tCOtN+vC8mWe+LN
HDj17nf+WVKeCfmVE9tkioqRG6jvoarfqk8eq8c+8e/dsMHgRdWbMacafpDExIPW
rtgOe8XP2EQshKb7MiwLWNpdS9e0Gll0o/vGg+ZRJn6K9rUDRoKrbt6SeA1HxXxy
Chc7mZBnRVtx11394F4dxA9SZwW54apBzMQA4/HTggkx+zVkv/hWDLzVAxfhy1en
RF/RtRgzyT6ylIgDs/tCCAWfKvFNATShqtt3HELWUh7wr1lpom7+j4Ba0UkG6yfm
DEaBeh3B4tHTrQULLWOSb9+5J6+I1wk5GsgDJKFGkyeiGRN/Ow/xLEISWcnGE7jJ
3qYWRBaejuz5YWvG1Qat/plzaUnanVo+P39hLRhOwJIfS/TE4xCNf3kt9XrmmTeq
3Xo1PkGwzsC69WYVjo7ylnQ5aCjL1HTlWpG7Eg+KVgQg8sKswKHAAVEB8YSQCyry
kHDUoNIO/1r1AB7KzKaEuY9QsG3yPcO2pT08a9e1FXW+x3G8zkbX2ISTx6MYOKdo
6G9jQi+md4o6HEfAMriKVxvc8tz73XRBl7+6NxI7X4YIIUAYkS131PBenJfCytVq
mxxlCNLSF4Aad+oEH8L7qtlZdSTjc4B+f/CmDVLuuclkjIrmCZWspYcrkMhEON+v
JmheDkMJunGkrqdCnmEC1QF9vMQWus0pWBIWKwXyfrlq88idOexqgZErTW6Ntfgh
dlddqVtOjE8pf9wk5VtXHliRdJLRvJXkcG/POXOSXh8RGWUTjzPE9KdroKx4z9AN
ClXn1/bZewAcLkk8wC3vZoF03eBamTHSi5L1r2Y6ez11milvNrOs2F7zLXyvL0L0
LNFUsO4OJD6s2RtXJ18SDXxQGp5dawTJu0P+R/dm5HKxzPWQdLUtufvpPg7pN6SQ
XuTq189FqHzkhRrjxSMd9nGv59NqHfRuspBR26j502IUbnfEOqewn6hJizzOxNMi
/wzy2IYDynOgjPg4Y/rkYyu6OLmRhtvTfT9G7mCJDinZ6qKUSFqlOy7eeVE1rnVl
lgo3gg6eGiK9x2uqScCFwGYAtJaINZijoF21NGR2Xro6vafrPbda8ZCe2yUfzAuu
VcYPwTbDkJyNof3KfV+rnN2kC2uTq24kn4u8JIojPG4ewbXpaaWXc7SS/SihT/Bo
EwY+wHDTyXWGG3QiFpZBDsYmi3QaKjfJT9KY0hsWeYql/fEpGuCerGA/MFUtEcIZ
tsg7NsWrkI1e1ZVJRoMfEfiSrt4CouOvQ9PtqTIKeTY/Q2PPz3cCD6zjA3Luwlh8
lXmCh41MmmRZlTO8ZC36cHGQxjgkGOp6sgNVgormU665e8efVW9khGtWGJHM7Ye9
g399y8/BWy03V6Y8VUL5o/BTIFkbHVH6tJR0sXrbKJxCNSy5bMiZ1ivYbLtoQSSY
v+6vtcEhWPkpRc9am95h5sS1Up3q0jWvGyBEndXXI37FVZ7jZFn0oLIKQGbuBoaM
E2KLpTGfkI34lJA1WtMyZBpvch8KcfSg9Ktfrec63AeYxOupEsy0Ln1f+7nz5au9
/1PU4zMx0giwwPg79M8qP8q91b5YW4QcTY3ZlgqbJ+1LnFYEgMVnUUP7ywRO0hXt
aIJBGFEisq19rOA8DdoZjxr/Ep/sVcYAlet5Tfz7ZeIDV/lxf5Ff415bNm+TP0sM
LLxBNeeUHKzrs9FHgn0mJbdGHcKNcLjU0hkfQwoYb06fBzNPBCWgE5iuxpQLJ02S
YfiQIDnqUqlncyLjya/kkuHJ34PsIDITFXY0XkECa4VwaWOL5U+bAjKwE9oLD0dU
GChWpzJ6yO5o9v1qMSxdkaXR4uWBiLH0RSZf2XtNyeNVuBZ3LTr9sPoaxggJ6g/t
W8Rwgd+Y9uxUHvSscL1oyTLRBdqKXTo8Dv1qppk2dh+Zz5+3ATAp8wY+5kUnTVVT
uN2jj/gjATwG0bcnsLtfLVfVpbyHeahmcvcUDeECOHNV+CrI2k15F5ZaJliHl8Sg
TbTJTRtXdk7Lf1GuszGCL7PUE2zB3YX9pEnKKEKHyNcUqgxB2vQKNUy72JaKI+YY
F34y91qUCZNfZk2eu7Rvqcd5Lpp9TY5WEWnVLAhUdz7W1tfGvN5U0jbjL9vIgRds
3vXx9YRIM/Iinx/gQ2ksZJ2mS8ozQOeT/2LrCTJ33+ozpO7ppG57LaLiWma9X/zw
PZhuPHcMG8X/mI9MkBQod6DTNQ/XZUlITEr6ikH7WILrzAYg5UlLfDQuKYjbZQ1+
wkpPlKldEt68E0Hz6hbxdt+0SWxL7sQAanNDb7SrNcjt+ccmYnqDFLF46jeChR8w
M2caQs7h4cqeA2xtVRYr2qE2nTZVF5Vf6bKZsnOAp7pyypP9Vlw7tdY9duUGN1NB
87ZST41p1OZeDZH21iK/8Gw3JYpawYJ4u0/CK1nkryA2BsyMD0K68IBLN+e17ysP
TtPBBQK1DFEHVv1BIG48dlqSXFi2FPKPeIOPo+MU8gROAylFmK/ocaMWItXJKnxh
Zpe5OisJvsRU9viufMZkTymE/xjdUe8y/K1JvYFkxm/c013G6UjDawJwEY5rl4Sj
2qNpqnUp9MW1hFHgDxWUVRujx6g+VLdqSQSZoJcXyJn9nbWpr1+bu4qh8agJwaJm
GGY3HEgv5L3hOif9kJXVduRdZsr5EBXfEjNhPtqHepWbA4ULiApICuZLgnql9bAZ
`pragma protect end_protected
