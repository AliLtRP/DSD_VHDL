library verilog;
use verilog.vl_types.all;
entity half_vlg_vec_tst is
end half_vlg_vec_tst;
