// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bdXos50OVVWz6Y0eQmh4DDY6AolhKHMOtGMokkbo77p3aPH53kp3lx2Su2aOspmq
9+NzvE2ScG7sCJSiMQtcoAJce+1sdd6tgVoh/bjEE53Xo4/0RWdb/cg6/YkqzcIg
FRRuSZ6vSgoRFXT9n6fHK1dt0FliPOz5ABQFvlvZEOI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8528)
5zQhmVxLTAScOgQNrSdy7mklz9ZkOnrrg3DC498IDogUSc8srwpAmSvTOp5WuguX
RU4R+wm+uVglkHep1WtYPDh89bMmkJ5lokNyLKAY5ZC0Emu0M5h4PS58YZ+rhjLS
y9KSptO6MBlZ7dqfvFR4Vw/Ezz8wRGYqKDUUeEq5Apb3XRUXJ+a3HP1AAPdodkRi
TCuM/UAc2aKtcQufeQ7jYXKzuxE6zRwZPLETLWS8YCHnibXYtXdUjvCgWToc7G5e
vEcHkkcCfYa+92E4G5l9c0JUeXvsoNkCN+wAGWtEpOeDyhiC0Zw/yQf4tSkjGI72
bJktmKYTBkt4AQlTUM7grzja4ImEEaMJKJYSYLVLFuzj4CfiXUvwXFvqgiNymwLY
aG3d5eQmbFpAbsqNTCY8uiPzEYMtXwJHki3zjzvKrxqNw7aI3zChMybuUnSC7eVl
9v2/a/oiEXG92oTop1oPewALg1bUBc997FDdmwaBDf5fZbeNxdZSJXhaDhxzs0Qp
ARamzt1mKSPkgUzxWjmPh8qvHvuYNLAR8irOHAx9pV3b41mxQNeQJGZET5Xw275K
+RMw+8C0W2Y/DfII+x6+nRV9ikseqKXgRfaLiNERPGfMMM4WIlvZKvgI9EEpaADk
tgX30I1f8tD1w+a6C3w96gpkNFOtcRBtF97pPiZ8xkUa46QCbf05ALBr1BawdP7R
k+xj8/Ln2kHlvKDR33xs2PYFJRbpl75Db67P//skWysl8C4nR+FR80gqT80xSGM4
KM/oppr4yDrWqa8Lk8ghspM5DZMU55LEnK5zptrqHPynzDxzD6aM2S9sTGsL9QWm
p7MUx3cM1+fSlMMfqH6cIVsDKNpLHbg8NHNNJ0D7ChlJGsHW3TEneYlCO/QCaaLy
5IHUdjMetGcZd5Xbm4S4H202fmtfHh5twi7GvayRsYRMHifpDKept+984D9mFMdJ
9OmBuFvfjo70ZVsriyP90UJxx16FRcz5ZuDDmXLbykfrgKXfWhggK0bk/R5YGm7c
1wmnU0yQGAKDWn8YA6ttqQ/gOYtkFHLNJBybFABM7fn3/gVO8kMAlmEAkPL9t3Iv
6vLLQh4Qx7TzGztHYTnF/i2tmKp2x4QDspJhehZlotcprwcNBqz8kkkZ2chp92yW
UySPziFTeaMyGqFxBLaxqza+Q53wRkV+akELX6iPgQrvNlm+hHTi7NsFk9IEhQ0H
hn0H/qEEf7gthQj9juGb9OKmCC+yrWZB3YWRmB9pa11IA9lwodmi/v7RfEd+IxQm
8K06+t1KVyS/ixA9GMYBBc7/Wf9CjRd/2aCDl/VgQOR90470jR1ajDcSulkwcMwj
5kRwBNUMhqZ+1X3KG91hyXjxRbC+X4q8XxWlFb3bxQJxZl7JHuH2zNtMVmc7ge6r
i1EolCk4Dx+CunERzlGbdzb8EXQ7PAX22FzKn8ihD7BErgKQYLflA35zBfLnAHi3
N/YW3h9cxD+GnNkeuynrFIxTpwHNVH2b4Nte8Fv9thNMQjHHu/ZKPEp70C9vKqpI
aARQtcCuBX01x4wNgQy+j/ZiDqmGnAzOevqcQzTp6LI8B9mNyIB6RTvIUr3Q88ka
WPxeLhz8B5yy6oj+j453iZZBK5dP+h2Z6EFB4EjyWe76eo0kbC6NWn7+CSypSWZD
st2I4SIqOtjN/WU5Ui/N4gClVRv5pPIVJuDO8CvDOH4mdI6InctBWWnaNAxjDrOO
Fl8ItP+9dPgHHRrxHbzVKN0CsLhucu+O646VfLncJGrU/lkLGcMTJ4xYLxHEtHQf
A9qqSz3MGb4aiAwKTYXrRnR/ELOUC+LEOoFktls9wC74Mnnfw5jIb60/OcXUp+sN
2DUhN00+ERiQD9XGPopDdVk6lub0dGjnt8xLmKNgX6f6MTlg879Mcn7xkuXzdTea
blcmAYjD3v3iqVQRdW2B3Y6r6ZMY4znNUS+ykCAqPK1m8DDApvjVaHl8tQT8uGhM
GH7okW558TC8BEIvHl7JSeHL0cnR8x+lkvMhOxsQeYmTEOC71M2T23Ol3ougzfLW
NJCAa4vGbRoEl55kfI/hJxpmg4g+dkfByux2qQx9SLN/dznAvmYufzi3G2wQlmSh
a7jhQZqaLtnkys8zNnGEluIQAJZE1iSF2gh21266Aa5gK7qsLmZt+PN3e2RDqv15
ieKPxjdiv5Jn4APBQIrmAc0wWIV28hVqD9TFmLPx9IishoNM9e+syovc+7CG03UB
JMFAMhFDNG1fcq1rBCUekdnRJqC1+mB/mhGdHc+rX9OK+JfdnhTuCHI8sQqi4Xlr
l4lh3J3qGp15WcLxhJyF+2zWe+uB1WsVZYZ6YEXqowS2mujtsGjXXHr8frx7v06t
MfgeursjJzcd60ZY50qVlNA6MFUNqGT5PH2b7iwap84kmlVzxwi1fMYednikvuAe
pyoNb6POKXHdbiTdFrGBaQXnydDCON6kU0h6lejEiYMgfbJ7S5nsQ+LrjRl4wopY
inpMxDVwDFtimIMirOTqkk+6Rl6ja9A8vVVSqHZj1ix5JoeGrXEA8HKyJfrnxEwD
qnkHsd+1A6jhPQJOpQnWfPtwv7H7k3mUeEMHB14U40Oxd/cL6Xqn0TC+s51QTdZz
2x4zTza4jOAzSS+eFT4ueyGsCYhgPAYUwWW7Y3T6JBbDkyJ0Lyy/Geb93XPIdV8z
3lyEv2mY2Ew8QhKGGfdyYhV6Z2tCCf1ax4rJDGmU7ukfauG0P+PI+Z3Rt/XQ8SqF
vMI/l720+L6dfFwQm6iYyiNqqt8jK4w+KmIK1m0RP3m2MoWAt2PJAZoP2wUE8JSb
7ZvzzNGBqcN3MOPfN9sMjYeB0NlkPzltpXPBsZyXWdVGkqU3rO+7EUPNzK9aUsA9
ix3MzMs2i5KjpWwRTYOOYnGuSqmkZbmbpjHGC10QYUT5utGlO81+UtWNVnt0Q8R1
jbG+EIXxloTubt1clLamILmQNyBs37xGFnZp8VAxAQkrmIaZBf5QVHWLOYR6Yt2o
jkfZ0SzkFIVymV6m+eruyk6lMJDPtwcHplo2TrwzNFFzgzvph35HUfvpNBMDU9Qp
HlgH44kXXHH+hIbUi6FZsU+li0krb8AKHgjoBbjaZC8SM7+LiqjrN9vx9gZwvOWb
rwpQL4r7IfH0hg/nw2uM7dF9XhXD1bx1Ih20QC8+mDpYfsGmOUSM/nmLDJT5mPL7
AJzgAex6h/wTBJVhGtPt/N09XINmLXeLCPCz5r9rsOIwLfDtNvW1y77AKc/opf3q
9pCEg6h8D0oHon3JHfT7jpni+vw8dQWomEyvJXxi6NatMeUQPM6PaMzE50h8UElS
taCpY1nlfVHfqVyrF5g3dy2Vr1Xmnh+8xPSJuPGvKgBVPSXn0jNGU718/8ukH8kC
N4nlA3wzTXsR4MTnfN0o01dmHCqfiDZKjD8DDx6Tj9oHpWNwIgfu9WviYIVQRm3W
xGwAa4KoukYqAwI9ob0LFrH1rp0g3/ZjyaeVhy0gOsSIXiuuZ/gJlI0/l+LMflEr
2Us7skAk9QGnFHaZQqLBFYeyRvlMoqZwGg3FHVoNAP5nh5mPTvQGXdRu5bnkOTO1
lIhb14ZB0fZZwHhmpumLzUH4QeHX2p9PL30bMxxD0PtmiBDJtlXEKzkUCa/5Il20
xVpH2q9/YWHBGg6LILGV8Unwue4hBKsSfR7DvTPVTMsz/q0KMx6r8V9ponrosXpl
9qwh2EILBGkFHKv1b6z1wZYs7ew9mF6mp2uHXj/KCRs3g2xoehQG1R4Q9kBet+3/
oYLAUxDnIFzo1yiJE5EDOO7sc55IYefx8TyH8s5zocZ1bZOSf/EYQ5SOvsPJ2WcN
clFYgeKTebQ2aaqnvvP9N3/kZlAiRWIGKPHC+hBcLkSyDMvCKFK8XynMVGniRNV7
shB5wg2qvQiLUlnQAzcR0PNySUA40RjOFZHJVjPoKG48VQE65wK7EIHh8Fp03Z6b
kbDf7/Rdu+rtC9GL03tVWcUtOKdx7WNbGcswKoHRH3vUiHaB1zPy6GfpigCeug8c
UlOTZo8NxdFcL13N4d9D1Qe71lx+ORzd/Q7DY3VApq0hnIPyoqaHAR5QVSDWQH4S
vIWqPphieK2JggEGNSdKZzV8sKHkEWgG++KcX/Wbss5/EsLvx2XwWg9pAJXKgM7V
13SRssOCFLZB+28PEtDAKZVr06ENdVrvnWd5vdz9YCs3EutPHx/95n3qKo4NrJg9
XocmjGlHl+z7dhoUQPeKPmGTOxtKcqZPum89E2Mzu91rl5OBvT3+uSdb8m+Q7lPd
0hVN+/FqkWkoRKakVeaPdN8K36DrYiLkhN9L9p5oa4jBGAcLkm+0bubIQRSxoiAl
prbErXxnwf9gVLyKIqzhMMo0O6i81Hi1RexT/52cSXxqMH4vxAJSaH1Jv7yZC2+U
90uoJSx/njx3FFEQqLLy7c2BeQxfVnC4LmJQlM3Vpu93uajFQcWNeAvbNYQU0rwj
WKMuRhAlafiFDw9CU6kIN+lZA3JhZhq+9cyn8gCNr01GvK1fFVeNmz6sc2faD7q0
3fuoQIpvaQjgVZJOyj9ChfnXiKuQe2jnufAhOGs+mwh45qMCbbBE7SemhzlOn8TX
cqADvbW7kUdeP5GiPJR4i5pqAzNRPj5odePUUgRhDcEk4FlZhSZ4N5d25TouQZS+
gC7U+oaFpWpOnYqUc/0iDkpFX0zB0oo9XRbovGnZFTMIl44GtZCB0HZMAB5Brqvl
xlMO7qEAuxHhBIpBJ0EKO/Q/YT2DfEfW4ZZ0zfPH599Q0l2apkIdLAWJv2febRxO
gVoLJOoY08v8nmTu5TIAtlztRK/H3KlcMyIvdI2OdvLQJkZxS+R2sEX4/owzwK97
eJkuPuU9y6B4b/HZMTvp0xgLXi5ZimUZ738c3UpM6QfN5kMhbb3E6XB38e7/a1Jv
FVvn3jgmYPm19EYlmWdzsDQ773KzcYw9qjP2o21Zdv3pSafAfUKW8KQeAnswZppf
uEZxmS5VXOLPJn0iIOBQuDr5RPV6vlH5RGUn0Lgvvtcek4cqXsxVVD7BQCx7C5Eh
8xLg/c/Zdn3M6ObmElIAObQ5Iw47l3SJ9UYE8QKT15He3W6n0NpoVKMFDc5yJ0tA
SLfiOEVtaOlpwqj6tmTWFd81Qk1QRYpTZz82xoUyQAo3xbnmU97mwD53QnynStms
XSpXT7fOGY4gZJ2CDRTEk6S39KTYRqzCfjioSaxHMWtiSiHEXdov/tXXqo98gC3V
8kks2iK7x9mbTlE1jExzjphZvK/rOkhZxCnqykMOlx9/7sDQbx0pKCW9TtIIHI6v
TbvTI3CkhTYGiwNH4+qqCjD5xvgcUNxmXIBdvt14oMizhyTSP0EBiGzXtfx9uhD+
R6YXo41VKJZAF4dKSxdqpSs1AzkJrwAa4fXrC0HK7G/o3ADDyAS7biZiQSQvLkiY
HPSmIR2PjUnyA446HpB2vy+fMvVXL0/3ZSDI/bnIslhOwB1eXJRyxYc+/qdlH8JR
jGDb8A3wnJN9H5x5KyHBDUBV53hBWeHJYx3v5cy0YQGPRdY1clDD3tRvOBiSbeP+
BDicpOJwuXW0sFW0Hl3Fc3olKwV7DGIMT5t3aZPNIJmsjuAwA7vQP8oT+Krfi/Zi
TWqJDaqOmcAeeeZA41hChamwywVNGw/Z70Hj52TLCH/TvJgJUlduCmh1kxRApOCv
kVse5gjvXBnI3QgEuQrSxVRvrRTsDxIm8pB58C18mD4llXJ9X5Yl9Z05TsaIAZsK
XH32NLvlaMRSi6CSmYAo4Wv+ByUmTDFZmoblVNYjq9TyzXScmvWKfQgD8Lf2df82
iUVI8d0uoXh4JPEzZ4FdT1EinNqhz0uQw/MU5BfRU+1Mq1/S26nbQEs0VNc/oLHA
f4KvIhqdCA8j1hRqjUdGyCg95Ep6wvRk2dw6wu6KK7BzVrP/VXtKdj6xV8gjl69/
jQImrFxtPHgYzRwPubwCv+WUCFXdbilKK1JF0CNsYgWnL6Uo+0AtlnPArRN9MjN1
uwTDJ2o/K/qRsWJnxz0i59CjL4nYxQybeDgBDKiI6WBepgQC8H8WaKbpy+Z9l7Xq
kos7GLFqyjWarVb/VaQ6L1qNmKCFhZjy8r9Z+s0zhBdGtrvI/GKv+TmxD6SS+pGT
d8WtOtXCZ/nIoqBtVSivQ3kfX4jmP4ZtPqvjYiWKsuc+MzJ5QjgC1y42wIvL0r0s
5XgfaahvbJrZpWoscsozF+HsB+QvL7nlLuRHYSGi7P/zSBJ14uooQ3lGIP4YQZ9m
i531u7ooR7cF0DHhMthbyHCzBt8A5IvgIX2LNoL1PPRZXtJRafFyi9BSkO4RTdx0
4jieG735gI/rOtGVzKFmwksfY1jT4BJXQdGsZuHdTVHgFo0MV5J3Pw7YD8IWFW1g
gafz8fBNeRAWBCHnAy0Nd1Fgz/EJut3HvU++0JDPatzj/N+/ZuIV1CHoA9z3qJV0
8o0F9D3apHz+gqhly8JMBy+faSpfH20cEN3WCUI78ksrmjB0/pFVHneJ+ncPEtsD
UhkfMuOz+6wSr0CLyMntH3zYA8uYVPU8JV43/U13vm8Lz0xv0oq+94tYNW/XS4oG
2etn1lFVMgj7OVZQuDYlYFtz6G0rjrhBTOjDRKtM62DoNtXITuheqxKe4DADtip/
4ykl8MSGB6GwzH+OTAPbXdXP3pOoX7L00ArgWq/LdSgp0W2MUNwL4otIRLgjbNLk
HTm2wM5+Kj6FB0XbW0ouc5mUBlLpdP9hnavxe9RIgwDK6Gsm5IZtnoBgd67V9iMU
BtFEYzByHWvGzzSCEA/l+Oh5wNkzohUDQpQQubMafhhG/7LJAizlk/Q5PU1BjiWE
YQytH2qfVdq400LO99EfjYbo8u+j43MTqE9uHlkROQwC3Y6foNmR/E1KmjCqv7kI
Czm6ywDsT/lyN7zTbmWnAzkrVQ8N6AjC27JWJA2vBM6yN7zBtaTs8mpgcf2ash8v
D8VS0CrTAAuFhqjETAbWMBxxZLJxCEsYyq+LCzYYSeE0+Ckt8GpsJ/am256gWFVE
RTP2XvV4auFauimthngAKeUWQg1FUZX3S+y6+CTtAvukoQOseQw/Qq2OUvvl0tom
Bwx4Lrcmp6ljNJtW+XpyUa26wzP28SdIJ0T8TknyHtTz7IVSl1zI/MbKkgKdC8fk
h6kGwQAHME+5A1ek1bDTjc2TFpym8wfF6bYnLsCZ3Xe3CzaHP8UQXLesAjO+6Rb9
ygKbFxL4gaS2lmNPR9BQE5y0Ylc6/gI9Ld1D1tGLxzKO1EiFy0rOtOYqQr4ehCWM
eiHKUSLqV/NTqxbLunEx8bHMciRmKAxh/qlWxdRa/RQul2zBhur5dgEVYekwMSxr
trMT3ec/8A0im0IQURY9OzpnKfHEFjWYIZexxnFnwcsywVOcR+WD7bEeLWMnM62z
eEuipEuzOxxpj9ohOpOHLyKdls3BhFWmEjiCK672b6Yd7I4P2hmnPAXr2CqhEnmw
dM0/F4WZS0nOT+HYWMRpXln5rJlBVTOji0t2GXbko2glBUYzvkEqGVdxNoNp7E/M
1EDTWIBLGBPsT4w1LYO4ZIygGujW5ze0UJ6rKw5rVnZ+wmH53O6Yh4g8LVp/vdnE
0vX7GuczjVhBVimU/XknMsZlfyKr5ZAoJg0LjHM8NlVZ5XNGnagpYIsMzbmkURcG
yVu+p/5fNjRLoHfy7dFhduu94rB+kNJfGdsNH6WKIlkvIhKXQoIcSo92ptgH/BK6
VOAYeQz5fGCfXMTCCDSfeBhUj17qV0K2pPCQJMOIwHLpHkByjWXobBFweLdNFc9l
40vpvSaF6sTc3Z78BdEFPJWSGo96zjT0tWJJLtsKq9mH4ocAly2PKTD+SU1ArIwl
2MzvDoGCGZmxF/MnOsWcE38FBWpqYQ0YiXa7/4TCSulXjNGMuvpWQzf74Ny+D+9M
em6jMpofRkKoG2dIF5Lw3BthtHbu/djxNkJkbE1dW6LxVqI1oSBeJ1ZWcIp+MRFe
tw7hTmiKWvGDP7FNRBMD/Dk17x+DyYp0TTAZkfOTIBhH7dCGX8CE2a48Rk3QCET4
PmvSl8CpBIEtfyNOHbaEHwa6Nl3LGtfRqg4HlFf1PnDpNc9gr/ZHRwXgmD8Gpx/x
ftHjdYrTPDpOByW5CJn1szKyHj3L/FFNQ35fPyMvnX4DgNR7aFIWy+OZzY349deh
1hpV5LfSCMBjJkhCgG6tagbOw7KMPsXqiVgNPhjsF89ym0CBVaIH8Tq5SZNMoOQN
9LSskX6YTc5lPtmedk1ypuapGCXG4YKnncAifNeKV74k0MeIm9+TJYVqWaUllXYL
ZVhOSovonifjEPXxE4yyeaNvIzOeX1PGk1+UK2TimF0Ydonoie1Q7BVS4enST9Fj
RKQ/9Kv0PjA8O/eU5sC4rUnOT0wvKlz23d5l7LxL95vZsohmVwfOZuRXqUhAn5pj
RrksgHiVImpI00TKdzcxHy1o6/CksBDTGGo4HruT3Fz+kjSWvY/fHgCSr6RyJams
ZR2/fR4EQefZbxGX6yBN7BqMnLHVxN+py6f9XVgjjedT1urj2HpbrYKNiIAZvf57
NacN4Ao701t0zIfujDnN31N6NdyzXmmXfjbTvG5njCldODvsT6kiLBinDfT4AQun
iXobJ24U9RCUtY/VyUSR+VpXP9BmG/1vEoJttTUwYGY/jU0qdWfYsPJGBJOlLxMX
3gEiVpDSKk5r6KZr7pzSR1F0LeVRyEX2b9KJM1mvxWaqeU7aDt8hFlvrn3W2+m6H
fAwXAeZPzq87Sm3rqDN5jl9qSTmy/ZjKN1jCCw7VGQ8L7QELtzV9h6FGie1pk4BD
QsFTiX1RFH1mpAgWc086td6Up+HpdNF67s8eC+hYhJULMJzzzChx/krsuT8+rt7l
CFIWy3EuPJU42UKzC+W7z8zPCX14MG2U4GJKJY09jkYnx26QiMnWVdyodxx+4HB6
KmbM6TuTwdpHoJj8JhlDsJiII+B21kyMPplT9nkV+WsTJLSefuOYaWLRtXBxyhzT
PBQMCoexht4Hd6J/96hfgCcE4PyaPowu4DZr0gH3WyORn9Dz7IybGHx9kGdgtDYJ
Xo1kZhfe1yEZ383bU0gi6WckHahAoC/epMXCFX7lGWNy0crp1a9+XCUGD4R+7VQA
2EAEgfmqqC130tHuGIyEFtI6/bKz7YI0KRwUICcgM7TKZScoDzPEJN4MTLoCpjZz
XBeVchgeThWXQ+ny97Cl+grzKKhHLRQxOaBJknCCljn3QymO8pWfoUeXArZr26uF
fvATVgqavA0X1k0TsvvnA4OO+1IVBozZ8xzFn7ZsuvYPraVhqB0kFTmvIf/Qb/CM
bUVMwus3ROU5PsDf9mIgGlxg9rJsZMl5u9Ub+fnfR6U1KZKR5RFeJ9cjA26byEV4
e2Gix5fEhQRFzns/52VUjNNrV30oL+8ji7b9SnKSPCTuUKvwx7SiG5dLxQcMRurH
Nyg6c8zjcCcQ0PGC1GSg3LhXsIk2pw4LFejRHF2aAP1EYw2CA/j7/graui51vB1A
0yL6BblFEJJFClBlCLoXAYIlfM/RMIoGj7p4H82EKCn1m3N9hl+je4IP3AyH3PE6
+XrPVNsEq2/rNgZa+SlZGihoNqJ3JrOeL8Cq1xZMEkibf/5uyYWEb4audvey0Hjb
8j2+tSvN2KVBZRapi+aNucEMuzS+fe9OrUBjAsvGhdN9wpAF+gqdwfE6qB5T39oi
gT41+qqgwdM+SqSzaZk4orzhh8xdtlftVorzRfUuE+OGe0KyG5ekmf+p55Uh9nf6
u9kHFNiFIXI2PMeAqUPmFXzAQ4F76ARWDpoxkYYYgLIiCsVtresG7l8RSR7y0hwU
LekkxvC6ZVOJrRV0VO67l3yq2CK3UlD9L0pkrYN05BsPGaKBxVuhpOWt8FgMqLdU
wmHxDF5BF9uJAgPlC/nSmPY0MLz8ik4XnBUEexamW55MtuJDYK3YEAUQ6V9MmkGO
JS0/Hv7jA3UeW4NYk2Bv9m2qC1XZ0raBTzHXtRNPgSgLV5RFkfdezEW3LIVhCwR6
dQN6ITsawQu7vgHRxhwRv5Ptx1zwSCPgRH0k38jHCBCPOBySLPYlcyzJ40X6cLaB
0CHp56seI6amW3biMBke8tuYBXpWR8qT6g7jZCsQ1FUBgI0LWCkLD0wDMOzVG1CF
RD2MHeD92H4qBFkcmqO9/wtVbkpUT/+wUAmSIIirSL6aG0H+4LUoIZklg+P1VoRI
EBQFRqmCs/lKA1FS8mnasC/H3SxKGcHRLGSzTSasbZrhHQ/RohSZixeCsFOtj07P
gptZXoygPar5wL3lLKjs88BrBSwyLG7KufaDlJiKepmzmPT2CVuGUvvhtL92hGcM
tHnf8abIONnXuj6XWl1hRb28Pax9ELvdaFbDv3509XG1LX5YrerpROL3i7Mk6N5c
L5VnwCts9/MCwb/IGkTQ5twhB8C0Jf+m4k7jd40wDM/XSUJM2fgdU6d+BzX7ZHop
iMh9u/JVeHBDIKK09Ibx2RE9EbUnUlukezft0mE8GpRkR/Gbc5GrpqK82DWBTXCs
vJ1qjWJ4amfb82zN/7xl0qzNSZKl+UZ01hlkUq1KyQ0jvKeeJLifPrW7umHhaOiO
YrLV9XSPg6flUNq/poUABKwXorJ6VZn7hYwdDTEuIYkTdfPrga8iQQxgMB8b47Bc
Oxg3zZqa5rgadwCjMabDOtHgGeUEePTkDI/dzYp/i1zL5hnJ0Uea3+ZEztqjNf2m
acu1fSuM2S0qzw1//hqnTmo6rB/vW8y2PASRPejfO8C5OzetPhCbC0/bI8ZXhbrD
ZtiHiz8Ae4WKOh3Kj8rPCiIQxhC6t3GXpZfG7Hdjc3+5VlQbcfuci8Q1RYvc2Yz5
oM03BGUzBpLAeTiXu/hrbbClXzmoDUrJ7O0v6voEmAws4+lrzAnbz4XUdmvrtGAI
Q9xRvx5Oif+cp3V0+IflH7nk5d72pbuFCab1KnXA5MH+NItfiwkjcZmKN+oq8uol
WBZ523ufX+7W+4XFmALMZqxBEDYe5XII3Vv7a4+bBW8yPLUoGFwH6alOfNm/YKE0
FN0wYMkxlU43NeDgZU2XyBD0NGVy9mz2oT0lLWiKeNsT1ARo3a/PIzwshL4fRPnM
l6TmCnv/wHxS9u3d4BAJjjsTZ9tplN8dEKtTSMUy/KG4SEAkv6FzYbT0GyPI7vJO
oJDfmeYJjGLU+zTbbub8bIsZb6QbqoT1bp2btOdQallYle3tNEDGFIAdjIqxGCaa
0vQ1QyUjSm7EIZ5CH2Gy5TlqZILsB9jPg/ZJspjOSacN0YbA0BH6uvX8AI9TDUCL
2EnqpTsyMHXKTjPjU4VTJ4XtZCI+bAqXZVLJG0GkccY=
`pragma protect end_protected
