// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OBtxJAstnADKDGl/9AI25sZ736giZ5dHFfVqTnELfge9zI5RZJcXtUktU4SMAfwE
jZk0CcLsffgdCZ2rOWIbbYl+eWReAQHcq8b3pyPI1j/6qeKuKU8E/A47xY8+/tRv
/vXjYXGLay/lJD2anhOj4F3fO5prGLhS3gwg8zHAwWk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13408)
UIXwBLs49jEW2SAlAfpsdM3JMShgE5jJ4oaEk31Iy9NbfP5Scy8TNVCcRiviFzpA
Z6zRc/7Er8UE/In45Isegekq/Pi9hMyILjU+ck9I2deiEaQO3EyDWaP+/jBpNPvD
YufEXLtHNqkPB3Ezu0YPnydsHCpTKwlaZDiVHo/iubf9GAkTUQ5Ax6oMV/qUKcKa
NUYVJE/RXKC7TXPobsmBczc5KPauvawqNW56kHaTC8AA7ZhLXuO9fk9Bx+BTHe0f
sd0eryfYj3qDe+O3a7ghQ/G7uZc7pTgQqP73KZgSxLyPoo+cU9Ucmnp1903SmNYQ
phjxLrPag86XoSSmo8cs1Rw3uBH7XzoQj//wmGjpPRtz+iMT/glDuTJ9sPLrQUxq
Oxb8XDJ9Y0rxZ2n8bmiDRLNVgDgQIcur6PeqBXgh8iJ1pI55P9Xp6lp0rb44Kbr9
48kd59oPlQumfu+VPJDMZC1Jd5G60J0U8fSPrwKGSgFHVdQH3p+kEQKti+279rd6
4m2r2l3iDwK+t9PhCuBI23YmDCCojRlMtLiXg4ZWN9cQXAzBTQyzlBBMEH4nMnpe
qhm6bauzt0MwT/KBbg2/MWdREfsKxQph555qSzR6TpgAwKFzSE1c3SoVWxlNkT6n
IVVWScrmKjZB5l28Ps6hwfj6K1MRQpBQmoZrxLsMoFJpE+K1XJTJJHe/zIX5AzBF
p06LK2bNx7T/+X6MHaQiaD+hM/mqJqNqNruoHaESDtnWBQRIzk7hqFw1ZaZvagqP
oGore2XVEIeGycgFXZghuyzo9mT9+JF8bjn3nfkSz3qudstWkg+fhp7lfUibuz7r
pm2UBw+CXZFoVpLo6hXyAxunXEEn6/+VKsKjyvthAjSKAjs7IgtqXgrKym62/fZe
SUj62J6jEeBS6qJPC2XddCRss5CAKzsOY4Uo+mKQeRuPgHo8KmF9h1latCjOUKyv
2Ios3hWlrfXOSIg0rPRVRnTMSaLdwSP6iVAST2S/9sMK4W6qOTnYNhWqEQS+V/k4
fZZ1MuoxCodaue9gaR/e+3ziNMe5lAuUI1qTCh6tKQLkeUPJq0VE+Gkky4l7VD8J
CDl+fupSiosRXnqwF1pRPSvn6XGt/T3YMWWTZARVqWRYCWPHQwuwXB2J5FCGPZcw
nOJk4XByD8e3LmlakuRK661lXv6hVum+7L3AxzflEGiwliWoQkna1Gb8WtrM9XCH
5gVq0JOy9uLYGHQP5FrjnaQq2txrS7mzDwGbbj6YsYm9CkYVveSYjrL4dR/Ym0aQ
SNFF60iXqS9BLxOCtngROplfBt3Y8wTGxu+uZaoZUU/2AOudk8XMwFYEGMHLwTND
/FeEdMIkuQiYmkAxvA1ZMT4zkusmqQ53hAWP6y7+h3+JasR4g9YUFoWW5XUtPT8j
xGUsmIikRNyitiyNuVYidZTlUmyCsNaT5dFLKOt2MtJFBGOtHSK9Bwl8JrS5fPxs
Hhm1XigRNDRvY0LBRaGCTuSHsUcRo53X6tWueacxoLygVOQdIopixIS2HR64vOaJ
U+lUDLyFOtNWaMT5enHXeSsACcpGBhiyyypQXJKbNSOfuj0Gz1oYaF/8X3IXqanC
Xo61QWHIOTtYsrfR1Rm/QN247s629SQBG+rToRjQ3cSLZFPiuXzchJML/V5fNuDU
64vzbxsy9L/z702CA1zoUAUNGxd2nPx/QHIyH5L1RcEHw6hJPRa1QTx5ZgjZRugJ
L57c9MHIwEaf0SK+eVHM45vDNLyF9a612c2tJBLnDqGgmb76VGGlM1joYzIY1rI/
DGaBIF3MAC45n2UNgTw0XA7VgBfCsZe8+EW/kMS0sagh1cT0JEdKqH4k7fvB3wYd
4evkZlnGcs9YV+KDMGMygIeQRJtA/Av0yaJQxrDE/e8WFF4C52mTVj6veIox8p0I
gNZstPTtBmEhk6qrHtL0d+8zbZcyvGR5gCoCPoZyDZUiiZQjzJ5A0DoCYfIvsJ99
kwb2zuHv35b1xSvzAQtHzQIkczso5ZWFHN3Ko764K2Bvp314FKR9t3GEkcOtbqe4
2DbbijdN4X3/K9KiLdBblWqUXz7+2aFQU7bNKPM/lmBA6INxROls4GVeuYDYQcQ4
HI3MTucTQdDz79rCxc8IrDrkHLOg6lXDijCMk/8EOPzPrF2WNuRGQdHkEts6koSV
DF10jibELNbnsbVFtXJEZoDNzRxIb9SvnmiqCYF75RrTUHArCdwZtAiTfvhIlUyZ
CbKk4Sa8A6+2GO32pPlEsIqP1DVJmn5W8YgUbNjDH1i/kCgqOoarNtmuROQi0OYI
sCd4eMbFk/f0jXUNsDlWQgez071mG3CWQQ0Im91z2ZlkpLVXZwy77CEy+pjeIN3c
cAD8RhSimJ9YoWdowlYTFS2AjoaxRvYE+O5fh1ow373j5k1vebW5OPI1aLA0dG7Y
8FaRsPSBRYQHITUzk+VDzSqHdx6wlO2K1e5Y+ekCOgXPU9MdZx5oZyk0+VkcY/L/
xFzBrzHkMo9F8oOLllSUUPjZENwW90aeW+l6fVG+N6CvXoK6z/P+gLSYGYXFkQIE
rM8b5fN3JTExtMATDfgJSbvXS4kl8e2SZwkm52N4m3CoTg15IBdDyDr5xlbkx6+l
4WXPgdt1NxGDMuCu6BcExH0nk5+RO0zjjyVfn8PKt7EdSvifjE+IGUd89KFnW4L0
BLMKHSWca1rFLdsY5hPDNspuHWcvwtLp9Xk77JBK/bmqa8GA1WSheKpmtbPUKaZe
xLzse4O+xuxE7fzKH6cLRkapCK82084pMCXQxVGAH5Wm5kEpf1LsYymlckOLvUou
ENJNGSPrvedK83uDihiDHS2RbBhrVdRWftThsbwMYDXNWuXP4vSoGXJL6h7Na8zC
uRr3fmgfX2ohAGrngcQjzkKn0Kc5hChLt0JGSzk2A3jpQH/ZcbIsBMeSI+x4mfde
rxxCl8bdS7pjmp+AHhJJOqJhrTXfqIh9Gb8HlXx6BWp4+2GV4ovVVJ9WoHtrUdD1
8ZAliuGpX5+VlIb+FMWH/KQalmIHdQJ40vxB2j4lJkTQOp433cESHMR087y/1y1F
P0gS8z/wKF/yD5U0DSCRNBxqVB4HJkKvp6ro85mJBQ9EUjix2EOX7AeaoW7PwgGb
MpGfziAAK9+GVqNXUn3N613vRXtM3lp6QaJ3F9xwde9iuhY4TXDcwgBItheDBy9X
SVGNEMa9xJczbITX0BAAcJgGFjp3xvjpNEGSP3Q34stOuAAUxERAMIxEPBXw4Mlf
skF+K13cf39hACWUKBqGoiBPUhyC6QvFCu/MoGrm8vofZJZ2xwejgQ7ydOdX/8ba
LnQJBjocfnOAFiIwLElJ0d/bIZraJqBkhI8NAXgjEKJ8nOhT9bqXshb4akbab3k/
vV08l8qixRWx2MDnEXG8BIKMXoTsVw8eXC1E7kpQDgAcYfmlUgCc3l9KiieRD4/N
HQsEEQAMGj95EmcxBb+yVtpMNXtjm8fro71pWw3r0PJhXsvmv+mibsfZ2hPTxkwe
JBAHhcxyVwtHfZoxqocWGX9E793TWrTHtbRzvqIWwrMSTdMuy0JUfC4vQ5WMW3Eh
Fxy/ld2DmkAT0sM+9XpmdGBGttIOdJoCrOhRmI7g62tNVMHjufFz0pe3AWPdCPnz
SCr5EbQ+iKu5Qjd1YKtWI5oOEZi2SPCjz8Ivi/GjWitXY4d5U3ivZDdBZh2Tvwwu
CvFmh7Yo8kPOByiucdzgjyvpJD4cwmrfSyoc6rPiYqi2mWkN4CAXADWGNeW9Xln9
4nqvMYqIOGvzDs7iNhkb8rT5sE2BGCWgeED8xzqj9BoFV/vp1hyRw/GEntROIXWL
CR0QzupOAk9RND+c6JY39DBPnY/RmI+g3T56sZgJ5kzajDgOLaeUkAQ0z3mMua8K
SBdhsxxF8+Rp5YO58DpYTF1N5OO9tvDTNfCIiFrF8nUw/luQMzKgNINdJA5/PS7t
1eGotzAYdcQvi5pawJVNfu6qZIk3SneOy5bzTr5wTQYOEBIYW95T3g9zylgWwseB
BaCCk4nWzy9qlnybZ4HmZWHCV/FX66x8md9YHxHCMdd5DOzZfWfVjdR5jY2U/Nw+
JQp4oUz/F8/ZP4cQc3ijLdLiQHIPBKagLUGlyhAxWm0n+N1b35JR1t7uyoHaUOVV
/QXbi8d/UQZLtx7B21foa0jgWRASm4YGVs4vuC8G/wpMQfq6J1MS+khDTMLuOPXP
dvbCdB0Ouogo3t951dD8Ah0WTPZLUxksQJHOVpzv7XppSu6GU/5Aq5uWHqDN9rlH
xaJ5zTsyXMgoyKe4sO2TrjUe1B0DqrCTJV/gkBIL7z5zHdDMlopFPUjc/8an3uM0
7PXFN3SjsxO69ZPjBWbLOP8ZNt5Z47UAL5LkogMfu0L44gUz3wcsXhtvaMNwDAuR
Yw68ntVN1CnAq3xQpWRJTSRF9UyyrXoZazKyOlK2AMFklZspn2RiOoh4cfMHvTnN
1jwk4iULJn4DjkRFS/H9tcO2V4mJ81fxN1/fp+yIJTQBbzccXQRpkNU2h/dauDpa
5OKLvmxacdrDEOupwtyoSkrPdWEiAEoHuNHUd7D4Xo3d2OoMfmnOwtXaTRTQRAKU
TY5ICg9z4xwc7AHeeWoENsL5OJEtOapRkwlOBWBtLc08SA5EQ53CW8L1Z8vh2wkZ
yOrXRvfnV0fTG1n/7wfj0bR/zEeiVNDHphIubFUJ/69thXNDn1fareyp5Dl/qL8U
FY9iRzGeFkLVMtyXQOQ7lwr5RTM0hfRLmGx4D9ZscqCxjOWvqvS4Bqfau9LMPJBO
jpMGkb30dttGFHRcYYKjUvIyK5MuavRkZcAM2STo/K/LroJ6+tc9l8XQsTjNDj1K
+7rlPNJKvmz2twHYe3jKlHxy7LCFLOsvaJzm2J0GVY8nCYoyuR2eS4Dgxs8mybk9
LbBXSZt50k2eno7717rhyz5MybwtrLURx4I61D85nq4R9byRNMtyx5DtQTPZFfaq
5ejPrIy7lbyLZNUFLy0Yv0iXOm/xxI7WPA7dZ3yA7OdT6dqX8hRVAC7NFZgkVKQ2
VGUPssiQputK2+Hg+/CUhP99qVb/titbgouPqGc+NkuCyN1exIHIdqs/vKdBV3AR
AtocIR9wfb9ZrQGOiAJEVpgxwz8IKESVRAj5JoXCoJwp9YJHlQLwDE7s2Betwq7u
TAPYEZ6IraZOmitvRsObm8Wph/czs0V/7f0ldYBcdy+qYqMFkCKVCg6tfwLXAX6N
9DGrVTaQC/yKWeYkBKYNCBYq8v+D26ttofHJa7Fx8nDzXZwaIVIGSe72bAcJf0Mn
e1fVxSnrnl9wWwqHj4Xxqhh4uNIjl0sAMEOgNy6tGdJ4v0GGobwBupdenEPhSVxq
8IWSLu8xgbbHUq4OZqvjP8W/g2J6jdTharIr/9jlR2vEASDZVDNyEfkjAyAg2RmB
KPVRBrTcx3uX6Xw5oO0obg3a1sn8Mz9QK0K4elc9HI8PgRJgLHOSRn6HFJM+Gupn
KOp5oXI8RExwJIR0fjWg7Tp6vzBBROwfiMUKWBaK/cYRI80CTS5giKxHk7++i56j
9ibnDTYPY+DthdlQCbxS8Xy1js7+LmB/6vrcpzjnyGggi/vGyQIK6E9SEO1raN/t
S6aFW26zxiPmp7GPz5Xsz8q2zHPErpuso7QVCbM0f8EHCx0Ah+3zYcJ59AMVsGul
c6IjZ3J7RKYc/siSQvQwNBIJN3ZL3fFVUQULaNPpYsRQX4CKLMdhziQKG4zZIH43
5aiRAERt+oHNezMj230N9J41SnjlfaFmKuiWHcNKidY4VO005DpUvsJ1nVoUz+py
/chxpVk80iiBKgHiiFjavcaoyyuyYsmtGEWzeeNXvfHVL/7+OifusXyig8HTRbHt
SSRFM5pzTQzxfT31fDLBgrJ7B8FcdQuTQDeSlyqRg+8//qonmbJdhggSPJjLfMuf
YhqAEvNOVKb7c7UDdY8gy7flVmKxNjYI7X88FMVsJyNi5BLG9TXqIQ8LBhmFK4pX
k+fOW+QfCRKnPgjL/MMF0XzuHjeQbWQe5L4uAnVqLpo7Wfb5uvcb5ZOg0InFgYLL
hHWMAvb+6ezaE3JcGNzph2F/ggItRKyphWrKQDvLOV8qeckZE0B1tnCl33VSm4Td
Ms3cHrUlitTED8/ZxD7+LhOd4vxa2T84N0ViznHB6DbadquAsFswGwjhYF/VfA8v
j9OrTPgYebl5wv2blhVdh/hMHvU7lcn8p7H0A7lzxN4uNDAR+qGa9GszezP9Itqx
+CeqjHr/QbyP8u0YFvogQWU2sdziJY5Kv1O6OBBE80sjC668kQoE+Xo3nv2JTpC/
/hAxmkCoiSZgm1lWJgMRnCcYyDXm+U9BKUdT9kQDCV0wNYd87TSQqqgePz9o6D9f
SZssWPN6pm+PKKMlIWvo4oiOaaPRT2oy20atBSV4alNXZLBZBlbujaBO7kv/A+jy
SdTKP1UTFJjjaiRyEl8mjo9qPXbievTtGwXjgGXNvSQoG/GWlNbsWC7lu+uIkrF8
qPvx1XV1TvUNbuwUkB/LqNA2yNcgiv7Lzj2jkSJIIjl3lnSWIUhnJNO0VQAxAM0j
TXtiutblJ/ck3NTAJFsY3EPudbUgxNk61Pj4H/B2IPiQcugajLz74bXrc95AMszT
1waAB5BBdmwrtTN8Jw8Ngmd9Nw+CMGYvV9whTV9OyAMkTo+3AeTgpk1+2c/O9PR/
7wHRQpUUPuE/BGzKOW7qLPxrXrxNSfcmB4rQfTRgOXyYOGmUQlWjMVeIfNeyPabW
vImAcd9OZmHrdggUZMbvXHdEc87oTMrw8DDrxQTB4Qv0xvJRVbwgYzvVNP7Xkd9p
9mO96hkIIXxmsx+tTWkmtBA4xDBgtZCDF1+I1CEP3fQ4heI/DHj9590hSdSUrt0R
jpnh4N05aDV0hHgYnuJjwbzd6DRZbR/nVljNd3PsfLX2/aqTiEUXq4M1ZcOutcmQ
mL/tuT22SaZVs9H+EKX/ducNF1Dx4lW5xMg3h77ef5jd9JK0cWi6Lr1IGlzXjehb
A+v8eVd+55+suZDBM84Na1VRTW+5dvqDWOsi8sgin4neg9K/vQ1rlt0z9aoaoDzF
U+fEaD1eWJ4+HPk7Uer0W0OjywJZh4rr/XUkYP1YlmSrc4vINOzLvTjYocDDxaUC
knBW4r6q05y/6y/mZyE/VxhVuX2uKdo3mI0o4lWNtk2fBjkQCMvflxM0Izqj0wjU
Teix5tAERmq+nUFLY4PD8p/gSwmTtnNxYKrrcQuDoPL7Nqi+rX+bNl00OBTaT1nl
6NFU6P/ixd7scR4Q6dfNxu+vBjTJISTbChsuHZYPKDgaajzj0Q8b1E+yHJ6rIOGp
tS65vFrbj6yO2UmemdTtftHn4X0YiqdAdjoE0ChJcZ79kwFhGAJDFx2outgK9XMX
Jf7yVGOQboTrA9bbXQb1jGrRq59Zc54igAacQMdfZDp910TKru1M74o0dmoFi24Y
GGw3aaDPMQblij3KjmkGR/2NzgGWbMWogx/AkGZyZ35nS0EwHbueXwQHFq9wgLbx
thVvk7zPqw/k9FHWvO0lumi/tRFoYXQSMtOA4432DyAnOstCQOdt0WD9KA0E2Py5
OKL2umNOWJw6Hjkhm9qQKc8QTZ/FT6qWwfsA/tFkZmt/kUtJ/CAE6RNCUne4fiK/
8BPqXk/y8i22kR6/u5uL1T3mFc0jOtdSpvjctZ0G56aWnSmilZRdIzT7AtP+3wym
KOcvZCYP+uZ42nTRGLFo1JSB+eVa0kbjnxvJCDrXLLv4gHYEPEjY5KxTnmL20JVJ
AFCExMU/m3p4sswoVPtJ62rDi3PBjbETmmbobo1wAgOU1RuwWUFFud5J3lpl/aJd
YP9x0hAoI4Tbmkwpk42ANykdcCOJ81UZScIgMxKY7S9XLFUALxD1j8r2Lfx/hcPC
pFVf4g47n7oY5NOIbRvIMOfFLG9wAuJykGU+8jplhVvxbX9XeolKolL5m7MmmYys
WxGVatW5P9zSNDjzxYqadJZobGyDwCTWcjqbmQhX37FRX0ZT+3BZZFblPQ+OCjtS
mg/PZbcILti7Dxu4ZUrY/Upjkz+qHHPkbt4d5Okk8tUnl92y6Amvz1CKHIgVxgUQ
xaEZQzlVHRJlhMH9YSowldPsj0OwjI7qh/XVyllx6EumYiiCkUx3D6MWs0BRs1ia
ewN/JzRIpiUA7cdWpxIsuH8XB8gmCrZyAypjKEL/R0TmHf3pRrGb/I10wt2VaQer
wUH332t5YBTA5USarpwaFlPGejieQxszDJMrwRUGOCHcUHIP20RExwMLnGNENqpO
egzZ+osv/zICsSafuLGBRb6Ffk4Y6ZLWpQ+hKYDIM5MlgecEIEnbCol/Nuxzp6PB
OtdlQk+G4XOjhcVYnuVu/02dMeVXs2Uz8APOhzkYihiB7l9bpK9lT0DERT1NPWzg
/C4jmMR/luyCQ3jDE4/sCarDu3RaZU9ciBmTLbkaG2N8AN5UbB72FNvWyZymp4jn
+KyojsuQ52S4PcFxjeUSbcSZ05I9ZBvcMDqIqRMbDbsWjNBESlU6tiK1MLfr4BLD
BghWFfcBkPzDVd7LeIzcH0c0SEaK3U2rzX20Pdjeb3KPsfFaRP51m2LoMbVjdxAb
yJTSwd1KyxHh/miHv0o0tn1YOy3cE2pHjNoLWEpWk5AbJEQaPx97wzxNn/zoJTwc
OOi5TAfIUzyGUIVc2uFYz/8GGJPklwS8NhAOM0aTfUDgF/vnlqan/vTfgQk6LIPM
7b3r1vK4f9hmwchtAJZ7gTOMr5RYGqsfxdKaU/dy9Mo8S0SEfBansZdommBO0zdz
ffPJJfzpmJ+kpCSqZh14NMiEpvGvrMQMVTPmLSm2zuzALOebbRxcS3JIglWFg7CW
fQypEbd/ZkBP5i0I036T2iIXJAE4hbjo7Tm0lmmP7qRNU+gllclKpMWVf6/sy7NC
cpzuoai2DyvnnekF8mQrV9tty95ectBuomjBSKD/yjCk5CJbJPwrcQA+eKbU9grj
7S8cNq8AKKg/xoiF6sJepnko7rBLOCxy2oygziRIUCNGTnqlM193pnSFmsF6RHQJ
Jx1nwCk4HKKuVdqJyguZro69pxFWcooBXTY9YgBUZSY1rt+GUpsMRd8CxF3iic1X
st3O35s5cYmdnDu/lLvxasFAf2LtHmXQQ66EoNXtlG0qqp1gZUhI//58bhsPq7ex
Vbt9WfdPTWYmbUK4jQWh9pk26PHpKes0ckRt/62+BQrSnX6qLEWsQcKY7EmETn/G
c78td+Bmk6qFvZ8rUZ8g0+zSN3tzzS3kfrXZq+4fTIZBgQCuDaKBpKFtuvv/WH/T
lSepf5MurKD5fPrIZM2ypgYWdewtG9jbKluDXKXQk6HiFPeiVF41wY6IKjbQmLSi
u7H797EHJ9s1iOTq4/3nzo/4gML0TLrJjSWabFZiLa7dtb0bm3n0UK9Evi65Mjvn
MuhRt95B3zfwh76cU+7hyb4vdkJqplJmB+7eFT9CUa7oqkE/2gbtq8VwToKR6HQi
Oe6LFLhQQqBFuUbmvFjFJoJedzYPhQc4Ydh5bpYWXZ+fW3SyB3ZO5q7ESdK6zLiO
dgk7h++5z2utDpq1Jz9oTrF7CLmJztIzLJY6qXT4ZXWzdL40gllHFZI8llbjgpjB
rSciLpBZ8ugU0Unlzun2hAqAppfFXl7KHqkEzov3DzkvicLe0ZE8+8mo5tAuZtlc
ryxz3pDJvjPtUkmApdLi5TFO6FaCwgJBfGvI8k0V3ksfF/YtRRU0LTXy/CoYWcQR
7sKOsZ/8xuQXUYORlaAzHFd/C15wtkLi/SuWo790e+GFW8hSa+IQeF/Al7mWm8TV
CAdY76rIb5dPPjLGI1O3mvbsEbDQcRZWG1wfdOGM8JVB/GG3EBuRjyvtnwEXBb5x
DSJyzy1Z0sCmpM0cRnV/An1jE5Z1nC9juFqFiwsWBMQvWgadODodqpD19uTO2DVH
WBMQt+5l7hEscTUYkTBUjYIzs7Y6gZpwu7iVaEirOj5r1dRMIVyk9SvEFDm7zVj1
MINeyhcylox4KJxiuRrH/HMQfKXQsnoeQspZ8ckPfR+Sq0DNQNsFqtqW3KcIaOXp
CGVxiL/xDg7IR/PjFwwDTRkOW0HQ26/Acgvn98ZBNs8F1UhVNtUNCKsZzkbWTmJE
X3k80nwI0ZWrpTnYnhF3WDchTPEtJIoO5tLl8rMbm+Md9D5IL04M30+YwohmhQgF
NsvciF9PHEfLgYyj2GFeSZRgOk0FxOqJizbn7qes20E5R7qIyNrJy3TCFTqcXdy1
vmUwbJhlmTKXx/6/IAAE6rrWQ+GL7OlJ7JQyEPspZyv9H8eDbY2YU0LMbdb8Uror
ZDINwCFA/PUBX9IZ3G5Q8iCRQk2qHc+hvVnipjB7vYsuYUda/gT6s/mR/0SwnvtM
RUEd+Da8SoLc4lidN1E/NprqLuHcOR7JnCjRWnSAq+NI145Aszjzwo60NUU+dQ7k
ESy3F4CBKELOPap1Nl9o+AheI+CpEttyMq8VZdoNzB1sp3V6ia1cQG6tAz+DGQoY
rHPoqsFQEIN6SNrfsihNRdr8D/gi2HK2dHvmQ/CAt4R7Ck2LoLHbBK3oS4AijZhI
QZiv9McGEo31sKYMvMV5tA851BpptQCFgNoCrZc/s1XNo9ThLmIo6mmY5Dniwc/r
Jt+/C7d16Hn0leL6nfuj0NJLj+Jlb1UwjPfRvSYQZ9mxckBTNfBsmghP/BOsfDPc
Ib2HdKkoD28EuBStgSbX28Q+WnONxbQFYH6VurK4zh8rMYWH2G4dUc+L/D7gKQPN
Gh5u8DIWoRIFQGf23MVZGNTnEL4VIegTeWkXnGibk5fXzXwBb+5Lk82x9R1N0nwM
RUiyRxG3SzrPJTtaGSRAN4XzLznKQA743/piZGXkRKC7Q3vwWRl4xCXcKJ3OUPA+
F898s9x6nlpu/WJZCaUwN8FdVYyukEw9vDQMdmPpYQIwyA3g50W28bqiudJwb81+
fvLGMAib14avQ0M8h1tjAQxFHLY+2kUqH9Zf42rdx307vJWtOjzcJ18Nc6yt8o1z
hBgqpggH0eWPtGZK31VLeCjEJgMUOdl5VwuURWI2aEIR4Nq2XqAPqfS584DbbEJv
GCVJnl1f1gTheWPiXJPxWV1p4S3H+1/QNtOobibgWA2suADxKzDiKUgRFvjb0nkR
ua6kZnnJkFAh6QoUd5+XWox4EUV6QxYAB18DdvkYVkZ1XbEm1knDZl7i+Y7mPsFS
lRkEk9BToKKoRBFc6hVjb8wkkPyYjwB6J3sFlv1yu0tmUIP1DE3tD1Y5pIuaWsfj
h4HXKQe8m9p2NOrUDYmV7WAcauQ5atBFZ9ynvT7qWk0hdbLU2KBgzhzkfyCArPT0
8nbcQA5dVOSQ3oeMzSW6Y+qoj8NR3fvTahWJHNaB4elgNtEb9/6cz8Mn6jX9KY8M
YxUKpGWn4lBtbj1L92l5N2C4bHPA95Z9Zdk1gd4Bf4d3SUm+ujeISbWtfEjpB/ml
YGAWXMJUOgwsos3m0NL4X7vzMEaZuRfPBoNdRR5VSx1viII/GQg3GGjHzT/z2lnD
+2jNi55F/wp0DKXu0nDrs/LOF/+T431bSSO2M5N/OYDl7BHSembWZ3HPs4v5u5c8
1hBO4F9T7eBvyEbU+yddKufW0Qe1vZYxnSxupzclSDD4J1jt+1bEtZRgHfUmu6KE
yzGFtHDDY8gIs9NOlVKXiu6ez9c3TwCdNgAQHPVHQLRO4m2vfATErExQXedk93OT
f3pspN66MBCSBkULcsT5qTfwVxchvw5V0ZIjDAxChSutsnh9PE9zLBB9k3kuAAfb
ox6IQeNI3QWIMmkqID0PfWs9lVPm6V8bJKSmrXKz816W9IBeaki1S15Jamjti5cp
rxO+ZQ+gz8MGQOZc7BkBNaDFAjdRmFHFTgRBoO3LZLAz6gk9BQcF+9deioeyOO7M
i6Nlkf6ONn1Z6an6hjbIOs5dcbjM230mNzM6n9Q+ZWrc4pGbx7uqI/zSs3tj8d3+
HOAtBYSB0dbI+B1/HBCySejblHWBjzZtaANMf+7Z/ohIiwTOy329EWnhUOhz1kZH
p6rts88aWittOlIsrqwSY1sYWbR9BuQ940+YYf1U81fX9/LCaIF5xhqW1mt8dmYz
0rf8nqts7Tcms+lVJK4mXcvayAFkuIDirzXbwzQ/vLmnFJhS3e7Zxt+W1DV2kpky
VCrQ3DhVy1UK0zUQg6TFfYcnS9UtHO0KZS8AgW1y3YX8q6A5FR0CMafuxqGA06o6
aalfRoAk6aZRq20W+CURpKg31uyNyaiShBbZKhQL0Ftu2mp8FdVr0Wunxd3AAAaS
DPEUTXBFtcZ8JCwcxJbRvraLfIU0O1CrCT5hIRkteyIxYYhJ0kaB3t33U3KTp9IJ
Oqk0If2yG/FE2J16tz6Kr/RUKTNrNbz32sDRYNkm8tt6TPmemfg82e1TsSJN38Ns
tnAMTr/JBG6xGXEoJ0TFYB04uZ26nGTSkoFFQ3fByT8o8736m+aI5SnH6cyWsKPf
aPAZ/MHirk/7Q06tZUHFqSYhYGyPzqsxJQ2q+Gd72pqLEbcZekMGuuo5/no4Nlvs
Y0aSEJ+TPPD1Jji+fzlRusEP42Iubljy9i98SDjD8IB9RzK9qh941adxT6hBKT0G
baugjb14ciAZHYI4hhqlLn9MUR4P1G6oqXHXoqUQHcb8OmZElk7CElimex9cUjNb
lf1o84LvKYJxZonNjNA19KyQv0abDJYneoZm0M83p4IAmY2QLlVR+MoxZK20sJvJ
zBdDMZGfcSgIqYkbKMznvVhrVp4mgYpP+JyKHql4uH111xKK6qfzyNwOYjFWJmKo
UPajPzbE2GQtm0Hk2HAZ9faC4hldvgsxn9LnYYjHqzqa/VFwtw4zisziJ0xWk/+A
5XT6vXty1D0wjddw8t8MPhwkbqeyChxrgFIv9ylrdu8B2+IUTpjSnByhYotZh+Y+
u/bON7u2wK08qaUH1o73r0ldOCCSvaPjBgwTYN5SGt5040/oGv4sMxwnwSEy4fHM
RUO7QHwUOtbs/Ih65qm4n+dS4XTEEp9J7XuGmHrbNx3PtNjuciEgdytPdyeObdhr
VYxAse525j8GoaqnoU0SL8jTJraKuEixP7uD1Su9vix6kqPzEXKVGw/Yhh+f+vVB
gL1lxizn90NiR8fYytGi95/A7/STeutHxWXL8Ea3bpP4zQ2+8HETIQKYwQpBFbD1
1a2E6yUgTXNJnxqsRpJAQ0MWxma2hD89Kk5lBS0AeKk1M6Tvrlsvzq3IKEEtAcvR
cBQbgC95HeJhz9C3S1pEdXEPaCVFG4Xoo58Q+HbziOeSVfVgfWrlAyYjhLNa1t0M
PNU/I3N/VW+15Stn+XRivRZ9c4xp4w2mmIpMC+zQ0SVTBp7qjqB0Cku9ukbwLg8j
nH8OuDjNmj0a16h71/H9PMQaxsja5m9p76EZjU/tusI7NxsfqeUEeGx7D2DVP2xg
Y0Q3uMo69Hvv2Q7S61IMaxs1XYzCPEU6AdRPiH2Vp8lfMS6S+B6Q5oVPGoaAYU4+
DznvtWJ0pG+02Z+2whoYArtoa67yF2aao0uH1FIvhU3Y4PQnmeznNg5RSdyA9n9c
gpsppgD74Hi6cg+DcYhZYUH/KlZOlOFQ5ABstNLb/bZ7fsdc2FP2YJ0oG0OWM6VQ
VUf2m18AHgxq76/XoFkUg4K13HvGCMpnRMVOoo2N2crQ+KoL4sxeGl7yDA4PoeUz
aMZSVMokXU6wDuvmXtj9y2c/EKytYKfaRVEoNRtywLbMfKMIlMdSvr29eV/V+5FE
0GbIFsh12g90msiOjKjyCKJLGRY6QZR32o47NlHffrY2nCBDTW0yDsRGWiSskUnP
VTWXTzxbpDmVGdGJs/TTbrJMqK87eEubE/t2XwBxBVOtHGfIxvg5U1GrEvrBkhIR
YijD0mto1oUN9A2PAmARChMQ4z6MTsUdmcZYPTCovPEwmmMHUtJHAS2tytGBWPEG
BTqaenGrRwbyjs6O5AEKrd48znBCijgrfzMIHDZn/CruV3xF218D1HYLMOTUpk9s
eUN9A3bS0PSMPPDX5p7DsDya1uIKQv0UZm27v54nly1rTJkF8A9YvzwmzQ5J5Dtc
YxXqf6EtiZff4ufa5ETVpza1vlrSXo99JKYCkOmvLVVMF7Z4hLrD5J2QKOv8Glyc
vDj7IgaVAVwGPxBRc0Qmfmq7nxFlfaoPauRbPY1xQ/+1sgOxvXsPV5C/dvXj0gmI
zGlWJz1oSH5kazcWG19qLfuPjBFFTP8wL1dLtaTl4ZxOIFZiA7yD21HQL27sErLo
PTSLLpRl4snEyYmdCeZY8eX7ikDfH0TWWZ7AbDQ4vcwu2OfXySHn2KkmAdrH0EAQ
h+xDopnJFUW46hXZ30kf/r6PrM0YwZqdXp8r74lEI5jcMGHaBj8U++ELzlF6RFL4
mw+q0X56diPL7V6Tav0/4S9gJm1X7BNUn0U1Av3r+NTSSCfcLgb+YGL+Vr0Ghxnq
T8fWfFk0sSVx/XrPJKjOZ35bIzK/qw5MO/lTCSS/5b9af8IF+HCA5aU+JVUUbpSf
rFcdfgNrzIn6IK14pZLD20ub9Y23dozBMfZUVADmhCgrjJYCgpdE7TjOPbZR51tl
OnDuxQqTmhQ9LUzegXEoBBu7NRCCPsE4zMz3DtpW8+T5lBJjz10O7Xsjdq9qZUqV
z1NyH0UVXLnPAYqcanLYUYvtVyfor5w2kOlB0lVcMux5JXpFcI3oKTXzZMgSiTyi
/AcCqTDUaZWONjYr0RXryMygzjxFNCwWk8o2Xi4j1Me7En5nrS6UOFyQmTb0trBt
VRntS8WX8HxB/jfAHK/THAB8wtlOygFUWcg9N2tiE+/2ldLMM6ap3Mls19udtiND
katEbpjyDD6zLs1mKQDyf8EDLH/bqrHMX8ZLBi+ugWGkZQ0+LEQjFeT5UP3yUVZD
O/0CvxQp+6VUFjkf6XJ8mrmhxgEJp5B75B9WHby8wclwPlxkcZa4LDSiRpHlAk+n
7WI+IiyBLBkoRUIMzu4Q2TCn5gNMrRc9rwNuaG+9JqP7xDq/3769KqNPShKrzmeG
qix4Ffgn/7WYd2eLjGSmFgJBg9DviypLAHEw5diKYHHSvVA5m3p4Q9zDgJF8tzxf
r3zd89IYhZYXmCK2LS3h9fIFBA7Lrgr1pvqJga6xbAlBQEtWWhrZx9AXwFhxKejR
3whjTD4yETdYMO45aryyEgDTu6zcgwje+58zrMg38uYKN9ntwafvx8s9B66blEu4
1Ry8igofKG2vJPYXbvu8wv8NO2N0930eLctDv9ABl+tFpQYF/5xX/yzucUy3Ck+U
+5reh6YmDKklB3N154N8U5UX7XZEox1IK2V78e3aE70+2NWCUbEMyfGfUH/nOWtk
vHj01aUsnjYdVRlJ5poQDxcYbXyixcLuvr30fYSIHnrXObVfoySwVpl5ubpAaOGl
efDaJCAWZyJlND4Vzyay6c42W/W69Zy6TQlpobi693Iu4Jhsrkyl4egi+vIqSy3N
NkjVBJ4+IyLkr+v9DhjFD4TzgkydCFR6jIlRMPRAe0jgrCnTU/8BjwVWSfMCPU04
n9T8tLRb+256YnkWXsJ4G8mpkjX7YsbOi/mSFELQrGEjTynEZSVLnfDM3sdKAKh5
vYOFornphGEI5xtq2By0PeBWS2MJ/GNYLR1BymEiQbS3OvtCZUAKJs4rmgaNQYh7
kaEqfa86tLm9u7qsp4l8ui7XYZDslGk+PHMRUJRe6qssMIiTdA3UzUEbBCaIwB99
hL4pZvFzagb4o5kcT6ZH/sWYyBBVNek5+Zo2Rlb3lTMBWKgqsuDe8IEvdBso7p8j
q8eCaLJsmQV4xoFbRJXdEJxMyY3n5YWFa3DfKQV15Hd8jBPBkDRr3cWCV2/zAxRL
AfQyAuOEZmLgi0+Xo9ZCno/l2T+7rww7+gEP3n+UgyN3B42wiklRnaHdXHsOSjI+
Dmlsa9NwvivgZu6C8pgzDcWBLfUgTl4hCGn308CYgWXru3wKrezASlerCsh5Yas+
gRk3iK9dO5GLJ8aPm0KEEXh0gxPD4Otaqkn7pYMdKvDj1La7tf0bOpaa2nzntqPP
oHn1YSGqfpG4RL2eLYZ3lJVSanUHLfSq6Z96A/NqCfyCYjaL4Il5yMtkAO3/N0BV
34zIdQuBakyJS0k7xrVgUIN3uJW/IY7uDUOiDRpR+IA4/xxh5BoA/3dgNyRq2jhS
unS9KZhqrAETdLLC9AdsVipUEl+U35YK7urfXSQWSEEyqc/H5Q/nT4AIGUcArMtD
xNiTNANQQ4egzbZxeN5WdvGHYiYJdeToirSaN459wxNXvc2+GcLnfXp5FdoCoipO
+YJPvJJeMMdIkoVpIoweGmoEp23brJ3XvAEeeZJwaLV2PIgeh9iBxwxtv7svMOOE
ePH2c5vYkTgvAlaTt7x5Udhol6dH18nucydH8FKvQWeWXjTXHJoC/jiFVz0iVH+G
Tpws5nrWuGCkLqHRZde3nGIDWkwLp/pjcxkULvWEC/7hswII+2cvX8fC8FM6Bmjx
g1rljT1G7F8urjfYlq44muV5gDdF3XGxg0eqYiuzBihBDrHPVWDJ/nsM07LYcexP
RTMGVOYelzROPIWrbIGIvPgwDJTaEEuEVd+3S5uZA7vDkb+3xBb/KUtqSH5VLyqV
Wua+YTnof4QLhmqCl3IXwkx2udVT1W9YAtnrutljhsxICiH+oDgiRWReAUtslsUI
Uh3MslQFPqD8UaM7VW3gF6uw2z8AYGO9LNtBFSrwv9q73o6aBMFq9efN5xKEhNwg
EXVXsqRYu7/cq4BtiAKW5UDshfRKA35I1CNBJ7jJ34vjBsCPdkQu2Sk37YY2Vtja
Loi5crsGz7q8eZlaM0A+jV7sK4xw3Xz5KlGnNGmaisdCN65rcM5zhdpkBDmU4rqC
6D3gfUzi6PrWUIrKBGuqEw0eOgABKXrcwm/pzeBludVIuwFcKzjJkAfVDj/ulMDr
Uh7VA4lcuy9Ej6F37VnuYuo9rIAqmLWeZQG5g6VywmqNOKjGDXqnyr9fvgndYmGb
E6X6VSaquouHZBoxrMoGuzu94doUVHjOOxSJGwb70c5ZleikyQM4JGk6J43s/j1w
gkzKwgxDAmtiBwkCNKNDkYeNlQTx+5B/Pmf5Wb35BES3y72VXdPVx4SqWxu9bl6n
YTeYH69qt6zZDsfJeDqbweV2I3MyYRat8VwPLuZ2H88v1XanfCCv1n9jF9kQGDRd
NXX2Hj5F3LNI8d/UddjmQwg2O985o3J63VOcRv8y0SRPZdk/jEkP24d99mssFb9M
fVHQ00OpiMUd87dHhClDq1h2GEgxXVpnRQGUk+QPnjhHgVmVjERs0I9f5RODQ3rk
QHVZ9A/fk+JayuQnrGhkmB/n7K1uS9yV9HCjhRH+5iWNqQ5Ni79sMkXIhQtTb1ut
oUnqxQABtNyq5QxywJrtZETrxZkxq4jgMuAkgpdT0OjLag2mNAvM2xtqsAxm+5Mo
TmW7pmn2jbN1wzMsqq4lZRhIjVkNCzJChPYc8vj6y5IMxpirQaBsVGDvFEzggWB5
XNHtAD9vUv8BqMSNvtwf/zalIbnuFsLFxQ485XOG2lu6zC0O3wH8U6HeZD9PN547
Qqofo9Qfxx4xJeuOh6K88GYbzV9qax4JMdTFd5AJpirPMUIIewOByAmh8Y9Pumd0
Sv8RvMH6VoZftR28Egkq9Gt8nOUU4qiifjW14ahUiAXBQntX6eSQEVW9jVHvKCmh
Y4+a9Ib/cJsaP4j/fVOoxqerJ40QdwR+c6LvXXl+WN27mYhVWcQ1aiGiTMv0oGnt
EL1yWr/MLHUSfvikm9Ko5Q==
`pragma protect end_protected
