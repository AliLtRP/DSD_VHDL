// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lpJu0FJSG17BPDzufBa2AIvoLu6BnoneepUfWE/IFcCrUL8/I0Bc4BotpVVfGeBN
+ucaNor+PnxwgWFW7xnUgUgklMk8RY2xsJTbNTKqW6yrRuIrEF/MWI64FHQS2BPy
vQ+hM23cFbmq9Q51rWtSL77vFbR+uQPtqWP61j3ijdQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4528)
OoBubGOyTPDR6Bd2jiDOize5yyeSUdZKV/ZjOVmH4VfLFryAbSqF38Gy2YQjNGnC
gum/Bx1Lh0evdRsc2UBsX32tgNMGRjvHalXDgsYMCTp3n3xDgQ+QmMFzBh/6hp7Y
n85uHJgQvJH/qmm5z5BMmSK52aiME46wmaVxGyfoTSC8BewjdU6pxsK8B5UFVb6d
upUH7HhJCJb0Ge6SbX4+4sgAWGEvZoj/23cxT9j48q4HcSjhqMHmcyXxC0Mgr0e0
IE2NUQqwB3Hb1HpPWTtraTOEQzLcDjj2pzsHpFuDK3d86gvrwcUOSTP1ZlzFhd9w
vUoxvA86O31vW3izB7HPupHKZubWOpCSq2/DNZmpviDecy+n5RMqTgEHpJ4urmEx
nuXqFdZnBe3Ta8uYI5j1LSPReHuIRIg/9tlUZHEdwO3sMZ5QAAplQbxkICdOsH9Z
sO0lFP/+XfpQYSt2pmZ0fmFAf8/mMFVUXAk1KPrGfVRqsK5QxamUYJt1JaFbg0zv
WU7S5HQnHCC6TO5/lITh7jVZ81eiw1asLQtGFxONB/tpNpQSH7aSIXeoeZ4EWvSJ
Az+byngiFNTe5FIVlYofzzHNm2vPotAQsdWekKjXeHt5EtW9jCePfpHtTYbprOAR
XCk8MQe3XjbTISHe0Q1BtPhOfgo3vHmtYHDUu8oOGsvdqduByRJ8Y8uvkZvQ66/J
kraCqseYIRbg5Jq0SrHSXe5eEYnE7bgIeLSbvBQQLA+Ujlr9jS8mCplkGbnOyuKV
CVzt/EJ9H9bkrzBeXDTtiTirmfXiBhRxp1a0+h78d6LVRYklqIl0biSWcn5d7uEe
ZmNpiqvQHgISVabf44tH/DsqfTg54LBlNYn27RvDnKhxUrdpICiGDMUFOCqG0b+w
QWkWF4URbLYWnYlcNkF5hT9saEGcW+al3zfhgFlpo+tAQIoQFWXxjwRxfpNG8uD6
J60NQblKJprtHWj7w79vwVpwtC/fpuW70D2qEi3r3ROSP5qu6kcNXefyrfLjZWtY
b4e6niCMoDvo0wicjUP6p/Rpj2yIzB6HwOO/tPO3dH75smwN6S/4/0hs3XRF/9hn
2H+AWwy09csu103GjhrNpe32Mpt/jh7Z7KRflXw3COLhoxGbX3SseRSMSsyg/iaG
0nWmJmzySUimTNm1+xTWkO9z2S3Xeg+fhWp7PxrCDnWfjco6dFwK8CzqSlxroJsL
kuKz5oJNdz2F7U9E6bYAzzwWdlSiA8mizsZxoJPcdLwwjjxa2yLLsuUshKe02Q/l
ZqT0F/3zC3lbdTrrZz/jX4doOVv0J7ZdqIIm6UKO9FkJKt8Ko2CZ+PfRaz5IWdSm
Z/7p7ZsM2wysJUIEhviq+pN8xD91uQLF4+rcjOMj5sBY4Guzgt6CMh19K9UDiwrA
VYE6HEhlQLlNBiF+0Vs0VY/GHnQjHI+mtV6X5V2K/ok9q/eJgrbWoILmvWyuMeU6
11OoLrfvY5AvbeKerfWZkKrBaaJdK/3GTX+J5078h8K/OF5XqUtwT9JmgLGoeLva
3b10jrCD2PQ0Jj6oMI2Zb5UAt4fGYTsYNEdINuZT8fAkzS+sIEPahmFqu7vvxgT/
Y7d4Cd/rXaj82Yhwy0lFejRhGca80M+WXNPF8XjvSEs8u4dGSJ4WuX1Dl/WkcWzg
QmiDWm3v6rQ/HwvhAA92AV5TQz45Bj/itfDEHQHG91k1AKc8ZssvTNwHVQkw/N2G
Pdf6T5czdpQPbf88NoWoV2+1CDbLSR49+t/QuKmwNh9iVb/DJb4m15rYiQBo8xgg
BNUvJiwbHPAIfUtBAVy9JGVs2KURnn/6Z8qbbeKKyr9oFljzuGjATme1DUR841zQ
KgdMkUKcYGMKxQDLYZD1bCK3nW51ThigDBqXcWabrEn5PcYpzCPxABwb9b++PzPj
CWoGLFFvrzG/3Hys7x76vnEE9lpcZcVrtwn77CLuyHMuIEXcq2uWWhlGpdfCAp+9
EcFyhrAqos72E0SDC2qvnwM+k5vmUHVCzN3mWxf18ce4a/CY5SFYbfxtt6s6hl+V
gtrm1ECwFMKd6h6MFjK944r5JlOirYkLJADsjGOZ3lqly1uGKyqZFwEghVptGnjJ
2M3TZKFZD5CYUB8lNrIsdl5oIKMh57xYpVhY2gOe+LF/eZdlD+bJ8uA58NYSJrd6
r4bJLWcB1lIH/tM7uJk73Wpr+76hvEDyKjmL5fG5jM5N39oAIvu7TZMneocktykv
UPaN2dcDg85pdGGQcaO7uoVqWkrj2x8Z8VpleZiVF3RKDN81IoprVFIzcwIuthS7
N7djNowzaLtkM55AAMB3yikP7r1Xpsk29KaZzlL+sWedptXOFuT+SJABX6A1xtjx
2qlifSZbPHj+BwWXSWBM+ppMYdhB23ScMIITmP/hqvQIt8vnsECXPli+MafnjNbE
FFmVu6EQSDTkl9/Z04B/gfJJwRI4dA5hR20m0SMk3lJzfRVNra/qlTyZ1nn+0639
3l4Rk/qxcHOH8YzHMa8fCDIvMTJ/RM/V0XHGIoFHIFWyQ785GgHmkKlDuo76J+ak
t3WaH+pq2RPFbd4OLLLMWTiQ3Yi8oXAeIUU8ivv1m76dI5cmhDhrG9Db+ZQ29bcj
LosBabOaA0BYXXOpkdyCdTBXinRDr0I1eixL1lqlkzkQT6MSZIenqzKLcURvOPpV
HqsAKtuvayNvf7bM47wQBPsjiTlo6B768/PqD5GnS0jU70TX5Ssa7I+86jcLGg6C
7LRDvH8qMZHnuqJcbZuAgRnok+gwggeuOzkk/Qz16n+27FpOwWEbicYNAZtjv6xG
HUNwKOpoYsIzAYnrXm8QBeGWxK2iJ8INWUaACg9C+tM1TMHtVuru4sfq4sqzwsG+
TQ4X1wcLXc83dAauBFgfqlFZ/P3md84rPbKFO4RX3hANMYZzxCGxK09wjPynQWHx
fHVwWrDOgY5H+dmpOsr3Z9fi8E+bzMUAzdICCiuVB2gwvC2KHpoVBDc+2nDYunGp
iSI8dPC2QXp+EA5YK2B1tJWSMpx9kEzVCK1NleG+PmcjPIE8sqZnWqn1aMoIEw9t
96AGcyZXjsab8vhOnKQ0lipEgNNfnZya8epvl3NXSgY4OlyJ3o5eReNsuJ5CFPRu
/ynOKeA7B4LVAIeH2gNN54MXSkKYhQ9EuANpaH3r30hy7/kXRKWoFm/dZoTIUQL8
21cWlKIkhG+99yAQlz6owhyN/3OdiuQYxaJ/DJzv6mVWYNqnlwRX6A5xsE3xlZ1V
tr1pdrj6h32b+b0Qyuy5b3XzRfh5zLCVfcJ3eNwkTgBX8zgaf7Dx+GPWdbi2mM2R
GVgW/wQHowQ0wD4fztZa6ZVQS3rqSLE+zqvomTuY5RAhqbjxYwFCfQ3jisAJh7Ad
x/DcNkqIH4SX9LEaBOVJdtnlVR2zmcuiXiLURRA1nYpjkav3PHy9TMSc46J36OSK
bSBvg3PAFae7/tzTaIGD1AJJEGgqpJuzsfVhEy1/Qb24WliaNtIdRx97H3H15EHG
K4aL5OC+7gjgSfWeNqDAQTeRJ4jgFC0+jmRX1TjD9NTPcPlHckSHIiUJUbPufGvu
Fm/x0KTIaQs1V3Kc3TXjV1Wd3s+kSg7FghbgbIPPm+nA/SUF/qn+gP2s/b8NpCPV
GaUbCYwUmL9bWjsuJCa0Kfqw1u6CQxc5li0enfz+LlGXPmgAfMwTZZ2bZLWoSYEr
FsIthxbc/gEZO2y/OqLey1oM9UoyWN6ey0WQGZs1sCMxFnyKdUQJUWb9+NY96d5L
ookewf6oTfOgyQskWir108n3XsWOEGC5i5TTZsnHrmzKSP746NMU0LHE+P6luOKr
cyVe65lYuwgTNZIjrGJGOI7Cfp6vbT0s9+caysxBEezAc7uxokhZ8cPsErCBUXn8
OdRzG9Zl2HrIKEhy6NmUwL29IRCe6KObgn1IOiG2VAtPX4xvrf1np19RIQ/I+Z0i
v44GH66J1UWp79dXdIgkxg3rxCQGWdxsjAM51OD9oT1mYIsAQlQ5uvA+O1HtR0BW
PRhoSnfEujV+WhBehuBCUosklRxBuCZtnar0YEsLfMCl3APAc33BQ3CWl0xjLcxS
p1WymaP4m0v+VkXKMG5U96Dh5Rh1jFMZTsrC+bWN4hB5/G+I2K7OBWbrGqYKrnt9
flyxq2P/gsJebe3TW5iHLhwQarhXKXiPkUPrdfegB8jLzBnQ2rLRg+Qpfuybp5KH
ObpXuOvBUn8cLVTpnLQse+0KeE5Chq+V59p9UgFEHpL7RmvnZYx9ppF2ZvObEJB7
JWJeg8AP+6B6/XgFsHu1c6PqMiMk+a8ch3FMToIwL9hb4Adq+xgWQTWf4cIDYGT1
GUF2JT7IoDx51T5tYa9io3y6YPdZS/It51KoguWYptr9TyxyxFG28ypqmqcSGdXL
r+weFAzCQ7+JthCQ8l1nYUzyPxPaylj0LKEClKxmrhwJfCFpxzxbqIxyUUModc5b
pySk7X4qft0LHzlvOIp9EePH3Ib/Wxj2acBLX+tdBWYgjW8kqh97sz28wAOXuZBr
5IT/LkgjH0jrs+HPkjPX48Z1ONDH/70C83/WsQRLeDlUlrb4ym6YtuuskubY8/Jt
8V4qu/5g6H1F6sP88PXzcAZKVKnV+gZl8HUTnMPxCJSbcdJUMPAnhA2FVgtOqjYW
skGzo02rvbjsq0OuiQnzFnfNHjOxVYkJDtEBa6NA7rNyPWYPIZZFbP9neCHBl7YI
HrWeP7o1P3dVzwcFmfEA5LEWzHS3yw6yJd2sENq+iG65p6lHUOAhGBwGHc2q7vZF
NBtHe5BLJV+thfkQBGWmdbK8prJKCl5oWshzuXaTrsEdMD/CZnOk8eJbWbON6lol
oBHDJm3xR5ng9VJfHurlPDASUOd1yjb6GtSPCgBKt4qMJaT3gzNRE/abJb3yl3FL
QZ0IMASU7ZvK5XQ2Y5QFJyi8xu0QSnwWWT4pD8aHGqVsTlGfwUVQTZXIKsH2AtjI
D3D7Ej8+6nsZ92xDJJHc8V9Zqr7n3aGc3n4wK+cnDpMHqIVGTyE/zCZ+ebi9/rxN
1KnZlM72Lgq9CqPNoAFcvRamrm758nQKx16OWfdCzJYzcORwTUJ7sFchSnjI36GF
cpIzz70zerB8h6WAsNkifIOY3MPTc1X4N5rk+i4ln5g7Vn3Yl0RXvDtQ7G1CpG22
NrRR3MviNf79+LWeTb0S0kPyBWaphBF3Fhha1bfYPpy9Tqz3vHORWNxy0/1P5qZJ
eKfbrMwU6XKODoAP15l48k3KTkoo1388fK9gx0xJwdWKcf5zz0Ncl7StTpUDNNyx
3UXbN9sANe/oqeE2zPRJo4c9KUuJPT83Aqrjy0hLeY5XA+yrC4RWptZ+gWM2IxFV
ELf5a4gt99WijFOjZNtm0xtjaeatIh/gBy4gYMLQXu6viF3zL5+ESirVxX1xcJmG
jWNFukF2UZ8y3V2sjyPKYlSiq7bu7jlX9VFIuQEYwDlNeLqyvmMQUjpIqFy1IBJW
gexrCHbOIGks0uTuePUCNT6Qrlo1pdpkUB7mUSd5+SPVB3ZUN0fX5U9jSHUlFBcH
ul1zuHWWNMkbrSAtNB2UAYus0269q47iBnJqCV/DEmHmE8SuuWnuHUfqp4FFnShh
o6ujpDWBTEUonCdIYX6RxMob6J0DCUEEeNqSnmaBzSw6123oYYgNIKxIWLKTJ4Yk
XBaBZDrlhmQIa/me47pGVzhGRl12EfniSCsbl3FCjSdiR443StfGniw54ux2xbOV
djjibcnkB1jmkAZQoedY6Hfi10jBhjduZA5Fe5jzDn6OOWTpCKZNxLOMk8uiXZkq
mkzsq0g2SwBB77EXi44163V6IFdGntvcBgANdL3olH1pqEN111d66gGQHNvBOQKc
uXeB8a5RvMz41KIgWYXr85gt/mZgRTfjbYsjhh9OhgLuHxwZpuiqeU4DWr1GsBqi
TKIeiDoeJMc4R7d+fzHsPL2Lydb6YxndaYmOQLnRJvY6RDB3MdQj+ifYJYipVuJ7
BacGUntx4QU5S5bA9wsftg==
`pragma protect end_protected
