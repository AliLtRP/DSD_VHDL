-- megafunction wizard: %ALTGX_RECONFIG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt2gxb_reconfig 

-- ============================================================
-- File Name: altgx_reconfig_cpri.vhd
-- Megafunction Name(s):
-- 			alt2gxb_reconfig
--
-- Simulation Library Files(s):
-- 			altera_mf;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.1 Internal Build 112 07/18/2011 PN Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--alt2gxb_reconfig BASE_PORT_WIDTH=1 CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" ENABLE_BUF_CAL="TRUE" ENABLE_CHL_ADDR_FOR_ANALOG_CTRL="TRUE" MIF_ADDRESS_WIDTH=6 NUMBER_OF_CHANNELS=1 NUMBER_OF_RECONFIG_PORTS=1 READ_BASE_PORT_WIDTH=1 RECONFIG_FROMGXB_WIDTH=17 RECONFIG_TOGXB_WIDTH=4 busy channel_reconfig_done reconfig_address_en reconfig_address_out reconfig_clk reconfig_data reconfig_fromgxb reconfig_mode_sel reconfig_togxb write_all
--VERSION_BEGIN 11.1 cbx_alt2gxb_reconfig 2011:07:18:21:10:02:PN cbx_alt_cal 2011:07:18:21:10:02:PN cbx_alt_dprio 2011:07:18:21:10:02:PN cbx_altsyncram 2011:07:18:21:10:02:PN cbx_cycloneii 2011:07:18:21:10:02:PN cbx_lpm_add_sub 2011:07:18:21:10:02:PN cbx_lpm_compare 2011:07:18:21:10:02:PN cbx_lpm_counter 2011:07:18:21:10:02:PN cbx_lpm_decode 2011:07:18:21:10:02:PN cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_lpm_shiftreg 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN cbx_stratix 2011:07:18:21:10:02:PN cbx_stratixii 2011:07:18:21:10:02:PN cbx_stratixiii 2011:07:18:21:10:02:PN cbx_stratixv 2011:07:18:21:10:02:PN cbx_util_mgl 2011:07:18:21:10:02:PN  VERSION_END


--alt_dprio address_width=16 CBX_AUTO_BLACKBOX="ALL" device_family="Stratix IV" quad_address_width=9 address busy datain dataout dpclk dpriodisable dprioin dprioload dprioout quad_address rden reset status_out wren wren_data
--VERSION_BEGIN 11.1 cbx_alt_dprio 2011:07:18:21:10:02:PN cbx_cycloneii 2011:07:18:21:10:02:PN cbx_lpm_add_sub 2011:07:18:21:10:02:PN cbx_lpm_compare 2011:07:18:21:10:02:PN cbx_lpm_counter 2011:07:18:21:10:02:PN cbx_lpm_decode 2011:07:18:21:10:02:PN cbx_lpm_shiftreg 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN cbx_stratix 2011:07:18:21:10:02:PN cbx_stratixii 2011:07:18:21:10:02:PN  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_compare 3 lpm_counter 1 lpm_decode 1 lut 1 reg 102 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_reconfig_cpri_alt_dprio_t2l IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 dpclk	:	IN  STD_LOGIC;
		 dpriodisable	:	OUT  STD_LOGIC;
		 dprioin	:	OUT  STD_LOGIC;
		 dprioload	:	OUT  STD_LOGIC;
		 dprioout	:	IN  STD_LOGIC;
		 quad_address	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 rden	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0';
		 status_out	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 wren	:	IN  STD_LOGIC := '0';
		 wren_data	:	IN  STD_LOGIC := '0'
	 ); 
 END altgx_reconfig_cpri_alt_dprio_t2l;

 ARCHITECTURE RTL OF altgx_reconfig_cpri_alt_dprio_t2l IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to addr_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to wr_out_data_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to rd_out_data_shift_reg[13]} DPRIO_INTERFACE_REG=ON;{-to in_data_shift_reg[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[1]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[2]} DPRIO_INTERFACE_REG=ON";

	 SIGNAL	 wire_addr_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_addr_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 addr_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF addr_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_addr_shift_reg_w_q_range1289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 in_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF in_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rd_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 wire_rd_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 rd_out_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rd_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rd_out_data_shift_reg_w_q_range1465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_startup_cntr_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 startup_cntr	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF startup_cntr : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_startup_cntr_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1530w1533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1534w1540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1534w1543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1526w1527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1526w1542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1526w1531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1534w1535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_state_mc_reg_w_q_range1119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range1138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range1154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wr_out_data_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_wr_out_data_shift_reg_w_q_range1400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb1287w1464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb1287w1399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_agb1287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_agb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rd_data_output_cmpr_ageb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_alb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_state_mc_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_write_state1104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_decode_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	wire_dprioin_mux_dataout	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s0_to_01121w1122w1123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s1_to_01140w1141w1142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s2_to_01156w1157w1158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren1110w1133w1146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren1110w1133w1134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wr_addr_state1286w1290w1291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rd_data_output_state1466w1467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_data_state1401w1402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s0_to_01121w1122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s1_to_01140w1141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s2_to_01156w1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren1110w1133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren1110w1111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren1110w1128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1522w1523w1524w1525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_addr_state1286w1290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rd_data_output_state1466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_data_state1401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_01121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_11120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_01140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_11139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_01156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_11155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_done1520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_idle1521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren1110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren_data1132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_rden1522w1523w1524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden1108w1109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden1522w1523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden1108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden1522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc1145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc1127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_11124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_11143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_11159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_addr_state1286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren1135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren1112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren1149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  rd_addr_done :	STD_LOGIC;
	 SIGNAL  rd_addr_state :	STD_LOGIC;
	 SIGNAL  rd_data_done :	STD_LOGIC;
	 SIGNAL  rd_data_input_state :	STD_LOGIC;
	 SIGNAL  rd_data_output_state :	STD_LOGIC;
	 SIGNAL  rd_data_state :	STD_LOGIC;
	 SIGNAL  rdinc	:	STD_LOGIC;
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s1_to_0 :	STD_LOGIC;
	 SIGNAL  s1_to_1 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  s2_to_1 :	STD_LOGIC;
	 SIGNAL  startup_done :	STD_LOGIC;
	 SIGNAL  startup_idle :	STD_LOGIC;
	 SIGNAL  wr_addr_done :	STD_LOGIC;
	 SIGNAL  wr_addr_state :	STD_LOGIC;
	 SIGNAL  wr_data_done :	STD_LOGIC;
	 SIGNAL  wr_data_state :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_dprio_w_lg_w_lg_w_lg_s0_to_01121w1122w1123w(0) <= wire_dprio_w_lg_w_lg_s0_to_01121w1122w(0) AND wire_state_mc_reg_w_q_range1119w(0);
	wire_dprio_w_lg_w_lg_w_lg_s1_to_01140w1141w1142w(0) <= wire_dprio_w_lg_w_lg_s1_to_01140w1141w(0) AND wire_state_mc_reg_w_q_range1138w(0);
	wire_dprio_w_lg_w_lg_w_lg_s2_to_01156w1157w1158w(0) <= wire_dprio_w_lg_w_lg_s2_to_01156w1157w(0) AND wire_state_mc_reg_w_q_range1154w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren1110w1133w1146w(0) <= wire_dprio_w_lg_w_lg_wren1110w1133w(0) AND wire_dprio_w_lg_rdinc1145w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren1110w1133w1134w(0) <= wire_dprio_w_lg_w_lg_wren1110w1133w(0) AND rden;
	wire_dprio_w_lg_w_lg_w_lg_wr_addr_state1286w1290w1291w(0) <= wire_dprio_w_lg_w_lg_wr_addr_state1286w1290w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_rd_data_output_state1466w1467w(0) <= wire_dprio_w_lg_rd_data_output_state1466w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_wr_data_state1401w1402w(0) <= wire_dprio_w_lg_wr_data_state1401w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_s0_to_01121w1122w(0) <= wire_dprio_w_lg_s0_to_01121w(0) AND wire_dprio_w_lg_s0_to_11120w(0);
	wire_dprio_w_lg_w_lg_s1_to_01140w1141w(0) <= wire_dprio_w_lg_s1_to_01140w(0) AND wire_dprio_w_lg_s1_to_11139w(0);
	wire_dprio_w_lg_w_lg_s2_to_01156w1157w(0) <= wire_dprio_w_lg_s2_to_01156w(0) AND wire_dprio_w_lg_s2_to_11155w(0);
	wire_dprio_w_lg_w_lg_wren1110w1133w(0) <= wire_dprio_w_lg_wren1110w(0) AND wire_dprio_w_lg_wren_data1132w(0);
	wire_dprio_w_lg_w_lg_wren1110w1111w(0) <= wire_dprio_w_lg_wren1110w(0) AND wire_dprio_w_lg_w_lg_rden1108w1109w(0);
	wire_dprio_w_lg_w_lg_wren1110w1128w(0) <= wire_dprio_w_lg_wren1110w(0) AND wire_dprio_w_lg_rdinc1127w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1522w1523w1524w1525w(0) <= wire_dprio_w_lg_w_lg_w_lg_rden1522w1523w1524w(0) AND wire_dprio_w_lg_startup_done1520w(0);
	wire_dprio_w_lg_w_lg_wr_addr_state1286w1290w(0) <= wire_dprio_w_lg_wr_addr_state1286w(0) AND wire_addr_shift_reg_w_q_range1289w(0);
	wire_dprio_w_lg_idle_state1147w(0) <= idle_state AND wire_dprio_w_lg_w_lg_w_lg_wren1110w1133w1146w(0);
	wire_dprio_w_lg_idle_state1129w(0) <= idle_state AND wire_dprio_w_lg_w_lg_wren1110w1128w(0);
	wire_dprio_w_lg_idle_state1136w(0) <= idle_state AND wire_dprio_w_lg_wren1135w(0);
	wire_dprio_w_lg_idle_state1113w(0) <= idle_state AND wire_dprio_w_lg_wren1112w(0);
	wire_dprio_w_lg_idle_state1150w(0) <= idle_state AND wire_dprio_w_lg_wren1149w(0);
	wire_dprio_w_lg_rd_data_output_state1466w(0) <= rd_data_output_state AND wire_rd_out_data_shift_reg_w_q_range1465w(0);
	wire_dprio_w_lg_wr_data_state1401w(0) <= wr_data_state AND wire_wr_out_data_shift_reg_w_q_range1400w(0);
	wire_dprio_w_lg_s0_to_01121w(0) <= NOT s0_to_0;
	wire_dprio_w_lg_s0_to_11120w(0) <= NOT s0_to_1;
	wire_dprio_w_lg_s1_to_01140w(0) <= NOT s1_to_0;
	wire_dprio_w_lg_s1_to_11139w(0) <= NOT s1_to_1;
	wire_dprio_w_lg_s2_to_01156w(0) <= NOT s2_to_0;
	wire_dprio_w_lg_s2_to_11155w(0) <= NOT s2_to_1;
	wire_dprio_w_lg_startup_done1520w(0) <= NOT startup_done;
	wire_dprio_w_lg_startup_idle1521w(0) <= NOT startup_idle;
	wire_dprio_w_lg_wren1110w(0) <= NOT wren;
	wire_dprio_w_lg_wren_data1132w(0) <= NOT wren_data;
	wire_dprio_w_lg_w_lg_w_lg_rden1522w1523w1524w(0) <= wire_dprio_w_lg_w_lg_rden1522w1523w(0) OR wire_dprio_w_lg_startup_idle1521w(0);
	wire_dprio_w_lg_w_lg_rden1108w1109w(0) <= wire_dprio_w_lg_rden1108w(0) OR wren_data;
	wire_dprio_w_lg_w_lg_rden1522w1523w(0) <= wire_dprio_w_lg_rden1522w(0) OR rdinc;
	wire_dprio_w_lg_rden1108w(0) <= rden OR rdinc;
	wire_dprio_w_lg_rden1522w(0) <= rden OR wren;
	wire_dprio_w_lg_rdinc1145w(0) <= rdinc OR rden;
	wire_dprio_w_lg_rdinc1127w(0) <= rdinc OR wren_data;
	wire_dprio_w_lg_s0_to_11124w(0) <= s0_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s0_to_01121w1122w1123w(0);
	wire_dprio_w_lg_s1_to_11143w(0) <= s1_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s1_to_01140w1141w1142w(0);
	wire_dprio_w_lg_s2_to_11159w(0) <= s2_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s2_to_01156w1157w1158w(0);
	wire_dprio_w_lg_wr_addr_state1286w(0) <= wr_addr_state OR rd_addr_state;
	wire_dprio_w_lg_wren1135w(0) <= wren OR wire_dprio_w_lg_w_lg_w_lg_wren1110w1133w1134w(0);
	wire_dprio_w_lg_wren1112w(0) <= wren OR wire_dprio_w_lg_w_lg_wren1110w1111w(0);
	wire_dprio_w_lg_wren1149w(0) <= wren OR wren_data;
	busy <= busy_state;
	busy_state <= (write_state OR read_state);
	dataout <= in_data_shift_reg;
	dpriodisable <= (NOT wire_startup_cntr_w_lg_w_q_range1534w1543w(0));
	dprioin <= wire_dprioin_mux_dataout;
	dprioload <= (NOT (wire_startup_cntr_w_lg_w_q_range1526w1531w(0) AND (NOT startup_cntr(2))));
	idle_state <= wire_state_mc_decode_eq(0);
	rd_addr_done <= (rd_addr_state AND wire_state_mc_cmpr_aeb);
	rd_addr_state <= (wire_state_mc_decode_eq(5) AND startup_done);
	rd_data_done <= (rd_data_state AND wire_state_mc_cmpr_aeb);
	rd_data_input_state <= (wire_rd_data_output_cmpr_ageb AND rd_data_state);
	rd_data_output_state <= (wire_rd_data_output_cmpr_alb AND rd_data_state);
	rd_data_state <= (wire_state_mc_decode_eq(7) AND startup_done);
	rdinc <= '0';
	read_state <= (rd_addr_state OR rd_data_state);
	s0_to_0 <= ((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done));
	s0_to_1 <= ((wire_dprio_w_lg_idle_state1113w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s1_to_0 <= (((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state1136w(0));
	s1_to_1 <= ((wire_dprio_w_lg_idle_state1129w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s2_to_0 <= ((((wr_addr_state AND wr_addr_done) OR (wr_data_state AND wr_data_done)) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state1150w(0));
	s2_to_1 <= (wire_dprio_w_lg_idle_state1147w(0) OR (rd_addr_state AND rd_addr_done));
	startup_done <= (wire_startup_cntr_w_lg_w_q_range1534w1540w(0) AND startup_cntr(1));
	startup_idle <= (wire_startup_cntr_w_lg_w_q_range1526w1527w(0) AND (NOT (startup_cntr(2) XOR startup_cntr(1))));
	status_out <= ( rd_data_done & rd_addr_done & wr_data_done & wr_addr_done);
	wr_addr_done <= (wr_addr_state AND wire_state_mc_cmpr_aeb);
	wr_addr_state <= (wire_state_mc_decode_eq(1) AND startup_done);
	wr_data_done <= (wr_data_state AND wire_state_mc_cmpr_aeb);
	wr_data_state <= (wire_state_mc_decode_eq(3) AND startup_done);
	write_state <= (wr_addr_state OR wr_data_state);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(0) <= wire_addr_shift_reg_asdata(0);
				ELSE addr_shift_reg(0) <= wire_addr_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(1) <= wire_addr_shift_reg_asdata(1);
				ELSE addr_shift_reg(1) <= wire_addr_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(2) <= wire_addr_shift_reg_asdata(2);
				ELSE addr_shift_reg(2) <= wire_addr_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(3) <= wire_addr_shift_reg_asdata(3);
				ELSE addr_shift_reg(3) <= wire_addr_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(4) <= wire_addr_shift_reg_asdata(4);
				ELSE addr_shift_reg(4) <= wire_addr_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(5) <= wire_addr_shift_reg_asdata(5);
				ELSE addr_shift_reg(5) <= wire_addr_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(6) <= wire_addr_shift_reg_asdata(6);
				ELSE addr_shift_reg(6) <= wire_addr_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(7) <= wire_addr_shift_reg_asdata(7);
				ELSE addr_shift_reg(7) <= wire_addr_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(8) <= wire_addr_shift_reg_asdata(8);
				ELSE addr_shift_reg(8) <= wire_addr_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(9) <= wire_addr_shift_reg_asdata(9);
				ELSE addr_shift_reg(9) <= wire_addr_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(10) <= wire_addr_shift_reg_asdata(10);
				ELSE addr_shift_reg(10) <= wire_addr_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(11) <= wire_addr_shift_reg_asdata(11);
				ELSE addr_shift_reg(11) <= wire_addr_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(12) <= wire_addr_shift_reg_asdata(12);
				ELSE addr_shift_reg(12) <= wire_addr_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(13) <= wire_addr_shift_reg_asdata(13);
				ELSE addr_shift_reg(13) <= wire_addr_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(14) <= wire_addr_shift_reg_asdata(14);
				ELSE addr_shift_reg(14) <= wire_addr_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(15) <= wire_addr_shift_reg_asdata(15);
				ELSE addr_shift_reg(15) <= wire_addr_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(16) <= wire_addr_shift_reg_asdata(16);
				ELSE addr_shift_reg(16) <= wire_addr_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(17) <= wire_addr_shift_reg_asdata(17);
				ELSE addr_shift_reg(17) <= wire_addr_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(18) <= wire_addr_shift_reg_asdata(18);
				ELSE addr_shift_reg(18) <= wire_addr_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(19) <= wire_addr_shift_reg_asdata(19);
				ELSE addr_shift_reg(19) <= wire_addr_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(20) <= wire_addr_shift_reg_asdata(20);
				ELSE addr_shift_reg(20) <= wire_addr_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(21) <= wire_addr_shift_reg_asdata(21);
				ELSE addr_shift_reg(21) <= wire_addr_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(22) <= wire_addr_shift_reg_asdata(22);
				ELSE addr_shift_reg(22) <= wire_addr_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(23) <= wire_addr_shift_reg_asdata(23);
				ELSE addr_shift_reg(23) <= wire_addr_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(24) <= wire_addr_shift_reg_asdata(24);
				ELSE addr_shift_reg(24) <= wire_addr_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(25) <= wire_addr_shift_reg_asdata(25);
				ELSE addr_shift_reg(25) <= wire_addr_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(26) <= wire_addr_shift_reg_asdata(26);
				ELSE addr_shift_reg(26) <= wire_addr_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(27) <= wire_addr_shift_reg_asdata(27);
				ELSE addr_shift_reg(27) <= wire_addr_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(28) <= wire_addr_shift_reg_asdata(28);
				ELSE addr_shift_reg(28) <= wire_addr_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(29) <= wire_addr_shift_reg_asdata(29);
				ELSE addr_shift_reg(29) <= wire_addr_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(30) <= wire_addr_shift_reg_asdata(30);
				ELSE addr_shift_reg(30) <= wire_addr_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(31) <= wire_addr_shift_reg_asdata(31);
				ELSE addr_shift_reg(31) <= wire_addr_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_addr_shift_reg_asdata <= ( "00" & "00" & "0" & quad_address(8 DOWNTO 0) & "10" & address);
	wire_addr_shift_reg_d <= ( addr_shift_reg(30 DOWNTO 0) & "0");
	wire_addr_shift_reg_w_q_range1289w(0) <= addr_shift_reg(31);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN in_data_shift_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
			IF (rd_data_input_state = '1') THEN in_data_shift_reg <= ( in_data_shift_reg(14 DOWNTO 0) & dprioout);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_asdata(0);
				ELSE rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_asdata(1);
				ELSE rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_asdata(2);
				ELSE rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_asdata(3);
				ELSE rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_asdata(4);
				ELSE rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_asdata(5);
				ELSE rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_asdata(6);
				ELSE rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_asdata(7);
				ELSE rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_asdata(8);
				ELSE rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_asdata(9);
				ELSE rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_asdata(10);
				ELSE rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_asdata(11);
				ELSE rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_asdata(12);
				ELSE rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_asdata(13);
				ELSE rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_asdata(14);
				ELSE rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_asdata(15);
				ELSE rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	wire_rd_out_data_shift_reg_asdata <= ( "00" & "1" & "1" & "0" & quad_address & "10");
	wire_rd_out_data_shift_reg_d <= ( rd_out_data_shift_reg(14 DOWNTO 0) & "0");
	wire_rd_out_data_shift_reg_w_q_range1465w(0) <= rd_out_data_shift_reg(15);
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(0) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(0) <= '0';
				ELSE startup_cntr(0) <= wire_startup_cntr_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(1) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(1) <= '0';
				ELSE startup_cntr(1) <= wire_startup_cntr_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(2) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(2) <= '0';
				ELSE startup_cntr(2) <= wire_startup_cntr_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_startup_cntr_d <= ( wire_startup_cntr_w_lg_w_q_range1534w1535w & wire_startup_cntr_w_lg_w_q_range1526w1531w & wire_startup_cntr_w_lg_w_q_range1526w1527w);
	loop0 : FOR i IN 0 TO 2 GENERATE
		wire_startup_cntr_ena(i) <= wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1522w1523w1524w1525w(0);
	END GENERATE loop0;
	wire_startup_cntr_w_lg_w_q_range1530w1533w(0) <= wire_startup_cntr_w_q_range1530w(0) AND wire_startup_cntr_w_q_range1526w(0);
	wire_startup_cntr_w_lg_w_q_range1534w1540w(0) <= wire_startup_cntr_w_q_range1534w(0) AND wire_startup_cntr_w_lg_w_q_range1526w1527w(0);
	wire_startup_cntr_w_lg_w_q_range1534w1543w(0) <= wire_startup_cntr_w_q_range1534w(0) AND wire_startup_cntr_w_lg_w_q_range1526w1542w(0);
	wire_startup_cntr_w_lg_w_q_range1526w1527w(0) <= NOT wire_startup_cntr_w_q_range1526w(0);
	wire_startup_cntr_w_lg_w_q_range1526w1542w(0) <= wire_startup_cntr_w_q_range1526w(0) OR wire_startup_cntr_w_q_range1530w(0);
	wire_startup_cntr_w_lg_w_q_range1526w1531w(0) <= wire_startup_cntr_w_q_range1526w(0) XOR wire_startup_cntr_w_q_range1530w(0);
	wire_startup_cntr_w_lg_w_q_range1534w1535w(0) <= wire_startup_cntr_w_q_range1534w(0) XOR wire_startup_cntr_w_lg_w_q_range1530w1533w(0);
	wire_startup_cntr_w_q_range1526w(0) <= startup_cntr(0);
	wire_startup_cntr_w_q_range1530w(0) <= startup_cntr(1);
	wire_startup_cntr_w_q_range1534w(0) <= startup_cntr(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN state_mc_reg <= ( wire_dprio_w_lg_s2_to_11159w & wire_dprio_w_lg_s1_to_11143w & wire_dprio_w_lg_s0_to_11124w);
		END IF;
	END PROCESS;
	wire_state_mc_reg_w_q_range1119w(0) <= state_mc_reg(0);
	wire_state_mc_reg_w_q_range1138w(0) <= state_mc_reg(1);
	wire_state_mc_reg_w_q_range1154w(0) <= state_mc_reg(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_asdata(0);
				ELSE wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_asdata(1);
				ELSE wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_asdata(2);
				ELSE wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_asdata(3);
				ELSE wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_asdata(4);
				ELSE wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_asdata(5);
				ELSE wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_asdata(6);
				ELSE wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_asdata(7);
				ELSE wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_asdata(8);
				ELSE wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_asdata(9);
				ELSE wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_asdata(10);
				ELSE wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_asdata(11);
				ELSE wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_asdata(12);
				ELSE wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_asdata(13);
				ELSE wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_asdata(14);
				ELSE wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_asdata(15);
				ELSE wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_asdata(16);
				ELSE wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_asdata(17);
				ELSE wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_asdata(18);
				ELSE wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_asdata(19);
				ELSE wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_asdata(20);
				ELSE wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_asdata(21);
				ELSE wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_asdata(22);
				ELSE wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_asdata(23);
				ELSE wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_asdata(24);
				ELSE wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_asdata(25);
				ELSE wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_asdata(26);
				ELSE wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_asdata(27);
				ELSE wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_asdata(28);
				ELSE wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_asdata(29);
				ELSE wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_asdata(30);
				ELSE wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_asdata(31);
				ELSE wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_wr_out_data_shift_reg_asdata <= ( "00" & "01" & "0" & quad_address(8 DOWNTO 0) & "10" & datain);
	wire_wr_out_data_shift_reg_d <= ( wr_out_data_shift_reg(30 DOWNTO 0) & "0");
	wire_wr_out_data_shift_reg_w_q_range1400w(0) <= wr_out_data_shift_reg(31);
	wire_pre_amble_cmpr_w_lg_w_lg_agb1287w1464w(0) <= wire_pre_amble_cmpr_w_lg_agb1287w(0) AND rd_data_output_state;
	wire_pre_amble_cmpr_w_lg_w_lg_agb1287w1399w(0) <= wire_pre_amble_cmpr_w_lg_agb1287w(0) AND wr_data_state;
	wire_pre_amble_cmpr_w_lg_agb1287w(0) <= NOT wire_pre_amble_cmpr_agb;
	wire_pre_amble_cmpr_datab <= "011111";
	pre_amble_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_pre_amble_cmpr_aeb,
		agb => wire_pre_amble_cmpr_agb,
		dataa => wire_state_mc_counter_q,
		datab => wire_pre_amble_cmpr_datab
	  );
	wire_rd_data_output_cmpr_datab <= "110000";
	rd_data_output_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		ageb => wire_rd_data_output_cmpr_ageb,
		alb => wire_rd_data_output_cmpr_alb,
		dataa => wire_state_mc_counter_q,
		datab => wire_rd_data_output_cmpr_datab
	  );
	wire_state_mc_cmpr_datab <= (OTHERS => '1');
	state_mc_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_state_mc_cmpr_aeb,
		dataa => wire_state_mc_counter_q,
		datab => wire_state_mc_cmpr_datab
	  );
	wire_state_mc_counter_cnt_en <= wire_dprio_w_lg_write_state1104w(0);
	wire_dprio_w_lg_write_state1104w(0) <= write_state OR read_state;
	state_mc_counter :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => dpclk,
		cnt_en => wire_state_mc_counter_cnt_en,
		q => wire_state_mc_counter_q,
		sclr => reset
	  );
	state_mc_decode :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => state_mc_reg,
		eq => wire_state_mc_decode_eq
	  );
	wire_dprioin_mux_dataout <= (((wire_dprio_w_lg_w_lg_w_lg_wr_addr_state1286w1290w1291w(0) OR (wire_pre_amble_cmpr_w_lg_agb1287w(0) AND wire_dprio_w_lg_wr_addr_state1286w(0))) OR (wire_dprio_w_lg_w_lg_wr_data_state1401w1402w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb1287w1399w(0))) OR (wire_dprio_w_lg_w_lg_rd_data_output_state1466w1467w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb1287w1464w(0))) OR NOT(((write_state OR rd_addr_state) OR rd_data_output_state));

 END RTL; --altgx_reconfig_cpri_alt_dprio_t2l


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=10 LPM_WIDTH=6 LPM_WIDTHS=4 data result sel
--VERSION_BEGIN 11.1 cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN  VERSION_END

--synthesis_resources = lut 30 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_reconfig_cpri_mux_r7a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (59 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altgx_reconfig_cpri_mux_r7a;

 ARCHITECTURE RTL OF altgx_reconfig_cpri_mux_r7a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w5_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w5_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w5_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w2_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w3_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w4_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w5_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (179 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (15 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l3_w5_n1_mux_dataout & wire_l3_w5_n0_mux_dataout & wire_l3_w4_n1_mux_dataout & wire_l3_w4_n0_mux_dataout & wire_l3_w3_n1_mux_dataout & wire_l3_w3_n0_mux_dataout & wire_l3_w2_n1_mux_dataout & wire_l3_w2_n0_mux_dataout & wire_l3_w1_n1_mux_dataout & wire_l3_w1_n0_mux_dataout & wire_l3_w0_n1_mux_dataout & wire_l3_w0_n0_mux_dataout & wire_l2_w5_n3_mux_dataout & wire_l2_w5_n2_mux_dataout & wire_l2_w5_n1_mux_dataout & wire_l2_w5_n0_mux_dataout & wire_l2_w4_n3_mux_dataout & wire_l2_w4_n2_mux_dataout & wire_l2_w4_n1_mux_dataout & wire_l2_w4_n0_mux_dataout & wire_l2_w3_n3_mux_dataout & wire_l2_w3_n2_mux_dataout & wire_l2_w3_n1_mux_dataout & wire_l2_w3_n0_mux_dataout & wire_l2_w2_n3_mux_dataout & wire_l2_w2_n2_mux_dataout & wire_l2_w2_n1_mux_dataout & wire_l2_w2_n0_mux_dataout & wire_l2_w1_n3_mux_dataout & wire_l2_w1_n2_mux_dataout & wire_l2_w1_n1_mux_dataout & wire_l2_w1_n0_mux_dataout & wire_l2_w0_n3_mux_dataout & wire_l2_w0_n2_mux_dataout & wire_l2_w0_n1_mux_dataout & wire_l2_w0_n0_mux_dataout & wire_l1_w5_n7_mux_dataout & wire_l1_w5_n6_mux_dataout & wire_l1_w5_n5_mux_dataout & wire_l1_w5_n4_mux_dataout & wire_l1_w5_n3_mux_dataout & wire_l1_w5_n2_mux_dataout & wire_l1_w5_n1_mux_dataout & wire_l1_w5_n0_mux_dataout & wire_l1_w4_n7_mux_dataout & wire_l1_w4_n6_mux_dataout & wire_l1_w4_n5_mux_dataout & wire_l1_w4_n4_mux_dataout & wire_l1_w4_n3_mux_dataout & wire_l1_w4_n2_mux_dataout & wire_l1_w4_n1_mux_dataout & wire_l1_w4_n0_mux_dataout & wire_l1_w3_n7_mux_dataout & wire_l1_w3_n6_mux_dataout & wire_l1_w3_n5_mux_dataout & wire_l1_w3_n4_mux_dataout & wire_l1_w3_n3_mux_dataout & wire_l1_w3_n2_mux_dataout & wire_l1_w3_n1_mux_dataout & wire_l1_w3_n0_mux_dataout & wire_l1_w2_n7_mux_dataout & wire_l1_w2_n6_mux_dataout & wire_l1_w2_n5_mux_dataout & wire_l1_w2_n4_mux_dataout & wire_l1_w2_n3_mux_dataout & wire_l1_w2_n2_mux_dataout & wire_l1_w2_n1_mux_dataout & wire_l1_w2_n0_mux_dataout & wire_l1_w1_n7_mux_dataout & wire_l1_w1_n6_mux_dataout & wire_l1_w1_n5_mux_dataout & wire_l1_w1_n4_mux_dataout & wire_l1_w1_n3_mux_dataout
 & wire_l1_w1_n2_mux_dataout & wire_l1_w1_n1_mux_dataout & wire_l1_w1_n0_mux_dataout & wire_l1_w0_n7_mux_dataout & wire_l1_w0_n6_mux_dataout & wire_l1_w0_n5_mux_dataout & wire_l1_w0_n4_mux_dataout & wire_l1_w0_n3_mux_dataout & wire_l1_w0_n2_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & "000000000000000000000000000000000000" & data);
	result <= result_wire_ext;
	result_wire_ext <= ( wire_l4_w5_n0_mux_dataout & wire_l4_w4_n0_mux_dataout & wire_l4_w3_n0_mux_dataout & wire_l4_w2_n0_mux_dataout & wire_l4_w1_n0_mux_dataout & wire_l4_w0_n0_mux_dataout);
	sel_wire <= ( sel(3) & "0000" & sel(2) & "0000" & sel(1) & "0000" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(6) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n1_mux_dataout <= data_wire(18) WHEN sel_wire(0) = '1'  ELSE data_wire(12);
	wire_l1_w0_n2_mux_dataout <= data_wire(30) WHEN sel_wire(0) = '1'  ELSE data_wire(24);
	wire_l1_w0_n3_mux_dataout <= data_wire(42) WHEN sel_wire(0) = '1'  ELSE data_wire(36);
	wire_l1_w0_n4_mux_dataout <= data_wire(54) WHEN sel_wire(0) = '1'  ELSE data_wire(48);
	wire_l1_w0_n5_mux_dataout <= data_wire(66) WHEN sel_wire(0) = '1'  ELSE data_wire(60);
	wire_l1_w0_n6_mux_dataout <= data_wire(78) WHEN sel_wire(0) = '1'  ELSE data_wire(72);
	wire_l1_w0_n7_mux_dataout <= data_wire(90) WHEN sel_wire(0) = '1'  ELSE data_wire(84);
	wire_l1_w1_n0_mux_dataout <= data_wire(7) WHEN sel_wire(0) = '1'  ELSE data_wire(1);
	wire_l1_w1_n1_mux_dataout <= data_wire(19) WHEN sel_wire(0) = '1'  ELSE data_wire(13);
	wire_l1_w1_n2_mux_dataout <= data_wire(31) WHEN sel_wire(0) = '1'  ELSE data_wire(25);
	wire_l1_w1_n3_mux_dataout <= data_wire(43) WHEN sel_wire(0) = '1'  ELSE data_wire(37);
	wire_l1_w1_n4_mux_dataout <= data_wire(55) WHEN sel_wire(0) = '1'  ELSE data_wire(49);
	wire_l1_w1_n5_mux_dataout <= data_wire(67) WHEN sel_wire(0) = '1'  ELSE data_wire(61);
	wire_l1_w1_n6_mux_dataout <= data_wire(79) WHEN sel_wire(0) = '1'  ELSE data_wire(73);
	wire_l1_w1_n7_mux_dataout <= data_wire(91) WHEN sel_wire(0) = '1'  ELSE data_wire(85);
	wire_l1_w2_n0_mux_dataout <= data_wire(8) WHEN sel_wire(0) = '1'  ELSE data_wire(2);
	wire_l1_w2_n1_mux_dataout <= data_wire(20) WHEN sel_wire(0) = '1'  ELSE data_wire(14);
	wire_l1_w2_n2_mux_dataout <= data_wire(32) WHEN sel_wire(0) = '1'  ELSE data_wire(26);
	wire_l1_w2_n3_mux_dataout <= data_wire(44) WHEN sel_wire(0) = '1'  ELSE data_wire(38);
	wire_l1_w2_n4_mux_dataout <= data_wire(56) WHEN sel_wire(0) = '1'  ELSE data_wire(50);
	wire_l1_w2_n5_mux_dataout <= data_wire(68) WHEN sel_wire(0) = '1'  ELSE data_wire(62);
	wire_l1_w2_n6_mux_dataout <= data_wire(80) WHEN sel_wire(0) = '1'  ELSE data_wire(74);
	wire_l1_w2_n7_mux_dataout <= data_wire(92) WHEN sel_wire(0) = '1'  ELSE data_wire(86);
	wire_l1_w3_n0_mux_dataout <= data_wire(9) WHEN sel_wire(0) = '1'  ELSE data_wire(3);
	wire_l1_w3_n1_mux_dataout <= data_wire(21) WHEN sel_wire(0) = '1'  ELSE data_wire(15);
	wire_l1_w3_n2_mux_dataout <= data_wire(33) WHEN sel_wire(0) = '1'  ELSE data_wire(27);
	wire_l1_w3_n3_mux_dataout <= data_wire(45) WHEN sel_wire(0) = '1'  ELSE data_wire(39);
	wire_l1_w3_n4_mux_dataout <= data_wire(57) WHEN sel_wire(0) = '1'  ELSE data_wire(51);
	wire_l1_w3_n5_mux_dataout <= data_wire(69) WHEN sel_wire(0) = '1'  ELSE data_wire(63);
	wire_l1_w3_n6_mux_dataout <= data_wire(81) WHEN sel_wire(0) = '1'  ELSE data_wire(75);
	wire_l1_w3_n7_mux_dataout <= data_wire(93) WHEN sel_wire(0) = '1'  ELSE data_wire(87);
	wire_l1_w4_n0_mux_dataout <= data_wire(10) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w4_n1_mux_dataout <= data_wire(22) WHEN sel_wire(0) = '1'  ELSE data_wire(16);
	wire_l1_w4_n2_mux_dataout <= data_wire(34) WHEN sel_wire(0) = '1'  ELSE data_wire(28);
	wire_l1_w4_n3_mux_dataout <= data_wire(46) WHEN sel_wire(0) = '1'  ELSE data_wire(40);
	wire_l1_w4_n4_mux_dataout <= data_wire(58) WHEN sel_wire(0) = '1'  ELSE data_wire(52);
	wire_l1_w4_n5_mux_dataout <= data_wire(70) WHEN sel_wire(0) = '1'  ELSE data_wire(64);
	wire_l1_w4_n6_mux_dataout <= data_wire(82) WHEN sel_wire(0) = '1'  ELSE data_wire(76);
	wire_l1_w4_n7_mux_dataout <= data_wire(94) WHEN sel_wire(0) = '1'  ELSE data_wire(88);
	wire_l1_w5_n0_mux_dataout <= data_wire(11) WHEN sel_wire(0) = '1'  ELSE data_wire(5);
	wire_l1_w5_n1_mux_dataout <= data_wire(23) WHEN sel_wire(0) = '1'  ELSE data_wire(17);
	wire_l1_w5_n2_mux_dataout <= data_wire(35) WHEN sel_wire(0) = '1'  ELSE data_wire(29);
	wire_l1_w5_n3_mux_dataout <= data_wire(47) WHEN sel_wire(0) = '1'  ELSE data_wire(41);
	wire_l1_w5_n4_mux_dataout <= data_wire(59) WHEN sel_wire(0) = '1'  ELSE data_wire(53);
	wire_l1_w5_n5_mux_dataout <= data_wire(71) WHEN sel_wire(0) = '1'  ELSE data_wire(65);
	wire_l1_w5_n6_mux_dataout <= data_wire(83) WHEN sel_wire(0) = '1'  ELSE data_wire(77);
	wire_l1_w5_n7_mux_dataout <= data_wire(95) WHEN sel_wire(0) = '1'  ELSE data_wire(89);
	wire_l2_w0_n0_mux_dataout <= data_wire(97) WHEN sel_wire(5) = '1'  ELSE data_wire(96);
	wire_l2_w0_n1_mux_dataout <= data_wire(99) WHEN sel_wire(5) = '1'  ELSE data_wire(98);
	wire_l2_w0_n2_mux_dataout <= data_wire(101) WHEN sel_wire(5) = '1'  ELSE data_wire(100);
	wire_l2_w0_n3_mux_dataout <= data_wire(103) WHEN sel_wire(5) = '1'  ELSE data_wire(102);
	wire_l2_w1_n0_mux_dataout <= data_wire(105) WHEN sel_wire(5) = '1'  ELSE data_wire(104);
	wire_l2_w1_n1_mux_dataout <= data_wire(107) WHEN sel_wire(5) = '1'  ELSE data_wire(106);
	wire_l2_w1_n2_mux_dataout <= data_wire(109) WHEN sel_wire(5) = '1'  ELSE data_wire(108);
	wire_l2_w1_n3_mux_dataout <= data_wire(111) WHEN sel_wire(5) = '1'  ELSE data_wire(110);
	wire_l2_w2_n0_mux_dataout <= data_wire(113) WHEN sel_wire(5) = '1'  ELSE data_wire(112);
	wire_l2_w2_n1_mux_dataout <= data_wire(115) WHEN sel_wire(5) = '1'  ELSE data_wire(114);
	wire_l2_w2_n2_mux_dataout <= data_wire(117) WHEN sel_wire(5) = '1'  ELSE data_wire(116);
	wire_l2_w2_n3_mux_dataout <= data_wire(119) WHEN sel_wire(5) = '1'  ELSE data_wire(118);
	wire_l2_w3_n0_mux_dataout <= data_wire(121) WHEN sel_wire(5) = '1'  ELSE data_wire(120);
	wire_l2_w3_n1_mux_dataout <= data_wire(123) WHEN sel_wire(5) = '1'  ELSE data_wire(122);
	wire_l2_w3_n2_mux_dataout <= data_wire(125) WHEN sel_wire(5) = '1'  ELSE data_wire(124);
	wire_l2_w3_n3_mux_dataout <= data_wire(127) WHEN sel_wire(5) = '1'  ELSE data_wire(126);
	wire_l2_w4_n0_mux_dataout <= data_wire(129) WHEN sel_wire(5) = '1'  ELSE data_wire(128);
	wire_l2_w4_n1_mux_dataout <= data_wire(131) WHEN sel_wire(5) = '1'  ELSE data_wire(130);
	wire_l2_w4_n2_mux_dataout <= data_wire(133) WHEN sel_wire(5) = '1'  ELSE data_wire(132);
	wire_l2_w4_n3_mux_dataout <= data_wire(135) WHEN sel_wire(5) = '1'  ELSE data_wire(134);
	wire_l2_w5_n0_mux_dataout <= data_wire(137) WHEN sel_wire(5) = '1'  ELSE data_wire(136);
	wire_l2_w5_n1_mux_dataout <= data_wire(139) WHEN sel_wire(5) = '1'  ELSE data_wire(138);
	wire_l2_w5_n2_mux_dataout <= data_wire(141) WHEN sel_wire(5) = '1'  ELSE data_wire(140);
	wire_l2_w5_n3_mux_dataout <= data_wire(143) WHEN sel_wire(5) = '1'  ELSE data_wire(142);
	wire_l3_w0_n0_mux_dataout <= data_wire(145) WHEN sel_wire(10) = '1'  ELSE data_wire(144);
	wire_l3_w0_n1_mux_dataout <= data_wire(147) WHEN sel_wire(10) = '1'  ELSE data_wire(146);
	wire_l3_w1_n0_mux_dataout <= data_wire(149) WHEN sel_wire(10) = '1'  ELSE data_wire(148);
	wire_l3_w1_n1_mux_dataout <= data_wire(151) WHEN sel_wire(10) = '1'  ELSE data_wire(150);
	wire_l3_w2_n0_mux_dataout <= data_wire(153) WHEN sel_wire(10) = '1'  ELSE data_wire(152);
	wire_l3_w2_n1_mux_dataout <= data_wire(155) WHEN sel_wire(10) = '1'  ELSE data_wire(154);
	wire_l3_w3_n0_mux_dataout <= data_wire(157) WHEN sel_wire(10) = '1'  ELSE data_wire(156);
	wire_l3_w3_n1_mux_dataout <= data_wire(159) WHEN sel_wire(10) = '1'  ELSE data_wire(158);
	wire_l3_w4_n0_mux_dataout <= data_wire(161) WHEN sel_wire(10) = '1'  ELSE data_wire(160);
	wire_l3_w4_n1_mux_dataout <= data_wire(163) WHEN sel_wire(10) = '1'  ELSE data_wire(162);
	wire_l3_w5_n0_mux_dataout <= data_wire(165) WHEN sel_wire(10) = '1'  ELSE data_wire(164);
	wire_l3_w5_n1_mux_dataout <= data_wire(167) WHEN sel_wire(10) = '1'  ELSE data_wire(166);
	wire_l4_w0_n0_mux_dataout <= data_wire(169) WHEN sel_wire(15) = '1'  ELSE data_wire(168);
	wire_l4_w1_n0_mux_dataout <= data_wire(171) WHEN sel_wire(15) = '1'  ELSE data_wire(170);
	wire_l4_w2_n0_mux_dataout <= data_wire(173) WHEN sel_wire(15) = '1'  ELSE data_wire(172);
	wire_l4_w3_n0_mux_dataout <= data_wire(175) WHEN sel_wire(15) = '1'  ELSE data_wire(174);
	wire_l4_w4_n0_mux_dataout <= data_wire(177) WHEN sel_wire(15) = '1'  ELSE data_wire(176);
	wire_l4_w5_n0_mux_dataout <= data_wire(179) WHEN sel_wire(15) = '1'  ELSE data_wire(178);

 END RTL; --altgx_reconfig_cpri_mux_r7a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=3 LPM_WIDTH=5 LPM_WIDTHS=2 data result sel
--VERSION_BEGIN 11.1 cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN  VERSION_END

--synthesis_resources = lut 10 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_reconfig_cpri_mux_a6a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (14 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altgx_reconfig_cpri_mux_a6a;

 ARCHITECTURE RTL OF altgx_reconfig_cpri_mux_a6a IS

	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_lg_w_lg_data0_wire1758w1759w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1755w1756w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1750w1751w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1752w1753w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_lg_w_sel_range1748w1749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_lg_w_sel_range1754w1757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_lg_data0_wire1758w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  data0_wire :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  data1_wire :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  data2_wire :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  result_node :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_data_range1755w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_data_range1750w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_data_range1752w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_sel_range1748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_w_sel_range1754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	loop1 : FOR i IN 0 TO 4 GENERATE 
		wire_central_pcs_global_clk_div_mux_w_lg_w_lg_data0_wire1758w1759w(i) <= wire_central_pcs_global_clk_div_mux_w_lg_data0_wire1758w(i) AND wire_central_pcs_global_clk_div_mux_w_lg_w_sel_range1754w1757w(0);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 4 GENERATE 
		wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1755w1756w(i) <= wire_central_pcs_global_clk_div_mux_w_data_range1755w(i) AND wire_central_pcs_global_clk_div_mux_w_sel_range1754w(0);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 4 GENERATE 
		wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1750w1751w(i) <= wire_central_pcs_global_clk_div_mux_w_data_range1750w(i) AND wire_central_pcs_global_clk_div_mux_w_lg_w_sel_range1748w1749w(0);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 4 GENERATE 
		wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1752w1753w(i) <= wire_central_pcs_global_clk_div_mux_w_data_range1752w(i) AND wire_central_pcs_global_clk_div_mux_w_sel_range1748w(0);
	END GENERATE loop4;
	wire_central_pcs_global_clk_div_mux_w_lg_w_sel_range1748w1749w(0) <= NOT wire_central_pcs_global_clk_div_mux_w_sel_range1748w(0);
	wire_central_pcs_global_clk_div_mux_w_lg_w_sel_range1754w1757w(0) <= NOT wire_central_pcs_global_clk_div_mux_w_sel_range1754w(0);
	loop5 : FOR i IN 0 TO 4 GENERATE 
		wire_central_pcs_global_clk_div_mux_w_lg_data0_wire1758w(i) <= data0_wire(i) OR data1_wire(i);
	END GENERATE loop5;
	data0_wire <= wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1750w1751w;
	data1_wire <= wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1752w1753w;
	data2_wire <= wire_central_pcs_global_clk_div_mux_w_lg_w_data_range1755w1756w;
	result <= result_node;
	result_node <= (wire_central_pcs_global_clk_div_mux_w_lg_w_lg_data0_wire1758w1759w OR data2_wire);
	wire_central_pcs_global_clk_div_mux_w_data_range1755w <= data(14 DOWNTO 10);
	wire_central_pcs_global_clk_div_mux_w_data_range1750w <= data(4 DOWNTO 0);
	wire_central_pcs_global_clk_div_mux_w_data_range1752w <= data(9 DOWNTO 5);
	wire_central_pcs_global_clk_div_mux_w_sel_range1748w(0) <= sel(0);
	wire_central_pcs_global_clk_div_mux_w_sel_range1754w(0) <= sel(1);

 END RTL; --altgx_reconfig_cpri_mux_a6a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=5 LPM_WIDTH=5 LPM_WIDTHS=3 data result sel
--VERSION_BEGIN 11.1 cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN  VERSION_END

--synthesis_resources = lut 12 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_reconfig_cpri_mux_d6a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (24 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altgx_reconfig_cpri_mux_d6a;

 ARCHITECTURE RTL OF altgx_reconfig_cpri_mux_d6a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (8 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l2_w4_n1_mux_dataout & wire_l2_w4_n0_mux_dataout & wire_l2_w3_n1_mux_dataout & wire_l2_w3_n0_mux_dataout & wire_l2_w2_n1_mux_dataout & wire_l2_w2_n0_mux_dataout & wire_l2_w1_n1_mux_dataout & wire_l2_w1_n0_mux_dataout & wire_l2_w0_n1_mux_dataout & wire_l2_w0_n0_mux_dataout & wire_l1_w4_n3_mux_dataout & wire_l1_w4_n2_mux_dataout & wire_l1_w4_n1_mux_dataout & wire_l1_w4_n0_mux_dataout & wire_l1_w3_n3_mux_dataout & wire_l1_w3_n2_mux_dataout & wire_l1_w3_n1_mux_dataout & wire_l1_w3_n0_mux_dataout & wire_l1_w2_n3_mux_dataout & wire_l1_w2_n2_mux_dataout & wire_l1_w2_n1_mux_dataout & wire_l1_w2_n0_mux_dataout & wire_l1_w1_n3_mux_dataout & wire_l1_w1_n2_mux_dataout & wire_l1_w1_n1_mux_dataout & wire_l1_w1_n0_mux_dataout & wire_l1_w0_n3_mux_dataout & wire_l1_w0_n2_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & "000000000000000" & data);
	result <= result_wire_ext;
	result_wire_ext <= ( wire_l3_w4_n0_mux_dataout & wire_l3_w3_n0_mux_dataout & wire_l3_w2_n0_mux_dataout & wire_l3_w1_n0_mux_dataout & wire_l3_w0_n0_mux_dataout);
	sel_wire <= ( sel(2) & "000" & sel(1) & "000" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(5) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n1_mux_dataout <= data_wire(15) WHEN sel_wire(0) = '1'  ELSE data_wire(10);
	wire_l1_w0_n2_mux_dataout <= data_wire(25) WHEN sel_wire(0) = '1'  ELSE data_wire(20);
	wire_l1_w0_n3_mux_dataout <= data_wire(35) WHEN sel_wire(0) = '1'  ELSE data_wire(30);
	wire_l1_w1_n0_mux_dataout <= data_wire(6) WHEN sel_wire(0) = '1'  ELSE data_wire(1);
	wire_l1_w1_n1_mux_dataout <= data_wire(16) WHEN sel_wire(0) = '1'  ELSE data_wire(11);
	wire_l1_w1_n2_mux_dataout <= data_wire(26) WHEN sel_wire(0) = '1'  ELSE data_wire(21);
	wire_l1_w1_n3_mux_dataout <= data_wire(36) WHEN sel_wire(0) = '1'  ELSE data_wire(31);
	wire_l1_w2_n0_mux_dataout <= data_wire(7) WHEN sel_wire(0) = '1'  ELSE data_wire(2);
	wire_l1_w2_n1_mux_dataout <= data_wire(17) WHEN sel_wire(0) = '1'  ELSE data_wire(12);
	wire_l1_w2_n2_mux_dataout <= data_wire(27) WHEN sel_wire(0) = '1'  ELSE data_wire(22);
	wire_l1_w2_n3_mux_dataout <= data_wire(37) WHEN sel_wire(0) = '1'  ELSE data_wire(32);
	wire_l1_w3_n0_mux_dataout <= data_wire(8) WHEN sel_wire(0) = '1'  ELSE data_wire(3);
	wire_l1_w3_n1_mux_dataout <= data_wire(18) WHEN sel_wire(0) = '1'  ELSE data_wire(13);
	wire_l1_w3_n2_mux_dataout <= data_wire(28) WHEN sel_wire(0) = '1'  ELSE data_wire(23);
	wire_l1_w3_n3_mux_dataout <= data_wire(38) WHEN sel_wire(0) = '1'  ELSE data_wire(33);
	wire_l1_w4_n0_mux_dataout <= data_wire(9) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w4_n1_mux_dataout <= data_wire(19) WHEN sel_wire(0) = '1'  ELSE data_wire(14);
	wire_l1_w4_n2_mux_dataout <= data_wire(29) WHEN sel_wire(0) = '1'  ELSE data_wire(24);
	wire_l1_w4_n3_mux_dataout <= data_wire(39) WHEN sel_wire(0) = '1'  ELSE data_wire(34);
	wire_l2_w0_n0_mux_dataout <= data_wire(41) WHEN sel_wire(4) = '1'  ELSE data_wire(40);
	wire_l2_w0_n1_mux_dataout <= data_wire(43) WHEN sel_wire(4) = '1'  ELSE data_wire(42);
	wire_l2_w1_n0_mux_dataout <= data_wire(45) WHEN sel_wire(4) = '1'  ELSE data_wire(44);
	wire_l2_w1_n1_mux_dataout <= data_wire(47) WHEN sel_wire(4) = '1'  ELSE data_wire(46);
	wire_l2_w2_n0_mux_dataout <= data_wire(49) WHEN sel_wire(4) = '1'  ELSE data_wire(48);
	wire_l2_w2_n1_mux_dataout <= data_wire(51) WHEN sel_wire(4) = '1'  ELSE data_wire(50);
	wire_l2_w3_n0_mux_dataout <= data_wire(53) WHEN sel_wire(4) = '1'  ELSE data_wire(52);
	wire_l2_w3_n1_mux_dataout <= data_wire(55) WHEN sel_wire(4) = '1'  ELSE data_wire(54);
	wire_l2_w4_n0_mux_dataout <= data_wire(57) WHEN sel_wire(4) = '1'  ELSE data_wire(56);
	wire_l2_w4_n1_mux_dataout <= data_wire(59) WHEN sel_wire(4) = '1'  ELSE data_wire(58);
	wire_l3_w0_n0_mux_dataout <= data_wire(61) WHEN sel_wire(8) = '1'  ELSE data_wire(60);
	wire_l3_w1_n0_mux_dataout <= data_wire(63) WHEN sel_wire(8) = '1'  ELSE data_wire(62);
	wire_l3_w2_n0_mux_dataout <= data_wire(65) WHEN sel_wire(8) = '1'  ELSE data_wire(64);
	wire_l3_w3_n0_mux_dataout <= data_wire(67) WHEN sel_wire(8) = '1'  ELSE data_wire(66);
	wire_l3_w4_n0_mux_dataout <= data_wire(69) WHEN sel_wire(8) = '1'  ELSE data_wire(68);

 END RTL; --altgx_reconfig_cpri_mux_d6a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=3 LPM_WIDTH=6 LPM_WIDTHS=2 data result sel
--VERSION_BEGIN 11.1 cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN  VERSION_END

--synthesis_resources = lut 12 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_reconfig_cpri_mux_b6a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (17 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altgx_reconfig_cpri_mux_b6a;

 ARCHITECTURE RTL OF altgx_reconfig_cpri_mux_b6a IS

	 SIGNAL  wire_mif_addr_cntr_data_mux_w_lg_w_lg_data0_wire1858w1859w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_lg_w_data_range1852w1853w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_lg_w_data_range1855w1856w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_lg_w_data_range1850w1851w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_lg_w_sel_range1848w1849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_lg_w_sel_range1854w1857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_lg_data0_wire1858w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  data0_wire :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  data1_wire :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  data2_wire :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  result_node :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_data_range1852w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_data_range1855w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_data_range1850w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_sel_range1848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_w_sel_range1854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	loop6 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_data_mux_w_lg_w_lg_data0_wire1858w1859w(i) <= wire_mif_addr_cntr_data_mux_w_lg_data0_wire1858w(i) AND wire_mif_addr_cntr_data_mux_w_lg_w_sel_range1854w1857w(0);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_data_mux_w_lg_w_data_range1852w1853w(i) <= wire_mif_addr_cntr_data_mux_w_data_range1852w(i) AND wire_mif_addr_cntr_data_mux_w_sel_range1848w(0);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_data_mux_w_lg_w_data_range1855w1856w(i) <= wire_mif_addr_cntr_data_mux_w_data_range1855w(i) AND wire_mif_addr_cntr_data_mux_w_sel_range1854w(0);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_data_mux_w_lg_w_data_range1850w1851w(i) <= wire_mif_addr_cntr_data_mux_w_data_range1850w(i) AND wire_mif_addr_cntr_data_mux_w_lg_w_sel_range1848w1849w(0);
	END GENERATE loop9;
	wire_mif_addr_cntr_data_mux_w_lg_w_sel_range1848w1849w(0) <= NOT wire_mif_addr_cntr_data_mux_w_sel_range1848w(0);
	wire_mif_addr_cntr_data_mux_w_lg_w_sel_range1854w1857w(0) <= NOT wire_mif_addr_cntr_data_mux_w_sel_range1854w(0);
	loop10 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_data_mux_w_lg_data0_wire1858w(i) <= data0_wire(i) OR data1_wire(i);
	END GENERATE loop10;
	data0_wire <= wire_mif_addr_cntr_data_mux_w_lg_w_data_range1850w1851w;
	data1_wire <= wire_mif_addr_cntr_data_mux_w_lg_w_data_range1852w1853w;
	data2_wire <= wire_mif_addr_cntr_data_mux_w_lg_w_data_range1855w1856w;
	result <= result_node;
	result_node <= (wire_mif_addr_cntr_data_mux_w_lg_w_lg_data0_wire1858w1859w OR data2_wire);
	wire_mif_addr_cntr_data_mux_w_data_range1852w <= data(11 DOWNTO 6);
	wire_mif_addr_cntr_data_mux_w_data_range1855w <= data(17 DOWNTO 12);
	wire_mif_addr_cntr_data_mux_w_data_range1850w <= data(5 DOWNTO 0);
	wire_mif_addr_cntr_data_mux_w_sel_range1848w(0) <= sel(0);
	wire_mif_addr_cntr_data_mux_w_sel_range1854w(0) <= sel(1);

 END RTL; --altgx_reconfig_cpri_mux_b6a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=4 LPM_WIDTH=6 LPM_WIDTHS=2 data result sel
--VERSION_BEGIN 11.1 cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN  VERSION_END

--synthesis_resources = lut 6 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_reconfig_cpri_mux_c6a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altgx_reconfig_cpri_mux_c6a;

 ARCHITECTURE RTL OF altgx_reconfig_cpri_mux_c6a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l1_w5_n1_mux_dataout & wire_l1_w5_n0_mux_dataout & wire_l1_w4_n1_mux_dataout & wire_l1_w4_n0_mux_dataout & wire_l1_w3_n1_mux_dataout & wire_l1_w3_n0_mux_dataout & wire_l1_w2_n1_mux_dataout & wire_l1_w2_n0_mux_dataout & wire_l1_w1_n1_mux_dataout & wire_l1_w1_n0_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & data);
	result <= result_wire_ext;
	result_wire_ext <= ( wire_l2_w5_n0_mux_dataout & wire_l2_w4_n0_mux_dataout & wire_l2_w3_n0_mux_dataout & wire_l2_w2_n0_mux_dataout & wire_l2_w1_n0_mux_dataout & wire_l2_w0_n0_mux_dataout);
	sel_wire <= ( sel(1) & "00" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(6) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n1_mux_dataout <= data_wire(18) WHEN sel_wire(0) = '1'  ELSE data_wire(12);
	wire_l1_w1_n0_mux_dataout <= data_wire(7) WHEN sel_wire(0) = '1'  ELSE data_wire(1);
	wire_l1_w1_n1_mux_dataout <= data_wire(19) WHEN sel_wire(0) = '1'  ELSE data_wire(13);
	wire_l1_w2_n0_mux_dataout <= data_wire(8) WHEN sel_wire(0) = '1'  ELSE data_wire(2);
	wire_l1_w2_n1_mux_dataout <= data_wire(20) WHEN sel_wire(0) = '1'  ELSE data_wire(14);
	wire_l1_w3_n0_mux_dataout <= data_wire(9) WHEN sel_wire(0) = '1'  ELSE data_wire(3);
	wire_l1_w3_n1_mux_dataout <= data_wire(21) WHEN sel_wire(0) = '1'  ELSE data_wire(15);
	wire_l1_w4_n0_mux_dataout <= data_wire(10) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w4_n1_mux_dataout <= data_wire(22) WHEN sel_wire(0) = '1'  ELSE data_wire(16);
	wire_l1_w5_n0_mux_dataout <= data_wire(11) WHEN sel_wire(0) = '1'  ELSE data_wire(5);
	wire_l1_w5_n1_mux_dataout <= data_wire(23) WHEN sel_wire(0) = '1'  ELSE data_wire(17);
	wire_l2_w0_n0_mux_dataout <= data_wire(25) WHEN sel_wire(3) = '1'  ELSE data_wire(24);
	wire_l2_w1_n0_mux_dataout <= data_wire(27) WHEN sel_wire(3) = '1'  ELSE data_wire(26);
	wire_l2_w2_n0_mux_dataout <= data_wire(29) WHEN sel_wire(3) = '1'  ELSE data_wire(28);
	wire_l2_w3_n0_mux_dataout <= data_wire(31) WHEN sel_wire(3) = '1'  ELSE data_wire(30);
	wire_l2_w4_n0_mux_dataout <= data_wire(33) WHEN sel_wire(3) = '1'  ELSE data_wire(32);
	wire_l2_w5_n0_mux_dataout <= data_wire(35) WHEN sel_wire(3) = '1'  ELSE data_wire(34);

 END RTL; --altgx_reconfig_cpri_mux_c6a

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = alt_cal 1 lpm_add_sub 2 lpm_compare 23 lpm_counter 3 lpm_decode 2 lut 72 reg 179 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_reconfig_cpri_alt2gxb_reconfig_7ba1 IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 channel_reconfig_done	:	OUT  STD_LOGIC;
		 reconfig_address_en	:	OUT  STD_LOGIC;
		 reconfig_address_out	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 reconfig_clk	:	IN  STD_LOGIC;
		 reconfig_data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 reconfig_fromgxb	:	IN  STD_LOGIC_VECTOR (16 DOWNTO 0);
		 reconfig_mode_sel	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 reconfig_togxb	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 write_all	:	IN  STD_LOGIC := '0'
	 ); 
 END altgx_reconfig_cpri_alt2gxb_reconfig_7ba1;

 ARCHITECTURE RTL OF altgx_reconfig_cpri_alt2gxb_reconfig_7ba1 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to address_pres_reg[11]} DPRIO_CHANNEL_NUM=11;{-to address_pres_reg[10]} DPRIO_CHANNEL_NUM=10;{-to address_pres_reg[9]} DPRIO_CHANNEL_NUM=9;{-to address_pres_reg[8]} DPRIO_CHANNEL_NUM=8;{-to address_pres_reg[7]} DPRIO_CHANNEL_NUM=7;{-to address_pres_reg[6]} DPRIO_CHANNEL_NUM=6;{-to address_pres_reg[5]} DPRIO_CHANNEL_NUM=5;{-to address_pres_reg[4]} DPRIO_CHANNEL_NUM=4;{-to address_pres_reg[3]} DPRIO_CHANNEL_NUM=3;{-to address_pres_reg[2]} DPRIO_CHANNEL_NUM=2;{-to address_pres_reg[1]} DPRIO_CHANNEL_NUM=1;{-to address_pres_reg[0]} DPRIO_CHANNEL_NUM=0;{-to cru_num_reg[3]} DPRIO_CRUCLK_NUM=3;{-to cru_num_reg[2]} DPRIO_CRUCLK_NUM=2;{-to cru_num_reg[1]} DPRIO_CRUCLK_NUM=1;{-to cru_num_reg[0]} DPRIO_CRUCLK_NUM=0;{-to tx_pll_inclk_reg[3]} DPRIO_TX_PLL0_REFCLK_NUM=3;{-to tx_pll_inclk_reg[2]} DPRIO_TX_PLL0_REFCLK_NUM=2;{-to tx_pll_inclk_reg[1]} DPRIO_TX_PLL0_REFCLK_NUM=1;{-to tx_pll_inclk_reg[0]} DPRIO_TX_PLL0_REFCLK_NUM=0;{-to tx_cmu_sel[2]}  DPRIO_TX_PLL_NUM=2;{-to tx_cmu_sel[1]}  DPRIO_TX_PLL_NUM=1;{-to le7} IMPLEMENT_AS_CLOCK_ENABLE = ON;{-to tx_cmu_sel[0]}  DPRIO_TX_PLL_NUM=0";

	 SIGNAL  wire_calibration_w_lg_w_lg_busy138w142w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy138w139w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy138w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy138w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy138w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy143w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy140w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_busy	:	STD_LOGIC;
	 SIGNAL  wire_calibration_dprio_addr	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_quad_addr	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_calibration_reset	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_offset_cancellation_reset123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_retain_addr	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_status_out_range691w729w730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_busy170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_status_out_range691w729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_address	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy143w144w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_busy	:	STD_LOGIC;
	 SIGNAL  wire_dprio_datain	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy140w141w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dpriodisable	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioin	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioload	:	STD_LOGIC;
	 SIGNAL  wire_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy146w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_status_out	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy149w150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_wren_data	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy152w153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_status_out_range691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_status_out_range728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 address_pres_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF address_pres_reg : SIGNAL IS "PRESERVE_REGISTER=ON";

	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_q_range107w108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range111w112w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range107w108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range107w108w109w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range111w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 cru_num_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF cru_num_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range309w323w324w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_q_range306w307w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_q_range306w307w308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_q_range305w311w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_q_range305w311w340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_q_range309w323w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_q_range306w307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_q_range304w310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_q_range305w311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_q_range306w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_q_range309w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_lg_w_lg_w_q_range309w323w324w325w326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range305w311w312w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range305w311w340w341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_lg_w_lg_w_q_range305w311w312w313w314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_lg_w_q_range309w333w334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_lg_w_q_range309w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_q_range304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_q_range305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_q_range306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cru_num_reg_w_q_range309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 delay_mif_head	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF delay_mif_head : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_delay_mif_head_ena	:	STD_LOGIC;
	 SIGNAL	 delay_second_mif_head	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF delay_second_mif_head : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_delay_second_mif_head_ena	:	STD_LOGIC;
	 SIGNAL	 wire_dprio_dataout_reg_d	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 dprio_dataout_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF dprio_dataout_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_dprio_dataout_reg_ena	:	STD_LOGIC_VECTOR(15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range457w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range489w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range345w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range384w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range476w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range449w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range465w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range482w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range492w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range510w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range403w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range590w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range353w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range501w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range527w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dprio_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF dprio_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_dprio_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_mif_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF end_mif_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 global_register_reset_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF global_register_reset_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 is_bonded_global_clk_div_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF is_bonded_global_clk_div_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_is_bonded_global_clk_div_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_is_bonded_global_clk_div_reg_w_lg_w_lg_q812w813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_is_bonded_global_clk_div_reg_w_lg_w_lg_w_lg_w_lg_q812w813w814w815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_is_bonded_global_clk_div_reg_w_lg_q812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_is_bonded_global_clk_div_reg_w_lg_w_lg_w_lg_q812w813w814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 is_bonded_reconfig_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF is_bonded_reconfig_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 logical_pll_num_reg	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF logical_pll_num_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 mif_stage	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF mif_stage : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_mif_stage_sclr	:	STD_LOGIC;
	 SIGNAL  wire_mif_stage_w_lg_q284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_mif_type_reg_d	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 mif_type_reg	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF mif_type_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_mif_type_reg_ena	:	STD_LOGIC_VECTOR(4 DOWNTO 0);
	 SIGNAL	 wire_mif_type_reg_sclr	:	STD_LOGIC_VECTOR(4 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w984w985w986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range844w980w981w982w983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range865w866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range865w979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range856w857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range851w852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range847w848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range844w845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w984w985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range844w980w981w982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_q_range844w980w981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range844w980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconf_mode_sel_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconf_mode_sel_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconf_mode_sel_reg_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 reconfig_data_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_data_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconfig_data_reg_ena	:	STD_LOGIC_VECTOR(15 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_lg_w_q_range824w825w826w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_q_range824w825w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range824w825w826w827w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_lg_w_q_range824w825w826w827w828w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range459w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range295w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range586w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range347w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range386w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range478w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range451w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range467w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range824w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range484w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range494w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range512w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range296w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range592w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range355w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range503w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range294w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range529w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL	 reconfig_done_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_done_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconfig_done_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_reconfig_done_reg_w_lg_q801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_done_reg_w_lg_q802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 tx_cmu_sel	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_cmu_sel : SIGNAL IS "PRESERVE_REGISTER=ON; PRESERVE_FANOUT_FREE_NODE=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_pll_inclk_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 tx_pll_inclk_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_pll_inclk_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_pll_inclk_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range544w560w561w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range540w541w558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range540w541w542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range539w543w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range539w543w579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range544w560w561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_q_range540w541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_q_range544w545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_q_range538w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_q_range539w543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_q_range540w559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_q_range544w560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_lg_w_q_range544w560w561w562w563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range539w543w547w548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range539w543w579w580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_lg_w_q_range539w543w547w548w549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range544w571w572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_lg_w_q_range544w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_q_range538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_q_range539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_q_range540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_pll_inclk_reg_w_q_range544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wr_addr_inc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_addr_inc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wr_rd_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_rd_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wr_rd_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_wr_rd_pulse_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wren_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wren_data_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wren_data_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_wren_data_reg_w_lg_w_lg_q1003w1004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q1002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q1003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q1007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_le7_out	:	STD_LOGIC;
	 SIGNAL  wire_add_sub11_w_lg_result922w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub11_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub12_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_cru_idx0_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_cru_idx0_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_rcxpat_chnl_en_ch_word_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_rcxpat_chnl_en_ch_word_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_second_mif_header_address_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_second_mif_header_address_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_is_special_address_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_special_address_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_is_table_33_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_33_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_35_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_35_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_37_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_37_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_38_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_38_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_42_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_42_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_43_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_43_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_44_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_44_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_46_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_46_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_47_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_47_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_59_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_59_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_60_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_60_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_61_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_61_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_75_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_75_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_76_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_76_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_77_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_77_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_en_mif_addr_cntr710w879w880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_data	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_clr_offset881w882w883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_sload	:	STD_LOGIC;
	 SIGNAL  wire_w891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_w_lg_w_lg_q741w742w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_w_lg_q741w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_w713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w737w738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconf_mode_dec_enable	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_idle_state278w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconf_mode_dec_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_data	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_sel	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_data	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_central_pcs_global_clk_div_mux_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_data	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_data	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data_mux_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_pll_first_word_mux_data	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_pll_first_word_mux_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_pll_first_word_mux_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_write_skip229w379w380w381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_write_skip229w426w427w428w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_write_skip229w414w415w416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_cmu912w913w914w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_cmu908w909w910w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_header_proc159w217w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w1078w1079w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_pll_reconfig420w421w610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch231w593w594w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_60535w536w578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_60535w536w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_60535w536w557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_60535w536w537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header829w830w840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header829w830w834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header829w830w838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header829w830w831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header829w830w836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w362w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w362w363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w379w380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w426w427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w414w415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_diff_mif_reconfig_address884w885w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain1013w1014w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_central_pcs977w978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cmu912w913w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cmu908w909w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_diff_mif818w821w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_mif_header292w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_mif_header797w798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch595w596w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_second_mif_header724w725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_60550w581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_60550w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_60550w551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_60550w573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1237w239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_reconfig_addr160w161w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_state693w694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_word_done1046w1047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_mif_header280w281w282w283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w894w896w897w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy60w99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy60w83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy60w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy60w61w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_header_proc159w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_analog_control154w155w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_global_clk_div5w6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_reconfig13w14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_channel_reconfig408w409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cruclk_addr0230w1062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cruclk_addr0230w892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cruclk_addr0230w1068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cruclk_addr0230w1073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cruclk_addr0230w1078w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_diff_mif167w804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_pll_reconfig420w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch231w593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_339w10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_60535w536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_61899w903w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_mif_header829w830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mif_reconfig_done698w740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mif_rx_only969w970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w460w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w587w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w348w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w387w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w479w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w452w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w468w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w485w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w495w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w513w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w405w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w356w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w504w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip229w530w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_reconfig_mode_sel_range51w52w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rx_mif_type1083w1084w1085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_read_address156w157w158w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_address162w163w164w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w894w895w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w1030w1031w1032w1033w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_pma_mif_type1087w1088w1089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_tier_11015w1016w1017w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip422w423w424w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip410w411w412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain_68_6B1020w1021w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cruclk_addr01069w1070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_mif_header280w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_59670w671w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tx_local_div_ctrl639w640w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip375w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip359w367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip359w360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip359w400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_channel_address_range93w94w95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_channel_address_range78w79w80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_logical_pll_sel_num_range90w91w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_logical_pll_sel_num_range74w75w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy62w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_offset822w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_second_mif_head_out196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_diff_mif_reconfig_addr_load889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_diff_mif_reconfig_addr_ready187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_diff_mif_reconfig_address884w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain1013w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_64_671022w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_7c_7f1019w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_7c_7f_inv1018w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_preemp1t1025w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_vodctrl1027w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_en_mif_addr_cntr710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs906w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_channel_reconfig842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cmu912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cmu616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cmu908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cruclk_addr0674w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_diff_mif613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_diff_mif818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_end_mif795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_global_clk_div_mode907w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_header177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_header292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_header797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_reconfig861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_reconfig721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_mif_type1083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pma915w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_second_mif_header724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_33673w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_35672w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_37665w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_38664w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_42663w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_43662w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_44661w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_46660w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_47659w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_5973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_60550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_61904w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_6188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_61669w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_75668w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_76667w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_77666w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_merged_dprioin658w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_reconfig_done805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_rx_only968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address156w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse1010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse1008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_address162w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_all21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_reconfig_addr160w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip458w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip585w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip346w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip385w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip477w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip450w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip466w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip483w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip493w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip511w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip404w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip591w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip354w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip502w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip528w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_done1046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_out_range1092w1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_pll_sel_wire_range361w370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_mif_header280w281w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w894w896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w656w657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bonded_skip228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_offset823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_header_proc159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_global_clk_div5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cent_clk_div911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_channel_reconfig408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cruclk_addr0230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_diff_mif167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_end_mif739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_global_clk_div_mode226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_d220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_stage790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_address77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_reconfig420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_reset_stage996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_protected_bit227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pcs850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pma864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_60535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_61899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_local_div_ctrl1066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_pcs846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_pma855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_mif_header829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_reconfig_done698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_rx_only969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rd_pulse114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconf_done_reg_out697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_reconf_addr216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_system776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rx_reconfig617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s2_to_042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tx_reconfig615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_done221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_mif_word_done291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_reconfig_mode_sel_range50w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_reconfig_mode_sel_range51w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_pll_sel_wire_range361w377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w429w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w372w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w372w401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w363w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_mif_header797w798w799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch595w596w597w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_60550w581w582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_60550w565w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_60550w551w552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_60550w573w574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div5w6w7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w1062w1063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w892w893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_339w10w11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_mif_rx_only969w970w971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w342w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w328w329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w315w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w335w336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w602w603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w460w461w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w587w588w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w348w349w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w387w388w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w479w480w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w452w453w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w468w469w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w485w486w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w444w445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w495w496w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w513w514w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w405w406w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w356w357w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w439w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w504w505w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w396w397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip229w530w531w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_w97w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_channel_address_range93w94w95w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_channel_address_range78w79w80w81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy62w63w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy101w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy85w86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy70w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain_vodctrl1027w1028w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_channel_reconfig842w843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_pll_reconfig861w862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_pll_reconfig721w722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rx_mif_type1083w1084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_61904w905w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address156w157w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_address162w163w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w1094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_tx_pll_sel_wire_range361w370w371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_reconfig13w20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_reconfig13w378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_339w886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_339w706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1185w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1185w215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_mif_header797w798w799w800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w598w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w581w582w583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w565w566w567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w551w552w553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w573w574w575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl1027w1028w1029w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_pll_reconfig861w862w863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_pll_reconfig721w722w723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_339w706w707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_339w706w876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1030w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_table_339w706w876w877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w1030w1031w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w1030w1031w1032w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w650w651w652w653w654w655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w650w651w652w653w654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w650w651w652w653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w650w651w652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w650w651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w644w645w646w647w648w649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w644w645w646w647w648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w644w645w646w647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w644w645w646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w181w182w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w644w645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w181w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w212w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_table_33625w641w642w643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_cruclk_addr0192w193w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_33625w641w642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_tx_pcs606w607w608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_clr_offset881w882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_delay_mif_head_out1042w1043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_adce30w31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cruclk_addr01074w1075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_cruclk_addr0192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_pll_address66w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_pma_mif_type1087w1088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rx_pma920w921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_33625w641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_11015w1016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tx_pcs606w607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_mif_header819w820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip422w423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip410w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_word_preemp1t_data_valid1023w1024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_offset881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_mif_head_out197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_mif_head_out1042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_diff_mif_wr_rd_busy612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_68_6B1020w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_adce30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_channel_reconfig413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cruclk_addr01069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cruclk_addr01074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cruclk_addr0192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_header280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_stage792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_address66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_reconfig425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pma_mif_type1087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pma920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_33625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_351061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_59670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_11015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_local_div_ctrl639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_pcs606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_mif_header819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_system207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_preemp1t_data_valid1023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_vodctrl_data_valid1026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_range93w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_range78w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_out_range1096w1097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_logical_pll_sel_num_range90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_logical_pll_sel_num_range74w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_reconfig_mode_sel_range51w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  a2gr_dprio_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_rden :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren_data :	STD_LOGIC;
	 SIGNAL  adce_busy_state :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_state :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  add_sub_datab :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  add_sub_sel :	STD_LOGIC;
	 SIGNAL  aeq_ch_done :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  bonded_skip :	STD_LOGIC;
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  cal_busy :	STD_LOGIC;
	 SIGNAL  cal_channel_address :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_channel_address_out :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_dprio_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  cal_dprioout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cal_quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  cal_testbuses :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_clk_div_plus_one :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  central_pcs_first_word_addr :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  central_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  central_pcs_minus_one :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  central_pcs_plus_seven :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  channel_address :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  channel_address_out :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  clr_offset :	STD_LOGIC;
	 SIGNAL  cmu_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  cmu_pll_plus_three :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  cruclk_mux_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  delay_mif_head_out :	STD_LOGIC;
	 SIGNAL  delay_second_mif_head_out :	STD_LOGIC;
	 SIGNAL  dfe_busy :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  diff_mif_address_busy :	STD_LOGIC;
	 SIGNAL  diff_mif_clr_offset :	STD_LOGIC;
	 SIGNAL  diff_mif_load_mif_header :	STD_LOGIC;
	 SIGNAL  diff_mif_mif_header :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  diff_mif_reconfig_addr_load :	STD_LOGIC;
	 SIGNAL  diff_mif_reconfig_addr_ready :	STD_LOGIC;
	 SIGNAL  diff_mif_reconfig_addr_start :	STD_LOGIC;
	 SIGNAL  diff_mif_reconfig_address :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  diff_mif_wr_rd_busy :	STD_LOGIC;
	 SIGNAL  dprio_addr_index :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_addr_offset_cmpr_datab :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_addr_offset_cnt_out :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_addr_translated_offset :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_64_67 :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_68_6B :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_7c_7f :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_7c_7f_inv :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_preemp1t :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_vodctrl :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_pulse :	STD_LOGIC;
	 SIGNAL  dprio_wr_done :	STD_LOGIC;
	 SIGNAL  duplex_pma_first_pll :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  duplex_pma_pcs_first_pll :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  en_mif_addr_cntr :	STD_LOGIC;
	 SIGNAL  en_write_trigger :	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_busy :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  global_clk_div_addr :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  global_clk_div_addr_offset :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  global_clk_div_mode_offset_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  global_clk_div_mode_plus_five :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  global_register_reset :	STD_LOGIC;
	 SIGNAL  header_proc :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  internal_write_pulse :	STD_LOGIC;
	 SIGNAL  is_adce :	STD_LOGIC;
	 SIGNAL  is_adce_all_control :	STD_LOGIC;
	 SIGNAL  is_adce_continuous_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_one_time_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_standby_single_control :	STD_LOGIC;
	 SIGNAL  is_analog_control :	STD_LOGIC;
	 SIGNAL  is_bonded_global_clk_div :	STD_LOGIC;
	 SIGNAL  is_bonded_reconfig :	STD_LOGIC;
	 SIGNAL  is_cent_clk_div :	STD_LOGIC;
	 SIGNAL  is_central_pcs :	STD_LOGIC;
	 SIGNAL  is_channel_reconfig :	STD_LOGIC;
	 SIGNAL  is_cmu :	STD_LOGIC;
	 SIGNAL  is_cruclk_addr0 :	STD_LOGIC;
	 SIGNAL  is_diff_mif :	STD_LOGIC;
	 SIGNAL  is_do_dfe :	STD_LOGIC;
	 SIGNAL  is_do_eyemon :	STD_LOGIC;
	 SIGNAL  is_end_mif :	STD_LOGIC;
	 SIGNAL  is_global_clk_div_mode :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_d :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_out :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  is_mif_header :	STD_LOGIC;
	 SIGNAL  is_mif_stage :	STD_LOGIC;
	 SIGNAL  is_offset_end :	STD_LOGIC;
	 SIGNAL  is_pll_address :	STD_LOGIC;
	 SIGNAL  is_pll_end_mif :	STD_LOGIC;
	 SIGNAL  is_pll_first_word :	STD_LOGIC;
	 SIGNAL  is_pll_reconfig :	STD_LOGIC;
	 SIGNAL  is_pll_reset_stage :	STD_LOGIC;
	 SIGNAL  is_pma_mif_type :	STD_LOGIC;
	 SIGNAL  is_protected_bit :	STD_LOGIC;
	 SIGNAL  is_rcxpat_chnl_en_ch :	STD_LOGIC;
	 SIGNAL  is_rx_mif_type :	STD_LOGIC;
	 SIGNAL  is_rx_pcs :	STD_LOGIC;
	 SIGNAL  is_rx_pma :	STD_LOGIC;
	 SIGNAL  is_second_mif_header :	STD_LOGIC;
	 SIGNAL  is_table_33 :	STD_LOGIC;
	 SIGNAL  is_table_35 :	STD_LOGIC;
	 SIGNAL  is_table_37 :	STD_LOGIC;
	 SIGNAL  is_table_38 :	STD_LOGIC;
	 SIGNAL  is_table_42 :	STD_LOGIC;
	 SIGNAL  is_table_43 :	STD_LOGIC;
	 SIGNAL  is_table_44 :	STD_LOGIC;
	 SIGNAL  is_table_46 :	STD_LOGIC;
	 SIGNAL  is_table_47 :	STD_LOGIC;
	 SIGNAL  is_table_59 :	STD_LOGIC;
	 SIGNAL  is_table_60 :	STD_LOGIC;
	 SIGNAL  is_table_61 :	STD_LOGIC;
	 SIGNAL  is_table_75 :	STD_LOGIC;
	 SIGNAL  is_table_76 :	STD_LOGIC;
	 SIGNAL  is_table_77 :	STD_LOGIC;
	 SIGNAL  is_tier_1 :	STD_LOGIC;
	 SIGNAL  is_tier_2 :	STD_LOGIC;
	 SIGNAL  is_tx_local_div_ctrl :	STD_LOGIC;
	 SIGNAL  is_tx_pcs :	STD_LOGIC;
	 SIGNAL  is_tx_pma :	STD_LOGIC;
	 SIGNAL  legal_wr_mode_type :	STD_LOGIC;
	 SIGNAL  load_mif_header :	STD_LOGIC;
	 SIGNAL  local_ch_dec :	STD_LOGIC;
	 SIGNAL  logical_pll_sel_num :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  merged_dprioin :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  mif_addr_cntr_data :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mif_reconfig_done :	STD_LOGIC;
	 SIGNAL  mif_rx_only :	STD_LOGIC;
	 SIGNAL  offset_cancellation_reset	:	STD_LOGIC;
	 SIGNAL  pll_first_word_addr :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  quad_address_out :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  rd_pulse :	STD_LOGIC;
	 SIGNAL  read_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  read_reconfig_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  reconf_done_reg_out :	STD_LOGIC;
	 SIGNAL  reconfig_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  reconfig_reset_all :	STD_LOGIC;
	 SIGNAL  reset_addr_done :	STD_LOGIC;
	 SIGNAL  reset_reconf_addr :	STD_LOGIC;
	 SIGNAL  reset_system :	STD_LOGIC;
	 SIGNAL  rx_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_pma_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_pma_minus_one :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_reconfig :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s0_to_2 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  start	:	STD_LOGIC;
	 SIGNAL  state_mc_reg_in :	STD_LOGIC_VECTOR (0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  table_33_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_35_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_37_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_38_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_42_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_43_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_44_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_46_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_47_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_59_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_61_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_75_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_76_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_77_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  transceiver_init	:	STD_LOGIC;
	 SIGNAL  tx_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  tx_pll_sel_wire :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  tx_pma_first_pll :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  tx_pma_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  tx_pma_pcs_first_pll :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  tx_reconfig :	STD_LOGIC;
	 SIGNAL  wr_pulse :	STD_LOGIC;
	 SIGNAL  write_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  write_all_int :	STD_LOGIC;
	 SIGNAL  write_done :	STD_LOGIC;
	 SIGNAL  write_happened :	STD_LOGIC;
	 SIGNAL  write_mif_word_done :	STD_LOGIC;
	 SIGNAL  write_reconfig_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  write_skip :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 SIGNAL  write_word_64_67_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_68_6B_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_7c_7f_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_7c_7f_inv_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_done :	STD_LOGIC;
	 SIGNAL  write_word_preemp1t_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_preemp1ta_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_preemp1tb_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_vodctrl_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_vodctrla_data_valid :	STD_LOGIC;
	 SIGNAL  wire_w_cal_channel_address_range100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_channel_address_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_channel_address_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_out_range1092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_out_range1096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dprio_addr_index_range1060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dprio_addr_index_range1067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dprio_addr_index_range1072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dprio_addr_index_range1077w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_logical_pll_sel_num_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_logical_pll_sel_num_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_reconfig_mode_sel_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_reconfig_mode_sel_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_reconfig_mode_sel_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_pll_sel_wire_range369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_pll_sel_wire_range361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_pll_sel_wire_range368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  alt_cal
	 GENERIC 
	 (
		CHANNEL_ADDRESS_WIDTH	:	NATURAL := 1;
		NUMBER_OF_CHANNELS	:	NATURAL;
		SIM_MODEL_MODE	:	STRING := "FALSE";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "alt_cal"
	 );
	 PORT
	 ( 
		busy	:	OUT STD_LOGIC;
		cal_error	:	OUT STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0);
		clock	:	IN STD_LOGIC;
		dprio_addr	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_busy	:	IN STD_LOGIC;
		dprio_datain	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_dataout	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_rden	:	OUT STD_LOGIC;
		dprio_wren	:	OUT STD_LOGIC;
		quad_addr	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		remap_addr	:	IN STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		reset	:	IN STD_LOGIC := '0';
		retain_addr	:	OUT STD_LOGIC;
		start	:	IN STD_LOGIC := '0';
		testbuses	:	IN STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS*4-1 DOWNTO 0) := (OTHERS => '0');
		transceiver_init	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_reconfig_cpri_alt_dprio_t2l
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		busy	:	OUT  STD_LOGIC;
		datain	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		dpclk	:	IN  STD_LOGIC;
		dpriodisable	:	OUT  STD_LOGIC;
		dprioin	:	OUT  STD_LOGIC;
		dprioload	:	OUT  STD_LOGIC;
		dprioout	:	IN  STD_LOGIC;
		quad_address	:	IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		rden	:	IN  STD_LOGIC := '0';
		reset	:	IN  STD_LOGIC := '0';
		status_out	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		wren	:	IN  STD_LOGIC := '0';
		wren_data	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lcell
	 PORT
	 ( 
		a_in	:	IN STD_LOGIC;
		a_out	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_reconfig_cpri_mux_r7a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(59 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_reconfig_cpri_mux_a6a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(14 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_reconfig_cpri_mux_d6a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(24 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_reconfig_cpri_mux_b6a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(17 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_reconfig_cpri_mux_c6a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_w_lg_write_skip229w379w380w381w(0) <= wire_w_lg_w_lg_w_lg_write_skip229w379w380w(0) AND wire_w_lg_w_tx_pll_sel_wire_range361w377w(0);
	loop11 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_write_skip229w426w427w428w(i) <= wire_w_lg_w_lg_w_lg_write_skip229w426w427w(0) AND wire_reconfig_data_reg_w_q_range386w(i);
	END GENERATE loop11;
	wire_w_lg_w_lg_w_lg_w_lg_write_skip229w414w415w416w(0) <= wire_w_lg_w_lg_w_lg_write_skip229w414w415w(0) AND wire_w_tx_pll_sel_wire_range369w(0);
	loop12 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_is_cmu912w913w914w(i) <= wire_w_lg_w_lg_is_cmu912w913w(i) AND wire_w_lg_is_global_clk_div_mode226w(0);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_is_cmu908w909w910w(i) <= wire_w_lg_w_lg_is_cmu908w909w(i) AND wire_w_lg_is_global_clk_div_mode226w(0);
	END GENERATE loop13;
	wire_w_lg_w_lg_w_lg_header_proc159w217w218w(0) <= wire_w_lg_w_lg_header_proc159w217w(0) AND wire_w_lg_w_lg_is_tier_1185w215w(0);
	loop14 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w1078w1079w(i) <= wire_w_lg_w_lg_is_cruclk_addr0230w1078w(i) AND wire_w_lg_is_tx_local_div_ctrl1066w(0);
	END GENERATE loop14;
	wire_w_lg_w_lg_w_lg_is_pll_reconfig420w421w610w(0) <= wire_w_lg_w_lg_is_pll_reconfig420w421w(0) AND is_cmu;
	loop15 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch231w593w594w(i) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch231w593w(0) AND wire_reconfig_data_reg_w_q_range592w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_w_lg_is_table_60535w536w578w(0) <= wire_w_lg_w_lg_is_table_60535w536w(0) AND wire_reconfig_data_reg_w_q_range577w(0);
	wire_w_lg_w_lg_w_lg_is_table_60535w536w570w(0) <= wire_w_lg_w_lg_is_table_60535w536w(0) AND wire_reconfig_data_reg_w_q_range569w(0);
	wire_w_lg_w_lg_w_lg_is_table_60535w536w557w(0) <= wire_w_lg_w_lg_is_table_60535w536w(0) AND wire_reconfig_data_reg_w_q_range556w(0);
	wire_w_lg_w_lg_w_lg_is_table_60535w536w537w(0) <= wire_w_lg_w_lg_is_table_60535w536w(0) AND wire_reconfig_data_reg_w_q_range443w(0);
	wire_w_lg_w_lg_w_lg_load_mif_header829w830w840w(0) <= wire_w_lg_w_lg_load_mif_header829w830w(0) AND is_cmu;
	wire_w_lg_w_lg_w_lg_load_mif_header829w830w834w(0) <= wire_w_lg_w_lg_load_mif_header829w830w(0) AND is_rx_pcs;
	wire_w_lg_w_lg_w_lg_load_mif_header829w830w838w(0) <= wire_w_lg_w_lg_load_mif_header829w830w(0) AND is_rx_pma;
	wire_w_lg_w_lg_w_lg_load_mif_header829w830w831w(0) <= wire_w_lg_w_lg_load_mif_header829w830w(0) AND is_tx_pcs;
	wire_w_lg_w_lg_w_lg_load_mif_header829w830w836w(0) <= wire_w_lg_w_lg_load_mif_header829w830w(0) AND is_tx_pma;
	wire_w_lg_w_lg_w_lg_write_skip229w362w372w(0) <= wire_w_lg_w_lg_write_skip229w362w(0) AND wire_w_lg_w_lg_w_tx_pll_sel_wire_range361w370w371w(0);
	wire_w_lg_w_lg_w_lg_write_skip229w362w363w(0) <= wire_w_lg_w_lg_write_skip229w362w(0) AND wire_w_tx_pll_sel_wire_range361w(0);
	wire_w_lg_w_lg_w_lg_write_skip229w379w380w(0) <= wire_w_lg_w_lg_write_skip229w379w(0) AND wire_w_tx_pll_sel_wire_range369w(0);
	wire_w_lg_w_lg_w_lg_write_skip229w426w427w(0) <= wire_w_lg_w_lg_write_skip229w426w(0) AND is_bonded_reconfig;
	wire_w_lg_w_lg_w_lg_write_skip229w414w415w(0) <= wire_w_lg_w_lg_write_skip229w414w(0) AND wire_w_lg_is_channel_reconfig413w(0);
	wire_w57w(0) <= wire_w_lg_w_lg_w_reconfig_mode_sel_range51w52w56w(0) AND wire_w_lg_w_reconfig_mode_sel_range50w55w(0);
	loop16 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_diff_mif_reconfig_address884w885w(i) <= wire_w_lg_diff_mif_reconfig_address884w(i) AND is_diff_mif;
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain1013w1014w(i) <= wire_w_lg_dprio_datain1013w(i) AND write_state;
	END GENERATE loop17;
	wire_w_lg_w_lg_is_central_pcs977w978w(0) <= wire_w_lg_is_central_pcs977w(0) AND dprio_pulse;
	loop18 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_is_cmu912w913w(i) <= wire_w_lg_is_cmu912w(0) AND cmu_pll_plus_three(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_is_cmu908w909w(i) <= wire_w_lg_is_cmu908w(0) AND cent_clk_div_plus_one(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_is_diff_mif818w821w(i) <= wire_w_lg_is_diff_mif818w(0) AND diff_mif_mif_header(i);
	END GENERATE loop20;
	wire_w_lg_w_lg_is_mif_header292w293w(0) <= wire_w_lg_is_mif_header292w(0) AND is_tier_1;
	wire_w_lg_w_lg_is_mif_header797w798w(0) <= wire_w_lg_is_mif_header797w(0) AND is_tier_1;
	loop21 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_is_rcxpat_chnl_en_ch595w596w(i) <= wire_w_lg_is_rcxpat_chnl_en_ch595w(0) AND wire_dprio_dataout_reg_w_q_range590w(i);
	END GENERATE loop21;
	wire_w_lg_w_lg_is_second_mif_header724w725w(0) <= wire_w_lg_is_second_mif_header724w(0) AND write_state;
	wire_w_lg_w_lg_is_table_60550w581w(0) <= wire_w_lg_is_table_60550w(0) AND wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range539w543w579w580w(0);
	wire_w_lg_w_lg_is_table_60550w565w(0) <= wire_w_lg_is_table_60550w(0) AND wire_tx_pll_inclk_reg_w564w(0);
	wire_w_lg_w_lg_is_table_60550w551w(0) <= wire_w_lg_is_table_60550w(0) AND wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_lg_w_q_range539w543w547w548w549w(0);
	wire_w_lg_w_lg_is_table_60550w573w(0) <= wire_w_lg_is_table_60550w(0) AND wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range544w571w572w(0);
	wire_w_lg_w_lg_is_tier_1237w239w(0) <= wire_w_lg_is_tier_1237w(0) AND wire_w_lg_w212w213w(0);
	loop22 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_write_reconfig_addr160w161w(i) <= wire_w_lg_write_reconfig_addr160w(i) AND wire_w_lg_header_proc159w(0);
	END GENERATE loop22;
	wire_w_lg_w_lg_write_state693w694w(0) <= wire_w_lg_write_state693w(0) AND write_happened;
	wire_w_lg_w_lg_write_word_done1046w1047w(0) <= wire_w_lg_write_word_done1046w(0) AND is_analog_control;
	wire_w_lg_w_lg_w_lg_w_lg_is_mif_header280w281w282w283w(0) <= wire_w_lg_w_lg_w_lg_is_mif_header280w281w282w(0) AND mif_stage;
	loop23 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w894w896w897w(i) <= wire_w_lg_w894w896w(0) AND wire_dprio_addr_offset_cnt_q(i);
	END GENERATE loop23;
	wire_w_lg_w_lg_cal_busy60w99w(0) <= wire_w_lg_cal_busy60w(0) AND wire_w_lg_w97w98w(0);
	wire_w_lg_w_lg_cal_busy60w83w(0) <= wire_w_lg_cal_busy60w(0) AND wire_w82w(0);
	wire_w_lg_w_lg_cal_busy60w68w(0) <= wire_w_lg_cal_busy60w(0) AND wire_w_lg_w_lg_is_pll_address66w67w(0);
	loop24 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_cal_busy60w61w(i) <= wire_w_lg_cal_busy60w(0) AND quad_address(i);
	END GENERATE loop24;
	wire_w_lg_w_lg_header_proc159w217w(0) <= wire_w_lg_header_proc159w(0) AND wire_w_lg_reset_reconf_addr216w(0);
	loop25 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_is_analog_control154w155w(i) <= wire_w_lg_is_analog_control154w(0) AND read_reconfig_addr(i);
	END GENERATE loop25;
	wire_w_lg_w_lg_is_bonded_global_clk_div5w6w(0) <= wire_w_lg_is_bonded_global_clk_div5w(0) AND busy_state;
	wire_w_lg_w_lg_is_bonded_reconfig13w14w(0) <= wire_w_lg_is_bonded_reconfig13w(0) AND busy_state;
	wire_w_lg_w_lg_is_channel_reconfig408w409w(0) <= wire_w_lg_is_channel_reconfig408w(0) AND wire_w_lg_is_global_clk_div_mode226w(0);
	wire_w_lg_w_lg_is_cruclk_addr0230w1062w(0) <= wire_w_lg_is_cruclk_addr0230w(0) AND wire_w_lg_is_table_351061w(0);
	wire_w_lg_w_lg_is_cruclk_addr0230w892w(0) <= wire_w_lg_is_cruclk_addr0230w(0) AND is_rx_pma;
	wire_w_lg_w_lg_is_cruclk_addr0230w1068w(0) <= wire_w_lg_is_cruclk_addr0230w(0) AND wire_w_dprio_addr_index_range1067w(0);
	wire_w_lg_w_lg_is_cruclk_addr0230w1073w(0) <= wire_w_lg_is_cruclk_addr0230w(0) AND wire_w_dprio_addr_index_range1072w(0);
	loop26 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_is_cruclk_addr0230w1078w(i) <= wire_w_lg_is_cruclk_addr0230w(0) AND wire_w_dprio_addr_index_range1077w(i);
	END GENERATE loop26;
	wire_w_lg_w_lg_is_diff_mif167w804w(0) <= wire_w_lg_is_diff_mif167w(0) AND is_tier_1;
	wire_w_lg_w_lg_is_pll_reconfig420w421w(0) <= wire_w_lg_is_pll_reconfig420w(0) AND wire_w_lg_is_global_clk_div_mode226w(0);
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch231w593w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch231w(0) AND wire_w_lg_write_skip229w(0);
	wire_w_lg_w_lg_is_table_339w10w(0) <= wire_w_lg_is_table_339w(0) AND busy_state;
	wire_w_lg_w_lg_is_table_60535w536w(0) <= wire_w_lg_is_table_60535w(0) AND wire_w_lg_write_skip229w(0);
	loop27 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_is_table_61899w903w(i) <= wire_w_lg_is_table_61899w(0) AND central_pcs_minus_one(i);
	END GENERATE loop27;
	wire_w_lg_w_lg_load_mif_header829w830w(0) <= wire_w_lg_load_mif_header829w(0) AND clr_offset;
	wire_w_lg_w_lg_mif_reconfig_done698w740w(0) <= wire_w_lg_mif_reconfig_done698w(0) AND wire_w_lg_is_end_mif739w(0);
	wire_w_lg_w_lg_mif_rx_only969w970w(0) <= wire_w_lg_mif_rx_only969w(0) AND wire_mif_type_reg_w_q_range856w(0);
	wire_w_lg_w_lg_write_skip229w362w(0) <= wire_w_lg_write_skip229w(0) AND wire_w_lg_is_bonded_reconfig13w(0);
	wire_w_lg_w_lg_write_skip229w342w(0) <= wire_w_lg_write_skip229w(0) AND wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range305w311w340w341w(0);
	wire_w_lg_w_lg_write_skip229w379w(0) <= wire_w_lg_write_skip229w(0) AND wire_w_lg_w_lg_is_bonded_reconfig13w378w(0);
	wire_w_lg_w_lg_write_skip229w328w(0) <= wire_w_lg_write_skip229w(0) AND wire_cru_num_reg_w327w(0);
	wire_w_lg_w_lg_write_skip229w315w(0) <= wire_w_lg_write_skip229w(0) AND wire_cru_num_reg_w_lg_w_lg_w_lg_w_lg_w_q_range305w311w312w313w314w(0);
	wire_w_lg_w_lg_write_skip229w335w(0) <= wire_w_lg_write_skip229w(0) AND wire_cru_num_reg_w_lg_w_lg_w_q_range309w333w334w(0);
	wire_w_lg_w_lg_write_skip229w426w(0) <= wire_w_lg_write_skip229w(0) AND wire_w_lg_is_pll_reconfig425w(0);
	wire_w_lg_w_lg_write_skip229w414w(0) <= wire_w_lg_write_skip229w(0) AND is_bonded_reconfig;
	wire_w_lg_w_lg_write_skip229w602w(0) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range297w(0);
	loop28 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_write_skip229w460w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range459w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip229w587w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range586w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 5 GENERATE 
		wire_w_lg_w_lg_write_skip229w348w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range347w(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_w_lg_write_skip229w387w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range386w(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_w_lg_write_skip229w479w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range478w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_write_skip229w452w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range451w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip229w468w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range467w(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_write_skip229w485w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range484w(i);
	END GENERATE loop35;
	wire_w_lg_w_lg_write_skip229w444w(0) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range443w(0);
	loop36 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip229w495w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range494w(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_write_skip229w513w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range512w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_write_skip229w405w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range296w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_write_skip229w356w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range355w(i);
	END GENERATE loop39;
	wire_w_lg_w_lg_write_skip229w439w(0) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range438w(0);
	loop40 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_write_skip229w504w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range503w(i);
	END GENERATE loop40;
	wire_w_lg_w_lg_write_skip229w396w(0) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range395w(0);
	loop41 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_w_lg_write_skip229w530w(i) <= wire_w_lg_write_skip229w(0) AND wire_reconfig_data_reg_w_q_range529w(i);
	END GENERATE loop41;
	wire_w_lg_w_lg_w_reconfig_mode_sel_range51w52w56w(0) <= wire_w_lg_w_reconfig_mode_sel_range51w52w(0) AND wire_w_reconfig_mode_sel_range48w(0);
	wire_w97w(0) <= wire_w_lg_w_lg_w_lg_w_channel_address_range93w94w95w96w(0) AND wire_w_lg_is_central_pcs89w(0);
	wire_w_lg_w_lg_w_lg_is_rx_mif_type1083w1084w1085w(0) <= wire_w_lg_w_lg_is_rx_mif_type1083w1084w(0) AND wire_w_lg_is_central_pcs89w(0);
	loop42 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_read_address156w157w158w(i) <= wire_w_lg_w_lg_read_address156w157w(i) AND read_state;
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_write_address162w163w164w(i) <= wire_w_lg_w_lg_write_address162w163w(i) AND write_state;
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w894w895w(i) <= wire_w894w(0) AND dprio_addr_translated_offset(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_w1030w1031w1032w1033w(i) <= wire_w_lg_w_lg_w1030w1031w1032w(i) AND is_analog_control;
	END GENERATE loop45;
	wire_w_lg_w_lg_w_lg_is_pma_mif_type1087w1088w1089w(0) <= wire_w_lg_w_lg_is_pma_mif_type1087w1088w(0) AND wire_w_lg_is_central_pcs89w(0);
	loop46 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_is_tier_11015w1016w1017w(i) <= wire_w_lg_w_lg_is_tier_11015w1016w(0) AND reconfig_datain(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip422w423w424w(i) <= wire_w_lg_w_lg_write_skip422w423w(0) AND wire_dprio_dataout_reg_w_q_range384w(i);
	END GENERATE loop47;
	wire_w_lg_w_lg_w_lg_write_skip410w411w412w(0) <= wire_w_lg_w_lg_write_skip410w411w(0) AND wire_dprio_dataout_reg_w_q_range331w(0);
	loop48 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain_68_6B1020w1021w(i) <= wire_w_lg_dprio_datain_68_6B1020w(i) AND write_word_68_6B_data_valid;
	END GENERATE loop48;
	wire_w_lg_w_lg_is_cruclk_addr01069w1070w(0) <= wire_w_lg_is_cruclk_addr01069w(0) AND wire_w_lg_is_tx_local_div_ctrl1066w(0);
	wire_w_lg_w_lg_is_mif_header280w281w(0) <= wire_w_lg_is_mif_header280w(0) AND dprio_pulse;
	loop49 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_is_table_59670w671w(i) <= wire_w_lg_is_table_59670w(0) AND table_59_data(i);
	END GENERATE loop49;
	loop50 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_is_tx_local_div_ctrl639w640w(i) <= wire_w_lg_is_tx_local_div_ctrl639w(0) AND dprio_dataout_reg(i);
	END GENERATE loop50;
	wire_w_lg_w_lg_write_skip375w376w(0) <= wire_w_lg_write_skip375w(0) AND wire_dprio_dataout_reg_w_q_range331w(0);
	wire_w_lg_w_lg_write_skip359w367w(0) <= wire_w_lg_write_skip359w(0) AND wire_dprio_dataout_reg_w_q_range319w(0);
	wire_w_lg_w_lg_write_skip359w360w(0) <= wire_w_lg_write_skip359w(0) AND wire_dprio_dataout_reg_w_q_range302w(0);
	wire_w_lg_w_lg_write_skip359w400w(0) <= wire_w_lg_write_skip359w(0) AND wire_dprio_dataout_reg_w_q_range399w(0);
	wire_w_lg_w_lg_w_channel_address_range93w94w95w(0) <= wire_w_lg_w_channel_address_range93w94w(0) AND wire_w_lg_is_pll_address77w(0);
	wire_w_lg_w_lg_w_channel_address_range78w79w80w(0) <= wire_w_lg_w_channel_address_range78w79w(0) AND wire_w_lg_is_pll_address77w(0);
	wire_w_lg_w_lg_w_logical_pll_sel_num_range90w91w92w(0) <= wire_w_lg_w_logical_pll_sel_num_range90w91w(0) AND is_pll_address;
	wire_w_lg_w_lg_w_logical_pll_sel_num_range74w75w76w(0) <= wire_w_lg_w_logical_pll_sel_num_range74w75w(0) AND is_pll_address;
	loop51 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_cal_busy62w(i) <= cal_busy AND cal_quad_address(i);
	END GENERATE loop51;
	wire_w_lg_cal_busy101w(0) <= cal_busy AND wire_w_cal_channel_address_range100w(0);
	wire_w_lg_cal_busy85w(0) <= cal_busy AND wire_w_cal_channel_address_range84w(0);
	wire_w_lg_cal_busy70w(0) <= cal_busy AND wire_w_cal_channel_address_range69w(0);
	loop52 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_clr_offset822w(i) <= clr_offset AND mif_type_reg(i);
	END GENERATE loop52;
	wire_w_lg_delay_second_mif_head_out196w(0) <= delay_second_mif_head_out AND wire_w195w(0);
	wire_w_lg_diff_mif_reconfig_addr_load889w(0) <= diff_mif_reconfig_addr_load AND wire_w_lg_is_bonded_reconfig13w(0);
	wire_w_lg_diff_mif_reconfig_addr_ready187w(0) <= diff_mif_reconfig_addr_ready AND is_diff_mif;
	loop53 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_diff_mif_reconfig_address884w(i) <= diff_mif_reconfig_address(i) AND diff_mif_address_busy;
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain1013w(i) <= dprio_datain(i) AND wire_w_lg_header_proc159w(0);
	END GENERATE loop54;
	loop55 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_64_671022w(i) <= dprio_datain_64_67(i) AND write_word_64_67_data_valid;
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_7c_7f1019w(i) <= dprio_datain_7c_7f(i) AND write_word_7c_7f_data_valid;
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_7c_7f_inv1018w(i) <= dprio_datain_7c_7f_inv(i) AND write_word_7c_7f_inv_data_valid;
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_preemp1t1025w(i) <= dprio_datain_preemp1t(i) AND wire_w_lg_w_lg_write_word_preemp1t_data_valid1023w1024w(0);
	END GENERATE loop58;
	loop59 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_vodctrl1027w(i) <= dprio_datain_vodctrl(i) AND wire_w_lg_write_word_vodctrl_data_valid1026w(0);
	END GENERATE loop59;
	wire_w_lg_dprio_pulse279w(0) <= dprio_pulse AND wire_w_lg_idle_state278w(0);
	wire_w_lg_en_mif_addr_cntr710w(0) <= en_mif_addr_cntr AND wire_w_lg_is_bonded_reconfig13w(0);
	wire_w_lg_idle_state791w(0) <= idle_state AND wire_w_lg_is_mif_stage790w(0);
	wire_w_lg_idle_state290w(0) <= idle_state AND wire_mif_stage_w_lg_q284w(0);
	wire_w_lg_idle_state32w(0) <= idle_state AND wire_w_lg_w_lg_is_adce30w31w(0);
	wire_w_lg_idle_state605w(0) <= idle_state AND write_all;
	wire_w_lg_is_bonded_reconfig19w(0) <= is_bonded_reconfig AND wire_w_lg_is_bonded_global_clk_div5w(0);
	wire_w_lg_is_bonded_reconfig12w(0) <= is_bonded_reconfig AND wire_w_lg_w_lg_w_lg_is_table_339w10w11w(0);
	wire_w_lg_is_central_pcs900w(0) <= is_central_pcs AND wire_w_lg_is_table_61899w(0);
	loop60 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_central_pcs906w(i) <= is_central_pcs AND wire_w_lg_w_lg_is_table_61904w905w(i);
	END GENERATE loop60;
	wire_w_lg_is_central_pcs977w(0) <= is_central_pcs AND is_offset_end;
	wire_w_lg_is_channel_reconfig842w(0) <= is_channel_reconfig AND wire_w_lg_is_central_pcs89w(0);
	wire_w_lg_is_cmu912w(0) <= is_cmu AND wire_w_lg_is_cent_clk_div911w(0);
	wire_w_lg_is_cmu616w(0) <= is_cmu AND wire_w_lg_tx_reconfig615w(0);
	wire_w_lg_is_cmu908w(0) <= is_cmu AND is_cent_clk_div;
	loop61 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_cruclk_addr0674w(i) <= is_cruclk_addr0 AND cruclk_mux_data(i);
	END GENERATE loop61;
	wire_w_lg_is_diff_mif613w(0) <= is_diff_mif AND wire_w_lg_diff_mif_wr_rd_busy612w(0);
	wire_w_lg_is_diff_mif818w(0) <= is_diff_mif AND diff_mif_load_mif_header;
	wire_w_lg_is_end_mif795w(0) <= is_end_mif AND is_diff_mif;
	loop62 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_global_clk_div_mode907w(i) <= is_global_clk_div_mode AND global_clk_div_mode_plus_five(i);
	END GENERATE loop62;
	wire_w_lg_is_mif_header177w(0) <= is_mif_header AND wire_w_lg_is_diff_mif167w(0);
	wire_w_lg_is_mif_header292w(0) <= is_mif_header AND wire_w_lg_write_mif_word_done291w(0);
	wire_w_lg_is_mif_header797w(0) <= is_mif_header AND wire_w_lg_write_state796w(0);
	wire_w_lg_is_pll_reconfig861w(0) <= is_pll_reconfig AND wire_w_lg_is_central_pcs89w(0);
	wire_w_lg_is_pll_reconfig721w(0) <= is_pll_reconfig AND wire_w_lg_is_channel_reconfig408w(0);
	wire_w_lg_is_rcxpat_chnl_en_ch595w(0) <= is_rcxpat_chnl_en_ch AND wire_w_lg_write_skip229w(0);
	wire_w_lg_is_rx_mif_type1083w(0) <= is_rx_mif_type AND wire_w_lg_is_cruclk_addr0230w(0);
	loop63 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_rx_pma915w(i) <= is_rx_pma AND rx_pma_minus_one(i);
	END GENERATE loop63;
	wire_w_lg_is_second_mif_header724w(0) <= is_second_mif_header AND wire_w_lg_write_done221w(0);
	wire_w_lg_is_table_338w(0) <= is_table_33 AND wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div5w6w7w(0);
	loop64 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_33673w(i) <= is_table_33 AND table_33_data(i);
	END GENERATE loop64;
	loop65 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_35672w(i) <= is_table_35 AND table_35_data(i);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_37665w(i) <= is_table_37 AND table_37_data(i);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_38664w(i) <= is_table_38 AND table_38_data(i);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_42663w(i) <= is_table_42 AND table_42_data(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_43662w(i) <= is_table_43 AND table_43_data(i);
	END GENERATE loop69;
	loop70 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_44661w(i) <= is_table_44 AND table_44_data(i);
	END GENERATE loop70;
	loop71 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_46660w(i) <= is_table_46 AND table_46_data(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_47659w(i) <= is_table_47 AND table_47_data(i);
	END GENERATE loop72;
	wire_w_lg_is_table_5973w(0) <= is_table_59 AND is_bonded_reconfig;
	wire_w_lg_is_table_60550w(0) <= is_table_60 AND wire_w_lg_write_skip229w(0);
	loop73 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_table_61904w(i) <= is_table_61 AND central_pcs_plus_seven(i);
	END GENERATE loop73;
	wire_w_lg_is_table_6188w(0) <= is_table_61 AND is_central_pcs;
	loop74 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_61669w(i) <= is_table_61 AND table_61_data(i);
	END GENERATE loop74;
	loop75 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_75668w(i) <= is_table_75 AND table_75_data(i);
	END GENERATE loop75;
	loop76 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_76667w(i) <= is_table_76 AND table_76_data(i);
	END GENERATE loop76;
	loop77 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_77666w(i) <= is_table_77 AND table_77_data(i);
	END GENERATE loop77;
	wire_w_lg_is_tier_1237w(0) <= is_tier_1 AND wire_w_lg_header_proc159w(0);
	wire_w_lg_is_tier_1184w(0) <= is_tier_1 AND wire_w_lg_w_lg_w181w182w183w(0);
	wire_w_lg_is_tier_1214w(0) <= is_tier_1 AND wire_w_lg_w212w213w(0);
	wire_w_lg_is_tier_1175w(0) <= is_tier_1 AND mif_reconfig_done;
	loop78 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_merged_dprioin658w(i) <= merged_dprioin(i) AND wire_w_lg_w656w657w(0);
	END GENERATE loop78;
	wire_w_lg_mif_reconfig_done805w(0) <= mif_reconfig_done AND wire_w_lg_w_lg_is_diff_mif167w804w(0);
	wire_w_lg_mif_rx_only968w(0) <= mif_rx_only AND wire_mif_type_reg_w_q_range847w(0);
	loop79 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_read_address156w(i) <= read_address(i) AND is_analog_control;
	END GENERATE loop79;
	wire_w_lg_wr_pulse1010w(0) <= wr_pulse AND wire_wren_data_reg_w_lg_q1003w(0);
	wire_w_lg_wr_pulse1008w(0) <= wr_pulse AND wire_wren_data_reg_w_lg_q1007w(0);
	loop80 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_address162w(i) <= write_address(i) AND is_analog_control;
	END GENERATE loop80;
	wire_w_lg_write_all21w(0) <= write_all AND wire_w_lg_w_lg_is_bonded_reconfig13w20w(0);
	loop81 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_reconfig_addr160w(i) <= write_reconfig_addr(i) AND wire_w_lg_is_analog_control154w(0);
	END GENERATE loop81;
	wire_w_lg_write_skip601w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range600w(0);
	loop82 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_write_skip458w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range457w(i);
	END GENERATE loop82;
	loop83 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip585w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range489w(i);
	END GENERATE loop83;
	loop84 : FOR i IN 0 TO 5 GENERATE 
		wire_w_lg_write_skip346w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range345w(i);
	END GENERATE loop84;
	loop85 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_write_skip385w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range384w(i);
	END GENERATE loop85;
	wire_w_lg_write_skip339w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range338w(0);
	loop86 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_write_skip477w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range476w(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_write_skip450w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range449w(i);
	END GENERATE loop87;
	wire_w_lg_write_skip332w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range331w(0);
	wire_w_lg_write_skip320w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range319w(0);
	loop88 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip466w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range465w(i);
	END GENERATE loop88;
	loop89 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_skip483w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range482w(i);
	END GENERATE loop89;
	wire_w_lg_write_skip303w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range302w(0);
	loop90 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip493w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range492w(i);
	END GENERATE loop90;
	loop91 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_write_skip511w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range510w(i);
	END GENERATE loop91;
	loop92 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_write_skip404w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range403w(i);
	END GENERATE loop92;
	loop93 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_write_skip591w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range590w(i);
	END GENERATE loop93;
	loop94 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_skip354w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range353w(i);
	END GENERATE loop94;
	wire_w_lg_write_skip437w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range399w(0);
	loop95 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_write_skip502w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range501w(i);
	END GENERATE loop95;
	wire_w_lg_write_skip394w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range393w(0);
	loop96 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_write_skip528w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range527w(i);
	END GENERATE loop96;
	wire_w_lg_write_state219w(0) <= write_state AND wire_w_lg_w_lg_w_lg_header_proc159w217w218w(0);
	wire_w_lg_write_state243w(0) <= write_state AND wire_w_lg_dprio_pulse198w(0);
	wire_w_lg_write_state777w(0) <= write_state AND wire_w_lg_reconf_done_reg_out697w(0);
	wire_w_lg_write_state786w(0) <= write_state AND wire_w_lg_write_mif_word_done291w(0);
	wire_w_lg_write_state693w(0) <= write_state AND dprio_wr_done;
	wire_w_lg_write_word_done1046w(0) <= write_word_done AND write_happened;
	wire_w_lg_w_channel_address_out_range1092w1093w(0) <= wire_w_channel_address_out_range1092w(0) AND wire_w_lg_is_central_pcs89w(0);
	wire_w_lg_w_tx_pll_sel_wire_range361w370w(0) <= wire_w_tx_pll_sel_wire_range361w(0) AND wire_w_tx_pll_sel_wire_range369w(0);
	wire_w_lg_w_lg_w_lg_is_mif_header280w281w282w(0) <= NOT wire_w_lg_w_lg_is_mif_header280w281w(0);
	wire_w_lg_w894w896w(0) <= NOT wire_w894w(0);
	wire_w_lg_w656w657w(0) <= NOT wire_w656w(0);
	wire_w_lg_bonded_skip228w(0) <= NOT bonded_skip;
	wire_w_lg_cal_busy60w(0) <= NOT cal_busy;
	wire_w_lg_clr_offset823w(0) <= NOT clr_offset;
	wire_w_lg_dprio_pulse198w(0) <= NOT dprio_pulse;
	wire_w_lg_header_proc159w(0) <= NOT header_proc;
	wire_w_lg_idle_state278w(0) <= NOT idle_state;
	wire_w_lg_is_analog_control154w(0) <= NOT is_analog_control;
	wire_w_lg_is_bonded_global_clk_div5w(0) <= NOT is_bonded_global_clk_div;
	wire_w_lg_is_bonded_reconfig13w(0) <= NOT is_bonded_reconfig;
	wire_w_lg_is_cent_clk_div911w(0) <= NOT is_cent_clk_div;
	wire_w_lg_is_central_pcs89w(0) <= NOT is_central_pcs;
	wire_w_lg_is_channel_reconfig408w(0) <= NOT is_channel_reconfig;
	wire_w_lg_is_cruclk_addr0230w(0) <= NOT is_cruclk_addr0;
	wire_w_lg_is_diff_mif167w(0) <= NOT is_diff_mif;
	wire_w_lg_is_end_mif739w(0) <= NOT is_end_mif;
	wire_w_lg_is_global_clk_div_mode226w(0) <= NOT is_global_clk_div_mode;
	wire_w_lg_is_illegal_reg_d220w(0) <= NOT is_illegal_reg_d;
	wire_w_lg_is_mif_stage790w(0) <= NOT is_mif_stage;
	wire_w_lg_is_pll_address77w(0) <= NOT is_pll_address;
	wire_w_lg_is_pll_reconfig420w(0) <= NOT is_pll_reconfig;
	wire_w_lg_is_pll_reset_stage996w(0) <= NOT is_pll_reset_stage;
	wire_w_lg_is_protected_bit227w(0) <= NOT is_protected_bit;
	wire_w_lg_is_rcxpat_chnl_en_ch231w(0) <= NOT is_rcxpat_chnl_en_ch;
	wire_w_lg_is_rx_pcs850w(0) <= NOT is_rx_pcs;
	wire_w_lg_is_rx_pma864w(0) <= NOT is_rx_pma;
	wire_w_lg_is_table_339w(0) <= NOT is_table_33;
	wire_w_lg_is_table_60535w(0) <= NOT is_table_60;
	wire_w_lg_is_table_61899w(0) <= NOT is_table_61;
	wire_w_lg_is_tier_1185w(0) <= NOT is_tier_1;
	wire_w_lg_is_tx_local_div_ctrl1066w(0) <= NOT is_tx_local_div_ctrl;
	wire_w_lg_is_tx_pcs846w(0) <= NOT is_tx_pcs;
	wire_w_lg_is_tx_pma855w(0) <= NOT is_tx_pma;
	wire_w_lg_load_mif_header829w(0) <= NOT load_mif_header;
	wire_w_lg_mif_reconfig_done698w(0) <= NOT mif_reconfig_done;
	wire_w_lg_mif_rx_only969w(0) <= NOT mif_rx_only;
	wire_w_lg_rd_pulse114w(0) <= NOT rd_pulse;
	wire_w_lg_read_state176w(0) <= NOT read_state;
	wire_w_lg_reconf_done_reg_out697w(0) <= NOT reconf_done_reg_out;
	wire_w_lg_reset_reconf_addr216w(0) <= NOT reset_reconf_addr;
	wire_w_lg_reset_system776w(0) <= NOT reset_system;
	wire_w_lg_rx_reconfig617w(0) <= NOT rx_reconfig;
	wire_w_lg_s0_to_040w(0) <= NOT s0_to_0;
	wire_w_lg_s0_to_141w(0) <= NOT s0_to_1;
	wire_w_lg_s2_to_042w(0) <= NOT s2_to_0;
	wire_w_lg_tx_reconfig615w(0) <= NOT tx_reconfig;
	wire_w_lg_wr_pulse115w(0) <= NOT wr_pulse;
	wire_w_lg_write_done221w(0) <= NOT write_done;
	wire_w_lg_write_mif_word_done291w(0) <= NOT write_mif_word_done;
	wire_w_lg_write_skip229w(0) <= NOT write_skip;
	wire_w_lg_write_state796w(0) <= NOT write_state;
	wire_w_lg_w_reconfig_mode_sel_range50w55w(0) <= NOT wire_w_reconfig_mode_sel_range50w(0);
	wire_w_lg_w_reconfig_mode_sel_range51w52w(0) <= NOT wire_w_reconfig_mode_sel_range51w(0);
	wire_w_lg_w_tx_pll_sel_wire_range361w377w(0) <= NOT wire_w_tx_pll_sel_wire_range361w(0);
	wire_w382w(0) <= wire_w_lg_w_lg_w_lg_w_lg_write_skip229w379w380w381w(0) OR wire_w_lg_w_lg_write_skip375w376w(0);
	loop97 : FOR i IN 0 TO 12 GENERATE 
		wire_w429w(i) <= wire_w_lg_w_lg_w_lg_w_lg_write_skip229w426w427w428w(i) OR wire_w_lg_w_lg_w_lg_write_skip422w423w424w(i);
	END GENERATE loop97;
	wire_w417w(0) <= wire_w_lg_w_lg_w_lg_w_lg_write_skip229w414w415w416w(0) OR wire_w_lg_w_lg_w_lg_write_skip410w411w412w(0);
	wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w372w373w(0) <= wire_w_lg_w_lg_w_lg_write_skip229w362w372w(0) OR wire_w_lg_w_lg_write_skip359w367w(0);
	wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w372w401w(0) <= wire_w_lg_w_lg_w_lg_write_skip229w362w372w(0) OR wire_w_lg_w_lg_write_skip359w400w(0);
	wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w363w364w(0) <= wire_w_lg_w_lg_w_lg_write_skip229w362w363w(0) OR wire_w_lg_w_lg_write_skip359w360w(0);
	wire_w_lg_w_lg_w_lg_is_mif_header797w798w799w(0) <= wire_w_lg_w_lg_is_mif_header797w798w(0) OR wire_w_lg_is_end_mif795w(0);
	loop98 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch595w596w597w(i) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch595w596w(i) OR wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch231w593w594w(i);
	END GENERATE loop98;
	wire_w_lg_w_lg_w_lg_is_table_60550w581w582w(0) <= wire_w_lg_w_lg_is_table_60550w581w(0) OR wire_w_lg_w_lg_w_lg_is_table_60535w536w578w(0);
	wire_w_lg_w_lg_w_lg_is_table_60550w565w566w(0) <= wire_w_lg_w_lg_is_table_60550w565w(0) OR wire_w_lg_w_lg_w_lg_is_table_60535w536w557w(0);
	wire_w_lg_w_lg_w_lg_is_table_60550w551w552w(0) <= wire_w_lg_w_lg_is_table_60550w551w(0) OR wire_w_lg_w_lg_w_lg_is_table_60535w536w537w(0);
	wire_w_lg_w_lg_w_lg_is_table_60550w573w574w(0) <= wire_w_lg_w_lg_is_table_60550w573w(0) OR wire_w_lg_w_lg_w_lg_is_table_60535w536w570w(0);
	wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div5w6w7w(0) <= wire_w_lg_w_lg_is_bonded_global_clk_div5w6w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w1062w1063w(0) <= wire_w_lg_w_lg_is_cruclk_addr0230w1062w(0) OR is_tx_local_div_ctrl;
	wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w892w893w(0) <= wire_w_lg_w_lg_is_cruclk_addr0230w892w(0) OR is_cmu;
	wire_w_lg_w_lg_w_lg_is_table_339w10w11w(0) <= wire_w_lg_w_lg_is_table_339w10w(0) OR wire_w_lg_is_table_338w(0);
	wire_w_lg_w_lg_w_lg_mif_rx_only969w970w971w(0) <= wire_w_lg_w_lg_mif_rx_only969w970w(0) OR wire_w_lg_mif_rx_only968w(0);
	wire_w_lg_w_lg_w_lg_write_skip229w342w343w(0) <= wire_w_lg_w_lg_write_skip229w342w(0) OR wire_w_lg_write_skip339w(0);
	wire_w_lg_w_lg_w_lg_write_skip229w328w329w(0) <= wire_w_lg_w_lg_write_skip229w328w(0) OR wire_w_lg_write_skip320w(0);
	wire_w_lg_w_lg_w_lg_write_skip229w315w316w(0) <= wire_w_lg_w_lg_write_skip229w315w(0) OR wire_w_lg_write_skip303w(0);
	wire_w_lg_w_lg_w_lg_write_skip229w335w336w(0) <= wire_w_lg_w_lg_write_skip229w335w(0) OR wire_w_lg_write_skip332w(0);
	wire_w_lg_w_lg_w_lg_write_skip229w602w603w(0) <= wire_w_lg_w_lg_write_skip229w602w(0) OR wire_w_lg_write_skip601w(0);
	loop99 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w460w461w(i) <= wire_w_lg_w_lg_write_skip229w460w(i) OR wire_w_lg_write_skip458w(i);
	END GENERATE loop99;
	loop100 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w587w588w(i) <= wire_w_lg_w_lg_write_skip229w587w(i) OR wire_w_lg_write_skip585w(i);
	END GENERATE loop100;
	loop101 : FOR i IN 0 TO 5 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w348w349w(i) <= wire_w_lg_w_lg_write_skip229w348w(i) OR wire_w_lg_write_skip346w(i);
	END GENERATE loop101;
	loop102 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w387w388w(i) <= wire_w_lg_w_lg_write_skip229w387w(i) OR wire_w_lg_write_skip385w(i);
	END GENERATE loop102;
	loop103 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w479w480w(i) <= wire_w_lg_w_lg_write_skip229w479w(i) OR wire_w_lg_write_skip477w(i);
	END GENERATE loop103;
	loop104 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w452w453w(i) <= wire_w_lg_w_lg_write_skip229w452w(i) OR wire_w_lg_write_skip450w(i);
	END GENERATE loop104;
	loop105 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w468w469w(i) <= wire_w_lg_w_lg_write_skip229w468w(i) OR wire_w_lg_write_skip466w(i);
	END GENERATE loop105;
	loop106 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w485w486w(i) <= wire_w_lg_w_lg_write_skip229w485w(i) OR wire_w_lg_write_skip483w(i);
	END GENERATE loop106;
	wire_w_lg_w_lg_w_lg_write_skip229w444w445w(0) <= wire_w_lg_w_lg_write_skip229w444w(0) OR wire_w_lg_write_skip303w(0);
	loop107 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w495w496w(i) <= wire_w_lg_w_lg_write_skip229w495w(i) OR wire_w_lg_write_skip493w(i);
	END GENERATE loop107;
	loop108 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w513w514w(i) <= wire_w_lg_w_lg_write_skip229w513w(i) OR wire_w_lg_write_skip511w(i);
	END GENERATE loop108;
	loop109 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w405w406w(i) <= wire_w_lg_w_lg_write_skip229w405w(i) OR wire_w_lg_write_skip404w(i);
	END GENERATE loop109;
	loop110 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w356w357w(i) <= wire_w_lg_w_lg_write_skip229w356w(i) OR wire_w_lg_write_skip354w(i);
	END GENERATE loop110;
	wire_w_lg_w_lg_w_lg_write_skip229w439w440w(0) <= wire_w_lg_w_lg_write_skip229w439w(0) OR wire_w_lg_write_skip437w(0);
	loop111 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w504w505w(i) <= wire_w_lg_w_lg_write_skip229w504w(i) OR wire_w_lg_write_skip502w(i);
	END GENERATE loop111;
	wire_w_lg_w_lg_w_lg_write_skip229w396w397w(0) <= wire_w_lg_w_lg_write_skip229w396w(0) OR wire_w_lg_write_skip394w(0);
	loop112 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip229w530w531w(i) <= wire_w_lg_w_lg_write_skip229w530w(i) OR wire_w_lg_write_skip528w(i);
	END GENERATE loop112;
	wire_w_lg_w97w98w(0) <= wire_w97w(0) OR wire_w_lg_is_table_6188w(0);
	wire_w1090w(0) <= wire_w_lg_w_lg_w_lg_is_pma_mif_type1087w1088w1089w(0) OR wire_w_lg_is_table_6188w(0);
	wire_w_lg_w_lg_w_lg_w_channel_address_range93w94w95w96w(0) <= wire_w_lg_w_lg_w_channel_address_range93w94w95w(0) OR wire_w_lg_w_lg_w_logical_pll_sel_num_range90w91w92w(0);
	wire_w_lg_w_lg_w_lg_w_channel_address_range78w79w80w81w(0) <= wire_w_lg_w_lg_w_channel_address_range78w79w80w(0) OR wire_w_lg_w_lg_w_logical_pll_sel_num_range74w75w76w(0);
	loop113 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_cal_busy62w63w(i) <= wire_w_lg_cal_busy62w(i) OR wire_w_lg_w_lg_cal_busy60w61w(i);
	END GENERATE loop113;
	wire_w_lg_w_lg_cal_busy101w102w(0) <= wire_w_lg_cal_busy101w(0) OR wire_w_lg_w_lg_cal_busy60w99w(0);
	wire_w_lg_w_lg_cal_busy85w86w(0) <= wire_w_lg_cal_busy85w(0) OR wire_w_lg_w_lg_cal_busy60w83w(0);
	wire_w_lg_w_lg_cal_busy70w71w(0) <= wire_w_lg_cal_busy70w(0) OR wire_w_lg_w_lg_cal_busy60w68w(0);
	loop114 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain_vodctrl1027w1028w(i) <= wire_w_lg_dprio_datain_vodctrl1027w(i) OR wire_w_lg_dprio_datain_preemp1t1025w(i);
	END GENERATE loop114;
	wire_w_lg_w_lg_is_channel_reconfig842w843w(0) <= wire_w_lg_is_channel_reconfig842w(0) OR is_diff_mif;
	wire_w_lg_w_lg_is_pll_reconfig861w862w(0) <= wire_w_lg_is_pll_reconfig861w(0) OR is_global_clk_div_mode;
	wire_w_lg_w_lg_is_pll_reconfig721w722w(0) <= wire_w_lg_is_pll_reconfig721w(0) OR is_global_clk_div_mode;
	wire_w_lg_w_lg_is_rx_mif_type1083w1084w(0) <= wire_w_lg_is_rx_mif_type1083w(0) OR wire_w_lg_is_cmu912w(0);
	loop115 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_is_table_61904w905w(i) <= wire_w_lg_is_table_61904w(i) OR wire_w_lg_w_lg_is_table_61899w903w(i);
	END GENERATE loop115;
	loop116 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_read_address156w157w(i) <= wire_w_lg_read_address156w(i) OR wire_w_lg_w_lg_is_analog_control154w155w(i);
	END GENERATE loop116;
	loop117 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_write_address162w163w(i) <= wire_w_lg_write_address162w(i) OR wire_w_lg_w_lg_write_reconfig_addr160w161w(i);
	END GENERATE loop117;
	wire_w1094w(0) <= wire_w_lg_w_channel_address_out_range1092w1093w(0) OR wire_w_lg_is_table_6188w(0);
	wire_w_lg_w_lg_w_tx_pll_sel_wire_range361w370w371w(0) <= wire_w_lg_w_tx_pll_sel_wire_range361w370w(0) OR wire_w_tx_pll_sel_wire_range368w(0);
	wire_w_lg_w_lg_is_bonded_reconfig13w20w(0) <= wire_w_lg_is_bonded_reconfig13w(0) OR wire_w_lg_is_bonded_reconfig19w(0);
	wire_w_lg_w_lg_is_bonded_reconfig13w378w(0) <= wire_w_lg_is_bonded_reconfig13w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_is_table_339w886w(0) <= wire_w_lg_is_table_339w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_is_table_339w706w(0) <= wire_w_lg_is_table_339w(0) OR is_pll_reconfig;
	wire_w_lg_w_lg_is_tier_1185w240w(0) <= wire_w_lg_is_tier_1185w(0) OR wire_w_lg_w_lg_is_tier_1237w239w(0);
	wire_w_lg_w_lg_is_tier_1185w215w(0) <= wire_w_lg_is_tier_1185w(0) OR wire_w_lg_is_tier_1214w(0);
	wire_w_lg_w_lg_w_lg_w_lg_is_mif_header797w798w799w800w(0) <= wire_w_lg_w_lg_w_lg_is_mif_header797w798w799w(0) OR wire_w_lg_is_tier_1185w(0);
	loop118 : FOR i IN 0 TO 1 GENERATE 
		wire_w598w(i) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch595w596w597w(i) OR wire_w_lg_write_skip591w(i);
	END GENERATE loop118;
	wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w581w582w583w(0) <= wire_w_lg_w_lg_w_lg_is_table_60550w581w582w(0) OR wire_w_lg_write_skip339w(0);
	wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w565w566w567w(0) <= wire_w_lg_w_lg_w_lg_is_table_60550w565w566w(0) OR wire_w_lg_write_skip320w(0);
	wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w551w552w553w(0) <= wire_w_lg_w_lg_w_lg_is_table_60550w551w552w(0) OR wire_w_lg_write_skip303w(0);
	wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w573w574w575w(0) <= wire_w_lg_w_lg_w_lg_is_table_60550w573w574w(0) OR wire_w_lg_write_skip332w(0);
	wire_w894w(0) <= wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w892w893w(0) OR is_central_pcs;
	wire_w82w(0) <= wire_w_lg_w_lg_w_lg_w_channel_address_range78w79w80w81w(0) OR is_central_pcs;
	loop119 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl1027w1028w1029w(i) <= wire_w_lg_w_lg_dprio_datain_vodctrl1027w1028w(i) OR wire_w_lg_dprio_datain_64_671022w(i);
	END GENERATE loop119;
	wire_w_lg_w_lg_w_lg_is_pll_reconfig861w862w863w(0) <= wire_w_lg_w_lg_is_pll_reconfig861w862w(0) OR is_diff_mif;
	wire_w_lg_w_lg_w_lg_is_pll_reconfig721w722w723w(0) <= wire_w_lg_w_lg_is_pll_reconfig721w722w(0) OR is_central_pcs;
	wire_w_lg_w_lg_w_lg_is_table_339w706w707w(0) <= wire_w_lg_w_lg_is_table_339w706w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_w_lg_is_table_339w706w876w(0) <= wire_w_lg_w_lg_is_table_339w706w(0) OR is_global_clk_div_mode;
	loop120 : FOR i IN 0 TO 15 GENERATE 
		wire_w1030w(i) <= wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl1027w1028w1029w(i) OR wire_w_lg_w_lg_dprio_datain_68_6B1020w1021w(i);
	END GENERATE loop120;
	wire_w_lg_w_lg_w_lg_w_lg_is_table_339w706w876w877w(0) <= wire_w_lg_w_lg_w_lg_is_table_339w706w876w(0) OR is_bonded_global_clk_div;
	loop121 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w1030w1031w(i) <= wire_w1030w(i) OR wire_w_lg_dprio_datain_7c_7f1019w(i);
	END GENERATE loop121;
	loop122 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w1030w1031w1032w(i) <= wire_w_lg_w1030w1031w(i) OR wire_w_lg_dprio_datain_7c_7f_inv1018w(i);
	END GENERATE loop122;
	wire_w656w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w650w651w652w653w654w655w(0) OR is_pll_reset_stage;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w650w651w652w653w654w655w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w650w651w652w653w654w(0) OR is_tx_local_div_ctrl;
	wire_w_lg_w_lg_w_lg_w_lg_w650w651w652w653w654w(0) <= wire_w_lg_w_lg_w_lg_w650w651w652w653w(0) OR is_cruclk_addr0;
	wire_w_lg_w_lg_w_lg_w650w651w652w653w(0) <= wire_w_lg_w_lg_w650w651w652w(0) OR is_table_47;
	wire_w_lg_w_lg_w650w651w652w(0) <= wire_w_lg_w650w651w(0) OR is_table_46;
	wire_w_lg_w650w651w(0) <= wire_w650w(0) OR is_table_44;
	wire_w650w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w644w645w646w647w648w649w(0) OR is_table_43;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w644w645w646w647w648w649w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w644w645w646w647w648w(0) OR is_table_42;
	wire_w_lg_w_lg_w_lg_w_lg_w644w645w646w647w648w(0) <= wire_w_lg_w_lg_w_lg_w644w645w646w647w(0) OR is_table_38;
	wire_w_lg_w_lg_w_lg_w644w645w646w647w(0) <= wire_w_lg_w_lg_w644w645w646w(0) OR is_table_37;
	wire_w_lg_w_lg_w644w645w646w(0) <= wire_w_lg_w644w645w(0) OR is_table_77;
	wire_w_lg_w_lg_w181w182w183w(0) <= wire_w_lg_w181w182w(0) OR is_cent_clk_div;
	wire_w_lg_w644w645w(0) <= wire_w644w(0) OR is_table_76;
	wire_w_lg_w181w182w(0) <= wire_w181w(0) OR is_protected_bit;
	wire_w_lg_w212w213w(0) <= wire_w212w(0) OR is_global_clk_div_mode;
	wire_w644w(0) <= wire_w_lg_w_lg_w_lg_w_lg_is_table_33625w641w642w643w(0) OR is_table_75;
	wire_w195w(0) <= wire_w_lg_w_lg_w_lg_is_cruclk_addr0192w193w194w(0) OR is_cent_clk_div;
	wire_w181w(0) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w180w(0) OR bonded_skip;
	wire_w212w(0) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w211w(0) OR is_protected_bit;
	wire_w_lg_w_lg_w_lg_w_lg_is_table_33625w641w642w643w(0) <= wire_w_lg_w_lg_w_lg_is_table_33625w641w642w(0) OR is_table_61;
	wire_w_lg_w_lg_w_lg_is_cruclk_addr0192w193w194w(0) <= wire_w_lg_w_lg_is_cruclk_addr0192w193w(0) OR is_protected_bit;
	wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w180w(0) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w(0) OR wire_w_lg_is_mif_header177w(0);
	wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w211w(0) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w(0) OR bonded_skip;
	wire_w_lg_w_lg_w_lg_is_table_33625w641w642w(0) <= wire_w_lg_w_lg_is_table_33625w641w(0) OR is_global_clk_div_mode;
	wire_w_lg_w_lg_w_lg_is_tx_pcs606w607w608w(0) <= wire_w_lg_w_lg_is_tx_pcs606w607w(0) OR is_rx_pma;
	wire_w_lg_w_lg_clr_offset881w882w(0) <= wire_w_lg_clr_offset881w(0) OR global_register_reset;
	wire_w_lg_w_lg_delay_mif_head_out1042w1043w(0) <= wire_w_lg_delay_mif_head_out1042w(0) OR write_mif_word_done;
	wire_w_lg_w_lg_is_adce30w31w(0) <= wire_w_lg_is_adce30w(0) OR is_do_dfe;
	wire_w_lg_w_lg_is_cruclk_addr01074w1075w(0) <= wire_w_lg_is_cruclk_addr01074w(0) OR is_tx_local_div_ctrl;
	wire_w_lg_w_lg_is_cruclk_addr0192w193w(0) <= wire_w_lg_is_cruclk_addr0192w(0) OR bonded_skip;
	wire_w_lg_w_lg_is_pll_address66w67w(0) <= wire_w_lg_is_pll_address66w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_is_pma_mif_type1087w1088w(0) <= wire_w_lg_is_pma_mif_type1087w(0) OR is_cmu;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch178w179w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch178w(0) OR write_skip;
	wire_w_lg_w_lg_is_rx_pma920w921w(0) <= wire_w_lg_is_rx_pma920w(0) OR is_central_pcs;
	wire_w_lg_w_lg_is_table_33625w641w(0) <= wire_w_lg_is_table_33625w(0) OR is_table_59;
	wire_w_lg_w_lg_is_tier_11015w1016w(0) <= wire_w_lg_is_tier_11015w(0) OR is_tx_local_div_ctrl;
	wire_w_lg_w_lg_is_tx_pcs606w607w(0) <= wire_w_lg_is_tx_pcs606w(0) OR is_tx_pma;
	wire_w_lg_w_lg_load_mif_header819w820w(0) <= wire_w_lg_load_mif_header819w(0) OR wire_w_lg_is_diff_mif818w(0);
	wire_w_lg_w_lg_write_skip422w423w(0) <= wire_w_lg_write_skip422w(0) OR wire_w_lg_is_bonded_reconfig13w(0);
	wire_w_lg_w_lg_write_skip410w411w(0) <= wire_w_lg_write_skip410w(0) OR wire_w_lg_w_lg_is_channel_reconfig408w409w(0);
	wire_w_lg_w_lg_write_word_preemp1t_data_valid1023w1024w(0) <= wire_w_lg_write_word_preemp1t_data_valid1023w(0) OR write_word_preemp1tb_data_valid;
	wire_w_lg_clr_offset881w(0) <= clr_offset OR is_mif_header;
	wire_w_lg_delay_mif_head_out197w(0) <= delay_mif_head_out OR wire_w_lg_delay_second_mif_head_out196w(0);
	wire_w_lg_delay_mif_head_out1042w(0) <= delay_mif_head_out OR delay_second_mif_head_out;
	wire_w_lg_diff_mif_wr_rd_busy612w(0) <= diff_mif_wr_rd_busy OR diff_mif_reconfig_addr_ready;
	loop123 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_68_6B1020w(i) <= dprio_datain_68_6B(i) OR local_ch_dec;
	END GENERATE loop123;
	wire_w_lg_dprio_pulse188w(0) <= dprio_pulse OR wire_w_lg_diff_mif_reconfig_addr_ready187w(0);
	wire_w_lg_is_adce30w(0) <= is_adce OR is_do_eyemon;
	wire_w_lg_is_channel_reconfig413w(0) <= is_channel_reconfig OR is_global_clk_div_mode;
	wire_w_lg_is_cruclk_addr01069w(0) <= is_cruclk_addr0 OR wire_w_lg_w_lg_is_cruclk_addr0230w1068w(0);
	wire_w_lg_is_cruclk_addr01074w(0) <= is_cruclk_addr0 OR wire_w_lg_w_lg_is_cruclk_addr0230w1073w(0);
	wire_w_lg_is_cruclk_addr0192w(0) <= is_cruclk_addr0 OR write_skip;
	wire_w_lg_is_mif_header280w(0) <= is_mif_header OR mif_reconfig_done;
	wire_w_lg_is_mif_stage792w(0) <= is_mif_stage OR wire_w_lg_idle_state791w(0);
	wire_w_lg_is_pll_address66w(0) <= is_pll_address OR is_central_pcs;
	wire_w_lg_is_pll_reconfig425w(0) <= is_pll_reconfig OR is_global_clk_div_mode;
	wire_w_lg_is_pma_mif_type1087w(0) <= is_pma_mif_type OR is_tx_local_div_ctrl;
	wire_w_lg_is_rcxpat_chnl_en_ch178w(0) <= is_rcxpat_chnl_en_ch OR is_cruclk_addr0;
	wire_w_lg_is_rx_pma920w(0) <= is_rx_pma OR is_cmu;
	wire_w_lg_is_table_33625w(0) <= is_table_33 OR is_table_35;
	wire_w_lg_is_table_351061w(0) <= is_table_35 OR wire_w_dprio_addr_index_range1060w(0);
	wire_w_lg_is_table_59670w(0) <= is_table_59 OR is_global_clk_div_mode;
	wire_w_lg_is_tier_11015w(0) <= is_tier_1 OR is_tier_2;
	wire_w_lg_is_tx_local_div_ctrl639w(0) <= is_tx_local_div_ctrl OR is_pll_reset_stage;
	wire_w_lg_is_tx_pcs606w(0) <= is_tx_pcs OR is_rx_pcs;
	wire_w_lg_load_mif_header819w(0) <= load_mif_header OR clr_offset;
	wire_w_lg_reset_system207w(0) <= reset_system OR wire_w_lg_is_tier_1175w(0);
	wire_w_lg_write_skip422w(0) <= write_skip OR wire_w_lg_w_lg_is_pll_reconfig420w421w(0);
	wire_w_lg_write_skip375w(0) <= write_skip OR wire_w_lg_is_bonded_reconfig19w(0);
	wire_w_lg_write_skip410w(0) <= write_skip OR wire_w_lg_is_bonded_reconfig13w(0);
	wire_w_lg_write_skip359w(0) <= write_skip OR is_bonded_reconfig;
	wire_w_lg_write_word_preemp1t_data_valid1023w(0) <= write_word_preemp1t_data_valid OR write_word_preemp1ta_data_valid;
	wire_w_lg_write_word_vodctrl_data_valid1026w(0) <= write_word_vodctrl_data_valid OR write_word_vodctrla_data_valid;
	wire_w_lg_w_channel_address_range93w94w(0) <= wire_w_channel_address_range93w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_channel_address_range78w79w(0) <= wire_w_channel_address_range78w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_channel_address_out_range1096w1097w(0) <= wire_w_channel_address_out_range1096w(0) OR wire_w_lg_is_central_pcs900w(0);
	wire_w_lg_w_logical_pll_sel_num_range90w91w(0) <= wire_w_logical_pll_sel_num_range90w(0) OR wire_w_lg_is_table_5973w(0);
	wire_w_lg_w_logical_pll_sel_num_range74w75w(0) <= wire_w_logical_pll_sel_num_range74w(0) OR wire_w_lg_is_table_5973w(0);
	wire_w_lg_w_reconfig_mode_sel_range51w58w(0) <= wire_w_reconfig_mode_sel_range51w(0) OR wire_w57w(0);
	a2gr_dprio_addr <= (wire_w_lg_w_lg_w_lg_write_address162w163w164w OR wire_w_lg_w_lg_w_lg_read_address156w157w158w);
	a2gr_dprio_data <= wire_w_lg_w_lg_dprio_datain1013w1014w;
	a2gr_dprio_rden <= (rd_pulse AND (wire_w_lg_is_diff_mif167w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	a2gr_dprio_wren <= ((wire_w_lg_wr_pulse1010w(0) AND wire_w_lg_is_analog_control154w(0)) AND (wire_w_lg_is_diff_mif167w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	a2gr_dprio_wren_data <= (wire_w_lg_wr_pulse1008w(0) AND (wire_w_lg_is_diff_mif167w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	adce_busy_state <= '0';
	adce_state <= '0';
	add_sub_datab <= ((((wire_w_lg_is_rx_pma915w OR wire_w_lg_w_lg_w_lg_is_cmu912w913w914w) OR wire_w_lg_w_lg_w_lg_is_cmu908w909w910w) OR wire_w_lg_is_global_clk_div_mode907w) OR wire_w_lg_is_central_pcs906w);
	add_sub_sel <= (NOT (is_rx_pma OR wire_w_lg_is_central_pcs900w(0)));
	aeq_ch_done <= (OTHERS => '0');
	bonded_skip <= ((((((wire_w_lg_is_table_33625w(0) AND is_bonded_reconfig) OR is_table_59) OR is_table_61) OR is_table_75) OR is_table_76) OR is_table_77);
	busy <= (((wire_w_lg_w_lg_is_bonded_reconfig13w14w(0) OR wire_w_lg_is_bonded_reconfig12w(0)) OR internal_write_pulse) OR cal_busy);
	busy_state <= ((((read_state OR write_state) OR adce_state) OR eyemon_busy) OR dfe_busy);
	cal_busy <= wire_calibration_busy;
	cal_channel_address <= wire_calibration_dprio_addr(14 DOWNTO 12);
	cal_channel_address_out <= address_pres_reg(2 DOWNTO 0);
	cal_dprio_address <= ( wire_calibration_dprio_addr(15) & cal_channel_address_out & wire_calibration_dprio_addr(11 DOWNTO 0));
	cal_dprioout_wire(0) <= ( reconfig_fromgxb(0));
	cal_quad_address <= wire_calibration_quad_addr;
	cal_testbuses <= ( reconfig_fromgxb(4 DOWNTO 1));
	cent_clk_div_plus_one <= "00001";
	central_pcs_first_word_addr <= wire_central_pcs_first_word_mux_result;
	central_pcs_max <= "00101";
	central_pcs_minus_one <= "00001";
	central_pcs_plus_seven <= "00111";
	channel_address <= (OTHERS => '0');
	channel_address_out <= wire_address_pres_reg_w_lg_w_q_range111w112w;
	channel_reconfig_done <= reconf_done_reg_out;
	clr_offset <= (((is_offset_end AND en_mif_addr_cntr) AND wire_w_lg_is_diff_mif167w(0)) OR (diff_mif_clr_offset AND is_diff_mif));
	cmu_max <= "00101";
	cmu_pll_plus_three <= "00011";
	cruclk_mux_data <= ( wire_w_lg_w_lg_w_lg_write_skip229w315w316w & wire_w_lg_w_lg_w_lg_write_skip229w328w329w & wire_w_lg_w_lg_w_lg_write_skip229w335w336w & wire_w_lg_w_lg_w_lg_write_skip229w342w343w & wire_w_lg_w_lg_w_lg_write_skip229w348w349w & dprio_dataout_reg(5 DOWNTO 4) & wire_w_lg_w_lg_w_lg_write_skip229w356w357w);
	delay_mif_head_out <= delay_mif_head;
	delay_second_mif_head_out <= delay_second_mif_head;
	dfe_busy <= '0';
	diff_mif_address_busy <= '0';
	diff_mif_clr_offset <= '0';
	diff_mif_load_mif_header <= '0';
	diff_mif_mif_header <= (OTHERS => '0');
	diff_mif_reconfig_addr_load <= '0';
	diff_mif_reconfig_addr_ready <= '0';
	diff_mif_reconfig_addr_start <= '0';
	diff_mif_reconfig_address <= (OTHERS => '0');
	diff_mif_wr_rd_busy <= '0';
	dprio_addr_index <= (wire_w_lg_w_lg_w894w896w897w OR wire_w_lg_w894w895w);
	dprio_addr_offset_cmpr_datab <= wire_central_pcs_global_clk_div_mux_result;
	dprio_addr_offset_cnt_out <= wire_dprio_addr_offset_cnt_q;
	dprio_addr_translated_offset <= wire_add_sub11_w_lg_result922w;
	dprio_datain <= (wire_w_lg_w_lg_w_lg_w1030w1031w1032w1033w OR wire_w_lg_w_lg_w_lg_is_tier_11015w1016w1017w);
	dprio_datain_64_67 <= (OTHERS => '0');
	dprio_datain_68_6B <= (OTHERS => '0');
	dprio_datain_7c_7f <= (OTHERS => '0');
	dprio_datain_7c_7f_inv <= (OTHERS => '0');
	dprio_datain_preemp1t <= (OTHERS => '0');
	dprio_datain_vodctrl <= (OTHERS => '0');
	dprio_pulse <= ((dprio_pulse_reg XOR wire_dprio_busy) AND wire_dprio_w_lg_busy170w(0));
	dprio_wr_done <= wire_dprio_status_out(1);
	duplex_pma_first_pll <= "010110";
	duplex_pma_pcs_first_pll <= "110001";
	en_mif_addr_cntr <= ((read_state AND dprio_wr_done) OR wire_w_lg_w_lg_write_state693w694w(0));
	en_write_trigger <= legal_wr_mode_type;
	eyemon_busy <= '0';
	global_clk_div_addr <= wire_add_sub12_result;
	global_clk_div_addr_offset <= "000100";
	global_clk_div_mode_offset_max <= (OTHERS => '0');
	global_clk_div_mode_plus_five <= "00101";
	global_register_reset <= global_register_reset_reg;
	header_proc <= ((((delay_mif_head OR is_mif_header) OR delay_second_mif_head_out) OR is_second_mif_header) AND is_tier_1);
	idle_state <= (NOT state_mc_reg(0));
	internal_write_pulse <= '0';
	is_adce <= ((((is_adce_single_control OR is_adce_all_control) OR is_adce_continuous_single_control) OR is_adce_one_time_single_control) OR is_adce_standby_single_control);
	is_adce_all_control <= '0';
	is_adce_continuous_single_control <= '0';
	is_adce_one_time_single_control <= '0';
	is_adce_single_control <= '0';
	is_adce_standby_single_control <= '0';
	is_analog_control <= wire_reconf_mode_dec_eq(0);
	is_bonded_global_clk_div <= is_bonded_global_clk_div_reg;
	is_bonded_reconfig <= is_bonded_reconfig_reg;
	is_cent_clk_div <= ((is_table_59 OR is_table_60) OR is_global_clk_div_mode);
	is_central_pcs <= wire_reconf_mode_dec_eq(7);
	is_channel_reconfig <= ((wire_reconf_mode_dec_eq(1) OR wire_reconf_mode_dec_eq(5)) OR wire_reconf_mode_dec_eq(6));
	is_cmu <= ((((wire_mif_type_reg_w_lg_w_q_range865w866w(0) AND wire_w_lg_is_rx_pcs850w(0)) AND wire_w_lg_is_tx_pma855w(0)) AND wire_w_lg_is_rx_pma864w(0)) AND wire_w_lg_w_lg_w_lg_is_pll_reconfig861w862w863w(0));
	is_cruclk_addr0 <= ((wire_is_cru_idx0_aeb AND is_tier_1) AND is_rx_pma);
	is_diff_mif <= '0';
	is_do_dfe <= '0';
	is_do_eyemon <= '0';
	is_end_mif <= end_mif_reg;
	is_global_clk_div_mode <= wire_reconf_mode_dec_eq(2);
	is_illegal_reg_d <= '0';
	is_illegal_reg_out <= '0';
	is_mif_header <= wire_is_special_address_aeb;
	is_mif_stage <= mif_stage;
	is_offset_end <= wire_dprio_addr_offset_cmpr_aeb;
	is_pll_address <= is_cmu;
	is_pll_end_mif <= '0';
	is_pll_first_word <= '0';
	is_pll_reconfig <= (wire_reconf_mode_dec_eq(4) OR wire_reconf_mode_dec_eq(5));
	is_pll_reset_stage <= '0';
	is_pma_mif_type <= (is_tx_pma OR is_rx_pma);
	is_protected_bit <= (((((((is_table_35 OR is_table_37) OR is_table_38) OR is_table_42) OR is_table_43) OR is_table_44) OR is_table_46) OR is_table_47);
	is_rcxpat_chnl_en_ch <= ((wire_is_rcxpat_chnl_en_ch_word_aeb AND is_tier_1) AND is_tx_pcs);
	is_rx_mif_type <= (is_rx_pcs OR is_rx_pma);
	is_rx_pcs <= (wire_mif_type_reg_w_lg_w_q_range847w848w(0) AND wire_w_lg_w_lg_is_channel_reconfig842w843w(0));
	is_rx_pma <= (((wire_mif_type_reg_w_lg_w_q_range856w857w(0) AND wire_w_lg_is_rx_pcs850w(0)) AND wire_w_lg_is_tx_pma855w(0)) AND wire_w_lg_w_lg_is_channel_reconfig842w843w(0));
	is_second_mif_header <= wire_is_second_mif_header_address_aeb;
	is_table_33 <= ((wire_is_table_33_idx_aeb AND is_tier_1) AND is_tx_pma);
	is_table_35 <= (wire_is_table_35_cmp_aeb AND is_tx_pma);
	is_table_37 <= ((wire_is_table_37_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_38 <= ((wire_is_table_38_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_42 <= ((wire_is_table_42_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_43 <= ((wire_is_table_43_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_44 <= ((wire_is_table_44_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_46 <= ((wire_is_table_46_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_47 <= ((wire_is_table_47_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_59 <= ((wire_is_table_59_idx_aeb AND is_tier_1) AND is_cmu);
	is_table_60 <= ((wire_is_table_60_idx_aeb AND is_tier_1) AND is_cmu);
	is_table_61 <= ((wire_is_table_61_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_table_75 <= ((wire_is_table_75_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_table_76 <= ((wire_is_table_76_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_table_77 <= ((wire_is_table_77_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_tier_1 <= (((((wire_reconf_mode_dec_eq(1) OR wire_reconf_mode_dec_eq(6)) OR wire_reconf_mode_dec_eq(4)) OR wire_reconf_mode_dec_eq(5)) OR wire_reconf_mode_dec_eq(7)) OR is_global_clk_div_mode);
	is_tier_2 <= '0';
	is_tx_local_div_ctrl <= wire_reconf_mode_dec_eq(3);
	is_tx_pcs <= wire_mif_type_reg_w_lg_w_q_range844w845w(0);
	is_tx_pma <= ((wire_mif_type_reg_w_lg_w_q_range851w852w(0) AND wire_w_lg_is_rx_pcs850w(0)) AND wire_w_lg_w_lg_is_channel_reconfig842w843w(0));
	legal_wr_mode_type <= (wire_w_lg_w_reconfig_mode_sel_range51w58w(0) OR ((wire_w_lg_w_reconfig_mode_sel_range51w52w(0) AND reconfig_mode_sel(0)) AND (NOT reconfig_mode_sel(1))));
	load_mif_header <= wire_w_lg_w_lg_is_mif_header292w293w(0);
	local_ch_dec <= aeq_ch_done(0);
	logical_pll_sel_num <= ( "0" & logical_pll_num_reg);
	merged_dprioin <= ( wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w551w552w553w & wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w565w566w567w & wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w573w574w575w & wire_w_lg_w_lg_w_lg_w_lg_is_table_60550w581w582w583w & wire_w_lg_w_lg_w_lg_write_skip229w587w588w & wire_w598w & wire_w_lg_w_lg_w_lg_write_skip229w602w603w);
	mif_addr_cntr_data <= wire_mif_addr_cntr_data_mux_result;
	mif_reconfig_done <= ((wire_mif_type_reg_w_lg_w_lg_w984w985w986w(0) AND wire_w_lg_is_central_pcs89w(0)) OR wire_w_lg_w_lg_is_central_pcs977w978w(0));
	mif_rx_only <= ((NOT mif_type_reg(2)) AND (NOT mif_type_reg(4)));
	offset_cancellation_reset <= '0';
	pll_first_word_addr <= wire_pll_first_word_mux_result;
	quad_address <= (OTHERS => '0');
	quad_address_out <= address_pres_reg(11 DOWNTO 3);
	rd_pulse <= ((((wire_w_lg_dprio_pulse198w(0) AND wire_w_lg_write_done221w(0)) AND wire_wr_rd_pulse_reg_w_lg_q173w(0)) AND wire_w_lg_is_illegal_reg_d220w(0)) AND wire_w_lg_write_state219w(0));
	read_address <= (OTHERS => '0');
	read_reconfig_addr <= (OTHERS => '0');
	read_state <= '0';
	reconf_done_reg_out <= reconfig_done_reg;
	reconfig_address_en <= (((write_done OR idle_state) AND (NOT (wire_w_lg_is_pll_reset_stage996w(0) AND is_pll_first_word))) AND (NOT (is_pll_reset_stage AND is_pll_end_mif)));
	reconfig_address_out <= wire_mif_addr_cntr_w_lg_w_lg_q741w742w;
	reconfig_datain <= ((((((((((((((((wire_w_lg_is_cruclk_addr0674w OR wire_w_lg_is_table_33673w) OR wire_w_lg_is_table_35672w) OR wire_w_lg_w_lg_is_table_59670w671w) OR wire_w_lg_is_table_61669w) OR wire_w_lg_is_table_75668w) OR wire_w_lg_is_table_76667w) OR wire_w_lg_is_table_77666w) OR wire_w_lg_is_table_37665w) OR wire_w_lg_is_table_38664w) OR wire_w_lg_is_table_42663w) OR wire_w_lg_is_table_43662w) OR wire_w_lg_is_table_44661w) OR wire_w_lg_is_table_46660w) OR wire_w_lg_is_table_47659w) OR wire_w_lg_merged_dprioin658w) OR wire_w_lg_w_lg_is_tx_local_div_ctrl639w640w);
	reconfig_reset_all <= '0';
	reconfig_togxb <= ( wire_calibration_busy & wire_dprio_dprioload & wire_dprio_dpriodisable & wire_dprio_dprioin);
	reset_addr_done <= '0';
	reset_reconf_addr <= '0';
	reset_system <= '0';
	rx_pcs_max <= "10110";
	rx_pma_max <= "01100";
	rx_pma_minus_one <= "00001";
	rx_reconfig <= '1';
	s0_to_0 <= write_done;
	s0_to_1 <= (write_all_int AND idle_state);
	s0_to_2 <= (wire_w_lg_idle_state32w(0) AND (wire_w_lg_write_all21w(0) OR (is_bonded_reconfig AND is_bonded_global_clk_div)));
	s2_to_0 <= (adce_state AND (NOT ((adce_busy_state OR eyemon_busy) OR dfe_busy)));
	start <= '0';
	state_mc_reg_in(0) <= ((s0_to_2 OR s0_to_1) OR (((wire_w_lg_s2_to_042w(0) AND wire_w_lg_s0_to_141w(0)) AND wire_w_lg_s0_to_040w(0)) AND state_mc_reg(0)));
	table_33_data <= ( wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w363w364w & wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w372w373w & wire_w382w & wire_w_lg_w_lg_w_lg_write_skip229w387w388w);
	table_35_data <= ( dprio_dataout_reg(15 DOWNTO 5) & wire_w_lg_w_lg_w_lg_write_skip229w396w397w & wire_w_lg_w_lg_w_lg_w_lg_write_skip229w362w372w401w & wire_w_lg_w_lg_w_lg_write_skip229w405w406w);
	table_37_data <= ( wire_w_lg_w_lg_w_lg_write_skip229w485w486w & dprio_dataout_reg(11 DOWNTO 3) & wire_w_lg_w_lg_w_lg_write_skip229w405w406w);
	table_38_data <= ( wire_w_lg_w_lg_w_lg_write_skip229w495w496w & dprio_dataout_reg(6 DOWNTO 5) & wire_w_lg_w_lg_w_lg_write_skip229w504w505w);
	table_42_data <= ( dprio_dataout_reg(15 DOWNTO 0));
	table_43_data <= ( wire_w_lg_w_lg_w_lg_write_skip229w513w514w & dprio_dataout_reg(7 DOWNTO 0));
	table_44_data <= ( wire_w_lg_w_lg_w_lg_write_skip229w444w445w & dprio_dataout_reg(14 DOWNTO 4) & wire_w_lg_w_lg_w_lg_write_skip229w356w357w);
	table_46_data <= ( dprio_dataout_reg(15 DOWNTO 10) & wire_w_lg_w_lg_w_lg_write_skip229w530w531w);
	table_47_data <= ( dprio_dataout_reg(15 DOWNTO 0));
	table_59_data <= ( dprio_dataout_reg(15 DOWNTO 14) & wire_w417w & wire_w429w);
	table_61_data <= ( dprio_dataout_reg(15 DOWNTO 4) & wire_w_lg_w_lg_w_lg_write_skip229w439w440w & dprio_dataout_reg(2 DOWNTO 0));
	table_75_data <= ( wire_w_lg_w_lg_w_lg_write_skip229w444w445w & dprio_dataout_reg(14) & wire_w_lg_w_lg_w_lg_write_skip229w452w453w & dprio_dataout_reg(11) & wire_w_lg_w_lg_w_lg_write_skip229w460w461w);
	table_76_data <= ( dprio_dataout_reg(15) & wire_w_lg_w_lg_w_lg_write_skip229w468w469w & dprio_dataout_reg(5 DOWNTO 3) & wire_w_lg_w_lg_w_lg_write_skip229w405w406w);
	table_77_data <= ( dprio_dataout_reg(15 DOWNTO 14) & wire_w_lg_w_lg_w_lg_write_skip229w479w480w);
	transceiver_init <= '0';
	tx_pcs_max <= "00011";
	tx_pll_sel_wire <= tx_cmu_sel;
	tx_pma_first_pll <= "001001";
	tx_pma_max <= "00110";
	tx_pma_pcs_first_pll <= "001101";
	tx_reconfig <= '1';
	wr_pulse <= (((wire_w_lg_write_state243w(0) AND wire_w_lg_write_done221w(0)) AND (wire_wr_rd_pulse_reg_w_lg_q241w(0) OR (wire_w_lg_is_tier_1237w(0) AND (((((wire_w_lg_is_rcxpat_chnl_en_ch231w(0) AND wire_w_lg_is_cruclk_addr0230w(0)) AND wire_w_lg_write_skip229w(0)) AND wire_w_lg_bonded_skip228w(0)) AND wire_w_lg_is_protected_bit227w(0)) AND wire_w_lg_is_global_clk_div_mode226w(0))))) AND wire_w_lg_is_illegal_reg_d220w(0));
	write_address <= ( "0" & address_pres_reg(2) & channel_address_out & "11" & "000000" & "0000");
	write_all_int <= ((wire_w_lg_write_all21w(0) OR (is_bonded_reconfig AND is_bonded_global_clk_div)) AND en_write_trigger);
	write_done <= ((((wire_w_lg_w_lg_write_word_done1046w1047w(0) OR ((wire_w_lg_w_lg_delay_mif_head_out1042w1043w(0) OR (is_diff_mif AND is_end_mif)) OR (reset_addr_done AND is_tier_1))) OR ((dprio_pulse AND write_happened) AND (is_tier_2 OR is_tx_local_div_ctrl))) OR (is_illegal_reg_out AND write_state)) OR reset_system);
	write_happened <= wr_addr_inc_reg;
	write_mif_word_done <= ((dprio_pulse AND write_happened) AND is_tier_1);
	write_reconfig_addr <= ( "0" & address_pres_reg(2) & wire_w_lg_w_channel_address_out_range1096w1097w & wire_w1094w & wire_w1090w & wire_w_lg_w_lg_w_lg_is_rx_mif_type1083w1084w1085w & "00000" & wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w1078w1079w & wire_w_lg_w_lg_is_cruclk_addr01074w1075w & wire_w_lg_w_lg_is_cruclk_addr01069w1070w & wire_w_lg_w_lg_w_lg_is_cruclk_addr0230w1062w1063w);
	write_skip <= (((((is_tx_pcs OR is_tx_pma) AND wire_w_lg_tx_reconfig615w(0)) OR ((is_rx_pcs OR is_rx_pma) AND wire_w_lg_rx_reconfig617w(0))) OR wire_w_lg_is_cmu616w(0)) OR (wire_w_lg_is_diff_mif613w(0) AND (wire_w_lg_w_lg_w_lg_is_pll_reconfig420w421w610w(0) OR (wire_w_lg_is_channel_reconfig408w(0) AND wire_w_lg_w_lg_w_lg_is_tx_pcs606w607w608w(0)))));
	write_state <= state_mc_reg(0);
	write_word_64_67_data_valid <= '0';
	write_word_68_6B_data_valid <= '0';
	write_word_7c_7f_data_valid <= '0';
	write_word_7c_7f_inv_data_valid <= '0';
	write_word_done <= '0';
	write_word_preemp1t_data_valid <= '0';
	write_word_preemp1ta_data_valid <= '0';
	write_word_preemp1tb_data_valid <= '0';
	write_word_vodctrl_data_valid <= '0';
	write_word_vodctrla_data_valid <= '0';
	wire_w_cal_channel_address_range100w(0) <= cal_channel_address(0);
	wire_w_cal_channel_address_range84w(0) <= cal_channel_address(1);
	wire_w_cal_channel_address_range69w(0) <= cal_channel_address(2);
	wire_w_channel_address_range93w(0) <= channel_address(0);
	wire_w_channel_address_range78w(0) <= channel_address(1);
	wire_w_channel_address_out_range1092w(0) <= channel_address_out(0);
	wire_w_channel_address_out_range1096w(0) <= channel_address_out(1);
	wire_w_dprio_addr_index_range1060w(0) <= dprio_addr_index(0);
	wire_w_dprio_addr_index_range1067w(0) <= dprio_addr_index(1);
	wire_w_dprio_addr_index_range1072w(0) <= dprio_addr_index(2);
	wire_w_dprio_addr_index_range1077w <= dprio_addr_index(4 DOWNTO 3);
	wire_w_logical_pll_sel_num_range90w(0) <= logical_pll_sel_num(0);
	wire_w_logical_pll_sel_num_range74w(0) <= logical_pll_sel_num(1);
	wire_w_reconfig_mode_sel_range50w(0) <= reconfig_mode_sel(0);
	wire_w_reconfig_mode_sel_range48w(0) <= reconfig_mode_sel(1);
	wire_w_reconfig_mode_sel_range51w(0) <= reconfig_mode_sel(2);
	wire_w_tx_pll_sel_wire_range369w(0) <= tx_pll_sel_wire(0);
	wire_w_tx_pll_sel_wire_range361w(0) <= tx_pll_sel_wire(1);
	wire_w_tx_pll_sel_wire_range368w(0) <= tx_pll_sel_wire(2);
	loop124 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy138w142w(i) <= wire_calibration_w_lg_busy138w(0) AND a2gr_dprio_addr(i);
	END GENERATE loop124;
	loop125 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy138w139w(i) <= wire_calibration_w_lg_busy138w(0) AND a2gr_dprio_data(i);
	END GENERATE loop125;
	wire_calibration_w_lg_w_lg_busy138w145w(0) <= wire_calibration_w_lg_busy138w(0) AND a2gr_dprio_rden;
	wire_calibration_w_lg_w_lg_busy138w148w(0) <= wire_calibration_w_lg_busy138w(0) AND a2gr_dprio_wren;
	wire_calibration_w_lg_w_lg_busy138w151w(0) <= wire_calibration_w_lg_busy138w(0) AND a2gr_dprio_wren_data;
	loop126 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_busy143w(i) <= wire_calibration_busy AND cal_dprio_address(i);
	END GENERATE loop126;
	loop127 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_busy140w(i) <= wire_calibration_busy AND wire_calibration_dprio_dataout(i);
	END GENERATE loop127;
	wire_calibration_w_lg_busy138w(0) <= NOT wire_calibration_busy;
	wire_calibration_reset <= wire_w_lg_offset_cancellation_reset123w(0);
	wire_w_lg_offset_cancellation_reset123w(0) <= offset_cancellation_reset OR reconfig_reset_all;
	calibration :  alt_cal
	  GENERIC MAP (
		CHANNEL_ADDRESS_WIDTH => 0,
		NUMBER_OF_CHANNELS => 1,
		SIM_MODEL_MODE => "FALSE"
	  )
	  PORT MAP ( 
		busy => wire_calibration_busy,
		clock => reconfig_clk,
		dprio_addr => wire_calibration_dprio_addr,
		dprio_busy => wire_dprio_busy,
		dprio_datain => wire_dprio_dataout,
		dprio_dataout => wire_calibration_dprio_dataout,
		dprio_rden => wire_calibration_dprio_rden,
		dprio_wren => wire_calibration_dprio_wren,
		quad_addr => wire_calibration_quad_addr,
		remap_addr => address_pres_reg,
		reset => wire_calibration_reset,
		retain_addr => wire_calibration_retain_addr,
		start => start,
		testbuses => cal_testbuses,
		transceiver_init => transceiver_init
	  );
	wire_dprio_w_lg_w_lg_w_status_out_range691w729w730w(0) <= wire_dprio_w_lg_w_status_out_range691w729w(0) AND reset_system;
	wire_dprio_w_lg_busy170w(0) <= NOT wire_dprio_busy;
	wire_dprio_w_lg_w_status_out_range691w729w(0) <= wire_dprio_w_status_out_range691w(0) OR wire_dprio_w_status_out_range728w(0);
	wire_dprio_address <= wire_calibration_w_lg_w_lg_busy143w144w;
	loop128 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy143w144w(i) <= wire_calibration_w_lg_busy143w(i) OR wire_calibration_w_lg_w_lg_busy138w142w(i);
	END GENERATE loop128;
	wire_dprio_datain <= wire_calibration_w_lg_w_lg_busy140w141w;
	loop129 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy140w141w(i) <= wire_calibration_w_lg_busy140w(i) OR wire_calibration_w_lg_w_lg_busy138w139w(i);
	END GENERATE loop129;
	wire_dprio_rden <= wire_calibration_w_lg_w_lg_busy146w147w(0);
	wire_calibration_w_lg_w_lg_busy146w147w(0) <= (wire_calibration_busy AND wire_calibration_dprio_rden) OR wire_calibration_w_lg_w_lg_busy138w145w(0);
	wire_dprio_wren <= wire_calibration_w_lg_w_lg_busy149w150w(0);
	wire_calibration_w_lg_w_lg_busy149w150w(0) <= (wire_calibration_busy AND wire_calibration_dprio_wren) OR wire_calibration_w_lg_w_lg_busy138w148w(0);
	wire_dprio_wren_data <= wire_calibration_w_lg_w_lg_busy152w153w(0);
	wire_calibration_w_lg_w_lg_busy152w153w(0) <= (wire_calibration_busy AND wire_calibration_retain_addr) OR wire_calibration_w_lg_w_lg_busy138w151w(0);
	wire_dprio_w_status_out_range691w(0) <= wire_dprio_status_out(1);
	wire_dprio_w_status_out_range728w(0) <= wire_dprio_status_out(3);
	dprio :  altgx_reconfig_cpri_alt_dprio_t2l
	  PORT MAP ( 
		address => wire_dprio_address,
		busy => wire_dprio_busy,
		datain => wire_dprio_datain,
		dataout => wire_dprio_dataout,
		dpclk => reconfig_clk,
		dpriodisable => wire_dprio_dpriodisable,
		dprioin => wire_dprio_dprioin,
		dprioload => wire_dprio_dprioload,
		dprioout => cal_dprioout_wire(0),
		quad_address => quad_address_out,
		rden => wire_dprio_rden,
		reset => reconfig_reset_all,
		status_out => wire_dprio_status_out,
		wren => wire_dprio_wren,
		wren_data => wire_dprio_wren_data
	  );
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN address_pres_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN address_pres_reg <= ( wire_w_lg_w_lg_cal_busy62w63w & wire_w_lg_w_lg_cal_busy70w71w & wire_w_lg_w_lg_cal_busy85w86w & wire_w_lg_w_lg_cal_busy101w102w);
		END IF;
	END PROCESS;
	wire_address_pres_reg_w_lg_w_lg_w_q_range107w108w109w(0) <= wire_address_pres_reg_w_lg_w_q_range107w108w(0) AND wire_address_pres_reg_w_q_range105w(0);
	loop130 : FOR i IN 0 TO 1 GENERATE 
		wire_address_pres_reg_w_lg_w_q_range111w112w(i) <= wire_address_pres_reg_w_q_range111w(i) AND wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range107w108w109w110w(0);
	END GENERATE loop130;
	wire_address_pres_reg_w_lg_w_q_range107w108w(0) <= wire_address_pres_reg_w_q_range107w(0) AND wire_address_pres_reg_w_q_range106w(0);
	wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range107w108w109w110w(0) <= NOT wire_address_pres_reg_w_lg_w_lg_w_q_range107w108w109w(0);
	wire_address_pres_reg_w_q_range105w(0) <= address_pres_reg(0);
	wire_address_pres_reg_w_q_range111w <= address_pres_reg(1 DOWNTO 0);
	wire_address_pres_reg_w_q_range106w(0) <= address_pres_reg(1);
	wire_address_pres_reg_w_q_range107w(0) <= address_pres_reg(2);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN cru_num_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (load_mif_header = '1') THEN cru_num_reg <= wire_reconfig_data_reg_w_q_range294w;
			END IF;
		END IF;
	END PROCESS;
	wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range309w323w324w325w(0) <= wire_cru_num_reg_w_lg_w_lg_w_q_range309w323w324w(0) AND wire_cru_num_reg_w_q_range304w(0);
	wire_cru_num_reg_w_lg_w_lg_w_q_range306w307w321w(0) <= wire_cru_num_reg_w_lg_w_q_range306w307w(0) AND wire_cru_num_reg_w_lg_w_q_range304w310w(0);
	wire_cru_num_reg_w_lg_w_lg_w_q_range306w307w308w(0) <= wire_cru_num_reg_w_lg_w_q_range306w307w(0) AND wire_cru_num_reg_w_q_range304w(0);
	wire_cru_num_reg_w_lg_w_lg_w_q_range305w311w312w(0) <= wire_cru_num_reg_w_lg_w_q_range305w311w(0) AND wire_cru_num_reg_w_lg_w_q_range304w310w(0);
	wire_cru_num_reg_w_lg_w_lg_w_q_range305w311w340w(0) <= wire_cru_num_reg_w_lg_w_q_range305w311w(0) AND wire_cru_num_reg_w_q_range304w(0);
	wire_cru_num_reg_w_lg_w_lg_w_q_range309w323w324w(0) <= wire_cru_num_reg_w_lg_w_q_range309w323w(0) AND wire_cru_num_reg_w_lg_w_q_range306w322w(0);
	wire_cru_num_reg_w_lg_w_q_range306w307w(0) <= wire_cru_num_reg_w_q_range306w(0) AND wire_cru_num_reg_w_q_range305w(0);
	wire_cru_num_reg_w_lg_w_q_range304w310w(0) <= NOT wire_cru_num_reg_w_q_range304w(0);
	wire_cru_num_reg_w_lg_w_q_range305w311w(0) <= NOT wire_cru_num_reg_w_q_range305w(0);
	wire_cru_num_reg_w_lg_w_q_range306w322w(0) <= NOT wire_cru_num_reg_w_q_range306w(0);
	wire_cru_num_reg_w_lg_w_q_range309w323w(0) <= NOT wire_cru_num_reg_w_q_range309w(0);
	wire_cru_num_reg_w_lg_w_lg_w_lg_w_lg_w_q_range309w323w324w325w326w(0) <= wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range309w323w324w325w(0) OR wire_cru_num_reg_w_q_range309w(0);
	wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range305w311w312w313w(0) <= wire_cru_num_reg_w_lg_w_lg_w_q_range305w311w312w(0) OR wire_cru_num_reg_w_q_range309w(0);
	wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range305w311w340w341w(0) <= wire_cru_num_reg_w_lg_w_lg_w_q_range305w311w340w(0) OR wire_cru_num_reg_w_lg_w_q_range306w307w(0);
	wire_cru_num_reg_w327w(0) <= wire_cru_num_reg_w_lg_w_lg_w_lg_w_lg_w_q_range309w323w324w325w326w(0) OR wire_cru_num_reg_w_lg_w_lg_w_q_range306w307w321w(0);
	wire_cru_num_reg_w_lg_w_lg_w_lg_w_lg_w_q_range305w311w312w313w314w(0) <= wire_cru_num_reg_w_lg_w_lg_w_lg_w_q_range305w311w312w313w(0) OR wire_cru_num_reg_w_lg_w_lg_w_q_range306w307w308w(0);
	wire_cru_num_reg_w_lg_w_lg_w_q_range309w333w334w(0) <= wire_cru_num_reg_w_lg_w_q_range309w333w(0) OR wire_cru_num_reg_w_q_range305w(0);
	wire_cru_num_reg_w_lg_w_q_range309w333w(0) <= wire_cru_num_reg_w_q_range309w(0) OR wire_cru_num_reg_w_q_range306w(0);
	wire_cru_num_reg_w_q_range304w(0) <= cru_num_reg(0);
	wire_cru_num_reg_w_q_range305w(0) <= cru_num_reg(1);
	wire_cru_num_reg_w_q_range306w(0) <= cru_num_reg(2);
	wire_cru_num_reg_w_q_range309w(0) <= cru_num_reg(3);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN delay_mif_head <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_delay_mif_head_ena = '1') THEN delay_mif_head <= (is_mif_header AND is_tier_1);
			END IF;
		END IF;
	END PROCESS;
	wire_delay_mif_head_ena <= (((wire_w_lg_write_state777w(0) AND wire_w_lg_write_mif_word_done291w(0)) AND wire_w_lg_reset_reconf_addr216w(0)) AND wire_w_lg_reset_system776w(0));
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN delay_second_mif_head <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_delay_second_mif_head_ena = '1') THEN delay_second_mif_head <= wire_w_lg_is_second_mif_header724w(0);
			END IF;
		END IF;
	END PROCESS;
	wire_delay_second_mif_head_ena <= (((wire_w_lg_write_state786w(0) AND wire_w_lg_reset_reconf_addr216w(0)) AND wire_w_lg_reset_system776w(0)) AND is_tier_1);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(0) = '1') THEN dprio_dataout_reg(0) <= wire_dprio_dataout_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(1) = '1') THEN dprio_dataout_reg(1) <= wire_dprio_dataout_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(2) = '1') THEN dprio_dataout_reg(2) <= wire_dprio_dataout_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(3) = '1') THEN dprio_dataout_reg(3) <= wire_dprio_dataout_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(4) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(4) = '1') THEN dprio_dataout_reg(4) <= wire_dprio_dataout_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(5) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(5) = '1') THEN dprio_dataout_reg(5) <= wire_dprio_dataout_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(6) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(6) = '1') THEN dprio_dataout_reg(6) <= wire_dprio_dataout_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(7) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(7) = '1') THEN dprio_dataout_reg(7) <= wire_dprio_dataout_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(8) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(8) = '1') THEN dprio_dataout_reg(8) <= wire_dprio_dataout_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(9) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(9) = '1') THEN dprio_dataout_reg(9) <= wire_dprio_dataout_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(10) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(10) = '1') THEN dprio_dataout_reg(10) <= wire_dprio_dataout_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(11) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(11) = '1') THEN dprio_dataout_reg(11) <= wire_dprio_dataout_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(12) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(12) = '1') THEN dprio_dataout_reg(12) <= wire_dprio_dataout_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(13) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(13) = '1') THEN dprio_dataout_reg(13) <= wire_dprio_dataout_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(14) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(14) = '1') THEN dprio_dataout_reg(14) <= wire_dprio_dataout_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg(15) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_dataout_reg_ena(15) = '1') THEN dprio_dataout_reg(15) <= wire_dprio_dataout_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	wire_dprio_dataout_reg_d <= ( wire_dprio_dataout(15 DOWNTO 0));
	loop131 : FOR i IN 0 TO 15 GENERATE
		wire_dprio_dataout_reg_ena(i) <= wire_w_lg_dprio_pulse279w(0);
	END GENERATE loop131;
	wire_dprio_dataout_reg_w_q_range457w <= dprio_dataout_reg(10 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range489w <= dprio_dataout_reg(11 DOWNTO 3);
	wire_dprio_dataout_reg_w_q_range345w <= dprio_dataout_reg(11 DOWNTO 6);
	wire_dprio_dataout_reg_w_q_range384w <= dprio_dataout_reg(12 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range338w(0) <= dprio_dataout_reg(12);
	wire_dprio_dataout_reg_w_q_range476w <= dprio_dataout_reg(13 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range449w <= dprio_dataout_reg(13 DOWNTO 12);
	wire_dprio_dataout_reg_w_q_range331w(0) <= dprio_dataout_reg(13);
	wire_dprio_dataout_reg_w_q_range319w(0) <= dprio_dataout_reg(14);
	wire_dprio_dataout_reg_w_q_range465w <= dprio_dataout_reg(14 DOWNTO 6);
	wire_dprio_dataout_reg_w_q_range482w <= dprio_dataout_reg(15 DOWNTO 12);
	wire_dprio_dataout_reg_w_q_range302w(0) <= dprio_dataout_reg(15);
	wire_dprio_dataout_reg_w_q_range492w <= dprio_dataout_reg(15 DOWNTO 7);
	wire_dprio_dataout_reg_w_q_range510w <= dprio_dataout_reg(15 DOWNTO 8);
	wire_dprio_dataout_reg_w_q_range403w <= dprio_dataout_reg(2 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range590w <= dprio_dataout_reg(2 DOWNTO 1);
	wire_dprio_dataout_reg_w_q_range353w <= dprio_dataout_reg(3 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range399w(0) <= dprio_dataout_reg(3);
	wire_dprio_dataout_reg_w_q_range501w <= dprio_dataout_reg(4 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range393w(0) <= dprio_dataout_reg(4);
	wire_dprio_dataout_reg_w_q_range527w <= dprio_dataout_reg(9 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range600w(0) <= dprio_dataout_reg(0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_pulse_reg_ena = '1') THEN dprio_pulse_reg <= wire_dprio_busy;
			END IF;
		END IF;
	END PROCESS;
	wire_dprio_pulse_reg_ena <= (read_state OR write_state);
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (is_tier_1 = '1') THEN end_mif_reg <= mif_reconfig_done;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN global_register_reset_reg <= (((reset_addr_done OR reconfig_reset_all) OR is_illegal_reg_out) OR mif_reconfig_done);
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, global_register_reset)
	BEGIN
		IF (global_register_reset = '1') THEN is_bonded_global_clk_div_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_is_bonded_global_clk_div_reg_ena = '1') THEN is_bonded_global_clk_div_reg <= wire_is_bonded_global_clk_div_reg_w_lg_q812w(0);
			END IF;
		END IF;
	END PROCESS;
	wire_is_bonded_global_clk_div_reg_ena <= ((wire_is_bonded_global_clk_div_reg_w_lg_w_lg_w_lg_w_lg_q812w813w814w815w(0) AND wire_w_lg_is_pll_reconfig420w(0)) AND en_mif_addr_cntr);
	wire_is_bonded_global_clk_div_reg_w_lg_w_lg_q812w813w(0) <= wire_is_bonded_global_clk_div_reg_w_lg_q812w(0) AND is_table_33;
	wire_is_bonded_global_clk_div_reg_w_lg_w_lg_w_lg_w_lg_q812w813w814w815w(0) <= wire_is_bonded_global_clk_div_reg_w_lg_w_lg_w_lg_q812w813w814w(0) AND is_bonded_reconfig;
	wire_is_bonded_global_clk_div_reg_w_lg_q812w(0) <= NOT is_bonded_global_clk_div_reg;
	wire_is_bonded_global_clk_div_reg_w_lg_w_lg_w_lg_q812w813w814w(0) <= wire_is_bonded_global_clk_div_reg_w_lg_w_lg_q812w813w(0) OR is_bonded_global_clk_div_reg;
	PROCESS (reconfig_clk, global_register_reset)
	BEGIN
		IF (global_register_reset = '1') THEN is_bonded_reconfig_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (delay_second_mif_head_out = '1') THEN is_bonded_reconfig_reg <= wire_reconfig_data_reg_w_q_range556w(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN logical_pll_num_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (is_mif_header = '1') THEN logical_pll_num_reg(0) <= ( reconfig_data_reg(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_stage <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (is_tier_1 = '1') THEN 
				IF (wire_mif_stage_sclr = '1') THEN mif_stage <= '0';
				ELSE mif_stage <= ((wire_mif_stage_w_lg_q284w(0) AND wire_w_lg_is_mif_header280w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_is_mif_header280w281w282w283w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_mif_stage_sclr <= ((reset_system OR is_illegal_reg_out) OR mif_reconfig_done);
	wire_mif_stage_w_lg_q284w(0) <= NOT mif_stage;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(0) = '1') THEN 
				IF (wire_mif_type_reg_sclr(0) = '1') THEN mif_type_reg(0) <= '0';
				ELSE mif_type_reg(0) <= wire_mif_type_reg_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(1) = '1') THEN 
				IF (wire_mif_type_reg_sclr(1) = '1') THEN mif_type_reg(1) <= '0';
				ELSE mif_type_reg(1) <= wire_mif_type_reg_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(2) = '1') THEN 
				IF (wire_mif_type_reg_sclr(2) = '1') THEN mif_type_reg(2) <= '0';
				ELSE mif_type_reg(2) <= wire_mif_type_reg_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(3) = '1') THEN 
				IF (wire_mif_type_reg_sclr(3) = '1') THEN mif_type_reg(3) <= '0';
				ELSE mif_type_reg(3) <= wire_mif_type_reg_d(3);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(4) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(4) = '1') THEN 
				IF (wire_mif_type_reg_sclr(4) = '1') THEN mif_type_reg(4) <= '0';
				ELSE mif_type_reg(4) <= wire_mif_type_reg_d(4);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_mif_type_reg_d <= wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_lg_w_q_range824w825w826w827w828w;
	loop132 : FOR i IN 0 TO 4 GENERATE
		wire_mif_type_reg_ena(i) <= wire_w_lg_w_lg_load_mif_header819w820w(0);
	END GENERATE loop132;
	wire_mif_type_reg_sclr <= ( wire_w_lg_w_lg_w_lg_load_mif_header829w830w831w & wire_w_lg_w_lg_w_lg_load_mif_header829w830w834w & wire_w_lg_w_lg_w_lg_load_mif_header829w830w836w & wire_w_lg_w_lg_w_lg_load_mif_header829w830w838w & wire_w_lg_w_lg_w_lg_load_mif_header829w830w840w);
	wire_mif_type_reg_w_lg_w_lg_w984w985w986w(0) <= wire_mif_type_reg_w_lg_w984w985w(0) AND write_done;
	wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range844w980w981w982w983w(0) <= wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range844w980w981w982w(0) AND is_channel_reconfig;
	wire_mif_type_reg_w_lg_w_q_range865w866w(0) <= wire_mif_type_reg_w_q_range865w(0) AND wire_w_lg_is_tx_pcs846w(0);
	wire_mif_type_reg_w_lg_w_q_range865w979w(0) <= wire_mif_type_reg_w_q_range865w(0) AND wire_w_lg_is_pll_reconfig425w(0);
	wire_mif_type_reg_w_lg_w_q_range856w857w(0) <= wire_mif_type_reg_w_q_range856w(0) AND wire_w_lg_is_tx_pcs846w(0);
	wire_mif_type_reg_w_lg_w_q_range851w852w(0) <= wire_mif_type_reg_w_q_range851w(0) AND wire_w_lg_is_tx_pcs846w(0);
	wire_mif_type_reg_w_lg_w_q_range847w848w(0) <= wire_mif_type_reg_w_q_range847w(0) AND wire_w_lg_is_tx_pcs846w(0);
	wire_mif_type_reg_w_lg_w_q_range844w845w(0) <= wire_mif_type_reg_w_q_range844w(0) AND wire_w_lg_w_lg_is_channel_reconfig842w843w(0);
	wire_mif_type_reg_w_lg_w984w985w(0) <= NOT wire_mif_type_reg_w984w(0);
	wire_mif_type_reg_w984w(0) <= wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range844w980w981w982w983w(0) OR wire_mif_type_reg_w_lg_w_q_range865w979w(0);
	wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range844w980w981w982w(0) <= wire_mif_type_reg_w_lg_w_lg_w_q_range844w980w981w(0) OR wire_mif_type_reg_w_q_range856w(0);
	wire_mif_type_reg_w_lg_w_lg_w_q_range844w980w981w(0) <= wire_mif_type_reg_w_lg_w_q_range844w980w(0) OR wire_mif_type_reg_w_q_range851w(0);
	wire_mif_type_reg_w_lg_w_q_range844w980w(0) <= wire_mif_type_reg_w_q_range844w(0) OR wire_mif_type_reg_w_q_range847w(0);
	wire_mif_type_reg_w_q_range865w(0) <= mif_type_reg(0);
	wire_mif_type_reg_w_q_range856w(0) <= mif_type_reg(1);
	wire_mif_type_reg_w_q_range851w(0) <= mif_type_reg(2);
	wire_mif_type_reg_w_q_range847w(0) <= mif_type_reg(3);
	wire_mif_type_reg_w_q_range844w(0) <= mif_type_reg(4);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(0) = '1') THEN reconf_mode_sel_reg(0) <= reconfig_mode_sel(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(1) = '1') THEN reconf_mode_sel_reg(1) <= reconfig_mode_sel(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(2) = '1') THEN reconf_mode_sel_reg(2) <= reconfig_mode_sel(2);
			END IF;
		END IF;
	END PROCESS;
	loop133 : FOR i IN 0 TO 2 GENERATE
		wire_reconf_mode_sel_reg_ena(i) <= wire_w_lg_idle_state290w(0);
	END GENERATE loop133;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(0) = '1') THEN reconfig_data_reg(0) <= reconfig_data(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(1) = '1') THEN reconfig_data_reg(1) <= reconfig_data(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(2) = '1') THEN reconfig_data_reg(2) <= reconfig_data(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(3) = '1') THEN reconfig_data_reg(3) <= reconfig_data(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(4) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(4) = '1') THEN reconfig_data_reg(4) <= reconfig_data(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(5) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(5) = '1') THEN reconfig_data_reg(5) <= reconfig_data(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(6) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(6) = '1') THEN reconfig_data_reg(6) <= reconfig_data(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(7) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(7) = '1') THEN reconfig_data_reg(7) <= reconfig_data(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(8) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(8) = '1') THEN reconfig_data_reg(8) <= reconfig_data(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(9) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(9) = '1') THEN reconfig_data_reg(9) <= reconfig_data(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(10) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(10) = '1') THEN reconfig_data_reg(10) <= reconfig_data(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(11) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(11) = '1') THEN reconfig_data_reg(11) <= reconfig_data(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(12) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(12) = '1') THEN reconfig_data_reg(12) <= reconfig_data(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(13) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(13) = '1') THEN reconfig_data_reg(13) <= reconfig_data(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(14) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(14) = '1') THEN reconfig_data_reg(14) <= reconfig_data(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(15) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(15) = '1') THEN reconfig_data_reg(15) <= reconfig_data(15);
			END IF;
		END IF;
	END PROCESS;
	loop134 : FOR i IN 0 TO 15 GENERATE
		wire_reconfig_data_reg_ena(i) <= wire_w_lg_idle_state605w(0);
	END GENERATE loop134;
	loop135 : FOR i IN 0 TO 4 GENERATE 
		wire_reconfig_data_reg_w_lg_w_lg_w_q_range824w825w826w(i) <= wire_reconfig_data_reg_w_lg_w_q_range824w825w(i) AND wire_w_lg_clr_offset823w(0);
	END GENERATE loop135;
	loop136 : FOR i IN 0 TO 4 GENERATE 
		wire_reconfig_data_reg_w_lg_w_q_range824w825w(i) <= wire_reconfig_data_reg_w_q_range824w(i) AND load_mif_header;
	END GENERATE loop136;
	loop137 : FOR i IN 0 TO 4 GENERATE 
		wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range824w825w826w827w(i) <= wire_reconfig_data_reg_w_lg_w_lg_w_q_range824w825w826w(i) OR wire_w_lg_clr_offset822w(i);
	END GENERATE loop137;
	loop138 : FOR i IN 0 TO 4 GENERATE 
		wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_lg_w_q_range824w825w826w827w828w(i) <= wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range824w825w826w827w(i) OR wire_w_lg_w_lg_is_diff_mif818w821w(i);
	END GENERATE loop138;
	wire_reconfig_data_reg_w_q_range297w(0) <= reconfig_data_reg(0);
	wire_reconfig_data_reg_w_q_range459w <= reconfig_data_reg(10 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range295w <= reconfig_data_reg(10 DOWNTO 7);
	wire_reconfig_data_reg_w_q_range586w <= reconfig_data_reg(11 DOWNTO 3);
	wire_reconfig_data_reg_w_q_range347w <= reconfig_data_reg(11 DOWNTO 6);
	wire_reconfig_data_reg_w_q_range386w <= reconfig_data_reg(12 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range577w(0) <= reconfig_data_reg(12);
	wire_reconfig_data_reg_w_q_range478w <= reconfig_data_reg(13 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range451w <= reconfig_data_reg(13 DOWNTO 12);
	wire_reconfig_data_reg_w_q_range569w(0) <= reconfig_data_reg(13);
	wire_reconfig_data_reg_w_q_range556w(0) <= reconfig_data_reg(14);
	wire_reconfig_data_reg_w_q_range467w <= reconfig_data_reg(14 DOWNTO 6);
	wire_reconfig_data_reg_w_q_range824w <= reconfig_data_reg(15 DOWNTO 11);
	wire_reconfig_data_reg_w_q_range484w <= reconfig_data_reg(15 DOWNTO 12);
	wire_reconfig_data_reg_w_q_range443w(0) <= reconfig_data_reg(15);
	wire_reconfig_data_reg_w_q_range494w <= reconfig_data_reg(15 DOWNTO 7);
	wire_reconfig_data_reg_w_q_range512w <= reconfig_data_reg(15 DOWNTO 8);
	wire_reconfig_data_reg_w_q_range296w <= reconfig_data_reg(2 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range592w <= reconfig_data_reg(2 DOWNTO 1);
	wire_reconfig_data_reg_w_q_range355w <= reconfig_data_reg(3 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range438w(0) <= reconfig_data_reg(3);
	wire_reconfig_data_reg_w_q_range503w <= reconfig_data_reg(4 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range395w(0) <= reconfig_data_reg(4);
	wire_reconfig_data_reg_w_q_range294w <= reconfig_data_reg(6 DOWNTO 3);
	wire_reconfig_data_reg_w_q_range529w <= reconfig_data_reg(9 DOWNTO 0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_done_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_done_reg_ena = '1') THEN 
				IF (reset_system = '1') THEN reconfig_done_reg <= '0';
				ELSE reconfig_done_reg <= (((wire_w_lg_mif_reconfig_done805w(0) OR (is_diff_mif AND is_end_mif)) AND wire_reconfig_done_reg_w_lg_q802w(0)) OR wire_reconfig_done_reg_w_lg_q801w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_reconfig_done_reg_ena <= ((wire_w_lg_is_mif_stage792w(0) AND wire_w_lg_is_diff_mif167w(0)) OR is_diff_mif);
	wire_reconfig_done_reg_w_lg_q801w(0) <= reconfig_done_reg AND wire_w_lg_w_lg_w_lg_w_lg_is_mif_header797w798w799w800w(0);
	wire_reconfig_done_reg_w_lg_q802w(0) <= NOT reconfig_done_reg;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN state_mc_reg <= state_mc_reg_in;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_cmu_sel <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_le7_out = '1') THEN tx_cmu_sel <= wire_reconfig_data_reg_w_q_range296w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_pll_inclk_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_pll_inclk_reg_ena(0) = '1') THEN tx_pll_inclk_reg(0) <= wire_tx_pll_inclk_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_pll_inclk_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_pll_inclk_reg_ena(1) = '1') THEN tx_pll_inclk_reg(1) <= wire_tx_pll_inclk_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_pll_inclk_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_pll_inclk_reg_ena(2) = '1') THEN tx_pll_inclk_reg(2) <= wire_tx_pll_inclk_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_pll_inclk_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_pll_inclk_reg_ena(3) = '1') THEN tx_pll_inclk_reg(3) <= wire_tx_pll_inclk_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_pll_inclk_reg_d <= wire_reconfig_data_reg_w_q_range295w;
	loop139 : FOR i IN 0 TO 3 GENERATE
		wire_tx_pll_inclk_reg_ena(i) <= wire_w_lg_w_lg_is_mif_header292w293w(0);
	END GENERATE loop139;
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range544w560w561w562w(0) <= wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range544w560w561w(0) AND wire_tx_pll_inclk_reg_w_q_range538w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range540w541w558w(0) <= wire_tx_pll_inclk_reg_w_lg_w_q_range540w541w(0) AND wire_tx_pll_inclk_reg_w_lg_w_q_range538w546w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range540w541w542w(0) <= wire_tx_pll_inclk_reg_w_lg_w_q_range540w541w(0) AND wire_tx_pll_inclk_reg_w_q_range538w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range539w543w547w(0) <= wire_tx_pll_inclk_reg_w_lg_w_q_range539w543w(0) AND wire_tx_pll_inclk_reg_w_lg_w_q_range538w546w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range539w543w579w(0) <= wire_tx_pll_inclk_reg_w_lg_w_q_range539w543w(0) AND wire_tx_pll_inclk_reg_w_q_range538w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range544w560w561w(0) <= wire_tx_pll_inclk_reg_w_lg_w_q_range544w560w(0) AND wire_tx_pll_inclk_reg_w_lg_w_q_range540w559w(0);
	wire_tx_pll_inclk_reg_w_lg_w_q_range540w541w(0) <= wire_tx_pll_inclk_reg_w_q_range540w(0) AND wire_tx_pll_inclk_reg_w_q_range539w(0);
	wire_tx_pll_inclk_reg_w_lg_w_q_range544w545w(0) <= wire_tx_pll_inclk_reg_w_q_range544w(0) AND wire_tx_pll_inclk_reg_w_lg_w_q_range539w543w(0);
	wire_tx_pll_inclk_reg_w_lg_w_q_range538w546w(0) <= NOT wire_tx_pll_inclk_reg_w_q_range538w(0);
	wire_tx_pll_inclk_reg_w_lg_w_q_range539w543w(0) <= NOT wire_tx_pll_inclk_reg_w_q_range539w(0);
	wire_tx_pll_inclk_reg_w_lg_w_q_range540w559w(0) <= NOT wire_tx_pll_inclk_reg_w_q_range540w(0);
	wire_tx_pll_inclk_reg_w_lg_w_q_range544w560w(0) <= NOT wire_tx_pll_inclk_reg_w_q_range544w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_lg_w_q_range544w560w561w562w563w(0) <= wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range544w560w561w562w(0) OR wire_tx_pll_inclk_reg_w_lg_w_q_range544w545w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range539w543w547w548w(0) <= wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range539w543w547w(0) OR wire_tx_pll_inclk_reg_w_lg_w_q_range544w545w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range539w543w579w580w(0) <= wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range539w543w579w(0) OR wire_tx_pll_inclk_reg_w_lg_w_q_range540w541w(0);
	wire_tx_pll_inclk_reg_w564w(0) <= wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_lg_w_q_range544w560w561w562w563w(0) OR wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range540w541w558w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_lg_w_q_range539w543w547w548w549w(0) <= wire_tx_pll_inclk_reg_w_lg_w_lg_w_lg_w_q_range539w543w547w548w(0) OR wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range540w541w542w(0);
	wire_tx_pll_inclk_reg_w_lg_w_lg_w_q_range544w571w572w(0) <= wire_tx_pll_inclk_reg_w_lg_w_q_range544w571w(0) OR wire_tx_pll_inclk_reg_w_q_range539w(0);
	wire_tx_pll_inclk_reg_w_lg_w_q_range544w571w(0) <= wire_tx_pll_inclk_reg_w_q_range544w(0) OR wire_tx_pll_inclk_reg_w_q_range540w(0);
	wire_tx_pll_inclk_reg_w_q_range538w(0) <= tx_pll_inclk_reg(0);
	wire_tx_pll_inclk_reg_w_q_range539w(0) <= tx_pll_inclk_reg(1);
	wire_tx_pll_inclk_reg_w_q_range540w(0) <= tx_pll_inclk_reg(2);
	wire_tx_pll_inclk_reg_w_q_range544w(0) <= tx_pll_inclk_reg(3);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_addr_inc_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN wr_addr_inc_reg <= (wr_pulse OR ((wire_w_lg_wr_pulse115w(0) AND wire_w_lg_rd_pulse114w(0)) AND wr_addr_inc_reg));
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_rd_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wr_rd_pulse_reg_ena = '1') THEN 
				IF (wire_wr_rd_pulse_reg_sclr = '1') THEN wr_rd_pulse_reg <= '0';
				ELSE wr_rd_pulse_reg <= wire_wr_rd_pulse_reg_w_lg_q173w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_wr_rd_pulse_reg_ena <= ((((((((wire_w_lg_dprio_pulse198w(0) AND wire_w_lg_is_diff_mif167w(0)) AND wire_w_lg_delay_mif_head_out197w(0)) OR (is_diff_mif AND diff_mif_reconfig_addr_start)) OR ((wire_w_lg_dprio_pulse188w(0) AND (wire_w_lg_is_tier_1185w(0) OR wire_w_lg_is_tier_1184w(0))) AND wire_w_lg_read_state176w(0))) OR wire_w_lg_is_tier_1175w(0)) OR (is_diff_mif AND write_done)) OR reset_addr_done) OR is_illegal_reg_out);
	wire_wr_rd_pulse_reg_sclr <= (((wire_w_lg_reset_system207w(0) OR (is_diff_mif AND write_done)) OR reset_addr_done) OR is_illegal_reg_out);
	wire_wr_rd_pulse_reg_w_lg_q241w(0) <= wr_rd_pulse_reg AND wire_w_lg_w_lg_is_tier_1185w240w(0);
	wire_wr_rd_pulse_reg_w_lg_q173w(0) <= NOT wr_rd_pulse_reg;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wren_data_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wren_data_reg_ena = '1') THEN wren_data_reg <= (wire_wren_data_reg_w_lg_w_lg_q1003w1004w(0) OR wire_wren_data_reg_w_lg_q1002w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_wren_data_reg_ena <= (is_tier_1 AND (wire_w_lg_is_diff_mif167w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	wire_wren_data_reg_w_lg_w_lg_q1003w1004w(0) <= wire_wren_data_reg_w_lg_q1003w(0) AND rd_pulse;
	wire_wren_data_reg_w_lg_q1002w(0) <= wren_data_reg AND wire_w_lg_write_done221w(0);
	wire_wren_data_reg_w_lg_q1003w(0) <= NOT wren_data_reg;
	wire_wren_data_reg_w_lg_q1007w(0) <= wren_data_reg OR is_analog_control;
	le7 :  lcell
	  PORT MAP ( 
		a_in => is_mif_header,
		a_out => wire_le7_out
	  );
	loop140 : FOR i IN 0 TO 4 GENERATE 
		wire_add_sub11_w_lg_result922w(i) <= wire_add_sub11_result(i) AND wire_w_lg_w_lg_is_rx_pma920w921w(0);
	END GENERATE loop140;
	add_sub11 :  lpm_add_sub
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		add_sub => add_sub_sel,
		dataa => wire_dprio_addr_offset_cnt_q,
		datab => add_sub_datab,
		result => wire_add_sub11_result
	  );
	add_sub12 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		dataa => pll_first_word_addr,
		datab => global_clk_div_addr_offset,
		result => wire_add_sub12_result
	  );
	dprio_addr_offset_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_dprio_addr_offset_cmpr_aeb,
		dataa => wire_dprio_addr_offset_cnt_q,
		datab => dprio_addr_offset_cmpr_datab
	  );
	wire_is_cru_idx0_datab <= (OTHERS => '0');
	is_cru_idx0 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_cru_idx0_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_cru_idx0_datab
	  );
	wire_is_rcxpat_chnl_en_ch_word_datab <= "00001";
	is_rcxpat_chnl_en_ch_word :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_rcxpat_chnl_en_ch_word_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_rcxpat_chnl_en_ch_word_datab
	  );
	wire_is_second_mif_header_address_datab <= "000001";
	is_second_mif_header_address :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_is_second_mif_header_address_aeb,
		dataa => wire_mif_addr_cntr_q,
		datab => wire_is_second_mif_header_address_datab
	  );
	wire_is_special_address_datab <= (OTHERS => '0');
	is_special_address :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_is_special_address_aeb,
		dataa => wire_mif_addr_cntr_q,
		datab => wire_is_special_address_datab
	  );
	wire_is_table_33_idx_datab <= "00101";
	is_table_33_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_33_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_33_idx_datab
	  );
	wire_is_table_35_cmp_datab <= "00110";
	is_table_35_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_35_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_35_cmp_datab
	  );
	wire_is_table_37_cmp_datab <= "00010";
	is_table_37_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_37_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_37_cmp_datab
	  );
	wire_is_table_38_cmp_datab <= "00011";
	is_table_38_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_38_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_38_cmp_datab
	  );
	wire_is_table_42_cmp_datab <= "00111";
	is_table_42_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_42_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_42_cmp_datab
	  );
	wire_is_table_43_cmp_datab <= "01000";
	is_table_43_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_43_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_43_cmp_datab
	  );
	wire_is_table_44_cmp_datab <= "01001";
	is_table_44_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_44_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_44_cmp_datab
	  );
	wire_is_table_46_cmp_datab <= "01011";
	is_table_46_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_46_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_46_cmp_datab
	  );
	wire_is_table_47_cmp_datab <= "01100";
	is_table_47_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_47_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_47_cmp_datab
	  );
	wire_is_table_59_idx_datab <= "00100";
	is_table_59_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_59_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_59_idx_datab
	  );
	wire_is_table_60_idx_datab <= "00101";
	is_table_60_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_60_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_60_idx_datab
	  );
	wire_is_table_61_idx_datab <= (OTHERS => '0');
	is_table_61_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_61_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_61_idx_datab
	  );
	wire_is_table_75_idx_datab <= "00001";
	is_table_75_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_75_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_75_idx_datab
	  );
	wire_is_table_76_idx_datab <= "00010";
	is_table_76_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_76_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_76_idx_datab
	  );
	wire_is_table_77_idx_datab <= "00011";
	is_table_77_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_77_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_77_idx_datab
	  );
	wire_dprio_addr_offset_cnt_cnt_en <= wire_w_lg_w_lg_w_lg_en_mif_addr_cntr710w879w880w(0);
	wire_w_lg_w_lg_w_lg_en_mif_addr_cntr710w879w880w(0) <= (wire_w_lg_en_mif_addr_cntr710w(0) OR ((en_mif_addr_cntr AND is_bonded_reconfig) AND wire_w_lg_w_lg_w_lg_w_lg_is_table_339w706w876w877w(0))) AND wire_w_lg_is_diff_mif167w(0);
	wire_dprio_addr_offset_cnt_data <= wire_w_lg_w_lg_diff_mif_reconfig_address884w885w;
	wire_dprio_addr_offset_cnt_sclr <= wire_w_lg_w_lg_w_lg_clr_offset881w882w883w(0);
	wire_w_lg_w_lg_w_lg_clr_offset881w882w883w(0) <= wire_w_lg_w_lg_clr_offset881w882w(0) OR (is_diff_mif AND write_done);
	wire_dprio_addr_offset_cnt_sload <= wire_w891w(0);
	wire_w891w(0) <= (wire_w_lg_diff_mif_reconfig_addr_load889w(0) OR ((diff_mif_reconfig_addr_load AND is_bonded_reconfig) AND wire_w_lg_w_lg_is_table_339w886w(0))) AND is_diff_mif;
	dprio_addr_offset_cnt :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => wire_dprio_addr_offset_cnt_cnt_en,
		data => wire_dprio_addr_offset_cnt_data,
		q => wire_dprio_addr_offset_cnt_q,
		sclr => wire_dprio_addr_offset_cnt_sclr,
		sload => wire_dprio_addr_offset_cnt_sload
	  );
	loop141 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_w_lg_w_lg_q741w742w(i) <= wire_mif_addr_cntr_w_lg_q741w(i) AND is_tier_1;
	END GENERATE loop141;
	loop142 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_w_lg_q741w(i) <= wire_mif_addr_cntr_q(i) AND wire_w_lg_w_lg_mif_reconfig_done698w740w(0);
	END GENERATE loop142;
	wire_mif_addr_cntr_cnt_en <= wire_w713w(0);
	wire_w713w(0) <= ((wire_w_lg_en_mif_addr_cntr710w(0) OR ((en_mif_addr_cntr AND is_bonded_reconfig) AND wire_w_lg_w_lg_w_lg_is_table_339w706w707w(0))) OR ((((((is_mif_header AND write_state) OR (is_second_mif_header AND write_state)) AND wire_w_lg_write_done221w(0)) AND wire_w_lg_mif_reconfig_done698w(0)) AND wire_w_lg_reconf_done_reg_out697w(0)) AND wire_w_lg_dprio_pulse198w(0))) AND is_tier_1;
	wire_mif_addr_cntr_sclr <= wire_w_lg_w737w738w(0);
	wire_w_lg_w737w738w(0) <= ((((reset_reconf_addr OR is_end_mif) AND (NOT ((is_mif_header OR is_second_mif_header) AND write_state))) OR wire_dprio_w_lg_w_lg_w_status_out_range691w729w730w(0)) OR is_illegal_reg_out) OR reconfig_reset_all;
	wire_mif_addr_cntr_sload <= wire_w727w(0);
	wire_w727w(0) <= (wire_w_lg_w_lg_is_second_mif_header724w725w(0) AND wire_w_lg_w_lg_w_lg_is_pll_reconfig721w722w723w(0)) AND wire_w_lg_is_diff_mif167w(0);
	mif_addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 62,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => wire_mif_addr_cntr_cnt_en,
		data => mif_addr_cntr_data,
		q => wire_mif_addr_cntr_q,
		sclr => wire_mif_addr_cntr_sclr,
		sload => wire_mif_addr_cntr_sload
	  );
	wire_reconf_mode_dec_enable <= wire_w_lg_w_lg_idle_state278w289w(0);
	wire_w_lg_w_lg_idle_state278w289w(0) <= wire_w_lg_idle_state278w(0) OR mif_stage;
	reconf_mode_dec :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => reconf_mode_sel_reg,
		enable => wire_reconf_mode_dec_enable,
		eq => wire_reconf_mode_dec_eq
	  );
	wire_central_pcs_first_word_mux_data <= ( "100110" & "001111" & "110111" & "010011" & "011100" & "001111" & duplex_pma_pcs_first_pll & tx_pma_pcs_first_pll & duplex_pma_first_pll & tx_pma_first_pll);
	wire_central_pcs_first_word_mux_sel <= ( mif_rx_only & mif_type_reg(0) & mif_type_reg(4) & wire_w_lg_w_lg_w_lg_mif_rx_only969w970w971w);
	central_pcs_first_word_mux :  altgx_reconfig_cpri_mux_r7a
	  PORT MAP ( 
		data => wire_central_pcs_first_word_mux_data,
		result => wire_central_pcs_first_word_mux_result,
		sel => wire_central_pcs_first_word_mux_sel
	  );
	wire_central_pcs_global_clk_div_mux_data <= ( global_clk_div_mode_offset_max & central_pcs_max & wire_max_word_per_mif_type_result);
	wire_central_pcs_global_clk_div_mux_sel <= ( is_global_clk_div_mode & is_central_pcs);
	central_pcs_global_clk_div_mux :  altgx_reconfig_cpri_mux_a6a
	  PORT MAP ( 
		data => wire_central_pcs_global_clk_div_mux_data,
		result => wire_central_pcs_global_clk_div_mux_result,
		sel => wire_central_pcs_global_clk_div_mux_sel
	  );
	wire_max_word_per_mif_type_data <= ( cmu_max & rx_pma_max & tx_pma_max & rx_pcs_max & tx_pcs_max);
	wire_max_word_per_mif_type_sel <= ( is_cmu & is_pma_mif_type & is_rx_mif_type);
	max_word_per_mif_type :  altgx_reconfig_cpri_mux_d6a
	  PORT MAP ( 
		data => wire_max_word_per_mif_type_data,
		result => wire_max_word_per_mif_type_result,
		sel => wire_max_word_per_mif_type_sel
	  );
	wire_mif_addr_cntr_data_mux_data <= ( global_clk_div_addr & central_pcs_first_word_addr & pll_first_word_addr);
	wire_mif_addr_cntr_data_mux_sel <= ( is_global_clk_div_mode & is_central_pcs);
	mif_addr_cntr_data_mux :  altgx_reconfig_cpri_mux_b6a
	  PORT MAP ( 
		data => wire_mif_addr_cntr_data_mux_data,
		result => wire_mif_addr_cntr_data_mux_result,
		sel => wire_mif_addr_cntr_data_mux_sel
	  );
	wire_pll_first_word_mux_data <= ( duplex_pma_pcs_first_pll & tx_pma_pcs_first_pll & duplex_pma_first_pll & tx_pma_first_pll);
	wire_pll_first_word_mux_sel <= ( mif_type_reg(4) & mif_type_reg(1));
	pll_first_word_mux :  altgx_reconfig_cpri_mux_c6a
	  PORT MAP ( 
		data => wire_pll_first_word_mux_data,
		result => wire_pll_first_word_mux_result,
		sel => wire_pll_first_word_mux_sel
	  );

 END RTL; --altgx_reconfig_cpri_alt2gxb_reconfig_7ba1
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altgx_reconfig_cpri IS
	PORT
	(
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_data		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		reconfig_fromgxb		: IN STD_LOGIC_VECTOR (16 DOWNTO 0);
		reconfig_mode_sel		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		write_all		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		channel_reconfig_done		: OUT STD_LOGIC ;
		reconfig_address_en		: OUT STD_LOGIC ;
		reconfig_address_out		: OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
		reconfig_togxb		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END altgx_reconfig_cpri;


ARCHITECTURE RTL OF altgx_reconfig_cpri IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt2gxb_reconfig";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "base_port_width=1;cbx_blackbox_list=-lpm_mux;enable_chl_addr_for_analog_ctrl=TRUE;intended_device_family=Stratix IV;mif_address_width=6;number_of_channels=1;number_of_reconfig_ports=1;read_base_port_width=1;enable_buf_cal=true;reconfig_fromgxb_width=17;reconfig_togxb_width=4;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (5 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC ;



	COMPONENT altgx_reconfig_cpri_alt2gxb_reconfig_7ba1
	PORT (
			reconfig_address_en	: OUT STD_LOGIC ;
			reconfig_mode_sel	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig_togxb	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			reconfig_address_out	: OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
			reconfig_fromgxb	: IN STD_LOGIC_VECTOR (16 DOWNTO 0);
			write_all	: IN STD_LOGIC ;
			channel_reconfig_done	: OUT STD_LOGIC ;
			reconfig_clk	: IN STD_LOGIC ;
			reconfig_data	: IN STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	reconfig_address_en    <= sub_wire0;
	reconfig_togxb    <= sub_wire1(3 DOWNTO 0);
	busy    <= sub_wire2;
	reconfig_address_out    <= sub_wire3(5 DOWNTO 0);
	channel_reconfig_done    <= sub_wire4;

	altgx_reconfig_cpri_alt2gxb_reconfig_7ba1_component : altgx_reconfig_cpri_alt2gxb_reconfig_7ba1
	PORT MAP (
		reconfig_mode_sel => reconfig_mode_sel,
		reconfig_fromgxb => reconfig_fromgxb,
		write_all => write_all,
		reconfig_clk => reconfig_clk,
		reconfig_data => reconfig_data,
		reconfig_address_en => sub_wire0,
		reconfig_togxb => sub_wire1,
		busy => sub_wire2,
		reconfig_address_out => sub_wire3,
		channel_reconfig_done => sub_wire4
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADCE NUMERIC "0"
-- Retrieval info: PRIVATE: CMU_PLL NUMERIC "1"
-- Retrieval info: PRIVATE: DATA_RATE NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: PRIVATE: PMA NUMERIC "1"
-- Retrieval info: PRIVATE: PROTO_SWITCH NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: BASE_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: CBX_BLACKBOX_LIST STRING "-lpm_mux"
-- Retrieval info: CONSTANT: ENABLE_CHL_ADDR_FOR_ANALOG_CTRL STRING "TRUE"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: CONSTANT: MIF_ADDRESS_WIDTH NUMERIC "6"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
-- Retrieval info: CONSTANT: NUMBER_OF_RECONFIG_PORTS NUMERIC "1"
-- Retrieval info: CONSTANT: READ_BASE_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: enable_buf_cal STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_width NUMERIC "17"
-- Retrieval info: CONSTANT: reconfig_togxb_width NUMERIC "4"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: channel_reconfig_done 0 0 0 0 OUTPUT NODEFVAL "channel_reconfig_done"
-- Retrieval info: USED_PORT: reconfig_address_en 0 0 0 0 OUTPUT NODEFVAL "reconfig_address_en"
-- Retrieval info: USED_PORT: reconfig_address_out 0 0 6 0 OUTPUT NODEFVAL "reconfig_address_out[5..0]"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_data 0 0 16 0 INPUT NODEFVAL "reconfig_data[15..0]"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 17 0 INPUT NODEFVAL "reconfig_fromgxb[16..0]"
-- Retrieval info: USED_PORT: reconfig_mode_sel 0 0 3 0 INPUT NODEFVAL "reconfig_mode_sel[2..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 OUTPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: write_all 0 0 0 0 INPUT NODEFVAL "write_all"
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_data 0 0 16 0 reconfig_data 0 0 16 0
-- Retrieval info: CONNECT: @reconfig_fromgxb 0 0 17 0 reconfig_fromgxb 0 0 17 0
-- Retrieval info: CONNECT: @reconfig_mode_sel 0 0 3 0 reconfig_mode_sel 0 0 3 0
-- Retrieval info: CONNECT: @write_all 0 0 0 0 write_all 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: channel_reconfig_done 0 0 0 0 @channel_reconfig_done 0 0 0 0
-- Retrieval info: CONNECT: reconfig_address_en 0 0 0 0 @reconfig_address_en 0 0 0 0
-- Retrieval info: CONNECT: reconfig_address_out 0 0 6 0 @reconfig_address_out 0 0 6 0
-- Retrieval info: CONNECT: reconfig_togxb 0 0 4 0 @reconfig_togxb 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_reconfig_cpri.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_reconfig_cpri.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_reconfig_cpri.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_reconfig_cpri.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_reconfig_cpri_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: LIB_FILE: lpm
