// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.



`timescale 1 ps / 1 ps

module frb_timing_lut_ram (
  CLK,
  SSR,
  ADDRA,
  EN,
  WEA,
  DIA,
  DIPA,
  DOA,
  DOPA,
  ADDRB,
  DOB,
  DOPB);

  parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  input CLK;
  input SSR;
  input [9:0] ADDRA;
  input EN;
  input WEA;
  input [31:0] DIA;
  input [3:0] DIPA;
  output [31:0] DOA;
  wire [31:0] DOA;
  output [3:0] DOPA;
  wire [3:0] DOPA;
  input [9:0] ADDRB;
  output [31:0] DOB;
  wire [31:0] DOB;
  output [3:0] DOPB;
  wire [3:0] DOPB;

  reg [35:0] RAM [1023:0];
  reg [35:0] RDATAA;
  reg [35:0] RDATAB;

//------------------------------------------------------------------------------
//MODULE BODY
//------------------------------------------------------------------------------

  initial
  begin
    RAM[   0] <= {INITP_00[  3 :   0] , INIT_00[ 31 :   0]};
    RAM[   1] <= {INITP_00[  7 :   4] , INIT_00[ 63 :  32]};
    RAM[   2] <= {INITP_00[ 11 :   8] , INIT_00[ 95 :  64]};
    RAM[   3] <= {INITP_00[ 15 :  12] , INIT_00[127 :  96]};
    RAM[   4] <= {INITP_00[ 19 :  16] , INIT_00[159 : 128]};
    RAM[   5] <= {INITP_00[ 23 :  20] , INIT_00[191 : 160]};
    RAM[   6] <= {INITP_00[ 27 :  24] , INIT_00[223 : 192]};
    RAM[   7] <= {INITP_00[ 31 :  28] , INIT_00[255 : 224]};
    RAM[   8] <= {INITP_00[ 35 :  32] , INIT_01[ 31 :   0]};
    RAM[   9] <= {INITP_00[ 39 :  36] , INIT_01[ 63 :  32]};
    RAM[  10] <= {INITP_00[ 43 :  40] , INIT_01[ 95 :  64]};
    RAM[  11] <= {INITP_00[ 47 :  44] , INIT_01[127 :  96]};
    RAM[  12] <= {INITP_00[ 51 :  48] , INIT_01[159 : 128]};
    RAM[  13] <= {INITP_00[ 55 :  52] , INIT_01[191 : 160]};
    RAM[  14] <= {INITP_00[ 59 :  56] , INIT_01[223 : 192]};
    RAM[  15] <= {INITP_00[ 63 :  60] , INIT_01[255 : 224]};
    RAM[  16] <= {INITP_00[ 67 :  64] , INIT_02[ 31 :   0]};
    RAM[  17] <= {INITP_00[ 71 :  68] , INIT_02[ 63 :  32]};
    RAM[  18] <= {INITP_00[ 75 :  72] , INIT_02[ 95 :  64]};
    RAM[  19] <= {INITP_00[ 79 :  76] , INIT_02[127 :  96]};
    RAM[  20] <= {INITP_00[ 83 :  80] , INIT_02[159 : 128]};
    RAM[  21] <= {INITP_00[ 87 :  84] , INIT_02[191 : 160]};
    RAM[  22] <= {INITP_00[ 91 :  88] , INIT_02[223 : 192]};
    RAM[  23] <= {INITP_00[ 95 :  92] , INIT_02[255 : 224]};
    RAM[  24] <= {INITP_00[ 99 :  96] , INIT_03[ 31 :   0]};
    RAM[  25] <= {INITP_00[103 : 100] , INIT_03[ 63 :  32]};
    RAM[  26] <= {INITP_00[107 : 104] , INIT_03[ 95 :  64]};
    RAM[  27] <= {INITP_00[111 : 108] , INIT_03[127 :  96]};
    RAM[  28] <= {INITP_00[115 : 112] , INIT_03[159 : 128]};
    RAM[  29] <= {INITP_00[119 : 116] , INIT_03[191 : 160]};
    RAM[  30] <= {INITP_00[123 : 120] , INIT_03[223 : 192]};
    RAM[  31] <= {INITP_00[127 : 124] , INIT_03[255 : 224]};
    RAM[  32] <= {INITP_00[131 : 128] , INIT_04[ 31 :   0]};
    RAM[  33] <= {INITP_00[135 : 132] , INIT_04[ 63 :  32]};
    RAM[  34] <= {INITP_00[139 : 136] , INIT_04[ 95 :  64]};
    RAM[  35] <= {INITP_00[143 : 140] , INIT_04[127 :  96]};
    RAM[  36] <= {INITP_00[147 : 144] , INIT_04[159 : 128]};
    RAM[  37] <= {INITP_00[151 : 148] , INIT_04[191 : 160]};
    RAM[  38] <= {INITP_00[155 : 152] , INIT_04[223 : 192]};
    RAM[  39] <= {INITP_00[159 : 156] , INIT_04[255 : 224]};
    RAM[  40] <= {INITP_00[163 : 160] , INIT_05[ 31 :   0]};
    RAM[  41] <= {INITP_00[167 : 164] , INIT_05[ 63 :  32]};
    RAM[  42] <= {INITP_00[171 : 168] , INIT_05[ 95 :  64]};
    RAM[  43] <= {INITP_00[175 : 172] , INIT_05[127 :  96]};
    RAM[  44] <= {INITP_00[179 : 176] , INIT_05[159 : 128]};
    RAM[  45] <= {INITP_00[183 : 180] , INIT_05[191 : 160]};
    RAM[  46] <= {INITP_00[187 : 184] , INIT_05[223 : 192]};
    RAM[  47] <= {INITP_00[191 : 188] , INIT_05[255 : 224]};
    RAM[  48] <= {INITP_00[195 : 192] , INIT_06[ 31 :   0]};
    RAM[  49] <= {INITP_00[199 : 196] , INIT_06[ 63 :  32]};
    RAM[  50] <= {INITP_00[203 : 200] , INIT_06[ 95 :  64]};
    RAM[  51] <= {INITP_00[207 : 204] , INIT_06[127 :  96]};
    RAM[  52] <= {INITP_00[211 : 208] , INIT_06[159 : 128]};
    RAM[  53] <= {INITP_00[215 : 212] , INIT_06[191 : 160]};
    RAM[  54] <= {INITP_00[219 : 216] , INIT_06[223 : 192]};
    RAM[  55] <= {INITP_00[223 : 220] , INIT_06[255 : 224]};
    RAM[  56] <= {INITP_00[227 : 224] , INIT_07[ 31 :   0]};
    RAM[  57] <= {INITP_00[231 : 228] , INIT_07[ 63 :  32]};
    RAM[  58] <= {INITP_00[235 : 232] , INIT_07[ 95 :  64]};
    RAM[  59] <= {INITP_00[239 : 236] , INIT_07[127 :  96]};
    RAM[  60] <= {INITP_00[243 : 240] , INIT_07[159 : 128]};
    RAM[  61] <= {INITP_00[247 : 244] , INIT_07[191 : 160]};
    RAM[  62] <= {INITP_00[251 : 248] , INIT_07[223 : 192]};
    RAM[  63] <= {INITP_00[255 : 252] , INIT_07[255 : 224]};
    RAM[  64] <= {INITP_01[  3 :   0] , INIT_08[ 31 :   0]};
    RAM[  65] <= {INITP_01[  7 :   4] , INIT_08[ 63 :  32]};
    RAM[  66] <= {INITP_01[ 11 :   8] , INIT_08[ 95 :  64]};
    RAM[  67] <= {INITP_01[ 15 :  12] , INIT_08[127 :  96]};
    RAM[  68] <= {INITP_01[ 19 :  16] , INIT_08[159 : 128]};
    RAM[  69] <= {INITP_01[ 23 :  20] , INIT_08[191 : 160]};
    RAM[  70] <= {INITP_01[ 27 :  24] , INIT_08[223 : 192]};
    RAM[  71] <= {INITP_01[ 31 :  28] , INIT_08[255 : 224]};
    RAM[  72] <= {INITP_01[ 35 :  32] , INIT_09[ 31 :   0]};
    RAM[  73] <= {INITP_01[ 39 :  36] , INIT_09[ 63 :  32]};
    RAM[  74] <= {INITP_01[ 43 :  40] , INIT_09[ 95 :  64]};
    RAM[  75] <= {INITP_01[ 47 :  44] , INIT_09[127 :  96]};
    RAM[  76] <= {INITP_01[ 51 :  48] , INIT_09[159 : 128]};
    RAM[  77] <= {INITP_01[ 55 :  52] , INIT_09[191 : 160]};
    RAM[  78] <= {INITP_01[ 59 :  56] , INIT_09[223 : 192]};
    RAM[  79] <= {INITP_01[ 63 :  60] , INIT_09[255 : 224]};
    RAM[  80] <= {INITP_01[ 67 :  64] , INIT_0A[ 31 :   0]};
    RAM[  81] <= {INITP_01[ 71 :  68] , INIT_0A[ 63 :  32]};
    RAM[  82] <= {INITP_01[ 75 :  72] , INIT_0A[ 95 :  64]};
    RAM[  83] <= {INITP_01[ 79 :  76] , INIT_0A[127 :  96]};
    RAM[  84] <= {INITP_01[ 83 :  80] , INIT_0A[159 : 128]};
    RAM[  85] <= {INITP_01[ 87 :  84] , INIT_0A[191 : 160]};
    RAM[  86] <= {INITP_01[ 91 :  88] , INIT_0A[223 : 192]};
    RAM[  87] <= {INITP_01[ 95 :  92] , INIT_0A[255 : 224]};
    RAM[  88] <= {INITP_01[ 99 :  96] , INIT_0B[ 31 :   0]};
    RAM[  89] <= {INITP_01[103 : 100] , INIT_0B[ 63 :  32]};
    RAM[  90] <= {INITP_01[107 : 104] , INIT_0B[ 95 :  64]};
    RAM[  91] <= {INITP_01[111 : 108] , INIT_0B[127 :  96]};
    RAM[  92] <= {INITP_01[115 : 112] , INIT_0B[159 : 128]};
    RAM[  93] <= {INITP_01[119 : 116] , INIT_0B[191 : 160]};
    RAM[  94] <= {INITP_01[123 : 120] , INIT_0B[223 : 192]};
    RAM[  95] <= {INITP_01[127 : 124] , INIT_0B[255 : 224]};
    RAM[  96] <= {INITP_01[131 : 128] , INIT_0C[ 31 :   0]};
    RAM[  97] <= {INITP_01[135 : 132] , INIT_0C[ 63 :  32]};
    RAM[  98] <= {INITP_01[139 : 136] , INIT_0C[ 95 :  64]};
    RAM[  99] <= {INITP_01[143 : 140] , INIT_0C[127 :  96]};
    RAM[ 100] <= {INITP_01[147 : 144] , INIT_0C[159 : 128]};
    RAM[ 101] <= {INITP_01[151 : 148] , INIT_0C[191 : 160]};
    RAM[ 102] <= {INITP_01[155 : 152] , INIT_0C[223 : 192]};
    RAM[ 103] <= {INITP_01[159 : 156] , INIT_0C[255 : 224]};
    RAM[ 104] <= {INITP_01[163 : 160] , INIT_0D[ 31 :   0]};
    RAM[ 105] <= {INITP_01[167 : 164] , INIT_0D[ 63 :  32]};
    RAM[ 106] <= {INITP_01[171 : 168] , INIT_0D[ 95 :  64]};
    RAM[ 107] <= {INITP_01[175 : 172] , INIT_0D[127 :  96]};
    RAM[ 108] <= {INITP_01[179 : 176] , INIT_0D[159 : 128]};
    RAM[ 109] <= {INITP_01[183 : 180] , INIT_0D[191 : 160]};
    RAM[ 110] <= {INITP_01[187 : 184] , INIT_0D[223 : 192]};
    RAM[ 111] <= {INITP_01[191 : 188] , INIT_0D[255 : 224]};
    RAM[ 112] <= {INITP_01[195 : 192] , INIT_0E[ 31 :   0]};
    RAM[ 113] <= {INITP_01[199 : 196] , INIT_0E[ 63 :  32]};
    RAM[ 114] <= {INITP_01[203 : 200] , INIT_0E[ 95 :  64]};
    RAM[ 115] <= {INITP_01[207 : 204] , INIT_0E[127 :  96]};
    RAM[ 116] <= {INITP_01[211 : 208] , INIT_0E[159 : 128]};
    RAM[ 117] <= {INITP_01[215 : 212] , INIT_0E[191 : 160]};
    RAM[ 118] <= {INITP_01[219 : 216] , INIT_0E[223 : 192]};
    RAM[ 119] <= {INITP_01[223 : 220] , INIT_0E[255 : 224]};
    RAM[ 120] <= {INITP_01[227 : 224] , INIT_0F[ 31 :   0]};
    RAM[ 121] <= {INITP_01[231 : 228] , INIT_0F[ 63 :  32]};
    RAM[ 122] <= {INITP_01[235 : 232] , INIT_0F[ 95 :  64]};
    RAM[ 123] <= {INITP_01[239 : 236] , INIT_0F[127 :  96]};
    RAM[ 124] <= {INITP_01[243 : 240] , INIT_0F[159 : 128]};
    RAM[ 125] <= {INITP_01[247 : 244] , INIT_0F[191 : 160]};
    RAM[ 126] <= {INITP_01[251 : 248] , INIT_0F[223 : 192]};
    RAM[ 127] <= {INITP_01[255 : 252] , INIT_0F[255 : 224]};
    RAM[ 128] <= {INITP_02[  3 :   0] , INIT_10[ 31 :   0]};
    RAM[ 129] <= {INITP_02[  7 :   4] , INIT_10[ 63 :  32]};
    RAM[ 130] <= {INITP_02[ 11 :   8] , INIT_10[ 95 :  64]};
    RAM[ 131] <= {INITP_02[ 15 :  12] , INIT_10[127 :  96]};
    RAM[ 132] <= {INITP_02[ 19 :  16] , INIT_10[159 : 128]};
    RAM[ 133] <= {INITP_02[ 23 :  20] , INIT_10[191 : 160]};
    RAM[ 134] <= {INITP_02[ 27 :  24] , INIT_10[223 : 192]};
    RAM[ 135] <= {INITP_02[ 31 :  28] , INIT_10[255 : 224]};
    RAM[ 136] <= {INITP_02[ 35 :  32] , INIT_11[ 31 :   0]};
    RAM[ 137] <= {INITP_02[ 39 :  36] , INIT_11[ 63 :  32]};
    RAM[ 138] <= {INITP_02[ 43 :  40] , INIT_11[ 95 :  64]};
    RAM[ 139] <= {INITP_02[ 47 :  44] , INIT_11[127 :  96]};
    RAM[ 140] <= {INITP_02[ 51 :  48] , INIT_11[159 : 128]};
    RAM[ 141] <= {INITP_02[ 55 :  52] , INIT_11[191 : 160]};
    RAM[ 142] <= {INITP_02[ 59 :  56] , INIT_11[223 : 192]};
    RAM[ 143] <= {INITP_02[ 63 :  60] , INIT_11[255 : 224]};
    RAM[ 144] <= {INITP_02[ 67 :  64] , INIT_12[ 31 :   0]};
    RAM[ 145] <= {INITP_02[ 71 :  68] , INIT_12[ 63 :  32]};
    RAM[ 146] <= {INITP_02[ 75 :  72] , INIT_12[ 95 :  64]};
    RAM[ 147] <= {INITP_02[ 79 :  76] , INIT_12[127 :  96]};
    RAM[ 148] <= {INITP_02[ 83 :  80] , INIT_12[159 : 128]};
    RAM[ 149] <= {INITP_02[ 87 :  84] , INIT_12[191 : 160]};
    RAM[ 150] <= {INITP_02[ 91 :  88] , INIT_12[223 : 192]};
    RAM[ 151] <= {INITP_02[ 95 :  92] , INIT_12[255 : 224]};
    RAM[ 152] <= {INITP_02[ 99 :  96] , INIT_13[ 31 :   0]};
    RAM[ 153] <= {INITP_02[103 : 100] , INIT_13[ 63 :  32]};
    RAM[ 154] <= {INITP_02[107 : 104] , INIT_13[ 95 :  64]};
    RAM[ 155] <= {INITP_02[111 : 108] , INIT_13[127 :  96]};
    RAM[ 156] <= {INITP_02[115 : 112] , INIT_13[159 : 128]};
    RAM[ 157] <= {INITP_02[119 : 116] , INIT_13[191 : 160]};
    RAM[ 158] <= {INITP_02[123 : 120] , INIT_13[223 : 192]};
    RAM[ 159] <= {INITP_02[127 : 124] , INIT_13[255 : 224]};
    RAM[ 160] <= {INITP_02[131 : 128] , INIT_14[ 31 :   0]};
    RAM[ 161] <= {INITP_02[135 : 132] , INIT_14[ 63 :  32]};
    RAM[ 162] <= {INITP_02[139 : 136] , INIT_14[ 95 :  64]};
    RAM[ 163] <= {INITP_02[143 : 140] , INIT_14[127 :  96]};
    RAM[ 164] <= {INITP_02[147 : 144] , INIT_14[159 : 128]};
    RAM[ 165] <= {INITP_02[151 : 148] , INIT_14[191 : 160]};
    RAM[ 166] <= {INITP_02[155 : 152] , INIT_14[223 : 192]};
    RAM[ 167] <= {INITP_02[159 : 156] , INIT_14[255 : 224]};
    RAM[ 168] <= {INITP_02[163 : 160] , INIT_15[ 31 :   0]};
    RAM[ 169] <= {INITP_02[167 : 164] , INIT_15[ 63 :  32]};
    RAM[ 170] <= {INITP_02[171 : 168] , INIT_15[ 95 :  64]};
    RAM[ 171] <= {INITP_02[175 : 172] , INIT_15[127 :  96]};
    RAM[ 172] <= {INITP_02[179 : 176] , INIT_15[159 : 128]};
    RAM[ 173] <= {INITP_02[183 : 180] , INIT_15[191 : 160]};
    RAM[ 174] <= {INITP_02[187 : 184] , INIT_15[223 : 192]};
    RAM[ 175] <= {INITP_02[191 : 188] , INIT_15[255 : 224]};
    RAM[ 176] <= {INITP_02[195 : 192] , INIT_16[ 31 :   0]};
    RAM[ 177] <= {INITP_02[199 : 196] , INIT_16[ 63 :  32]};
    RAM[ 178] <= {INITP_02[203 : 200] , INIT_16[ 95 :  64]};
    RAM[ 179] <= {INITP_02[207 : 204] , INIT_16[127 :  96]};
    RAM[ 180] <= {INITP_02[211 : 208] , INIT_16[159 : 128]};
    RAM[ 181] <= {INITP_02[215 : 212] , INIT_16[191 : 160]};
    RAM[ 182] <= {INITP_02[219 : 216] , INIT_16[223 : 192]};
    RAM[ 183] <= {INITP_02[223 : 220] , INIT_16[255 : 224]};
    RAM[ 184] <= {INITP_02[227 : 224] , INIT_17[ 31 :   0]};
    RAM[ 185] <= {INITP_02[231 : 228] , INIT_17[ 63 :  32]};
    RAM[ 186] <= {INITP_02[235 : 232] , INIT_17[ 95 :  64]};
    RAM[ 187] <= {INITP_02[239 : 236] , INIT_17[127 :  96]};
    RAM[ 188] <= {INITP_02[243 : 240] , INIT_17[159 : 128]};
    RAM[ 189] <= {INITP_02[247 : 244] , INIT_17[191 : 160]};
    RAM[ 190] <= {INITP_02[251 : 248] , INIT_17[223 : 192]};
    RAM[ 191] <= {INITP_02[255 : 252] , INIT_17[255 : 224]};
    RAM[ 192] <= {INITP_03[  3 :   0] , INIT_18[ 31 :   0]};
    RAM[ 193] <= {INITP_03[  7 :   4] , INIT_18[ 63 :  32]};
    RAM[ 194] <= {INITP_03[ 11 :   8] , INIT_18[ 95 :  64]};
    RAM[ 195] <= {INITP_03[ 15 :  12] , INIT_18[127 :  96]};
    RAM[ 196] <= {INITP_03[ 19 :  16] , INIT_18[159 : 128]};
    RAM[ 197] <= {INITP_03[ 23 :  20] , INIT_18[191 : 160]};
    RAM[ 198] <= {INITP_03[ 27 :  24] , INIT_18[223 : 192]};
    RAM[ 199] <= {INITP_03[ 31 :  28] , INIT_18[255 : 224]};
    RAM[ 200] <= {INITP_03[ 35 :  32] , INIT_19[ 31 :   0]};
    RAM[ 201] <= {INITP_03[ 39 :  36] , INIT_19[ 63 :  32]};
    RAM[ 202] <= {INITP_03[ 43 :  40] , INIT_19[ 95 :  64]};
    RAM[ 203] <= {INITP_03[ 47 :  44] , INIT_19[127 :  96]};
    RAM[ 204] <= {INITP_03[ 51 :  48] , INIT_19[159 : 128]};
    RAM[ 205] <= {INITP_03[ 55 :  52] , INIT_19[191 : 160]};
    RAM[ 206] <= {INITP_03[ 59 :  56] , INIT_19[223 : 192]};
    RAM[ 207] <= {INITP_03[ 63 :  60] , INIT_19[255 : 224]};
    RAM[ 208] <= {INITP_03[ 67 :  64] , INIT_1A[ 31 :   0]};
    RAM[ 209] <= {INITP_03[ 71 :  68] , INIT_1A[ 63 :  32]};
    RAM[ 210] <= {INITP_03[ 75 :  72] , INIT_1A[ 95 :  64]};
    RAM[ 211] <= {INITP_03[ 79 :  76] , INIT_1A[127 :  96]};
    RAM[ 212] <= {INITP_03[ 83 :  80] , INIT_1A[159 : 128]};
    RAM[ 213] <= {INITP_03[ 87 :  84] , INIT_1A[191 : 160]};
    RAM[ 214] <= {INITP_03[ 91 :  88] , INIT_1A[223 : 192]};
    RAM[ 215] <= {INITP_03[ 95 :  92] , INIT_1A[255 : 224]};
    RAM[ 216] <= {INITP_03[ 99 :  96] , INIT_1B[ 31 :   0]};
    RAM[ 217] <= {INITP_03[103 : 100] , INIT_1B[ 63 :  32]};
    RAM[ 218] <= {INITP_03[107 : 104] , INIT_1B[ 95 :  64]};
    RAM[ 219] <= {INITP_03[111 : 108] , INIT_1B[127 :  96]};
    RAM[ 220] <= {INITP_03[115 : 112] , INIT_1B[159 : 128]};
    RAM[ 221] <= {INITP_03[119 : 116] , INIT_1B[191 : 160]};
    RAM[ 222] <= {INITP_03[123 : 120] , INIT_1B[223 : 192]};
    RAM[ 223] <= {INITP_03[127 : 124] , INIT_1B[255 : 224]};
    RAM[ 224] <= {INITP_03[131 : 128] , INIT_1C[ 31 :   0]};
    RAM[ 225] <= {INITP_03[135 : 132] , INIT_1C[ 63 :  32]};
    RAM[ 226] <= {INITP_03[139 : 136] , INIT_1C[ 95 :  64]};
    RAM[ 227] <= {INITP_03[143 : 140] , INIT_1C[127 :  96]};
    RAM[ 228] <= {INITP_03[147 : 144] , INIT_1C[159 : 128]};
    RAM[ 229] <= {INITP_03[151 : 148] , INIT_1C[191 : 160]};
    RAM[ 230] <= {INITP_03[155 : 152] , INIT_1C[223 : 192]};
    RAM[ 231] <= {INITP_03[159 : 156] , INIT_1C[255 : 224]};
    RAM[ 232] <= {INITP_03[163 : 160] , INIT_1D[ 31 :   0]};
    RAM[ 233] <= {INITP_03[167 : 164] , INIT_1D[ 63 :  32]};
    RAM[ 234] <= {INITP_03[171 : 168] , INIT_1D[ 95 :  64]};
    RAM[ 235] <= {INITP_03[175 : 172] , INIT_1D[127 :  96]};
    RAM[ 236] <= {INITP_03[179 : 176] , INIT_1D[159 : 128]};
    RAM[ 237] <= {INITP_03[183 : 180] , INIT_1D[191 : 160]};
    RAM[ 238] <= {INITP_03[187 : 184] , INIT_1D[223 : 192]};
    RAM[ 239] <= {INITP_03[191 : 188] , INIT_1D[255 : 224]};
    RAM[ 240] <= {INITP_03[195 : 192] , INIT_1E[ 31 :   0]};
    RAM[ 241] <= {INITP_03[199 : 196] , INIT_1E[ 63 :  32]};
    RAM[ 242] <= {INITP_03[203 : 200] , INIT_1E[ 95 :  64]};
    RAM[ 243] <= {INITP_03[207 : 204] , INIT_1E[127 :  96]};
    RAM[ 244] <= {INITP_03[211 : 208] , INIT_1E[159 : 128]};
    RAM[ 245] <= {INITP_03[215 : 212] , INIT_1E[191 : 160]};
    RAM[ 246] <= {INITP_03[219 : 216] , INIT_1E[223 : 192]};
    RAM[ 247] <= {INITP_03[223 : 220] , INIT_1E[255 : 224]};
    RAM[ 248] <= {INITP_03[227 : 224] , INIT_1F[ 31 :   0]};
    RAM[ 249] <= {INITP_03[231 : 228] , INIT_1F[ 63 :  32]};
    RAM[ 250] <= {INITP_03[235 : 232] , INIT_1F[ 95 :  64]};
    RAM[ 251] <= {INITP_03[239 : 236] , INIT_1F[127 :  96]};
    RAM[ 252] <= {INITP_03[243 : 240] , INIT_1F[159 : 128]};
    RAM[ 253] <= {INITP_03[247 : 244] , INIT_1F[191 : 160]};
    RAM[ 254] <= {INITP_03[251 : 248] , INIT_1F[223 : 192]};
    RAM[ 255] <= {INITP_03[255 : 252] , INIT_1F[255 : 224]};
    RAM[ 256] <= {INITP_04[  3 :   0] , INIT_20[ 31 :   0]};
    RAM[ 257] <= {INITP_04[  7 :   4] , INIT_20[ 63 :  32]};
    RAM[ 258] <= {INITP_04[ 11 :   8] , INIT_20[ 95 :  64]};
    RAM[ 259] <= {INITP_04[ 15 :  12] , INIT_20[127 :  96]};
    RAM[ 260] <= {INITP_04[ 19 :  16] , INIT_20[159 : 128]};
    RAM[ 261] <= {INITP_04[ 23 :  20] , INIT_20[191 : 160]};
    RAM[ 262] <= {INITP_04[ 27 :  24] , INIT_20[223 : 192]};
    RAM[ 263] <= {INITP_04[ 31 :  28] , INIT_20[255 : 224]};
    RAM[ 264] <= {INITP_04[ 35 :  32] , INIT_21[ 31 :   0]};
    RAM[ 265] <= {INITP_04[ 39 :  36] , INIT_21[ 63 :  32]};
    RAM[ 266] <= {INITP_04[ 43 :  40] , INIT_21[ 95 :  64]};
    RAM[ 267] <= {INITP_04[ 47 :  44] , INIT_21[127 :  96]};
    RAM[ 268] <= {INITP_04[ 51 :  48] , INIT_21[159 : 128]};
    RAM[ 269] <= {INITP_04[ 55 :  52] , INIT_21[191 : 160]};
    RAM[ 270] <= {INITP_04[ 59 :  56] , INIT_21[223 : 192]};
    RAM[ 271] <= {INITP_04[ 63 :  60] , INIT_21[255 : 224]};
    RAM[ 272] <= {INITP_04[ 67 :  64] , INIT_22[ 31 :   0]};
    RAM[ 273] <= {INITP_04[ 71 :  68] , INIT_22[ 63 :  32]};
    RAM[ 274] <= {INITP_04[ 75 :  72] , INIT_22[ 95 :  64]};
    RAM[ 275] <= {INITP_04[ 79 :  76] , INIT_22[127 :  96]};
    RAM[ 276] <= {INITP_04[ 83 :  80] , INIT_22[159 : 128]};
    RAM[ 277] <= {INITP_04[ 87 :  84] , INIT_22[191 : 160]};
    RAM[ 278] <= {INITP_04[ 91 :  88] , INIT_22[223 : 192]};
    RAM[ 279] <= {INITP_04[ 95 :  92] , INIT_22[255 : 224]};
    RAM[ 280] <= {INITP_04[ 99 :  96] , INIT_23[ 31 :   0]};
    RAM[ 281] <= {INITP_04[103 : 100] , INIT_23[ 63 :  32]};
    RAM[ 282] <= {INITP_04[107 : 104] , INIT_23[ 95 :  64]};
    RAM[ 283] <= {INITP_04[111 : 108] , INIT_23[127 :  96]};
    RAM[ 284] <= {INITP_04[115 : 112] , INIT_23[159 : 128]};
    RAM[ 285] <= {INITP_04[119 : 116] , INIT_23[191 : 160]};
    RAM[ 286] <= {INITP_04[123 : 120] , INIT_23[223 : 192]};
    RAM[ 287] <= {INITP_04[127 : 124] , INIT_23[255 : 224]};
    RAM[ 288] <= {INITP_04[131 : 128] , INIT_24[ 31 :   0]};
    RAM[ 289] <= {INITP_04[135 : 132] , INIT_24[ 63 :  32]};
    RAM[ 290] <= {INITP_04[139 : 136] , INIT_24[ 95 :  64]};
    RAM[ 291] <= {INITP_04[143 : 140] , INIT_24[127 :  96]};
    RAM[ 292] <= {INITP_04[147 : 144] , INIT_24[159 : 128]};
    RAM[ 293] <= {INITP_04[151 : 148] , INIT_24[191 : 160]};
    RAM[ 294] <= {INITP_04[155 : 152] , INIT_24[223 : 192]};
    RAM[ 295] <= {INITP_04[159 : 156] , INIT_24[255 : 224]};
    RAM[ 296] <= {INITP_04[163 : 160] , INIT_25[ 31 :   0]};
    RAM[ 297] <= {INITP_04[167 : 164] , INIT_25[ 63 :  32]};
    RAM[ 298] <= {INITP_04[171 : 168] , INIT_25[ 95 :  64]};
    RAM[ 299] <= {INITP_04[175 : 172] , INIT_25[127 :  96]};
    RAM[ 300] <= {INITP_04[179 : 176] , INIT_25[159 : 128]};
    RAM[ 301] <= {INITP_04[183 : 180] , INIT_25[191 : 160]};
    RAM[ 302] <= {INITP_04[187 : 184] , INIT_25[223 : 192]};
    RAM[ 303] <= {INITP_04[191 : 188] , INIT_25[255 : 224]};
    RAM[ 304] <= {INITP_04[195 : 192] , INIT_26[ 31 :   0]};
    RAM[ 305] <= {INITP_04[199 : 196] , INIT_26[ 63 :  32]};
    RAM[ 306] <= {INITP_04[203 : 200] , INIT_26[ 95 :  64]};
    RAM[ 307] <= {INITP_04[207 : 204] , INIT_26[127 :  96]};
    RAM[ 308] <= {INITP_04[211 : 208] , INIT_26[159 : 128]};
    RAM[ 309] <= {INITP_04[215 : 212] , INIT_26[191 : 160]};
    RAM[ 310] <= {INITP_04[219 : 216] , INIT_26[223 : 192]};
    RAM[ 311] <= {INITP_04[223 : 220] , INIT_26[255 : 224]};
    RAM[ 312] <= {INITP_04[227 : 224] , INIT_27[ 31 :   0]};
    RAM[ 313] <= {INITP_04[231 : 228] , INIT_27[ 63 :  32]};
    RAM[ 314] <= {INITP_04[235 : 232] , INIT_27[ 95 :  64]};
    RAM[ 315] <= {INITP_04[239 : 236] , INIT_27[127 :  96]};
    RAM[ 316] <= {INITP_04[243 : 240] , INIT_27[159 : 128]};
    RAM[ 317] <= {INITP_04[247 : 244] , INIT_27[191 : 160]};
    RAM[ 318] <= {INITP_04[251 : 248] , INIT_27[223 : 192]};
    RAM[ 319] <= {INITP_04[255 : 252] , INIT_27[255 : 224]};
    RAM[ 320] <= {INITP_05[  3 :   0] , INIT_28[ 31 :   0]};
    RAM[ 321] <= {INITP_05[  7 :   4] , INIT_28[ 63 :  32]};
    RAM[ 322] <= {INITP_05[ 11 :   8] , INIT_28[ 95 :  64]};
    RAM[ 323] <= {INITP_05[ 15 :  12] , INIT_28[127 :  96]};
    RAM[ 324] <= {INITP_05[ 19 :  16] , INIT_28[159 : 128]};
    RAM[ 325] <= {INITP_05[ 23 :  20] , INIT_28[191 : 160]};
    RAM[ 326] <= {INITP_05[ 27 :  24] , INIT_28[223 : 192]};
    RAM[ 327] <= {INITP_05[ 31 :  28] , INIT_28[255 : 224]};
    RAM[ 328] <= {INITP_05[ 35 :  32] , INIT_29[ 31 :   0]};
    RAM[ 329] <= {INITP_05[ 39 :  36] , INIT_29[ 63 :  32]};
    RAM[ 330] <= {INITP_05[ 43 :  40] , INIT_29[ 95 :  64]};
    RAM[ 331] <= {INITP_05[ 47 :  44] , INIT_29[127 :  96]};
    RAM[ 332] <= {INITP_05[ 51 :  48] , INIT_29[159 : 128]};
    RAM[ 333] <= {INITP_05[ 55 :  52] , INIT_29[191 : 160]};
    RAM[ 334] <= {INITP_05[ 59 :  56] , INIT_29[223 : 192]};
    RAM[ 335] <= {INITP_05[ 63 :  60] , INIT_29[255 : 224]};
    RAM[ 336] <= {INITP_05[ 67 :  64] , INIT_2A[ 31 :   0]};
    RAM[ 337] <= {INITP_05[ 71 :  68] , INIT_2A[ 63 :  32]};
    RAM[ 338] <= {INITP_05[ 75 :  72] , INIT_2A[ 95 :  64]};
    RAM[ 339] <= {INITP_05[ 79 :  76] , INIT_2A[127 :  96]};
    RAM[ 340] <= {INITP_05[ 83 :  80] , INIT_2A[159 : 128]};
    RAM[ 341] <= {INITP_05[ 87 :  84] , INIT_2A[191 : 160]};
    RAM[ 342] <= {INITP_05[ 91 :  88] , INIT_2A[223 : 192]};
    RAM[ 343] <= {INITP_05[ 95 :  92] , INIT_2A[255 : 224]};
    RAM[ 344] <= {INITP_05[ 99 :  96] , INIT_2B[ 31 :   0]};
    RAM[ 345] <= {INITP_05[103 : 100] , INIT_2B[ 63 :  32]};
    RAM[ 346] <= {INITP_05[107 : 104] , INIT_2B[ 95 :  64]};
    RAM[ 347] <= {INITP_05[111 : 108] , INIT_2B[127 :  96]};
    RAM[ 348] <= {INITP_05[115 : 112] , INIT_2B[159 : 128]};
    RAM[ 349] <= {INITP_05[119 : 116] , INIT_2B[191 : 160]};
    RAM[ 350] <= {INITP_05[123 : 120] , INIT_2B[223 : 192]};
    RAM[ 351] <= {INITP_05[127 : 124] , INIT_2B[255 : 224]};
    RAM[ 352] <= {INITP_05[131 : 128] , INIT_2C[ 31 :   0]};
    RAM[ 353] <= {INITP_05[135 : 132] , INIT_2C[ 63 :  32]};
    RAM[ 354] <= {INITP_05[139 : 136] , INIT_2C[ 95 :  64]};
    RAM[ 355] <= {INITP_05[143 : 140] , INIT_2C[127 :  96]};
    RAM[ 356] <= {INITP_05[147 : 144] , INIT_2C[159 : 128]};
    RAM[ 357] <= {INITP_05[151 : 148] , INIT_2C[191 : 160]};
    RAM[ 358] <= {INITP_05[155 : 152] , INIT_2C[223 : 192]};
    RAM[ 359] <= {INITP_05[159 : 156] , INIT_2C[255 : 224]};
    RAM[ 360] <= {INITP_05[163 : 160] , INIT_2D[ 31 :   0]};
    RAM[ 361] <= {INITP_05[167 : 164] , INIT_2D[ 63 :  32]};
    RAM[ 362] <= {INITP_05[171 : 168] , INIT_2D[ 95 :  64]};
    RAM[ 363] <= {INITP_05[175 : 172] , INIT_2D[127 :  96]};
    RAM[ 364] <= {INITP_05[179 : 176] , INIT_2D[159 : 128]};
    RAM[ 365] <= {INITP_05[183 : 180] , INIT_2D[191 : 160]};
    RAM[ 366] <= {INITP_05[187 : 184] , INIT_2D[223 : 192]};
    RAM[ 367] <= {INITP_05[191 : 188] , INIT_2D[255 : 224]};
    RAM[ 368] <= {INITP_05[195 : 192] , INIT_2E[ 31 :   0]};
    RAM[ 369] <= {INITP_05[199 : 196] , INIT_2E[ 63 :  32]};
    RAM[ 370] <= {INITP_05[203 : 200] , INIT_2E[ 95 :  64]};
    RAM[ 371] <= {INITP_05[207 : 204] , INIT_2E[127 :  96]};
    RAM[ 372] <= {INITP_05[211 : 208] , INIT_2E[159 : 128]};
    RAM[ 373] <= {INITP_05[215 : 212] , INIT_2E[191 : 160]};
    RAM[ 374] <= {INITP_05[219 : 216] , INIT_2E[223 : 192]};
    RAM[ 375] <= {INITP_05[223 : 220] , INIT_2E[255 : 224]};
    RAM[ 376] <= {INITP_05[227 : 224] , INIT_2F[ 31 :   0]};
    RAM[ 377] <= {INITP_05[231 : 228] , INIT_2F[ 63 :  32]};
    RAM[ 378] <= {INITP_05[235 : 232] , INIT_2F[ 95 :  64]};
    RAM[ 379] <= {INITP_05[239 : 236] , INIT_2F[127 :  96]};
    RAM[ 380] <= {INITP_05[243 : 240] , INIT_2F[159 : 128]};
    RAM[ 381] <= {INITP_05[247 : 244] , INIT_2F[191 : 160]};
    RAM[ 382] <= {INITP_05[251 : 248] , INIT_2F[223 : 192]};
    RAM[ 383] <= {INITP_05[255 : 252] , INIT_2F[255 : 224]};
    RAM[ 384] <= {INITP_06[  3 :   0] , INIT_30[ 31 :   0]};
    RAM[ 385] <= {INITP_06[  7 :   4] , INIT_30[ 63 :  32]};
    RAM[ 386] <= {INITP_06[ 11 :   8] , INIT_30[ 95 :  64]};
    RAM[ 387] <= {INITP_06[ 15 :  12] , INIT_30[127 :  96]};
    RAM[ 388] <= {INITP_06[ 19 :  16] , INIT_30[159 : 128]};
    RAM[ 389] <= {INITP_06[ 23 :  20] , INIT_30[191 : 160]};
    RAM[ 390] <= {INITP_06[ 27 :  24] , INIT_30[223 : 192]};
    RAM[ 391] <= {INITP_06[ 31 :  28] , INIT_30[255 : 224]};
    RAM[ 392] <= {INITP_06[ 35 :  32] , INIT_31[ 31 :   0]};
    RAM[ 393] <= {INITP_06[ 39 :  36] , INIT_31[ 63 :  32]};
    RAM[ 394] <= {INITP_06[ 43 :  40] , INIT_31[ 95 :  64]};
    RAM[ 395] <= {INITP_06[ 47 :  44] , INIT_31[127 :  96]};
    RAM[ 396] <= {INITP_06[ 51 :  48] , INIT_31[159 : 128]};
    RAM[ 397] <= {INITP_06[ 55 :  52] , INIT_31[191 : 160]};
    RAM[ 398] <= {INITP_06[ 59 :  56] , INIT_31[223 : 192]};
    RAM[ 399] <= {INITP_06[ 63 :  60] , INIT_31[255 : 224]};
    RAM[ 400] <= {INITP_06[ 67 :  64] , INIT_32[ 31 :   0]};
    RAM[ 401] <= {INITP_06[ 71 :  68] , INIT_32[ 63 :  32]};
    RAM[ 402] <= {INITP_06[ 75 :  72] , INIT_32[ 95 :  64]};
    RAM[ 403] <= {INITP_06[ 79 :  76] , INIT_32[127 :  96]};
    RAM[ 404] <= {INITP_06[ 83 :  80] , INIT_32[159 : 128]};
    RAM[ 405] <= {INITP_06[ 87 :  84] , INIT_32[191 : 160]};
    RAM[ 406] <= {INITP_06[ 91 :  88] , INIT_32[223 : 192]};
    RAM[ 407] <= {INITP_06[ 95 :  92] , INIT_32[255 : 224]};
    RAM[ 408] <= {INITP_06[ 99 :  96] , INIT_33[ 31 :   0]};
    RAM[ 409] <= {INITP_06[103 : 100] , INIT_33[ 63 :  32]};
    RAM[ 410] <= {INITP_06[107 : 104] , INIT_33[ 95 :  64]};
    RAM[ 411] <= {INITP_06[111 : 108] , INIT_33[127 :  96]};
    RAM[ 412] <= {INITP_06[115 : 112] , INIT_33[159 : 128]};
    RAM[ 413] <= {INITP_06[119 : 116] , INIT_33[191 : 160]};
    RAM[ 414] <= {INITP_06[123 : 120] , INIT_33[223 : 192]};
    RAM[ 415] <= {INITP_06[127 : 124] , INIT_33[255 : 224]};
    RAM[ 416] <= {INITP_06[131 : 128] , INIT_34[ 31 :   0]};
    RAM[ 417] <= {INITP_06[135 : 132] , INIT_34[ 63 :  32]};
    RAM[ 418] <= {INITP_06[139 : 136] , INIT_34[ 95 :  64]};
    RAM[ 419] <= {INITP_06[143 : 140] , INIT_34[127 :  96]};
    RAM[ 420] <= {INITP_06[147 : 144] , INIT_34[159 : 128]};
    RAM[ 421] <= {INITP_06[151 : 148] , INIT_34[191 : 160]};
    RAM[ 422] <= {INITP_06[155 : 152] , INIT_34[223 : 192]};
    RAM[ 423] <= {INITP_06[159 : 156] , INIT_34[255 : 224]};
    RAM[ 424] <= {INITP_06[163 : 160] , INIT_35[ 31 :   0]};
    RAM[ 425] <= {INITP_06[167 : 164] , INIT_35[ 63 :  32]};
    RAM[ 426] <= {INITP_06[171 : 168] , INIT_35[ 95 :  64]};
    RAM[ 427] <= {INITP_06[175 : 172] , INIT_35[127 :  96]};
    RAM[ 428] <= {INITP_06[179 : 176] , INIT_35[159 : 128]};
    RAM[ 429] <= {INITP_06[183 : 180] , INIT_35[191 : 160]};
    RAM[ 430] <= {INITP_06[187 : 184] , INIT_35[223 : 192]};
    RAM[ 431] <= {INITP_06[191 : 188] , INIT_35[255 : 224]};
    RAM[ 432] <= {INITP_06[195 : 192] , INIT_36[ 31 :   0]};
    RAM[ 433] <= {INITP_06[199 : 196] , INIT_36[ 63 :  32]};
    RAM[ 434] <= {INITP_06[203 : 200] , INIT_36[ 95 :  64]};
    RAM[ 435] <= {INITP_06[207 : 204] , INIT_36[127 :  96]};
    RAM[ 436] <= {INITP_06[211 : 208] , INIT_36[159 : 128]};
    RAM[ 437] <= {INITP_06[215 : 212] , INIT_36[191 : 160]};
    RAM[ 438] <= {INITP_06[219 : 216] , INIT_36[223 : 192]};
    RAM[ 439] <= {INITP_06[223 : 220] , INIT_36[255 : 224]};
    RAM[ 440] <= {INITP_06[227 : 224] , INIT_37[ 31 :   0]};
    RAM[ 441] <= {INITP_06[231 : 228] , INIT_37[ 63 :  32]};
    RAM[ 442] <= {INITP_06[235 : 232] , INIT_37[ 95 :  64]};
    RAM[ 443] <= {INITP_06[239 : 236] , INIT_37[127 :  96]};
    RAM[ 444] <= {INITP_06[243 : 240] , INIT_37[159 : 128]};
    RAM[ 445] <= {INITP_06[247 : 244] , INIT_37[191 : 160]};
    RAM[ 446] <= {INITP_06[251 : 248] , INIT_37[223 : 192]};
    RAM[ 447] <= {INITP_06[255 : 252] , INIT_37[255 : 224]};
    RAM[ 448] <= {INITP_07[  3 :   0] , INIT_38[ 31 :   0]};
    RAM[ 449] <= {INITP_07[  7 :   4] , INIT_38[ 63 :  32]};
    RAM[ 450] <= {INITP_07[ 11 :   8] , INIT_38[ 95 :  64]};
    RAM[ 451] <= {INITP_07[ 15 :  12] , INIT_38[127 :  96]};
    RAM[ 452] <= {INITP_07[ 19 :  16] , INIT_38[159 : 128]};
    RAM[ 453] <= {INITP_07[ 23 :  20] , INIT_38[191 : 160]};
    RAM[ 454] <= {INITP_07[ 27 :  24] , INIT_38[223 : 192]};
    RAM[ 455] <= {INITP_07[ 31 :  28] , INIT_38[255 : 224]};
    RAM[ 456] <= {INITP_07[ 35 :  32] , INIT_39[ 31 :   0]};
    RAM[ 457] <= {INITP_07[ 39 :  36] , INIT_39[ 63 :  32]};
    RAM[ 458] <= {INITP_07[ 43 :  40] , INIT_39[ 95 :  64]};
    RAM[ 459] <= {INITP_07[ 47 :  44] , INIT_39[127 :  96]};
    RAM[ 460] <= {INITP_07[ 51 :  48] , INIT_39[159 : 128]};
    RAM[ 461] <= {INITP_07[ 55 :  52] , INIT_39[191 : 160]};
    RAM[ 462] <= {INITP_07[ 59 :  56] , INIT_39[223 : 192]};
    RAM[ 463] <= {INITP_07[ 63 :  60] , INIT_39[255 : 224]};
    RAM[ 464] <= {INITP_07[ 67 :  64] , INIT_3A[ 31 :   0]};
    RAM[ 465] <= {INITP_07[ 71 :  68] , INIT_3A[ 63 :  32]};
    RAM[ 466] <= {INITP_07[ 75 :  72] , INIT_3A[ 95 :  64]};
    RAM[ 467] <= {INITP_07[ 79 :  76] , INIT_3A[127 :  96]};
    RAM[ 468] <= {INITP_07[ 83 :  80] , INIT_3A[159 : 128]};
    RAM[ 469] <= {INITP_07[ 87 :  84] , INIT_3A[191 : 160]};
    RAM[ 470] <= {INITP_07[ 91 :  88] , INIT_3A[223 : 192]};
    RAM[ 471] <= {INITP_07[ 95 :  92] , INIT_3A[255 : 224]};
    RAM[ 472] <= {INITP_07[ 99 :  96] , INIT_3B[ 31 :   0]};
    RAM[ 473] <= {INITP_07[103 : 100] , INIT_3B[ 63 :  32]};
    RAM[ 474] <= {INITP_07[107 : 104] , INIT_3B[ 95 :  64]};
    RAM[ 475] <= {INITP_07[111 : 108] , INIT_3B[127 :  96]};
    RAM[ 476] <= {INITP_07[115 : 112] , INIT_3B[159 : 128]};
    RAM[ 477] <= {INITP_07[119 : 116] , INIT_3B[191 : 160]};
    RAM[ 478] <= {INITP_07[123 : 120] , INIT_3B[223 : 192]};
    RAM[ 479] <= {INITP_07[127 : 124] , INIT_3B[255 : 224]};
    RAM[ 480] <= {INITP_07[131 : 128] , INIT_3C[ 31 :   0]};
    RAM[ 481] <= {INITP_07[135 : 132] , INIT_3C[ 63 :  32]};
    RAM[ 482] <= {INITP_07[139 : 136] , INIT_3C[ 95 :  64]};
    RAM[ 483] <= {INITP_07[143 : 140] , INIT_3C[127 :  96]};
    RAM[ 484] <= {INITP_07[147 : 144] , INIT_3C[159 : 128]};
    RAM[ 485] <= {INITP_07[151 : 148] , INIT_3C[191 : 160]};
    RAM[ 486] <= {INITP_07[155 : 152] , INIT_3C[223 : 192]};
    RAM[ 487] <= {INITP_07[159 : 156] , INIT_3C[255 : 224]};
    RAM[ 488] <= {INITP_07[163 : 160] , INIT_3D[ 31 :   0]};
    RAM[ 489] <= {INITP_07[167 : 164] , INIT_3D[ 63 :  32]};
    RAM[ 490] <= {INITP_07[171 : 168] , INIT_3D[ 95 :  64]};
    RAM[ 491] <= {INITP_07[175 : 172] , INIT_3D[127 :  96]};
    RAM[ 492] <= {INITP_07[179 : 176] , INIT_3D[159 : 128]};
    RAM[ 493] <= {INITP_07[183 : 180] , INIT_3D[191 : 160]};
    RAM[ 494] <= {INITP_07[187 : 184] , INIT_3D[223 : 192]};
    RAM[ 495] <= {INITP_07[191 : 188] , INIT_3D[255 : 224]};
    RAM[ 496] <= {INITP_07[195 : 192] , INIT_3E[ 31 :   0]};
    RAM[ 497] <= {INITP_07[199 : 196] , INIT_3E[ 63 :  32]};
    RAM[ 498] <= {INITP_07[203 : 200] , INIT_3E[ 95 :  64]};
    RAM[ 499] <= {INITP_07[207 : 204] , INIT_3E[127 :  96]};
    RAM[ 500] <= {INITP_07[211 : 208] , INIT_3E[159 : 128]};
    RAM[ 501] <= {INITP_07[215 : 212] , INIT_3E[191 : 160]};
    RAM[ 502] <= {INITP_07[219 : 216] , INIT_3E[223 : 192]};
    RAM[ 503] <= {INITP_07[223 : 220] , INIT_3E[255 : 224]};
    RAM[ 504] <= {INITP_07[227 : 224] , INIT_3F[ 31 :   0]};
    RAM[ 505] <= {INITP_07[231 : 228] , INIT_3F[ 63 :  32]};
    RAM[ 506] <= {INITP_07[235 : 232] , INIT_3F[ 95 :  64]};
    RAM[ 507] <= {INITP_07[239 : 236] , INIT_3F[127 :  96]};
    RAM[ 508] <= {INITP_07[243 : 240] , INIT_3F[159 : 128]};
    RAM[ 509] <= {INITP_07[247 : 244] , INIT_3F[191 : 160]};
    RAM[ 510] <= {INITP_07[251 : 248] , INIT_3F[223 : 192]};
    RAM[ 511] <= {INITP_07[255 : 252] , INIT_3F[255 : 224]};
    RAM[ 512] <= {INITP_08[  3 :   0] , INIT_40[ 31 :   0]};
    RAM[ 513] <= {INITP_08[  7 :   4] , INIT_40[ 63 :  32]};
    RAM[ 514] <= {INITP_08[ 11 :   8] , INIT_40[ 95 :  64]};
    RAM[ 515] <= {INITP_08[ 15 :  12] , INIT_40[127 :  96]};
    RAM[ 516] <= {INITP_08[ 19 :  16] , INIT_40[159 : 128]};
    RAM[ 517] <= {INITP_08[ 23 :  20] , INIT_40[191 : 160]};
    RAM[ 518] <= {INITP_08[ 27 :  24] , INIT_40[223 : 192]};
    RAM[ 519] <= {INITP_08[ 31 :  28] , INIT_40[255 : 224]};
    RAM[ 520] <= {INITP_08[ 35 :  32] , INIT_41[ 31 :   0]};
    RAM[ 521] <= {INITP_08[ 39 :  36] , INIT_41[ 63 :  32]};
    RAM[ 522] <= {INITP_08[ 43 :  40] , INIT_41[ 95 :  64]};
    RAM[ 523] <= {INITP_08[ 47 :  44] , INIT_41[127 :  96]};
    RAM[ 524] <= {INITP_08[ 51 :  48] , INIT_41[159 : 128]};
    RAM[ 525] <= {INITP_08[ 55 :  52] , INIT_41[191 : 160]};
    RAM[ 526] <= {INITP_08[ 59 :  56] , INIT_41[223 : 192]};
    RAM[ 527] <= {INITP_08[ 63 :  60] , INIT_41[255 : 224]};
    RAM[ 528] <= {INITP_08[ 67 :  64] , INIT_42[ 31 :   0]};
    RAM[ 529] <= {INITP_08[ 71 :  68] , INIT_42[ 63 :  32]};
    RAM[ 530] <= {INITP_08[ 75 :  72] , INIT_42[ 95 :  64]};
    RAM[ 531] <= {INITP_08[ 79 :  76] , INIT_42[127 :  96]};
    RAM[ 532] <= {INITP_08[ 83 :  80] , INIT_42[159 : 128]};
    RAM[ 533] <= {INITP_08[ 87 :  84] , INIT_42[191 : 160]};
    RAM[ 534] <= {INITP_08[ 91 :  88] , INIT_42[223 : 192]};
    RAM[ 535] <= {INITP_08[ 95 :  92] , INIT_42[255 : 224]};
    RAM[ 536] <= {INITP_08[ 99 :  96] , INIT_43[ 31 :   0]};
    RAM[ 537] <= {INITP_08[103 : 100] , INIT_43[ 63 :  32]};
    RAM[ 538] <= {INITP_08[107 : 104] , INIT_43[ 95 :  64]};
    RAM[ 539] <= {INITP_08[111 : 108] , INIT_43[127 :  96]};
    RAM[ 540] <= {INITP_08[115 : 112] , INIT_43[159 : 128]};
    RAM[ 541] <= {INITP_08[119 : 116] , INIT_43[191 : 160]};
    RAM[ 542] <= {INITP_08[123 : 120] , INIT_43[223 : 192]};
    RAM[ 543] <= {INITP_08[127 : 124] , INIT_43[255 : 224]};
    RAM[ 544] <= {INITP_08[131 : 128] , INIT_44[ 31 :   0]};
    RAM[ 545] <= {INITP_08[135 : 132] , INIT_44[ 63 :  32]};
    RAM[ 546] <= {INITP_08[139 : 136] , INIT_44[ 95 :  64]};
    RAM[ 547] <= {INITP_08[143 : 140] , INIT_44[127 :  96]};
    RAM[ 548] <= {INITP_08[147 : 144] , INIT_44[159 : 128]};
    RAM[ 549] <= {INITP_08[151 : 148] , INIT_44[191 : 160]};
    RAM[ 550] <= {INITP_08[155 : 152] , INIT_44[223 : 192]};
    RAM[ 551] <= {INITP_08[159 : 156] , INIT_44[255 : 224]};
    RAM[ 552] <= {INITP_08[163 : 160] , INIT_45[ 31 :   0]};
    RAM[ 553] <= {INITP_08[167 : 164] , INIT_45[ 63 :  32]};
    RAM[ 554] <= {INITP_08[171 : 168] , INIT_45[ 95 :  64]};
    RAM[ 555] <= {INITP_08[175 : 172] , INIT_45[127 :  96]};
    RAM[ 556] <= {INITP_08[179 : 176] , INIT_45[159 : 128]};
    RAM[ 557] <= {INITP_08[183 : 180] , INIT_45[191 : 160]};
    RAM[ 558] <= {INITP_08[187 : 184] , INIT_45[223 : 192]};
    RAM[ 559] <= {INITP_08[191 : 188] , INIT_45[255 : 224]};
    RAM[ 560] <= {INITP_08[195 : 192] , INIT_46[ 31 :   0]};
    RAM[ 561] <= {INITP_08[199 : 196] , INIT_46[ 63 :  32]};
    RAM[ 562] <= {INITP_08[203 : 200] , INIT_46[ 95 :  64]};
    RAM[ 563] <= {INITP_08[207 : 204] , INIT_46[127 :  96]};
    RAM[ 564] <= {INITP_08[211 : 208] , INIT_46[159 : 128]};
    RAM[ 565] <= {INITP_08[215 : 212] , INIT_46[191 : 160]};
    RAM[ 566] <= {INITP_08[219 : 216] , INIT_46[223 : 192]};
    RAM[ 567] <= {INITP_08[223 : 220] , INIT_46[255 : 224]};
    RAM[ 568] <= {INITP_08[227 : 224] , INIT_47[ 31 :   0]};
    RAM[ 569] <= {INITP_08[231 : 228] , INIT_47[ 63 :  32]};
    RAM[ 570] <= {INITP_08[235 : 232] , INIT_47[ 95 :  64]};
    RAM[ 571] <= {INITP_08[239 : 236] , INIT_47[127 :  96]};
    RAM[ 572] <= {INITP_08[243 : 240] , INIT_47[159 : 128]};
    RAM[ 573] <= {INITP_08[247 : 244] , INIT_47[191 : 160]};
    RAM[ 574] <= {INITP_08[251 : 248] , INIT_47[223 : 192]};
    RAM[ 575] <= {INITP_08[255 : 252] , INIT_47[255 : 224]};
    RAM[ 576] <= {INITP_09[  3 :   0] , INIT_48[ 31 :   0]};
    RAM[ 577] <= {INITP_09[  7 :   4] , INIT_48[ 63 :  32]};
    RAM[ 578] <= {INITP_09[ 11 :   8] , INIT_48[ 95 :  64]};
    RAM[ 579] <= {INITP_09[ 15 :  12] , INIT_48[127 :  96]};
    RAM[ 580] <= {INITP_09[ 19 :  16] , INIT_48[159 : 128]};
    RAM[ 581] <= {INITP_09[ 23 :  20] , INIT_48[191 : 160]};
    RAM[ 582] <= {INITP_09[ 27 :  24] , INIT_48[223 : 192]};
    RAM[ 583] <= {INITP_09[ 31 :  28] , INIT_48[255 : 224]};
    RAM[ 584] <= {INITP_09[ 35 :  32] , INIT_49[ 31 :   0]};
    RAM[ 585] <= {INITP_09[ 39 :  36] , INIT_49[ 63 :  32]};
    RAM[ 586] <= {INITP_09[ 43 :  40] , INIT_49[ 95 :  64]};
    RAM[ 587] <= {INITP_09[ 47 :  44] , INIT_49[127 :  96]};
    RAM[ 588] <= {INITP_09[ 51 :  48] , INIT_49[159 : 128]};
    RAM[ 589] <= {INITP_09[ 55 :  52] , INIT_49[191 : 160]};
    RAM[ 590] <= {INITP_09[ 59 :  56] , INIT_49[223 : 192]};
    RAM[ 591] <= {INITP_09[ 63 :  60] , INIT_49[255 : 224]};
    RAM[ 592] <= {INITP_09[ 67 :  64] , INIT_4A[ 31 :   0]};
    RAM[ 593] <= {INITP_09[ 71 :  68] , INIT_4A[ 63 :  32]};
    RAM[ 594] <= {INITP_09[ 75 :  72] , INIT_4A[ 95 :  64]};
    RAM[ 595] <= {INITP_09[ 79 :  76] , INIT_4A[127 :  96]};
    RAM[ 596] <= {INITP_09[ 83 :  80] , INIT_4A[159 : 128]};
    RAM[ 597] <= {INITP_09[ 87 :  84] , INIT_4A[191 : 160]};
    RAM[ 598] <= {INITP_09[ 91 :  88] , INIT_4A[223 : 192]};
    RAM[ 599] <= {INITP_09[ 95 :  92] , INIT_4A[255 : 224]};
    RAM[ 600] <= {INITP_09[ 99 :  96] , INIT_4B[ 31 :   0]};
    RAM[ 601] <= {INITP_09[103 : 100] , INIT_4B[ 63 :  32]};
    RAM[ 602] <= {INITP_09[107 : 104] , INIT_4B[ 95 :  64]};
    RAM[ 603] <= {INITP_09[111 : 108] , INIT_4B[127 :  96]};
    RAM[ 604] <= {INITP_09[115 : 112] , INIT_4B[159 : 128]};
    RAM[ 605] <= {INITP_09[119 : 116] , INIT_4B[191 : 160]};
    RAM[ 606] <= {INITP_09[123 : 120] , INIT_4B[223 : 192]};
    RAM[ 607] <= {INITP_09[127 : 124] , INIT_4B[255 : 224]};
    RAM[ 608] <= {INITP_09[131 : 128] , INIT_4C[ 31 :   0]};
    RAM[ 609] <= {INITP_09[135 : 132] , INIT_4C[ 63 :  32]};
    RAM[ 610] <= {INITP_09[139 : 136] , INIT_4C[ 95 :  64]};
    RAM[ 611] <= {INITP_09[143 : 140] , INIT_4C[127 :  96]};
    RAM[ 612] <= {INITP_09[147 : 144] , INIT_4C[159 : 128]};
    RAM[ 613] <= {INITP_09[151 : 148] , INIT_4C[191 : 160]};
    RAM[ 614] <= {INITP_09[155 : 152] , INIT_4C[223 : 192]};
    RAM[ 615] <= {INITP_09[159 : 156] , INIT_4C[255 : 224]};
    RAM[ 616] <= {INITP_09[163 : 160] , INIT_4D[ 31 :   0]};
    RAM[ 617] <= {INITP_09[167 : 164] , INIT_4D[ 63 :  32]};
    RAM[ 618] <= {INITP_09[171 : 168] , INIT_4D[ 95 :  64]};
    RAM[ 619] <= {INITP_09[175 : 172] , INIT_4D[127 :  96]};
    RAM[ 620] <= {INITP_09[179 : 176] , INIT_4D[159 : 128]};
    RAM[ 621] <= {INITP_09[183 : 180] , INIT_4D[191 : 160]};
    RAM[ 622] <= {INITP_09[187 : 184] , INIT_4D[223 : 192]};
    RAM[ 623] <= {INITP_09[191 : 188] , INIT_4D[255 : 224]};
    RAM[ 624] <= {INITP_09[195 : 192] , INIT_4E[ 31 :   0]};
    RAM[ 625] <= {INITP_09[199 : 196] , INIT_4E[ 63 :  32]};
    RAM[ 626] <= {INITP_09[203 : 200] , INIT_4E[ 95 :  64]};
    RAM[ 627] <= {INITP_09[207 : 204] , INIT_4E[127 :  96]};
    RAM[ 628] <= {INITP_09[211 : 208] , INIT_4E[159 : 128]};
    RAM[ 629] <= {INITP_09[215 : 212] , INIT_4E[191 : 160]};
    RAM[ 630] <= {INITP_09[219 : 216] , INIT_4E[223 : 192]};
    RAM[ 631] <= {INITP_09[223 : 220] , INIT_4E[255 : 224]};
    RAM[ 632] <= {INITP_09[227 : 224] , INIT_4F[ 31 :   0]};
    RAM[ 633] <= {INITP_09[231 : 228] , INIT_4F[ 63 :  32]};
    RAM[ 634] <= {INITP_09[235 : 232] , INIT_4F[ 95 :  64]};
    RAM[ 635] <= {INITP_09[239 : 236] , INIT_4F[127 :  96]};
    RAM[ 636] <= {INITP_09[243 : 240] , INIT_4F[159 : 128]};
    RAM[ 637] <= {INITP_09[247 : 244] , INIT_4F[191 : 160]};
    RAM[ 638] <= {INITP_09[251 : 248] , INIT_4F[223 : 192]};
    RAM[ 639] <= {INITP_09[255 : 252] , INIT_4F[255 : 224]};
    RAM[ 640] <= {INITP_0A[  3 :   0] , INIT_50[ 31 :   0]};
    RAM[ 641] <= {INITP_0A[  7 :   4] , INIT_50[ 63 :  32]};
    RAM[ 642] <= {INITP_0A[ 11 :   8] , INIT_50[ 95 :  64]};
    RAM[ 643] <= {INITP_0A[ 15 :  12] , INIT_50[127 :  96]};
    RAM[ 644] <= {INITP_0A[ 19 :  16] , INIT_50[159 : 128]};
    RAM[ 645] <= {INITP_0A[ 23 :  20] , INIT_50[191 : 160]};
    RAM[ 646] <= {INITP_0A[ 27 :  24] , INIT_50[223 : 192]};
    RAM[ 647] <= {INITP_0A[ 31 :  28] , INIT_50[255 : 224]};
    RAM[ 648] <= {INITP_0A[ 35 :  32] , INIT_51[ 31 :   0]};
    RAM[ 649] <= {INITP_0A[ 39 :  36] , INIT_51[ 63 :  32]};
    RAM[ 650] <= {INITP_0A[ 43 :  40] , INIT_51[ 95 :  64]};
    RAM[ 651] <= {INITP_0A[ 47 :  44] , INIT_51[127 :  96]};
    RAM[ 652] <= {INITP_0A[ 51 :  48] , INIT_51[159 : 128]};
    RAM[ 653] <= {INITP_0A[ 55 :  52] , INIT_51[191 : 160]};
    RAM[ 654] <= {INITP_0A[ 59 :  56] , INIT_51[223 : 192]};
    RAM[ 655] <= {INITP_0A[ 63 :  60] , INIT_51[255 : 224]};
    RAM[ 656] <= {INITP_0A[ 67 :  64] , INIT_52[ 31 :   0]};
    RAM[ 657] <= {INITP_0A[ 71 :  68] , INIT_52[ 63 :  32]};
    RAM[ 658] <= {INITP_0A[ 75 :  72] , INIT_52[ 95 :  64]};
    RAM[ 659] <= {INITP_0A[ 79 :  76] , INIT_52[127 :  96]};
    RAM[ 660] <= {INITP_0A[ 83 :  80] , INIT_52[159 : 128]};
    RAM[ 661] <= {INITP_0A[ 87 :  84] , INIT_52[191 : 160]};
    RAM[ 662] <= {INITP_0A[ 91 :  88] , INIT_52[223 : 192]};
    RAM[ 663] <= {INITP_0A[ 95 :  92] , INIT_52[255 : 224]};
    RAM[ 664] <= {INITP_0A[ 99 :  96] , INIT_53[ 31 :   0]};
    RAM[ 665] <= {INITP_0A[103 : 100] , INIT_53[ 63 :  32]};
    RAM[ 666] <= {INITP_0A[107 : 104] , INIT_53[ 95 :  64]};
    RAM[ 667] <= {INITP_0A[111 : 108] , INIT_53[127 :  96]};
    RAM[ 668] <= {INITP_0A[115 : 112] , INIT_53[159 : 128]};
    RAM[ 669] <= {INITP_0A[119 : 116] , INIT_53[191 : 160]};
    RAM[ 670] <= {INITP_0A[123 : 120] , INIT_53[223 : 192]};
    RAM[ 671] <= {INITP_0A[127 : 124] , INIT_53[255 : 224]};
    RAM[ 672] <= {INITP_0A[131 : 128] , INIT_54[ 31 :   0]};
    RAM[ 673] <= {INITP_0A[135 : 132] , INIT_54[ 63 :  32]};
    RAM[ 674] <= {INITP_0A[139 : 136] , INIT_54[ 95 :  64]};
    RAM[ 675] <= {INITP_0A[143 : 140] , INIT_54[127 :  96]};
    RAM[ 676] <= {INITP_0A[147 : 144] , INIT_54[159 : 128]};
    RAM[ 677] <= {INITP_0A[151 : 148] , INIT_54[191 : 160]};
    RAM[ 678] <= {INITP_0A[155 : 152] , INIT_54[223 : 192]};
    RAM[ 679] <= {INITP_0A[159 : 156] , INIT_54[255 : 224]};
    RAM[ 680] <= {INITP_0A[163 : 160] , INIT_55[ 31 :   0]};
    RAM[ 681] <= {INITP_0A[167 : 164] , INIT_55[ 63 :  32]};
    RAM[ 682] <= {INITP_0A[171 : 168] , INIT_55[ 95 :  64]};
    RAM[ 683] <= {INITP_0A[175 : 172] , INIT_55[127 :  96]};
    RAM[ 684] <= {INITP_0A[179 : 176] , INIT_55[159 : 128]};
    RAM[ 685] <= {INITP_0A[183 : 180] , INIT_55[191 : 160]};
    RAM[ 686] <= {INITP_0A[187 : 184] , INIT_55[223 : 192]};
    RAM[ 687] <= {INITP_0A[191 : 188] , INIT_55[255 : 224]};
    RAM[ 688] <= {INITP_0A[195 : 192] , INIT_56[ 31 :   0]};
    RAM[ 689] <= {INITP_0A[199 : 196] , INIT_56[ 63 :  32]};
    RAM[ 690] <= {INITP_0A[203 : 200] , INIT_56[ 95 :  64]};
    RAM[ 691] <= {INITP_0A[207 : 204] , INIT_56[127 :  96]};
    RAM[ 692] <= {INITP_0A[211 : 208] , INIT_56[159 : 128]};
    RAM[ 693] <= {INITP_0A[215 : 212] , INIT_56[191 : 160]};
    RAM[ 694] <= {INITP_0A[219 : 216] , INIT_56[223 : 192]};
    RAM[ 695] <= {INITP_0A[223 : 220] , INIT_56[255 : 224]};
    RAM[ 696] <= {INITP_0A[227 : 224] , INIT_57[ 31 :   0]};
    RAM[ 697] <= {INITP_0A[231 : 228] , INIT_57[ 63 :  32]};
    RAM[ 698] <= {INITP_0A[235 : 232] , INIT_57[ 95 :  64]};
    RAM[ 699] <= {INITP_0A[239 : 236] , INIT_57[127 :  96]};
    RAM[ 700] <= {INITP_0A[243 : 240] , INIT_57[159 : 128]};
    RAM[ 701] <= {INITP_0A[247 : 244] , INIT_57[191 : 160]};
    RAM[ 702] <= {INITP_0A[251 : 248] , INIT_57[223 : 192]};
    RAM[ 703] <= {INITP_0A[255 : 252] , INIT_57[255 : 224]};
    RAM[ 704] <= {INITP_0B[  3 :   0] , INIT_58[ 31 :   0]};
    RAM[ 705] <= {INITP_0B[  7 :   4] , INIT_58[ 63 :  32]};
    RAM[ 706] <= {INITP_0B[ 11 :   8] , INIT_58[ 95 :  64]};
    RAM[ 707] <= {INITP_0B[ 15 :  12] , INIT_58[127 :  96]};
    RAM[ 708] <= {INITP_0B[ 19 :  16] , INIT_58[159 : 128]};
    RAM[ 709] <= {INITP_0B[ 23 :  20] , INIT_58[191 : 160]};
    RAM[ 710] <= {INITP_0B[ 27 :  24] , INIT_58[223 : 192]};
    RAM[ 711] <= {INITP_0B[ 31 :  28] , INIT_58[255 : 224]};
    RAM[ 712] <= {INITP_0B[ 35 :  32] , INIT_59[ 31 :   0]};
    RAM[ 713] <= {INITP_0B[ 39 :  36] , INIT_59[ 63 :  32]};
    RAM[ 714] <= {INITP_0B[ 43 :  40] , INIT_59[ 95 :  64]};
    RAM[ 715] <= {INITP_0B[ 47 :  44] , INIT_59[127 :  96]};
    RAM[ 716] <= {INITP_0B[ 51 :  48] , INIT_59[159 : 128]};
    RAM[ 717] <= {INITP_0B[ 55 :  52] , INIT_59[191 : 160]};
    RAM[ 718] <= {INITP_0B[ 59 :  56] , INIT_59[223 : 192]};
    RAM[ 719] <= {INITP_0B[ 63 :  60] , INIT_59[255 : 224]};
    RAM[ 720] <= {INITP_0B[ 67 :  64] , INIT_5A[ 31 :   0]};
    RAM[ 721] <= {INITP_0B[ 71 :  68] , INIT_5A[ 63 :  32]};
    RAM[ 722] <= {INITP_0B[ 75 :  72] , INIT_5A[ 95 :  64]};
    RAM[ 723] <= {INITP_0B[ 79 :  76] , INIT_5A[127 :  96]};
    RAM[ 724] <= {INITP_0B[ 83 :  80] , INIT_5A[159 : 128]};
    RAM[ 725] <= {INITP_0B[ 87 :  84] , INIT_5A[191 : 160]};
    RAM[ 726] <= {INITP_0B[ 91 :  88] , INIT_5A[223 : 192]};
    RAM[ 727] <= {INITP_0B[ 95 :  92] , INIT_5A[255 : 224]};
    RAM[ 728] <= {INITP_0B[ 99 :  96] , INIT_5B[ 31 :   0]};
    RAM[ 729] <= {INITP_0B[103 : 100] , INIT_5B[ 63 :  32]};
    RAM[ 730] <= {INITP_0B[107 : 104] , INIT_5B[ 95 :  64]};
    RAM[ 731] <= {INITP_0B[111 : 108] , INIT_5B[127 :  96]};
    RAM[ 732] <= {INITP_0B[115 : 112] , INIT_5B[159 : 128]};
    RAM[ 733] <= {INITP_0B[119 : 116] , INIT_5B[191 : 160]};
    RAM[ 734] <= {INITP_0B[123 : 120] , INIT_5B[223 : 192]};
    RAM[ 735] <= {INITP_0B[127 : 124] , INIT_5B[255 : 224]};
    RAM[ 736] <= {INITP_0B[131 : 128] , INIT_5C[ 31 :   0]};
    RAM[ 737] <= {INITP_0B[135 : 132] , INIT_5C[ 63 :  32]};
    RAM[ 738] <= {INITP_0B[139 : 136] , INIT_5C[ 95 :  64]};
    RAM[ 739] <= {INITP_0B[143 : 140] , INIT_5C[127 :  96]};
    RAM[ 740] <= {INITP_0B[147 : 144] , INIT_5C[159 : 128]};
    RAM[ 741] <= {INITP_0B[151 : 148] , INIT_5C[191 : 160]};
    RAM[ 742] <= {INITP_0B[155 : 152] , INIT_5C[223 : 192]};
    RAM[ 743] <= {INITP_0B[159 : 156] , INIT_5C[255 : 224]};
    RAM[ 744] <= {INITP_0B[163 : 160] , INIT_5D[ 31 :   0]};
    RAM[ 745] <= {INITP_0B[167 : 164] , INIT_5D[ 63 :  32]};
    RAM[ 746] <= {INITP_0B[171 : 168] , INIT_5D[ 95 :  64]};
    RAM[ 747] <= {INITP_0B[175 : 172] , INIT_5D[127 :  96]};
    RAM[ 748] <= {INITP_0B[179 : 176] , INIT_5D[159 : 128]};
    RAM[ 749] <= {INITP_0B[183 : 180] , INIT_5D[191 : 160]};
    RAM[ 750] <= {INITP_0B[187 : 184] , INIT_5D[223 : 192]};
    RAM[ 751] <= {INITP_0B[191 : 188] , INIT_5D[255 : 224]};
    RAM[ 752] <= {INITP_0B[195 : 192] , INIT_5E[ 31 :   0]};
    RAM[ 753] <= {INITP_0B[199 : 196] , INIT_5E[ 63 :  32]};
    RAM[ 754] <= {INITP_0B[203 : 200] , INIT_5E[ 95 :  64]};
    RAM[ 755] <= {INITP_0B[207 : 204] , INIT_5E[127 :  96]};
    RAM[ 756] <= {INITP_0B[211 : 208] , INIT_5E[159 : 128]};
    RAM[ 757] <= {INITP_0B[215 : 212] , INIT_5E[191 : 160]};
    RAM[ 758] <= {INITP_0B[219 : 216] , INIT_5E[223 : 192]};
    RAM[ 759] <= {INITP_0B[223 : 220] , INIT_5E[255 : 224]};
    RAM[ 760] <= {INITP_0B[227 : 224] , INIT_5F[ 31 :   0]};
    RAM[ 761] <= {INITP_0B[231 : 228] , INIT_5F[ 63 :  32]};
    RAM[ 762] <= {INITP_0B[235 : 232] , INIT_5F[ 95 :  64]};
    RAM[ 763] <= {INITP_0B[239 : 236] , INIT_5F[127 :  96]};
    RAM[ 764] <= {INITP_0B[243 : 240] , INIT_5F[159 : 128]};
    RAM[ 765] <= {INITP_0B[247 : 244] , INIT_5F[191 : 160]};
    RAM[ 766] <= {INITP_0B[251 : 248] , INIT_5F[223 : 192]};
    RAM[ 767] <= {INITP_0B[255 : 252] , INIT_5F[255 : 224]};
    RAM[ 768] <= {INITP_0C[  3 :   0] , INIT_60[ 31 :   0]};
    RAM[ 769] <= {INITP_0C[  7 :   4] , INIT_60[ 63 :  32]};
    RAM[ 770] <= {INITP_0C[ 11 :   8] , INIT_60[ 95 :  64]};
    RAM[ 771] <= {INITP_0C[ 15 :  12] , INIT_60[127 :  96]};
    RAM[ 772] <= {INITP_0C[ 19 :  16] , INIT_60[159 : 128]};
    RAM[ 773] <= {INITP_0C[ 23 :  20] , INIT_60[191 : 160]};
    RAM[ 774] <= {INITP_0C[ 27 :  24] , INIT_60[223 : 192]};
    RAM[ 775] <= {INITP_0C[ 31 :  28] , INIT_60[255 : 224]};
    RAM[ 776] <= {INITP_0C[ 35 :  32] , INIT_61[ 31 :   0]};
    RAM[ 777] <= {INITP_0C[ 39 :  36] , INIT_61[ 63 :  32]};
    RAM[ 778] <= {INITP_0C[ 43 :  40] , INIT_61[ 95 :  64]};
    RAM[ 779] <= {INITP_0C[ 47 :  44] , INIT_61[127 :  96]};
    RAM[ 780] <= {INITP_0C[ 51 :  48] , INIT_61[159 : 128]};
    RAM[ 781] <= {INITP_0C[ 55 :  52] , INIT_61[191 : 160]};
    RAM[ 782] <= {INITP_0C[ 59 :  56] , INIT_61[223 : 192]};
    RAM[ 783] <= {INITP_0C[ 63 :  60] , INIT_61[255 : 224]};
    RAM[ 784] <= {INITP_0C[ 67 :  64] , INIT_62[ 31 :   0]};
    RAM[ 785] <= {INITP_0C[ 71 :  68] , INIT_62[ 63 :  32]};
    RAM[ 786] <= {INITP_0C[ 75 :  72] , INIT_62[ 95 :  64]};
    RAM[ 787] <= {INITP_0C[ 79 :  76] , INIT_62[127 :  96]};
    RAM[ 788] <= {INITP_0C[ 83 :  80] , INIT_62[159 : 128]};
    RAM[ 789] <= {INITP_0C[ 87 :  84] , INIT_62[191 : 160]};
    RAM[ 790] <= {INITP_0C[ 91 :  88] , INIT_62[223 : 192]};
    RAM[ 791] <= {INITP_0C[ 95 :  92] , INIT_62[255 : 224]};
    RAM[ 792] <= {INITP_0C[ 99 :  96] , INIT_63[ 31 :   0]};
    RAM[ 793] <= {INITP_0C[103 : 100] , INIT_63[ 63 :  32]};
    RAM[ 794] <= {INITP_0C[107 : 104] , INIT_63[ 95 :  64]};
    RAM[ 795] <= {INITP_0C[111 : 108] , INIT_63[127 :  96]};
    RAM[ 796] <= {INITP_0C[115 : 112] , INIT_63[159 : 128]};
    RAM[ 797] <= {INITP_0C[119 : 116] , INIT_63[191 : 160]};
    RAM[ 798] <= {INITP_0C[123 : 120] , INIT_63[223 : 192]};
    RAM[ 799] <= {INITP_0C[127 : 124] , INIT_63[255 : 224]};
    RAM[ 800] <= {INITP_0C[131 : 128] , INIT_64[ 31 :   0]};
    RAM[ 801] <= {INITP_0C[135 : 132] , INIT_64[ 63 :  32]};
    RAM[ 802] <= {INITP_0C[139 : 136] , INIT_64[ 95 :  64]};
    RAM[ 803] <= {INITP_0C[143 : 140] , INIT_64[127 :  96]};
    RAM[ 804] <= {INITP_0C[147 : 144] , INIT_64[159 : 128]};
    RAM[ 805] <= {INITP_0C[151 : 148] , INIT_64[191 : 160]};
    RAM[ 806] <= {INITP_0C[155 : 152] , INIT_64[223 : 192]};
    RAM[ 807] <= {INITP_0C[159 : 156] , INIT_64[255 : 224]};
    RAM[ 808] <= {INITP_0C[163 : 160] , INIT_65[ 31 :   0]};
    RAM[ 809] <= {INITP_0C[167 : 164] , INIT_65[ 63 :  32]};
    RAM[ 810] <= {INITP_0C[171 : 168] , INIT_65[ 95 :  64]};
    RAM[ 811] <= {INITP_0C[175 : 172] , INIT_65[127 :  96]};
    RAM[ 812] <= {INITP_0C[179 : 176] , INIT_65[159 : 128]};
    RAM[ 813] <= {INITP_0C[183 : 180] , INIT_65[191 : 160]};
    RAM[ 814] <= {INITP_0C[187 : 184] , INIT_65[223 : 192]};
    RAM[ 815] <= {INITP_0C[191 : 188] , INIT_65[255 : 224]};
    RAM[ 816] <= {INITP_0C[195 : 192] , INIT_66[ 31 :   0]};
    RAM[ 817] <= {INITP_0C[199 : 196] , INIT_66[ 63 :  32]};
    RAM[ 818] <= {INITP_0C[203 : 200] , INIT_66[ 95 :  64]};
    RAM[ 819] <= {INITP_0C[207 : 204] , INIT_66[127 :  96]};
    RAM[ 820] <= {INITP_0C[211 : 208] , INIT_66[159 : 128]};
    RAM[ 821] <= {INITP_0C[215 : 212] , INIT_66[191 : 160]};
    RAM[ 822] <= {INITP_0C[219 : 216] , INIT_66[223 : 192]};
    RAM[ 823] <= {INITP_0C[223 : 220] , INIT_66[255 : 224]};
    RAM[ 824] <= {INITP_0C[227 : 224] , INIT_67[ 31 :   0]};
    RAM[ 825] <= {INITP_0C[231 : 228] , INIT_67[ 63 :  32]};
    RAM[ 826] <= {INITP_0C[235 : 232] , INIT_67[ 95 :  64]};
    RAM[ 827] <= {INITP_0C[239 : 236] , INIT_67[127 :  96]};
    RAM[ 828] <= {INITP_0C[243 : 240] , INIT_67[159 : 128]};
    RAM[ 829] <= {INITP_0C[247 : 244] , INIT_67[191 : 160]};
    RAM[ 830] <= {INITP_0C[251 : 248] , INIT_67[223 : 192]};
    RAM[ 831] <= {INITP_0C[255 : 252] , INIT_67[255 : 224]};
    RAM[ 832] <= {INITP_0D[  3 :   0] , INIT_68[ 31 :   0]};
    RAM[ 833] <= {INITP_0D[  7 :   4] , INIT_68[ 63 :  32]};
    RAM[ 834] <= {INITP_0D[ 11 :   8] , INIT_68[ 95 :  64]};
    RAM[ 835] <= {INITP_0D[ 15 :  12] , INIT_68[127 :  96]};
    RAM[ 836] <= {INITP_0D[ 19 :  16] , INIT_68[159 : 128]};
    RAM[ 837] <= {INITP_0D[ 23 :  20] , INIT_68[191 : 160]};
    RAM[ 838] <= {INITP_0D[ 27 :  24] , INIT_68[223 : 192]};
    RAM[ 839] <= {INITP_0D[ 31 :  28] , INIT_68[255 : 224]};
    RAM[ 840] <= {INITP_0D[ 35 :  32] , INIT_69[ 31 :   0]};
    RAM[ 841] <= {INITP_0D[ 39 :  36] , INIT_69[ 63 :  32]};
    RAM[ 842] <= {INITP_0D[ 43 :  40] , INIT_69[ 95 :  64]};
    RAM[ 843] <= {INITP_0D[ 47 :  44] , INIT_69[127 :  96]};
    RAM[ 844] <= {INITP_0D[ 51 :  48] , INIT_69[159 : 128]};
    RAM[ 845] <= {INITP_0D[ 55 :  52] , INIT_69[191 : 160]};
    RAM[ 846] <= {INITP_0D[ 59 :  56] , INIT_69[223 : 192]};
    RAM[ 847] <= {INITP_0D[ 63 :  60] , INIT_69[255 : 224]};
    RAM[ 848] <= {INITP_0D[ 67 :  64] , INIT_6A[ 31 :   0]};
    RAM[ 849] <= {INITP_0D[ 71 :  68] , INIT_6A[ 63 :  32]};
    RAM[ 850] <= {INITP_0D[ 75 :  72] , INIT_6A[ 95 :  64]};
    RAM[ 851] <= {INITP_0D[ 79 :  76] , INIT_6A[127 :  96]};
    RAM[ 852] <= {INITP_0D[ 83 :  80] , INIT_6A[159 : 128]};
    RAM[ 853] <= {INITP_0D[ 87 :  84] , INIT_6A[191 : 160]};
    RAM[ 854] <= {INITP_0D[ 91 :  88] , INIT_6A[223 : 192]};
    RAM[ 855] <= {INITP_0D[ 95 :  92] , INIT_6A[255 : 224]};
    RAM[ 856] <= {INITP_0D[ 99 :  96] , INIT_6B[ 31 :   0]};
    RAM[ 857] <= {INITP_0D[103 : 100] , INIT_6B[ 63 :  32]};
    RAM[ 858] <= {INITP_0D[107 : 104] , INIT_6B[ 95 :  64]};
    RAM[ 859] <= {INITP_0D[111 : 108] , INIT_6B[127 :  96]};
    RAM[ 860] <= {INITP_0D[115 : 112] , INIT_6B[159 : 128]};
    RAM[ 861] <= {INITP_0D[119 : 116] , INIT_6B[191 : 160]};
    RAM[ 862] <= {INITP_0D[123 : 120] , INIT_6B[223 : 192]};
    RAM[ 863] <= {INITP_0D[127 : 124] , INIT_6B[255 : 224]};
    RAM[ 864] <= {INITP_0D[131 : 128] , INIT_6C[ 31 :   0]};
    RAM[ 865] <= {INITP_0D[135 : 132] , INIT_6C[ 63 :  32]};
    RAM[ 866] <= {INITP_0D[139 : 136] , INIT_6C[ 95 :  64]};
    RAM[ 867] <= {INITP_0D[143 : 140] , INIT_6C[127 :  96]};
    RAM[ 868] <= {INITP_0D[147 : 144] , INIT_6C[159 : 128]};
    RAM[ 869] <= {INITP_0D[151 : 148] , INIT_6C[191 : 160]};
    RAM[ 870] <= {INITP_0D[155 : 152] , INIT_6C[223 : 192]};
    RAM[ 871] <= {INITP_0D[159 : 156] , INIT_6C[255 : 224]};
    RAM[ 872] <= {INITP_0D[163 : 160] , INIT_6D[ 31 :   0]};
    RAM[ 873] <= {INITP_0D[167 : 164] , INIT_6D[ 63 :  32]};
    RAM[ 874] <= {INITP_0D[171 : 168] , INIT_6D[ 95 :  64]};
    RAM[ 875] <= {INITP_0D[175 : 172] , INIT_6D[127 :  96]};
    RAM[ 876] <= {INITP_0D[179 : 176] , INIT_6D[159 : 128]};
    RAM[ 877] <= {INITP_0D[183 : 180] , INIT_6D[191 : 160]};
    RAM[ 878] <= {INITP_0D[187 : 184] , INIT_6D[223 : 192]};
    RAM[ 879] <= {INITP_0D[191 : 188] , INIT_6D[255 : 224]};
    RAM[ 880] <= {INITP_0D[195 : 192] , INIT_6E[ 31 :   0]};
    RAM[ 881] <= {INITP_0D[199 : 196] , INIT_6E[ 63 :  32]};
    RAM[ 882] <= {INITP_0D[203 : 200] , INIT_6E[ 95 :  64]};
    RAM[ 883] <= {INITP_0D[207 : 204] , INIT_6E[127 :  96]};
    RAM[ 884] <= {INITP_0D[211 : 208] , INIT_6E[159 : 128]};
    RAM[ 885] <= {INITP_0D[215 : 212] , INIT_6E[191 : 160]};
    RAM[ 886] <= {INITP_0D[219 : 216] , INIT_6E[223 : 192]};
    RAM[ 887] <= {INITP_0D[223 : 220] , INIT_6E[255 : 224]};
    RAM[ 888] <= {INITP_0D[227 : 224] , INIT_6F[ 31 :   0]};
    RAM[ 889] <= {INITP_0D[231 : 228] , INIT_6F[ 63 :  32]};
    RAM[ 890] <= {INITP_0D[235 : 232] , INIT_6F[ 95 :  64]};
    RAM[ 891] <= {INITP_0D[239 : 236] , INIT_6F[127 :  96]};
    RAM[ 892] <= {INITP_0D[243 : 240] , INIT_6F[159 : 128]};
    RAM[ 893] <= {INITP_0D[247 : 244] , INIT_6F[191 : 160]};
    RAM[ 894] <= {INITP_0D[251 : 248] , INIT_6F[223 : 192]};
    RAM[ 895] <= {INITP_0D[255 : 252] , INIT_6F[255 : 224]};
    RAM[ 896] <= {INITP_0E[  3 :   0] , INIT_70[ 31 :   0]};
    RAM[ 897] <= {INITP_0E[  7 :   4] , INIT_70[ 63 :  32]};
    RAM[ 898] <= {INITP_0E[ 11 :   8] , INIT_70[ 95 :  64]};
    RAM[ 899] <= {INITP_0E[ 15 :  12] , INIT_70[127 :  96]};
    RAM[ 900] <= {INITP_0E[ 19 :  16] , INIT_70[159 : 128]};
    RAM[ 901] <= {INITP_0E[ 23 :  20] , INIT_70[191 : 160]};
    RAM[ 902] <= {INITP_0E[ 27 :  24] , INIT_70[223 : 192]};
    RAM[ 903] <= {INITP_0E[ 31 :  28] , INIT_70[255 : 224]};
    RAM[ 904] <= {INITP_0E[ 35 :  32] , INIT_71[ 31 :   0]};
    RAM[ 905] <= {INITP_0E[ 39 :  36] , INIT_71[ 63 :  32]};
    RAM[ 906] <= {INITP_0E[ 43 :  40] , INIT_71[ 95 :  64]};
    RAM[ 907] <= {INITP_0E[ 47 :  44] , INIT_71[127 :  96]};
    RAM[ 908] <= {INITP_0E[ 51 :  48] , INIT_71[159 : 128]};
    RAM[ 909] <= {INITP_0E[ 55 :  52] , INIT_71[191 : 160]};
    RAM[ 910] <= {INITP_0E[ 59 :  56] , INIT_71[223 : 192]};
    RAM[ 911] <= {INITP_0E[ 63 :  60] , INIT_71[255 : 224]};
    RAM[ 912] <= {INITP_0E[ 67 :  64] , INIT_72[ 31 :   0]};
    RAM[ 913] <= {INITP_0E[ 71 :  68] , INIT_72[ 63 :  32]};
    RAM[ 914] <= {INITP_0E[ 75 :  72] , INIT_72[ 95 :  64]};
    RAM[ 915] <= {INITP_0E[ 79 :  76] , INIT_72[127 :  96]};
    RAM[ 916] <= {INITP_0E[ 83 :  80] , INIT_72[159 : 128]};
    RAM[ 917] <= {INITP_0E[ 87 :  84] , INIT_72[191 : 160]};
    RAM[ 918] <= {INITP_0E[ 91 :  88] , INIT_72[223 : 192]};
    RAM[ 919] <= {INITP_0E[ 95 :  92] , INIT_72[255 : 224]};
    RAM[ 920] <= {INITP_0E[ 99 :  96] , INIT_73[ 31 :   0]};
    RAM[ 921] <= {INITP_0E[103 : 100] , INIT_73[ 63 :  32]};
    RAM[ 922] <= {INITP_0E[107 : 104] , INIT_73[ 95 :  64]};
    RAM[ 923] <= {INITP_0E[111 : 108] , INIT_73[127 :  96]};
    RAM[ 924] <= {INITP_0E[115 : 112] , INIT_73[159 : 128]};
    RAM[ 925] <= {INITP_0E[119 : 116] , INIT_73[191 : 160]};
    RAM[ 926] <= {INITP_0E[123 : 120] , INIT_73[223 : 192]};
    RAM[ 927] <= {INITP_0E[127 : 124] , INIT_73[255 : 224]};
    RAM[ 928] <= {INITP_0E[131 : 128] , INIT_74[ 31 :   0]};
    RAM[ 929] <= {INITP_0E[135 : 132] , INIT_74[ 63 :  32]};
    RAM[ 930] <= {INITP_0E[139 : 136] , INIT_74[ 95 :  64]};
    RAM[ 931] <= {INITP_0E[143 : 140] , INIT_74[127 :  96]};
    RAM[ 932] <= {INITP_0E[147 : 144] , INIT_74[159 : 128]};
    RAM[ 933] <= {INITP_0E[151 : 148] , INIT_74[191 : 160]};
    RAM[ 934] <= {INITP_0E[155 : 152] , INIT_74[223 : 192]};
    RAM[ 935] <= {INITP_0E[159 : 156] , INIT_74[255 : 224]};
    RAM[ 936] <= {INITP_0E[163 : 160] , INIT_75[ 31 :   0]};
    RAM[ 937] <= {INITP_0E[167 : 164] , INIT_75[ 63 :  32]};
    RAM[ 938] <= {INITP_0E[171 : 168] , INIT_75[ 95 :  64]};
    RAM[ 939] <= {INITP_0E[175 : 172] , INIT_75[127 :  96]};
    RAM[ 940] <= {INITP_0E[179 : 176] , INIT_75[159 : 128]};
    RAM[ 941] <= {INITP_0E[183 : 180] , INIT_75[191 : 160]};
    RAM[ 942] <= {INITP_0E[187 : 184] , INIT_75[223 : 192]};
    RAM[ 943] <= {INITP_0E[191 : 188] , INIT_75[255 : 224]};
    RAM[ 944] <= {INITP_0E[195 : 192] , INIT_76[ 31 :   0]};
    RAM[ 945] <= {INITP_0E[199 : 196] , INIT_76[ 63 :  32]};
    RAM[ 946] <= {INITP_0E[203 : 200] , INIT_76[ 95 :  64]};
    RAM[ 947] <= {INITP_0E[207 : 204] , INIT_76[127 :  96]};
    RAM[ 948] <= {INITP_0E[211 : 208] , INIT_76[159 : 128]};
    RAM[ 949] <= {INITP_0E[215 : 212] , INIT_76[191 : 160]};
    RAM[ 950] <= {INITP_0E[219 : 216] , INIT_76[223 : 192]};
    RAM[ 951] <= {INITP_0E[223 : 220] , INIT_76[255 : 224]};
    RAM[ 952] <= {INITP_0E[227 : 224] , INIT_77[ 31 :   0]};
    RAM[ 953] <= {INITP_0E[231 : 228] , INIT_77[ 63 :  32]};
    RAM[ 954] <= {INITP_0E[235 : 232] , INIT_77[ 95 :  64]};
    RAM[ 955] <= {INITP_0E[239 : 236] , INIT_77[127 :  96]};
    RAM[ 956] <= {INITP_0E[243 : 240] , INIT_77[159 : 128]};
    RAM[ 957] <= {INITP_0E[247 : 244] , INIT_77[191 : 160]};
    RAM[ 958] <= {INITP_0E[251 : 248] , INIT_77[223 : 192]};
    RAM[ 959] <= {INITP_0E[255 : 252] , INIT_77[255 : 224]};
    RAM[ 960] <= {INITP_0F[  3 :   0] , INIT_78[ 31 :   0]};
    RAM[ 961] <= {INITP_0F[  7 :   4] , INIT_78[ 63 :  32]};
    RAM[ 962] <= {INITP_0F[ 11 :   8] , INIT_78[ 95 :  64]};
    RAM[ 963] <= {INITP_0F[ 15 :  12] , INIT_78[127 :  96]};
    RAM[ 964] <= {INITP_0F[ 19 :  16] , INIT_78[159 : 128]};
    RAM[ 965] <= {INITP_0F[ 23 :  20] , INIT_78[191 : 160]};
    RAM[ 966] <= {INITP_0F[ 27 :  24] , INIT_78[223 : 192]};
    RAM[ 967] <= {INITP_0F[ 31 :  28] , INIT_78[255 : 224]};
    RAM[ 968] <= {INITP_0F[ 35 :  32] , INIT_79[ 31 :   0]};
    RAM[ 969] <= {INITP_0F[ 39 :  36] , INIT_79[ 63 :  32]};
    RAM[ 970] <= {INITP_0F[ 43 :  40] , INIT_79[ 95 :  64]};
    RAM[ 971] <= {INITP_0F[ 47 :  44] , INIT_79[127 :  96]};
    RAM[ 972] <= {INITP_0F[ 51 :  48] , INIT_79[159 : 128]};
    RAM[ 973] <= {INITP_0F[ 55 :  52] , INIT_79[191 : 160]};
    RAM[ 974] <= {INITP_0F[ 59 :  56] , INIT_79[223 : 192]};
    RAM[ 975] <= {INITP_0F[ 63 :  60] , INIT_79[255 : 224]};
    RAM[ 976] <= {INITP_0F[ 67 :  64] , INIT_7A[ 31 :   0]};
    RAM[ 977] <= {INITP_0F[ 71 :  68] , INIT_7A[ 63 :  32]};
    RAM[ 978] <= {INITP_0F[ 75 :  72] , INIT_7A[ 95 :  64]};
    RAM[ 979] <= {INITP_0F[ 79 :  76] , INIT_7A[127 :  96]};
    RAM[ 980] <= {INITP_0F[ 83 :  80] , INIT_7A[159 : 128]};
    RAM[ 981] <= {INITP_0F[ 87 :  84] , INIT_7A[191 : 160]};
    RAM[ 982] <= {INITP_0F[ 91 :  88] , INIT_7A[223 : 192]};
    RAM[ 983] <= {INITP_0F[ 95 :  92] , INIT_7A[255 : 224]};
    RAM[ 984] <= {INITP_0F[ 99 :  96] , INIT_7B[ 31 :   0]};
    RAM[ 985] <= {INITP_0F[103 : 100] , INIT_7B[ 63 :  32]};
    RAM[ 986] <= {INITP_0F[107 : 104] , INIT_7B[ 95 :  64]};
    RAM[ 987] <= {INITP_0F[111 : 108] , INIT_7B[127 :  96]};
    RAM[ 988] <= {INITP_0F[115 : 112] , INIT_7B[159 : 128]};
    RAM[ 989] <= {INITP_0F[119 : 116] , INIT_7B[191 : 160]};
    RAM[ 990] <= {INITP_0F[123 : 120] , INIT_7B[223 : 192]};
    RAM[ 991] <= {INITP_0F[127 : 124] , INIT_7B[255 : 224]};
    RAM[ 992] <= {INITP_0F[131 : 128] , INIT_7C[ 31 :   0]};
    RAM[ 993] <= {INITP_0F[135 : 132] , INIT_7C[ 63 :  32]};
    RAM[ 994] <= {INITP_0F[139 : 136] , INIT_7C[ 95 :  64]};
    RAM[ 995] <= {INITP_0F[143 : 140] , INIT_7C[127 :  96]};
    RAM[ 996] <= {INITP_0F[147 : 144] , INIT_7C[159 : 128]};
    RAM[ 997] <= {INITP_0F[151 : 148] , INIT_7C[191 : 160]};
    RAM[ 998] <= {INITP_0F[155 : 152] , INIT_7C[223 : 192]};
    RAM[ 999] <= {INITP_0F[159 : 156] , INIT_7C[255 : 224]};
    RAM[1000] <= {INITP_0F[163 : 160] , INIT_7D[ 31 :   0]};
    RAM[1001] <= {INITP_0F[167 : 164] , INIT_7D[ 63 :  32]};
    RAM[1002] <= {INITP_0F[171 : 168] , INIT_7D[ 95 :  64]};
    RAM[1003] <= {INITP_0F[175 : 172] , INIT_7D[127 :  96]};
    RAM[1004] <= {INITP_0F[179 : 176] , INIT_7D[159 : 128]};
    RAM[1005] <= {INITP_0F[183 : 180] , INIT_7D[191 : 160]};
    RAM[1006] <= {INITP_0F[187 : 184] , INIT_7D[223 : 192]};
    RAM[1007] <= {INITP_0F[191 : 188] , INIT_7D[255 : 224]};
    RAM[1008] <= {INITP_0F[195 : 192] , INIT_7E[ 31 :   0]};
    RAM[1009] <= {INITP_0F[199 : 196] , INIT_7E[ 63 :  32]};
    RAM[1010] <= {INITP_0F[203 : 200] , INIT_7E[ 95 :  64]};
    RAM[1011] <= {INITP_0F[207 : 204] , INIT_7E[127 :  96]};
    RAM[1012] <= {INITP_0F[211 : 208] , INIT_7E[159 : 128]};
    RAM[1013] <= {INITP_0F[215 : 212] , INIT_7E[191 : 160]};
    RAM[1014] <= {INITP_0F[219 : 216] , INIT_7E[223 : 192]};
    RAM[1015] <= {INITP_0F[223 : 220] , INIT_7E[255 : 224]};
    RAM[1016] <= {INITP_0F[227 : 224] , INIT_7F[ 31 :   0]};
    RAM[1017] <= {INITP_0F[231 : 228] , INIT_7F[ 63 :  32]};
    RAM[1018] <= {INITP_0F[235 : 232] , INIT_7F[ 95 :  64]};
    RAM[1019] <= {INITP_0F[239 : 236] , INIT_7F[127 :  96]};
    RAM[1020] <= {INITP_0F[243 : 240] , INIT_7F[159 : 128]};
    RAM[1021] <= {INITP_0F[247 : 244] , INIT_7F[191 : 160]};
    RAM[1022] <= {INITP_0F[251 : 248] , INIT_7F[223 : 192]};
    RAM[1023] <= {INITP_0F[255 : 252] , INIT_7F[255 : 224]};
  end

  always @(posedge CLK)
  begin
    begin
      if (EN == 1'b1 && WEA == 1'b1) begin
        RAM[ADDRA] = {DIPA , DIA};
      end
    end
  end

  always @(posedge CLK)
  begin
    begin
      if (EN == 1'b1) begin
        RDATAA = RAM[ADDRA];
      end
    end
  end

  always @(posedge CLK)
  begin
    begin
      if (EN == 1'b1) begin
        RDATAB = RAM[ADDRB];
      end
    end
  end

  assign DOA = RDATAA[31:0];
  assign DOPA = RDATAA[35:32];
  assign DOB = RDATAB[31:0];
  assign DOPB = RDATAB[35:32];

endmodule
