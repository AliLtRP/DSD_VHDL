// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
OTvT1M2KiQrIfiz/0uwMwCls5pLjFu8UiAbeUpCbOVjIb6fkCil/e0LPLUnnGZfhq64o57GdO0c1
LzqmgHCFJL2UtxBbczKQs7OQkIW9vzsxme1fkMBuFkzo1ZKAR86vvX2QlDZBYf4dLf+CwtkPKXO0
UmJ1IlBi9nwt4GM63+IEqv35R50q+dcd85m48va4rTVJ07ibhiHNHuR+z/uVmzTfE1AAvX9Ycv+/
tVJNK97O3dwob1sLF2dKYp1liBmEYpCshvvnfF3npZbDh1rouzizxHwryy+1ALpgMgGuekdKJv3+
FW4B79AoDbpsxccnOjBOrcNSk5NraelCsu0M/w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
MUf0ghqapq0+tDA/5JvlUsRTc+6Q+SfsCCVlq1rtVTbsK5MQmGducVMhWlpa/beh8sx0O0Bk3CH7
vB2x8yLsdQL4g0pruy0sI7RHXndW13aQsI64X/6voSf5BJlOAut9g48hR6f8KQwMHsCUUyEa8Qs3
mFgLuoqBQhQGdEbNUCcPaAegZYjhkxogYF/8/Cu3A2xerIkiyf5YtpQB/9GF1HRjmBaUml+2YnAq
cGmCBejI2ncLs5adV2Lw+gTAFFDnzqzkVdZJVG3RmTephq81JEFaUukLz6AEDKXgxcPZnYJ2KHK3
xZmpUiASv0pndXep2bSHWskFWrDHDXxM4Ja39U1TtVk5lZN0KKoTuoHbqq5VYHZY2b3IcKvtLAtY
f1C+FZPnBPU+CC4SqywbMWXNa9tLIopUrucQoM/SmyY+GbK59FlyT3fu35irFzSgcG64xDHzyXMx
rTw5ZqAb/6ZxyL/C+b6PE4XknSZUbTBqnzl5ayte3acOqcN/cA5UUTvp/cnqJN2d+Thnyyh3vYnJ
91l4Yiq3JaXr/gGBpRqY2WHDN3o0KhqtnbpIyGKxEM/tsL6pg3QRlomD1CSFNN/LDCbMyUG/WPqk
Xm0h2iqBaOGi4ZzBAaklGS3n2v6RRvkDFDns4pwhFAA0ENXdSGLmN3U9ivJl7a/qtJIqQoOmXs+b
NG6TqmpZaTWhIx12d/mOO+77KTiEJFw3DnFrraKnAqyve+umQaNWd8gpJIhPP++wa2t2McVg1Uu9
mr25EbVZRY7HhrKGI4dor6Ew7adkpdMumtoRvlFCP7UXc47OMjdz9HREgOKnr2uQPPkTWBm5tb4g
dd2TawPLJdwxRm8GwcKqNhq+rbgV2pSFiRfqlQwuecn2sXcfH9nLy+ipo1DfjliFTSMxhApEN26b
4EyZ5TNmxv2iQc6qzqHlfkjl6wdZjg+Dvi72nfeqE2Ncau48NhKrK0P910AXZARbL+FpcVxa6GEf
jNPx7+HOEVfuvhke+EmInhyLqb2ttn/1mM9QdQgSzxT/ZYleGj+VVG1GAvSZ+bZhU9McnYdUxhHd
McU4eW4PwAfUl9NY3vFwC8zV98e8V3gaOlJOtJaQZPuPEpeMHZup/ZLZpRZmr+TQfP7tE5YcenP+
QojC6xn3O2pfU2qpkz+TK3zTL2IvJDbmW5MGK8X4B0iptYmDC/FV1gZg/SBltxEN6J3OYSGmrWsY
yiIcYCqinepovcYBBFnY6t/4MVkvSC3R5oeO8KSpe4Bpbde0IPYhOjoVYkpXJ7kYsroU4U3Z64NO
4zbhe03ZFF8hKu4H9H1272ISyKoMLhq3IYC51E8+KtmFESo4TIZkJWqhtglRzZju5qIUCHZFDiCf
dFsez1KpjhyjaJCEwT9lw7sWMkZWTvp6KlCVNAaUqn7qCe38TeFNDhvnK7hQV/ww7DMWkGf3quV/
pIyr/pqC2S6mUvowKNQ1b9Pn65bxn5PFMUwPS2Wl1RmqiJnU5rpKAbJQ7awsSVfwyaaucDEiYqTg
hihdbNJlk/i7j8ii+HXXq0lQv8WpZ/08k5qzIG/XgENbOxE/98vGNvRJAx+ngX5DQzCxlDQ28Lvf
O82avud+WHzAwnVAjpL0DZMS3M46rQq020jJocttXMQhpNgcN3Qk5okJmp2kQnq4P8VAHE212dEs
6hXHNIqei1c8/UOlpCK4o0EBU66++LJzOqVywlE/fhSrkTlbsDjrN20G059A5sLOAUXHI8HzE0bn
nMNxr15+nfb/nX7l2ic/+vX/jSFXNk2YvqK9roarv7SHkFVqXYUa0cinVooYrTeIzB3jpEjmTNIj
oPsdtAvFXIQmgIV/LnV8CUqPHFKc2C3s0SEYrcyCqzZfrpM6Nt18hoAbm6ioAi+vbHS9WEzM+rFq
OYLfhQT4+LaIlMcnbrjXWQToqNKbSBWbC60BKrcg3cgS8l3t6LuFHdiQlJ8OmlCAvUC0HXRK2QT+
Ryp/hJ9iD/tMzM95hiN0J7rx5yQ/QKF//NwiiEyfF9Nsm4RN8+Ucw86cco79Qrx1PWWBSrx4PNSi
yauIKDLAvolRaGnf+izdTo3iduILjbkjPxK8bn5dbhWu1Z+JVSZ3bhTXxXEBjS/jKkdPFwEec8wH
BjAmkgIDGtpWRitfwz2SpjkHjap4FoZ378D1GQ89EnW5dz3B+HmDFUiX3AWTdET4G99DlChPP+/C
MrTf8LM1UCu3+zpQ5r5zzyLg9ko6MdW7KycQsBHltSqi8qPEAKk/Zg1/NYEGA4JRIM8wSNFnYZHS
b7AGm1IJZ49GdmlaoY6DGcDxnib0vdEqI7z3/JqqE3740SpS8KmRaH5gl7XHI0CDUfLAlBFIsQI3
5zIyys7s9ELVKVSHMK7SI6INbm14qRn3rkQA37JA+QeX2AYu55pdkjpBGdqfeyCsKYHkdBP5dY7d
obQNybbnvl3WgvfmgXq7HcXiDo/jHnA44YlpizCccuz2kl8bxQCPkwhfOgyKjmzzSK5/QKKp4b4x
9iqgtArXbKr2xA5WfLzq4LqHWZ08I/mA5PTRbERxm39WHhW+5Y0fzhZnZimFm1T4pRBsZTNHOmo/
jH0QcNW+PPWzbjYqCAtPCduAVIoHiZEpGdK1RS2g1TnjGvvZ4lJvmWUfg1ysnc0KOJ3Yh80jZF/X
MnvP2xikbDcJTN/R048TOxcGifZ3Y427Zw1i9DOqanIZD1PqQNRORCeKILiV3eFyyT/+BtA4TKs2
K82iFU1Z3Csxe52p/pUb9oTGgbbK4qw1N3rIDMZuCfgsAmTYqSFevy3QxbkwSLFGIyiH1XkAjL6E
TFDYMUC3movCklU07DVnypomDd3pQIf3d89c5jvcJ/QkzK+7WEVpoX+fwcr+EPDyiGjzQPKCOPaI
zVqnL8YlrWZkTpAqssTgg7TXEiT6qIbQdtnA7z6SL8BW7UPHsexK+5mw6HLz+/igWsL5C2++0ffd
83vkKGTvzxkPeDD6xcQp92et53ogyUtVq6HtmCLd3TotIEzqnxwnyU52zc/GbcquIvVSccwbQLEH
/u0AqXIOra5bpb4aCNrRzrk6iA+LGbOZREyr9f7h1M3g/PVSKTd0PC5r0vGZ6zqCD7mdvP/DERlg
ylt2FWG6fKWzWi3Q37b7URzU2QcKsr1W6iLev/mBZOg00XhFG4r4ePgvmqFgx0gXOh8+hQGQiRs6
Lo4IwJS4QPLaRYopvjx76V2fRhw0f7IyhHF3NM+BWV0fK+VaUipZPULM2/B23n8f/maNofATMn2P
9GtAifjDfceFM7fasipPOkV0xUbPCm7rKz287CPkxryWiFq6xKZjhcCc78H4X7LPe2R9wS+OuT59
Fpk+MioaEdOBIHXN/UdAXKGkYwVa96X0C/4OAEcXcT8p4KqoIinw/rDPCoRb5Vbjx3ipI0a2LliY
lWpt2BTBZ7L4lfsW22vf8ZPnOOkDXZUAsAZdpD27OVeNHwAnjjILlyPTVmrsLG20LZ3twWanNqph
8iQmP8ji4ypj2NwTcQwGXvlYqwLW5I7Rd3R4mmoKbyocRwdvCHkgM/3sFtn6XrQnLG+KzhgLw3qG
LTnuFwDdkfJEmS4L5F05g0+P3i+8erFFryfPsYXe9uO6Ql6TAB1RtG0eIF2jP615RZbrRbAM9Eim
BjLKn9YltjqwF+vdMVxlIbbMej7r4Q9kQz4hAtb/JuYAB7cf08UhyBaGei30HQTxxO7aJliPSKwH
66aI94vnbvAHGCxY6tIid72ZJg+2TA+CKr/sstMfJ+TucAbdhQ0Kquq2l2R3txLUJwKi53hmzlBB
iaGZ0WsiBnBXacIo9aLhGZZp1inlmdwY6OSP3S8HfQPeCUhgk8/2GNdgHCtmeOBJgjHhGH//XWDs
UUry1yROoKeIJ7x+L+K5mLhZdSAVVAyA92TkH814c869emLkdz23nihX54K5sa1i+7p2lBHXtJ5u
fOotMu+GhyHh3LHZKkYcgrJtNX3+X/1VbvrispDzquUeX0InXgJO8OmEsVC0RL2C7F3dG7r8HISC
yERUIAyfFMyfos8CvgCTbcdAzGmCS19GbgAyH470ErxriTQsjZ+aGUyIZKNJV4rUvrh8AFUMvRDp
OEmaaok4FhOf9WLv1Bh74h3fGViaB9898/u6LiKJ0hfCDy1qx4xlvCe1ucUTBrRP9Na6kLfIDIME
QV5jmzGAZO3D8w61DDLBPHHdsGXCh/hvqPRUtUJV3SJK9rUbSSHNlqJd5yz68eLedLIvYN8nZ6xE
IQ5NzMk6+NiMdCCJsNOE64eC2N2nJhCI3BDp8rIzyCiDW3sJ7nPT8TspKM5Uzvul5zp4O5egkanE
A2LHGH6cieOS3wfG7lRyPDuCSrzicDwo0sSnyN1N1+vA8QcnVPXZWtsOLCWXJB/Icv5hapQLXOzp
4fZZhkBU2ti1xsllyLFUHkN8c8fSN7QcSRhwzTrtAHljYe+7mCj9PaqbJfGuG3hZz2Yf9az8jOAc
BECA73ZgQrZYbu++ArZMJec2JTBfVjdZUeXNUv+jIYqswULPcnFHTpIi1UYbPm5fqm6DJOdrwuZs
koUDhPto5uFJX+m2EkZqweq0lC2/HvGrCHPjBa/wXpYXaNGRj9hnKCgdbk5hwJt6ImyVC+5tRuwv
wbb87VcXPKliBncjarVj8tNa0X2jTjfQ8FZiDEhCzaRp35b6lwegGHPbGsvFf8A1QUIOgEK8bgUw
j5FUPNYk645i8MH9u3CUp9FHWJLi228yqaW+97Mx2tHvQnmEz1AJbx0mEg+/WN8/fs7ORDPkyt4T
qdXGc7HvwCqnnJgW7WnDu7nQDg+gi4GOIwXb+aX0blaM+V1ZF3yBN5XREDIskk15sgltQKNytaLR
o+yE9sGdxw6vqObUAGikH6q6GUloa/fz0AY3y33w3zeaDTj2q5Fkkrlqh8W1EV676wPZ6WZgWDSv
SV/32dqxx9CCLRvE0SuoUe+XYTTXEvmIUxmEOMI96W2YTQyMVJCdbu9MHFk+BiC0qkHonVpCKVkv
Ci5t/Epz3mmSIz+8yA3JuvtcWH7POworz2bg6yVcHRN9syIABfzK+Emd/npYYRq6WIPjel3rakdC
cgJw1htYMdnIv0XFiQ7lKvI/ZBuU2P974cSVQD4BDR2j+gNV3ZdPcJPgGSvNQGiNZrC8qNnhJ4qx
6yqoOtYk6L6hnaLxthCPgI2kxvYxlrH03SA5dqcuv4fOxO3jJU12qiwmKO22BcWFEKOYaKQotu0V
3M0RSzUDaBbUyOI3Kw8QfoIcAdE/zK2ZUULdLtNFDZ25uutOXfBC7tE+fr6YXlNTzEYLbT3XAP2l
RK9lWbSDBlHK6+8scfDeQ6dewrIVofkHVIw0A64InJD2AJOmpzTBaKPKc8vrADR17mrmKDPW38hF
ZvlAv2Fwne7au5QZCZMVXpJKnMZCuAqNU0+iWMhGOrg3Q2HogzZRqJ0OvvR1W7kC0MRuqYBRXohb
K+NnUCWm5/bGtHLv83pcHRKx40PNUGDT2NMn2LYMy7warKtjJjO/eRLkVEkm8UChVaRpZk1dPO12
v6udqBrLBuuzB9zMlAyG6bWmxqJ6ff4OIlqCGVVyln34VH7Zi4DysXxCmyV7z74+tPThdt75UMoS
+GrG7sd7nC2MUxMphjtKmbom4Q/2YAZ9jaGSU9uuuLKAYln/MBx/XBQACVAB5sbaOsm7MgVRoZfE
xXBkywt4+PnP2NEwwfeAoY41Q4mB4BaqvdK/QGwqR6wBeAW56huZseJKaY7gOi9oaGyEdqQn0bnb
JDFg2hjFSd4VVGgBJGQOPv+mSfsO3m7Z0/0n6oLtv4g9dgd3WN69GB62KU0RGbQp+RScMI3n1dV0
3stO0QeeagZXkrB3wvuGIoyBvFoWS5suGBDzXp4ETTF6LfELbf9O7xcAkE4CzPbBVoxg27FOGHQ0
Dsru5IxLJJ6HdPMpuMXWJ3p/YJK2qJLvUgrovL6tZLO6b6G4Agoh2c7uuewo1AnNSjkUnCPxVrGZ
M23X40Z9gnPdH3gzAw90aeWXHr0jIx0Fu7/V2SdS34QVsVOrtukP79RQQ3+yhHA7NceF5Phh1XfO
hoFYpuxm0Y7I/VRmzdLaZV717njbGIaGRoL4+9z8yPMbHqdpJ+u+WqfuJHlBZw87+YFEI9iZ3cuH
NCHCbe1yk/NucNvI1C6MFr/ON75oSjY6l0BxaZpnh2DBVtWAim6SJVnL//QVlqvO4++SHfdFxvLl
3R66or9SIDkU4B8N7gu7GVvMLg76SkoeztWYqMXaowI1xISa/iWELR1L3Ubf1YIIsi90SxxJbTjm
v4uJFK/wUrIQxp6/1pdCTi0dUM2/8gmC06jtqiFd49Bt8HJtiAToo/tc3qB8rS9fP78KIU2TLuGr
HOHqQAFDQevoFjr7cPxl0e1eBSS+06Lno/++E/mHoOigW6iJP2pTkuDOcaWwKtEtYmvYa34BvmOT
A/X/jz+Py6zUss3hMG8lOUh684qBp6ov7dJLf70fSnVxlIWMTpWTh0x2RobqQhNoww1VIbsVm7hD
dZE2zmj2c7bn5mLPZIQuQZGZTqQxx25ODqwZGi2AskWm0oORXP1pPwyShN9AfT0TVKDWjXWgzAc1
DjmZUDK54oykJGdiXJEMy2hgsLO/efwJa2w/1a5Vsv6X2t5znSGXRdezwGQAW7dejZ/k2XkZUa0X
za6ZXNqKeVOWTj9Xjha2guVs/7GNqmIJLN8RwYwffEGeV5Tr3j8Ym/YT0ezdA6cxUa9DPZ606NwR
bCx7umr8SP82vsUqxop0AmVziubenLPnZghmE9jGHeRJoUoh9oLYlAASqDvpVvCl4cdRQwnPOX8a
8Ecfn6Q1ICs9qZeFlZODp36ZIwmZ5RXEFg6k3LP2cAvah1LhwquxlBpQ5s3i4zW7iMQwd5BXexy6
FmDF7rj1KYf+YqNlDXZEVF8XwURUS12Kpl8gA0Ta1zrG5hi084WU1Aokq/kzaDwUJxAGTXwufwLL
NWaeWpxBnHkC+chGuk7qx22EsWhyBJHD6Q6yF1NF98QkuVV4nj321vos+9A6DK5AZlB+xOiMKSQ2
uDcIHi3TnTGO4Hc921Pnc5WhYhLdI61m7xbwt0ZLZ6hkvtTetscKpJC6FoAjpcJjNNX3UPXwr6FS
WKQ+aQNQUeD3WwgrUss9FKxxYWN9DzSdZ9sFGtQVJYFnXZpFUTa/EiXC+oUO1K4Jmm9M8IZ3ZSqG
TLB3vSbQDJ+BVoq4pvNKK0tGdTa5Onr4amqjcgtws0LljWQ9DiB2+q+dGfyDiQIYf5KPV44wXcHv
AiMe7gaw28cksd8QM+VRJu2cBwRuv16R5HOJc8HXK4GDQOkCQlZninf51FQETQppaX2SWqMnCeQD
snv7WaLtDZeZGATr6S24CzVeiZdftZzoelqgBuHLj05gwGqeGif+8vgxcka+w94kW3tmTOY+vbEJ
47v2ZDyzzdpbKqH7ybA+RnhmGqBi8C2qSf0iU2D629OZ2EpCS6sj3Uu53jsaPEDuFJL/RnE8Pz59
kE4rS6uHY5w+Ss/fkysOlGH6VOHbhHoL52AnCwq2iujZXKIrqWYxn+9+1iMQwdV1jJYADQTyPLSE
6ERpPB068Ujf2ZojWrPFKsKi3HFpg7wtaenwGKcKK+ayoC9mSIrOyAte2VtOl/sXEuGQsQB0rI0Q
HpsGeuBLHX/KY0v6QMaLPf7UKK+oZdxY+o7yugY9QNwdjXDKigrWrZ8DqFPaGhyIyyTvGiTZRwus
3dwVxfwPqpbqsw9QIuw7rs0/6skUpammNfitzgmXR3Db6Tra7Xp6i33kOV+tmPt1tytWvlhEYae5
Cmw+b89gUvRz/h+4D6GxtYQexBk3XNgwtDN+Kk8/xn6KTrCx1YvzDgh/zg5d7XVEMfN8sdqG9Use
OjD929Rti5ZN2Ovw6ZUT4LggoArS69CLZtfo3OxgUYMzNLi9EKS5ryYvxiF4XktJpeqi2B4xHMKn
VVgBmFP4ndEWY9chOuwjdiawkmTnoNFLu/k9M0QoCyyqfMGIlsJbQFblKOE6E6gDzQSs7IB6NCXa
jbhBdhQ0uOknztjbWGeNHZyzfAcKs4BnoyurRoooHH6bonuNlHsq4V5bWawINsxALK4AqjIdjbZP
RukH18fMPqRjgHsJPWDiKWoJJLJIvWUc37Gecz9BtWgJvspUFg1SK7SLZusBJ8gosiSQAtkcdppe
sEO2dWTdS1qUJMTvxZrMFoCA8jFbQPtql/jnrdn93TdmFspI/pJboHQdgS5YNDspSN8C6Ghg0Vva
htDBXlvoHH6CBeqI595GObg/gt2X8hbr72Yb2CxOkjqfPhIMqVmTGq98T3Ng0WKkTOJwd0nrcG0A
xC4BtPPmI2RIT+dNw8fz8M+MMkclTuQIAYEMCqwbVjUEIjZuRQIbFGnC00Pa8ILPfWt7CTTCnpEa
OzAz3UlH/xpPjDFLnjXGjOS6vrAQ8IDkJBGHFrSCoTqEWlofAhm05ChKzDGANhFcAQqeXRV5cPHh
nSAlFdA/saky3sRU1igHe2IjzshIYuJxLMPXu+pFljl3nV9PMpnw9bvm5e1KilB52T6xEpcSdt5Z
bKFrXnoQuYlcub/RkZCdUWK8+taQeUgd1L2g1c3I7XKXZbOMtoghMC7HABngzGojcWcR/FBPKD/c
ZeCilOmj4uA05C30YHe3LkM8j7v0fhkO+8Qx4IDGhH70iPhbF2y8mcPqpuHRvsL1A+jPiXz5ORqt
/3vChz3stkfZMBE543e933kG8eegrlmplq2NIo/nkG17MWQP7L4FBotiqDgs84goAVC9lpfQxbEW
dBJqadT8jlsMBXCe7U1ECyXjeB+zsx06YANjS+9eVVDcMXyivCkXDfkuiJYqbiP0m5KqGev4H7ta
3RLlaC8mZRFFdRE9ZsiF5KjQRfZyp9ZTNELpQ+fFUpmgGxCVE7rRxQ0X1ovyUbrLbmWatzB3nO1y
1lT4HFPoMveM5agsgHkKb1q+s3uaD2Cx2h+dNJ+ytsTHY2WSB4Gotc/0rn18Nzk35i+wkPQEYQEl
CdZ3PtZcwkrX4kw0nlq7azRWgBV7L2JzLWAH5UuydBugkZ6DgAsVx5HqMj3+XzeKbiHifxdljusk
ZwsHhUg3poatrKKksTBjdngRKmbB5I535JMmXKgDHAs20fj/Kg3kxe1Y/K7IQ+nOTV0CIrh9VGrn
4pFxTvm3nwuOaTR2TtVjTfilPbhG8BIdQC2/g6UheoLnH6W6YslG9c4ztqZYuaMEO5mm7QRAxO5F
MqXh3ebVgBDC0YTYPcEDCuCkJrFy8WD8CfOxA2utUwAU9GuUQp+oEO9dRPO2kubUlub85hL4JGUV
wJZsKIPjris/iPbtdHiQsIkgnQjNMkarHsZ7JIZBmovVBM3S+N5Bwd0AkVJpyGJ0DgrE4MLdawDh
V8d8+pBtyslnPkddSfcONaHCOa9FdAaKDMmbC59n8Mcg8U/LsQiOML/gSycivbI1VwssFT+BWzj6
G4etQGM2qXipZ8PPhVAItCemoSXiImRhabkjwjh16mKs0F8ClUzfShiY2isMXDpova4B1NiGszGp
hdU4zXsiD26RZc10uD8we1uYPuz6+EB/HjdT1SLiP20T3DAGmStmBcKI0K9Qw8k3pghcNYU3jI7b
GoCGiejVOyHp/VabT69TU3BJ6GIynUgegiXikcvWRJinlTR9ofV1/Z6h8ujDYOg3TmM6lGDyq5rd
iPKnASPVHs2n9/p/G+EXyARbynJeGbz3jWHtp5bO7LsfoGoqSzhztkNGe7aNQMIf+2kFT4vERqRv
KXz6Gz63Y8rA5WVkPlUNU5Pv+lbdP9ktbaN067jaBadd3qa1AhbrVRiK96Kx463bRgfy0ra0XP7I
KseiZ3FY5U97zfz3ca5JarbadLRAQdB8r1whIpRrH7ab4VaJEezosWVlJEHjSUzYFu9Q+C1x9wGT
wTnwd6vpvH+R7swMb5dnmWrzfeDGG5xaVFlragMA5tjdtLeUF+r/bcjImflNCsrj8bcIDKJugmVG
KI2Es7yr18SF6QdTDEUxnc6vOF0mGGSD3FpjFtQT5AY6DbAvyyg9GFyuZRGulWZTV0PcKhtZGw6Z
BXTmLCrcD8aL3gItn6cbkjmPXLa23Bo9+Aboak3UsVLVB9KVSl5c4kKfGqKiOWkHxC1TaoogXcXr
F+1uIVRM6K9D0ObSRDwmt0inbhi378CFnSstaOT5BuxJIXZmlNPhauqaH3KBw9M2UeLURDloyVLm
BjFEZfz3opAmxvKylqC/3CQm4Ld12PEVHSTFztQUm94HvHKs9ujtWExrDO1imRvOEZYokFgcI1AC
tIOsCgYbRABTPfvsxvxk/lixzX4tXJyN5V+ZERIJBio7fW7iAM9wjRFYCDuyRuTpYxF/P07Ajyjb
U3i/qn3fHW79LWYWA0sqCOx9u6mZBEKi9XahhPb1RJMf8WY++FPiO+/c7STUU7tLiybXF2FR5A99
04FT55epl3R6QHDdmy/wUep82gvV31SSnOy6WmRNjgAWaFmaNGXm8/rxwTX1SZObz5+9e209BvZE
FXOImI6+cKUu1SG9S+s5VH3UJnoBWLX/kjihElZ57loV0fcMavMc7UJfBdQukAJPGXEXcZlTJFha
WeXKuo8mQGdhjbHxx2hr42bqfn+eW+5lk9pI8N1R2Z7/OSFXl4wgK8PtWriNoukn2oDwr3WbTuUR
1JGSd81a0vp47DdOGqYeP/pS7YPtvDGKG4JtNw5342Vge4NTlyOtLwUSyizhBuOnrKBqnxaeSAzx
D0Hl3HRLSPHmMzRh1WGvRNnSnQGk44WCxgkRA84TBOYUnlKkUPbGhVjcB4sRBsFF+qGiCuggnA8l
GWH3aDTvz30ZF3Xp8LgKM/1KdSnQ1ZRtgPEwNbcNZF8rNwM0ePMW6wjTuJKGkD7UBVWJzQTJmpDc
o8bNnBMXSVf+iusfhQuIPbz4Jhu5EcvCG3xZsyFqk0IKlODhTFZFmpapVmwuGDvC3bE4ehRhLxBN
6s3X8A0PrEKJYVnj7Xl2Mo4n8tzOomK+Mqw50Kbgaq8BzVXn+FGSPAyVxz1ovlfBI7MSuSwkNbbd
4sIyt8/obVMbH7MCAuSnI5DT97QkDjpi5qcgoYnU0EIOG4fU5qaJLhHstETiO+GxBK9EbbLL58h8
FPpcfgtHfJZvIoZTaV76R28GfIIE8jiYKAghw2Io1SColV0Bddzsum764Mvmk4LWjPa7hrL5385c
jOIpzDgveTpD/2as6uVpzyBAPZAkYzCEteOAekDHeL/K+u44QsFGPk67qkcTGw5VBG3GzepsMTlO
8wQCrck4rDy+cbEQxwFHeN+vP2CbIlXHkcCjpWe1UMdwRw7suQYPZSNwti2GB3ysr6Ros9dUfxGr
e/lyDDF608wmJalR+XtsfMJtM8ltkLBojrJ320Fm3spq8hNJKfgbKrEzuCu3V0cVDj5aQLaBd5w2
hkcFBl8k3WZ2pB49+apF1nerom0wUWJm1R5ss+bmyrqXE0UwUuzciKK9+HAaoOxQ/lDh2b5K/cOt
317rizSqqdSHZO2oJ96MwP4hHRBoLGVuvxLgJvMNre3Gs1q6BGEGqs5lNwhJ46MqwCUnFToxBZRg
0aUgbdttmlvXNeppzFxzGUznJN25fv37bXyvBcVPP7Ufh75Qfea5Wv0hlvBhhqQiGqchQV4gB0EQ
S6J3EJrmC/AIePb5FtvrEP9KZKhFGiGg7eqkd+nCWXN6dEoYUWWhiBGSUHc7J4MR+wn7OUNhuYws
CzpjwiGCfsTpvDFPnoUQ7MNsrPI0FNCzYvsXo5QCZjJupai82pDwEFB7+obpMTSnF/6Dk8N3dGnK
bNm9HCvdAIP1nwpZ+we8RCWTRcuQwgjoaYfWsIjMbHyEVy+dnDupUEWryNWaFdzpk3ALRmp16Yvt
UjGQRGwcRrdxuwY7svY5WwprvD/uHiOqzeQ0JFLMDFrs+ENvyoK9RRCEgP01KEOWVH2lg1FH+WOM
XrzxBD8ATwyJpI1zj0MYE5IwcxY7unXnJejyOLufheWyC+vD133B7JwFLPrAS4dMPCK+crmv6yk0
RJFnng3wYAc4VcRr2YdsCFn4t2JkBjgrFfIaYtDF2+u4rMeNEWIN54h2aCWr20tX8XgU4rQh+nVc
Bx7z8LdpHo6UCDT+ys9KVfC5Jd8dY+IxPPY8JsQ4Vn/gt7PoRvGr2lBugHo8rCCveh4mR2pMdm4F
+wjR9UTK6yW98o0OoaXNRYJ+F3dSUBBqRK26mh1lciJDinGVJzXqV9Zk20zDe/Su8NFsbsUsZaij
7X8sylSAqeOX31Phq9Bcjs4HrRcC3bWDldoXdOvk3kA60AcKZlG8wyicH/2Q2RFEdole6I0UChPb
KpLJJd4qBjjq+gmgs6+XVpyiNRxJpoyVWntkGJYlLwpXzMEwykPYynr96QvYeBAvXS4rhS5cYwkQ
u0o1U0jLJ5eomY3vSVOnG3lsQ5izk2Nlget7zbrjvxXKxF8wogGEMAYQxONyfFp0rJ4In6B8hGPb
BCcqLfv08UKlZDtf5zSoBfiR4jm1Lqd2CHLXY9AuWzrTMlk5R/ZEo+5yLb+Gyi3b6xDZcQrq7c/2
Vd0FdCMiOPdFZUyrpB5tRfSJYYyuPfNrKwk6xYPFwbC5xppBUoHxWc2rrRlcmNhI8V2vmSqpCRdU
LnnIjGmTpnCbM92mYQwdmM/vJft7q4ILrduUNLbwlaSs2fJMPi6zYvDmZvYKh/RoJoJKdHT0IW9w
0A5RFLmMzvCdddhibs4dFZfQZRmI9+d3QhG+qtK2uIhzk1w/77XhTjFOSHs89TpYrTVQa2a+yKq3
hExFv3w+FXW1u6e1NUibTB9c43sG3D7HXdfoxvPCX0h7wMjwQ+Qa0Rj/nRVSRLBPBP5S1FCl0Zh4
U5ISfzm4FauKG8vNMMM9gXJ3pPjAqEgMQk9rhSJ6PXDM4AnpwtenjgGMptbDq76IBXYQZB/I8jtt
726WSCrTl9yZG5x8jQq5B6FouBQLHcmB8XPF8Qegjj2Ey+rdEbpVG6RoWH+xqTnq3Ifz7D5Gf6Cc
WaEXoNe9fZrLNun2u6kd0BHRBdJ2FSdOZZakSBzvXOAB67RpaMbFI9JnNlJNY0ciiktAAATBL+To
r0CboVXM6UonJO0H4GLLaqQ8QEE2l5nN5KYsWkDjw2Nxva10wzyqs19FxQ0Ghr2Jx0PXHXHESmJe
oJXJULBjIw+/r2aM7lDtnyi8AUSUV8bmlbmiYLRAbAMGkHEi7NSNs4z+obp11i7xR1tPeEgRWDSD
ZHWYujqGsbIKMuDs/j34XmyTJ1gWVNNVtZnSFfMldlq/VztiQCm5940d7ajJ9UWgZXKB1jL1QXV7
+Rm7cy0W5/Rv3zbCdbYYA7gLL0Q8r4SJc/VqFBNWCJb9P5nlo8xt0A1vZu0zHVy4q42TfEP0x0Hg
XiEZeLuoQ5yEQxARxEWN32i7drg46326+dpbw3mp7z7dCBPii8YV6RVWAu44m5hBpI+SAlP5RJSR
0O7ztNh+6pk6vQ4/sbeYiGV3Mh2RbW0zvp5cJ11oGeNNjt1xN84UQU1gVuVgiePsY4VAFi3G+4lb
MCFbGwuFT32BGyfD2l+CIfxeT1dh9ljA5ewIKFkA010gtmbT9vLGFJ916R2/4xEnAY1gnrC/x91f
tdUPoqPqql4KpAcUO7NGotwO3Mp3npeCwe+bg7lKYeE8Xd0h9v2F2FrrnN5WZkAh6gSlzE1Ssbsc
JgesS6M3wp1pqs2SG0xsLwFNmviXWyBUTo3XDOA+RltREbZCVVn5+Xz4CLvgAp4Yr4OhT7a3kpy7
leAuSJtMh0peaZ6vLlR53bRvd5sNOioD88tmZWAwqKc4clSe4wOloPRyjBFb++xY/80QT9QUWSBC
9zNSanXw21vFn5VUBp2JQpc70RweIeospt8CE+dFEe1Y5RmCOu7lKbGC/+krgBgWlY7yHdSQCzdB
1whpY8Uvyk3d7hz4JgutNxE37Rev0/sRVbd0A5C/GoAczpKTokEAXiNUWfU4a4JY/ZsehALQ+Uzb
BGDHEDrWgHo4LavqOqBUA0MHATtI67+XShu9FX8VCWb5n/7Nx5UJfZCepMK8v4v+l9q8lcaoWTNe
jBkMvdBSnA4PXqm0t/eYevIkEcyEBhiIuDz74fxI0alezyAXiALeVsJWzq/RRSP7K1KhL/5czcSw
ZEOyCs8e0IYOv4IJ1V2p3xIUTnMXt9AqQb+YEJMW1kJbPhEoEK6IBRcqVIpbj28d2SABgztTJq6J
fid/BDE3g3mQ4/hyYH1jJ/sGGxPRiZ6v8qFh4l71Da0Q6cEbVhWGeSI2wYF/kik1ZxoG1ZwGAUFL
Z3vZBQIUsEWfg+DmHvjZMwQZvTDxZhQyIJcGlnaYqYPLUrWENtMK9K1P0l83OFhbeTCMFS7bKv/p
xTC/BkQsDvZCXLZsSBWtSmfG+WdmK2KP6pF2vRXxqeFXCgEaZDK8hek9a8EWxCLfdiWVC0kyhsld
M3kxlxwkx77LpuWk92XxpPfJQ+OcsLc112733augBEW7T6LURinhha4i8mwthfrJht3qnwBVvCy3
v2Y4/PBvOrJm05spdk7JX4FS1WmV5NyA7lV7VVkMpMC03RzEziSIavx1mU6Jqh3POOF1Zo7oecRl
Sgs3XMR0kmeEb9o6Sk0FpwDfzCVvLMecoZZtw4nFKp46uk6r7+liuPtf0YKMsfm6oVsC6G8omcSb
Ozx3vj42nImS31BBGJwpttq8r5XlTMb0ieDf777uOQ0OjBw2OlmxffOszanfnrvCqheQc2wLlhng
nwwpXvhunaRfjHmTr2Ef1N9Lc6HjLUDdDjrHX/Bfwn9Xj80cz5rQyNUE6Z+ZidPPQJFZztkgbCN8
NKc0sOwYPOnqu5ty/IEfex4dhPzfDuIYNbtGpzVle+uGIWqsmPmBSaclq+ChMP5YBKsGxwdseDwx
i5t18Xx/5stEDK49bmyBuPUr8WUEh9nZho4OhnTG0aOzBHVFC/6q2LEnyqtP+/Su7Xm8CEpcrFFw
+5++aXewCDmMy6u8gXDTTfUnHPZoRKOjYxdmEac4zO1fwY1K8ibkHKQNegYxPaWgVcKsdiC0U37+
cqL7LzJ6IN5zfBto6B/ZlQRqEWCUMc6ikEfFgpC5JcdZzkCl0VFObEmFxv2jvsV7urb7iySJUdeL
9j5VXg+K8ldSGULFQvaq/jx0A9HpPdY3RzOx6kJ92LhmFbRgFYHwOvoDmLg7CojsN5wgFIHc3IHb
urxS6juylA6kZBW347c7nvFCP2AFcsmqrJ4sHC7w8rZXpIrMQnzBKKDEjzNC1vyeJkXVa9kenfVj
e/cgxXQeWB7gp9Kf3kVL7enJr1g0xYFld/KhmLKbLm8G/gYXdAqPmvTgZMT0+7NJfRrSrZSotn+X
FMyU8STsAtD/SxC2S3ooTWEWoov65D5xF8LKx7v5ToYHJ9YeOjW0oLb/eL1rk36j8aIGnZUVBy6/
q2GJoViP05HIh9IpuGd4JNBo235LycRFLx/rEYq1sssfbr2oqPfbG0p9zajk/Y6+yuBBAjEXdYqR
w3MX0/wdSeGKqU+g2+yBtFtiTOp3xRHTDA6IngKZpPdcrTDg3yd0JS43EEu9+KAfwylXB/MprTsz
50Zx45qgevAQp2FYVvj+K0kvfNZoY7BQya3JC+itoingXqk8euIgz4rvjrF4YWkbEGezQwbLZ6Yy
d3yi4sV8FegsDZt3w+q13CicEOXLRsKeJQptDgja1tE8EPmVRuivt3ssonDTjmFG/0JfVNj3S3m4
GqTOEmGg5M54+yTmk4BGAzajTOrNXsxNG65ZVxHBzMhqPkz2fop6/rJVvuj/ATuH3gO5YhJR+PVA
9Dw9er3vzmhVBZ4sps4NBHvmNud+Daz6Od5O9UgzZlwlxfG3uXqu8/ib/6ZxwZ5bYeaAULVgfH8X
QZJsY8TjEZ71F2Dq32F3dR/I++Q21yWQUWxbvJZpm/3ut+kp3OcIOUGCF9C4J/y+Y3hnpkI5MxSs
tuPPnL5j5GPHec1mMyMmUxaCJu/k8holYw20S6IIKCGMObHlTjcxKw0K4zECAc/otR/SxD828k0W
51vLGZDfjMkg9rtWmyu1xdXycMsg3/6mOWR71ytks4TQDRjU7oPHf97GXZsv+GAQ4xJTlR5RMfdV
LXiAsVCIii56tTtW+5i0eaMD004deNnZU4X1o+1cfjx9W3wkK/W2++9fDnEd1kb9hBykOkY11J4P
lJOAD2EI5yUoMjfHqJmSDD65zM37Dixb7Ek=
`pragma protect end_protected
