// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ef7pI5/YkI8q1dRdftWJ3PUXD31ZkC9fo2R7zOTvZ6gucp4G/5Gpf5vR/TQSoQyP
gUXZpholl8v2JG+K+kdlnI0IGXpvVlU2+FvPkKKDhpFm1+cfbYoDtcaraSXzPMgZ
mCRqzijlr6Btg2fGl3wHMjpmgIjin0vb+R/kTW782Xo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28816)
LBbxPa6s7OX1X4xyiWblimMKPPc/IoojRLiOafGf/eh4gyyB1GHUvVk65cgYLd/a
CuvPPjyr/XHpWIYMLDtdCcMIgFUIglnvdvAGAk7FyZF3ZpzU2JbX3wKewLpLjPmd
HNmHy7TrZqaOM82tEIOGCxzRELNok05MzCMN6lx6XcTCj9ew3xGYSNcsNa6gBwlX
+x9GNJ37DpV9bVSzaBr89PWy34qEyl1fdhCTqkDROFjfr+MzVSV4f1SxivBVePR4
EHgptTAYwUoe7hBw7j9ctF6la1TaclDHYK7i86Dk8K8+ewGvs1QwOPaeXnzPhaYj
y3PjH90YXTh4AXIfDeDmoW5lz/6uItHeMLQJR+hbt1uNk2dB5ErrGVEN5xoHxNmQ
8saVb8GPC3uwmrKIXOGyGIDMl0nThJ9ztQJNngCj6Ao0JwXhN1PYDJlwcdyTQp/0
rj6F3uOsHU/VUaWqM6FpfXKYc/91gF8lgHaXG0ZmPyXPyLXZ99fxNbufwB0/WS1K
Np9acopJAu2PjTfqaH23CEZuq0XykaIGn+k9IXhaYVItKV0+8T0Lt7wAAbeYicqe
0zvpCtV2pMjxOd2yArxrLkz7e9+pI1H72PxnuJRhzPps0FaRe/EK79wG6MTvjzP9
SV1kGQhfpDe3reNOtxtRpX/3dVvsy+KLj/lSA5Ud2Brxd2ijXgqwxeibjtOVsj31
Xdy1jXSwQfvGsIlMj5kMucz3hBdudgY8GJpzEL2sbXY64VXGEKuZdzK1je8GdWna
c2u9Xj3AXQfT55Irn5JmguhrseAe1XLLlFefzTK9Sbn57fA9TyzmgMHTCEO8EcGJ
/w7604uMOuXWXY1thg0wAbKzGWCkDMcAxnJh02M01OnD59x8Xk7Da/OCBI/3G9IF
7hSWFbrh0z+r2zJNbZZNmykh7u6p/BeJX73avpDkviz62JdcphrAIQpZfQlrlA5F
Ugyst4BID1klCeB2ER1p1UsrtfZ2jqd/Mqp8V6oR6MA7joqrex3aMrSKuaAb4Yox
/C73KXJ0Z3lU/YSR/sYo+vF7R+GcSr9AY0jdKuvAX/W0QeKTJfXkKsscA7A5hUoL
Bf3eooa40YYcTf6/k1ytKdmUDlRR3xTmvfHfuQ2uTVEfWiqHch2yOH+HvaOPvVGL
ECkPh9+aQdRtxt9LwfIc6eSDvmSWZaGBWLr8Noi0u2a+vBxddk1YYZQ95N1bkK9P
V9X5mNFDeHbwlsdwUAT5WjDSb3nsKeq5gBRZRTuQoU/x8V39DUilSKq3bManHUuS
jo2s9f67uITEzrsaTq9MJ2LvUCG4CJcnleRkahkYeFKoUoyBwz5GKZVBxvDsUXBz
royeZuJS8B/ptzLrgXg+OjtkdZ+Nbxcq56+dxdTKwMICTFeT0x+b/mqnRraLA3wI
Z2xpf4HIOM6aJWEFgXJSK/zldQzq0zzI9cv14NCqzJ8bHM5V2AVR0DE82AAYs/dU
yD+LsfCboi8XXVjA2wApDSL+vlAkg1F5U4SVWae04sxhaJcPcXPqBaZ//hQUp3/P
MEuaYGcH51JwcZrf/wOg73WVkjc/WGlXWN6pNhorBhTc2VgTTS+5aOUfMBlWOOS7
YM4BobYkExkmwxWiEREXDqFrO/OK1xFlEiwZa69vyj9c1FyPma+8N6bPumQ5lD4Z
nK9ZDKr8OjsZogw8FROWC2mQK2T63Zd0i+w9hsjMN4CM1kudJ1eXrgPfQE0we56w
I32UomdADE/msc3aQpwacTvLW907N0wG2BdGpIPWl0e1v5If+nNOAc12+S2ZAzzb
4pE71Sf24FHgcuu9rf+4XMwULs+KkkAWawXUcdsq91tW50ZG3dWIrfiS+RgZ8/sp
bEZYCNMusz25OItp9aQnr777G5+xTwVXojLbsVJr5dF6IT5sdtXVdaQEklVGgKDk
l0rfscPTXdbd1ecufYLf2pl81VriwnD7x4uDJIUxHnbzXMK6hJZgaV72As8lVOgk
K2gP7sQZppNi/fmS+DzufM8gZxqsQo/RONijnr6UwDayrKim07ua+yK/RDk6ULvZ
nJXPWHQ0/2bbZ9JosKf+wWPzvGs3aW/pXVWDorw/fN0OuT8kEf3HVHNHHjqBuTjk
8DdjQxXrmclw1BNCepkM/uzqg/8C/BlC4iBdtpA9goNIFOcv+mdS4nRJEmK9k+Y4
+1fPIbrPj45vdCHcveuGoyax20hXdHd4s45/IS1EuFJHOOFuBGeQDnFQOUKDJNrP
gtW56N4o7vFzj1G6qlPtVOdZQ9EPlm9x8M5Kte3b5+hP+QlGKML3Lv85E/m6eWAI
pObt5Ii6Wte4hP0tOvxfgb6lOu4sWnXHkA+DZW5qLfzi1rYuFjyNsOvyfVQ0idwL
mUR+IIeDlmKCoWBuxIVJaaCUgGb2h/XmWy+jJ8jmyEfjqg/Pd6+7vsvidSZjyzav
JZyG91jAObNWTo33z2UpLHeG7jqkprdZysdtRXxxB8aBCwYk1Alry9jruj0IziAF
74LmaEBnyN9SaX3edRQ7239VNmMoXgkXV51VQ8D9qlgNra/d/BJlHv8wMtL4+1rW
X7q0oRlPI28BEs8Ku8H4ikoD95e83UEvDsdFigEsO2yt4bBIzO1jlmUZ1fzXiiI2
OobU1knReTDMmp2DC/550PCAIYe2J+pbrwndmWXEv4IKwApsb7437ENvjyuJBYvw
HcFtzmmcamI9YWHkCFh30W+YHAyvZmpKGZtBtNm5vfo42HyaB6aNLAgZ8Z/JvDOk
uT6g4HGtg5CA/URzdoiV1LPi0cTi1lQKxvbraqfk07Onj74g9yVPUQ1wec4QevLv
WTQbqNk9CzbgEYEMlSjG/zXjW0iEYELwkny1s10B0bJnjw8B9E7vpd2aSUSZ4Lbt
A6Z1wTmgZ3mAf5EcFzIUME9WgNh+9hZSEH7yHhxd/U/6d4Pu1BE5Z58z3ztoHMhb
2Wbvt4/xicHgEzMTa+CGHZtnyc0hgYYaOtUcJUhTOU4+H7H7QTjCXQ/g2I+7OUm1
qfp1xKbpA5SKdNBGbCJvJDRSFSPWUuojEprsQgc2WbqS+o9aE6MwIaW7F6eDOpy6
mLI14l3gBFEWNPImZHAh7mQ6uyzXzy/w8oYP63SHQiOSXBXT2IuKOCW3zI2fzthr
/f++4FX7wPmuXKZVg347tL0jOeG9aOGuBN1yqzYYh/E93qHYPLEzhr/yngXSkTVd
kv2UP1pDS0VLFlQDvtqeSI4AHQi5Sr+Mg56qP/UDsg0gnt76xK5HOTdAVllKHGud
nvVZkuKFU48CuZlK1oADrPCLHMjuMlW1NszV1bzgSJ9sWMZt/TLnpscIIzl76Egg
SvnAD8Vnv5+ajrRUbqswOpK/bc61PA9wBYr82TQ8i5vs5RzP8s6o4QqHs+wegh5m
F18f/H+xb0gmWCf+Cg3GndvzLyw5EbNbtis1GRZFpweQTg59jCPaRRwMoGOR7BGN
q/Jp1v++0c/GPXEBrDk1T1QkVOIVJ43vLCS209AFM9yogO09PVxmd3+8WMBOaNoI
gyDTmufthE0BGA68SiD7j0R9drn8KSPFirs/hLOW+RzmtZggB7HvqO5jeEE4tX71
E9byukuhYf/mCEoP62uxuRiIYf6kotTrVtdsVOglL1hwE6Kp+ETCljfs7jbEO8Yb
JvD5jG4xg54f5nYkiHOUed2bKf1onJVSQwgnG0ARHQwwkjT9mu6MxH00N+uIJVbt
gyz/PpdGcl4XxSKuFgkhoYhe+UmALwqKef2bQkbXcTjWFCovx3KzfMw0Ucs8uTlW
S3Qx31n1OrDrm1+tmSSD4WfBaikdl0eTsJHluH/2crwwSr3h0Yyoqm1EoX7uwrwC
vJon6Vw46Gn83CTHH6B5OVK5ufuiH9L2g6SdigEZazVDDfdG8sLLCE04WByc8D7n
3il2XmnDctshCCsVk+9uZDoO8HYHLpPYh0f9GkR1VAEv5FQflNLTmLDR2xUEx6Vr
BmEEa/oTvavtqD9D4vR79X+wBRboOIb/6e8Jewqe0JNwFTBcoddiaGE5cXoRFHc2
t3qrO7huP/5XB8E1WRGvQCYoA4hwPg7Nt8IjgQEqsoTdgEPlqYcENnZon7XSjtpd
1j4pu+tOwCUcXZhEE/vNoPfeRFtSX7bjU0o3CYxepditQXGyxvwcq0IqZNEy/Vgt
vr6D6GGKR9bzneUiIS6bo/WTzwp0bk4GvoF52b/W7y+fJ2+MC/MyzP+Jw4zVM+XU
MwPDsUW/3w+DLKYpnFq5ZMHNybWfVw+yYMUq183spYoVc3IvnA54grU6RwQRWrC+
JqzTIYKUxOOfvrSCH/X1gOGO319FJhJ1eg3OyiZulRpOMiA+q1A7bOJmi+cRVIai
xh5VXjiiOx4z88Qfgl6cE1zmBWYXMj60niMxRpoENVgMtAOxUNvvCckbUQb7t9X2
XDF1afZCQQMGI75C05LH1Lh9ZWh3WPgwnKFYoHBTjmbfrUQLVLSivem+Q96h5gl3
Lae0069xSXhlPNII1xY5THiBfO3Fz59kXVz8xHBDGHSnPJhrAAsy6uBOO3UqelEj
/XmtFT/ZA97ujFlwkHLjnP6OAm8UQdkfsFWMD3UKqAwBj66K5jSxd+HgwKInjhcZ
aqyXYjGAwBrehrbGiLPM6sbHiWKWDII8zm5W+nBOZ5SWWJyRb+cWjCd8g6rVhPlp
6uIrytCRXEYtceqQ/wejyRfB5JkuHPHmIj3nU0WyVmiAhRW/kpSGcHyYwK8brmbA
ZFLSaq4C3XkrgTY/VYblWYZ/M8mN03P7G7xJ6TnMAZ0S+H4PH544H+bWx47r01Y8
UvgVOicq8R9UEyv+RT8Ivdh3Am4NCouWTn3eMo77mfIvwoOpHuQU0jOA47xqIrPg
XlkU7YMGKdyZl7hFcXfpwQ5Va/pphU1HH5geb2kmam4dwLv3+Nr6jVWZ9bSj9BT1
sDHAQnDRSFTBN1zliGY2sh7s8A/ElYKL4lm65mfrL6YM6vbZnBFQL9c+Gn4zieTh
/3r9x9MvwoMjqRObeHHL2p85e60rkZtuqvFNpmKbe63tRCG7gP4gQPoZMi4p8nJb
D9RhD5Z+MhIdmMllr9yqVgmzDr53J+GJmL6ufyPp2gn7Ovx3ZdW8wY++GSReGoWe
aohvSVNRnJtEm0v6iPi9O2J6Fw50D+GbpBj8M4+KXDID9wIl/Bb05nl4+rAcAONy
ZNKCy4IZ/grbQbDNkqjmZZXP9V4mPMXYKH7Z/52P2q7UN8K5ZdR4sq7okcndwSNC
mEotVUqMym8W4nKlBUFpCMQuRaornPS63oU3uVPZ/YIDOop0tl7RwkSdqFrRPmlr
FtmhbCES5jEYw4cO+gdgATxleEuv94BlvgfxxbLIIHKbqqPKXn6WU/X2UXgMUfXh
/vwUdtUaVzcOkmmYC+6CV5nVSmtL57bHYHiVbbuB8YXs+PtUQxBWIngVWPOKl6AZ
/R19tECA1MqEE5pW5mP9HCWr1Wji1ooxqox54D1F6yTHcZkIPyzSkqy8lAeAfPEq
Re6eFe8a/ImvsU8mqVGNruW2FlmN9xVDrctlo/POfmMAUuxoR1z6bTn7l7f+CwGq
zU5iRn4Z+BSRiqp/9jUBuZAQnSSQZbPJvob8R4xlGo0ljZ04D4nswlVJaeD5I02X
QakD0Xu7eFMBWiVpb/s2YxEhbuGRTyrePZF5DxteOksKb/FPsmqCl9D7TKVe5wbX
0+54bY8o2zal+eBzE+whEN4jTfKoTLQjGyGKEp1n6r7cfMi/Ax9x+Z5Wrq6tKnTr
ewWc4B7MBIx1CQUVQGGkDP9r6PUMI/ztZA1EmZDSH+y0kPhsid4L4tMqa79rdCv9
zRxNHrZTCLHsixNFM8FadCLos+TlMJyrIO1QKnVazTxK7wWqo+zZlUIYboewncK/
XmX2QduuuX10TGqKxw0d2DfMoWVf+ZJwU5nB/6bzr6oW8fmQZEcXGUv5gLCO5LOF
704KpXBHH+xS6DUDFhmuvwL5wf1/jjD7UlX9iRshRCF0kCkss2yOlFMOtSYUwzIc
jH2uol6tOAg49La4Nywfvopk1AeMe9h3z5Cx3OCbK5jOajsgbbvWxqMulBgATOzi
Z+tDhiBxxFjW0kpp1B3Z4c0ocMuBvLMKSWU3zwPyonOaMY3Ku0/yfDPytYFV22aW
hbBM5+g1Ybqzvmj0CRaYVoItOzOTp7/ox5gvLfGfuFk4RvB96/s7VphwdpZnLWUu
12Qyy5uhPVt8F2SsK5nre8sk4p+V3GZv0ST7s0tQVGhaUocGc03WNlYdQLL1rRUc
mIPVunHBtwikGq/xAhFnlKs6EFsRvEv3O7zlPqzrJ9oSpmebMFJLXWOAZtVMCdQ0
7mMfBQ7tYec/NeX2ltBDjNFLqeVg34Sb6FbObdmNKR1TGNZBmd3wYc7pkBupOWCr
ocZlbiH0MiTh2lf0+9x6jhCOsUN2NACGyPL5fvh6hBTbOCiPpnEim5DlWQ1XrZ/H
ED2qsb8BT+27fZKYq5zY8mxGJCoV0h30D8to4Y1H1KJOQ6DjwQEGqmDh7OF/Xd//
XkKKlg80wOf3x0GqcPe8AI2ertuoxx0L+clpKhEzgJD9ZV0mYyzSfS7gQixfouPt
sYe7XwANORnks+DkaMOIPbYFEQGZ2PEy2nu/6Iisj54zvCtjlpffSj4SgliRKkVW
rSUOCG9BqTDg03fZ5mw1k/IzRdmKbPyVVk9wKygLx2soMcmjoST0WoO1QbSvXFet
pvQQNfncajLTKAUJjtAWTZkoZyR/TcgvixsL3txkYRiwRcjduMCfuvf20GqyAdId
7tWBH8HIyDdp+zcv0Im3DPNZvZ8JwEMpDHxMaPE7fruPCnvTULmNAKra0f8UHqUW
2pV+DHsKfAiY0p/0i6CW4K384gFfmx8KxyFqxGCkKzdpVniQxUAZ32Md4U8+Sh0Q
XEu0QLM3JD86sUxZmYHDBFFvRI41ybknq2Rm1zRxCoZiDPoF9IjRFMKLCdG7+sPL
Dzk7ZErO0hjoYNGqX/0Z8Rv4EHqcAUbyQsGMKwhqjPpgPOxcqu9HvwheLXki1m31
WzlhUdUlhqi9DlIBPyes+JGh0J5PM7+oVoxM9Xt4FsoBG9LaS9Rdhpi5Yo01Owwq
HwSfWBcb0bjC88ZOOzhGUIEZFAwO3d6GJQgmSVSNQGMH43qqeoHBOMx3ytSF4YTr
1rJW4eT5qvC8gpxobR5NzkBIV9099fgBls8vee9rA7s6viV8uIElYeN4nuNiQh5U
w/TrcKQ+QYazZERnRYwp5kYDebh4rmVY/xUUmHkrdaYBeQXO0V13ONYpEjyKSmLS
FHRTRBfy6Ph9i75NMv5M3RxTYNSI/aaw6dKnVuv60PwycoMMPxymsXPxZ/KtGNY3
izaKc26aSGwVRA5KTAO9QgJ0EAX0TWfNF6Ogqs3XLXAMUIxJlQP/xQEfa1vpTw/u
ekW444Z67UoFb/ya91sC+Ize4YthoVpCHCfVZS2fws33S/1Z+mRrugwlmAvzNM3T
EdrsSlzJ43b//3APED+TYVN7GKyoqV5nBhnmFmEJrHzNGty1J4Jn1aKA8Nfs/cm7
SQzBY05KDChd1UQfUGptAQoFqkoamsY070wXcDoHmCBIMqWEpRQD5O0JKMmfLKuL
GWGK2nRrtifDicV3gIOvPRFNR4YPjQbeWLVPcxZAdWIoebutJFqP7GnL2jbP3mqs
rNjTgQGO05j7cAGN4K1ETZgWsLZvy/31w5gVYoShM9/vUkkUO4Z1vN04ydcLcnpV
Sbll3XOtU10EklBMvfXer5hN6h+56msdi5J0kNVvbfrhFPgJEO1tymGW7I9PCcns
Z6ZtXLpTa88CUmj09UuqXnxHwbc8cU5Z9xGOOpkKgFhyMKaxYY9kJn+KJsy0heER
cW8VqD2WVclnrMhMolapf7wnLA4++bCkf6YWPJD3kIGa/ltlOt7RZsHirSvIvt/T
QOtAlpZxuRhJt9wG6Gafc99Oe6FFqmNIH/erl8gR+J17dhWluiEJ7udyBinhUuou
KVbEzf7HO/A65GeLEDj/ynQhA06J2a9f6s8SuNbnzZXTfTLsZVNRdqEqhvtSUAUY
WUND5KAep9NnarMMNXXYHr4w2aosXckQyw3z1iuIe9sUUP0pG5n8YgE+YChQDlCO
X3uLOSInzOw1J5pnnTyJhEMRe5bBew2wxHJ18OGGHixEHInDsDatdbXCTxHzsADl
62+bHOuBvdexQF1mK04GssfXGb68KDiQ8EkAuoLvffBCucEIhMvYNRubP7IoLqjw
QEBExHVHYY/KXPiumZWt2tl6n3uTc2NtewoNYZjbvazGqBUw4Mt+EZN4iPSpdoaG
jVFGq9GkIytt07jjT5VRJjoSrcezx85DqWvGQU5sijaBy84pmq/jqW+52UV3a374
pZ/p8JBfEwbusk0oowupQ9E34MFZwV2jJ3HSG5DdtN3NDKxbXs6XQ/cWDC2z6JJV
niiHp3F33RFkzVklPhro2+pt2nYAuCj32pcClxkEutHH6Bror9uUcfTOdVVhMPHS
MtNI0zNqLREU/pnoVQFm8Car6mU0s4hQAaude3C5JqcjOOaNJ2EhqafTAnSrHvwi
n3sBbU7LwssRsQa2tTqW2EvIUu7+zUpRQ2i/lX31j1d5NLrmWZkR2HBEfidh6Zdy
ZYTl58U92oU8F5xRY/nMfjaJrbxVu63StoSQW7zT8CJhdN6f1ax8lGSTkVHKKvbU
kU8UdOmaP5lAEI9wkBtD3Q2OtKQOd4roXwBjjKig6gaJ2Gos2398YC9swCeSyh5m
zw+GzmkF+r7I9Oa1TVSysQGDpi/TaYU0DU2cG1/wCtbt4xh57RprFv+FcXhpAoVW
ZNcChun8vax6J56vrIWlSOHPIqfnmKLz7f6fh6yMhJn/n+LGZWBMuwCvOsII+Cv9
igjbb/YR4MrjCriNf4XF6XYctNDWblsglKA8UErONFOOqaZ4Cjy4uTchmIyCs/vO
PxO06vn/ICsqo/TArQA4efYeJHr1HqoM+9VFvxPOxbywBjwXRTEvf2l5xKRR4Lhp
AvLetcyrpDS2ivJ3NmOsZ81+nGb3BlAt8K2WkTnU4+CwMh/56bmpz1kkS7XiReE9
I0uDK79yVYJbk2Y0vz/OhttIDY7pjS0TTEyRVeGiOluxPD6FVmA1Kv2QXfD/PSF9
kRkTMTYFM7sAA0HfpcFeNR2IDVm4D0IX64HAtfAkQ8GSKLDEWjUqP8SRmntq0WI9
pn80nslGHwa9KLnogIm5ufeTNjyITJadLwvXraL2dDVB+T6ZE1hBUDkx4wVR6hve
gIPXSuCVIDzIFEOIcOP3Fh7VqmKdjsPrQlfKA+UQ6Vl7GbO7p21zY3TNhsmUJwTX
5Q67YHYw8QCaNapxqrsla39prGvtiRAkgrHKpjY7M71FyPn7ywd0BLTGGRCuxnVy
7MQzctO8RQGD/KUd4CrI+ExcMDhmwnlBGoBcep+/+UOeUIxTgZhJ8ySfyNUn/xMc
FkGU2PgSYf2hFJCbXvec1izbdrHkSVP7S1x1yqf8vKNyjKbC7zgr8lAywDxAzazo
9nP1u+DKr8C1ZD2DLgqB6L9bdP+gGUWQnnQ+kbeX+rYRHVVhOrLU1Ilpt+oCzTdH
m0BJX49SbQ77qTc8aCQqLvRgdoGamrlsUt4FzA4ckLOkns7jnHDtQR7mhyiO+KjO
oZ7AwPnKOtbgzRdsX+/z2C8Vh7rgisbHefHjfBqK+REpOkC+ozcFcWireYrQgIcM
x8iOaogxpqTD62dWwg1bJDjgbPiTr+lKycdYPqb5FhNVWQwlnGs8UMZzcS9yWroP
UV1wKkN5uRPUJToZIg3kL7GWscEmKYy5s9s9+09ym3rBWvaV3R7lHfJuUuvK0amX
pVx0V6BE5zIYg47J5l/O3RLuCKMGYD25jDKF0dye9MjAwosqbIqNgg79mkxAu58t
qaNFb4gj6Pjx+07Zy3MqBVLaL5tk6tB4F94bVIIH9iP7jIKgzx3fhuSLEmDWSsLv
qOuZftiPO1ORnEJkZJzmD+a/2WuZ489E9NFILYCj+sBkIXcfC/hwHJWERxaWky+J
3DXlFAsLis9j4R5Prs6fAqG5cDgl9yHl8bZkpRwdH7Ir6OfS9p4nnpCIWNdhEtYD
UkC3EfKkSQbBVzY+dgc3TllCJU7CgnAHNhHsV9KeV5shzbsoqzCss/vJqCQgJUti
PA50FMe3P1V1coT8nePUW6t4VwQlpnHiIiYa5dXFvL77KLwal6H609uPivoLgVIx
bP9NFF7QBYKQz6mSpfP3QpqS2PRaaDQjtfonZ/P8vDVNHn8bJyq4wZWY1OnSmq53
cmBMLw/ZPruQssj9sJRlWqALIetXTMiWEkyHCI4vuKckQ/9U8hYa2ELsqPHEjJN2
gP5+O9MauNh4YFibJLTHt1rl6DntUb7ZXgVXzLV/CKGsnQqpJYNys4f+oWWDBG3x
ZgZbHat782YNnVdWuZnj1hsN3q+lPmmO1yW8sZg4cAvlgBM+zokXCuz7l9nFhDes
wBSIkvEXVIc26YkESmEVe5W3atFlQxrI5l2d4tBz0ZfjwAltfufAW/Pa/mRGQ24m
pKZ5zkgF6GXMtixTXoNKWK4axcy5TxtArsaUHD/z0HoDGzJl+yDgtkeYAE14NssG
cy7wgyVoEtW/edTe/a4HVntvOnzqittmnAg0TKcy4Wcpfjkt907aUSqZUtXbUNNz
3CEGd3VcOg9ZJhC6n2IRuvuakcPFlmcxiO90dEa9Z2yf51O+Fv2KnfsZYnjXkHM7
9ZCCmd7U5seb1NDxWP7XugGicDHVzRN5vG2TgjHB81vs+Q+UYe4X6bJgSZE2/v7H
ODAKxRD6InGod0icKV1LqcQ+uPh2veGKiojNEaCGGEpwFfPtSPDMD24X067vxEC4
GR6xXPU/VAzDkBZrqrYaYjAs0NEUMjFfY9SkMR0L2El5ELdHkUqT1Sye7PSr58Bk
LRYO0t4Sf4E9fM/8FOe5Hgjh4l8K+zt/MqcHPNo0z1RYPHzUkQsP+z0lej6A1Wn4
2ra99AvS8GY3qe3INoVBNMKmzVji1yMW1f5NiEhnlRyjM0nsxG0ksLmQasmUC7Ts
9Wh5XNGynKMKx/cJN5CnRbfYXF8nngbOR0tyDkSPOmsrBvFfnqN7JvPaXJ6EBwj6
Hj0EW97W7Ocljl3HgeWS92mtZUtJ3KB6F6ZNzSCphDSZfRm26QuMUBuEP7i1+by9
Yoa0ygIE+wpyyhbpdIR72nptHOHbRzp2KPLfMpsV4ZPdrrWFUY/GkNk7veeEP0I7
6ZaKvGkXgz+GFYtZwENE+JEMdZIe8s6zoKBA+RamUwu9ziJyLgGVfGcKfgka0bBS
nn6YUgWbmYC7IbZk2veh3kkIVPdnCqnCdIew2o+y/5VqKWwjtLm7HUzYwzOUGXJu
WBb6/aiEobyjjtZ+H6yll33Q0qI6EjThqWVzjTkrx/3ulntOx/7lHHK1sW07/NGq
uNK/gWpn0ettQ0tojC0Dh4z/SiQYKtBs6wtUub/wc7a2gTbvjhOynbf9e2yqT/Zv
839NzsyatOElp3u30W/loiez+4TZ173wmPvUEUWfit8IKSFrGArASmf7kqtwiFF1
2KCIqV+oC/BIrRVlZWRaLmtOPaqPicS4y43SgkQU80L5OGwg0Xl0ce15kG/oSSnv
17DFZw+hOt5vUVpeO9K1WY/huwxBfO36jFsRyoYPL9AyYJIslTuATrF6FN2xnaWL
paNJKKoMu5dGE+/OHTS8VcbWZCNjs5xf1R9tqPUYcOSt5rrJ63jAQPC/W6PnzWkn
a5gFT0wa/yjkYcNzSZKPQjlPv+4St8Htodr30CnK1BeWIH4Eckjt4boOBZTrTgff
uuQUGR0lrUhdb3lHbIeR0Eydha2uYc399bFH4dd96oqsKB1/DZH5MC+Y1gq5NPBG
fO3kYJBpkrFzD7HkDJlEPPcBQhnKUISh8avreE9fyom9dRh7kPhwlXQwwcHIzyXM
4Rjx8SJkPe3sLpsYQvP3KAK3JC7btRKFFvpXCNY94qlfsi0gndi4k+bH0gjrfiAq
JnFsRrNZ6+VxzyF1zGzkoKa6oBKmQw5+uMn8bPIirKCzPrdyi9FzmPrB0GvmiTtx
hMizOCt+GjwFw2/n3MrozYv+D6I0wbBvzq6gtd4tsfanP23Aeig+iWt304MTWQPG
zhkAmTEz97oXWwal/zWVpGTxlJek6mqw71PoHhFGbx3YofOucJXQXyuOOXwsdCzy
QSGk6OeYX24iDgsIUmtpQJ5ZTImOJZSGaMihMyCQqLWnwgSoI4fD2/8OGCbRqsgD
gmO9m2pOrh6iGJV+WCms4fVZh42YCAWER2vY1d2kAbnbXNrJ+2ucxhhJ/q9N6pmX
LtOj82fTGFPErpvlGq8a4l3uZxraFzvbA5ElR6siuzWZ6HVHe99c7G0uK//VbBIW
DQ32kZfQvvLjKARjm+L+eCwuZWh+fYC33TfMHVqQglJBLJwmcEsacs4p2+l4UCpe
zeFCPs6CPpjIV+IaLBBBfEP/1UvhxHBnpGFwZwRa/nJI3f61PgCTwS4jSlOG/n2w
OrS952Z75f/EmQc5CdjlTKYL/BQvxRjh6vehQjlvNyWxf4fom7Emfz37A9Ezih+Z
Z831vBRhNUHYqlGBchhe7Z4dn9l3ZWJDmLzfx9/auLlYpkV7En2NTfllBw0qww5K
zizef1sqJGuVE6gJyiTqptiM69t7b3mznzrzrslk+w1Hi79MU5pisFyO7clLGvOe
G6YFdGAhQ5eh/CLWgn94bDhRHstbRBeHm/Ow9OOjHbvE0Ih67JMt52ga7qo1Wh1B
sGSzwGJCc7T9gsbpFqso8f4Pkc1NSVDBVPVaBIByxH1/jEL72nnx6nmgGHQWTb36
cc9Ilukz7x6TTExlbVL2GF/YulwzTgQwCfvl3tLQhJhzq9AScCYy6nua7yga4l2k
GK6dwrJxT1+3GtOTKIQwxdtjH41hU3n255GJ6PupSMWhV3hP0lellt07diCHgzem
tj5eRV0DkJu9LG+JKQqlRSStHUA3vdd7YawRz3neT6bAG66tp6d6njX8lMbNrwfg
uMSDtHK+3a6pN9jjgwyygkSIa+9xoAnSFiTsXCYEIaMQe+WRSaZqpSC5ZR5Olhoh
e4wqQl1c49DKmWNlLrghsaRFAPRQFZ8CCh3w/e9tGKxRTpqRuWv05moCRMcuAVJO
9y8iVDTL3s9utCMZNpCvtawdzl/OpWRWyvV/OoKIyinu90VLWdkIzbI0u6TWBwAr
BXMfTB2yFNqUA/eEgD8st5KDzr/Na6octfBtkgHm9TLI4EPhQHPtYxAPD6OKrznq
iyuPTBrGlo9hln+r/SzEYbdbrfPVrKvrgIFONoeIPo4pkjYnoaJ7oCQV1Ly34Nl2
O4ptLm6NNoCTcwc7ReaWUTllcIn1+NT7iK/d3sykRQ03vhwLn7tKk0uQjdGoyOx1
67jbvsur6M3jF1qH9oJDAs4oNCkMWj403LMG296baue0GeA52taeGBD107V0vHVm
RXnH6yMebCOliWItymUzkHp+kg+y6FzODsIxnZH6Zq7tIp1hgpAFEdrdxeRjE90e
7SAG/F8JgS2zffwKORnSvhcZUDY0mepSGnHXx6sXM0W49z+f7M9Yyf4BizHCS4T9
fSQWPggOgkNWYo/L+tNWkZS+i2KdO7F7flbFYNo6kUaG0TDxdd2dXdup+yvukcxk
1WEKUxXRxImLtFlnPFN4FM4wjLkZoK2XtQ3s3YDyPAFvItaYSr3qzGtp8YX9Bvk7
2k7lCIsC128MLf/4YV+ZP9fM86xHtC/u7Tr72sZvU+Uo97pO2X8A5LY3bCE6lp5p
k8Sm1GxY8Tyb+qqiHXSjiPB1Y1+GnGs5OplE6zkBt4axBxMNcaLniv5ancE/GRnI
ESFFfdKFAMC5CKjbkVFEfCy999Z6/f9w4tyf4E1Ddy0MnSesZC+5LFOSe9J6/kwz
4wccPSJe+onNltyf6/GXL9s+26Y6FNQULkdRg8haQe4ZDW3iz+BQVMtUY6ye78E0
Pwu+9rt42K8T5kWkqWwWvlaroZ8JRncjPz+be7I3Lqajfvwq1DvmG4R17mzmIHyT
ciV1Rdq/zde7xt8ezBOWLXHAgdfqiIlvEAHB1c3g2i68p7bixa7dcF3kbUwPloN3
ZIFY6HGxKLohG9UREUlETGdPozyuL2Iycin1MGLEm3n3qNn9MKuIflMy3t1hWM90
WithBGFEJ3EsOKLIb/HsTaBlFiJAm70AzUNKZUleATpQax/CgEKGrB9Au3zhBP4N
UWqPLpt4Kf8DmiVO3df97Si9Q8DJdIw5KJgMwBPPfODeIg+Q+Pk1xwnkhjp5izQk
kUbCJk1F8o1lspckcnZe9NMgblsb6BO7peCU4Jagl/w/RMgHDt1t0is/5dljzUFX
aWm1q7e1IVE4UVG+wfGOjlER75v0K28eODHpaFd3RHH77K2DZovLB0dP6iiC0GP1
0gc8llKsJYltWOqvj6UWIqfkVSMWVUUQ9aw7uJs8qfINvyxltOkFstNsx3niz+Ew
NLqbNLJ3a5VfTx/BhojOcoXAw1A5yNOUxIkf1TyPJZ3tOJh6j2B09+g+xJ5ZuDOk
/P4veLGsmIz6KbNUq1+INGxLx+sl+Tyd4qHoRRdDWahqjKjInOODCUe4qfFDVdWN
R4dihPOHCwNfSdNxZOELQ4arpqm+6YrO453KrQggzWiGBk0hxdEN4bxEF3niztJe
8g6TQpAQKjrvoLwnMCYYgNlr5nbkjfFLjrnFU+hfGQ+LJ02RcKwkqo4grzGX2e5m
O03cPoVI5i5RP4jzHNLyNYb8+trcolIKuUVGO8i6Vzr7TQxP50mFE8IlDu6wEwIe
XMMOl4e4Q90eTgRVXDMc+wcx2XfkaBYU1sUDF5oamZra1H79HdJ0OOkaHqDYon8j
EgAgFDIYp11FyuwzxUm+9x5nnnOUb9ojGxojIAuAsz09z4EcKlcejnWOXpj/VnS/
SFqweicSE5/2QavB9wvcWk1NnvKTa1c1JbwBK4lO21SNFQXsNwDks3pDMTXeo3TN
sr1t0mbMz3uBcYEpmjuLwFT6bcTjZ4/cVxKSUf5+fWz55s/Ooipj60Q0Lw/9zk9Q
P//5BILydsYtCyUlG3mV8zvgcz0PncE+hLLzwArPQ2D6Ch3mi8X9o1BRx0YL4ocm
Sk4Wg9R/W0s6Z7aN1v4nzKAwC0SwgYLfBBq9s0XBC7ICO1b4wqiQQvRGNgXdl1g7
LQGFC2JG0jsgyhnCSDvzakVO2RgHgXOgOZg6e7cdTHDBjFG2xvYQcpknl/PjhsrZ
3tooQXfM9VD/1jmb91lDAAhEIoQ22dLyjX52OZ9l2e4Lopd/Et/G2w8C9A6y6SBL
tUzx5V+f3mao8pkBAWNSfUokySObCWZFfdqFDepFA+8Jr9vi7xjtNbh6731VIz/T
fM4/dnSlvLoxajOYF9Fs4hB3S3cNcIbSs2dWH4+xjnMbMdzwtjEbChN5LGE7iII8
rIVhjLWyt1J61jqzh/f9aWb6oqq3Sff0mLXn93s0Z7uzadlgcU5zWWEpIVX+WUQe
H3JwWJmQrrUU4xQIMEcHS0v52cPqQ5c6z4mKILq9gvc3uMdft6IMlbXLxfNrEQ8h
TLG7GiK/+C1CpmOIAI7u0mrTMUJq24kVRfep4sucV27OT5wrBe5peiELwABuSRct
PnjNk3WZtzNf664+W+PSBBsWHES1GXXdyoZzdmVbXCQs+zhItEG96LAmHydG3nQt
wDEmV68Qb44JidCHu9RkF1frpIUJz9mWsnBL1qib1aBS3qYaxJ8e8UAIWnV7p9Bi
zaew8zH9x4E4L+HX6/VT6K1hAlfIqxxksnwxkLLR8tRV4cr0LfBmtc2NkA69chOX
x4eTN0FAAxLKvYVr2l0MvHRQZs12DeseQj0Q6/x6aIeguZon6H4C7HLxT1E9dd0I
1MfhzHjrXsU0hBu6GaQIT1PSF4dWB2hu8map2A68wyJDmCgyxgmXf+9MYwbJ7hMU
jfqtVvT2EAq1aX6xHIaHT4QlgDOLpmPAv+DL6huz1xFweNUtrjlvzbMDTVW5Bk3F
KGFEVPveRK1pIpy3fLoBh8dqMqtUn1WbInG1FLIxydBIW/y8TQDyy0/KWBI0bCcl
eIN425ca39o2apjUfGmwIR9XQXsUvAwl1jSmx9yh1MEvW7LetL8De77deUU4hPrg
anlTXLpECF1tW6PqA44iSap10UQP9/MdckhRvBN0KQo17koXpq0LYqHHIqSmdwMN
37xcXsZerX10DYLPzCAolge6OMr4EMfhiV56N8mi30pYRXd/GNic5STv7nIDVHpK
L1VPl1NUYbSYy1UMrzg+2FRDQX61dwTPXLNzgCIne2ECql7rja3HiOQ6xNERI8Qk
h9ESu/CRbhZemcmdml3v1AdPwuuOS0UwU35sJH3/hLR4V49HtDyEOKuObTFS3vLC
yIqHR5lTRbDzfQf80AOp1LHIUz0EPrrf22aX43ty0swFiuAzGMF2Edg620plDmm0
Q7OXiOsT5nw/UDPhNMJihB7fym2DEANlIQd5VDviVlwKcZ0CaByd8swk2RhbyQ2/
RQ+SoMqE2orEjR8rR6KkHidluLeAwosX2EfvSeI3TjLlb2RxOtRDl+Fi6TRBJnPm
bKzuO4W/eiSqOrlYW9nWZ1uY/RY1mq7qXfuTMH/PKSg4Ld/1gMhVDvcC3qBd41fK
RQ2RKLWhZ+tDpG95Z1c/QD+L+d4zWOv8ZAmHo3xf516nwSdeUGogzyxCHpRwJ3Tr
MRbsEj9w7bm2C8B0t2Ao0hAfm/BBm8BkyohT1KEPt7SvIbubAkXi1QUgiCtCn9ia
ftq5e/vd978f+jCvKgSjBQFcs5m/djlGlPaTUtt9XK2AYN8dlHTQzxDU2n7uePvB
azX9FP4kq5bBh7pApsmVwsG7kWpVnDOYI1f7gxJgUfppAFcwuL1my/JAxg2klO0n
3Y9FYBq+udwgMoCosDpie9RPnS6s0hBwttg+zC0/9XsTL/hNC76ejyP8CXsLuFDx
3LVDLDEtsfKFg9L6EQYmaFczLK0JWPQw7773lhpoBRLtsYGeEOXaZNyiuMAhu2sh
dhfIZ8CJbELNdRiUpTYHgP9ssO/YHMIoM4HEyVTHAeTDHOZwneMWXARcRrsHkXjp
DYjdHWbd3A2dbNTq6iVL++I4k29+TpfZdhMMvVIpPLhVBea7f7vgNaMm6yaSN+vS
4SK/n8BMyrck64JEdd9JcqhtjdfWd2Z216jcf/iINakK056aWZOHkA6Amuy27sIC
D5B18fEgHEi4Qr7OGOb6dpH1q+sHy/waIgeSsNRCarh0yng6dh3o467L5cD0xe/m
VfbgRL1NeqkIrg+oMlGH0DsAm7rNBeaSO8R2UQqERI42s6sKJZj1aj7cb7fPRKix
3bzrnBTin2XPjh7/YQaBOvsqHcQZdiMsIcC6Ld00gyL/WlyiZR5O9K2RKO23hLV3
1zg19NjEVS93fVwsCLQ3BzxWbCTdGj4qHljjQ3H5dmsc7QukIqOSzclRomGEl8JA
GSuPSGEHiEXWVYutA9qUhsAxKuaIHNAGeSW4CxqOwvBWmi9Y1/7dm9AvSOrv69zu
O/s9MDQ0lIMuLjJCtGtfHoyaM/h5DyTxPJdNNgJHOxDR53z7jpxtJ/X5dzXoyF5U
BorK/Gb5D2JcF4Txgz28YyYdYKN8+p1xv2/1hP05BDUcUBGQZWewES2osLZHUhIp
EnVZedvz/NQDP6XDxRoSwEGMow1+kE4YTMq0TWerH2LlsMffbGtZXIietmIu2S9X
U+lgYz7MzhwaCdfSGtlwWF/vl37YnFLa7b51S2/EAGLH8WHkjoS3bPRrAi4t7Esq
q9FRUDwCVekgGdWJbad/w0BKgkaep4Ro+mc1hSuciw06Bz0tVTJ6JoK+Hp90QDZC
bgJjtIqkY0UQwimnoQ9XX/ZkoKmhPu3MNM6PO+SVPK+CiLrjvz82ItUXRy4RNrci
o90cBUG61jw80bAV7+AdnMGG1R8YoosXmsHIA6iH6ij5l1K0H92vtfvOcPHYql1a
tVJ5ltZWVrB+MFWmkoQ4WBAxBc7xaf9Ul/pokUunTpsQLJcWQ2RbGTmuTCxAfohu
JU6sopi/Y5j1zshVBYl+xphw6DW1gueR7SzC0XKcgmEgFqWBiKhxVdaycsVfF2Z6
NGT5RCBI5DflVWitlF4m/Jr+5Z3edjLkH63GCmlbZS1+YBOKdwd67ut+oYBIEby5
bsRhToOmnW0CQ+9QM2ffCmmx7cgMkgYMnhTRLTXDuWOoS0ywBXRuyuOQWyLRtmX8
EYYJ++U2mmgDoBs/Oo39Itak4K1+/lixvG/j7CViKXPovECCsTiEwrxQWxg/B+tF
ngRA1r7qKc26qlB9jiK8UT6LGxg8q0uhDSoVppX8XmebJeWX4A5Z8ztlcItXWqpz
G2YQTeqYQGWVlbZRpVhnq0oGT4SjvhB1YXyXDg4HoYz23hFNusrn/dTN/6oMPCRo
LKhdiJKAWyiahU3oJYEkLRapN97KsyR7DpZQRrF2kY37KPm0Wpz/OtBFlDsYXVfb
3Ukw2ezHTHREavjZSCvQJccqL8pqbnm47zIguYDw9GN0iSsPesXM5saDEaHypW2Q
tcBBKxwNrF5dzOhn3hfoEqtnNGazhjLkb6HcBm0QVKx9qcOjYrayoPO8Tg4GOT/a
6YaQedmUDgnoc1meR0RYgszeYU6A41VP7CDXTQyLOLwEnqss0wGnz6Pjxp+r6RCP
EHv8o7EWdQUb6T3ihCtGRSFBWo9OiofkLLhGeQiuiXUiV9h3QRwND6rwuNhOOJ9m
0xtbnQwaRIqIgp7BgFQLMTc2BO+NdntjmfggF+m69R7dF0Jf/2/mmYwR1Yk5/JY1
B9ALxGCdYF3Dj1VpVp9feXR+B5RdyBd8y0ZXzwEKrIYXaa4CMm7424HBoilq9s+a
5TxsQCHD0GdWiy2un5Ekgw1J10T1B/+1JMdAfZxV/dsRdNcPwOAWrYqfQfFjbHtw
ypqqfBkOKPJhEm7t1TrwOpGmjTrHF3slWyxq3W8EzVxXu/+4ppcOYVJ2yHS3yiYz
n0PLREi0gjhFXG2CKI0YXO+A9UdSgo4bXmb3YU3gcKCqYQoQ0OAWudYtTKeLyTGT
jgskRpCyWGD+ealuYwktZJRVKwh5lE73IrsrAadMzajo4NIhZh9pN9mH8zfP2QKE
X04gRmSL62HJgoxmkrmQgktUsD2KDfNysd1yJ7LmGpZJwh3Nqa+nesOtanhq5yQn
ixbMv7HorEj2jqf/Drau8GxCldr3UTqLy53Txoej5g6LAi4VSS8mZhTyybANWlVu
wsFcXjOVs5rNk24+zdclaKd9A3W7Q2o/A3r6R1JsU8eTB7/6676vxGda1mTIPrQU
aflILBa1oF75a9thVwYH4Il0WlBv9MoHpCAqVTqTibhvqzd16nJxqmVzA+HqgcLN
K6RyWjJPReK9BxSiDYtZNiU/D2MjPGMTSFZyJky3s1lr/pAfPri8BUJ50oge6PzI
qYCFNPP1ldT9EczlAkSycuyoYmj9rArlr/utvt8y2/1DkpRH1/WpUcHVhVazP2Vp
tatBe9JWp4Uc+reFz/DmdnGmJfj/UtLSpWOhfjayZy9VVsfzaaiDqfLIhtk/MnvY
Al9Q9LBz6GmkxslkN5vPu9LE1mrrOO4SjZSHnqrm9rxuLAFTrzrsXoY2xD8rJW+q
L7JC5b78d14Xq49G5EBn5qm4Z9I45D5y3VUig9Wp+P8z2xpVLk8Ayyf23msunK5n
3DflO8ZzXYEdtRChGKkeLXqnE2/wZ3rznZbxCr0Rij/W3PKUq61rp26If2sC6mY0
3WK1M4/4Y12hrOtR7doYT4ofizGRFwciNmTeaXNa3fBSFcGQLqUdHlDDNixWLs0S
TN3MrUyoWvyvQDu50aoIDdc7j4OiloojhSKcn+O5jL+GMMsu6GFmxxNxkysHdLQN
VMYGYWCAFcCrURjN8LLvyKDesZx8EvSGFbWnDo6jQ/6a1cw/4LeUMQ00x8v1tNvH
WtkTPEEoXLDsoRzWNvh2pfRQQ6L/A/uA2FbU2G7Ng4jSpPW3N4FB3MDm/JYVCS7q
sIshqirfJVR1sPnZ+G//ddV5H35UcgtEAszn1vpdc3uBSjMe//PwjDO+fb3RuZgk
uNRUHOtWbuvdY+MxYZxlnXuXJF80RX1Nst3P++CHcS8eDafKcvLNUauKsbtfLKUd
56S12Shsmxr6Uatq4Y17PIwOi8gUDm3Cfzextq+aeN8aHfYrtAV/0a5XHZCSLM+v
PbVEcI5JyD1fk0RA6waNRd50gryA6sajIMsclH4fVoxgEj9MnxhsTeR+Z2x4oNrW
88MhV9IcKO9Hxy9vu2r8QzWgrcoWKHjrRl3KST2ZNSIeIznwlaRfeY5jfTTRPck/
/aCYhi4rs+rqmDugW5FUg98Z6JE6YHUIBbPfBgdSQ1u7gQhh5DVfTiuqg22QJLO/
0o5wa87vB98dE6si07X+3xOWNi3KhWw0v6/Ydi0eoGpJBtZmGm0DnS0RMI744zsE
w0Z1bN6sIedC+y/hKydczcqgfKNkCsWOB9rdTJ3ZzcnNN9KRgZW/nI3hXsfkhiwM
R8K3Qiu3nnrHi1fmRu4omv4+ydiu2j5jy89g4yCVZxUktVaUyvCDoEgUpG3bdaqV
Merv737XmDxWjSiMA+MCheG6eIFpIzVNr/2pDf8wqc5FqiSY38rn3UrGSvk59s39
kW8ekVvc9BmHhbijfpLv2jllt0LULs3FkxyxFN+0/y1zRA1QI/xLAXTHj0wtsf+H
Q3Q+hs2GbyvtOmx+8vzJj0dpis0EaD4Ro74v95umwiNb0hEVZLLRZcTonYCN6eyQ
zir4FffRwR0iqCwVehdUz5RswfQ7yZ6PV/jsLCdrIHHBm5Ru8ClE03fdgX2r6jD6
XrikGn1kOftACYw8mMLCdGIy6ODBcOE1jnLNcmPVwqGsgG8oy1g9waDXUgGIZwnO
JwnSe9usb82Y9PX+6BjIKzeLvNMQWweU+opt4Evz6O2E8fTq0LECipwueoT763s6
nsCw/9AOLIspAJSK593+zJ3DFYhV0lAKwbhj6+y4g4tnYRHf7daMgBhZw/iFO7y8
8SR71Xwzp7oNJ7xSyF519DG5RdEorbg+QMezjGM+8M4ELM3FlSne8BRgIYpOXkOU
KfLvFoRi378IQbVopKsToYWMj0hZInMaNs7cWCOtprA6FG/1iQ5qcWLV3vPPceb+
outtMxWEey6kJhsUvP03GEGLP/Omnys9ZqnRULsgjMUtqG/9I25rtHDAj7ljCOqN
0tuhRmDRBrut2Hte9A9g6r56y4KIbPJcekAdFFK8Q16J/92eE4XAg2NgKoOc5jaY
jZ36yWLigUpkwVca0axVFUXXfKXk/jOwD+FAfgNvMGmjkxwNohSa3r2O/PqAKrnZ
fe9H0WGIbTb1+hyHECi/UXDPwZK1dw4FVGAXzBXcZlSgyWxdobKknt8bTmXtl09N
LuBU5AVpJBAne0Gwq83VriiCzBKvkGw0C+UxoXCcgaqXLOq1mSpAa5kDfW6So4FI
IhA7OuZ46EIDdX8t30iLbFY42hwhfJb58XNgZFWfZvXhLmrRIngNZTL8lX070zVH
e3H9RI5G+aCAAuo2fv6L5TuSuMyf7/oKHh0POaus6mluTYqqMpr1QXBxypeu6F5H
9bOv9Jov+h+sSiz0Oj1ilBwA+NoYR+3ZvcDwcE2sKePISEiZGMNGdlIENPKxCqrY
Acgp8q9s6+yB0hGvqTj47fiY+iGGyVp0eYfTOz2rXPLBL9HWMreu3Fba1kZ9cA21
9K4WMeGVbmmKZEAkYP3IVsJPaGXrVlDl9EQ8UtpxN4Shd7Z9w5uyNEFTmRgYjwPw
7W+L/TgmiBnsb4BXWdAN+npZ8k82B5PcRTnHV/Dqb8tXAJeph6pNMw6AvM0jbFhM
fygp4R69xLRs+V3d10TxvNI1SQNK0eHV5bijOH3EFlVoT5vSMUdO6wGi3ln5nDL9
FMNYjTFQk4WkwZzLSXR7mf+fxEucW14Ve/JGcYHUYIEADbO4i1MWQ2jv/QnLobLQ
D0190aqYl75d10nlbT7hRBd53UIRc2TUPe+zMgkd3SEeUUBUwcBEuIFeQMO2uuxk
TM8gQZIH1QXz9ZvG33Qi3a0VCQy6GgNptLTlD2TdT7gJ7M5nydpR7/8K1weiZhDN
fIP2PMFFEZ0ml0Q5EA9FS3yc04qooOINK2xVJmzLe0Y2VBbAKAo4YSNaGB/cUC1J
R8CQqR31kCk5Jj8j7WZojsbT2XdgxDPVRnJYMSt37sMOKWl71emJR6KL6bf+AnkJ
5+ZkQKYZAZ8Ol/CKtZBstUnRbxQnBCKd8pAn24sF6UfcUcSdEDreazsAZdTwk+s7
FH3pqX6lsGY91e2QE3YDrELSHpUjAThMa54swWNA29bi/GtGIGQZLI65tkaMzg0p
k/FfMM2vlIkLotFcTMryAuN1MW5weAIkZotNlb0FEV5IUGiw1OZi0BuFCVl8ZebO
yNg0S51NP5XBTbD5tli5CGbr4VzB8dEaQXmPkXkRBDXhUDGinrh97dlH1XolpkG2
Xpyc4GOjfH9uabanrvjIt2qO0FzF642jMNjXyKbpbO7Wfix+RTMiBL+uhtiB92j5
V1xhn5BmJgIAU2XnoUMgBIhfgBCccQJp1pr35gPZJILxQS+mPuyTni9ubK900pgs
3N8tptMaoZGIrQSL0najzMwolyyLTcMu5gXRZ3odSA9NOHJuw9xtqCr9phza0Va9
atSiWXFI25y9D9ynn3JVPWILTwSmvZypsqnjYt8PT7CI13MNsEw+67FPDV3g1Uzv
poVq3sQv3rzpdjGZI9h9vCfztnuUYEupJL9GfUE0xcVlmAjhsyTdLaPALOZn1rsu
4qcXlBzpQvdsSlb5O2tj5Ox9wDxIS/owsrUwUYa2KOXDOWRO4nw+W3dsyOYBf7yV
7NTmxoiT0NJTpX9+XAIcajukce+HRQ4sMWP+8hQ0t7TMTnIAlY8+j5f/495frtIA
vNd49yIGVmrqcpUbUjQPGJEcVJyPSd8+HQdLux2KLw3vZWtXoCdmQtHjIKksecoQ
HMoab8PjgmtgT0uwFLN6lgfJAZMNS5ZeawuFnuEoKw0bbVM/m8MEV0nQEBRHrrNM
8nNyEITM6Mx0c2IwdU0WQDLiWWoUXbb830R59wPToUj0AIGdMwnuWVAr7oYH6Dym
6wCFQIvkAEA5SebmrhMx028qe30woKhJi+/hmEpwA3yQQ1rB9D/ZpFfo5zrfHnWW
k/5c1p10ypxwQwEkBIqwK8eCm412OCoVIh6UfNwZH53TBi7dnG4OA3a7Y2ZtF8Oa
qrVcC9qF3AreKEvqbbEk0XQPiK0UpzT7LO3TYCPrGLQIJRLepA+SQeYs64McKLjB
XVnTpXmbfpKfBsUcpHYu+vMT52QM4zR0vN3B4LcutvMLRZ3cJhfmDeC6KZdlycr+
qZ9WogHhstdv94bYc01ft5Ih+8uztQfCZsYsOPL7dUKhyRn8d1cIgnNvWHtvJmS2
LKpaY7ya0nt+mX+Gbjwor3Z4z+NSCYCyUQEUE1IHIxriMNWz4p9sObzWytJKTlpz
+qVnf8O98JnzX31WLqM258wI6QXgydtgQHoE1htJljmCNXvwJnGmDKPfAcUhzQrr
swOHZLxRaUC46xCYdSd0UJKMScbMsMDVZguk79KzmFNjHe0kS8qOKMXwRSjkwKGR
ttyKx3C+52yw003gxA9l/Y/Br52aHGhAXzjpGa1zEuDZsTrczx8Duz5s4riDofvT
j2rQPDuZnqLzZRYmn/nZ4U6+CAL0+08LVRkScnjSInRM7mv2SSE/QGHxjhEvtxFh
XvUQBg1EdZxaLxXoS6yXUxA8l7/4mVc/VtR9qzahMzI2VuFS4jvMRBAKtIwtGHYB
n+3UHpIdRuUthxYrpOdZq1a2t/NW7c4LFv2DNKMLfLHgqH2KYsE7k4l187e4LNpY
Lzq5wmYue3eDu/PKDai1AVVP3gDNBmjsWDJAfHK/3P863ZZ2KI94BM/R0pXZ73NC
pGvDB/xafvisQCIDIA6qzxfEzakV6fPVXUY0CrcYsIQ9NXuuFETAlp5DfNv6ixZw
IiSyS56JKNRrynnb+PXPPTEf4BT68NaarJWLapCcyQeKwAyV+7J9lCzCX0sw0vXs
zZOoIOUgZhgyjoQg8+YevecNZ7VKRKfGopO/sWW48PItWBLEuS64Caxi/B/WK0Eb
zGRhsGQiJIywdSkmk0/K94bOgCrEE/bKWYvPqZRyVu6oQTRc4bMuObFFB44m5uwk
0SleaR5t6XYUELrjWeHsT2f/uoVpK+EJM99L4yaF8N3pA7k/1xUzgJxR6c1yfGwi
WXmYQ/MYEd09ZBkSa5xl9Nj3j+OLmMQ/qLgJ4+UM0PqrPp6k0+fFQkUpTm7kqLZf
iJwvOaseARAdgefkkrLPlGGgl1yymWhJXdauobdYK/OP/4SY7khBDqrhgcEIEXMT
RN/CC4SFBwiysHSKYOiO3MXDA8uFbFmcE6QZRLhHVuIT91fx7r3bc1RxkzdEVbZ2
+KBJPgGdUYj1TM8nSYRGhgxkT7CFIpl4BLGdn3nYTNtIqRnmH/HULp0Xq2Z6I5BY
M6Nei+K9ACngjbjeD//+GEtjHZadeCNhaHdeZO97UGwI+87Lsm9ORKtGed6wSW1Z
PaWgVFWHp0Z9i3I7v4Mgbu40YVQjfKrlpu2VcRGF5mhR5u0MbXYcbndn5AfpPfEK
H5t3zcW8KuzktTttGjTpA1IvA8rBB8sAxATJPQkzH6I+zqH321kmt24RAPAtY9cK
ZtcRyg57p9hIeWiiDus6ETc2wEtwoJK7N3Oh7hKXxBGjyo5cQSBUIUo0oEs6559t
T2Tdvf7XP73nTB6OA5TVKWrjvUG2YSyPm/00CzbBXxRKC1JEvwHlwrmW9B4LIYSY
1GFRDTm5zVx2+g8XUyurtQkgDeHmXWqoYXTW+k/Gz0DMZ5Q+rdLDpfsWww1GOJEK
X2s58aPa4+MWpRrGCjEd55XNavRpo58ariryl10AQk7qRbZpwtkYZRPnE0QM75rj
GzwuQEAcJ5/Uf4xJeKdY0wMZPyswVRGCQhCOKSlwYWkvqhNqFP3769EXjpUr2W9S
A+iC+W2E2hQe6U7j6eFNgthleGERCLnnPwufl/rKt2dXsA49F+b0xmzkzBJWZAwE
Vq9A5NUBcDEZwUHIBa+Jwgf1bflIK4Rm4+znB8p3BZgWejY8DAfR42IauyLtW9d3
k+d3haR2EMmn2xWIIIonw4VcSEdo6YVN7I5sn3VEu/B5vMuUoLQaG9uxvSXDgc0l
3sUFR/Cl3Z71wtyYJoIPG0J94JXZk/MnlrP7Hkd29KV/765LupJXUC+uIue1tFV7
ngi5Qxx4xbPG0IgJJOwEajcNQsXsJcapbFGJbsl3nk+vqJpEUxKzsi7jC8mFcGEl
ed2nwqk/RFya5w2qpApv6e4M7E/K1xDltyfbYOjJqf/Gby2jimhvpplqS8XjE5aD
8BgAOGPfxhzXnHoJMSbon3hUih1parRdvqifm/PeCOstREFSlQYY8wb9ppq6Nblw
nxWBVbA0Gur3LH43UoHnRtFkXHck9TqSKA5AuTZsvkAegBuDgSBRM/0nYGHMgJso
izilsV0hykUgPpf3Yx8/PWzEC70fq5pBPj5OxBVwpLSSNMTwdG+5Iz1nF2EMQ+HY
sFDwZiMkoQXn3dqSRwa3yPMNN4bTywyZAdZ4i7iUgqtCSApwIey59QOGJADejDPp
+xllm762ItbbH3i2z3G8gVgCoNfH1+D9oW0Gbb3POndFUiuFvcOFtNcI8807VrTK
ZPvb6J/6JSCijRxBtyBco6uDWHyPw+uOSnjVRJ79wZz82J4Rb8+ZBPkLnnY4vUbS
19ykBkmFz5+eEQdxvAJ3r/Hp5u8dVvpZEJxy+HEyib1m21976Yk51RU91rCRnAAt
5tmgtcFU3QH/VizPzSAzlqQSr0MViY7A+s9Vyf1oHZpGWXijqnwt30l5fhCKMkPa
pkq5QOpw821KulAmOqTbCwmmdzH8m5203Y6HySMKz5S464QNib8pN36r9ZMDgUaW
Z/lpjxk+U5ksspW0efL+mD71dANFHXQCMS3qJYFnG6tAvmvH7edSV2XfC1sWpNiw
7W1CNr11i5yXUBPUf0mx1pJI7geI7Cz4eGoyJ898UsqhZB0TK+sdv4oqc36sTO76
MHlKTAb0Z1yjxMjq+bLXimYu+bqLSE5FknxB4PcpXTn3p0d9oi79A00vkubb6lYh
8zVexCWSHVDTjdEVIfWt7EqzGAb4U5WceSCfJjofBdOAtzVvO+oI9ue3ngp05CiE
XASNRq0bcrd9NDWqs5lnrnVMDL8cHV+nQ+BZtDdo0CKpjPZlt3OlwqJ/kQjNEr4T
d1wJlYo/FI+tZshEyrwUdzlyW10eMa7c7S0MSFBgQnyw4kEPhHYU6riizF6AppB/
VtJ7Q2Yvc28sFKk3b+hJM3H0f4pYh4ekpKPkKmJYT0peOl6Yf2kCFmZ/8LUYBnSW
G5YILIvKGZipUY7yRK051UBnFEpairO57fxEZvizaD609u5ttV45mz3jpV+rDYUq
UMu5NTRn+5j6epwoDLqnQRq887IAoz+nqSSZ2fJJ1xcUovt3f+ayQADKjfr/M3v+
y7ga1VyjEvzxHaEwCxoerTXXuk7BDN1BSJFbGeHXkrfNJn/+maHYidfApC0pOvOi
sQazYZYMoibsoALSzLSmB28cINc/cObjZBGwYxx76sSCQlvYd4p3bEsLSNR4jiWe
b3sbMCfrtFYGMos1l7KY/uRzcTDMLVm84o3ag/ax+j0ECq2NzqHErUZsNHoVQE1c
3bwcqwCSU+JyB8ddsQ3QHk9n4/DVJL6ieee0TTkq5oYRcq6yuIxim96P1PR/ibWq
uUHcGYbq+WQsM+WFzSRyHQ60hfTz3k2Hj/Bb5UV3n2H5CcqvqoQLfaG2nFWetyOy
ARq6/sNwqxP3sRHfAvbkaywqJThShN75n3lVvWL8da9h5Wmot8V7/kNPdSBNMzc5
LbGUR52IzDLquZ+WgXXbBRAdq5tc6I0/jPmzR9IXwglQ3RbYVl1eEYwbbCWdhNuH
2SMaXKuVJKPMmAIirnQYX3ChkNlFMbNUbe+wxJgvPLoIDDqUnKoLYqtyoA8pgTE0
Zj+jWeig83Y2zAreB+iN/ME7A5Gi7Gf99vgsCfsL2E6JW+9bVqEaUPV1IByLG3Q1
OJHPPEsjMMqp4m1mUBoVmMXkqiykvytNH09aZLIl4BuDj8ruPmRyrDWqy1PhTl8d
BfeOW6plSQrKZP5IfLvrZ+E4nSP0nyn2k+Ua4fyrHqaVNj/YVJ9h41fCpjaJGWbx
ptVQpW6zoDH7EZdNU29/Qt9ydg8o8f94dOg1s6NfIzVhPcFklb7goEHH4O/hHrij
xltJH+a2/rHh6IzLOrHKPA0E8Di8zTpQUkZcwWCk4cAvC/aqsxeqVeZzBlsEKdGk
1AxO4+dF/1pwr8VcFx2ZFFVTghMTgej/gavv77Hy6GObJEPmxPEh81LtG9gIo0ls
7DY9hDaA4dVYh/Z3X5T6yhN8HKkp2W22QYHIQMZbYnzTbY0a8cPi3p+K7txu6Gc6
qYD+k0bJV8pUfPvR8+yESjv6lqpIdSPKKyL7f3jdkGHAq2X7sAH++O8IW8xnoFYs
8CA6Ow+Ao0oG6nJQOgCUEPS8qQHnRV77pb+SZWE7WFg7CF38TQJTlyBcrkWRUt3s
zDSMMGYleca4OFSoD6wqsSnkpmOthr0UV7oCeQiqS7Ch1RMThjHS4adEG/JOC9W9
56gUM4N4v+TnPMjkrdjiEfFaM5BiVpwdnUM4CAntZ+PbnS6hMeFAS0/ODXqh4HXn
bRm724Uj6YMU2veeRavHEKBVcwouaszYOdIKaehd1XqEJ9LMnXtSHusCu/Tis0BV
YC3Hdpho/IagnsvUu1Au8j/CcnOzZ/r5kIiNr/axTAx3uIgq6ZfcULEBne0zly0i
IQ0Fx/vtsYdwF7vaC9UBqs871iYmgTdeDjzuptVlGcXiql95Fg1Fx1iv4kzxZfdn
zZClaAJzQB7MvY8mxG23v15YI7WgpaMj73CM6XVTsWTzNLOsiPC78RRvJ0qNhs5G
GEQ/GOvd0UViZ0EuEBvjlYsMvy1KRicS7GVDsFBwBwwm6MbhB6A2wSl/gaGDEADI
t0hY+NS9FzafRxNEP8P1yo82QcK1vWbdIs2+LfVBUiew4chl2H5ZzpPaiZDvoVa4
UBcDB/ol9gaMrPNZTv4Mvf9wIqDTajXgODrr/lSSXlfy/QzaY9vb1BKU8kMu9V9o
SfhRBdhoeV3dFiSpQBuDI2k5sBgStCwEBJy7etmgs6ugAVqjd8uXocSXiAt6py3i
NH8GW7n+97mPynXLx1gJljPEqdbnBPex4sgzmVsExMCv/3S5raG4QM1IdNOxKjES
YlhUC1HgqvVNb6kJ6AFuTmEQCK8FzY7PDJfGU99tIex7MdYBFK+L+0Wr1GIQn4ST
1Cu48LV85qhrozSY/Pu26oWT6SlCbLvzaXkgWNSaWUahsPAXL8acY2afS1QotdmZ
/LAJ0Pe6jIBESRCCLJPZzb5SCXGFYdpjafxZvKiBYuYdWArzFSnAjRcefAikp0hu
yNsVP6tf4us9nzF360GHyPkjXNQTfAkfH/u3Cs3kkzAPNp2fSrWFHxWm3aVKUyIQ
eaJJjniSOGU03g3Ln/aXmQpOnYaF5SPyqUnXAmC6h4hX8HGp6yIntuC51pHtbhVL
fCJ8fZ7+HuQcJRvqoAa8rEQ8iXiLhEQ++lY/VpujYE4afv6qQr3mWOzo+hRzvlvf
C9px7AL8aUPUs0PVPoKLVTmH6S3mYmLCpbc1zfMNxegxEG8/3tEMBxtfi+t5tP8g
dlnSQ0dcLyaXgJLUgaIj25ByrmR60wtAMvRZRSDPJDUUjzjUjLxZ4tMWDxLQQ7u9
wM3+p69heawQOgGoF37/xaxwIYuHlpf3k5sWWYs5nFwpsMoz0Ux3781j+qt6CYh7
gDkRTEYfcJl3tKuwDcXiu7cB6Yfcz/dn4m8SGb66O218Qxdjd3wu7ArDx6Bv00kW
4hVp5z4DIEwCu9UE5YBrcBmPpAamsOT5QKzFk7bneXBB6NmYmZVRnbXOyxBta8E+
uxH6T2bQobxdUAlqXhW2G+d7VMrhfCEM/OYv8kPpuf6VPffB7O2Q2td+27O11SNq
vKLny2KzldQoHG7vYaLclQvbQgAH2RqHIksB0h87ac9Oe0oSVHEkpweR8oO5pK4b
QcKCMuCBvIx5ZfYm2eM8n/Imm5pv17DCzuplbT6mEQKY5O9Xq3s6Db59Tk5+723N
RjBxRxCfnKtCM+VaNNXcjWC0qHBXiFJSthb81uybwiyIcRBtbvh7i3hVnBna7PQE
oV19xnwxvnqkmT/wLsb5KNczWWus82H0RvkdFQ3ah/BCUiqMIIuEzuI+CkeB/cUi
+9tgepD3HO/F5Vou55f9SjzNRVe0j196yBqQAI9Xw1GI/NrTJm1Pfk2lqDFdlH18
fwmO5nh63YmeYKEptn1p/SD7qJktV+f24U8Rfm5FSrKK/nPEGv0CbYghKGeDsN1c
jLd1XcoeecDJlFK+5sRcwOATebpwVtuUD17qbnfpv4ELoAbxSyqrgNt5nQF60h8Y
OHrQvQ3BImlCpZtZ92CVuX3xxiFL2gqFKrgydxJ0PzznFgu2P8waBpjM0tCDRA/I
3PmDYIgHu1GIpWdqIJ8Vg9cUV6LHb8B4PuCJTf96AHtluoAJ61tvAst+HsrHawey
OEUDMBigmJnNVjmz+w4svtgBeN4T476IKaHpk47sxUgm25M2ZZLAMrjZ8GlMIaVK
yTE5CAB5k0/ntK0ciID6KSDRu+Xc+eO2LybxZKmIfaNNQX0JPOuhitEIyaL0jL2G
/39XmmgfISp04DPPFwYx++/wwlInpjnkoQ7zx5et8vWK4D/YXa7zwWIO8WEPmbVZ
oc/D47F3cmuco/qitfhgQw9yZWCPv1yzwh13P+2ALJwxJw0smhy5qX9tOrkCid6w
GtnjBEweUaabMh8O/0ROaYjGZi01DRCdmWkZ4eJ+zGbTUVf2VLuJmwd/EUgU2UTX
HthyEYt/KzgMCarDE3qRPSzmhtCOSxz1lsUX6Niqm7aqLetLrJAaZwA7A3z1mJyk
zpEiKKbSij2WvGVM8Hf1SLxugDYd9pVsNPiRe13Z+86I/hLN4JzquWfoPUQVhpWw
bgE05atLstyS/cF8STN0UG2lPaExdSQi9TGor8/Zn4o219vUbEIdvceHElMePJMu
OyKchDrooVTH0+wnSSAmO27j6ne8o7G5YOuJidDn1Ne4KHgDRCWorjnyKII+WOvx
nc9z91bc/uF9cxNrU9FqAF6fMOGPpXL+34POTcr1RJDY/WYauQmeEirzSeOVt5ME
TAGzPDox6aL+uDsM97TBUxnTwW1YRnlZYoRJ4DrMvvIe5eA0RUErhd/kVVgdY5Y0
jkoz68J8XaLvGN8pvPnDNGAnezAEGywpwKsutxfKjaPLp1j9QkhG76nkhfAgX7R1
DUhYIjEc+lKSMUPca6GNkKb1EA/KKv1nFIk+CaSsxJHw2S3pF0+76wOEdKuCFdf+
CzlL0P+Z7URrt+4enXAowwi6x3ZYWYoSo3sr4P0HRZkP4UIQp6qeKf8ILHkOMs2v
YijeDkYtQYoInMzIeRDSniZqSiIBkmgFw3Orc3VNPTpMEplHiQGf+q9tiQgrUBTw
6kduUn6wYNkrveigSHT7jmVJeYSPJ//bVGmjDUEPn7mo02gu4IrL0LuXtJWDKBgX
gujSAEkeYMpqHFG1HSt+0z3GLtluX0DPUpTVHiS4GT9UdRJZFloG6Zmfr8ObbOkj
lndN189NFZARw4mEIAysYx5MuZaoseXu0cIOP0EMqX/pNtGB2MmrRQgo0C5lS7XW
nhMqCrdtUqQVlCRDWT9J5ICFszPbjoXmn1jBpgu+kCpotqtA1ZQLsck+agnt2mpK
YCzhU7xCtDnxxHnrPBVTU20dt8ctrzi6ZnRGsouWEb6jUnhiBZzjEa+WLtoSAy5H
G6FRnfTksxy4lPWkc6nSE/eeCntsZeUa1/emrtkN4JTE70+LZVLnE3hOJJZYviQI
vEDtz984rkzcMqNn9vl+4uj214kFjI3lZzLq+GgdI3dg59ppDu+XBF8H2W/biDNm
clNl1M8mhxFoZz6ch17RV3+kVZz2hF2yqiI9pBQ34Y3GDdiE7TrfFPJ+IuSFSi21
qW68UR/EM6xa5ryNVUKxDNapUaV01fBtYzTVizLRok9+9/lt7HzPHQVVjdLrsxpo
3IbbIVbyRq9r+h6Kid70tC9SEnGMszDVgWT6wg52f/5gmE0qmXvMo/khhggBh0Uj
SSzaTQH78vnqefzT5mWCE7JJdtqYeJ2lEqI1ZCvABCWqvsMNBukHIgbc183KQ6xU
Jmvyd3V5Uiul71x6p56ds8ca/+wIBgeyCUZKeY/1X0S4vwzsIIDtvRHusb6YEqQz
kULLgsCFyCVqrJo88/N67xvqLfvMQkRm50Qf0RLKAv9mwYP6vX0+rEf6DocB9GeN
rZWTtOCqdVbuxZhenQSyEVfA76roMjJdD3n/GuOJ6asrznqH0lWzyYn7gVZ32vZJ
6jBhs5sk82XlN41YQUHIOAFUvPCTVjnngqgWM96yHkSWXAxKGn1fPjjWgRRAvkaa
OjcrRB0OMztIsSP/9tOxneCRenrCfgWHupmJlEnGZJiEDt68++xq4QgOIn3d7Ci4
9jSk9ko0yvaBrMkkgTr62qOFVrB2SWKjbIwtX/n2S6U6vOgK5yfAZJjnGkxjMiqR
Bl5Lqz+RbDmzaTiQeD3LeJt41ddX5qJCXMWGlvOJdLIeuirzEMy3mSkuW6vbuNeX
VWjHzihSeL4yr+Jf2LKAMY0rAYN22ETprLGoSxqom+RwrI1+DSGKhLEPGPzOJNjH
LAm6uMIY41K0/qGaIVBCaWvI6aqIcDB08aVhrAWTMlP7gzkaZd8ZKuvPD7JH/Unr
uoX/xHlnXmj4bf6kEmRdUecJpa2yr7VbwaANjWFbQ3BDFxZFSXHhzRzwfVLN12r+
3M6Kb3XDpcwxR4hay5MqBFi+H1eY3C17Bn2UwNc6G3msyROVOtIVUS7i3KxCcDaM
8YEfWi+LWsjSAWX2/0S2i8hue5ZQG53uEXF1dY6zNnshH1l476iiQ/j7ziGPFlsJ
VufKXgkyib7ScYas0095nVRsy1Ww9MmZldcGGJRKPVIh6B9VEHX/89PZXP/uv0Y4
vUracuR4KSi5x8v3sQuhGq4JU2eCTw8EoQUaPxJFevzukofe8jVJ80yQ9vUS4a6j
NN7lUqQGSg57xttI8xHz68aHdwQilQJ2kY3fM8lHCfCK3wIGxpXOHwyC06Evj0U8
TX8tXkIz7RMZk0ZL5B5U896KcRyCFWvuCDYjz8FK49MPK6myfphHRDsoTZDN0rt9
uSJYTTX8V8Hk8TpUs0AYyRdonHCQw81QZ3oeIqDa7i77baUSZitbFnH0Ab0pw4Rb
+HMQBU5hp4GjeY8FCL6KbTmLwjR5hN2hK0KAia8lUIy/vw9BaCy6RzNKIeRXekhL
q+JtQtjOVNrUkpPOt2CiGzt8Yt8CO4i6c1n8uQPMZLz0hPOfq9yW9bMRfvR29Qc4
kp2lKRsCwOKce6K1nY+nlB5Jt0iBVZ4ysRcTK2xFq42dkBeJN3S1sxqqaTcBFFFI
KAMmXHfD2wnDr+NDvCnF5moMul7+oSaBNb0DRNg+f9wVbnJZERh7NTtYSybYgAY6
2W9RVUaCH+Gn9Ume87k4qSaGcKRDlTL5IbXv/5o9Zv7lQ37ZHEVm1cyPL/lRRMnG
mNBmgiccqGe3l9lC0G7tILa67JVt0dJ62WtSRpRw35iBsTnVl273orVlmH+T9Rqf
8hX1PddIqSi6qIFIFZqRdKUToEpeSZ5pG1b9oB19jBWvFk/mD1CZtkUPP5cGakhy
nEdDL5Ra7uOB9f0fBN66/1qXaNXUJ2WBjTOF0MLsojvuVNUm9NDi0wgjbvM5ysvR
lfgincrIXEl2R12gODCWOy3H7SKBIOiTwhjQIT1NoRYGTh0KaW84v1T5v582fUrL
9mm4DamBeQ0l1J4RToXcavt6aBWjN3RwIZU7b/Ru/0YKTKuu621Dhoope7w0iMvF
ARUXtrF5AzteKMQAGW9hVaMwM2hQoeTMFWZtu+hMpvSDgC/06VbD3INUV9I4tO3Z
2vahPYeLxeTe7QT3vhSm0qa7Zz9rcVWivWZKpt0Y9vxZuqB4LG2IWCBOrh26nxeM
e17zWMYQxxH7pwCVgMglbco4yEfxhxU3XpgxPzS1wvZwVY27cSBN7MgJroJCOHmE
pulLlxi4rK7VFPPRbIuGjNn/k2D2YiqrCrn24Ra4kIcEOf813cT586XN4e0t0lls
QqCuLPwyD+dweygS3Dr2Eo4AG2osaW2aXynOM7xk4GSHU61+UMlFheDV7kyc7dOK
1L4UKme2ShlLeB8vMKHjYmx3Rp/PLV5fp6L4jUnNEkFftN2Ri91XqecXz0hFDmOZ
jKxnL3pZDaNMhJACbdm7fBhTMJD/8zJnO2Yc9o8WM4fvFuYgUfOogel3WFoKrHKG
zuFDCPALF2KhtJr/QpT3F3aMumlE9276n4wkUBfP4JKy9gzm3c99pJvpt4oSN+QY
7ByCWXjljLt6+EohL+fgNk0tLi558+UZs9qY/p/ifzUk219yaM8DTSLdRJQyDzMQ
vQlhEbQxPST7x/u4wTHSHVgg00uMTtWZX1IVUFLs8xD7UEbc1pOCNIzSpboS67ZE
3XEiOBTZAPFXcAw8Rki0vxOdGyiPUI7gN7SUC7Cy8Nr7kYuMvGVUWNMDNvaiIKZN
mAXhZdspKO2nyIbkJWSfynTEAbkdoBYgr0ScV1o5kWZV8eWVhT4j4ANr7ysyBDky
HNocmrzVFqkGVw/Ltl/mzdkjHhQHC9fgtm33NDJKV3jfS0gv/zH7rmvSmTJYUhyF
4Xt7dc4+TxHAgh6hsc1+Z8R5GfqqEn5/rWCKul2pUAgXUVG5xNSWzmZh32pyq4na
8zIV4SVusNbd/Chk9OqzYkbstDUL/eNSO6oSkLW4A8KiClCdzDTmVdrIwmM0vj7u
XB5JiWdCzzJHUeePXz0ClpBNCGVdFx7Zskd2jbxTggFsfV1NYQllsZoMWCRYug9+
sAxF+GsvWisuPFCH8GZtOeQxgmcBWCQtOFhmMSkvqk+3pUQyEejbkesw4QO9paTd
DmyXZjM13DxDMIno11HUXZTFPW0lZgPp2VG2nSt+lNC3gjQYIA/hrMSn1TqZGAFR
rlvcfB2jHH+GZg96OxIM9Vhbm+DgqrMyk3u7NToz8Wipkt4FQeewLppvYSXIRkVe
SBp/asak7oDYUj1g3m+sVo94HOkDgtoZ9LZD0hm9n5lL1f1IYwnEqER840RGS338
zEJVQtEYe50wlyzk1r2YN2LN4Q9YX/pWQILCKHU9L1LTNQkS5LHccxXEZTfm66bZ
bFxqJA2jDWkBgLEAM5DMBg7sHewHIudiPHirRHKeF3N7lwJthmBfwnPPzckRRXYp
tQuXzueyacMofTlXr3GC8psUVYdzLaNAs76Mb1cV3iFCXouF0brM6GTg5/ZxO3aP
EwEzMSZuhNxonSkzAtc+JlzkX4YeU6vNr1zzI2WRM93hrvEm2vdhZnYDXpFSRvqH
5zWQtQ/lH23bu9c0ospjTv0Cpkp06VL1K9NDThvKNFAYntQHO87l//+d4j0qtorE
AFnibkVZoHcVSm3BJaLW/eQrl+9WKp2Nt2mYk9KZtNcF/5eHZvehELumylbWdGWZ
jPpjmeokJrAjGhm8rgb6OkZSxvo2vP7A9icbHunyYYrQGpliq/9ImfoGo6y+ulCT
QOLK6vBKlgseIhLIvLW+H6JxKr4mY8NKzty8++B9gTAS3baG6Frl53pJTAdlgCaz
a4DgXhhvb+XpExP9T+8WQbpwvK3nxN3iP12FmJLEFzxhi5ccDy8cc7dE910QbuF/
u6IT66wXHCLkP+FwpBD9IQpzAbxp4kfI8Rt8gRaWamywPQonlMFpSYq8HJn8SSa7
HEc4d1dqqJ8blkGrFKKoxa0f6v6eFcQ4GqRXn1fQ5X1LfrE8SqjxNi2+n+M1p7Hx
QwRtjh2OALbZTkWRar66UkVkXtbZPqTpDVxu6Nr+teg3lhb+mc+MS63T/MLzZsjL
BUbOJ90xc3bE7WQ/A72EPFnyOgGd+ceoqouoUJPvhDjs/lvH40PF+z0mtar5ksRH
qTee0bo5Tst02ej5njYZJU5OhQl3nj0hXrZ9jk3NAoHI7wQh9KGUPxWo+Ba+nYUC
MztJnBQEQ24tAazuAl7GEYdYW79p4dO/E9mA1kEmzhqJdX7Y2OcaFS3lc9Ui7uYF
L8pbdk5t07tGfCU5JGVHFc36oQ3pGjEusVG9J+xbGzqlTI7U/9//duogCWiE0s+p
PhXg+kC0lbg3encY7W0anniv8MJ/Rpfv4pT4rDYqjVmcfB7FSlcHuszJaELkkr/f
BdR0PaPWMdvTxjjBwH1Hbs2cBm6yS61WMOvGku2uo02AwmocZ1yjAIOKuQh9tiAn
1zkhzjSe0FMM5mnLgMbzDFU2ai5TtCIS8IDTHtNZHWtOP3+f6AYhQtLyF0/Zfvjc
Z/67Bkbv8lGA++q5IQfqY2sPyncqJImfqBGNrLjUNAUZnI76m/ztL3s4iCuHk8Mr
hjcwKuSuL3c9dHJ91gLs1uEskimsPuVCZ6exu2wp1kXHz6XjSY6aC8PogK87zuGD
dTRODx8hSTV18m3ZvTXoipdo1/WrPLZf/HuKvrr+rBi0owXhqAp6nyxOrv4xcZ/+
PQTEFFGNZqsp41PTYdvndOGDg6DO1t9gO60vqSO1ykEF984cod2PaZm9ngGZYt7k
fWA0yEcol2LBmvpCDIUrHxd8ZGqDSJNGYAWkLTu0WMrHxdHMmP0g3bhFVJZSyl9D
/VBUDtUnsIYLdaJcvH3Ufyfhj7HpQdEnP91YFZsDFCmAMezDy910HPfM5g+Vq3sZ
rFRRek2LH8JKQGNJCXmgKzd5qT1G+8lp65h9r2VzbrrRbNYo5wPKd1iNcf4V1jSQ
qe9pk3zRFoWhd39FJWQuTh+z32PRspRdPWb7BUEMR9dfgIXXDQYC39Zx53UQICZm
X+QTAfqTDE/+TQCzikTFdSTq+BrQSscVSap28N5jbmMaHVdU3NJmDqllqR5s2+d3
GlpxBsA96ShNMqKZ4jTz/Lc+xZpHpLe83YeE7xGUMrkpC0u63k2Z1uW01NjaLu9C
8IOPLnkiHdvrDTqkTkcTrXhjU7MNajOuKLvgc2sVucoKYpjMaFdaRAYLkw9EvGSt
Cw+hNwik9aXl0+CmOSgh3hTONIhE7kN2EVnBMMSmWF3YhdXpdlO2tvxVidasIggY
t858ixpzz/7yr5XUnzm/FOp+G90inhpb21P7qPH/E/410dNnmt4AdqF5OZyvo9e3
FZUsXY4jdEo0BWP3mp9xpdodt4SIUnuH5VK0CliXvs1nZP7ujstJyiu3SgWeZZ3g
wx4rMAaERGDb/YIVItbvXPBsuasJBlaY0ZYo2R1s7qsauIJ79oIdfq+h04a4I5b/
aUHVWvYyrMblJJaRrUKvITjuP/0kvwYnrU9vtxQKYTf1dR6pa7cRGiNTljkQsIOH
K8BselUx5Doo54wHicO/i+G/tvf2+8ZIGW7F5yLB2ERtQ+yf6mq3HeihlBq5neNi
ObrYgTXZDGxAmUYVfrBJTzRbXTHOit0RxUc2GusSOjVz9VZ3TXVKhndBZMQWTTN0
3J+lBJ/UUrVQm31fGrVSHyCefVqGFSoJXwFV6Z/U4ddB6ukuHgNPdoqZkBHfHVfm
Am8s+V533a2gHLsl5BUPvWFjdClzEkuNsbVcJ+2tyltkB2tdu98NZsPzpljs+Kvh
oo+dyozwU0lhhj5Mn5IB+Acjm0Xg0AA2hXCfAJn6cotN8f1FfQKzh5Xcz+wPNfaO
lELYylc90xf38xKg4xfMBzMJbufG+jW6HByKkSEDaNFyJU3junD1yYFhGZprX8NZ
MfmeHCxk6ef/YTyRTScnvKSRVq8OpfiZ9hJECADJtSMXprLosR5LX/y0fwn/3+0D
40ICAO6DhNu5OvE5ZyOyOv1tucDVsF2ZG8REy8r+/pbo6incahgim77bsZd8OfeA
q23prc7gWeo72LA+pN2+CHvbwQah6d0c24S76ttWBQyn2M0SuRglIucte4EfHsCC
dCByL0cACkV6I5zz6y6XhEwwt43amz0bu4b10kJaDwLk6oKyROgvpVCJ2YDBrnWu
E0Z67zLuEwvTqi0MvH2DI1OF24wmAHVsPEkmxMsH/wXefbbVfwBEYV9MXOIT/Uq/
nNJVb8NKdsLrwGzjYtiVQkKDVKHQCRDWdArnaAPCDuq6C6/9AXLllq4R1HpcYC7o
2d7oOZOyhiMoACLVZeO38nU9YRulk9CPIW+YpEcNS8B4RUWBydbLnGTGB4R9Ff3t
MyLyn0GClaX60chcluUtU+SSNfFTEZZ+UChY+0Z+27hdYTBFKnN3x7djKzBJN4mw
Jpe5SASIPbGWoelspDhidxlP/4UxqB4MZB/1gZxFypXm4N56DvXXkg1AndtOGa9t
TC8Q2JPxvvPXhQvUbblQnMX4gZZq0gkkLKHM73iFL5c+8Cnk7RNDGfSgeGEVycOQ
acj4GIlq7VBJWeOHqWRbsfBGtSYxskinV49RhG1SjasZvfpZ+efPCiwljrdrq7is
AQXBWHiw7vtD4zUO27JDubYEHiCuk3JWysaUtDvt6b97l0tgWy2pNR3H97fTONsy
D/v34VCptqWQagJalgdQ8N9zkD50YKmgM1geLVdjvw4AuM4nilgXlPxC1jcGKh77
+W3c+86y9gy3y9Px6BjI6kZlLaKON8D9jem3iKq1tGILHR8bI1HFp07778Q3OD+C
SEG9JpjwftKGa9nMxNUtcLL08fxE0M8XAaUzUGoXYL4cPDa8V3LuFUGBc/0rUYV1
ZY+ytfD2Lt0ygsIFmSUPalf4FpYagDPcZoXOCQPsEbYFAEEHdYo4Z1nac2n75RxH
VYPaysO1GEkNoBWXg3Dc/JQgnCUEtxUWhoyNofH+JfLVfo4BEQrMAZ6Ledz5IDDy
Ewarcsn8177wc5LISUlhyacaQBc43sIRqqD1W7u5KahOXniBMadIYHEYNeWap3nh
oeAmowfFK4NxKZhS5YtpeSVwiKBE6hcpYyb039UDPJD/haZO+07aLMbqjO4xcTw/
o2AEK89BYL2yHrD3ghkDdDVfFxxN0GYImyQt/JHP6FDvLGNFC7W3v+7RbxirAue3
lioXIOnQo78NQWs8cYHKeg==
`pragma protect end_protected
