// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HClk2xwQGvIdHViH1Z+fk+pbHg4JRCDIuUnn+K6vNiW+jhjahxHKqcTyP2r0Sftb
BPdVsq8pZDSz3HhObYBhvU4xXTWidGH7WyXKB2JnoEsER8Dre1KTxN7mltdGX0uF
ENcioU06Az3zHGQi2l0anlmnTNj65sxnKynWEvBWZ4U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3152)
xqnuBop8Jr3DE/WkZtp+yg1COMyJQTKXZpYcVse5FEdTh0qusrURI5zwbD0mDMCn
Rhf5rFpY0UoNGK1COA7B6TVvhHKO99HbNCjVJSUFUMsczjYLGp7dKNKAlQ650SAQ
SI8Nlm+ZYDuKjg9SoiWPtPMU6E0soGkZxr9iLHZoxbj0jSuxigVQe/yfaMck90PS
XzwiW2W6xVc8gqVZDd/89Y3TJm5UHS1EkMDSefJA37ikn3DMtif763epDUTNGA+C
UIcJy+KUk6IERDz4gBDqBREkoTXz2jDol0gYpg624QuQULDg2SABK+cDqNHyViBH
Gba9VP5GFFFE7nwpOv1Sn05qLb1ztE5SH/MX1iknbeHjH+1n2sm5eBG/8Z99+1BA
Lwfso1ZgUSa+DyLojwDphSOMEFAQhu0dsH+XqtK2iDGsLnzYqOMQ78jOgGqC4Xft
fZObMktE45/TyhWwGX0sLCR6wpPUQS/YGOuOnCJhRE0opA41t+VuOT7Jo3xzyQFk
UACUxGETHZwHSQFBZYlR0pxoSJaFW/3LG8IAzBzjAVW58bnunSs7kn9izuwnOXMy
9PgxaONXI/Evfnr0sSJ+VtXO3Mbs5W73/rOy5ZIVO3+0iFaLJX2BrvLmNzfuV36T
Ar3zXr04M66YNyl68PPdRKSjyM6B8uHF1i7THXLfv5gAxSC+ZWBNUr2Og/7JdAmQ
u/biF+Cqi0NLL719fEiN5gOYw4NbWfs+jwKdWUtIhfDIMPKrqB32SVysKBuhpfql
ztpzQioRLgVkj1LGXT1yA/saBSfMr60NFmwKZd7INKe/hOLoPT/PPuHFgKgjrIvz
Pfc9moJD5zOyB5dTvsh4lN8sbzFlyE/Qye/RCV3u/ddB+rpY7J+sTk4kvgcEKppt
QzF8gMtOssFNu27nd8JZif5uYM7NeDuJRKK0gvsQChKrC57Ubnfcu0pvlDuk4Rf0
c/txNoJFVY3JhyO8krkxWiOJMKRYgKxa8ltndiF8I+1eKZpakHcOFV90JV66xRcy
2F2XY4sCc6mu4zbxGZZ/lvCeWhLKcHyqJVM2daci9Or1Utqa8Ni3/jwoIX/Ut2Cm
FY6omey685k10MQVwm+O/ewQItQN7SnbVKb19EepPpPIluc/GD2kMxS/qqGVLf3j
NU10FvuXrRQ+0HrTUTgX46EihslTVsd1SWWdDKNiCqT/VoUV6RS4j2nqOUCXay6X
5oW4Fnup+p4Pp8hOfoFGyHdaB89kqeX27mD01OIkkS67fhNFiP2T5WCAOdlyd+Ty
LZMOCqJHfiodIr+feESwwGKSrHYOKDi0jqQV3PPtCXjii+5tupePtG8zI8ZfvA8B
iOxZeyAyaaf7ZBZRofV8tAWCbbpkl5p0++m3ON3zcIzUlIkUWOpBZFtZKmfdy01n
PepbtB+NL8oLBAOHn+BEqm/m7u3lCSFt7SvfRYv7FyOyYcPknx0S2GueItB3nwuo
QfdGdcfwRu9I1EWQsKY6/oAcloZmRjAxHkRQLqLWVhMkRrhJ14G8nXCl2seo0db8
o0e7HJXIwgBG9nvIsPn2rByiHRHBlJVOrUk2Szwd/tYKcikQrEM0L+BehnLkI8Cm
BdC5GRGXC+1+EYXplQIr7h1LKrUxJrfk5ycL9JjREpbAp69lfhPh0I2X/puuUuZy
IG38lDjklQokJq+1hcB8m7nVZmHJqEGAlAybXfynSwzfRQIL8APRSQfWSZD5IdRM
o8dDMkvT4vBRFjFToxvHvp+ipkZHhvbA0JiSd/YlFwrXpiMLv3ZCkeydWEJGusP4
XjsY0KzMOjBP2PwEwMrtkcgtOROlK+BzCzTetqhDrrF8v9SNriGDlyEsK5S9/ra4
GUJfRTEI4f1+bQxam8qvLCfJsBRzldo2i0BYyA3P5wCIue1++pMAMLR43BP28v/K
4SG/4toZcZwJCNcbQPZ9GdcKxhCaT5TMab8kipZ49JVKRAPrjDc37qP+lVV2e+2s
0CHvOwsqG6KmlnDizgZ6J3WXjLf/t6JHJPiuTKJvFoOcJLy6gYkTTiNyyBAW4WCZ
1ma72/z3DKJU7PV2f6sVDcGPokUypk1RZL656Eu4BEaA02ZPyslYiTMjdhOHjUUE
sfXRRHPsm+X2w6pBYsIDF0l1LWhczJ0eBObcdXnxAQGwwC4IGltY5kRT4TI7A4FU
gfm/dkUpKM7h5QYfoiowQ+XlgnbUScHoemj9A1t9UOYd5BKI64zZzUos10/TPGKd
LXpP/ejfBeqmHCwREwN/xnHbPF5yRjdW5iat+eOG7SYekX2RAyYxgZM7Qlf4vFX0
GRV2OBzNkX6TyaJOYwhiW5/n7BIvw7f54habF0N23TBLyaPa0/CdVQKyQxzPYK6I
QqzsmMyFc97vgKIFZ7Nz0o51UgTAZgz+8k1BZ81LdUNA5md9UVF0ipxncB++CrvF
mmCR46xNLemk5/HfzAXsj3zr3hGfvacKPdvbw27qtqvN9G5LLK9Ftihh6eYu2msl
sHEANWLZSj0Yyymyt2ESlqwiSEVoWm5fUNriMt1UedY9tXNUMLr8CMmPS+WUmWP/
vOYrKZ6jf/toRSf+m9IGEQBiMPlJBCXtW4t2KIobRJlpAWWsKpjJ2y/8Tkv1koao
xBt3WLMJ7fWDZhtI6pbTGXH0lPB1DsMBVUkXC06NLGRhgbPZe9xmkCWztUGilPel
GLOhLA+ePLGklikfh4KMCM2KTnRStFGjHxZLZe2HeICik1jDGJZZEsReCXUfkd54
GuNviB3e6L71WwA72Q8pNLMR/FbvF9wjcV4RzvrVNGiWp+xFfLb80AwLblEc4Fee
lPJXxYqW3Yl6TAPplrC78r3UKln6HgAfWB8vke7KBRJ2sboXW3NLkhcYKT3KScq5
mxinW1bBgoSfA2YXwgpwlLrmiejcR+RrcVjK02oIml+VJ/DaIHX6vpxBax4GirCC
Jm0AgjgLH10nBiMHtOuEgpA8MUX9mwC1o3fJhwtrr8l7cAllfyX6wkuAws1oAf9k
V9T4R6oHECNayNa2Xu+Tjj8xKompOdp+dXkIskjcCYyOVWcO1L9Wk4cWlorNkqE8
DRARNe/lpFmQJcF0/qldz+xP18X1VzsnvFcqGpY5aHw3/sbbZKvXD/R2gG819b/b
0v9zyd+LZOXLv5VQbK33MaTx5b2XjVGFVZLkzBhe1PROKZPQgD5qfUvnXrLvDdwo
dwH8HnxxwepaE4eJcPOzv5Wo6cDH/lmlR+LR0EkWbUAlXOA/tq661EFJDGkl1k3p
Dl406UfKbNncBKSEBNQ4oAHykb6CanYpT2Fo4DmDGpSj6smq4UJFG+WYd2VjAxyH
puxyhIQ3Cu+3MdgsA6XrXnMg0WxSVA5WdG5smr3wFZDzJcLnk3MLqEKJcgYiZVSa
xFgaQ/ukyVBCjGG5iIqSn7i9KI1/Cke6UAlHl/+f7SLWk3C5PW11i4Prwb8q3xfC
Iiv9JcclqfhG5NZsPWjLxNDFRvgl8OeyV1luyIDYcncgY0SKhIFFyleYmWe+XmXH
TZHeBzlArycaa0BxEP+hIrcGjkSNohgpjhg6Q48fQHF+Mxpe4zZQRz5gRRoI35Qc
hkyrAhQtLyfzc6/BnOAS3a2Yxe+cIy7/n9ygJanjosKdEoaNRr4zcKmfLuCjIxDI
+UHVe59104m3shRP7WzOeGG9GaGx/XKcQ6LcdMdBct1UQ2MjVo469DokUAorYEJb
F+m6wZNje/tm9azmSNQeaK2tcOWfD6zIBf+6/PUJgXi5jUQ/wyK8uIW72gRZGe38
lVbKTCdC3fs43mP4+CA6gkrJxpRAj68aSkPp36Z+QsnNlXJ1yPyY8wSB5ZZvznhk
o+wwdb5IkdcML3B9WOMX0Yxj5bZVbNPi3ybhzAsxT8BAbS9bd3fYdvqdelxB2B/r
+K7DnOCMqW6x46IG52cTxCpHBwAp6rsCyC4OdB2QeMxxFa7LS/VT+A+f6lgErYas
Cg+mgzmAqQ0dAYDerNCkGIY1z/JkXikaZ2f0PBdmND51RC0KdV8n2OiOzYuY/Y3T
SH18Oxx7+8sW5pZe88/HBqGXFBWj52kelLBM4P6/XVsj68Ei2vPVWwVuyFRNS39u
ekEncwZzkMQIuA6p539V1IlUTrA3GgJxJdOS1cd1apACHR7xkawN6r8GECSodkbQ
+N8Fo+kY/CZ9PTrgs15hl1jz2i49fsI2LNuOGD61NJ4=
`pragma protect end_protected
