// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hLgjJw5FVYfsDQ0G1Jk+JYp3JeWPIG9jPKPwW5cUTXMqpI9qt0F1ZQ/ImbeXYrjk
iweR/T0gF0M9G0CkjPRAcqUAAeryOmJvaRppzLOvHr45VRGmErkzrKbOIbahVoKQ
XBdM59c+S/vkIAfmImp3Z8EiIQJ/L0FdB+ZL22zaUt4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6608)
AYARP/QYuFa3l0xfv7+BMUmGMy9d95RJHzdiiX8ExZoi3BY4WcwZh7ikMHhR3GOF
UeN9v5rJgsC2o88+PF1l+2didQRX2kwkulDoNbzDSOEKYsN5+hAd8/pAm0SJpKCh
305OGmY8dkPrFMoI68625/wX8UvBPsk/ghxsoBzerwSB3cOAVLeLZ0ONOz7ylCWQ
e3BF+NNmEqhyi3CdBaofEGeLdbG7kd2T2l+r3+msTABFJkor4b5wXo3Zx/LttSGE
IrZAP5DxKhqS/bAAg5RHhBZvCRk0OGirhYvnRE+XIDKQqcSrm5Zwx9ngmLD+GiPp
7f8SYy4otqF1/gc46ksfprAWGB8U95gM8R7VhCdTIs9/SZ7m00HPJYMOgPFQyybZ
GRj4l8RcvWBrJU30xSHBtoDd2dXgXUZMn8/jhF6/R0D8T2ktnHsBvXSE1N6CCCWD
TRX4p32Ft795vjNPc7gN7/3hNrytZX7B1E/h5xh1zOlVJKjFcgTWe/guagQGHG3L
k320IVAKf5JVIBweFcK2h63XL3c2MfcRKARyqX5j25Ppxx6NBUJctXKmIZZFDpoO
f6XqyjVcQz+TvOeP+KbaI6SDaWdWaIo9CaYpDyWgJ1+Rdhh8LJn3cld8h5kIj8eq
DpdimZPWfL5ib2r38u7WBzI/VRphts/SWuxqnAOnt7XghGgCJXKAyjgx0OCMjDbo
2F+AKv0Mqg8FARh7MHsd3cQfpAKf+lDfVwXb77IOPz6ieUZzAMepsaSx1+JtJA+u
gAy6BBj3YFFCyLxE27ivTd5kJUa/xZGLqzoS1TSNgOdFE7LYEueCyhYUw4AKaEVH
uLEgZAqEI/jToPCT5Z3TE2RVbgrokMlTjKcaGTbdr0Re9eYuY2EN+2akwb760NqM
VGu3TJHe3MSuud74yxCPjtC9LFGWCIjJJrHmb7pUp1s0o+DTRxDKqvjyvMa19k2h
n9zcvKChZcxgiHigLpNAQN1aSFW+MHnZlUJ1HSwU4ZidcwOzb3g6rjgvks8122yz
pw1wTf+IQjSrtIAZWMBVPYij9zkMi/fjdVjfSvxyhuq+vrVHTO796ZxNPg6QOYGI
5+FTwPkn8xY9p/pDFoA0NeYUZN4/X1rqWxfKqmtyWgQ+k9idKZZTHeTKyBbXCiFs
Xl6i3fs0MoN2LvHfJ+DI9XmBrafHCWTKAmeGmztuadOr1r5jx7fkzXmWJEtTvub6
0NY1k+NlFpx+t9/qo6kOOAH9nPX65efzPh70ebgdThivoYA8jf9aauuY/Wq8dzEW
5qBpwBFd6E0Xx4jdx2og+UfzvX6BqjYViJLHNHW5sGos2I4N6FSQ+b5deDVHaDLy
vBMTjAvp0fzf8Te3Qe7I72TUaDayRXR8K0ojyj/uFUOzhw1RXgkKQpyeknwBPeaP
Uv90jPu83oEaDGg6b50n0aAf/4hRyJs9YeXr5IocGjZcZkKKRJVKoYi2Db6Y4gDA
ZeX4y2GYqWs0quvojWQARvk8d+Xa6DgeOYsInf0f/ROZ721GkFVOeb480VhOWyWV
17yuvSe0F1PLJh3Rmu0HIkuqSouoRTuQ1uFIQ9fN5TWYIZqYpfDyWdT+SHuGzJ3n
pUFpNu5dEifeupQDZjxDjx+0BxaMRo3UKNtPG9n4xQkCo5MwxfgjXV1ndq8ij0Vn
WfUt94Pw7tTluK0MhG1VHdjay2H6cwjt5AxGwnKxaJvf4lLfOgOksbr6vr2cyv3U
+IYW1Pxp5e+mm7fwf16nfl5DywDY4z/EtMsZ/lkzbKR+orPd/OyfbpTN+4DHqmwQ
nRWnf/AvZI9xqOb4ZMgyvMfhK0+kM0Ko5wgZxAUobv9SVrqWwOPBskkzoTOgA0Ny
BJFFVtRoaKRNIjgBWWYWBK9X+w97ujzh60KLu5ju6GAlxXK9/H3CbxzbWJDMC4OR
uqgHBkcnXMZyF4Eds+9+GbFpx2NGPVDDfv3m6HJ8Vkteg3JDRjtyk+Qp3S7lG1gW
HkQejMxqp0X71uQ4nZlhoaJuaGcxqp728nJfhxcDpxc6CMrj4BXMlcB6PlvwsDxT
R6rWLXxZ8V+5dboW8929txdxCOx8ua8Ki2b1X6QWKO+hnwxwe2+Ao4zIso0oSgSd
od42g+f8xrVNwRGeV0k5i5uMxVceUgzZ16seCOLswDyswI4VjIfYnB08TIY/06P8
O3LD9r//OQBjSbaGUmFobxcz9YXX3oenxWwfwF4k5Da26HC7MoqL9EKj//60tKUc
u/NsckjHAYCnO6FlR6ipD6XRZYzcCTo0oZrsbna7oweC0FqnUkLYp5O7gTNIJOe3
6gRgWMuTrUKsPH67PynSuxXHcPsMHPkYaWdJPQUJ49IP5mQmU6d91a/AcZnlF/Sg
oglsiN/L3jnh0xcWM2D+ng49CNkN/xYpICej00un8MfreMCedZaRLehuJoT/ppFi
uxVmPJ6l4o7fXfE4eMRMkY7vyME+kx1G95rrSl6/xUaj5zmAdrdvJS0SHZl6aBNN
0DGnc2XutRACt2uBRYhtaOwdeo1koUNDuLSMM95pAMMgzdCk/8ckGTSIsiLrbdEv
/xMWrVwhVxMct8qRUxKgEEr3EBnfHffy/gQr6/aa8Cta5MXJSb5zojZr4HGHNrMi
KleTf50BqwxcmdIOtZND4zFtxM40o0SUJudeFzGuKflLauGsk25QDut1y7ntovOt
VV0qNlytYYBiFLKmQVJlWXWZYKEcrl2NzWRALAEaoDjR0/zwpaR353Oe5r1Hsp0Z
efV05lQaIJwdQu+eyu/OIklppSA41rlmOrWY9JakZXTRk9pOtzHjChYHnXvSA7vx
qFkZeQdwecl1J6Ove6W+E78s1ssNXq4zTYtYLdmZCXnEYsUdKiqknlaty2I7TUqi
WXrEevdl6z5b4aou/4YHWj2eB7L+SLmCh3Ni8FCLQsCI5fx3MWi5flDmPDFiyNGF
cNnTyGKzVLzWTZuiusKeRHBwTuPiKUA/BEQoZ6nhhi9JkXgQgkyNuZ96UL1JrGK4
VYcaPE752xiL6aES5jn0DCLu1CyFHFHLTd+HJXpr3zIHOY7mFWcZD/Hc57m4Vzrk
/BBy9qQuANcY3yF9PqeG/qnbsa5YvVKv5DCT7RVq5TdDQeqQDaLNoDxdsg9wmVhM
NOVqtz87IKUucASWS+PDwzYhzPRoFbVIalmR3UuHIwcpKf6CYDvD5Y36qVh+ZwFa
18edNkgk3LNHL9WQ+PepOTP491KzD6D+mVcGHmLN0SZLVVyQIQUE4P27tJ7MmQ+u
itYzGxCTqRGopiMrSuWNJwp3zuL6FoVlDnLPD9NRg8rG3jCkaUFXdlzZHztqlAkh
G55X4k4p37sF8wMy7g215I4eOVxzxL+K3hupeo76MOP+y7bmRrbGzTi060f9VKlL
/iy0I3mUxdut99ME/UPawTX5OqoXzysyPCHCcSdgc0lpQtj507zuZPSDSdZgGiGt
d3/TrVVLWNtZyVj+8CLYMYAGV4PBv0E2YP2kvu5jIeQkSeQuGhGEUeH8yxZlXSqk
BX4F4ZjiW1y0dqGDtjMnMdMAxvZzYjWetfBzvsSOf35bsT2aVrV95fARCl/PVtNh
atT7Z6YfXxU64+OGcDY34ncrfEVaa3vx1asP65GEqwD1tWw6HXKvWhpJ3PZvi+9C
0LnVt490yrXB7BcBWrgGFepghq6xZJ5gnipkIoJJtSsZdVP3xtm8ZFgDaxXwQA05
RUFygw0u1BWVR9b+eUOcfRReZXs7UExJonn5vPYyn0qGjhvx9Veuv8dGAAmwCdhx
rHOtGs0/3VNAurQOSiTT9t5w+h3TwvmA06uWgunbvnzrijB4xEXj6GdxN3VuWyqm
nGP9pIMMvotoXAdfbjqaumJ6eQClt1LrtBNV8XcX9WvgoGvw826EZRd9jiKCG9ur
yt4nd3Ba4Pxw+UbKtskkmLWdePuGrzLjqwNnh90i3lBrlU1hicM3TDP3Gy8WUwaN
tNAIRu8w24Dn1pbF8B5Fadg77XGiWCK7+JlLbo5zx7irAoe1ablCOuZoY+y05Rf+
0JnDLokalQhk0y62bxSGdy+lepczUvX/+K9CS6YP3IZ4Se9yvkyaFhm9L9SM/xa/
lymXLDvrwmyaEPOY3327b6lVDIGTU9naVIfVreP3LDH6xcOfmui+pAEmKEourLiV
PH/MDTQl+J28sIFplcNLmayY/k04AE0gzvrjSaZB43e1Uurn7N9UMOWH4HbEYTuf
9CJhH1D2aHqbLXdJvb7oEHhcWH5yO3a+FG2BwO3DiPxrB8yMyoqRP4gYUel2jHrc
WaDox1WQlrlPtX0xZCFCRInalrUbPlNlSvGpjaqWkjAgpc2COJRe307S+YGz5D1h
lpXzbC4kRdGOZpHHcQGTVnSNaX3v8OtTF/rhvdsUwbYdrq+9E77ESB87x8KXRdp6
AgPYHvts/p32EzPBEiJr4TTqLnt2/xxw240oQTpaalymDZBsd5ET0bx4Quw6TBfV
g2awUmvjs9lHmhamD0a9ruNTrninplHMCAr/v+n2KaQgYKvebpwrW4f9rRADd4rv
3OmpSn5azBWibhUud6CbpYoeNv53BKIJIvB0yGVAHDoHEKGf8HI7DqcRXBkEf3eG
LTCy4Fr8CnYe+mGHYd1Ib8jKXsQ/5lxmofKLBHoUVxpIAFgOFwPpmLwTxH8vRg+U
VqKuLPkem22BI/H/J3QuQimwIjvVveJ23yPpZnyP5EzVSnNPGJ5wRr0QW0V9pD2/
dwmoZgTVOlLOvVmewoSuWbPTYdQyDkQti1lpRPgbOtMAFa+5CInvVSvP1v9IOg7c
J/tWVEPeV5uWe0bzTSUtr3V0PDh1svJYFAaFEkQ/JYx23sXuwFfcRzOMCSYQafKa
UleS4RI7n9xkxmdTXAdAXIVEicgdAJMBxY0JooWiemMtvwAh262ybfAOy/SCVKj9
OQOfQpGouYbjTgxoWeHd448Sy0SVOcaKk1DxO0AbJlS6eg0M7tKh8GuRpOukgaxl
+V7YX2dHm6m64zju/BDS/X40I/ctdu2DrQTx/pHGSkqtYlEpiUU/bwX5kW8/M3TF
RtHs6s5cBXzwUjsihfdR+APjglcqVyKMuhKpkr7ewT5SY1QC+IBZmuzApb3ymjmv
mMFgVV35emfSdzjTT7sRR2dW5R9LHnEwaiFPSXMVXWat5/XEsSIYzsYGxGGO8vWT
Uxm3PJOONAGctWLajfNnGhJbWFjdKo4+iw+APBal8W+C+aptdWSDebleb9nIRjnM
UFf+ELCRqNK+66Aj9PEyLCRHAaBAnixKRwOPANkntRYgoBF4JDxm7gSOegaCwMbr
eN8YIQCyrBdo9mUAsMDCyqZQrNUQ/+z19EKvEJjZHm6k0aOOTpkem7vIgpbw2VWg
uaSL28+RaNywOH/M0hO9LYvv9c7YHoGjky8B5Xta2QSdLBsEsUGLAST46ejOCHj4
/Sq+pTXD7RqFtuajhkU+fzgI2+HvMZA1s5zHBrjEBimp0s8Zj330JlZR7aI7uNjP
nuFhy+VDnrgi9SpkVhtBpxDrIKpHSB8aWIfc3dIQiEgVsNPGvzSCeN0slDb2KK/v
QD1P5MF6WHI6JM5YmaJqym03LpdpYjxXh4YwvUEvo+qv94FBAgVQdFcVGsNmv+oR
MuCWEtNcAxjDQhSeuCT4rT04u3o7zUzMCfqWwvA5zri/BMS43ugSvISix24zmdzG
0E8p3i7vuwkLp2X3+gYxb+gZSz4tQPHhD5234S83XXmduRxZ+x5RPHr5vfKLh4SH
xJjAfuRfDdXqtp2fgIwBq7DY3LHEWQ5/Q74fBeDWW6FQFv5qkw/4ZgAjGF4wRqjs
Vo+t4APQsrQjXxX1oO0nv8sedu+ZEtfhBsRdg0e0tIXyErHDUq5B2XHOYkar7Vho
CEh4bieC1k4GxkLW29vQAqh5fevnK0GpT/shMTzVBl51P80UIax66xO3dkHphoAC
rSzrYB6oi/jiY+cMjyWCEPIUVWO+PcuFMpPi5wFDs7/AXFqpMxk4GrjMDK3B4hg8
+3M8n4xgiEvsvsVjYS+WsvRI+GvvRH020EMXr+cx2ImnftXV2mKmdeBeIQCKp/zP
eHqLokjuRY483f1B9PZTxKRfsHnl2SnLyFAhcBpe1OgLdsG0VZ8r3vO8hJKdz8cc
f2ma4ymBYq/UF7fJZl2uPFUclJp3Ba88tscb9xobDteVMaf2PLq1e8PDGtlZDayT
Fv9yhTaeVdzBeOz5lF0Hg+753mDNSEX7mO7hOCdFwB3oixl/wtMhhUWVt9ix2u/u
hIgLfolqJx8XHJW4h/meJv0c6XYMwxsWZS8ZskSA0FjCd8rV/HCgkhbOqH/BwkGi
KlxWjLUJ82kCHR61YlUjngm3qP5LnPgYqmQJQfb79PsxTheYG3XHvfXhfRmvbOnJ
7AqnT+dHw2Yb2IQoW/T2QISzj/0gNRij2Ic1aRMJCN3WpuoXx/EusqolBXryq4AR
2CPHdwyp2fEE9vkDVh7oIISwFbkcTAzSJPQwoCAh8sMM93LO5hzOdVcXGZq6LGFP
u2AK6VByE9qHtYzV3aWWk/vQ1fE7Dw1SV+dagfFK5Yl0W8Jrtxqf4iROGsRV0hkm
/zJ4cevFkPbHKJDbsk67JPcf4lBSnUEyRFqO9HsrbvSNrf/zNbGgh/sZpQ4rSLG8
LfKRG3CAOR996G68rvQXyawoWmFwViJUonl0O7et5d3SYxsMLhl0knt1slTqsczs
M/V+N9YgnVIazRiF1RSEsXwCxoDhKDs6tYGEzOr61uWKUTqLNQorAx1lxvV9Bc48
8E1mEeBmeAUoRCGRk4F2p2cuh8qIBVKRzhqKiDffQKhVqQ7ICS8eAe8xZD88RVKL
eVywG+/wurtF97oy9371WXzfdjlYndE3vLlca72vXL7s9/RcRmXr8T9835MetzJI
SceTLLjWRpAcZwKg+ewg19L0tLFRnCYiRPJMGcWQbvxTWEhTAFgB+RZuaeZs8oMv
XZpMCMrGOspQ2WU36cyzSLKbDF0ARUCMPqoKZRAdyTKn1fqaW4OCWl1T6gBsHZNO
b3PsEa2DP7jyhJkdaXgrOGvYyf8cRWG+nAY8UfWQP0ANnOKenTCCmcUvfb0IkfUo
d6S+KR7kC7QgsumUvhHuP3aeCVppvVQsNqwm7OeWgAmpGOLsLuCfDWWdkPAZKw5I
u6fymcywiFnMNYBs7iIQe2tFAM3KQEn1fpMEkucF33+GPmN5sjAYnlaLvsgfrv7H
odgG3M17HoJR+P9NkFpVavegtDBXB+tbljfncV30vAxoIhZDZL1635iGvBr3M7SS
HUo+FSis40WYjef3HJdMEqDbLPEDT7m+9ZfLPAFgLabaPrf8soQBPQT3J+dwvLNE
xfJXXNYYfL7cyXCH7txHrqa2cEzFIi+vxDtjaqXpUX1zJHVTqc6yeJFSrZjV49KX
n7RuYZIyYWAvH6DS6rZq7emI6WHfsjQU+tGem1PZr6dbweTw/ddk50mONj4uTrvv
TiROELZUqqT0qhvcP4pFyVGt4qLPzyRYLJ9Xqgtb8p73/1o/2D7P1rUZDo9lWstu
rFQfJ6ZEffw7Pxy4g4Ou3AEWZW2FJhYG6ycSHUBDeOYzbhVSL8VcdKSi+6iS1tVC
Ghxrf1gRB04/n1aHsxkV8tTl4g48UGr1mrjHRyyeuOYCVWAeCthH/G/l7Qzmzm8Q
FojyKOm4lOhCwOdvHwlasT0jjruyv1ajzzunOIsdJa7BlY+fzoQBFfcg9uF3UF33
44DNczYX72poePqfXk0yJhXET3/7wUjVoYby2mfynYwyxsWijFn8/34j6aEnf5xs
njQTLHJwj0KWC7me98KAQ9mvPsisY0uUOS8wWXtqCV5P6NO7ZwprHVUL+SFAYNuo
N8JgGfryWKl86hPtEdnC1eFUB4U9b6Lv5Pi4GIlHq2Mr2dDopVw2uxidtOCmscq9
ZfLlJTrqAdhHF/W0Xxq6K2L0FVgcexgwIXla5DjNWpf1SKTlQvg/C1d1ALGh6HON
e0umq7UupbMU/IoJxGgKjdnLgC5pYkkWx2cKh1BBaMb7RKoQgQcHTDx8g67ThakS
caIop8a9lOAWU+jLWch+KDq2AOprJ1m+RTxCu7EKx3lOND9j6PKDauMDzrC5ry+7
R0oWMXM2oalwuzod0THTgZcyBJBJgCrnnhvtHSovH8Twa2hGsHw0sF5yGmvAcU0m
qQwJpBG+A7Ym2z8ZkZSd5ckg42ovwtcFyAZIC5kjSan6p2daPJuIeKhKcd6SPSlj
wEHOgSUbSzLa5wvfecGsFgBh4KQ5ZH6QNvJcC0XP5BRfEXJqN64R+Vfyhod1gXPn
S/DTjmRIiL+pq+MG8uchhsVQ586MMQuOK8nAqd1p0EW2EDqb1HXM6jU0qIkeoM0t
x/UX+QEVOM/RsejeaQlBrbfjzpu+yg1yr5RNdX1eInbAnV8llqu/ltFyqjXxpkqQ
zliTueTIwVflVlKjdY4WK9bgHh5X31tTVZANxzgELN3vBCiAG8H2F+PW3yaxw/JB
s/tYc96Wb3oKHtJNv30H+8n3kkcOnb8wvuaDPH2UzyY8oFhXioJoUnXMYEYPL61D
tXGntiS853FKdv4Fr17J/KI5AhKemiBG9PpaBjyJM/rZl/tgeD3XvLDArsSfA6An
Xd5A7fASFZD6kmOIw12O0mVcsPHOXnVJ+ZlByN2JSorVBi9gH4ZuXsAhQSwIOEnj
8MEzflhd5evazlkr3A/Y++OB7tfbHBG38fTorLmqOoXBCEF+b736fkyTjAf1xI3v
4gzjg8Qiqt4RgxWFqJNejV2VPLURf14RGOf2PpWDQbk=
`pragma protect end_protected
