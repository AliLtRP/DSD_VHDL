// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
eg5eS2LPIJW+xkELJb1RdYlILjle3ur36H7gInYY/4ilZsuJUgtV8YbVmyc3EZgPfIg59NAMzpuT
Kv2AwEdhar7ubfNBidrV6E4iONsCLX/MF8fy3PvxhilVs97Ii4d3sF3ggbvaWO/OBj+7TSs/+F+F
pGgHAsPUtPhnVe1arXVcG38WLecaxrbBRvF/7hvdkwJ2qhh0SN76/l9M0MTXyfhnsuYI/Q+cUI8e
cG8FAnm90kaBIvRR1N/DKYuoHftD8VppRnFLjVnwXuvilUWoSvGC9Na2t3PM8+uo/FYrtMdSlpbA
5NctEAK+Ls5ziYCJKfj8JBT4wQD/1ci/a6CwRw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
DKT7OAlsqlHwQJRGoG390V6QmzBMm+6xTLxC59bRua6YnIg+/yEY1IrjRgCkW9PbziSP/b62U8vt
d7VhjHiuVHWOWKu0XXr7KtUtAFJeCcv8v8ER4QlMbiEsfazUjlHOGZHb8UdgMQWZ3bvrMwxait4t
UarSl5TzEjsHbeRyG8Vpc3yqtDohoN6artjeXQQo7V0b20cRKwHKAtOE5Ifq/yEpdpcvngtBAeHo
o5LBaetRRA1l29tTeycS/Al/KnrgHFrhEFMRt+SiEUGhyQL3dHymmRPUp6anP2YB6W/6boz1vU+y
3wq1pnZnHnvlG4rH6VabRbqHMBFARDBta14O3UmkDHrU1MUdw9KU0ltUAgOx4w+u+jwdxj5KJRwg
p2A2v37GLSCmvfYowgWesd+HPJ83/wEqXkxB+5HU/UN+ogU13FBLenT1pmgu5xUUm8haIwq9tRv3
VA50VL7cF3mhNhmTL+pTKYEt3npuFAEdnAY0VS4b7JkiHfN0PMbWvcHugXVNtfyvkk766TcjPbcs
fdVD0O+5Y9ncTw0yHwEdY4jCFAxmyDPtDDVH/w1vHB0HjLmNvVM78h4k2QiwtAMCtGyHwGrZzJ9E
siXtNzwH/CRGpD6mCGEwUwKqAfUbmL0veXG5lTVfcnwalifiGa5mQve/WfyS/mrOOMrHjFO8Bzmd
GYcu1Z5TodIdI1G2EusA6qRpqwv9VikG5BxRjXcvSU4qBEmi94jbqZfbmr28hCh93yfUpl4kApYo
Nt09zfADBgFF3Fj1YGjZ4X6aIvuK5a2AlFzayioQP+p96l+yHj5t6vBembDcp3hXxM+TUjB5r/Tu
3AHTi+l9DDW/JxbF0t7d1glVQNMdRvqnzQrseHugH3YU5Of/g+vxr0N/8URwmPoF7eK/a6NIQiwb
ZlMuh5rd1y1zJqM8ICGiRsdSD8p37kLLVIi8dT1Ud1oLK5af73/xqlnAZ22pCwGrupG3Aedafnw4
os+GXCSbY7bWWNBmF1Q4D1u/b2B/SH0JDo5kHXsgC+htGRVa/IwmVyeJemlwGQvaPh7+dT7QUyTo
v8/dIznlLUkigv90GllWTq38+04mU+vq0bQA5++FQHboGM63ozvdQFmwq6P7/xxSd0XAgDr5ZuXE
zCkmWyEejzWeGCrHM0syVotcDvZWwZK/CXXR8keM3b0mO3mNdlau+qyfyu7GhZ5W533uQw7FHsbu
bcHU6eoH3Ps8i9MNMWNKhwcT1B+dcXRGUQQWPPokLP8iIi0hn0tO9pmEwA6K+UmAOWFdg/cpZt15
hrQgVmdZtixG+nPC0e8JoQfvRb/0AomdQeObWAg9QIK1sJ5P1gjcL2O1EvIPaXsamG716cyq5Bgp
+LdOizJDIRO2DpYPBoE1YV8M4cZr1l0A1/YNX00iOBwqXEM3tg2Y73apZIF5BNjGPZconvnUSOvH
SG9Ef+EKDDN6UmZ4QkTJoAYIwwKrr66pBYQiBXwe06VVjUCpiNsDg5tM9F01W2wkiN79tkBf2q5D
7OnVldnK1nMdUL8FsmG+VbP/7/rjswk5r8nponfTjXcptyMo8OF15MzW/fm7CCJLEtg0gET/UTL0
kKS6UoCAa4H19yeXvewgTVMstBSTUdfj/NEWxhJVKSt/+M+1hjAFsFT8FlsDuiTdyw7LU+egUgfm
z22eK2oEIVMrjT2EIg0bYxsWwAbsVtVH5dBr/7YdycimeZxdPXEP++YKy82udhc6S7EHXLTVuzvu
AqfJLTP+XD50+gUtypkumoupd6tygKs+9Lr/X4DT7smo06eSjuAJ72YhCKO0d5GpubCloU3WdNZP
LO52GelprFEDmK319QxWeI7q1qq0troxbClnvENwv+aw25TEQZyK7nhZ4mmFhp2loGXhiSL+SKBA
KpEQwteB/OXcdL+XvupRbPkHKHxKzQrarXHfVyQNk8ZRLhD9AfehGzbjVcdD9tk2EOR5aATz5xR7
1AMSQD0WUih9+ohlCBdc2a+7hHOQDwGotwF6Bd/ptn8N9+ltwi8uL/jLV6xB9Kj9H9ClXCrEq/Gu
GSC5L0AozUp4j4F31M9MFH5S3TfUiS6c2+gvaifZWQbWZa6L5VIFLpvoJUfmGjbaJafvcF+MVnel
dukKkUGG8HgiK+3KYYYyC3Eh9xqDL38grSIE64EIStIUPnjZzDEezCUQMZuhtCNVgHUW/q2SUxKh
uLw2w1v9z9mPTSLMi4JaRlzbdbSWlQ7r/f/qEvfLEdGv7z9BKW6jl76nsMqI4vgvhSn57HcH0CHL
UIZqNU753tOBsZan+I82s8pz8QxDaY4vmU4pc9tWTto5aBZ431hkszklmHspNWIASYoau/n6Bmub
yfD3t/rqWF1q3mrlM53+Qz3PJxw3/x4OvBx0jCpNBljQxtXHHt0haQGu6n49k2/AV//fm2ACWyST
dMuAHQ1CnqwXz581KlKrKH2aFAO4WYZCQrTEycJ8AGzWiyTVt29hF7BL1Tmh2DlX4DvBhJr5YffS
a2QcYUDdiJRzFyiSUHE+ITLdxiNkn3X5XTr+UOfky9H2FRJC7X3onlXxZAlWcOkb78mZO7mYPXFu
2oAEWKH+0zFqrC1YioQLIP+qw4N356I6zRGp23LDt+eTKguQ5wfZ9aihDCC32OoCONDGgzCZXfuL
QlLFtIsRLQC9Pd+R2czYmT6P2Eu6wpmGaAen+UY7wDjFIaLrYQtorETdnSZ5LZLzDAAg2gCXel8m
9rs6ws+JFS66Q5tzgkF6odYUiRQ8WqiX2mq/UPQG8gdn9HKpEmEcOPdPIdQC97Y4Ym3zRAfqvXMU
JTlfLwGyYv/Wkz9DHG2lLFng443PuX1VkHTxZNtVPOP0Emia0fHHf1ixBpZojm+V+Nc0FNkuOu4+
KCJMekaL2GO/obXBO4M4YGjbSXtp0D5y+qFngXpdh+eOAwgJMZiHFu0aJq46+Lf8evlTFGz0045Q
LgdtpAMrihRFPv2h9/n/a+E2HLeSdH9zQttaYjWvIxXyF2xAHgBu3RG0XSM7UAXV65obdHSyj3J0
gsJZXjWPa9xBsYvP/OQE3YzHYrrn+MeeLPCUvzTECooymW+IkDgvMJvtHx6dzuJEkv97lVKNEDIW
ZuDC4XOy7WQws/5iAKOs/hO7m0fDJw4lQPVx/kxS8sW9ECSIoS9SB4MrlFHLufKofysdmw0si6V3
bbQ9t0N5mGaNcWCaEZ62YOwKLCqGZ+yTbLr8wofAzGPmUyRJWfvChFjbb/QzY65R2j/yZSzYTJBG
47PykuD/q5Y7UUP6KFJ6ZuLmLkyAfvHOxgKemb304bplmYsX66NbWIBg6F75oXHH/bUkGfjExkAm
euVZDxVGyhzpqmxSbN4aAXXbxI9fjnRqTveoK6g5wP+yxTl9LrgdGhj4FWmOn10ljN6aPkUbQIbX
F6Od/N4lOZWoGSbMpRiY0fjdZe+6HlHX1uyLN397+jg0oGOcNEr/Vg1p1eaK2yI68qDIUiV7/jft
+nsR3Cv/e6vYypfkftDeVCbT/atXqpz/lWUT3HbRHIva4HiUHHwyAOq11531dsN8xgk8gBUZeEq+
fTp/au0wom0dBoBNnvI1T48avZIILwJbH1sLzMG7Wj+DKiM2Xd5c8XUc+jfEXfO1xmNxboJfCdQ4
5ULll1lfCkkOGfwkK2+v0KbkkKkQoF4Wzrjz6NLYu2uroF1zMHrH1iofrldEKXzy+jIAV0/3hb/0
50CxICID9JdM7WsSdAq7ppBq2iF6/muAlGTFTu4kS4XnbsYoSbyrXC1bmOnfxU5e+ZwHWulXUN6V
pIOaTwyXbNBBGVCk1mXp/GjoQjI+yzVfi6Gv/MZuHnp9Z0FFWSJnYjFofVWV5wEupcSXOCP/23Yh
Lp6VhMgonZjtwP5Dt5napBx+vhgAkIj6rGln3i3XiybBKAgGeZc4mfgMwwmq020CMv45bnALIiXc
Eu5ONCc3Raa7OSAp453kGPGhkkKYq7MA+zqfpVfsAO+DZGEYqDE7Tunws68+IC4lOhVg5Y64tCN5
pG7mXepWAp8WkneojsuYTDeWyBKcuq8uEGi+FhgihDze5c9JlnpcXLmqOriPZpcWjuyzo+8KP3Xg
GU/iDkN56z2akPIsRmo4w+Kpgqn6hGe90FXc+kTDvSBiaU+m/MvfFtIE+PeBiB/oGYdEXrirhNzw
cLuJcLGh5v77LY3p7NGGZikfJ96aLBQ1yFtipiJLcn6G28bWFV3iN4378Xv9avbQtOcc34sLsjyZ
WVI2RINP5GJMqMOpG5FWHT+4gyVG8/fJ9dtfJihod9SSSbiDcQXTLwdIYuatt/248Evz6rpuAkWk
K93svbFB9cpOYm+qdfOIv6hjjFHLLXwrgTBTaMweTgdh3MXYRiesmtTpv7f2JNCks9HoPTR7Ldw0
4vfTrX3nquk0h+aFZn22dDMalCUWPHKbklLIVvhKzmqfbN1aGo0vtnmH+JUoxeylgvT5w4bpoRN1
Up1M4CQBr/0ku0OriakhxtOoOT2q7QB0aAxOtof1hegD/dx9+Uuqf6un9fBOJBgCXkqHYM7tZdkQ
XQpvinS47KQ4TW15+ZseNxufcOYkgaXbK9fuOGd8xJtuoGJEIa89RdTUmRE5jXm94Wyb/lHxXGpd
rFL+OmOB+7fMy6GzbSjKwWJo9Rf1RY4whyRnqx8COje+mYnU8ZNqDeBXP2Yfufhxx/JAqX8+8PG8
cB8zbLGfBzZziH/7xfCYftar9BebY3+hP8qb1XwRtct9Th0/euDvORVkJQ7eu6f22gBQS7yApO9f
zsGyWL+WYeKMvCN0B4CHcyhcTYurr/09S/ZwOzW0BaeIyDUAJ8JkAzwbzZJdWjeSpbwe4ewbeZsF
KnYG/T5ERM1GApm3IEJNcSffN1DYqpcpuDjD8jckGf5oflIPadnJYO1MgUslinqZKjVNbrDHAeb3
Bj5P/kefilZsvSDx1FmyeD/JRdSNbuUWXOZv0kyUYsORuou2ffbrVkO5vPfUyLLQsN+vxv4tDF15
teDZAtNHy+8wlcDXe0zZrBDD0V5XHOfgsqslwzBdSF+rp1UHu4uG7buQIK5y1J3ABbh/u1CJL8Fl
XhhshIfy0kKSgisfVHjVeglffzpz8yoCK9q0wy/1P1CBmJC/UXOXNd8lTkBeUdxHjcWsKiUx7T/L
3L1FB6bJ1cEAi7K4ztEJR2KFY2QNkrG+hkuDx9PlfN8QdA4oIGoKo31YKhSpKyiEvpPhXrp3KD63
SJe2lNSSzq1So9v1WRXLsm9CHMZkllTsRX6RW89DatAWmoOSOKEPgKAGtzYf/Vs5SnvsGOP4HQhz
qyDu3H2dQDBTy1daw5qZVym9PfKp4o7we742oDnBs+mM9d9MQ52w4EIT+FmPmIB+YJq9YbTN2aMw
SCyE+ywCv42+cc3sjxVgUb77eu2/4mxXMi1jwoJuR3uvnKE3RT2LInrV1k5cBxkCG9eQLy4rbrby
lsYFbfliYyJxRQ0bJVG62PkRizSwXbDZCt3D23NvVQ50bSmyNkzm5uL/o92QYQ3j1QROMdHCqQd/
4crTNeJN9Sden+bT8FD59uEUOLn5X0eIMSMnPbHzgI3hEnt3ErAFo4YgTRJ+PH8A9PDKID509QwE
4UurP8tjU8bJWxwhlP0gtq+BTe7exQ+Ext9Av67iJWtmHslLIVvlgy8Jk2uFqvBxD5YvsTPh0vyB
t363zj7FBZNf8fzny8wVcPKoyljOIGvJYamkeTsehvM7tiJZug433zIJnTZJ1IpNE1PamEJ73pgL
3JY4kUvTrByluT/BgVfCQHX2ExrhnO1zwWLiXb7yuQjh+1MmU3SQx9KAj7u+I4aq+1OQyvlWlXv6
hxvfWnAIvHd0koopJ3nocIfVaZ4Q2dl9+5VG0gsbfJdbESKL9yZsiEBaHhwJa1CEqHfijhNPcZxL
VQmE22nJzw06KBPn+VzD9h4sMic13qwhISaknm+sFIDoKjOQV3l2BmNoYlbCFuUG55t0QQrt+I7R
KcfJgI+ss8a9O8saeS5g6mj+J2pq+VYPGe2/W/iN++AptZjjJhuBFpVKLMs3ynzKUY4HLJt2ojhA
zlxk5JgGPnL2icSEpxthehla/jOohvLzAFAMaQJaEefHgPxxCUWh8gaJ0EEHY4Hjr8IZVE03eK/w
XE2M7cx/+QMnOnUvJV3ratXDnt3YEAlpgHwHvBfRvx4qfzjVaAsBF7UNkEqEsuLfT8gLa/a47hqM
NrLAnRZqb+jy186sWnu+aEhFY+FOoZtJE0sLbAYfqMOWTIkEHWRe1ry454/WmhPnBwii9UJZHU/G
5EzGOM+rNE/JJGQ4kya5zHtNfRuCvc347Qpk44M68bbGBwMXrp8EtOXSQLSUzjiqjeVLL83qkfJO
mTWv9FnwqkAKVmfqQyO2XpGp5SZ3z7acwJfLyzLic+rdumdfIzZQfAsCFe3pzfTLVEua3+8AFsBN
RyYK7ddu9oyQb3V/N0GCgvoZjsYQNbJMGLJMU9+dgAPPv+pFLcJ4kG3nAnF7cMww0PaZGO47PVa+
OM8e43tviQmLvCiGRNu9wjTnmVgjf/QftDXrSWyB2sSy/I7RwaxBi52S0eNpzqrDaX9EPJRkfe/h
Dnf/jn5TN74XWq7G+OxwppIkVLqeFYQwaEkKRzleHJVoD0ky37LR11FJa8vtCWXOpgUNQupG+ZB8
lua6ONoeKTVqnJPI3DGFQbGhceMXy3xtlfO02G2YARqwz9h+j8SWc82JQahsIqQPbMz05Z9Nn4es
6dTP3CAbbuhXDFT6E30ZegGRMw7xCtTI6RFNIM1VGlogwDBeCQFaS4bVGyI/Rhm3BD7/zUz/OPf4
yw1oevACwHTJphtnY/s4zfPMYhPhFYDUIY7Bsiv9SyJgtaalOLuTpTOdIZzaNwpBFtofaBG39+G1
JGJIz1Id+7f+oncykUI4fpqcL466ypgmM4/aZ9GuWc8h4DyvFKufRkBU6Ngf1n03dLDpWwfre4HN
9R2OCAJXB8VckprBv/asEuUCP8jpByjLocQfY2BoruB9xx1RYOAMniN2ZOvhkEndwkcUDxK91ri4
WTGSFSgcz1orlKqlq5Ms5dfP/FkNwYhi1DTkDHdhmGA94egncxxcOK76NxnEbfYuYeYGEwZs1rPx
fyPiYZ9d8nLhxTzw8CmofbxYoG3ZtMrlL673CTKbFKHNqoH5f7Mcjys1Tbjb1pThllepZWHzkxma
iraSyuMaRV38+lL7+B/soaYNnDavNHfKgiLBC3FYZd8jq7PHY0BEDe8/2/qLr/YPQLHj4NjmSgxi
+9ZwiJ6EliNPNwlH65H9fzEZterl+3SkLlXTSgeWMLtWiNYyqB+r4P35zpcyqgPFcBnYRovz/Sd+
+C3vLxXNyrlSP6aNwf8CBqHWRPfGSvwFv+yeL5rYhp8EFy4JZEyPXOXvmhD+PYBIg2B7kVdOfAll
DCc28V/oEMjzxsYjYvbO/sNkPHBbnVLfXTAbCDJXoBl3CeE5HT1STF+wxUwQ9gjWN/wRXJnyyLlq
qDrU/qlYJR70aoyTxkQa2hTNu/yjoSZAbmUb1p4uzNWEjY88+zd+r9wdJEjAvXBM7f7fTn3SFnVe
NA47sWhJVT2sHlWTkWA83M3JkRVw+PNP40T4wzf8TxlyAIrJgT1jbwBp0ImAuD1KQYyJBCJUEvve
TkEGtAXF1WwTW8vtFz7Qfl1WGNQSBXRwKibyq/5LCAyNC6/A/EMFlq84rhz35+q1+90QwAtHil0M
YSzGcdGpaH+c+2duV//AxEwgAs3aV2A4jV78eunqNbxPzlu54qQ2yR8X61tmAW3iBHD7z8VBINcv
4EuXhsRlMYi8RZo4dL9pB3N4BgGscJMzrWnVUFB0JA8ykUhSheWPEI1oh7O7h37Hr9PlHPhngQei
T0KxrRSSMBQ7HlJRPzwV1o/CJIriixfczxVVu7aMuHo0D0sm+INMZF3mAj/xuzmeSonuI93/YSnA
4Ux8tCd4Wmx/kyMC9aeL5Y0XPoMkzVISST6uXBFpYPEHDpmMdnqfKC7OjrzPeKRf8/zWejHU+Z5g
+lqNgw4auBGT1hEIW12W08QybQL7Ii3E7fgllGdNDJzI5WsPw59T9z1w4Yq2DeAFg0RZXhwc/Som
gQFzCe6UJaDlOPq4jquuFXRuAx19d+MMLl/QMSWXTlfU0crR+cvRphT1UMkizCOELnEoCn0PRdfT
WsvBGICJ4YByYc+p86DWLjAg3r4r4+KsnSh/HJsD3Bisr9oFiOeIEhm0x3fPCKdOYiI2phky4KNm
+bKaa6C7Vqgd51jcEedekZmlQD+bDhV3AG0+Vq16yrfiASzxygk0QFL6DA/4lUbM9Nfkp5S69SYg
oEnrAxR2bRFTy8THZBsFZ4+CZ16jgUZ9aD9+nojwTov/Dyv+lvGE2OLu+zAQ+vbn9uZG5NBLpR3f
xEcveEAihRt4WdNfM0KQoH5adI2o8ANEuE5+sDglhHLMj4BnQdwAkQexi6YADjjpGwNtt1IOEJ/1
1pMcr00RjjV0IqbfltYWqQ8/n6l5FZ19/CSRpnSL4M2O+YgVKdFSESIBMJh0GqFiUrGwTkwWe2T8
vaba2y2PAeeA3RA+R3RNmdd/KX161iqiUGmABtOmGyNLV8x36RY6si/hRnOEgGdI4uTFeJWFR15z
du1kyR0RRW89atUlzKqMPrG40Gp6Hl6Yy+F7b5S/N9Y8A2o/wEoyY75Xf3R98KEkL4eCS9RXlOvc
0DNLS0pSSyzmPMRz/K1xUn0/fsI0YkjBqHlJeumL1gKFUpCw8VyxqZmCxmdRqbXUjUVfSw0+W/Ns
cIlgY5n/9+8D9HbE1IqoTnFIDP64AoSEXSt0SqBJ+/EB9QsLu8FNXi8DDYPRLdtpkWmZGk6eWyyw
xHGOInEISMkalfwKu/B2PaDcS8O2sK7xm0jpmfzUji/keS0nMtd6xizKt/+EXFIecxCrChpUrZmY
8VRSmptz6T4HK6n1k8Zh7XKJ0MblqgLeZHxAoAYVxwA0owPMJ3QPrlUdKpg+uvmTmF06jwmvFo2D
VInECGXFahxIBM7FhumKZYOoCTFf4QTaWU/u6ARl8Rm6L85eexAJXxqWmFZ79q5DLZFNt2hm6S4Z
CpKvCCAbQcFvLHH8aDuWcK+STr7J6PpYE+qTsm4qZ2y6yELz8960bTA1lQD5tZYGvW/kON6qL1VE
GpocAGnzFguVaoarOcVJzKg6FJKn8518WLOYAdSpynj8bIoGjrsFQd9t8ORrlS5ri5zck7AKgi1b
zwPOcGGu52bhMceg9UTsQsLGdL0t22+PAYV5G+QvpRYDR3aXCNd12kAt3b4WtXpJDKhPrWQE7RcB
4TbCVvCv3KO3YhuwhldNfYNUuMR4UFi3yuD+fas3go66qPcs3lHCYc+S7zGSaLbbGtlN33hfHGn9
3Trp/yTpVXU7S3vuoxDBBwCxuLbgdAk+DiPoNLu18AXde+oMXS7sH84JmCSbLqkUQBZWTVZBIZ+G
qACrZFIu2xuXy4xFPvf3pdoDJ4eVDuA3/upKRKgGjLsIUx9a6/TvVwl9UM1puxT6KvooEk+Ylotg
5Byq4xJsPXyI/UFrdnPEVc7uN6y8m5tyYqiNgEqXLJmrNOxwm7stnxg725n0ggfF538akbUR0+w6
5DXlAG5RCtiplCl7stEz3kYHxXWr/XEoZmmaVi+KfsA+76JghsmlKw533BhU4wGQ/7cZY3XYECFQ
GpF1kntYQ+9lt58yMIw6GVjph6yHT/9iXxoEHOY96VPuLaNjiqggXsQU/Iuzq1sQgRO8CGJaxQk7
IJmaCy4gYmpMr5UbGy5xHO+zmBHePeXQvXUoHk1Dd2vmamGDdT0ebbdCeTioB4AvYAW7BzCl7Z6X
i4Pt4kyKLWb1abKAofAtojO+vbbbh3b7es2cihA3Fy+ZZ54LMHLW7knFROYABQJCcc0Isv3NABzg
e6YFIcKhpjukB8ByJj0pQUSapPG6vxydLc9HdIHesTpWiWmfj97SDwvFA+rQZfYlExk/BYK+Alm2
Zqm5dX0T8qIn6KV2g6myHK11+E/2hOj8dlnLiAnVaPpdI3uZ7DgG+WkRbDerT0YfmcbQL1ffAuMf
QVXXO+rI7sbHCC4lofvGcI/hZqyQMyPvVUr2w6GrkmY4yAMWQCRium5CBBpRSE+At1teHjc2iL86
sAb5yhy/rVcdzEQnIKZvlOpj2+GDaC/rOk5EwQuKk6avytlVIaXtrUukGCmE65Itpd57cEC8Dhv3
1dyoevrOF/XWUM4fwFvvCBq+MG0OvqAlmelvRJAFFpS7z10eIrjOcJdMo76a5KkXumuv3FRltxzn
dhuEjcsye/uS+2TIB6c4rWDFZvoihiXEoZg9ICehyPMFGO6JenU7xlW3zq2U0/SRmPCojagivJSb
uSE/ANX8oUGBf8Z48NLIagjSQjqf/WsyeYpfVDaMhrzCSL26zqaQ7jZjByRO+n53vYbioLjWu3+I
ZYzhi5nJFJTt75VLewRf0LFJYSwk66JfStahgYgb/TvETne2WdCDXZtgZdo8CL+RfstCsjeCTaSF
fIawyDhyycsYFonVenvGY/bJYFhHcpk2R1kVjObANL60vSB5FG0n+78Gxxa5DI5s7y/MrxHDD6s2
b6q7hfwlOmsyGDv04EaP7BKmSSgY8S548nuI4bHJeFDxui3r8I61ACwsPtUttsTS5zsWLWN2mckz
r4IAywvyDh0tGlSu9KFrKEsYUC3G3lbpJxZy52NNRjZxzbTCb3wkEoAk3s6V7XZDcAc/hnqtAoR5
2bghD2gwxXvH6ae8yp7w0tFxFPRfFbwLsh0twMlqPPJGgzyVLzNHrp+iogvyS5t8dpXG88+2fpm2
vPG9VYeXIwjZu6jgg/+C/7XNRTR85xTgTg8y2WGNGfQhVzU8/75wogkfvB23uwgkNTuMB0EQM0NY
1JRG+fSmNE7fL3GjmxZFJmXBHp2Eq3GTjF2QT9k9Nn0Rg5jvvYB1IxHoHnM0s0ahxMnaEWXcW070
4Kh+WHo9D9XhxbqRXykD9OuhWnVB6tJipJaVxVYKzIuncjIs3bZ9Fud+tbsit/yk/IUCKj5MFwSk
Lq5SgOR8gDigFPaeGIX1wKPio4mhLOj36yRlHu0NMGF0Nix5aUCyq8J1w8qQuViCd7t3nuPDzv2c
6F2P3Ws/qnUcC9lL27q9QetuXZ6U39OXryAhXzEk96jsdi6kqMn5JImZalAeE5giEBFSxa6Ctrjv
gN87SvfEhtqXg3YI91Yn/8GTfZGG1TIFshE0OBhYDf88jSGQyCFYnYBngFdA4tDt6C8cZ4xWd9Bn
a6djr/3aXw2l4XHKud0KXQ9ZWdJVBvKhBbMM+sVL7ncwkhuqfAIeMwDp1buw7bloO1e7s/AXKFx+
/0QIsroaKK2ff5RHcUqxGbBJy0tpBSyIX1ZuRuP+jYoKXDX/cH45WN3Ev0TJp/L2ZTT9S9ETe9pS
7LPF2llQO1PEsBpf+oT2q5vvcUeF8nbO32098x2fyLvlCGpKK80nI/lEO34+qSQp7q1VZHLRTmG4
nbdaMaZqGA7a+2WFVLdSiNuVUJ8qz83NCQSI9AItY7pQmAfztxC2zQKipxAUuQMBbd7G4NX9qFD4
M8xgklL1yizxk0DCd9sJugLYm1GeST+LHrPOYLbcpk9+h4F6lH0ebpjs6uZMXQtyrtUb94vpU0c3
ocRcB5wesrcLZ5yRY7G10kSz7PxcF6bYvhuCXI+iTt2xegfJxUQ3rZ2jhhLPlTO4l2Tc+4oHoHn+
QXQg/fBI2qjXHqJe4jOMwLzXfFVwW6XdqYxZJ+qqkiyB0tf8ZCUItdZ2U1IefguUb7tiVcjDeyrk
dOBrXHAc4FfHfZnVuqpJKEkgPiY+usdPSwzJv00o3akPTNy7fCVNJ/dKvIfzlsmGoFZLytOe5Z4p
vAp2LfslDOz7ltgN4Vol+EO+KgWgNPAuSLLdu/sLbL3Nzi1vsl4UjE2dvEbIgVluXUW4bhuBmtRr
EssfDrA4/qF6p0MlSiOm4PlnZfrOJkwdUwl3DaKvA11EjsC1h2siWAFDvOFWRH5Br3TjeG3+4Lm1
pf/1HgkOfjf367mnGumbuqxv1fhGnUXYphjvrdAdzGpVhkrSpR74zKBKmtKLO41MCFKYH7JeGpsK
/XY6U/GRiMABMs1wSjHGDUFmatcrq50zzE++83httVugEh09/SWErQa9cSkoS8v0plVGB8nzh2BA
veHyOVlVvDeb8yK27Mk13pKTDw7y1YuT6z8poMBpHkmROtx364WxH8zM/ocpLZK7EqfypzZzV/WJ
ayEIZkKt6vrrPa1AMiCuI6nxxLkgA1nm8yKEH/f2B17fwMHd5vqVvFphiJwqQOkvv76tMWaFbj42
4/foQB7iVnb6KRqGhnvP3BQIwNXIPJczDjXWAj8G/kYSP3a3o4mx2BH5NCHexLXu7i7eybwEV+GN
EOs45OJpfGOaKdVDr5VOx3xxcfeik0yrC9uonlXKSEo0A03i4B5jvjHKoM0NeAmGQfiprCFxwzbL
s4Vkgxucuvh0n0WOFHEo7e/aRKtf7pQsCbQrs/Tqu0NlDzrUHKuy+5ivUBDPvHnMLdzw1iraKLBw
x+U13jsSVyMnt4CosGZnaIN+HwUiB0TBlYD4Z7urrf+6BOVBOvgGR29GtuYKkip+4O7BF2/Ut7Cd
rvqNrg8k/1YuMehHZqh3yDtrEtMZ/VNMz/a+Ecxi+sWXP4sqq/yU7UEiUmRERK2QCuIeSmylVp/a
abo/0xp+WAkY1WVPwZfFStBQPj5NlfepiWs2WkAmvFECa6CAakcTQx+w4EpbYYCNPLy2nyCKc/Mc
jQQUVCIqQUHu6xaI0Lmk2JGWag6ugriDY9hWl4K+AH3PuU+Lq8rDvJU8ms0I2ymgTIS2Rj1TqxFH
Jyne6fOJm5gSS0qIf23wCopYplArLDGd+xJS4iVaOcQND1MmE0z25bhPK+FtQtdiLpLN7fGWOzer
yh6/AEzi6dAhvx3wthd1KZedi/589UEQ8biugcCcrJcAMigp2nYvjQ98fvoxV0hIt6tR09x5cpuB
GidgSkOHqOgPI7YIhSbyf4iPLbSXFxROM4G0PJqWDqmFbD85asl1EsgdJ0VORMOc64aYig+2E+y+
BFlcyNm2K1VQzDKQhdq/UAdCBIVkRrzv88LzQGq7sJz2TwELvcjF0GPmG9/NyXJRSrz674D3Sb1W
pZjZgmIoP+QVsSTTHQoMpiiB+yeUEKdl6smAe9QCFFVucU6v/azYwqHHfnB4dI5soryDoJiTGPlN
THwCYltkOwx2sYeNEuiJHFfCTAs4kdKoeb4pYGiAeJO0S8DdeWm21oUaDGVJGNGqU9iaM1198e9u
2W+qvOHqNVYGB7UB44nvZMbHPEY0uz+mW4MJGSW3wsoaw/YAfmuJYIC4oavUMZZYTtkVlvP5h1Mp
tl9KyIJH1POokVxfCexC+CFMI7wm/2uu54LnB72pav66Ounpecyi3Uj/m45fryriVyuBlOV1j2Zd
2ETfG3iNxxYBUr8pgGo3y3LZcXGKCiOKFVgOaAntBUj1StUDoBhpqn1lgAO+UBLLuaEd+IvoUTA3
9/luQKOALqrmRvu0KoAtw4tqhiztFVo6GHr6pWWPd+geMs1yze5YIKv8mXP7fSwb2Dr5jHLQgnFq
crdTVPIKI+76LWLqONdrRqwvfcZHCe+Q4b2pI1x1mQnZUA+IA7ywGt5lUHcq/KWlFyGZkARTGLPH
EjDHNoy0aTg2n6N9PTQ8yH2WCxBaS13EhPbkvLUUQ/nkPfE40MSo+ZUTaguR+d0se73E2hrc7xAH
ZlIZn/hzfFqTCbB/QaXL/17IlyRB3UE3VLQxn8/y3ciBEyxq/IApeOKMZVCDmRzIL4FI+9Ydccht
SBEbFxT+65Zyr2auh00yIZrRFlCkavBGP+bXvzrZAeQC45u5Hfi6D0JttdnkS0YxsPyFYdYndsVs
RlbykN83/dbsPpdFGTXvtcZhOrfhAJbqLa6KRpMw43zwrDg0keQBasD+wlJYQfk7FavWpO9TPUhw
lFctfP+608DdGD5uQsoyqKjRd5FegjIVWoXi8oMi+XNgxlJEwrLvezVYORyv8jefKKJDNoluomsh
aql17f80H/AEHiI6mYgoAv4FXKJ5/fVUQrOfox/I+cKK69DDzscYU0/nqX2zwKhTfm40w6JEhkCj
6NF7NAZk37ZAM93ttt2gJilHav+L6qwL6Kzr3cLBHdGNkuF5apUuyrRG7xvyJ4jafM2PNysGHY8F
7oGLYbB6Rqksec0nvLVgxpG9/w2lzA9zrXAfEaO9hAslAG+q7lm1J6ndPZny43n5Y6mm4e8Lyz3/
K753t7EAzu8ihZ/us8TW/NFO1OiW4QmMoJnfTt1X7AZqiJ2qTksdHDwwDxGG+9D+8osSv/ZwIxTm
wiliEXd8jj3PaDjWvargYvItLJiJMIessjd768S+ViWZBq3NmEoIPCM7fprqAjG1hWxx05rJFowg
y10iEw626f8RFNCB1Lth2qv3cDzzkRTnrL4LtPRoG3E0RL8Swe2YawMzsaeo5rhoupEqEIuZIMgC
BMEMDoBwkvPoSGtpz8SruU0FHtPXQDA+OGKZ9ctQA/jtDQytz39B25uI/0llm1wj08dMbrQFUzYv
y/Zq9fNINBm1Y4m/4gRB48ks6QTggRNxHtOKvPdk+p/rPhxeNsL6EhNA+bR8C2r6xAm8qTtus9P9
kFu+DdYWKVOfyAFbpCCzvCDmqJX2G8vOOt0KB7UUPnJrd6FAhlPj/uncPwgz+2HXSKqMgL7TI9vM
REhKoYOp8xIqPpGm7YqbnmIB1IpXy4RsgB4H6uEOb3X0C+zszFBDPxm+6W35+5tGI5fnYftxwJ46
mZTyGHqxLKNfraGgBWaNCtHy5VHJaZHnzYd/JcNLDQicdIPSjh7vG9WwMppPYujmL/yzMNT1SmLG
1jwjQje320rSbLSiOFSwb3KU8MSdZIE2s5ihEYhpbHsZqb7WXe0iB+zAVQEMr6PgNEEIu5qoqkJa
3nq6JnfF7Js2oiBSg20Ajtwi/6MqQJ+EE+Qm8r0x6/yKeVDq+Qli/WZXcX8LdnDMkPFC72FTDMNi
M+TZq3EEEYSTdQqHghnqZtXuz79kHUhp0lrMYeSN91F72hAl3HMPiMZfW7T24EjuEe77P/fxCSLy
L3esz/Hymtp+P8L/0dWNzDIbnK0+3MnVzAx3zsYjZJf2a8gx3H+U4zoryDQTado+h8gAIHj59l9a
XM2uXxREdjNvr+wfIUG6LFFlD8ysDvAMDwx7gW1xmCzamEtxp768YFfy9mkBr48nFnKNcCbsSwWC
nqoJHvcVHaoa7A4KUStZsLr3cVKfBorjYLzsuz+eoZTxdA7fcvErYIuC/bBJ01YeSaqJ7YFJ5UIj
qrb5nKBcYU4YMbitANvWm+F8DdktdyT6TEtrD7SMXUlQiJf+/HGcv0yY73F8cOUdvG0nPV10yr5Q
LAJXELXsx4EH8qRLRjYI2vBIztV0IH0GKxKbKjkoxGFAPuI3pWmGF6MxtwGex6I3rf6IbGCMKKQL
T94fQyI57nlT5rsBlBpOp9m/QWqsz8krWHI6WFmR9BfysdnNnOWLj4k0X987xrcAw11t5Y+0xsKQ
lCsLmRVBeAm76sBiqswAV5i7w/yrwSErhe4BEmkNFxoUGK+s/LqkzFrSep4rmmnlHgfkXlYAsrNu
vftZ3d7Xs146WJAFQLACZW6yftsQ1QIp1p13zQMg6L8QV2ucw0jcTIpo4bWDafp/zLk0hGjwiKx9
j7hdsUGJIVy+ieeg+OIxwhEfYe59n9ZxPBUXtPmhKAIde9dVBsVgif/Q+OapFuJ52v8v21FApPcU
sAoOS7GpMYHRUGdwdsReBZAdcvGelL0NEuh/CwkAgf3vm4pmuLA4k+Tdo0rI4S4zJN2lC2O6lNES
4T7jjfD9+C0SkhkcG40NHZtTqXfg+e6v2KTFzPUNXT4zzCJfUMf0ev5E02piZj/DNmZamf8+8DFi
QYb/C/zfqYjwyfDjH95IOhEJr4SF2JUgbU+U5NmYCIlMLD2fy9f9zeaSX5JLxv159MVqEy6W8+QS
3YCuZYsi08a+ijFWmDLXq12otnqCbB19e1vySjfkZoJmjx2sZFyD27LwD2nzVm2Wbtgp9xF1KHGG
qRsZzvhB1/fc09V6xZKSBCTjN68k5cnEazspdl0bntH4NXn0DyejQPpiYFLVA2JdD/KoKCW4maoO
ZxVgJyIgSNO0TSJOceWbAr2rJylUkp+Ng3a8BeMlEWx584dwvdplMkv76JsudU1EaL89rzszAvjn
N9jn6VoGPfa8tylmkg/QTpnC1b83BmUuVaswXHeWfNMq1HSAX9JuNuQO2tBWHz/93zzjrqcF8oFo
89jzFFF3D2+cYBhZoCtp2yuzpH+pjPTRRp/otruV67ZzTjSoQieIcncDrDEamd209YLOoJhkZuc1
YS8ly8aSDspKy++v7yrToSG5ZBMRNciyagpaxQYYe7cK8q54p8HLxx1lKkQVknPwN44k4qlcFH8Q
vRksSMg4gQqz17GSE1JLSqJMiMYFZ4YRSDEyA0ppsgKB7vH3xcTJ27C8a74wput1z8qaggCYM7tn
dqyrLBNMialF9qubeDvyv/koK0uXu1tCTQVoTkgswAXcfzvakcY+2l8l4Nmt6ZuQHAZTYd8/7gAA
LirHJmRpYzkiNOQ4uVIJWb/En+b3ihgQ2kE4vgdFcWV1yZVLviUAVsy0JxXwrQaR2h405+cR7SLK
/Hu1dBVlkc+JWV7Gjo4432YTiJmboZhfRbhUTmP9b9fWHoJ5QuEkskt0IofSLQAbVnEe+wsk0wsE
LAPD1gMYPmQ5dv+dCvHdvWTKks+AeIGKQmHfQTTkV/sQr+lVALXMUa5LiVJBFrNNuuQ8QSdzG/ZL
ZaVcM27NOTvNqvhqOTzWUaGGrQJ8GhjWfKl0DktkLepGUb0eQXLtR8nQLlqO7QLwG58cUsNvj23F
m2WwVL3Bs+s56w24OgL5CeG5DEHxPrptPt17xnGYm/EuXQ5p5BnKUd7JFQc9ze9xoPNzvfgcmrkX
IjCOH2eCJBvo3+aBfwdRYzDG7LjM7y2qwp9XBJ4eFUMuFUPbbGTXmFfVImUzxFozzQy8i0OeEDGf
M30ubiPrGz6isSpSlzrpSPpIUhgXVH1bBH6lbe3+rEUEE7wuiitK/QKG0NjoXDnwotiPVbctSHLL
kdBremJACkzZQGEjnxPRPscOj6ju5R4kZ1sDtpeUPe5qOUmnQiMzFY8LrSXkhCiVWTvC3L7reC2f
256DV/TaKoI3NN05u0TMqtJ8kaVYCdHr9oM0pcGvk/e/P3ymvNwBvCBsknNBesgfhGeEF0hW2TqQ
8mQB+d6n3+RJLQcbJZmxuP4Gnw/5tr1gaZripINmB/cxCViWRMVL99SddsgqomMSTvn+lVXtiskF
9H7PzAd4XMlOPPBvlgCOR+AwKZtcyoHsRkB8iHZ9QZV7gigJVbvq+N2Y6dWudddCDHzjMT9CeWd1
0zjcqEMw/fE4mc5uKde0aHwXrPSKhEzFTFjrlHMG3Xe8Hx2I/dm0JikJ8u4m0yYULVLfs+rB/6gH
c/LQ9iMspEBUEAlmMcT+TunesyplIARSWCWkuRdiEvG7MPo5AUEtHnk2rn9Mv77FkSuac0jq6pLH
sPfRd+EbULgzgWHfbFXyEEWltezCeb+drfP7dV2n+MK1Gz7kQvpzgL1oNIyhSxmF//bl3EWaI28v
PV44Jk4PyJBY85o1dyc+HCCeyAeHskVLR6JOBuCwjpSYzm0rBLdoW9Y2cx3PAxx1+ajS0udSImwd
xsDfxYHQzfo1oNZm6nxkyaUVY0/+9FiQLHA2aUu6QXnrGOuIpvhuBFmcqYC6TdoFFOeTjXJhJ5C2
sutYvp7kvcvp9dOZnKlvgNOVMNZROrz4e+wZAAIlFTFLgpD5Qekxi0i7M9tFQF4OvkwvflVsg6fA
nIzwMWCI+OM2UDAVHMmTObOrH98W4ulGlEeTveBms5lnDsmT+ATunt4WavMXIZKfhPz8+wPuWsB5
7aqygLRtWqpfVqnxmsDZ3aAJX3oGO5US7HmTDACoADE2m6It+nkBEBZq5FKsoiiaFcSEvgfNmxRk
RCFoae8Gl0ejp/1MDURrQTVoH1uLNetxvthbGtG7RgeIsoOem++WSqA3+i+9lQqrJSsWAQV001rF
tMIiLt9esVrYrVKi16sqpOglrJnNx8RE1cpPyRnNpXpI23eEfA5toldfALFnbprCb/BUdTaPft/V
scbUfI1a/egUsGCbESRFVYiw6sYFJ2m72ghTQXcr7C48zzAzowpny5zXhxvwC0+xzuocKr4NiF/h
CPZDT97gM1MIyeCM5QgHUTjSn5VxWEC+Nt+ouAyTf1W2xrDxf+M+UHDx7gUV6A1w+yRkGN5W5w+q
rGCs0T4f2tI1VJcpLk2tEdS7hYKsjPQ7uittAaV78N+PYdMspdW8EZULeg1U/WGdEDKQeXl6D2tk
I0Yl73UYZV5y9NE4UZQdtw/zJpv+MoF+LwirHGmfUYth0nBpgRnqZoPwikK42hpEnreEjTyhwo6L
LJqzJFBpuFThO1FflzQpaHoSX4g0Hie6dNd2tmcuiNXIazKpeEdx8zdDDC0AaTVjkR4tPlRgoAqQ
IZdmciJYO2shEYfJ7jRZ8n+obG/SRmI338Z3p4uce4lZq+c1+ypUgSYDqKnpBeMkLB11neXRaTD+
T+HpLj5BUAc9A8mR9v0CORYzKWeuUuy1w4GdNvTQNFUrZtgKAhZsgreTJXWhFTcYSltnmKs0s7wo
F6YJIJEv74bwV200eBdLAqxOpPW6ZdxjjgU3LPql5VUDPo2/niatwRvAYeCIGOk4JOvYqcqKbcCI
bl5OlhnpcOo2WAQJaTY/wM+UVHdRCL0R6+bJDgrdQDv1mzDtHNDd9mciL/7UjXg067JhW+nEySbS
2s5rNT2kTNmUmYzjOJnODluo7aSK2++i5YD9VTR+LjVRiZPAxE0GZfW86rBPYNKL4t42sv0EKGVh
DyvDfNp8mvYikm+35gQvjuEqp1ebJ7G8UWYLThh6DOI8GsQGAOSM9yXl7YLcIqbrsUrkBawRx5gV
bEpR4RXVk/6E1j2WAo+1j/RpX7c0HyDs6ltb7HGLGwUO6PK0dZR+6m4IF85LdHe27vXQfFQYOYdt
BPi6Rwcu4z4B4Nh3IR5zp+LCZIZaO+xvpIwZteiXV6e1uQICUffaDb2getrqLYcRnZ1eFm1dpu51
MGmo5D9QMWd1QPAp0BZMUUVKdNrNx3ksjXsEsSTxTPKtUMFCkZPsHIlcE/8CoOswt16FOrab2KJo
mpgHqxRdIgYyEJMgIx6XLzfCxbWrbeHn1WTzMdfDrDMkbQQx7KDqxs0omfGPWFlEAQm8bZ5Kgn75
L9lzs6P8XcrrSMOsrXxIffJpOzT0zFpMMVjdmUJpNW+AZq244r9xNP5WCBIEaGsnC153TbUdGNpn
GOSzMncvzVFbS4+iG9583+LPK5CrlAjcRHQ/l2ZewWUIAobnOIpEAGxqYNpGRDT0NQPX/EcZRry3
tWcMgn5aXp9Bu+y3cY0FRdu0/kXuuRXGOFAGY/PSLWbi+CGo61QLAdezDoQusP6WM/h+1ydqtRY7
VLGmcreMKjMCQvg49CdEQw82kSJ2X1X0f5Ce4Gw5XcgzxNwiuBA7TPE99rNtoDftXWc+CHKKTzgj
GT/R9u0Ccuiq8lYDvCMHqsQXdJkStxIMa38TkvZNS514XA9ovlk5jq+Bt79Dhfu7ObttuSJGn+aS
cOA87uG+ymtOOyLKbuC/YsYKFTFx2GocvhJe5OrD3YUfJaPFv4Tq23IaYXtvZ/YTMJy/rAKdEmmD
DhYxaxyF/3IZYUzZaHM+619LPA4u3oPEAgsX02sM+0/Tib/jyeg6f4RteRjedXdbmsdQJHZ0YGll
yP/poh3MY91P7caCJRZbL7HW/+Ty80vakdmCbMTrs+4jEvAbuBq9l5HEoPzojboHfR9HQvq0xZW4
ziBEkEOoOcUETASs/IgBHDdzfHb5sLytMWhte/fDwaj/3P3aYo4N8iYvjXLtKL3fJ0SU/eatZGoK
VQtNOxr4g9vahI1iPkiQeFY7cz//lEXjm3y2NszYAaUsWTSAlAXPF2AauLZuY1pDqcyGoHR5DT25
CBp6JMb0SvgqQQaZpEKA10G1M0OuXo8k5M8hqwrW0SDgfzndKvQrgal1gPonN6fgzR3x9Esf3KuS
AZwMQ8bSFaH3tVLwqtuBS0yiWO9zt1jh8gZePGOdmWgLcHjPpYUhe0O7ZS0smPAfJvif8JhyGvlY
RGcsvqftiQQo/+7GCmKHJzffjwkA9Qcwo5cGO13Lrc2Pg0GtAsv93MmzCSWLdfmOdTM0in1GFisC
Fw4qXig2NxDwuLSWdU74/Gj3uTXJQIjFxHQWJ6DaXxlxp8C6NyXbvWPv0qgdxfjVKcau9ZY12eET
nEQp3TzyAp9Uv4Agm03KIsqq503tIvwqLLsPK9SilDKNKJkCx46o04R1LnWCXjt3kXDmcW2DrfV9
m0GuYtRGz4hqXtkXLWEoSMd3AYm6j0yWEq0DZVSbn77QqqEO2w60Qf+msi3t61AieStrspZygjpy
UqW8kar0OJZpLIIbNl/gVD+pqN5ksBq7goqfGsrD55/pDW3tFO/9M+Uol5MwGzcfcw82AKYo2ZeA
euG0IDD5uWsvly0rnmf8YcT9Zy34O8Jvk6hd44GTx3QjVGhuZ0TF9688EMMEJ2zm+CPy1EAICKUZ
5gGaeER78bvs+bsE9IZ+X8hAE3ykNMtMufcO2onf+rYT7F3Q8NdVvgerAI/QYHCQu7LE1wDhiOh+
yJFXGY99fmbl12i1KzeRurjdrNrOdm//7Elx2D3CiEFi61O19D8rk0KTq2dl1NehNVlfNzi/huPO
ISO3gf00CQw0wqWImOfNVRlIX+8rHvEjFLcHwTXpYrbc0TGGjen78Jp3U5tbpXAIar7xSGnpKauZ
KIQhYcJVp9M40vKhT2rsNDZEOOzGkRkaTGBr8eH4hr+TwOXe3M65oDK52u0oRODyOFMxkyoJ2keB
35zUvRnP++idDuSDvjMS2JljBVRKacYIsA2i69GlGIj8p0lfP9SqKcwktm0VeGlw1famC4vzJlxY
U6VotcZhVL53agjYY+hV9+UXRUWyTJe9DR9Orw0TzG/lwyQVs6ZA5/Ubo2ifM4+T9EsjFibiVj+T
Et+z17vQLA4cDknPf3O9Ht4RYF6NQbNctzvrgMFdoLHhdSXrXJd4r1hWYtKeJoBS1snyj+dHvIUo
qmVGQWwwneC36IY+cwAcVK2A7rib7qaGWJUhOp1SsSGwYaNPhWeynKgCvnWU+yFLZWEv7TD4942l
cu+qWndkoh1n2uXCXvqQvgVd4Z5twhyRGF+qi8qSl7fW7x9+Ep8U8ebAeoVUAYfA34lB+IN3CmkM
wC8mUqp26YmU8LVn6LCHg/W2P9MiOudti3a6qLuCHwS3mdvFYZWDnsoyP6/QTAluEV7ABXxKn/ue
nzb4qC7WfVeUm9zjR9/tuAU5B4baU1sxnKHgMzwzsbm4Uqs8Jxe0aJz/5O/V19g2LM+08NqCxJzm
TJNORNILbUatPjAIdIZZlbRYZp1iBuPhTXoZnb+MHQkQNW/Vq1i/5H0TC2eUaFKUpzRxEyKBJ8W/
OeT9nyZo8iHfBvNMORI4a80zcIKo3K1mEjIaooc7YdHBZPZPwZj324QdYRJbUJeCz0QwRLZQ04Gd
+HoDkfwFWdknLmuP75LSmykbRNQrIrhHdVxGfLi41eNu4yRhhoaO4vf1plpm0RRUgw+KLNqO62zm
6PClHwsOVOFFA87NildmuQcJ5XehiEsePsA2xxNpA6r170FGckEFejxDw1ls7iPTev6DnQQpalfx
wuzG/hzC99Uhixaho7/L2y7jVH6xsEnowYzFTZDZP/BZOIcVYLmmflQADswzFjMwWqrOGAlIMBoc
FaxqfQp15a6ZiWfDK9qtEl8wis6aSLydTf683dYGzFQIyPxDSdQNjnFE+SgnfQ9DJyLLnL+TsDAm
5th+Fig48pfyOp21w1/XCBBSHpdttnLxko1a88+CjFpIxeLAJXmEC6wSJ46M9icYdhccsC2OI5or
YZDcd/j+A8bTh3L4bHDpqoHoqsVVyoplSpvuey/jpk1ZHXuIKMitwLhbxVYd+Dip4o4wUBrCmx+Y
+GSHpGAAHA+JI3ZCJMgz3LuVBQFgwhbrfReaATqsl6VxyfhkYyO1hvRU104WbQfkvpqJ3imLl1U6
9QFqYKDC5FiBeQqorK9X2s7Et1AHH1l4jLYm+1nX+vXJhOXBkuYnmWhp3rP9X4eoHsZG+FygxaAu
QYikA1tqDJzBvAXSS7VRNe5tIGtn0fBJOXstIcetBUqZkwDR6uBFPwM3o7qfLx1D97DRY4zILcYs
RwZgKRrD7JMEp2YPYuxUfJfIl7wH44lg9I7UR3LowKu2/XZTxYLCnuYQebdHPzATKyDhX6I20Ulp
6jRWuylat0eHnXhb23vmb/CojE/7zhH0VdJv/iP1Ba15EoQt6wJflSSkqhyx1hYeD8tswksg3o8J
wgfK9B/1iCrVOUY2dOWWJdKLT5egPP/9FutmLYlS9MKbrD3s78dP6Gclw/rSsKcFNkmzuH3Rp4Nh
cT6LP4krM5HptXlmDhhFBXNO7bkEF4bDbh5cCXEZ50K1E8JMeBjnorABN0axyzG+lwYQyTmvBIvz
0O+qJPKZiR7xW2o9R2XcRH2i3Ijpg/YKJYNKTjHV8CbOaXZQJl7a0BZkRPtGNRLZlXMqTjMkZcyL
DihJE5O823enJczwUia0qFkud96Ptp7YTkKSwa+qZHTY8TA3S+FUS1JIID/s1IFzetcfWofts+/8
N6utBgjlHdmiNjbhAN0Dj/oxVI0LoLXcT13ILjh3AjdY9HhBK/1Zkv+jzPPgLebIApDs8sZI8Mm4
kmYOomarqVIgDMxO/pOdn3qmf8ot74xzcAuE9RsZzhpnhQyLQ9MeMUYHRspZX0R0nQFyKAILJWsx
0PR/tJybkEG2LhQ+eJpvIHXnT+T391xiFI1LC0Et5BWGNFK9H+VSz+f2mUFIZy6XYY4l4za2KYeS
KQFIhAiTcSVQTqmFV2OQX7TPZDsPms0ybQEaAkZ1ek754+S4IB+IylxGatuCPAk8ySgR5au4kr29
WXnfxK3g2hgIeRoKwv9IXLywnjkMcnLDeyfLvgbR7Kt9BLPzKkkvNXK3iOT9dV8uC/Fa6sM3WDuB
BV86aCdgCOg3p52kKliRgQ3v3KUZxtIp05LZBhTlZYCAeELk5KghKW9PTKptGEqM15IhHpy/Nx+2
ppl1Lbfh5Zj9RW+69g4+qfDnaa3FFZS7sICItceHUB/usTK8CVJYMnNAEPBPMZ8HWt8aQ4Fh8vxh
x+9KYiWx93ucytNqGjEF+J/wLRYZYdNLd0mImSm8m7DT058IAdbadKt9NJhdSQYMNss1SkwAjJG0
Uu3PKZ0VE+iJofdowaXQUP68xV5ovLzVmvpGf5/ojmetsOPqFZ7QjnTzErA6dfDSZHahA8+ZbVvK
6ALdc2IJRIH+r9lbdX3wUWwJm4w92CuH2f/D/qwjNESt1nR8na2n6o69ElKuib/WWqO45U70a+in
T/guLJDXrToO00GXCkmItnwB6408yVdwm00FlJiiOEjrA2Nt6NCp6QVGmOCQhXrzZ6igNCIJGd/l
ZQaj4/nMGQ2ufRW7oqgSgUcEveTSCY/2vxlBF2sNM3PiuMMFlcES7I1ffzMNeePDen8nAUwRC5OM
Y0gwsQ1u04BeQARIT24QfOr7Jer9tSPARDinpy4P2JhMbBPwGvPu3ePTUs6Hk1EUcEMqsd91isxr
HltsEzDygvQhKWByLLuUu9pROAKxdLaZMdDdzXtAtYe2zJ0wx5Hl7nVfBb/JyRJO/ffTSpvviDR0
5pEmIfN1zWpZwKwDsI4dUK8ERtTEO3Ed4gsVMzdcfe3LqZx9cZA7C7S9dcZ5q8moDt951MMEL3Gm
Tar2vzCt3gv1WRcf26BMGHwF1ID62fo8UVAcnQJi0Sq3YAg7z5QWdpQQL6pISwJj/5yKCPvoR8p0
lgKOxBfEAyDC8wP63e8qUI9FTrQYNFkhRDEvJJafnXAdWLiaWporrs49LkhR6m1sas/Dfx7euNbD
L9/FUfjjvaTiQAelNRHZ7G7jml1RoUiRFEReC6Xdk65TnElOuqoyxzbOfU9MKu+l34/l2s6Zv7yn
8Rq7bMGvsR31+nqZlDyICrCH/MHJs1s6RDZDgZvnHH7yn6gM7Ry7lg7QbN8Kz6w2P1PkDUccdCBY
9qK4Ht0uBj3JyGvDqV0M4spcF0Uz4/Zg5n+ok8WJF+TUfEIcwJf+lUTPLSltDGZ5JoBZ3wbQEPdm
WKtL87gQz7fq7epZ06gklNL2ue/gvzukUdy33XTaVlgE6kagOVZyRSKS6ZKZwgBvU8CHcbGcsvfk
g3yAB3EefKc+taztfemXpSFhtkDa3u9WaQ9gUuvpjlMHzwL9HWIEKR/bGjGT4+NwGBFU7H2z8G6B
2EpyvMHCSpWqbXqkhh2mz91l1j/dbjlI5Py+KB5YuBhZwvSEaJyOCW8kkRPcEQXBbozpFpha6qby
UOlGnAGPXgVWpFzipYSjHZZcT+0Qv0p9r/BIwXFomldw51/BGldibXiXZXpTM68wcUPiS13QRQoo
NrIZegTtzeTWfBK9OlMN12YET2pwAADfjLFA65zF0VXL0TlbhEkdnS/My5jnMalHwXWuzmWzOEtU
4HlcQTtN3qpM0K7DTGC2IXckFxjVPZBF+cbZOnIrIq5Oeqn9Mhw1eW5R4rQ0iyDYgwK67Sv3coBI
qvzm5bmmszqEjK9723KiiULKKHweSSuIUz0PEx+XI9qP4Px8Sdc6SVhnJJNPQum1VHbHWpWfMYBj
7Mz4H0mdRcc2X2EK1KHNYpZpJUKEHmUTPeYX2ROwuooYAh+/KFlwa9wBGjhqVagGAfg4ltnJVgRZ
romYTwPBS6zXw9ktuAgzzqSWcnANI13rSbJAH3hWW9Hqlc12GllQcP66zr1BLM415SRZEpmLwXgZ
K+Qy4xYYWQfXmJyC/iXzy9liZQklEGwfQeKQ+GzyMNsDAoj5oOVxMG7b5KCKcjhIGYFSOONLcE3o
cnSq7JpwKHRzWvIIk7s/CDPzNDhqKBZdAKNEmVZPnaBazti+CZ4itCsek6kA+zSOpc2AFpnThoVD
LOjEGdbIBtW9rolbzz6fKtqwf96WUNONbHNcGaFF0nav7tKBqrpNyJEHFuG+ZSSnBt2yb+b98fZW
aNdUdUQrQRy76+c5qyqXYr8N3M3WE8ZGisR/roUpF9NM+yhvIuM6S5/S25I/qDtt+4zh8qiqlK8k
zBQMgbr645Z9eq86TA8V/lhZCKavzSMOviX5kPAMZ+ruUjmGdpe4Zoe/Jk/gsEPGhREA/fhyGZnj
PMOaFFzKp1mqSY6MnEDue+yOG0BcqEttj7RAw2V0muneBQCA/US34qCspYoq6Mp8AWvYvrAJbxB1
XSJ6/UBol9b63IiN+NrCPyU3d2g4Jy14IZQwPPhHDaZF4QWwuI1xmbSPpUg5o22wptO5aZUn9D0H
4jRqCYwZ+NKfIIhl8Vho6qZkLMYBfoEVkiQvGNEgqY3i636i+OfE+jC25yKBLCZze0wd6mgbtGkw
fny5ggCsMQ0u2yFKgbXmnHK8e9Ds/Mp8CBpSEkQl2GRB9+XZLg7q7mYlYcAY818xVhg0YF+4hKsB
m8NIshRgfDxTKWgSaSx3uZZbzXRNbEZYDf99caac93wRmx8QZX+CIoPgFW/5P7ms0V0SRoVSXPq8
W7E2dZaJ4LVhXA7eQixjfQhDvPKZnpKzDLMuGOfo58lpUnL//46ykX3T608QuYKKFspXrMo358yW
2ICb0bwaEHTyT7UKhOvGlzbxgt4IOIz7YUe5d0OWpEwWnh3IBccCkzBMv8ZEauN7lwxltNkaNjeD
TkI3pmOABEwGo+k3a1NFjVotrJvlKJ6E0hPeh4TqeVu7GFOisCct8jkxOD09ko1B8nlubjK+Q0ls
CcnucYQVOtuWjE6PZlwPTlwGfHkr3MhDDr6ShfYV0vbM9P1cdw+cyCjlqzUS7mfq6jklhptJZqDf
6oqw5cwuA7iXDgayn1CaDP61R4hD5iRfWJnio6zw4CQwWStbaZGnaVv6Zt3Ih55EthZCvzJR4axK
bPMHu0/8XwwO1MkCfy1/J2rLYOZR4bBF6kGRH8NKTbv70t2wI6wkAzRhjpFvLMtmeXWnlk1RlrfV
eozFje0vkem198c42LiCW0fuVQP23bdhTYY2Zc+Qkow+rKPAqNbcTu2L5huxnaF12y9y9XYjLTVo
bIZTWsLmsmjwy2BjVNoQ5oSvZ1zEaDU8ecb9K9KLjPan1bawT6tqDe77F8YWnavucqIw/NfSJdLW
FRfO7g7aLQ1VUbCGV7ko6Ft08QbdH3JTuDfDf4YuA1I04YWgUZsLA5kloPqcl0Drc8OyPs+WrwiJ
qyDqJ+1IAbJHUrSoQO81g+3iV4kjwnCfu9mlUA5h6LCjkrapYHomMJqxNrHjwcgQmEEDKI+JtH8m
w9yyGJ7Iagqy0CSi7CVEJCgVWmWfdLI5iXdcHVZHB/9MgfzBDfmGGd2h69d2r6Zm2SBEahLuwkEV
EjoZeAq25Xd+HTNIUOqpgSyh9XZ6yTTTFLiUhFZlK33MRbUfgc7DEIo6fMWCmPFixajdxmUd79XP
mc3ccjNi7bbD1jG8/Z2ur5BWoqlrGCBV94XHXqHDVV+nUFeBr7k7IYH0U9uH/lMHFKrSTSSgQvM8
ip9o9Fiqo4RLcEnMEP80fy8CEs2WJH7toYrvXu2VFxU3W8u5EYj3MDtWjWj9NuyuOY4t3HGiY+6l
+TgOeHXxE+GVaFZsWVJp15jX0YInHDubmWBzqQZan5+5d2g78kcsaFDCXO25tfcEfw6xiTgwvY8D
0QuZIKU1wUbuE1zqly2AcTor9fNsHYA4Knr1IA1tgb/nA/OwBlTGdVBezYygSWG7qa4EQuZ/LTij
X9D++Tb0+9Drj3wmboCsSHu9qneAwkt/lDwXgFN5cCF3DarMdeSl79AvW7fbl5YsTsvxrgowUm/P
RO96bzPSAZorCuN1ZrZ8XKR0DfWUkhAavddMElCupc89a5MN+umh+KK/UL5sYHxjObQaGatAZkNR
eaZ1nNvIlMAhbI5Wb4bmWQt9a7VcA9C8cnIUaTPBmCohqESSWURgonmjzGg33J+a1999Pe7zCkpN
1o/3uZAKpxiDf8WoqSJDQszHEWlJd65/vdw+YH2hDuHZugrftHEfsRW70JLtXDF4xr26jM2N8PgF
NhBIrlUtnhCvANcHN++qs9xBp8IH9Vww8w6h14bQAx/BlvUBUZ6G+FQvr/zjULl5qjKernZf5CJc
EirQuTtYC92pEgAA/F17hyF50g2JUGDWKrL0cMr85yBa7noaIJ/AMLNZB7FWteo5F8rV7xs6BANN
8oH5c7tNJIcPQD2RIgOvQAcpI3Gee+QzyDoPwRlS1yDqf6REKp5fwZLdwVz01cQQLLrSJLfpi7MP
ZXFejSMKDWzEjkubaIWX99PIwKXq1t/8C7xhaTx7z0gG6GFK4Z5+t1OFy4lOuHcqNTKeQdCF3gxu
2K57LDHiiBeQUa9PSCoDb96RD83vVE1zKqB/QYfik6t2kdwicifnBlcv+9++wYK5CVpOFly6ZtOa
o+9G2vmoUTsiCFv2O3M4723QP9uDl6k9nUx7boNu65e+14+dpuDBpXG645sSAdi49EQp1hYojv9I
ATuA2mGiBYj888uouOqTN8b3gGGUcIiyMsx/eL1oUziEbUT24mnQrI+jbuVMN3FLnh5NaKgIy0BP
a3XpwtJhUFy4bIQjDBuR4smPAOqpT4CN+5e9XnwLAkTGki7pymN8P/G9488Jt0x+zcoRjH1/m08U
lODeS55p6dm8ssDZzFLy//8G12UImR427bClVzjWf5tAdb0CgtPq3nDSQDRCE4nK8YPS6fOmkMrr
1ZXCKcK5046L1v6meS7fvAPIdLHTS0cczplsNEpEO9KppiTOhiuUreIWDtRxW2MwL9Psp+o4wix1
SHevxKEd3cljaUDD9ck34YQWQmMrbK0vguBIOhCrjK8E9oEW6aDDbdtMvywc4ZkIWFzsXaEeUh4u
FcAr+OQUZfO8W1KkNzJaQSMllTcYN7zmFrZg40N4W9irwYw+ayp2Law79MUKlBShfUmhJshYrcWt
FY0wSELuOM7xi3ru0fi7optB0LYxzwl0Uy4/r9PrXHkdzqsT1gE+W69Yc4U1d15RLf+WJ/2E4sf2
hHhy96JKsfjzCk2ZxCy/kSSsgnozS+NzBXjRLla1PAfqE5V+RDLYkXrMKD7WycCEPOPYMcQnt9Px
G1Ua8okqcS4BqvaB/1DFsCuR2ru+zJVHCRtfwIxNSGJKUiZ7iUrHCnRWYfEkldFWf2BCI9W4MZ4j
r62QgwYMAqG+u47yEWW8UzFewP4ZGK9hR+wUki4S+RrLF3UkXrgumLqWBZUuZvu96+egqCPB5EKc
zVtanP76smuTeGzjrFmaJkRRAISdrS+vpANaLgBPOqCKfTWXg+nAudh7ruZnuUpsD7njzrxC2pgL
zeCKGOfs6f4BcicptIQwuMnD12o3FH5gjvRSJIjblHbX7zSClYxV9hdXRmPZIo0gaYYg65qfVGlt
dQ/SXAhLc1EXmpnmAenYDTAKz1t0k8YDF+9mX5NSAU7ukPRKr7ei5uEWm8fAsN5oi2fGWfZXDz6n
/rqhu4tFnxEW5+Kofuo5dEoP1miWdqe9wTpuyAXBgH1TVzSy4yGLQIR57df7gOL54lxMNaAbccJy
8LBannUkPbZ+8YVYNMG5wfkMZBBplxkvGnU4U+dSKTuBOJro+T4DZprzni+omhlVVdDpQUxv99tL
OhrxvguFCEElZI2iDNSqAsp3d364L5YAE+4c7/ojoMD5dFcJF/v4hSsA6CoLAMMivXYKRsK8K7aM
nBIOAdRMVFriHijtrgJm3g8GOawne5RSukc3e1bp6MQ1luIri5xqSxAPffOQgwPHj8Ax1ILw9S30
UVyuJOzuaorg/OsMHgxYhpBltrP6w5WUVSdg/lEad+WGL7lw9KKP8i4ajey4a5+kUZ3KB8Q8Em74
lw/MBCN3UN2lm+LcGH5tYcEl05wsrWg+jjopedaUz5Nnb3wI4fnKxh410comRzCbyKUfXCtWOoeC
iUPu05dK7Hpe2MXcDNC2maJF77405zlcGb8IHUnxFlVy5gElDbCNjlvhhA+gMJ6F73L5vswkKNks
fvgTbgrRnRYHvVXyMFECVfBEMQBHyP/9wp7IG4PQWgbO1IiYekpVygLu1hlqGZOoQFH2ofhq8QJ4
+uwsEw2mzJK+/kyRTmbk3XxybxXALRDynx1OZHHL2LNQXuAzG8kNGZPd9n+17JXbfvwAwOzN3msU
XB5IOMncYeet0jshoGK+jb7FBgGMcw7Hw2dX9Xqq2sGYVJ7qFuhpl17BR2xpCvs4NKKpp/tdHTEk
U0fmTBVv1Sc6XQxxwK+IsGlDYOr2ugBXQ3FBAreHbkuusOa4wydAj5eAjG0Uwz4aj8ADrH7UjVwA
GmoMRge3Dr1rQ2DkpumAi7CptYGoZB3T9w1cvF/s2M2VSx3tlYwoJ/Y2bsFbRWGWAh5IWRLo2CwO
xesDe1fK6H6me4I3g/azGHD5KookC859IKja6tMo7QZK2o+yC/5AdEtdWZY3WvkRnJOMjYKDAyLX
SLD0BO+Ub9+PSWCN0ete+jln7U2TWQuMnXq8aoWuEdoqB3cB7fsneeX0f0rcsZS1pNEe0zOMgwZd
X4esurAR4a9iWMjj/X98nSsqFTYQ0iRshvLbhSfI+1tcfdHtllZl3GWEtRbQ3/yIWcR2PaQf0NqP
RNsG/5HUm4XFTf3WVsFxt++mmNR+Grrv9pDjffqPJILRpVRiFD5AsG4kwwEHUJ1LivZYlh7yqZMq
uejtILQw8xVxcPRMLCe9SJfKg2bIJYLy43YJt8r2mI7uUFI6amr5/3IJdwNkjufoQECtSCnzG9wW
M5ea9nQLIheH3gHdMG8aIhFrMpG2oiEkl0LGro/0ZauVK55sIiL4HjNeUsXQauEliPMzCou/hsSv
fAF7V47Ub/JkNUJwOVHvoOfsTQZDBVqILgLY1t7Vxj8+bMEKNb2zRgQNvZ0orsoQVvAb1Y0EqKy5
uRzRym+6NIdvs3PPHea81qiNKISieFI72xdFvQ+pCInFYHQWULvqYEDGZLVDuJChP9YKBAmez2sd
zzsx/YHb94F8YBe4Ipo2CRn2kNCCL4wBPUbGEoFJpS8cra1dTpIPoOOQyknxMb3wlng1Z+BkfhkO
Et25oyU/7aQY9Sfx5Iz9IYicedDy9XoUjnOpaTCkt410PBI09b2KMWA1E6BPw08TDR9oq5pynbjc
BV86GW/QW8isYU9hMFWxbYkS9T4sgyCbSOWo8UkGIrAuGop5BaK+0IoP4zWpsufnGi+qUNgDsNXy
qZ80kSoME6ek/S8H3RmtvB6m9cSLNLqlIMAVo79pCX4qkkFddlzxQdJtsxx8GZPy057AswM/F74G
9c79bb+o7dxEdybAxF+k0YIqRNsWxx8umcCO2+RHzpySZaiH+TTcMpWLlHUwNgX7q+uS6dE8g6tZ
LkOBnzTh/xA96xAriSerx7i56LytOoGVRwVaAbvr1FtKrfI6OVAZVbDNj9UlzZcPc2Qf9Rhbj7B4
Er58NhGc67XTyartwJLRweW8jsW1dV2u5VV21zZKzHCjyy4ZiCPas0ABoHrr/ZbLp4XQlBsmndt5
UTGlpHQOsZKou3fKPYkghaHbRSUVgeiKzcVe4f3VA9zy9wAK06+xxQxyCj0c/Z7JcFtZ9GIvQZid
ZfjG2SXbPg3PO+bJn61DwqKFNlAyyScRMpchaHkAOWvzqxFd4D/KJv5P1FIOKf+Ftmz+i3nmloZO
FFu8pXjN9oeEXiE20qdQV+AU1j8E2AkGCwXW8KgkecfphwYSWaiGSMdlf7MMCQFBhHKN6XmRTjhG
zaM5SykMfR6jOV0mgzH/pV84gX8uR1xOm7N0MsySJtlumvnDFegcr2zoA8jpp8fbuDMxcyN9HQNs
s2mA5Z6GHXumwAsulGdFP83v4VRAWgRUNbe/DroicijKVYXPyHM0fZg1OtVol752eiClz9HZOFhC
aO0vvZqa5pn74rYhBsII43EJtOTKOno8S5gQ+P25cKtpG+CeTalrivwUE+lz8lhgK4A3tHxi/pp7
WAYeQTb6otGHPNZ1ZofbxWmXmROI4jWkt84nCTCxr2VuSooVyZ3mbkMaKJ6JvIcU3QeYRR/ZJw9s
V4xKuDxOTUIFv9vq4rx9/C56ERGZcEwYh1QXy1RYRNCz8nh0lgawxlBt/yM7q2BkHiQi4GxW5CGR
UwfjzvEYOXwH7ohq4vH7tfUGB/rcXdhbjBM4W1A7sNUdwhN3wdTd0s/QbRDFZCz8+IUjUSsOcwKi
bd1ZAW9h4SCmFt7LzeEQr5f3+UTlqkM1O43wAZkqkpUrZYsWa7K0AcW3Lv7RjrSk3pA0h56peHpC
UN4YzHBoE8Xe21KB4AzbvDYV663X+sDIDHkiPXZzmcQceiRtbPs+X1u34mhQXuI7L0T8KkMAWI0H
iti5O77DQsNuf+mtYuDJj1u8QdmxOT4dfSWqt2FwI1sRoJdZg22LpshXf8n2rGEsO8JuZnCCJ2pa
sovx5V/iASP+ApML8TJ8uxWdsxzxO2VMgxEzluSqEb1lYvSJJkE7qOEMzVQzfzLrQb1fUVwSVOGm
WXHT/QsSLS/DrQnEyxdAFBlwYV4QmG5wdKfi2kEqlcCijBEgMbq6AFKYsSY006f6DgEOVX/Klzex
Zb/xsAHwmFTpgFk7AvH5e2a0sQ+QILyjSOeI+Ues+/W0b4PNyZtULtEbgjkp7LLEL87iY9Ld/q1k
/04J8i2UdEJ03xXZYP+OLPY3g/HwQxtBZ36rfSwnVRdZ2RAEhYZq++jLpwpWn5Zyt6mgfW1zD0Tx
ZHRjnPtZx3JsYPiNHhbnMxNydjNPJWkLC5CKisaDbP3jkotnKDHyuTHggHUf2v8Wt2lklXqPuj7z
RrEzeTyl0bmfTbxR0p+Voo6Rx7ZOtQ4Vgg3Z55qBH6whQU8Kx4qMegbVLvNYjP+us20IquoGEDQ3
hWwOSQ5j2txB55gILoyxone09G7WRi6BQNr1qNOn74VCe8XhzvM/sQmzoZyywlkzaH1pOgu7MORn
52kfyueU3OJuk+Y+NYw8nWSN71ncwxrkm37++3jGaBHR3NaQMdJr+nBEdI54qaoQpjwF4GUs3EPL
+ntc2n3bPJQ+nPtG+5ujG/PopacqMYmPbILhABqUagwWJ/9cZNf4Vqu8xeEza9+hp2pBK/USVh1Z
dXR5bx6DRlhh5cUKbvxZf+11/Q8mAbZmPzf03+7plG0z3dAw4tZ+Lq+tSvbBKwQBfoNbnq7lJk5d
RcEFKEcr5yduiXJ11+Jnxy0Y545jBvITuLJjlcDpyPcZMu95Skpg14phYq8/eNuQqz7ZGXAK4+BJ
P4bx7rnnsZR+IUiKn9QUocBBRvEatxEbqJQxwXPq948oiiFJ0Hf7AVpswAxv/4fGwgeW1u4xCHge
PENKdDFG/uCgIWtHJ5iuNhxXFJbY23Dhza6GrR/eMQC9Cl3xZFhXrynJ4SYR9y4HoBmJcTEa4ao7
l4Tpf0G08obb3YcXTnA+bGXSqbhco3miL6HhvT1UlpTbDqCfoUumhUUhqW3VnMSfq7717J5gGJtv
HUUMGaIr8FEpF1pW/U+q/8V7ivdCFy8ZzeaSSCIdTXIl4D33CTkbBikklxJW5wfJa4twuTuPWVYG
MmX2PuboY4RwESAatTsErgEim2YAymjspVgfAytyFSgCBJj0HN6GQ0Q6tu+8iJwlUbwZ8CajTPok
5OmXg9pR06sRQ6943yZ4BQEc+/8aVDb68Ca/O4l9QzdFx5rjMqGtwk/Mgon8xko2XINssazgcFdD
B4VQE5qs+WSkBqoClPfMPYkGeytBM9g9MEJXQhq4e5/lxFQ4ws8E0dfYMIYDXNTYe5Pgqq9ylZm1
9bF1CSdvJrCT7cIbYbng7tI2pbpmplpRqVQ5H/STiurcVxYyNDUh5kt9Doz6DxiSFyuB0MfrJA+h
HVOjjm3S5I0jo9BArCi39hNDGi3t5BGS6PkLBHJ2w6NFF6BlwC8Hjbtg7ysbwor2XMDhKEE9p6ih
O4f21SR5t80IJmcqO8Ox1FCpzTnaqUvzJPOorRgxxXrjDRA0VzuYfB98ZXMF7I2ypAvqt1pZUxA5
+53aXbxTbCzuctubULMcqSEH4JVEHbZbC2uRZWSgiUAuUYJdv8/V2vQWV0Ci5+7TRI8iq3jLudx7
b3TNDaFbAa5dRcEyhRfVgzuh31stfSzOTbEjXDFCj7f59VbI1g540U50pFfN6HEhelVOUvDvBrFM
d77AQ/xKyEbx98oG5yTUFmYT2BeOaBByjJycnzeLuCly/6v2mJmy9dXqlqYTCIoVVtl2QNlL3NvE
nJpnR7KYbiwfV9WVNWxZBtqjumT8IOLKTiJ8vvejVf1i04vZyTsNs+00v8589/vG0YZkXDPz0eI/
wT+a1GhMoMRRbX7wPLKEliM/37ItTBJDVNf9pPrmgkCXQBWUAKMk22RkqML3vajxC58AFpnd+Hji
fuCxoYjS234b56ayQdEj868Eg19e5ZM7+jv5m1UINA5oU0TJabMLWeAhVDsKX+6UcHnHhjqMloGA
I89PpRm8wcmTZZ7Za6HnIzLa1nGe5LjtQK5fDxS8N7+nsJ3+yIqjjEzEWofdzG0kLsFlkzFTX2AT
PErAM3GMOkodAqMalIoSQKYsjvAETx7n0y+OSX+gTQlePgN0465P96d59dYJu4D4xhlutu/XX3dv
uVZXGjURI+XyR3P6Kv4z+EyRGeSP4XIScGOEN7zv6EYAekRAcEQKHkNZ1cWJHykXSl8BigGGgHFM
oHF4k/LEoSDXtZ3P+jjYbJd8v9DFpv3/9/uQFfxJuhf9370l/I1JHki/wlPE/tuG0ygcUiDU++48
HFZxUBsuDE5UZZwRzY45V9XpT55o+jCQqQ1PD5vqTEhQjFuVOobBdOnQnpfjxlKOHM9JrMlcD8Si
cLU5BVgUqWzFBcBMp4uKg+Dh/z58+PVu5CnFjdP/87+b5bglYXQ8s/amikk55KGucgQkB+zAJz0T
Px0jQMhG/+9ybmHLJuzDm2ATUDVhx4wSmgZQCt2VMhdbR+N2FwTrI4rxeC5wDgzJQruvQyKskoiM
xjl0BsgKi7GcUxLPXR/6f3mvScJX7SoIYFHqGtZpGGlzkEh7NCTtS1ZgXfNsb3g6UL6MIemDUsHu
O+H3fREM/Wj26e5vvk44EDp++uVKzdvtwJN80ya4qmeh+usOSfELWd33SGlb/nfFykT0tNzmxde8
f8ii64YT/AUAZkKxZq5OQd5LV/hjBX3yWLxar5V8aMDAfcW70U+MGTWjhZtY1BAPVyXSp3TYym5I
8v/Nwg1uLgM84ZP7FRV9j/sYb9/hd/2KI6GdSgUI+JR9JNjF8vvqhhe8YhE0f+yOxlDWge55FIFD
ezmHnJDR73UBu7GanitP3LJpisjndis4ORW4vgu4MZKBt94fCSJKAcr9j0TAu1MUl/0UXdRL9i+V
/vSkS5uF1Y0/J0gJ5WyvF9xhU+YBSZ24bDZ3XwKu41JTGxeoLjqBvDDc2VY9C/Flyqy7vMNe8a6x
5ycGszxh9anhMUHV+bBrfPR4BSIEpn0+lmn5zKWM7hL7NSBvWnqaP2efO4rNMHxBpYToVbEU9E6W
zqIVfIGQbTxh48A8zboLxZM3EH0RT6XLw+u+pHZhbqBDmXD36JJSOZT35JzaWV8A/NttVwfi9Cnd
YuHfI0i4YdI7Fj25e9NbMqW4z471mSlDuS6yBmTI+rm7IFY/5+GSOTneagD9piUj5lg3VwauF7PP
GzE=
`pragma protect end_protected
