// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
tbA1gA7SmU4J9FuRz6iG2OF/sSvj4azgQdr8Pk7TLQySWHEyCI/xTS0eOhMgHoakI1wG4MdsimKN
x2t5xtal264AJCUPcDooXR8cNM8leeOv/xmyaPb5XCIQcwKU1w+PUslyzMxvpsJWYHNk4aVy4bjR
3m35ogHYYu5nffNRRdZ9BlvcBa8wBoM33KXvO6ZEhIBzRS5y0JHX1zrO584iaJbAplCzRRUC38hH
pOP5D2DKyVmCsU73NFDaCkx7cNJngmySoTR5YxTAIx6k2fXLsiRZ0e7r48zPTjREqeYbr8l3nwOH
Ya7KEi4bfKf58Qf31BgFpVydw1T1LEWDAogW3A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
tYf/Hec3iSbOXZgoilyAZ0GsC6DhrguFOZoj5wqO88OMqd6nctDeo2joV4T4T9xC7Eb3ATjffTzH
L6NNu9uEfpUPpOpdWGOUppQ7SndYLXGxK5ptgQoCjXAs0Ttkcvb14iRUR03IFhmCmeKshPN+cXSV
xgefcxz0KwUZzahoeO9uOU5vzDp76M0nrZJU/DObZKC4Sdq7w33w0QP/a+3lxR52dXk4K7qQijRc
Ek49qM/lSg37gu/wRQjyJbmupn0z4A3qZri9n9QOi01N3uBDKzFmyf2GRk5SxKCOSIxYayJWM4va
61htXKzfitwKOTXU6AKZVqILID3Y5c70W70K9uwagKnL4VXnkzOERPRHJEcOOK9y/VKFGwOl4bcl
7o4vKy+BHZwDqmRFpM+iQqjFyMeU6qJbDe6FWKubhYMvUNgIh2Q0yHiOojk0kigCOP8rTm+C7lBb
LvI0dymOEclXfy4SXDpf9CflErRiqQAkJTPtiTIP8pQKaNjSN3TvF/bnRdl654kBAXbXIekXhMq9
DwKPzg2FCvAi/D7Oh1gIaxJ5bfCvJ+UaenrzMBwupnGPFaA7AH7ueTj3S833Z+797l9IB3YwDp8V
rCvT7jpGiPhQ0Qa5Cu6oLHes5e9CEoYQXZ9yXizFVgehoZT2rKd/fmEKA11bSAsc6imKiiM5JTbO
goYWnYyTrjltzMNrkCv03W8epdloaff0NiiiRQFeFRyCqXesem/xRIdpq9G3Hx9kfpz98mS5Xyk6
8AmwIotS5HHIjM8Bigf7SQW4BSkUVQESDYfGGFj9Rj4sa/EUPwp0iqeMB+AZ4c9EngyHvObU4m/v
AK9k+qceY0CSdTMoN12jJizEEvvSLSvq9va7QpET2ECyxBYJUyHTitgiKTFrLeL8JcOhecuaE0ze
H2wtBGJbCQllk/HMq3CJK03+DEqMuuyZIFQDKm4ev/SzufNBnn81unlBmsG6LDLnh5b8L94ajvnH
GDw6+6LZm3y2UVGZ+1heTfVFYy3CeP56pXYR0tNUoL0V+MR4k7/XR7AeevecSvfbCLd+YfODeFzO
qq6nMMCXhPcWjf8ziq/OrCk5cbFcxROcvgw/3tp0e7Ko5xHG/wGbI4tTj5yKOimdA1YI7x8xwjRG
vW42F1893LQEJ8mDnVQA8t3za5kvDoa6CJP2v10Ho9z/XeMVWHWidEKoyunG3cptTBOzbZGtcQXI
LuARdc3eMINGKcJxldGYAXfRzhZR56Q9DXS4Y3MjvYElL40om93hMPdshGNJ0CQI9WVqudB99nUT
l6tfMFg+YRJUCKltJb8dPEEc2AW08J0WAatYpVbrEPhUVjHQYLEF6+0NBOfZMX8CrgbTZUDIn3/V
4OMOjyPDADn1ZwaMZvb68DIrEuWouMZLc3yQFCH9YakI9n2MybI2neXnmMaxRV5WmP9DDNttn8Si
7eM2V9+JPGPbld1MC23EhzVFK4nl7DL3IZvyFNkb/vgkaRWIH+MnYE1fgdkAOZ/KJoU38vxPuo0G
jw/tjb3N2ApES+VO7GTPgoCtHn56SffIlAvC2yyqKE9VGVNqxUtC9AxGPKBG1aQdjJb2hBXBaq3b
gabA3WGGnD+7K+6GzUYSVQ0ucqed70B+w0mYz1w8/ry7j2Cr3DETe9B/5//E9sjaaMqhAzawCmYI
S8JNFqBIhjeksBS421qs+JhAS0uMZbDGlZqAD+hMYgdzqB1pDpxfEvzZHFYzYBabJAsgiRZG9gBm
CQu9MObcdwdI2y4Jd32w2ol0RljAAWDC89AC2eCj39u20XhO1lGr+7rA1172ge4zgmWYLXi9CKjT
HoxSDVcydnFUvk42VaZl7/EuS5jzF3smCwFgTKJMk/15k/b7fEZMs6G2jPK/yA7PHAICNO2aAHi1
UuBdnsfFAZ6bQaGj/tXnFLiQqVX7YTa2+r9N9TA2Xx0vRFvie8gxk5P2nAvZOnv+9/LhQDNf1b1g
3hPWbZYk/HjBcILK/i5rxRalgRF4Duv2ayYXQfdppb+o+yv9olF/fOEWd70I18z73KbP4DoufJUU
v0uZiA6qOEyHkrT4GE++h0A7duLLO/R58xMvz/6e9nMMI5KTAZ+hsBExdlkkFu4kdxegZ8k+TKu4
va5LejkK/K6i0KTwyLUilFkJfZbtHk8+YbF/i3JLUdvzjgjWs0AHOTQIeCYrgIU6IhMe0h0IZY2M
y4X82NBxa5cz0z9UxZeWLja1nIKRLhiDOEF60dCa0YfPFuEfuRGMnEIFU/hsTtssWRbmYEYDe+uA
1GcXy0EC+av3lh0VbA7ZqUHjC4G7/FmqNbb/ma676fQa+gQOReEfwsGjswNBLF06+cBJumeK2++h
+KUehpXP5frJ4/p7cQ4e/6lns4N/0INxZWMNQxHYcJzUg4IJnPLC76ofAX5Jl/kMWVur5JpH1VA/
eGVQdjJFdgNRg/YY76HxIOBEvVBH93zlvk5VXanETFKpBlBnKI2VkAvaKmQbBKo+NW05eEuH3MAW
W5nGXfAQRjEFigFn/PQJQwCmHfNQRW7PEygpRyQx076J7yU7kkvf0xrnlRNxf/RghzKu2SgXYHSN
qJfB+VdFsLBuMByp2xlbbgAVpbLDYdlgChpr5MJPdWSZTtnrSohF5lxB6wTh5GZ86Cv9VS+NycE/
yDBgiRf88ht+drnL8ncWyWkJgo7wOwBJlrL9aEzEhlFoJefUG7HXLkVXTq2Ssghpz0slrRImmTMs
xhxKMZ3MNlGMX1+kdHEXs+zT0dq1YNkyVQSH7J3O+BBfieQS5lOvFSNzXiyBOxuJzhtg4yAn8eTO
RD8yYwgG11W7UVvsk4Bj0jHFcLDkwCjjZLOZYB/fkNt2PywWk0k/+Xu2H1Xgru6+nFmlhDkBpL2J
burX6TERit+dGHF6fTVlpdec3DhpNy6AEM1RbAAM156HahWcFGURHnOjdKH52poaojfxxbMJ+YN0
X9XqzN9BRNCGpeAbuJU02tPFdhMWs6WH14qQx4JAFTFkq8hMf6oHPzCCaYe0pjFGXuhDXdNVl0ue
lb5DbuE0ZWXvDRadIdeHjsBZ4uSOpTl42O2Gfo2SXlnEkLBcz6EaNmsKTRJ85//siYoWM5pOIxIG
YQPOXq9ZzG6ZmkGyfk4d+CXNIecRu4x6CR7w72RSzo/iVVhMGZCAp/IY2h03VC7AFP3MjV+b8SOQ
ws/Dr7DxFXBTVUB8bFZL9hqpMkABUEN7ojVYul1JMntRdFOegXZ0Nq4NYRhkYRQLAZUe749sIgBO
GZw61PguSLXKRgAwvRMmoe5x+141fk1ojBNmvKydUnEpkE9FPqBP2ewtZcyY7CY2lPEB6zv5bR+A
Qk7lG8OrTvxlzn9Bf9Q5e7tk65aqbVU68ZK2AI5kXfKT9lCMGv+rx8ApC10tPvrAXDGk3IWrqngj
b8BiP1SmUm527Z7ldfBb8PIcURnzXYYWHyXZWZ/rHA6WJG5rUsE842FSlGne9h1eZLp4tLskX+KR
rtToKLanExwAJDL5xOvz73U98ASDARjCmPaO10XUzhK6ssfECJXHcJqBt1ti3ChsMw1AgOC+FI9C
DumhWarsGS9Iy/GMfEDHSzuafvFOTm4FgX0ZqKIqV9XTLWxH0yVR3nXgon6Iuq0/hHypHQswBJ9H
Mjf8+/jIElkIt3DrxjL4K+WBZAtj0JIBmlzw9oqMffWPh513Al3+sz3aIDZ/9IEpb7/5Di2U0aVv
6mn/EmDNmcXoQAPQDy6eqVLCsAeRZ8eUul751Zf5eaXCkw8q+Vdl0L4ODhV2CvHPBwzrfXBtUk6s
MQaq7BvBRlnYFx9cVZxDeMejEVu00sY9oODIJPSFgjzAvj61RgtzoBrrRCMpFSvZW7fwnr+9K6Yu
Y+of/SdE00zwxbaZsUC3ur47SkW31pnQrnDCW+kEhQY/tOzwUPN8ZmcsJ6lZai8D37nFW1zT1n1X
qtqFxeJdyjyGRB73XgtWv6ttzjjrnzPdfAkfy7Ds75MzKInrUhON042Xbafmpox54wfFKxmcE2Z0
c7fktvlWs/dLVhxKAgONj4gae6mbiEybFYEA21UL629ay9jyn6l2uXeVJiBsIHqqj6fARDAlwcTs
vCrCqQUxGNn0Rq1HCocIGJw1qDn5Q12A/oCYyg3XXdhTARR9sKbXz4waq0TwrA601cQNPcUuxU1+
DGEKEA5A3Gh2CAdrkNZopFpzgD0WbyVlJ5XdLPz46BxTwRs3G334jHHinDkjstYyOQ3lwqldwGDc
aasM6KZ79jlilOazruCLABDsHAE+LUVDCdhla8gj7/yXC5lVOH10qfF9Qk6Q6Y/ts6wSYCWf8mz9
HAJwo5nlVb7Dhn2H1mqtujXA2TXntnAE2JMeqrhmBBT+BKmStO8dublp3VHX8rB/nHoqmFf5Yi+m
aJP9byU9/aUNaiWfHiMwG3eKe5/BP/llBMvCnurgu0pwZrnc5wcs7vEvDxYnAMPGGzxk0EL3ir1h
jPdydHvc/4J+oVFrIykg3hUkIwO6UlnhOvFNNYqHb/9yUhoMz0P+jNT9LuxGsVqa4NKxswkYugF0
A6SZ3L86JZRojIRQjUrJ28g+CTO8STuexgxytZYH0rldtSqrrClR1il7ttVg3sXGBbjLxkjuEl5N
bSdfhc1kdrsberek6SSL+CqOG00dsyADfOY3urPVtWGLrQKRVkYaDKfb1Z8Ffv/e6RteQiXAHhDs
gAnIIgF6hPSZ2XNeCMbQTJG7YXPKAIOJH7p18DqEBbFLgbkkLAtvtX/0dtND/2UvuqT29nSvYAUf
MCsKE4MwXiGK9/8JpmBpqYq8EgO1NyBRou5MzqH2EdMqPuJ3HcIq9ciGZ/PAoCqoiz4dT0/rIJf9
6qPum7Ir5FUUgH4PUlNuC2miGiFN34UCqKInVu3GfGlWW7eoh/wExPWy6t2px8Y0VB5FwIJCfYRg
zbKpEf6p4Om3uPxXf7lZPqx9h2oJAkLWhD6RrmYcUTjqY8T7jbeOpOjx5CxLZpyaAESVZalLaQ1L
QJno1Lz5/fqam1L/qJPOOWo0S4Mr6w3VE1jG5MocO7aTQWMjgw72WB54fIiedL/ofQCqaut+zDaz
IDZcH613nQ0zrA5TIABUOv4lw8p9pXzqZRh3XgNprnZNZucXIVgRfJW35SFbo9pFRX6atPdpiqT6
cOmT8XMQa70qneYqjhxY/+cKkmzZAiUq/5tnqAp7vW6yvR1dsAursgGrnecPkrmNsLQ27ur4YINC
reWlJseRos1M3JDMsQ1uoQWDPN22GI2XjrI++PtUdCFA3ixoNbBSzqZbZ9P6iNAEPAPvk517V+fn
nvbHk+GTlKKmOhtY4HMQtOiNn7ZfhuniOE4T7j9Pe3/J5u7U+ApOgSWmtCoMxwEXRKWU+hgSzxY+
7vuoZ+41rmzhXiS2uRwj6VDqEIYgFS9wGFNZK2gVMhtKmQiGar3uNwQby7KERRREaZASAwHD84K0
617h4R9PghrZhFRdWUI80CQrmQD8Tzzm7kijkwfVDcho9WYWmKtmIkJuvJFzUX/Orj9gWsIi1J+1
Va/Yjd+vBHuuuFaJTw+sldl57xSkn6l2oU4mZ9iBUsa/t4ColKgpft8z7mtymYtGy7CIbiNw3lnm
pz3PP2NMF7vPsSZTUy7MEgJS5TUxaR1qmZ5kPIHn1pg3iHMQxmuv5eM9Eet8LuMrq00JCcZIi6dm
UJ73Teary+Z61l/FCQ==
`pragma protect end_protected
