// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
OotDWzWCDerGobDn9Tqa7ogoSWkp5vo093Mdv8DFAzu6dCq6EPbi8x2HTwUlks5wyOfdeodgkCwP
OMxhD7Bct1Y27c5mX18Q5THWU2nHLaMjo+gPxxJHn4YRetkHKRFBIROjVbUihgJJqoa4E5/RVcQ3
0CfXOBGarW3W6/4BOuns4ymeF5SFYPRjyuhn3xPkC9+FmMvd5MoO4lHJ2a6w98rIWMrcK3xoloZw
W+J3vouBzZIMFXPo8a7qL88+vjFpgdlpNKInG6EH90tpuE6TVgo//stlS1S22ZBf+YFLLSo871sV
nYtnrz0c2ldMvdePEn312QxcSDa6myOPWkJBJA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
xUUyJ3YFvxYfpP3E1ZN+VWd6i/lDmqRoPt0ZlczGQtTxo6VzF8VOEv9zDUDto7tOPsxowkDUgBRE
k3Hn5+9aF7ziZfQUajOtKfs8SnKLY7UsAzoGfC1Fr670RoOwQ0/Ahe5F5T3e8uOSY8lMyelwETUm
708xRAHT3OMG5iYRjZN0wUSZ5lXm+yu6KAvJ6s34aT614VD/7BgKTu5TfNxPrjz2+qJWo5vUvRa7
wiL5Ut0KgRIqbYDAJfzRNKWIleWQQegFylr9jv53jZS8CSJlO3HQFCmohhWiZRE3GNyfrZ+Mkt29
LA6cR8FPt6YOSqQHxXjXar/Mgb75NUlEsVrbUYSSruD61DmjK793fbzvbDhb0dIs0MTniMZhvR3C
Zj9ByRioTynp3ilrti3/1RPak5X5onFdDG3gJVIYGvJ9KDZxM7lxC5mRA1Qq5cjeiToJBPz5EpNm
R92EcMHFoUnEC2AoFz5n+QUWsVsOCt9zlVN/7E2LtoCeUp/k5nH817/NW61MwOYVtlQsxB2tfB8K
T10Rd7uFGkuBmBLcwwkZ0pm4hqpUNbs0iqTQA8pJ9UJxN3LQIqGblk7+Xlt5JwdbQjsTTfqXmXF1
9AkaMbUUUX0NGVbb4YCUs9iGMdvIl+/ZXnJhs7NvpBQKGgegIC3XaLOoyt76QLKt2dFwBeWEP4ZT
OYKkp6R2CHcz9Q8BAnkbXQiWU8uT/+OgCqW/JP32YospRtw8FsD7oV6Kq4HOr/OvG7C/tQuM5L7j
+OP/QULD5dBu9hckLUtCqBIdz4A4OGLNfcyeKpeRHol5PEubn82RTHahYYJKwjT2M/nu5H+r3ATZ
VVTDiq83V1DGiRnw5fhqtLKuTD4qFMC1q/+ClUFwtaGSQ/0ti7g0hfW2I3DtfMb9Kei1utoH7I0n
tWXLHw8cmX28ef1g3q3JiaA8ppt1iY6zPPb3ZhWWlvjSHcOk5kt4KxgMC/uX10IKeIIyzvqzvn3d
cJXvfFKMe2GdiLj41YC8yQZZ0MxA2Hlt9d/QR4wPCyfvA2Pg0ewuLFQgJ68arUoxqR6/bjyhH21P
Kj9FtT3FGBxcuLunJIT+uy5qqJuvDKggsNDgR9bx0NmmrvoBHgTvA+WsS3m84hOsDmfvxZwTedSi
M1moK3wPZCfxLpCTM7agXa9MEISIyayOaLBzVLopMjZwUwGLe31+sad0/et3s62GGLhIocyFvFL5
lsJlPn+tM2hLlvK1Ja7UliR3gre2u6nKzd/ue+G8HwkEPDiQA2EnnREgeO689CrRWrLoEjsBN5GW
N/sCzr0rlsgI2GkztwME7LDbMcbBAtBhOkCCiZ9yfAtx7+rdynDoXmE5yqNDUs3vsxMxyh2IyfZi
okYfHY/zQS7p8iHknNET+UB0NwiAEy6+pUHR0xm0Okzess2SHFo2YapaWq60XlHE4LnDXexrV4Rd
Py4ClWgXvtpIcz/40kGT8YfmYDOPffSHPyyaj+O0Euv18hV6a5hgUENcSGySv5W2sLJjsWmzBYwt
hCAcP4iISHfm+aGZYrVGWd3/MED0S4NpJo8dnArJgpjsVS14GcYL11VX4BaKD5IHBjuyGmO4IbCK
Skk7jot6HKHkdWBTje0DOtcQuQumKXyA9KGhYMZsoXEsAhIWfFN9OiEASgSWQqPIq06wS86fMctK
WeAT1UKFs0/C0tg8a4ittMGMSHEFiB2k15AWP0RP7+s2rutQJU2G9Qzws3R/BjPXCswYRji4KOwL
gDd14G+OJuK077WbxoQWonTRUQNHjYxmKgLoMiOTXMgzHK2bLX0VB34ZwnRUJyRLk6Dsj/WBhu/M
PmpWIp7w516HloNJlPswHyly8HZuaFVjReaVBVQgxjhr3x7WvIP09Gg6NWwiN6yIi6nY/ZIQHVjm
AK7CS7hsbdCRuENr+CJrNNA4oPOdkiyOwkhnUCKUBBT/Ka2ifkhKxfK41rrGZL1g0+fngv2WBMXB
tGXnB6tC/gFWkTDyc8gn0hNnC+v8S9OUU6SlkHKML8DMNAz/UFcZM+kQZxUgvJnJ/DS/VU8MjvuY
sqXPAeLI+7pci+2tFpXa8GUbx0yMkWxswWUZjykE6EdftUmEj5ci9fJ6TZSTCTJMJC0x/WFWdfDr
z6tMUTKz0oD0yYr+xxwAKAnSk0PZ6PeUzwAJJIZ35TwTW8vZM6KToJgOPUtSjAXCmvJioMuBUhcT
vAxI3JhuA+TBWSYqlqEgwwVDitm/26hQAsWUU1U/zdwQp12sThfTrROZu+h8t9t0YBHxiMBhMxdH
12LyD+loBxkuqmUPEU3RWkbQZUDhqj7s90c89slzpIFmrrxb22+KY2Lg3+9l0yGsMR9gSWCHmVb7
bDJKGrLfzc8jVQSI+CY0jZppmptsbHonmLG9HRoaEp4stIi2mJ+SGNBlfPk5jXA27bta2vSP2kU7
h9JcE0766SW4kvJ6d8gb0DVN/eO90PQEB26wTZHtEqUcpJDpmVJzl7Toj0hg/Y5hShg2pHPm13rW
zpN24cPwkK4ORoUiMRLGCBawr5WlgMAuYWFFXvn2aARZmupBpEgCMKQPXjplKTsEa7LGIiRL89CK
mg1MHIwY6hyVgfCs0nmmCAwNfUtrMksVyYYPFB/XwMsh6iePs63n/jSrNCjS2VgBHr4b5+7kZif7
ZrSW5ztDdo9O7ulV7WVFULhEGoXAnhJD/CGU73mOHSdxCTkgch5qVKoUsGuzgQeLdX7mYQFMhnuS
GTmZGvMSxW7K5syYzH7SkeK+nTO8PDkQpJ69g/QKAeS7Y7kczFMl43mIS4Bw4cUHgKWWuMoB8DTb
ZsQz+3zlGQpmSQTA0PkyxunkIWe9TblJYYvNAB6zv0K/d6+5YBoh6n21GcV1Ln38H6rw9ExBLbfU
GvafTxBf6ys0joXHLgpjcKKeBcO/JnqQECuLo1K8iJrD9lNBs7NEhzo2dqepFLTnKCOd4TkjGM2P
YVb/k38iDIcB62Q8Jd1DpV4e0LhFDLGye6gco4Uqhe6V52E7R9t0JU89G0cXbkzG3D2Q3ArLYqVF
yUGs05RuDrr6te06Yhm2CnpgmIEI2tZJ00LVGhfaun7MCyZUv2Cy7B7KRVtZ82VDkrsDuq7a+ErU
ueC71sUqer26YGTOOcEfB4IVAq07+Kabe4XazaTPigxTH5u2al57ZwDGzXlWW53C1abW67LnLFcG
hrWl+faPu++4Sg7w4HMEBIxIFRIVlN0m5xHsFFz/CJKfJPPFsuF5RHMpXweqkgq8821sY+hPpOf7
G+nuW+4m1a/bIPn/sXwkULdrIjK86m168Mh6GR9cEvCdglFvxyuo2gmd3a2okuiHa5FsWYTOCkJ2
OCyjXgqHwA5bUWNHJJUQBWHIWmz/WFfg+7sUzq7r4ZLmXowVewKfjpaHx5O1YXJ+67vbvyMz+31N
DhQTBa1i2gN2+pP8T4Hvxx9G4N/4qKvXDci608LceYegdvHOVWpNugDt+cZXvGN5pryZwKOpNTbm
7eJxZWOyZRMAegOZ50KLgGXHRUYdQYCGX6XgDJ4Sw5u13hrGVSW5m0rsR/mnDFFWBh0yizj5hY4x
yTKfLI2KVP18JnnsjdAc2/S7vX5OLryaVteU+DlIJlD30J3AwTOVqp7UudEsAv+d7VVBjtx5r2p3
DvpS4MePAj2HFzlRBFBMhXpFJJ/aRVhJ+yRa57GVUEjzfd3R0+0IE9CMsq7ET1unpdvAWXNH8qwz
nqRam7Rn28ogMYO9T5zKDstLuXx0de9VMBSsSCPWbvgfIqxN69+yBS3ITR9Af4lGdAvrxySzv6du
G2kwgaVRqXHcf6k9uQk6D1wKNYKyEBhAm+TGs8cSMXFHZu5troyYOz1YE9ELC1FehJGxupEDCuLG
GLeBNdRV0wRB0hwHWR/DClI7jW/SrxoXjQgS8pAiTPYuWA8JLNyugxCLJeA2lf25KtNuqqVnjzgm
YMzw7s5jcKf4MDMRBs2k8V7nadK9Keg82ZRLlrhOtatSn0r83AQQwbpoMrZ8iEYHZiwbS/1jBSf0
3HHRjUIEz9uxc4nMhMrjdghR8f909ANW9bwZsJkELv37Or6YxHpOTExkQPGqM9QG/zu2Uyawc1j0
HKHIspV4XjoWnMCoAXVXpKNbtorjOGeZE1YkQ/Fb7fqGgUlSHCQ7bvVZPTzYJ2HmI0Poegvbmfav
IsLBQlwmLO8SxK7EKmzS5l/VwuxDA2vkn3w1NQUurVZDRCQLa4NP639zp9s26z2EzrFVVJDgZXot
7kYEqvmf1vOEzOTMiituEqCxaSfvdHMBBK+YR6bKmeVnkSQIPzlkmWLXxAO85DJp7A96RtEOTeqK
4iIQayl8IMndxvZFrXWUM83gQChlEaJxrczcoAYZgIgENXWKUtdazUjkbUSCW+MMBMjzRRA2aOAn
Bk5g5HX7tih0rHHGXWsLWQ3s+Z/UmCURYU8p0XSpgOHD59EmrgPWo3znHh2IDZUe/1CWIRTa0tmy
BZoAQUvcsoR7ARJxfzV/r8L+Sd4CsewBLpfHmiipsneb1RGoxWPb3EKGZfPVSjmrUf/+ReCcbHQf
uXOfVyXht+4yG4r62WvdkOtmKEQYqxju/geD4FFPA6ifqqZLOQw9CUt5tMzV5z3CjPyxZgf7eosi
nyI/9RH5kd+nAucjuVaOoyEu9JG0zHTIjM+mPhOQ3YipAg3gqGUqM9Wa1gW4PWP17HhFiXlkk9dM
hiY4gWmLvHZzTwZM86g9eVB92A61teAFHyo9T6tostaqUOFuLTqD+GgKhPDbYYfAE+OWQF5MoV3T
+gF+lsy3Zep0SRLs8vFcgxKfGF8vdy8N6MC6cQFEaYsTej/RLonWgVg7ti8MBbSQkNMKFywAQDsE
TpEpT3wQ2nFthhGDLf8xaFRetotDbpfzneg9/iAV5ceC6j+d6DwWXTh+wnKleTmWw/Zt3+6VZxnx
9g3ppLbieiX26gtqVWluphqIOf9C0DpQWW2YUNwNqx0gbqhTUEPBQ6UqjZU4Nxcruv4XNTvVIqhz
PiHR28efILdE/p9Y1muNEGfhQ0Hf51k4LHekLTPvu6gPiVBLQ/PxQ+JrjmA20iLLTRj1t8tJ/bHH
Sz6lFzEAZGLwDeN4SA8e2Vmbpbzd6FkF48QtTY+nfMgBlUio0T3VDQSNQ4dxvFxftwibW0hiJPxx
LWCDdU3M/4cXW+e6L+0VmztgH+vKfApJXotFUgRenRTkm4r1oRCLktybkDb5aZz+AlEg3EJikb6/
imUoqJq6zaQqIV483qhDUcqDONTZS+4L16Tk4FkD5pMpoIkhccrH+AwaEzZlCtgDyDcoC5m4igb1
9SLMCUqWZBYK/6eM9kMqg90zGV9wnMwencd+M3WEtZfegmr2q51Y0T0PSsNEHE01zdkS186w0kUr
cT02/EQzAGnM/0PX2RD0Ph6qer0fP8I66S6vzSbfxiQlWapOoQmSryvBkneTVukdveSHpHGCVQ6K
LrKPjIhh4zew9AzkvMDNu0EkBOPkwr7GOVJLxZs4+yPasPnN1+NntPZw+Ef/5RTq5zkLbzvPLnIO
MX7pj3eoNRRD6X6ylUmt0weD4P/wxSYQ0q1w1q7wi/Z0g4j28BLzoMfm5gYM6l3toKPdHKffHpJd
f/XgXU3yoGutZnpNK1uMs5O5OoYJsjNnPhwJcnDXaFNX1nflM/ohhhM3nkiFE//fqXNPgN+wSyE9
HsFJ2QoTiKGNh7ab0s4sRhcBslhVJfwzG5IzXDM/qeij8CPXTxe6omlb9o/gLeZYYMUJvhfM19Ij
iD6nyCQR6htx/1gL2GztWMNB6quo4Bv3glXC7Wtg2dIbhjCEXTq2YRrHLoLOBYk4aE9XskGBp6qQ
jyRPow9ujh+vProePxQ3t95l/90KaexRfHX33WoCJKWe6HW0bxdEWnXBxH3WqWGgrTfjhPQeeE5F
1E50ohNBKO6yzLeIOzsSK0qTr7hG80re47Q9LtoH91UvldHffWJYN2MhjnaUA2swKg2H6RTO4Wic
Ydv0xtRoDHjzyrpULi0YkDcsRTQyqbpwIdD/m2Irwo3yNvxtHI18MHKW6lhMgBLXgUq1pD92Ld8V
L27Q00j14exKHb/nDU4LZdNue0ONiWKHH4BxUxNE66tE2Dw6vTYGWpNhTtmsGv3sXtgEk2wvpL6+
qe0gF5kGiPaUc3VKUjF1JeMUT944HPEpsLgtXRYhBg77ZXQ8e6IWHk99SdKvDrFxS/p3txno3mNe
X2EVozUWwnB7tzO3FhuVk5nluEBgxUu1jEzoorWJgLKCz7wok//2P+PcEIGwPukf5Vx7lTp4yNFH
VMKB+BE/9+vQkcc7RVlidm6W7DBZGfxsA/jA5rNdXHVblKepKfoSDHPXm8f+WLWtblkjd1gmui7b
qlKPLRaKZJ4bT6kuQcf0QRda/aWzmdLcMF1WqmTqH/wrzGoLn/irsXpvwn993TdyhLy5wmnOJ9yd
EYy08rRYUUyS98bK3bDGnoSI/+JsstPuH5qjq+4ZzQDHgfxVyLZqvSVgvassLR4YV4aITWJ+m97m
XSptTLtjU8tRpVLIRP2bk2fovHlm4taADS0L9TGk8LFrIysWzDFlxy2QeAc7qdpwyLElx8JguFyR
WaX4IehX//X1z21x+BiFTbKxiMkZpspf1Cdd4m6tt0jTlVBoeGCgVN8JwC4nDtdth07uYFiSVC/5
TbdmWYxZ6FqjpAFi/tka6s99Vm8wgpMcbWzDLkaj8oXkp5pw9/Uex8wkEIo7rJ53IZkSxQCmhPPL
U52eUqV3xJvg7SnM5HkS7ON7x1CAAR5deKCOSGXJwCkR+pD9PnAvaznK2NHkSmmzD56NSzHNfz89
PR5dtqyhHJrKT7HKgBGarHSWKHwM82YDJtYQFubZ2NmUHtWXoAUeu3uaW7qXnRxwUe/pDpBlaYOl
Q6VfciKeZan+EQhK6H2i83yFx96VPaF/zgkteQjACk4twn0ainxUEVR0Jg3eVwTMCLrJ2eki6Gpb
FkttF1vgKTpYPYSNRZIN/lxvIQ8KUK4097w62TIt2J1Jc0C6oYYyVem0y0B1iP8UC9qXsJsbMTNU
FVq41fXy/artJO/KV3bM9AvQ+7mjKmaWfuzZ4sTHSKgMN6J453Twt4m3Faze2zRswo3ZeC+8q7lL
rIFIR1BMo9NJypx0yGbohQwIvxgi35NhV9F//tf0ejREuslkkXIleK/QD0AnVwCjk9BWiJ+Arroc
2eDfCFqUNYV4VhplyxiU1VrJLTZXGOPQ2YSEv9qXMn/B/krjlOZRUNKV7WpbTJOcfjKGmSINDXBE
UsLL5gKASJWNUvZN2ETi4rCkuZCd8b0Uy3W7MMCVHwFAk6x9nKb+JeF03sp1fNWLT22Gbbb7iDzh
7vPmlBNgVf1pfvNGiFXoC+5o2iTiVJsy4SyIg7qKUc/tYSMDkP2D77tHVvhM7oeEVWu2aMCbBS0s
KjBT540prpxWQ0VhvcjqwrKLdxxLtF2J22bEk0MRbUnKDxKvMPl3knbZm4+pOdNCGghw0lJ8J6dE
KF3t1BQdreQD0B9lLEUw+1s+ZxrYTs+MbQXk8I46iqMWsEgWnryjmiZPBuzZ02j5gsL1XWmcpNt5
w4JsGPJjUugiNJqKN1ZCvLhGtS8N6IlZk8VSMwJ1vNbXR3z91Q6oqpgXOD8FmptyM8UybkBkJuqZ
XZ4wP4ZHRpkxGEzXNAUu3R/ijA1AJYwfTynnyNg9xo8JmU2+CHMn3lVdI5Sgqb/79In7zaZO5ZH+
s9FJpgZ1fODZ/S4CvFg50Is7pbzUWJLAJs/1a7GYrQbBLQZL80IM8IGDFuja0RunZuaFH/RFTnIZ
JLM6RxbyRbP0liPiZLTf0glQkNRTyO1AysUG6JFSeYUSbUrv85RVifUhlmlde7+kAjJxfygnle0/
UDPw0dwTQtzC+Hqr4OT/lUePSVMmiyd3Ra14Kk0KhF2oaeg7443HsSi5RMlESfTjLxG8M3z5fDw2
TZbObPjxvH41g6UWr2L+FHT1JHQWYDwCmR093a5HV6eInkVud4G3aQT2rHPjRr9TVonSVwqzOS33
/Kd9x79gh5/3VtXXyIwi9Zt4yujYQm/+9MpOyNa/lzvgZ7KGAHvWwyywZZkK+tUfl2hYH9JlTEQJ
gPulV0p82d3jugBZABDjdWI3uh7zSBdxXZQBePtG6xv7iCKi2dvZji5FUx6lUIxogQKmNXX9ue+a
vX0AbOS3XTWLuDcmSdgm77Y0QCL6VHWvX+YvpvQm2dW9n8Vhrqf2h/KQsv7G3itJr2SZL5U0pyVh
zU8b4gOBrQn0yABrzIy/8bnXSvKlDA1Y4ltiVMvBsDjRzXez072caMPSLed093UbVp/E+gIVqkiM
9AWEFGPIy5H9W+Vad7CEInajQWiViDPO2SvAklL9eWxIccI4AKmyWMs4ginJSNYwymhPyRA62Qz4
6nFLTjuiwTrzquuc7xmavzSHmpt/kydVgPoLigKtYcL/D4hWjB35c0OouXFWi6j+dN4NJEoFCPB2
jf94LRKBGuYVxHoDgQd8OW5XjImQF1oKxCsW1D+Gk6mS8aH0qAOKyZzZnjnnJLLmRy9TkFof+sjY
nKxEt5TFrIYnmKnfu55Vxtuw8FfUK8aBfST5KUEcRgE0yV/OA2Inh2cKuzgN6vnJf+o0Mi8hr6lA
EuwUV2AN5oGRfcX56tooDZVug5vc5BMUdOwm8iFkHiBjosAtvSj/+/ToKERLYxaKsIs1Nl7cL7Zf
B3wn0n+JSURtO8U0tgBrQpU1lazWlW0T1VgJd9bmk4IQhyhZAO9yTBRcTVH7CB6FhHUoPRPy+oPG
C5O9rNpCqPmnk63e/Rj/ZpBgfNEZc+7eYLdA9zNtrQknRNTTVQh2LRX2GrCG9GA7d7zrWZidyYJQ
ToMkgLqIpEpdxhgvDD2eReSDH+ZknH3e9gGoF6KaP8O+0VT8Zp/gEAc7vh5ZODfHfex+DsUdJmpe
T/Jir7u5LemIOl2MEOfRL97QYsaiO7IEyGG5VvlVtH0C6F+wfBvWaKptl7M9CaGciPs4mgpX3dNi
PkCkrBMCBxdnfMhH+eShOF72aPJG/7vOnbyCvUg7QPaaTizW5gCGz4EX7DT64aZVb8Ld7IbFE3HU
RYq8H/sU55lQLagOsgROT/BEKXGea60gA2oVWeIp+aIA6nu25E42KkvRfmlB9Z+/vsNCCp5F7HnX
5aOFviWIXjUmXcemlwosVas6iXYwzznGcG5cyy/Rw6d/S6Ra+aq4M4ReK/L9r/XwcD8uoFYRr79t
NYLt1iEfOe0CNAp4McErLsRLnquVvoUqlQjJcClixj20VxBjMvIixQRNTZsmejwpjJYRDc6iTKxp
pADHVAWfOz9gXMEZw7CfNDzvPT4kCat/IX9oViBTagXVH5OBc2akTJKdaJFTF4MMTmPRiKEwB77p
2gGld1m+n9PlNWHudQGbgMl+wxWIsh8IfoXGmoJ3Eiwm3oiSo/iU7mzfg+pDXFmpj5xIW+NT+BeO
uZRtIOHZqrrFdrTBJj3M+i3CEdPENFoIneK9Mk/+nPR67XLmWeIufAgGwRTiHhY5pEJ2KXlqPbtB
hSbsQae4SbUK2n4r+Uu9eDk4o5cYmVMhXsWGHmFHqDpfF3QtNUH0rMR1iXMDxY03AKyAvbeVRSZb
e2xw15XgGLr/sCLPHSgZ4y4aFZcPF0GtMvXz6TArxfJhHfsEAW1aF0gex/JBztC0XfqTyBcagaWS
3XlQDm6GUPWhCoSYsF57QmVFYdmWPZsUGhb/GWuGsmMro+I/fXwZlOtOMRDPoA05QcmFTCM0fXQ4
jWPob3xSoF9nRCxXaFep3QiZ0QgBUJlb5cjEtWoyBEy5K2KeleDtaelSUI+AdlOFIXk3jywpISwI
6lWu2LYcJVBYhHNeRSEbegTICBcrxFtnk1TpPsrYbIk1757KUeL9pM/Rq9TmsIcXh3D4vWuPqYip
5pbLnoUiyOTlH/Ij0C6KhLL7kGQzr2h4fMZ+M5+DvgGrR7sRC5kCItnrrrDnm4/cMMtSwWN2J9IW
lyF67ojSEQSX4h2fV6f88bXmu8TfTzfQwqHeUeQBCoWVzF237Dse7yyjNcBMQdBlTu1qUFBFMHtN
SM/e23Y68b52VY+mqRHwoaQRD9BVtjFOpBRRJK5bejx68g8YazTRx60WpboxH9dc24tyNVibajsi
IKu/4AaA8JgYMzxOeecuTsUL+VT0pd5wAmHiwR+We4YtyU7lMnk4CSryOHpJat9x9s5CAKJtKSC/
319ODjW8ngw5wOn4roIXvJrPoN117MUCVbdDo621EbIKvJKZnCZU97uoearG+BygxHrO3gvenEDR
Oefwm/oM+4ku93vU2nbaIqJ9B9S3+gogjQgbIxA6ALOUai1wLlj7JcOx9T5pHINdHIKdVL1pLYpH
FBs02DPjVSeYEso9SzthZZquFvsmGhSCcUvsZvC3j1FgJTxWfQ5+FePA1eaLnxzyOz6PbVmLE/36
8g0/etoY2v2YrYOsX8uwGxqV32NEyruV2P0WVJ7Mq4nQDqs8pphSNwDIyN/TZohujbxYq8fUdISL
VSqHbVsZrjbYbboKEZst962ePsbVaAHUe0Ej7u//qGZpURvsmZyu38JhzHGwZpnMHsmQ/5QwivBm
3U6ht5lLrDZ6Re436BWSEfm9R1xkDhpc2hdrxj3Jgz/fR9YTzpZxt/aW5ufyVboKUZg6SmKf9WEy
IsoaAiN3DTThRUUcZKJ0JY0dBzbCZ+Qhra+ygTuWUcLq3EzbrTOnP+d0BFBQGYReY2fGgp4h5L16
jxY38ttVhHpGLylVfLtofLX1UANOFMw1VUMtVsgeN08+BY5BcrFG/0UuTp0SIacdOuyImHrrow6i
oQu0J8ecJmAHe9nf7VW038r2jEf0W/rF1FYHANejiAM2NFm2r8vwZWQed6LkleOsf/XUmoT8/jfe
aTLqdPVDk2HaeYBtgTr88zFiRPYzWk58Fe3JNxVaDl4vrKSoqM+mr1eHKf9d5BAeGd29tU331LTF
8kS7YmIXHQ6qtcD3weWd+GS7/TtoyZ4y8mI/PUy5qi829LjmJ2YPlVPHabaRsjrNall8aECnllDZ
SrmkbWUuMW1oTUud7X17mxLJGHwBUf3Rsp9Tei5RUytW06aYjE+Pcyes3HutuFla1l8RZJw4FQI/
gYZaDEnA1ReyZsG3zojhpQ95v/qvo08vCKrsIb0wGfALTAgxjWZCVLcnqaOQg7fDhJSmotda/qKv
uic1prjn7wK3dhzW5Hzy8Zwl4TYibV9yvSxO/G2DDL/NnQ2plNFJDFbNDvTb9ETejdLWeftc3N8D
L3XAAyxaNpT1gcRcjSp3/0vY/iMYvJ+k0dZ5b4QENJd57pBNVBk76bi94p7ylaVdqSsRbXOugxRA
bwhzSPWibjK8lkKENVoFv9FQFUUW0N5DsZTjQ6kNU+p9CLbr13TZPzNtskfQ2+B3oeu1m8CWst+q
MEqyvMyRW/KEiQPKWr2BmWJ+qy6ggWOoqgVCredB31WN/hTnVb5OCrvFPTA3MDj0D/Awb4B7A9bq
R6cNYdrgOAvp20n6lJvaZuiu4Jco8v9qD9rgmYupoEdQugCxQDVZf3ICBOnVtoTuowwOz3+/PHex
yYgrKFpyuaLM+5gKNAt6i5BV/xXEr+vYijYMGOOzzUlWk6chraJN+i0OdtexXWNZC3O8laRydfFM
CWPS70sryjgVa3Zz5iRtfILRVrtTaMp2HJixwM1P4qmEbz4CVPPo7i8Y6g3szdPNGHBpp8vWSTVb
R0JM1c2f7aCATAb3Yn3OUXWtUJ7HLbzVckmqWf3yka6LFXNAewBHBwFB5ey/+Tj3JzOSrInvc42H
JXtp4aHcOmrUC/YhOTqRDVj0JbGU4KTHw/3kaO0LQJ34Bogxh7oaM5vRZDA2/lgnbsz5IHfAYrqx
hdksvH6PU3bJax259/xIulDx3Okr4bdz0Se5qP45PYPYbZoK4DNgy7VEMDZBJJO53g943Mx1u7B3
BLCVftL/Y3x80T4o+OrVDWGDBC19NHQdC8O+L2MkrZVqcWbOrrZIpF1kMbZ4LBPTtmC9VhA9E8NC
sBo6roVCarL6IlZSE1XmlFhkW7xBfqTwlM+aG7XBaUF98EU46jq5IBBixGo/fLNh0ciM6kF6vWLL
p1njEX3CrZSlQtQ7bATN+q4AfM51RP67DQh/HAiPVOmbTNW7Uqb7PavlPhl/p7ve6j5ROJR4n3/w
X4IH3Chgw6ow77gxdvlAZjsq8UZt5iqvYNm0WQoFEdHvcsDYQsIkyeHLt6GZTL0LxaBI1f+wKCO/
4dffzglN6M71LWULAIUgY80nz6midm2Qf799ZGkGeOfXFZx1btBXegH6nMsffokAwZPtDqNf2VTT
9VDomY2jW24k6dxVeF88D6+HzieI8/w4MFvdX6uxG5PAhNdepBrQbv0TADOkYElJ3N7AJq5Oky8c
YE6RkvwGjlxI1MruTN24NVsHRdIpa0IyX6aHplJmAoXY6JCIeJDzifo93dD/+kfvQ7YPXT5Q3BrF
m2E3xDf5Zc1sQOH8FoQrdp4VcRryry/0JwJcRuxA0uuucDYKi8ZGyi7a5ZPngytQFr3BhZiG2wiZ
0Efsh/mXrKtGBGwl7m0Y2xr6LDgh0i1S76sueS+qUiGMOkzIbOS+1KHHDig7vAKbtyZlM5cQs9hB
/tJRbV55QoPEiWvk/DgCq9qwC1lnr8/1KCNfdHKR4/2s+8tJ3gyhzUPbSN8uTvIvdzEkOV1ib13V
cvOiwdBsWcwYZNC6Wy743Vj/mF7SRaXiLgXSbz7b4yy8dsrTny9QVN649Yua68gvBKHkwUob+bhU
kvwicRftkcItr38rslB0AnUOfs+oHScOkQ0O9E+otAHn4mZOeK3lLFILdpWsvrBiGtiZ+Uok77pF
DjdlbiFg+9AxHjCK7nP1r8xEbWA2yhZ8F3yKZjmex/DfMVTaUys/C20an6+zJHEOTs8N6eZ+AAtm
3Yzt/IuUPswV77cvzxorgVlgc5YNXQv7/a7czbZQ/shx0EJO3JnhR3omw84+x9PjhI0SCTW3/1pj
fHnl0ZHbMz3YVq4wQ2aukHmdjYQ7BKQXFereBFS1R8EyxiC9JRUgP5tfXoVgxDjYNk5SEJe9Np34
tSsA98MRh34dRosnzgEyVdSGL1LiS57gMkuq7gjkYrralbiJmE/nAc9lmODul8Mr27Vh7c7z7U/N
IVMGFWNLxg1W1IpLTB2AwyBn8pKOckyV/pQCzuPqqA9tlIgfKC3Q793C7zNajB0MXiChEHeVYFjU
Xdrb2ocUdLebpQquBPOJW3RsEIXOANCzAQ5v7I9+9vdhEQ86nNak/1jod3ObDE2lHZyV3Z8zVrhD
VqMF2dsHSUXuzJCjACCd/JhJ0eKy/d/6TxOns8X2wTh//64024iyar7JoT/g3yYJHm1qdGQHa3qF
o5bdS5qjimbDx9fyXiestFp9aRUvSNdq1dwbvvj7DrdGK0GBNTpMUSZt/tjatC/4NKfEgGdh7Gfb
IG/T3tsJTYfXqUmLIMw7mkCYu33birxIHOSgurcAPnxfGyd+H/Mb+DVCmEJkmiCGU3d8oJIUV8gD
0UxwBTZNC3JQJhBu9/TrhOXKfq68hoSGohggalWfzKry9H3qj66I6viWatk26x39VgzUBiv618wr
7WBNj1tWsklNOUzH3V07rfrDTsBr7adhU/KXXD70bGRK807yNSWihh2nKMT4MlrOdMx9EE1QHFVz
wHft/2fEjnlai+yrkSeoDbhwMQbIT+n5W+WYrSKP2R2lcslhG2fa8s+1bxIEz3JyCxa5u4nr42/d
NUdQ/gFm2RfdXJGsC9fIkOwD47xp/DfSVamkunABAFki1MSczvySPutGllagH2B6pHWNbz4ccD0U
gkTXJP3LO4lk4KV7n8zvgitKsLdj4bWE0fhs4LSrjg+QOqK+jun2wVXLpom/uJMi9HwJSmmNWy3g
x5MbvzdfCzAtVUpUsLbwqkcUWfwK/iRt7HvuJrwFqJXPbh7UQ1/gCOku/ZnxJ1Ov1y2/Bsr7q4Wn
m4xj0MkIUFwBeA5dXDZsILmzPMDzZbtprnxR80fE6NpzY2wUsNzGZfem37dmF1WQJEr7nD4/1EC+
mdq+VJ0kJnkLFkKVdMdDdsqcRakDDiT0LU+DyN7dXp7EoYYejT6eVC7GXQIqKCrbOTKydRjkGwPJ
/oMUkMe2ZJrKTsl0SZNlAF1tslhsdbbPEw03GARpr9X0esUVQ/sGs3rUQ2DBFl+Vu1PwjWB3DrW7
2jxG1dOPetghbmqrLKhpA9yM7n4CCviAoKI8l6MKDF4QaWr15/52Z3CVBanXDCX8KP+2dmienHDX
sYcGr9xozFs8IE41jH/eFQVZSLr+o7uM9F5p1M09bGQYqr1I/N5iDFICFbr4i4Z3JUZ6ABvb7Ri4
n9gkw3+viq3V1JHGGeohMhwfQhp59Q0UajyK2isn7AT+Qm1z2Hsn+CUOrwu0RYoTxdUqyB1NWhOJ
YhkMWWZWE9y+lB8KrspftvgUiLJkw/8978HuwuqobyEoTb8EA7ehQSUHUoYeebEgyiqJhPu4MnD+
8voLpUY2/NFHqd740Zig+lIDKu3feFPUpR0dh3u06tKp92k48OoCDuxUwrKMK4ItPpWqkbqKGrSz
HUVpEqTSfBtPM0010FAcMP053hUkuZ/MUvVYyTPKhE1Ah7IhDAzM/Z6zCUZfD8WKD9DyP1hnCiHB
A/j+7sfCTzEMTnaKVipbToEgs6uREJG8W/TEshyXA2t/1bGADgsmNMyC/IMqeWn2M5t67Z9rtkHg
qjnPzv3J9isjZbmtYHydt13V+NgmXr9CQ2i9R4E5dMvZO1pyzU6/hBulNSAX8d4uu/Xeu94ut/IT
erC28Bq59kDqFc29k/TtCjfSpHw4WAIrl+XXm5a+ORflDh4CNTTkV4+3QxE6eFCUg+rb4vMyvR0n
YYbAsIBIN7uDfVjPSCfOvj7bB9KMGNFx5/V6VTnVypvyeNRqSSTFU/T2uxa0e72vfow9ZRKco888
nHC1v+iJmqD5tV45sYWxqXpizR/kHXlWMtHOYFOKPAl8cgmJYBIpDReZLfzpcuUaqVvUuo09RIoX
ZMbuGzyLUDSOf0PpU7K7bPqqJoTLDGFzzYLvxFq226LYbzkHu+bGNN0RAPar2Heaw7D47oUHyldY
1fVW5N2o7+foxAfZorHn8pEHnudKuxAh751fFhYFJp15Gqrx872RC7sh8lYVGGAoNzXBmJAUERH2
xpQTIkawxGturKQCo8H/4LgOHJGPlXN5IxyH2bZ15jijzf2F+Is0cUPL9msWVraRrlq5s5J9ABn+
bEBJ79ysSZuI4tKNfVN8R4wdqdGS+sMv8P2Zu7Xfk6RJx6SpmvjNQmCOZzdsx4yXjgfDmq7kvSzf
vPy7jETpK43I9Bx8isp5LfjRr7L4wk0ydkxeKW7dePjNt5vGNicwave7dsnTe2imJLxob3Mme+Zx
kbZuAqwcfZ6GkK3/BvELCcrkq/QUri8Fk7DkWsAkkEu2ir97M4OYu5SsWRBpvs4Xnn/G6nCTck/M
cnNJsuptMKxah9x546BIsr7YGbcMrQYyFYb2iqB4KK45VmM38fo/6GM7faifb4Dmmwv5RZNYlkBi
4bXZW6NOrgjPRio/tlsKM6Y73pPVQvPkCWKW3HqNoclCpkzGTuUQFoOVBHM/uG2n6dpx1FJ2BzkI
diopJ2btzdxbJlgMKd7AFHPYYE1ws7FgNBOD/lJqgVNroNwMejITAZJaSCXGjYaWkhDB68YigzdY
8/1aeS2sRa5z0yHz/Kc5JI7qfCpwWOLzER0sdDFjfjkvoT01rLvpo3wx7ASBYdsb+WXJmC6YeQ21
G5Xq9xSf5Q4+4QDlZkqZ6L9Uccpw5EeKa8KWJcmty2l7Ti/mFtV+fZeTQ4yED76azZgeGi2P62i2
JLoDx6hqg8qVBQ0cbh57S4BH7NZ7jYD7em0RsECMz0lX8undC2DYYkQ9GA3IgLH9MW7uC7qa3dFw
WXic83vrI7l5w/rBSHuhhUU4kQCUXE5OlhL/Ve1VLjBXgmwPKmpivqruNkU0865OQ/Rbh0DVse53
CZtCn5WJZTHac/plWaxCXYxtZplsKOtfkp2yuhKp3gkQSNj+tcevJX0zGgxpTE1JcnAcNlxTG2Nq
COlGBec62EUmYYLp/qr7F7fbpISGppdhhDsuMwVXbfX9FpTQ7j5t4A8bBoG4f7oaeSxwROzHm9kP
sHalKYIRuj9J47aEIBztGnSu5Z0Wxqxp/OTKfmTsNr09CRAsAkHzZKXZUD+P3745vondNKDY3lDL
4B00qPfNedS0CvC/+MiDllYNkfhtAqulYfCMPkte1KNgVk6VjGpR2LN+CEE0S6LAozLyuX8BgevU
DNhxD7ga+2xw8noMtuy0pHXsz+4W4dTiWVvIeQT39M/7wRSjsJZDX453JwPB6FeDrkVJAGi9h/90
hDs7+981SC2r+emozu9ng1w/CniGy7EB4DkKAgjJ1yvEXgvicWYKi2D7mrTawDxJ+mVNgGKYVhGO
4IIYMuvB+U1Fkz02t6Hf6TAzfYxWjlO4UywenWURfr9ab5lLJgTXqUZUXJLLFiIJw9avvJO9t4K4
00nyv1u1//Gdli/hH/TiyP0NxMTbGeqPu6Qnjr7xxYvRL8p2LhlrmzdAOoDwp3x8UI1efK8wQBwi
v3HcUj6BY3zTKDUQGoaV/oFb+eucR6V6pCQPj9m1sN6vpw/2MCd8Bo1CdT8QIiMkXyrm+wNcQUXI
YHhKPUr4OKbKu/XRoq50BY7I7Ssr+mNJnBvShSvnssLRz27qTm0pDPPWDSqTL+/ja1xe9LUR4BD7
KJ4sHP0kvNIVq/c3wPjKX54+oPsdKUIfT4NRXBh5v45mmk4ox05HmD5zxJqywnwpOkf5Wf+vA92D
KgAjf3InAX8J34GD+TIekUi6Q6AsRLvQyq0Wqt9MlnAmld+l8eBnxknSTa/gzbq0Dl8dc/hPdsms
XTFKjZRd7i4JGYGn+v4J2p6pznv/mXz5eiuhUAJwGe1l+D3L1cD8ItzKANFwp5k8nZZFaSdc27Og
Bp6uTV7wDrcCRHaiiwS57yR1zvn3aTyNzIIn3/aY11DvSauII9ZRtJHuYXkmQt36e5tXeJK5grDF
uiM1iAVWyTZP/rNgdp9LE95MC/BexSeuhHsbSEWMTWxUlN9b+GeqxGAXtW0XfZUHEQ1nw1ikF5E8
bOxW57GP1+prqENqLo/2zdxijILCih09LEKoyo7y0bbiH5C4YPHW2HZlYakCcmOq/4EUi/nvTkgu
Huw/YJAf7vmUH2UhbGQd+hMI6VFyqeSS2LSAlG74BcP0IH/Se60+888+pZgf/KDeTVatRt+qKx/U
o4m4yS27yeDmALZChnE45u4meiKFBx3nKglYSVWYUe5fgSxwoicRQJCvvBhSGDO0hle1QqJb8Bx8
dd0XYkRxFwnYDe1yfJgaSbySE1jpYZtIdbb1GfCZPzSB2+KoPUeVWGy4s1HIVsxWGrr02wZis5bi
FjpA5ect/Vn+txTJfameELmQiHYVV/lpGIy6AFqI8/60esi7AjWeOaIHJunHfKxID1eKPO2G5yIO
/1zfPy9cH3cdkKgi28dS9C7mWVvTFn7yUysKKIkFlxIH7Emzq467yz1YLHoSIpCKd8t5kvYIw4Ye
5bP5RYt1CJojdcGmcsrvmOah4kjTicdjfu2z6ZplN6b2l0C8LfgMTncw28KYlldbJPFE6yrVUxeP
Uzm1nkUj6J2oGPtTYTjdIllIUmH9MKoQfT9cfuZrSce246/vs/QaZ2PXXs40i5qCEO+p9xAlFHb0
wlN+ItKeCFqoTz/NumEaOczhq4CDuHBJX5K9koW3r6LJJIdY0VIVAaLG5khNsVeh+9VssvtusKhK
sKdU/yjj/njfm2zix+5+9TlI+Gp8zP/kvhSdj9e6A6tvcprqB/PchiCrzx4A8ZpG5/lU0ipg+nsK
shEUoZnCgIl0lryMmPHcywEKYot8ufS2OteyOIzzJ8yhOHmEp5vDIuDnoTLTw+pqalrJyScwZ/j5
jftpImBWLPG19HEJvDVy0aVGtjVDK2Y3YASZu6n70VrdoFd8NBpqLpuL26EfgH8jklphkF6u7SPn
atjf4U2CfW5fr52RjZDLtKgXMfRAfLLCtMqRwgdtYAZiJxtO8yN78AUJszXzI3qGrfLaJ7sMRFlB
AMELQ5jP+2TMQtDlmx+mR73iVcIuogw3OEqU4qUO5TzNsSAkSvOEECo6dK4jJA9ml7U5eNFiRaMq
YX8hUCprocRDeoucLGJnhp9MlvGNGCeiJAztyj7Kb1R6IkIfPHfabpoYZHI1ousA0peuZLrnd2wL
mAEV0jYm2zekbseoxgTxNseY8TcjUxovShjAeoef8mSbuPEjupNsPN8mqX7cyCimSYaFe4THqXTD
M6xa2uv9h8J0QkcjgTBj66rHY9vjOF1bMG6LOl2VkefIfbR5J3Vb2jyPwLTP9s17JPGofttAetr4
6Zi8j+tDKCVzqDP0z7iG5RjIHd0wfP+GHcmUgz88NUr68e+tIjzZd3ocsrcJId0bPcrk5SNI8TvD
Gz1NWgS4c0GrXfSboT6+frKsEuwwLJCEWgO2gmNs7E8b9ZuIZe7oMLt/dcmZzZ7c+wqp4uP5fhrM
u68Z9+9a4pAireUvbW/oyDXnUOTJK2WdXlGu7syDHJcO3F60s/dwX/0o9ALhMoK9WsYtNLWoDpa2
IX/H2uCm7MfWle3XuGeawtr1LXd/vxdyuA1Z+/wvxQVmpyQYYZQAQsj0VPmYUUTNoiP5FyM51MiQ
D2Sfq+cOAH8kejJxxkIZgO04LeqkSZelEwwvlgbMtEZY6Sr5FTw81HY1IviLCr1MaCxypiUn4kVf
fuO+9vAPPgyMSxhQne+11ImCLTkAywZBoNEnE1kcr0ld5uuT4iw8uokIp/REJBon07zYbU1G1eY0
A5AsrmGSXWjcSxrUp3YGP6V7MqTXFkSKq0IXIZ8hel/rVuy96fFmHA/8gftyV9TYZi5qfIkBQHBi
i+ftgrvW+YpyolmtdOPf6CuhgwjdE1yFmi44h4dQNTIyT6G6JC5UtZupwI9JiI+AjUFFdKswC3uM
XDi1emnWXeuHwTU8voQIzqWOs572SEiFKLuHOGBykP4ErM7xXxvcxNeTJcI9+u+g1kJ1+8Eh7GdZ
2Vqqi3rAtkT8iRcJEFFDUxIU35FvrCRBbT0szT6/SFGnFtBaZcPw/mdT5ZsPVeD423CucstQJwKg
C1ZdTJwOVJGY0pPRo6uJEbFzDg0vgNitzoy3OntIXAv75RzYjyJbvrPug3ZjFsuDpD6fKKG2y3Pv
pIjZcmO0EHDyuwFORSPaSXhOaItkGyBr74wRa3uHeRIm1erRoR7KLaab3YJm4dIudlzLp5lwO4Fz
gwwQJNjB55nsaqWyxTgK3XPvEsPuyCG6Mty2/Oh/Wp6NARQIq+rgUpC1yrjPY5E+qt73098zgJ1v
fq9rPrfOs9KZa1c15rKRW7MY3E/jFyLiyR9cedLMjJS9r3DEWBBc3l6/T/Lozwl1+dDrP/WHQS+P
J5hd58dMnX69ZvFd1pMnkhh13RkT5a+4Ax2FREfngmMyBjfsd+21a0YeqNrmgJeNch0AzZ0F+zpD
AOjmWXdowlNxUI3+izsk4bJI0HN7MemAEbHjChp3BWxEO2JvLRTaJMYtP7wfjLNN+XohZRMFcc5O
8DwHqWFEAadjngGa2e8+Wdjn56VDi4claxNG8o7vuuxXuHZlSffvt4pY905Wdtl7gK36u+GOYwrI
WfZN2TyJemxedKxdRsT7jClYYLuUXZkiUk0fOIBRVEdSzjLeKK3M+JPM6lQSZC7FQ/pb99ri1WZn
9+ov7XxF6ZaksCaCfUj05Fk/eMmIZRUU8NfL+UXobFm7GpNfGWXHwH1fh9eKM9/TjGUcWqhmxI8N
ZeHBpebo5Jx+nefP5X74kngcX2svPlDFfxtlH/yp6ivDJMsY0E+6tFPnlp+2Q+qKRBLPSa9KPsYd
rGCMBn/8EUzjFOvQdP+8okzCyh3ZU1JALLxQ0HELsqhA6UEX/YMDkbS7bN9imNadDIyOMJGhUMV1
4FBA8+5w8D8OVff2UEUsQuaM3+byAAFvegO6y+C81kImLQvVHRTQQe9d+kMwcxPhmyoFSXYQCVdp
Y/UFuItdvlxB+nuYsTj1w5o0pUyzsMMinx06f6wUoy2+21BrTiXF9RWa9mkPxj+K0+HENzNafAlI
50+YWRY+VksYn7VLbdSbvTvjDCGG4Z28aZDX6Iqacv9YNklRQJLlQNL2Ne7TByYcyz3GK8s8GZV1
ipMjxq5nRqHzjhNtuKhvhBG3XR+G17NKnGuIOTjME2EHGuY9IoCOImUX5pB2HT5HrjMALaE2nSFY
7zW7ns0IR7jQ24ldH1gJVMeR96KVvczojr0M9RVcOFrabmLTtoMSWW89wYIIt/RJXrA/aIgqsQCp
Fsc81QCZ/mUBi+I2x62o23zySa1c8bXhxAiqmdLM+WvGVX63NbK2cW6tulePYD82h+QcjvjOudsv
gGekPDQxod6iJewdrTY7CkWTay3h/QyRdXAAAirEBKSmlHfc1lOTnVGi9J4ZEAi31krnNxhRkqOj
kdQTwfueF5iEK6V3VL0SfzVesczOpjuLb3y2r+6QZ8q/t5pTdTIjlc0OV+mQN3c3TKk2Ah3y5BGw
0GwH3z2zGxGMMMck6stwXDAnpnyVLgzC1s0vi05il2AXCG/Dgvbji9SbnJnaFqt6d59wHOvuMn0I
PM3Pz6TYVTsx+kunhvnMYCI5UtADGVtwIA/pV+gDM9jxFS8SwOpnWTginxy33mgId4ViQltjNh+U
Nyoakhp4gNPQg7XeHn7DI6uIfzmqrqHNVaLFif6tcxf6i2pPZcmx7AiRBLvlUUy2hd7sz+Q/p8pQ
LErrCnCI/4iQRjTubZpyvRcLuPFvYkW1FcNvsalYkvYQ/Su5q/wf0Erph5eAhf0AamNa6FZtNzGr
0IBnXi+QA/PzEz1YS1TaFhISU/N5qBRebt7+CCZ/P76M27TT3Wn+uoKiuvmt/VYDsj1SaC7NrZ1y
MHwX1SUvghm6TcUI2/MnglWwL5kz6Tt5f0h8qsxV+0khKekciqjjd2AOIHaUr9U2dJZpeBQTJgYp
FBu/XvWF0BVEkMngRCoiPzYtkkQEZY+4vVpR3fsM2q+/SswXffFevDd91HmZD9GxoeBc7SCsF/U7
kisUTQgN/BK2R072iU0Cr0ozP3LVT7oQrP2fdjtIPayXxLt2kvWdLSsQMnIIBSS6oB8E3t2FeQuG
sY+gDB0kKig+aW7gLbArcsSjtck5gyD+XRm+ZWEjwjPepg8USyz6xcPiJGdkU/0QCFM51QLlNMrI
NUyw2dImsKOP2NGjeCeN9+i6StJJ9wk1bswC0q0A44l8HAuAa38lhYILpYpG02G70RhzrB97cfTq
fjbuLWdTO+oquw25Nn3D50gqmeFFNYNm+I7CzhfOjVQXrrrAol89/mreEfsEh8otw57vXCuYtE2c
/zSacIdmfWBrsta9IaPjww/4y4LaGKlblPILaUbHvu6vKWAJL4ZePzbGeyk7l3+vnrqZjwxT2dtZ
01/0HtEJ0pXs/yHc6FTB9zpticzGrQJGOEj7ALOUX0/IyI1YU8hZL7y4z0GWa9qOfxBLQWDEcQ59
vqxbJMcvzSwaQe6QR41HolewwZYHJbl8uR+oLbKRZ2YSP9piUjhTBTKQbP7QsIQ7NjFYqlavzPPj
pWOGvH/9NXhNtfpYy+Hkc5ItwIQgLJ4RYjEa+E5CW/VjQuQSaSk8ZAXXJZrnZBA1XPA4gCZWF3KV
kheYHdeFTkxmmR5KvDM8y8v3GEjlGTjVO5fUoCCihaUdPlXZd+9Pl+x0+msmo6NGQFR8q2Gd/As8
TY6I8f8tgHpkVjJvv+jcrTJ5t8dGVKEQ2ENR4lIMbj+pUG8dVV+n4fnXu6J0ta4CoAu4lCM0GsZJ
00AEif/1AI+uLL9k38TcisoxiVwyFk7amFIVcgz9QU1UJbWZ17TB+9wcPAiF3KxV7J7y0wMHaxYt
R+2ssyo3kJeA+XZVRJTVGrIO0+w9Yl0l4pAhbuawsOaD7nrPNqVrd0JjizhFDb8kQsEFUBX7jdB4
euv0ZRvNRXb0r3GGqmAu2DBLvKk42mnTrscdwYIVX8wcxrKjEe1RayD+59mSoJWUrDVhtmp/d/HN
cDH30NKnsED4gjlZCp0J5WgE6JaNN1cF3ZLUYQXdvSyUPd1F0Qa/BwH0LS3n0NQlbZcQt90JMd44
TGzD7YHumaSOTeJDKt/CzemSCDswZTmy9zzt86p9hY4VF0S/bAsKZj79vHkxnUxCU15ju+CyoFdJ
8c1Uj7a47lxPNXRJjwm+f1EeVeQNxDAxjNV3pnFHb3XSfR8YRveduseJjGC8Nq73+o6/S9p5sPKk
DcNXM3YLpLuo5AzDXks19KcmzmstQ677qxPdCPgUZuAPp4jzf5r0F4/rKow78Toxxc2him7mNyOe
lfBRZjMx+RzpduvH1/s0oFxVFV6bX/DRLT7e3BoTHXWtvoJoJa8XoJdWw7mE2ItylWMIALqTgfGf
IQ3O5rj11YYSaZT3Mgnao7XBrzl/iVWL8FnTXurtVWpP5L97ds3rwVOxWXRuWcRYgI3dvVE+bvbP
PEzUffOzZA+tAD49PAaS56SbiE2eiqKzBGOec2c2l1fFLmrI6BccUH4YoF9fALouAcTeZWGhyfqv
7qMki6HTKrhLt7rPIMFmiY7b5U1Xtc0ehiZgGPUADaTwZ4p/58OyGg+ymL8sKvBKP5epKx7ijCSU
Ec35FzeAa7dt5b5DiLN1ByEzPJCcIZ1jUCI6UAsvTArIytiW3VlFH34ViqSsAFRViiosmEDwGfcB
be4CO5TDtDJ0y8tFwNMoZeXzlk3kK0K+9pFxBOu3Xq1u6nNmOgg6EYiZwVaUcCfppElchdsLyKd1
iprwy/2KTWQaDWPL+SpvBqrsE+P5BDU6OH5ckbIZMuPHqAorK0I9cHvQMHbpwYxYtZhyxL3dKIC7
goIBvNRst4NI5FK2Q7JNDzo/g+Pj3ZOtVqW90rqW/+d7apRus3ZUXUqOkbQ8PGrkR7HOHEPWT73t
n0Yyqa785JM5Kc1abZQo8jbhhWLd8OitiXz2gv2N7qJThWjsv+tF4hLJROqsus7/5AaXvb2KqCOH
4ua3/UfN08/x+6n1FgSw+bC75ExM9G11TsZr1CJom6ngPVY7/7eOQTaK9EuWFtrBcSY590gZxKRm
foUnVFIz0HTZIODtgXyJk1ExGKsWUzgaRce/9u1RIQEQ/3D1DxVcldbG+JKpCkz5riHXQ0xakJHe
Dk170WmKbw7sk2hy4kGf+8K8qD632cOT0W0VhQD8z7AuRZ7Im865TmeARGz5IRLIXtL/BJ+m/U0F
6TiBilON3CzOSao0Lyg6DaJHMeJ/2ZBO6HfeAkFMZ0ZFhHKjQp6QW4xCXHfXM1C8tQQNC5F19MFY
bWTcKqCGtEBIpm2R8Vsr2eRzWGFymEphKR7EdOWLc57yhoHmKWarO4izzLaWCLvpJsR6h5jFqSa1
Gd8bv20Mzr781+dYqJ0gN068P4exLynA8fARnYYsi552Lt3papk4yG14XobrUEmUAHmpYqHKW0dZ
gxlkVd6wd+T4dUaImZhU7Kzr7YwobAD4PSPxKz4+H9EdegqZEgceDzslSOSNvMyqoNduZOrX9Ymo
AYNonzRRO1NdxrVK3IOK8gwy1X/LXTsFn7ve9I42BgGIHH4h1qvNG4hIzub1dq44RvQ8XuIDqhII
DDwEC2KGTlKQB85GLjItTpu+/NXZBQFaxcRAt+yipMvt1ylOpaSCeQRkQGxMpuSfr3ObQCxa/6Hb
UcIsTonwJfQGB9CEO8m2/tGA1acubnEpFUqu7sxsA5imD3CSiYTld1rl1NIF2+a1HjBkQys3cvdI
GhC2ayQpDM++aarJSCa7uzQREqD6dC9qdGYUjsn+7+3eoiaeQJnqt5zGUVnLLfjHk96SBJLJl172
ltb9RbFNj78IU+2WQ9aU1KwJwMZo01RRxEjQ58ohiPVdQt8iRbAa43vtS4dV1X5CymU4dyvSHdBS
VlqBtKcgMPZ9E+POjFXUm9Rx/+57hLmIFbwDBHRTNhXq9cv4L9P5fXKobeEv0zIjfra30NYwiuyp
3NbBJ+2iIhbxR/081DqGi+KkDVemishFKkve+1AFbLPpfLPGBHLqnO/iZNJOC8aGPKv/QnE4PhcA
dlQT8qXaIFh03TQlOmIMaqbyRcnxBaVoEAQkR8LSgo9HZswEgS1K4VHva1ZTDYE9S0+ZiThHbgL1
7Whcp3h7OFGtwUb7TBR7sDu4qgfu4rLDTmgo9hwRg0TXVhOvBqKb/YRvikBVKkvxlktOZGYvMV8s
EMvNLM4gsYVHvjtnUOTDKzddo87FkO9byhc2vh8yVY4w4yx1BTxlmdU/paQ+tCLkKfLwrN3wTKF7
jYSSm73Um/+ohKO2tk/CBHqE1H6WGUUOylwFQdI6JFz3n84eAVIWbPLt3hDAHJSASJ4soUMc0fhf
WP0xmNtP+ld3twkmpyRECihJBo6xnWkJUkGCahPd2Rab2oOh9m3h8k9MwT/JxDdk1lysyV1z41zB
bXj2C+MFhWE/1d5APwbufHZO/0+G0iTggDFYhRIKaskcaWOExhSNcyE6flGQWwiVQczcPaSKVMcg
rUc1Ef5u6NRsikCDYruwxSyR0S+QGwuff9JdFZk458MwNKCufp7CnHJDcu8S12+qnaahAlHDJQvs
j91d3zORSmoKyLDCKYeBRJvAqa+BWgl8HsRO2utxGEFeiDYOScAArGos9DwZmgbHJkC8IAvjYdyT
+u0/4ZaWVZDZur9NNrXOEjI0W3ENMQ3F2hRWztjNrXZVe3Tqhy+wCPATvOTlYbiJGrQtBgPDHYNX
qy3gGbiXYY5+9u66T/kAXDPNTQACj4XFpMWjR8DQ7uGcSWlLvnCd+bHvR10SS5tE/yfj2Xg3kSp3
BP0ZongNBRHPkGOPnF3jWjSPlpeiK6jWxmN2PG5jg+s3LgftOhzAmizJPX0eo7PyR+RuCN+gUJjN
s0RPgXDQOLtXqy68D8sHiU5FrmhUA63/rzWiySVdBHtngs/FnL1fk2B7QASXquVmPuc0OzRywRDl
L5hOAKso5nwbSxQB81b+m9Y3ebpJcRy/xM4BhHDV7jpi8NKiKWcjt8BEZvtwER62dqPlN3iKTeJ7
wHNjd7Ghm0+O3hpkELgNu+jclIRrBCYiMRJZ+m57xz+hOLhdb1ksl1e5vb5fxQ5g6OJbCNQK4Np6
rkheHrOZ3wlVYWz1H7PPSEZHd7dPHTNcuUPcjNItiJ5HMHovXLHJJ+SVdw4O1IBUs8yvYdnCsUyK
fnTqW33wF+euZp2yQ8miLxCcQ6rcP7PJqSt/2t4TyLLzxrzft/lnCmMvRZiGh/L0O1RXpa1SsiAs
5NBmrlshC2piZ3R9fTnLu/83ZbP6XWQ/yeCHiQucL1dXUP42G1dW5i2yYRMeFfVO7GtazmO+BdGN
PbHxMhztAGWE/3PK6aE9AC+ibWL5kWf9wC6/AqaGV7FUAsPlYXq72bqi9P6la7EPiTQ8dAEYnDjI
mjE0yyYysAfO0yRVb7NBmk0QUeuwaEgKRNlQGNH69T0FSwtFONCt7Q3T3+AYqEcMAgyW5YPAnsFC
v0GT6pcBmRQdQm4S22NmMdsIP7tU72yrubvLDYV2buJQlH0mU4sCphuAZHjhkSzbjULTMXzE5fDh
VqKQLklzp5HRMzbE0ENYP3yTFYejovYlB4x2wtMGg6wYVK4WiJDD6Ic9AVuyYEwavLdiCDurw55i
0CESt5EfBhqCQopMmGSMuBv69YvG6sov7zyhwUUCkgO3Wiui9AmwmCR3eY8QNhf2Ux0PsV15srDP
OpAFnQhSELUzWD74l2ayaXlnN0RBpv0BL+EPmIIF78UoX/3jYabiV2Zs/8pKCLuRbhBXj/PqMH80
H2qHsczxTnOKhAo95GMjWx5+R/th0e10CAhUTUjbxmqTPQl7sBgAJQuoS5PK1bG2AJJ2VhwASzcn
6OVUL6KWsfrse7XWmf47EhWXVg3HVma0houtXBpf2zNk8ms2flke8YvoWRY8WuvVL0hxvzy1U7Ku
LlDDY/Rafedpj7dKPPtgXYsbUvF1RN+MdQBSB0/01Sjkjlpw0FdjmeBAfsmU9/kDZf6t+epVUIfk
b7HfgAyeqOMz5fW3OoTKYtf7yrF94uy130/UAEwvDWWmmbNLNba3zhKPx/7LZMxCaH7numdOIUTj
ob+obzVissZ+Mk6MXgQBRTwqv74svAxbYT1EgOW8NedXYk7K8/qLub+WmFTosj8TtPYzxwGPcc6c
z+jLQSp6LIaZ8rzSNsxVt5a3H9z8iLXWfgV4b7uRGKZ/s1PsoowLmFur7/jXABnfXMjxGL6pSb+f
OLIw92Lblh0oypGJgNoxKrJ8fr93Nhs6E8Wbs7Dgx5QdGh3ian0EBmvAsH1qmtTfOC2lMNADZS9x
AjVp6YHCFzzYE5jUmdOGPJEPXTUNrWmHNgm5cFqPQcf9NB6iIHlEoqEQmEOimHspuNk0szg8xZhS
g7qzzHwFSuauI6TZFuSbOv3QAL+KV5k2v2JyLOPblaxxgVGZIgUtSCjDvlJvzLn0LrXLVAYaz9Ar
qiLku6hhZfcEwLiVDTcPSkO/YlbGb63+jy/eQxqf+deSEBNmvB1Q7p6FhnOOGVNjMtD3+5mEZ9Qe
+Z0uTX7eFm/WrF9lRaUgwXDjcIUZpk416aqdV2HJ+LPzQDrKcY84dTBFJBBK6n3gVLako6DigETS
Q2IrOF5cSK1SH77Rh1jVCxQHHZlJsixMyjO2W+FARVX1+SikzxTwLUfxk9ThahJZzQTzhq9HovoG
8d9gG5ze96EQrkiVzdVZ/m7jdwkN/H5QheGT+xQQ2YjaLmRo7IKE237rOk9LC7Hd6abkRuTe7Dt+
81U5F87qVR6TCpdZOTmAl/6k2iGpzqAJOFp1m6PiA4bTIXNBVl02ZThfWaYUl3AsnCGXuTBmx9wQ
BEX3ISxr5nVKG7IgvZHSINauQza5CAe42urURAXBOD2DIS3c3Ar1TMiOKHHk4h+8umri0FL4S1GE
sozH8sZLLLJT10iOSzH1zFrkZWfyrFZ7yWn1dAzu/TZ/rmhnQprbhQW9U8c1uQ7ZLZkr6WeQzDLW
Euk3mcI51d0nLhAEZ54bXooxGQgX7C3MEJpeGtPynffR68TF7WlGn/AzFuGVdiKlF3eR6eOYH8BV
iguSWP+vpPK7UjtrowskiJiR1XB9uYgi0bNQ9xj+pbPL54dgLQN/q0zCGzORJoTRgx6dkShP8Tir
p6065JODTZYaG9SdqhjtqDI4Rtq0g0UEbXQ7WNbiFx09/E2nA+sMLXqUJgigWqFX1ZO6msR9faih
lXkVRPQDgfiTvDcsTxHaYEvrszxPEYdjQkGruW8S2wIEkib6xNS+bOdfqHVFGuVWF7Ya75BcgblV
cHiYH24InoI+rVLOYYLPyzvEd6KUhXGd/0Md01dBidA7yai+zz4YoISSOWYEiAoz3UmJIpcfLlyb
K9BIApzJCzW/vzp2iUYfcloC4DrIw093lZEOO1jvqmyM7E4IAIWOxzy7Bs30XH20mRvgmKQ2+KD4
ZL9AdHMCZYJaJa5xbwAZaDRtYrzdZjcStiUlMTdMOLVTpgFrsgFQ3WnkoT33AextdXrEOu8ZxdG7
NqmttWL0eUVd3zvAnXX8Y8W7fZWXkef61Nb0gTfwVR4/p+Zkw+QY1MyGFXjq6KliWrrgTNNym2IQ
DfqYYmzImfX/oMeaCt0L2d5yGDZXOJwlaRVcwo9N6U7jlzWXpbP5+26RdPDQship+HVkxPHluriW
hnCOFk+9bCQVPgjxOaV3jEzRs8wpatiJaN3FuIIsyD3xnloI3GKWMcfZpj8CG3CTIJAaCfh2qdob
S7ypwhPIN5+pg7bOzbIgXmW5d9qf9aqv8lgSSW0HCtyIbDY98nnbc/1sSv3jijaEn8asadJp3CuK
1J6DGeaAAONiu/1z16PA4Q6g655qkt4xsT66MTAe/RTdqOLUp/7WHGoshbcQk9du5XWKAJ2jZ8uU
C+9DGX/KjKhbP5uXIIk8vnHdlYbv2bpcwtbJ9qVXUnXu0JogG3pfQnVUilv0fhbW56Bg7Zoie9Yn
ntvt8rlKyGeHkffT2lief4ZeTzjlvsHqZuq/j0e389+HDa1fTqsb4e1ClwIUOZMf5QqRjn/Y42oX
CskIYnS1IthlTr6l8tSLtns2Rs71u2dvZNwqEx5N8pPCcEIeKTSC63DMriTNTV8A0uhNhSXBbOTe
NBSnpJI/wWIiSXCt+4SRAaWMO3Ip+6Ej0Tz4Q1Pj5DQIDQuT8avIGmUJPJZqGQGtXDJ/GLWZyISG
J5BwrQScl488ZLTclf7WNC5TLaUt6h+CItFhd20qFPjbl/AjtQFa6oo1YiNE+xJ4U/ozptpwbMJY
9ATmOMMpEJ98NlUfbCITrL0fDs2FKNEVKzQ1yxz2yN+9cI644mFBm5jbutNoJP4qQQBs4OERl9te
WPRxHg5mbh9NkhvoWVW5yvtopD66J819Da/sg/Ev03JibMVyKxc1hP1NChMKZOAk6M+XQDUqZ1Bz
0XPOZoWp/9iMfoabjDGiRmx6f6Zw5WI9fsZP72WT7qGQ5Z5t/aoEOJ9qGJ2Hxh0WqJhYWR2m9iFa
RWDdikwl8V/9Eo7EX62xswfdsJfSrNEo8XT9njLNt7MqlJa/onmYiVSyuVr5JhB+uOnw3Zz7pIxT
yHUZevyV3LKzKjkV43fqDzqfU1PmBQ1NVQYLDBE1n/E+43pFOBx4HiXXH4bunxlEB0LuD7/3s5G3
DkimHzSm0nzjbtpmQg+T5aV8DPUKwYftE8R2IqkOtx9s/XE4UG4i1AJM48nzOOVVG/Axs9mvEcwY
F+wiprTgdpC639Se+1gG0WPmtUrSGE/3zdAMeyOW6JV9vwKssSn0ElW7Y1vdGuY2thEOWvsX8mry
V06oRfq/UU27estqp0Ln8OKj+NwtZCyUKvHqUrh0X7e/kUzBQqGmWr+vAXHJuo5CFYAHBvk4EFbz
etVHFEcdO96/0F1c65jR1/3cqjFtGcprfqjpCnryS7uoKcUiKB5eCQHbZgkqGtmmrmMpvzNT+4UT
sOinXxOvmOdG6M1wnlzYfy28PiA4VkTTpV3tm1LTdZJL8I4EEgAJhu8BRfPVzXVxDncL5AX0j2FM
MZ7/9HM8+75vFulREZgF4vNcNRdCNzYoY9m5wlp6m7AvZt7HIv0tbcfg9Up0pMkrc09dW9gE+D6a
X26DTkpWRqXmZVOBVMuoU58KI5GRDDPbqqy5NP2nvzOkfXkwNCnnzSOsK1fd70lyS5JP3gmeJv8+
EmYpZ2dOWQ+f2fA2a4iFfirZo+RIpnW5NHUg6zGaT80CC//cAXtSDao7IjsEE3S5d2WZE2n8qurv
tOk3bB+oW6bQW+454bsTa+GkmUpRSIamelgTgvsej5/HdQHR4eHjY38aU0lju5QD7eBytL2bpZoc
9lz0ZbD9XPfMcojBvnMR1dAXJP9vymcRDzUG+g9UK48e/FT6Wy16XdcRA0FMG2iej7GPVtqh21/V
DGj1CK/knSEyqca+twTYmTO+B6etiYvPWUvkXzFhUsmWaKeGjc6ir2KyQN2o5ZsRVWurZNO2fZMY
uqFGU17lsshE3Pz5cBo5onjevMlthsOLnFDyw+FigxPSTDxBM3wGrFj+BgV1IIOgfDBu+xeEPNcY
ukCjJOry/MNqOZLLOWJqhwF7G8kzo+0tJb5VCy7pu5I9fuc0ZDEYM2gS7NLdgluSvQoIey0CmXkm
U0XatFeBL2AvTKxxcG+WrAuWKF8TpuB82Yk1CSowYCz0zhFPMhJ5VXT+y7HHPbYsy1TI1VPsoWOu
fHEC8cIh2KaSiqR0paD6bo4MoveznAz0eNmgCHF91wSn4HnMaHIOze/a7AWdSgKZ8MHtZEnxxpbv
3cFGp+8LIukxYsFx8bOxethicb3sLCmMToAiM8nmtqcYeyVvk4zmGGYnKsFSqrK8j+AJelIrWrsq
5nXbw3FDBdP9bkzdpIzKQODlag+kA3FN+63hwpAzYPj2U/nwOKr+ff3Ta4c0wYK6+nlgyrgPVOgl
F/rvK8TJvLrrdhhqb6IOxh05cp17cqnLP8HcrbUXFhi8PkFy7LF8WkItnlZnvDuUuudOjjiTuNTP
i6TAp/xLVjyzVT31Se5b2xetVzUt/SNdmlHI4scc7S/tX4EmbG6IQQlDmFd70WGcSRYhe12loHxK
RT45Up8NpfOMqv60QQsF9g6sRuxJkLNHaxHk4Y1QpSxw5lGYzNZpPrL1sLYI6YzlBVur0DY8RTYV
KQEv/84XHk8lghqzRrUS22yDdKVQAiKkVNoPuylcia+sxFEny7uU4vCIXNlIYyiSmiouvvCrLWfg
oyZBhnKJWLQh4K8JkVwrwWXPW/xE/DzfGA6BR05xnQ+VEm+a969T0XiRDbzhNjwWsZdt6toURiYX
M6VNvuVgj8fJdwSlmOrtPK+OiB10/Z04P71Aez8dqQCTgBYhTy8Wiu7vn1fLEkhF4/ahckK/cU2t
3eXzdim4VwRBsTeWzLcGsIHPVA5jBDqBjzQqJ92tuXOI+E+LTWB4Ruz1vel5ncqlBm6xf6AztlBX
NN8vhjN8DlquP4UxAGL2vHcbLq763ItoCIvwP1wkXc4VywGINM5CsiUgkYD5tnhyug5n
`pragma protect end_protected
