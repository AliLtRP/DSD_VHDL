// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aL7LRO+g0BayDZkK1q7/t6sTfQeYwdJczetrN/E8e0/Grhj/oTBxLv/ONnPKA4v0
jas/gDJL2kwUbSlYkMw3juUHUuV2/FsOusN1BOnk1ngeVH+0CoheL9Wz0qVCoaNe
oLcBlBZKRxPEE5Z2FvYEJNKvfz1xMr209RmVcz8Fi3k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3920)
pn419749af6DJUXBLBT7GRBh4gD3u/ggdpECJU6lMtSwRRFUh3HgiA9jXTjGWgWq
O7Skk7lCVf2xSV99ehvfFZQUDHzvb064CqdSn2m5GRswjzl4Az0xrBDekjDoeePg
33rN9JBEqM0ANm8PQzL0fwac6E2r2NhLVr5u7dgQCwKTw22MyEZhusgFrMIeIUtR
bY8TOAwZRp0zVvTnu7woj5tyQ/j95NhnEltfLLZyPt5zUNtJ5gBGVyiTsPouHYTD
V9FKKpp/2HrYgSYHhXWOXi9VEgfUa7DjRCxkpKYR94xFpXWoZcW99vcLEilXbb3v
K2hxlY+dHO84WSQYd+31UigiuaVz5eEyI1bt/PnhMOMHiFLv5G5O1hscecPy3hx6
9Te7nf/LnVJ5INK9rtCQPhWkpmGYcFQbVvCXnlRRHG9sFcdzzqSxGtsLqnsS82+k
kEJoU/DuxzNJujT5H7hnN1gZWH7T7dqHENaqwMhygmrkkKwmFxB6cjx09Q9Mz3X0
gW3jydUhXX+B0siR3zO9KeTuTzDf4UrOHRTC+x4ewRsa6Zp69V+RJlwwCmCRpoeQ
oriqyUjnBwdp2XUDn4EJvN05uvQgBmv8xv6OqlG1/YLMoYmQutkmuwbET2963o1c
B0hh/6vnVoHtE92n52WCcY+CueXkgd9SHZDVvSZF1ayI7uT8lzuF70lDDuRVUf9J
eTteH3G4YbsGK7vro1UF4VhpCX8HKeH4N9YczpV6BM/Q6967tQ3fF6LAE+gR+/r4
bZ91vAh+x+jJOvSnOlrnNVBxmTmb97E95kCjsys+2+1jlcQ83A9UmglDE9H0ZBq6
kwrJEqoA6vwVk/s2X6sYyOdEcQYALNTTbyezqLlGudPOLGMixrgQJbBe+aIpmdRW
QPICgcQMHDCvLIKVJ6Vimcup9cLarqUym8AafUTAYxt0DwNyQCHEpkTVcyNr4cLy
WNyE86sZdS4mBqNtuGDslYk5oInQFP2qKFDhQdkdhnZ0ZK+eH5+tXhlQxR0isnFu
S5JiBfdQIcF/a5rU5XXPVGArvrCklyrI5WdFXCJsUUEeXkc43ED3/dAO1VZnYRR0
RjbWpay2CtbeAirsCSd2cZK2O26nkjGIDzrOi5hIjn9Fa29pAkjy53tuHFUV6dKH
/6z77ElZFy5QJ4GeqeNWSVCEwt/3AufzT/rJUEeseSGTwGIh+GK7WpPTzKdhBDS4
CaSAruAt3q7QVFoj8oThNGvp8D4asKSRusdBoEa10aKxkEE4YfC3mpa/l+rcMfRJ
ITcHjzfNm+4Xe+lVgRmOJgRpfRDECC8DcKp6zsNpHiz7rdFbGXDvuvs9sKPX1lN1
bGCq7dNXx3SHCxy4nQTayrXRqXVOqjnuJ/bCtIGdQJR6MNwiGMKbdF9o1XMdksak
mchJLeyUxrIgN0hEZrhUJEWg7IsrLDwwrZ+gkWIIOkyY5pJddspPcdDP+rZK9aUz
MnKN6jNTtWzlUBWUQEh0tGChKpY5JTE925ZbdsDNGLnUBgs40BVO8VRyMxiOebkP
v/4p2vT7k3eN4oLbj1KoHovLiZ7jLmJ6LOWiZrHx3a7SLGrjNXBANSIYwgS6UvJ7
O3dngRs3QrZdiDd435l1W0jR9hkvLZHnL6JsA1Nm4JlG7Klt7tTOzT9fnIYCj+xm
rS2i5MaKvq4MsH8w0viRydAPQgLMjUAE7jXbIjMJ9pQrSWmH2IvcKL1Gx36YvOg0
o+TSi6x0tJPa2G3g0VkjQ4CelgO/CWdOFQhbc6HR0SJqpkKjvN7WCv+oNM+OuRh6
/oEGrJkCeMe899/OWktsVI3FJCiTc5b+Dmn6m89eEtjaAYEHbEuqKp4z2egbN5hz
MqjB7E2uHGF38aLTLc3KLLAacXWRcDFHfB1OdUOzWTj+Z0qIm2jg4o8QHj111BHl
LCZp68NKFb+Nt/L2LqnwSL7/UvX7kH9satEPWM8IaJdzP9blxYU1a4wn2vI0gHcI
9PkQsGujreHWwbqLp5jH94R47QI57BiL5+7zExaf4m+S8hfegHKYAwaGMnF0afuF
cIamAV9zTF9NRW1/fwOTuXGWdKWR46Q1ipl4bmKRriu7e3Tb9eOpqlp3ZwbCM8c9
Tsa0zPxbHeiu95wgO4rWYdE+eZvUb9bNtgCmoB6WpFJ58OBYgMyrNcacFHOM+0bb
z4K1xdoGCoKTUhn8wlQ/U42YwtZNBf29iCMLyngMW6KjliDcAeRLb95jDsjfiL8h
k+UDKLTAKPN9zP64fPwYvBBzYf0bgIEEjfuOAqDQaGzRuPjWZI4s1EzUiGYuny0W
ZDUHSZSG89oTj3eIU91xR1h+KlQC3WBHETm8rM5Sx5FB6aMjry8bBmqoTI0C6Kf2
5dBxPETGI5nFWcwfvahhBEfSdVt3H38qFBCA4RtCBioG4NwemBClwLUD2x1PP6EY
nwJrn18NdluO7CbY/bC5cqr1FZnPUNgbQZ52GpjOMLk5/AQA2O1A9b35UnPngCEg
ue0eJjyjZ25frq1H4OXoR2XRpVFy0BFOk4lVTLmUYM3w2Wp7khSprvPyE0Ib0lAR
l6Zc/XTGgAZz6sL6Kr/y9YDTcfC6b24lSxH6C8Ei7Vsmjj7UPRjdcgir2VRBD1Ru
kmLlYmj+j1Atk8e9bqsDfJoTLaW5JgV+fM8xSlM4jX7MlOG68b4PRkyHW6kVmpkd
80v0eo8SLpz96Lp1N7ozJvSOm0z+Cgzf/GJV+mtuvlf0H4Z5xJaYGe14QWxfZP8Z
t8ZspbxIA9/LSRGUnQekCy+WPYAEPRaZ9SQweWNh1TqR5OOclGPitb2Vok2qAQEM
KHT9U2yd9AExquXJSHFhChyGkqMT8FXVBqSUpFPCmlWE8S8oJeC1s1PH30f81IIG
RMI+Rc/NYJ8jYiavNyNQDkNEyNZC/gAyvwxKOek0PFDUj1Hs9cZe5Y3P3F9hiMBA
NW2Hu+NI/8JlEdBjskm4ukEQIyHhuaRJgwwm+WGDW8iZPuT6GLnoGROb4j4aT97O
yg150lOpvRmU8GeN9pnLfB/Rrhe9gdYivFsBOv/uUqNlG0ieOe+B2O6JY9CZmNuY
xXLnMtYe7KOp/7KdR8cr79YC7wW3GrOHCP4DNfoyczryzF+wmxg0zWWvx/aQjg6I
LHoOksKpCbJspN8O25J1GQonIWSwexVXXrc1/stLh6+FXo3V7+W84UJ5XIq6e4RK
Dx7iOpR1HzpCT/pTmj9Vs7QpCAENpZmZLMuUmvEmAfTAEZu8rEHBdOgBmiFmE3M0
T7WZZj513Yby81fjDnY7y3aw8VfcvwN+9RJJz40kBJvyK+SIUy6x5+qopfYb7div
A5ja+jO8ZXpEua6JO4BXuFZN5CrsP05los8NoMli2cCr95Aun7i8eomsKgQdsVFn
zycJOKdtB9Q7vuH7WHudvNPn5xN07W/HEsR7OxiAO3lYVl0ntZOy9i/vmlkrCaW3
RkKlhok7hQSKSCY4tWAXc2JA+FzEoX8iRbDDibP8hihS092aArIM1XDg8tTjsC/6
rQKxkOvF9VuKYCa85c6Uf2rZppC5cc+o1fV1NHf0bM48Hi6N1xWgqSU5e7T/MxNs
fECURGPb4Tpyd/09BGNJwV4oz10CzkilCFw4vAeNHfgFSX4LGR7TWZz1qJ4quGoS
fu/KBn1w5xISEZuOoUOfQnOw38P2ZKkpN/7JB0FyXxqncUbeyRDL1Ie+l8VQDCj5
xTy1gaOjejCrYcSzQMhYZU2xKEvl4MHR+wOE5AgCBkbckkc5bh6/BhYgCjD+gcjo
ePGARUm+KjTpLa3wtrhZNdOUu3wnTz60hPUVlUVeaKwQlNjhLXce3TIr20HwZITa
VC1ZZ0aWse/Ajbpt1ZvtJDTZyKoSXDdMsBFgCfTSTNn/53VfRik8s6kJhAgFDX/j
vIdC69+jTXE48LHxOFZFUyFDUk72C0LKdzcnHALWb5jfEb1jbGulCjEXJOIKQdRe
8M4HuQ2jgbtoMOrEr8kTb2CzptNLU6fwydGtT4oBuU0HaUuuj102x5OwlZCPDCfV
YX/dYtK9QHubyT5L+n0s5P0QotM05zwhRC7Wf4TKE/B0dwnEL1VpTcWSud1AJ7Gq
Y5xEM+EfYELTQNzSLYle/6HsauiFox9CTam1hoMEWnnuQjTVMPlXYEw7zeETG8cA
M/xkXjecCqfBoMIvhXqxyIG9fMVa7ZyxMhc2yfpeNwRWKRxr8NZa8/pKLQZmDmcl
X+oz9dw+Fk2UOnPb1wbjgBQPhpae1Xx/2o0uUYzHsL78HROuPFciwdIPoj5xL/3Y
QUPl/xDxAvq3CB0mbWulOhdD+wN8E4pAx/GDZgqpm7v16/CVtwCDHdbEQtXvahC1
WG8lYxH4VI38aPaiWzvSPT7vZFau7r0yein+4dS0nlxq0F1XrXBc17z9bnt5s8ur
umQr98K8DE8P+tGJih59tFPWAEZ2iIYIy6u+aYEQyR1EyiEmaOOkVdvYibHtjOoU
kPBYxbWvbXa1x2iUH3VUai2pMUXvpD2LSjnl+AodxEOmCwuu5OF6RNmCCZ4ZlfLY
em8ADk+A+FJ60pbZto2PxcfO1QBcluPeCE2BwYwdX4FBoBfPX6GcBj76hVPweeSV
ONfdt0MqQuIvyIZZYwzum5hJjw9uK1YbeK15kbtgnN1kdHPt5nPcfR5s0WZy/EnJ
o2Ritt75mmxFD2OBimlNuLVe1+beWeq/SEExZUhcq4s4SN6aJYYzONVca0Ev4W5o
IhuAOseGXRusbWupvM6UiqGRGavF2YWxIkozJJSBPJvl/FUYfA/b9nhQNqo92djE
xh1GuuNBXOA/4wEedyNVLl6lm5zT5f0CYfJER3Pfq7UVZ/oe2wXgm2YCKSC+uQlC
US4sbtQ1x88rdBlTUrjPF6BQwaCXWxdYGCpVVRDUL7wOGVV4QIFO0f7FY0z4Njpt
AkCgGMP5ZoeME1qCP/fZVYYKrGsrx6Ks0UBZfbcXKUaQSlJIi0r0p40CRZtT5NLZ
RASRvq20yqYz0bSKAm2QHp7P3k1VZWMjJRsoCl4QBTgcMyKv1H0zZ652Zu7uqU1B
/Rd9y0Hg0HBhrHyzxDSP9OokxPTAJbtzaac6F3VmdC2/alo/OtZccAr3nv5PF4TS
5xgY0WTqSHmWYREqVar+2umefJ5IiBwsGGKIzKcH2tMbKsq+psoi5pmrMuW4k859
CjrqectppRgAtjvRK5wE/5vsMK4Udp8XRmeHHz1pTL4=
`pragma protect end_protected
