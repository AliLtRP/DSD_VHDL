// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
nLcgAeYIgfPdtTJsrxHxtWyp5oAsyJIXNvbc8Mcgf7CCI6ti+EFWPet4oBHuasVha9xlUHEvJYly
0UVULEHg/mC+KL/EeiPDoBxDOnjxjLdtAjYYvxNZkIIaAWTNoL7SDgAZQ8VWtNLGNPHDq7VdMg07
IYT7KI4OGT4/EUkLw/FJRjFkPk7wUQswTnqeuZV42R/UVD3PxnqbpIVoJ6IzROL3LD5PUnfwNXQt
MF6wXMrzrolQEx6QFq65Dt2NhK7UIZ7pFwI6iX3MA5gDmrj3JMRDnBvEA/GMDDJUJ0VY+votXt72
Qhn59RzdkML1JOZmVcNvwrbS6mKkoNzqm7H3TA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
DMa0ARXai4zEEIYpvl/aKG7GNWWYPrMTXJPOLuYlur6XXyaPWabET6VfnGMJwmGuvABqjqlXO3yv
UDz0u2uZuYrcFCzD2yx94jDM4DlCw8eqZh8ZmaqqNOE8FxVNTNJppxjZzZd1B9g4UJIBuG5HAZCs
0n/GJm/fevWggMNoRV0b/tUSDK3OFIZQ7lbcD22D9tZqPCrFFo5/rIYc48bdWQtNryukeYCxP5E2
pMqlKGF9IMvZ7mVfLNIp9pvKbSLMnLFejwS/KHsT7/m5hFssWQXDQKhBhqpaUGyQ2KzgSPZz9Xbd
GdEMHPHfqAKHBnchAHkw7RLCfi2fDtWvrl25vVug7p6dz+AARGshNouEwSE7NHbg5TpVsn8Tk0+j
YjDEMt9FGPORE/MH67K5wOhl5qLxel12Ag3P5yCVFi3falavljpPwR960SHuM9JoNkLKh067kat4
PBEN6GvLJORyT+Fg7zym2sGkJxby2rKDHUgcjFUoADk0NdFU+ufX2dVz2hY3J8765K8DZnrUPOz3
y7X9d36sc3XyvQhrfiXiL6xri74DIPNfen+mCXPitwbmyBJuicT3/uzKP7mvHgJWsFgvubslKHdK
ejEgQJe+e+4lKTadC786hgFUokirzWE+K4ogoRSdqp2vzMPJFFyq85WUHfxxLOUHFT69Sdy2OtMc
qNrV+lNSnof2vacgTN7TiL8f+82KrRxzcs00JiCoyzoHaid44UO2yfnsmkFqEjCN7laujwpDESYO
jzk3IWOPdC7bsKl/1xuxrJ6mTOTQjE84G3Hax4lz5WhzUMw7feCx4yjl0EAgriQcWszBF7RjgVLG
8YJ9O6K/lfG1AyBf+2MJyoYQswj2WOKySzKoCYh7ZY9hOWZjXaLUjvAlcB9df2IAIIzibemfwHeH
d9Pga8R7qfX8DRYMnlK3EUyDwalq0crHGoWnfS0g5NDnnOjxyJGJq15Q2B+A2Cw/FK7/DTEJ/F9H
5eeIY4UFl3ov7msMnnQEwnDVXGY5BUbkR/sNG1GXCbBn9Qnf4erj7Bee5nzjmSf5qZOCDDBsA9it
woAnAWbox2Mhx2YVB+3YntZQ1IOSEL6DX6Egj+JiZkZlSPTlwPHeJ6mEGE+EGe06k3on9PmRVmCx
nnokpt5uMoqrgJnMUH8Ohhz1sEaWW8k2h/NUri2anEdyYc2v2dh2XZkFyUZ8PruUlKt77FroLsrS
/e0Bxppl6UBFtlt5bUpjmW7oHrWGVJt7WZz9DdUOi4KrGl9ohC+ItqOZTzt/1nQqPpbDJNyOgATC
in0xitDliZ3eEw4CmEzegU4720bYRkk2ps8zztaqDVaGngYo3m3jp780SUMb8wo/kphdGGuL6D4z
b2MEpNOEuc8rj7u/ZCJFpq/2XlWIgU/LCOchSA4nrSFhr4/MQQTFqpJavVm4FyK7xnBaDe9owRmu
ua3L5aFzACJvgnM31j4MVDLV4aWDsxomcsiIK51dac8FetbP/p0FMXrXneH+1N3QXIXSHLfUPuYo
WKGSdO9Cx9gDPRxuagx/bcmk7ntjCa0o41ttajCeHpGixeb8Hc7m9z1hrmsG/l4p2G/n0Hbk6M3X
uORh3IAxQTM3eGSAErBvefI8/+jRqXEAE267fNUm4NERbGpsdTXvCpF2UuAcPjfP/0Tu1S1w3MHb
zlgjSKstRz2lutwRrT0wonQbWV3T3BMViEpwsaANQ7iww9fsqFMNrnN7EeKUJI6wXsD+Hf/U7Awp
PRh8KUwYPzHBOpw4j/fDpn8FXbt/oVivIXcCbGG2N399+mcJNRDZHp/3r2+5v9d+4sFz88xJ/ZD2
DQvbve6BW406XAwOm7h6yWPz8+h5O4JCjyvO5q3r4RPpJwsBpWCMe1i1KR719pJo9U1nnQwBGaWY
fCbncw9CPhdMl9cIR5QMZQvDV6tQO6uS2bjOMaCtna1xxUurHzhFhE5QKeTqQ9jkPiMNB1ExHjKs
a4KM/fUML5nClHx9q9PQMVLdHTDgddG/PvEuvAi1ReedPnZEIcFLbLzwzFkyvFCsQAHIjUyvgR98
GDFvgOQyOA8cEhz7No6JiPnpHZNL5yzlYLFHSZ/O0lbpjrr1nANgF/RSDE1stbQSEbPvbv2fskIP
YBmAF20cWyrDmbiBWYOwOee0am7z26xqrpUbL+SmplhUre7SrzSUzRoJOO0p204MlCMXnCiLJDJw
ziY2JMyUkJy3tQvDeC7BWOKIFcKu/oe5dtmvPLNy6nZ8OcWiuSl7rPCN6jtwxc0hAl00+2eWEKkT
umxSsJWulVQ/RG36dCDj9XQ7D7UZPJGuyNCXKP75jwZ/aIJeitnhf0++gdhFFeJWW3KhH/4IaPlz
Ab3A6FBFG+OrxabJoJUmKdYEIeDW6jyUrYnOD4AmXMAMyHbHHkDey8qUPpnN9bZ9aznYSR4qhD1h
l7O+dkDrrvOA1w4/IDAzSfOzFwwGgGtJj6RlmGnQ3fXAAW3YkrO4nLm8g1zgaimPAFpAIpRrZgly
Xdxz43F7jjloo+ZO0Z7MBp5SoonW3zPOB9PDC29b5A8plwWiT5U78lFfMHYGnpOPNq2XgRntV2XU
vxBBHCWIFsjpnP05UcUBRbcRNWAPZuRD9+twklZio0qguztFD7KebayIpfe1Jqgl9EuzZrg+axXP
HSiIvCReQ2DXqVAVLQUFmZgMr4/0uGv5lPzF+JiGURTfhPWROggiRY/2X7q8Uq56j6BPTVOFcMHP
Tl76DzjY5OoTRDMyKSU11EKm27DAY0cKnAdUQPziqNtZJ6mdE5rjWJrn+D44gIpjkdmD2ha2JnvR
gCNaWw4eo6oMwN2iV/vWmPTf+Q7TPr69ZPfinFWf3uxwp0qyfzawL82S3T4yFo6iJ3lA+bxqCJtF
WyEA2Dku4+Ok/s09E0LSkrM/lEFx9fhzNzxdikPo9Ju3qER5vV7R6IpJVujLpRU4BY6n+xsh7HIs
oEIlg9O+vKg/WBxMsWvxJ7vje2QdQ7bQZ/Pp15ZPYdoJRg+aYBsn+yGaLigD7UwBsjSQUd+IlfmN
7XDHkln/m7r+H7zvjhvRB9wOd9U1/J39nhpk/SLUe4Gu9lK2Fb80QZJmriO0gsq87enqEFwhVOeI
zbI7hgEKyM0+Qb7bZhWGyQc7LkwTytaUmrPw7638sfMoM/9uCVLrsBlBkTqeoEYR0139Yu56gIcx
boq6KCIjZ/PPnUWb1mI9fAcF6VfVg3nUQKnrmCt3MP+VQpBvIp8UJ8LEVLBOurW8LqsJBp8W3GaY
2q4O534d8MYcwuIMjeEhzLXR1Halnooyxo8fcoWE6SdocDrBKw9XefeYImUgZenyvIJlZVEKwl3t
uqM4abkPl2YGvn2vgfgOpXxv6iZvKBKO921yjmLrEehzF+jft0QN9GgOolpBilP/I2UmAtA91IhJ
vso6YZluV/yhZLBLAEMzuHkCP0Y1JOpY2nOEB7qDgiOjG0epLrO/ZXV7loWIynjy+HZqKqGofdqY
nfT3gmexM88AjpuWrPpg6JQxZwOLrO4lPqOnl0nPVlVUB1tHmJdExys11enVcwBdiY8UmHgL0EVa
IFsdufYATnsTaZJVvbBwsOi7gaPMT4QWnBu33Fva9bQwpBrXcxkbKS3EZGa0djqC+KNvu0CAGNE3
EuxJJaJnABa3slkro/DfgCyboCxKXzUKq48L/in1gG0qPOvmSeCU/eH8IVC5YP0KD7W7sj6R7IEQ
OoxR9ezcE1+E/+4hSfSd6VpcBKbE+9SFhn6ZLljRSDETUX4mbSxgs483DX/r9OfXYGhI8l5/oj2F
iszNmjPnu2VKaau1CtrhhtXO9hGn4WO4qg9B4t7BzKrDcjIRxIQ7q1wJ9JIvq+2c+6zFAmErhgRZ
kfpeASK4sOtkmRGWa144twID59BHiUr7aURAXtSJt5rA1nKd2XPRyipxyTa98XDwmaUU3saV5Kwe
OJbKAZUWUvsqt0pMslUx9C5bRo8GQDK5Xia3tvlX5beK7lMYbJ52zW1kbgMpMbegrrp+rY7kv7rh
g0FT5LgHEgENtter18TmPS1eP8w8U/HAOqGmNHG3oPrY85aJ0DGglThUSYqtnpftTYXw4N8tCsL1
lgOZZbp4RtUDWLYuG3+mQJ7VkMjFQU1AUtlY1lnZdtO6vdeoZtf4m4GKV+b7lomN6rUSzuUDOw7X
q67QoCkWODhZUDLt24SwKfHQ7RnO7lI3L2l3r8nB0eDxcIM5BYFJ1AhpD2RQl7cIpE9Uxjm7e5Qx
NH1ov6OVd0ezl9Huh9unOUjto3ezpQeoW60ZF7j9TMwZS5pmemt2z6XGQZNcRMF24F72rvHAL+M0
o6us3yfCSPjA7jNgTSrZKJGVI6t10fkJagnrdrKqQVEgcKOoTWCs+8+V2YWnmm8laGKIEd7pqciT
N30E7s0OhnFr1gpk+nmUwH/Gm1lQQ/9l0G8ibEgCGEeF8ATvfTGB9DIzh+YlsLkfBKvVgIVGeEH3
9DZ30u/euCFGUTBtQSVJladzsY6e5JHZMS8sIF0m7fKIWpPoQyrYbXXuSnHScmN6K3X4RzdnrDho
O/yRXj3NPR4e58es/JkjE19EQRE/KHTHxg4HR7GvkpNEBtJD42jZUh3kA8HBS1hfvbQAxUSCxwx3
tOgP/DZJFUjOpudGRVlRY3xGDvd5Y1ow0eFZeOhKB59WUr+NGLPcN7RWjTCm94KeM+Qlh2BjGBUb
qgoA1a8ZWnfSzDdzEnAY0rTAhUKAD4aBnXvhdoocLSCuAxg30uBK2M2Nzi8hCAqOdBvfViXz9YPm
7Wscbv8Fb+XfgB42nEg7G8It1CwUZ4IN/zsgIqtRPpSSyNCY4PSbv2huuN9n/GQ+JEUjeft0+pvJ
QSIbEFdjUaqwUBbZdg5BLHhWlTpgztNiwhIe0+peSehjhnm0Hb/Nkcp7g7TsfHRNjWcpTXizG1Rn
bPw8PBYzoM3RBQ3corI2d0w2yEGP673+VYhHJB/rtikBIxIts3vqSs0NRM+9Eq0IFnQnjxuaR8ts
rQtci/2dLPSp/QhvuyqpPwc819kv/STDRRxvY3bbDTHOyJt6urfBTVHSVpNyjDLV5IhGJjl8XAJu
sbEvZl+rOFJolyGhPJWf+WM0ik9k7+NY/pBJjZz/I64RfMX2O7GnRuUze7udWJ5/bSCkihH6RIA/
gK32+cJcK1ahmVHJbpxrvqbWbUZj42mpdDnxOOHincP1kWkhw8oN/uNS/ZsMpuyRBLZ7tnicR6ea
cDqZsY4n0TKwG0KStKLAVa6yGlb3I3uKcyRrYTbvmnr0RTa1LQGhSWUEMpRTKtoZ2Xk6EJit/aYD
YYljcPXROA/vS1Ii79R62H+bsnVPfYogBKschD9VXzeZmVQKLX5GA27SwrQVhzCG0aO0rvGHBde/
kqslGGjgWp1GvPwD3VExy+bZbnmg1hPiArcMXQjey9S0df96vepUMTiAYsKLu9aEbsXJ1TE7IVmp
CPnn8ioUOfu6iz0IiTWIWz95c0X70egiJpibC9ivdGCJ4DrRhqITFRc3VKU84ejJx0zxt7S+/AS6
DVoslEtaZBCFuIDbO2eCqzmSy228ae14MgDqrRxLjJabKSJ3A3hr+Q2yQ8qfqrGfL7/1BcO5PFGV
TBSaNduSOjgGPmNBS9PbPxrxBP8hxYMgA88qMJtSJOF1oJOBU3Lrb/fslNkhMJbISm0MWkNuK2Y/
zSd8LlFiCg75NsP5dEZuIYDFtjkhkere7ss1/gEnW+k3NFaKTh6q/CETsOlTzESwNVsypEh4kH33
8ikh+SeJg1uU2pXMznpxbBQuPsroR0I14ZyIh0XukRsMDY1nY2LcTzfDZq598bnWgd1zn3YhPNIe
Ah1VqAmlQmttGuMD3N7zjvRqXm/9xD3WJkK70woHdAvpSoZKEsiuHzPPMvmR6XnqAR/Vttn3rjFI
pqQWdZkbhe11ZE8wUTDJQsJRKU+ns99tCMoiqA2dDnbpmpW9MiRSd//vFau9p38pvQD+rmPvK4Cg
FXIxcfrvEcjJZc1azMusl0M67DjnOestYo7AGkeMxONWLop5+G0SWMrz9sgtw6ZlbsZwpLz5bWiq
S6e6xe2lyZv8g6DyAInWV2vG+Ajyx4BwLx9Nh7voGFNC7cncvqmaBy0mfroA01+dRd+7BQEKNCM+
NH2NFRhctHzeqsvj2kKHZXRgrvmE/0t7A0gWQ+PEr5yg5M50/aVX561E9zPrUKQACqsxKxTLJEP9
upzfCRqJurOti8JG7r5in7ezPl10dGVKvU0Uq2hrMkCTkJ9m9xw0Uugjt96Vpx3QBxVC5qr01Nd3
NEmlYPZoL7I+60c9MSP4kTQwJN9kj/vgPGbL43fGTvQhFFzxXNXiJxdYPwxIoUoJRPykWLXMkxtA
soBl1keWy2V5BdaR1D3MxpLD3B5mOOr8VdfBCAdgyqwgKTQLymxdNfRxBknCpZgOlaVY66/Y0rc2
EW6FAtOLocdY7X9xnDoKkQ4noglG+KHgSbOctrd3EEb7VOTm0LbXa85nQ6TlfAw7LtNW5/UDfB6g
OMd2U6f93ZqRAKvjJyyztPMJQAm27ZyEkQjx1kQkrnwQmK6AeDIyrj1+KuKIG0+LySSv1vS1MV4A
BrYoRKSgewuahwh5VTEldYorsSO8altksgSYSXBCqGGcH4/b5dbYBAqq8+sht1az3HAm5AIrUVPT
yFdigkAfnU3NuDucRsoerki9AzjOv6tQCxBzw2ghlMwjRuMwcFduHUxqWFwfP3XZTAWV1+p1ktuQ
kvI/KNddVCZ9kMirsispaim/sEa5vA9BHLl/09tZKJRilANXuSryUyn8ZYJPiG4dHH+GbvU30lt7
ajqbJ+4tvYtGsFaaIoI5oekvQoeYbrvdD4Z4V/Z2WZSzb8oHWfU3tecPMTL6dBwd6OQDTgL4f45e
aJzDwDgaPGElRqIcf38MzvLpOz2PIrn4488XoPyn4ROyIrp4RX0GZST4Pv8Zcm8XLnDYA78+bB4d
AxokjwRPuD7j2LUf7UR98JqTV5i+lL0mX4XWg8bMzYVd/UHcQY2mRsjR4ooxCQsSKwIi4+7qWxfZ
i7Gyd5TO/T3A6zDadMv4x8yT90Mz1MwyRektMD43pCpogAqz/N2zLWKgiAZv0UY9BCpEM6xkAbS4
Zx1C5GnjaE58g+UT4WcZSqPnlhPBdugdQevxE0kNCDYISxptgSaMKmagEvSI3mNdzayAjzhsCpL9
BsRymCUzw1eR9+VNhX0kwT0kxnK34d7DCFCBpMcfB+9dzCOo29bNGiyM97Eh6O+pKJYUYkMDr/FH
m2lAu5QNV2r8VfgHernS7ROVcWJ0w/C+BEnU+UHxAMsG7YQjZR/ZMZtHBlb/erW6Syqev2OLi26z
AL1wAM/jnMv0MqwEo7spcJtBfi5kTxUPouEwjaI3LKo+kYrb4+0eETIcCvwH6ZH12rhkJ0701vK3
auigpAjiaSIS5wW5PYVgRzYGPe2Ck+YQnvbzNifEosIKYVHZeWtGGwPPujQdxz/0kyqDPv6YwJFX
nbut1UBMEjGtX+/4KveE3crY2IRz0PkLjwu+rL/9Bk2QNOCe9Z/8CzCpV+7+RP9Qczsv1aP9n4CR
CkJNYa84aXTdwopP2rM65VqNXuDDeT7dflrfuAFhqfNN+3ZoUkExgoZtQNMLRlnERiM66qgsCuu3
j/CaPf7aCY/BMBMQ8OpBLnVsmr0o+16ZRjw/lGaI678nn5J2O8MYYoQ6iej28iaUrKJcSwesLKCW
+kOmdjtZZ4m5UQM1gO60165Jg+cKio1OFFBW68OCNT8sMHdoYFpbJPDNObI2SfAkhdA17zqcufki
LglMMVyg9IJ6/6iECL6Bvjpwm5IHiqMR9pkud0xT2e6NtpWG4DlaQXFsZ00piv6iMppkwsRdQ2yL
M0bqcsk+3A+ot9zaiq779EhKI/7dX1e/KFJSIQvzgVEi7T1+GDxbnRr1C5HxYYxb+N0F9EB+HtBd
9z7RTNPtMuX3M9aw5KZyJg/MKWUuIItbRF9SlWoWuVntlo3cOdykY5ZkRe+K27V9982ZmIIgLHz2
DKyah3pSU4BZX1gnxz9AIeS/87OoGSv0YfPRVyjf+p4XgL4WTr4fDfSkao16ouNQlQKPjWRYb1zo
2PvT/NE3U9CqXmVkvNHVkUJZDgzHLwjufattP92OQhToof1gxxk+1sH6Jg4yutjfZLIjAnW4GihE
yhCo1UTgJYQlf44Hr6Hr7KAAXHI556B7XxN8rjo5fEZpTMBEvy+OsgZQ+ng01a/ssTgzqyO1Dz4v
ojTAZyYuFZBSeMqUmU6EzigF9Y2Mu5+jHOGvwcYTqVffx9RkhSvC1Sj5R7bnqbs2mciXCA8SdzUk
4P8Uc04cTi6jpJr+d17ERqmHS20C2woYp8kaKc46DXwqxDAOHiY5Mwy1yOSNd94Ry76aI+6nQw5d
cksIK89rExjQwC5i2mj2WIJJKyuL7Jp6ca/fv1Ws1g9yZa5B4xaW80OF3RIwaKZXCJ3pvhNpWA56
0bdA+9TJnXOY/xuiTSCOEsDr0af1yqis0Se5781rFay/+Xj0JoWoBndZpA8XNykLW+74tY5rv+o9
4n6WFs1hwQ+ztpit6EoectTcVBunyGcY+BCEjvBJY9oDH0mA8gvk/E9uZpZkII+UFup44BWnDosK
rfGdtKo9Jb3WX8pIgERK/FqELepWT+Q54YNZPf0dKAFywWLCVB4QBxZWi0Ac5/GeXjZQ8w0UYdpr
yTqcgm6GATf7TFNUVmuYI/Mg2XM4o64/TV3+RDcAqwqw8QatysVWP+XoXry4Ugwo3J3H58G5awbS
jeQRYK3hO7aY0ypRfrMS3nNhm40RdmJRpf1MFHXxzF6HI4j3kzuutfCQwLCbKvdsP+ipyXfBDkae
1Y1BGxIwtn7wA/Fi9RnwsR6pVH91SJcgUqEpqWSCwNl6rucqrxlPwZTvoF3FvSMJaT1WJHPyyrv5
JFjkKEeaPPMAiSVm9xguM1Xd7mtvt3UTPIeqExkoQ9RwmJ4dw5m87EYdNA+F0jzxnLj2qJVsDaoO
pQhJUrUJJNSd8jy4gV9rGpWwnaXgtOvYJ51fnvcpC7GG0XXykjAIdLa6VHyn/7kgveAZD53PAsD9
WGYxDICTZcp0PtDh6mgW0VL38H7iGGA/TXMXG4HV5EsFbARu90v6yEI9VpD8PbfNjwvCS3oCftV7
v/ruJRSZ2oSgWNcMvkEHftO4xFzEy6lmnJ87Tk+fao76NwfpgrBacHyTj8YMkaH2YMXQPSoS42d5
c0uFs4uY8wlzKn4fEDxcH4bIpVmSmiGBzGgcrlzlYpB/deHrcS0eiDZlEq4lSwXYWUo7UO++vVH4
uExH9zdZ3js/a8j2MF4FAFE3OpIU6kX6wC95ARkLV0O8qfF4679MAUN42uLlUK2MKklC6jsALgNM
QUQsoFR/0bYw3ZQqhnIMrEt2S8YYKR4eKUiupTGeyIW1LxACRjVtz5loASvCdWORyD+L4dfsHANF
b1Dzf4+TrWVWXv0Cl4Ghn4KZtXwOg0W7SHvBfMoGJfl6vzSwJq5NBKW/63tVezFlWcUsmnwwceL9
4UG3IQUG3unOQ1QuM6ClPMSqpcYXKKjQFAnYHsxYgV1S1ZbXlgZlHEg2x4B/4kKchDeGsToivNRL
b7hMRgHi8lvZCYec+dsec5NSw6niNGWPz+ixr6Wzf5CTGtOpn7xb1yGv22R3xmgDxfnZo96KoYYB
oP+pLV3hdz/4oG52iuG4rioLx/RqIDH2xmh1AoLPOXNUKNcR7LS/PJTkxICeWVsPKzePkL1tAgfZ
tbvpvF+MOq1YE19qHCbTSeT/JK/J6VIAdMf1nacPIEKyJMjSfRKVW9E4+Dwg1nMXkQmbSqwZ1Dpg
NWPPXsM00s++OtXTeGNdh6v0pAZYprTK/ccqxZJ+kyrJqXP3HuC2EKn8IUBYRzr7JMpDvG9PlnrA
3Ag/Eeb+iYzCBHrp9rjj4n/pb3A7/gWiIVNUkQGvbLm8CdVjNjin+9D6u141hhm4d3AGDqu7z95V
IOyPadDXiI/c7NsGoaKPrM4PEO1BmVJKfbVfI5q0pu+xnDKNEvpPakpFvEIzVCWEDALnRePfbrD4
QQyrDFUtaucNWY+76QizdcBCPxxc06ieyFFqGW8nKOk2mNyXzWDqYvY1kcWMw6VXwm3qQ788nNSA
jj/E2Gq0dimAjRLMT6TlCS3dJDv8BQ9o5uF8T4hnYAo7vt4+wyJdFSpmtNGNY4uvtGnAQ0QUKxE5
548Cxe/IZ29a0hIkn2yWKGDUZtWtqW0LlcVYPRtWimFA3x3i5jUTJQcJIR7DbciK0AFcyjiVHNeT
MRpMs7xnR83ZEMBp9rjw7BO4lFDTlYfK+3GFcHEv6Dg1czJI90yEt9ux+KvmXzJNNs/VguHcYxET
UyhNNbNM5C8dqh+bKEuDwYv4lVCpryHbAiy6jpGSmj5Taoa9c1TPEE5Kq4R6VYBnCG6bUKkZ8K5P
au4EIJHavqcERlraD5P8Opiq0lNEw5MWmJ9fo5yebu1f3hccGaaBOydBUBU7VbOYpV7+IEvmTV2R
hRfaRejiw/EbnW2fVwjQOZhwQAPq/wNLhOaq+oyZXRQNZMjXRIA40n0/nqkQsj3R8fA8eEqd6lQ3
ccA2guzJ5C4eSEOUGHLHs+mskgFATvLxQbECqH15LmNLQLmAUHgPKvaMQCAPzV4IaUeTikVremaP
p0G1oX3D5b5vHyHv/TTZwCCL9VrCaAWZuilQzCxmFVxH9GVfRAF2ovP75qtPqmNmzxS8zJciJ60u
C5Dxni75Eyr2cCf+lgeqQIDdKy4wXklPn9CE6dt4hJn02Akk+TJ2zz2fkxQMysEL/K9/tagoNP4h
oq0yBHc0oZXCcLYqei6R/XajbdrsmYH/cw/yqeylfYD/p55lRhYduiOJNdfr/iCV5brz+EgIcIax
lygLuYO3wdLpSVUshRcyBXXakgaWqVeAXKyxIvDZf4nq3rVmbL6Iv8tegZcM2Lm3/yqPGaMys/1X
xJHjGeR+41T7mQR/T+CEr1ZIi4W1FHsFWpTcLgHnFMGk/mS/GGkqv/4SBR8YduqJi/I4HOM8VVw6
cyJvUslrQUGF6xHY8WzXRjcGmwVVtX3eBE00NbivNvNQc5braJdgOC6uboRErF3qbMeogZZmBTO4
tMso/lEOCjGCx2bqi7PAWcKu/kqMnnScgi6ezH7pxKnD2X83TjiI7gUbrmnSiZzBu5tYh9PnGLFo
MNjgLer8KsrV8fdD3cRVBmBOYn9HPLIDjegMejFUqnflmQnRVlS39YbCAMvAajHR9k/z6Kw0NGTj
yl6gbRmStIIoWNbNHCUiFpcYwxitYyDf+vCUV9utlbL09jqoCsYH+8QQyAt7/0Ore9ouUkCawI3w
KwJXxe+7EMGV7S0XyEm+qP4o8i7oAjxjKt5p886nsqy2oHSgdf/OFOGBT/yJNCT5d7xQ/pePIfDs
8FL5YJW3pp00rdwX7GT5mXcutJG2zzGf3Ge4ip/55uvu82PVDc8kPX5un4VVnNWxWj7qwXN0xqeZ
zVsAUxGo9IeiKed7gk23a9i97RWqIvmYRL1W8PYElD76EaLsSc6eH0Ut/chIReQDlP4PvupkaIp+
X2/UZdCuz53hWje0/tsxMoGUlfCyQZJ0a7N/XgfLXWt0NNZbDu7dhu5nKcbCB/nRwKSsDYZjYzuS
Is7bhUjB9LnO7/Rifmf9FfBuLs4+hTnuIjTFFz/tZc/hr/t17XiNgycmvo4UqdVs5UgkD//UJ/hY
33VSaRr0CyW7fvxU0zQlzwAfX2cvDq9D94aQOcJXVNiZVF810Ar0ZzuC72SCc+qhZ0Mx/DHnVCb5
n6FWkIhoCs1VkDI1nF+DImPIizUKdOf+a8Uwbq+TWCpgWDBUNo5MeEio1G5kUPcMrNSf8ypA4lLe
Kx+EexXXYJIYxQTV4ariP/IpURb7zJ5TKEVLBEHs+ZSxUWrKdz1X5nRfxIcRwAmHJ3fN8AC96/Ec
plc2ngvryVQ2Hk6RDYjf3jax/rex8gaBohHTfu1LtXzKfr6DntMOAnNIP/lT1SUctW1zzI3OXb7F
93IYNfEzeMDbP5fMgYIYeKUIjL9ZYQM6Nx/JJPzdhVMoWJg3s1xUUnG47iup7Rt/MzRi7Vz2jzMP
yFd4dEIEYBv8YED1O1eopnvCa+JGxdoyXZm7La3vemSILqRmYPGKO+WOBV4uTnnQbMyXkCl1NX1o
9AaT5r0lcZugjxT7SBiwNF7P5UnymrCje2k7R7Adc3FRyW+IHWn7cY0Rs739nvVsq2WIywB1K6s+
MKH/sThbZCnLc2lffK4k6JD+qWDAH5wL7TPpOhLOtPzrdSPjTnxxIqOHsy/AYyKj85y0hcwsBFVr
Tny6IuhnXAKcHIubFmjqnSWVgqH5pn356LLDLu7BjTIi8v2WwQykmcwCkeykR6K7FLFeVy0dLFpB
QwRKb7OT5Bm05FvrUqcQ9tPCJ9MS6zsUuOwxGuNF+2XBoIjh/8eNMYGPJxJZDCEAyBzrhCQEXuLS
djh0u9AeWNwMIHGktVzgDamt1zFn5QtHf4fQBpi2cp4MGlmmDhwJgRGnEgLTxabNo2SPdz++Ur6k
6BqwaQOqu2cmX//g9hbCns0Qx1aCrV0AGAZ5Q8uivNJ65zz0wRnNGAvW/zOSZqmu+KW9eQe4HhPI
dlzECLptnp1EOpFe95eUxOvXn6WcgfY4MLNVf64bAwsb6iZt3nVmU8tGqERxuZX1utCxgLl6am3m
dkKHlsQPDZgxFc7xsHeaoC0wYfGRXuLDNcH4Va8AWMYLAOUy/Cemkak5n3rM6iOG6deGxgb2SYBz
ywqQkEqwJXk3d7fcarazg2bE6kgGHIsoyImAgLTZs22vVswtUL1gS+zibbKFtgGqe3bRhDW9KSUg
5PcK7+gwYlSUFCwcS33ZfRqMChkVOqUU71tkw3514UewGvum4zM=
`pragma protect end_protected
