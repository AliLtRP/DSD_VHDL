// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jiUXhdsBNZqtcAdSqxa/GDjPvwzPTY6JJc0eaR6ZycxqR8uTtY/GMhwretOdnIKq
TU9oaJpHvYJ+6h3d9C9F6nGFKoAYaJjT9ZOV61TFgnMTm1oJctyTSsZYLRaU3leq
RV9g37yJOt8Q7s8JI6Qh4BFKw0jx1TDzBGP+bDVesY4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48896)
WfHDacvPdI0Gbtl4n/nvOUjRVJIQXPE5YY+UEhvK70g260h5uNsDv+uFtrJWedS/
pUlxb3/lymYH1LnPi7DAoHXsNRUclkeG/T7Q0luPfI6B9zADJKyjAu4yWuXO1Jt8
rLxoisnSkbScOqF9dc2eysVR1vyMFSt3UDUJvLEY9STbnxnGDjS3fqjT50Z9u9hS
K0k9nbSVvzrM1/fRjJ64DDGYAAYLeXSVMgrsktJBS2MDpQDmpUVxA5CWsKpWwzX0
JPGJT/1E2Ge2hWuYUJcJTCBk3kgc0wK1Ha1K6bRlLJjC4XhKNrIKPGENTam+p7uj
E2LxJu8m2EG+2ZzxlTTEEqsJauSaRXmwq5t6gdSYN9/zLyasuZgJvvrnldzb7Hl7
X6in/LcjACFTjYq7l22T/MyqtRGKOGvna8YfibuyxJr3kWfXAiN1F6gCDNJDFBGH
Mhs9A9D980b3VnTtputghyodtms8FbdGgl1dkuydgLm3twcYRPCgoFhY1qynJhg/
/nj4jfldtJf2C2vGz8r8b/KYMZvtxee1h8a42MjvkhWpWtCHwzsac2U9H7ipwcp1
KjG5ur96ui/LY7GEOKlseWD2nnG+XevkQ8stK5ATSZZjGZ0jHzqpFyKHU+rhM+DD
D7KzMzt9dDdfqHlOr81RzM9GUwdmPtqmE1P/aEEqsrVo+b80OcbfD+GmOHJC+W0i
Ypqyng9Bk3tucyJqO15dFL+LxIKIkVL/EIkc+bM3IxVSql/FaRqgi0bSuCS/wWkX
FWhCNb+6tgad3Sihz6SDChEvdMRbeUFQNYZzvqpWvuE/o8tDJbTslx1mi56Hr0H6
k5TtOZoi6O5S4hlc7bXfjtKkLC7037x000bZoB+7p6Xccm6c8jL2DJ6ZiqfKvNUF
JapDFtYk9prbpuEaQhmFsKf2tw5jV5OCoIuBWg3ApK05OoBDM9cx1/OBPPISVHD7
OkPS6gcQUrdlemes5hQbkMQHJPhQyqUsQs8878qu1sGlWW/pJmfHJX4WoDXKdN+b
Lb5F3/BYE0pTtKisnLyLnDQSLYJm8soPlEsd7qBBzslYhyz+uOy3axRyUIVOndML
jr0BzU3diyG1q/FlXF9he9Pb0eZ89UmdK2GtwXEYcovPBxlDfNIYd4FzSfvP0+DY
zARTse7NXLh6Hr0A1HENQHH+sgwAdupeME1f/KzAidbUoRJJYxCbdYJJex3whnYn
venAWSu4F4tWbUi4H7hQJjL/x5kiujBBXWhZ2t9m7p3+djxE14YKZZ8j4E94NhrG
T3rAJHZb5uLdg4CL2ejXzUAs8/sHOqrdeSMFigA+kI2wJmDXv+5mnh5aGcVoWORN
j/uBWzY1Y4HgSJWEq1Hh1uJXTC9rjfFGmmeHxvCoVP6f8X52RzuA0s8M3L1jBw5b
yDodXJBY2CCX2ycWbFJtSEdSDyn1kMgi2EcA4MZMbGb2ubvg7e6G77WZm7J3O59W
UaNuQcYmZZex5NG42U/wf9qHsIKBFBqPZVQRJEJ9LLgJME5zOZQR4QtVMMMkjG/D
cABYgGADTVsMd/WR9Wl0X/TfP+dOLxu5bPKrWmseHoAJ2T747KlWpvVethz+VmVV
GGOrtsSDOb5ll0T7LftMpeEwqTfkqG4pM340pi9ft8YvG/UKP3i+4VEbLaXKHsQf
IS5FEpeKgk7eR/hfDCZN2C8KkxHMUF9FMLr5Gnd7X5dO+sVAMt1P7qD/GnKr2agF
brbUcubZC3ZUwmTIsmJQoIxQnR6LvKDXwwecwjxycJVc4VGnwQYG8sSwOMN/7PAk
Swl81mxOF9tfCK7HS1da5fLD8brVulZyK4b4KhPkgqgpRmDIg/S6gmk9v0fc9ctU
D/jSUqea68ee9jaKJd76KQOnHUZ7KVOrRxMSgmzSq0fSZ2DwiFJuwImUuOuv4wEM
qss6IPleW27yalCXhvRaHVRDjNZ3vbNeQ3yao1STtEAS1p1e8v44aIzD4WOWFPpX
zi828u8FEFimm/BXRNpccNPFGGCbaLevOt8Dd62TgFxQbHiaVcej5iKy0TFYF9Rx
YRFsS3vbQ+gKizUoMFVQnT5z4AmKKmsjAjqXsL68REB5jIXYA+CfNQVpBu9BCzAp
m/ErqC0/Y7W8+/CedoYebuN9g1P8a2jvkjcodUS+Cqfmz2lqg2P8D0L2oqMfQdih
I4JXuMxIJ6HtYs0Z0dn0l5KmcAPxptaBlAO7r03cI+pO/dOM0x1P/ogbhbvZlgTT
4P8zB8rv3p6U2nw1dhYqOmWzKY7g9tGZEcZucavWWU2bDYIn+zt8IUcIcNQn5OVc
hgtdJjuETmLGtTU7UVl6fwRtvDt2o86yQ4OWIpX9DIHe3tkGs5PxuilyyiSWWVqK
ol6i4n3h6eqAAUPd7U/nettIDkbk3CYopUCoi5Mb26KytQU2OEWFpFaMmufY2y7c
l2j5RbtyysoDoHsrJ5FEOIELigD9n69eEgPq868BJwWWgycGwnriSUblZ9z/NvWM
0RQH3MUb1XE/RfuLos83o652EVhctm2UZnUpQk1UKfTfID0Ep3P3dGQoBg1l2znk
DUeVaI5IQ/y9Ggl2Xwdea5WQiIBF0itsuYwffMe3yVH76tfsMrjv89GTiABphkzP
mm4G/JpvHaO64E3dQ+ifb/SK8wincM18spRDcRTjdfQvPVECcAIPUMU8n3mKUiEk
JVcFIJpzBjlefsxNYlo0sVsSIH6AQoXZljifa3XKp/5xU7nuNKOADCWOU6WU7sY9
cSuWM4Q/hrr815PMKeFBNxYbMFX2iAQJWdHW7CMOwhQYiq0zS0EsdfPPBtaHozao
5nXvrCg8azhVgrBnga2z3zjetUckXbIR6QsYsHynUxL7WjFrJVzUatTV2uyX6TlT
QEXM4xTc/d9ItHMNhpnytW67tzMOvcCfkt1H5KDK/EGjzfkjw6L2Y3RSiFKKvOXT
FGqawBVSpe8M8945Ns9p2X5pCOtS9z515Iu30j9iF5+0E3zUcdpF7zKDgFrq6lDy
P24+mcHmu/elMlvoa1BrSq2/4TYLiYMtvQz4fxcYJneqzvtM/pa/VDCjQygM3/KB
qN0DGxBSIMZZ40ujxXkunw8DICmV4eluGfhQm+H45hkL7NoJEhaMC7eKiBaW1DsK
qG9Q+d1Pi7VVG/hdL1wJlsWFlOtuFSqMnilfTTSpUYFdR6FZCA95zWAFfC/LPlkx
DJjr7dfbjZNMvOrzCPciBawh3Gg63PQamEFK0XYqw0lhqk7n3IQC/DKkHZJVqdVb
Fm1Jq2oyuNltgs/BeqiYv9D6JXBQG0sUdgCOXY0TeG74wnN6MAHkrGMDiV+V+etw
FJZGWp50PAXmUwTFYlrAwVzRWwAhG6fVcXxuXP6LFHRhlEvNU/kh08jkhyqZVOit
BfaAgJIMbA/+TdLITelXu55FXjKmuUcW+3ZFwFJsF5PnTiHgKP9OmJBCWMwmYPJR
K/yWHuYCH0oumgi5kAoig79riRxTOjTYB1XQs3Fycde20D6uNqboDxpxktTWFPA+
PjgNJX+K6x+krg4vKVv0XC5Xtm6Cd6t3/WNIg1rrMh9arqKHVB6eeOJPp1svEv7t
Rror2C6nIz7bEO4/arFIEb76wAbNW/nDHU3rK6dDGqH2dN6Wu/unTzl7FdC556Wu
oWNwsCPiqdFhSaW8gwkrI8lNhkO7EH1MM7TkyxDHaglQqp8uBZFCWP7BS6DvR8MG
Nc8ENDOz3+P5ODZlmSAkoWmQ7odFynsMeXV3hz8e/9aVCNOUz0VDL+s2ZQYqi4+T
7I2/gZ53KZv2gv9Rjypa6NKI+ou590SMQTwtywHn8pQ3K2LUbVLCIuUAdkYuapTV
qpMqv3vmnp6MuvNA69JtqotaP1UYa1rAjUPXNgaTWY6euT/uk6wmO3zRscpucNM7
e42EW8+xmzv9sRj13zAjfijO8aEfacIGVw4T0HodWMAbPHdQGuWWO/1hnIuiZ8uE
SVnEq2ZmK/CK55UqwFs9dVhI/u0bYYWNjpXEdWRSbxjtj0diutX41kJMxfb4HLK+
7VvxGUA7Zf62L8AYvSdHLCouC1EZvaiSVX+CjF+tGZzLMyVAK29Bk68FH7YSKWrP
JB/m4PN5DESeOW41KyvR6D5/F5+HVxCaz1s6WI+W4gZ4vnZLQQOfuy0d9qb4eZXY
VvWiqNokUf7aKLwWO2wGUoW06yZYuqLTe1dKQ5wyVhyUtB8T61OCXXcJrS0MPB1Z
0I9sI88uIDycR/pV74US52JMQhF40RQYGvm3bKQtlK2q4lzsuEfElT1BuhqOIH0V
V6qkUUHC1B2UBDymfu1UllaWY0TdCw1PkU6utRoHhDmxlYU3oXF1EGieYEgRsFM3
sTBbtIlt+Um8qH6wQcWHo/mGxTPtcFGMoqM9vlwx4SurlHzfCjW5MNKgZYYvECkO
EJL33yP5WqFWfNAXj09t3IuzGqkm9Pkq3kQiT5+KOll/p+e7pWUv9VjoABPTN21q
lmBVea/6YOGY6mXmaEQ0Hr1PrE0WgXow6/qgCPyRf7MlHO3p8o1Z4vaCegV5tLPy
Ig/fOX5iyW/dI+xnnDcdQmZZthfMDBRPICi8HNX4T9lw/5/HR6bxbb9OKb53m6Sw
JYqUMBpsHWl5EUH6x6bS5Ife3dRhsc+QvGe+iroDehLgWS/Q+fF35FFlgkQm+lqD
Hj4PKrDaKZrHBDNvnYwY9JG2aBUbrK3x2s4BhuiLuyas4mUn8Ywry4XGQwRBMgm4
Dc7ThzmU45N08sLhZKqj9QwRwpFtt8GyK2aDDeTNNh/vYkbSCPa4qpsq55DqikG7
OhFpmBZ1hdapvPnz2JlqIgxWvtGv5mXzt5nPqPAXSJg5WT52MtJHjIqz4H1cmfhp
3vvHul5zLhrdjcx4KTjHAQnm8pJME4/VANhrF5Q4ss8t5QzSrzf6B4l0wOeNeneu
ys2mU7/lv1VvS2Dxqau/8BoWD6Vc6xPVVGHjQ8IiDgivxk3T9rAF7i+ORtctdap1
5zE3iZbeKrUainT9QGbddQQCdaCmqElaUebYTtTQTlWixj+GZZbx7JZ7JYM7L5hF
hkvojeA4BmIcE3veViNtPl+XZfeUs93WveUdAGmPlEIsWkyJeBWLnv1eQog/Qiu4
gZqwn9IMb26uXUdOm73h3njbGPvA6zyrrpMa7GS2BBztJ7XYP5iLB4quW0uhQIca
rnoeqbdy4/ZTuTqD4GAn+yQTNuAh8wvaiyDH7m7ntJu92AX1IeHwHr/3QwKFnS1Q
PRh9yod2j24boJrMT3JkMqZNulkMlMlD4QWq4SidNnaZFB13BL/ijGFFIB8XJyBw
5kxZeChScv9WbairGo046NoSKhOU8kvJ9EJ5E3TiA6s6sc7ap3kJCJENMMFe6Xt9
3WLnlfwskYr97o0B5pi+DflBSI90nD9ra8dkbRLwU1F/A3Qfpr2pWKI6UHMUIPQ1
EpR7/RtGWlshaB9F2oIrbi5xkp6IzcJnNAcdT4ojxhrPQvixn+qa8TDW92Fp+i56
TI0T2h0g+rhm5QNGWZ9nQzcLeaaQLKnBalCv4gCLrxYb/bPRzeSg3TmZykHGZ2Pn
kBWGe0vdlBrVFOKzcwxgiWyNbkyqvtsHtfzpbqWLMYvApesnvKjpxipgMWzBWEd3
J/J5TnXY251fLXOqAFOKrsAB+I+Ijrpb/LVtXej9msKU73jtQX9Jp1y99y7NQ1jZ
yX9iHzJFLo0Qa1jTYDWJvm4FqBWW3OJX4piNTG9/hTmWNqOTmckBsWcOrLbvXa6g
kpYzy6STWIrXw/PipdXcuFWiXi+U8N/U5eUhXpVdDo7Gvov4OqcJI/7U+uhZrdlm
bA3OSNHCFfUozLm7z4DYqzhxazCyfWJvJ0L5kX2FNlYL8I7VA7Xwa7Y3FCloUj1p
6qnF3lz278DrQMyufTwiuzX+pIF77LVBY8E53K0STzdIE4LMOGrgugY2NtePEfy1
YHG0Z/Mxco9UCxjvsjNYVEiceVHKLkt03ybQmmq50S95gIWgq9DOdSOcZcjFUkmG
0hU99mI22efQ76vHNHIq8kIssGjQsPTWr5nSvbBXdLQ0YCDXCbPsBgTqHlYR+7GH
WeHSSWgf1ehIPHcSdm6CxTV0kxxfYMWFtk1q2+dOh88Kv7QFneaHfNy9SdlK6K+4
1nIHUGN9+JEza4++w/ClH1hxdb1Ir7KkVeOKoAkLuBh0Qjh6rGmiVJU5VfAPjQ7x
GRE6pYHIa0B9zWbXJqqKgt+zm+1CHCtjSv3rpbJ6Dv5fts+4p32s7YLDPE2Ma7xt
AdJHMqiMADn/LA12t45xM6NTplJTktY1QTK8iHVUiyuBwtBlf/Lkuh3ksTjUEMyp
+LMYNAY4XinhgWNLpKj1irLXWIsRnvingruTkzgJJUgCrylHpKo565Y6+7VC+SwQ
7ipmwB6khh2T8ATaIgWJhVjjDigfp4amvuPaQfcW+NTCWFtEH7qNTxuV8DJI4oEH
CpesuDv+bI5fqXS7c4Ft4ozGYpScSbbZ73euEO+5fneQv8mzJh6T9FBWOL7lKOZx
XAUavHjEJxr9Le3py+lPix9OlWyhyXRu5xaJdCDSHwX1bCjvpLTCqJqnZo5rGJY+
zjwsqmfxhCMCTxmc/9LU/426HEnStx8PKYABo2/bfzmENFigbI7DFMB1EyDX2u8P
F0No1Pqfchjyu5F8CwAjcoc+ced5d2dzjf+HPaNUjsTOiUGdn1xUYKFo4CvfG6aW
2aRFtXwaEegbLIkH2Ao2xNxnZNzT+inalG3hxGLsK0wlrvhXG0lw0BroF9v2f5Ju
2P4a40YHPYi/QTcwBOySMv7D3XuoIf5IB23UmND3Cr8UctxjrhuNMfapOAkuYRMI
8Wl+brn1pFjRuE83O7djY6CZkNYyS+/pE0evNZIvnLahWtbazTAGQN3Vu+K4AQbJ
wfkfgl0Qj+hce+sKtj2t2ytKsfcO9KxOhdRn6hJW3KFdJLZ5cVnqUcXhdEKgyHqL
OiHKLIyDj0rBxlAp2OrGqTupssgo7ZZrO9aDTN6SwsSpe3Gd9l6DFkrpHENp3jK0
6CDga5h/70Keobe/essH4ZMbTxvjwohGvpQ09iEqM63IAxWGuoU1UFsKEU59lmok
jf81Xfg/OZM3IKRTO0YQuhyzUHvRY0v2ec7qeBhXP9KYuYcoAfOgTAUOZ8cZ6My6
EbqwJ66+epjWsQqGXX+sh72+8IikKCA1r9c7lcOkLUYXtcR126tlSrw9qEZrF60+
YLqZY/eBOAnVJqTswvr9Bjd5eZ1UGMWsnnViGNHPkmjuPHj3L+6He2s2PEEJgdfE
gx1sytUVnyvVIODseuyspFKT0CsGnFY+jG8bWcc1vDj49qZl2eks8e3cxaU54uJG
MRCjyW+r4hc277scv4gQCduRc1X/mL5aiVDh75S65bgGL4PcNAvyeQCDPWMfez50
SLMssNOAM2oi6thfhQjnNAvFvXoEGJj8maRraWPkRt85FSt1Cx3Ou9fkax8LrdGO
Oau99D3EDGcFdZpGv7t8nXX6iJTLqcsw+xphtQSQeLYG/xiIjIRQOiYhamD3fhSc
UTB2wT3VhXz95JcMVeIR0zQVwYzvSrqKq1GaYVzd6a+mgnImfPx8G7k3XaPtlaTN
u78cJuMjyVKQaekVPl82m+rSU1oCofQJW6njaXm++T/jJC8+rrZ38qa3M7B1vDsd
QMdj2vOm6oPfm+YckCfTUk/6gyPcPzSeZCOGuF8fb/ChOAM7QQaBDuiwGqjqg10d
0F7E5HyaLUxWs/w4Z8OkY7c5rWmgkdPytAeXTABx7/vyTrCirMO0GteRc8TK0QVd
mIzJ93QrIC/7k0hPMU/DUInrX4ybTx8oNrvHb+dAz+XYxRRWchX4dfs0ZBnqxaWN
APEgW8xC/SyT+UjqiiKnH4IWzUUlZlq1KaysksSbeZ1uvAsh0rBuDYpSaa8js7JP
W9cNTVnId4ULEK0XiTFrFFwJFzAwjosyMsETlG843SNgRFg5XNN3+RPq+rMm0PM3
33iqNOtRVHbpgsT5TLZs9KTWEWDqaJr2JixYD4ld3bK8MGaeje3xoyDXzUlzXzum
g0Y5M5Gj4+DeAvF/WE34tF6sWn0I9/V/mceA53nxVimWlgqPswLmjEppmlx360Iv
ETpFsNEPIIuXrW+DcJahG4EcDmej12YOx/oVmaHzvtiBbK7UeM4h9NYlzee/9TN+
OAn5kyB4EfryoN/vFGr2Pq+36T9E37QaV6z7nlxK8ZCK8ECbtHKSfYNMHxtCXxBl
eVGA9LcC3vZUD8KakWtMw8OouaXBTGNHLzaPdS8PAJQcvNvJTYWKdp4xWFaig/M4
/8g83U6C+zalfU7Zo01W44V31lZrRUhVV3r3AlQRaMHkFNCzOKIMFSnG8meg9EBz
piso986sa2y2t6ak7LSdlX47MNs+QQilJCZT/JXRF8u8PPBjCJvpNpaJOlOkj0qq
L9Ro4LgRr7wn4J+CRxDqFdxW6jb9sFJitKSoAUl8tzQtJghBX7JLxrwzpE6cuM0h
PooX+5g2gy2PIcHX8JFmmTiOMAYeiv7hiKjQIxMVGc4TBezklqnbWsMjPK7zYcI3
nucOqlIrjLW7L/7Xi6um7dvdX23EBXgBTM4kULzetQk+1JxhVEqI3M3rV06DBvCA
POnRFP91x/YHTgzOKdWBE1Xzr6IXB2WnI7GAD3QGXtNDavgSvozBOd4NLDEYEslv
rJwLONHQtT2Eyf3kZkj/x1EdiXeS2iFN+RSywbbbmBpJ+hj/dmamTBRw6APnDYwE
9EgYZXFReRCwRJ1+rZ+zVwNJzqK6gc3hUn0gbz7rjCR4ImNGuYAn0YUHBXJVB3r+
W7uWdIIaclBZQfLzo3SJC+iJxJxw8DBE424NRwNsRaAlvVVbiwK9mzOewyrfI3qv
Wm8jjsywrTPoWg14ChFMJ14bduZPdqgYKkiGmh9BSg+OtWqYshFEptjXSQ9TZyEZ
Imt5cVRsnXA9QvdLN+D7WEz7JGS45Mj3FONQdKdGnazxrvD9g0O+95tOn/BM0HNe
vSus+wiSDHL2RwsgL4pTDyLeZxPuQYaERbgvoA6KIyt+muNMwkCvROTEWUBV2z6Q
iBlOwWPCMNz8fPEP/cQ3BMucLdwyxpWa7NbOFnj6iGiWWLxsvpPw7HNsvDhFz210
xVR30KGS3w4sAF2GGUcATFHpjYCa/bGd1x6svxD7ffAJeGOzdK4Q7fbx2oG5R8T/
KxXvr7CF8Xn4clWN3BFvAEYjnbh6jpFXpEc21/tZTegPD6MW8LiPg/v3BrMOB3Vw
DA5kBoIXKtXYoEfCVpJ4eoqplGQKTJN28XTDrgoVQEX6ht/V0W9dfJlCH0FaCjNE
TVFjsh3RsN/RO+7KSz5JFzpSYnA+qfz4n4RCZZ3SxnvIv2HjAltt4GBE3GZUACk2
xJF5kfVTpjD29HJ4jt0PzNKoTs4PIuldwRfkboogXjZKhDQKkNpRVdGgMEoyvPQR
ROVXNqJyn2BArD2V5ga7aOlpD+AhH9yRxd6+7EiaRqJepYmOZ3jNlWAUwRLCdnKH
SsgyAXoyVi5mjTGVabvaDO7jN9pKScs1EJkALoTHX7YD+TvK0n7Iy9ikfKJPsE3E
e3ofmSmEseTidlSqCoTPRIKrQHWQ48GtaiQ2Y5Atz7vWi/+ckPDDSklzQQFxeejd
3XDxql7usq1nYAWPLGVf9Qb/3nTWO5Xu0EUn56NWfkMrjNC2QCfjBF4QxyJvN1mL
nWObPOkdiBck6vTvgE1DP36DewjVasp/ozx4Vh1qBU5Eb+Vuc5VAfeGj1PU/Uyd2
vWfBnp9gFwneLOAg0UQUeoP01SBnYfmwFz0e3sJUV9hIc9xxm0q81p36NaCUtR6K
ZnrfC5cqCMPqbka/wzZknFoOBbxyUBN1RVC+Z2oo9SYPYjvSaXrgue8LEP+GZqmK
m3CwNaCVyWOzFSNkAA8Fogd0xbfc4kjbN8WezoG1lRExy8KUjObzb2xrEAeV06Yu
Ao8sVqU5xWmcrofEl2cM3m3EDJ4CcMXQcCVuBOcEoyIFzyZmHA9H2JHGO6ZOxGPa
/vnD1nfDyz8z05CirJZcVpqa6Kdz2MvN4ymdVm19vjlvQ4aVy9LiydZMbdwpakil
Xn7cis9Gomvln/nKTKcg5dhlW+js9gVs7pkQFJmxzBgmUvX16BtjZhW/b9qc1GGO
u8fjwOumRSB7939HyuBuvbTtWCpeLawgcJOXW+fj7oW0ho+WObd0QiN+Vcra/kV8
2PXGt/7R6C2IjAOHLdx4GS5Q1bNPta6vzGwEY8QaTiQohOPmm9lb8ORFR72D3p40
nVrPTTNYEATCdnYECsO+25DgvbhDhdUgWVa6gnmCIJkcMst7w63acpx/ASWxn2pq
IElJoD4QvyTVtiL9bjyPFYDq3K6RDuVc9UyYY7xOYMiRSePKIKorU5E3ShjIZAAK
uA8qC+Sc4w3gVV871aUXFKq+7dgjOgDJ/MHC5IHYNkSzdNwvUveeB9cWN2vEjdMf
lMBh8y4peEY5nYWoFDB+B7DaFVjwOughfP3Hjk2ym83WA5SGDXbBOSFjOQF6GZtk
1+A3i+vD7PTJDz4PT7+47JMQgNwL1weRbkL4T6P974HJr3uI4CewKJugkF9dIw4E
TqwPF6zvwcXNHrpIywyOLHdwjNvqZh8Qoecnw3Lp38v+n/4D9fnSTZY8nnlWQ976
iTFnNl2HEzSMiABq/3JKfpWtzn0gC5WmpkdibajcczkjFAQv7Ivaxw8HOJ0u2zQD
JDjb3saPG8rTkFOuvcF/L1/Uz7Z9FNp3GML+IqPxs/G80XzqkDe98jxsiBC3tJL9
XTckIuI+zbTrqDWHLglNJPiAr8FIN18KBvzn7LrhaeA5ohA0ryVbYu/anm9lztOA
ec0iMt4KkLyUlybsrcSOHcJagdNlmwniASGUrE8oQKG7Ub/vAKgFvRc3br32uSBc
A0Do5yrliY1dzDpYgxc2Wr64DcitAn+pN6eeoW40nDBCjmge/wJTZP7IduDlDEpo
XrpSO7vH2GxiJFndzdv9wbUz/eBhUFjV3hthXDzF4MuXG7U0acAMTXmib6nk5eTN
Z+gEOtcUqYso7NkqktnPu7jOBOziLoVIJO6Wn3cf4QyLopbGffKSJbcx1mJ64Y87
nVjvrfyCbZgI5jnhJ66KcZnBi3Jxp7/PejezFOqPlcjP+IULsKVwvg5jUa2u3Wk0
b4V4D5wlX67hQ4rAkFF2Ub16Kc4bcqlUFX3VXiO+4btPCOrNACfXHYb1zGYkh/Rn
eyaNNdE97tZy00Ds/3r5l/EHo4TOpejWtxm6ox+TyDc3Bg+0SiW2Mq1gB37xrau3
hP//Mat52NRjOTglcoXWTF8rdMD1UPKBbz2CdjIj+UnkwnIaMSL6/naFljho/ziz
d2ensK5fbnoRP+TBUM2vr2+w78rkm4KQo0pPVp/OBuyfXg73fHheD0HmYr4oVIsf
GYVH0Zpt8+MdgjlPI385IetK0nMqdYZZxd3dTCgAywraXLfX7mSs3uw9Q5auVICT
nTlX/mxpOWUSiDiMvOH/vKSah8FqHXUG1ZxwRKDAJjRtWjLAciK3WON3RApzypHO
EI/1Tng5VLpIUeI6NdRUcJc6JiCvN+1o+mklqNy6KNdpIHyQE+rjQDNORPrOFX0h
Nb+qasCHr3VO0dapOuKm/AZMu7okBzdRGwn2DzbAwL5my48bnj5tO4ps8DbQfGvl
BKOhmsSgQimcnSM/cMymHAKrdGsFFEvZdYb5TClYPJ780WnCPorIKvd2w67ClnP1
Fx7vy0Ws6CYeASo+XXBhqrJEx29CISBrIQyiWVM8ORRiq0kQ6huH/rstnFXu77kw
4qWI3BLoaaJqKPcYPp0eRlN7nGG9tF9jr+9QrzFzGZvuQB+cg6XJh7EmengGoUn1
g6RLOJvxLh/tqILAVEzCK6tM9NNknLfyEFEAx+2WM1W4iRtFxp3jgdACKA1DksjA
UlgU48BHpt+tSrN15HWUf2g8c+JosD3fTKy3MwM3JzAMtQJjW2x3DVhfakaGhLb8
eKHZmCTiuhjlm4E40NlsqWrYYnGFzdzL+xrFLmYS9ADb23PVoB3j+D8fpBLXvERF
J0Nu+mVmzHjcITLYPLmrtb/zINkYM03yooeAJEma5ia356oSJ2CakIsHnkJ0akZZ
rVplflZYEt6+oEO/WQv8Zv737ITo2ergTTdPSsIHgvfJPPQwPK1lL3y77VZ4iMnA
qJY6NWl3Fwc23UqS7pA1OtFIaTGViNkxb95/qZg2J0EdlQf/jL5XVHRWWemhI4F+
/8Lxo8UIYi5VZKPQuDbcUkEgSLEaTh2LnDdQExMKswltfo21rEwd4pR2f/EKj0rT
Ks7j8D9BZy5oirnFBrTy7Xh6Fyu4LDm93QZw7SI/bKfIHLTxo06sg6rCoHElCWrT
fNMc0i34z3dpHqvVq9R98fCj4Pe+8Su9g+fh28uoglrRZt8jK/qMCvb2Stg9dHgy
F12WExw6A2n3kdB3Ivfo+56pOQnbhpwAMj/C6pzB8dtzKgdAN8VNUzVw9AsN460g
8FISFTT/GPSTOD5HWhQbR3Pm7Ep1ZgkKiV3EnkefeJb5UR7xms5BzFEMPCVi/GTk
DyaAKrcsInzgGmFnR9UGqYvCKXjO3upEPCPgSkfIFmfd68qiHNcYNtsH+G/be1ry
o0v0Lob2Z71joeNaBn2HA7OT4R34dlippIvFa2gJs4hBJZdKwREbgnZjlf+r2fTN
g6NITLaOGn+CDdDBiOQa3+ja49b8r5U+UDoqN/OqG9qjB+vSZ40oHxa/pjfPxfL9
QxkEyXKjmrwoMtBOxOVRXR3p1tG98BJwSbJ0enwBFSLlZ+1ldg/VPDcqANXxmGp4
YmdzHC/KPiAwcoyn61pH+J6KOh9IwbrSqG0oGIhSHLFkvLyhSey62Oo0Repj9Uw9
7xxjZ/xBoDrV2nVcfUTs78yd4+E+oE7UPO+0BDt6rA4niu1I3Sij1NAO9E6br8h0
DfQld07pmIbcQPnAIqIDaPX4+rrovN3EmNM/AxeJhZvzqoi3Ma0NliY+sh3e66xM
DSDEYXPWW/2ABFc5pcs7loBEiC4m5Fgx3qeeLC0tl5rGyPvHE/KljxK8/7/iBBPf
qVfb6X91+3DieN+NSmZCvn+/kap7lljs5kXIJ1KLCXG8w0ii0kZPrOTfzC1P2pmF
OieuGB9MdM+SNxHKKAAQWH5agLzRQ0sf0CgRGRF7TX8qN0LnmZyYRspSe5wIwvzk
HwqqyJhb3QKDuA05DXNihQpkc4pdVIxwGzhYpaBDdWS1MsKMgZ5Qd2aJ8EnUo/z7
F/Ee38DKGrtzAEsnNOsQNbw4DTd/uOaiG7uRfBw9THwASl6dEJ3wxe5S/pJXDS0M
uHNxv57QTMNpzNUq5uM83VTCM0EwuJTzw19nWdmmnFtKyafYxwOtddo0A74lzLFS
HgR6tgcdUUdW4Cx0X0GwrIyL8sl8EytYYltZosXXddtUdwuCVsFzHCBIy5tjzibZ
pmLFJ+mfVjiFNU2VVd3QvUEqWvcAOyXeQ0E+fV+JqxsKXhJ86I2yWvebC2uk3kgb
E/E8geneqWdfPeUZkzOGva6LYXlPJPqJgzWl9vElSwAaTtPbPLlAdT1ThPNTUCR9
cBoQdpnX2rrpZ5wpksphD9R2D3TriswLJBM1ZdRXZ+vfA2wzY6rQ/b0Nw959n2xL
LGiyp3zWWO/CG5hjnTyOn6T2Fo+wrOJgQkljZAlH0+yUWHyUw/a7gwmEkkhu2zX3
yfYRmYOCBo8d3IhR3ugEtPIs0ByFr46KgRxg5ATrWOPsXnMvEC680n8RXtKidsaP
sgh1F2oKBiGLRo2/tYFeRzIoNCQKMHfe64lzy0KYVbAFyaeOyFximBmvePH2VfNO
ynKp9Jk/bJ7gJI3gGRh4AOEZGj8ynP6vuXEA3JZE+XkmqgQW7f/Ya+EWojcep++v
+xQ8I5xDireQOyehiHIcN4XIN2o1KWK/omlg9ziiBtm1eOAmvAtxc8IJ39amN2W/
iP3Vk9OArxFH6t3m9Dc14UI4Y4Zoo/KPtt/ywGK9vmT7b4rhyHF4fzakhbe687Fy
PaU7DVUSoiaREiaf54q6HlltehMQ/o1Pt5WbhAZ8fiwst+UUJwRBAU8yGlrJjhsV
uArdR7VH67zUiqYAMU/ZyLi3rwqIcvc7z6rsjBcR4esCgu58Sdh605bgRCIKeRch
NPx3S51aNZaoix8V7IYQMq+4KQ4WoZH8APd6vJa/7tEmLYM9MIarp7lHz61W8pPe
2AcbCSrlxWymNJ0Nx0IxPdququImowLj/1L4z/Bo2tLzNXQbbxhD+75EqlN3tl75
G0i59+I+fYM6CyRxaOFkDwAVEZLPqSZrhMFGwyMQaXb0kEYTA0CNV20mHv//hKgo
80F+YNSC1mFVdviGQfI/jUiErZoHO/dGgrPc/x5/E0q15k56KSl0P6D0cg6Vn/6R
H8BNShDQ6Lw8GP+L195JpTpBAWD2hWO3cptNQ7uxf8KvDMbOvO9mWGOTaYXK80gM
OW9k9pVX2SBH+mbRWt/kQVhGdxUAYDPn8pqm+Qkj9quaM+xHcQl7kH532sM11z+q
p1XAx61DtXs9r1KPHRucpY4Jv3lJJw7RWxTT1e/pNQyugbannOcQxLYV0dDQefB0
c7B4FwknDEStlv/PJp3fwOGAyiiKguUramLU0p5T0Yq+Sou1pPQyTgoPO8yPMcQd
C7aygXoPu2M0hnXoxsigSUgc+awNcVqEe/GswFmFQmo/e2S11v6PBSGmOHmBDYKH
wVVC+wVEF5WibNhN+J5sI4NCSckefBMkDfm0PiU9ArecRRObuez/8Elh0ledR0vM
9Pq+eVIJ6uuE56VVA/TUSsMyTekkAVCe++Kl1ZU8VlSgDGvC/hb7l/Qfah/CpxIQ
kAdf+gl0P2waK9cXo11OjuME13iqYmuAKo6csGVW6ip+Kj9XmVNjhv9Cm8fgL2Ud
696931hNk7Bejgg02oZe+AdeZsixixewLZ2FU/53N2dsUP13d34LS4BEhOoFSIbj
+fCKbfTlSDQBXP1tf3ul7dV+7KLo55CtP3fdIX8r7PjRbQDE8DVNGqBBd8vrnvoZ
4pyrvHujlco8OPX3jvnKGGtos6MoI+RHT2GzUTKFSY8PwMlTqu/mAKWZ0KeT8NLi
rbyIPXQL1DLYftTkeixhYqduFBkvk94PMnYTzL0k1PJRnfuRqyUKz7INrLN4wO0I
sRiPEOfThb+prqh5Th5U89C8FnMPwYNLB65F75vQ1NhjI7vir0veeYVtgDqq0UGw
bHGqvSNOCwpDvDy4bK/MXl8DT57/XBUdrZKgGnagIGB4KMT807L30tMINAc9Ob3M
nLKIBIppr/KbOLSPpQ1sudXgQzUP9ojhSniVhhPzYWXVv37xrkBxjZTeNN5z+N2a
J+dmhBDFSnhvPPEQSoUcrS5NzpvNGPrSNwLduXkmW5ZMG9S0IyyIP/Cgfv+TbKRJ
UTZI6f0UHKBC61IM051liku+jmTZOIPbTwfoFn+xx6Ih03FZxXbL1j4zGA/qtdr0
ceqpH3dpcfLDIx/UKcEz1+QgBqyMSGnJyo6cQNWnaLxeKIII+4mE0GI4p/Oe2/7x
hoMca89SfIResr8RGJW6IXBzA7DU8CizzLLVaLYS838BVwHezqnRo273jVTU5J4Y
8bFHZ7t1dyFJQfQYEGjZeM7t+5DTC8LuCfC5RMS3Y+XNCV0I/EqJ1qrIoCsKajuS
Tr21E+zcPyGnGwota6ELUS8Bp1+QAVT548tOUjQgGipX7CFvobWJo7mbRUQLnZ6i
/4wKNCegp3w9hfmoVLSwS/9qXXdyiVjctqzl5OcQhpJLnnukHKl6WSPhrh9+SNZm
NCIGaa+qDegdigGAV4LmqCOsHq6QSALHXaNuqlvsf+czZ8wVn4ceA193ATjm4eMO
YHarlP1zLH4m9NJbd/vLRqQ7wOO/5kE8t7qXRLjjPWhGabDCKTgcXfwjzTQ1fBP6
dfTZCdfDQESe3/uH4+SX4DxUFbrRqaumo0PjRR17MP+q9ssSGUaQBa8XxYdv5eSf
G7nmZJ9OZO01mM1ourPbA4E1b6Z8p/fYb8zunRZ4HpxuQrdXo81l1RlxZ7RmU5tX
G6vH03VnlnL3ZSWQpsr8mkZXk5M93JeQuk8ty/nfMaWOM8nSoCyNuDljkuj4y2Z0
Mvk9Vn2/9Y8aP7jNyCA3R6aBkClVKCBsn/KPR+AY/uKYAyrLSPTTC1wk5c0jWJ5m
ANPvO8vX4iQSzxV5xLlnEr4aPsPmw2QCsd6hwAtFqhXhwHx0OSTpK2jzddYt7/u/
3q09+jtIdrMUzjpFOlJXH0qSvAbkVj6XyQEsHqE31jyLL1IRnwqWalNrT7pFWWd8
xo0rxsCgIVxZ0FhGiq/Dsjb2TjR7o931SU3zOs4OlbjBeewBp5FaPJqFCNKm7EhG
xw7aPf7zv/JK6reN4vyGLBKOSTcya8NeWdBZuDT/cXltYSNVP08XiuHTKFGja6Vq
LkOvAFEYnuc5eja4fHwp8oRdUsZSMcCg0UA4ZK4n38x/IyTwBwHOQL0M+zSZ6ust
8NkBDK5ALKSQuhgotXtrCkN9rEdanlyIey8iFlmCinFEzkCGbVIcfmTrzs8JsDBb
ISKA47XUi0hVVeKTe14qtg8pSKTEmLM+2+JDVVIR5nMw78LzW2oXwEHjotv+SoVM
6NbQSuG6yUce6LciG/2u3vj77vXSEIrufbSxwPv2yNq1cW/nZbfusFiVOnmHZZ7p
oz+EuJSsPWLjyV1sNhbSW17uyadrQQVZQ+FOjiNP6C6v5AcOoa+wJ5tJikiSLYY+
xTYKoz1jCQeAYDyrTR8JaMw6UG/Zseng+3vXTDlrtxTTXBK9BJHovJdVB5i/F5lj
4529IyQMRqhmt0de79WQ5o2R2+zPkmRxWNdXgxyTk57q36Ya0tgfIA79YIo5Li24
SIMNza84EB7kS/omR2cSj+IljKEl4atY6NouEZilJPhMhUf9Dc3UKT1socNCTA6o
fysBPtZEq4/WberM+f3VKhrUGaF+tk3OkY5fVH1HsyTVFufyTP0RM6vwRKU+A6D9
bWGfFu8hFdULd37k1PSsk9f2nCwMkki/XiSgpEM9f+HTOTILNg6KJTg3p8+QQ55C
chZFTDP5nGKN4KkhRggQQKb7ZcV7+3tpkSEqpCyJiNP85D5/Rti9qMn1xi00hH9H
dwP1SsNIgSaZLWKwo9DN0hXrOemOjJx3OtsV6HHq+nKABGTjqaf8qwEFNNOvbBIx
KzM/07Vxgj7mKpHhTJumaIk9pGl687KydqhnA8Z5zPo5XFZWwoGpXiAf84R4LHAm
p0dSefHdb/SpEHQquM2A3eaQ2gJhcCNtyhNfyhFUPtRW3qdw/5a8V6A2izGwleg8
fwteC34jhneyoFgJZrtBZj8JRBRI1j1HWcLnSKjWRs6f15PX+3jE+b2dGYNYFB21
0goGVQcJcol55Vm6HjW5tSc03Aj3kQT1gFFQDKmjzcrnwYawuV/rJ8iN8N+kyHuB
8mXfMqy+u307uwUuR3xqVwieenmDfR7ST2TS6SKnz/jVJPttjMtHlrLPb+PrhqDh
u+8+m4P77uAYXXxptizC77xDnnyx1qUyjipMGTjJbcOCIO0eqk1XM9Kr2P7+7Q8h
jL4RH2VtSAI+923arqLrEuuZm8epW05qPrNQCQEsF5rNh27R6ylC3AufiKvSZehw
CCqtxvknIvfuq7JPqCOgBHMwDtdEUdvIBjaxq02/Vvhb0hLYqDgwHfUAci7Jnie/
IQzZ8vmTb+K/hrXFD0E0jNbh0wHbh+sLxULfjYxB1FaknypTIqeWJdr6VWUCM+wy
syB/z3OZkEvUu5g1p8oxhmHfwcYt2kJXL88hlu2mRoQVETcxOiwOQSAHdXLUDdKb
l8U0RZaqe1mACP8A5i0RbgPgXFUe1eIh8PRmrQqOsKHbgEsBDLp13bKc2kWrz00N
bUHsyxrUC3DOXTSe6cknUxqPqXimDaPVM2wXu6wckny5HRBdciQ1rfatUraW4rSI
jvsWL6Sb4BxMiT7jNwOvspZkpUlZsQDlzrENPbprkr8nMquuSnlQGiV+esQOcc+J
sTXIUR5VrOqH6VmLCybw2VZN5WfQqwkc/XiuAYL126SfA+uRlY48+Q83MHEw9Pyr
ym4X8ymcKFshJFaVnoJhdHAHEDgQt2x1PIxRWTmDC4EMmrFai+pgfkcO06wAm4Jm
VAzhKJx7bG2ipZsAbWIlZZurmncXJYucoZPxmsS6qHdLCNQiKbauts72yw8VQkes
CFnNyHZmNsfURj8vYWcb+DsDmaGZB2/TFZRCJyDdKbvUDG8J/pamIrygFV8IBW/K
Ku/IEYqgZDGzlsUCFqIJtm0ARvboa+cDOW+2ncqEOgheaje63/TJF/x9tmUqRo0M
VgTp2psOT0KJoteywbkOx5yy5VM3sNhqDwjjdFKeY1NpOzNitQay3lNFYdwZOVvw
JaIbWbxlRo9bks4b8BTerK4wRElUveIPW5Kp0vA9dQrcPCKa5/bDm8elDJ+jJj/k
rCt5rGMYm/0W7NrzvAqcCL/elsEUmn0uIp1xHIXtJrUkH6+uctSRRPVyw0nl5WOW
m1g3vSAya2fahb75ZiSxNkEXInwAkMkoPXb66q7kam8dKg32jTXTRrxba8Q2+rnF
yjqkm0VQJFDyUEPyDQs59y/MRfUaYmthAoDJvoFwP1Z9pXKLKs/9Q5ildsmy12Mq
I3L0LzOzgVEZm4FlJj1/GqT+Jdh/4kjkZIZ7/XqbgZCWkj0GQFNUeg6DPXOjLyAY
2yRXufLTb473PagTmwuIHb3+mUp63QoWthgxOcCzMDpXNDXBv/t55lOeZxd3S8Dp
/qJRz0vaBuMnulF8ALv3zZtCf+SJInT4+oHHyZzwEojREMAItMZsRcZks639P8BK
sQlyG6Wru9xB6oeXFTJzJTI5+7hOCwUAjT/XaIB2DkKs9TUEcTKYOOb7nahY7wxU
QMC8z3pahq+XljeQgj31dMSna+z3KxwRN7KzbJenX8wXGTrMPN7coBvX+53xA4GM
h4z2Vd+24hM/DYR0iU90XLaaXUDSbNU8zyVpxLUkT3PpcqCM4PXrkVqAeN5FDyIo
FnH9W3bP539/98fTajsktq5kwXDMXLokmNuA6U0euvJB6goatv3+InLAQN0XPIpM
RpVmHB3wnCQYqkQMn9uOQEBO+TDokwfPJE20deqCxdoAoi3ZOL/2gxAhqemhJn+A
HTjeLMWIvsFhelhLOOSIC1nio4PKOsl77rFk156Sey9QmO7Lsxr6da9F0E1Va/fA
sV29spnp8gq8Mwac909UiPBBnqNSpCz7RwQlcmY0ujoSgRi2B3XpiIqEX/vSyuFW
OkJVqWxJWyQcPAPC6MzMtqRFXEIiTAt/9I7ELZ7huIZuWPi+LzypEz3mbB4IZgV0
GIOA5pGXsHfaul4427OAO+ZWDPBOBf94TClH/J+bhQ6VKqsakdI35mC3psilVtXI
o21+KQe/Yo8Hyzk+9rCGbXfuyB/hkj24TOg08+XkufCP32p3CpXbqgAfcoaULcu3
NPOeKMRBgw1gd3ZAv7qqa6iNNihoVsuetTbmHpTuCAM/7hVOQR7gwrtQprXKTxsM
nZ3FZK9Y53AXy6SrVhq/W8LKho7mul7LnFT0j+tD6yNsmLS0q3D19VfaetcqdjPC
CxN0ARRwkQDVWFTaabeoTXVelcm+gbn83o2Fg+q/fjsZexTzn7PFpaIf0HfnBoMi
NQpSrrwTJfut82LUrTqdJt50tIcFGhjWBJGdH+J9liviUtvyHEtynkL0j+rWjPtN
mloSzNgryw6YWuGczyMzs85N2sD0D3rPqjb+cSdg6LD8nVp3ZlxSOM6hhJUZxTlo
AQsaEfzWbXIflpaTIPbN7cTtHD7DopdswpesqvoTd/phuN6SZaYrdKT3MDQOZ5yK
Q4NW8FRE6JY5o7RzDpUKFrDvaXOpyYj8y0deyCPOOYsbBcEG5XmRUPGzikrS7mk/
Y0hj3tLT5q+bqUjOc4jk3ePH5OkI0FTxREToAMJKVcBkdZAd3px9+4A8qp1gxaHF
Z4/Ody3bGYQBMrMsXcBdpV4nrzEWiNup99y/72YJfgJ/0qVg8cNAwZ18JN0/5tAA
wnV5MgNqSrWRVk0IwxcOrdjIXVgCd+3Ptop6zsCsXjE7L07B9auAJlk+J+xSx/mU
bCognElGaJlupBgVRFmFlk0fRnudF9OsSA3Zwqd7j6N60xGYuGKwLMjy7X9Yq8UX
QN5HzuzuVvMwI54yEXsMNGWbcq5EJ/LpHHam6pI/FHI1f3CYVlm92YNDyTfzykrG
JosXiaIpGaCkW5P8JQMzHLGaX6ud8Tu6dy7RF3lsU9geT7WIyuCw9FgSZY3fWy7e
A6n6UmPqyRpAua0z2C/p3090H1qKCpPUs5rwxFUNEtoHPj4hLVzJoZv0slz3T8D+
X6cd8zpq7U89RAefm0lNT22YlnRlyXioFldXJk/x41AG96aeAQVxqHoYRtB+q20W
Rcca9UkuC3YXtTClifYWH10fqRJgeeHzYE51SVQ212urG/yHVkZ838962mNFNvhT
7nxXRbVkBMP7+yqPQm81iGoxd8a2FC1M8IP8qxel5/jeXduFy1qKjRcxy4B0uYCQ
HeOqWpK9kWEk76EW2Br5HLfthD+0kJqVUl5KIjrLVMXswM2PCs4Ri3cYgIyalBoL
+X1O6HN77ot4o5cmjWX1H5v9Tw9JUUDfnzN4NfE1ngJBLZTiS9PyWAlt2b9Uk/60
QSRVUjDHEzxA7MhX23A+vwd3qzOKBRFoq11tnBVQXLVObRrgUE4QfvI8Y3XxMPKi
hohwo2yjSxXP7tU7JVCn8gZ8lgn2uE1TQI8TPEokT/tE4Fq3E+2toUfEQ6DTKB+r
2U4yp8ioNXy+Tce01X1K4aP+2YsN+GmZbjzCBB1Znb0lNF3fN51Vkn9mgdpdfA0l
b9k5F2ifUnUpAryxrvzFkMyKRI7oVjCkFynlaN9iQeNRcZsseVdrvjaVXLAFHQ8B
hwEqSrRMwFaMzsH1LiI040cBLGde9sJrBYN94lY4SWIGmDhTD6lXP0p/Av1ksYfK
ZJdH0GomrPZP4c2XYr5TIQCg5BeQSaiB17+GjdBpos+mCweEGdL1OdqJgSpyTajb
yiux+mjSWE9cQRLVAXZDBuzD45iJnHipB3tet1DUZbhX9HSvYWiYTZG2oW9W0pzo
wodTMPWWyDqpH1YmdxxrwDNjpJbTVMcSCX3/1ilnqotkM0Uy7zULYuDmunD38oiB
Gd9vsHVu62yzWeraEm3XQtgzp5KHLjZZJusntm/p/cO+wzoREZPCBZ1spJv5heeF
VRIQkWU/k6gkyHDp2WxFOuASZUf8Fb6N3k04zWxKm/AGR0W+mGiOIOa451EcZkXq
U0Z8glAeIpADcehR/Z5wtcScPlgqG9Fp/ExP7gzsHUAqlBhNu/omSYTcHADnlwG2
/l4qWFWxtOoiyRZWKqTLGwXYKD1BlJASxz3NPeyt1ioWLKKG/Leuis650DH2GrYC
q2H5Q9b/1bX1OzhrvHiqWqZGOsJKeDmvCh+4E7njzT1f+fPJRBwiPZVh3vkfJny5
tPFdQV/gH/jk02CMANvK74zfh8+s32MOfqKdEQ3L/njKBPDMJ/tM8Zo6RsPga/zM
mXxoLqNDuArWIfguyS5LRm2lr3JY+kRPBIbBc7AtEfXtV/dvYa5Eg9zPY22D/zEb
Bi7C5riceffhcXHcbdHPjFM/jRXEIsA+olCOD0/rrezNzxDhYJHoRfS5LYe+nsob
XQZidjO+GxxSi6Im5M0xOweuwvdiWtZzuyGuI34/x65+ZfCpJfObf3uBplFuegmH
4zGTzZo+C/03+Y+FRPH9IHbUF+phqwAsUN+hKgQz3+X/ieS6WQaJqYIKxW0EFRI9
rZ4U59tlYTHQakhCI+qDiph6NKTm0ZXCX7i+Rjgdld276ozRthjCg8C5iCFP0oGj
Yq9x8/w4S6KVgSH0JXeTlP+y1C9BYpxxWP/p+KrT//jen3YNN2FfW0jwj1td/NzB
iYT90MFtf2A/KnlVX8odTEVRe+VJJpwn/IoJfDZkHy8i+9t3OBW5gwN+72M1CqhV
Zx4gz59651Zimko6niKPDTpXhZu1MeCvKQpF0LfH8ciHX6/myZ/oCbyFtnyT5lMl
ijqolnG3IQy8YFnIzrB1HymaOzc5s3mwwaG/hK/ct7oBuxo+Sbxl8z7NlI4ctTG0
Xm9kyGq3tMKYxVuLoO88N9qlfC7zludHgBG6OQWGYoIj4EPl/w2LukQX48kUdyAr
76uOo1VtTMwBX0IdUyc78YP8OPlBbaZCUgIu4L3yi015BD8zxrumqAzFDOmxW+k3
L4ZakgK30a/HpN4boZGp8aeBd3Q15QmQ1ziKoRDkW4R2VMkN/rt5TAZcZr3R2Qqo
xdRL6F0W52Z5/71g7p0Shywb8oOGxz1mYJagSVzu+zaXk2xOKnVrmXMY3rKA+QfF
YclJz8TIYgYrhB4ev7RDV5+vqEi5LUuo7f0dLMpcXvOyViH2yeQcyCb1cYtjqv3F
TtyilGPOobAzVZDVsnJOHKL3HR0H6MuL74keZFVmb6B2FL2Hk36Sj0XX8P3pcsrc
K8tRVAxe0NEzIcp3I+BuAO3IgGb8mqZbi5Ul4q5q/UiSL84WAdjtYfAhTNtMLj4v
uLCL1awA3e7s3hPgozZRIb9j/nTiYowXI9GRM+34F+8tJDDsSvo1abg5z5MFRCms
UNEn598TyLsazAySoUEJ5tYonDHM/4qjEOYAVQhC6T8NXfCg9G41xOmYjK9PlS5o
GxTVXvfKnhukYnO1ZIzbJZAq1bymE8c/z6mWgg+IZXIEfg2vtqBmaqFS9TE8C2w8
TjnqK8K7K6dsnAJ/sN00LR/IHXJS0Hbe/S+zj6M32l/6UqFc91tdq43HTWses4Nx
zAvhNUQRhLEAHQI4PKB6F5n6yuzvjAoDZVQ/V4MurmOvrEhE6qXRmQsyM0bJ2Z8j
xIw5PNjRjueEP03Pi9fvFu+K2Q8F5sKqjpK1rQ+A2CDPD8QqEkFWvJfYclGlN+9e
i2DzaWs8/vC+2AnY/wipLJ4rnCEvLJaDIEXWq5PigB+ESC/V4drI5oKsZhDLZw1S
B6fZT3WGHotxsNPZQf3RXWIH+ZrJQc3ZrUv0Ufu/5aiIjOQJQIVZA2luOdDDmJGK
T+HSv2qXyDEs0VezRBt6Y9khJHQL3XU3ECkE4f/VZLsjDi4d5P3QlTLZwDzly3Cc
7eT8C0FU6uySJT5zhFaSG05UG5auYwDAvFaNDItCodlvmVha5V1JVv++Ipo11p1i
YA/hcMJjhEE7NelJbraizFdWcQTbI39OAm1j+in2IcpdCURFHVr3wOoiYiZunRFw
XJeW4Hk1TGPXdjdqR+H6x00ZUAeMLu8auUvRBX4rlFMVU/GokkNGA4k68Pfh02HB
5saBk/PzBnypIyjmZ42kq6UcWkk+qVugNkAcC0C5Qt2BbN0xIMy5gJS4sfC6YkIj
fQhA9kOiZqOX23WugoHuOZj3Mw4zbX7rAIoCTHqG/jRkswnTJtUtPeNTsic5Yzp+
4oDEUEe+roYXrm+IIWP2sS6rFszNweFJW0k4nmTIa/6LNkTBYe4kVmnUehszs08l
ZDEWpFPbwhybyuQFOH8f2gv9hWTPsL1Wyb/hJHRFcFlasffwp6nRXjGmnk2yWiII
hDje/j+jtAmSaTjtEc6MigMbzPO51WFEUwcKouDo4fVA+VWht4NoD7SoqjsIkFrZ
McbkZo2APnnMt5C5c5bHTcMvUPmqGWiqH49Jgaq2i6j6qIcFE2ClvhQxBcXu9SoN
pyd/vDcyWgUBhi+dfTYeLP+uhB+beh0AJwd+dNqJSSBdjZQV1Ko8bj6VF+M2BZlG
0LCJ2i/YThWP36Lp63EqRmgUosSEZ2wzOqrGj/PMXbBIrwyzLnF7wzNXOs4LN3Ke
jmOXFoA6Cuhdf+WepvM3bbLSpS03exHbbkbuKAwYP/9VQz2B71dB2QqyEZB0lMhh
qg4MmxDjQQsnCl4KQzyZdamgwP/54zMVodaL4B5v6IBHegCaoun/yk6jQzqslC4n
7eVFlWIOF0DArP10ebE3aPY3Dk6VlSw1l0tcLDlWcWgLj8F5NeZbWeKrmb5MYKEJ
Rm87Kl18nZfNXl2e1fqg7GALn9ukiRx6Kai45BQDTqrUNjtecd7r/YT+ixReXZZz
yNsjZ6Vch5l8Xf3z5jVgVE0jEYARhF7RikrljXza8JYMgAurnW/uwwe+GIft4Ndh
h1//GBtDgY6XRIbwsQLTW2/LNIst0HcxthsYvw2rNYgBPyhvfJSMlrgwd4plwEL+
vpThGF7Nf4YqIGQ7qTYgOlfz6tMClto9AKzLWkvvH8MsNuvyL7g3dqYkc42a3Z+w
LKI+49iknZxbelsb8Xom+Qi0OXPZSsQaRLgi1bJktCYJkdPFAjZFJU4onsRmhgeo
PpGNB9TZKFTCmq6csVNS1Fme5tcEoLVWl9D7x/iwHe3u0infojdOAS1nYAW1BjZ8
xfs7QfM9rp14/Gj7jGdY0qVer4V090QH8ouoroQZIWYrknFN4rZcom5SkeNKacA+
hzyY4faP5GseUOIt/MHDDIeuH8S2OSnPir3wrwGlWAdmRoxjHdIHUuAyGXNKo5/a
1pf0o7mR0H9bs3+xW3Snnyl+nWLCQdSlbSap6A0HmKWWn6MjDFodcFr8K+2Gx/Zc
1oIykpe9Co+CHp87lm0zn/MKjw6V83aDGtwH+kJBbs+XTlGwAEhqlhpWjVZ+7CSB
jy/OVMtAavisCqEaWotNDb1EKvM0mMY4INBDWWEoUCZ/UIJepTw9MbmL51fCas3d
o/gy34ABw83Qm+Ua/bJlwPIkYIlVI94s/4Diuv9vgy29aiFOXrkYSK/BPrS/zw5r
wz0oe66g/FMLk8FaojU0bnMKW7UmVkwZgEuL/56qdepS1z62S+wJ944xIZw495oH
KtxJzsqsqbAuTUSXMorm3TSYyTdiYLBeQjxxQEqiOAunYT87ABM1OhPx+3mwen1i
QbYSIMjOhv3tBZ9mn96EychXy3+HIv/fJDhSgX+o2hOJSXe/anFMaxZh6m9hFU2k
ySi/shcQyOC+dYGV16K/M+f2cW9PKh1FlvJ0FNhpsM+L188EtlvhLdv/Y4nZ447y
HJrgGeWh7pP3G04M4sZmlQ17KqkkGR9sF1pGu+LtTyVT761BUTayBV5JYKiVh1ho
qfhk8WMlBVmUd6M1/XS08TGti8w0wcF/yWfQa6jjjxiThYyz4eSEB6A7e40QF922
IJvCgqvc4eZe9uYgWzP1UST/pi57IBJg55s5WIyCseNHKMC12CqLBbxDVJ2tviHM
nnud4ZjKgmHI38krlzV/7sS0yVdmt60oqs1M2ULXkbWmaZzDKm7auSeY6TGXp2f2
KHb8uLlG6GBXHDw9V55/ORqOnLlUlSmvt8i8VtQBzQfQYQdVWZoxNkXJp8FwrHhp
muhK2Z+upmX3jkr5LWESNh8lMdr1lNWvezWlLLLYcLszwvcHOvFXG+GrbnGxhaT5
uE1CewSEQ3FR+ejMBs7WxklWIPJjKK2F0jP0CJJ1J5yZcUiQAwrVPNGtdJKPP0H9
F9vTCBrpkUacm5XIp1s2JcxubwawBJHDgixWhNBdv/BHMEhinf2PFkhfLzTlu3Wp
7peoqucWKvbtNk2rrXKP1y83HNirNEF/jWn+7mgi30vsPXxPzVwimzwBirDmaL9/
PWy2ONSx4tsrV2hr8BIYIJPoW6mJ0C5VFHUnsFtjXjUYIguipN+GRbPpfW852Tps
yza0mhBpmGjedq4Hiczsvz0Nym8pEX7mT3xBvjCq9FyhAO17Bb39dGBmVdo4MShu
ivAgZCPqu+MfoE509ty8ZfkhLBjnJUoxOPZCqpP+Pb6ezAPGQ4UI2LLpF29Am6Nd
RtTcx9DVKbtO6QU3o3hSUbdgszhGzP32einFkG7ftDWAJA/sZf2rWNHcZ4cZkxIT
cEw8AzMZV1tCYypCmNBg60Gpbu+lzYkKUVECdHUvjO98zVYSc84mtd3khZmWU+z5
oySPeCLMkRDYjnDgpuCGnkR7YmM2BgxBd50VRxF3EBNpK7f0dIbr2tHrJ5T6ec11
jMcxHeSdpWaZBMT+jc0pAagehY7ycCWOMsCFkd/4VnGBbFeeHz3K38GO0ggpJ430
A64Px2XtJkaJ8pHWewy+9SdWwU44N6uG+IZj5KCia7UcKyL3WP5VtIHZt0AofxZW
L/LOa+UpWhHxWGAfpYFUXAZbCRImplUrtis3N7gPlMw7L2SnZjhyE7Gog0PJOOFs
bGaK4KARWya7nwYXHcu2ewTtMx6jHmuUUhR+2c2sGUiezrtUjofqm2NLvgDsNEwS
U2/Pbv64Wbn3CawX4gBRTZQ9hGAG8XDmzNf8784xWKT+LvAgBDTW9oKhZTD8s5xi
XiemAvXJnKznFBBxZcZfpThH7VI6xTkxe/NvWm/15EO70ESHM8BCE0rTaBUjVoks
faaO9cF6cb7deCuyZ+KQhbxW505U38E3q8996tGBLDa5EzZDbakMxU2yRT4zkegi
se3mp5qgJlrv03Eo+qlfelJHQ41FSgw6CFA192FVa/kQuYnbvANownj53aV6EyTE
IQ2KrXZQV6kccU6lDitgdufqw3EA3IAOVv9t4HFLX7u58s1CdK3jvftoO7XJeuC+
hP0XdY21cqJumH5fE1NhwOrYDMgRsXiiay0zUq74EG3yKWx04vWUSA2e1ZYLgzTV
ulEByJPNnks8XpVAgYssRaxcOLgBmLfVJqYGqPNk9dxOrr+4X7X25MVsiOkVqfX2
GRtYI1QNjCg/mqjUZyosMFBbIS33ZRh2bFDsBx/lkrQim3gIiIk3xphHaDF9p/RH
InWBLZvFl4GzoX9TCIpkM1GTCV/ptrxn9/yL24m/XWvkyzvkVoNhnc3m5O+RwHZ6
KyV0N0wBxmwquIHd3d7xxh8oSg1smvHdZTagdMQI7IhH9nq9KittHoPkbihfuUJi
lk2TklnDUhaRdPQRssW4WWwo9Hhd/bISEqBiFYr292V4ns+0TjG2TIc2CQMGNIuQ
N7JPO08xlWF1Fs1V+NH5JLZX7gRzV27B4fuz/RMw2zRfvaXblUZ/MH966OY/p1C3
BWv3/7Cz/KigK5KJLyB4H2aYTo7LLtCeRCXkOsl3vnobOK+Up4jvCIu49biK8Ga7
RGjtqM0J/+r62/bQ0QISRsrmvy9i51A2Q9kcSd471NyjgaypB9QVA47oenXEQRQ+
2WmC/EShe3IHnlrywnWVTObuU5buv+jbL/EtCJaktd4Yeraasvs6/qqZqeVaDqwt
TF6HXXwCHhsKENC2uNQNkhBYnq8/D16T+CUHxn/FatkUu/Ux/Z5eF+azlilr7fm+
rtCnuuTzyPRp+s3HhzyBibrw9BxolaTwyvHZ3O/nDe6touVsynxb60NyDRaYAU/+
RGhWBYDkblBdkmL6CUOPnCf3UZpffzYs0EiNH5YdSgfhfm47q4Scrgj2jpAZ/tfS
yn7tHU44ZnqVbPJsSyjeXhGEz2biG3H9cxsTSyZf8g7CAnu0EBb1cd+JQmyOreFH
zgLTfDXKnw4Urss8T46haOJ+5nRvlLDt0BwPBsO3BbvEs0AogVpkjfdCQiJbE2ob
9YRpGZ3yTm14eDndgt648/0VHQdTzUpjQA6hu4BhAbIZHR9tWMat/ZK/fdjuOJa/
AYOc0Dc6rzJnJLzNEeLDrVkhbT0PZO0igpDhtyi6VkKCiH8mQyR1gVyTgoqwuyXQ
KTWwE6cPOP1xuvXzUXMmjzqXwqgtWr1U7Q8of++DlRmJ6O20mr5RWKQ1hTVxa9AN
tbhd8G03pAbtlZ4sRCzoK8r950fZr9Lvw7dNqKmJPrTxL4rePRXuTG98K9W13fL9
sZ7RCIV0M8QxfI8n6v8WZE70yfPXseCSztLYydsFL30O101pVatUDYODiUZcGMx2
qgQ/cZEvJJjmc/J2C5yojShne4VhvFYEJZ2LR2twUfPDVGq1Mz2UDF38a0SNzxPW
zGiF/T1Oe8hT9JnFoPd4vJu1TL6Wno1OsA6g4zhYzQ2Xc9GNK+UwRjUaepI2lKJv
3zWUaFdWp2jXPwa441vrarJR1hVWRiVvtZiRjItyMw0O0k36G6iUsMlZXKUz2ZpM
uXDMn7TMKHAOJnlgaO79tnrCEIfj+R54MLuGOv0d3jOZ3P7Et7eKHgfOx5MDHMFH
hiCU/nbd5VsZdFo/36FNIyR5s7kOzgABauKenKc21OYZtBfP2yNzeDmkFWyMZ5sD
zQ0oVI7alSC7yg7PYi/FpDzjMGugf8HKvyjBwgwzm2Rb6IIZWELwJg+IM1XLnx63
Xt7nAyQVzdMX/bXG44bhO4ImlwZhKQY6eeHc4CVcrGUmH0O5X5vm0HzFOxjiBNB+
gjNCUlNFzX1WwRA8VGmhcPKFlAQTy53l/yErHotj5A69TjRDQMcLVnALkHFv8tSI
p3/G2yCfsTCVbTbJt08vyDpUpmJqgMKt89FqTwpWvwcKG4jjXau4xUd08rkrFhpp
u5yM7vqTTKcXcjOsrurlXzWoTbomDy/Ka/kCJjN2DAmBdynjSAPbJ4o89qyMwnH0
J02x0a/YciT6mThbhtT3vRjTEP+LKumAV0YA/QPKhq50sUY4T7ZePsKS8RfZdDHi
vi9G7LEy+rxY1+A+8H6QAzhclKVxI6wZp6+XMurVOlTVdX0NjPaSJghctjNNt24v
PJRVNf96r9hNoENgmMEV1JjYN4uYcf1fNiBwHj6yYTKwEH2uf8f3IPVYXftLM5cY
WiKP2NKaNr+fl91Fzzn/a5EZ868wBkyGA8bIcbLiWa5oGQOkHMhblePBPxsTlxWU
IgYmg6bF6uwVT1vinNyRFARwZeuZKBjszvtFoip0U/QQBu86jSP+qTxD8tR3Yxzx
/3UDYEL2+P3SAaZ3hD6YRYwWy55l1J292EpFjaIQ30uYJqQnlHO/0/FG08aB4Rh/
c82skOURbOauKH0WLJqp4Xe19hB+ae+HKc9BsnTGj10+xKjoB0XABBAwnBlm7pCC
IYNH4amO/ZQsz6urAcGBK6pq5urccZZicm1HWjmI0E/g7NwzFcSio4SDVNsJZTY5
6O158sGw0UiL+WBUu4vcdP6nNiw5BdDNjX/esQLl9cSk74frZkKeL2B0SvxyjqQ/
L7KGbjh5YKNJd9xDy+2BD4TYXQWicGQk42o5ycsB6mJze5s0PjxcXnMEgrO25I3t
H+nYTtHxs2Kz3nYnFdDw9CklsAJusWORYWIGtTafTY9CfOvgP8Siw4BdsLkEXWQz
+dECgdUvNeqjUEjok0Uwv6/vkgoNp26A0iGGeiowFQfHIEoK8PejL4yVlK+trlcO
dN0b/DR2IqFAgfi7K7w5iRpDzaQFc8y7emc9A8RHzJ1cJCVXWQIBVj9yWYhCYmGM
wQyVIX+YvkUFhqG078hw9nmtzh+g2mcL+A1hpcDLxarFPYcJCa/so15930hBzOC4
PrDN5vKhAFGMaU2lfUhtIm9GEWq0kfeAxumJ2Ot5fYcDYBadMeCRurP+qaxnzsbb
DgeSshQbPrAvrEgRr9Tm5YWthDQ7X7M1T+fc/44E06YyfckvugMHUj7l+TZvLD2P
cBvIBh+zr/gTEb65Bp4dTOV5KSvkq74lPTdsJFA9LpTKQRmGPoroTtMyiC68HbLq
1RX7DKUaZKkMWqZh+PtzYx09x55egJDH2hk++SjyEHqWN+yoQjX20tAchzgq+QSq
4y6kpBG3WCId3B7UM0IxCEtcxxEWO4/P0/zdIiaaUwM18ZBJTpBepr4AJNI/iWNh
UuvSDs/4ll3xH9i+n7xpsNdZOb6OoefNYFytz6Ds0hjpoSiacV7MB6Tr+wVuW3dL
bTVjNGLizMWO3ra5m+ZLexecu633XaaTOityRUcbaflFnLCUlWEuPwWXWT5KuaBk
vbW7hBBqmIrgyYfGQ9qkPIoKNmBeHEiK1Pw9pqbaeITjQwMqVD8M9o+YE+ohFItL
0aMnP0Q5iu+QgThLvD5fV9+0M3cvMl9Mo1Ekfik+N8Fpo7EfclATMIieEApqGpg+
NmpyjKkxN3mDIaxQhYS33eu9+w6BEvz5czQ1iFheioMgHNFErqsWX06S//Re7BIV
8MuvBiW+54qkZjGdP6al5lj+F2Zpb1GFBGSCJ3IjFPyw8VEk6ay1dV5T0I/pblgF
dtWFEYbE1+r52xepijmxE2zoC77KO5GqbB2QSFManED8Y+P0VMU7ZXuVCAS1+68Y
86DMe0Yo2SZ3tWNuWMo/NjtwHcWPXKgjZMDN1suU/VRxt2sQjouTSdwjQ4/GuC8e
o5O4ooLIXGy9216mACgq45rurjpPGRKoLjjMWDgNnjB/d3xODyEJuMkpF7rKz9+I
Wn5a8hYJXe6RA1f60hLTE5kGN+ab6u9ovMkaVCL4G/ErFNuZQ/Sv/Vo7qot7Nz2j
9eVN+EKlkUGQugcDUHq9/CBYrnp/Fd9xhihy5rJ4QFN2qlk4iOB0XgnB3RTNJ5oh
YE9ZOpwBNWe109ZOup2nWRiFxNSPsWAnjMF6TCBxJKogILu5IE49avQWK5GD/Uxo
MJ1RUWGvW9UJlXyPPfpowSYOaDBlsoxBMM7Vy6jDzG1I35/U9eQp2YriozA9OwK9
Bo7qMS9fgmbUE3F5HOg0BDYoS6UNrIVKOJ6au4Rpk79q7B7rQPtIpce1Smv7GHHY
REDk2yIpkJ2AtySCPMQXjooD7V+BzD+MiKhakHG3cfVqo/6L+NxW8KgiRiB1QGY9
gqevmWcZKQA9jM1qvbdVf1TYHBoi0c5pqIQcrVbWZSsuUGwKDo/sUiJSdDV/EgTC
MKVz31XUBiL3ERKsDLWenNFcnD08N9B6R9s+/N+MH8ZNjwqrglEwuzYjRj7/9J7c
9kwaNoUbkiPK9mdUBg5VqgB3WRV2FjLlxnx5YIecTppNeyfBuO+leTVl4nz0LjY6
Y50pvnpliBi6ZDrIDKiO9PbnZLqoS9ORDJZSaxl8lby7yDlL48UnzIv+iavPUmBi
p7T+VsGkMNH70oMWv9Gt5dO6SDD+j89xGJJooWKKmzo1KXlf0BN+3tLFFXjWxOry
vWajNorAoptHxldqmeYsqXWLUoiHPGb0ZyepNlRXjm58giI+zrfJAG59/cSLgpxD
P6fI9NJo3Wpka4bIukDP1w0o/vhRJTULgz4yLHPMBE5KNqRJ9wzRHJhsWa2XEVjP
6bxFTrLk1HcoFHTEO4vMFPIrHLid5XE94/yKO8r+VD20ctnEczGMjdwu21cu60xP
eFlhj3hW/X/RRKYdQCkY8ORWZcPH00hlSkDWFERUIlDj8ZuvUXWuCyF+7MczcBP/
UcofHck3BXnY2G6/2aGrzaoIfOwZs7WCy/AGvMLQei4OkiM0wjaqPc1zUI52ez4Z
bBep0ocBZx1uwD9iQ/SDY2ahEq6kG3qcxwUCe0miQ+1syi59APZ5Pf1eMe95rUVF
FNEyWUZfFqMgQJ5kFDuIw2tX8y8B8zYnxLJbDtUdHCnKDaWpefMpGkplLlmTa5z0
TYNn6TSiAoEzU9jbbtq9mddtZA/iuDHP5+nGHTKsqkXyIdA/LWWttY0d+pp0eiO3
NuM/OMhtaZiRp9azPcNGJWTT1BXiIOa01pl1YErzvwejHi3NT58I+wwDTxJ2kQ+T
aLKshuDDJ64Vskw1WRs2eVyi86zcoJ8cYc/YUUpJLKJfrzG1t7Fv1RT/p77g4CCR
/jbE7M41SrGv9NRusPiaeBr6VcQdsbWFl/7q7PozpxhOW47atn/SYKdRtj65TlrO
/HrTbZwmq0QlPorTciOcmi28UEagfPJFchX9Nsp1xZUnLM1+b8KW7Q2Yf/nQuEzC
Mfk0064BLAxF4jR/4jEqwf2pT6fpCQRUau6wW0EizUs1m47mwKVovDir4UX/EZ1e
uLN+nRtRxi+KRSq1kkUtwT9U6HFzsnMTp7c5trvkD4kQJBX9xQojCLMCi9WTLiY3
ppG9XrdGoZBKP63rZZQQavQUElr3fuU1C9bW2lkc4XN7x7YHIUjsB6arPLOOHikq
oM+Xk/HNXiiLdwPrzbmr0Hs565tKnCBVdx/DzXfIQvRKxU0bhBFmSdCZufqavPu5
fgH6udOQB+t/uftBgGyCP4eHBDJDTQkSMj982EtZqdOEXP1M7ovhMIbRTmEbxNm9
mm/w9Q3tIoLdAOzGco6ajKwOAQ7/+wJg83V/LGLxCzbP0ddhY0QBZ/eu4PpN/WXp
7XwwdoGtYeRy+1V6mN2r37iuspggjXTVD7qEpz6qYjb5oL5SF6yCJFxSG/krnCfX
87RbusDZ2Lm+D36LKujrLhkJHmpoGtCsWCUcFYGGI1lzfo7chZHggOZK7aiguBFm
iIM+HoG/vANY+p0bqwRa8uOy+2ASe2CBGscBXVSyIqQqqcH5QE2ivECuoRphWcu3
nmQ5shb4cvcj7mARCTn7OCwgu/j7af65rm8lbLrhFYPz/J0qGykvMZ47bqBm0dOX
QElL+d5XzPVvx4PGcvO0paPM3vMNMLMgaMvcNlDf2YS086W2nnpQVEJIZ8ZowORa
oAkYQMNQ+xizEvB/LCcpcNIo/WvPThx4ybsrgrZswRlbk0eAQukHcy3j+Af0LAtH
A+gujdHQf41ayaToPE32wVJJmRjAc02HjLHxex8M+9R0W8Qk49lVAabKZj1YYZpZ
BmpWgxoadmCyOTQ48SlW+gYEsIkD2bkBXse91zDe6SMCEYPk1jBA2RpjzFx9JL7/
BfKvkl+TmcAAp7JWKLx3EMX4nGzy0hogjA/duS+K7U1HB6Sz2818NEdNu/hFqmxc
Y2kXDKSYPkZ58cJYE7ZiaFDGfl8rCFWqE2xRcs3WOA0OoBQWCt197KVqbhdtEvEC
LKOY00WGMkwRlOGuuGh4Hi5cwyPLXEUjz21UkeIAzpKd9q6LJ7kdKUPp9waAXhnS
gMhiGcqC7h0XDlyz1WfRwd2IXjaqzkYtwJLZNUwscwPVgjqk1eIZTBspkHlJ/zaW
wNz2AES+qk4fRM6+DlWxkP0WXbU3c74BbFD4t1ATyJ+EAaxKOQiWrzQToC60Pirf
yc7IQANw/aBpAviilAw9+YEIfkpEjPxa/tURQWCz2NhFRZAaBYHdLLfKFJT90Jve
VbvUB8E4kh4WMtOBp5H/4jPs+G+Q3uMyyHntKyiE9QJoGVZAy66FhfLBywFFg4ek
c1XWoASJT6yezBUmS53TIOckPY3v4B/prEqNQucRDa7027Ie/lMeNdfJEj+0dh3V
sB24Iqw3/neraFTemgPl+m88yFnB8aC4jeu4JBoFXvfEWQX7Y8eJgm6OaTEMIc3Y
lYxWPYVvKpda6O1oZYQf5Eh19W1jaC11exSdIh+SVf+rJbU3rbbFZv1HSt07ONIH
uT404CDOqYdJIVtTPm8kQvbV31uR/zqA82czP3m+7m1SQnIWJMpV4nric4MEvdOG
93Ml8nEgmBG8bChHWikMweAJpUfBiTQaSSZRsTC/u8E+tSVD8hXntgs7dA09shFp
KwRdXvrU/4NZ789F3CGXVxdy5H1K72HS0Sz0Y+b1g5ttn5Tjfv9QFYYRtEKwtksa
Ud9IRAI0/UEtxBqPAz9Qxk8c3puJeFk5eNJtk172ZTfTRuJmix6VvNiuNHE6R8sb
DwqsNG9qN8ssimjFQ+UCeMaxJnbRfH6cmIo7rsbYGHnfyr60StXkAyhQm6VIV4j0
A4054mMbQ3S7OHf5WrOpPyGTNl0JlvNOAqFSktSQtu8hnQbSQrocLH1TcBoneym2
YSRDGKUOz0CLhj7tEOQ28kiZng7Vj2E96eU8pVxmcXkEbUQznjRzlB5hUqtKE8K9
yoGQNeszzlwoC+Ew0hp7KUf+Gxp2ZGy7ookO0/37SahoAY/wVwExWBlKSz6NcBQ+
o9S4SmbMKXD3f5fXXuLXmzFFTs3s5iowQun05uwdbK2M4FbMKaYfoWE/svGAlF+V
MRkEHuSEE3zGxTWOLTC+MB+uYNiSzyn6Q1AOm0ZtTlSNXz7/S2I1RoBQQFn4zD+P
yokEbu4mL/bewdqFRh9gvgXjR8xfpzEyoR6Z/16gfwjULiSTWeD9s2XMm0h2FRKj
34inlnXIUIahUAFJ8JJWeUM2c3cDy6SdIEPeNi+evduuYGnDF8EN28WyqSon9q5i
sP1xM/r9S9oF0eV+/etCY7qim+SUTQ60MDB7Xe/x62aVBB86vTk2QTSSCokrLNiC
5y7F31XrlxJeF9skvaCGMdJxKXt9Ic0rcCE2j23F9egbqn2y2cUIIXaLwdWUxXx0
GtcudJ3ij2zS/EdvL9WhR1jAP/8Q1/kQQk6GE33Kvw81HW8DLBzN+wR4rpdOSaQQ
6O0aol/i13gGD4VhNQbtZneAFWDNbXFPOB5Cs9NBKFQ6MG/hHTs6UvTD2i9ctFVi
zgDsXgJOdsQuZHqISTgNAZyjgvzEQSt0i8j/3hCqOJqK7sTCVOJt91TY1XMdJSHt
+QQLwjR/FYXkDfoo4QWsBo10vO+HriV5H1ri0z7jdws+B+2p6Oc7vP+yG42IZUhI
pI+bkawU5Xc1NxKGVcjT0PuNTSmdVxjNR4i4MKP7rfXiFng1qo26GYhXbxNU11J0
t7HMZ5X9/2xtHgDIqc/y8Y8Bbo5U5mDFUtCH2k2bXlLYIh6M2M6UM2Nzz/npcQby
b2icUeKCFeisTm1PMCFIdaU0zhpXKy5kERblhFqxYSJ1tHLmYhOaZbJoGwk++Fe0
6fXS8sqXZljw3aUKolUmA+cvsKscBfeZphgH2h5vvXDHYzuukec6rPynkrP0QZu7
neeVMtuG34N9o/e66aOQTIsRHK37/kWIiDCkxWHnZMv1EhA63m/IwlfDqJQOEl77
HMpAjm3JtOU4nXiUFlplS6fCicYCneE6o0/tN//Ao6xhEH3LDu91VJiISqZzsI4U
q9A5K/5SRK8bqQi0JlW84+qDeewM3Oca/SUVaFgdS3CoKGbd86Vziyj3FUXwhbVJ
rfdiEiFpEvUL3c8xgvNqoOHJvqUBsghULz0FF0DApqooAIDrIHxNkOH0NXmM+9jk
t+1yRcKLzhj+HHLj91K1g5HzFQ6ackZbCVaS2rsEX6+xireYsfgGP2lR7s4SC8LE
aJtKNLc8nXJPeSnhrBjqIgVc9In5oLLRnjRD5U/g6IZjprZf5t7p8lVTFYIMAgPA
jh2i9P75HsU/5uoYfND3cteIjwnXBYw3lzsXE+UXkggVPd75F09UCsDBc0wE8Mw8
HEus+U/i0BjIBaU5NAeSgtli5R8UCzZU5M9WC9DOl95K06QTNivthcVG5MdkoJZx
7gEA1u0cS7MDHHrCjXj7NzAQL0F6GdDt6IHU6VksE8TM58gMG2PHl3jndM/oM5EK
JN6WrRSMdQ4+ijAMmIUApty4iB1N+M0BaOa12TUmi2ZjrWR/rBJNKU2g6lxLzwL0
PjqMwULKiPjvQx2w7DZWUaxQnB/DjqS5aBvJHjHeC3k9PKI3SBCuhoahsgX5mPzI
1cP13t6mwr0gnY4SfY8GEZCg/5+beXtrof7SrSXVQcBT8t9y9YXla41KPEwQZfF2
KauVwPihhKHVdiuVHtMTdZ/+NhJw0Gj2aTM4Ui2+OcQB/aLHUqskNq2x+m93mLBl
yMr8GYtPoabYIVaZpti+kq16+hNLsSh/XsxBJN1KBm4NhuZwWinFxP7vxDG3uwgv
zPXYidMOehjJ2l10JxCSDH7saxpe6Jj3h+8N9FVeKZ+6UnroMq+B5D2Iezfu64v/
aDI+742kFIJnceumHN0PeGjmrIAsJZUGYSl1rxwHKmnBKOz0uCRARgeuOlQpdASr
VOlgB5fOBtFtmYpUABAyIvA8DjM/lX//YRRtj7dMnYdHojKLO1qU/bkt8k5RO5FN
0WrvWbEW0l+SoZ28FpieVK4ScQeGyVOxMEnGH/upsUtm+pnzp4Bme7/XV2+snHko
Kdk6yCiDeiPXEJj+yOM2GhUhrhqoEbsIezFY0YYX+qRxDfBFu1zBJ07RXI82PFad
C4HukAE0aqqBEcwQDgXc6lZz+5FlID/mljv/Z3ooUMR7l15u6pbnn5JUFDtLnFtq
fzJPKE2iBzwQA+ABMNmVio5UrLEHdPbYOT4dcRSdMWVTSkg+NRK51SYSMXaq0AwB
8m4GFmgfokUXLo/BFD+ZfakjHWTwvHg2dpNrpBz+m0J8JQ93QoueggLsOqozz+Uc
SENtcM1zd04GtAlAFE2xfsjIt3I0FlajapmeTumIqbP4C6sIiWZvqY3hGKYqpBV4
pI2kvN+yYAgluYrXVH3giICa3TA/D4D/qUP7/1WVd0WJ5QwXaTGq0hBWs826WTnI
3PAOwUb+RLMcROSCmJ3V4B+1RAHWsEimYVTX3J0NnVAOzeAJhYDaRI9sPdh4rhx3
v+x+t+7Z+GkFacetwGxDVpzkBOUNT0jslw1H+krtoLq4VaHojxnAEyMTk+5ANRw4
CMdOAyKtxpEV2NVrcEM4WKrLHfhda0LVSamsCrmzqM/wMtp16kTaDC4FQu08dZ0d
8asO8LwZcBfXZN5gAggDS8RyR4bPObLfhYOoCG4Q8Hv5+87YoRCZdBS95zdvwpvl
tn1OuuKy8Nd8ybPk4lT/CcqIZCjqSruJY+GAUcLAw8gWdeai3JaiEFAyslTRa55j
yHkgo0FWhx5zP9qAUo66bIUdM/IicsHmf6m0SX4avCGm7laDcvpOMWpIRtKO4UzP
UsFF/wY3HjtKF9SPKVsOjEyS0mhJJVgFxqzU2rCY/Mp6syO+ydyOTe3DTEf3B2RW
QgPY3dKNKeBd98GefSCuNOAigbqLiCOv3EkRsOa9GR5pA7NIst5MIjYdDEgfwwbr
JoBz9dH7NVLYXh8B2quIQy7XOLI7qXqtWl/F60pTZZwcQPFoPPegGX/BCoe0NIfE
59TKLth1dTVBDKwEjyn/auzlkwjaGoZu3+9T1e5zUPS9KlViwYe3zQCceDIFPja+
k4NI27p80NfJJpOVJWsCXY0B/FnDLOSy3+4A+q/hM0sU7Me67VnVZPJWEWJt4S8t
i+q2Dp2PuRKRaU7qr/luFKZdz0wsRqaAZlqwU4Y3OhoghNv2lZtXOUHXanztcyxO
ZkLWstGKF4otNSetgaOKnDybdi/5pTQvpoqWj+naZ6eNTacqSLvnev4sulCnWaS1
yrdHTj1bRe+xis9e2kXMIXFTQXozIfpc2WJdAyCpnFwyyQoB8zh3PCbPwuzo6owC
hkN404Ul8ItSFwTLeV55jp87KtFhDeMxtuZFlqNPbzasP/OqGK4yQ1DRkG8B1mip
9VzBjEIg/NGzi0hqq4Mxyzjej7A0xXKcNMk2am5eWZen3U00H80sYWztRQ1dQYRp
Qn6tUWYII3atTiEUVtS7NAxx1KEYEW/UQC+tRrtgGx3uT08iA53y9busZIpKjQDf
JFyazAI++wCJjUJU3k3SevVHHR78fr7JxTY4FEODotyGYlYzRrzdW75E1r4f/F1U
UIwOZLV0Uw4JmQSwM/b1TBX9iZnCEUTXJHGsWFC1Rb6npzA35OP6KFS6wQh8INpH
kSNeSH8nFRnMJN1mq93OyQkCYdvnYXXKlG/wODdVNuUtAxs6OEoy+qwXGCV0no4H
+NwpTfk8+WTVgLSjMWIeNOInJN5b1BxakqYMjIc/OQe0bPxeKZFZ5hu4sGBulOkh
eUNVlOgnh5/4uTX2EKK/78s5kg2QDXuVAh7QZMWxVbV2qlyNx4OTpOsvx9M2/PRs
GBOweflcFZqahIHrLQneY9n9r+y4KixsXd2H0hHe57RbNRFmSp6jWm0Ga4BSTjt5
fbpEJrDq29IU3EAG88xHXHTBdZmZDTYknLpQ8hnIHcQkXSOXx9B/aA97TJC3SgHt
IBRKfxM0msMl/PaURqmZgrrdDr+mP+1QFOh22g5xeuPcNDc+DzJ08Pdchazais9v
HoyjZvnSXu7e2fELRgInG4JP480F7H64gMfduNDVroegNEmPAX7BKsfueca4rnrU
2t+iPrFMh2UQnzQQ2UErhIOBqSP+C6nHac0wNhPXb20sru2eCahLXLXSy6q9L+vZ
Iml63zYO0NV00lQ84CgCCXux5opAlahXb3uGZJauRraBfsKdp/pb8tiPgTfUfLwu
79/IZkbr6cGpvN6ZhsxD2S/CYDR8F+qWZl+x/dRWkf+x3OlDOHDyk30XjbXFleYq
/t3f8zo5CC4bi9kdA/xCYGH24W7rF/R//Wx1KMAvbVkW/F/EZEMrPGrEosQNL8cW
9tubNEAC3pDc5VZ75CIISFQGSgzU61Bee4k0EfTrR8I9fvDry19W89B9QFpMSgcU
ie+RaM0Jc5jD8hCHloiK/OkKZALItSM1gJ62s+VuP9Zjb5DqOwpoFnpXy2a+EF7G
6ra/eHJ6IJ+DBJQCgRsFmMoXpeNfn9V0A+fla4lMetCNO18IpJy5hh1tAzOLedAh
KrHql68yrnZCtyR8muLLlc7N9vow35xBWq1F0s2Ebb2w8PbLKKoRHLoPxaiFx1tz
OBjzap9rSsTdziNe/ihXPGO2xEESZ2ugf3cP4SRMCwn7LjG59d3PyJg69imOyAYz
IzrEb6ixMe7DgEhSGXDZWBs8hF6v+IjssXgZQ9KmNJZ7fpqZvmWqCw+HwQjbgcKG
l0iU+YO+3245kV3ewzGsq5Pp472UoYeFjHwnDPLPGo7RZG7swDha7NdZRFrLypY+
0eWbIZHSElqMoOgrvje6v0O6gLrguiEyNyuEhEhz9ADIlAMBD1P238D4WI7II+W5
p+YA4OgrrCXhl+b+NDQZiWzip1RFa7C5sbJaVXpnySESENBrnEkoCrxQzjGbslz4
wRfAPnKaWyz77Jr+DwfzItFOBUiKTAwky9mpg/6OTMGOkvF5hwd8MFaTobGKYJv0
DF652kWhtzv2UW/zPvWwY+oz2ojUgPmYr/V3wAN/L4lYmuZOi9f99ARN4gvAig3p
qR35l58f/3MgJurnvwmPgBk/Sm/XAhp3QPggb6SenwwCEsF88W54lzkX1zHLZSLY
xizobp2k2s/RQ0M+CYZJsVl1krIVJR7cJoXYshwY6Oljm7s7/NcQMJjCr/72sXsJ
LbWtyKV2btivsdoObaFeICD0h7ZNvxaezN1mkqhK5AiBz1dpq7GT/ap9lLsxjJKW
djaPaAYLveYTXuuPLPpCISJyU/R4vpjme0Z9S1wRKxjZEIkE+BC7DHY7mX7LLgVK
FVwiQ21kV1w1DXkr2HVG/Z2IYxdtFNMrsPpC6KvpyXsSK5VVN8Utwi3flDb7Al4E
EWrWS8gvX4g93Fyn/W9eAY2sQTVEMssGItUrmEnXCFhdn+CF2S7FHvkO94n1qM5a
4nE4OZp1FYqBZcuhxF9bKmRE93BltyU7BmJwqE69Ad8+N9SdgARXiBZHqZ5iU8NL
hSobx94pz6SMeR+RTV72ShCoNAes757bAd06fIAi8OFWFqoDacyw9j+mH6eUaSzH
PpfaeCgdin8CmX3Xa6a84P4ynnwyXh5wh2kKNqKwB8sWf8o+DD7EBpasRs3ZJm1T
b0SvAWyZWs4LEbntDbJgVBf6Y1HZnpoCVgIEsfmvfIy5762I5cmA50NUB9P6f3uo
1oMqroCadsetSBAG0YiycAOetvo0Zjr+H5V7cPUgQUJjQbPfVEI0O1eoAG35CpLo
eG9CDf5a+KTNzOiQytT2vGhG+ag7Dej9nUYWl7zVJrnq/1PHKn37m1anV+7vsL+C
yq7Ob6o2D5BDrVTVhYJDRa+/J4W2sUaN6pFXEvYAEnIx+pOSow6u0sHrxacgNb1K
+6K0HQIuzlE74xPKMVposfVIk5c8q3p0CTLhePnHq+M4EuHLyNGgVjMt8wYbvxhi
5OYhxvJIVYMxa7enEVe2DRiVU6YjRDb6tLDPHmSEwnyAEmfGnBNFHkUcjBoQCrVS
ceUeH9eETKtbAPnseCrT0iMKmFcghkwq41LdsGg9TGzR7TgBcnmHotDbeVR1oiyQ
XrFtLOQhbaVtd/qEd8K4Yn8mjpCeb09WcWOqJAgd+PEUB1F5CSCkYL5zkI2VkNKG
BFqAC78x9/WeoFBRkVwZL6tR7e2rlVIElPkfFWG+/RchF9kOelHXlhQcNqE6EOet
ldJrjdRaNtLe54TlVrNmGXT4OQ0BmQxilWhEuwQJwYoo2Pjx8LdbVi5d6hieks+F
6iQGZ9lzxxe7OiwT4s3523o6ANgg4KmGj7EcBjwGETCtB+rc5v4Uq9OEukHNfAIf
1BqkO3S+o6sqCP4qUT6FR1Q6JZp51QypYdX8jOpptHgl4MgRJwITfnm0Vb9RhD6t
3fFdLvMWoG6ghQtgy4W7FkijN73NtGRIn/5RCI3826N0cofIrfHeWh4hF4ufgaoU
7FwwdMqDrl6TxS0wI3iaWN0KEt4xLPo7vJIyGRO+pRi7VllfGu336zJ7JXE/rVGl
GZNbdpXiTHpggYaG+dBnJ20qADQm0yggUn6mSg0PqppwGBLlApRjy/4YYWK223rr
kgkebABFgYX8mHwpmEq21yyazRK/rRX06/3JwV1QTn7nBZ6bBVKi9fZOd3k/Zmko
7m5s/cGjGdyhvtVLNUmVlRdnViQa9WLnVxW5jZAXEDdXwtTna+ibElNuvwTmj1QB
O2G1POHC8+uZx0/ZzfFpW2SUsY1ZsPGVOF6xi/z3ZXPYL3WLgHJWWrCPPxbq+MG/
A0pTJR/RU2BTnGX6ui6w6RwmTwWwKa7DWIrGa24T83NeZ/yFo85JAPLcY78mlw3B
245xfhyujUMln1AnEUIa+AocoK/iCJOVbk+F+6BYfRzkdql6XDWxWGjPnvimXyer
vdAgPP6x6t1Aq0okaycutz15Z7AM5IKonbpfkQnWcKnzIiNF8VzHUozPSeUtWqqD
8X0xB/gTmb/HqPh+bt/vQ+KuHYX6AOagpJx+JEX4d5owyGBivWu11Ghj4s80gIWX
6hYynqgr6QCUIzgFExfDlTQrvpBbEKA9zoBK5a9vN36+1d0FxK1JreF/TobuNLk4
2DUsv2co3GMOTl2H9bcx1f9jGzqSmVDMSoVs12EHNCviB0+yjyLZ78K1UhnweHhq
K8O4jT5PIvSP59gqdwm6gS8FYobIVTepaOYA7/m+cAc7RMTX5+wrIfSwraSDfCcR
evsOMe7n5T7GkGmwNODmZwPhj6AycxL9k+rMvjfubYuX2Tp85UyrAFTUzpa9PmVO
gGS1IKFP/Bu+pf9wFEJQ1gcj7qolCZTkkeBi1EARFS+Www2b/627MHGIvJZM6WgB
xLtqPsRrKjfna+vMVjN/ttHUek3hb4A6IYLIwxMwp5x1LBbm796G3BhyyliuTF7M
2KIeZWNJtNcOBjWvwhej/McxpTRJ5RnN31IbErtL9e94NHjKr+f7LKkm+/V9ad8Z
H8gUqv0B2IHcvBXBk5JUGN9lAMBA17c5FSo5tOs0YLTjldM4wzloPRruq6o1VeFz
G4p3FOWbTGllKfHkEaCz1pUOgwfheFMRso9Nj0LTqMuM/Y3aXnzemkm/xsmDrjS7
xYHv3EarRo5s7ELARho1pwRx5gTwgqgK07IgHaaoY7KU4BAu4U9pmozBhzoNkDCO
/cBgKOeCKhRbndp9g4jI1BvRUWCKuXldRP898pS1K67VYWTtRFDCpZx0BynLPGtg
QPgUusTsqin07M/PZeDFDn0/aZX5xABtJV7X7YZO102faedX/Do2iUOng5NJNkPm
Td9VxjckGhTVR5LPP3L30T/M4KbssrNVDYNNhbhNCz+OnYu6kz0SICfHAK9HjwMZ
vt0xjmaAR536v+OjOgD2HSdJGqiUo4cM19RDKcgRArkDdwEdUHnroRVug6srAbNh
6mv51fmfm70VJebK7rHJRB/YkoeXklucw+FEy2DE/RnPy0FhuAMRUMpWeSDsunQ2
nL0MLw/R3XmBFGuKg8izzb0KYJkdP4Ms1tBwXDbcSyGuuE8Mys/04xbm90E1T6E8
QHY4NlIzti6TZ9qhUgYa3fIere/RcOJuNuVZJ/ksA5I2hSNj0voi9LArunhLpYo+
xZmfiRRUovOH6IjP+L9F94qVeetxxApslNeRyHw+7a3+F5E6yIwTHZkZugps9kRy
i4iR9gwqd2LlOD4OiibH12j+/Tzd4G+vl25mBgpNAR3zm5YUp9WBTmhDrlw9ncAP
UGI9PScb1VYN4Klw4FR/MMTARQrVrWmR3x+AMFnCSpZGhY478Gn/Y6a2/xb9ovLs
2olHWs8wvoaGqQ6D82K+pDNvBvQzHoimUobVpCpHTtu473048o3qFmOW6GW9o0VE
2EvvIT849/gMZyvNwPMwpHNEp/fX9LQijN+fxajmj4Y4MPeEPHfGJzCPpBIvkrYB
E/hc1zzaiZNEPH7bGbjpsm0b4XDSqVMJ0ERYnn98ZHiqlZlkCUkMcjYEXzvsrk6m
e7idXHP5L6wzKS9uEP6tDeq7UKTnHlqNDGhTYO7KSrPnAPFGENc7bD9qhRrHGdJM
OZ1QcrJumoppV6ZeBu3yTHEJRyP30nNJVUYolyEH5a4a7aflWbApgjPuqriT5Mu/
3B2B4g9oOA8MJH4ip0IMGuABeyaAO5a9tsaYO7mgA4q26B3zYiYCrywNyXjJWPZ+
x6Fz9A/KclwphV0DI/dHjh5FNVx2gkz4WgfamC+906NvDWhynuNnjBN4wBjKxuOb
YoDIziXgd1UTpQoZt50UD8PWgXrpVRq7S0TX4RlRRIBdNmSe9Iaw4PX3SK488T1m
AAF4NwpSRmxPFilF04KZAuoDACm8RlFZpnkeucFIM4EtNqvcd873eRLxlAHQ0OGf
Qerd4it9WDA0PphNgM51x7beSVj2/umOm7EFYm4a60KpzsCgbjKYrxSWOLYHDSEO
xBB64i0g4pIFadELjSLAitfvXlo5ym0VGcMwwmwWuMrfEwKN3rTn4uTDkA94x+Ev
sCMQUmy7TbSdCvWwjMD3grKjwcO5R3B2NyBAEALtcY4QdFZFik0ndgnWexag8gW9
PNVaRQ99yS2PeLwAeWroULC16eFVp5rjzjN5+PWk9UonTmbOCqdVZpyb57KCnETx
7H3S5LX8cL7NWxHZOJ8yu8vezEH67l/3dE4WogM1yMdfyxNzonuy7Ac3N+rKTh7t
6cRz9UoWM/3MI98AMwkvbU4wM8gui+sW8Cp0sKItGaQmCuEovFy4hIepUnjDmIR1
gRf7eGGTe0l+reFR+Q9qZ5J6lYsdGzaggj2Oc952iQh5xNV178G4InZpc7tcadA8
yxTn8SE/T5zvvYxne9YNNWYd2FD4BAU1YPwAlEFUzKqw8tCHDsDQ/aulAIu3uY+F
vPzKTewZfk/je+7Pg4hMbJzHKmjzpRRbQaG3MHYecd2/Qk1ZOirEgQqvBKQ8gNrz
O3IMpBCFeuJMJGlrF2/3oJl2s8eXLJjGsiXw30ihdRirlmI2Mq3V38rhiVYPr0hL
YpACEyPEc8QbUdvX5nUw/FdGF2gljxQs9x1/6O5odtjU54jcyxkrkejtcc7RCGh+
38RtxCSDYCzvqC00OrtK0PDoGJQNZL3ViPwIwzkdPm+ZJPlqgmWmeRoVOt8RfCjN
PpjATFH4HP5YXpWN2yR44uokxMDy2xMCUaNvwc6roCmArftVM1G3wxYhRS9NJslU
3smMF+6+iuS2APo2KlVU3+hstUERR0mxw8o65MTzfvJdwRe+cw7xPJbzKDtJ+EgE
bO0eaj5weD9KB25YbCK4nRCY7QCF/jwNu6z4z1yh4HI8vNVC64508i6SuIWvAx9e
f96MGUpTzPvOJWm/Rac7Tap13lRtL6uBMmg33PEiDz1yuGEYjoZQ8cMGar2DrBk0
nokZSY0pEc85c5Bez5GtFSUqk8ivUOlpiUAD3WOwHUy9AlvDVyiHfRV17+GmcmOF
auu+5BgsGKbG7fIk9e3IW3GqO+lp+gjsdDDmaPVBw2G1BU5LQfdWemK/g8B9p2Kw
rnCFLBJXrUe/WFdHHEzehapMknUaYQqkV2bKyQVvOw2O3zM4pZGw/4WeOe6Wl9l7
H5Y7Cf1DilgxfFQ0vpzq5iFa/9aZCNEnFM6l5fMnlnTBHqzWMuX6o7CaFK9rCfOK
jNGm6kWpj98ndSyHIEdGFm0g91cUCEKW0yH4iDuiMN6W4VsszkAHnW7/Uj0y3DqL
UYW349z69gO9krqTovNEFtzY/iPfAwsZcMeXMjosfch0c+lRXzdPc4rBUeJ1R19C
NcOUmYOPc90N7bh8oQUyHkD1DK0j9t/F2fGA8RpTdrL+3JpB/7byUmKhRywxN2I/
3ukrfoQp45Va3rMz2Gu5vp6K75kYlB4gT6+/Me+pjRoCMdHUHzCzA/7z3w6hY+en
JTUBLL0JoUu1SRfCy6EDdbfrfXpkleLNw+oNSKlqKm1EhReOQHDv/deZoF3ae5Fy
SOA4fYwljDrOVw5Tu19P0egf15owdW82aDK4K5iwhH3uPn40sG1KfV++sMVFMm4j
ZEF2hAD1G+odZ2aYjtu/GJj3peNZqHI9VjhuLrUOlJrLX3/QHZQGEQ8JlOYrBVA+
BLrocC8UXJg8N/vD9fvlnfJ282VjkVae/3j74VL8ZYrSwslXwIcVavV+WGvAyD7j
RgPGNGXFxfvTuEWIbGwkoHcTPCvNNmZzzuq+Kr7gsQMfuf+9hmok1CS9mBr0hhge
mMCtVFCSXDk7H8/uM12qH1+LCe2/n8sUXSuPaQDtBavymPQ0ifaw4XGfdnUqZNAs
GQqk4fZdm79H0IJBcAXC1h2Xc9izdkiKjnpgwttPveLCtZwOF5HIyInBzR+I0U2r
YMhGqmEwl+PODpEHH0tLlmOI5o68BG0S8F6/KnVEL1/Zhogas5+hhS4AID2DC1vX
xy0Cm4ABxWCiFYCYuHFNtQAKTFTbfYD2zAoGoliW2fkzQKTBSH+LFeCpWgz8xk4V
wq0VzwlyLOUuO0bmgFjvZ0wcjISdnuPK6EGT+CZY+v7bRbxbQ6kJufUec+kdAoFs
rj5z7TkFyMrWFToTjd/AnfbsC6zTdkpVi3q6LDODK9d1MHB+tiIqjGuaP4l1EIgY
irC4yY95rrdMNH0BulhA6OiG3hht7Tbf33d2OoMTCVGlDgnmFgTxnnuYVkbIPcP7
W3+V6/SSjIFKdZk4ax4aUDuqIHSfPLaU7I2Tz2MyOzZzLBngSIXV3wN7Lcqj7iAV
THhqlG8uiVJ6LUhpqCmn1rTFgcN2oRX84dfeoRGoUMjegFO0kAsGAvyz6cbE70+4
pSK8BKO01gOT4c6BG6gwGbQ6l3ehmPReP5zyMW8TduVNrr1sFnKoJ/Zzf4G4QtzK
Gyt1Kd4EFViJthQ2xj3F32wv4uXhCDyRq1hFGPdILgL7gKDJZlttWYCdKi8DHx3R
28nimPX9GolRLakYwmj4tQGfHUxUsWsiPAqJ3GXFMgXR+uklWeTlsw30urUGrS+E
oRPA+hlky9RJRUKG8LUfGitm9GonEVlUGXObwqtQE6FBPlPD90jhz+mMKwaK66Bb
J9bRwb6leZPdfaBSHKUrd07b9+U02cqEVMknFiLybehnvj/gi+8Wmw1s5kKl2OPP
T/3v6r9Ga+XzRpP6bTy1BUcafyqvKD10C9Z3AFXx+1KKbDpl/P1t4gJaRuir9Pj1
p6Y2INXfrZndADE/ff7p04iK9FoLp2zhu/Nh86fr6lGfQIfeKcRQwkaO6hfZ9y1V
Iz/4mkEUlydSn4UvDAEate3+buk7/CEHlK7wTB+qJsklY3lOWOgT4vC2/VVsknzX
bDuY8DUleYCZzzkFVOFfjcQq19ZnZjyEcVM59LQwj/Z0a1Y4LhgOIm1Lj5wUhTos
Olg6gN00iIl4plu9B3qwZCuHpOJ0Ra8GIRTmjXTMrraziqh0M8HKYTXYLcEGj2Qw
/8gwZn6MyGxzBrTkmypCe3cShH5B9Mm1SAy/sEWe6HzqxFHWjmC/J2ogkKMB3D+x
ovHfdZL1/Rw9qFX2OugQM2fzxumSXvc9kN7IrVt5q18MnbeaQ6FfEbYG73BXrDMe
iDZbt2AV2tSNNpmQYccc8iUAPed/+zxJI89ZD9yu3LAdiQymoG+k1A+21yjTOT/m
nNc2da8KHT2MZoiA2dbzkdpRzbYtgp3uJ4k1PsxA466GJuplwNubibA+txEoECmh
xsf7L+FGLJUmKDGi/uQIaL0XtnzGHPlvsUPtMGuR6JsX8/sgt8G0GRHqfUeoLY4E
153IKh2M2DtUEXo38SHcF5adT7tbAgo8/cfD4MdUrdLLFrPGRaf7libwNG3ZT+Hu
q3noSZ5hm22EwrcwG7hza623ervoNlzGiUFQIKsOsBn1SXBAFeKVOO5yttqT/xj6
rsjmmc9gK8DSTTSiU4b5uijL2IS10ZAUrze6jxeflBzu28QcRtK8E8iafDMpj53q
DBFeuh4J+S+I4vfLbRMWCDdwz7aWNfKy11rLkgp2wSYyJrHkf3g8Eu2U6ra0XLlh
TjSRxI8pZiNLHGOfszroj19fHI8NGlsWl7fWjkpmVpplrKar0F4eOGJPxpxVO+8F
zaqMvr7+3d7iwNraknUltyyWFjviquTw8rDLIdxqqRNntBzwZldzHj4jinKgDkZj
sMTuoUFAk9fKjNu1whbRzrLgZCNG5DHjkQCzDnbi1Gkgcv1IEmwyXYd+g3sauLyE
T9Z7Ztnkwd0GpFcIycIXi05TdH88oo5v9GKQPJionnu7mE8qlUYTNND7upytstBg
vSFiLeS7qnu1Ua7hZEBfIc1GIUjEUaPxiIKUASm8bd23deywNEvDdXzwdw+BVjPB
f/1Gibubvz5rmguGCoZ2XDx2IvMPsSiu6DETZaBhXuq+zNJ7i7BA7d8lnPE1LQzW
Xv7zw+tlH0lvquYqut4L54QQYcwpOktQy1AE1wa3JbTzygrb/HSC5II7ZIkgulae
MZjaGmxNczkGBgDc4J2QWa4bHperAKYK6KVgw2Mk4CMyMVcLFNg5+Z6QrZwidvfX
ML3PfnChADY3pq7mn3O2i0ejbK8xI+PZzT66NrS+KrVk9n/+VWS5TGTw8L9vueww
acJhIppDsfrXm9eGKtIMPoQnNRQX6YWi2twT2HT+n7Ui9xMhwhgY6Lj0+78/LaU6
Blh836GaaWTTthHKOXtHEDJ6NUDbC7eSraQvOcM6if4tuwugEIEKsMmUIoJFYVf4
JB3B+JnyUc4gNIHp0FrHNiFlBJQruio5kNsl0E7DM9iHAVmruRvgitk1TyIvv/5+
z4GLEU2AYGzQu6lBuLsA6W36OWtytU3QnpWdpA1FWkIP1OLW5JnRjEbAJ+8lj+D6
2sQA51ugnVE7+7fqnnduWoUsOtEeMyg0WK501LC/SCKYLuDpuDb9j1ilW0pgqwC1
bRyZ5A2SxaLbTloszdgkkX9SDj57BZYo5/n8FmyTHb2J0lvZkQqMalz4NUttrnTx
aSSJoe5vjsDGiDoEZdIE+mrcsAFgK/lWrFXiXqFsYlV0jA+rZPJHoYJsU47Z1H3s
Sd9pXLMAsZE7+o4SqGQoEOqf01QKBPqAt5G3p8dfdxbABLPhXztz/hg5Y7cUizir
L9IHxhPxfay0Wa1VBh+h5aWJOaoN+FR4DYFpF+3BDZvkvhWB0+vel4Kj4M7Nx130
3wHtff/AxKMKnRoB8McbqGLkWr8+5xQc017vfLkf6ISMrS0JZMc/IIx3VFJuDa7L
mCpMtLvyK276gpmk6JFJp31S+yw7ib3vHC9pVkhLhimHl1EISadlz4FKm3ERrOM6
zvznIdS4QrPpU6ebAQllk+SSsuAEeh4AGxtjXpdMhaTnVn5Itcg6H0zjgfzyJlSY
24Sf56VauxUmoiAhfdw+bxg8rZEQc/PCe9o3cRJ3bhEsGEJuLQlgIog60B06Pvd0
HxniD0dqq3IgOKA/TMj2bg70cCFYLQJ9cCrzMaCZOaMsZE5vvw9sgysLGrLzwOH+
j7IhNq1k4JcNehzj4fqeEQsIRwoYHpcVUi40/sT0Ek+LVy4PO/Cy+Mn4JW9EyaLz
5hHZ5N+YYJAgW+WuxHqpIaVQuoPjPb8Ez+VXbVQJjyTiJi6MCvKQse2VYGna+U8Z
rCLseLGmERg+B6empPxvvN1J2NSGii+oxWHoNTCfAt1ThbToQOGCOhKDPVm9hBN7
LzufnyRjixZycOyQ9kAk62JiLyIgjG5ir/zvKnkkvsXRQpxS36m3fhQLakTRPEnR
K+A0vq6HJJFe4J/OaWTlj7G9pMLNBUiRYeBzU/JVtOi9O+B1WoKm5unGfjXzfG+3
X5bKbyeC/ojLYqNBgz5kleHn7LW+9yyKYt/6W9OT6wYPb60yPmMSD1EM3XRd0HcO
xhQZHaA6PunmDPLUi3H+nglhNXk8e3q8wH5pF8zt9xfZxWSp6V3YPkSMR6ZUQpV6
TB1xpxNaDnfn0z+tdy8J5TN01NTR8vCFZwLPOGjYTjpaHUqYdmkAR4/Hy3NiF5rx
hoDBlfF7LxOxg/EVBrLB7QysAN5LxRe6Yjw2mgP45w/Tp/93dAj1e4QY4FsMGPlq
wQuItPeJ7anpv67skWuf5+sh99UtFyVshYW8P44i0fdZ7QzdKTpgASKMNpk2Miit
QtB0IyCHVypsuo75TbdJn9NVwFgQkIvJqCugb+8ZnKfvb67U6xoqrF1Cw7wLWdDZ
KNwyA4zOiWBclGjcIibBNDHlGt2SdVAs0NxRZfP/4SPDH6N6zth73Q6oAzCkF8gF
XbTp2KROoknQcoin0F8CWR214RTLunwokoYLPe3iZMC7z3XG+JxTS1BzP6JnVEiP
/l7GnyMHzwHLslHMrn9iawV/qx1YwJn+4xfUbyJYikB+ihlAnw1qKWWrrX2PeV//
ikCHvbp6hOIyjsVrHUKPFCxIIML8p0NwjtLkdmYWJ5lZPeybLSxYLpbq7Azy/kGq
7ETGIX2+5tPAref60BZdl3hUAqUhGZ4KOmMyXwPriU/dlyc597LlehuMKyM14qTa
u1VUcUnEhOjW1Ns0Re4aHtkpxW9oxwFFYUNR0I2RhopUeYvyn0V7db/ySlhmi6jU
D7FUU8DYCAh/xisJkTuuGL4L9WbbeFJzflBnUPQIX5zt5mZOIiNwXcAhMJCUdBoR
YDS9LH0VJW48+aS1ev7GVKTKLXq8Qy+ZxCqYES2PRlySeVdePm+e0niND1VSnbjz
aPZBmeC9XAOyIvmiDxZOWSvuom9vAWrVvgPUoou6LKVBL95LIhi/C0sFtdJs5MMa
M7CPYryt5bPS3ycH5fRXVrZU8cvrJzKkb5UNcr4L1jq/nnVkoesPuyDNsS9BKicW
c2/5RLJpJSlxupy8/SCviyt7Lt3c8H2aNz7rL1Eco3gBXct/QdJVppfmtskZxsoD
94C+S4E+OSjfosHiFJoXK9ubUujuWqXExYlBpPP41IRDfycF8ujbZ1ZmXo4Feq+Z
nUxeP0mn6gh40bk4S5vqm28YODLnHpwIRpgjqEueopt86LkvFn6nWipuREf3Jsgr
3VrIaaDyru2bbwFMCBt3T//p3jcd4UGStijTuw/CL4loQc3j3dsnM1EE7pvZ1WUq
kHwt0s8SVHX+QO4ijyghpPbfUy6ddAKQlwH0WVpKvQuWVf2SuB6eGqs91m/PUv4z
0GUS6qnQaP1cplusfkSBwwZJeI1of50EA8c28ENZzc6pavEQjsw0gt3NN+aYY1zD
J4/aY/eGur6t0dZBDvK0+pavbw0Sq7YZ0/57crQe9s0HKXPlWhLXyJjd3JReQ/ER
c7UbgeedfrKyJ5xTZXLxAXJ+pYLxQpROGU+1pb7lvZleGNqUgInLcCjtQ8ujQ7PP
mFIZorbvVt3l7TdFrPImeSM8sYMpuyLTzUfXywOxLe8PDkH3xxkp7Tgf1+jcHAfP
kjI1Gk9qkHjAivziRTRtqNm0yX1UFO3e2bU+ApTN8z2pUBNYub8rgpZRYTR+NV7A
ISu/jmUaSBIO4vWDfepb39X6fEMWgMvUZzUR0abzAjPd6iNH+eR8icH4tjVzWmx9
pQgMn6n6TfC1YyAKasEAAy7gXkYWVekGpDow3RoAHfumQk/RVMa3UPTtiCG4uJ0j
vvumVhCWFC7JMFHGtG8+1THzyLOEhFNUyNfDnBQzsVF1qdtrVym+IpR3ZS56NY7g
49ncjwfhS2N2DVYBB7FxACU62lFkegw5r+fGA3ZENmKUtOJxixZEmN2oLkBD8DhQ
hS8hvgM3zsafOFWaiaErgf7pqrT5KwkNjfTuc3pwM+p/63RZoTjb0RgKlSOG7/bN
kvH9efM7usK/iLIWEs0ETGpaWnTxecfSIRkUaBjoX5+kgud7/7npiEyUoHKC8IBC
CtAc8SOcuu9YFbLkq4USvgThYdUkTTGcLb5DPnqSY5djMgl6lytQ69YfYDQIIJO3
N4/jfS/xXZqGal4hzFgIkyb3BHoNg9NWpY2dKN2P0FLoQlOvC52X9AhXx4hZIWtE
wCrThTM2ZdpVvIGT4i2WUsbdScv7f6cD1M0i/5MeCq3L5ckyHDjVZ73GBzXPHyoy
KULb/uPCjpQa9b3OAoBOGZjhodNlEhu67+dJPH24EwoVoRf8H8HyuVV4HH3BRQGm
jvTwkjAN76FkbZTRLdgGHk+6RPiJaE+j+wZujSKNfqE8jate5CbTfWOrlRczPu3v
eL8vrtHlPCUqlfOAeqxbK4448nJYN8iSiNs0t7PqYWNfQVbRKx4TbcG2VVmZrGFd
6/ZBAxlk+CFMK0yaaJAQmQbAf6C0W1RZFXh6Lymccv/5H5rZcdbex4zxTWXikdbB
cNzl08+YQ9tnfms8Lnn06TclxKrxb1APl6CRTE1ZVin9wVm3hP8JS+tv/4y1e9+g
A7VoRjyFhQnFqBlWufo10VBE2nXOWXvZBmTwD6gmHu7CDUdwK/PVkkF8ip+LDqsH
hni8xCP5PaDYqGmdkptcM7D1UaqJPMxSP3qGq2zc5F5CgwCsxquxWyDlrowa3EhD
Ma9b3NKhPpBEvREn34s/oChpVvo4ISAQRUe7FeHTZygkFif+3YbqWfU8V5B6Znqe
fsnqYJn8CbnR8JuhA/MqSYlTxz53ZZ93bwGa47KtgJbhpuUKKKpU9KvbusXDu9vG
xWsA271JY5BHKu0hQNl0/++mewa8/yvIhd9TVaFpM+8sliFWe3tGUG808sc0Rg2c
BRbRCrGSH8swG0hJj+l2QdxbagLdB87cGLxtnIRpCYMORRYGEFoaxmXnepwFDRid
dXEs8xXZV1yC3CuSgeHHfkq4RCbotAclxC5tLefbq9jnL5O2nxKc6PUHukfmPcrR
SKF35pVEQyHStZu3CCBlK1vBiXUPefBopfm1/9Iu5vuNlN5kYuLV8etlhlGgtYip
G+gz9ny1lPJNRLUwVWu1rDNKpTa38zVkHk9GdveE4UyAeJvTwIrqmKMmmeSucEsB
G+HxCSPUaMJyeuBUKO07hT/Yzt7poRwB5IqiyozSeolR3E8mazsXHTIX2D3u6PFN
4cUCv3jN7dSURvX3neb9gtD6IMpJMVR12Rd0w7erlh4H/0RwhXBpO7Bm10ldh+Je
qGjxj/8LFQtBssGOZOtnECW7xE+juuloudJ2+OPGP78IeHvK5/tWRfnQlx6qioSc
czZ/YFvn7Dr7v7KYcqBg0TB04skecN4N00Z9M4Ozu5nwGLJj+L243g5LRCMcuEe8
mWCXWxJ3BXxthQLckzYeZ7GwMJUtjquU6xKaFcAz1lb1AoNDkt0SFpBFkSZkHI+Q
h7OpL3PE5RMUa3LjzF4E4DH31HHWMNPqasHiIUHieW74+liQyMqfpo38k2+j5alO
OAPy+0f5MaiO5sr5m7L2tQ2/7Fcx2wmAdlkpyKQhtFpkK3wT3fB0W0sJ8AJ2xwcY
G0BQECZmai4AdkhUn0gOk8xchehY2IdNt5Tu1tc+m96MB9ZEtygn0cdFFqIvO9eW
6kRD4AyFRm4KeaU4s88DW7+PCPE6BdlEktNcB1O2K0fQP/bwM9phn4G6SuqIkFyF
4vkOSaxgzZvpKTwKcuLYP8l0S4lGX+Yhori3VtuzMmpMLrhs4CXgJLRXHl1YXDMf
qX7/FqSbjLykHaqw/it95jM609reSaLttYN9aiT5X54Ji92R8Ymy8tPEEUzgYtZ1
TCDaSxYShVS03GklUkM39dw3nZk1hSGQeI35v1vfbqWNeRU7PBm+3ZCu/hoCkO1F
ZZIHDZ2bDktqgo+gTc9Uz9ZqFcHzzSpnIjwYZjQ+w+/6/bTbVaqZDEqDFY0uAnrz
FMwr86KnS9dmMpr+LUxGUu6UvyYytzIn330Wzj4yCYQuXHontzHEz4THp90uKC4j
bPJfOG2EDZTleNY4pmydjZcYw4vFF2wrIR/371FMhPloV8KPyWvoDgfgc1EsMIIL
BkTxZGD1uSH/nRLEwcb7SUTVVpcC/Ij0sicogIOnMT6b2VhMLHyKjmwjz5AUI0UQ
1ASla2m7NVnM5xak6GD4y/3VEliGC7YetJyMi9BnXdRNdoFXRdQaco3UWeDJJ5Ui
JlrE8lsdUwJmNUr6FptCSKpXHCeMcYMIx859TKjMNqfkUQE1jIMHM48KYp8BjP6i
otlbvn7xnyzkydtv58xkoYTJHoj4ARAsqCzmcvqNCV2K5L1yBPegdU///+Q1X0Tv
cJl0i6qUarplgzhw35xDTrUFiMPH+dM5qTWV4Vb0ZqcydZE73g1XnE2m2f4qVCku
ej2KScgn0Ix741epw30XW9+yc9FH0MaSb9Yot1fw3+qzZeKAGPmtIfOhcWYs8WLW
dIQ4VEInm6Del/RDmk5WxepwZTCV80PikztysfCjqLpwEmzoVt/iUXLNkby6busc
pd8uHpG57uX97Aa4tD2oCcwT+juOhGDSwvz1xq+rizeKvmRqkXn4+V/jQA7lHFiU
TNvdAJl64sKnqhzHHUuU01c8VxHgnvY91X4ufLWlU2dUnYhaG+Shx4qfoaaD3pAl
cczC5uqDkNatA/SMdOhygHovKfgx1YVLN1gH4w2Q+M/bqPbXnDtaIRLzU4qX5RkR
atKhlPLgtvA0AzTsv9f8mtKjKm3dUjCcjtn4pUYoo8Sb5blvkTeRC0gpJ/vi/4FH
sWGlkNBnZ6K4cvC4KMMZYqVie4TXcodafee5tIy6SeM8B/11Tj76h0c3FOXtOu3t
m4QGdCx1gZ99SQafelFm21QE3aW/4M0GiQz7TOAVxx3f+Pw5VZCh1sq6qPIXpQH6
aDERmy/pqE6oOQ2h7oisZOEjJjrglDajFvlD5gB2VyWcIXGNWKGWmnLWFYbsoBSe
2MpBBqbrTmZK95Zm8fVNQgmZFIlFs5hCYdHwV+NMDn/EZua9/uzodU4cctTkOCT+
l/JsWwVz6O5SaNHC1uuKFvu5r9cWqhj/DouWnk/Txs1PR2zupvD50AM8BN5GEX2N
c5LTCF704dkzJWQTpE40bDrEonNXF6pYzNmMt6qNJBOSEISlgw39K3O2+VJtdg47
wqhmn10GRXx4pZ0HI5xs387A42y/JM49gf4xzH/7PacaPYOT6kLCo4OJ4KFLIjQT
a3GQ+Vf+OmBXZfq998fi2GFZyPZ3FKmcqtDqSGiqLG7T28DxEoCJ83cL3+DmsA/V
0x/z2UvIhYe6XIK4FOICK4vDdHZXSw59YSTsgUnQy0dz5SH+Wr4WM8Bk+oIc8P+V
OBW33s64DRQYnwSZjjfm/ltus+if3hANehORA++aXpN510PzhcLAzNmvnvIBMz0y
Uxm41wXjYFCQc2sFFCpwp0Hsq1oai9jlHi5BlIYE06TQII1yp3Q9KuT1/Qb4+gxH
k3g8hyEWHHXpJ4ULXZD1ZI7bpcgCaqT04VcGeUc0fsGHShC4Rfs9zGApHiLEoTDH
1MB+wR/2JlisMCBImVQSlraPjcPPKRrQFseS4H9ibtWGbe99cuzmLOccVUL0PrUY
FwEqsysmJx2zKKPSCWeY3l52tFsrZ0i5tkyTlLRiXISRxBLo4gt7+RG2g43QYWGT
lI8VgXK1HKnNthaFDmdpDM0Fb3jW/BedG3/Bqb1wOnJ8F7wbpR9uJSD9WTVVFOnG
rd5mLGKXd7xGvtcE77hrHUW5rFmbRHNk9jOGcTrlSwBIPvxKSbvBg4jgv/Ce7pS+
mZlalrkxQFet07NESS6phpj4KkQhyc3pXeqHa2SY0cx36khszvKnICvL1yN/BrA7
IB8SYAkebTzzzF/lAJYacE1pcZhcALswu3d+Ti9b9YqOoxiUzRd4H0dHUELTUIDt
W2i4JVlJt7zAemj3IrjxqbbnqGR83I0YD0i/lN5VHZfOEqgmgPZY9tptOa4BO9WP
eYbKBr4EWCcCDf6IrwHcs/rTMGUFKXrJ4sEiQebrEaz6kUkCdDtHyhosCZy7fZV1
qFkbqkfw0hzQMU06DQRUSjJs3yeQoFa1f19E1pKA3UcHy4MW2MOpBL0NUPJH79O7
8/ccYNPwrVDHXky2Z9w6ZmVoM191VpGGbFqdH5qqls6jaLOvRpBdIeXV6xNYZzsF
Pwj1YaTzu+tJDjd6kZtdDYXmvZSXQ0f459tDZREX06bzx81Xg9xI/BnNQu+SNiz8
UBp5elHoBM+asrPYQeulRyuIGoKAB1jxzOUhtIIR8oaewC2myG2x9VRY8U3l0QEI
MkdFU0YJyBvOFpYEdH3PDBrXVJNoSCbLlBTjIpq8NEjXWPtUvkUXaAbuv38qWl0/
x6jS1OS2Sy2ShDyLMyJnoKEiYocyuXu4m5Kjo0U5rmJt+5VXJUdD8f/KyvgY5jHp
nE7AHtN3Y5goUPzsdFTJB6sMVPAvZNE5U6s3VAvMzedjIH5RD60tQ1zFPYPe/U9k
eJLIO1g5dTZPfyN2dNzj8K9XF3w6k2VPffVHO3WLEEX0FSy3tE9vCdGcsP3uYtS5
yWK6jX9W3NzSSPe/PtOOaQC83dt+3Z9R9bsCiu+JMeIcOVAX7pwWySdrj/wasIsB
M5vH82addbtXmNKbTTBXkqbmFiXZX03Cg6X4qwYUnSq0I6hQQhJRbocIBz014gfQ
n+1FjhLitoHeGqCB1BYVqXBCr/Dy4OldqUJ/yRha5/53p5heOp5QojI71y1ojN9p
EKL1m7wNcOtbcthU3uoQGH7YyKC+xPYAgB9l9+EYmPddiMguJG60PbCSARzltNJ/
JjDGFy+GPcodQbl76nY8SU21gQeH5cbn2QLT95DL9b9kE4c4VKIn5K0GzCZs1NKC
uU+g78UjiUNf9t5WLQTWAjiQSPVDs2jjOE0/PymFlkyWhfILYdb1Ii/0JmCS0f7/
pEKQVRglp35Fvnj+VCWdMNKPl24Kt0cdFLHW0gB7AJ1Tafd3QXOSKyyFnjLM4e39
/k5iYFBDj2V3H4OApeIWWTl3rjewzdWlXFUh5XiI7EDs2Eun2Q2/1IN0tI5IKL2+
kYzRTKFU5Rk/k4cb36SD+/USBrZ7/HtTEaqATWtAf86Yu+Al9weUGjICwr8v0QfO
b8woeQKFL6Pda2Vb9+v/fzFU7fbxgI5b3yWYGpKpWpE5GvGgfT0tadgRu91tKrRO
7po0/9cfO8noZXwHMszZDdonInIkmdTBv1CJdbGqUmHHdlwmFF+ZzTEsPyeCa20e
Ht+KJvKhqCY0UzQThs5yPq/gIJ9c1AvWw807Slro4EkOcfZls0eD4COgK9QbfVJl
T20/8TsBYvTcn/wGvZutwcBcwBN8dWwACwO8zW0c7I+QzSflGtAdKwyHRBQkFOgF
K9CLcFHVzkT4iH73gT0WLaz+qBanbXPQjy4Hm0ZZJvPlStLAzI5vdIZVQb4li1Zt
uy7PGaRCADfts5Q2vD/0PZwowoTHP3J+T3h0aChIlSsPgDDOCXvoBC7mO4vm87s6
x6U0j0DlzG9JUGoGCKKHiybjvFg/SV75VbrP3AMp+Ue/w9EF+uTXtC62XvSwwsdF
ZsMBa+ZbHsh5+1ZV6aZt13XMoyisRp73L4f/U3ys/WjYLxaeI2a97abM03pHEWkZ
y/wO1mXbTJW8gOWWpYr1eXVR6i1cRnzJoXdfL22+GTClfmNigxYldnEPamFb7Hjz
IVXTxnsJuqjuEtetJdN0V4baowSypWlRoi6E21bUxK99BmbiMWxWMPtbbuTomO2v
mR+VYQEciJ1UqH5BN6yl2sabsq8pRonzRLaG0mxJuG4uaT2YoGedg+aXmRBRjfEq
GTRIHiXCVJbFJ6p1zBpg8F6paWzBo3sdOS8XvR7FFLD7Li2r321iSj3ftSJatZZZ
fDVbINaORQdT6jFopSyKXn84DVSToexaPaWVJtEw695fGYes6loZPu9Bh9UF3JPQ
LruMw46wDd82aObgUIh/oPOjjBQNsBbrNj9Adfi0Huc4hCYL6kUzoByvEuxKiQzH
RrYVOv8b28NFYyypwxKoaL/pXh8IRRnRIqRfL2PtLFW7R7no6VyYDXcCOLxiMDwK
4uBrC6P6Pbv5yXWoxqzieI2JAXCEFOQ/qkfLIPlm8hTwR3ehSfCsxNBtZaRj/54z
K0jkTY9C/JHx+Ha4hRyh9Qruq9vAmiPbIimhiHoqa/mwbNuj57tCMMdOogHm3/0U
VfcuyVWvgoNw72k7A+qB3h+4+jytQnGXo831lijlmN+WjGRZ3AepnzY5vZtqj86Y
jdo1zTbFg3KcnmCAJGq0oQRFcu11wAeMY/60Db6uyr8S2zc6iZM/V/QCEDKW68sf
qLleec5DHkmAJOHQaYCmJD3XBM8XNLTscj0Vhq0IXO7swLoqo6Jz3yCBNlnwmHQ3
hWOPoU8vXMHnD4OQnt8FKTuLkjh2OCAgmxYAThwDcJojOa0DjxCs6LH/YPa8awTT
rv9t6KKtv6JMzPE6TDX7aS/uDimQBo/VUk2TwHSSesFffoiQtA65XBnjS8sggg0G
Oh94F5etfu3h6tibkQvbgHS7EB3nI8KsnPChli0/mSauAQ68UfvAbS6o6bDmtPIu
RT2uM5TSIA4s26KfmDalF8Tezj7/Ht6ERS3ZAGp00YqIJb+lfWKBQOPvzxQRmXCz
2e6hfVwKD8xb4P0iqTrO28pGC7krJSo3/fW+XLC2r4oWBEjacTJYXuXPeXiQJxbw
FUtlC/d0Fe9UDBh1k+lwE0b78k/BBW92doVBHS9clGpCoPpNe6O58advCbw/xEus
spOoHzOGT3pX50pG6cDtVW5lp6B5RgSHrEwsH/YhVX+AOPEna9ZXdMcfQWL3GiJ/
sVC1TLTCLD75gaYCO/BPysAviSwyBuGHQ57ny+R2TGenx+7cjgkbCZjuR41SMuhS
HCgtUoKD4Q3wbFVnMwNvhneDo8oMmQEyGNiCwND1xuTpujo6mgXLEuKIWIztbshY
rBUyrfdGd4VSKts/VTNb/0HgGVqbFPd98hPg+WDK4tAkCnjs+aoBVqwd1XzJEdbl
Y4fF1DamqNlW93x8Hiq/blhGRiLSOSCD9CRnHQJhPVXbmhHHUgiZ1WTBOvsVPfj5
cu9TSynUwI6JYjmbE781j0X+PvfkaG/+lshaU+2bfQiEDR7Jqh0aGsI8QCtDlFDU
+fSMQsX6xY4ezu++IgWcWHJqFoRXxbooMrWdBKVAftJDhWagNOGmLDeYe8n0DHNK
L2L01NMZLVcEcC1VKetAXdivvwAYutRGX6vJ1o0e8axgGsDzCKfIkH3j3cAg5QEe
+dKp5NksrzwIvJJuDrfMz6fvpjRqz8kZLAhQIDCru7PTe/HCKMdU07kY9J/MVAGx
FC+vefyY7am2YeZzWndIcAn2IfL7vCaMKwzmwdoq+ujClBQhRpGmEBzCnkyDsevr
DulzirK5BpJFYAufVx1Las+n8jMaB3VkDOFYRH248slW4jdKx4we4sWMvlR72a0S
17yqZ8muLqxTqPeVe6AoABjEjxxZ43Fvutyahh3JIHc3VnrAfIJibSF6hdS83cGz
pUyDehOEDmxXo+Q0uD9Odp/zq8gLiGcFEMmQtLMJQkH01afYqpVbVNP8rNpvkiNC
2N1l/BZUsGCFwPzD8NMP0kgXjwJFno0I0D3CWy0E0xFeu/9C8QXD1Dnq0F4GeFCs
/JJ5JwiHS+e/E9+vqxKzLpb80vQxoHEmZEpvmtostX5OElUYL/iUnUwkeS7GsFv0
9dQE6EeyZYD3Ag6g2uSOcCZZfIl7bpFv/Igeqkdo+EeAuUPkEDgjdh+1N8DO45Uw
211a38Sh/7GH1YYITflmcVvHtcIC7xgIAgZdneWaDRocuEeQ0u7vTydpdwmtcgi1
7EDNiLx6hvJ9K4SuksbimY59nd66VjGu5qj9Vo2EB8MjclzZTzESKXTGyMNv/KNl
rPwm8aUA94blfF4IMExFdtDETMNrkgAD2R9gG30xoWf40UruAB1XfWHzn1OO00N+
mTVih3nxmwQ3EXScNGeHdRY6KDaPZux5BfhjF90np4YptSzm1c9kjybkvXSgscDx
GnxPpa4h/b1fwZX9njjW1PvMB9x7V6e/jPX96x3OQsW7EEkNT5O4JAHPHwNzKuTO
jUdrkB4iW8DKl03onJfPGynuhao7dRVr/DfWwk+yGLjDMcp9qXxwXWwv330KZsNr
AkW6vbi14pzLQchBZgk14i5JiHMMzQElyaiWN5NDi422CAXOd3OGgRncqbBN3D/S
rMuPFlR0fD4VlfGYcDDyyv51tjMjvXvZUgdFxDgAqj8fdg51Kn4iA9tLCXSxxQYx
y/Km7mU2JBUCIh+frhDxEcEfbW4Hq5BFEzjj0xTqu/dKjnJ4b50Jg5EfZuZfCbAR
37JL0g/CL5EHvWpUsRtqm/vhBeMeaL8aO2FxO/7jtxTS0N/x9DbBv90c0OQYMs5c
ih/UMRZ8yC4RzRj86+/dbg08xX1gIyQHDR98F3g8D34WozFRRVlzaTCj8R9GvJqj
pKn0E/ovNEoVwNtYjzkg4smgOIuqqVHY7sAye/VlBtbMJrroDWyqZqGZBqGVuBw5
I3cqLdUKUB/MyZEyOKjx7507tzfBJWpt4QimFHMBW15OFrFMlHi3EzHIe6zfRRIP
VoEeNzv5ZPOW/WoNYUm/wiG8wkHTfP4Nz9FJ3uvDn7Tq3gDeUong/ZVut2RCuPPX
U1R4BM92IuzRx/hscfwUlw/pdA0YNls+kkIgBeZXhc27YrKDEpZFHvWCRAtwOHUp
cjS7r/Lgta0gdXTh4nUE4D05JjNNFjfq0eQhK8yaFjaKa1N72zHIfb1PmVREKLMD
kVugbw8iJs5fi04YHtfnFAE3ghFh5rRU4iPsRoO5ACBNWMF0eSG9gwdEJEffSR5L
SkvC8V0wUTgkb3J5cCkCKvCt2AtQDZoW/fFkR4Glq9BoedjWsOrJ3sZSuKUtNOxi
3AcxWRBxdnN8o+hXPJ3uypYYWxFPoqincdDBAG6qCiXVwJ1+kIXR/q23i7XBsBWm
uq7Jq2xLbqPghiBKPXq9T/kzDgyZx8k9wGXnWtM4Hin5MMBshm1OFYEP7jUS0mqm
iyUeQYpf2biH9GbCUU1TYT60j2Tbf5EyUqvHACguYUK/QrQREz1CP1aaGMbitkEL
+KQlrlXVNrPZa2xeQ036BthESkuqLkYYZZ5VyvsQVrJMfkMVpt8VVooiYGB+I9ZO
kqEf+UUY/PP4Nj4wZlh7ImTEMjYJ80yzMFOvkVlFeHOzd213gtpK7itg1DLga/bp
3HOoJXhVtV0t0PGmxHkJbJRhPsfMIcUMpAfrnCUp1gkblLpFOF93++nj7xq8yQb8
nl2aEJX3Sv0CeITpLCVLO+d/WuHxhbXCniExkh2fQ0yjQEzeyR4rGus6QLuClt5l
fSJ6Xj7Is0a6vIzGjb+NB/Ezk8/JluuO/EjcUyZoZcnzV3VR4H6eWdb5TF8CGSAr
vdgRSp1dPUfSmVao0itYyXQEpsSQWTZqFb0EdnwedAgvLHN71rPbu/4k+5hCrT/7
0PpPTvRtdQAt6q04xWozsg6qC69bVVwiWl8yFAO7ibtQ1wMB3JTmQnA2emXfc110
mbA3U0Bijd5bwKRkGeLdVo6W3sXJncF8B07WbmgN2QGggK/R1YUIQI2jPNd1T2jB
oH8USyh+AkisnX+0/1jrwrGMk2tyq5S17kWjmoPOT5EEjok9iXGIs6/yp4zsWfYm
QKjLkf+5baTAEzllRA7oM5Lf+djPtM4Qk0cbjD/obrUqM8dPO6GDUraoFAx7TAsU
bQHRY0sdmbESjA85hdepnJlCkM0Oydu5nXE5RS61Yz7LJaT2/hu96z1wNNLiGtWM
LRRVdACKjUyDmFiDx4p3B7xO6SwAO8ddXJ7p7+QCHxUAnwwENdOUNMCo4xXdRvMT
p/EsTwbbG+/PkZ56fS/bQTw93pWvJYxGYC64GKTLOKpHKc6pIq/1y/VRPip0A8vk
1GEYkU/r+8m0djc1O5HK9npCLr1XpDhQKXvLTqZ1/8yB7ulvI490eDdexI50axjp
3z9iYadXahr1Mn/RFvqCg1PxlEtI+DVpE6PbrjSVycZdmDOkYB380T6GRbz2q4gq
KOLEHbjZlMNpPflDGTBxh6YJMtR/ZcWr2st9JMM5iseQ8QgFuBvJuLKBxQ2/fQ0d
1VWIeFWVpYcFyuG5ymo3Jv35TFaJTm3TXbKriT4s8RADMWEb9XYBx+CgoHCiei9d
sbU8uMob5xtFbgTgu099XmhdtqPuD+yQlwehpzfYNHS0YXuaOYN/Q/6e25nDMpUV
FI6Mt4ilky6xTILTlK2YmD5nDmnFVKStJizsOvTGocGJjk6xjQ9Q4gcyh+fTnX/P
8aoSbZg+oHElRoqVKpITwp1d6GeNnZty3Pq3xdDYvBjHVbPulVoQBmxG1//6Xa3n
QeBQnI9dfFWabrNqHY9NKJA2Xl0YmXxHj7vLIcPWOlLrOKLtQXJqwOrEzPFpgSXD
AYT9WN5xUZc6XpRtx82bwHKwh1kJyw6WTgAemIZdVOF5HMS4VJAZs/HuRAVHXu2C
0VYOOgXBBObWbXlGNU74W5742WoyRTCn9GXWQpLd8UmksIOO/+WJoJUiukViGuO+
YVzLTtE/TVHLjEok0U3FliI+0jLmfkweeOUzWHSLsvXiQvDxP3ZlsfNJSfCeLJTu
/mVF2JJB23wEK9ppIjLvyU+swcnthn2oc8GvXNZFM7GuTDe0CjLK7BY5jlUGEd+k
Vhv142ztPQadxUzR5uVH2jcdxeoHJtJIWGtgmeR2xnYPrdUH9IHe3pc4E9m4RBl1
V9vknvrXC5f7xYbp2qT+wPpKwq3if1A6qK8ip+yqlkM1Q4QnZlGbfn0Z5WIt5MeZ
AT/Se9GBUcnA5+o5XDfc3s8Xea5jbLpUz2MEoB1B508NNDbU8X7pUAMLkShogyt3
yOLadaz1MhjRVpvbTESL9/K8U5Vmmjny8dmo+lu1BCbZQY6xl2lxgzYPkIGNz8wC
mrOMS1qk6PNQzHhFh66TKrLJjNdbKUXEMBL/9TZr/xOBrJyCSXZ5WkhaHHWeSFHQ
MseDEVKEnJzrBdSs49xbSEno035Jh5UmHLisP103uaEzgSrMMvRKzDhuvyAOWeag
GzW/2+C2Mjk4wRQwJUB5lwUE6UYDS1o7mIvaxz65kMTE315ZiVbhquZkMBNBX7FO
/KB59HI4rRxfSs80UO3EV3Jds4jOFKPXJ1EDdnq0jLoAqwjtuBzr0ZOsm6uAs+TY
CEqt9AAMX/J75ZeRiSsL6Z2ij/DdsZ0ecafuj/2G3D4gDKq9Ws9gBOPINRzfMOUS
D0ymBDGchM3NUG54FIBCB3aXpG7Himi08ritQvLOx4Qxn4Yw4fAM0WUJKz+qP5oT
xkLVKMgrb+dpMXGHa0R9pimJk0e19u/bFA1PgTEjf03XF11Qsi0hFvSojbwl6YEO
zs2eR3v+FojFBmrKIXK7Tat7oK7lihF2F+PJphuLi8ZepSTQiKzlC7NhbNAb8VAQ
PLTEPt1rTCTGkEh61ZeX07V7rKB/tqYs/mfcj6ns4rGqE+GJWh+thXhLMgw6GSbH
bgSyVm0nw1soGQxfHUVii7PQTTek524Lwf+CwygWBHVZ8irCjLTvIsUE4ha2uj4x
2TI5AbYomEYW58/cLSYPCYIkpYgv4NU6X3uh5PBupx6zXjEoo9Q7cWzxmgv68hiA
ATqS2hNMps2RJQ7VUZ9aHUjIgDZFgvJ0wFDHJSgV9j/eap7azhNBhzfc/R9EIyPa
OC41wyb9MatuqMYPO13Czcysfv+5WGvqigMuaSDfhTCrO9lmDT4XGvr/KP4uKdfU
VMcM8+SsWGWg/lB1Vm8WUVfUyi8+kAhV+IjhRKUME0GLmZmnRWIvw1UeDZrTEwZL
v+csp81vS15M0OHAxWwbYsYLC/afyDBMNnsVC3DAYZ6nB18HvxRCPgnjdiYJtfei
s6N766JmNaZOhuUaQEwC1fskmg5Y9lZMy6DYmA8pD3OgZlEEkB02gGwGMzD/Xf5A
NgKRed/XQYj1MgsP5gY9jrxUsy5khM537VkYlGjEbo5HzybhBhD1HrWtgFV+IQV4
0D1uK3m5sn2bz6qKzyJ6w/6jGqPOmiOaO84lzmyHC6WVY8vHirM1++vv+bmj+uAN
/vQ7LQ+0IeTcNcOEeyDc5SHd2h4kzztu14NWw9coxKc5NB9jarO4aVc85jLtAUG5
mrQz/rKDKscXGVyzk7M/1SA6XTqZ1iBNZHh91it/RL/XVB52CEUOgvSEbqfqyMP1
rgVX/rmTU4NIhZdU/j9TdRpHrm8zWpRyPDT3xZTZRGr3opAND8fcqsRznbJ8LWpC
fdFn3Rip+EuFkzZoFDG+DREDYtwF9wddSju5PzbkXYGzjN9WJVPZGl1T66oWENu8
/UzFGDiUvG06IBeEC4XGijsKIex+8zVb/erSiQvBdIqux1K+GyxavYFjrzZ69pWV
8PKG6ysG3lgmRlXq7cDywRaChSbIb5F5793Sfn3vbqefbBEzGxg4t4O1ZN1v0uoS
FX4wExVkgZ9QVaNWnJe9MFY0h5tOXDpLkEMRieJRTYj0dGoOcF0tgAfQf99zqmjO
LWzCmVVOefzgOHCMqM4n/SqgeYHhvS+BJ4e3iA28vkxAk/QBPMnkP2aL5upMTfKs
3ZkkvbabMHl6/seb35z6Apq2ZbSG9K6XSLl+iQDXcyXNwSRRl/6Ng9LYeAv6PIMs
94gcxev2bH+fSMn/i9rwQPATne7aBOU3WlkDe5sD7SDbE126Po9gU6UhNn8U6ijx
mLlQMe2CSxtJ92tyxbbcXO8Nw4p3ayNFwAF1varA411ZFoHpDYu1w/0PBs2Gntxq
u+V2stUA8XpZ0Id480nw5kqACU6jwdel1MasbeSfSp5/1TINxrlqqipbn+QJm8kL
VZf+eAz1R0P1rTx4thsT7yqCrw9Vw6gY1QhxTvLO98i9drtj1V76SavTIhcFhmk2
FEyXbcqd9GB0cRnQdZYowCX2KSvQxxVB3Y3mrySDhN4othAbtgOQxGYHsbY4x2D5
GBahFF0V5BAuDQew3xysNLHINll4E7X/GQQZNNn0oSsk9uFJW7hTsXKgVhV/BCId
VZ75Gz5LunoJmQH4dZxEpI7MnyvTP37nC9OWNNFAPoSQDlPx686NExKD/7eR37nm
ZCPnPoCfsTbaFCQWXGPJtvZlfNVA+8I/gb8Ck+k9AZIhBa7Alro6W6fFAY/flbd+
XsKMufBC1BeT/ZYOJw6XEzm6wJNCSs5B3tdAaOqH5ZaQeeW6Y1+JJHmySJ9bTIYu
FQ5ntEBUgjzVuLRV1TDVR/ig+so0yZF1ugmEXu7veOnQd3cKZ+mdAmNAHhMbMiBR
NdWkbVKPZJzu3qF9YiQ+sCSFka4eqO57z5rXd51duzkEbCmd7U6TNvMNMEu6pRT6
Cbv3ilY3bYgm0F2fjUdi4DhDkddaxIREHfPHou8q51k5XP4VlJdtEyxH5LjgiqkA
vNW9ATr6nXyK9SrNsroe//XCkmhQdmVcM/vX3mUfqermUdVKzKx7NBlZLVL2C0vR
bYZMJR1M3YPGGgOPOwHuHPyhiijru7R3/raXPRCRLmRzjQwzkVkAeot+ePYfYSsT
NpBVJ0c4RkkgmanqybY7RqqUuWE8jyf//G0VlNQe7XPEMEevEBZNZmb3+OkY87UI
pGYe7KaMr0pFLEv36me9iTUPLpg1G+Tldyhdr/sfs4Q51dLP+TRSkODVxyNLnTr5
9RdB7Xqf0fOi3Dgy11vE3hHC24jYWirNnY5Ie1lk9ScpQZQG2zk0mYHHX8XYv25m
C6SCv/b7MUqwRknY5UkhKO4U6yXluH+0e/Abx5btXvtoPmikan6DeQCnmyucDs4w
at4THekxuDKqgtvxqZPJQvOomR3iFDHFb4Ns0fDjsBBfDDg7G0SL7KwqzmkJazSy
5SfJjMCgtO4l2xgXhr5+13dimCoZqGImXwCFdiHd24nUMca/9z/R0y3+H5A+5DQ6
TJfVIjI6f7qwHE7rViHasS8D/G+Y7VfzQGe0UvaAIfCwrM6yqChCXD1P0O/iBRLE
z/zxAHLmwi3/FY/xcpAhrioNgY2IOF2efs37n4tmeXCHf7yIjIdVnxfiyDS2KaAW
A/6mwYShre7JlUx5+JDkxGzIiOm9Fhx3Y0yN+noAAL82AMiym6qcU/FD6QnCsv6U
gvgTBGwym7+kexpTCOU7vrW+4eiXM+KeHcsmW6742jGNyS0OsxF79CahVnK08yj0
33U2kbZKiEkYvuPptOYiUUv5ShH+pKcA4RvJcd39e/JW7rWcL73Lj9sH3U3h2NxC
3n6GgahmxU7iYIK8m9tOFlm3GobJvJq2cR8JwdgiAugpSZDhxqF0IqZbz7jmqD2h
H9mtqKTFhc/rlReTnxuM0AC5l5K5BAAbL+CDJXceI+Sf9pLilDJdww3v8chtfSPV
V2Aw3ZRpF82YLSuGEXNJw9IXYuXT0gWkQNuNV/a56CVTSCsKeoyQwsfg3HqGkulJ
aKSsayCcLog4hUC2iRxxnnV04QDYexprsK3Guhykjkc3T9kpfvycFhX6a2lvC1/J
PGV+gr94ydul1vQ62A7Fh3TvJEppsL1JVFSN2lHs07l+QNudpBKv2Vg0BY1qyWlH
no/tpfXhacEGfWua7TeH5nPvO+iSkUvNQ5LP9i6H0aGCicNpq0B8jCRSSrQPHW6K
men5WRNtq1OVm9FtS529XZKjz5T6Q++ar28x09NCE7lq3UnsWqaQ4ulzk8OUokV1
kzI/Qzwg1VntHQOv+ucUIplYPyyHSJ1DgIBVbaKAJFQ=
`pragma protect end_protected
