// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Om39A9G71Jx2Xu/sPMbYTMAP8x5S4AIC/rrtVPnsdCNcEK07FhIqOH31HTjBNIzV
/nfDLqVbgq+9NefwldiTn0GDKVQf9z5wXvljW7IO0mxemDE+GWaTct4NQhLXq8rh
O+MK0lpet2/OwTK3Lr0MBw4r7rmhi04GfSjrRPzNY7I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8864)
jXT231OvHSTb07uk5RjkLv5qtpXNFpWMOgIQ+wxKmJvW0Avt27p01Xa9XtiZkqIt
tNFMsA8N0Sq2adv18ZbZO+ETcJ4xH08e246xEHcGctMvMphlOlZtrgVILBUKNGNn
zwQIF9UaMJ7beEEhw0VrXhQ54zrtV9oTlr5HxY5WwRIbi/K/c9bUwpEdAzK8WmSi
embdZ2dJ2KmVXecKG3eaC/jEICVYRWYuZ2NYjj6rDYwgnWZdLWfq4VMvjSBloO6Y
xwQbWy12Hjp+uhwX+Lx8HGEWVWYW7SRDOCUvs6CrGTuF53+2p0KmKiYvuPm1vtdy
g5h74dBlTCbO8u1bkHtSbmR+HWtfuX1FPk/fXpws7Yrf0joQTmBJw4bBPW3tfbDS
muFMFYuFMFjfNj2r9KGBVXtdLRZrdDUVUla3npkCBekDbD6gdCDLr1uldatqhTiv
mRoG4FtUlEvYHFv86fUonXsTGgSVuxE7ifzDXjSKBhjTDl3UwuMouQ41/Bs8ZrpF
U5rZ4DJdKwfs+0x/v+1No9mIgq+H+E9x/5aOaQzaeQYLsKW5U7nTK/tX1/sJB9tF
OaTuxBq6FGA4pRB/ezui1Z0DFIn4CceKIVMkz2Y+4umfR9KHTu8+etrsudOK/KQm
sPb7t3RGibH5ctrHaCCdT7yWzj39w9++sDj2G3rrJb0lzEKbOKN9aBpzlr8nrdZT
93g/IQmoG6OhVs6nEi8CfJDnHq4alVd6eXMKuYYA1aE6ed8jnswg28aWa68qTCYn
ZjvS4OOmAQqYQ1Fgn+Tzfa1rShm/BxO12hkUCIna7dGihBkrhzqm6zl9Ycf7wbuD
9BdzFm22ALVKWSgjOp6M8HBrdZ/8YrE6/5fiPbeTaOplMBIEsLBnZAZl/ErolxzJ
DgJqNCdMVbjYf77BLGsb+6crTqYqlPJwyAw9oVgItQHE/0OgkuuLXQqB6eHqLd5+
jiDupRhxhwFolDLHCj4nWsXkkAkeG99Y/LZ8OanuHoPWF8Ac09UvfWWV9gW2EVRS
gMbytn4QDPih8ybnWhiQUim5Al8f5TbFshN8tXBM7vgKjVz05lUWM254K7fZKYN1
ogFg1oUb661h4oSGzsURJBE/qeBtwEu+WLqIb5Z4Sz67O0n0yVAdp7hWZk3sfHI2
6GxermnP71a63uPnEDcocpLQ1nvlQq4KvcGQYaZq3JyY6RhEA5jYIaHUmprA627U
jmLnzm90X2yfZEL1dmK6w2n07FUyW+TR5Z4KQT926OZrVfb2ENH2aGYaK7UQcjgR
+3WP+70bv3mGk7JyRThib1TKSSkwL2V2sEsTp7dN1Pp/fnHA7YjkMdR14UWZiC39
vkh5yh/uIcdj1uaTfX21bSu5MIktio490p+S4Lt2rAcYtIhqQpIrsYPNcqbFcbMZ
hV9wqtHGUC/5H7ATKrcG2cKITxrb6GEL7+qVsvMWySgGaCgLhXFaArdLsPbGIwHM
4qbkCiHj59WmRInlLHjsrh21Pys9q1Ce+su268avtIttzOVTQl8aNV1ioJuzw50k
WbjorY1tchWLiVumtDQFQNLCqdT4iuXJo3olzV2nbbnsF/25T7ymOl9/o2hEfmk8
SFxlV4RiPu//bH7u9N8TnCbEwbKqF1Ctbt0vjwbOJRQycyqQJ1KgeBlP/DTAWUbZ
XUuYVbcvTZSZ/qoDGH6wZNSN/QBEGvZ8IwBvgfzcNfRIkfN8ku3LhX0aXsoSVcXG
y8G8r/Cy1+obWn/5iTgejvnVh5+uDaNJeliJxchL0OVyxbGeuXd09ZEJJhi9eXJJ
US30zY45/rZprl7RanqirMoIqATWhRRGxhKqLcaRaqrxcAP7AzNglA4qMwGChhf6
xlZivp6rCj6Jo1z2tioC95IaVIGlF+5s5KT1ivsWYh0zpcM6IFfhA5gkzD+96IfL
trkAZfHfHS9UL2RIORGPyo+p4QbfxkTT7/8rXgMexsTi9wFrDpyYwTLAwYaz8UAA
6gj96lf0mviK5m5ommr2aoDnGFgBlhbmzR59ReZWt0+Nzs/28OrOCuuPM7PLyMSB
lfEekRjZBEt5XJKpggngEegtA6ThYFh5IPzztFb4uuiySI95xKHHJ0RNBbfQyL+A
CJJbyedYsvB/hKP/FloWS/CBy3CdL4B8lhytaHkQODnyeSBn3sP+yPv7BZYABzJD
vbKHu4GarvMVagxPeiHI0EhQhf2wPb+JzglQu/zsfjIuJeWlru20UcIZYSpaLv+B
JGuonitTVWmfUtMuX7VYdtszQbiQ0TEYabUbxdMbyVXPubuPsasT+XdNMHTpCD+D
UuCLJgI68M0HWAL04vddkHhW8yA+KUbJgfAZbvPW4v6kBd3TqPwg3HyMGEenheN8
N3IyAv4+hywNW0XTfS1FpzJl2BvkJl1JhBFTaAS29YvBSQqeHPLgKO4SbPYKDv9P
ClR5+tJqOdUEvp+DPz1WSGBNfYO7FdV4jCFnUla3vu9iB03HtJjQsTn4GaIrmu5a
OvtK3z5Gwb5TNg4qSDn2OPndwzOhXBoiSyJOZ8D+qpGVRKzZBdxh2uumcQwzXFE1
ypzYTQ7uDHGviSp7JVMQgANpzM/vjy03RahDzG7RwaGQY3sMLtjX35v6jkkLPKQD
cVroMzhqRizuMeHJqUEFl5bVnVk0UBEMJf/hXqliJQpGYu/czuZbXmuOOxm5/6NU
VLg3WjOzG0vVnCDNR3feTVott9+mZPOWVwHZosYumnwEqg9BpJI1OrZMq1yk+/fV
UJjqXfiYm9R3iBGOZ5yZatSL7xDFFscPV/wLlDyCyNjJoSfI4U2cuvKUOtb/rrqH
37ugULgWJuIz1a+qT85AnMcI5NFDA9qnAH8SlNkxpWPeyaMPos13z92BZy5uXJ3l
RZlKb54xhON2FPx6ucASMVzY+J4Efx/WgujpuTBWPU+h7RFOUbKS6erpfqR+dCPQ
hduKT7MtPmtjbBsVMxtM8ToRzaHXIUS/b0kSLpZ1f4VkMHTWUGQKgzlXNOSMPNeZ
6gqgesPI7EP20NwwankClPu000/TYl1yBOcxrMg9Vx7Q+pysYfzPBwubVuVdQtjJ
/YXoheXu5GDQW9e6KmNVR+VhoJhGYzzkjQ6jcXeCQfeM9StoPMkLxGT7bo2tujUS
TJ+ULKe3fqEzNU4xjO6/TKr9b7oKteWp6ChnhgOmBrDeRf0iW07+NIaenqiC81x/
QizEoSzDWYXf+qOflgmMH/7zf+PUk33UI6OHnuWlz+Saenndfjt0j16c196Cdxxd
HKgVHSGD6p9y6aj3eifFgt7d2bLZVLKWeh6exYj7fW0rNv2AgAonoarVrlIbMVOt
wm9+IVWIlMVYxcMaCJi3lOVLxi66yjzEddrBSbVsZpZlRW0lWVJ0SH0EOfhchWsg
htc8nchA8nRZWsXB4OWsWZplE9h7ccoZkb5QA3dx+4DTizYE5m+TJ21UlA+S+cMI
3GtyzquZ5lxaRU+yCbCOnGM7xhsc84vGVd2292hkiUG2va2jACTwtxOUsc4ORg8K
hyHT1UIg7tEyIJAJaZxbDf8VLawGgcLIh+cYoivKuAEBLjY9xIxBfDDItTBf5i3h
oXe9WSmnLxwBoMHd64YDbJoJ4baIajx3XlUHo/ZV5+4f8syDD0XaZat3BXN5ClBq
8TiNni6kTiVD+mdkJZdFQ/pGyYechCvp1sPnGe+JJw1/u/JqI2a7GvVz7cSzZezm
cBPLRKPjmPn+KphFJVJVIRN2oUuQEX+PEfgfScuIJfSHIcaHbQLaTlMBC0ZSLLg+
5dl9rdpnPKPIPTgwKjdvQavrTVjzlxFO7QfmpDGhEYoO1FMYfKkfzChTGdEEhOCu
jAmhm8Ue5XQmxc3rEFtXt5HHNJtI9byKP2qCVIVcTWghYFr4t5XaFPPXE38+Shvo
yTdXXVpV8N5mKU7bqvq7SMhjzY4rt2s5cKq5Wx0iSYF9tg9mCAP5Y1ernnsNHE3K
LsIvLKbsK7WEKbz8FOcrHZtNtsJqzF1OcGwaBcuC+vJAlAVU2AvQ7LwHOojm+y7o
jYHuKHi9Nfywwrg7Xfy2JLJpI5LHKZcxWuLjN+lGel8P+IolNqkg2A6VdPeHFPp3
lNTwTmgqPBp+wzxuTUXfY02yBPYB/t32YVg8LCx0eQfk61lbaAfd564PnsIMI1DY
+wMPTlw++4z+Yp5oGD/CrJ4A2pI2Kz+IOIxcU6xvFrrwmjBqfaLEJTvaKlDvf8U6
0cDXGil+I28c+M6pvKsDHj2w5Bq5O5meEYTSGnIBV9J+uo2sJ9MuLJCCLGXSCHGm
iUXtU/fdp+jyvATQLzd7srqrd4TAt6OYvWO4KGnAxuwANGHidaKf6V6ibSbv8HSh
l6vaWMDEePCjgaoZjFKTu4zprkM+Xcw/wmQW9f40pg5i8c3+LKAVR6AdduINTMMJ
IwU3Ig10j3k+ARm1xnvPETvVH/fImBlG+ujXMUFfcxeuJTMGksAkctHeiv1uaRy3
7L37Z3ee6FNC6r7PIXSeb4K27e6gr2lSGeO6eSaF9DQAtTj3WNAYatpmX+2vKpTc
KrQ+naWrXJxW2kZVoKx7t7ITtDrDCsKMOtc6/Mk8JuqPm3MC8S5lV/jaMubHnsf1
9gzRXYRJOP80IRbFK3WIVcFA1FeYv7YZa4Aw9yRNDSsUZDNfrpmgStP1XH4DEHRn
kgyFWKcRx2fKtl1vxFxv4iIbZY7NoBAyO11r1i5eD3cnPY+mslkp2YlsESGHDbGf
BT22IkUNyIgav/Dv6d3cDBSumj8xTa2nx6DVcjpvCWUikOQcquCWr9jZO62O7b9O
cWr6KWwYHrC7tZMp9PlUSk5+rP2lwyroXNXWV8cES1Gn2WBkbt5qdVksg0Sz1OW6
5TKdz7ZFHBX7Al6egOASsCwFBxRae47+SGEvCAIM7WOUByn1nacIuvKMxBmTE7lp
00eQeaBl6W+k3raPgYif78Zb4yKPrgQlqwWfGKtCWSuxZuD16XvxuRbUzT3SwbRB
9XmcFOz2vlsSEjNXoQ/Mq5+7+/5Ub46AtXBUYlpi4IfVtT1w+8/PLlj6uzXRAq2l
6TjIsOp/UaX+8eV68x+a/9j+c5ecHACsXCJ5vagnHnllGEsskGlL+D3pDy3BkMaG
p+NK+mgzjRYr7alU4PXPg87+lU4RN8OOUQKQsfNSmXHxFUkkz3OXK+QGYjE8nPwl
+rnTShNpVPLFVrwIfyJ+7owufi6q9N9dZEbrJMqQ/Cqrmf/YjS1NsUsMlcD20mwQ
N9rpPiKQiFOgUbIcmGfAcJUbdjoTd0y6dcJ6aReZ7F8WFPIJ/dMKo4SFMSfnd/bR
b70J5iJiGimCctL5ATeedquIutfF3vq+xUeRQfTm1mgOUJpAgF7zGa6k2Th/G+cX
nTmLUbBBElIUoRDV7XtxIXooOjn6MY7J/3d6ZTdDy4mhSqzgvOEI1WkhEaj65t/P
NWStRQsEOl6GJmWTsTnthxm2Xg2jryr+5Tet60fnBz1fcd1/Sb8KN91FFSEbJ1N4
Ifb3S1067ka2sgdSaN5h5hxVfZDw8XqzMA8Xmcrp31YNZAhaqDJ3Kfe7j0PRWvmN
r8zsPSo/4jSVS9bV4cJMKITyoJyIO62lu5SoHVVmfHMsuC1+tMFvqzAfIoDw+3u4
zTNaukNMINx17Gd6D6HtOyuiURFg8sGE2QLgyBQSJdXoLvO+zTq5s1eYeTNFwh49
hTYojKtBVJ3qpbJph9AdBslSj2/LT0Rm6C36VudP+Lij1VAq5E758moJUvH5A06s
LyjlFu1z5fAFnNcaEQ+37UOoKXU6s8/AIHUkmZe+/UV2GALa25APu0l6nF+LHDSG
jtIOSj2cHtbvnfm/D8nOCcguzkIAt9Vtb5DtF6nWBDUadVIPtlnUvc0aL1lXybm9
6GHb2pR5SyZtzzCaDvx/QWVbcgY5jJ1dpUUCYyKjdiHizzefTB1F/BkZtljJT+qM
2yacqSfF5uOIHoeFZKe676gSwEiGk6uJg3uOA89IZGvpVLEwaI2FuWLaj1OPTxm+
g5H2vzMuriIz2K02jOY61Q7Xj5IeJcrXN+peplLuQ4Cs8oT+THpuzxTTdyW7ibvc
TbajNwAlR5OJ+dB47Rnb6x9KFyYWoYWVU3fbhWv8fU0HbB4joEKakJ+Otun5K/gX
O2xVO3wlOZiSln4kLPq+x/ndaf/zWJtRLdhQw+b2GtKlEGCGbJEm5EpzTnf1R4gn
uac9aaUBdBwyBbNXQU0pbudXkiaauFxZgfNfOcu/eylbGo5DyrPltyRSvW9I7w4w
ZmjoNs9DQAtll6HaObqhAOcI2nA7vCTPeGd/KzUNlXogykY3kbft8kY6vEyNcxD2
+4Vjdj4PeUsi88RK/GREeR9tDEWvC9lFjKf9CxV4ND5il5BFvUp2PeMkzKGjcNNB
bcLW93kU2iAilbyTz1v+KF22xlCMe+lJqWn06lwPAJ+3OXC2ZxElGA9CfrrRuC2M
Zx3DCJ9G7yRX3hXSndRAT8z+b5h8CkiS2VDrrY6LZpWTZ2LoQB2GykR4aM0lXXHJ
QsraM6FZUsCRsccG7+ce512u79pgld0pBjHC7azCHJkUFIAh9jF9XMN216rS5rmk
bXS6nBd8GDJBXIUidrvO3ln9i8t9qJYlsukDv9XsavjHipukjO2Er77m04LyWNWa
x8fPNVagG38ezT8hlvnLlpcYd/UAIXSdeuEiga45mIp5o2EZdRa5lA8b0IS5RosY
o+tBoRFfs1/iCZZHAXKUaPx7H7c3Pc0vf2tEs3ngvu+zX5FMOlzAe+WdKCK3Yghq
G7WUSZZqjakcTmjsB+fv8ri9R/HhQMCRD7bEZPgh39Mq0HvobXjk2J2RTOUMYiwl
Frj8fMacpaNbY1NnCnXfjeX0dKv+lNKuSWCS2NSiYhrH6FIYDTCbOGVblGEsA+8r
6C+rHYpbgjn+UdE/jyvJbWxfj4QrQyH2TsRlvUtJ6r9f9ipXxDQPGG/XkzOlGgu1
CJrzGRh/KT5C3Ry1LI0M4tXZkcbZZqH5Bh5b6U1ZVgRQbmGdkUK1P90EiuXfL7D+
d2qEfn4lGcZAOmNBo4QtczeaiCg0KFFhtqYuzwTGgicRVkHVatkEr9q1RLzVjXyj
LnYSKDDKXyxaB8Fz02wI3smFJNIe9DJml69gEBXpTD0cxaD+kC34TFmdjRB8t18N
Fs0lpQSFPvDnm4wYOLMfzyQz0l7X5sQ7isXBXd9eDD2y6XMyCXK5tEzxRMkkfE2K
mbzv5RaEDQlsJQioaWZgD+eyf/A6XIgA4HO+ugOyZalTL2C1CxmuFlFEaLCgs+3s
Mxnwte9cM0deEQC7KirhpMIiJG2uCccd4sIZPkVa6Tm5WUKSDNzgeBhjhras8uJa
Mlp5BwsAJ5+D2fn3YGxuAdG8J//kXjP3OezG4th38B1sioTypBEOJpWtP9F3/fXC
60ggEnC4Y0E4yhjIM1KSeKSTzFcsvD7nh5Cd+TnFNIrvPlzy7nP7cfFWLDjxn46f
oirvr5yPMPioXVt1GcxhSBgREaxSb9sQsGxi8UW9n+Xu/4AHQj/9Iq7TTaWIHobW
x+5+J+1ti8AxeKpQGdWE2USPwRoYu2Pk/RBqy3p0s2J/ZphknckBdTdU4MJ/wGUO
FkDv8KfhF9dsniwgxtSrjvjivmSKDxcl/loQe2WQ3CjBewCLXiaLtbDs6vupaQ15
cffx0PDPsaZ6km5wXoNBIIjK1Vwb10vQebFZfaE0QjRofXtmIuzBH8r3kWbRpfgq
40JV33bbVL7kswdF4u4QXpJ9lyuaZLy29NjAMkkf36FEiaVRiNfx7VV2rNGwq/r9
niO7+s1hgX+FjJjcOB2TY2zaBx7zblKroV9WCghMJSCzZDYmOJ6ENuT8a605Kxta
pae6zOQDU4Bb+VgCgXSBO3ZNVUWRBmtrWL+/58o/kSWtbIniR8jsh6l33Br9UD/4
c1YXPxuGa2J8F8ibdDJt17kpxDp9mwAWMAtCb77hNB3+f2FeWajKXdEEMEwByc1D
4Ew7J0XrDxcdyudQzn9h5ZEmS6vAnG57fRm8L3UqUF554/MrvofXZyHukM9LRXDr
qnCOiwMzaxLZcQ8enC3xRIZGGHhwec6rD2X1gKSnMougy84dX2cbYKPIQMpQmCNn
MX5+G4DbIIerhTVccBkCasndON7ChfBIIyy1Lt+MRSp42fIOwjfdfJjfDTZVu34k
d1WAmhtUNIl19W/a+upN5nodMYkM68ZCtgum9okZeVh6WSKNh5Y61zt6cWevKHMp
eLIVuqJJxaW4ESRVwiAmtE9T3zvkiS8KlZHgUpqJ5H0zlP+AHlJFECVrxbhWNcfN
G4YyGbAeaBDF+Rv0rf+aH4WIUoPN1Ds/55j7Ci+DxanhRKwfTDjoLJ24TcRHgCI7
JcJbUY1LnI2VflCL0L9kwJUpI0E8zFbwK7mwH1XQg3+tctcAnaBeyzHxQiOQrOhr
4wfSdkMfWk8mjFZWpwg1sGmCLTCe0h1gCUzD13P5qQ1FPV4hacP+p+7HArhpEbqb
c3z0gaQPSQkNJ+0IHZQuMKYRK8yfFeGNYY1yu13q7SJkhrEsy6Md8P/6Pm/RmNVD
+8SGkxrWz+35JhSnd7e36KFzy9ncDL414dIsFNPx2AphMv/T67zqfVrPPOfuokma
bap/Cq2H00Pz5vTLJd3lXH0KY37VRzwr8eIOu5lrA1oEGQLooCG094m7xKQ5Y4Ns
iemViBc7XOKZly9AxSlzwkTjSipnxtDRNcp8uH2jm9JVLJAzDAwsha+D1a05Mfa0
bTqx/CPJ76qkvAbhkDp2L5wAMHPd0UQKc58u9K7snf83w1DKsPthDm5+fcMEjWL8
JWxofoqe93MaajCMElaBHQMvBFmp2s0a1jokolT31ADzEZYDD5J8Q5rcY60DICc5
TtkzpoDtZ0HQwF4zmPmIEOvyAj8lOm82xvZfQS8SJTcGw7wWcjjgzohs3gwTlQiX
FuaSrcGxWH/c/hGjDSY6mOomVYYVqRGRjljs5xVm8DgB0XXsQAO5EBecl2N9sRbk
izOeyxbU8qNwTYrqftzl8lRtBAyBsDlfOZdppyjfRPLuRS/Dkzx/MGJs5JsD9KlD
xlGqOtKrwA0P1TdQj7qu5MzjgyWOTTnm6DombuA8ZyXyP875dlVWEHJZzLk1Jkkj
XBfptI4IimpTOsXX6VBv/jMp+N3YNjWeGTpgcpd/BRW0Oh/Bki7Gm+rCUG/0XYb4
ARxcUqEbuQojeTkbyvRbexF5HMEanJfYUXhKxomuuvyfGzohipFObuWRjYMe0A4w
M6zKELJgyW2RIoUac8rp1C4D7JV+mrX/ngswiXtX1rMkN9hYI/TqgKqQcIPKFzob
ZH7mFUJXQNJRE2LB/TUkp9ApwRJ7+pPUWy8LWYyWww15jwvecZtllLGxuvL38ugv
6WN1r7foUiSRfAjQNuzMGqIV0MrQ2nIYKuupD25YkEogTfM44gnBA8WsOmAoA/4t
7j3cee9sLT95rBHHh5wXtURNjcIl4zQvF6qoJ1Yel8LS8hEM/aflBeRSjFk+rFsL
ruKbKjbE48ke+AC3WLRcw2vwZObi941KL3y5n5jVXwfQDUa96eE5TTkMT2Q8PrFF
8PVmvknm4eAF2PfPFYb7+aOI4jN0l6p4gKXMPEA8qw6Qa9r6pxoUrru7HIt+0f7y
Siu3DPXYtOggADxqqkvNXX0Ne1loCCoIZwyAx0TMOdEaReinEgNI6PeNwO6gy+HW
CKfgvzU05Pe+X5eHy5cr+B+QKiBmlYvzaAuGpyGmqigBQgJPHpCrs+vkPdUpKWU5
VE/GLiFWEz9w1lo9EKAtnhJ2Slyvpq4Y9nQLVL0eG7hO6Ob8ryYB1HwHf2PJ8aJB
zAGSaEI5DGVEinBlW2TOFUm5CivaQXLxgWrFztJjzJwlkC1S3GNbyBXQ2zx7u2+S
JkqnPMzwWrXll4ho9TRsQc7VqyxYY1XwCHZ6NG8H9sYMkGDn+kIiZ2FhaBRVoXBm
LwziWF7imxIl5rTZvsFMhTMCK9rOZbWE6WGnlqy5c8W6dmadh/MhPh3nWJ6XlsIZ
zgb7bAYMl5rMGsrUhPRXBHE13mWPlgARY36xYDetUgvKw/59SvIzmDq5WQGCdwXn
I92QGiR8rg2ZBz25EzdBkZHdjui+DUxlfi5dW9ndD3UUkOGuDRJWxKsfddP3QNEi
AK7w7qqOnvUndh87yswm6l/BkPeupNK1XXFKhT9QtlwnPs+wMRh1fgMYAn/2o1jn
6j7IVqVXa+S1u0IiJDStMNewZewe4k8rKFNleuoR9YKe2aH4pYg2OhFi7Pb4GTPn
MjGWsaUfDBaeuhy+L5WQGKsnYNxV98XBmEYu+wsbWE+bcQZ24VdqwZk3DRwX0m3X
y5YVkQs/RPQmjEBLp15gDNsuUvRO8XhB7IbR3znEy4kgyyZDsKKurmuIAjcYjjcK
Zdo3wOoSJQmPYCptOCsfziV9V8bsVqIbaCBUqP6GgFz376If3P3qZoJFXTP/2EhT
X2MO2pyxpVyXeNPMesEcU14c3T2r9DCuw6iHxmVJVpKE6tN3rwr09DUd20BGnGUX
jfs555UDylD+EZsC9WDwGmuge3sZJR4IK1ZVm5xj7EwKwPMLTJIyoM5GXDnKlrDb
8/un4Re6CLLb3cT3KpOVikL24zhl5TLuo4qU6Gf+1VKypVlnGJdmJWPzgs07t4eu
llVxfQvA7FI/6ix46NpLIxcxV5OgcM+DwOsRMLYjCfh0STZlwWLtnnJI5mbwDplH
SV5euB+7BYaG0qwOjFTPwPEIZ5ccihhaqKs26zl64BZCtdTfZDmXslMDKvQNwWcF
AUjs8mrol5JbnYRvytz5Kf/odLWQnDM1j2vlgJrXuvyf1ZP8vCpSYJpi+SxdHm0N
wHfhIx8m3lxgLgcv/PqGqIi3rnptTXnn0K/0rbQfby+eVyi/iH5rwYcnxAyk/98M
g3El+urMao11lkgN+WkpFcUOGB7lyXMd1f/14YGwjQ4y5mD2/npXTW4/goaMhwwk
jMh0xKCSRBRyd0s74QU7lzb9z+JjeAsqH+/XQRisugyvxtTvoXl8z26sk2hGeH5I
tSTiAb57Bx3OmZd5II2s7A3dp2MJobC66wUXGkvkSpYDfcCV7x1McKk1rEkvB7zr
zSRBTbevJstiQIrpvLO+rfmiImfxajkKwfhXT97b/ZHLJ/yNEjNbac8dd0YDumSE
2NStFc/g1Iz3tsViht7kNzWgwHStJvfuqtan22H+XaQ5mP1Cd6G44mejz8GsBhvi
iIRmLeNBSJhQWlzBADlixxz7w4ty6nsK1rLV8oXH2tBTmvVNie8WDcYvzpzGZYgK
RcCUx6oUN+ahEf1vQnqZhePU9sNZ8MjCm8m0cEr/c42dsLy/jhOkAk1t5Oojrgcs
P9fwNJhLfe0gbA8KCKwkFhOz+8wHxBXByUkjGwTJO3/teoN+hzJZhWEv4cYhAq7e
J00gErqGuQ8ov8Qvob5Na525U6Jzz4dIQqovqGJIj+/gOfBqaGrH+4EFnumgDTWS
RPXtYzOnbqtMjZuLIZbxYCPCV+GMka51pBPkemtGCVFoa0Fren8d4dWfmlO0+oTg
ubgHxZfmGxzkdGfC/YqXe1XbImj11d9TJ5RaRbolR2q1RRvvb9PR7DzXEusP3Gqw
8VIpvPlMfyHQT+IDdLuF/YlleI+0Mt9HhNmDWDrp1zGpoRXQJVjNLZFbt5KraeSN
wScfAii32mPtHyPFEQU4O065knU9gY4E8u0/gZi2Pvndv4zm4OOB8oKbrdh+DBe4
AFnshe/WR5HcMl+Pr4rpFxq10xjLurbtUim7FXv8c9E=
`pragma protect end_protected
