// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t4lf5SmuUO7QSZ9H33TUGIE7/rG2e9uTTG93KRaXBLMa7uGNz2qo5uCz7dr1Vr9n
fHj7/PAtrzO9wjv54mTty5ZZhtD6N+Z5Ovm1WmOfflN2mWX8mUIsFB1f20Wy7OfG
faRyA5gwFgd/kyJhFlYfd4pi+pv986FdmWve7ynPjpE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3312)
yKiF3dYytAWslaxcx02ZvZw5ZiSW9Qld6NM78qYIgTC7Hy/nOpD5QClH1j8Wk0BY
1Y9AJ2HxNl9RclQ5J5htDIdSMU7tzin3WOaZqLQq1M3uu8LukeGlsaTlyU7tSHLy
Fdy6ruPENDbEZ7PmoOiminBwg1VPrbXZCFWu+CycMU43X6GW1QWHu/DtTiQ6Qf3L
SDlH4Ouq4N3EFDdAdflSBHBFvYrKWmB4oNipWIr+/G0bf0U4wGLaYUkm5yCzdu+G
p5M14xC8jjqtID5ss2yk5AytQjZamVGVG01U8HCUT4KzTaNj0gRxyMWrJh/JwWPT
j72blxQ00ak5fvN5mXipGpwsm+HOnoTXba7u2oy2uubypnWI1blJfQok28QZ8kF2
YSBqfgNCf/L3S9jLbGTUsDXIeRb9K0r5L35X9PWjelKlCv0azFCEo/xq5Nfh4Gs6
vYqFRQnpriJbVBbbc9QvVYt5Jr2reV0daNvAFPIeRaIqZU7Kq+Scyn+TrC8Ob/c9
lDOS4X0179Pe135WtmhbxXV9tAKoWbMzHJsmW9Ug9iE0Od4IbLEpWy5geM0FvDxz
NXgGR6/XNNBYIOPg4FlqQfS7GzX7Wxc/OiQLyDoepbJyT3nTZQMKBT9oz8NGLfUS
3KvL0fxmLX1RYgNl635ipLWBw2WfnxCRArvBj0Z9taiKa0CArvM9cTh/U0JgMrkT
nwEFqItgWnDTA98ucqMQ4dPx2Es+stI25dbvDiMsGhEWI4rEiR5SnUFNCn3l4dTC
89TCduVvyjusX8v3h9uQfSMn+/DWTO0opNxGWmzD2N2JSql0oyMonhJSqO7C9ZVU
8+rTS9YAhC2atroCsvy4CheyYhjZTdmeziEOosU/3brQvWl7l5Jtb4P/GWNkB25L
uZ33sl1nCjqKPzTXtngkPLSxqsQygnkJn1jPztLs79ENb6vw8NpCvRUxp4AIqF8r
MpZnQELmBGOMsAum+My3wENOuVWlCNMDX0SxWpwU6k+zyPKErkHPnP8VBlivNgMZ
4R+YPFr2RVGHu74CQawjw5Ll+P7F6KAO4VsggEEtTPdjOQnfIxwZ4QvXJjj9Uz0L
kbX4/jhPjz2sA78W1gcPNUmLYr7FOS+/f9bc49xOfh2Q+nYAx4ws52xuNTgMFo2f
fwIZo0vph9WN/XsYqHZ141MbtbhmcK5RuXfaeMjzTsHBwzqHB6YK7ya7HONx2vTO
XWEzM/9kevTUGbBHNaPJ0oZznQtfGFyZphxDJ2HP7CRczov15F7uTEd9VS4IDh0q
C5aUNGwUd88mUQ/kHuHMGbeZwQqouwPbdvr86Z3qUb/B474v3Q5cvjB1sVX0AX4z
rbdPVRvBDKiR33k/gMXxRI1CfDuZuMJ937eYi7a4RCWOJNP0N5ZuDYh+OTniqT49
R2hHZzvO35ctD0btdTSgouvnLpjgJlbBxMTUZ7sWSF2o/27TCY79BTCjgR0AW32d
yx0MiayyGsTvGUngIkD29Ad28jD+k6YAp4B1hbORFO2ETRoLWM1rk/k6xb1BkqQD
OByPUYx2rFT64k7CDVcgyDYFR3uhZUlEGVwfFoM0N/f5NEdiSWXo9is2wG0aDQOF
2vIaZHQJO9UbxiKOlxwLwuCfo137SB7yb/fdkvbnepkm4c4xIhzQjn4PgSHXJasU
vPZ5KR+sfPqSJ+8BdG07XI/sjIeIFmn6ujm+bUX2u9t2aMUh6X3dTxdiJLv7GOX/
Nq++NoHvOrAGRggdSsZKY76PGFJ3Vgw2ABRspjjmRCkWaGoyT7C5tVUIFzvpv+T1
k2cDeALO6Z5sit8mXqKr8koON0GDkBVkzvxazwcWiP21pQWBwEqJzZuI70u5kq79
K+G8l7uXgtim8ALfqUYanvSxhfARjbGweBVC55mP3rBbMgeOyymdxr1MivFwt9sI
qKOXNEscRLeZZg82GWIkq56/IKWILrFS0IsWpxweWP6ra0+z5UO+u2D3JXY4Ojxi
pXHWwCS+41uTusAbYEKOZfz8wwW2/DTdZDOSfpsgbskt2z6QRpyYESdpwj2zCXpH
eGNmKdylDMXCEhYP9VyZWc8fCeWxPEgopjxgnsU7Bi0sotZKSiwb/tfV/fNMnu/V
YnkO05ESydtdjgmPE7aoCiBc2GD5d7B3hpdH50l+yaZQDAi9kJbQi5ahvfXbwyLJ
pQD+BPRslVwgN2OMqQWb77zTHX4XrCNQbfpjlalgab5WeUh4I87nvDZ4Q7qZZYL+
DM9wGQrH3osq+q+stYNHiAv41waig02rgZsBn6ytW/exfuUsWRZkiBKmL9kKgsUm
Nkor9Xjg4ApLkSb+fYDC4BhapvJwjfvOMiZ/E8hnsFqTC2VtzyktSKiG720dY155
xhxcTFw+jj4sExZXDyTmXl4hNL/wjCy+W13om7R5G1LPE5HmgEYkTkAOwcSHiB9A
FVsDuCAjjxoQPr0kTHlG9xHYGrbJBYsQRFwKiv0Q4Vt5r7bsi7QUmuTAyul7N87B
DYFpK05wgtJEK28CstMGd9U9jZAXgRsUX3QzTWg5ZOr5plRg65x1pAqVdcV+/CdG
CYYDhhtfpZ0+wrkCisA+ZIv738lw1CMmbpIT+KmvNg9BVKSzZv2m0JCqU7+p4yqd
P5DdfotaZtc9mufgoAKr8PJOyA1G95fgztWJrwiFOte4KLIRz0CzO8dkkrYTMEC7
oRB8/A4TdSjgsv52pnWOS5gncBoy965kshqvMolnAmFA2ugXg6X+e6F2YQH+Mhnf
XW//uRciMXXAvpkcI1W+MnNwCI9Urn8IJwi69Bnz/HXAkJutEo76IJlcRARFDQyI
AfQMz29pGeN2xtja5kR3S45koePwzxd1rQ2+2kkAEDTzV0wO5v87oYrrJEm81+BS
wAKctfD4kM9Qg0lfpI/aAY9gK+qqMrNgiaosxj3QorEVSqCtXXgoe4TCSIyTLX95
7xCZhNYKmswb/tG5Gz1p9behErjArOz0g0phZEqyw2FTrrYUfRn2dUqh3zlDDvnR
2Cl5hWUEYRmqgbkKaz23Q2fVZ7JFOCaIWIgKIcvWcUaDIEy/odr9DLgYuD+7EzQB
XSzwINN6RUevJYKf/zhSelMmoKX6CzmwTg1t4dyZ0LDq4Li/kezGxIey6bYS8HAM
y8vbNNlTYQE9TMmhO48FDPA6rzXrhPwXsbsmeT2+qLUUikzxPfwx05oc2xaTzMBL
9NlI/WBwtmbRpic+sx0yVXLof9cffEmPDmEMUAOf+BKE7Dl1Dxny5ciIoziQi0FU
IoNxtFFwbeXCuusb73aIm1cZxk2cNsR1qRv7IXdELZ0biwGN6VBWLPkmKE6Esy+X
3+w9b8wN1e8SkZK8Mg+CXPa7SNzzm2Cs3fX+g35+se3beylW2Qeytmun+CmmdaHP
UC2gcnRXNfvFc7fg+9vnsvEtiJHxDbiUJBVDoGeLNY9h/vnxrFFwNpqpzdUh0OLc
IGtN0vJ8BznzLcElJdw0f2h8JPruIMFmWcwCkAb6hyd/1CFqOihag1uPDsYi8SOk
EQJ6UK+eq5HNwFyJCGUAeDS+eOH8HWJiJZvcFo0/PufkwtkeRtpTebyytVdGm6Yh
lLMvTgyyg9VKwRP2TGwF4X3iCNTXcv6bjWJ5BlcZlO8ST+JU/mgIsOjYyKMWGabX
sFQsYTmAUpNX9g54wU7ggtsGfqRba+PhY7gYx3+/45mz27ur+NcrfofjKeSQ/0E/
MzB3eTteHAG0bUm+VgJN2rua1JGtSgE/K2ZAsAQ3BTesD1Lx3ezs2v8wmjYTULuS
IEvz4XFhI2bDx8HeqvGmU/xS50xdflRXfARwCctxMfHPXCP10zUDgzGY0eHqgwOE
7q26uS1aB/gwVSUa1x+qnDjWAd5fzVRHOPYqJ3G2ncWdkwWsuNf6bI9oqvGkmvkU
YwlQaW2OsltEjelDJWbXPORlbxlpuulX0vOEJKSm2x2Ql1xujI8DUhzOH65qzz+H
cwfVM5LE+HWNLxm4LOJc6NT6GsXkmLwbVUnKb6OAThJmlT9VuOQHEfVKkbYnUucW
uGprHmV6bgZovhJTBkfFpT8ziXQgjPME6iT0PM6uS+pVTM1j3NkeuaKS9K/M2LFB
uQxK0TCiaXT0q4CNuwH5QFKs255sSbRlxeAG7yCbCs3+baGztghF7jLlj8V73/0+
UgckfjhKb/nEWw4V631MHlr0oVuckahkthJuezH+5eVv0YjWXJWODFUien8f6poj
UvjBcrWLOg0+3EW3eSvYFETHm1MGqOpmkJ/HD24lEWmHBfDMBtce3NzNUNdilIP9
Q5MW6prTIq64iOOdAwmv/Tz8YwE2sZ7AlCR3y2djStkyG+iWpa9zyGrBhTOyfx4W
fcYy0v3Fmrau3ub0lTB4a1yvMD88S6k6d0HEu9XC48RZDi0Foiaf8NNqpkn5Rx4j
`pragma protect end_protected
