// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
XH2Hkk5VlH3TgzagjNKzRxIYZHvl0rAmbqBZrxdB858tA3D+sUq1CBu41xnWKkKsB6K+E3ZQK6h4
BJpAYi3g7vKuTlWs9DByigbRTy6xvXH1zL8lKUkdWJv/qAU8e4CrUDNFpC3t2RPAAnFBNARNOgyC
47smJ0vo3ntbwBxI7WLUD7tm9dvBapLvDjSDBxH5QOOZVv0y0uk61khM3kZInmbNDVnwjgzMgV8a
MC9qXatMCG+6Z2NAJ9x19kaPlQmT6A9hgqGqxt9l7C6DyuXrM/o6vuR//Ird+tZrbOWdcbTQKawx
LYZ1lR14dRULPWs9tCDvweknxxbj85QJD9IWjA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ZXCrxBjsRa3N+5Cs1dq8+m9/Ukz0cid4gqWJ0KiMVdLKUfE+8cDjeZSghlzUQtzRi/XrN6mBNJrp
lmIA29b8KrI63r0dP2jzP8bg4CMzOdothuPvICp4jMfORPqN7Eoc3YBBEe4nV+w7kW2q3mZnhlLp
TqtrcwH5k+qB1a189/+86s7LLqG9Tue+rxYJemILD+B9y9oCZNpelWXeqmIVNx2y0gyTo4bpxtVh
c9Ilk/VpF13hAgcCtBX9Fzh8h2SbLOVTSMJ5bNeZL1uh47rwfjzmDoMA11+NQ0Jei0tQKjmJL3OK
UD+bqdxURRZ1XGRGL6SVgxYFl36MJsT1R7XeP8egsqGudCsYBNLc+47RJhVhG3AyFeeqcei4wWb6
4KNaiOo2SWyZ4bkMlCaXQUgjM55gTP0FiVMMznhNocyqGaWrBeQ3eCTmbVHnkN8WrF4L0E3N49Fc
ubRhR1Czh5wwdI+bwtw/yhF8rRMrnmmX6Qc7soVIr/2Fhx7S10+s+646Ekj0W7HymrAYPIZyWL7w
U+5ncAQaBKnYmNsHoD/K+y2B6YHrYQXvZvyePZnx+exo+jhtQqaw6Mvh0q996j9lUV0xf368Sceo
b/uJbNJMfwjC/re8boOPcftipHy8kDAnWmnwSgb9FEYNfhuqYeouwevtgF/maTJnHkjPrRqpgD9+
jJg7V6OCEcP18gA2cRnGg/2Afx3u4VX/xMKanjJvBh1Db5FitTLPN58UICyqYeMMQAUa8OfcO6Ms
+xIGZDpV2x7pwZgfKcrL3MH+jF90TSKT26arMojMF4AqerAHSRGc+aHvMeWFHdVt4D4LIChi7qXX
WQ2h2kDK6oSDZWTom6ZxlMO7Wo0bM14ApG1BIGc7dyU8wuRJlzChEe1DJpzYRdesk4Wl9JUYTPkN
Ti1MDbcD0Ntyq0XYnQzoBpu3cmDWoOnuhtbCOtZ1nLdAgQdmiB20jKBGN7WLz309yuZ7rqTWlRZY
de6XEHf/levbYWW0DI5iMht8MLBcqut+c886L9i7wRWkq3f50mgFMuMoGiWJBElzBa5JC0sVQquP
BW84+Xgj5SyO/Ldx7vAI9vKFmDFPjUF72C5N5bgsKElgv23UrL8HDHhvOjmJpuJx3yI4SwFgkOXL
yO0P5/FEFdobPL7BUCX+n1YbpYmoE/peER4v/HU67y3qPLQKQLgZTfCYthvXvZQpgg9kRlUOA9Ew
yLrTOhvpQ3YzUYs+5CnrZaclBDfKXzx112Nn+cNSIktOU5bF+xRUYqsvlRZ5IuSxrOwIh3l+eEPN
V2k5FRn/MulnHRkLxOb21IXKRj9EwRyFhJojDFkEFqffklSm69yg2YMeymjhM3Z4xPIlkE8VyHf2
EVvFoSAQkx/yV9VNnI6bi/1xrq+jEEeXBvkwj/LYowrMBp3ZYsgB0e/C2dzTi2pxwQZtCrhvwCX0
MKoamY33pTZcn16+ZAIy0uC2GgwMEERPdN2aWHNKrg3QJNxwxrB5WM9KYEIe2QsUlZvww7ddyUb9
IzBXzdjv//cPi6Ir7QkmMkdnMgCd1iF5rTzZWMPDOgn60kiU3E+HvFgSjG/nJiYHiTe98utkM9Dq
rJs4kWj4CgDDnm6LwipFMEKRDKFgGqHUCX5Ux40xfp/lOG/CXW24Gf3uiAegpeeDUkgtKilJw3Vi
WKtdjh9mSYQNGtZ04uH6c8/1nQZCev7+5gwo1ezD4BM0Q/jWgEyrBsXUcJgIlNIJ3+0bKrOWKwCe
pVFBCRf3Nf9ZvUCam/HEyFbiND734izIgC2/RKI72QbJ2+VoTf5GnEXPZ+X8nbtx9CjpppEV3r9I
o9swwqf81dz+QN+vQEMYZEbiP8/LsUrgjuDDdn83dXuWilnkFs8grCTIPDXvrmrVgInDKAIc27A7
VIcOGH7LiqkejJ4wjehZsP8CZI0y4Tsw5CFptfJEJKe94so+Mz6/SXXYocfoXSuen4EjgqMMPOh4
/6YbqSeYZKkKZMyjgfFwMPZVUXWYsn8fVjwD0Qe5Ho2hAMdgAPiBvcgcRYvB6c5oq0+yJvLpXKzQ
uBLO+WLThrYmEjBaqwS8p1iaoZZf2xUnaYawwTGm2RnCYZhgNao34GyLTmXTtMaa2tKYk93p3z2a
Kuchu758Q4I/Hf3FydJPnWgzdOm65p2yka7XlQ4/hK7VMlSyrBR8wQMjg1AI4jFAxYjhgxB0kXpa
1HNGZuH9LV6ogKTOmO4rIjZeCPs5XGTYr7IGhmuXulE+8qdhlO8mVkhNUOd56tOAg+MGOH6k6c0h
j6KfhCoAibUTTeIqnfFcCjvWp55SGR35ophlvNspJkgKthOUZlAS3CZzkcD9IzGKEz/S0+gfuWpa
Bp77M/SuSXyLL+TtznixJSpqoMzmWN65NMw0QEb+3hSw5vin4Wv7L2hVBGRnRXR3eCEtkFL3Bx34
l16Ec3PlxM4XzP2Sg/sefUBkMSYtt2gh2IyYk9fshEsVl6ULPxk0Dr+zYm/HLc9uaoY3KodcoXS4
F1TJYN3rePHbTKEwSOW+jQoM5DwQZsq5p/7G+pB02VpK3xkpMRnVzJZv3UBYMMI49vYH97oqyWoE
l+iHu5XFP/ySiscVljMUQq1HxISH1qTlVMCGuSaaxCCWzfKVQcuLq2nN6ANMzYlXmJAV+AmbdEnG
eQCdgg5lG5cwqlZyKvqi4me2eBt8ha3xpo9xkoN41Un1sYI0tsVEIVVyU8vcfp0PxrSsboidB9fW
MjDqvZTrTeQMto+uT0uGWBVPuQCwVa+opCP0/yWQkhapaMS5PtWTZj1/cQdN8UKvnSwKLoTmPXeM
B0NLNaZ5o+S+j11+m+9UmU0R69nGAXlyDv18WRnrCVfBpk9Ep7PgPWZ5MymE9k6vcXnXCQg3QffB
+d3DXSzYfEoj/WXQ4fkGmSWN7oz3hzDhQA+FKMAY4UMpFjyRsAiiaijWi8YdYy7XZ8sCJ9XMMKKg
ixbQwxesU75N+R8gIjG8wBL7YRuzye/OwrsJ1IjsXYsJtYFdoMrJB7TgyeH2Qm9mgr09llQSAj9Y
Y1WapbWkROE8rlTD0A1NaLqNuojganl4jTtPi1gi52j0SS6m8956S7OaXzFuHejOYP8gJIuC8Wn6
MqYDlLhre/vTtzVu0PbPEc60ht9GTzfrsUPZM4ObRbI4ehcgK44vCQBZ9qSMLVOXccWX/3gS5+za
JOtR/FiHQqCqixaMsncJ1D8K0+wt6z+NYpHEyv/CGymZVXevPyB36Hze2yR3E2ybnF+cdUaYnE5f
YfE57iaSzGa7YZKz1SWaSjgSqBonXaXGZ5Cgfx3UiseSujabFQmZngSJdJTpJI6qenFs69bpmLOG
tnw4XKx8F4gWIt782G4RRsdPLUNjtgz8yM78LfyKiBDDrgdguuLX4HIEOPN6pgafnsW4avRp1yJs
VJiHRoihLIbB0fK64ouHzMElDu87PZowIpxEDYr+zWwCx2E6mL36tpdJl/vz9luyzZBhJK0gt20S
lXqEJOI9C4oyK+KgWsNteqfL5+AzpKvFdix55KrAPVhBQ/LP0InvWePhnvosiqeoSKfT9PTG9jsy
C6BvpAMi1FaWl6934tRpCoT1MSrzPKX6FeVAYNDUELI+xPW/bKY74tmL9RFMMC79av+/dqEBoHTT
A+Clh3Qn5+St5a+HHSbZaKYEsfnyj31QsXPh2erHD2QVFUANYoU3UwbY82u3PlyvR7ST4EFe4lvF
bQh2Rr1hM+3kOpGMfs8Wqj/F+EN51cChfV7hMhxLYZZOUX4+KNIzxQii6zRuXXifhuzEpU+H1nI2
W+kWtSbeRbv1zMN96STWuxKpGu2Y8wB/ZqVXJRwjru633W3jxRcmfs7UhdcLQMCW4+HZLcnBCv4O
t0Iccx2czN2bK9teKdERqvoRjeTytsWyKZMUQ9mShs1OG3qoqCgqksRXVO5XvACoERiXmJmTMaRJ
E5yzFVAzXonah6MyfFW0nQ7lkrZM84ff3hOpUW3P4LwTAbMLpljgfjUH0VpyDLJ5IhKNymsX0xuz
Io3fqMjYFTOJu/XzVciIXy/gGQiO70DYAhzjh8arN/xwMX87uv9d83VYzKOM3hlhzCiJapyn/SG6
45blbFASog8Dh+R3M/EIfDQMiZCt2L8h7bBPSPJTF8MsMrhDw1Ynx6swA08MdsXrvzwfsIyqCQLC
qUwGSX+JiIpO1U59rrzVHxKeaNZjHykKXDtXDuYQ+npN7LUlgaYGlwXd9cQNBgy0wR6edzp9HIGb
ixpSAv+bsFsUzb+7z+/0PIbqlPWwDEDXzZQB6iyCShF7p3IrwB57VInVdUVzlMzjOcjMH+2Lv4nw
IAQamDMyzhcJNsU8reaVX4PubXUJLb4Do8SqB+Ft2nzfqqENgZCZ6lCsDhRYzg8BSeWrMKrQYk35
YnLxPpxy3N+dCzlec/uC2Xfv/vwJQzUH0mjDCBOLjCMpFRQi0stGDqNW+U6m9QKk4C78ugyIk5cM
J/ueLBa4/lEE6R3BLzzNREdXTEZDR/i1iIxMBy5rXqosne/BRWlxqJ9m7NKzSw7qCKx7OWVgr0ki
N/nC5Qt9ojl3lpDGfRL3Tyfl+BdezOi0MsdTdY9FXeAovLMuttuYgdsTEGbCNNvBI98Dfli+rp3T
1a9qrDYCxlYHM8Nh8Ue4RmnSxtEhGsr2V/88yrPBhmm691AqZlmebgTZbL52voopJrvztF0gree0
1dxFh2XZptku/VabAMM3bKX/p4/826pb80vw8BM3ztaOc8+XTXuektSoy0GstI+U5mrZ098So5Cc
uaFq4c8yGcf6mlu0e41QmNAI5foEY0jcKhCmuMHfMG/V4Ud7DKiriejt3UHM5L3gxpMfE7OIGXAT
B9QEUmZV+QLeikJM6Zzy51JwP2CRdm/k6xA43NCHt9r4czfmN8l57uRbLpSy8Z3Q9bsn5WVCiFEM
c3NfXcKt2zppIIDZe55VtnJMFzW+cFAkoyCw8X3IipyMU6sSI17rfaJOKUuNagu/KAyWsoE0x2Bw
VWADL0OKpQsv+NeMGQUGsaF+L1ndlf0IU6vHwInwv5Ol9ZsUdoiOlG6QwkrO56vLEJZ/03zE6NOa
vDef2fvUkpSzEg1ewv4JqWrXFK2UbGO88hqp+CIjFIUGyVnddGpXT8QqYdko3oEcSF5mtICjiq1n
6MwzU8dUvcPygRGVU29qdqfr22XxxnQjQmgxOLGj7mo+yMkzzkzOipLhMaZryS1sRLHlKEqaYVsY
2jW0sguHLEDls0x8GJHqYX3CvQNgdtYHM1Kgkr4JujgXsFAYnQU+v9gCCeSkX5mEGgtRqP7dBRie
eK1B8mtFd/l6RRxA/61lOTdNY/fuExmzLW3tvKW++3KPuCHhuX+Zwnw4NtIYWr8kGU+w4/de5nKA
d+1EcJRptlJtfIF035zgp3TyeW1M5DmYxyPiPGxyJetPYwL0N0Wu3nmrDc2llldta7iiItxiWqO9
s0C/wwubliSnUACsGTXwbVUPO2jFWFwUXKo1rs9JjVVCITIjqENAqVJwIoLLpl+yqtDyzYvx2hux
tXP7VrCG+R1lTf+3cyWryDEn2dc8tAupGBtvlIcAVk6tblVZGZSsV2PoPsr33FZ0Rcgu3n45ZAPD
tKSqVJpDn8BIxYsnD6oioKbpr9SrGuLdc7skYDiiCPhBUww4aAwkdh6BZBKmIj7rEol32QOl0hcR
gPlA0OfQxj8A7fGkQ+xKX9tcd17tuCYVI1xI+yGJyzuz7YDdvQl++rCmoVDJUjINV+Nao7n4D6k4
WcfvUnbiefMX0SylCHEXa9HISSe4YKWAm7uBsSc4XboWBaokk1wOxxezG6altrzMWn8yB2biGLYS
I4m3P6zdyyxR9jB6k1dml9oVv9rLlWqg23ZjmAfjykWNmIzM1Wr7iAVfocNBwwAZXTn9a0e9Wm+1
IQthX5Eu0Xg1Bs2oe0zXnAUwCGkv23JAv1flLqVGC5B6U2gDLX9XZiGdZiOUgiAcIZW48YFP8wMG
cAOq2UvsBxFF57REeOF+H4v3lpH6S3SDP/Rmj9FAuYq7WK3r+mSGU6lisA4DLpWlu7qt/2Ysbe72
EHGLYTMf+AzzdhyZ24n0rHTKx8inqvG/RjqSe+VrfNskF0C0/NwvT2HJceIyXl8yXpc3BmGahjSy
FfoAzBHSbBb4oLJc4VLFD8aE4c7qaFaZZPoCBdk8l4CSsY+Bv00mIO9QMQ+LOg754h88CAMqmLgd
zuzNQEldrT+fbaJm9+zGvbTg5nWMm5B1PFNHQdBz+S1UZvVYiH1khmXnQXOoiciigiyVLwKW8qL+
Q90BuYPuQvs4oZ7RUUfBzklKWSueHfp3v/uK1taSfYDMkUvAZZH3IsYUhxpgwX6DDMjCRm0Y8J9b
p5uG/ghK78mMkyuDB1AGlpOJqZkuKRpHo8gAVQf/hYDKlTENl8BGVhf7MrAdes/ElbrHfMMgId5m
67+KI7IcjjampwfwEEq0shrYTdWRljUf2DvoOIP0JBdgazFocO54YO6YqvSSsiz9WnNxf6yAZ4S5
SvQQlYxzB4azYfUrb/zju2WqZfBiCbTqaIiSSFfpQ2RG6X2j7C+e9qyn+HZ4XSADrWsT6muElGMs
/sZpmNL0YCMiZ9O6jvfn4gi58eonsIdImd70dbYojZPkx4IgI/rWoQ674s2O28nYR/xTHX313Gjm
4iGZVsrRvx0AtxOMWBrCOH+6oogvnxD7pOINgW9dqtmik0CMjyhsGy/2rjVjpn+iKZ6eyWI7HWNW
mSnxC/drYhJhLNgEg4qAFUvZF/QOn9GrWpB/P/fKUlpmXbhH0uWsVNuZvYIipphXahOBOx1WSCkb
sJ8jb9HnXTDwsRVOT7HU3QGS1XLNVLz9Sdg6Z1luoEk2aeDn9R6uprrvKZmSGm+1IgGnzQ9Y1Pba
LEdmWncsCpmCYv3wtMXF8z4m0GjZphx0lIctqAuQvt3ptCT0RUWQ++XPxRYZoZtUJlbcDWgedEuz
/4mf7rwMRfwGYqHVL1fjVdz0v8vKF7hf4z2XDp4gngcjBGuqpFDv4YQE0YEHbaBaRci4dFy58Mj3
pqXQaqQW3aMJPlJJDnrB6HBExA2Uikf2BdTBwu6LB09ObHbCVkzJSc+NEJxB9l2CJeod1PM3WncA
t5OK0AngkN77iG9gAnLHYtWEsaggIvc6uSuBSZYS99/mWyHbucQ1vmvg2y3821/W5bi2LqEtBY7h
B7WiJUujaKycaQp2QPjfCkri0S+wnm4q3YoP2ZlH4qp19c2Lxzv/Oe6KzZsJD4cpOhfYFua6sGSm
CmZj2BM1ISatDQZEredC2VbxYB5/Y86LIaMjjGy4v0AtK7z0xbWo6Kp+fuXF8qHKDoVA+PP9URS0
fFSkuKZP3PvVeoCrpij/fxBH2PWykD3W1VDjCz+eTRvzodEBE58NebDxGOyVE/XjvlQ3vTeYmiOr
onWhxzUVsy/k2U6Jhf5iyZjjU3X8Nwk5kY6mOmxBGOvTlgmcirnCzqrLSkTpYpq+ikieAKJGDYgy
CzbjOYRx/D4nllOlW1+pqWzbygDs6IfdvlU0JD/VFXGuT8C/Xp+z++0OB+vgRYjPtCj4kbVHasiH
1TBNblMQDZDVdxk+8HWo0peuJCzjBFmw6kRNikn4cUnrGLSJVKaXSP/aDAEOv+sXtjwhHAa1Y3zs
LEBgr56T8o6B86dQB3e6jEkqn6xIJr4e0NM8tOdTA492bsSuzyPVIKdHrXrjO3dErnCqHuWpsszu
85EVsMF8aNGo2VbOrt+7FwFFOOs2FZ1I+uJARrCoUGyiai41EYBsjm4EN0BX2LuUY8eYFthXz4Jj
MeYxHnV4LrnQepmOdR85Kz6ehm2WSPyoPCrzzUlOlI6hWWthq+UzMQUNJCp1rf2o6eELmCFRoSHZ
3jDCKCtKsSCzrMojV3V/oUskNOSGPRMA85m5RbAaR677n130nbCVt1Z7vETxizSPZuRuAqj5e1pW
wjCT2+nGZa6tujvdiso2jXKzzAkq2ygQmR3l+tsAhiSIXVgV6qywcWv51KHBTpmH/oNoh6HPPwil
U8+fmd+E2R4pa13JcKLpgg4myXGIv2ELQTfUplzSmj8DJRf6RhBKXiQyuQVoRXxT9xpxxi01tWrm
oKWA2Ed4VNrGZBNt7+o7M+Tzq7lQr62CZiQC13EByiUBh14+HANntkVIvBtKoIxgB93vjQi3S18u
gu/lvOHVcCJMloTYOe4Ndnn/tg+0XAWxlAqGRhlW6lvVU3LUXL99Zg0rCtHc50yCkPZOvqRJvzub
GmAHO/t92YQm1W16D/EzwEcKlQHe87ZVN1mQDA7LsIM6BJLoqr9oFGDeGFWWsOyBlS7a+KHJQdQS
VHEexQwrG++dOCjweW1B+TdyBqkrbk6hYzgaCHpvZy/sIQVqXcuIRLdOJwawSfMYTEfb//Ml33JA
9oZtCZzgysk/Ma7RWazoF+ih7T6DjaOwHLn9Z6FOjeI9jLGdRI2nGhn79OvvaKB9SzNKGQBHDH1V
zP1pPl3+Haa+miAwZaKJv6Mtd+ahw0f+kynw2jKymjd+gpSse24bJywnaoi0LdAtLKxJrWxmclOz
dW5dRl0elQoMHWCNZTCwHhAk9F+nAlwr8kjBX2EEQCN3yO5NvE3mzdzTb+G/LLlw+Rax6j2QWSo1
soKEeQBSBxYBQOgRtuuH+zGhcTXj2IbyNU/HZLibcI9+39Ziid0ghlFETVjTVM3z9uUpjiiEvse8
OXX7uIgs8J00sQYRUm3CDo/SNWtiQF/bhJNtNFFF49Gv1rslhp1ynVHllt6NNmzyQGX8ihJlulSJ
i11cU5jTAh1PwMpv+E0wrdRGrhWWuqU0g+rT7IxuhpeFyxZsJwgoxlq5DLmKFMJEOJXZHfhvIo9o
XIAx7m+exYEEFT/t1nSz9YZE1uCn6RwNQYYoPFMCs/t12WjWK1/7PatcVbAEHP4mCAJPj5Y0lByM
5m6ltmT0JOc5pPzPpwncpaKWO2i20XqhzUhKSBKgrX8qU8GOgqs+V+bL3QdwDb5rU3gCil5zQYBS
MQ==
`pragma protect end_protected
