// alt_xcvr_reconfig_cpu.v

// Generated using ACDS version 13.0 124 at 2013.02.06.18:11:40

`timescale 1 ps / 1 ps
module alt_xcvr_reconfig_cpu (
		input  wire        clk_clk,                        //                    clk.clk
		input  wire        reset_reset_n,                  //                  reset.reset_n
		output wire [9:0]  reconfig_mem_mem_address,       //       reconfig_mem_mem.address
		output wire        reconfig_mem_mem_read,          //                       .read
		input  wire [31:0] reconfig_mem_mem_readdata,      //                       .readdata
		output wire        reconfig_mem_mem_write,         //                       .write
		output wire [31:0] reconfig_mem_mem_writedata,     //                       .writedata
		output wire [3:0]  reconfig_mem_mem_byteenable,    //                       .byteenable
		output wire        reconfig_mem_reset_reset,       //     reconfig_mem_reset.reset
		output wire        reconfig_ctrl_reset_reset,      //    reconfig_ctrl_reset.reset
		output wire [4:0]  reconfig_ctrl_ctrl_address,     //     reconfig_ctrl_ctrl.address
		output wire        reconfig_ctrl_ctrl_read,        //                       .read
		input  wire [31:0] reconfig_ctrl_ctrl_readdata,    //                       .readdata
		output wire        reconfig_ctrl_ctrl_write,       //                       .write
		output wire [31:0] reconfig_ctrl_ctrl_writedata,   //                       .writedata
		input  wire        reconfig_ctrl_ctrl_waitrequest, //                       .waitrequest
		input  wire        reconfig_ctrl_ctrl_irq_irq      // reconfig_ctrl_ctrl_irq.irq
	);

	wire         reconfig_cpu_data_master_waitrequest;                                                        // reconfig_cpu_data_master_translator:av_waitrequest -> reconfig_cpu:d_waitrequest
	wire  [31:0] reconfig_cpu_data_master_writedata;                                                          // reconfig_cpu:d_writedata -> reconfig_cpu_data_master_translator:av_writedata
	wire  [13:0] reconfig_cpu_data_master_address;                                                            // reconfig_cpu:d_address -> reconfig_cpu_data_master_translator:av_address
	wire         reconfig_cpu_data_master_write;                                                              // reconfig_cpu:d_write -> reconfig_cpu_data_master_translator:av_write
	wire         reconfig_cpu_data_master_read;                                                               // reconfig_cpu:d_read -> reconfig_cpu_data_master_translator:av_read
	wire  [31:0] reconfig_cpu_data_master_readdata;                                                           // reconfig_cpu_data_master_translator:av_readdata -> reconfig_cpu:d_readdata
	wire   [3:0] reconfig_cpu_data_master_byteenable;                                                         // reconfig_cpu:d_byteenable -> reconfig_cpu_data_master_translator:av_byteenable
	wire         reconfig_cpu_instruction_master_waitrequest;                                                 // reconfig_cpu_instruction_master_translator:av_waitrequest -> reconfig_cpu:i_waitrequest
	wire  [11:0] reconfig_cpu_instruction_master_address;                                                     // reconfig_cpu:i_address -> reconfig_cpu_instruction_master_translator:av_address
	wire         reconfig_cpu_instruction_master_read;                                                        // reconfig_cpu:i_read -> reconfig_cpu_instruction_master_translator:av_read
	wire  [31:0] reconfig_cpu_instruction_master_readdata;                                                    // reconfig_cpu_instruction_master_translator:av_readdata -> reconfig_cpu:i_readdata
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_waitrequest;                   // reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> reconfig_cpu_data_master_translator:uav_waitrequest
	wire   [2:0] reconfig_cpu_data_master_translator_avalon_universal_master_0_burstcount;                    // reconfig_cpu_data_master_translator:uav_burstcount -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] reconfig_cpu_data_master_translator_avalon_universal_master_0_writedata;                     // reconfig_cpu_data_master_translator:uav_writedata -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] reconfig_cpu_data_master_translator_avalon_universal_master_0_address;                       // reconfig_cpu_data_master_translator:uav_address -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_lock;                          // reconfig_cpu_data_master_translator:uav_lock -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_write;                         // reconfig_cpu_data_master_translator:uav_write -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_read;                          // reconfig_cpu_data_master_translator:uav_read -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] reconfig_cpu_data_master_translator_avalon_universal_master_0_readdata;                      // reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> reconfig_cpu_data_master_translator:uav_readdata
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_debugaccess;                   // reconfig_cpu_data_master_translator:uav_debugaccess -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] reconfig_cpu_data_master_translator_avalon_universal_master_0_byteenable;                    // reconfig_cpu_data_master_translator:uav_byteenable -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                 // reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> reconfig_cpu_data_master_translator:uav_readdatavalid
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;            // reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> reconfig_cpu_instruction_master_translator:uav_waitrequest
	wire   [2:0] reconfig_cpu_instruction_master_translator_avalon_universal_master_0_burstcount;             // reconfig_cpu_instruction_master_translator:uav_burstcount -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] reconfig_cpu_instruction_master_translator_avalon_universal_master_0_writedata;              // reconfig_cpu_instruction_master_translator:uav_writedata -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] reconfig_cpu_instruction_master_translator_avalon_universal_master_0_address;                // reconfig_cpu_instruction_master_translator:uav_address -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_lock;                   // reconfig_cpu_instruction_master_translator:uav_lock -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_write;                  // reconfig_cpu_instruction_master_translator:uav_write -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_read;                   // reconfig_cpu_instruction_master_translator:uav_read -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] reconfig_cpu_instruction_master_translator_avalon_universal_master_0_readdata;               // reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> reconfig_cpu_instruction_master_translator:uav_readdata
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;            // reconfig_cpu_instruction_master_translator:uav_debugaccess -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] reconfig_cpu_instruction_master_translator_avalon_universal_master_0_byteenable;             // reconfig_cpu_instruction_master_translator:uav_byteenable -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;          // reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> reconfig_cpu_instruction_master_translator:uav_readdatavalid
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // reconfig_mem_mem_translator:uav_waitrequest -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_burstcount -> reconfig_mem_mem_translator:uav_burstcount
	wire  [31:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_writedata;                     // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_writedata -> reconfig_mem_mem_translator:uav_writedata
	wire  [13:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_address;                       // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_address -> reconfig_mem_mem_translator:uav_address
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_write;                         // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_write -> reconfig_mem_mem_translator:uav_write
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_lock;                          // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_lock -> reconfig_mem_mem_translator:uav_lock
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_read;                          // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_read -> reconfig_mem_mem_translator:uav_read
	wire  [31:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_readdata;                      // reconfig_mem_mem_translator:uav_readdata -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // reconfig_mem_mem_translator:uav_readdatavalid -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_debugaccess -> reconfig_mem_mem_translator:uav_debugaccess
	wire   [3:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:m0_byteenable -> reconfig_mem_mem_translator:uav_byteenable
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_source_valid -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_data;                   // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_source_data -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rf_sink_ready -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // reconfig_ctrl_ctrl_translator:uav_waitrequest -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> reconfig_ctrl_ctrl_translator:uav_burstcount
	wire  [31:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                   // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> reconfig_ctrl_ctrl_translator:uav_writedata
	wire  [13:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                     // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> reconfig_ctrl_ctrl_translator:uav_address
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                       // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> reconfig_ctrl_ctrl_translator:uav_write
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                        // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> reconfig_ctrl_ctrl_translator:uav_lock
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                        // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> reconfig_ctrl_ctrl_translator:uav_read
	wire  [31:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                    // reconfig_ctrl_ctrl_translator:uav_readdata -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // reconfig_ctrl_ctrl_translator:uav_readdatavalid -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> reconfig_ctrl_ctrl_translator:uav_debugaccess
	wire   [3:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> reconfig_ctrl_ctrl_translator:uav_byteenable
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;                // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;                 // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;                // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;          // reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                // reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;        // reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [82:0] reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                 // reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                // addr_router:sink_ready -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;   // reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;         // reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket; // reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [82:0] reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;          // reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;         // addr_router_001:sink_ready -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_valid;                         // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [82:0] reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_data;                          // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router:sink_ready -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:rp_ready
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                       // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [82:0] reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                        // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_001:sink_ready -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                             // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                   // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                           // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [82:0] cmd_xbar_demux_src0_data;                                                                    // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [1:0] cmd_xbar_demux_src0_channel;                                                                 // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                   // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                             // cmd_xbar_demux:src1_endofpacket -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                   // cmd_xbar_demux:src1_valid -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                           // cmd_xbar_demux:src1_startofpacket -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src1_data;                                                                    // cmd_xbar_demux:src1_data -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_demux_src1_channel;                                                                 // cmd_xbar_demux:src1_channel -> reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                         // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                               // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                       // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [82:0] cmd_xbar_demux_001_src0_data;                                                                // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [1:0] cmd_xbar_demux_001_src0_channel;                                                             // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                               // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                             // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                   // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                           // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [82:0] rsp_xbar_demux_src0_data;                                                                    // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [1:0] rsp_xbar_demux_src0_channel;                                                                 // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                   // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                             // rsp_xbar_demux:src1_endofpacket -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                   // rsp_xbar_demux:src1_valid -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                           // rsp_xbar_demux:src1_startofpacket -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [82:0] rsp_xbar_demux_src1_data;                                                                    // rsp_xbar_demux:src1_data -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_demux_src1_channel;                                                                 // rsp_xbar_demux:src1_channel -> reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                         // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                               // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                       // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [82:0] rsp_xbar_demux_001_src0_data;                                                                // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [1:0] rsp_xbar_demux_001_src0_channel;                                                             // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                               // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         addr_router_src_endofpacket;                                                                 // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                       // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                               // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [82:0] addr_router_src_data;                                                                        // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [1:0] addr_router_src_channel;                                                                     // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                       // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                // rsp_xbar_mux:src_endofpacket -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                      // rsp_xbar_mux:src_valid -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                              // rsp_xbar_mux:src_startofpacket -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [82:0] rsp_xbar_mux_src_data;                                                                       // rsp_xbar_mux:src_data -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_mux_src_channel;                                                                    // rsp_xbar_mux:src_channel -> reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                      // reconfig_cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                             // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                   // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                           // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [82:0] addr_router_001_src_data;                                                                    // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [1:0] addr_router_001_src_channel;                                                                 // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                   // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_demux_src1_ready;                                                                   // reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src1_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                // cmd_xbar_mux:src_endofpacket -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                      // cmd_xbar_mux:src_valid -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                              // cmd_xbar_mux:src_startofpacket -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_mux_src_data;                                                                       // cmd_xbar_mux:src_data -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_mux_src_channel;                                                                    // cmd_xbar_mux:src_channel -> reconfig_mem_mem_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                      // reconfig_mem_mem_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                   // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                         // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                 // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [82:0] id_router_src_data;                                                                          // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [1:0] id_router_src_channel;                                                                       // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                         // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                                   // reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                               // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                     // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                             // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [82:0] id_router_001_src_data;                                                                      // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [1:0] id_router_001_src_channel;                                                                   // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                     // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire  [31:0] reconfig_cpu_d_irq_irq;                                                                      // irq_mapper:sender_irq -> reconfig_cpu:d_irq

	alt_xcvr_reconfig_cpu_reconfig_cpu reconfig_cpu (
		.clk           (clk_clk),                                     //                       clk.clk
		.reset_n       (~reconfig_ctrl_reset_reset),                  //                   reset_n.reset_n
		.d_address     (reconfig_cpu_data_master_address),            //               data_master.address
		.d_byteenable  (reconfig_cpu_data_master_byteenable),         //                          .byteenable
		.d_read        (reconfig_cpu_data_master_read),               //                          .read
		.d_readdata    (reconfig_cpu_data_master_readdata),           //                          .readdata
		.d_waitrequest (reconfig_cpu_data_master_waitrequest),        //                          .waitrequest
		.d_write       (reconfig_cpu_data_master_write),              //                          .write
		.d_writedata   (reconfig_cpu_data_master_writedata),          //                          .writedata
		.i_address     (reconfig_cpu_instruction_master_address),     //        instruction_master.address
		.i_read        (reconfig_cpu_instruction_master_read),        //                          .read
		.i_readdata    (reconfig_cpu_instruction_master_readdata),    //                          .readdata
		.i_waitrequest (reconfig_cpu_instruction_master_waitrequest), //                          .waitrequest
		.d_irq         (reconfig_cpu_d_irq_irq),                      //                     d_irq.irq
		.no_ci_readra  ()                                             // custom_instruction_master.readra
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) reconfig_cpu_data_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (reconfig_ctrl_reset_reset),                                                   //                     reset.reset
		.uav_address              (reconfig_cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (reconfig_cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (reconfig_cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (reconfig_cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (reconfig_cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (reconfig_cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (reconfig_cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (reconfig_cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (reconfig_cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (reconfig_cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (reconfig_cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (reconfig_cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (reconfig_cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (reconfig_cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (reconfig_cpu_data_master_read),                                               //                          .read
		.av_readdata              (reconfig_cpu_data_master_readdata),                                           //                          .readdata
		.av_write                 (reconfig_cpu_data_master_write),                                              //                          .write
		.av_writedata             (reconfig_cpu_data_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (12),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) reconfig_cpu_instruction_master_translator (
		.clk                      (clk_clk),                                                                            //                       clk.clk
		.reset                    (reconfig_ctrl_reset_reset),                                                          //                     reset.reset
		.uav_address              (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (reconfig_cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (reconfig_cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (reconfig_cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (reconfig_cpu_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                               //               (terminated)
		.av_byteenable            (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                                               //               (terminated)
		.av_readdatavalid         (),                                                                                   //               (terminated)
		.av_write                 (1'b0),                                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                                               //               (terminated)
		.uav_clken                (),                                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                                               //               (terminated)
		.uav_response             (2'b00),                                                                              //               (terminated)
		.av_response              (),                                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) reconfig_mem_mem_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (reconfig_ctrl_reset_reset),                                                   //                    reset.reset
		.uav_address              (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (reconfig_mem_mem_address),                                                    //      avalon_anti_slave_0.address
		.av_write                 (reconfig_mem_mem_write),                                                      //                         .write
		.av_read                  (reconfig_mem_mem_read),                                                       //                         .read
		.av_readdata              (reconfig_mem_mem_readdata),                                                   //                         .readdata
		.av_writedata             (reconfig_mem_mem_writedata),                                                  //                         .writedata
		.av_byteenable            (reconfig_mem_mem_byteenable),                                                 //                         .byteenable
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_chipselect            (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) reconfig_ctrl_ctrl_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (reconfig_ctrl_reset_reset),                                                     //                    reset.reset
		.uav_address              (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (reconfig_ctrl_ctrl_address),                                                    //      avalon_anti_slave_0.address
		.av_write                 (reconfig_ctrl_ctrl_write),                                                      //                         .write
		.av_read                  (reconfig_ctrl_ctrl_read),                                                       //                         .read
		.av_readdata              (reconfig_ctrl_ctrl_readdata),                                                   //                         .readdata
		.av_writedata             (reconfig_ctrl_ctrl_writedata),                                                  //                         .writedata
		.av_waitrequest           (reconfig_ctrl_ctrl_waitrequest),                                                //                         .waitrequest
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (71),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (72),
		.PKT_THREAD_ID_H           (73),
		.PKT_THREAD_ID_L           (73),
		.PKT_CACHE_H               (80),
		.PKT_CACHE_L               (77),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000),
		.SECURE_ACCESS_BIT         (1'b1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) reconfig_cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (reconfig_ctrl_reset_reset),                                                            // clk_reset.reset
		.av_address              (reconfig_cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (reconfig_cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (reconfig_cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (reconfig_cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (reconfig_cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (reconfig_cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (reconfig_cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (reconfig_cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (reconfig_cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (reconfig_cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (reconfig_cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                               //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                             //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                         //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                               //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (71),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (72),
		.PKT_THREAD_ID_H           (73),
		.PKT_THREAD_ID_L           (73),
		.PKT_CACHE_H               (80),
		.PKT_CACHE_L               (77),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000),
		.SECURE_ACCESS_BIT         (1'b1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                     //       clk.clk
		.reset                   (reconfig_ctrl_reset_reset),                                                                   // clk_reset.reset
		.av_address              (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src1_valid),                                                                   //        rp.valid
		.rp_data                 (rsp_xbar_demux_src1_data),                                                                    //          .data
		.rp_channel              (rsp_xbar_demux_src1_channel),                                                                 //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src1_startofpacket),                                                           //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src1_endofpacket),                                                             //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src1_ready),                                                                   //          .ready
		.av_response             (),                                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (71),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (72),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) reconfig_mem_mem_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (reconfig_ctrl_reset_reset),                                                             //       clk_reset.reset
		.m0_address              (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                              //                .channel
		.rf_sink_ready           (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (reconfig_ctrl_reset_reset),                                                             // clk_reset.reset
		.in_data           (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (71),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (72),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (reconfig_ctrl_reset_reset),                                                               //       clk_reset.reset
		.m0_address              (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                             //                .channel
		.rf_sink_ready           (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (reconfig_ctrl_reset_reset),                                                               // clk_reset.reset
		.in_data           (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	alt_xcvr_reconfig_cpu_addr_router addr_router (
		.sink_ready         (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (reconfig_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (reconfig_ctrl_reset_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_addr_router_001 addr_router_001 (
		.sink_ready         (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (reconfig_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                     //       clk.clk
		.reset              (reconfig_ctrl_reset_reset),                                                                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                              //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_id_router id_router (
		.sink_ready         (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (reconfig_mem_mem_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (reconfig_ctrl_reset_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                         //       src.ready
		.src_valid          (id_router_src_valid),                                                         //          .valid
		.src_data           (id_router_src_data),                                                          //          .data
		.src_channel        (id_router_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                    //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_id_router_001 id_router_001 (
		.sink_ready         (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (reconfig_ctrl_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (reconfig_ctrl_reset_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                       //       src.ready
		.src_valid          (id_router_001_src_valid),                                                       //          .valid
		.src_data           (id_router_001_src_data),                                                        //          .data
		.src_channel        (id_router_001_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                  //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),            // reset_in0.reset
		.clk        (clk_clk),                   //       clk.clk
		.reset_out  (reconfig_ctrl_reset_reset), // reset_out.reset
		.reset_in1  (1'b0),                      // (terminated)
		.reset_in2  (1'b0),                      // (terminated)
		.reset_in3  (1'b0),                      // (terminated)
		.reset_in4  (1'b0),                      // (terminated)
		.reset_in5  (1'b0),                      // (terminated)
		.reset_in6  (1'b0),                      // (terminated)
		.reset_in7  (1'b0),                      // (terminated)
		.reset_in8  (1'b0),                      // (terminated)
		.reset_in9  (1'b0),                      // (terminated)
		.reset_in10 (1'b0),                      // (terminated)
		.reset_in11 (1'b0),                      // (terminated)
		.reset_in12 (1'b0),                      // (terminated)
		.reset_in13 (1'b0),                      // (terminated)
		.reset_in14 (1'b0),                      // (terminated)
		.reset_in15 (1'b0)                       // (terminated)
	);

	alt_xcvr_reconfig_cpu_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (reconfig_ctrl_reset_reset),         // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (reconfig_ctrl_reset_reset),             // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (reconfig_ctrl_reset_reset),             // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_cmd_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (reconfig_ctrl_reset_reset),         // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_cmd_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (reconfig_ctrl_reset_reset),             // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (reconfig_ctrl_reset_reset),             // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	alt_xcvr_reconfig_cpu_irq_mapper irq_mapper (
		.clk           (clk_clk),                    //       clk.clk
		.reset         (reconfig_ctrl_reset_reset),  // clk_reset.reset
		.receiver0_irq (reconfig_ctrl_ctrl_irq_irq), // receiver0.irq
		.sender_irq    (reconfig_cpu_d_irq_irq)      //    sender.irq
	);

	assign reconfig_mem_reset_reset = reconfig_ctrl_reset_reset;

endmodule
