// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JtQXVPvW/CX/H10TTjF6cVfpNxpSafA5ws9nwqdmKPnWE87e/ug/MXUwkXDLQifw
yGhilamZoxN9Mclt1ktmqTdOzAEuSmQwJV8p1RmAme50wSyZyT/3mZgpL4RwPCCT
q69Q5qz9aNOZhgHN6eJn/URdNzIPCCjfrte24/vuZus=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10240)
Vel76jlWrKUslu7RPQ0EnI4LPkw4X3eCrwN8/XRUWdXjRZV4kU38pY8cHWb2qUdj
qiHrj4XV0UxPhTLyE99/ppsUpaishETHRENghsPgrf1FPjvjxoJ3B+dkNW95wIX0
CTfzx3aayLDQEVmWWc5r48aSgcjHgRXDBIWXdeYVvqC4QY7ZgQv2OuxUaZXKcjY+
ftocxWYbCq1KEB3Cox9xW4R8zHgrMAvMjNPp7rOopfy6rsyXlzw2RUNBXqDPKHsy
d/X69ZPQDySd9zMVoEKSBc6KFOwJSsGVmdY0spb4nr3O2KyH4OWxRQ9iVZLJKqFh
oYvOhkGIhRJDe9g1CeYJes6GP43DuedyWVn+bKwXozykaLqjkBDdo2aAqlAg8oVZ
H1RQBrd2CtSleuKaueLYPIailQgO7v1AQVUbkyy//cLpGxVJGTzC+Hssvy1GtLDK
BrB7Nv44ZmZMiJXc68cDoKIrziKLNfsIDfYVVTdob4kX21MifdjcPaVKuSUvtwFG
dfdPzw3AbTqh8Ns8jtwwmGWcMJtQjEBLsxJu9F3pTvcQ/hsHgBkZk200XwDxWqH8
mUw9UNfF8SeIj6xyxd2EdDyj6g06ZCng3Bw0eCJQkPBiVG2HujwjlHnSIvUG2hwG
I/Bh2mgO2rd+20IxNN4ejRiHZ28e1nkpTEl6ersb5+wSGoWkmr/6TvXZHYedHjI5
LL0R3LD3CUr8qViqgu9M1a62JLZxQkJUlcd5ztkrwythJMfL0C7G5fctNFtSVT6/
Y7MaSi+dz3f23VoFIjXDCggZOzcXEYLQOYN8LOLnw2NXAvWH78NRmSnw3F068aVh
SheamdjcCyD0Kxp8ygKWOi8XzfYNxTfh5opNP8bTHVvIhRm2/cnuRXoKhFwWPPLH
RALydmIJCISkGJ9C/OfESyQ9qe+mKNMpWqBhDiKByE95fCOSnkn1U5b2hocj4Zmz
PI34zX+2PDqwUarziV2rhKVnIvUnvIsgM6RGv+Ps1Cia0M1ShX+KDGhgONJr9sXM
rf9C/qoyWaKLrZOGPgm3FSbao2HUEWVNatt5GTLR+LkykQYu3Zr1/JYhJpDmVN1I
isXFxGJWnJJfIRo4m9W6EW+hmzBNn7WTx5W+lE8NnxDNB0n1oJwqI0bdzf1G/u65
MzfQyxJ+d5eBVD7WtmEAe6dJ2ADKCAMOf/uH65DjbNxJO5OWmRB1NMNMZn4a2lu0
wlr15xL7ATAOg2GFwcWvHO+pwy79/16f3wn0CPtM/NgBzOEmlsUxt+Xwem2j872j
PvjdKin7okX4M1R6o74P8CS72JDyODhgnv0qQxPQd7n1Xz38FHdIU3fqrRJnNyRh
XfIby3F3gwZ0hALo8xENykHeZT/jclbw6MXxdXiuduLuLvDkHineewQrqLIN9VNw
jvQ7OJmOiBvXFTGuV+cpdmFe5BxbiQ3ULI0mek0OFAz44iO0Mzz+9PsbyqjGjiPm
+Jt/p5ECHSHRcFTute4t1ibGKWDm3iVdd+0jmjd24KYc51rRUXyWrZcIyrazy4xk
f91mNEe81nmhqXC3dH0EUHUm77pLNYo/xVoDWeDei3dytKKaCnnn0IC5MptKFcUf
MTU+o2PbZwMpC9kazOvVXRu4bIVJ3EZ6RBD70KS8OJzUmpXptPSVHPFvnXMmLUyV
Gok7+WBuJaP/QyZeV9WNF09KfVAzhPuGAEdLPQZVn1zURILj/hYYJw2pvGkaPuun
TS17+DpE3rsBfiH/IS83CqeE9Onvvgo0DWxW0hrTl/+YWqTvdoR7mPr9PHqXYARZ
oEje2AY7COcRvYvAN4NP37XOrdAXBf9sh1kCw89GsAVNqzJf0S/u+RfozJfa6PT8
QHEpf9TW6KpZiXFPPZdV9A+j9f48gAvPPOEiG+SckHz4GpKG9FnDi/TNnBKFQoCD
MkkuxuW9f2WK/P2lv932+rNLvB1AOn0az3s6AM2b3ggK0HGDqEgC6TpZJPBoXCsI
YFI3a1lULIfbyhQKBNRruvAXPyCcBR2SCT2hSRG5ZKbNZCm8DhcgNe5zCZNSKEGY
mwzUzgVqrQJElZkq8tW4m5v+wAfc2DPHR7VsC1urPttrhfzybxZMDtw2XSyWNztx
kmnOlSa+oPl3/A+JQTiADiTOiieCdsqpGcDXtaO3GSuQGbGc+E8ROt2brqboSe+I
dCod6k3w1aLmGTg6ruvx/UoNaElEggPm6LDMbMEv7+kBdDcGuapsDAptckWQBoFX
7unKYLT0q9BYfrOsgQkYqW4z9EQLIvO6dg1qRcw3GQxqJBjNmXDfRA1hOwYaf3tk
g9Mg5ZMGovcX0RXovQJz9JwkeXg+aohUuSg5tbRc7w8/Nse7pNRvjG1UAlwkOld9
onAEgXrH6g3+o66r2IYYWkdW5qbfH/z1z9Gtrs5nStPxJc+Oy7GgCLA1l0mj2IL7
xE8uDSBd+/yviG0GGJDCGFthXcs04GSbLggjKodLx8xnVov3Nirj4ZKZFfhrJ1I0
XrzrlDYZsM3CKaoT8i+JOt70gKL+qOaNacJWqb0R5T8dWchCZ0wFWZYBEK11Aj8+
/wld3nN34a1pgTqIF3uptJl07pNMqDwXEFYwYL/TA2AWGu4ii1o5E0r1bmVI2xQ0
1GGOPpChGEhSa/U0VH9xIcR/aNHvH+9SjIuDj3k8PEMP8HmNUGuWMOC8NYG2NCgh
E7kLS7JHgoes5ttW9Sbck3s9MK2cBiybfmqTzVntlsDI1W07exs78XJP8J88ZzE3
zJyJxEnluaBIJEMGBuB+RLHEp8POzH2M79EJ6LB2TKl+b/wjah6y1kSv3e3FADa5
ujjyQRVa+EZjBJxS2mBG8xvqvbn5sz7LF64zRKjHmaOCAwWNkPIRInnRzPTzqwV2
+7ydTXHXk3Gd+BWoni5Ks1nctelkf1uL4hfkwlTjGnqJgAKlXctbE4ShATN5AzSf
CkgDPKwHykIpU2wjlFiymtl8aCzNds1q3ur9e1KjH304HOXJMMz+SAMr5N6536rp
gXsXx6OmFp1H/ddRXSUeBffSrFQPYF8KqzlETmK0CT/dtFx91xdNmf8HCFapb0zH
/4ZqMreF5y2yeDmCBIghvVGZBzny/UxwjxCE3sFILGhBQVyCIB82fAdXXv9DG6uo
eAPp1TzoMUSUaJGcXNgJlWykeYMIfAcUCTTcSCrwtvF16KKw2n9fUNvCyOCJVAds
nYiL/xYIQllymHo+8SCTuPihkOe/aCoIiKbK55Tv8U9XJ4OuywqrbJiJTU5Bcq6J
+sAn6fee2e4pPoQSb88x790y3C0U6sBZvIJUaGWPuGu1YKDYXz1r1r7B6k1g/2sF
BVSRm0KLhW0PKyWlg4ww6bQ68JrjWmhDe8Xxl041adsvlC8x0RZdihR50rb3PoLd
x4DZFIde9X0ASCAobGVkxYlJ8kJCnCT3U6BYS41atx1YbCqf6b0r0SHRwCjUZYJV
UgSIT1W4PHozwsSnhkkrmSn/W81QKjDT7TpSDBadBQ1RRfVfm9chaxN4gyy87gmg
OVNhLZn7UNCe2ygvgr4KUXBdrt14IGwilKb+upyIuv0+LQRhrhZAW8BxMmPt4p0L
w0xOXWi4uFMKNy9uj/0XFlyLLjlkNeWEvFbyZNp1v4BKOGwgL9a+1TdJsBfkdvRg
5E8QAW2FLLcd0jw6gWerHKl3y5hCdGTSXzLksik3AEYI29rIKWKmEWYyWRksF3MR
cFiF6q2Y2ULsKJ9u41NecxDwwh310UYDyzgd2sE/fygZJha4w35sUzcaTklAZzVC
zNcyG8ct6V71MQgWUKAP1lm/UHkGnvaS1H6nIWQBXi/NyM6pg03c65KciUlEerSH
2DsxlkNqFBwb6eRoAntfYxhD/y/bmcuQr9P1EycHS9b1UZFQpzVA9hpJ9WvCvGpA
W6Oswx+ylsIlG5Ll3hsB0iNlhrr5TZBJ7u6xp7yIk8gvN/iMYz1n/YhxrQ0vkrcD
cVePeL6ItopoGgs3XOz/nItNg90pjqmESYqIHqFFa1lLAVrEpHGY2eWFYNiPkQNi
te99hu40TouPp1YBdcdeJrcubbtwwoI0ebGZv09+29FwwQ2CMpKJBZ6I9I/x/jIg
m8pixSaE85fXp1e2fJM530E2A5evwzzmeB+McPNJxXSncwF+4QAEKRNRQMgJzVGt
Tr8Q+mpUwDyPJ3JGZlkaTa1lOllTgcllmwvDUZr69roe17LXy8xXm2wZQQRlmIom
kxtOBkwsv7NlNYPN0m55uNC844BMJuIBz4TAysw5RljAn+bEM1vSkUZiu+59qVvC
HHXkDUgXpyQbaQJdhdFW3JdyLwvUBPxAJ0X+pfIxbNXqUhrKSB5m1F2+mJdiNjX2
/oncPLmVEtOcklndx7L800WDYTQl+w3EdYBd+22k5x1mr8q7Ecs6IXvuNuebtNjh
LSD9J9ito2zkROkKPTjL4RQv18izdy/WnNwjSJy7Ac72Z7iR5qw8BK6b2hjC7TLE
rCnWnH+1I6pq0Jonncy7FtViFOXQqDbVLKgg3L8vSqz+1t5hzecAIe1XRxeSxWrO
61a+geEQ7tZ3IKy4KTc7bsJD8yAYcNj/JSKGQRZOpeTV+nYqiGlugkrplfGGg6uy
oxs5JTCY5lLneLOUGND2YTHfnBTAilHFZrAglJvaLZJ9pRwsH4bAfhniOru3qxnV
q6xA9JXc5wc469H9Ydk4ATFo8lfEAclC9uJDXU6NEb6zF6AE1+GTgK+vkd9rHl23
rbOc4MTUpkQ5xRO52lgeE7GwdJLCTS3V+h5V+Xq/Iq9cyd8j4b8TSwdm07xErOEl
f3KoQ7NCqt63WnAKXWUPbQYZjvcGlC44Udfq10UoILfwV+PSyLLi+tUdoPjRfGNi
YHkdZ1QSYETjZRwxBjlkb9on/bmfFipGUeiCC2R7rmUsP4acm0kHhy9vYEzbL4IT
iOzG7CAY+uCc4ruX/89JBi/5mWX8ryzZDbzeUJaaRzOZNCebTIYlJvSv/VGwhOCj
2t0ijZ5gcKpKlq4GxQ17jiCSlTjmDtLzFsB/WT/OUctKYvoz6Ms0H3nBkWfEx04G
9aGL0P7sHf5QdRJgRIPInH8lXCS9eefxuo7Ml8I2/W7muNKh+WyFy0JTs1ATsycz
bce7Tg2vcT2CnFZjbsqYVknGdda0ZAlQihavg63L7oPdJVgKh9MrqJH7DrECUQny
JMYpVZ2lmAN1gmbtARxdv295mDOOuhSzBIHd9D6VnGvS/dreCiqF4zpz6D9TjZwl
6S822ghemsMooQ81Wxc+jp22m/suRp+MYf3dq8t5zcnOeTBVKIxOucENH6IjAsYd
1c3CinYHLF4sO9bFrCg2s/hwpfYE4Bg4813ecAvfLp6LZvqhs4XEwB6x5MHWkzxz
YhEADTiOClUQH95wfYK6hy43isCAQ4BsUHKubAtIZBZCqf4viJ03n3Jh+m6puRkd
dnCqT+9zzjJMICu4f0yD2kqYynlyaqLcO60+nfmGDL40kXOOS71W2NwlmlbR78Fe
AJxCvdT097hCB1PIFtAnaRLlntScizDdRY64eNnfz7D+I2ciA9KxQHQDEoduFP3G
/QRm+JxYoooC2pZIuPXOHIgy8ozwhDC49yvXyv9byhaIgi7928QKTVyVhQ8osjhm
yUdqgQ/tuoYLVURSC+SH55K007XPic+w5xMLbk9DODjJlrAwgHfF3hs5YO1Mpwpe
cXpPDhEJuE14J9ExZtCe4778M54ojYsRj1fNibSEVsTDiEl4JCJ1qf7bWUuWcgFo
H2KTMBCLn+7JMpWw9+J9SaXQs5IegPACShbySnbC7Hj/Y99Hh8vu5y3ls492ec8l
XRQwqPWTHvWggtOm6gSMIOO88OG5KSigz4nZ46MJX+YlrQq/Yfml7WhYVOU6LBOm
Qk4JvGZavvsziZV1AEgYaVjSqFHAacPBhZYe+1NS9uXOzSIVY8SQH/8VLyYcQVdP
XZKjHfUkgD0eVIAxRnADvA7u9CXelgPbydaYE84xR2WJ86cMqXRgHzsSgAm7mzai
BleHHRB5I8+knAEKk8i4rWyOyfaD8l1T8AuUxK1+o97dm/xbdmXFMECQoW8PYpZo
etD0f8sObbiC46/LMp1kIP6pgovsWq8kxhHs7OLeU/iVZGkx4B1NWms/DEGPjmEF
oeyj5uZ1rilTBAkfDFP8Q8cUjNmNb+F38xa1szeohho4uFKKE7809eiN9S9cx9wo
SQS/dFDEgPe5aMykazaQoeKK78hJDZhFbqutVdBhGzBUDGa1O7bMde2BkulHvbDF
3Ug6bxlk1z7cB3bgKu2xYPsPIH0P6Wu7YNfiu97NMjHRDV3pvn/rEiYsyDcZTQs2
MuMtxsgmAbO6eouh16z2VHhP4pMVNsn0F+iq27p1CG58NF9/zWEwq+3PLWLC6rpM
PqGkqsJqlobpnJ0FjJMzZrXrbm+9cKKDlZONLLiE6ayrNQhHSfm1W2Sfopj4+3fD
LGM4RddhTfyqGWLezsgn5bsiFF9xzdDiQcr8mLj65OAExEy32aA2wVDRqIru8wKJ
5JhrLBMG2j1ibn3ysc/ivm1qQq9CCpGFjTILMEcM/1nngQUZjlAwa2f+MV9nM3pM
R5SiJ7H6EAJWFQ3u7bjN0dZ8jj0RahQCMTclAOyM+nfh9Q5FeBZYV10ZY20gouC7
ZKYRiYZZmw6X4GEd+x1CMHBVLwYaWk4PVkD0fx+81Txgo8KmAD/2LylgLIVHIqLt
hmCx81hcpp9L5cCFSKZcKz8jAj7vDiRBdWL9dcCEDyj38EqNvErtEAl/D4TzBfp5
8b3U9624aNgPLzklT/8PGce44PO9+bVIlGoSsA4TeVT4zUmknq+QokySUo31zC5F
YO35LyAOFCEK3VQLRB3b6hqxsKikkYflZSNiDiJoNAMTgGs/af4hBFa0eFfOJ00p
IHcaQ2UFnWkyPjCd36weNlgJoExzVBZqCoSZzmC/jLL3SLK7dYBglLs8TjmFEePi
11mntBS/5QFnByFCSNsWPDsTLvifbJRNXs9C3esnIXrveSCyFl0UkqZMiTbh29Z9
q+gBvzE2DlRKjwgDzzFnAuZYwSuuC3+Pg00HmH1ulyw+0C6i2iKJf7tQo72WTZek
HzufooB5mSm3L1qPSy5IYvGC+YRZi0dp79jfK7P2X/AmhgzoiohIDmAJ/emcNUpc
GAzPDMLt0qCXYDbtFjt40fA5gKpZ3rTNjtNPkLBb94xoPOKQs1ToFY6+Bldi/DN8
I8dXYDYKREIOSjYQOiJ4nz8egSubLQfOl+rv5vzavITm8oNqFO+uz0ShnulwZ1JU
zV5ldB5lSml5bz4YiFYT5ATce33nMTxZ6YtYkyJfihOBtG6jBwipDYFmvcGBpPOu
7zNvNrUn9qyXlBjRudevhetGTNF1dn8sf5o89/suyu7tTnUx4SWbQTlwy0rAR8iG
bwc+g04A39cFV82y8x8lzROmGcIgYBAUHqWpHR4+eVeO4cLGWUDdcd8IY7gqa1+y
0ZR9RH9FMtovDqIdwd2Tgz43Z2DBfmnDjwxJ6F+r9aXw7q9zqqCxSgb9Vbxnk+P6
u2mIeTcKCobaCZF/0nZtpmWYht6qmpIALuXTeIyE2hw98J0MCdp2kCvGboj864sV
UA2G3A0E/8kLPYujQXFk0z1Xl8hJQTS41jBIAnRXoXXo2nsEJWZbyjUgbTpVOiNS
L+Qadb8Gyk6N/OzKpLVKN7ILg7IjzswmSyenlp/oHy0RJAXJcuzYdoT0mpdTsUu+
NytjwzYPAXv4SnWOcCgsOmaJf8IjWCSKRcDFd6kaHbsEoiZL6JXTeqATBuPYc1jA
IqeeOgLonMeU/ir9rgU8nmfrvOTJ+jDdkpKkcUiNyZsPppPBGTJhbZDOJXS85fvV
KSDO48ItyqCZW7EzB/rnLeEtNOba0qJhKgjpBaFt1o0kVx+ZZyMdp38mNHE3Amcv
RR8wE75j4LalZzNk8P8PZssGxMhcAbpwnvMUlMV08Oo9U0HPdH62wNQq+yHCNVCX
wUoehEWV0B8NN2weCZPguMq8dQfA0QqLXCmkbUqiyz5obXxZWzwLBUAm+g1b5xeq
wkA4z7WgNbTOqRZOA5Mz5QMI3Z//bNsDv7QJjUP2bvsxkZnOAR4a82h2+b50RCQC
ogAvBsk5ReEKxFV9W0wIC890LVB5t0X2lOWbdiNdBPG3XNM5MVUnZu6ihRpsogTS
/Ry6eIMzjuZPXwL8mYpdLVkhk8UP7wuA/D8rkjHSNb0DTNbyw3ys5R8s9IB+P4ld
kZ1mNDiTQ/djO7E1WAzvPf9hs9MYvBuCkawunym0awvxOTYP8iWeyK18pyX1xV/k
h1/m7lfvMWwm4Dd4fOwlUJadzmYqvYstneRFgvhqQBsZsPeDq5mgWcrm0bP97nOv
k4EoMOPMo/73QpxKlYuUKc/VHBI11uCsjp1tl2At+tbzFSLyjg2igpu7tpPpwbEP
Vc1oeeTSglzwGL5jJhMAtTQpl4sKUESotZ6kR8A3ZMTIdx7OSCC7tSeW+VAshU+0
XUwJ2yabtO9nRGslUmiIPUQi88vyTfc0kayR11aDaoEe02St0K0d9nDWH7+R2Rrf
AGm9Q2xq6G+VGNnZVigDE78wjhmUpk34hMYetORGHpwtFUnC9xzUIaT1vFvMewml
ji6gTCTK/D4XhbOd3HNfitOx9buH52QWoMQ1/BDh2O3s9OE8PFuZEudjN/GASiIl
Votv9VlM1Gv9VvrTdGfcJCfpl5Cw1UPY4/v65RHtauntNF592YOjSV9buDm/ycfW
1mtDJeU0TUYXsRZiYl6fzxJJ9yCPcpFr2213KfdlWecFzV8RQnzQmffoueBI2v1/
Ie7wydJuZ+9yxsM2VsfHyczDn2a0djej12ZZ8Sa8tpvTCk+4oEBB2af9JZz5jxCG
2MPRqhzpVJeDvfVX+PvakXnI3zDRpJwAPggCLTnF+Qba5P8szS7LH0BMYIQF/6M6
rr7pD9iONh7FAnbxDl6cZk17M8l7U4bq0KGOCd/dMQym+SM+oYMR5VCur7yY3i8b
KE6s/98K5+KyxMUHYl6cZyk0kZYEzPkdVkbpdP3TUwUXEhI0x96RyNCLWdyuA5Ut
MtKdW9Inq4ikRAX2orobicJDyuryUUGdU4i6erPzftdXY9uRElGV3lyD96j10w6d
QerUumhLaPQHCYHBbkLtXvRTttLu/wxJqTYU7o32SpP+r1Rc2II6mzxCsQvlmVV8
6sjX9xSWYooTDpSBEpCZSSyjWHnGVpDESTzeYLI8G+o1NWGmAGgCrGY2v0Jbvha+
ooGK8ooKLqvIZjeH2/dDVcRhXa3HMXYPTaVbaqr9Nn+7OTQ1ZGnfOQy7jznKnV+B
AykLhGuK1d/pBdXRCxbTtf7aXNWj/ZjGv6toVgUdm/PwnoF9fXGZzAUTVhFfvos6
6g9w6WVRrC4Cm3W9oZ1Yubef+FW377M6tkIop4kYt4Zb17Ey87BC2tOPj3mEG6AE
0UY6wrsy2WKIo5OmUdh1Ht8Ywp17vsu1T8kYjX9Jnuu5BRy6iRiBf8/pYlaeC+v6
vmyStuSawzS8JUFYGADBEjn0GIxgCh7V/GNsOxNccunhkZWbJiorINiC6p69M9if
XItXaBfuRyfD7oIlsHcKA9Z/QGi6Eura+QNVFT1OBXLplH3OMYhNXaNMeJjroBBV
lQkXHr222z53BiAX9qb33eSVOp8gLU6cd6dlMTWjXtZNLNkctYzu2wrPdf5UG0wV
1LCBYvzgSmHG5Mh8yYgqoVwIcEPkO5Ce180MsBrzseeWxouMRAGRB4Oqn5hv/2Xj
3Z5wrhLcGdK8Nu5p09+RW3YBRM8p+zxeWk0ZgHWgRBpMYpA2dxcj0usR9lsh+/ZQ
UbmUOkj1RNtaV/VPVerSA0SbFK14aTQd7WdVBn5gKk882IJhkgm4twPZedqJ9SXn
IzLuy06sGIbrVq8h/LwBg7aYCACa8vTWvgphj8VZGKG2G070LCuCJIhbFxsuOQsE
LTHAqCDmMVp6de6xeHEK+cbe+1x3mpUO8S0J0u5GyzHyYvhgUIu1bybijAbIOGnO
XmJVIrVJcgIJ4zpUFGPOGKEz3bNIUpuMWQCnUaSNA7vwcKJllzl/ctB8qmrdkbLt
ElIy5Qc3U/4fLKRJEj2eiE1ho07VkQuvVoF14sV30Pfd8Ha6azSZWgGSjPkqGJCp
78BYbFy6Cx1u2h+cis8KqfZ6RKd3fktKwMUx1omCYrrdi/bbGaWxO2SefDht8FBe
aBgPXurkhLE/shqNs72DxyZLKaqix/kLhAQBPD0QaKiLN6YG5KSCPtrYJ/6hfBs9
ndn8Z8Gciky9Y1GiPjF3P3NqIJ2b1alIr2ukq0Bc8haESl3/Q3qlFfQ9OBpxTBqr
qfvohv3tR5XBJ93H4LXfafYGP/VjIgl/GFJPkxx7vcPLKwvOM9AiUjct+vkDYIGM
+VlUkwshb4mIeFPof1ff3Hxq45QCpww7s6mVYTFRchRWY3jeQjQ+IPfcB7cCHBKn
XDsvY0Nkj++dfCTxPozDmDV72lmTj4Y7AYhxrNkp+HIEr9ShnnuqGCfISHp1Gx7U
hkhMFsM0ZC91omhE3YG1mnh5Ako7Q4CcYkIlS/2Z6l3Hx901VGC4MbwLR40c+q8z
hu8AsYz0KE5t0WTL1tkmkUUQW655sKqR5gjblP0+LzHtrCNbdC/fs6kbA5aaJnKD
gZB9KTlNkb0bSwmLfyIGJq0qb+VCWSyrtXmCHos2b/+1JI+66XGqWt4qjC1+HNE/
rH2WyBbpaNgcj1Lk+QccMPS4yO/e6LJbu4GE0MU7vlU39TNSTYozkXt+WSPOMNl6
OWvObndqSK+hk6WoQqHdQ3GfxMv/cPg1HUS/WT+/MM6CpfnfpqLuDe0UCueEJ0Rd
2AtLfjeveoF3NdHL1BRpDUGrJgt5A+YOdyBroXU4H/v/j82AaRna+4YHfyc2jqo9
FjQiW48oYg0morJkTXV2ynoxvlWaKVPqpLn1UOTi16oRyAyqPyWSmAhhN3vVBAXw
ngr9gHl+TY3ZcnAjKsmnNmOdLrsDfQ3EbfaL9kfHvWsusLKx/FV7YEGEazljoNuT
wmRWqizfxwZcP1dIiS1fymNRRl+8+UTB505KX77G4p+XYdtUcDtCj6YCYt5nw2sD
RZih+JB0bdgs/BY3b0P/OltW2iTTXyLrSjGeM2JXu/PhnbovOiXBMYhFvbzBzhT2
vN4Tc5dYk+r4YqgrGt/BSULemHoOM+BMO/wwec6X9rWmcclu41VajX8SCdTkPXSx
sYfognT3T3iHvj7g27vTuJIkU2ltA/+1d07r1eloY6LYCo/yET87W9bVOYe9J/5m
AorMrUKIM2FIE6jFd7QPik1oWMvdqoVeXt4Wt8CKK8H9ioAR/LV6lEOJUR37z424
GbwPfBgwPdltWnFkQlYIiGPt4eVQ72qpN6d/qoQ4zCkfee+bW6MDKKM8KF5m0/Eb
C4WeGp2Rng8xPViqBcFl6NiGLCjEk/yX1MZb5cnm2pQmSbGjd1YR1v3SOXqgKIrv
JZe9JsnlK7ME8sAgsufGkP2RroxKgXeX+bVd6IjAfflEGvoBy8pc12wAR/uJCc+D
LCBAu9ZH/Zs4Qd+v6VGLHIDn7TiAuW+gqIPE8pF/1DUHR5pNtznKTVB3xTA5qaYU
VIiyJXx1ywJKfEHWOy6wEyPUCUNQOy6Tb5WeE69KEZJgoHXXizIsZLSiuKmrLM2c
ARZX/j5RiAbxgCLxV9fdiRQ7oqitaBPiZefi9ojtqRJcNQz9bLOVNBvXGXJkn5+v
JML9NfrVwMkiIMk22LXlxhcCmzy53R9hVDP9faIajWJd72pgmKK3rzj/fNxvbHG3
6veTIVy+OKvJnGh/RLCdGDYo5ox7CRNcwD7nmQrUui2oeukvSvNxOQ7lSpwWy+JH
X3ZLwXAXbQ99PLNpi2vKK/0pZDTZQDSnQE49OuJJBd3ChXwlTPpGX+YcRmkFejoU
m1aAOoCIsCFmpFcMhsD3X7aMNogTbqOLQE2m6/3rRNyh+mc9apj9TuUZNBVhmM4W
+HMBt+a+Q01KDe21ZMkem86Bp93pipnofgua3U1wuA5SLKSxLbSAOkt2bEykp03s
kOMTVstKc0pg4duGMCzZXMo9LZhwmIN2cW8hzVgmAaWx0S63zGX+wOW2jkZW/wjh
/PEKaGNe9k79rXskzGg81RDp1agcu0aLOgH8a4uSPZ42D77lAXQ3iAIVZcsYHru+
1XMVvMC/yjlHRiq2V+tS4u7md8odQZP8/CEIXjeMFXcERh2jN2vc79DiKmP3/Jam
mvHdhbmamzXBgPX1MPNZraPVfD0HeRDEWt6WH/CTEaLGQaouHAUIS/qvidc+72aw
miheDJIlnGvh1Xyd0GIF7Fe1FGiPv2koBWbxP/fnJTreHqXD/j+wJOBWyZFh9M3K
IyNk8CcQq8TXY/x/F49Kh/6cENWfAHBoQzSgv81oj+1PnFoXHrkFNtrI/8sBe5Ee
EJnq+39+OjKuN+jSIZrIylItGCe7rrrTmfZfULrOlwV8oVJd4B9NfGsdGX2GaveR
62tqd9/356rwKSWf7wrvgIfvpph2mT9ddGQo7bTFPRebWSoqOQ38Y6u1Evu++FZK
7oGGR+xdo1vaD8sshCu9DzxIHZCEO4ILRPF6AjJZVwCzbj82ItcXqJxWFMPBy9bY
NoevE2pZSTI0S2MT2qHqQFgvM5VjAiAliynLOjEsRQRV9BGGuP94LpSw9+/A0t+G
3PGQbmlUqhlAxwcpVAxlwxOarOEcvgAz/ZhyzBI1NN+Dctayrz2zWF9hk7CKHnji
CU+q0EPal1ix+RoJJtj4x/9LNYEUbkAULlr2O8SVF0zQqNaeLMHZz36+q1QFq5HJ
KC842sKBHwfpR18QR+xV7lcq7wsTH709PsaMaWknqXsx58l6MT640uiGrxapdh0Z
DMb2211CbHMWkPyfwR+Z7saUV2Eokoot5wneyRDRZvBpowm7yf7QbVCz2Kk0cT1k
cVYmWQHbT2WksHp3jZcDtDp6HM8KMVko1xo2HK1OF1LRHrcBhqO2mU8RUzF0pkC0
P9fgCpBCx5GKzwASuRPshIBlzEFa1j0BjteJ33319sTP6InUGa0s+lpzFs+Anl57
W99t70BBrRwjjXhCzYYKf13t98PEst4DtvNIV65BkbKvuJYR1zIpQz07WTGoQoAR
ZITzbzlI7O9Dlm2kq01qjH1QZMwOm8jQkeFV62zJ+XuoTqmCNI3xuznpoyHcBvR6
YrllTuE5rswr3iWP9pvNRNCrlYpHW3MP0kHnXBmWztQxmZ+QpyEK1WHxF06wNp5g
p6uMElLrViVpdZMhD8nt59kv2fBYQBngC6v+nF6Uog21Xuf/4ymsEhad6k4j9hY+
mu4ESue0bZ3tCU/sCg/OC1IYJM3JZP4wJU9w16y29IlGOP8ivhSSzo3CmxJWIbGQ
mxGxY4CtXiGGcYeHO+yKwIa09uOu/NLpDVUP9uAsQqVNuf7Dn2nPq7JqdTzi0cjw
EZLTVTvXEwF3Ju9HHUYFsVrCqPwkIO0mP3R5cl6iW75ziaWAQMEQD5E/LI16CPem
rFQckb0ml34y1d0An3iR6Ub4CT2NylChKDE38I/l9Y7UU1O1GCbf3qcKfofkJFcQ
1K393cI+DnWITUvMBm/anQ==
`pragma protect end_protected
