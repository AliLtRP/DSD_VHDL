// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DYEgmWIk6EdZkZFoQQdw3q+q5UwPqUZfbut6CoTy1d45VvRZZKR8qMUt61bmABDA
jOdrFIjWYt0CahdcXOEBDaDNGbnYiZ3+16n2YdFyRXHwjTmX/Bdc/tEMcTqONz3k
qraX4Re89ZTi8KlajZl1q6/JUZYCV+JX2m54U8r+t5Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2320)
5g430WyHezi/TisJ9t7RVVfN8RIwKDn+w+sarhPRSbrPsOpEYKOfr7Ng5hlIyGBH
MXchdSyguJhJ6RYhEYk9ZHEH50Xgm+5RmDfBXvNNFlZVc96rtQNybB9bjllUZkE8
6vTtqwSjZA7EQ/JYpsP43V5sLTvhYZOYOkKYeJwSanSEzQKavdnZQkKBdbSJXLWv
6biDtIe3VeIln8DCljw8XyxcJp2UcaVA+It1JpsrGvVLcKT5Boli+ysyu4R6Ci9B
DNF0NwQifo5/mBu4t9D4kXe8N4SWDoPmO6WzrsnwxhVaHMIQmSxB0OAKkYNa3Nrg
4muWsbfCx1QCVdl64gHXbzu7YkLBCzBc1F9LQm9QCSYov7PtMLi4EGNF2Xh2zbmd
IYv77zb0msyLA81h3atEpog7lU9AVYpcB5KILcqmXcCKj1rYktlAclCmITfymOIZ
58JkkV5KNU1YHOtQ8421wPdDXa2Kd6Ninn76WDXxN30Gi+KOckzfA8nRrBPbkfxX
fxXoLGBPoXjsUgxzD1nIuDeOIx/L6V0KZsm7NbfKLyE02zGhZ3kxvo/mR71l8XvG
SuyWITqK3yLiqxBJXzA6Q8SvcBf50WT+ks8n5rCoTKnsFagqJ5SnjmNNh0SaDAu9
ThxzAiPMGkDuv8I3W1pVLNVmw3W2O10EsxFMXe0V773WitDR1MCwSUa/NQo3zlNh
MCuLO5vQZDuIZWU44uwUjxNj6nAWscUNM21ueNVpzmB4Wy3Mz5JfacasYz0kht5s
lkFPkTyXVxfZHs5oB6GvG3Yu1Ejjk7QufLq25lqLdxIa/Wm/6wEVIcvZTw+jfkXQ
g5CPSPMJEXSCH1/PUycXEpLlsobV+0ycp6RlXVfBH+pyW5oOWTBUo9zax26gV3LZ
gihxK/2Z8qU/EWHKZU+Tg0ll7lOPR2dqO+mAOKYmn62lMTZy0M5PKt8ctLLShPqi
xUxabksXZRD2km/n+7/b57T0HVf8PcK0l98GXWqK+W5FqwanoV+EL0O+r1cgX3GA
moqAOHl4ByOVSgDEn1sBA5DPVURWZwC5h9B2d/b6PGE97HPnU2BFjLDzQ91X0z+0
Sv0UijtHgIzGGOWM4lEGEwbz++ZQa5hHJgd3K7dMda56rcuhwNSY2ItLwY6JCFrS
CNCOI+7TuNN8t3OhxEW463/fQ7XareiaJvBHg6prXem+l+Q0GU6s3z/YSql7LPGO
8Fl8PkqiY88jvUxeDERBqxIIaV3lm590ax4yE+6A+1QL4csZXmLqJluouHsRo0GO
Y5msJ0J69ORJH2FcD4XhAr4/iJcyZR+QfVS93wYoX4EZkhCf1hgg/r4M7IArgudG
JVoo/pddIYjhYjFHj1jMAYUYgjfGaFvbJ+9CMefBUmZM1gYP/En+cpy075/SputC
c63VXqGMPQn4yeJwjw/QkrjadlQjgBbLxTBAfIaDZ2ID/hg7c3abos60YzfXviaf
noG34ceiBOHcN3TaN10F3eGd+JKJ3Tu5d6C2AVqn3HVaEsj+QdQb265JA90FcNdI
R/zuPZkndGTTIAGd+RPGzI45JNGtFOamNR8/gpERArwk296giTRe7Zy+gTuvwjgI
gQ2qjd3fjrDV4JvjZKVmGz2IBErkcd14oMvqb5YfAiAWGC46Ve+1bMkPqU3yhMMp
F+HWeLzWgvtrt7647iUtsDhU1D8rkj5vvzGl/MZytxQOcrdO5yL05/58ynS61D6N
wkWjMDt224Tkvp6+c6fhjAY2NOxboAe3G1eHvStgK5TJF2y1cBfXurRQ/IZc8QoG
eG3NJyK//W3O6YTBidz5yv+mq5M2bLqMouUocDgkCmQZ1X2aXWds++d205ob21X8
EG5uQUJ2iKRq8MQPl++T9EBmtNMwzv2E1mi0Xukh9zWU94E3HccbGcngHu9ePHSQ
0IOffiH0A7mvW+uBJGi8rIH4RkHimJkW9jZkk2BmPs6MtUvno+qGi+h+oGgyVQDP
neEsIXyRhVT8rNBQiqqjua7bpNJ10CeMO/M8y8mPfrAKTA4ex8+IpnFBJhI3rJjK
bA+MyHpi/VdiSVwaBW+pcaZYKEhfU3zq2vZsBtJQSW3kmPxKPXvXu3rNzbezgJL6
HATsOn50vtevETfs1osa1lDD6muSnr5G1njkjoL1MtiTs4c/cO9L7YPl6IfUfr91
Jn0m2NRRwp78S1Ek/VEgUp8Y/GMp4qaHl8Idl5rguFX0BgbEjG9bXe2zu8SCZhSP
fVUc3Z8dEa2DQxMasJcajXydKAzXSORB1BJNYbgvK2W8twRYGUajuthmU1ZQgUoP
KwuiP+I74ObMOWJ4IpQk/F0nMfirFLOtDdn9IKLiYzmcTV9WkhMorDGgtYGg0OGD
jG7Xpw+FoNbLp4CO+byHiYNk8DghLUnhlQJ3RghDN4xLpYmziVEdl+vJ4lTpomcE
rMZw72ES8UuwkVzMaj9OPtV/HBj0B+6nqpnBIsUPbYrfQ1Dtu4YR/s6+8bVmgHPw
ZXoXpfpx32jFkDdRRhRXsZN1WxRS5yxlpPJUYveaxLNJpRdzasfvkUlM9XIERPpI
rhUWoD/c1huI5DEFuOFCBD8NJg7lCDdTIfhsrcmUOSm6GplQ8VAjU2Urgmlss9jR
Zsr/Tfrcfci2e8LZ9KY+7wCafCgGE92MVbxnE634m8i43hzM/59f9Q7WCI8vGSx7
VKpmB/pGurPIxrYFD+7c1kmzXLQuk3LKhQhujgMkFFe5DbIRERI4+C7TrZW7WSsk
7sVfqq9ZXWZX3Q3nXPM/E1RZS1yMsiOBXu4jXyW1C830NpQTg8B36SqVmVC4dgoH
a/RBSXH46gv1iU+crabEzk0QBTSenFHYDyH4duLFuehgiAtm1Xv36Ubb8FZOi6Vp
+YyB3FmOC11gYMLuMJcS7+StGc1NLlC+kBtoEmBCl2fkjWfmETk1e64iW0/BpWiG
/J/BnlhGbzSI1tD0H7IDgAIYRHyiqakDiSB3s3sSpv+OEmCyMQfznRczqoYFY3Dm
CDrhNv5nJleTS+x9MakG1WFPaWhZURNrhMf++4WELipyOXnWWDKqrOaoS1pfhPY+
YFds+LQPorr74wRWQRZUGQ==
`pragma protect end_protected
