// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Upxx6naF3FeaRP5ajKs4UvG+EN2NtydrM/TaGlvI3g/aT8UMvsaT1GxidYpfl8bd
pvj+XKgSphuSiGxHOKTC9XjBEE9ALbrmWVaUtaJZjwg4+QpS1EL1lRNmx5g9c90S
0TAl8l053TWq+NMVGmYZfq7+fO14kBNaaA4S4PMgdSk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 90288)
590by+e8310XymAWgws3eE9tz/5+Ol18brhGNLMSg/zIlqRTconSaHR+BbmSG6PO
T3rfsY/rbcwwnr0FuiE3iKoVuu5R0IrU8sZgwSAHBA8gKyp/EyaP5I8jBaomzoAF
kS4ISJlbgRh3QJMnxEnq/77EnBqg9fDeyJessBXYylCrNZ+sTED8lazJd+e/vFSp
xow1E0wTgucfzZ/TF0OjsUYrLlagxpuo3p0izgdmjnz70mU1PkYjCmHI4XMWqOmM
/mpW/vzCG7DsAM7OFB5tKbfimXVnJmRirdugSCjYfIrU3+fIIjCeFkZTrTPn62Ga
2F+UNUFcGmoDh0hLtb84KxJLBd5s+1QB/SCGf+pFp+tr5YTfdIfHLOncZUuSVzCr
GPphYaBgZqt/uApnnlW+hN65rO4ehpjzdZqLbWv6FeEIem9E1KKn9+badmzsH2+S
CuoQfFg5DraJ/yEMyAkMHfUxG0T48RAK9BczOo4xyqCxPkBqyGE4TJRNxtRAWyx3
gH33gmy1DWnCGPKyklMS4CH9YivxP4Xz2Cy5IvQZe9OpCVy1GoHvgjhSKSLbDpin
0iuuJEweJcFpsV8G0WoLJhoChdfdkZvpU3F3KRpE6Q3Habu8i8u7n7QacdJ+JlxW
OmoMdXIAyRa6PaEB4VQZXbhxGW6zT3vWWNyCbdyB5lx0jdUXsYVbFByAsq9vfsJ4
FfHHceYvBClMDCMCEG/IniX+xsauA9oPDwwDaeQZnmImlLxpx+UQC4w644t6TSgc
Lul85SuhgIFAjLynPoyl9rjvxKVQeIn9+wd+RKdcJ0/R6R4W6xSD2G0ssi/EE8f9
pvCAvERE/uErw9YREskVoFaQL1ue7jAG2sRYH4Ov5ObAEEBQAhdW154tRYIkKqX1
qune+un6ukmA+sTcX7kMLBuQmYBPI/Bv0TtT+2EaQaM0w02DBfxso+blwiYbucM5
x1YO662X/+4aUQ/rN1B8wtqDffs+JrS1moCPvoRqOh5uw52t17p/7E7Kep2/CILH
S3UlPMq9+DMiv1CO9AtMG3mQLbCjSDKTpdOZ2qqcXQdHW6xnegxMS05TBhHKoLww
jkdW9eti66aj4S5NmtLTjCiHC8aLR6ba/dCoLjhT5L1UH+URxQjM+tPqh1ObahYM
Go7J1cLN8Ryqu+v6ZsV7eixkYOacg8H7d55aaPX6EVXmaNX1J0hC00nTZBb8xPMF
2ewXCNtRkj/AV8/mp34ok9w5ialYUJbHIk7MSA6znrXZMH2ooyKUYkqFWcP5E8rm
ZVRF5XrdiCjaRPQNwZ/3GD7xNtlb2B3T4lUpLXGhuote/Ej4AU9L3CT/ZSFDMK6/
wYMKcPNVuvnexLtQYJdU7QVwoTX0y0TQ16kx6zrXxuoMavomaq7lGrVZYcb8dREq
x8A4ztakrLkG7zKof6LCIkysyP5EUmWxNo4kOnfbRPdobe2FkOgUi7Dmm8qUD4eT
Kw3c+oAM6U1XLfFJu/9gqvW2idvygIo5uRCjwLoRI3PaFKUQBQ9RbDqKrAos9QFB
Rsevd1vbwvNLrc82EOEnZ7huA2rM2/U9vjlq2O+wWwYS0Pqqmx6OngQCfwNabt7N
HABKdNS5UcpgKF7o9hkLTZge+oRJOIiNXJBy+fLZMeZTToqvWY0LGF05q82x+jac
bdtGR6xvxCwMWTxcrNT8OLWEaD6fFS8ANEI6Ms7ia+rS+jppC8L6BhMOVdw44Wtr
9/0SiZFMQ/kTJyCs/3gy0d+ehIXbyjuwKHpKnSCyxDS6tjFshDvirNq7LTANcVO8
DraMS0Yp4lPQcK+D+S3ycZSpeLWuClhQtmtasWURsVbx2CFw8SHy5lUD6Rno3SOO
Q3y8ZbdyWxKXVA61qI6JrhSARADQ1SVnRgvp/CrFoKL4LkbZNGSaPzJvVXoiGiGy
28p4caz9sLekZQp78kayK2961NYpXpakFKKN6X/36DSArKbvP/PHAoz+EoSOLIiK
QdkTd/UlyBn04bkecQ4jrFyveyPJii8nXALvWqK4PFPzJqqIpi7A9ryCN0o6AuCA
f48Enr0nvJ6NbErzD2x3izHt7PWed6jpYt1FvIyNtupPRTPQs9qp8FWo7yIBEhSG
kYzmSfZ/ZpAirjotxEaVyykquI0rSZ2TOCV37J4yfFe1QVKW57Tb/TzQ4jDW9RWQ
G4y4SZNzReqwDyauMhAbRb3eoMXLGlgN4QxCkug8rILtA0Mbyjo3dlzFXZCdUN0w
TRBoHyzkLKqzxMohQT8WgeDBqQBQlTsvdYR+TtqNDBqEQWV/xLXIJJZCaobPwzQR
MNhgy+P0OFVobYsMur6mPoKgpQ7wmm5XXRy0sGWNE4Pl6MlcTIkCMN3J22vVMz61
DKw+ZobYbRaij1zT+jMo0FNVFBwjFmFZGxrPPqHx9HuOpLq8mhSRJozcWNzyMv/W
MtEAZlJdr0lQG7Gmy2NReLw14QHXwFZ4XKAJ0MPnVEi0pNCkyjzU5J2NPLQ77P0I
7+5w7oOLYfnDQGwTI6V1ksWhLGcuFCCqAKMfXIHch6b7C5C8gI7r7giWr034xO1R
fJUJ9/2jHGvGo8j1Pt1M6lbgA4YJGVaQOvSboCOAULtDVzBg1R6GR1K5DSgxyHaj
2XRl2qScT4QP1aF2Ohl5L6t3BArZzf2CRGkilW/j8x6R8Fgj8b2x+XzJyIgeetZR
roY/Ysk9ajHvXio2GO12k5PWFRXguigoY8mYJFKOWL5xnMs9ISY1gia+2kCCkfvI
c+ZDzcDnRu7Xg8f9u92nfOdIewpI/qg+DGEKeKnHR+RWQhcDcVe9wVZqHSIbh91G
96LOYfQZy/1u/e9HuVWIKDbiFjWo4jfadwlny1BjpANzqm6+2aW5h3nmHjfbl6Eq
rGDoVJUA5cK9te2kuE3fhrcsAM2UvxSIxb7/ZYyf2vkqXW1LR7B0NE/FPiTxeaPr
+49mb1oJP7ql0pOCjdQBifaRps3/pVvoz69U+x0YJtBHu20MpMogEu1TeIsZXYQK
6gboVdMMWMMBIfNQycMypeORBZJqkeUU2S1zUJNPojFFCmGCEN4thXqfah34AUov
0a3QUQXtAXUboIK8muXBpiX+GyOVIKZlndcZ7A08VSRurNtRD5q19ZRVL7LJjH/x
Kv1geE13/QCIPdQCFDnpYIgzkFf9pAc57t8TSMqF0z0rG/tCDSe5GHnpZz3UHauC
B4rwvVmocEISyvIuuL4KOHYql0eTPYbKbYJlCQ8MLSylIKspRu0t37BaPqNjbXFh
0d33WjUDdD4JRkRF4eF5kVqiHxUYZTIHZXQ5u4qD6Rb3OEN7dqVpiXS6q09qMmCy
ehYErT8bTt8mh4mVJfkzNf9gxEPmT7pjtCuiOJyU+jlLwB5j8SUf0IPEpK1bq44C
k91JM7v5yQBVzuhyFj7AS5VEkDNX0ksyoQpMihCvlsLKffVEgweDZzZJ4lgYPzGL
5nF9S5Z+oGGzAqwXJ5V9X4hEAoAMpvei8Oy/QTKuqMMvMGKkubzDQlJf93D8Seu3
5ubj8H+cVB1hA2Lxi99XD4F2BwTj6fZ/Z3qdLoly2HJOVXUlC0Wvz8LTZx8XP/UQ
NVMC/W9yrcGCHtvEhAAlAoZcJpfF7PVsdcrWIt7npQ7sdZ38M3svXCo71Ufi71WA
D1D8Crlv44zdZHRkgSu4JCCTEaknnTEGpSkScXuI2PlJnHbNOfD8tWWNOYwu2LuW
ZzdDZS1bBt6Qlj8YFpwVuPaT2Fs0kablASighEG9Uy7PBxomO/bDXjtEdA2X+zqW
E7Y3QihyEcWL8seax4yxCDnhx8mDGq8mOHtGkZoH3F9/Hjq0za/ex8UgeTqAt6un
a4K5rtG0GHw2Sf702h1YxzRvqn2Z/AuDnGlMo0/5JuZYco4zHQ6E1u3Dmst9tPwo
VQ062wFHNNoGyj6GiuoNQm/PqHR8zaQ2wd+gIWQJFkJ2vqjk/yQsUMyWtmBJ0o1t
weB/5pezYPNnebPYQeWxdkIMQcgBQecapYbyj6k15qlT+EZ6FzLcvtiWl0JJehPp
UnxxJE9Mxeyfrfkj7BrokBRvhJ6mIt5ikwrcN7Z4EH/mC0tA1xfhvHgWHLkkDxhx
X23tvHkUQIlTZWYrWbZ0K+Py4dMccHa1TbFq2nOVmxrHtgzcpply8sNCp9H0jIJY
wa0ctV6Kkhdg5sdpufD4upXBVE2jqwD2ynEdNr5hA2X8WQQw59kkFZVZpysrRH0D
f4iht0P+yrguqDDlc5qwzje2TM+5VMLOr9N9u9tx0M8+SpH1RUb/sW3XTHwdQrxV
YmlNG2mro2zt7p2YAJ5WFxWxYbxYjrRoqmPI7bNRygXo/Dxl1jR1sylDDWCh7QY7
cbAib6xqlC1bdLFqOa9Cs+JmFsWxt/nA08X9RFBG3x6KptbrXKgU+FQ4dS32EZmi
MvWPbmIf5aQFHACyIqOyySW0p1L8/u9gsBylQxMerZO2UhYQs93vzJB+rOsdplI5
1BtMy2yTFT0ZL8Qa4HtXym8no2gVuiek0e5hO6+R515YXg7QJfsXosvoSwJcOgB5
N+SMRdl7grnEaNE8ZeedrfMi3WaAU6U4su3sBmt+RvBkis2OHapaiifq1oC1NqmH
4wjHLjAGearTKe3fKjkS5QGGIRKakHyrgV6dTZfBULtmfwvlou6E3Qd9G23LHJ2s
iL3Ish05Ord2qjlhv9xBVaYAqxKGZdZglRBnl1r8Y+FFDTxPZhQSMzjsE6D2iJMP
b2S++fCa0FBkYz18ZIIerS/gkzyflj4kTnB6QnueZc1pvuviD6P22cYvRT5hV2kf
a21xSXKmFSW2SM7Fppc5kFQPDRp4ESaV1+hQqRTRPdY//K6OIIv8/OuqNzXgGwh7
sSLJw2WxuB2ugexuXU4Mt9hhC0W2xsvf8esBZfkb4enRwiehCLAgQC0wR4Qcy2no
m1/auHkGyRZzUVUBZaTwXUa9fdatJigQ3et/Ehpc9assC4vDWZf4A0Ajx48S+uRb
gnyEtv/4P0mUcpzWdkaYz4yQf3frNeSuDPhlsi+5Zik4+ZPQChaQ2+8fa2BMoldm
TtFe/GH6ESnPXD9OIE7u9I1bkrYfvk/f70Usyp0B01c6t+qEMJJyDql52iWohYki
PUnPnpzhZ6rJ6/R0nPEUmNNmTSCDRJdNncS+ydMnKaCnegoLMlvOnRirztllkE3D
GwWxAoRgagOY2cmtMWRZkliXPdJuo0DcIPeIyE3z1pzWr62ngwD2TWAbWn6I+10n
xIt+tVMGDYANfExXc1XCCvpKXD6CmJgS+4zvSQupAcQYR+M+i3gjtpgd4xXqpPRC
O2HSRgLQqloOGdsda3A8QtkE4zRkdeh7JJyoo5yTYNQIh9YbfL5iLMcZNUe8E2Jn
jtUlj3spNAUJqvDbJYwdYr/k9q//ynk+dHNoYy+GM/qrU/kwgpJ9FvxUiAQMw5tV
f6HQAx5LocARFfFwN8HKlVkr/PTNEhPhsVw0CVg0xwx7juNkl4DR2Jfo2+uBihBn
u58Ggqigq6sZLd6Vp5mqLF7XqV66cLCUyjyUw1awDw7kB1Lqx5Tb3aDtTcZK8PRM
rTupub9AB0gYohM2Ou/Ejqpma7eraMJRxW0qd5gkHLXJAJ4bir0bRVIw1DYukBeQ
iZA8zjv+dzeW2jyGmu77rYHlzUXZD+3Vk6sIVN9JhU1EoQGdB95imAZ4e1EnXbx1
NuJoX/hdSGvr0ypQE2j1qCs6QzLhqxOwrcbYQfUYedZJqGiRq+yLX9IW5x/2YSFr
oZxKm8g828IrUHLZTk2zmyLN640GthBeFbmkAYeXvzUOEZSBH6cD7ZKFhKIh1a8y
71UFG6ows5G0SleGP6C3UBL52tKGxfulVUSUWZF7WL1bOw4DAEMEA9y7x2NhPCmB
Il9yXKLJT+/rWoiLIpFRppItCOkfMm/5NUIic8r9L/wt88g56rJ6FMAAoNNGNdN5
spxw1Fv0rlyGzhJdJkRgVzkWxDBpLdoGGmmR3wWTB46PwBjQt0Y2ufETpJLso+P2
E/tTWPoFuyyqOGl0kmAHos2utAmLp066sCOf11E4pMyqZFAEh5XyTz7SNx+03Dn7
2oNycSJ9zjQ+H95cLlYvaDXKd++9GltvlsVTZukkxZRkWRRRVdV9MBxFD7mvlYAy
ySG0h3t7/gK4S7LcG+AfNGTtSV/Be/HL3MtRBTuXs4a+nrDx5eifvFNJkDxUFQfv
z3roEony0AYD9regE19HsLTZhVwh0R3fys78KWVNPyIXR2CZSabSdC+jfTZmAGxk
G4MOGkL0hB4k6l62+KkVDFYwOSthUh/LM9MZirGvDnVuS5g6qm0k4MSWxrwGGjkv
oA7BUo+QfqwXp8b2melNEGmLFt0Gqu32uqTc+81F3tQIscnFjgEsHMljx1VtLa70
blW3lu0m7VRQX1GXX58E0QIXPFXxslZHwgXDa9o8uMzCLAZXiOCrscgohLtunYN3
/YyU/8alHoOrYde+yyNCgcUCygnFWTwLJwG0kEaQ6P7ztj14/IqDMu63kkmeWS1Z
cVvESMx7uTxJxkhI+jUEceCsrnFd1oJ08YsxetN0q66JQt25L/sc8KfrP2fWz0by
fV801KgStXAjIjdmLDXbGyX2iTSHGk8dhl4hA+g6g/KxfTa0uQIyroexjkdD0TMz
sZy6x3KcD40SV3dxhRloAfKE1yvz35TWMRlcyuqNXoE5sKx4FuQ7nbuKVepDVuzU
pO7Aiwn/mUo2nowPCEE5dFuv3eBXnCn9U3j7AvAexTdYKGdGPPBcB99mAp6liIvj
e8mdsqq8jt0c2Jo/TEb3fbKfL8Xs+Nv/4MMsBTkPrsFWYa1uy1SrlLALFmdx2OdX
pJ3/ZHh5do8szfbgpNS0NpKw1B4YDkvegbL3DOYWVwRU9JWipjAmbfd15kMb5eJd
8xATi0w2Ugjj+mIFSCMtHTHwDbLN9J0VHs1axvNwv2C+EVs77Zd+3Gjx4HlRJzeB
34NTBwkgR7pvChbyMBeKunCbY7R706UncS1w2Ru0LfeLr4mMrrP8lFBHDjTALZ0H
y9mGHKmjXIQKWIzTvRZhWoEOghKRxvmU0L/RWy1KNFTYVlXx2/tSmvQXgIMimMdA
YJm1KSDKElkR7ASC+9J/BLh0PQdFrZvSTB7rJcQYuIgaYg7oR1ce8wgPrIOhpJ6G
cUdSMFqenlOIoNBpWfQVQNkhM6xHdLyT3NusawTD2dWlWcZhR7pNzzOEYBw3n8+P
XuRz8Z+JO6Pm5oQb7CIiUewvKAYWCO+u6n5kakzsi2uYV3Uux8CcNR+Foo7LOmeo
laqqVyYtsYCHQBNiv3RnX3X4aR0G0J7kQiD2D4iOJRMTZiVWZRQIFP3X5lwRpKdv
6i/RJcI2TLrTFGIuBHZGa/rrgT9ozbRH7hl5YMV0e4xDFUCdXL9HfcM4HtpMcGLf
4L/GViqybigH4ZywqC9iKY+friqWyO6DFWkEErod+Xdxf12YljFqmFObmQ8wN7io
+DrENWRjEBQCPE0fT9y54hWAnDY4HxuKRJ8gLAy9oIcenjVVfx1sP0yOqCXusU6P
2YOvb43rxpYBAhcFdk3iJX5vo7BNm3Vjwgrq81qxPb5eMuUGDWr4I0ODk6NDqury
f4BHheW83yaQvfsxpT3aux3IIerF9TQUAgWhK9MUtJB+8y6UFX4CLjYCIu1Wjh/m
mR5/YJ5AC0HtsVX8nAPyhgQofb99hgJU005FYNgEYFLv1Yt8o1OW4/cd2JXjXbqP
QD3kgMti76tSG+BfkEhKOVRksBqEdEpksekOOQ1GKXfhLUkwD8/bCtGRVq49VmSN
aJtRsvET8pkVrEQLscTUQZZC/zk/y6GbdedZ47L7rUlxcloZoz6QrQNASDlMY03W
mLrYDeBJZGMsOrjOWntiFD50LkmGFFROWKD5NGDpJzXekdSXIFZi6OrA3hyuPQGk
QDdYm4FsRRAlulf9aeeDlVOldFCQq+O8lclIXAFjFHmWHl/K1XmE5do2V1GfOUDi
Wf4KTFz/5DRjwLH1RGGuin39kYqIcoZeX7Y93TUgkB+rHM84fbO54Ha0tN4vPpST
fPYYI6e1mudYYNwYvXrLSWd+eYJXfXa1Ogdddv2Op4vRCyEHM50SUMB0BdMjPTHY
suTfa8s7BsEDErCyUx01BTn8ATeq+RcfYB7TBOzjtvJLs4pEychwPIdv7b91GjKn
YWpT4ZwkiZF5S+Qy8OF2fjp98bWdh8oAMSWM6OmMssqicWHUnZAHpdSmrUdC4n6N
o79xn19uzRRH//E0mU2Yp8GzWPaGVTQhBGxZ46nOVjVRSoojknllx7j/PsjA6FH+
BrlhvLFxI1alWPxbszgssJxqeTmplUYA5XdwwEWBpqhQQdpf72srgiVe4HiJiDxv
pp8CmghDFj/NkXsxIWv6eb9lTdwSVHDBVUUCgecXocv46cefaAmAcazDkBPh9hkv
iS07UsPx1TzzNnN+rv9oD7ESSxslj+Y/3XxmEVEN3dhLddl5MHv/kgWM3Sz+0mbN
qQ4ZWBCm+RuB2qbTspLB/uJ7+h+75s+uPiO72k3AXwQX4aGvJQtDbsPVmxMI93ot
4B/uXbQF0MLuOjt0dJc9ANr1ufWfjOEHLW0uBmtU08gwEDMDRRLWh5G1XDAsNJQY
ZxNMdxP33WhzBZxI3f9ahAzM38PrRDobTlUZdh0/OgN0psVqkXKyB7mJOI5UHkS0
koL8duDHmJ9xwQw8Y4gnIqzW0tT2gBlpGwkI8svMv53NdLBm6JxBDSp/VwK11P+G
IPc6jP4L8iCLXjU9Zxzwn+AOxQ5cUhhQneE20v2GWIG1rtq+Qt8WxgjMifSGc4Bj
XRNXN/YAZNovsoNkwzjUPubX2KKuyOTS4xy5Hzc+b4Jai2ph3bCKwubNsrKOlqC/
SnXgQ+wLUsNTADNQ2uAvIFjYZLm6n4iiL3JhKR8eJ9InuRluh8hwEBCvHfw4UQPU
rg/l1R0QuXK1Yh30/BP5bnfNId6ic10HZz7VGIy+HY21n9u5uztapRFAzSWhulCz
J6IOJhQSETdNZU3nfn90tGLQ4JPlPZtp4tQA8gzDGPnVoGtkuEg7dXPtjcbmQMJK
2DXAcGi2NCOvW1EzL9b8GtcNJVPETkDtciEm8780DK0IJdJMFXqNTTsKHZYNp1E4
YdPxjWVaXkV80lnEl/5KgFjHkOAC0c7Gweh+q4xTlJr+a6s2wRG0bWxdMqFTVTLp
1D6wJgo231u9MkKqfs0yEhlNl+TnkpKxHmvzerdFXfLEyichm3ray5T2Uy7viNAa
QgRGc6cZQaxTzZOz65Hr9SDKiez5dSMOErY/U6UH/KvZoBiO+O0hbez0QjXOmaUO
k7dI4piVHtDcf+qNwrAGbKQa1zrdQryLCiw3gUk7Kme8cCUG/7Q7/vNPL42EYORj
TXnyVr/juzvY3+FQ87b4LT8hPfXlxdH4RBTAoBEDrTMQzyHoOKHzGRKrK226nIDr
3pHvcZzk0Wt1GojB4ptdmgpks95e3nKWyY92lhQBRmGST8Qo1qjgELJxNB0Ks6uM
MfuK38EVsuIe2L95eUgV2WCGOItGIoBeWvJbLAl9zqc/R+RY1tvtRGnROaftufPG
Bq7drpwmnFYaIYs0kKiL9q6jHnAnsSnz7HC4URHiiEJhxGx8dZIHPo9o38Lpsi86
rdDjd/YWhPcWSlW28KuSnZJBxI+kShsOy5St6oIYySJ5xKMZHtoXrQGvhpn4mPIh
z/N9ILDK/pAMNGOm2Vb+E2NAEh1Ct7NRO2rj0gMhKHmnz1qS8DEQCCKfKOi53WI9
5aL/OI8FC91r1aiu/PYJJm+QhmvT+siBmvCvlp/FF5F4XGbpRluZtCVJiAC4aDbg
ksfY5RJVehRwTy4YTsWjyRChzO4iivL6Pp62ofTIFykj9TEh/Zb9cAciUUGwtRC9
tfdZLY8Hggjc36wtCTbjW3K3HLEEJxU3qsuv7U1nDRMV+rnLBm/gyg8fDj6nfHxf
YD5ddyWyx4j9mCdFJDMWeKp/FLC11e9IDGQNy101Xaa9y2bU/+W6BzYBNRgd8WqH
CsDIkHF1tKKc+qW6+3rzzZ0M3lmS6cewJeWqCcTQzdizjI5wsCUS/W1hRNNNEwR6
9zVQrTLH2eMwuqIlapIAuijCIfHobfqnsimIAXoBMx9NWfLv48q/sTGSRHBh0wRc
b4ydi+dDMhCcrXJOsm8lRF+DTQmiKpj4DlVVs6GQE/+q47AGOsB+VRrkqiHvLYP8
2ctS9+flcAxuL5oC3C60oUF/2E/ORsezoe7gLdrR2JbkXs8YN5rR7NsBXulrc9zx
vMahRBqXJW1M7KAZDzeKI+fTaVmbE/Tvx1HW9iU4j/ns4RAujLWMopOfkZ23tDeV
lbALcVyMQ5taXh3y3EsQc+JXY50122BQhovgrlmqazvBAe14NjkqCpTatkFSDqOz
IAb5lO/5QDJy8H+gChjvTDAlrEB6NzMz6PHHjVpHaSj424wrdGikEabY+k9GRmK1
gveSb6YyApib1RIYk96Ji6hxAOeyougbtB8qXhTiEigXk/wZ0WhVNRcjvKx8tvD0
ka1pGh7DbEKuniw80hQC5EwpzU08YfF/WMu8S69ARWSYLEl0SqKMbjJz6GbNjw30
TK6hJfVRTBU0ouUJJzYWX7q8Skv5Nl9n2b7rSEY9uQzZFXT2YAFZSRXJgOoIs1mS
I8EMLb3HlLYBfoPJ34xA29s7mQy651783uKoSqX5JTscVgcNzuQ7snIFyC+er1Wy
+Vp7U9TsPCuH2yG4S+wP/zv2Pug40rcbAco0t+4UxYVU8ZE5ia20ddI6cYE+Gj63
nGAOC6gP7gErUC3Mc1DK+qIc/YD1fZqMbrPfE/os0YbsLKuK0N4PTuzznUDM3fBe
TFCnnZ68STiDSlHHSh6KGFa6MLPBNz22w83G5P/z8chtTPLJA4CDJfj0B6doycAg
T/GfxxLIVxhQvDwsYuxoSRdHgZF8otE8/54Zi3ZkkBWr+b8tyM06ZeNcEp1oP0is
VPRAoUCw3WbE7UxMILCEtWZghHxZzT8km4gHEr1YJK4b3FbLsi+fv52nCPVVQrDq
HAUbHgfEdUG/lPqZK+Ydb3yTEwy75wy+AbFs5k/gnrNt4ZNlzmbRLcq9Ym5Y8GTW
ibsE1KRSTGI3mm8zGmc+2PeWnNWygu1iaJ5GY/r70Xq1Pbi9uZ5FfaFvH2LmqvJj
qBOOzwF0tXAuzT+oAXQNvv6x+COJxupSV5/1s9wq2q4hZQxljMG7tdcSIMmM53gH
RwpGJVXBrqixRmUIYQWHpTfKR/Lig7agfXSpMowLZiD1uKwhZXoL7isCOfz3o7GD
Ij4xYeohIWYl7615uUiGWcHCo1WhrfZkcKA0ypp6YjbO0r4MH5fy1xyNUN5G3Gai
EX9DdA7PNvCE9CvAQo2EJYK1WDpzw5uOucgL+raSAPzUtDIzibldsuiKtzAy7/q8
Mhxz6v3qZbNlRzF1+mWSSugVC4m25Luk+FTdEEwMxDbkjklNxI167AJVkCt6ZHau
eqwRAsbUlhQ+1YSc5zPwHJSXhM3ij3cNHS3TKnh4mWWMNBR838Cs9ezel6huACHe
tS7Ruo1bZ+X8Mvpw7Yh1VxygeXyagx3R5BXiW4fICB90szxIIV6k5ZAZ8lUVvcpb
YMLqeZve2WQJtROOKaQk6zwY6lFNNlOaN3hu46JWHapWVOlkCoh24+c2sCEEQecV
PvZoc1qSgKmeVy/P3OFOgK1SBDt2lLH21MJPbqj2GwfZxuq+nvA/rrXT0VfjOvAJ
cQZZ+xSAjdrqJM0LUEwep9KDGnfiRqn9ot2MKfG6WGAVXm8pVDpmHN5rfS2Ua+22
GoQ+DXEzLIP1JpS8PEutPdiix8zabFNLV6iRUiVzMNB2en438wGftF0rirlA9zOV
MBbVhuE+MhrA5nEe4yqTVN78AjpALSMVa+RZqE47SWXwxl2egd9+9wkeSa5Mwese
FaukYH6MkuhOpz4AN9q1xzRZle6pp/Uxrl6h4BAZKJ0v0yAPoAsaDDyCAwbqC2/Y
4sI+r3OlfVabQpKTj1/26++NeInC9adEpxV+05SCelDGZvHd/7l9JemzwU1S7Hiy
5a4UTG/Yuo500++me6vKdD4GkBTNJYtnBBOc64RYv4R60J9SImtguOAMOv78lHzt
jinQmtt6bxoYywn/L1IRGYi/WZJi7td+vf5ZqrvnMS6vD23iILw+XcxAzYvBZ2PG
94i03h4Z2ybJxr62lN5Vvpah30YomjdexPmWTp6WPpMLnOIxmm9pAJA4fx/H4Khy
jsSyD7Kk9+ATsDe05F5JxuNzc5e23kduWuWapGTC8geLg870PD+BRa87N/Lo6OQo
sztp17UEdPOJJ4e9GGkrJJPDS3YZxM3EHmkqyxpgfYjrftgqbg8h0QfPIaub8RN0
iQ7YmJKzE0D68auKcx4b0k5rjrdXyi3hXTSQuh/XaOXJMpAgO1K2U5/G8hLjZEZw
HYFaNPXbA8SZpzIIEqJ1uS6eiy6/uzTg9R9enXQz5iG+kQVJecywGlU5nWrDEl3s
s1yupk+WWP5zS7kAnarAMExIGB6FC1BGCKpY9HNa3dzaaq4plVDi7vID8KFTwizc
Y3sctE+bpzHkhTZ+a4j/BHpK495FsyLPV+EgVL7VXGUHEwjumoOpmuhNqPTLAvTq
sPn9JIfZ2Fh33zfC7PSY5an7qk6Sdf4bJ9FnH/zcDBxSHcR5D6k8wgY4sJjvDl1D
njI04/C1dnzgLBazUre3s6Xq0IgV1DAMWGT3UBVFE5mzOjJrhRDcD5m6mYotGfa5
CwA2H7n3RKTMNvSBCC25ICOFz0KP8scg7d9zLIJMHC1Tshs5uuL3tGYeiXVLhOoH
o/afJxZuR9wH1yKB+qdR+y58mfUJrDGcSs+Hp3aUj7fc5L3iOI6kMh4gIY0/34zS
2/8Pwgao9VMFjPF8JjvLvVgEGoDuk1VEI4RhDdkWxddSb+J1YG7Ip3yV6KPckOo4
WB5I9mpSFXUqxpkFWXJz3JSzso+nOE3BnZ25OSAFFkfTt8RoaBwDuQIs//KVpWBc
8daB1Kscz7kAKMNn35tx6AM+S3eeTkm/tzs8QNxboZ54RrGvAH0FVbWPHOxz2XZH
KWaQ9Conq2vrmwGXpEizoD2tKw6cX3U+m0nmx7MkQ/vx33TJz6gsTD+3oXHlTl+r
NDhAN/R2FjKABPezwPF5ZmIOcJWweHkZb96QTNAbYAhXWF5c/lTvP0jXxcSlgMe7
8j4P5ZXwM1yIdC5CyB38kmJXFxApxqqsVJ7+/IC8Cjx5MOhZJ4dHXQ8yb5sX0C/7
YsfcdOZkQQ1TSHz16irK9mcor+TV0u0uA7oZDHjTAMV2q+pc/1lZWVUTA1MOCeh4
BjOFe5WnvKm1WyiFTwVwTymQvwJ07zdi4X1b9MczlqHBdywzfaaeMuzgU5gYq6CS
uMMOS9hnJmVLH1Lp9ulicJxN9TOMasK7ZcMoKgQvoy36enM3lQhFm3p5vdGkMY11
Em9FMqhd+/wtlxLP25K0NpUxQal0CisaaGHRA2smhtNJcr62Z81T3FWkO/f3p7SM
7WQNHGT++bvktTpro/HXqbElxvXdKq3N6O5yJgBXPalG6orHhjQ43bloPeDpo1XZ
iwykjrX/qaS/x/LDnPmBYy9xhkgxkQt3S8UhaYcFhcMSqk70XoaodcMt30alsf0W
zkWVGLnQ0CKuTnqD6U4X57pdGA/PiL3AxKxD822DBxmy4gURj/y61uokNqRrxmZT
fmb6sG4YY6pyFJlfAj76SI9jZt6T9jV0/oAXq3IKH/G1dpi3Ko9fJzINjc/65TPY
3x+jKL69F1W+IUMHJPOqmNbFNxT3f8iI9OiLOYgOc/sN528y9/1dY/I2Cobq43XU
6hFvfxFV+fIf7E84SQJkg9g2e08DE0TEAI61Ik6hHu8g6PkunQWumdZK1gWWKG/G
BPNYWKexCtPkqjLGx0vPFAQtZgcDJAzJJySylpI1IYg9rBrvXkzezqDg8ArrCSfS
/ARnQtKNt8CvcoQhDosQPukqfYl7/75jNQD+nFqTCCvOLiP8SSOR3NAg8MQDL6A+
0n9Q6+aB/00Jdka0hmWRVnruViZjiiBfGKmP3nIQ5Sy97pYmkdPH+5xQUDKXS0++
kZrL9gbeDBRfV9iISXTdKdAopZ6vzgMXxDixXBXBnE5cOlC6MXqFLAiEflL32sy6
FFq9bHHV4I8n7gOUhrD983ioehylZCAEMPddGZJk+Kdk/8D2OaX0RqJ4ILvqu3Sv
/Jvt3PQCBpQ8+ge79p4K8YAb9DO6IyF8gap5eT4Whsf5xXXkkF3A6tF/BdWvfEJV
/D/qWIqbIR+goLDrWKhwpUlN1YO0VPFIrmYYPxzlU5ByRxCYRGpycloN7Y+SBneE
p4oxmM/k8x0zkB8TDUgHwYWuCrYbU7k03H8bqEg34arLAEem/n6aBbKUDyA1xPgG
aqqr4cLSWW84GZd0lkSKoSzUbPdwhxAHoyeWm0dDRbEAx6X031c71ipkAUghNZ/n
yoCOvFtE8qW0bBBv2c6QCdOpIER8L2e7YxANcy0XTlqJBHcObguN8bOi7LFupn3t
+Pj2oXiwcM0PxWLBTd/9lpcazdk+BAFiIds3h4uNCeojSG3ol8ViKaOhlKzLuVkJ
2ZxtK/xsVSB455wNpI3ehOl72ohcZDtl5CL3qaCdDlnw0K/nVRsYzrBkgjSZR5yL
ZJVfzE0qtxhayaJw+J6O/l+yLjTRbLwEoOa5S4fmkTUeOZp+b3k+yYg6YyxbUSIr
RGi1HAZFigd4QgPD5gf3g7ksdFx+eSnpV/I5N2+QO5wUu14chwwumtns7tFgdU+Z
98QLvscPXMsZM0M6RaxLcLxYCoA9UH/mMjIxCt+/HJZ/AWEtSfvRb66nEsZ/lqNn
nH2Pxm9Qb5ok/JzwVx4mXL4fkP8gVqAyGRKCtREjtQgBh8/WKMR7a71tQ7iItt/e
gTs9ckC9OtTqJ7cddmbNcrhOnOEoQiQPkW4+5vrbJngKHDCgZ6GeovzSVCrxN5Xg
AsLg8bWUB9LC/8hn/dSHOnMaZ7KxgIp7NAbentuqen8O7pn6QT8jBE3R4VrQv/3e
MbniEFexEaVRdQ48zGhOwxnJjWUMvL/2t+j2bCncPHd3i9k73K+ITjn/tOnUOIfJ
er9LEQjXYMmE8DvZx9wMhrXC+sYw9afkGZr7+0bQNIv+42sZDlVxJdC3XqvepnFg
kzd37QIGHZ6u4qjs8ntgNxi/yN0xeWUdDvg2cgGfXGAALDwlQNG5LF0Cun3muh0n
ET7KI32p4e0oShJ/Jf0oxh5HkBrqLD2jVKNDl9pV4a6sxbu0Q3nXVyxqezUrGIex
6Hwm8EUSc21qM5U4xN6vwA/xd5LUwukoUEa6Wb0F8qEpiizZlwrv4E3bMdLJGGuL
ncpur9Ud6hLqnc9CgVFWwKw/QrM6tUiRJd9uh6M39a12DWntS8Xf0fRRYSHQfhvl
4ktaemk63WEuhAnLvj+6WawRFqYE9gCdH5hSYtc+mNeMBOYvJUfWRxk1Ye6Cy9Rz
4iC4Yj4jC/A2v51932I1pNv2ka7hAVxJ+nnT2l+nwGJ6/Ccr7iTMQFqwKSqQprO5
cg14EZLfYVgp276Dk8wKuF5zG4v/NKwnfG5jH33Jm+pfY2oY5gxP5AKgFmwVDt6Q
H15QXRKnDlmkffUjU03QZ+dUqVWK586dxiggHpOwfIpcYNx89c53BnSIAMKEfGBz
qUWbJ6kTXKuG3Ff+L8gLC5d6Knjv9pYFrsAARDxbHMSCV34Enww9CNws86cRzO48
qEOy9R44rm0EZ1eQXqXgSL5tyMxDn+gl/DKvamhHtIT5ANZQi9Uxrn+sqZVJ3O9P
pHRIGy/d3LbpAmYNRlKjseqhS/Ytz5M3ryF/JXlB5l6fca/XtWKwcIkMHn9Rw0xK
I36FY0+X34cs9lg+QniqzzWsNMMXIqOzhcO31tJ4ZXsRTWtfRIg5lWyIvjPYfTQH
lRSbILcdlKQkSntqHO5UAYPrUsHIzt1Lv3Man74FjJxvg6YeInleMWNQdNJZ5npm
bj7LFIOXmweJ+/8MDCFwuG59h0Rlz32AitPuBSsc97IgbyixCDBib5H2/i0qDIfY
c4AEsLv1Jl3MdEAJ90BPmDf+wmIpEvq4FgoPOkTXuU8Lup+APBiE8us1aF7uDA17
+eh8+33sCTUHvPxIjAnLqNffe6BN+UU3Ktt9/Ih/XAd4k9mI9k6+pAjBJhNEY2c1
pPrY5Wz2p6dSSAgg5++K49dgO3XgHSN9iLC3lTj22VWQmkjlT0qAnpR3luEOAPc9
Q7vo4tl9VNzT3/Jk6ziU1UX4UIlF5Qso3yWckfKNIhV3w4sR8/oKb2LFdL72tXh0
50PjRTKAp5vlsJVrhO34v/u/1YF9rGCOxItKRrNlOIrJ8lQrKXwgNgWG2Hyrc0vY
qJEWrDaORyxhkk+hz16tXxYcSJDxHr10XR9kQ8rpj+t9IRiFoZi0A6SGtduwtWJt
7O+N1n28e15PYccdbrHYARboIYV4Cgvp5NH6cgpazYoy+Jc8sWvszC6dWwbjpc0H
oIhlls78lHAL2fMKuzgiGN+rZyU3oIVYNrB1zwmBmJ29teWy0wegzbe0PcqR6HL4
R0Pc4NiMEHfZ3+zaIUfZfmXR7zl06KN44KG5m6oSQ5e8N4k+8eBH31ceqBdcOCjf
niPqvQA+1Yar+yeatufuWt0ps2v2F/q+GJmELHAHSidRHvXA0zwTcc+ZFm8VCPMn
DbpDUPcgxrCWxmPkGzP8sB7Q9tiWQOy2B59YmpXA9rfIb+dYDRzMZTuFD7KCvuNp
zM79nD5OK+VdoR7QtBgW8hxXNQNiVskHpPWZXmaJDsP9khoTjFzk8s6rY8CHXcYd
PrgBsszXvHn7+AejZiygalAD+VfuR6zPenikjGdbwJZtzzMYE3qC+nzBJfRqRcEu
tzcDuaoXkOzYXQcpRpSE52Y6lokaa4qktJNR+ktcIlbD9VU/EzqNi5kPwj+QDDnv
ilsuxSIy0WYVxi50ZkeSiN95/UB8gVRxM3zXxhDXb7rTl+YWjXjBLGhNvcuad09S
Wtx0tJaUdOqOsLjXLGWlj5GS1Zhdqray5nRYhimE7/CHln7WDfnLy4u6tHG+E9aQ
GbDIKmwWnhfmiyW6+RHPgL+2ZBQqb1TtIy6P1HxglafWmiAe9HUI1/YMq62xRPRJ
eWdpxJAtmNwsC4ty96xe7qDD+FUYZhBblt/6UyUYPNpA2NSBlEwZQ22glfDIAGPO
oxZeCd1Ouh/34BHxK5dqoQVe6yOVyj4IHqsLGcWlNo/tTgto98G8aqZz/sytBjs3
hlLzm/ySDVdu6+8x7frl5EUI0wKCnSwqJvohm0hgiKmmc9s2CnfUvrNoKjBy5Zxv
WL+Wd4Bv9J6wTj5NEqwZjosvXuHLi/qVeCmEsFxbcd351xYpF/tEkz2q/OsQe9tm
3uxPmtx03HUiBN9NXYLePMBVnltOwxu4jASGLJa+iUY5TKQgiPZbo4vr0HTBRnOt
850DsxiVRZShlWzHoLpNRbEY9+jMtHbcSGWkEVTN/PJqlsojIxA73Ctdoh0olQJ3
PNrvTFWctApZivdDismwWhEtTwgdwlLdDYBaPfcSsKznnIVaWy9bzwSn7UekYsjI
Q1Jwd8C3kIq+joN+qwD1wZ14amitZLoIRgIi24UiyEPvGeILhDPUXWEIzJxNQD8q
b4NZxURz2Zg1xNKbLVsLSWcxKimn8wjL0qlVSaqYut9rsEG6rYoyoKqALG4hWqEA
iaicTBq21pyJdBlo+8waiwfflAxTwpxMfjnWErbx5xYqfCI+z+M4i8kNxyR5fWBG
82mY8GD8buLlhXhTVMMVt0NxuaepmX3BD94/DzhXmaeDeZmNpm4UO3qCXnBiL5mC
TWgFGsl5xt8iGL28HdDXRhBHiaVVYfuTGFPBHmjUjfDfgFvl5rSfxxp/CVCasnNR
GBIFkSwiU0rJ+lPwkv1wdz8m1JW/jX0MKTrC9GuG1luVPVmWr4TlLCdfqOKDU1mL
FR6pdQBW31qiMhTJfAgXT/MgIwUZfEPCVc1iWKQzVLilhtyRGXLwQ1B2Oeiln3bb
+VHu5mtossJLoX8XLL48KLfo8s+Lf4KLdmxTRTxKy7U9mCZ/5xa5iFgOwI+KaZmI
YhiKhwAzxBt3LZ5ECQUXbzsb6No7nWafYzlr+Va48+OX3gJpDBCjhieGVGrh5ljp
fSxYkMsTqwLMXMoTYP3D+8yj2AYQcby1y/pCcoem53MKEvPe5T4GwMhHCD8J7MgT
BFbO7PPcmUzGQE3gW/xsoKUJYR3ru0LlVQv4MHwLSbOlOrYv3DRYOeHTcZglPH8R
jydKDxQmQj8Z1MMyTboWpso8lluUPJ6Bt2RUVXRoOmkFXKf+ArZi3970r9taNT92
+OWCXCfcBkmx5Sn8ZoK2/WbyCNaoaWJZSBsShJUYAnEk51rtOM9PUOrerh5Y+yGB
8wzhS9QITLh5TpIpVhm7VKUeChhcPjzOXl9UQxb/kKyFhr7SvzIHe0IDowxB46zM
hkgjW5guOZCS/Din+Cm2Cp1uYnQ8X/5dmGNTxkMTiWHbD6c5XN1+FQTTwEHaI81T
d72Fnfk94mqqatL6gGuSjShB9+8WWB9YPnaSYNk7CmpxdoKpDPdmgTjGg/kaviO3
IucsbGzkk5S3+WZBnGQrlPStgtRIqx21bHZgXF8SsoBb38Swj+AywxWt2OBWjAbI
47EBwFt170luKdPTHu95/jNipjd92hmD/sIoev4m48jPWUvvvJfuwXz7dImHTFm2
YEhlbKCHn+kKZy7yuAK5ZsGwMatrHiEpvePIm9VFUi7BBNcnru6sGG/lYETYjnet
pWuv4NyKb79UouZyv2DJXHa0GGtw0Nz1f183sPdljft0Z0fge0Rq/b41A0l2usKY
Hr1EAr0uNkbw9yvc6R7F/te3/fTvtlrAKeRxNHu352OTNgijzIG0tQMl9KX1DQqe
cpccoyEQLlnU3ZrZ3Yj2epLQ3wfxKvUqDz45RqWdFdugQHuvQ49GCCX5AQgAcnw4
Bof2YOOaP4FkdzmsZghwtVcIcmsQ3CjjKxo15r7NgR5MtKAdQCUP6V3a5cczKwrk
QZw/8Dj4uuk7jCZ8jbH56tnuCJ+wJZRU/RlH0U57zdwQ7F/LL4uErEwlaDRvkaVZ
u60aNWvSqpENkqI4Un1o2S9exafz8NHRds5wXyBDHxlEzvQ39FnhjqJGTgCNlwNF
q7oKNzwfr4eLJWkTXWKBFSMG5ktQdcghDI+oXiOeWFHRxTHqdJmfL3aWVKPx74JR
WDEGrIvvA+pNubCTpKlYfqk4vsoQD3T/hTkweP3T16PbRGfeq1gbQ9l2bu8G06Mo
5xgY5Bzb/GcX/CkFxrVVGPfB66rcoWf7ti28ZVD23vWRDST5wfgnMMWfq/XA3jpG
I2U0evHcwEzaGiSvHElIY8AW4pKV+o92pFFmT4OC5xyn6Fh7yfHb84e5O5yWh9te
nkFdOraJasmreq2HEAaTbBvqfrjVaOWoSG1KS1wurCoiIE5Q6b9cFEOXNDzdOglf
jrUTJmekIk1hKkoH1f1dgUmFotplHRtvcW964zROUttzHd/Yd6fa/AUi9ebRl4TB
vcRBscoe4YtvzrHYL5y1OHTbk6s5RZaePZOuqXEXv1siIR+vEcDFd/zz8ZWNta/4
KWRmEmwoPMeZdf1fi8GVaWHnQ83iYaC2YuQ3WYdphzcG7uZzFnIIPDtcXEfJSZbv
WKb/2aVWzdvGCySH+eMFDWo8WatfUNz/MdNrpNPklVKaj9K7OYRNRc0YkQeHbHLp
4NIqvBApiTix3Iq31R2MWrMHvXb4YGjNnb0Sh56AeuaXHYmRuSh8RpCEkaWRLSTA
Dx9b1y1e0oHqzkLb3HUUMq2jxG38+3xrUutsBeytEZbWHlmgEQs5x/eVi10zYXxP
3VPz9q/AkIcg4vxzNd7Rn41YAROJscZVlyDTNjbRcDSYeUJA/6GGD5ohuwRputms
GLucCaQmGILRIKvW0Ywni6M1o/mYmrBl5NYax/zj1N34s3XwGvBizHefW66Io2Hz
3d9d3kwCH0ss+1TZ4X45v2InPzRyxPS9skTrV3sXWQWYzvJiRu4iIxZsX0RmWWDp
1nZwhZylbdLvODiPiU5paxW+JzEegiMPaAE/ac9z7nuTU6pY5PMxYl7YH28QuPO8
PspREti15oOkK4UFVhx6rNXibUaReGfuNQ67UU2X0gXWIwvIWXuHvarueri2pr6b
8VjEr9PKF0J9vvsFYowrRrPxEu0fqcAQwwqjsiHIlHjnTXQRWNYDl2UOtv5v+1mt
GeLteu1gCzUMitkhErp+X699KTGXe7c3jqYBlhqMNa7HMTDjtA/CII4Qx7huaLaE
KIHjBbEsks/n4RNQmJgJJpB9raAbqTC5v5cL5Cma7zRb/6ZrGUrtDYRMwNIlLy6v
o1j5oYh08dHbyxeEIQmhWkxfshJYR2uKHrKY5+TPN7Z3BruZyrBhnrGH9wZqAw7x
hxv009mMy1tyO0aO8jmAvlzlf/TTmmz2dyFW/c0lMBegFfiIaoYjDSZYlp+VtErT
i9jPmgy7nSoyVV0QO4fFAGS/Rg0LcOj5AH2kWV9x3LUsf5BssP/NrVXQS8IfEsvy
DNtyiopASKHHBHvzhe20dKLa46hj4twN3a0DmDiXSxhmthwZh+CNjMeQ3y/gn23u
glzW7YzIfowqs2MQD4NUgkxlWfRLgySadBeMyq17zKUrzrb/ZnKPud8MCqqMpxVP
/XZnU6+j06X1psofgBnWmDY1kl66cWcIaxwX0881rrMNVXegcUz8NPzeCCLNF3vM
hk/58VaM7hNz24Zq57WCwW6g9QxbiBkxbVxg3h7ocr0EwmZdUcvjmQd81o8jnuDW
SRSf0jqdoaK8MDKJD87YegBqNk7Kte2JUPpY3GBlr3ggTSC/EXthYMRwCh0Bo9WN
6u5QK1kl9TsBHA1/uC53a54S1hrH7MyyIMsS+zOEFc5v4dBX0pXsGCmqFoPh6opy
PNOfnm4h1h5B48nXdlYoies+rueW6m/b56A6GaKqQ1YbWa7N7z52n2n5LrDngC7x
Xapw6FfmV9NU/ktmapxBJdb/F2ZczRuNRT2+I9l2N7+i/bew9OnYAJ5N5clFaHi1
zH9C7/YbUphhfy6F+WNk1qxAYYco+Zl1uPdYUmGUbM4GYyORBOfrKesn4hfFmRmH
MnCzOCfolampXQiPRLKvbe9sPblpkajYMPh0VoUgnGQWu35qScKBes9PhfNHE9wK
1TRC9n0vccuKPNxRcgEL+ZJ4v0V9UBvxwq2DgNQEqTbt+iwjNDkWMWwmbdSu06yQ
r7i3v/dMuroVmtPuWAqei0ta7cLG50nZ/WH7hyoL867thwcW5UsdOYR+JExILaCN
RfRDPd3bVaSqVoGuJbDvh1yzufT14KyPDYDkQ2YaRicwaU9BHb0NZuTukJLINAuG
IiDzWo8BR/s4txXOdwaMIoKpFJzDcQzxUYHNsmWOaqWih/K+vYz8Y0fJn4pz7JPV
v07VvaXRwQxo/Ue48XfFTbVGrZDUghsmvuBUwJPCTz5GrQ02bET4jWTDcJNcG3fE
JjwyiZ6k3fMvdUkJkAkG6Zq2TiijcSemTAPAI65x86uM6u00IJXVlQgJDFZTfPdi
mZt9x8QhUK7y1nxG4qXRdn/UrqiptwjTJQrdotoUR1oXR/KuOzsJaV01LD/Q4pmd
R+045keyHegn8Pdq1m2bW3hOdCQyvorEhDwySZxspiHP8Ipv35iwEpJnAtiPYNFn
6pToz+q05stlHYiYQ1AybskBOBS9rKwLTg90X22ulRauzMvwxd1BpM1Kg6uyn20B
AOE2s/G8aguiKidC8bcBFcrIjmEEmKa2J4cjRVdh6az+48v0ecixCfRz+iprCLjj
/7CugWL4hRYXHycpJoQtiQH8uSXs1pe/nlI9vXNAKL8+1Vl2Lsknp4UmPRoLG7Jg
JlelFWj7Fr8vH9Iq2f0Jl7bW/7L0gdvIGFtvBtiUOfuxt0Tban793wAjzUyO7N5z
YNrS4xkF9cMxD8TCVl6i8FA8lxWUr7bElXmdmXB4wWHvc1BFdnVd1JzfIM2wglDg
l6jzkYolVp37CiA/blfoD8KCPdOEoJIdqIFPYKfEhbYqi5r2QL0jBFRtjPe/LNcx
e7pBYay+BXCFMrqt8vSAti6rAbGINHPmHBYxTlWRfc7/lVXvPheHWoJ0gvFtE+mU
nmd31aYBUKgq7xyV1AS8AO3jtP/97kKuyvYBSqw8aVlcIxWi+WsOd9HIVzONFmM6
hsA9/qH2XEHc2CIoe+FUpYpomgDAW09mg3sbw1RbljqlcGZ3wnmJwNNWX/k4vP2z
UPYNEQgjbex8URRTe4mvAhKqgVSSq7DmMecJwqSozJWcEGN18syFpdw3oyTPCZi2
XHQ6WV9oQCyYgySDIoXNpK9qQma0+8vC8HmrjkN/d1aVlB8g+K9UIQpBNBJjPpPF
0uRXSaLf72i2IUkXOnEJ5ag9jL8KawJbmIh1dbZFQ8yzpD4FwMP14mKfZijF5ClA
B3OUbpUclEeJsIQnKwtDUExxPYf30CvMrU78nI3tZh5zCrh8AxD9Y3dPPnGqKcCZ
uUusnEjSKCaQmm8imZibXu7Y0meQJ3nYLG/olo2vpl4FUIYUbmX6aaVdTlUBxUVA
Tj5w00PmoutcxX9386tBjwT4Tl4xN3xoN6efrB7igBdNzyWtM4+44GaI4ZNvLT3q
wkcyyOreN92V/DfaC3XYXzYdZb4QL7LILE/wZ3Wk/vDPgNL7s8+cwWSD0fZ85OsW
X1yTfleWBrpwlcBweF+XIIoG7bhdaFSub/jRrh+AeiRV79ueNVQS8/q/unZlSqiL
K+x7knGZdx+MUy+bsa4uEzSPcmnRVFLq4Qy9oe4vjN07S//KW2Bh+y6WUfQ700QY
Nh6rCXvQJNH2T1Qr1L4nk6ROZ8lEn8zu4vzRGXwCxELpQoP6IeGUU5xRKPFvx0bC
O93ZQP6077sk+nCcmxt00oxjs6sfLJWR/bFrqDgjWDk1LnyfEman+RGN30rjHyiH
6oq8CxnoX9o0byBxXzLw0zJBKngmO61TMV1LVOhNHijINzex6TaP9296gjcvnE+5
UGpR81U4SbO+M3nZMPiPY0CbHSBP1t9Q8Jqm1REHq98PUcxzMZVIA0XwAgwlu1pp
a72rOK7FoViWLFJ6kD+LyS7BmE8wBdXxOfdjhZetg+7AjXtZNcIRf7GTuin7ZiWM
nlGqC4DF5fZfxjnFbHacu6gCxIVockZe+JzSyArNjFLcegsZrHRMEOx+s72u+T1G
jZOEqv71VA3Yr6I4x2T1cWJvCdJ7RSsRv6OljV/YKHvQE86c8xnawfLxpVYqIKpq
0N/HaynQIoBMHqjNLQYMiqFIAPyGEMPWY8MlobUtes65ZVgjITbibkiPOKWIQQlz
bLJB7qWr+Z+bQAs4tOWjxZcNWm5ABe1UxoB9Gmfu3W3gVNq9+BN8rkyH5FCHdDEs
QKQSZC57zT11MCpCtZnIjty7Qwg1HKhnOt0QxlQQlEERsdXc6i7U6yWrx9TRaBYg
PXrJIMxMdVNk4yw0jBbee70o+qc21/h8CRN0Nr2MG1BfEE4t5i/G+mQKbIrdC++8
Sskuz1U1taxzJexdFve8Xf/X0r/GUa7NhALWD12vV9irthE0Fww0NlFrAXHlow7I
lcMtfIoSpamYAMM4hAhnta9NgXu3Ttzlo0WzN7tVAB9hljcvDyHGQWmps87s1Kj7
K8myeXR1P+vb6tXwYUmbTU/kvot1+6WQvllrq6XfYTfjlrDFeMmFAhU0KzVMDG74
Om3vUtP31j9V1xMCj9DNN8qiPLDhn9xs/plFz5pg9ArfG7Xk4ZZwWVXAEHi8aDbT
z3RdQazayLMf4Vlhdi3C0jQbRQ8/4KR4rtwJVuL7oS7ymGWutYOHO2+5r7w01H43
7Y9KA2gXWHllTEIhrzOujxVS3hUcb1/KlpUj0uaNUSMxSeRnYiDd53r8We6vZzy1
C9FBWiiTj3wP+MyRm64f56+ycrWPV0s3M9clIYuEof7PyTg5Tsw650mSlgSCHyUq
JUSfwykbSG66VaVc79iBRIHZQOAB2D4TNHZAbhnrZYx77wwd7y/sE+2NXEYKhvMq
wFgBa6eMAJokBYTc71JBaNhWQG7vnNGP+f4srnQzC18ZvOSYONjp4j1uaa9QF5T7
GFEzNn6UqUjKfgaH3QOHcmvou3kWO0p4FvC+1jKOjQDVxt00GluTelCmpoLVw61S
mdpzTJZunjGgGYaLCmxAsWXrhrQlsUswRnpsVjgRNZbDRmgSHQm3rC/DCw7J5sLg
fw/Mc7GURPoc1j3eNuMonZkC79/VJHQD5MzWms8GFH0LO65DoKuQ0IOY8GdVM/OM
iQbro8bNJPJvdw7kH0FvecArqV7nnzTAZrrEdYjWZtYJrcSsCJ7ncqIDYnSxZKCa
L6fpzxLaiGs0Q8H88rcGKegtYNTyGbwSi6h8K1xgvU6SeDpeV3LSqefoawAMMrfy
0y6dptDrNPJKMXNfGjhdp6fVaswICtmLlGV6oPItLUWRXbENa3xNPjYS8Z+512uC
gSqVX/wb71MaD+oNbpKYnWxSLx8lk8x9lvsBAnbye+cfQJF7xiBrBHtB3b9rx1wy
aOk9IuBhndksKpnruqid59OdJisafW2B0AvL32hVBvKz/eXCzIqQA5DJMjrmApbB
IsC/QOs5COzRFAWHwQvg/lkofg/GiLTZMQVXaqSR8l7MFduDpNJgFYGa01tLQ+yP
pAS6tPNoq58LtO6jpGfw7vnd4uTQ3RTxlm9HwOGHe+ag1C3++D7fqWzpwaiQW7d3
O12J/8yHyvjcuftwnRpnjBmOzW3cr2xO68wviNuzUoGvt5qfab2sKyyxlJYoOikM
UtyUAdplDVfPa5MafVwYGcAauVAunUwrCMdx2Nh0I8tTd0Y10LjU6PTiY9/cwI4S
r9ObE994sR5ehVZs5SkLGDeEg5rXMb3kTxeagq9CTPf4JT9EJnHBVhT9hnMo9XGb
f66dG8RZaS9QcQ14RqPEaKOXlE1QuzSh3gQX5P3ZDTBjawWgHpUxdNLYBRDsKOAc
6nAxXVS4MDbMBHiyiaUHb9wznBIco8ZG+nlYO6y1VYHJYcM217nCj8KANPDDZdUv
6k5ALMOUx26r52Mmr3r8lqbRX+AGbrE9Iju+8SbD+cfiU7axHYE0knOp8+cqKTCt
mLVvQWz0xlmHEub8VCT3V4ghZv3EHorVd12tFvOIQzCBiazNbviJT1+ZQtWsWNuo
urKCpjisxEpJ26LQZ3dQig0H3lN30PQ0W1vgMB544G0o6kA4obKxK4EWzJ7cpJ6D
VSTUh7i4Cls/sGVhmgjMVUTXfzU4VMj0Z1CEOOJ87Tyhm+2MUCS+N50FFiXODkLM
eQdt/rbiqaJYAFEqR4jAw1LJzhcocE2bxY1zarR0uEryQzzhdZQR0J13zD++epPn
b0p8Mv4dFCndykeoe09pCQbrIUH4kcwZt//WLgHFu30pRrfkILT43r24RLlUqpR3
S7V0ZWFs/RsRq8LamWMwXg/zx6aYMiW/GolYETfc+D8RTY+a+nFAbu8DJMrB462H
q035DGT57Hha2/AxYyUnkvvL8Bm15+AeSK5nXorMFFzXUHyDAc2qfjj3g83hfAUO
vBMF7MYa+J2YBEIMuw4pwhzdu87YD6CXRhEYysdyO/e66pXMWiVLrgGJDgorLpmd
yrbw+RIL90AxZkY/bYc0aqaeRH5VrYFoPELo5/ThDd4ExD56MxMmGW7cM4FOEAZy
8GmNpG9N/rjvAXzmU5QERzAe0kRoQBV5xoQBH97FC1pSeActBGaqTMEqsk633vGJ
Y9mtQUV7TIJUp1DA2lYmjywb6jVbSfYn/7JDAA6UQeOh5YSm6uglaZa0a20EUdHJ
xWvWUTIlFdLbmfvGaB3PWlrnAVDK/KYQIBYDkfEOInR7j1dpUTIjifyl8zzQMUfa
QevsBrolIdDckCI7LsyOhegSl4kEVQkv/BaDBRkCwHm0Yq8s1CllzL+CHdYotyMF
XjbhxgbSXx+mOVLxHs6jxdemnM+QQGwcp6ie5Gr5S638dKmj6KxswBmBqsq8UNgM
KvneS/BC+XgMr/oLi7594agQBBHjdMpfXA3LV02t8hGXJVVB2Yb5HOhz9TlamTTa
2/t16RD/JJUYX+pRK/PiH3LZunJpOu/zPevsQOqrKY/D0v9x2YMy0t+YUV3qTyrE
w/PuiZRHF2UhdrtK3Y9F3e36BqkGoDjvPf387ebR8BDduv1O28heZYGhKBwMYyPh
5GeYzm8QfbIWaS2QeC7kkJACzVn3SL4Lso9Io3jpGWCNpdaw4UcV0ozh3P4Jqu8/
SBz0i20rGQMBd+7XknAdW92KvVjA5+FVBDwSI14k++sdx50YcPwdCsfYJ3H8LU1Y
fsH3i0SHOe21OwIOeM8dYNL11FmK+mwGL7OyVplefMZpF9hKEGrfb2iKnQGVL94Z
M2DKYVYBQryTWDW5RZVnSU6tk4IoqNEYQs/8RSS1Cf4Tsys3q7j41oItyHMMgPZa
v7BFRGDv8QTSaIoZLEcAV56EK0R3/DblpBfk0slH7pdgR+nPiYIi1YR91CFvXsHu
71sOEH/2dIMxa6yDGR7FhYuGfdpu5JDpe3h5Rm2zR7RgQ/Haw2fE02sOTjaQnCjd
+tm34nRhcGSYDHODeFu/xqFwLBV8IYkVZUEbm0xm3oZE9Zr59XeFLQgMB/Wzw1kv
pG90WUjp/OMpWnY/6v3j7U5YhVSyZ6NtjkqGzaQ5qv8kjl196SWblbgqm2qtFgpk
1ibv8s58CAq0hZERWRSdalnwisnC94SlvE4Eq0xIqwRVQ70BBmPModmHawtS7B/2
EFI3z+5TZ6dyXE3yo3BY3s73jmikegY6IAmnfamx0tUIaKi/H3FghOhe6eL0kkcT
k3h2nmFzIiUB+zzBE7yBp4L3kf1HsV6mNoxOTo8iX2fWvQHOQ9kIhv5zIiF92aoZ
Qt95lDT9MdOwMnPEoZCtxmIqPaMEcyFj9QIirVljgOTjn45Sc+w0n2zW3Adt2NEo
MiNjWOHveCUnwyjWwj3NFy7q+gX4DAgIWqmIikONCPGuMGhDF+KaUGfEbR2w5IIz
25q7YTV9QWk42zDALfX00y0EVjzvwHCoTaPYgC488D7fHPKodYhzSqhafSj/5IND
d7Hg4nDdU7uix98pJ+V5ey47nOUjxTkbRwzdDhqYUhDbn/Ke54gFzbkSrxsCxHaa
/RodR9HM7MFgZSPuxtFo/T6YnRxJSVG1FWzT4bxjfLJTsFX/lRZJ1WnkJrmvb7Zk
3J12tUav1lZ8vpSOZIf+hYiiU8dFHxyFKa5vX/i+WFcD9dV8SR5FVH5Ht2EieaTs
sIPdNRrDt9XmiwWoRUWZY88nBW+YbFI5V+rAgReYKfxxU2vno0dG967JDF9lVgSs
kD/nJ0tG36FxWebNt6CGWZ3OHgaYwbJfqjS5JWN4SVQeHU7TB6yRUtG7FD5lw1YH
ZKM1nvInZD2s39YehOjKTmvMWGwInWbwcKSRnoWvLBM6wc72zFn3AX8JzjbS7K6p
h/hfdMxtMthso8g+V03uQj77tGRGVXc5CSiqlXc8OU1ehaHiILIQxfs+u02At0bj
X5qesJjURNjVtqwP5OsAGZcJwQ15Fx0Uuol2QxGJeHiGMW5p03dR0vWlpAmL+Z//
DCTFxien3uPi8YUukfD75RT3NERjyz0U15j7zZrrhi3atm1L+5tbcNUCFhRbStoY
ovNYl7dFYcNqWtetPabC2Jsd7eNXO7zdAEApAdF12XuvOTVAY9O9SBGW/lDfOcUh
+ARMdJaQEl77N/kizTSZbPlVfTiodLJYRP08mRC0iVUp9+HO35rRJTa2IqVed21b
I1iIul15aWaVIktwDpDrmIB+UexnZso3zpUXA+u1SpRrkZh9Ux0BcbXDiDtlZfbA
9CeF2eGSTYz9E6U8L15GlQqcaQyXczH+OgPNKYJ2DPaL7Eu2Xqm8YR7ZXoiohXqo
TAv4MrmRZ6qLHvkdJqjtxhsaIEg1mfOULup5X1ZuqHyMgOnxzgnS+wZqxjgtSXqO
r1xr62ASvb+3CMr7NavL5YIDgYrSY6kb0wz6yYcxrXdomZ6ICTVM4ZnGRPwGeUHF
N4p3qX445dmM3VHIQ3YGfxrcWaZfCANKOT3uE15AHAEERM72ASd44WBVLQLctr8q
J6Vzfq41YSzg7993Lune69w5Ub97LU3HXbYFyCHhnDl5nLjRLkOtjkBk6E//h/42
ViVFrS/XayN+YA4h7uEU0JMQXx+RGmxSr237TMon/swxuVV/zp1MngfRXb0VjUXq
a22OYsEu8RYLf97gQU9QcdhpLAJLG9k8pSHNhLJLPBJow7+BXgaWUbcQ5a6kBled
Zl39unl4W31J6xWSg6fIOPtbgQxQ7V/yU41k3lcb4G4gKEbsaGuiXo34/W89Gohp
dO+43IosgEIyGwPsSDvX8IIj3ux8lu6rB6I5OGkUG/l3AxVrLGp4Ed5ak24O8KEa
pZ4NuRKUDQx0ndpU95lQwiZ8x4KFU7DM4irvJeVnhuG/qfeYG+yIPoZKEnp5Ee/7
NWp+4eQ1eNA4LL5X3+6vascUPdEZ4Gj3cy2ij7qstsP7qj8eBh2E7PcJAEhTK9RG
paf6eV5yoZIGD3PL8q1DMUjoW2rR6Oy58TPfV0/IV+E0QHru1wTLPOS4FJZ5ODcU
Pk4zfzOl2ub9BrzHYQTdhAvEJqjqpLLhIynn3DIJqu3m45pCRcoKUL6liPjp6HyE
CKEUrpB6Nh1+9CZ9ECQe4cpUawtAfQ1rZa/63GHmj+0ZrJGC4BStUYghdzCftu3Y
K0C5fX0c/7QmmCY8ma9UGOBn80WvnyDPphkC+h1a14zUBL+8x4J8PZCWEE0t2Cjn
pxzIOcRkT83pF9ee6Gh61Bg9vWE6bsFwX+fkopQHVvYlEip9bkLRL0jGnhMamZwp
Gh5mqfyykGZjz8vq7KmB4fTdruHhD/TcRhMrJ0Jm577Pg+xZFVyYp8yknbaHxwc0
Qwb53udgYnNn74RhzR+1N/unqQUhUj3LZBnjU2AlA5PxMpaZCQFNpnSM9XtD7Iot
WKEqq84uDfWdByigktOHXo2/vJfINcJb+coT6eB7n6RwHs6ccoLiWXxjLZeRpmhz
WZg3hoUMPyDc+1d/AXkyRu9bZxMwXgAfiQjsBg2TOkTPH6h+blEqMilqQcXG7ofI
1bO0wbgKL0Mmi17pf0j3WZKo7GX1xI5MhrteM6V9Ivwen9Cpz3H1gXUMxZx2/4OH
mTMef7UDyiFBbu2VqsPHI0HSMh64Ir4z1xzU7pBOxSkGmvR2dteR9GQjHUvvIe0Q
+pxL2bO80qNI0vAMSag61Sj/q+VIm6wezyUGP1FDTh+p4SYgFBvLQCfI/bLD6Gom
pgx2CeoUjy4680MiKfTZE2nXWla4IvJxhw6quFf5mt0L/+/0F1U5LwJ5WtfvyRlN
hxG9RZiLOFJbQjP4hE0vcnxM7yTLZnvWvJdDBluNSDwmdo+f8ppvrR/ik2owRWRW
qbxHRHURkNiOTrYcfC93A6xBiN56cG9gEUGr8138kNuiu6DrFCP7WhIaOaZoBI3f
RcXcQdM5mWAiGj2wYbUDf+zFDpu+QyE50Xc3haRKHj3X5W1/gOD/1Pw9/1ESLMUh
rPgropnIb52ljb3Edxb+vkDg73f/WvP1ZFA0vHXiFERHD2juV6UJn9r5DNciaX5n
bM9+Jx94AM2mRMH48WpDfwKSODrw8tAqnrwWKU4HfT9p6kzK1hRY8zd8+//bfHGV
rKO1uStiqB1XM2sNJBHjAnbyotjPUMT3IngRNqhFQh6B3+xHmFe3FWg84zDh3kdm
SY1PsgJQpbqyBAFeR30FGIavPzijnwt3fZq6UipoM+0Av+vJWDx8jvKkq1e2Mi+w
AOq/Fq9wJp3/F69oxlFpxrWi6MjBQD0Lv52j/rERqKwsqJDmxn3cOy6ran5TM2ad
tr+zietJzQj1xh90g1M84TjCytUf/WSkdD0PFo/M+frlLR+HdpcY6GRSAgwvSGr2
WVsi0GbLVm0k+7XjKIV1VmgfVtE/d29vYRLtjsVcTbgGAchiXs6vpBM0qhHIXCu/
wtXCUfJGC3O6EuKx4hCwl3CCl//Jo1njOddxhAz0bOTkxy6oq7VBSwL2bAbz2UW/
UUaoq1rPmqfHYu352ulyxt+zqhoUcRVfR5vLVnPTfPAIsRhVsNJ7wDGyKIrCqVK7
a32FJc8zCaJ6gRHoEuTgaX9yP7BqzyxSlrONAAolzogbDWZ0NeFZfR85F+4a1Z1N
UkHOcHLYCmym6UldAv9Qf2CUjAutGvoPjl70rT+mJA+lWgGHD4QvwFrVR3/YSgYv
ZIwxymp1qs7EEWdrvLVbDMoOxR3yqEqcz1aHVQCFI2zTemY2MVYFo7SsBal2wiek
5uQFcrhwDMrxDedfFeP8eKERd9re2aoiJLz+8oBHVQotOKybTxaZsBvLkSYqHTLF
JEQdbqac3qc31c6EHT52P/2OKSV097HEk4sUy2gAphFvi9Poadg5+HVfYzlbAbSc
8RYxt5xyu404g8WptuISqdZHg6a8JDUKOL9E8LzkYB4XA1rKC79F7Zuq96veMJ3N
SZov6cx1cF7NypyGb5jGfb7oSfqadWe01gLhYltHVbG+dQ14SxJ9FnPlY4WyzxKQ
l4Ql+pdUKynaXqilZmN5r+FqF+ClYXzV2zlvPEywMfm0M5YOG+sRCLI4XlV/9ApL
qjqH2TKX8A46j855v521qTcZY3B0Mg2MZdcuqMCT0uaMeOGks/rOk1f94ahaWSdg
sEVbF6O39rAICavLUEmYNYdpPSRCBRnpMtPCV0BQnzypF5nGnsbwSbQeiufwrutr
XXqOsd5xr0vSne6rMU3NxnpHnPOYhaDKS9KnSOJ4UBhCW8zM/3NafysA+l8VVokx
XStxS3Nmlxr83Z9+TarouXg4xauwrloPK8OALPcrg9auXgQBgN719C86d/quKfn/
r6HP7EZJfEOhHmjMGWF0JeP8EOUWenp9MXgybMOwiR9P5xc3glnuuJcKvWs1uk2E
32uqEtvBGzflO6Z+pRqmIM1RzX0c3ZiOrsrXzQmEpA8muVvw78XfnvcYhi197pBd
gi9iO91Xfl0jYEpd91YzGCvDtRggP9rb4BITxY+/IjHGG1soJ+YxCAgFr+eio5J4
pt4jOaMhB+z3Ic04ayqfn1sH/hOr/VpsC+ogCuLpetvgpAHgvdMBiodd0vaBBxjG
0S/bILR1g6/t+3n/YeBvSNlq6nS+ujeDYg9Ym8UmNJp6eoAyPG1xijPiWxl6C5SX
nrQ+CrgGagV155pWbL1cxGr6fr7lTeGtw7dXenQ16iN8rFhjZ17KYAdUjAO5u/Zk
8tgcwgX2jWMBexj5Qwb/sd3UvmZU4J3p5GjugFU/hhNDQ6WwTHjFaKBFTm7EuzsZ
9ZRx422xpVTOa3PYJ+k2VjMhUVm8++myUKIgrCrvjkzpJ0R5nebCpLQTS69VxVnl
2u3cThIrTmt/IhJXrW9Bit8aeg8d9/l/OhrEH1ZCSqJfW1qzl3jXtJMpfjR6QJpO
u0FQcU/5IwBhZ/bDL4z2wmwbCmA27AqNduq36AsaI/GHEWJZMnQi42VyO9emX2zB
NM7v3AfYCMx3y547szfN3+2uUVMaafX3sUfuR2Un5x8KcO+P0kli4LVJ2Cbs96nz
ft6Fe5WX9bRy4BTKOWB87ttUhgTd4b+E/PHr5ki+yZub7HdqVvzXmYCeuq9552bp
2IbFev9hIIRz6JEnwtacqDOp9ULlLwaRb2+iWw1TZFvX022YCZjiryu6B5TlE4oP
94phlOsyeiGGLgTcgHzBazPxJrK60YEUBhfoDcGMiQn6vQnjVAAtfNvKPzd2Dy0D
4y++t5niFVnPVSAy9CG5m0rnnXaJAZBZXiEOsFaZY5zCA8MurHnxve4wRvxX70QV
UIj+DlXBfiTe1Bzzmfm7F5Wtuao+wJOl+H9Yh45pcnn2DIpZfzqgsSFPopuaC10E
oCSLkCgBuQAJr0wsKa4oD6skNSy2VBSEHqPLY3q2edr47aKikw1XrHyXb6M+bBeT
swhEmEF9/jvow+Ia6BMMWe1y4tmtaLjo2e0TNxjX3D7z/+aNWu3Kribk5X4+X33U
k5tbFleznW3wzYEFe8BrVjNAud367+BAod1RlfeS7QpD7TfVrTCHqSL+8qc7BMqk
nAknZqF9/4IDl+SbygXugNyNFySZ+n3K002m9bxwYhbDDdHvGd37xfF8gvNuNF9s
QS7IW+qMvfv6NtFD5B952wDqnUQGiBqpv8HgxcXPwY0al/vir5niMxGeSH7KTsQy
3dxKkcEKPW1hMTMTpvxzLtksCeAers3YI3EPhXFZubTFXOxCIi5sWRH2SR2jdO3k
HZkjX/0Esm/q2inGH9Kz94AINXf7kPQj3Fqnfss6va0yjfVkvqIxJUDi7lpcDABb
uSVQd7sKexNHKKlhM3C9hzylsRLp+AZaJUk6LYXmoe0OK+ZGnkU9NLRy9TDfLTbb
VLtdczxetb5NzmDYyUnDQafnyvaiP4pkid0BYcz8EalDRiO46gnsyZ9/ck4WF2sf
gvXRupU/ECkkCYCxT69OvCLOaNKjP8E+PKKHSF8+zqsN39tkuYBURNa5tCULbQbY
c1I0441MdMxt+ht7yfmzbR5QAzw2vAjK04eJC4BstYk1hQQ6rcLgZbJ6+Vaq3lsD
MT4sUDyfsFyLo5NFXcFkCkZzji3lR47KCRFB0IpMtlLCUyTFMWqIYLKEINSOnc2N
RU+q02/j7WAuCWxUKwNhD6Aca6JBPGUE62M4DAm1FrgxkccjWt9YpniZ0EUTQB4z
UalGro8lr3+j5FD9FU8K/FR/Z7Y3YFuUQi12G3Zo8C0DOPTBBFyDLalCzb5knauS
3TCdgYYUdKjxyxCANj4XIjfjD8sNrQMqw314S8ysBqpSYHrvtvcM9Et08KMkVFQT
NrrCG8rXiioBq2wWr21yScYMrTUDh9z7qHpW4s4XZRRgZD5JCM6DLgwIcTGEju8w
/EVWpUrFm6J/Rn6lBKp57t5ski4y3Qq7Dmjqtjik9Xzq5gqOSkx9qCAHRcGBMDP9
Ap2+RH+L3My9S+9Lfboa8MIzm+v+D2TZeduXRjGH7MjS89Di3tAEJFaUr0lajRCI
MTDJEcj344Zn2w/xWoXbhtE4dqKwzjOhD3lOA8PWe2YFAteqUGmZ90exi4Tfyl+r
3S/zgyEbOYvQmKwP4tvpP73hNY1ouRQzdhZ4l1q7dCd/K5R3GqytyLoG7A1KG5Uy
u3C3KSRx/qSiy7j/zjpLYmILTJcKgh+qeWyNPWNh+cqYhxPI8vT1NiuZTNxD6vC8
SESkiSE+k3hmHYhroJ0FesyY5OUkGw7/kcrGjxAbICXLVyWI21yNIfg7UR0EHYys
ui39ttKm3VKkaOXYASj5TURCFhu5QKA5mFxFXcjI5owV8I2wffcBDSRYMDpFDxCt
bcHdHcC65VFISbmkyfjZugLrpGAXcskPPpKM+F8a3Ezqwd/lJ8NtqeXqfAvlIYug
s0l0rrlJWRsv87RQ1KS7UCgsXC2LmbAH9lsLpniWBGF7tneLKnsaVKd0n2F/+bUs
Vk1J4+9GJj2qRpYgFcjdX63WFPCjl4J1TALn23fel/e+qFEBLx/CmALjsEwLmSc0
2QNtdbmMPkFEVehAyP9iBUlNmZ6FW2dQjIORXQRKp0G9GUwqksd5YzPG+2B7bTfm
EU6l1jU4zghO+ZF1VyBnUDHZYxHgnMDvrYbzuajttAo/tlChY/pjTrQlOZBgqmQa
dwkWF5aPSuFWTiSmK1dBpNJwmUBtayOk3bi5jN2GnGplSRLsAksblc6mC6QBWT+/
MrRNvnE0zEEouXA26cyRAQBZFnVFN4093wP1IiOnHTEccFg5Fx1fahodlm4Bs94X
crbISyCcZPaoZ6ATe+pmsT2CdptqNv1aNRLd6VXDIL9V9nIjGn4TrkREFd6+5UK3
Tv/zzxBAsyML1YJbv+T2U/voptS6mkYrnI+puCi6DMj3Exb1rhCuq8y1RVAkyiuM
8r2gwc44XpRZQ6EaACj5VXiHydV3AYp7JEVZSFblJnDpq6A3STkCf+sdtsuiz5GD
K+E9WhUzISpA6fooT6qTg203CsfXwKpJNEONed4H3DQ+J678u27p6S0T/44RZbdD
i0p2VFRjw2d1XeEBqAR268AE1E2xxDUT1dYwPzhxSqOwONdfNFi1VQ1nXAYTEsTd
O0OTgfRVR2MCcfrU/W1b0mofHwQplGvF9CHdMvWBPRuoIXzhaMN/1PvnWNuP7Bhn
nEJGHkfHnWt5ryIqI8+6Wl/aBsHH5lj6JByjF3+xs/8C5lKu05fHpAJJ13OdvJOw
YT4zwJm45XwrrcsGXZCNijSjCW5wRA/vCZTMcmzlUZZxR078NqybkVd9Qqq3IpB8
EdoadgSYR2HTHor7KnskUL73DZPUYQR4vGcy3JIcr0yfPGUsWOnaxcmsdHiUwvDa
d6qpHEhAJyOemGFzs7OAAscHgbX/eAcH/94047xpC+t7e02x6nLO7/UIR92uWwSE
PI9HVQM8ZNY6rbKFm0PxZ8fBDzbgTDyezMgew2gVDb0X3pFsnr9BUxnkE2j4qujo
gIBn/KTD0QlMcgxsgsmZnW2lecjQWo2zBGDq1/wC05e8S1U7Kw5g7GQC5T8H1JTO
bORQCmCt6CBYZwUOPzp408TSwOBo8U/YEf8dF9WrqA6D+KDk/I2l9YNE+frY9Hx2
vJsU95CpU5GhYBq+BbZN1/MeUP/RXoGJ+onrVFBtrJt+OGwqQQjfbC2VIhrH6mW7
fjcrUKr9LWptA5xMBP9Wtz3kFEWOPLuoyen3TSxO5iM2WlrYa8uAz+Y761Bk5qwR
a6LUPKja/1eq/h6Y0fqXyI9KV23T6zLod/JScKTGe1bYngYwj6eE98o24DPg05ON
w4A9Q+S09VSZkRNTt7BFG+zo2VnCEWo0VT+mgfXb4iF7ymxLUHkebYJ87Z7Sw7VP
mYyxK1GpcvMmc61C0AxhbhZD3jYGyAcdj9IYoqvkmtKcend6sYvUQF8V34qVjgeZ
6m2bwAuWm3EIsdEfbvhHSzn5K+66BJZYvi1ais28De0zlS3KdmGDoavCFWptG+et
W07M+9xxig/naeB8FU1DqUR2vxefYQVmPua8LNNZoxXzFoq5VjCTtJkvzLSn4IbJ
dpCwFVwyqL3Kof8urtGwrI0kdoF0H7ZQkGlirJCflCNcoNGxc/Rk5z68+Z1iAVq+
a0Dn98AzsOMUfbRxWxVb4UW3wHRSaNtH9EwitaYwgM4xc8tCfZhcwtepc+XvJAUZ
pmyoYcoOOzSUkgWNsLYnIzUvGGuJy4krJvQrmpAksuwfZ8DZ5F3JPkCw+/2YIKFm
Iii2qANaXzjS/qT4Sr0t4YG0TJJ0b9PkHDO4gQ/3hnQ+xI7D5HnwGl1VvZpMHD+D
VZ9XhSPyV5Sh6byFDCCPEvJq2mRMlXzEhuVKnHAU/8d76VuM9h4o0znoY0rVrTUj
lpE+8txSEyOHQhwyuEIO8e2OBxGPhdaC2H1QJVOBM960xxWp+qTtGNxWYnaSz/CT
n9hfCMs9lcS+Evnlbukz+wBLgySSPRoKDpYppwzI7kzEqKHmZCySxGto2TGSBBkQ
WgexNkk0xzpcnX74y8eiF07vnu76e71iV9FgA6pwYPzQe4I1sXkUb22xczvHpEHK
vU/DeNLyjsj13uqo0KAZb8qgYHrZZhzR4ruEhB/oNPwVIiBQ6azh6HxxzGlisghE
ua3FS+ZKXcU/ski2givXP0px7J8Kmq4AuERlXa1N2qY1sNxGad0u7uC0rWD2xr0W
4rP3DTp2fE2LR/LSG0P18ICnFQgf9VBnUO48cv58uZxCZ5Dw6usmc4eqOaBkoU3J
VEdASE9Ld1dDytP25YWsG/4IVE3JSp0WVC3gKx3Z91+3LqSkeJ0dQM2PrCTfvBTw
cEepIxEyvKuNe+EENQ8H1nja1gFdHgQlp8DxNai0NGnFlhMIPNiRzuULPEDcNlmi
2Zdm7/w5XhNUYb2JmvRPh54q85NNIOSiRj+IEUpK3s/42G5GbWajn41fmM3RxXbO
Bu2ZP+GZhMnvqXhSskGOB6UCqqqnBdpI99dex5jMGfAIzDfQu3eiTqd7p5CeqGQs
/7gooLQ+LUZg94hvtLEMVxje6NpCChdoB+2+Kjak5OT0VoYM868TTos6um9w8462
Ux6IFVgSo07cUuQ0gPQaqLrb9enW4V2hFfcD14ZSjpqqkHPMKy5hdbbHOgGY3Ndx
8+p+UgoslcEgQK4fa3IdvUmQkJdvco7CMZXHdICdGn9bK0kldoLFVx4tiloUIY5u
KI9xg3sO8giMf0D9+PBqHlC7AEg+BeD7DQtbU7q2UWaD/aabWyk+HsOX0Kagx2p5
B6N9EMGL933x5Pix6ekbSzjDRtJZz+evrXDnSUcox+bqT9ssNQq6GmFV+756vJyA
eVz7S4+yyScAnjcorkQrHVj68gx87y1Omeki4abpigztEHcZDfnDqbtqhNTLyyPA
W+R5NKeyTX2cFCKtoIFdz76VhzW0Z4M7nQErJ5zIo1PHlLUZJ/RLuTIvieaobakN
GYfCYW7vwUJjB47gfzNIoBKrsohyD/g3wBsU6Nyy2Y8FKKPUYTYLuRQBsBM23qmG
R//Yjjx6iuYrE73zLJ/yIGZjc64rY+FwXlipv13mtSoUrlCYbtseE446ldpmHT0+
SMBsBe9hfAczf2CKaRY91PkMc0oMhpj1q3e0NsyieBK51VknAziFkG+tRUt3sf17
e8bI9SgjzMcoXU/VBwY9IN0oKb/iJUwLdhaowEQxInrnckst9pB1FAIbFyWb1KGb
ubDJKOguja/vjo2MA0TbGHW+m5vd6UkseihCir4Fux2yDO8s6xmOI7YF5Dnclnm5
oanTegARhi5pOY1XfY44S5+oDXBqlGrP+ybr0NAPidEvupreiCiHXjf8Ku4K/3EA
/zjitwWS/S1gEx7LtpdxLq3hUXYOe9BVYBlT3DtkyEDTIJ3zzugw9QaY3Ym+H0hR
BU453DwEJdn0h/h87WxwtkQjaBTCv44nkaMxbP4+jtN52QKs/J61/ullFJjPxdvV
QOg5eJuH+Tob26f8ZWI7PZqxf21tYOFlPLKLV6x5Njj5mBVXEtiR2xrww6ivRa2a
SNd7djgSlhDzYpfiQc+yE7D9Ic61npVSYGSMmMa12PnRHz9o4pHfuruUKUm58owV
r5l2RqryQJMNpZ2QYK8KAbO+agl2UmTJG1TD0gv/aXlwda2MEI1Xtw2ecdi2+h+4
s2G5iLt60FD7vuUVcKKBCoLSRUFUO5U0UqGLgu2LcbhsM1UCJdhiz+4UJvPslKOj
Z/kXzY5FfjQQnfm3qZeKOLoaVjFeYKA5EdLTpUoK6FDrao5a2lqyKd4MDKLjy20P
c4OfcEwJmsiYZ/TtGGGxqkXzgv1cQfkLk/8X2ID7uo6+LusMI/i55l06JEdqZ73M
PYut+v3WKoOmLLWehgovBQmgA+cOuKD9I5xLSVaA7WsmmfKMvMo3gM4P/ztuccuK
3OEdtyxyODVppF3GCCulDSTOxXojOxU3HRerRcuoIWZ9/w9gKy3HHa62q/unS4FV
IP3VnxBaScxiYL8gZ+ugmYX9N+Qjp7Wtn0yU9+vEDloywMO/Ik2bTcK4l7Llqsw+
eW1SPQiYHp5KTjj6iUSil6VwNWZFXzpoAvubyl9gm78TeVa2tnZpdn2ni9+/m6Am
+oVXxMser7Bmnzlv+Ok7XmRRQI938k/TJPBtSEpOECNxbVZmfMftHkthxan7PPtF
H5+Yj1UNxdGo4t6RMmLVGiYRhIAwbCHEcK7T+XCSzEd4OzTAcKWaXQnVX/PUD6Pj
aO+F5yNlaHlvGPDPWfEg9ZZ3XMlF8zV3YDGsEgu7KQlNOEy+jJ4hSV/3jpd3CJyb
7J/Si2oLaMKvHc2PC3ZaQgGDfuAntX+SKPK7+UC2mZxd2hXk6hTQZGFvyeuHV2E0
SdvcJhUbyxGf8AIoqcHC4k1uBj8jcQ81Tgoeav7wzno45GebeFeqGeuFV5aGFikT
/r2LyGHtdeP947XHa535ZLDA6uZp6xNwPLcfaj6A9flHMgaG4CpBI3QnmCWy/k9E
UkYStuOOQc1j+AMX5wR7nSJwXp4R/a7u1OkdMQkK53tH0JsKg6YsAcmMIPV/TD1j
VPfwbKlD2lVbzflYLJeASlW+6R0bsdo2A4erLr9RnRdr7N8zY1IAqAs2gck9aNQj
Z6WMQdDa3WGof194ZF2WZiOPCWIz3J0Rj2j/GfT/EVsxkJEzzVp0tKumKW7VeVb9
/kYD24lSpPQds31O8pjr9+W8uWH/yzbKTHiHiPnOzrI9Mu6O7NfDorj6cA4dKdOY
byy6iK7KWnSOek/i3DafwBT+se3G8Srdujh4VHBHRjHD96mc4o+0v7XvJiECiHlQ
cGjMzWEgYbwW+8w1Id75y8nMMGaMykONCRB1NBVKqcB8SUJPjFm1JYrVhK1t4Mnt
aTfj9PV3ouiSVIl2nHx/mBonlQtvO5/9xSBPjtOwPZOfFVQagc/YyIrVadkiuBGF
osxJQ841Obf+eX0TtF4PbZ1Fh9wQfoH67/AL2LXcFPWApyV2pcrcaAviC1P7bTT/
6mpgrTU03H+UKA/CJcUONZP2QobU2Pwk1c/aAKY+FC42k/eK8yzK/NRTfGRmroXg
ygqGcleMRqdiAeXrHc0hSMPdJELL2yq6jQlAp/MtKIVH/y0Hc8QnYHMGZHj3NUWw
zD8WAsjnb4DeHvMMWGo15NkXIiixQL0AdQgD1uEwknMiP50jSNkVWzjJBrur8ZUd
y/Ys6mT5gRgmSiD1vONjmMgpi2M5bYYK63qW03hHNoUKEo/CoOTLCv0LRJ8S3QiH
3JYjlPUNCY2XzQdk8nwQJxlQbl6mw8TxgwIBc2m1MOOx76UsT68CeHAL6oWGKC21
Va1xq7FlSPFNQ7+gSTdr9mA+biJtWe6kuNMrTv0rkV9WvuvjM5V3uNlqiNiRVq3D
zOidC8MbuFc9DPXF7gO+u7Zchq7t6ACmYq+uxGJqbLiWOR6Mbc5emWsQLplifDZC
HE0VwjiZMLgrSNVnL91Nh8LMPeOG7zSypMhecuiYrfrIsdwiwbK9LOvWqf9AIoQ1
wfvA/1WbfrzKow4jzmUBKWLkqiLbnqCa28XG7GBXNyGkvaa3IRcTzjyWof/KjBrs
J1TazIMxoZ8UY7+qsOIIJ3PJMTt9WFcmDyl4cyI4bEYvmWFU40vsZBrdKo2ZGUKA
vt4SETcXLLy47FHS+kC7yWYKHxi8eEAAGqrA7m3Jq4JIU642INeNaMEWqbu1v5bd
PlKuikHgJPrUa4eM24Oc8PPMV+IrDcoQ0Iz9W8XNE2YW47JT3R1Km4ZryG8wCJXj
ivDP3WBVkFtadGiRtaZHAW41FqtWkPnldd9lKNbaQyYiO9tMAkbStI47rIP93WCS
16k1Tmsb+Oucjvlvk90a6maTVltYdyOxMJD0ZQL53NqSn1QUNhUaMoAyDxatzhAt
QQosEbQtFo9YScG8ZRWom0JO43azcXcXH0uufeiJYW87lQhnkGeP5qIwRtPipBvx
AiDwBhWxZly07iocfyToV1rtPmB/focaNSpYq/hTsdyGYp4zV79qA2QQ1yPsxLf1
EzRfrsg30Wn5DWOOqMm2UjEO9gZIigh+PdUCnYQey7s6VuIJVAu5s3oglv5lnlqw
CXIsPRFJ7qLEokEuwgPRj5EixfCesbPSGY4TPWv4Tbl3pdoVhGrpeNyn+yoF3Fk0
R52W+2SMahbyET8wYLWgV/n+6ZeMJ/wpqV2p6GkbLrZeqtgLSpFfqIFysm0vmet9
y941hMX7ifN5K9K65Ac5DqqR64pojvGA4qCD36w8uQnov2EbsEL9zOSd87m5TBVu
fvYnPHC2wKMQEZ8pDsuYLmkch0kij2wVt0cpvaAFiwW6vPK02zyYZCphzoxJFPB7
cSXJTsT+58eGTGV8UbXg6wJvgRZffxB/np6P1OK57asJhIgHWP/Xw6tYgf6njz51
8VovaTsV0/zMN0fj2ufcJE+/FY/ZQcwGc+jxqi/vjsYzgUuhZ/wbLihqdODVyBIb
zAD9I5OPkFNMGBl/54J8rtSYNnlips3DJUQ0yHUxoFRT0N6s/J20QSGKN+FLFoyC
uhl/zFlRm8bNv+9CRZcwU61+i/207k64fhTeoVRtSeVZs3IuCALlr9t7tWE0WUuS
iidaX1HRsX+27zxXR6FtnjuaTiXmO765LENZnQo+tSf9wq2GJKZ8qKqYxCJzBU5u
c5Dn+vyt/4LaEfeqD18CggShQ045a/tlPb/3l/qHhb8xxe0WzjfrcFKqpft5a6rj
fXcBy98BQRAGTJBsc16H6bOzA8neSyn+zmZKbKL1+eD1jUYSsLFxO12Sa1GStgpq
PVQkh/ISNTcK7t5c1PsJmfamhzn/wLtkjsTEJVyzNT3tV4PUpivSrJa+rhna5P6X
Lc+t8H4uzaEeRLar0k2PAHTlXRFxXgUsIAWXZJCQdrsDQhP00YiRZ4DKYJDsDdgG
78uY2I+GWTajPbPE1jyabNU2EmCurKhbn114SXUwNgbUii6clm+nNXWbvN4NBBij
fiXGZt9fIO4UDsgCN/m2HVhQAMjTJkk9KZBvR/etDprI3oZkMa5TRgIIGI+rrx7x
5kDVU5EAabmOQvUuozK3g8fU4RquHSejXVyG4oXwAjLoHy61EQiEEphwk7r1YX+B
8lu+NtXmkhlKGiJXnkS5Utlu4+GDTW2wbQg0I1/NpgSDs3HW/+eUVDZ0fKkzUtye
CFZ4w8MYvc+VocVs1CaHoqU9UsIjGq3hTSX0LIEt/qOR7xO60wqo32ttD6gV1PRQ
zevBy+ieLMybOzleIJT44N83o0ONUqcrWvIamXyBEfI9qFtOYFUxZp62BZfh5K8B
MLWu9F4VFb5v1qqMWenX045AIDI3PK97zY3xv1aJm3FBdgt3L+1YmsAEd50MmmUC
N5GfkhLKLFvKAdlFhelmA4KApeL2WACiQBvleJookyz6azEueU99Qv79TAmwSiIZ
cd2+1EbALZ9bGtBSTnTLzSQHWH0XUxhZzJgauoskTuX0xg6NgGMMIZFua2iKQq22
L0Kb7zPjeB93ze9tRoxu+YrPMUN6415+NQogclmdKlxVtINvGAaUB/WwoRssDeVb
fRTUY81jnvxnat0BcoSO598osHIdvz679nBV0CRYN5V4Bw7lkc7FjfPmiia7O6vX
313OpVrle5ecHxevA+9VK+sD9+csJwsrcMGPKYsybnGwWRk1D/PqqXIwAFBa/7Ke
M5UlAnDcNc1E+e/M6NBNm7SsbXzh1eRqMs03njXxZOeW9pl1Ki11yD4i97B0vpHK
5G11cLHR8S9UrBjRwrRBce3qvP9MpXTdxC9Dcsm/Gqpm1CYQieTVr94+XAOt2sGl
7IdZyI2sGwPMs3rFzOqg5jcOQ0jA9BfCugf7PjR3x9F7Hn62RtqQJpsuQiomwkeJ
eYfCpfUQe92QjNLxgU5JJ9TN03eEaGG4qr2BgCLxs8WK5duWAK5x9gP+cDCNi2LW
60+ia9OgdJwP4RuC+/0t+9NsjZ9BaKsTASo8/Tl0d9T1Qq3oMDwPqet62QZfaxeP
knCqfoTASHEBMKFywldaFlnTxTIDOPIvRfjpc/SeKH5ruxCglAYVS/o9eUNj8K1c
G+HU9+txr/sDq8J4mnDEVAJGcoDO3KtuEmN9ETsr0vUqr+bFcUKLrF57HOdTlPYO
4E2f+FKGqRse6vGaudYsD+Ivar+AFrIM3reoKnM7SIpJJ85qUTEAQsLZCHp9H+di
AD70S38xGUYqgItIBL+PpHCEykVMLul70cILA2lqiqKd5KcDWt64uTX+FQwS5gBa
4Hga1p10gSQRtvw2/vVcUE6BxOzVLPTVY32AvuTooC1KmtlatFyM8yFIxQxj61yF
2lkkfR6Q3/S1fLnXgV509pp+oGD1rz81bnrPKUWGy+um7X+DKpLaZ5R7RB4QATqF
Dq1gGIJ6InD2XRGY+QZaSfjrcVigtGkn9sN+Xpxu3xzaQPh3gvqBp31WXidanYCN
tsdmfzH3FeHCq1veCvqzyVNAHOdG8IDPiI7/hRWxMkZmnrUD/u3AsuSf/lgK1j4H
WDaCvpjwMzK0Jhu4firCvuvPUpwdhXbSVIlpXhO5268KnXma6RESoCPhJy64VhyV
fEzNbN8UjstHIT5o4nsXIJDaDK1hN5dRz6Po67kQQKgLiETIcPUM4vGqHeHi/46l
84U685NBdFQLDAClTzpuvF2TQaUgvLKy03QyKiLHcbifEaRdQVDwuxRvUL22UCfE
LvMPJE1j19puKeRfU92++b8ubdzL/aLyyR4op8tPsZs/pxJ3D3p0JYuKoxxdWk9T
egXjQwpDqFlHF+pZQEcuJf7L4mmu5zbq6AwLpI1WpNhwCMo88TutIA4w9WGF4U5l
Qzda1Hj+ZqtSQz3GhD5QSo9UAti/MaQyrqUlgeQEi2RKE+XS21jcORcMN6SI06gY
y/gsizv7b2A8MPQLN+AonlGsnEGidl2oBTDB0PZD+DK824paLRwwaZFM9SV+xmwE
N+Fj9cUPZvYECZcyFrFRJvfhmawczmRJlbmttNcxgvcfdqoG/YLdMeFopXdXWeQa
0IxJGf3MMidxXrjKzJ7J7xic0QKZKenidVz7BUcJsMWHvYwQ7OuS9jHp4qBFEUvZ
7wjbFFyB35jHjPP7Ze8Yk7kcwTCjk+ydnJSRnGkCKQD+kCzZsSc8tKIbz5UuSWdF
RJty4RC5VTioLKopDCWv3YwAJdxpO4f4Yj5L85lK5zfEbA0fu/aShYR0OT5XMup4
YLYAXp6Eq+mvNYe8SrZbfaayycVaiL5hF/vergoZzn2tRY72e3dFUIsZDgdLIIVu
1vvED9SYadcO5TxBtl1eD6Usvx2kdcBq5yK0GfY2JTDZUbIAtGkVOH/4viW99MHZ
sXpnLRWjP6nZU1qIsgVcioPiT+q+uCQNNyQx4L+qaqA5m5fycMfUOrNTWRGH/VOt
cbKJEiW1kTGDmllIwP6lLakgnrJPgxZOU2HX7QIFUQ9/IdeYnlVWN+mQWVzefWIT
au85IPf1Bz0TaqTvuxfeZ5asnYB0H/kk/pozt39McqMAXnhykIfXcsr/tOmxB8Hc
sC1Oj5XQ579monpnCR6bxlXOXIarizc73ZtUTaCvj6aFkv9AheYUIEoEBWCmVbjZ
I8UzQROFHQ6wEitxesHUcfNTXg6hLPddjxZMtEuLZRmjiMVox/vi3Awts0L9N1pv
+VVq7h0wVsFP0fsVg7kh2r4+Yxe/prOPFYW91TBT4bS0UnYRTojST/Qf/EzdEbZd
iOemIcICRkL48b5mJGWLzj8r46OUfI4xMrxNbgtzWC1GfqCKI5S8G9QyhZxGAVkc
OrdynwBupRLHFGzZwLGeeVIxrUMOdY7s75yf6SKVquW7GCYygU7vuNVmjA81/2I3
Q90HRXFjnSoM5rMUuD5prQrWkIxCCdAXopuslFTmGhE3zu2YAYj8bZjH077FuBCQ
eTva9Bg3eAT0b0YCvYgOhdgZup6+xz2Jv4e0U3/SFKhADl+sNzYMXARUpejiwpLO
9resjHsGw27rLpjDmpsv9Em5VjhJtwEkmClGT0XRqXjh5+RbhsE7rjK9vi/+de9b
Te/NxDc1TsVozrg1l/jjh/toQ53bughhWa/ngRyU8uRF0wW0rKcYP0lKB8wZXXhC
JuZS3AkufE+eESp35DkHAep7enCq7EOMB5tuh0lwy22e0zNNsvyJif+cbfcFvwYz
Ueq1z3tq72ILm0Jx01vKuJQHZH6lvVsB89A1qQLSTaFSwZUseXealifdzIksTWEq
DSCeJ3c+rTcvw3IqDp2K5aYF7pny1ie6r4GAbbmcjwfR0sp8yX/MRWk5Z3QSh2OZ
mSvDBIGWtlEVbVm6ozBEMQxrsjecVLUXmxZjOZg3wfW0iXMnJN4DkPOFyitcmM9w
6PQH0XsEMBkYC5v08sgPXeXt21gQFSAxYspJ6iTigOC9nLeXDVnHawOY11YxXC59
re71x9AEiWMWB4KEEde+O5asdW8ca6RwYYjWl1D/JwcWMAHNitDKE68jmyUob7fL
nwVAxVnpV/YUBxt10eFR0ehW0beOlzGlqIZ4InrpAgrS4nSaV8urJvk0Jy88k4Og
NfLIBHGcol+eyEcxvP6xUXbJAtsYmGbZWinD2l/17fS6E8MKwl9OESdCJR553vyK
WlixuTUHMY3bFTBsV5/t/ho9uPVPYxb/VzbqgZk652RhUCJWEvKeE2j73BpJnP2S
yPe3q0LhB7xSneSfZqupY5w6cOBN6/YQ4+WpZ4iXs6Cf1WsoPOiUM07yzu8dyrrp
9eJocp5ExAij9q8kHi8tSviFuF3FDEev9f4TBQiEBG4HS1p/Lvh0xc8MrdarRaXP
UC801dq6FO/g7eHzL/G93M6c9NaBraWxA9Y1Kk1cQ5CcZ9NeeV2OAiS16Xi5sfus
tAurkSZu4a4T5AYF0pb9AJ9W3giHBm9QUU5C2jb3HUaXwZRAsiZyLvnmgNZMgjGh
Vj1HNxM2h+9uS6dAKp6lh0+9VOYCY74txbEEaQfKI2eDLwLHVzI2xUsWcYJGAvGY
N2oy0lFNA71LzI1FvPP4/Z6ZWFcsMFSFT/0v65c/02D4g2W7YOGJMH4F2SYLj+mr
jLuknRicVqfNgmO3ojNN2O7IohRh+6Lig9ARp6jDbwJhSDZpizy+xTDvQCPY2GFg
1PIbANnbpHquQRwM4zAlrdX5UxLyb/4gr7FCgl6w5OMbWxNWyt32p7N3UCK+UbSq
d25ZXRg8di22L1RbXFztG42JD+hJYhpBfQg4yTUvev3nlexfTC0agG43kfbVySel
GbOJSxm/1gkET6STarMq6LwF0eg8rI7r8nlksc9MFnHg0zeXdiuxR7Sbhyd9oq8q
OnPjlU69XIfsjE13VpWEK+ecNfdfGitbU04DLm4Z4fXtPEGazVdRcnLs6/L6jq7V
aNNiA/0Vd3dQu7nlDyEF2Kb10scCM+b1o7hrI21CercPK4pMLicKZN7pCSGxNV8h
fXIRJO+ecCdeNgCcNOTP/kWMh84ngiW6hM2lGiD1GM2jsBgUoCVJIQrfqHR0b09g
AIsnn7zz3LzSGoQnpZ+B4xJtWgGsspBnQEJxQ/eKnGZiACWAkSftKW0Mmo62QPjZ
j4OUDo0XMRQD/dq/5sk8NAh3V5on9G8kZZ/P5s8B54XPXhAtatRYUcPXP23KZz5K
K4rPvF20TtVu+D0dLAR93QyD+EkfScusl9BKcTkoNUsyi4G/yqKGekzFba/IEx5M
oBnV8lerlHYG4G76vHZqvcSRoL/eFutSaFPuLI9OtlYodICVm7HWkRkW2z72s+Rq
Ccf66oA+oCXr3xiQ6k0X7x4QV1kugZocxLxyG9F/W+VxprFmxbAfuuPzzCUVYebK
y9zeaBCZsxnU9Z8EfTKEAj9h79kJIeZg4aQj16vs+FbvJD9gwIAFTvHd+9uYfGWq
Pr1xYAGSG0l4fMBdYp8LQyO90TBRLSYoFWIbv8dmOFeG6ywsQckrbCQ9lIlJ0aJN
sLM3FiZLCVex3ABy2eC1kTGsOrhsouGuJC9edc1D5ap7gkOH5Ay3i9t8bPC5F7Hd
Qn1uwC8EZpTx68BWX06lYJ56MhOYFTr288kFdOQ5h7E+gzyMTF+7hRgv5xJzfg/o
tOe0o+vcrSkrk6neBULBwVtu3QYKogTOUcYVzyPF1h2yfjbxrBMpL8efa1T+qqJD
K9eLwiOvheC4MNr2x3tOEvZwqqcfokGYVwWUYImHZtoHf7GneJNnTXMfnCiee2rh
7DAbpqXcs3ACgsbfSG3ufE2ku0MFL+oYFVgz0sHATpnLcZILX2Lew1w4rjqY234o
zCTepkrV6leomoLMdSsV7JJxxKXzxbsNnerThRYhc409jsUEbMSmjzu/mlFccoD3
d8nu5KKf/Ft9w9/xCQK19VpYuPAE2yCtay+Lx6AMI2DDwoAruoQMb8ngmESlOPab
FQIyNUDmEgoeBCWvKNh7igKp2YsiHfHdhPls7spko369FYhRb1B0Q9ymNYEXGLYD
GP1n70lzMaTmrAH7A/kefxu43iy01fdtwUeRJJwm0hheAWOK+8oOeXE/33m1aU3s
9pby+GtxCKWN2ufJg9TMHvsvSSbGNoAc3I0kCBbogXJ8Jy5HJrKMj2RSbomYCj91
nkzcDPGVb44+s485CeO17yeOmMVbw2HMVsLhuySws2klaa255476Nj+U0MEIgN0x
mTQB7KQzKPQq5KQeLVW4h4WcklWy2gJMH2LLUxssSLDdVl93kivrI4M4ELmHtzvg
M4XMktsOWdYJXijvQ77RhoQaDECFbrBiP+H2TvDpm/Momevo5KBlMNDH+V8JEUbV
abGSuseqiz0ms/g7yTwSe+sAuOfB0+oyWVplsExNyIs4dtArt4HOHQFAb+WRppUy
s48jTeJkz56I7CzNDr06h8cxflm9+697oqxwr/aLT8AYQqVRJyTGjQDnlQPyQjEB
0oPaM29E8gGGzGjMyVMOdEhWPrXq2TBWyzmNrhyA8ZHu8wfPJ6WQESlD8QhP2YGl
vkCO0yyqkC97T6yeSuabC6LFIiQktOFnnSU8m2FdtFZCUYs7zpmTqHTh3pnAqXv9
3MhqL7Ci7O1Do0mcMclcKuwvIPfwAvwe4ecOS0vPDo3rBjnQzc4qYyQ18jZhyek8
9/MMXkHMIeJeIx5fLbTYwtoir/CHOmt9TgMrmQLtVzAKMDk3rm5rnZ++6/4FL0eo
HveqEXaEvDFEZqNHy72hfzMkDHKImF1FrcTbiIo3yoqyGNXEEF1g1SlbYY0mdSO7
P3LpRNe81Ii+b66DZXoDzKqpxA75g/rq+f7ffwYeEDbnednz+ECgpHuQHpch1lNS
hRrKb0dlb5rVOgcArJs5Mv8KQ3NyYkEO3GdjmsiYotM7xiZxRSVXqZpCgbxmykUg
KObXKQ2jGGXyXuPjVY3ZfCsftogouPYCXWo14qsAxls+lCWJGd6Eg7DKupbb3MSg
b1A65aOk34UwjTjAqpeGPuS9XQR70rp4O54NisH7nkzzYJ+txVjaX53bGJHpJCKZ
v76O06g3rA+saN9QOufmbiZ9/lYyoa5Mte7y/76ic/jrIkdppks1GCYComsjFeAF
N4g0WQqbVV9UfdnVLDx/5gP85H7CIMdfG7sbuCHEOBwG0fohib6DO9BD5tJ8LVvo
gibLdrelYyU776eKUzvAUkqSRiRbgvl1V7V6xj9eB8jB9mskZwiCmoHWv94Q6eEs
syT5gxonFBk6fcsBE0syTeJzbreQ6x/TXEUu+0bHadwrNephYz7X3kxhQYv2niX2
9SsWmvZW7Wbj2PJvVn9MAcQ4eBc20g2FjgkHvArg+BIfXKT+iT30giNNtpo0xFwJ
rZSV0GeR9CLpOp/CFfa+h96/Cq9efqcrwMI2AE/5Rz3E/4m8hogkd5qhBSp+eUHV
5adHdvp2fQ77vNgOmX5KnAjIz0dIcRzhf6Bwgd9DepcjOY6FsdZdSGKbCVXXiowM
dXtRwFHxvNEW8Hinv+cdAmnQV3qf+QqkIJMqo2BQbLRosu8rLQe9rXJ0J6AuGFGK
OLDqhVOiMsKSFeTFqr0hag1L3QoPr57CoJrG8tDjh4yaO7Iamh93DY/eoxYUuZAK
WzdShIMEN8KW4prDw/gVSl1H2cD1ee92S3q7cjcriys9EvrtLqYQvf1UghTt8amq
lCpIZ0+tjuGEb+07XG/91B9YHLQVD7NHU1S2p4s7E476lxEsPuoajOZWAT2aBzcU
jf42X3cAyTpEvNHyB7xyP/my+ofcbQlzq1g2SSN69HC6Xb1GAXEQgfbMCIVG6OYq
QGlgsvO5kh6ePPl6BBX3lWJvjQZ/QNXMRxN217C5mABIKwK/O7oa3ScQ18oQPzk5
qis8NHcBBUgdIWf5lAvfST0yJgxJ1ihHuJiIqCy0J4fvOL5quVmPOL+jbkxuGcRR
QmWxpvh4/EvlgmallzG4oTv97ejCpVwjURDhn0qP5sPEaab0iD2TtBqi7IL5FZ8G
2rCJ97ge5Tk/4D9R31YFy45F/70viU+xeJRE8cDQQxdECCURMQ9VIpjyK9U9uMN1
pMcmbZU5B2tfaOfAxN4DgRscICYt1L3sv+QWG+8QwSwiwNWqqaTaNK2jtKKZsWNV
QAzD16NRJMqxwZklvq+MgBvmuC1AyzcMG2lFl9s2r9BFB7MIDXJOBdeTzr4wKtos
xB/thaujmurWNDUIcRMbOHy70L4ZJANwv/QpHImgZPpoVD4NnVCgC+CLcyJXnKwC
VBc1aS0KTd6PqBmkwd+F90HswoYerH3l8gjw1TQRcN/Z1mjgZzLDROQ7kuRqMKI5
23Ca2JyHedOV5SiMzPBHFOUL5NiUMhICVNRPCp2KyfzCP2nq/KnpMjGlrgeQjObz
CHoDDm250PCpcWXt8BBEX8KsEheVmPOwEWh8keIO2yGg+TKeV6LSegiD0USVvFvn
h0zSQJ+1cDsbUWGALOvGOIZFBvBPVpVFNlt1+JlPs5AugtTWJR7akX38tJ2SgTVf
qYrjQvE8Btw2KvPbibd4gn8wavX2HPW0ZeqSn9xlQT+Na09LPC+gGOCfZGquxPM/
tTHwiTAa1A6O2TREXgOaPuUMSLsDFJAXz6bMco/4KmBSNhCh4gc9gl4ENhfQdGFp
Yv7fm9Zr2j1yD9B9kW2ms68YsblkJeoPd+jFdmC8dcIoYg8M+pnqogNycAu2IzmZ
tU6et4+NOinQsCvogu1whHg3/PjTKlQJFZmAyHYVov3QGWQ5p68Z8JLH2/97m7TR
GVxLq/8MU6nvdsgsJs1KsP8dsaOGnF57PUYBQUHpBg+AKG62NpCPqX+mmjwYxOpe
+T9I0LmBL3jwO0xZQILM5vxSw+/e6weMcAr0s2YopYeBYZon8dn5MUe8IlDPXckS
jjiMIBatMBx4kaOMAMQANw1Y/XKJbMPc2DdWQtvElDqggBHdTNK1KyuLsVlQNfXi
l8dq2tb4wE3KWCRtT3atoPe9lp/ybXqlNpmmAHZpmqiWpcZE/F3RQCm++D/a9VvJ
bqOH/4NN22VXJK3qiL5gGrM3hgxN16N3EjN2MgdzeOYpjSIDfxpwwapN5YL9p0qK
rOApcqG05q7eqhZZX5XfdRhNBApQx7Pi72xgvoBOOdbs94zMMxhK7df/A3ico7PG
1urrKRYzYTWoqF2y3md4MZgia0apC7jkPILkWZsxwQXQfR1IW9GBBRlzaAkPiJM+
LHBBkbyvn/6RdDWwqUCQyYUQ8tZwOnlNihinKXn+mLP2Plfps8ln3H5rwl8K9A+J
VHUnFXuYevybqNVLczL5/gVLBbabiAWF4ubRkwV1JqYnMPf3EaLbGdJpmdoZWx56
d9uYEJkuElvE6sn41Fxn/b88kGNFKNVvEDhvT9kwiKI3d7vZ5xSdb/njSBpYPwD/
/D8JGtJg+groThQ0UXIoohEul7a6F0Lp3RE2+tn6PVkBfA9wTft/V8EknoGM+4Xn
9AYAwHu0EzZhilIDCr4PuyaHmgI16EWrcUTAK7dnwYLPK19zuuAQlKiWsREqUcOk
KJVBAZ2JwmSEz/zdOWCCwwo+DvQUmsqpZArPrGCsVNl8IbYeKTxnNKFvmSKleK6D
KjfL8B10Q+CZIKA4hrg33wkiV/Th8R+g5V+1wRqICc/rkCpBLi3zPs1ib8Yb4gcm
u5lai1S9UsDRFif1pnpcW+vkM6QzucdgLv4J5cy5ahtqawNzcSb66Vdb0xf0vGOJ
AVlVZVB498h2TvwXl5W8fCTe1WDKfXtO5rDiYyfwmTZ4ET4nHkp3m3mVgHwDxvXz
Arw0RLR1ECryLehfV6tLFJQU1dW+7fa/SKDHLbyxAhGd4nwvjgFXi5pWdNCovQMp
40tlKC2Lms3JWUDyEUyzGqMpYRarRwh1AR0KwW5qrT0ocPI/RPc4do1vJERl4xkz
Hwiomxpah4UAfJsG7XIVpbiQ/XzvcWKzCVNNgFufhjkIAIs9g3E14YxOdvxrGzpn
BBXUkbeQ6UpyVgmT3j9jQY/lfbRFmPR3F3VMZDbiLt6/Rt90P/wm9+NztkXZ3Jsh
seGTgkEq4Du0zJ1JwcEBxEnEYpuvuArku/JsFFhvbTMG7ajfVRwb9ettd+3zGjgB
9n0cUwLiWOr297/92Ne6gFY9pbiCUHg5HjOUEhxkxdJZ3vatg0bhN2SyjElkz8JH
gwWGD3NC1WYxV346yK7T+akUHfHCmBjw8y0fu+lik2fcXEw13vVfBvX9qEFt3rMi
1cTIetJ+yGM5nengDycZNYi48vJGnwFfDRawgFZf7IzpubR/PfzYiQnpudf2/C3B
zvN+s9KLav8ELV2yOFjevtKaLIe5T2bS0RfW6U06ge5MmZVYjcQuLfWNzmXs9evR
f5g1p9jc9rmxyFvuErnL9f2uZxsi6psaP01jv296S42aY2+Vb2vjyo+j/KfDVi04
tW4251cJUmcfSvyAyY9RD+SAdJ5KMVZ3pJC8S2dSAh32r1+E5afpbc7M8ruq69ET
a4++Rm5mef3zXiEFof2xY97ahVhcBP1DDwlhjzVEnaFHyywwqTCZPQuxn1eLAdwc
nLIey7P+wg4gUJZnqrbAo1HXjRbOZGEucjdg6Ryrshw/tt6/+UCxz+mF1DN68nRI
vqvd+nm8+FjN5NLogVTcCWwuxIicA3fMf+yYQWXk+KYpOyQkxiRM31bTKDg0c2qk
sr1aDAzhxaZYhoUMlXx4Ikt/ShC5YQRLQLQ59cYsDFN2cwHQ89RjXK41GtgAHIyC
yDOIBQPycY6qCglp9XCXx2bFd8Ay3a+K5ARx/tlVOUPIB61hrEC3HYh/KlrKAIFN
hmRHB6FrFZjv79q9bMr7vGriSYQh8olPKPYz4FfQ7/jZLYGzFEvOmk3r3MNnLVjb
zQfSsfnJH4ReFLMCfcX2JLf+cXQnjI02DuP3JEubtpBfq2696RVOUd/8K68oKsb+
nR2JRqX1NfdK2bqSMJ0n1nIsQvjAKvRuy3po3mWl00SfNLf49jxv8ZF2nC1hFpcf
9RGV6xGUbXX10Y44x//72viVEbWgk8MEYxDGNT0oAmZJqQTZgYNNqdQjYHk/IkN0
QoOTEr+Ad3OCgv3dN1jAKXljMBfLWERn5bUaTpfzZZ8QDOHKgsyEYsgO8vbA98Bi
w7OaFCIIYrvbFPyEP0pktAeoB/XEYbGtEiRYrSJmLEcGuuhYICVKo8hKM1/B1vs3
e4xgoxXc4tqD1vG/5UBfFbJnyPATFTcDeVXSfCpqYdeepk8KtGeY8vPo53BQSNX4
w1KJK1168XRT4zrz83D0Etac4D3quqj91MnV8vJ5QihyTWXmOeAMDDHyTgGyyscg
5/HiWzAGKWtVj4Xd/0T3p6vvSwg6QwxgBSHazX8PQjwiFAskBbJHLDizUTno2sIN
EaXeGbQ25/nLiIX9CRJklpD9FphvswP5cG/9dTzVGlHa6MBZeYXcbeoyAU0icWqH
cCajD1iMRj53CIyHSuuXE7CsFKqcHmiu7vE1c8R6u4ynN85AdcKj0aPgjmTIUlAJ
/hvrAhnyrU5KNTd/sxD3ZbZGh9jyUpYvGvKiyBQwEl1Wc/4xSsNZG6+qj/UPeQeW
cIpHP7bUxsKXOcnYrLOIlRRV8BVNnAJVbunggdgeb71C6agiQILVO9DQxa8jmjtN
p2NgUQ/+CWPv8Gpa74zoZhsu6tNrGWfwY2C4f6wg0qXfP79sUO4cT4T3bkFRU6BB
NTNTnZ7MzGaku3G7GBBr2lx+xAAmsfpZXDuPQuhJQ5Rsa90YXl5OrXoYoplSd0iK
sYoi+4isKdsJUXI4TH/8+lLEK5LOBbjV410aBlqIqtEvwN3Iowzwmx73eET7LRs2
UPgAfjhnPYbqYdnXkE2lMnxsOKVtInJOnjTxEiPh89ZwtoCEgSSCEQHzzhYl28Ct
vhcVn3qWI7K+J+R873krX8yJ9Bj/9hernzVc65of2LC4+o6NF5LQyCzcSBo6YcFk
HGIiEeTAjDG1lsRUfbVBPt1jAAAOMWIv4C5aORq7ysnPRvpADHWBbvI93w/oc0s3
pC5nxG4V6YBEY58tlN5hK4Ayxeq8RnDGduLeFt1/Gt60DdSdLif6j4OJUWn3Onjc
qxbLB/n6kGOj31yJBtYj+zbJtit6HTj3IwwBG4LeLeRAPfhXtCvKr1Xm1WyjYFXQ
Nm7/KYn+eqeJYG9EdJeebK8Sp9WmAAk2fR1W44O1yNxj/vLYjvuqNcgfHc55HKy3
QMrc2i4jzEZLugJU7UmZmo/rSszFRNlIf9ThF3VvZXL5P/5EDJGAT88FtOLBIXtD
s/59x86/KtlFbvkkv/xmAzKA0BIzG9xzXG7OfpH4SU699qkXXr5iFuNM1fLJADaF
cxitqqtuQe4vZK9aJCZgQS/C4hyJL3ZCqNCUmvzMAfVY37/u+nZoE1QXtNhfff1d
TYVPcU+j7Of8F1WqGH+qCuPdYg2sBIRSvDtDlI3zQQz98ExF/0TlUxsM/CuxpcH8
vpPEFJupd7DL0lhiQ5QVOkaUC5KBwkijZmOi0ZRrSeLlcqg3CEeXWzioDZjF+O9x
PK62wuw22YW6EB+sQ844pE3przl4mz9HDAdgv7S0sSbdAO7pUPlWwPByRN01q6Qa
glWbEHELpLihIf0BoBJkihorEFcuNPdawiBgENPSLBqohz2busJgDviCSMAhPObz
oRPc96UnC7y7IePcTuOi8Esu+2A0JyNCd3TAkQVv7zeohLsDjrcynn1d6Vh0+Qju
ZP7mdhJhbCQv4qPUBe1fcDgfQ8gUDeGYyaKOSyTSGkFdp132TrKpbReU17eQVmyd
K3hpXgeR6GpTz7+tgdSrLcbX118gnVUrIl6gwZbW/PWwwvtNzlZBDdzPEEfq9Wg0
lpMM0mlMdCBb8seyDtYInvFuXGMu4f4YZ35XSfNvad6UD1OukkDJMUobZCeKn2Qm
U6YH68cIADtiwkK9Kdu46eDwcNCAn4D5PBXYIlhaXubyDdNMb7utJWWkoKdXQibh
6jqm9jWYc1KPmA5/5/Ei9vTPmJUIvzKt3IBAYfFWzW1trK3sYEwOpBmUIGyIXaTR
eoorXK+85HJVD+c/QAPzNsz0xNYjrkmkH7gdqDjvvLm0ZTWspjtTObUMcfBiE44k
3289mHjwiknH+69n2vLk+lLlQ0kjpbLdZjL628CYj3IonVDK3NEILgT+8mv15IRZ
wraO1rT4kMQLzVjIfve+Qy3VS7fL/hPDsLDe6qOkVQYZXtsJyv1SfAogCtFhaXef
Z15D6jDfts7DpH01FSQE2Dl4ASCBMRSZac/Y/5sWk2GbxPU8XJf39WF6RSH9Qppc
UTEje09vAz4wWOF1NSrJhktuuPYGRObBEc4uHCkliaegAq2njWlbAg99r3euMO9y
Sjpg6a7kWfR05Dn0NCChYM6lLDFE9a7G6WajlffR3Gaa5opWI1eEG39kZWFoxxlS
k/SdpMBDxjCJRn5ZL3T8qbIeyWqn/eAk0k4pIzsgwRnmQCryM3Hpo5lIVv0e47IP
+AWZEx2HXLk/6lfHJTIFGN8I5obpOlOOcrLqos4lzFye00zakp3tMoYMHWKvANMl
YfDyFaC4gd6ue4SAfbMZCe9IYoajSNFn3zC9SR+aHRF6NyGzmBZkxs0yBzUJZHhB
tMzBvc7VPEWVAcrI9i7WZp2gZTH1gcaOVcEBwEi3KqDEPVUi165EUemOom5lICIR
BY6eKPjRTTnXJhwCCv9h1SGz/JkOj2EI7oY5UiAgEtzoxFj8haMrpWv9evDrU43/
CYF2aBqlBVNXiSjA5GSbBiytKVgLqxqHstxVDyH3kwFXhKpGr72yGqO0DqcmZwoA
NdnVsL+N0yuIymXqluvDQu39QeVKkM8Svrzm6u2mIh6AgLmK8ddAOMeFp522N/hZ
9hWOiorBLdAOW7nhqzbLv4HBgMWMQQAQtFTSntUEjJz4wKmW+IBNSE6pi18BINAf
6nhatQOuf4zU9NsxGQimXj5g5RI86LkvHbzhqb1QkPZwFbGfiN7ZF8YMI4qie0pq
x21BPXYRrBgxyoumEiiDy986X1SpLQDNaf7ROIOoAN7p10k8LF2KiU3WAI+ijphm
YfJbjbQPdY51FXNMSF3HMnTjrZ4kTYD6iHRZcRxFd4gQ60Mg79szxT5viZUj2KG9
UpyW3vWCZbj/jr7KabZsjAYZ913dcUUP9vcqXntfnAqev1ulm435S4hTyweRh8Jl
ibEgK+/9IEBhmGgQx1Qd9FQnKnZbav8IkN0OnEMWo/FiySUhN+9fielnETSRwK+H
X+KCnEfZeRBJuNmEB10auF++0+1WoH39PXnefckJCf+CgSniN/B2+vrFTEbiYAQT
SHcEVFX0QJ8pNfNQKcZsbmui5LlTVYBVluLna5aTXZSexLWLnL0/ws+HlBeQSfHz
HNi2Ho3kQNKaR1zP9z5JGbANtHyyBgAhJk4j0/ibYel1erCY7+2IjDsAqDTTBg2f
xWzZ1lX3MMl3m6p3TkpbiMPIpTd9g/4u8hNWsv7v2nD7/OD4OQ7DIR5hUwq0N8nH
mez8Wi2jiQ2J8Yi1JETzLFUYr/RZ8vo0JOUh361sbaGWDHOD2qpLPhkxL9jh9DWO
sCbII/CsQM43o9ZgmAct4nFJfncDRvRjN8CNbfA3rvA9VD8T1iMnTW2TvOi7loH9
grDpUUuw6lt9uQux55S4IOte0MhJ8UUKAWYYcQ+9eTXOgKypyjKiLwyolh+IXLDi
UA/Kz+b92typuFR/HtxhSNvqtFBjgG6OQYq5YNq80d2pg6jVgU0dgCo0orUdFh4v
svz4/tNc440g4DJWPSr/sEIfYD4edHJ9hiKYj++uN1Z9iS7AP6H/v/jaGupY7QyX
i4zC7qTP4Et1X7/zecIg0WqSDZeHttzUlzqKxjoVyVz8ep6WjFkqjV1zAWDbLG0E
R8CB2yl4icInwAZhiXl3nar904hRnEmGbB7p6pc5hDWAShdUNxUXpJOvuFlo1VB8
LtYeUw1Rre2QnAqZyBkcJP9W8hQGFQ32vehDSPXQAC9+XmoD9TAJwBJj3nF+kS7F
1V6tWhpPnsXrQ1uUz9RHwkZMVBDitWRqF8Xao71jnnexiUVVr7uq9mwVC0zjeE8j
AmNF7cyhJRQB5wBw9I2Gp0EVla210wzj40740y6GZWm0cra6YpaUPKZZC7W9mpso
krQA3Fuo//1eddzpEHQKhTrJdyZyQKHS+bUEKDZ3pOaaO8HWJAY1oMRqJpOA1MyB
CfjBpOezrb8O0MvlXNam5n10dV+OB6r+9BIDjn4brv3m8t08L65zUuMjQ6nPhNGE
ixlbuh3xislgVb1PwFuOBuJ2gJk4qHNuS84q7Q9aD3fk6HIZT1aQk/IzRZf45hDX
MaiCyPjdKuA0uS9NWTttoR+0MHKSoEof55F2QsTRLIVCvYM8x37u217B0AW1o2J1
S49vJeglm5EiWxhg/1Y+VQOYtWXZLSYAOZKL9yo20FVx22Vr6+aKMLQvuYEcJdXY
q31Pyf9/xZy1G9FLT2/CK8K1B5IYQSwyWTPmwWbxH3PXOsewet6X9zFOZ6VEfJ7G
SAAzWpiYDysyN+BIrDeBxqZTtWldRhH4Wh5fol+lNLX+NsyzN66K0Ih4Kacioitg
jnkaIr2mebZBQiunJxIu8eMBwCzBO/nBPJHcGwM8SptlhROF/+U9zx3xRfl8MKEp
wHhh2t3FmPSotc4sVXUHUHiWU7W+a9izfQv8a9PM/aQzPiKzZEYVyXYycy2eOq+1
232TsN0KhTYcQ36snDohyZLTniwmTYEXccsAdIWYZ6DgSCNty6kXV490FvULBn2T
bnfV2BYt1VFcjTX9PxfZsryKeejYUZWclk2sXb9pTpvA0pLUFdAsNZ7Yuc6z+tSY
raSSUw2YUv42VuTuKh2peXrNNUqHpywEj/yvkett02kEkSq7aJ2vW9iPrC5/xmXz
mB9AOTgjKpJVoCvNY8AudVjdP38U2it6HHNT17Af4lySEpOZLfuCkATsf/HIIvH8
KM+FxsKB6cPnSC2+BfJ386rzfCFSOykmd/sNbzw3Y/wpTz7tpGME0zB4cEHJdR64
FwfEz+ZxXsSDEJDK91cF+GE2RA2q4RX/phY53V2P7ouWKWjolHV3JDBlVXn1JPvX
+8NryT8eKLvANFkRT33mrxPmlpxemD75UiAn+la031EsqcoVUpZ/UDsv2ztPPNaW
mNB2tsGzL7BM3RG7TSCbUaI4nHWSMdwtTs81TNEcZNVgIAu2QdvxKEI0gjsqtqwQ
/C7iC/f/LrqCID+g3Gc017A0+4+jnZxnXvVPBuNYEW6H4InazVh7GJoRyzhNqtGw
hfMjak6f1ULrMrY2O2TbbVW2wAY7dz55eFx1bXUveNzDaxW/MEvUZNCyX2bwR8R/
6fPqKqbx/p8CP5iornp3xdd4+dkKASqbc/kZKJZX5tOhJHRTLgGUBC+B9fJBtAt/
W/B8mDrH/7krIJn69dG0KzUjE6DAKKvdvcHsSCC+STMz7Pf6ICIXGBbGI6l9I5c3
EqXQt0p0OdbgakyqSmsdxR6lhWJDr24V39jC4HgWEsvqzUoYWPA1Em7i4671koKU
1vLPY7LQOmLt7P0Z7v46BaQtMsIdKqPZoDIW52FTiXagnmsEiIFBVxt/Hcdfn1Ei
S0CixPnioi7DhTF9jggmy2qIlp/t8Ia+W3qXw1/LYHlWrMgvmM2sg8GjiNzgU7R9
IwUfuxJY0tONwsv+rnScl2zYS5f2wCPmUB+DzCbcg9wrTaQAX9ea5M2Tfivj1MfW
H87nYnegsMKMxqYpkyTaphYv4qEJPWtAoalFdulcjJfFqql8Va7NNaX2Vdt6iEla
3B+hERwD6RWX7i9h+78tMgVr1d/kA4fHVHagmMXJg1hGZ6+enq3aBXNl6J1orVAq
YtSjymAYUkYUNx8IXotwIlQRc8b0i1N5L4QGpddMGLR/71GxmvaP0HuF9ufFlqeB
Z1ai32fKYxaZREu5j9H5tROCqvTYkC9byrygzE19CpmHJFDmmp2dpz+K3liCDk7o
iWHzT77tKHPVK1dj0K1lGJkdz1l/hf3QFSnDUC2YcnMN2vVsxnsxiCBnfj+QI4xw
a8tM2gqhKVtTKviplTjJpk8+P5jjL4HoHZQ9uD2e37hxZimL/ZTrJArbnA68tuhX
vPOjRwOvTjKtP9jt2KLA6A3v0HKZyqNefaHcetnQVLHpNJDLb/7R6kcjCtgMhdB1
xQ2GGDZzGL0pqVomoZ7GFp8u+td5508VTQvtnvF/cVKspIENZofRUTDbp5QUnKAD
qBgur9dYosdvRfIV3v9DneUGEEkYXlqtLioLTxGZwXX3hcnZXkvudsRNrFBFTva/
Ho7xxX40E6wpa16HWoBkewJEmU55RI9VNmftl7zkIFi8dyOgYrpC8CJ70M3Hf5/o
H3G4SuQ709NvCLhd6ggfLmhDuEHoCZtNz6jvbiTTJlwEGRECTevhfF9bWbkqaZ9G
dTj493f9kFJHMwebuFisFw87Jg+E8rtHml2g1aRKIQkMoteIPYzvIRp7HGi1cWkT
p9nj/32kVoL7txceXJnm23xUMgf1iO/2iRUV2nnlakmY0pwG43ltLXBERI2aH9Qz
FnAw6vbqlmO8kSFPSSNcUlmF40j/OLmGnKjziWnLeROYEq1iFOY9Qj65fvcDAbpe
59/xfDfHB5geHIl9MT5NqiUQyCLybKUufIWZzCeu6UiR8iQfjVLXA6a5rmQ3cCky
r2KQUs2zKQnVNRWu2US8kz7N6JpaYT5cTw7Ya+/VbHxpaBgwWQuy1ZfmdXRaA0nL
775+bC9+f2HiL7gS3ed4FnOoF7ejB14n2W5pyau7KSPbFQEP0LNIFYB8OHiMWXin
VgJSBGaNEOmKirWB7eBGZqfHayeogzCxLwAAL6S/rtibMG9X3x4gIxAUvdsGLqid
XyB5Y1Cl3et0NnP8PVlrwihEWukVz+9/7Xr3JfcpwIKzpf5baGvattdvF+c+gN6d
iFPuO2J/EupouMjaEW1cl0ssLujVp3FpGbgVk+mv9UbK7cJTnhZECnjuShm3sWYA
DSt0VKJ66sf4UGnow/CL4kAo8YLQYiGR2BVst8LXEjG2HtISl2VifH0xOafCVVVP
DBPyOCi21zrEr+RWdWgY2vJm2YndpsMeIag7/XLWPJZX+CYpdk10ZAYmRzB/pGzt
SSnfseEa4xFS4QvOAzkUxNB+8jT5ebSCFPZdWJLv5VcLNlLHfJvEgwRM2f4bjpbG
kkY1/85/Sya71SD75pWBGs053lIus+77EkqpF7nt41JzvuZa4czixeQnbuuRSwZ6
phvcTlDBxYraNNzNtJOJhMt72pukgMk5cPjtkcqmmQJ8Zl1rfzGpVt7muZ6rBWZd
SbK3TKfVXx18iyxczISQ80KMfnKPjUxaJfwRZ+bJsVSxpNms2jBemaeac73ZER36
G1OKlZrWfA3HmGkAA8bvbN6cKIkO2eg+1RrdZEealsHMEHhdjLNTZquXJLzdMHaK
zSTbO/WsE6hu7LKpRzxIIiFrTvjINSXIEU+TNPNb5+twsajYhCajJ4UCrvawbOh7
nC3rw5bbH1JMrvcJMI09A9VIFxFoo13YDdIOBTJK1c3kWoNsnMZhSViZuVqhndJ+
EmW1MVOtklCHMx/BtiUpqEGXdZJobod9/yhjZq+ztFyYJ0UgSWJlPszG3jguY8nY
9i7dbFu6R6FzkFflXIKDUfEV0znN3DBXtjAZ/Gsh77ffdcLYS551bI5WlSqzFK1E
Jmgxv/vo9i79yuHxs0Wo1/yfyz4EiC5uhxpo7JQf3e/OEEYaIyz4EwmTDF5hRKg+
9k0Xm/Ify5lSqBn91Z08rlqdW7XbGdsf0ySmi9rONwiVZK6fvfmX85WUq/EJtqrt
qMhIrRAlNCTuAD/AvjkvZh83O5uPNGvfr2zf0i0ABVcXLgihyqA5v7KPB4dYtRZq
2ubAPxo14x5Ojz84NxpzKwXlZ15zUYrT1Nk7VivJ9I/Ts1a58p8KIyfmyhJkdKKe
hCrfO8y1MvLfsiAU/3GB7zglz7kB0eW9nl3lLcl0hi2yVrQKUW5xN6DmfBWXM1rM
WW63sHmm0ZGnp2BR/t1zPssleQ7ZwLygrsASa0bJPXuMItPY68VBNxPaDaxNK+Oi
3tinFFHaTapcQ3gana2gFedRktE9ultfjag8peaUC7MUFx3nct5q/DAC0S4uqdbk
AlCPFw1LEOSCBS4eV8B3cS5BUdi891wQ2aCNmOrjlKZ6jHBO8k7PnrOt/MBDdtOt
BK6bh8QqVEuH52IeYwNgKjjWrLLtKo7jhsoVIdighCfNVRVt0srHS58H3ptvtvmM
rKN3LSFrS/8dlHXufLq/KT3a579jkm6EKTJxXFAxA7xxjT3XVngYkTUa1yncJD3x
RmOC8q8nv5aYAQs5UTqB+OniTdDShu5dA239L6SyzBA1mmiwmX9nikGeWR1DSNtF
FHVpZS3SoHpgt52bmQFzuE6HPx+LtxXoiS/SYkdOxjP1cCQk4YWHuXUuurIZXq9+
CQEcsOs/RVU/KLAd4Twlv8ZhtKS+88MhHZoQhdJwL1cJ9S2fieJvGpTijn+1GCSn
AXuUH6faXD5jGGz6Y7zymMbiA6++/2+Jw8Jxz9CdfLzBB9rjanyeMl4M2SvtSqTy
JWwzwVkCKaZb9G/ufzSjSUQJI72oGe8NmxWs6o0yaIajmArcHKj6aM36cpNA+kHj
DwR+2pIHc02SmC5Q13QNccaYX0Dy3bth4YXsUPeUfhWysXI9gWab0HVQevKguCCq
EEJyH0wVFK+BMi+7rIWMxXuTwifZDte7m7q00uh9XqnwB6dF1xumFr6TcePGjHG1
W5Bb/1mNZAVu6iN0lnE0Gzdm9puJBGLFyyqOqrKVvcN5JREPpHuEQM3b1CQoobAh
EaDvyUqhuRYu4dC0+0bpuwVYgKcW72/9Bwt0N03r79UB+okHh1DG/u4Op3HNK1GT
gltvy3Tm4h/D/k3/mfKbh5Vj1k8gBhci/DQ3j+P7F8dPYxYTa+z+vA/FAiv1lgT/
PH2ZIPVz1hI+TK8Gi+0DbWxIZskU7UGcqNHlrD8noTTEgTjmhAvfU0Yhht9E7Lqt
gz+v7TKf0n4AFVFF+wIg6iLSqD4/48Xl1iBtgiy+anoBldSNa5O9/ZtR3oxz26d5
3qK6XRKYoFBEwdjZE21zvIfiBHoUtEIX8L96JVg/L+jJNOhBc2mZeU8UTPWkcAAW
Lhtq4b1Dwo8f/pDlC/Z5/khR3xouUYhjrcFquO+C5Pb1BvlBB8R4k7Q38gi2EwDs
cLkOICalpsxIMQNp2fsQhhY3vjPt/5aTzTE5Qvnh4YfmFwX0OXhLw9iGcgFmj7ce
rD+boXzzySSXt/pse1BR4bupKbGC+skcWdSM/6zbiTdg8Yd/qdV/fvgZ6oSFyPvU
rxDlYFdMcTOLZ589I7pXK0UvJwXepQJPzrjhOUGnkeexO592nDVnSncj9pXX/lDp
EklDsvCOXGMUYGsu30DcJsIM3zjmagEHbvSwbnYeYbFNUApQdnkIxtdjXTVgKaue
rFhwzcRdt7+bQUqEufw7Y8HEoyvwqd8ItVy0VXqxZP4NXPG7v5XHt0Iqaxc10e4K
fjhdFlh+iK14xKEjP11odSLLvMxY9Sg5wIBOFLtdILduA/Cs+Vbktda2buxSMQ/F
7Bt34BfugGlz93QVvGFd0FnHl6/aBlFB9/6PKxmyVVSHpfgZUvnN7LJGs33D8VZd
Wwd8AC2nnhlxFNor9VFZY0qOEhPCNgzxKZsrDETL4psGxMl0Jrotyq4VgGUiU+M9
VYVItZ2b7sFUT0Zv653vt2sMGvg0FkBIZ3F2NsRlYhzF3A7V0zTSY5WegbhTobJJ
UhKN2Po6YMcgADX42vf+eZXjmrgqY2LtHP8PScMB9fzKch25oyevLJXKsQh35pYq
UO5lnS003k9QTyGqoWTsZSzlFUHbNmDqEltxBSk37eOiDmn5tJmseHzMb36UnMnm
OBmMt7stJXMe8NptDKG3OI5zb6bYCPemE3XrbyJkzs1oUoSY5WbLaB8+CIXYmAeY
z03zQdqmPK2ueHsVvI7xuYlYjtSgzLvfGLo1TlBgsXEAWIEZ65Rr78LdczHeSeff
TOUmFaBd/G3pcYip2K0Yo+zdfk4kPAYv+KALdzTuXmgTdNAKKMMGKtvxvJIM5OYZ
5yB/VmdhAQDs1SSt+BTtFjY20IjGb3fePoVfKziU7uQPcP/zAMmVi8z0u569z42Z
z9Xaa7Ei4w+6Uv9/mLX6lf45NDTe2DikJbS3IZMeHFPNU9X0ccel/i8hW4BQXA4M
6SDEvz/9wWvJE/USOrqSAM2W5R27YEJ3KiGcPN3jYjA0/STvL/SiQ+1pUARs6Ung
/qI38Zg0ukz1Oz3wHNJdZULuUd9y+ampoXUmQg/oFA+L8Bsd9wlcTcQVN4Msb4eK
HeB4ZUMs33K1mKGgp1SrTr+tzQHyjCTWYMUd6tbZPUoCciwB+0wTEIbc0yKqNBur
fcp7LSmPuIHNwy0aip4eBZyuWUZWoMfDdtN4jeJ8qusB+IIoballGMx9+s+f5dwm
g1TIwTFRF/R8QeOOdDJXA4M8FP/wytfH4+S4NG90GQmoAz9h39tQVd8Yky61omcK
NeR+Pul6aPDnms/6Mg1CMGOiG3YOD57JoNvXctBHchm2OtgECYfSBZ50Yg53NUBZ
+HyRHpJWL4PH70jg6S53Qb+rO63WFmRwusHAAYX5qHJoyiD1ZFiM5rRhuQHZqTox
svIkjttEmgc8y7ZRgLSQwpDqvN0Tg5qmTktbPL88Lc5yXHFDMcs0F2nqtpWP5/0U
ipHx2jFwcjCnKBdpi1A9AX78VnVxZzalS34uP0gfblMqOc1r5m9yB6CGitvzdHIK
H5ImyBAmcFCJnbaUNKu7PE9ZI/GoQgtcBcK7TLo3vDfWsl5sGc7pluzEDdVkZ9VB
AVVBQoKis+KOg86vAoznuw26y8WtYA/P/RJrxhb9Ul1oVRKv1O+nUeiNLEdTcjI+
mv6dj2Bqb0ORF0ApUYbDcytQKcQ5VXn+j5cBLDOzKCEvw6U1AvfobK3/3VsEQjmT
rmFrZjp3k3qLZttAaBGhzR3rL7B0cbwbcS/y8MyBFcTjScUxQ6Gu6/BOZWhEGRn+
h9e5pWLQRrpHQK6xtPEq0MTBoWhl1cKIDacWsZaG7xIPqoP5VqIQvL4BUg/QZmQm
ZJ4poQtuztQLxa2oUe4KFP8NCw92iY9h4eHvxrwWlSAX0XO8fhwM+UndwbIZlHwk
gJTvzqc7VVn4k9MHkEEIlvOMBc1yJ8FLZuxVceDFOEv2coSi3eyrADUbpgsWU/WC
kj9ArswLAhYyN9DXCbgGRkTM6mSQHkfceHQusHTc0FV+anIhOm1/1wef6nS25m8v
XpcDv95HNbya5pgJ9N8xLg+av52OY9vucLURlQ+XL3GszgcM/3GX3W9TccbM0TA8
WBh6Xj4blgh9Dr3nP0qPbOB1CeWQqR6b5ogfp3oHUZxAOj7nU52pQsTUUE4lJaNV
r5s5/8Z9OlA6HXrDIeLLL5ObRSTfjQ4MAR5ww3sf0HgippVMVOEdAqxWVDINuhA/
eVPtoeI4Au5fuDm/kbf2pHoOQxijSbl4ih9/mqXJFXtULJaIXeHXMefOfdPEaI+i
GUZnJ0D0bG9WbKETDVJktKRzOEBu655PmhUWXQBY+0ZEkzFfRw4aqdvYxNuQmGx6
UN11T24iPHNb83mG3QtW7VLEtMcYiBGhm+1i/Ms2sxaO8GAuTAJaWky6H85PFNfJ
RccdTO+e/JjkW4XHdN0slACTRLkLwbQoiv6Y9RFvLEqFfgl7pGDvAEnIh8ohafgv
+6GiPQo/Jl6XYPSAGGNU65VidyOoxZm5yRpEBkFw29hoxU/X1aT06GcmR74KsygO
o7XUqqlyDhOJcXppApryMFmLGc/UDS8RnAGD2txzSrJRHrwkLCCa9xe3XrQ3g+fM
dKJriy0/0mUD3mdwWAxKpx780Mj/JDVvJqyclhLhhSNEBL5YfcmIy6X/1JbNVkWm
FxSx4ws0jrq7V6GtBI2Fy2l86nD2MLRekFVvvahjoPzrwkhgAAxWBKWeemTegSOz
0yiOgBLw6uQ/hMG1vec1xF4MnSGZ3F2JsAmAzt1zZ5UD/KPHUpXcwlsJXa5dW2VZ
PeGofMRu/zOvsljNfX3nL7oy8hnC280/jY2zeB4PT+j+XOrd2Y67I7707QuYDyOo
Mo22CYoKiSBdEu147kMALxvInuvFkvFZdiTFJHXFZZ0oTIMKXcByWTUXXxJFGb6Q
/TcBZ5Wx1lKrfEukU3/cZHJDEIy1EFTewumdIKuhv8DPDDXl8ZOjZ6cnqmMrLkPR
GHd/g5yjsyaCSi6ZiTtMFv55jQM3DWfOYaj67M2mBYonj7irRoyTYRIUWN2/9VNk
JxOiLKQh7atNVdYzC/0JkCd5XlNAJAgbQm8QXLioxMCIssBiFvtXayLKs0ARx1Ya
QbnS/6c4XXXuRkttqKt6ClGV+hKQbG/wU2bhJGQdNChoDfyt2vDCjKYBJFWdz6P5
gUIySvDMxCC/AdA0zGqxDpg1A0I2htph5APwuA4hi2tt3fJCC+jlfZ+2cHNZvYu9
nEpdJgKaHVrcXwz5LpruBMN6mKcRq3fHHDDVIpqtUOtdENgXu5HLZAG4fCWb+7RM
hcR8xfo7qgDM0p9ZelrDHOKrTElfA/3XTm9CNX43PRVW2pDoZzBG7umUQLiGBZ7z
UueNkrU1H6yOgavHFvQz3J/sjaYZ5U/5O7tZbjSCgfCxwDFNU2JqmJVlNTvC2MuO
KDk6rPIrbP5uS+j44TTklC2odznq3uK0IKtT7PZ+IGbYSp5aHU0qg+rFq2PJC3Wd
NvjhGsEjGD05BudJFN15atWYnpwDnB1NgezjTPm7X0gk8WZPpWUEP2iRb8d6X9ZD
X4kJQugQVnLUPVIvWTWarM39G3+XqzcmWVyUdpYiJo8/gOQjSDdA03scNYI6RDXf
PQyWIHVz+X4eMOrXkiEMqtQa2+rSgaqarUfNUtwVfxNAoGHe6jsYfJbYKRpszB7b
KZhmu58ccwTtgWEKISSNlVoZinv/oyiUWEq63sSwwP9q7YQnpZvtDQI9QYURB9yD
9izQrZR7OoQFi3jcyruaCawUOP3RO+UQcuvWT0tqfB9q2LIDFLegKXe8a3YtDMKa
pZieg8CWUhMUguuCKwW4Wb7FeiUJnVmdJOlcDsJYKlkmka4E8bRRFN38pm5TCum/
T8pbACEG6oLRioZ+vV/D600jgLQBz47RdR2oO0praQ/WEBYTyrrv+t/pP7gt0U7Q
sUtOO82qNU6NXAdhpvPvSe2o9IAOiIR9KoBXefrfMjgJC/CoqymcaLY5lgM/N/QI
Yg65pquwQoCDB5KaQKwvrTlxEFe+65GXBcjfZuuC5Hk22NyHxfiRVxUCIZ44dnOk
WmWKSiqYiGE24NJx+zMCDHn1XifJE9uUCid8s4pa+4rojm4k9TBUcyPnSSBbhToA
/9dr55EuLZCC2rGDqU6FJI4ZbLGj0VGHm6hv0exxv7OwJOxumR8+ixKVzStfVhEd
iQvdjGH66crVYGrIjVNaaEjCI9MTS95cZbm8oiVHiDxNkUjgBKqZSDjETDP6fPyV
GiJ6YxDXW7b+0Npu8EmIjoGOvlF+A86eF4T+fvTf3V0StAytAHUmC+j/MB0JZcOy
JWLIknk+7WMQidOokyTFYjfIdMt6jHl1DODCMorrvqnxrblQc8zmZbxnuui6YP/N
W+yxLRBGRdTuwsdCmE1xsEru8oNqBQF94P3N62bjTPw+5WZ78HuLAEWWM66VhAAS
D+EoTycVrEeHBLMPIETuyYHluPewNYFiEM5njihFq9jTfxQC8XBNfkmkwcOkYgqd
6NrO6eST6/9tfR7jewokyB+zF5YX0yMDWdSvdXwlyKfwV8YE9HaAmbmaEIlkhWoC
sEJmUJZCJC4rBN8hWFgysR0P9I4kDoGu1cjsxR6EzeIFkzE/Ca+yY3+UINgAtEG3
NoK1XRorl6+eWn4KHKE3xDHBFIX8JornEVz5klpGWwDN1tK5APbm45cE7xpphcdz
YoH4j1EyzYdwr3p2e/kGIpJDysEq6ttidqgb9PvaSEnjnlZclRE7EPIu3l8PSN9N
pv9w5iWiOLLmJAd6Q3uuux4aO4OSzPTxx1Vp+RKEXhBFw2YbuLkzwSpaiMMHMbQb
P/R8vJnisQf3asg7OZsQvqEgZX703RxnIZfmOIsK9AwgV6LdX6TZhTkvPxadsL+y
EeS7EVViY4rvjTbAs8uVQ2hOHhnQ7Bp20eMdgvlUU3LsG94SYa4XvsS0uBYNp0/3
XIdh+cCdOTX5JGqH8sBPwbIUeLeiKJ5cDrOPKVSi+JTzimFacT74M3Q7ZyOuHRGM
/Gh7VMYH3gDUxmYYXnAeLxJjAwAOUjZSigAvToGETNnJ8oDN4fEyBX316PyNkzkQ
7keaMZ/u2g1ajx/szHTBoPqiWyAeyY4peZ/QFPPosgicnPviABLEY9h+9I+JS2vi
BkFX0dj9gJU+xkbik+mMEXwW1mEAa6hJ4jP5GPrhixUoAUHzMEY56PaPqSDrgMvz
juGOj0oE9QgKI/g8jc2O6dNgy0e4YHSu4LkctrsbQjiIkMjfDh8WUV6uPCX4JSzf
uKqcvFX6a6KKmAalpabSDizbb2Sli0wmBnYOFX5NBetNk/b+enXQl9INYD89RMAz
ICPGivC9iCHnVyBbDw6xbN47KRHESw0kOtVpcY4lOn3hT+VENhf0FTpgSJ12drdp
oWCBCeqe0neEKfbV7ZDKmvZiEjWmBaQPO7uVFCh9EsqZA2r/kFvkjcfpwgV4GGjb
0kXM7IFyoz3GH+QHhviZPq6Tf6I3ao/uVDaMm1Fhypn1YQltfRqf5LyV7tDsLCjr
ULR2myUZNmMjQn74NDUbZiJ4kfnz1M2kwUQ6FDeHtMfBhZBHvEs0hZmoIS6w2N7z
91zhFwlv7oLKXjw5Fca8Xf20X72z4w50moWz9RrWoHEb41ztKGuTZIpDinL3cO3J
P+UwJzH0UvBB7E+VHZ0SL+wJ9Zs/yq5x5e+tggLFf9dAdJdLn/vzpvDDCUSmnwbd
txKL3WlpqbM968y/e5Z7wnz0XHI9W4FBSySxPBp0JO0VZsgJs5ZFDG8Evk57Is+S
EQPS3dk5waHBcHHOlWSdFYbjrzhIJ0uJaQQLEI6jaq77B3CC6UNJoux8wMr45BoN
kGottFYTRChLwzLk4jMmp+w16Oho8Dc62mRUpXUz86QA78pwOlEY9fms7fuGbmyf
lZWfdvUCqSnZiXPD8QubuB+SxW9WIfPBeLQebia3IW/Q9M1Rr+2dsBIr3WuIDDAb
63aIfgIttfm48ZhwHP8lBsPibUXuFod1QhR+4h9nl9GQWrs8q1OTZ4XIIGZjB+7G
PxsWKsuITl9/pqrAiBDtSO51l5IEo5/Rrq+KR6EKVuRL2cqwNRReRAsKrmSqrvYg
BTxQu8g+qErWDzwzudOR7ljgQcUF41/pFMJV2uZw1FbnxGMUOEknHdPp54tV+Tbq
gLA5eYtNXiGupZVzrsWRfbOGq7XMU62YGLr+opmuF6EHYZgXn/zqtMi8U/ZKIK0a
9t11dLfuoKDCH3tmELPmllmNLOJ+ONS8SnBFfyp0AJ/RoYnVO0RgsFNwa8oSVUHL
lm/63OCkdB+k1MCjOJ1LPS1w0ayMB1TG9LxLjHEDS9SbX9MmMtsnw1XMlTmRu6WX
Tsz0mWRJR4nXBmlfvnUHom7xwsUErGIMzN54HJFlEzBgl/l08ziFy439agMxsoip
wMnWTPCwpm1iPPq0pvc7q9TDwL4e6l+1JQL8pAUH/dkwFBbNLcitpTdYe+MXIVYw
uCLoNNfV6AGbGmpo7YN5ilZPZ3TjyCse0ImoWHFqgm0iXBibRsnIO72xrPL6/bAQ
BwbiHqxhTt49H3dHXNvdn5lb/q9IaQ8Sc0Ybf0R1XRGSQkpb5vRpd1XAmEaHZogx
NCdDa72E/ufoLqt0XkMK4eVvI9JVEkMWpSFYWm+vULWTgvS1VqoW3mxSnZI9Xbe1
PGje0604yOjDMh7xq/Wd3PcSDlUHRLuGHUpqzki2gv/PLpW54p95lvIcoyWISSGf
oljBLNCqhSOG+ArLZrPR0Km9PfAxOJ8+AjMjj35RPAj4IYEgpWkUpezN13ShbQB+
0v7P/qz01+bhvzXg9OctbVSPHs16bHz86Ej+CEezZtn4UtGa4i4BSHDkINvn6/zO
5kyxShIV+fLljyqhAGLhcKWZ+uBkOtpIpJBtNs/cdNSCq7TaXdkwU6kG2NZP0lju
sMTndyzWu3WT63OHO7+iQUFtLFugCPfAes7SJ5yRIboh+uuPBQD0FFt/07JCSDGJ
tWuRDNUWMHt4RcQq9M+LBM98oNzfTIe2bFvw9Y4XItM3m4qlycRm//wgqWDlEaoG
zIecz7zAUE/g9pvpxF+pn8dwmo2C7OS52v/FjKY2h5gS2QPw/uLOqYtO2O26cl/B
ns01FzwaGmv5IxdydEqg6gB6Joub73HKC9G3jVbdq1s5k7menCWIidrvCc2MKbTn
qFDPuHq5IT/h1VBe2uENlX3H1ZCi2Q+lUyiFAhtrvghqAV/yDxAER1erwEHca/n3
3qYTmnpn9noZdqwwWTH6GUTKWk2PqUjWqc+5QEbkKJGCI4FBuwAtIN0nq6R73TnD
+NmnVM7wf/khLH4OnYmr+8D9tAuh6alze86hX6dqi3C4a554cOrQkNv02Flh8yJk
XT2X1H0eG/GhvinSQzox1ovACgzXp1Jq13BkPxtcdeTFRgQRkOAI/7crFc+9fDuu
juHzgyV/qLAwZE3Scn4JvOJus1Pw+9jogYH2hxl3xHfAElrat1AYcmM3bH2Y4mew
S1lLQPM5fOUDn8Ug3ghqSxfgooBw6uAia7bvSpxO7cOhiMYgnbjQXXf6n+5wL59y
ra1gL08n4UkUt/68QPaK1NNbxuN5Sne5UQHkWvIp8ceMYYlrFXtijK6EB4Ut0v9d
qyseE9NQ94dDO03sLoIA0uAQLN4EX1mVxWu/JYL+nTcMREDAmV0M2ZMIW3423nzR
vVx8CxaES3lNWm0DcPTjL9/elWA7xU0aQ06BjD3IXwbkf74BX9TmqzoQe6BlTo7a
THFkTUlc8+vt+gfIlLiUCAjy7rRef7Iu4l4X0BobGrq/vZ7bJBTzIKx+A1+SkoBX
0JgYM3YV449qTnwKDtbf8KRRpmrPYBh1PfyXzGB7tE3zFZInv9/lQm2/qFHMVhQJ
5qRrUyWf410a8Awgm014+m02HPzmmhIPlHCkjoSmyjJWWZ6llZljad55eil2f3Q1
HFuTTrQ5bNancZ2CYdVWVcCnEWaZVCDrMTLDgfBOVehyDdjavpkg5pnI4IqZMzdo
RE3o2SCrXfUwNicooLCZTCALmmbYigObOcMkatAy1dGuN4ercUuHhZ0aALXvUt8s
RB66YAO+bTqs9s6BCv+iM+chIkt6Db7PzT9Uv/kRT81az6DQMEl/QHfxwg73lcow
02CB5Q4BIhzVgfFgmr28wLRvoIEVp8oH06o1qspvLwzw8ORquVNBv1DQuf9dCYwJ
Zc5AjW1vJXDvFM2/mHfqnsE8tjA2L8zYSpWmP/5oNtwpJpMpoloVPqQpXvKyf5r/
+eA8rzuT4nMlDPRP+jV/kYhwmofI1WgL0Pvu3vqHp8miQ+RyN2eHe25w82O/VKL+
/n62JDIVb2WBsWj2/GMCWajtcKAT9bG4DY7v93JC7C9mur8X8XT7DkVyqevbJEaB
hjCCdIPYPj0+j776G+a4MhGRAp3t35OAq+9TSWj3OoYnaC3HhnqCg2QIfOX//iEa
LkqYdnbkj66NOWCfiBAj8+SHI0joskxtmBieORu+eYz3PUBhkYH4YoL7PG198qiO
ZD8NiA7vAGA5pX1axWwesW32aoN1TPM2dHPHYx0Io8Uhm537yq3UVxtxocYaRkCu
JRrWzCgPPclgBm1YHubCtEAV4RBBftN+oSLZOjwnGYU3HMxvUSxxfgwsuEtMi1Ik
bI3BdxX5o07e7ZHNEXWFvJBzWRqW3aPVcceG2dsqJVTnJJxNLGpBOgM9ECWM4mHT
A35UPujOZQybfCSMiIRHTzMNzKOPUsBvzcwhZWBjW8L/hFKGr+zEw36IjX9YQoKF
n7SJobZjwqTz9ODMp/tNSXgiYR1DKl7xJYPG5JRS1sMZpOrZuMftLImY5g1IFRUw
5YcihY/FNXRWmvjhy5qoiXJU9zCxnePfubB5fTZqmfkNLxecR6e/oeynb0pLbAHJ
MKATCLqJspcdZy7e7bUpKpzF86Ys20P5vS3WIq/l61aCCtxqmPeUoHOa0gS+hY/2
+uZXsYrCQAAUc8kbcgNZ4lpJoVupOW1TTpZOODU4xSeLio47ItLWFhSifosDIbgk
BAwDl1lqYO22eb6yqN8qTo6KzLyByY6slrIjSSyPQYxzFFR6Y3sQuQ5H4uPaEx+V
VkkIcow21s+GexeEtvSp8MxCdSy67VBStDC9uDE15xXm3HP4iHoGBCjLsHXp10gO
1VAChjS9723b0wxxM0ZWUEObP5lhJ6jAg496Mu6QbcmSG4rN4HltdWYE1Vx6Ijks
7nUXGhe95jONgJfD2lszGdgRq46lj8s2BUIOGsrSKVvWK+KGPkQRfaaNKHgkMvx3
KkxiDHOi+61uCFFIVN6myEgeJsTaEIj8TVicaBBvW3gNBNZPcUV9yKm5o6efsuXK
uIj5BjxwEh1dKsewU3TTZkZwpFgJoOvQMD7TZRMSZuhQycDDp6kCIaTeyfHLpDNl
wGFO+fhKCO9dbBASJE6IMVvGrlwfFIBGOWm1nXJvccxy7gcljgJaKSdqo+7Bg5oM
LLEhNfDV2Dn59c72/3LykOQKZ9AufcWWrefZ955PNS0h7Z4mmaLnZx+8szwKNKDm
0cxd1tazmJlr4Xe21kKr0HcExKTjiSS+z5RerYxDyDEEQ3cV11z8h041p6EVpPTJ
MnsnSlSbdC/d98Afh0nt9YRORsY7D/kDkGxYlRJpbvHfkt12tuquXrIU1lfdeJhj
nz5bR2gYogtMDFOfnYrE8AN/YjCdVTbzIKCfur9cugl2BmdLk+pmqFlPRGrHSX2D
Y9T/0n4RgHzVEMsUH0y1rdXEpgN07d0y2EBXBcmJwSgt9EdyzI/gkybeuZufvaWM
PHyDn01fAN4Ny1c5hxA3Cm/HutgAKWyP35JcEFpdfhHkZIaguT2VrZzZrbx2midf
6S8WVIyWusx4/TasvjN7Thdz9vGq4qoAypWxqNwHVavM41OCbXXCldNazQROpvEY
RvbDvPFuhNJekqwSVhkwrquID4lgslaphn7vNJM61IeiNss8tbrnK4CbzjeFSyLH
Ti2Jp1RtkNokJ6KW2NXG0sqKYdl1qT1EuX7Lk3Qr60SIh+PGNn+Z/6Rv9q4qSiQS
jPXqiRqqgWEFsWjKCqM3xUqrEVQ4QcQ18tuNpVvUvm7Z3JzqX7hn2oTCRdfw7qWb
Xd1g5lav4qzDRDtxVk/qe8yvf1xY7KneL6ixTgF8DSWQVFV3evS4YgONTlnPwsu5
i63lGIJDdLcJrwl43qpVIG5gui9sl/R4Ay4mNSmXn5J+n9kT1xZuscCz9ox5UYl2
sBFmme3vg4F2JZfnu6HXV/HKb1GcJxV9Xc2U5j2WDBjI8etQeJT5W2qLajQH4oou
vNjF3xbKaIQiQFGfoAjreR1dFjkCUtQI9hNPaldCLxKDzhRyvL3xa550Cuk1L63d
rFNikMKkLvNSOn2ZpgXAXhtSyNfmmoaucw7H9bFM5hONj6UwL5U63jgrUPFD+lIj
HjxyiMSFBQF9eylMkhEs2BJMAkCWgNjxx3VyitUpP2b94tZ/xD0CFKNssNkQerLV
0RHInwN9H2ff5CbbZkJ0EnuiydwAV3eyV3OMX+KSdimlxjGEz2YduLjFgHv2kGf6
CxHep+KOjkjnnENhWGDx4hEvHAAx9cmpO0G2n84rUySqKWc871Mk+Z0nRo1aVrwI
Y3Ag+aEZFefXIO61wa7o9bQKzXNURZ+JqUxRYLqL4pOBUs2fa//fS4L83wBMHVy5
yaV3OfXLR4YlQzdmz3F/qyJzWMcxN/w6ebpfkYc+VmzFG3N+2Rcw2AfW45QfDQfv
HOEk9uajM+gIpeb8KK1NJJtqp1tSebWomEVqU1/zoY5319lTLT4kMb4hrGFvOxKP
BE+9DxT4wcM0fwqbTMVhrFJ3nV244WRtyfLU2D3437XRLZsqmoeY6nQBQ21R9Krn
BrXIIj++Raw9IQM77lbqJR0giB0r9SDNOTHNGYSklxO3AE+7Q5iwpXw2Ur/843WT
yh+wNElt1WydYxR02uux+KdMa1ArJOvjwPV2umOxdv+0ttJbjYTnUJO8Z7PIxxkw
yJDOiGHSEKXoZ8yT+hAWWJqhMLQq0QTmqGsY2XjCH9KQJlJL61JP5PMhmpAJ04Aj
YXACw581RktMM8fOnojjPzJqU5wVTjt1fOF/jPkK+O0fq/t4Gzq7LuEJ7Fj4XikA
jRAgAU850Nxm671D/GDPcZErlqz6WWNwE+ddojd4YOynhqMTemmPiG+yN2MR1zqq
BWBs3kjgQh3OpRicGDwsO4d0+YG2bgJRUcp6DGu339gozEBTXI3RRYrjU32YLuxy
Z398xMFII1xSIOVmt4XkicHKZRdDQW8n1B3EbRyYDI3VCcNV0dH3ZsFb+6LnEkjN
N4RcGD9y8UEJAdCTvhsQBH9D3vg8gJo8yeful7kuphl1JX031TlStxX1K8nrRNQH
bXI32GlABLRm/pNhcEAasFz1McBYjGbDTACi+J3TfPRpl2qyROJIkOmRrK6D2P/K
r6Tkc+Uz97Idz/FMBgpQKC9KVYghLGM7BydLkCIS2i6DIAOrOFNIlsEhMsW/L+x1
FB8czKmVcj/aimlW6V6ror0n4orbEMFPh/oE3XbhmFNj+Gwkwik6N0ZhcCxkTTb7
CCmlPdRSU1CYBjNva9WY6ARMOuXir/xOth4XnuxSSxL5XtEMgJlkoK+M/pDcEcDT
E0rQ0c40w84+bOunPXQB2ryWmDHeCxOU+RCiQCnRp1aAMcDiy6oWQt48IY6tSWLU
jeRZ+H6O7Ebj0mh/TjqlyrlLnjumaiak+7gwnbAj8ajCdNcRdPpxLp1ZA6n53lCF
HsAHdDza5qk57CMmcqla+nz/le5KK9x8jbPg8gG5NVG8RmU5SQecP0eBFrp/Gnns
Gp+YGmmNyRhippGEk9LnACMWZAciXfBsYGSVGBHjgcaNYEg05b01YzoKpAzezNga
oI/d25S27/dvoNTjjjyfA5uIjk6uztA3K2J/OUgNU/QKliZNtVqisZ9QKf/evKs9
9w8qxu20ZnF9JN3/zQUNc00kC4fQSIj3nu3RXUWp3S4V4WqR4q5Ph5xyWs+EfdTp
4xFXYGp5rB834ervBfNoJ8dayWh7PwiQZO0jC8q4SJJ7rGdsAhkzqpG269t84GuO
nXAbl2cMF+6gb64O+xz74GaFWf2BouPXL9XbCYrZKxnj/XL07s4afkwYxcsvCz/3
ejX5ssTabE/KAmn58jGMNjeB2AAHE06TY939Z9G9oOKrECaodZjcvTns5j39OTb0
dYWbNbAPZpfZ2ijSnZYdmWlx1iBYwDGb2wZbS6pZ9xrwAwKG5/8uAB9RaLDlKH8C
YIDdrwPaAm/FFZ6ATzUAw9TlA0m0/Wdc8qIyPExtiqajB9AA8dfKdMf7XINtfI+U
kDC3ayHgK7bNANZgG5iSGPXD+uXMFSNohXaoOEiFjhqJwwTqv8H95KKc7uWE1ukO
SFlkS07n/ZknRCyVYXrQleIYfU+laQ2TlP654EpRYVAP6c9hwTo8lqR5sxLmeMKv
L1Lwn7skp6QKggDF6JKyiXk2A6v/FRQ0Hl6DPPXriWw8uPWqypmtviybCIdkr4nN
A326oBerBnJz1+RVACZ0+LwimsqHTaNrDLoF5qOmOIiR6+ix99sGiSar3B7r+tFB
Q+PoBd9XVh6K0MbLpDJULykfqusSG75DOILDDVrNe/TQ3YB2Pavh0gTB19MIkMuZ
A8vyKIftk2B76lIomYJo+/5mFbNdCNmEjkfqynw7Gsuvdcg9Mtm1tRUYo5vrCTkz
ucUMNNN/Ak00/bDmi9cNggCgygkmvNvWa5RaeE/3kLXFkxMnLGn+Odnyo1LN2Qgc
FZ7/VmEL0fbxH304I7zddInsENHS7qIzMGInPbLwk0mbPAK4pAMqfCoPbM2pt2Kb
19WhAZCMzR9/Aqh2iXuDCFV3/9it+wxXbx+H/pCfWjLXJzUJEEE0asekDHdUgUMu
7+j78xUbiXnWod9v6kSzWgPo3VlRi+WS8Ln2UKT6vki/n3ZGSeP2z0hs8tcp7qd5
NOzc6eZ2TJf1Gr7FECOlPq2FB4ibSMSIF/mcvtaboWInJ8n5zUtEjUaAJrcAVfVN
FTqedaoF3uEmQQdAYfvBH+It2/ix4Z/nF7L4AFxmdXVXIv6jYr/1/PtDQc+xW07K
iYkcS0GwtvnzrIIca67D/V3WPI5fCn5wri1WvypwZwDFmUAnPgfENf91ESBDfk+c
nnodRO9eDMEHUIRAbJWLBMb+uYJEPiWAeXeRxR8nmRsncFCOTZKKMdIjMFgCzvmV
H952oDmWfsustMbO92yUDzulXPy0dkGmi9NsPa4AzcvyRnUhkGieZRzN7xcba2a+
W+b6L65YzXe88azMYNa7ENXcyOhlmzp9yph5SzLTgmruz3M6plu6Hku5F9Vzt1QI
ky9uOxwukz+pJstpMZK6g1oSWKlDbiGNI1NJQhy0gI/uUUs2RmrZYxbc2DUe3q0a
qSrKr2LkoVQZh3EENrtcXx5Q4XXBOPlLnBOPpP0ySVbc5zCpMUo6y8jA/QF0V1mO
NUyAzM9o+qnmnvfbJx3bCQ2pE3IJ+hQ/x34Gf3KXxvynoxcNe5l8EK0FEOC0NWsb
1Tw9G8QEL4UOvs0ktjJQkLwR4N/7IOB5AFeO27T8ge4NLGfxgOtP4vci4bsILbvR
l8QpgJFgwwwtRVf3HV0bN19oTthDR3OpNWpCxd7RSjgrCnnHxiteyzvcDTMmYrZt
nZ67MDI84GuVT8Mkhlrv/9pcqALgekvbuI10HuX2Mj4rS/YHfJ4y23FU/wWMQvjk
tbE5VXqGDZofC1cuFlnjN0MHlLahKf4TBFzv8xH0hJNcaSZugNrNBE1mjeN1S6EC
HKSAbCBJr18fmIF6jGOoGl5qpNdVJsXzzqngUC7tal0mkPv6BeAiO8X0i32JthXv
NJxgNwGoTZf5xx4TNTOlJAJFi7AEqbdwtr+pgEhfufVxOp/RfAhZdiwmxjpfgk7l
AuUrfmXJdi29XkYxRBS/yrShOW0OxufQOwUv+22aJMoj0YiC5PujD3rweseVOwf/
h1nVb/WL7SlGB4BrSXEupIxPbfeCWnadbjtAPmg9DomKOHHlfqcCaB1zAKmIo0GL
7N9VON77Zd5LbYZxi+fndOQRXvM2XT0m31At2r0OA2RBIDQjnZQbXBgZ6WnSMHpW
ioPD5a6z0O8zAZQGoyBQ7q5RRCUQOzD/g2GmhNW6P36qYzfGiQQo37aI3gSUjopf
rBgikmrWV7swuzlbZH7P7VeHY48GSQ9f+fYFRxjnDFGTCYl7wSm30uWqiy/FxWuc
nqc/q35jTnAX0JTwt98BMYOZc/9EiZeCoFyPJtIZq1130KRxy5Tc2m8JGL2hxwkA
ZvXJkPoB+m8N2+EYoRNRI+cFCmpIutniPVrTsd6npMYW+f7hTe1qBaogI/p0KHXk
pewA/INPifeYZbA5T343JZL/he6+0VY2YMxYhL02ICM5hK+gzX84Pzkzzksd6YnI
hwQGgg4O3rbgu2SbNYRTtp6+Tfmz9gvuQzp586k7kw6gBY6i4JqBC3IAWy8cauHO
YhiGD2BiskYMfc+agY7O5z5vuEeeU8Y8n3vZ0fT9GzHqY/1eqSlY++U29+5LDtXB
U40stR+M3K24u8hgMi6N9sB14FHti0r9vQCJBcTLuBXZWWM9Hmgxc9D0v3tHLW/G
D8VWFJiijswJ7lCZRktw+GxcgXZ6VprHIiaPqKMJy8WYv4cDvp8Fl4yREVOVfufN
4H6cftHUdLTkaC2SmjwJrZuuJ/CoeTrQI1N1oyCjItDOQrbPkWjL8siu0ZOdLNr/
oAu3+kXE7YW0IiKyVSgOxkFaTA50fKgSwQqGjDSNLJ66XOD/V8d8T5aQRGysgZhZ
OBtie79fV/DKecMpv1yVCvf2mk3AsYCmWiMQvGmKtoMikPIm2Z+XQi3ha3R11k1x
LVfCSRh4WPZT55rDxiFiZ9dbN+Pntvfjb9NxePwXSy00MOSqLavftsO+FLGaI1bM
pC3BqbdNzAPiigkgjk9Gs5O4npQdu/WpNYZ2f8TbOe3qvUHUqvMmlnX11O4oRCSU
jSp/G1VfDNYv7OBG6kx71pY7TzYNC/N+q9W5BAnWRRoDjoZpBDkogYFnR6JLTD53
FR4yxLF/P+pMWk2A01OrvkGIzXjrpfaNPg4Jhh4KbTUrKunqUS8L7EAs8J2O7K2y
1PnIqJRdh3rq3MI6Bsn0fr1k8h8Qf7TgS+35Mx9aSErqAO87hxTej8CTckHE490h
VrwUY++g8VINFU7RW8MLOKRqKQ4JDtLQVZ7pV302Faov8DatjCICtjNt5KGBogcO
3IvEv+RC/DNE6J/ZCuC47fueQNtJQd2aUCbEuAPKRnvAKMBbv6VveA/O5GwBURvu
xd3Sn2xaonC9n237mwHcJyYeHNjS4t93XNLChrbGy9TOhjUfMu5Qpd4UUYDo3g27
hj3kj/RZwEmRaUOJ7LhV9Y7eHa2iKcI61MhO3naeIhES+EmHhY4lZSUuyMIdvPGv
OJ35BMZkTbdpLjl/jUXe6/nOuBg6B+l4LcV4eo+AwQ1ucAMCyqu9P0Vel8zA0Y4n
L5VLAMlkjzRmIq+jbZIDVVWNjfUVKy8tRTvgUSH1Ptid3jLEPJ1ErV8+Isy44oP4
K91bTZRgvpof663j8+Rr1+dZK1pWsDz0DXuzpnOYyfhclD6yx4CkMoMhPcvzNCoP
Sa2m4Hw0YrbdLAV3CK5yjBshS0FkrnV5iXbmJF+0mNIoAQLG8hsT+R1rEjEKJe0X
0Z1SxWpKWi0EeldDx6SMqDc6olf5xh0Rol3wwj5qnvDCyrIy9t6A6ES8IOm+J/rJ
nd+eObORHibblIFxk1jCgqnaACuEuLfH+2m+f4jdoUhYhZslcnjupN1fwunVqlVM
dwqFLH9pI5traS2uj22+3vjm5Eoi7BKPclB7r9GXu5w7cPdcrZL2w/8aHPCYAw7a
bYqnJL5BVXNYsbEDLQin1ecSk/dbWSWpclSy4Nx6AIwyojbD0KsK29noMrD+A4Gz
BL+VP0eqLzzMNtzjkXChdlehT6SDwAGYKLcEsZdR3cKdl9zwkXsoLv1x9IrQKQRT
MIoVVnPDLzicQNtrPVDQwYh3QCXHp9ohCazBuqQmC82xrxq1pbfLbCZ9I6bbvT7b
nLsX7j+FbvD0u6ESGolm5yVsoWFYR2ZUNmP/0Evl5kghLsENB7H8d/gALf9yJWrD
BJuQ9n8tZRZGCjL71CsiF2Se/suYT8jHumMP1PuDqy6uDBuvGcApcsUDhtd0YDT6
5FyKgDoeJRD9zeMAmKVkFL7CdHI1ayRv6bNUR6ZuaD6sEfgsLHelXzdxVSnLIXs8
Yp+j+JX+HukaWeYtWEdhfvHGLaVCaOh94OjRSLlzrbEoPGj4QSiU4EIA7tX7GXfP
cjneZARNKk1nPqywO7SrNHqVUKe+2Y3xq1DXhi5eQcZMHhrTl7SxLEyDqKNEoyLV
ENCShKsqX8CUqQ2NI6Hk2SfVV+Vnao+wAev9LuCTpXbFibfmMMVgDfhs0kmdmfNF
p74bYa4+5MUFaERPsJEIC/j1xLGGI9OLrHhADk3Ki6Uk+n/S0Tw9cOkoqsyo3TR6
vuRFLcJIkWwy93Yft/Ym3g0BvvxrB5aYDXXn0N6N7BG64/xMudCcAD8O1T7E/ESn
e7b1FlUhIlu9vSDdl/wvF61vEqREHN9sfsr0QDL46nCprASgD1A+8ayyaKP+ORW0
K3D+1gznVq7YMrGrvyqcQry+X7wH9v1DaEYhv5ETKKSJC4+0zWirdC4mufHZ6lSb
A5tTiMgt1UNtu9Uq05sSjWR4N2VEmfYNemv5VAybUSM/hfPBdh9EQ0xM9wwTWYLN
PPAS5ur1NetrcGY6RbJ3o603vIFTbluE98cHvjXkTxvu+obwwJZSqA8NXK9XB3qk
UCRDk9kU4BgtMFgaK46a1Hpa03sx++65tyE2n8EjC+uVL0QlCW/0LS6ZKKBsTbeK
4WermMXPrLJT1n2vSISGXmDlEDUUGBpH1gVXFu5lTnGFoxbrL3p8TqxUypejrsGR
N+TOdnShFuX3HHSFpsoqAlChCUzweVvAUTEz4cZ7aRHaSiIsyKyw9zqVfcOH/vuA
ud//sTCzM6pAUC66kCmx3xC90ey9WGos6TQjOdQwWMvBqcmpDW/QbXCzc8SitSbN
ZcJB1yKkygJBJnw071U7LJXewQQlsOPURQxYfAXqg0oYcekv40OyGlAAZY5CXYzf
kGvWal1+YoEvhBEvHOKduxjdg8yvC9hvwn7uG/TkhIyLwzhC61jJGpxxAoJ7Hqd1
oozHp0K11nmrJOu3Ud7INIjpgfMiKBIbWH2pgyjPleNL6ZObbeTSvxisqPC+6Gt1
0/FdB2ILCVWEWof5M1ojo2oC3I1AFuXU8PVGxxgA9ROxHx6Re/R12WfQunEaP1za
RazED5/HTihHAbg3TfTk8kkn/7qpacqI33FUqfM2mdt/Cc2MtquyVXLONOg0Tc0S
W4FlCmFE3CGmFTy0VFGvZUGHjcY7QBkznJgj8KJFEusHriC8joMQvAhQewTKpNkj
jfbxGf3wIFDBvrHSkl2O03WoXbTbxlwgECFOIOCtJsPMLPj/jkeeXp7vzr4mOGeh
2Ct9+1NW2wQYl07jcDoSRn0B88uDGrpVWLgd1N+DrHFUX+2K8jbnwLzUf+bWH98+
BAYS5iNaU8AaZwaL3KBQzzLpGNIKa4TEUhu9j+1LfSdLMk0Iyn01fkpvKPOA1K+j
BUXeI16Jfc8JRS6KqyfRRNp4wuoVaTLUu7kPIiLtJhndnt/cyFonwIXvCbJVmhUa
emISNNUsvu+9G9TBXUgPQ1zOqOEH4yCrgB6deo8O5wSI2Ji1Y7Cogx/Abucfn8AZ
p1J3gp1CS9ddLBGXZM+jFGtyv0IhU2cAgxIhj+csCL8QIvt3ZdFSOkNFQK0Ojz4X
7aJdykJNvbgUcV/vxaT8JMBEOPT1uI3SOc7pCbt+BfbFc4Rqut4V1h9OFJoeDuCK
OJ/q5h6sROSABPIBDHCTA8+Eis/DNVGR28aCDZaQHVMuFYco6EDbyRYPnPisoQHM
WQAGkHZWQ40N+UGq7jw2DUi7k6mHFXGc+G5XCWDQRrAseBEWeSe1EMtLuIvhEF8J
rz4hr6MB911Cq+Zr5lzjy0KV9SLLpQyb2MK0s4t4BQTThmOu/SVUj5OxXFQ3ZEFQ
E/zXemIsSWXrGtYjRJamb6afVTHuwkEdhgGZIyknfTTBmxMuGJXMkL8p/5nmmqwF
eVRS/y+evLcLvw1BsDnHh8/IyOOYWXOOfDfqzn2MwhEbJYVU0KAyvObvKKDN6diV
QSCPMenMA7OnTDiBEd1ymwORT9Jic3KEkCNsSAUrA81cKNYUKbA50uUvs+V7UDJ1
5PEKzsWxxGhkGv7ZWU07/o/UpqEstDipAY8g+NA1bz8EWty8R4tVO7iyc0M9+MY9
w1h67nSlc9UVy/MnLYItxqwEnBtBCVqxa1sVkFYRcQyxEnRXZPVSSWBj1uYpGoyB
o3zYPqLdOqU66exA+XjyZxrvs032kBYhJsUeBdijx3/Uhg8tPSd4xF4moCQ5Cmea
sDqPP7MU+dUIz39iufPmfqL0xXeNhVvll+eBXlNQ/aToIPWdVvBuOaq2kht6N3fB
tFZZBShm/dSIjCF4QRWos7t2QEBaiXSQuSDgyKJJr6hqPdv9Ll6UwuJZz6lFTJyc
JuVIK5n3jhdOz05jaCwf6/t6sJQ6KHOu1/akDtk6XusXQyDJjjILQlHlxEIpRtiE
BibktrIlA9za7TqKYBK6CYrNaRoV/+8BFDX7WOn5UI4NHW+6J1JxV0hEoX+MMiX7
3OsKpKCwC7KUxqRmT6L/+OaxVSvYF5lYdI4jz4qacsl4BT+ngj3/A6gCG0IQsPTZ
nuYYEoNCIe1q+Za2Wciis+O8k0WxadNdOTxxoq+Y8IRsHipRC3V2+U45W50nlAeB
fjh0f3Flyj2cGCxEJWMb3Za2YATPBuf/3YCW3YY5BqTxeB39ZkhDhstvSo4yeh/i
F/8Ib+Sbd4bgOSzSl+RTGPwh7avPCmPEaOIms48mkYR58cnZj54GjNZD97AboVvs
aFOPSHCi2L9WejoAre3Fs9/+iY/L7zKCmdFVeOv4rIknGmjA6XNHgQuTmDQQm711
VANN4r86hAldrZmzR8fXghwPa5tmmuL+OOn7G+7Ji4LtPyBH8wB5QN/9Rebc/BB/
uBRp/YcmHU0WXl0s1ROoVp+3vb6rsrBusmnrR4wNa41l4FBb/G0nPr/Qii7Zf/gw
8IuloekhBVi0z4sHA8dl81uyFA5ad5htOeLnw6AM5MBeItYgmiaVEHkhL9MEcqoP
PSApgXuU7TOg8SnsPkdh0i58JHNoQI4gaKXnXOLlJ10OCQ06iwyixFxMOZHodGgm
0aD+LwKQkEQHie9gqBSd5vuc31/IVhgPXqcWfAr/bp15UjXbpuwq3eB4nxTKZtpB
pAUDA7FhqwqKwtAHvDZyFSNGi/zPUH80LntcbOGqe5qCvzYWSdVeqaCi6YplGUa2
R+pChySTVSTaBOXXBHjhrlje4rVF7SOOjFYL7DY8DMx8o3Rc1005iR84PQNvToMG
p5ZrCffAafaeXN4jku7Qao8zYVyBJryGcCtuksPj9WHwLBvY7f3Z12THb8ub+4HG
RBB0qdKQKDFpKyaHdHByUoxTxf7jLelRm5rKpoqx1Mt35s8pmHHXzfEvkOwj/Bbp
zkPLTX3GJbL745uUKn/zD7XKufclrLhp8z+7YIDsYe7QGqdgNmY/d2r8yLZvOwbA
bOPWE3uw/uNyKxPSIOGQ3tWQOutgpRtdfq59gXEF7MC7HFuew2rSJjQjecK1b9k9
6edTUV9ldrxHm47wiX4TwldhFG3xaxkUGDiSYxZGlc395uyxLBrMuB3zk053oiLA
vxT8mYJQGCClGjpYF/Mgn+5yOozFZNRPlSmbS6bOQKhSY5lziKzgmr0tmBnShyVi
3KOHBLeu8o/iKH6T1/vzJQjR6g8+2ArLi79PKlc9IbrhX+1EJS44E0LmPd3rMJaS
u4CsSjD2dFdb3V4UQ5ZAemK7kKyqjxIofEVj2c8s/lx52zbRBPgl6dEia3dJSzNQ
sdttR94tp34CzbCcXHNM+37GmyvHJXrtjlE8MpxmnzCFChjCFCHMZcA+nRM7tXMQ
yK6JocJiSYW91KSqSkmhzuXfB62Qrg0gxud35IDzzTo20Ib4HQMb6GI62CRdjo5/
GQI9HxXX7Nf5Op5ZpxHZwc3yMySL9ThGaRJeP1DRQSPjtsM/Bc2+LxLvIacRTvzw
WJLuK8HRfI1I8ImnVY1yWJYEWcLxEZ7rSssc5TqX/3/zVIK/O9DzmF0KZAFHvI6m
b1GURDhrc2ucXuGjVEE4XrpMa1tSLrdbkbe2bQx9MSxCAoh0D6Or772Mk3d9wxNY
jlGFkzTOYeFzleWBzxioh1xuXc8ny9llHBicGxOs4RD9EuK3AS1/l0vSfqziN0mU
cE8yeNl/Xgrx1farQZB7tcTvXxdQFZ77MQjkvFeApMYFDFOKNsZx9rsZkHRPY/Wf
Ywc9F+/IAM2RxQPHQ7KX/CZkr+xO+oqx5dzWral2ACiWGDRafqYIoMR0pu4HyT/H
84J3zlR0pakPfizE9RR0aT0Xc9c1wLsuFOUSERC/SlLzqkSRtWX+BIPRHuMJht5o
6p5ujF+Lt3mYegAXALWNDd5pzA2/A90eXgodbk0qGmwgvgnb3qR9iFV37uLqbp0N
jM8pwjdYljYols17xidJ1b7e07y9tS2qFa7icdYxuLvSydPGYrquAaq3O0EdmmIJ
Sr6lQBRkEwugBJDi9aB0U793S1dfQyUT1SzptPCcHDp8cA2atTVZWHv1aEfmB4YP
iW4mB+bPa8QiMh/jDm1MrOueqXwrXxH02DuN8ObwRjK/ExEVeZJpuFduOmJjoN4O
Ztxo5lzuGZf3WBxLZehVK+XQ5m9UbYjIHny5fltY4w1Lv3NYS2SRqk0fSHc1FOLn
UmjdAazgZE5so6Cwmw7nGRPk9O5VznWF5rVO5QMZmCwl+j1BnuRmAUzWysQwc+3s
j6ATfXtIuWgUmgDxYdqCPuGdH6xZW/F4FO1jdifIRIEfmN46BoFlMlhKIvrtSe/L
kU9DZIs/Y3NAIUcTbxem8OTryKOMk5xlrQYM/nhGPJavDnGuca8IHECHVA1klqRg
NakPuuP7xvAzlw+uPyVTFjzTAex1jVCSrYV0SJXA3CE7OQBK+39ciUh5J2lhIB2t
A+sjb+gbsDKq23WkIlbex3VYfb/YSZs1pFpBY7w8xQicR0fx0WidUmXxV6sqLeij
jrHE+ihV2kTx0onHOVs/fDn6PwIJEHxTVc4koPJgcoq6P3dvloWr6J6WISSIo1bP
AkEzydFFzGBKmOWSGFLCFxoW+6nIvaHLScFk/aiwjovRn4KWs9LPf94irWetiYAr
Vx/ugvkFkDbbkHVxTtT0Aw3iFLDCu6PCVN9YZaqwiYFfhP/+sfT9HCnTrjdkHdQD
6PPk+rYt2dDoG5YO3FgUkAcUi8wAhyNwo4pecNlqm9BK0DKgwU4ymr3rnk5ieMH/
rki0EFKHdr8p+4M2TYDym5UZo/OzppBSmOgj57eCy8lEMdnAFsfXZRZytxszWP+Q
3SZiihSd76ZjLfrX6QNxuxo/s4abJcITleix0hXCV+hq0fpeWd9amcowAtAlUpvG
Qov7EZeCPviAE4ZQdqKphePlhXl4tOWKVhrNwF9XJehzYKbpsJsTE056dQNwQQvC
O2J5LZ0wPzFlrIK3IbKvPu7Z7O4X5M8PQD+pXKKK/p+nAXVEo+fad74IVVsfZHKj
efGTqGwCi8VeW9/at0NCIAegqFJWnZ0u+oDHpzc1m+myZ0mYxJNYnKHq//UMtiRe
WqK2damD/KH+ENgamSeF+GKmRYeiKlY+dzDeFBZXz6/HB/tImk9397eVPjpYgaX7
rx05sanMtalXVNA2xvWjL0SFdZCHJazbLVDqMts2e5bz5GpAE3yaq53q78EOgiS/
n0/o2OovLsV07xlPmDut+G8X5t80k8E/+J4N6xuCSqvPLFQxnyCTVtP5j/qIxu2T
sUKx6rD6dcEwvK8KdpNIRq3ib2L6ds+d+VDOf573DWaHgcsVl75XjfkUZxpcRL7y
e3jFXOSF6rc1MSgaAsviinzczNeH6Uub32wMgW3zXgcB/7dpHvxeifjW3khu41hM
J/3FUFcsll2poGwengOwCxk6e7ZJ+4W65whG+8dAp0lkNaeYwwbfp5Kk4WHCXT/L
e+otrsuWRuN3to+D6x69q6vMJEwHHP/4lPE2yYfJaJqM3uitKOcZb7KdB134rfng
+CWzYvPh9yirYsdWIobVLTb4aUA08V4qluzgQlmEjCOLJ1sRCYaapEY/uik951qf
xjmZ6OQF0gksjqXuUUmWhG1hpgetyT+Jom5FBT8ITIXD1d4Qhfjncaf5pe8qAPkt
pysAklhLnAaKuj256R3BIoJ4juQkKmkW/MkE0r36mezq2gPv2KuiU2PJhLfKPAGY
jt0LSdSD/F0Axt4sAUVbDp4WDLz4iY4594RPf1u9qtPuTVKOU0kBDCRMvgU6GuS3
E8T0ylgxOyHCztSFZ1OkeUOX5R3V29895/x4fupQMY/Ku8VNZWgT+19kfai8qQ1b
PWnFjd0+1SeKJVPY4pBu+chH6bA4pi94rGWOw+sLpY0VjQ7OVDlRC3/nAR8Bvjez
Qdhuc5pjUgUxvfXyLC/BemekKKdtTzWMPH9tKSBQyBUQT03a+l8kPbqBgcuFvUEO
ZsC4HJw90yFNMm0ZGT7ByoqO9vVPIYEIE/W9yhrpVEVLq9zTvECdz67hYW/GZJTd
jYB/nJcBbtLaHg498rUvpUDjf71PrO8UI4ICDbRXZ3hJrEkQNE6mu1KKJZpYuaVb
1Zflmbx0jxvk06b5ZN8EWHQY0SfOPlK3NER2LqImE0v3jtXBXw4LPaBXS/8JFGrA
o3rNVB3S23YCFAQHCly1r06m0DqhyvFXmQGGAFEpqvzZ/043mKnB7LFHVtGyfOjQ
FhcV3ENfRSQPj8INxNRr74BYv76YfBcf/vi6A+Cn5vjowDKnVLt+qD3WOJHKSxgm
3s+YP3kqZ5cHfdC5bRJOaEf2w3vJIoUvgs1tLohrXSwy5tWf3YLjhvHKM4QzjVWF
o7sDlhEF+GZkTddSR/EpLdSfsdgc7PICxYWSisD4JkreSbGKe+uVyy8EY99LSUcz
X0jhgLMRqwtHZSugdzQ+dpzNf1q9idEzC1rX/+w2loIFI0eUayszoY1QhZwBZ7FN
E+CKwrDpVYGZoemWGBCaSVGeDP3jtvPrh1HkwlB8Z0JnLdl07SMkG2bSYcOukSUb
1zu64U4flqvYG8fqaW48TfXCe66+rBbn8HSf5sKsOwwPIACNuGLCnuTrQ5YKiTCs
Tu3jowcC1kahUVGl742xfKnyUAdVoliJ9VOYWnVPmwxmrJNSxqGp0QYPUrxeg6ld
X4BDO98GZxbAnlpvPh6KH8InvMzFIKlXCVDzYcVBSMqoNfbTXvHGO3/vTG5iBtX2
BFzzEcbib+D0VleSB/CHx8/KpqP7lq8Jm1ib8icZ4yAKpWKr50fIjkHbGygs0xLc
CYCqZl3yD0e3K/+GuxXAh7RKvmnE9OEh+uvDqIWgvsflpC1yRXDp2p8rQzh2FnEv
cj22AepjeMzcjZzcHC2DyAwvmvL/Fv9kaoiLU4MeegRfXCzX1yiWNO9pL6jobjPM
7qtYkmbQWiwFjpBAywcOYv7lcxEIh0hP/IQitJ+5lUaNoAjvqRQXfZEumx3t+6sK
T8GI+RkDgVpaOJxwtz6eT33kFPjbTRnBkIFcgKtZfwD0UuYtAAlzAVXlF4w/qEzK
DDWbebztGFkmJQvayf5otLV65iLLnZvJNU7WMKcWWCWF5krIhLVuJEFB1S0wsBTL
fVmVJ44o60J6xaW+Rtv6IZgx0CiLARejMZ8M6OD2dljRtYmRZMq/1nOnsGPGxzIT
1ms/2SGmOSHY2PlI0FKqhq1XfLHtzGj/eGFb1qxoiYMJlZi0xzb+SoBpp4/r0FrE
Aix4ENmpEojuyM2oLQExYbhbV4+Yh2vZIvOMZHEYNU7V6I3oFIoE/55S92ccmKSm
KZztMBwpLIRmKqImKxGtSMw5rR5ZBJ/HW+z13CFG0qv5ol1dxyDZbTHsDsAYxvgT
Jr97RzH4Dh1fZdCzr5qZpyIoWfmjbuUxK1QQrXVTyRS1STx08fMP+MI42AdOw+yZ
WWhnks8ANEjBW9zz/pOL9TPqJfslhCFZc+J4pii4CFftcclibH4vD/I2Lhh95ldD
F0Pqi+vufWMbFA5zLf4U5cT+ArPsZ2KFjiq8Bw5AhdY+rcOxeNiUjV/Wxwci/kvl
af7X2SOPQ2fgaJeMJzEHKK6b79Xw68+5PeJUY/ITQQE7Y0O99PoN0KwNDnGfZjqi
GnlqeLuIwPMtlQ1kGdySgQbf80G8SchBgguHAUw2bcCJH6dfMKXj7xK9K20iqHg6
AeA113QWPf05m99WCZXdfI1DbbIMZKVYt+5bg6qRJBOzoadZKbjKeA1yxoMr9pZ3
NPLalnWFrJuegJ+Sj9dcVD3quIxvNu4hv0XlawXkRC5T5WVEwUdgv50ewgFK9xmT
ZkYz383nWERu4CEG0ePX1T0lgDqh0BAmGahw21zPIKN6fSHx3y0iYN0GXgsYGQmO
aSDfL4um5EVMkRyMYc1GAEWqjsb1nitAcKyVxTJWbP2V1QUvLLjmPkrLU8Es+llK
ivqxRZzUpDPv0bPUBZ84wLtcadPe7e1eHHyK4J4ubCCNnlk7NzH7cXwXHiMns3zk
0Xf7Tvyxo8d90ugTo33yhBh3UN7f/QcPLgC9u7H4Qtx8zfBYXFWBlo4yDEsHpiDd
IPoswtb7KwdSLVVIxFi/DGmxiP5dQmGqB4NrBt+vs0BvbjUa5ajdTBi5NhAVulWg
gHAJdI647351s3RGuxcJYyJRQczIYd7UT5LLtmhhWRMOjXFoLlYYZxJdbgeyd/J3
b7yFNrjo51HNArw2oOQYfyTgii9oHIBsVrw8RoN1GYDPEppAyYbdmgW7KNSk7fMn
n5Q/vQwSbZincpqGkQxHirAXnRwSUlIAJWf0pMJgzQDQZYZMgS98/gEKDLeUkZkM
Ys7U80R2nlGn3M4LJmSfujsmChzBSbzooT+0oeL9jBwTrCZgzb1YSi1HPHF9+Yrg
bdSaD4lZ7N6jNNR3jwjSpdrSuP7mxGGmEg7WF2JjWErtac/7YihjA/R6u8yKK/c1
ogeLz2u8Zfr7ral3uZ3NlIAnTlKo/6uSGkT0iFgZtKCuE9a09LyV7V7B8vzCwoeu
CJudZqNkG+NIoQ0IcRbcb9vVAMGR6VWb2t7fJMvZbzIlpTg2sY4BsO5m7w3mTIwp
s1Rn5j74m/mwjnFkJKmFSS/LnJV6SXhgpUYdXaamNSiRf0kQUA4cAQ0+AOeU7QcU
wXmTr7GXAaAYWpsSSR2nFZKGbwCED3vJUGEhsu+lrboKXvZHjCKSdmRRBqWVp9hU
x+sjgHV1B7b2PL5UqumuHd+u5K79yoxEpYgtJ5A3/hiwIPkkKK1/rtbxMPIKIs9t
Vjf6AWuaUk5GP59QJQ8HN/M/9N1F3kgZvZEvAIiWMe7j5G6nq6/cCFhndvFxU6lT
9OzezJWOTOtwXTjwv5HG1buQMvUnfjRlNPrH6qwgmYFz50S+hK6cjUT+ui4Nd529
MCBBeQ35h6st/inbUDR3Wg221DJYb7wLK2RCiVpOzFTk8COCBiHjKv90tvaUx+9Y
5dZMWcB+I/Vfw0HDCo9wiknFqX2Qh3HjQA3CVIQAMDKqI8SK+p1Ulvj1zuYdjZaD
aFm6A1VIsToEaMnrAm+uyYPCt7ELgnUqv0CAcn/trFJXl5IHkI9WDaO77baehj7S
3A2+bekwvTJFpunIEHlGfvomcEMCMnurX1rMsj2sti8wQJap51tTq/TIyQeSWjlK
5GWXsp16JHnc8onMgYGBi7lU2MxO8R+7YwKAswgtmNJC4XQE/Z8gdD5iSg39rY9h
FUWESzHaJM7h7Z4bCCUI08gOS3qOp91lkJJxEbXJe3BUQG8QYAP9iFYHyld5S77O
VL1wXwMt4SNdgwY3+CrWXMt+fHEUaMMmQpIIjApiDnev+lvMp5Utf33aDSCUKq6d
yETswr+53JcAWv3EYUSaUYs2GsMLMuYy0xxwnzIR8KvitZYrNPNke8ss3tsIXN0c
6xh29P4XHttbMYHSKaGqaUZUy/wmbOlQ6b7D4MIs86Ujw0qGMSFN2cmhpg3W2ybg
Nv6MkUtHFfK6H0WwfIL+BJxv9TE/JnaAD36EOiK1/gquZdP/oKANgqBFnl9nfaZI
NUEwfpP/4dkgxgrew/HuqjpVgHJdTYc0Fz8XSXcKsNGuZ4jPy0L+i9KPSG4D7UVg
jkcm8Fovh5Gp1DAt8wgmhDJeAE4aqLOBYrzK/nqUZKOQxjj99uGMVwtXWl4UV6ND
mUDdArZ66NzVk3FgiH3f9yf8XPPeZfIPV6DvhMYu3kAtbXBVrXm1L6mrvXG9+pFH
ezmfxx472tKnltrIuA0QCD0efosW4M6tn26j8UoKD38jY2xRx+nHYa9ZCXz/qVxt
FO0FPl0gIw24ga7RUJQW3q6MmLzHLW9vFHjGpczUOZK+zIzX3LGZxpH2eA49sarh
X8AhwcO6EKANd6rgWCJ2UiwQ6WWnO6kea7hYjSJu3vONGdXZJJaE/zc8hyZ0PHTj
fEkuBLoVhZEotYyUTBv3ny7LxqnlnFV1LkkQH/zSaFuJ7RPEhtRRK64T6MoATRNZ
oTwi+3n4sIGUXXHvNAL0eX1c4fuOH3WC9akiL+KPCi6JA2dOXJOwaOw/FSGEguXB
1s0W9Ofmq/kPuUdXk2IksppSSfymXIg43t9jwzkCO+xnlNASe5eOnUbNx7+ZwyDk
VsKWfjBnT+reJVPJFymN33IV7VBbcaU08VKgOeH98sN1sO4VkluIK/9Lmw2ML6tV
53W0WcP0+MbQvjv4I4olbNrUXxO7GkgtshPZI7gV7m40/oTF+5vZRoLFIyOisQkM
UXRs6abBrl5aBFB39Qq+h0mxaDQLNgRycTsrNIQLhjrqa2Es5AvkYRvQRwbz4G3a
Sdm1QFncbSs72j7GhS5MOkqhPZHPc6gZ0qYgLC7XheveZKYY/+Bb8XLDxUG4gUJk
RTZEe9U6v+rfr136HQ9dC+AUaZYSt1xH2v4lmnlhqBuiLmU1Q3Mlr/xYJ+c/PS60
8saZlBgo2yIpqFfrlWdAaG/sRCMWAVLKZwcvwTk5yv63U58bJORd/2V2c4a23k0S
Gef6cWxcJuMXKKbG7H3FfWfB/lvf4i2aMrfjHVmeKoBjget8iHV7eL1tYnE6yH0O
2CgluukkuHYrjPB4OxiihYnCpaHi31QI+fEOR+3ugBrwu46PZA/x/HLKsv28Ba/D
kc3mgJCLtgsWd6eu/mjI0qDrbX7rhpuAlD2Inv9UAl0ZMmfHebTwjVzY1W0mJW5H
k2On34vqmUUYSuc9QIz+hB9EpaKlB5LNcS+T4NKQAp7EUGYXpZucNXBh2vlplbkq
x4hDK0S/rbDslmJSSD7+48yzmOeUACB4feKHnxZwYigHiB8oqGlEt7EtW4Vpo8Yv
ySV7A/MpB9uSQL8jn9WM3Jaj9dhPH7wqGXzxcLoLYyVG9CLyA2yDZGXTsCiuR5j5
60ShrXtn9UDdRZvAArG8g2TRsLB4dnEKmZVVKSiSsjPI1VcDAPpPjCfrWqx9fHZe
Vr2o07Mh9rVJWqC3ObJvlKvypM2DtbCzcqlwkhPHVTdrDFANVWpETjcSgSc7VDQf
XdAgG2TPRXTifPoDTtreVw7qBW5uFzLp2SNglWlJdpF7pH4XuGHviw8G0FgwTF5f
f5m0IfXd/GWtyzgfuM84TVVyJ/NUwiME3LIq3vHPmqQPJZaPqIZTU6aI/i0Y7NFs
FIs1g4xm3w/d2xLdLyR101J6iMwXmIev7ItOoYEixlU0I6xhz4jdXn5gjTFXH9Yr
1PN+gDgTIcjI8ep3VY9Is/gMno/en6fp/DHr2v10DG5wgYzRSj9LFolFNdxWhI8t
8Y5kgIQDLtQp6mVQIy4dZ6kSjeiE/RMUyZxxmfg1IkJfwFFzpZDa/1+ZI+EaFv5R
WkZytBmGnvkj5Y3qxVupaY062Z6kII7CcvyoxAAv/wT+f9awUIzn2OMaoEJF6tSI
mwNkw77+OnJxMPSxIFazc5CRfxDgCmNklqrvENt0I8mAoVHl/pF/2vhS9T+YUqcU
fTn0NQg2CXlBpWm9iMyfdB0UQeYGEBpEzK2TQ7USzZFXR2O5W6BMuXgBsgk8qrbM
pnIszE1mBXPK89oMz0pN0k3W3Llwj1TQrD7O7/EakwJvTLv/8RNDxmwActQueleF
28lNYDEMRdAZ45bfMSt++knVAYzfO4ZuBvKBtE7fJQBUaDm3yQYUXHHWwzh72gDK
rNjzGaKnF9FwL1zZEBvGRPNUeI1kPYSjfstGgARgUyYDm3hRTYgl3gnRH+x9kziu
7n5y6u02DNSD9Z+FgN3ihlIb0AvncHsSKuK4H5rVdvuAegDrlhl9zmWsw9PDeQTb
kP1wovMplbpiE2iNoFXbWQko68fVTm8r9ee2bHOWnKUhKxwEX8rwRkdwK/FOwAMy
HACHMsu0sGf74oEfM8C4PeMF1SrAZ9A3vpfChk5DSnRUmU5GFXSvz0JWlr7CWV0a
8CXBYkqu4MFdW1Zn+0GWszUwP6J1p/T13gRvGVMSBR4uGdmBfPTFuUtXOtLgHlxn
JTv14eoFM8jcr09XixKLegZO3b/Vis8gLKkfO2E08IJMcCOtutq/2Vv8z/Wt69FR
uR6bUQ6Yq5Mcs6XM5BQQZqkeHX9MBZKeiGKmKjGMbMNJtmv5M9wwXCVt9BZ9YU3i
FU2eKkGMI4zxVFjr1Ir2WZOQ1+Im2APteZZAumAHQAVU0cB3BNegTRbxeEp+aPSN
bjcUCB6EPyxjMy0i/LwdU/GkceiXZhf79NXCRxLlR2hF59wBCkvHZvJLuvnU7CJE
Lh38N0D66g3dfGydOfb0yNCbdXO2Y/UvfpqfJfhKMC3syjxz60AmHhJclHYXLhQ+
FN8Mf58oYxlrJB+Vwx7RzFbd25IWLopRpTDZXlQj0RCl28oRWbGMkXILeUx8fjnP
nzrWuAacx2NSbUWCyantQaV0yxM+FvuM56LAYKEh4O+Q8xyjNTNhiQO2/PtVboan
3rGBKRNEZ52Hjmgl/XIq9PmUswG8INXZlrfPpJzDCROIZIEXghzSLdfjn/zUvDPd
vdFguqe8jSaeyNl/ZuFlTEZlHGzlxNVRrdNfCRE8HnCg3Cgsf6j9VOZMxcbquJ6R
j3bd9L5MosqH7N0TfUGYQIXQ2nXKhLtP3tKf1RjGbcs48kqNVv0zAJgnmh7VET8u
luZaV0fBgnacYRjtd4A12ttttjbGX30EUuh31/UYeSR5UTM1+KdpJyodPVXNZL9Z
RocidLsgxZqNSIXuhlCDLmAhRHKZLMzctMDrDRGI0XIAKtxRTETRPlpYHz18kkqr
DbEw9N1+Bn8O5UeIZepIYnwpEGVOX1wNCm/GvqeMebmJKtP4J2kuODgdtvfjti3f
fou+eE3ttLmxqk/iqk0+i+WQIyWQX2Ik1QWGJZ1nhVps7tr4q038uAEXb7E6ZB34
MqBBjaPA1HxfOG2JXFxmau1jOmtywauW0Z6tgkznq1i2WFSxVrfmaXIuppdHzLUq
P80HetuAHs1b0onfAfY1o7WHSfY6jLPyhzfwGzWGFOpl03cJpFyqKSs3HI8qyxi6
i/Hkq70fHwfJvY2Sppi3zHl1eFNRn/y0PVCafsEFrx4+QCle90RD7kpgQr6jIsDg
hvLVjZjfN+u+94nl/44vgqeR3m/k9pzkCIV3ftlXpg0tfXm7nG5fkGDRMqpk2qM2
VE33RxlpujyiJOcvy0fSvu/KElUGCi3ri8j60tTYiUKxENRlXIsxQWTtmeTrc1nX
S+Aq5pcsqNmrQns231BgF5oHx5QKlc/Bt5k/ehOWyhJ2La3Cr6EX8aeXzYL+8PD/
jddmJivlDfBpG6Ii1ycJIGkIVSohDp+c+IulAwSCWiI0sI7pYI1e8dDFOHYxOo3/
eSoha1ms2mGzxjistkWBbUH+/T5K5h+1QAOh4fpLAscf0DDUZmNgmpAvFdafq+c7
T9+9YEkdAsd5snaG4ApqdOeQkFqj4aiWU0VkiiOZsAX06Mxm/SZNRcelpAdOunHJ
YDK55djDOdUpt+eaoHRcxfnEVQaEW6o6hXQNjfzrsVorKrho8UmJgvX9GUES+dFV
vz1by+5w2eYSyi0PE6QJLP9jeq6y+MEnkFoXbW6x8a1Vogsj59HC0ANdr5LfC3WJ
MAONzaM0S1eS5wdulzrfqesCM2coCOVftcnfezIq5zWbZQpoMhIZy7m7lRlFgY0r
p00niIlZa9dwy9vWcJBBS+7LrvmIix5JfKYh3qEwxgoMO5/wIaAClfm8sBOxinI7
nCy7/GuLJeVIVvGmxmSsOZyRuNPHM6nqG86HNVxxy3EjOE0/7uKKbSmdpq3bz9CR
a+NKajFpk2iAo/Tk1PdkOodTe/+nJck3dcekfOZKfSvTHHcHhWn+TUrzVx6x2uhS
Or5CpzwbI6e+vQm6r1s3Kh+G5wkMAWI6toZBu6bh1OpSEF6bPfaanbt7OE/ZIkmX
4fTT/7WNWm3+o0EtkfQSivFYTBNbr+ga4+hxEivWYOKCuWzFH5AbmV0OwFZr+yGd
uqX3UJA4QFlLuUi67AKfE5lyTzIa4HOHQ37n0CjO8DPkBpTUnYtpEc3C8/XiGC3C
zbA9wblE1+QuAexJJfiI/EK5KcvqUlFFJfNhcKAbew+HcpU1KpHwNZO14LmBs0c0
DJfArGDbKrrWuzI7DzHzuWGeFoarQK+0itB6yPtxp2AJFK/JOm0MAB67xSYEsI2/
6D+0ijpkPL87UIsDMq6msGDyrqRW4563uoFRA3o9ERX7jGOdsMqCFxw7urs/v+Ko
utNQipoypiq0vqDtm1Md5VM/gl97jgI8rrBeu+K0KWpwyBery/tn1nC5aHvy/07U
3haUZbOpQC8V9qxeId/weDt5TLoES2Fp+kvoNivgpyOhcoQoePyvJMPBdwiSNV6x
zhRFYTwQdrB97ZHIOPMvZJJXxbS/9VG852I+FAl7CZMn0hKph3zvKwFWl8R2J6UP
ma/zdQz4TccOkbe5xoqXpdZ1HI4JKhpZokpS7mqUBakdX8yQs3zp4HHdKBPo/X3f
oJHiHbKBeax2fNweuxJqwdulb7j7kPp3My/Nd65227hoA+iCYnyobI1jkAxXRiFJ
CTUFCs4uPhlQoVEHtNhbdbT8FHEgHf5LfETHNjSTRjm3WQIQzNjEwR96sSYxGK/+
cEaZcCUloN2OUPrNXLVzf9fsWkPfrOoJflMsLJ/bsIOSan8lpcOn4G8EoKxRF3hs
ZfczgS+7mlDgPWqaGAppo7wVQeh7TQuU/o2mCUuYhZTeC+kvXy85yMPdp4pDLoip
iPqAHkjTawxVKcNoMm+H7u2rCV3scf2RnxvVRloH23zepfKGUlYaWcZwqM8xC1Zu
W6dlj+qDnR0EwY6/oUJ5cMLKo+Y3b3W2++0suOwNeeyhqAzNOPBNlngr+0R9/ngq
oCAGw19rRHxwQUEPgJg/SJR8NmEy4nUQwD+qo69qmbotoAq7eUrbHDrVWqM1rIDY
SCvfJaPqR/M6K+tE1XdMTlFqZra9JmPJ9Sq06MMFSqXUKS2kHQdScCnCrtTO7cg+
ZUIdd7aKy/NGWkzYH1n8cOCa6tnBkuO1fSqgAeDyvJ8t1h5UUnVEj5LTmKYHxd3h
QoJAM4WaiBj0oldRRz92agcPbIlPMx6OdbIPs1ETB7JCxmrnjFBTPpizzE0d8LM6
JXl25aoIrExx1PYd3fWrOK3gdsAwKIBqUATHicXGzdJ+cpBQ9DphVqK8OAnkrki9
uRMFRgivf56YsqFEm4E4t4fDF1ArpFGxNGURqJee2EwDldrC9/HYc5B7aHEo08sm
J8qbihJrMUdScGIo44Kzrgt7ibB6/BWyFh+JYNsjB2QsSY9LOb9AgUY7cTlcyJ4J
GMbMBLYBTUW76h3iNkdgRDixc8nXZ8LJMJjdrINcnwPV/T3aAS/c35TUEs1gSCPy
xRdDIKwiXjWw5rX13c97RUTn2LWVRGE+iZx3yQ+GaFuJo6DPRh/IJLeZm73tCqac
ly8OUSdbWF8/2lOyHDw4zFTaCk82nlw97gk3PfXgyWWj6TVugmQ6sWUJ8V9le93R
vCawGEzcNCx7poyoERinZ2U3nrdneeWFmN4IRp0YkNSdhyW1EHmTCHDdU3cHRnFp
3TuM2Cnww/8+SrT5I9cEIZ8+bLMV0cGurxyI/h4nuX75IwbfBgnYlIMSbZXQno0w
iUz78gDgKdeXl1gU8E/kOoKNneOX1dZPfwEsm3BF04ae2D1H1rPYV+0l5C2wel03
apPxGOyGwkfEFhWCKhrWGrUcQwFBpMwkJ0+etHKrc46mGv0MXDEl9DKxAiSISrkK
hpGQfOPlwTTsGTNQSNRZrxpUQuuMKSgr7D1x365WNnXi6UOai7iqMiU//X/TdUZr
r5sFgvAcqf6n8NPtvzrln4y/2Xmi1T1QUTBDTzrvx/yzT4Dv9n8fZVku6ziB8ER6
oTvB5pyYK+Wna/xT1F+nFCvEpQ3Jg5K55qr3K/jHj6P4bzvyHqr5e0C4rc1GIu4P
TgNbfY8ULnpmub0boS5kDqjprYuCg7Uj5Bd3CZgBxPgbS6+M7bVVHg96IY+lD58L
DBloOjwWK0Ww5GfcnY+MZauRYIvBnYreNRR76W9aLwyDkO0NAAUglCYFGG7XGGEi
LBm40AFYQlbskZTahCOoXftUdKqzQhBpEIJvpLKYNXvOOa6DWzLO+YfH5qXhhlFW
AMa4FWzBm+hQZ4Ql9wPL4/NKEFXJTb9lgCgGON+pUlXd+7tULicf1YYwXEF6948Q
RSsv9HuMe38P+pPC2xicZH0XuBr7Q6hzXK2Fsc5YDl2anJCpb0MBhduZ+LoxbCl6
97dXRaGgdTeFAgwb5E+igTuwxA4BleeszmR+BsbzU3dgQaQMYkCuFY4mjZSG7HJf
cZcdJ2hwOvvpGA5fdtI/T+I67/MxE5ZctqmL7Yw7c1jgtzwPNzXA68GvdKbVgHxi
8z/vqZSJB8s/4GxWpaPxXJChHjlRb0cvKzM7xgpmw6gNtPNSAE1ZGzWAPSEJeVxp
vNRHHd4cLYmMsR/RCguJ+i41cuYr2jVRlcTvCabXEro0NzM3HQLpAU15cx9WVkLQ
cRek9OlNexTq9gPSt+x3iWMq0waTI8K0iMGUHh4dGmZjRkrmiUsaLwKtc3VbpL+J
BffnvalKQfPwusaFC789SxYeDVvo6zEZE0UrQKP1m4Y8MCr/Y7pdDiobtbwNJvXW
g9no69R8ZHxZuDTCuqwlJVbv8/9Y/hVr0D0SEUUpRsvtcM8KJZqn/hl5V6B6s018
P47TMpjNn7YmigGA2CmZNh6/raNaRjjBIs6w2z+pIpXUjSspAvWvbaqCE0NOMarL
iknEZ3fgat6HFJhnq0IbdO8tVM3Lse0LNzbs00pwXPlVkZazmjEoxDaFRmgBIE6r
doGKXVwG5cGmqgi7XaX+mphIYG/Ojzy2BsCx/Dse44xWf2O4AvriMFR4woAfnVjb
kn38dym8zFrPoML/3vqdLmQGnZfRdjaockdjnA2424xtnu4lO1MXITbJOzL5qEQZ
W5wD8AbCqBTki5uXwMGiijN9JAc04MW456Q3Z9O3WdMHWKyARhqOoolJS8+LOmDl
jDo9gS4JG3TKidpAyuha125F3slLNe1jpS9TmjCG8059el74+78olEwt5HfJLOA1
JqEgA4Zv9/MZoBFKlqpOZQpn/2yqAa//w1fZ7vnwM67ymZkHTXnBJTBuWy2EiQAX
62vkkJdXqHMOVa9RcoGVAPI1RazYOxUYUHK5vKJ1+dXbk12CwIzC2Mkn93ERImej
cPITcl2EzltWBiuTHSUezosLZMOsJ5yu872QaLcn/242zrPeubqUMAJPWkZ0T9K+
i+4dkp3RG1KfIaA6yXmKm2GqRROiFgWbvxaSYGQjMi0om0PonaxEy7Uj1bWtkgES
5d+b5L98bUPt13h1vZq3QETo77MilqLqnbYO1Aqax6p871n28rJjQHvV6Lcr4sGh
AGZKYwNsDC0ofGY4+yh/jqFE6BLB5U4DBZ5mohTNEgM9nBJTQufU0G9f4gpryZgV
gEPv6J6uoTiBiF4Pn4XNgzpy+WuystmikNE7cC6dHycSdqo+LblKIUm1aRKywImt
Gl6B3uRUZWR+2raEko1yFgztnT/igJZkuCWQEYzTgO3VgHKF+ra4lUdnh9vpZU0Q
Pixrt9gs5NHA+KrZGp7c/I+/Tm3CqCbdG68FwATwXXjlPwaxF/e3bffxpHd/ff7d
NoreLB75sZQGaK11CsbNC2EHKUGcrchDD9gual9Q9jzePla+tir4XsiyJVlk3aY8
cpF4MABak5mCuHI4JrXBEml/Mw7MsmQxXUcBlYW5D0LOpYEEDXRhizWPvTsx4MR3
L95GgEicJTO6O3f1Y6L2Woz2xxYN+UeXoTVenZrjo4RoTTENfuzzGMFMYlIg/eG+
bmoK8xpYmrig4CqO4mKSs+/RiWU2J3H4KIH9KvYjtzzCQJLpBT7jP31R+Cmz02fo
xpedJAKoCAtsoNgSOJBHlwiokSQnieGyASByCvLvipdC/oCoBRABDb0Wwyuf4tAs
xSWi61OPtNlI9wTK0GatLJHIXZ2U7HDgZ43UkRfwRhl5GKkLf7UXVomZYwFtyjmh
jB5gAKcZgZDCW4cYDFP6F0laH319ZGcJOzc72Gxe3MLFFcH8eL22jAouAYm/d0RL
PHmGm1TSpTTsZZ2i7PKNE6QqXlbygcbqbVhP/O+guaxjMGeb8cE5t5KEpGgLgWq9
eEhrbMyikwvCk6KwVqBEgo5k+MrJiUoyuMU1/6ha9QrYhdFK6dXosvf0C1A0wQDq
AJwaR1BrP1YbPdej6KAG2ynOSIEeRHsZO/wu9NEuUu5ZVxfNLnP17rMKamzkog9I
V5TWMbw6gPxzE2Jrk0IgvXP42Zfr9TucHCZoaOkdYUmYQcYLzck0w7f0V56+I9oB
mmSLe0sRkEwJ6ZKsru0f0lNcJZ/z1cuE6GbLPOVdBFMU2SdSjZv2lca6dPSkVn+9
ObeOKf5ob6IStmSw3bayWFWjiD9xihemqdUPKLj9D7LfSx6M4CUWMOJ/6WCD+ng8
4sjUyWA4qQw4v33IeYLZRmPTHmlQIrAyHkHZzZ72GGtb/UlYKAfVEyHSBPgi0ysE
sVGxr9qWTKkLrNOyj1JOabn05kwfDO3BaDplobJK1sxU1usBVKSozwUGD5r+2Q7L
nV+JHGfTgbyldqB1VGUVvD8Rb2XqOmxM1/QT83uR22Xm24iBkIH0wvDOlEPL/935
ieHwkagGGlwitixf6/HkFWoXSbhuTNuUXueBHJE1/WSWWrHHHv4/15NqvVZCznZ1
gbODHaSApwm/6w+uY6TdEbU0O4+Wyo0wM5eWlAiF6ofoUpEShAA/cn8AFazAz+6g
H3l+H8+hVrIkdWOkuxmG7cA9R75G8cm38X8huIlqHcu4NX0fJUesEo4K+atGmGAJ
DyQAomXikLgHs9Gx7ydEtBnFiaUGzoj66dQuVzUqeIbevj+Q/aGd2d/moHcL1MbY
/rsBuPa8+IOcpTE0+YwwI5rq2c0ENpVu4Z3rP5BF51cFWcjBheDw1jiajaAYDpNd
dnNY3h+so1TB+MVYjge/kJmCNL10JOehowpwLvHta5+zgU5z+swQxhOjevLcdYc6
8dvj6KUxkptb6K9KtB4CTtEkNkCxFMESz1HiTdL50ccxP9hLL4YTeOAixYK62cWt
lx3AqAfJQznejAXOJG6KgOcfGZCj2OlPd4yQ4Lsur86b4CsEpGxutFl8mHsTGmiH
S6incQ46yMHIaLhj2LYXgstJiic/BGgFAi9VUfqQiPmzokPDNRqr4XnoTDEiArJt
10z0anxZlXTYlhu5UvJF7HjuAA6kgf7IPMUG5P03BqxLQmA/8V/GjiGsy23rqNiR
7U1CFJb2BjoNikePVIgEvXdDfHoNGtBhQ3dbFKvIpYeatvTvYvzfe5gIl8hglFoh
QuIr5DYyFsah1ne2x8wqg0HAg8nrAZtDKMOQaYoV3QVwGmKAtPI6G3JArxUrHxZw
JogzwKMC8zFzAAGtQaf5G3FKrePwRHb2LiEl/RnGjI/s1+RwCwfpQcZhKll0kbsh
APiLfRzHAsU72MKMQ1QYd2wqzWYolre1lGSiNnCPRZNO5inQlq7xRXKuRUT0l1tG
ZAEfjKysQ6Osq9f8jcyhmZfL6dDhYUOVGPY2qncaPh9lLXzYI76tqThF8k4BRJig
eelnWKkbwWPxiDsFi/wBOiiriWFH6TQAJstGTXcHjqqzVZj4FEk2SYuJhoykttsN
emNAuFZ6gEPC/YRVbZex3OQ31aFch3+daZGjyC2VMVf32gzTB29KDrrmGABJ9InL
2s+75Aygat0eKOp3ps1LU7E5BLtkXduOU5rEsl0SBN5i+qhRZcbu7u6QeUygUEOb
MDFjHK1gUzVCezoHVNSWIaPzPBfZMP4x6kdmRxcAcQqSl5eaa4XNDjzvwIObun8J
tTFoajj9dN6QyISDtlyliF8TWBM03GQsvapmnSOafVtZGItxbm+t6uiC4nkDT/Zx
SxI0SoVPCwhsWsztjVgZCUrsG1mltFza+LSsykhOVAsCl31oAyRmIAjmUaTxOGsa
M0fuwoizCWEetZfy5tIaUBDmaAZD6QFTrm2e34NsGpSvJZM6n4Y+9g99kNVVz1ON
KN8BonQBV3j5Nz5+YKmh+4/8Qt2QozTM0otznEHqdEd+gIKlAM9OehObLrBsl1bC
76s21hlxAq9nk8JZRP7mgqL0fIj470lpDAtyTuOhe2nGhMqmf7BDX+/zmoKFeeU/
NtqO02EVhBEW36uJ5lth+k9gO/dch2zklLpvyo4P9gUK3o+ShmXzt27Q3eK7Rcdk
QhB4qAfp4wUZPvAsDU8AUOE/+9pksD4iwNwa6QbFOZ/lj3zcjlOsaOj9FfK/quC7
PcfEtAmkS7hhgSBkBvAuAV6XFDjpU+FvYexgwfz+82BQvBVUIerZXucql8UYQ0aQ
1xw2yBLYGWQlylKDGT2x6Ngs3liWG2YhbHfFZy8U/H45TsPYnAmGEtsC3qSPeUv3
NG+uSUuNcs21HtirT2mNlc8xMV7MinFDbUymf+1/9krQzt5/Wf7Mt5yUGWCfnvoB
3KFA8f3LsZp6FsyMEr/gvIQt2Zm41wjXlCNiyyZIIjHK4dyPShRu3BI6UVbq4iyJ
L8CllEoVi32Cm67uJORURWXRDsnCgZrNP9FbKHUc8H3ffBAo9xytF79NsM9UzS6r
/AnatoCxl8K6zLL7/41OlXXqVapPcqdfU1TJyScm7RQ8y4OflWLhdym+MCBKIlxt
3lRJIP0zRbTGQPZsyLLvC7tvZ5FKnfIaTgQHuaCYB5sflfr03r8fVuSOimwdaCa2
Xw5MsbbDk1Oa3gsspbmaaU1emBUGMmA8UG7i99cIuGWGz8/1rMKShVm4TvQqaBOp
y7EOyt3OG4YjBQ18clPAMYjN+Ce7oORjoGIESUc9HLacSQnJ4znxI/M3mRJRRCTl
f0LCIaxhNr3nr2g9NTmtH1+ZI7cSUWYJP5HPzLn0o3aJ/25dxFEmVWGiOFe1yxIZ
CdXilEwjAuqbPJhYtenW+N8dskdtgVgTBCet6rcImmbohHU3HfsiHDEoHHPAVA4R
gRkxBnd159q0lydQl7hkYIAZ2yKhcFcqPnRjXxZo3fID2NBZWWWQW4ezyEUYgOji
/8Cb7mCjy3amwUuw2PaZ9f0uOJK8nA8Mq8vdYeTbDBlCBHBue1vQZmkLTkn0QeRa
RqWymjHR+i+9fCgNRZy3zeL2auGfGGY0tXZ6H+AwktFcKA6DP1wkqj2acb6Mau+6
dtp+Kz20txyZDO2c7SjANW1Mt3cmMOVbClxrdE8Fk2aB7GSU124pS9MwPfTtXPU/
0zBXO2Svio5C24f1Y+i9XM9mf9nPiV4k8HWDYNDeuqh1eEdRuXO8yzsj6yljDzVL
u5SiKxgJtfP/P9dUHExaT3Ey7byh4jwW8F2iLI/fzaw+vlsexmsiDSprMwgsHKM1
p3vvJF7/vLHI81YvL8gV7WLVRHcMLJSr7cDsFgX0iMLxLcQ5luh9XVFs53ijUoFG
i6pqH6uzzBVv7W0Yx2TLQGY6FXIoT8wURpjy9Ag4dMDbcKvDJidpk8XK0g/pV65D
Fq1iSpyXTwK8ZJwFQk4CuLfuQxzXZo2qxfffM5aPCT4/qmoOj+uFLd4u8Kiyv9fn
+ycuSX/0zu2Bipo621YfiyGD8uRrbUYCZvmaJyqiKCQtEHYq6agabsiUf82NQCW9
eWWQzjAVCfyG7jF1xvEhJAfTpSKXBkKFXzSAe6PMrtLCksz0Ghakkgg+1f1Jm5tz
ertlgVlNiKHm8vBUgwmaV4wyV1L5A8qLaC2aW2fWnA1ZWbj8K6GXuLZ8EZo+YGND
6sj/ln8/lgA9wNUBnktXWCB2xlKrk3zi7WQwcPLkH6ijO2IyQ6Kl68qg1/aZrpXS
yans1eAdREwQydE/FmswByXy1ZJQofqfnVHjYsj4rCZqwnhMalikeiUHHk72/JPx
z/xiACik+8kkBZtRchQrdcwEoqLbBLD3RTzP68xZ4e8xft0LjlywW3lF0VKfiwBr
JjsQsFTGFxHZboePVQVkqgfcceK6YYsXfwDj/wspW8ftWOkem6Epb5P5CNSzrSge
DSF+RE3ErnvOqoGJ3rn992v0as8ein8GUEzHu/+1EUKEffOpwz8J5s3qx0PZ4Gxb
Ex6TIPgDJoBZ9ZxbtfhSlivXZiOQcwTlxv/jbENbPtA6lpzsspSmn5sikvT4DqF5
guZpz3yALIMFnnT1tPbiuMgZ8jiCvgtzd3tVXbtZrRE398lqVUdDEF9y1+y6sIGc
7E/dK0TW50/YHP98HMESO7/Z0ZCFap91ig3e4ATRw8F3zd9DNb/l72eBF8Ts+r4a
lIJeTEsEI+3Ww6+hua7hB/nnxo1re1YyTq08iruHclUirLht881Roh9hOICNmGPt
dlzoKQiyylvqdC56k1YPXzVLBrQPaM6OJrpizMLBCrXCyLTxFh7YgshNDZZUzWdB
l2jHM5t1/6VsW/7NWuQIKUN7kx0wSjWdiunFD0dfN5hjv+WwLV+KO3cxPHUzl5wZ
ICbugndalTp71SdOaKCuzxr3eoTEh+lEkYQoq7bozI8OWmBYK5HCfFA2reUd+5SH
v1OVTt//WEzapuJng/kEVjfB6lFyhIB19qxTsla9C+6vTaK/xG1EP3G5mwuqNd94
PD9lrWdInyYtEwhBMQApiHYov0V6R/PnqLkeehAgq4IFtR4eYlZC4VLMYHTXr+YW
JMvio4ahLJcFXB+AZCaGDicVNlKjZW59fmApL69VEUYgH+2TTo6ymEjFEJWVbkif
Vq6yWi6bwxWv2sCS6404L63R8WLu8aokp6dA7pcy1LH6QXhUPJCEMwthRml0k3HS
OdI00SiSREZrVPcMUu+cxaRT3hU6Fzw6Cot9ZVL6NCOl9JqpoDHG9uiB7fRr0y9+
C2c+vcIQio5l0UxIbnDy4irqraLuGWX8fuJCtq9dZ+CdN6RcYoPN50ovFO35tHOh
ToO7wr9PXInJ4C7JByccS/VLkovb7xCXFt+H6hswkUk53s+0cQ2XCQxDLy1mL9Xk
B4MBlFfmJnGzKf64jW26Jd0CtDcdVP4DheguDAdhsN+JVf/Z857rCYCCggp2j0nY
cLqoZGKP3yzOwBrN0+Vb+p7xgHP0WcLG345n6F+Aq/dPTxe3F5xIxnkVIdwrBFXn
AedGm7H269CIENdk4B+Ee+41zrchbT6G8h1y32KWMzmz7QuTlA2gUmz8QbZekco9
XTXYdMfdWhXPYYFuUUyy9iZK1iXKtJV1TjQ+2o5ZkFlQzU0y6FXsNfQmscwfjRMO
huXH1Je83Z+2I3vuTZu7kbLOIwEbuyF/wh1o9ML1hMp2EliE09MnLGAs74/iQNru
+QrRr3DJnutjFrHJ8Igu4pgwpIEgn2Cvihsbjii2551p9VXyQHF/nTaQCeajP3ty
/ex8WW+iIz7SNy6PGqDE0VzsrPNVlvRUb1a/6N7LrYCbW5KiO2DrWVlfWZ0FxfZS
u7SoyfWd0EUifKXttTcfoLgnPNqVnz6sis4AcZVnun7jFd+ynOYMLSAheUhmFfa8
MTOQl438gXH+REDpZDZviVlPfvqVe6LL/J3srLffuYBX0MG46UcEpzg5rJNoyotZ
KU6Jdr01XyozNf5cgbdWE3L16hRbO6e+G7fbsYlkGXuX7dNpCdAQvtc77/A/4O0i
uOmpO6I6+Rkj/ySyrbffhBJMISdKh4MdGt1wvdR2OPiwmZNCi3PhaTCDpKO8To6u
LcKpeWG77UnEcdZBAqMdXwAOty/qJ1HwKWpNuxvygyHwut4Q4lbs0jY0g++bMnaP
6dWlCGjOkdWnGg5w/1vyCMb91VH0YyOeJHRL05zmuD33Dh9CLaUbnD90eL0r7OnE
HEpl/t4xlFs8lar0U1GNOXh8Gc7gyZXCXzkFIPfyhGvHI7Fe0TLLo1vU+RrXD1gu
/zchveHQQpDfH4AfCMuWTw5J/QN/GO32hMxNWkY9gsjERV3V7c1IStGXQb2AaooP
15XR0xc+l03o1b7e/15QOyoMt85r6OY3a0fu4pNfksDKu0pSeOFCMl+ZnXhx173R
FwZ80P4QsaHF3L/5n3w4i/DIzoLYVpVREis/Gs40Vt1nU7uQ+re4HvY+dw3kfBFy
3tycdyWed3z94WmiN2/VbfSDi7rgUCCVG09BKJtxf678P1Cnoqqaz7dnFmcCpOsg
9mNusk7IojNsttmVdSIH6oT4LzIewoFJkn8D14ngMFbdNYLqMxiy+STiuzeGyvG1
FrEwwdRFnZNm55IN/2cjmPRrfIoWHGszr7f75DHoDwp6uiV5GKtATdmlgVXGu5pY
MIy2TJquZAiT6EaBc1r9g8BZZAzlMLSHRXxn4rlARvbtORPIUoWna5IPf1tjp/or
jUBNwVAJ3fnHZ66q5tFPdRDR3t3m/OaDk/+bE1FltaE7ykJkqHw6np1JuX71pizG
fsxIOrAg6yxZITRDmsFiRR2lnH5UYzNBoLk1cj/wrRRO8MBsvvnkJ0dFibYVlgww
uE+fZzPU6Qc6UP6gcEIPBg6ZtDXfgGuk5n3uDayvv88ySP9RXWFhAqqYgEae1M38
1lRPpm8ezOsjBxraan/kRqLvtC8oTYaWgQrtRRem0tWK8LFTfQmflOkXtkLwfyls
qnDx+YYj997LXa/EhqL5nQqxi86b0gkwhh4n/qFPiG3rdF9mFHf3OYTV5Pg2jQr9
H5FZ5WrfynhM5oS7fztcugr9WeDDofqlVBMD8/18huqFhg65viC2wp2Gt0m46ZeP
/GkDG2tmZA0lte0/FPnl0tqCoeJgi+eKinokfGUnSojL6WHG2MT5P1WIOC8NhB7Q
O0e8KvI7pYJiAYzXI31MsMcIzkUBaPwKXcOUEVwoipUe9/93jmhbCJRgiPR4o9lD
vMAVEMEm04qznLRUYBvXTvIJ8MVizmTtO0RxkLTftyueGp0gfP8EtCK6Wd1ZfMp6
Mf7o4xZUqT6jWJ8lt0M+DxayNA0M4aLbQn8CY/SI9RXZ4J2ZwBL3cRVclmXSa5So
L5fGsMNNafucdcSBYyPrm8tHvEi+Kbym8ik1Qx7xL2zNjsxPI13Ap2lLglcKUULI
MmJebe8WpdRWTiiOU3N4d8tXPZsg1fgZT3eJ54cd7VqwddJ4QGeu7ITMCx1U4o7B
xx9LjTqAN/yctojcNDIq1VKZJQ3epcQiycKRg2ZCL/n63IDy2OB+J3+puDk4yxVP
GWRETgRe4nKXJ2gmORsZZQzXBjGmqaOcwK7WpkVhwm1DyAJ08LWbDs+MFdepwZkS
YcPNurMdUwohoG/cQD4CyXpIO0lKF7XqXfPh2/yBqMJ0TtuxPiU2c4lT0ceihWUv
ZcJNhHx3X7u7ErBz/JCNj1OX05tSaur1UVHdHTJGrjlxPoqs4FJxOrx7qQ1SZjuU
VoYMs1+36oNPuJs2QNOqDVwc1y10p/gHtT6Gps1z6P2yII6/xYC9UJqvP6YRe8E7
ZfSeMfdGl+V4pwxKUfNhC1WDygUtSj/XtMxZD+CDA2ZxWIYE9BBnj8B81lWtxSp0
SiylOiihEmZGPqPppo15ohKS5AGs1xD7JXSVvjbU1bPa/x5JeKdEpGuH2a8SsMxC
BqGZFzHhzKDKMj0AGevnSsZry2WtYY36qN5at5oXdhHnwOkhGnUHWpianYS2Zskz
HMjUwA/xDAhc8erwAftbMTuL5jvI9eHlMTbdGFB+Gr5sm9mC5aII9JiueLdpbLZr
xi9cJ/8FXJ5xJMYtTRXS7ZU5aVIfzRLwBIQ3TdcHXKmqE951/LEwS5Op1clMkHQ9
z+fXH1VljbwY6zq/QfUM0yTjPuZsrr8377zpFPcWSbYLlUESppwyduDcGaFmK9ga
jilli1TO/vqJ7tPN0IeQYhR6XapELWZmTvvoO3tVN5PhJVEedxu6zOHmoCw8XGGn
VUpbD7zXNIoDm4IEs/RTEDVSqmN6OrPl6q9GrwIIbZJWI0fLtwFEapiJt7ta94FZ
0LGzx6ZmSpsJl+kW5tf8UVyIdd35iZjD8+dWnD0Fh78bEyRZ2rUdYRomWb8sPlDt
T50DJT8GIMqRmYqkIhtwQlPJ+Iv1DFjYS0O9mZxOcCj3qqeKtErxBHhV0nzrZQkV
i66imyR+y4vA7ieftUD5AmeYKpQkGc2CgmRE1xRkedpsY7ksjUcCMsvnbObQ8pb2
7+X8RI89JE9gzkkUMMulXCudDQHhfFc+ZQ4TaywPoN1r+4JskGFR01SR8dKu5z+t
Rb4TfH71XhzzdSfQnYVPoyQ6LDkB82f9gpOl6znHDSgt3ko21Zmi4e5A+Xo7FM/o
sPMt23+Xb3xinZqhCq5Rv2rgs4qVmv4qVyQrT+DEkC9/0yNqP3uxMT8KcF7wI0Zy
jKER8SE+4QMIYQTyFmYFOLJ7TwZ6Ys0RFzKgSKPwBE2cjB8GWhmshuGF7EB0Oufu
4YNHqbcf53hFkRLILE6FXSH5M6zOmaq22+swc4a5V7XaXDXdn7TeYE6fxBzxkitR
yvIlVtuEcJcx55Hta7MGsZa6r0Hqwi/EpQAI9etrnk5nO/8Q0njlGaSQ0Z2Vsml/
QxPpvBzlL+1K4fpC0DY9J84T9eA25583C/Q2/kHHGG2HOyH27HeGf/HFgLiS4/sJ
gCzWgmyeWFR8x4DeMWKUfaSgFixiwmn4El0EQ9BlP5husCMYFWliMhcwi79/tApK
ZqjYGB48i1BAH5vLsB4ufxC7JdRu6uvqI5Drld8BZsvkLesBmfMMGNIBwsFiNFEV
JpjRVYxt4XCARxBKFGQnxfwQGjumxJHsuM7mF0/zsK6TD9qwEhIMBFCwA1kprImt
Qk8qxFyf8Qk+mLPi4hbOgq8uSqdqnGFGSLtmI5MuEbmogpK3b4LMwxsJDZPEWVbJ
GUPNRjfDefTpSxJQb5ZEPjYiC6rfEi0NKJP25H01N4oSGo7ZTNoatUVO29aGeZrI
ZMEGnDU2NY47TNhwp/q1IF9Ch0HrYVjKBnQZBIPYzf4LU7w0dmdZ8ubhtgjdIypJ
DlXgN86tDYuRyKSQuBkzUmk4xlLmBm5MgT721UmfYp3Ca44mo8/ilh6vxyGndfLa
3xQ/QK5p+FdpzrS+drEezeDsU2hIyDgcUkJICSTvMxZDtOONQc+uiQHKkw+sUVhK
Qil9lXfGFe4niPeglG4pe3YZ1gF8syGubZSzR459uCON1yFwnvKC8Y37weA9vIF9
OEY2CNdyyntcuYScIotghrJuEZT1U5nptRUFqws8KzgIBjPz3yWhVB3LX36IbPoO
D4py8hTzoBK5z9BaJQAwd26y0tO4s5KNBGieMPJlLytNqaXkCg+H0hWvXebdtYl4
nni2H6zaScGKBBt4+UriBFo2a94m5kpW45poF1zdusQcm25c0qwMIjcZh2npt/pP
Yrk3M8JPFT5byufMWsRpbkZdnWUMWAXIc8BciXNgBnSjvVBsREzqPa71B7yBoWIt
ck2Y98SiSQSLGGoKWML4qBKK5j2Yd7eL1wD7+0zSNUVS2f/ZIZaF7G642GgDx3qI
wXHgv9BOdA9VK9aw6uwPnzsukQyq7wr9mLBnKDE6IawYsVPCjhabMT0rlJY46OAV
g342kq0Mwg2QYXv2yNwt81XV/UjXjxDJxsitQng6HxMZSCU4CBn/aWlN3VcM3m+C
X3K+DKlPk7VAlWSDEFXLaDSYdn9UzsM3PIxWXtQ5KPiY1xBk25bhs4zuvXzY76MU
GzqpI4+wwAFl4BBHseC/+EEzURTKVMx1Z50OVHvpbrQqY87rxeG4WvAHkIitzjDn
wtOuhFCNwR1zhmQ07KPnWdXJv5u1HzBvUt6wuwFCbCoiYt8cIb0dPjfruqJzUJIa
eGGBvUqHkCO+eSJxMw17MO2jewH8YCs9LXGbbedu4Jd646d9j3uj/LBz+MAKpapB
eErfhYnx7ilHK5tlcbe+Z1Qwpg1ngvzSmmWEOeqmCNd6hazWcZDT5DkGF78R9A/6
HlLkQNUljL4pBr0rTsSxoyKFyl+fcIeUfbXKaY4a2ex/8Fb7f6xfJwxZfUlpkuVV
lbYhUsoEQRbUmSIsOVDBv6h6penMQBgsphSe0pETnWWFpt8OhD55sgtBkIIRQu86
psIdG8vqy4BE2gKtldCd3jfnuYHl6TFq/tKskWEV9b+WiD2/n67j9b0xaMuc4B6t
y/BoaipDyZ7q5ht60JCNJi9m9TdxXw/xZ88E4vr0GPMGJDMcC4VVfZ0450AEkoFr
aPZara/NLikR8bpvp2knH92/HipONZBS/0RelKT5VAjkN7DndVXWxrhzYIlTmXoA
iaMJAnDK6VHgEbYhTlpaX4Acf9laiLyCqomT7TpICSkNLItcef9M1YtspPaBfycN
HB3F4zv73F3qERCb/89beIYZdaabxXQioYzgha7F2z0ZPBKv01z39a7Waxl6+7Up
qJCoVEbi/ptp9vML5H7w4x9ZY6lKIPrO4z1f/o3TNC48SFTkLuUo/q8FsJjfQZyd
aUIKIahSmggeThSpSZ4bO64+km7ofO74jfc4Sb/Grbmud34fXhRfZWPRWn6Odv5S
gxP/5ODf9YavVZDbhY9q5roqnw29s2uJbwy44ym4cAf+EGYz6SSPIJ7riI81MdQv
R7+KV5O4wRqDosmnkPGKKeR6qRzHJQxQ69WMWwPnWCmlIHFWDQxdyOkb8QXeJA8X
RJH5YdH5pX/34HSXUTO+o4GzsP/s5LRNkNM+GN/siW3pMF1J5UA1m4E7AZPlftY5
rE8KcPT3phvSCb5aXlM55hFciuphb63bheWzxrUEMusqFjq1EucNA5PBN7ZiYXIW
t5k3nEGXtyYWp5N44Js2B4L9PziFYci6Y3BfFwcLaEBfJe6Mq/cdD1dmOqQWCq1I
4qiCJguVSxxmsAusRRnogVK1qjZSpn1IJk+h2cSttkcSpD7jh9RlUTTBHi55E8CX
VU+9/x0k+WseYDbKsuEL0JuFWuhibPGrTIT9Lp9qshIR6Y+IHXPR61IEWREKX2KX
fWVEfsZ/5vZMn+FTdq/Hp0M3PnQkiAkmnmXwf9cEuIuJ/aVlCHBTyhgTD2t33+/p
bed0MmiWPoUiAUhCWG6KdEtLw5Fp/jPSiHrR/aGN6eVlGdnJmkSxUUbwPF8d6mXM
oZ2pVEm/Dyi5X+ksHONCSYm+YjOVj26Q4UV91PZuWMOLULYzzWX/GAbKN6hT4xib
v7/0QK39cfwBfSyVUzwLgftAagtQh8hBFz/IwY+bfXdbarIOJglQly+dhLlCM+wN
RGx0eaFQ9iZQjSZLyacETigHTAF/Yt7wb13aSXHwOaH+EYJ0BVmycHNg+X6izQk+
OJY5eNJGBvMNq8MylHTOUUyCohpF7H9ULqojEM3OvL3CasChFkgfenEK8JemQkNr
Mm5h1VJwJPMuuNt1L/vDbJUob4EScUa3Z99kHS6b5w4IfByGwf6uzBW2Pf/vmKrY
Fbn1kFSMfHECq2toZndjCkO3U6EQiolMIUkUG/NByplBTIm2HqqzI0poyMKxTYhA
4c6H70C89004+Fj/6AOq2SLxyDhFB8FTNJROj7BkBztWwr08x0VCtSMzvg/Txsst
tNNFkjwVYyzZJ7WNUxPVbv5w5GQ+yZcO62kpevRYFwyYGuZvnP+s5OCeAdlIhNVO
GHtnUnqNcHTzV8ssfTQs1/JQ8PEM2qW3npJgzAQZovQrus7dVXjUSukiCX2URbQh
FXqa+zi4nfxMIHm/l31/Xvud6Fevok5VER/CMCG5X9PKQbGxbO0nOq2M4/Ox94BW
3SmNpUrBJk5Mu019ozgegJem0Hu4dOQ9NFeC1pr8tetKzDVQxHzNgWk6HzROogI7
LJNHxYSpq4OFAjHFoWDbvzt4kMfZrZXtsL+ficRpoyPkEMmpykcUdUyy6C/NqDOL
nXwNKB0e75BaJ1pa0mKepTz2vV0r0ebwcna5GVIhk/W5VuTIZhiI8E5so+pXU93l
JJHZfShaLxAcwhoUUM69MVUxtnYdWYgxGyTKkuL1GryPeXeeWbK68IkpVIuhKoG4
bGoxVh7B5oottQRqW2zQ8txp9cu02b5+0KsFTO9mE8mZvpC0/Od4Sav/SdKndSEw
9zPq7dLgB9/EqLDvSZpCkLvQhIA/1hbiXiH+mH4TTkmvGSMcA7YOYEp4L39SGDna
9YkcBx48DJ/gV9BhgZgqD1JDMyUCCBv6ChowiDCgbOVazdZfciDXMzXAerBQaD/H
9RZltnRJ9KQRFgZykgX6bwYtqYajyCA7JosUVVFKwx3v5aa880VfvhzHXRIDhjGC
aNTS6zgMkHO5T02PFAW35U/k52LUMs0OJ9jXjpuyAVsEVqebXI9u2TYy5HAi1uz/
AceaO/q8Uqi5k3+hmtr2u1eypRlyyNdQ7oRzmWX9VGc8GffLY8atk74STP12+A/C
GzHbvGgPohMWJC/6YVrk2pilXA7QlfYeMDSO4m0H/fP0658ErrfxftSsdPgPxtJN
Cu7WdFhj2X6ixvhlqKzrY3jbDbRTWf4oNEaGKKk5repeN/YtzqM5ogigVpkd3WIE
UNquzP9E3KR2++mvc6tcQ3eZ4ek1Vf0SphxiZotIxFoLml2lPT5P0ofn7tCIW6ea
7lywTLswy50V6TRd1PJWwgyxqf0p+VKCBDAdeuz1AHT95ZvXqaQi5O/waKlAAETl
vMzJWcc8/vgUhLZrJQVID/r7l61FaR4lldSqO9QTQDctOq9x2Rd2UTJu48w8f5dS
85K0kxMcMvr4suecJJIJxW/nxHCarcQPLuJAz5jN+6dwuuOmgfRMQcQbD85qMheT
KnDELqr3BDn+cgMksFisR+zeTLizgfWJsgOXNAxTjBRcJg4+bwoofiuyqNNnwv+E
u38y0obo+LEKnpaHuiZzzMjxXVCz8GPZ5whdai3q1eWwPE2Fz3JT1Bxb/5JRdl84
sGG3lVU0jkkUK8cczi0k2Dq8/XkVE5PXzUOfdvUF8d/hy/TLXBqrmYGRErTHW/2V
Che6EDVRjsDg+88Y+8vgqm3zalsoHVbL3haXzIg0ZV77WnXOOdw3CJpwlrCGCRyL
ZSiXTpt67dJRjJ5KJ5f0FdumYvKSV7d/XiiKjcn8NGHdozfvxZHyv0OJ7FIdXUYT
B7iytiCnIbVVNdm7CsqHHdB0cPXLaxcq+yKHUw09WOc4Je3HbDxjXJZUeSNEB3w+
2//VMBKWVnq//JFn2Fitp6iSaBtHFbNe1T3Oqizp70aQ7hfAypUBNzizfjRriGQA
ZDXIPT6gd/am0SkS16w0GvXy3vGnDPwSUOHgxSAGsiCX/N7W785CvAT8l5Hs9NwS
F2F7XVU1nZUvpEjNWYY2LFB7v/CSdQEhavh8pF7LCf0u88m58NORiWYbVc71guvZ
AXVWtj1DL+dYVd3QNHkyDUWwvVHOV7ZF2Oi+odBHwCOTVkWRVJ1LLdDFLHKJaCBB
5b5QPOHBvxuxUiLY0uXIaBJ+6EFaZFZpb/JaLV1FdO7gjMroOg8DU278apiEo8cn
Oq9JDJi3pFt+vooYwAoPMjwKXNE2YRfMGUOnPFLoaKPd66MMOy6IDqc1ph9pRtoh
jFSrAVR3qM4o6okPIIZdidaAA4Sm/zHD/ZFBxZ+DZXanZqg39ZDOnFfD8G8Aam0x
KE3FjAAvlo2xOCqqpNgcXGWMndby+K+YYI3g8UTWLO2CNcyt7xxUYQINrl6p/2GX
KsMfsyFdnun24njbAv66x73+motdpzp6bHu2rymHwN7Kr4LvtOcXaaiJpUlbKwyn
eR/j48GYw+JFlc4pLW/Qxtrg2T2j4fTz697IVszpTbqIOtmdrY+ijbgomhG9+9bE
dsiKYI9E1/6JJeULajK3iAVWKa3D/O1rycnBowfpePjgbck7yot9Ea7UGro6eYPh
BhkLTSvVIyUR9q7qhTxcFgOTaqAGTg6eHEh1RSA0gRaSFutBg9xnpiXAZKCeuRXH
l2P1CmCI3bR5zabByHBnOpFOE3MTXVRAvDvmwf+GMrPWnBr55MXsPYfxmClGfCRX
q1WJXNYescSI0mWfrWOYP5CB0JT6ErZlELwGqTP0JP1UA10sF+15aa8/klqyF4cZ
HTktF4oRUnUDkWiNWfWm//njYYYyteN7FsHcqzI/JUV6L0qx4GfnDUgw/gOIYMo1
pLySZhTVrRNqs28S40DceB4YWR4Jezq9PnyQmI6licNph1B4g4131fqJbuDpFba/
aylGvzafopcyl9zcBWFJQ39iEZ5rujnxzjMtoGvGvK4SziepR1vHzqrU3BeZ0dv5
KZptdigfo5cr6AreFU9YVLV9nuH0hzUmsxKBc9FShhV0QZe+wz1zsk4PNQtvgfyz
0AHcICphBV05a4edKwjzewzCQAdGWzKPNvnJb+jZ7+m1VH6flzqeXuDeO8zRruIP
2a2Fd7qmKlys9wWCb21B/2oLYS+2LQlgOlxfGPUe9f+cweeZUzcvbbb3AfC80Nu/
llcLK2tD3Ob509YRJVPr80a3f385XmH4kdIbiFy9pCUf5c3i+/S79iBGgSw4X9sk
djiXoxHPMGrV3vrIAvGMuYI81wPd8bTYfNAUrY1Q+OAOPivzual8b9fSC91KoP7a
8jeUA6N4zhGRhZ6tOlz1u88OqNVcT2UXB8UWNk8qa+If4PlwwsL4BETCSwXJFHp0
54+B1Yc16U9O2UVo+KbHEXi+uQ42F1WTUCCsLHBD+Tos+Hbh2H/pM1U7EL0aR3bQ
+u6tGt2tbFqpE0+zJpD+oPpcy17swIKtc5p0cQgkG4+Emq/R3ETKRbWBESJWcRzX
1YJcuJKsxjMs5NQNWkR0VeQG1VM4vIdi6qO07FhIcHMzVwWi2nF22FlfNY+mheTX
AC1MiCvT2PMm+VmsCJ/tsBvNYSHU38heLgDrOYaUFeKpXMkTHEs/7p8ZkzZ0T+er
ejCzSvJmYEcuatAkdg98Dhq6HxQ9DIl1FYsozd46VWfriEU6y/rzI6+sHAzmoFdE
1WSSMe18gp7gBFUoabhr3emLHRmmswJoAWyk0N7Mmf3r9GUIkfCD//8AwJzjuOuZ
JfD2OMqS2Sav247Dk8e+rli5fDJNFiKv+W2tM3KIdrdhnX4GDTPrIvCvouob/cHg
0DXRjde/FR6hMScLbF60l/lGs52OqUhQ5UiP0H7bk0Z8jVrdi/RjUrtZfIhZk037
ia+hO4LR41766bVFndLp08galPsxVTJ2SbJg9KqNk8TF7kqvw7Bc4RcvBRYmUTgI
ksHVWbOZuHnHPgNVjHEN+O1/anBH1/qVyG6tdpoLDLWt9Ly8uSUV+rOlIL3nTxc+
HK2Wi1y1jt6hU+NRvKBOmFNlYqfzM2atmBvgNV/BFYVNzG8X2MVfdNP7YmiAHu2P
2op/3u/OsksCjkTEvV1UFtXbD/O2SrApZ3NQAj31gv7bjMF52tgU4ueMaavhMNvb
4dYs2nSrAL3XPnOH5rfPOzSyoBnKTvfEKHlntbDvDJjOt1ks8pxASrekK/gP6n2C
qCrdXYzPYFeAQDHMwa+ubnQXMlh/w0d48CCbfX+haPFrgfQTWVkmzMZ95cEIN1tG
qXh8C0Za2zYvUPBYpzPRRroO8/iM/6CApgS91Q0HHyTpEeDM9drVjueOqcagIW7s
s1Wd4TB99ERhexExRLVhpyg8i793Kf0t7T6MwR/rtQEJexDzjOgow909x9Ow5/+u
4ClmxXRk2JqGDNhBKtUU3EEkqIaYhDi6+36hkZa8tlQg+fXyGMKMDZ87JIWjB+Nx
khNbJnPDzJwJFDgRbg74cx8G8Aj33N84389rX/DVTCEw9kuqdmd3OZQCAKXFPHIa
QzQLAdaaVvBKvXFHg6vq/fHYEZHfOf3u107VUWmRE8zwQpmQttwYOKFu54JbJr94
CGsll8RArQi45R8a+yQKJ74uWrTVFzlzdOD1Glv8aOOcFlU5M3uiwjyIDGnxx9U0
D9QbqdUX17JAspn1ARV0WQcsWrQQ8M8OY9Jic7C4mII3oBuzjThC3J2DVMmM7grD
NbGFP75CQON6szDR1LW9O/UcBR+5E0tFt4svSUiFKQRYWPa31AsW8Yo24sPVKs1I
KvXF8+OjtHZyBdshDDy2MrS5Tualbk2EOPh4E2dUgch68wA1+rGmrc3Pv7vWNQ03
xw2j3ybCP27DHI2W+Cd06Bcqzl7Htimmo3JwW71QwwQgjsdyoj32FU4+pff+tpS5
Rr+zxuWWD/R2ABFKwppoNglYIgm9pTnugdTIfVH3qc9/Dallb9SPuqs4i1sGSltN
8F0X1qLuPb5wLbAOo4SabsbU6TO5c2PGLLYKNAdsZSgfDTVdNmRe68JEp59xU4fe
hf4/Ah20ZClLxto5kjAvwLvkyVLdrx7Em8k2XPcpgTmRo+37ZBqNYHbee/kWr3ll
JELuErE5D//1qrraeGooeuK5XEoMMdbIJBA2CrhaRo3hLyXPtsb2vaM3DZ0+rtQT
aEaRjuVH0DHkk4Ig299HK3V/A4FBuG454mJTXkJCCisL7qX4c89clBaI2QTJgoRy
LZChU79ScSfkqFNYyYb5HT9hZTibiErk0DLwuvKO/QLtHMdc25f2Y9Q+vbrG8HC0
wts8fcR2G9Fy42Qhqcaz+8YLLjBaGbaVEDUXqy8rg4XupxMg18EV8iAhIiJZUOyJ
fXMeVCIOc83YqqSptqcwXR99Yv5Kgy1CVPmP0w7bcF+/5+lFOJckgW7xkpWn2J3X
fkGlRGg4oWMSpr4bcbE8de+7PczfiiSAxog5Nqk5KELrukcIRFDxtbyyd86uSkgT
urKJK5wtosTA6+vpiHBKs64iCE1bUUY4RLnL2hSSd5oqWgs+cTx0SY206njCxcz/
kO24nJ2etwuZ7K18oafNIoD2L0OxPhEuLYDabc2uboa7AiAcgI3bknwZjOwcgAtf
QxxMBd4VSPJoogPSlxPda3MjXJ0iWlw2TMWqC85GsMTlNux/gEeNkmxA9QTPPlmy
muEnHq8iII+hco/HQCOUyDrfgU0DLVtaOiK4bIjoPgvL0VRO0/1faX87oqQp2ecY
oigyusI92DqEPm4G+MQF0fh4kyBcpNBJwz5hWb22EEpJarKUOtumUDItjv5HTZ4A
amrzVKZjMt1IYKy2lcoXpN7+3VhBzyK/aJUpn7QtS7n5GCPBig5rOlWggwseRjXm
ZppZCZwN3nBt4eczSBxKaX7fdopOaQ5B7zaJS4WIfELiKu5rh5hiURf5AurSVhSI
2vjViM1rsfeN4ntbvVJgGKcuCLFFn6UIrSuerLA6o73Wp3qvzvJEEFCgrKZXeBmc
k52F+kVDIFCzAWpOZIWsd9b6CVXRGhF7mN2+1EEZxZRmg18A9mXBX0SCJa3SDJUp
XzRepJYfrQszS+Iu6j4S4pcS5RCN+EfyTVldLKMWvlPbaZ30lYcMt+t8CXLBupYx
CPTmMZv+NiTckUlzMPR9seQ+xL9T+6njOlPi9+cgebrEE2G2OtmfvW7+ojM+0Kf6
00pXs3qYbjJAKj0g2GbSCXL9GdKrUk7HLyq0QCUXWKFa7pKSLzO1IS0dJ4YtK/w4
Xp7zK7E+5N4wQn30nu/4sQ5aMYOODrLndV3uEs/7XB9gpSMoEuoAAbgxT0Ukpf7r
UG98vPqKucidDkBecBJ9OGqob79V5cd5hnxKODroX+osH9m6hsSxZorKG4/vfIb7
UsBS1hhZrp7J5IGF0Gs38i7A1mXiIut+nWaPLndzhX361gtYJ2hWvOHxltCHPhh+
uzEg8oZONmU91rGiOakvV8c5ULWnUvEH2vcA+4z3BdJYWi4C9hqy6Woa2kWzSU9B
RsGrtFGGgN3FPoy7kr7IjFHt6ccWOXkNZ36g6/KsVJP30DJjSVBcO4NxHnLdbGKq
65vnUgA+Cvp9aIG7kPDFMXD7qp6/+gfW1haT/yf8SvNmhMXpjuSzUUHWfxC+UqHH
XVY9W4iPCP9Eg7T7FTGUlSbs2dJtTPpDBKa3A1x41QJPkJ8ZQJ1boyG1RaiUkHR3
cVImKBFImdRthOvkfvARGkbxI2RA2QJtbeisswBTrqJXrFt8iSSidIAPeKWkNfKG
hFYxZROTIRYBV16ETTmXoyyV5YSAZMh1vxpAOjRHZoAbYf9hkdzlbzB51eD6oLOg
g/Q/mb3SWGz+iMjid+iGy+Z4+IbJ2sC09QUNawD6MKubh+tKKgAF7zJNdPUBglew
BlVlokj8Fs28xtw+R57Kp+N41OgCACIssNHbVni5b8LRrR+rEz4FV+uYZrnjaECS
daE3aAlUoeLBFnn3V0/KG1Fqn6XbHNGPXwiphVu1eJuNZkgwAW5sRDrZoOVkB/p/
0H4cp428RNCsQLGk9UvfmPHaQidiyqKIZxE4RerMES7DAm3NxbnOZEp/RzHhRAnK
UihhHaySZuS36ogmatVGLmgXNsKI5Ut3wOwonh2a6D0F9MRTejY4AI4Ydqr7PyKH
UNBTAj1QzrX2xZhR8iHpOT3SiNqPKRlC1Jv9A4b+e7hvs3VWoxrifnuDQvwcomFO
6h8ghqJgBGMpRGDK8rPeG63m3QbKPQRA0/JC8Aau5lIlwXWjGhKO/KB5Z2HuggBT
JrGexeXxrHj7mEYfNfUVlic4nl9EiDYb8FzWjPntPTKAIZYsZoAZSOnfO/yLMT8r
vDDDYp6aERi/FI2iEEhP8g0R3Ea3NIDfScuJAJZXH0a+OWxcjw/K7lUza/r0lAhN
XvsCEmN0V9XDG/bXQYtOIPHqQ5z5Ay2DF+SDWA+c0iYh30iL1hSHzqapF460jSkd
oshBiz6h9JYGGh7Y7XJWSUbD3CzOFqB5RRPNcA7hxgHhQO4vSIHeGkRdDm1a2d4N
EivHfPLH5Cn1F2zgDGz9bjGAKEwu494MUeQo+bZT8OTJ5QTVZT05XafNX9s3EgOo
KiQvkm+bRmbaVSkkLU0eJgHnY4MOE5lRawqOuCHxHJVIUL7SL11+Y1TjzCOrQapr
281cq3DPsmJCYI65aLqiFUC/2RFE/vIOQ8Th/Cd2RIMVBrfP7zK0z8t+aOxzaZKP
Ks78iT3x0eepzTos0JLzvJS9Re+oQCjXL7RkLZd5eBEvlowrPx1YvLuFfqokBYb2
YH4Qhv8t4FtkQBz1781+KW730K2xpCpbSxD+IJpuQzWzoH02DR8Qv5wswPgz9Bhj
ZDqKMd5A5Th5iyJfNgusZ8blNOIhRt6/aJrSdSV2iXJxRyp5rQHYxdrIdFJ5euyh
aiZKV20+JoaiVvzv57CQjWllb7JZzhsQzQbYxh03EpAu6d0YVw6yLgr8WEC5EDzI
VaoMBkPe2QMA124bYiBmSBj7xdPZhLvEPTrRzcOMs1KKnaSf4pr18mLKdfig1v8G
U0cVcvY+FUwGd5ip/PetfYG56eEye9su+ltlTzM3O/G5hL4cCT1l+Eovo0cG2U3i
PBB1mIBy6B8LRB97+kXl6oP6bez6AiexkLhTkydotFctvnJKPsXJZvXDrUz0KHnX
ABVxrw/oIWmYYC/ZL61S0+ZctSj4FdadHr2FYNuy7FiCKL/smBg3hBNk2r1Fiwbe
ORIpED4JL/5NlsQRYccbrAMji7DAhJPRIGDEoDlMGOjk2my3cHMWmNNMxv8nS29X
UIQbwCAJvRIVhiLOMVK28pxtp9Hla7v+69YNZKIBG8Wuc2xcClNwknW/CD2t75WF
c6bgVuwihzM0CbN8sIC2GRr3rJcDlI7HHG1uLfaTMxGsBRlH0QUfbiUMHWRpzNo9
f3bta0o887xM5K79/FkuQcUljZejwMSzcMLjRHDXY/WlOe8Jc3vE1oi0LOWUE2VA
8cPh9y6jvlZZAIhNTSZt5uYBTSMDdhE4qwmeYKjNcCdPSADMtGLpgED3gprVkE5V
b0qxqvqNNyn6Zq1/JDna/ZV250FTNGPchbNOY2UNpRYMnxLyR9fbsVsOf0iUw6NS
cJs2JQ5WjJjT3Gp4l9qtqOQ6xqPPJcBT/waK0zr6e+n7VytCDvdpyBXm/sNp3r/E
A+4WE5jaVpIzB774LoOgAaHGbUTF+a6g2Q8qbit5IEC0HKkWj6vlwU9IlOv/UDoU
gkzyJZNIh1qh6fNBK4V77lbQSBtx8rinDrK6k2bHwDl0yBYnpPxGqp7XIQFZ/Wft
yKILUSaY1uxkwilWgQD8ySwaGczFKhundZJKyhRMVzkk73XZeGyEEdlExoeuCGGG
JsxM0sZtlmA7RkHaWHde8+pZ2owZiu3dfqdnEle1fDedPNRRol3DIHrRgOcT8APu
2BSa/hCv+y4FvPkpHzJGhmSKdrYfF65KCHb4W47e+SOuW8khABrxT44nX1tZyNxW
+pdZChcISdhMtLOCWb3t5Z6C2aDpM30d0B75JPRRgUW1K0QI6YsHunRo8c/DPTd6
Imcc+eWZVy7VL097oI+SqSEQ3yekMpqfapCXWYFyGVeWUrB1X0lH7lsaQhgAfyDX
2mlClXvYrh3TOfvyN1R3WlmHwykBdGOe48egJiinLrFUwKGTCxjsaS7pKQGmETEr
fZgkJpu4039Ln7U7f3R62uvk/EbGfK/mR80FK1yWwPXZuvlM+pnwn2UQGV0HWaOk
tQth1DxLwGmUMILcktelwxwFHJzBKaL78lBJovjLmmGETo0bVlcfCu79NKRvoFmQ
GgRSO2RFGRfLE3GrFX7y2HTpqGFQYFM0wr6n44xVlxc7w3W5h7KMIm/TW6yY/3x4
bFKAo/CSW7EFOXzGxgf7rpLQvH46c6+M2GNEFyjb8uzwP2skpfVbX2vnILsoEc3E
a8SpgY2xI84gPbzSQXndcoAGOjlOxlBY4R4UN2dV7c74Nj7e2/hJVv8EuvtOBkfX
7HZr6qmART2yTD3tR1j3rny35JtOlkyEqaRW5DPaQufRev3j/Oc/jVWT40LZsP1J
DLRz1CxJr3S7HARmjI9ZXGAv+ZVuIB3Uf4u90GBy5ercdvwsU2AX5F1jAl1qnVfU
cUVvqCYjRNXHi0H4Svv/8hg6CSMoJds7SoiwZAkHl3SxnrEknaXD7X6XY92pSrbw
olebtAE/B2s0ovAt8fStcoHAk3x36EAauy5y8OS5Wj8uOcMG3/ACxnkC2IZc1q6n
PZezbsF6FlCUhM3We00+lq2uinVD+TIkWADYolz5YVajVt7B049cf6TS9DvHRYxg
V66wk3ShdXIAH9TxkErHpkmm7f7wNR1lE01mA+V1vH+tHmjM+7aM7O5bhmbvdf8C
uOfx4iHeB8/Q/DHzCRXYrhMjcw8fZOKngUqWG7ykPp0LfeJ+AuZyiB/OuWCwpRLl
howmqnvro1+ZIZ84ohDTsKp/bdapHMrMkzA/IDWIf1jB4IWZftaFtUbI2qubBgAu
1CnwL/fpfBC0gmNoqO8rlOa7QPzdzBwky1dE7JeIcaPTGKcOR3cXKjE6mRANJE3b
fqX/D1fq6/p9WW4+nwfnnKyMSNtDMwZpE9DsB4ixIEN7u/EhJTvi6xlRhW+Y8ATJ
l1bJDfvvCtGWLnpVAhNqgkg3k7xY10MbrXWoeKWneEIn/Rp1K1w92UUCEfc+mWoP
zxgwPTq9huzafZY7sw6QV8gLps5wH8QuMRbExJK6OV3wCQFvJfRnELG1TANJd1o1
LM6dqVS8zqUQRtTFmJekvoj1ujMs0cGrZf1G4DuAqXDyIgRVxIfTnoDiiRaCMqis
OaGO5e5aSYAZi05mEdYNCyiwNzFmCoJOWoHtQW6uWTzAx5hoDsPbhoDWqofKniic
U9C3+3wf78MoFCDamaNok405EXUgjG0crEANoC9HnKY5RUKIphvAnEgb/bN2xE+f
5yQyUpxSlNG9mHuIxGeT32b7Q/8GBFBS2uTnNeVNJv7vTaRM0iN3+mBtoJ5VOsf0
1Av/ditKCgRM09GRZmOLP0yZV39QirrGkxRCvCzZNwUIGdXsIub65aHZ2aWVMjps
LZvQQqCkGdWXDG+DKd8EaDXj+eNbzqRGmeFfh3Q4L7zi6jnz4XIdBOCQSdtYm2Ov
et9q8gM5nPZQJUV7vfFf1nDQAUw01+RH257ti5zJc/5Vh441oQz1rQZ4BT43S5Nz
ok+cjr7T+84BSlSPi6+85wILEEeiQ8a+98FqY2JCXDSJPTvRtzmng27j0n0OBDKB
krLKjP9fdkbzqWC3iymprlC4nEEkCgzePbi1RNVfoGsVoMy0IYyG6VMiyjqPtNg2
gC8w7/6R8VsNDvt/BbPgC5nGJmQNtK9RLIwWJq/UsKN8GtYMS0XmwAFPSb9lK9wk
tIGBE8Ruy3TKoUdzyTG8eIEjLxBhOnsVl6YTCiuyzgZz7JVibaL2yoeQOesa6Gxh
+F7bMgbXxF3qKl4Ks5TQcqmR14y0xvtAdcc3J4pf3sclzFqTU5nO5wghG467zq10
pmh3HNXDQAaqid80ZJz/0LfNDyYalLwsKRP2FYo6no2bORDDbldeiJKQfrQq8zPM
++zkSlE00owyLqAxxe9LuaBukKciLaCCy4b6cYEaxGm3rVvM5ssonIfnEOn4iBxl
4r74nyBjFNysqnY1s035DYZRh6sDD61KAuIL1u5LNPOnKZ7RdgQnawYN+IJtU665
ux1kKy/dstM0ZTJrP98QdnwyZPp6zeQy5/0JmJHV9yTfmdwC+vHLNW+JYR+CL+yO
cpvZGt+rspHRk2MpdNyn+sDv3zHaV0RxBChx5PlhpZ3RY6DsBKAdT1bQwJQwj9mI
ssgAfk8hEBuWPa+xu/MSJ5eZxWxz7tLtSaa2Cmm526MbErW9WFfKBujGKaH0YRtj
+FbRLJdax74+dQ6MHjsrqiAcexpLqwoO4oHdHktjR06/U0pXYIlHHGO9L5AhO06z
etTXKwkknTT0/aFuvoVEUVd8I9Z50FCAY/y12Yig2XZnykcO87W9eCA3MbpSMF9Q
m0jH0OUU1r5kUaxAr2IHIuAXcsXtNTRPSRHZikvE5FUrzXuXYw5ECtCgjTtUAnjk
/m70lUME8EYHBIi77UaGUAiVXXuH4axUXmu7DFpjwkxjhhBjaLs39pdbBSwH6cm1
MZey4rCctk0UFUqMTNHaIfnGNLRqytzidGvFDh3t3dC4GR53gq7/YW6mI/I2/6zl
I9mMEA56DJVCyFQimi7de+UjdEVDgvHORluSZiXQSbk5C/WGqN73LIE5p4RQoYAc
TrnAdsAFV6Q7YfCrsUdGWN/7fJ0i75du/27w02y9cb2Lo8TrlYVJH4DKkavfbVEV
RiBEYoFTd6wcpNF8+0HBdC5J750r5GafQ/7t5WiLWu9DJdlskkQMEzxJoF2H4gJy
s3s5H8lecUW8unXJA/2wqn6+dDgELTQEU7OnaTGOKlrp0xaL5KjDYLs6x15bY2Ut
oUm3QnHrIBxY/XXSG8FcuJFpGgmfoTh7P3S+6cDCiGHeAqLo9A+1lCvul4SwwY8x
dl8KtCNTOIroOLtAag/ddJPW9e8MSLiWF4C0RsDTbVjKs8uwEgD5MvDYVPsIX8gD
RZu3Ar0OEMenJ1HdCpstpAUjzylSO/v8A3kqQQoEKcI2WRghV9BcMxqFCymWq/Vd
w3Aosn0nBzxJL1a4SippWRQrXpQ9CRKKIKd79tG2iBPWg7lfBgMM3TuB7R6G+b+G
zNa98nWkSmiO7K8Gqt5mfNisldfsXFqfpUL9dIuigTRYfwwac0WVk8CD/ctfTzTj
dtblES1R+EzrPNHjxf1KUEuz+6ZM76e4qk6yoDVAsXcCALgW/bUMK4Isybh6BqWn
Lnrs/ZnwMtLgBftGTfXKqoec8MQvB/EZJ8h55BcI1lCEMo2QBYEr43YIxDNvoP9u
wefZ2h3D9Mq0hVGZJjvpz40OBsjETjWIGoZ6mIOPzP+tj5R7wjsyPLXC0ZX+joEo
prjPYqNy3XbG0wL4VgXInKR7jVcmVzqtAS/VN7prZ8oMJ4ATllnVAn4DyiUoMrsg
F0AyemQOxOugQqIu4yR+eRTPYio82/wmFq6x+cxyzYUqwHD0CJgxebQyB/GhZ+4b
t4WtUi8UIqncZImXvPDEdLmfCDiSZfF9EaiE0p/M+w4rDK03LLbzzLVAU2zeNhW+
dplLNIpnQVveaNbnQ6mFPF8g4elXZyg0HO+kc7yLNxvur8HoNhMDsSrKyzuh+aG+
JvEbuYjDRph3nakmJW9N0yGqWp4C3ihLcoLgJPjKG2psAflontBSyckH7+wxkI3I
2SbkAyZ4KZK3kJ3C7TQd1Q7cZfbW912o98XFtBlGuhUo8rfgMQDdP8wIyJ2XXDF5
cme8e7Nq2+qkSVQAu4esOIhk54gOPU/jF2bOf2MBSi/OFemZSarTFuc3yRCOUujU
tnMGxwbfU/IY5621jnC9tHZ5JB3wsiAnJ5Ouf9Qdss/RpwbIRRey1HxprKr4LMlw
jeXPiZANzXd+nlJX0jjLZ2DpNOFAP+VvKJPYAzIO6zcvZP7bwe8YcdPIm+9WH+lv
30ybsRGRbjDagj+yZgkpAzs/JhT4kyPxEsuGf94zCBk1DJt4O7bif9Cb//UC1ZW/
Obl6J+e1GiYnE8yc4Xzgu/uo6+ox+ZDUCS2GBFO16blzoxLBaes49XngjQFgttPO
Xf3JEkBv3FiZyfr0KqCVZddNhn4QdykEBaXrK79fyvkLeqK55AeH8bEnjW016Dri
81pLrSUycbyYH45xjnIfadZUq33LmY/1ribwKoLOJLoWC0aT3IICzjK4Y84jpcLi
x/G0Ni5txA6Ot/FfC4PZdUSHUePuu+esE9G9TiPAI39AnDSLFnNtPiwP7eGvnRnM
gOCCqHvAOKHjiWTaCzG1hoE0eK70SleW4ZtkPBz9o3sg+3qaE/t2rIJnAyq99ZDo
I4PNlssRjxtiLsthLKZUNh3zO9ZuKrDZVECV9qEK01YOdemWF0oGKkYS+SghSugS
3DYVAuhEkDTeIfsoZHTXNffg1kHUY1DXcyL5QOSmNPSJs4oPM9CbuEaziKDSiGc+
`pragma protect end_protected
