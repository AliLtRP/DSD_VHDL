// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VP98N+OOVJkCayz/1vpRxF6Rg7MWlzRHpHMjCnBdkAjQAGgukdDGgABk6xr/qkgx
Rt4bWN0QXI4QYMpB3frKNtLlePxh8Q5fzXlybe67ThjQj3wFGnR2u6suV4EgMIiH
AzwEmScIUIp+5pnnH8nahip8sn7dFGwYi5sCWc8MmIQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26608)
DSCIC3c05ygV8pwPzgDvjnbFF3cwACmZ8iE6qcbJHbrJRrxLIU6fvHJRZw2z4ks3
3hdjREr4TYEpNAEjIyBQ4+1wC+Qxg6ZR4FRARSMS62tB3YPa7cIyGc4EEBx41Jwd
2lx1IbJJmEZfHYEtWNOPRcmot30+wd6+DuHQNHsNVqHg6EXdREIFjmNY/XKjeoCi
1UkWicb0C7UL+vx8Bm51o1w4HmstFhAo2FSjXQG5KUg/JUnnQYpLmlNKd+4lfjlO
j1Bw4iF/munEK0y1F+ceI1BEdl9eqjjUjUOejT3cn2voCHBHJlgVsv/zUcZEchCK
67Qnvbq5wUT3EjqAq6F+wHpUmTJRjGIx1fprVwhK/Q+DCW6GKdHKHnENOEvDJVlN
S2M3nySdnvBYvtUM+7mMElm0GXVyQZxhL55t8IL7mVLu2P2EtdJN8z2kRhrOllpO
p7TOz+DRilt5MdErWDrSe9Er+O2flVIuo+jg2HnMHCUIIoLRSNDphEUk3mPenW6y
Lfs6MBkLqpWwvF6cDGQkiu6Ojizb6J5gvIR/DrEoK9swez4AKQdQRiU/Qkd/Cncd
dGOUZ4K4BNC9pVahhX4qBs/wJryFSSoollm1lG3Qx4y/Wijle9lmI7wEJg+ooZdl
W5gCyLu9mvWKdX1W21LBzdqXcDUanEleYqCXTvaD/QO6BCYJyz2KEnI4L318oEuf
hnNfcUHw3SUKlN0lRFurlwlaa4gk5bjF1Fazz/XvlJFU6Sc8AHC7ozUxMxTMH7+d
Zz7h4e4WaSUlOH+mNgcIGdu+HZZmdGOQOePrJRv5VY0Zor2Hufivs/Lvb7WdJQFP
VnFptqPPIJxeBES9hEDFR2/f9C0v6xKPvZsdC61KvmeRYJI6mDWbxrJq0X/kMlgO
qUPTlzSuMUdEdokryPrWRGD5FgECnkO2qa9YDFaG2U6fCMNXqxjmJtJokXc7ZjIf
EIIejTd6v2mpuSqex7krZl5og4EVtizm5Hv6mMrutOBQzdLJYg9IjfOZJ495A1fQ
otskuTNwgLVLkOM+VBCzmbqX6RrqEmybDKoaDquHZjiDFlncYPM31qpLrTICC3CJ
rtZ72MtFZiK0alDrUfcDrIyXfaHCkrbET4yQEn+7B9RPkn5/ILRo2Br5sOm7HuSC
d2a85SkOuFbMmFzQlxLZFJAznj6rJFK6d1Lja0FZshCgqQw7prTVJmhelRxAPc+h
y9C2J9FQDSDWAz956fdAncmDC5VrI2ezQUk+u1PPK+DYCWEmFEsfxvwv4uqw/iqW
L5nDlN5NfJozWigJzS+k8iBgk7J0vpBZWaor6OLCiqwx+H5veGaMuckrf6AZi8pe
gWYrDAceCOJZsD5d97+vYq9p+NDg7A0lqgw8ihf/ZrnGf47eV0Z137oj3bzBWtiH
joAbG0Zkeq6gh4dwx0JAKnNUvZ668pst5o8yVONVLxCvoAWS76XYNT9HNhX6fojV
/jphwhusBEN0NWAahN47PQn1wvQLA6/537jQs0/YKw9+zTpCFCAgcIh8isk3J7DR
aakyiODRC9BsTxUQNQx0Uq+j3sve3hT41X8IviYXpee3zkEgtu2lW1oTOSME4N3O
nnzMxrZijDEKbOlxz67l05vsNaQlGxT99Bn4PHhNgjKrpa+nNwXy3+nMWfO50MlE
9tQa2Jyjp47p/PVTy1Ws1eg7fsKDI+wa1yabSFvDNXJtk9AoIDVorgK57+ImPNLs
nO2of3Zp+VjM4OG2wW3XbM4QESZHISB4TqKbPVuLWo90xdRw/bgxSdu7p4PhSHZc
C3kduxz3fOgabAa3LwsZWrJaGMrU/M1QwyW6qif6ep1f9BMLFc1xqXYEbAKKdq1j
K+0aJqGhT36c4JiqrqywUe7gHhHQ0n6NaKxp7sfI2IcZ1Jj1XefXdGgUF4PWtnrS
6tUk1Bv7bfPtUSvXd8b3JS9tta0LgBIQ/ulg3wNPW0LUG1Lnjzx5rx54Rh2fvEQ8
s59PxwH2XE5iRDQMRJCeCHFd95D7ze2/p8jp5ZClI2atrktCyeG2ifQHmb3R6hMU
GOXDUcxk1sSOGiaKW+50F8wlxM2dwhi9axatUPJmmn/1mK1SiExXmYw4Cj4pexpe
mNgeXpnZ+5zi+9p9qJQofLwd/Jz1aUg5vwqda7lHGNcla1hWsbptEpc9AXODfA0e
pgCIiuVcHSKRCO7HmDcumCp1fMUOO+519uMmFritzCuDjpem+9SZMD6sGG0vVSB7
i2/9/4Nz2BvqbecM1w+/22kfJFooKyOoPTLPWq9Mcd9D+6FwiYmBTc1siYs4aoKd
FjXYQeC596g/A3bjg8sEWnDAbLl1n0qzXpOSoyrtBHfGT6gEi9eS6B2/KUDe9E6T
x693jMBIUgjyq9x+UhrUIQCVXp55RPN6/mIbqrNp+/oLW24a3Dlds+x64bVZCf+r
gDoI8S1T9843ApD5GydpeKMoFFRGMTE8JicAivtxAcv/gcMjMfZXPYoJoZfxvnF6
keJdma8SuRqp8lxcx3EDLcC2aD7eKpKOo9MQJV16l7vhakzpxgSXyjfUTQY0/1B+
cZDGAgJ9+PCVtaHFDsLjUXc8nVIYqKS6X+bDrAUxavA3zCjDvb/mhh7EBF69hcP1
cVeoHIhgdZsvD0CSd5ulHyXP27ljEr9qhnlRA+qODFNE9VVkzwhaiTOL9qmNuoah
TYlM5r18XPhtrY5Ht0tTk1j18T+g81/2ukv+n8v8KsOku4oU6S/LX71rY6C27I4f
oRSpi8lVrrO/LuWWtFZ/KpErAqWmr1DuHHKmERigQzIVoksuMK4HYv3BitVXhZMi
5VhE7X879ivBUGL+nmPS7f1BP8Eib2MGQ5UTj8oayYmkehipp3Fj5p/E/cjel2Xz
Zp4TkBznNgLW0iDAqwC++ZUHlrk4oVlJw91pEjG8TOCLfgUdLNU5jlKzSSJanm3h
ewT98KsHXCLnEiqBokTXyuTlB/FRlocb7yrDdZDkTmFw4muzjSe730XnBsqsw03a
3E4B2P7lab+AIQ8j+upiNkwuJEwrogEFlJApnKKa511eOspZzs7jVeNHXe4J1JdT
UpAFkHa5GJN6xG05Z5Cms88EH9CQkQV8sMvlkomsk2+y4OqYGqrpXBXqbPPj4e/W
AwAVbZE8luZ83aduachubfWEwnTI+aeZxiuUrrT7IJ9ZnLIxbm4lWMfBzJwLqMOH
M5YSBnLNfMqtl9Xf/7Tamyarop8AJH9qeYaHp+xdNoBLt2O5j+W1aqDokLfr3qtI
Yjb2HuwmQSJFmm7e72zCnSAkvoMo6IWeW4BiFj+NxbzELsOCL0Ak6fmp68lwxxKO
LfYwi8dP023fML7IbblG1NEvHUuKC9ryjG0yrYjLsoy2V0EL0L/yxwdFjiSblidh
F23M6TUJtvBsq08lqlBAQ00dyZ/iuAwwvDafVN0lpoHRmxIXTegVa1bVQp4dq0Fu
T84ALCI6AZJ9ufoSliwkc6m5fYTOgoG0g05AZHuAeDU1DvW5hcf3T61/kjE+oN2o
cbOW8k7M6DyRIbem1Ml5ruK644IzwaO+/mImfZZqR04IUKkRBkZjfxGkfJLiPQk6
ae5occRun62cSGK6gf6tmRUi67iSZjO4PpKbI9ZfoTSrKjWQ0yZJjnGWfPdr8vaD
KGsHFS8v7CqD+dxsdMoSYW4uqg20+tHtA3HYH86cMHiAzDHWYlrMF3Id72NZrQOy
pVV6ZsvrFpGBzcIMU0AOiJ2CedajvQbAflTPFo/Eimh0aZcVRu3W3v+D86sjAApC
gfrJyUPYebk5bywrOCznc9ZBSH25ErDGw6GE3lhd/ZRWK3w/8K0UQS5kV1s3mZFk
3BHqPuOf2UB0BLz4nJEaB/W3nwkwUV9Tjuh03EHF+z9eoiayEfD0ymobC0XhdI2y
3DQf6SyS+8FqZ2EH/2w331UcpwAX0aGfM/qR6cdAucOA+H0TkWEQGlUGrL18vzVQ
bqRjYUI6aheVqHkm3AZRl7f61PwgidIt6QNrcW4fiAkEglhsfB85u3qARn0RT8Uc
POc/Vgem5QhB3mPPsOOn+GRnOchGLYT+V/l2HEEN4fsT5p3rq+byCkL0hvGowStN
qTzHUVS+vv6jLa+yzctivUds0Pt/5MjMoqle1KbdNHLhQJQmiB/jPfUIaJGNVW3/
unFH/nNM157h2BT5ElQAM5965//XZup2ltda4BXpJzii6pjRK06Da9xw+viM2ovM
3Jt0IPknSJNbNv+FXJ67Yd9A4euwPCaokDQRpP351zeyR+sWFFxkmjPiY9SQzYBc
9HVlo/fM5O2IgBiKhrUHKshmwB/qm1n1x0Q+f3EVcFZSW8nSJw9Hq+RqNe+MZi+t
XTzZ6bSg8TJSALUGRHtNjzZ08ZGwji4xkYrzHm0zFuMEuyWGpnHsxu5Prd5XaLV+
srgaeOHC6AAtzzNlNYXh73WvQG+xb1I6opHeeQ4vBDSZr0refiGkCLHfqecVJtrd
Ml7QsDrVVjUXtxteI68U9T2ehI5x6Fot/IRaA0kOyrsbQEUO5rnKZTZ2iDdGAm8A
pRfbY9Ub+G1jOAowjtdYutxGJiCfeIzYJ21BCu20o/4cIJWecyZ5VSmPrJK3V46Y
1j+/qI/eV5ZamPJV6vmFO3hKG1kY3zbdXSdRRthakUsMzr4lXtlbl6dLVDRKqTtC
ETputpt3r4unzq1ip5azqJoXdGZ/2e6dDpdoT2ZuyqGTN4/pEoYf7vNkhfuZ2uzx
AbCX9s25BbE/RUqz/DrvhS3y1cj9O20jhVtihefTF85gQMKSjpBV+KRTdbWVjcF8
ceu+DVXnjmU3e55EZ4k3qd/J/2wh/k8Kfr4uT5cTRRDFFuLoLJje9xz7KT7ETPem
/LpEtjRU39tvg2rhHfK+/ayU1gm/3zGr3CY9EO5Yyym945AZ3u6sW6KPPaXjn/zM
8/b1r8skD79SGWHRGaJqVHnyN4IQeMItaQpHVrcLeiHkI3fa78IbaMZ7RoghZpfp
bLz8XhjyMc+Uy9s5NOKedEsTNIrbBQz1hQVNO6z8aFP2Lm5xorWprEWCD/4N4nzg
O1lsefjJIrnlutmnzpet1cjTFE9Tydl4iJaBYBK2GY8TLo8/c/3BimytuXYAlYqZ
x4BQyxFlRDemAPSBxg+OET9WXQe3noyZDy1c3td4wDQbn5u8wvBA9uNpXum/PXMu
iAUu9aT4wTh26PGkzNrNOVl7tJ0o3Wi0cpEUWvotCvZxuV+6H5kRcbbUGvR2ZTal
0uRwEpAH69qcGiPbEWdgsVsMYZOJ6W1yQVPHNnleC1YTsZeYb6csaLW+YXz7IV9D
1SheO/5LqUoYneYBAEoqVIUg6c4DhJqxN3zoHZQQkWtkD4SpjrAoq9Rc8Pifjnw7
O2OIMNA+EMrUk/Mmg8VkcTuTDJQc/USJIiMRhtuFFU0c43jsWqZd7VfElQtXXce2
d0wPpF9Jp1DIr8VLlLtBf6o6pwwdDbXOfDGCjTq6rY/1u5GdDUZGwLIUEzDG7mWT
5xOAa3/ozEmCDUdKwchThT5G4KRKc60pOVO+pnF59uJl8JGs9QmFbXyaiGoWr110
c2tGnowyV2x59aDmNx7In3d1cRm2flzvDapt79ngylqmFXHxDs893TBXrymei8dD
TRJLOZ/EYnX5jx8iS3biYj2GejdoemiKhCl+yVe2Oe1uRKxOH1cYMrHvWlWbDp6g
usecRHfmfqjbRbq487GLEX+tpOn1Lwpd6U8WwMsfoAxYIPTg6Nlnaijd8Dx4+9FH
S/cpI+aVWqvMTSPUIpQdL5XWn6+v8srsXe0Znpdy9o0y11e+lbxtRpl/8hsOLnjo
ErJdGcGjoxV9NsJvJB2JpGlS+u78+i9vQZfHtajEMxKU6axf9EDlQiwr02W9C/yN
/gHhdAOCrxfcmA7Lf0e4kjFMkPxuY+ewrDoenSHs/uEkCFVrjqBo47PyOYcbWghX
FlvjQ9bvg8RU/8W1wSLA6rVqJaM7RWRfJHV/bu8lAEFZw0fXkappVJPoF+RonY8V
eTeH3L7i7VvbMUwjEUOh1IH/r3Qu9CdrLgwLsgqp7KbeNIqH5yOm2hAmvV0fT3eC
g8Hwr3vnvcrF0YjUs0Mb6mrRj8DE89yQT/0p7DCLlgYOEEaoiPAKnfPJfro4BcBD
XLYdBBaYN5IepfDGzoca7F8Uosui29nUeVSSfQecxFJAZCH+OnFysqgG0lzfFiDQ
JRjoHvaZa/1Ts7vNUuxW5dQeGSBTtN2/rA0e6vMgr/WeZ+e7/Ac/uTn+OVQ+cjun
COGkZ3KuH9VA4m4NJRprXTckodHB4IIVJcCY/gIFDuZ7su4M9EdFEgmAGyW4F6mZ
SSxGOGe//ZRwRNro91tX5b6KBcIl42MNW3ecOgIwm4T446PA7RS5dF1yyUMcKRrd
I76AQEk8BNERdrcDqDIa0BWV6cS2YjMICxVm8+3D7kkDIsUlkteMC0sPsUT84WiQ
PF4ALXw0L07qzCZ2XxN5r2rrXh3xkxmfFezUBhgZPPlJG1BP2zevXpYB0LbSXMWv
6dcn/dJ1j/489yC0bF16WGZu4r9w2WzqrDWBoBy94HW8Ma3DacKQ4p8Mwk1jvSm7
/HUPXyxG0c5xDP3pCa+/4V/i6F8IvlzW6m18+ZMqoIbedYHM18eBSOiANsrMT3+B
xaOOOW4EibSYX1702akMFE1c8dGC0YAHjD3yZ5dh6UKpfMGfXGnUd9Xu7VT1VjrZ
cjkVTk8qeMZ4cxOwYexMWIQ9PObKRFcbWiOXufrW/ddNounflW64dmHhKhwXkya4
nmo9RUa0g4JhE4fbQfHgVoNWTb/LO9zCjMX+8AOLDAOyWvTEXBMy2EAGsPL89XGt
xXCc2gwg8jr6faDM0jH0SGKt617wlYnx2HcUggGfDYA2bjkw0IL4AflHq79u8OuR
VT6kzek+63lF/k2ImrxT7RoyArxlsxTVSlBdOlkbjFocJsdirRrCeP1F04v57+9c
JaUCRrAvQtYt633ISJDzWShp8EMcSRnPnKhcJ3ABgkr2NohNLCbaRo6AUHX2uv3L
4D8jj3Ra2vq3QmCSh1gJ6VKo1OtTpvo7VlQwEq/dPcMMWVvOzD+F59NaY2ydPzEx
Jul9S/a8ZRyYDhKhcNWFrR+qs40hKgSu5FGWJ/9opxKaqk1kohKytmAcFJp83YPL
J0YZwPsH9RilXs8G9IkeXwJEs748SVXcMvTKLGVKqVg1Yffm5C/uiy865v0A0MAz
eJRJVS87SC+9ido3ptYNNLBDXOt8/RWHFTCtICAEOzcsx/+yIpsiU3E9GHFyNQ1v
8Yi5Or6SBFpisfszE3jtJ9CJGcABYZlx9yuyqzzYPd4vbu2IwLFANDpJsJoNwRP1
BmohZ1DsGyaqxHgfKeAzPD8Gm6zIrLlyRKrwMGs05efSHGd0rAngQP+UHn85lnwi
l8/qwK7ACqC2nWv12F3YQqtcV4/sCyLyvDTxYBqmtfWwk32XS6EcfXrnETYFecsb
aEc2NqWsOQMopwbFxyNDLVZikHkMqtiKpcEZyzpSqs1h5zl6B35TKrE+KVT7sA/R
ItyegzswuVZ0+o3sSPrVIGsOLejLEDiTeb3lX/hXCRjLi+3TjqJnP/yK1sgXHYux
WHcWJooO3W9c/NiOAbHoqje9PmUqnqvY7ygzkFUlzxFtDmfbHyRAXN74WKFC1fUt
kIw8uWNI7UAT04gAb1pEmMR8NQoYBe1mOyRGOhfc87ek/KIFNAsbcWuMA4NAVx4S
zCVjHY/OBV4xugRi0n8mcGv0yUWb/sBLuy0FcjTE/wyJMTKZmcuEGihHvbmh8uR1
F4i0Loj1T1zeQcpjWqlFv8JV5J/7/zWoo6o9zU4fsHV+H8O3WblF8NnlPeWNioU4
miTP/S9ln1sJPTKrcwdcd7LavKfnvGhkl7lhHvPL53Ofr2YmvCkE4KzeqamJkdG/
0BRtQxFPLAD+WG6H6ZGvsHs0zj4bw1ZNARS5roOFOrkJ1GJocadDVhRLKSm+gYph
3UWWm++Hl47Y003YzuxiitQbLF1l1nK91wXQCFXLsmHWbwcFG4+yghnmiQijIevl
HiH1CgKyZhBBIa+tkItj6ZGKSClGj10oKEhGm+bcEPA6sNAEjVJCMdWlx+ozFxV8
MF5/LTIlH73sjiUSMLh24rcqX7/nL0dRITqxaIa2uXNFvB5T8OIhEnF3tuhAApI2
aHYO4zGPeSdRGDFqtuqcnnwaJOCQjR6QqkTzuBdCtprpZMqCNIYNQBgX4j7D2bUY
9vHDckKZOdwmPPELyNxpcyvNHMp/co8wKArjgybIFaFUiGvdwgOmNhy9YCOElDU+
O7N7CqGppb1sZ4TA2olYdBB1cqE4q9QfcAU0xEhPEoTKbkyj+K8T0mitPuJSmzsv
sTahOCE0AtvSFijoxrC/jMb3ef2FuAWfAwaLeYOsWA4YfBpL9yZaveyT4nA31vNh
Q1z/qjTKW8gZk0Ewkw1fmlj7YELfnKGp5oZyfKxow+2PYHWHsnbDJFgtOa2OhYGo
II81su5SC9CkfMNjAlWfNB7MVhGpwfaJxIHQN2ggxdtIO1MwMKFK1/Jkt9jbcUMm
IzFTmy59q8LWIwZgsT73/CHGFHqk3SdWg6zNi7fe4L7OhShq3dlhdFbbJzrY5m8M
LrdPjxMNxtXxWGWLaiSDX7iieAnjjae3EsxlTIiBlRX6FCZQCSJIapgX9j+1h68Z
3uMITBCSxHkt+bfIcqQEGfg4s5mizUY/YGTSDKD0B0/QfivWYY3PuFhds76GVHVm
e3+dMqI5DMh1Gtt3dF2iPsCyaIz45gro+fcx59D6SLX/8DW8rO2EfPYx+QI42OWZ
0IlTxv7Nb9CNFIBYv/7Qt5W/HlWFfgHVoVE6JyvFlfZDFb43+cvrwP//XcanFf89
/EPInKEh3iJWkgvOj5653OMTcd7R3UhyibJVCX9AOOSsWjZpg6i/z1RlAahaxCN2
v2m5t/3Rk31ggpLAWskzm3Cz2Z+1PVEhRKUUauEQXvGXqLiQc8i1U1BLLyMTjO3s
YupKoFyB5iuAVQ0n6Ls5M8kHjX67oAl4aIx8ateMu2fqjWKUCK+eundHzpxpb887
HBbaWOv0EsOItHYYcRK8l0tRIlHIh/ZV6ZyniTxmp3vwO8qGLkPKKd0KS1+jP8Mj
kArJZzaVE8JMoxe4J3I6YLSgCgYUEIrGMMso8vUlF0Sn+q7Ew57vgQTZf5tgcBSv
QYaDvADsaV/HjfKRwLNhcihVlP+6qc0s4Lmf5IOWm1oOiobY+lHcFG0LeMNO+k5p
C7hwU/ts0kRagKi68BST5rzbmbKBW525JOqR7Y7ps2xrVrds2lIePAs9Lj2cKVaZ
QdIsV0dZVHl8ynYa+9xI7uibJYj6D64SygldL9AKimqr+ziquzxolH98cGJcfJft
+Y/hrrY4oOF72k1FHOZrgqB7memHkohuOicaSXp1m1sNQ5zGDaoMP/3p3O3JMnPf
b5Z6YsG6PuQ5SVTmdoDqMI81jhNs++5G7QXWeLybnG2thmL/sM147kfOYUExrPba
zI0w2CxJN3QoSxOBaa0OVBk+iiK42B5bR/8YpPShtwLi8hfuWFWSB9uLYgUJ2qx3
Tr7ejSuuu+vb0kFcrNf+ploXeOrGhVQhXR9t1rZT89ntjBDSAqktPgm/R3oPacq9
i1E69PgrQSgMnXqglXrgvr6TgD1a6Mwl1svr454ADx5kNoNvon+5BbTGoECmmRZQ
hVFUDD520O0UZ1yJcRDVgt1rt3kuLCSmuO+2m6feC+BPM7lXvQY5rWrQGps+xIHc
fgc+9EqdJijo3whrthU8INyvDwifLAD3EMv8QSao+qDUfxpriKacDmo4IEhzM7Up
PfTinumPGqgPPWUXhnttSNi9AatApkVFogbouYOOnLSyZV0Zd1J6NJjJ5qa4SnmW
22jcn+9JessPDQ+2mD0YHZACANCoxf79snHYE6703od6rcOXiqh8evQeOldfjhSs
CD1u+Yzt1iy2UMIpqu/9NzV9J3Oh0oCqZ1BuDW25hQHrtvwP/MwVF+pQC7gyuE3Z
3hduxEJZ8yHCi/2cwrahw9YdVp4FfnpZH9A9ysR3qJYYTixveaJzdhEHoHaYvQ37
V3jjLcURti27ScGRQkfsVFR+ckRXASoWntH5eOWGIwTw87Jkf9l7Sb41AA2EDPub
pAyJw5p7wvJv8G7Hc62IBR8IpsO2CuJi/4oLX4KceZ9WhJPSoh4texhjKeAXQAuH
fdPtDgsUxxJT2kNSQOtXMLotG6GFEX4Le3gfqpvMXG2ojddRVujnPbmVHQSiCrmy
KDOfjjb85rVmTSvnsqdDZpaP5x6PQS2K4317+JG/iQvgOOiElA6JX8DUMbxz6nuX
93eRCSpc+XxIKjtaX6IpBN7anlnhQX1+QZMfF3C3TCxtnOUm42OPJ+0Gt+LjCxJd
hQvMKyr2PgybYKTH43Dp+D5mM2g9rGkTwT1NEFIMJyrFFNzGnlhoqs8pRxzrOuCL
E/3jwTIcnuQSh/iA4bx72vSdBjBzNZf+K5Zkucl0T4Hw7eAHP1VEPZklqhq11iiG
ip0wo8Ot7tke3yFOKjjfNwgJEdjag9qEIAH8B49IAAMKPbFKaBcskfT3tS05RNwH
XTkPFSwME90fk/8MU0zeIm6WRq28vY4//fqxg7fVIFr9Gd1dVX1Mzdu344cN/jCI
6aOrq5Gb+rxQ0A3uKalKu8AGjmq+4iQ4tLV+i8MC/6d6aFlb3vKl5XFi9kzWGJmH
wrch5TurGo63WpSblG57pT0HFGyY/vSUrp7N2Dh5qzLMRzKeMmqymDVcCZMHu2UD
KxFhwoecwd5zdRse2P9qMwJRjw90vvnTfFQaYGTO3lA5J3bjcmQtACi/6oq7V6U+
0vVaPU32bZ962R98OjbCq8dPcaR/w6tRbQPCj4ERqpXKO9eN0+N8HGvM5P1P8rxo
RGxYGSc8wq8uImYN3AJaP1deYLeQOBfgNhx/HV9HOQ+oxVw9dqeIsdkasTBFiSpD
yqumzYoAGTFKQdrHSaOTNfoFql5qDLMILEQVmn6ML+BoXw3jGhs1VX1TouCE24yr
IrSoT3ef3j5klatqU3R8GVyoln96UCcEMUvUWAWCut3VM5s6x78skTW53tsxcs2E
OH+cDGkqoPwj29PlyGY3Ac3OGHihvlg8h/JXFO2cxLJ72GBKVb9XuBviTXEnzj4H
9krtZKjB7OBpdQbiKtedxUR1medZdbvoyjTvJd6q/TJr7lPMbIlKmYI8OydV9CgJ
Bw79WoFs/EHKmM91pKQldT1OrFqUd9xGKD9S/9FAtq59OXe3jhmgHcU/ro/87Wcj
54mc4Dcbn+3kMdhE1xrw3Ux34hW7PxilI0jHRcx2Bcn7odpe8S7S2JNhP7r5ZhHn
eLNd0uk/EQmd/Z3IbWfk9gP8kV4YikU+LhGcb91rfLGDyiX8OGI8YjP14Gb1K00q
PzHDcETz82TwjS36kIzKrPwByrMG9nkx5HZJfGU70A29882dxQXJzHBrQGjexBsi
3POMQ2kS9MUpPlA1PdGfy1Sl295akFpZNIzJBNU0j+Xu5oQvH2JsEkJVanC/25fQ
tog1pX3c6UT6ic5N2wAXwzJ7IV4V3vgpW8YXkM9wJlyZycstVxym3b1TDnIAgASL
zZFbfnuRmjYiygpXPuR/O2sjXQoHIvvGpw3/Sz0Ssn19cT4DNfe8IIt3UdGzr928
/OSxDZ87NYtrOw4ekxNgqCuRK0kKH56ckGjgWr0CVIX5WqYtR0JeJLQnCEjHzX8F
y9ZPye6ZsyNSq2YgueNso2BUqHEvu0sa0YP/GHKAZyXZ8cM7zLg8kZL9fS64IyDg
wQxY339vV4IhF5FPm4VTD1FIc2duKLcudyfqBGoxanghR3d5hmTsGURlVhQWfcTW
TWPdOA7U2qo9/ElWuBSiackinC+zRewyqsxEpT84HrnF0OC7YhH1Y7zjUPr8vDgt
j0uQwLVsVW4VMh+nMzP/wbwmH/tmG83SdxgHciZZK7AHkC2yrKTq2dYMQzE/piPe
8hnHnf6GcJo70BDq8PgrPqVmaDEQ6HUBj7iMnTj0M57qWb0vZLuKHIt1bJluJFNr
1HGnjqfUuu4jrnFhwlsxgtYSQe1rpak2OVI4tXOPwnlspaI19JL+AVnnzf/tlqJC
cwlamw3IpUxYpQxdpJVm+wyqepppNJSRoMh5ZVTDaDqJgLtk5UMh+pzNnwSyHk1p
0W8hqGi+N05UUVVpNi59lljLMQP8DlrxEtagC/+apCHxKZkGT2K8kwXb2Km0udUw
OHfZq2i002mR1N+imMzwaFvmxwzXSB2Cuq/T5X6aaLeawhBWGKpXcTBxrQ3HHAr0
qo2j7mVjImVdqj8BIgMEDNxvpubGbpN2uz59fqlFlp4PXUaZ2PEZVYRw9JJLaR5u
iGvpeX9t8EEhM/CUXv18lpUkKLmb0rTsvfRqLSSfobLN5Su/VNi6/TrEXN2705U9
sXIh8AsjVt6wDlYLf+yU9uie20GUDi0BRNcezfTEDCaDru4nuoJ7qlCr8lFA8zsr
yFTf+aKv7hO4l7TfmccUKD3gx+iLybKDGPYHSioZh9+uwwIx40D5jDx+q35xAwzF
0d0HaADOFpDSc0JzPi+sguwIS69/N+dlX5WsnaIyTZdAfKYhlyemk+ChyifLR7Rm
ecUjHe5OpMJDTES1dYIdfUA8tb72I8wNZNt4ZHjb9tL3WMyCV98G/H4nqoLeL5FH
T49QOqDrWhS8FACA0NoF2dE5mLc81R+NrT+m5ZEnAPC3vZOE6oeRDtByzH//26iO
YH84IMZ9wNI1WoXidDyCPLuayDkSwcfcGnD6puhxpHG330n5lBZgrJaNasiHXaAU
OvWvu3k6TgYUhkrOtc390mVqtJdlcYSMxy15alwQPqX9b2noYwD+d8ynfxEs8eau
UbQNpOZhrRJsZAvdA113B7osveRIaQshpfiwoAffSHo95Gz7Q6cznO2GoB/1G/nM
KqRDpPDMeNvO7iWQ1ZQGvVvHmP4wrp/9JB9kTmUGzM3RjNlu5DZpFOA9l9GKXmSo
hNkDIWMSwYIwnHUculQhFmkOoXL2bxCrL94N+2jdD1CcGjbVeR+sLwLvjJYhrxi8
LMltlUjjAGAZJ7pSoWNLz0Rfn2YH3vU6Mg7JFrtGd5Yv4sEBJYcVw44rSloFh2zJ
DSTI/ranLls1HuRLfuzr/yaRpDky4A7jLPR5NLkbhWkAYjNfOB7TdE8sPrQzjBV5
mDg+Xwr3PRDNQI2XL2byMlP3hASkkdB1dd3+3KBjVRPy59rUXpkINoZHbSLQSqNL
DGbTt6pKFFbi9aP1GxDk8d+O4bo9bzfVLiR1JXb9OEQazPui/bf0EPrkKSbm89Ew
JNuJxId3qucUgImuzvqryD2VkmG80CmPj/7HRfYA32U7BAtm4V3mkIqzfb0sEo2Z
EOe+0B5NQ9AkuUmuTys/mZ1CxNLZruk15orjynrsecmnDuLzEby0y1ZNvZXWYUdH
BQ9KCHgVMR2LxBEZySWE+CdaDSEeQRVLcni6TGyUCNVGSwUi3jNwv7ycz+etN4BQ
em4AZYi2pm0P6xOt2s+TjkKjadrEl7RtQeFfuzpQnpg9nZs5R2hu/BdVialDr3mx
84x0Wei0QA6LqSVuEPiLa6g19/qWigOBkzNNR3Qw+nym6Sbnt06tPymBUvR9vV9p
x1wXxLN0ry6mdC59Giuevfa8B0LRfJx04Gv+PCRRRjb+JSZG/lNV72+klut9IoxF
x1eaY4KkkbV+uwwZWLCsRiSc/XFdHPsZT+b8OHNiVA8Xk7LH2Z4GeizBZjU473kp
8pda9bTSowjshtdOD6y701sHdIz0PxfMKyScOzMgtCU+0uUKlcwF8MZLusVsWKGO
AEGhpNxqdth1w6bB8DAvimYMghDH6H7qKAxo23wmuUNGbBPN9Fs5dJttuF9asCze
2pvPaav+K4boQmJP2qGE2Q3wjeufckDGUFip50XaPih54V1bo+BBb58y0214FdJP
j58JmQCz/CHSdCMsz6Y0h1bfRc9EqdjEXriWPIpwST4y+9sgAkr/3qoK0NDvvDik
onpqqwWw9PaqpRtNWspL6l0z8tZV6Q90/hWdtgNMcZbkln5nXxXJwTN1S/crx/xp
lNLnGHR7pdykrDhI5RyjpRUJ9tJ29ufXmGokpD462mNYRPwjyQ4o1MN7OmdLXGq5
jKWWhMZy4My96wl2Nf7n4Ge0+1WRhNwtmCM7bO8Tybi0laEnl48JYVq2LrJPwP7z
arMHkXlZP+u2PCQh5LWyWqnA/iBJ+ffpQxtQ+gCh78yTqLtPpcyZaSnHqXxa7tjC
rbt3RvrYwgexwLqmdcdmT81ceEN5q0yfMYC4YVxrBqvmADGu/qEwttkWWIIvGeeM
7Af206y4QlcdQfGCchIV69R8eNTMtwiYxWhNue8TPUb/dHhOq/nr6xtggmg+clUr
Gb5thVpCywq9oHfCc07lC4kX65udnfwBlH6JgrdDbhR4ZxpKA6q3uI77qWN1Axjv
rSvo3w31SJ9tTO7kkGP22dPrxYgbav8aPOq4u4ucZHI/fmre62cdaif+s9vzVrhM
Ia955ZTfe8k7piNoX2zpMfcNxpGn/v7y24L5O0znixZlfwwzu/jKjoNlpyrrr9N7
6WkH6IREwxI0a3WS7ng8AL/bLUEA0j+HUy9Qjao5hR8rprGDti4PJ3MlQWOpAYAt
72Qs5923nwY5XVJ4X7MI3037TE2DUG6GsJ71Ufv4JqOvHZD1KDqs4JwoeRKFpSkK
5VNU2jbHxmU8Bi8Ewjo9mPoVG3TP61c6qd9oEULEFrwGYzO2+KJo9Iibq1891WUv
t3prUL7HY+Q2XEzcfEVtdHjGcgm6FkMiTe6B3YfNrNcCRe8XUZ/WY633v57BuuuB
xpVXUzkm6DbAObkVhTs1Uigj2XpnE+AyY+UJggKJXFdekc0frhAMaANJoZyvUos+
Y/ku3oH5qZRb0Ig9PCdmAV+a/h52GZBjic7sdgt4HsFXxQTzHJVMUFIQaj2UU/OI
WssVzyaLvYk0AOS/qPB/Wc/eyjnfX2Xf/24RjuhRMgcEpBz0fbWSpdyiahK2lFC3
MlcPxgAwhNDdSdxkbqcE4AqWlCJ11SN/wAlDK+JZlmDWWMnF/4teaIZf0aE8M5Lp
LTqcSUDwZKJPdwvyZcSCXodwLjHZZLZOYiNku0i/iYSAnliAU5zXVQ3CAdB/fN84
9MBXtoQ/jI/UKNnpHj+N949RTrm1IZhWccykphrAnmeJ8ZK9Vhsumn+ykcNjmieu
QfoiSyGP/ypP9XUoyXI+OJ1++V2U9bw2qC1iX2QqwyepP6xJpRLCRdBm4JZoqyrK
n1c3h53pSmwJAqDFx1/eGaYiW18iOC+H22AvzG8+oCmzH6cQ7hPMkXLfzxljLoDR
s4WJ4KN5F5eFbI986NVckvkfFfjcT30XenFYXjICHZjYg0syjTYqP8nPHHjsK0FO
JHmTuOyf651NURLoUZn1yCbRLBlCF2Z3staXhUz4vZpVXzfsIeDSVpIfkRyYVPm0
xisKvMiP0F/zIR5tqn8Yry8pytqqnYdNSRA4KhOYsbCNab4eOrUfiQOauFbGBFxC
qstLd0FxMeArRO5898w7s1kW8HogXb0BKEYYKXSEKenTs3jJb6gU436euxNxbkgJ
GQMM8SK7DkupDJk5izoQzX9dG2CL45ZhTDjQNckZqgf/NeZYQDQByyG74KiJlm17
Ly7EMHIA0dzYz3bLsH8+fdh2kObVfCLv8TPCgBNGV9WGf4wM/CFRwEILq69PTlyH
Eqk4z1NXdHcflmEBUKB5gilRjnJyAjPm54csuPOYWDoGjk9rx1Hci1sC00DmQH/S
jipPTw0VFoifGPmiz5acxV/3AJWQYZbRMqSLAC01AvssOstYnMTEogE6G31815Hm
nCD2RDSkHHQKXu3NFvwmf0ryHuN9a67eE2Fj2khSxtyxZB5eCAYqWB8Y+p2YfU0w
8OUom6L98HhJkwF/pGoMlbHCc2cQ4Fv3Jo29zpPUM0g7VXSG0Qv9lvfEtBEEz81x
96cRJ5DVwoyJ4iJdSh1O1aCv9VMIYa+NPAALBwSkfqydHdkQrifkyauYEaIkkdfS
FtiKYodqnikRaBPqAv5uGd8I3M02iIavfq0EKtCvkcssYCSeqhw94/I5NnUDdzIY
x4nrzdQCI62k4rW73kEkoY0QFWRtn+3HSqTRUsO8gnQDthAt4yfh7nMPG8T+lDZa
GD6zp9x0BFUxPmzYGTmAnREfIsdQ8wvUO86dJQjmpmdagQ9sZ0jpkovXtAhsnKPd
siUP0pz0f+YpcEON04UmY+0cSftImWn4neoh7ln3UoCLmRQkJ5yVWJTmtVfPk7F0
S2XqwWNs3QrmBlvPOVgzA9eTztbFULhsaZy1rO14r/JwRtB2NW7FZ/bsREGKxq9N
Vcmh6nXDCeaNFRGQJXdcTamqVjVbToZrEUCsoZ0eWVh1xWp/NDaFcnh8b0wL1b1g
D8Qu+jzR2WdZa8CzhovsuQ9kyOFGGj5CziY1N/eEd02p86/dL6P3Ag7NcGAIu2KD
5fZ5L3s+MV/SIw11jvKLhz58novJV5ueMGfWzSYGupKa61DylV/i32yUlD2XZx68
AM100T6T0ugfc3Bl3xgW5qltYuHOk7NTc4FNBQ2kMpViKN5S++iufvrc32sxG22V
DADFziNJ1B4ZG6+kdBRGXdlCp0DAKLcSm3WeO/W5LZgckqZmUaGtBnK8W7ySJA9I
FUIEgZb2CtUAY9+2oIuRwS3ihn0KKJs3RScMMAKiH0/clVb1SmmX5lHyg2D8CxTi
GJjPOuVjcV/SN2EgC5udfa5aZnh9jsDvXLa5/IxYPQp5nefwb77wjoTwCMiQyloF
7/Sgvw1bZVkwlN7DEZZ+JQWtRgfMqPRsLnRZxC6UJppctCbynbEkdoL9JxU0eaT7
zjzzwlLcI6gujPiOk5iHpjWEFIh8psRE8cjzI67lgYTItp6wvnlOwHEP/B5Rmnam
x4DaA2JNXIQWfFB2E3K7mT0M9v3rzXYwSg8rAIbzOQX1paC7fYRgEePnSIZrT4Pk
HD4QTJqwM6gxHW7CC+4e1FgJQtRnrQFUEaaCkHX20ejU58aMfGw/fFESVFjPs9oA
d/U/LX2DD4uQDEFQBq2WjsSubpSIYM4ww1NOs+T62m/gzCy4UqZUsTESPYgJ3ZRy
ScgI1LdTOTeESAvb9q/gE6OGRLT/8S5wEU+NimoKrcAOq9rvaoC9ApFurI0+qK3I
9d6dR14bgSS8c0kTHCm7sjWP4x4ZSrEzTE5o9Oj+JdBHkbDOoy4rmynK4ZBS2QMi
B9cNmfwvXakGe9qx3yvf6mUHCED5eHep0ucDMz9pBKKKY0NXMYLYiAZGduzsE1zO
QOYHwnR9Gno1ZE2Faqnv2s6NNDvMPQbWy73CVfFBcZJPWKjuAgrZSrXyWw1hVHVX
0yZa2ah17u8rMdsblpjWk71xb7gyZEDTB/3mfwQcoPyDYrqUiY4HBLt3enM/zF+r
17MZJGOUGuNH1gOWXwp7GSW4Pgs0W/o1psHpxaJhJKX1lPkaCNksWS11Smg638op
sU30bkFmVdv9OeYsyvQrxYbrtBikyHyns1aH1TAj/2k7T9ZDNoUVyVVWVj9pcinW
kVP1cGTjJZN0w0BBYQqrg3tBf8Z/CmPNjKDYB36M6blTGqeSOWhzeqwIBtAINz9r
s4YLCccamDwTnDdwW05jtMzRo+6pGt0BiEvSDQZPwWwhWlM0gCH5hflaRL6xP8aL
cKdwk9bh9oaGU/pMZwjuA7JCL8upadwaOu4evBn2pEY892VXhNxz054+fcz7M8AW
AYWSVmmbxOm5UbhvAUWfVENb3cV3JX7AphObsjTYmR7VQZjkB97Nr9WcXvdEcdr8
Qghy+Q/jd5//hKfdWormqfdWCLOnpgv8Tl7CCIievKFA+ODIbfl4sqFPVN7OzUra
TAduHnhLOFIVgrc6rH/T7elgaewQMWN1lffnYCGN+ECMzEb+HnjWROttKIVVVN2G
IySUODsPyEif/lY9XFAC/o23UArzeeKKBzcxr7KlXi4LzFqtq2bMBItqybtCYIeL
BUUn+Li5xCgsJ592hOh06vNXW8u80wF0KTSNzKIl+/Bl5kkbb4Ry0IH3RI0GhlLL
qh0IH05z28iusfPhce8Nq5qq71YfVDH0fhpt+aY5pONT8p5W5zkKzQgWlKsN4jGI
3cbRFLazk0lQhqJj2HBe/ThqAacuRSU+eHqEgOS9Ned4RALh+hiWOulbck85BXHH
iWw1MlOmIwfBZ3O5HQ2k2olN/Tjxq7FfqtwTRxhKdA0YOscvj1GN2JibmWRwnbEf
HR+NL879o0d9kzTrGc9xVj8R2meluYz3IX/M16dlE6Qa53f4G9OAZJodQCgYMzdp
pDuUw8MBr1G9wrrHgZ+Fs60Cm2dD8tngvmep/+S8lXmrkFMV0fuo55C6vY7nXpcb
KfiNtafvSJjZD2nSOefdmQdabRdcy+Fyq9kdM5dS5WSSIs4B4XZ8575hebv/VwsR
5dLyIympzqWrfGkMJQYw66Y5AF4/l42pY1KvUuAxOvVzw9Qp5Zj9jQ2mDBYcNKOB
f0gMwsrGXUgoxiA1TBwcuVCXJqMccaTHx/ebllaeKZgVxcaNAgvKfUTWvtGfXAcL
MbiDcFBCU9/eoPTR5X/Fgsd8o40AoxXYoyQluaq29XF3G+ivRRLm2PPAZlKmuiXO
9BlM/HF7/8bbUn4c7T0mLyvuzzsRW6GOkSIf/XiLwGZTTdrcP+JQ2uocRqbPVsJA
92Ed+M1jReEKnP9xiHKuv3Lns6lZLn2CcReMdKzD8vYFux5yosBSylRCZBevJMnB
REa/lPNDS+3Uxs6cLfvEj5emVMdyQNwQxw/ZQuyJYCvaUguQCBDe736eiM39RsXm
WsF90W8yeuxFwm6yOJPFEup/zSt5lxEhlnwjuOOZ/t0JQ5fZvln1b0jx9NaoTzVT
Nugsi/AGXm3b0WNT8Um/EQqCZaZgIN3tLs6+Q+49UbEM2hqJlqSZCL4IcATCFE3f
X5IoeX2GpziE78Xc+okMc7J7vXlU2ITJ4HLEGLOPd87GcCkQxiE64Tf5K/eXUxxb
mXFGhvA1K7VkOyJR5cVpoRHynm0GdWew2D+MmQmaTXsRnVtvWc1+R5mBr5hQ6jsh
HivIr4OHAjjXgLxRXHKai3+ft2WNat3TK6HC6GLSFucKsu+dee9rEqC5jDLdRheD
Fxjo22zrXfevFRj4I1INhnPDi6HdK0hlkkO4IB0UkTOEcgmoCWJE3n6cZmPlpXPe
oQqfHufBnD7hgaiH0ITRysfR6WKYGZNmlfoRLM6KY+SvhMQmihbEb+B0PdYqSL/V
Gba4yRTNpDnz5hUovYHSd+z/hdxSeH6CkIQwUAx3hzQutSw+IUlbaXiuZq0x2kMq
9b9uztPHspnNWHvmaj7qBf+IW+bht7Kb0ClrlR0DNQUP525Y0GJWZYOi9VaZ50RV
l4DTaVGlK3uiTcwRaitL7GIYx+6uiDgBkfHB+NfW2/AjbrGpqjNs/W71zJWyjBAb
Z3spiDp3CwXgTE/E6keKOcxzNFb31f4eFbcNp4lm+ikTEldPCSJR/ToovWf2U/wM
DQajeyfBRjovbThkc61BypWGQ0XROXGRR9vEwGBkO1v87dvtCXCxTKd5kEO5g97T
xNkyo+E+AZf/PwhJTaiaFLC3GAeUXc5pY6mMAeP8rsD45XPuJw8NZGYsb/6+yGhY
TWGgEktW6DcS6hojsJXdwrIT7wt3xvonQ/ADSJyyXi7W6LKqK/5b0zO3w8jMwB9I
JT3mAyM1X0+HYVC3/J/mpl2ESY/i7zqnyzUa7Zhft59pFVJteQZDdK4cFZ8WxZpi
5JEEYyiyqr1O7MjLx4YG1xXsSgFGFITZ4Z7a+uJSRI1f7C0riNlPu2XTfEuerNRK
xi60Sk1dd3X33+Sm7zx3MDhOvdES+KW8Fn3BfbQlFS/Th3ijNH7SSSdZtN295mDI
PhZ+9P+JsZ4WcgBu8Vw5GaU1nVlFImlWSlvURM/ztV4CDAM95WscG9sa1Ik+t1m7
vv4pECBaqEmdm9V7iEUVQK3m8+6yi50OFxVNTT804mFaH1kwREZ2hSVJW8Pg0hBi
G+RVMGKSTNF3lJidlV1d6q4eZ9vs2ssGGs7fWvFduPIYqvUnlEwBuqWV9NlOyih0
Uh8qSueWJqH6h04l25bmPpjz9Jg/EJMsXe39gFe6n/iRuMfKro1TGxKmHAu7K1wo
IoAYGhAgKjlRX0f/01GyyBf2peKDj/2HwyWUYr1mW77prD7zPnfBFojkUcwIFnu2
dzr3YIX4jahgn6eGEgIn4SM/rbtBMxK5UvCNOWCfN3Q/Ru7MaVKYmbhI2x8uz3uo
vCzmfR1VR4IrKu05nqUvWEf5Rdod78uVzgCvhL/yKEeyaG5PRH4xEMV1rDXX/mFR
IPeceLQkXRPYwxQXOCf1Moj/K4qrW/qcQ+Bis8X+Ttt4hwOD31T/V9A1EUY9cjNM
gduJFZad6M+OPSkTb54CRGBFPwMUgoSPcn9VCJQYWK8A9DMmkLOn8gGaEDqEL2sF
QjbxPiADRUu/YaDDHnXlEDBmXE2uVYOsng4AtjdtgZI9tDflMWjejcfvftF9b8Tx
mOq3hMvFr8MbyNp7HbFk3MxvOpLoA5DtCuL1NCASF2sjELP7TqDMWrV0gmRwhndZ
g6ePXJjK9Mtd+3jouMu+pzfhn413sH/xtj6dsLTRyhWyQhCFPJDXXzoKAqyBMLb8
izjPH5d6oaBlYdt7B09AuFxc2j1v3cnZWHCfOPwr5NF/H7AtIIQNSYXKM3qz92RR
K1lso2KIDF9pRbzY8/P8vB2i6lFiXPFXf2FJIRdwwNgdO9L3VZVojUo+0wbf+ecB
OUwMDhP+eM9NqNL7faAmrGGyc8iGpCSHGDDxibbRXZ/rzyQNdYvQ4uTWeEdXVUpN
2uXrN8BqAK/qmSg7CtE0ecfdzEtOfE5DnWttgsqC3JlhauCymUqAY+VW4xXBorV9
NliWnVRxO9cJ5hPqsDMvc4RpOrlvaYZ7GPgl7y/6+JcBAG8B4Da2R1KRAcgZrJMI
TsyF/YhJPViDvJBCo3TH5ke/OqwQuubfPPKutllb3h3AZ8jd9FspDnHTLI93/HmK
9KjwN375KM/D8J3uGfskwEd/lJ1QiYDbXQsijxyrUSly7QX+DLJ9VAHANeh+VhO7
iHt6kOLCtZVw+KB0TJ9hu7vgQkC9iSDA0+/H3eJz631Rt3xP6tPgsQ9kq4E5/dw1
2o6jhaMgWY+UhjFbdbGZbGE6+3wmuixdJd/RDZSpW3BCLL72WD8JymBytQUGfgYE
RjEnz1BDL46Whdj4AnNBMSBlxcglxSEi4drTVMXt0v/aIZJdqzksG3LzIz8Trfse
6AK2Q6EN/t9PpGcFkswQkkpLORrIDmWQpuRhYfxtYFREL7uBx9vIGByWBmWZmvdS
b62nCoj+72oAxggsFYTadHOnwCno0slO8UDwt2uT/UpQSjcWnasALAzyD+xeuG84
Q6OImZRArK22VWhEfLzbjEdxRwc1b/8h/GtDI39qUcfaRoq6mJBUldZn96Yqr82/
JMlb4GlsLLqDQWr9wvd16HKbSEobp8JSnfSnE0Fe/MtTHCIPcRRmkMsezZpA3V75
aePc0Is/j2bzeaYQJRyTKv3buqI+5vP4iMuE3U1B8YEyJu/DZyqkwWmfmToHEk1D
mi+TQKU8lsG9PTJuC6fczVKIOqQc7+/CR97bcb7DVJJR82nWe+MS7hjijFpw+MLc
JYqfEkPxFFZDo5oEakpzR3pUn6GNZ2t175P3pZzJJjnpNrwwexiVa2yu4gqKy3Tx
e96zMXIIAt3oJPkH/0mc1ZE4E/kbobziL4ogC/7I5KdE4xbvvnJh+N0QoDTkG8MB
El2uyxQigrfN9G+NJVWuGAaVySqf1LElVxGZxaoXgLJtxlxyXmxH0YHhFcttq0/5
ZzrkXkBsoHbuocJ/SmFL7yGUkeN4vKiTw90n0D/dQ9UCqx1OWnQ2XRFSOWHMcLrh
blUK6CEugZi4WY76fMZoLx3Ag+X77DmTVFD+1dP5uNhN1e+JewBenFt5tHoXht7n
INg/Q5JF02X7k2+zx7G2//a6XsHvZpZUWQo7G5cQ8cUhqbbnXar+Oe7TNvkrNLqX
tTLasaN5Xk43ZueUUoutcpsWOXMsWPUqRqVP6TdfRwCrKYEH/jcC2FNrypgx7WJs
QBPoQ1BU+e/RXtP1fKDLjBiBT/5gztjovednp/I0+Bc0qEy4jp36G+Z8B5vEHuin
ahIDH5bD7JHZ6IAHXkXgm6aIS5HbQ6N1R0+LizRJrKY2nj8F5P/mcbdTyYZ9BoMo
LssUh0oRszyXjtaQxn+611NP2TEZUhO1P2rYtRcGHcs4kwX3FnWxYdL0ouW9u2jm
53owIAPGURkJiwOJbiOa5Ba8QFxzgvgHykavCSWvaFOblTZFmzHyj8erzfS4DIjB
uvzUJQkchAWjcKHgtwiyFXTVdfZ7eEggu6lIzjQvCpPhVGh6pLSWdj1rfG2QD18+
OB8BKWemtOishVJWe4e+3RWFJngDkjgedoUL661LnxkT/yM3BpBKzZqnRYhQkrdZ
0F51uRRYKRf8NLJkHzdo6TDAN6ZCBEkWIRmZvMvK9J877HtRxYXkAK2mUYy1+FPK
Vg0mwIFPyg9smiQEQrCgkLSBLxqR7JQ5fBwV69KK0pkBnMK4SNIO3FxFBSW0ROqx
DIatWQcj4Tr8BEseZHAeY0KTzOsmE0yzwYQtTPBvOx+Yg49i7boIEVExo7VcjHIt
Ac4NXaXFbEBJa2dywFhfmqz6IfTlRk/KaoI6gD2Guhar/tpRmj2wxcZCowUv/irW
9+gOBtRRk+yuDG39K9tWKuYyaznkFk/PkmGM3+Sw5IMUQKDwZe63BS8F8Dfu+WoP
8gabjXFuGynxvyGQVnqkfBjQwuKh1o4AipJE9cE1bsIErnGcaTHN4O+vtHtgQzx5
GmMsuzy0l95ojY/JHiyEurXiXIC4Q9gmsiRCHDxQGOfzJ5YPR8xwgLsV0F1QUvNP
WBJEUGkuB73JR5nJVUxrzWM1vARE0vYaP51f56U5joJsKt9qNzvLKu+xp6Jc/TZQ
BgK1vNm2ybPm3WX6cDY+E6G/KmZKy58py8SkHzN0+8kpSWp2PBvmfuSV3lVZrX8I
mo9G424jG/U0Q3jg94f0/9C9jlkYYy0D//SxGZ0B1EnDYR6UeqF3wRpROcMIDCZJ
Jrp5fuXVbFhuceMym5o9SNC2tqAcTZ+BtmSLjkTbcPW52cEBiMg50JZT0tc3J88Y
3OGbtLvy/zcFfwM2JtCoo9n55PuvfYvO0cKH4Yw8jhmjCgKdwm9ZVpXZnYuRbAO5
1uymPKqjByM6yVDdScDMIeA4owvjwKcknbPehzJhAv+Vyj/1IodAxVRRJPXu3rNP
uQZwXj0jyHU+duKH0WcAp9UhmHxeX54kK2LyzrXnBMs9pbwn1yt0GioGDWZ7RxUb
LvCAgGBltw0PvkgUVnpLIhCQzzD87X9qnnSE87ll5POCtm4ykewMmuZCxUH9I3EB
gr+uz8hOQbjLM2Bdee7Rgsp28Wy4sxNjdJ5i8a6mif3s3EHv7JDvdhuauNSE0FlE
LQG/dbY9QfEl8Uib9yvMC1QSn5yr4jj6B2XCTGNz7bdSPr6QDhDZ+qiZ/oPNFLdg
MXRrQubC/MxofvpKzHzrYUgNNa4d7OsQae5jcPyBvQw2qLHGBLXcAnC7ifhJnpNg
vcnMo2ga781RWGrJBsT09epXaVRyNgScv6YnDv1rcykJF4tXrWOC1MUydhr5K4CN
lSNM0EBNAhQ8PwOr+JXP3eQejS23cMmuNbNHGpc5EXYVBtppzOyc342QN4OZ5IW2
N1yl9FU1xLm0atkJVULcmDsqK064crIAfaYtiPTtxDg1Mtw5rK92uGKIjMKMP4Yx
9LXAagDDt2spEW+Igw5UFZWRnd+xipDFhAV053qHdJTgZMiMBp44e3TPsGR64eUl
ESzeRxuPaWFAnOHH9pJ3ccwjAJ2Gv0ikTDaHtH3iUNsvY83ONZzNX98vdmZoKkN4
w7RJzoDXtxws8SDnjfJTpQo1v++DEPVhPkYLTpO1xFGqt5ad/e1lKkl4Dbm/EnEx
TkOSGADxp/CX3pi1/PR10F4EJ1gtyw5Hk/bpBvDZgM12pi/1zrFcJN6JofHHl2RV
YI0Q8eK9k5eon8N3D0IBUwDB2x0bkeqWT3WzuwkUGq2k5Y0oRsWwlBkrg7kkvJXH
mKPJUBv1ZNdfUZJdYl5bA2x6sOghjLw+/zMLKeVnldFjT1uX716bdVsGbrP68gLW
1jFul3ybMXWvoH2vK0TpKQrHNlFqOKhCHMa/35iw/AqNGcBCXa+nebmxcIy6Bv8U
a6c/jc6InlmSuFuZ8Jl/ZzCwHbX5uNlWuRT4zZVtkG/IIAiYYHFJBLwqnEchZPre
IDm2qrpmsDi0y85qT8Tq9YLdfBDGe7Eb/U12WJ+PUcHgqrgblzb5dqQApe6a2kRw
rWXzNwSquIfNV7CGulISeNqvvR/vH/6BqWvCwjSqthMrFrOTHonDtFWROPIOnLlP
zsULKYRpyUGJvNinlUh6Fdm3L9Z926aNIxoz5GP57bJcEGjcBq3fdabqcxYBeqmV
KFlfx4IsGLKLtfVpBeTjtZevWrlPDf1ACDZKrjMdM1BpYPRmq3vRnjmDPBfGXi8C
OENNWlwQnQIlBFGTLsLCJYBQy/PVUHloI7ZMMCU3BtmxMCyWwWZNU5HtOExJ6CtF
akUVGndd56yDP9chMUY0/mFM5xIwZZZp5zoy3r5PDcfBPzC8y+ij+g30vtk563jl
tjv3Lx7KoPY1iyBcPNNyf2eCB78a5h05nlAkDBSNyp0660vKQTDEWaYfb14ki9JV
bJ7Pzba55SPubpRhpvbH4f8UR/ECcTt9qe2NGtufzJ2dvLgUb3FZQBQjcXOzI2aJ
EAolCSMaqmdZAkW1pTzVoQbwZ2UXbMQWhl6b2LQ3xQq0rr4nJgw/xCZqWgyDDIyQ
9dVMWBXWU/cCUoPKp7qMJXL7IqlLTt6bDAFEx+HXUsCdju+Ptwk1npGRk8OvBMxu
plujarKoDpyBLIqxg4678aEFi2ECzeRDk6AGOj+BSmFNNb68pDO2Wenac1wzDDG9
QfyPrvjnogHZ9EJiIi59bF0lK09L8BSrcOeOCvbhZiCGsslTuEkuHLlHAVe1hZD6
U2wKDdWhYVVF59uvxKAg7rz9Mb9cHn3zt9kW2EBPE8MsBCRK+AzrDJ2hx5uAIDqR
XiwksfhpcLGHQDkiJG4XTtjE7xCAtf5mUPNnVpmXzN5dw7r18JO1cg+UC25Dh7bT
e1NFzLWI+AukZHN9QocqiNkWH3TbiHGy2E1xLn46hgbZH0hkkpsrlCAvPzYgKGoW
swm/vesFSOziuWVvPWmBOwWSmhZ4N7nIClBfCNndAEQoacGQuKXXzwcPONX0sldY
/NwdJOq8Qni4G4wg3dfY++S0Rue46JPNcTDkoXoKHdl41UbqgObfvWyjjY6fv1bW
MD1NNF1MVofub4NrDCk7It9j5ZehGpFt9YZ0OLyw7+emJViqbFDFJaivQSyhkUkI
0RLAnOvshcUsKCa2rKByyavbjfWn8Vj+tGVSPM+lxQItr7pzyclOQDUEdsXwBHzC
VlA6fcAOmjX9Pi4sK/sI+RAlyyWHUsS/M0ssJfu4f7zoy7p+wEjEq8/Taw/ymxsE
dfnvoWMI7SXdrrI/ymtxD5hhl7oeB5Zx+u3kd+AzjdEC657iu8Q5N4qW8k7gwZVK
pHieFG9KMX8juMrSThwYPsksKufio/5GXR3HC/pfpyuzaHGJtGesXLDkh6f9MYJo
s5GLOVjOLSynLrGyP3ge+7tYOqzJU+oQN+Jw5vUmml+UlbXG5uxK9n8ODO+deg6s
Lp2xCCmceiAXLele7ulZZTwj6zI82wvg5Nn2g1W47rEyYc/x5uLdZy3hTYAZpY/A
Vr73pfg3oG9j0wKGz50OTUddds1wwbvHuAkQKS4mhrNdrFRcuk9L5mcPo83I6HvD
7yGrJHQB7riD/75dNZHpEISWCaq3h7GtGpI2xEF3vEcENGSMG2bKBWtTulZI1DBa
ixd4NHM9akKC+Pdxv6AtGs0nqw/WAqJtAZvz0B+Qd/rQuJkBm94qMepnxyU/MLBU
tR9C1RJMbBLTXeKwAt1pg9YaPJW7v4tVZrhB3jvUQxuUEhanFxV95DGEMt/moY20
6M5JbYCEIkLdssq7skIOSnTx/vWarvX0wS/EGo8lS/uvoRWBPV6MCd1m7DitWSta
56Kj0FhkB5bHycFCfA4m3bXVm5De3kxQzX9HHyzUh4ZHHteJN83h/vSB/nblXnVr
IvfFeLmw4kJAIeUA7JC682TxSyC7V/iM42hSt5utcSpHlw8hQg53oYOIAYziiD97
jQNX0fWZHogfoSY51KEqSO6M1TyVJCbsWePDhTYOI2xv53xKQVssDQ77q6GAI6Bh
zbMX4cBPF6N/stGsCmPWSfBRudHryHfr589FrVQentJejLDYKmOaMyYPd5rPioUK
DLKwq+kSw4EsbJqMYPqiVSGz+LNxt8SD7yDE/wOPvA1fkJltzUvuxXgAwxRra7T/
0/1w9kVpBv7YLPPeN2dV185S3rYX9+gXJ3zkQoghVoYi8LQ1NO1AQpbtluJkS0FZ
dIbkWJh6uZnjKMq5rAaL4nzsF1Yjiifck2vPIJcYG4FmTbJaRyQJjXZlvNWa/dih
zBgm4nWCP0TEbXH7yosPmrwZZG4EOMZSOH241+onyni3yk3tAvcNlMr1CQDOcyog
+qle1nDcO8ycSUARhxBi8FVP6fn1Yw1CZylpPiT1RyLpn6rlueKPNIk9p/yrdu09
9k+zqKak6cdOSTu8ZOGp90m5f7Q5YD2Mvd+kXkuh9QwipQ9J/AMZnrH8ekczmzZq
diiGgsiQGLy4EQwnoyDAMvNDaEucUhWlnUkcBnzB9B7iXGUqAizsGLYcBSqT5VT2
BLnKs01OCKLQceEfC4OBKimmYEnzaJ3whNw5RZJXg9jXpTiquW/qf+gBffZeLo6d
Ub1y36myB7Eu18JywjjVAa7Yb8cKR8uVV/01x78e81zP8m4rWphB7KliOeq+4X7c
I40dAGglkfQku8iJRXmn1SkjjdaWf7YwgmlSw8DYNEY1SOen07CzUuNMNYZxVG0i
mPF90YJ1uNNbst1IDqrLlqasbCjaRxuBgu8Kbmx0lSK230M7Hd3IUXtt7EpRfIKg
o444Lp5ilgFOE8HQnKqTXg/R12tpj87cLnOAfS/P+O1FLJudbu/tb3iO79NT28lv
H8I4gxZQ61E2xmDeimcKUnSOESkRiXzF42HnYlgGe4DdDfLu9jqHeSrIMU5asg9U
9hp5TPZ+rV96pnrirkcIOkQNjpLhZQL8sIeqNZU2f0WT/VjoYpBqrXMnLKJwicmI
Tipfju81Yx/g0CfEiEYHiSgBaVEjyBPMrhh/6RUrW/6WM+UorwTXn4jXcuH4+8Z+
wGs45PIWvH8+6+NUUpqag7rusKHvGjG4UpugigsbBCK/Rs9OsCZMG24LkFXSQIS2
EvEi+E86nZvKkmNr6aqccxLk+IgJCPEtMdgiqxfDgOPHs7XI969Wtw6EDgRqXwww
zystbxhYCPOD8uFoARJeOYp1uX2UCLeqQkj/5p/rPi1pQvvUzDpM/wlSCB2P0uoV
H9l+T8f/JwHZZanCidSZ2J354zcOJa+Bp+Mn5zrJfFXFP70QV3bvIyWZqTNERpZD
4ZEUhmoNSbz6KTXmrRK0cc7UNP2ZnfBcgQyIR3MR6H9UkOCyFDmGU1OsOTp/ILJs
UV/ZLho3Y4576uqW2D0PF96y/oTPhjk7OtauZHgX04ARf3mL4jRj7JNrJjFZ3uv3
MGkQ2yooWQkFlABpDFccXnDkoI4V06zbmQtZSMBHydi2g/7AzmqnGeDLcCzPjSMU
RtjLnKXOZA2Nbij4Xhk4OoNTFkVfM5070ukc+20nAvfYwwzqJPcu8BmvqPFm+Lb+
q6K7XihWq/qLZxjSy4DH7I/0rw7uoWPUvjFgNL4NhBYJXNc8LlDIdY6WkmSsHduM
Fd2PVV2JB0/Iz/wHaZGPOPOFKDgN4iQzmisYKIv+j0+mTadzG1N2S2Qo8IJ8WDzZ
KIpjatT1i+zg1U7hDURSFGYjJxMLLFDdP8bizNlyaDeBiYbqLd0MfEnTn1F0+472
1eTMrKm9avMZ4jLyccT9CR9L3H9R5ytPYBydbEH4knOB88jH5LwO70TByq7Dz6JQ
Pp5EbAXZ7B1qtg/gyXjsD6vpZQ+Lzjkku7TI3P/CdrQb/O3QUENTatNGl8H5wep4
SQss1GBKuPPUrsHSDPhiLUlxc9rN0d9ER/Xrcx0pSmJbvx2pQEU54MJHF/HPuERm
mWIoA7In8n4ZHu3VJ2UgjcqnbU2E+roLM1jVFeSARlvn3FX+PCpLbLPCpZwXlN2i
B91OAQ2w4F6eyxzUSBF/hVCxLTL9S533gpHXCkWCaBQqg+PEFELGAK5m055Z4EYQ
uJw/Ga7z2uqCjcBadJgizjT7O24Lg+yU5SpTvj/WCqe2MR3cMMUhe74Ss1morJWL
5UZzxLLX0oyiaxD04H6JGJXpkS4hT8BQGL6hyyxmGphPQg31Kxs7cwgUXrjqSS/B
n4Ewyq0JHMGmOvhy86/0rsho3B8rjCAIZUEdrLV7y389IDwfTWNEX3v6xIldbl0z
olW8Yw7CSoQgOx8ICxXISxVvoN6dkOhB/c8mLLYD+Sq/nJ2GIWGXtg+xb34vFnPh
pjMUakR2O20lgJSnzTX0FtulSOz2dU7OI0cuqOwGPXoPHTMFoXDYWN479WThO/h3
5QepeZwFwYkG7WBXuxPuhCSPzwFZ9MD2fO1O8gmT7bUUAfTHC09Q6T53RjhOv2y/
iRQxyBOBJNxdj2Ma6bPZ9Jzf+Y1bi3v3cylYvSjFvjk2ll53oIZV7Z/bIjLg+KD4
rGIgbn22DeMqWU58xakGWFW0KhpdUIijvj0XL3iV22XCU48CKh7ZWyI0BhYbmjGP
WGMu0Rv+AwCbU6ZtzjHu9DWcMdUmQWIuRSIp29kAfL4z10O3ii6Sufd9WHc3LjXf
ulLEcvYWyalbtvIDoQ+FKTy5YckIUnvhzUAftkdTlgZusPaCe2/8SOQnqDcZsSXD
E9Nw4RaGSO8Jm0g0AJ5powKQoLs7It6JwmEN3c35GkSlyApLbgzS9+RlEfJCBdVx
eR5va3mf3We3lx7lXZmtYKFx9ETUvITemmSe60ndzwFKITXH1ZerMC8wgaYeQ0XL
A6pfcgjDviAn+R7NQEJ1UsfUtdhTj09jStWcWyTlI8qoydiK7uY7MF0CKWIrJ4my
KF57Hvlv8umiVy32hak/bHRntG18zV37HJ9Hdhr7E2D1pF1kQSuujxwwsAyBFAQr
1D5QKJ++6Ms80Uf6Ci5zis+z8B87LORTYhPCWqQAA+g/4UITpRuiVr7Eza2EcHXi
G+7Ja0H/rbWcyNFxc3NwxAr8W5OrF7bORmVvhoJ6OoDceguUkjcHwoB9WFqIgkOg
RFbYplztxA1zgBZ5zxl6pi1K9NMjnS2DMR1EH5vLwQr3I3vULhs9okPYuRREP4P7
5ssp81fye7mq2xzMkfNgLH0KTDV50aU8HeTyw3GWvkpOB2266Mui0hKd99+XDluw
Qgbm+EtVzsoopNWimQ50xUj16fw22d8HTCaiLxrPERpzaKb/6yqew2tpmpOvSVbr
e4zH56J4GqmAEORr0zF8pmToJq2rv3DuR137BdvOIujCkUbwUWlEZWd+DOq/FiEx
IOj2cVhboZtG4uCE72z44RZeET+9NMXVEhSZU5Veq1A/mW8l1vOzcZ8NUw5gHUHR
313DLB4VYN3LsYsTpJ3qWDL7gs3N1jNGB82F5jd8unh5hyx2L+XpyataRTT+f1zB
HhPP1i/dlyKtbcviGQ5LsbMRU77Lg1PvcCIeR1Vn2qKz8abvtDD5g+y9tjQPkWpE
X1SKbUTQVxnmpNKX1nGYZYsVsy4uBR2QPdMJd0l1iiybPD9geZQjF7KY4fuzQeT8
3+qRyJhJX/IkKCDwDEkvZbEwbwewJELF8dibbv65EI3Kaw1X0WiAjHFhQZ+T2a1y
MqFTD4a9PMKWzVRe+dtkWI26Mz0WyvhsdV3QtJEQJmhP3sB35O0nP+clPdsiTGzi
DcVlTqhCgXTOlpB/cECmtotpe6RyU+NZdS6mqbYC+YsThoqVpXVLoPbwha1jznKV
ABKMRouPQD5blZm/4TFGiPWRGWtaQ3PEZbwvWULme69VcDggDz66V2nNcC30jwkX
l6Q6gUqNdfs7bE3nEWfoMqmbeK1LTXGhfTzUBCwrB9mj3FLs8IWn878p+lChvFqc
R603xRio/h4rih6EtpxR9+qh83GzAwYWrOTjbasoYD/6fjrcuIPNySIhJWnacd9o
TtL24lx5ZmmnjE889rw6q6M7iFAC3+tPu6phZ5FdOOuXMRQVdHE/h6xaXBr4D+CX
vr3wcmh/asFICjrbVbAcoAhKCG5d79LcrgYb5rWuJ2TKeF7bt/k8+nzhDfmf9hFc
CUsEq1Z5vyZirbc3kVY4zEbOXCe1CQBWMq7JIsS4lfI7itpNK11FDzOZ8gA1pBpA
DCijzaTnIQ2awoPHqr91dAmLiW//uQM93zDcl7I+6VWvnBK9Q1K41Jxhz60F7Ati
hRDTY0dayKhcW6/OhzyF9ORI9963OEO1tztC480zlDNHqjpGRBVtwaCYBHgs4v5v
ofWtUtL9WXv+fBqO4tBN86cCU434k/mtG+2NWdA5cUAjlQvJi5AszoN8UMZF2djB
uC0167+08fx8kXBPEslWMheGr41AQ7zafoUzFR4UJizZBKrcux33Naf3fh8hgz0U
I7DA5h2TU7Bs5K+uNAO66He+rYs/W5/TkHHMftJMG6JjWuJxMOcM1pfGywISlipM
q/FjPlrEtnWVB0FRxhlvl2pwh76+elHuYlH7w3WUVrZccwj1ExwFedwK8CFcOD+R
NhqG+VHnXP49O8wZVD2lnAiRw8ciIuSHjbjtBcjiMj0xoPOGlGYOB18ZwI1XODt5
1TceEbRylTBAo8/1ZqlCNVHY64HEuqeBPlBLbd/hHdGts4EaLI7n+uZwBZeXM7QU
BYLioEyRXRw3LkBkY1baMEu3JafeQWWUazzeCSjT0UPkmN1Gcsh02lyL4xHNKbTV
CJ28+anY3PJxVmukZLvzg8ASJV9a5eObYR6TcYtYlzNO1pZUHExeaaYTu+drTfDl
EXtbiBjCJC1n4CNp5dBvcXF/HVUVABD7b4HBAiYfwgnTl9yL0oXGaSijANqZmT9T
YVpNGw2SRrZaTcrvKoaVsEmWBbs/g5/RUggoMVATh1RYU+mOWNEf6KQ2ErgG3mfk
t94ZN7IMhrD4uXG3Dzvavxx+dWEQsAZU4m/0L90URh3lsbaHfXgMuffIMYYFF6w6
dco1bdNok6xfuJoRDvG6kqd6AZwJvDMUXOR0sTRTQq9fF3Ebn+mEm9VHviylPjic
KtXruwMXaIFxKuukvFQwEXWDw3T1RhbnMNQR80mDfmdXotvkgYPmRZVX54SGUE8H
j9bM5WE3DV1yODewYWg1o+X+SLpPAFmcc6o77sVCR1A/NeOZPABkn34KESw3FVRJ
fIhFNxhp8lf6Pkd8XzhOpRoy7HweB1WaFuhsKOAvPxtlj47xK9lCKhNU8aPKT7NA
EexKyeWFbxp+Cz2mN2/bkb2HvjViQ6jSrDAJqWHUIlqhmA4jJKjh47gG4NYHJrH3
dCmehbEGiZOqIJKgqcYpIcGcloCwOTIokNJDxFPWnJpDfnjY8kED+1JYj7wilDZV
0BOZgqK8rMPJ8YXx3q04H0Q7u+8R7qxcw2bbcgpAU96bCvebY41B93qi2diUHqfp
qtntGhHAhqUtMjv5IEfVMbY/bDyr0hYoTT8aHJaqElsPBiBmQPfvdhPck/oQjVCw
9yMYuFqnPs1HaDJ9Q7VXDhmXbj1GxF2RLlb4mmHJ5Nv1FmPvsyKmsaMK3/kgSa0S
YWhIt5+m79Oc4RExStoRGq3W9nJmyyK4wsTirdYheMmZGzvsvhDiZg1+hb0unG2a
fCP9+dwYpnhIhWmjthwrh8xGTO4NHY4YjkAxEN/haoL+6W3ouAnzmEPzX0N29+V+
cZqlEKjLEDUbVugyR0csGMoAk5Bzc+s0cN+G56r3ZUgODnTxPK1sMMrm7SYW19+K
Z+JOK+cH67DBFRvNywbcZo0O3rLhdZqXV7hIiUp8dJ6opqq2EyKFqY5eoE8lcdgA
u25679W+v2crZuKTEFAVNDw5K2VNrjlqjIIpEHRNCpBIsfHajs1Mb6Irf/O2OIES
gQIIagYG0gTG5TvrUPTnZYqg2GTpHkFbiUCouhFaZFzL3HIEkTXmDQ+6tmDDUnjE
i4NgbfzrxQUoDbbcbVICwRfbhWJw8/jeZS7H6RO+AcXmROYJodDCqKd1gaqvYqAZ
+TTmuQ4sgL7K5xVEtplyDaYs56ytssWgl8Z5JOJsOlld7Uaf9/qspTiHawIzhy+e
zY2HC7LVdu43aMGUEZcJNBvRF7nSRZ7opXomnNF6gBfkUQYq1twNqPpz69naIa6Z
srYXp2bbfDM6ll3jQZSGgS5LWcznd4wIoQem8yhY2SQq94FSrsuKnUEVU+Wksv9i
P/AAXbHSX9+TDjSCtnIjG5k4qPjPzrDKfb3IIAyZLxj+NzK7/KDyA7SXHx/MmtYc
TsOUuDNQHBFXxLq3Uw8jCfGkAPAA8uGaPIlAg/a7+ismu8YJcyaXjdQg4HUjvCKB
4wF8OtjbTU246pVLnYO3Q6PyPHW5VhTaB6ScN4KOxyHhD/5zA+VIJldpMyfViH8b
yqY9z/dnv9DuPEo0B/OlhxFgM03wJ23wfk3UYOo/Fn+XGZReypyOVFq7+xX9b0oA
CACfeF9HqrXQeHbl5c6xAnWWXDdHmIKKqikfpk2Ln3ap3fcQvV4FW2tyv8ONUi6P
i9gTZse2ol+zTnvpp2aq++I4EPsAWxFpvAGZJrPezpq65e9HsevPFTd/DxkbzSBy
V8l4jD2wCSjQDGltagybecpOugQSwkl3uKMQRvZL+Ynh8PGEVE1rkzNG7a9h3WRI
2EfSDb6sOUBNG4Q0HHikEQ64KhX+s3rB2Mj8eg6vjJotX9iieAkuNzdX1nCBVx4P
dt8aPFWQa9D5NXKhcc/n18drfbk8VlgqWDdmbU7udIWYjKe7mvUDQIw3x8+Q3CHF
fhPJaUhh3A90cctnAG9qMUhe3611Ih1NwUD/FVtV6jk7fInmvgSn/AA20aBXI+FY
CZs+7ieukzyIsxY0phlmMtKvQCNRQfvBwXU+svJCBEZPq3VG64ppkIMjJvE+NQl/
n0fqOc+Iyb6CsTfmjxruc1K+G1x0yPlYQmnsMZ28FH5OMw+qr95geDMkpL8PEPL5
csMmQr7N2OxX6MBG62hXws5niZInGtQMTYeMGI2R2GHfLScpLBcxa0An/0MVJwtE
ptLXQplSJACOu9vb+QXagsIp/QED2lURuQ6QC92KmhlvboS/QJHO1tI3lW9b9UcN
T0036dIP2sdkFdN0tn1mCxxw0pCQErN/pUMhsLJEURGAVnOcfSNhDG2SOPaefbc6
535aZlQr48IGr/O18UNswM8MMlwawWivT2B7T1KNQlXKE0b4fd89/5otmnliJpY7
GDBUWLEnDxuHWRdWq4TT9jtkgufgOL7VoE+l1gPRZq1u231OXZiZkshhwR7b+dMl
ga9ou161kPMJH+DgYXrr0RGg9yr/RGgbf5EJ1eKR9G1cfetGmtOKdez7fVM9uJu1
PSLoqvXnaKRzWS6i6ILG9W2mjfvf5TucYqhuauG3DO2/rzBdTUXlvhrmqtzOTLa8
2Ibr46UMwzKyoY5Z34ValHaA5apaJGOovgD7ftsf/hQ5BWzDnGz8sNdAlEcYjtc3
kdmM1H5SJ5w2tnANsKG468kjYBAp+ElKQe/y2CbUE6Pph+YwGtwFooTCcHmlV4Pd
xKjhXvprhwCD2SZaLkn6f/vhLBMFtXEX+uqhCwuF+oBjzzJUAJsdwiPTNw3A4ZKO
WTlnh9FoWLEIaLLWqpolIwpYyZu4X08KiSSqTJb062o8FRZt503uaTWE/yezQr0R
vIppMrjZZIR5xkDU6WB8zcyv59/AVUAK0Au0W2pwhzQkwokwXzoviUG05sKwrTAl
7L2TgoFn8/ikPBuqj9CN/XvpCyqGamjUjPGBMGVVaZi5zmzLh6FiUshcUELCzMUi
0y2te4RATegbcCc1ESOPRsSiwdlYiruSnqSIkE8tcvOhcGHlLMdQhJw5tG+0gBAZ
k4jaITqG3Lla+wmgm2qPitufuRbuGttUL61h7Cvifu8F6ZhEy/4egVnEZxduslYv
krjNIIVrDMrbFlgQ1J2b3tDjysS51rGNy32YGT/1cwE/E5jXH0Apmd6xxS/scREf
6JDrSBG+8ZRbCAeRKsV5EgqYxn84rLlYee048q9XnwdcE2jCwbnJML1bYxlmC8k3
Dub3f6HD4SxyX+pve55ow0/SG1KT89XPgzV4hhYx2X1WUcPXZhio5+Drcuu40rmV
vn4RbdCQqcw2opHgnpkdlzNW2aErlAGNG2t8keOEcYQAL7zkoL7ZB+tlXk2uZ0VG
s6h4LLXVI/g2eiXs0kFLl0bUU95Vf+6WlADk3jNjfbvfr4YArrZ09YbBWpjVpQ7s
ty4w36n08aSyjAqLc+t3mIXZD5JImgyytc6fcGcw6ZxAvw1xHxH5eZGPvZIYjqha
rm1jdmQsafr0OCWpdzkn6c5+/04xViuRr6phZGVtdHQD0ek5LKANujpn3Ed/0UAu
00f3FAQ5+oSONCr5KJeUAQP140IczH+8UR39keRZy2Ar3cg0lwSNwkjNZynGzTQB
J6DrSOHoWVSHupB2z+em3jWyB922kcFKqxdcqDYDylqEvyZO0wxNtjl7HrNbWktx
hO6IscLWk5Mlia/+ucfJ6wM20V94aqVHy+R0jaOAKCG7AJOrag9zVnDlFjeMl0fy
xCcqDSWiOSxre0bBh1rr4WjHYcB0K/u7Gkr63YzCilPRqsPadQMtyXcJrn0v+CV4
nejyzQAx0tNx73O/zWogVmjV2WZ1YTwH1NjTDSQw+FEWHhUJBVc+Fh3o+WkxCirB
RxAf2MwUEa+nnlbYurk+Wq3j5CJpQauIvViyBrbQa4vq9vk67d7Crn2eN8oBKqCu
jBDhs/0QeeddF4EQLenY8ZJVrtsqn8iIGjd3zA1lQ2dcaNaz+G5RkeJSk8yC9Owd
V+JYv/7v28EWKuDmhW+bVhyGzCDUx/GpP92MdUh9pA62DgQidKHZzfTbGpIbbG7l
bQfu5dQpDXj+EzpD2Pu1uA==
`pragma protect end_protected
