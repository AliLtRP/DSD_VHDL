// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G/zTeZcpZMQ0f8nTakMjp/NWjSDSie8QMvWvYJo0/vJtqIztj++XavKSpm8tWt5A
JZy/ApBa5yIM+EKG65kg42gKY8DxFmKKT+SEPnX5D7AV/j5CITZSix5YXeeOxTTQ
OUmxh7wgEqDiKV/w8tiLhhjeEUS1ySwiRu/5FdkchkI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24752)
ScRt6DWOptt5i17XGhZWTGEXM2dmhVzINLsGTmj1MXfFmQ7Mm0npGFYQVtCn4RGU
UYJeDORyhasWJ81ke4GchkuCmuqQ2xceXFwAs+fUffUqdhQ+pEcds+0uiSJewjdv
XJNTVg2dxkVjgxAbzSERDx0ahG1NSSsILT/Dzy/X4PJcuG5GV2yTCSa8mXDrFI/X
eyghUKiYl0dDdUlzqIK4qJSVEaEZrsWgzqit7BqIhH/fM0e/1rkpu13nGZUDTHj2
bxhKL3kGVnjJ7Hs87R9C20p3qRmuHYy5DZi4hywJYxVhuX+RylFDzTv/tCuytu3V
/kDYq1mMNLMsBfHRtShGmyKQtbEi6mDq+BEbd5qoTUELnCefvwyJVxhoyaGxPDih
hlWkUtigx45J6ZMoAufE10lTs+k5yzq1v8pG/zpHWU/znU4xlrFHTOdg4GSl5L+Z
AZhTw8g90HpKm8LK7pwY1F1MlkXo+agMstVU85ScQCYP2nwAmFHDuJSEQiFA3PQF
gzz7MjlLzuc/dkXjKGBbk4hm9HaTBMJ0VpQSFEybE6bsUcD0f6RD5eU6ZXEeZb29
9c3Bg1q6JDNUDlQLK+Ymf9cxwy+UZAz+b0QbFlvjyiDRaR+jj0CQ6byhrhwU2rKO
VYBCGqxLeX3iSEepuAlz/L6PT7Dkz56cWp9gUBcpljGxfqS19XteEentTmIT2J1u
GRKxBeO98YiSHNn9lM0Gr7JK3uAHdV7MzpfV9B9PayEVNpLr/ZkmEnvjk/Aiwrsg
u0b92g1u5CAVAPDz5OMknN5s9XTtFkh6P8JpUbg57xX0NCjhW8A4QSQISz+KTjUm
BZNNgAP7W9v55zs6gR2m7wd7L+KbFBX1NIRejYcUd9eusdgUvj1QSyoCcpQH4GnK
C4j6Hb5QdAQk/KJvTuzHUnk1wvkJruxU34q2HGPgyAV9wLw3o2Uk60fu7/yC48aK
WwtgTQeM86pBi+GOXKw5x3GoRqpxVgiW6xZiAbj8ohzjXdllL0HTjGMWgXxfnYEo
ltO7ZUuMeJiHzqIZ0u3kTlyt+gC9oalLovTLHnA44s0xg7yN/BvNiAXZTMDSfNuc
BKiW48ojGmDZSR0jjTiCS80Wh0h2yOL+060KPsW/qn34poyxVvn1a4BYt/+iAIMw
DPmSepOE04Dwa8lLol/8Cbh4SsTy9fQoUjlFoqFNLB4H+2KAJAyodX2emor+xpEZ
1/ItdGmnjpBCT3j+4hVe9EnCTcU+T1oLQ7ITpnnSzeVru9vYwCGTmC+C2Ahm+3Jk
xNL8jrYOXIQ3C2v8zGKnnq1gR2jnE30XfhXuueabFVkY7UuhqEg5a5rMcVORP7do
ffGiCjtn7847cgc9FRTwkhMTlgwlzBxzmthHBCoNs4KFeLcwzcStVkyrJV19irpr
PlWbvMSBNrQqGlqZ+cwVSA3aDMI7hDJdxnlh6wfSUXsv8sX1mFcR5aLHXmpJTnyL
1FVgGf12zI5AcnmWd9Fh0170n7h90EFkwYOD1QLpSI1vjOQByoRFB81ICXGE16+R
0eNm/eqM1rQEnnY+e4iShFTQxaYnLNcio35ancVaCSQh5jDdHCjutJjF1JP9lhIc
4DZqZIjz9kLhYWNbFzPdtBkAAv1dMfF1hc4Vrx1IFjZfJ/RFObOTCy0pn8d/HNEE
t3ClTMP95fcwwGLBi6zYQenAhJWdx3XomJLDJ1s15d9yLlqAmsROYSr7Gzu4P42/
/cay58JqhzLEBSD05HFpONE2VNtZRXei8dv4daBmNKg6NOoE+dHadvaGbgWsSKkU
SNgi/W18GFBmIfwwul3GZ4YNBtrKC9t3EY9DniFr5XaaPll8FV3182UBKi/tut+F
wp+r7zJ20wmcVIWPSpHfzAFCVGKOvfqs+5nWlu7smJPpTj5oz1K1r52/rnwawH1I
8STDurEY9/jZ0RX7gFftcM2mCD6AeMIAUFcf/66QhfrzTwh34gJFvdUEsuhwUsei
xUmksgorDj6fZccVlS9puUmpY/V+I4cR0VLIIg2hQ/ZPTZwRY5XdLwB8/F8gBwjk
LoABzArVjATDY58R2MKwt74aEidU8vsmDv4QpII98rgTSTiR6J5TtNraSBlBV24G
NjIUgAB5awPmPXmVA/Gc7Oh8SvLVdiISG7VhEgMvNh9jQuRqrTC7pAECJCPN01/T
sRufAG9ZjaIDYnb8Ig0MRdWL1JZet+t2HqdMhNDWH0/eyGO/7pMz/OePOiHK7CZi
hiWC/upmH+3AdFyQu+F2g9JDku0G6c09T+oNra6W5py06j71Y0zvHhXTmDiAQppZ
yx/ULlXO9ao1pdJXFkB/9hQ0Eet9jWtKkohRD1o4C2/ilqbO7uO40NZUNkLe7yOk
OVxKjyo0NMtBBntut1b+QqKq0Av/BRlALrphvEFte0SPiMUffra0ezjiPJQnJKr1
VZhdzUnLHhbOqWL0x9BXCXzHJKKtD8bik43fbQNuJOQ1zzHTfHRSxIY+pCnfG+gA
1F3lSRAuPXCz2wrRpCYnRXnWP9wO+WMN0CtC0Ffxn26caVs1JL+KbcpzlXD4ao0t
XS7IYBwM6Y14Q74vX8ynyXeWj2pGfTRhe+UD4lY55EI73QOoiKi1hZem1vhg1ow9
/u2HROzZ5JUhyBU/yfb3aFHzg+NFOpm4PHHr32pWZONDbgrRweFZKMxtXhmmuJci
x1mKDOC4UsY63sCBKOr1yqzCR+EnFUU3kZ0+zaL0blAlyHW0RoInOtRAQls/ZzlM
rTC49WK3ySxTriCD9dWkjQxMbdx0NRjOvm0PIPbBG4AJIEUL49QXIxOmpi/bZKU5
SV/aBCseYexF6uUa1h2OYOw73ZJTxZ+dy7QhMHv+OS+JpobPrYgK7t+zgS8kWtae
c9ZoAl505+irmkimVFe8QAT12KjAU2nAMHLtU1yd7wZhy9wd4+a88ovtn+gng/z0
h9W44N8y6SpEttsT8NmJQjc3PzV8/AL9M6YgvMs0Waf3Oa0nX4J0ht3IUqzUgqao
0u39iAEkh98KFzfSprQXDnjS9H9sovVgWDXpDqHUR2HQW2tqNwo8nmyCq3WQjPAY
R3K9MZV/NIbs0Co9fUaAmI9jQrnwz9+zppZ5+pMPRztNkkxTVJ69bFGMwhKDToyD
SWtCQoIHUN/XoLnyu37vqxuQny7dkRgIU4uNpVL1vtQLlPINKEpUypvC92JrJjD2
A6dMG1v9pqC68/lhQLRC1Vp2chagCTG9Ayzy0+NxkvuonGJ5/xwK2LGvbRmBX/om
rOSA8xYFVZ5Ocy2/pnuPGxNcrcGznYs/GJoWO2M0NxveiXcMrcetLht60xIqTat/
DIQuMscTeLUHhy4H7GZgsB9S1gqZu2JfP33pv7NMA9VTaVOCI1L6x1w1jCTQz2GA
5DZPa/zP0xiMrxWxDYS4crcjtR8xOg805UF7t9zFJkVXj9HVYTBgB+ZIVdXbiKah
BtmJZRuHie0UzORP6vvzKaSdl/CgYZXWEPOKCZZa2n4tWbBnNlJmdNrTYP3WuP1M
FyRdOzqg+mLVlK+djb3cLdHECaDQCf+yK3pE0e4gwh8oBWuClywPuEmQ7z8fwkuH
zLh2rC+DeStF8uaOC8rHuSkotCjv5M9ufZZneEJeUKHViUgJ6T9sq5wj8aEqzFp6
zyRwNKWjzHJ2zBxtdk7At03/9RXv8GUthho7zs7k55tMmjHaBg6mqIE8hZ1BRyD1
y6H1Kswj7x3arYHlRt4z4KZ+p4AsXNrgrz+CKaOsjcIrefpwTlapIvNEp24r2CL0
gqBOtd58x/90gzmskm2aiq7yq28iFBP9GIarXdeVGWviYbICLmHMXl1hMtPA0kr2
GJIOM/IEpj03jVkZhseDyQm/h8hMPNxemkROMfYK0UjPoWFcayWdUJN6MQEW1CpP
hhEU1eN5aVyx6D1wq18Wd9+oIguplOEi9zAFyS6sjF85Vdj9lKTwS0iWxAkn5aDY
plOGXEWHzcXgFUHHCU9h35pIXqOxYKro/Uvshi3kgmpNh+YYqGQoF96hQLCaWniP
GFjQdobb0wD5lVQZN63iN2Py705V5th2v0qUFvJ6TvGO0IBhqyh0DdDqa8LyNGKg
bcB3KW8+q3eRSQh7LuhHZI1vund/RANT9cKwz6mx/p85YJKJ2oiD0wXxvf1gaETm
kdmqyJbr522Itl2DmZbGorRlrUbZh0p9qpuQcV2jPegADJs5EarSaCqScpDQUWQM
AxwjZTX7YBf116sa0oKcyy8RDdTMTcNU2OCM8X/xuj/qiEbVAgpMyOCU+HI53t9g
F5i8JHGI+1OUr9Vy+oAwweWjLSEvZI8zV1wvps7mf2y0QIFidOfdYp4toh5WcXtL
tZVrIC7gPimHlfpwPaBgU/lKPlEnEwdUGL1Ia/4NAH8H8oLNBhtQJKK2QYnh5R4a
ImCD8FZZBoA7i4js5MzM01HSlM5xx5XIGoAOiAeDIc4fj8r6Z8YOleW0o6WA0HxU
BxyDl/n0S6W4zFGc24y7RibBCueVbTTQGYs/bLXRMiLaqQUHTTNXapSSB26QIhHG
6VFLb9qtWG58293li/AivrkXMfJfyXOP+IBW064lTKE3c1lHlXmQzeyHSfjYWrek
0iv20Ht9AG2Cjk31UJKkE9jmsAubAMezXLrhMnMG+yet+j14k0InQk6k0GT1zJ+e
frbhOVP1N+JorLrvTu3YERU6Z4EA7kaCtAe95f0ipJv/GRV1UIO0B/4/SmFUi5nW
yKnS9/8EGgr/EKieLafTbohSpUgd5iaA4Je83iFWpwaMEooLPHV759T+7uhKqlZF
WxbyOmoXdMrv1HjmN3Hb1iWRpX07Qh2kL8/NEj3SdLtBIhSGnxj7EQIWnkrh+vI7
uFkUM9jvo+Tn6bJhR6Lc/B8BIxKeEXKDgFO30e2+OUa3aRRFH6D6pLyvrU6I+RbD
9ysaocSavUbudYzD/L4YBzgXvGscYeQTf2opc5ZlWGCt+se05FRCfuWX0f3EX8yR
fosvnUII390tAAh+tCFhipb5X8X4sY6ZarZHptGHAVEC39pc1vMwYjjI5zS5s3Gn
GMHbPR3jm4Xii7hGwI0VnC3Xdc2xvXrdNaWdGZCxm6Api8Nftc6/273kFghkYuic
VIb9AYd+5P5pVPPPhe99xssaETV2LHTQ6HgmsJmIQui6W6FVgP3VMITQ1NVp7FSV
mhFDGf5cu9Jc429mcY3f37905krGLqXLI8ID9FBimvCCVdegQe5sUwMKuNBptmuP
epKTbhM29tnowUG95XMHiVNtJqD4XotdqUjprpkdbmjXu8CFwnwRR/tbaY7b8+M8
CgDoW+UCZJLI5UhD49XStovdqeZfV2JNmP9Z/nVjlDuzrFg1l7dc0MviqdQf3vTU
dm8gN6JLVC76i7KpJICTKuiPAtjWxN0ko8ciG53FvXI6MJ7nAa84q/sqNuuTrfGX
7bben+7VdW0uhRVgihXHnICkkK/gpqcDhV7E/ApCcZUeMjjYREMXbgrmnFztA0Tm
VI5uDVKPBC2XnkPq8haVyIrcU7qzXQNkN92LAHvJwWA4tqwI/gtdsM8CVDRzr2G6
QpHfF/YaplN3mTkG4crIfJjxB5QpYTZlZocwSMdi/Yj09cesvzNHHdsmTfBvefwe
nx6jG5SGG1/5IF4ylMsxqZXsKPms7QdIVKk00Rxo/yPukxCOjO4U6P6fhx2H5YBf
cMz4LynM9HxHqqxxyMXimQ2Ij+iYP1CYxDkdc/JUVKS3oVPo6HJne6TKDAl8lNog
+j11GcDVXvfgPwyvKHLFqcJ4QkW5QPCa4dW8KRYfNpSH2zKpj7g8gMc5vtXN5BPU
R/bUkwLQ3i0JuvIcQGudRt30M1zEQJAVqFIAp2wfrCTTuZwPr7t6Q9FFCa3rO8X0
BYoyyFpC3SpAHPho5dZ+NxiRYL5LJygWY9cRHKv7NIXp+Kyeu3IZEl/q0HlRdjyc
8FTVW5MjgwdUEowWvAw2ENb+8+VCeMhYB20pVOaVKuG8PjADbO3P30GOcSCyGrVp
5UhmJrvfVv4IEnm0pdXIY34FWm96pelIdYzp5RdHuzrfLWo2646twEDGvw7nQ9FQ
EvScJEz4Zrk8DrmAsHy2bKKJxhvi/96xjuptj1GHpPdZ4C4eNPS/9/lv3Y2IL68M
4D2knnjx1nAZaEjQSvj397DszmYBtrC6VASlzeSfxZm74XZbZARs1cTRBF9AxVAS
udu9514fjIDzGjjzwlmaTH7JnshItn9QXciECByrTWWNsbUAxq/mHa8L38EzfJ5v
LBwp4rcqcXxzn8fsurY1ZTPoAOXs2TMTKSWtcd1EWS85ImtepGOjhEW+DKqnuNnP
HSzKGbAQR9x3jSnZyNpy5rer1jRO4VDpWIya85EvOOhGqtyRM+ZsZyFMvolJFJ/f
oEx+Ddmo5z3Lf1mAAkvqbP5XpshK2ORSUakPiY+iEWAzNu8gtIl3Ezu9t3ou8OYM
4WHJFAgiPOgFuYdOVLK+NSj8IYvpofcee8YdkH6+bsyQcqvEpYKoOwDjI2Uvxud3
ov80OfDP/HWZMeI7MiXD/hTS3JuW+cYjRAiovoYqnWoHXbecU4Tlq1cEbzkh2quV
OmThSdMaRVqRQg5ptq780thIT0CtLNaeIOIbY3QIZksrsaQedBZFo/AI7dOiSrYi
PIxBuTUcIYzCDrebPmeKLtQuMMdvoHfPeR3RsBjoafV+bmL1hwzXpks+YY3VnR73
wF3fk30BBKkOh2psuJwjiBc8/gdlJqE473CdDH6fPB0DGmC8nkmJGHia9Nls8QyQ
FVHOmxzW1X/Q+S2Xeuz2pzXRZ34reZW5QDyCB2qIlidZwlChBZ101SbCmv6KUjak
mjV0eD5ZKEwue47bAwlTEhT2TSy04+xJQsllOSFvIBB7LWpp8TY22HDIjZWWIWg0
RquMPxyb1m8Bu6v/t9nfREBavvSmR9xykXpp4ucs0OF5+4kaWMO3MTtWgbCJ5y65
6ClpeXjkVUJdtegYvUsDrZgQLY5EFCbHDqviKI/xZabnUX/Il/zsCQ6CJowpodK1
sFXNAiVYXltyiR3FBSBj85Ch8LE8WsdAgY8MvrZBH4r6B8cFdDh9WNdk1Fx2Iw4l
x5cmol0xJE9xg7Ee8+1CeFmUCI5l5Q4g3LNfwIG+vYK0qIrSVfSyYK4CAfjrCkLw
XHUI3XJqDgMoDCBKGA2ZnL5ZIsQlip5tEDOYwokILRprTEFLl8WuQItYdUDtRP3z
VQ4dlqKcxtPA/zamUZn7zrGHg/qhKy1m4XpSKSsZVuO/CMeZYosQXahfYmY6YqKe
spODEjg0HMql8R+U4UWzrrgS2XCrwcYawejnSXC6z+5MBdVCLXD1zqaojEdGPXzb
dwWcx6mFOamNlPbtxxo04dxe5alTMmVK7a/SKBxnLj3FAiTJ0W2KWD2mm3f8b1Nw
hUo99GGnuoOYGHqQFArzrGqPAA2mZwYwrl0ZCYZLi1w3f5o7ecpxSAvWbh7xLX/b
ePVzlM9vheRkxajm+f07tK+XlgpQ1sHrbQc5V9DXyHr5aLKKIL2O4PqzF7XqgsdE
1+IGKJgesDXNGJbIrVIIYIxo9MyUDXdZqYUWCttmvkV2ebvaFZCTVQMKGeD4+kUa
mQnV+jcR9TJPxn/KLWNZR+2IkfK9+PoacuIjXceQujwa+Z5PJTjZVZE5XvxbF8UB
ACSLEp91g0kLFVPw0niMTxAhpfbn9ZtVfVeoiGGkGgp6p6aP4pMeiczU/THvJkyZ
wC53eg/QEkjBsa4Oyz9WIkO0K6C38OGZ4S7C5Q6hf+1a41aqum2WvDOqzGsRKSRG
mnFBP0gZPVy/YIR2gV6phqOf3HIOPMxRa0GQRY9SPu30a14p29eQTkmmx2ThYpMV
VwwB5IFUvPzekDDAJLVq3y3HRXDf5jjSujh53pDky3MVXrGUW4tFiPlosMt6oIPR
J4hau2JUzQFrX3slwQjhfOgr6oKw+QXZ5Jh4d2/LgWW5EcFNNl1vZCHeGposXUd1
UdnYxUjt7l0r1GcV0AqwcAVnekWD4v0GtS0YncqY/hme6dqOIP6RDRB5pKPxfTlz
KpteZokDGchXaVhu/HkAjiB/ClX87SChNf1MQexYB0Y0O1WA+m0Qd8dHteFebf2G
SZfk/OtgG2oC9Nuh+ibrDd8Qzyy/Doo4TWZA8tMs1mbWZ013FcSNVZT1zKXxvS+v
KecE7QglrsNueSoZ5JMtR1MiEA+4H220IwRYRzBuijnKsy+QZByZaAlYK8QSvtHi
CmoSGt5lfCXLPOmeYHAalE8kZlGsOKX3zNaxQnOsg/X6nsaSCeP7ydIUYvoqSgvz
OQRjCDkh7c+3YGckiSB8qVUMMIy9TwlEaz1U/ypJByacVPC7phmbrz0qpVL9FxiN
DSY6UDUk9rCkcTOBHwobqVXYVCS//bUiSaMN3H32eBJmJt2wtgrcrYtNPCF9b1gq
tyvom2HcIVhPmuea4QGN2qeFI/eaIQV6xk/ia0MCET5ViNXDtfACaczt6+4FBhNc
O9RQDW88tXkqcBfyZigd7b7CqBS+0xKKs7aRvR9jjrjTHJcYlB+0+7z1HRI3ST05
11vMMcak8MocPB6ZpaiFeSOzRe9YPgysGJCwzz9Df58TzJx0ioIkFMs3uXYsGodn
cyZF+1IHCuAd4GUIVvGnwxOwgAemrA+vHCchCkFAp3UWpOtunwskPtVEm4XaEGAZ
ztbo+L86xAJj9L+dn6ZBzj92lBE6wq6thTdeL5Bw0NKRz/ObPKfLOvyMBsZ/MQxM
k7+qx+0ank/MIxsyM4zkS0q3472TUU+Dpmu0ArUOomf7PtykQ7gRvkwZSiVxA+Dy
+gG2WRvK1P9HjFAISbKGnkfhXHmkAPkaGvhjhRDW+p77axN1c6DhN5UNFvewVwmx
irAMa+my6d7Ex8MoYSY6qaIYC09aqi/cwWH+anGHZ02pZ4oOiTN7PbUfodsMzSVT
CqE+xxM6tjG2Mt8kXdiWSy2VIGMDdL0csdgqWcXSAnIbvsEsjW5v0h9RZOhvG5B+
rKaBVYR205hgQmeLuXqIWjb1wVVbyHSfy6cIXtC6c3ITb8BJrXg/1JyXmraoCeG9
fvfR5dE0+RBXmOkBKSlclP1YpVrS3EWyB1pfEftu9RsAZTXry0iJ8nUeCqLW5Qh0
JvpdB9Z5kWojR8j25iP2oWq7SRWCNhlYzGXPCq1SJ0ZFVNmt/k0lmItjAOgIfIZc
03wqdbEQzl2YMKah/R04tqW6Sw6h5g/12SqSs+wVqFd9KaptqRfX5FZDGv4MKwBb
2d7/bmrLWM5t2645fcVEyHl6CsTe1YSsientA2SlIxyDbx9VO8hC5RCvjOq3LSYA
amQfXXQKDtmsqGAmo3PAawH8yEwu6qomz81DnfTatD1c51m2kQPBswGQBAppIcnu
DFa5dOnQlOd+FkrPpKKttIDCBTpVaFee3FHRi7OVMi6+IqnglM4GJUDtHt+IaMT5
k154LnN3ujiSqLogZaXG5kaA/AMakso8cQrY6RA88OeWzDfurdORP+ZWEP+dkU27
ZNkDvYRyfAKmwXdIzUyZCoWQ25TZOOrNvBT2K573SVOPTsSBKHKscdvei8zVSWSJ
SyoFaDpS/VHOActo+EBuIswOlG6lxJ4hU9nPdKVQ/mQTrm8WtqP35vC/Aow332Gy
TwRU/JkGSQLFu1y7dfU9fPR1mIQDtCZ1TDzCC2L++0SQ+Ms/fHIP2fWrtbcWVJww
nN4C6HTn1VDeg7VSG+b9HWhAgpy801Uo0tASHVXPMEzfTNAEFpteWHkoQUulaRaD
SwbEzU/YG3ClHArTSmeVhXQ5YZWal8P5JKz9c84V9S/PakjJsdfBHXNwHx5UjDEB
yl3WuQHr/4BWm0YsYF2sjbs+P8NSHer+GKRXVT3F6lzgO6jvWOEN/q6lQtutIvwG
87+cq6aKFZxT9ou/uMDYigV9AHIFmuVXSWuM66YZV0QyZeFJoXzJ49h4dwWEO5f9
5gzuJf+uW8Knun1BxCc89y9sjtjWW+Y/zK0Jtx3MEvvCsmZdqEpfjAJPzAQEncd1
GyCVTfGX0BtU7f0kXiDorzucb6PhJOGYzTWkkzaXRtBpSC1HU8zfBQPIfNNMrZzO
ukrubBIBbQzwQ+xrw+mfkCp2jleu7JagMIxg7wi6hjVpUe1lzLeMlWQipj2QWlFM
ZO724Aj0lFYsqAeoSAiJ7ZYn9C2vyRycI31NPi7vq1O39xZCdIGxh2DzKZY98Aig
04e9ZxEhpl/mVnm9dqY6CEXUY0tLnh87wtkVRiL/vcHu5vhRMCcEDPBVfWjn6neM
Bivt0I8dzSLM5r0h72oMiDeHV+i1ZmD6wETBgP32u5oXWqeonBvRKRJZhAShWvWr
Ze6+NYL4/D1sLuDilE9Ju6WTsyQuaQY63aWuuMBspx+atD/wTYIulVmrr8OwT2B9
XlXgLHZNisqfm5DcygXYvSagxlmgtMzNuwkriXjUDU0pfFy8I8ILp2UyXdle8Enb
HqCUYyyBM/ndQz6tXbkmyu/GAs2v9HFIt/B9h1l9jGaH1U5jD97eD1nWj2erH/tn
FeXsSsyd95k8wu9gXzW/QPRGtBcQnAfV9jH/qh1xkhenKVauv1A+rsA3O5fiFbem
rQZUU8w1heuV/34ogZdnhBCTYacMazOAPqhXu+8n6oVZPMGOhCx3XnzEcvuV8yxI
eNCRrSnX5KG7r6zaY6K8nsFDjYFMgJ2FALCgRHUzJOZJ1KaVybWDQD5p/p6+zTFy
G1cQWrVLEe5/Xb0o99rsWA233AOVj8Qg/lgFxB5WQBOivS5m6c0svqSlj22FGICx
3RV1OCDFmPpJkYTiKzODkETTQ33Gj4lx4H01zSgvtjSr5J3sAw2DKHKMXwbq74xq
MlVuntIB5EPbL1xMfFgtK3oxwhJ5m9P1k4+rV5AhKzpjQz6DUi3P1gSTd1woZCcF
goIy0A8S50I1onTrUPaDKO6aiBAY3R0XKcE54I9GK3oM8km9KcSXxkUPZHb/FzLF
dkesRC52PSe8XFG5sijNsunDLQdkcRZV12u7EipiipHmyTfV+3GJpp4d8nSRYCOx
nRs7fc0a/8CYyu57ja4xL4RTWJOIfWuwc+WaKKdolAPP96sckPmb984cgtxCSyXS
uMWUSOWC/TP3Fu37Z/aHQzlrtS+As9fzp044aiLZdGTyUN7nduQUCHKfVQ7ujkp7
g6jOWp+DE2DGX5Z9IBbOTCWNnlcGhDIqh3YmmyppOAt5oTd+kKB9THScWZGGHUBl
cRE9y1hoTpu7Wa2sf4ZIptbwBQT5v2xHgNQqtzR1+fo1+kkFvqA7VFuG1NPXTN4Q
gO18r2l5w9DkFt1FTq40Dt6Svpr+FB0NZd8w7npXphatDGjBM0OIDKKxVDfjIa1B
SLJFySu5tQy2474snnTYI3GYRyMCmtGAflRovceiw3dV4I4WHN4teUbUshGA3LHT
qMnCEAxCRWvb/akvr4Tn4dz5PQTchum2MWLohVu/Yq89OZPH6iFEuOYPjTM+/JER
PaJZTCJWF6gmN7AV3qUMBczPdJKGTJeey2znpGDcslX/66dbF7ijLXWtAodDYESR
MnGPc5MvgnWBFTXNOsLtSyKIcROGu8FLBuU19hQZw18MFsyUVt54QvLKlicD6byu
x0kKjMcS8g5CLpxc7h6zMoaRusfJItkwht51xLcTJIRqHObdqRwkj6ehyIRvb8oH
0AG7G7RQfC3L279NSiOr5CPiY/mAdUlt7WaBb5xxgpBGMgwD9EuPKcFLzltY12Gl
cjDWqWSmPcv7Ub6vO3csL8Kx/JvcIf9tvLIE7T4EZmb5j/P2rVJPFNivJYebe0ej
O6SRXxejzBYSuMUFJEyftNjAw2fmQFM7vc0pDGyQU9CklYDHERg1NK8xDCGzcFm8
n517+U8XkLSDj3+mqywXSb0vAoOlazmGBxgt5doVAhBOyluC+o2NKKLhq0n/esvT
9ojb45H1GC5vsHJtfdA1MKgUjjEPhtsHeznI4v/C0dglepNC33tCgHVdMwiYWsCj
Lz1eszbStavr6ZAM7u8EFt22+HCe8kVbk0d/ntpqssyMGkamNbdpwYIdC20/6Be6
MchVD8Mtq/kAc95mZf0PiY3aT51dLj4ebTFnK17nMNvCcnLmMOsdiS+KAaB0JsPl
mKHLc3gZS1N0g6oHFMG3fN6y4jW2B4Ghkyyd585I6bfjxHdKIslXDR1Xf5UjFYNw
8SBzEmd9UZsDgKBaPu5c1sB9nBmec/Iaq+UYkSTlAbGoSd6nDvvenwfaUepBy3MC
ZTwa+2PFFBb4/fnyjmfjqhZ+6pYew7X6yZNXUqqzeoRNimlgc21nNAVtwkC3XlnC
jVVyaJSC0IBsT6U6d2vdNcL5Bh+AOR+kjjTPghnEIgeQkWJjvcoJVrnFIMWNrin/
YOaIt8Qj7C6T5J80jsixHpOeC4uKx4RvX9Q8yEYZyY186PECYUSMV1j59NdE0QO+
q6OGRyuFAwQqyrxn7VW1Jl56tog3S7hlmkf1efX7UQ4jr98BkwobRekfOmZQuhpn
cZP2q9kJK7wQ2AYiAfpjYs7y+Yd1sasnGFkeyjE/ULf4xmGaewUS2nGeQvj+uGoJ
qnVutLewBDDml9qCt8hd4X6ZJ/2IL/g6WWGe9Kqn2PNye3PVsoSL/vZxAXs4csHk
86HnGctlxknTjGigSa+WMOONO5yRCH52kPNzsHkD2O0m13Q4fu6F1XmyPXUltX9L
977zuyONPFMoualHdHRuVGaFhKs+dBlkabCOu+weC6F31SAQe1rlTtaYrHLJSspw
5QxuCPHkTI7V14nPBVK57V9oma98yxY5csC9DArldmBhJIyzRHofnlywkA3Ma22T
e0uq0++aTe0oCDtHilYyoguAUSnfJLlg+P/jdXLGlxmFVFouAnT7PJf8krJsLP/x
q9WMDhyW/nXdrOAeo+R/nW3UVOvT1q4/HBRLreci6arxQ5bvEbC2ZDDESDpzQG47
wLfK7py9vjksLpyQj8JLpx/2AQU/U9M0giVhoCETdZnrZ5cCGJuoWESpJd9aNeMk
eDk3xpF9m9DDWT3BrrkD8ZEB6BwIdEKAMo4qIAVW47bzfru2TkTvHh4aS0d9PMU0
iqu7iia+OhX+QYJtsraVf6xJcZs0GUAwhqhi5Ee3D6xFxHVbhbjfWC8DZ14HeEVn
X2fNpoq8IxWrOrjHWgCNtr5BLiaiCozXnzZJoZQ3xgjGsdNc9+iuPsxQiU+slcZf
NPLicCLjan2pRJ+fLSoiiv4JSnMSbnIDlDixoFNYnb69B2U+eZMH9FkpZUPB+qVU
EJJGrj9yqEnwW1k2/J8O4RlaP1tgoQBDxjb6SePPzbwvYRfHa0c3i4SuSOsw5fAC
Xp3f4iKphgqOfC7uKpU3LD2gsjver4CjzSnYziMWUeQ0MtlDlmmegbrfIpwkNFA9
9CAzhT1h2bVkjlRpdZnEm1drLyVrMDNVlMtUR4Nto6BFpj5B+HXdCXoKCwn6vZnz
iHToHwln32vERvuTSEbUqNMruG9JCfD1z2t+p5/Yjd+5nZgYo+m3j/1lo7ybrCNr
ZNJt2hhIatTQ/knZ4RejPDwoV3LpmVq8C5RA25d+TrQ0Jx9ldMhvq7WEiWC/eZ5x
RmQHmBQHVK+trfjGcN1u7lY/WznjbUh6pzUYkz3v5h2Weg0ybCSh96XagmcsbaWa
PQP+ba5G7WfOBBvsEa2xqMHIem+QWev3gD7YRcLd7Lav8z9rgWOUnh4+0tjdfcna
GQ5H8b8JOKXhtyRQuXxTYwLDVuK89x24TxFG3aZe1qVWN2qWQNmLuya3ddZRj3yf
xo7F0sPqWCS3HC74u5+rkSt4Y1+6T9wbtoLGLSjG8IOvFFiI7bTnltGLqfzqbYj9
Rbb7BnXZciS19YIt6n4ko5fdZlqPhZqinlkHGUiz9rgx+0VTZm3myVxHZkGqJ9V/
oyYT0boSxcu1OGI02+BcT5nB7mi1FvWxxNheCf+DKZ9BtI4eI5R9LmAQhqoqrYxm
JSblUYmVKPfNA1dGuPLN7Z+oK/PXnUnjiEe6cOnE719+v2izQEDPP17lgpxt2KhI
fzxt2Qdgzm8dYkdcsgZsY9wyDDhfAZky9gjZ5AuI05mMVkEdR8oa00m7duMJEuDS
Pu+whR+xhmNvp6LKwedErJmqVwDRKrWqOAUy1wfBzY1ZKOSjOTINyxQSbrHmFqIV
lvryof2bUBGfniOcphVwpNmZUPGCpQ/mIhQ5onxDcLZvdl0x44IC8/heps14BqdA
dDoiH2W2VVKJJ56mRPQ4T+q/nZPXpucHtlaaEQoOOhgW/jFZ/8qDWkeZPS+4+RDD
2UHazslFMcvDwO0WnN3N3rTQ4Vidvl8onLoKiLKmXglVPUowIgnGtKaqHB6eVS/T
179zlP7jiRz2NtXD8N8PTsCe91IWNzqmLUctBHaJEXRW8JucoVU+ZHbVKMVFavyx
iCcFry6T5g8zHFENM4j2UecmI7N5kaW7vDVf7CnlzINlCUaGcdzCHEir1/u4ugNd
WS8BB9YHno3rsBrhbQCXuOG1MiW2z+sJlNk7+BnWKxtYg43FKkGZR6Vr+YcokSoS
NMbbOlpY07XGbhyEYalFjNep4q/CYR3tlIRiN4RaCRrDeGugeJFlhX198YgXjGr3
jvs4tcZ8+bVd3I8Da+pm8kHWpFPn0SOW0LY0l+aBJ9Ig/hagsxZR/pgE6j/Wz3eb
VsaJxh0cUbkoNmkD90N2G8dE3gAaZz1ybenLUaCQZ9joCYxkgcU5ilCdXof14epi
0V4NSJGEgK2bP63tF0Bje+28d+hz+e1dyd2K9tuLBU1ex9WF5vH0FYrkkt+TSQLa
9KJAX8W+VnQAs3pem0rcG8xiKore9VYhvaNGim2bBWqSir2HeZACLtewAutktbwU
2lSCb5nd7LUTHajmms3R+LiCfup/xGdvMhenfDT/kbMoROMCdQmYhutNEjO/b/RR
Zbhe/qGnqTycpXY2ivJcMKsQY0QQJ2n2FNoorONJhB9RnpV0cN3z0t7Df2CmCEMc
VWRMfzvZqk44aA4wFXU0KfQK2K1nFO3NlipiWFuiDmSf7UkFjcF67dqLlYrR4E/k
SKY7N4BO74AT7zLdo9uCQ8Hyk2+ivXibH2kZIrtMQol2vcgc5ribCMWvedeCbkLf
2E3AEzCvAwltqKkiNMXEpDXEkWFj7N1qnv4fG5MLJguVIy4CK//IXk2AWeP/Sc8u
UlE3RZcI6QLWOxS6TqwQMpnRDce6L3CF22FrrmMa6S8Rzbk4AgL1UfYdPXp5YDaq
T1LGCMJCTo1jAym2rAhyYvX3uH/gUrZO19o3Iz6biI+hVJeDoNP/EkNTuyvXevXl
zDrFPpy9o88SnPUYL/xwNhQy4VW+rSm7gtofjjmGmdYFh5k6txfKwdIi1R5SpLx4
9itDXTx1w/MzTZvwyDpsjBMo3Qusfyb7RS+TzUuN1cF+ihNaVAfGuI4nSv3N2Cpu
YyTTXZ6uHwYty/M1D2CeJ1SydQwx1z3ocueTsaBgUXZ48IUfBXklXkfgMaAReuWq
V6kR3mopIy9n8/q9y8/b3OQ/gsotHmYd/hpmV4j8xOw6F+j7uIG0uB7r2uut2P2B
1RZBwY0iJNVTUZtTtvoVNZEFkG8br4oX9aOS+z/3+eSV/9jTvXeNzB8lTr0/sfes
cWUFVQvPTJ5iMxePkmR9GyB439pv/CHOsx2iugFFsei/H9pG4cgF5dmCojzXGnWf
ceY8N9uPOI+ct6Qbg2PpZMMn2EVpc10FwR6kMbZQPtihk0lu8g5+PzdBy1t2OkYA
YHBjQrIcs5PT/pjGa69hxxlp67VVkyjR5K95iqQohyC9QK5YRj6ZJ1DoKREo2vpq
2/zx7T3EJab/eS1oukSlxL6VGe9hl8h8LJ+rrSHeFoLeAzqShmlQKBNzIqC8Gwfy
t3oVbp9lEoBkZvARhYWXW6AdPH+r2NhisX1m7gStgrCYNbMepWns/LfOCTDMSzVN
IZoL9GnDKKqQnMbccxD9jdCBVYhJYaj2473KbHLUS0OUL+uC147+aVE9ghi70Rse
gapTrMisb42KEXrfqMjUfLk+IUecEkwdE/Iom8kt9gT+uyj8KGteHR6zCNI8GKwo
Ho49W811zJgX+DBHOobzwYbdIlq17+o7x67rT4LbqC1Lft9k9B2NAs6nuQK7LHrH
/N0CCTpWrI3iq77rPTrzaVrPV8VII2wxrvdYW+ByD4Q2SNZ8uzB66salRMMOjBNB
J3F2yvmVZTWNFI7zhSeWgb9UgIHL7NrMHr7dTNSvZt0+YTIuH1zM5zumh1hWbQFv
zYKumT2+9svVDUvnrGiRtUeMpxciDjiVTG01IHO7tg7SpVz44HGhfydTZ+zBNtFk
VgSWa77fJS0mGUTqEW54h2LtpLwquos9csejtcT255GcuD9aUo5mWGBu5cwW1I+s
F4Db73a5vQuMIwq1tbenM955naQPEptkSQ/23Z6ggxZM3D5/8ckBMdKh/OCeA7+y
RjHmO4FNhuoLzC4mGMyOGSLMb8ESnC+Uf5mJUnrQYpihLIA7l3BcpoA2CMLiI8dK
/yMKK/iJeUG2Bpwuzbv3dXDnsTCLY69ZUCJ3iYgDUYDNBotwPg1AWD+2HZJCLfu4
h1pjno1R9L6tViEnLJadEOFfD8Vx0pTK1PW+6+U6lutOI7FvTaROQGQUxliUQW/x
kIh0lfp4jC5+0Ut39PqBbB577k4ZXNVz2gA8Zh0t7K4t8QRLw3UemaxvBIt554Zs
qnm9UGR6Bu2oY7nN5LiMSjcsSNfCjutbqvzMkog/1kTTOtXpSMLi6omQms3rResV
O2Nn+BO6kS7f9szYzcmKykqa22Vs5XFlppbkzMYTybNJrGX+rLJBsxNnME8ubYrE
KB8kufXvUE9BaVjjYz1+S6hafAezuKZ8VPQ9E5JXQcAh6snbn3z0I7DliOnXf0Ow
sPwhXA7r02ZjpwEL86XfrRkzC3FAhN9CgItx8aRQT/kZXLtYD6aE+e6x2MiYUy/3
8D0HD0zPz7g7L24JX2NTGFzKXojmvK4Gj9q796qaYqNpm6wkvtNI0jRC+Nyd4BTx
6pv4U4w+fNtPLBEyGCdqhoeLnoGp2KZjVUE/L5UsUXnQu+fxEGlK8c05L0CrTpHW
r7t7YA2dNxN/47nfb0yV4u7Agjb90AH7OlYxKwXHdjXgvFXpmN4+38T4Z7DiwXSi
4iEvJ6DI6LBJOV+2tUrIwHc2Y+h4nYa7XNGOsjn56NOX2M5ZLs5eix/v6TuxQ5k+
6iwWaiRFvssaiTltXj147Zi/tSM/q2kPHX15YdxaTKBbQbnBHrjXBTWvmbbjWjvR
XBdEMtuSHuYse6X5JOSnUmOGryl2oIONd4cPqKgoJMZAdnQyJY1VgMpTowL9JeMY
xELIuy6vozN/b8np1Bn65PT7dLWomC8HY9ABS6Bss65jwsFhXFAUzgki3CeRDYjq
ZF2Xftl6SbpTp9IoiWfRmi7JbGFkKfNAFmHr91sg3qEp16bZy9D+ZHpfpx8iBkp7
3996jelYINC/QtgCGuqOHwsZsTV3BlmPiOtTcf48CXKablvH5XakyLtrmVAewoVG
OxQVDnkjeZxr+t4qzydXbBEocgZt+9N/ZbRqFMprJCFeEfHc4SvynU/TfwBoqk7a
x7B6ejBEftC1gIZOdEOuZPVGM0sPrpt3rOegNJZuDXhMZp1apItfEF/TJ46h8DQ1
e2pka9pPmPO2xCM3SdC+VYvZw678ZZgDZzCGUxG5jpboT2ybaVRaoAl/ZxCfTdQR
QTXpEn/NKphMnGG59sAI3E967dCoSjbQbE+y2uduJIFDdz2MmM1RV0+Jk4AusphF
u2cugTU8HpuhuYYzWj4Q7j32B5U5rwlNpQ9a8Z8oYfWw/0t5vER10OL1/jGGM7BX
P7vmHhZ1dPE1c+asNdkdkAwj7ZpubpzxOExdzM742NH9KdcNzyUP0azpuM3wWKIK
QJF7XzEOaGRZuDtOshVN7KInEwAMSOD8Hm/KWpNnGl2jtgQY0OzrovG2AAotcHMl
XKGt6gPdcs3GbTc3si43Or+MWv4G49zo49U8UPJab1nz+Yd6biY3ELT+BRjb7QT8
Y9RGYuVFzsqU3hlmGADnm4R2TUtGR2kqkARuQXzAW68pjd/pxoGOGQTWSDZpQOge
82gQ3NjAKs4mdIGbPjZGCSiEOIVfTcDvdBYYDFLbUPPrX5QJZJ8z0Mnn5rU/XVhK
8FG48hbBKe9nyawRX3+NJSxhxKLd4+8oMscCT5+AJJkLHqh15LI+u1vjXBL2Rkot
3jnxT4fr1gN93wCa4V0fn7nVsUwLdSFlR29Qe7aXfCUJj9ND2e6QF6DMehaEordY
XEW3uJGm5cVSuB94w4mLWPn1BcjHK8823JZV0RJXe2u/EOCVQUdTqymfZNEQTfZC
lln6T2F1Y9VuNZ9U4av46O5naXXTnH+A1YocLVlWbLcmmTcrqp9pDDGmsxmZEdjQ
P2sx9HLauW0zLq/PpkcupEv5WbqVKfmpUTAtPpdvxtSCkulHTRisNvu4ql1Q+RkI
te9JdSF8ln56z+u6ZgR/AQuMjVQoByqjD0u/K38xeSH0V5fXwlUbeTYm2QZqPan4
SfH264Nvq95l27UIauwrsWKzILlCCHuMq2k7DvvOMBGOo8rBiv63JQ3RH6EcQcst
FWZwnYhARe//IVqK0PxbAQ9lXRp+aVLzIybxSBo3CPZmZWporgFUgtt2r7CnZGAF
2y6gwLW05dHba0X63oAN+dxcPSA1UaGSDmBex0lZ0vzxtB77MhWcNrZxZGOd+qUS
7O1FDFz0/jBXyrKnUtkCO6IC/WvT94sw/IhR7ZY7q8Sd72NAP90XVChJofzjaBlY
z4gQr/jA4Ki7VzaHl7PuXl5EBfX5bj6w3rCinrja2Y0BxZvsl9o57k1m/fCOxOtG
/6hb3hgYHfFOWjTmkotdkemsTjpVCI7sZ9InG50zXLKztvcJU7fFw1BJRKK3vVfI
PIy/ZbhVPgH2RdznwNOfppLddG2InpmIxlD6p0V3d3goet0HBcCjve9ScKIWzKLb
Y8iQva1wyJgzl+4MBwL7l2+uCj4GiWj6L+vFZrvM9T9MJLYpQtsSzDDmaQ+rXDgo
4CUGEH/vB2qe232gaXEGv0xMJQGlKPfN2hIyphEc+lxh7/5hO4rD4+l/TXuHzFck
jSvdoUZLj759PQ8TdfDSuffTRXxF3+KagY9/M9Cmwkf6D0g4SLelttimxHaYiJr1
0w+AMbQjGKi6ms5HgqRaz+kBIfdbFn8qHg9cVY9nqodK3OpgMlaUGLbfv+f4q40I
PizZL1/Y265Dln6GiZdIjid9kQttNpEI4FEfiBorRtIUvOLlHEhzC/lbi6LxMcsg
6/L3c6j9BOpXbBQ1d9vzDRp5wBUUC8gMTfjJt24kSUp++iQfKSMEQAoBoTtdAkfx
GIbGMUOnYGWFYJWdZ/0L72LBTNpWneeQ4cesp8xzIAv6469RhSR4qAzuNVZjAZOb
s2S3vmmnXkdt2WzBluz2z5q77TBX1Oa4VXA0kN2FPcGjdIaLokhUyzY8bBuaOZLH
nCPBaG6mCaMOGkNrPcUVGD8X6kchBa/PdDllQOGSUPIaFBfyS+qNzSb0PA0kX4WO
KI7RyRj5/eMI4wsG/xZU+xWmHUMB8/ZC6BIN34SYx0yCp9Nd56T3/XfX8pbunjUM
h9hK8ghSKRFHBBqIWKAFK9k+1J5lY8WrqX6T77gw1zLhzNb0W7lO4OkwNHSi/kPy
DmfNaw73VDDwukJVBTwiVm8HGO+sfArSVSKOFFyLeuUYFYj3Ph6By/8sY3U/6dWZ
+AnSa8xin7jGD9fP6sfnu0gkAZbwuHVj8NRj5YZ4+/v6Qk5OkW/YFtO2QaMJRtcp
on5paANfwLRuU6AD3H1GIDSV6o/oTIuT/y8Fld1I7bDlweqp1F/MlraaReL6rm7V
VwsrtwqDKEZXTwCb+MYqdycrv6POv+VLSAw0A2LLXwzZLgHBTAGHmy9yzoGLHATc
IYyswRZxDMU5H9Utlm/jTcsHhlfCYUZakgBS9zj2SDlFGu5qOZyYwxZyJtRssZ+c
DP9xrL/7XYiNPejlYT13STe0odOYn+k7aZdXPBISMR45dujzxGPW/GakOrNAm6sZ
gAaRkN8MTcPmHQEUDr0bsa5ZP7MOEAW7r6OMP8brbqHTJ8RSAByo9oZehmW8JwrI
9Ol+QynkSwT3IR9agaf/UsLhJSkUhmKfiJXMJ4ozu7NM2CqCem2DgSebRwSiZ6Iv
NApZFWBtj+YiL3I8JO51IogmPYbrYviexCnrDMXz5rO7IMd1NXyglGOYyARKU6n2
IyisSDC90TZTVGn2jyCa8FZj5T468W3uSDp+SSTqmnBKLQJMIPOp0QSv3e5RKR1E
dPFY9rhm3B2kzFeyJrinDajhpHZnmoHQ2LQ9mMom4Tbpd5I3RTGXE8KpCs8DeaeH
6c6pW+3SS9ElROIM1fNPzrw72yXTscV2z5nmt1oY/8P1PnVaMOnYFWRpqlKb4ZaQ
91yOcsPBhcrLMGf5nW1k4RrH+lCFUh7gMsG3Z4UaeLIhJjhT9/+KJf2z1rU5NAlj
m0+UoJWJwtaCE3hA2LjkaLrsHIDj3fqV8ESxrDzULIMCqvOxunbUwmg7wzc8O6sH
bQIERZyeGHBy29PhBKbHBxabeb4E4Ov9ecoAKvZxCC/aKV/5fqYZRch5PFFq/+id
685vk4ArHY0WnWuDQSvgc5+NBtQscAKNk36eFxUVqcdoYyjlb45+IK5IBmftIwsU
UKL2tR0DtxWlSL1f8WH04NJNJKO1tyY1MhQWIt3MdPwTrLNwt3GO2Ln3NxziWSe2
IkctHRXcF5k1kV2Z2h45YhxJA3jOXreRjaGa1fMjK/F9mSVNFp6ctw2nWSYukB1Y
IgG2uN/QWIHbpq5sjiZx3PfBIOpr6nUNb7tpSZWxm6gFht/pYPsCzQjntld4WQQe
6E8HFOdRoybEZy6d0/5q8VDZdTS7a4YNQVxob2XureD9NFmIfuy8f9ZKD2Hkulkn
K6DNSH5ksp+oTmflCrr38k9ep9cMcmdKPtEYxesp4XyLxmeOCHOc3IMO9P6M/Lfv
d0SB1kheOnli5b1CwK6lGOaUf4y7oSV7uBEDSeUWEdDZYOKRJia9hx6n6o5Vhle9
xoB75T7U51CwjRgqmbdfGsj5otp2k7t5i30l8zj1wVrRnE9xfvXjt8805WWTRGK4
HK7JO1btHAHkgclrJi3dZjE1PWJzTV1rAYJLCfOP3wqVhg9rtZ/FDfLkDLbJZGHI
tEJW5O6Xf2O40J4+WUiWzIMRG/T/jaHgQDMdoOvpguWevG+PX+o7KCCibFsu5pW1
uUag9p5bb0jsnB1nkDmvSOKrRZ34t36t8TNFvCuSk4io0INuyte+v8D6QnpowCoW
IegM2CB5dYivV50VKZqPa87ESYBkJPtHTBq+MwhPmzCswY6ycyhVulNTwHYP4kt2
+BiTVhCYK+Vfa+WTsSDeAppvOBsQ2J8WMxzMjPBb1Rob2ws/bP9hC6yDT5egK2+i
U2pCdUFdzPNETohNmer31f4kj71SyvRBM2Kdil4zJhsdcstu313lMIrKv7LJU8iO
B/OjUMvdevantJjVbVG12PHvTtEOCpeiryFEys2o9W7xCD68L/4nJ9cc7MNj3S4h
Vq1t6F6P6N0ooeiILc0mDlVRQu32iwxtOp6hEEXypc0VOhlMXIhM6t+gVbYynxFX
RcpaPUFPmuOSgdHVpnJHz2Xe2Cf4LUVFdy3Bqy4lMC4Puzy2fUGnwoBqlxf39Xj0
rxElGnSWJ/SXfqP+E68Jt2AQxT6wYI1dn315bahO44u4a27YfwL0Qi7EXiT2pAEi
PGuV7+g4W2Zk3GF5OaD+pwuJmS9+0Li5j6Fw7dQj0yWTedSKVVsK708bKMALaxVP
Da8XLFMAv6QME4i5VOOi9Ijbh99tpyoga4vuCLZr8sHavvGI+sWNv20r2a773EuL
9eLsQdV1GIMxZNz/YHB8wn0uKs80whma27pfEVXJssCztRzS8fVorWuJxQCxTBEs
bJtAfIurN+J3BXEcfooXKfDGhdofNkuC8/59KuiW0kNUoiJh9AF2zchUwN/fiuhn
vXQyLx3tw1vXTzPZp0m51xLALIZu5iEKUskjFzL/J6bw5G4RFl8kd/4SYFDCIouk
49dcorzAYCGNs8DMYkSrZGmNF3WoKIZ/jgQaum4z3M6n505Lxjawex50J79zyVQ/
BWipNiHeH3b22dnxQUpjikNDCRq8yVaXdU4ilrLZmvzG6Wu0dVUvwyckAxzR0n9i
YkY9KP/tBNh9ij8aiCmOJYnT/ilVUaYXtiH9u4EWLec73OSASBQDMdLH+LlbowjE
oRFRrCVD8A/9sIxBPeoWFj+Y3hzWfMT0I/U9LX0nJqEsFfRPy5MOAdKuGBItpqZf
pyZCCCPve0kAY75Tgt3QlIzLQC0BikU+5G6bSoOe9VsJ4rvVnXPkkNDbcBJGSpOd
99nnMXOb+A2yhG+Yfc32L78TOxrdN0mjR90TLwhT48ink9ECCswD8qZQJ/RDwulJ
yXM3X2l2Rq8Z8hkuhJfWlKbMA5VaUC4mIwsx1oLwM5Kz2618GNmJgIQNp+Sv2I32
7XCr8+hUI3uaZozwzxAbu+HZaeghYwuRor/p2VDYSFvUCm5E5SykDH2/I59VM67X
LqvnMssoQn6calhWtnl5N0MIQfX8RM2Zj+Dc9bOh9dPQ+h5fssFZvsQ3LkGUOpKl
8bhbuEv3TslEGNqexoSv+FWPobmG8lys1S9n/EIRZeojLR82dss5ky8MUh1Ztwes
wVzE1RdRbmFEa11M0adhG0U0/7IG55EuypQgQyh08blb5YS9Iw2tW55yQhhVpl2Q
YTds7/L9OxQ5ezwT+wzzIm5hbPcwLtx4uTBDm93QYkH4ktchVNvnYqUKKno5VAD1
QvoVzlSrnEh/bk7hOF9ms/mofB4lsk69sW/Sf7Jxl7+krgSPtnfOx65bMuu9YtKa
EOAcAikOegg47cRiH/7BWxe34sdnNhiImqKHJe+xO/OX9hTFTt5M23OUF8peK1e5
YE8mK6FWo4cQmqvjLRe97JKP51rPlP6BgsRUKR68zB3flwh6cUm+osUyIXaR+47J
X6jIZdO3dB0nLwZkYO45qFTIZVdG6OtZbS7fccCU9t1By1NIdCuAbyg/3spUiEl1
LKwr+FoXqzNn3p+3kqTpqmADaop2vYjbpOZw7XpY2R7yipaq/MTBI7xdujYK4qcA
09rQEYpZJLvoUkt+LXjh8nTWwEPSaa61T1psxluKAAdXX7KANpNIKKWj10hbQJhU
R35lcVCb0paat4piW9e+1fqa8b44RpoySznFkcYfwA3WBamWWpvLUHOUFAoAeSgA
JxpxLQZdS8ZSXqSwz/wAiJ8Dmh4KXfiWGLaF6tAh5yVvOkp+cLpe0N9lJBmS7uoj
BgAmKlnCNcqMj5hMFJ80HR+l+Y5SWc6CcYWHOy2yEq37AwBiZKonmvZF/AohD6b5
Z85+4twrWqnKFmkycsFwSWCMlP2ktKAwtHtCquBkmqGgO1htdJtmEt6aFGlvGhDH
B5MDa5M8Ksn2kejeTbpuIUIdskwLbmeLo2bMh5vMCzrTAN5f91JTBKkGPdBmGBWN
s8x2t19gYGSv3u6RFmSCA/rS/L0/PcpVOjmaNHl+6LtOyCaGu6IDQODonGuGXgNg
/2FVLWTqNOFiRW9jotQ6tsrLNo/jRKeZDilfQxcvKZwypWF9C3D8kDZu65gSjeSs
iV7fQjF4+sK67n5097F7d9wyv/tsMiZTt70l3KF63J82vIdXaFDKaju35yq2cwGD
W9RtAL8DOiHNx1/RbmWfNYSdMVqngZV03LzXKY5YCTwGE6s6+QFWjqmaH72uout4
9AcVfjxz27MAvFUfTAUSN3hyhfl9syDYYVyn2LgylcsrG61+5D0BT/amQGBcZYk4
xN0xFXgb2/pcGnT9O1ATHSMdtJFZzzQvHjLKorMstsAYh0YWl7+LfMtHRQHCbcnR
pC0qG99di/pRzPvZBUnvs3B/k1rAViZQMN0KWFBnudu7RRwWSlzLEfVosiDAlg5J
9ABh0NXjIiVNpsO7B8FrqPEFGjbrcpROJY2u6guIHDzkhFeElBccGxLVeWNHTHS+
KvkyE7DyYsuzUugs9n4MUQd+k8+axBJ8mL5khIQZWBaof6VI07ah2uslUqB+nulz
MV5T8a1MqwqzjVqWugmURjkDHlURlJ5VMRwbRJ4wlWaLYyxVSzvQe/3anEWwk5s/
u9yAXRy3XH5WWZRtj7y84XegNp40+Ecuuyvof9o/8jFIxgf7OBS5Wf3xkWkwkJB+
efprbjQ4u8V2YjgGwmhenPDs6m5Ch0+IS1EDnV02O5MdiDtKWqbjlOHMp9K7WWaj
cAFTPT9g1yOX1RQt0zr10sKZqLSew/a1dXAlulUFZSOiDibAeTRS1v30CePoevV9
TBCdxB/vAn6rqb2pqP0UjMUYGz6u6vnnu8YO7DD592IZkkhBOsbuOyHM2dnz9QkQ
4Glk/634V0W/AFg2gOYbRfQVN1oFOeMKv7dvW59nX7PzcS5ec1YDQ0j/8+tKdTKY
FP8Wugs2A8amsqK6GM4XxQIPXJc47DrsMcD7aGBFfbs/nDuA1LnMhVfwA2qhRKWu
0krqMWPiW/L0hMOIpRGfaUN8/xlQH/e1TAQblWUkQthHHHJk1xHkIRMPUrKr75rt
WdxpFxc5g3LSD0r3UuDTZf0MP3Mcm4buwGtrutMHkx/G5ZYAc+WU7JNmso9LR1iu
zauGSGSoUKl4I3GDGHS/zTwJiP2jxsJK3iT8p9Cvvo6P8z5liQ7w1g6/5UwUYnO2
7mXQDvkWKjGa2P72p+Ee+0z4Pu65uk1ghJPzRDmkGskT96TRim6UMZcPIVy7d3Dr
3MI0Cjr1uEDRMeGLSbZ3+w6wgbOVe9RehNym6RTfOb4ZEoYuGtLLk8v3r3lwjGkU
1iyM5CB6FqieIvvKAdjUajxk0siayKiQDyiEcewsgNXYI6XFLYicK0vfRpfL6bdm
WH/PinA3O++XlZ9et7zX6heBazAo3rtLCjk/M+vxcYiXbhQd+DlP6t7uFEdvukXV
0FQe2z+VVnOMtDcdmR3k7g2IoeCRq6JasWTZxVAsOwy5NWKBpEcIjELbxt6PSgD9
0cfDeV/FYTM7luo7/G8JXNGUJu9aFcHAB1M5Mgv8kLD62DTxH76320ga3htVqcEO
zUnKd6/Vqt3stCfO5KkrllbJ4xOhA33vU9NmWr1PXgatN+jzlxxgUNTIg2+w+ETI
aHbRrw9liwoat/IhmqaQNLkvoiNlOuiUSyidK7ZtounHjJGHxyNvwXXPblhBsGJL
m1shdh6SsNHTYOT5xqFoK8cX5YQsQyGcbpzuHM+OL8csazHNkfp+OnwfGieyeC40
WK788IdEuFtNiIvhrUQ+NYcZCkz1OXuPr5cP6HsLoNJohwbq3Fnqps8inJvhj1+U
vIrAQlv9lOmsTStYpHBuOd+E3DNcA4tR7bJZlB/WIMyi85i71a30zt6CN+YuTPu0
UU9eMM99ndA7gMwgFHpocxcl9liqjWN7PyF6yw5ySoDdplXE+VAd6ZzwXO3i36gN
47w3Y29Y6fDA2fg7WO4ogkcxrNQi4TZ0TN4idoiB4TKfAzVz0t0qWXEwlRl7o7F5
XDUq7rgtIVaHZXzKL6SiOoGedGiQ4NI8P0mJQmhOp+1I+P7zVMbATz56lzd4q1/F
ykIVHAYUo0KP9NNM4iAQzz0+I0BoNSMnJWkuEhlWpmKtpZ96eweVTYDDqmKDlzpG
f71au8gK5HXsobsALbGorQmliaM9clJ4u7O1xNCLu+3zlVceA496K3Sgc/8eJ8il
87Wa5V0RZ0dtana2j9bLRj4F9ivGXtcvMyw6sa/MnpvsaDO2zimlDtD2qciOpPiV
HJW/X/E5BQtiahBm1G/D5fTSeYVH6RLSgP3l/rP5b/zCBx/8266QxkI4dM9n1OWG
Bs6MYW6S92zSYPnlZsDZB5BN6ng5mP+/tOqWfD+88ibeqQpo06/LbIL3/qbetAz8
d5PaYiiwnpNjhyPxSr6gA4RBzDU9CYnBfXvn6fN+DYpV+IbRvbA5hJtiu7BMPmVo
7F5klY6/WLXte18i8mGKSgX8flTYY3AXpfXb2ER0dS1+Ix9Vwv5L16PLSxYPEKmz
iLzms1eTxpXfQ3rXm8C7vFA9UBh0Wo68sb1qTl0kZZbOeNUbEm7beKbomNZd/lzk
bYYzARrSEiqpSBYUyLnAH7pPzWIXdVfFJafsZo6ovdMcPdteuMxm5oavApoDikr1
YgW0oegIp4bi3VlBGk90pARUe3QHhdIMVqlnfjR9J3+pE9gwOcfh+HMVe2M//PC/
WWSEqontMABouwH1Y4Y5Edi3xktgZL44ZvTUdHVUqmUGFeIvgUZ7jh3nmm9zfON1
ipzmTCRmDmH831o4IfcIZYTCLcaA2QDFQi56cdInQPwAYestpvev0xJj1zUEMJa0
Hg0F7d1H/TfHTTAQ62VJgveswaJ3UEjYDnwAJGFtsUy+yDxjRJ1fbr24T5D/V75u
lUroU5BOQRqrz9PwAU0CozlV5eHpNrGY7fFsSt5T9hHLetq/zfb3FQDQhsQeJs7h
ZBC/UD5PIbCDrXjY5y0vpnIq8zxxYKEitKVEqM6yr8a6VI5/fh7kl1AQc0ITf5GY
8q9br3DhDpFRTbIVJEuoAwIjXgG/2I6/Av05Vf3HD1s8zPH7PA/29tHwdY062Yog
N2pmsvhKb9bEUviQvxxZQ32FEkNUD29re9TmBORgPblRW4uGl4crvljHt4ODCTDv
w/Dr3cxto4mturdowDbGo+5jKj53D3a5c3WOnI03JQkqwAFM3CGzZpt+ZJI6Tsh3
BfzlPqyqqYkFpDqxxHgpRVwbUmX1SiNvi5sT9Ur8Eb1d8HNr7rW+SgKMBU6ya/kM
iOqyLxPHqVGjYf2vBWC4XQRaFxltYokyTYIheMiXMctqy+Seew8uOo+mjSQHgA30
ZkBpgp3snJxEl8nUSGpmqzTRPKo0QuWSVGzXrvJ22p/ghbdE6GD61M7fYTYbXxs7
H5oNG3xmbK/+vnCz/kh29LOXX7GvxOBCRikDq8lENOVtQiI1DBtZrPCVxWp0sPl/
nU/3K4cgPjHzAG1d7Rda/zWSKPMJMPEHTBnS/Uob0ZkHxX2Zty+c+1SkPF+reqGf
EJEhabAmiRtH4Mnwcop35SwWKa/wGsDCfBUuwg1paeOk0JcKClUFW0yzaQqXOGV4
DzNqg2zh6GWc51kfvbqH4ypWSiCCFSSeq0MDYQzeipcXKmzhMpg5jEeScmEKuCQH
K9/Azch1w8M+V95dSjvmISLk7mswpbSuypyvyGr2dQU0cIi+r7drVnVpUK7Aas4C
7tTxN0icrMtQLvH9SOj5pVt5gS0+t1Z1S75AnomOVvED0gdsnogonU5BgpeqRM90
IC5nCVHYPO+h9k4H9mFEbPVaF6fGNssoDbZIRzjGCUOXeZ6JrtR2Zy/3miISts2q
xPTyg3JpNvRJ4Y9ILrdt+h87wZThMMfRhTHPnUOtlttqBrgtzbNumliTtuv0B8go
r9OVYeuk0YZ4eB8Yn3DrnMYSXjIGYtFtv/Et9mwSFp0R7BPYFg/6YsRHv/DiYigr
/sypiekqEWeoQsmKYCO7MtSgGIqKEL+sV6iluhtlvO2Sb0TSiXRCrvsGXequfvGf
+Z53sN9UtaH17W2PzNjH5fhVYuABss9Mo5zL8xxmZDYt5lT6LhFT1OUiQV7NsPuU
ZWPOPFdBnTzd8uwzdVQhHlWIunSkv0KQjBI2EwZRbVPu5rdmm7baQ1lvRAlCKce4
h6HTDw9KuEDpowO154gGP7/dZPi2COFDNOZw8+/Iw6/bHxofa78kIBeltPZR/yi+
8OaIptvxTcj5fnPC6oIY+a0KQCoOjPxFK/GUpIR6p0wWmYBpBXlMcXO3E/fzUApv
cwHDi8ByYXQ8Nnnn4E8eOdsbmmHPT9MHmrPufF9s4GDoWoBGCq8N5D8Vkc9B7CCg
EWj4SH7hnwbNrHrL9g1iJ215ba0+DwSxYRej8Th/NIHO2DyDx0KF8oPpH1YODyZZ
pyd53dwuEAv19DQngRL9j1ycJSOHK+c3rkFNlUaVNGSHKIRdNDXkTvRg1PmZnPSA
sCTSDwad7DH8lyRbGn5ndwXiH1uvRKhuqmkZEgrQr/5avNFzA1i8l6i+F5lnWGRc
8kHxKM7wj0/ct6Wl1wNMTQyGRxKxU3JeseSf6OGNc+gjK8Ozk5hfrwTK247mPXrZ
6W+GNp1C6NJutt9gidw6cSJaA8Wu/jhoKH4pZ/7Au5KXSV8g2l0fQQPv7LF/bcAW
d0Lsy0CyhRJ0ZeTK0fOTDvHVNUwfMI1NiCPBvXERYGscpBk1QH2NFu726z2iCekl
xYWo4QENROc3TI2G9e8NfaBxVjKnU082E3h/fsUalNXrVIEqTa1feyOpIg6g5+JZ
85WNkOIU96sA5XzTeANJtl4i6tDwOutnz900/QWIADCcGr/YiJH5ide8RN42Pxud
WfKNm438HRCDIQNvz4Q2D1sp3RPZuKzzOZkAq194rfkTmwn1paz5NY9Mcz1nWYKm
fzTCELA7jTGdOPEZkw4vTay8hJqqRprm+G4q1g7BmeElBJzHUS1eeQle9AWukUio
GwbiqYLHTupVtIQemKl4Z6nEL6LsoONwiGpW3z/qrmS0cuy+xOx2wFxF72H2zt30
AuIHY5ETjMK2sLv027zysz9bWoH82EPzpB9WRToLII7RKx5rKgPdlck998XF3qt7
fKY8iCZTOOQ1Tc+ITZEZQY/KxSIkrSg3eSMyIqvpJBMh5+bdwfBdmIO/KI45isWt
/9hc//7NAh84m9BPYLXSHG9ov3OaCF9rbHFGw2RhWI6mnoq19Ytggtg69v9DqbJF
B+vaf8ClSNXsmszMO0wuMJEqkk3NUziokX2YEv/pz84zSshpZdgP91bm4rTjtJO5
AD+Nc5Gg3eHMm5SsyT+AxxuSGJ51GHn/3v8H5SOCAsTwhIMDSZpPGr/W/Wkx+iJF
B8cvpxBg++X8YAb4iI93iODfEC0gjKzZ1SWtwHP/9W1DQisPmP9ju59e8ZssmarC
BwOY37uYmFn5PLIBbaKWRt9p5ouvaPHiZn9jtoUNxd+JMLKfov0CsvAIn1Royfup
LaIP15sIFSVClzLV2qejOOMHXaaeT6sgxc/HsVqL6AGC62LP+UjMGU/u342/+3a8
FERShWt/9DApqIdMEQQyv9DWSA28BT2pbfYGdmmtTnGLTEFAEQbxL574VxnZRvgs
W8pzAjqYWRU9/rDvw81kWo9hZMnacCUm/AmyxEefqR6Ht2WfnQ9FIAiVKtb8TlEa
X7/dLdTfIJyXX6ztr+vFHJdnvkU48r+1IHXYAXc6UVmqhH/+RV0ZIu1c/NfVT+Mq
1LY4Tij7JvIGK+SifXVnV4Clin+/DTuimEqjJH8WyuqLNCcVLQQ4lscF0GpC1ykg
SBiydAgcpmod5Zv0d/g8a3r5ZKxgxAmfU/Fx8xG21SfCydzuP58x2sn7YXRkhL37
V6BwxVIPuib2Q3Aoj9Ndc14sHc74etptf18t1XYOnIu5UEwGKUBQ1jzwFFy3xwQA
ohH44denXNUPkOAoYaLSp+ZrAo9oP1hck97HfRqPDMgVDHbXU6cG3JuwK9Q50Q/J
tBZMvl+a39dNZ/nA+VxPgVau59EJakd+HaRj9fscvBoETpAjX6m8E+i6/binuSIx
L3XMFLfQXrZZuzcJMDKDTMbSKQHIf/mpdAjjmJy3qc1JO2PpuxAKiTE/QzyzYXJN
dvAbyTUVwTiPYYh1Cu2/Haioz9PvlXEURNUuVaKGpx5rG7o9hk6x9UwoqUuNi8vR
2GgsAuaRo5l9gSCyal46a1YSSIPVO01zBVV5LFX4V4aSzWQofxFtiKIAwuV9pEU/
n762egMMjBSHDQTPBO11DYPZkpTLe7QwFfGT8913icxQ95EQ51muDcjN8h33PO2U
lUq8N5gc6aX3boiVE1Nc+sKunsu+Gd8zrTsnLn/aAg5jkgOyCN0H1ED+EtofRK0Z
WUoH1TCYNdOXWFAyZy5UMRjYnIMiWny3F0BZXYy3ImGBCEzo+yZgkcikshqQbfIp
ZAWm992714iskYo7xuPYBRTPj0/7pjKnmHfGAHQ52udRKtH4ppbFq3/pqn/jOUQ7
MX7H6NXy+xNQhz0JXCFjddyxf1x8l3oGlNoLllpO9WpeOfj/prZNWH63LXWf/GG4
inVjjaD8vs4lNIfLN83CTZfY5RRAdJ5ui1t+Y/BNAx/GoRQVZSok2iv7lu9R+298
dwxuOt9ehipC7jMG5KfgDspRkdxIYQnH/n+EY9/u7e3xKwsSHvoCP1NkmbV9kg+L
v3BkmHVFLARl7+Ln6KZHQmmMtcNDJSeqpiLLjnXt2erbyghQzRGN2rZYKVEDzKhW
W0QIJMehXFnMw93VneCw6qEhXde5qSbBcUvaNxqMGuRAKxpTn2KeTmgahU7tcsYO
qCxtvilu6o2prFKEvt172bKbokdwS9rznP6CSrARGnlxCZX4UmIcuOSuvoSOade8
/t7797RSb6zl1rJmUNTttKrv7KVfAT6VQNt3+NAlIRLLXSVynEJruIihWM4jYKur
tpbPqijl90f9/2dU4h2rzZmfNw9UyLtC5vhzlGQ1Ged5zaRQwPXxcHQM+YsWZLRb
Kg5mHYtO+H8o3M8fJI6i8lfgUdc5irJ2gSWTZ++LoLYaxXCsWHXrNQ8GJineqWOq
ZTyKmJ80ryovmj/NzRpjmUUmk5y6Yx1TasRMlsECwPlnj3BlTMtYAzU+PHPITq92
KR5f5ILxBbPk/nRmpFrlHt4ywBEX7dbpGWGm1x7fADU88sueNHON+ML40GL320oF
xM2Q4Khy/Ilt7YkcNpCAmxi2pWWX1yM41qETh+UGWfK5sakfPe9RbkzA7OTT8+TM
irVMHTau1q7QlzaqekLytV5D1w+T0N2UrnP+5NRwtzaukiePtzAOQ4WofiTlRs1X
2q8hbaSrbBSrIs4+v7Mv+B84rWPds1ZaLyJe9YMR+NO8zDzoOpXipJ5k0jibjKN+
HgkLPqo8qrJvmMz/yHf4M29U2FBbTF+bz6IMwmKx2cv36h3jitNrixgH7av5kWWu
+5dfESyHmXvdmvplaQTYHEHGDW7DYg1e6699P3TX20oY1N1hyBzqG51sWb3ZcHxF
NJ8jYNt/QyhETwNy1zj3XzNJHqHSgNwAm4zH2kasHKdRbuYXC2877ufFlYNDKGhM
5kXLqzIgT8AaQUI1FNgms1a+iuOnruqUMUTxkqcC7ZVCek6uWUp0QIpNLhDJfMtk
Op2RgsmFgR6mn0Z4KcRtTV88rap2qURuTiTJX7E9slGLl7EHYO2iQMrLVrSq9v2z
GPC3+Y7RPGRD9WQM2+3FomlJ7VC/VK5waYy4dbBckGiZ3tqorbcAkkNBuibA+IpB
tSSDEkigKqd/Wn/cIrh74zvcvUAtkal78cx0BfJPEF0/LFTpA+c+NkUcUEns/qif
TTZR1uo3eVduaCJguT9N7PIR8MeRCJNoaDFnjT/FAaiC3ZEJa/mHopBfjHz5XiVJ
IyqIFZnBtadHg5G0JKp46KiKm9KYMZ5dlZx2g2tZ0mAyXywFkPHxqtYZo6RtfWDR
ospyYoRoOZWIfuybjLD8zbrvKhd7thD8DWqNmucGUPHO7Xdfp7xQxFGkX1qaBjTV
nZuJve0vlVtzfJPQtW2ASawpEu6By8H0/VEnheoH1OpVCcvSEKdAQc1uUeZWqQqT
iYyR0cQ4CkAiSnSbwI99Fy977QSNsz95QN3hgYbtkh7PYtmDb8TNVlcsC3Keqv0X
mNZQVhlIiR226SjuidnuA5n9ypwBCRq6oq7qtx8Al5fAXlQi+FNuT2iTEfEld6DG
fU8gM1+TVLTdt9PSk/tBttEGbX+Con+Y9QntcwmVpV1oZ0fy3zfsnbyBMQgsRjjH
H4lANKX69/J9aWL5Izpr0WnCWghUBU/LPhATA9zSWB1FCh5VIkQo44TrYUZa/jN2
4DjwHevpyF3WxolMFQLg3/6hoKROM6CCbQfpQeRiA5tXsCTN0358KImEhbncXPzM
RpihL53y80jOqT7kMoOtJLtEsoaPnB5zevlcgN5NqsP9V9xf5lC8PJuZx1AZgnrg
xMWVHLVE99hxTdlAqKVd//Rc+jNPmNoQaQ9XrqA+bHu/xQeZF6Gw0NBA2BWqkjUS
AATQp4wnFbeIbZrP1ttfUedByxBxpKKgfnEnTlaxn8NzCwN6HjR3JOtcEudvAhxT
K276tMTvj/ehxc17NtEDfRJLeXOFmQnomkg+ax26J1n0rRYzh+i5SUxTyG30aRDi
CKYfdCotyLtVhhPMEABj0iw41JBHO6VR6oSwmPFqKF8JvixFtkbc+hYl6gk5wzLk
CdUW6tcnHfgRNrO4eBB2ek71HlGv/gwCoZ5u9VqOFaXgMj63fL/yoNXbUXHigLPH
6qXGT5UUwF+i/9CBX25xdIXyR1gGrY37LoaY0UVJWT2ZIqayAkHlLdnyzfLR8/0g
EJOk6IdJhQTpuykOkN+Lbl8ms4C5Zyl6ONLyuYmdphNaSfMy2vxoQrDgkuQhH+s/
kjB3WswqVsmLchMHyn7CS84Z2TXvFEVsITEGP06w+Uwsst+j3um9gtbFO1c8YZuN
36uJt4p8f/F9uv3tX6b3GJ1HBRP8aVNTt1NIxPH+IQPMU2wKbL66B1E0h//RxsXK
xDd53waBtLAJEiILV9UAvDtf26ADVp7gr/bziXnVLkgZljZkyVNOH1sQxcltwpTW
bOAsQhPpaEYxDOdWpO2jukLRXBjqnlODhRpqcUoXHpiYaVGHebiBwvD8gC9a9+6k
WGdE4+xS1kSZttamw8No04c7xDQPtf8xrKsKy/pY6G8=
`pragma protect end_protected
