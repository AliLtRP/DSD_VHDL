// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RL1/r98HlMTL6n9xuRG5UeGhRuXe3kfiAGgmNTDPgiw2UkB7C2M8s4rSSTNLmaam
7Dht1O6rlAIdH2dHOlTXDIIdsFb40psSPND7Cz9Z+yNI/XGCZol0lDUv02kbPMfE
YeH+PE0YP6wLAgVoeSbYrs8qBrIqAyhUutStXc712Lc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29024)
XS9dGnOWoK0voEXOqPWYDhnkW1u2kUKV4WYONKPvohXH+RhQVqjYXPshzIk1jPQl
Z6nTMP6HANfbKNODB2NjoW1LGm+yJ8NjWRLRcRJEAyFpARB9vQMNiUroQCCxm6GK
zTo0+2Ei49IYJC68pcDJKn6YNCInSMuICtWRzvI5Xj8yGP5pIJ0Hy/Y3m+skO8Fl
S0EyVzZnTZh3+3gn4dWg4jwEuPD5fUvmaA33YVoJhE1X/VTykxPcoOSJ7z02h6fD
7y+DEwRSfviZrVE1mcKznJeXPyrC10CeM/DgLWfl4n0fusH6PFKiUieJdBY9G0DY
AfKuN8TmYCRYv+OY6mNlwU+y9/jgBd9UB2avlas+rkNqHU6NWcCgm3A8qQsoLiK9
HoUNccyqNTPBOSgYgKCL9R7Hv+acqIbBdQHOYZ05KCBhnIoADxQfYo1dg26puIY/
VGFPIAYQUhMZcznc4fXsweeGv//oGokwzM6QtuzAAZi38aUzdtrUv2+LCa6HhF8R
7YyFHVMTX/6U6zqjZnVvRb9X5VPc1xc2XnUy6vjjkCHSh7F44ee8wWPJts1+qSBi
LOyyn9L6G6hA8a0ARWW2NQw/BgkRpgtf77Hn0rJ5quYNUEiPLLRMRGJd1q4ZSICO
TOC8YsTY5PGIIXq0W8pxkUOcyE+/IeheVVRtaFzfNob4uDrCFqfDmK1nZ1x1fLdk
XBeNQCwgwjP5THUY+24rmMCbBrpnt+nkkyzWVcyyRGSXQBqRQmtipmZIwo7hVpKe
V08rMVFcIoM7/5umz7VArlC24IG5/x3jZEjR2ZHo23WYXaDXEvr4jSJdoaO82IGN
GAE9OAdTqy44n3C1Lc3Hr6WApndbb8WEADtRM9opfFnbDDlghdiXO0LlR24uzDbf
oOTjZEX8LOtWmhmesSQqtHBUqu2JogqJQDo5Q4ioFpDhhE6cWmiu8mdpakuWK2eV
dqxVMZ0bGucoXk7Q/HXUfGXDe+HiRf/eeUdgBFMnQm+zRQVwXo3rj8eFwR9UBR8w
Dtg51XywPnNeGHYzCQi2lL3mpr6SJuiQ6o2xQ4zzNYu+zpTgItm+IeA4uWhSKBXD
Y+wmia/ky/GzDvqBi5ui6Of/p35lhcUjM0YNJ/4FS+YHC1ZfneVSJJMKdw1mer80
mNILtypz1tpNQdcXi4N8KCfDnR7NnaZ61jfNxQLRpV/7GY26awtFjm8o61E7ad7q
8XA8XmY0+lQeSomEABypROAMXciSPIx2g0XjBv2TQxDmZO6HJ6VVRJifn88uCn0e
tu3u/Ff0dxQExw7GlvsE/Zu9tDSd9NU6Xn3le4y0tii9cRguz4T/GrFZwWPuypdR
kHRh3dBAzgPzyoGlphJw04TQC8gGwRb4ZQa0RTRuV3PzagLxcsaW24ruH9U61+rS
GEAUEv1jrc6viUG12HTyqPzeKznQjvaJlqFm1nXJcy91YIAito825j+GMOpbVCJm
Uf4c8XrF0v2dlJ9r/Nh3yj6yNyOrhaVNRQquHNwP1lvJwI/1K3V+ZgAcOyBDdsry
7NKIrTp5FZ33gA3n4KIpVirH1TnpU5AkYy7bh2wlsYTQesxVWYcf6JSI2DSMjQnE
yZDLRxlO9tTwKjigaYlswys6HI5SvLnqajROBvJ8l9F5l+s+azQKA0rXqvcJeFPY
PSlE+zxr/NFTLK17GmGQLxDTupX/pLwIoU1rWlsgZWMpUentcpTUyqQEX7BpiWtT
nkW8LCBI6xLss/ULDELUoFNsN8rwvstvrAylxWpt1jK19lpFKHRsovlQ6Nko0n5A
7D4bUorgbgD29r31DSJbZSR8QDY2Q9lVYo0XWFlxxvfBrGAHSBV2w0C/G3kvamVu
5QfaxhNodU+6DHNdqrTUlSFNhZb31aRMoEMlSKT9U/xI2R2379BK4DPkdj1pe/w5
qALtXbQ6IexmJO4qi7QUhrElAt6/2hczzJI0ACUH72jEKCu3NL7l+5z7dW9X3tSZ
T1BgUUgUFe2SCRmHcHVUWTgS2ty2DF+9273KqmZEjNwGhEyc7iqAMGUfgBVdZmdV
OKHwrgTaWxIXbNYXvYeoAPEZ3rjASGJ1NVMzoHcfQd/9l0NkqvKY1bay0LDFjYEJ
afh2ZevmqMuROFHhktNA7fzIXOyQPy6f1qGb/HBxRkC/19C3FF20xDNUMVmV069c
FKKc/nOOAaKhv+3bwvWenUi1lEzwLt3mqp7S/4wrukIF69Qw+c9lgCnNhiwvE9tz
hr4uhaDpwp5EdDYpoQYfF7fPBhqG/8f34jRiWwkOt9dmj6uKxZmLR4eSbOdSO8tU
Vna0+Q0y7lNX0FrpbMmM3BQ5Du2jmmL5p5UdFlQTvX9Kr8Eu++VTssjhtE5LOOKD
aUWl8qAsMRnXuMclyzt6CUsyZKS0AHFRvJ94RBb+/nf0ItyAAPIrmrmQW4tfE5xd
Y1RuFNVsOFjrb9b6LTVvCaGzT5xbPzQyWXy0lL6zITBm6HxtOTz0GKTwl56z6rai
nFWtZDXHj6qm9tJqJJvG5T25OE/5kGiRWLSO4V57+Zh4MUmjqyagpvYk3YoVe7vB
8jdx0woyXiC97Zu19C/eaJgQ6YuLhy8AgIGq+UW7ImMAlRRd+d9IFx0ozaxOmkWa
csOaJn6FMbeOVR7pFcbpQS7Z/zuEi4btkPpZVxbu/KBuD5wJohOfO7hrSqFrRvUa
3KiJEN6YFpUjcIFlWHcxgDG6T4pXynZhdKQaAVH4Uz7HkBYYr2h85QBQaBia1HDF
qiB9B06wIdVxxylrrpEUGL/bd0IZwvp1mPc/bUVjJSWOTUoi+GDyy0sCHkUfgy8s
tP8CiXSJvx5q1bgsC7JNWm6upinaRi2HWQNR1XlfTM7/PUAc+rxIp5DXm8sQ98Dg
0WcIz9n2LZhFn+cFcGgy0JLBeZMdtVr3bpJt2orM2hHeFtzIzwQ7RBuH2tZ21d4d
fmfOHmDWOdsgOjCE9ZLI38AVhn8xHEPiT5Caj0qtVycscbrFb7Zoq7F/CSe7IIXY
4yOVoMOCZsWHzomUde36FYoWOvAts+906Ov6t3RvzEtEccD96DCnRk4BJG9r5QFQ
kS0GnmsC9OQHzB7DXkLIh13+62aVnTF2OBgUq8NoGcRt/8Sg+JjD8gdh/1bz2uFr
cYu5tgRkZmG5BOEZJaLYBr35z27QJK7LbzhCvUNs5mY++Js81ZIh5kizw0FoPYec
b67f2rh15wFg0y3V/ExulD9Ig/3JmX7ja56wthn1SBLHpVBi+YEmRkxMgcEaAbmc
ySs5OUL0OkV5OpyGCiJrr2PPYG3FkGXHkcNnk6b6/kri+WUdJ0j+TKexhipPd6+m
P/+LhNBCNBZEuEIlzb8UaxTK4J4HvZh5p21/8+Lxwi9v9Nu3jxBU1b/EY4C/tZuu
yHhjOS/Klu+Duy5wTzHHg0WwHAWsmdJ4216C0LfBgCZEnfGlo2YFILHg1OEFzTof
mJMwkwBzBkvHeRrChgXAi/uuSTFAvWE0p5w/v/O+1HFM8hLmxYJrj+8GnoRukSU1
Y/KKSMN9vAnqaTixFCN3PXn+6tL6zSVW9F+euA0QEBYte5KSDSmAwqbLgibl0UOU
I6PsXDTIwQAjSbkG7ykDLQ/IvKgvIuKO02uYbWFxj0aM0M93K1aYfXQAkoBe6nrn
gceiDsObyrRmoPknhu90mWujSklV8CACdIquNBNUsOMgZsFvPXbk303mMMhfZdTo
0UX2rh6tCu74IYuzjHAQmL/lcB+Q6zpHot/xBrxY1a3NXZSzwOCr91min10nFcJf
kEkOgE95VqrSlSnj6j9jZPSh/YUS+VTm43ZqyU1z6qS7ZydkCUwDciozAl3gMCZG
P86gVbY7k4rFMfgUavuWuDQQQhL2x9ZcBKqZV4SGabrOITJwYbRWqWBwGVvhN6O2
kbVpIZ2rL6eeE6clKvFPQ/VNFhcsrZjHmBWD8feBJqvyM/lDBlYjKCfkt4nUe91Z
cPt57vupPabIezMl5/COH+RC9SFMDT6b7R8TPgcsUdqXFfkLMnoIwIBbmZDn7m98
g5Dp5Ft3eO5xn2Dm5QUdEWu2lV+odyfteyTOQ5Q+TgBPR02yS7KOdJgyvjNahBzH
fAKP8gGqVr+jj8sow4zxk0nmoHkd5TbElqjIebXel+ZDxtQIQ1YjDb2rYdJndTgp
vwYlfx84K2PqHKoSChQ+uqWR4A5NV6faasONBzyIBFBypNvHFabQKRZ6y3K53WUc
If0UBtIcg+W/xc8XXphBk6/V5ncsn3GA1NFPOe1cp0UU/hF953eGtnvg7p2UG5ye
Fp0k5BrtQa6OuicHrY7fvBzLLr2rNeYQ4rDhEXYtCR6GYWxFVXzPEXQfjVFG/vj6
gAeRAdUfaBYXk1QOCX20cl3pHNhCs6kXdfVbUNGnWhxKopKTKlmfiKPaEGUdRuLF
TB3HmfssXObTCoX6fTfpB175Os3KCnfUb5UX97ALDUBcqOjXW3vQAyZCWLYYH3SQ
IfzHk5T6py4Xz8o0n6CPgg6l/HOQ4nNaIMIuok5MV6Zz+en1t6WEFH/niv9z9GGK
nkedeMEz1Tlq20AuR0iyctsC0yqMeJBZ2jNiLZTr7svGlYnTiRR4frjeBHAQmYe1
jdOILg5IR9+0fjGTpMV4KxeotzRfjvWUrsqf26azK6PuqNkFDAuHbKwoBmfwz7R1
R1wDtgGCzJZgrlF7zEC6asEKTOwuLktVl5t86BmG0F6rgfdqjMowLz9FmWOR8tuo
6HF2nNKd01x6FFVLkNdXlCb9hxJMnizW+vGwfwRr03XfTmrIDRHfZJWh2MdT/3pz
eRO8jyIRNjNElD3lhOn3ZVeAjC23p1Ja8poWNy1IgmxKCB7mSviBtDCat91h6KiS
5o32cv8rAP1xHiyav8iAXFotTvV/CjlFUwyStpWjTxhSzQuzQMfyf+GefdhEjQct
u1SV0bpd6C7t6wewan94jv4dL33ohFK7Nz7NXY5TJtxfvovPMT+jeMNu9qD1DfNr
/aqYg61Uah1ABfvoYXPG8vRUdTWlmevcqSybOkqWAJv2b8Gsk69w4CV+Q4jiDBaP
FTi4H9bPyvwAInvpgOhTwOOdzDZ/8YAvYIDYhpdIXvCKU8tH+5ObGIEV2ib8z9XL
YjzzilyV8h3D7hR+74ZGOcKhkiEDHKsX+zYonScmVqjctCpXmaN6fmps46i0HFO3
D+NckzVVM/Z40kVxWTmylgBN/E1SkT3qD9kwwN1Cm0rpmzhuMXfVlDjhUj5jZCx/
b4Wb4SbAmfKRYv1VAXvNG20H/2PaQ6yktGuiK6I0TgLEuejjMS6Q9m2N6+r/MGOs
GINM9lO++i108r5+oEoHv+2sckzcDagSwiVGNxC9/BK0c8cEh0HRvXblOwr+5Kzo
v6KlN9gcHmT77fW7N3IZV3V7oho5sNG2ba1yvrJwKNfMeK1vu9nFWen560gwB6BP
rvfltXRYnvYsRV4dTWzZEWbdm+O1ea/HfBlM1BRCE46yAeYeJKBGiOUcu22lrrhs
pgiq9GSknYHObqDpJ3cyUkjW7AVClMb22GUjLr0NkXg3L9iwF/OIF+ZoJ9807kV7
Iq6izWnkwOB10LbOsWB0OdQmYvbAUZqXjeJHDLx0krhhnjou8UGCc9dpa32R3I95
0lMPIWCpsP+rjV3j/cXz1igaCNUv3kBAyDWFoRKCb5XdMNo4+Xmsf70LPvdft2aO
E08N3Z9pKHg4xVFItTJcWHStizOpPgAs014kwcRwAtZOGkSoEAgTFOXbWAzThkqe
6h0PgVbGlbxhppjz9tAiAjN/a5lT5GdC5dOIm4Wz216/N9nY1qAblx70nD8dpTm5
Mz8dmO+yq1N6PpBdU/nuxBtnchmNvvMLxm8r22g2X28zUwat0Pmmjv/RCuhXCy/s
GdZck4PaEI6S8s1ji1QPvxn2a20Go4u43ON6HlKj7rum26dfGpzFk/AKXI3donp+
JC7S9z657KS0pz/Eqth/BXDuvWlceA5qNWhQDee+b1Zc5L/KsmgS2VjYCLu6Uk/H
ZjQ5xfFC1o7oyf2HdOfsv1XiJ7Lk8GnJa5OWERxGejb0E70nCPKLc8BLO8WOyuti
C4aUl3fCfp8risMPJ+2dIekNakWSE7/OA8WERDy0DsgK4QzCryhNdPiPoT/tnyO1
R4jvP2dKMU/NHTrejeUGKkXweqQzVkXiU6V8C0zaijZeFCEcAqzE+dUz2y8KDEiT
3EuzMBMc89Rm5nqN1icJb1w1YEVWZzztiELcaifovTAH53LyaCfCdiVfnentGZTQ
9kCz09ngiG0U0Wl8JX4OXflhFZUxIz+NkEvx9l3JllqFbeJshvXV/IjvXmZvyfsS
tKY7WkJ5tBHNw1lpT1mluFztOmxS52IwZ0yBL4r2zfEsaKC8nIjnAZ5l4OlnhWHX
xrbRplqeWksZbygNq6JVY6oMikfvNBWdwqPtYVFdRixVIjP0Ggc59yeDvQ17xwc8
2SDS2+tKBcXP++i03dji1DEWCcT3tvLmWortadI78K/HrckRmHdSSFGOn1h7d9q7
yRRLf9c5lz0+jQITbc6Z3NEioi/iGKEzkBwGekESJIuo3rZXldKoTgj3GkKtpH6a
M2rjRx2MQNbM2rRFxBFR6V5jsDF4unJvHYIk2Txzk0IT93EGoLr9Mmnnn5lnVU8e
qn+riB8vwbF2yaqgjCmSwpgHvb1yKvh87d4fhgwkcZjmA8XBk5FwPWUrUcPQIwVh
uRMld9ZmznvLtYeiqeeRWhjk1eWLlQgVxEQsG5BXe8renZ8P6UxTVzzGShCfH5eO
RzLSfvC/RW4c+vU7acREw14UtTcxFpCHdRFJiw0DFwMwyfVc1OtmGIbZxBdTa+qX
PuJxsSb8raK0T6f8X6CJANEiU7FEB0xArgvPQ7jOkLJlM1DW/str/glAH21sKU9d
xGHbOHtPIbDzT7nEJCd2ehkv/aQv/Ajv+xBrx9hgLB2EJALDtune8uv+QobZDS6X
OcIDTVOrg1xUI84cyYigNryGqkTIq52MfVW1G6eRg+pkUYV5WVxyoQwe/PzanNVi
VF+b+8mcdzqTRotVjU5pW4hcWc+2f/GCjTboFlvvWuJEw5asNylMOlWzsofC5r0q
sPsJ28iQJQ01As/LKH44x0NLt3GHegABe1dT0E5C46xer5Uu5mrqGdxtTjJII9rf
gzMqJWIxVjAYl3BRPKIxJqfOV59K1Hnq1pDrr2o2T/cFohamp54uJKX2AaIXk6CQ
etbhUjJNEMfLBUizuYD/M6/T1scQzCL/gHxOxk7S77s867VJs5DHD0PUPNPvUZ7o
50INtaaInioxBT50aASiz8B5XtoEz3jfOg1/wRhJryyhcXAf1/hsltRZzpP+a2Wp
4A+t65d48Y+2yse88tZU0thwFRBvnRsnMyx6oRjiYyNq3rpP2lz9HCP4usS5PVZm
ZQKaj80Qir6ibm6JNlXTOUaHEhEHwfDlJM2rECQUEGdQzkInl2VnVE84LaEcqb+A
ddqwSqPwpro8O2SdX6p/OvKsg4YN97CMJlmXB3ukDZcYtAmp0rtYrYsDnT6vALng
gM+8Ud1m4CuV6+TrHxZsaNHiwxpcRKwBmaj9Pe40c4pqm69ZYtVKziRN+O+UP0QD
/8s9styg0r4G1m+RTEQZw6zv2jcv5ulmkL1D+g+CF6I3wjlOrQic/24lGvniAkqJ
VMb1x7H7yVWytGjxx8A5tyWyBAw7eWvxQJMxfZHDhhXSSZvS6fzOEfiFRyowhBxw
7LjjnDow4tgBpcy/ub4v3b3ENb0+JvUu4ASRMsnl5fwxSn1bza4JAY+AWk5lBMoS
vOnAuPAZiaCZ7bgbKj3gx72CV37nmL1aKN4N3Q2GVPAYNlzolLyeZ0YC16Vz6km/
fLiy2mPI9GdGKGeqzXQ4hRZ+htUWZsN3AAUSktUeaJkR0WgV73mkidBU0xLRdUue
Dxt/TxM5Kj538Ine/y0HDQggDGeBDaU7VZ+wWuDuX0Kq43sb9QGyTCAsy+NM9zEZ
OpJYX0Bp4kE7Qr086hBhR4ws4IKS9z1A1iJsxOkk0zArAHEdBIa6awkqdVMPAhac
5/hBorhUryGKJV5TYFGgkXXGOzVnKRCJSevJzjDUikInPj76gxYzGPFxh9KBDSJm
VbgIC+X69XjLDJvIWebEwvCHpwW7pgKZdxtpkKZxRHnyQWEeKr9KKkdHo/oE3H35
x4ApvNiKssjh3R1fCFyJxAkhDC1ErNqoUO9I93UPetZzBOTqnGFplNt8sXzH9lnK
BXrT53bWayhUGEhCmaQ0ZzKE6WRzqbMg/y4WU0qW94MWn1ZCoX/H7ttC/Iaegaf+
djslfU/7NhvJuKISxdiBFBT6izDsWW0gI3eWCrdvETPyA8+cXt9PUJesq+0g86O5
wEgVMWEPRdRIwqJsmeP38fyIG8p11xCuOCtwTsvTMn3Y+avbjYjM/Hro1C7Go8l7
jwzkXqgEqZDW2D9FOz925F4Me6sNZ19jvrCoJpUKT5J/+bw+XaF3Ly21T2ENZj71
eTt+QIR37Rrr8n+rlXh8/5yxm6IX2vYrk3nO7pJ4Cm9UV1uVI0KWqhihe0pWEKBN
9QdLNSidAnwoOEVvgWOpWPXf4kBE61VZYoi3r77CPevttdBSbvYCGTo2vXbyOY3+
Dvnh3o5S/GyFSIhs5awQaFMxJRf1rJ8uxyt9aXfitsHfCi9f7hZVFk6DiN0UWb2a
3zVrvitd7w+HCi/MaxGObzaE+XUzbHe5AlfRoAuDrkQWQ7OMxc0FRyOxUTJXetcp
JM88sbITXoCio4wOU7nZtCK51gVEX09NOujfeZrbR1iI/rtA1dPknr35KArowGwn
bZU4A03S0hpmRbp4CwE3TZhiIw7CUjwGE9jXmypkFdj50yg7brI/7bkqcotChMgq
Qa/R84y4Qr2ZKfDcYU9l+bGU+p9TRYjyXPzc+6sCL0VHTlvqowWzxUDHnwNDOeCe
NDs09r21Wg/fhuumPFuQ4n9zNnsF4ohTUlRWGEFtPTW2pIdCySI2HEt7dGRnMgKn
Sx9JGUNsH7RCyvAhZE4i2iBXrU/Pr2RpKxHN8MaIaKxfJXWQyuabQfwAVeibTAcN
y6eXD0Pxa55FhOjN+iawG5lzYtQfmcjy6izJGB9vTB5Aa7/ivxz9XK4KBjyx5iw4
1HWvCTxlZ/sh8ak4mLvLXyjkqm8WdL2gQdyBNeNveDy12xye2OZ+93IOR9hcqTeq
/SDbL+AT1ODdhgrMi29Z1irJ/CGx3hY5PxKanZ+qAMs9iqZrrg7UgKg2/jkwMFxY
uESZICR5NJKbPFeer3xZiNAQ6grE+HrcKr/hyWLBJjOfOdTzfpmnmcLWWeaZhTsb
V5ioDfemy+vWizw6AVFmxClNh612Vrg+jCmKEinlumRay17Bc/bO+JWqf8+Ma6iQ
aZR5r+gHfzUxSAVEC1rE3Fvx/0rYhXSsYoDzOSjnsl8xObDNVyjxhC00UzKcHtD+
OrduSQXDWse1EQqxK5bWWSqrJfi+ZdyhJFuwIBtBaiL2MifAGxahIUuMPo0EVCg9
B7FEs0cPk52oZ6oMScZmABBA14lLEHMHwpexF1fVnEOM7DMqiIQGWuLeRliF/Sk1
Rm5INbScdzMqCwfmDImMI2F8Nz1LV6FBvB8ua17dg6b6KOGD+ewjU9tcobvsRA9j
5WYsRiJiaaYbpNcvzStZa1QSdMrlS1+TGKQUH4Lzg6R3klG7x5WIFXpbcNLPyImW
ItRPuAh3j1XDH4BSZaPtzmNk/J4gnO54RIQ7ZhbqAvvrNZms51FygBoS/nJihY7o
R8DNL38sMSzDRow7v5SUPpDH/37/tblHlx1M84vk9CKqcxdK5dCR/OM0vJMKixmt
qmVlnTaUlnoUIqG7nj8145oqOOrvxDvn0gEgBEnHOkFyXu1VTCd6h1tN5o91Lp9v
3+Aq+GJf9hEq9b8XcrwMuIFjCU3c3VEg+1CgFWdX9biJsW6yi8K461KKsXtOVv61
TgmCVEiZbQ9e00MhFHhOpHmy3yfvyHDD9684nTrpguShaNFeveNJ9cH0xQa/+5yM
L/A0I89dcBT/c8J1O8FYi+KZ0q8/Hp5nzSyo8iAc+ndhcuJRwMaaEyl9Z16o7S/Q
hB+wazIjhyUTTzEBFvHiJ4yJWGi0FGeYlkgFKByjjOUi8UvB4NxN0IhDkwOYetbP
s+J9T3baiXTxDgbjnBkJQdUbe4H9PN4wVXJaoz1mbo73ffZVf9Uii5AeSL59wQCT
ysT/gMxduQMud8QQjzA7XDJi585Brh7v35QwHg1npubAJitX7zCSIutxDl+Uzozy
c7206a7zPFx7HBSlZLnud5CFMVaA378coLN08Jti4bojFrplXyWWNmLnMsM5T6y6
EGneB0J4thwjG0Pki4SDcnVrd9w15vkPlQzleDUK6oQdcbphGTp2ouVj+vi8LdUt
BG0CVDzlGx1XUMMmLL7jklDoOqVPLyblzSi4NrqfBvoiByyq1XxmiAlu0lYuQ1WD
A7Qym8OmuKSmyI5QL4ZYPavLYcax6EuIdqQL0+nAbhirR7DMneuFWweHJ1i00sH6
WuUbnaBaju3tsQ7tA/QVV9qOzf8UJb3kOYoQwNaUEAz53XMkMavWhfX7ULquuuxI
a9avlOh5aDrvefGggl8o+fc17a+cZZdBGtPu2E3lj6XW9j4TJUUePXWMXHQC1o5s
xreEaI5ypo/EzsHJqaju/8RKFBU85Z3K8kfEoKwi9SIxCEXh1g0HWk1G2ZJaFwLV
eqGL0sGPCFtdU5Ftrauvtd0PHE3nJeb+bvFnOlBxNFAELrK6uT2g3WA8gJVOAN+S
98XnSubIAuAtYa95MxDMdA9a7INuCmoGbWnLVTl4PA5u+uj26+KDATgIjwdKi3KJ
w9GalPdyJclxF4W/IeNJnEgd57NrM2cvEmllRIQr5j9cBe0L4lvlGFEhXPWgxZlW
6OfjvS+tkeSoNu09/OftMSND2cy4OJrqUV1Y+Yf2cRjt0p3xK6B6cbf2toRKabsL
APEvApfCbcg/xN8dRueGwjuOirsU74DRTS+MGVTnjhvu5MG/BFlumOj2paUAQv6v
65Yzy1PvxQk0mLi6ScGJO5UNlg/iQ+jmXkAc16Q8OPsywULAX5F+dB6Lq5G/Dkyy
obeszfqZK56Zb3WYwG64M8PN8Q3SQlIbTH1StyfdQ8osJwmq1Z7cd3w6N8Rj+Lte
wEltjsG6jQ7pbxZs8TYp+k360cOVc5Gv9JDArlYPAwSzePW5BuaYHhwYCgNSnrvJ
uSK78RTk9uTjMuvS/h+knvZnbLdZYrdw+wU5yBP4CjhgBn8M5siotB8jUPJlqBs2
C1R1fU1790c+X2qwB+oSxxgypXMgtVacskFnz3t9HNfZBB0Ix91ubAy4bYOGYDdN
kzTgf/II9WvsJ07U5owe2TIjfEiOvcdmd8xdro41wtgh9Q23GcoCThWOFTOPih5c
Pv53U0eTNgj3kwHArCjNqoSn8oiHmYF9oSmtpQycD9iite9BH0JogSvLaqY6ZzKT
uYDsyN/DH87quQHGSkUMVtung0rq6CC/0y5y/9YG85fe3/kBUuDxjaG8EOSf4/o4
f/e59XzsP61uP6QCMOWKZ21E5Joyu2CDJlGaUTR9ULCkhhS/ucrqJusiScs+ofF0
J8dVuE0ObOQApTfw5JTmXW6Hn6lCEjC7zl05aqVMib/CGGEa2+Aekw7lKh+hLH0A
i2Pu278x+k1DKTdSG2Vt7rLHhRHHtMz5UkZE0eibhyS/0dzx3yfojczGwK9vRLG+
vkHnAI+au2uK8/C4cby/kIIiOa+EH0B0DJE7E+2YLxpAVzd8Gx13e6PdvyfdoCRX
U46Qj4wdNVRT/dI5J0vhGjX93CFYkydXAsswBLh9jlLZDSDVtSMeC03gz1qqqeGp
lLrk4TdjeRrI36UzaN3h1euDH/Phpl1UtyOz41cad/D5j7AmUw8zOyXC7SgqkZ4m
9/g++ojX7MlNJwx1yoSk/e61a7ZyJQAyzV4Dj20lR0bPFcuSy1jI5/jb+IpIsn+g
j0Lko8672xw/HAa3+B82iBMYBT9f/kcKhKIhQEj0rDe1mRwWwA+W6PH0PVea02Rl
b6LZJ6PKI4j5M0/asq5GfeTudWQZGC84thKAe3+BJFR4MY+FSz8CwTuZDpMaDFmA
f51jpOebJwmCGpDoZ9hCzQXImtjCCtYJE7aCJ+xb3oB5eImDOnaA1c+q/fXD7Dro
qnqKpifXb20A10nZk03fIMJFBPdOj8N8TWA0AaR/eycFLmXO5VjA2AtF5P7YQsLt
P80cOoWYeLCu/esLHf/zCUrDkXcaFJG+pcRf/RR0ZDdbAAOPukl/hN9VaOLS8XYA
AdPenv06K2QJiFyObr4x3wcaxqWXwxXFKmNf0bOAlwSZopZjvV77qIaXnA2saoP4
KlHzS9rayE5JUgRCg0lKcsxZspHFIggus+qvEeZ8mBjtVz7U/w5J1/z7Mc6MSqEp
L/tj+evbQXsTSDkj7tgZqT99OA9hETaGMx4MzeWGjhVYi1Kc/kHqmiSh+TxihRPx
4mHSKXJAVYRz0iPsXSrAiVT2pvPYhXiDv0O43wrVgHHOO39G/ftQ5v47UqwCabhx
sAAo0spSvulegFnzTb9zds4n29ZvrAcrL+A65UC4mfQnd5As+sovXUGouLhFIGUv
mhFNbmBHMgBSfDQfNFdL3X1WXqe9NacvfCAaor0iCU8uRGxM9BOYdP9d+Ctrp7Uw
TlOmyfR55QmZ/bw0hM7LW8o74ysQrcixHkINI7bv1UV2SSLq8n0qbQkfgSeY5L4u
9qmhPumby9R5mTMjEda4AQdzDJMNY6b38G/WQi1a4UJfXjRDarfFp0WqcfhNAFzf
l1AKi+ev9blbFmOmFdmvll1Q+h+vkyDt1GvF94uNSvjl2S8ZTEdEt/1OkhI7cyHs
4E+s+gY0WgpdR2lc8F5EED6OAenQUsyZDGcC47j4nSt429CkvBGTMC17E7XLdrEL
+LxtyAos8Oy0rT50uchXEjUCmez2U/Lf6CmOqMG40U5pAWUjwOmM64FPhTJ7iEDq
ZI6qde9VnSEXQr4hve8GhttdBczPl3+fvHK3m5kG9Q19VUWR+pmC0ZhlIo3G3SOU
aI1ZiZpThl3lXoQyG4RAphUvff6Y5s8iHZXdvOB41b96nYq7Yw0h5N7/Ohft6SAF
XCrWBGgBbuXgSB3Y9VPp0kpATYWqahUWw3JGDWOVCCSpwpVYN2ovbz3xnZRcbBiF
RBWuwrmIzmva9r2SiPR1n0nsl0a99p1eYfVNcnVC+Aq5sqpjxk5IApe8iWnyEmUc
BiLsTGCbcM2dbk7B/HOwaPBAI9SgFYSj4M+3wAKCpQunTmHa69UEOvEYflpuTsTy
t/JplY5Z2vDI+lIl9JuM4Ay84OWYDJjU386Y1E1pHbhx2FPDZjZ2n/sA3QYNyOXb
KmYyFgAu8YNBbW/xCKLwHFnyW4sbU3Rrx6QZB5fNVFFGIR+FJrM4UoJvvlx9ELHW
+HUcr5ZDmkSNxe9hNQr1NJ/0P64qxZJyx7hPoK41Eo/s54ubmJ4+YezmWjFvDYWt
/qzJFjYG02EdOWSwA5dp4gkfXr1zBwT0fWP+QHkSS7aQYjIXlSe2OLmw3/jM4pXz
IYRN6ualAHm4vXqOoJT061NvajfBX8L/xeCSfOz7ViqJH6BgihcjY1tBH85R+lvk
dhAnICXv/rVD8vGfH24Gm7X2ODJVxBwcGZuCXE+F2vK7CzzD7v8BUBIhJO2sdkKL
4cfLW55F6K2OdH2Nk5mUPt+wIVoXkaoXVPdOUOZ9RXl0sCABeYXm0LHSzuDUnTY7
F9wzUHNizpTtUX0An1gXZC1MXa7PwtBbR181z6GAKE9N7wRXU7ekA9J31GFeFEXp
mmvLIwM0jc3lK9upUwf/s7HddemeFrQYScYiVFKuX9/8i0IslbC/29tXttMEV5DQ
tRra0tOPJly+sg4FkyMKkkKVM3gHXWH++OTZWxVMdw/RjmO4VLoaCFSSUEOKjKPX
+645Nv6W5WrnxQeN9xTF1pPTxcJZqD8QpnYlFzXWt9HuFLEuxtp2MaWqyg5ZvAaG
AM+w8/kF4/379H/o96u4cfBiqiQmzmT00+IcjUAsrbwLuTBmjYBtPEhFu4RbP6N3
TCWNKTVc00xGN7vbJKA6NV5ZE5lI9zEF8yaKENZ3+lwYAIR5FI0duhllNjbMcZjB
FB3QF+ztXLF3uCS/YVPeYhop1i6fMh/59wP4IdHk4D/eyCzerVKf2qQ0YKUjCUmS
Ip2+bj2dRZTSIPipI8XEpkDkiv2Zo+VrAuTWwuYYhGTcZg+pVh9xmRVHwwndDjw+
hp+EciZzbS7p9GZ8qbSTDtTZ8ZTYATcnZ69HmhzOPvJoxctFEeQXZxKjWvfTzwXk
+sKvJ/YNCbdJ5pYSkicGAQylbfMOYjP0lW75x9YDpVjB09H2/oNcR9aHJXSbC32Z
vrmJTAwBkV6/aw99rXUlhOfwO8mPvABQe1HgsmWObW9ThnayevpCLOjLvy9WyARy
1wbgml0RJA5KMdij0E3UHkRhU/TStRektoTe8oF9DVK9JvDSZSdEp+sT+IuJvQyK
nNEwa6LIOfl4HL4RjwbM4jrmwughhoU1pezhdvzQv4jmfn45DMc83zukWCSNF4nD
7/IXziNY//3sa56R62pC0DQQtcVHEoIgegUR5Og2GM2M+fhfADRJADG7DhMu7X/3
ILCH2dtqR3xqhKQp3C0eNtko+aBp4vWe6jwt+3o19EMzJ5ZWCfsmkIUosMgOGVI+
ITpFdUDoOUDriVfunTGd0n7tQY02U/0T8jvk5G8+08JunSEONBszijfykFqWr7Uu
rw97AP1lyrxNCkFyeK4kMEWwkCWboKv9mK/LHsQ0s7z0R5GW+QX25gXa3Bu2J05S
PF8q6hjZRpyDP8cjS9+y7MdbzHJWN5RZ42hSHALKxKe9FvaSd2m3oq76eNlfGRwh
pS9fgY9lRT53YNYBh26duiJeK32mJ30dsWp3i6foKIX/R9x5IocKYA7RxbaA1sjv
EU1Bm8MEgo1KIhBBPAhTCV623sz4eMt3u/SAGVlz0o5VeU6WN7cZ21g7oKWjXO5r
+rXKDO17Q5+SgBqPPYryB96wHZibHqp1FB4LhQZ9apx2aBge03Lj6vNKIhhg9Ult
eVv34wKG56V3xNKY4/m0eEddDkAtg/cVa+lpvpHuw1RWndiNueRBpX05QY5UeinA
rvZnj50Q4Vv4m9Lie2Tudq9jgyId8smZK/SG5XdFJIp9bhTaoyLcKzTnHXMdit3M
6Y4f2YTM1CbYMcfEitCrY2383AkoUhvXDtCXbF3Dp/0A0GkC/AHlUkQCSz6VZHXq
saQh+gLuRFwLRLVgcEjeUaxfAl56eZlcpvEFn0NE4StxNGCEZV7ceVKZBgAxMsfa
g1IRbzVjN7MTu/pvy2tWZCyctHa00icxHAYXBLLrb2Tkgw8uAXfGHuu2vw2+R+mg
8kJ8OPfssQe26ycfra5ctij17NjcOPCg3LQChEMiFpACwYjSc0UxQXLyq73TEUvu
7j1HZPrUoNF20ue2r3PS4bKgu9eUHwOhwA8PVsNicZ7+NyLvFLN4gsF0fTUE6I3a
3l/gM4ki/NVr40icwdYBC6hZDfqBOIA/dmcR+Yaaj1O/bO8pkv1Q4j+iVP9CSb9D
6mpgLUN/ZTCYiPb9eqO1LYj+yYLugFSkw7Sjc0JwKh6E3AeJ+MycWd5iQQyGe9CT
gsAg3iyQTIIiQgZmecuj+GgOwjXTazBumhFPlZe043ZiTzjaAtdBhn4VeE8QD+S4
bGSxNhvql8P0akBD+Q9KtS84/LSGYAqOVh46GFxUrsJbSjpYGkHzCcPANuOzbX7P
qFUgXGFXVm5BKixRjc6DkM7jK7+ZbxPemwlL2vwP2ruqk8Mggf7d39XGNl/028Wz
OFjkYzc6GET0w4GyEvNVP3h0tt6jP8Bn4+f79MiZlqHRwfZd1DipGnl9E3Qhc13y
+9pZbAx6kya5x0g7QsqO9/c8eXRAXb9lBRRzrf6LGOt7ojhU6AbPjHsx/BDef99u
T9cDKFHa3Xa2KlAY/LoOjj8sYG414Uf1xd56Yf+Oixexna61bTCWhVl0HHGmX9fW
32Ck2zh5hs2UoY/HlRvZ7kZTgtab0NtNkCL23O+7dqw/lT35m8JcLNE92oWzyVOY
bgQaowwJM/4tLsHDp5/WtpJNZvzRTwQF/MyUuBdjy/P4h9lF20U0NI+ZtbOQL6je
RH8ZBCFx54mX6ezSCOHu1r4MVFTeCk8iXicwJLUwpK0Z2Zx13WSLkqbMwbGpXnDW
zge5uGZnwNgz0ysdI70NQM3wMT7sbQ4tavC4OfN2vC3vvU3kG86ldiuY5jKCHoJh
9vv6pD1MVbziEpwL4P7BdFh5FQYtQduQ9evBGMuDRA7rrUUalR5DBXWmSPbOL/7v
zEW8+7bXv8m7KtsmKwhU6wRic0UjK4EIxa8I966+EB768zcZePDJAWM4jOJhBGLe
1ZYoSLpp4eEnakiQg7DheY4KxwLr8u1ZFCXR9YGIrhIgV4ms45W2GZp5Dpc6hFJM
8jlSFttTqZiNj14izJx1IxvxrQVpbs6gClkblGyJaJB92eCDuc3d9jIMQCl0ZZK6
PVlOONMvqyTuTPI7CN59AWTHAfPR3MZSONC0aJAQgaqDg8vYe11qnbjqOc6Ez4Ro
KFelL+4onOMlo3yIni0OTsITqjQ7M1EgNkVVcRLrqzIc8JTQkXRfBsrjjYqJvDAh
+rAhCrdyKYc3BKyjGGM2mrEscNskAxXFET7fsxJkCf6bXXwa1RU0Sw//argNLwK6
RQG9eJilydF0KOVShUQjWZbyAZFgxxsIFoWd/leZ28xHWwYYi4YInpvV1+XpuwiG
WUcNhxPTzMNeN8OoUJBST6ovXLxUnxmF6Y+pqygIMmyT9K5jNe2DVLV8wGV+7tvL
ribw70e7ess8E48DxQl5Cp1q2mBcbhELDxo8ir7fACVYmwA+Q5beUwEK8N6BmR14
Zzw8kw0qRdRwORju4vJea/MF5Ql5SBi3cyLdp6G5A4xnOliQCaQNgQAYY/Ijghl+
5UHARNbXne5bl22k1+F2gfZoGoW1VxdYAayCdYsYTI38HvcZXxvT6subXDbDagnz
e8yHMaBP3vFGXl/8k8rU+ZLwb833/l/zs0sOdmdmJf1xeOEc+RXFm0srPBoNsoZN
jnrPMBfg0buFDP2aAGwxvLoP5Aa3foM48Tt4toxkBlA87wlgZbbiAwsX3rGIHTaW
azpNFF7k1CwtWlzJ2jWjs9JzImflHUEUCUMn1KixI3siZeblHyjo7n98l/pJ58gh
gTevBoo0hc/q29+lc7YlTGSrY5Avtx5xJpTb4kxkNu7iEtSHEtoO+HcGAaEc7aWk
wpwrhL3E+tXpQyHDLkSbCem2AzTIwlCgtUQL0aRyxw/oCgB/pt1+MJ6KhaAy0jCI
dn5g1oYMK+vnwyxG4jHWsiMbDM0UlpF7obquLbgiVIGyMgcPiEMe4xAL2NZieyyt
PywpYRN5UKC5p1z6QFdvdlonihpDzrVedPj/ZKEfYOfPTin5Kp8K96aAh+rQB8Nq
uAwy0TWIKcMaZRUmxcmcT/+esvJvRyQS2u/VQWuKgvJ3Q/kSB2SbvO4CzxhmtoHE
/Z+FjMLjRcGph9cYeAFr29TQZzC7czjEv8Njz91pyP8tMKk2Q0+e60a+ke96URPZ
1GUtDNAAGaSvT0gNkf4XLPjqniDCqHe5nRPWC6haF2hsah5XovSFtIKuGiOkvHJh
z0RahkLVGygswmtojqyxZkuaSfb2x1edqH+VWtzYxdRgyclVhrzqtMzGqe+A+/bo
e9aFcjY/nQVc1PDmDzkyfA82MhYUfM7J47iQVDkGR/l4TfZAKo0EBIGgENMMQeiI
0XFijeexqLgHnFWc/XWbwmvI6MwthCs6ohrZEv+9CVBhJRGDYW/U0k2IqWxDZVyt
BoKJYXf/utnAPabDpnkZzGnrwJQ5rew+HpmHVcYbUzSchAPfdjsFYLb9wZUIdC30
kK1mM17RJCT5/pAbpjAwXVy7jYuBCfxNr/XqWUxCCc1Xnr2GmMx4itTXhod+M2vf
BdHH7eerjmgZXM/Pas1wPBEphqoGVtLtlnII3HfJq3F0jlonJMqX7Uo4NUpaMENT
LJCxc+loMK0aNg0/kjDtkyAgvJ14rtlBSbmYLWAoRiipAptqfbt/Ba5BPGJFzBhq
nmpd1+SgjCmKz9dLpJBtorw0CGmiUgopwqBxPVJBCJ3+m1CFsi50cAH/gA2ZA46i
pxRVAnmcmsnk9hs6ySxg96K5p5EI1HGzIllfsLR0uICwzkE9VxWvvcgxEjt7P7b6
sO8jooX/FY3AZCbmn8lskVa4bbrajTfrFpnVQCORqUmzyjMG6JncVEas5rIx0PPe
edeQ9k5eoIXRsh4c2Q3GSC1IAMV+sYPPpElIXaLiZ+awJoURBNnrej8eplMOjr/S
h9LkHZnS42Wkuy9gVnHfXtqd83gduGoRMsoejyfOZu831+NQh2QJXjbO4SD27AzC
DxJ9eGtnKKbGjzX/B2sYZZjZKGwaE26zh68xjydrTMFhjnf9EbNbKQeCVlJtFLIB
CKRj3dZQ6k2aOJU+Gp+NH1cHzCpeTXs+0jg8/p85PQnyT8ei6zUXW/VdVJZ+8k6c
32dI25rfYKGrmidH3/r129uMjBR+KKMrdnkmQtK7bCP/vtFW2/uNJpfBgdSbSC8B
DUZmzQZ/vhsRLSulXprGqz/7SW5hs3YIrvOrFqmZVAdYbq7W3zxEiOoff0cFeg2w
EtQKambweZCBPng5j4tgKSHgDMncyVbryi64OhFSptBDKxAbY/3ezOIYXajs5Xxr
poS6m+QY2bVEK8CC5KVTsAaFt/L9BK5MWu5fv9aKbizSk0dqmmdKc/+femhcY02A
iRWsAr9gkCk7UEpWKjsU/9nrofAvggPi1qejVopt9Cf0ciRoQxHGH3rFjuPvZWa3
XXTIhKQ/mWODx86dm8i5cy4cn+EslREO4cA374SfTRpFU+AwpSpCo8ziTvLSuv3x
4+jkcCgVLJrsWpSoRtoV1zFLBB0RSiXupPsskrfHchELpPYHXi9jvnuP4fgwQkiS
OuPO4qrSN911RC8Y9XAMvvIe/ThDCRjJsdvNZ0ppC4QyrPSMnf9RwJTKmMKvprjK
dUEIs4hGHIX0bK+ldov61Jva/Kbuu4MvMjUg9O5CTSFZiBXXb6uLSZJapgn5PLkP
tyytoGcv9j8ePo2gff+M/5yzXaVnTwBQ5ohRtA0gG5VDbiREhQdsw37mwQDqxqz7
vL8YIOBXDLt/Cq/ym7E/p4BhdVXJvVFwgLPRGsNz5HWkMtX7u1aODOPybKmgI3kP
mSCQsZmRkAFcPr8qHZaGIPA4ulz8ee2FcFibjjmaght1vxEUgQoNQ8OkVQPPDT/3
9Q3fY5sCqKg5ZCbU7JOqpajZDeP+hhdxVvNPI33N5QwnZ3dEp6tpgFRc2cuFggrL
AnqRQrOpg6kl11wPDpOgVyjy3DZH/JYK+qWq51BT0vAaVF2uickrM1LsXHrfKy6z
k5mRH0KvTsuecU+CEqZu/z4Ch7J47VWKH4N6uWLVVsXv9x2bh7+7T6LKa9QFq2VH
XtDLl5Adh0pDHKrSf4rsi3xJeimCiyc5ON2OGjE8JiglDFWMFY2ip9nqbEpZMUVc
sXHgTJIipfqGZcX1hnIpM1BiG1QBqtQsAPG1eZk2Dx5Zbwy171UySAgkEmytEirY
qS9dEdTCRkz0Wya83Qj5PP+YQBPAZnckxauuEziX093Gg5A4G3yLONgNhWD5I9ZD
ipSx0+JraaSjIW8pXu9XW3aAa6aH/6DdRkaB4C2XppfEXnubWSTis7V+XTMkp/5O
gQ83xqnCiwrBu168rw+eiTay4r8uODlyD3PMcamkyv8Clg/Vrlbu8hKWoiruzoaW
RRRaMNfBF2imGupRA8vDi5klagPHoQ7Ut2sJgmGP3CgdgH79koVEkLWI5gOm1lxN
4jT88q3UMEuMgs4JmndVAwjejDd9HfDqkD/76GRaClR4rMra7n8SX/ed7Dx9V3du
m6KJw244w66eKUnhBL9gLAuuyR4yh9azfQnkXuRpPG3U3nCqsjQHNuajxbalowHQ
f5jk4tBM0JDKTG6MuQBONMPGHTCV1w/WSOKb1zWr8TAWqY9R2xt/w8hijXFJm4X9
CKeYLU8lq9GSSOcRXW2GFuSidDq8dgLZuTEXanFMd+bos+k4mB1oxtJ4xbu5cOqC
9vo9tbgFqstaakW++1dDUAiUwcyOoUtkcTbw4kKCiLBz5MhGGqItnJ0RD639B/go
Ke7CBSdfCEkgFQj2KvYctg1W64jBOtOEZMs198yLB8qW7SO1Q1sjr4vBCIU04k2c
HovI9BqKT1W8Fv9Ijy/qfl9pPRxDyX8SzGJpBW/kuo/oteW/QgWT8QtLf1WNxL3U
ao0J5jqneTzCVviu6u9vxJg/iVrHoWreXa1NR/xkkxX4hw+aUkVmxONJ9TERJTVy
Ydx4JD3SUEY666jK55LDznEsrd0cMdh1f9/iBxebw+EaS8qH0UxZ/QUPd4ldQlZu
fLFYPI1H6RjO/GqTQgpXAAjjcRFD2zQpgvHt6YLBxanGQRaT7yMZngIwEnYN2KIV
6PUl7heIylirvFOpkNbR+SI+VCYeu2cC/2DNxwdpQZXSxPb6voq46XjUKo/t6CBJ
UATk4NLbr5I2ddQc8l4u8nNt6moig0k67dzJJSAtNm+BaPRl17AWZ9qSmzFMkwcl
9UPGAUR+1ToYl2SWeKcUMFIZvqt3WE0ZaEKhRfSHo9nh5CMsD4Tw7V/ytYFvNIV0
cu0no1IoQljHcJzPXUUqCgiPwQjG7yz3WUC1MEbvgmCegjzzMoFwSYAc0AuaneQj
biGCMBK1ZEEfFHyDwMK0IFcl5erFVNnEUKpHKkEF7BQScEpeuuR7iW1M1GpzLF3o
2wxcdUdhydZC4BAO/ZmN7VntxSK+ZqEmlw7UagJXkB+0rBEXhSo6BIFaw+loKynQ
3JoQ0rCpkvZ9jGN4N3ASAgi/wbscrLtT9esD2nALbJyBkzJ2G48JmucDmAKLj9y1
kJMTYdOpCUWSlDGdo/Wv6ckg5A+S9VhFjYqnsMKybYMUuvK77zBQFpHS+7MqAT17
oMC097bztl7AEl2xwFdxpGkSanwVjnwGANwQUSQ7GPY0cPlcpoSlAZRtOWrd/uy8
Ve46Ke4KPOLwqHwRsFdeU6AqxB2FgrvCnCrUv9TSaKA5JBfPoKJpj1Ej95W3IaWm
GZOEPXG1lQroE5gyFvjIr0M+cKH0YlvoIaF86nvcfS36u2J+v2+tOdK5eFWgCKKy
MipQ0QaA8qUNk6RgGNtyMY140wpu6xpwrQnNKEBj2uV0S+fGtYaPyOc9pLEpnI6b
iq3PdBrenKsXGcvyGx0suxWvjhqr1xIoL1+aNcKkntUI/i8dwfTzLQhgaYq4etyZ
1f561LR6rfmQgwIAOh67ltMbq5LYW1x3n73riPcoIWOuciC2sW5RtGc3ZEjvF0kB
rlLvJ1ArYZO62VncVEDrOAuoAhqkMfIYYk0kteXuttM0O2hJ2bwww9/0Wp8gcx9N
5wjcYGCBe7sSEwtPgeZEis53l2Dnb1Fs8wg7IQ5LOhalhAojkmHYkx8QHrdodJmi
XzZ/+fO8doRa2y5j5lmc85T3a3KoPClPfMwkRJtlx+eA0a1ECAeKLyVAo5yt1qho
bU6DSm8WCgfVvNM6Ep2NW2/KapeKlTRh9X2HPgxUiwHXDqHLKC1YPms+ed0iNOPF
Kz/5sRgKPL0/5PQhvc9cWYXT3rWhfV0ofx2vwcM+kCFtWQGcLBCEOA1/vHJqoSdJ
GhaFIii71f5kuyBEkqG8IiXgshcTcP6J5Dynifj2wMCcL2fGls91yoCEDEm6X1HT
rOc3waht6y8hncMdLlK/yJvdr3l7PahT5uOB2qLvp74bbrhnOOp79sf7Q0dOnFum
gjSg73eXpy8mWkyR84rs2t+sDmfl+tpY/dF7p+NSIXnM250ChIGpo72HInY44nPo
jRzs8Py0h/Aj3DwxsvYST9V9ycR10gUCJrStKeweece4sVbH0bdn0VhVRv08E8/h
4bgWMxMCE6YMcyko4Xp4dNJv/J01W1A6jyXMbRdlISAirqsG2u8+JtEnvUWeEQB+
GB1XaRkFGXBri63u+dM/c/HdWQ7BOAXpEdqgUcm+lRJopansGCUjjTbkrWjmX1vw
5v/8qIh9gzeajhp5QpLRk1ibbrpPzKltKFUvLPNLgt+Kbe8kaqeScVAJG9xrJD9N
pwW15or6JnEMcATqPyiErQcm1Hcy0rFRGDO7LnVSaMWs7QKIG9nONOD2J0AJ7Cnl
3jErAzKhBsXpK7pqnvbNBQmHxM/CBawIO4bN/2oJzBvg05KVtH77nqTiACz23ZbC
Mvsu4b/iIhxz7G2gHH4TzIgNwx8z8584kmue1CxZYnHKxYKipJTbcNeN5jySselU
ek8wEKZBchgitNYkg6qxOZrtvKG9ZTV6WQL68P3Q6dAZfm/6yn7ZZOjWjT55ofKg
YIF90QNvdPd0HQ2EN7WMNq9aKZGa8VNuzphT5e7dnJc1FJGP1/YFOyPEc7hU7As9
em6inVesxNI6Q1Sfva5sphl4CqLaX0MpeXY12E6CPU++pOl/PkIXLLLbSeSAvEi7
XwbX4OPj8qsC924LWMlMzoUFEai6za9AoHlguZBjaMSxFayAcCMQzbFQ2RD1gbhu
pRuxPJUET40+Zd/Za/kFlLbExODNQDzjSmGZEo5rYr/VNvEt0tQ6mZDWB2CjIG4d
fBRS89ZUiboW28SU3z4IfTZSohjlRJmAiX2CS24DsjSpwyTVT2uYH4kr36QAB2uA
Obfypb7qD49a3PGDjyFHRYPwaGScGdb5uGIvnrXHT2r5oa+Tjh6kYuY9SdA8q8TA
D//SUqQ0futkkdRIRXMPF09vm+GhiNHjrfpE3puWca03gvycbNPcMh+1C1ClNc2d
xUp28Q+qU2Ho5RRyk1xt4Dw5DCnB231JAAmig9+IlyRx2IRCCx7VDCXua8odQbZG
BSpYSNJ3kMd2Cw2sifnAgri9YU66IL8EKcW7v++lL+sTzCEWkWHTQ9SJ8XC9+p93
Oi/c2sfcSHJ1QK1mMS96y1enLvQs1sx5YS7gGhtCbKG96b/n01yPiOxRJZ4OMM/a
MluPy2KGHfqMSGpgB3UlqV6ITI4QiQ7R+3Vf7+j5C0Y5LAhUwhe4eRaQFXcI7LSO
qQ3GlkFPRtQJqNudfMthelz+lcwJgbH7RJynaj41g7yE3buKowZ5WKwqaVXtFwXO
gpIi59k7390bxIgLSF8cOhF8bjAG/h/x3mrfx7zu7hMAYn3V4d+faf9sN0+PIKW/
V4ABmid8G/aHi4wHFryC1hbjp1egSTYkS/wZHH1t0yOTU98sVbV0/m/BCFLFKRJX
wJAl5kIeA/TVj8cIlm3Yc7ukyvlKfpsyfqAkdA9oFijCwBXGeUYOZjebmSBzN2fb
+jELkqFp+5vb2nl4wCl8vHS97jywHkIF0CrEafqFBoxUIHJ5vIL4ZBV8EEr+NVkY
0zD4ULrB/+ehCDc8Yvr3fixAypOwhlDH5IQVWiFT1qxGLJEc6lT9LfoE4DbqZjSz
J54FosmCVgfwEvgnOg4Md9Zx3bCJxmISmoN1TdCRZFn9TE9GCV5vVR391Iy7YdG8
m7xww7PkVS34VZONyHYi5g03pv0kXnzuUT5RMWgZCefmVfib6y5VcumRUP8Wkh2U
Goabuzzma6wtYYjshQQ5SPFndWsmM0GIWLhRrLo/0KlYH3Il/BynQTQPMEqLncJ8
C3pXsFFDOQF1b4aC7444p+xxUn9xBou1UmuQEJEuJI+VzeJC4PxzfF0JLHb04S3k
EZziL0Hw8dPS7Ky3wHQtocmd/Jf99bWvubJAFfX85F1PFFRBN1ywJQQH9eSGEr46
eXmIMnZxL7w+enYhMwz+BVnNOwU5latbeo0blNqJ8DydpHpT2SN+rSKYSPfoWywK
/DGDqzlUt4b62ckid7rwGBixbob/euDG6BELSRgvq2fjTwPNGdXTIiQw6lMclVkX
VAOaG0xfOQn7/pvvbRUb+VzloUMjfK0tBvl+1wsePrwyqx2EMFuB+6utRTyIPBGc
v4NnBbJjrxaFy9xOt8aLeCX2m2vIWrVyrcMRmgt6SzYH5yjbpm3IYvKd17XGQN6H
6izjA9gs6qEvghevWkCd3A7RsaC6kjGeIBbky+KAh3oU/p7trw2Xi5HtiqPFrP2y
lhRBJA/fvSDSR2k7AgHu2LbNWc2UAn1+TpCf27kjw886DXKHyjU8tSec0ru/I//I
bxGKMTPTzXlzFoMvs6dEwIaNh2yG2aV2uZEkJY7/eBZ6sDWUlbqQWkOXxO1KAd+h
QmyIpVXm3th5B//AZ2plzdFW2bSWOCCQZb3uz+HBz6G5bwV2RLgnA92U+szwtV8G
OROseFJFlbbx0wVCPD6JHNmF4p0vAJEGcwm+LDxzK7rblNQ7qhDAslbtCgcXxjV4
YlojXnYrMCGDyzabYDktvaaTbnlCLQ/E/hLZRT370lwAXpbCseuPj8ZdSqvktjQR
yocPgMKAenIWa0sk6KEpNr5XQnRVWpI3fFtFBKSbBGr7pIv7OyEhVllXdqzPdm85
rPOzptBPiXywgKjE+1+696dARidQhQJVoVlmDqUyYLlYuXwn3hXelYYjioFkyMYV
XYCbj/x3dC8eEeUfaAJNzZqF1tton9+xt8tKaM7luNIGM++khP2Ouxy8s73Fkg2l
A9rgZrlSG8v1LVf8z00a08sdeIkSepytM6d+gOATT7OfbjhGVs5Uo53QOy96QHT9
NEtIc2OBA3+Y3LTitT0HoZc9i62rmxACgyOu9LRPpaWdtjICkUZVoT+nJX05AJox
qqCue9ZVZ2TwvjuT2htnbyiBuCpkQ3Hz1BTbQB+klhBeoKEqF3wh7RGdeYOOA6CW
8eqcZoNn8JEzX+xJ/KkVLP0ZT0kWTynGXEdYAXOkoYjMaE1XTXECzzGnHFver52H
LeLInOELzpDo0K++VvBWf/K6tdFWuufoAh4V1/OAsk+T6YRchp1Jm7l/zlZokcGN
8Cx3/52IV8BB8LqFeLmE2d+dAX0pzA/uOOiCr5c5BoJDeyFcjMKi027gEWL7gWo8
d7mTXDBia+IgZ1cid2SPN/Tp6Yrw3wadaKsTZX61QYXPtwsq0+EBWyKXULg8Br5b
d/zl69VnhiVEuduv1t7hbV4y9g0i0Jq8MBzdu7y3vSBfSvUVHSHBintwDgOfr/H1
XUjH5K9JwC3v/tSnh120PKW76NQ8dRKsZdw9kDg3pWSe987r+jmN/j4PNd3H0Tqc
2GCgjCk+Zp2qRZuN3bS8/OlXHaBle1uCSgpa4jc6FYSf4zuSP7JlQ15WzYDawMjK
4pnjx5pkJ+pbqpEXcvRFhjeakYuBZqmBjiS0qiTSvU6zg8qWY3K+zR8l4laabcBm
Yt40l11gN0AIcQQDnlrMK/hpVf1Uw7rzSCsBy4hh9BH/dVAsk6LOFabyEtHv3XkS
9BajtylFWQ/+7cbjZPYN7octArnop3eq3BrdYFAPIGpMenb+4Ncd9OvRaI/OJR4F
5+4zFso7u9RhDfyryMZ8nYEHr4F/y0m1HgnaqWUfbvJg8N3sY7MhvxrFXGFcn0gc
Aq21ji34l7xBLgDTUnkbL157tMPyST8O9Y/5VAXaSY0xfJeVTOTcpBu+jQUw4uh3
2SEWhgfo2rIj54zf8CuuBTjlSIn8fRhjDV12W5dtOtk8TD8qS8UgjY+GkBMrbLcI
dEjyvYlipByOfoyJIe+HUE3jxXWhEmviT0R9gQ6/jPwhNDD7BV433cg5rgLNlwru
zZc2bbsP8w4H2vLyi23k9HUmFvmD3RwfD/7z5jurznz/Z0eub2elHXnV3tt6on+P
npEASQmkvdS7vS/qZDpnh8AL+czIQDmbp08jCYtn1nJvFdoypevWuSWx1X4pT7CH
RegmSHBzkRjifEW8xbo63/6CRyyK4zPbNACBa7VCTLJXe3EN9JY2SdTwfFG0lFKp
lYtqXcX7yGmU9fT5TOM6dfH/Dn8TEZ9Z2aWlOMv2Btgi0JvczpPTTz38QhV4I+Dh
UF+ejuRUo0SagpaLK/AZAHirZvbdNGE1DfyX8hOCe7p6XUgkbxxsTMC1sC+Cv1Nd
Mn915BBSckZdlUeT+cJpmg1524I4i7Ms3nkeDyIg+yVCWaFXs5BuXkmxwhoQ4wA+
vxXirKYGsvS2NNuuDHj4onVJ6jrDys8JWTF7ZYpB242BJJSqc4KCsWzX3oPyo5cm
vprZ19g1a6tXg4PfJsp1blfA849rb0NeK/d81CgJKluB8KSQwYKq1haeK34vctfe
7wPCyyqznCAkO+wsgVy8d1lEbXrW869R9X2yn+fkrgl1euD3niVsjGhx6zUoKYfF
Q/NLCBijmSdPU5jKorPzprD+/m+yeJwMr5RzX5cvqYb6o/4TVwRd6b+esmNwbnGt
APJdY+RDeC54xyflQ73qaaGVe23YbvO4NJilLJ4QvSqwaqui/kxj4zvzmGx3cspA
0E7qPXmpbWhs2dcvaHHxqn9O9qzkHXyvvlPhyruQKo59X4stY5XPNgNnk1TlAbnk
vLsgMzi2QoqtKLVRHIEZl+PlIy9+J4tXhxWR4x3+9+1G7xd+gPGubPpHT6YlAQs6
ymkq9iFHDlNKm313C6cH6+xIgZglnVWVPpq5i5835ddTP4Nxc6yBl36LoClwzBMg
fyBY0NM/QNi6LPTYagJT7O3URWXzKDc69iqUS/c6CT1xPB365e94VeKoWVRaon9q
XUb1PqTRPqYG63Ook1LFdv6yOmkD+ssUrfWMxpdZe18/YjlaUpeoG4kY+OcmeXOY
D+8N9dROeW8+aZUP/UvWvB6EqvfRR6mqY2V3XVjykvPtLhQ9Rv0tgBF4qznuuvQg
12cI1c8vshgfSSbxe1bgAt3Xs5h3VmSB2aNtSF94vC/yl1xdQKnuE3i4h8ONIa1u
GCmy691fW0MViiPCh9B73qwpO4ZK4SfO423NV/ogDgkIwrewsHxzti54+5nYTOIq
e85Gthxk3KaSNigJkvqHpFuuS+5HJFAn37sRADQW35/EE5xg91T7zl/p8YChZdtU
xELnH12tf/PSgzEMAx8hIgVjE8+S2DrLnhkwu89HqvYvQ13ue7PNtynQkzv5I+Au
2Fk/TM8Ops0yjK1S/x6qS3Ye+7c1NhF1GICSTtLPknGvVTSp9Chjr5sbfSLuXqp8
pXD8I9881SGi41PkeL9mDWQulqEdTOkJizNXsYN52/t3KZSxOZexnD6oEocKr2ub
WjeEJYqpnBp+nYeukXI3DuBMpE7l+g9+GVKyhC7wj8UKFqGDc/sUozsoyZz0WirE
T/3/vaja+vvLP6etyLZNq/j34MxGpo1gzAK4KkxKRE8+r88o6z2c2hr7HlcXVz9T
R90rq6ZuGI2tzRn+9wtySTKnnQLFZeEp53edLhXzZnVoUCPr9vG15uhQTR5NB19H
9NGJdqGb7CU7oE0PblHpkXYmX5gnbmpcC4tHshcUyabNM0Rf+110gKf/iODOiIdH
ncfa0dO66cbU1FWOJ1+JO6hYH4eE2SpYBuUrmjV/ux+SsIKbjJC9YXSVASZZUPmu
Xv69Tvaas6NwqsbHTejHaFkzz2YXlCEvbboGzY8nEoyisM/Xx5U6YnjHFy2vI8Gd
aYoWOIg+dLsNYr7gyEGeLZlfkTsinvn6jXDWl1GsoOfYyX6J5OGoGtV4aPuDjnpa
bFF5U71gVPHHpQ3IUGL+/nJiNgCD6IXueqy4Svhnq1tFuPKRurv/u5+gJJ+IKJpn
6nz710xKz8GKBF7lN307Z8zxcMk2C0sTps6ir/NikSdUoBaSIE32RHU2byTiQK3i
F/nnYtbvHOh38auII2F4o6eA8sC2E6Xoa1UdRoqZeDeTgbGNDbEi5ym/AA5u+wsu
cPQsPiX7bDg18VpAqX7A1Mh3Tb4us7Vx7pr9gbYnaAZzQumLvFcXHOFrxCukyRpz
u8Fj+skIEOeRHgNf932Q7c5BhqlHjDS5CHbB1RlHlOfNSbF+lyEgT5fexjfN1ZOX
V9m6eDMZgQ+fXK1Z5ps3hAgMCxb77J5+j3+eu9rP8kznp+QEwSD5b+mnWf8PjWDa
VOOD65sujPc76Y8jRgkoqC5LsjAQjgcnft9KWW0S+9iLhVFWVPRhmB8zirWQcbXa
pmWKt7E/u8m0pM6wJRKm0yUmUdRiXwsl/qXbNk7Kq2CsWIDQ1ObQ0nbXu4J3tKMo
5anLbNGAcxWZc8gMTX2/+GwmiV4J4OXbZphWJuqd8srkpE2l6eNAX4ybEbI14oqe
If0SJBdZxW5XrcGQEzD8HtVVkEFUJ9qA3AYkRhUxBwpc/CEyGiPFLxK+gN+LJb4V
Wvq/kaQ07GDa7WkNY7K9FlD0GDWUiavVSMJ4KOsx5PURET/Xdyon53WL/ktrwCya
BYuOQYAzC04zTuz9hvAnSz6KdMVigPntT7/H3eIqnvcUfxQliRqEvbAp1B9k0zfF
8Qjb9DoE6pdUA1h34yoD7mHYooDHc7zCIn+3J3v/qhZ5lLKqnOeQ9NQs/V6hAU4+
pMVmxwaB+p12E33zyFlRDZX0hxYk3/wtgmj/ErENRZdSS7NGfRxmb5Q0/eVKooAT
76DJKpgyJQenyVgFaHbamMcBrwz37sdtB6u28GcT8GluT9fecmlG2OrFxJh/884C
9uGiX4nyxryQbpxNKzUabae2sp1TCgclAlMfPdpcsAO/b4OYrTeFNwVRAlnDoDkB
0cC/jpr+bT2DJadjs30lc1XOFFdtKSiqJHuvnYJ1qSyEzn7cmXHL+D3yoO/IOXig
DD+zEqtgZj/OzGwusFiQYJ6VnepLjuaNVemH9BD+IBnFinp0L0/7ylDKD8/cK/5c
pUBy5kNsCLdjOWW7y5u+pqIRR4OqV0kXr25GrRQSH+QjDJlZJQANSFngNoUOmA9Y
pUGN7ENV5YYRZbNGzuRoaSGiJu/QEa5XbsZ98iz4fIZ7hRilaP6+NrLZjpVbc8tI
8LItShZb25xz7aRGA84pMHQzk/N5inNMyk8q8W9n/VVTTAcSoxGZ5D90rLeH4dOY
dLEZzBXizQ4UZGMHRh+fZ75sh0KM9uKwq8q71EiIGG3jtZi5wR/pLDlpf9tHF/Rv
gpF/juXDtOce5bnHpYVXI44R+Pw0r/SltLW54BfAgvur/GEF/VpCctmAFErcWcpo
XjqemnTNZ78wyqCPYlPxOvhkDD3KNlScmlsVPkgdtUlXZMDqymbbTizXt3Mthxc9
XAqugXtUPK3XRBfLVsGhiPiPwb7zIB7nd8Aw461kMoFcb/vP7WxPaCf/ZdrB/Bls
waj2mczr0SylZDrTTiM9OaoPSr2pycVKVBk4gRmBBfeWMwgZYY5I/juJK9WnVhoo
9xahjaKc+n7gocp3YYT8ya2YyIrGT+BBFhsLKTphuCeL9kMk30whc0LjG2aXHaWG
nZJtN8NUqAi5tR2ipY6GYaprsVBTWCgDFan8SjcFNyEWyyihFYYeLjdZQkTYmiRs
hCyjW6zGnRcSMQ3aC4mWHEMKVfSWYS2Og4iXkUHC3Y/LXgmWC5hmMa9AB5fmRlzS
1uqFu7amB8XbDJXh8b9sV109YAEThMknx64dxKy3fWK/R2mF9lBNPAUvZ1BFDfkc
8hIFaBQT8YwGUp0A6wfUxzLN3BArj+KFh7fD7qveHgk66gsLAZ3BaRXi5cboWubV
5f/vdajs5+wSr6Fcwu0sBdyZhGQ4UrZ44Sp22ShNqfUwGZeA8zaVrEMRowKgzw+i
ukEks0zor7gWI2VNMbi/d3FwM+a8v4XJOGZ6GLEFTWdhj555Ie0P0SFGOu6q8+eY
otWWm/lPbt+lGWMbQGbBK605NC9mkcfzLtcTwKi8VEpLnT4aS+mm3Zdb16zNLBxJ
nzMsuSH1VLoJxS5MaB+2h0dO17EDfaxZC8H3lewPwsMG62k5dN/rFQGRDyEHuLea
oz04QZLBhx3EA11eau5t65cI9qKhphJC3WoWK/k6Cps6qKE+OqqOokT8co7UaTRT
UnSwzXi9LLg89BINgJzK6NAhGNEWO+RxvYvQj0fFpEg93Fm4qdES5LZOsRWZVf7u
JAjWQTnpyZ0mw/JGAbCH3rzfnjEIB0dRW8AjVCzQIt/C8CZl8+IZu+Wah8GQVRjD
A4ZpZ1dN+P80bfi/G+qpgsJM+2hknEuHAeQ7oPIpM9+3gG4wuuy0LDIL+TW4K4AL
AAkbxjWoIswmAR3aizCcOCvd4s4mERKz9Hf+1+mvvH5YwqfI1aKm6asWORPGSkO1
+9gey/ciZ768k4Uiow8Q99nHGMm4q3waI6VW5SceICOhkvrV9+9vuDmK2soY3L33
17Z2c0WuXiaGUZ9rekHnjqLc+JibTx3216Qh9LOI4WzAWiqF6cSC6XGnsEhi1Omu
p+K93ZmN3q8+ymX4imZq59woghUP90bhUwNYMDLrYJE3jg/ee8yF5btE/BPim/d3
/BorSvhu30eFfy4gNVdleI4MqDspq5jbhQ0C/DHC4yRMcSgHpiPq7bmCKHg8bR0U
pYNOVZD2BICNqt6s6ZOiIkpky9JrNJqw2AMMn0nQ7Tvg32aHe2r/6Ttg4WG8qrlK
O2O2OSDN2W1KG/kqrGLQVROLVGWUKRKUR2+7KfBFVGuHYK3qwAM0P7lTFxtZELiC
PDlMJKwgMRzlO2195vlFKNKalmLuRCrkHwaEqd7okkXA28lNUpNDkc9iJEIH9sXI
RFU7qNdoDv9nYgTmNQium3mC3IcjcYS1vxUwaALOdxs0+U70Ly12JuwLTgUN97Ok
XDVd8L98u1lv3M9PFlghxGGH/cdgzZdd2KmPwb527WlelFsYY6FKK+vK3A6MlPzY
Y7oBSmtmKxfpGzTQyHrmBtyAv7QYHE8xlUl+rhq2+iUOw1mrmJ9P6HhZeXoVBHKN
p1hYoA7X8yboBcNjLlMZyjWFSrWEI2c9KidTlFYJJjusF/HbIDjGrjz+fxWWj2yO
8mQKrvMBBp8z16DHvewD/QGtDC3SlSv9wjK7lcNbTP6TFtpCaL2uZq2JXgKVutNz
CgOfQebofkHsv0IotgYOe37DwrDyHJmQGdRAFs2BbowH6wXri8+fsl0/rDk6BQwk
9BK6Fzqe8Zq3vXml90J6mNmHfSgpXmGM4zVOB9h2cwVkogbdopDiA+nlnK0MRDXH
VAnZ4cjtDgwTiKwYLDuB2q3tXN77vvLrmjkwfjb55fMLux9O9gDa9v4582zKXNLr
j1kCekRJal8XpGPhybIMmWBTsvQv2waZjTvxjkGIxZLpJLXBGicy96RS1ypLeC1a
ENAIHkL4Jh8PRhmoOlR4JEJg06/2yIfhMr9po7UW8il1bpXQwvWQIzLiuewPiMK+
1BSIyup+zekEUOQUyj+5/o/nV04feR0bPPPtveUw5MXxZYdOh+6iclvXFcT1nJBR
mN4pJvSS7mQX4bmcFm4HFEH4o/B/ig/Kd0tZWNQa6boerxDzhoH3LZakCktp3CkU
VjQtyCgzfWysznAjXa7EDLC7SU9szdxGpMXKBNeFbRneI3nT8Xkfdpn5FoZCDyhH
KymW+AFcfFZVEVbTkpAZgo2BjWdakFkBEz9Di8zbIQXaNXcpF1Lv8c8n46XWTzBu
/rVd8ftmny0tSpcUJQNBbo+DUkS1jWMDr71r0rV1Rh5QYRRWGuoL2BD9nSI+Bpn9
u8rbG87MKQ7jWJVACpKy/N+MjMVs6PSReE5F/hwcv4Kz9bERkFBo5LlsEalfJUyx
sNuNftYrZ7CFyS/XqhjF2n64zacJZT2I2NdOC2kuHIygFAaNeoTXc65QmJPRQ/Iy
l9h9nT0yVJ4pGcJT918f7qJKtWzi2Uq2bjWYsjWb/k70Mu3YS7Kr5Q2T0puaOvi9
LC+qUmzT5/oYjkQFvcnMZvb0l3dHEBjYu6CGQn5WuF+hJdAEFqIiQVrWqySvzqVf
/t92Uo/aexsc3hTct3RlGUtwRDfv5Y4rq8DljrUDaaPb5FCEXxOOXZ5O2J0fkwbN
8/VAwawBbITpT41jBlCDW1obx8Vk4YPklSsOeAMNeqY4RSFrRMdsCEGUQrkuPEIA
pc7fv6W3hsJ24J8eB0/+syu3A6DXmMgnk8myRi8WXwulwr29/Q5KoCScCpS52tIe
YUon8sQBibmpTOIFqHaxrv8QP8kfpSHosBLbOr9jW+kI2DAYZUihxFHK/ZpacWjb
KTN5XyDhh0GLLK34cWUEgIA8cx4Gd9LQz3JkKBZwV8p8gavY0Nqw4DySEoIriusp
/RdzKSr1rowgdM0qCzwV1JN3FaXMNOJ7y/2jzmZrw+BntTE2Hae5OzaBRBrZLKW/
RiQzLLTMEjJy0yB8hl17Y2g5gCh6WfZFPeXBe/vDyz6fb5jATtpzGrSI3fH7IdsE
nnhQqQ+TKTKBPJEpTXUBhvc5vywbhzBn7YHgsFykYpg6ydjg+3Q3FSRiD88vH6Sz
2HC1McUXWm8H+SJiM++HCogD/gr7IwPjOvA61nlYIbJihrJBZBcgdmtHVee+I+Vt
30EkV5QnlCIsZNv6vv6beN7x+A5f2qRP7GqasBLUye8zS0mAWb1y1FlXCAc2Q6s5
m6FTqxx5Z5fCOgLxYWXusV2LWZmYaFWNIsRmBiuGPWbVGZEpVSF6YIMI3opQ2rSM
YWcY5e2ONVr10zBP8F+3LAeW5JxGaJtpdLmaqh4i5yRy9wkLbi1PWG4cIKlgJP2t
ut8hV7fkBrSP4HYkwiqnoytcsaQqmq65pyRM5q5Qc2bZ37craFutFLUNCjjKfVaR
EHTjhuidl1EdT7CTgixqu/30PSy/Sz2K/omzx0ZJy9BKz0rxMnYV0sXyrdpgrAzU
U93RaH+E+Du5y1X+7J/cfykUph1HOARs7FwiRg1GNfgPLdfK8e8+IQ5Po/0+sigP
Ss8LQymSoipIrgq+4EvV1vXMftQO/4tUwhBZYM3J4osffwzehXlGnoBeu7J4qCj8
QW5CZc17F0twOfA/ZFndq8EWnyI89t0PlbZNMuUYAo/a0BYPzrmSFv9Qa4dItwWx
7gsj7kfcVErl3R0UI3VY6tMotPIyy8dpZdOb5RR5Q86Afh+NjedmdqSSAY741pnT
E0yOQ3AY7LuoPIT5XHEJhIl6y37WjcoOw1SHe3LMjm6CZXWeq2T6DBIGJWdUwNIe
zOkS/trPfuumllu+r5lS5NP4HUjq+u3Mzqja5uvQW5Ylc8TTfaKefy+0PZlofD52
j/7KcFB9cmFDsQC5r9bz0PwM72E+5Abek7ygvaeMULtoDoMdTNd3w+DL32/BG7m2
07YAZW0TdNeOTi4QaI7BHu0i50UVkIrkLltzc9A+EsbCAUkfVCO2rF1SlCxJQ27N
bE8rejXyVf69ueHnkIJWW8SbGmYRVtwZFc17c0d284ySAMvRjxNHxh/U3Kl+ao60
KIVz6mvHQ/8q3jUdDKaXGBwZrZ0JQMmvZMb4TYj+KMviBTtnl2hRnZIrR11gidRI
/3AJLImZbzRJZQ6B69etVul9cWu37lT+rncctzD9+tmG/ukx93AYqY5nN7f4wEPa
zLXRBh7cRM0P3Slz90KxgC2FggkVmMenoBN6QiCWh3i5RLQb4+T3p7D6355K1Rbj
hD576h1Zjxe94QNF5xpoo0Ph+mPOiPb9AzITNXxS5p7XsEWiE2KDxB/ZSv4i0ajv
pejUIVLHGmECwtq/+UzA/vfuyGPQTJ3qb602biJY+1ytcnK48r3HZ1vJI2zOnxk7
R6/Ay9Bnoz+XBg6HoEkCfckbmUmUEx6uKg34yBOaGGW/p/OosMu+C+47EouwpXSf
VE2ok7GX+OARRvYzkdwp4Y/f1dam4CjXFmvCAWe7MTNChUFvbZNA3CgJfleoV1JT
o/lVb4U9OECpcoz23MfgcU5nrEodt2tCnmcXpjIp86QYk/Fnc40kdfskpeKzaGt3
h0f2SonGJcFNLTaxjBYnDtrdkPoSwkwpcwwrD6ew/b69XmPpRPjtmAtBbYPdBvfX
T1vjqIpVAT5etiY4nKNfwQ/idyxthJ4wwhhEC7o/eHgoPmD1wYOmSXqDR5TS1lWI
64t6aUDT/1wRjro2teDmCM5l4Vhl6eHvX9U5bukk/XapC1SteLoX12cOBXgvcdgh
fEQSrdJxW/SaK4QuMKnzXxS/wQKAtahUa6JOGjkFKF+5WNkyXBaGCKUkSxTk+gsf
tJPjat640ikkiZCpADjd7w0yoGVwcEd/XB5mE2zWuXdjav+omlSiKjrOnsRTcED8
Tvy2Nm+E7iARKt5yVgrNJlW1EemXmRb55RRyNaW1RhPS3jMYSX09lNaKmP7WU3r0
TnQrsOhBxEhMzZfJ1MkXJIv78xXa6sXusrJOmp/Rli64FNo8/KfKJeDkX8peDjeB
BPkgQ5twWIqIoPL9wxCLqXx9VOkX5WOBkbq0CRPilb8BqppsPti07s1HIHXhgY5r
olELduW2A985YS2f6O0tpdwtkE/pJ0aDK8oB97g+F6CzB2TXkqfdqQtEt01r9cJQ
CUcukcOxMQlvHgqJX88jPlj4hFRwy6/X6ZnjYXJcVL1YToGYXDNDrBSpvHfmu4Ia
L8uecVIzvTdSWloA/4xuhQcQA/MMWEB3FE3U8GfNSzrOkEQ0Uq5FF4wEFDLvvErE
oNWwHPF7rZETv3hhIguaemB0+g9jT2RszbsxHi7kBTX6rd18Qk5JDbHHzEMqPLmX
5hG5F/GK/ewJtvImzU6x+22yIKYs/hFDtMC78KuGKSmCqGfsO5TJJeVk0wno8RQe
f2R2yYwty3/k5FJyaysRneFV6T3xkMRQODPmYzSW6bnrLUCydF+NsAzl4b4GnhwS
koVWNSAQ1ax56zGTHrE7Sshvl3tO5m4VyClTBdZFiJ/7/Mhbxg+fz3z2uJwQYjIS
mOB482eoLwpNuW7QqVDwimyNq2RawbFN++yUpCls3QsSetsM5lFXNh34p4umrdX9
92hjB+VGSxxtPglfej7cvBAO92S5H88VdbwacpwjNI5a778b+q7MfNSwNGCfj3Ds
kUN3nzjvQOB2VNhXa96Dk8mJsBUqnI2K8ZNdnX/XVqHp8xR1fBan/m/Bl7zh9Qv8
+86NXkh0XbFW62w48ZCFGHZxzacFDhQqs77iozKMV8odwqlXPT2uYj3fmF+wNtHm
TbHYkEq1wU7ciXrU53Oq/2ivkcJP15xfKbzDCSov+qPblBiOyU9kM/DfBsHLqgEz
Yvs1n+debsb47XUCHt0J7KWYtxajg/3VCVm847J9Jf0NSea33JoQhB/VyK7WeE5j
iCTO43Qn8pEJG4YU/nKY3GUbMBBsQbTftBf1SXmUQmHuspwK66DblLL7V3xrT4u7
jB7hPGj5hEdTX9fv8CE17ln/v6LoZZub62aTLH3zoD79BC1D0FzSRWmTLosKWtNM
zNqC6afMoGb1J3QQ3Bv3oEJTij5S4d13FIw+VkcP1Ft6Et5cWhcPzOzx0PTZlwqZ
6liJ6NGs7mYvG8f6Lp3LLnJl7jiTiEWZWFJpvDtT9yhZ0aIQvUYexAD/HdHcnfWp
QTAd0q49+NZLza99kfWccXG+RPcqXhjkHMQcR/qgHU0Y4Slt0b1NUwbiKcVM9ae9
jroLYKIj/W8BEZ6Y4tLx+jQ10uQB6SaYtudUwQ0GldkowMtYnIqEICj+JhNyjLiv
juTXF4b7JfhS8IcWdctoE5gPcBzPJZDbR1hldfax//pn7owZ+6g/YZQN05/RLVmT
SFrm2+lgQBPAzd1CJPxYmPZT+3n+dUkzwnTkmEef4cCHoT6z6M2AIi1JGO+1JWiz
whPFXWpomybLlMpCANslDNMGh5N1DWCD6/VLtfZL0Y7lIZs8xLkIcxTcMT4Fxoo5
Y9BM6Di81E6YagmcLiF9rSnjTtpPZPSawcfHS8P2wWd+VIzJxe+kXvll6O5xV1ME
zNkr6vK8f49P/UFAyy3fZjSAybGs4RNR7+KN4E7IOAnbxZroZ0TXEC9dCYF55R31
ubRlpciQ/9SERNva/0o33AmGX3GZgNOFWcKZs6DMvrp+fSwKuZsS+74jMSWFwmE+
DpdhUXCJowYwqRTgTzcpcOl/mMoKWZgA5+OVv9cBwkvsyIwi4o2+YExreCpUiagQ
i32mBsqSzdcqi6h0NatNcbmzjqjtM2K2KQ9Mjc/gUKNXlppHPjmwE1MPYYYr5B/D
GaueLEpcjCoCFzDWogW6BmCLRIm9Wh616B9/MMXPxgV8P/o59mvnB5/I1fhqqBQH
YDwh74U8/DZqy2gJtG2N5y5KBr1+69ajBJyC06iXMQh2oKWy2C5YuVSoQRaFT0Xd
xtunXxa/u1VncdFbCy909K8SZEbkqGWLc3WXtFw1X5oRasd8bfHUCrlGuuNozoPE
xAikhobomfjNrFQ27TCGeSflSV4Memaokop0kzZYL951x3xu2IvW8I7+hln6Cggo
xnoNpgN0LH44URnWAx8p1+WxByypoIF1QzgYK087DEXPjMTr4uEMK4NoXDHj1iaM
3269T9G0tNya0y0Kw0Y1mQQ9RZbLiQySpmdZaYzVfe+qnNTZn32KLyHRH75cTkNC
ILekxHcPD0WIOWGbCGRI4yawL6bKp7oTyPKb8nz3leIC+E/iwsfeBVM4IKEoM2lv
FSUUzSgX9D1M1YV3CbVDJVMhz4pEPd80j9chM9KCYYp1bYFiv7M4zWsVE79k4OMv
XHVVzjcZ+5Mr3msloDGEnphKeH366aPE7nTc44ASFRQF17t+LSf5jYBZ/th/JgVU
lA6IOfT+FHmsoqShbuE3uIhDvVU3dLhQhHPzR7lvOxgHBRvBC99N2z8Rt+nobg9o
9geP7iwtRX4DufejIWo+6AMoWmPYtuqnXapUo4HjCHCJbHlWAJSg4H3pTMJlRse+
NOq5vWWxJznfYTe0c7eKi+4++x7xwyDMOyaPgu4XfQyrbrq8XHD5aCCWpDj5zWJT
HlPd+NUzi4MXOg/r5nU3MO19ZcJ3302iGwUfBUPe0Aa9ZizvSPMe8R0tLZ7f1cxg
N3P3IVVCB3e2M1uaVKQzRkp+OZhHgU+R0VQ9J2rNk0TjaWO5pVUvzXt59MDMER4Q
SAZFhFsTmuaiX2rSfwJHxUwp1zloHkhgUIKF1emGgyC9lK3lZtCa8vM99t2FnALn
0Lx+Jn4s4UTxnudIweODD3HSJy5uc8E6cVf0pk5U7o0RrAI9ALdUw6DRk7Be3ky+
4e9QVvSLkoehrxNiV2J7XEh08pPer4PRVikjfnxqfa9kJIE4aPaq3PD2r2zJ129K
N9U9lL6qZF+dMktKt2P30je+HBIY7/qrrV+1kvJRG4DrGrf7ieMmywuxND1clW/N
4GGgB0PgslbbHLu5/3wPuANVspbk/YT8iE65fLufvmPwhp94t20UarrAGNGAu7rX
cW5qE9VaL+8SnjJf9iYp/jvXR4GwLhzCAYsPJGYON1HWQfPkUI1ftf3KBi8aI6kb
emx2LA3GGbh4jEWRGBofs1K3CTRjH/fRgLzinbtD3ko0hJlx/djYjdfIoqDWqmY/
pSfGIiWMQhEAbIVN0wPzr1ltVNjXdWPIn/Xvpyw2OxCXtiZKUNe6XnwGcslSyuY4
huMvnG+UBcPy2LmTxW+r+EogVzMtRAlWRwXkH1aWiZVBzOHylTo9QTot7wYDKbDM
RyzSSMzZAX46tpB5kzARKyOdbMLm5/37OzkZhCL52kCvfo/Yty4ZPiYieovCndt1
8I9LuOB3sGu9Jda/bo0pypBf4BBwlpxVH8rRcRjdTD/gzT85gksDKKwTnc+ARgwa
kbqEZ/W38W1HR9Ru6qdu0e2KRTDiXAHGQl7SjI1siMwSVDyxNSACH58wyQG15Ma4
xH8C5UfU2W9zWrlOpb+zj65QDaqG7iHyjpaWLQW69Kef8hZyqOvZyMAgdW4tPmb1
Dy46E1M56iyoxc6utboNtfIprr+Pj+El5rMnUfguJo9yfRMOxEPczQMwxUBKknbA
pNSQeyZxi1tEENmNvoAGqmpktOOyK21sC2qKvdZfoxB0ZHRF/nEGc7wZw0K/4OAc
6UQIISpVABk5YuUd5mTUiOfZGNabRSOoygNoNnVHwvrNqxd/zSgaZVcPk+GuMk01
eSejbAhwczee8wSKIDUMIx9aHvDI3IqekFBL1bqHW4r6esoVTBghcdwxtMJVDDCj
qOt6/9gmGh05m/9Se2DBpYlBh6F5KfXemv0es9AhfYhl+x4iZBclPplYJn3fEjBH
ddwY/riF1tCswB9F3FjVN/qDfcf3EdsYEYXoV55nWGX6WAcE1XAsGE5Uyveh9Sh2
Qn4vKbKmVqbW6upIxc7zZvUQ8/81cobeN4NcgwBWKwwqgXN/iG8KMnMENN5Snqjz
XeI0KdmDEM8h4LKsdb1zJdKczlyMOXBE4cNERQkeuXv4cO/oOWM6fEEjdTDqxqQU
YQSJ0DHkpvBvCZ3SEYhfCHMDaqrbuRhP/raZM0kvNbzOOjqHQa8jc0QmKxogtHzF
rpuTmuK5rEnythbPCPjSoXRnEWUOJnqaa5IMrovht8ITkpS2pPrGkkI6rQxaxTYj
q8cPLGVeUDM40dBTJzoQ58iwfyoGc7AovNBX4haMHVk=
`pragma protect end_protected
