// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hh/RvbEWg4ztfp/mVs+pRLZmvJAGUqG2ZM6D51ZGNl4i5pbW2c/5CpE7Ckm6CqF7
DzJfiwpKPGmJa+9QVisCUIgPCNFMdl4P2+aVfiYlrbKCEH2dLoetHOfa9ri6Jios
x/79tnnuekcuPmLpr1541X6/SS0KFCc/zWKdArEJq/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26400)
76zHL3hgZA5jDb1m0Pa7qz8r57F5N4lKx4fF3ycl+3AABIOQ6b3+qVjzB1oTX6/y
ADMTj3DHBVSYeMYX/KjrCXjLVPjz2eRaAyYfO7NLQep9DcG+MVarfk3NNSoudD2a
pPHar+wYYQK19p/+dp0vpzqV+x8ONKbfMDry6XtMWcN76cPBrubV4p/GP9EIqyZO
gFwM9HWF+GRLH2f42OvTNBlsZhJUDWnL3n4nPFY1tZD7irPvOzpmQszUNvghtxLQ
znMuCABs7Z8pmVqfqaK0TWteObvk2XYzh0vBNrbEF42Cjaac9inBQXL9Qs114nQJ
E0DI8AjMXrr/x2/+OATlMJqwaZa/srwB+tdC1zlgBMJLNv1iqgKzjKFWBVeyq/Oa
dojv2Ir4A10RR3GqnM+8evwMK7bPWseiRN7gaRVQNcZb9+mduIVR0Irp6GXs3MTK
SjlxhkA3SzX6227qf6SE4jYcwIyHHq4CxbNWCqjEW58tSloSg2yyjgDuteLSlQby
7fSXjd/AxZFikBHZZ+MZMZx59zK9vRRQlrL+38hMVOYVcQaYJ3kWK2CKGwlYIWq0
1re3Q2C5/+ELi74rWn9kMJ1yz6Z1jEhaznaE1ik823YKxROt7f83Uiz5SU+r5gPl
XQGD9RnX5fPpt/vobN4Nq1CaL3rVs9h30yoHG5VdBAXvfx9TyKhZZohp8VpHCsH7
djWpGxbBzekdKDZMqLA6DRKY3KZ1jT0cfCcXOgd2Zvj5uScPdNcDHTpEKcyeMIUN
tkBL51FAKXL5Zce0b1HxMi13AMq7Onj1uKBbwDuGaWAlqXHJMR9Kc0e3K39D1TTG
axy2tkfTA6OTLvDjwghEULd2K85w3f1LNM0e4x6E3oQ8ik97/gcQV2KkNWDsiNei
VAi4RWEPJF5DV9cSqWuHKXbbXDP/dEX8GiG/+++R51OqDWmrNfY8FA4xRk1lmroU
pvuXPr1WlqNdaBIegCLNJ7E36dhhaf96NkJfD930dzEImDJR9TunSfINu2EFTPLZ
FO8vFT+XMZQuipg7Je4EW5LbDPDlHqZmXaE7cBO8PqHWPxWVPp5CwwkLxhP8qH58
D5iXXNCmY0bser8EpsCVvrSx5fYCk7zuQzSK/eisgTzFnWfVXuV7IRHxtOgZTCGF
T1zw+Zibvb5iAyOuSHRoS6Tnoh2XeVMad2vQQ4e2xMz5U14Lxm8VsdA20V8Kc7dC
+lqUVFhlggztnXF3a3UtFqbIB9TLYpUmuskeXbYDyMpRAbidF4w8m1VHGhJ4hRLr
Z8WRoJavJ22hG+GWNLTOuecdk1eEd3oCCEbFnSjsrBX5mLgZhxVGZrRMbOvHzkWg
5Jq4YBmuM2R2gl6JHvr6wowvg16l2lCuZTMJB4YQch3zGMqWiRhMUJkmcW/w6YaL
xuKz6MSwemr+kNLvPfyoFY+lH6wKQUyyQaQxEKyghuAGYs+IU/2qfGmC0QHx53fL
b/Xf7wu+p/yIZmF2Wc4oN228I4vthVjlMykYOWyiaUGWiG/KYcP12bH04e2nxSSy
SkZ9suAT74mVObl+wF7Dz2VoO/nIkIfuTMBlSOLAZ5I3BxZOyKyuAAHzzkGWozkT
L6iaqNRn0ORa+jqjfoU/LAaG+GI+PNL/BeYS9VVnR5ZVSHbYTg69+7qgnpxokvTH
10m8bNuXkwtcRowiP2jg7jN/2lGsyJJmW+iSGMJpG3Qe+zVmtnFYoAGpnQ0XOGlD
t41elpA2Zk4BSnFUv2fKi4raTFdn9HVWXGkkvm+dPzuQ4lkhv3wzpznD2AX8FZ5J
E+hSnxco7sU2n2+V79MDOUsDDqBDsuP29uSPT0kgbOeG1zNq+w2OWNtmga72k1Y1
9DOUyBp8HJda4NYlxdVtDCLwftcy0k2qe7L8j4kygk6mHVz401GxGMOFwH14Fvoz
ywW2C7QF5JPYmokkJY3+Rj6Lvbkiw2o3TT6ITodkecIUwWWIZWO1ThbQHqmz/G+U
0PXxNvbUfOe21ExG5BTQQixjhwVGPlbNMrBMpKYEvZTA7ZkfxwtS7xrgWsO8oWwx
dbCKH9jW0e5T5N2AdvF13GezDlSDJQmwr+k+FOnpywgKIaXyGTP5/F59GauQq5uc
Omvh6gwg5RvOTiRd1ChdeywkCunwAfCvrMHfO5v8z8ZKaotdY457SZvpaCQ3OJ5M
z466EZSa8nMgYyFCbdU3+NmTIi+ZyM4ufice7gnv84jHsKhwM77DtXWTdFDlvCXb
qrSCE/Lq0IBZ3TcvMAKi3wdpFP9A2Gv86LcOYS6gxq/4I5LgNfghXRat3ZcYUQFo
7NSby9GU0fZX1PY5zdprd17/TkjCPszl2Z0TSDPSDaG6q5vrxUaV50yDcWA0oDnO
NW1yUqzs3wMIw/phZUfB0ypwOCS6OqgsFIQpF8M4uZ4Mc/8an1JKp0qNpBtqHsEb
k1FCAA9cwuCeawQ+zOvtsN+z5JSouojQWFla0K8Vqd8TTECKONSAc/WW2QDc5H3C
sIFQKNUy4/PxWwh6h+06bjTbpeW4paYTFQvKL6TfiUsRJ01J+jCuPsovxN/50fYM
JczJbNNsPDTc8fW/pPWEA5VbVZ6Q8VL8jfgLJc9zgrh/WaY8LtcEgbQeHy3/OJLN
yINHcSH+I2HfiBlR5uss6IBIOawCfpM3jw1TJ8XlMiaC4erMYnps2OjFDpWXyASD
gM/8dnm5ldM7kknJDuXTlLcBnd2U/dcyiOZncICfE0Nlsm0MgadJRDx8OeXQxGzH
nIdxSKzg2xtlFenklJz+47vN+U7KGMrEfMgGOn0HjejecpPkR97TIYQNrEnt4vR3
sZBk2UoBnXIXUCxnHa/PM32Wc20Q425FMjLiCDDObf6/UWWTnRRTbFpYnpwiIV8X
Byp1OyWWnsgkKh86FA2O4HgR4glQIAwv1DDMhRTnIuHFVresKk6FR5A32sgw5CKP
8eCm6qYVQy1UVq5cmVFIJa5LxhrZznTZqQqFjm0eTaSHFrCblcCEOQ4BOVkUKw6u
j4eCOmZxOYH4JEZ/PILQP1E+bnSMwSty+CxrPzd37J3jRGNdSLhk+/ToIfq6QvP7
JonMsgosm+nxIfhTj3LQ+Q8dBl/GUik236RqrA/ezNyeBRcHfeleBzeRijSqFzK4
GcMmDv9DquC+i2Q6bhMgC2sAz5zV7l4QwMTEwTYLxzfTjGyZX3JejRs3e25omA/G
kKbDK7ihvqAJReQt552HNne9G+O/UjvSFE962HJWB9gdRNXBQZ1aY1ie2FE9ACdI
uwHZZ7ujaexm6//m8xAoigVvEEZS/O7mYkAYjikeaJyb0G1bp/7IJ7mM7TYYrlAy
fFsEKXvyavaAEz4U2fDtUIzIuNnCCzM+FxjByhUyY9TB0C9UM7up9GanCyBjcV1e
AktLWt13GrBQjVfnrg08/tr3yZE4fz8o+EQ1/eixZz9o6BJYa2Lr0JtPjahBo5Fz
SyzbR++cuf+A6wIXzrRq1K9WtZLWWmk+J1OIZPLZBgib0QnPzIwXgPYPJFwzbhFK
8wTVVA5CPfWlG2FDX/JZNYbQof0RmU9UxBgtN2Rdd3cftcHU2hMoXdPZapImx+Ns
6VvE4S6YDYyEnjumlRUtb+CxZwDYptSOMW3/kmN9+nIr8b2Zx1AoArHTPhJ04MMC
eKpjlPGUfpyhnSkAG2ZhswQA25nfePW5UFd/U82mzLMQA8qyfemUKzCyI+UZ5FZp
iDe9DqP4iO5d6Hue8a9X6JZ2bwjMgtvokMhm8O4oI8g3Mf/NnWun0ujOfx0pEWmI
DaVw5E8evRSmTgb4mBmcW1fUv1j2mHDPI+1HLTH7GWUCpHPAsymnk9iyu9QLgGxl
fEK0Ar9LvjL381ltJkcmqdFYyEq+0zIeENuneRoV13nc4xKCu6rn205GbFn9bkR5
NruLkq00/giNYkZ7sMU979F0zY08WHDG+UsupzTiiBT0UtSuFVE+1sVvgkKXNN8V
K/0R1m9GmJYj/g7ljkM0bx74+dEJu4R/8PKhacaDJxx1jiiDQxWGo1z202bC5LuJ
AjOzdiz5RjlN5cZ22FWQZj3JEpxzJzi0QjS8j5r5gTcp5UnLnlcq1bxGEASltq2Z
GBhw+c0S8BPOyw30vNxBHVlpz8ol9Ok/i0J8r5wpYYCNjSoKxHQpayhHaJla6lvi
yAy0IiQ3tCqQLqf45hWDl04LtgQ773cvZp96k1x8xRVuERkCyGqsHuvtuihwnbnd
k5qzq14mWj5IvBR4ByALybAMhUYeHqd1to7LrrqoMaIFsQaRPxqPILyF/IpbHbfN
JSwPB15fJJ6lEbvyUm5V7s8NzegJ0qZoz9yQEvGf4aRD2ZxPp8YhO1kxLdZ3QQZF
wOFOEyZ/XJQ4XiNsISVeYPVsOsZO0FNcaElu3Amr4WD5kYzNcHam/dYfM0OgikLE
AumrfFarilOtXX/HgZDHc8CaDNiPJtB9U7LbzYCFyybMOjl33q/jUOuFjvXTDDzZ
omVgNZ7YeNn7Csfi7QrsbPbHKpk9CgPTpajURHhNU/YX+2k3Nnjgwo7N5skMSQpw
YFgujryzDczRoJ1Mhtte8I3yWd52lKtCfIKi4YwTl33URzp3Pg+Lved6z5kP2f5h
DDvh7ZfD5RqQAh2rPxifPywqb4SQWfTiqwRTJXvqBvAalhdx1ot4+ZQhdhTDt0Rb
0FeRYi8yMjWrGT7PusnSpMQLnzLNy914jtGSMiwqTJfq+2KVijkPnaScRcPWSqeR
hs52WfFb96PhPXMEWoPnGMOqFjXvz8ftmCmsACcSTeZnWTlnbSVN2ZAjsivxy5QD
3B9BP3/gIsrJaniWU8lZ2DAX6uXznyeCt6h+FQC00lcmW50157T7o1C8hxKFRnAc
Kc5X3isVbUbKXdkhk76TxmJPgTA4ikjbqjak8WkQRO6qN9v82mdGnyw62ny7d5VA
PdrbshPvQmihdBYPReYC4HszlsL81UBtc1oheS+XVIlpfzO4WWpDxFYG3aVIZpsM
n/Jg2ll7yF8xz+RnhPuuMDf4IbLi9eDEqLXsMUvHitjZ3E1+BznBnAH0wcLulMyx
PPcevVFhHCFVRvzvjD/Bbjs17oByR5JsoNAYUhRFqjfy+2lSRI8Ig7amEMJrikeo
nNWDzl1ktYNEPDk/KAtdWtTUsgaYoEsYQO6xrf+lOvVFYqWuHoukLmmGkc+dVFUk
moPce4upI84K7VFKqYowzzFlODghScxdmrRNz8amB2+ZjrTS+7Au2+Ktd63BzERN
1L6BfUtMsOqU4NG+5UhxLevVo6L+DkIeJCpZHaIUJSHsKCFgX+CB+vKYFO90wMEv
Fq3EKwJ5Ym+U0zXq7jEZyenDApf4P+Ovd4ENpLjak7GZoBIUbol64jAf5z2f0tX1
t0HRNG9sHFtJ2dqAYbCkk9sQ6l+vi5ty+JG6JmmPf6hogVYjqT6BvNcD6rf58Agx
YUH14BQms8eMJ0dP9uOpqvoAkbAe9UWaiRjkT2oCNBnJbpR7C7JnEN4mrLLSaM23
FUxawlJR+6dRC0DZ/YcGuIXCNxDXhK1Si2V4NCDChpkohGVM85o26DJqb1L/6bTg
gh2ayXaKQ7+xR1I7Zf758/Yw1Zu9PR1VAYQZTaTsNvQMYUJZg/J0UP5SWp/cjINc
eGYsDdrruxRC5F9Urixa89Gteq5omAkfIITxtFoTsw0oc2mZiREUFrJCtzWfpZf3
gfSiIQAiLqs36UVIwh7m2RP0mQXG9JI1ez/YExWJQefF0fOMNtcFU41iUQHouzPF
XFsvbOwOaJOZpPiEW3ENI3Dc226mnD8RJAvWWYM3r0Cqq27sq9B8lmCEeCmrepUv
86r4DcyltjyN3nhDUJxYZ8WRW/NywicIDUjaKilQARkYLI8IxfXmfZ21eTNH4Oyb
EZVydqfpEtu4HzQpFPvsIUIn0BfV7citKMMZUxKZwrPm7eKvs6khCscv7uV9pC3P
C3x1YdMGdUbn9rioYl7OK8M02CK0teTNKKTr5VV/x6XMjWAVmjHDEC1CLWv/SZQ9
OJt9+Sl+WyfAmXwr9cKGUIxzZvLkSSxUtWDxl51wX0rN/S4P2c0K9aOEFVp7aSus
eAV8Jp97WrJGXrVHSvIlsXILt8JYI2kSJHG+WT28a+26I4rF4Lv0XtdfykJuEGjD
Ob4/j9MZr71X+6oU1MsLxeIMY6csDuBYT6gRA6p3W54E1VajPTIQ/UIJYn298axB
ZnNf7D3Kzt1NwieM9L/2Ee6kH7oPqczfh5UH5E3pwnh7mcv6+dNXV5kabFq7gAEv
gxNIXdmtDUaL3+QN+8HHNgZ5WXWWOjxwHnTbesWWkeKX7zSRij+T52cMxnYpmfiB
fo0t8AyYhAvkkvUdtT+szpM+5rXrGJ1lCOPGfdhJQ+z2pOzxT9rZfPj0Ki8VDOBB
Hh6zQqstPI98iqQAHksJwzoS7iy4TKzylQ22dVNGio0BuamDsN1RocQg5ZYI+fK1
GvreUYF5YXjs3ECDfcHiWMMRY9SLGh5MO6YvNxSFcAUO4iUPhFmR2AtX8jVvf9s0
0va4folGwLYCYBJ0FADesuefq/DvXkT7EUwDgyEdP6uvveKcEEJDpsXY7mLmp7Xh
OQEYr2W162/+4pOy62DCqFLGSMO8ugUzZjJh26mFMV6ObcfZdjyxibJY/0MuPFQZ
4rK6zH/sbNo23vQCbfZXxy4s0De1ZqwyiuTY0F2nJ5cNyYG1xWKI6ODu5leDo8NT
lyT+/98ZJl82EfxTbboSi4YJBDkA1hDZ/gMPuivZ8QwJkdfGiCi+U5FD1gjSe1Nb
VNG1Yn7Xw+UfJDj2czyFKzLETRDMzA0S2x8JunYlGY+p7C2J7d1LGIppw26LEZ4n
tsNw4B2hRUqPxPh04VY9U49/HPr1F0SPeo6TCbTvZ/BOS08dUgbSWDdc42/eDAq6
n4VgqJ7WoZr9JH5hHJYNLj13TtpBineaC4ysKB+tKyEyXXcZKV6kO0Ebi26DwEl5
1jmgd4cVIXFnYwgSNEG8jQ0rG577iTLVZj+bQvMutWp7mQrskwuD2noypjCMkdVq
CPu+sbAQ1G8cgPZ1t+5fOmDQWbD9QtvRH9tAS85+QMQBCDvPYt5xkU608AlX48XY
R0EZWnL4FZdt91PEdO3ZxmTAA/d+OeSpwt3Oy+XrUBUUq47He6q8wmXKK4MOJHcf
JGeRm2GduTFO9kDPAvAyuHbAM2MlvJsMEx1fzeFrC38M41iVQ6x6gTEzLfG0uKAC
RZCtUMkB1RLS8EsxRxSjDXPHb9NRj6kTYKTlFXyHNYb0MgiWV06bIaC0LpYEuFrt
TUYJynsG9XivlmAQwzxWLmVmPBeQxdLgjbD8p0StV4tOLd5CPstFJafR+kDm+4mc
q15TqSwG71GTaAZN8xberA3il2Ea6qonkfq51gA9YLZBuXxl0wnB5+b2VqK8Q7eF
KqH1KCwSeoWliVD1tIBkGj4biODpl2QZs9oRVEpERFqjP+NFf+zoAttlqn/HzJoT
z6WNcA2o4b3k5zuj9T1w705jnsuLEtg4mjMUcLz66hZ2ISP+a5nwg9rUn29zFXmp
j1qqlvUbnhqr3Mhp+Emalsl4en3ccFyPy1/KVNZ92t299bhSTZy56q9IUTXv1Su7
P/SVl58nLkD+ULrrzLQuebXFiAekj7c78a9vcLHsk5f+bXibFqV/8wKpcLmnTGVP
TJB4P+0xkUmY9MUzNZQai7QUq84llw1Q+2XICwyjFWG6+4aNFojlMSoc+ahSgBty
CNW9XOxJqOQuAOAFSXoUzVr24z5tnBQiZzu39OSyf3jAurDHhQ+mBhlRrP4X9rZK
ynotJNJ1XL0J94RxIXnJCGntIt99ecIYIGQ4Z3AfEvQ6nkVLWx/yYLC42h0IkuRl
7wfukQyp2NyParwkNCE0Hc0YkJaT6nCci+3UKzMGPgz/pZc6+meNN7ZhOr0vfADM
T4e06Ns1T/jSP+w6o2rLzozqFe3DymQgQf9qorsW02uJzIE/BXwe/9pr006K9bXJ
DeMXPbEE0UHcZIEm6NSr2pU6VZHwS07Av3fAKlQjfy3mqzdPDFaH08pha+fQh+cl
4QJlROyz/MmRIrQWu1sDFhmEwX7mWf1LR1E75fvK77mOvXyABHQC2M317n8Wnt6p
NtyjN9iNk4/9EeD8v1r3kC9VpmgvJAmZYwAerLYrAB2gFfma95PZeIU0aplQmjsr
yvGGnSPNgj3It9/vTLzqTTsodtFEv0QfTXSWcUK6AXOVVfyRSDcgLTd+90RHHI83
iZzg+BvES8UZ7Q1Et9Qk5S37UegTJguwAIvAMQEGmQnFDhidGh5YG/6AP0pzk4tD
MssBI+sZYTwVuTBQx56uVQPAMIxs7hRgL2Oa63c4ToPk//L6Yj2SKNECWm28uYTr
mGpHZ6T4Nhgbt6SmUsZdBL7E/bwFHUCM/JJldcVgHdzai3D6a5G7WaMRj51IBXmU
ryQLxUrmrv7heaekvTYH8bkGtGXNYjULxsUW94xWerlhsyMahGleg3azMh9AkRMs
oMl1yo8U7HPmTiFWsT4FRLI+Q2IRm87U/NHsL8j9uSNt6jy9SVIZinQ1Em2/pJ5t
8Ai88zphHBvKZM7slB6eyDSLKZczxnB/trXhcpti1JqEky9cD7kdSLu11k/y3O/s
Oiwv/YvXLf3XZpiVyvGqHTlzv2B32O84XjHwS180Q68OfiIG2kUTerF4NE5j7qp8
YB4xBgU+gIkNHcbHsE58lOD73VmmM76nlFakiZaejReA2j7uxwL/D2fW6PZxpPVX
iVGef5IcN7H0s0tnNv2JOnaSbM/0xORfWGmJCz7oVCoSFtlp/4H1SY14J9DmUcJt
XIAmGmhW0kYnNdIvWy499LXbZqt9vw5JYKVmr3HcrV/3euGMyBR72vFoqGtgaM/N
AILmuIk+sAaNhFK/+ntxdzmPjvGDov+pQlUGCv9l8Y+30JSGaVvKnxS1C2Wu5tST
5DZoogHjQmqbd2W/PPPsJdfWvF6G9XVGmoH7VZ4pk0kAw4mB9f1oKbt+yYB7hvKL
WU9WuHuld/jBAEJ+newa2QkKAlt8KAUa09ftB4wyoomLQwQ38Z5bK8Al8zUNvAqS
1yPzhjyNhp27jSHwYT2JIeetxIvAAoqTVph9utjywr0LaZYWiOJO71zK/pt+89j0
bBhY4fEwXNzp72oVMgylh/n3zT1DopQLaD9sM5qcRNvkK0/497uqL7ckLQRekOmv
KdqyV0KEO0fIVeb7QXrRMG7/UeY7nrug5A0wyY2CYbt9FETAaudnD7fz+lxKTrO4
GFsIUmOuB85R3VGYBSqyT6x7V/aJ3sjeL4DsaEe5cON2muHHVllqVSXSiSRVM9A6
X4yBTv+8Sf/To4ktC6nMsz5OWuQ0F631ZgJ1RDQCUHdKNe3TkKuV1KfKQXh7aTRS
7N1GC+e+MfW8WJKXWm5pH12eSCqBsKsrjuuGNFzlPwPMJvS4l/6K6emMuZdK3BaM
gvUrd7CcIRtY9cTQ3zkc45ROPOkLuGBy0BxEgYOH/DzgfEKWCPCbpA0qjN7x9Hxy
n67ukCzNwwTYb03qwhAirXdpV45puPXs4Xmd+zDTL3l4NtjpY42JZdbgHcj44Jzv
IanA9wxNyfTkEeiYM28XboIHP2CCELYvxJiz9zV2DKFuyGe+ugUkZWvOJ5MEpSMM
Bz74vV/CIdc/4AtMZITcRS667dqhz/5srAbkGP/B6mWhwgEGOjJLSSeAXI1+luvW
whzi7xPMeu8C0izHDJxvZjSzju776Gbbix+wiQB00xtvj01qv17FDNFeDhR18Fy5
zIEPUPd1m9UMMlUdRt9m5BLKkRuSLgD8Tds7z9uTzp3mvEIyozGrebGxX7oYubpN
vnykiQJkdyBSkadQoXbPwQuZJIvKrpxO7QAqTqKxNqi9a2yWDT9z5y26mvIdLEie
7xqrDLudGZwJn8GxWLC+lVoWVFUkaDiTnplJeGBKUag96TpvUp2mgLpNO0JUF8u0
TID5bfkZJSL2nW4xIWV9Vo84BhQAe84UzpET3jRo6NUg+X9C/Ij8XQYR1QF0Hm/l
eEc6K1ywO189N2RNAJ3CPfVLUX2dMdsZSB/v0n0LrK5NZpdNYoyGzVpPhRstYZxq
CO4YRECd/fsqqPhR+keQM+NqIypjuDumoQBi8tvGGQROhRFheyM1AXvAwtuEtoqK
UzdfX5yPSCdfPX9FHNOMjX3VlaqfOtUend6jX3QEWyuoUk2SlY9GAdk0yoDPWH+U
bJGkGCRa6NW4CbElwoPNz1/5yCVzGuzO+0o9dpnDpDkI4TDKGZGa80sLkoNGEf17
tMq9o+29iKyb4t6DIX3vGRQWQdKTg9084JrZNcHqmWY11wOGUYEIMzmffMsaOKUz
M7DtOYjq/NCDjN1aK8OPHrmYcxtSaT89zXzu0r6SbL0p7ooT1H8S533eDjUpQMyl
NZnEnwMCMtsQda6pun6yBQrXP81N03510soNhVYBgueioOHbHWD8twJ2wn6iANXb
/FvglySmDw74aGcCbF36g9Aj0GOm7Uxk3DYCC7rrATPRPLRjIT+oOke7y4PjOFbv
amSQiPiLFZoa/SoHUtQWEselGIfbpRW7qLJyRACaEbeyHg6jv0GTJTAYlYIDPbMh
5wxThH54b2Qwm9Wj+gVUnjE8b5pHJbFIX6CSl2ExTXADzltTJMQZFXZ2X9clF1Mu
LbYOvgc1cQy39ss/htifsLhtfWWdt0RAvIVukL4eg+GvYH9jjFzLTdIm9DrdoI1t
URhFh+wW7WYrgZk80hngSClQJMjz8AAFPHFT0SvQPTG4mghTGFBE2baShSyToKH+
/0BWi2habKw9dq9f1UpEH+1blZXjiJb8Hlb7P/I5FtwAOikphcbeZOo14FJU9Q/W
xTTVFFw68jD3EDfPE7DUXImnd9yEldAzsPWafWbhqIdD9I7ObGnhmy0g89Lh8SYt
OZ2LFRFx6uw9u7j4JmX7wG7igESxqb+o7rfFjJu+7rNScecUMlTE6vUlu8C9svVo
V5giPljiX3FSFe1nnFbi3UCkptdS3VLKPMZbaNUnmF7OY6DWpWllVtStZXlDNdN2
OV1bA0WdVhiNA/IAboYivrMaJw+Yaj5zi23sDfVuzKHwyWyd7xPuVsur78hV692w
QJsfZ4gsuvGRtnS/9HUlmN9QF2cUmIktMqUW0M0dWc4LqVYMpp8spO6BBDwhQQOu
g+EkRScCFV3PaYxmplCTbknAORvjtcQcL8t0HBDK+2PagdLArK1GpRhsP3a6RUSx
deRJJP2nBmNzmZxIpyno4y5266fHF2r+i9f0qdmgwm7nu5W1MYgG80Ra6HlQBlim
dI8//pkaMEWfAnjAEGx9xICQUYN5tJP+VJgEedikIDf/7QN6Rgbdts4Kfx2YSVix
MYjnzFtWa/FIrpK710VXg1CMfsmznWylGLQR708SxddlRH28sMFnkfol+TbfkE5e
1HdiM33ZZPmSI1ixT2iSx2R8E+reR9zyq1pemQ8J7comDmmBEYAJKh3TSEc94Zwo
VdvV17vYT1jmxMvTlPYwIqnXz6rgNy17nRMge8k57q+nptGQqk1utRlGn4ZMzuf1
omPryM/HTvvgofgz4pkFEkvZmTeVQvYCIh88KyQJoWpwgiX2FDNGZblnXApWyahn
1qQc5duG1m3zuG6QRABUygpNIYzRIqSm1+YAjuQ2hNq/aOCBA2lK+/okId0QonQE
MgLiwOOQiI+b61LyxHQy01nds0Nj9IoeDMeTvv13doYT0rIWwpADuPjiY/5HuG6c
qEc8pqj2bltRhc/e7Z/rFVuivXGFNMu9jrDmCnxLc6arW8sN1F+nRqx+R62L6DN4
vYpk8NGEcmvxUWpyjuV2jYemozccQkMM8EgRfW3vzPlxZr53dhheA/m/W0lJjcC7
E/ug6hHA8eJhkl+QfTkvsL5HwdHDselwt3qqG/y5VAGJef1YR/oKeDFYOTgadPZZ
mb6n8g2qYq7BfLIQ6lp/Sxkm2QOeUaQVrpq0GyawZaK3XFHXc2jeM45CBRK/evgz
HJRBW2PD1d1tg4ybTlZP3cu/KfRSf9wQ8MWHOr3/n7KHQGCLQBWwvN5j8aNX8+7w
nQcT/qZ2+UpMOiBJt2AgxVsUqqb/UT/lzKE7e4YQxwwj2bdfU/RGNPsjzMB9pHgx
laX86pebKpUiLEQKP7C3WVOkN4M/SwzxyhplUGWii4dJ4Lamn4jmDvlcWbPj6RhX
uQjEcbCqZAJMkLYhLj35e6v6CHXPesffNAZmh5+uPj0W+aF2L/5ZG6RnYVFyqE4T
LFj4AKdoHE8IHkgXHEBbiRWwNmo0ta5xGKGqVUrpFIfFYg3A6eGamEBLomQpzyNf
8/UlG39MxPTwojVWRd3gdFIuvN/QrezURARJ86bTlcFon4IZV+qWprjes7UHRCy0
aQ4HyiwaznYujBKR3EDtboZFbyySgOvieDzretBYFp8tlYw72fCJl86UzYK0A6Sh
ny2pb+UHzOzKS6d0CIlzewBge4D++U7HsdzZ8whq5tudrhvwOOTlZZqTBQtGeyaJ
+HKt8dSfsKGvExm5ItaGrVtlWWW+fBRmrdvv/R4/uq7Y+sy4zxPjRx3FIYqHuA8v
mt3SAR83fj5zdssMlD3mo5NixET1KLVntuBx2VFHww+nykEbeA3o/Pv0F17efUAB
5ppNkMziCPfjzAfzY7SijBDZwGRpS0OquJzqglvEqvjlzEkhxh4/QnAtwySH10vO
LFGwFUx8idb3DozkCX14Vvh9XH/tNJVYdMKAMqSnjqvHCaZO+AncHxnebtyQP2Qn
xD2PccEMbcd4Mlg0tPi2EOYi3C/JOihAD0ayzgdSkcxh1Ezxvwd4SsMPWszoTOtG
9dkVfOIJPHG2MPOi1lSJCSYtKGuuu6lIsVAby1aQG2oI2RLqYvE1z4YYYQ+Iie0c
HChMlgfEam6KPqXGtd9lrKbX7B+E9utZWX5Mr7WxOEQeR2CIaqxv7/+Xu04Dkqhf
J4m7+1fXULJRcaQlDpfg/DIZhyon6a0TDK9KTPI8It6N6LNHKWvYYMAlu1xZn1Wf
AjsFJvWni9gPwvfjeMLcMLMlS2C8N2oNUzfiGgPS5u2PRD53x222uFKZBArQzPud
tTeMuRT5eqi5UFShsY9FrZxtFFUB5tGWaA0AC2iNzKGZlv+nc3W9jId9yi4jU8hx
OZsdpNwbz066XCSHjQ6bPcKR9u6JMeMz3DQnTj9H9rijzPf8dY8LhEbPwTrY1DB7
ZzHX/LCkN+ca1eK++V9ue53eHwW0BMwcF3Agmw46Ohf+3VZXbpUK1dCNwOFstNRm
97J3cA/H3VhQPUaWx6ZL8W16dv26IcJJPU7/6zMv+DJOnI98TVRYSKP2UrdXmQ+1
jbGSsz/V59hvY+T2flHDN/l6BJ1Qlkqgy/L7aA77MIyuM6SKP5yn6qQ6HV5cFBQr
4/B+XQs5ntdsc+JAPC6u6Ely5tOidoKs38uewHzJT7Nmy2xCD+Lyd4CXx+RUXnXx
g9NBtqYx2tL/k7MDFEhmSUZAuEiFaw+FXizOmPttp7B2h3epWMbY0ZKOVj5sYvl4
hdneWydNW6LS3HnMfzr/FAVvMJpfhxh79Ry7XOtdxAvI4YkkpYvOpj4eDpQIR/fw
wINblsbY10ivCg8UEZcMF1n8ullloeWC8LJSzTsxlv/AQ27xp+1AO8/N9Nps3a4D
2WZ18I7lqJ6rYjgpz57oU8JexSrG3FqOaZcxyb4NSUzQV9/yfbFIM9Bmh/bWHtha
f0gBGdl/AKhrG7PU0kt69NjGS2qb/Kf4mCwPGd+nUEtYMB4gIc756g5j/Lpgz6e9
0qVI4kKLAAkaxjd9khqfimVxmAqsK8tMfqZk2/EkWsOqm5MXx42b6jX/+gs4jTRm
8m0Ago7A5zCTLX0b/26y3hQ2gqA25wmT84LNVL1vAGic2mvZ6M9zR3NtmeS1i55x
GB5GrmOWmbtUZbAFRh5/fnOOHRHr/lqLauroKENqOXY8SPOAqXUhy6aosq9RhJKy
NDEPOoT64LWhLGtt9uriMHKa2JbPZ9uIGp6RU4FUCDBkUQXC1d8itI7yr4DbBnc1
dxGy3JVpmh0u/6YDb56D1viWFr8tIkeWEswDHdr5Cl7EmJkJPBqqEHtm1J07pNLl
XmlZPnj1U8w8yo5oS1BbWQNLdlNdBVYMFm8EM87ptM9jodudMh3rYlsccALNykqP
llAj7e9wkoRC5o+cnMUTtvMpAXy3QYIcSXfrJyorn8zewN/vC9P31kwLC6QKF95j
ODyrokA6mr8lI1dMKfXeNp6mLwkmgwP6f/f3MNW+0Xeq6UgB3leArPMKMACIR6Wg
OAIUoDALUHlllHjOUas2s/aYN186+f0/fPNRQoq7qpk0WaHy2sr0eSwrqxLgzDjv
shYzM3Pe/sYSd14TCrgo1nlhgleff6y4Kb65pX6GcB2djqJyiJEZXtuV5JoKnPiK
+pwinD2ZUugUWddOc0O/79fJTVfNZRQHi13tgAJi0BH8KZn+SpmXZ3bE8xroJUCX
ePi1anKFqyb7tGsEKR/72gV8cm3UIAXxF5oUvjqEFQi5QCDULyFFnXgDIbIW7d+1
B2QvY2zd6xGyi1UawP4TKHQGH2JvmB6SiwLt9ocYjVpZbSkci8/cqfa45hqAiLOv
2HYfl7YlaLoMHQjo5jVQ87NP/D2rVsXpGXm3pHiCUh3Z8qRtl+kjjvxnNXlP9IkP
PgEv5735Q9kvPL1FZ/IBK0fDn9dWFchh2IB9o8SACq/td5sYQ6gBMoTsANsPnQwJ
Kv8WylU+pXyrmAEnya5HmHlleStbVPlX3/mWgra3vTWNxnaI6w+A2xgZenWfjUvK
wiFlfbWKLDzaEtVP6glSIwn892ACh/Bejl8MWtn1APOfA3Hv7saY3h2jyzwfy2h3
BH3tg84lfhfBZ0SLXrjs+2t2jbDfFokKhnIP9nWCwusRNJBMFEWWR2DRZNG+t3zV
CPdFx6calQNlSBiwpTs0EE0WcFjwnvFPJWdIaHgUMhi6gnIPz76XLc+OfsAkwHQ1
p3Dn3j2qxhJxe+B5M1oSKe2mfn6X3ZvMSMKrU828eT11zCw+F+JRwUEFP0T7VnSv
nIb8veeqedWlEW+ocS6Ummf0hhfunud9ZVNJ6lr6aJzH9qZ7Hl5BTEr2gvY1rzOj
z4bj+/HehWIi++6WI6HNJP9Q3C3HRh5VIFSoGlacixISTW0fWDRX/WSE7IoHpHCM
wGha09ShUAtSz4v5Z78gRZOmJCATYNOpYXOIe8m0E43xPAC+KUt+MDXABrmmPRDp
aBTPLSN2UVvCHI6bGQB5rHgD7oNWX7/CWhOuZj+CU8WyMw1XgReuhebIKCuTpOdu
pThOr8u6Gon0HFE5Y0HhPMjIkl8mxZV2xlESC90rpykJCBkjnrDzSR2rygvu2oGV
0gqlJ6Ju3ZhOlcD+khsgAEJuH+uO/oB468jwYjrkR1drWc89DLR0PT/ZGV9O+lQI
V/NtksIbcEI7n4LC482qCXsjErVfdGlNV1tUShJiN+ZgtXa+ABqZLltKH29vZU5h
F9Xk9WGeTH178tik+7KBWHKOWrNBNRRTjAAVAI+ajSqUi69JFOo+7Hp5UqMUWtrJ
dAkemxviH83dJ2oeDfXry0Jh51MkybjWg7UcFX3PbPToJ4t8xAHAdKjpYp7s4SL1
S/8QO2safak2bQXjl637qNLkpiYrkQbK3bicQOrrDFsnEERHibPS4kheu81KDh/L
2StXy2/YsWXZ4mzI4DUoTXAT3JfxeWorxZ270CrkH1mklDYffLupiYkiW6njhMCf
b8NiaP6LrLdJlOZaj6i8zExSVB8Ngv4A5bgDgY4/PqsXCia5W63IppjEAxpOh5Xg
UsNRkb0Wy+hUwFl+av0SgRqh/7t5RT9zuJaaJhHsDZi+6BNoLw3hMMwm1WjtpbXb
yXRp+WF+EA+9dZo7UAtP6Ss9BVeMIsjLU64/3wfz/wVtak2vKyqOCxuYeYgw3n9f
uw0tlBlQmfX/6vSWiG8L5SrR9R8+yzBv+7DH4S+YyVc8h5Ff/cY66Y0H7kBoows7
ZBLNQ10e82CmAlnlpSG2TCfA2klwqCD14h6Yz+Y6x5u6W0YvYA/LHImLeDuWAUN8
oZufc3ZUSKTfUKrzwJjRsis335LIGyfhZKDgKLa+wLLZej70+nseN/5+IiLuRfhp
z+7OOKOOFmxgGrc0k4+qCeAl6lCfLRvvBqTjKkXN5JtQZQhBlQUSCj5KMA2vsuIU
j4Ldit8s7XcOWL5xlL+KgBvk5DQ3OcGm92ppe6GKm7SBnBGfYHQEYWM/KiZScE6U
szMP+eShi4bIbfXLsRAUpsiUruGv5x8F0Q1b6mLc7CQi6yCYnNPpz8fvmlAeWZBJ
55RYo1fxxQ8iqHYSG+LWY/nVb5Lmf/zMMHlfr7Hg6wSBf4oBQaJIdVci5a41YPSA
c3AXkFHw54YkNfAieusW1ldrTN1St/cLsKkEiHSTBthmQGadNVVA6HO9nmbehSpA
8PGn5+EVqd5/H8rjZtQUBRxcLMJcNciS+lAjgDnwYpAOM4K52oYPGDa0Ip79Jdfv
QVu5Cn2u2Erc2Z7DB8y/r5cSgRbCR6L81+BPC2CkbxV+2g1L8g5PnLmm9v46mRIJ
fJDQ12tO+xdMlhy4C+c1gxQd8bCj3CmnWecUDnuFG7ASImyx82JlkaZwwqy9o9+a
vFYQAgVOmli2L8TCsOLokKHNwvL7aNAw5Tkrs6dFoyjFMoUyHdnUqI98+43+VqYV
7rArHY90kqSu8q+rxSYgqwX18eqmB+rGPCHx1udzeB4D4DJLe7ExIT1O3Eit4ppX
cFJVHATTPFzjbivpS38GG+g4xiuwy+MESRGn0JtjQ8M/5fhaKXPZw3c+WM87W73M
805HCfwQqLPrp5ZruN2OQHIz1aviUL+IXJQYGXP4Prx6hAdqpIAEuYPF3xy9veCH
YmveQCNj4ipadw2qf5bH293SQXw3AkW4VeK7xvZ5SndoYprFSAb4r2LgqbzfFYPC
aHGbi6UeimVHalX6qbj5LTPDTFREb8ZXlZi//SOFpFkll8HrwEf/a6osn3VnRWQx
FM9oS0+tG6NcBymYzhFBwkZwrQgtX11n3UlaSAXC27+ZqTW1Q5IabrIVC9JMczrv
VVYE0l011sE0vvrWntAb/s2jqfXi2Ku5JfQwOTd/QqVOGBadN5wJceZA2OeEfOI5
hj+kJfHNo6ZeA7AZb4QqxLvDToY+4SdzB7EhpMnQ+hEAziU295LSH/Wf6+2AIDmf
G/I4eqQZ2oLsCZWCL3xcFAbDxcmFXBAGYhTsTw3zgkPlBlnTFTIAtr+Du67kBVkC
RTg4YzrGD3wnLY8a3Y4pfi043dMDqtuSUAJoR+atNbMUP6om7JAT6SYpNVVrJV6H
c+oCqfum30IJP9isE8tqi/DkmR5v9l1oOHzr1ZF64vYVPKTf5CxAPps89g0mQlZ5
q5upuSSS+NAaoz42m9hIwKzbOpUN2KoW8W0YDlwzTLoE0g6RQPFqswcrVKG0TyBg
zM1/xxVTjZVW2DvuM2WK2l6/ESVkJULFFbofLp2v7PgxV0XgjZP3KvxHW84XtRjb
J4m1WqxzjQmJFyP5JRfaSqm64wgwaln5QfXB7AV1zpK1eifxu3DnJZYH0UFeYz+Z
GgsrFu4SPs1w79PXtCAGgZbZIakgZsH/HsIuezuak764ZE8M+Td2YN8tkSYWK/6R
AyncSA70eniliqVKa5tCDficabvU+35mxUJav8wrAO2+S3M4pgsWyClKNFllLVW8
XDCyTWosc1uJSxuQbtpDw/ooTJCt37yQSLPFIG7YW57i2kAh4GaoxFsKa6SgNrU4
3NQA/eArSde8u7toYmz4FlLfqiOFFQ7CP5WmbS6bt3Ldh3kDiu6QeM1G25w2GPYz
yC5Or1Gcu3lvBSBqIz5v08OQBUDyu/okgTH3CnnAOZ8ytmStZsAgpnsJBzPViKYt
inMySXw8FADTFl/Ah273/QYwa6uGgEBGSCblEIcvKinOdznA62aA5pmK9Xf2tsui
g6zE6Ed0y4XJ1+8DQzJiD3MOG0Nusph/RKFTIpoG1uHgyvnkLzwOtVkrd6UPgaAu
M9M2DaZ8zjDmXb2X1zoJmH4sU8G4axaQ45n3u/ou9IkfWkd70rnuwOs/YsEJm+Wz
lJhjEt8FJfjQyRkmoziaPw3xduMTpFauARdwchf8ja0qs7fqWJH/CQOffMsx2wbr
4mRh5LmGednbGzU6+Vv/HGRayNvYShHsCyGi9pO6wGoe8qlpN3OjEHZDGfNzZj8E
LZpBfWT3ZS7T8V19ebFnt5DifHQaes1B+e+xKcRj6PLHe+/fK1wdNnAvGZACYgQE
/8Jc+KnWdawfZV99F6EPeyjjdsxaJ8qfr/bmWXtOUGJjAz3hRnVisOXQm2Fp9f5R
8e4HBxuwP6AQlQzCdAnQzv4UBzV/5XRVF9a7DS372qjI7kPEwUUfSN5swATP00SP
jM6blkmN51BIS1j83wixPfEoJBzJElpZ0PLkh+Mf+wORbChvkaZI02hNR/QNZKr6
3QQUEgkSEdzz17yIWPTd085jX+i8CbtMaR65U+UNuj8cr5nxaU0CYn/q5V7ccoq9
vng1fDgvdkjqmJtgMBY6CGNU+lktaKfua7gNN5jPXFzW/Q5dwbVFYCYRMDPCpEfl
pU3iYjCwYGidX50ZXO9t/M30NFdPhT61iRRvE6VPM96Swh/+4+uX+p4TCf0iuND+
igTSxOKbTZgDD1tCck9YmiaGD3uOE9UUG+/jowIQ9AgW+vqaqwvgHWByodnj1UKH
zLcBI3q317qDRj8EjEioM6abC+sqFWIcfmEfAvQ//MkwPbQaSs3FWyvJ5zVJHoGT
aytFlk/XZfkqQ/wc1pYluQD7jxzqh8b3wsqzBsZ0sXALheITYeGcRDApNRJXSgO/
6qdm+Phejwb8C6GW5sXk5NpXVB0zo7YFd5TqW/jvsBJXnkGPzlOFJePhTO+VlJ+Y
P79ypfU5uSEdd4upwpQCRg1q3/MeWfZ30t3Fv9bPqDHdUPmVTgl+Ag1goSHb1kan
tAYN1gjskct/jhDylNNkLxAw+J4O/7VO+MaTAMMZsBCTMqllo8mbWQrbww3Mnsyb
h6r6cTOxRkQ/XQKt0+7VQzY1qmDFL6jo5V31L+pJj/dLU7q+QIGM1xOIKw3aIlph
rRC8j7BO6R4PJ1NaVKPHd2ZVDJl4S/7ARPOg5oC5xp8hp9WMrjANWlPEVMhQVcra
8ZT6JUNSLgXH0oL8Sm8iskjVtQf50bZEscpSixNHaV2uGyFD8yNJAa2yRhvu/KEk
wpJ16RTr1t6SX3P+uYQDeUVUWL1SG4+KIY1Oyg7VLDReFH1LhKYzCIwtQ9MnLu3m
RHixZJ8j4vzj83+XEMperwECtngN/dhW7pKvuvX36PLuuANTcb3GTEcvHK/+Mifn
gLJ32KISVkuIefDGLJDnxAsmvwyl9foTvhfQolDfwhST7J27MNxYX5CjO0QcrTAp
8WoyWn7ze+KqiqePdeOKe2/xrGSccRLWbQKekdiGxbD70+IRS3sF8aXe5TCqKAng
6boUFq5vSe+UWoddAimsyR4by/hp753O/G0JI+uz72kDO4DHltiA06ypRvXxifW+
SkbMKkjI777rNE6f5NxI4EaaqDkCEKKymDjx5T4YHCmXzAlUthm2UbaNoOVwbdOK
njO6zYKLqTyZ0svCtrwVRplBovadrdWNYlF6eM6zrCQuL4gk/nYHmVVYmy45AlJl
MPBWt3COsQQbGjdFCDz7T1WnrEUejVVmKM7hUwJE+vYnKT279I4Y923jGcM6VqDm
A401Skz0oNTJwEDM6WMfq1SfGGTVRVp+aZntSWvkUdrpnp4IOhYmt5Id/M0fEK95
tt2a75H5rEtxs9KBcmRsIOZAGgSP9gFjzrX97g11KPxyqR4J833hJGFjZ05kDsxA
R4N3m2T/V5qYUMdR0gfWI4PNEde1f46+S7YFVxN7Y4oZTznzKIYi2mBzUDXwDnRh
Ag3k+w2PjRfe+kR2YG2/BHDFp/L0PKUgjOqoEG5T0ecw4FfTLmcOWJCOqihUxF4p
1B7kNbU+QLw23eYk97hir5FxMKu+2q0mG4RUoqqLJdJhN3ypd+tDlvXLM/PcA8Vb
EFHTJ5d1eVqCQ48Rk12CDHNibtQOVu3C38HSZO+Xhti6R+rLXlhv0FfgtZuxwc7A
ImpgDSvH7jPM0okqfco+3OJaBdgslbJnoI+hVeTIOvH163TncykvEVVEvIHOZDbZ
4HtBlO5wwqLR/oABvoglhpDwWw+SUuQKsXwRJwHcnjixQRTIPx6eGIq26CamSVm/
suxpF+k7A6xsXYsqQvpAGx7jjGmWvehJVdhGpktJmysCcOxHb++w3XaSQZ9Hyf/U
q2LE61Tc9XnXaTnnAO5mKtpLGKIxEb+VxNAEpRsIiGrPiDHnwPL1H8lrTQ0B293y
vDsMMf4TyoR7DNC4dRL4/cc0DXahHG8IWnV6ObU3btsl3ExQcieZGHRx5ylGjN+F
8BpQ5uu67JFcqJZRKrPGjUfLcVGq3GjdWhmboP4DSC5US2PpX93KjhyK/GH8Scka
SXZNrjCNQQVHIFKKkUnLKmvQe/PrivyIc64L71jOcL8rZ6XpF0RvEqG4RkWTlqqm
7zfqNVm3KdTKRxX7o1tMwO2TTcdXGLTQr3XfLEdMK9/kS793ERtwv07T/Q6vurhu
PIs66WS8onugLCKrl6C6V9AR2pWYnNwxoQx+21mdh2ufkT4KRuaPEw3POpVEKlew
EHJNQSuPtQwQ2310xd5nfJsZEMI4dOs0sk2KyEJy6yIiOuJBUjYJcD+Qh5fKYx8p
DiwcXjksQwneeuhjyGAY9Of0qWaQJXn98dzjKMpq/68uq4C1u69eoqcW8EmWhLsY
S5+POSDHzYK2xsmcR4wAtE0Hz/160rgI1Hf1TOOKhdYLH+aYd1FYqTbIDd8hllPC
sJU9SW+sU0Cll6RFl6Y1PLYhf1onLcYnYZsdzaP/E+7eKpZyNAXAwMRUUC6Y96Zo
crkAqRftZijMQYx4JHrRWMQe/2Uoj9lLBVQjrnNxjNbXnKlfiC4P6I+tvOIwL8N2
UJNnXQozHvlQ1wPbi6x6Cy5vo+w/fJnPl/pX8Sim/nAqU59eoI0VxmFe4mdBcI0J
Rt0hfQAAXSps9d22NabDNuyYgETI7w4glGXlvJcALfxvxpDbmYq+suq8qtNLEvYx
QTa0UAQ5jJi5KqvVtUWcq/SsI+E82k8C/XddzG3qcb+zH5xdipifsDC43RsdU8OO
vSwhD2cPwel5ynmgBsZwDzkjevBRSevbri9KAIWiaderuZW8z92Q4Wf99C+SUCeu
52pNP8TWfSBkGrxW6S4SfLijbKiZ79xxII/Hhdf8cFISQF+utRUidE3ccxPbeLvD
ZWzSxOULrsJ/gPqHpPJkHrtwf8KT3i7i5eZIfceY9c8G/gaMxy3R1CJiIib+a0pg
fgT+xi6mN4touxsUUBAbREm4zNEwfor2hkuv8ORX7Efb0AQOIE6afMg0a0yzkhW8
F/cbyLRSqo2J2U9ZwUWf1rrK2qn0FqCLIh4EHFBlbzeRB7HkmzKiSf1+xGT7oZ4K
OKJ3bUBekGYYvpSwBAJlU/z/oKVWt/yIlIdU9bS7Zzo5M+zuo5xLFtN+CL3yK9jE
TdogxdjX1Wm9Tw7mXjmqGyyN08IFutTGRHmIs8HvSj9bVPIFxfUticoS4E1sghi4
IT0tnqZgsbI1G1otehX64c20ZeOQwto01lBXEVMqef1RAWlFCCleuKoiHpkhBGYW
jeh2hzfGhCyVw6kcZx/ngSBgw4Hg3h18wbESSlHxfgCloCTrr3cuGIHtIRNy9miq
mio2pa03zpaGR/tYE5/iSEavKqGtUip8MuGZ+fdWhgexdkeFZ9ef7hD+D/x/P3Ng
czPUUnRJAYO4FbcStDGQMp1TPMbI20YeroB2z0JPCszfl5cwdc3AZRzEaEdcgK6Y
F4wtrPbqfHehfWtna0j6Rp8TaB5bkSVFggVr1d3vMkrn6y413MHTYchnBoKAlEkj
ZuL1KwZG32ahYn+4NB1l2J52jFGaGPeK8j4b9nn9QOvwmH9A60mUadyRUAJuP3Do
7qNvQvaeON6UWVQ6RYmEG7hgmkWJFVPeG/FUxuLbq2OkR0BvhNOZmSNFy4yPH+nQ
rnunklze92nLP1S1rCi8rwSZbk4FlBlbbXQqoOmJvGZMFDF7oLAclmMIKys1uS3m
WtQlfqCkFbaf+N4ELhoffym7FVUSZ/HBABoXLxoKQA/PDQ5tvjQ6O2hij8vHOVTF
wHd9+K0gEmFRcnC7TQsMzq2bkZV9tv4mKCbnZYXmpqea1dC8y+2u19sJZwv6i+MY
VsMbnUZrn7XYhZ77vGZZIrz8crX9e8wZlJvc6kPGBr0mWYDklunGUMDiY4h7gfQX
ZmxhoBqwzaC/HpyTp22F+ufm1ukhXoOsEbHrkGI2zyh+aZIA9oBN/t7ROJPOb5hR
SbWJhR3Qf+2a7T+ZBHa3iJpXfQbpNILKdejikiIuXK7VgQqRN8kVKMQJfmRX5dND
uJG4aimGDaIeUeOFHwmVpY87uFIldQ7npKdnQ9irL5be7Jh0BUiYbh1FdoX5Gyrt
kAZI19ELDb7BO0qeC5wTypisPOeXQgUXmf6VLZiiqKfH0UXNBDtnCuJCy2PoFK+E
dWctD8OtqLX1nOUG4/FA/cnYeoLEbNEQJ5iRJjL38FH5KK5DhtQwYjEyvFwBlIxY
y05f1RSoTrlgG1GkaqQ6Czxei6ICz3S3BnqqfpVt12NJ/5cnCcuKmyjjX4Q3sgr1
Ks9s0MGlEVK7xM9HLH6jNh+7ycwin69OVe1vOzpRBISjCp/jZFQG8SWTT+FvqYhS
6B7WXvKii3XslYUvkintjRiReh7aUJmm/MpK8jaVr9uBJBppcUa962BH8d5YVI+y
o24SjrXI60F5rl/izdm5XVwlSt6sQ1FpRCrLvVYm4gWgRze9z8uIHJS2t775m5Ea
Yeb3nVolHEdT0HDZvlIsr6/Zl8CX/SPmoG5XbYj6wgmchGErxudaQgbHTMzpUdde
Wfc2lG1nFJ5n8e3JQ19WO4scLkanX8OuKnJUaSVJX2cbtyhi2NxmL4yLoCfbR21H
0SZ1Eyu2BsoZGmg5R+FYwqNEOnBSe9XbIMHNDW+nqRnv0T9fqQXUXr3/hK+BlXU3
WyCiXby4Y4OaeFs1qYpH/HCsHR39uggsH4KpPvRGj5TBTf3JD05DtBi4AUss86W8
/WxnX9BUEZzPCW/KhNB4s2/Ltkbl9bNWZFL5v8FC3xL4hqKMeWNUQlBWzFZZrIaZ
b9M7J6F2DsGl0wLhvHt1x3jPeUNT8JeK/f7CcXPkw/GBs5JLUHFq827jrYskGNBf
SCKIVJAJEM7WRA41wqU5Zp3mg/ucnZlB9w31OPLkJS02yOFXz5kVK3swaK0KMbGn
ikDiHjWbrOtwX2ZdBxzLpVBj1n9gYAxGTWQCNY0f88/qrb8rgRE0qCjaU77AqxSV
MTC/nHN+lNcVSzC+9u+4IZhqiVBDhHdJkr+I0GK5D8qKHWvbDKg2u3wNQnSucuvd
qKbcqGNwEkh27mMJEwIae1EGPWKYpgggRVmC8zGtX3MQhM9rQ1ih1m15rrAXVOaS
rTS27tGM6ucRi13SKtMBaNSSi6f/TPzMQXT5C6MVqZu5QxZkxHUiNRZE8dOgLAR7
gcbVJkxO5RHbrPiRmuKvqubwS9MAIZFWXFol1GbuS+/vhTC23CfOHOm89g+Dq+AX
mP6B+7yxpS9r8d/pegb5wZdmo/fli6TX11vXIgEcb/vldACJHQ3anxGj+5KitH+S
x4s/JsNgx9KADvCpJbqIneoisduZMbRYs17taUt6aaC1WgmT2g7s8rV0dogvd6k1
HgQouWmVrq9GtohevTxOedGuBhjUxobaHVPYH+UB9YDdGxyqncBlSIYHpOs2i6Df
567AgbIarqXetKW2JfzkK3jTPjKxaCtQHIsWJLf0PLmYD7566MKoZSl53kuxREIi
10mtu8VdluBkJ262x/Z2uWrfjt63mBp5v4DVy/y1KqpITX37M0SFbSQiQW+Rd0y5
z7wS75NmYGRmdiPd2DQGoo0LrmJOdF1y87iLXNn8znjNxadLUPPVDs6q4m3Lf2F/
hm/lUsWIU9jx6oY1d0MFK4h9ISZJUujyQ8sV6PQZmNcj+ej9BgfrSmGzWjamFHUu
s+WZLVm2w/WlldXbmWEe23027dYxR8Ho6SvNuMmZGmSO0gXtZ0MK7EUd9pQGq+yO
rGYBSPLcDqaCGL20+2xAESqwehRR8zqOT7PaIQnpnHQ0VAp0XDy8KecO7p04kHJH
xv+c4GAhGuaSgcdwGArGhxFzSj1OQMj2FQdR/FHbPb3SB+LbAzNtWk41N23aXkKB
GuDevHj0cL9Zb0U0rZGm5ylsm9jtdRvhWAffOoNjrepl/hJ8XFZDi/+Um3+MCRGT
9iJsxeMr0ynZOECBRafIxzgv2JGMGW+oJUmm0Js5COEo78mrd1m0OBQ62XXb3AH2
dRRm8Ouih0Xewz2RayJT3+M0Zae4t5ZCJhzlqBIWAZzmmD8EHx0g+hm7lmL9lCuD
Zlf+DVRK99xFNNexRL8R9fOMHrFWtMDt2FLAAlgXma8AnJtOqR8s11BM63mVFEZP
Zj92Psn4x5sFCVkQC75P4L6pKK0jOcrEQ8g/4+j3fWUjR9HM1BSiXbaOWryvn6K/
LYJUVUG23G7H1egO1xdokpeivbpFYdDfU0E6zkii4peif7RqcSvkyiUOO3/sYor9
FcS9Hfsmrx8QIYxkyNcPcMCjM/0vj6p6oJtqafrSsoJZp9RWSVMJ6X6vtjldupch
BP3NCN8FhZlFWYTdFB3UUTU8SABlBkKATCisC0/A5t0T3BESHkHZ1tKnDVwo/qBR
ehYz+DBKtgiXRH24VCP6hPr07oIoPCGWKowNiKz10uc9tA2nJM66yjYSa6XQUtIQ
NASY/JnUnuU+AJ3q8moB4XHGWhP3vwLVYqCtuT+AuWM3p26Tpfr8Xl33QQAMjJKv
32y1Yuse5iKJSZn85cFAz1ub6GVhZGBce9Wzws5acHOZ5sOpVEbCwXpjrlaEEVB4
L1P+NU3WvFt0XrO/lqNRfVQ37vJu2WjghjKRbhqeTz2L2Hr5F5p8KKNVnhokGPGM
w/4hG/On9mrcLCr3aHLX7BgFJn5hsn5T69uVXzmsj74QZ7RuvXiS8NsNQfsmiOrZ
SSiTJyw5lK3tHboQuYDt6FLsn0Q1OMmwshkHT4K/k18zRnegZOYjkRwte0E81fDB
4rdUv+A6iF7eeabAFvLMEQSjZR/0Ufu8c/QAQYrQxE/IDPX/1ie8bvw7zHW9SWrs
bLQMLdE1h0/gKQvvorEjLAlGaUyKd7YOmHX/uCmGdYZJZvWxL5ayZ0o3TCvnnYrq
nt9DquRtSDSPHwOEE15Py1yWU4qw6gh4KUfj+zcD8VRX6Aw7mJLmHhv34RImurFb
FpYuM/JC7bl+nHwjkjitsx//WTZM/8kTI0IvnRjLdypxUi0G/a0k20E1+VhtWQ3U
xtlHQ42pdH7OYeeq6jwyhJKlLaruWvqSzAUSLcObZhIfstAdCRAgFEqTbANa5qD9
hOv5U987K8AX38AvovLA5yyTxanepqsfNcAAxTsMimCPNBW277uF9V1dDJ49FLwC
LXKySDcW7Z3zmQtAcSkhdvAg7AGjO4If/xbEvcBTxBuvmqFYxmmKOaf9ur1PUcqQ
3BCu61u2hCv7Mz7NVZzfQqs3RrlA2VgH+TSJ0fsmhlr/vvy6giMF/rV61x5NW88W
j4GDRUZDQTUFrKdqWwzQsVvt9EjRV0opfUIVhSiBkdilioa7SOIxRa2noIxUz0Vv
jFDekFyNzZHoh0avgOWw+IuNcnx1MyV+nYD/8EF9ZsC5mlRRAYAbmpqcdUAfhVCD
LBWgpNYnhlrCzzByZfHFZr/Q+vzGjWCWIgdkL7WJT6njp6XtKdj0u6CNThE7IjQt
NkTd0nsj16J4+dSNRiDkOURp2u3aH6+b/fUVd0bsP2xNRuZ8pHuAbczwKTN6JTek
IBmR52oaJv0OefxdvReynrkX+NrtRyTcKVn8NZmjluankrF1UKOpdgjk+bF/jhDp
vi49g90yqO6a24GLLyzjKSrsgbveeMQS1bncWR0BP3CF9Z1+vKIOYIw/N2ZONfzG
PuoxBBzsVq6s0iWK268Ig86gnDCnGySsu2LuQJ6UgKjQwWMLlzcxLmvNCZhGh5/k
8+8rXC/3SJFvPyPgGqlnoxGxasfpbQwMHASA/OysJkp10ImbhpM7ZzqHPE342pio
KmMCrx2IK2WPC97Al4Y2ZpwMhkoIQ8kmwnomCeBme1voTeQf48Wh4Z3RwzrVeJuj
iu07KlcDvuvPL+/X4iGnVBj3/g19rulekeaoj2ktLpNuVj7IhENQilT96aDn7FIx
nNO9STcKXNUz6kH+m2+fLVxLjwG8/1cc7BWIwETnvwW9t4DN+jERHN6dsWlrf8u/
nva0Xdb3esQsUg4kLddeh6NdkFvPYegeWffYv4wAJbbr6wbuhGNW98Nxm/BmxSFH
Ff/2eVRBDtydgfni5Xb+Sbdr0mkeP2S+PpDCHXUityY2TRJk4d+eXvIaM30BdaED
9j4Dw8iTbs2xIJXOVkJWYZ/GFKp/XfIf3mCG7AkeqytmT3cKFc8SRTBJknaGDYmu
iK7Y6sa1LwNVOOTrk9OQP/F909nCm+BFv3BrSgZRWU2H93QKq/rjR2cXx8oMI6Rk
+GJvxI1QYNLqpflaaigSMqR4WlkQ5dQMno8jI+sqavvjaUdnLBQygHo8hNJsNfUL
eKEsbhO/830g9roKIQnJT8RwNj/5op+la503wG/WUjd2N1CU70ted4Nt3aiGhAIj
v+pgN0rtVQJV3JBvcQgaw+EVZgJb8yZyw0CBbnjWbeoi/3X1Fxfzg0e/XkZRRkbK
biQsXYGVRLPFDklaDawVfLNYZQ3dQXmMsQh6wd2H/F47Vne5tFB6gMWuPHyggzXW
fjY4GVwvQyWwcCDKTxMOtCNt0/HqHPTIZE+yvwRVjcplyw6Ud21ruH4uLPS4EdtB
sb60q570pG/rM8k4xujCYpwsAV+W6LcNe14Hc4/2SbDbyJZFgCsl5cqARt5hbiHE
h+9ouyj+VoGYryuGmMmMnxi/JrRNVfJOcuBJH6V5MryeRKJn8pLRYdYxUNZ6QTl5
FJvFnkfS2+xCxkByQFikenYmSIyEgYEqVjHdE4pINITFSgD5afPV9rceTyhPNwqT
Tv2yHZPPg8wpjTgHYIlvMSVvhGWOCaBhdF91bnhrzYj7sAK1Cm1o0IEaCAhfogIA
3CETKmp99UEC2+2QcfpM+2+hfCESD4RPH8mkv6Gfy/6y20VABdU08pTKJbWbG0ZL
WL0EedNjp8izPotnn86HBsPMMJAbn/XAsNYEYEeQSyZfAyP4WSpRlozCvdOYDkXO
xijTP8sSlG7jn3BSkhFRgqPzxllNofRv5GZbfBmS+w1HZ8QVbZ/mMKRPVD7n7nRR
0LpENaQpNgcz6OEKMt0+/RVXeMPoeI7ZAJIKGgxaa2SJ54HHChFWzP9v9gJS/y+Y
YEgNEw8QaqRTZbI+Inb4sziydpVTRZq4snsmgbj20W6Zb497fFx4WiHj97OzHX7C
S1t2fjcJ6joxedq0PGLLGH+NNppYqnM9d+/oosT9KglXBcU1hZi9b2NlpYk8NcyN
lyB3+5VpHHa4fAx7l6xhhBZ/F6/zD+9tlbMVw4tsAOmtd5k1Jz1fmx7BrB9YTGjD
eMTQIjeQL3Bp/iavfKNb4CJ0hkJTdpfzthVW1E5CzVHT1qirywsxIiA7taql2G0c
4BaE/vTQXpOdxQagjK7+hY4mPEKH6bpDcow5hFNjM7Dt7thdGOHg2AfxMs1NiwqM
r/Eaht2NH3gPjO8Nr+syeC4LCrwYvEBM1WpgxRRtpxX9AqnvZKzS0yiHzO2s4Gg6
WyVkmLwC3n3K2+0J6f3EOUeZ+dV9ZH2kA2xPj9E/tKcalE1oQBZ2ZEw3bfuk3nhX
napB5zvCQI1o8/HaNB0RE47tZByioptfgLZHfHi0/4Jb4nOUMvfhb2lIc+DiS0aY
yUKpw+olY/3GKuYe8qafFWbBNLLP9vzcDVoq5s7Wd4IyGWRF2ND5fYkWNECrwjKC
2WTHYmBoR+GlH75ceDPA1+tXxva7zNC89O/LYYByKn8btLgKzcD6QwOsJe4w0xn2
FVp8PGTEUvxnFj1Bd/XaeR84GyYlnQBN3S5xBvx8HCokx1EZhrauwVQ+vS6bMyb8
Y3Oytgd7OTTu/jWw+hpYRmOIJm4y409+Q/sCosdqVLQQUTRt5ub/7vwz9vSQDSbZ
RQ0DllMZtarVdEu+wv+0RtzQsahZQiljBakwJmvH9ZKMDaSf59Ie7NEETdqZGdEI
z8DjG9JKQDmqGY7hf9uWKjEGvE+FA0TUOEzghjVsLwxr8ZFDtW5OQS0riYwECIo7
T2UeJylvogXEW3tmMzSOM7dCdyeQ9C+5P1DBLsKHA1cf7Z+3vETop3Bc42lBcaq2
X6KbG0cj8Z1we3UeBhpntjC2T/RUT20OUm3Ojfaz2sp1IkvSs8uTygOwDeIAOnm3
iqVlaE2buYqyWG9RSUUkR4dcctzHHpY3o41QlBCbME5pZTSsPCNfAhVRtP4iE6eZ
1qGXRfDy55p4ZqLVCM+okCGWOz8trkPwpYc0+Xvl2ci5H0/J93w3xegLqxL0Au02
+5C97Sq3Vv7HcL8UshBpaKU6q7iSTBQLESOWizHq/Rh1EPcNkCQ0ckdULwvQclck
v0DlyE2OM1wtgdxifIZ8zlT4MwX11g4OOAoFzKqmQjxlh0+6EiyCcgz8NENPpbeN
mS55CVw6Jq8gtYONzvy6aDYXDVROOtWkatEj0hTLcn8dLfTX+fyV8o0/LadVMm5p
v8xyvRqd9ZF2owaCujxTdd7ZyG2n+fA67QEciq8za91ILjzgr12l/fN4SOtx9Bv3
Y7bRpdWci6tc32bRixmiaRJphh/upZ0hluuaSWtR06DnK/bwBWMuz3oIhhAPonyA
/nmM7WomSW59j7iHwgkNEay/5MHKLc/nIoA5d2Bg1VNla9eyT8GAKSq7NqKYpTGQ
cvqcKJGU4M11+zzIiCqRrRDtp8Z4akYletv6/tehB1o/vC1JsR8RH8jFCaT9SVXF
Pf2Oo8kLfPqwPNJfOpDFfPXP/kfh4C8IfkMfcTg1e0NSZPAtlUHWn3Bheqg/W93u
B5JzJwYqlrSWJHZ4fpTdauMzQDcBVVzh+WEppJLYDM+VRk2QS6B/5+4EDHqlXAe/
Rdfo2ihZUsp6Ott6YYFdhdALiropKDWtproBTJmVCpm37f0/bsHg2q6Ly9LwvSOW
2Nk3Wj/ZxdQBs7Mtk0wSDmoo6X6z2bA98CG8vp/ZWG8nzRZ2+0YV3YhT5Ss3ZYvb
G3HpcqsMhjes3IH+yLgRVYblaYC9ZyMhJwZFcUs/f1WNEDUR46x1JdenUKyO3NVa
HHWCCK4QMzldFeJ4A5VdZcVR9mWx+PQtM16QfFllDRoQM6l9jHvk7kbUQI8juzTh
Re9IBwOMIX646PG6p7nUVOaS+tAq48xlSqJ60iFdo6cK3lvceBA8nyQsyMUhHMMt
8gpX10ZSYxirirSjuey/LsFF7cT52wue5DMkPi4FqFOoMa3D7YS/TpIujnPEfqxh
sjtMYoOgpE26OaJEZGCxcmN66q1+HuegdEkp/UIzMNoUv7/Ap1rydPnPjlQaU0Wl
P6quyBxl2/5OPqUoDP2JYN+vKRddWEEQe3ZlYzyl9bGKm29t6tVw74FG6vHkJnIg
H2gMM4WpGyiokBQwsWSYZEYoD3RiRnvfluVAW3F+1lG7+Y75w+cjoyOXm0X6cWIZ
BZkUBy/eLQY1DK+12+kHhc3dhc8byBPAi+5qd4XgW9fhbM3Hrhf/LCu1tBXiLRRa
pu7GrAWALQiCaoR+thzxv3ACekfDr1rfe0vziJTvIKX9Qp41zeHUTeOa1XSPnhXh
+/OEUPi8NPQ3VJ6eF5MvKu9nxs1G/0noTrwzLVnX/Wy1oT/sYNillu2CNoAZYhMd
mm9FwZ0K6qF8g72k9h7FulZzRFyQGbempfxc4CokH/+IeoEIbYPFxdpSJsHAVJ6E
LmRIYorbA1GIo2c47314SkSNS32OrWPVgvyzmLHwm5HsIeDG9wglZINCKtWqKhV2
IcKlvAE4NzxgNOE/oe3x7QsB0H3u6E8POZWUyiiPeP0DKOqkc1lWzqWGCoQK4Cii
bXQbglit74UnhDmAlkFbO2FIHZkwOgLEegKicB4t6QyIATnu1HqTU3YVZObZaxM/
DSVwvClNArBKAo7FA6dpow4nFWmx2HKJCr0t0KGOsqzxiLeYGioMRn1d/x+faeTN
TBYsSSS+JF4MZWXw5Laz6NSj7YiNTJwR63oGWZLvZWJ0/9fCMdIFRPxlpd8GLwOu
uR5grFfYa5v9ehOV7TM86FWd826pDPsiyRsPMiCszD5tLqk0ajehLlvZE8B6c80n
jEcn6hq0ZnsimZieHGdA+VIUvPd3AAiV0fMFzAtewe7fcD+Ds+4nlC7d99rQnlVt
o91x2Nqes1g7SpE79e4miIa4O+6jXWYPb++NRPVOPIjFU2AZ1fOVmSuUMGhVAaqq
7GDKslIg3zOMiFjEny7vstXRizCUv0Bbct/6kwcGB4kudxtF3hfjzRj05kwLDiDi
4n/QgeT7QcRPHWiSdwGnZx+R/xn/gd9D1a7Ef31uo3AYR296aqtIOhul4H5bdyHc
Jck7d1yFdPtO40k2ECsPb+PJQKM+TTNSeF9p8ntCnjUlDhzycF3yhSpfRSn4z0YY
GpPeagaiVv3BXAG2+97GRqhscGn1CK/JSDonCHWIpHXSrMT4d3a5uZg7YsBRqn1z
W72diV8mLWJVRp2n82Tzt8FL6yKJulIY/bOkRfHZlzR58/igpgiB52Nn3p/cbhSt
O3TwC125aNLHHOBWYst+0cDDMH9nUG3hB0i6FCEIEQVY8bvrJyvUCxVSt+VWlCQ9
H2MfWMB2YfRMyeyBYsrixBXuoH7Wx9gbzwDIarmj2VGDKaxy++3WeLl03IDo8VOQ
ZCfPEEq413UFm15AV2rTydL6YoMPcpHHInaBI+0OT0sHbKvwpadcgLfUIrBbdby/
s1fsKEB8nUtspjNxPqDj5id6f0B04B7Ix3Tz08OVIWDki1XXd6HWkg++V6jdFF19
Gd/foFkm2Fg+h8H+I8rMWHTIRog0JT6rQWURzIsAmuGmsS9e2Sbv0F6AezgUt+K2
zX8JeLJIAMx7ufQqdmaHqDd1Ay4tCd8hUZvjjNxA/azmmaBQUnEjkMG5buZolySk
gQKq3e9kb9h5dsSQh7fjPPePQ2I56vkonBa7dRxDzAhGMwoCLAKJ3KrdsQ7BoZi/
5KLaY1scDRc7iACO17sozA0VsWmZOb/bQyhJObqK5PCLBKz2WEyonJuQO9wq/cTs
HcfkDBCeav1OQB0gRsn9BBQeYsfbtJxo11bpCs/+lViuCq3qfENyI8xiapCP3xZz
wIYuw8hUMy7LhKUQEQ3OU4iDezlHO9wh3ztrYzgl2jefQcZG1B8MV9xG9AFJk2UV
4QebiYQCi1ynpKMVLwAInglO8wovifur7ocjaBkN1osf5FowszcSJ6wUJwJNAW6K
36j4zagTbwCRGCiDnXsNG1HGuCZdKiIG7K1hWDKFAx9w9H3PTw9IRWGKszikrt46
7HOLzPwF6ZtfVuTYIay4QwjdUq9zExCWvgCD2kQo4ad6Vm29fBqn9zzdz41wm4Pp
lxA3VsE7cxGRGhg3DHAe0bR+k5j4BpnUrW+RGFwhbVd+rvD9ewJTDePhnhc53hzP
HnjN4hTLRgZOYHl5oMcrnk7ydpGdCSRQpxf8KGsk3aylJ2izJnc9egBYYSL8iBY5
aZm7N+7joQn216OcIG/vpBTUAMbyMZL1DmlIXJzpQ6uMZO/z28BUpx0+rhMdNg9T
m9fOGmiXWUgSvJU5wv+cjyqh7KOmCdURTD+EelfFOeH/h2uB8O27UM01LGwhxers
sBtbhNRmK5EujpTyiTS6UFGBr78qmi9C/2h+72+dKO1swVBPK0ZmO+em7wsCoCgl
PnOq+6ngJY1QEqY+wj4j5vD3LAuHGtHBszk3uaW6c77Q1B36SbPqDJiE2kI17S15
RcQZfYNjPOSmRudwAXPC+KRp7Wy4bmFVr0+uyX5S6aOrxxEQd2suU0UZSA8MsLwS
71RLNfdkwg+DqwraSkUEB08Vfuh++s0GQvlvanN6+VYDZbS197TWOXx551KcR/Yh
qF6u41P4rdps+Zu5YJGS676SbFrEiaUTtvgkcZcqsMWBj0duegLIw64S7DxOup1w
Hr5TW60heAXvsO+r2b10hFyy1S3tAI+TtUXrfjwr17xobILDXPcHdkn23QuOuiX6
IJUYQ4MD4irZ8nC1Yefe9r2zBaaB1NxJPGQreBIOkm48ts8L7o2o9Q0/uqLyJcaW
Ec0bc6oTMptBkTK7lxe3DHY/PDebXCyRU56Pg2/7Dpi6Yy9lNeYx5/cNq2tLs+Nc
5YDQtwCZMTNNAolxzwzHhIqP9/xFBuJgPu1QnNYJk/x/xLO6kLlyMpQEGxq5EzR7
ozzA1rSBxgYhOriMG05XARZUEWveYxlsG0aMcDn/XsWS/gqGfEApuCuxB5fNk7Se
C7Df+pvTFpINuyzB6cXwjB4tVB3eALAjBgNXsi97iC2d4QgFmbneTytRhydJ6IgE
h7S67rL384CtcHmGPHhr9dizdUcCU2nEuOzLr7sbdJcSvCYMFdGhsJjhEMhUR+YM
7GBereSV4gytJTZ52gwuqVQ5YS69DPP/74Sp2QrjAXzdwgawdM6TAkvF8mJ3cTJx
cC61upnXuFzMvz9JYwUl6AMnnHmZL7+74qR39v6mEWvoYK+AABOqOybRKGedqkJd
DmitC6neGyGkB/EBz7WUuis2+R1TJVAoaBx/C0xnRo37PQfVsuChhvYoEUfZa0+2
hyj7WMWmxM3SjmpAss7Wxpihd7sX4++sdumD4f6rIJZjc8xvQDBEjUNn/e/aDYst
avkEBkvofTU1Fh0gOO1toDBBGTVL3QznKbt2Ug+okh90A1JkO8IAwx4VoHElE86v
lzhzWm3KQY7N5VL/pjSpB8FMcLu6LI9072I2IuzKSNXaPSNdtJfxIvacenFV8Ya/
L7sUZux5u5ONgAC35/1oiYlXl4FVjxIsSNmsVUgScpqroIjGUSI3zxcWtcqd2z/1
JdRztPDI/9YDnf7h7NG41MG58gCCjzRvU4TMIxKp+kVJa7xBPyUOkFQvhABoCMiE
TuRfvqqT43v+l6K7mwokAo944h7xsEhTqNZObAdauC4ykhby5K7ZcGyrSx9JfN1i
IBjJYtp0b71QA+MLEwV+R/TCDeI7fp1VOoJzNKWO9wpSPnP9ojh2rG+9G2YSaOAR
8lqIfMy4I84zqbIE0zZGmmoOw6e/j+bPLbydkzOZILBbzNWjn9l4MvE1JOOGsdY1
Y9+xZ3c/xlgIzUj/0LZ4KUwECr/dtTMxFyu6GVd2xsV2pRf0qwOUbltt1kjC/r1m
81oGKB5Bdx9OFEgiyhMOyheEGflS6b/Ww5PIp2g1LMCfEGOLRGBJwNCJgga6yN2V
YW7Mg36TxmkFbWDc7hDf28vdP0m0QcfVpqSsSx/e8eaLzJ5ajWfP0rc9IwlLMo/1
KHLEKU4Zrg6jRiCg0o2kIQtJto+bwo9SsJDrGxmV6Q7Qsqsrk3/GVu3BegLNcMoO
iC5CuJ3BeA6cmtmAjqvNWRBu7Gbvi+3Oljx0NokMVaScm8TCFiuZ3yQs33QO7PNE
75gpzqa1LhHNwktBYSrYlmkrVjHa+Bdt9tD9phxBZbmarz3lEINtFyTfWu7zP9K8
czmfXt7of1yHfcuW8SJtnGVqZ6RALSEfF0CBIC9tGaqKCLYpdCxNv+/P/Ha3ZfDX
Gv3m535xaSihH1caKxEfy9g9sFuWgQ3hu4Xqa3MHLDDJBuMa27bKx+A37GO2SjGP
L9Dav6OBxBrzUqpG69A87SSdiWF7YGF/yrhetXOglcXuV08zvSKF3gIWLtASi9Zk
kci5ovZHsgSggQwy2FJ2gMSH5oV2Utv6kQMyGkbhasVVAOqCYEvjT/wu6zwudNlg
hMC9D/ytPAQ7ltBql2F5k0jaDkSKswBCXGgys1USItY9z5/P75ah94NNFhNB0psj
cc9SbErnW15nKR+4R4LWRKMsei+v0JCpo4YrEu2IINceBiLVuqSoR/zudR8NU4Mb
qsY6fC1F8PHApVTGIdTgkl98kCDubLDpov6EnNi5/7K82oASYA9Sud5uFtz/BEhE
N3ThVNECB7WczLVF9+kf4+s5aUi7XpOhK0WzsQdRsMLmrJKwt5qQRWiT4lEuNrsT
bIxEbr13XqHHJmzNODusSPyLto+j/NZ61JthnfogITy0/uqCVvqyoJMpEyXv37Cf
LaIoG0n5sE6CZGup+xHIXEeOEwAhzO5gTdIqY9Bv2wFo1jlnnUxPRKHSAs6DSLhZ
AtuL+yvMaItc+R5eE1knazgJMZcrTc4Q/9A9CaqTvHCcgrxFps8QJztdjf7iM8zu
ypRKd33Fxu0yjSmzd5e5bEB/+cJxzQnZr0BnlqIVC0AnQX6lmGygc96Iniv3RuLE
oN5vKaznKBg22OiqjOCkBPtMY4M7dp4DVGOud9IslUg5RfyB2By2pjd/+Iew0Qve
+ixufltjG1/JirfnV+FMkIJWyHRr4bc/smsohLTTHTJwDg/fY2rJRaJXXOIP1HrP
ZYYDMp5mdJZENUltuXz+/pjK/B5e1mV8zftsdmvjWKnbsv6P5RNR776aEVOSqYbG
Z8vn4LLeCDtC+fPolAze1bxk0cn6Wy5hjHlVlY6LQMQwhMRO3nxs9VJBvaycL/bY
9zoNzQaTXVLPPcwWaQySte/tQiiutc6yEKhxN4kZ/hqeCPNPMPv58qo5SwsjNUYz
w1dczCoQL6BU/FfL0zJ9kqo9QrJVYGl5vC+CAQjE52l3Q8SoF38nsmjDVdQ+uz8o
7R9EG7HuO71tLxvXh7/pEnDjpTnM6Cs3f48w9zUBhBMTjiLmbrXavY0v8TtEMaSQ
`pragma protect end_protected
