// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hYYDYhfGV3QqaTMHAeIcyyeuNUxAYbvI3C8xY9X2YbuoWpsIWlQZZiD7uX/ndvGz
KdaCyv+6AHCZOSClP70gaMQVmfQ9ls6NZ3AfBrVo0qEoENg+zdyP+q/WPwzKSX15
LHx0GU8eajoo37hU+bgZL7+31htJ8sV+TfpSBww225Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9056)
4gvHD+9HvVIu446dyb3LOrDwalpElAwrkg/bxVAY79IIVu/cMTfYWs20248O78Cg
rJPP/FNd9YT+d+HScrJVdrMB9LMt5Reb+dnNBUI+xnjBZA6fNYtEQ1eGPNoxYpKu
SV5u6vhO7WWKQr+UIHt5/tSvM7k59yaeCSjMNjIjEkjDyfkoqdV/8iKZsHxF18Ji
EKvTzibXwuchuAJp+tD1EIdmFIkDsy7zf8ZkvgnHwGyrx2FuvRjVtjV8U/ncYp47
75JM2Y1EtE6mKHabFo7PoUWYDujkFnZcVwUZBhfrPLDnni2vcW8flbCOxJvTkZTH
RJB3CVPoH2ttbKsUvP8mBZHOc8FQDKIZuAcJT4ogTl5ptyY7X59SLmRN/Zt0LvmX
uQES+WMW97Qx5UCnmYxdK9QaT0bXVhVpc4a+fvYqzhSGTm8C4MBFHXsbgSDZ9+OZ
R/5cDqlJUsokveVnNQkM9tp30hGH8ody6qJOsbWXzoGvOnevAvKOvvQZsBJO3a6H
WdSwe0/+AXuE9gTHqC2GNWmYFywt+L9O4X0wSMO48VPEDwAAGa+rJOBrrB2Hnmiz
56kTqSnll/K8tQ0ahAd1MdCUbDwCR4cF6hG8dMXI7dH+L2N9cEn+WGu+Gdl8KTcY
ZHMpkM3ay1wBqPEg0lS2Wx5b4srB3F/rg8IEt0Jqc7xiuBHQG6qV2JfYcGvG8L+W
0NDc0v5MQNFMY0oD7Gd7NEYOO6cxInzHo3fHYgRMKNhY6E6m29kfQsXKqEZrL2LO
r7/kLsnnN6AfkRPuKcJLlUIoGRlLTxo9N41FirzcDPhjPY9lp5ar0dCoqKc5ZDAz
UbSYgE95DZeDTpIMHBCM39SPOlYcN7lnp15bJv0JehdFjTn9A/Bf5BzMbRfGm778
DVpI7Fb+oi0Oskv5AiZlm5rMb37Dtc4xvzeGRquhhE+hWuqecEQGRsrmAh6C0o6b
cFbTwR9Tl2ORvzklLYuhU8Niuezsm3dNGbOwllYTI8pWFYdOBtScXqN8ycM7PZqn
F+e2zKJMyTmUmidCow2OHbTiRg9WF9H7iP3ie2/ITXeKIGrpQtSLaP0d3rtFwEjx
6vgis/JeojU226CiyZnXeXD67gy2q0gCK0sLUwYfaMVEteXJdAei0SIZfdubMncD
Oce6CYeKbDGhtX9LwMJCtMgIZym0iVovkXIemdUScSHgrzB7glKiWdU/pp01veUe
SW5Ta3aBORIDC51YGyL2drIBbWIF9SEjzEYK2gBVThX3I68JI2dVDtL4luRwl9JJ
UZOc0NkBNP5nbWWkoglI3GVWPQdpbF3oYTpNLDeqHtqJ4Pwqn3y/T7DniRkuEimk
cYV2NsTOclmTydAxTsbJKyeUSgLRWvO0Vo/aJthsYdMxvKJsOKABRX2HFkCl11w2
H0ToefY1MH47swh+C4qE4H9Na/MEH4UH1rv12PYSeM0cTPrf/ye0AlFx2YnlTcLL
tuhk9byXk0riXNyODRmTpVcA8/aqNsdUs6evHMyhIhKq0VSSd3fRwoRWSLl+ZHxT
PX6v1iszsU4NDPYCxuyo5FhDxlqbZvarzaPYMmr86drf7+KWC1Z2grPBbKDVtWqF
pH00/4u2HnN+S5g6HNSoenIJBNZe9J8BuZzYt79mkkTRkpVgNpSmp3wpfyMu/s2b
HMnarro6ouM3Cnc4al0Rl4Cw9h60hnWfwe3mI+iSgBkWzIeqf1+1Aff+zDUZqGpX
Bgdhvjf5KG0mRsbsAavqCuJDL4q3PqwIik+qMK+admcwXzOBfFQ9HjAZzxr9Kqf8
BznlWTlfZ9zM9x7/TVYi3cb6ZyYivC6Zab6G5ZByhPI4BHG85q7AS+N+CcP6DDdE
4MfKu9ia93n09Mekv2TKAT4/Bg/dmtdY4nqsSHfV7esbCaRV754Zrd8W9Wdy/URb
qQVIvPGw+umYFHHSHj9RfNjxe75omG5+Fnbx/ltZkjzR11xlcNbqZT5TEn7Wo2jQ
DLnH3kAG3PFVeJ/23/W9W7dgzI60650WW91FUaUJGNCSH4GHWbcSNpsxJpeGj2za
oWindQJQeLD2h3U5SY/UHkfBtnKqjt5ICD1I0np0SF1cTasvOetXcqX+FCAdhRc2
GCjYpXC0ow6L+vD4EZbT7Z4nMNuBQZyas45d7WXspGhE18Chr2lavlLhOc21Ga6C
MOkRistbxd/S67CKkSEFy/P4NnkFmKLXsOQiRFSsfVo9zpHPCqBzyxamWYHY37OF
862SHsAz2QQOJtw9sDu7j1UVLHM9irf+brD1za7PCGU2jTu9xcSZCJ7AnJEBoSc1
q9pmk3RxzkQLoX2I7q7QxGUiSXgCZVtuH7gCJb4T16hl8t62Zx+AVLztKkzuwG+v
emze8JE812aNxQnHusDcng3NflCH+sJ6A9wVLJAIFVCVXAqMN1PdbV33awyWB+eQ
aeVOWirZY+SVAvk+Hnckuj3PaAaUm8UPgGuIpOnR1AVoTQUlZjbHfANcRhKs9/dJ
wV54ovJz+i2VhgI5CnerMPjdP1ivRw6JknwacWmwah/AfDbFJo11tSmUvH44ve2p
MzX8qLt2RqDfFT+k15FYCGG/EOVBq8xdMici7QEJtukWrJoa4RGEwcvzxzS1NvRg
DCrZNRiFpDlptAstKrLhcuoKLZ1ACvnveGnr9qtcrGP7voUx/brfOWgJn2gy24y4
bkKsVTNd/7Zmq364MyiR/Mi+M1ZmKLTlRQmhf3F3v8fDcDC6kam8HKJvg+5UtrB/
CU1q73ceYLyNjGrChatpmaWR1nveL7G2NmeTg62mkU0ohLAtrVho9Kxk7JUCvx8s
8Xgg7YeM4CziEWTWGm1+SsS/dDb+RP+XLTmr8U7shty5qdk5N5rs+ydbrWY4PhJR
GI+uJRdVfW3JXjWpspFzucKZ6m2cR3k0Z+W0rRoK6iHtwXaZOXL7oAdFipwXUCgX
jKfsyeYvm46ISb2y4xY0H4HEkexF3x3kSPGIK6evW6sDBc4r/jPzuXTMAehQc8kJ
eRb1ghSkBVFwFPhIxKsYqwwTRvrt28IA0VRv0jgzkWDGyFjvVBSYkNbZZEHIWMKj
OushWVD/z/dD4bfoTmOzvCowM221K8bS/QIzbUWU7AKK2YhlE1Gv7rFKVvSAZ8QM
8+kZ+CxkaYiWy7yLbuPBb0TNLOJRU7hh3a7QfcMK/W7vtkmCSri6nuTG/Da33BXl
4uuSlznj/fDfFyjIr4g8md9HqRpeub7ylya8AY4NJmcmv5xFvMvcDempsvdd1TJg
muUJd+Rrt4lLp5XYHPOa5hjj3OkN75SYZBRIl4/ur4U0OoF+n9/Tl0IJ8l9UnkJz
ADHzCsVcO9EGPR9R440lG0k9rvH/FF5aYKKJCyE266nEPi/OHJN/3fVisKerCDL1
EfkFM0eXu3GZaVc2LaHdtcnF0R/FrPeXiohSoVKXuD3aTtuPb46aCar4BjZZznvX
y0NntaSyqqA5SL5zdmN8F1ycvbW7zwILEdxttvjtrXubgy8+6TfpcezgqU3YFY9c
9HEudPWly5EBtzxuYZXFjxSODqMYsmxoY62BWXjOxZMTGubw53xYeowpsUQYwRWy
84g23rQDFu97oJxT8FzOEgD/8vRRDdVfd6wlGcPBjf3DqNkFnVQwIOtjhA/7cvxq
JKffHU966vj8M/0JAFhNFwGwdEEKEYN5GQ6995aSdVGTp6XElDJlXisHiGOy7mBV
ESv2MYwAx9bWefpV3OmNjW8w6XMcPlin84xlQn7aSpE42N/G1T+Qr3UMEP5VyyeL
Me3vsWp3QBBYFSWIN3O/JNCSz3dNVgDBjDlvGNhVuM202iQfQALITr6sufrgCj91
PFTPT7ZjWHpEdDeEf/4LtsxDhBH43sh4vtWpV1OCLa/fIs6rNtUvdspJM8bwOK9a
E+Nlq0bcHjuyAfYQHSdFBa37+Ve6/bZf4/Wg1UMhPM9ViZWryOMZpD9sj2QNWzG+
Xh8JQutSpDr16suDOnGhWBciM3WzInxyzGOnF36X22Bt/cng7DhsIW+cRY/4VW+7
aWsJAjEbPnFI8b8DHMqL1E2SAKGwjSpPr4MmoS1OrejenSPmr937j/xMGpjfj8YN
MDuoDl3L151TixF4RvtEYs/7kM9k2NJxOpQswIzEDmevu5tWTKZHbdWC9bivqDZ/
PzIWSjtXkB8hiaWKJvqyKLh2+jOKCE+ncRO3kPUAUpOBJxAD6VtDNmDbvm23z9BT
tmZg1ULN3QW6aY4alom6qBODjzKKTTyiq5lKrtFtXADZxlqvehWfQJM3GIeEgqAa
oeq24LGrPkkKpK4ulgNPMvWCAVUZdjGmYTXSvpHVZ8wD84M24kDyeK2yO8zt82+s
qqHPuGIYQzEUQOuoIA76x1zZSE57Z1WRaWuykcND5RqwQGteBCygrMoJe6tsjJk3
vGNqVyBH42DwTQ76lILbsXF2ojDKDjWwJSKvNspBhYW6lGxuqS38kfxES6DVBjNr
J1N7Q463GtZ9IRmyR7vOS31n9S9KNhlnEgOHDoP37qBuUV6CCLPr4DGhOmm22JTx
ASnlNl/OAz7sY87gIuBht+Mq2lw/fIqtldYMAle2BV/K/0O0yAcoLRyWvA8S/N2w
PN0ccrwpUfK4t/vmtmaFYv3I6R802iN+L/MT9Umhqe1hJz695wDhrHr2mA0JFr7F
L9JULrJrBr+QILy2lj+cQ8ostos11Syki3LWbH8ReUo8wYU7xCcbEN0kobAtTs0b
d/xGGauMRMWV6wagPCgrx5+cnMBTGMZoeKs6Jog2unt8hr1ojjEts6pN1FeCjZop
s7CwOBsdk3kH3qWK5Oo89q2tTCnbcz4kSpOMQmbhV3X9t7cPCeaK5bQBaVP1QQ2f
QM7ZGGulrKjubaHaB4uNTmgVyCl9gSS/pqhkwAdsfyWVjcUZaRFiXzTVmVLSLt74
CihIra0r3ICJ7FfoE7Q+JqLbYvDmczdOGQZWn0cIhTYgnumTuj8j/p8GDY54rqA6
m2ZfxE8WEKlOVsoKxNJ1LroRC8u9podxusUEfVHNIww29KJbpZN9iN0TGSud8NTX
gjFaGvvEaETQV4zjYSSnlIBlu/dAfVbMtqos+ACvTHbNj3IBb3CRxM78okUhyYwG
DC9z8FW3caPTphvWuXjVHF+B3NWmJyhj7TFHuRKcb1v5t/Kqx5HTL+J6DyW/WJqd
ipvIa2f2JLKfColFp3fWlxoad76aPK+HXSxFkSTtjrPHbXakdEe+VPECu4c0vPzw
IPfvz8kw+3vbanJmh1otTCZSmyQu4RWya33KzFTrcSAtV+mshMxaur8dQDHARify
gghinTa0FM9RLU5yBkcjPqq2MxkCjFfept04Vb4Ua4GSoR9AP/7PqtKRXm7FSA4Z
1U9446mKObT/lj+fl0RTTbOu3nKkVzVUPxIixb/Jz4gN+3czWfmUPthKrbZeDjti
pXdQMhdNeaeRevwQ+oof8pvxOt4hwtwL+sQvM7Iu2lDljSvKgy+NOrIZBO/MCovx
tdgBD68OmLKPru1xbijg6PTenOjnSgfWorXfrxn3RJoPWz1jdXinla27xtJvgXuk
9limners6CA2ciVbIrRi7FRAE34gM6cWzuI/S2zZt8y8LbVu8zRkTXAnIqjj1Db5
lfgyRh5twIkFm8UShQ46Hk+7i23BgiF4k7ocyY7RUwrYxTbdhbdXMHnbAgU/cjSc
xpkdgsWfuE9ONzUZWnH13Rz4dwGJRvfCwb/Dptat9xblMQ2nq8K04/WjxgsmUcEc
ViKrLlt51JgNuYGofuSO8Ls/xe4iUkZtMzF7uCRv7anmUTYQDFBL9afxbBEfZocm
wuXlFyBooMIwgHOWGGbqg91DHXGTC0VVqDBAR2eBd1u/3R8aNKpIPkA+yYIjQ5Wt
OWR2kQyjoKVxrkTdMeO0HKhxbLUbibDPKDAq++dRJPH5fwLIGcNUSy9IRtWMnkeS
aTWy5dtT5mpW+/fT6voL9iV/bN2AGd4EgSuPoUC3LoqYxmYwFMV78jfA1gGEcdGn
L4W3Qpz+RR5SmZqMjqnrHGTFVYNagmgBjXRmYn6zkG2VRSlD/C3ERcWe6P4lWVMm
PMOzWx3LulW5bjB95TJ5kY5NBhvMsE4X7XnxeQYbH03mQKapWDkzLB2xFypboCMJ
v+8HRav2Sm1LIndxQ7lGVaC9EyKlI87Wxqfcop2KFLH8DfvXFeRBc3TQE1FdvP/5
Zz9Cb2/RUORUhGdKY0TjvHQliPUunyf0/R2fq1GimgrZhRb/kBYrMqb0RaaWCpF8
RzYA4YQmUgaJIdOLwEa4cAhoWx3hLzS5bE4qNKRuw3asoIGq0GWBRPfrzZ/8lkV0
0AV7/tQmUYxi3Xmw1ccNjIEyPDaYGuvoBeBvhKbIvZEQEiqL6COEsZIMnP0CMxwz
AG/e3hlvEP30+9HmzTAfr4zyXC1O+aFy+02M6GE3a5RZiYUGgt65a4i6aKS2UFKU
Z/wbsn7f6k/lQHlQYKmXrEm0waVj9PNGKjvwReQG7IdK5EkIOEIrwnEbIC1vDMdI
hl5gykgvdtufkz4evwULiLuYX3mtSV438pmF87DsWCCy5UjI0VhPG18bavnkkKJX
d9srgp5pLtJoOw8UNkZKEfmg2NUzXQuzT4RwX0ER2O7nzhmJykW1CVxqkgv3Gljr
5ph2d9ytnHvldmn/SN3NEqJOOD3csJqd27RUX87mX9y5W2K7696pfAY+cNK4Jd0y
uUkb8Xk7BAWXBhfsv0rOekDiNzjmshRMe+0MdY6s1c/NahsK/1I811nfT/5eUPpw
wJ8XlROaKRzj/36Jg2pqSbldeYM2DIb+EPQxotWHIJeNQJUXwip5T84XAu/7FeoM
SPUILUanOcQpoIFBMIP6q92h5sZkACwp0TOIw+Al5tmWBKFWBy3nnwwn+CKVI7b0
BRG3t7qjFvX6GecvT+TF/PPFnkI31NDFtJPyH63KoKoCMFJznb7yUnuJoFQIFpHi
2ONnpzlpHj+DowtNmrn7Bd9sjj8Dy5jbDfNTc9xsf9X75AJkVsBAfN5KVdIgNYiG
ZIC6OrY5I3ahDsqNVZLcYLNVlI8v9IdLKD25yPqGcsGrA9MWfpsiG93JtvtnXU9s
XlHQkjba81p+DU9M927CsJr9S4+B+uNbfGQ9wt+NrYSIHgVSlogg71ZVLJGv2JP6
cTrJ7NXGxBjw8FjO+Ex0kmpZdIYDSLpT7kmQMKsOPTVT9xicKdOZPMfZxsyo7Mdr
/vTJrtg4ajSQ2Zx9m/phI4cxqEvsOfsvWVgBivIOhQAYMoxE5/rLRxsW/S0iVlat
ufJme38t9Pz8cqLzv3vfyEJkir2qPEUhSQ3jrWJjHWtxzANE4JqP3JoAj9RQKCE7
gWPZMZez3ymTsXdVPmaBxa+ZzNiZOuSXp/Q9Dgi9Ul20HACzKcfVvkZOd+9t89/D
6WblUKRLdgJA4va3FxC42dWRdEUTCdr6OldaRyLMzcI/ChkbdONpzpmQm5a5WBNP
QSG70UEiEPHLWeXPa8mDQrwZDB8cAxD9tDmcyi3a21zJKpcxLJi4s/Okc7bnPU9h
cDlzoN33JoqdddDfT4o6+AQbPh0Fxg7Dchh9hb1iyTdwA4o3JpbCu9EZM4IIshJg
n8aqdhSazw9i1UQezk4eFTkcKqkSZAUWTSrVcvd9fueKcyjVzCRVnRLM6E3Gd9wD
zc1o0gEOXzlyRhobiQrt01pEWcMfimSp58dM9ysbiBZe0nDMTJmv7K10hFxL3e43
MWQ2FU8jbAQtX6atRWhuNEzx+PzDBHuFUdDl4Q05n6pD7n0m2Ocfn1zrzmGJySFH
sE9VWnWic1MZycMCU5inUzRqOwnY9AIUyDqEa1mfLvr+9+Wi5MqSPcO7QwLhhiPk
ov+GKdtYmE8N4Gcirp3LFm5Hma/zaOZiJSfLpxCW9b1Ls3lSQeSGrdRLQJvFk5A/
+0wDYVGox84n9PygKNaJb9V90QCjDGSWByBcTRxESflJKRg04rKvyAM/aWVSfTfy
021R1Oub+p1WJVUyjXAn9so5hnSrMDiWF4rQ8FHdQF9aq7F8r26UzuNNotsxMwDc
bncvK5aOd9wMNSR9Q3mSmZluUWizskABPEn011o4BfXoNL1IfA/Tc4edSwKtVYYD
2xfwU/EpAGpdRNZgnkcxZ4ElmVDLskmLnRlyhgrIYLLR0yW1j1dgQ/4bfCOhVEGB
ScqS6e5zDJfGS617hmEmCtWwNsxOLONbrRYCeVaQLP80eB+icuIDqSA1SCsQC+/d
3Q6qoqJPtp+0COKwgQqf+UbtFXb+asZnRFnn/XCuBlHkVAyk8F0ZIXyGBfZ51ZWZ
1FK2+WTabjQVoe908P2vtSfPBwIQJ+9875+jNRhAJwI0zKMUyxC+k0m20i0aKBDA
TbsV/5g2/Ib0DYXyuieRYQe5mtaP/O/7ngJoVdDQNfKBGsxBy03Qjuq5hL33RdG1
Ph9Mn2DvYSKM2sf8Nl+tufk2yaOVBCQJdz/GAMTLtF2ucUi+p5jIu4dpPsRQZKUd
cyuDjkgQn+O454KQogNh1Ir4c+6QHwFw3p831JaUGS2e9jY+SAC2wV3URIdQ6qW9
EINzWM11qFf3XqBbVSQMJkUu8S5S6h/v4jkpS2vgAr8jYo7Wg/JVvsiGQSWMOl5Z
Jp7d2KQRG78qICZAr/UE7zSBVX70ycI07XlfeqL+mzp/cNAdDwSRS6vDZ5Wf5XwL
JXnqrDxQ8i06Jgjh4jF/TajXMlto0FjjK5wnaZTT+RGA09aMVR91FvFRp4P1M4MT
jjBPZD/tyHUzI1KBqSAklpE74pwohE4M18BCEZI9FeISNRKQSr7MkG9SAqC6Ksmr
AOC76Z8Uc1kzHHdFEI/HDa7RHrTrhAEv/mHAxYxuZ88mt9Ij3MUWYRMRJBa9GdQP
MiiaBIvsv9pWY8Qz+rftOAmUYBYTyrLV+Qh8GJeNAaSYfSGE0i/b8xBHuo5yxe1I
HGHzRarf4ozmg7HXSO4DeiOA1ctN9k69TiTZ/AxUYF/eiUmQRIdsOvuXcecwgznb
10GACMsegV1R6r79yB0zuerkohzCDDgUVD58l5LaWkeOaCV1ar+ZPKHN1PiuUcX5
YOaoQYbON9Adq0tc/cxVfGU42Ydq8GgpO79BWfq6IpXJkLOXkZbyioDsinB2ULdz
ClBdRcbwgGixREh5NH/bvXEWo1+lfsPWPUCZeT7v6BtnvRI94/HG3+3xh6h4qiKp
JFW2bpzWIXsFIq9h7DNdM6qQG1WXTd77BdBZEtSu3OX36tcZkBaUVzT8Ua8bX4yk
GHTh/gM5/nKSx51OKPUAYIKmpt178tg8FHZ+sVgTovfStDJtmGkgYcpUGpYjDD3w
duJiIa2yamX1qXQAGNa+YuwJQjsnybylMJVZxW6jesMDJlFQGzRIc7SEnq9ee/8E
dLG8IYXGNNg3j2JpoWnAbLOqUnnVUvtHR6A0xsj3YH1NFTO2CJa6mtpfZiC1f1IW
h65HHCZ6J2KrkgLUuEOcfR5jF8FY0F2ed6DZlxTxaUz0A1WuNd2aQECc7HoX/ORi
jRAFrHck8J2hueNsOZlEgkQ3SgKwK8ZMtAKmV6yRzNGX0HHA4WQn6GiWcUAgP3v9
g66M6r+th/CQuVcD63/YsjDQBSGIbg3epLR6YJYLf2kxq5BDX4VBukB+1npZphHu
JSKbq+2z3fgktCU1H8km72xPeMb0+RHXXBvmoANA/K5JI1yKRBsv0156DrAj1okS
eclKWG1XcwE08PDss99L6YrkMyK3lWL6jlpv8Ch2jCwSekkfpf0+YPLYr9gCCLB2
Pxarvcqc7P9YzbStQnswknOtWC5Uzy9I395aL25ZGjXxng9qrNXi6Auy6hRfOGgw
jGW/2iJ4L12HCTLE1fZW+vWHJZbCA80JIarBh3dbhjf3HBgiY3SYd3MR1z0LpSKz
tqGfOE9LanwOzpsb6WX0KpnMQqRDtF4VmzsONbPKn9m9IW1+6qVgwJ0I8BdnQ3qL
WpnZQStt5z2qQ4KOz1PQoDwYCqGsm7qVkKdJ2zzeADDk2/eE4lriu/CGwKU1OB8H
Bp9ssrTYokHuPt9HJYf1P4k8FCIq9gBNABenA9qHlis0hEM1Y5/jJ8vT5tfKXNom
si1oizPWRrOuEgxiZcZ8fC64mUrdJgxEzqWGBHP57scZCHoW/R1j4bBE13DdwZsQ
aF95Az0vBrDYGjVautSekNPmveauAbpxjiDm2h+b+Dbl+5CZyu0+N5aN9Etn7yQX
IRiNbfBG1OYLapxB8RtrLSco8mtA72BnFQel2vuXeLTa1I4OribEt29hQB/Jd8WQ
B2pnXJXup2nUYVsTw2vlXlUtiRquYzUz/EolTCxD7nE2cf6uEZXDsqyyQtukXhl0
gImZRWeINTK+BAJNWvEM3sHje1/oOI/52ZYDdBdxSERIqv/jDZ2+YYczf+jFDLY2
hevezMpxa9JgNiIOaPvJBDMQeN4ysQpBks745oECIb6cCrR46hD9yQ4Wpj9jDqnl
c/OhioKZ6RuYxUD3AmmzfasFrhFPlcoif2W7bsqnZRDIl7yJM/TQK/I7yg3GVwo/
iRdcWsC9w5MsKzUumASEb1bKhKsTUufiuyPMhEK+FQOrtOybVJi1rxTicUiiFVvP
/EwgMy4glKKlE8Q0xEuCQE0l8yeEFHL0m09KcFo0ZB2+5pdcnHA2oNobT4o0kZsb
taOCNuAyr1pd5WylLttzfaXhElsmZMcNqNy8ZLgGBN5D+5Co0dQLoWoKNnyK/+GN
XaCRmsp44jAbUEOZ7Nycr7Q0xcDDQ3e7rYqlYjx6mqn8iRJ2gcUnkjbzN4PQanGb
AiM2SRposm8jn1Ck/yxQx6nr+Z7xD314GGLbkk52uDNZz5bG7+86v4Wvf7sa1ftE
jGFjt7LvGH2Pydql5Ibq0/aRrZczRyp8fbwQfQqBuPfcC+QgIYvu5DnJsOlNC51l
SwPV4v49TIWVgBOuw97VrEuSML4cSMUdoilE1Zj/kEjvtMRMti20VbRJNVF4Euas
MdXve2I12EXDHXP6DFlKqQdVpIJvr0kYCMOPAUcdScGe9A46KxJF1kDrYNoxZG1j
utOWB4KnOh2yEb4+JeXNucfmNEa+TXzZ5RYKlB2GNwQf0tLXKatMyRI4G7QKWdzn
/3sIS8b5FlxMJ3DQk8WC5v5AVdjUBjtOc+WLnY44hujz+0+Btom0z+4/4qf4QD2y
NEvJZHkSrCbCCCdu0GQaTVM3ED9mDs6kLUOQ1T+cyC03mIaVFPsVsUOrbiCT/rst
Ngx9Ee4CgEbYSuFA4pbwuk3xXCEK9MtqvHU8cVTyPq3g1OipomYoeshUtNpc3Ubr
LWgE0dCpGWUNrPQf+LoRgx622zXuB/egA/HojWpQxqE+dw18GO4BSVEPDP7c/4o6
nbaQbZ1KJ/64VWv6RZ48lxPKsbl7wjJe4RuHYgqaLIV4VNOMrgwgLFoXuXSu9KpM
dX8Ii5lrN2ayB5+7fkmftDUZpU61NOiMsebDrH1ktfdfvcS1n7g3ACETJGSyGXUL
Acu2DbIqYdi4E3uB1EZ2a5x2O4PFmEI1OxDoY6NoRNCzKBRgbVV2kQyZF+6W3R8V
SApRQlCRK7ordiYaXcsN2/z02gjJctYHOPvh78HuPbZwDVWlg0WAd5nl4LrYhy8h
s9D1GgmUAq5ZZqJZxj7qzS/2O9WGTnz5DB5QEw2LEpK1QH0SaHLfPr53fvo8VJof
4QZTYA9jcxi/ukgRRmyzTuh+3ab+0Uir7+q3QSKHF2XSEq2ins392VhjYgWCb2lr
WYxZWntX56nBp+cl+5sZTqeTIkQ+PIu1JGDzc6ow2Zz1KEjI2xl5d14LhuvefDF6
oFnIC5ZOUZzEkOrsDdsqzaCIRZa58YAybIrRrqQaE0UavLzg3fQFzzDUqj4UHLY2
unvsNTaLgA/Y1j0jUejKs48Anowk2//JLKEudYSgWAcIdDkZjDN4P8aI1JDgXXCz
fWA/5D609MNseibFSlQ0OeZNqwzbDBJteOzM1L7owtZPthI6STtVEmxJg8xczunx
eJJwg0XQ+mY6JS4/slPU9GTG0eXGIX5NTUIrA+IYCqM=
`pragma protect end_protected
