// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fqy+4QwIbmzHZ4ri0zFRUJz8zt8KtZWbrDTHwsyQO6V1GPlirnOdiFzVRkW+fMBv
eKL+ZdmDImM9PCCQy4BfvBRZhdn2IifUeeWBl5xXXun4IceywGYujEgGb4nXG+SA
rbdoXbpXKMDUKD6jlmgouaA2ZfP/1gqPGwISRDpnIfk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 88720)
NnWGg8mpE1ZH4HNC/J8vNxlVhdjfQgJZvZWmMzprPGIOoMhST2bU6CY/Sx+uLsL1
SrDGsqZ33egild4En8paiH3jMoNWs0boNe5wvA8hixZY34SnasX6+YWYX27Y2bc3
QTzLO4pRFy6vy3lXq042fyC5saszQCGX3ssR3ibm68zZYB7Kr5GfCfKq0TgUey7O
0WRyW2CUQRxCAFVg9pQasFQky8em7EkvuOc9xcMMmmSX2I2D1EDQox1DPCrioJ1R
dSF7HFEf4QMx2Y9d6Q+y36UDzT4QnNZGCsgKxudaedngTPCgt9KK0drHmp3kKk47
aDvAwh/8/ybvmaR79lNQdQ7QELO82U1I8UrDcRPjS245KEjyXdO0YjK7j1sOD5MS
rxybarrV8EIkPUw26W+Yeuyv+YPAJ99Yj0P3rV+re/CRDmoQRFXsqC8gCWCOscQn
7Gx/tOtym7LDM/hQIx2812iw0OemF54RNx/IfX98EVJ0p1kNo6GEHx2yn/u0koiW
+Vl2Nzn3AqiQCbMICGirllO2kgX0+JDPWY01dPajQbwjC88eLQ1OMIfhC3KBVMCl
dHS7dc88Xq1OD84BqGK+0TiIRf0xHlpHAZpEgClMGCVS+Ohp6fvWFSdmgGSbXHTU
WMw6usMkPc7wfGQaJFU200+vu97v0K3Y8wm4dFP0h0eV+2C5/wOQyrYJUu+rEYZY
yOjQfZAxYD8wUyUolBtCaNEKB6aDruyqjvDgEU3GKk6DHKK4AQiAoom4iQgdDQhu
vEt+SpU5TnzkaI9T9F1EGwd0L71mYrZ9l8BER+kU9uH1FTUVT2AcdfLeVjwuVlOt
A1bFS25w+ifAUrFmdKtg1FMqnjEOtsr0YQLn8leOPzigJVJeeIdmtzUgxycsdkqJ
VvmjNbmYTxvPbU8t5MYBAsoyPTvPJXoHaCZm76oXYcDl7ILP/5h0Tsl4ncUZ6Y4Y
9U8G2WjrUslNv2sNbSd5SlOUjt7Oe9QWp7wEUxQT10kygZGhB3exL88JkYKmFoSS
bj4IdpIawLuvj+1mIGkS6fHKkPk5QeaLOIu984q6CHnbAx1z7nWzzVtJ459T7oKA
gDt0swFWx2+wOmcRIhtaDd2PwZchq+2fbYG/ghtjxDPoCsVpLlJenSj1s6CZYXT9
NpZS/6AErABdluZquVV76bicdh/6fm81eZpmklX12C6DIW1Bf8lMgjQAuWtbUN4d
XofSB7Pemx0KymL1PjsAr6Bq5IFhpKuZj6MAdtfDvodnUPHSAolTGueb4if0bi3k
dFuqN9sX225cxmNCc+CsYO27ejrmCaa63l1EtVm4VJLLtvK2YyKfV0t9fFWb6Yv6
L4YUlNgMK1XpjlpvHQzEmNE6jeqonJ6DTuA414z7R4r5+dVjqWgJ8nm0bhT17xW/
cZDe/OFIKHrBwoZDIfWnXy8ylG3Bz01Z/GrW5XGyC//NWHR+xxRqJ/TXdp/AAQ/P
6MtP7Uvg/GqiwnGy0JnGolrLABP5ASGYlt/PZLD3as+gQ9K+jX9kwzvVkBWJGWJ+
eWl5gDE0CZKCCfKXP3KpCxzzJ6Jba9/eeqlEG29vUoS/cUdWMl2AHfS6AmlOSkee
JnV8/2On0/tf8Mq4gGWmPUozUN25kvSkgPGkWQPJp/3SmvuEGH9bjKfhMLZ7vt8U
f/QIsRQdZb0/ad70NNfuwzEmQIzW1h6jSNvNf9FLZnRgwAk0Rw1c3s6+09+8pc9U
DpLM7Vat9BBtn5Qw8qLhISttwfDJqtMYIKuLjxtyx22gUisRcNaDF9qDuQ+XKgd8
czKWOqmfc0MC1mv1CZg2rEJFQT1XlrVleouUAg77fQ3JxRAFMBb9zZQFMQEXi/Jk
nB5Uo/UdZ5XCe29d7QM5DnE8vrpB04wE/Le6oroeLwaCI2xy52myYjNvKC+bUXP4
5Jp01vTOgiyk1B80YglAjRrUStyg5htV7BZjcJb/26Ogr+FOwF+LSp6FDLmJLcsb
rheYGyD303zV2ZcLdhUMJbLlB/W/Wjyqby2B8Q95LOBVC/+PDBTQ6Z0jQpALKKxA
9ES/srv9bgFd4iCpn//toFxUx16Gw+xccuOG81fMarQXh6HV4xgoOArKADQu8KJg
XVlvmZD3Sa1LLPPdoIelJgSuN0erCiQ8j+gi1FH3SIj7L8jgj3r3uQ4hm9ZGMR6J
G3WyTNytB9qv6k9aCw43Lgj9o81/RMvGdbCeqMD2XxQ1ZPhTARR7rDJtwJEeOwyG
1YdsVae0GYZ5INJHvw9jtNGpWGUJ0TtR5PsXS2+lUiTa7SVwVFaqVNelG3rII5Ou
O1hHv5Y7jHQilbw/TpdmrBwm1zlVVZBZA3VZF4oqjoLCkn4WmIPwIEuRfqexCtaY
0gCRc9iX5hW3dA5ln5udqEr3lH8pm3KQ7L4TaLWu/2vLuHCvmuunIWQjFHQ8BSW6
98TtylBKFYNCkag4Yjmm0Ha3I8bKMEpNaJtQSvzwKfTyXR0F0rVEWnFDzBhNnPzU
7w3dQjklXvMJLuk6C0Ixyc7u8Eo1lz6gQTeCpWxdEKH3/Sjg8Z5aEw4/UV4eYyzD
4YOdgH4R14I167WP3o8guV4HLhUPVPItT7f7ksZcXuBMtXkpjYgdxtTZGoGpC0ae
7wWh8MKh6Nw7A2THe/lN6/+3VH02cWrkzmhUqckKu/F5eCi3lKX4Rn/gUGLpcDQw
0JqR6j/NccaydBSSVu4p05wzgb98tRH29WiVCASUn0yK/qwmHmlI35MBgTyLPTDV
gdyKI4L5odrx0jCOv+oW5JFTFrpw93fx6aILsOKKKOvcGs6V36nOCLSHeTsVyeu8
ZkOH+vPef76pa6YbQlmOdcMyGQuj8GQK0KOH+PwfmwnV4VVCpPzipLMOEvTnZp6L
Bew8mEWgQsv4dbjgHhlLCkxnRmj1eN6arhofWP/LLUdm4ZQ2O1dBH53oMAS6fvri
b56kUhkuItpFOIagyxWuC0xgx/40Ef/8ZGFViyhtt2cuny9lYuerzllVaXbqqz9P
cYH/F5VgoegvmqaZJ7c/AsxAsgHdiX5hpldYs5J+NMXJsVU1x317a9kpDYR5X79b
xo2mF1p5AMgN2mub+7yKF/tkjQCicLxNUjjHXGBkdBMX4YDAL+7yupvutiukvJkB
OKVqC56l7IJE2TlzLYnwbDa/WgzDAqlttqnhYDFEqOBJMBivAcMzwc8mWuTdWOwR
22krVyIUfeF+hzqTip84j41wTU25F/UhUHaPPdgClsu/mT7xfHUrD/9/As2VrpzJ
opeYP3T1Sp7M6WPoFFRP+vYPG1JTvcatF/WsY5zJhAxrg+GZRuhfXhXsYxkANavR
grzIrE3CYlweyA1frJw4o8eLirFt4EqIxglo8pArp/IsIpvQnux5RTFtr2dfCQF2
FXvdRD3P90Ymcs5W+5LToGz12dXaFrHVsFKzDu78LZtvBA2nZe+jEoRUh7zl1KFV
Z70bZAvonUFbz7/DlRGGMzBvu5inIk3OdiyaoMblGgZmDqEpOZv4lLRtVNBf2NLA
yWTCb+7mLsBU2AGaS3aFW8N0d4WxG5RM4gLV3tHp14wvbgeYJXzvMWZO5cwC65If
tRQa0gVpFx/Wp0b/YGo6r/l2H6NwliDPUW3V5cDQAB1lWidD2DseNOyTuZWV9EPr
fZHSr5Q2TeD686VlYPYU1h1ktQYrCPG1ZEIUSBvNpR7X6KDmK0ZjfL2jC0tYqoZl
u8X6RgvNimP+ZcO/+vZ0UfFfPv4gCFQ37LPpXPw1Alq0GDWFEWKlBdaAGFf1c7vE
+WZEjbPaqxxOOOAUg/jAkB9f+1d/k8kVL75MatfE4kfEIOwIaUjGyJkbSpU7BG6A
CFQdB6lsdDrcDs2g2AP2ZukpksEt/GnlAGwDR6G9LUXek0Dlh+Sagle3i1v+LqB+
iSZvUNSd8ybLio/VE8N4rxmDmUNC5TACimGZeztAY7pLE87QynWvbWsGYNOVH7OE
NKrWfWLKEFqr5X+BcxE7+8cdHMIlOeeeokVY/zj5XXyQyxwJCYAIa9HN+638dnw3
W/hSK5aHh21myC6DYsGxyzGuFck87zVIeMkFm4J/tKdbSfckDVo3Qv37JCkpwu1F
jdHAh2MgjxF+PBrXouuKx//bKgVfOyuyRCwCJd9KzGra5tyCO03Nhda2WOguXlGL
c7f6FiUxelJ19UFcbw6372ZhheRtnOjqag+r95BkGmZWY8AbCG5dxGXNSuRNHk8w
Z4BNaJlKJ4I9Lz8ar8BblXwcamGTUI8STO/H5qxOYgYnQM8kRHgmyoxnB0W0yqPr
YglY3UCzQkLHgPKMz2WzEiA7YSuFX5gMDKO/lKpSHATNXMHkU+mqPJcs0g8UFPtY
3uVaDbmw79F1BW5PAxODikdOFHN/EhXhIZcJD2JxIWH0qASRfzf4L3OrzRxdPyqL
m+WnAoUd6XwGU2XRoAKKbM3c2gA7F8FzaqNW9ybLgYXcAZS1+B1mhEPw85dDQsyR
sx4/em14mefxtAAgOvsuhdZV62AERCiBqPOqm7uPj9nrvr9gvt/OuujI33HJZAax
7+if9G+IGaR4e0f2Raj24rZ2H+edmb6hTqc4OdRwFJptwvibXzDITnXxyBZ89fdd
wvih3DhUrU7vGHCw0EqgccLMycPjUiCSauWG3j4REFgaTcaLtN9yaEvPhNjD/28a
wvB3xBzdLj8vRISe46xpbNLXp/wUoopn+U9AWTbcbNRcwA2luf0WYzTkGR/XEZvd
pl/Hleq+YG6vCnf5qQX+VbN5HZFrId0enyDlcFVDYKdv5OZFWKMLuNXhk034jLDt
nuypfiL5J6FlnAQp6P7RQhyDbuwfgqDGkVBNuEat4orGb+bDijJPFokP7IwI/wIH
rpObsnretKQ0+wwGn1BC/3o673Vpq93i0KnnnCso3xbce7W9rr3SomNdFpfj8qDU
UyhhSa+EQesibgbSwsIX9nuCoROvuWLTBXyzsjXHi8AEmGi4eYpRXBJk6qcCgmVI
/WSVEpCivc0EJjdVffwEWJxebEEfaC7XDxGT1cQNjWPqJhYAB1s7nRlfz+dTkUDs
xVpE+Y+IvNdGEeWVngUZ61vTs0TbNZacFjJajUNWFZGNNlRjAU1qAFU+LWa1XnEl
DiaH+UWNb8gxUEWmM9eutnBZmw5zHNrnchk2TtEgUL3uJ+bNywuNsPwwrZXI/oZu
aZ3etPib/aHtAMrnwqiJv1i4KpW5jftDXqSDIYm+sUgfRQQihdUe9U0qSk4IKTln
7S7aMBBC7F0Rsh1LmjPliuRZ1v4+6csRF4oeHJ8HHvUeRWI7nLiHMQOKIvPyggfM
afG2p6OuUj711QJN8C/0XdEH/L0R00nwY3yKJO9WTvoZJEfwLAwTnCjSkm91u4aa
A/z5lELyRo1l2h1//4Wx8vxt/nfSVWeg2zuNOzgxc2cYCU7Ymc51GNF0YHgZMcV7
rJv4SV/4EVZWQ7E/ecq/qAjZO9pi14fqwTek39Mr9lAypvgdUPMV4ksv6zyrdGn6
OWRcQNfELIZ5bKF9Z6LFa8nUiwttLCnqV0QmX12ruqSeBYnA90/xpWAvZKMs0nXk
K+17F1cCtO12X3h/boJkvwyMUyCoeTyWZMAPjP/T4FRmubUWctVMCdUT8r36aka4
zdPBNKKyuUyCtXbXN0liQeNV+OKTkfVfQ1cZ5Ki+6cLsY1eR04zf5mcibD1PsqwO
Kf4NcpP/6hznKXYjp8OneVRkQC0bpdhDDz8UDnCIVd21lNe4+kUn7zOYfJseluhy
x5twOPmTsa/+48/JbjKHVe459d6eGbHuX9EpXVbJ8ywY5qibezoSyVwUN7a8bt1s
33aaSKPh5cek0JvFwjsUtkkiINX1LhUqwS8UunhdJjXDdtdNXhucxeVSN7AQHN2Z
ZZtMdq++/FpHucFx69lDHo8JeqMJ2itXIY8XcK6/xk3SlxXtXb3TDM2Sw5IfFjjZ
A4dyCF7F/czTGQ8Z9VPQDBZR9YOlkI3wApA0b8Dug5BtmJfh2GaGUaqFEXjpssHq
RgaPtjQXfAY4thA8itwXfecRiX2z+kQ30JDa8t7+4Lzed7Si0HH25w1r6Y0hUn/m
ESDj2fszSpfm6a6wK3TVswrGy/b51LoJAXV4soKjYqNqR6/3GVFoT69IJh+Vqi9I
nn3lI/pQNoY2S3dzovnMh0J4kY3mFVRh5tq9WXfjHbl0wFiHCqXXEE/DTRIdjhJN
r6QX27nqoByXa3v7k3DqaJHNLG+vTe9F3IeKgTrtJu1HPEhLvygnfgIZlx4nnk8g
B9fEdKeHdy/0/+lqO0b3EALnSj5gy1mYqbL03OJ0f1cB+OwNwLelR6ft8X3hZbMf
WL3juHGCbbYDdbYZ3I5yvHmeGhhb4ZzZIJLny+HI+hqwJE21JSnHu4ZtOoIGrxXf
0wYrm6OP3UsxwAC0BRoFYUyrtCrg1BiRP+dRCmmNanq/uZmC3oslL9ZcMG27y/Ps
WGFSLOaEKZkVGT24P52yxdq2DVp8FAHznNRi6RIU6RI4YbwZH4F1YROzahnGh5pj
jOIzZlrL7SWCpu6DPeI4l9FEe+yd+J0ZoaL6U6mG5wbv5xFTJ8EFlma2YAwCTVae
5don4EO9RK/I2Npep4R3aRxuazk0buzHjIpSkqmm/+gYL6AIDSMFZZ+A264OC8ys
uHflz2Dml0EGsrMsdfPmfnhJQDTECwqzYn6Dx+PwcfKW1ALw4p878LDMK2UZYdkH
aSXr3nHuE3NN0VY5nPcjH9bM5ufu67z861zoFPVsGDn5wTyLjipBqRgJEbx0VFGC
kBcnew1pypBjDRm/fstOjEYPXgbtwFneDqykbi+8jbXTyu9ZFbPNUUIaywUpA6Gv
xRiLYcnUSMM7jHhXhp1kLdGhSfgTeUyxgdXfjUhOjj0Tkm8SaZJNycV3oU4Ky1RI
DI+08r/Enu3GUKPUkSaco4Nx4Odiz6dDiw09L6WMmcMldK57pz222uaoPuPpX38J
wz78jwbvf0B3h6hhe2my3jIHghD6N4ei5gaeFDUWSDFbpvszHCtR8NAo02pbQzLw
uQ27+9clOupAFWXKdT7v0v0rNhJCEB+InPL4hTryMSJ2xmwimO1QOKkue584mizr
43xBsedZeLhuoPyEqr4pvkoSphHq+geSEuN5QQsC0QdXs7k4cGywXlRKDRsCmIeX
zcNnm/DIMkUWumA2gynElxLkUpcUd1SYE6opvaw0S4UxvHKGooYjVS5BRFTbtGto
3k9Mc1phmPB1Dqm/lYC84M3+ZIRjjm//OkT1wIAE6Iz32lZyRsA9A4e7krWbgXck
ilsOQQoMllz2Q9lRre3LYTEBCpJQKwEK1gPsBvWFoUsTOShWU8QyyvXScHl+lSDR
vF5nMZcOIOg7n/jEatI6VAqLFDRB08JWAipqVOEIa5vUfsL4CE28s+gStuUZsRW9
n6RY91XzBuaJ9aBL6+SFUXdgn2s1UV40Fk+k2gC72R5QohozwxeqICib1yLQerQ+
3nciFKbOjfXsZ4G0c0eVUmQPwTFwvWM2bRQu719PkGZ+KWHGPgEf8trdp4wNeHG9
YM8oCcjlQZdoJhturGtzgkQ8nXHO42IsShl4BjnKOBZ7ncfFhpp8/HIQgPXJ5MmI
uUx7JRrGDdk1Bs8lBC1UzV4gdUJTfABhbcUXpBIpPA4476XYzPEwHOfrqTv1ofig
2iRXFLSB6bLjizz8daUVf4VD9xnL9eZipsE0SlS1KjCaetPE/z/ZGYLsy0Gf0z14
vwSVv+L4E7iRTI30erm8WjoPCXEddlkIYf2PlBwvs90y40bs3QOjOKQcmuisfev4
xhydc8py8t7yAM2+cZ3IQe+eJfUt8PEmtMiXh6ZnRXH+qyTmK2M3+pJhKe7E/+cf
fIW6asqLYHQzRwSvUaUkQSEN0kSDe4wOdD1I821WgeCDFmsfCnabKi3PEHOEHK7V
12s72Ir4hPqfjxMMLFDgeDM978K+UglVnut3KD64NPDQhoESy5oROmBHjjt2cAza
Libe3GSENJcTngopYMk+dtlVQytZZfIdw7UfLsa4orKMrGRj2+yA4vWMU+Xxx8PD
PBaYR95jPfxvdepxj5DistUP1L9ZOW4C0/KG+Q7zGR0/3R5fs47DRhymWgJ2A2C+
TK8HWQi9QcpcfrN+9jhwJmXw79eDCpgt89B4pyEhVHTxaTfjqlFxOgSDpsR7nou8
q1wITZp7S/4OyHEl5W9VCIF4NyA1YQqBZF2coPo2OnxGuXajBS87BKWIblRobWxd
xXRRtO6wL2e8WX5bZEPckDYDUYvrBQvyIHNAEKPKxqDV2GaY1Mv/wvVAw0YEYaQr
WjTvWm/tJA4R5ywHTIgIQaJAY4oKcbihnPATrnGBIf6LO7tI5EG9YcZnukC00Jdb
Aq9YO73pD7dTsW159bDgremi7ZOg1WFjYNT7/M5W/vGIwiHKK7ljyAzmZgkmMN3B
M3h93EbcSBPFA36LOI5BEXz5/HumH0ekC+916pkMs94wI1H9mIMO2DoMzPe8pDMA
5ou9a27fCs98gNtDI3CN/mD1k56dwLoxKbKd82aODqilzS43sfLmeUnfcFvnNs65
+PybOiu1BBzYj0C8ntArmIh1uTgvvhATnfeLXlbJ5SJc2uMH1M3a115gkIqnayV8
KOogxkfcEdBwoDI9UX3bFei+Nsw5Nd++U9VuNGF2CSFypMty1UPpp3Gv6zA/GRop
W2inHRtBFGSSXwBZoYwZaAkARDe0W6psk2eljAemx4FN55cjWwcIcUilHRB0f+Ai
w7VOLJSOeCYziIXeB+XIxkycWWTqO/+maAgjn6PmDu9+A0PgbnwAupo3QGh+7ihA
5Tcpb/U1gizf35n3djYYK78PP38xF/fmyZojjbaRann6yG6WosYRhG/M5/lEIeJ1
RtJ/vzXhXSxDmm9Y0Cq5PsxIrD1ANq4YJ3R4qa/NnM20JyDDFrgmi/3tYamoJo4B
xKfNOoxBuXXz8qT6RtGPTzOh8cGNmBEJMnSenyfECvwOrYf44zkc8lAIOFX5Mw6x
AlQz1ZpMEeeoXs0xhEtP4R7veux3rplPktH0ezGNENkyLanR6Go6ZmHAVHi33iVZ
A0XIMn/K4tGWQRHLGnS2U/V/5pc7FdHtPty2wxIceRKIBK7wdgtdL7Vq2JzRoFFF
5u+aJ2QU3F3N1wJ//QEpkb48UGRAJ0GaFNYHWRLWc/AkQBnTnLNaNzYvDQIRb6kT
ofQQveG02PwxLKdFJSsZJg+NrVyKEJRf1Ttbvan7yRU8aiECUL6UWBRlHNZrFxXC
EaF/ISBIUT0sWHLKHlttmb0lz8K36rrTnSbREUpfM2TLzjbY1hoPY2EfqPCSGTgT
Qyz8g3N6GSmbKgZEzSce7SIqsNW+1DHGFneewHGNF5yeTgEMdC4fU2PC+xLoYK+Z
KFAipZh6nxzvompuoDSsNOt1Bo2QzPGnV6Ep7gYekmjfIfAz62EZ/rY0zevBGBC0
8y13YO5AveDUDMYNmv84O4YdnzqEzu5YO6kiPr+Es5CAwhd99IwPx0BlwUAQVUpV
AALPyihpEfhUS3oNnIOCdOiYqU18LqhrHvOHXo2kC0GMMao3s2/ZCbCVYJuX9cRc
ApUqfE5RQPlSDrfshYlhpOf78KudLoFCSdTBJKEINX1sacqvZapRx64hc310U2Cu
mjpG0T4JNGnWZ7LPScVF82vkE7ogUvqtjDGd2J1lHTI166Y2wZj3yOC92L6oGwTt
T00hhgIscwkfLsKalCWUhqmGNviVXYggLcuidw/6ZZrCF4AvFe69CyvSKCiw3Odl
8ALOmf3iKkMHWEMVf1ZnU6uRYzePPaghwcoH8iOFFNkOojFu5WNXyXRod0WdK0od
04D0m7JUBHnGL4rXHaaY3H1GGsssvCaSMmcOVQgAe+bkpiu8dI7APVyz3OQH/OnQ
4GZe5ScnAPovg8+wg+p7lnYtDtirbFGarRTUY4twQhTBEcUdBreeSum59dk+laTV
0ZyCuLUJwASGmnplrj3vLA3bDuyN9nIOaE4ohh2VBisVmxtyhvY6YHePjFv0xH7F
zqIZiSrEEhckR+VFRWDQFXg6/JkroBXRAG5iG3pbsPWH5UzPAVjijlR9P1816cwn
ivKVr01OpcQ9Xi3Y8Ta+XPDvO/G9OIFa70aQo2NXMLtB8x8XwwWHc8JZgQAqrFxt
97wvXB5ntY2hSUieo9qRCPyBaZq6XsbiMs/7JeWvaYBV4C8L/0yncTqTCvH6L/Q4
+LM6XPiIlSygR65RhiN7XE9q6iM/v9YNu+GNDxTDuvOiBklAuKezyQaUM3XgC0A9
PBxPYn/hs6fZkmiJZWoT5X+E6Kt2sw1YsUBXQiU03S7XjEwMI+1UU6EqVCYV7fzL
UmcaY1NxYY5sWxygOA/m89rhLsV9qrWaNHFbnIRL0PaFKRaL+Z+jORXlD12ou8sx
xEYwNRABWhRpHCZFlFjxILQ3WTPxstvXsj0XdSIqkxrT+TWRNUFDSVBBXGQJa0Op
pclIUKDq9GiEhHC+8nQEmF6imsdoXxyxqcy1jsJFm0BxHQxSog0HOnoxOcSdMWts
o5UTLwHh7PKUcMMSh9Y459afOclRtF5+hokC6R/BQTfRCznJvCwE3Ab5sbzGN2QQ
C5X+3I8abRDEtKV77c9MsdRKySDLVwrSetnXQX6CO+CTjj24EDpFDark5sWis7eq
TOyywokeYFoXczMVT67vNK0ytUwoPdLFM35S36dTDFQ1fsv9w016XiUL265RjFeg
8iC3e1/m9IdoDA0qeeiiC9EmTKab773kCMrl0MK4YEtrDZ4Uu2RrVZ5iYOP1g1Vj
wTdZGb6FrEoyW3NHOwb7QEelrMoRhcesIOLtBS/1U0SWI8S4s90WXvHJp1DrbKeZ
rlPvr237wPT2pE1EGY2GAYGzO5EXiyJo1kGmqZyycFMSYxxxCjR8cZbIV6IEmQbh
r301ML/O7ts/6dPgsoLoJHqmVoHpEViy38VZaz3AIF17gYl0D0s06mWkLVr4/E7z
BUqYGx1ChYFZf6AE2/m2XQADSRGaSGoOhlNNdFWkTkh03mnCs3sy96+UjzRrI4T+
+ReQqVWoL/HrwsKac7Urg8fNL2lENJlOwpVrfTp1M4vABfHFeJRL9D4EGfm0uyEf
kD5v0PsBJxSzrp4qLLi6BhZc0jgn3v5bBcwJIYpMkIRBqBxF0WZ8B33wBvKayCKA
DnsP/YqleMLKK5NjO+VS8tU6ic4AHL9QoM1tkOF//FHeUHQfmKGCCnTeDw2eaH98
jvLKLOLnQvzavER2EsKer6IhvTFh4REn0JDyZWAkvoDFYkb34aM2b/SaLn4j9wXA
HpaiQ7eQSSk3nbj0CPwgE39es5swwSQao6v8p9ewd7rEkhQn0llw6IJyIcazyo30
2oUv/AAx0XHDw+bYLNGN8EtQY7MgpMifCA0DtRUpZi21SdUyZuOyt3TBvfW3rgN8
BPrA1igPNR/ybXVzgZXpYHkOaG09eMTsd4kk3Zt7Nwnw9avXZE4GiYSj9mwepfrb
rPV9vJVmhkSvGHzmYunw6rywZ8+2tnx52CUP/ydBGVihtXtJ+erprN7Or7qZzajB
bi9hvZtQ7/46UpfeVxkPWjrnMsq6GM8GlQDjbT8Xu+rn5VEZFzQ8eZvC2U0jQnG3
HQLfq7HdT/8D+hQQ0YKNwKgul4qr32HIzvBQ0Nc6doQ6JgXqVvrDh2av4q1226IE
/ezD6CU2/kogs1HEABddVmcStPH2ZTBX7SsfrROuEvB8TUCOaXjusjKDlxGHBfer
Igx4lsPcJlRZeUalXUCI4Gq7KrF4ByNvU8zLIXP/uZ6gRHrePKdeFIHtNw2QSDXl
6K8Z128EyqhI3zgPgq5h16hrE3LLztsdICEv23C3dAv4sGVYNrz59mYxmDrzQH6B
XQzIny4lkDm2pBJhNDCyVSjH+4HenfSoIewlmQuUUgr1RxAHkqQoCG1r76e6cjiz
hk/mUvpaxFXP9yjJ9JGjWvyBadsjHpE/I3YPuq3EzDcfeAwZ6qHCH115Sr+F3atk
QwJ8fjF8xzuJkFyhQNJ5pIEv0mPE+osNbqO5dj6UuiLeOY2n+iFXulZmSc7b4of3
gY5U7ao7D9POMo6ruSpiq6fVxP40ly73s8BnoyXhSPGF5q3+WwIpS4ur1HwbZSvV
GrqAgVHYbBGfd0q1NKGIlldRJHMrKlY/WQW5jRdOBWXqf7CnzzpN/QuoapAGn8BX
fC4j3ROiSn+qH4IFSF3ZGA0mEJWkT55SRtbuhyGSmG/vOxMkhGCAQw9yojB5NEE+
0dJ6ZIuDFL/7VdaKp0jQcQ2X+oTY6GK9DfwgTuZOKhDe9hOpOHCm9bX9ei3Z1uK2
E86LVVDm4Ut3m51+rL9v2oEzeDV+XgZ/fU/q8IdSpK2c51YKmxFYrWUqW4KMgDt7
autgJ/KHe9wPhHqVTe/fR2TxoBIRy9qzX1u+EQHqaeX+VtFU+Sp5f8rY5+3VIU50
/Nqx+cypoprAaSVQxUZbpLebw+S5waUlH9GV3vV82MZragF7jr1WLKh27YhU6zxl
HlArJR17+G8RaPd9E8WJdZhUI4/YiZxAQnn4y9KkQaxLNvpsTEqoT5+geOr84f5L
MIe4k+Z35t90gB8Zzx5glekqR/Z/m2S9DA58LhdMcq7YDedffORLa/4RR4DEO3ov
0i3gmpZvhSJPcM+xp7B+kdFPpBl/UWr2RPsyhQ6pTzN6uJAOyd8XjCA+SZVl0XCD
PnRUpqnzQ0iun5NLnfzQgd/lMl3E3MXF3DtYe110zo9irf0wjsjpJ+LOnbQOlaqs
S7hRWYb/+ea2Qa2Q7p0HijQiIsu3wTCDP9R6yGwYV3NjyTVITHvK4YjU7Qtox83v
5dwiotCmFScVwEDIer+wnba3hTrqv2lJevE5PR79CinHoN+Sigdu/Su8guXRnwg/
UIRGrjDfyNzTEbE/XAt2sapk7IqzSGwQS7zFHF7aUt6AmP8Bj6am3N2dBGhkfX/O
909YOCpvcKGMeIacrmuAlN3x1XPvUkbjLhwVlrQb78LiK0mGrR0iJas7tRCqK1vi
iTsodoVFlBgyujlhPn4tzWvu5SlTIWKdIzFZ8dhsMrwtRQcIcOPCIduiikJqbkG+
Jf74Vil9RMWuDYfFXjIDYQm0BGF+Q2v15QOXyuDxx0CSMqgAxZh88XJBislbGLGY
0IP0HGMmUMBvafkL3jj21+SoRZG3muQFUfy3r2YS/gAvRFHwUMMiY1DIlZJHJgnb
O3/hWpMezffk751R2zLcjftQ6xSiuG/WGAUigZNElS1Haw6LhyunoMMnf8EHTOfD
mwXT8L/MXs0O8CLFs7Mza0KRYYcHYgbl4a2bNKOfse6qFwiXhVdkrk6sJruEsSOO
sriaB886+iN1zDx+kBZniOEmnI9WeD0v/jdU7vCJuryv+xr9fyq0BmNU23kRTG+4
iMsfuUFlJzyS4idXQGynH5xP9T3dnhNJgZF685yfY7jxq8wb41RFnIxWFefMgCo2
WvvRG5UiRS+8Nokl3PB96FPazGMtskX+7enlXS4DzktJRoZmFjrPbhuEAbXJFmNV
vPzbuS2SlaWva1HxkFGOLqcmFpYXOeFYUDOD54DGrN67t/V7j36QprUwB2cntbCo
UdYGgRPOyU8ZAc3Ftep4LC3Xo5Cp3gxirLYTZJEKWtTuYnONjZZomVSnixNO/A0d
krpiiIri0mg7TqUNZQTy6rOYoUMy8MwxysejN/Q1CMT3YRroBWALoX+pWlKdYOm/
A2yMoKzXg/DAYurCT3wVD0yTvnLImwbSPlnAafGo1C1yK3U4V1YGBmhpMWF4diPz
cR9NnNT8tGVtpTKIjx/qbS/W2/PAnlhZ8y3z9ok1vjlUs3IYrSGic3YOJa5JtvT8
wy7lk/UgIwvXSM0e6TWMgr+q3ZXFDdM6npv+sHVaMJmSs2j59silGUsRSzOhzSus
KFZrht3QY+jBXN56vv9U6C6iYlusm4TuOqK/Ajm5RmGiWmZLrwi8c0tjgZGtFDww
rCOBWsHvPmFKwBGCOzhqTesBpZJdH6L7LvoKlBT4RgDLV/sATwzQD5RlCPnYgWD9
zQfDJsHgwGEqiuOIeNXQo9F57Ly1XtwkN7F3CbiJKVWqTAG1kM7YnUEzlSm7SsnZ
NRQERjAt4ESZ/OIhiaWOV/R6WSlbz16IQRzBYdJr98V7ps4kSR+adYD26ggochVn
n2N6YYdBtPUPGv1woVWVojgvPV26K+Id4ZGHVasmzwuJ3n78wn7D4MNgA8eCsBcS
u7vI8JAjZXo7tSae6eYSHvUCcvsd9eftSmUhB61ygT1Qh3MW8o4g5zISZSoufUf+
fDaDcgKcm2mwkFkKosn5lgT3M3YbQlxfYhvQKTsi9wYkA7b0jGOP9s4UviPRywPr
1vF/urMoO7NlKEpbjcOxtyBWJqdSf6J/Lkw4HEBNOCJQeyj1FOMsbIVk7rTWgdbQ
w3RBA6fXjVWWn1C5DmJmoxklPVEivyDGE6SVeaUSLppV8AtvayONQZKnuRFcgTRf
Cgv/8X5NMYihCVQL6iSJQUh/OGZxzwZ18uUbJ0KGCTvA3yITio/At8glQmLKGqSW
PaNVAnLcToZCv4MC0Hvua5O7gpy60Bz8CqstFOKDzzG+coi5OhslpXgDh2zl/Ld3
jOj8d/3UEtwdI7Z2h0FpA9IWt7LHYm8wq3yXu2Obid0qcXVBaw90TM80bKP8EF+T
5+kECP2zPsq2RD6KtlieVMjKmUkf3HX9fBQzqhAjHNgOxKCh7a7F2418JWwH07wI
pVgoHpLUP3zLdO+oomFv1rDVW/Q3wOAFtNyYe7lmF+3aJAyb9jresX3ezjPM1VkQ
lyMBuAPKvujz+fjT34p4qMLmuJEPWXBoNzNKs9ETo69KrF6tqtoDTm5GiscLm8/k
OBHWvOQ7gNJG0R0cSp9a0SkA75IXa3lhFJGaXtPjp9hr/EpJXHqlbQA94yrjizIA
8Vfxr+3YLoHPVj6ZUnDHVGjnpjjZSTlr7GbXr5J7LOH4MR3ySEDUKITAFjPO+Wrc
yThMaNndbd7BqjNTZ+Lz1aXtD9nQQ6a6/x+vM2hfzkpxqhzxzioXIqNyrFyhe65n
2X7lCwPRetbgBCEKRdOphCH8gRVOaUvdpDPN33gp+vYRXYIU0HUWVmv3VmLC+hXH
TO7CdccOw+dnkUZwFjy3oL2RwLd62UAX1pQCWaa1IZJXo0VaCD/4JOliONxjNuEZ
ZQOotFtPu9W3E61b+Cqs0Venue+LSCqXoNan1uaYhiKptYSvBg6DgzEm2+MN0tgb
lLACmdftMUJM7/VyBu5TK2jqN4HsL2735XLy09p88WYdrMp8mRC/4JyNiSwh/BUf
2qJNrMgUz/efnuws7CDS8SkZv0K4ZWOmjrbN6ul/XKnuVSuxRNtZ85gUE1GCmmI9
0806Nl7X+4GuqO+PYp97X08PtboYlBJL45+kn/uJ06bdDlkDM5j8vhcaj2sDxw1E
dktqOm3xrpaHRqDD0v99Akiu8pNTF6ktX31WjTx199aHwiF/u1CZhig4Mvc451II
KXOkBeYTIOGBx9Lk8LsxGGf/b45dPm4WFGmpVgSL+uyZ1UuLfQbqQ4ZMnlJHnURt
1w8hRwfNhrqWXXpH+cXXdDXXvwWlqZ9ZMS7h7C5ygnLqOvrqeo/HPuzjO3/vW4LV
RRQGlGG7f1qXJCoJrDio8vVwHXiccHoYHvFDPKT42h+L45O8lCCVci03+m7bq+4a
HXayeoxRHjAIxj7tc+S0leugWt7XWff1bxqNwVyHnE3CM6MKBhAsFZnBE9eolq06
xAiXB247zTm3aUWV05DDjALO+bdNhI8AVl6c6z6Br0mrH6y6J4IvThMEPONG7I0d
+T4E1990cbDHlj43z/2qv94KaejKCw5r0qDe3jqsofLtqeGD9clsXtUZB8OQdlrA
t964geBO/BtE76WR8XwWBPuHmqNRa4jwZskoWd6tfU7gOPtJwt+7kF4QBQK+ZEQ/
1zK26QZgxDs0987L44kHLT4GIIgtV1aZw6l7+Htvabe9mfEcisFL385gwJU2xS0d
EBrwjX7ZO/G31NkJCXCP62Qckbnrg2CJb8x9hWXvoUoufuCYUgpA0IqhvWztbVYU
m89qEa8MWdAUxllhnuQbsY/6cYp0xHG2lZdKVAZSyWqp6K62QYCoA1PxQxfIG9wx
niSGhmsXLRLfwkj7iupqGmbv4/uz1orovGJBS9+NwOC6jWJRbP7SDbTXJaGSCziU
v8whMuv1mGtKqfhyYvOcO0BbhE3W6DkunTlXYvt1q91nFfGBhoD++fmlsCfywl99
ksVLdqmtA0XyhvezebviHHmwoHZjtmMtkS4I38+0qIrcohik3h6hVDVFWeUSZnoF
7GDL0V2ZwGmnFq+wsLpdnQKwuqlS8uUV8HL/0dFEzywg8dapXetyC+5ZsaEzetHT
bHp1BNWVgGt7lcvEC401lKpimkJHN8Q7Rda3SJSLD12Zfc+LzEsPlCy6f++WTbNJ
uwckS08dhfAebe3o/6JWLGVRK7M9+fzC92q6acPhMEGidWIV1uj/4zpn+tUEu5oN
Q/GUKwDRjkJnwjRZgzMPEd7AAevAPrBhFZw4mwcc5UA1XlSoVVCvMj0+dTy6JxkZ
EQTnoXvpyWPSkpCCQvk3P+0XaA+oDwBKeBhUaeiAbSqf2AxnLyzgbkkhj1kMMoXD
5LEflEsFFJ8VHj2arHWoFpDBjMZjo2v61J0dmKAOSDHlGTgnj1KyroGMiNchZlVh
Q2ahPDbvSPMeiPbUhBjYVB18T2+J/h0AHOPQWIeulZTqusGfFh3XIOH/P5UwOHNw
8n8CukSKuPU/ruwPg2sMewAey6FoXg+AkxqDamu/H1rhcOIQP2Z7K5btkJhWZfgV
93hnVScz9QMl5lI1r8X3kIxHDZzg4IapFDli87l1YxysU8lEhZ1ANE6GL25PVFpK
7Lij1dmLjIXsB7LFGii0BHHK5nTOdi24d0qRhKsDVILK1TIzkEaXyQgA4zLjMIFT
yeCQSgBIqX6As60wAVx7n7J0ICKx1bKFUZ1oWvNy5eGz55uHSLjqRrKAjM//P4Bx
e1PMUP1FFCq1flxO+C10HYZKDbjggmztSU2DvV8zi8HUGliXyoPfSQuX8+iWGK1h
tDxd5BEKSVec/jODrEEWphBiBOGSQ+LVDRuRtP/978a3vD51qqNzfGtsHO0xB9ID
8Mc2AsaUoPNJC00Q6ZhupmXP5tqVv7krNzSiN3TOFqalL779U9+RrCZ/q6cbKwfD
3B13kau9hYY5SkbB9gJD7grxLrwsFdrZ/xMOCmC0CBB4Ddm4maoNgPdQIwdZFDp8
UDyzKxM3aO14x1pSiaiGVkJ8ILp9zqD2Th1UDOyZESesNVrF4nUECNwMZX49RLY9
JJlSbzmAaI5+Vx4/7KV5BmJJwz7/sx6ZX8okm14UF6RTd4rwcz6wdEAMRSJj8I5E
HVzLd5oJrVHVXcWLWKnu6jIBIto1gBlhTzEQp500IJEr1fXJV0aqVsRQIG/tqZy1
BEcdPOxSM2bd2Wb7cd0jnxq7Iqs90ME0IdBO+826rxmC+yHq5x/OsKAooM/z+6g8
C4rE2KCp+MIwRne/sFHaI6VJrN+i48Rh57FDJkdU2A734CeYJ024K98SVyuAEY1C
ItQ+vbpUZ/rubHeDMJ18CH474OVCDgnMUQF3L47e3dh/MQ5do1AP0Y47JPrOyepy
bQ/uZRtwQgJICREhSujM3TfAnVwW41oLT34iGUtJaJvsjoY/Ki1IKdXBK0E0UzG/
AXCA2G52H/Oa44Tc88gVuEmtc4TDM44v3f1QBjj9XXXCbqLhGZ8+c+NgxntR/Y7F
ZVK9muEPRNVWYzwm+a1uDSH+7ofFGlkAMyqcXgst48G7ihBSa0czoW3JC/XyfPyU
nVWPoj507SvtoBwvfqJhm8pbHnZhUEShoL9hx9Cm1XPQz9OrgedE3F4J+2nReqo9
dXm3St+ZOp3gljl/S+PWaCwsjDJCDh5yO6upTIuo8VwIxrDTn3xCzqkC9wFm4yWV
2mAaZi8GGn34hc6QNQg98IKuG1oCDIVTiCFpYeUcGdAiB7Ic8lEglCbaBUIWRvBl
ytZ289vYaj8QAZLSMWZTMiCvenn1JtskONAA8TbrLtiz9bu2Xfr0RdhIdwdCOnxX
tkIolu63wFf1ukFYLDxaaf1gEgW1zfh617hAFaScSsSgWU5pHR5HeQr5r2ZYQEoK
yXN2cu2L2fZTBOtfSpxOunQdLcT5oFhhs/mVtwtBad4xfYvV9Q26CRVQCYJlBuja
r5mIA0zySAsi83S0M2KcCfWlKhIlIQD8rLqBBdu3cuQGpJMZqoUvlpJ5AuLD9YHX
r9MzuvcvuRflyGplt9TmwQ/rceo2p5B4Oe2tOt5XRGNbMv6Hg6aV61B9OjDyDyuU
6zhqkYdjS+2TYPBRZXoLFEWKXduOp8cMX06iFPMxDgM5rvXBUJgvGo4QV2wqPtOy
NFGzTZUnLEUo3hReBKoGYdMjfy3ZKWRzhJC1wYm0FVCzyAIHHOSKO1UajZ0QKM3s
U5+f5w5F1Jn30gxW+nU4lSDvYwo+Ai7NmA3t0cVi4xPwSqf0pFJmX74z4rGZO6qb
o8yKNHakKhYIGcQPipUi2A+GDGyXinFm2Z1rmMuLas4wgA7DlRtQR/DQbBCCMVVA
oqngIxLW9IN6A1HLn2PO00JX3v2UHsN5mEU9isL+5ICDIOFonV+U0tIB7sjB2+mc
zym/6omY/f6ka3SjUWc80tIJEJwTKEDwIpxW4+Kiss3bWC5o9s+BWhDHcxdFLLBo
nmUtMkjcjv6bY/HBA8ILchNzAocBTr9tbLcf8rWfvQ5oidDcjUGb2QZfFuKCV8Hs
VkJqcsOKbFi5IzEAFxd4hTmcFLM7JT59HMRegzXLgU7rQaIqarERkENhP3f/3Jiy
ux91HGfTYKR7bK6AuOS4JmMpMgk2LmfPyUCHL1y6PihR3upAJPBOqkcnJjt05rBi
uA0qAB/Oh58y0awLL/uMAlXMzOpMDWfmN2n979tp3l1KwsJoV0j4+dafHtY/Weq2
gyhdX3mCUgUCAE76B9UIP2N7Bgfgxqnmk1JKGTxbbnVRpYCiMqDPBxPOt2wfPCEW
j90OVxel8Amh0cZ0L5TzP/DG/kmwMtqAF9758ZXSqJSL76uAUr2ejhUg4yL9C9sk
j1w9pDbWLZQHnvVX7gwuauiHzP54J7iC8/ZqRU6Io5rAqNWwSnAjMQ7JCilykuz6
ETO9eVratRxfyqGmSBW+7mvf3yWAL/eWUmj1JFszwicz9PWu6i8OMTp8Mb0d/lfr
0lh05a8tA95S1iV94FiglAOAviITZiionN6uJ+1qlx6JOPMTj+c7NKWxrqUOjegE
zrWGBwXxSlSRqB78leVtzrg6RDE7r0BW6vj6TXaKaB91o7GBhOiMAXWvSQM8/XDS
4OxagBjByUoMUoX+tykCPpeUNsQo6rXAGp30MvKVZwVizeLM36onkrmDe6bO/o75
cZsudE848K+qQCDQEaUWzMGxVng0euz7ZeXRw54xR5alX2hEZAxxLe4CffvtPlxO
T5DRcrtmPRxXmUJ3RFloBqKvmvwOelwNG7oMZkEX8CUoF/HeN0pTJwZhLYzBGG+g
+YED2mHilUj0iWE7ds+dgoOmHuAUUC2Xn072AAzk8iq5t/vghD+QDGoV+Ox/32r1
cI83Yaykb/fjcwpdh2Ka+e4YV2tdcDbgkb0ktNgkC+OwTaLj6t1zIVlOPWvNefNn
hyij7/l3+DmtL4savEDb5YkOXnrM/+45AXRPbH9kNwUV7nnWl0XA3+gJjTYv9MBB
oFovNpBYJbabQbUim5lCQUemDT1Brm7FCUCthfdIt6wqylQ47rUFV6j5X5jbNaYo
KWSgF2PWQO8/blOx6ybnq2+76aklawZ8Nxe9TsODKb8OVOOLF5Cz2nn9D4pdKuDB
k0K9Se3pbWYTamB0hXKCNpWERLl459J3Fn4wATU8U7LKMOb2MS1PvSeydZIdHe0X
VuxqWCNN7g6ZGsNsEjgPLBsUxtf1DLX0cJOkZDipNqTM0BWe6MCg/Io8ic+q8iyo
OtziNOXth4Su3hn6oTyupDF/ycLJ39fD0K2xaVj5JGsh8y7V5md2uzkQ8t0lSsYe
ejrzA4F9ZyW3Y62WQYaefTh4EwKYhAKRXgduGa4pSuOLoHdmDwBnGnCLsk7vrCKl
SDNYH8kD7MtfLa+adkn08+rLz+LE+aRjRUlSueQC43Sip+trj9d2vJ+pKpsKKTIU
6nYm9jM9Jv+CKGd9COHYZ8bezA1vLdYEcLTEK2qRduLJMqkuzXuJgZA+1AZnUUAi
Pgpmh0SwzxuyBornh3C+tOnH+42WCGI6465ld4ASCFPh1gaHiwCL6U3CasKiipCy
OHhHpNQ1qiWl4w0Wu65DpDywxmkjZkDCvc155tB6BkbvoNzagOHfak5PXVGEWtI+
UUmwOwtXgQCiJGjfhYU6Um6uvXOUtRCGF3SK52OBUGqDCof3gKM8wLOiGrG8FXeS
rw9DqTfTAXUkoZJifu+jqM+OrEkAGZcJamxe5FUvUc6yoJehdmlp2Q8JoXQu4uOi
JqlT/Lzh4h5B7mMPzLCET5EU5o8AwsSKMUWlm3cU7FnunhVyT+0+2xmDUCaeDPKH
V3e4ehkYeQspOWL93rIbnE6ZvgVnDPViegZ8Or1d0Ue7fz57lKFZjL553fEdVZOB
j59h2dThAVba2hp0m/PDJzMDSl1AaGCgbNlyBqG3i96vwkZ7kffbKhyCb8Nfcrz8
iUPuFkWe70wNl9bDpw+bDR/xHv1nUJlUk5em6pReH1VVT2btTA6YXqI+dv21M/Rj
cov08itwTSm3crfeAv+sVqalBzCGhZVcr+aypW09EGysTk2rrw2o17f5ExXLlFAW
cdCM70Eeo4x5cWUUwbRdgXCB0RT5lNRwHU+Wub+Nr06XNuMK5edQykvjb5xC2d19
wme6zZLBH4IKdx9x9EoSfBHi2s03Z0v4lGv22HCKegfiiSNOlf4k2ADfr6s8ttMH
rqIUi+tb2TYGI/t1YEsUz5DzPtpneUw1zzNufhU2nqbY+AH+U/61tw8r3SQSEOGS
GgXFgYfp4zdpfOyRmbG1MIbhuFQXzFS2xDxErLYw5b2ieI6iJeIaAYIULTTWCCVD
/LQNf5pOL/EOScfY8vppxBIt4DW4uvMzkSCU6dlOqsD+ukoqJr0GCqSkNoyQJNC3
H4ayu2h1Ap+ViOdz6pw0K2bv3VFaS4SNIkl0U/JAIoajThiW5HoNla4rD0O21iCh
Ft2k2iRceEIRNTaatqmxUSJp5mt/W+aZcIUteL1RpzwmQGg2dW0jEFB0ZlGpiwYc
b6PG0FW7b29hqTeDxT8A/BqVmFd5LdBUjvlC1hXCWKwGhiSLjycggXJiGv9jQnMV
U9icKRVrGwztEKkx5Tyr6bX7RqX+QPS4504mZStM7uUcy26RWmvs3gAs2JVC8JAh
oE1X0dJ4DXtRADBBCmbtD2MgzycL+BHtT5caFyJpzU+oqEMI9PrSUpIWxhkWYrQK
zflGsI97yuXrU27HGtLd0yIsambQKYiRbKit8c8jgkOAfkwgS/HCtJMoiogwKK/7
KGh2Sbh/Z3o5H14s2PoTzbwgJYMFgGZrBQeuvtmix8zSE1D5iscTG0Y16IdRTQIp
2AAE9iAQOLAPF8jQRsUKnc2iet5c8SlV9oEvSeNHN/FeJjzCHWRyUwE27JSE6Q0e
rlOuFxHK0YCHqIqrkqEBAaDAciO+KwvhG4SGYujykfJhKs4tRHCNxIImDLymPK+x
V5dAaAsqM84pv0m5tuGwLTrfdhHEDUdOueDhDr0pGUO3O5WM3Kq0qxZVvWnTA2KF
AN69zE+2T/bZTTLJsyLgTUPbiyTwV9Pamqj5QHS4O0+yYJzKY2MTq7yY8vFcHEt4
B7RTe7IG0Re4MIef9zkrgq6+0ieKsj5bhtWXyd76EwknieHJvETjmH/TuDCyTX/4
qOn1zE8OPllGWee7lwKaBLXNULGecRzOgQq6ZRP29y8PjRBNN7e7EniLM+Vsbikr
w1g2dKdDckMko9LBI34bTWgbV5/O59URIpxRHvYWf0NbBr13AsB0AlwJDm4QYY1d
bctmYTgdM36BtP9jfUsa7IlQMBf7yuwPyE7eKqo9KGWpGyr8pP8pq7X6E0XgYsj4
dYUrq52cU8wP0GPBFLElsgVtB71KOnH6yQkL7X3EPDfn7UsdSPLjisajml/grEra
FXzwfFb/gS3Q5BcICgyWe9211fDo5LPQOnq24xridu0esN5sBCFdwwBaJVCq+jCB
6pfDRglWW7smra2GBHizIlDqbfDVpPtz9UceNqMuBA6+W8XfpxfC5AzzhX/V24Io
7jW+h7E1Yn/NVny+kWlhLzrCY6CMXKB/VAVGDkbvUSn0MGEUZ1OmgOkNtp5njtAs
u9UwBBac5d8HHxZP36/5JBPcliF9pgXN41Z7w5xyjB2G8wE5xuREMWPd147I0nEI
9qJvgDDYI1cQuOktdM/8XQ8V79bHtv6twUjrLy8ornfRT/HM9Qe4OgQC766zk/JI
49kOcnRqSjpvWuT38S8cQDZ4VkUKXJdn8AbvmN7NiBwq7INWN0vYfEdry4Gmo58Y
D9YesucCq2IIL1c8clHUIO3zaEvDrSBFd7AGYp+FaX6W47wu91xunt5cNE+7D0DN
PsNYz9ppJkXE/3CnTYIGY9wsefhZqFWIJEv4+gTx9cF+gCEXDoR81ibSLEFttl+j
26pGiDO+J0IljJh1z+L4R3A3K3NUaDMUwaEIo9ngzIj4AyMNp8sbeT+rwQX+vWRX
reyKRX5scmBf5cBGF5a23FyLQ+iGr/18kZO6rbJOBuLCvOQJGtGaWszOi0X4Tto0
CcLIQ0e/9SgcZVFkK6h9weEfDDuFovDk0S2ekw5Fwswtfneju+NgudvUWYNBS1MU
mlXWeFQGmhBsMiT6jqa331qIKW8oeLgvHEEm8lFRHion3qEkROvEfDzRH1g2uJ7F
HnRUq6fEo6nFoROT0ymnDIGgfUTbGHP+3DvXyCb7dcYF9+CvoFTP3RYAxb0TMHq/
yyWnL/qqAe282DfU2XCwAPBOvdZSgSdkOY7VAmc/rRBBYok666tIsmSWQkrtuWFY
tumqBiwCeyrs29Uj/9tJftLqJkrhic9m5bTF/i2XNdry1rOVAfIQnbdeDPSbV/eV
RBIEcjxKvMVQC7i537LgeddZ5K+vb8Y1yqTUGUAQeMldubMuvRAfM30G8qpgU+Pp
V/uO3j3ayyR8KS23rVHzEF/3K7uqStmOjLUn8e4+zMe/SLo0ehvYhiT7+tNf6y59
4zMcuBeaECKex9iHCgX4EKLHyz+iSqrwfYNbAohlivZKXXitaCprEwD85jgD+k9W
FWDEQJSDDcFfTCfQkNdiVr8E2tDTxrIdxo0zw237WzSW311JLOZ1BSdnl3JRRp9k
FkN/o80JWAUAOHpAMQztI4yPqalp8lqurDGC1fUruExz/ZcOtWkgEPRjuoNvc8KP
q0KbPXz8TvRpilbX2PL7Jm3plwF8eq20aeOP/I5RYN497jBemaXVCa7qQSvJvjYp
mExxZxEIXG0n3Z2tm0ShSqh8dXjqNvD6mymZTCfMuK9BwhnnndG7yGhsxnTYnFnR
YQgt4682daqab9EqJ2NdOvDyIRv/s9INQZjB58FUsfUbhi4mAeoVzrE1thqMQfQH
LMlPnw0XLLOSARSZFUso1h9sov40PmGzWrwPwLBpzls3B/myqfi7AdBbUmNwXIOa
0rvBkea3+xZu2qm+WybdTvYBakYe718DwmRPseWVEi6Nsg8/n2UvuqZf+C1oBFdn
fi4j2N59ApLIn9g7TBhq1uSyNDXzNMep9y65HfrvD1SlxNx8Rsd/1/WpXyxLIrO/
6zommtKurBN5ak78VYy4JvALamtldLFOf+LmPpfDUHG57ADLuWYmHgl/eMwHkpom
Rhh5Lvf3KW/9C+BokW2DC5Vbn3vt79XVuu2T3NAp64h6IYWT4HpbzY/BhxMnhwf+
CripwIuW7VNn4CFwugJ7uOkp9Qtp4pJzBXHOmQGktz0zqFiXV6Kbi8hBL0CdcOW5
XppkMDnrg9WqBDrOBIG+pKVkWigQLt9UTpL61n8fegY9lo94XFKNB5ufrMhjkTKA
bpjmuHUtVikxgeUNsBo59jDpdHuFFUPXTswnanRnM8ykeSr0barsax1I8jHFM9I2
9AW1PVsWAG1LANu0oHadiMBYEa4D5AUIcesbky7RY3hmLCRnKL7C+HyCEBwC2WYD
h8Ak2+PcqZBhgQxrhygrVDgdjgE4E2683X+9GxjXD5j3HPy2ONFP4MM3fIBlvkOR
kS7leSsMBuN7nFhEM0kq4FhG9Jk1M/1AF6gbGkPP/aPxv9ft6R0heECtgWI70InL
x9nvGHaBz6CGQOj0DSjq+/wOdJMsNt35Es++TuuiP6zALZn9+ZZ1HJLfF/5fqJsl
QcbTK40fkmkAX1CJWn3TXb+GoejNBHCeyjLhH9NSIz7jfff7w91sM/gB+RXAcpjP
3Q4hP67TRg5Iewk5Pw6I7ybsqAFd4jZVuduZlKgWLSrnTrzwV/4p6d7aGtq9qP54
xrDBkzEotCfOy35fGdO1n+W0uweFH4tzsQHJLy/Iuxf/h8fsh30zYN35jAQYA/Kl
7dJ5ZxzraMPtzrU7oh23r95BIQJllv4ky0TcTPedxXMFLrD5ZGJBETy0kjC3OhSQ
u11Kwml8hO1g512pHG9M0OmIkiI77pje3TUBsXn7A9U5PwVfgzyeh19y9TWir6/m
YUqJqSlnqNxJS9uCPajf+K65Dt6NYFrf14wpgKZ/F5UxdSJJZjVoraFpW1dd+KlT
SYcJNwJDYsmGBBybahqcV2kVKAiyZlB2PaPdhdKK14YSxyHHtnpmpxU1P9CGpXxe
sIKdaoXz2V7xlhdn9NlTPsuB7GgaKA1mMCnS+s24YvzrzRumsybKdaMfipZnuAkJ
izpOmDcML1C0UW3+DCnNYvKRE1f+sJ/IcmENhNiUqOwSe6NpxkmIGRA/5kwU33cC
5nDX63Fnx7tSh7t4O2WCFsEWpah2djPq+mIVcyz2F9DJ6Yr801RORzgpnx3KIM+A
8dAcouqHMh0WZt7lJLym4BiIgV+a9UYPG4S85revBjcTx12A4C+OIVTjk8ZZvOhs
2b8urlZ8v9htwvf4MKPd3Rt0xjHi3G16RFPZNIpniUEV5W4bEG1uTPfZzpCcaQbh
zHKPMWMiI/WT5gEsAT++beN9vzAhhTomZjR410DfSQ4HNxO6kzJKgY5if9ssyY1l
tKmH/VzhxM1s6Ag/1DwG/DsjU9hhjBH7WK+tMYCAflypSd7NRXpGyPmO6xYgWEUj
fMOoOkG2KdKPRyGbHvX+lx43Y166RTiACj16QQs1Cf16cOFxLV3MIb4qOET6Hbk/
D+Cx1WdcUDgtyU/ng/8FZlGLgub2bVRC5AB2N5O37pw0n3FkZrKeY71hQ3sGrAN6
NwKnHCzqruK0HytmlpSq9ZZzAbnBFGS2ZkX+PJeXLrHJ6wXgA8FioZrYE9OhpFNn
l/P2xx+ITXVcYaBRM3Pi52apK3sA+/SHOA1Shq8vdciPtGCMUpD4sy7PZOZma0f9
Zkv9f6tw0x8sFfbUvlc0NXgt0UfZtjenzTj+6Bc5bG2huKlyey58Oh5z1wmzS8vh
0PGmFIlcvjrS7q7q7adscIPSZlIQmsJgwMm0dXEnM2yq2Fo28qS7Zok9lWhjevZ5
ClVjVcTPOD0AcT2n+3AFfO0r77GCBWqCOnlzb9cHRrqO8k+6zYzzppPgUuTGp/4I
3fbO7Kw02SUHxcird1g/uqh+TqLXMvQ6c2dK4UQyDeCCqoHj+wpymvLRNEcLugaX
/fuIR1Ja8TU2T5b8IqcvNmD5Cm1B1AmPZYJo3VTPXLbHPtg9us6MuMAndLRPkylj
4MFwIEsG0tiqPO6dAaEsbgLLAj1c/Ry0zGZvJo9InUShc+qgd2d1Dd7dph0L6UTI
IbHI4zx8vOUBSsUS1P5Fvabsp841JlQVkkpEn/fVA7zemGFGX9Z1acNaRAL+CtBr
lXJConEHR/SUerVZqVviC7F6gFIC8Naez2gNRHD27vPXwsKZTLLpOmTIUpTUYOKF
qyBAXOZjaXcfn49oTTHQeadLloofnCjkg4LKZ0OpFl1BRZMuLp1FNRM4QXRQDwJF
Krv9T6jnbf8mrlcAZJlSgjXEWrdJ+WQVsuTldvJ0VsQTbDRi5ygEtN1hU3NInVqQ
WJyKShq2MPqqaqDvL/Lf1mD9AwWJx5L+/U+rVC2cLQ8DIUKUlDlODoLWqQkt2i5m
BOVaZjqBHZhGYLn7TAX/JDMKEJuyP32hTRmVOsU+qSD/TIn7sSptkmk461WfLjN2
EGDyJqkJrUjrA0ExXyxn9tdQWujtMYYh4oC4P5jHqk10TVHz3DQx9KFwUNvMRyR5
0iUfJyuMWoaB2Bz03Wx0qSmR966wMubt8bpVgaAT8GpxGPinXsNFP9ZsfFH+Y3ok
Y5ZwFK8/OGIwqpiOSnM7IWJiqYE1R54zMOXoa82Hbt0PUYUqFChM2iW2jLc552X8
qHs3j0QlL2xgzlAbw5+22AgbbK8/gSDkhDQlF6XKhKejdEQeTYmlbW616eqI/FcS
OzoRomWDkhs8RWcEhd17t3WqRYd5SMoZa30njqsEqNicrmsWh7cyp/u+qk1kaH7u
9C2k8b5A7bT5bLDLgrfmo/i6rxSdjX2CCjPpb7dFz+0hwyVrGjOIgde0Ysqcz/ug
pq9zlxEc5tIQZAj9XuBTLnCD0jpxu1bCpgIQyM3wQ/II2muIWTd8cPQ4sLKP6Xiu
yNsE4szoiN2XX/U/A7tgEbUwxGH+0GAmbPzQ9cDkQFh0ds4ct5luf8Fc8+i1mAWp
OypA8oF5hwmQusrzRMcFG2dPCFggH4mDNM74FQ7wC4ouFsIxC/Td130xETcYghui
tuTxwqYfNxkPduoM/j+GYyvUrskIBgJEsxrFitsDADRbHS95fMCNNjZltHNO2He9
LvV9MdZACsKf0AxCDY3CSbfmngqfnhvPuhY7pDazEByUDOnTsQy5nDX1SYnqQesI
8NdoOVdeu/2bt1Z0CUZPAd4mRu4eX9c70GEcpd3j7I+HLgaTnXTVjF2HkFT92nie
8rCurLWovp3T6sAjgm9/wO/bkWZsqRAd+4dV4ZvGLX7S+l4VMy76Zmfc6CRATbyR
j3YrzWhULX1KYJhx4zSlOd2yQXFyfu8xEArXCvLy5YhNcdTq8gKhRwssAamDU30V
B2BGyvO9hQqcUahkC4emg63toJJ9z/Cw9KBKU+xYzj+hYmJy7jN3idKY0TlOGE8x
wnc8AMCUn21MLOfWqjoy4CtcU2g5k9ZMIx6N+1xDqSNDIs4OBAtbWwFJxzKOujOU
mCT08c7+jDecTtb9JN7m/nf99tNq2evqVSMCgmfz1lSf0nD1cHuMD4URxexRbrgm
3tvFt68qo2qeWG5g7Fk7JACMuNSpnYuPXmiWF+/MIYCtkAIMNqlDu9vBNgoXvYNd
3MQ6AJ2JDdJt8frrE4mpF2f8j8hBEnSNIb17pvpBTX8q8DIwQ4/Et/8Myo1kosgN
YtdQV5vz7e+MFkTnmYcSdVV9C5UsQl96hwtKMPyhuNC4MbOC2WO2XnCMAnb3KubY
TGu17T9RlSn+ERJReXYjwoqLi/6XVHKM05I+rNuoRmYnVUSJsRXmeHmeGW6NnKA5
mHTfEa2gnPwTCsI52mkoc/imGxn3mHv1bJsubyoAuP1Arqe1BmuUGVqMryGlo4gI
qtj7b9uwhku5JxPOcXBqMs0P6/SsYE/C+7uiqJ/VJY+EvUQrPmlbzvTL6HCocxPt
fsgPOF6IH/KuJG09qkZXopi3SFGN+6Ebw8zkhEW4//g6Q8IJSEPgqQCwUsRk4rhF
19V2JMzeAJs09TVrWpzRWgBza18D2wfLptJrkU/G1Q297Em3zfwY1VxRms/8OkV4
m3iG7ktzZNaGFSvYnHx8vH93pl7mvUm3JcFBJNz6vZA2/eH8aBHN8ffMfy4QZZSR
2UcSBW9UjTtaFDHrDztUKoTw90n8syhPWUPrDTQtwWijTBNIZRDBNnoIODTp8svG
kgkCjJDTGkSvet0Bmf4xq9ghossCb6Ci2iu4GhauJHD7PyjOsjD8SA38uLaNZVvG
LkjdMZzTJvYsOpD6gE8783OTzp2iyl1gNL5p4e6uOwtGgiP9kSfs3JRPJm/3qxQy
L7MpwOsMRqNnWqg7xTNv1qPy7RbdhhkOdIBRY1GjnHbL0bHvcdOhdkLsde+8d5L6
qmuQ/rJ9i+scw4lEI6bMw1DM9SPiOME+gnW3geS5wM9aRSSHZGOJxtJtfORGfDN+
79N5x8aOkBETwNRx/lrZf9zOus+PAGb6zc+4X3O/ez08FMHyUpr6tAj6DtDMDSsO
1cc+3wbRSr95bmaR8V60ls1a10t88gdEZsYke0tAQgBPl4gKjNUr5qY+L3icSO1Q
vXgx2CKlGHlUK8JKkypAtXCyBXhGbmMSrnnVfrfAmSGHwrPc0/xYqo0aZs8daXKr
OxBazpEkFUcR2GrBLUxu/7zFAOYpW4iNOkd8dGMXoiAJZe5tmC+YFsxcsk2LvEMp
MMLMt4Uj8KpNPGv6z/dKZXp7nqncn5gdcONsYd+B2qGfsaFej8jmiHDT/GIw+4u+
4YhyxYMpJgLSZgBUKUqaY5U9ReAnoiQ3mEbdaW6vkuEno+LHHjOXI3aolCvbJsIY
rHyojb+XdDe32yoBb5stlj0uEDqZqAuCO8Wezt9UwWt5adPgu1srEHs82SFB/EoQ
XA3Kjcdb3AhbvKpH5R2UY7tWFcVD24Wy/A640OG1eycukM+4KWlp1+78+6vJcsD5
7K886IbIbL+ZECLaetpuw0RtErSmq03BEaXV9cRGqEcH15cgP3ECoM1NjAN7LOmc
ox8+tNq3tcZpL/kqj8JjsVnn+LWn9e20mJEWph76c5EYdeTlXt4hV/aConIcIGbo
nIcUMDsndAi6tFE5iDfYzmwhQZL8fsHtWrKVhM5XiGzXOBFoU69/pXe/wt+oPuWA
wChqhUr7HUk3S52ldqsX62aySN0o7YWPcwKdpGLmHMIR+qUomvOiDBXhBPjONDwz
dx/7gqbAnDBnKLeqNzrAbbFoLukvmVfcOK+J5MJrXruST5IqJ+Rj9ijeJzaEiw93
Y3fUpMfxMZiq5YITpZOi4xD5otV0uHRFNK86EROi5UDf3PpuEfvhxqv3ZnOZ5Td2
Rj5pxO0ML0/WhdC+VihD7Cfr73jN4++52cLLfO1UBaBQ0EyJ9ZenzS+RInxV0LP6
jwvpwrLVS0qS+OYtGCcHbb0ah6ny8MPpRAg/gHL6+fgT+EppjnfdZjHWNqOTf5OR
yBrMvdT+qAPOGBGT/sHEagVHtKUGWhd9Qk4u/Vt2HcKzkXV0GFP1GNTM0+LlLtS4
0jGeT02lha6J9n4vSd0nBDH12cfi+EOwVs3A++jn37yilcIhpoOn79y4KRuawrGT
BFr5bIkRGaT/KsYyRdQtJg5U4/heOgojzU42NwPQeuhRMwV2KX4EXfafW7SW04+L
8b4UCiQgpNkKsYlyf3TYbwx08Y+oF3dVlPSSIhjeKntapqupvVcLHJAXT72vypRm
NqsOk26W2HxyprqlnKFGdrgVfvex6WpqpZk8hKp85XwFriDIGkzdw17A5PnziUDR
WnbvKotEau7/H50FuwRrczh4ebFjDimsWOoElSgPofnTOSRL9lMOG8YMH/Pily9g
MV1m5fFZZv8XXgL6+EXT2FxvlBqP/deP+JjjVwJU7dQdgOyohj1e0oxBikreC0m2
vtdQ2bZU2t1OokZX79foqW7KK5LYnueTSpspMVZX8/znElQAxgiHRQhUhKO+rR12
lmJJysgSpjVlPpqCjM2l2hxilD3hUgPUr5yzdYMV3N9fyhgwQ8Ygev1MeOftbmBt
MHlh13+R/TrRidrGKVnxD72Ad3jRQEHR6TWwL33/6SSHr52wkFElVaHBc605QMrq
VXtdWvtG/L0Y22DorplWejgjitcgbpHvc7Qiz0Cl9KYx2Rgqx81dzmK6wfBn29mo
BzCVhsKjsGf5cY4IjuBIMR4OxBDz6SD5zynHRNip1xptvV3IJkWAZM+FrYVlDG3J
lSBLG1El3iPeqFnXemvZKiQNUVYt4SbgWWzmIlgNbk8b5Vz16uHY08uSjIRvVOLB
m3vWzoL2QJ06WCUFkSOsNfz/dz2on00uQ6Ys2JCZWXjnpPsZEUEgC8W5mXN7oQ2W
l+0xFk7PVVZj1mDDpVrZwdBkaxyac4hPnYPaTxp6Ghcukep56YyAVQiGDQolT8bT
DlqBT0kamqLKZ+Wdpl1hSV5CYKSJrPV9tUfuMAq8tGD5qT/gqlnneu6gzPlztYB3
AiuX92DjOjPLKfwKaPBPkYAKd8QRS/unWT1Zx2eLxJJ+vcdsaBlAkFBt4sKreB+b
OHDAnIfanvD/Ut/9uDp10jqNbsPQ7kBHgylNso7PR4ijPcs6JGpTNjtXG7K0MnBc
+KB4xEl/7jFZZzJmLj1uPqHL8bx/Ou9ngLqdEtdyyPM4a8AmTGwsStkigxJERlgT
7ZBxpV1qBihaoe+/Mxaq3+flA1T4dGdn7vCu7xQBQitY0e2KduPUctzFl64Q0mwM
4zUZE7mbZzrannmwRvAZ3dhFe/VUuPf2P99JPZJLJAy5JJbZVwDxrfZ1efBL7gmN
UqUYK2ZO3EhtVVC/+DvdR6VJG+4GkS2L6mjkZCrjYBj8Ya8Zegb3TYJQAotpfgVj
t7yLnS0/m2oiek8Hopa/i/gvH5rcKrBIISQ0wN8SLMhdIJnHEZsq7ovc1drdfP5X
qRaTgr3B3Ilk4NFn6DjC/wRguZ0FYcRKOS4/fmvOVH58hfyr/jIFYSM9xhHFQ4Fv
35ZL7dH5NOHggbhfCu5GdmCM36rWjOEuWABjsGv9M/qN4pkWOi6b3GNybE2r4MfZ
wlSgT48q8me/BqtRRwuURQal6sPaiuhYfMqkmQH6+KY8bjY8Oz0WEvjaiiRllGeB
d7B5ex7aNtoVLSP1syE+JOOpZ47VF7I8p1jw5rQTJ++oB8oKNQCwlpYV7crxpNy6
P6K6e9HJGMMGewBiPRV2+xysonAkh3eXswYmusy9RleVCC4cdHildOEi+h4PGmeh
D9/U088WNBC3iGrb9v15RmnTTPH2LrW8OmvCbL3q1t3FB7jnzOtmMaQlKsxjNRei
LKZPQBY29/d38qZwwKHY6U7g5KSaShTFsUjbn4RpTxaNZUDl0+KobvVFPLzlX7RK
5giCUCWQdoo1E9PwPetUesjIx4OvDUBOufBGjQukNQyvsPoBC94TIKH7BJgl8SBA
Oe1CeqyZuy2hyes8Uo1nxcYVEQf6Q/+jATvQR4hYgz7jt2+Cvu+48wGCN8yWkgbY
nyqPZcMMob2W5OkVnwLyjgx6IQuXF6YL2bmnXe6eduFhgVbk0wBIA1rneVgo4JPe
btfcfKVml7opziybf7Yhy4eWF+vzdBxJr+KYPp9J5t9UpaiUKr0U0ium7Nb8FXTY
xPxu1zNFbDWQRb3/dk3iVaXXf1EjVvSI3Q7IT/Dz77Krnn2eSra9jOY078T8pekX
v6XB5MQT56QNOigh3rhSx84kGRC2ZLt45X1N6QBGWZA8JY6Nb7zKxR7VhRuTix/L
gVKrp3KtDkOuWWFQgb6Xezr5wASKrPcOeOQYglUw0XezQHzgrvkf0++JA5VaI3Rg
1ZaDPN/VnVEnXhHHyZXItJmHPm/SQhiAyy3xCNGFzAo8RgWsEaZnZ8mr5Ogk2V5p
iODGvHn61M6QYW8l0ravtdi4N0K/NSshZTHs2rIWpmIqaYosnlCEACQMfKeiqAFK
FHPbc3MMmZJsPqrzEM+lDxDey5+UFPHuZvBRBj+TPpna/OdM4VmCFl9CIhJ+l3MX
b2U9rHoNYR0n9spIZxHjdOObJ7kZ8a694ETpbJ1mp9Wvn/GqAFmDwSGDvgEe8YJB
cr9bYY2B+QFQ1n3lxtIg+H4IqfELyAZUaMrbHtsC4QXM2Q2j+b7gmSxvG9KCgev6
pCNUNfaUu58lXpk3s9wFfQlhUMLFMv7qfT1o7RELS+FklMPcSWIPE++tjgxFqKKT
J6KgWoWe5uNrXgANLgqiIuUlR43Sy2pPeYY2HQjKgzo4XhoSI7+wdJq2y//U3O99
dU7oJoGVnQu9lNJrEn7Ttdkd83E9fSYUHQt4nGZZygDepg48eo8OU6uGwje1lQR/
KHdv0GB1LWKO0I19X/+6klyqb7DoUflcQxz802QUkediFAX/8tYAhp/XedflZCpZ
nBTxz5wx+ikmRvykubjK0FP6CZkJLACPG3Ko3d84JmhY8d+Gy9ZMDZ2lppL3xA3k
lUre8ZJRbCGxkPKEEFmn97PV+zflB8mX0sBuy30lCaQaYhhVll4YDUdjc8NAEhnU
A+GLLYih4ggUi7QyjIxSeQ/1JLo26wEh+oBVV+qbUgskb+4NSBp65EWPuEeH/TaW
Z3RGxrqevqvQAL6bt2/PZCbXpIsQpjuYIdaaJ+7tMzhARud4akqBvEq04iuKagxi
NUXOB4MU/s3N1VBHoGRg3ZbFRrw+QrXppN+RhXfLzsRBijqAuuMX9lyCYcChv7zP
3VN/5dcOCUnze4GMXDQUyhYHKA8D0y62PpfiQRWbg8N2/fufBypZ2Q7gOFYtNVSJ
MS82mt8tUTGJ1/EsCCl6UqwoBxgNDSB4jUzGH3fDNuZhgtNcTl9+h0lQvZFkwcBj
5XV+N5iOrdv2NLI+nDLcdHosIblLhA+WNFrmyljIsqf1geOURUMWDwNUZyqE+cIZ
eGJ0B8Q+2qPwpewQ+0rtFuXnXbA1j4CO1lLjnI573yIOZOVTwy18vKL5vU19g5P1
gV1zypd08eiidgkGvKNIz6UAi7QDS9Mo5meQYs0O7Ski7qyGGbN2H2tPqI9e/fWL
rSN8HvR/COrArHHpHccFanUCjptWe7Ez814kjkr9KZWVkF9/QWb7/a5Lzi+mXgj2
Hhz3x6AV07bHJMOA7ogjHSQhbQyKHRSsZE90oxjWDprd8NOuicSPgLavdb1f+e8w
TxV2UZo7HOhdMALIbGr2fqS/st3MHjXVo0DZ/lisUjP+sIQkPHFcVrDaWWF/hHB8
1Srmv+UUssGxzdaK1ECGla4OjQ5Tvd34aGER7vnU/bY4ICKp3hAE+HlGo7zJWyMs
KdmSjWXjQqD4/zI+I0AN1jpGfPIExMkPne17pRoeUsT1+I4m+NXlygyDcMJuUWEm
Zxyv7HfzS45VL+7/glG1GDZ860Bglg8sc1h+krlmvNsiZOtLcu76jfSj1FwJetx+
EbaqllJBSJxZdKPpfHEal0luZ3SqjSEld+5Gx5erHi8D50uyg4ncGywhsBklSPe1
Vb/TqQOMefHs8gfxJtTDAZvc6jf2X96OwgbF0Mi/mKhK2CMv4zax3g/NEWv9GrNG
XBpJNhBcAgwmB7JaBe7JMQ+6RA1+7NjKTeW/uKwh+Y/nZiiAYGUEK1ATdns3itIm
tr9EOoUJUgqiILhUmxwhk+KF5pWs/toYdfOLOem8mDYdbHNSjb8VimKZcu23rlxN
rCe+uoeYEyO/kSbxrzjDHJJ58qMMzzi2FfJlXUfQ8eso0bHmDdldltjyKAOquHKn
drokdNWP92n33vIbYS7HiMh1AQsM5fbVPk73OXVSvRQksEp3aCU/3arexMtZ5GDm
h31ZwRs/dKt5QYf72mV97T13Bd/KJNl4++ZeZrjI3Wj7cHDNK9jjhtPM7SjlILQp
gFgHnqGx3O0X6/fYCl2ikmmUI5Y5HO2QTAiYtBSsl5H9HHlqu4WZwke5op9zsMSP
bnNkZ0F66bigVnDlPpVJoiVzzNaPXu2/grDSpOp8QncIT3VS64T6txScj8aVdX48
wcKqLfEBbzI98ewFccaRHIoTJKE2wk9InrVJf4IlEx27XSeCeLGVXVcjV21RTDEp
n/9EJk1WgrKI07qccLp9VfNitmiy/VsEcE0JDC6M9FtH2OAbb5I1LGUzLNjPipCM
TexAnHzbQnVQ7wJsSpbRmXl3fE9oDDfwEsTDfDAw5a+xBlQKwbmjQin1uhCjjObr
hywlzqp63Obsz2p1xb5EqDz0zRuStjuqsp2/evANXqHl0q0jSgTYp3dVzaGV8IYQ
AOrC1W/mHdPs7bX3jYiqmRSsg2f6ROuhZbe/9bRHmya59KzOuSFkD7WP+PSsyUB+
zFE7hacTSGrNcO6rP7IeXFAHJDUZ8NGAx22n9A6NRbGP313S6LqLWi2VOkQ6RoPq
f7URD3+92r2C/sdlpi4+q4CgPHVKxD5+6fukKUazuFucw3EqJMjegyvuBmLIKIm4
aLWz38NuaVzs3gVAckyA+/OjBF1B7jT6+AuIqHAH3kKWOQ1SxiuDX40Suk94fbi2
m1pOZG4azegM+dzI+CkCF4WmOHwBwDUZ21Vf6fCr46zkzS6HyErUgpdpwuoihANi
56qFRG5OoygqNm3AKuVDesyeR/jpKsTzCFRORncQ/B4cJVyPSHyDebLXuYzuLu7Z
ayOGnXOq1bUxLj3eF8j+P43IcSZ0H7RwJaVMdqFiZ5Iigd38O+kuMl2sF3iBpCv9
WOuYvEAfRsO9pmGZZU+wwfBLdSybXmd1pwP9uyzaCzAjMvbijGOdMixK6wK20MDC
LzjCxvVL4mOe50ss3xuBGURPCP9IcZAwZ9zLnoO5btTQRRCivRQ0YFGtN8F2xhcw
UrHQJm12CuxR1FBW4yHPl7AvKcuX67PrW6nbErIKp5XBDJHilFhzVZHWWaVTtHor
QQ/HCjVDP0xcjo/H0VbHLPsOle9a9dkiCHTuACtpun56ywKyEo50Tkm2WIpNjQpo
RJQyNMI0IEckJ5gv4n9B77oNvllwnp5ptPYuZsY5nY9+0iKDrYVgHOD52viG5gO9
au4OJRnfXGgT36952cg+m7JqJ8EhqhvYVC43ORKGiUCWdMtRwdFrUsRQemxGjtKt
LeTCMTDDAB+2XHutvRsIcQoD4PFxRGLExcLr0tEn3rCf3ij8jcLxNm2LQnZXCPv+
aLipc9rKKUgILv7RCww/DelMG6L5s85wPdGHRWZ1EOBvCy8o8UpAfOfOEzlz7qjU
wuuV9xwpEGNbEGcRuhLoO3X75iSIaFgbIsLMc7BVPmoXiLOAgy3Afv9fb9D2ZJrH
NBdDD6QidhuWvooaLRMBxUsrO0Yy/yK0c3rUOzbnSy3vZs9N0Y9xC+HzUQIYYb6I
DVMPjZfDMme7O4hWVEnN0s/0LT8xzEWN2wwI6qYgTQmx3n2s4gZXe8/5MT6WhXbk
HwtrT5w7DT2ZuqagEYFg+hqnJlgJh1BJI/MZKBkowIVQi9Ow2daXTJPrsAHy7hMb
BjpVnv/Wr55te1Av0YmzicaGeFessI0MlZlWCPAX+XNAFOrZ2uAhk4fow3kXkhXN
daxTQ/hBz6I13cNwtZ4iy/5S3+FP+kmaDvEaetQg924LYt/kD+9Q6XuTTOc/rKiw
QoFZZUDi1duAvM6I0NWmEbS2t5QaKqrWCIs7BOkqY2zZurz9PULW89okMigH08uK
KZFjZksxMjNKPZhHRdjJ6YVSLyc337hRXdVmJJiZlDl32QSY/17LiFZ+hu8EkY/e
lC1wz2DcfqNBgxC7GGAsjSpy2iPtdLcRd0kTcgWTDh374kgNSHWdKrmsnWZkIoNe
LhMe7n13PD0pIJvA9l8xuxBKjGOWYq8AXsD+9dg7ArsMz4v8yBj0C8mTtqI5x9g1
caWfTa9m5Cm8O9OyIZVJCqKS0sFR4NcN2QTHsgRfXsgNiN5wfjsveyzL/msjv1Or
2hbrUHcXEFMhahTagzwfmzbrzhf+4aFMPmJq2f/PzbkUBrnn7Fje7IsACjGuyn/E
6VOhAHZ2UZo8AdWl3E0LUkxa5uRC+KFnaXj6R58FH17gXSlsJLhANRhRFQqTKj79
uWYbSYfdEdbv2zbJSBkNtKTefhSdHFJpMLOyO6sABh2ey1F+Yn06QX/fV3BKaFVi
AoGHkMCC0SLryei+KmRJAYFvyVqBZE+hbUfnS64PSgGmtLxBw0x7RNSZC8EThi40
2P/i6pmjkfSx/6/mQ1z3R+39becQm8YveU/l5GWsmtjUJkyiGWNEgR2wDOY4TZXa
Lr5T9UjLI/uHNlqu6l4WwhXePc66dPQor9Omg4ZMMpQJsbzxpXomGUV/LaCmHWsF
mdUxZ4pmiucSrMoLGOKhbMwhd+V/Ou8Dr6ANN/64ifVfV9bLBNptoyXfyhLj2x4c
pXDkjcmtHdHphzJMMjxgwpQHPEq/iWBbQL8V8b2ReLP94UOXGczOsVOXMLkFhOpP
OFOb4XjAazQdn7Ah4ovACaLfjYFpX05H7+xHFOx60TS8qHXgdtChegCLvN6VVQ0B
L/Ylm81zWiD+84+oRkaWbkSIWJZ0wH0F4TGgZk63nwbvX990R2u2+ooxOGKaIuTg
dWm+FqQljcA+J5hmkPFdi/n1Rw5guSyEBm5HsAEsDjIO6TvLMx581G4pgEyO5MSi
iH7ArWJZ0ZTWX1DmTmJzKPkMd/uQZ9xtSVlPlwlWrDSLLqtloCKgfUCJOaDKaBl3
4Lccf7gL0rjLk5hIEGL8vBypbgDWQyDeDB3onf6cvE5pnoZvsjf2op+grZoBZyAc
pETPhyUhwxLonM58eCTQt7xYLoyNlcy6i0Lrvy0EGwSQiKeqytBmqbaWiKWTWflU
wqqUMmizPwyRJxY3a+uQB+VcWHCG0UulF67+cMqPkfYqRd5PQ6nSJSjenkDFQW3l
2JveIDl1WkH0FzReGYvi+tTAhJYajNuZFdpazc79tl8YWbvzwEnTi+zFqlp/v55J
KnUIjvmEwJLP+EqwyI2rUB2Wp5a1CIBPCDsxBi8qlPxQFh7v+rexNG7u9rbnfhfb
dDm+NW8CBPpBGvTPDrHVkr3SODuWNcsgpLJyc6kF5q/W8s+fd2KmTJd4Q1GqLkVU
TK9Xi8gDyPViu/vm0tIpmMN+b1ALvB6Wh0UVeDmCPMGA0yO1rUI5ybHW2hrQzWMf
VKSHQZtRQNbuEGJPL2YZrLpCQBVBkT/qXAZL2N0/mWCYw+r3Eg9HYO5i5r/pV7ZC
hbjv4XTGmoJhkbSXa/xU26MDS86tumykC0rnYuHZgh/jjvRTQF0IUyXzCABrG2ma
0//IMbJIF55OOTHXo1boz7XPjemdzBlZR9ksxN5BC/OLMQ/u4gCO87rDpe23i4NE
MFTQhEvzBDX4MyHjbqJMC6sr6MQ7EZTn64NTjnNwpx7S0veXbPCQ/xxD7vae3h9z
g9itST2SZpldgLGENltDiVX+60ierDT6x87MRLPl05ocBj9X9Zs4p2AxmCnpX8B7
BLd0nVqK76MPyRITwFGvqe/SwuOq0PGchvIRQImYeOzAEBgcoElnpRe6QxvnROk9
upArvLUdPFWWT2oSbVWG4Wci9ryRQ2qRG4s5DlduG+g7QIcZAYbBEG066UFXgLEX
4Ftj2gS24AzEMKYShBM3f6nSGRfBgFF0CX89nFjSPzqO1woBz7lM0eaIMX1f0z1A
7KpXb6GIuHM86o3pJtbAoPhWd6/6vqgDD4XxfL928/Vy2AxCCyyk4ttaGJJVeaLO
/G64y/G0tN39GIxGI7dWBePddZ6JE9AWOhGs+/90fW8P7PtXjLYBV3K+Idd5ncfh
v92blcvrES9V2uY5bPDiodSl8XeDxVK02aqWtVM2AvKy13VmlhEtAqw2sxm58Yjf
JErJVwTE+VRQiPeZYriVK6tUcgqFr/cTwS7uarmraEM/YRAhfHVPJK9Afuc/qNYN
HYi/Ln2Pdik70/Nqh1DvhFDtsJlukSr+CMF6doHJg0RKC3xJTIfhfd8kCl2TAOA2
WvPVq/vL/BPM5QFmolROpM5vgtjcEkRLXPAzYaAr9eDSTmlV5mwnuf+U2/ypBP8d
qvoHi6xEAdRzXzRN4hTi+vF6pNFOY8AGhpaTQY/7f4hNCk10uu6w2w/Q25W9Ce7+
aCaiqdh3sjbQhVJZFNpLgdko7JFGgi3iykrItz+5Yq8xnEvNw86vW3VEVmj8xx3q
51bbIB/dp643jyw3tbrE2yU0OBQN1X5E3plOAkrvjqzH6xg8Jp7iHU45SGXNkaj9
gNt9c58QrotZgea+gnlZ9Rl5Zc/RPnVpXfXPocTSh1dtfXmG+J70kJaEXklhQ5v0
v202LEzpaNOkWzRIkazaEFuLdqukXo1h3e1KTBoO2dHX0WyJ7mmRM+jVJubqbI36
uM/Zrq4xwuSlnWlvCuigqgCfUxLMYN26R78zE/z1UZ7RE9QXH6F27k2BG74BUZph
/z4j50oxEi6/5KNOLkyhjp14DXBexjh0Pd4AX2N/Ep+A/KAXffhE3s3JRlj3xw9Z
DEQ/ixbDivFBlnOw479v6zl8wVKaYeSSNwSbnHQRGh+/sBwxPkPU5PrE1MVnWh4G
ZPN9ZzjZom22HcNzMFJlTVAi0QO/ToTnw1qexm5ZKIXEBABfIpa9doUgHZMehaX3
z9u3rhx+7sO0WIO0PIVK/istIicXbEVNnFkT8lCcji9cQi9GbMHQsp7uSCCJYaEV
W7/mz0HyRf4P7TGSs53RcpZnsV7ytN0Li/eSe4dlFqbthfdKyjx35K2x2PfFN7XI
yK6r2zU7fWBR8ompvdwq2c5IgF6klufGhSS8nSFvlKHeoKFpNOMm5MBxjqjBRBy7
gBpE0J9Eb1jBCAAeJGgR2r5k/WqOUfwJ44cppPAfUqLIdQT74oEut0aSLosKTOmX
OEUKPeb0TsfmHYifhkoJOqVss5Aui+/24y+F4U7MXDbLccm0zw/eDCEWLmK1ynpB
LKX053TTdwsCJkExmQPQnsqQ2I0YYmJNGQISUBt6seOIYaX29SFi6zaYqiT5G74q
pzHbYulInAGQcblYE5wbE0+6dtpdoJyX2LaQskZO9nZVAPQF3DpmhE+f9Sp3PyRF
0Md3XGGanhDpxt/Y3t2stcgc7q62gSa+XjhCjNacgXZLQKIKM9jlNBIL6qbjlVZy
0c8DQ0t3vWVsFKVj6do/MpxEbNL+gafZjmAXpebC8shYo9zp6xKqwYmOBJGUzMjB
cNWaM4ksQZYFWTUecoCbAEO/N8JEWUVbkm2JtQUNCAeI+yhLG8HYs/5+okzxA36q
287bS4JPHPARt3VEPGL3Sqy4f/0Krxv3cQjuCMsufcLIUDnuKcE9PhFPU2bbqe4a
eW73agUSlxcEIuW7AAYQKLXk0G9bNZO6Lo6nD+xUFZSN1K/d4ifH+trDnIZMr7k+
HHuLOwMNjXUhYLoF1TU+SQqVqyiaRLrgwnWPlQ27wGLv4870zs8lZc46gwhADlV0
mh+Yn1vL7ctEMhpJnLLgBcvc0/XiplRPexRWvNgzF3zTIYLqGO5cSOYMI70UDqGC
2Q0NOzR8NakGyu+M4YZa34z0r2XP0CF5SvOdjCaUHbcipDEakw3cfSoaGhDxTIVj
/N2tX7AsFXkitH7iSlLdcIjzYKeJCYrWgAicsjAo9t1lh+gbuXBTAlS73WilE6n6
7OLnYl12eX+1fberJ4hIG8Llk+JDI/fVA9b9XBoUyMpBBE4B/h+e+ly01PUZFMpn
SuaABKt6iPmTdZ/jxfWyT9Gtiu3STgpyb26Ad6ad5djaq+qTOQu1/8s8IECHlxlh
Gaja6D9e6GzSAgg/+H/839KspvWnXzpwJuIsPqifRc7aU2wPLQjaxKY47dW1oGaG
ugQUJ1y8Sruf0a6TBWuCXukgLUy0X8aICskhaTROPDW9M22AYRc/aEFBFJOB5dwm
eH4zj1MGpJGeXUmzq4/XB2Lll80W6OUNt86b3QpqGxg5xv3Wn+MvSqQ7Fke+Y/iy
nD6FWlcVf5iH8rZreIhVrxRT/XA1Ih12XWLLWEa4yDnDWvXsbG0v40kTw2vZ+EsO
C99raBKBypwmRmlT0qhhbStNaCKjTZp2vYDFHmr1DlJz5ybqZHEbGIk1zYy3kPdY
eW1ZpZf/F2Zk+w7RQjg16KwiuJEYA+afYdjTC1FTM7piYrHO3Nb5AJEAKalZ60I8
nQxH0oRSdXqCW28iAx0M/AM6bwpgwDY6TT/Q4uHffMEX+NlyINNdvYBTZm4j2kZh
NASiAO9ntNHsDREoHfTjYM7mBreyzywHyFConl9eboOqHWsffBXKDcmgQXF3Fjrx
KJB+b8rueLiKPnE3P3FHJoOlfqqqmo12unokLvouKL1nvN9qgDGrtT6gVcxJHlf2
xjUAXXP7ptS4am+eGbwA44KMvIw+GXFsb0+zSbm4rMtt6ep1Y7sMDiYb7FS5jlSz
WeqzlMlxaMGqOC2yDFLnWDzxxV+eyqpDDebm+ak5whD7Y1sqlleMGi33jbPOkouU
ZnD2FpEmwdS3oy8bE+RjueGIvBeZXooOEdYrECqBToxLwtxM+SFLkvoCzlUFFaXz
ffwhUxuiCS2LzsgTG+OqJXTcMxxADdtjNs+6ClV4tcz2O/6G2EwjfCK5wuuYx/QF
rwamMdZ667XxbAVUIxD8ulFJYRw9/hlanIxL69YBDJbsI/pvKQmiyQv7/3KOZ04s
/4UnwrMGZlJaj0QcWaBj7MRnfaG3JGSjeaBnANZL3/CKJJhxk1qOiBuiGYOSXKEO
XnxO15yqMGudKb5jDY4BuufW+ZnU2Ntkr0aQp0W/TLWbvlQqnHBHeWEK9j9Syh6w
qo+Q0ZTxthJcnpsToxIxfeZIJinyFFxrPB/jPl3h48aolopeeYuE9qWuKVp3FZCX
5WArUsLwD8xslW2A3xPx12BBYs2dqCkqgf8+G4i/v8PpMPPpMTF4FNg+YUSTny/c
+LbkeWbMhFe2wYs5A9JCViUy9dGELeccxsDbCmHguSZIqbpMrQZyOQAZIJsVT0Nn
embKOIhovUUsIbuVmkS85ORe2KG6qKED57WeqVVqKgSUZ09pWg/xD4xpJUU5iBLW
JKh7a14xFQVKhN8k7fs3tCwS+m8NGJws9juQpfPl4cPAdJtNMqUaV3Q0HAtTFG11
nBWoZKYtbBT+fV/1aJfnO9k6fGgN5kfULU7yyrCJfIUtHD3HZnBVYk6nttQr/3P4
PHkWoR9k8xX/y2a0c+TdHh4/MkdGMzzeDVk7Gkl6PgfaMObipuylPNS8KTyPROG9
extgdvyPlibJj1OsmvZzFM5LNn2Clm/yQ9sOD8jVJ7WuJNhgisFrrvZ4HZW3QRKP
pOdcwQYDF7QB4POhwv6nqo/EgKu5bXKBmx45YaWOyuiiRSSSnQ408CbvhKd2nTvI
T9BZV+75hIQ4oVSE4KF+cKNzkYMhHEUctzfCJkgFOrfLtLYeOruNC+IDiW3HeIoN
YjVP91vOtlZ6ZNmE9iqJW0zJdJw6JB6ujtqj1ct2ffSNSe4EBgVGMw+b5Cv9n+wo
uQsosKnV3jbyse9hfjY3roRAIhuFhY7KZf9yQ22MWHMBdxfWXYbx6HUerIDJsSiP
te1B0cA+de0nAhOroRZgMWmT7PqexoG8FnQkNFtC8gnPX6FsMyrT4HdlJJ2akJgQ
feDYZIDkDctIBs2v1HcaG/GFYneFO34LQG1T6ZieIk6YQfraUCATMpQDWckUbwWN
Wrk/ev1R1y0zJC+Wx95A6P8Tjb5zVnLACet6LvRzLl6KS7k9KIzomNurgoUdIm6m
vmIHxqtc56DQglbLDNLWiYfb9ID//V73+LNypqgHor9zA40MtKTTqRbbcxKO+P08
sidsTOV6sVeVtHXWhwdKnRfnPM1DdfRcLzaIJMOKLYHeIJre0r7Woxl5JOQwvSIS
EdpeJbwel2praSd2hh1+XhRpdyRowJYISekJyzR5BkitRNw2ktQ5/ApltBw0BWEq
jaK74FjLEXO8J7HFtvxuXgEm+B5wDMBkMIuDbbfzCuROJjSEb2ld4Q0icO9cxsKD
8/CCP1eeX8X7wZ9GZWhSXabnefK6Y/u+1RgnvOQ3iFUUqphBFqPjb4byPc3iHK0s
2n4S5CABoIAz20lXlS0LZYohGi134YMUqP7O+bBA48bRDPH4M+auL3hhZ0Xf3qd6
LUXlA+4saZ5yNklD4pWFxAvxzQdNw3BFGZo9d52Iu8UAoqxxC/aBKYYVTLtBi+zi
DlnuNx7bKU5JPP1IxrldmjheCSekJ5tNqQv0FVeDji5CZrna+9oFO1VkLFB8be2l
1TY98HUWdZ03UMfiPiPuE83Bzg29eNFs3DtL70iuTSa/I6TZYGHpKY5VCjdpYK36
j6D3ACebJ/VLkvjg7ZzJSqTFC3NArUJRvgNznW2r8j0TPZ5BYmdx+gFVFl9y0EBE
doUYAvt92GrZ3wWY68mzEPMMqGb0fu7PCE8E4RR/mtXSmzPo4HJzdsdbV+Wo44FP
8haHrVAxZZimIEgtbyiB2sGuRorjDSIOdRkeBBJe7ZyebLCmxoZrqz3B0Lv+uhwp
XSEMccObBnJjCfJn/eH7EuQkS1GCFvJokqm9xzJMbTcHqc6E0kTmh+64qBwIJSv2
C8PQSxZw2HJjEe2GNA2tCJwK2ZWK578PwnwnAOEq0c7MIfDiShbqk06AuPzh3hYN
DgDS1xW9dzqXaRuTFBMNhcQk55XeMlp95x9bRF17btIYcqUf4GeI7TjdyHGkfWqn
hcFh4PiCX1YPPPDjWYp8NSKwYTToIeHAN3hQ+0PLZpVRq38/dgBaYPaLOy7hbPSE
5Wpk9rC/oyCArvAgh6LujWzkLPgaJRBii/K0RLfviAdUfaeKLT5rSFPjBsGJ9i3G
JdnYzHdot7z+0z6rm1/2/KdaWlAO3s1jCYlYprabgBFMDi9V4BrH9ZrMX7oPoVY8
y/mnbjKjOb0eqQiGXcLMXNuu8JZxsfTkHNOOYHEvKI240ROLpbibo/3H8rSp+Gd7
wwu50S1z4mLZ/VsD1WJF05eopGyV8Voou6lSizWQtWG3gIoTTxgDazs+h97OafNj
NnakOSf+FwaGFJm8rE2pmSFALyoIHHDQdYsUTutYd7P7FydsTPLZL763mX2/Cafy
DnOCgcntWy8gM+WhrLbFxMSXvRE2pLq6NCXbkL9RpkO+/dDmZk0a1kDJ6dYCwknJ
DTDZarl9kOcCZuFPriJ/67ik/faNio72DSsIvcH4usPVGFiHr8VS3Q+oF5/9t+X4
WVx8SQHBAyVh127VSeO2dScddSrBHpnt0RZn3Fsz4Pulck0NxLdxLtrndPeuHkfc
b+zKZVNjAzhOJhE9KR/YEUxl86RFFtRvHFzaoIFHssr8tcBlyFCO03o+o9Mv9a47
YWL3JqSwKeQ7pPNB5Hzw1VB78T5QQa9KVhhH29Z4GNcLEhXhbm+rArLCs9S3Q/Aw
RRbF3F3WOzBPYkQk7TOtsdza19cDgS9tOAjKASb1nR82hSsBIlR/CLY4lMX8MNQH
rRAQPnSZpQL/y/ikVBCRxL67sUck+mzZaheZJvKvCUDVU7vmfWSlNuv4NwqcsVHl
CXH7SVAHcv8iLsaHGevpi/rIyM2zrWSo8Zn0smzvg75T3cYCBPrJCbKDqHeAvhvI
LmleMFeggXA5heTMf40xQayzOdqdOZTMdQ5RWdDxdRyHqGkFNptQDY6sVzWUABSZ
FKDjX+pDyv/GPpF/NeeP6L10sn97zXuJixZ6pCs6RTXVPRjEkDzk2iGAxmuykYID
1MiEF8PfjmAUfOiDAyvl5zGc49lOGSiyH6DzNaMpf/VR0Cx5el3UzaJ3MEaZipdo
GmkF1CfoospTofLZ3v5fhOiEiGIe6l5lr3nlLU3tvwRam+mZRcqKtVbT9Qum4Nx3
OM2Epcz9RTbWGSIlgow8Jt5wd8E3WOmz2Di8/W5UWBr3XgQBiIVbkkCYowngvQcZ
fg+L6GYTVT0WjjWinPBffFI0yEFOiVL5N/y4hgYuJucZkKQGYyngNpU5VtlvHGK7
ZQBKT0sPuq328QBx3K/yP+vn+UkSHU5tRm1kOVMiu2cz2VrjeROdb7wQn1SlWpuP
xJbV2ZxgRg/5kvrHnRclthnoBIa86B0N/pP4zDx78s0ILxweUtuiCbGssH2CVlPv
I7WK6Fyr4mzMbwvXcR2Rc9F5HX61gqVoWepW/ics3QH0utuGj0rzUynqyrlon0nX
CdTFh0ABjlKv810b3Btdhd/60LJGDugymvM7HKGN8BA9D2NUt9iru8/yxa56sQo2
5JCJCdnKvtqewCSxlXkpD/Li1WVlgyh0g5wX2GOlv+rCnJoxCMdPAlSJdXb/o17P
tt4rSMBpMpxawY6dAOmWmVmCo6fqUP6NYYpa6FXvYD40E3x3leX0abzYco5vO7P3
D7Ai7+uU89UKeZuAEMsPp8gdKX5Po+xc9Ar25yTkLgd5KiMV/2XY97IIex4+NnF1
xznUEb+t7SLhy49M1coDBxqT/l8IKPPdRZdH+9ZMD+VspdVz1ZVN8ZJovvNMX3q/
oKOD8Bx+RCGxFZDKh35/Xw58egyavvp2teUU5qRhThVYoDitxwBfAKNDBquOsm9+
dGdsjrTjXBG1kogCv9KIHk63hvvShsOCnxeSWMQUsNCROAvSN5tCuzOqx11phXaj
7XKzn7WLzDxoZdIC+O2WGwZrHzaunRYnPE+vYA6vCDX0Wz37HxUuAf7vZWjmaGRK
OH0EbeRkfym2+QyR9FYaq0CZXWMz6ns2y2h32pEzmJkVhaPWDpithEFRX1fSUeds
tfXE6/ljHboWUciR0dP6axQSO7xsZwYLuFGMxCCHGRUFvsQiEj+B9vpzcRGZTIvp
TLER0hZav9TEqP5UxHyS6OyOBRjGd+Aqbv34NCNvb0fSYhA4v1eiKG/R9ZR9oyV2
VClGhDG8syGdrim3DJdDCGuS13nIe+FMHvWtAAhU8TQ9CmB+fqPFdT1UFof8NBLQ
McXPaIwNy0GfYTkZmM+L/Q5Z5LcrHDBfXtsUMpaJHFo+ddID6DXMDoP6awyaBGrP
2fSmHgkhd4v2tbrUXKJH9oi0HRR+i7KA1VPPbO+DKTXbrSGS0vYknHq4QIzoz4IC
yntgBNmLmit/dfxvddhkiXFwRPctJzoaWiK6avawmRsodRtosrdtB4YssSDINotA
6CKRFY5X+/N1UAq2e3hbylWCBBRoGKt0/eJPpfXO3nA91S6wIG155CmIEVPNNosW
kLa6j0LSxCBmyGRzpJkfBAtrf3z96UUqmyHEh9gjF31a4Qi0rBjr4uAdh1muqJ1T
8/euUgq9JjuZJls9uKWTsZUPMR4odSo86DALd14IVN28zDpCUIf1tzSjlpO13qDM
DLk8yQZLmkaL/I6pV9QZpoUutvIbsiSxdNE3T3zBC+87gGPDiRA+/LU/RxZ+fDJI
1p8g7X+Lh2gd8ksZ+ra1eEtU9qQsja8g/tHQPc0mpULJHgNy/65mkIEg15nQNf85
54UZ3TRWoCH6ZMYmOVJcr4VOQkrPmawHvpRJ1uMLOwl9QTkE3P9wPbT83iRaC+RT
u3XqYOaYiz0pFYBCaePflMUUf/7PUS+7JryprDkOs3KrsA9Y+fhYvUBHrKgFmpQB
/cde9rBT3cJi8zpdmfQsqkvEGcN1qnc6xfW++HKMi+nKHFh+Py9ADEsrKSUI2Z8I
/TgJ/IU6aZ772f/AlZ6RxmtszCo9fvUFPCHfGU46h9didAawWR5HSFJR13AVNfQd
l58vBGpOHDFaxH+ZFTRNZ3rK4eKfflt5LDhKuVCS/UrpCddunPF9v8Dyl9pCDYqM
tCZN7AXyrtAKc5Ydiqvqyb4vsfpGeqoB9L78RrlvAXEqn7jmzlKNRRe8ZX3xjHF/
mXb8dvcuSohSmzlAxRkBw/9AMpYyU7tthV4KrbbwYcgaIZIg9bBP8LlvAvS1SMyh
jsHWboPQyGNyHZ9xwFIurMje6sZ80IqQUFn2vSYKUSK0R9GbFGTGHx77NX14PrKf
xZDdfdr23ji3BBpyoQWj9pdf2cX7D3wNk1PPJ6t4mI3lsrUna1bLbqJT0S+/2fHz
spL3/+ga/YOUpYDjQHIGzM4MwcQIJPeOlYVDuAl+GWboGEwW3qlhMclZJUfSqW/M
lzk+7HEi6ZV1m69TmRFtYrN72GUA+aHfzTdVe/osRgW3Uz0e+U8Hk4Iz/kjr5XBF
yWkduJ/WaiBbBtCNwmzcEDxpuRURQGUT5QcDZ65RnRHRBw8VPB01jm3Km4wMGZYt
bNAxdCRIWuoujY+HOVgLhhbODtHu53DLRdO6MVDSckL/wq2mgf/JFh1BM//0I3Oh
L+c1cjVbayhD0RlhMlpVM3UgXny0vuh4JdJv1kjBqILL3A3uqSXAwTdS3Th9aZgJ
k+cVw20ZD15nypkuUTbvaXZLkITJ9xOECsyaHp8o5mEBW+JOYVPiJPe69c4goIYk
uxkYRggLFGX+ugzKl+Rx82NTo7q85kjLSrbCEnxyWz+ozL8v2TyV1K9096sgTnry
jkgErfbCaijypI4YFEeoXTydC7aoxacSOyIfRkJmIaIVool0WsMcc6/cWGpTQA3G
gJMPOrYGZdFPePBQlvNnGIoofI3r+8gPflQzgAL5dKuOEXmJ+0W6dVLfJjIAnmkI
IgmJiXSln6jILtXcOZyrZ3fIra8ZPRt6m3eAYKeiD8fiOK8jarvpBX6odG3cAOtl
St9kiXZa6D3unujH4SrU+WYlY5tMc2u87hrckBJsrk2+0ufuwYraeefWnIDCtVnN
OG+7n9YQ9jlKak8HA2BrMRtR2QXgS+yMWyvuim9dcdhiSm69uiBBksFl3zPjfN+Z
Caeb0dtob0D+SUmRRi3S9aT3auKBB/l4Q/jniE7loExkE27lD9prhwC85MPWopdI
2AC/h//jpwy0vRzhBOx0PGVHPAdHpLC7KIRzE4ZTVMWZT/wxZGdyMHtcJoAMIObh
B8sMveBirL9jEPPJ96aDQabEe/VAE5baw4kzB+zcgagLuqHycvA5UJb31UzjAFiA
7fFKD5piD4U6f8RaB+7WdsPFacF8QR7oDA/BEdOoD11Dgt5Sex1TDrceaLo8yVtX
/a5MUmuj/iHK+xP96zpOgguHsyU7q5BFRUTDlRym8X30tgLTPBlbOPCg6UvSuWG8
nBCXhxvml1jq9Nk+nNB4qnuXYxG6+qTsBYlrd9pSerxPYM3Sl2VjkXMmfSMv/fEL
qKH+9yRpeqGLlPZE1xglcTEsX/u/GkxObX7LtkZICZKysGtBBoms0X2CRnav5Woi
b+dSLehI8yxF5ibyLcDTcoLy7tLXO5/Xlvv6mksi16kL+5knwJalXPQTW173Fwtg
orgRVhgMcxCn2l8hBTdo6S3XTZ34aFxQExoKqTadQMdVafCW4uBe69m9+MzRIB01
/uWIXZs2bQuDvRJKlcK5B8SzX3WGL1mZtMoXcFvb1VrX4UuboOxIQcPVldagqt/B
O/iy1AsR6clRpB6E3TjcCzTedkW+4Fgb55oq5ZLDFx6Y/FBdzIHZsEpZIztSj1KO
X/4L4+SEGJE76RfPCISJcITM6EWuMBVR25dgELHmXtj5vekG+dpK62L9o6NDn38G
R73U/0PukRXeg4Z3KwIbCQNiydnqUIT9ygY3Xc2eVCxsDvdLRiHpu9gzbftqWqcz
4xPOkcjw9+52GvJyc3y/ziMQ165l8LKMTo8bsR+CxXqDRSDVffdAu0EShZlrXmit
FbBuvIR2ujYS4HY6sLJrflKlkOgY63ARyDkrvuc45RHJn7ucsh1j08YCKYGYp5hd
R2IK+USxmUXfnn5Tyj15HwgzQ68xNkBZj4UzHj8TSrb4Oj3h8CvQm5p63qjzR+DF
Us6DsTwEfTJiq2j+PTwq9gf0TZ5JzJM368HQKHIUIiG4yL9E7VfhT23d/cPDWtvL
SXgzLxvLA/sHwYURzZZXvZFhCu7xgV9EEXcPYhXV22kR9orHTnUoAYQwX11G/sX7
S78vBeKDzANT1kRqTtSL81F3IUhLBR/T1bIrKcoJ/XH6uvQ30aQUUIiy6DkNEPta
wJnthkiYdWFGlpK2Wj5ewLdqXRFokvvPkvFvFDFMhbs9UGZRNk4V+KIZhZoT6Zc6
SzXqI4u/zUI15SJKJuDpTDa0stx6CHLVSfAUo5b9sZ8Td6anBi0Of8HbicMUwiM/
XNCDU4GyaN3YxGYZH0kkZycxR3Iijio9v1aBKMk3C3hVFXgG4+w1v3mg/1l46m9t
GyaQE3Xf9z52CzpsGPhv6i57/6sWLZDJNljq68JId6r2davdpDxxLap5wOZZmW10
9rBAcm6r8zOZtNaYhcs1TrLCYDTVoTZ2N5woM+mIROprqRwqKFiDYidAf0NzoS1C
b1Wc80HDQA6QW47cS08nRGS0jAFZpdXa4i/1uG0L16FjHZRyntg0+u/wcn1738gC
4Qm26Z6eMSZgj+1gzseIyy+eAzcd8bAAXHPtWTN84FePw/KwJdiVoPVtR8oijFEs
0+IvEpN2p9IqZ5gqawdRK5kDGfGxyY3M642IVt5dwEnLUDLEgZfNN+Puk4/LTQdA
B8hjp6oM+ML+3T7X9568++xaLU5qOeH9Eaz3Bx/Eiqp9+3ulJrt9/1DXJnvaeNlM
VlH08/om/eC6G2ANJj0p3FN2PGjCGTLXndXMRepaLBo+32mG+M9tpZ446urD2dau
72j/Sf2NSeI28PQR2NQPbuieWztZhtYT60ZO2mBPPPaxSg0I1WrZY2Fdu8pxkzIL
fvWzplmkUtZsF36nl5usSYTH5f8LdA+7SCBjC6MsnmRDK3VuCz9qjbptJdjnRPm/
Rn1FlXpWtt9rPpiMK5dURY9HnQSfi9yz1XW4qrfwhKdUuzXP0QuOBJV+7HfCkcb9
rP9rrBZDVvG4fwkAp0FYAaM8fgUwYMotSbrRvhtnWK6gfRLW5xZ8Vgsfn77tAHtC
GzPvd7pQ6t2V6IkZ2dnZ4XyzUaN9NAyHwcyXuqQOGg2tzWYsHYPlUM6Pzq0syT/C
IAdyW/ggo+wT/zOmsYo0vR5E+w11InKAODPoFJxuPcea+bBJxu9A9sAYaXJrpz3X
KDEki4SlfcJxbAMTYwm1n71/xbLnm3B+bBN/Fl/aWs7+nanlv9yYEJ0tNYxxcRyR
CcjojWeEE8HaKHNGZ0OsETAcxZCBGQkvSmxt9CyEoWqYhQmUZC0oxtQa2iD5s1n7
sHiuxV5egaAaQqL1hVcy4oVIpp6KcmDxAkfw6xnAHJqEPM3zXp//Hjw7/D0tg6DT
Q7C8+1UjthIwQvUAHxfFFn5mR1F4T0CrhnN3Ow6oiVYoHsOFk56XY59R+0E+/NFk
uDSKdknE/NKpqBXL07WYBp3QKN0Cxq1XAx6F7x3WW9u/1e6LMS9LzQutWnwFAeT0
/D3MR3VSjMPt3lSeHMgHM3NCo1VDhJXyZ6p8ARaTdgWpJjHCW2wK5XfEuKpZbE6A
mSX6O0x29tPIkSU+U8hjJvGiRyCVHXQDSs3qeSeULVoequA0KXSzHUkh8f8GvAxF
NDV1DgKsgTIhGac1LWmyNE6bb6r0cwVvz8lNQUwCEHOLu2AbOxiY60nTdO7HH6bN
JDtskmhLCzRSEviM2sX4c1VsvU51Xk5yi7CBJuOD8CqQS5J2xsbYD3r1GsFWAXUG
jy3LM5I1/Ha6JtU4awe71jDyAlinJo7cOY4nuyJlIR67brMv3uPY04SV0OeIuusH
EZfmpMSlqwG2ynkez7vtcrim5mNZ5tsl+FMJ/VGe84j4jiI8KIC9jKSYthb8TlMJ
bCAinQ2RLblku/ZNkvmeP66QbEFwauHLqFngDsN5pOdGWGLVvvZvQItwLRnoqLSb
hNly7njY2iOw19wSOSM+zKlJXQmORb3cc7EGXc/IZOFPkzKXZP0Bc1t6vrC9oNx2
X78br4OITAShVako3ri9g4jweB+DeeGzcprcy6MjEA/ezba7TXStKTno44oO1uYM
1wiod0qP509jv80QDJ17uYryi1/InFt8ZctKjJggns25aI36zNnzJYC34H/opwQG
O8KSfmaRzWFarwfjxL+KlNtJDOdx6p+xeUUhb5E/4BCSjaAUfK4d7lCerhWbAL0K
U8hJH2PjJLHYc/EjQhW9DYilXOdfKtpoLV49CcuisUopCwuftB+DRvxl33RPAYgO
Sq8Kprigp7Xn6RxQWOBAR/cCGPx9cAkGg/y+5/lxY2Gfeg8wwfriY6ffQoTkNH+g
suJEh1Xbr0i7/986XwXqbwejE1BIi78O3T1I6sWoNCGm+FaOAN9PzxWDGWJ2ADeq
Ue7QLhZ8WtmZLE61JoJ/3ebzUh9YNcCcoVdE7RDRoPM/5OHWXeUcKti/EHZmxJXr
GQCv1P/Ws47yKz+QbpG+8nwu6w+tythaURSrhNlsjRTNDjC3Kk2Nz02mPM1Uqs9K
7V6AMZ592iTVVgZs2JeEsvcQxDPl2yERwkMw2JNtbUjFi9zIwq5cyJ6ZiWeCeve1
XDniGpMq+h1gB+Blhexzr0q4REvheF8+AGWcxUegcuxXFV1AMlIa5PmdQfR1GJoO
xKDvJXRqpU3R6Nxu/jOgpYeKIBB9vqWq4n9Q4f/5wAPiop3wj9JiOLuGPN3JzGN/
dae/OfIekiFR5LoNGF/vbTQCLdBr/e8YQvCfSPO1TJ/V4DvgLee7feLfBd4lRRmZ
DxYnGyGx/hWyvpMaSBQlXVTzFC8BVKwOBwUEy4dQKPIKsh3T/wO5auUNiLcZ0Oaf
1qkNgLbohgNtfOkTLnzUmCPak14/PxnjTbJVudDrg3X8PwlTQHxxJ4suqvVMM83f
K61Dh7HlO4dwe88NmZHlp0DHjfd3iWoSki/yoJq25ugZZVYlt9wctrnqq3Brll58
FPfHc6/UhzWb/BRxh9bL0tRlVJTzB0X6dt+J6NoVr4cnumLGy2fZymX5pVW1Gv1J
IHlnYQn9xYwz3hK1hEdr3TaLA8zFL6Ph1gmzlBE0arABlrLLFs8m4eR+CzPWcQmR
lXQ3toq0irF3WxFl9u4JzP8G1G4MKEsNQf53hKLIT2tdlqbRbUCSCMf664S2iHef
ZgDDBoJeRZ9Za+cgkPa8MzCP8jPKbYLRZmYbXcGl3uBFrfrj9ypEY6C9kzi7rpWj
JvJEoHwwkMuttSjbzOsYs8BtJl5pVMHdySVIx9ZAP7zVwGi4eVE6HCoS4P9JgzZK
J/xdgF8GHXJJFDutq2Y+MWpHgu8XqzN7gCrTyFgV70xaMZRMmHic0xv9s/VNabSC
bg1FlTAtPVa8P36Z0MpjeOutz/mxRld249MWLySlHGa6VebvyxmMeqZX5Ua3Bfps
iXj2gZVG1jJyvViXwigy0TfiXZ/dE9H2nU8Ri20Lgoch+QoeFxki1Q1jEo4+0dgM
4wq3YN8Qa3ZkoNaVluoRDXIlzuX2gPzF/GYKwg0Dg0mZIUzV5JnnhgRjGDkTvqEz
zt3DaXmxwA5aqAf85/nd+YR4LdnMBtUKEVEDaT6fD5WA5fObI1TwwYKptvz1PGSf
4yBFBgFFk9XGJ6qi9y8UOdLbE4tUpO4n/GOjR1FkkQcF/tU9tR6TrQgvD5g+bUkz
ReZjamK4WhTTRjIZzfCEHMZCLECCz3zzQdHTDz7COt1kL8V03zoZgcWGyxjjICXU
WgiCZbxnyXl2+2toFZXrfmjZWpWYkhbLb/DaEwaNRZfBCLb7CtRU59sxi5JJZt0d
ykPlOdxhaqBzXwJ7S3Kmrj47wAcYUnySvg/TIk6Cln4SXJRawZKqT6pWq9WYedMe
zsyMOZ++r9cYvFRVvUeTaStQSP04fsubyz7gn/gj/CgKRjICyLRYaoiUzay9a6zi
T7sFWieHUIML4a7zmkgQ2CuuJmZ35pZNCD5mzQu82/KalRPcu3Vv+yjqGZQUiWc1
Im8v9bMFmH0gWUy5CgwpzgdciTMS4LD2ecO0FhF6umHq84XOfufcySrsKK5/Co+d
rW//cGL7yTBitjiSWUbcmzaGMdf2EhkJMvc+6jJfd7HYq0kNPBUZyjSYF/qk765n
aOMKLYRT0qGr94Cua4+FYD4k8Aq61/dVUMnD+v8c0QzDX+A47Y6YMSWn25G+B1gY
A+fQFYSndSHZ1YUJbtMyWnjbnqVG97JDPkx8CmD5BB9d7hw7gjsRe/qxAp0DpeMX
/vrxCraqdapKy3Rl8lyzfzlRShlknRZk35Gv6DKHQLepU/OXfKJtcnqrrh2qv0rG
1+FaS3oOvep7BwqJiEOjDnuWXMGQu8cH3/dLTadZ+138mJ/puoFkD/RiWYoIHvjg
ZxLMlsf9jEtJbqR2HO3YzqZxOp5HouvomtSFtxsM5H7mUN+hCw6cG5vRrSftCgcn
ogfMH10bE8Y7BRvsd5ttQX4yByMZFmUPwKnSYnpFFORn8qO+c6i3VS5hCkHJGZqN
5rwNX5/Uat2YM21rfxkCIlaQvx6pazJ4dMRbRxmDh6Csj/5c6IOqe1WqAbgrAnuV
3do1uWJMDZD+Chm6hbwsk6jOP3My4z1tWs89ctT+YZk5nkwYLuIyYXgJt/F6rDNc
Cf0tEH1pAIOsFhz+1RaM5W9yWqiWDLCIk/aM6b4jYtp38LLornsE/0uoGotwIne3
XHe9wn+DsmKEuUxkOFsEvrT7IaRZalOz2Q2xQBAvg61LR7ETSJ7ptrYCGxNGJbm7
Tob4EPHrV6jdrffweFZo4/CUFeaQvnKeZ90viq6MvPzmtH3eYlbPu3yS2oFWnwBB
EFsxXnSR136JRXUXHveofToiTN0/+qxpOnZQKCeTLnbBp0a/AqjGj1nwat+03OX2
N0se7GyHtISecHiqcos94ZUBta/TWPn1ISorf8hfMFSln3qpoc0nCT5GjzVlOxJd
Iqw3r7Kp+5VFBvNUag6NoPsWiX3hkx0MS6/k6DuRm/o/84XHqFzTZ/kZ4y62RYD4
k8ro+QSaigrQhr7GVu5cDx7AyR0zdeYkEYSgG8sCDMWkv+6RMYzZpP43AKoWNMio
xD3d99iAolPkr35mlK/yVazDGtWOmqpD1zS8/mLf1ihwqAl2taw8LtwkL5PxENOH
JVX8mmlFM5UwtseDpAplpe8xGG5mAEHGzetxkq/7KahlZVkAIfTbIHNptL+w4AxP
uZDeLLZSeT22YEHWsT4X/J9MQDAQ2pqvCGZf2HSuqvIrXY76rtW4H3Biq4cbv8PS
ZCe3c1VAQ4aT8VLwFyirIjrgLOxHEWaxnP/lpaSLkR5qvdezlbflGC0y3uJGOgOO
E/ojTwO7x9bZfKOmMBk4SHH36j4Fj80Wj7sdO6hTGof2hVnpUxSGdmR9vrQ+qtWT
BrIA7WvDPVURcmuCfqtcsVZkPYnUx5hY4iBvqC5pdF7W2DVeQNaW1kFyuZ3Kn/Oz
M6Hyrtst+5hGm+pcEgUzpcQM/sGWuOa5rDBCvnTtrNDaFflKVWvr+0nGEcOA6luq
NMdqHP/Ic9HKxYXsIuh1NoX0UIpSVQMk8MeWbELcxgXvXBc+LqYqqPpwdk/pV0eq
guNIm9ZRPKha4vU+Sd2NdIEMpe/0XNzckuurScumCgEKdopyQzSkjXZYLzPiIrpA
0GE3wMXQS6w5/QGi1RZWN25cOkNrPq/fILveYGYI5bRnsArUuAqIAMu2IZ7/Zaot
dplwSkI/pIG3rNorNfKd1j7sYNI4/IbhSCRm7dsda++nLic8KM3EvkQiu7L5BvvG
+vWNm5smrI/KpuzW3Mzl0AzqW5xWZ74aCnCnovVMkwdf1hu0ltPpxGMxADzkb3a4
Z9klMvY/lncUHRVvr8ICXDzV9vNJsvFBtOkzaj96rCA9f5NwTLfJK7sQkmVzYBvs
QpaNw32ilI3nnqEuGHcftptoOE7qg060OUUgz6VYiQGlMH5QEzwuwUPPdCE2PKQw
1cyffm5T8zqdz0V7ahibJAjUgd0kruPEKyRtUzN+GlkKtwasnPvpRNOdwSOHA22p
K0GBRkdg7pEcj7TNmbPEd3mp/Prrbpp0xbojRYUBzFWzCL6HnynS/jqLEwzyeYbn
KCRkpsIN9soXm1eex1lTXp4B23GFxV2h/TmUe9LjQQqO7KOi5uVUY6MlQHTwXhLv
lxW5Y75cZL90tZkmt85HpgYPvxBYG/YioMijyLDyT2QlRjqomRqYPxAzU4Wcl2WY
IH72s4wPOGX/WlvvMCFyiokKWTi55NJ0mt09muoxSvln/XSIlyZsrs/LhN9ZBj2x
vOqhasFhAYzfC6xOaNicG86/nhRAtzlJF2JmqCtg+DSmYYIBXwl96iKnfOiWrDkl
SkEDY7rG73VFAVm2pz8XuQrkN6dcXSqp7SJ1o/XRoahetS9YaCACaz003kFrTXVh
gogQIIco/WC6imedMdHRASAG0aK4bA63+REoCHWv4vQh7BItgA6Ns0yzvm/pMCmU
NrqBjvyb38Gk+nCR5S/l60wlJ52J8mzle6t/ShEv3SyJ+nIEZbmYZQAKg45JHyQ3
wlZMaIlnpjzzKDK40beALBggcfILbkhTAzTZYwTgKbIZNET6Qg1xOyGPfwwQkdLT
YqIxKZ91P9wgiygPS5n9PtCBYZVSHEdRra89PXev02H83rj5gVh3CpYAzHQLCxjS
9ZQp+J4ritCcy26Wi41LR0XbmlrZQZKCOSEa/0d4L1E2fsXDXcqgxl1xPnIOBd7X
OHLqi9SjCLRvhmwQostCpyrmQ4UQXrWZBgPJAzoFASvjWLSVaQbXA/NC7N0q5aS5
40AkjxvtzhqbfkMBToVWUdBEX8dy4OPTbogxIRmMOgxq+rxmR3iCc2BFuziM1Ijg
fNWeAXQk9SUIRdu4PmxTYMzN5MdmNsoiWeOwX0R8Z/bvzjTKyJJYbOnLFSNc5KBg
PkVgsL9eWOpmilSxZyRAOyYa+Nl9v755UL3QDFyVEiV5yAW5KoMBxq4Z5L7lHXPW
IKEEVVn2REh7jBFewDR9OzlMe1Wq1rl56PszhoDdJGZj4bR2jJ5HD6/sR7sZvHwC
IPZF23EuTfffiIt+NZTAu7NneuIyCYcj9VnEPSgIpBg16ch1+VXvbIJ1qGLcIgnL
E0I8xFUdwvtb5pAkSZqctCJQVK6lCp3shzRq/cEpsoLqDpNadO4O7YEa17yEamG2
paoPn/rKdALpGonxPEbeCDMSaZK1yauSI0MyvhKqOWCz8+7gFCtYI48SiKbBwtDI
wXMujCzeYAkS4OLKOwrBU/LPPDAx6lO3pYjsHAi2xVdd8a7wuNeC07ksptsBU0Wa
Jx0hvnrWdjsopdc6TxI4Hxc75krEM6R49GDr8Ef/0zrc8ZW6yQQ3HYatYzQ5MPFH
ezFpHtDySxoh66Am+w6FaEqtPa1DogavmipYQo3BKmbvsvz3QpYxFWwZcVd9zl9u
GgGkBBQWfnwt7MPCR6tbeptegEevi4cKtQGTUK1KPa4heLFCv45ae5/GLz1oInCd
8ZPQuAA+3Xd/PMpBixout3OTKd7/ToMKVR+ZooogbQ+QspP2RfLEHppbhXOBEU6J
j0SK7EaoepLPSQBKB51tFWIYw2q842phPhqEjshqD/CP+DelcNJ1HKHPKWHbJI+9
huSpL4rUk2xMCNFj26SKvPokABdLY34DQszQ+3a+vlASI5yB17KxySxZSNHS9rvr
cLJLQLt2zE1W31GIEcsD8NF3aWK9ScAOfHAIca2om5Ym0O9CjAs+q5SqNqQv24Jr
59Ck/oydq/dfMBfu4zH13UFtoL49836/jS6ZZ6m/vKoiT9xRvIw6Lcx6IOvLcqmE
nEItvBbOGaMX331TuWc/CilQd5P5EULsxXlZxtS+7Sy45vzBUI4TuZuTXLlBOEMW
e+cJoxqjjA+Z70mE/0XVIfzTfBXkilGGh3JAjMBbpuYNKs0YDOVs0UEMTX5ISHna
+3BIPMbt3+YY75Zi2CMOEdV1RFzF/N8J5FEIwy3qwxxXGLIb3bWxPbvShs3zy9Ad
FIfkT4ilfeYWhJAmR9QPM7D/7qxGsOM3kYoH/mRQOdP2IXiYXx9cwdPcVQOkhyRV
JjfPgfem/yqymnp3PfeBjBayowo9+YS6dWe1vrn47huYngH4xURVB80TyeOGsXwi
D2U+6VIPh67KwNRqxLcy4l2MgwVsj6y9spkTesQdddBVdnJzlfV+C125S0R91E7M
d13GMmByWCi/QslldtrDS4IQAANzIWCf3yRUeXxVCLd+Ek/YyXqEcVnJTW1k+NX1
uxFd4cfCcngeLJ6mdQ3fY54S4hfwtmBgR53QYpN+IrDALqGoOwh9f9dhFzI5Ng5S
yA+IuU7pnKMQqsnXniDAEkeuu2AnnqCpsIXu4k0mP4OT72wrwWwLidzOjNx3gPQl
YUTpJgwM9j2BdQLWcXsjCd4wbxOsLxt2gOlzOUG6nmhnaWI1+94IsfqCtOY09riM
WjOb8FRW17rVMkeETQdELtaNvy9wsDvtOe3Pft0OVDeHgdfmgkISi2K5lqEqCtXL
lt2jOzlrHkS8/0sdG5WIcpAghUJjDM3FLX62bOCTRwt6/px7lVolBVk0pgAoBRUI
dmFKZNRdgW83jKtsbFoMSpvpH8cJKVKwEhiqJq/EDJt7X0E2Y9uBMWOu9VwXQP3z
8j+KXxE9e37FGf/kevOCh7ct0lut9Bjy/Qjr5AKQ+ndVuFT5jY97iyiKjro1fe/V
02TTo3HWTGSjKltxNy9ogQOkz7tT5P2a1d63MdAxtW7wXjo8JWE+zmZPVnKq1rjP
r1SOhzpmKb3LcskwQUS4ir/MOTkW/AYxCMVihoGA8e0mK7YhqQuUhsFLWMEUOFje
ugf58MptoLuBGWFNngS62fKpMfpkPC5NJlGQ6oXw0VOk4cexdePOBjkYEBf00Z+3
7KNwekYwSvAgPGSGHuFksciwWFD4N8pMoAVmGRBmLiY/n/i36fCqU6a7PlrJk8yI
MfTxeCIwV812Bt8ks5XlrrniRx1/Zbr5bj2ENOyARmrIu0ammxK72krL63sKGaio
IBB90YTpAd25uhlDPBX5M74o/vRfsHiV0EhKgCFXUkbWmOYVzIlFY8mJtXzBdekL
YpIsKkgaOcdTq6ZMTzdz+T9jjGfh7TnpZFHLAAnGjBDWTueAGll8BBATV3RjGX7Z
XaLz55OqbihbaR5fAorEuSWJHdolW9xpM+VGtOR3o0qByodHx6/s4omJ5s3IgxBj
zAEQhyWjJy4piAsTDx8jTbqsPtruZrKpjpzVAO0rkgECBGMBKBOw/RZebXWJFPbI
x0nMa5ru1L3jD345WAZ1ReJ9TPwT0QCpKnXKuABwBf2vnFsDkmwbE8+n2vO7Sk2M
Cqv0JX5Tk8owuhD2zxwidvD6NtHlDgSge9z8VHdN8Oz4OJ1pFKEMeL9WiDR21AJZ
eVCoz6vmC//R8kyl4zKsg3cD5OStR6qm/2+I4iqpRhuJybcHr3D6a9P24oHYlbR1
520fHootxJkCqqzPJvtjCw1bcDBpqoPdEbLnGKjng+B/oHj1yNm3IxSlgv8Cv+Dj
x7yIhCAncyU0y8y45V/qe8rt3Nhs67qHz8wj6j9frWG1JYtqDWYzl2cF0A+JmrV3
Ffq23lg8BTYGIIunvTq3EwFqHJuqTMMYrrcgUqXwXDTu+DccHs5Bq1uG6fELiSIF
XKtZk9R4ejp6Qr87nPpkFMQTFn3JmE0fd/ON6EWQiAOtjrD50t+D3OAVSy3Efcle
s0dtgJFpcgHmk9Lnlp/6VTylTUu3mHVqAmM1zt6ZFjwOamPM2VW0d2RRL8uGn+UR
pied3dZ+taLXMTsiWTL8tYM0gqJ/rZbpMD2cqmVJLg9AaSn4QpTR/PL0OY5omMl2
QPrPixAJwlV5+6ifpCJ03dVHt4Dg5uHggnrxs9qeJMg0z1vgToKACrzd3nd0f4ao
6F3EVd52N/4wWAVZyH+25WceYpycJ/wHKP0bNLr/sXWXgRGi7I4CwXopxW2VP+2Y
8cVgkDNx8EulGl8U8nnWPvryRruAEDqYKxbprN9nz2+C9/vEO3ty06+nZMkMPFs/
FpTNzShQ5y0H8V2gHyp0BDpXgM/9fJhh4XO/JgH4MHIIFV5D1P5GQIz79q493Ada
ALo795+tfPTkLzKlAyupTjHaqvs+O95WVu0i+UX6W4VAXwCSZOgHc1R3Jw8q670i
MO3QWkA3JyCP31sEiyKzyG8gACWu/pg95ft++zlaDR+fPrDG7+a/WNSZkmgDZOaI
vo3DvykSSphHBPUafhEzfPku292qdqzcHi53UQYYkDxqA86V8q3bhsXAdvbNH1Y7
1ZPf6LUTdpDaj2NGJLbUIpN9bNbBfO+bB1Fo6f4Zk6t0hndaKD0UGDyzBFDquu2h
2mNe+ElwxyBF1rEPWx9ykmTOEh9g54sjh3v14U8nSBgtWQngWdmBIkqj25yQBVhW
EcFfx5FSl8NmZxa6kSPZy5BhW0xDjsquPug19shHvCw0gpP66cIcZ/ZqtgPaNH78
3GAJ+zPXP0D7SqkBL51klemrdDPSs1LJX4OtwiRT10qV3jIcEcGSQUICQCbjn10H
he0c3Je8CKll/lu/2k6e58tSTRG9Lg+x8a0X2/59VGyi8yVU/T3bsxG7EDnw/x8V
cF5SPTDZlTuL8+pP5eOobcAUz5v+LSu8zpYPG1ehxA06rfydgwZaxZhg2EFFJQ1H
E0GE/0zN9/Dn5zx1NFlhNfz268B/YmHXOLUl30kzZUb0NwAnOt200z+Bh4/uqCUM
TQow5wbB82uuevp7yRhPbqp5rUjgGIz3Q3o7x84rOFm0zhtuuwvV5TzCl2OOI0Mr
TZDitjWZI/MS4Tn5mTMd+hyBZZSNTnnt6UqmzczSAxyWj8i5/zqt7Lym8DiHqmFt
Dthe6haIMDV390V2T+Yai9uUBok2n5h4xTMFZpSDw9zhTug79FWhVDkfmTCTELUX
PP806FvCu/VPjb0da8F7v24wdFo31Rv04F+5mT0iwq4sY59XECjCOyVAYqRkfqec
3FdvQUjP+v09Gn016mfdMa0eflRiwG+fQN6CJ1yWpKU17lQt76JeOeEQ0Ju0axTg
icB/xORn3fjOjpEDsAbXJVHvMKX6RdCmZfh+fY9pKpbfMVnvxcEfrM4ZKSUo61WI
/v6uvEX9TyrMw5/HODwKF+QY/x77vWxsATKg8le/lKbb1+rL8h9f0aYO+t8K8SCY
2ZV3UVAvKsJL58FGCjJAEs9/1JfF+Pc3C7p1FoTFeBiN1qvr0Q2e/SWhpiLl5g92
i3TpqCvsMR+3saodyMziwLbSzqNPhzhqRNPrngYt6qaxvoYtwdRjIueqWYDPBcgL
F8MOsXJpynYcvuPu25/trF8q6ZDl7tVtLrALts0TJmhwEJBQjLggUmcK3iUJe134
iL1LqAFUaZATqUicUjk77FpLWg6XSGiyxJiD3h4V1RSmjhmkRWyW/HIKzOn6cm6b
QsP3cCprJeyPW/MJ0jsi6S9/+KdoCakaL6hfeJxXoAXgjCAhr7wTEFu6PokiyP4G
gnJlbiQVplUTliXks1DcFs1MGhPzSDJ/1cysBRzB2lEAk4BJ7J7eSQAiWXMVpPLh
Yy1i51sX3dOhwXE1YfwY7mmDM/3bC6iskwAyCWaAfdxc0Ves4VqZeJkt45Cqu0g7
IYTWrsAL8BS0XJBsH+J6I/RAO5YTUcPLGN7iY8BL3Wd2F4UbG8ufyiTlnS7JhlnH
+4Tg/Xw8XBTKl6FzxalCzX5vo2FEzq7WO9glXcnXN6u1F2OXLzKWPGScrO9SmwUP
f2+urXR2uXlv0HrHy5FnRSeDk5HiHZElg6J9qig7QhnddSLN0DXDKPD+3yTOq3Ua
+cBQJ8Kv3KQsNrN7CmKVHBQJh9D2/Q1Of/5TLccy4rkr65Uyax/Gf39KvNEnqtnD
SHAAVPMWvYlgShg9o1JcYDkZprGdppkyFZFoU8MpgVecN2i62ZonhDyV/lfhMgyg
qekszw/F1k2FK87N6sFW3BJWjhCvb15GtdF6qdGfxrGMdgLS+20S/2VYFBdhANKY
6fZejSLUeJsr0w0VXWPUK96RhI6exU7WWMr9HA47927wZkA7syu9ihjIkdytaDhr
VmaCyy28wKJkx3FfEUGkkUj9VpyWtxfBPg5LWs45+OZdAZInjTviwYo4aB24eZI3
Ii1x/UowbYjbENb9m2eCN7RFOFvk2GR7KEqZw2JTIAxxPUNz2oxETunHEF4CeXdD
TjCK4XhGediGMTAI/5whhvMwPYluRU99rNxZtd8fFXNi0EI6HW66dHzYxP+EkHYd
oSMLlQ5DBp8c8ivtce96sI3H2dpEuStwaW447v42n+iLgV2G+qzTQzStpMppscIk
PAP6ZKmvVErFM0NTRpqncDBSWg4Yk70jJdEWuIWeTDYs8J5uLC8FQmJBRYvidriB
YKEAceL2KyBHhIJgjEkdQOw436+F8Kqe0Wn8K68mge+2YBdGYF+DpaLtxRUzks65
ogVv88t4zciNyMoSCfsPYc5DOC/LonSQof3xPmpBOhs+t0GC1FbwmPj0D8Jj1XoH
i4+mC+bm6Uolfgj7tFhmslvSgucI4kVAPSiMG8J1xs5naZyfu189eKEN3sAkTW+O
4wUwvz9fbEKKQNSbQClXVhpeNt7kTyahLjD6b1gI7hmV96nEWiZZliZ1wlIJY2SN
JU5JovPfIGs6nd9zc4AnBQS7ACITjEn9WqUdSGa0ehprYX7VvhXfFpSabJ7nZyfs
mtBWHgSxxQo4voIvuPmSIxTL+phwVeuzlllTYc+ARA0Ok7j6+s4hLi6zMnhmc7ji
jTqBXepaeU9FmD+y/fIzk3Y904EcF5SSiaXS3rMuTa8tkev+2OnS8zqgVbo5Kif3
uVYVjt/QPwLmj4JJpyV10PLLGEluKWFYcD8BkAWYx2k7vVQauGF2CLbiZprkffjJ
opk67tUpZPRdYWVc+dXdqjUqlyEDN7gcio8Cc9lVQC9eQ8+MajH+ew2EJMdy5Kgg
dxkXYmUuK0/wZhV2EjkPyWh0Q6KSCNzJqLx4wpCKGe18zmNeFvgSW6VBtkrapR73
hv+1CTREA3RUia6AO+5gl0xn0prME5UuCghTbIUNnNV/UJtXiIWEbGo1Rs8Fk0SM
gS0la0n7F5t1QeqqLhzTfeVNTcRHtIzj9MUVW4vNBO6iSjdwHMIb63vSsb1UbU3g
uWXxbBwT5hzkRgjuRaHjTDFnDmFxNm05elSW4pSnEIJRrx/fMq3cfzyUEkxvNgoD
gw2S1qSomJFq7QQxvelpfu/bEDaf0QGsEOkIazuH3T0SASPkZg2IjWO4s9G+SgLE
QoXTXpaJh0JE4+6bDm7zp/BbzHMtFS44uuyjghgrmtsTajKV7o0yXjG38rTgfz0g
0j69sZkrW9Mybo7GoUjPNPuOASlfLaF63oqCe4BuAOgTY+wLqk6/BkO/sdSmL+5v
+vYi0CLO9Wevv5A5OhULUb1VA0iiBYpsY1BheUsVZrWFMUiEsjG3WjQdioEmaAr+
lXzU1D8yCqbJvR8Jv9dQSoZSZf/05lrPuL9pwlRcu9QS9KhyXl61Kz0FsydvBlOR
Ej+KiOnLKveo3OtW9nhhwAhxUbAuI5O4K9ijBZ63pyHleKwy/hj/aya7fqrCnA8a
sMOX8f4pWLEuFdBQlLRCvWO50IHzlodyFHtDNT/uiQxgX0tjaJxUHQUW8Ab3kOBM
72K6faHeVroEsCoCZfEZPxezjbS+BeU/L/njL+b9rX3Rt+D9FLuNTG3NMEAskuyL
aPw21fy9RsSxCbIvI/gbZOQBO+PDU/519PFpFyqChq06WrL9VlFE/HWoZfMNRakW
kHMi/P2mcRsbEA7fixiv3WwaJle7+W+vvJuQLBemt90EQaDHR7ejfdXM4abcvFOQ
F2SyMWo72jPgYhbebNHdrSgfgR2qjHgQ5Sx30zCSD2yELcGoAbO1c8Y7pd30YprE
agYBL+MRbAftUNck9d+nAJgSS5fukvQfNfW6cqKI6aVqsDxJNcyPo2r7pz6ob0Um
qcNyHjsw+em3Sv53LuVDd6t5hdbb+xrkepdRz09ix765OJ41lPiqFstgPOADTgbc
GFkXiX06UexfiDk4zUxubk463doMlBvFW6cTYKmqaC4+Y+ESpo+IP8lGJ+3ZVgoy
Vudis/OqMfdkbl6VpjM4bh5FyCqw3nOnu03TYqHLVWp5NwwMx4llTZcZzKKAzc0O
e1ppJoYzQ0pQd3/gIO28T522Z+CMZyTb7WtmsdXYNSosqGS8yxbtzod7oWGb4EXf
telWQ6o06svx9QIkGNtvbWZog6iJq0MRFrE/nOiR9D/ePacuop87M0N1YfFdiNOW
MhQhCdJXbOv9thqc92eTcl/Ee2GvBXBzh5gkA985z5EN9S6m947QCzrI9vA3gum8
ltwcNi22KERq2a2HezxBJkUDWcrRjeWF9FvPxMsr2nidC0IEcNDNBozclI/ZCVmI
51Bv00wuzacDvrVUn3yTwnZMBuTnl0LiVUkfvw53RwYLmGMcw0mk+i4aBG0t8hPt
EpeOLNBcLM2QhVguBHvMCfldk3UfoJNw7Ge9IHn9rE9YULI70BwO5ZcFXqwz5qwZ
+xQ8Nu9PaVoN5+nYwKigSRvs7Z1tUmWG8ymeCdBfFPCDnZRXwAIT0SNJ6uIboAu2
MYDhwJhbGd5PmavIik7OZqRKOmmb9cCcLn9Klz+zsBpsOzV88UXTEWMv3wQggJYZ
CyokiT2snqDMDAMNR1dBhDM59CkrVjWkgj9MoWEWhTj/6spCloahSS4MEAXesUqn
zG+wDXrFTGmMTCzPw84JqWmREmQwh5sutslwqbc/tX+VJEFYna9zys3shXNrnCpx
pbqbzGtJatEv3mOElivicmuWhiLQGQdOyLX3PZyRSdin7knLwghnQXuIhvimeTOl
wcubXwD6+HF0p8iBrm9Co7oEPR0rBE3lpwDUHW3ufp5lopcGij0rLXnxnI7vJMns
py6zYh2gopThSyjI0dpHeEOI1ujPc3obzCMTgw8S8voTEhfuZ6sKwqglpX5q1GIS
kNxpKj1+AVKadqN0TI7SrAlWwm+qCC1C5Q5KdA7roGoWtjzxxCa1qpTPYUTBHi7L
b43As+HwwGZZTd+zt5MrCy2N5+/lUs5rZTrUMyv/FH8hQR3SYnIaIRrpfSkiIiO0
HgmLaiUiO8rvcxn+N2Nqya3v3QQLwfL8NoogJE9yzFoS/VH2DGoNPYIHoHdIzh+Y
5xp9+TIQkYi7FBdT9vuqcsNvN7kJgPMjctw5g0E9uhSVed79NFkogBViK0p0hQSZ
zw//jHnsL8pZ8C0AwiPs+wcD4NHPFF52NnUuMgYXZbpOXuu6mwAPDei5ViHwUJYP
7vmsv5zIchKXmCl9hn4hmzerQYq/CD6/IpfCm3ODAznYIvDpS5UM8ZzRA+PeKSXI
wYG5cNyshjR28D16yUnIYtt9C53z6HJ2pEmq7PKZOJLOdXIM0LCmC801F0AORxaU
GS41RdPuOqQq7uP/lA2THmOFhuYyUq8E3wjWWYz9AEAcudgGw7CEwXF7hVmrq+St
NDNM5AnrxZ5n3wQmLqBjahKYeSYF0XjTz6P112KfuhR5wGuSaPEyf0Bah67afcKD
EeaMwuFxvwpuKQ7uDngtbpENP32R1tI9P3X2TtkMwLHyLpD9kolYp+N55qFSidNz
hLe1TysxoE1u56Wd9xEJlOvsxV4w8tDccqXHlAPBIajgFQl1TY6Y2hjfCE940KFj
JNXaZXL6eDN/uoolmD4sIpN+OuW6RJBan53wOgeptWobiXrV2XyU8idsSmyQp5vM
6CdGOCxg0ZpexfotPWg7JV6aF1v+/kIwjbUr3WxpdfpP3/a+JzYTSMqxcdg6MPI2
TrVUEc14L2OkTjPAQgey0MwIjV/q4mg5hmnSq/QBd6c1DkdCwmZ0AyMMMnInfujE
pdU0m346jpebXkiF3Vs/N7njgCMpJmA8TuM+RMBmuZePE62AcR+9Kaj93xER7ODe
YHxNMRU/zDv7AYoDeIAPq0euIXn6caLfg/CAie6Ev8+uLXTUqVoIpzFtnyNX7nne
sd7aKwlhwCgI8ShmKvrzKM9ZOUxi2IxkJT/PNNM97xx4FjMaCpOylsTo6/jMBnA7
T90s6BiLZqaOoPm5dp2lpbkRt4CJV5p4pUvZO7UM7Sb9XyinfYIQPQQnLMa/7Z4j
yn+xaqkm4QKI/OfSh9Ydl78SBNVvyGtNKWhWp/uePajaLNb9001/Cvz1wo/i0fZb
G/NKNgQkDfq2nHsa9YYcOhXBoiO9PFvwQTDHMYXLYl/9dPUbiXEVjdpBG9O1bci7
L22wTy7rLrDw/bARlztyCJ0j89GuaeVUfbhWJmpgTu+JwauTZtgA8NtK8XaWOBLp
YeqdYW3lqCay/wZtIfZcoirLBmMhWWejzM3VJ1tij2iJ9NYS+mQ6nng/iwVIrhol
U5l4HH0FsKm+C5sqI/TAoaN2I3hcBhi1/S5t+GwCmbYk9fHkLkTaAaY9q91A+P0V
0Y45ro65bfu4lCVgjTMHzIvXVYLvR2W7+fLRu9qsxj5hmHNFQR6KJEZqzJvIGlSO
isdr95sIzULHgoms0cKopvvsdMl70tatJH4GJxWrmbVfbPG6G7Dalz+POQ/brAae
5HwozcYH4K/SwamHmVS7nOk77oyVhhjvx5gb2O/MC0QyXb8L7j9MFnezKS1dNSRR
qAaBUC177p/0Kt1gAF0k7CSZlH18c0nB3Ey1CF8XP3aoWjanS/WpiPyFAKFZP/fz
x27llDB/z/3PWJeSVfRkWCpZ0rGs6l5u7AOB5PKLqA1PA+ZCdjS312e+jJbEbW7V
vnAealhxhNV8NqeJqSgxOODk6llQgKPX5wDfBXTYzV7k8ZRXy57pOdFP1GupHXv0
h2cevHPnlAua1i+ivyoBgFIhpjq6xTzADaTJlXxdfBjxlkuIsDjgkalrWc7wqM0d
lrbOEB/97quVVQJe8bRV4Utm0Cw19Q/0l1TMn6W+Y1SbnYyUo+/mCWoY7HdkV9uf
q6uvmXlm/lMdABr5b5QpUg4gBLCFbbtp+qAlLhbBkO5TWzHOQgUbFWmdN3fXLF4X
m+3RDss7f3Yk5TXaFZuEqKPwC43kx0y9q2QeXha5oWzYSYrBBY3/477RCLH6PedS
MB4wqN2Kz/LG6ZbFvEI4Ja922aq42Gn/GD/lzDHxOVOhVlqPAjsC5FBxMucbSO71
1/YBaw+PqBpGtJEmzE0w6IPBaESJW13oUqqZW2gT38tmkJqxAHnmIwAU9Vh2g0kH
5JBPuGRnbxBHjwRhPV8HBvRABt65v8FslxEN25oOANtSTo+TTXefuHLMlFFwBEXf
gllW18SY2SNj2JR38/KL3nbZwTYEOMg+m63g8hLmzNMy3wjcYkzh8xd26FuL+nt6
Cb70BNULwOuWeeV40PZrohXRrWURwCHWckZAMXyajj0xjiK0BJh4iBlMgSM0TjtX
Uw2+M4xp0PMBsCnHGXXvmgJsVmasd3ywciV4CbK0paRMMWMWkG8jkEbOAzldsw70
tbzswLINXkaVIbYBIBCA+9PTVljd4ztbPBTJEA05bkYS8QWKnS3HXCV2B/gjwbPm
SRJTF3lrY7+RxaO6adMMVWDPHbHdgSJTwXar1ux6EudFYu7zoPIVBZwptZBssBQP
myM0HDw/rRhXqcEuHdRqnBfPSk0Q1pCBZW05eb19fb+knHIL+27E/3fvw7xlOaNM
chOMr9lFh2e/PkObvGWe/j5K6s3fUtzBEzOBysVetrNFclxVeZlA18/MwkL+0AW6
VTfhKgquE0vc8mTaBo1v654zybV2g09TV01pSUFBK2DD+dFKH/DTiDT8VtrCOMKA
lySH1CS8pUuN9wRJnoMoOJigKHtoGQg359cjYgrFWnOEFQcwswaZ9Bc7ILhVEdtb
YrOPrGDywNEL+GSkskrlaHtSBEWIolIM0L18gsyTxJ0HWbExQ/gsEj+VAomzpNNT
d6NCC82ePG1SNsziZQee+JN+/dI1o4T4QVGoAo1Lfj1v1hiygQrGfdYk1VpQry2m
4CPyRoyChBAqyaM+Mh2630uLt1jZRmt8I+2nOCu4u/qhT2rzX4/atWUGl5ASGrI6
oOwDZv5CQDov6YZFILjxup7/Fb42NesIHASRqXV7avRyBuUtNMBzI0gXU5KxynH5
6g1KJT7ENaQo8ClaAbIfsJAMsC1UkJqdFYFu5yYQq9aSQuZ7v/wv0XdmBP68/Lpf
Zy9MXyCTq9DFCMjCrjLeNQwtLVk0m3lwwtwkAeDNEGpjwbxA/HTPAzpzPsGVM5NZ
BX5/DcmbMT4yMxfrkjmtTPQ194KisKH7Qlcp3soiHF81nOr4yvSPfQzGa77IOfCP
BIpY/SHEn9vI3KyQea4HSo45UAgbAR47/Jyw+N+IATuvdEc5QLP8aS+aCLEWyaW1
pYpGt1seXeAzMFydAjU+TNIvv8nSAtLQMjVy1AsI1PBXEbpbtJWoDKJFIvYEzB4/
lnZ8KVRhw984MhX+VzpUmP+LbnMMLEIz+bPTcz2Je4DkrpG+wA1ji8ax1YQAwLim
1kG57ITo8e/vtNMCMxYYgY1iHezXuSj8e9yxopdx25n6/DiR0eLSMgyJkbQYJvoH
iJj8h3vMTN0/5wWsCA5e1OQgLOh8trG0b32DOqoD+ijvcUqGsHeBu/7J6Kql4Jhq
+28VVOKxzzzyNyi6WxXexhb4OCHVgvS6Wm5dGuQDsLdGXc1HotLS/vTu/Wi9t2PP
O8g/0U+/XugGZTGqv7ZKNjLI5tBoq5vDOyBt705227iBaLKjJRAxbUdsSJHloyFK
asYmnygjEBjimXBzDv4snfqtLiQJ1ni5X+cCbx/3xnr6rmWmOXMVfa+tKyMKUXPy
qTnw3LjsW+3OdqN9zabwcd2IebRGtPwwSnUYSoNBcgtWJQeUxBb6KUYDWcolmPNI
5hyJdzVyrT37PdT8Sukq3UEA8C7FdzYxUuzIy5dH7/cgZuc5bT0cvB/J6s9s6GSn
/gqftfWmbEFVNlmrF35N8eGPL+ddi2f3HpFYsGJyZRuv5Axq0BytwsbJdNYRryIW
2j+glU+lN0WGKMn5XimtZX0INsRrRTnwNLw6QbJoLCRZQvrc7fe/ZCRz8q7IdeGJ
sgh9XF8nLHszpNHZ5LogYCRb6VQAiiI7QkLoKEx4oepJtXj0eZ3DT4QFVT9v0wnN
64JLvl4lDjBUV9XJrg9PLn3UZIGYw9byDqvKnCaJB+5LJMxEXvhAxN+7EMxlpXuH
cUtJWX19Lt7o5oY3gsNhO5XQVR8v2HpA3SjfN7mT5ZrZdZAGnxOs70J3bb25gooy
ZBKrQG4J/V42MRISYYPCMxWIZOgKMcUBXdR2pdcAqrQ8P2YLWaT8GkoCRtGYQFaj
fGKgENdflSMZT6zOhI3WT0EE0QMs8Y762q0WFATiTLywau0CIl0/A5/TdX+UIO8Y
hR+0DWUOpTRykthYEpnlxjhV1z9WOj9AL6Pb3boVdnGOPH5+hj3hpeEAbC0KHm9A
JlHnf02z194r1EwcofT2cwu2ztM0Mf7SFqF7Fq2qd9iWW+dmEdqXjuO84gLq2pCR
nUUl6PUGCHFCQh3pPUv4OeKTXbhWQLTfP3+L1p1oLffzoGUNiv8OtE98lMREo6VY
2RYGsL5v4FFjajulXMy1G/awkiyfuWARSLifUg41l7PrX0HSFYT4eEGsKVADae98
iS5OF+OHHAyk1sQ/3AsgDaasKAp9TbPpHu4U9A5St7erlVW2xVm3wFDZrhqrEmX5
mSwJElafxIwlybSPsXz18q6wwSh1brqAHe9m/sKvviasd4YRQbHMrCi+1L44hW0Y
jHW2/R7Q/jHGs8B0K+khUBgdeLCCQbpqB5R2d8jaaeukx34V+J/mBv27hMCUDM+/
24n5fTF9Du4SNXbKEw+zjsCLkP4bnuJi9IoxbcH3/uef19Fjrk0EcwVMOiGeO6am
xRaiAJSk0Fl3jux+YO3ftvflQ4GyBtdp60hJ7B+e4RfLhomukxEXI7PhR7x25Cpz
i4lgXoB3I5GbVXMDwpwkpBh1FDRpylGc2XYvqAnKbcEEj52J37HQNKthyor5sYkz
MMdTHvc2mVGHyEM/caE49b9BYP1fvXpqmG5mcTR8DbzCZvlR0dfA3lyir32catSR
8G/5swauieF0FhgSLpwviPRG97kzVnFvBrutexNMW2IXowVNm1iZaAKvdOe6Cy27
404JyJj0u91Vaxa1MnuUrro/TPuxMM16fQNXys1q34HSYtVBm6ytCfAec+epGIyJ
p25mKWpvHoiRC+tbD0pxv4T2qIAcU94rzpNqYyresAmm9Kgoe3PvEQ6oqX8mKix/
N+BdV7TMjc3N9rSYoT52BYTlWNwZIo+Y9HCQOJEOzorpPM3y4TVFULSMn8Gx6OEC
RvyoiwC7sxEz1Ow9cpBeprICv1Auvpdu2YhidD8PAxbg1+vHamZgkxS0qvzbmb1H
UPkw3FCfDJLhf4oKroQNhiuR/L89Z1Z4BlawgzwS76ZsWOz6CWr6Ys/+5oEZHpVW
HDGq57TTBmA6p0wuu7xeGIypVj11cOx2Q2BhqJRjBojDHpjnFAH/prRsJmZXfxmb
kSGYY8IveXb32bxAqPglYHkA+bvmDDLHwoecP2ZZHAOA3NSxM0xzupufWNX1CoxA
/ImK/URsEMLjsW0vDnbOI+aq7HK9K0vj0wvmgl0KRDEIEDPABDN4QzXyiP9ou0lL
AtDtFIt7z3t24S7f8iVU1qCWy7i1UVjbU1iBp/l+WjxrlLb0j2Vv6nt27BVAUM75
LRTW2I4k7qGibRdM6ibUoFw9Cl8oH9Qs6P08R75mlTNq4l4bAD/+QbASDlS+OQsX
2ZtDzKF5Q/v9iOIG2TUC7PU71HB6RfjcQPAhe9mkQ+ytlkE7xWo3aL24fkMHQQLM
Xaud+vj1AwtTBpaX+dkQBc1tXypE5X7C02Kw7dxOtz4l5B5v/Yd9ki0oBb3EEo/3
QI28028oPx04JS5J5MhHWBJeOfirvV3qLyE7v46QHFAHfIg8B49Z0rVEFkW4huVs
u0RYAqVHGfzQM1Cu/tmc5UtRLxS0nSWQ1PA2kjWZblYxs6zgL9AW0TnxVO2s3RhO
LNskUFLGf2C5HMHMailjnvOUmR56vRYJ0le+sFU++InvB3oG9SHOle5OcLHnMTsM
mHeuwyM/R9PCjGQy8HXrK7TOLLjLY/kNXIsaPRJzxBX0BCQNMFjyL/rM/lzpbaIW
6aEwh/1tYet/70VUXrmTsUAhStqHE9/MjtH2uPCaSpsI+XMedraNaoNWlgMUD/8w
k4chW6TToKJjGt/OFn6nQw0yEAeimOLU6HUzFdGv4qHJiVq/1yiRAZaA3g5+Wiu9
Y5V8Pt3X6RE5pQcyHEl+NNR1Mkh+TddXrL4bB053eCVJYTJ70dtqpsoofi/p0OEw
exPpftCUmblLigNE9eafay3dTBHTgZAnwtQRyKFKN6+gGu8i7QkmQpr3zEUNyP8j
O13NadYZ+MMqROiwRllBOLMHgRt8OWMwAz9EgWNm8nBs8xwQh9BTHNjCbpgSJA46
K3Ptnq0lyEW3x/7MoBQPLJ/JGEdzL8tIXjWC/WyFd4XhRTtyv4e970rCQJj3zUgH
Bg1A8cUOl5wgQ0zbvCwobNcfOyJZX5ll1N1DE1OmkkC9qBAjepVwAfl5QsDjVrwf
7NRZO4ngZ9y02bhra9wgZ0ALt+nAR2osFQ/mwH5EloLow8bUONf7tf/VTbGQ+CAP
7lgaq/Iw1NBBppjz9Ooed/6mUfPoRp3b7nmVaiiQYvdz8t5rvOLaXwFxqy2ooDLw
7XTNOW7xxiXggQcQo6ibVRu750ESbFHjeFJCUY/bkNWv4KKkRhNdpvADAI/4ADlh
Sl6LzizR9LugE1QqN396wvrqtxWit8V+CV41qjKcZtypYwtrXb6MQSQJwiGn7x90
lqXYHU7y7YlHldBYHt+K7dmDZp0Rvn609+cLwwTPmOoXAGMNxXB5k3w5wP8bzvrL
uCRBNOFs8VzIdkl+CMGZiGc5f1zSEovHHSDlzt1fRJDlXQ4PB5HSTbkic4x+omtf
t8IyUNHUoATJoB/37LcWlAH3y7PPBwMRsHMDR56iAtuOzBb9a0SNak/XDqFlXmXR
4N9yhemlvr8pqCwu99r37t27CB34VE+bfppM2p9XB2uPVnEjXCYPaF9Pigd6KMFU
WaPijl57LDpwOW7Zeo9CYrVzRB6SLsbHmywnnUFCDLXVvHDVCstHU/sFVGn2yGND
W5vjiaTCvlktFic/INcz9NtBy6f3NIBD/4ZH1sp8tq0ybH2GM8J0Q+5RfUJvgvWu
DfJx23dhgFcspnUFaF9ponUu8Y5sjSo+eznxYwBDmpm0kcAF4pJ0nKJRjdoKQK8f
qt0GFF8g7SbM9QpL+ZitaCgeB2fH602WQj4WEeJ9uSlgx+LJaTYPFQDbEfXGIjao
hrF66yygmhd1jOU9dHQryq9ptXD5QIwFTw9xf28exBFhfNLTYzB/IKm5SS5u3bBc
EBcr5Rd6QBSF2KXKSFQu8aMggB9BblY/gP+kdT3leXhKTLKaakIf1oKUeGl/Ciye
CdD17ruviKKltzGLp+249cDYiVzHDo3dwE6RwG6exPwCLZXi4qGlMtCje42F1OTg
UvzKq+xAjgrbGr/lyOZPWQ6oMqBwdmrGJf8IX2Jra+SmVBjFUXUyfhq4NY9xL6+5
Q/izW8O1WzC5DLxWQ+zswcK3TK/KuGnpDn5un4qqjQstMw4aucxaAKJ3btMeF1pY
Xo3KdrsVzV+iGpWzQbMoH78T0EJ84W0CRHNF1edjK5qdsDRXuLUv8jUIRSzYqmCV
wpTFwRKF1fYCNgCCWKlML/fTIqHK38crriIwokRvlF/JVkAdZ/3QFg5awdieQNcA
q9UapLyjE2ChK1UfQrV2613myu/nQGkwvPHDOfpuLIZDrnjIcbUpsWmHgqgYWkb+
im7f+wD44CrxYmAqQo2qia2TrCeuOPvhZNyImuudN42ZzOikfbX6kIcKzS3qvBSt
AbfKACFuUHCP9sCmJi9haEU9IG2PEctZLO42U3FuBYx6eTTQLIsTpYGjFlSk01dS
RxHjODaSbpNt6Q0oCKDH6qAdc/6q5WXHIZQfnX1s9nujzp5sipQ7JRJKO5Rt0Ky4
UDd8KO9HxKI4KmrgdxCTmgVlrB2NsQtTP5Sb3ro84nPmBOgbNnPEtsEtNmCU1xsV
C6RJTAZmEO89/zuSXmsrLEkjmdypwcQo3VN5TYIW7ZEVaZ2schTb3jvaZgLltpIB
DFaDiwemkSyYCdQT6hiKs0zUElHU/2Sf5Dp2PNy+hEwQUy46CBrThu6OgJOLszaZ
xj6/CUn4cG7qVOQxRODWeWnZUc5W4P/7hC5FQRVfbh/AJI4RaSJmtvqI908hVIWz
91QbERP+YO+kv2ydIn2UUT0ZzMzKF4zq+XthNiesTrLkdFTnGhrRE5IG9bmNTeP9
PmtZ3f7wKnXPjlETbYjx5SYqCFM/GIEIkdK67RqSOCMHg0OQVriEHJQwd6VFd5+a
V9P7UeK1DE/hLZqQ5lRavyrj+Tqste8aQdInaJmFMWCfB8aHX0xlipB6DePO31V+
Um058XcCkfzCvkq+UecMcMLmOnotw8VzxFV1jlHhPSzDG6X0ByC5YjmTmlbaGdgU
AnEqId8e2zVaZ03rFsJ0m+Vc0NsK1Z/Zn95whxrci0tMPHIIn9SsODkp1Lr2n2oR
J9gwWpK3ppkWdzipSWEyQJRDqWdK0HteicR75Na3mMjN2e3kjExFe7hUgWF85Y3P
phFUT6JKPjD9t+ow1nj3gVpgKJxNPDwZJT9fHundiyWjSjl6rYMazZj4OPfPzr54
Nyv/P0JyJVkL9P7zu6b6cQ/nD5PUjmD3jYND8wedHjgDSQMn3u+IHAQaT6wnH6ld
7xlIpf3XIseOovR0b0hyG42EDnZB9uEccktQVena9XzYR8vQK5Wcv/8HbEWh7yQN
2+GE+3GXoC5QRmkGdnc+fJqCVr1uNRyz1QCmclMGHCRPhRYon42+Mm8vxe7YFyTx
cXcMXqy1e60hBDujEaj3y/kZqzEPo9XVd4fPYNl6sMSerr7h0Y0SAItOzDp4Y74C
PgSLZmgMrVCf/61eO79AFhtySZcAuRBJiRB/lJaqfOb6FJwOV6b0XG1nFmmuF04P
KfSvjyC+OokUZrsxUlDRcnm8Obq6N0aisd/09DxfF83hrTrCW5JyftZpZ98yXGsn
CmjWzeeOJNCtyvEh7pmLiWrso8xk+5YgllI3bboe3/MFO0Od/tqe48C/GX5SZcMw
4d3am/iaP3ufxlw7xDCgOSyvk5BCkf1ItyWZ49hvshodj4ZNGANV3IH9K9aQis2F
KGWUM1IYseFAmDkSNQCbDACsye/v/aFTfu33cAPrD10uTGRaCtGupsQiH5Qj14KY
p88JUSUzNzv4uCvnTnSoXHRb4KoMmG6V6OAlToK7jwOKCoDmFA1zjkVmdKF4qiPD
9cxL7kQ8vTUNhWZKdJHdjSgpp3XLPXR4B7xxD/5yToMrMlsaVF4lxvmwr382SNi1
GSKzBMCkq8ulAH1dPxjJsTphqkQJnKYL7tMr3SpM5Ru9NmtRI4XQ94H48VOX84+p
Dg1J9KOtXzoXZRK1t52WYrWrkOMBkVVtjajnzAL0m2UcZfKY8DmiJpfNy+hb1697
1YBgllGUmAvKMsUNxf/3mbSpY0sQ0tg9CSOCJbwBwVGQlXOLZWqeks0Fnr+uNLSn
J2qZ4edaT/tt3j1sJDhOYwYnvC3etct3VAESfhfpgbZ/KhGSrs1kd1Vu4QwKc+Mr
YHHLOUlPHjLyxAFImu+N33oAUxDya7Bs1zulVixLNpraonb7yoOooyPrlUjgmz6W
sWvIR9jWZH0Rv6pVJknhDL7B+9jXIDspSdUnYjdkFIov6WXjW14d+RIiXuCGQplN
b6Dt1OBURhSFoPY+7kxE9qiw0zuIMWz14xPOua3mjqEwNZHOWIt5i3cT+/TqYANL
1vUQh7Nx1eUpO1+pCxTYYlwG0eQ34ETXvGPWAP/cqCitZoUSkPjAk2O4ZcXljh+5
chEcolZnckWrS9Qx/bpU+MKpAVl6uDee9+th7YmUiT6M8EGdbWzRh41ZHUscpNIe
toUQMQxj7+7Dtvr/JeIoct3aAMB/c/jxIsBJ9mHu4FCQeZreHxI0vVYh1z2OoSTW
HOF3wLjE2UdspDBUYPolngjmZtVNjwNfj4AxKcOpEjHqG5sGJ24ZLPBNCRH1q8u9
72BNKsjrgAalkTD829+Y8RlINTsL83cBCXpcKOvpdrhoyx8zu4aGdREYljrPClhD
HCj1AHaWF+0bsbRssXGHeHyB7ig1w0BOddTaZdzaWHGsN5JBsWAbRrG3uzb6U4yW
NJuG23veLhE/fuc2WGkZ7EHVrZQnuzKkA7hwJ1PwXVPH6LkqCLjl+/xiYRfASTTu
JOTwhRalKRn0cX2sBac3BshvDAWBrqC9agd2BuwcAwej15Dwi4h+fdNOUxvfhPC2
73DQJuIirhUYwBjA2+syMd4015vlzXZXkkidPh/uzAn0mkDVv/B9f1N6HBA0SSwN
299KYlwvH1d4I1PDrK9lE4UuGWOOefNBCrTcHNkanmapCuhODZ/4HNS1cDxDqTvJ
say9hCDU9XR4s13//NQ8lj6nW+AxMAgO1Rcnjq216q76NuNKNOhyLx1CZWUVuEAy
0LlDZUNSYxmKsjcKlXVR0HnZT0qA352wF4kHHrNft4MWI16ouRGe/E4KyEryZ85x
RLUNqsQmqyHyT6aKvfic8ekEtyLeuiaS2a2WL2ZMD4UcF3ZcvdoqBilxLYtGPQmY
Jgf5aR4d6SgbDmuiOGTt/HhyeQV1wGzVPXUJxB1kzzoeVMHQF3qs0DvRyvOh5s0I
4UBkyi/58O4zAzj/86787iaFo2gsHYDURUUoHF7mgU+QSzUcHPTrZ2b3P6fSwBop
WgiAaFs9MH6Z+lRrv4hcQt0M/b2jYtG0hUhxH8gOG8x2Fg/mzoFXHayS32MpQHuj
KnVVnJU0ofM04jdLjm6aPSSKd7ENt4eHuaOhJGNDiLKZ4RIlPuza3LykGriK7O7q
5kXgkpbdlj99CzjQeSIRuChM1u1T3aEHEQioskEYPY9lo78nNGDYy5xM7//N7MPm
0mHyQjPk6kjeePCG5VrU4JhSnxMmxmApXgx0+nmYhga4k4vNuCtC0jNLSNblkB+k
jYTWL4wbDMA1fzpiPLJgNHd6MyRlhqtRP4CSf99mY0gC2GXWoMr+ZC+of6X6wjgy
s/QroU0mu/Z45C1BdyTOSHj0wdFQ5KVmDOSyWVadANhyDmecFF55DvyHiz0vR0Vy
kpYDeOd1QgpwUaFdneizU8Rk9sXABA86SlrQIC82GW9IOYGlxOtrZLjWCwqdciIJ
YItiL3XKMVqmJM8bpJE/vU2qXl68veG9zrRLEIySG0UMYBoUgrock2H+JhY0LBl3
U0dZeS20DM2dM8jvpNW3tjZ/1D/G8aEke9DBMhE3VH6dZMom0HiALCxtKgKPsqjn
flLZUdecT8UmeezwhNOwtrpfUkcia9pIqRpaqQ6uK0GyEal2EUx9GgKHkcBXTJTu
U6UF8xIxby/zUENcEksK+sZuyVL3TaabmEakR/HmmuYvIvX07WKe7kiuUlQyAEKH
ERuLIo0iQKGA3t9ZykCu8imsZQrdytAbnrsR/032DwX55Nl8nlVWreQwu4Pj1eNK
B/W5ZQUiWqwrsM+rjQfE5RpNHoyUBKpJ9uZ1v2h+ClrOTyI8+yJDuyjFL/1WdhPF
f2KhEXeVwJnzNoVbJb9Duj7xRdaOxKZk1H4+//KuW5up0xBLQq+3EsSXAEQTVuuF
xuPWhAjTRTFTyz0yu0B5f921NgKhyuQXABNyT8u79qIIadAmGGT9Gwn0307sdJZr
T1fqhRx8VqluULQzIcSb3OBcmfbI+pXQ+9jiSvkcHA8PxBo79KSWvI+J4Ct+WGYw
1eemnXRty1WOZdey5uTFdgaOnWrm037CtBbrtMW5KDQP2hXmhsFCn69eKcXAJc8m
AUvx4UGh8WUavVVIE7JcZ9AXL3uGTJqxlhRSwgn/GFaBZemKlu8hzcA1Y+3LMj7J
ByLWGTEIg5iavWyjJrSXEPnzDDQ9I6TvwG+C31x3Klgo/YyPgQ9EodKylNyrGXBg
a0L30W8wf7If6wzs7K5uJFHBCIAxJQKBGPPB4+QNcxXPx+5b2cYbYOS/VoT3QlU2
fs+qEzM0ERywUmnmD9v0AG7vGe0JqP4EuLjlc12rzCs/0lywZCZWkMYLpgmHOCEv
R4cv95btXikgunV9rTXGUD3AjGW0r6jqY8X3n6zB1nwIQGRqQFDEHWt8q9hDR4EY
4wsTZMfkwe7LkG5AmeDoUP3rz3XmToNtKqgcfY9MkdApYWTg7CDuBeUc5zsnW9xM
LxsQ+8hun1Za7Am5wL6mWirXPFPxtdATOMQpWKmM/gqdRELv7XzmbLEuEEW+x5BV
2U0vh2G6FDX91BzUwDXT/entjjcMclMKfPK5YvmM7XwxCWLOm4qkb+6aZpYZgQdb
xnUFuYoJUCwzrVk7srrbjH4d5d40a1F/OjeUrbroqCx3mGiN4iqSINBegepknVB8
fRK7AqEYFMKMkV6/wYU1bb0leP9C4iFOrPYJ2G8yCqB/wec7QcseLTDfFksJMgeC
yrzhcNWzjMCGXWmqmcKO8YFPOtItp3ug5aqX9b3c9IpIS1hKuachYRHUA1QNRXmp
XXiN7Qe11+hndorKDP4nQf9iAWXGDTR+5UxTRCFUfQrUhz4Wj2IvqTvOFAiLbXbo
5HCEQ+y6/xlrw4OOIJY4rSeVr2R30sdh9p4pP5JQBXqsYKyoE6aWZ2XJezaAgqqN
g94OPivB17XC6XNz5X0vnaouPj1ucTOpegtCCO8KmHyVYVs/FvL38xkkIS4BddK2
8tX828PwdOmy5RBrRd3aaxeIG9EVyrzeJIy6iylkgohaihfcBVwTSGa2HnG+2uf6
RbkkeQx82xCux+PdV32qyJgGoOSK4ozPEopxodIJl7YqVu5RmcYhGdJP/5DQFy+L
6rzYfWYHDDV7R6W/nvX8K2oEJesqvSYg/ENDjzovlZgi1YALIi6JZNZ80y8tKA0G
byEpWCwjSnoJ58E6WtJ6rv29vtnGEw4k3TZ7Q5eci9paE/2+o5exBlw3QdQqEFkv
6q9sbfgtOOAMgFdzniORuOcDd7ayUz8ygzYEaEXci70euajzsXQ3ufZgBzy7HVyn
bIxPU+G5osV+404K2Uf8pT99tiJtsQUGY/0wcC+R6DXxQjDLJPZ7ZNQFm+pMHLmu
IkkZyO4NnSV0/Rls37nykQdJCVHCLrxxpIC+E8KzWY1+SlqmUzJXeqKz1BzFLRfv
TxDoO2qzVVG+7I5dkiX4xFdq0KjEC48pwkJ00RuiARoLBSZh9isM7ov34YFhuFAp
FjSo3ftbSJ87ymgprSK0gunnLhsicEux0pFX6u18iKXvK0KYPPGiX35ZyXo63cPe
54YWIiFPOoGAv1Dv0AJwUgK3l4RLO3j+z+0U1Cc7AIqntE5bic/ERryeLNqZgEcV
SJS0nARzkbqmeIkQ/Po5+1ZtluW/Q651nG6go57ZzKl/SaGMjgxVzgeoV3Sr6FfJ
FIHcOKaXeUkgOY2Fs42/llNAC7GX9BEF3AYEanWd9MbLmLxb9FCJs3Kf4VlOK08r
i97RPvtqwFJX0hDUCYhVOh5R8gdCZKaE1emvwxqyjtSn2pkXeipkNQ3o251ovi3q
61bfoj8iQmGT86Fu2SCqDeTtGvsAEhFQ7f1YzqYlznNWOA9BJKdRCV+mGkfT3m0e
VdBdZVEj3wOCkNLNuEm78dfPsYXdyxyESrPzwdL+aBXyQgwC1AtJtjTdYR3DTUQA
osXSWhjEc4AkVcZXraH7PklDRPheEqwyRPs7zPYy+toneUkH7e8pmEhXvkT7Nd+m
N2YISIhqZWe3G1axthzQ8RpfC/De+QkknyLR7PilHJwFI8vdgNkbxpJ5Fe5iv31C
Ma8gexxFDKP8V9RooWe7NJdg5Eezdjz0xT2q7yrr3FNxz9nsZLdOFE5C6un4VeaW
12dlJaIbTTC3rFbPi6SJNuCffnBMOnmQKz6hZvPvdrCfhLF62MisxcNInNROhHRl
o7D7w38djUoI5RgnsErkMtvWNgCqwEc7p8je4H5ppUxFxrDOi+xyvL17g54Nv+6x
EXsVGLpMhFHbjSUXg9R6uktUjSJS+HMx7KWP4eo0Ose2qyYS2aBoR2mfKAZYODCT
8ATvWDt8dBH6FHiko5vtQt+/CmaviiVlSOQ5Sh4XEp64i+6b4yXDNhOgztzz093B
cqXFBowWOTKOwiJfPEh9TxYPVwnPi75DiRCBHtpYQwQsrf3Vuu8UadnM9zZkgXM8
ZI37Nmr3YPWdef+qKR+D8Mogb0Zi6JM885sM/YieGmrijmDVTFXr77/+7NIFNOSs
LGUr+pxef0P7ySO2jVv/BbuuA7/AHmR/jGKVg/pQU8eFjg8W3cI9CJB3QFxrBwhu
njk3291CxUApYBvy+z5TBNfExRj1IcjSqlHH4sOknnA0kgF0SxQt53gGHWV/rCD2
dVfrH5F8unJCB8OmpQCkdDtskWUoI9FiehDc8X8gy2eBF+ilc6aDh0yP/F1Ifdbl
VHv91ugGCa7WW+uzghEGPt/z76Kl4mlQGsiywTA7iR0hfE8PI1vtkoevN2BVj+ZP
1y5gMhuf1jBd8ESzhAqMV0AfbETWME7fcgOahdAizqUyOvkkgqYGMQc2YuPkZesT
TaaUeTvBLYUX1yXeiv7rV+RvTI8LaLlkKYiYr2f1lfdojXA51pEuAZ11CgCNiZ8Y
tWIU5dJ+b0spX6nDRe2ie9+DXLv2tPfv8vBHCb/YqErToAfC16iJpK7GfoJdCKNu
qxYL4zLIllBykRJFISUbAMt5ZlzINte8ZA3sZuAQrSZQIB34k+CSKeImdAiS06Tm
LiJEsKhupufDvcZZYR4mfS3/SXGpZBcekSt/SLiZUpLvpmQbiE0YAX414j69GjhD
gSm+s/gTYSg6mn8gMA66YU37ByTFWbMn/ZepaSkqsWZ7yexLuwdq6YzGxtx9Nnto
jreyciq2JaFpo+/dGdQ9F5oQk6I3iFOsxwbnbwMERB8G+sGBL6Z+bszxFXmVa32A
NbyKWihvnOc1B7hTgcc4GlghHvRsnDV2zJB5p4NqNaYuQH+pTJUCUzAq6RYj+ktr
h00zeVAu7276LBRVyteX0VJid+hU5uT9nfGBQGu52BUcNRk9zOPDjpjHElUI8Y8a
gPNyisbfNuSJhxFfvUmfp58Uqpkp6V68NW5naF4u6uXkvYn7iRwsWIisV5O8w0yv
hRalI6hwizLd4ysTVBcQfQQbxo28rrRLjDPtkp0WRiT2229GfWRpO9fnflJqN9Kd
JHqqI+5eFev6vzbnQ0bvB9j9itpbgzqYCj6eoPZfCr9xmlaNqgq9Z1MmruWruEt8
HwxxpaGaJIvZuo7PR3WZJKVmEwguHPFWPZZCBUq3DlE7jkqmnoikdhj8zNMBXaIp
sR5NGVqtBBTWj/cFKPei1x0rr1UsRqAJaHdlP+K5USz5RSRupCvLDggpHAt1+ikx
471f79xv/+IGbNRGfUmvKi/Hcpqf7Rf7SqCbU0mIbJ88nN3wK2Wlz92j1miW4UTR
ExuqRYtic0nuwXPhDFNtonuoHPpOD1I/P/gtZxzplkH86v/L+858sSTX9mpl5f7b
RONZdNllBuaVui+F9zGPy5qw7NGRXW0rn/v9k73C0VSDkGCapuMhFntHt/2S6MMm
y4UNpddI+XVJ/aJXq0xR4KwwdMnzRybfDFt+trCIn4TbjHbbM8m2BhZ/mXOEQq0D
LtaFAKZfhFZ7HWmLqpG4jNOhM80ySXuNkXF/4iEAW1mRBo+tvkXevrMM8r5I5KDX
k+LsYucj0dFMA03pCtyhqC86/EFnmZK+tsGAOO9QawXWIp2iEehlRsMS8prIrdrz
9AxiU4x3QvmNYoHqxfdGoFZSTD6oHE+1R/DGq9kH+lqH+q0fgFWRn9fUIv6ryGhm
JJc5xn5Oc0qreEj/ZeLU2GTZPZ9Tw+z5LNEGOrV5wDnu7I1Jrf9zreBNwhU9EXzA
bdrB4FbiP8CHd1r2BsriZqSA8Dkld8WGSS99TJdVZoflUAYEsyAx7elf+YNmZftV
Cp5d0Ijg51F5Rx/dr0+Bw4+E6qmNp65HGmGeQ9ixmUa29f3VPE9+JfErhLGQlUm9
tuXmHnG1U8fT+l4w7s2ZAkHaoUdEL8IYlAtC7DFhIYm/NXVACmc16uJHyHbSC8xt
MozqtFugvauXLlBIxUid/9KJ/vQtP648SZbu1pwssDF+5D+N8CVxJFcsB/MLN+mv
GAShGmzttx8t7756itd4LOwMjEtozSpxxOZvtrZFO24Nww1WnPpGeEswwhj0WA96
tP8Cs57Ak3FsSlE8K0HgJsiFFXGWFNhv9LcdhebD49GparSpOFe7vZZ8bhybiG5M
X2oBihgK/4l+u8pezHlpt2XKar67pp5LYJTI3b9ENs3NkGTQedyIy+w+O8OkFQ/2
SJ6XmgwuRHcQdELZW+flLV8N7OizN2+bij7giWSHyvgT+aF+MypAVdZv3oCK8UFT
zC3hi8I9ycef1e0N7SKYsLPtL9LHx8eiCOrMHtx0ChzEXPTp/UFJZW0wWU8NzGtW
nvwtQC2TIgKf73fVM7dowfTxx7rLKJK2K/uX7TWCBXobJWKbhqOmdhtILT+J0bqh
b5ne2ki1nKEpqZBAcrBs9awDuETIGefBvRpuli8DaT0uJAsUgkJQAzZBOaXqQDnA
+/GByBHQfg8rPh8RzHLB6Ve2nuff2Z0zCsy42XMaOmtoW7jKUPvYYWt4m9gt8eoq
sRx6t0f4oqJp2alfgXvuyBMMBm9UZjJq75ea17cx8vYOhXO4a1uXRU8/at5xo4IQ
eWpU+QT+Coh4PbLNgpLd3E7L+yihL/aRyADOsYL+gsHI823Ln6b2SoFjI5UssQ4g
cwh2CKqSx4Ny8CQGpQpKGf4xehw3MkpU7JZrqPbMALC+GR5day6Pl+EoGqnc+bb5
H+FuiSDpEWCHlR1Q2KcxL39j6HUiu8MWKpS/6lVjk9Cor/MSHQue37z8weB7k6tn
49P1eR+tyWe8lAPp56nBg/wPGUlpnl2M2yzbG898gJKqoTTMI5x/+mFtTgXPLO41
oTaBgG+DDMeQcrDnoTR/3HD/255JKlKFe+pUKoO8/HdVUyAWvZp15mFRxIZAj1DR
zJctjGNfLEBalM4B5lJIjXkbfflnr4EpmE+7yAOWtRl8XpRRLhiNDP/jwXq1ALuz
lru5j83eDd0kq0nhgw+TioSfcSiQhNOjwTgmXiO/9iFt5tVsFdwHyGbWpFuSBKvl
Kxb+5im1KT9FAPZFu1taaqiV9DRQqk1ziQF6Hcm706S/qVl6Z4IYaRngWEZTdHYs
R8MZ7Y6XeFS7xKzvsIK5d/LVryAWDJr5wHAC7flcypWtstK5mu08q0KnoaHdyQ6P
+DE6IHxZAHYm+Y6rUbo936QoWF0P+/smWtRl3BQBuJRA0lGkVGolxDFRzn00XbFE
pm40wGpzgzdItwxJ0EFKqDA0Aydo/o3D+cih0RN8pLOZMX3xzVFyHk21fubVwiEA
sbd5m/Xms0Hb01262zID9HWqw20tkkeWmt5J7u9vG1a2xiOC1fa5JI7VrtEkIejt
fKGXcgPsdo8DpHtupuCKBdyZUm7qFu4b51hh5wdr/R8fRvKCmFhln7NWvrILIELz
ynssqAdVwTY1x6KhnElE9FBpkK/EFuntvcUWQF7GfeaEg4xfau9Lz2rp4fnhXDuH
NdduNMTW0kN8/9OnosxoOKVtOjnqv0kfhE5LUre+KHymD/x3ex+RwPlbPJLRc8GK
8wXqS1AEelvf/f7jdjjYM33f6Fblr4kj725HcvuPVl6SwWXXLD6hFuEcCR5/Q8ay
c+Bj1otu/vOSMU6YjGZepeDvvaxTbXp/FCNz5D1ZVnXVRbQ/m7VfKy7fnVGr+Idk
4zs0P3sPz+y/iqCYwCMEZjzGD3vLb18SBV06z8KsBVufCxE/4jlLjly4Pemb6t0D
DQL7Utb71R38KbYcrLv1KTgRkKuGfuMw2DFzEh34CtbMIPQAOSE3UWAQxyl6sIZ9
Enhuic/A6gHb7gDw9jiFR/xTN7Boarpu3vtJ/xZpjpgzF+jr1NtlsFqGLAOYB9V5
ABdHUaZQn8hx3DKIo5koW/QiIKaV74w5HIaDK3zbPeZ4ed0eNLz2k49KpwIRhuSp
GnjDYkIYZv+GsjSCI0T8DAlptg5KPL7Di3BTxdgf8yUs/Xjk6I+SPt+Y4yg33OeV
1BVZq8Wuzb39yGoK+4t+M/TSbWKjUYqRsFhZjyKfv6M3RoExCqm/WO1dMLrve5QE
jivBmZBvgCIXFnse0JgKp5uv0mF4hjRz+VtYMNA1tHo36cRD8cu6sjnTs/B2AO49
e+P4mR0LfWi9U1bkDNY8zOIQMDLi+SO8ua4vBJw4dp86Uz7u8BEu1yyA8HdmILsf
y3RyMCaSZVHbkJUEoX73jDB8RwjLPKjo/kXJFzb5HFOckpDQ1OSYn8u2hOfSBvKK
JaFIJV4uoMUiwuXeF0oG/uUgfnJ4ozek2nhBkIhZVqvzWjDm3I+3O8zSpU6RizLd
8qektMrlsibbKFNhACkOUF2Vv7nhOgV0prs1h0izrKLXU6Xd0z9DfCkrlpWPZhvz
Y0PNfDVQXtNddAw6SAlQoQB7XAT8clAhRDMeFl4qApbwHIx17DPvXHVTPJ3qtqDH
lvsqAUq6nSNu6oDyjxshim6XLM3C9v2hvcyFUIAzu5RoaIkjoc/EVszrskKijJnQ
zv66NTGeXuhIBPW1bKnQNbqlL3TleMIfE7BxK6oVHBi0JaK250PuzSBdYIBJ06Vr
eN0uGyVTDmAOlluFzrbbJ6V3+BLZwDgy16LM/OIX8xXe3mbKweIdQSbQ1UfJSHXe
0HlQUiYcmutETzv0OuYWlhViyCLvfduEuWyjfLhhLCv3VaYkaGQL7obd8gCUVkWP
BGxKiW6KHKIvD+Ld/rxK9qnNyP14bm9vRv2zDNpP6L7yiTYixUc2OA30usSftpZV
QBR8cBXcspxN/vMfQM72wyBikP28z9EUofFm6U4gt0tmyvq/EX27E9TnKJV3L0eK
9flsW5ZbZR53pK9PjGd5XmqTw4o/yp0ZEmgVKt7w6SU0bJz59Po8ytFIBxcrlrc3
I3AF3nXQA6Jxn0uYI+YwhsFu+s2Qm+cXM8OK45iCWa8fzQdvA2zN3kMCQvW+Y/8j
cRSOSO1YjreO3VvIdmbtbz5qKYyDKBqz1WQbUdtRpxFCqwjEjDneUXM640BUGi0L
DdvYV/+CV8kRutTTuVrjL4Jp9oOYl8gemDoN0eug1qA9m+9/c6uA5MWoTVNNTAOk
rDGFRD2aC3ob1DzQDbqmHJ8QZgF+yhjppYphvMMfxwhjgZF7kfjyCBVBgcexediy
jyD87rnipI7ttq/M4XlTTPtl9GtmevETZe1rCn/PyNuX4ky1BC/kA7PXumKjsRVh
qd8cwX4kQu+J9a8v+YR904TpRveItjEFqKZvf1mcg1uFcnqyNu+CdEDbuAggwD+s
bxluphQR4WyQAPc5zxOH8e9m/uXvpK4pbzjdtNKWvNhqtj2t9S8C6e1D29m/a8x7
v5wDmPuYvTJ4xQ2glxgttDhmQvImeTJndRUuHI6L9yDoARcKb1qqGaHOlXHtfoSR
Pn6Ve/3GWpPFfVkCmk4NMlX107jl3qK1lulxwKVouA7QGVUtzvION/8opok5ZYEM
RstBWjW37cHV6ZuhEQa/hvNzoWsbCqnokwxNTTCfrWvyHGYh/95sC/y3OwmEYDvM
sg5Uz55IqchUeIj+LMsa1yBK6erS0Orf3n1tfKfgnGrcyjyC2FvoePDmQI48ZURQ
VwFQvOVva1aVPSM5OWG6SwNqUVNrDFaXwnjI/RK0iYKuNXNFGe4440dz7HT21aiC
Ov3h8gHtqOcSpPhxnl7Uf/27OSFLWo1DZ6g943P78/HW8ECbcfIcTwUEQWRIu36c
7ExkXCPoCu3NFrf63p1BYri+RTe3XrZU+z6duKPFKjGxNaV2GWth2WSan256Pafn
pdiE7Ace+pyUdMnB9tu+hi1CrOxuX51S08+E9rbH97PHl+g2t2gswzsVw2McSq3z
vv0pC5Pmw6ZIE6E/djbqcuF4jKlZKXxvRuedu8QzVPOvxtUsGOnvnpcAbQHQpk5S
IsWX1RaWMghYVMYRSAv6/K1tK3EoF5kGMPPHOa2B6XqETmZw6d9hxE0mj2p75wyV
Y9ZgU5vP+EG5Z2kCRVHSLHyPdtZAOq8suto8oIzX3+O8TbKroKxCFbwsWpeu6Glc
Crmk6fppR9lhxLns9Q+/q6BQs/of1d0tpOLy4rim3nuIQnPD++xgYos/05dPizj/
+pda975rkCMDJcSvalfokMdXKjnLYyMqJiTV5gco+p16f4TJG8S3C75i9PZjJtY5
t7VXseoEE/EBoYTcOzlrETLK9Jswug2olvR+JhYF9yB48t9S2caciC8pIU58NR2R
IQPrlBqZwIppYjnXqbA6t87KMB2H2UgihkuuxSGnMAHRXnh6JikWPGb0vt89tWW/
AuuxJkVWahQxQtB9LJN99tLE8DRYuC+5LI1rewuNP6klIEvRCXj5F1RU42pjHZVI
7hT0bJgfANIAE3ejvE8DLNl6ekZJWVt+MERzh80UWDGUDLcoJfrR8ujUsko4uYIO
qDqzZ5Zbetr0LOpGlR0D0rDIeiqrc+0MFy56Z43NcDrfRYNXTdqOZBvp5+vUsdqV
n1kt7FB9HgFDWZgmMvwIvQQ2hChxPDjBaLzaarsfq15O1NBF8RUbkj2py9C39Syc
ls/wkn8O4hw6teFSUPnXtUKYRmThLul4vCWgwrlq049ICtVDvx1+xHq7He4eafqC
Rgyurq91s8Gzil6iJYpo9oqDDIqE/Du1F+eDLUWzO0amF6q6qgBXTL9DBiIln5kp
GyiHnGMAmCiH5f5bGIOMqtej3IeIy3UquMH5Z73xEdr82Ks+gu391odVfyFw+zc4
PBRE87RW+7Hbc4vEOWgAwjF0pfCasIw6VSGpkh/52a52jpu37qAVhxkW1u0Krlx1
NLsY5NQF35T96A4B9b1ExB3p2wrT+qQltyjBbyLxffUNmP1j84youucW+uPcaWlP
hLOqK2KTy5bRP/7W3duwJewP8phuI0GSulQBlIaJ+7ZK06LE9gGyxiSfJVSqlwkC
PP8Oq5hfULQo9qNo3e0yVe5atkfOSQI0wnMVq9QfaXEy0cMd5wKfrMkySruzikEZ
6qbrDuVnxSOwzZFi3ntzaq7FM/u8sXIImGfzwGJ1yzRU/xcDzIGrkOWG00YLR64I
O5F+NuBz6rXmDzTKgYJZxtrugZ21KPCh4KQpGtue1SI0tX6Cvmrk+5PmwAEMTAub
R510e5ed06FV0FS2MdP1AsXo6ite/00SVx4vak9lLczD+zHrW9rJ9WfZcwsc/W3u
I0E2Bu1xD37U1t9CAlUpaloCmE/8rtavYZJSLeKryTxpLVW8fP9u5IzVAjUuJ+zf
4PUEVa/Y3sQMCsNlvILFMNCgiEtRBkJPeUoUFia547NMYtMjQwHbIsGzzTYJ1vVA
DOmVpJUS0Zxulu0VeUppoKaj8yZ5WjhnQudbCulzqtmY+c0AGcuO3ZWWeArUFIy8
CpBukAevleujZWqa1HksiMVtIE7U+2PdtzpBJ0g4w+sCKH97huUNqfg0oZk9v2to
y81bnfAqNbKECK/2go0LaXGGLeDeP58fNVQayn6aXY/DBj0LT/QD0R7sKJglA5m2
dlv3cR+YDSzf3Yn2rhOm3S9yAc74e0PKefiZXwZjzt5bdZxpWirjRM24PzZxfC4K
MY3E8O5qoJlqSEl43qRHPZwOmVCqoOPoXUgRCGDYxlt4qmN7z2wt0iatT20W2xei
lxPEsp3BQ+6gV74/TKs2M2GMdu+tKi9isCDCvDGo5UtEYl74WlFQn3gUeVAjGA+8
y16lEGBz9KZFh1aHOtBLQSOBByOiqM57QwWp4XghChT9f6hJM/yF/ZuEF6EBA1nH
jXbrO4Jh/y9zPd6jdbK983mJQLHUtoMuK6hvSmtQ1lAQE5eqR3/pX4Xq50Y/JeKQ
KVb0MnknR+qR6zq3o3E1JbHcqEgosjK/nkXfkuEkm/KuGjHufHZTLcOQaH1lTpVp
6pvCn3wj787VYMw5u2YbL/BG1R7qsvFryx/JZgaVM4nIaLESoGw4UrRsPiQiQYs+
Yk+/PdLqVKiXQnBJUVcOynETqp3JHLF0l49/cNSSGVRsVzWD/eWWXQSt82+QohCu
9bcAHNA7U/D+PDaRMRyhC89OEE/1pZhr2W6PBN34m9IYYF+R+DjRhvyumdE413DC
jJhlaCeTNJsIAtWig9Zje47fugjK9OivMDYf48NmbZJYI/g5h5aio0Ia9WE55gIZ
YZn8meYviOmWxx3wO6lulRhtOSM3vVqTncXKzLaecsUWDL1kc4osxG5WK8T4AxRz
LwF81Ni/3qoDF2BcgfWqPg+YdcNGL1fXahtBE/LgL6OQUUoBwM6QxR6jWOSPWTCp
ZW11HDcP0qiq6ciUw84mmTEW2Igf3QlYQRG07SO1UqXuqiYXqrQEJCyuRdvlQReL
fjR9H2afF/Sw1MuNIUPpwsW9DX9edI4k8yaSeKNU/QH3+1H+h7y5SDImzLUvfYVc
XicRlzqTqpUiyFhc1GYHR/c1OSbQaoDwTKNbeY6WO5hw9SLzNiJVs4735CHTSOQJ
Dpau0+ePmb/B+LWGji1X5uJGVzWpdvbUiy3lTd1ZjK5lc9Z3VCTlLXGcKf2W8sEU
g8LTjPrjSYsVvhkFki3xtP2ktO4v4rdbgFemHHq05eqjySKTVs3aA9xVYqix7hZL
6g+a6QgIIUQZN4FxDLNmhuq8kuozKEt3q94mJLFyzqPvI0NsVNg/lUiO8thZtkSm
DgRNPmn7+GRjlZ5NbIn00j6YXiQqMixH6EYwvHPLYMpBZ7KQIFnTsA3cekVPnBhv
+DqZ78XD7ef3Cm+dUKb7g/+t7BW9tEwacN35F9P7nAmQ3etav9nDRemCCpI+EgDT
GmHzCGvfRIU28hdgfxAbCVIrmEsX2yHWSlHKe+R9axuiCUDfoZsX8NMo0iPfGwok
1JQBrn+Ixv2RBb0j105qLagEX1SoS4k7zIb+Du20KkbP52ousfTblHeygKvzeJCL
TIoVRxCd5I9I04rWL7qwD9dg/a2yLtnpXPg5cviUiytbr2gPpoCbmuPf5GGKSVZM
Db7GjGWjwaHbcNmXLBqvD6aevIz9LWZr6bSPaHVn7i/I6nPIeD13p4lX7EjwZrx5
jk9K4S8eKelGvHwuRMEmOheNTO1G8rSc+3eC47qgVPM/hVONkPpFsuTFZ03W1m1p
DzxdGddEofgVK3soDditXAWXXZVRY6OUubJ2DDI4k7cgSSvX/TeISyUah4Ar5iNf
gcGrS0zz/IjCUG68ZmOBXGEOf6w+/Ai0tpKiDiaV+ZYbnm4+KP37fzplospZP0Zi
EvtUx3w5B8kxL9c9lyuAvwftpTPnxfU6OJtkXlxwuGYL1J7n5GV0BnMwtO+q4GPD
PONFoAdhAo6nwI3LUr9BJJTJmpO2t3W3j8FylvXEzWFwPPmr23LVoJVzCeij6rlW
d3Xss2WLmoqBpe21ZPC3WHux2R6t/5ICgikxKnM0W1dySu+4dwNk9plh2ALQA2O0
be3+zos1w2pHCT3gAiYhYVm9ZmykfHDlYnAnrDDWv6ra97DorYqL9SVgLSw6tg/f
GtJ/76BcgrkQO13WME1tG2wQUz4Wih6iN94L3jEn4TOJk+0mYR5yi0s8KM21C/Vm
qawhe8bqPB2+dpjIPkW22GQC6njUvFP7xR3knV5etTomzzmy/8kyVrowLmkgDXTz
vVT1ITIf9Up3voJh6I/K8bEQXmXAECbl4jVcQ7dvALpfhqJZxcMWlDK5Z4S6lMQZ
+Cf6i0aqqMG59qVwjIOgj6ItR6EXb1uENOqQXSsmMUM5d9wqw817ovMEOsNkHJKI
DbBQvFoFy2uIVkRSrNHIaerG9zWLOukkfUN7/IeunxzfaaOJler21+v9+cv4LJIB
b0CXrudOVasHGeYq/oIbp2tLbwT8WswzN1ocLDmeF/7gEobOvL1K8oHp0WeznXmj
S92aaDrFQywiTzo3qgW2HCemDO2Bjx9omsNmjE2b/nFfcDbyAwQecaAOBovJPPGA
ztjhKiub5X0KIuKS3k8H2LDMEfKyqyLKr9lFa5lKOHXrp2DVE8OD8jqqsbypK7CV
O6sgH+ox65uUKZGMlMu0yKwEAGOdUyZI6AeFgYdOYqqPQLh6CojKQdlQ5f1HO+u5
K/kN1y6xbrPVJwpzmoVG+UWDvuoh5LZtmfc+MISmI30G0bfYvzN3pesBo9Hck98J
m6FJVZLz8hR2aOKzD6daW8AaZ2RwAqNQDHLzVYthkqDJReCmViZYf246tVBxv/mb
xlYc3HI+lLbV3KRa/wU14K/VVE4HMCDEWmAYbMG6wa79kHJbELXBvFtSZ9vezvYr
8EDbizwlM+JIc4xU3wqWotf/QRA4kvjG9+aic98seSJYuHN0GOOpdt/atuuPkRD+
fvWdoE0Nzj+KK1hyVmIm/3dHj+8/1zLZZV1AowHp4xx4/YdkkN0+TObiP9wU7wWz
xu0vKpD+QDKODhXnO0UEDm6JB4tmJPhdnAoyM9elLmH7i+bpSmdh9LNmUweKXjiy
lG1QuL1slQai8KM4yTQfbYjEhfVkGxFzl0pq0bZeb0deorpuiMfsugpANJJn8ZVG
VR+J3Qe9/rK3bBz9aEKcQT6PdMTdsfZ0wxkeovI/7/qS+sDfnmleaq2hrFjBqdkl
ORIhYttM/vtpON/Eiy40ET/+Xl64WhFhmE+WlBFqQuMDgCV1/+uOI4fAFdZIAznh
ZQzytjzk/BXI9W/Ssc00E5zcEUsbN0a7NR1djMkxJbcw4wphDd8D3dR0e8nulvjJ
BLRXRWp4r3/LVV1q6/uq7CQcbKP6sQSecsdIFLEjCdejgtgN8K8DoP47ou4Mh/w3
KvzKec69UKdGh85zuRruTm91Fz+wpQ6KxgdBivMa14P2WPMmeUgu17xUHaV4GXY3
6qZhFhlcu9++vMMIuzdaCChOzQmBfe0xysak+SmeabIOTfUm/5lzKsFtddUlfsRR
j3dXmJYpPMFKn8tg1lAHbCA6jo6pV9noHsbW4M/dQ3aj7Diw9yQRdADjAOuiAZvs
mSqVLb8/GhUbk3ejlzhaTEA/H+zHObzI6AcMP49M5mVht/ogdz2i4Vt/YOFHyO2u
T9aWBQY09o+yTBmGW7W61sOkpPXCbggnlF+40aYCR4lNDmfG7EmhchdS2w9fFtak
tWCXzmj+Zq2jDfg2HXPe2SwjoIvdsr+Q8eCLXLvsCvoWMiMFYXHLlE0fl/hrEDFc
fUj7lLM3zPnr583ijI0A2EIBtbPakd6raKrY25lXB0Jar1i465U4g6zSe+gTmYIm
ypzNl8edRyd3Gj9uiHQgdYmWsqPAQc67v8NsZBa1qZV3I7AYBr2WTVYMCUQ6aQPV
mp5cTDAal4bZzgVNXZcEcR0Cwca58G+/fh/lEFjTYulLdw7kcVkABS+FXZcVhRjn
7SL9rrzlSvCXCC8aoBbzFC3bUCGjsL0+8ugNvBATnVNieENaCGVOwO7Y+4qNbXDH
LaBxb/8oNHq4vXUBSGiMBQWDILUUzxDhigIH7N0l+MWDVw2OgRkEAVX+PuXRcqVj
k5mL6na1v3AG3nKKkA3L//2TegWEk2l14HljstImY8Vjt/Qauz+4v7EQHYQOTYik
dMgVZrii347hdIhYqGi/KCk0ejbUxg8Cjuq05HcfZOKVWQb8IPXWvwKYlcxn5ASG
2kQGxH3IUkHtj9XE6Acd2mIEGrh5OO1JUYBZriaQJz6Aw6yIrsXZtye7YzoJSd7N
At60Dl9zAV6Nhz23gv1AGZibt2BXjia95qd4QDAIOZU6DjQyeyZJiHCKfBHGdTwA
UH1piANc2sj59meM/0J7ty9HOGTNu5jFXTqwhHYbJnzjcb5CuVrKTmzc66VdVbhM
2zgvhBnMleOAAtL7Pu0BZVtcpSAVGiCTA8bxDkdN1Hf/La4/vLWvNdSnI4+QlnSm
P6TKpIOcGEX/qDRBdhhcZuOoWNmA50XFMMS7kyAVVSpurCKEp20w1efVKs/94f+p
yLVq6yVonlmk3BNK9K2J14x5P8aeSUADV0wizraJ7SpoOPhm2rvnW0UjgLNNAsyS
fdVlnxIPWW8KmUpYKkHZ5K8//mVpBAABKbKnY1Hptnt49+0KY+p+7l62w/jb1O1N
yILwzjjB16UlsZkqFzARKtgnHe95hGa0ow/eqEcdNG2Cm2Bs9ZCw5qSOJNnbP2op
+L1uA2LhJgF1Qm+qjg0VCISVmWufc00V/DRHJrYGQX15C3flIQ9qS3y5wx+1jcFg
XOvIpnHA9Tw2p4MaAHHHyu7lC30rs48pN+URgCTiDe0Ilhtg/ERBybG38w5dBQfr
8ENBZZK7Um7ovnagM1y8vHjf56NNFC/SXSQ8DaiSusX2nAnZ7co+cvgODeWS+wS5
W1rC4wTWK/LZMBEyEHdXRSjIkwSLIbquRqkzT3LM2DlLh4T+dX80R3igojeWG0bC
YPCJFSHpXdfmWkUjaiUMj1x7QFd8XoEWLJ3LNSS12gv1/F28zrQuq3KOZnNDG5Q7
VeuT3shA9sD7sivQmPdMO4XZ24AL6CWcU5P0zW+OfnfWnxshI7bWEoBjKTLwlTjT
hx/xF/TdVEQqY3JS8RN6eKKGddXk+SecOoLKfyMLmCaQj4TotKOkMCPvo6agLNcD
lktXAsFdILLD40sb9A4lvfRduGr78QoIXiEWSg4b16C8iSwk3XacZt1H8J4Qqp1J
uKnCe/CS871uVlmbSLXO5uqWv/8dl2KIO2Qd+X8lDeNT/Ba7zvXpHbEqv3Mnki4H
G/cTmciRr3r5IEdwjthH2ta6kK4hsX62ccsZFxfotFaImclkvGOTevuqIxxX8bJy
XN+lse+xXUiin0B5i9HyX4XDo3IPlKsxYuWMZY1XB67i7HP+sDSs7gf9RFpCxuOD
616ELokrIzoUz+r1gbPItmVxODgv8zeapsp8msZbH6f+Pns9t3BhL/tJw6ey9veh
omq3182ova9F+wIQYu5HO4zg6IIHqpVXRIECKGjxHQTfZykZR22SSeMLv8pK6dvK
Uzn/JZ5ceNvX2GC7tjWBn6iTRomvyZ83PAejoB7zr1EElxz9fW9sLe1kXRUYlFcd
Qvy0EG/BNiCad3qpoHGzT5OZCHIireaWb7i3esPLRDanSMlE32D3kZ8EfrhLjcW+
vHKIncf7Kk9oEvVayh2ZF8HrpHLFLNSlUleLTwL6fBZjkOOqb8RA/nYgvKNu14nZ
njbGSoCHK3lidX+ZpkvzXb/XXGugA+QZJlbIprlYw/28e+E1duFgCxiWF+L96VUt
bCFPbP7Kdt0gl6SMaY5lwn4oAX4Yn3qoOrqFMR7cwbTz2XcoYuVE5pa/xJNtPjdo
G7+W76WvnlwSzfTLB0lv8HcJZrXszt7PBJu1yGk/z6cNInWMtT5BBxMLyAeMZK4f
/xCwMiXqpKuxWOnutAiS2NPTi/wWCiwbGtxTBCFtIKEfi2WxudxWpOSdLaSlxqGq
YrjzN6LsO3x6OtdME7uvaH4Wgrbq8SFsX2aMz2A3L959YkrVE0tz0pC/LqIEbVMS
XA+Eu9MjquO5T/gO57yCiz6dw/d3gqXpGYazM/iy7ogWqbUGMwAJAlChGQzgWeug
tVTVJnystXA1lVLpwyPbx8DENt8k4NgbNtWYJOf1tDmIZHmF1Tg7UOp7ScLcRG3L
F5nCkDOqKptsqEg9gq3BgZsjFT9smAUOHiXTrs4JuylUZ+m/OlbMbpNAbFr8yuM0
582EzllL24ldvUAtieObSDn2YsSzfg0yaF6POTNz7lg2syF9ikhsFoAtZXm3VEvi
AaOrxXgFdm6/yNp/w0ZJy/jpBISuPZVFOTuLbRYDVPcdihW3YlRrds4GZFtngiuB
00ZloLbTsk8kxUh9BJVe9pC8mQeNdcAM0biF5Sxfdk1JzZCgFEMYaeSF43BMD2Cj
hhkiya6QLCLuJ50xjk6b9Y1QqoAqK63IXvCTVcW4POHbpeVMhy75wQnPfhxpIYCq
GG/PoDmdrYDki2ELKS+Ng0TUFlVca/5WiaqCb3v2Y1KqF0aujDd1yE4at0hvQuHC
uS7Ix3BLo0YMoJO8j+fVCMmcRt1fb61xrf0a9HPWlk6nnDNQzeQK2ugTiS2jFMvP
49MNj0LN6BQQtmE5AXNbCiyW1jKW5W9XlqyV112m/FNpeYTYYOnVIwlH6sTS8085
4urYAueO7r6baBairmVYc73VC32UvllpRapcf+hrsyoU+wQ/bdm2htG3/LmtC3zD
73haC7LgBRnQ26RCRSEV18jxcJMSfHZYJQN4eIR22OugYkx5vlgUyuaUs0uYB73F
KNg+9YOB7Ybilzf+1ZguyLvRufufzUpXCHb5z8D3NImkUZ1VmvBkhFI8iNTxXbzY
QznDgpjpO1s5Wh44SDGUzPqDPPnsemBp/svErygB3mPBTRuTjT1Ou74z/ZxhEN3F
fIkJepJerKsc4wSMg1OicHvbp47u5JG/Pk3HbRH8IOWRkYXMcUlB6Es7BnwrMOvz
PtHu78n9gx1xDLMMGiNKyZCPB1BYak2DyNRzaVJ1ceiif6xU3kCQ1vwkAvxUVvNu
Tjo8aEr9u+RgLazeg+wWpLq49OiObDY/xKLdXxipMeyRWsjclKkic7/umX99Er0J
SYdOjvLwDB23TU9L+x4WTvgGfvZgrWg9YGX20YMVfTFPf0jSD97wUq0Ygsm+q3fz
tx22K3qwnOUtf+VE9QZSRtTjk0ixEdxuG0Ci+GRZOKXqDbu0WIztJ7UOuCeXHiOp
cX9mFTjh+gpy9mIcIGgbc/FkA7Lx430Hn42ahMEHAp4d6TqrY25F5sN54FKgoGmF
hrYT8aEWhjlo7rebwQ+MzHNlRcSJuUT3VGTW2FSucS7b2eAGNOgv6H0oYTiHmaJ2
wUDDNmSENN61DNHQtnrvpoV9PBIbSuMPpLdQaAbTVxrdH2Oc7ECCIC9T5Dacibxn
z1dAYS3z30Y5dSDzpcUITOE7eVKqwiiYk1XPVwA74DnSgbm7R8tBmE41mrMq3+E8
fMy2vzBr20Pe0erp3jHfCD/T5CElsZ71y9E/s7DdgCzZC8rUUuLRJjq663c2Upre
IIu+Js5tXo2ffYmKGl5tNxonlMbZDXtwOAgky8tlULK3vjr4uZq5PUcLJwXUUc7Z
he9BdCHp+1DDXtUOL84cEPsAmEGjBwVFBaNKLiDn2nuaIUFe2g8eDBFfHNSwBXxm
dZen/NVA7ZKqBpvaWetbrkRu2qHr6WewHiHJpLcNkEhBXDSU3zvxkrlx3Dw93a3r
a2FUl1d4y794HhEx2DM+sTRcC0YwKV8Fr3vUkFwkr+8AnnQ44c+HL/o61ZkDvCag
McaFI5AXpJ1HcUSPTBEaie0sBPfkXPjoyG8jcpkeHxrM1U0bPRcS5YoRKLAXkdfd
/EdROwFQ4/dqVNK1xSjAVa4hwYmhhOJ3x4MMmTCwsCrLiqeSMTmDISl2Hc+kFXm5
lvuVUgbHUibkgnCPwC2IhXXNDs+SQlIyft8DOr00FGjuQ2ouoFGgc+2BtTocnbXH
Atp249EQbijihjDfvUb6gX8axBx8B3a615TvQ/eOz+6Fn7IOHIeGmntNoi87aID1
Pa0wfLJc5+t1QQdO3J1bXsxxUZ/ti86Zn7n+b7bU68e9Mu4fpbneq2AWykGlEUuy
stHxRDd9I3d3mYWV7TNFtP70F9rdnaitEzzX/oO5PXPJ35m02wOszQ7EZBsKcHRd
TRzLmKchfmf/Q5dM/Jdnb9uEfsv+NnRrRm3YoVpJ+t76oDnahQx5fb29IU97LtrX
etlPuxt7JZmYeFszX6RcNj3HNFQZchP89t1mty1W/j17WK8pCm42YU9zN+Ctw9OQ
TQJ0HX7yL+juWfpmL9KCoq7SYBh3tqsxDG5Aosb3hMSYID4RfiHHH4n/BYLnuaHk
uBPIg9wu8bV6lj9G2tGDreQOU1qPaiWrDeLPkSFaEBSl+d6jOHWvtzKNSS2xoYdY
E7pg/3sMTmusxwok65f5Gq8UUj1AHIKW76QtoNnfmDLFepuKkzCat72DpdNBdUAT
KMb5TNsioebQ8IIoJHmePzK0T9fl3cSLFSdk3+kh9AwAzmY4RYOyzmY4tW4103fR
qb4q772SZ98rfwswdUvun6I08gqiiOaflpuuN3w36NLrLTWz/xEP0KrPT/3XCaaT
qR+EvvSZnOaDQkCuUisZUZbhXK5JOLUrBcj12gwHF2phwzIEj6O7gVpoSXIkcsM6
42MW+Z0tkxEL01OvyUdXLTl/UFHMoRq9sgez7Jz6xLYSkeBmOG5uCEpdSl2/dYZk
5iJIVqTuajmmJfgawdXAsTWSetubylqWtdTBD8+EhBmf9jXd08Jc/GxNYfaYwxil
qmTMI7sDc3XPa0eIS0Y2nFc2+d0HR74M4w3l+0ovTBWgteit9MOTLaEn0/f6K/Et
U+2bozP82e3Ko9PFdIEG6obe7BdAClKfvNsPmqTVcnIv86rPozRmOTwercCkQ9fs
d4egYzN9fQxIsj4uzZDfVYQEdPY5P3NFXzBLoSqm/XbFh7aTZRtqNc4nFoE/9vaG
eRTNTjslUtyLvKH1sHgtnC2CtJA11bwdFKivEl2vp21akKa7YFojNkwoam1TiHda
QK9lUEDDfWKcUN/QB3dzzy/g4r6utHvdiGOfbfZMKZNwofLx9z5HAh4zUetfj5Wn
njOvsWa9/N/PR5z35pskGTzHI2E1XtneoWoMgYyqo1yLhPsu8MZOmYxpjr4Y4CdY
9GG1IzE6Nmgg9BA7np9uSr8xJCR3aGXB7ziKLIhXmpU8KzplNzNe9EaafzQVdbKE
av6clXgw3IAb7wU2dzGfigoQXPatOiXiwUwXgfnzX6dXxYH1oPxa8IVQt11DryrY
xCX4rzMqiTYter9TIM1efoqDO9ZZVkT1v0/6I1SEW/afjgkBcAoZqGto6hMpDtaq
D8BbeZqRJrfryO+W2lDrmUCABH0dBJ1/3OaMz8Awn0W/ovYwjUU1bb4AbLqoaB9D
gd4izNLRBzw6teC36SToXXuyDHUYxmfvGuJRhuMuhU7EF3qk99UpTqdKXbebQkPn
g5PZJpEJ4+9JcxkVi2e+B/ABnn9SuQk8SWMrHmxukXre8HpZM7z7kIklOPyiKfO2
XpgXW6VPZIkQ9ljY0V6I9fA9+k6nT58Yyrcx4vs2K240K69c1zmGc8v6BslxyYoe
npHhAXxpVawGGDb2JEUjOr+BPjb+tVrKsCbricaTBvwaX7jSVTCFn+YQnJ/WCD6g
hjPkLVWNVUV4f7WKFsfBPRxHAj85+gAYOWYwYIWJ6JU5GEpa23umgU+ucFTlPfCh
QSeRSm+OoSO5zhTx/Lb2xe3SGXJAjM6kh1dJRAjWr1XcHWcKFHuJpKdw0LebK5MX
Dh3pp6a5yNehsDkesJ6aJMSqLtnLH6i3Bzc/8ZjFv1QBw1B2DlM/6aOQIWlyYRkY
tzaTmwkIkdE2A78No+lsZgsusNP11Lb2Fdl+FOOCY4D9ZsnEABTOFAUkyqxbX8U4
MaLiuW8RaGDfxZsCLguS09IF8bJ8vYesnhtc8vyXeC/RRAtV36M9f12tv7pxtK1K
7TaRAQyX/4r6CTs3BaQIlF3Q96ORChg7OzEo6aDpwZvlVbH01z0zo5uvVbh9Yvct
tMqm36IhfvHT3MMm4+1jrM5VDYoG0yGl5BAJR0J23Pg4vKC+PoYjnydAknsgWdfj
xMlxAdyEtZkwQXbyBUhTmn0pJqtDtNMGZcnU0Hbce/cVVA6Zh1fv5m86BGbFwPqi
/g0Nwfe8slGcDPB16nDwWGosaYyPYYjtjSMXymR7233R1DorHyibT0ICTvO5TIjs
j87kCwBQjyNTmKeNnd4/KtwwgjvPf/8ANl/HJrtCBWXQzdd3nnfgSzRKeTCYe3nG
ABMJpGihhv9MJeF0n+Zhvs76lrbc2M20/1qpDDpfjZbxabhklfMMJMRvXILKVsns
KPVUsnnMQ4QFUPaUrgK3srMmvww796CD1wA/O4atfe8zORt928jChXSGRlDfipKb
KWoKhLl7ItbiI6eQLA9YdKUyF4p0n8IzITtcCxUrbwscKYNwWuxpQSO17zJuS5rZ
hIfHQSpbgYLHsksGsKVPhee1IQowgbsFuzpKaRP53m8HY7ps2+uSDawHQFRw7iPh
FXLgkfEZ4zO4IM44YU1ZOjQ+18A3MV1eOdNEivW6RLMTJUjHXPwZSfOv025gdXoO
lTLz/UL/SrGfD3B/yLO3XaYf14AY1bqaPNdLjF3ONPraydymhbpBuUllae2LwK5e
dCAxfigxUgJUF8oaGWPgHdDlG+mCkrfDjz/0hvqL6dzQC0qg040xdl81Mdu1jmuc
lvcP7/0HH+ZCn0xnreZ0ZSKBhfOyc5GIHLtP9xf+FolmNwznYwXJT12pdV2TgzaA
PhgfGKV79Erp992tDQIpqD5j5x5sELjlX6K6vUsvpKjEzsL4lqor901aueMolRtO
aHVQbDlt14yQTOW7rh448z59yrdYLHqLzOluHSSOF+LGPZ17UCAJVkae9f4vUMoY
fCb0CVkqXUltD3074xbFrngKCkHqUypKSgUpEl+o+31wXXOPtdSKXSJ10OGcE3CK
q5Ls/pcvDC4Q75LLc/1Q5YKz8T63oVIbWHNpYLCVB+iGj6R7wXS5WlOSU3OzNJwp
VKE1MHQAU+CiWTDub19m3dtcNgN5aKJLnpM29Y5bhNOFnhsPLrRLUuOGtJF0gM/+
iP3ZROcvMt7tr7ciWngMQGrpWCN+gwTrNQgsiNl4Ay5sQB1Sa35zfN0fFICqOwvB
8Jq7wUgMp5D/lrQKxw2+z8b/3CK5vQzby4JDwIKMJnuRKtpw+OS/wNP5eQdlQs2Q
RxMRJTtdVRs4mlxSqgomwXAQEz8oBS2e2wB6pS1qdMhGAQg+U0oAIGpA7dtzdRJM
KCvEqGtiXBiWrj7OYzsTGjx17HUfXpC+045yDjuqvgjYArce0Rd7gdPgmdaaMMgC
4uCyANzptkTTdttoyGt0NNHE7RLsCZ/qCtOCcaBwkVmB/KPRqWSmC6s3sTuQ5Ric
9vJFrq7E9FrRiz0jx11zmThPGTgZS5L9tcrgyWvVmGdem58KHea75QqH4tPpdByt
kCwXA+Y+sGbdfM7W7VS+xVyuDkajNI7EsGSwJeRNc3gYGnPWnPuaUAORIwmLUheN
/TpCOGPwQcdAbJVeVHfwxSE1GUfK+rxmpJnrfGYJ7HbcZjCP6k24Eqo0GNZ7oR56
3HlzHTAvvALzbRNnrYzBUoe2UcpNBYpXoev1fszVpMH+fAW7Qniie3IWezkOMc1S
H5fk30PqY5UzZwqPtVxexs1WeJ37GW4rc0z8iUkzs7J4O+DRj6SoDOP34bxFk4BH
32AiHFc+bCy+gqcbOicXR9sl9YDr8v6KWrpkBEWxBLAV++fZQN7Uag5up6wm0naM
4tF4dFKVL8plt5G2ISBbsS5ALlVisQgybqDbsxcfwgYYZfLJVgDWq5rT1Qkls/yw
1Bp8J4EoH+PaFu5Pb+sug33N/3zoFDtOTgfXKH1NuPuxVvoqJlg3NmfbokZeP8b9
bAYOjCY3iNFf4GXKrsIUS4fGj3pxQ25e+dUEJ455P9jvd1yjlWQ3znOH+SXEqh/W
jufwBaBGaIQxVePi+a0O+LoDyPckx6iLdy8JS0Anx2dGMQcjaa67HTJ7vNeCcows
AFDQ6++aU9AQS6RQKdnG8OL/RdFiEIPfOjthTDVgiN8cw9PPADJ9sUjG2Ec2EUCb
TFF/let9bLlKUbpgEqaMwKodcEP4LVpTOFSEoTwU7kyFQzdFU2gd2EKZ151KktmA
4KvsF6qoeN+K9eV4U9QBxZOEg3ENP8NHN8h9qAhomxUoFtLSI8YLnuUbgw7rrlc5
5xh22iSN3Y8tdIEakxeMKaLNttYW14AstzGSbq7I/qOFpS0PuIGqEjTKaWcFOSQr
fwUu2OrhoZN5K5zLTD9YCrv6rvtxwRKyB4qXLRCM/RNIooJV+8F5l1UGya34zbEW
ZqBQZ2eSF1O6GVbADTuRCzncJOM/tVhjvt5CWm6djUVHfHn/KfqE/bFyvsFkUBhs
JIUAc6/zeyfXaaxj1pTfRjEUYL/lg32JFNY+ha/AFMSMP1XTPsxhzDmcys8HQcP9
HBbA0GkUuAZKXR0YTtfMbh/tS36QscNQ41OZcyzxY6X97/znEsyKQ3H8CiVZuOEl
U8Dx9YLCOs/Dh+JkoX43yEp1sxxpcfK+BIlW+mp8DDOiwG0AOdsvR9bhghDKlKg3
7oyf6i3vfoMtC/0xgPPn0IU16SA8eB9HVO4auqq9zVXWU8tCALbOf+UDd0DHI1NN
fBbWVzAdwy2Ry9vTBeyM8ox6VR6vFSlHi+xpiGejQAajvvEsQb3yQhW32F9gtSaZ
mFGoc7l+cRzEHFzlRDiP3VlXU2xztJIM93uN4LR23GKArza9IBEZv5I5He7mIrx+
g7XjGR2AVZQUxRFVxCzvZAiv0iR458vN8Xj6yvWaDROg9SIa7r6xLNMKljTwe9B4
VuxdL2Unb2J+Z9uaWbA65d9bCTpY17gmO1sPPi4DwLZ2XDFC80Qpt0PmrdptZZ2a
el9++pcq7OYy4i1rM3DCwG7aOaqDA3d65bBkRvUadExlNJnOzDCaPx5ecYL9xP5E
erIx9TZPE9TR5ovRub9+4GAUUMvK5adMyl+Jet8fFJ7cMDbEu1yL0FJJpeyMFmfZ
rtxtNLepAPAiD1Q7GwYBe/wJwxj3zCijzDKtAEUMNJ2ObYvk6C2gExUUm2qq9pde
DZM/x0E+uNOmugp7/S5IydsjXgz3izW3Ex028Dy6xaYVts6VjAMQr1dxc6xaPiAw
sZGfxK9eLzVjLmkqknwWTuW5J4sktmGV4E2lH+/X8/swMsep5RixNgfaowhfOtnL
z4nK71VxobPzr8IVfDWN3c8xVTqCqloUENKpa/NC9IoR7b+oIkc1atfH2cqaky7p
amqoQUjS52LYrSfXQABixfkIGK0CIh6fsTVXuYqHqf1lTt7tWwYuDzqPXqJ46hQX
1IR8Qt/rAwUs63P8oRW17VnnneMvhq1xAUbxvbxMzPvM7BF9LFyryokKD/wWFhE4
IJUFkkDwA0bNAHMGKF1RHqkN60/RHz9XmruYbRMM1GultGfUBmV78KaY7sI8PjS6
5DEnuHTdulkQkKuujMCz3ku/G2v5+3ufLhRJITvuU3KxFhPrzk7MZm3BjQbCCaNr
UxZ1+e6fwE9DhSu4JBmKByW4ZsgumL6F8U9JUfhByEeA6R4/QBsQWr5GKRK0Zyq5
fuUTjXXFghlpmud+EPELbyvHKoc92qgi2whPpDOorgdZgx4JU6TgxMlFXW1k8qQ6
CagUpI0dku6CK6gDVciecnX1aMvk5GCp568UhnKHHenDJbv1gsEEdo2eK5iQsigb
MAV7Rz/R/WCfRHvvl3Z2twYGL8GLwAreKn5k9xzTf/m4QEQ2HETA3uiO2ElUNi8p
OAThLSI7BMgGkqR9YRoTu31BC7rCFI3VY5dPs0a605lxVTl7T0DSETsnE2sWP6zT
eBcsNRsbg4hEd4upo8BuiOsQHH4cSCgRn6SYq2uDsFAtoT/zztKymZtJrkomz8YQ
ohYKHRDmi7xZVNxCTbRZbXkt7vYfKtK2ttPX2okJFxTRMFWfEWL/sEXoZ6iCJ7LS
xsyvP7+ZkJKL00Iljn73B/PKWMbB3UiFT9ett3yF4BIsZ3IU1M3pEGKyBfTunmWa
CsMxFjVZlUGKri9f/MR+FuTvIUWRXIY4kln4cmVujV7seKoolpSOvPkzUpa5qW8z
F1UMNPue0jMxDHj5WH5oTzJmAQ3TI4EiboM2B4ltnfA60jQUCC4Exz6rEFErQ0dd
5AxjT/UUs6YtGOXlxHg4jtkJAjuk8d6TUd7TKO+sscFvqA9WVolfd2SeJXNmOSFt
4lYQeVawhszjuCs691x5lIdfNC5fIJKiT9dWjTwDT2/DHuVizSpI2Lkt3Ll8/439
PFf7FaOkTKc1BmKA8XkVXfkJHrZ7mLdoO74NUEr/kfuWejnjfgXKsoB1POzqtjuK
X+TyMOEhTS/bwW1QYfAWBdeb5Ws5iedQeRx4AbVWdCGvTz2aLcITI5c0iWc0g5mb
NcvNQ6ylOycUqFkorH9tbEknZv8YVdo2IyucZ84+KVFOx3zAq5ef9/kNmF4sv2wD
mm3ajLIvHoRrAZCm1tSN443RnPHXFT2VqBSKyCD+kgbSXVg+INjRCdjsUE4GQeRm
Ib7Ig+6c1d/KTus/wTFEi6jg9yyIVXeKm4ur1FNDFdqV0hNyuBEWWYKTOYSe8wep
qX4NM9vf3L8nXHiKNewhzXAnX9YC7T+Pt3ZOvyA6ljyXMruTlv6dkDmy4s7btqeb
A2YafAa6VyDE+3IVS6kQ0CPPHJaUxczJu5I6t6CG3wKLA9RI0gpwo6ZWIOL0SbE/
mY2dtZjg7HSIU3nmoaFE/Du1TkGkghQzDQFuoNQIGrrkoy8gskHbKPmf6zQd8TDP
dx6OW8Uay33gYvWlAFpMQs3PPcLUfSLp3PzkHgzMoSrLyR/16Mls/Hf1WkD+6TId
ZBr2MF9Q8bds0lLiPWxd1Z/7erU9fXZqK/RwNP1BbcplFU/McLK56/CXaM0HbRnR
efh3YQtpJw1rnTcBJgR8mD/tJVu6xf995wefKRuXUpdciR7K7JeGQ04/9g91fWei
guOYJpRicaHoQnopt4HC9110hRzwy3Two4YoFBenp4M9aEaBMtu1yDCG8hEDgqRW
2H180v+EK4vw410iXoalfvvX04UUsTwZiWohw/56FQLF7AnOCE+8g/9KMvjZ4zLw
jiZitxMvdqRggOGvbO/lYqrILWAsIlrX9PapAk7Ke0G/ITVTSENNrT/rJrKdPfz5
r3keuWSK5jfn/HHH450iQ0KaYPNShCzVLyr0XoPBx77x/HrUIHtZl9cGoTR6a8qM
LPlFQ36mBmkYEFWIcmIVb4x+Ns4JPfNGXh3cfJSQTNdjOYNXyA2gn1IWH5etPftA
aB1m/tG/+zXzoZOHBfr5oHBKoF+rqh8PdOWQ3wEVgnuLYO+sUDKHoa2WQPR4ra44
l1u9bqkHHHT2u3wCjks07N9IDnj27dH3Cscm6pWO5z1egM1fwLbq5cImI1Crz8js
4rl1ZDItv25RakuiTucNQ0OAkGP7xi0CaQKa3FM1llrHa8OaFczx2lU+0Xh2y3A0
eyrqBQZSJoJ0vw8vNbLN8uyKZRy3lptqJZ5Up+h1ErHRsN7oRIF9nUeknIW8oVEF
KBqlcrecjndQFjhrYqyzLznYK4aVRzZYRQnLZBkPOHOpVO6Q+Du6mLdh9ZaJdKcH
g7E/SlCiYGbgbEJB3VS3GITgboVSvnPqrY2XbezfR3nss8aMKhv/rW3wPvAjmy4P
OPzV7VWdL9zv0n9yHk+wLUszd4qjLdeuo68qDXc/0bSYkGPsH+4WwEyrweN7vKMK
lfITCG7fImfGtm8UhCa4robkdZafMOlQ5tT1zOiEowyyq19jURZ9DdwwWie995DX
3KC3EGff2w/PdC4Me6wiw7gTTe/DpLp/ySl/D0N23uZMl1HCvPyNm6sbD4Kk50pD
95TlxhrPVhloYEs6XTBBfSMiC9kJRxbdotNg0vFr2wn35cpapM+eo0p/PyBj35wQ
XeQ6bT2FNyt6HVKDQijFZI7Dv1CpZmeS/UL1D45jBvYA9rJ8H5O1k8POC0QucHr/
lmdKDBM/EVyWzu9/hZKaVer0Dr0HIiH6YcqjqpEi5+9BNvtm9OJQAf52xGnKrxjj
ensI6+RCkQP1ob8RKZxw9g1Zc0c6blSRsBPdK+jKZ/OA1Q0JE9l665ip2tmctOih
EQEpJ7fOhhjEPTRbLESycpeQa8Xe8mbguTYdTMSdZjalzVhoV9Bd/RmM8dFd13VP
aQjVMRlZpL/7REPbJZnOWBY5QkolIOyJJ8whmOJs8TjdTO0y24abV29EqDac9RWe
04KR9s519ukTrlPViYb+3CykrHzzXKOFnkBtGk+BotM85dnlrV29ib9R0ftYkbgN
ojjyvjRL8rZ0h45v7QOqZOOPbGtm8dNjExHEcd/ThVSzfn7w9G5LLuoxIDA+Y6zJ
O6MvAwVHs4NXzvzMHTAOFy9NYz14ZgkydyO1SWO9vkAY/OfhQT/I5sQ23OuEdGaF
2m6m6gwKc55Ncl/1CJCAQ34XGz89LeOKcEzCBlnkn1r0vrdeyZu/efeN4nNCXksH
/nwatqhvS0w+GJoImaUw+P2wYBodOGavgeEzdfDjH/Ol6FPSIVi1lM3sBs/vFEiK
p3vODQeQLU3vTRAZ0GB4B351LEz18bogCDIOMJ7Y+cK2hc2M/YhUS1Agf/HGbAQZ
nGKXPMl3KxXZCbVBL/0ybq59qtipggmG4p1ZK8ZpSfQRbFEA8P23UVqVSd6OlnlL
qaZZOA5EugIP/YfA/ZJcDCjr/9oHrmvochOqY4tHqe8Kw2bjdFlPDhjcdrH8sgQn
xF/6F7AxgabLOWnEq1Caq9lHm4BbE8VmfMzpm9Jc7lMQ8pg7/eTRCWe6Zw4mnsVT
AsenJI+lHU9POorEjpMMTNP+/AkxDUDnWVKhBaetP0vufcrON2IVWm7wAb6VBONf
5EnDdzdIkYtN6zNTKX4P8vWwhXnzjpRNH8l/pwMMb8kPsXQEaSOaC0Ln+WdtCgAo
evJd7FZjVz2s8s/jiwqo+HDle13LTSyCjzSc7O+VrKsqwY0RPS/YDJ02wTQPAlWN
0CtMyaCHWnTiG3bs8FHSyiGUXgxF1gwmM3gXveXBG2NwCUWEJt3WjNAZ414ehOpI
EH6hEh/jseJiZXbpqQcaDRH1wQdUX9WVabXH3T2tnWX811W7YtrCb7w6eSASQz+c
1q5VcnItdRsNmhRmVLlEElcTr5SU5zccG7iQy3NOkMCzv1ZgbWWmG+a3+rXfIlPW
2Wa3I9flix5aRUjX+pxMSvXpmX0arlOjHsaaprQ66t0RzZXrDVfhDdc4P+uF2hvW
Nu7preuU4VLPMPNv3kV4fKE32u2YJ6zR1BvsgFG6UO1VZ1xF2SpWEFILyGf1VPE8
hxclmEIIinfj4hDhwVMUCixY7/ViJIWdaz4S1OgTDgTo/q2xXP1Xnkn7DA1Az/ME
SlOfOB/CGdFfp/OgypQdz+pcdPxCVun+YxowGFHRLU3hu9btJJM7PZLbthZzRw+J
CB3ppKXH3u2ec/tZwr0yj4zrM581rmWIGDCfMYMV/Qv7dI7QepIlf2Z+vO0pHtUe
DAI75jZRpKQQ+YmB/3btTE/9nAFLk+TF0WeLJqRLd45Q2EomZlyhZUMB/iVOD5d8
gM3JiQxO2wmze4yw2gz/Ol8xydbWsUd42NoMGD/tSlDGwLakWAClwcYU1TyaQVqM
1L4iSBwOxcsSQW3rXihBDI746CPpBOGsXulOw2EPFF98K9DnLahog/A6Gc6kV8q/
83+XO/TMQkGfLiFuzLhHor4U70Y5SmjnlzHMTLpWyh9WinaFITkNglUtX5aUFBgW
DMVTmLByIi6JenOFO7msDTB0pD0SzVhpV63qCLa4XrkbdLvPxFo5Ks18HVxWgfGx
60y9+2dj86AnFDiEeyoq9f2yCQEa5EE3nUIxMBbIJYnuSoKHB/8yUdvTl2Ea/Df9
NNyZOb1vsFRBa9mJ8WTkrJnYW9D1p8bw8v0r0pA0D6hoR01coOGLSdRiGRpyF6AK
unjAWgABpGZSMJXQvnjI1FcvGiw41TMpxcJrCjoqktDI9vlRqHPRDay8bMCvQiVU
/uO6qCTbV2s1gHpEKraC2ZZyw9PlVYOLAhVpK3DyNxuBVwpTTZF+giVRf9Q4bSP4
Ba6vY3RLE4z2yqaSOrQm8nAv3ulxsY3Rxgk3wDWljn3dXIZsuuH3C+KcMjkQVsGQ
0Cy21vY1BBIZkeGGNyjGaf4gcOow0zC7KLYAV9l/u/AT48z4lSJBC0M4g8jnMf81
9+UU29vTgwUPI1CDdRkUQmRpSXhP17gbofRuRFlSn2V141aQ/LuK3JXyFaybgUsl
bytVKBy0RwSHXIrOClbt5aNHWawcACze5vrVIJjqiNFeha4PhrZvtwLo+Lsz9DJ6
zBHa68iVqMtTGu6zpyIARjdRhdk9PAyaFeO1w6Pa2Whosci5USP72sblwgFxmza0
46LXcwjWgGmmhS2SyqnAph9JimtPBETmWx9hByuVYftn4jVaFxYRr8r8EgRTRuro
Uwqp6g3/YdVOFBmdJ/aRqpCzBktxlRSnw5VlRRXCfNXaFZyoJsg6VUe/7oyoo1WQ
XiN95dRLK/l7c4hS/Y8G82hUrmi0QZYC5peNvihMVb7fLqW7faWT6wq4p3hI6bRK
Bx9FEy8lA13NZoTrylwsK0A/A3JbWBLKy1Z3WHGMMu6VC5If+hfHLbZMRcDcreEs
+e6hVZeNzGVpva2kcAZg5/pCEd8gQ5b6pwiV2VLMRk6N/cQrRXCoiNUuX7+6TWd2
TOebvlkAsUA4huXVxL/NwfzbXZOw/BmWUVqKy7yhBnpDi9PaXmNz8hzVbEmmWNpj
v18jojituObMgK03kWvC8jKQ31WQGedKLdbf0R4+PqXUfYiDS9U0h5Fda5a/eZri
jaxsQahXugL8b3t5Q7HV8kS2sxFsSzuC9tah5U+qa2Bqdcnfc1FsmpndFab4oD9L
aRowbaDo+HHIhRVD1eO/0Mr99oAMLDAWvgsPC+MaZieLutrwT1V+NrJi2xHrAvQf
MY7xrr7r4PiCzZo2wiol+EHcX+jtzz6VP8O2xsOlwbtZHGIgqrzxcU0Kq83FCRFC
KgtxitEu42pOJ356rfampRT9HDQzBHop4mZvGICXvSbJ2sHccqHkJja3LcL8wjY4
/M2aalEDTMSM9ciTdz75YRxaJPIk8EsqjC2KAyzW494B7UA4qV/lCF9XsHg3llpK
3s+NCRbXUcz5elCPROv+AgMUBrfxjfXMyUnI2s38JSz5w1YUfI1h98qoZmUUhauF
ca29+eKCVWRN1Shjr085lEgTvIlEaC6osx0OGFyigDcJvSjXrzDCe5lIkgdHPfAP
1mScnCmvR4VBJv9CepDAx8nUimwuMISm7DvqUuv+sZo7XXcoGaUvVKrPrKbkfTdv
TTBXG8PHDkMU7qrcUOUUH+20KDoOWVn43IcQDfdqPB2Qg3pZq5OD0UA/OlprJxBH
Qsl6GOJ/oiR8KEIfpIrTo5NxK6RFrlq5hruG0181Epbb7rDFerAy0/PUqRE+u+wU
AuZ78Er7evbtirWCvEC+5kOIv6ZdO5ynPxD87cSYVH3H9j5oIf8nHAt3Yx0hPJQ+
GpRcqM9uanHovyTVZuBveVSkREe+A8ed3/IRXeVUZnJkEqbzdK0Wk+twC14Egy05
SvEbEJJzKmPuxBgII0vQqbL0PMrtm/dnnfGK+6IbRzboqumh53KLUJdfeJcUV7Ez
MybXNCliCgEwf30LiIlgph+16COv8G/V0KXVS5vTgqxB2L8YLx06g6Qn2ZJESWjL
GhstWCsH5Lu3k71jUMIv+n7PbCro5lRjJ30KQb4Irw6uK0rTfThgSRgnf8ugeEah
tehJiFtTCbB/kjwl0MEPaPS5RXfcKgH7Cdl88R4pMDnxPU4ZY3zCcesAQkdFSS7U
Q0w7qwSuEoTP51SIxS8Ud4blMjSCXW9So8uXNOeTTHWwVTVFESyOn7apLMYnMqqk
vAWEd/19tcq2u83tHQTt/OZBzMA3NIYXCeiJ3ENdHEzia6+fawFQ9MinMtU1a4Yc
0Jy3EzDYR6DKY/WkOQMe0mxKUAK1rta0/95OcSM7ZJLwh1MHPr6AM09RuQrS0lR1
HgrXvDWL9IpgC6uVx2JKL00LdbGRLyp+CJ6W3Cx5xRWNiKgvRhcGKSysBnzCrtYt
SiseS/a4e7FIcHyRJfSbkAv4IhYKJMHMN9SIo3I/zEKHLHqvTWoXSnvXDpySLNCc
f4ePoEtoIZ37X4c9wWosmmAS1nzgxzCm8tQjoVOr53ynV4R7Ls5UiuIWFXwvSNml
6eM/fYZ6oLvJBttSNfM4HhkLnce+rzdQsTS0MQkrrOEwMfoh/iwzH6UOzeehCTP9
kU8Qwm/zDJx+WxITJH+l+zOP2u3yfnH1j5WYuVtsG32opFCDPJBjPQbihQr3ybfj
4SGBcWp7zl48hKz0IjvIADIYIyfYDxn9GfMcDywR5TE4NTOyTUDZ+oEBkkeNBC3s
lqU+e7rZGHOqE5pqqTpvKxkdghA4atHZ6xn0+eqbf2PX46ZRI40P2R+zGjbiKYrd
3ndVdyjs1hUuQJSZIY/1kxtxiCobR4Au9+4/B6PuEphD51sAtsE6g30x729zqRDO
+logBI37yFmdwyVVtKKHAAcU28oY5kJsKsEDVbot4kTguhJqjSkQIV8nkyRO4dRe
eSQqpQaUul54mIlMQKBCHqFb3QaMOxPc9oXrkbw7TS3nwZiIg5JLHjN20GvCLz6/
VXxEewzLmCKGTDoDs7u3sQsqWNW7/hJ9n6HMOzhlElqzpW0fSAr8PxDlOD0O5ja0
xcAke0le1mdp6ek6GxF7iMYsMkZXO2Y9plRPIA8bjhoi0BzFrsb4/1xtMaz+MRpB
dVeV/1QnDnoGpWCjV/S2bWtTK5LPvGjvqo9nAXx6G8wl8H1S8zmWLVXJHnlMHuKn
KgTkdt3hcRQNGRTrPd8/aTZN7S2/KHnfmmTBvvnh0wM411iCTOhtgwEMwuV5dC7j
8QGsiV4Kb5tvMi8T8BmJLbtYcoVvwSq82wzFiEtx148MyeIH2tkKMOnw9WTDmYe9
1RtbmFEkldeUq8yoh4kWgUuyuuaACvSpQ18yP8lsyYQKr7fHGpAmS/JIUmBmHfHI
JdBMkQPa1gbppsZbTkr5oaHygeUonJLqxfpK+y5Ob+PD5x5fnmbvu/aWG1GDZiZD
ZGEGpWXJAhQzR+N4SSNumvQ2jBttMha4WAqisG2V6+jCXlkRLYqrsPQlKmPArBcG
WnrOggKoEdf/AUH832qcIBVOBeLxBc5ClQtb/dFj2qC/r3PEnpy9v8UyM0m6Kje4
PRQamYVgqSHw7Wicv/RWZuhyxN5tXmxcGnlLje0p3LeUCrOCqHNWG48kOtTK0Dti
+G6VUV0mJYdeQl0MfjXBfwWj3mgFLTm0cjbl9SwRoieAsAYkyG6g8jAfDT0y+ff7
LiU4hTgIFUewKBBV6o0/e4Odo2aNnEd66aAxQL8GHG5UFECqarRljDXnusWXICzs
bapFMeqIb3yp2qo6Ybyw/Ys7Ft+OdBlZqRUUjz0hT9g+FwZNKEVkjOJXkSI9Bmwj
QXY+cwwaw/HIEEh8Drl7F0AElbOYK+XZqscli+/RXLc61a+OxrEhmtOaAyoT0WzZ
wePMQWR6/KybWxG6OdZh6sHUdc3iHfOH2Dq4YeCK/gHHi6HuDOQaVjnmt8SYiOgZ
uI7LdOh7TXi5u8kPx5MjnB1pVQMwkzFwWVGIGgQ5CrIvTY80nq7ZsRXjo8B0hfaQ
f2J/cAabLe4DdvL9R37XTzkcrGfNrj2Jlw1bmO/fV8Gdp4Dj/ILKt8Mep/k8WGVD
7TPkO64KZyVGSNxubnjB+YIYRHSuWLpRPG9HbQrPA11+xc/UvWMzJ3qvBOR5NU/V
fXkeujtuiexnXaK6tqe/F/Nyfh0aLvdAAoQVbKs5fjEuxfgS9zNMUmW4hWqvM3PL
KIinzuhYV5p8MRl2quIZyk480jKCgTOX2am1BVf0tVAF11yYMyNru6IFN5X6Ere5
kyFeOYav3SI+Q3FvUeYEwY+eNDGFjN2etFOUqbsistT/pnL899RgC7XDLyhOjunl
hPuZvdIWiIw93FITOk7KOhU3ImJ1LTo+Z/0dqZOkrwitZzjyjNlnOAf199iuqobL
8xcZJKAvz7q6/jXrHX0xSnh4GYIeCVQIyxHGRiZbcm4QdLvHo+Emk03R2ZJigPXD
Eaj6CgtWfR5YDXSr7mJbKA2OpH+/fViUKLz1DQ5hB01X18Y1btA11/BLg9j7tipO
9/X82pI07qeQt/2ivozOsQf6WJbfJhPjLvt7LmhXV+ARKZmbB8S/It2wlwM1+tgd
yAohT+f3Bes9wwRj3qtnXrSMKstHGwtcJ+m4VRT0yXmYodCC5gJHb6wZ1t3K1WSk
XUtgekrI5ieYh1KjxnvcVHvlS0/ambaAH3lscDixH+bdIHPHj9sSCa69JpWAReoh
vIaUSJOXNOEI5zSNeN8qUqa3lxtxXwxZgvhD4OrPe+GF9WdaZ0fuM9J8qNbGMxcY
Y+igrMFH/Q6pQUempe5wlB+BcNIxqqBQ2Z4gxXYqVh0eJsDNhUjBwCbcztvdrjs1
gd+cOQttOarZnmAD8NEma+ykc0Z8fAy3IxzOgnv2WsUlm20tqdQKpCJ03DhdJjP9
pgtWFV2t/XXLdUzM5iZkSZexB6gr/OuhDK8cXmAEz13s1Wbm8g9CObk33Yg4GKrt
XpHlS4GyINfLoo4nOCUA69ED5lVCUhkBBPmZcICG70NmYfXnFBo35v1WVhCtcnWX
WwpKOW6iaaNpv3ZcIG2PzDi9umOTmtB2tXrDSTA0Zrw55x7MLv8ZclLaPTmiViOd
GRuv7gyzy2M/iC9ejwwRy15F19amBBhVWSGptALV3aMMdi/LFzbjjXzc0A5iNLA2
RkgTcC1qdSAc4Pzf/YcAgS13IrMUVKlBWfVshRuxhxd8zUqNFNpCqxJQk8D90goi
QiP8xk+RVRQlxQ+M2/VrlhJ8oUbTgcYZY1yhjrJ+OHCkrxK0s+ORYy2jQw3HsF6C
j3I0LB+Ct+TNONXRs0j1ss/QIiho61TfUePBwwXTnvFhy6ER9CwYRXNQetSuzxZi
zBcoEJAjPHmR1EOaPn5enwKYbeYfV45jprp+rgpUcbkKP3ap4VF57uGPhC38OwFN
gUv6w4EWFZuf8P7BkmcCwMCvfe+75IS8sU6JdjVeq1T7t/ZbjvnH+Ee+y5H3HTlL
rSq9gKSGDhKAHK+vKlm9ruH1CpyX/8Hiijg/637ZTj1iZ0K6EnKEDx2g207E6Gk1
FnyjB9FciQJMfDjDwFKTX+67cidKQtuv+P9G4ivNL3E14Hi9hgIaTBHgleSXjbUa
AERbaS8RZqDuETuxtKjQ+LCSeX+vqteMkPeo5H3qB1sOkzqGXBjckyn5AG4Z5Pr8
1cYujhkD+KJr/FKfoz9JcD8e7HYneDBAlWAdQcjc5plqTKyS801b38y90sfHuGmm
jJADiFkFVKq7cbvOpDf1qQascPs87Z5g9Nbx476hMNhbOROOJGicPfC9V/Kzd5gb
XEa7pUeTCqUp8vvLWq5G/S3csCKeYzzUvJNi6rQJ0b43nMLYf77XwtAPunVbbwus
sti6Yka8H58jBk6Z2gybPq3DiXIECFkSMfedlq/P6M0cChz+kQJ+vIDw+hDUQF/6
7z39uLc6FRUO151dk1H8/raHlTuL5A9MI5z5nWk4nOKvFKMPp4Jyi+32YR9Ul+B6
kAdFqXwNeQS8OBZZBFKu+v/OBMS8q4NO5MbrVIGzEcDR2GwDDP23gbwuKBJszH9/
6DWTxQlRcpIoqxYcj9LBM439XTAiEayxOAOgg7zBV2I/wyJNN3fb85gzPEZb9yTL
0GAuKz5Z6uYP8EOaOkKAacDiGL1V3ljkjTwYF1kdLRPcCZmpb2v3OG0weIf99Gnb
xnRoHrV1cEEWQZgXAKe0m2boiSsbUYNaMHAYvIZUDv+VufNTI0j3v8gqu+74OEfS
pv8gpTs7MH7eQOXXuaGtApBeexCmFkSQT2K3aHFEADsz66wkzC82R3cPoEoXN09E
w+OQENPKBleDzJa0KeWLxDrhWbzeI6GEzRZOpCaTT0aGpUjrGvJQRTM9sMq5FT9i
GEMTFDHzaTwdgq1yZ1uxSyfeHMXxDdUnUKIZSJzm0uZAiFw4JkAUQJSPGP8NdIGM
evjvjmH1w5RJTP0Iy7R2fHK2yXTcjyqJODKmlLYpxR2bty6pTLWPNh1grCBmQ2LB
liOsmqM2OGHHDwr97Z/B/0dJhgxLcCT/CZYTKML5TkwoaDULb4tkLVNdd5V4Ccit
Zd2uzMR+R5KFjqhY/UeXwZaLjLaLrMewIpfddiybWIjxAr03V0hp+cEJgX0zsWj0
NghfeYiXCNfgBF3/LGCB/UxEew6v4QHEivXz3tpH6QuSRQhNNM3XjBfdk7JIdRzy
o3FUnYsl70HPSlpD81pCVLBjNRWSXcQuGGsR58JiI1rBrfCJE7mGpBYSK2I3PBZf
1m8fJ8BbwX4yxSNHbaR19WQvqRt42ucXbjPVGW3Mjl4J/NfmnoE49jJ3SxT6EA3w
dOVobDnAHea0ooRzH+KQTVCUjlVYxqbstRAqGJI3JFedH83Kh1nI/8640rBDJ3Sx
6XDbhIbv71Ix9/g6ghp3M0bCvnvxUzgZMJIXdsc1/OrwHheba8h87LFNQoCDUtyW
Wt2gWo9DZIgLfqxxI9ryyOGcRx+UuYwFc9usxoldjnV8CYGaxy8Rz/tflT7demwi
IgRTjWia/B1FwI9P1nLxcNxOX6HkxqbimgdtsG/KWF43YdY3K2tJfOT7MV7Mr9Gy
Wh2gqod/DSJj0a1RFOJApnakibpxGro27aPSnfnnj/yqSQNVLwu3aFRjjEIKgahc
B8ym7ZEPKvmooIex0aKzLea50J4S0IkZNZJd/xOXwUl64fcJlX1O/MpzePFWIHPC
wvFPqIaEZhSNRbMLkrLuB4qOtmj34Urg9FVnzfhLRyGtBIeCamxT629SCyf2upb/
H+pfoOGyneEQDtrlpJFi484Y3uljD0+yGJymyc1CfYYTIKu3TqMyU+sUOWRcP92z
LUrOznpq3skVvkHJpk88fE9lqT7qyG/GE2INKzf+weyoIAzO85Ww/8wtpkFrAVhr
QNyEmFkIXAht1w0UiO7NF20iPFAqIKYolgfk2TEfhrLRNEEw12vQW/ZhD1UkVgRD
AY0neOHDLYCF/teR8rPX7uv2YuNj5MusU/giTmAAnoEvhKL98g5Gsfw7ZvYVrdsn
+yRZrU3dJpHQbHSooJWOAuppNcx7UWQ6fQSZKpJWpNFV2mBZ+Fk9ZM0wEU3XSNQc
avzXm2q8LtI9xlHt9s/Vd4q6WfzhKyXgPV+DWGG43w9CSbxkRIbK301LlrXjFUd3
oaYejqwRlkhldwhl2MxAiUeML/KtcBQH67IRE9edhhkSu6DC6moJK6x3ATNiwctG
nLrhfa+OaFn73W69E7DHDNvwEj25+CsfFMBPN3P0uxCNXRoPR0CRj6v8POzZ1OdM
2aMa5HvlOom2OvvAk05H0e4tMQ9s9eJp/oDCAcNsmCOknG8hsPB/jqxRguOOMaOo
Y8Z88DWUv3RQqPYwJTDeHMn45j3OiKw2fBG+A8dsatyXCfars0+gsoxVyXPspG1i
cj0Yeq0NuzxgmxYYjulc5+NthcbFo7dagmJQ3etbeI2VY3kD8p+Ft3PESHDg+yBH
G4Z2nl0vfmFCzRHsKdQKfe+YqGeHKkZPaxkKod0/PQPZ+vxDSPalGc4tGNDNj7Yc
NVKqaOHPUErVqB+ovMOSIpSo5Xr6WRO9Y71AvA/euvprACC89yMj/RHSOzFTHqOj
xbz33wRgKz7uekjA57z/hYbxJ2B/ksPAUXFEpVnn/s1ffi/ioASL/Z+Ov8jKRieX
OnQvaTNl979XHbbg8F0zJH13FkeEk/+zHIiB8WuzduGFIAWtAjrs/F0h77be5Mfy
cvNHhAOXoS0IYoumsFujGrvV4TXZ5GxspeFOtBYbeWuXnItcQXJSLEcF4/glv4et
i7qJr2WhMTbvr3zRLD2z2jYA11iZ0fFiaQFQ7SrqYEZ96iYEQahi8uE3NkpCm1Vj
OtHrcm3nfJJN+NzAgpQ4KyxTbTL38oNaoIFIFG5HmzwzWITVhejrbrbYzdwkpyCQ
k/iw8OcJESaQpV5PU2U2d6DZxOJB1NH1mBYEYO0giy4TKOJeXfKhdHj83nNJrJKJ
sM01B84KDoeYNYvZCnZ+CYQjX1W0Z3GAkZORi16COge4uvgWVCDA1fyd7dqIYhcB
jdJWVyirN335aOJ/3FfiBCiYpHfA1bWzN7mMAJf3MwcVuYJ8a46Zroj5ShcBPCDC
gvXumlZK4IVQ1tLMelm/lX2QnTiwCjEGHpu5AEfsGjO5pjfY4AFZR/VeQoh2pDHX
AtAY7rHcdiKCvON1wSCxtwNmbIKx5PAUr5bOGP8EKmaJXTMOdCibO/TaoY/ePkGC
lyxDqr/SiyEn2qnGOLEecgArlgdT2HDDJTRU0cKvOnsY7ZZ9E8I42vZnQRJ3fadp
tWY091C9jvBABFzPuAqURjwNA6CueNzU15JrZODI5qHTTp97OtRa4S+2akrnA33k
sDpMtSyfpTjXZ7SsbxR+QU29Gyx77qkA31xOq7XpsNhRRliJH3ccn2dCg3uJkapS
BeJQ60FOpaypXRotRgkLojp/sEzJtBo/fR37E9F2a9g6w9BuMlLPuZZTSt8ql5MM
xX4Ac4vg5e3uO4jKb+T51X7ohh6RgunToSnK9SsE6V1TjRPQt/hX57CUBgZzP/+Z
gwvWZiqwoSfA9u3ubr8P1GAce+VhYt1T386ixmGZ+a7G3GcEH47krPYHJaNfnvFf
4wxgAUa8Bbwfe23OxDbfRtuRyDs/NfPMWGDkRmqCujtuopuniioE0SSuNBTn1MiV
v/c91Vc01Cv8cMj8SwlPK2nejWxt6NnPJ8VXaE7OSW6sLzox1H0L48lSJKYC5VAJ
WsgiDO6/Y65jfEn1jJfVDLbFdVX+QzaUsLTBJXlVdt5Vy5eqH4dbLNTXrgv2PZx9
7iw1Bjtpi1q37QY6QdIRh1LuZvgROT2waPkYjtIqiHcKaFiUA+0z9noIarND21gZ
izNnSJxx2Xp9NgZYpsQK3BxZB7+cgWbcrZmmReJfMNz5E5wqAp1D+NsSuVOAUCw8
zVddaKBpoNTSMdLKg4Gakn+AsiWvXPqEsEWCmyEzGsLMsEFiiOtkBjyB6Eg/hpJs
EXAxHxE50xYdNiOplckZxFlnSwritzrUkU6pUx9vLVdzOaKn+9GJChI3dEtxX2Oq
/o3b6e3qMhExvky141IxnI4tadizSmScMV9rgP+R9ZpkQQdcdFDVV3Ar6VZTHUhL
oNAuoZKAE17PhdS3ztm6Qvbj+vRn34yflhh92QbQ/ZB6zHemPlujOGXi7ekd0377
yXZ9kWoDtH7DOWU5XlTPkamreGeVoelOPphWwMCzhyNvE0x81lCXj4kjuRYmjBOO
2ujhO37+lIYyZFl1Fdhrj6NZBGuhCMzVghT3iFsGKuwd09hootlnts94wFWikFiC
Zxy+Li9q2qWeNJ5QSJ3a++rfK0817YRee8MELD3herTDT1+569sDmgzsrd/lSv28
KNyR/A+ZmxWqHU9vFuBSON1EaWqitVQNP7D6/UBQ06fD3lrXWufhH+rodHvNIVlp
qw4otY0pCkcPmqeyaVdE/y29zJVuHdKEdhHI2GDIt42OlGDZd2mtFLDGO5HQrX8q
waCboNJ/wZEiFehIgZmf2KlvZmSjFYdEGrdJI8nI85vWWL/ZRAHDGOb/iRqu7Buy
8x5ircgBQ8hIauUSyTWr8oTcJTxExmT2t2JRsz8E9OZgSNLtCLYLDQ6j4lY+uUvb
NiLdseo61rNrUXep5mdNPmQCIojQTc1h+eetc3tTexiJPzSN4xDhqgb5lw/5y9GK
K7Lff/96i3PNq4RlnKdnjS/vWrRlhJkQ36ZSkKbWd1ktTY3zvMEvTOPfoWD9UxPC
5IdeOB6D3yL4dKSbqlZJReHFeOus3wYEEEZ5Br2bWJSSgrtjpEKT61yidi304wR6
6PPaxc2R4SONybJRsAc9NaZm3doghvJ/pVHV6Xk2m5XSGImfUIPRpGdqs9vpCsxI
D3xmiCWAkV6kRryauWBb0BVms6iAam+6hP1HNAMQB8xPZTvyg1Q3SGiAKPxxS6+8
t+urYP8gL5O0fz6tjVglW8p3fWR6gBQODYSWO+DGuNWLJYW7uC7dRNaMydy7A3+v
qecXbGxAYZVbLxDUdJn2WLpf3WUEFnnHedjTjTk0z0GaAxci93IjK1WukMz69vXA
X6ivm/g9BXOGRtCnT2hg+JUq1gSC57WJkMGtifXBbrD0GwjvIJ2euylA7POHCcdQ
iDLu7bX0KAidi5lnoeP2OkEUH1lkkQG9GOcw1LqmkqMZBWqCc5RdzN7QTUWykeYZ
KlLvb0MXNZAAY1e9iHDfoFfEu9mhrK8nA4M7eDo8nFTJOdxYmSIN2NeYEhES3mDn
7hGv7it61LDQa6Kxsz4rzoTzBOfy8Ku++maEAbocoMXmOwMHeD60wD8xWG1AjDCX
BrhcWJVN9//QYndezDbQdo4Ek4BHk8Ml655HMMedZJYS7H5DIReJnjhmT6bYnpmj
tqpZSfvVtXLKd6uNhOqP/gqoyi8Nzfjzv3mlmgJuuulCuNNf6BvDlaKDH+oOhzHk
tSkQaYSto5YrOzmyrOmz9E86U6pmHTGW0knxPP59Iy5e1g9Vf1s3DjNtFKBghOlR
UsSJoI6WJ3E+D8ph69olcyMbvpAK9NE7bJ8MtnfBlumXDt5wrJ+ifczPaKRdvb9C
b3mQrRunJlDF3en4Nh/mlTIgXWXpqstuEKGQR4cYbHywZ0khszJyLhUbaZgotDeD
69Lq94N3VO4h7yWRB+NXGpX0pI1RR1BOGd0wugIKaZ+5JrPHd1DDxyht4sPkvqGG
buv4CURFtrDdllARqRebIvm+DpVmG8L+7vNhAnfC+s7IoFiPFUUYcoFTQTXVtR6K
rfqZHQAvs+/BcKwYxYWJl9+aksOcJzNfWXNIWzTRPIDKFY48qEDSJEeFK6NGMCoH
ShwlakklqU+sPoz+9L0QgYmrlaIsdgG+HEDubMaa6LRzFlne09PnA9CUm0mJjTDX
KaRMkTVtIJ19MEu1yigT5YZDpeAMYMg05k1m7LaptMgS69nRMWElBB6Xcx3JPvLK
oHzqW4rXfT3pDDNaQp4vbM9an2gkhFUg+yYcsGvoFqn0naCVlEyKXr4LZD2Cn8qr
oFJeIHaXmZdTHsPx2+FeWk7/uv293ltLsLTYwiLu/BAxm5nqeio/FtDMltBkZlRS
l+HsP6A0fNwB2u/PDLTYxH53M/Qshuo4TsM3o63SOZCc/e4KdBhBtqpa8CczPZOu
223KxvFNsfp/IoCWJl4xgQALgfr3khU1oiUrdol/TuquJB+5byvHQUpf7vOXQ3QQ
tbJrzJyNLES2n0V1glP1JfTHDaQXoUncqKndihBgHXlavEhnsjImWiq6GKPzFH9X
BtsU3vVEVgqS4ia8qSUv56WYjGqupiIAv1yyks+GCY3wKrVHT9nkQrQufQEh6rwT
ZYAVTXpWFVX/TWLj/KO/Aex/qFnuyZzKZgvQ+kpnXMCLuVO8W+5OHg+o29y+0URS
fEVHRjCnR/Y0KWyLYXkd4pOZscEQfo8e2hWz5TiJjth6lPHuJsdH1F8mXQil5XrT
3DDMi5SyeJTt7ZCgNNX+TsvADd+tNw13FMxZBCztfWgd1QcaS1r/IF3NvZQ+AhNn
Au7GaRdsRa9mVqmJKHXL/p73/hQhY1sm5UjhMgzs8nt6HkGtczOhSYI2Y0tj1PWD
HB/GIIvoE4POMPYfvZi1gfL3tux12ILqMQTxi6f4qP/9ez5SuQ6UNNWoZyN4ZReA
kaepIL2vIfhFKNebbQPgPvAGlBLh/SW/MaKKlYj44gd2pzsvltpWSWgdgQ/8RkPv
m1G2w3jSKBZE2PPbifXYoUiUsm/Hh6JRDGj+2vqYoteLYxhRZZmhKtugHoAeQ3YP
W+KCG/0mqhyAYqDcQjhM6DsseETKztJFirwqdVyDoy3CDt3TJzVBA8EduwKcLwvu
RchbR3NCJiv/FjfDQkk5G52zc+Ph9w7UOWNZkcdYdVxEkEK3fay3/YAIKvf51laQ
CugP1cwZujJaS5Ymke0NuXEex3tEY4QxVKp2a6qoPI/QTUPeOlh+CATd6fVCE0CB
kyJRJyImhfe7ulZUmC2FkPXlWsBn7veJt40sOxhmQgOCBgdUm62TDM7go9jJ4tXL
rwsl33/x3RXdGwqdVEac/KPVZ8AqI72MSNwK2KfuupDbMMZom3BPEE9JEjfoI9WY
QteVZ5tKqidAvFy2kkHtDxm2wGqIwXNeQVIuXw2L13nfaFb2M4zkjUQ0pENOCCzR
09DR9gGmuaTTT+D9i1hLt1o62cvE+te+o3V8I5ItsKp+VMrepXnlW19TBW5xuBiv
nZgB7hbqXAjQLC2dQdRd7w7iWRJMI+sGuDGu4roEEN0JRqE8uj37u5DP2DX9K3wx
IcoGj7SBHrA5YSkS3zO03kPKw7PJtvd1uyW29DWxHrUi2dKi22XHD70Ei68hf9BZ
nD0CPNqehRgnO46EUdsEV0k8O9NCnw7LTFAJn949qD2EDCvGlXkl9lz7qM/INEY7
ISWIpgDidkG+o4Ya9tG/r9vLRVdKEZlMgeGO7IRTKTUHvop4INuJVUESDQPRzklh
Hd/IQZmnPAOfMVo6CP+exaU3q1kHzd/nY7vpURVyuFFvgpTZdymHftXF+yIeoDOU
1vdl4TQrbfo6WRif/iJtGkY5quxODmkksvFqnCOsIpK3T0NB+lk3ImM/MXlbcWT6
K7EiOPKfqhmOMDLHfyb+EN4s36T4wUSeYbzdF4brAk1GuyDBOvJLEqphmduUccZY
Mz4jDZRmXKmt9NjOYz7cPqrqjqEyS7p4wD7rXAwZ+nd6tDmjiL3d6zBc2hLzAuMy
j/Ku9RQsf4p4UizWR52D9EbHrY4Kbs3hcLglUlN9k2/df3VxDkecWT4PxQ6MATiS
VWdm9nAVpVpZWtjcepTbAfd3QCFYSc8G415xhHv9HaWch0n+2sAp+up2nHewbZiW
/ljuaCY2PApKNsmsbvZlnIfZOIutDewfHy8KbpiOk9PtxxDl1/TiEWG5DO0Ia+nX
gPVwF/Nu9VQw5Q08hdFyhiFlZLjai6lbYpoKGTK7ld1MrIZJxboGqDxdf+nKYMtO
u6U9ZLJkitIFsdVG/LWFUbJKUewHNoHR9sqAyaOur0jzf9msjuJvcxmuMQ0MfqSB
Td9egHtslRIOjW9pQu2L4bZynNCb7d2KISHU9D/S/VH4IfhEztu2OTt2QtQcyPEb
kjk9mMqEB4tpU5fV0+nUlCRBJbAPhhGY2x9giOWSV0l6WH6e1ncrKSdGU2s5+euk
G6YVmdWbaCAQcW62YPerOndfokikoNyzXrqwEaibY/tWtEGHWGopgvz2Vy/ZS7SI
hSNGPuxTlvmYChheiCfqdaUKyQevt7cW5Z2DyiJ3tHhHI9ScJLadC2n3shmyo+aO
QyNRksZOaJpM+dWWTgCQBzbWgqViHE7+B6DASsD/Yl6vV5q765b5Hx+td8MR6AoY
SOIRl1ft4tdkmYfUbq5RCPb2CyKPrLASlncOewHiFBR7AabEAEiqu/11JSpKBe5k
GtEQyOMiN+dMYcEziORCIz5I0gFcLNLEj3EfWsVNJOeNDPjDqq2h99X6ov3ncl26
4280Flba6aybCmxuFz7DT2Mjs6mZ9YXuuXCfWxGmBCOKioDxBviyx+ho0VStawMX
FEkOeeKGqVuhJa8B5pyczWQd7oPrKhxGddy0Bt6A6fpJBheGNXrNegRrmQOcBGDS
wNqNSNKhPhGdIhDvGIS9LTkMclvn+b8kf35IYBa5XI0W5WU6IN7xaPIOx9U+R/iw
UvXs6EHQ2w94CN2aroWby3TgdS/E2lwh3rJpVCx2ZF5OFMxw0SwmlSqf076uz8kL
RrDxMZkawbP2Xi1OzfHrMrmAG3A5m/e5ITYM/WFXWpN9eWExP0J5x91AMqSxDuiT
+AxvC39llWO2Pjx3TgEFBlLERmIQLVVFw3s+0pCUibbmAECslIh/7Zn9Yv/dKP6y
zWwN5IiQhMzx2QKK82DIqT0IPuZhFk/74b+QkNYf1z2y1nrocCf7YpXcI7V5OvmQ
4KSC+VVbGJ9ohLtVvmg5V2ReaagtfuaUdfuwOgdL5oUggywpn3Ciqmcb058R9Pu9
7gRgAcrxGfHaOTdJyEDZegssccjCDAelcW1Qo2YfIt20zVTmOXBG1ZiOo/En2POv
FtV3UIEEMSxT/CzxYP/v5XJvLVGBf05vVtA2/y8qMJfFrqpViFHyD22l82MG4qww
IiURQoY30KLHverow0ovG7r6QR+yi5iPvZwV8k/onggXPVSWpEHKcfRGJLAV078c
CHSCyZKoKd0bf3uV5GKuQrRP0EtrXiktj+k7ZOy9bC7u0jODrbO8Yq5z+TYdbsCc
yz8Pz/Z56OuYKgwz39tNDWvEsXVJ0VCvMziWVAu55UYm39ossd7fkfIVJlf86UCV
wfbNr6oK/L5F22OmrCFIHjweMtm8e6cciBz9d6lofwYA4M3uaIpl2+xev0O7ot5D
Drkri7b0t+UVKQaCk3A89GzlWNKhkQglYm2ciF5qYIkFDVQm70696R8nkr51pawh
A5fC0NPAizjdsB042OryCh01N2JJYzTiGSwajpLhVhM/iH4mnO1YH+vjzcwAmf4y
oeZXc0xVpO/4+hMD9L5D9qw84BGGz6g2wyu7sUrpqLFsOySSs19MkIBkG3Q21IFF
zkEHeVA//f/oIdTDfZ1X/OKwYhfPHBLXkhPgnOgGkjk+vWns0JrIQ2WBbdtD4s4W
0CWrrMIU5+OLK2zkcYkg+W1AipczvBdawKW2LUVANykwzOltQpYpN1cNBhJfH85O
8E/TTUufqVxA5A3v/hAyGnh3wTk807dYWXKYZ6LaSfgF6mFg4DYpt/JdNvuPjhqg
r93wotw3y6B/zwYrEXSls6sEV0WP7faIAfg1WHhRzl9XXIK5BcR95AzeJv6RtKCk
Z7haeEDVjWpQidpeqSvz1552m+qGJkEeKwPKTJxHoiFgheZYOfwEVEntDO54mGPb
V0zk1i6jODSY58Ew4RbPJBxn3AsNSBvhX/w5wZlZLA3OeNWKeddzPY3bVjWmloeg
ERS6GW0HqsMowYFJrafJZrZPe/uAlMVszKpFN8JQW8DSktiA/C+ZU6/QsF+erjIw
QcBZATkrHgGZqLIqZWFwbg==
`pragma protect end_protected
