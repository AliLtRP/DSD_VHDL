// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qg34mViCf379P6FknEFuCPNc4haUWVvxe9kIKjKIwvHLFs9nOhRnnelAuASLN9X18KERDpo77RcZ
h3QBzdWbyJZakktPqsub2qfe3k7E58HFt5eyddPbyS7BK5tSovc6Nb8SevlhFy8qy9Rs0or4Kz4e
xt7AvEtd0DSr8nPxjhoySlzis9MmXqRmAI4I1iYuzWOHDF50XAWGWB7bk2m33VOxR02dePPsagzY
zwJLNwNE496fbnDvHbwm6NcUtv4Co9B6gsQw1W741+9YGheRtdSNWR2C9BabwGVfIhXzP120RMVp
oe5CnxndpWa5c8qjOs8KG3eqqo27pxeIc8LCQg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
LzEBjmjdkxM0oP17/u/HQZep8djbV1G1px83wUHHx1WcJbHL/JTAXVDUbpLlpUpB5p5iohPwuuCD
4/M9y1ps2/0Wcy+uFnxaYoOuGHpSzFP/9HapYZ236VihLNpibk9LvZxe2r1NEBIzz/ax4xeF3blN
DW59IknUXSlJ4q4gcJ7oXWPZl/mb7C2DeZ+MG19HmPTugM6Vs7yrJ2pek96ehIgSUzFGgdhn1Yqz
Xzgu24Riz7kqRVMxp1DJxC9LMznjIXC+G1HvL5pOohB07LTDosO9AgTEQ0zLEuGEedeN7SoOjM7j
FP2eV70JIukKiUQe+XB4vqyYXNlgyjkSeVpkVJSNeZPiZxjrEG+ScFDidaMD1ITjHY+0D9YOOSFJ
mUxO7ftFj4LO55HZ70o6Ks/CJQlWvQW0DxTv/BcsN+OQ8rH7mkU/soePOtze6i+SqMazg0GjKCnL
Zlxe8pa/KyhUkkDSXnZGeODV58kQAse22s/bKjb7yBq5PmcExgSq+4N6bR/SWXOxWjM5QxWo6ofi
BRPkbXkAhms5tdNTsQx61zTj0vEV9SFz0jXVXE8N/WrqCG23P2vDUFUjLxFbYCMSTH0zb94Ol0c1
pRBEfsKpwIK8Zn74Awgn07iiAvzveY78s4+ttY6aRMyLyn0b7VKA4dZSIrPrUSR4jxhimNgTLIhZ
xAWAx49lSKoZAw3MORpq4Si7XiyNuMlzMVnmLVosJ1+Wpjrvl6v4q9apxQUXJHBw5V60ydfpoBwO
ntfzV9xKyG6OuB7qBK3pPaLt3f9a9/UakSEBnechnXBr9F+2b7A7usToJKrS+6YTFBblU+ryyHyc
9gyVjcQ2gPIGMq4AO2o26TB5lDp0Xq7flIYdePzwJ9FSfPNdjR+7rEJGNvbDkHGyI5jzAt95tLEP
IJObM/CLPELMgBcZzFbHBd+tupAo5lOuZPgmMAHyIEdJLOMumqiG8zdqNBgQ+s7uji2lttBV8X+R
YAGHq3rt4L/R5nTiiSEfW75JB/uCKZ6Gsa+zPstsfLfnmPEQJ6jfHZ4mHMgHnLNIMUKdvHGrCB1P
LvUo+9ViJMVfD3p3OcEVh5abEfhRc6lDVZ23ErSGS6zorgL8AUh7S4gaU7OG0Sx66gGF/NB94KGm
wV6vrufxJAHIku53ic00TCUNXl6V7QJTp3XI9X1BuqjfBWO2FouIHt3BxyapAHSVxqqdk955tG6I
cvAaCsE/dGtrlYlpLN7xR7ZZTVbNlpUhmyytrKQzSLAQ/m777WG8YIyB/HVlejl590vlD41fUZi5
WyCPQSQryfktDk6TVFnV4D6jHD4Zb4XSTv5BsTznRiCJEZ12HglTSgHmpas13CS6uxkcMfu049N8
XYqZuCXyEzJGaKstP60EUD8r6ns3+oG8tavZHxT1dpP4oF7s5wr09mheKnvw8Tos43aV2wTZn2nq
WguoAWr2f4Gt9P5htueE5p3+hOC8QXb98WVMSJLxTjXmfAX/k469D6QQDjRtrSiWmZv2Y8P2k+Uf
mesrEi1kMNouuZ6VjzV8cfK5j4tfq+ZOGJ3C6LCjFvFiBtbKbuu8H+UpOc08P8F3fB3ceaz5iAbL
9kkVG00TvynfLVCXC0LgYMSyPSaOPMmvSJ618RzfX63L4K7SC79VA1pWEf8k+4JsjVJjvm8PSU0M
Z/69qCOd3kZ79FmeUl0UG2fDtGEAS5iAQhDT8oO1gAfeCiCDudng0MbO23cmwCZOrfJaczkkoi6J
YE7mjYGeelhoiXezYOp9Nlka1PkwwYbmB5ENR71jzIydsLnTaVb1tY+ucuftAB+VSY5qGVU0wrNY
M/O1SxJPkbcTnCphHwrxYlWbisu5JRFtXSm1Zn9+x2hX3+L44cCXx0zINBjgTJzagglu5XlDaKIU
Sx6GodIYzdFNYpaou73DFrzaHBhAfYERZmLjYwHqfUie5b7mBun4t84xgeLvnd+HZdZDCF2cObwZ
MLn9T+5KwXRQiByWzLWPat25/yTCy29GCbiCfm6CNHW0zkerXdJXtUT4Yu8PXwUL/6+233fVPvza
ovTIhtzZpQz5bCSR2lnQvdAYMQyYqd6Re1ODSKUYHK7T0H8QfxorA4C6lFS0Z7xfPcNQOYrGguJo
YuD/Hzvt+kVnHusSNlFlmYxpXzvYq9qBdhnwf3OXRLDgE5LPDhzyFHy5OUOIlU1oxz86cQR4k3uF
zwbwEmt387eUjFHOQGYIb+WZR57SNPSjN63knxv4QEekc26OrNQsODfWEGKcv3096hv+BfvlOA52
hhSOlph8O15AZoiuB0l5RoIHO4zhEgNt5qSy1vv3qsJAi/Rxghg9I6/8hAyYrb0P5DLpALQjPBG+
3A7CcVdsay019msuBsaJSxSLW4eyhjYLN78LgTzXCAE1L3nxZ+gBXQM6kQVWYE4mM+MrEDywm08q
QxjuvD3986fizznovezMBTBHHXSP+Bip93U1XVCM+RMxY1MQYKOuVlkheClwgpRQhrrPlPmSFAj5
deSXjySbwy6bpRxWrc7hx0iQXTCjCZJA2r14kFjkhA7MJB3sDsvJSTHWnBzherTPTmAcy0IqEtmc
1cBr3DaVcoK+37iS6vnhbAO0Q8znzITeFA/nSnn1DmQYP/HO0R9avRCUWcXSI6yjecPJbxJ///xx
Sx2Dmdeaylfz44A4TFg83VyWF9+oQnGiq5XS98YUAuNN5uMipSHwgqurmi/XggYjjPVflqyL3JHs
okvTXbkkfre50Fbid0vlpVr2g1wM4sxLWRLs7kAe9l55rAcN4fMwxtnh12z39CfzX4DyQworpdRX
KZ9w7oJVEicmwaKE0qOCgF1Heb0lYFn16vUgrKHCk04Cl5KUtzCW3h9hdx9nvHs640g+BK+KBMw5
PXIlie9NATX40werd9ObyofEPMMvAsGMS13Jk65n0vLg6WGNJvwYyHTqeTHFWe52yw57uyNpkRHs
CfWSv63YnUw+jkISI7iROpSlQpnRw5GLc9ZGDInxqKU60GTU8bgOdX4agi0KxgCGBOXy5wHi9g3e
fFMNW7Sl84g+A2BztONXkBxsa2t42fVvj68DS0EU9RFmSAY1WuMrVRbLoBwfp0mk0QwSPL3Rl2xb
n6LwSxeXh6GwghHVF5Ar76un+I5KnfjSUvjV8d5gVxPd4W/CoqeOSuH/YjnEQswVKZvhj3TfSDMC
WP/h5ysZ9dJKdVs7vU9/bPmHugIgUgMJCwsNzGUoY/Ml7bODWo/5/OXHBS0HdUtkqn1nT4S88DKT
8pWY4Lt5TN+atv3ObjJJcg7KqZF72TmuKQUjuXzt/g+VgLZa/ig7qbmnXMjuru9jOtFy5Eg1oxr/
jEfr8DYUT+X3eiksYD8ZjnWebM/c53EnF6bYbBsdUqPQUg01Fd1JcKPsjUPzkhbQcjhhZl52XodK
v6+TVUqv83BtSX8aJ41IrpxHTfiOdYYdidIyFD6ve2gL7EQ95FZRQdZKZhw+Qp97cVwyEHW3/KGU
tP8b3C4mbObBLEWMj2QAGwlDJ6B1SSu+dyLPN7VrB0EDWTz/9Fcn+ptaXQMThm04Nf9iU/zTYpw8
q9JxzFJAB4n7FHV/jgg8z3hEHRYC+r/6mHPO8ezj+AkvUifgvu0CeYKb87eLqGXSNOxdVRQphuRE
Mwti25qBecpcWHVpV4EAHKEvujP8b7hPaMZXUYpIon9VIjEL9uinWH/zRKshN8v4UvUkLdJn+LxX
k2IOvkYY5J8oqlbwBo00wpdVZG8PNUfJ09IDBVA2BeX7Zehq5CTbHUxskVz2Zt86ZJrggmjeWzGJ
TtpiioT72NEQqsMy4SN+HtYl9b6G6YhMyWmmDJMQSnSooaCkoZh0BFjoCJ2PxxcUj+cq0rKKM4pf
lFUo6N5YwjQ901utNSnEai/iBIBNMNaGTFwZJfgRfJsMbmmlMVLEQ702R9BZcdi2LptbvFa56yDf
CdDmtT4w3R9WY1F/gKkCXIP2o6CeFabRODjxszLPEcTRQJZHSFwQ5eMbcu8rwL5WIVS7syzFzGyF
XKunyhyO1tYl2ha/cxqS9XrEJgWn0p2Z4YYq5bGFx2ADrmH/jPmmTLt+MwRy3PlqkYOINMFZvG0y
NFCCIaz1mR7007KC8RIljp9YUozFTemid9UoTDzL8KurvqUDe714LcCKTFZwe+8m7Wk3Rc41z9II
Az260FXqgYBhtzoYY4CVKGoQWFScDUiW76rLOfCFbsnPLjDuEpKr+F538E0kAbrdb1SgSQz335R4
LIFC5XhXO8T9b9KGnTU1pxTNfgw7V6xWdbFajTuGh1SJQ1hFrQM3jCJHwkKXPMef9SsTN8KAv+Rc
HcULcITFsClhuirskRkTVYN12wBFAaA8eJWrRcOFF8Uv/i+uqp5mv/JUAxoTI/0gEMgZxnemO8tp
eCW2Gi54MS7/hGu41ePD5rJRnKZLkNntnXQEGmlatVgtyoXwJjpxqllQ1TBjdZN/9rgLlUz2g8lJ
WCqiTpPVK6Yn21pOsjxxPaawwRDK5T0IQFb5eGHZ8GbvUIIg5qbKzR3HZJ2L5WW9eeB+JUbiVg30
nZWMZ5pl9TfrDulvNcNE7t/Kj5gcw0Hvb2U1QD50cFNlxXp4EIS5hL2Fbp7wfBvStoYacSGmPhyS
5rCV4ifyX84FWgGleNOCn1ypdXBBODaVxN1rq5KzHPvXyoLiFRAF95LllCWRe85TblD1t/DcMQ8y
n/tR+YAvartWiWI9XwOH0UgjoMMmbx8HbYlNUuuXwA11Pl7olZ2jKnLcX28mWWRQJZyeqfTZ2z9i
EeN0x53kEb+pdKT9ZL1ZOIlxSWgQIrRtnIXRolz51sF+BiJwwCVlEn5zedKvM7eo3FqxpRZREWWh
ZaYwhkPuvoA6em9Fms3cwro2/WVWr57HC+4GYwE/7E6GJL/FPztnQgF2qKhEk5rA5WY9320yjfJv
eycCCbjecGfoQSXqJikqeMEVtWTMj2UUvYcJYLwOD9SUP20pE6nLi6va7jbUP3RNeKWxyCAYqGra
OEtrEIaBCs9e6MwQv0EWaTn0L2pIzpRnFOWzew3OJ6U8FoYE9Ps3p1SEThlADkcwx1ChlHl3qqGf
RtmMagVn6dY0m07FTux9hB7NI1U9F6yfTdFvUdqWRuYAfgjXy4SMvEqNhAr3E+1ffTpkzr9otPVb
Mbg4wY6yc+Ax/F4WU+AzCWnWxJZWBPTYoXFRwIdie3tnUzch+5h9LxnJhiSXBeAdXcHuXuvAIonG
pClYlG0CNo/0Ll2Yh8wjWG/lnSVN6dn7T8XlTYXRIXag1Ae7V8wKdE7x4ioE30p1CdGt0rqfe8dF
TlPEIkwc1NZj/F6YmNM18lGAPIxLgyhIMlEx0ilVXSCcX5F0YoiNle8Z9pVsR82TUrPtfR0q1g/m
iMEl84PtOEuEKjn+lp+BluuaCjeFmhIGcbr9FSMMO4guibMR1ER7q2n/keJ1dPFMjzuXOvpe0H3M
O8/UQR5VwPs3UlHIB0DCe+MCAfcgRHp+qJfG5ZrKNZ7PRHNyQiJUqyg0v8tO8OevYT1BsLBsDKfY
mNpne7PDSIx/R69UeaaigZwxRofSriPoT222VDQq9kteSfAds5V4QoyucrHucKGNnozvWTM2KgQo
81Po+5Uft1jxOiGpmf1aTJU7JNP3W7H4WQGWWvbeJCi/jGqWz371iU69l9TSnKfo8d94/F4a3KMv
s87nrObphES87BzYqhGtQu+n1B2HBQ4CuGtFpjUtujtvMZIkGISifJFqHbgmPMXNTRET19RV/yyX
2ZLOYf+P21YE4oif3OnuzmveLxB2CpfE5Idf1rJMnrQDrTMdCn4W4tkhkrhJx/GJoOo4cG8a5f2y
+q643leO9vIo9Yf1fUSKnG8bN0yaSbCPkaQnU0iIlwISSsuHQzFZT3SVsIQLijYrk5TqKnE24v9r
8VyAceAgCKoG7G4acMa6K4wiv7FI65F+DGndkkgsiNqi3dyccwuCkfnkogjr8oc3vNo4wyobt7vO
6wnbs51TTMdLeaDmzKANLZTZveuRlbzwZQIwcWA1CkFS5HuR00Lfu3NyDzlInDHmAMRjhFzbQ1Qo
iw5e9skHwOfPSTUHi9zi7iSit0XA4X3k3e52kYuS/AdZUzpCWq93rMS3YU7DZ4DIwV69sNeAjKBC
Bs7ZhtcZg8YbTcxkuScVmWVBO1qk4WvKjEs1ND9Wc2f+d8emZ7eqBPGHh3iyRdxsBR6oAhTfMWvq
NyCKLZjj5SNtEcH/2NRSZU76bGCikC5urENFJG49RdqQmy0eRrU+rGoioayzPAIRt/aQSaf+Zjgi
r8xgLgbKpwjZ3EdY0/lmWH6zxSqxAtC1BUvkr8hw01xIBnNH6ArjgcLDlnioD5r4c9M/zftZIQVO
CvgwoS4PKnNYdE0aU20F+BvQZ4wftiDKqBejiveYc7Vw+Yx1rb4pCBE0+lhQ+Y6PbB22zEx7Tg/y
4/+gI6MKuMwF5xO22Y2zdhufrmFnSW7VqVxpzJSdCfS/JJleMmVDjhhxq862FEpdgpGnJChi+wWl
RoK8MjvHmFh+pQtnZ1H9+OzzqQE5mHPkGBwYpQe/l70so6SIIkX9ts8Fd1LHa30+HsOFBVzMsCzK
yqI7fD2lHHRqXTB2Frilqph9QlSrxTqX2Yfb8ohGQKF39wG8jyZkIJeRas1dAwbEvI1rUnOmCxH0
BOOZw+EZ0nvhXxIZvxwdvul13Oz2UVpCGZgOvEjUD8rKbHboLYHuUEqkReMjnKEHzyVvziTgAw6p
THInmXFU+wCyvIHCM7MDumcMbYxdt9QA1ZwgLX/L1DFvpz3Un5zM9U+/BmGkNMusA4K99LQpsAuX
r85b8uB3rKLFBOjBlq1dJwTIhl1mV8N7tIakNAvNT8GPlbzfSRwNmYifpFEgBuPZD7DmM20fW9Wr
PScVQBB0AbtBIdwAU3ipZES+fe38nrWYayXF+1JvxxNW1rO3NfU2RkCJMZCXFL1xqAZoyaSyuOBL
QbxN3yoAGxnRMi9rYCx2CbdxQ6/7ubk+XNUIUnNUUzOA/89HdPtT4myjcbhpkIbdWgwatLY0e/4V
A2857Dsx3wsZPd++G+RtVb/f7a+5vLNOF8zQ91S8f46tGglnTFaU2UUv1VYGmoo834hxEtKQJZlJ
7VXla4PdDi+fcwKeSizC3ibKIHfazCa80nv3hroPK7uEmeUePzEk8BZ2G/CL7u48Cti3V7GifiBh
jZ7CbQyoJC0Ck33pnarMFfbzJMqnZ0eYKtu9QsI09UlAarsF9YekgvY=
`pragma protect end_protected
