// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A/49IGuhsm/CLbZPhTQItamdbMqSNLAiVa5k5nuWdbWf3K1GB+zWViAHxc4MPHI3
JIuKbKE3FwokJpkkDMknOTIjsNYcxrFtStJOnfgulnsVOFNGFPa9nR2xql+jrUwf
Y5kAft4G0tdnhsV/MiFpnZI4csVyjQQvtYRF+LZJJwc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13744)
5eLvp1dLQZEH1pbUAzntsJtkl+L/t6zxzxikmRjiuRD0HfNO4Z07D1DbgneWTIfd
hfI5C5InNNV1B9wEs5Lyl1PIcSYlkNpPAKcmo2LTU3BQvZb3f0A+qNpmf57xleSR
B8dbnXqljCjAeHYjnLaegi23SUdAYTNuIzcS4WAmwkCJtT7zfslZBimyAOS2rIFL
1nKkLBi8rEgU6RVCEvvPsp8Zxl+Am41iZ00IMsyyk3LdpFrZAhvBMuKtAQvSKJqu
hvkcZsieLh8RWMI64vsenvLlurIQxmXxZ83P/2QCBa/uzTspt1PXETtv6UD+MvDK
/DfF4rhO4hfSnxt5pbxNrMVPJe6cROInAD7CXzVm45DS2UXp42ds5TG/pI2d4ygy
M5+6ChuwFrfNcgdBBunp22NMDmEKSLlDDSWAbRIIkdX+roQPb29Iz47mc6XrtM2E
V8osPYZjnk5TDBsaLAwyRKWCoh/dCBKbnuv4TKzabReJr1eEbcNHcTWRe47vpC/h
TD4RzowOWbEc/kKtheROvLgxL9NkSO+38Vz2PPHln4q6d/FnwPjC/45OMg4Qbscq
5vSArUuJ9drLGk7emx4UgxJ9ZTTOwjVrWcdRVU/lhVq87seV9ZJ9R3V+Y8l3WLEV
apgXCGwAHTMC2QuZSehf+ETM0WBijkJN9QGjIKOWmkpOL8S50A9oNSaOK4R0p+/a
iFf7TLOlhR/rBPKoUjALV8FA/U90+mGvAYEKL6MJ8C1UlOHCF8zA5jRpZct3Jbcz
fW126ke8tdsUBVMQAHl/4CzvF7UZOyHHrYZHTBuLQPLHeMkjRu3duKiIo1O1jAVo
xwR/k9kpvJELapZZ6YEE3/XH+tVezRYHMNLPFOQIxOs/ALYFCLuTmOkIOSbbCCmV
6gGlitrhSY0QHbzEviJhBfIbdw6kDZUwew/F/BKK04SciHIItK1Q1GzOuICBsAZ2
Kz0NPrzbKZRlGL9fgeKJHHC4C56GtZi4Idqdp+yXKeafNvtqL7Hu3Jf6WjP6WKew
FRDz53IilgbjuS7+ZhaALNw8e3QM7PFBA/dZNdhq5CYjVK7th4UxgHJeew2Cpnc+
sCRgXLkFZB+ZLdB+hxgrMUSjmwa1UbGWARd0lpXGbg8I3Cx1+88XsuMBjvM3Kyoa
iqmxlS+OARs/ixUrp1LiBrQkVJf7J/ttYbxvGF+hjt4AjqzHm37ah0d6yLN9aBN4
O2CPlHJn0hMHN7KcQRcYPmsiNTmNXexaIUFG8mSjKuCC/WE7RpTBTNEc0Lz8pqNJ
+7bPI25071jyTxm6xLOChRWouNeaDDofutpetWnZccU7yKxteUxxSND1X2bUpxVk
zyfFMlLIbS+c6RcXJD1ThlyWqt2Nx75kcRNRlcqWiw9AYTC3ibAaCrmmuSZRnwFn
OwGOONotpXCYO/qDO6jYlxdBDfenYeafQFCGlQJoEwaoXvlgOYIqaKeZZaKh3ROv
oj+Oqif5oHDFqm2ESA8cmFSiaZBPmXdu0xekyCCPgx5c/HiSu0GT0jY5h9GG5q/n
OgYUn61ROu8Vt10rl5oA8Dk9lf4a65yVQBRSaKAaIScVXqW5N+sLIpW26sScmtjp
WfSWhF5o9rklsaqACRGlsnMVrComqQSqn/rUPC9RWKNNB1XjgSwznwCuJvl9OG+K
GMI/4Hpi/RDLi6mAOZrJeQU97CZonNdXEr674hJbD3ROb7MVdW7DaP2ZJdkri/0q
vBKWqKzm7TuzWs1Opnb9ESBz20PGSw6vtcJ9H5qLxTm/Jdgt0pJW7PAnUU7ccw+Y
4V2W2G0hhxI9FpxH84JeQWWPKVhDfiTudTM0qd7cnbPVPIPm3gXJFxi5TO24qF+f
XuEjgXe4qeMjHPPwrwekyKNimr9obrTTbam8f9WA7u24R1QEh2TMk57oaM94h7af
NriVuKVjaE4TwenElA3vu7SNSLwbfnd0eCEEKuwP9eyQlHVekmJVoJYQ2Mw9EVC6
t3IUX9tUNczmJwbhAxTpd5FiIY3IHp1Der5tdb8c7dq2fWe4t4q3T8Y5hjg4vGLH
averU2i5FDXfjGibLLmc2nALiWO7xKlvDesI4rLonH4XMgmUF+3+vU7tDPMdZdaV
a79EuRqiADYgGUP2ikNyU+/QyyI6+3+j8lbHkIjzLiovVQkmyAxDoJ6D1FKHVOfS
BvXUcl0Cpyv/0JGCMquAlapDZEJMCNv1trCcF4pR6i3FIfN3c12zgB9DbsSkzDiN
3VHwQiJ5AuLdDOaixmB21c9Nt0nBsdfxB35h4yfKYOwv2Nl7F/FUFI3I50kG0afL
edf0fnAP5OAwWl0qHSh7TquzSukxm1XXVm0O0C9bPLjOqqM8xw1PL8XRTOBh8rYd
EEBP7m8cDGdrxeX1pePiQa2gd5UAJC0ZXf81NlrP2/MFSYVxy+WfRC5EgMxGx4SP
DEVXnzzYIh8bPe/ZE1tvXYZuRy3f6Fem2G7BYajYQioyQF8+YugfxoABr4tX7tNX
szbMfczZvVXd9+hsjmLla5mxrMCm0J5iu0+l4qQLESq+fy1w0r/DPhaY64gGZeHm
AnAAOOrOoXTfB7fWH/gdEN/2s4I8Ts+ktB852ohijqTkGfJx7fU4XnnNWrIARPD9
7LilcIzTZ8SSRcNPxwv0vhMhsYo69p5RLZzymC2ksYYZJjrCKl3O0Vod8FcmyPLI
B0BL7bjGsjNjyu4O/StOEgIIC4ZnC4Z5IkE49+adh+lIJo77HNZc+f0+JWHmsAX9
uhQsp0iQLAbMyARAfDODeH/eJiqCJkMddnF+mFO2DQqOOqwh6kJ2bI2Czb0uDxC2
+9AYnO7t6cenHn37fUhJsmoJopAZgSTsxXHvZSO2+Ed0CHWEDJBb7XxWrI24TG6O
lW5Le81F2Q7UkRiPMRnzAFYaKik6fWWoMSExY2x1g94i1qNou4fkUJOdFNZUUn03
XDPGYCDFPNx2ie51b91wFqQEDb/T3ULcmrjjSp/croVJI4CEH0TV9D9mJHGG9den
Sx8E+rlJU8b6vh087IQEBoyAQ/5Y7ttxY17FyoBG8bgFgmYpg+eEPqqw2WYmsECw
6dS0UVfDcw6Fc4OoVUO+x5NaCwlqSA5HueediDWkourdPWf0iGVuJN/+PhCmDe68
zTIENbJUHZu3CSqwzcN2aEWqZnRYqQjbUb4dre0fNvpW9yKb0j9bx8ty6qBFZR+j
5M7KR0jP7LGezqThyBIt9wSsdK7+piOsv/3JYb02A2YLD2f4R/rH4t2v83Wr/guh
wNyjt0M33ViKYqKwXvzksaCDyqaExen/7R31+8qYjl0/RZciAAal1+ang1RFpgS0
szUr3dfkh2VpwAGrmMnxbSB14XXqlRJLoRxcnxukikUA+hZSoNeyxjvmXLGD37wO
KjIQlja07DS1GgZnj/dlWIDRuK1a1hXl0A95YAX7ySazO7I8DIrYgJcmYdbgEJu/
/yJ7BbcwZj41qg0Q+CuNUyx7jaEqs7sKHqwkCiGgy5BT5PeO0yt2CIdXND/gLooW
LMUuhIK5IS69Gghza7MTZFFB+uUjWOt7hF6Eogzs3A0fP9oFuYMdTOKCmA/gYUmn
1PDQs4pd7nmpUjOrPkN4HPekKpIsCMstLlbLvqo0KqJ4gmPBAAl3DoMgfnmaSv4w
mkuzpl64b55ucnNakkyePGSa9+xMY3mck1yOgF4E4jLXrSm4ON/8buPo/eo4yFRz
zT9Ou/2+vh3FdFSlpLwmswHVMvB+24MdNUTNJ9LkmAIOkCsusUAyBTXGkTmz3R7c
Kpq2Ey4WmG0LVSgHPifL1OPN9/Szw9pI4PhvPcnKpsfFYH9jhLcy45a+lfFXdwos
waK09K8xACpXITi+aXwJeGeOZjI3PMChrdsU3R8FlWYFzCSHgo7jN1rXlZs8cc/Q
QM9GzPVV76ei4xUnFYy4kiUuaXE3wGb6dxYfpfoSPHFl3rLDVsbyWM9iFY79ppFk
G4tNUOP4Rw8Hka5I2001I8WMpIeeivIwpBr/cecRo3wHuSPErGWTEfVnshZbz8zz
SNjOV+3RbZ3IPcFQ3GhVcvfFFTJR3GVq/fipFHsF/RhtgcJobRdV8AxkhzSSsb9x
MwQsnzebGLWnHvys522/eEkpeqaFXN8b+dIVV2TY5Mks7WQ3WliyRFLe0eEp/1R7
DsDhkR6lIYhgk0TAxyDkZqrBtaMYdUAJxLS9x5AGPRzefDSBR+elP43Pu2mm4JnY
LPy021N2d1eptgwd9ze9K8yYESSi4XtLmhG/D/PD0buTuFPWOuSMC03PLKkP3N4p
wCkVTFhKn6/4ZTMryux+2cCAosw2xDu/22p3hVW7RHr2Qb1J36wqHU24MvtmZO8F
J02jM9Ie9R/cqzbktvluBoF7viHyRQJKYW2Q5UFAE1iOkeGuLtGkL4JZgnYGVw9c
B2fLkm0pOWV63F+azyCfkG3IVMFtzVH5E/V8yp5R29HobcvfRnMuPav/Xta8b5dE
6Ie9XFwzJMA0TEBPjcAj1IV4xyfpYY0oC81Zfd2pnVBakhWwjLhrRAjislaYXHR1
RfH/+WAXkc1mV5fsmmv9sWlzCVQaYYdftbGdHv5ZXfLp2zlYqbsweaaCxall7g55
Kj4EoekiXCVnDuD5Y1uMiMTYoIm+ohWtGN033oPxYXKJE5EbGJ8/on3PZvIm+H9J
4QHmaOhc5UQkU+SPbnIFef9GZn4Q3SJ/C+u/VkOku0kI9Cv5vv+HCnEusZaBNyTP
wK9sT+ZJqiK2lzMnrhcOA92a79JWh5OfopgBOjuh0pDhWcEUH4vvH7Uz/GdVsmHe
4T2XtZQ0XQZEEtZl2II0w3yB8LbrqRmVrebf2iwYsR6bar3Z99mQt0OkX+Kp94U2
XlWaRO0pj1TgEAR9GxLvGp0ZaqJqH8C+xR8O71OX82WwAlGnQJiG1Kt/mVg59n9x
FNIm+Gd4K1Rs1joyh0ZWRGgAdM/WAAi3Rzp9QYMGmAOnJA7dyglf4Ba0jzF/LtjA
yhIpNFfxXmW7OLVcm4CXuBzbUZNSAU3rxlHNujD4LGKViYzhb6Yc4PwqmdYTfoaK
MDrULQm5XFtdntu+GhF9BLpRTWYC52RD/y32MohZB7BrveeMDbBXzaajoslfu9fp
4s4RZvtkhEaeq+7C6JzTSyEH+fJESDcCIrdzP2KRWmNEu2uzTcMWzlYLB+x0edQs
pqrpQTFIxE83gULdIO86vWVs0k2j1PDbYc1fAIvfHl8KRYAkaB1IIydslNbRBO0F
zZXSr+a6OYIxNdTOqJKKtWBzPuC1ceWLqEV36c3pyWDQShZns3knRUkBIIC0HypC
MW+sx8hZoaBc7oFNSZT0GAgg4cjhidUeJrUtuj22nZPu2QGRgeuYx+0hP8FT/blD
7ftPYNu81mFSgpkHCrvrHrH6zGuP+4Qx0trYNPaJo34Fmd5RSeV8CuRu0Hy/jsXh
uySvSnrM4J6JCQnXalkxyc0nDNiwhuCtVFfgQ5Aqy9Xe8N9hImonLWY3MNwsdiOd
4SxDuPZevW+8GCxMRlon0c3Cb31VVvbh8kO7H5jdOMKQDYKGCUelPVgKfuXpA3iM
wn7Lb8xu0bM8LN7pC2/G2+lAPOCyXrNl9A7CB8jS0uuA+D6rEmo1FvfPonUDLXnA
D4ii6MmJum0wI+hsGe4Du1GCFanM4KTnG1e+2A6QQPDJr6hHDKdEIuFtJl5kfKki
SpJSUyBxJ611CQ6rdPlFB1mq+ntC8gnozEo6JuB/R72encOU+QcyZlBGUMe0NWCq
G4RRLGoKSv5BYjA61sNHYbpnaBX9wTOM54ZoS+QJmDbaIyKRZdt5QyPUGuUvQIGK
mhXy6DC0lAV4M3EDr24soHzFaWeA67mcqhOcUVhjI4948rvcdOcIS2yZnHyE9oTX
p7juIMFF82JzI17a72Yi69DRDFr5Fxpe2vyvaEN5CBqquROxNx4SqlmVeZQ+mzb0
gqDdhHEewWeaDDXoKAjLaTW4zz4RKuEIBCqhx0YNC2vhD/XssHUdv7VAClbinLby
PIodN5rSlVJjeFTh8LTLRKwDykYfrFrexHI+//m7BPatyCoT67c0EomI0lcSN/nt
AxQQYsR5ndoybaIawvtInlWQfQjubKrJa+6YxzgM2HPZGpf32kQVgnxnd12lDnUc
QrbcSaMYZXQNZHv8QET77vbCn+aa0uxI4ZOrwPw7vIo0viXPeHFdktCRqCLPOvP5
CriremyV+4XLx1GNUu4D/j8xJv/Cwmg3xiDOAmUSWMTHy00Z4gMpLFHPxUdVZmgY
i63O60GKtuliC3SHC1xA7ObgwYEsjhs73LJFaTVwrpYDB9O9BQCFA107HjD5shvb
ixyCayLEsH96//zHFqI0Cb7kyoSSgvJ0D70p0xdAXcG7r48Evc8Oni0Sz8OikfD2
xZIcYpZAEeLkbj3MgYvxgEtmFpRnEIRJ+GbwgUiFmEsdwB5cQMju0JKsUxP6qN+7
XCw2GymERGODI5u6Bkuz8Rt1yyP5n9ajCxEqiAv/eCHMHssHFtZw+FcOEF4x4K28
iVcA9CtTXNL3a8nZs3exnRrIttRs1YF8iDXaRRceAYfkNszuRq05jSy9/I2e0eiP
+ozuL5mnV4uvTZLXtCmjYGLbzemDZYRqes4XCZCHpiP3bpiSmfrWFK7QHFPcYbpK
vYNqHaStDj4Laym1GjO4YbkQDiayNgVA4eSEpuPRIrqM2ZheCsDeZQNFv/9R+m0Q
2vLedPE9x3lRStwhJM7tf/8YNpbrUEBwSUaw+3+kptHYS8UQ844nPyfCyiRAiI89
9gjvz0raQFKwQ6yQvuVQXL8/kOPqhEYn/hsXjDyKWKAd3Yt4FNfeWALkwA6C/pWG
hRFXHgHK43WdBd6n46YfdMir2pfY8pOoZ2P69OkK9b+xl7c+SaHAuRT++52n+mZc
g1LLhLQKJDZUlcZ44pYU3E1VoOFVQTyxyLw8WSgDxvQIBSHSyDlFQ4ulKMP8LfHP
KqZpx36Gv/HKXnxS+cuL1xzFND/R8l/j4EfYX9ptk7SkS0qfoYbjrqOK8DGFwD/r
Ld4ma3IEJfrcW3mQcjKUyUXy1f9XcPALimLnZiUSiAcJIyEATFyas76bVlYzNQHr
HV6S6ujwhNI/+kQ6WMGAShwtiPTCleJVgG0lTaJqp2ss6qkWltU8FTU+IDHEWqnX
CSrebUblGYLYPkP509EIR9R0ars3AVPuOJmwI/2pQq+n2f2kVfmTYyG7khIH+CQo
OOha7cEU4x8PGRpuiw13x5yEsRUjBZPC12jDsrhXzDp/NLRyzWVmW3k2diOshiTP
ZOkV1SR7v32293LuxDPIk4ISv4kpGdATzHiXhBGo4Rsb6jqDFU+vd2LqJWTOP/ss
FWTgorwKE3ZJhA6B0AjGNF0Ve3nI/hsFinly4/fULplZj/LQNTUi21Jp/4Naj+n+
NIgs5ql84TJqf7LnNiMe3gfoxa+Xaz0JXiG/IXh45dFOWEXrtX54vAopFtXYJs6/
pLtqc1I2ztomrUj7GBF18kNKgeNqE6TmoZD0zP8a1DEZN2Tx6FotibXDknxjU2OI
RwUSaVa6KZK3BrbYjJRb8SpzJLX25QNZ+4OauRT7nZK3oSJJIeW+vTc/EJ/HilQb
egrA2bpQUs2jJhXINKVi3ceVeAk/TWH2hbyqezH+w4ZHtEWmouKNg+uLlV20K8s8
aO8YQmCSnwSjljS/uk/PQz9AnSoapi1Pa67S4SQklxfkJU08NUBjTinNBLIUex4Y
BpKMdMjHXlbaCCR67MF8IJZ2FKR/wINPXBSZaD0jQUpBZDMoRZGATUsNCNDtdRIx
/QEl6FaVQ7+xVo44jyK5B79GioGxw+pdhbpxOcWFancAtrmqAExz0Lv9PNuZcb5k
59xrqVmvrDdsLaXRxRrmf2/uYYwfb/E4WOeaWIOccynRhFQG6bFrkwRTGuf9punp
9tl9KNyQGZTfCb6te86NYII91cvQdDKLqYAxloJH8gYIutPgdZLRBG87xmeJ+qss
tvBwmu1Oldu9YjtAINajksIIwF8PZKSp7YgPi5eBP/SIzYWoLm6IzElpmVuP+izI
Ph276MEFeCaTZ4+uLvs0FMuU/43BDaxWxM0V2pbKlE88j9IMY0Ku8Swy9aPDagjn
JepwsQiTitOKka1Ylike9+IvVg8vGhSGh6E/0XMovLhsWj/VrYi0p/cxXVTKMc6U
v7d04zsX6FlWMzTidHxs9m7/hN5XwOxJSKZ3DIVxLtKQIgu6Zg6ghROBoUEhSz5v
nUs+AXCNFhCnaRWRTaEmMSvtny7M0t+Ht1Ts5zealI+RUaGwU8QOQcOmuVYYHWQ0
ti3/qyN8GiEAhu58Va7y0/Z6L44xEvnww9T8wsKYpnv9nQ4V4TtioPsnP+lSO231
Gkwp7PqyvxkOnWLg8jhgXPr+96rtZdBG+Hqaei/9LFgO1OJdvSuoWHxRBOg3QNZt
J7h9k81KuZEuGjs7DTBwOTtFwWMdt4EaS3NcDOeCHvT6Sy8JuWUGKOGG68Rff3DV
h1nVIMF6LzCpZc1CTTumwa4HF+r8BOPqFnmZRgqH9sgNNxouwaYCuxIhX5H1FCc2
nQuo+3iP/zpE7nkRaKauJXTPoxr3vdyHlV9rFWnbeVaqI3tw45dH1GhnfhAFXneL
EWvNHWEcRJ/fzMniNkBmDtVcVPOTBYh5AxmFqPz9oJ849Ofywy1pvaIkaHrthJze
njijXLf0Q79bWR0pnJfDaYpjuQyWM385fkTjmvIQMNdst9M9QDLuCOdRWJnU3rvO
l1ERQE5PIlFFbCwOpMTUdKzDUvEvEKZQPGDW1pEt8GLrF5sfjIZO2j+z0J/br5p7
LY4/jFH6HFZBIb3V0UhHaAVL31DY43hVg7L80HrSOFcmAfpgykf/DG1CUGWOZY7T
13ygXuT0s2paDJCNao5DdogKaovQUisdALW3hQyY5akoSObaKVbFm5p/idJsL5qf
mQGkw+5sHE1uQhDx8VXzFlA5IJaqGcwenZhhvwUm/FcOe0zAz4ZQftjXXYxA+fFp
qUj6gnor0RQ0b0aUCUvYBFTmbtTSmhtIyvXfvNCyR2oIfv9Xk2hh7dgZuFmjcqO2
yvNM5UchuhNABbc4NEHupNje5y1+7I7aTycFWdSnA4ntHemRgWkXa2Xww4NI3DLZ
KVqlf65Qxf7o2uvM7+6vuEMkw5JSFpehJXFQSTsYx/Xk/bx+piM6DCtaQemDG6lv
dGmh4QoszBXxZgMIxk2lyGzf+fGcVsWLNiNPq1r2Cqxxu5YvuA+hhITF1tzddFEn
nwQC73pHSsw76brZ6NdfJbcaXg5aHzJpQWmVl35TJlmzPFd1h6JTOlkMjHjME4JJ
qECgi2JGmfvgi64wKInjQZz8yEwfnFTJHMDzdR+znpY9eqiux9j023i3ZUQGjF++
5XaBj4fGTzxDNrMlysfbbfPNENiTQDlBE9kvUZNAyp4pf99l9bDWJz9PRgkI4vE5
kaHeG0jN9ofxPrKJu8XifeHRCJ2ZXYX+FjN/08P3nEd/wWMIHF1gP+5TWtCmdOBr
P7Hp+svpCxlxcVi3d+Bk24iSFPJuhYGlSXl2qc+yJaGGTZhzWnMRrH9gHEKTycs1
6ZFPj5lhB3hlF+ZeYa9bhzcTD27SQ4bDMEAZgFWl78lpe4+Tc48q/Q8HtPPgOnvh
bwG2aMxFMmuBaVjAvU8Eb6oXId4YLtBRUui586hr7OsXK/0nruGCnkya+jT5rW2i
oyuVcmENiWMxQdzVSVOPsCaqgdLZk3BionAN7xcuzLIj81LPi95o1R+/CrlUXDEH
j2CGKaJ78WAeketxHKmDzy1zVY0Y7VE+h1J1t2UJHJpZBID6F74BQtMqUbvfwQBl
YNdOssYD0y/0hs5vSZd5JSuEa33sCsWM1p+PNGIpVKowXctERAXbNSYkg0wZzSHi
CB5qAL0Emp3eDAs7VCAtjReQxkD/zvFGk9XSIMmtYAAfL6yn08WwAqh54E+bUblk
x5WXiIDy1mHtap42Rh0d8xRa+u6oTjcGkd9c4LAAfnjnWQB0ngmIvGWF1o+N2+54
o3JI3UhtAOdK+f0ueREOXE9KTiVfgM0Oi1AtfpMInNX7a+5WFEpTRR69ARu32BtU
fVOphwcyeK9c4V5KuFPEk2UEcYhbnebpRrNkQmvUiucsTR+BTjxLrwlgQGz0b8SB
wKp/7vYWL1aOUuhWcqF3fNt80c5IXe7cFDNcUvEkzk3brENtZKUK9Q8Bt4OOIf2I
VJUbXnT4jvRpOTawJsUwKJFpvEAKrvEymEB8i34D7Wl3an4870htZNUWU9ScGGy0
w0hiHrMlcNAKrMWW0lEEJx3jcdwn8PjObyB+vBvF0gSx1CARW6DDV+FDsi43QlPT
ms0chWEMbNwEYFU9FbZ4Wt8ioIR3N3/Vatv6/06U3TmnUCpnjcTJZUGeZz7S36Dj
Z3RmIDkG/Jp8K4IE2A+57zisCz7X7q+c4RMmQT2ojsSTMcsfK80We2LJsNCmDEO0
sjpfZ/T+zYYf5u84Qwb8CuqYYR1uLy7/jP09APjKTMxJT2s0ACm2UWWpqXfqChin
i7BFk3LDy1E2q0DUGpMarcoe1ZxadMgi+Sr0KtFud71Of0Rni3Ab9hFKUqGgez8p
th9YmTidDfqrap+nUPc6UchgS2uFmVx3A62r65+pcfxnbMhPb3KDjXrhchgfSpLn
kjPCx8t/t7WjX1yajdAk+wjSf+vxxUFECnRnMOKodw7hW4A9VsLHWWWtr4LpO9aK
M3zU5yym2NE7Ia+wArMdOuqcsRheV93ZZJXXx9t2rxb084hHK/lj57r9Aeq23fRn
JNh4PyAN/j+oM7hEY01YU8v92hBWX4fbKSHf2EnmyfA/abmomjVd5r1/lQAWDa4i
kS9icRtLvnnfwqxXG9X5GiPZO3OEe6Tg/dJbkalxrftbUHTMkkGq2B/H4TsoxSMV
AHUq/j2KViid0kTxO+hlvPxj8soXCmPdqkh+c0fQHxiWU7Nh/YInNAN2yrPsoQHD
yKJn4b4T5firC6IkoUQywgCPGCOEFC9Np1JxbHzS87c0mDA0hWrx/4vdOucEqh+R
SFSWUOnd2I9i7SWDCkmYQUlWXGIU6rLVkNXtqEcvzsDrantjwbmTgn7exlyk0sQM
4X5VQpqceJEdHTYFPjvtnfifSifKtd0fm2nuInOYnKt/lQtnB/CXSejJCh0wdB2x
pgr/O+Nx9+Ye56Xtfr863MIB7hKmeGSB3k7Lw3IdWLeyNdQiu6UGfMkVNR/Pbhh5
QS05veybozzqaf4OrGyPnV2LIq1DsVSMOIVg9SOIROufZmgwlnz4HzYKWuxJv7mz
6bOp7Cl6cepKkFug42sK/uIi0X4+/nZeaK64ShW7iMcwLALLOi36zlEDoV/YH6ow
becoYC/ekL3I1AAY4h5LX/o+2V9SP/qlYJsRRrULkL5gmoVjoQdxidp5xCfVqsRU
ZUbwZUaKdl9TB6h0uYg6iwONi0qKnA57WMTJJAqMCxwQWK4EfirRhn005NWtDeDb
KVzhXy4pT9ERyBigCpbHBHAaWZX5EUVjiOAdbltGcalISoDWUXznOX8TVGwZigSy
m5YoQpkP0UulnkB1/IMgfoWLEVJk2KOpfQXjqIbZw+KQooIjoLubwVOrq4sBt5Rp
NzW/Nq/OkKzpEMtxarRMtUjnIbijJrmEVbbdJlkBN0y2zTYeCrZlU4b5OIvRtejk
uqrPGOxbRPLWUSj78c7mHrYmALGk/A7YVdUA0oc9mac/gZn6ZHC9EFulNQYPdqUb
JdfKk7LLVtBzzCbCUSU3s6V/luFonD7YSVTYbVJGJccCgKrrtbAXulrAL5aeQAN5
+hd9pLCj0nhCZPNfQI2Ljyerp9Xpuz9mE3vpgDSZMlL+LqMXugn44xyA9nlcEiF6
pZ0ScGhz3CVQtz8FuBpudA5qHyCF4C/7+bstthtubaRmXknu1JhOPu78Q7B0kukE
lHS0rIu0Zi9hHwpEaNl28VjcoTyK/PV07xFKGyvczRiCuRByHEKAEMlj3T/M4d1N
sxLUY5bEXcR+9GcIhKCoyTHo4+kiS7ZOLpvpWs8slITkZnscmO7WQ1BygDL4gB18
NDmz/0rrB595yi+dMXkvlP36XwxhTetjsDTvTQAOAlVNz7BkHInaIhBWYLQtHRJI
PwrJswRHcf9T4gRQlNqTY9U1yL9zNNhJOfTtDjlJO//tqm2zUxAhKUGZS9TFHaFd
MMR0Homfhic4heoRcgKaoO0XbzdCIpazhj9SYZ/izj1gCMo6LOPgQm4bdmGM+z1F
zAix6xjfqKKAzkUaQld5W4DrbgKLBKtmYGGwWpSDbhTcvoesx9LW6tjew3t4cqTT
F3jAxr9iVmnLTLQPyGH2RT3/QxxHk7SiWtir53dC712ZO7YScNrZr5Q8l4yLZpAJ
O9AtiIGD0PCZoTL/3RT8N1V7qwDaoaHA7SUp8b6eDqjfNQrMIwXWbYo0pxkyyAze
52ATVby16GJBk/LdTUSdVyWqeLt9pP8BELmEvkklgIw8dkQZp4+cffvcKA9GzmcQ
yeQzW5Y786FgL99uyT0MH+caiz8I92OduWbCeLj5RJUaJPKCDso7bCYHjK+8Ict0
A8vVmWNlPh0rn7sNeKUpX09DhinGUst2XEOaoXVmcz3yHB/jKzHqrb1BDcPsAY7a
vGowCZtzK0UGKZ+WBDM+lUT61dGaXuKBP4gTkslqt4Nw8pGNidOdfOZW6F6V1nKa
a8Fy6ih74/Gsh7vX9NOzjDi7Vs0m++ZSxxdHSKQCW4i3Ph44KccUVgBStcR5WYzG
j1dADCEGn+NonHG+T79aw1LhJb6ENc4qEZ8q0hg1ob7FhpKHilydB5ldptuu7Pmm
9NBRnzOy/s4G6tRgNxFf+WVvEYV/b4QWenoLsMEmsyNH2SvcoQxOFvYjkSioMWtI
cDqscsPJ9OqYKgnby0+GqC8HmkxtfxYW/5sEOOR9sItKy6IXuXIXIe0j8nrVAydZ
UDZhmRG3C7JGuCcQPs6z57umxgniV/3Xjyye9y3qEJEn+g3R1tUKbWGlQ/ktCnrF
sMdPL2ZLkwePGDXUpjYUOqoHflhj7jTScCRPOdA1Ft1SK7iiLkBRFCCPpNbr/Ffa
iLJB9JF2kmhGypEUdqYmfq5W3GNGCY2iMiHgVlTJMaiaIFwJjMbpiDR3hpmsUQWM
bxL8dtWe/SxZjK5MdR52uCCsaTT+SWnIthwFHVtdLkS2AuiyGd9Kwwld9TG5z0mO
DOEq7OptRFrCFwW5sFcSg+pufk7jF62fRdPFmfDqAhISPU164RvzaxxYSL3GAS6V
K0qcaPYJ8J+ydMknD2t3AGSIrcAIymS9Bz5zcwQ1meY73+IzQIh7zzo2N+G7zsog
0Sd9WZFax5KYQb4GdUeCoMz3F9WecoMmGfCJ0SIvSx9UexfumgmC2+OJ5HX0eudD
Fza1m8jCBG016iyLP1mjbpuR3wLtCCM5yZsYFseGKwzInWzQC4gb3zzjgp+ZljIw
zen7+ZG+tx26EDcYIklK1I8eiTrKeU6SufsIBh6wcYQKsrF8n9i/efLYhUh7Oo3K
lyIUJ90jIBERvJNeUKgqp/DGJ+v3QKe+aM4G3u6O/PE1jqIKClGO7bpB1gqjt2Vm
p08na4nKnqAhYWuPQeiSNDDPG14rj6cQHN3+0Gep+PHtQBU/BGUz0/PHLhTixfND
fq4OM1JFMcti79rxReXDvE0CtLk9YH8+2uPmJ0f6DyoAQv67NCxz6aTdKruRBnJg
udlX1MxCzRWEvFbtCKSjZNUIh81sH9ycw4RZeYq1eCx+huYa2/bkikgWhTor9f3D
Ejz1Pf8agzqCOEX3JrtqMd9NKdxQQEITSfhJekaQ8kZEvAE6VFOhamsS9NGlXhmB
Y04YHQCaxCBzrpGyRA9D6erweDEwUa2RYnxCpzNVB6f1Q1hlLP9qZz8sujheHVZ7
RoLcVsbCWR4oF7Mcl8MqbNAy/AMLqiuHr8xsJd9nNZvY4IISyGa08Oo3poQIZuKy
8RxPywNc2z4jqDEb9+LCmk9ZTUyDkaTiLlGfANbY8h59HVUPytNj4PMoFLrd/KRb
vssUSO5mcLc6QVK6ArV/FOWVjf/P8ZjYhgOxPvdyMo01hBcNWouoh/av6AJ0BP60
uNkEoKtsjqQsWt/hPcJDlZX8uzmhb2aXjLelNcs8dUYMXjYTeHhqwf1+G4HRn3ne
NW4s6o/4AVnKXpMv884hjcWSqRf2M993UZ+82PXfdd9Gqf8FgnlUUtc2QLYLs7f1
xHPBxImdkq1AN74BYZFcLtJ6BTgWr/fAYXPkTsSPrpsc7MbYBexZXG7sjulis/tV
faHUgcukGMz9aBA5U1YavqoXm4PHm7qI485HaKQlhsk8sHYKeOHgjAStFV+8Udtq
1E0UJTpTsO/IArZm5f/lcNp4hIMJwnTVW+s3VUwgrkta/cSQYJSFmDNydQqylI/+
x07JcK1uOUm9MfXvTZKHHYUHl9g2JScsIUh68JvALAmCgylu00l+JmtdWD/FV1DP
dSdkandE4a8FdwTDRRhfpeWz/qBxxFK12YtBJgo1PiG+n+4IfMTyFr334+Y9kSzS
jVrI+Fw2s3mIXp72+reaKWmKTdsNnU2DYWqVZQ8wjNLNQuvg09RwfN9wzYfqHcoo
DqNqofOie5HvBj9rGAnedmTqWWlH1DoEdqaMmkK08JSsIGOyvzqt7CXYctiY5xaJ
Fop6hWA+B7AphZdbeoAHbghDcowfOVCI3jQIRQZTa4ZprVdehY1oCawHfJSRPRMW
970W43MuTLsto0eKKtctmuXFQLltMAICd8Pd14iCb/Tb7tx7qj65s9zSEMo6gkY2
u5raMengjMkrcR/BFMUt5t8QAXjr3K+1+a0WkL7xwLCxfIRwaLpvGO9uQe06Idxx
kjcBIbO/ySzATnVwtmJ2+ebJLZn0+seVkqHeHmdOlmLu9M5EpCNh8HhJZ+0Ul/5d
RMZWNjxF/Rr3aahtsm/EPB/2kDzU97OBOoJnR/k+oHn/MWbhroUzfXU2+20K/rJ0
dlprH+ya7fXD9PT8JzlEzJ1uOpmCqkS2dROtYsFIwe3Tg1l9iP4BWxhAiq00dHQE
OEv3AB6LgkPnvsdYAq+p94ZU5NVYFRkenaBSguYuRNc4fYAqDmo3Ljpmm+Ff7HQY
k68elon/gD+o0L75UW8cKUYcffwROaT/tt5vd0shF93HKwOoQsRiQ16OHh6ijgoK
Txxg1+96zZAEgRlp5ZLKWVnt3K+S+po0B6uC8zhBqeF+SYskM+iZhv54b3/7GopA
OC7IX3vEzdmaFwqTZjqvD6tUD5hZbfbYY/pAn5cEuBY+8uQT1oCzSCK+8HejuVwl
12Z6hrOYtlIWXKBZvvVs/bzYV12wEuemAr0UgvQOVpvlnbS+3OTDCiVhwG4N75cC
3+JbWIXgQx0SraxVe2OqUSQILuMM5I+tpQ6iqRt1eFnxkZCvI7M4EsKPq4uTWGHz
wKIGyajUL+8aqGIJSCocHw8lxogx7qMuYVnN66HY1Nj4wzxikmhwEeyLfUsz7JkU
6IAA3wD5ry9op4np7Hkvhq0FcVP20DbvjZ9SFXj5aORqaoc8H5TC5Z3VCHKoYCCP
gbCyiQ2/gKu4Ozto7zcoHvmRlI6p0SsaLlIKqg3ihbEyZ4KgkhLsElciKEz1JBLO
pNy3bltK+KVbfa6aOFzGJAtCRvlElLBlZHEsiS8r7+VHbAFFgm1sQW4lBbtLKgKy
o6vcxhpzH5GmJHDvTuQyGCVwxFEpZplHIeJu3i8KgjjTbMTIz47BPk+t1jhCugLW
kPAsDWaE/FbaAUnwDYO4XRhjsSBIIWuB7v+9LZ+MFZb4zzNaQbLLUqohh6GM4GZz
20UKSlTgufs7om8Zj2HkHYkUe2J1U5usIJvpw05ZY+s4jet+KFZiWOdRTA9fTEGN
lEWw+FcLTrq8Wc6IYzeAFVAN3zqrEi/mGxcbRdNjreRRZr6iDtvloMQlk1s6Ffn9
7RXwugtwUay9WWTvjGLxKmC3+4/RbL8n9EL4kkPYxxRAARSmY1vdIMqJTfiS3YUL
hzs02F/nI/M3bqFuC4GkKRF0rigOTSX9PqWwobJgxJH1rDIvL3yuISL7biaASTLl
1y9OZmAkfAZScCpg18wgWQQh3XmqeSqwkwFr443t8fVCSxJlBoXlPDu3EHPg/M50
vseaCAhKeVm37I4rBmAtUU5TkEtIVDYpJ99YcxO6NUITjZIm1Nwr7AEiQjE0zxVa
jWsPds0Ws57EeioxplXSDQ3VOP3XWrH8atxrBTvNN4UmAG956nzFNf7m2ogQvfDt
XOm0aGe33Ijsvk5FBLEiTyQYfRt6G9n7euo/nOxlNkqqxAJkeoMuAi2mMnVVRUNn
OqjW9bL25klTvYg9b+dsojF21JYpX6iXEzXs5ljhFCTYbzWuEXfeqpeoXBbVkH3T
M8wfXKf7I9Vxe97xGLsqOZ3wvRNvFLHd06NT6+SMoSRmUsGCFJbsc261hIMDSAcu
MkoxjOe5jO+usBoyk1lcQIM4pEDsUkcucOWsxMeRomVi3BNzpgUbuXCHeAE62vQL
VFqlP3Xdahb/6SFGHg3e6bkF3EmqMmRlc84YnecKF+QpwZDt2FP/XUbCwM1h3Q2N
SFW6mcvrv/RQi2gvYsxqEfPZA4tvMq2O3ugPxOHMGjhtf1zQ31c5Vt4NpFzjQr43
NMr9LwLUDv+/vI+oqg2UoWRJjLfw0OJSCNUqWHQQSnsFGr19mN8uFZGFt3xrp+hq
zfY/shURylUM9tZQjeKHN81SSfYrNvCnHE7MlDlfdod6zz2TrGuOH54qcbpSuOkN
VnAZ7O8FJLtRb8Hgoim0iEFSD93mgC1fbgvFYFzZl4rhYDOx/WOtXmE+hlnHzaY3
HYek5WijSTBAwQOvv7ydwzyDzBrFH50rhilBTAmgE8moyKUdwgRYgQEbYIMu5s8Q
72/l8F+H60XEyOi2I/6mV5TNjc/RH06axM3AatI/nA51LrPDmGuBUxVSnbbuAbzN
uImAXuO90VV/G9S8KMzqU3kxIaghYr87hmpNZKfb4r8wktX8s76mB81E4xaBGdXO
XCM1pjiS2LaZF6n1+C8Lzhw3xtR0VxRfl0D3WmHYq1szMSEt2iif5Mw1MkM4xCE4
fWAQ9/40E7mgvCCNBEd+gM7WPB2Jiwv/JMLimoZ4AkNgbVGX6iTCOfwH5RqgbZyk
QGq7TnGCN2U319BxKcX97mEbQ+6HbuxK+PnEUb3U1LHLkXzu9BhTIh8yhuwombEV
nOYk8uTBm+COB5YpGc/1geAo64WiIwEFd7679hhnkaXFW1przj/4rCjiZbq00OMd
JXgpvwW/20xie8+pHmOvbBpqaYT7YeKBtvECRwg6dodJ6abHoLFZoflSy3k2IShb
qa1U1rzfF1/plwgJpfgZkvQj+Tx0gadhnPbLenU0BfB88vmo7DIERbMLIGRFWyyt
cgG/GwPbYczydPztqnaBg5zWUqqlk3YOZ0u3445ex1ATxusLMp4pwv2/x12Atg/u
XV+dcBGDCvykIg+lPUYvNRXVsPE3Fi/4WcrmxVbf1m1KIL7pm30rgAqpzzFAnnnL
fMUjHeuiEsQVapihQ9M5ILfL/bJBlYqo7V/URmdia4B2THzLIRh/xxh0tRBjnpWO
EaQJ528tob7VfY6G8SJnTCXLw6rBqZocK5PuNC3cSR+oqDuWeJ+LQB2f7sIFfOUF
VQ/skwLNUgIROu74d5ZI0KBhhW5nbflV+rC0IXTfZw5/aDot1aGcUuDszsgzbPTt
8EzBT9WGUf1Att5vLfrB8UexyDPTfKWLP8XsZBWPOHAWkQOjiryVkog2E5tdkPVk
27Ljm/Vom3LsJHkIPKEddmUJ+uKWWKlQ1vTIrK7BMDQ2D8z3hlbZ8EF9nb5dFaOP
/2ylxSndm9L3y0WJUf2YUR3wIMLx5yjkwEIvwc+XhyuJ2+xzCJnHBGP9p7BLoVp2
TWRE9jKCXx9TPhBiuOnSG6qplKljMKNeMsKNK7K0L1njV+pOHB/ZyiDFdXcUSRyv
nqyywglyjXr7xsowYM1oOfQzm4ZmdVY2ZWm22jNXUhnwE1+cCT9ltal4tBd52D3Y
WhchFsD8n0T0T5/dqm0GUhyOkHyjGjKaoe4dFx5vzwazI+ow8nhGM2/Wx72LVQ67
ugbbtUaDboxw2fN7rA9EgZA/jndc+3Kw7KYBPfytZ7ynyQT0rzxFdVw6hn1NDdNt
c+EllEjtfiupJSWFDajwgt7NZq5gU49ClO57NEZPr6AEhWg2ZXE6zdff5N9xjhMP
OCHMNftXhpoM9B539Ph6vg==
`pragma protect end_protected
