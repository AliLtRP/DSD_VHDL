// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gvF3npcYUFKV5DxevRB3kukXAFgM7bcNEYYoqNK+/BTeoiqiz5XqJq0mTxC1q/v9
RErgasZt4pdq7q/1jvDyjpJhY3uJEgfIjPIDSPSjzo2/SllLPcVKIN8ayrplRiJG
snv6Oh80zYZwoVxrFBLCWM79psuHV4XAA5yiQz0AeTg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19264)
f74tlTGBtXwF6xmVSIHErjh4eJgWQpfJlRkEmTh1Xf0f20N5Zf1EuicY5gFoHW2L
4D1SWVUqICLlkSzkN+X5o1snqrSSiFXBVsgD2mwzzi7m9Xi2S7LEDLOVTSAa6wUR
d0+JMONofE2yHsLaPFMZitsPrCeGDXq3hx3am0dwdBzTPIA5zPU6QhjrkIu2UHGB
Uj/9fc2+cK5eaFXpjk7H7M+a0vNRkoE++F9U5Dr3BQqvH1uEdJgiRnUfdHlM0gk3
CL7zl+1ILtG0L/Ndp+jnDoO7RrZueBmky60lRzSFhSMn/eUQ7Bib1OLhSJ2PeG9f
pBsPolhAgWDI1rB6EXaSymlz9lQ9EuqroQSld8pLAX1z9N4LO//uHjDV/1flk+s1
VzVoDhEjvnbICpdmKiMo1OGX6zcvfenVLILdReNUmwuZ/ZG3LwEgCsbuCrPl4d6m
HYhRQBW8UQJ2DJm4YOVD8KSMrI4YXyUy8Xl6L99+aLRb3L2ktIy1qJffdUdCbdYs
l9DlXD0heayFE807LR8DEIZydzmHU3b7glGXTcrUXzGGdPxQzr0rKxM73QYoC5v3
1q4RySJF1Jcsc8Lhi3X1xyAekh94AdAztayoUPaW7p+zT2uL5K8U/8dHdfo0RFl0
r7aRBI43bTnVezZSNAIQDGvv6IDjCGMq2UC4qO5xixzK4f+IE9cGOUeYn4tCjA6i
/BSYwfh70enT3xqJtxPsuMgTUf90ZVlRIsxbwPU1nmNo7+kr4XH/OfdhRrGZuPYG
qKTwPIK7+2g5RUo7RR4WeXNjDgPqwwYHKdANKr+PkITFc0uCJ54w5XIdBUUFxowS
MsjW5LUEACfpJPeA3VNOeEmdk+zDeOnaIgL2OKJyyG8ZcBoEGaFoZ8Ff2jUpqcm/
+yVs5S8eWzQyO2GE42A3j4t+FmlsW83+rGSP7H20BPBP7lqctmFsaZIA76zkv7iZ
a2WVsF4RETmADogYg8L982lv3Z91xTQy+K2FSw3edADn/mxAKmQS8RcXe/T4gCQb
cJvxifMMF1F/Nz2O21c14nHPdeK/TGljIEhiSv4RzeUeuXOX1h3Hu3xI85n9TRVS
E+oWpOlbFHpfA4VdvmXas38FSeb3nF/FBG7yyiz3/n3hHQIh/+Xiqx3YDLqN/Fc7
cOyueaOtTUQtQPA4MkXoLQwfn2R7QODdTuONSO7O6tHrrEhMMoQDm0DLn2pYLeZT
jla6h4FcjSulOLc8hRt8cTJ0u8gEaMvXHeHsf70VltyptXIZw4m4gQxhpyZAqmRa
lhpDU97YHHa+hLahc/9vp/KYMloZhKP4V9N9nanOV12/14K/xi+HAkTGabggmvNH
h6kHIy1wHaGlUCH96z92Sg5cDasXqOgmHgp6mWDENMYEV1gG3MLxErHmz3C/XMBc
bYxUp/sTmp0xj9rLNKnrvsQYVwMKxjVg3vTWgZJH71GM+9R2KoQYQwhvegzcydpe
uJlZsuQjSKU8N3BIEtHm5LZWm263yBobr5V1YrCFjGEqkKA1o+H6ew6GGFOhqsV+
p58Z34rlpMHfh+mFfKyF+Gdq3EYZXKq4gpb4tUcrLGvU/fbEvvhwpbC7q5F9c1Yy
RqoGmGjJ7AHLXNUpEjIueeQr2oaEiYR+K5QfedkQz+vW4umqU/TkeEeqWccVID9l
kUsVg3ZEMd2RLnHo2QeXk9gtMQJs5s66pW4NTGcOcO3WT0ClCXizpq3GCsoR1Sl7
m6D3yzumwHhvi39CMzMDAkdvLy1MpS/mPC5UyRaVtBmG88RcKtFnVfItlXlGTgRA
gpHTeNDPYuekmgdTlwC25/5rVHYmMIY4ks6xKDBSjeVJNL5Pmbub+z1xmMYkI5oS
yiEFDDLHchA7hdC+yoy8KAWyegHW9QF1rBbRFuRsECEclfU/8UdZ65xXUEUZ50aF
16bqeBooSaRdBAqh1l1nnlRRiSTu/T8Lq9tivZmqNxht5PKuEBSoGz6LPBResUjd
Djroa75NYEuNcfX+/Uf/dRfxLSH8VlNvvtVGOyl08wuU35gpjIxFKFocC92pI4oC
wilskmk8eRoyGz44fq0+L7rVma2h7f+jJvN0ZqHqAaK1tTSOJaMxtAsvBPimGttn
jrBFSUOOXymexu0XXGks/VZrgVIzUZvWxCBZoO2y980FkriaiOMA4s3g68QN/CGe
kTHpBZ/uANiun569MxKzfzfk7gSIWB3ytWuFkSh1cvOI6pMfLGW0XMujx+gfI9Ac
Uts+7CgII8DjBZFxEeGVqek45h448Jvi/e1wzDM5yM0Ja5GxGHECWcXQHFb4UlEg
I4yggE6QORxjuZoEBNuWEeq/0OuHCSwXFM6ATIMfbqc3rKbxvH7oJU/0CpjlZfTE
DM5EHCvaWV0i+8WfpiRylZY9oGPWK4x4gLoSNQzwEo3usjrcfOdaFwGCS/vNi0Th
MFGkIRHxGpUuAtfOKr0sQRywoJffE0abueiggY+iYpc2VUuJ6HX1qyx+WICx+2G8
BjPhS7F9SudHK/edGQmWRbtK/voOD8/ltijOIWERLE4kvQbHY6JdHWrgRzr6PFjd
ysAqPlP61JNQ+rKhCFL5RWUdoxn+AEd+zrJ7gN+hVauEuR9Z44A1er+naeiR2WNO
ikJjYBX6PjbE+uzr9gqxxh4M6O9MKfH26yPavR6pNf3d0vcxtjj4Dm80vy+mBrMR
CMZjjKFcosZT20ihHOV7621EfFiJ1KmGWzHoVca/Aop8TiAY/AS/oQ/XmgMG/bdG
Y8vRtctLLcKo21eOWcApVu8VVvF/JbwpvkY5Shwt2FwrJ7NOzA2D9lyzTn3GGeLh
QL0tWh/v/nzJ9obSHROvxwk2wuQeVweU8ja6bmvPL/NgylkoH/BU1dEPxlRs7GPY
w6WkspArUJs6zv6aDwkUsEOpN3yEVJDlEgaSDrx1bFdtBxyXleYkrzOLSgoWiA4D
Eu/0vk/UCs1ec00WbnS4DhMy8agVhqe4dtuc23IMhFo0zYaaLqz1O4xdN/JMfJvb
Y56+6iLd6gIC7fEEfk0aL+bPYOAhE1op2BU0Ydcewxg7kvCuK4zCS+Du8hPtjXs2
+rFd5vCItecW3409U2bIbVYIv1xRE3JClEtxfvkxjbzVyQKxmDnaFs/cTtXWwcWe
+ZYMe0hx/PxSNHauio8pV8O5T/kqoegqJVFrDtWB4ReMtZsLUmzRPyq/m4q5tU7Y
g1rCnbYMFlx8XTsPqTZWZyCMWTr0VN1weAw5eIKhAZZ3ZaaVid196ry19pt6G3s2
h8cq30D86x8OHLCCn0yzxQTQT2UvHuVmu4T3FIUdB+AWgUEDAcD2c2gXkivoX86e
CFXAEvuPO6yqNJaWB1QmKpCE7womQNKgi0jfNSJKsKatwYnyNnhfwUEtxFNAI8HB
Ly5bUv0PQ4KwO9xlu3tPRLj5s/9i5aH4Del99Mz04lSj0Io8KBJay66dMmBAZjrE
GZ7CBARTyhErMyvlv3Z/v21YrgY3JZ5evliSt16OwMEqu5b41LL4RL46+jYM4mxf
VF+4MsLogqDsgURTscyqkcnd/aFGwqtWURMCpTTgBR58W1y42Srou3BKCN94dOWL
ajWmu/j8v0s4issh6oH4GJgkcBijDz56HTk2u8el8fAowRaVOwYNTZcbadhyEBwJ
6f27AfoguLrs+2WeHJBTtWb6tH2ERs+hBROWProIMNBT/Rd1xe/uLaJE1hBK7r/+
37hd2bmovQo/vIhMwNrJoTmg+sXnvK/QVePVDME1CPqMQQc5vkDJ6cF9zYOTvFFR
VJY9NhtWKzj+Nqd8aRJ9NBmJNBui7cayst6HT2rdY7ekLUNABlPctU2NXm51myGI
+n8vXl8hNhQhz28EsjYBSJkAkO6LblVCmJG9fgoKVmU1E21+wBpsd1fEPehTU7Hx
a0NM1GgSeMaXtIBEdxs26croMcTxRWKkiA879sVW9w/GtcQw3iaZwnUr8Jnm9UIU
JNMDePVV8bPHwLXA3J8u1eXBiFK2jVo8Na2/Nze+RzvVdyy0tzRb7vUnnHX9qk88
zbiAFqMhxJF6LxA5vVm5HRgST2oixqDqvKQ6Fkn8tEJswI0q35S6kuFPqp07Flva
wme42dORjIFM9o3kROfNWSfZOQ5sEqxvEcsqDZXaX1P2jPsPUoty5ynKWdHp+84C
wM6cwp7h45VYePe13V6HCkoe8k/6tiNJaH3ZR8RTCJT6vrTNm7u2rBXEfFE+KOPT
dWDA7oN8OvDMSgauIYSxJ4MgBKDAM9bsWh/QltJCDLCYMnn2pzuxT6LYJCWH/9lx
1/SfSoU7HYqKeVnU23VOYIz3C4cMo8e97pf48mpg9VTCcqo/OPEjt6m4ctPzEJcK
UJRa1lqxCPL5cZSs8N1diisHJJqKCiwJKoM36KGKE6kcdmN3YxCwQDc9vuLWGy/n
zNCsapnbJVUjWlInUuYz7V/VJRdIZcsNe4f+H22x48z7kRa+oXz89awWn84qBCR8
nqxa2f7tSLrfOe+KtbPb1CqgxKvpJxVtzThz9cnjxKlBHagaLP3hlSms74xLmAFP
eq3GixOewET2UjLyfqWKYhdIvQpmE/yTGdDx+u6p1wyWxJxB0Gjv095Ud1ZmRCAw
j4yeORY0rIO0wWUOZ1W9hR97EJaQdsJgA8bGzn0HDMg0LDR9WHZd91E3HUqkZFPD
pZxCF674xZl2Ur6d7FGA48aNobNVhrpY0P6JBwoKDcpHWcCuj+hZaEDdEJFTRkWt
gRXLO/alQgQKRF5dvnnrqqfen73xt7J+S5eo1rIy+fFhPN3/1ab1tF85s7fSK6bn
0VeEaX8W4AjviNj7o0eceLUxaFH9zJG6LDbLxUNerP5yAsd+arxKbOglD8RUFa3A
GdTydvTeFaw/3BVOeBTPAzNO+aSqfZGSJo00B3NIyyBYtn/ssgoqLmONjWswEZk3
sQidfYixD+sm7tWuH+p6wJ+r2/ZeaiI3g0+xvpgh6dFa4p11hOM/WUDiypVTT7AP
RBjqG51in3hgR6BSutc//dUcUaneiDT1mCEB0/0Xpy3OSk4+aEfszWENzblYsisG
PLT2HpCo+s90n0DEqaMyrXd/SZ34bWgPb/+tl91zpDppAhE5l3YeAauHC7x4e8jz
Iywyv7H/vGdX+EHKq+OO6wIg1MnWHCJyIDPVvfJi70xTPaogQE8ZUgiccev1ZFt+
2Omt7j07iMNYLdMh0nMqb8aEqbB+rIp/u+tuBwHCMtXq7BEnw0CSW9F+auGxzC2t
MdY8tSxo2HbBcKUSh7mGIsu/jt/Ti/fJB2nQls++zCWG8cfSMIGcz2z0MAOAXaEj
rdjDm+qk+P4F/hHpVPZQL4aLT0BFkwVk6wdkFXo/WBoXG6MasFnxTk5mEf2Pg36z
xvolmhATwtHKXJlGxsJdZc2WxD2uFZDBpeJK3f2mpDtTjOnHN3KQCzLHfONMTVa9
zqSvJebFEtldtyxVEkLLSguXBHeRyQnuZPGnY0IMk6m4eiXBJTQsO3h0NBlVGX7i
5UXSy6Wt4R9+v5z6IYwhzoRlohKPGkpGeaLZU3EsVobjwdbYbO+Zk5XoBKEjQLGL
U4y+ekWusgFgQCOf3UJVxyPO13VWNdXUAt6HA4f18Qllsd4RNiPyr7q37EClEuR5
bCsjv6tkAteZoGSJQSd/8WomQJXbmS8Wf6j6LfMU0QGxC+fYd+oPphvO7ieY1xyL
KZ9/SE7Xz+MtK7eHUpTHN3qWpM3WEceazyuz4INzUVzsYnXX4qjn7C0D4eiO8kOn
UXvLL2kB0QOGmBGyFTVq9t3PEC6VZLyMvm3HLUtVTh6KEnPQtzYTvNeuPy67VLEQ
JQB/Tp9mYGpb0loukyBxx/XSp5GV+XzNVeR2rfULIyuHeXTjGpPR26EIgsrj/NeP
1gDyu3miq0p0fq8j5HTLig72HfyfRZFR+R8d59SaXuI3iWJpI+cAne/ISZv6aatb
9KaQKwkZvyt4brbUKAwZqVyk/8zdg1nvU/1zvOCaHSn6FZrtQAwBPJvKBYveevXA
joBhz0qKeMI9p9DoHw+fShsfm5cdOUSBrPVBKquyblgnPBRA9n1iLVb3GYuijnDc
n3CLZssjaLQq64jDZzS68u2hza1AvTn5zQ84sj3NRyTfHHLWIKDKxLgskm+uJMI7
1+BEoJCNyYveod4QBTAxdhVx19KKfb//2od8nOKWdLfmDpL7oyvSDxqCZi12FDju
G+ONzQoOQEFo9uCvDAHrLPl86Ze2OIxqgWusIZ8RGMKsiBfs+97RXniIYXCzbeLF
Zlg7w7xHlhXjC13MHYrgVbFIY1S8DOKKyan3fa5Mri2dLN0JZSvASfRcxGPaemXa
ES5ALG77QFKFzZpHq80OAsQYdc1CNa8AgIlgzMUMfYle0WwVi/uB2fyngUXCJup0
QcmT9fU4GZkQ/8VE0zJit0hYFqn79cueX1t7NuDjdeFv318dpONgJlcYHVhdSYHg
hYH9pvDtSSJkMPZbLpICSWb4pJPNaOUemEEe6OgxA3vpEi3+UtDjg42vOmPZUHp0
P4mtDP6nasQlYXGIkEBTorkJuENTIVqfRfttMx2nJB4D3wVAfijK4Pc2aioHZcCe
SjQj/jxqPwRvv4kJbkFt0NRU2IkS4f5NdicwSzWL/eVytkDXmDA2T0QUGsPwnKp4
234btRUcO28JER1hdQRSUkCpZN/IhYH/XPOcpMVQHtXZRrE1LJwpmoU9TKY1JfLz
2J3sk5KsQfUSqCvWwQUPEUln0hFR/vvBKkhEGuSQXWlihY20/seAXau0RRQnC05U
i2ZFAhBbr6Kg7B+eeKLZSHZWkyhbKr/w0kQ54WNBiPqY9jtJDMmvj0zRWzxT4MFH
ZiWUcUmz+XAZ3f2dUknhjgpj8pog2k+kT3OGSO3lVeCstZuS8CmZunYGIEsTb0Sr
vrngQ/I7YnTiNs5nUFkuvOOmbC5fQ2bHLAHza210XcPK4a8Bh1pn2O9bJ1LvaMG9
Gh6C26dMcAUrn1D+9BpI1Q3Ow4KENC+OCCF5rzJJrzSGUch8yl8zv98Hywu5kIvC
VvksaQTo3T9SkIMXZluS1Cv/cthkKtcOAhvoueInvMh9h9+tLawEzF1GKRtp0xGw
ODUt8S126IKYLEmoEjdBiNdGMXHSHpFZ72QilX7V3b/fLD7fTyC9+Fdyl/PdLniR
/64DviD3bm0bZ0le1KVnBI+xK201QhRQ2QwZtTHtjql1VXG3r+YZ+usu+toGR0i/
lrZq0DjeQy9EHZ1kfdm9s1xxn6B1Y6nw1QY+EsosdfwcgIsbgmXIF8C0OFaioQ4R
ydaJPnCEc2mLmykq6jxTY31E6uohzbJV/M5D+F6desMfWwcdS7pjLg0TQHulG9ci
YiANzeXXsEzxJFD+KR3cfr0FTCsLrpv0eRdYgkHFPT7AW5yvpL/xP8q8eJW0IPrR
ou7A4B3Ii5eNJ5FW6Yx7jvQ6Fwr8thKqwymfb1nz6aqoSINlDhN4fWdIDviRQMd7
8gygPSc1IIIrezhwLzGK8Yl9GRZCXSocBECXwsjHGvd3zMWA0PzQUdsAX5npDWw1
d08IGXMFS12KK2t8CJIp3zW/i8ya5cGpty8jzVg41yTHscEa22YQoJaJ8HSKNKEw
Mk1i0rSyiuX+BE2hDIInj8ayq25qgZ0xe57jfd34hUceBaMnxKbYsLfc19PgjKhY
FRPQlFxQ6V3lvhnnkYI/ZrOx/5lK/js+P71jV4vAKP+hEsN4WUZogsyxmCwhDHvp
4kkmCtSIwnN/FXHWMCkPt6etMPNOH3rs2wtth/ADDf0v+3udp0BH0jbRV4GEP7AT
XaPhqnuimwoF02lbeC0EcYYT0JhineiYDhx1UsWdIjuB/apI/sEzAKA6eik10pqH
ba7Hvi83eyoYFIMHgg2Wuzus8CUQIXDT7hXRbJ67bRKfoRc/ciP7CocktaHS1KW+
Mb7PDHb4volUCXkhDgW/mTIDGHYD8RRv8wmIxMcz7l9s+ykJOO94W4t9f82r0no8
/tW5NXbxOPAyvKzszjcWCNsugetnP9h8XoC0O5kvkItv2hXZ1ZSTr1kGLiX/UHf5
8dcqDs/nFp11kZkf3fOAInin+qXgXGLOUZ/S/s4N3lnzSglt54WhiXEnp+2EarYc
ef72VnFXMhufouGsV/26BMzUjFtOqB08389c6p2ACCU9sc9SVbvWbprak17hpyt4
nhaPUcX1hFXmEvv17v4yUws97t7dGqeVXaFHNsiEWyXpvafyPgIS1gSGwwQ21hji
c8cdP1ty1fL4LNaNU5w13NzAbILc0vL+ckVxePl7IhDCmo+nGJTyRrWC0yagdZG8
USuBNA+ZdMXhgnLEt+pwiU4P80J3l9Vo4qfg0HW8qOlnXC/ZjyqIjaPKmxUhKPzP
slVXYUAYh1QgfUH417BI7aOqBmkiOWsU0mgjm2GmiO6fW5n68MHhKuns7foS/Lj0
U93JFC/JdQbIPCsIMF5+1+yZuThgGjm5Xwku6kQgJtxU6lZqcsrhQY8SxYozYKcu
M8LBSVj6VYAhXouZVUnEnXzf5FbyUoVfr4NWj6T2Vffiexzxvgtcxt+2kOQ6iKZA
rHzcQ+YVHmBzC35JowWSX9t5QdnBc27xbAahMEjdV+df2nDRyidsIrOK5i43gCYQ
s0eCarYDH+tlzNmvmrA/ny0depdi/a1q2wpxMtgb6/xtlE1HPOn0b0m1Eib0sID8
vwcx+71tByOySWNOyuHvYJvss8GzXtcB0yiFUkkjsNRHPFONzfFm3yJPDYf6SKoa
zqEO2XptwE587+Kj8iYCP459c+VGOkM3AP03PGylrgAIq2Fl/pgpuxH8ee2OYekV
rT0t8PinewfIkldDErhBb2To2Q1pY0Dd7y5QhgePwyLpmJAn8Y5ZHA2SeF6dZG6i
R1GwPF7vJSX7V8Zey+SvAwXAVIUxkWoBeCzXNWciAxAW+wLJzAfk3pYd/7ahP+zz
peYZxOiAuyg0hQnoxpR39VmobU/X3vPq2xyGJPd8OINzlgooVSp5LJjUGthixQV8
RUUwEuiQBpuqUMUoUX9eEjWx7O46y4Kf6dzQDZk/EeVYrj9OzoRW/lYGk/JNQleM
IalR2/cb+0fMi0eYIblC5BDgMTXK/vQEsFJM5H6/JV1f9fCvjcdc1FfEbKPuI1LE
VC3yzhNSLic/RwPAv9tFNSaDsGFX4MJ/EydcgVpFmdt2r70z1e/s/FssqDVrME0K
IeOWqLMYANrVz+yNAOEEKndkXWo+t0gFPFxo03FTn2zVf4HNptLNdIEJ/BPFf6/0
fhIdaJXMxjPfoR8O/MANjE4ueb3n27P+ryDIEVwWZdVbYofqT6/f/N7ZYOd7s0g0
X1y46Xjd0CmgWv6k73I4B+QCj4NP7pjrM3sPLOublMDHLYEj4ACGLSnr77UzRCGz
7o22gFhenzlW8XdUSFnGAXs3+iwnrR3wKvVCObpOCmAB6G+yuQBHK2nBHvogcjSH
3KFeUFGIqDExpKkPaGKMTWekeSvs8ea+3ChqssTOd8TPth6/802qJEfaVAXUPM9c
zG15Qm2tMPpb8XfPPhDQM3z8gF2Jy4SclB98WrV7i/zzatnISa6stHgNLl1ueXCb
0sF4nXMtkMP3NfSa4giEEv5HLhVvTjiajkP7VdrNvuMdcFLcLwajTo0C1lltonih
0TUpO/leXoigFCfwpwsd5WbOFoMIgTPFIP7oFMsScBtvwoupXcMOAhi8PTYTlAoU
Cz470UGkSLMnvS7dA6mrEywJQaVKdKQUo3W2Ta3g8cnQ3C5J05zGrJoeLTR0mS+u
cwP/frWq8Gkx6+i4ho69Jctvh/eC1AWg+eewpNbmcq5EUevAxXVbFSJcjxAULThQ
z6xh5eRTWExMtgvAz1ishHBTiB0tn+2MOBaA/gW3sOLBfsgIhOVHSOEqczPfLHLZ
ethwVk9T/XZBgjaEYKdanWZhM2V5BzwHmcFZ4o42DxZUiKHfhcLxZuVBpRgp0ErU
+n7UKckSfE6EXsQx93Skrt3xF8DX6uiwgO4lAkFLj5HZIkelio5o2NESzbzfWgEw
DQbwhAIx4/DbAok9u85smWTjHM2tWiQgi6nDjKMgs6mf6UqH9RXxfVdg1CHyAn/m
4DBurNsGiVtvQbE9kPysX2J2Yu6oUtgVtWXvgKEPgBJpnKGqshkaoxLWR9KR6hNf
MvWlda5I9oEF8gQsOiuaGaERqDemmQEPr3ueKgtjHe5XI4JoNbcue1k+HMlPufYg
juyac6hk1546Xbk3AC1ulb71ZePx0xT9ZOtPwQXXJ997eWgXPIdJzW8JzaRT5/FC
RQ2DggZ2z39idd35oIUNuhQ2jnr1Alw+hO8v/W1MER1oQTvwcLI53FlD5bEMNDsp
D0Jfy6ABK/cOsqSfTaWKAFcdMQBeuQoi8UgZJZaNtaV8SH3yzL+zgtsWZEbzLq8i
89yQjTtZaNj2+IctAYIPOKhsln8uQL3WRd5CNgJFbm4YnUmDIbBCjnhsGOx6bEiC
Xroote08d+efY0zBa2COhWeWM4l1BS9AsRobU9fnj4jn1fYcPx/ZyIk9qllLc8x5
nGB2zpiMDywpgKB2jyR069/rEjN+oJgK7oIQeESBpZxxhSOy+KE1onZoykr5FlW7
49ChxY6/i7AAmqSI/YJyyT9JBQfsqdpZIIQYLWoGffDtouxsb6OZ8mpSwQK482cG
b4sUa2YQ3SaTvhFI9QaG3ljKNVOY5FLxJ01zM9WVC3kTju1EinI7xQIFMeZCmkg9
b4eNDRqFLfM/P98v+R7/gCCqhA9mezQy4Mj33UuhRUlCr5aTlSN0SypN6QJVvszu
X8P+8ls7S9bKH9kNWSeB67bmCrRQyRLyegNZcOZfG28KGBAMHtn4NVua2H7aWXjR
emlZRYWwCgpuyZ8ZEaahhsSIHBty4++ntMdFCVDnGpCPG6AbQ1Q5OGem25mXWXsL
KvDGw6wnsjDYaFbmSLSxwa5d4S/li9gFAJxdyWGOZw5Lu/cisDQVOXOQ9KB3MBuK
dps9BKMLn5WqoTsWxPC5cV5FFDUNmTR7eIa9QnSEQY+oA8MearMj+KoDMh1ui8yo
Wq+imONidj4eGb8Nam45S4t9gNGcjFWHx1SdLmQeKJPmCFuERk1Gev6A7RfuaZnZ
mbwhDQaKTvZtLkMHDNh54jff/APnCxCLkLUwAbSSiT4ByQAS1+sHhSFlBzfsBs1M
pOT8XtfG1o9CMK/V26y2sOI3Q3r16NTONBt//dOaVogB4yBSGDDmMdRKkYRoctPE
5tYn8hqJiZxj6Buk4Yh7ESlyyqHXMRo+Pje0pa65LJ2cCq74WAqISgUA+F7gpnBF
VOe/2P6tjtnoYhuZ9ZH+kJAMAC5+N7NGc57CKC/9RErJ8u54k7XEPNyJt2c97JZ8
WW/VbZtpIFpsui3x02OVQhXYs/V2fsYAu+6eLz1NLNUBKsrOUx/DC7SubKbiun5k
TDRsBxhUFiCiJgcHjFP0i3CP8XARn1LvO00DIecU8Ti8ce7mRbu1EtTdUnJDgTKt
tDLHRLI6sc3Affq/Mu2QLJ7RzgyEwE05AxJmWnuDlJV9s5gV5eSm69BUPHlQSJmr
4DcuERUcwss+b+hJgGPXM8RWCmeAa/KW1ssXxFcprNinNZjlFBxH2cbQiw/8ezBZ
xhrgqww5DXB+oLo+j2U834KFZS9Dxx2GtT6J9L/Ig+Qrju9FTZ8ghOD83Yl79M03
Aj8XctaIju6vQvcY3YsU/4w1+/sc96Vd5nkrxxlja5W9xGOc4azz4eP9zC4s111z
9dRu17PtG2FUq3XmBDSSqPxp3F5IbH1/zQ07sFcI3185LqD6fJdHLHsTCM8qmUDW
zh8jIngox5NI62hGk+seN+rGmydTfOw3dUKkvZdw3iVohbv4FbXMYqauhvJVRO9r
//5jXQ+VFW0ZdeffqZ8En19LUgoAC4smeojA13on7XhLnK4jwiajb2dpwU8WkG9R
QarHc62EPTWl9Rtd36MCmlL+Kc9CRQPDDxzPbQztVUvgcEiqzrbvC8jHxTBkQ7dT
FC5owGpBqw5NjtYSl63vwKKfjlJNBdX3BN6NGZlfa7Wr4YhffBecJP0O9QpVvYjk
SYRSLI3oZ5OoKt9xMyRP2Cyc4qsZFDYyot8qQLBpfbzIBNucyXM8+024DxmxNsDt
G6gBhDBVtd/G6mB6D1Jd2yAUhEceedzTxu8lNePhSoZlg4E4HwBMxXeZ9azlWBwE
zsmBsgqbAu7F+okuJ5oNTpYeNqkwesjzo5kYSP9QD/OC1qptFYyCtkhMhLxtd/is
RMC9sVHHkgq01kceykAVJr8G19/lG8NyHWiMAE7dGp90fl4L8VpHYow5FY6WBrAE
cwjTxMW5UfUoy0XyEj0ZNOi9u3vufFK8Fwb7xJY9PDQI+jMWo2V5TS+gUPIgHwQX
Hz2evHhf6KBFvMUC0I4h4wzLiHgxANZoMzldcfkXTPucxHfNoORnxaG4Qi3gREpg
gdfwWGBOE7pTvzpQwCgqrxULxsY43QomLyzv2cUlHk0qOnsRVWGJa+TGYtB52Xdc
2Jpi8kPNVLl6IfzZ6IgAifqDcc0OzKyqllhd0fWPm+DfhP/CybWG4zr5u5XwT2ce
Yb4Ipz5xlCKURXsqzcUKTZRZXG2IB7Xrxt6MG649zicuHUaKeU2oPbnIheCHayX2
p0/GBWw6Ac3dJ22fpb3IoTm4S6IoVBo9SD14CGh76LI2fJDkIEu/MxCtoAA/lvrA
GRKuZ0PzNpeWaNalqXzVHDHtwqD/XHynuZM1CCXvsJhEHEeBGtuG8qIu8VFbhEyY
KoECGzNTz8uf9Ilz9YLljX171j8g56Q820OYQ9uGXHH2FxCZBdvEloP56XvM/Tnj
GoRV7aSnR2PcARg9gWUWcZWfb3VhS9i0P2n1mYOsMAyiTk+Jmi9veEWoqj2icTSz
b1IxcyP03e1bLiEhN6DVDTid7n5joQUphdBlx8KPssJpKB0P9BRBtqwCShKl8FXo
p7EdhDAuCdEb3AaoeC8TSiqokJjR+AwHgyQTuSZJLtgq+XG1nGgu0lk4O/WeLgkt
UmrTcd6ogNScSldYBH8IYwmXbNQ1o3GwCyq7LA3i3BKXJNYkJmHUnBuMhQUY5CfQ
eDzFy0CMKOBL40EghQQPvS9qtvB5bLmkp1NGzbex+/SNnd361KRorCHOKWA2quuR
ejVvWoCBXzPaAXphFYhlhkMLprqqLj+3NfAG4OypeyY6TiIf+bBaAbgMnvnRgmPb
vbeUSu21+20Vvpip3zRp/E6qGGmMCBhLVrcfGQWbXoQAvbpNk5fZuSIxQSEpbyJK
OTVlrCUUDRHys/TQ2ySHpa0VMmZzvsFhPhE/Nf5APXrecRJFRpItG6yTKN3Qs0ZG
UuBsh/FOR5LISHiyge971kpT78gf5+FNnXCQze3Jd4gnwW/XXikeCioJnxc/Zigf
uq6SuOV8sL2pg5j9XmcWlFrteMJldFsiXizEJ/ntbYnO1UBxszgiivsY2WZlYx2I
1XkVXeNyg63UQS97cnBBJxiBHkjYJ96k/HkbWkEi5g679lX27nZV5Xs/IvwBRP0n
RTXMUUljmw61bYfGaDy/ERZ56Ob075SvjYwpHG7YwXMbiDedWWLvQFm62dOiFh/t
PfqBpMQcueklnD2xL95DkGSZNIxQE1IGF1HREC1USs3CN2eIRT0sRLUdVdcXWXtI
x+t7/o6tUVV1RnihsOAn3gZd8uYUHAak0cKfrzJfQG3dwcSp8K6/vM2MKuhW8urg
ha0qZe/bLqhFQ1uO3xs1dCCGUVL/zVM0sTw2lNoYnjt0sytlDIywClns5oMF/qi4
rHFCCBm2svwXEAav6pPOoxWlBn5N/FN2L4inLlL942BVRv7gZJXy3i+KNyHqjAbB
jHYzEiLNSnDzh6VBRUtQKpFpjTC2mWZeToUR61HQYVKcLCKMUd4LBrO2bWdfQEn3
dnN/gnxlbBlPta/DdhVpNelPLm68fC7t+qasrI8dh00kQVDN0fiK8iFKaEV0IF5p
ehWHkB8R6KO71JPJjuPDx6gFSgBrDkbpl123aN9zjiW2l1oLkh+/+btUx4Niz312
Ef9aSWdw35WXg8qnkjtb3dZ97OOyTyR++gKXSn1l2e1DgErhheZ7fNGIVVjqr1Oh
OA9ym9niHwJIy6c5/1/aNFoOorcqFLfPUYXtHuJdUJbfEPeippG2otwke+DZ3AJT
QdMy1Wf+MycfIkXhCZ1P7PrLvb8/UFEBNKMDsmwWvtdNQle1+RfZictycEDurYw4
e2Pa/MzBdoxDZRrcrUgjKUgT0fGZfkAiC4DQh23jY3xUv3Ti/6IU55uyYk+n+1jl
nELmX/fnoeZSbuufat4TuL4LCic+nLD+HqJwdS2Y0w/tAM93qVbi5Q1YyTdqvMHl
pX+7tF+sO1OxO0OgOOYJH+mxIgK4Q7T3JGu1mMt90N1LwpbzJat8ttu++56Ta8TP
aIFDX8ii2QKG9AhYquPV6OyqdPoTMiHbqaVBzqKwbAldwnJZ3wXWMugxt6KtXqtn
AikP/06Fe5mZ0v3YJGjg1Ru+s/YnBtlH1Nngi38dNZ54TqNgGKu0de9/XjPO3hPV
M9n6uG0O4sjHBu2n1H69RgCDX25PzboceOt8NJd9AkuqXhJxKZu+SULM4ZyPlGsT
fInMIAKuM+9PiIjp6S30nViunLYfTFQKMLZbLTFk+J5BDyjgSM7EAEvqLAw96dUM
SM9JA9yoM40iuYpyuNXHTzdpOaqAuPSuBWyMhcQklJT3ZbZOVsExpZkQ2ApF3wBW
qkCMwonThtDntlwVRMukrW9iLs3qKtFyUiWnLXeIty3Dz6RxS/KdRyeUNXdkxT+Y
zid9f/QxJVpZ6Xt6uL5w55KPjIdzWkgfvgBTVcTMY6pl9gO4kVAIQOB+egteKiMY
3/Gtx5fRMl0O5nr84itD0ySGBb8FITAtx7gQDrBxYvpblhH6s+PABxhpp/BMq+45
5Fuhu507SeTtVNsGc2G4vpbkEaGC/68k0B2ddfq69NzlyQOsv1UOlFieJmolV0gR
VxWnjMMpAoIj/lCLybbyMCKWackNIbZWQYtWg3Q83fSeGKmA3LPnlp+omOEJglrk
ArCBAcv9kjv9z3jaI0/8CmZXh+dxWGPEaTDUIdMhkDSEGlDS1DzZs4gOB8lrEnMU
pj3YibX/dft8BWcpQo1efv+YVao/QWP+hFVcBTvN8Sbi//OZ3GzCmIH8xIb22zZM
VSgYAXFfv3SvG5y2o1Ssfno67lfCJrocNIzSEQVVHlnQzeEk/0/eyc3hu55Yv08+
aQ/n5Aj7P0MA9UVmBtpO5mzjX2yagNEe8I6fu1aw2hnxVu+p/6KN5YvirwU/puR+
SUagWCbxC0PswoCStzyqSi/ctLGaPSd9oD1SC6z6Zn7racqMC+tHiLgOjGJXTJ9s
eX2S+HQPEsJFjprJEGlpsHgEhQSfYNL87T0C+iTbpmRkE+5hdeDiJYCfTttcFCut
OJf6z2fu571Hr2e7Q/l2+pKDbvUhgoHC9381hHkg8E4uvUoxwt5m5iYTeOL08q3m
TxHy67Hch0qRknMPMo1h7NUKch5lustNreKbM0NDcOntA4ib4zpbzWy0HwkllhxG
rgtieHo0baZOtahK0OWUsawtzQs0V9pCr4huymHIb5FtkP7YLJrpcPQTga/xnj1F
RwEV5fDLH8BwjD4X8eI3yygWVYEv2tk20EHbz776LA1lJD2AbFi5zxQ7e5IYRzeK
KYozbgAvwcSNQ6LActQBoaVO5mkBwkOwca2PnDmNd1HBYGh28eJmZWlYymuWCx7X
CNd1DNEILYzCHl+bsYJbcbNRu6lxFdceyyylGPsVYz4qezJN0cG4pZjhakwoKWtW
ybxo0qw4l8BfHi8v+IhiJ03vP/ZLennZv/lZqtwA6tMfJPsQOm9foPKUuulPIQJY
oCEdm1QGQTgJDaN4Upngu5okMMgos4N6R+ar4C9Wz40pCTRxEogTYig7ipF2MmXz
l190c5pI8mMP0/m5Faw1KEd192PCmMhFwq9jT+3CXuD4FhhQphOR/kls3dpAyv2x
5MNyxXCBeXRYW/TYn3KE/kGyvIbmXg5m+1lpqEQDtG2yKR9flKyI9HRg4FZI8FV6
T63BGBundoigabJvozCEjq1nXF//B0VvDRiTGbb5/mzqy3se1X8IY4QN+C3BoH7j
Rsj+i/9ep2xiUA6CEUxqGwXHdudWFzCwDf9iP8VN/1vEYVyhblSPGiTGO/TT6IvG
GmJFHWNrQSzq56f8rTp8LzoKt4rDy2pp56jsV7Fmv0RJYcAF8Tg6zn3Est09KQij
8aF+kOIamrvH6yBz75sTWmLkTC5m44yy0YMhj5Aj5R7QP1HXBWgr+DYm6E3wIXRS
ZrFI7JG4JGdmXVlfVbrHdcx2cXXdINxhKHSBUPXDmwxK+3LbtuxR7yZRzlNVJdot
5TdGOdfuzN4vMemWWRt4XEmi19vCfinHVKiBzu7/e5CGVkK/QVlcoYMBQQ0nshS5
0+DORkE02CWCXeSe8Br9rwlyKTIaEZSCFoN53bWON0w6AZsFIxz+CA+GryNAtX7/
vF6MsGuTQbEZxarSUR+tqZuEYdiOUKWbmzHF+jQf/sdNxlVvXgxmL1V5asnR34tS
79DT9ao3ur+vho8Vb/JbTiBMM7/PyNW4vm/p/r88O7QP07nlSoz9VxEc2EkMQr6t
NOMXl50lrlzPOetsVSZPV7VKeC9LvxECgIiG6Gbfl80dLNbO4jPbblOTvYHPikNL
lGnLJspsrDZXEBJJpXPYm5faDuzwmN3riOZqh75gZsu94398tqlezbWQYCxeCzdu
y/2FQDdKFmLkIDDnHVRr6PfveecZ63QU2AphPnFAiUSs5PjDfXi38RxwRqdqqbIK
rp+XsMfLa4JtlOyImHarJm7R0F1Lp/2jkAzM4KGDsWdwgxOqw+3P3riQAUD5MzQf
yVs61Ib+QfVxOvJ/Vbr5PMU+9QmkX5M+S/sNp4qbarSC4UZ4H53fo83BYOAI2aaN
mc7Gn0gjPTldpFUmughUOZZkPizE0h6/sQQ4yYVAeSA+6Oh8qI95iWB7lULUY75P
3dtPjlljWqs9vYmpJAw7b0DAcfV7Y02a5+3uS+I57c62fUh5W1ZMTgeSLDJRffap
uYYja8GgYMsLRaKSYgimFNpyBWMerSF8dxhtnkOWrgb7xELd54wRDmJsFT2VziwT
OTlpDOmXzkA2Pn51HV6sMHaCbMKhqQOGOK3LoUO3HV/4FJ3M5ypxCjwNGgzgCB2u
AhuvU89OuRYMNjz0d5JhWGSqqEaGAHIriWymAhJdOKdUBjqGwI/0ZI2wLbZWcwzZ
Jt+HBXxImtvmO2c9EDo0/ZZLNh04G7jue8ELQxoB7OQCkaWKAKSl3SVbCtSa0QfU
PoS/QR6YU4mKycPEh1PUxFFXALBtx9vQ9jVDQ21qqnG/7R2f9kGB/SygAmjQrM04
nDunU5KLpXVaThYg1690EpEJrVhcPdLUNl1PwZ3l/mgtX62D5uo39ifROmviC8vL
XPbAF0slakNYzAGmhiitTU99OVpTaEMdvyzovb5U7ouy+p9hPx1wUYybI82KkEdJ
xMAKiVQDn6lVXFgavYoa2cnT/oqdHMExffBu2G0ZEBkXCQz2yzcOlKaVdthAqBiE
fFWu4JTunfZHK+6o8jPQEXj+IJfpMOsp6ktSI/HDIqkvkARVO4wyzHO5urEhuewD
LPuHMDfoZqYfu8/pF5VBYWEZTPljtYeGWgWPeL+3r0l0zU6+Y7Wseg62lm96Krv6
SNUrQbQWRYXtCyATcUy2EdXPAYGm785C+TBezBhtOuD/ScAyU/9r+E361hgX8Uis
0hgyHH2tUHHVuxtAJGC7yWXXvNnXverf4v8Pu+hWaQQ/GdraiPJBgRo3Y4TZ9yYk
WCnus4xqVF5k2N1H+SgK/43EtHZyNEHm2FJLwinbBMa8oe5OUBhf+yJH4vo0KDMm
Bu6egPavHWFmQk2o0w/hk+oWYfjZdeupBfRBHVrmgNLu1jlMKLHODw0Uw5ziAA5f
iv9fv/7TyqfPVD2n1iC8ONYF1onzPuszre3Mp6W5uADQXvqUFZ7guihDmTfiBWtv
1xMDE1PUq7qREaQX+P8DgJih+SNIp/1kL/zrckLlBh0Mo8MQJT7qFyJOFGIDuPjk
KA3R8nwRsKb1yuejxsn8Nru9L5lh4zG2tvMupWXamUbuHvs3KBHZ6HMLm33mc4Uy
BBtlaRRbgBb5Dscatba9p3t1B8IKaSJVJAcFrhr7gv4FxzFDUhSHyY9Ys6vDjn1K
Dqxn13r4XbVb0UoleePPqcEzFAnUhJw74Im4BV9opTv+HaK2gkcuj7SYIl0QQgt1
js0v1B7tKi/kBTyzsp2prG0GUbXF7O4SLIZJIzWv7txFNyci8I4qZVJ61BiiA6fP
SYBdo+cmHqqCErs7S9ineVpYVue/TtCzVpKBVC6agyLsFFyf2ymUO/zq4svclW7v
cynhaE5BOG0aUEhIxyKO3RhDJXoD9woK6pMzrqJyQ8oVWraKeoMmtw5+66PcVRKQ
2bIL8A5HVMpFM2ezHisgmvo9XJtSul9R2PGc/KutJ2glIw2Ds1vDr4OCt6+RrcK1
Cho+mIorpwjlQpWw07N6epOWqsF1kWqP05paeQWfHAo8nFPxpZctmFNb/fX+WlYC
zEo+ZJskORVoG2FXZc8YFiIF4xn0FXg9acV5xcb5WJPgU28J5Eiaowe3gaDJEiqS
bNSErx7NGrP7ATy/KBEevFJFEemMdxM612ezScAqR7l1BM+I9oJuQ0ow2bJwQZ8C
NL3SAs83P6axXRirlhNFaXMZhnmOWG/6RjPDRGWJnJOXlj+NkAyH5K42CAbVqzR9
uxhLFJv05ylgxPmS5OskNzVRBmMLLqAaDgo8b7Y0/hyn+FF/4xgvqm6l3S9s4JwH
wE/ATZWUdAV+wQULv6+JjKIoidQapxXld6bf9CDf2BZLbqVch8W2SBvXdjq7wkck
+arXVgRGm75gU1bHoRwDgoWNQ1OojVem8mR/gJqm4FtzgPwW/erdif/90TSqt9U+
axGCJmHHjppmV8sPJoI7/nqxxb5hT6Vjkmr0s6OUMtBN4dgd4oafpfA4yajRB9f2
8hsXLcMztAqERcyytfJ1LZ0+SHkDZNGqKKslFD+kuuUKiRZ/lyJIoxdE3qWMbhgu
XgBc7kRZGVQP0m8DNf2izdhNk6eh86f9PwoJU/gwZ8RayQScOaKhK1Zz5xKfM9FJ
/YQaYYMlOiTjPiRy+8FZmqjnKDbnTBmSUKNBLxeu61iKpcMnlP9ruUo8gkW19rHY
CMdhhp462rkXsYa/nIRWsyEgWRAll3adWm1YUsmqh7mgbLS6WmbUAeFyLx5FVnjj
H86g6GB64bChj/kLmC5sB/RbH9pkz4sqLXlPKz4lc++BsYLawxR96ZkuyCt1aV1J
wEcJzS0u53jgpUaWIDhBW02BMyC4OyWcxhf1NwBGLeuyDNo7LUwxfCFUwfZjhl8J
R7XyujXBmYn93O2cjuKgdPUjoLRtQtVbzTt+vTwWcAj3QjdplP5ZuJcW5YdJmnfa
UTsds6FnVzvoqduhyjhpdhixpg6m530dji5N10hXTfYyQ4l4A1C+hRt3rI0lluuZ
bQAJvciQQj0AFMw1XVMs+G20Apo92bT7EYXMnEs2LTjQNiZpOhCNca2AJzfESWuW
I+jzRFLK+Ryfcut+akml09YP9OT/NJWiCSRSSktHkfvP48b3oxcsolU1R+m3U+uM
k6EAOCuwZix1eSJba9HOAONiGuOgK5DjlTcjtXDAakZl39bZx7tEO0IEUoG9B1WU
FFSD/DAIKRszabfCrI2CrAO+me1CdnwTWubIA4BaSUBQi9nHwnRq8qXmrC+VVUY1
rp6uZHyQ7VGsBDV1kCr2QSFZbH+Ry/glUP++FjkwqNR2rHD2nMFQ5e7F5jl9kLX6
TTiQ7N7oe+yd80PPfFP79JgiBjwpQIab4k2ItbT0DGmiTkI3Xs+iDFgyknco33g/
/F0onw7iBShCcVVKqnxg2wlSX/9x+75vMyp9jHc1shHK1Ym/vXtTA5oQVooRslM7
5q29z5dlyy5UZMkbjhgRP1JNSB1Btuf7LCxLOWjqzQsHdKF0Yx36rFiuyW0HMt0q
O1lTkYt3nRhpAXYBmd/r1hwMlDitYfgMoZbDoyDw75lyPVNaNRR9oX5kIBwaHu/4
rnUrY5yUYNtVtQo2RbH3ulNbo0YTAbKyLH8T4LzrDTL1jXaRkl8L2OWUzi8Fyaai
dmkK088cYTP1F8fC9G0bCTtjD7NleHz9Omb1U4Z2OSPExv2fCLYGY6x0X5d8ikzn
tRMCVSIvrZpdQqtTXO8M52EirNO0WlgaUtbfgzgL/+thTr0s/3Ywe0S2HVniT7d8
S8JMC0y692f2+0xabmS/b5GkUwj5+fh+wabijdFen9CGKALvP2BKykIE/Ua+brsZ
LSSsWlwwpEMDnoSG7cPGDBTsXSnqH5YEPt0BUs/EKwbINkVFetIXrtAR6p5k+539
yBVG2coi21vjYj9dWpP+iEcE+f4S45oNBxPN/f/E3FQL4KxSFbM3EEdYlGRFWQc2
7hqrT9G+4jdFBfhpZ3DzZYYKgfjj3I2Fiv4LIZb4fq3iMQPnbjwqV+16CeB1EeA4
iewGTBmd6Kiykf7bA2e6s7xIG4FLg7t/c5MHZkrp5CLs4oY9W2OnfCgj1edkZeBU
3f4A1EqYcvORgqdgBx9dYsY/QKUNgonFyxCzN4arCilUJFrOuiLN4N3kpT7gXto/
fDVe8dOWCIPVht00EV3U174vKk+Qgw8ucDlTzvggLY16v3+bYJFk+X7xPtP9/LZc
uJFr+H8JrZZyCWB1TMRuJ2dcXlvvdJtRjsDRCh2GGoF+JRLi0M2K518fPc6YeY1N
c6at3gD4rwYztfDOhhLlTF75ZfaQMC3uM8EnYYhOh6ikVINS543CAC0p3LfFKDcQ
GwzKGJC1TaU/bMHc6sxRHFZLJsAeB1WY1B0DgsymLtRNY5flpwaJ6LitqeVosKqi
nMkn9Ss5Jg+xjfyx/6Fp3cJ8pY1rkqAqaVXBfyhoOmCK4K6rl8StDdqDAkK3C3lf
sLIQy9LtPdJ0/mXmDjdz5qkogd/ZW6apZErBpxM9a5Vxa/J1W1k4w4/rCTn3AVci
nY7Hd5RBm/xDcxqOvrywyc8rKPli1xW+Xpa01e+pqmFopIiovZvfNoW7QEfNuLgI
zA3kPAydL9HqQgJAqk5xGe0C8cnHgg2CXUyGMl2E8ZC9vg9GCCH/5BvQQjRjpW56
y0pTdPd+KbXRuoqoyLy3yCrIaSTL4zO9E36GvoD7iWogUwtlcOIacc0+TIUngbom
UTkWxWwpRzp5qIyheFF0TbGrIoUV+pmlsS3JJT1WCaGBtirfy7kUeVcCmRz5Iu42
mqH/20jzaQG84wcNGbewqVctstcun+3vK37euRIgmxpk/m9NGY2X2E/7SaqsoNma
T0MeyfL0SspPMeHMsTe4caTNpsF8BUzMipLVI8pdh++F0otVc8x79OLSX/Uc0oas
SJ2N++vEgCkh4S9noGqF3vGRTbzZlutrMGHYennYBKxXPqnmssgkHhhsa4KAsoFm
h+J0mBW1rt0rlAqYKiMm40inZF5euAP3C2zMa6LO8roXVVVABeCaLmGtKcXm1hbE
U8xa/Q11sB55cM+AnixkiE3Vup7wz2OQNd3apEGdSRBPBqSNpJvxP6G0ZYnqdpyS
k0sv1V6WM7mFcJ3RRDRRmk7r0mDGS3MgR9uVKi65nD7nXIUVlut/Lwaau0u7HswO
zqXSMKQk4u31mx8jcsPhCzlAxb0H3gVUg4+8vKm0V16PYQQuvnMW6ZanX2iP2q4W
sRADH2LzbvnUVpZ4TeovzMFTPxw6yff5F3035ai1MRLRRepZQarh2IGur3aHy2ai
Gia4XTjhxX1YjrcqTh+Kew/YEgc82XpcrzqdJnU1YANKWIryPfmcY9YZQLREEG4A
cZvFtE5JzhytRH7RB8XtixDa+WPO7dL2t0t+7NEMKwSLJBP6OLeeIcfOS6QC9ane
Qjkn9dFZEAGsMEb9WtPwfj96lhCDNhAoi8BCm5/5UZN0fL3GpPy7lI/JUdokVGCA
FVyu5s8WN8KkJHuBAu70zySI/qMkiLzQaANhDGnwqDl4z5FYMt4GAzmqid4rQwmG
J7xMJb44BhIlwlicCNidk4gdavko2nIRylj8xJnd56ggw/cvgpJ4wlmFRI4h4tpJ
IpXEkNGDfiUmwOzDnrMHwr9ejiREq7YlEUgskttIin/JAefZZDdQCQkanEqlYt+Y
l925ZbdkXQq+7z7CEcGA+HCkHlO5OIG0uu6oMoSXhPCDbYn/ynsL82XFzttEggAh
UoL6KlMSg7v9IMzQ0SUvHFLMHVbXurupucDkCHNuT1vsYMtFXeWeWy1jb7s+S3ae
ILUzxXTWDQrO9os+BUSs1EwHhuZETX/GN6hznPIZe+zQ5goZLfIKnNGiUh7zk2nA
odC7g/26Y828LQ3MHvP+Kgh1BkwM2Gpez8MCzjfjKk7T7M1I8cH71Pq82Fta1xgH
aLqe4i7SZ3qVtOZOf4YR4TbZiW2oaj5pVpgW5v15GbrU1Kfxff8QL8K6fN8HhHLD
ZuOzvhpwcxNKL3CXP+qH+JCnahsvxi1gBx8cKi6+1wY/YnATG0Xpa2RClzT63P45
Hxlv3+r/v6Fdga5ouD039lRY1Uz4sRJvRJNUHiKkVpYp2ccZ7Aiz+BidPUZ/Gi9o
WoOzbOjQWAaE2NCIdzFOLpqxnWstvtunnNlRRY2f30wEp1Lc6ZL5CQvTDoCuDpKq
3eFLPnj24buymDPtzfvAyei6l6w4Kgq1tknH3htnrcI//BNaa/fBTRObA8ZE7xkD
SuYsYSrpjpahOlyeFaTOCTc8K2JPTkp1i+7/A425l4Dy8IG5ha76LJE6NZl2Yve/
lAbK9wT7v72H4kxPmzZKAfEM31iBqHE6w2k9JgASPK7As8KoFqbXTPPF3eDshGps
swqfJyYOOCQzEWulYh6kEdipEA/CS2C/KSlZLTRbR6xfUeEg2SExt5e5uMDW8wBE
WwCVpky9Kz4bi9ZrdzHUASdGqKsTY7pgc2uZ8zOzzwo+NuGDRVscZ3nfOr7kEQJI
HcP/TpVO83Mz5IdxQI+jDNVj0r7socTfFmNsLDMfFh7BqW8Ka1fokMNYeHcWflcn
a0hiNsAhdey1Vf5MGYBZFdVdT+4IIUjPnnc+sVdFUl7g2E1xa0bzTMrpSgZy1IR9
wjp7kGAmbEsD377G8Une9cPK92vHasmkJoyWH5bI6sNilt3AYRqodcBqsQtKV7kS
ORptxvF5E7ReuzFVLxBG1UnobqGDtNeu6aLaAD55u1idklNHd6uEeYW4hfIpoVmr
4u0pO2lY3S5iM79Lz6cFIS3hvO65hNaQaNLkGFfZEpGBpOV/n24d/8lbll8MsfEK
nLC2CEU1LRRnSF03aTKTbaRAsIqGx2p6XnJlPQCfYslvVf/GOMw9MjSovEvzn6Ny
BDHj0KzkpJ07Uv1esM77CipASYfNFeu2rPffL1jomT4p9FVui+HbTRe8iaNldeaJ
YgzYm+bVCQpRDab8QRnl7A9GCSGFXuUhMB/p1dSynMy8D5OG1FmL1O5Rzja0BVd4
QPG4PH4oDJfrRXFvoYZIVdvdeiIT9x32KcJDD9/BR5iYpdQGoTbDnrHxD3F3cgtG
KwHPb9puJjwuhJkYuVXshGzLf7EAo7cJGTuSkpmIAduwdx2aLwLR4CTFAdlypeW0
mKZyznahB6Tkz5KgUZ6GeibVRA0VB6tq3gU/kQlmd6wZUfL96PtyHcJKfh8wsrag
88ShfZctRkNfA1+X6X0AW/3+q4jWw/uLo7acPzCCiNnTkXwIuP+v7V67BMojJKPH
FOevXLukwRskiuOex3cf6Ba54CVf1a+pcmakXdWh7YLo1daIpLoGuMm1PTxe3JXf
xvV9ZBZj79s7Q8J/mtXBIjTAigIjUx6WmBfrBN1V27W6SECT9foSWESJa/ytaaY5
6YtATaavZ1+dO/g0/wL2nkcQ9giepnGgLNQwr/3t3+SWujAYZx2DQRFJdVPjTwwR
ZNcD+r2T/U0jxUnlaQroaFBuYAWhXLPqrEK3LR4uFwl+qPpK90sg8ocD8roF5v9q
YzoleUGpXTuzEQmTyF+DoCXirKJUHTQ/SkOlJ6wdXsmmHU/MFTiYESNr+wXr8IDn
iwVgU158gSKLl6EiBYo7kPxDiu7dC5PuiTX3uK8ypGcPBpo0a2QqBk/LrP6vQYFq
/ku3zgV8I6aE82FKbUPf8gMjkf5s91bazPjCB7TwmwY2PFz7fflYe16gBNGmouxG
VKLiSNLzMvoUlnucCuEqesNi4VgVB8XHmxu3RTbRj6Xj0m9Jf9Sgqr8HkIJK/Eks
gnNIr9XXqJMf6Ob0fEI/Cf5bwCOjAsvKtPQurMpX6qqV5B12rvvaXlNAs8RJid4J
1uuSq9orzBUENlSWHFq5pzbKN1ZbCSOD+dqIk2dFda3zidADjR+6IDTwvGGSd2wh
xeN3HMN8SSyxyI6U5wtoScQ3TSSQfWH2OXNpvMoY9mkNFudQdq6eL98TTTAjCyaa
nwitlnyVdFn4GHDIaOlsCTh8EJFCo3aT2F99cxFqSVmkljXy3xkxlbmsAqptzfRN
WXA03DasA8V8pYbNIPngHGULb8OXd0Aii9BI+QD9p2zqbhrKrBf66/4bJ70x+//7
nuWrKUN21pSUXuPQ9nApH1FvO9PvZG+4uJPPRokRpwd+dBpBWDpzZHiiLxuMax6I
SybBp/+Ab496+VUby9Umlv4BAAXMxOi237Y4P040q1tOyWyZlCtVwOIOIRhl3nFO
hSGhHvo3TaZiVr7ehraGYjwL8Sn+vGu3r8nZUAqS3LTQ64hg3acX9v6qpnu9zn39
SBmw1/wKRNJp1GOHO4ADPvmxe9nqHAf+lidz6AgaatP1zJX8BRo7Vj7qMfeR/rFK
QpUlylvzSphRaq9vCtV+VZkSTA2V0X4NGpGd7Z1DjdY8hT1yC62jhU2QT72hgSJR
nPcx70YRiWLyBQ2E8naJcJSjFNy5lB5GqkHGjau3TfuQxVdGZPwpVO5n5lpRc4Og
PxrN61eZQfcZHYML0fGuL+IhPEdqmgcmtwlYVA6Y89t8cRARl8atcVGcc0JFLuWu
J6pqeZrWryJtPJhzyAoYR9yDjIBF1p2jVcx4KrrC+Ba8Rv+Vx8EBquF2whDjSl2z
nt7HaUYbNGEmun1GeYNpFxAUca4lpG0tL0F7XrmUdlZBzdoSKQQJZmj8J4CGf6AQ
CH9mWdlOVQQtAHr+88xhleKTAgwo8voo6wlYQw7Ah3pENshGjGpnxNcJjWnaTm0W
MwxSqX/tNyaFDl5ofza3i6KZT/f3XzyDFp6u9Et/7r+qh2lZTNQ25mKO+3maQ1vg
gyaExsSDvYMdfkZBmSOx6Qn5jHpKSOengcmVXbkuBN33NRCrtxN/SzrtFZEpx0KQ
bYnUtkDBECKvZQqLjoSujUjvBHkTtl8EyIW+ODjhtVAHN/5mQjGnsdKdjnzegsJk
Tq/UbBDOiKDgIDYIPOtp7XZei7Jm/CIwCHE+VRbbLijOj1/KdB7fl59IGzRATtHw
vDaqYT7NdW1/uLP5xWeSzQ==
`pragma protect end_protected
