// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KjPDS9E6xlYQxN0WHQewU/HCy8tUzkNKFn7IMIEmbJc9iD87UEF7U030BzMdoegz
pj6GPNEfO5MrrC2VTrP7bEM+J17kKgxl0ff38EPO3aEAlSaeUwamKBo1igzJLudv
s9QTLjBzfPVCdVWfHOZ3GAP/FX7p1wDA1VggtuVRre4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24096)
aVcKS2o80PM0fzqnO23McGmEt66x9ebheir5qKQ1DCIMBGNjAOnKWPOYXr0yzyYl
x9SaqukLtqAvg/+0dpfOPHhDuEr59tszlYK/AMuj0KNW9v+5ITX0ZjvaENn67c9m
5SUpMI/9awyWIWbpD9xFkppu3yVz4lsfU249qbkKLA6WXl5B3oUdLEptqnHibvwt
db9D4XpoMYzEt3ajF/IoYpWQPemiKLuppBZ4O1DRLtD3ySV23b2Astrvd7zrQTK8
NFYCYiuB/9WVxUxyRJH+BFcsMtMjavSwEBGoGZ4Jnu2iKiBaubbrdEhiClyCvB+3
WkzlrR9RT7vq4tQ79cZz+eFOjWQF2BnGCBEnXmcHQWX++HoX/KIdTUHcmqDO3Wlm
M9rOzKbJV2wqDZc+7E8EJ6ufTrFtEyJHpxTC93B2vjMUiKMEQpaGjFYXhq2rBVz+
kpulL9MJQgPLj/oU52W8TCU3TYXthK9S3COFf2gvgAYeTnjv22GilYHwWx6Zrzz9
uRtNXOThZR/r6PJpsyWUdOvTkDIcElIxt5Q01LjNL0h7Jao6KSJ2KoZXVn7lVW45
kKVntAzamz8EBmMkaXB24C6TqaEalakKkxuGDklEhq/LZB2AId19dNrXZpAavMEC
vD8HSFpGeNe+TyIy7oIoagIazXJ36nDsJWINztZaixwc+MlWgvC6zVrqC5Zupouq
VDSMSAAv+fEfDV1VwhgARkNbkJ/SuskqWnj+iPsnjKnhtKgNs88B4oEij6MrGmcz
IlJ7rdmngAp3Rp+K62xSjxp2yJsNtuDRF9B5yhHpJ6jCgNT5QB5UXHHZJvOpzQ8u
v+Nnt803cKLvSaptVL491i3pZpDLMizzv4NKmE2nbBaku/JHFoKkl+HJXjeiP3LS
O+iy5UKC93SrGBDhjjnhlBJQcUX1+kJPpy2FT0EJ+7DXvviJ18HKIOn/b8FtGg2b
l7FLpQk0I1GGEHJt818eQcGJeOhkeA7HZedd1L4Ffv6/+Te3AMj9YemKDhp1Ii/I
aFngwoE6LJ1ONWQfPJxQeSNHvIHCrNqlq8miFVwQ3bKAwFwBq3e/5YnmmqCtujEV
tGRw7yGxOq8rIshB46iYgTchtHssMTwKTUj8JU079P0zx6x4fjPaqiENBvITUwAQ
ddqrdNXNkNX0Man9z9PcAvMUeyuZiIzKTijrFMEvs1O+2GcPOMK4X18DWfXR2XVi
PUY70ycAyBUxMeH2p0We+uvu7MR1zfkqHqhpE1KJio1h+F6cjvQJYncYMEO3P6iU
lkGM8mLNGGV8RyY7CcfJpjoa2E8Nabb+00zSJi0EPLVIlTwAVh9bnhfZNd9pge/C
7WzfoMK6uDVjzZ/rXAhDd/0tQDC0IjbrnPCNcek+a8zFBfgh7kloqBmkyX0FaALJ
CCJcBNWtlPuxq/BCAuZJpG93fUFuPbkwaBZeGdXlhfRKXWSB7g6nOAiIFcZydQ8k
Z01ud0TMWsA7wWvk6rxjRJtzNqQdUqKXL03gwkCJ1/MFdjNg6UU24jcm7Vnwg6xq
VvN0SLjKdOmopq0jzrx2XLg+Ass0wo+D+68qhFx3rYJ3hT/fv2+oXi19dAMJP7Mz
JHmFAOLL7mSkCkYTIaNO+JwLwdASVJsPYI/jpitoH44UsZA7I9PwnDEf7r0JBoVY
y43iabK+EimIsg28nf5IZZNN3xxu4V95XnPZS03l37rO/0MunEKoC7b7jiDChA6m
V3/8LHNXQC4ScTwEQ0HYFgP68C7OQxmK3hbkZV/UwNZWosYTHAq0ZgkgA7SCpN1M
6cHy2X5frWu97PvKsRTUC2RuLuFNYJD1NwUg5UIWogFfuZhzpLjgiZ2SK6g9uep1
ndigbuyOcBvReqCIr87uBnGZ6A5tWlESeFSXOQ0d0/XMVoUtlUnKOVgsRTqNkTIo
omtf01R36eBmTLvq3o78dmBQkVpr4JTBBS2dfjeYaipsZwB8rVFcVxYSiZIVID2J
OQQ2nAC7JbeQT4qWff1/Ae3ziI7lxo1Ss4wtRv+StqQBTHlUg8kVIlWoWaOSgUaB
Bo6QOKJ+uBh+02t61e28sy4o2QfkqygA4kuQGFVpuKOsDenEt63IJ1A/2u3hyVlX
qn66w3p2yR7vw8TjpeU7o8WGL/IsS9Olxz50PBwq4LSeBHdYz99AzMltksKtvamD
HPP5KsNtjF8HRpUZtNkfJnYnwhV1gL9bWm7K/I8ZQpKQQOMgwbx0nnngI5tJtQl6
gkOB8oDw1lYDfDBSvLv/1jXeWXnJTQFKzJfGiD0YWDOAgblcHAquQDpGv6pvA4d1
DAXBv+dWr5u1dQJUJYK5Ws42RsJpByLoiG38CfEP3xLDCw9ngVzLd8Ia9ycvz3Dw
+jQRlpGL5TNCCs7IViOl9HldvRlj3N5Q+CJe4ojlAvSxcOxva83CBRzBRREyWWzk
5TfeCRUW+zzNs5gG4WW7KrHYW2cn/p+Bq+dofUm0P+zoOvKVVDD+L3zxOiHWUAaM
hbgxhCwkortBjbvsWs5bw/d5X8YM9DqhpWW5dHgCaV+FNagvFcDPmtAMc2oEexpv
W6QiNCX7U4BBzubeqZQ6SX48hjcI1WSmpuVU1lakaqd9CI8Wl16K7XXr/Tc8N/LM
QtkOIRCrRU/TEMSZnGP+m2HYx8P5rGlXET8M9h8WiwOZ+w+M33IYZta3DizQmrac
z028f5e2yAS3KesK3bk7lVTCdVCQJjZHoENzB+jgViH0uDjYxiRrPM3eMqp1QF7y
zHnhu+t4cH7yDy8nEt7x3igpYMcJNAVm1sewW8LXcXvHbqZeKmaEMt8XxfXPcJyU
GmoKpLK9vxU9bo37eGr/KguuUfKtLMYNJ2PPXK7YFZYQgDU6yJsiTAjzwQWZiegq
+tG7YaNiSBCehjVL44MVPayknf062ePzWI51ixcggUOn//sHPhC6qqoA/uzAKEJP
5dyFwwqOAD+cu76QbcvVWGZBxFtjk90iCVkg5Ln4Vm9+M6BJMUkOU61ypNIJqHfA
ROyw7OEEtwq+wbDrPCsjxDnKJoPTsZbAfiGX7SVzD2klI6fZXbCRe9+3YLfiotDX
gBJVjGd/ZL4vENtKsvxcN0vD/3YYqT05bwoUrIuwrx3EruErk8Wm+YeTtnjOjste
e1r4uNkz80dEHWCI1ywuwNXRJ7lNGibogiplAom0EjhenJI8eKNttUSqgJqqGG43
uyZ45JRPtepfq9EO0Wh83N0pkwubPbwlrD4CqIjMxXbC0Ss8Mft7tv7/EGrDgmLB
ouhM/NVV0oklMKyoiZnbyEUJD4ITaVscg1ezO+EZJ0hPYvCMn1eJGFm+qH6wyb+K
uG7+eRBzsb3V+DJUnuvsNTr5HJFGY6ludsEI06g0qSUpmMhU1VR8H132qUSmZqO+
QDFNI8VyfdbUfamm5q6QXQKDVk8ysJhEx551lr8nT9uVtA5M9GhLCVpj09kYgk5k
jLkqzuYdJvV5rgx0NL7OK65YgzG0pcC0+xECt22MRaSJKXLE45njxyn+VU5tWufb
VGWXSiNs/QTLSZMXWD6/MLE4vtWV46uUwRw2Vk/2KAgycc/vasZbquDOz3kZZBw9
bY2hJa3mWdswkURhGnaR0mb1iqOhMTGkU+O7kvLIs3HHeo5z+2y09UcsJKXmztTL
4CifZL308wKOJGg1a9iwTQKW1p8OryPb70rj1feqdydEIRXA3wau3fUPcburDRXa
MUcuN5p+Psr4eZORviDuNjA4GHKvtgSsiekLsic4V2RbNLygNiQFEmRYEBCdG62H
xd08AFqlKtsrED+Bmt9bvK502SOhf9yE0qopb8SxlSirYY4SVG07IIuCV4agimZX
zNt9A+lSImlAGfwtppYjqVXKbgMi/iFCgnYzaLe+LPRiTgxy6MWT8G2e9iYjpEhN
9C6Yfb8QMdNIRNmwavbtQJ6uUOI3+e0HvIPINwUgwMTkhBFgsiNRPfgRnCEy+sAH
Udynz0/XUNWRB7obj7n001zS9ylavw8iYgvtLWzToC9cHNEuOzGiscTDLtYc1HLy
etphUbbcZNHDaJOKah9Js4PKRkIz1393q0Tmpg+BkilCGcSwdCyZu7udNnCzQXiC
D5iAJ/SnnSZmaYd/G+N0Z3fTm/B0nSacdsp29zFEPFfekdTG+ZiZKPaIKFL3NH3U
b0tl5BnEtQALFfEyQccdBZgLo7mcWmQMEWbX5baMs1JQAed1XozJwXEpwNwIa3uL
95gyLxxibj0EEIEpZLUjMcEDaeAkHbf6Vib5T6pbxQKkHW5hOM2gzc/27pZEaRwp
898P8C0JLTNil6IXucbP70pDXPbB6hZ1Qm25XDA6lWP+dP7PROlXuxUbpIakiOwG
5rrwdkq0bHBLiIdZJVagx9ZlNHs2hrpzFNMXfh9ym4cHUoXrTcAoRC/UALhbY4wI
rSydPLZzXrH9tnH/ZK9kY0ljVLqumZawWGQrBxrUPmGxrhHWycxLYVXFNVuJ8D92
Pb5pXducmrzO4gSh2tran3O2O3m1aymz8aI5LiQkIfV9A9nhp5W0fMcWGKILYEE8
spY1MlfDfLW0oDvLfjObVpH3gzpnQkDllcYc9xgnqot0Zg4D+Awh0bZRiFIzGjUs
W1MnnbPuQzHrDBMJ6rp+cv6dH4KAiIpTCeowlvhXheyE5qYOgVxDjYhabuOf3TTj
5P5qoI559XIZeY6xLWb41X8TwpDeKj1ORx2KrKdFkyeoMg1u5jDm12PhK2/RiWRB
QPrXPENlWvZvzY4jIf4px5N2IOkQesYIPx+9GDrsnVm0F2lPoiHSwN6RJM1P0TZi
SIY9v4PCEpxFuOCRQ0wsOP00yARPb9ir9KuMuNbHlIWHrwQSMoEmtdV6LOIH+f6O
1OVPrcEeS0MuK8eV85T2NIXmyyuhFuFfgJOXb5YUSR5R/xPrCDntzS+LH2hr9lR+
0xRri0/YOtGpDIUAG2GIt8ZyCrmQHcstt1UE8Fmb4Xd6903IJ2KMrHK+tWE7IaFh
plF11Dlfm+t81xEYGjQZ155eT0xLarPmhZpnSQxPoJAf4OOrt/5fI1oNQ8hHuKcj
1elAldd4OEy1OqDWjRCyzfUglrswUM5xLegTzZAtvZ/Ao6Wt/NU9Fg9bnUcVhuy/
d1I6jPApDWmM/W5SFGkk0rn3DRbBrtA09Dpz8hMKZhW8vgVfCXGnleyRN324kNbO
U+mw/x457kN95xcHwyjd7Gm5lKxsoSTKQYp1SYq0Uvs5oQHyxsuoZzeYoYs6Evtg
CQmkXAzCIU4k3LJGqy79QsjGF95HX21way9J2GpG31cjfJTMuRRplM1m7+ky3Ld/
wBR1cttPcL124SWXjVoLU0NQOpP4EUJNtQGtXclY30xd55xxc8UJQlaNIP2aivnd
qmn1xpeiAu/JH2/Kypu0L9HTWvHTIUldLCbSBr5KMwUltTDih8rfv80ftJ+3mqmo
6kx3KpT8vWhY4oDw6A95FlvF1EjoE+Jkzh+GhguWq3tbAOtJHa6OUmCUx4l1uYF7
8NlfYArQYBPnhmi7MqV+igZ4JLam0vz917Oc+8GF/wyeeoYDZ8Xu/FHDPjbH8qnv
l6c39sQHCTPjaP8cBJXOAa9uTtbc2UPPzhqpu7d1siBOvuv+zcF62DczgppQj3W4
F8XQWrjhrTEjgqYaSDsWzL2hRhdJ7MHtBSYiHfv++5MleKJZkmzxeyo1Lj0bsSep
U7HqNx0TybEeyqlhKCa4AeZwdPAMkMyJHfB2Z27k/El/ZLgcbds/U1SPg0bXVqd8
tLcFf2nuQo5VlSfG48C5FsVg00nW2rJC7k0OrnhujRlJOOC5swNi3K6PJbx1DsbE
J37xCfqPhTq9M0yexrDY60/F5EqzwhE2TS5es+BC8Wy0HIu7N9hntqBO/toP5Bw1
Ap+b9RgklkuGMrVrvBkxg6FevINs7I7v+9eL+XV8Ngi09r27rm+DXzADX5ywkxMA
wytB49vjRUoKlb07Q7/qYvKSMcUxZKADvkKKvn454hJTo+0zQ/HYbRsUXUfHDhzR
RXSwBMek3AibJk6tCILdWshL2d95UkP7haoSQdM8lEZDVM9TZvCPTTW8+zxr5nks
k/sQxaPjVvO/rUesWxKfPy7biKteXAVLWcOqgTBQ4YbCByDedyRMwauZHxHTz+4W
UopBzUj0JM9znPrKBAd1uOBbviD+shNuCWuUo+odLpPvYEmvD4tDpNA2FQof05zU
WNmbj10omW6v8KasS7rbqz14gGtMk7RVWqnrQ1lv9cqxkejJLrjTRNz28y7AaiGv
lO3LRbWBZKlcp1NKNtpaaiyPr0HwQQpJA+FEfSceCfO4ZiewCVPGQBV93mbMRedz
yhMGLmzAVQ9cP3q4tYybY8ukiUMW5/GSwo4QX+RZJbiizDYbecCmqWqG/pi3vpN2
tCr4S4MWy4QkiOd2JPPA96x9VJAkFkRme1gBwjHlJnEoutobnLMeluU7343mpW0j
s/Jnt2J6tOYc4cSBwZ2ENbOyKvdhCTQiLFZH9SEY7FtzpoSiTo5ICLw8A9Ypwwwb
EJOvdIoBkbgAzXTrtjrO62iZvGmcYaGRuYy2i4Wun6BnaZBBgJ7kNE9Igg2rTDht
r9tvNXTbJr361MAVWcLq2bPL9hDgMkltRkc7wIHRdf6s6Myo0ZMBHFTJ6ecWBLWL
Z708QgfNqqbFJAQJYF+ha64YjLGmPxjydnkutbRO18dFoyldpp4R+Ii3Vo8PaVUC
JMN3a2cUcyfOpEr+hy8rvENbb6fLw7QvWRjra7DH6ZLW6jLTCVvWvvpaq49set2E
7vuCnXvceOySVNmIkfhQ/ARQPz6/BpcMU/8b5k66Wvr9DbNR022XIrBz4Sme3BUY
HhianfW9b40zGD48I4IzRdcadTGgad3GpiYD/UuEf77ISZn5aHDugwzHxO/Y9+2g
Lu8jWYl7sScWRPyzDR4PE5meBM2/VMcR+yF6Pb7mFdGi31jzomvw5QHdyQeEOH6J
OLK/wtFeESA4urcrnoNLIX2FORzeRktw24+5E4/bI689ZzuC5LNwnVb2q51i4X/V
ANBd3SsENetJ69dtAX7tPGnr7LqpeFjOnoQB1Y7pMItA9nDx0QIAfh4n5ImhSjAx
MXOQsZH2pyO2501t7j8dn70rkuuxMI/M3PjDOMKQvJvLkzcsMeiTNhtCdy2AmjIZ
1tHC9zjjRHHbUxGYTpi49ox3qrOCkOQ8JEmzCyHWtOEeiX2BOUp+UxxI8PN9kRe3
/xdFohP+x8gsKrY2tK0frQENM98OeqzSRwcjw46mrHlltNi13DS9AuXB9OQ1fgmw
ZerNcNvkY3Xzm1PZLEwsP2z5wwMTRggd4ILgIVrgpPqo06FeqdDdKa8hRoE2W36O
xDUCXC0ute3XAeK8vpvkskGq5ghJv4RtKtnHFXpXMOI3/PJi5x2IBySj4JaOdfZs
YAzpTo5glWibz3ZQ8Jr8muQ1I9fm+ZOv9Eio7jEu1CcGU1LLEJ7F1E5dXZ9CktZF
XJZltp7XQmu7S+xUdOGr8LWnjRCroE+dUIOKyrbrKtMVOwijOciVmyrDOkNIN/WH
yWaZ3VywzaYTomjChVpWeqBR/ONOY1DcyNpP6O7zfFZ0dxyJ8vjWgcFEHCDDyuzN
691BWWl0P1SM/urTDvnqBMuTuD9eA+9ixB3mq3IiPKm6x7QUFGkpttONxzbhys7T
yNVDN7iTjVzQ5SQCdgT06L4en9/jmT0pMFq5ztYRPwk8GSQcUhgIeAdVb1qmFk+B
tNlrGVSRZkmOo9bx6Yqsrqhs3/CvAXi97dpSRpbD/s38XtKzhyQdxS9efOy2/n5C
tLiZ/dJtjo4iN1JTGECtLFSsDC1pRq6FbrePwyBXBVXcz0dPArldSXh2vVpFJQAV
L3zz5RpVr7G98RjVztPpxCvwMyubSrQm1tlHPbiYdyCO2S64QP+PEq2MJf8K8A6n
LHNJHYWtQnQxHO3RS7OemegHHOhJP4lqWLOFdtyrU1Rt4HuFuJBambfF2ZesWypt
0djk7VzDy6s213TiPg6xhYN2IrrcEnDJVZ7KeqFVJDnqAKVwPQSP6kVRSJvwo2+z
OXHfZu7znJSNUCTLdlEHSOaK+Uzv9T2sWbriAJ5WhOz/iyj93ml2FpfDaE8P7r+b
e355DYa36qpHAkYjI9suQ9i1yQsL6WgMXLNy6+46j3Fe3RfPlPk16k2DFhmVNNFx
732U6+s3vadoeMYXJvRNBgwnLtETHrYGvnxgc3AZkQfLtNeUTnX8DB/YQVdKBvVC
j9vJPI+A0Y0arTepWTDpR38Zq8iWi6RzK0hqfdG7QXeFu1KCbbFXCuHDRD+s6uY5
uvsohezty+iEMxrPXWxfUnQwTb2jAIZogoHRqfYD+IoPBTH0jZyCjOIkKQlnQw8b
7NWgG2a0Ydb1nGvGbaw2G2LUufnW2GXgtlmeAtfkw4hzHxaE5nONH/wMFabV8sD/
y0YMj9TN85/KrJf1n/7I8kokOXsMCROmlZo1ABQ92rvsfm4RK1miGaemedDEvsn/
PolwLpmTcrfTG9rlIJ0a5EGk4VHLqtF0ZsSC9/LjUpvMcPgZFNVcZ8/Ky4UgTvY6
x2U7A3JnD325cxeo+cUiasyoJbsAKxatrcM4qRPmC6K5MS5tjj4aRFKgMmCGn56U
LWOS7yTrCVO/MORW0I+vdzLwz1qiDVcKwZOruRvT19ymtzcj0HKPvS3oz85krP3I
IZ/RyKqW0WtyJ2xDI0Zb8T8KLx0KiadiTbbBCHe/UhBEDzfSgibLuEXs4JDZlUG2
VFeG73zJxLd8Cwg2Q95PB1akQzdt0rJ5PcG7V6Da3VmkZgBQnC0MyW5Li0pF5hKC
z1Qx1QWgG/wh8k18hTtIZ/78HPqqhIPw2YYauWmnkQwh1TR5xrkJWL+icWU1Dll4
5xsEw0Uubv+kyhfIPfdIL+LBb5JatVuALeln2RYjSy5rktuIPo2KPWRbhI3dT3Wx
PDFU2vP4WO2uKuMWUtRd5xgpL5Aw6u81X5BMt00oGwjd5Rjv52S1MyTSI+CzGKWW
5R2p2lk0k2duGmIhRsudNH6Lozsh0GZEF5M/kqBx9UoiGGDfaQ1Hpt+PZLmBIEmw
jXG9d32fJSUGByzDn2FaWHatFNyk+kT4AklJSsX7ofcm5QuTuGi8llR57L3ybhgy
NxBWbI9WZRkK8y2notaA9kkH67lw6e98KVkysjtezlzrl0GpcJbwFIh2iOC1BUjJ
gYD3YgOfPXBBYB+KxJPfcNH8I8RYB73BXeZPKYJ6SyR7fd2IWIVjOaaLX7g4TeL6
0UVwJis26z89uOAYEPX5CxQTRrRb9idA7Q+4XqotVLivUrukj5o9D6JP8KRSCLRp
wOxDh2aeHls1pSSD7m4zMV3B7wrVvLmDEA3LeDD5VeAwHeez4/6kj2MvVVd8z8AV
vUz/9hZW9Olo95qrWHEm1r1SjjOGjaQsvfnXGUwQQHDf+88mJwuw9WyH16blKt3h
tnxW7bxgkQaagk79RBWa85x8am0Mv8Euf7TphHe1vHHEz5ay1RaORo7v+qZYsYUT
3rHMNIG9YnkkUWqrEQpcDHwSXT8YQ7t6Uf6KOBr+GDk9zI5qT2zqjK3ItKCFn38r
kFG5SoraYCYAostrce0QEaDWLGH6qPrVdtbh/jeiJo3/v0Rl3R1YSY4UOk4Abin7
s6JWaeqct/Zamq3KLe0BY6iSnF9nEvxB087rwMKNDs8eQI37wvYPL3YLBDGUu4s7
Px6DYLFnHkslGoAyGEkRdfmeq3Y4Y3Ub/zGEbeguUbZWhSgNq6IDn2UgDzH9oirs
ODsT5/rg0RPSrLNty07nczlybXtl9jJXXKknL0KE7BgJkRj5aUyiZmdnrjbixmrB
qP3iJG5o26o3pdQuC5UMixeuj9wxbzhW0PmJPRSLSYZphrk70V1uNFl8rA/yto9s
U2ZWDJhzdrk/jwstD5QBiQG+N4Trj3GqMDjhs2s8EHBJcZpBjzn+TyB2MR8QMk+l
9I29DkaEfgaXrFweZgc++vYkHHkr4VoH3abWvvvBHN/TXW4Zy/taBVay2sVCe9EB
Sv+8TxYQOr0qj1pRbvk27b8RC29u/oFKOPyOvD0L3Hq/s5XwiSXVdRJWJms+OYqn
E291FR9GGyo8xGRRiouDDXcJ0OC3lqmlpFqB1EaRu97AIMedoTNbgradzuLeb+XM
n01PyzfmzFdu+E3arlztpmbWxidOe8u2j7Q7Q0uymgflBuWUWMOTk9RPyZGFFxv8
GJxkE4ipJF8d/2gxd+sGWQmWNr7c85VRT96aazDUwcNAVyjHvrgd24E6Ph4yoKev
TRwS5iXrG4I0rN653SCKZ6V9sbKpWbFi5AQ1gWUPnbZfxxpdJa/LOX7L8DuVfxDS
R4SvH6WTaWJomsufkzOGan4XwcAq7u24gU3Q6Ffa4fPrDQgiYfTYz0Q847U8ZKaH
RB6pLYRYfEsJSmuqsxgPFLeZX5Dj36HaOLx58UPuFQOyfr+SDEjyxI7yV0jRHb+v
sgJi4izRLX3lgSkWG7A2jxcyZbOICiFnV6qUQg77x7JRzyBAsbiNhUa8ct1jGatP
cGkG16ae10H+lbrXwOf2jO8/lilM+u2p4xsL8U9U1rvSoGHIEC3q3BlSgBqdXdFR
LiBeIcrefoGHF1p/KpaCg9GMzJZGb6NaUSF/+8o7AF842u4pj9vFXoz5eNBTb7GA
Dko3fZggrNgjhZJJL7bwsL/Ky8+DSnK0aO5GqQ8EmBzc+vIikzAZHOrbhb+D0N/Y
ceqg0ppYZslZCpwMNoZ7grtfwKAr7N2xwFvAvteRSOBKWIucgGMOQQZG9zlMLoZW
lM1vs76ZpzUD3Xl2yq2hXkrKketphyKGoeuNsrZBCQmMD25R8Lq4iCnKsr6mY3Yv
oYcUcPKcnru8UBrZPtLvyh4YNeRyHgT7eNzBcq3r+06D9P8HA8sDqKEV+lWNWX8m
VoWGg8afN+aWJzY8/gpXdH1tU6pFehvX4cC3DCPqdjsDXX+5V45yIN+POl31Nw4l
Ga27GroohAUUwZKHQamJ+lxS2rQe/4PiN50gMetrA63EGM0qhLsfZRW2v/WOdW4h
E916vNzn5ukyW7rMvOwEF6gplOKQh1DaWc0XacUFiigfBwzYZs6335plYcnaEuZQ
O54Ejc5hFfmQSj24ZyDdhJmxP2EiZIM57e9dN+oUoCmjbX1yH9cyEvly+wnYK77U
Afbq04gqjRjxC0rDusI2qn1YXQP1ggfeRruBnizQqIFQgYPOVldRS9YpNIQE0fVn
SyOnpN7aE/drPa20HNZWDNpTRDVBYLZUFQcxzvdwaYSH8J7uZzNDTNIkEdqRdu67
AkIz5Qgq0B32AXA4MORlPqQM9VZ0QJWQI/iujSv60q+3+yDg3PJFKG290VhiyHmu
bbUzddzOsRM9ZCUEBrLyxbPLAFztzg3RmhfeAlAUomods03MPuVFoJOdb1zGtrgL
eyyHzx5oDEvNQRMLUTSPVq8Gx8i70tjDFnV4MIV2YEfRdNj2a/qU/9vVwU0+Dzbq
ZPSL9YKaKJmjjQIvOw5jlYNOA9ByZWtVqkU2nnoMVuQM0hVhByeshW3fxFF148n9
Q3n0yepEd1YMwHIH+/+PW9sdjQqVmCI0BfvyhPP7U7F7RrBjRr4bp6f481Df8Haa
HUH+gvTP2WgrU1KEObIDwwtOtZub8L0Uz8+c/SrEMtt8+L7G6H2xdzLyxnKYieO2
dPccACszXcsBJAOPAvIuGxIRMuJGNjxCOPtfqZVkhVaB5hyZv2vLI99IUfiV0JbL
hxBjtXZmannZoiGZ7yIb32T+23Uf2X5T3gWSbq29CymqXXhlvuQ00RMpkmA/qw34
aLpbnsTXsqj4EhDdKk7IzgELngQD1ze85nDg2HnX6suJb2kERKH6YZZqOhWU0lbX
0KKjT5Pk8J6aqnpvhLDVYHUh4euhmRJN6NOZ3jgEUtlbwlT2URJBKLR0oyVjXf1K
eJf5bWQ25rp0tXTqHBMfQRFN+8BobAvFyJJNCKfiJc3O23aQIbxfxi1MDewMGz9a
CSG9ZGC84IYVrL2TJMoTZEFRtTYVY3lbeJgzMQwP+EEQar8iSphPM1jZYKXOFgFl
rtV9XStS6IDh+2jvuVoWJ6mTsu1bpq3VuFYci9pvrcZO8RMGhpo8rxL1q8fRRQrp
whz4ysFxCzZyQEd5d5vFii6ErSO6XYmOgZablqUH/VsvUON0ue/It928U5jV1OMe
HAi0WFt2oUD+9W63BaTviq4VCTpQn3wZEbY3Rnx5qtQ1uCQd+gwFuwKc8K5TVrdD
+2tEsDUO37BvtP29XjlLeupEuYMmXWyiRBVOmMx5YPLzYndJV3fGThfz/dcCgZVR
ZAfcD69n+pBILvAjJqxV1rzGZ7Tjx3aL/b9ySIWgj/nyXtIcyeUp5qtqkhWzzY6z
99IkxkWZQpg39ys2TISNkH7MwbqO0CCGsannRzXYSMB4zaYbr1EajD/rRvZsOE+c
Lkqwhggi7EiJp6q33D0KAJbSZW/lQVhzaYTUnDT1vjNWBsubVqiNsy+SXixpwRcM
DO6rF2H3bk6xV1WLjuqTS+Ww7ttrxa5AT2dAieUmKVjNysEyWp7r6zFPe9j2Hl1u
DJhDyqmdYmNeSBoF8TfO8LvyuPQKUM5lGSBfZpD6heioAa9K7S/T39wbJarIQjvN
+eGM/GRAXkk7JNLIGN2kd2h2BD7730HUPn5d5ifIqA2Vp49yzXMuR7fG3bkmCh5X
98Hlc0pkAP8iK7ViuefongbBBaZIU5oEQI73OduWrXVdANgXGmSbBBg0ktiyuGpy
xPCacBQu0PbbVVx4xL0I6U0jRa/aJq/CSu36HFZ0Mh7fGSeV0pkhUFXB3Ag0T5GG
xocqSmv8LS7tV4cjhIzdylj2xT+rOcdBcXgpNvJNxH6uwh+tEkhvy1aTtFhu0oR6
LIBKVa/g6/Hf8dEF3w1Bzcy6Fz196UTcZ77d4TNdw63GhhDe22giUBuUN1HqwMyG
Y/RzHIBcJP9zcgTyRmZZbwb46mHalCQAMDkiAx8ttJpigqE+OWfU+9IyRLYVoWqy
aFhjsudIy/mbwTmbvtopUz3F1NrMyA+hHggajUlXOuIrT+uxTuWo0bB6EkPj7kYs
a6R1jrtg+mV7k79FO4PV70PmoSlzBX3EQjlhn4ES04U4EI82onaEE18Kst6W5TVp
4ztxHQD47fCiUowoQy/4DnbGD8RFHcjXwvZXfnlP1F7N+uKSj8rusMXV6/ptLnwd
Dj1Qe/1fx3Ka1qI75Vwe1WX66efO6RTRRN7t/gmiVn2guL3UE/9F7VJTRoVAHXUJ
2ahcu+YKllmDoXc+IxRy9MJqqU9u5TJ7QO/JQb1adjTdMDCdiMlPPb9f+TL5mde0
EnhE9DG0k/2T/3DcYeHWmUYTqpP/aDR63JhVG2VrQ1Xq08JAuEwQV+03m/VFtmt3
1B+jV/HD28RzNrZWck7VTsRfNChrfNlQFBHBABA2yBaGHvxIBeTSgnsFQrUKoImw
C31R7AVkO1mYYkkNk1cyagVCgYiuFsIgeIKxU0157GGKlZDfAmfqVnSUh7tpEaHN
DeNOAVYBQt0Qpep7AJXmG/3euVql7s2UlGgXVPvi6kKfZUFjnePwQvGQyv3N8nqx
S5X/7lb9N32ofNcuYo+OUa/kwyU4q4mAWafUk5s+FFpK0L5wVYb07JjW1QMV8h7G
BP0FzFwlsqMwakWI9LWd3jRk9YetTTrknpBb4MKl/0LU2v9sNQwb2euNhXSrxsvf
g6xY8ucOUzNpzDEUNkVOOUepFRAWlNtGHJmQ52rp9lAlEbtYRjUc5B3WK2kn0YZI
FF0YfhE9YCUIB6UgpE7ySHZQurNJzTYO1OqFe0S+KS+rchIDvlunV59LBOrhh1AP
X40t0Um/02RSlgx1kb83AeaAq/TEMYRHyXehR7peu9LvDoHHsVlSvR82WfbofJyl
nsHSLqEERd/JjUk5Gl8OTrutsvyqntz/bUdUBocKCDy5SDLxl/2lEIi/dASGZv/L
Ub3psuGDpItmJU0kfIeHQZbXy7NoJ8JRhsbJCFslWiRHiInICrp9EgojKd+x62p5
sa8Gu9SefywTmFJIh0ImcGyJjQ5Zxz+0wPebp10pPqfc6uksr8yxJ3nP9sDQ1P34
Yy+Thywhv9gBnzeczXpvEhqckUpXh0P+hBp3Zew8X4plN5wS2eLj294JzgW9p4w1
yV/02EofIIBakccJRywG550nWZNvZmmgaANGl6TloOg6xNnZvv3UNui5oZXTcd2Y
X3pD8zzX9/XRpRg2DxDTUrdAXCfyCT3jKDreTe62YQVfTYyGtHXEP4dlrVhsEhPC
5NXwm6JOZYJrYeJa6CMm5o2pY3VSLg4stCLMxRZBDM7A3i9YPv9/VxKbyPM0eRgC
wigeD0TByLi/WiMQOa7RTOGuFY75y4/Z4ByPMwWJYpMEo5eNyk3dVmvzgmV0gMEj
rxUW6s++dCHUu9lFIr/gbSUx4pHiY5699M7DXZ+EDQ0/uZGKjzggLPYT4E5bbR5n
sFveZxE4b6xur2iI3UXH0pE1+moXeEPSFxGQdeSn3aVTxZ+3mPXkdjlFzaP0T0ay
kOUFjv/j+AjpbOeCYIPC+FgUZB+6wtaIfX+7D9PtaRtli0K7JhHF5w7Hv9+ElKL2
2evLaL/4F9OTlxef/fcvzE7zqJ9EDaEzR8dRU3hbIBKmrqi2eym6PlViiHtftiaI
W1zZi6zkocpXcecI6uORvGBn7NzJxJ592tJfq+fDKQBmFHGLpTr7gTtjhoFwZaar
DNJ4lvKCFdjD9KgENz78iv27OwL4F0Dr+zNKW0A1PiUD1qaUnP2WZTi2KodjZ/TX
2rn6gtMFQfYNEa7ZO1npvh4A9Aj8ZLqtbN/mTrsmG+uaMsZG5rcwI6Ot+4ERqNsQ
MOzQXlphArZGJ6Nc+KgCkLwh/Wm5cxafkKX5qHrw/Trkpc909ZrrNcNee8cbhKb/
pL1x71KyH9+Z6oWrVpL7NtnlLNNbCOM6sFBIMIGzuKz91aEOOJjDHzXa5ei5TWGs
Kd/BL87f2VJS2kBagj6QOKC8enE3XAMdNrCrX+Bfpj4a11TPmYfgiU5IsK78G1Jp
sJOy7w1+UO7hJgcmi6QCW9d1uQSgP7Uho5FU/aibv6Dgf9LyhthgzXapzAoa7NG/
8+40wNP2LM5JM7lL7FbALHpWzmG02SevfEtiBC1YaikKDE830GCw5Y4c1/m05+x2
oGBTQdDxaw68FuxWR+Zntxm+o8gYxB80fhXHjP+4PFKjA62+nnbH3S+G+gszIQdd
Pm0hIiMSAt0Cih2Ch3rp9SIh97WtX8jHjZz0dny7zfi9+WSOWT+QslxGdZCEMrep
m5uPEu4G7VstAJkZYeL93GLg+LNTLvA1xZ9tRULDfUAOwCO2oN508/jEp2Ycy+2e
qAK138aGghs70/OgwO4Cw/nBSutBRJpmCBebbTxO900Gm2ymvszqz/cCOqWuqYmZ
11S3S0tET6+382nd/TtUz2qu8qADkC2g6OOZPKvELlIep9HkN4PyuGKEHXUJUzch
QPq2WYGp804LOwaW3KGHvBYt6NOO1uGhavTjUkJJqWZjHWCd+0ezaigRPbSx6cRo
T7MlDm1Gem7SPeXZWZhdTWVl6e3MHLGd93FvS9BxZsN5cNeAUBCB7vOM58DquexZ
jpqKsx1Zq6wRcpOdt/CrU7yD+loNFXLg73+e91aFQISkjMQvaGa55zEUVJzHEBwy
mXY1ngb7DkQymfZqxFH/V+ppp/eu2SfuYgZPqokwVh2ncg0wdBMAFs99V+sL+96i
vMT+yL1nvcIC33YQRaRM86OGcQYx20WI8cfxDU0MzpGByryiKz1cZv7RhwG5sZGz
N2dLCxrdZTAjMOkQT5mzk+UGYfKqStKMSRmx4w3KqRKLjs67Njqkw+twutgK81Rx
D/Tu3JwQ/nuMMGDliK+/72i4wsDEwnbvYwa6p+fN0BEOXVm3mXb8XjzHS9xHtVUg
xY09I8OoM9l9pnzivQwbbCXcNbBi8GFyzOUp1l+bl5pUXL/mHcBJDotWkuyNLZtE
buwvOrq1MIiy0CRE4umwUouG9DRFEi7nmD3ybugxwSDTwQbyoCOKVrAh9ha5xoMp
SEgnmYJMRgzsCfOoNwasjsLrln0WmI5BZiCvVLraBDHGCRjuNGtkYd6v0RcaVde6
QxsUyaCPdN72GEZq88kH3OGTn/D1asg8746A+YKTSYuZD+LHm/HyfKaLIPJlt77F
WrR4yUoif9BSouvSh8efy7v0rnIc1Ww6g737xaTYJuhAbGvsWVm/8ibtMUWLfIKG
pukVJ6VQEMVKOSkDdyIHnKwi8en9IVWfUBkBW7MkuN+0vguCE7WBWrh9yolsavN9
E7uh18914wkmES07cCUZci2DGNbJQ34kCAAeI6et7C+Mgo+JbEJr6r3ncz5FhZc3
cWjmPyCFMD27Oz590vsFjGAQYFjhhr/QS78MI2H2zhWxGt4Iz9wsfY/tWiRWB/EF
163LnHh6loIotfW/G4LrrUXmXWraZctqK0skz4wxMOVpkMd6awaqhwsF77UaBLBD
1Rl9nplHZ2IvcZXlbviEVjW7XMd/M5BoBqKW8baisHPyd/eTc4uUFOwFwN61yoNy
2MWJQqChBhVgih4BGnzSNIVgsrFwbiWx3UQp8wVgN8kLvQfEHPDg25VtViSvyxSn
OZufTOCNKQ2i0/U7ZEWysA6d8wXx6eArw+w7wshVv3bs/yIYU3g9tn2lc8kAnagb
Ve/FSSOYWdnNZMSl/ftVJ7cFGjiRpuP6dNrha4skZEBzR3c/yvKBKOUkcQxWX8dY
fSsVldDdYT2lUjr365O4StI+wEPDnKAjpQ+Y64/W9e/aW87CWADC9kaO7JFoMt+C
rdBSsc60SsBKY05eQ8xaa+uW19KtPIvDuDgKb31u3Kf/fPZ9vCx+Y1m0bArRSX8N
OXPOucrW325drMC0bN09LPo0FTw+dQYfzzSyTFNQTtHhfi3AIk7Wq0SZsixoa/EX
ZfMuNxl4YvFnFNdVPHa55ocu1j/oLDtt5hRuVsAejBr7qtkUxuMtyZVxrV2VX7WQ
43qEN24qUPh/UWKkuF9wLqQBqnoZrgnmQdPkuK7S/LL4PHXih8GkeL7/h1tiMBW4
PAbrI2r92lxvuPuo0Bl2RjTiUECOUXeHXqTv2vqQPBOaPDsxo4LPUBqrezFdZwvu
LNgen3x0LREliSkUhJlZeEZtep1HQnlTf2aZe8udTpmO2oMyO4lALlQTzHfRGhDa
Y+XzB3h5xorlL22q4K06Idrqia15WpRRyvaxgRe/XmbGCQpztGybWDIf6EA0ZJKf
7MTKnfJh1crQcIA3/7OkEGmD11BAY+ucVvrfr+AXPzR5SaS4tUZAPJJ0M4j4qTyU
cH3hX9BL+jfTl7HJ+wzTtnYX+FrKwQ20hrt4yeq4ljHKFqFjUtjCrzqg1GzKYfwa
8wVzOZwdIi4XXrANcYu56wVCDZSzHb6Pt3Ofn8NfQ76ndOdhr6HiURj2BXLFh3ze
Qwdg44wxGl1A7RndFCyx9udfM2bEiOy1LOUX9HduwIErBb9Y2B0HAtLHPIHVEofO
OmMIauQstw5cIIoTD0q8H39WUIIUyK5an/sG9EiFWt98rmEJ9pn1wrKB7imXG4ZZ
Zsbi7Zzswpon5qw0LShfwZlgaIjWbrUPXOe2x3IJzjtJ8494T+YAbt1/sZObZV2N
GDO6e5pcN58UvNJEX59VVY3oC/sTbPpY/qUsavvHg/CioRTbcHYu33NDxf9k6xNK
kHaR7JztgHQpYMrCL/7wQ5t25C8eebeQxUGOXNN/PgTqThqDrxEZHQAv+r4YU1Uf
JTeh134idkRdyHfKdb/76ZMv34ozpPUAgsi+v7P0xzQu44Zwgvur1/75DW+AP8ac
b703r3gBgI9W8nLHZ5TdMuwNc2LcAZLLzChgo9lS9XOxF2D0zePuELwI472jzMnP
A+5bj6lVPUcGN6OxmoBVJLdisTJfbtrwJDEZCZiE8qzBpxFIM+QIT76N1EnPFt32
7Ra88nJ7CMaTOq4GRf38S2Eu18WDITQtFvdP44wANqWklSEATYOZ9ulYgr5OuhTA
MJkc6+aDPv+q5g/xxp0DmE4fDhGLzqEPKrwVAYPORdgNVZiDTYekHbEZSpgQUWAy
gJBDXige3UmdOoNkzS2PqG8dUcuYxAoJI/EvJpOL61fI4/Q3apBj7tn/NFfEiM4Y
1kfBD6S3VBqoIBhy2SZPEZCMX+yDJuYXjbe530zfbV2DIOFGGuhvXa0UK6fAMtW0
s1e97ahuQ8DsJdTF02GrTpPYaBBuI9XQO6C2s3rVQXauAq4wum3Y9qcI/itwlTbs
pXSJWCHA+RYhcgmceLS2LjuQ7pXk0ddB4trS0g3VlA23pEY6bZux1NNq8mFqj0r4
HIP/WTZ090pP1xpm3mMRhGgslxD2WYm0i9lsMycgHTPvTvqOelNxOE+DxwYJ82n7
kkXRTYFgEV010+Wov9K0GWkCeidTUrIlC5ZpG0aHiO0xRdDFUG5aX5zdt6FH4qDp
2xQNyRdpDSUqiCPZQFFWoffuq6693kcUvTsEblLwO8pLp94HzwvjuRWBTZ3tni7u
u0UScVLL/XtlsuQ8JMjjWUf0r3rRlmuEPQ5JISmJVD3FeMNnLzaNZdlCcCnfaef2
q1UgTIbvPwzbi76uGh+iQkpMY4T6jLTIUKGWBl3cOho1+HKmNlNWrsAyNyS+xRyq
WjPEgrfPn7TysQcQ/d4X0WBWDw9IbtDptg0F2R+aYjG04Qj2QqYMd9qHbfiFV1tH
CQrQdRDCnDFAR96v8qz49qbwXo5jkIDXxqky0CCaWuGXjkbPWitgvoDjF8OVWfmU
EPY7rx19HUTkrSGSsC5j6el62z68wc/wzxiGmq6Rt8YIXhlnQMrFYzPFL0M3dQXt
HolDDOB4OzNBwAIacWQg3AR7i40IFoHUaZJfElCnHKdTqMuunZlxr9Hp4WlWcApm
2wqpM6g2LbkhRuG8FsWLvCCbofypQm/32trE3hc7ppFHIZI6MQxESUHFj7IyEDTX
zfbQ8aDCs50Q3m71ZYhmfcaxQFTPxHl8UPXrEYs3uf+BKrKXjcfcTlLNK4L8xjYT
/0WRZnnkrHcv+vqO+GovbZSeJhvwJ7sMWiNHllowOEP/8NTUxKPZ6kbXJDh7QdFx
lDZPzUKCgbbAlSJxgVHZEnkXpMLkzi24CFNxMfFZykVeHOmpTXvNpJxCUfWHKv56
Gixn81jKOxGfxX4Jb3SMIswdsZOCJZvTk+wph0VvfavqpTPGCgIjfQv2mNAIga8g
rqXPrkF9dnBUZiYvXA26qfMeUhEBWdSNwbaa+N+oIyqbRwcIdKZ7ymoKWlv5xnPV
vOLEpbovJpjWlvBqQugXixn+p2IdDGsu1eba7rppENwzEcS6NPD0f1MFnyhXxfwY
Lb2JJJCM4FAbHdjmNTXAeamAZJDBJLmHv1PnNtQ42emzyPLFQaYrdY+49WvfREqP
ow8HWcAwHzwRFRGqMbvLes22ZGnn/lWCmpKZe1w3cgKQORe7kV9tUjsaxLnbKW53
61JsiHu/NeSbG4Otgz2I8wg8jTUivs5elHY2oEX2giBYPzVECrX1+l9b6fvkDUzK
f53ck20N5LmLAz8jfIMkHx79YKv5ypUjYoi52Pyq4JCLG2TRGI2Xx7SKuO1Q3W2Z
s8EshSLV2bvzw1POir0lzxl21K0731J9SYUWTZ/8suEDmzQ5z72WosUsQfstQZy0
8TpPQbIJQgXVdiO6XuWSquz7BeZJimlB/6s1OsIH1wkr+5wHPHc/AZX3g2V49uMU
AAnuS02P406lG97TrCL6p3laPoFNJEmRyIQbe/Z2wgYbGhJm9WI0uNDlIgcBAzsG
YMg6aS+ZQJko5AtzzL+kysmZU039dqQxsCRdySZ3p9hUEkaQKMlTKSOABvL8SFMM
6IBvqnxKKEw/1wfKx50xbX2fMb7O25IcuaetsgfLpFqaxIL8yD5gl7hDRj8JqwMS
on5EOpijzuRWjL1f8wh7YakYN6BYQI4SApJQDe3FVb7AlWWYouREoBGqRUrAIPn4
ZVP/vkcuMFuWe9YZyGYMezB+wI7trTwxJ4jSMEG0kyDOdl6v8ggtiNWOukz4TPiK
3sXw7dDGuQPFf3R+rt78mTsk+InWxtVdCvNgi7xJ2KcGq939VPyRzluuuoNTdFSq
8edwa0KK+HKESruixf+FKkHkFlHF6d7ws+/OPJG60SWuIpJopOciHcGFFsHuOqub
7S1at3Bymc92JYZCc0mTGRE96wI8ATNaeIB93tDoFg3S3RLa1Zlly6LI3yXy+un2
/WA7/3TdzN7lcSSWw2Y/kBpYenkAVcjjj0XO0ubXndbuYbytMlEjOS8HP1klrDsp
A3LwQozq4p6fa3RgIo6zy98Ih/s7PNWuagEVB+YEp5dMC2Rn8+iZ3gYW7KcZmyX6
Ik9oFoYb10bPAznkCznf60jis82LpAayR9Degn1g96HRoFYY3ZO7ND+Ou0R6usf4
eQyS9EyzSK2qornPpXLf760/P2bAEMs1feW85KTFx69aEwlw6sJz7x5utnL86/6x
ARVywbqtdgiVuDPkcyMMxjw5VO5HPIGKygCqOVq6B87pyPYshFWaU99Q0V1b9feA
A3ExHIatCyy2c63XkuZzZvnabVxsNu+lPjW4Idz3J3bU+4N0ou8IG822Wl84poSN
wEXg2kCoSbrZPgufWMKpf0fammDC/lpTo7qjEyff45qUSp3nkz5O0UrKLsx37ux4
lKr9qCoNEulCceSShqU45Nb83XoxToCmdvSCgUWZT4RT5T65mMPM7MhdPLqW7fZX
LKTQlOd8fL3GbSjpDHgpuurjX8dCEbE2Q7janAAU0MFjoj9wQbYjLdaqkxPV/sVr
bfCKPEM2OQfmo4vOJ4S/emf++B8Zhp4VN0sBq6oaAnC76ncaUqKqCFirAb4wUFFB
QNXwLF3yoUl/DSP9WGfTnuAYNVdZ8pQMHd+FzgGMH4mtlfsXG9vwpabpiOPkudiq
32F3nxOHm7NnXcrQQy1/1rQxfYs6unH7kLmVQuBe/YcPgpVqx6bVHx77+BoGmdLQ
tVt7DGewkZCrIUtPriRw1h3i1c+5lacpjeay6lngwpUZqPQJ/nCnq+mRqjaGPs4e
rgehs6dMEbn66Q1/qSdnny59oWvGYW9ZNRY3pDemey9X4FDnhjmpByRUOZ/7MyVU
OjnQQYo5R54h3wuiv5+S37K+AWr32Fy4Gx1eaLiNXtxLGykJ/zFnmTPw9DLcymiD
e0I8Tk3JXdZlXYxQ+ZfOaBnSHTiPUgmeLdWpZIFoaARZwk/dC9Z2HtxcFA5dl+rx
pxjwiyIjIj/koTATyTyWd/Trm1ej79BUenDnKUQKNpa90GbU5sY3Sd/NV2mX6XPa
2loBNujMIqYUCQZQq/034r5RAc8KpsV3vQL3bu/aoMx+7qhDAT3+4GC4+zUDR2Q+
heUeUUj4JGHVV1BRbLI3HbwyV8lGWXpmlakXfI6qQDuDhviV0L6Es6kER7KirCwP
PQ5njsdOUCDQcEu5F5Xg+00aPIjje8Rzc/JPe/TniY3HrDGPks9MwDGgSB10TQgx
dq0ny1p0U1Tzinqha4LGH+f+3FpZNjiFG8xrYMhC1g2htpjxvvfFt4bU6bqJYmHi
aUGb5gFXZlispV0F99OQIHlsOndcQX7QTS1ONGLza4nqx4dSI/AR2T3IClAxa6rs
MoZvwfXYxb2X3A2DXDoieeV0jWMmR6K9rUTx3q8yqzl4K27WWzLjKRxmhQDhfbVg
x4f6cWsdl8gk2SDixV0ykQ/PbZiEfrCjL2KlnQR+XNhQMd9vIGJGXCzwr93w33Xs
M0C8kBH+ndz275OeW/Iu7PkHKw8Y9r5wVxkPOhbkaUWsH2J9hPDsk2HTqZ5UYJNu
azxwh6G3KlRXOY5DKPtUwVAVU2C66Diim6KBszzsYrFkcLtR0OnChKjUOOzn24SW
EY2XwtwoWcXeXyUIrH60exJ6Z3m4BA/jDU/KKHlVlFo7e0F1wxBw0+sb5PFHcjAu
/jeIuhoB/9nzrGnFQ+TpdCGhVcPAcnSKCosMPF5OsfQr42vzXQ5JiTI/xoc+mm4z
+ogoG4uQijl1bWVHR9nljYV7gtgMUA2HYeBw3aWS7X4cMiRlmeolkUPVgLPP2ePk
PKimt2It2jZbWecW2b4868jXEzhrrr7zqcgakhWNswIPRBLFpKoiWZRp09OuoZzu
68CBW/ZADvHcgptK8Vxod6hvyweroPhA4bLjJnc0LO+8SXfOu1gtFyt2mTrxxkHw
RSkYhv+RNHB+iB/zFe8uuoroGZJ6CYrb9xzfIUFMBRH/wFPrWwGq1zkVl5r2WxPu
gr3SkYn5bPn/aRxw/m4fsJQAmJ4Yg8LzYDfh2znucd+w7YpGnx1V5gq2LpvMrfmG
jr6HcALFh9xWPEk6318BBANDbiwICoRLJyXKLC1Mjt8lWuYrniDifRjcIKHfv4JC
Z8YtfrYr8YBSWHPI6XYCRWhFWZWloxQfDO2hOC1Apc80pDpqLFkESAunachfULNY
rS5IQoV9+p9cLefL49tk24o8qyO6ZOIaqO6PyYu0difXZ8lTNx7QXZ6q8pxLS/zb
fWfPzvsj7j1LmWtXK342mYDyC+1c4OUpbU//o0QsI6U0nTmS26SqcDqh/DM6cQVy
KUI7U00T7myEfQAchIcV0jW042sddEWFaL7nqMvkg9SbvXQRhy5MHawSvSuFMHg6
qr2E6Qd9MNO9nPONlHeVJ7t15FdKHB0PhCmYylKtStdGI6k6B6pgx0VxLTAstqLw
p1KyxP1/Q3qThezWAnSFkwVQG1l16WmSOMEu49MHLY99e89aJT78gkRKQNF6l2C3
dLwrD38DS7wiSZEqoQSnypWsK4NNcFsA5CJgPQrp1nzFchdpkBUnTFT85AwdWGAy
9r9V6t1DmZOQdEWdeBpkahI8K+VHr5FsbmEZItxPO58Q7UDEPOYwQumffhV2XLnx
WtKuyTZ6ZsvxeblniMp41Y2FDA0+8ejfb+mZDI6CPni3L245qnVDKr9G3LDdIFWv
DDVSt3FzTYwvNUK075a2NLOdEXJMySaTfQMFGTxHUTXXKsE5PeSFP32xmqAvUB+T
OyjrDc3RfNwUm04l/wTkipifysfeI1o5LWQczX4DPvMDA1mUbltklFuGLO7HNSIs
Y+ThyN1AiwZtpp6FP1MbhIt3jzXNaRI0BCFKcPgsVJLWW4zP8ZpsQ2xcwgwSYkSC
6Ys2QwZJdd3efhvf7MCGFndPCDJf5q/OTR6FJIsI3wFGS+aTP0Vj/dB3oTDWmFtR
cATFX15gV9KUX77esilu8UM/hnZNcFdaCUnDDfRwlkk//BIq1yXH1/2ew+y86Gfg
kx8k0GLhucWGWMxtUobOq2iMtpyAinhqV7ykOhRq9W9NcWPFfuLL1gwcMqibDhvN
CG8zlCHv/IX3trtt/ZLwxEbleUi4Y84/236klsBuJUCxKd+P5cds8U3WIQLbxecV
Jo2YYslWEg+3ugW8UT7HVOqOPYlrkVlsKidldC1SajR4dJf0k6kuO/wGbiJYpGfA
cfnKPAbbPcWlBoTkjLZ1UjHJRE2QHcQ+v1cGnMNb0K8YlUHh09YQzG+SendODrY6
UsqySkSOjtTAaQbykGhKu8ZTnYTG6LHOhCiqdkELTm7l0m2V2M/7yJmwRauVhG0C
2ZV4868Ci6Ec4DSGrs9xcgUhEOF3LDjQmuX7SHV4H5Ug3SJx+CBzjKDkTmr++Wmr
wa+S3cPVmmC9n9JMAvAEgAbnelCo+Tou7frfHnZvj4pbr5GzuVafaq5m7y/wm/hT
rpcxDa3KigmaglBHYUzdGDzVBM7O4/zys3tFWnp/4ES3rasYNJF+AbKHCJAp5VAj
0/YQF/vmxJa0m3CdXC4yiHlgzTYVwXHtDgP1WMKLtVCxnqkBJbQmtRNOfJ4h9y+2
lWQbN2Ol1vA0XeduMoGZE3F4ubP6hprBXdAQfLHbO/DiGXIfHj2GwIU1dHKdPvuU
g8LVQNgB24niLGzLkIA8zUnqSObxBfVlXs9TDxjWofWBo1NuGWfo5zPEOGaM/ggl
BQyXjXR7wmoaDDF2sA6wUeX+A82G+9mTKtn8XpRUBlSAXEr8RIzMSAIa3m2bimWE
RbFnTzzgkXPJzgrixPGUsYdrrg0URMTcg9JGRbPpSA3n6focj31o6l6ZFv23QQwh
EG4mjP4lF9bMxDRkDJSRp7GLSkMi0FA50mKZeFtlQWIM0+jPPmBp02cXjOVDd2dg
6XKNjhGDyDovODwYle6hv+Gjl2cQ9ajJp6o/cE4JKDxtTKq/e+lwCrS6LbXZQAOq
Sx5T+/M9VNhd2YCQI8B7iNwTjQHawGs0sAi6YXWBhN1oOQBEzddJS3Tx4GuBs1zS
g8ldLLYCXTbpul52LSO80jXQLV/IxG5kQQgDBXtndeOVY7atvr80yn4ksRGmceAp
zrI8VotS1nuBA9HbgBR7IYrP4CM95Tog9jsNVy8eIbQmnbkgB3/sXte9pPDq3sjG
jhnuCuQAr+xBDgEo8ag3mk8TFM1MQ0sjfgDfW9gi9lVdLDlYwfxb/FcOdHw/SiIA
KTW5PzqMjFVoLtSLi0BE4hiDD8XELCpqqrhwj57kLxhB/6aMDugcDLoX6bckMhZe
4wZz18lsahZ+CC4RBYlej+in2dchpEdHaRJXSmEFlQnCgRVTHmrSXrqlJV+LZEj5
E633BUD0eSaoGc7gHOdh3AauxcsfYSSolQ5jKfwtF2k2Za0HGRXezwtjjvCuwWiA
DcWoOty5JUdhd3TQ41mYK6oFhZ2mw3GCbbb0sRwsu33k1am+H/3QWGkK3jB/eb+p
ETHvVGxfiRxVk1dvJR6WU+11QPCl/Ux1y9XxtC3l8XkH3zewhIb6xkMOYLxR/3ML
/h79Bddyn1RKYcf6+iIHlqbe+FgAZsMBb2UywBPs4G7X25af555eR2t0WPDbii2O
91quoUalZgOdCEsUzfdljwwWBpL9Gfio4w94Ae5LEsDLzFtquHoLcHn/TX3SN77m
8f66L9DeJ1nbW431Rj0g2rR8nu+suE0m8j+7QhcttDOmshJPBt1eeCSnexMRxzSZ
RmkOdEjjc9Zx7YEXPHJHoLxaUfOMzGo/CwRzIgNYpGPzcMQZAsFnfFTipkbIxWaT
5f+ZE3t3EgxQJoN6+4XKFKGGt38BIIomIku5siFGMf0ry9mWftL5GHxGqo0TBsiv
oInfjg1566MOf8xbzC2Ga2xXr3oLFOoM8zNWKZ61srWVWY7snXsWVvQw+ekwOKll
xmVX+cdXjvTtIWCNOArmLdYq9uoVVBTNz6e5aEB0pkBnKovnWpuCvurQER/mCSgq
mlw2Xjxwv7WsKrfmfEz8HDkdGXYVWvFIwHm4UWx4yuX1jfDakd+vGBp6Vn/XoDjS
4G0OvmxT2PxGL3hwzTp19sMOihNZoh5TqZrp2G3Q0s6/mKBCmedDlJ+yIgDWOC6h
BUfmMoUBhYm+isVUZ59gw6siDNUdY0aE7c2SzxX5b9kmQQHlRxC8IJlo8tzMYLoq
6Ngd4dnb6ER2wA0N5+JhgLMtGRilBbwJPtxdxP06r+P3Rc3XbWGTL+HjYoaHzfco
fgO7xkDrWN3GCURQpl1rNG6zaS0lTqnDG5fqkKfhsi0F3mcUMB9MIcTI8Ba+myXZ
5B/Ohdi51LUBS49fHQFSJVWGE5D3xdhO+Q0KD6EgRDO1aCkNPDiDzubsxfFDUQDd
EdlzJ4eneziktY1QlFvkvPhhMrr//sTggtDNYz1qzJ+tSXWkSNvHnLWWarFnqORo
FXOyKkCuCwxvVeC6VIr15Prw9VGnQQh+VsLVj0TDiOyDDM5uW3BrHy6tp/gPtkjG
K8D9veDlXc9PTrqUexe5Nn501snAjmW1LDPtiIqFkZYsMXK6yc1WJcRJu7QfI7Tg
3eus9iCphKZp7K/My4xq3DuhiXUKXwkRdZTOn1nar2LPkAcb7ekRuGefEtfYSObG
z7gZvrsSeV+E7rmmoxPwlY+UhhM6+D19xr+QEhuGVspT6ViKZKcAdaJFqyqZhtQ9
CnHKMdjx6M8inU38QGKKVGZFDHwFgGTuV8RUfDTeFnTZLtfHd7ugNIcG9mmBpwub
mBc8ielzm2896AR3E75sHXnPwf6To6Zr3ba1q5JQB5mGmd8ehoeUHzhQnQ8CJWQq
NA4UrN60ntZD8GNIqQ5614ycb3z7YgzgcimTyl4piNK0Zd3XuNfx0bv34MyhFk93
zynkCxUYvAkUK4BcQQDqyZTTMpSWCJusySPH8AI8XzE3FSTdkzv8c+hK7cCEjhlb
ueoAa2yLFM+saOX2T5A9qKOI9kdkooh1nS0pn4zn414QIxjheGWkIotxFqw65U9Z
msBIjH89b61+o/wLWJL0PI0n+lA2/j9zQaKUN8IlWGc76c1Bigs9rdb/YYP0aFUU
GaDIpfDYVUh8uAe3FU5J9feQKX9HgLQKu89oEmhRp9WB9XnIG0m6APA9I43eSwhv
naIpzvgSZRdrDA0xOqWTJjyfAVgrKcUTUytDRkCithkm6O4KZz1g31u0MwhJLlw/
6RzIKp49y86MEasqhDnSQt+fpobqSyNxBi8AhiN6kyD6dsm/W7RiyzTtUryePN2v
53ZCDoVVpj0YoipyYK1exeotfKNtE6xg9TvfRLBx4reb1n8SbCdw5ThGGDeY3Sa6
nWyAaAlx5oZlXXTm0cQf6uYyM9Jnuk/b3ZObABtigMGlOoYOIlMI+Ar2myeRJR9t
Qhq90l3OpXMu1VeWLGsa/tewuvRu0NO4EliuOGw/r5mQWlr2qxYlQkxnjCftDuwM
f+xS/d2I//pkEuKSAHFHpoor/yS8G8HVr8WCKNkygqKa/AwatmCWVYMlTMhVN58d
ewDT6VsxD2dtBSoD7divDXSLRn6/Ngyti4a3yDVVy0wRu8L5fobRrS3ypOnkynh+
TQkMZm7ibGEk4Q6C11+4gsYv8HVNKI1W9SV6ihn5BNuGzXuomuwr4aqUX/5gc5wP
RV81DoarjrZL8pIlUNvxTIRRmVhMt2UbQ+qVbtv3xCSoBJQAF6S9jX9KoxfjJrll
gPI6M6CpXI7XKq+67W9FVCX/swsUgRzFgaT1cfdOvpUv5WgdAf+v9w99xCx4y/O8
fPyAz4hr5KVE2uKlNqLiTojGYpWpfirbDVfjNu03AYZXTJ2+/s/8l/8G5Og+iiEa
42fy1OlYY8NoafT0I9tbmYp8TaBk9E/X/1hqmlxFL1BAyIfgMGNigGWs0Xy5gNf8
GoPoIaOiSTHzhVIyBBsXyJZqp0Gm4LFqfTY1qaHOQ5iIpcj13it8SVOwTnkHovVI
qWmxwMxWOHNUg70ZW497e791SgWLvxvoHwx/ZRLQgaOT566Cf6B7vKd5YWWP5CRz
Xlc1/2E7W3W4RraOGzks1ZA0bMmBprmI7JbRx1u1m8Yfl1ccuykQ3WUGEjS7Dnn3
eD/dlHcLfwxVIeqDHiduGEdiYpTkU7SlSWFzNKIlzbNLUutXV7oHAGJ82XspHh3x
TDKGbusa/PIOq30WfumXyK84iLEghm++g3w7yo4OYKlPWnwQYv9xHJAK3yhll7vY
8DW9ieKESDlZoQfPSWf8PdSq+9bTg9vgCN7VlFEI03ZCFBqoIpBfH9iGLRPPsn1y
bZVoC9c/OKFDTA2BnmRoLK9OU6mmanL1ZoFWX2CxRNTWz0AhkckXBy9aG4AybrPZ
hhKLfPz3jzPJS4QRpJ780YQaBOnNXvzzH/52MjkALmXB/hJAhHypOQFjDH76quNl
OwMvGWITNpvNObpIRBIJu7QA/ae2theatzvYF5yXNHZy6BGQsP1Ikf3IxSe/JBDz
ZrtXpiEBo9OchxdvNimkhEjcYdJvexyxlPfsdIsRkh56bkzDvBYe6Wsb41dwjtcN
bIDDh342yKkxP5Qax0tpdXCLQVG9Mbv990V9niT7Cz+G+Bbtw2wjvVBqqTsmMh96
99Scw2uMjOCOVPsB1R7OHskre/1lH93pgSIbFbJV0KRe6gfha5MNnk1neFwrlAbv
GK4t945er34qcOjg0itCkV8l16aQc50DYz7l9LPkFKXtXldhySsXbgdY/C7ConIq
iOJ9+4nkHN4IGtqUQVWIv9VJSCeNBlYGcJRkTSNpNdAfBym0AnskFbFS2BD7i6WC
XjzFBK3nXD5ebJWbhN0Aw76JOYr2c3sKbXPN8nGic5efoa/2Gy7QX5H1SbRVUXOS
7ZsdwNGccMex2kwllnBKbN1QSEb0rJhnRCq0go+22WpF0K2NtlDQxK6FrACJbs2d
/POnbmJKKbPfBqvLd2HBeorLeMvrx0q5mVmi6fHJwzms2UOdX0Jpe5yNsutmrYfX
a7uI2W9S3pXx6yqVQcDd0ekCNcWqctSo79QK6vYlcHoi0SNKBQlafYpLbfNVGR0d
uosrqOMebdqbgoxnRWtIgMh9RxUjWDLOEkv/rriMTBlpoyDQZ7wKrj6kZZVwIUsZ
WCOY4NVJRPUE0lcAKGBAJMr/67YliZ17z/eylVAUrbMUo+iF0Tp226KArO39G7TX
XTiNbbk48ypmUnyOgCqi+7qApu/N4mO2gByNiq5sls6tirjbvKKHrz0wEphJCGqp
zKOJoM7mziUh1YxkiXrQ9sTWNZnUrcKmqvvS0rQcFmBfJpWK8AbYqFNQ3/N5DNda
afHdfjPNFgPLscaCCgMt9VAlNsh7855e4gh2HJBn+9fHAeayE/7oJBGcPXG039gr
LDagw8mSfi0r5LYEpiImBj9EeMCEacsU8japU9yqvdns9LDF9sGlTNtIG2CgXF+i
z19nP11Pmpv8yh0tSG+xGdsZ9ryu2qFVnx84Q5UOymakuYmct7srLPiiQtqmbXJN
WNf+lV1Oz/bb1VdLoeBVVpt1jyYZHp25LeC1OgQrjeae1W/wNcAUDW7LIOb8kJl1
6sPnABp2DbOb0ZxQK6JpHVGPsCPODiSO3l9Y+f9tISQyely+Kh+CqVRksSVjHWY/
cgEBN/cJGeiKhJhm35dRF9J2tWuYqckCEgeb1J/aeOCBN/Ij9EkkCpZ8rtCSMnil
M+axqwYhdBddug3XWHXKF4rHX30yP/FbI8hc2RAGc5Vh/h+zBe4SMRNisPRBn3yE
Lol/unv0ZzW/eDxvqh6Q1VdFbVbQhJS3vmKqwvShBczwGKLlTA8yvtZQixndVCj4
9mlwdoZPu00aJughqFQ6u+/Gfsbq3VccS/mGDHcJkmn+KSSkp7A1B+6PRduccOPY
aYOhKdZwGb0Nf+KMts/AiGFZt2TLGFcJTWMop8Bkp3E6yFYKhcwyKuVnsjfLKmvn
OAGq/DOH5DxAFFMbgLKwucTqfFjNjHzvw/YOaYMnt51k32+E/z8OfiBMaWU5uRN0
2ST6/dPEWvNQP0HD/8bwTiSWNYZCqSro7qbnX5JHnAWTaRsD9PFvhcyyDboh98o8
7mIeaqI6Amw5NLCmYBD/ODrq8K6xYFyQp/dJKwPQsPWIJ09jHL9t4BL2RHmpfCJh
p2CrEbdaW+hk5+mHHss1a9BgS972hCo0Tmaz0iRplITrjQc5BhgkrPLlLJx3LnF/
UEky56Fk3PnzroTFk9a4ufbtH1qC1wRDhce7jM+ruvFIWh59wAp7O7hRzyqR1tiE
bKADVuzwrSRuokpCRoMIsId4EWuXcWTOTfNtCzbH8kjrW7hzPjTHEJuWen/lemVN
YlCx3YNotICJWyEkJzRQSuMsdCQM9IOflM02+tv66rq5K/MmqMqZUOveuJzAs5Lr
1VVx2DL4Q0vg/knUz2koZewFNZwfa9hvOeTE49XepjcwcSlU64KS8DMdZ69aPSOQ
/ArprYsv8IjxfZds9CCEClFyvVbrYH8b5TROXgL5bqNAZxF1rlWj81SPe+6eWe54
Hy8W3wuLBlFWiLYsNa7nuf5qXyhZZMlSL90D3cgRmiZfl48oSrH4mQm8P1oY/Tak
lSsHFQKfqPVz7PZZ+6x6WT0dZ0R+RElRUp6miH3z77wye3lmuHVUGiwk6fP4Zs+y
LXzXexYsG6mdOHPX6S/J7b5WW9RR88GKHR7TJLnq7QkKl6aYFeDKkQo8762NVPbB
fdoVomGgMA65s0qyiqtRaE5hyQe7eW01lRQxfOa9ckT44F0mrthIBBBpvqvCJkIW
OtB4713YNRLpgB8zAqN4MkpxZGmYLGsAQsj9DhAMiMWRU2YUbG68s1YFwgs5KwWq
6yevEtBSftbV0LuXhXpddtZZboV6PjXRT8XV9GwLEYPv3bCA6V9hyFyFlxnxCgcL
cQL9NO4xgLCsetXN9vUQvczx+hV6mnDGt0MUrsTmCr7XWYuCs6mYWfaLk2Rf1/VF
KSXiFsK60jS7u5AYfOKA+YYDA2aXpbqiqTvMv0ASxUFfLOa21HrQ0hqRqbFBb46d
aL7IHIQ4I2FF2WAOuADP5HnlMhF4qpn2rcwdMrcrxhwUYev93uw8bG3GeDFjODeC
WfzSMfuoMLPRR0G477uVBTrK8w6oocbCckPSppEPYaqbxI8jylMI+u0UZi9sEPrp
+20OWzO/4fJ1ClPcj41+VC+vywlqTeZ+B4aOSiOAzSb02DsiYBBN3aiv1ZRPErdj
UiaKKCMHyzY8pxCgcszNr7i5AMlrHVVpdylU9NaJtR9+PMo6rTJCAG45UwsVDsj/
JP5TXXPP1Kda+mh4+eqdoP+XQdGQ85dNggMxIqYgycIMS/VY+3UcWC5H+STFV7Ie
3I/Qyh/gZQKoB4NJOag23rgMELjQZ+hiyqRFHY1ZyrOb8xJUcq/0Zq9AhkZSug90
EcQ5Qa8xi/AVfkRmUM5BE5RHnfPGy1RKBdL6jL443Z0/hu3jJhCp7SD2b3VO5WwN
miyuOvBe2W080y9sNwPciHzOoMQRa9WuU5K0Ps2TCl32cCCuAxZ8PPJV4wgzKBya
nquaunkeUN6jTW0u27CChvE6wFEZo455k8OK0MPWwSOGFnujyIrx89z3hY7S1vzY
DddywAo5RDW9KcBgV0DJqyjo76NSgw1viQX2l4y7T9KEsQwuWEnA35zDNweobiU/
Frbr3z+D0BF/hpRYUD1P0QasDXoa/ZfGEja2z5McMonrpKR2ZoKPK0I22V/Fe9Un
0ISXccPfOK4/oudfef+NCPSjouOaEYxN3Pl7doTMMcVtIzYeRM5gCo4iv9v0VNC8
NyL7PV1Fx5D7gGuFJleV9eDfkedcUy9CKAP+BmmOmsTwartKVPNhFgtzQZ+5E0TU
22mLRM6vTZbT1bBQdzKq08a1nXspNGuEtLPt72u50Mdl6dBFvsL3EPvfMGHzrZGI
GhJwC96I+RynqIGKa6ncdSI85fYWAzTIS36dOv9RI3CDKEMfY2Aq1yLH78/x0ziu
SOa45q1D0pb4N95kewqbc6ZiZ9Ki+SbklPT1V4XecIdrd/00XDFQ6laZDMyQHC8K
AHJdUocDkSksuAyYTXzOgbxS3XcBsUgkS1wF92ABiXIKYoTgv4qvYMwHqA3q/6zW
+q0KHH2EoCyP695eiaKqBIMwxLQFrb36XNeMMnxpPt0UyrFDZiSpuW2CF2knMSHO
E4VGxc8PZMPhTnuG5KZwslLyG3n3KcO+G5oBPvyWiHhh6P85zCIi5hTX8KlistDp
vcOrTSSJ02+vpLxK/VvjtwIDCKbZGt/zVqFhDbO+lHVm4Bpu+iFfhGOs3DrU4BF5
QA0OcBzosbXXPHE6pdQiwrPnCO/FknGIbsyFW/xXCUrEHgEGovLUagAHedPSmMD+
RN0HTLsNUMcUj5U5LbQ8KskHoRIZekQzP4hAc91r1bxl6838jwVUAE9of1B0MuIX
/fklgGcAfEpUYqMwptYmW5riPiD67IU1RjLSF1v9rbYG7XtHb9qV+X3uTIXh1gvw
cOn6/wSt/TEm3PSW5d4RzJ8NtqWwh/aJ3v407vEhAneodIagIlYfMNmeVdHlT1zM
SwZgE4dO0bg6+kUm6khhuIjljahHg4TEaAZx6MX3/qkTe6Toym7kQWfZzBzwnihO
pwMcc44z7LCLcjwr7CEB3KEp++7t/LmKEnDLLlO02fRQajTUhnnK/i4xPwGi7zTV
`pragma protect end_protected
