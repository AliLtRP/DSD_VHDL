// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HtWxW/Ugb3cVNmhRa4B4tkv5QVoJvXgnVYyMwDI28Bii1vlt7jKM1vk434NnzJag
12Smi+eXxib4fKJ2ZD5cSioJpsXxmfi1oVg6Xzn3cBbOPynofuaoHsRtintaGFEd
7bo4dAYbIqWSsyq4DG5hkmLgmR7DwyWJsgjL7niq3KU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
rUF3X2ISbg/enKWTqhLjm7le0Judv4kV3pMrdJKRYEDgcABpIK/UcTO5JllzPnFk
7zbVuiyBuKxhNaEP6hQzkV2q272zJc5E4vBOywNSP8X3taHWWeuDY076sTCL/J4N
tuXwpJLiLpkWrbRtvAbpEpbcDsWIUoKrSD6r0Z2JRp+BOt1/L3H1aL5oIAd1l39d
szRwAnwAeUzG8ISiNOCyOYFdMJ76Gjn4ekQd62l4E/eXkZqqL5KguPJMesgtezxc
K0tGoYcwxCrUPl53KODIN+oRRiN4oQ5I0f/jRdyV09zhwjuZ5M+yp3UMUS2n6J/K
cJ+XWBrfqwSSomJ1tClKr+WEfUJ+3xzQ0RRz7vjyRDazIe/WzcA8sILJ22C63Oo4
8NPVSrC3JX6F3UmtEpHoG569nzIE3W9gBOHv4kJR2dpYvfvTOFw2IhdMB2fAS6fA
ypWJpcR8wXla91LC6HXnel0kvK41WfANot6spoN8I6JBRlzjkp6U67tvXfJrGtVz
o7rqGxiOwev8ePYmnwepUyqOpMt3jeYduv3HcK0bBYs4Gu5N17Q2Uj+C88l0VJUw
sG1YbQ4Fj0VJbPh93yS3P3TeEoNKw52ktZsZv9DqjlWYHaip8UOcUCjYV8puxebh
j/dMNW1bvkAZ4GkMQnxPsMkIpdKdGeMbE01HZJNPTJj69urcniOKVK6QTq/AhgS8
OWADREWbhJN3j04wNhPuAoGqKwi1SeuU2y6tgFKAg7y09yMALEbh/j30d4Xfz/Qh
4Haq6fUC1LfUk6mPb60qs8JzNSp0GhleOzO6xFlr64MCD5icOziRy9yTeA/06cj2
jYK+3r63U2i4ETlNhEa8BIf4Ela6EjraV0nk8ysmoWgDoGBbVo8NXlnaj3NHg7g8
2yKbtPnZhUVOqH7imyp3j+KJZf/iznK5FLFzPf4mMvpkBmrqP3CIWtVOYREbH29w
Z3JwFMzCyIBG2yZ5wIAa4tSEs/lYYBu1LWdpD341y151qnvcmaTUdL/iaxRngsfs
cBopUn91qIHOr9uR9WT57LQHX1ImLJmmIYGG20IXg7JbIGydxFKTh/9MKvRw2ViK
m18HvaHvCc1AlD7tw2skSQKxvfE5NxZsWCiYuJ85WM8ONwKZjoJgnw1Z2YrURUrA
eqjGEILvpVt4wOFUgSb55jEt64liP/bRKf1Pt1DXrGLRvJnr8cGD7jlTfQIOZ+h7
K5kn2hX3kJQBUkQ33oxOeV0QDtrGQU9Ygzhgqfz9qo6gB4gaiEyyy3ZOfIqqVZqj
j2+YV9PY8cuXs22dhPRRpIPItgBkBlj2rlHBkxnntx53B0n9bVEFJifD6Cxxyhkb
mTdxCzomE+aNGCrh0I/SPOplv/h/y1NRrT0kqDyM+HZj0NMhd4YExFcruzOn4LS/
fOcvD3XlVW5deAOHpK2j/YAcucABH4Xr9X2WJHYV7BmFpVvdlwFUJfaZgU9xLzTj
NvucWjEUQn8H880Xhw0QUDs5aWWM5syvKeLOowsM3ZGb4ypc3lT22Wpkz5+2Adx9
HEWpTUrL4ahr3fw5S6cROY8VSWhZo8YoAVl8akM6tWzC5Mn4ugCoLN+WQo6+NCBQ
M3POqyQB7RwTbxkpf1rlplSWpBzpgcrue7M3w6jn8Iv5UMz4W+NswVuWujA2v+YT
FR7E8Pbd24C7tAky4q7Nj1USRai3V3dquk+6+837NxNoyh5Ru7o0UjuFuCJSnWnG
DGPKX2AZMxM3HmcjPE1qsLw4t8KpL+RclBWW0rNJ1+71nujwXT5raUmd80ahWAKM
0ZrBV5cX4rsZOTTXUalI1TMmdMWuJuU+3UhSTdRxlbWGn9Mh22RJJeKwCP+6Wq6J
UdnMbMoIMlQsizkSLW/eaq4yBvjSlbJAKj4g5+Jl7gsV0TaPpu27WK9P0l5Z7d8Q
h3gOu0DXlbebJTelVRGteri/jq9/3ZIp2h1slvPPHUQF5r9etZwkCAtaH88p7SqP
t0ZFqqKrBqzzU53YluxtpqEZvdToYNqIY6AGEbh6CehAmxL8QD4HbyBj01UyP8+S
EORbW5uyHqV9YJphME9BSbozKLSjLGDchWc9X5ts47Wa3a+4AEzolsFXVNNReoQc
II88nj+I+dc+kJDGSSvszR8cy0Of5BAUTPmkd6ZmuUSeL9UXTOv4zkRAW7joQqum
ssbh32zIDxHK212USJ3XVYVeIi/6oMLssfgNkmyhKmI1oU5CFuVdO2btUUN0s+dM
S6p/lb8MorRbLsyVfrcluN0XvBcdBIqk96x0Cmt316vxt58OFv6luCQVs3Cbmn2w
umMyWvg8Wpoy0pDNPe0EK81kMNQL/Zxq9ffTuZGgsSq3eh1/2XZ0WcKnHM0pQPV4
qY/Llyuxvz2G+lKm//8qqwzbhMFGULOpBlFgHzHPlf/2/NSA9w5+Wn9tOZaImcbr
PuJyeCuGTczFjY9UurcumrTg7Y+XQWhn5Ho9GIGUXVK9ETwHApHOsFY+YaoDkp6B
mpMh2s0odoS9INWd7xBhlozLfUIbosL2MsW2N2wY7gPwMHo5IF07k4hezK/6uDwl
ROUOgvrWYcArlEe+sWXaQT0Ad6u0HVriCyJIMJkX76yn/hNpsr6H9uVjZc/i1AjF
mkOOkCoh9jRSGleRy6R2DaypJ+tVaAd75M55f9vFqBFSRAfUSVgbJfkMP6QXaq3s
JaTRFSKYzYs099La0Q3s44SXPKY/AZYjF52xEzdSDtvgEZgAn/wlxAZPYn3wQoyH
VAjt1xuWxjCil6foogALyH/LrPYT+BZx9Yv9lRy+0sHXoPPvvQRiTMf7fmGVbJtG
/XQK3QcA+L9TWeT68GA6eoSf1+6UCOhDiNllhHqwqZiVMbvGIh3n9cxqn9cuDo4l
6Qvc1d0XCzZzfmaH0gG8A2yrEozgRy6mF20DQKoaw0NlXe1GuMMY9rITD/WnxIeO
+vst+p4OumTFYiIi8MO9cqKcDd02n9YU0N0aDwh+TW5YKLkssEg8XlzgEmB9Jtvo
f/prTyAQBYMt3UG6PWmo9ebyw88kTzY3m+snqOFEMuU2WbOZEAzyEPTx+GEvN7WH
id6Y1oDt3jdfaEqUdKG94PuvvJvReABHgfFh+D0Px0ak1EtFN7wdJSnKUcIN1YsO
v3w44S6o7HvxyTQU1hB9N5VTIAn+wAgHZChKSwsePBj30HhBLR8wSFNURmJJjD78
QHAKj+fa95rNdzihDAk12rsxxpBhMMyhFR8PDk+64jI7Hm1H4Bf80Vz7RdSdLGDe
BKzY4mE0iulpRyt22hCUljQJRihf7gSPCLj9GaA98Nf6eMVzoZ5u7S4zLFqxMmi2
WQsTns/dFKVxRbr0mBVy+KekVeHTSri8nJOVMPK4mrqRjmvu7uyt+9C8Ac3VIrDA
d5SFtqT9GJewrwiIhXuHSfN6mWQFmHLb6Z+OH794CGL8e0tTyrmTY743if6AI2g8
3KOmtzMw+snGQPcwS650K+HFJ+Zck1t6aEG4XS2bqdUbOWNqZr+1DIbgmoItLoKR
XgMMLP9wO9mE4mPpv+NFpS7H75vVPGgUAJphvO4IF/UiKCh5VKWSaohHrm1SjZ1Q
Zl8gMQIGJHJYEkDpS497ZcSFcmBXq43wML1YQoxndYkmn9oA0R4R8VKz1Up60RHr
9pVier+FcCSvpA9V3Tc+5eS2VwMEMCF8LITodHqmdaF4lEzAVfBv5tAKpwNK8pGC
zCo+aFOJhNdVIjLubDQLeyoDlAid+tAuG00hmLfxgaPh62mK58BKbdT6YQm7vF2D
lAWkF74RRvnTFtft3VsdRx15OfijDNJMS7xK/Z++HOjzr0gQgSsT39AVuHM2hyU8
mBPfp1NfZqvrUdHjfZI/cMgE7/jBDYN1Mg1Vh5DgpTvpKzR5qazQ8AS/JSsxC7Uv
QcGe7e+sVy6o1J5f0GyXA4r+EvevTJ89wljmpq9C9c8IJvydjmOjakziKUOzYtnz
wi+JbN99DgfuJ+B/3Hk0YAOSawXCTPDZI+XyB79b2jCjP85UfzVo2ua8zgvZajEV
pCOA4r+ice3qOpGFkY3D4q37r7XZC6sDBVKae5MlBaF5hUco6l0065ck5Jb9QoaO
3Uoy/0M/jd76eu9A17fOXfQJJVbWEw7MYK9UJ+iFLW6olBBoMWJkidMXvN6ktBCN
htBX4rj6CqAp1Pl0eF+7k8Ij803dyhULPXTCJFZFa5NIySAQpQxSYbee86xWGwHD
AvYWQtcfRY5mZc9+kOWQ0o3Mc6TFSd/xHrCjErAy0YOiKurlBM079PWe7Jht54UV
dPrnr+/4pQq3lHFsqvOE2cOvElz1/UvO+8RLyEsl63uD/AK2ne0WJsLgX5S8pHVr
zpUelA/+5FB77jGYCA3VCJyHfXksI7IHVrfQSHiFJqdY2pQq82EufGrucicz8PZe
QbwHfMYp2Whprd79sq+cWIemgmWn0ZBcKjc+2X30uxQKoicCLRdu6NESv9kfyxds
NINB577WhrJe++Ek319qwiao0l0U4Om3sPwUQmtSo9ByFivQgd3i4DcncDhXAPno
DoVEI4aDh74gWrF4XJE3pe13nMsey+zajNlwX0ARHdo4Eoa6kgdoCMPHcfoY8UC8
CODt6YfRFRVjSdlrVEeX4WpTiWFEZwgI61YUhV/L7bXADHmIdMtTPklyaMUFTAwc
YQfju5dCAixlkRFRr/6AtAcdiG4FTIsctGmht2CzGhSBz5YNptvXjMArB8e/S1lS
ILsEfi8kqn3E7G4XOnLvsewxoyGydAsVZgXxh0tSJNNV45huKDqU2fHRGiJPVmvs
wpnKs5WFWdnBCRbz7hLP7DaG9CsaFu8TKMIVjyJBaiIfS4SweAQs0p5QH271Xz0Q
Y00a+MJeorS2BBc8BDgJP4oki+JHLXwEx4aPplVbFW4BzM9EIgtzJPcQz4BQ5Vhd
qElgaB2cstykhPkZqaOYA6AKUY3yAeANfBfNB8o3WpjfI9K1I2Kb8PKKsxPhsbmW
ASqFbJS2bpiOsDQrgn1n3VFo40ti5YP8B7Ml8vc25BFevo0vSdcrZ9Ed6f1xMnNT
1RquGFx742D0v+u7BcEIMyCliJJVCfdQyv/yEdhv3/If216cJxJvGcsZzvC4IiMG
1xc5h9PEcrOviUgdmEAEpDsvEp9nky2eDkJOJI0ZEA8OPRGX95zbQulfXPY8hbYH
PZRvaJ5S0+Gr6SF6k8oGtO6+aPmw+F+dJ1Oc0Bd8WfPzIn4AXYoCp0wt5k6vT96G
I9taQz0Y4QIafv9ec8YE/yvVZvX2mOP6MRwKAaAW+4n8tmQmJVSZbQVFxk6SIGPB
BZxPSC7hjJEevJ8cjP+bDMfkXvWzFApAKkqtLuxOPT71zfepStz3lOLFup+TZ7VZ
YEDldUIYsgexJYD6PavqsBvkeyxpXiFd+9IhF0ZC40pntZoB+U3xmG2cg23TrOBH
dTg3/Pin7FMt4SetMnw8pbgPKsshrxBR0P96M7Rfv3hJ9rSX92nZUOctuPm8hKqn
slPb5c8FynMLmM1IFspgZc7/rM6gS5hNkLek1UwSdXpdNcjgonn32/eOPCU4L2td
AziDfi2t7bkSLCLGrcHIcvTDPr4Tpj8GbaVy9YyLojOokWCSTIPbNv+voZnq477t
JVh++t1CEsXespE0VzhU2ihCI/vB8fIR0u3jgF9Md/0dJuW4tHLXfkArn69aCRGv
zb5GkQxiOWdrjfdmjuLBGZAZf7ynZiSbSjkQF5W7Stj29ebGLQ280l9Q1pS3D++4
rEYcoO59Y7HDd7x+G5IOSNeaJPt1iSfI7g59voO1Kqxt56wAdu+Y8NUD5YEtoe9/
IupViRHbCLfKpdmrBtDWldZHHAFoxdCEUp+1vtz8RcH+kfJ60/DlE1zVpbBE2VKD
wbJ5c2oRo/2bPIiplvCbm0MQzZ3qtVVtCdbCWLJdpmzGJ9TzjR72O6NbhBHdFZsO
D0QjcaCJ1VzmJ4doHzMP/uhU+NFBsR+wCKqi/wUr/neFqmyKRK4qcDiaZJXxt1lU
qKRbSGp9sjqNyPG5e8TMauuLMrMtTBZikuH3n9NM+dItud3ak88oo4RExiNpnoBW
9i/X/8+AGbsywF0hLAoIPDpyaRo1ivtz+CKiG0Owx60Z0v8ccwy9OPCwJWyIV9CR
yH/uEbiZdboPvu0c+SNHA7p5lwNSqHq/uhXk85mEmhrBVeox2LXf8Bkf4IM8ByNC
5DkpfDXOx6rOQMAl6FUH/zTrH/9wjkClsavswh30LKFNSKwhsOC4W2X6d/Y/2G53
pi72XyYSD4jvu1b+K8msuVGN3IFd1ejB0lfXWd8+Y4L8q4XCsmK084CFNR4uq56n
Vq+vR01r2syDJhjLDc6Rn0Iy39XISkRJo0ALt+sa8DDlBVI/swAAyilmkQOJMo10
ukr9tqGjEQgc0MTKDo3D2EEv8BvSu2/PBdezbWqOX1lKlSzA3x1T+ijpwgfS02lP
POs/LynLyVWbInrzPM8GP+8kTImO6+DPJg8kQB+IFtOyaH9WE5kLdiE7lnscpzkS
omJUDrs0Go8WY14eZ3aqCJ46dNr3nY1IJ0QQE5eu/W56q6nyD7YcvCtwBaEiicKe
yx7nPKhBq0N6nhs2bu7OGcFy4H+bz2t8I5dPIJavfp6DWcPtpUWwUlIiGpzBZe0L
DR7WEwTpFlEQqDKlOFgcFpVsn2590xuBJoiPVHGbFbhtVyK2HX1M7njbm4RqEKS3
ofKVu784ZJdllTFgMRPacLDBnLtCyEqWxZLfuf+xcaUxkk+SIwueh04YF6M/ivOm
8xTavSDMQ0uU23b/ZIHmc6/c8xMYxrHQcZD0j4PfujZqgQOGyx+LZ7kvV/zqQ/e0
1gtCjbPIs+vXwUvg+BB4GaEuFBYaQoNbFriu0+lAVfQDWol/G0Sa3E17T4EG1qem
oAZmusrNyjg5tpn1FJ6Kwqu7aZbn6C2Wug3npRbBEZmjI4KJ0aPBfiWnpBj4bgCE
XKSVwvUtdltNYwsfxeT/2oPnj2NaIyGqDgFxU8A5hv4wzmkWRhiggZ4sixEMEdtc
ks6c34TerOnrGskGhUH3RCN5BUYoDyTCFrhgcJXrd6+jyTbOW07vOIwY+fvxQDWW
6FbTTbxDcAjI2vMN1MUfj6akejvecE1VrXgDvhL1BGPo3tFuXr1RBvvBN1DDYoeQ
diqNOn9G7ORsUVQtw5slHtzVWZy91SX5VrqtqAQunXy5Jdn4PXj0qIgMTVns92fO
rbjF7YVOhDbWMhetHnxU+yqt/UFh1NV8FozoaYtptvzuszghl7JNVW8eBraJQHZF
+bv53bUJ3+pblAuTNx/KMo4DLCvVGLjHOQwVL9ZIQjKqcLnv4DxKoF80NkavHKqz
KN/9c2iQNrrVybs6955aK4OoG/eQKlwCB0RuHIC0YwRYoX4MqYilBZuTf09t9kdx
3uQxWjZB0RzvhnVnaELopQBtdNiKnR8OBZSEKTRVIntjWEhA7xgnLNL1NnX17smq
UNpJaQJTDac/UfznKN3VBftWJh9ldBumYFx0TGry76HD0YchSApU0p4Xh8v5tHwr
pHltRne8ZXxoPChaoQRT1Z76z4NEOXuWoyjmmw+SnqVtrGvCus2F3RUF3uEHSECh
896c3zGu9V0TYc41iSr5WLqsgi2b1kV3+fEKTHou567752/ozZNIcOJqS6/A5mrk
cIvObr/EGDDIX3XyM00v0dYz1s0kCTKhhK91YSTTDjLx6MYQMyZ0c4KYpwOQGay9
FpvZ7MirHsmEHauzpG4CgMydWEGu7Y2cAiBtPDgkTqXfAj04lDu35AZktK2k0fCd
St32afWG+n6vzk8kAPM0JZDbxDAgmPw0/KVC65oHCVmOTdLji+DtHf1r6ycKTd7M
RnwzRJcl86srV11/SRBHJ1a9qkX34Lk3DLdTCOBjTprpwipI6JoA5JJ0DqHRNjcQ
0vytKeOk80aIreHPAWEUGS3EGoImrnUk1omx0meA/hE11FwG7jsGT7YEEy3PLzPz
03G2pHGa5VeC5DyaWEfv2QXnHbkc8qq9VP/NXZiGI/QauDixcSY2MMdUTymS/QeM
zyRVojfx5ekYHYuEcDjMj22VP2XKimusl6U9HFpt85sq6wFmwWF2EEMJYfctOH45
FZ/uieaJ1d9viN31MiRP1ikNBgxk5kpn6GP2aSBHM/eXolyWSYHGZeY6KvK6n2Lv
udZj/rmppHeZbZ51OrwnTvam5W8X4lEi/Lt39CY4SlQb85kMV/Bpz3hkbWcTJ2CR
ulmxtrDX5n2XpnD1+0nqGkgo+GDWP6lEMqJ5QSyfhU2piTjFTFSNy3PI7wjl0oCa
vdWEGlJ7sexq59cYKfkLR8ww5ci6lwffyYZ0axX8YOwKL94d3ex9cWN0n2dDaoZk
747Rvvpso8vqciNqlyIyP9O+TKGOtTVj2PY5gq+W6V9QIFllRqCAh7CiNcTJjl1y
Drmd9ASY5QvMsdELVdmlk920LX8gVRLJbWdpfV8HB5vIh6qRm9AOclo8mQ+EXNi4
p2MK6B9LlqjR6LdJntBTcORNFbH4SUTWEpGFo+WCzjJT8igWgOcsvbyBv1CFf0JQ
OklHqtgLcxrNlFkmpyyUjjExPC6VRR3a4AejM2/imj86wf0gzv/GHTZ7kwNxMeaH
9hENmIL/BEvVXs3SnoDGVzUvFde/oCblmhSQMdowjIRU/OKBeQQfb6CAXWvGI9+X
Y/9RwrRwgFvBfqTaDOcCk1nHVL1jn6khItdypxoPXvNu3kT5YVd5bsogDbigpC2V
mfVeWva8nFWif0MhloYyY7nTjqbODxZKveJroj/LyWkM1ErQMCGFErYjjhBwMGqe
2EsraDIHSnhZ3GihAs7z+8oDHBBr7pAnN6WhXYnyr2+yxq+078dMRC2+0kZEc1wd
KU4OoZRz4HSFasY0ycDAXjvT4XAobL/i4+AfGbFzTt0Vt562u8a/I/ThTvyZwcww
vmEpKRc33Z8NtXHUC7MLK2HwmXL7w4YFKYFt7OAnqiY/gWcazfoZPAL7xfgrlmyV
gPuxcsNWVUo0iPGSXlPTqu007dhHfeaoW6yQs9pjL5ApI4EG63uJPmqmizl/5zsf
v2CzDJt6+NDHkP0hXa7Yiq8qLBKEF0pIFw3EoQBAJm3A2hezVrABR5Y7kfhGC/a+
BGDiTGH4u7vmIC8qrGmVckkq2oiWpeq/bwpFbZ5TFnEDM1VrFqj5m9ZNgNEO45OU
keApulghPgJLmotwNuZCaER2Fck0n3IfPx8aYEbfSsvUCGBDLdBe6o/qOkoasE0o
ySsPAk0b/p+K/i4QJNCwPEiyNRz4OjcHWK9g4HLNbGQfGuiPiLx3ELXkQy6rgT6Y
VQBGXsRqwetbi6jfudB6jiRbi5uj4Jtjpr12Snrmkoz7kpkRdLj1usSFyyj7obHJ
LTQbvd0kMQfMSNMYWP3WRK/lHWdj+UKHiVfc7X07YDUm/L2K+p1GhweWKvy0BG3M
7UZMomkhBw+pcSbqh2Q75n178KLd1aoZIjbQk9+L12kn7bnbGJ1aZvQpXGfR3VMg
Md8v2OZ6YW1vn+DZnWehsnjknvSFtjGiv0xRw7AaoVOqw5Mi4v7bAe977sY2CuXb
upEYCwaiz4m53dv8hJsyzW9t2nIzg+etwhSCfu8LCGRn4weJY16x8JDR4wypK8jO
tvTYxH5jnEhBYbL4tnpBpCFZKVKyS/NO0H05ONsi0V6dGRU8jTFfmhv38ofEvTYV
g5GOJoce+PkCXAJTqNyw1tI3SfalyoYhZ5NjRicfqb7QK5pGYhWY6gY70DYSpQwx
jOzKlWcjXgj5FODhadqq8eI0nUF2fDPhMHFl3vDH7iHYs+754AOeJAC3WonrASBL
a540Oq3srqqfqAHERo5D9cCeovukTpxr759uKQWeu/5yvbDnnoqod1nPmGNHknkX
tRzW4ieCkXYC4ETPRMZRyR9dxRysIIwOySDazzfgrMuBqdicvG26SYjUYix86K1G
hIbLxEeVkjwcoNlSgxZkAGgP38hw9e/yEomw8M2n0v1S2ogXbW7qjUuZFF6Gqz/N
L66jwGJ1R01o29pQrfW3iA9XbZSExnMrB8DA3+GTy9hWLPq2AO3mqJnmWhqJwML5
MaFaZ3soz0FQWW1s4NKCuZAKKs3zYMjtbcLs6XmxGWRbepILbrs/tOyVysCX+9hN
641g+iZOLwaG3TIWMMzuBFtXNLz2WGcS8+PlSyFFn/AmfMTO8kGvFTj4FFlBtnF3
EgnNUvEI1qz5MuVn20Ib0M8Ftr20rummvK/ju5gqAlQF+M5hCNYGISpIgN/TWGNT
Q9izC9Sd/0Dngr0D7WeGQi6bwotuZGMr0Gce6yOzPq1gNs10sisXNeZyJR9ti7Nr
wyKsxpB9Xm3zkWLj/5LqT6fBDTFfWimOqkXmkgU37jhK+YQz31diylWcGxUN16Bt
Wr/RvCeLrg58OUzKcIIjVkseLMvvepMLP/Ice/EOfu68y20ua3Fol8cDtXA2O4OO
scViaO0nMDHFjyGm/rmoUEQH243+ajazZAT8nniTl0gd0Eh9SV5p8TNfuYFOKDDG
RL2y/WJojm4rwc7W89tukaDPZKrNEAsPFOfTucTz7Q1KA4C4Ax3bfqBJoU8zY3gD
ZzwfN3XzIiUtD41vGE8e/ZSx7NEYTcC1yYaItN3+HhDGaldeENXStQby9R+/ostx
Iy/LYCTMKiGA0G4UeX/7eSjuOt9g22pDay4PRKr5N/XOQAxGe4TvJVKqutW9Cdde
Xpo0CR72q8Gcx28V15L2WeXwHFAYT4RPl4XO71UisF9hvyfsZePVAYJrdSr+Sr8q
L+IiS3ko35R0R1cIyZ0VwvzBErz9WWOtG9f1GT9La7aox7Ybf64f2IMCJfDnClEF
VxwxRLJCT3slZ7txU+ELi+vuNv0zjmewpQ4tueKZBHY31ZemLphvb26EbmoqSa9C
3P64srSYQQ6YlrvGEkqjxElz9/QMNpgUj/iqMrGI7mQy8rr+HSUTrAzRWW5QkRnz
wvW+lwqp8Ina0pekqbO+KTAF/NUZ9LNKi9uDyY2RXOl2UOamdkdMiDc2MEzN0e7F
tXqdzAcBQLyKNBBgJxJs6Yf5cVT3B9WkFvU8gcIoBHaPWWezLftwMeU9Dl1zzT64
zUrHSLsiI9M/DAk8ASqEUbR0pNABCEW5rgmoyYmjuTzPU6oDZT6mw6daFOm8dJPR
qGK9R1OKiGhi4Dm2x7HawQhUVTZL28HSDNcphdq/LK7FmuoeN/EGbyiIkP3X2Iwm
dCtm4LCRiQabuQZ89i8Mz0grlRANNXNkutAuY77wcYzND3uJV2mrU7ALJSKarnRq
Aghid15RRK80O4PcddZNlT6g5rXhGZkxucxeFrkl1kXajOMCac8MDflABQ4l7rbQ
gN3Mn8qOR3QsvJE0Y7L/TrUbji83pYqHf0NXVgxGFnvNs6o5NLtS7Srk1cwmC+15
+vhC6tNMhAnsNg1F1ty2+3S0uFT5o9fadR4JXC1fSZnMJOqLV1Rm1McO4WMtAXae
WewcCGQ+pLj9a6RNh3EekpRfOYgKtpX/8X8AguFdXyiztwphpJ7x8hDG8X7cMnV6
N73olbq9UUEQ9iEIzeZx93nFPRee1r96kYh8SGh7Tnncc9auhVPRYRMabG3qMAOm
3KK+o4Ig84a1eArva71zZVYWp1Q84iRdT8c7cwlie5PkXeBbnBx123YwRhlTHCVu
qOT2M83b+JAVdhWz22/bwGVfWw+6rkSXXNQXhFWjsPmGLpvMVM2ZVkxXYRN8NjET
DzCYJFOSsQ6Gr4Iw9MXNhHsyG5QgADdkYA0YVBOGw2VqNKKg/9vkYehkZIp7kt5f
VCI4yWG9qxP0BY9iqy664wnKVUylDxkAwnQVMK4T3ttRia2osA+6KYQg8rMCsxpG
kIT2Nlbh89SJaz9ckWsjadhWLzTIo2YR4K++UDC78tg3N5x5UVxQf8ASiOrmse2A
GPufL3xd7zDT0m1opIv+CC4Id3AMLS+8/vq7T+8RrCAi/nY/eNiGYRg9MPgXi0vr
EGOfKMEce4cmJ336Cz2OiGNmKngyzNWKx8avUY04pPJlxE9XdWB3BIaQehPzkfDr
j9hO8ywkWTHOAL1SMd4BJhwuZwZv71Uryw5ZMwyIvm0phWAQQ92T9n7jpuYzDaZj
Kr8EOqGc2SOUNF4n5oOFsLlWPBdcWj9ugDWLTliJv2l3l/7kyNqn9T37uof7uvLe
d/kA7WiIg3smMWU6+tOcwrQ6PGpleTwv1GJrTbKwjBMKlgrkfC/sWXasMc+WE1Bs
yzu/Rj8e5WuGYy9u50edd7PEdIu0C2WjQkx1wpssVScSBjZXfpjbXsdwBmjoUf5o
9u0lFILMmb1ZPyshvSSrUSvmZg0IA4hVA58m3HqPnizgYC8qxgsJjpKXc9Zl7CVV
CPzzL6a+W9cr3dU2mGIn/NaWqAxSZ0fbDmNC3Ay9/wPIW16VinJJ7VffC4tF8m6B
vYr3CII+qyfbneM6CC8kZsPUd9BNrsOaX00BUntPPleQx3c0bfWVJff7CBouvlPs
s2tU54WjCGvCXUp25x47w4S3yVmLCpYKz+E4+FlhA5edaEGGw12YrLZXferDYSh0
hLbGFoIUTyo3TC502/jyAuzu/d2KDHrDDT8nnxDs7jOK7qFy9L5p9BbW3G/ob9fr
n4wLoLbaq6V6wTcoOE3GvzKQ8mqTr5P8Zu1SrFag3WbBOgp84JCkY7vNaH2n7qrj
18VTqGrejGnAVwNu0LSHqY5O0sjUiJHZ2mUfGxL4rNnGR4+B31GcusfmI4XW/LNV
uBpZj4ssyvckUSrOh6H2atXz5L5qpCQnt2uN/eSMG8YkINNO2jtpL1UcmRrvoZmH
X7Ke+VzWE00utMz+s2K9j3UgzP7qcqoRUtJf66HribvkbLQCEyYLT6YZghmxRaus
lOOLbFDs1sUw/bclluuimqjnoICKzXLbS5uXgHVwWz7RhIbIAzWQgWO/RprMnHb3
m8LytAKurBvh5ZtYG5uElDZ/z9p1zu+UmmpnOMJbkMuMVMIUw9K0rG5ZjwihY+Y+
rjX/t2fKTV5QzAlxcUYUpnK5RzI7cKNVp6O60K/HqN5P8zpNsy/A6XOhrV9glQ9w
16jEFb99TXF7CtmSzlgnG8p9WcfFhaH7X2DUmhC4nmMl3219xO9G/OuYxm/LTNJg
ArggTVR+66ZliqkZn+q0AHSkdhCumZd/aSMblyJNEokfqSAPm9H3DVNSNCp/NhzG
wSo+ltRak3gzZ/KlPY/NvSz8/9afn4Ow6s5Lq57CQsGCSdcFVnTj/+aL7i/e05C0
FYWglns8R9EJNJwWTUN6Pyv3QGWmcpy2g3iwM/fdDNHlgc3zzbu/wrkgPXxjZXMQ
pAt5cYULixWqbZiaMrExx8Q5LCzL1HIVn6HZG4MIzea2bWbAQ2HdpqSVWDL8dJJB
+LhLHir6ER91oJUqA8kez6ITTT/bnRH0sjg/OnwDgCn2m46/wjmMWiO+33M1txhh
+/AgbTTcjqKlPGV73oa0huBOhNOPHNSmQbQiN3UkFfflKULCXpFUP9Sh0fw3RvVf
w0jMTcLq3dHb2NfOfw9/B53lmRDGIv8aosBQdGJF/MTOof7MAUY7kwnPRODPREND
3fcMe3DlqYe+31eEoTTbzZ0OsC1zS6mIa5d2AftC8vAmdPNTgW5QXuD4+4k7LdkH
cBdW1KK5IhdF0XhvcAHJ2atAGuuIjLYsTOBammeK/0VF+MY8/VpCmREy5N4/k+zu
bSjO4Qam+4ehcABheucPnMSNyBsL6Li5bgYeBdoguMuLSXT88LXkUozWJcqLkohu
yigIKJ/fbsfAHCO6iD0jhUoJKhASOQml0crOLokKLfrOeAjLq4sMpcshLnGofjhv
RQFJlD9IKj4Ytz2zcWMRgXb+WW5cMepPBqcHQKk31/T4pMVCCZZQ2nGCAMaAdEba
EC4DUxvaaJhybysqUIYVyBWnUOJK9HEeDvpEaUPpGU0kD+e3sA8oxfaC9m6q5e2x
m4RSr4+GLQJJW4dagNlsd9kd4TUfyflydlv2Xkj1QkZcXpbdbB51tUfk0acw0G8o
RpevcPda7YuOEtubYvn8q1sus3AZwrMsG60GPhwqv8+pC4+MwA4RpXd39NfiWPWF
+S+arILcrN6+N3+lmzms8hkHG/QTM1opjF86RMnJQlbhmMewhXNbT4b+mSBye9UV
ifvZ9v9ErEpN01GNAtvRYM1v3M7V775xs5UUBcBbSaEE/l4dj07ug5wzM4MYgsEK
I7ttRxVd6DObBqgD4It5eMwtH/jF7Qd4XWGcdF2tCXlyE1URfMi6dMQ8zkQhiAxf
EyhQW+wTWrXG0i7R6Z4Kpd777ixjZwvltxiuoirdqG4Uo6ap2XRazqF4pAEter3j
5ju6wCcT+nYHNl06QgEQwAIhkkyxfm5qEUsj0f+LQoRHegx8i+hiOF+qwFspavv8
FPDlc//wrEAO18Nr4R8br8jslrTlZf8XmixF/4pWZB4Ih37IaDTlq7FQuxRHlQbu
9sAtgOX0rmzNJsjsLU9AH2KO64FPKb1Vbn5DkS7AKA0zOOGWdqhBQa5N18O15fbS
I/T9nn56GSDxWBbV8jYC9RM1sf6vGhbF7peyWTT/VcuU9QEnd3+aYe4G/eUXVeck
P/qecw0n3oQch9gQhdX2wHz6xcq90gwg1WIvEIRVBpZLZxGrsBJQPHn5GLNZLxjG
vi10420GZv+wpEl6Ejmtp4/66XQ3zRvfYWw0cCLrVXdqWtJ4/VrO+ahPJ6ZK+mVq
/8ynUxImtruELXxnB3czTKerWw1wyQ+0rN98/9sL4Cnu/XqiryOfhL0hyUIqVPRp
azxT13we7XvvDJ1ggph4hLvoxQnwaUv5rxNg8CUhRho/scLj5ypFKRMvCsEBatw8
kKn1xRePRwxAdg5yOpGvEHuAD6Mvpf/FGE1yQlDCb++TmnkNguXKEhNEiQf0gVZG
Y6zEbrm3za7Pc+SiCRBS5eDuzWP81jGcE69K5GF+4wXDqtufGRgaV5PbfXE/DLPe
vMWg6Xq9kFRUbqyz1z0e6nJHD7TOtiBv48CsuizDJAeKWzMSXOGBVIrfTDzi4pbr
MhxvC7E3c1BQHvKSKhUV/+VtTPOkjxMzWGlvuc3jxFxevY52Y+HczmY2OfbB6e+4
6h977ET7e0ioJO7751Uff0zMum8X8AElSMms+gegHdqqhrdZuwOfBLBm/wiBdSiW
aBMi9nQt/3ipnX4iuZSaCXpqIxNl1U4eGqcH5FFHWlt+ONQaPTQTzameMNmjkC4M
1HfyxVswTzlIImLe/oSE4+cMO6CtwR/0iQXXdlNwX/NDAqztyo/C13YFbtpLiESx
yDr9XdWN3sjiFxlKEE6aQAROR+5Jt+KZ1FOSmHC5qmZWcgPQxTNm9/g5KGVQmyef
GUzM39OQCdWTemFHScl3JrBUcDrSC22wfv0yj2dERM3l+MiHRFdH9+7JEQi4jBHR
j+Uf36pLQzVhyu9X5UxP0m884ZATt9N1zqNCgUHS54NRwuuKN74l/QsW/T6Nebe2
8e5IDUPlVXvcPXodmEECZP0oekJd9p1ER6ToqKsXxQk4Ni98XAGjX1RwehH/hrRB
b0qiwvCXHRpoBPTIiXbFkpunYuwF8SFTxygjP0laO09Fc3KEN58ceXhuHqtIm0j6
uLS8J8/LSbKuu8CorcMwjDQVtUtprxzPGBYs5dx3k/foXfmUT3J1xltgqWJsB39j
63ZaRxyqZGLMD+QsXokzZ5Wfyx5I/dmRPn+X9wQWx0dQ/firNu7BiUiv80O6sZp0
Evf3gwiq4NIRPb1dWPg2Hr64xUFiZvVNbljW/emeYFMy0gpi9L7FbfAxve/fMbT/
ZpqH4FxZdmXUQts0IDkI4qzI6MZFEMeAoKwqDis3VSHZkTcx3GEX1C7Hba2mGstX
3nlWlHv2gbVaBHFVPvnjAqap4y8gSrUurOw5OgARDF2K9MUhZrvvYmzX2Dkqzyxh
9NY43xc+yoz3U2owitcmPXr5m4qhM3g8Mj3KgrO2LZn65q3hVWN3PkcMtVKsOAr7
FTxouHQWrrMVY3FY2LA9cFseLd+CeGmCKAVMRzLfvzsV4c3sekJAc3AtMa5Bkupl
vMgExIo0lmG6gY9AH5tXmQ5nlruZzA9kI9DgiWaQA0XNLb798UrwZ8MN/WBK+2NJ
Z2p4uhocZCZNNs8aAIEpqspK5jipSQw2t9NRcl0cI8E/2BzfjwqLGT7rcUqevSPc
EkII+d8pNUvwQPLfjJ/gggV8tLBbkPYEsmTOVg6nI7XU0TOJ3vTpW1T8egqPHWeQ
kUyJtE6fbyLIPPDTM8eju423xatscdy6N20ifyQnKKXQ1B6+NY3ELEPam1pbqxBA
wab8vx14xugYPKwlp5U+E3J7SO5iFHCTXaYo09Vlz0txA5EMIJNETj2Yf7jcGB5Z
oxbqBNRNzNKqpWtNwqnaryKZz1aFWxP0002NGwKESYaS1MuL0ySAH20OPXL8ZZZg
ve/n/hWW8M42lDOEa/qF/DmWWVHZa5CykgCVWlPe65Gp46QnrI87uFzClQFX+ceZ
k2AlETP0XyE3Wqj2oKDVtMI6/ROPuLwUS5Tg7AS5X/qQnOKYuUrVKAVu7BojO86t
NQJeblBcV6cdHbSbwVeD0ETUPjfVooxG7DBkXY6YKLHZwdg8Ugm1SZEU/vc4yCBb
EQieILwmXw9wJX8sOCCdSly3Z/ACvFALRNlS1L87Hym5hJsflxWrMIswu1tMo/Ha
ZAwkH2SEPP4LLx2VMgGfhjmfJH5eLz++94m4P1S2czbwFozex1hY9BVyWUsSOrXH
Q+D0eYXvs0pTJxqN06f/y8YYYSQ1FPCa1bclW6/M3+2tVPGyqWM4lSHk4c+QO4Tr
QQQ34E4pTacqMhJlV6Bt3heEBw2BSoXcOlqjLKT1sO2XEgase26m2gSdUtMhKcT7
2QCvwK7WyJMjRpEA/4ma/dHEGKMvFKQZ6Gnws/Ft/0UsmoNkf3majEZFb/YdjRqR
2DJVB6XNwPkNmlsyGoNPxRmHkF4fT39niziUK+2UkcY2hLOR+dNk56vlE0auGt1P
Lplot3zeRMH+eVWyudExTBL5ICe8NuX1uh0b6RKFi8d2woAl9FZjNqnhmFjNnQWU
agPmicvoSeugjf1ItP3fZGoqloBWqo7DYnprYtm4ziq1vWUqXz5+1pXIYW1xk4Hg
xZlGQYvmWhgeXHFGZtM/KXx6nxykPZUFDikjCNOpup4Sqolf3OZaFChAwA1NP6ei
oxYNzEsSmos3JdjxKize5RSCdHTXH4APBu2N/xZooJ8+RSzQjcM6aGwW1nA+/avv
1ZYbTxC96bRodYRKOQkl8l7KADOUH7YHrCr/JsB+MgE+ypWn04rEolIcb45hQLBF
kECmuAlk8fdZlEuneJEhcNbPi6TH1UJoCfvALM01UEb7V/wo6zv779s6HnULoDli
QbszSWMqOipiB1JD6SMibSN0O+PW65TDUsTDzs1sc4cynA8Lel8ldf5Iw4tcFv8B
fRECygAE//oMtnQPSRoqiZm7/gQI5UXipSe+vfLwFAv44cFhsfSTSaQhziuxW0p2
kyB8O2MQKpRvGnp2yukshMcAsHAVFvGT9+UHv8g2JbibfwZ7dsrPVj/1K6bvnnMP
9np2csCDHJ8MjURgleZFtz0+VEp6emkO8v9WbdwppbUYpsrfDDS65/aYi7xnk80Z
/Fn1W9NXW9QM3sdyiy50b8V11AZ5UFZj0j+pjYFXEaDjjouRzb2mDF5i23QqhhCK
+2OBHZNTLshOn5mhWtaVuI0kqz5do/BrpWTg5JQ/1afiiXYVH5r5HuLq+vmQLN4q
NrBEU+fx4IwxxpzEWLwDSS2CYrnmC+InNWwx3zkHFII80ojGfhyuysYhck7jnLLK
fl7bUWMsNNE58zc8utW7uaCxLjhSAjLxFzWhD+XFotNxqqhxbJf5Knosv6XEM65Q
oDskBriIleIs6ItOHvUZazJIGTwCud6BOBOiOD92bCUKu5O34jkLitlkrEqn8Tql
fYeWSqLusFpFOejsFwgwAOZX+kRcoNHciztuXbyfZP+xs6ZdNMSxx3RtMmRJQzLH
k9Ul657K5K1rTD/SaQMqKtsbDECVUXaSFWXlpCcTQBqlKY0WW8293vtdRwrXY60T
N45J6D8f8vDru7CrAHzdE/SY4zW0Gh8nbMs4Oe64Z8a2lg7vwCoGYUdIB/6EZntu
03Z7GyNepie/PVAkrAKsH9aEpw7lO39IP+p4Ntc3p0Z7wKQ0gxLOTn7UFAwI9lI7
BmR4+HkiiiIiRTarn/RMTGlGGoy7lb+OgohIvdQJivnPrk2XsQ38Hc51nc67AXdz
WxnLx5ZVwmt2UKi0Lx/2hQqSgLHgUPIDazDwOxfmgnDIyJMl94CQjQT9cgiNnCxo
Xz7QAEZ7mnwyF8lXaQ7iWz72/oEhzb/kDNaifsFtvNj5E3EPQaPl/fX9px4kf78a
xQ8WGoH8z91LUYqb0BF8jkVJTZeUsvHTr4XSrt6chetCiXreS5FbzMn4P3XLAOc6
I9ciSd2LkEUfdZjHEV6EULYBG50A5RccWbSaJTaZxdcbVXjSX2IPk0IbzswkDHSJ
pQFB8P29JTZFzbTdGuBGP30QsiUJJpQH4LdROe2i47aPsfUr8kAptIrpoKMnsF8a
cgPYwNXtR2dSxYCuNzzSgbnr+jURwvW6OrEdNyVvdwBqsdE/h09FfPY4T50rVIMJ
hRKR/aw9giX5zLxH68RDZDDJhV5Yyp5DLCdUa8zL3iT5rRAroGuyrBmfsSBwDeQA
pRdImjxNGbyBfpTBwgchrhP5g6co9RVDDg7632S4BpvpL0+XHFH4o4F6IHs5Amr5
Zv34MRZhRS1XGBk84s5bB+Ls4fjKAQVfWmZoTjob2MV8tDpsl112n/607u5zIy7F
esyNTbiz9cgHeEiLMf5QtP/XvFbh95RGaiHmwoA8aB1NZrrMDXOct7hvCGkBn6MO
F++CV1Z0X5sZGDXsg/SmCYCha/mmhGnW2Jv5zw5l1K3sqyLq37+QkLmZYfSDfmLV
+PLxs+UyB5tkxZPVxMvpUgyLhPH4HxR55OVx29psjKrCp3KGwUvlLRjCBvuIIMYO
wpHGUlyZy6CgtcZ4FyA0kYrM6oJdvHlKksASFMBxASVJenV/NhpQ9ye050uvBFal
xNLJieL6IKjYaw2n43PeyfZeHzcqSkjYxfdRpzkuZ5h5uYcfmGuDdldw0Iujvi5J
TNhpSfM1/RNNImrJWTISjKUAveaOj1O+0NmzqXTXYUtTDJllFBis7DPG/DFU66Qb
f3wauuOpncBAsc0H1Zq3mqFiG9ygbZDGb/44MAbaVNoNz13pzyZn4P4SZExRSP4d
TUXJfhDvDiMD08Dal+qn/zcy8DliqQmEOk5nhAr7PpUbGSlXqLhKPY4q6z2fae3j
n96rPMT452Kqh6nPhgpwo0xB2V48b2hSe4J904NjQVPoGC4H2yBumdUHNBPgxvox
YsctjwOZIbzk3+6KEIw1+fj31kmdtjvfnzkBrWqS2jjDT4RfrtuoJX9+AcI922Pm
feBWlbV3RDEPehy/6sYDDSSCG9LSBxPt6n5D2Sng0JSHrNz9qMhDaVYRdtS5dq83
HHaclWh1t9BCvErpdbMB3V11dwNjwDfh5P36gjs00kVvKQoAKftxxiLUYgiTiR70
JNQ95kIfisWDdiB4l2P6tC2pMb/YTjcvb6XKJBV3T9hkv/B/KJp77c+1LMzftyR9
/01W1M0w1EFKH1DPfrUZh4sTBidJTwnntY3Xb1TZNRwVC0CxryJUM1ZwddEGX2Mo
VMZGIysEhK3GL+KXpo0/XOrlfm9SqdXGTOmpF7UwakJUsmdHs+wrRu8mUxS1N7AE
uKrTLAR70xLFtXEx1tEeMIc4BNitGyLacrPJsTHglVEbufWb6nRcsx7xs3thAAFl
3UjroARLrBZs45bNLhwi8pHA284J5hwiYUvVZ1VqOCAKY34Yty+Ymk9WZIDDbQm2
xLIxVcYFuRYpGF0JThr8reqJeRDX8wOPoZeORl5W7aQgF605JfUqp9iZpvPbwVb2
F9rZZpt5ii0YKEph6i1OY+mvCmwDmvvn2Npat8v++eC+xeK3PNS65AsEeLew4BLW
Df2ikg4EkxFjTHzycbiRk01bJOPI4BImQcFovYeaCOSmiDlt+PKduomj9XPWfERW
ozfFrgWbDvCIkXpgRq6XUZ4k34ANPh8fEtgwHIYN99Q/K0XV7Oou35S7DKDkmvHJ
JzFy/uJjUKm8vNZEqCy1FBc7OOZwHyiGe/jXuXPui159GAk898qDxHd1e2Y8S3LC
2ux9c7vAuww0pyNO3W+ZPBjvKyCcp5xIjc6GV6qwbwTaNLmjO72XfmvHl8T1mMJW
54p+CWhdIw/3x/Z0+9L4HLkIitxnNERmtUAK3CxKtDcuGsE+VuoNSTBSGzyN1eU0
UawNq15gGabQyxgm4JXcOpwm26G+QKFg5+rwZlGarIREmkUkuvprslJwvAp+jR7i
Oy63fvurbVgGV3opZmPLjOGX7wxAj6A5BM9YC2r7VrLw6oJr86NaZNSMfq7lc6Hv
K6cUX4SKrS+KwwgeKla3qOgj4s4zcemC0Xb8amEkVx1d0bP5HGxFSfKz0uNOi1R/
6nZctjWtdxPNxYeCbooPJptNwWM5Rd1lWUsAbXhrdMeDw1s3LlXrHc5+p9QYO+DS
kSDca/toDA5NAdH9Jyawn1kDll3jr7xmOGRkqFF65T2d4iphnTek7GKT1TPpQI4M
O8eRCduLI063aINaXsYOaH4bQ+C6lzE4v7U//gSac7tkTi0wfI2gHUtSZQha1Uuy
rHOeht6nlXWWt7Dv752uBm2Uh2L4vyjbw7ElwH6JxiDGyOb3VqgjR1D/4C3EAdXn
6IgtQY+lsmBzSCAyVF+mZUfxWyGWrxdSM6anwQ6UYrW1WzwFq/l/o5WHi1ZAvlGs
pF7kp30YSHeZ4BEUthgpjgh3brSWI8Y1loaic0s7tKCMTRESY1/jia1XkrUKgGZg
sPKsa4Gjbzys6eyYo4/vX2XHJC1xXSShgmzgeQRay4bGe6dnRm4sPWr1pngykrO0
NfTL/lrRLCDflm/BzEKA3+qQO2yO1TL587nKl2Lu+FUtaN1pg5R2h6ENNm101qUS
m7meV9ZkIuqg4KfIjDCRn+IIysllgNCO4ePzNDF7UMvQ70Qk400s2cHF+v3Rdoyq
nxUfHJ+fX4hvCxcTcFKKwIoeCpjWOvMc/P4fKhiU3efLEJxA0wG30Mj8aHgxeOVm
npVTN47qAl8Q1BE7gwOlnLdAospfXHxjhDDA/8UIXt4tziy48WADZMZVYUWkoS0e
Y6yjDukoxUgmDN0Wti+spJNsyG+SeVuLqK+hyMP8F5rQTbWKOEN7RaFG1rK0+TJD
u2UNzn4iG8LRpCnPIkK0GP6ylMUDt3zu+dU74f4dDWZL9FtVSlFDBsBnZttQkS76
03Oc/QVFZUTwr45OMN+qy1XfyAXmWvyPv4oXnKTIlgboklHlpavhdZ26pB3NGs7J
1BfQjtNdKZPfcHYViyc3NIuE/dYj8I9jB78XGM/ZfS6H64mxQTZoVzjztWnTTy03
kjx9SewWhiSP8xYmCbjr8J5be5Hx/YghjCUGHn8Nh1N6QR+LfgJC/FsyJgc0OJwz
yRVtXEhUWA1+zF6mn+MoLTHsmYNTG6Y4W5pIH89kt5nmvL51Tq/RrDfDrYyPlkj/
sViu/6Yq/wNj9W8kX39vtzVEgPDaNTtHZ6K9ZI4AeRzBHjjxTl9tqyUUMlyVqUZg
nTP0QTOBvEq4VwNiWNvKm+FmRh1VM2MEWx3NsW7e+HrBLEV8GtJq0e+oRP+W3i80
APUb8M7do6ZDs9WMvv/vmFzEh3qhsmJPQdIe5jx1CmgASk2LohfmFdEJySNFsaS0
v1DNt79QBLqNC3tdYRvo/ZEtI5R+hwtBfbPomrZXTQrY/Pv//uvzNoguGtHr/X3m
myC/+2DdYkzYU++ZEjIRcli/z4ziI/WarUmSuXyXubqM/FgBZbFIt4TvM+CBtCXG
VbdiCWsFIloenmnCvGYzw4U7ObQz6c1vBrFGG5WXoXJIdmOrYLZxxlOkidxOxR+J
uRsvne3L2MqH7QK7EWkSfLucOzitE6TI/jcLxPBwrVjZvd7gbA/Y4o5UAmMfdTdl
mL+O9gmTHRMkA2CbAtKf7A2YJF6W91lk7TYxSDNLAQgLpJkprIvYSuBCzGxIMwR8
pH/ZMDBFvJf5W3BBTZ7ZFPKtHzVSEmhlsyo7t527/4zHpl0Bi3wrkbcuWlhfmQJC
rXXuU51V+g4Cw2P+h2/aQeALmxKZMpXz3ec9/4tRwh8fexVGYTHyUCMzLLufBcGi
V/0qceQky9cs8s5jt+TRMcZ7qXN9ZQDpxu832bVeDw7J9K9/JLuKm7s31PyNVlxp
w8hZve9oqxWCCmOLSy+DqTQoriXSBphX7GbRoSmen7dN/CPds3tJ+gzN0UYp2Ghk
PPSot6b0mFOoFt/T6gvlEMNf6tQpxFbY80bmCCcLU4l7vT6QVtDNXri7mwKbjpbV
ybhpSUtTwjxtyEEaupgXTU2wwH6ovjPZe6/11R398xuzd4vuqwIvCkeEVVuof6e1
X5RLx16NX6fz5DYxVeysH1fjCDirK9LOYsilt6wABHgvxXuIV8cqwr+gduCsOkBE
1EoCQPLqvmRd7mvCvU+uMDQiKeAMbCc/O8fmf3voGQOFowtxj9X1ulIDN8X+93BB
mLxJogovdSyutrIMdQbDHW+Nk4i6ZsSs5lRUdobSvetY7BLU1A6u+32avRUii4Aq
3g8C8hH6V/LsomYkW+RAgZsBvW/GnyPxwZ2FD5bbiz2CtkssoAwMRiDS1ev3smNv
JPt3Ty7ASEPlTkP8Al0xT47h1/Y4IGQvUlUOAD9avBFD5GJFbgMrQXzHceb6y2tB
FT8hBu+S6mQ+fRulSQ5PdXtAzR1j2ioPl55QKGxEIcW6sL4rlzwmEn/0lEZsd8nF
6vFv0AmDFsiegYpz8iLeZdEBH4J9/6i2OpeVGNfv4f2vpJ8BZcve5sBLnIN8OPbl
IYDy+BzSddXmb92LnRaclqpIE/fiwi9wfz3sC2UaPqcCgGvffSXiWfh2WYpHhK3z
VpmkLpamnm7G9EBPs+Ld34WTebRn6REPqDOozJ63h2xQ/uz1mFEbFT4UEmNgbWan
58O7CbdrOIYS7zG8S9vgDtrEG5oTfFX5DmFIu0H9dedDN8cYVOeTuQswnTf+8oPL
agJ5HpDdHJpzRlK0aIzNtf323sZXo0Jof1UriLt8xdySZjjcjZg1FShD1/44rOm1
IaqHaw+Bql86ChfkCa5axk5A2RZOwsgepQYfszNEeqTwv8ti2u6Tjl06czEUTy0u
X7aghd8vGQLCdU44UMShaqxxjLeYDyu4y3Oy7Nk7pwd4kZo/W4cQFTFhMoveIcT0
KOgUCJ4nG2FmD+f8daBC4dVIrh2jeZKn0y5IFWIMx5WI2mAh3IP26W0fUk9YBdII
fUUd9n6/TFG5NNQqfNg/FIS+7VfBTG4aWjcDuKZdVJSc9TIcvjs0YXZtjW7V6hVS
hdGIe02VtK+VOnwIA7ihtVn5H1ptzDeoak4khRg2fq5tQi0veNe/e5xWPl9qPQ2l
7R2K772ltYFBhSyHiP5I4cks8aMvH17BtLEj3MGVr3jwQvdyJA9dVQyxtCq3SxoH
fIbHkHtvDpHK850WT85YFsbkbftbyL0WT0MRsih/RD5aKfjwUfJHRagl8RaAvebh
rbGB4DORcPaPRwIot5ezLJRChqsKu5HB7/boZqNZVbpHo4fvqJaN25+1aCKAWEpm
emx8FxbYiN4pel033KqrJ36yrm0td95xWppNMNHab7ItTLRUuZDfUGZVrLBAspNC
KYei+ViIxujs2eZpYwtcNUaWfDVWCcKfeBOETWUNz2qLZrhegWThTGOJm6px2H+D
f4UBI59qQxSjsNg+Tjlz3UeZSz7B1U/6VpCXIHS7CrwPInI+ZqIwvKypLj6E2qdn
8hD5Dm9SViyzDNk5573nHBknUizmlWQzFm5OtrcQD+K8IAInqdDLRAo53sPT+ohm
OQgxVHo6C02Ve3ZOGBSvDj570s0JEpAf5sdXSUXUPF1CauhXznQfDuPayv2poJj+
PM6i27Xp+wcliNyTIoKapUZOmNqj7ZiFspgd/CbUr/5VCH2Ts7kewEJK9Ilte782
Iydy4lh/d2gtSCqkhzkkmrJxQP/ZaLMzUcSvbVSiMsLbuLOKnTPnWpg/noWSCPGA
YdX1q7YY5+ULZGzWqahkTk1Xrq3ePNHmWUcH2/q0FZEAqMgb+wzK4HBjrCINQTzz
OtQeTtUXdsJtny/IoyNg85vUYQgFtZQbqqTaaS/eyCjhR1fy3EuBOFhQ/e++JZdZ
KnKFtABMkOCU5WPRPpLebF55FSc/3zuioWX5NBP/rkaZx5DH4l/g/7dPKSXsrvAT
OMsk6RqFRbUtxZmBMq0EntDyecCZY6Knefv6hH5v6QNiBsvRKXMSu390I/lv9HN8
plp+PsDRFxBI56YXHPPar1C0BLj0EaL3wl4vdIiGbHcT6l0c02Mh82SbNcXA2BVT
wgk3tycoi33mN4iaNtiLX49scYaPGS5oumzpqwqqL9dUsIGgIjENiEhbsDXtMFvX
yvwNDz9xu7k0k41WUSXRh8zNv1+qmJuygDSXEYTmMtoxXXlDmsCcJA9ItuN7rRrG
6hqiMAgiTwW1ZVsny5/d0yDhdcEwpVN7KpJB+TyG3f0XWMbOTWCrbF1IbVszoNs9
59M0phS53Gq1pFjP2+2zCI7C9TQYDXwiTeVaL+wArJdJ41VxdF9EzQP0icEzqlw3
rU2FnnanEkFwgAdPHVMcblbUntF7+wOGa+v/AVG233o+6h25C+elD2p0obEYx/EE
9mobgk0HgOwBhxaKx2QaRVKGNzQ1an4dBsnvQxN0Rexa7MTjMwphDIkNepZMZism
x1xUyYHw0YFJyZLMecHode6FV7FhXgxQeudZzWBvJ5c4odSz0cwAVdFQ1RXBmYK6
fZ5+qKD3aGwfoVALICOiKUlyFQXzK3IlRA9i4mhTfrHt8f/00iyhoz6XsS+Ifcaa
3UD/WcVVziLtQdABz5fJU43El7ZBShcHmFQAsWw9VbQZE0p6LTEgbWZ842OGRinr
mPFHwBk6ZggmB/GMgLVgtH25MzusRW8AVYng0iog3Xn5m4wJutJnYIjNIo2sFsRK
X6/bH2KReN0drZ5qjuabbdzWULRYfDJmR5qqGeTTh6Qb7I4o/ah2v97QUpnPvZDE
3Kyn6nHb0Dn4Pki9MI4PdrV7NR7WFMxLjxz9HYq2qSi0vOeXkRjODNXSh11KlBGJ
W0wzcAPyDeGOxbcr6k+Zflzi7LU2gKQF3qsIXQGMYpmhOqZ4eRi5U973G1ynB/2I
zWeoG2vy3RjgRdnxb+w7C4DcWwJn9K+C8tMS8LggiVpQrLzhMMHF9SCoMRi/icJD
R9CYsgEjiqlzKQZl5Hp5rF4Fe4LSfIE9ZKJHFKozwOg+ItLV84/BZoH4MFaOSRDZ
lf7ZtEF5eIxTufMeC10rfN/ZHocZMPoyyNVIlkmobKdqFmkzr7C4iLRXNfvMcH+C
+Y99wb8gdncRgqDoga/yrIwGr0kWHTX6bkhc/X1GerAgAOfe0KokAHrpU6/jN1ch
6qbaW55JwE2QtPTSECzVUPSZ1ho4UGZz0mXjPr0LyTbJ17/NDpCSqguKUpPnj0Kp
WSqSk8wfBEtvBXiM4gNBp1mKs4lmtSzdntez5i3g4OFtLP+E1iKIhpPi4vzjJzzu
eU3mUIYwb8JHnAbHf4X6quZhi4/Qm00dxgnu6RlCkBef51GxoXPi2iHND962Bgbl
Sx9bLnmzZ4BUj3W+IWzNBrtwKhoqUwh6O/OqB4GG3JIRUXfhG4voI+1fiCJiJ5Ck
ed5aDIhiwqJLmxCZoPkCx7sFjn64ffbsFb0jYuaKHJsOXhJUX0jR5crc1zq1jCTz
cru9BS7aIMzSwh3dP6+0bgrepIdpTNBSufsvWxd5v+H6t7EC2bU0QE+BNqhbrV29
Ur7pcPMxjzTLMBxj6RvH1Wp80wVXekK+Ow4nulXUuBltkrJDotNEiSdxAi5QiZ4R
Nb7KA0FKW2x2jNrcVrbzO4U4J9OZ5XmpRF+2xNVpayhg69nJIKmpGwv+vh2wOwze
cJ+ezjc1SS8DzI6EwPYbVGLpfXj49/Lit0FI5EwOMe/BoKxIMBIoDhF2CrMYA3we
nC4hJw3vTngmUNeTQzeZ1dk4VnDMEvAEWancD7Hj5jfW7yoww0dgsPQATv1C4iWm
aQusLtDxOlArB8dawxbQcLG27rAkP5Nnx9Pn17yrvzpaOeV54qEc0VupTWBsMGpW
W7bAX+BBqI58FNt36K1pq/OKK7GiD0BlX8gwdbA9pWgfK8om/TYMiGbdSS/HNeTo
cDYhXtr6bp3M2BM2xGVZWGLC3RIVBJFNMtbwcZAj2elXkBC3MEQ1y1Ig1nIs3NeM
HYPh3sviZrHkUegmgtwrKDbNEcAbjl0krc73jBoaRU8rbcwIfZYvbNGGeTHjA0tT
+F31shkHMBNAZ8YwCvl6qEA2c0BFVWhDfe89dJKPM02q3z7wb9JhyaVVyku/1UPo
lmSADgrzwMEDikpBx5WcCAN71K9Il6dA5M+qEg3McDoC1aC/hlNcDfbAVTuDAHgb
yG5E8mOyOJga1dUWjdaA9XR4VVls0FAcc38bSmO4X0F6bcnpinkTmfehqUlBdARc
OEk+5dKQBZKl/qhy2pGWpJUSAcNKnFL8WTKmbo3XlII0en8gFwdVCZszymTR7zF3
OnmTA6sq71l5oye6fOKI/s1+Szg4J5GPCHocQ7wYQHf1Ras1WZxrD2NWFIRGj3Qv
nfOZNSMMevGonBYDwvQLuhpCg9be52YISFaVngvCeEw4HOROjiSCPAymzgbnwyv4
9Q4bGDJWK4Kvw5MvQH76C9pVdt534ve5YxGxPGFWN1HtugTNPL4eIdNWzVbjNijX
ZaUoYxvducbtv6qiCIlAqy2AejeMdHzwa7lKTbOzQufUpNo1Rg+LMd6ctJ54Rfo4
VqyApAFO5+LCOB1otu0azJ31VDZQW/EDjQqkOGj7P0IJ7hPukL3M3H36bKiPxKlB
4AzFy2S+1/q1p7D34SbL5v66rIXwVN9vO0WWYoITtBu6KOV9WfU4n2NK+rwGpHiQ
V5SRrL6Q1sOcn27LysjyMWjF13hg5iqXQBNI/+gOzbqyiZh1TTQJn+WIIu8Awtpu
Skknu/C/ZRdFTPVV/Ix0JTwM8ke22VbW+RDB/9J9AvWBSu0wqwgQk/AbN1EO4L9/
rkkHt/XjUm3fVnAdTqzQ6WaipTuO8y4v7V/D+kbV52iMeFUEV/CVd2EcHAjNKcEr
QcffS1re3goLFKi/xDamDsdS0axg15SP9In4U/EquJQdv/0nSLZ5kTQKu+/TwPdM
jPKvSWeRmfhtPx2mFYpHIQsOD0Fq5APZ/PP0YvBTnXfDd+NMrToo2EaNEqxTRaZK
KaRlEou/UW4mpcHSXnMUC9TNzCsLgWJ4Owkp04IVrHmp42Lj6NaJj03J1fA5uROV
V8NqubSMq6YvQ73S2Pf4iF5VgW6ZUrUS6a0ZFSKzVegwpi9IbMVt9hGXHqA17+X7
tqllEiRv1rfMyTw7aDrxAjUI6LIcvfN9h6xlhhUzq1qVLR6K50VEbMMlYNKKmHju
5byf9NFHIkX+yXq57fdt4WWw2MetR7S2Drk6Ft3oLKphCOtMPCWGYOXRMG8sUdLI
0BTl4OXHk23QSq52aHXAcVtiQdQqvRjLrRAAn1ysITqS3KRZtEDvL6psNKaC6IEn
YJR9XBllS0WqlqbA4GPLifKozLTTnCHWEhh7LKiUYpj2ljnZs8xZdqPMyEm79Ngo
eB81DEybz7LVoRR0Q6EIho1yUtfHu9eZ4X2eNKhFz2hEmtKaHr6009n0oDBlk8Hv
J+UGuz9ec1oFn7USQe4/5zBq3ziVmDJWCyvJhaDt+tWoe5Txy746zV+Ow8r0cSnB
fPI2nqoHXyeQ4hqqpnrU1EWLHX0wfTSCGK4+wknL4jimNgG+ZNggl/i4lOXEEGWk
J+3pe95IvYBOfEiGzCE9INfFnojO2xz9MhTQarWFfyrZd6090qhEqWPhADykzL14
/KoVYlKPyODbHoQxvGQvC+jk5BNcTbLj3uYt6p7uBsYA5M8RCQY8uO/dKe0pwkM/
5rMd/3W1at7KYFL6saZJWm46WEqNBDXzhnEgSI04RujhvqmD+wM2vCzGc3iXmFyr
EfCPapibFrVnRu6kJ/nNSpLQ5m8KC7PKL9zZI39A9VaKqR/lkoJ+//y+SqtetzEf
8FaUTA9wFKp+JKJoUKMm13VfSAliRxQyG4WNUuIshLmid5utIrroxztw6FpVQQOM
/GOFleqk0hO7ZzpvofOMSRlRwlPUpjQBRIfEJyrHx2YRH/DRHf2vdUCZeHNG8R48
J7N7uhhcLRPHZFQ7sx/X1p8WgLRkKzdERPdWEJkxYyBJTcG0t4aLughjeSk4wzgs
YNMw+P8yRQ7OlcD1n009jf0ZM0ZF+cEyGhl7hgQC4SI9jwYdZEVkXMbb12l0jR+Y
t2lzmp3jojMQ8LyDP7JwPJPws8EJdcvB2WJm3/omouFG8ICZKJxfvvukvGFTsULr
oAK1R77/z/M53rSwbvkRhDaiEQMWBgh+X2AX1buiPyXHR8qI3WwoW6a5szRlqY7p
zgqqVNgNLrXs9F8oS0b3M5M87RzR5Z6b7MY7YbcolYNbH052Yg7tstkBx9jj+ZTT
EbDGKotO/tc2JxuV3MictS4ttvbBPeScO6JcAa8fTCEI82h6jhHXO+ZZqA7sTb4N
C6boTVMpahbiljKVPjxdMnu7XXr5phDi/1NFWhgRnjBwMTBAO6QmNWwtB9kFY62B
GkAxoL3HTdPsh1p3JReZtOhTQkz7YgchcLusIkPa7trvwvgtBQBePfigLBUzZo2D
ygIfRELmVgItWhGO8TelaDn/cqVZB2xUGmflPIxWKMup7ORHwzMAgXMbEtGkoWKn
gqfH+Ocfok/V92ccurW/lFLjKBND+Ms5tZ8T2M6I8hqW/nayIW8tbj7NeXDitaS6
OoXbo42Z2OPQQHVRWIQGLlphW7VeM99WY4yxNvuyqowyZ0yJ4mLs4QxWiFgOZt7W
6dqOS43OXIJG4XuoLcW3J2WnNnpldTLzZwBe0Q7IZG9DN8zcqqnnfJvv9v+MLB8o
drH01dVUZR8ZsBD0i1jgTsWk5ih8uDoGMcNUr7WREUuMX0xZg2Unykybd4fRQkHG
3ffQvdWuxxEOe1++5/LdjB9oKONogEF5SCxBg7VQqVASvOybq19KKwin+dLlDb3u
HKaMz2fS8d7KC8qaar5vqqIyTCFlo6tRPyPAoU8a5+IQ3/AfunWRLyJkf5/M+R1A
iJ7oYFkiL3/JYzj5sYaHmyQQpOK+wqWV0y5jxEE/CZk4aqu+gab1rS6IRjCEy+7o
MkPwAlhNeHJRQ+VhwhH8et2L7o1FIWHx+90XnQJB7KLLx7BeF4LsRA0I/wod2Vcn
FKOFxrrOlHEEUtjTF0g110pnMi5ROrHB81H9281ry4+RypLdZbJDTruOz6QhQyyg
hA8RmgnTFFPDO2raTskUuwhQ/0vyuKjyN1rq+ApvDuk6l+NhgwX9EFlumtsvwgJA
cHfgSOYtbq/t/VbZk5vau0MxhzFz/qR8o6iY6/Tj0Uu4PsrbP7Gff4ao3skWLuSx
zZS9BDylYoBuoZAQP4dUi2D9a8WgGmJPC4l2rYLRym5jm4Hht8OgmA1jDTfJqPbG
FNR0mw6lJb4jFNg/z8RC+zX4J0wUAOMfYk3jD07g7KAefHtTDsCSyPjm+Qj0bozM
GmHejV9O11WsLjUM7VIDpvIKQDMktvhfAjgl0K6A3EeFsrJOUGF1rCvWx6q45Rl0
35IIPSbXO/l8cejLlcyIwrtmUF9/lrWwBUGcf3HPcwVaV7PBF5Ar94TfrwT2sWoh
8sXJFKBtOpIrSEf+9vyYx/Vz0t93KnR+DmuJEH1YdY/6uh0FFlejub0Cs4u5HQiL
MgFR09egO6JEqQlFHO1PjZBVUO3cSgx/+zjYDn0kGRVU7tR+VXaghvV5gMJ9+hln
30XV8pb6ggiQWvyy4mNAf2r/hiaBBBHrc1GqykXcYAj9RXWITbAMHef84565PU7w
O+VUR4JBU1opEEL2egnwVRKZwAx5GcnLXT0eFD+TamhUrJVGyFqnTVCn1Zrc96tE
9R5enWX6ezMUcxf2Io7KdaJUVq3wOziv5A8DlFOUaqs/ksR1JWveFw6mX7uJKt4I
cBn4C9JMhuNQwJP8jlTZmy/kbxrHw0mipZV9BXkOoJ0enq6yxeXydAFhc7gTiJlQ
qBv9XKViDJApEwoh2DTl1oso6y2pxgiurCYJi1/SARxMrdlUNEH5+JyhWfDZKSoR
mkxCA6e6vXLU6rvp3QDL9qJMsc5H3cTkHpX/wieUZRBEry8wO8E0Nx4Ffi5dcb2T
HNdCW41zU2kQYMxTdRc8N4ZAik2AdxnqD7vn0H5TUO2qqVYHpp7gWFD+1Xt5gNpc
kMJnNIdPRkMjvXIhOqGVmxa8iVZJg5wXBZwJpcHOJ3SAzzM3lpoqzsk9T13cvrKI
Mzs17Ki25SuAn/Oqtk2VN1Ll8gF7mQUXTwoFVIxdf9qUrT0+uWt1lsHQZfqdDveC
nDazqI1UCvDrRQPxbWD+8UXhNXbQyL2cAnVlAohPl7wZRL6ZB+eCEYNJjxHZiWKq
tDWjy7TOSMGzi4cOdrEvB5sq0FfjbTHl7UxVK3zNCv2646r3Zc0nKTb04M0fEyyz
XVs7hgtpgyVqkvF/zdiabgsV1l/aKo/QCb0ZMo4fXnNv20tYk/zPckPuirDSsygw
XsmKHHyYmCgJ8JCJHPIiAdq01mbUB1em+YB7U7AYe+RkwFojme7cnIGxX7jTPLVF
jtICctTNIHG17Np5+6SJk/6yKmqNBfFW5uZ/z2mhF3rhTTJy53qPvXd3quS7ysZj
hMaESfRkUet3xHTt8dhyrFAq7+KDfUdh0JkvI7B1B6hX1wQ43WwFcw1y6IGNTLXZ
OwbZ0yal/MczJKRn34ARNvh+v4aSuyJ5Qdk7H/scIDEEs/1eJ1eYJZJUhQHKj2p6
9bWJTTCjBes5lsf3m6Ngj15n4PR5BAvvi5FgFVP9uMICaXOT7kTKl7z1OtSqnZyQ
Netg7gvNPfBXTLv3GzibK0EhKG13q7Kt1ZHZoRUWU6AOZWS9bYgXaJHLQqaTnuRp
DTfbhIJARGGVfNXn4GGLZ7xm9cb+cqRgOwkvr0yS7y13YGBOZCMhWnPXuIEC9HD0
a/INkCFwz0rce69ihKxs9x38HnJzXMhYCoQDW8+jd+XPYbl7Z3hsXrrpyYO3cnh8
K+CbEKuJt3nWDGTy7ZnmgdzdlingwcuQ6cALQv0fFycgQ43CqMrEp7DyCfuaDijv
HTlE5uu7uOkswnI8IogyMvmAk2MyS4mkA+s/BCS7mhCJijyzjVyts4Gtd0NJUhCa
UMqiBHUl9zIMS8oz1S6PlzW9hFpV/zSUp5WrJk2mG4C/tnN5zjcAzasb1iVY+H+8
Sxi9CkZQJRCMi/N4I//iTUAQr/FqrZqOhSoNK+245AdInBSz/A13GkBHi8PeJlnd
ZEKnrPVEiI0dF/cEHEJVrn2PwGiztXmzwRVbKDf/eLTY6c2ZsnkOviy00CfDapw9
0godrdNFKEj4Za9d6SmBHNmcnHL8A3/jQsw5By+tzE00uohy6HVM6Ta91UPRdYGR
/wpQjlWPcW/ihkQzfqhMZgtciTFBKCBRAOeCGnOpt4PQB8AetqThT9Uuoc7/xkrk
1YhByDI1r+6W75cOxvD9r4QA58qb0se1XpT+JjeTUwr2X945NzLYnvGiRD3MvxpQ
TsSD32f0HfQ7VylcvoFrkDwYIDhvb04uLuhY8SvdX2QgWFD/9f2nt9di8+HlnZGW
hju64R43saCoh05S6fjfREX9/6Lhx3bDGhTKaO5SXOFsYfTswJE6eEwKv7ONvvql
OYUBTR7l5k6gGi6SrmxCT8+s5w+hFpIXDLwei4aWpeUsuS6jdsnDCRbalmYt7DZ2
S5wsBGkru9gjlFBnVecjAcgQaq1aVXW9/nMC8w+C3dRp9CqUo/rijb0UwombEiY+
MpxQZJZ53X8Cz3rsNOa22t3yM60LVi7gnJNtiGdAQqQtwZEXBBK8enTV5lEDs2OI
clS2adPb/HmaxMyQ7rozA2v8RNPMJXb7p2lkWa7St2cz+3kw5HuCf0uB9Z/nPRCg
ZzJGG213/4KrRRb0iZgKXCCiAzkKdg1TFHNFFeP401KkEtZSpZYsmMt1i06VXdU7
EqutLxtkKXJP3fNKNyXBgKyY9EMlTWd6MGf/cUOWrbWOWwUmdAbvnWWdLtlPex1i
oJ8YBB4EsrnjJEH9jn+pnw0SjsJDGuecyPb9srvZM/emb0qbm9drZB9tTx2s1/Or
AtgcSagN4p4yTpILTHB/hBN76uk0AQXbsvd2tRCEnrVvVQ2c5rF8EBmNZiyBsJ0p
4IvDptuKJQzSiFWxOEflhvbB9jAobMqGajqDV8bzuOj+x0HmjNZ81oTxaKK7EiUX
qqz9yK5tyZ+8HQQETV3CcmqmOd9dU59oHgkRe4xNKwQ2tFXhhJr2NKiGCHDfVe1C
oo/78KqtNn/xNwQ9y/vNI5HjuUdIrcFP+rQ0rYaEaxK6Cy5o6A18xS6wx5Yg4DVK
txQUVxjr21u3ZFBkKfQeTk9ekR57HFI+MEqxImUSWO7PR9yKbyE9C0immIN3i6/T
UFGp2/W/w93I8rARKa1XzPCk9n7pXRL4LnwxNn8+lH+VS8axo6K7f3AWpgC7GlOz
inLRjkUYkoURnneC0tiH68H12m5z2WS6yGbqIngsx05+IrX0XBiTUtUaC0Ua6Mc8
td+wVSrCVIHoC2V3jnBZb30VJL4otD+jc6NDucHrdW58OBHpJBHCQd1jWpT50aGk
darBudOYyOGZx1a/3tbPAIbqBA4xBANXaDAhJYN/ApFvH8yzRR7dNrJVzY7LyJie
BcBIC/A+9xXIbEHgt6VfA0rAl0g5+BhMFfL52zHaFshMwf37RJSUSEOI2LHwRfsH
f+F+48IOHo8g4fyik23e45kPeR8/9a3DD/vs592SN9TvmQ7OUGxPeAsCtikNw8eD
sIXGYVTV9KtQAjJGuB8ctYr0Iu7klCSoxZt8J3InbilBMh93cPrTlKcOPqbF3k4y
voZJ1AenJ3o5BaYWDiOtdb1E/49zspeeT/ysOHul10jalHHu8cOXZZO2/Qw07uIs
ZeJJf5wgK4GjFbtouh0c+KrDRRlcNhg7zWaXx8AgtknLhKpQ183QUBFboXXFdJdJ
4AI+cOK4r8iTeHKhUXhUXepbuzgUZkinkPL+2vP9z2V0iWSOC1lf68/WYUlLW0dE
d/fNVkWHi3LWCDLLbz2yeMX0pSRuYKxAEchgeaBj5hIJ292fcGgXxPjH8xCPYuz5
N791r4bbn9RVaDKggk2Jxu7tnmKZq8dBbHP14Dfv8DvpAI8v8/nR0LID115xk1DP
hgzWPxrIrcOFfn69QsN7eQznuqu5DyqbGdqGIObqOdo59ZuX5Pn9113oFFfV8Yy6
zflUFVdimDlMq+DO7HbDU0AYsPlSiEgHziTcUHJVPi9/YPMlxgd06HI2O1QV3OFx
2tMmm0I/2pXmzVIHlYl1rIkDU5ZTtHcuSGRtwpXC4Rlc/3++vgAur6CFnsHkL3xK
kssB8AlqEDAYXOeYoIgCXLzqONLOE+PJnKGXEqCEX9uVCyjCa51wwaDGlqU+wxyl
TjS5QTcZcffCWfqlJ6j8nR7SgAJK2/HCtxc/Ajrm2/Gumzc074yUGqIQgfA9QX0S
PyxyyPbUttJOMsSTzFylIF56JjnsCfNE86rq7//gkAYdiO/rlg/ShxU7QdeCk8OL
fGfpbagBsXN6GMQb9GllMyGkrZjsmXbhVjylZvScyp0qcafjb+o5q58d5Vpb3Vv2
MmDeQJToaB6+ikWuEJDIeltDNB15BGnwwqLbrNOLZcB+XlNRe+v3bec8Q3md4lh7
tXopieAEz+kzD3+Txtvryfy7Tu91VtltBEZOLvirOI9BJBwfns9PbgixhPG67gcz
/V2cZk7lrnqh//ufeQI9qjCSTCQjWR4cdozawBg7nweu4yA/np3on2PbfempC153
uryXjv1oI589TVUPDcAgJLoRwpWDcY/ooWiplytbjZw36HewT+dMyiZ1JVeZctgy
zEXsIDPhaPgLrDQOAgzLVna57YPshr3rOIn35SWSoqFOyc115P/ArHk8wynuXkkd
fJBhSYRtV4CWvgCRHhANYHPNtvo0831YMz3FDWPoVL+yMWez1us8wRCVEj6UJQAl
WT366a6HTDR531dp8g6UunCjR3HZaFR3eK4xMdwqqWfJAL5DQNqMRf7twPTRAN/w
aWW5EwVwnUDaWjkbph9TB7g6h/9KPXDCjwMcwrciGgpo4m7WpkUahjIZGCm6ZnpQ
pVPulkIlLZGAg1vWthiw6TmNBqXlNCDaj9Pu2RDp2wgH3MRyHpICXe8cuPbrJ+kI
ET1LndvaiHJd/r1M3kG+rgsncz2jjqwpnRsd5RrOWFZhTvDEUiQhagF7SKb5ovTA
mvey9nuxoNMVY6WAwpeTLJsHaeJxygIeW/0TlMCWdFmWS3rMkx9JwHNgXE9UZ7Tz
kyids608tJiV7Zd0Gz5hKff+scrt71e8ufovzvkJe1LaHxrHhZIpQie0Dh85ogak
3B6Uzzx0JE/XE/iQf/P4gsiML6QhVskFApoSmNz59kBzDoPTzMb7NktRJBVKJbOv
to9MOt77VdVKFkf6hT2ZJOoTmwSzdrcuuT14mHH499xRW/fmVAOyJfT8T7s8lg5L
/sNBn8GM/u49pl+T7imlUzuKg5/oiCbpUavK+bwxEhuMjoKN1f/7gm1rFehUYYCa
CPtWaADl/Yn45z2Chu685eNUGJ79sSE6NPwUYfOnR3z6++EYpYf+cBzb0s/BATqs
sr4/f9ScQyxjl8fBNSErJrxAlCHs0qHSR8JdflyMnlzZ6jnYF4RepOJObFDJClAL
DQfMOWxWhoC2BxdMktWOyEAXkXfqHZ9gLNb3VGHq8s8QOT1Q9fQnDA9aCDkAA4UE
zC1EOUeq1yWYTRjz/wPQicDkxjwBl5Nd9QWPLxswdHUyCCHiEu4lllCIbouGs9JO
HRjPTo2MsMSCC5llDqtlrbAJkETIBDt1Th4PR8a8dQj5E5SamG/qR9g0gjxHT189
4AiVd4Gpu11OSpLod3aF7NnbtqQBNjGYPrEplAerLw153VUY+tWMpVC1KFSHssOY
Bjhv/Eed0kzcvM8onpWL1y5N660ehzecrGoLyNkzFmXZSyzPm9t2fNHljsd8qT2j
XMPgs4fvUGf//CeqZLf7LCgsWnB7VCoPRy97tifU1XdcGrMAxCT1HttQkA+6N0Th
1thKtMgAkF3dODnc7Zlx4knU/1ZWa8H6mBvPk7OTNYqdbvXdD1LSb7516gVaFGWJ
92B9XylhCsZCmE53ZmPiMiMj+R7ZUbabB42j+cwlW6bBmLiTOaeurddXS5bxUgww
0u2L2BXeczN54mzJERpqfIOby7fXt949ebqWWjVIWx1IsD5UUlKRHuUhWXZPLdpk
oABzKLhU2yOAMTNKwT5zYp/5t6LvW9m5NCbUEeo4qZicZf/hjbeqBSg4cW8gGvXO
HWDhRBC+ULpK5oEcq0xXBqaYNeH4PmwZN7tekHXiTd1sGxoZy/eo0f9WFHFucgU0
g9fHP/sLz7+XwxNHT/dUrMArdAx6haJG5YCgP8vNsOJQPV+Y2hS/JbHYq3AadX10
axxIYY2h5D0J0vG+1qvItGHiSTN0DF3OaD8wIwh8Xc9TmRzQx74+jnFUAbdQXEyh
uIc1/3swbK9Hy6yxzq2gaOUFZlrIyto7HfAFXNIHW+lJvzRoZk8+jl1gWFX3ycXn
P4cK9l/dNqFmzzQZYYmsbTQ4Atxj7dHY0VdaN2rED8JVdrFe5D4vtHqbWp8Un+5R
hrKHxUn4l7mxZROOohQyAAevlObOS/lGigpiyU+lcxrOJJMAPriNz01Yf6kQQbRr
m7nzDBSAw3mIADG6SHp9Z0MqKzQ3nmYrEm8p0PZYoC7wyulUmrAMONn9HYeJihLo
Cffcb22VidXkqEYlVtYWRQHk2Crw9ODJDJSsSF3CQxsZDO4Kku7GNM0Oygg2w17L
EyOILTP59kJCBJqjnqWdunihTNmRfytsSFOjFWmwg0iGKLThLRrjXosU/x0U0SZj
0HraEg+LRMlvlrnzzzydna3NyzFk/pQp+tAnB8CY0eBztd1wxxpy4MKlB4ngEYTQ
Gqn5LkydVv9LrKUCFyVJQ//c+vcpuzW3ue628JZq6pLtlUdN3pKME+48+yoxYJY4
LBIrbvOTlT/XQlkk3vNEmZLYgLGJDJg09HeteX83bLKR1AS2t6KckaHFEbNsOzzt
ipo5I/boZ+zADbQTGmXfMMF5y7EKbLuyQ0dMydzoxQP9TNiAG0GI7M1EAwYh3mnt
1bvNTGK2XpPbW413IEMNgBKMnIDJKSVKdL1bdlzOMqR2SN/R/jZeJ3j8mRaiQV9c
WoqBw9Z/+a7/jjQjKTGF2eOy01x7l1edflv3qkb2x0N01dLWb8VyHuxz/DUUtOx3
Px201Ihn+6UVbX6lJxczhvUQtKPwZqDAcPwCbioNcNo7srh6uxv/7qVNTOXel9v/
OZmBSRRVlHPK/nOkWrdBitLY51R7YXKmjHTQvE9dJoLKbSBX4RfH+KipW4Ryr6gW
KMNUvL5wwGK1vYk6jGDHrd8PB7PcQGIMTBtc6rGw1UiJm6FO9L/LFTJCEm6cjqWh
VMVAWNSI2A5l/wToZ+mGRWzqintuXptPzcDZQ1cci8UDbla22uo0Ccy7J0R31sNJ
4aAkw/mu2W0GUmC6i5Nbv++o5h6Oxqn2Yz6aZYWU/hkz9tr/XWzDJn9wkPLqHXoo
mpM/xWQ4zzYBvBLdcRdgtfpsmgktpoF5Tu9CokipYKzjTo9eASiERqwvHsS3su9H
lAfswVpu5agcbnkFHl4br2+85Yph8eDmkQPH62DQBF3hvkqk2Ai83Y3mTwCGCoux
AsCtEzRU3HzWCGAuUagjJ5uLCCp91bxm07/La4UK+75JXASzvQkXJeyr0+qbEg/c
x0j1N4zqP7oCoeF9YzdW+cBuxDAOFt1Exxtt8IKXn2Tn4FNCEJnEV+AuA0Qek33U
MCMEgmr3+kGJu7RQJ+SH4AmMe3GCydCgjjMSMY+XpS0qomtw2zEHWL/KN2L1x7uK
aMknnYM27zvfILROobYscaAwXDW8mQwv0kvcGGCD2z1zbi0hp0tI18zyo+YXqkDy
rkERZkIsrywHvkhv4GkDM2MUzPNPS9SwF1BSOHmj0v3dSi++fNOrQUrIEHDcOESd
aq49hKwiraAFOyLWAkoLRNROA84+0JtrKzPaE8CZImIYM1hnPoi4gXO4zjOSyT/B
zn/7gYPmD0t1kre4l1uztQn7+vBiOrLwm7tINqenK3JZl12ucdCx4DaGztw2XG4w
n0NqNWFv7CQ6UmUKNhy7jE34mPvvLGAMltS8kowNMke2P4Uv6kGdvNGU4JCVuDb9
mlFwiFpu8loYff8V4v7/HjW0fZwoB1+WXtBZpjaz0I1hyYH45Bm8wQnlr2Mvm3de
C2dT8FM7ZWegwwRZtYZIMU1UazBMSyiEMDHy9eSGLBkWV1p1NgQzrmgr23jHU5S6
LrpXsH35lsTJBCM/66LOOL9t/cRyZuUHR/65DoMvtrEIY8si841Z4KcewxW9IR5w
2fu4io/C7PYdm7Ch0XcFq9RQoNyVYqbnAmakZg80wvRNrg883Q73UPQt3IMwKhOx
UORDM6CXUxK25neNmttZxyzqEhUNeTMpO7CMuFmExd6X1086tnSIrcRRcPH/P055
KgVBAqIVTrnuYI+9dY5iTdELOyirULAV20AhRZ+5r9b8UCtuIaaxPol/nUhyl/R0
TSUsjuZZCwjpOquXP9athTRONX9Sm5tnamDxzDFJf+2fRVyga3oJquy/3OXokloE
o3DskHHZR4UtEb+JhE419tJP2K86eSrX0hYV1wSps7xKlpGW5sjGpNJ36HUzOrwD
qInTA9MpHvq2q6UNS7Wn/QYY8eDvDnGx/J2QDhUke32fE7jV/lJIUOlNNffJpGaq
6f+pP5V/q7KvSF9+9HlKtXFfMrfq7C08oKZ1eFyKr5HbBz4vZjT2Dp0L+IKWPmsC
iiEdpBjtqyXVTEUjHpCrBm6dN4NsuMxFPXWO7v837DsXr02aMcOBuZg0V7j4xWsx
gvzqVF4fvv2DvbFr4gp3MWWj9+e96iS04alojrNi/f4FMgC8B7thNIcpnQXZrFKs
Rn1lYBVG2ALCs7Mb0Pk05fK9s8/GvUIdrpcuxeYnAUrf27pPzr6XrQhBU7YhaeuM
EgndOicgmvYFPFxP76cggYD7zYmsN7U9LIiL238l8jidpOEWuoMDO73UzwJNUoi9
paOp3Z575H6l/+w46CxZ7rCnr2IiEoZG0JKYkkCzlTxqgsQWzSuw443+1jwiUYB6
`pragma protect end_protected
