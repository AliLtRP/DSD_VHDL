// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g4i2JVdE14SpyWyU9OMKGG33euTrNiGxOUNq2UBs/VUQeayOjOPty2oBxYubt/BE
5mox/2gaAkTOCynOiLGASA4xAdbbz7VrvBVdak0nfy/bMBAZvNKLBSgGprCMO0e4
aKfSOic15VOODq5qcorAYCi666gx7CEe9+aHayVHnTk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23504)
XZqV//uk1m5Ry8OYiYAbhNL9eE+RsWBcWuDJjwoPlf75hqOWA9N8x/qItZKIxJ3R
WT+qOsuN7LALvV7+2uMJPeXcg9wnxNYmncJnEJ87YndKo8UXfPHnovgcbqRZI9db
ltAnq7KagxFZWgaA2I1rcvbsz9Xkc6VDk8DNjkiKNpDt/6j65v2z5ujho1PijU7Z
Q9GUpeG+ReYQS/bYJK0vLWrObU8covWuIYXzjoXhu3Q7pMa/FjBv4mcjRxr0RQnF
DVHjX47GzSjGTRwpDI/IoWbKcDSDdla2TpdEfdwREIwqv6teY7PjJDrX4F5hUu9J
gvyAnd0+cxkdnn2KJSLE+nmPWz+wiwRG9BJaEMPl08Hpu53w9SLV6KRI+IgI+mqO
K+9GrHzZwIBQtj8P0Sge1SAiYD0HNUSFYXWGnpwaG8L7UuVsUg87+rxetd3k3mlG
Km0+NMHO13e2q+WL2V/ExKwRaGbXDdTp5/OHKrF69eZ/t9uqkUOAuL8sh0a4YD1A
I2ETyf5GVpeeRK0c/KGDksPEYoaDyBi5ndUGMaC5beccC91PdX/klHrf8i37N1Xx
kFDWBtr5AjxloovvJug9tv/y7avswoA5uqC+mzvw6a/4EYCrvVqbjMnGNjYRPM5l
tKqJ6GQu2DmFQtUpc5KeV14kjqHASd7Sr0i/TmzEZ5lB3f4z3ulgZbrTVT/PWkcU
ZWSwdLPwgWfZFznhhbqeL3+MJltokmsMadNmfwgS4O8xc87NNF0yaSje93Q4JVE6
gqQjtuJe3zhPd+E3A9APVxiGv7mftHaM3JHWgDkIyzB7rMyDJWJWWdmdfvDmMB5Q
qFpAjrlLJ5uJLBBkIjziBj4/n4orgWFDIlbQgeDgxt2Vu585anwmEaTp60ZE3Z80
SRAESpjiEcEgzAvVn+n0UntOPIrtkXhs6xkIhhAeOWkx2LLO9ba+c5JI5ngYuGO/
CZlnB64bv7dDKXgdOLgnFWeRFxsErJxysWlGTUJEPvBVdVhYZNUMMuW1N8WkRPXu
0DQ67+OKbY08+cu+E/4o+ekvIwDpEos2tRBhwseki6bwH9hAWaYaOQHEAllE0fpP
L4P+wzC9Vvv50ADPtaCx3DXg/jM1Fd6nKBnyPOJY5VzWEu4admt9pzG2qhC/OCcd
HCLBpkS4zNdEVqPo4ACnG0wuLNK0klqx0nAWAK93B/crxNhFwkUzgmHbPMhNrtu2
dlmzYq0nHvycLfQOZ5R1+/YqneU4GOuroGDpMEE1jo+i9TahXiDiyiDDWPnZAK+C
MEoVO2CoDbY0/XmhVwS74Vzh8jhJKsSOjzCMl95psEFZVoK6GWuTf47P4BLyjYG/
fd4NZQzP+KB0OP0iedzvKg0QQkpx3KDxgj7QetVYhcwa0cG+U1x/px9nue5KW5RW
2CRUtBvsu9Ciy6Ie/9Fdt49jSTRGshGw7gLyand3ZW6pC5Z1b4dXNQzi2bkbn0az
kHxYDCcTVpprtqf8/qeW2GQSMEyaQDX2jcqlPQifOTIFRMs7cuvtlEdUIqM5xoaD
gsUt4H/EouRFNAkwKG4B2yNMTdtxVyQNowmHS7K2sJwo0cQVxhJPW6fDPPn2HfGJ
SVu0IVasyc+kZio/prP1ipVfHedV4edrmRlCDisOmgdkwGR+t5I5Vtatwn+wgAAO
nSON+wO04df+o/SNJehn2036SNMwtDuG9St9dHzNKze1sIDh8lLgUQc5Td6hc7te
PeKYK5BYEHaiyB6Lv/eL7J/RQmiirKY5VT0mTK/f0A2Q4oscYSlq1tRVuPG3UHEF
18GIcXsfHtwfQKSEvqYy/qUOx4tx92pRz8lN5XdYX0MfdrfBLqXLJMb5gCL0cnaF
9r+yptH501y0Mn+j13GMFSEfSc1fXvChRuKnTLYB5wob2uYg8nGD8xzgEMk56+m/
4dwvuGIh2V4XkoxmL4jbWDkBL/c/FpnTLyiFMMz2frQPlUqkRepKdLZIBQzlGgCH
ASUBvSyn+K363AmH3giHo0mb9SthmFpr0ro8kUP+nk6S3L7kypAVUnfvatC6SxI5
zSeS+xo6KFN4HMHTV4xEGsSbYpTF1N6J1CNcQLbJOg+u1K8jBTQ1Ks0B+H88hIFI
2NvYAhGpzck/rZKZIi8jVBU/wRKxCPbmkUeMZ1zOWZ6b4zCphcZnQPp0Tn/e61XQ
MZc2kJGgac5MgP8+cjywVf9wsBRcZLYZQxk0ZcLGDlWHbEVTwVHO5VnwKrHUyBIf
flZvpaI1u13OLGleqv18uEwCBlNRRKqpGikraXt7vo/dlV4m6Zz6jWeE29C6f0LW
SBAYNZzXhx4WQsU8Y4I/eTbIAloqFn0VQe81td0sRIwaqWQ/U3FEig8H8rPFibMT
22KurxdyryUugcSrfrRnLwMdJkLh9/1NSQpSigpq4A46B2jAz/5SrUwbLdGRf4jT
YGTAdLMabRbA2+O75bu7Asx0WuMj7I5siuTaqmBUb92LsYIHBDGgC8j6wQk7/7Qz
+qcMcw6KQ6/hkyp6rYjd5JQc6cHbWFJA4b7kKPUWiloOu5na37keE8VQPZ3x+s3p
pK9zLmM9H6EALGX757ujRceLy0jbeoUHy5znAAcq0kwHQx7Li9pn6LbWcVMDQPlX
armz1xU4GA4/apCjgbyAN+CUrkVz/HYsRJo7Oydl6YeCAltWy/TlmplXzQn5O6HI
f+SKttUrbbZAXP7gmRI479t3/xdrrNN/uLkdDRIMJ5LM+W9YX5pPz+UPughvjqcD
PU6aGpRmJkzq7bI6QIAopv2qRlSiiGpo/HyGoZU7ukLBfA0N2FpRj4+jYVvCPMlD
G699hlWhR/g6snln5AB1haz1Qxfs/hozrXGFKi2gjVDjDa1EXh/UmatVcQ5N6Zh5
WU4ihVHDLQCYit+IpzQ9KbAQp833ednP8v6TPTTMndCHlsml/vtifNiVaE7rGdvn
VJudp3ym/+kgZtHUSQ/Rcg57edGFxPrJqrD2pwW1KS8b2F5E6n0HeKnVO7qT18Ca
2wKn+HZ8xfMZnTmsqEPwov+nHxcAYubNZylM6C7eL1G3zKmbWMrNr8nJD85fmFpa
e0zLMQj/cKTimJJgSL2IIrwiMTIRavOgT/oNHQhjFY44DOH0Tjtaoz4CgVGIAngb
3FrgaJfRERfv8m3i5RZIhsfVRbniU0sfcaoPDEHmL37HxzA/GP/M3jJZcDYnQtq9
hiNrOpdJBENRLwX8P1B+Z1a/1c0/2j3IbF4ymHrwcsB6HJQZ9bLLvMjRG/jigaPX
1XyhCtqyG7W18QWNcUrrEB5qpi4UpYxIZmC4j25SS192bfSZYUpaLqdM8X/3BlZl
4sb81SyNutThnTfRnpRrJtvqeRL9NndvsKcazch9HoYyRt60tzUI5X/BAENORv+J
nwJvLPLFjpHhpWwmdzmfylNgp2gm9rpCGF8u1ZznBd21d4yFZE6/xUoFmTneFAbw
+7b8aoymFw/8T20PJ3AI7a9SUNdL/UR0FALKE9ymD6rG9Auw9zivqkrWdA7SrSp0
t96mZh1RM/Ob5+q7gO16cMfXwg6zrwT92dF1jr+GH400GYQG6axDzLiFsUDvS8+P
MTW3z9d/J0mTxgoDqoQbiXiU082DbezLBpDbjQ1OLtbjV49a9Jy2tUUK7fZsBCOs
dW0tpL6l4vN4IqA+psbZ2cbhsMVmXKa8RfvrvHH65uz7DgGbhudD/dypOlaQ1I8b
8oF8nxNbO2R5YZPNPCMxft023hp9rozO+Ah2AjPu3yYsncV64GePgv+ACfzRG4lE
ZSGzngtqqSO0VoNBF8jfnjf22XVNsJQd6Hwl9YK0AyzuZ1817Dh23B8hlW3acltP
ppiuXysgc2uSQv16uVPDkTvE9MfhWmrA44NTjD9st6o0LYcnKbTfvH03GZGoKxGA
p2g2Vsf1xI6XuXSqWz864gRgShlUnoma1NP8A678d9ycLFdvdLQaeXbQkFDg0cQF
2IfX9KSp/uvnZxzvCJ1YQvWJPBtuoo1y0lt/u0BNHlvnSCLvXkYy2lSz9DLrfwnz
Mply9diptAU1+sRsaY+0rYIB+iLlxm+yfjs3ua9PaNtEplnrqxnb+Wg6KD2URVfA
mDQX9zbB0Jjzq9IQJiIDvODr2Gf4fTAFoFq4DNvb/o7ueAC11mzQ1sZkUYreOZJ1
uCO0j2EWL4ky2TAExJLAGQ2cWpK1o/B8iklf3f+JyWw3o/bQ+Bz2QTdT0ngwwGKK
gNGQyspxSJG9IAqBjYxSix3aM1q3eEHF8BHYreSuBxwnR1Jgz4Y9CsdGAVtQdjHh
7AryaOsSKYYrASQwLxU7J2tVuoZ7GzJuxRB1ISKHiNQakwf6en7nCQOzIyhH18Y5
A8VTeyu9KX3e1aA0DLbEt2U8EWHLAZdXPBQv9E7G4Vddr3wMlWJ85YyZnIp9/gbV
4ObycHYP8eMr2ngXqOfiYQlgZCZSxgXLY9KAOTkeJBGh73MdylLvYQfA6oO8G30F
6qQucczl5QjDwMukjjjpiso9puOeiVS2dE+cSKGbOV854YY+KXEHlEYdTUKsW0yI
mr7VCNef1x0L12both1ikyMLck+sO5awZvd0PHrgSQchf5m4CXH90YEV1jOcvs5B
4lpJaXjcOROqaSLmkhxkpeLpJWLlC0cjCB2HSyDxwtsqcPEcLTllTSH+qGturw3I
4aQlIOIKKEDY2BoBnQQQmNzpigzcrgGwEkwDXFacc7ukrxz/1ZTFhrHIEBIOwXak
7L6hsGWj/ejeSV7d4o7NPzzDkkX3df201BK1pEiPqnMzUcoNeZnv59zN2XyNSl4W
HDgybBSnTwyXunr6fpQbyExtqZ3rVZ4+5FdlmWTTEhtmaK3hJ0XCDIp3GEXfGmf/
53l6+cS7gDIbUlJUDdGBOoXA3RWC0VnUCePNmQ0X1SHgfKViKeqps7yGnckbdvoU
rAI4ZFVM33lkBo9JP7RKDXHtL6CRVVQvmffxwOMGA+xHCiFez9QR0Rvd7rH/19Ya
+wCWzspDGNssR/C1EhSuWLXwdg6IlhxkPRv1hKYgPoEIaJK2PW3aOHEPcPs7xf/m
cJb7YstDDu8yBq0Y/ONKrhDKl8LKu9gMVhdS1hc7f5r+xXJt9OHZoZDNyxcUoAKy
Ls0n37B3xNa5C9Z1YrBt1soALuUP9W7j1lE8LtFwaTs0XaZMh+BRXS9TAlUVP79H
/DxDSxMqFzQpL5FbquDHykrTkbGouYJDY9Ez8rkcPz28MGEnC4rqyPtZH/XL9J4N
9m4HgloabkTpHxv87q5xx1P5u0bPTVpM8F/RqOqCMaP0lLD0KlG270hN0IAgAQ1P
gQiRP36O8YymVQU1FxVxA/yOhealKCqNemtscckxtL6Ojl7gU6ty698I9+b9MchN
fGLXFJ58rn/6oEKBDBjTfZMHV03YbuZ/ftK0mAXPQlO5P2zP8msXWkkjRVjkcPaY
DCpURtn8nYi4rLJA8b+E8XvSYXBLTOO/nQ72ldgD2vHZCxXaPAoIrXAX9UrTT9NS
Cm7RVtnwSdhgd7+hWKHoiSDVpb7uI/9b6W2GOYY7KrfsYgi/Yc2OM/iVeQ3Pwi7N
cdP9WzUrFLSe9r4PXFzLj3Ch3VwA95up9avafEEpSkwQ6m/I8Tkxj6LDZfdiH/ho
y/w/jKXe4irYCjd11ijbh766hovJ13pnj2SnQvd+qaGIpE6oDHHpzBsUhxQUm1Pv
Cwr3RELzqb+mcP31MrkJB/yDCctWTC0fl9rslpziUYxElB2wUhCdxRa8JY3WxCbB
LsVxltIPMsM1VGvA9ve1MFsyHIL6Xk6X53iVCXIL3/DqpO6NHivDsetx4DnvkziA
caEQ1v5zNGHMXRQJ0bQ+Po6xbvlJOYLj//ybVP04O7J4VYQuapIAMwXc9lKfHDO+
Fm6SAIRM5Eohoim4HMfk3pUflnJsFmLGlbn6j4YrFRLM3Ia+YsQgumz2R1Yvgjvo
/mIKkKx5v94Hn8zj1D0inYRkUkDreS3XQW0sBjjkYroEt4KqV7ORuH2g8qr4fHEO
l1YQbhcOdeLHbOsxfpoB/EpBpG2e0ms4Y+EOjzqhZhabMoK/FC7AslAKTFI/mCLW
xwmFfzK1PYH2aEMHrnA66/WyMt4kyByQSEEZ2Qc5VUqxe6fUijBKcF2+vQZ43wkE
+PUeLA5NDJE6aW6h05bNzFcW7vMjNlvRk+hc5egUTpCmMBeSlaopN95IZTUqvgdN
PGWc5aY4csR7KxXyAUap1xAs2tEUxwsWCTbsZK+DCbeLHByUeO1fXY6tTWTEjROW
tO98PvLIktgEooXgmaBMz1x13H7NF0cXCF2fYmU9VN+Zbbr6hf422XzIw35cnd/6
P+he7LtM1MW1+cmb+ASeteTD1WS5CM+hXo+8fjfko6DKH9Viz1Cn/DFzC4ShKV7v
/xiIQIXbXY1bv3lTkbX5QiNMNPbwf4ca9Gg9vHnVSrvwcNAbt5N7ny/SOxBLZjd4
90zJHgtZhslY3uGjG0SkramE9av0cVy/7bcciLSxGMbyov3kb4ewKI0bC+P3OWs+
bC1Zr3vqAGy7bhv1OQK5rkaLrrLbGyI1t+tQ6DMgvEq+RZakYTjFDpJ5aq1lDaU/
pmnPQh+uFnC+4tknS5SJLwoQR8FAYDmVKM4xQUxqiJIMtvdSm6l+/AswtrWo5BcH
wBO9TQOVlmI59wuB9hKl/8nSSiRS5ZcvAGvuMo5Bm0d717HI2kW3KhEHVj3ncby9
a5KlZzU9qMS02j8ISV5p3BVyWt0/AZAL7HZRbGQyQYMOzzydSIOIwfLuvrZwJ/JY
FZ3FUGh7JUMBUblRQJDwQ/gDuZf9Kni8bKRIV1tZ4xz+77447tTtLkxzBhnyYI9S
Egf2uOjfa7PEkoMWXkjb9KtyieAKv3MxRaoxIE+msSebiyTnGVZimHDGzY+0xhM/
0l8hulGRVfDEaRVAs/QtZEP8WWGhf7E9XJk0nqb7nqrYHElI9anKbQNJuZ0NEsOo
YUWelxV4aASxeSHHNsxn0DZWaRsJ63BlnDrEKTsyFE3B/yNhd4Xxtg+POUigz/Bg
5F+QqXOpZQKxnhkTJf//kKuc5g6N5oItY1Rpkn9WNzj1eM9E6jpx9Wn/xCMwC9gk
UVVe+FdGrdov9rBLKkUgYTediKr+kVeUrcqJS716gUDqrRHC1FMgvPtJqFeqWFUW
DnlS5csu8jHkbPbRM6rzY2SO4DWX3LyW76NSMSJWcg0Buq5QpCq7L5yv8Y/n3tX5
R8yqDFN5JgKpOXIvWLDAR7ORSwLP6K6bMfY8FVdM4qI72RGl59Sk8HWuTy7SrO6O
lspsqSwgRltNbRhB2mRvLVHktmnj35/xwKJcY0sMd5eT1x5teLRTpC0FwaWyRL4y
FkKPgbNHNGTcu/M2C4oY7nkqNvZ5Lc2dz666uFnWugYFeNXfEMGx4jyu46BImrje
VpFQylJlHxdEDm/QsTERJwxcUodjdfbdMLxRJjEvdAAlgAxsDrsf7PhYdvQePWe1
GIYVq1bh89vkW9VAGLEQ3Rmkh8ATdar9r6cFcoSq7wiixZZPAiI39GXQa8EXZzuN
kHKP7sVRzZXmsnsxM1CA0AFu1wIcLofX9J1h0rXsM44uqISxNtqdzs6/276aZmFn
y1FJNYU++gZ6PwqOTwPl/7yhgk8j4GPDtcLcZvk4jWgBLsjYN9fl/mYS5cBaL3U+
hyoRSX6vLBUl9RJEQtyNnsWMgkuaNdIvvKy8ED3hj/vlzVh+3dHIDKFQ9h00OuWx
wmOVUA8UYZnGSVW4HMGRli7L+CmxRzR08zEoNr2sqEPa9JOiqiJGqohyS0PcibMd
yrOTv98szcJcUao5d6FHPcspFbfd7efiYFfO4uIuU+s6jso9XYvI5+E/JJm+o/u9
65ud/yAzxuAfvNPjHjTMpv+ijB60K+z6Murky1faDV5lE0wZ6b++bQDCav//QWt8
djYW0MdqsFahAA/i23vnKdUsx0pOujq4gv29DsBFMsis9kYy66JuvpTtciYFQ1ZK
uzW0w7YidTdp7s/6kTfu3mb9U+g8gjokpS9eMDUs0S1mVYJ9W7oq+QXrv3TML5Ym
QyQNI+BtZH9kdveuC66zGlembQvXDAWbrriZKBf7ZgMYw5d70LHrayV57Loz8dsv
dZ/MsfrCq8qpfGZsVjAJNUMxitAFnFenFyLfRhIrDv/paXCuvY/4nTv3mbXxT1C4
dZm41pGMsiYAsJ2gX1HavL+5m4wcClGvuV5fhO/K3X80Peb5+TAKC3NM7u10v12W
wc6eD4nVyuVUa7yVzbhi9MWjygHlsh44J7i5RexhOc/OK1SnTewUdqM0ffsMnsGR
al2wbe7ixzam5mQ4vDXpNqnaLduzjol3NJ/bVNZNgLSsu8i0tsVKWSRwMaF0d4qw
FCiaru35dPt/G4XM5bpqXrITtWMvSlFH+i0qeTy3rGUpgSd60rsAdHhhr1jTp3Yc
rie1abZMT61Hqhvr3uP294MK0B7KLzB4/ukZ525ZvD6+Srp8uMdF+fwUBGQUhXFo
NyslL970xEEjW1FhEj4IvRoAWCK9WwFy0hME+o5Nn90AHCdy1ydiKQgOaYfJrJCu
3F4E8Vpl3L+/JnjlvIiz0F9ud7XFlOmnsfrivxLmuutYeBchP4AiJFF3zGaoBUjB
KZpOBrwLkiU0yJB5pB7+D8ZDyjWF6Yyok7L+/uk7i+n5WCI5LKexjhtec5ZcNdYc
8vRQ42kCxFjbidApxyx8urcjsZbQ5mrIvjQax5nUcE2nRkcvoWtgjjfTxaQub/84
P1i900Pn8YQ2wCWMHOuncIchQCUGYFn0hBwPOFrSLB6NB7I73AcmIYcs0mOZ85dS
HM1akEOLnvZfJUkJwzlQiuA802jOYmh1BuMJQMRPwIsHzr0lIPi0Kq5SccAhk2Jr
9EBUmEFGuHYhGnI7/a5SxgHUgxGXYySHtoQ7onHPLFM0WvY09KQOFvjDtKDkjCyD
Q7AZDp9GRnoIdos5OIaQpKRiBg1U7rp+7I5DTnUo1c+dqAUDRn/tiljWwUOChLxc
e+FALEzXdyEsKzOlNtuZ7eBLwo0TnrrF52G3xIGfytYDYkamp8sknPeNEeL0a1GR
KuKFRZbLa0AoftEVSvFspOryb+pIQd+uOEExP75QrLRswQl0iJeAnHhP7Jhsy1ql
Iqarw/5q0IbhgukYDXx4hHpFqdIIcy59rF7N2sEcp7e1IzDDW9lnkWloJo4Tupiy
0Kfu2Vr31U+5joRjVQgGpBv+PqYaiWHTgj1JAoo4P6KJaFYYh6iEhL0JAiUMGNnz
H1AOOK+pRAO7E8a79JVclqGjD3WPIWjHpCAfYP6dIK+fDc8o4MGn/KtOAoGP7CQ2
M/QOvghSMwxu54i8xdGRpLTSSTRccyZYo+jntoddkRcACFoxzo9Xl1D2eBgxl+Aa
OsmapamBrInoMn85S/eYzZXZch5tCvxVBLvtO1A7ND3blGLxM09kwuuyrds52r8C
jWE9zE1KSHvYU3aumSRfp3RRA7UnRMangTgmki+eYbriF0nVTaXSW1+4w8w2nVnn
G5qJuEnFwfTitM7T/GS9Ai+LxjFPaHEvkIeSAsNWGMC74nXZpY72VXyDnzndkxfM
0cF8EtIQfpL0dFPnMtdn3n2m4uiDfV2J3ddrC46nMahuw+zbQfPqwFRjx+DWfRwT
2+E2p8qNEAFgb3+0PEE7A06gHbPfsjYTMZIe8SFE4gDUGPeen2FP/YbzYaQC9UD5
Z17HgQjrPtu7NsZDbfjKn0eX2oVkhMtIVh50Vx3LKyFMttS4XSzjxqhBGwCDjKit
F4QSq6reLhODWgmkpmcQWO7Yp1/F0f2m0ZmP9fz+28coyK8409xDHfUn1W3YNdfI
w4xogjk65QV6Fl0Lg3xH03PspZrvXb7pSg4iJXkJFVxdM3YY9y/c+S1s75snvPtZ
WMCGEigUMpSQI17TwQWjEb4t6KB5GD/gM8ECecjGMk0RH2NLvAT8csX+87BdtsUX
GBiQQAUtjZW9TDnJDmhx6tdiFGUwNPEI4l6pRqtJL2tPCNGEpUlYAzQtOWvDPe9B
4x+liwtevYJehsseiiRDSvhf4huAtQlPOjGK8IukjX4GsoxDIhvCnGcQA83ySoTn
inDgDd6fNoQB+6W8jP0QUH22wqdsrq+GImnX3z2kpYEtc/aLsC0tjc+bn3urkxYh
873PNrZRVin8sxtTfwRgnbri/I1jYj7haYbRK4CWmfue58m4u62R/CVx7A3qASai
XLlLZ+8qAkcgFpHD+XH3TXW48QrdOZjw5/oJKQc3YGcrGkfhLK5St3j+KRKDs6N+
irUHHgh/SJyKUjUewAQVK8JYFpgLLG52z1iM1jUl0lr2DnvgWAYZF/on9e4EwGba
zVuS96cgd+cggegC1LLpiYA/h9ifcGcHHmfnsc+Q8K8xiGPJ8m/vHi5i1ao1Jdgo
BJCMge4IMjdQl2oDkbBs+coRtKIg5jT7LDzlNREF23nOGumElMYEIpTTgLeUbLQb
b6WNoARzC0hj82sBOCaCy06CGvNgXV+2WGeOM1rnsj0SoGveYDvY0Ve/zx5vwT17
tmAAetX9UbaRAIBu9f8gNzGgvnfNsNnYDWjxjfmkkvIyJelUuizjGF/ZcjsdOk7/
YlCTQDBXD/KIFv3N0IfQ7rnAZeY7F9puJTM4JVQ5duJ0KfMT6XTC6Qzy3Fwh/1tx
Wpj1rjpCmLXU3oeLm5wTzZvLq9qSf2Jy0CfxRTBoXy/JBEnZ5Ogt5a0RSwSxSZgG
OfPiMlE9RhtmaouLVBwBe/ZJ1JOAbxW7tx05HaQHd0AYLqb1piW8nWj+wKugkwbC
sdkR5vfTtY2zPDs4nBVkiBXxXNn3QMCIetB144McZTaJBOTgwVsheG9OG3aJza/6
mn9OW89fSx6cL8zLWHytRRYH964vLqrRir4e5diZw22khxMuaBxkhN9hQO8JYoRA
N91VopdyQLP8zmhGhNpD8nJ0tbgU72Ys4K9TkDn4eboC/sKKIMxnX3iortwgD6wq
pQdxY86iWGcWmrZIhvsHj95a0Dw6oqpIW16xl9e2w6gzhm3gjf/pf8y6aLsx6NP1
6Me7KMMBRFXu+DOjsUhujSgXhWfvbcqHN31qV2ZyqcNpvqHm0hzfH08fP0RRbB8s
BF4UbJMl/K+O+kTvT6+VJwVLJSlHl8TJptpi1P5eCuskO3slFP6nO2mwhXZgf8LD
sV6BS+2EaRrhKeu9m/5/nwGpmZtHZ/dTECKy1xuFOKpE93ji7qSc+rRqCcmHtDDP
ImQ4fYcs+CNED0xhY0+BjJa5Rj0fCW9O8ftwv4JgB80fnMe4h9GCiqAYQfSyttBd
6jUp/J9VvN86lzKYzf6asIvlsHvRJUDogkW+FM+SOXcAd6HMuZZUKW7dXu0E2ws+
Ns/b2oWIxK84CXQ1c+Mf9ZxZHafzaxyljstVaAhsSAj65QTp1vOkL7Qq5ML2m8ar
bpFuBow8bY8WTCAcI8fSE7RuQvrW93bszOOG3KTrjGyFsuG4uqEYGBXZOGPmct2s
JcLTGv+TakBbShzu79WKWbDOQrwR7a4D/9p3ySWt3m+A6e2/+puXccN4Qqtc2S4o
oA9DooojEfSh8mOITTDSPLOQDFz1MXODa+bkNFZ2Egfxidaj3D5yivi83zUrX1Rf
ly8FCyd/AIAIQ0MtQkkSttYP90Hv4Z28QX/pvjUb39oXHPS6OR/yhCAuvHl1I+P/
WYicHvZjVXy2nOrHOQOo1EIzYspic+A2BoGhkk6ppWqyxjralvIyzi3nhrbSPI5n
cm588oSnmleuJnHmLsCtIjRJCtbnJbFFugFPrcrMDQFIEghVU8s28zs5/nCf9kcx
XgNekg0KzH75iOKhg6y3NfRsMkcrfbDqnJXFrxK3y4V86mqvDlqMrJbQkUtPxRlJ
pGmjTKRtddkQYyf2WxfJh1sn1BGg0mIXMEZuZASahpbR7Po3huSmnWNAg0LmTbBe
gsPxKGLKYLEQnTx4wn3S8RCRe1YdOuWDACSQSN4lDmqruc3aC4OL0CS29teee2Dq
RpUv/ttumL1SmkbdiAgJC9AVPqHi6uTRlY5thA2x2XjnM5KkndeWr/J9d4rxYVZ9
KWABMHWSN5c2TXAXpKmZeeDK5LcaadskMJhwpdR7EhhquGJikpMzfUXvYsFDSq32
/6F38D36qpHlE0Dkdwqaf0/d5A3apGtozDHrndIg15qE+WBElVdeUQ+x1RqUKV2E
qftyUoTt1RxWivVaCsoz9dn38+mtPasIzFu5q3dLLq64dYtOyGb5KXYU8etOWjLW
oY39ro0clCpGS+MiUPDrq7X2f6ZGq4+Iq34prbeJLoAMphaOBQUFLMenZhhni8RV
ZXU+ztSQBCL/DBFZ1wR+QNl9qL4B3vH8pw/KR+6aiXjkqTgloswLSzOkQl+j2bg9
anYvijzVDUoPxv+yp4EvMvuO8UIp8bcHQ0f3g+d27zjW9iW53grgGlUn2vdNu8GG
qeErggDpZ3qkVtq0/Zwc8Uxfdlb9Xyg8XdnsLbPFDBF6KQRXnxszgvzrgn57FfQW
iDwOiQHmjATmqjGNFKd0QUp0x0Bj/h5GhDFbDL+b/Lenm1elwNi8VDq0ade00Lx6
YHt9VEKaN3sqRf73sF08LcKGGojlLs7MJWtPNVts5JXbUNtoZfYlcjpor4H/fy68
Z/gyVv0tHkF6hENuN/D8WsGbQHB4ETq9b3XAMvy0wImQg5QfjcMXwxs2BVyfYcmf
pFxDi27dzs5JV+E3ulyRDuvBrqj+8NV3eFxqrrpQ+DnW84v1wfvcET0Y0gg6wwRy
B0FNTypcuVG6ZlmmW0BNp7PBvchDDWV+8d9YLcTgK4V7p5heCoEBkEeQhF0ikM2L
zBvFZ/TRC4dgC9Q4tiwX8Z3wKu/7JaKxitNhiX/fqKhs5BxtliybR7P6I1AFIRko
gZJBmuOgchSh5W65Yz8kxbjVI7QVpZAH4s0J5ufZBFJgQairzFSOVnrmcHoISVvm
T/cDuVuH8OwanJNoofGWYkDHGa6fH9QRJYB+e5Oij8kp0AhsyuATZb96mFX452bo
cndUurhqRKRJqB/ttRlUy3k/f2/RdaiQfaSiInFu7pnZGuCLWyrupIhjyDpvtNLr
2GjQz2UVw/UfFyV0iNayMe0zhPgCEc9G/1iSJjBm4b6c9WZF1EH8fu9i6+h11EHy
dU5qaFz51Ywxyk0XdtWNMc7Ip2xoPIVjkR+H77nnE6LJy5Kpy3hg26RL3j72qVyx
WpSn6LNhrpV9vds16FWgHHdk+HcQmAN2DXhM6QVusx0iEsBKOut+D9Jn7Yw0wr6E
0GmlWdO9007qpZDO9u3N0j7rOS8DHrImJ7JYhpk/b1Ez+6D49y3hiO2xlAeLzFaH
GYu+xTMW456qof/S5VxTnDRg7SXBINHIgdmihtrBKYqIQrWy9gWxmNBJqtaPEMNf
Nn9r3zkIwCAoJPD333Aigjs6aW0cVS4Ngk3Sq3SXtFlqn6rTCOPjUC4jgKNHFy8Q
Xx/Lq95ydwTr3WRhGrabdMxfpL29svtgtm2FudUXDWxjsEEc0PbJwuRXINsQkvRi
LmklvnsgxKQm6gobx3nmcg4EU7CUfuFZaZSilPuYMaFeuHXj9DltuUHmeScCj3lg
2nJ22bhxSF+EYw/fubTy89/K2QKlbVC62PeIUoMEhXK81ySfYPjN1P/9sLRFScSl
/nVp8DXIT2HnrOHmkXGuO5LoLoCxVzEXS8KcfOMlSexOJgobDOSDE33es9e0Iek3
i6BVt/HLIY63S4O3C+O3VFOEhk69MB83XGs6Wpl6sLKeGO6sGp++u1TgoZ9gCOzs
NByYGEk7ML3aTlbHBrTv4UQg9WkMaPYy6rHqeMMRaVBOCtv7FQ5FzSH5b+hHGlRE
LKnpfMDwXOCUoxw53L6b8dBkaiR+lvGM2gxId1u5uK/pCrqad1EzpghskiFG5isj
J6Mxfxb6RmZHmT8CvVbKXTP4AejsWycA6G65XLLbAd2OuMe6LwtezJp23IqZePFM
AGEUJy9t7AbowTN8cUkWEekeInEmMoH6PoOMcBsjF8hm/Eg7AmvyctUeUnsp9tEv
cPHQuP+FeeLhtPSGGB1N7QN2qrqL45yoSkBJdgwoEE73jMLW3YtFRcSTSOIW/QWw
pNxyrYmA4QBKDtmNkdXeZvCogZ0KEj3P5HJFlPKKIdkQRmkS12XkFmoDfxIeVvnh
pmtylBjoBSR+h0CBZR0y2IkXVPUrFkNtPOckIZ5JcAqPHoGlBdCrlBWYiMGqNnxq
JhPzKCB5nPGMv9lPKDmaZvKAmCULpyxwqsFNkyQErGoRnRd6/fReELirf/PiHE6Q
bcPpC5sZiNtrYoCV9gMdNVc+Z0jYy6g6vIkT2gZrvm5ujoyPxasI7/DaNP2Au+PF
m4hDsv/BwHwCEICBnCOgfZ5yxSWkLuG3jm4s9IAIPtjexuu1195aVVvlETcoG3KU
v4MKVZVCKRJZLOrwXiJe8l2ZLshuaXvUx/+G1mNvCo9yj2H5VF8n5HeVn+7TK1+z
jxFFTAETqYjBTlM9tydFYQm0/twPmDQ6aQSYTsF4Wpm6hMMFVHSsy/dykkunz3JT
OYzkBbNBd8o4nNIb+naaldoW4C2VAQ08oYy+OQaHHjioLfE+cplYFvRjcUGtm3/o
SXDXpwZokbnPeCOV5PiMYCft2j08oVBRTN2xUmu8tP2Ln3TQPU5paKyGg9ZR/egx
91cpAKCPimtlzDOlk3pliykjpBgDUWQzF2W7yP9y4S9ZpxB8n3bC3v6gFUwoJ1Hm
jOr6SsPWDmbDtuxQVLY0pcSQHW96a9ziDfFtcvPnjvSg09OTMP32n7/TJbhupuvw
ZrAmNxyJM6x7xVcN7ofJVfmnO23lpoKbvwQPDJhGFuFjbFCmA/T19Hjhe2r4okLF
TfNB5y8oyfQX7AiTdwLoILyKW2JM7nCgi9Fem5O2mOG3BF/GlkYEJdLUoSt+lEaS
PGTwMRdZNkyry4RysWfUBlCpxCCtyxI3nRH74TfKSiSQL+WM1DRJnbe4DeZwQiUN
ALEDtPHwO1KnT5/X/EkM3MfzzV8XCu0mONqjqiVuspzTepaVBSZqK8GcGR0AD7kR
irLPtGYYYbxMsLNxc/tv8tWIEn8jWeNfJQMPgt/flSbKeIwn6Ar8cK+wnt2gewtC
cOyq0LideX+FkUuorwL2emtFiJZ6M+9f+eGSjv+EUW4CctMWIucIDwuIW6aTcmdo
WPtLp2QbAObqJrL78i7y1Ar8ucLDG2L43GY7IFltJRRHp/W/dqKxXnvMXPgc6PcX
RBMzRaP9uCgUV+Xh0obtUwyx480MX0JW8PYfXmH/FwImzbMSRei1jGsX9UDE2oA4
CnnNu8E6PVzVJaHC2pQ74wyFDb3c427Q5dtUWlVpj0kg4mNFhqDhGmqsBuzqNFLV
uOkLgtaboYY9usf/Ar+WLkhVr1EVSpAZ7WpRSCbQ4MIixdgE9s1DO1Tfczhc7X+n
hE3sacwl0wc+bZL8mzG8IEQlxveF+5dk98oJqzCm6SClbub56ufHiiUrpj5dbjr8
u1jLHnkO713kFFWgyRhf5iam16AZZEyDd4d8ARCwfgE3aoEw3TUoR6591c2TFqSf
RWP9Adey9SFeb/zCecyi/7eBCb8jZfGtMcdSzOcS//5UujKHNrDxFvjs1hTHzYuO
uozT0/imAEh8NLPkFaJK2uBbYJUMrbQhDP597YNOiNZdJWDWw//008U2L4K5vFYZ
I36D4RYTobmmsrtyonZxz11AGkol4bGcP70D0RfUysd4dtVCPe7RAc8hR9W377b1
r6oUX1yUa3QIb7dwghrj7C8j2r0UwIRwO7PKQ0ygzx1puqTFqQfy3hAIhF6qYX6k
pqLGANyDE6jboOHOcgRnpQrNK+1WamGlvY7wZsRrxVqjF0r0cKRiovs/RJKQS3xF
eZYc4C2DbzP7EXCmzj1483wDHgXFeeH+hGDD4deRo3691hra68XgCZ7TVoluJXPN
410kvgoImyhW+sfweHUymaYKGGKwAcXZcoMSAqCe3PTnq4Ofzvmwr7KZ03q8zcHI
KmR2qSh3tJSTI/jhlXOhxcVXnoKtobWjsv3IjlRnX9kv8QPAsODJQxZrEZWk+Cab
mlfC0t1LwlFndvZH5DZyGwXJUh0ffJLqMqdC+duON60BsCr/EkZaEdmAEXs0WIGP
gdGvz7yGZtJbZxkZDJ+eVxwdyw1xs73Y25kGipaI9jGdbRjTNUVbOJ6+A7PElJJc
Oq7bAkAEvzde8h21feMC/E5ZOTqeMunU4dGJTAhkwM2uaD9VHeacG9D2LVJ5vqLj
h0MS/4aklvll/q4ne80WLbt2/CkAWiHoc8QbQNzGPkpFGXHJIZRfq2klJKnpMXQs
SPV3wpKUURTaA8nZ/RmuBnfQyDcc4pY5MktpKnSCjny0sW1dQPGevfwgqQ1eLzEv
7/UOUhgcEwfhVMhC7bKjP/wrtORP6q1T10qKD7l3tHrMLpO24HJDpA98886WpGE3
EAD8zisGSOLGlxpPhXB/GDtcz7Gn2cLBesHBy7EFVCMcKYhqOL0Wyz+DKVJXYvQZ
fYL21FIOedpVCgDyog1i9aWwkDkzdToYKKqu9iIO2qGfdYNbWq2bZFEyS/kB0o6S
Z0V7dOJ0ClLHhBXNV8+CrVjKF9mCfKw6wkEt9U85+fr3509kCwHl55CLVDniHSRR
2j7jh2nGIW9sqlHD8RWmRYSFH5j40LMWfGf7moCm4H7F3i8pOxSQTzAYNqJ4E1yx
f8pfSbC2hnizRst9GubCh/hmOSr9UODj8ZCkuPgwShwPpOQIYebSyuKFu8BGxnLt
3ra/0yGY1UHf5uManMimgcm6DYQNqryV+Wa7sfH6h146j24T0qHf0M3Qz6OaX2Eo
zHwbi/O7apuAQVlrwRN9OecC8jLC1wUsXGjFAQtbhnaeLE5svjjrcE2rae9mmJkJ
cWSr/q3MglORw8XTvWRppOIa7Qi5tzC4N8KtlXOiI+5yPkS9mkOnVm+RYl42uK05
I/pKPqauXyQyZiFSN3q+ZWs8sO6AEKTjcbmC9xl+w1m4k+bH9+o46YnozhifjXUV
0w9Co6R9XunvJ9iIygEaaS7G4OL8zyYuplVEal4DFAS2bpKK0EzQTOZvk2Gb2U01
f5f1DescT1EycBFgtQdpiUYO1++UnIm8OWHApSmMVSywJmc2a34yykYl/RbdJwPf
DVP6/FwAdh8GqFniyT86n9zofTLcJtClxIdqqyAkueoW7zD6yXu/3gnbDlGDX8jY
Y92MqFBwPf5oNNssBOvY4u/g/AFU7o7WhiEplRNIIZg4d8xo7ApGi4UhC7JsjYFo
Cfm2bFcN6fCd2AS8AAaAKvJWC5Z5aC/YjTouzDj3L9eBONJuHTVwicXrfbA2AP+Y
SJx5Mgo2x07xob4NIv3HLT3GLi0B7kdaivj/D4BwDbSeFM9Gfi4e9zq8QTF9RyiK
ze+2tzsTcPxp/5eRoe1qIBgONmsBGrkhc9syXpZNt6SU9/oC2q25Uat1BSRdKnYc
P/kffjI7IAZR1XxZGrlwV1A/X3oBF15jx9J10ipRQAHc8955vGiWu/lj1mq9LLQv
LNDVLrS3aOzRw+Y1J16b4aKqxM8RqsmGzkx8CEiUL4fO+NNs6Qq1Ua+FrCgY8DP+
xjawNI/4hD5CkUDykM1Lvq5lbRv0og9rgvTJR6ci7ru2HIGG63cD44IIQu3zBqn8
6KGBEgOF8kz9cyMPH86IYzfp9neokrSjg3qbkFF22zIRW0/cVIri09oBH1Mxaiqc
fFezDXB7D1ckONDoxzy+1HQaLz5j8/+dQAwPvZy2gKQkIyA7zprksYqqEGx7t6A4
I7Xtjndi/vA/csAWkqbHgRvaUHk8vm24XJH6ZD6awelpGVZYp4aHY6DQL6LGA9QH
JDXVTbq8aBDGQx+TOYAtqMuvXb1+DuVsv4VYYX0k2CVlXxf8JHxxb3Kd/N/FdRDB
aJ8DF8uUjQvFAT9MNKixKKcfBFlXEdrRUS7mbxXfuQoU9ixq1mbtHeqpEnZnlzzl
a1KE/nmVS+bFK+WZzJ1R+CPsbP0b6IaUvoBEEv7Mmyo6Sx3fW+4XJYyx91KnXDl0
hQ6Jr/Dn6iAiPqykTq+Zv69zl3awt3saGwYnWG81w2Yma0MsfL7zohwZSA3w/Gqd
V+1nmdv/7Ze2GlngCXkSdLf9CY3w8Z3ZCI59/iaOiJDvoTYsqieBPr0x0SIF8ge3
oykDYmqfcHPmaPbuXv5+uOVh+0VMgTFLCu6VoshoKp/cmMPk0oikXNp6uDyRTXwr
HfwTq6ZbZkCQvuEOp5BeekXV+MIQiMCdw+aAAveQgWE8NM7KooBi93jGEQvAU9PE
dMLc25++4Vs10Gc/3UYAkBhuJv+09JddypZSM5oIajMFCdTf0QI3xzElZkPSydwV
mfJT/o1X15xDxo1MlpJavDSH5VG4TKsfzn1zkJeFDij+6DwMExibsyJWJJhQ8oBz
VZMZLYy+CFxjFo8xsHSWrSRrajBYhLZLEfzGnqGKtqAvris2TFpQ3k7BJzCPzV2J
2pyI4poj8Pw8qh3A+x4mc8GgT+49oceCANN8pG4rB15kDeIAshBpnuM5ABt47Z5Z
bvfFn0rEzMvERoIPKDTlKkmyXqw9NLD91/knbXIFk/n461OqFN4zeNKC0R2GSUWC
JYcyQgGRrOo4ZkwrnK3yO0nXzhKP7OqhUd3687OwFLPhtvhSq8QCpjuEipI/LWCA
ERJF5yBi5mtnwIrjM7iahaGZN/iqg/3WCVUs7a+K1AGpeTU8z+yfiRa1irMIig25
sWgHI4BgM8hIrKXIglgao868vHzekmax1RTDtd0VTjFUIlXMTg9mZlPJ5/WrsqUA
qWOV6RRXoxeCFJKRFalrmqKtaGTJJOD5HK7gPcLKWJRV2hf+LRpwi+Cmb9bFLNJV
m1evMvSGJmvjFF0K4ZBiABJomBYbi/YI4eu35Y7Ftd59c6LoF50buKyhdx/cB40r
1GJOjqZCBPv3xCgNGec0KsquxxQZlYTx5wiqp3cxg5iJ+VvqQ3vzwBSxPERCPMaQ
8XmK0EpnnJcWnduOvGsPbygc6cYO8RrmjIWqO58aSvoiLtRoMqt9SGZhE5tlLi4+
sa87X7LvzAbbv8Zr68hBhiBjuqmCLHAkFv7HhCEqoJqpN5cRI99rzF+dil0ZsWb5
e+M0wN8lgxqfrSy9Bd+CdseRz3cvHaBoZ4Vav8Q+50r3Xd7txOBLYc6PY5RHX2JA
0I1O7rvQxruxRdY0vrq4hILPLaoSn58rGyu21jsfe7V/nXpRi2Ic2zjJwwyPywB7
nDpKPc3qPntQ+EsbgT4ImgbjseGWIq8b8zUZc/9nLDoYufoxRka4fBIxt+IS9TxV
AXxGell58X8GyRcFo2FIOZYmV8eTswoHspXgQ4dU7Hsy/Gwv8NxGXaFLeZwrMjrR
pbYdGXJ3OWy13pbn5S686oNjDtQ8FZfpic1N1e7FwN/bpf5J07KpQ9npdHO4FyOg
gYml6viMwVCWItaWhM6h2Uz4RBhALstojVLoW5/gJmYMqGrZMjbCDWo8S8zOo1Xm
GgwJkqxAeAsenx/VvnR6W534/Z0NPZx/luffXG29/K9YyEtSIHiLap5cK9IKDoHH
OxL6JyXy0T3u1Y31abtkrrLgyM9q2m6iWo1lKO7hTiaim1AHTmsByWzh/jBLUUGA
6V1kmc4P35NqDDIVtPUlsOw3jQR1hYIeAIxqoUBBGOHqzZTWMEpnnbSr52nc2zzW
I5+vBr6Rz7vux9i3XCCuVCD0T6Yh0TIC5jXLeS87uVhW3RjJew42tgDmUo9m1Y5R
Hd2FGQaKE1ncvuwye63ajHZyO2T5C4tXNoyA0JU1LgXM7fDIMLwh9rJIbbZiXWk0
/oDehestANTQnItXw9IasQz0AUnGZjH2wcFKHurL8fzcEujpcKxJXfN8/RqQUZQo
P7woPdAKRLrpLE3NEnPZESqEtYck8WLw4o70rgWZACIOvuwYG6WfoCsUYeVwHqUc
tWbRWTByiTRwGAYBg7LnKToC7gxuUdVNILAf+DKscGijHaP/M7oSJseUNYWuFRe/
XBDL6HtAe7LZ+20WaQUzTDgXbCAovJtZ+e/Wvax7oyiqGpJ1I0U8Hd3alod43lxx
tPtn51rYL2Rsi/qpsgnEMmB2pbvqiUccWLGGa+ZUtdtwvqAktuctCL03Jd635G9e
l1bnytiKekzlHxFogV18zlz9TpXndwLSzX8EUyPJzzXsw1A6g95Z7LoPTLurZeHB
NJGwvQhw6rB0QiXr5+XpgyijqZjpZpi5fRx6KriXzwXIGvUYzGzR5JX6m2WSyzzK
hR7DbhUuX3I4aLfw8g4yYj4R/ES3gy3r/FKSboHZBUvOq+4ivQ0uzw9/Ob21W3to
5ytFEBBMJHvBSKoairC6lo0T3DUYC3bQE7mWv9cEZd8BI2Xo9odNOSJkVs1w7fKI
c9z4a1uUvI4uwwoizLiFlHshSIlhjpH64wX1DAyihI3mHXwylFocVXZXm2gmlQeY
m/g4RKPc2+XULOEhZu87p8AYG1qyxJIWSrJGEo2fsdNq/GMF85n3M+Re8USfNRUJ
gE3lFT5HpJIc8hAktmPPf7I/fEqcrCbqlA+UIdFZDWuQ0/TfBJ9R2VfDfhnP32H+
xjQTzQFxDDpkwxd/7HxzSfAnIFVFHY2LsbtMxsMiVFo8fMgQJBLD5EeZ3MOvksfA
cNJPvXhitgAyZFsMEL3ZWTarMf2ho1J6mH+NzpsHK9an9XK43IzBY75EVmZYNZES
3+rdrkD8+b0jMANf0OHRjV+wGGyt4doq1GsAPPcBva4+XGK8oLBDODdJ5Mno68cx
zPIBdVsCKYV2s3ge+k8drll1KNelKQXS9aD5yCt7by2k35jlNZFGWF5XQlaiYK4Q
dXVHKc9s3j8AGpjQBPX9QAerEn2CuKWsDaaPCfINzhcGwnpdEU3quSykKrinxrw0
KhvHHdbb/KUkrGEFPdsNP1sAxV+ftcwgrRBWUcgLn/m/Wb3FCZa1rliW+KlTYedi
Aqcr7AmfvAAdYPR8TBbG1YIwOGcMcqR1G737g0B/gISb7xJRLIN2UODoU0+Y4HRo
KmDmis1aNgvmltkUspFFB0VbidJj5gVAQC8m/Re8p3hH3J2LO6tpmYH9MlWDZ0Ie
jBB+6t4fLNtKYGoiIE1ki0tgJaui6ga4LzHxRjdzVOff4zi6fQ8YGKfzpZQyHQ8C
r03cRpa5SSPCGwDzD7dl3RWi9y0wHZ0h0HF28HbQOLLKExzbT+QfvRx0l5aE2blc
ZXSCmjg6triro1q/UlYXKaPY8x55CpK6apdiCOgGqN5qcW2tSSZuoyfZ1u006bVt
rzL+bjyHLeCE3aSntRPussOxB86juI8dHelor7nibg36FVCsw5ayaJhwUqnpq2iU
r+WzQ/vN/o4EN79d6SYvwc/F5xUW+Gi978Y4XrMgXmGhzkcRLkJKG9n3rRv+esdS
EG3KZhEnTHyDrrp9FRBrLqNujM5rLvhlz1YcXI+4gnjJDt1SxZSh4m7l3+x5yqxY
3UfPy94QgWohNaSemWOkFAQKdOgynmTSnMiqt+m8G4RiiJtYFt5+0KWtqnVLiWFq
uWw/AgtzAQvANOpZI+09EXbgdld9ab0QMUZjBNVFDeYjpCWokeLyYEU6lWFqrjU4
yt2CIgCdW1/Z/hfVH8ck4hK4CbFkjkY/LkaMsH6cnjaUmClU529D0k/TFoaqISkI
xZKyI/SNK13ymio7vhYTWVUmbr99SbwWe7l7cGmC5Naq56M0aWvKOZigNR1yqje/
ms06vKpH90uNiMpKCj7bx6ATcxS2Ycnv2JbJOdvVFECPxxwECJBOugaLWW90BTH3
rd/GXboi2x95y5JEdmC46lufEnLm7Y7yMFAmrhjEmd71xBK6DHZU/4KQgrUkorKN
qJZ97eBcaKzcOEabzd8LKpM4aCcPAUtmGDju4zcy7BEnpjx1R/q1b0btMtBJE5zl
ua5uLsge08n6t/1n4scHgBLRNnfAn0Tgk+qbsurP75B8xg43mA1yEXUBQKO/1I4G
VEs0VX8SqrWUORNBxi8icJgukOaEcqU/fe2VOmdBNhF6bZ+deUUbcMFrBGIC51PG
l2aZaP22DeFuCeEuMQuSxW/zYwi56e8qaNxXDjfaOBmOE4F4rhDWVGecdKOEIPNc
D8U8TZaQSGuCcuOrRgcMp00iYHdSdGkuclowohW9TUVzaDY4dP1u3Hvnpj1qq/EO
BCfTHitGALIiDG5b4KzkVqEwcs4SD+tPVMsXEiohU26UJkVlC21JX0MJEOghdf7Y
DjI34+zx+B4HsBgp/GNSt5q8uDIqoyUWUwgwUrOmnxkFvjiDcY9gK4AoCR3IfXnv
E7CM+2ZDO44FLmg+9Ap4zS+DOPBo92UkNLhZQq3kPQ/Wa1DaVCJ5IdgQSIilUYIM
vBBoTqMN8S4gKqar1qygObHSu6u+3u4ByyR1A9ojlhEh5aqmWXtU3joKKs4DsHyg
8EM0kXVHB3yW7W1vhXcKSZ/cB2vArsD0FelhiqtmyGi7y0VrfGvXmC610qivnmt2
8ClQ5pcqrA3+h1RS//wYFdRnCSJ3mIIJER6cHZWJOZrLH3M1y/8JhofSBunDzED/
KZTcI3usrD0gwBhxPH5tA9/OjOH7qDARiQAnZmCwU2YbZlcMT6yhuyFqxOez8r7p
nKLM87wWEt2/OSEAWpdaSfKNhVEAHadh4kq7F0hCxpoHB9qTxyuPfnrD7dlTQT96
UIR7Cd2H4WtqCodcbBQaVBscN8kbsR895blOPGIalyl23e7XeAmZLl2YbsKejyq4
qznTfWaLhkn3jytzYLRKBhW5l/dmXontr0QGnsnajkSSlXnhTgPidrAgZXyIfo4n
vq9hCwP488zyfMZAXTJbEBZLkqKDjAA5b3FVNM5EpDbWsRvRmE5nbMUXzyqA3JIE
1RdMs45JNMjh6hItAwdSGXT2QPV/XEUBuTq5fvtJ2Esc0li9miDnuR71uEF6rPHH
KIHrrQYL+k4qz1GAg/SQT9p/tl3Z5mw8pHHUt66xGHFs1w76Lrc6m06fiKI1Wztp
Y+Y/FvQP0R98Gl4KdHZXwmiTCcmvDH6tspnRRGQ2fmGPIMWNCXLPisgoIZE08EAz
ccuqvc/V1HYc0utOrBpd52pMurExSocdaae2Dba18cK7GHwkmTlteEOcagUjiwEY
9J15o+CyU+gpqZaJfc+0WG5aR1gYbcKAS5tX/u8bJBn6wkignciEsgfEGZbkQrVm
vTjk9EbN1bCxAhq6zW90eMf5t8ahWf2whBEangqHOpVD63gDwldEFYKOCJEQRoVv
kmQtOgmc8be0mhWjYhno23RYpx+yCpBeDOBxZX2ZBzTuDLAFrA/6LiWPx7QvYbQo
LQNVDdVffat6KtagQn4gTdb+eYjRhx6yWVAV+TFWwevb/x4Pw0UKWlIQZIy+zVcy
U7QVsccXKgoXs9N6aOnsR4oaKI2FPQjUVKrxGn5ix1G/2MduxBG9tgx2nwohv2O+
AJpKxwG2TNcYGF1Q8+9LDidmpCptnP9wnBGJuPNoqDBAqSPmpqWoML6kp6uia2zI
agWwOftWgOXDW8KZAccWqmGL7WRMu6/X1YNQlLhY/YOyM+r/kif2K4UQd3aHVMEb
xdE7BxBSMpd/Lv9Cga58RPJuOgz2lag/nal/H4O98MQef7k9SVENGQdi+5iKPm6b
l0VOC9b94dUdAbJFv8MISeTmu++YDDmghD5ot3WhHHONWCW8OuMyVNyigNl+bsD7
diex2Q/HWVaMDgwtrTCB6PyAm/V6kI2czRcygH5wIIDA7JtT8R08SxG4vG6piWOl
eJRfBXK2aWr3TqRNjnFbkuF+A+L/eDvht70rNNnpsvpZPPzxqsv0WMmBxKLcdIsQ
9yrVpzREmQ/bmy326mQp5uaXejmYM0HoUywrB2YIW9mQIbjaxU7mSt85Gv2zgIM8
M4qgMrLfDvCx7L+G+31dY6freRqgsmTajLX6onb06CR/kvgpcST3kf3fc+kSEyIk
+ahJAPo5a8j6BHQNBAu04g+gz/OhfHRQxLh4EUnWEtxSYBOZkbyVpNjAYzGLQ+ta
DIB3mlzTL6VwqFhpdWnLEzvnZDzZvb5UzR/fm5vf2CVba3VIeBdjhWkgVKJgkOw5
wLpsMWGBgucJseO5bmcytiCSthhNiJxRSXiL9uPGD7+WIkMFvpoa+eHnvZAddFy3
cOifWM+U0jZfKiwx5eP5pwojMXeGD3pp2hJbwlh/tFp9+cAG4VxdwGXN5YN5T4O+
ockk9J35ErwY8RDJvr9ia2soSHNAo/L4FRDcuQY6zp+BgMrVAojP41D3V0kyCOGy
xRkAtnQTwFCfg0/oiQfPLw64ORYa6Ena1x0Nm7YjOIlW4Aonkmutifar4mfM4d2P
u9Q5kpEISMLY0JXzUtgWqAcGhbeWbiCrxT3qdro/EUfY7Mz2DZzJfa7KS+mkWM5G
KpgVVLYHlZqTN9r7xFE2XiNZCfKgY5bHf7A9Z54c14xAZzP0n47kKgkNQZjPHayP
azyunnaQ0a93aUT9MIkUEtlN1Eml3G029dMUc7MxqBiQ4YDe7BEuIk2QBE25MS5n
5q8xPZ7zOCQsE7/910qn+vBhMXGtaWYjgPgLd+3kU50mrFI7Hxt0VZCZy5QAf5sM
WJfgJsiYuKSG+IRAvNnLgrmXue41cepM2/9cryAqNu4ltD+BZ4/rCVjBzJd5HpF3
SotNsdrAFaTrpQVWrjRWjAkGxTpRuBlAkJ6ZAmr9YwSa+DVGI4kkCEhxRtIfmTAV
jjrlMYcK6H/89K74tsvRebltnecIVipVSkw/nOWRMdhGzGi9K9yxDpGmZCqyFXQB
JZqLCi3auO0nDnxxfhSYnmIErN/J7yHSa0xZQOmbFLMTj69Wr8WJer/BBEu5Yq0U
+SZjGl4K3o2DOhzR9oZ70jBx4Y8wU18yuLeZhHi3w3Ew52aMf9eUsMXGX6+OD6tf
dxNwcAHwOk6fB6PGSq151eyr/yu+ZGmylWFTdbaAeUevrtcpM6UaxW7FujaAaK6k
wsYSd1PSjPQSSt8xfdqCdvaQCtdOZ9dDzudl4BLkmYVpS8QDgmBGZtJT3QAcwsEU
qSuACyK3bf9nexpQ3rWJH/D+cfkSS904LU+ibR63jEf/LcFr53UU3uqRvVSMhq8R
1MUjs7KOY+MMHkWbPZibsb66mMMHft31KZZ8Y207BtGf8+gzOjbUjFZylV3bOR5o
LASviRItA0fFlrVGksOsxtu6z954R9oOLCkJSJJW78f1a0eceN5vOCptZnLGow5z
hQz4KqL7uYJ2zF5IvuhSh8xiqylK0l3SDsuBxPYHEynU0pI89aQtub82N+a3ZoAW
MolziaFRyissEgweRJbmw+euZAep6PkFMJjosGdwxDKp2QMYGMUcIsmgwNxnC2YQ
/9DX1qZrNfzf6Hoj7XqNiVx1AnYSmJRBEfDk/2YYYSxDiTIvp7Abzli/qnseu/Tv
/p4BxU5YZ2qoJXFs6qO9pir/HanRtASRE1v6aIcQBatLCl2vc/XBhvLqxPNXWSZD
rMbPBcuwy6Z2ZHbxmhPIDabimetTnof5ZXxH59k9HoNGd26UnxUamfXS0it6A5eL
OppAZIqAe8K2naGWGNQkvL+uWw2HYvdoHqA7msF+T6R/E4/PnhzFTpXJp24JwYOL
Jnre6+Y1mPvEGbtf1EzmmhqpyfVHLNP6GMn4v1X4X6fpKY/LsdvdHO4hpbZPhPUd
BOBkfIxtpN7IQfS/dovlx8fThrIJy7TtKxhsCnfVgWurS/PVcsxtme7HgHv2IXA+
/RHg/Bgy/Sz9oiHQrxKaOGwPkQUhXQVFAa1965gGtDtJb3+6K1UOzQ/l41uOXeOO
ZybM7pTdbfYoGpvp4vnRRlxqfVKdH4tPla5HG1FOigeZhu60B12qxto3VkXWCqp7
ErjzN4Q+b2clnAF00nJbfLVTYANbhlQvJHZs0EXK9iWKPjtwSxEv76+x5v0v+g38
5EYy2rbECr+48hWgmttLxqmXvUppMznTBowO6pMwVuacgtcacHQOgps15q/wKfw7
HnSDmft2I3tHAH8kni14dmhC3MTXP/5oHDBjKwC8+E9jTU8gzdTaqSKfn40Hhur6
zysl6NW54+LSvC79MX1h6vcEL/ZOSqasXVvkVfxJdmqA4atIBeSVWFLRAAymFrF/
UJVp0WhnIriGeSiRUMkDlO2ch2FUCCZZZqGPzuiDaXiH3XqxroQMyhQ3yrqZRiqS
vdgns1oNZfTpKIJGy6AKh8kUqv0a/sQwpH7inpxaYzGt0HZt2cnrso6jW7ziMgW8
Q4vVQC9KR1p8wAxPw9DPqdpIhezHKXEYQBBSlTUDn0Pqx2P2AbJSLaNvoKd30z7E
yDJDW9gpdoKqc/TjddSHcJ2THd427rGmVuz10tr3qWKavsJKmT1J8fDvmyFerHfx
2d9oQiMp9VBlUhU4s3wjIuUzlbeF9PeHl2RcYpOt4jQjmW8u39nWrI16b55guYbZ
Xry1sKmwt9898mMr1NWJo3v2ZLqzrWkLcQ+YgRjiH6QXE5Q45dad+a43H2fpLOru
RsXWqNVSGgZkrqGvoCUK0ezOmcM+H2033nE7l0o5TgTKfJnw69gSyTZxqZkvMoof
v33pTqnfqA+I8Ew4TG3dr3k85otcgDPoU7lk9jdZIp2lG7W/ZAAUkxxgQaJK/fia
pPJQmSv0ODEEz7WdsGdvF8xePioMMddktBvrdo9ga5OIWy8MJ7r3r94WXoRnkvna
96xvIMzbeZxJ07KvtkpEZI8G/O7zDhYYG+jZzSkZyFXpZDswgf15Zo/RkP6mDLRs
6UnCqgK29FoHi9Pqj64rNfK/uNR3SQVaurkIDOU41e3DFqbblGf7gqOv1e+0IKto
yS/fKGpC6z9aT7cPOzo0tChg5phNPQoPNe9fDVpGsqHSJuXEQ7mrykcKunv4TZ/t
nHx2f6C6tj3WY84Seot5oLbAXdy2CNhUsbedzHkC2sJhyef/dBPb6DejBOO9aqJG
HPFdasvx775IfaAesShx7HdUWrxWKCslYHt3/b+IbczIvdn6OjDgX3vqZQGY+OeV
CN86zqWUCKN+4Ma3ceYIJJW+Q/V+fmuAXcsu0hmjKlTYtHg8UPTexLJrhJpxOkJ8
0oEHOqY4z0cYW87u/cGIcxdWqfAq39mlPyUZgE954V2TbRjS2I0GQ8QIYxZkxls5
lqrTszaJD13UjkJNIQ+U7WLFbY61lVQbV/e/tVqrpVaK99IntbGPVtuHZ5aJ78hj
Ds0AR8ny81KFaSZv2xqlrf1+QMbjDtrPTlhsPm3ackyZcjisp+YoUCmME48iY+JF
NpKFaVRvD+aIt6uM1PCxqBjeyChuyr7lDsKXM+UBJ0R5dxtrcjYgnzDi90Hcttq3
g+XNfc4neOlTlSM5RQhhzbzv7F0btVJiEeJLJyVUqnbm8S1q4RSjT1Cg1y3DWRRd
CG7ShpgRRhD+IY/KyXxr0P3Bw+9ib+7nd6AaYqh0i6nCcM/fsVM1hKkCurjMlf6Y
97n6yXAhYlhDrPIjnJt1rcT4WTlTyHGKpjtB4wKpTRXCEUZsWyY/O1wFGFMKnYB0
znwy6ROv/ezoaaWkR6VDJa2orR6LFuKw1hkovuCkZKMReNOIKLAaTqbJtiu5IpxQ
CTxEPEY/OqNAX8G9YqmBI3UFYfW2hKVF6nI538sYvZMDyjn+j9qr0++gqjcGBZAL
9kCrU/mYuC3TC3jK1lZYSZtJKmW3FXn7hsWrymcmRTbNukBxl7A/uuqqEl9AcxYE
b/mqXb9olceTaFOxQsYrt7/tFbTCkvoB4whUTy0tKdif9lw5UvQARdb8uCPmKckP
tL5Zou+FutGfOICPIMnq/sNhC8M3bi4VtG3emY8EJEZfhY25YpE+kO1/Wouo4qG9
CeG/nWAZunEpKaTw8m4Eh+qAV544niVBFzOi45X2Wpnx+86CfoVFuZh8AyUj6xTR
cYAypAwYfozd/8T4CTVgEuQkBhr9CQm0suiYTpf7o5gnrtxt8ca6lvYWboRt/Wmf
NP+lfaNejSbl3dp0+tE4oL+rRVqnkFdGIw5VcHbxL9vhvHqGCGkzvKb+GcyUxppg
h3XBSWpjYBJcoCu/QvqIeg0yLzCdQaN4Be5/AGbvtm1K7i4w2IdRG6Q8UTGf2Pv+
1kms9k7qnynxcF9beKroUovYw77NZndZyeYvY313iW3/BAEBu+s/qeOwTVtiFxl7
+QqMenoj2GWtxSW96hcCRkAjTbkgvVvXTsyYKqU8xLPSjKNXJK5yj6ARMPE/HTEx
PifIofKbFV1BY2bkx78qcDzlBZeljpXtmr5pDvbae88Ks33qIdMwuiCPAtLTQqE6
xVH+IvZKL7CnlIK7HOIAlgsxRUL+TEt6vxZqaydai1IAXRNCIa73ZCsQ+a4o7KzE
bsdfpCpFGMxfsyZvCUL4SyLzQEBvXirykIPr9KkpBnDLbCVtCvH2Jdrx6sZfvudB
0R08iNdRjhn/C+yxcNOuCwOAtftORL3Bk0neDsdkKRZ/CXWcOwfBnvXBbY5wQoTT
lPFKF0pqybDiXHO3eMP1/Vjw81CrS5LLOY0pOGJ1jKHCtLkdyZ9P1yh/J5uDX2zI
K39+bA6Grs122M2zrttYiRuFhKjYSjwlMem+/aDNnl+dapQKrKvEEZp3u0oK47Dx
WKReoqlyS0KxnKZrVfrOsD8xO2o96wh6I0mQahPhcg64R/f5BEVv08ZHOtVRdb7B
S2IV1Z1/UwOAaaOV4AUfjlHEXt6hrGA1QaTl59OtDbfjVr1sL+Fy6hVs4kSibj+q
g81d8zUVZH+04PtlUhKZY/poV0YA1iJK6ul6AeLiya7cIc2yjXky0k8fMUqDzxf7
T0ayj7rLfD4VDBIA3AGsG1egnSndHfazVKcd2vqyXPxpMq9AtZqm2c005+xJcR1l
NKSJfb8Op61HoD/IZc2pEWjP+vBeN6LhSqk/iwYZ+h74GDieLB7P8Z/fRLJp8/jz
xA+zQFip20vahws5oLYN9CW0EVFbvZ1jPHCKJEdvue/v6eLJY8QD4GShCkvOY+O2
hzqiWXqmv3InPDyDkkSgrqBp1kepvhzsaImQML4LxU+TmYQug0i2Y73lsIQWMyJm
9SzVlOMF5C45/Q+gnHTsI7hqEl8aZkEEAk/U1+xs2qFnPOb0IFnRVJcWfrRDavSD
ecn4th3wdkzngco6x4Wi1gM+8msXTKLgYuArwksy+nu6ZwyKlt9EmjzYwxfOGwRr
ikwkrIOEJUmy5Q5NNslXLKkuj730o5Xel/1adG1cfnHeGxLt12i9Va2m0g0WULwp
xgyWKdeh/6hwX7W8QDGNBVg1ESP36X2HJIqPjUJiun5DekfEY9MCCLR064jHaUkp
Twli7NlwKqZq9rKfhVwhQq22ZXk/m4ZuMfrFubTRwVfh1v/3SN5fuR9Vy4IYMNe3
JYAu7pdJes0T3pJRjv5f3fRZuZFr4Ss5S9Qp/2EyosrrlBcjhX1tnUE+z13iSbeM
oH2bLJ07YmrC/MK+6cM8EYsIEGHRG7tpxOOAQTbaX0JDTfv974bqOAJTuB8mE8UZ
Y0okfGmXJeAkaOtF0GJP19EdaLWmt+/brQWSBKHRdtA01O9DAks0q3pXndILbFuh
S+wwsWZnDTp/F+HxKLU22hSxmsnQBYDH11dQ/h5cBznDfP59lo67nob/sOjMdb8d
ZgW5WV3g+zMW8oM021Y45HH8PwzuBForL9cuo3+b2+bI+TcHKWhPrMD4KDRVqzdU
0WZvcinORCbWrmsjJrgFUP6RclybnLuyr6t4KCKNOfAhEsdxrfJb8Ai5C1mX2KAf
ulTA1F/MPY2zw84UZOPllHjrOzzeu6VzJJW1kubu2QVTz6QXq+CrYqy2wDv9KNft
yBXZ/gePNgmZ/FfCn42r4kiTnmiN38A4JZWvHTQxHpTvdTZM2cjqRxJhfYIzszg5
/5VkhAM6hSwbYvOtWWHs6qqBisGfGYccpwtXHwGNm0QQWfnU5xi4cQfBS2aoYWIa
yfZDJmEu+x+RYutI09TR3aV+gNQnwDYj7ryGWc557IpfHISWzulZahG/+dw5Z/cZ
9c0RgWUOhDgKZupWdqeYgHGlID+fDnrwb2ys5FCOVOVLSyJLye8Wy2TWTBHIbo1G
iVUNCzbrLhHh+eD+eYiSmwL/yuPgKOfbr093UL2x4phwXRCCWx2kgbl8RhxhW9WT
Z4gdRY7f2CPDfiFF8x7jVmM9qKhxk0Z/r7L+bWp87GJYkzBu2yqZ8JPhMQp2CMU5
coKW+leZPVuVvjyNTgj8TWtXA3raZ3F3da45gEL4MzzNUu/w+wdgQlruDFCe9xzZ
aY3YgZKPIoAKdJDNbYwtcpNyb3E3SKvK9ikFJvljlK7qbXcz4YQAy+bw63yMRNJz
6mnEdUhSp2P+sVH3Mer+TwWrhCMSN7MuLXe5jiPPivlrqlJaLBixymyCJBPt7gl6
htbPIuE07GJIvgNT20FZtefLcS52/0ccT4QxPMihToViGQw//RdMCjcEydnJbTW6
BCbjDXgZSOzpxXPvsSevvpMFPA6KT+Ukm/w8yJJTFiM4t7tjlDi6xADwW0vUbyxy
EtASL+3weV7eLhuV9RT48a1TNIxaVZeSIxkRML4IDUNHCXVo6XMdsACOiZ5HQuKG
5Ys2s6BrdcCTKaLL8s3lkdQnzR/gk86189ysNavjKttaavaHM1myo5lIDjclCVVi
Kr+vA+ze96ck2UUReDOJ9vprvXwLPIR40zot8GbjkKgANefuWB9ABxfdhXsp973e
JvOO3NXtW/pcOqmMrEmRdxmIFLJWW3kBRccWM4hg3z/35YdsnHuuvVCaedaovzLP
cKDll+4XmZC9/kn5Bavpw82v5BvMHnmuzrdfpUVWhEemI4a0L23LqJDQV/vKGtRJ
YD9i8SV4BpDvEErTz1gDO3sXQapTTVILiyfXTtTp0mDmcjfk6cEds7gBGUa8urt7
hkYH3MF4/5Q60pHk8HNj/b6fiDyykdisf2gfccTRHgipl8KKdUz51+gYFl/w9wF/
INs8lboQ6A7SWvy/q3hjHaYiIEVHIAyfhXGqSEr42m3pFukupJmI6M74Kdbb/Fen
CGJyJMGLd2gbgKPvL0OE1YvuyNiJZimsjyNC9pqrste332TX17fs9bVtvkcGi/oJ
ZG6z87Cr4Fg+RTLEuYosYa/180Qleb8JyjHaZK/8rAHqLTWoRYbmtTyc6lCb8eQs
WR3JfGA37JCk/Rn6pMM4Cfzf1BGRmXktQd2RaJYTByY=
`pragma protect end_protected
