// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Ru8V4osoFYcHl3FPp0+dApyFIy7KD1KhK5VzkyEaAra1UjsgBRj6kpKTv/uUdQTxa/8ula8oK1y1
XpyIoiVgCRMd5DervSZLOi3IYcEGuGVLqDJR1qvfTSfl+SS9qt05lgWEBk6EiMu/M+3W6unN7Ksc
YK7Ut6grPfThQR9Lj1cPQ6ohPP9jeCtoS76Yq8hPIQuwmp2BuxgiHh1/78UOFRJgAqEfEVoCxxGx
MPyijHWwNjvGYIcdaMmZkY2agkLTP9hfmA7KI3wlZ86RFhTe7eTE8PrB3AZlRl0uLGiCColzXg6j
qGFo+byfPBQ1qCkIPBQFLaz+zu7bflxr7wmBYw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
E09hkfPXTFjXnfaRNGdu6Fm7OaJBx16i0Xr726Ute1VMAAQJRCleShROAcFLV/sJ/bu5s3G+QEVd
lZi+IcXQLQ8N1CRQ5Gbpoxfv2epxBuvxv9d4CDqU5e7U7PCJPXdhLG/YsiFNxn5ClqQavLu/2RbP
xAkidkZkVvOaOs++q/r6r40rjdVw3PickwrcauHS24xAI6XDCpaQhuWcOMzu8BG8LGqeltFi7zai
XH3HYvBVtbv9VufdfWnMyiOsQQI5bLP8UWHkTvLrjmxK/iGRcjhUJYB2OeK1uEVicm26qDs3chzf
P5uFGdUtKPc6y4GuCI0Wz2eBvg0pXXOLUBxI1SD2U48prcUn7aPuX90PMOABZEzFUbHJch9IVeFf
Ggn1bjuoYe3G2pKV3SYxBWj339cTX/VyxgcPEX8QflH3kTu8noQzF/jKTQ35IP2URTZhwqV1455M
C5TIETwivQhIDZLXEuNGXr3v3fI1rUDP+sSUGnapjjZPLgehFBkajL6q27FbD3HE/+HPNWDGLe0L
qQMze2DHtd8aeJMG4LG+YuYeN+GZpHGVC+nz6Er+ezO2apensV9DfxgXu/YiAT/iBxskwXubkrD+
2bWWjUMQh8kPID1FeZAshhUfGN8AfqLR/t+fZO3POuVRT6cRMvDyWswlH6vKfF+JJF2soVBGXYbW
yuIt3DR9bHhJGQjgSnlI4T/bE6rFPDfSwIInL1cQdwV8Dkbak/Lw2jwacuHuBfvQwwBLUyzYf8tM
dlxDd0fyPu28qFad4D4iJYPQHcC5wpDR1C1dd1TEpUoYkUX5vDcmPenXZZyo6w0ctyDzqspJA+Tj
sfXgVodpVBpRCWNdpy2MJECgWOdvEO3yVLApH8yjN4Bts3Vl7mCT1fKGC2fiCBPV4KObGAZHEBRu
RM122dCf0GIs6mIptLefG13iYCBuu+wedexvtimcNTE93GvyTlAGo6ciC9G8YEUU8ajRapOCuPyi
X0TnBlzJskGVtSWSuaTUVzwcyHe1wW5H5zY24cK9Wy8ooBuhocDa74l1IGfN4yGZdk915/N2UXSl
5buNpu+F1+27Ox+v8W4NbK/vBiY5F7hZpilmOSxifZSTIJE0L2MUC3O7MhTGCy8/Ncjm3F3ORgbe
y5nqhurbbGkJZ/Ac1kox5l1XZQxoZd1breNM9iGGr4OAjcejBbwNXlcDuKQG94VWbe83iNESWleN
1HAC0d5b1wSO4bUrqL31wpdeotYMwKOQ/TN0S+3dYat8oPb+O5rjkFVT9XjW41bXO1n/67WjZZRu
rRrIlF6/DMEZGp+jn1Ne6YYfCJSSKF5peAfFwbjag0v4w73pDNLLjc7rjX3ehMcMPe8YL6LALEV3
Qm+Q1C2sFXynHm1DsEVTbwFAG3b134fAKLQfDKOrJ7woFrhkxVI1JCuu+fbutmrnGYbidc2t1iT3
4q/Ho3YRdcGHJV6bCHLieOqP0oCFOUXPDdzf762ru2MJ122AMM47m+Wt5ed/Kc9+W7qywvu5AwWp
wDSUFptFKdyAhic3Cw+zSeM9RlpnBHXnbaz/mWBy+1+d38ifJekzPc8sOU56pPNYP98/NHqWJp18
iJgTwDxtubFBODFjHrlrYmKrZVu7jkuB895IgLd5zIERpIGvs4FmmYhKvWWUehsn1aWEwPZZ+iPh
NC/dpjm78W0I17qW13/IaAuaZC95CixjulDRJIW4sqxSd+t3deB5ge6/A29WfIhQF4mwovlcUpzy
rZ2sWcryiZJVsxPpwOmVz8t+Q5ubkjvz3UvZ++oy8deB9nZxCeB9nzC5RrmKU3lwDSBVVpACY2zj
xAgmhxKanFmk/ektKyl3iNff93wE6q/wEatw6XK5i7RaHyL2Z+nN1bp145dCy15jUjsnImFBywQc
dY6YR/Ykycr3OV8EhurYQuOlbwZRlvGIjki3nmgHv0iaJzM8CkTvGf2a7A8XIYrJ+60uxlL2YIDv
DOhjFYZ+QCci8RLe7ctAppdzO/Ibhes8gbjhdFTia50ICOZmUckPgGBGLr5Sq9Yzekz/i1OqLfFh
5PzjPBm3jrKM5H/HtO3DCDo8DixeulqeAUxeOZVjd9i+iOvi9AsKL+cin9nMHKXYAWFRt0B40vhB
rAtyrVhXhRCdk7gtdfnvfS1QParRP4WfzuF5QbB2TXqSDdqGh8jy0LWFR5fby+8n2FkPcz2oNCuB
k7VDm7I0xxaamwHZIbNTOs1RtQYfHVco0uQ+8nX/Tv2KK610JuFUFT9NvCUbLC9Mcrv6hG5NoW86
nu6r+EwhRmMkNhPnD744dHyhhZ/jjD7dgSdt+jBa1sXU2NQha3Vs+DGo/VQaYdef9vrS2NSeppHL
ANQtKOSMWU0VpegNNuGusJS0P4nwbippG9IMaB/EeBnpIP6S+cmK61RY29CYGKjO+ifM/XvrqBnT
7ffbhvF6DZxiGgRid4ZRUsfSAl9ZZOG2kD8e82gCz5XFyi2/nBQfPOCJl4NU7Q3gAK9fbtKSFESH
PIL9Oicz52XKwCLG3cOsf3oW+kOHz8ZfKiZipGkc/0UpSfzlwnMAzl4c2x+/UbvizJY0yag7lL72
+TVsZncMvI0K3mjtkf6uuDEh2+u3ky7OjLalxWgf9wjD8Gd2nMIFYc3iAk3yUN6+HVaWZhZtQNKY
vzbZsYT+l2MtYAZV9CmMPT6Dx1o0A34T+vWA11Vq521EUpsiITwSXe5KYbvhIw0Y/oKIqeCC4oTZ
7ZVM4Hh9jtYKN+XpApphw/e8y4EZGsPfNIoMGC4MNPlhZVV45BUg8layVxSZernVN/7QMrJxwkft
9lz2D2WQr2/sdbmSQvRoKaRRGlayVFkIlEwNTmxuJ638EzyX+BBTaNu3Zk3HxFiB3OMVbaVPBd5U
AtJrww8q1YlEWOb25EeS9+4lwbzBZRy9lLlEY4Dyy9XaUX7pEALbChq4Kvm8FyjTVJPbXCF+ba1N
p/VCHG2YSr3E9m0nm6KG3Owg1BbrRNS0Y0hcXinkPBlzsSBoo/q6DYGahZQ+r0t3eXi8ScVN805l
M2t16mAF8xXxvB1aNUkvCJArsBzMtkhMTKaly5IN7BbycbtDnBOU04iOd1wNEHDfOtMB4KwNMAZm
SiYYB5okDQj+SGA2AkfDK6BspunBr6grVWPVLwL1VRL0B88kL7v3lgbs5+ufB4q/QMRHqeI8Q/Os
tTQT5FrvoHssgRBszpwccNR8UX5CXL21V5u3gJzhCH/UVT1KpCofg0Cu9s6N+VP9jVRXCfKSUZ05
xuBZD2De2eAXAHoLT4l7pZLJPXRQjeG3UtR1SBffZ/wccuuRD6sX/tzf1iB/zC+8Nbukzm3Gm9Bd
BmNDtqYlvYXN0GB7iow+esXl3s6k5Bz6Kb4TcX4KHBNbGLF8M/zo5IamzkQP+w9qcLG2N5uEoqqz
+qQ0tPGrODSDngYKCPhB905rjkDyFuiaSijxs9f/MkXbBpFGx42kLn6+9204gqHNd3kqBZkBzUEM
Dqj36tzHtBefJmo3OZTjpwDR/OnnAtlizXFfRIJle+nwDDFD0JqqwsXGU7/ZrG2upmRPoKy95VMV
ewexaCfsWDVwLGRgylKajYPACWA4wYTfnF0Oy9Fz5hxnZHl2zlaLXLftGHUbrfZM13Idck+4bqoq
a7wzSKodbbOpvWQSHHN4P6H6GrqbJYvvUvNBEjYoYhwNrm9n3qJLqb3KLDGDRfximb+vL81ph3BB
e0uzcyvmdYA3zcn+IL7yRGVZPwkBRavibg0tbZJodiGqRblO3zK3gl9Talhc7a9pmP/3KTcCyWPm
ke0GwhoDPfAtCNGSQwjz77qGOGjJUCg2IVREXYX3gDEokIndosNvALF2PVGUXedJHRxwuOsKmrLR
eN1RCXGcbzelPdTIYfPgKITwvtoMArn/NITDAgfjhzQwJiOjA6pa2XDof/687Yf2qr2jT/wWk7Xs
8v8ZMAG8LU2a173JNQRxP5sLp+H6/UzlfyJEIrFqHjHrx6IEYpo44pLH28CmpYHOQzU5v1d3yaQ8
Z9zhbr0zNcU77UA3goGy7L1PBZxuKSPsDhOuQRfgRXio3TsWGzjEN9h6BSw6dyr7gxk6VbtWBePN
5R9JBTgChr9WEsCTfCXIKjLljayNTzoWJLdk8IxDUjNT8dOL4s8QmiyIWemlrwXQAYzvEKrztGRl
v5BSGnGItGr5GHFSgHwvMI1PynTpizfix/zZdbDHkcJq8dPfunUbdYFWqbFSKaeli0Cp3+Cnp5WL
jjPsXkDECvwzCeDU1TWrB8mlsypJ+yrzJvZG36pcZlyoTvtkS3gu/a2Qw3YtvbY/UP1E4zGhwsAM
4XBt/SDVoPgSKM0G2xLXkN/hmSOGiBYq14FgFXeJk83KNP/1afyZIYRLP/H3en+gbHamyndJciTA
uRIoL3l3aqhF+B89xTgWOvIoEU//8TcpLqL3MpBb9tz8ugZD9jV5JbIuiz16RFIohekJZUu9NcFS
3x56nCKfKfjkqLffpzMzb+6j5XTTyRxWMOK81qIcMTLGxynveu8RpzriWYwD+SDpFePFzwBL81DD
u+5ZXl1a7jTbuW9PI0ILQzrpMZd/W6uBMP/OaTlCjvmopQKYUiHjIKsFOIqs++DnAS75kM+ijvfP
7587lQ9Xu3SXktd8Efw5zjvyuoHyWm1uGYviAGqmL5BCHvmuqPF7hChmcN7qixjlwn/ZseY+stEO
Ht0vLuzPh+ur/Y59Y3+HOQBOqZt92Yf1fDan9v0grEREv0lJ7YbEwDk7Ju0MfiVO+NAwr0qoFfsK
1bW37bitCsNyj0pB7tnhJOSQxKZK46KESZOq+dwJYeqMljnTfi5ZnbZvucerrxFas9e6e2n8Sqku
CcPTVZK1AUQmmRVviz0UKsEdwAigam7mxBLaOn71H7r0vN0JVCECNhMqkCVHQelrBWrlSJgcMtfs
DI6wp840ST9dId2l7/z7TuCT4tnCoF9UnkitPnQ6P8u8EWSneodYVjyAp3Y7glVSNS9g6x9qE+Tg
5i7EF4Bu3KjvG0tM9n+ol/NSNym14QOeOnSv61vryqEHvVfJK141GrcMyB5BpNfuSTAafjtZBb/e
wQdEj7f3nb5EpbuS1vX+7sV6M8cPEfofWQJ5hGBpEdHhprY5QHtLBo/252f8V69jA0JODk1oopR6
VnS9nIXwvSdFdWSE9E0ZXEdApw9nkAtze+VvfPkGOYyRnMiPdrDB7zCyk6CuRw0eUTLIEWYRF5qe
oNi4pbDr/jopRtM0tpOdzdCrBkha0ZI2sjOfk2WEV2WUcbw6oNBU4ijgN2KJPUginyqS3CtVY2Yc
3/SUG0sLO10HudbHou56RUMBR+uAxzc2Z9rP7qIrbLzHjSuLpv5LZWu4G/JxLY9i/glLyIhs+aRd
CVyr13RZOIlZTFlUQSJ5PYSbnsRfbVDtjv5XgppAejTeQDrRPGbFicn5Ik3kynRPMBvoFVivfjg9
fKDHb7Cu4lFiM6QwMdA/jb9rm0NHeXhYdyziCmzsu0GjjxGyM56sQM/yCua4jt6i5aY9UU4XAOXc
rC69D/1BMoXc37lqXV+2+a3dm8W1Ge0C2xF/JK4Y9vPx62tWxRGdbOo66PIPov0eFj1mwqKOJ586
GM1F0MzB9bUW9XJ/8ZM0zZNWUUDZy6OWXOoe2wt840NenlTewv8t4999b2vyI1Vo/gXmUhVek9e6
5usZbYJ+r7TwdMLfGspaHLzvEJv8/Sl57IIeNcYh1kKTsq+au4eJn1BI4XZLDqGmAOmYEwqUeojV
d6kyygedXNG6D6CKzdbEuh72byIhOox8oWkG9OWWVQ6wWZt4t2AouniBPmiDDpPctlcSjlRYJAOg
omP0Ll6gdtTyf+Y+aDYm6SysTnndfA/fRHs2+93zJyPjtHfxCJdJWhiUYSPwHKKqXiFmA6BEexFo
jAZTTHW/CLfRuJNVkearWLigqi3jrQ0K1NNUt0V3C+1lmW/o6oVloyDiMsZBC9sbzXbRFd3qoHl6
hdj8H+EKXUVLnZihsfDZnyGjlsRpo4FP0l8dcUZ3YD2YqUduw5yIZEZHWwP6C3DCJsKam0IAyv+9
MbHWASgmYFD5BS42EMoUdmuuOPSMCv/u4m41f8FD65zq0pxZ2sMuKfeUkomrjN1T+UD7JW+HLMN9
ppvF4VJ+uFOW+F9WCRaRIM6Rz0Mkb6M4B32L5zhZqLZOZIa+oMgA+mdVbFEGT60Yk8BNQLB/01NC
xYHFT49zVlWuGillKPCflOpX5hotcXOMRjuvcdQB9LLeyg6EvDs6x2+xSVTjlMsOh53GU/9Tgwhu
rrW/rUZpgi4b2jB35QWvoPYPqigNAlWoywjbugU8t1dB4aqB4+oP4AF/zZEGvO0CZjCCB9LrqF8W
3Nw14Czfv3XDneA0ZpWmtkcmyBu21eyFw+TlE+gU35IVdHFJXqJtFdXAdWLsePy4Ef1lRAI9dqeN
GlMtP/vnim0GEP4WC8Uhyz44XOUtX02fbAB7ngaDgqt5Vs2cpPyut8tzc1PZZx1sMn2GdX3O5PTo
jeo/HE+UBX9OzZxFpldp32O75ffIAZF+oTQqb1rQh7SPAWslXRUt5cVbNV4zgszgFn069/Zt/mfY
SHj0FeMGMl/O1eF8YB65FcBkUe1y2JYyFos3EBYDlYxJQU11lRjB/yPKeCzJjlNEr4RVeKaEZ30s
UpJqGpu2J1OaSGywYOCaSI8At7X2EegzlFfPR/f+7j2Lkg9A7TdhGffExJKvAkcAyuc+zltI1KqX
Bk8BTZ5BLQwdPBAZ93+szrUvNVWZN8MXD+d+AmfxWCPkUEeXRogGf6qa066fXY4+ZIJV/RKH81h5
BPHlvWmDDQswOYnMXDqf91Hh8yRWnlhtyaoLQUi/cARk53+BZf+1XhXg3fT/4gtilI3CtpJt5Ei8
VMZBY5gqM/gpSuEwjjsmxKhSzApX4+oxZU+b7rRFURpUZuvf7o6AfnRfx9r+clGg6W90TKhe5Jrk
lr48aw0gHdcxlCFWTdv3q5FO43f3Ee+Do26Fv/iMXZfmu0HI3PH4flWK+PD2fLzA3NYj70pOjQVF
vA5nhBs/Yl4NoUJcQC0+SFu/I+2GqtCNEJ9AbqloiWERZGZxIwoWUrtw2RHmUimayPRjl9JQbdOF
OS8o82oQC2FOovH3wTBuK37cg9Kto+hqaQ8lfRoRABA3MjhilRec1TZPs8R8G8Otw8Kkp1M5QAgK
sLvyyf67jJAOcjCucPYvyX3UINlcwr9uPChPkEzEmSAxeVJ0XKERlJqXX+qY+cIrFi5qhAVRbncM
jwAhEQnB5eNZwlZx46YcMSzNx4pkFQTFyvXSaCRtGQVpV9C3D8bHDjUyLxM8rc+xTdFPze7It7MA
d1LvrLLkpn6BsUVKkbLTHVMWQdVqCeOeE6JOk/35E9gzMRPMhRhX+DZB/+oBpOPABOe0B618wMtH
wsNSul274DX7XKglgJynJCPkWoQKjtpvsFSozMlfvG4sRHq3pDTzJYMvsfOdDO6Pi+qpmfQVmzSP
52aIi4X5YPwoMQkNPny5ta62mC8Ekw5ehO6P25FNfY04da/78p1TiZ1tIC2rN9vSI7O8+WXAZj9P
ybhtpFpuS48qjuNZzLmd1CiJrmi1SlnUywxx59F93ULucwJ/id9zT5qPnXen87rrvj5W5vdnvVK9
lh7lu3NsDURF/f//+r+fAye3VOY5ZLObR7G0nib5g5jKnFMw7OBCcLMgjJFZeUumfYDPNlkMEFyM
u4zZgpoHnCNE3quf9vMxQdgdzjsWbCa31++mDbvZ3+lFgstVlH34shCwddSl51cFu5CK3qGW+m5Q
xY7+77WwHDcNxI5X3VwM24aHUVGJtrBFO6lJN1y4HSvjFsu1KWbpm3g2HH1ax3kHsSVgcbBkf30U
75PRmuFIo6CCaXfAKo+El6aCpPaAmu4osWMy6jxNIPZkZlm6X0j+cXZFa6Ti6RIDSF8/C1Vt0YvO
KJ+I6L64a38eg46ssazA1O0BkOD6FcXjhu8Mtatzk4Tzwr83DudA/eCG2mewk9dcG6MjOSaLYQ3Z
gzVqZFYHOjibtA+1PKVWvO90LBtHXZ4W+JbZ1A/etQYz9dtkEWsf+JCSa7jnyCxx3FQ62eTOKztM
Leop/n3ba7HZOxdg0jErGoIMxLyT0ncxW7l5mQf95rr4XsTnEHGfKeBUAARbkdDH51Wsp1xcbyP/
f/a/CBhYWfNkwguCD2uv/xFccU9Cusl2fLdbGHf3VnZ8QZUhBd665tqFtaNbOpV3K/9aMiRpErHE
gkX2oDFjj04tAqdGYfGhsZk0jsuj9je848FpQCWo3kgChAds6avR4kTzeSphirSr+M1qjIzb1QS7
jYxnSqWKWRC8GudqS89Y145mCnaddSvrAHkU0Tu88fHxGfQrScWQPOS2rw53WMaunzUTFVoOyFRb
v0BWwt94db1QY/4gFif5WZxCe4eCtmtnxN33R7LTGZzo3/ormFThtgjXN/rjgN+r+/84R8AISXF3
kdbKjy2zeOkoFkAnEtxmJfgPACenWSKFsIPHZ9S0Syfl/MHwD8yy68nf5CwZIIFSElFd3Q7CdnLQ
qBafF9ipgBZX7PLPC0KvSgCrV8xHEau58qs3kiGQXyEXI/2Js5QnP5brLqb9ohjTPHTlDJakougX
65/Kc/aPvqDOfgvwc8COQDXdiiCGUgC8lhvLA/uZWhoxanSJZAe6R62MCxHSJEAMj5WLSDPvMUCu
viJn2VZZJBCOEKqRIrOJEYDmQZT+sVfUPEXzbF28ldF4UdsnfVAaOWfj3SHVvGJ5M1Vz5y1fI4pN
UhpDKVdgFUeH8ycWf/rrNcuc01f6cFVErqdV2IT367As3AHBC7n3Q0niYUsGHLEQR3K36tjQdUKg
6MZBXyHt70HhmtvCZFcrr+/rFGXyJlHv64zup3k06T4wY/iRcMJKyG5qwU1QaYtHj3L+16GpPf+B
jwV60SV+qJleV6uMjAJv5AMh6vnDhy79iUL/08CXXYxwzY0TUspS/XCTuKeeIeOAJRWxeQcyiOp5
+VWpGwV0HHHHrmaOXYIem7Gi4il9tba32GUx4TAphM3wO7tLdZWy2+VeW9tHK9xUL/sN6uVxQkVg
V/D5zCRJEbCuNXsoKKRD79z0GWLF99rwM/PCkNcDM0oEeiPta2i+fhMc0oFnFfaftd8JDYqtjzXk
2Jj7qQ0CQC79J7un0iLdq+gtekXs0ijjo9+f5PyPHS3ABG9K0Zi3gZut6bTRbCdxwAzQ+Vgr/cp3
N1fHf5neWaGkP0EjU6rY77qaagCWKDkPpcPRCmcMZTEuDnlOyaI/SXDC4SJm1A4am/FahPE0Ywgb
3ayMhMPqXjHyox4JNkXwixFBb/DiLqL5tbHQPOwzwCmTjs33RrWs/D41zByDZ6gq10WHpLAF1Uwm
fUCA/pi8nFRaMWHF6rbONfLEc4HnnbC8Q15QwCNs8d0DAydqvAHChBmtjDS+ab/2jmGVeIElfMK2
iD6srxZoEx1W9mHNibbPZnTTTuxBtVwivSge2FXysZCG87SxB+MQfGcJEVKjHUUemKLwkw+D8e/Z
rgszUE1a4SYyH57DzUof6Aaw6ObjTVI+eO2N/QN97WkZJwjXOZV5YXxC9YdyXeWLvtEJ+/eMezeQ
6iAC0WNVNMs2/jt9Qr2r0OXQ4RgJistvgTppg/9wsQ+rTe3n+uul8H3MHQVFYXXy5Es9guNt/75G
pyQOXHLQrbrOX264uMCNmGK/sgiMs4chIpRLuEuoJMdzznomZJWiIZTQHaQExLJzJyH3+IYICcOs
ljXVMPXNlzf552dpXfdsCGEcxPi2Czr/QAGZ/84WRJBzPCAZWe4x+oR3rc7ZpRSUzSrZrVUnr8g+
t3svjLyEyrT0Q6HCGLgK3CWhPUHFDhXLemsVgBUQ4CHEmlGmxUu/xCqluXnP7/0vwi5YmvAMmi01
bGyBAc9GS6TgVEq2tprrHAJD0tr+uU3p2ILA3BY+ynoIccp7snZnGIbTzBTny76/kEDK7SS2xhiI
I7fTPF38aXQnn8rENUu2JA5cTvNeNZ5VsNRzRjtZg+iD26SX5mn6VlALYwC3iGuUcMspD0cRLIr9
7kEG7JizmbglYGegmF8nXraJIUXUpghUNFU7jYLC6L2/bLNqs0BRNtOfS5xEL7Pg9cwsVKPGlCpa
T288WBRI6HyCFTBPhHt3Evu930pJPmNAdkEA/CVf85sQIQmXK9zDPJLvFsqpstb791Fxcgedmifp
KdjkFiure7z1fd3zNErFiqEYras+6y1b6Kw1lFUwF8GwvSsIReZRcIyizvlTN7OgCZ4sJbJde6vm
Fi4WtBIVYHxgV8IKKn1OhdxAG73UZNdRBF2ktTi7P/0ZDd6t5PjfiS2oLSV32npcTrTnXQoz/g6C
rs+23nyahl0WDPm+I42mBC2RQMK9aENwatFfoUFWQYhTgRlc7aBB7+eInO6yyxPJ2FAT7vyErk3e
QgaSUe/x/O0f9AJ/C6KXbF4hg/HbUpeW5j/pOK1h0iGRGwonRDYjD2iz6YM388+UsySpFc4Kokbe
j4FC4Ckeh5I+th4fxUX77HazfE9UEwRdBjY0mBZSJHm2HW3Z1lEajevXbad9V4x5zsbtR+dQv3es
wqw+D0OWQUAAjx/DEI7fzvUgxvo9LZTzMFLbxrWi/6f6b18eM2e3lT+6maFWHLQpUyvjpFsNHABc
jjlOpbH6pLbJzW6XUfEBwcqyAlQvBgTmyQ6m1LT1NLmQb8+bccM34KwXNBibfTtp9iGHWWbQw1sm
BqxVxAhsfkNqBHQ5BARP/FwBjaqEKy7nZezuCvuzb4EF+2jAHOVIbBKeHhudHuW+krZc1L71ZhH8
8rubYlvGeWavq8gPbglogOu7KHGrm80Uep1aiM7T9sQmAf+eBhmiwgQVHgLBIOnekHom5j19ya8k
nZtxoxgzUehPebmbJW2cV7KoiNpEBurWo40Ou6GBkb9W9OiHGi114x8RLMRujc6w1OaYCFH2pBqu
+Y4yj26UKi5H8HUw20e4iVv1fdb8p8UC/bPeUpLLtifNZxs2UvsuoVKn6KHy34HzqCxKikv3YJ19
QV2gQiWildXs4kmrS1Rx/PasxQ3QtdguIMHkO136a2e31gahAxAA57T3V4HjNzmyZD5PFLp5nF3L
I8lQy2+iuJSc3jwiWQHmvtQRd41lRKngQ5ssZpoc6AqFO26lOm1jTRCgHTdy/doWNo1Z/Jl1cL6P
UKHugyecys75Gfe+3cBY2oBD3dXDc6JLja7RFyiDu2c58cBPSs43UWDZydJkeGecDBOwknG5QCel
Ym3+e3Nmnce+b9IErSn6sGOi84esA1Cnyd47W0Fucue1fOw/Ky3W5/pg/BAis+/1XPhGN/pyMSge
NO7EUKKDgB0tsZ7/kAQbaqmqwwz59HiYbmkCd3e21EsaWL6+JXvdmo9te3splFNYTWvyDMWuCnMS
fcRiSqRoTGBq04QSpRvpMTwLbVsFQa6hEZISXJMQowfaoJApY/1BLRQp64tg2MvWdFR8W2ntSJJm
NHhjpFqXTdHGHLviBXfY86AXMzxtt6brHzufFu7r1lE7QKzmQdoSdOBZx8vuRWTnWHYxE1hMMGwo
LYJZEM00Hx2oC8TzTTq8ZxZ11bYQVlH3npdjsOwAS7SODJ3+ve2W9W9c6PUVNVIPsvYlTyyFhhdr
JNLkhTPcdc1cn2hWM+SbrG9iGOMPLzBI9kmwOEbxfxz+4AZEv7/vQh7rnyIyoWdTATRPVF3cMEAU
wOqriYecCzflTV5PgfxRdtrAw+bsOad9QdEDYN4yszUPKPbLRvAiCKO/JjSzoCfLwnhPzNtaNjFg
HFNqXxS5nkriMN3lT409PV7x9le4Oq+qOaz6e4kQv2ruEb053XulB6visH4LqG30FpEOG9u4Rop6
rMZjKS5zblE4cq7auBpQyrfKQdM4HnJKBKq38hl5mcLedZspu5jv/3zKkPJc5wvmQtgdi9rC2j4L
AS7S+ogBO8yIc4zoFI0Agj0LdZWnO/d+ko71mTBteT8BXKpNw/0m4ERSnruhUDLqoPVKtEpK6H3e
6lxcGo5bQOPlwrVyhkJhXmU9wkGWun/n3obdTP72IOldfOar8aneZHbuQfXmo0cqd3EiD2ZlgPoY
sRcXszr2Jt1Ell5mnsNC9pojOV4zijB47xUEz3rv+92t/C0HqDLgFXm0CeQ7FJRYG9cN6Xm9lw3n
4USayZtDo7MHpa63S5UYJn0ZXO7dF6/rnkN0bwXwBuLdWpu6WKC9BxjAxumz++bpAFHwk3qfjb8x
tKvvnuXYLpmCpP0gLAGsJYXMlYHFjpuGtwhY67z64hSqP5QfvKu5JpkbNXIU3qlxRem9ZmdPfByi
n6uUtnyntkG8PsXFTVIknpFlfGEVRtRpW4unP4uQ9H5YxST5up+F4SEFBcOiMY1nl3rT724yFfm+
GK2z06DJ7BGN1XGTtqvV9aYMTqu/dfkH8Q6fR5c42jwzf1wC7ZWc2IMhMBv7WMziw+LrpfC665pT
hQUmbVFM/t9esQ9wVAWWtlcPSm8FRrIWXDNr9tpltbHiqjLMCMznZSIhhmq+35uIOB6sxSli0Evz
QyBEvaajvwt6fZIAwv1NREsFtwRTaawYYuaoWHBrU2nVt6xJMq1wFV6KGwoQ4lGyRoVeDreZn8ot
QhYqIFFUcPIIYRiOyVyQFfG5+2VbYMsEV5b1gytDZzPEmfGMGTCfZFC+r0nI/wn3eCElVrKkJ41b
s9Zz/H1hlEvloavSAZFm6WzLRnPd7YZPDVVpJxPTi1Ls/5K8zU6qmMGO5azS+vfPvWtX4lMLqTJg
T1s4Tfd04sN0ynrUJltf2DA+pAs/Fk7xH/Cc6LwTlumP2BXq6uADBxLNeGKtIBTBl5k8gIl+yWKq
RCbJtGMVqLyh/JjLhcMWUo5o+kyVgeVsSuk2T0Ie6xQjC4rsk2oIw1S5ymn9TeUawzvKiW3IkMVR
rqTjDJECqHX4GHvOMEWpVn6ciOpIzaP6dEbVUHv2ME/GjYqUt/1/rGqMD9bppeK6oUd3fvqzLzZn
/Q+COgkhe4irzvw0gRO0ZDRfvTZHgoUmTnxVAerGf6kYwF197rskBijANdDO6PUpWCtmU2WQazSS
/+Sd2B7EFypJFueAixnVyn6o/7Zk7FHdxR/SMG7pOiWnulaQqq2BLyiyIhDQI3KqXSRv3q+deu9o
Lq0NPL8V2VGnL3fgUMByLXMkXDyrnT/U7TL3qrYGSfg39yoKzzbj/xOIVTXeZ4hD9BnHXBsxJHpq
LFRIDCMu1z6yUJRF3+Y68A7vyf/DvAO/zmvZHBQZZL/juNfSyxCFgFzM7YS/WRbWKBMDh2J7TlmX
yFdlFpJ6Q/vwFbvipiSI10xRKAVqooZj9aPpfM5aIZVNTN/G7hg9eHjx+1WIsdtPy+/E5wMRfneN
j65nh9lM4uJfzWxc/SBErzEE7dU2mtIS3PghmNs/FG7JFjH3yPEiT2cZ4yyoJzGzMGemgHI9+1KH
Zb0z8oHd6nnXD53oobZxxPSZgbFGsPxyIiBtz4pxwY8R4VnkKxpzqa7tcc4flYEV0VExoh1dDNBE
awfTcbFp8XHwjjkXYCqIGt+TWxO3BGTfquZ09Dfh7HjNHiH6hlS/LHsT7bIxEOd+qHDsjIlrLjDA
BlzYjm7pz18SRmVfJXYQFzlXpR9CDfP3YP44IztPX8pR0CYL15d6fe8qgb2mWohJyxLf+VeMY6CU
l0zAoT2gk+PRoKClfLRgFCPVYjAVaksfoM+sl565uS42t+grph4YBrzW02iPn4Kaa8RjGoY2au7b
sAkTa+eADaiDbQW3wO7GHBuJKKvWPbsuHH28pKBo27OQJJGNnmez308FhC1p9cMlwkJ6gGOPMMgo
26MBYUFRvkeC+AXz03Ac6fSIrPfWHKo5zb2aY7RXT+AgDxOabJMqeSWM0nRTcuEunmHB6Q0mN/97
B+m8yQMhQ7WMTG8Nkb0Jwt/3qE7gGT3PBqEYVbajjFxj/EuE6/etclYoANWw6wVopfG7/PxL31Id
KmX4W78rHw/wUjlFAC2U1I/t8Xc/dzFMfLgRCMEObBJRWyZjqJi4q+G3zK9rZIv26TjGNtcyzUMJ
dDT5hgOqLuWwFDewjDWRou3Zf7W7ET8GSpHXmumoc+xnqnsq+uXBTl0OwbBoLvUXzzUBGQ99yh8q
4ajE69uBSH/ZqJmFRckXwLCQAj3cx56p3Kk6VKvNaOzb9o4sMK1TZihyJdEhZtaUFDw2lRTePoDV
xgNz176DNaQM4PT0fVkbCpH1P5EssA/Xwsc582QR8AgnjW7Q5gVM5v6U/RXUudY78+J+JLy+2Ljr
bJ+qr/ZhfsXBOhmn6dqG98jH6m37fUNY0PGrQOqvwYZvgKP9WCn6JUEiqRYr3urqRC3NHSfYwtOG
1/sC8oAc+F+4/BxJS9GvrAZtTAFZXL1hEf3zkbuGEJXhHkbusDDlT6q42T65BBvBDI/zBFf7aEXa
uZoa0wnuvR3mNL3tn8NdnnyPgX1DEkmWSS5FanymLPIa/D8V3ZQx+mWYySkJBmBTDsTZs/eu8eOR
X4jntL3MNFpkvHt7eAp/P66FV9tICnNh3l1czHkJ4WET3Rlx+6Uck/+Piwwmh9VHzr0O8+sIz/S1
OlJeoevW6cX/gSrll4rVbWgDv9ykVAXslpEfwmR74ZF4Znshs4C/pfWMtH1xwwJyK9hZDvWT+45u
FhYpnAC/KWwQ0h4euamtHJrf51+SkAfZzFPC3+Nlh1E04KCo0fZkfNlwXnrkSVHs9bqDVmn+CU9t
hQihdbQCoYx4WXz+6FOJKwM2xoHXh99eG9HLhU0yGkiKvZN3Gx7R1qqlv0r2ggaRLmr6Exjaa1Xg
DE80aSNsvT23J3kx95+CcA85opGSwBgErGd2YZbXwNbkAIctZWJsIdQW6E/ct0aCSlXXTq+XBRnT
DIxM4iE7vtDCNX36wvwoaGR8CZjDqWREZLY7jS14yw4Rpvu2VYFSIcBtKH9mMYon+nIRbFyWmnjN
KzymH4IxYMg69A2eFT5rNyDNQzRj+Ts9Z5/cWXAdS+7X6OesPP0vO0hlHzRUU3Mcbu2cCLSJsfjb
jiff4n8zhVzACBLBjorZnueNY7air5XwNsdGkztL0fW2/NXNWsLiBdkVqaO0r+tXyM7niiRcocS4
dFRqSF7OSppPvRGOv2XFuGCYnCs4dlZCzpKkT5uTVHHHAKQD/D7Z5fxUwTTMM/fuOjAauAUoDuo3
vEdWstwrvWPk5F9jNRBKIHbfuyz9NyE8TikZ6YMBtqeQXDEuJpllUPhJ73DVEoESB29hM+zIYYOd
hhS5Z0B7NCCzacdYUduCJwVfrXChO+j6cy84TEjlCGpPbnLRpOg7AkoWZSqvfeoDVlSd0hQX+zdf
6IFfjJQNhQqoGU8keJyec+38ItMwuSa7a3mBRK3ChQk8EkDbWZDNZFXPaNYrJkjGdt1mGgAJm0ij
YmHz/OG3uKu+NJdzFsYN9ErQ9rP593RSclTfZXd4/VfKfSVx8dLVD9S6OSt59zmSR3pDIR6u33Kl
RsxIOCglxLbnVESMXp0x1YEpXsp05PbXMCxO/FiOMwQgWiUegPnkfdT7jScWGfFq1GnNbQViDOWw
q440pZXiD9nk9tsuAv3DJWt7I8u4gED5TlRSfsut/klV3x0mzvnsgmadszdQKRERTbON60YIcuZX
7ioX6JediZIxI/labrqHpNhStmDux9wQAiEIXXTrl35EkIN8xnuvcYPh6OYB3pMMNOWy6ix0ivDu
pAYNLUTl4zA74Gfo53QUmS65D1B1hsoGf82u3QAr4ICdDUCrfdBwfEHhPKw5w9v4NV/kTRFCbRNc
6s+OFZYWOmRPVOM6kAp2zKXr7PwTFZGVSl3/m+UyUeQh1ns30idnquI6vuof/H72DWbwU6e+PcXV
f7BbLUaU1TwVao6B+GkPJtVwwI+1NHktUqRKts2K+ZThs2DyyXycgfB+jUfR94MUqx9LCGOMRgPL
WY424ElJaGiYm2Cfzgf17B88JOFzTHeu1XX1GBy/EWi0GPMKK0Amr2SQCz5UdoAFU0k4QYexx1o0
CdI3j83zmQkO7+FpSf+KyokbuANWRAno686Po2BwCf5gnWCK0MCed8c+T6/VrglAdBxWIc8NMBmn
x9O40dwK0Yz4McTyMfJkOlHu5fCkCsu7wjETnm3KgUiIHcPkxn9gbeIhVIAiN0eN4HnGolHSYrWQ
zKuvdgwiVXwCUMOnFliNIqkqohpU64IVzkJ9olt46TbsNGAh4wzQwQCws6z7Z4wXFBfgLYE5JkT3
T920MsNXwpfDq0+3I/j0OOEt76LgB/IGUdTJTDkQVywWULMIvOn5L3EUp1SYNMo4B/fD/MYKSG0j
E1JUSudHxghj0d2oCGkniEiN66kmn5dqwt9JCNtxdoXmcOI4ylHDzROKsGR86P9liPutWll5opWt
nhPEgMyT3vXhWX0CUmqHxn8HH+EXWI5uhsOOTi29upAvNTCOLAHOeRHXlA8IwdnMTcx/L1FO3Bgq
VPX8TrBLyi1Ua3VtLs30ejXJGK1XmIsyM4fAFe6eBl5bxbx1ca/TwjzA+5N0/37U8hNSqggm8t/T
tgp7lS0biO5MAU2gl6VxkSzU/8W8ZmPpf2GGrYMzzv9e+5rlhoDp5Aay4vOHHW2PJsu1jnK8KOgS
CDfldqxLSkOGtcU06Uix1Rpdi+kz0D2bsYJUacXMkFSDUFOQavelsmBGGV6sUm8eRxQSi0luD/ys
B9fKO71u22u+vU7+XPhql/OU7bDOW3znGwXwRy63uxhnv7mzKIK2k0Bn+RYZpj+xtRE2uuWLGJ6m
if5HPo74+xGxOTIxLXz72fm512wGRGp+b2NEcSGhXYdyv7gm7vBh+TFHV6rP3Jv1nbbuGjXVBaXC
c1vnN97P7edzrsXQbYyANQMVRgKaBbmNMA7rukewzC0v3rYtsxo74ipFlBnrVqajgqcaQLPSurhI
QCF6ftsdzRtoVArmcXd943XT1qGL4uNVozJ17odG6K5psda7hF9bCHZPDfsiy3YCX1XDx6dUNklJ
oTyOje+cMkCo/MdQqmNTnUIshF58fpL5LmFJ1PA8UAZ8H3aPfy0NiyVJJ6qUVlKDcUhTqzJxMB7U
ndV3c/D65wOLWerEKvZDUVY+4T4iocgJ1xsv30unv00wfCYCAviKVi2lXnU9nXO8/Adeyp7FnTbM
0QAz44LY/DrpEpSEDeAPE7sdJ6b9xEq1IgMe4XzTjc2Nq5bE3P7vN/gyzEUrF0rJsqOiaifqqbpp
L/otOJlYH6fUNng2lhW7KHaf8Yknuo782mA/aF6wdog/tBFXkQ9HksqLC610Fla2GBlMlCdk/3RS
JSAowNAe6M1jf/BEDy5Xq7eX4JwDVuIBOvshq0MOmrGMQnql8rSjpFi4VsKlXCnjDVA+MRwkjCqB
WoIh0/XBFeXJTqXgQSHeDnpEDwJAfuQZqSYhOzAxjwHHCmHWgkgjU1AuUo0zDJ/YiqKryZRd97T7
QTG7Oq7rKCnnV4LGYxX2UQgEJddMrO/AKMwCUrmM5aiH7QLoP2c8XaGAFVRnng68+L/Lk77qXCjz
3BrMt/S9mc82f5q051aJhPE1QMNDXIN5L1NGAZOUW7Wllnjn5Aqm46Q2aY1hlw4rV+ombHAp1byS
buBQutFS9wm4F6MnBhwKgRKaV6ImLNFDxE4YV2sQzLGwNZ1PrAusDhrfXqDj+ecMZtXxOA59z2KB
b3k08/iUwywjXWJWL9EIoD82w1F8cFr/uy4+qDpXbU75uwpj79yZrxeGXfkV96u9cYLX/cG+9/rN
DhNRAp4L8VhMs5RXBHSKXwaN7KB0vzCP7IH0SJP2Gqp4skIwwOExNYIPOfhY2cKdCCVDytMq+ojV
K8Ud0vSTgnnvoeieuNV4u45uon36IyNWqCOhj56DZqXLr6v8/6Ohlk/LT4CvNYCZA4fGiOEna+iO
69LNLVag9TTZx3d31vi7RIs0lcYBpSKKF9Ze1xSp3K9DNjafTW95NhMv2vIukykstIMiDYCaB5Nh
WSkSH+phmI1vJsYyh54ZGmxkN8FPQqqVFyOEQ7Eo7J6JbYGaQ0I+NwDOKY3FqQFRXyygjg6hdWBZ
Ckci4kmPdL0J2u28UpZY7HjbAvbVFosPMTGJwj4T5kbeHHfNE2E++szjb9fNCbS94TgNiM6220C5
Yvy+TbdbYPuWSWtSCzMvlEdRLGULSjSKIvOuOPWu5K5QzCoidL1GYp7ugZQ/m3mwJ8GESRcNYUUv
g47n1JYiMPu1j5j8mcomQvXSPzbfGRCPlvEPP981IMLcYx9jR5zGFQQGoK/liavCumeDuxNsxB/h
V88VQ4TGe/SlSEnhGeS5dIYvkss4AWWX2YzCA7lPrSFbKqYjddDNE2gd4B+kXQl45TGBEkXZ6isq
I170dzBZv0gNlCqNiosvTmkAx1J5QyuAl9YDMZEgmhRivh3mqgMMxJO2fXoc1TiLf+HoWsA0Fvbq
QTr0illJi6J01JimkYUGQZ1Z4NJFAXpjaWaHjNSgzPGhWFDmmNwXzVNoObIOTV486mtaIztjt4T8
a8/Izaeb6B+5aTPmuyohlYlFYmzzgsfhltwC65Ld6JlAvTOoGsnxinBR3fw6bFnvokac5Xllt3yQ
UThU9UuP3lKXLP12O4Dh0ThM3rruH4M/zfuQbd0yUktyUZioB/0Ek2irqiD0H5bgEhgdeS5ccitT
4jFidQYuaHZIBqkMXU+JsIsFJPULj48FemeqB6nM2IIfG6ProPTyfqnbtsMgKrLAmFudFtDk4xnR
PcVkZe9WjCEs1Fqe4smlu7MdxCtOTtSRtHYTs0UGra7eLrtmJMibulBX8g2LFQBKWIg72gEU68wO
PudvnLKRObI3dJUzgFaoRKDsT2XpZ+PwoU4ugn9MHngvgJzpVSJx51c2MxNRCxntHGXb9w6WMv/y
X2TaGlzU12QWdxnSS53dmylrJaksBGexwUaOFUHFC0Yk53oL2j0xuQVOqZMCucNpdzNFSM4Fh4/W
okxrgc62lNhQ00bW2F69BaUcpizdgA5P97j4xFLfxCFaLHnKf2pvSmCUCeR6vDCqMMCaf9G8uD5l
zbcYkGbqA9lP3/bH6zemQJ0kIeBeTXRvBdAMZhFGdxaW6Rq9G/Yoa578L/SpRaWFhfTeT27rrdeZ
sNOTSk8+NZ4AI0et5bpQqqz5eoGPxt95hZADCGF4CqBPrWU1g/+NEAANb++W6I5y57Azv5msgw3Y
S1iq5mVy5seIGdW/vDRxVFeXZlIzEjfoI55i57P47HndWi0FkY+g2kA8JHCoSIgV7SL0mMYFXUkL
buiqi3lsZzioQU5c/g00QqD1ay0dDTtX8ffBVVDZ6EB5DadRj2pj/5FXvkliiTcAJCdQwKz7otls
/X22Y1r5pNnGjJAGFdcr+8DfvVxBWZ2R7XaXeDmfaUQE7uMApd2QfaVYKYLq4tEMthxaOwoJ15vO
kcrqd9bgIlZ4h0tFEWlR30hrGg9ZXbVoOsN4Tk1Kte+oYa8hi21G+9qhkRcUgXgAi0BJNauToPZA
R8nIGS1oim7o1anFSLtHLFOcYXlTNDHlJf405tiCYTIMkHb8mTl0DqIU2mKZoBYegcfhh8vDhmFR
5KGr7VTHsFT6Xn9jKmiz1O0j/LY6vn5lqxgk3DEQuNG5P63yGGOTXT20pU8azOASfsRGoA//6AYG
5pbvjdZeSR8Q4iWCL+xH+X5kYwCF4FCbQm08Vu31jXYQtjZaF4sVN6Vk+hRC4gTQ6zGa9oMEpA91
azu+VfbjFzgM61iYDw9PvYrFVQxedtZH86r4UhbKohaN+YSeAYOibmviHLrFNI7ui81etm4/5QkJ
zIV8pUAAtT+qFHgl5B/xd5Y2pPlatCcFp5BREY43mzUQT1lOfSQH6hBqmy3uAy8zM5byAOoxsu2P
YbySOhBaFJgFES3N4tOc6uY=
`pragma protect end_protected
