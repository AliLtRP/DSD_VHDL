// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YULvE152c2wEo2z+iNd+NQe1fxYFOxF1AhyuuVSwqYjBG35zxhLpmFgUw6tkyfR0
7ZuW28Bz780VOdWfwqCbw1Z8+9k/mnak7idTAEx33WIU6syt0h06Lai3K5ncmvnv
YOm3bOkxS/9wD7brZdcysdVthkYOYzXE2208ZWtPiI8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
jKPkgt0a49QhlyclQSxVHU8xtB7Qyk9ya3Itb0AYAjt5jHxiI369Ruk/785BFW6/
wStVKfz02CZp2aAe2yh2c6oZsqSYmbOkNy8X6oQ9AFUzitYvzSpW34YH6DNsPB/y
Tjc23VuVO5YybDgSM7u+DNJ/Wk/tIIdmDXnHMJig74xwMEVAvzeZhtiQ+AlnJ4Qx
V8KgeawQjykWSLxQfNSGXBOiL7i+tL51Cp6o4eNNX0Xy+PclYYext85U+Uk4mEZ4
ZNRAbCCFuR0jqWIa3qSXDkxpCQ4uwLvaJ79rhtgSnxhRV9MboN1dQaztigwV9KIl
ZeGAdGu1rTaHaddbz5QKnHUL+aGkw2IybyzX7AvzIAEVftHxY8qix8VuvPov5d7j
DbanNTNlJ3/qVvsuvmicnFsffQ9BfRCkDy3JZXQqQWgnPW9wT6aYTJTXV3s3L06I
EivImvJiw1//wSk1YeJFwJBcA2sI01iruHyN+5AKNUBA4ssQ+c1DDYB4X51G/eIe
9spBi6LUTaX4Ga8njejFwwGiRXT8WF6FwQrG2Iz+SX0tkE8oBeDVsAYAA0SNIIXh
tdISauDFd0VNZfLMG1Vb2GFoc0Ydr8AaHn+Qbtq28Ywo+RNVkEOXEZwCcmBzhEXn
uwgVA5yeFN4YMKto0otPlmHIyHR4804nm5kfvSJQfirmwTQSwZvuRg01+lg5Gvu5
4uRE+EhZAUXVPYcAQz7VbE5oJKb7odPYpU8eaWjM5aAYj9418Rg28e19D5LwFvaT
scfJBAlw5KEafEe8oVJ2MXIimDfeEi5uP7lwWNajUiNQuIHm6WO0Zb+tdlftuawR
W4EOFWRTH5d5tB0kmcWSpnNUy79V5nOb1XMAGD1ngbJJk9yxtOZWyVZkrTyCVaXO
yBts43uj8wNIRW6ZtMFIUPfqKqTPm2RYBouRmz1oGacFkGJI9X+GTavJvXP8jxmy
LvWYBkhQnPOnTb0I1LD3AhgKSdEXQ4xTzACpbtV3y6ldJL0f0p+//I61ob9+4O1J
FDL0ozrTLEne85a7h78yG5KwetZbQmxVnupM+YSS6T+PCp01aYRgcBGeWvfmWKFK
uyNwLV54ToPiHV7/U6Xf13JEmiqrYoNc2E23Vt7AHgFPuTTMyFV8jw2esr82exp1
io9NvmmbboHuwdqI4CWT8aybLc7OG7iz7pgqUNeq956lo4IXECUyKDpZuC5CBfgW
iSdiwKMy3lAEEv9tRoynHhpPCcCmH582xEWdmXmkC1qEl3XduDDLV9LDUTXSGPDc
5fYrhvLQYL5eSaJVJVGFOfcqNoOLpELpC34QucPdDkd+yqI/6t3w4jkLPJnFsZlG
aPPzPzJu8aL38Pjs0hOe5Uj1x0SW3a0qCkcDxfeic8cHJOg4XWNWrhodGOAUD17d
q9MObG1urk9/SHdLtHsWNRQMIVtoyUedUFe2bf0MvJ+Yfca3GnkwEXkyEHtRaz5f
2vGHogJVG3qX3CiMp4Fmv0hthqyZTbMh4M4pSuI2ImXwtTQk67V6PFAp4+ucVtPW
BiGdRzUQsZlbThR82BZhYdFRswmnwoGRnz/ragXM5pGi/uL+M5Fj62Wqfq3/Ybu2
m3ziutCKDy1p7P+2aJMBEBWK+mkLSqWZ3nQLpxVrV1S5AiXDfj4YrWECf7ZB8RiO
V+XrhLGYXRYlbrPPWc3B77iotpqOXSMVLvSMZePNTQUxQbuco23Yak+1JPKg2Idp
thd0+QSsSmpuq1CQJFFEfgVE7FlW9OtYj6H3s83zCnAsKkX1Zxh6kjfGNelN6N/L
DpOBUb0bjJBaAt9qxRpZlTrX1stye77P2xaw7sNduHg5bp6FNl2RrsSD9ZkKkuv9
SYHjNym2I7f4X1s9MzuZWpJoloMTJAX+PziE0dvghFoISXXuFY1UGoyn9plgxJ45
ZDMXUu/xKktyo+C9U1vH7ShibIqbHks2TA8R4LShjgFixsVLUKHTJxPY7tewmcpI
RBpSxRstTs5fWwEYpOJJvsaH8cieux7umD3+UPpEZXaoreHxDmKwSmOCT97LWsf0
AJFcFaaFmT5K4C0lsVFdJ5Rekw+2m3c802sgfq1pMNPfZq/heX/Bv5QZO6cGObgo
4dyRR2BwP5CLpML5myX3gJjRojbejsIrdfGpS0psUes3B8KtoCwIQULTXHsQqX1y
ODsGa4xo7O8HD1jz9Mt9+iSlRIN8EtmxRj3bxVdGtfU2ofz53jt27brusBozuIvc
g4Vsr5o9fv4hPPZPSxd9ZKucV3vo4vwaj5PPyQ4eKeU2nxOSo2dH7sxToGj1LeBe
gTHJMH34a57VkEIteM6ZRCNDhwp0vpoxK3xTyNyvDyB/oIbFwvTlCNZ07A6zY2xE
qZKgscON2GDpSn4HOIAbwVONfLxMChhDFVoQ2r2JhWl9AUVBk60RWC4uhpJm/lEu
45zCYJ4pfzoEQpe4gnR4+irkQkakpTYe6a152syJtXzcIhtv6JFMMPaxWly4x12a
OEuZLiPKSU5j9lb6NCc9NPDMwPED58u9taAJncVuEjP36xl5BAoluPEAjrXduLCq
dJ/nQPcyUsNPjyr5PmOo7Y7otFxTQ66niEuPscOFq6VO/+JOHZIHmp0aC5YXHbm/
UDJUqjDlwGF34Mu290MitZ1xXaoq3S32cZeju070SJG1nc+hafLlORF5Bu52Offd
2wOqHgMuwBWCoRxx79fIgzdTu8PIYdnf4P+cBKLrVRe7nYm8J5nPLTJ2VS+PSasc
LCt2nS7+OxYN4HESkqSnvP/sz23yAUU3YtKj86lzZYDtJfc0MyXgUy3GH9fsePQW
muoVObbNG4mesBmpMQTTylpO88Glf2LDQr72aQ2ziFkdZXhlzIS/zPWBGI9RFa6g
rUT9VwFIjQVjgOdnNzpA2uKwOJvo/PYh9yqYbxiNBZqz8pu1wNSKPyNmN3mge5yu
1hzOrXgCYzeZDHuRZEzzK755HS9JGgeKk33nf+Iu3Ilq7mHa24YIETcsxdI18BDO
6tX0g1n2hS0hFD0Eh3wQjo//VR3v/jZeqrSTpQTmZoSLGqvBKWEAUQJ8VfevaycG
ag2+EYvM0kTrZH2oi7mzKvmTDfIGn7YQOzOpMATCpWuHxmnKVJMjViWIWjIAHy+H
adbf0aTphY0OkcyX6bu7Lr42raIYra90riw3Na6A5c8jDlujpgwWV9j/p3p4Pbi4
pJ4G1HStZPJ+vW11iB1eb4Pld/+PzM9fcFywBSjdTNQorXKfNVU1DnOqWL1JAjeh
HJuz+f0QVZEfdkDbHjXLP1pPygkgIoUpdGbugfzvPYf//BFRU6p6n/XJfAW1vciz
y1A6BDoOUAQI1HATcTPqkN96HAezPyOOuWjy3J4qPgjYXk9p9nkovvSEfmMMhEK1
P3pqnQroIHJoxBejO0qd7pSXUO2FCDL/Myny33moJR0RijFoNVDEC9gGCytnoeqc
o9b7brVJwr5NcG1L9Nj+fH6i2bCbtkdMcF2BtorXWIKVvsPzYzlKG3U4gnh5JSGi
68Dz3s9LwqugimEDkSe8DC4bH5YINpRpivCDiyv+uZ7GfLjUPWPBHwEQXtP+tzDB
no3Di32EEGS5hCgT+lfRu4QYxmLWIHLvhxC8ENym+272vZ/FZhRxQQlgmaTrXM5W
qSo6Ojpwecx7+EnWaVqrel1l2bZCoADHBNeKcpUZtBxOdz6pcJ2HVrc0oxEAZqhG
mb0NEY64Irr8EocgYuKTGhCt3c7cYI5ZNvEaHPm+Tyr1B7fcIIWmWW+kvN9VmhB2
cnT24HLbvhYFxBixXUhKfMUN94YnCuVMFtUF1eteQZDJRC/Wr76mHd+oYHQsofG/
NPl7r+s8vD4GxW+9NzJp5pWlwVujzdt6d5pAlwYIroLyg+ZIyN+uEuCo1etF0p7t
GbydUjRKZITJRExiU5mdVj32q93WKFHw/lAW+Bow6y+cLNHxTqy7Niayq9WUjyXC
IZPGua+XBj6DhE+PEztmlA1fX04J8wm8AKrUApA9OSyV5MwoxepzuzNo37Jdpagr
h0X4Jj1UDntFtJYgt0gN9LMAHXxVYNdtN6DN8uRG0qLSsOxzx/4GJX3MDA9JNsVA
t4iALm2wKqS3VuyTnHW8W6ScZYIgUNEWIbWnVc9vIYt2taf+BxcV/uzZogtDJhub
86Ha9c3jJfa51z8NpBJaHwcdalRt0TOt5cX0K48DOGLV4P5Kuo0TbHjOtDW921n4
BdaNSlOSKfpa5ccwtIJObgwRquEUxwmwZ/dBynmTQdd/+52HBjACqLdkf/SuFBOk
rG9MiXfcBMxqUEde4/YM3TQtwevsLLVaZco1psFl4Sl+4R3SbiAZMaZQd3AB2d9q
qwGiKrCYhOi9b96VGXTE1BkqF3AlEUd/Dwy5Ahi7NqGLHhdRstA005lrMK0jp50d
lbf7q4Dyf27pGJ1ihAN7RFg4w+VhFi2rqTT8Yl6dpoiZMbpOIzWqRIbh+Y0gD5He
6X9DDI5dqtog7qR+bPXGacHgG4bStBMIxRnLWyADOEq1Zeg3AEql5s47wXZoU18t
d8o3GxbBqekSSXzVd2HQBjTQaKyRPS2yjlWQVD8Orf619PZzP97V4DdpRyAKWn1c
+K1QAFsAMhWqNLFI6xEbW8kHoQVqb0ccZ335BvgxIQG/h8orl3SsbjCPIuVPturG
l/E+2wf1sLrd2Lz2NzlCHKbkTf6J4VinlRoX6p7+dcbgmCNnMM4NHGz0ypFaRBqR
u11xXjZfqWrkCPrgZWwpuB2BQQdui6bhrckyqpC9yT514kEIMr3M00ILakvM4DxW
O02z0fH+v2VSPU79hw8zgSaLcXljfEEssHp/vy3BgWZg+3jdyjyj0ppmTA155Oi0
jIKJVqhr7x7x//rFH90ngg94rEwlz9ksIC6NHygjHewsVWVBwCt/yQzExW7xjQjj
fqNsg7SpleiIcSP/tIM2bVJRsHA9ZBi+FnoIjp15WSNKFHyCo4/F0dKZYJRac8mR
RjB//mH3ptM51KrzYT5ylg46q4Hy+jPIHnuFZCQJxTojB7ZBD5Hk+7ytsCgYj5Se
WKUFIo5ujTIWFj78FQ/r0KQRIzcZd/3va3ypcBiTBfJ5JGNfmel96tRA0YhfLw4B
8LRKp4uTzmCwLIFr5P0BoXzRmBqRZ7dTgMqU2KnvfViv+i1H3v6Puudqg9AIfmRC
ur1US6IgRdcGhO+jxBVhV50XcxckUrTd9R1eTx5uNy5VH5FGe5qRfDySrD74Qcqp
tWbIXRjCXnQOxOUdmH8Jfj6zQxyAat7Rj7oHBH+BqIMVIVlJQ7vSEmY10CgnOpjk
nIdg1JFh9q+uslzV8u0+xTzq6APwWaWDT4NSD6TGG3NeX4zrUB/odBy+XfvOuXCP
tGyQf9VOxNlbTSBlfuls9+qokU+oZ6r39QZ2PvUK/HaXT+r2/js1D8Bz1b7uYd/x
vFyd5LlwiDniOIC8CcrPTT5jUHDn5S+GzT0bZJC8tucECvtyOuTvyJ+iEIo9wu9H
jv6FWuKWQUNmJYHkv2bgvzJu4Y9DTBPYVA2T4Q1vb0wWoHn+bfjOPZ7dQJp6zQBJ
odWvjs2fESPQidbAuJXjgrJJTg4Ncv0PpThZw7d2+gFwgzHEY+s9BzIBRxxQOM5u
A3RKdUsbhUBo+U2N/sVjqofV8b+WB2nQN6GFH3+nOFYEeHLIpnr0xCmPh7wqSe/O
voDAAUAGSZwDByHh/3iQoV/X2PHNhzhMqz+bsZMI+8uL11wgApPpE2CKw5LDxokU
AIxybbCwwKsy7mXEGX9HXILXBGfXi/cLhCM37dY+WEULSVnr6c8p22oyAfnvVOjZ
ARWsK1FNXuaOuAtz++tWrpwk5i+zWXPm0gre6S+RtclkokTWlzlxW2LB8NSRDDAm
pvKza9sS3W6WDgNYtdE/4dc5aTxPr1vn6qbfGLihbeDdEbciJMdeWRQB/HTfbAwJ
BOYynJ4hh03UtJz0JkvTHsWM4OmENAoKdFLfIWMf4spP8GeZeNv74VVNr0qM+LI+
VFPT4NNn5yHwRtD5lo6q59VoBLVQIzQ1e5dwyRa0ExJ3YG1C1kREg54CGzrFxjgv
GGW0ul/qlb+1m/WO9RlYzXzI7lay9ST2eLBflMRQtbBpyFYHs3dyKc7KcFQAkmxl
jGXHecaeambLK/dgw5wA/sVBQekKXlpL/iiyEYCE/weY2nZKAFHewojRexdNhTCs
QeLOoXo0DuV3fBBUHeVE4/Nj6N9sWO7X6i4dWDPMiRPSd4rc/nNdI+vhFrjkCgw9
TkYJlYCPcB5wvFDXLHQKklT3k0pU88pXVUaqQVjkluLRL/cf8DKiTZCR6e+6YEKy
C8KhTupMUeNtDVgu/L8iE/6mKonvWzljUO3m5PR7vC91l++3n9G7AfWAnKvNLpV4
6kFI05R2ygqcmxMST1SgARfLkCV5lLGaBgKeNIIB01HhNczmN/qSPeVYV/I4zWhp
RGbIzGWjnabI1Bsafxj1xzmKPo0eVB6soASTRgq7LT3/e+pVZzdRaDe7lfOJeu9c
ZUfiufs8j1R/Nc9ECfH1H60qWkZ3J4IXFL7aH1ANjGnMShmwfDkUH46yNn89mYWv
bT3E6f4wIULTNi/nPwz6Z3f7qyOuk9QEfEmkiUo/yJRRrHPJ9dfFQx5mpqM2KUnO
jxrL6/dcRh04fHnJHggl2t2ILKLpvC1UdBEPTSLl8/siP8ibNto/BQAiCUO63d5J
Tc9Vnx3njlorprbHifr4KBODA5hcUK4wjYAsyZAm0GSupS769IxkPP+ogeJ6y1ao
CZj20EG5geTtVlKq841JY6aj8LxBqaZ3WH+U4qZf+YbD/1EuHj3OXvOkhDYVnAHx
Clty+unmwj5O1wroN2opfiWE7D1IYJhlhHNJqbeW0XQtBBN02/nyllQJsPmU/MQd
9RJdhQj9rGDhP7itFAseGP8MD5Pl6txhZ6hXaqhLmpY7H3TUqBbe+DqRFGoy+STL
aK4bbLM+u6W8yWUsENXzoIS2Gigkrsf2bIKv/9OBwzq7pb8O05nWv+EXoU4CLbCk
HZQJelhSQIxnWl2K8JAhmao2AHuDnvsdMrFumgaYzB7BhgKNmfdqVign8dzFYD5f
ZYZLFLOqfm0G61nOkhIIfkq4WR+jWW7igShkquNhv0QNDN6eg9uZt8qJvj2YMWDz
pnLUAmhH0HqiUxRYF+NkqJdCp4pRNL3/yAnctKstiiDQksV5YSu1luolaKtaU4vr
s02ifYyGoRZwbtO6odWHle24ewnHCi5TZAQRWLzJ4zE71XZYjoLJ1EKhcxQszzdW
fYaZvAj58argZjoxmQch7gg0DHlZG8NRtf6I/TXyQamg3LIbE9jSWwls4d36nJEd
aSefrtLqxcWbfir/5DSg14NqmYrGteN14B6IboTa0MLbGg9WaqVuqNiMY+aCCfUo
MGR2LUOwZTG/SgD9cjEHNSlurEW74CHDqs81XaO/YNKEti6gp7Bwarmyf8O5032T
ZY5f3ImicKLRYNTHNnVZY8y1vw4ceePM1MPuz1sTeC4B8vBH5eL8Mudv3mz21opn
Mu4nXAw/Ly1ka+V8LszE50xj/B8c1ojMqEeYk3Oza2ASz89gC0Br0zAsTWtq0f+S
um/3GhgLxIo+VGKdZi/Az3/T7XS3f4zVzFJM9qVXcR9osDHnccEA31+VPkq4BM/M
7ov0P6NOPc9gE43n7Twisx3UNXC49S5U4d9wb/Pvh6kD9y/TPKO+KmLzdZHJbabL
DQSmMTggtHofy2hXsAUiazSNy8Br258vIxE6Xur6T1KeBXz+tmEpvWB6kO3+1Z09
+4duH9KVd6ZEX64bAzC+JKxq1HPuYdtPAOV01YGk0YkUVSoHDh3JmUR62AR8eUEf
YI4TGlhM+c4/xYkd9urZC6b6ncBsIYh+Fly9FdcXQdFX3S+700X/QFgImPuXvou5
34XrZSbLJxyiMvVJY+yUnj7Bov7Ddx5sN+56Q/4H3jejc0qt5YzL/CsQ1WKU7glW
xnds6cPLSmZC/vB7QTa2/IIAqtFiEl3S6nqsvjEamdnoIojXTdjzyWg+25QmgXgV
i25kaz11emjXVXpFxS6RNdiiLZdJoZZ5736WbHaD43FGEe7kJQ7GPDTLXA7uW6DM
JOIw6phWyZ/DT1TEKmS4bvP+wGEpPOJ0M2KoxTc6Wdvx1pSe06jS4r2H1WKp8gls
8kEU5IAFpwqbNtY/gKR6RYUUvs9P848rR+Jgg6mXt0DtcO931qbojmQDYVzeNk+v
eO9J83TwVwBVbJekcx6Q3ws3DOIUDUw091i4+09HYIj/FpW6pEMZDEkbrnY8DR+t
QbfKFfFx+QjFmqr0j3vKa37DrplDDVVeBhWy+b6wfwfHkPbuL90SKw1csxelvj0E
3kDgai4mWhGCl4+2vBbuz6q6I15Bx0owryQvgN3QZCUTJNNz0fBP623XIPAct8xO
SpmwqgCkfQ2bPWffWdWMk0eUN33l1GZzhczyhGygaiOv7WUh2iwlnmFu6XSc/vIe
zMbYmf8M+Z1zLpun1EwPKg==
`pragma protect end_protected
