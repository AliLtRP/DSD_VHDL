// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DSUq8iU7heiAb0c3Xxo9P73Muhkvfo1JOQum2Nch4nQ1pDXk6Bmoh7cdYt76HMjD
pJ3l0b7IwoIdQ52RUUb45J/U3Sh6xzUoKP4VN6tz7Ki4lqIa4433nyi6P5PcQp3o
uKjmkExsdXIRU+l57NVGc2f/PcDAiHrbMPjLc6WkGIw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19184)
p1gbzIS6DwEJpq/SfYML1YpXyQrK+pkk8GegSuqcbz+snaCl/dUUPMJhtbBZXjEt
nzlO/I/SKti0OGZiIN8H6E9W4B8i6RW/0yrG9h3I/nm0ZT3c9r9k/2S3J7E35mrn
iOxtaeaqD1Otx2IUmnsKEZvyMHRd4BBqiLnwqF9OQ9oMN4+JcUpb89mVzYDqgwko
am0Uw1xZz23Jpdvb74TOW3KC3LYeH7GbGwcf4/LjwOs3L8gcMBQrsIS6zHvonYJx
eimFM5PGqL1EzvHasmdiIbysGIOVhcUuJQnRucmJ7hKnkgpR33TVPXT4ueD4ZYgG
dd2CzrG67e7mxrgnL0NrKV4bq/eWH1DDAchELycH95cub0yaPaMkh9qhCFExmsOf
67scoLFD7fP+22Cb2VaNTgqcel8BgIKZeJP3gBAoDXkbiIdBk2SMlbObaakoYunu
cEpVBY7q6Oki0q0f+XiK792kv9/6C9ZCMUyMZZleTu893wCVbrT6Tjl3wbjuUubd
ZyuvkglfJwkTJnk7mWXl5e0R+EmIQOoxoXilvtdQ0BPjLKsgczCnrbKdGyadDXAw
MACdEP/4GszlSlx9HukzDUKqnen/FU2Qj7VFaOJa2leo1y5MFQGOgdv8OxIBzeiv
d5dTxNJwXWUInXgNJE5Hgvy2M2g4Oadpq6uqCdZHJ4+C9zHvdkDuj7TF1aMmfqRa
dzZGUaMjdtgoLy8Kr9AzLUXNcjZ9BgEe+EsqW8TVoE3nl0PnA9f2rTfeQ2xNSWQz
WCWNwOBpEV1s+2naQEKw9IRkV4A2EV6NcbURjHKaePCyiCfuGv273Hlk1tFSmYdp
JEu2R3EX0LMEqBnlr8bASt8MIjmM6vOAhLqAdDHW5R6VIIZTuqimwMbA1/pwBamk
MKGkOORIiTHEaXd2SSHitZ8xnVlrBTh1U2PaeRzG3DI4TipBqMl/ohG0lRcZ99dO
/Wo0ybz36ZvE0jC9sr5VLMo7nemxniIt9e4A9cVUUl4N+kIaihXKZwZUVoU3uVq9
oOYt63e+yBSLCDO6EJiC0OI8k6dT/+0bHlHwWo/7RkLs9ZQg4J1glGyb3div68IH
q9H2cG9L3NsGWkvw8NR29Fo6kLPvEAZTluT3S6gc5XXe6hyRIuuesNCX2EMUXdsO
FqSl7VlGIekJIb35ArMYNLh7Xcw2+GNI6xYGpmy64M72Q7G2axkPTjCJDSxFAfRN
hKi6OafZMeCbJ1ufNBQ3kkrz1UJP5IrRGeco5gaEHE2cSarAbt/xY4ObmqoOXGrk
n8LQYVCkQdY3bc/Eu1C9j/vfw8UdfccrTg4UuphrI9IIZhbGqeh0uZyy1IMFwjML
P2+7XF8mAxIvUnlZrQXPDqa2pEaXiiwloZCJRGY0GaLJM85sP7yL19fYnK06/doK
NrivLhb956pI1Mx0yCxKZ4tU/ypQaNp26ru8JaC9YmQNXdk6ZSEWkyRd4wSpGdGL
BnQbnK8Ko2/VrSU3KmeSibFJg525y8wNLTe/ZrrWfv2+FSH+meRGB221ImIi0jwp
50PHtk7QPFqhq3IeIj9qnPEZoSm9jUSYkyQcSYO2dpcEGukQyeWsUPKHAoh2F+ye
nBTLlcQZ4C4zK2sXS8vI+iE8QD7WME5+hFPLFPrWFZuNgeHY94AD/IFRCMK6tLrM
B4X5ooj43hcU+hb8u1Y+GBJgI0KTJny/GsTGRNUhBpxa9ipN2+9SzxpLy6Rm9Sku
T8ATkUx2yLUENYlv3cIj6oN2V6z/I1Fy9db9jm3lLXGcuzxq76T4ClltI17HeLvA
iEHJrSh3dlzoRxout5iUPK37SXy6EN3SvcwPrmI7OpGZ5e/MzUifFF6oGDjyseIB
lPFLs2hStCqN4iTFI4T7r2JkTHYm1+CAtwGuifhiX0ur2FPi4CmSH6bQ+0WRJjGf
G5QHX8KeuwgKl4qaxJaH8Wmy6PoZg6g3/zLv8N5HboZVTqCysbS7ufPd0zsyn2la
6ZPGms7hnGnlCLhtQCTZBr+fIW2nXQuNelVKq4YSLa6PFDJaxcrMmtwHaYzEYCeE
+jvVVQeIuxC2w94KUOW9SQIyWslO6B+I99h5gXkYFoNFpDc2qiPI60oSPwJwuC2Q
XeX6JaD2+Ou5QYARTw49DLF1H7v2RDqrGvE1RjfG8RxZ/4j70XWPfV4+5iX+b+gJ
U/iuDMeKAAmLo9k713Z0wMkzV97cgcIsTMx7O5cfqOgamI0xTB9UubYk1qAArbFi
onY9hDRmSPUDf+GyR0vBKfa2o8YacEfYKQmZ0VloZlcSGTJdBVScyklvJJadFp9/
klPLMyVgh+Jq+vKNRIDwNKeNBnHb1l1yozPGPA/cMr2hhenFJWYw8tzyuJl1OMUZ
vaMfLEh0vLoHUHSoF4sCYmqs3u0/a4qTVWgnCecX25xX+6pkmtPUYO2FVF6cVSsr
qslOYagUPlTXJpSvZU6bxBNH+nq8I8vxCZrmBe898kwrAVDPoiXTgw9bk834cLhV
uqTlYlvITAbo3IjW6YCdgyomHCcKMH2LBG/VbyefIcaBRqXh146vWLZa7ChkfMfR
NET4tZJDUqDDhjafoIJjNIGXodAQtHMeAExI2M1b0MjgVnoApE1sRuIk9HvVfSR0
d3ZxpstkjPnVut4tij1ryZuSOX8+8+4wjAR8VqpuJjKr6rvDP13sUeaLc0wOVobv
Zim9gND7Go7dM8L7iJmSOqrDLB0M3MgLt1jst64A3o0VeOEzP0Q3zh+v0x3xSKgK
L0ahQ76Lj66ic80Gr3ZxurbEJcyu8mPQbgBKp1F3be3/tHPWSZx08argb1/59hWX
2y7DbJWo6ujZDuwApBwNAAIh7xtnWkkYHz8yNA4o5nZ3lp7WTKq1jeih0S31BRle
viAXzcOlC7nkkw/Vbm3Ml69fx0Xbf3P3btgWuWn9y/qhQk8Reqr1d3cdHbD3SFnE
P4AB8Hmkw4cgSAyxDFrzbtbI7FwJWi+cXPF397B9cg802qYiElA5qMTaFaqbMdQs
VAhTo53CflJNrm177byaTTxy3LZ/MDT8SuG7+nrg3AiH5JOfBIRj00AbA5YH5ClW
oGWnWJKQMbXi8DHKeL8PuHrl3U+fXe9lZgssPaDD8SnNIeN4wMDQNuHsdURSbAAE
vdf6WsB/q06GMy2JEpLrA/26DSPLzpym4ljGVArLg99IJCKOdwN9ROLxstuzGRLX
ZTdGuzPoDLuZGzwVwVzJesK6QLgH1o5Mz3gBDH0L2foNuk2QCp0gLXgrvnesjCZn
TbWGfdBTStNnyr4NOyix3MEUwfzumkvd+5NvSqIGkhlKX4+LKS+AmlDp3xtwxlAM
NJ69gtY98gQ7v7N3gofEMW1kx+/kbdzLDIbmSQoJq9E7dgEeU5FEdXR2lZRS4Q7M
k6UaxwlfG3XCryb6T8CCT9VNOBWHeP5NfW2FbWcgSmDV4yX9VqpZL4UNIXsUBUbY
2kPEJoO7hi0ux39eMukD/mKnrOrV9IB+N1rJvRIOmlt1kwH0Igdi3rmhjfIm33Wo
B5eZy1rtEM0awlV9XVcu71n+4H2SynEew0Xb94dMHGKoxVptgMEgQ6PVhWcRNEVb
08VW1Z5gCzkw5yh9UJP4IbqFE7Peug/doU1aShEySck9ky661MZJ1yHNMnzMNL33
OaYxrUUJaP/FSXAbBu7dZgp7KM40k6mAONJwy4ckLu/nO7x6blpRpddsZVu90o4D
gCqlCcxc4Wis2YyN5jtCG2eAGseg/hXk6hmYow2xcCUTGrnPzCcwwzi3klYeYlfl
+H1E/N4TiUJhTd5o5+2qelP1vh3eweV9uYAtkUwgambfD5XEY37yBR4V8sM24ENf
D1l17tnWkmHLFdX3TCY/ejxip/t7E/4ZZkZopFg/RoDGyaglOxFnOflIT10Krpf2
7e57a8+XSwUSy0nFZf6nJfubzCRASLSk3iTk7C0pQUlBwE65JR+11MRkbpb5fZoj
TjUbC6hWmpmApQmnOKvoP32gLKxRgn95emHKDAdY+8435YQIfzvUZpMM+cJLnNGH
OHjk81s3haQLwWKihIFBrMy8G0tBzNT//yBUsguS7UEJ5HRw9NNYCs6cwDCaLIoL
fqukec9b0WTKQhaVcudwDII1nVf2rGwpX/mFkABcq0W4DhNTUX6oL/5zaj337ffL
2c3WTvtCtZW26kEAGq8BLThUBmqEmMo/YFppa7UD7Nuic0x5Lg5jYvjiw9CSnP2c
ifAfFd7Iui1nbpUKKGds4WoqplEHQDicR1uKjAGzTnZuzyU8pP2h+kHtXRYEY3iB
7zGyURSbKE5y/1zAYl15kSUT2U+htodgqGeFYRAqZAuwyLFFLFzP63PgJGo3c4O1
eq+2WG/mz/Vcp55KNspMOV6Nq0y1BTKn+iuxsAlf4vyGIeyjE7Q8HZ9uKbQ9VfET
gpAyztbGqn6zf0EP6ImXvj8vcKru8SmwjMalAo/6h5lX/ZAtYLlMRw7dbpDVim9i
cQrBXCRVSqF89N0uwq7Q9tl15bFXarm489m3KIrdFt+QTV1YmMKoFkz2nIOrmbO5
4qMY95B0PkNh5AlOWWtnIWl/YfYY4t7YsHECaJFAL6hXHa1H+0LRDZBQpjvL0maK
Dd6sqDR+7hDwuVy2K6eVcLH9M0souUt+AB6kbYGPwSiY2Y+ocWHpjKoNbXhmy4eB
W0x7/DtuAhVBKa7KUpO0X/SbDh9/FQgF4mlmR33obk2cQSj2yvsnA+3SmKmwr60C
vr872n+jjYXZGzHE4JJKlnDU7JAVs03wyWsot3Y/7uHyboJ33rX/sRNPjR8DGGwJ
LGgL3RBRoArwcyvZ1f67+nCDFXWSwso3jwSJ5fSjgv3Ig/uCmeLwp37BAtU05nSN
5mPOppDPvohnVua04+Wuc53hCysByxWVKWyiWpDyNOMrAGS55XgcwePAMAmhqv/C
sLjKANmSeD/uUtFiFesA4779MZQ39k3GK0CKufyOgsaUHVS1SQIZgPxYj+FA+xoM
OvpugqPcxekCjlJl3Q+88E8DPZGrld1flWO5y3cNo1w+h75/gWl/VQ/B3G8LZtQN
/+bk8jLWLuiRvVaCkj6ihniuRNHgMbbhfzXtBNDOOA4vBAeLxzMBTVdaNG+IEACx
0FI289u4cTKiJbOtbJiIoT4606EXZkG/807DxvxpTJObkNyubIa3OHRN6MtM/d9x
VAzIgGGkIWcgu6V4CiWUqjfUENrmgRYYV4+BTKZZlRu5VTJSOLa16IA+SE6G/tJe
+7f9D7KND0HevergwXUlsOj97IAKvN9ou5i5pVEtszbf1F2eyeRCWt/0jxKy3tZl
fMPWaqmvulOz8nQs/nFPNsWEG3Q7An44eO/aoOqEDa79bQvorFXtlOL3nHPh5JXR
ZkYdVNFJkW/nPt7yv1cBW5+7dpqkSROGO5pP+G5tE0c1Ovn680tMvH9xwm/myLet
eYKb7ZPGXPOdaOL7zQKWggvXpYHkJ5wJHTQJqTrZBHW1xyrhfD3LfRLWC87n5BUm
5PebNQVBUxnMqvLHcjSKxrDuLinjbsGvWoL5PHKeoHTLLKlJfu16B+lOTts6ex49
5JCCM/EnDOswtchTI5nKq6zkse5W9g3k4ivG4f7lZesWjHTcs+dGn5fIB8uJuZNZ
udF0SBnQPrwtgZYZsEFdRwp1dI1KSop0yPA4iwFjVcNXjldw8JFq1iH2b5E4C+Pa
hrhU7r64QkzaDpFYCO5sQ6kFqYNcVjAhn6Ble9z6FwQoQ4J4wyQV9Wg7YQoEEGWl
ryVvzQHZc/QGQx5A+1O/8nclpYKDOz2oWWSCdCzvp1mycMusKsIkUqkfCz4TKb8x
vEzksSLWz1hWqFcLuww4HjQ/6bHuWN6O4nMaWk4W/HLuFxh7nZ39iJupIFVQqfZf
UCG2ABNb7bPUCM79JflpwFF4tYJupuiJ/ilUXuoDxo8WxPXNRxSF3WB9wG3QBbM0
9Pwe/ngELCcaEL4iApZsqRs0Tzpnj+t+aQoT+3mwJx/7ewRyEQ0/8TQ+/RK7pSV+
/NtXG2PzlzfEX94iEuj9n2+L95p9zgjSFuGyoc2gvHA7WwrUAkXYBIbNgUpUkG29
rrik2OlqZxSGFQ4l9aIVu1rpYLi9XbgnJLb9rmXdbsbFS10vEURgP6EkEB3e9Mvm
4MsHxtTPRkEC8Le8OhMAs86bXKHYudvoaa7gP+V9ClDigSy0sn8prV5cajDmouSX
ePOZnQkJjiUsuF5qV+ptZSe9HTizuDImH+rWK96Fa7Rnd+2Sbfs20bmjXGAcLxTi
bfAn9q1NeaSjJ5oefWJ7kySGVb8toVAUsF0eW4/p4shyJ2+hf4YbUW6U1qrk1Klj
DrQuKBRE1XV8JbD19MfTbA3MNl1DvBZJmzBl9ZhYcY21ZCIAalhsrn2OFC4jSwxG
VjyO8OclegLGyyOo62Ss+lZFUcwQougzSPR7QzbbBizJpBKfvT6DsB9Ip8ddCLo5
kzxh/asdXO/pBRzP42pWqyWy1qU1EnUV6fmiRJGL99M8g9lXivEfCIozsomxzfhV
2GlGotxR4fkyY/sMWz+/WOC6XUSyBU2VRUHDhOHWhbUxuQ3wc9aG+PhMgPotIsxP
5V6BFmrSFz3hAVJI4G7ag6X6NBabJvlo7JWDgV6qFImL1/UFyL7SnYwb/+zBKidd
P7tiYz8gm6G+oSerORwvPMr34xnM3PJ0Cgp8BrGA3GxV+6fp6y0sSzGLFoN7eI1K
Gz9T2Tocht2vj03qXPfWqDaby5kjQjhiN2KOqzYNzpp1wkCyllc/yMfIPe7ftom9
W1fVjB7ZCdCfVv4u2XVLSi2S7Gzs4GM7VOo+gyadiuioTdKsHi3gjXl37UmVlfVg
ex+JTtt3SFxrLujO9f/cNnpOzszinSKII2ohEwxCwNTaxdnH6/+DM8ags1GqZrM8
PtCPRpNymKHOYRZUs6QZakqU0GFUzTElDcidOgLx3rAYz+m063Dp471Px2clKfeG
FicICGvJJ9PhXzdPI5BwFgKtZNfZx3PD8GoRnd6CJlCE8G3eVrJPFzbn6Z8rMWPB
OWrjFti8jDL0Vck0IySCixNOOymRIB4zwIap6SDAMrzlhykWaEQ2Fw8yBGnzNipk
h6zXQRkisqTKWFqKWZ/MtEjUNdllpb1rPQvCYAjE7wZVbpObl5Epvcrjrqj21iZF
Jqkxn/Hl49qmhje19bk4PT3xCoilIyln2yvErNhE7rZ9SBN+bn4TyxqUrlbJLqiJ
VntoK2ppyINgFiFQC2BI2vqhsDyFlD5ISxRl2183l5YwHFlCvvB/phO163InmgyQ
QJT/im1XzGckF1o8HDrI+qisq8k8KeON8ad7uTT/e8mE7TMOT39NY4vITyglPKor
qtZCHH77lJAC34V0Q/xG4noVkAzxmRu35jGpBK1WhIloNkcGczOV70f+maC7N+j7
V9mUimF+o/V7RKxAVBY3SdY3kFTLyu9djKQ82IWoqpuTcork/4mBZaEOxhYmhd8p
neBr6okgetd/iEg/R5kK97gqL6Lh9vPvvnPJv0h60qDEyeY/De0nbNS8R40ukY0F
hGkznHUTJthMY9huyzdzqugAuiSMVc/bvo3by8Umfi6kdt8lPAdsVPvo4F30AdrQ
BZ3+H1Bc+1R2DQAJILtBxXmkmVUWK7IYIKbPDpyL7PsH1O7WwRoSSH5pIDXcVTqN
PUcDVEgApMdO+spE1xaSaEdkt8FNgFsB9uU7T23Nn0zptQ+prLbhHx52cZEpXW/5
1nVHpAbVFJDmEjMhp6n47YPTOHCHlF3Gmm7CEM9B5IXwrhvRHCMfK28zO1egtc2o
C1Y+ntpF/XcM0BScPEZMWFu3G2WuCyUhF4WuIJZueoJP42JOCm+BRUMDOz2Gfunl
eNE1hw3k5cj8mjIssSxp+BuBW26yDXzoWhgmmoIwoEEPUAHfZtE4KGA7rGpEo2Ny
uIK/fAiTCqApHLdrOydVyKncKItvxoMxVzEOxpsZvnU4IPsiax98YxOsMdjPaYk1
KZUODAelnK4sBcObXL7Z9cniGRyS1iMmkisrC3NLifouAQCH4I3j5XE0/goAsOjf
fR9fOEIwEWraZXXQEsqSKu5gisXG511ku5uO6tS0v84RZYw/Ri6rLPfFfZKIoTHy
ZEWavNGArg539kO/ufgqdvo+22ZjcB/mKjcP5txeGT/8w8lyw7yT+UvkSsY/PDRJ
15LGi5pG+JW8eY+vYZNdzjusklO8M08QRcaJuGoK+JMI2GvS6zLpfaLtoEjyNIH7
OJT7Lk7LaODV94OYYeoKff+ieAIp9YzoYUqxenbiNLHotz9phZLiu5EttmCM6k8x
vf0Sb9JKI+s+hCygrRYfldPfRNsOUqF68Syh1Lp7jj2PbLJDJZcoGu3sib97i7ic
iTcyrT92Ja0uT7FqbLR1ahk+Wwv/9jCVwuougCW+gz4xWfq4uBNrC9Kk83Vdy9xM
1vfIt1RKvPsI5GPsOg36IumJ+F7HT3MLk0RabAo7Rc7lkVHaxwRubzWoEe5hhf8U
o0MqC/jkgYhwE0jBCm26HCl7aiVp4yYPfEbTj7dCWjnDmt6HF9G+uCiKdoXWADoh
I4FjurbHSYVAWdNwzyLTxQ1VdRBusUB9Slxp4xwwWqG6T7mNQ9YEQnOmYMfmzaVz
AYw0Kg46D9t7mH0iIT9U3Fxej4zQzkO28Eyy72tSg+n+dEuHufsDyo37mce0ttI6
D3oNdFNrHr/set6EjUUtpeZeIXoK6YJCoMfCdHtKBvKtVC6sdmeV/h5fOB5Mp5hd
e56SPOfLvbtnPqtOBe7oloHpGJfqsROdN4ityxTDoFHK1+KL/diYxdG1MhRkPh2Y
lK3FSe9kAHS7lB08NV2x6OSHxZNCf7J7IVFgH4rMvQ4Z7glzGD51KEi0GaE6Bpvx
RgFqsl+RvIfdtAB6GKL9RvarJADnVNlU+glYw8MyxG8Ua1zvUWv7iaFtM7u9/OG1
DugmEyS7/OTAu7DmGiQJcAmzY91V19vqRaQOsy0rahkrV1dYgvHCNhyERfVY9gVp
kLBQRsoPHBR8kkS4+ghUJCnOZ5QNf1HcsEkhmN8mbWGRlHOWxMy4mY1vrXFXUq1o
kjwpkPIu52Jov0VfVdvROCXCuemA4qPOfm0xCrnmDjUE6RbSmY/gv0Vojfvfdl8Z
G+6n6k2PpImr0f4XfNA+A5h7f0Ytg9f8D691xiWvsZB6x5ZNJbcjOGOtPq7ZcJsp
iwAHazlq8gCDp5P01scjSDgVz9CCtvJ3v0DivP5dWgi86OSOgbI7APPyhbor/Dv4
hRe9ZRoUBOECx68bKXAOo5GtQZTqZKQ0AePsSES9xBbm8+V1l/gRcfuOyeCXBnMj
3GxPNbztRZlAMbZYdOp2MX3KGWk7TMlWfF/QhU67DgLw0wI2fxtPRSoD8dTzkTWv
VMjnoPB+6vpn3lutG7iaJ5FcqG40fX1zS6gdZwyTEHys/GoxBOrARhPohUdzT1Kx
uEKM5Bxixu8un8W6UF3/YeiVMwMdWt08a3ZUvUCbhhU4Wd2jUneRhsPIOJwwLtjR
wfWs67fS0JXIi6DGTJbgfjDArexKDUfGInUi1S1JRdHYhEwYV24frhJHMGfegwx1
k61Mudq8u1CDdNE377HbE2OJEvLsT5QUmmVtFVZYsNj0AqV6/W1hS2kj7GAiSmAm
sQQ8ngihpA1u6IqiS64Gp+uEuPBqbbaryihURHXVSV2ewij/jK10BejKyWYYJAIw
mVzURRvltS6MyNgyzCmdHONCI49IZnAu7wKzDUHk6R9MiSpPkyqmvCx/bFEn8V6Y
qW3JT/Zpt0RFGStsd98rc6ziY5tTBEJ/j+yjeG9rLi980uvB6yptQ9KU3RptkcP9
3G+jpm5+8M6Us7X305cRUuqdDElJD400lcXB8mJAsXaFCn2RTauJBGYYwQEqW77c
siGcle034DhRvE9w8DEAJc7xQL9ekwwPN5PA/hTbhs3Fv0qiz/HdV+XKY60h54at
shCyGyyjskLCSbRx+ju3TA+M7L+x54DAXxM0V26c1K6jL1vfSJclPL8NdEVxEJqZ
UJ9g2X6eZn+K/fmMHaxHoxzjVXWYHw9b9BIxQv3KhzhkNkheaF6ceeXbDzK6ig0z
nfVcsjI2cgzWT5gak75jUSJB+Qvqeo06Jc7DONwDVc8KrmiM34ew/RjMXIF+uZHq
U6RLDBEkmOS1WIl0vyKfxNLdURguQwYQI3E4TXgVpQtVrKd1Qvn+mfa5jbvSHM6J
c0V4iAEdNur+Aw1gNE3Ug6D2bTEkJjEQvO4kfJ8gLgAj8zKXvsI2OOo489b7KVR0
g2OlLyDmAb6VmgRqwv2RXJigaYfRSFMaC79w9Hvh5wcrSMeC8H+fYG8Lqn/NtNbH
t+yK2+BEJkdFB0FzCmchUvRrrJOREkxozxM+1YAMEs6XwEKTD5vNexg//xED4Bu7
+fqgFBWbn6vFY3jHO2B235hyjk6ZLjjwDNwKj2ipUuk2wr2ISZGmfwsQpsXezEdg
Zfntk64/iTb1PFaBchapgBVBA6DeoX6i86h8KOR7VX9oBollPWmtGsBn8DTQyAf9
k28mlrdaOYFwk/ulZBD7f0HkwGEzc89DQm6aPgP+pC6Ye3BspUXYqQSzGufALMPH
/KDxx/vTemB4Fe2EHnPARsdRFX0CJE76WsusR9Cx3sJEf1IPoOpPygwvYM7Fz33V
4ftZTzbqV5Rb7lCstoo+AAJK/v6tH3bapokou/Zl0hlWUrtXPDYsdcZdKp0QOtUw
c6Z7YSDOCAPgoWgQLtC14EE/+G1rgfhnKROO5Z5wJb3OX+cm/Qn5v7YiyQU7OSVu
l7t64FEidQ93dwKVk97tADg/FG1h97yRr8sE0ZSKZ6u1RZ1kC3bYVkmbmlI3D9Eu
bOuoNgPYUL9rAjk7yuHfGkJMzY5D5KogQOcf2IQknUcwK/vWHxSm7izCQsPYIBqL
F8pDc/ERevP2XQzi+tqdddoUhCrVtYClFAb0yULNyhr0q+7v0h274BS85K2kxRhm
AfM4o2kQfzDWB/XxeNoCvbtkN9N2WhaWXSPTLK0FuDFt2HOjjobIhYr2OlHC9vFm
f3F55ErW9nCNO29yG5xZKB2Oxt4D2VQ9r7aLKZ6zGnZNAYDsY3OslbQYd+5LP8ND
PB9KpjH6JbEwIbdnmA4foo7T3UFKOnR45b5ThRXY38SBRGrK+lW2/t9OF/0h/LJS
aHPALrzd9IaKpy0EGBh3lcHQol7GwTbJEpJJ7g4dBIeOSmnOTbnXTE2AudHpb89V
oY8Ku2dIQ0ahiftMgneyiKGiB3Bk0lZ79jT7OWYkIOcJCPWMVfH3f/NFefD2J+vZ
lgAgO+LWRgNzRzBZu7Ad6cKel3qSZSkmDbc8ohUDfpJriHxF2Dv4bJJquGz6IwXJ
hNBLiJ7Hy6bXN6hwY9FN0iWl0CbM89gLESLIPoixxhw2tcXyTxNyzzY7NIE1RImB
g9RjDkiXcNzFaYKvVgUzzoCVQPyOE7l2Nqb/eYbSaGJDOijK2/UxetIN1hFZSvYZ
pA1P9mTR9mViCkE8HD69bpgUyFe+GnJHFti7FNPOts0GrYQiKa/cg7Wc+/OnTARJ
tnwKd1GyjvL1+R6iy37CMkckwbmSXuYeWzvSd1nNiUruSWjkk6IuqhpDNKi13hrR
l3bm2ysKtsqGVVuk4Foz9Q4xkic7bwBAVweJZc0Bq4cr+wiyTfS63xpk8i9/mVSx
xDye/b2VzF5Y7zYaEnd9N5znOtQ2tYZqIkn8vzTaOxQcAfBj+AkgRcCGWx0Q4k6N
Pa8WOkLomqIxJcQNtBDsxioJcW/bSKTUDAY/ld+s0Nf7ax0u0eIP1bKTjHhTA6B5
vFv5u02iaLIeRHaqXHT7CQ5P3algQrR0blqrZu43mDVtyqScv0OarMeikXn/4iD5
9zTeWDmQop6olwU4gZ9cU/M/NlDxkRU/v7riBf/Y6C/itmrSMd28z4arenIp+56Z
TerS6gI992T8kCev2PMCSScLFuZjgwo1blCNyERFjbsGETWlpTole0zVzquTbBGm
99WYd9Ur+I8L6cSjbrlrSsbDwFdZgfT72W5m4qge8yfC/GS4lQgaC72LrUdN2kUG
1o2K1tQDNvpLXhEmAe4ODU8etMHecy+X7eIdgvSIMk1AiiKPjnw71HYEIxM9WbLY
sZsJqxJcQ3EAyScjPZwCa5bIxHK8bnj0unYz0JczZWnwW9//kUxt6FyVCWq4dqUN
0FGWqlLV2ABK36fO4JmMd3/Qe0/uHSqT+OQHYgVXuazBnZZFC37942IORF3fuiLh
vPCB8AIe4GXmgn4F7qnOsJ70/kKfjPde4iyiLrvmefC5bB5xZvU1qynbUAz+cxZv
+Ec1JLTKVIf1E1VhesEzKIMfPYML/J/WL08ojGQQ5EMmGte6BF+CuEXjLL/3526J
EWt9eAu17vtUCBx+myBx0KPyWe9h+SwARTuaqc9gCJvUEdTltEddLajNivPTKhsE
M0lrnhfewb63/LyCRACPUT5FkYsB+FiuqYz1MftNPl354D4flzkbizFzlUJjksTX
RcJOyTXU+UkMYClEOjwliM7iJnEAltoYpYEouBTSh7QEHa/Z/XpY8hbFI3KDL1GV
d3G1Lu0QGHN3bHMZU29eQqhtx16ekevvZVKXC4f8opHXAPRhi9chnu9dt7jKD2dM
E6azspEJXFHKq5sWjixtcfLZUCRxW76NypCNmF/7HHfwhOvA7plakU5yzdJyaWkQ
IO5EN3xaFhamd9al9juOCG0wrpiGjYzx+GqVQw5yYNQ7sFOafn1QwyniJGt+/zts
xmRguv8YgfcZgi952OdsP0+a8oQ28KI5oVU11VrLmZW7ayRvK8QBKv7Lumy+g4uO
efvt9Yj3eLw/Njq1bwWMbcGI5i2eg9xMwnuPXnu4LybMU+nPcX0xBF6lUw5hUDfv
fThzGjRj1bqx7+4+tNgK9b88SeNm/kDUYr8vShWA/kyWIax9A5IOwXhTwFeeWnx0
UMeimr35N0mBe0ArMbUkSZzIYst4PpjjZJKcj/GVsnenaavGnQITKdKIuHZGU+5B
FqbEUotB9JuEUx6SxKgWzF5FWFuBn7wnQq7Cet6xsJtyNiJpdHC0vaV/iL6V9gRZ
ARx+6mLtrg+1yVuO4flTZzEFzhDjAIUTBdJyqtY5OsOPfoaAP8u0hmhzJlkSsdBP
5DycWH8ckEoDignTY9OfhRxcLUL7X7zc46Db55Ie7kxdioajjp8dEvwJtHKGhs7H
WdC+DpcR8Vh3Lr4uflpnAiXKVBJbLUqickaa83LxKYHAPQOWAN5mIBcPJtL0JFpv
M3to8MejNzGUSS44oRE7i0fvlvw1NYd1ndJO/M1LBiP6HNz58R+SNTQtoDG+Z0J2
C3aKTrkuUZEE4UECvqOsKY8zr1f+GUTsgwozy9+Wr4JrRTz7g2AFdv25Y6rwdFTk
doAFc0PI3GS8HlHsVPxmFPWYJNtMLTiRkwJKZ3yh6kOl8XazguogSjUt7VSZk8cK
9DYvMqYNOshpp6wDSQZrS/Q+iCyc4eX0Vy9pO+bnlmqx4gnTbg9d2M5MndeAmoRc
drkdxjJWhCP+EZ5tx0D8aKzyWWI84BSU969R5zBCclb4JA8+t47l5tL5bdry4KFn
wDqVHCN+A1/B/0hB5CofnFvUDrmF/9fGb7jrPsz+qUZVh2SXV9yrwYOTIRPmWUjC
WJG8QHA9/aTyr7lkAfNph02XVNdsXpVjMg2RPztLR0D+B9neTQng4apG6Z3Rxjhl
4bs539SaChMiyeBk5hC2MFPJ5Z3/QLBGD/kzOwiJoZ1dAVgPkY8P6C7PLfqPChoj
5YIZRa7wdRF538xM9NKvSQ6czC8dkX2w5L7DSXKwT6lg58vgOyFkN0CmM0afKL9o
4MH7a65XgLR+jsWceqRBbFAdwn1oFXeTMnfrg2Wf3RHPE5qkPNEx59DaASCQddXF
Jf0AuysGOCtTxAD5O7V5OKwDiLFU1JHFM/+aXEDzWqJvWnncjj7Veih+lGKiz3xN
0j3tuqvvUwfRvb1CFsblOtKf6NRjD0+DEryTWjKkfzl25EglFCLDLSebbqXk4OMN
N5fnPWY55R9aOjIcoYYKPWryI+0vlEzvWBIDeHe4AX0Et4wIvMpOrEg70uVJErZ8
42t3oshcGKqQXdfP/5TZCDFI4gzdXzDnjbr4xwxg3oSK0y70ym+e0flFhz0dShjF
klQF3g6ZeIC5pvfj3y3pgRV1tgVJf7v1kT75MsrXQnqEW0ya8A4g9ORmxQvGTPHV
+FaP4TUFV5xZK50Infyx2EMvS5PHbJTVuvVPgCtpXk7ue12lk4Oej4c/UyIuAcfY
LCNK1Rz7AGxg6CBfPAbK04NjVlK2N2kFfwk5Q6mUKVfZlU9ZwcWKXs7DVrN7Ct3r
rGS43B8X0VITMnMmPB39/sJcWfLISgETkYx1+01eJSnxsirMZOWJk2Pn8QEwliiT
cnqjI4HF7fSu9oMt+8sUjTHOH6SF3t+OicOgK5z6f3nhQDWA0RXPRSUd4iQN5JUI
2bh1RYWXYtBNjs1ZcRGTxZ+t7WY1ChtcPHwjkPNbrB3krGQZsweAczCCbJyu8+XZ
cYFc3MMnnaOI3oLpjNEQkLvSUVm0JFPJfjYaD82gPfpa7tN05/OEdMMe6qvON9G6
HT8XE7bVzzQVsTcL0mniCsG1Zl4h2Zc/BD+nnaBqSXClbtuwtAs3RD5VS8rrzC9g
ZAwL5x1fm8OMfmu/vp2iGZSyuBvsiPv2mK30RrfV8g25CXGrPOC+na5KuP6dEWP7
u7a+s3hIzw9Qk8JRIxWwJfyBlpMAamXhqMqjVxYIyRzNHE0xjy+HBWE/QIZ8Qo0c
ej0PiDcQNXWCyD9LO2SOBSwDGj3fzcFOSLsc9h8wuyeAi5cS4iWsX07YyGzbNsuM
G6sOhXlo0Dt6UZPgGl/oi8h0fcD70/Craia09hXT0LWEThLUE74KWqhp30yus4Ac
Bf//gOW/bBJ0zbG2l6i5iDmZgZsu9pxZBIM2OX0QvxBrfFQ2aa4cl0rULTXDA7XL
0mtsZ61/w29cvdBDKeH0uys9Y0EgJJBHT41qZx5FOnrfjrujIM/k3yYuw/N71+rA
tKjtx6+Eyt5IBElM60bf4cuYY5hPpJEei8882wzkvUm2ZXR3pqhN8g9rXdUnpBrz
7PZCOiNErx0jEx58etvwSmd2m8l/9xIFSn/Rh23g8w4RNED79dSHVJszDtYgkMDe
f5Baqstx4OUE5fYRWnXr2I7fbL+xRbUBjPUny9d0ExDOtrI5KK0v4xdTp9l9r2Hk
kpODJIpDMt/GplRfcdps/cvZjHFq9jermWlxdn4OROHg2i3881tWvDvMdqD+gwA6
i/MFJy38jZlF2z7Gbft9LRzi/FawerjC77tT3AwU0ItGjrMVWK8fOrB3EMiYoN8J
pkOvlXtmyVhB5ld3XPXXyd8AEpMlhMA6Hs2SZZ+0hvW6tH0z1Yqi8NGhUn/y6FFT
ZZw64xDgc1ZXTkHsflqqucWfvsBcsNiPTjKQR4AgUet99GH7bNS8mG+Oq4FR9m/Q
vgmFcUyP6jEtcoI1ozaSamnI7szOyYzUUPj0JXHyCUArllZymushVqrk9XgFVf2d
vyd1lr+IelZ2cHHlOM9h5a1oNcbsrhhBw++pS5M5Y4Cmx9mBWTpMy75q+Kbgd2j2
DgxPoJM5/YGLMZEqUF3AHiO7EPDQe/JNl7IWnikmXLoL9OlkpxoUUvLy1yhexj/1
mColRjQ55fLFK50LkOGkAejU06OzBnzEXWR1BYglpfnaqJPdNXBrkDiKzAM6yn+f
SYn9a3zHbKez6XXzpDD5cO2Qc4z+jjqLy0As7/FwZKrMXTRqHVA/10teDYLYy6U6
cehOymKH7HWOMLQNpXw7DodVtuPYGqks4lDdxWGGnLTELsnZyF6fnTjje/QPMF75
KfJYYpbmzAlNeHLbMFtgJvQ/AspEGmXOKUe5Zoc1is8DRhaePDEPkRdBv2mTn30m
TkWiemODorkMVjrsKQVkgsns1BvXN6K7TJ034kVsEPBA4HubKizvqKTUVgB1qlVd
+Nm1eOMY3oYP+IDgbOlIHsYV1v519XdmNMvnaL2BpfE9wFfIBQ/5Pa8ICuKPX07q
kN54H93UsvCv7SiSVW0Uw9JTBdy4oqzpsv1Lbgw7rLKI3//tPbrJaq0h3eA3Vmjf
9zlqxaPVbYmJPyt89kPglJWXaFFTAzfNJgoUU3qumKldfIDMk+bCSvCcmf84p7pt
ZabSfhFkFNaxNzssYcYQ5iC6oADGVJofbjqeBQKhAipVHmYgXHJDmMP8rD7szPTp
iW12E4OkKx5u8Pjqt3V/pO3KMO1OJRmP4DldGd4sNSUTZQ56yw2ZV45pp6WpUWlL
XEd86AQcippo1mXzp/ZnkBIuDnP9rMGvG9GgZwuq/Db8iKkY6L2etn8NpcrYwpUe
TjpAP3JQhrliQqNUMsMWp1HFbhTfeGDxLjt4OCShqMfm00KPAjgf6qxXz3GFpQyX
cV+GZVU9Zic4Viz9Nasc9Rm/VnQ9vrcwjjnVZusoZtoFKwoV1edoTtA9skkIAibw
0wIZlc/tn+yqXFLyJ3afVeRXufWnHaIFZqfu0qX5dimDdGY3Gwp9r2j6G9OWCH5S
rOHF7jT//xWcbb9A5c6RC+tCGvYYIvr4iK7oOvbd79ZN2ts6euO8kL6H7TNedXwb
CDEIAwTNGVnwT0T9V4jWP54XEr8N14Q1lWDLXxBdOGs/BWyU1zaPSHcGPdutnsWj
sF3AtBWBJbPS+jfXxc2xgdTGiYaH3Vcwr7ayL0aLkD45zfmonv+f+3ax8rkr1/IO
BZWhnVhs/WewiBvxhB8coiOCbXfhAouqiYx0DXM9ISkCUK07c8NYiysHrY4GhQqu
Y1+EqiG01KGnwo+cYut9OXTNXsSwFtNuw8vsrta3MicY5Ybx8lxL/komk3GnZxAQ
X1wFfQioVOutL4lNI5V5p5v/1GF57kGqLgMJR7obxRxyqzHn3RWaVdRiRKn8YJ6W
X5gxjMOzTbxWLrcGv0in06jdCQ/ELg9Vd/exn/fGrEdwxWxqvbI7xl1oZztyf27c
9RmWkLgPktiqiDsLrc7ejVqpbBT8+Jma/eqgT4kf6VDiBuKKfj4CHniwYRqqZfE0
cRacNZVIX0GP4qfInrBBIhCeleKzOjRN8bOe7JVPVg/BRPI1ZhpnEJklEG8cutUk
cmLk3AaJvZt3geJ14BIQHPJzDgWme+az2GXiNDFszgURe9hHb/i8S0FwQqplIulU
GfzLTFXEUnphDWHjRwBd8hAIUYx36VY/w7j/Fvvp9PapIQIcg2cu3YX2bxm1D1S/
sKN+eJIjxtNdKwSrpajGDeYhpoPQ5zzKvWuTLTHkZKvvGa+5se8FiEVPXdcjwNeq
JCznhVCW9EbS6xGO9JYzm16GC7CVqRiXKQZzvFp4BCRPtNPwR0GCCdPU+nkXbMMv
c8Iz7wfCObLRffJ330+9PHwgJaRxToS0YEtfq69Cl20J/yBek+brIEfDwe71tOyl
c6eiqkjqLYQ68AmuQdLt+iVUM3WWmG4MMh2q7/DwfSQZVVLDkB1yWEQ7U4v0AlYY
SxWuGTpfc9lW9vhNfC3mv6KV/yxBCr6FrZ3tq2SJCGABBSAuqLXAUlUoXKqaG+0b
aHfEahROlYsoL9W+1kfFnWD1Ku8VszgfExFfPQA/OWar1hqq8EO0ooxg0/1KfnfD
62UPozJM8MhPURXDPgoJ7yw7Zio5/GhGAKIsk+7qvfHYz2j+MRe2tH4f5L21I/Nd
saTV4cZQKwB+6CY2u5N+hSySFQZYEPlOVGn52W2CCgv+2K/hTB/Osf75cdvWwen/
Vxo04UR34siQl4dqnJNJFiKb7/1Rylw2HxsFwYjXbRP7xLodPqEiAlARPIcpo/JC
ll12+k0tnNYv3gPNk/fq/fgqk8trFSqU2xaZW03107jJWvh4yePfk60QuWapwn+Z
UlLKAT6IBNiWxj5gHgQeMB8tBb2hcnlXOLqvAQ196sGKfchIPQY7uOESFhFmiXtg
Xr7M+bXe5t7LBbO6d2+jmdHBVE431vGf1ZcTaMn31FzgjHGmwDtzBm0INKhpBZp9
CTLm7yOsKLUPwJggr3rToK9y2PWHRzsCSHsQ/UVXpfW1/g4Zzm6WrM5EU0MsXXet
JPMTiHBnmAgDpNhFriWtvxaj24Q5498ob9vEBPSSiQc42RIapLR034JmGqLEVQir
dkb0ier9rclg7WiFEJ7wuWSesaT33Fy3Ca4nRIN8DCSfdr4eOLZhdhreW8ics/7k
t1NFttOuH28AHG8yWuol87FgU/0FDBmHJXHRxHNluUpc6L2gvdI+QY8tMH93S7hD
icsqqRJXwaihaQ6AVmbIkzWfDYjP3PCEDn0TknimEQ4ke2v44Qe8tJIPd61ZVbDv
EUyrUSAucKLXaeBYcBfH8tNb/IJbjH0k7Rj5ZK+RrXCSonhTVd286iEw2AuFctYt
H6njZLD2afc5lOgfIQ3LgxLBQHH3GpNozRweHxscV/CBnaIVPbRr5rPdFqocplUA
dKCDUNH+DWDjzB9wTUI13rcjwn9w7xYit5jjJFlHewb6lHl5Z868HCKM6AgWvOkp
c4YUxMITuJTGPv4ZJoE+1y9UzmAiCzXQ9bV4XMOwAx1W3oOHNRsRBqGUMINzn8GB
Xm6/mBkJ6A77jXQVoGqI+SrdjN4sg8/eXI4l1QUCBJu88yxnWE4O6h+IV6GCXLZr
J7nvN4JGHu1suMQv28n1mSrzkjwAFoyIWe3XH98UE0rglhDKmExOhWzJp3qDeuc8
rs+/7WALkmEdv5mUZxQcmBmFCCfnT1eZsahr1WxnpqVTG8pfyknKAQCJQX4lnFZ1
tEnZnBnYaP/f6ucpGQnw8WD1eoGT9/N6+JPfHe3E3kU7u0pLXOqknXP4cAZthUws
sLSNTb1NZOqBnRnCUCi+ORUCIYa4m6SC/Wfja1aE6IjYB0MWmuIN7VfWVeKl25/p
mQDhGphbFSIVQHK1a8YwDYW79eK6u/qVmb1QHkeLMum0jvHV6PqllplrxCtHRMcR
gIwZKNTN5ecWvSUFs3mNAs3KFdKV7HjRKk2NSVRZObHmdhMOtxUa/MJcablvpoNl
imqneqWhEB7TZaYMYooJclrdUf2w2bBo/OkxSPVhsQ4mJnoyIN1+88g/MvQH70ta
/qEaTLvURu23Nmz980kemC0AQQR6GVwfWNDV8BP33MApHa7jib2ItXePS+NbyBtd
kswZJBusEexWk5VdBSeXSb/tx+MAuF5xEokIiydkGOhZeT3/P0bttHNzO2VkhZHK
zc1x+7KaoTT6/OWsG8dd9r7M37h8bfjZaRwO7TpHjJ+jazjl0Q0p4Tg2PlrFeuhn
RTsU20g298qs4Pgr6+xV29v9DrU/pDUIWTvZbYFXpfx6DGSKDbJt/MWyzJNdf796
qR/c1sj+iYm3DdfH5k5dl6MPXaNRC9CLMdWMmeO2r081s328zpeVv3mUrk4xAxjE
hQSKPnrOlCdCqOTJWaeCWxEg3mV2qQ0d1DzG2gZsZIFfDWcfKfTao2I4AnTwYToO
qfSteGG9R5zdAn8KWTll6jWrchwK+c0Sq7SrxMLtXcSvMAJLGzLkoJuZFWq3CuBK
7djIugvjRU5bg9va2+9HorakTS5zZOua+RVP81PsQoptRvHPEaaDv9L43FSGw5bq
hmkNP9jpCyxkf3t87Ssqncs0ZU3UgZ64yPR1zVKbb4a0V6AW6vSXKUrAtBvwn1GJ
8qGmMau8HxEeB8GjGvU7peFxvKNE6thZencbFuROnsuHateyXT/Bv7j2q2BGU0VA
2fZ0e3UH3BFq+4cUj8vYA30yDsz6iBh/eLhsge/7BBtLGzc4cxeck0GGMVl42ADm
zAQqlIQpxOQqzUlVNuORrFmtlHxAlKhYreHagCQmrzszVmcEiQnWx6A4u9+qkj1o
cRgZ46tdX35SQtjZBlru0P6zBZlcmd0mnpZkLxmpCZ77lXdNaQpoiOpyxLIDuWDy
84K4YsNGO9WMcvx+phsmNsq8B2GfcEgMwo86aeGiKT2UwhqXW1wQg5UE34RYYQ8x
eh+7R24M5PLx3OVzBKifkrmwa8PQ0DcFg9WHmcCVNe3NowZucF++6pleXF3xCYkH
+USt0KhyR9bBKKTDL3bu6OWiQOSzthkLDJ222DZ1JAnkcNJ+BnBNbxcCvgYQ4g0E
wsBLQTUYI7JIpoh7BM8dW3oNKFep9aj+mxjeg8nFThXutn0UiJw8nho0lsfGVQ+Z
7nqsjF0Ogxat6S5TWS2vhppsEltNwsA/KhOrVbXTTLlZV84DBbFKdS69BMW0f782
AtSspW78H2aZID79jz6z3bUsCIuO/Imn2CEhk/595zVNzHUSaAeH1zDadRYrmh1c
iLdXA75tfRP3jzUHgfWlPU0iNMjOwADAlcbVA8SDnmPl6JHD8HTsVlI1REYBPGl+
quD8UVPLTWzawTK9owFB+NtUQ0YGJ5N2O7dsIosogyZDZE0SSsEGINXXaEsqt/5j
gTzTaiccP2pVwQuZKT6A8kWdAZYZIIUWFw0BnRvn3cqCIKPfBat4LucucCERUgiX
PZPBW+T+EnYF8f/jPKxBKupmNrX0QQnRgsyrEdXZ7BlbWZATmQluifKpZT0vXLAE
id1iaBO9HNJWsz8C+W+ANZuaIPCQZFqS87+dzQlywsE69zh3sA/AoRzdWMbEUO5a
KOrfzwUVNvggF7Wf2UQPVB9VUg/wzkogpKH/yC37RgL0G6CIAtZoplqH+EcZmoal
1RePb7ksC8hYsDTzmrWRD5jyncrRBe4PdTHAqQdg8PHF82VzZP+d3mLsPxHIoCHd
Ui0gDndsbXH8EEPFsgw10twSVOMk+6LnLNcKs5gdwixbzIpyZA0lxZUKjdWGepIy
jsIPtwaPadXEob7hjLe7tjKeprTmhIPxhJmYfHU4Ivri+ZMGvGVzYVuR1knK7nzb
HfV3KswK0dmtudHshEfeb9RkhvoW+qP/mHUg6u3nabzNRpKXpVniWxMYdBDXSGqN
pNIH3LidinIBVn/zqyesfWDGv+QmHgKAVKm+lmiBfocLGP1ru/lFvG1soLevCC0L
7DWyMqImxLl1sIBSdxkLPdC96Rp7au+v0zCsE3wcUJv2Y46hh3Ut30Ja/3a9zbcj
bGwjJ3PRhLTRDM9jIBb4vYtAfccTjridsrl7L2EU4ta/6Arw5oIhy9gxD3k00Vcq
NC/4LkIB3t+iMp8VG9AfYzHk1Th/DMgBMCfw9gEJl8UJCd+Jdn5bN0RzTXWKuOB8
01xebi/887E+cPFSJOZl5ZUZCBDW5fn136ha4IQ1LheJTG4CBoysMgv925j5nHCz
sRrjQfwdWMTaxI00+2XpFiv+8CA5sU6N7HSxPC4MzuwvsCwgbttS+S2J7BZFuTau
BKTSH1j5swKttK1qE1lKLCBTset+O2Hw96T1ik0AuAHptken3pgYMzcoyDgqQ5dh
Vd5otrR/rTnaMZVPG5omdjLs1/H9e/IiRggKiB9bUSJlGHEnf+/RQx9+ohjeKYHm
phlm+uY1XBtfQ82T+VqA38wlxe8bl8ES6GUWlKttFD2yMC7KE05ANtsNWYJgWBQv
cxNLKPOPzVmIiWMGZu1XbEdareNjdDQP8lKnkDGgmzBZdwRgGKQ4jszNo8qRI6+A
LkoyYwZS8CKd9ZZxqBxXUyDVSTu0G0ukL14H1lzlE0oYLQai2yJ6eytn7T9CqgB4
qyU2nlq0cp5tiWshEbeBrKFxnzLRg4I5CwC0ixMMcs2Y4p7C1BG1IJx3Terx/hil
BfZKWpRQSXD66pn3fNcOwu1VZvqXV5Fn22skx9u/3sRzDNkO0h8u8FXyrKzAaUWr
LOT5wQWnKGINy3cQTlapnIvGFZvlJRqpKjPXMWtfWrWNSvpFSFXraxLPMkswGWC1
ofrVqa4Dxm9cvJObkBxy0OnvoYTzeZtpcReMJPYd3A40zmPmApF3Dh8kukWMnD9A
IEp+1AO2jVx4y1L94CshvQZy1LglomXLPb1IpdukY9obfMv2ZPfqX+VX0uymh2XU
02+AmMakltZxuzZQEnE0PNanLC9utZiMIFOhNyLReFbsgt2RsgjkAtuNePec7qof
Id2MdMh1nPLRhceaGVrSNdwRfzAdfQD5o3Q/TkaGdio7Da/2zW5VEAiLYS7n9Egm
Wz3Iqypxq3dCNVxNgKHqD267dQ1k6Muewhv5czhnm9yIkqkOkMk+ZXhmG0uG58tX
mqLeLhEgPocjs9sOkdGkEJ1KkmGeuIMboDiJcw3G2etMmK0MpfAUC3w4z+XdvnKQ
iU0BwxMextUDfBS/Q/GBCy8IlRLZ/tWEwb+k2kuD6fHfdLLYSR+qrMRhLYhZiSJY
0aP9mQ8WYYrGXQLW8CNcR9pD3dtmtKNX2lY1yPhXL8V9OzM7mVsY2pYZBp6wHDNZ
GyiBsXIFQYDFHmkN1mSKbUKYm6/t6VRINnPZGg5Wsb8EPdySDtQcLIPt14j3YD+8
Rd2odyi8afeMBTxHsp5kuLtshwVOYF4ddLcKchO1wGzTIYRfxKbI7i1KIjCx4y+K
f9Du4RpM4gajefY40LGoI0de/Uoa1AklSabVbZ7wCAcoo2AfUFlrk8nFti8jckTy
bYrLpTWlHGtWsMf6itPlHuYBy4gssKlT5et/XnlO4886z4TAyNuSwLA/N8m2wibM
Af4k37smOz4nbpm7Q9I0T3/LWHOpMkMx+7NVA07dD4bT4kShnV+s2PeKN9mbNFYq
NGoLJrjfQhKdJYRmqaTm3Kit2SIB0pOjaUgOpj8Jb8Mf9GG96s6O/1g5YBava0AR
LS3cTmHT3mGvrxvoflhji/jtgc+1lXs6f6aEqOGi8RPrVoDw4ABoQs3ZzDCmdJqu
rS7+3QOFSp3SayzuzelK6ihE7jcCCFVw27Mp4+7QjltLqjpCmOmDfD4RB5FaZJsE
OERx7VQGEgX1bHMGEEfnU3S3OvPxJtsmBOcUTcgZVBCVrEUfUExPF8kO8QLv1pVN
DgdKZ3L3pcEmkCFgdWdvA9R77VB528bF41d3ESOB0s9z9YEGOqtJyLEcECGQBWso
pTCNAAANcYwXm4ZvTHxlJryov+yBgoYHyEYmLUsy06wbUSA2lrLrsbmM5vsfSRH+
vQl5UMznsYHvMQ8agDtq4yzOiqt1EG2PsFVkVuQiflb40QJTqCXvcEYnuOzk7bqw
IxAdZo+ugTADeHRA7L+Q1K4ohZEQ3uWFiTUs0ZL09gWOJ8VjZIgKK67b1251unjS
etwUyp7D6IWKIfxrlEoxhWxHJRoT1JCZplx+4VT16SR4Ao1We+O2ZuqTFWsET7sF
PAMdIKeTV/HHZgCX2fd5QAMJ/rLEzfjyDJ076PKUg/0QMMqZ2hilFo/qrsSdMdap
5762hMLUMMZOQ+x86xeBePXRThGj64CRMuTeT5nBHu8mmWouYYvGM46qE7WlayBt
I3gUANmXT6YdvywdhtIWMsHmShqxnnDQ7dm/f91LM/CT9jGaAnZJuXSCBZmaWvWq
D5m/doT73qJQDK/Fw6OHSuzl+25ov3Y3eqqjXl+qwezRikAOeA6Bsh4OeQEkU8aC
xIV7lcYG4oW0qqwNyP54kGk5OfYvjscfgQ+CiLkoHNwZS/XT1zuyw2MksxjUClLs
TEKkdebX9PZM+wt0nlxLU902TzGps80kHT+YD9Bm34rER2rxyzfVWMAsomiqdKIL
NETNS1uFE7aGMoGwiLYMeHkDbPL5+q19jz8Lzi2zlZ4NumSduxQXhf4pLqZPiVWh
svrX5rF76xCE3GSgV/Lsq1BKrx2msP9yb8MK5/03wn8u5pZZzMb/qsPvkIvYVJ+o
3s/pdz0aeysurJBcCfO5OgzSwVeCAvCYF1IjaDBCQS/62hqeEhZ+ShRLSHptVu2T
M81eBXRhW1j66ElFyihSmEkYq15q8gSqKx0b/ixwUY2wE28cAHmfaoTSJx/dnqKN
DXVkeazLRfTJop7dSVswsjq6fWskAGoYgt9YS2fASXr4CC9xsWetnfnBWzZLmK6q
jVLwTKHj6mrK39F0xV63cG+K+uk5g+sy+tzpqExKjPpVkxD+Iav2dUUMIle+TcHG
D8I26Fw67AkYxD8W06jn4fFl6Oh2rQWtAxZM22yu5U6lPmPrj0pHeJWJhMGvlqUp
MJC1lpfKAM1xPb0kGlRd9av0uhjOY0+z12Y4WHNBN/KbZve5Kmbeyf4BS7T+d0MM
iHhnXRje7H/K3WXf2SmBlEJAwn8XwRORNgUquoL9ggv6FKxLnXx1lJPCN5ZVg9Kc
oOS1am23k/81aAJ9KZxTgzIQBZ6XpOpfBih0bLlgKX3pKE47VeBfblQUZlR+m93s
21YM4lUAfyDwcyj/GWSul1QlT4NysVfnuETqvHNKztPxf2k5M4VRk2DJK3dqzekP
8qUfXwgccFVt7geyypqgWVpBrXG06WzS1Dj6mykVIxcThWRHyk/QMQ6h/5imJfmD
pG1ci6p61/Eq2XzEJ6g1peFCg5DJkGx0O7mUEV7dyjU+B/a1Ht1ehElgvXcHP3LV
mUHzto2hSPg9eA34LFpfrFclGrIA5xcH1ga8q7m06S2tVdSpw9OKOiV1Sc+vrq4/
mLq40oObspBjQN/u0p/n55N0iueCWd7GDrAS+pm3vv6IsFSghHEDCsI5AfkH6QRo
e1WRALIoBRXxH4cI1r4DseBBMMMO3Ld5SKmCo22AzZ7/qXrCSQfHjcv4Z4J3VN9f
j+g/4swWHYNF13eyNzwCFWB5dhSfzT6YpV9Pnem1YtA261+tV/WI92kJHBFytEVs
itdVOt2QE6Ttlekw3sdb2gCO2AjVnLeW5PY+t47/BkVAGyw1a4yMgP5wx0Y6Whle
Dsn5XcvaYRINsfTnj88HM7XJ1omLsoCZwTNFQE1iRYSQrmBh5q7mb4tlDyn1oJKm
fUPoFMQW2qorUcEMF942j1chxOPoYhRx4FmbBeJgup+v86NrEiIKV+6UJwc252aR
TmvQijpoM2YybqsrTX4GXrOMZJwfTP0xuwbfQ9DErLnnSL4DD+JeSHUUkbqxwBB5
Rc2ap0UEMzpyT6GMykL+75SRzES88NlRIiMR5e6mmCVyvnoIyYfEagTGXDoXBGfA
9KXysjUzzjEZybiNDEQtnwuV6/1ezxXuuQcF3jLjH/9XfNmy0FoLyvijLqPr8Owb
qbIQIdl4jntJy7EF0O+Uk/bflycZUh3hah1IN4cl6AGlGALQDf18Z+W8CmS6zVPO
wFTvEZpJSbrFvm9V9U7+l5n76rYlec2VYfcFKgJ0KQp5YnjSSHimwHQu3Hr0elRE
r800AvMyY4sYGLkjTQp38N0pVkLiuT1WzErWrPWe61pNjusfbgEuMj11UasFvjlZ
jDWWu3wG6ih49FQrSWYlTIzjwmeR+2z6vMe3Mx1Ibt8pp0+XemgjaNObZiyOxkHl
pxVe0JwsqP8U4Ip+Yaxs+7pi7s5DebdC6Qj2Z9mswCtdNQOWSaJ7mxgYxShQYkA/
fcIJtoD8a34BdvWv+3gS3fKfdqk/D033tNpRCLBiT0U=
`pragma protect end_protected
