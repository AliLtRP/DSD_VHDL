// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OAthB/qIRbFdtWKf4BPhaQwNadPZj+L986IG9syrxclYBV5b83aIjskQJs+NLSBf
ydwo8unzjVw1QeDng8YrXEHybpd/nvedptIM6nufmw/hW30F81lofxQCJsMCp79E
J5LKmT6Q0vWn0ZsL7vN+tQnYSY3fc2oquymWz1zY/To=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 80720)
h6x7XauKWjbN7CL1bQsTH1nyDESiyIfHGtXJSTjsDQiGtNM6PeBEiWs4BTgSBN1t
UQvKbdI5AzgNkIpu6GHwIiWvmM47suIS9y9mgBwMzTLUNn6l95zDGWC3e8Cy0Brr
vvOHgvnu4XR/q33KLwHP5kxIS+CMMBIMW+6WtqAD9869JO1lK5+YZiktLMcioEpB
4xW89nPYRUqrzr9B5NQfU/0sO9ZOiFrfjqsUtGt0BgVxrSah/0zZbB+K6Hn8nOF2
q+nYuRPdNonUxeRp45fEkrVdimiODm6Z/dkGup43I1awsQ/CPXuVyQLo8+Nie5mZ
eGrQqvH17j+45+XjQ6iBSmUE1FbmvHWH+QrgTFadwiIf8G4mh0Z3Ifb/gBSyVvJ+
6XsrEhu8kGl/5XIlqotTdweFcL4/bRnHUiR9DkHhQIBBBESIlnnwR6mskKxzA6oo
XREkjtEr6B/KzVQRFOV5fDqJjM7vpkgXUrQtr43EY2DbG9UNx9DqHl+y9I0vKR31
fs37YENnF18DHbXm0KrC+PnkRIfg1vIUWwb+h3FjSPOUyOx0VRfncYtlK+i6hBHy
B+zhkO3Hvj3y9CmoZkuM3NCwjg2C3hEf4j+vRLGQ1Zv9S9DYB8Jvzjnh5kcMdNAa
b8vqwUfVaPS3EQjIWynwG+BrHTEMuDizcY+NNxPqICxsREAc7f1x/A4ZOwEq/Iez
Zy9qdCS+XTVGG27v2+DWNFH4xk+bImngyG8ppVYuq2RAjiW3hFf/Eo+A1Abp4zdu
sa1uAPxlnZbBOqTYVRxCaYL7jRHRa2INscln1LKGLNNZb74+acoJbMn9GSfZ/eUr
KClg3KoTZxDEqO0uEdX1BBbstLebrTEzboeE3jSEPcTBsS+n51ERMtp/KG7VFC63
QX/QTwAbGoBFFlv6LbSvbxUv+VSJ6nq46DKjCEnK2/6e2Yzwr54hBvc0sMlwe6Vu
U/wa9ba+FKOfEETAFly0Wnu4xc3h1mYVLml1mF/lR4kfLeAPWATfVT1WQcnnw1dZ
2X1q5nvptIRvE8czWiyQ199H6AqUOMoyWOfL07gx5Yyu4N1JSc592f93d4L6BDMl
NTvka6r/PeRqnGNaIw2fZ3Oa3z0rwua6qnWDapXF8PKX7ZgxOc79qXlv5PgcDLoX
0JcsbuJmOyzlirMn+2bIFNRuvABrI6Xmx2231nLtzMRmT8GE4mPchpRjF5pe2QkI
XYyl4PWNuPOSHIySJSQ/MW5c5eWXlE2Zmfh1wTPM5YVNrr3Ln11YwYMoSISmHjH5
m0mimebKXiJD4HTnvVIqVoqaQWfCe3nWixV9ckjh7qtHluppbG+PeWm20yJSQ+FX
gtKq9kP4QoVNcqYlq/ltTvAB7yZEdHAPE/enPuWh/bdmF+yVwrXi3oAZwmEGmHte
mIVwhZsyFW0hI84G6PKZabJKevKEO5pkud/T/rRPAYfGP/FYlRcM2OACPci5WXcu
h/vP3IZzKZD6WVzt9+JCXsRte+8giZC9PtV7tA2oqgTXc36Gcep9+hTKZPnbbK/Y
7zhcrBCEUnpIhAb2CGb8JSTQ7x8RnGTqWsyM0Ho0JQ6+E49PY6FOaJY8qw5qbotD
uCazj+BuTTSxKW9Rir76E6GWDrcd4ab9dpP2dUDjVRj7bdQpq2eT4OF6CSqKZFCu
QbgOfQZlebsThcdvqA+9nFK0k30QMNU556lQ5SVgD312Cns+pKHGE8ChqFdu/J32
rcGNelewz4BMSDFIu92tDHOWcXYRsfSRnzhzBsHTxhZS+82oSRzfQbLD+XgCaUa/
sUXwUKaqXxZwcT83RHii479sn26lPrOwzfJeR4K4NtrTzmNpO0bKj6f8rnGj/RhX
5fx7wt4/9akGwSvpZO47ycM8xgC96hx7iIc5VV58qys2cyEmzHlG5c7MvuApQz8b
BbhZSrSBEW2HfPG1J4oSX7vZVcFBZapHbjysVyBMP+gZ9usFkJZeV5x8XRbHKakb
Lvt0w1z6iLZ2YE+7K6XiOtc2jml3uHwMHMSBspIcQfoZKIoJDthPfdivuD651xm5
3dYlq7N4qxPQavMSlDWu2h8vNkEvLPKQm0ta+LhDc4C/9UhK38wg8a6gZtfM/P3I
QYfXLUdVMVDrzszF73AwY+1LNFFytYroamK/yspqFYH9E3fxqVdeEBEZveTqmXQx
mEVTADTf49ISckOmQK0uhZ2s9UOG9fMSAHoxNYJO2fUzPsYVDR6skPMjSwvbqQ9Q
UL300pPc6Wfx5IsKkmzwnMA3c00hB9mQ6NgBlHJYmVty8mwZKlJY7oaHtlVO943U
Jd1/kwBur77pcTSupzbBlw0VjMdQXTWJzrWTLrKYmHsCk3Y5G+6MSy/xMkihIQBI
+Ua9PF3M9UWHIxkpfQ+6Jrihlbgm4a/tp+6RIl0f7XncAmwlhtsHbGrP7nujhYCs
QYWBbabS9EzxC3Q68LR3zPdNyEaFu/3pXwTWbD94peGaC0Y7ljqzWluDfPtrn9p2
5SnHNM+LOn1/z5iWvhif4uaTRIx/adZYTuWyTszhjhjk72sVbFi/OyXgl6W4HvQV
kANbS7CRtOoyOkHY3Jb4FP/yZXO8pIxwSbfEKeBGlE0ge/vUixhUCqDsNd+yGkI4
LRQpx7wxNhE6/XQPp9VwwqXGktF1SEGTATYoWijiXUsTIYliKXY2ZKQwWEu2IlI5
+IqT04fw7avkqTBCKP89dRsap7Lqb1dMhTkWrjPneic1Y+aDdvr6p9ixZffyiSW0
7btYvJMbt+Yh3bUJmjVvCbxBVO3mhPMvxaH/WS294DaPZHJn6BWZSa/GnXJEtkf1
+6kigoLr9hwZQmqrpFeQukTMGhBcIngtk6I59TuBeGaFWmdwe+BgKBhJI3jQHRV9
ySLr869dhTARa5rtNiZfkJKXo+gAI33vPDUNK7XzX72aGTtmkn9CMVP28JYTSgN0
HlOQam43/o3thZcFGj8ldpZ5qYYQi+TcFrsEkwhSD6DRDZZGVXkM9Pf0cuZiDuZ2
RkdgP/S8PkrXXX7+OkreBeR9eo2krkZ/TmuyfTVDewUYkUKperXMIxZnCeoBgTqC
fPcu2O/P2sAUwYerh1azmzLar6a+09J2fnoYn0ItkZBpudkP7e0Qr21OSehWMG/d
EH95nwvj+JQstXJZHOcBVe2tdZEB9RdsJi//fLyZQLjZsc1vKQmO4pZ0NcgueugB
jhRvAXZmOBRFFcxAXj3uSZA5U8drkl/QIKALsXU51mbMFxmbnJvuviKH1bSHohnk
vreMPbaA8EcwZuuAVvLts7eCpK0PGfiyOmLvCp6MN46bGWujwuapI5hkkYb99odk
r0m3v8BuErBOGI8oaX4xkubTihUkRnRIDlcTGT6vD5G2T3VtUTyNNavtg6gotMUE
i13BLQTBOyyZc9mz9YkR46/r042wNdsTyeWMr6X8ADH2IcPi8TId0yLmbzW5s0fr
eB83Dl5NgOzzUJ0NHjd5ObVUoeGBRJqke/92ZuSc5Uw8RN83aJm5+Km8FA3rMxPL
TIlrrRmmciaU/IA3KmE1XRv22tHmmbqgove2NOOyVCL5FWOCFVn7tMviNmVR+Dzx
QHlgGzcnoN2wJnxnE4FbSVDSsZYyHUa3kg8Yx+3RW9bbvhpbALQkGE4rnCHLPfCd
WBlMlAXhzfVUu2STDcCTJd1oMpi4AZOUheLgOqHC6XFswSarUBIj7SA/lhJkA1ti
/wmaRiTEpzy2bjGWyOV6AtQEmhbFDN9+vBwghMzdjquDiOwhm4ApDzRTtr1A13Ul
4bfRbMV5BbWdxiCmfloqrjhGuDgIq3+bj1bFcCvaieG2ts2mizGnE0IR9SoU+6OY
dk+FdoO/HM0XJjTWCfi7kpoPkHF/WtF3caBMzm2QXwhpkPaxiotvjMgOiT5shYIM
FspbH5VGxQZWh+ah1a3UxM3gAWKxWiYeG0Je0TIRYQZcmu7z4FxlJc3HQxx/rH2D
SoMnIYArWnZuO/BBpY50qcQZPn/zko1bkCicGlRYXyjk0+kJS/4vhKaLgdYrA7sE
9BlgL7YZjbbdqtWFcaA/fk2Lu9oRxFQ+nUlHso9Vg3wyxmoee0U+LojNiCq7kktr
3MRBYb1zaXhF2sxgyZnjnT7hAR7YK0unL999suCEmo27EGaeScx4U1nRdEd3/EBa
/auYQ5V9BYZ/ZN1eqOXcfthwpxSIU21ahpnSDzNOiTOgpJc3gq7LQCtTz85oMwDm
UoY68cBi2NCijq4FXm0t0zrDdj8B9pEWNoY82D0HZ7Uk4XsORj/vMpFZJToMmdsp
0Nx86Y8GCnYaYDppPA58qkL3yWF7T9bT/vAYR8Eas+zeEMYP/WAYRuRlhQgtrbR+
YLQXpvv1ZHjtx26RoGQvaLYWenfs9Fng2EVhl5YK1YH57z64KxlyYDJFTOFlQrC7
DQwOKYfnbvPzYC1rZMi4CFhNcPx02wpeeafAVhWsPhjSpam7impSF3m/7r9Y5CoK
nurjjRVtK0SxGUeWEd9pqzTmp/mxrGy8wHEl3Bcpa8KfgD29LGGil42alRIO2j1Q
geiDBYTr/AiO2/e+c+ITVap+mbp45iathWHZsuG4zoTiN3u4S4zmC9P7rJb4PV+4
YAJNnYjMSqklThxqA7h1Ivzo+TXtwWVMB2AhA0+vtD+9CqU/5lfDuHdkLQPFmXpM
w2eZfe/QK8p65yFiUh9XSH5BJCKG0LZ3Ha5OcbOvk8rdtnHU0y7mpkCA2jvQSaHr
WnmK+51uXhseDsKCRpDJCi/t/Lk3cuDI4zkwIrBksml5MiD27OffovYDyfo9v0QY
cC+FC4kcCSZ/eC23Zz8R84xCHR0qP7h9qwij1h9j4vF6IV2itTec1lCRUv4zhW6C
uGZGbtyfUhzye/GkVaTwKMieoQTiPfaok4r8Gtx7QYq5FSqJRaOnQ6Jre1TpKAv0
3PpUNsHLCaNSttz0s/CsvuT5oSgPxZBBK3r7RosEQLdt8ZkoDse5d2TOyBc8Gb/p
VZGT2js8t86R072ekfgO4wu9V5Dn1XDfSdErRm5joSTj9WRVJBBlnMv4pl41dN33
IhfZcjFutQepbey2SBNSh8L60dA0jwekoa8IzGq9cGCamIa3uXRW/XoyD9qSwHtb
tmdNL5X/1n6wgYz2UwR5Nnvuv2oROoTAo/FW7PYaYiM2t0S/qzGrz+9jk6Is9KCo
7AltRcTo8AaXaXJN10BNAzCp9V+ds+cGM/r2+BqWi2gTtKnPArKfAxsi+qsRFbK4
I9VNU+L4Ygr/McewL1QP5CPBaSzoi+Z/yVHM/eSlurtyXdxNLk0Wno/Nsd7po0bx
vkIxjmW5DIbbjWbiVWhUCOJwQiXgyg9LHQyLTcxMs18FnJvLRKdb4Kk54lQOTx3L
/xDFZqkaCAvYc1HdEJgbneFkskWrrZr5eDTLmHsJk0YYmIh8DI/K6KI/+zSsv5e5
8J2LTETaqEexl4iRrJh+W9N5IyGTBf82PSFdAJFE7IgwW8SmRBoeznBVuYHSTQP9
UjCum+VZbD0EcgnYKf1Liin3rRKdkOnHa5WZGrUrgR7jh1UlMCTUYmY8Hsg9W4Um
mxk4Op/QVj4RGB8IqWtznQhn4FlG1WY+6XhWUAnIAY2r0ltgHpeeSgs0dOYdJReQ
tHSOaGVCLh3WZLHDRX+6wOM9oD3+wlh7wGp0BpKiD48PAObyWi9mCsoXS0ltiX0w
J37Ben//Tx2jPEMgvDM+Sp56d4YuB2ycXk32ViMp06Acs7bZ3b0iLvuaPcrXMPKL
OtKRkMEA+ifBu246IHifJ/BQNF8fFVabLkUFFI7tFPxdc+GEcegzu9VYnPbevdEO
CW5SrfyBy8zjmbZSNfB+LG9K/O89NiAeRkpQrdNHLzUCAhlRMXaAN2ldSEXgniEr
1LGTahXg/AUiK8w0Jyq7hhjv4eWSt9RSYgIMsZOBQ8olmixCMsVi/7KNJqcRvCdc
ypyNrCszboovnx4HPHjB2Lb2fcpWDYaAkLxahgi1RWInTOj1dpG4CxYvenxy4sEd
OuPYmB4LjL1K2UkWjeZ12UMdJo/LnXcclPk9it6E3PxmPTJ486XdKGojVJAZMVBc
70vsctG8BAsvy+Nec29H1hncn93FSlk0Fz6gnlHPN8Ir1quz5gn+l7njCfK6cRDf
UDU8LYiO2ob4ZOKdpVh9gjnzFJAaa18I9C5jm2bCQgkur5hrXuNmWCFOzqd7Eyn2
x6lGVXPASE1vKVxgDLnlZeteUqORKaDweVVMfDNihEv4fIQ9zIFarqRCtd9OkVxS
vaTIpRwzWWZd1xJIAo2CWFZnmrzS9rJTmGuBtWHTzNIgW+Z88WIbrG2/PcDC4LwL
TNcjjT0lGWKoF/CnrrDsFIJziGqqEqTWIuIl7hmPf/lhSGzl9elkrONEZgaiF37g
ADuQv1ZLa5rKnNu/j0g97v1J0ZtREdIF/We1AHliO78LGFk/AjUtYMwSpXkqB+GV
5FCfAhzogsJ0h9FrKxpwqtRK65tDlL0+h6DuVd9aon1P2/q7xw1GjxAVq/H1bPyy
SkWcovcq1osq50E15ZXJRmJ3gASiZXzEVqILhhPRYD7PLWA3Q8CLdUg90lVmJRNx
X/y+hXekTRZTW82TtyMqxivzU6lYmmbjeB444IQukTNKpKDLApyisSwXsBSOPlB2
rjtGRJRXNBXLVruRIN6lwai8jHjpRm2DsZBxAyJpmK3hJEwMGt3tZcAT4cG08vUM
xnVtWYX3AXbzCKp7ORV8fDdm3yAO0YHvsnmkPNw35ydh6J5Ft3LJP0BsekPtAn7z
F4vD0lraEpTL49sujnFFGc48SidYhulOEFBLrPUUP81agDemLzw8t8JWe5JyjCWA
Upc/vutueoNqsKI8pznr5pHH5B9qK9EeI1mhkJs6zbS9Q0RnWR4fKUiCeuQUAFE4
35kn66fpfIWKjegusLEJFkazTt+0QkME02h3+OCnmAGA9HoZxYjOWSJ9pf//gahA
admq6/d+bBRFUB7SJu066vA9al4o22pbkcoco2q3NzZzSvANWulRH/D+vZazrLzH
MCnGWnKz64uDP/8JqyxbbmJ/K8sLe1mPQzFS4VH2T3gurUYax7gdT+tO0SEAjX9S
argF1qTy5FPCcJaXEoWTLQDq9yEt5EGZVnDXJIu9umtEFLGYL+ph2YaSDYoPwqkE
YNtRVVjU5s3VDctO594oi5FZqyRl3mdzLFXG4XQU7xYD69QYCr7Nic4HYUiCSL2w
I+UBXW+sSKoPKjqV0aZuSecjyO8HD+0f8ZdtWojzmheFtL2CVPnPlNQQQcZ5BwDB
Df3Co3+dIMind69TKenzmF2RiiXC29Chfkaipnk9n+a055t74B8Qyfhw9eoy8B/U
cKNM3YaB+aKZM1dLTJoo968ibHgefREMWat/EKxFFIf2d+R7WT42LwYqkT3cIbhh
wiA0fFAygmQip8trsfn7wETPTCzOcLiB77XyVYd11b91fdSeXrt0mmm7EAMLHdmX
yB3l1bjF2jJgj0SOTH3uALc4BUwGziYPKLO4wkqu9EFNSAyXf1pyyetf7MJAho9g
/rpa9r2oLA30n/XW2nnpKupKH4012XKemF2YEGYTeUFvBW6KiDylQPUz4maSApNg
W1YxsP3sDQ40eFDM//YLIHNOYle971YkhICULcDy2U56X/1A8cKmHhdixcvi4rkG
JrdfWyJ9AijHXZ/Zvj/nGnv89HaA8SJsrbk6k2RJR60ljZN5S2GwyrPJsVQdmljE
+79txeqkQCzTVWT630tsH0rNsKpe+3qhNMnFEbVr58+cp5MXfog5IuhVCh8Xb31z
Ep5eqbutRpWmbecgO7Pshum7n1WDRD+q7NzoAMl7oyjyVJnE2cO3VCmuxnYA68eg
CzgAenDCEsMh0A9+I/mDkppsOfiL8NrDkhQNZPuHuGQjPU5YM0e5ajuJLILzHeK/
b/wYXH4x39HQt3q1gPitCkpDz73dkiC6qlVLhqa1papm1iqE91WhomEP5x5A2qdB
QJa8TsWF+3acoTCGbFawgTT+mkJnQs7ILqISA4QMtFkPOIRFSA8etlBu1VwXtrST
cdbaYQVsQwyvZJJzuc9Ei3vYTkzLBdXoPidd5Z2kkCA657zi9pdoXcunF+A/wTc/
jY8AJ0Lj58P1Y3Cuj39LdfZrKp2Cv8dSyowPU2+6w1l+w6mJSFlrtejaCnrUnGqu
Dv36c9oglWjexyavep5hHxp0w78A0vp2FKaSb8Zx+niAVuBkZDBX9GkSHTcyGTZY
MtJUK87Oh6wPrBgzVemDrq2InhcYzVZZ329nhCLYA/RXv4cXBd6if88L2JthsK+V
16IFHCllgi5bVYhBi8IqhHBGwdgX2rUB2vi268+0kAwtREz46ko2cT7Z5Bpl62Fs
vF73WR4Q4R2ehWqOdW79wv55E18RDxJZAXFU/CDGfM39/UnPUTCRUOYnAi64BVk1
ADbr4vyu3qWYM0w9n2n6HJTIQWZQyKXC8IXS0bmrFmt8l3Ms1ZWY4FVF0ZToD2k8
tQU2gS4onU37ej92ln/UL5AAt61npFdSLsyE0LhFPNOernKa97Fk+T5PRZgbV1bo
IjiFJ4MRsYZOhTgQv93y3DTvywM8yrmsaqiUrlaBJMzNZir8NRvFzfAMKzHqJhno
zmvhayQm240larN4MPODPcE9y9yiYaC9MsEPtMGrkw1feKstXV702IF2oaUDCsaC
bZgHgNxfCYkm4mrGjUWZjV5ExsJ7dib7ySW3Wy+X0e4bAwPhhPIOT6r/um4vTGGr
hz1gr+6ycNjlU/mHqNMYqcTyNzcda84G+nJaxTP7pm0rkp2xnHppf+DMS2PWhq5U
MjK4Umv0SjUp11++r9Dc5QO5J0cpNeDFGqS8CxAJ2qUHH6YJNhjv+cj08HnZSAW8
iUh4jgCRS887W4aOIlxkcLoYkr0uWieJCWDhZ1hkpSLMRL4hWX0x6ZrWKQaUB1BN
SS6aaMs4Y4xQJmwU52zW3QerLWFlaST3d/LKA/FMNa4YyDACSGTuPnth5ATM9zyK
DeAHA+t767qpD59jzvgeDHZVJM7wwNxcsCcLw3KFcZNOpQWQvQT/5g/20Pf1mXbc
R3/tdCHyBakkQXjqIDshutaWBxz8VR2EgIa33twLJAXF7WL6pcizDBucNl4k61U/
bY1na6pcmjgJP5YIoW0ECXBmXKCuO0F7htn5nb5fvTswQBJXPMSx3oOzYitud9rW
Vp6vmRiRq04R4pacTVJwld8vC3My6H6UOU7CuwPOAq6MXhj5Rtk5qhQlxRnmZuqD
Z5/4h9XMygk0kFZTjQ/m/ssx7UtItxUItpb8jTDIkSGAXaJWb36qeWIyAHDHB8nC
PN3SCXFmA3OUyWCYwRl0hcDIepZZqEquQ9pdIY5Y3lJrU7JwxuNmTS5mgdilPAvP
gCV7xM++OC2zGVHhCBTXyAMPdUczKOTsIIvD5FUK1C2knQ7OqBzg4o5IS54sTJ8R
T2AY1b1z4ddYocMDIPtWLoCbzXlTxeNQYLL84jJmmog4+wbkbwe3LsrCfiroFlzB
T7ccrIYmXJc3Rs4zMrerg+j2d5lFpnIFK7KCDDEvEgJbjixr0weHhMftMRCaNx07
YaKwMWENcioAX0603fc72xEK83+Avb8XMSezqM0mdLskhf02kqK32hCtb7rVr0nI
etbztI04iBnYHq2TQK8+IJARpr0f5341H3RbviTlKCm6u3Ff/pDvm/Aw0qF+PMlU
l2E1SutvegF89Sl4iylGbJ2fhh9a3W8Bp+OLsl1KmVIEVKEB2bxHbvG/Hb0U+4dC
AJO1C8nmccGActxL4Zj79OFDDWb+ZQ5s7AnP16UL4Mle3xpx/mw9ihrZzlV+9BZ/
vq1d0XKd00wFQFmqL68/EU+VZRlSfO88rSHzKs2wWrKxFHDiYin+cPIeErk3SPqO
U6i+OG53Tb0wIu7GnIHr6B+4q0mnCsUxT6XwGrByssfu9d85CeRF1yIFSeRKubl8
jRGNKTrysXwXC5+Ga4JkRjuQ13Pb5BUZ/BMcXd1cq8s8A/nBLNl96hXnWN/Vas7i
T59vqtIBcBucIHcORmewZKUIBYS7Y8yMIiVwxpJCNB40RYF/oyD1z5a4Y3hN5mhE
dFDmZfQfoiZL64UC+hd0l2rMJIq/o+xw17NUzPw0/PMqM2Lm0/jAgDPpEGm/ph/r
b3WwPNYxJTggP1PZWKKaEpVJu6m2CvTr770/iPSai/jX1D/Sx/k77H8bCAWDsrwZ
YCricKBAwoE+NjFxZrXbUXD9C8LdNftkB8SA7s5unqhoouMXHBmit5sPyX+D9jpY
7HAGcpjAdO+uGFsJYBKtEcceXKxlDcC5E3emo4fm8qNx7yqST9DzxutSqWFXa+3d
bGS1mckfCKIqhwSjSZSyOtXIb45XjN1TygvWabVTO61ZfnxwAEF3oryNNP5LTggF
ee+s1rJBWcZtuVqMGOSoVFgXVlxn8qo5KxNmSlaWB3C5hwVqlbirAi250XXeHr8E
uDzl7YcMXcPTMiRn4YRa9yaKsLq+v2KcOhNLIkQHb2jXYULwYS1O2rStK9SGBFmW
PUGYdxwTZYTmh1Lrnn0G80eudAcYYEGIXtL4I7tqIiAa4mYOvCEQgn1QNjG+x1d2
ripitszRoSWZv0PfS8e2FfHUTNarPpyKCY1QgwAOrMi4cLwRn45jJkXX6gkLvnpT
cBBmvJtaGHBuv9GJX0eWKhgqyc9QM/RFP0g46L5XpiZfyJ/lvzRHqdxNgq/gCbZU
EpVKvKo7oLfJVrBWY9rCq61frhQSngspQZqS3GQS6LBjZxF14OTkOhE6lDr+vlRS
l48K3b6VsNM7aXNnTUufmwv9xwMfAgrLSlXv5zfrKYe6XGD7DvfqtcftLWxgPBi5
83QYuoEj4J1PQh2NaEPH1CoeOiEorsRIGXPBOy1hJ3TXarZ05KAf7WgrAprqnnUY
r06qV5NdLvx6L2c1TUl3iiMeAc3Aw0nNdLKgS78rCrvpuJ3F+bydedfxugutFfE8
xJ4N3zxhXLYFkG4vWo5/WmS8D5BVsZCV4mssPeP4R6cEID3hZEgV8p6DjsoSMgLc
5VZBNbV4Fqgtpgrir8KFxbHkI7OgqqJcQHWqvfIljti8y+PA4/+g7l1QbcwyzTWe
YFiD5dZ6ZHw/wSf6l1zaZgnr1eyNIKhRPbTYndPu6gqGsfp4Ec8nKYJJeCc7EwqJ
LEA9C4RhADeR0AC9r/MeHuQCHzqzZZTMWv/C6+kmAcvAMF3nUhdWPNPO4UqQroko
n8LmehsV6I62bhPIQAqx8WYdt0zIrqAexF3CmWZeZO/qxJZ2fQtxgkuZtkL0PTGH
GSWkX/rGjoeIT/lFgD0XMt5UmD0m1GP6FwBYvoPalYVbqEk2FqK7Qboi+csKAN4p
MhAm2CFu7U35lQCCzB/0efpK3VJuAHYfMu8EiVue14z7jgcH3wEUDS7CRUMswdMh
ix8KEnOb/A3+Q5OpVYqD96W3WnNjNEJp3i0xwTE2qpoqTPTytZvoekNw3VH4+sFE
9p0wL/o8eoDtNI63+XBlDNpeoYquzToiL1mk4TkBMkyHCCDTBUTvMqfbODBNhND6
al3IZlGs1QL/H9wQVIjfZWzho0hDqqF8P4MlNXLAdb3blSb6ox1K052UhFcREdyq
WiL1lT9XSqASqft4aQh1zKP5AOkw7y6u6CJ0p/x4YPKlvOLRCVQTeVqOhmmXSyVh
JsAQrXTVs452W/qc5eoWIzPjxpSJXhLZOghuEA+4NdEAyY0DgZ7DU81f+r5Ioyhs
875JSvBlXuugpz52t/5vlbDp13IY8eF0lx4cQ9u3C7ovLxHa21MNMVvwfmk+egmp
G76PcNT0g29CFAw6z9blDHhUlvByuVGkrgVs/cwOTEoLs1SkMQc5SlP/MNnl4n2F
KPr+TjfH2Ukz0xC82RebdoNS83nb6OqatTn/ud4h8zo9g76NyxeI5AKYyMIjHZUu
zFMMVn2TJrnHPD4VnFD2RW5simrLzOUNc9xOui0l2ZkiwZf8LnnHm4/qG7vkuXNq
YCUwWRqDtg7u9LyKVEiIrkfs2wY/0F82n2MEXw2FZENbAta+TZ7G7y1sfIa4fsai
C2CVHH4fxbWOFmGc2eTplibYKyuGUoGhvF/IM/a5PLKA50eUARyogjJxxqvKxMJP
y/NtB6iRsboL8rAftIH/iOFWfneO4lm8KuOm21zWrjS0x51KEb/S/W6sdIp2zA0Q
A0WiBwlPm+4sNtaQ6dGDxtytR1vJXFOfIuWi5EMotgX0f8Cy99iSvelrBKPzrTds
QfJpeudX9xTnckZUnlhLKfuTtgxVIozV78yE0yi3OLFoXEcjxRRS2JExSIgl3Qmy
dR43IYYXwjnXL7lHzmfl1351om8gYw1SeBub4jaBHNsZC76wqyDM6jK8/Zxx/CQ+
3xwV6JmOQ3bVESKVuu6Mo7j0D22NwpuePLzFXdBZPDh7QkdSXthbZr9TnpwA6VEs
cC2ga+QcNSQp4PEb+4BFGBDuj9bVcooUoe9CfvNX5PjGzqxnzMdlrrZ+D7rI/vZO
PJIEMi3xH4bRwOKFv29myr7c426mqa53SNnw03R/2l15Wz80INhgLw6T+GJNFRVO
Wy7pGcLqf8JdnSW6+6SCRO3/PmFBYfyYQtwqDLACuH4nw932NN0jAOX1qgHQWqSC
LkP5mMtURax+H7ReT4ewbpfe8yGJQF61+6g9/ll3LgvA6KdYBZ5a9iO9v4lqTbRN
OsNX5pT7+UG3Vn9gpjBjqP8SDmpASrYm4RI3SNSpqnTb6mzqw6gtzQH0gVXE5DCE
pWSmalk00lgWPviINosjaeIrIboYZ+U8rcz3JKP2DlGfnflGsp04tNTsrNpvNILV
mlzrOpqb6izuocnmcuUIuWjp/Ux5UpahVjuiNUwpYStMEXpZgHBmkeE2vMEVxgvp
8N/mIiMuE8D9pEB1dvOzddvqdJkofec2ZJX++vC6Kru7HLcTb716jzCLAtv7ZJrD
b86sWERKwGjIVT/XLcx58Py+5TmMKORvqFQxjhE3k7fo6ymFiz8C/qln+agmaiNM
CIWdH2NkEar8PCoKx75Wrzb2mRgQW4trhP6Is3EH4yeXFwKeiPUZNpzr9vOGAFrk
xbJd/r9wZyFSZ/66RlDMi2zD4gJb5l35GoiDcoUAI/LkpP5jvKSBfbzLp2KfxKHf
s//noUHWpzJPFqSOtZEHBcyq1Qns+PXWxkJeI0TMKbacuCDE05gxyCvGs/rGwHE4
s05kJRPRZA0OqzDHiPjV37vNcVMmaGwLvq1lU+8h7iLmFevEjTs4a5eNWhLhu8Qy
ju8UqjtgBzijUFnkdBSoshNS/USqJjgFMOcN+aXOyOjPvfCQaBCCbISCfhgLFspw
enOaSK9mfFAcItdEFdQltdCy71IELKQdw8P8NLyQIoWoZuQrtQcAdlJSMdWymw9d
G6ntRSBelspTLq4pw4PiH8DV2Ize9e6Vx5wQI2hUtkI/T/5vk6nKeA4lEo0RFQvk
M0WYPXMWI2G8b+jJRodRO6PUTiURpXy/Cj5AyxITwPWoAFsOBTplGP0nIaaIwXub
id2DWdyAmDhHfhWXaQ8Xob6DmorkQVZGjE/1Onybt9cldCr7EPWIVt2G8wLyTfLd
HoqwyUF458Oa0PgtHpPLryucJKCczuPXleKZ6wftjS34WVwvhcyDY2XsgQi+aPCJ
2jSIuRXUHwIi24MSXLQxEQz2PZCn5H9dAbJ88l1ISizTsvWng+xATPqz2L2+mdzW
vIBBV2WPZuJVYCbIwWbNQaen9dwrVSoOAthR7yKGZrwBp7U76A/xfRVXgm2p4zPw
v+STGi+P/YR96ycY/GpDTVNeYF2RqTlC3h+7oCEGf9ictl2w60f+by00oyOTN0Hx
dq9hADBZNZAHNMtS30KGGGodjlLg/PpdThm4+JyKWJRnLZmgIzznIks9rXBtP0/A
lX6DPMBG54efHYFNPRWSQFH/pstfEdAW/pFWEuY1anzm/G+Rd7UPZzZxfpwhRtyW
I51GJHwRdF5oZAdeelYUexVgG62clHJQ1QB7jvHIzNBwzlvF2G7evtYQjjlJw/6E
D4h2Jv/SEwuFWE2D5dFaDv1qQ9gSZcdST8U4glFWYrj8gfkUzBC8xgC5UMaW2zTG
rxiXShJXxbZC5j4q1v/MZWZ1ZEcwUx+FmEk2K7bkf09/+UuCN8jgoywIpqVD0RlC
G0eZs8iDBSYry1Ih/M/lrRiVaYqauokyiAVoGUJxB4pGjtXPeFDMg3vQgZCynvQG
mTvU3vHBd4UH+dN/46/Ksurkw8IPfHtP4BTaSfjhI4kuGW7tkx881deFZwVupBTr
19vUCjedKOI5b5mLqPL94y/uqi1ArhJ37SZvWtSPFysUa+1GuWcNayelF5koVSpC
sJ7MMJX1uGAIYNnAOOVuz6ekfhYfE2a40av2rSquwXgW8UAcbcUJ62QWC5i4b5DV
IX6ZBSad5pkcH0Tz39gqoD7r2dl1SV/+V6Ff2a5HYvfijrRdB3PV20lGkp5Tf2QH
z4e0NiUh2Gm8tA6BSV21DSzcdBfUqrnYxtP1tFaDzQIrmKsSa1jHqPYrN1dNxpF7
7zpFj0id3YkNMKG1rRmr6+BgmZMzQS+dspYZMThG2uemHO9zKoOr9z7mSpCepgW/
po/1oe7gOBMhuERqtTDyXmWzHXleZE/vN8uMdfbvZ/BwpwPARHkkiQzovyRLSpEN
BZBuJlq9tO1A93uNcCZ26in1PfF3Bayq5R12MzbaV/YeqVZeJF8Ldfrw4qcma/qt
4GLpiL+HaX9dOLczgtbgJOF91iQIDpYeS7RIKyAiN6RqRnhqTSHt9pxe7b4ClYyf
Kw00S4DrKLX5rSurupgn/92sVpjtdRdEGHqog+7zEZDYCD0FQMzDvTs+T4QMCphN
R3CjPwYALLU9dOR8fIvtDo0sy/IdlsxVqfXLYm6mGfkTYf67W2nCgvYPcPbEUdBA
1NvR1fR/VG9qJNI173cPAAyfpnJEzvO3IlBvfJKawQcGNWAkeO3zLnVR2OeyPMGh
exKBI8aqwucDMcykGUjNwlkPY4BrVpRnoaUe4RasxWpb+ClIBy1kA1Od2zTCuAaF
eneUhKVdjCCLg2HbP1zVGnKdW3j4EN2iYOzzBBVFXKDhlavhk8rRMcX7WHThRTxC
klFcguyh0W88dNtfDb6mKye2fDBRqvoH9xX7qxFDMLKLTNHTBvqLGtTfFY4B2/gB
O97PUzr0LzehqY9LHmKHpDH0bjL4sOtauFkVtF7VRhxXQDiMqjCMUd94fNpsi0dQ
e3u3W6GPJrJ7R7zYwXRC2L3em3PXd96+C/L8IudCr3gmbXETzjMfqZRydwWlLv97
+PA7cdqLnqywcRUKjYH8E2JTetVsI7xQoyIOUjKycBKFjhoZG0454lZBkGsF2faQ
9RpIjOEW4lKDqZqrMltVFfBkV0kqgl0V/ZIYHQa5UhqMETUNZGiwQNhNWlpkfzV3
O5r2jul6f6sEWgYbaW4EsqSBZO7XIAM8v72uIAxOUQxcO+PnnHNbyV97Jnfc4UCJ
uSE8uD5BgDKdX7rnwKl+nKcXlC+Rw6zvtz7Nwr22EYuskj7o9j5tLA8XV+73kpQC
VwalrOcyqhVaT8NpLLmUdcNh5IsSlwyZoWeQxMPAihBHkwDNrCt0ONbh00zAFga0
nnkIwR7HUHGWAY+NNGko29ikrQpuidrkhgHmQxnTBKEDHdLSAMEFpz/kZfEYNfS3
rVcGECyHHn9aBMd7nXtmMdm24o9E7HgO3ZJDhWZfn9NGLjKNkEA5qxXb/dFP/O7k
Wo/0b7HXH01bNf0Kdzdud0fUvPIt3d9jov9l23KzwletBeLmfkk8iwmJbO56XEeK
FvTRByOrVX4sZTA0XQyY3rOpGXLjDV/HVz2hmhoJhQvn50L8jNaRCZYFLv+emmJ8
qAkBdCyEKcoXnQwpvi185KkJrV86clb5aVC5V0NugUCPG+EJpvzcrzPnYPYQJyEi
YbLdb6My3Rhfn5KEpJ7YG4kKp2Qot904BzX7/P2wF7ByNCm7li8l5Jqf2r6aoT8p
tkWIxm0d9SpJbt5Au00jZoW66lmfI+fDt3pBjpzdO/9lQ5plZYykFzi1fLwWSYTf
3HqiZa4BV0rwNaKGQQVlCTO4ImbrQuB2oZSqvKUgtqC5w+Srs8s7OMeexSGOnQp+
UXhdzRKtcXc4xqeNT97wOeCVNqo9tLsrMoC3IermUDZTrw/kZgbNUIIHHgoLu8af
esCzU7TlMCgHLD9+AV3WoLZ0gLjXq7QNnGaaxyU7iwRksphr15sySarUpvbnJLsF
hcPficsEx5ROpi7mEzncU+VDit4R3jNdS/pvDQzXIrJOX30ao4Sf57cv609TDoNe
nOHxI4KAqSCX1nakfvMhm7rhbM6Ia1TMLpbGJ30Y7+wPIkvU418omxstaxAg5cJ6
sI1RASSh0e/qUz+egk1UAWsWKa0vxvNHQq5nN3yygt7OOJ3IFKQWl9G1JUE1ug9J
NXyCcSraOdEch2PV4FRmie2Lxw6auKPW+5vkXAQlyM8xAYaciD6XnkHuGTvi3ZFm
XrnBvcyoqHBqgPT238sDaMagqPT4FKbTf+nSsh42uD8mrO/mOtBWdNbItZ3wDYsj
6guT+C4NF0oSvc1P2G3xZ8FAxzP7/VrLFkpIH4GpX6FlFXp7d4nuR2btzNqJ+8tl
CKLyM2+U0SAFHYpxBTmPO2V++RQM7s0Ub3u/pckIjBQ9UQdPAIJIzt6Vrj7tfH2U
KZfFsFwEgNmnawR3x3ZIaD/AKlwro+YOtQOwKocSDevW225zop4lVsurG8C0Pj3T
dR7WuwSbx3e5gXk8Umtxdx19mYsCwHIv5y/9n9CqU7/KTp6LP791TaCWUkK8/yS3
dUcO71UsmuzA/De+qt6zzfB5oBL26zRKzMahAf/zvOpDnPMpbbQj1MZLX3mkcbls
4GRnABlmtCowZywgKQomTOuBkOItRyntwOcP2bIoKlQKXrtIXvnJnwsdiYsbCem6
rdCGa1eYhOIcw4LDADy8LdHCea3x9Xzb+D5KJ3QVK6VqvwTFdPdV7XD526pQXhhh
GqlAWagHgLsyIt/SNmhvG1YhQnEXTczjXmULSvV1wu1D/7mT8ePbeYp6L7kb52kW
eUOKVcIwNXZcxn3jyCeyaGfyRfvq8LMJ9nL7RCXCImEoEVLdKQapHgAJKWifBE87
Wtbvhk2y1e0uLH+MV8gurnNhJXQTAq1oO7CJuDF74T8S4rJaGXGGjwIwCRVIrakC
oARQB4Y8xsEMFm0W4WzWj/HePCJq6Vh3gAG/4RMg/CvUxIzzKuVr14xhctkYujug
XzG2UVR2cU8jvTI71DgTTH1aJEX38QP3TSE85Gn8UsiTKyY1Xyb2obD0F9vPho/+
kttiPnEFqF6z0B1OBoKpBcpQqXzNmREamfaGf2iNxs5iW0YpaXViZPIWm71tZ02A
clr0ZA/1I+noCJdNJRR8WdJGHWnrIszmC8QC3wyE1UmXx74pLd4QE5o+d7hWpHLY
QL+RC56QQp8JHIdcO2+d4OP0o7wNKqm2vOuDJ6LpL4OVv8O5zBbrsugkI5+S/SLL
Tf232ACzCk5ixCfjkOAZAlJxMm7PUSQJ4djPnlC7Bn7Ekn2zc3MJtS/DSve9y763
YHlY+NHNrsF4adLFU91CvrCyhbDeZNiWW8+tEjNIPOx8jOGlnBrrAOZk6VviFwMa
zQ72nekP9VkU6HWqgQJwpKrpUt122csqps3iXZFvWqVaWqpNlocF7Goqdv7RhAtU
0hdlof8Chh83MWMr5qK8Vk4GZcvXu/bcd5Ot5sjAmEot3h7P91S9sm4xoyacseDX
p58DQdObNyoU6d6pOH6DJPWI/HeTGnQn00u000LBRY6sySpDlP0EyOfBzYeBWOLG
cM6udhDb5Bb9b14AA5QE5Ao4+uqMng/FZlwAbHXkr7Af8mDMLBSsA1XWS+iTKzEO
3KsBgeocMM+l8o7hoMWJ6WkNtw0UBBRLOKujxq21aOCmIIQR2xyiVOoC1eRvJmkv
pzKdk66cTqeLWVnjb6qXizttlakHGk12RrO7u8WBg0UOtZFUo5CxAq2yV/+NnRQW
YWeYCN8m7jTzafgyqeKOgBBL8oyY5WroZmp1u1eaqcUxE/T2V1sKWjaoP91MX619
d3LUzMxhcl/mHDKp1S2fUFsoEnWu/pPctfmKZQK0SXObZnVil94DLNqPrYd11wwE
jdMqaCe7gS2lHmR8oMSiZBZcMk9ZU76jGgdaqUnJuG74bou94oZo2WrmPNBD7V3Z
CTg/QKSLN9nyf/KSjtNeLofO6TheStp+mgnBD2Li53CFL/Iw3wQtWInIh/soxldw
hlQfnhVIZvXmdUt1XiMXBITdg8vCI8xx2Y05OHHY3cFDHkhWKWEQJ99ucY5+oQB2
/j/sfLXLgDkrPtEj+lWA8fp80ftWo9FiPDK473NzGE3+Irb/SdBuC9rnyFs9Cidr
LjPdDAhR7gfot0WOIX+8az8AojlP2sYnNdyT5O9QSoOK7DDioBRiHxLA1JhA1A4K
DkW/pFRx70C/MJ4byngxBIfCRCkKCU+pIeEo7Kr8/w4bpaJXu8WwZO2hnxQjG5X5
JSoTTW4DqMdwNWtKRqWcLwwTRN0b42/u3KMYco3uta1uPMWK5Ovve0IIeF4tA8b9
HH1fWpANqxsaA0D+jDOcvRg7h3qS5ib6xNbRzl7irlY4//Yfa6PP5swnQ01rfraz
+DtXHFvyP0lZjD+j9pl7nD/NbDsy1jQ8kKbTwatVXUGiW/EbJAj7ntrLex4nzFHi
Jzybb1+2+e6sg0mNe/v4Rg48x76+mVQcfbhJ0Pkvc8amKQvhbrU82089OjynUPi7
V5N054+K9e+iYFiGYZPJgFFaidPblJA0cGfiyA6j3ySAEIbPPdm9t695l79bMUnT
xRb3Ia1qHrnVFyzP20x53DVJkS2VCUOYQ6jsdQfxrQ1GV6/d0yA/9qKhAM/sQeWC
rb2dBV1iVLw0cW+veo517dsMhDMLegQcBcaSPVEQJ7vYXMMpoHya8mcCkJ9smtdQ
y0Jm3YDEDfzSGhmoxXsUZqtgdp0mVkAFxwE3S6T91C8z+GjDrn/rGGEXcLyjCHBr
hOzMlkVyoLOzq2ZVjEpfHBQGvoNi1w001+WnrwN9U6VBAaR0nANpo+hxX2nrZ1Cb
h7vXYYG2T8OTYkUkdF8SQgWudqAlhS2RXdKZSb4vwPC50LeVUaH7CaJCZzVv7dxS
gH06OZzk0tjFWROvxVq//PLXB4ZY2ZwkRfrNX+oZsGppc4m7uQINEZJAv7XxCVKN
K3nM3+2SLbBPwnApSVvKbpsd5fH7ys3/QUw4zzd18Zcwtsj8uS+GXRgitvR9a7Y3
LZsk4UKbpYejrvcdCtAuM0/Q6Cli1Xb7qrQWSknqoL9FAR6T5zR8jZo7ex6vIMpP
rrmNJOSNwBR3xiSxO5WqD7cOK8hoiNzcY2v5YgLfCONI3J2Hl9md1SwTyoqKg1my
pDU3+2eD4uwtCLv/I32fDKjiWjXzr/TSbuB8PxC8a0/TxShSayu40XiLdpo6HF0L
vEFB5yX4uitQQjsGX+neRuFJ2ar4AsYdw5p6z53ff6ymj54b4WmvHa6YCdsWB98K
F8IClp/3LtiRF4A2DcSG8P4mCuuJE90jv8hjqocMZZasvwsQxsR76JnliEYbGeW+
6+uYgwqA87v6rGe3U/re665u1B0haA0kJfK6AskR262qgBb3Bxk4VBCB8s619scF
W9BsvFIBq5LArSoWYeqP13xBxTWx3470c6L7chh+YLSD02e77OeuWv8A2wqZ6OMK
pyNPzvDulpdc/p6YnCjDrzs2/r/sW3c+ov0hvs1/5py0jw9Rix5O4MU5a7NDgL2N
iZbYLsilJKfk9a0vtkeWynpkQ+EYrq90dI/G3vnCt2zDELLr7Hdkj2CPZ0/f3vy8
qoJveuKF9yk6uZ19WAzYj2+6QKZr5fflkt4Fw4GwnTJn1eOE6kTU1cWdD+LzzuOb
58K4ru9pun7puykFLYKeSNhZA+fQix8w3hTvSEPFOWwrvgYc9aw84MHLfRJCusGy
MX1Jbuhz3qJgZ9dJQ61XaEmNb56HwpDCaU/VOYpSVzUy6LeDZbYm+K+NVQbyNjsW
E2BAdwOSlZnLS8nG/XV8t5IjOFZAjK00OElTjXUV3Rp7AdTZux0dk34nrOEqCiR8
VQvQnrgzeJm217wT15sfRcDCna+OIY7syy+wxYe9h/kQKiXh32L4R73tD7Lf/pI9
f2RHTChbqQfaWyq9vpuFj8YCsuuzPMobjgL0gyx0oq/BNhO5eNAHlXufV3vP+B9y
VHgO/BUrMy9+yQl64fBULu03PVOwvfhOaDqjRrV1W6Nh2PTGoW/mCr+fVH48b5Jm
6NK3eBH9DZM0szh8wj8Tefg/T11tZCJTiymu5AN51bTrZe/QSmbO4E1M6+98XNJV
VrsyoHqM0icaEoAEiibN08sRFYlTLV4187lGFSifRccAEaVuz7J9ay9XgREWF5pn
BZFSaPwZk4ZF8dvslWAHI0rUJ3ayrXyCgC36lfTGBlmFy0kyZ9GTgcqUs5f0VlcW
4e6r2EAX5CNMyDZiICHXh/KK0iraDKpH8NTVTTupUEi3pjA1CqiuAKRrfwOaR5TU
SUYLtkicG24Ov/7vqHJds3SrIcCKOY5+VGwRI1gNDOx2WETV49zqSX0CFPQe1F5k
lSt0ZbRf/KYa/e9X2r7UzqHmx3Mx87/82fW1hiJ7ZEgbTGANe1EEjRVn/mjaUYiT
bmWuXDugaUOp8Vgsbz59kcx43zGgya6enq9nS8qfbrRT5CAZRZ71Jsa6GiN/uNZP
WScArgrIIsH4fyf4tH8fiee7JIBzx+W+Ih699a4moKPOEaKdreUwS8HcDwc0SlQE
PzaE6B2XERj75dQlifEHS8pGb2soDIbXwE2mc3NClZW5wzLrHO7yIvQNF5ldsaY8
BRe7hEV/1D6/oyrtoz/mdiuiFqCPB6kB7UE/UmqJuY4cPHvAfnAzIcykn54qovj7
7Svr0N58mvmCTcbCjspWDjnPhZi4HYnr//3B18jz2C9FMePVa9O0j8GwnJMrhYK8
8s37pniJKrchInxW7bAtLMxDOuuX/5GBtlLtiiYOxh8NsI0DDJ+LYcvB2ddL6ol2
Oh+YVbunxWf6TGfDM9cMJHTDJVUThauCF/GanXc/PaaPQSAImyvk2isn827YjgK4
gd77qveXlViJwOKSejzjiX1vNXRZn7/W16pcdBko4AtH3JOLP1AQXWqprSOr0qwg
Smn5EnwvYTGPV4m77Favdgzu2R5Nd9mEh/f3E8d9k81jH8+sRLX1OO74yTUJ+xlw
J/tWOW5hIh7DnkZoc0Pyb1ebdPRTvinxXB80XEHofEj36n1MYuKTh5wv8fRO9lWW
CLigAtSW+CjOeKQ7czP8tX1ZmaPacifhscMGIgDwfSQ6URl5dn77VZUkj+nVo54V
TCbfha6G2ipyqZ1y9EWEkgbjoBxWXnv6AJqvUV9DORSNDOWl2DDGvahEkvaNQsoY
/Ra+Y8GpYnHo0LwESP0jeetCN7Q9k15eDStx0OjLWlTaQRKMEiFfk82Csp0Vxz24
w7HeJkNh33bi1HXWrOYHX1ZViva2mLpY48GPEc7mJ2KlfHUN67NY6mjpJtDjEgJu
dtwa4AcGbxVxU2vcCuxswZoOq24AvTfXE1wOdef4O0WwZJmFL4NSSmchxswXXQKT
bJ7/iE4US+U3wndPqSHVKWnNlJxtYjVQP9bIvAoBnm1CTSByqmrIdDKXgb2Lne2N
ahylWROVxVhT1z+1FlEcUGysecZEZw1reUmJPpxFwemRlgBC+65Y41lHerbyh4hL
GBWsQlBsQnACBRH3I5xsfPROKyK6CK7ksedXp4MDgxB/MAD1LSpabdKVk+bESzGU
vh1i90oaeoWTZtcQK0JfkzedC93n3+R5/CDlwQgECWS/wMfj9d+WSUEaJFnpKNka
MUay0pmE8/VpPvS/+9CfjfX/Rdsx/ktPCyRcYKB6KxuM0+cgKDOdvmAM1zHvgsui
O9K0n7miNVeDZXqS3uWhuB3yctPWva8HN0/y1l26HgPxM8jV4kqvXj+1ARN5eT//
OTeJ5xbSCg+ydhB1KhiBEFKdo3K/f4qp5pJViAB5XpA2Fe2j4zfvV41x5M8Jv1DQ
qx4hAhBM6UD+quts2DVIwjpUVWuKPNTMNNzdGRZr7jitSVdyJEW2BxVFgEZFupR/
VtCQaZw+2e5QQCwxZLu60rFVnW5cOQnz+nXpqzy9LAb7f7TzOF0tHHGCHsatxgoa
1vXpFP+nZM1Lnov3gLaHgbrNWPzApmD1I3Q1hCAX4El51IxCQbRVi5CS3sVMmjB7
pvBZvSUygUr3aJx/Ab2ClS9t59HArmWOd4fVQ8rGdNsl223gfjo/etFoonyidmaD
zj+FiJr3hL0nmZO/m37u/Xyp0uq4G2wY4MQg24TlmGiv8dPDjiE48bjOkuBKJ3kR
5+4B67QX4WhNaQT3SOLR+Z+en6gk0df1SBKyAU31Ilzv2mdMNiDsKd0zJG75lWWq
w4VX5luvMh7K9hRrgo11Ft46r3mlI52QnJYG1qVmsVDejd9+5em+r5WHd6Whcy7c
HLKc6fmV2b/0mV0qmTPKY/fyGbQxYN+OKlzeRMO/HKnfB9VKeX932Ebmi7EQCDv5
scMHgbmL2cEDb6vqbxpQVcNDQA75Lav2Tfo5pJcYIHAvHdiSDsq93UMrcK9HTqpW
ZSSHL+Oxvv1y0GaDoZld3laJK3JYqVryVLJcWURAmh9vc2mYOdJBdK5+Ut8XQ0/F
4Z7iu86vfxDhoJQxzQ/r1qq+HFnDZtaRpQ35udnAVHek+OYPbQ6n2M1OoUNjjCPY
6bBmih8qWiTjgzmyL0hn36YoDE7zwkf6prbeRG6NqvFiauB/YeNUbuU0pXJPwr0W
D7lX+mqlaC+llX+P01XZoa6HZGMRAJR/mzGWNh1k8xRC2SdglDFWIR+QYlTe7hCo
R4cOPhhLd2ZJa/x4+uL9PJOyXRfSA42R/NvYOTK4UPCv7kTbXOHANLxFywDnKzlU
9nLzxTDduFsqLEOLAa6kMKbj0TjCzdbvi3NWO2HOjWSGEKNZkJgCED9Mq1Q1FkA9
lk4Y5Qt/xyx4VVWiaA1AzoF+YlVBB/vTDzOdz/Xa+3r8Q3ytB0cVN7AHv+aiBPwB
2W75rgtwdRJTfDFTWPhjJnGKBv5bjHWE2ABKZIuh0Va60So0+PgcoFZ177YRdEcj
2ZK0mB50qc4Y1TbvINZt06Q5xH+n0ofrFkpD1rUbLi9kVy1etFeLg22h3MPRK6lD
nylF87Y7Fye5xIUWt465vVv5TWQHohPtIpM2aLtzfAz1GSGwj194DxlZWg0/PiZ9
bsff6ij+mNgHr3Hm0BMcsbsw6mRvMwitjYN/aPNBg+NFKlh8wYWj2W1Txnp71+px
CdIcRJNjxE0UPav844EbsGkjy7lB5StFwQXF/xeCpqL8/n9LU3aakz2yiCQdrSb7
mNABujbS8BGrBECrfmKGbfWW52J9gJ2cgCvMFyrNjRJpi4liNX50DRzbMNC+JGrB
HAfBf8+iygSyThX2HWGv71/L6uQnKsQBQvakwYZcanrQsbVFrSJUeO9+jQcQxsdI
+ePPyQEO38sODWgyCzUH8qFXpzcZY+oMz579JhG8MsZO72l4eLf93WkkVTUrWQdp
JIVT+7P/h9dOfgZTu+3aaZ4Gw3FmoqbTxj/tnWB1X2hBQtLJR47GsrzgLPZV0WIm
U+SvQmnwDTlMNRcGr3/TmotspTMlRYeDjV3r6j3vC0p+6ZDGiphiqzV1LwiRq8u7
cMQKwS5NZ+FFaPKNd4T6XKHpgLe7jzCGXK0ybJMTQJgvD58hBeIM8hA43AKT5/FF
2WJPi5PDfYnN+eDgZeynLchCtPMk5AHxFg06gzOwGQInqcLPNk/ezua86zYWuI5L
XSH5VVnMKULbIwgd0bzw7OzHGbwY6HHzVhRbDvGCkq8y9PZjzOGfL/m76x3oPCFu
QdzX2TMYXrgpSFPtgu3aeps4xv6s8qVYMiuRHdGX51V++8lojwy7axP4A3amve4n
QhWKkQtEDzL9b+06h6Yk42i1MpKjDxrHkgkoy+cE6nnqca7B9hsuvKHnvNxoHUA9
wOOTpw+EEja/jN1fuIykpCxOR+NU2dtEihvyjPvCgHtquoE5OxWyLVoRPvhKTIJi
FVuw+CNgHevwsuYERXvuYSzQfkn1xEhJsheDYE/XNxyNc8s9ntW2BjkFk3yt0mmt
necOjpAuqmiG+ArDahbVOqwquNB3DCcZikbPB5UgJrSt2lcu5XwEiHMwqkD8b4vz
m6kqtwQqWDWtdU9CKkAtGJPibuny/o2Fr+Yv9POhfnWwtOp2UBCmldt70vg8fLQ0
jsUIpDX7Bl/cmY9Q1qZG6iEVo5SXSoGW+Ud6jVunjfsgMa6S8dc+CugynaE58XMN
M+qIQto/cmnHkXLm7CBodmNpkG8qawTUfVFxBw+ASiQN+3AIx+FxcwyhrYvJgKSj
n2m7rnHc61D6s00W98QQqwOXsJvMiCE8eD2Uzp/KxgROdw8D7Oj6FVU1qg0Umqsy
xwgB1/kW6Ma5RQZm95cLEgTKOkhAb1FjP33gPdZM7R/GDKojG0o+DLfEy0uuEvH5
QpTO9D74JW9qyqTZXfnzlk4NPzBiL0/3mU+5bQ53GAw9DTReqdq+K1IVTqKPviSH
mI/7NBSO9nrxKx39BUWqtfXtiFB29SJntuFKUJ7faGyLgMM4oUDtvFS2BVcmbjp1
729kWemocDnvoEqLEdAiM58jVdSP1LnUh1HL2tKSuKGqgitDZE6mlG2JbArOebjH
vA19zCbfBTZHHWLy9Fe6Q7YLtPlnRQ8I9iRmkz07kgVnHXSn8rDcR169qbqM6GL1
c7ikAwok1XR2Hl4ddP7/m34GGBS7s2M3vSW4x1qjHwSnOPsPBNLOZ/rc8pWongZg
KHt9hc6CNlyHRbAcZotjV8lJ/UPpUAMbxFuOfFT7Jx5lLav1G+So8gsafbctzJ4A
v0whNLk1JIMkjt/KTzkjyUpISXkVITRPlXB6ipNwB1Y/1hLMgvIJL5zjj0pkTIfI
MUfl5WKHD2dWjkT2wFoWIp8XgFmLzSVDalj1bJKADSnot88bfJmV2+wluzJvoJ1c
HyTHThlwhEvmtz0kGh63Pl8dZwaNfU//XmWiKRwNdYdyzn/YSy34QJJzVNzT6iuF
ZKaMkJ6xuAr2kWvDThDFdLVdzgzW/ttc70PsSymt9kRctVebQYDmzA2yLbClylU9
F/cVJH3+YaYa1DEa94DxSrIipw7khTVHSIpFFwLP1NZmDM58iGg7ByXt6i25/uet
CCh8JDYqN5P36/+tRv9V7JD5I2L+w/aQHpJj9RMLzbztvBV5dBeEdEZErlIsFNrx
Yndl1BkhdqcXYHKZRN9dVtCjQgj7/7FHQmDumE2amFfiAMWgcHNJLxLb4EvnYB0k
w4DLj2iQ7hR1ecrk5nFEr4Whe/Job+c324MRkbl0egdPiNwfSHr5hx6/lN2oxHIZ
G46hAx/EeZYWg1NC9AoqwdmzcYhS6vWeKdUYmdUp0jkD1ogr2J7SNzLvdMB8K5zj
7j9Si1MWNIh49N1ffl0h2ByF/22E/3HEDfcdkibHbplyi+qogSUgrH/vEGuUNsdc
Tzbcy3U3CdHymTdpzLaZZXOa+tCEi7nP6VomR2ZVJjmMfSrlVlq3BekFdW7/LOBB
SyLNAVGCRyp+XWGc8Hc68LnBBMyfDIOX/tW9aCiWtkjTj4xFCrUQSacJ0so/V3/D
1KSat3F44H1rRs5ajJUNt7SVRpgeanTru9bCj/bwjiJFJaEyWP8qkXwb7OQ80M1N
llL4PCNotv25ZFnBWnxx2tmraD6haNVXUZHrF+ev0j7e9OTIcaBC8gTjZCwykPO5
5iWexIw5l2cO8wDneSKdsQ1V9kXxkp6TqYodr0j8N+vjtxWs4j9mMjinWaxT6zae
PrvHrqDKoTvtzU+lRuPcKN4D9+6xLdKJJVCb622k19ro5UMmLgIYGfAJrjvWsFGR
R8wh8CXapqq0YYHAUlwVUd4QAy6jPj7ga8l7tPNBuBTTPHYAx72mvioelYJGAQtP
vM7pw83L2LHCbVrpCXYrSKNvtixBdICggg2l73pbuMEW+mxuEba7Ma3IteYMA2e2
yxw+7jot7uGlqQApCScV5OHKduIpNqSjyiPyVIbc59NP8NTiunikMf0A1JY2UIuJ
7BwTkloeRQpb+OWplM26U6lFY1Xb1EcgcTqOlCIPIl6yY1EHVvi4wnHLXg+V+RAM
Fx0WG7nFA2G8rnvtvqcB/ThwPvnjYACNuwjRZBVb8yrkGuERXZ0CKtOH9eJLj6kT
V8GXnxP5WMxp4Msp/rp1j4S3fHGNMsUWBjYFkFYAMsjUQ/LGvWH2brDpjyjV4ARB
lO9fsXYoij7ZFP47sQgstYL++y7p1XOZjKqeCSHv7c97FYF1hn3nLw3XNOCZ4W46
AgRdjQ9qNDbpphS8X8tRKisKtctyXTixnzu/v2nARWVJMrRLIYM7W81m1seh6b7q
88e2e+sHZlov8EHZBGU2qWFwy1OjDwp9GJtaMiy0ann5YnCoAvzPZTLS/aruq7va
cDubdkRxiIj6Is4cIAKTLfCJGRKDMR+Jov7c0p0jMBJEAtUeKzC/NK8Ke8T+hpAQ
5BXC8kIuaTxakmItMM3NWJBwQBncxRJn47L0TFuc1EwbPhmQYGDRy0F1MwKh79aO
lPacjISUNQRAwq/F/CtB/zNdDS3xTJ1dYqRUyIgJNCAyZ/I+kQ1PBabwx7Fzd8WA
hAmLNVWMNFSX+082c3Ze1egAnreYzifT9Rdy7njDe8etbWE5fBTXzo1Pg6jOuDZe
xvD4OlD8hvXKIyi9ziaBzIX6yW+cm186jKayNXl1DpNNIWshc16xBM6jl4yY1vgk
5atBzF7HSjlbJpUtCEOQpXnvNNaOx1K/eCA7zjYDxAlmO9aJqFxotsppAGMsPRke
D39DQAowyjuSe0ryIGaIWMMJo2BJcv2/1l/Nt1GJPZ23e8Lwpcr88g5OdOhzZ674
HYbqx+ZeIlttIjZDsh4icW1MxhY34u1ODUTwfNYABUJE9h6ogLAwuffYxBq8WAdO
HogRQ5ZN7SwOcXm1IS7kbhGLbMjSg/WNfqNk4FleY2AsjmmTVnwAeoJRvyOduWbY
60DTu2DyxNCNnVnG5dUqlDcpy2rGaxifxn+GrcLQILzaWzXDKpdAgoFD8Dpag0RJ
PkFGMNkZV1zQdxZflvTsI2voFp/Tk0kzbIuhbn+VhexMWSZ9bYUyICGnKKJosf5y
fZC6JwgnfqVf1y3clJ+U7x3jPL79CzFPg+5gJsjZUYvdt79lV1qLjjBkoYGjyPbb
VJ5tMvRtsZKo3Z54QghfWhQENvDO5VIFtCnehMBCO/gvoVgXnETre4nQSgK8gAN6
Yn+b7pOilHRWNvmE5wbYAiay2xWU9mGP2Sfb6jAvHPltGZ2YlW4izpdgL1e142ht
j/a6yAaQgiqsu6MbCa38KFBllfPf/rAzY8UlOAEgn6YavReu5gJ0b/ZMRDS5hKnK
Tjb1K1i3/uigAhg/B3GrcKoROWCrybjjmLdWt34G7m3MZMdHlq5PXEFyWhPM0885
MI8o/Nv2zKKRdYoO2XqSGSETbB0ZEW5Z98sb4KHC+aFEJBMOACqVktdWHvb5a+zp
g1D2yBZT5izRvzw897/jVlY9gsVmZt0Qqct6Qyfsi3PsR6NJnMCOIPv8qxf9rjS0
6vqovW2Q2iFS0+wIFF9QUqCOjYNCdrtTSK7lvZMr33PNdez+yONpI0ksRKpJuqBZ
2wq2++pTXkXgOTbSclRVJk4PdICKS5e5DixTX919yi3KXAwNGPcKr949pXn+WUjy
qgTmP2k5OvkJ8aCvHZ6hplLNDGmnhuyq2tYPoeoqEv+16h+Oo7hQdPC77/+GWeTw
9tC2q75fzxTOo81CPkU9ZG1JuXbzQOBS4rCznhmMJDDN0I6w2ed8abo41MZ+PoJh
CD437TTELXzOnpixgS6qlLVbn0JKvXyi5mzdBeBjH02gQ4MO8/wx94/O3zLTNY6e
QLqBq/pn6zhKxJelx2y9jubj8xXzfD2BGne9dLffWqIOMZz8OlQYWD1xTCCQGuhf
dziSmGAOQ4oE9gNpnYpiOZxF7tZNP0E0waQSvLq9efQTZwFTqm49id/qG/eRcls1
JWBEMBCX59uKXv8znOrp/GCGORNipHhKjLP+Jc5BY7g3M8t3/5SG83DhWUu+pnYG
mNEOTAUv5FG/IXIYGwvNWHXbqytfWciH90PjvnnzCNLrDmRqiBWqSWyXp1tyLIbX
ZQhzEFUOUcJk2n57Zs/ie8vsYM4YDazRCLSnppXTQ6jyNjYD2H0hxM5KFZJNur9H
4291xgMsH1T4pO3Jsx0cD69cVCd0ZkDyiKitLH15UXvwiyMObBNzoyQlYtHkCHit
xG0dbbFknRru/K8PcHhpydOh8HLL4KIv5P1EY0PTW2cdPTLSZqPo9JWYUl4hK38m
XUBhnu8TnleO4Tclyc6TpXti+uBUjdZwPAa9zK+6VdyW9vm5aD8KODXnhEGiJ6fB
CA/awWJqnX2SCkWYLS+Yil3wJMFzYZKCH1j1NkaqvniijK0VBeOSt68FlMpTGsGc
t4QYA4gipLbWIWk4EpWgPVgXE3STqT45+S5l8IhkrjvCz+M59cMeI3pQmAm3yX03
8gTmLkA8yfv5rnTFXv0rCc/2IStObgGkGc6+C2lI/vsn8PVEsuplq7cg49hwipZ5
rw0eZZC6oKIrxfauq0c1PDIKEeNeJuZvKkzwNjLix5Uh88Rdkih9XQBn2ghg9mEY
R+827EQ0U2Fg6mMNYIKBwZcaLMuhRcb4XDGViP/kRc+kLWfMTmep+xxQmhBQXulu
LDqnt+vqwSdBwHRWkrx+7PZkh6DzsPBB3WmyzXwjSmzyMIuBu8zzeSXzYR67nyWS
k3id5ECLNGt6RfmoZpp/IyrUobAT/GgRnn0L1WuTAKjHNwez3Di8v3BzxLZ3ffNL
hbMgochMa7vgziSHLzi2NrvJL4iz9D+WDyI3HxwkoesavnKbdEJ+41/coCLd7WUF
hC0Uc8OP7yE0scqZIw1/AXViluXR25KAk7oC7NWdgmTP/Myj6xKum1u3nO8kbMxl
5PtieNbQnmz25jfQ7kLTfP/R858khzJSH9PVZcyyBTN6lPuhSOaHMQO0sOIQi1Zr
X0gGlwrTrxfu5jktYiFtY7VH7FKcabsgDViDD8msRFWvXi3+bDm7VR7fX7eXHa8s
+TQqtxkXezfyFRVhTa9j++b4MTdX17yriaThy5rX5xYh7FnGhFvQ6JuqEd5AQ4U0
P6xfXs9IMv5bu/8kq6FOyDzpiIUjH8LCeuH7mhGXVtRVG0N1LaT0annB+wQ3xuYu
9YESGXS4Ct7wf62I/9XPN7zwL1BFANjDxoWhjM+KoEAnp+o74TZxWszUH0d9MGSR
v/aADxLvGjW1OF9zVf8SN2QoAJfFJ5S6YkA7uVAg3MQO4Di03e/MsJnaSsGnQ2ft
VEBxZC8/096KmUj5Yu19htYJg7d6q757EELAcm7cqkVx975rMU7Basm+TAEvL2TA
FYm12mL0wZueKSLCZs8mwQBSt84gUZa1qF802uz/1fVpCQsjM7w7+1nAn0lVUx8a
cPptXCH0ptJld63mU/1UxPGfUMmXFESiJXhd8lAUY85Ay9PeT0b5VyxBOR5r7PPx
Ue6/DLnq5rK4i4h8VDlEQvuruMJbmLVH1HiERwg3bHswtxzQJcz3UPOV1Wzae+vh
oDJic443r+i+RUWzbYEUqVq/cVks85r0V6rttyvudIkj9fNot2Zw38spOWvbBma5
1ru8X88cN0ib10o1fu7BMqhdsMuDzY6+zq0tsdJk61HD1RLAfvGCYeCYhCImw/5P
QIE8d7Z3GHQGKBq57xSKGoJKr5TuThToyi343e9Bb1NY9D2dpz1f9/5SqOoCgf/A
UYbc9dh+9rv2I4mEqltvy5e4mBhX2kUXwVk+WRtmwWPLUpCNYJYVQa1Y3s40jaCX
OcjalupancFWcrDsWmYv5iSXc5tyYpMA4UA7+reu6Cmshneel4FJfcVDpR8wdo4U
SlQ6DBZWE70ssWBU/gZw4vziR2WCATQ7dLhh1AtLicBRsOsXNL9E0Eg0cz52QX0u
JtYQPKOAQWu6sCSZnLW41ke64Nsjq+DQkJ+VqX9RgXbYnjci7X6tvK5oEedtveno
UIlyyswciDRCUHMNVMXYcfsLtJ6m8nRhCBgHY6OTIvJgAyW1GKhP5h4nrjwKeBAv
MCYtCytF7yKNl94DsCDlO2WpxtZipNJHMpr/3iszJ8aDkLNlOHmZMqh64OECfvp4
Mb9Nq5TLnm+An4OJx9x2ytmo6Y+rQjZkRMWYOJ0Uf0b9jgUvq+WcevnR0y7D/F1m
u1KZAkmzGyM++VXHBsuPXFShuaLfXLbuJ69E7xL6mRULBkj8woffF4W6+zzuzSrf
XBTzLCmgtz5c6Lxpet17kmvVCzFm9RoRRNAoj9/ceRqgbB6biXpA1Ip2PZh7CZLL
qkL/VGpdh+A/cfngL/cGqfGmjJ+L01iTOGGfqR3ZmzoSlICfeXkzJyYIUcaN8/b5
ncM3v/lnONXnPHKcbii6KehzIsORCt2ampJWTdPTasWEJ/3xL4rO2+2e/MCovsnr
oyaKwWAOxPiYeQzQLFPy3MKrbpqmmxbnGH3yB/XxZf8rzTZ26C5lCtnAFZGu879u
fMEEP1ATAM+TgWenB+6kfl0NOibEECFQ1HL9k5tw5ncAzRdEbhoiluMFpjKPOEaT
sScHAVOkWFAsu0Ubxf3q2o6vify8+tIZyDCGAuQDybFplFndoXV4qmA98M8SWsJd
o/H3ntDszXp0j+K9Ii2ereox43W7ixm8oyQb2qpFYT8zpnm8mRAI4RbrqJhrfeZ/
7VJm27fIjwonJL/J/0MjKVjgsjYbup9RiKbcConJq0rsQ3NR2dmEjx6rviOxNLlO
dDJY2zqx5Go5q5ks8sYQ/8PKyNAWUCB1rojQOMiEzbYbQoBwW6AX0FJ5LNgLwg1q
SF3bkJlNOeDsFSYhz3Kbl8buj686QdjNBVNfy2YVrLd3htUlvqY4kEXH57ezbffB
ew7zH2BdGY77hCZwijA/SnHtj/Em9IHymNpBoZSJ0Y+WTIDnUu6bYkUqEY2aBFUb
pJbjWQ6GMrXqE3143uWDUAX1K8JJX1x6cArzM32U48zn5z+5kbVz4JEVBrnjlG4f
l3DkD3GAyT6L0jr2Duk5ez9bBYiYHwCNWuOffFfuuJBKNMVVYABnnwO2duqEp6La
+VdO3TRo5Zf1aSxBiBYa2tA758Lp9KxKF/wjeqQDSi6VNqFGqwMNJEqTj2kEDVdS
1hKd6MDr8LH1GWivtkNZfAuJ7hok4Wf2Tr4jaK26GQJbHPgQ3dznoBOMNU/R9f9U
2aD6sfjGKgX/ySYqqdClIrtG26zJFLrGa7yZb/O83AsKn7weU8HsLgZQ/b9Qnvos
KUkDTP4pjeFPnC9csAngliFZ/jOExMSmxI5EsOT9uwjVpfhpY1reenZO4koZhFXU
sm8kgNDjuD0vdLgzhWsfHjf/U1jj+Ucb/nkjGoihrbEpD1JPhCUqbauBnLWYIFte
Hh8L/fc+eTDBzlXGip93xRFHYQFFWgiWKfj5gOzvTH+t7HN2NU63ijHwkLDv0J1X
I+AMikbfdAfnKXO/t9Jn+ODNxSYSddRhYyuXBL7SN8NfcNMUiqyzEQyTjvmOUCsK
tCzNN0bCOJCbO+J/nBOdLm7fx9yFGXapwxAMXId/nVHFxUHW9mEqCkWP+bw5cF8J
U1Mi5xoQbb5pBYOEn84hrYe/yiparZaAgepDkNtOAr5ZUzPTHoJ+hejcvqcnLvV3
77bAQK66xiX+k+h1u9PAMKAXfqtDIPVmqtXrmkRp5zdVIdfJ2bJe/0jCfdoILr80
jRNrdLR8UJxKvXOxtQ8km3RAh27Z6rK82hPNWy/8zmVY1inSI+W6GttUKVVzICdM
aMj15OyQRSawWYbRv9f3KOWBiiBJGgV6WcQrL36pe7Bo7LjD8oip7Axyk0Lwzpbe
v0Y076qimrML+zQLbA6tdHFEIbLxCUxib57mL6tfgCJiXPiHQxyaQUO5hT34n/tN
2wCiVNdUnrPERm6r+OiAn5cT0AB0+5rqjQ1sZ9oG1UEtuqk8HxI2NyLwJHCbIgtJ
LfNXMBjY9i5Jj1Y+1BjpEr+q7kGQPQACWsrTz5iIxO5z7bPemRWeMvRY4gDtHIVZ
Fj/j7xYujtE9ZPmf0XPD1igzmBMY2/DcXAMfEjxwATWhRoIKvDEWzxIEGqlZ6x1R
WTnkxvM3vnM8MXilXaaXUSJ/334W+A5ldh+z84NulDiz/2JkDzWSkwdqXH5m0x2W
JMInhZA8yWal5RJfsjW+1syUHwHJHFu9LBgGK6tB2XVGrhpjn0SXFKBSaJrbk9ZT
hl4+yS8b5htq/vFUzJqZgzUnYefsbYLUawnbYYhFGQDlEPK0qgWKfnkSmw4gXMH7
y9eOqoB6aZ1Io1644lH65jhTyF4/FIh/AyRMElizgJoxfalVcrWmxwVh/ZF4eRYk
NVZtQYRl6CiA/ijUv/spVCHYzblVxbBhB7E6+jmhVYBJeETftUh5yuFdiKKtPCOU
pUS1UKgcKnssyJz52JDZx2pTOQTItFyfcJhGbd+15q9swIGl1iD7xpMDK1eGiwjM
gFbrugI+xTODXJf6PphFHE7kM2nJE60qTCi1MbB/ErJkedPgbn5tneeRPI+DiUyy
Mt852u5s/B8AfeMTbwIOtZ/c+OJ65OxPCP2NsED89eV3w3Nz+S4EoKM1twZeUtLD
u05bhC2H9tb6f1UhsbBs17tP58vZChOq+ON+JJgGjulbrCA12p8m0tY9pk+HcM3U
JaIYPIO2kUqqCOb2+CFcbnP3OEkhY+cEzdAOWFoVEYj6bA+9T9+rjGEAC2QV819M
g+7qmMyL/sYqP87YfB+lu9FgFgzSK4DKOUrSkBcOush3rm2nPovaQ2Ki+GJK/kC8
SvEbcZKHOZ/R+u6zZgKH60jeWTXIiy1kF3NboMMlxT70+En8aJb5SJCrWZFrk02h
NlzQFpM3eNbOiHzTKy4U1LzcrUSewqhYgXwbW0m3bHAzVBugSrFd0oI4jqoGs6fb
7Vov4YgYjyxUsBRZh52Em6j+a1fpx6xlt3cB+6Vxvri5nD/UcDjCE4X2Z2PKofoU
HNTcYbxkNGRp2Y+DL8Mb6L5JuHcgStJ2uD469qhxcajb9a+3sV144edBOU6QMYJz
PvBf+c/qE8clyhtY0chxQIFo8O+r3xRyYDqPmax5EvgQzwfL1cJipa5pt9olDBws
LJ+ys0e3iEsdf9ZqTkMG+M0HDZSoq4CtpJmu/u6K3jMOnynBngMYzFFeke9eHMqp
AlgLKYd9mtgpfdhGG6N6KXIn3E4j83q6NsEv5zyVvE2Jioit2KUk4QM+2SoTqrgA
+RtRBZ9L8Dha3qH33uvK5ET3I5Uwe8guvdraWraephcaCs5XQWHHbg5JEQkrqDAs
nhIemgzcRGQVJu9XCIXGBdPZgKgQAJ157pipiCmbY0/g2U65Z0d0vYDkzwMynNHM
KBULE3dSAB1qyWXcr44tdXSinFnf5D3F4ge3rrG6pViDhhvxoxmNWJB0ihYmjeGO
1QWzsQSJaXcawztRATgx2s9tJQSgAnyuOqx3N8t31IHoNRPslEjzx/7QfawrUM+k
ajPSIISALShkA7AImXzoX4yVNsVaAtuj7ootyPRduLWFUUlojk1d02aMHylFcgNZ
aw7qflSpaB15Rnfn0E4achiXAg8FaOJ7NN8uwx4Fx2zwCCb+pTFfxWqe0NrrHFF9
NV2ff0xaLWXsYPx2FY57C6nUMBRA+NAhTqLlJ++jeCxW850TB2O19FLXTRAZ4R0/
WoEc7fjhgLTwAXzboVMPE4Y+/5NpqCVSQlrj/s+phwbryJK23YnLL6TFms8I8fUD
fdSldywClBHcA+cmGSCe7gDYFRqhLtEVe0PArbq38O+HSBYEhN7bubrTmxNp7dtx
TKrKatKbJlq/Yg1fu9GB3pOkL2ygdSpponNNFzZD023JMSBkBypPmr8Z9uBfwX/3
myUf0/hdNH6mYbbo4+Ao1HWjaiV+pwgaN8gT5w7TTUZ/D4ulZLrtUdYiZPYoXLq8
gRn224MgE5ERNTf7VF11eTXl6ayrtrYRNmwkdHcfoR7RJfHOyl4esw73Mar2/feT
MbGAkhez6q/mE4/w45v/77Hd3dY5D6/nGzt/OgF4eS73q4O41DQI3Oj95SK/1yRz
JQDlUQLw9WsJk320ZERrW0FqxxsKXxEqj/3n2YmlSKHbn1Iqlv4ot7ueU7SYqVDj
E3LNSOrePNpAAavsWJOGBpWDPuuGbw+R55586nzLO0allCpumomcaNVpWPCTrDoz
HkojLx7eH/8b1la3n/6gBfV9T4MD1xXNY8VOPGhjPskt5Mx4moVAkeWn6y20zPTS
VSfEFEy7ZdmkNNhvMPcrw1A3smDyqAVzgMXj3k7VspPXBg9ogwloA+XCoi/w3Rh5
biWn+D4fNpkjjEfOfls6UdrrPHqUwQ/cfxu6WrkxGiR6Qzmva96lAKn5/yPH+kb4
kcDDLzYK7iNJieWC7V0czLK7J5kD+qVMO0iXM4h6nmFo15aQgIfHXWsUpZmTDdop
XUi0DSpCPoM0XQ4evSVcwY0sGAVOK+kR2lWgEGeLui7oLtALvyrlQ+AHQwSQp0yW
SZNlCV1VdbRE67OJprt2+RWXGyzXRXemnPnolOTBwzE9hHmA9n44g1Gkp+3539rA
quV15qggN4+CekxhDlhTOqsPErcdG0wqwLvq1+OJOVot7WKM3DPk6wQLIWvKk+J3
MDwvc2h79R4ia2lFNeC+Ac1gBPIxeQaGw5GhQRj9WUYX0ZVnpLz4KhL0Gw1eFrdT
6DhX3lBuIvq2b+wLsSPMsio4QD5BXylPvc/0oEnUuAU97vdQOoGZkngHUIFejdvL
rBFh6XANN2ZtyRThzySZVjXXOFruWK4j1WHBCoBgmL3h2RvIfctsGer8EtDgrDVY
tQuMrVBqX8529uTMzc6yAPxZsnMpXZ3kwD0vXexKd1swf5GD3dLi9MU4QNEzyqkJ
fRkV/ZBVcOlLzc06G2NOW+1XhlM+8IVobr816BUr5Bnwu4M21anvpU9Hz6smGEU4
F9lcn9cOQnlykW3ckJS62fEPC9EQDKwtkmwYGoQE83ITEJf0WsPB11iwTzWNeTKW
atclDfOpgfUcVktc0pPxJUFIPe+aTq+t9wzuAwOp57xE+8hSQDk0oe1rZJ7YZUgO
Q8goo2ViyXTjCYXVufT+2HJvnICadlbzaIUiQiFOJ9T4loTjjK87vp5jVs7yl7ta
Ifet/lPkbEG2pYeY6BNMGhPXUc0MLPJfRMwBhA9VLGN36sUS/672uZ2jJmKmc61Z
sc83u3TltvAEB6AO8rmoPsKGgWVAg8ChQLiAOJ2G3EbPzZMRWy9W+el6GWj4ZBLz
XqM9NEnQiHwzLJivw7pyUWGORR1BZbrZgv2jTB/aHVqygIploN35OvL5d9yM/qnu
NFd6c7oNhTeetK6FMklIrmwr+T4DfOLem6NboqgTUf1dCZzhgkLKeDU2G7Pmqxoc
hjEPXvCTpzP0jSE+UAUSFyHlnIJZ+T8gvu9iPS+aBdN+/h9aQwqHnWu6H0bmEWPu
+tnQKKUF6Su2VVHXam3RS58ecwDQavczaL+QceMHorz0EunDGaTkR1G9N8GTH46f
LOzfG4XH3KxsFf9VsLD02hD738ZdNTxpilc+pZBD6biRRlAioI89QzHz/MSQiiUn
q1sQ76NQij9sY7dCLhzwWv0Mz8uI3E2O/7l64oiQnTGFz+h6SAekBNk3W9KR+SZx
PPXnjQshn4+f0DHcjuKkOymo7J9TSqzkGoKiyrI+Hrghx6q5VTxF/zGXuiBnDKrd
7cPQveUEL47QoQM4j4pO+q6svRO33hn+Yn4SaVuWEsmViQHZ/J7W3pVEmfvaOX59
dGfP7qPqwQPEqpoKtDB0N3/uISIaRuPolKYl77i198QmeioZrI0OblDDkCl341rn
GOYuOMoZCpkp9KzfAWjOwA2sVRDwdsHT6iMmFdxqRU8P6kpC0W/etAEe7rpNnKhf
On8BNhNqw+yktHnR7+MsoxmAmrLuFTWFxqDWkpHP0qDEQ4cRAU2PXL5oHgdkhsD0
kpvxp/U+xwuRmk4/jMigZYASBKSdJYsaA5oswMQcIYBt1zzMpas1IhE6WVC0BKnO
C0KYOl4QIXkavg2+SpfTFfrOTE18TywqgrtaipA/q0bL6UNNK7KFS3RtYnPOIKr7
kcb+/1+MX6phqqnamDD2rYn5PG3pjMTkj6roFpRzTcdampP2OJaef2Xfpx8PPuXT
73lFmXbpRCMISnIkpisK2uIu+x6OwuizBNGexOq6ADpKR+FYjzb3PbefXHPPQUwJ
NiJ5jtRdd/+YwhyPwFWbbLrMNppWoB81iFFl0LXXoHsZ1sHfM2ycdQGhzkTf128X
ORoYhNsORN47YZ4Rod8HqxoVlGYV20wdkShZgCaKPZ7QDfUjE7g2LlqTF5Cgg13Y
ePIId3QECenyN9Q6icR5SA6pqSvyJU5pBu+/ikRZZ92itrS9TyT+zH2uexROkYh5
fkHf9A8hYNrepmwc5MXdEq+kezv2gzah/Zap/xnyj33tbnIVr63OWt+IWvmxpCsv
sk3TCOF1vBnXM/C0Pb0mJjFmUSgOSkgmDSJCbfqQs7x+KfSuScmnV/L7SgeEzxNJ
kjZe9ClUUczno3ztpGfSFES3J3VmUkr3E2tdVX9QTt7qUFigeG7l6vkh4fqCCvyB
EUf3eC8Tkwe6SyMhe3GFqzaRGiDSEcEGmXltN7cH9vZb0lcbYWbMc/QNQEUKSZ8u
P6ufcmrHwOxHd9lcd3pTiuy44vcDgup+o8NqWNpbJ69s4hxN9Q2236suuuxH9nMX
7/q6wup9neSFqLjeYgTGd+6df2OUERoVkCgBkHl4Cu9nlEGXuw/zhmeVuddxLxny
yxSQ8x6H/4VDQWZ0T1JwASsRhajiGVK1S1QPn7msCQ/Y5QGX1kuMy1A5AuwZK3+0
WfO64LbWvR0OAcS+td54R4Jq58Ijw9xOuP5zgOIGZdAOmWQ5XvoHxkFYr9MkJK9U
BWJNGZQ+c8BzMTeX6xEitud2XupGxyQYbphAIuMFdMdpR2XJEZyg2VSUwRwWvEFm
MwAhhtPBi+8ZBkdJWaRKvDpizssfEKJQ9UhV246bVBbKXDEabGpQ4JVxT5iM3p5A
6AppsB9UkBqt+lLQF7Fcb8VpKIYnFc4p1YXSNaEf+d7H0NSrKm5xy9XYaDjMOfeV
d/VXLAPV3B/7sqUWQo7dgaHK0fh5cYm60liMU3B51iJ+howrfKIOPNilunhjPn/P
Y/gkwyBtxD6PWolM2dvMXBA2AksqPFwnNeSgj/rSBcxavmr/AVcm4lBshn7h+gi+
splBBQ5i3mvt+vZPu+1kDrf2NDAe+dCOFqMPMI4JEW1lelktZw/E7O/c7zuw+QBP
2HlL6zzQx9vdVfS5Hqk4YL94iXkRtdbiN+h3T+z7IoP5BUIzWGbLZGv8Jm5Mg+AH
jws0tWAfV5hQK6CTSwepWiYGvm60RveEdYtN00WkCQh+PMx6C9iDnavq90zs5uV0
pzpYAgj4QnpyL9beTLBu7VVWyK97Zx1mZsob2WivFdACOpTxFCFtj1/WNyZQaMpI
Na7YXwe97GC/KDBx89f89OuFcIrLH8FEt9bd0zMVsW12etNJrP2PEcLGcqaVkiV7
y8So8OUlV1AK83gcXZ1b6dkCCLZB4fUPoIGWh756+gSgJnC9WexU2KGLMD1zgDpm
wutf03Pu2YUZ2Q+36BTKzqjvIByX8iMrxeD50QOi2HkT4U3a48GGpHBGg413jhOd
tuWTxGj0eQb3JKxFv9xZ+kErjqVXRFsAO5/9mlw5OT1X6ixBSrurCENB1yRw+yWL
B1IsHr0iOGe3sM+qEUq9ViWwiRLl6Y/Kc8OT4ydUoBT/omcJA+4nvIS1qclHMeBD
7yNf8V/vVzeWkqa0M9XI9pGwBX21b3JvsMyiR0g8QWBpbN3HKKpMiGsVQNCWtbKh
GFSfUxYzc256KSGr7E/Am7dpcF7PsL4l+3XXLkWAjYMH60OX6aRSfmK9VrMkU0Jc
UArRFVjI8IK8dU3KNxzSCTe4fw2UqUI6ObDoRpLQxBGwnnMBZPJzKdBwL9T2y2LE
6ec9/MtZpZI1i54J6WPLAtM1iYDixJvinT87tKRvk3IPa1shK3lkGpGvTNYg04v1
Le5DoNu7caFO9gIMkfWT5n3+QIoL4CWm+4dovpfKxu9JF95v0zNKEn71Na1AusDU
meMiFKwoe5ivDcftFxHkNaj18ohFK/dVuHiyD45/ztQLN3YL/eo9qXw8buWLvvb+
6jZcDZwwJXts+5l0mYBYZRma4/IYbbm3Rvy0jD6h9pp7wJWP1mhv8A7rCEiMbQyf
Ym3Mx01Rm2kqVG68qymCL/MviaU1o5IThqaltDQfMQmw+RwTvjFox8sVu90OgWvs
A43qZXDCkMU7FR7BfvrLZG/f98KM2UQ1dxRZWcKEhWSoeTa9L7QXR3C6OYZ7bBd0
1yes6Bu9hC3wxyUesOIqTwEv/ZlJwcDcsbRCYrPMFOEvenEEjQcnJ4R2r2uNnClU
3i8a5zynsnmlSPNpSB+8R3TlktGEzt4M95n+INX9h4qLVWHtaxp/5JKWJBnwxGRb
hQWKjuZP7JiFBOj6c5mx6mWz9onkns5ArWWSPM2RPsba5O3eA56o2GXmal/AfJMy
T1p/jY1BELbyI2Jnf3JEuCRuS4bpgG1naWpbUq2MpqlwahPtIVdb6gdQUdtDorti
x7GUMOo1Km61mqYLqQxyUAJ0b0AU7+RrIoEyM4lJgx7kepzr7j+F1+faGlLeDNbK
Ag2ZyUTXLt1V5UQWgPAfdU5E/nvuYAQzBTZD0kdJk7b4pVPGTO61MfRDb9v8jLYp
HZn4wCZfYvlCjaaUc1OZWC40q/U6wk7BgBVznDoeiIT7hJnLVXWrlKyWDNLN4rC8
sTdc5Y75iu3OCGA6jJrnaPgBy/xYg08fgaKJsZVBz4uYE7OaQpJe5zI9uAjnkuZ6
79BloC0eVHyAxCHfVqDbsCZW1H+i3dfSkvIKDtIIMHcbfuMPYxchkOAYEfuHm0lS
lmzmfZnb2mW7kMGmL86cddv7+HWyBWsWA/BbQc8/X5/S0Nxr6rXTfaPYn/qW8292
a/EXK5RGtyfAf+gNvfUssUUN1YEm9F0IiAtj+2iuHE/kWU+JPdxLPsnvNy7Sp8oi
XnT1gpZMp/cA4/bAAvj9I5AlQmY0oEI9zipLKwrI8Tix5nWeelPPzsPHdBYxZQ9G
uGgtMRlWTZewZbkxawG5bkyK5JnQcfNUn38kR9+W025abUkfSGYxZPU0Yxn9+A7g
qupFAXSuIHaKByU0fbd1PEQv3HPyfFysvarnzYharpiMhnNsP19dudf5AjdMoKCT
wKMBehSlpXr+KABkGMC3RjzpS89rBIcpfkiGY/+1+vN6GcHsjxfm5L/bg5hWL6QU
FSBV2DDnm7BzUfJPhyinPO/XH9d+ai7JcE3S9fWDMcUdahQgbdE3LHm9U5e2x+2Z
05E1JHEMg1dZ8BYAtDsqhUzWhQ5CC0rjMWtYs30uPM2OmRvp1l+h8xDu3PR5jGa9
L+fqFjf17hWVZGrygwmrHOkGHzUKqdmkzscrZyNDROb2VOhrfHlHtv/JfIF+hYf9
qlwN/HMQExoZZSg6c8vG8TZr5jMnyW7bG5ArbicNJgRcPffrlXX9qjo1UYW6aDFd
EKaa9RfqJnJOrFx3zgv79xDqr8QtHj7RCk8dC6Ry6epP9V5cY5fSFlC3xuah5g9F
zf14AWS6R6QKI8CIiLK+hUQYmW9vxbYRT1SRXKLkuvm+rb2gYeTsksb2Kqwxex+u
9sNnxvcS9ovITyjA1z+Nmvj2IGMiccCK4axab03zTt7bXuD5HRESvzBLPFd44osF
4rrH4KL+4EQNLnom5oLrQOftT2e+bB/8XpVyV2zFu6zjFXO39PBSqz9VUftRx4Cc
SuU3D4pSzyiwxiXRuxtFffPbJbYdu367KRfGfchUDTGKpZB83uLPUP+UJEMqO5mn
KiHFntTaHx7miTh5XgjzNmDhnPIEG2ufslsIJhUKZdQFRmAbj6MazgCGu38uI24m
idJmGSMJBIm76p4yPxGrpL/KI/oLH8D7IXc5J83Bzlv6bo0rAPjoFjKpzban2pwg
lz4FmTX4sPtkz8E1xYIEGYlrmhBZO+fKcCpOofRgbVbH6qF6DUf2Syl3PBECfUZs
u8XgXDK71sYqf4VMYiJfcwNdMsWWQH/Qq5csExoKWeGTIMBF2Amu2aoTINDz0lC6
vZY00UU/1luv6Sv3p3bNpr2cj5+dRE77PDVPn/6tvSYBE5nB1Gg/bJQa4rp26EFl
9eGQvmhxDflMvLTh3imk4xCYKO82nap4DVNt4IITSMybkQIO57RhyJuyMOsy41A4
nLQKG8lUgRPY6fOzC9kL61uDFDm9qRqhRQclhvl8UTi61x8n7f3mv/QwGOYh81D3
K5T3FyPHZOghNXK3wXE1s3zs9iZWi0i37t2R+fzghbfcXsTZe9s3MLwooMq1sKGT
qN1sVZi/6539hiVS5mXgmHAHrh2HGqXBvzmRqVBI+X9m50/l2qynZ3WoNAnurfZQ
YaVNmDIBV2No8/f1QF+o3S2hB8EGlAwcOCSL3/0cDpFFtlaYX9JOeJWomYJIGh3T
2e+PcpBspFne/EWkGZK9+ItYE9IwnkSWsWq63lNlIOSybdjvv6MBUjhdPb8Hz4Hp
nN2JNo2kv4ghwTClPzslJ1QJ75mF0ApXhSFxXDknsO3wLAShkbNgs2SKF0nfbvWf
cyMkDlQhvYHusNRVRrgN5HyHWtNhsopFjox5ZNoepFQ2nVT4mst1Vl7HboZD8kjm
dusYptb+r01vz8LToXECKo8TwMiB/It5SY1M/W7fwzAfcNXVAWR9veGHSDLh+iHg
/7icle15+g5GvcenCL8Dghp9cJoQ4yDe1r/90qsaF1ryY28tXDWiZj0YxUkPKTys
GHDoi/EpKHrwcbO1AQ9y6HPE2vmGABRpViEWjItzmtIsvidznRe48coOE+2Bjron
E1M/xJSp9kzjz9qRi6/w5M8WHDcL5zT9apBf75WHKotb6H2ndBaUJarG5ekNjZet
THz751KuHbGCd2kxW7KUUm/ab+WfQ6Y5eLwd2Gf1V4xJLC6bI9xJ1Flqi9IfJWfg
E6Yt9PbAfa4zWHO6GlTRTcd1pTlAc8/uAh+vNqdkKuVgGcfaR4vQplDPU4g65RbB
YNTLjIHFXJ0kTbSJTEQ8S3y5ivxDo4WJx6ElZBCSBjdklRfM6TAi4ruI02/M0MXX
VHu5uedKUmjeJj//+6e2O0c1d/sElERvUOj339vQnsHbPYKeVE94QPtD042TMNjZ
WrDAoQCCqwPD2TqvDM1s9kYAHDiFB1LBdFy4IkmfG16YN6SwGZtgGV9o8u8mchc3
R+mzllGzIvVi+YeLLqSzAxCn4a/O6KEuL40ADiHavzCM2JWPvx8h2n9gP9Z97r1N
kctIxPEIlmM+tg0AKZYJwgF+qk4HnSHfp4mHr3xjKN8qXkv6uxdiBWVoNiBR7yNe
KFzRIVBuayDIC+AopVrsIfIRx+w52eisQRf1qHXs+gSleROij6hHD/lczUqp7MND
RTdCi+t+zWkSrhZIlBci9l23p/vjVdWrl0zSbE1LQ/3yQhO7r7fcej+/FXuB8kSC
KmjCtbU3qDnMVszgkX4qgzEx7SsjiNVHACzS59orfS4QdUqZSZF9nCmU+76q5Cw2
i3asDFqj0NnR2j7+54VulowV3HBTnP6gpkCvpe6TpC7NiPFe5RCvi+CFcXcvclMr
uxSGmtbGwwPgcG3wUd3TwMwnp57qRcXlu/dGmz67K00FTspUwERWsG+fqBoQZ9Wx
i7J+89fw2trETaQOrpFs/ZDKCrYewco/N12JZclI7XRrdHfaWomcj/XHo+2oYAfy
LaLabWj4U65d5H3+Zn33du+VWbw/sG9x3VAsr7JlkuOsSOv6EOr9WJy0Ylmaj/Bw
p6BIcluebqvAQ9Cr5pW8rCV973yikG73vutV/XwfthP/xQQU7lef3SFS2V+JI8jh
h97y/5KuD0M9NWvW29G9eZW2gC4cIBu7CWJQctkcg5c0Rng6PeHIFLdcvBqnbEwk
Ey5c4fl/wjf4frAuo6wpkdt7/j5MZj82tpFmvjb6pLkdw0Rz09uqLOf/Dn9E2NOH
Pa1qUYg4KKWFSh93ePE43TxBGI4WHVdKlOJDDIb286W4ys+sv/0UmiSJZpe7UA5r
xwHifT99Up5o1Es0i/efD8WnVnkp1+KpKKIjQqN25TQNgac10R1qmOKfCUMM3ikZ
4DWSlYj4ZV33+VUJ2fBaXSvJ5CG4N16ok4t3gaxexrSJQsw61tibcJEglwcLVHoR
RpQO6vFDUQ3azUaJQhzgnuXED/yzaR3aEgu4XnzG2KFyqZy+an5w/MJy/KKywkUU
B/wrEwm1zc+pNbz+1FEIH96Cu4avRm/iy9DFEUqbVAzvh7HqDLBJ0PR3k8Rw4mmI
YFMF+US9upjbWs8P1MUSsCVWUQec95I8Ca2NVOazQIpqD20sM2wEeBkTbUyZ+jKH
F5BWHYjEzk9CDJ/ciN1j8ERxt+gjVoL0mbY/IQHDQxNttBou8vn+j8sn2jZcabbf
FMpijAHC3MKVoTlLXiTtNSRLPIOF/7T+QJWvrM7JP+1/WtoSNurC/O75Is+OMbYH
Eyc7BVYLEIUXp537hyzu5Qs9bJ871CC+6AT9El1hyrjXzunawj2OicvCf+EF2YKT
kg7O3n9sEs7TKwFYdQXpgeFf/30rW5X8XxwopnXD4jgGmMfkpEuFa3dxCylGak7x
y6YZQTSEywkYz58OM3PzcDEbQbYtIuFVf0oBwAP7DKDuJAXNif9817iKJS9xc3yk
3lbiF3EPuW2CHwBqXKlK1jZdwf16NqcaY17RVxBXgbt1kGVjcYfuG6ESyC/KGKe/
Dn/nwBTmgO7iHeSobEnhNrqPSdVgbkKvgKtXQvoRNgcBybqHOO6STiBnERjgObIn
RFaj/ZTOIKTug7c4ak71D3kOJJRa3w78LYJMYpwPJ/+qlM5LvGI9vjFbL2d+XEei
SDcRUL/WqkeNnsMe6alHXUi8ap2hXXC7glOou//uwOQdjyXwFK0KXOXoOH//e1F9
Q7fFwoRcWRVQW1kEaBKUnLj8HM7jVp5Nz3fH/iP8WE4Dq0PI+IH7IJVIpGeHu4Y4
PLrevP+UHFNmoSoFlysKBzInTj4uxSRBuzgdO0CWXABMC7UkZQvvS6An4NX2B5AX
Wqv1RJ8DvI0dEze/aOqBxkpcJxjfNQ1PiQ1j6HTU25ywWXRgjuiMUObSzx4ch56V
lGc7GQgXwKInZSpD4qo3SVAe4KX1f+GuOc5uy+RrEINHozJ30gR0S4lXPq4RIOA6
iBcM6Bw3d7UtSg8HYxzgdGxK0WpXngxUBJ5gm+qFlgFaPniB956gW1CyMSZDgLsQ
0qQl6ykp+CCBmgyZRg2AJo9NbHPE5z//A/YU5gSF2cb39OXXHifWJQpaqc2skfXH
7jAcK9iHPyAN4j8ArqG20glaoCs8KD0J1qRsLAk23VSqiXUrkJk/livoLldeygBU
iAtFbmU1GjfNb8FdseNJ8Z3brH9K4SEVuuz/iLwzErax13HB0sz+PQmIEza8Xur9
XTmv+tUY+M4hRoHtBilT93t8ijQBX8Qao8Rx+OTqBf9yxzBltBkc1C6t3+UFpr+O
VTyuGEE+x7olcFf2KVLPqoaqpKGt+TEA/4Lydk6Vgi+XrxNo76kntXa2CJwonmzI
e6y1AMyC63gaRixynPpG316g/VizKYWPhbqpN3XUj+H1WwduO+vmH3rkdwvUymvK
CeNveSbxI9dVjpqo4DDWiArDYehyqgMBUqljkEFDw0WW9BkH7xn1l9OV99HJjm1w
BJEyQtb16+yobzNJ+F8YNqJysq0vH/7Qm+gwQg4MzzirrF7HLkzsj7Jd3yiill5R
vZZRzL8zsMYipOiQFhP5Z91aL7ItV/cXD8eNlsD0PoG4CJtZKH0TyPZcNQHB8DQV
BbIK6ayHEvzZq+lMdoOW9HP7U5tKSsN29giGqw0GAmQYo4nhOnRoJHHt4BzOCsAJ
KmX7szpO1vxyWq4k/dYM42zzW4J053IvSKiOp+QjCMlTAI7oAbhwVAy6/6oTOLEE
mFuwOlqfy9XEBVhXOeHUamEFyRdUX1Rx22ePZUx8NzFB+MNddqyZgXEpRpQ6BoCQ
/3+k72VOz/DTz9ToSHzt9q2eELl4BbkGXgXgj4joHEheUNZSnNeDeDQpXjRQVDr+
+BSn4EGN9wUrVsAtPdIU9A1rldIS+q9My3jy1q0e7gOWlWNmFKp4R9m8kaXeAlVj
6sOCYR7qNrMr21QeRJZrnHt2jwRpMfDbyXC4llCo2PzhngU4D0hJlphTvTdc3GdZ
hPaHUk+ohhIumaULXE+bPpE8bEaTm42ynaB7Jo5G41FZlQDXVHeHEVgnsuhthC4p
19klPkNGpF6ZWAA9YAPtda/JEGhOwWZ/rhaxzu/R1Q2CakZVup59vsXeimn9MhdM
SXZL607EXzIN+jX8WZfUhGxnksdPmzcHa0Hoyml+nhwsjNBgiBNzWj6WiLjLUsos
3zZGJJfxtasCzdnzQLYhS1CKXlTFQmtS0cnxivk/lJxH1JvmFvDVa/F9HX/rnQ0t
thODgiG50yzl75MlrPdDGyJsbsSHK7uuTEUeq6knXTvIpMxLzwVTk9B177b19+mr
84sU8HydgApshlwACTWWsl8x2YUxOM1OPtjPAXYE3qbFbYCOgT/vKlynpy7NhN0s
9D0csTJI6evDXMGEflcbPSTvZfx9Kju4V/stGQiy5EIVp9RllkQfVcabELJMZqH4
jFKXI9tS302bzr/54CFmgmA5AAEbgrShuLYusm2h6UDRntkWefgbvCLSUwtZz+IZ
HodBbStkZ+IM0L6sYoc1Y3pVC1/nKC18RU2N/Dm4mW5JIYkHBiNMOXEeAzgqQ6+p
Earoqo7CB81oSAhbX43LtZ9ux4H53Rj0f0Bg2l0c3HkTzvBugBWAU0ocesW26DfI
SM5B1/2qBQLO51wqgEpkkfZf20H54DB25HHpfSmaTzXYRIoEqAKE512bTiVc1MgO
2T6T0am3XRfnCr9Y1SGTDyFkfb3WWNNHxVSq8k0v3hXTcHtj5TIBMDP8ttAhLqvH
vVaAGPMRpAHjlX9tN4TvGJb511PQkmOu/oPJqMo8kYHB+ucXIR0VJkRwlShlC6iO
Bg51f5w7FMSZ1nQAQZgrF+mJI/HmA1ROvZMeA6dbpkiKOry8cgeNL04mrMcdyIFf
mYcp1KjCGTODKgzAuF+ymE8IqvYWrlUFORi5aBMj/BmLs9E1JNvKxbJXwtVmqSI5
iV8r+o1hTsDzFJ3Tm4Ug6c7aUAhQ28AlC7WY7fJ1q6MWjGAsZVHqGhaIt0sUalfR
pardwQAHAD7hrVt6GFj2oDxRpxN6br/O2ElJGCTR/FJNBHy8fZ0IgXVJ5YSs3qCJ
5UCuhh74TcUSLp++n1lQF6Vudg3UG6SQrCExy+xsF/A1rVD3Mh03k11984bz1NfU
urc+moShbJCMZIRyQt0eQcT/QBVPgwYonQDFTikFxz7fky9xIr4IUkLPVXb7+N8w
yF1cdsYIMgwXC5FgimcGDGV/4U2fFVfA6sYgR3GG4GDvhILhBQmHXWpXdrvR9ARr
tJwCYxcbVNJSmHgjJDAg8t4Z5nbiN5yCIgKsBvYCgCgVsu5HGaxlryyfm9qsEswe
a+eR/41Zt8ZG8+HbyL6BvZWJ3aIHLZ2n8264FkZuSwgVO9PpxcBtde25reJQm0o0
2TiLh8amS31gPcHQKT/qmQaoN6kNOC5V5ushNa6N97S0RbIATKSwy0oyl1f1J2tW
akeY+ADc7XKM3xxJHwtYN5e32bIkl68qKaMGvwTe5BfFRq4uu8xe0C+7ABBTfdB8
NTeV2lS66xv33UOdcQgZbbSHjBWFXdR5TdRoPdcBL6WVOy4r7KJ8EElQ0xU9oY2n
4pFs5z04PRKqqZMvfwXEnlMFyG5k30DL3mhZxjeVuS+BfsD6ECRmDjh2mpJctf69
FzzAlwqZ4r7RG7wqF6GMLKmaCRpmgHetJiOKvW1+LAbIta4HYNVQ3GxVQAs/yh5m
bVhavvi72QjwU8R7cv0roSZqyurZfadzMCuCFLbaLFFGuV4uF6N+BhB8z4amZXQR
5SSHl5AKCHpM7qdcFaUx3J35ZHQsnXRgk+hbc84YC40YjOt9wejynIQ9rB8i9t7L
8PanVgMt6sKiZD5mhP9yr5F7Lvu9GkYpw1FiL3rb+WKE0SFIQsDGzu7mMn+s13Hw
e9tp1j6WZ8d1Pao4WEDyE2wFGAmHx1N+Jw1rlAhuOLhkgzN6jEB4HnLfTjDak54w
SMx6gsEq5pXqkmNVNjLa6uaIe5XbjV9vk2z6rgOjKWSrOh8fquZw/nuhNZRWCcnW
ehy8HwhaZeEHeFQOv9fbb8DmFIYT8vQeZFiIIx/aRul5cYNaiV1Tl+/Y7UnBDaYg
t6FNLyp7VROaqZTfYPOxEtgAyJaYI8iM4SDKLnkfTokgnyYn24IEinEl1DrRBHkm
IlFfDHVeu+Grppz3cIy7wSxRRtHKWB9RppPmzrRqu9j9uRtmLpK1FOZzqYvoRsbY
3nEpT4x5GhIq/19hWoItfsdh2heB5w1mRAMdjHKh7xFCQpf/k7WQB3YFEbTCWyc7
A4OHCsARe5UIhOg0j1HDaTopUgGUi0wiWti5WnEeloe2ymj7Xd/WQMU1cCiQOFN4
ga+QxM9rDE0tfISyKJ2XkrZEmFLtV8iOYEq1vqgJexZBq5C9HPcclxibeykNZWP7
XsMpbqlH8AUFmwxvN0W4uql3i10R/BCKys9JzTd/y8X0iG+noNqFFZZs0juR81x5
BGDv6batYLHxEUQjMxDFWh/UkFa37iQGvypXQMsg8NzikRgMdEU5i1Kry9xqUrya
+SZaJEr+TreVxP8JqAGXfmyOLv7i4UBwBDj3fsxkO5eMvyN6PHThjqy3lyIv+9Dv
EL7ozm5OAl1tDhWHoX2NEJvv5jO0Pp5TXDyOihWhXvgBqpu0v2yIWBZPWuAnGhbD
nd70c/eUzk645Fwfvs/p8+XGVGTmWpvASbYn2JdIT4+saqf9hW87u1ZskhRzWJrP
qxp1mfe8TKhJDOWvtJhsmEjXuqb64Y24LO5XiSoGmkNCWuR0Ootxh11ME/yn3/Yc
Fqy0OTrKKYYgwpydTpzKK0fx0340GgHX6ds4quVzpWf6rDTsOMyZAe3Jd3oDgT2v
xJwaZPte6flD30ZkRz3DMzGenfrJN3NExcFhyYludOytnSorSJMYGB8BAQ7UDY3Z
JY4cXSPHXE0z5Em8QHJVCZRZCP4q9uFXksY3+EWi3P68YTAgyRiDO0/QR42uP9PK
vF02YvVZtJn+/OMWTxp7PhFWU+DyHprRA8EaoxNlg+7jjX30abX/+piGim5QgfOo
MWO6+/pi80iYXOdSjMzeiCyKAKEduuCEOo5O/VuuRSXQAYg6BawCzmp/V0n3og0E
thXOY0wQiUpQqRJgb8KOp9REJamTvA+KXOiUkm8VQEjmPJHs2g1LSwekeVnwT7q5
Z+a0zrLFFLF60PiV64Vh9VgO7GivCJz/31uFv271yyZemThHGMAMxt9yl0VzbvnZ
VY1ZlzZFAWrrre3lUYk36zy/LrJqP/ACw0N5H9Bfy4Wm4/NS9RhnhJPO1WuhxJ8w
ZUvayKTNo5+Ukd/EGX+XF5thVphr0IklJFwrs8qxdg4n80dZGedqhgvyuQEx+bkV
AooFPqOS6wTPxrqdwPQrEsC/8FXuWao2D0IwWg/5wX8mRSDW2VKt1/tT4BZ0pagQ
TT5L7laqp3boE05+S3FefWnuchPY7gCoaBoqEn6m2XY7WjCXaa1ZekFF1HNYzGuu
r1qMg+e8MI643Aa4eMosW3mGevSnubsMJkjq5LBrzSXwUFectwOK5fp8V0Cg1kbS
nkN7hCY2n/q5FYEIl/PwCr1ehyX+erAGxI9GH9lLfs6xQ3uZNcLCtg08+XqPAgBS
vWZ0U6+4GmBOV14SmmExLPuiC0iv1WBT1nQ0tMCpCotHMYcjOtpEMAmbbB16afWc
M5AZkNQ+goULE6tCMqtxCr3mGpm9vCQE6FZW1ohhv7Zn8o/XboaWI9RXJttLoRb/
jb2jgIcQeXwy8RSMnOHXTAaYrJw3+k0q6MRhrH2osgG94lsiFQtGTvxzQ3LMO87K
9rMIGBu6f+ebOqHTnvGXsLdN2euj+oH0umMCpzNbzt1miE99PTMmiU9WystCWc6o
DHlFTcDHgeIkOHenIPo4swzpR9mmGMMe/Idhq1KR40p6U5G0A/M18Yr1IV/1cqh2
dkXfRb5qmCwhH/cYECCdGu3mFUquTjldfgY9GLoBcID7TMmw1vFYZkr/5sYPllv1
MZASW55nm96FbuVc0O4tC64hMzk5wnRzGo49qCJ3WpUL36hBhmR73yY/P9qzo/c3
gV0hQfvdxQJDNetOUWiscmuF51/aXQi2fAWx6gGKYRVsqIpir82VfIPqToqZnSVx
kTA9XmUJBvqeb017qkVJxWcU8fXWOjM6srj89QuWEJEm7SXaDpTo1rkMMI3p30Bd
oysY9hbCcn1DpmVRsrU3vhrDnXRmfM21Cv/GI7j8ZqC7TbKqMXsVLy7d09t5rDyk
SoiH6KBboVRkaJcvCBkQkc7ajxPYMb1nxvB1Iqbu9ee6uArAjMjh3D4fp1zT3WeJ
X0ScnEtaELEytH4l//qYYpyBltHDLOzxmLd0UrHQGyaG7kT7XBc5TMFDIif/h/kc
EVhfyFOlCi6MAPtr9Mrv8+APjffuJghtVr5qbNXZ0VpDUUonXGFm23v4Fa+N7wUK
x+Hx1qqsbq8bqJ4/k9pZ+6LW8MHxHosY1kgaCbkMlWISwrvvdIBAnfrxfposBGnf
r22saDtuptW/x/DwbCxIBMA2GpLpbuDtrJXPQ1X6GPe7zi3/Ol4IoL/RFjRvV/e2
Om2fWZa83VhIKIc67k8D7PKLO+RhTyhTR71ltX5L+ttF8o8V/SPtooabCkS4W89a
w2MmpY3P0xozKOrQy9V1mJLt4VS2VYXAm7hHKoOa6v2DrSv9zamDR5LUt9wvn8ZS
S3vVjiTL2B0F914bcBLmevh6yZHaom/Qi2BowNQldPEpqjCMTW4pbw6IQK+8UL8l
+sWpox58nVgA19Vxw6+tDwHpb+kVKt4GMhNb++pNuBujHnNs+1vamU+5XQg+aHw1
vDHa0xwLc2oE5/E2xH64KVl9Wt6sa/TR5/1ho6T4eG0GzwHYhoaNnCN3B1YTIypn
zbohouxC42aYGHPxpb+wb0H4P76CSFoszTcdQOdS+yLFe5k28mtCrqh4/syIwt0M
9NoKRRjz1cPjo3ZlJmV4p7mrFa7mTfdhPmeSb0KtWYpgmb1nXBsfTwOd1pyLRWbL
2S4Q7CLL3Y4eIFJVK3dnvKFDNWw3WoEdBg2EvwmzlHzRO/gKR5Pe7ShqrY2Uk1nN
8yToXOZiF2tRXraCA9DSGw25YMmNwA9QxkFsoSPYZa0rtcnusucFCj4GfMfjfZso
M3GZg5vYdP4CVYnJLm8V3Ez8VNiCRAuMi+cftGvcimq5o2HJhThA/vi70t4n+wm6
kqcMGEk6JiYljj0peY+5wq8FrPYld7EUo1eAVkwWUdzwtP64wGegA2ebAj5wsW1x
XeM+pwBeD7FydDAC8jV+AHdCbrDpxmJ4JEGxZ9OSigR9ghg/k4iz0SZLdC5QS9fH
5r2diHIs9nMi8L9vjF+HeBFU/RpCua7PNbNbFAaeTwS1ROwZ3LABqDI6Oi8tsCsJ
9kSfURMPpPSHIItauWL6iApZMmxD01eTNQgJVyBOKgSqeN1F1oYhwdG7uUl3Wsar
Utau1E7ZmUsHLBihL8fqTbXnFNvdH/tfITAwsc3Zhjt13/hcRXyyenNfJkNx6sQs
sf3IhmTY1s55ZDW/yUOw8mfDGge4SLFmrSyJCtht29k4HrVomsy4xWC1+B7dQC6F
N/0C8BRSKqwdHDm6xJxLxFjNYVaNkwtRHHxDPXUg3DIXYzupk3hnjWz9DPbLKHgc
E3Ngkd/G/JfpjORKFd3fU5wg8ykLzMyOtYxwfGANba/nG0UZdZBe/CzhIYZtaUX4
3Ck1peilleAwBq/OdeSaIN91/mHesFQgyUbaW3UbIe+4wZViUZT/kAlZGVb4aKgT
OTfVQ1nboWaW+uGHVtXjvFnBehgLNdr2SKtjrTAZtZYkhzU8iKLzWJ5dXi7uNusQ
tx43ks8Fz4NVxU4ZbZFH5L3b7PMW1Vfx/a3alohnJu7OJEeBJt1VdbW5Vg+FjDaG
RvNDSCnJWOPHSvdncm3zAZNd7pazCW50rnrgzNXvuLRJolEfIqsuvkc4Gb2NuvVl
czhouZnwIAJa1jXZt4HXWFpdBYHrixNzibUZFKpLDHFuuQ98d4z1t/guMn3JuF90
21vq1TB1S9dYmZLvXUYzlC19jINhKVs2elkTZjCvx6BGUvKpTubR4MeabrnuNddG
xOz1qz+TbiFg4E0WCL4Te5Tz3MA1nRuk9aSLOt+20u37H59IfhCcHYJ+idA03HXX
INkxkEJK7HxtifS3dB0tPhE6kHAXQDPJ9IU+iAt7upmZ9ciipC6TmNZf3vBZDpVV
rxL9UOMOlBcr2iosaUfq4p4vLxg6PToKiy2awpkElhggMU7cmZQbsQr/HS0eOFAd
msQKhTG99S4ukfIzg9rg0ZC3dgNAa7wa+r5Olh0BXQ4nl/woH/hoxyI2yaQod+3A
Fkwfmp1OFAUSAAMsXV86KU7BoZmvejh/GhmP50GsbsJdDFASVikWoASf0cDbvMBn
IXdlC741gWL2vwNCLeSq6SjFuZoAxRk4uv2UbRdz79emO9+xapJSUJyTNH9ZbtC/
XDe8yRTe1b9cXrjBaAx1nEYlCSpDzMa2Jh0JqmQnhXxGD79L+qaaXk4K2V+RTD3x
V23eWJPcJrVzkiU+6EI69kSJsa4V5HiVmoDsd9nwdW5S/Q3PZly+bME/Q4vlQ52G
pfNyUKjKyF6dntu88AuDzsy4xf5pkdG0dDzrKWjHIEFNpibQZynUhltmEshQdhrj
LzusdX2KF5XfUyKtcXVZ/WYnFFRyVl0EB1PVZu4PGvk/29vF7cWkOBx2zCrJCjh9
7c9USXDYm05YZvNE5BfSMsX42gQlNbsTRQ8P/mjsiVFyT7DBjYZ+V9Lw+kDPyFxf
Lf280h9p3HPrnJotp4H8JizxxkS5SPVJYtlSjlOmhjE++8Dq9DdyEsTzu1gDnyTX
aUc6gAnBsmxymLm/s+m6xK7eQ9P+LLWnPMWcxFWvETomiLJUvEZLAnuwUlxkc3Ff
HtyWCsYbEd9QtOOlKUKHwW7uIFuRP4YUGo5NkCuchL0Stg0GdQWk9bYB5qJWU6bE
4Gh8FS5+ojX5RaqIt/1OL8wVOmaU4eCWDKZeasXpH5RWC2HmWQtzAYB3oV4+wReg
/liaX2eIoEX3MmNkScyMiM+ULhdn6QKfftQWO3amjGhCLVCeQbs3AkNJL7wnktzw
3SJj7NhCz3ayX3ZSFb6xbrwkPJB+9wDVFVSpq1OSBdpRLiJTt2t4IsvsD0S+nKGF
i2vnE4zObH1ZM6meka8kFq3zN/TOjUC4k8P5jZdbVYKjLbH2PEvn9yOs3JWlGeWD
RWfrnqEhRgfo2YWaiclRIilt3GqBMj58aweOC0VVVLMXiXMGX4kuyjw7BlRZOyXL
ZRvp3n3r037L+hCjumB5LKbfDqGix/kNu0sLCR8BVtfzoWUvSN4x27Z/U6W8p/4z
p9Z2ddwfAAyBJJWU64TJzugds4VZSiL2oDQmcGf556pUN4bPlvLMn8iiwCXiREyz
x1sVRtTv60btaEO/csHJfeJxnP0qsgPN5BZucV6/ozE0D2QzWMdu9P5+2zzKTpiN
zfywtfXTxhQ9F8CRPHnybw21at7NlOvDsAklvIx7WgypDK0ACX3+eW/6RkD5m3Bg
0/w12+FmLr2Hk9OhOQfnNDOixj7U59gGweDCDJGRRlMqtnuJZEhiQBhai4pcVpL7
/Ca7PUQgC6r2nDmUBPEtTnja0HV2eff4r5bFsdQEhKyobmkUD+as/WIATL1Lg1ga
GQAX1NYJ+zLt7vODdpAytm9Jy8DT2zk94132K0QlJCJsEAS96fZf1XyszDRs9PS/
Xx7XmJLt/GjL11IAme7l0bA8cITz8M0EFdAUtpNObRpvAID4ioUQboanW8cbM3So
03e13w1fiDNdZzEcFJUU7qs7bL4+I3CUdSJZFA8Yp50dAPDWHKnuQHLazMh2ffLL
pJWQbQnsZmL7Thw8ldnqRT6p6R3DHmNuSz+5OUvXmnmImFIke0UbvbZ4Abc4qTOz
yAv7XakkN7t/RA+gWjBGmNcl//+LRIDeLeyzQsiKCY3zoDGexYqZA7rQg3x6r3wF
pDJFf/m6hVC5wCzISNyh3tNB8NZUX+91TnUiEt7l4GwEwGgkxnuUymbzfJFlXsLg
OMlwnRLEpyIlevXk2SFj0TuoyPETadpazRCzeJ1b98MxrYWfN3jYgnoQsg4N13Q2
DwdgyzGPOsRixQf9EiwKw+abuF1oqwF01d1Pn5GLZUzO9IWzW9qHHN+7tbfLZsmz
OpcXguAgbYoDorx34TBdAOzxRn9IGAgO4rI9kZCbuQ9UNrMKar3ZmyNBbr57gIDw
4x/IlHVA0DFc+i/pWiZtXzoOjVuKOaOwPNXaSX3LndlXBfeTa+UNSZLOKWQ745AH
gB+SCbCKCttSElUBdASQWYdmRHjiS5saKi2xemu7a6K5bdKJq4LrxjEj+LF05NWx
/xXb0JBheYGeZu6+mntLDKPIZSUUi51qHgD33KrHVOoWI9qHVD4d3EVi3OmSWqNl
IfYdx2vmMEB3+VIry9ICzanDV4e/Rm6IzvNZhgkTISAMENoQ4sA7FbJywwdMCfTy
F9FQwBt43vn6ztxhw8a8BhX826KtinK2C/yuYJYk0+gsD7ll2Qulo4Ad61+47++J
pU7iA043FYUxAX6WPz20b3zLc8MrhKYoHORVCT010CuvCes8mJWKAW2HqvVy0i8b
RL2yN2wj3sVk4Fho95iud9Pd0RELUwuQ2hHe61Sd9YSY7uPqS7pUEed9LKuWHtRR
qEVwj/LmCpknxm1XUJusJNIVr0tmBXH91h7U7XZtnJKJSIBWrLL/peWRC5J2AMws
HxVRituLl/rYxmwu3AIBu5Xze6jRacLkgiqjxn8swaKw/hqPrTiLoR9nQCwlqtv8
sl6w/1PFg0FKRlX72hzIYQ8ZfBqXl+HbsdGnl6ignld/SjQxzkl24toBRScO0JwU
KjRwIWEc5eqoSAOI50/EyYPyhlXybLuatfRsPI5mZ2vQ6dLSoy0O9Q/Y9XJEkFfw
ZKaCi6OG8TUROuroBLOW2kCATNNo+mhSvswRvBp6brSmSPpO3CGDRIOLEYvqzi1t
6LbyFFKDVAtbliTGh5GlE3sqMDh6qMxRXvrEk204jVA7UJziENQr3VJlpyl74c/R
PvpDUcHPid28XJF5KbvmUquEsC7PLZUi62qQrUhKKz7g50SOrGD8MqRZC1fg9WRZ
/Ce7zv6ghl+Y/VZXHCz7xfDy/DMKKXMM3/77nb5O2Bz+/nCBpj2Ym+05XnZ+UUYw
JTwLonVuJbL+LPBruUnOY2HtkESrbBw+6hUcpnjxfVHzSCYz/D0dAc32w1bn8qXU
gBUroOyx3qdFl9Im5gCHagxNb3O6RY/VKv5ar0z9i4veSbU73reFsB0d+8hFTDUZ
6H4LwYzAG7L0Rl90hO2Ieo5r0QsgUSFTlXCmqYXj8hOFFhShcR7nXPNNGw27TGzv
rzHl7YG+vfcDx9KDdEnpcATSaUf6r/L0jgUqqceVhZN4Rzd+1E5wNjqx25wx75QT
AxYi5bNlV9y7bnmh/m5PIf2GMUgLOCFGeS3+TNOct9sh6ParM2FUpfQImpFYf2vL
VxacKcyCWoLmGrpmzTBO4661DEKav6ruiwuJ3quAr3JkbIwlw3V8fKrWcQA79Tk2
nQHFzBg04dBSY+VrkRIHIgd/aa8/PTD4dFruXPoh0zL1O9044+xMjIQYVQr5u095
lQFjTKYE35axMDu6maMWue64JO488QRUpdK0RIedrdrRiQ0eS34ZsgZia+RJG0FR
RSdgAmt6DxVpQC0Yqv/wBLp4VWZE8ri4IhpPzjepqu49cCXyBbfNvob7qICxpeOx
Y+9vow+RkIdY7+Z69hZ6vcC+30/uc1fJd5rpAjvhN7KSBEXmITObcYh7PCcFB1vr
KuCL0Lf0tuhb9qaaBARdVx22ZhHiduxyQR1jP352jCEDmcOjQV5Zp0//WAhZe4wi
Coetqt0e3wOPSZyOm+PzMPPeqwhqUwECYQTC0oTjsm5BdmCtjapTOff0nZUCTHpw
WK74rJ7EeQERc/sP2GxfyiEv3iKQj9FGnn3iAuotJPIe6k0hA1oOmKJdHtdhkG4M
oujywpKvONbH3TZUa8jRfxTGYI+3lXKGN8JBgJlFaktnKyoKmlh85wef0UMOnfzt
DeZZQNiRu1GEv+0eh+HqIwOQz4OtOjVF0fhDSwLbT/MKcik0D85CMqbvHdn3+4lA
yFwBTW6o42YKuQfTfGMBGVbZ8p9gG62QjVnzB1uSBxg/tqQuNPKR4kVcH6WNYZx5
I29QLqyTINn/a/bOSkklmLJ1iGAP4MstHdaogzEg08cBa835HAYsLW+x6s2uoCyB
lKu65yMy/coV8pjmdghzkPxrl4WLfjdJx/yALKVmRjNbF4QBAG4/JykeFN58OO3s
8C6lFYjcrbpLxUxV2jM03ufWLOdEsgM+9/jKCxGbzhp7yK0TRqvXLwYRathTXcGz
c9fZJ9EW+tK3QN5GJkfjNuIjWtPXmBV9t78/ooO3X+T2qjJe8KaIjvq6eFjq+op9
2ktR7IPzTsVyLKBjZ2JCMnCXabpUHjtF1+RY4CKdCzyz6Qj7LG7X/VsmDDdYybkX
+i6qqJhyx/o27cXeP42BR55iaMG3sIO7uLL5I7g1bmVFUk1N25Rxbf9sIMEvdLCj
U/ztcIv6MaWDgxT752stNwuSQRfF77rUL1iTmSNbwwsjjEa4gs8cwMNC9kRic4nT
DMEALEFi8O+KBUUMtEjPE93zlLtvqQd4vvlo+YDWS8S7jMYVCwpXXQeRqM1Cno4f
LnuVqKyhKwtlZ4TcKsWfhsBGTLPjKcTNCK/72NqWq8iSsslPWsVrajS/ZQoUV+pM
bAEOWByGexRiYgn3qRI3RVozUT5S/7xMna9J13gwH1GgJ9d/L6WoZtgla82vM9p3
/YWH57VQsoChYqxZ2c/coyusWU4AOzmn0EWZrufLYkhBrrCA+A5qaaOThVd9NPX8
6CPSAptgfKkxXVJDxoc/bDQxnewXLfw9OxRVguuDqRlQ5aKsXV8q0abp+ODPw4Jo
u8iDtONzO5PUHr91pfjDpuIeqJYOwoOEw006fRfszbgV5lMJ6YcY4GsQcMZtO6hP
2xmzFRfah9lQABsgUWFOwQb9EPerbRZc5NYlISaPWyj0fuOUlq5bSnuZprQm58ut
sj57MJPtxaFHq22Sm390WMtq0pKnIK3xbWuTaiMnO66Ht2N0YvNu00EFfXu0Uqon
sZETI4sUUufWtBVw9+czaihd9KzmoyaNu1oR2O+FmHnrDkS6u8bqqgsfqZfxK0To
NAoh+5FtYCEmG3h2YzaIj1adm7QGJtenLVjAe+mb9tnYTJOesvbyKWYPQCRZlJMS
0LP0Iy6fwFQtGQpKr2C7ToT1idbheII/GXctL2+sOZIFqYk9iggYJfsiIyjahLQP
TgKtY+HkAQRB1c9gSkzPFC/5bGyZ13i/NMzrmV4e+V9Iw1ogmCGEMnXXTzzAz1CW
gox5wj4EEE4nsOAhbKNspiD9XavMrssWcOfrf9h7sngwMFa+9n4X5W3Nd1PD4cIy
73Eu0BdMFx4lHLxg4vQKyQ14BQvpis4dQ/iMjum8WC3mRbbHOODNg68Vhjl0HJvY
z4RhGOwiErMP4zsLJghtl9rJK5y9cWLFroanmtcitrBh2cGfijP62GC6XAc47V+O
zkAzyP9K+oSkiMV8LDTJKwED85lY0jg6iz2M8TGPAVsAQBU0v/Lcr+XkiyaUi1VQ
E3p0ztwIDQL/veDiQVwD2JiEKk+9gK8CRup8KxMXrLwIbmwL/hrciM/Z8eqvogwi
5y6ByqIZsd2EKG3Y9KrJZLD2pbcVHVN9UXzP9jYBS8APV8u0zRPfft7qpn9x/IXC
2XA7VJH5Cn5DU1TewRkKfwA3cEYwLVaPdZGFYlKrdKBKV8f8gG8GtZ3bBTyAbmjX
ik+2YPJZYNcxxUaFa54HA84C1JfMgaL94oxSeDptHRspSYe/kY5rcugmr9CKBliQ
FMD7ACb2dJywLwPe5823XCVCETZZsomu8aQaoU7Us0I7zi9WlAbwwRGNfZlgxSsx
Kz191f8KKMk4HK5Phbamh+ktFO5gQVLbtmyjFCLLAW5eeGFoaPtWOHYxs1bB9JR3
13BdCKkh9V8l/n965WKXtsqbj37pBKExzi9RioKyorxOeBBnBaQ5oBqt+lborrzn
HfWZLZl1p5YIsKyHUAobJY0q94krMVwcAdKz2ZhXa4Wo9EbNwo0NitsT+GcuTxkF
JD/ZkupoX6ES0X7eq+kWlaGLY5noKfEu0Whhr8k/sFNq8AkEgAsJHSJqNxyxfMtL
jn7WImdi42cwAKruEeyVTDBWYvBnAaqKQt70z2Af6O5Si4xx8X5b9m5YV0FcFh+O
5kK+TraxjCZCYicqMroZ6xiBWh3XYsi9+hjZ1VmUDWe5SNUjXeRR1PZj4N+wY+BW
zSzB5jVdpTU1uO67EduEuEXOOOjz9H4Q7GPJOpjCc8FTtBBATU5Qb4d5LjomU6Mm
tkyeb59GuQIWzE3MF+lV7uyGBNcXJli81vBCYo2Ttg3F6xqzoO4y9uIrGA8ueJO4
JndFrWgRVBytKA4ZSUdQPeNOuYnaRM1Rm7y8qIqab3w7hP9qwCFz0dHpRCKPAXXl
8U5NSC1W7POdvxrr4kRENSztqrIL663TsAE6orQg9VztpMzIx+o1Z5RQQ6//uElO
y+yCnw2KvoFG8wj+XM75LRisb2F9o90xtzOKcn07uAVv2BoqwAJdahyR73O8Uvxd
6WUX23NGnjyQGDFzJzWa3P11wcx8jQGtiiuhBX2AMXbVvImFPHDYpk0ZxvQhKs4/
vN7B2iQqhk5cU4A1htRAHsXxNi0LPhpCqWBZWpKkTTKGWwtVlusvqf5rvhTKmzbX
x5tTyHnY4PqH/ALpPnHCq38+x85dN0cHnJFbwMjOkbAfRDqkxGymbDWre8Cv4Tfx
4LwQR915ptK1jrfXzc1m2Kyc1C7tRcKHm1U62TUYxtaIwQU4ZpHiXnFdkBdlsZ+4
B4N3IGNhtoQDtLThQuxu/o3rPUhO4dWLL/1e0H0+OaTqzHjXx5mcdH7+k1Ltvdpq
eMn3oX1Nt0liZ9DnIwuZrN3FdnAvHbWpHSOs66cw/CVEpt6JInL5dqXtFBe4h79F
EJUcgz4sxZDOpRv6sxc18KGmeAjG0Kk1CGx8YW22ME3mp1rMesTwA4Dv5KtuuRPo
HnHKSLRHqeVhqRL6PXf9viZOkgxTAXAZsTuBGRCdvz/ZDg8/L15DgjjXM28UyjXB
FRdp5oDtxhmfPYZoa3af8iSshEbh1ckrrWU/e7pRNgfgieVpE4Ll15Nxrru/SHAt
8hyeha7wpckW7x4tuLp/l2Lkndt3R5O1Ntzp1Fidz0qbyhkRfE31zmk5ALlQvMKR
f8W3p8xFg0V+aKF8rymwRnx4WZ4wCpr6E3qVHBsGxpm7BAzxnln9S+DXWnDADKFm
fl6P2zrCtgobsVMCNGDsLk79Ei/+8KhzqM7HNbLoFfvegQUSgr3B37xlcQlW22hD
iXzCfdvAo80tlBGGBkHKCGXCmw0oU3kzAiIdr7PWa7M6pqvMp3GJkUVa1/HAM6hx
Z9DSYDHd7GHeeTXzURX7qHdLuwlX9Iv9GdVh0MimnhYWNOxpiS3HvNpU8uv+/r8v
REBYVXfsaM7qZxjvRO0h83Cp2N0SmWllSwFXiu1TgF/W3a42ts3656FPvwHFNd6n
dhKP6Tje/KR1L2wuOokbDZg4ZM8NvaKMh3pfi24txB1scgz9kIzR6Lg0iatWeeAS
LutHewIosyxUoKlLl4pXbzv44sfsydMzBUPTdr8dwfqfMSg69G9XrtONTw/zffUP
rpV0SHmS/D32eOe7SZh6BHl2bnctR431C3jwoeWFAv8yyYnMljpjxqi0hdkbu/1q
Yj0eaDAPq4/TAUtKYbOii9ajhyRJdYlFo9ImpikLNmzs6hgrCU/J+AC+vhYEodpD
sJwn9yV1Kq5cIp9KrSHt6oh5x5BTsBSoy8NxFiFKh9QK9FWsQG5IGjt2VVQoPxz1
X49qgL4f90zLS0MSEm35DoiyOT+FUDBVS4GLjliRgi6rrroud629rwlQOyIe3PCK
M9n8NIydyGCV3wNQ6/dXH1GliGPcjIyP3kWNzFBUNqvOfPlI9nDRs+7pSCRrcw5E
gz4mwbPn6OYrvOKZJ7w6YzdC1t5RoYruvG33il4fD4jj11qflqlk0LBkpTaHD6A0
53VXChMv6Oe+3T12nfZB49jSJcojTYZ/MR/APrQEVjlDmDWXcEt+eX0xwoj9ktEy
/lrvai6NxEIAbtEyyUjKI3rXe0Tide1vy6U6bc7PHyu08pXnkoFetNg3LI/GnTp3
PlsoHymvEJCCVq/rGWehn0cpF7Y+fSBgb6gqgm6yeWG3G2CSohIar01In6M5wrgx
T5NuhNPkLkGRbl0PPgKL9bkp5uLSc9TSpl/Ox0LSHLP9UrSibcHzuO4I9fLBNypr
Xv+GR6C3xAkSIl16c4mXoU3ArLRvuImzTkdlWfjKsA/YQVitsZIBiQlS6YKzGUSU
d3N4yrpgujn2WmQBpKq1omgSmVwtdnkrP6YFHG/lPA7/aoJiI124cptyDcAEjC79
CJ/+12cD1/duHG9ou/H0W4e/rjpTfCjqlKcAvYh3rSmrZR8Kx22qULLnlFBDXai4
GK/JaD2Olz7n0e7h8iY21tqm8rFGSrQGwI25tEZeFmGssasgp89+6hvTtsz6RNE2
0fDvmVv+1mvW88FEfbtS78yQYWmpE7e0+ILK0WErI5dmXs0XJ6J4/4r7pI/BHVUp
y2h1SIvlfpUy18CAw3M3ym2+JbgbBTa2ITwGy6ajXl8mjYDDoDZzUfJDN5Ura3MZ
gXkFWEvHHqWfSCJlaeEYF87TdcdMxMLzKigU5/hGn9qYmBPew2JUgD3BZSgLuIui
dcVpPqwpjsO3+vpLR0H1nKdcCGTG5vm32gf3PxG8h43tvjgyjMYXqq+MOGRip5sr
XTadH2hvA5vPqd9hRqVwU9ISoVc23YtDnffF3NpBlkCLJpxDC9972axocJpa6MEr
kZ02PC/62OpIIO/6KGODUnK0kwSMmQKG0f+ZEF7yeZKTnNL3FoEURW3BqtIMfZeq
4HLF6ZNt4NykFWlukGUVFc+HCk3u/FwqL5hdGluXAEFAjzsd91KSvQXhT/uN7FIy
q8TPeGXNqspy0JNJQ7TSyRjrP7Y7ZAzK0cNd+QwwnnU/fJqX1CJWtJ5WK87Obncv
3yhxi/gTeF64RzQquh8gAsz+aETCueOHVndHw9me/++O0IFk7C/Ayv4ftyM6K40j
3r99zoSCGZ4fUBUNOIyoSXfDCtEPvQ/yIrPcRieVVLbnL5ej9tmNZbnTVJwn8sOe
nvLswR6Ie5pfGQ+CM5aKNojJgIg4KItvKuVqlzQrye47vjITR+ExWNZNXLZ/aqx2
hgU46nWLAOQShpSUaZtmh9SewuXyC+Tn1GvjqZFknFEApHLmjSbshKoxBAM9LT3v
9qde+QzD2hLI1eqj2/62Z2bGidybXwRt/XHmfXPM4tDaq/v+PFY+oC6R3aFURGsW
RtuxLp5Gss3UdD2GGnSWmQyxZlF9pXpiMtI/xDtIk9VeeawCd5cRTeBn6XQWl0vf
I00PwyGHM6aYTsFZSz5fF3TL+eRDyn+YO7q2XlGsMK3YUEHiGeJliwg3l9eScNqY
036L0udFiXAxmtbUsgwfpV1OpIaxFL3kDVKysfAiCLaPw6wYYkB8g9PADaf6bosG
MKrTipPbZFk6t2sJyDCemjqWRgj21EqgCqueOuQGzr6bhDQMqYE5cwhNcuaHPyjk
hd5lHqT+feC9wcw/E2vc0LOFgfpgB0iUgmK4EG4r7XDSNgs/f1sOeZTbGxLs1Nrc
YUmZvdoBwqQXFR/bP5q7ttSD6bOaUpn/NxcO+eiDbIezbuKBLxPb0CtExEuqRfU4
WB1ZzyX7LPC46l9uMhRaunp3OmP+nFccZnVG52bkoU3HnzhghbikuI4iYFSbAboI
rsWmlAVLAjjZWAbWFoLZaerHQZedP76RYb/KeObByg4wf6HfGzIAR+u/2kWdIYH1
qW4BzWUjvri4H4VnYHBjM+EJ0wYzd0b3oGXX7OX1PThUZd5uhn5dt4O0qBWHn5nd
vgrxsXDDFK6MlNlgQ2UTRTicqefMP+0W9CiznCrMcoRSCWVr41q7HHhgnNoBt7YR
G9FpkdoHuHto96kseWvff03QTluEA4wpAxgidyJgXl7LrBkpOib/cErW9IV2ix6c
UyYbdyQq2C0PNa97dGU/HVBs4rFXxxoJZgAObvywI4pWJVOtWGhUSuJYQo6NFRSb
Y8ng1JNt5qcPV7mykr5/zJXOxi9wqVzQzkoxUNZcd31vnNRI22NvgTA3o2y9qRHl
gdf9P83AHdupmWQgM9sgXrYafEFdFYTwxaEO/zgPy2/tGGD9GLUtxSpPAEN3EyW9
kLAMTOY6V7b1mvq7SX1Y/H+pyo96UNNz7mXRLKjDzfisiZWnRZkBtNuXq5TyjVAo
JOgC0hcb8ZFwbQ/NdzwcoG0EtQCkc8gj15gLeD7a/dscr28WyT+hArHkKrR+rAK9
sgL+U2XgZm+Rix+GAr4UeIhiTMJ4Xz3IFkhTbizCengp2pAgDpyXVl/HH3/TGtn+
0lIY17t7u5tU/ayIs05zahjn6OhxIZDxEafoWK5qavxlevTzzWDYLzySRgoBvE3w
/bdXkQfrXkApuaJtVC4nDz/sLavAcLzI6gICBkYyY12a96rBoQ8OAg1kvU1N6tbH
LupnNSQVRu3pyq2l9orpaDMqTQQ9VPITNZUjWkpBaxSBywpz2xAAwMkOrjiywhdv
G7kN0FRL2Ft2vdDLHZmgP/k5hCd8fbT/S9du6Uon6gIpcQK0jRLF596lFHbEDiYs
VjWjakGfSr8SGfyx21DDn76wY4ScGknZLtqLCNd39R8qmDRYnJVH3uYdJtynFv1J
uRDZF8c3X7P4X0df0wVYB/Sify6iKQfBRT3+awT6RPudw9dG3V90hMQ+ibEZWMuh
SuN12PaPILB60p4n6QmWyokQUcNawpvTzbnDOV0UvuIdUMZEpQFXQsqNlTTYNIHH
o4j2etGOeut0U/769SkDrM+Yiesz6B1ByJFtvglingBHK0onuag/naTisoCggeWp
ReGCGrVhi7jGWySHR6k0yASXRUYMJu6r8dI48LjvViOhuRzy03xTjxd2UCWNPQ07
esxr3gVSG0R+lwHwDWaDcZt+gzKHr2bWEOKOVK5iLPhvsstf5SwhFVK9DdDhMlFJ
ZBO1sNAZKFnlLWCm4tU3cA1zhCiwWRdsTvShsnuD7ohwNcJXmZFhePg2C9WZx0RC
/70OvoeLFYY0Le3c+ZM1l2YrlcUO6G2byj4hN+PyhVKie0LWE/fjhPaDVBVOfPYW
ULaH2C1yJdwOBxJ0ezERGpcUsTB+tepVW9IcjMKMhHw1QDioSo4gDreCVqcAylq0
GjSLe5qswZ8+AzMgMQBSjl3OpbO9tBbJ9j+aW9IWJYxNL7PK+sVsiv3JITtIPOvP
VY/b8wwkoCTAukzW6SUqPgT4aNpjQ4TnvxypRhJ8BUaGIclvzVh0kb/oQzl9IkZW
tZMmKOzsdHitfInbDz17LWthg3rVOEiHLSionuFTnbk8niGw+0xPLQYlhfCn2ReQ
cFkGvIxtSnC2GaNRjpbHgXGEZJ0kkb78sU7HYlJG0z0XF04GuX7U/xkIY6iYfdE0
yrgZ7HfFMMX9c115YNzRUx0/UAW+UliFSU8Gr2tfB7qmHser9pqdc1+YI9x1/Ri4
DwHYTvRIZTbYucyYiZOvU24j0NEUZ6DefKETgz4aDEWYdvskg9CLdlYXfmOO5r3P
5SEzy5wHt83fTMNBPvMC2YWVJ3dFhczd4BXzm11h55gGwh9OB++eDC8xB2MA6SJj
A7aa+8m0u/7X9YerEJ6sf5DT8Wcw3nqCtJkGM1+puaNNcrS16uo1iaR+UGnQYjZO
UgcwJ5I5hrdtU2J7bukIxeCewULIZRbvrxVMICIFRQdbntmj0F6lMlM+85jV/Jka
H7qBKCEbyX3ElI1YbVgKoAgOFXGqgRXkWtQOsfVlyOLeX2io+XmV+elCYI+z7jVL
CYn1LVkHikAP6Pb6rP60zOSqfZvO7j5YXxQZ+wjkRXaUMX7DrV2DLPBT44ton/v6
DofuyalaPwUH0GVhP0EZ9BmZUqAHKDTbcYbNpKthDO4yXDHpKoa+P3CiEjVIJ04w
uhWeGzX3+jiaYlRx9x/0+KWv0bWJ9KI1XU82GDLnikEVMi7B7rfj0n4bsG5tFVcJ
rz8/x7D4Sv8IEZ90sn23vzj/MixpVi4hHImC8zruBJ4DwINRhZUiSx3/I978JLG0
ptOukGcliPf/yutDqGtQaRAj2uP1vz0wz7olD6XRPTSIKs+6hzzMtPF+WDJo7vpd
gcu26h3W5r+jSZ2aSKaKkOEnQ8j8zv8jPj5wAJIkyN/+7d8/0fjZRBaJD7M7lTJB
Myc98WtIa2dodjh7ofGngh8D92krOL7cG+fBTB121nWk3IDJRakvi0N/vC2NH7x8
G/1snGb0V8of/W9h+b6idH4Nv1Z5fG4gfBVy5Pq0BHdamqyobavDW3ZOI66K8ol9
4S9x5Z2/gro/5r/7xTME/i0RbxQ6/sGcUgrrevQJoteM26gv0x2HoRSsw9R7u6ve
+XzRSf0XUPgkN7EL7tfCNKyAiTadHfwTcc9GjGkxPXSHsy9wtKTcsDGMo10+ff6J
W6zOEyaOOj34EfhPXQ/Qn9QUFnYFoX560UxEpHdFnMYjDvkfGZuExu0fzxT6gi/R
nyxGhX4JVcE7SWF6UzZZkGLV6RaPJCZcKrNvkAeUiYgC5o+66Od90tqf8g55eUDE
OHWFOHLbx2am+kVJqOkJyd9SXxYFXcyGRfeUU1Mx8EXVljgWEP5cv+hIWTmThmxO
EadRImAeY1ujGudhH8s+lSQ2d+mpS/lxPo6kermwQFkV6f/EE5aS3Qkqk5A2OstR
Aj/FG1/d30AwI/JNZoio2nx8Pv0QP/bZ5LNd+YXiqxCMekUc8iYGRKWhP5+HLd9i
x4224jW9iI088COzOTAEbv4itGmquO7E11amqn/oiDUsEi5O2BHrqHWcpw18fDKG
hlbktyd1F6oIYEikpqKFVj2D+jvayNYgmGQcXWMRv/NSZ3U+oHQwoRDu425l6pkP
Omt2AnDYKrKKHMgKXjxC07YlocLtNmQxqxYVHv4PAf6xav0A7ZfoDpLiNggCCtLa
/2cE6OiQsrbIV//GSGT2HNfNp/oEilKzHhouGyTXCDXsnG7tB1HnC+fIt7ebofOF
3G/Z3XY4cndMklzcvOpFeMHFQ0ptvei+NZm94Gk8G1fPq9M30wJypSMVsiQdtr0m
0z3kspcV8M0llNFi129qIj7dL0VF4sCM95sQwysSlVy/uHe6AanyD2jepMI8XYhr
XCD3hVvU+oHVbCM4MAK/HVEmnYj8VpdkpBS7wVkocFgnCg1zH+c8Q6H0AehTPJNe
k+Pl6P4BUjVe0ENomeKyPHZ7iUD1bh6RyiqnudhdfgY6mb427LVJM2YRQFms7A6r
MPJpP2cNEx2/L68ZeeXIQv7vvPiSjO52q93WU36fb4NiFEu5OMtdfk06RFtfr3N5
zWIJD5r3juVt0C0EZfmY7a14IXlVtHuBN64N66Bqf3ll2dlN2rL9P1mzrKdeuPFG
W87QTIXPrJkZiWvB5FKjm5otCTzxcyAHPmM4h66+bUxNV2bIEcIX62RGecN3Qxpk
jvFW4tkMc5rQ9RE7BPeeqhbv7FNHkHSOWOE9cQLe6+j2YxyhIuPcvaCQfdA2EKJ1
iG0R2dqLwLJLcFK7fSHjffi5ZR/n85zbgJukKyTd4vhPs6ZIROkShcfUAVwwIC6c
4zdpZhxBm9tDbbvVnS8m8xdTfKomJr+spntHxqzBj0IfDRaaV1YXZHdcSUu82sme
C+DJHbA4LpLyN4w8jcbJZJ2MJx+6Sm/S4bpirVndN/WEOmYOzR19ymriNsI5WI4u
sdnbmZx9LTZAqkg9faD7KWVuqKKdvqyvoH92N5ypuWhFJXiII427dTNY7DZqA7Pc
p4micTF2JWhyduJ46FTaBC/HZG8cKTSxc7jjVDGaHZhwii+Nfko4avKLbjE4vFim
KTqco6fVRT8veE8/0gEjc2WGUGQnHx93cvaSMlxQ+UT7T6unqX6tAwdorMbWEqjO
Gc094qYKZuwUbneaWc59M6qtjJoSS5ZYsOpyfQ+hx59iiVskNb5qfbtJi0OpKWni
yKuofonaqN6czKhIhm9XD65rvSPuV/bNp5sJ3YB79h5eAAL9UCdmG1MyzA0QWyf3
mSAqE8diga4SZz0EdWw40OPIU2+6NtFsaInUqjZ+GADXSDuPSYa4cpbqjJAFpHGD
KqdbJCM2urICJT1fL42DCpn2TBQjnY//j53DCJfPykNMn4C9T38vc1rSKFOzTjSU
lyu8MGkt9FOLsJA23t4hvTAoiMd/6W5eJF7EnBTahxPj25I7Ge4wLxMpZ07/E+Ui
fLEt4iE675wl2VIfv+JgN0X8C1c+kvRVjgxfAxNjGkvuCu4BpcvkAYTYj3JGMBj0
BfXXgqT6R+oT4exZ9Ny1mOZG3rxpLtGmPNEGrYivq7DPpHu9jMuEUQ51eO80gqew
gihdCG4MwinCg10Y0tppmp9VXy2p6DTB/PpsZG0h3yFXx2cgkOy+dITZSt2noLsY
U4ZoUvYfXexQuk/x0hOny0vVh0PGuYA9M0NvOEaWKJBj/kpm8ZKSG1FUf0D0JyMo
DqMlDm8OXW4lAfPP5OIqqw4cUKTb0OpfBmR0G+5aJB146U//EyCET/mJLB1GXTTJ
cODGxOUpBrf14tnnp+329RRcA2XPJsVK2DypQ4H4HLkwIkowdUE9OVIA4uQLzQhS
KCTK6sm+6sx/o+RcIzbXH+esasGPjo2534aHiUzy2ieNJ881J0o3/IODYWYI+5yP
b7VpKAEeEWWrxtIrKsA3FuTTnYxZ4Nm8FbjcWW+eN+ThHN+YNIPkaFTo3lTF5FHl
Acv0IpPt7fjajt1/aQeNp33isPFdkBCQvsQZ5BP6Iec8EsVcVoD7txAsxEnF3+bJ
RvBVTi03bjyebS3MNPEgBrnOnAbgx6TVqlQWk9ggmdL53ftM8XGmeNh3LaBz1395
NBbew2B3CiIIG0olAyPe1nAV0707uVtcOMUTODxnoLaymBjzWP3uYQL5BRZ2Sr+3
tyJ/6mk/+qCFLAVLJyryKAL9BYmYKbHv+wd0obCwcCbZhwy1QECrJUWjFKQkvxYx
tHabG9zpz9HYXIBUaeSF1zKeTaPEMfQO6hNMuTkp4J4K9wjUijBUwrALXjwlGgfN
zTFMqvWigyyoyQOw/m4sUi5zyBpMAWky5HGxzuhJBLQuKI6a4IWgnNuNpkqLrcBB
eihK/b24TDNO06MMFzB65jRVL9JzpgUu9VjuowegDSItTgn2erjWnL9QKmsK4dp2
3VN2+GBWEwAbxWwbH+Rmms2APnIAdVRKfUMV10Ymue+wKoLsXgZ+VZ/D/fJkGA1a
j5FHNs2+3ArfZf1K8VlBWZzOYjTbukV9bU8f5g6yGHd8tGylVmUuo4oTHbG7PRKo
JZ+/vVgKuKoLat5NZEISFtrcCJhADzJdy308Lzl0Bu7AYjTdE72fQaGwv/hkhD3f
6irdq0OcsAtWCZoGvvpxWmUHIDttKD8ol9+v8v9EIp/sEu51hkw9+SmWTgmsPW/o
63nF1oBCnG0Pevbm4dYC1ZDXqBUAjwmWmFT1B4AH8bgZ92+Oreo8otGybJw+GLn2
xK0LngX3IwyNp5LaJu5NEHYrotv+cs7RQB7vKLvfZuNpuBQR44hNBw5nv8zodmlo
AjB8lUm+O4WQ6xFTkUZvJ1a7g3U2N6/Oi+V/BTq9WHBnFe8+C3rq7zJlLiPGs1wh
G9xIIWNhdchNBKYf3qOwv4LSX1+BvTLTwHx9Dk4j9FSTlOrzlCWscw3qfm5LKeBJ
j5A7FqJmyt1qpN/DWI9e+tDQi8R/RcLLf5hd5j/OEonKyOuMTiAkBCD2IVTuwe+l
rVBA2prEGQPj2F0wS5oE4uc0yUlUFETrsGcQovqmEZTdG+XtGQHnkz8uBQsJRItS
EhCQU+4XZ0/Ss5nR2AWbHxXFAEnE/In9yiFQRUijosKjuOXql8mA2DEQkicJh3Eu
f1Z+L3FZ8+PaqZ4yY5NZ1vzliSNe/sLdzP4xHWlf1UIcMquYHltjZn2JYPfXm1fC
hihE8LDnZc7OPbTx5y+3JY7DrYX3iZuDrPVLpm8qLEbMSPQtCuSK4oIUUQFSDVVk
8vcutFKg5yQOaJpsJ4fxs80szjsfQ9J4At+w7vlsfixonkg6ns/eJV79E2v/qJSR
DRe428V5pjA+8vLv+pEeMN+By/F1v7u2RJPpnnbdNx1d67LwscKEsKBxAHCLQgpk
+qjXmKiI7zEJSkm5GICIqmquPNE+wDnEhSqpXgKyBn7fK5TG6YwH6HTDF0wob1LH
o4FcYfj7G1OBl2fbPUM2QVHleX6p3Hj/D+moeIcqF8CXbGZH4ehGpGoDGjf5uTK8
mdYsam9BuYSPl7XaRTUpj4v4WhwO5OeZq2DWvhwYFl5TItgfzNRgeosd3LYf3U3p
uKfBG4x5eOL+q+IjIjvmABXxESjwgT8r/PRkwF5ngKhQHpcvRmUtrNljLxLWgD/a
MNjCG4AQSvKUAa9P7sCRmqLxEAOCiKNpzovA782tzeommbaoOmyYG9g8IRN4wsvz
q5DF3NjxUhrF+hAH98CueztQXi2xNe9fWSzyi2CFktp42iS3cqk+4fm2spcbZ0FB
BUQsUJ8qciEJbOfSmfbe8J0RbVXyvglw2riEyivIpZ9dunaVRud93wU+p5ZecqQ/
GTMKqCwxw3FkhgGtmUOSHRO7PAxQKWzZrgptvN9PozOtNKv8gntCeDUK5h9F1Fli
ODODF5Th5BmcesaTJHp8BA9y8S2WZd54aR9EFuQZfNPpL6ssxlV4Sf8zUTqaUk9I
v0DD87IMg2gAoIlsSjlg5irN8SwWCye1Z5phwMZhkYlYEc+4Kz0l1hbDwPdo/lhx
nMySovbbMfBfXcAc677Gnbg+awU4QQr4bqXVyth1//pUO+xYiR/fRDgYhD0y0Bdf
TVmE3CIqlDwNV9sMjTST+Kw9F6zjzp5Q9I8Up/Y5RDX+GTs6yhQdCSSHpl2M8mNW
CwboI1YxZZBrIdAgl5Ws93CZlk+SNA411qn+LCBss8ZM5IxJvalZZsh1xdgvdYki
ApxkRMiJ5ijxin6RbQsY/BFE643ksulAfNrqYyKkpJpEhLjLBKzozVgjTL6i/Ee2
fazms5hkV+n2v5oU1zOiLXpH7sF0YmJq4a0iEngjO992KPL9m6pO+hftoe7g7UWI
eaJn29u0lyv2lDw9foAlBFt0YihkWcSzKmhc56IbNe9YE5k01HYqmb4QmbD3zA67
ZmMG22Ob7vbEEz+Gj0/Llbr5vRqqQPMB3ZTK5s0LWnjQvTJWq7G1fiTHgDCPzaVj
O3KYvoaT0CWq8Kjw5UTiEnDS+cwAbeWdL3XVHM5k1K00atzw24sEMwfWpvzAbhWS
MP57nFFG3M0sfdrSvxODuCCQXxD9EEYCW5DtVUj5A0AhLSL53crgj3Bp68Rvuitk
ftZGUVzdSW9D2v8j79rHHzi2hv/iIUiMeyUsh4dfygQ2rTyHhUd/JiRdiguVdRuv
0B1qsa9t7niowT8iYNIYk/z4t1nPyYXzk3+DIJ6u3uqdKvQjpicbAtYRuUoN5HCM
m+IyTyFG7r5RTW1bDXWoi8TSKnAGrWtqNs8RW9b8VYNcXyP3DQT42scFQ6fRbAo5
ba7owAD19hN0iadESvwnVB3YciQGTVTKKYKetcuQwBXGVqGIBg1wbHxLL3gjaP9w
4FV0i1ARCelC89imZdc7DFIK5yXhkIw1VX8h01m95EReEDrByFgT0VALxMhp/AoR
m/hlXeY0RRyT/Wfs8oO2ob8WwUVfW6tmWNv/xBqEepicFkcOjLPQ1ljWlXkw87sI
cBgV10LuOKLncUdYAw0thLDKDwkw06pr3Ds/znyW2N07fI/MQwh3lypCY3g9hxOe
Ux/9e7B9MdFwX+FNJ8q8wqrEdViej+J4QuXpr/xAmPyRGSN9kB1OtGZvH61Wmtvw
nt7JqOBrX1awgaBNjA0S+wfby5ECIRVidrOtHzgQsZzDc4Z0FN1m7h3TC1vuZFfs
o9/dtCxhXjxS9RMNYAGH5Pub6I695mdbBptZfiSy6XfppByDu9ULrf5NfMDljRor
vZAU48WfyHlBRV9eJoDc1t+Lmw+Lk+lUsCjH2FQU/X9Dw57gKNvwvo7NiszUXpMN
2DJXFKGwzW+MCV60LrarBxwlqN9P0khvblreHXxPe9slfRIcj/RTnF/D7ElReS6+
EfHQjSDGiMwuREMXM1DGE60CC/h+s/9LIDaNd/qMMrU0T527W9D6tKCuSeSVSmtw
/ENpaZUSAzidNNTpLrq2w6MdoMRkOor14tHmb6TG08DY/Pp6q35WjDFUabJ3ztbx
g4gcAJAmnbTIOxm7fB+Z0ZoNRssFa/FjVkgZPoAFOjRCmJU5DGGPJpcnJrQcvhv8
GQc5tlVnr/AqUDG54SH/4ArTSjvP+OrqZL0IPwSNQtz0sIBWsIiA30cgX4gL8w3Q
AsTEky7B377aPjYkoFNMhsqP0l7+H9kxCEZD+JHW3lQ2CBLn+jKOOGswGboVIaE6
rkj6p4g/jRZYdmQ4XtEo9asaMILEJ+VTVpalooDTQ/ngJiIj8/xmbjps3X2ciS5X
Qi7XZbU7gTpOnUwXYK73fLen/JzHeDbW9en6tqHf9OWRjvK+4qNNl6uhIchNAaIa
kaZXf+bN/U9G1tJRopMY2pXNK9/nKBNgsdMQAuMc+sdqchBApr3NSeqcg/zUJeMe
kUfizfkr0bTDtriQ8vgST3W25rUh+sch1VRV+kzAY6YucVpMiuLS9RyxYwK1zBaM
1cFYh83JTUn1eznRL8HlMqKFPo+z5IdCvNS9BBmr/RRMs0vvS+2xCxjaOaDDjyvd
xIK8XC8djqOd80SeznOHIn6yvtOvGH/7sutryUtEaO3u/YAWxskYTfNed4FGawtF
H0dJr155JWtLIky9QAwTsT23YH69CtpFXw7WO6VIMJYmLOmRtI6H0HqS7SIJl0sz
5qI1aMtEeZzVOm1MjcxR006VPJ8fX6rVI6XeNE/vBUTc2U7ugFjUZFyf8D/KJn8x
xDz9Dy4+CRAS7lAmjHPgl3Kp26iTPJrivyV7O6dVmkhJiWTCWSeFTdMuM9F/lcA4
kmXKcCC30mzmv8m+udUm2WBgBmaCm1wFRgpPcrfPeSmusZYlUYLytM7fg4rvo9UO
q07As9b/EJrkyPrkkO+gaEzV6Cq087iCMmmfw6cVfDRTKnacCXXKmtkw832CI1jM
h4neytjZ0ARbUtgs2GihlQTqv3PXx7BO/tZKmvodwuMOTlYzWF0dzwBrl1vA42W7
qoMDqNmo3tMjPTbOnf93i0cN6W90W9K9DyApl2YlM4U9xZ45ey3zFvmCrZG7jhwj
Vugm3UqpdaRlAQLtwjQ2LLy+uImpAMFS/kVqtFNlFLl16Z8Fttn4mtE7TTZnAwPh
j/BMYFMJfTtXcSFJ+nhpFsjUIuMn2XAVFc8HUmdv1dW+mPoXL5rg5/TTnKma2Bzn
1tXB4CbqxBGaNIVXyZDdj28kX3cG3afvrwUD0bDUFeRmk1LuNTslBjZfuszjTfwy
jiQcIptuUF8T/R0KvToi4FrGa1Fe0DQp/5Naf0eNaaf1zAGHjW5hkwKVnPPcUFlt
HLnXnNyQjW1X4skzJY00KDIQYjzEyzo8np5EgLjHIFQW3Bq6fIJ4SpUjxxRNE4Mh
4o981fhOASvMsphuWIfbiU+cfEzw1AYWLxVDLheEm9P3vzNmLhtW1rekwoBOTgBB
lyNK/1SCMxaKZkJxE/SQBfN3GBTGiN5CKcCmx4WZ5yS2i0t1nQ3QmRMIapZYbf5z
KBfLp3EEXMTFKTd/BtrRRn7+GMqE2RhXUbaYSJS0zsNpcsbBhik8+QBf86TkvFzC
6hl4aWPSrqeekxLgyof4Oa+v8CZZFFEVFicK5uyYxHOEWbXNxahot8arMJBGGJPE
kK2Lb2hXigJMZJowgXAAIa7ZenH8fKq+SU4mY49nmJy5io85EFLMHJeawsAdYY1Q
h6T7m56xXH0rqfwWAHVXL+TaoDjtnX6WaIxpIHShQwbHVxjOC4ydUjSZRni22PSA
fIwFaqHBKR44QPTlFmRKGQSV0e5+P3ZFcThiE9aVwRxi23Zf0tT53+0A+rgEodeo
4l/DKNolEKnMF5cLr9GoPoGi/xj1+P/ZfTP11zYmdzat7En5S92a7RYr/lpViRbV
HM9p0Pr+29cR342CGH0asUSaFssa5iGv/+zZOSSF1xmjKnO0irMfkPVHmGfdPqFk
3C2SYDthT0FwBtiVJyDGmmpsZUqBD/oSOPFwNUBgQVvG4rViI3z6OUGRg4aaNa7F
Y+nDFZCWAZJ+E09j31e7oEmek4i5G0kJD+fnn3bzcNUOCVmhx45g4ltGXJJ9gerQ
Q+TXBmlcLf3YXA6Y3FeJWKfxpFwyjvqcr3euMw4vm0ROMBN3usEGMk9vUm8+i8BP
FHt043Xap5iapWIlT7RX3OYSh1XfjIuWnTGHPR7KiBrzmN64rdgfoSYhdV3LI1g2
Y83lO73xUERhMJt35raX2JH0xAflnsmWCYnIGciNl+t8fVcIwZyq1amhJMFi8xdZ
xIMAM9jruWuDoMnDxcioI/RtGX16zN0s/oRAIzTqCRylwPcItuxtLAAKPo+9AHsT
45VCaO3G1QLD7zGJqVC7s744LHnjwa8Usk0BRYsLgGOJPe1ASTtkV6Tu8nEwLnif
+mBVdkKGLlV1gBDO/TSiNP80h190HDYKe2nBGxyz5ihEa1TP3g0vyBUf901oh048
ZR31I8ihzR/QSiuzoSrNYGTBnWqsferbY6rgVyrn1X1kZx3X8ZtpczqskTrLJ4nD
MvxIo9mNWkOGS/i31EOSf6OD9n9+nuaassUyggiJ3sSMqLUfN1fKazGKmFz5gd1i
Xeisco9MgSD7lO3QMBWVDtFMlJJUbSkxraDWzDI97BWGF1Ycw4ntdt3PN0Uj3HKw
IH2p20YrdjDBV/UakimpdWUmLDx/Re1oQBqzgS5zE6XMLM5JLCRlLfopMFatzLks
cyJokLv9gLDWtA6TudBOAPumxHc8FBthTLatztXvdrKvPS8tx0llUnMf5sxNdxZn
a87ftkToxNUq9Sdt/cLmZY4fD3rolBSQz8dcEhSs0vQOnG7q71LIZowk1UD4W4zh
ZpPwDDZcweTnM1ukRrWpRwwrXI8aaGUV9c4cWEc1uLpC0jWtEzVEveAOh74wiQSA
UAFpVE5K73h++Ddxt4CTq9kGnWE19+TeJgeQd2qrRhbD4HsYRAnsPS6Hdlx6OYhK
K/nNHsA9P7Jziq8mIdUOs7GWnBN9dQ+LPq1lX6zruuLQtWVmP7JSk5HHo4xiEoow
BPoxuhzfODko85992G7lfzmHFWCiOqVHewA2M9qabqTkgqz8faG1LGSK40I3Fn+c
lZAG8CoBToyuzsJzcDsJRQZDBpt4pygKxizP5F+d4XRciU5dwf0Oz0oxEMua9odv
fT47Q1NXKuCRtKzuuW3+LL7P/ZubbASYRFM9kb538PI51vvTN1E9Zi8+7zTeRGcr
1ulXbRzynFsd9a7HTf3peZu+8ohw/JUnrGwZTX4eBCH3IWO7JbEXkeuLDFHkerG1
pczK59ACM29SqxcR7T63yEPWoPArfFe/dIe6wgIrZabgLFqd7Xw8BXSchpqrrhPT
H0+SKSwx2XaZl3qCmwBASC9ozjOqNhZsX6Vc6Q2qo/eI+k02a50kC9bUxw5Ilg2S
b1qjNyoAnEvga1qSkani6KCRiS0mR2zxTPT3Qe3rSDnGjufOPh/C28p0iUUcbTkN
+U6j6EawLGrgrvb+tFlN6UNkBgAVM4+d8zSUmhxso/uqVE0qL/dUAdKHqjbasBDf
gVRAuaMTqnb/bkdTA6PcFqFalI4IouyPm4CkFoNxXcf3GEnhfuFgF95oZsyc2Tcn
RtDIFVUbBBt8Uf+IxYR1DkYK5Hb5+fPVnCwb+4pG0S36SIOIJxkDy1N+6RyENs08
kY90vfjddykSgY/Qc4iw4nQYKvUyweBWXtN27rId0YQaayMpXIxkFauqTErt+N7q
GLL78HqEwVk/5IwyetFuRAHlZgCsEbTVYeCnvRyQMo31g/3SEQvyooR6xSbTkKpl
4NOXGnm53TjoAaEJyPZxEi+BMnyJ7TZR2rqoAA6IPT7jk3LlZJ22NqleNQscbjkv
XyIEq1wOaJUMhAZYzdPOWnL14p3FipoGuzKvOdwJwdz1ayh4USgS/qL3L30xMzd3
RZeMTHmoikWme8ZdUhhoAdSq+Mo/AZn5fR2A+7olkq41AyvzlGoYM6FoWWnYiumZ
RvFWF6bgobZRlSwMnKC48P9BCYjweOXnzxUqNuSvIam6UOU9PqFjwY09f4L84Cfk
ECLnZKJJYkwjyz36/FUALJ8Hvs+q308/Y/Vko9VP66paXW9jszju/7JJwl99quKA
7oMrbNAmgkVj8fpovZztyvBvXTZbRqb5HY+JfBZ4RPWyyoTrWYW/Lnt33Dhi8igT
KIBLBHDozQFNbVtaBpSQs/ip6PKYRV9UMWxG/Sfb8cTRFIscw1yWA2AxVXEr2VAA
IgJv7Hzo8W4UenlPxWOUo3d0MGLtl6F1MR8Xzh+OF1RtQ4yH2GOcvVO0M/a6y+Yb
I7x3s/huiIKthvI60l14Lf0wFy3tAIO8sIi6VOYRbXwhdYT8WV8vm9OComcugSqC
OyVE77jkfufSIAYjpRJZU/XXet0P1JrQVoHmCnMv2gghD9STR/zaEqV7/E8rXfu0
8gZOn3SzKEiUXkkH7/z+pvVWXVnewarLCfen+aBfbqXyhLsQti5LFVvsoJMN8uQA
ZOV2ySlqIgjNHLwxltW0942XWV4Vs95BzuuhcpqjC5eES5ydlMPlwGF4TaiRlO3x
X1Ux81B6yeZBCoKWlx5KxVo177WzA8NdCUee+cHHXoNjTBjPY96BCwZW2GPPhcIt
BOhCYQKQ7SWWfeqz00xijTyh6wVNF9FZwa8GaGRfFj1kFKAdGNIsZpY23diCmKDg
/xgr7dMuABvICJv77PjmsybYN+MFZAv3/JrDB5GcP7yGSFQpQ3oiF3zdvdTndiNt
eu3WbPeIqfAaZlYYrQqObl9sU2xrEMM9aFPpZoUScwfz+PuCAiXAcIw1UHRjdSVm
ZEfQKpWbVRj1pKDi/IQRqiDdui804hIVi0yLS30IuNnDsjNDTsskG2r3IdwrO5Wi
TboXF91ilSRusKKNzKjZ2stAsUQ7a93LW/fKpQCVh5KSlxoKEeWmYwebil9bwSfA
lN6EkDNlt4ftgjO7Fh6gz2sP6SFZWUT8EeSkKll5A5tKEelbjnS7v3djfAGf0qfo
Hq/OHgGWwx2Kq45JgQhToeCc6qtzxJYgMyDw7OU7uElKNK+gaWzpChIFUOyyWKOA
SEfk0FuTqo6ZqjjeiQSQmWBk03BRO5owPHywRXeCe/DonEETSsxeWljIspAyQOxa
6GMlhmJqZqGDhYV054w8veMT3YNyqc6fubbfG56EEwn9N9TrPzlXmQxJnxY5wUDZ
LHLIfO77vkLXlqdAPTyJn+/5dYC02cIw26wRZYQ+B5Nct5pw0L4iJbKdT7guMfg2
h8ywH3ud8zNXCsI0XzRc1np07n2zBaUnuTL0etwQUrU5SBp3GJgFMmklDS5dw4PQ
DPxE0Gyr6M4/Er23xzwSPxbEeA34xUKLQkPex6WaKG3lNfluC3jqKLGMYln5Y96Z
BkR7ea+V2o+8/QXw5cZTlmUHPVzUyQP+QCeNZZMJt4+EjMmqd8idBM8uyR1cMQl7
zU6ymvX5YAPPlDtv/xff2wosW9heYZL4hvXRIYyeK5QAE2zVsCMgSZTPKA+Raw/d
H18GK3/1aUcF7TiVJBbEnHN3S/ALu82D0+Y3xj3NCf9b/zJqi9cP7WnpnR2UPqsO
sBcYopqIrMy1iISqtjXvkSEQgOnYSmb8/KcX4J7eJyeJzk9jS6T2sT89ZPeP5Pjn
jghl9AeQj99CyawhkWuy07xdUxVx561sUfh96LYduZKjiJjz4kLI6j74TqZ/3q0C
LY8Fdu+ByQnvRD3TKs1X9LrjWrLKl3Ja1YV8Dag9tjSWRqvv+Eetj7tQVv/wHtSa
DYV/KUX/DcnppBGMGJM8XAijQ2VVSnd0xeK0DMcXNO8KNjkOgz38Scv/sVsZglD5
VmYrg1YXrsY5qoa4+YeJK8MxbpcsHvWLMSntfOGjY0XH9yb3eU/5fdtRhm+WCsnl
MS8feeR6pwf0smgBLBgy27/s5+OvE/AB0q2DJCtoOIG+sppvbEzaWiIfqSmbBJpa
/CiZCMz97ctfgAyGAx9yOkSSbfgzxmp1drc0bVDazIH+2TUn7JXtwXFxpTYr9kkP
ib1uYQPP0cFsuriODOo/9QDAJ5MOil7gGMYzJ53M+wL3PRMk0kGF17JoqQm/mH0p
mc5wHpWXiA6kgYNXpH7gSFYpvfNuGcbs3JnOM0g6qUFwQHteuvUBNiXhVjqHk5hU
qLwutYwCVjpzBbGturDcqGUCTdA70w3+VNv8TiBFLO04CXYdd2j4HTGzSaTT1a29
igyGxArQlkZ2ZxvJsrhgl7lL+HlZ6sVNIGqsYEn4o4plR0PvsUZraapRHqA9QCVu
OKZXCpLzW52x2o0KsP9bKngyuB9Rgmr8pyBSeWmz5MWwTLetOGqBGiHtEgNm4glt
qcm4aYvW204ttEMaHVgbOnitigmTIKHyphz8V7ZxS2hAwu0DR0wimFvGi30vhBv+
y8EhtCkWO2j+UJ7bO3Y1hbETcH35YJx0wk0ubT1npVuIk9NRpHCv0Xgp7I5ME8t1
EnJuWvMu/BT410hhE95Yb6MWymNgSvl5atWVLN6w86DuQMu5Fn9ZwH9vGkWPOiZj
BdmrSaPz/D6TgXRqCklpDkO+Aj5y3cf4yj/R3EkgtI+bAV3uWTS85uAwPgjQReC3
0ZsALYDOowTZmY+/7w3cyr2tmrb8+oIQ1rGvT5ig/wjbs60Dz6HfW1zY9hO+puhw
7gUsjOGpNKjJFXhgSe4q/9Bw2gppVoFJp67arR3P/XG1rIbbgb3tyFl6geASWvW4
4oxu7vgkTbpvIKtiZTa3siRyqZ9vs2JXF90+gv+cPf06JI84gDecsxtzil/D8UAH
ZamwXKoAju/fw5R695Ut20mRCioo9jJtjMR1hBM+KC9uYvcAaLDh5+DUFLMGclbn
U+DDjdY1RGmPWjNvPL6SUFTFP9a+mgndaB/B8sH8hzlnZDJhHHYpVw8XV7KYcJFd
2O0sqvg8azGTeB2RJ0TiKDFRIHd90prl3Mtiu98XjI5blwvNPmdB0qGpCZ9M/Yko
W+Ttcg3CsMYOAPJAHm24osCNlJpQM6lYbKC84l3wMU/Fk2z5ZqS+Bs/20E2lWoIZ
I5YMs6nj/q+fn39U2feNKj3CCYRbojc/MqEpq5c0ot5w4yKittA2Sfr1BM/4LX68
hFHz0wIwX0MjpES5Xwia/i5k+h1NTP2X3672h9jF0FVnev1JCDdc52FGSspEmsG5
FiyDHoCTs1goEPm1Yoy7Z2zelBs3s73Pbk1+WLycpL0rLDLnX2DFVjFFs2eM044j
PzTTOj4dAg5dqAdIRB2jEsWeL0UcKdZSwnfSB3sLfsUOJQqzZi2ZvRSSLj+ZZ9yg
XUnx3BrmBUr6tq2ylavGWdEg3nFtFHaUVchGYTH2PnyPl24fzz10T+lJVGpb8eQK
h56oHG88+fQHWiISndnfWS8hh2qmYf/0muPcNaKq0vV2mMOq3g/DxiSHabnEwLmi
hWHUEH8nSjhlNh0aRoMQq390/B7GCp3+Xk5Wh+kdpxAjtQA56BWj+5FYBMEsk+Yn
1ZEnPMWqPdfRpRbYMCEdXMfpBOP03qV0/QH9xYe0s2oSLUymBiJQIzp4a6RAjW+P
FNL0hA4JnDKEEyct3WVdykzh5E2xs4tukAvrRUARrBh6HNTcJ5w5H07fzby8ONmd
Dn0fu51ns8Ipr2224kZipWhEQEu3cwc12h8lpRCcwRT8kKWmBkquJTUmIrPBbQQZ
MBrBGH36BO6fW1/vo2zg4paHRxXRzSQ5cZqMHlglpEbbzIe3S4H1z9+iq5J7ebo4
tUECU8QzcQBt/ci38jr9RfAcQjf1Mz6uhjuJ4eXVAhrquMEs5CY8rd6MVVc8mQVO
KAM3mqdfpLtxV6v9bmB9xDlZgDQpzQBUqzPlmrA6Jzt3XkUFYbf1oZ0cwcisasN9
z3OPQ9kalhwWAfClNmb9HPyG3mQRzTgbgPHWaSdNbAJzpTW6sgjeZUTVEbt1+HL2
v76uLUDKxaRafQIZsuYjxsnn+Rl0VjgXH2PNPLKkBRzt9pBgMGkeCzijLDVJrNkC
BKs8eRud6KRIhjipuvDDi7Dg7FRotjvOx/be0OlTQg5KgPP4ybp8mHT8rbrUvbOF
3PH9GNd8sBUEneWxihdrwnX6NoAtF0NrDuvjCGtPxTDN/cx4cyB3kZBtPD/6ra2D
O3q1eun7B7iuzAGeHHdAg9hY28lF6AvvhdriMYVGDnUDedXr26lslJXR6++zibgc
Ng3th6T6prYY2Wsw/R3enkM44k6FmiJ9GS0SKQemS9KarvnenSPA/sCvDPswUCrw
m39kSqYGQBiRbuEAD3T5GVfcJdoZ8Pp4ON0PvEZDCblJrlynULpw63RPwjNgGa4h
56bmpiII25AEcXjWKOy59FYp0LLkhdiWEZOuGHsI0aeXSTJUp47sFQ1X87YFQMpR
CA+YdkqwveDC5sQZn2YUyw0yVgXNdccnShHhqPAFkqEawqnOzwh0qYWE6r/e7ka+
LApYdA8hUI/h+IRn5n9XMGjCmiCUmxjHGGPdgr/n7btOKtaXINbz8su1abT/S7eD
exorG8CYDiw6gyraJcjqNRycI0+j69dKEwpeGzpFEy9+nHAEHhLIW1l3XWrtUmVP
/vsTU1FT3728TdrWtkOP80Xi8Dp7QLqOhA9WCU3aAhxfIyhhiYPQ6PfNrUizklXF
vNWLCZSxq492XnvT4frYPjUNgqQbKmD6zKNqG4498780EIanytDa3L4UnRtCsCy+
UnD2tCiXhrw+S/R/lQep+RwDtKJmlUXwMqhAIVpL0KhG3tJS9mgjwFtDETiG+ks1
tPKDNJdv930Y8p2qQOzRrpAxrz5IPKUKYl62eRacJZj3npiR2J+7nK6aegg6jBE9
yA4e19MfgGG+YZclZPkaS1ENf4zWeQyOwYJZHzkByvfyUcbxs48ukk9xgYel/rYW
H2Sd/Pg81+C79VWiJY0x4TtRugqNOr1IlIkHlSATSP/9nwy9jIUkmz7CrAOrvFrz
c9eWh4jKvYBuXcuGDRxoLMCZ65nvR9Rsn9nQs+dlylmfeQT7MCmQpSFsF1aJUvWs
/MbohDtcoRyNaXR+K3fEPgceDozvVcDn2b+3BomN/QKn05gCEJ6WeXRz98bJPnm7
QOJXCQQuvjhHpCn9ec+a/a6tpT07ioLxGAQ8/XSJ2OvoHLBn4OgSwwx9CCyMozZ4
bIAOxxuuAh9hQEmuLpnONHF/bjn1rkSSaie5aCezrYbD4pWhE1Kmj0/+wDpC8Mts
noPk0/DTCmxMPh3Keu45P4CFqxBgIyCYrgQFEgxJUQJkTH4W2CL9Dcg0CS51iQ/n
LAtoRcST71fm2gepZah2/CXYjYyRZ0CA5bPw0JU/UhAFTXzpUY0kbu4lKM/w7I/m
/+qysypJvIxNzojbxEcawdJEnCBaZyuqcUcbQnZ0rIVfq+klEnjsVp1ybNKuVUZ1
2W4QE6Ui0U08fW/hdnViMFxl4ps2zQ0h56HJ3+9eFGUZvs+EfjEoFS3oNabH52T5
cBgu78kK+oFudGGKhLEcWm/iu0pvL5Hekiss12dtJpdjCqORHF4u5n4M0tdur1aR
O2lnu6mu9gr9sVAJ104B+SiamUuaqzuGT2hhUKO+tuw4/SSuys3En9RFC1c23yPj
bLDuQi/S0ZjNmJBX0Fi5Jm7vOGbfFW4gaaktcj8SrDcJD+mc1Xj4MBg6MNI3vvIW
uVMwqHKVqukwLZE7XxaxmnM3+k0eoRTAdfl/8DosVpyy4u67nL+p8rTSoNo3v43G
z9urAmMZe5Yb1S+ilHh92UKwdp1gflGRgQL9dIcLva94O2RZD00sdctE9shjev8D
zxorgdFwjHiBNsKWzaOGC+TcLjnbeM3fyBI7mIqbp8xq1ZXljZIpqYYLzSOfeHOt
vuiQ6vx/iNuhbgBPFaCoiPnP7EMWQyIhH2Yrh1TWsSnx+KGQky78/WZSeYTZzNul
50FF4h0NyXZB9I8gHU4isgnAIriqjpjNvjKkNz2a5i1y7ZJkDnptjTpGUn1T61WG
VOaMcclnJupFoj0hjg1zm7p5FfrJhGsneOkQHwO4hu8oAgcvu+SJI9m6tmXj2mrP
zYzfAaQtRxV7QpjdShnNvgkojh0WdKbtG6vT59bz2UkEMtOvSglKPOfPHwdNLx63
mr9kKkum8JSMM8c0bN4ldBAJukWpKnKVdQI1gc3oaJf6pCWAKxwxQ42fiiBzIKpW
7TnvU1UiqdAf15096s3/eADn5cKhq4IIZTEurDuOlAgs/E3UdNWPG6YEuXZs2wrN
r8QtsTHdNIKGVGKM/GeXmH6vN/OiFV11rMSJRSpZg2petue75WyZUjq9osPr6Xrl
8SGdTI9QlugjjJOENBU66CJtgTUTw16CIZ0UwQb4Ssc8vTLbKFu32gwQTtSkC8VZ
1E0Z8RiXakLvlA+HIZHmb2mvDuPQTQlaxSqE5d28fGBkbESIY772eLXpBltbZEd7
g/Nzl7red5jncsammS+gWDxC8BvnBkkSmo3lNwWItuvRnU/y69cqS81syMTxopdu
Xh2ba45EqKxmWOFbIvBqm/wTau/4keUBU0lmcDk0ZvSvJVn1Qq6+MmJBkjs1W6jw
oVKFhOxvsvCrBI3G3uh6LgHI7D8PMutDNdci85WBQQZYjl7m+t2PvU3AfBzz3BwI
O2bVt9klPfnNDyeqj22HcrrAV9fErdGncw1vIQOQK/n1zSEf7WTBTMpQHE3WJj0c
mFV3/Ib5y6IoSz20KEHsa3ISbExycDxp4ImtYnykbdVBOJJgJOWl+MFFIVPH2Agn
EwYsBceU0baOvQNfnzeWfrKFZRhTVcEXFLdBVeFFk7c651qSS0y/Y6O4Dm/GJRHf
ZKk3YKoKNwrYTYreVExpRwfGUUtAZ75Q3djGza0pTb0zZWeFYLJ6LQX1MZZg4sv6
ZFJed4ZHSTOI7zoTAkEH0n6771QbTvyEgQXLxJZbh5+HMKy+Py4Jt2YRuXu30OYL
+Sd1BvNUuF+kfZVu/UNFz74U5RrDz6nH8p8V6Y0ltanxoN9mQQpWXCDkt8BpYmfK
kkFkIiXIGxdNzr7fAnP9h08lv8k5XrpmGQLlg9WZbx4vcASLzZYIXi+bavJ1lnok
sIPTeQbJirZFscfnqKSieseoFKIf9zsTQf0BIhSEhsQW0MVPql5l0wcKc2GUl51E
OTfB9RvIqrW/Aq/dNi4dkCLpjERSnsXQktaB2Tg6NbMP/P1ERLamJTFKfO2S/RsP
vxO+lebrAFfu2gJ0gPwPQmMdI4m3PeFTnhiRY+Cnzv9BkodABJYdgzjTDGtl9yUA
DIF9tUMZoDAHIMaGm/uksoPxduCoJBNGGRoE7js5rqimc7dPXIRGBR6drPuixKYm
7x/nnuZI55rkmQO2+bp+UMnJkN4RlqIsOCCLB64y3HrRNxGQxpgNJL3ToP48fQnP
Oghb4Gpr0Qm/qIc/zAhErokIZThbm08iVcU1eYth3lf0qFXAT38/BF5s4z8BU3SV
MIyYIbFS4xkKc6Fc50rit0EQ2WW7s2SMFR8OSa8WxcdvQRUjAiXpIALH/QbUzFQn
tasCbgcKO3cd/BxuxVsO/JqYvCqrdHqE5not8yWn9BgVYP4MQFwqumpGawhRKODc
k/T8PB17Odf6JJP8XO6HPBjamefBSnot2DfPsAhu8qN3G0v+yjid+2XATdij7cZp
bmKcqN4Fi7Mx964SS2i+UQW+CPVketCZhZ89ogLsxm3aye6DrPfabn85v7wx9UCU
//vjwBYyiCYFobrOMJzeTu9OnWnu+RuGEdXnk9spWgkMY1vbBmUDvjhP+B8x8D0Q
fEdai00RXIVmYjnEdCtG9r659+pN5XhtXAds7agij70vH8PQ0RFam5AkcmHP12yn
gpvePuImUzJL11XLKoTFvkkscvxh9d1JZptb1MvkeOIjFwp+RxO2vjPl8IL2ZPfx
9nMR7XnKrKmqrZI/MvF//fPKtLCuQPdbSDsYOvs/pNxOPVnYH7lxld49VZZTCSD6
sStc0HuVvRV7wMLppcrzNX5DgC6KEX/9AtHkc3CX/4wCQNuaIz+k4BGoK13NQSNf
L2IR/B+aLU/d0yFn3c09yAQGZEvpQ33vg/Ygvd2jsvN/eZ5/coeFwDwuHijWSsDz
SdO7jmpYNwMibSyqfvYJHx0O9x0sj3R8OrVO4RXTjNaqkQ4tv8EZXXqPc/0glt4d
6ixuZfwxZ0mgnzBefpA9BocTLRFTq1rxrkK4Fgubps2/1V0m4vSAGycw2rbrnrlb
PphQCV10w+PIVa0n11gg7vll66nVhXyhOKmhbm8NXuqRUQPOAe4197V6z8QRfiB9
Vi+Z1FxZdRJKfyM13nL9DiOXrLAZwfMDV/wycXNwUamHo9S4lEZ065aBUe8nFYH3
zjT+3OrkuCO5b85Hsx2stq+otLpUCzSelVJNJVGRbMlAJKSF5FdDcZojURwoC9jZ
vN32JWRiu/kvwyLEIXzQXBjtohJemLvxyA5LhosSYonxcLKhfAg47zlEaAQ80zlq
jb0EgTkDKAKwFMoPPVWQxWjSqU2vutT1VNfwOteVXDI+UAjlgv4b7ewEu5wJBhBT
H85ie6X41hnD3w4I4q2WtZIwEEvrnxYh9DNXjSKW0zA9H7FTOwv74kxos9VajvjC
X9YVqkl0KuATwIZbj3jVCDAJFbxfcUktBaZj+qb7S5AxStTSoBSeCo1cSGDqtV+B
osIp0P9KJglxkxJZv9rD47qdndT2CdhWdaozjnOfZ/42LGi7CrkeLZdEBALtQKlL
CGlPi9WsfRYwbrddpK8QUpbmGxfvXySWDGK2lQlbhpHhG/kdHYKxL0R+SQ1ycyFg
KqnVzmqZFMQlM36qrvxHRfMDAxzMXC5Ku2h3PitusjB0tXo51lK70+IgbFMkgxmA
muxXyDe3TxzFbdOewjJh87uKm31+eYNrjtjC9Tvd/ukXcUOC8yayOA/44y+FovlT
kc6zea1GmQiQ7RJkUVs7M/n2Nz8SqRILIKCc8Jl+O3t4EH+FKWbeUEgrLYGq8Vzi
uAsSAuQN23fq4alctCH2Y2oE5eZkemS4fy0ibSaVcqAlWrcZHyOKURMjnUzZvmXs
jl6IuRqlvCcmM2ks4oHe9SkBSE8Mb6Ye44T6VWCM1i3EBz0h4eDDz8bRu1edp/8l
QJqmCKBdtCl085jvWGcb9ZiPzfnL+QgVkZlexRU282Lf9GWKuZUe5P9r+eC1F/C3
fecjQctxJ1b7PPRLGXZumrozq6vs+8sVqK0chcX4TC3JtfjF7RlaPvp6HFk82XNh
tUDZtMUmnUHQS4JE+kaEmUFNxaR+7hq4dnW2Tpv7RG7kbhjjpuo7BbB6hBkmEegv
y3HMS6hYc6TleHo+NwohMv6if0qoIkIwjz7OzzKEVC9XqTvm9NUZL2qRRbDVlSan
myU6O3vjwF/WL71okrpDgvk+AhI+BAjsNNLDHJDzvAxe8ESU9KH+h1J+3gAipkvE
O4E6odyAxPhwNQpubonORZy50mnrkPWzksgpR1B8dIZrMCoHy4jtxSYurVrRQPDy
1CccT/po21kSaH0Qpm6d0vnRKoJCJMQQF3ieTdF4AYWkFPp8X+LuzYQIrFXKlpMY
axXp59OjbHQVIIvRi6T6ACtRFuituF5pp8wk6agz60s5c/jv6saGRsqyO+PvXJ50
NR++UEVZsySXg4SuEQhvVbzdvBK0UVQjyT7uqH4qKly5z9azvQNDO1uAoctYKCdk
nva2rs+ELT7EEkhDeustIdxN606t1yQAjmd/HuYRgl3bL/+Ho9GYuKByDrwk4TCT
Cl+cOp3Q56hq7n+H6d3d6T7Be3M+nhAnRPlSHUOZsR4D+5S9f1dMjsmBjJQVVUdd
0bTarzIfsmSUCe5hEjyyhggE6h9gS9oeUWYbRcj1uXD7by2+D46Dx26I9sv2nF6T
+FlcoGaGw3ZU/vYGVVtMWwcCNTJuAYwOO83nxHh+oJR94ZEmztkuUEtUTTEgAOnL
1Uw9jHjbk8lcRwOwXklwEPZHFjjZvypcb0LMa5zjlER+A1J8TeY1VsPbhjijXYnC
uMqc6ypqsg+F7HEAEe7zQkyD1MDs2IFKHxmbrkp8aLKGjuMExONQS5XM8orjz2Md
6o0g16im2EGWh/fCFPcvNj7fhmYZEXdeo92vPEMjdMuDJUXKS3VUgkySB6JISnyu
NM6HhnQ1WDZFvIasm5rXXykY4MedniSoifUJKvKXWpypmnCaehCh5UK7RcjeezKL
KBBkiulitS1P4kCzCELidAnM45D95xBzcownN+D9Lw6TymNt5sPtFUbN8S6sAd/6
KKWLqJo+pj2pJoGFUrGrYaaI2x61JkNwnJZZJvqh38x+6OiMHEhfE0zmWTVq9Aix
VW9nHT3Ht8na64lWo7+G7fjcDaucSmQelfV7vux3l2Ishw0WzQlyPjDXzJzEI0Ql
jLZDOPeGlrSREmGrSxzZk5lzwc/1sUvU/1BVdN6BOVymM3DDgxcfX+IEA6QERPpY
p+fIS4RYGtE4DprnEkkivrdLO+697D+Q18/kE6vpaTaHcQBwk1ssrOHBbMS1gdLb
uWCG+Guy4qpsOzZw1aIBRC30eaJbCZNosyc23y5SuwuyTHBgZx7Ca3+1tE+pt0Er
3xFLNVDEA2p7M96deuEcda8nrPfjXUCalWT2zifdJSmD791VTAO9o9aeGSKkrhlS
bnjK7De7aibzGWhzyrJ+ABnqftpZ2oLh8FSMXLCxcgxrbkReJ1mnxcUMaHaBfQKp
mU+48iRqUfMaCU4m+TNryvxZ/P+3DQuD37OfI52Da57SNSkX4SQGrxFNgHiInbRm
VjzD4S0KBPHxtXKbzUDbveg/1cdkt/U3472H/0EHreVc3lDETwd6bS+3Bj8WaCMp
GmhOxH0ZkEmHlz0vLWJrMksC61Bxp/E3rHJaK3OUQ1f8ZWNfBqBvB5aybgx3Vlpk
g8sjtidMfyshEOI8SlZf6+eJNXoWZlEfwLzvwsHv+byvbrZm2HrHj2R3oOZvkyMB
9K3XvyeaMEBaZO8I846Drvso4BJS0UJmczZRo9dZAPPEcK70kqVkOQZvBuYii0gv
rKDoNi46kG6cNzDUKqL3im19gVRgBkxMUkzNI8mYp5MmoQeoZ/UxPLDJB3YQ70o1
M0sL+G+0zORrXTjvN+k+2Lp4B/LdzXXQqQ3ismpED3cf+Mg2TADchRLRfAlOaieh
jYQRmEhWOt6uI/tNEND19G323vV+XntnfnYwLRpU95s8IdbA5w3w0PPnieOkHbFW
kaiAmSj98AO6h34jG+lSpWCp6rKqoA/vHGqxQKjvLQK3VvxyjYDFVjo1axom0dPa
Jv6+ql8elzmMd/tZIUYb4qlT6zZqpdY2ob+rY/ynMGHJAADEALcpVKX12Zmw3HSn
xDKPwnC62bSN7NlHapJydW5MOdWCMmU0gG6X8TULvYdRiXQ7Mef2MTEP3verC4NE
RkTTY9j/drPruvUe/UBRVa7dJyPTXSa/LBnxie0XeMupqs5gCkXNgzbqxee2+jWt
kGgADff+S1tpdkwa8xh0Q7nKzBrS9Lj/ZXEPW9VSGuTpBTV4/TK/3PzajNm7ncmI
nkccyImR+WN4mYrCGNz1O4G06iFDdjS6fkcuiOe42zvTSDXZmFXTgXeMFOuAU2GU
eWaIjxVdI9nQDeYwVnAGucsjOMF+TCOlY7NJR7PwtsZnXr2bFJfHkBQx0RVKKiMi
PvWV8IE+fh9e1bQ4TIPKggNjtwNOsP0cYtXz127WqstSOs0vvQ9PrpNxi1g+o3AZ
q3XL+5doR6M/IvHtOD1DPA80bU2kOxYaF33QFQGxB7zxCRms8vQMSSNcbv8SLcnd
8tk0ygE1vC+5BcEmFUNt4m1yS+0jt8hhRWo87Bl0hDd01IHBShmvZHOuRDbnWiQw
bPcFmNivBve8DI1IOwaRAWiJVuonn7NdSOlwWPi1tewN0DfS5e7yIbbKhaqDVGZl
bI2H8O5OkXkJMtBj3Ry6oJ+pmRmfUVOJzcZRrdM0lQm6tCAVw/0PkzQKaaNo+Nfe
uabtuSRNmtrsao9fK3XJCarWFWX/ivXcoz7RVu/YHkaHvr/V2CIxw1hV9FRC4vCW
+LUou9SBQNeYIZ7kvZRfqs9BeMYtY2vp+azZLvBNDrurnCrKJJy2nyWfjwmPITmD
PNNmal4sn14+lplDWaUMaDD/ujYo0dS7u6p4sIaFu5FSEi2j3W+bHKJXwJJgwKOs
zUx4DUi+wgPIaW160741lTjpkAKU2jNFqrHqPseGZ+cZKxISwJFrGX7udFPZzmxT
5YR4j1nL1G8Uxid9tIEa9jK3NPPOvKDQNZmlV3KJ0pkzUib5UHwjdBfx0/Hz97ni
7MkQX7XdyLJF8KSyU2Mns8NHrIoqbaFlFYTxPRY2acJ7cpdyTFLkiv+la8btDgpV
FQxIGIQNKn/jQ6x/J5aJaEtB0kxnVkzMLh5jXW/cHrucYXTq1HMGZtudMS8dIk9O
rYx/LYvzBc66QDR3XhUHJck5T0S7C7KSjTjX73q7iobH87T+kN5QiMqA2EXXgce8
wnItEfaxou45K15mpFdncwmVS+GSblbZVn+M+f0ZBXbvCAk+8Qt8aqjpd1Cxjtrk
9THFHk3XKep8tod7WG1QD32UveSoSSFFnYkKBEuxDXZl+r9r66GsNq8N3O4tl/hY
1gB6FXcrr34djV65X95OXstXTIUuMQEpexjSjhCgnHms3Fbz6rP0rBm4p6aemUo1
eIPmtJvaXxszYE1/4qKnrVxVavPeae7tzftV8t4cU5HYpmsTX2HYmp/U+hNQ7QEy
uX6mW9/MBl9tc8ScMn7O36uUaWbJH5DNe2JGjb971bd0Z+cYcnVwmIMjjEq0XTAD
AFMW2ClQDQUTl3haHfbLK+XuZIlNHcWHppTQK5fYLLmFZg4kCXS8GdrbNjL4BzIV
0wHMCINej+v6an+S4PMLPN/zpQvab8aA2Z3XW+x9FUixZ+fZskO2vzSEQGXYTdLw
0yHNx820sTyaaHtAifLMzj0dNasE5wDCCpF7rlg9YDdVEuBWKEebBgYeqYq+VcwI
HBB9Qb0/WT0XvTfr+qLnEJGZa5raYhdSFHpBe5/qFt8mur8sI+cMQdJchO4rQc5t
4gMi5ikEwTATJXWFoiAMsq0vhBjAvv6f3i535n5q+p3em5+cEYAgw4XJ4E9edmoL
ezSeD0nVGjPDcYuskJWtDpOWWr80KnRB9T2cVhAUj0aTW/hy3RdqQ8qwJTFPfytC
aeJ+kGSFsRiuuwKZ/OIXn0Yrrfevt2h85ZghXiJBKvlGa8Dsavyi2rhhX27CyiFP
f84zWf2uufv1KnjRO3eN9hdR8jSNObY58wcQzvz5nLI0sBu08VfwCTv5Q+hAuQK/
6IAS1gCwYrwdTfz2GZZIL3U0wa0agEtHH0VWVSy11usuQFA1xey6X3uheyBJlcJi
pZBNqk0tTmfgju/QzIPFpbjzgJ96bdCDzRxEznVq6FlXf1WMAaVMCD6+EHtZRmHU
TSYnRK0o40xXr0xVAENZ9UmP+vsuVLLu0yFFFQW9VgoxZzcIi5qzQabDTe2QXYta
f8GyXzy8nwjutjkgkpQ9Mj6QTJtHiphSGZb/KWU7QeaiG1xf6hvbbZk2Vy2dyoDO
eLlQY5y8SUWKu84grj+wr3dlAE9+3kHvabNLa5P2CJ7w39dlOwIzgqTMi2HhYVyG
jS+rsQ7ovWQjJ5b5ycbE+wm1mOzBl4LZBC1F0PnlxkPTWbS/G3X5HgLuD+35v9YF
pAGurN3jY1RWpreL9k96iC3IiqMb6X7CQBa2ABPNorlr3wS/jW8GjlWl5wgm0yGa
geMS9XwBroaUo8sUpT8SvynLf+LnELa7gjAb6nyENONOkLeU7GDLuleiucILdBbe
4EVlrGS4GT5hEHWFB9c9M8ByhE6pbf+Sc+enXVzW0CjTIEr2557LxYAvx5qDluE/
8zjGBTA6uLkqQ/5getsLrcalWKG22fkAjV9f/zDsiyEDcYMibI1HpXLdwovoYlur
+5wuqg4E1uspflmZB8tBVjJcJbZPRYne9vTrvhoGxyR1R7hSqJGZm27b/AsrHtzK
xrc2Zr7yLqiRmaxe7mASaJ5T1X1MVw2JVH/clSy4jEdUcTGuQJeK7KI9qe4Alt+u
gtxdKwN43aoJKkBtLdkcoCa5HY6xLZU7hiU92UGCO8l1pdCrZ0h6Pd+8WmQXKTrC
B9uAC35Avs1oVeqwT5X+T2GwZUqZpsXEdOdagNzovChB01+TjkQN+tnZPZr0Whqf
GdCE4v3Zymqc1yN148XL2mpSVKeBDRXII+zzA6pHVulSiPPxkKlsV0BasMV4ba/u
UE+5H4NiS9kMCvTlcACxhBhWHyQhVqCTeek8AKxJoTw4qckcSOUVIen7xUehaWP/
PBqmlP92YB208kNHCySrOofT7hV81IAXokdUWtIwlIe1WYYLrWBodAmDav5AkRxv
theslXkozm87DJO36KLJitlaxNQEiJ90VunATXw72JuYJBseOfzs7j7iilDtWUWr
vTNTkHulVk6xFS0PFQpVF6GJV6nC6I1JdpqbPvm12ovLM6T6hGAq2l7JyT/Ue+Hu
lxGQLRYhu2jNTcyLAy2rsNcYp/clVVqxYzm7/r+I7JkS1c9DVGRiS1gyBl0LBNPY
53Y+hZLaZtV213yDLuG0UYwUTc3ih3WefZX1/MhVmWJCKzyRO9LYKABllACC7RrB
/eSQQYPOEMYZSPqaFSN65ftVIcyK/g8YdMgmthU6N/29wPfT9R3hVLQUWhYOq1kj
6kQtLZQATgkuRsYDrNacz969lpqryMkqhA6jrR2+vZaDeR12q+IKGKywcxzoOhCm
9z1Qy106sqJor7e+do/9wB6CuLo1SfFn01UxGLa/fdPL/lVxyLA6JluJnNxvFwQO
hjx6NmRbFR516llxDjRf8ZKx1IifzrBSQyHmXfkJBCv5xCErQWWkdBUorZp7aFoZ
10VKdgGAHL+cYyo8u4+FqAYEY1i3GDcG8xQAAkWxi7kf6ctFyZXkl4LpdNTeD9cd
EKF6RFsnTLouKRGVaZ4RiLdSMjSe+8Apjnqs0R+94qWGx486i3C+WIHwnTGDo8Az
vUxmli9/t+T3lFZgPeVs/uaX8wxxBJiHBQ5lGf2H3MqmusIsxEUGBuCFwIsDzB1m
+19y4/SZqhXF4EVcyQJeChp7QQHmajNUZeSJto4Qyn30o8yEwwScr4gpbnsiTTNJ
MDdBROYfjfnQWAHIpD5a8/6td6pO/UYgbqXBf2ENjxWG54tzUv5wscKWUl9cl9ia
Svx/Oah+5ILKstERuqHeJZFTy5CFsEikeD818hiDzt8+Rtj0+jYNgTp9fTpj1+9G
2+M9DTBZDlG51oOycpPDxJWogexrVWUpxbSjCGzIPPFu6erTeVKGx9CDMYLiiHF5
VutMsPiGqcH3NlpC2hopl3BtStpWx/FsfdAVE1oC0BLMpdBNHPhOBKYJ1GojlOgn
x07ljGncYJYrLOFiPubOhgR5qC2Cl0OrKDvr/JSrxr1g9K1dzL+FZrO7PdchCTCR
8yy131IQmkCNu6qtGiuRFZivgXB1KSV1XHQWuVkUHLEm9iDZHEny//IvxKX3WM25
3Xk6lCCWrkpE6TVS4NT25kQBdjcvjPuS7WTJ6/BmkL3jztfyUwiyQeeDHofCIoDn
1Nk/DwKZWRLn0IzY9yHFBmtrtQULDNBvr7N0O8n9zB9YvWOeDwGpL7mWxfa/XvEw
q7qAM6+EmGUfp/m4qCyRxyvdeBOBWIKwd6m8BiW4U2BTbjYYilGWHLBtgoL+UMvy
CITRcOOzrZBkT3CH00Z7wk4ljUw3323B0YkJ8nk143/tP+sH2sZgqMKpA7XHn+4C
Zb3YmHhYzWbIl+izBgp84He4EmZzCO4O4P8L20lp2WI3MlDTW3ieNNAQdFit7TJB
yPbYIyz0xEvmkMY24Dhhh7D+OvDywGoB+CodYSXSNYSM06IZpj74bSMOGk6VFb3i
aD/Q6wd+5gb3iIYLe3i+wQB7T50bK85Eiw7UPmHQaJt1CYMZS4eXSAiLs4Fd5MIv
lOAvG37dk4wU95t+azelKiQxYXOWMikNgYztKSiBJGu5ywtSEeg8rxwM+hilwuz7
jY33Ynxt+7aYWoxrK2ynrd34dZ0zuNOBUm1bpXRe6+V3L2dglpgQGsoF3FCc2Xva
lhlr22tPBQCqoe9VftUag20q/ElDItWEFepAKXlZM2sn6nqlwGXII3d31hStQqoz
igusqnK8wqVKbB6zgFbPLrXw2+b3ZgMhDYteDtL7PVf3o4PGgOcA2YhpkB3kG1tR
3izb2BWRKaN3vBf8P3KYtjtpMCR9OiwL60PEvwD7BDTdxkm3uMhPp0pyEj8dty4n
VVp6Iuj0JF16NEUeeJzGJPoFosU9iW4agt2xBlp5HlLGQEjcfGsZdmXUwmtO3eMW
AeusrFmNwEcSwi4z49mbh+Y+ZyLahhtLbbInGHmmBsG3z39DFjYU4xcM38YVEHJR
K8ek7cl2QlSyu2juXYyS7SpjMl2+pSxKQpn3gDPrZ5jv4K13PW4QIsaf04Nd4MVu
oRLQCaz9KJE8h0PYE9IepAykDqsfzSCbTRneUVi09JlMeXfYQbvFzQwq3c+6u+lW
stY1nYpkH71+G9caqjNhzxydrSs5LcVidSjDAFzqyMtLRg35zUej84ontF4Bf40J
XE1H4cSgz9ti+bcaze9F4poSZ0as3hXulfGGFSLV3kdJc5nHmQpsRR3Xeki2nkaS
iLyH9Ja7YFpq6qOjuNLPb3Eg5tXbT8mh98LIoNNVSZkAk7zNG1vcHRdtc6zIFffL
QW4C4utjaNh/orioEOtLsUj3Z+Snz7wv1i3v0efSCIRDhqAThfPexIleN5esNg+u
03YBgnEilK4nimI710/76SyLEb9fmHdQpVhCZ4rERjOR/fMIhlr+WH5rohbjAZP6
5+zKWeEPhSSRT406q0g8FH0Wio6AEY4tLsxw9JMKa0ZhObprkh/KMrHOZ7TW/hRd
/q9nQSr8JuydjCjDkFfRtB0G5rfIkn9t9uDSkKrbzmCbb+WaOeTWfmfJS1k5e0OS
SwYxYS1jSl3z5kQaXq3IIElqK9wSSi0O1wnAPlg2GsVF7q9adpOR8csHxOKvyxGu
WywU4AZZOCpOHgJLtrh/HhS4/NvVxRcEcZSQ8XrDrmV/ljktdTDh+hNOJDRApRZs
+ONCL7fGoKn9hDSKFafu7RgAuofJMTXhkm6/QqukxetuqPxddM8G4twIkxc9e07/
fdcXGNNhmEpc+MXpc8MYROSIDEblYRc/sjpmszSn3MmhGq7ykFRDXkx799PxZkFD
zS4TVJv5k1pYT6n9cV47ogXWFAley3tSoFnQH+CyWayFbOZ5/3laOHg8W8ajU/oF
2OzaXq+ZctO74JvceBtdHH9XagHgCW9aC2Lymna5vujS5FSOLEnn5Ri/NRLSJkNr
/AfZrn+PEg44hI6D5B+vk+Jh5Xq2oDxRQUXAlCO7rAHab961c5DMEglOgakPJB+I
sMP6ypI3/ItvoMig+Un5YcYjs7ZLgq0QA2jMatnNKUc1twyX8BWNFcTSOGEd0m1r
oEaH5iHlfINp0mqXVuQn4eY1QV0MOLjFKDqf9qzEBvUPFBSSt2s9TiGN+K4+G43m
Q5X13/W71sIJWxRuLs36roE0fajO5cdxDfDcbraHHGnSACW7l6cOc+r2Ps3COA7Z
/ECj98+Juvm5LDzfKvSrSMGVE/RSXXPumuEJMivc2mzs18TYRQPy5vbYYA+TOByJ
WevqHetVueDwlKRwL7OxwZMZqIH1aLkYRiaWnJYkHreWtrb19hl0BH5pBP7hr9ip
ZB+2ZEvoBe3q0yXE28KHQA9qpapP60SKpQDYkj4K+9S72VSEztXgxulrUPes6bR6
Ku3QhF58y4GtnhtNWkFMxVh1jIu2kCedn+0cyqpiyKk2YW7umgBGbkCei3YMUhIy
0gk9ppvQTxCuTw3LnaNu/SrjNjlJNxYOcD6HQUyBsfG6C2RoI6K32iX9jtiQviEs
FvvWERR2s7I9uGjDwk7Uckcav39I0q8pIFS/HzHjZ8b07n4jdTnujdYT/QCc5yYs
+PJAa7UgFcsO9zTsuG33h8hnsdl6Sha9Aj6qFqfCah8LzAplL6pSrhCQWkShWdJ6
tJEhcHfg7oxd40DsVuDQbaex+ocrMopCkWUhG5ozbNmA/+VS2USS8jdWPqxB4Kcu
molR5ahChC11k47kTQGs0lPrdlgyJQEJ9KF6H1mrSIK0WSQSubj2ehlreyLJ1J4+
wSnIWCagSR7APbjFY3X8+nnmnmmXgs7jh0aDeqwqgRg7HQNyyg9av0lH3+1dlf9g
fFr8qYukLMjKBS1H1d8Y1u5BlK+thAs79KDjdd3lQYQ14M1SiC8rydHtrufSJ2Rf
xQQPhp0FRSCo+yeimTCV6Pf31CnVKUWDRAGmuSOyuEVOJxEtJ4+sqmBlon3yi6EJ
terTtlj6LdvAnzH0ViyOPQQao2xQVFev4cxk6aTHpbqQRrQSCqY4k9bJKhlxkPl6
B4ETUdDKVpgH4FJDefueFPkR3BPJ6ELyUXxtOJYeMb5N2nAHLEcJL+C/VPc8ydQT
XiH5RAsEPKPgBG80o2p77HYIFQyA5Yo+YL2ju+Uf4wH2EgLCqXUx6mjkbwSxyrSJ
ylmvaMSCUh4DtroBflnnE2wNvUxXej1kVMWkt5jB5Jzks3UB7iSUVjFUp1yOjvQo
H+TZWFFT1AAL8BNTZUB1kpNf+XGeFZngwuXv/GhFJRo5Q2iTYxnI7N4bwlZJGVp3
XQ/Av0F6BlC9+EZQ+PKsrLc5c0oT5PSGzSL99CT8YP85ILqbPqQor31gBsCvSXOA
LbVywjITHhLYbW9KtF1UzJoC0pYVbL+N5FVQQbIwuewFLARzO6/fyh7D4xO3cxrn
aUMMl6Csm1ZkuiwKy3Q2UH/1xupnIGsUT7nh/+WztaVeVGcwhBnqsELAE/PQiZG1
FPOBMdBOWHhMM1Ye6jYwHwLuIZBbj74Z4RrfWALB7JAYJ1CL1AuEaYmJb5/Mf8i/
3tbcR39UrOdKtiRGAMlITmb+ga0ZrTz3cTb6wGD9AhNJjD6ZX6Tv1P4MTj7HaArI
fCfJqaKtI6xVx7AjIXhfEnCkkx3QUf7vdA7y4Do2vHV4L9HWmterK2hXeCf/RZp9
t7P8gUsTmwNLkS35I3aQNFIi3I48I0nheMjvwEa0qvi/E2w56AGTNmz2U8gX1FgZ
3NQYQbJBXu7Nh6dOqu14cg2aqv7ETsZAlohFCenAh3BTNJKn+5AClW80hTTk/3N6
Vv+pNsmy6DQ3NICRDf7fS17oVDThaHbo44H+vmraBhi0c1jYtXkHW3nKOe2BS0EG
rdZoLLyjkP66cuorhGS4ptzOeK/1tdkxY/BqAn/WEuN1C6RpVxzS0xv5qr+5xe3F
8PylHYXoVd5Ie+HJ0O3PimiD6hWAkTH0B6SX7EZtPEi3ru8DkSSOIxgM9//AqfU6
gT/5qzUITO+UlwcJdw0Pl4WzWgZlGpD/RAhHtC8ugFK+/qs2NNL4JGiTP9+ekV6M
W7erI5S7yupiaatEzq4T4PrpjsNUwXnl84geU5qIQVsIdW8pdjLUaDCFT1OjVqtf
f6Ckp57oDOa3T2cUiDX5/ROppQrram9PfBsnAczmdvS1QBiB5hga55SU44sxxjDY
LOIFk4VcUSAJi6PFOzZaXSqOy/mWK31Xpi/Vj+xowg+uAqvvKyNkEYRiR53lmrc8
MVzyVAysxsndgJEe3eKLnF+DxNEj6Ht/de0jRApO7swIhQzf9ZzC0Ztf0HgCz/mj
uRne4jmCyEK61fgEkh2qBuvr1N/Vtfm4G3WsaOoplaDhMZvebWIIQklkQTX1r+Kp
jrWM81ryIIxVVhS4iCDX8ZZGwwDNe3d1cZ0vk7Pylqwv+LjXyNBPUjPNqXifH+AO
FLhvhSFqmhrdA350TXCTAmV/xkqmEkA97d/aZ75V8Z55toE/QH0YVi1jQOLQ/O1M
5OhMxEXvOrxtGkPdZS4K1orMiAwKDZDMO+1jpi+IEUcCw2goLg5HrRTufxl7ZM6r
HARUwWp/M0WmwIvTP7IQviW613uSHvQ/yOGxOMi8qrPzV8E/FocEzOEfMunruT4A
gXLVlywfEHx4VjYDSl4hS1tkNF9YLfv8oip/i0g5hyNL2XE/c4HoqP+xl4ZK6P00
wNWY5Whm3GgwtikiC1vM0bDFW2GTDlh5tM/BrXcL7QM2ow77WZhebPoaidZt9D/z
7mhWj/iXm+LMjmLwCHH0Lk5dFlUt9B2X4oHLgIjuxFH1/oEBm0WltEuMLsg5o7Rr
076miRH+kpi+7do5mRy+pFbMB79S7UIH/WU+D+DhYj022KZtwpgb4UZNoZLvHjFN
seBxu4+XWeQ+nFRRRpXZQyexRqYxvAuCaLGXnRaCymdM4EUdKAUL33jjc+0HkDH0
JhhT4l0wFW4DdE2UuR7qyiJiWF1CDaMwU3LhGa28RHAPBHom+vtL32UXVSe804wX
BqezKAnJGJ10Pv3iit64YJhH8PpBPcePU0rRCAvcnAuPavPvcK2Erpb3kW+XYKRl
Lj50jHa6McFiF4tU5BndjvkmF7JldAUe0JT6YYx0o2AFOMNCS/jhFBliGa19vBxx
wZEoWVbrKL8fLEcvBU1clPTG1t+sVHD8eaHmaGxM+2EypAhU528mQBoXoqXuCYFw
6VzkJklrpdLZGD12/kh0BM3dRF65OEXnrm0sn+8jzFMnpldgvcXZlUmjoVsxTjNv
iyCFHfzM+vL7rPTh9+H9IeIk9ABg7R9re7hGAyMJlfjVoP1QG9YZyxDtQi6Q2Vu8
BrnTqF6kl6+8UX9KnvQLetPL7PHzgM7Hi8hKxjOHE9GNdP8OwS474plw82J7+GKm
VqOgNoxdhKwhu7w7HlTz8zyhg1ZLbFpj6rVOsv5oGolUIVBACvRGoDXb6PIyHygB
Mam0VaU3HnlgV3RwDj+ZnUXga/rWrKOqlIEq7xbG36sw9sIezBSGGQKKiHmuMtZB
htm8IkY7DsB8vFs2K9OMXYu6Jn4NAGI7CKYOz89fZ1aGLXSDmSnBYdzJbtf51y2s
QD7rWkpMCc6d9vaKD3bRiGWqZ9dx96rYzXoQd+xyBFhFEtER+n/QWLNbtV9gsCmy
SA0W4VaKYtO+ehyIYdtzpys8QRq12Va/APLl65xrUkwvI2N6xuzHVgDedEuoU7VQ
JHThUV5DcrqyJgrHwSCBYO4/IQhO/hcZw7ZBY+NQNBRoPh7yQZs+cZwfD/tPJkdn
u0OD7PGvumxgW5DlXlnRonsgUwTKt7zqzXtXFGLatLMrjw9FAfjRXxNiKPWTHyjx
w/zpoQcUMm6kEX+HlCK6bQHhsNqTA3M2vBSYaDEe2HzhTUsO3bTpZFPFnh4KyoOZ
yISWNW/m+DmTcnXCwaUuktvKodeNeY924ppKjSAmhG/yyvNc/n+gkCIlLl73cWtM
LJfSHlKSMrnftgL3zB98UTjIYFImwVcQsSlqwniuFyBzKhsoeXD6tk6ThNI+6DTQ
j+kTOoZr781h/iTIYhotIFjnS+nnL5EXGJcUpcokbMxPE5MESgDbJ1OBd3DGLOaJ
mKDsRNfyDsIHeGQE+ZelpYwQY9nlUFkf97QC/gSQ77cIM3Z/RUDnOlcjOpYNTcXJ
kPTjk1HEwp8IBtKhiwCtul5ioBIjiJufsCV3+CWMmRIByiqdMnkrnmGC3ivqSbUp
8eLO7xbFehNJeZdQaCyejM3so/+ifQaHTLNY6J6N/GUkSXIl9nMqOuvCpugfBQyn
q2sr2utSIKhpm6RB/0A1pk4NHG5h7Cr1qw6w6+f+Qh0k6V/cPcs/qngqA2xtAPId
vPLJvKOtcI1z4gBh1ibebBTYKFFd6WNb0KBoYeTgkTClQtZ6GMIF0/3HDo5Bs8qv
jgY8koI/oZ4ewQK/KxdcUg6QirA41+EzlEgnj7l/MjjA2garfFIgVauHisE1ibp+
GmYitoRPXA2idFvmRYhO8qZjOuxyr35F9bvkzwPrzVaaqp2XgkPwew0yeMESkz3u
TZuNfC1DsYSi5UQ8kMlx2ZiQK2DSNJfHSp6CPNM5raGUTr5u7ngweK4PCrMMB43Q
DFQbDHvCspl9z8s01hjhenK7t5vPwR/jA+5ypekDeZChEgNn+LGh/6vwUneeDNF6
nBYr6xFePLz+8IgPFv1+b6R/psJzwyKcqJ4mzO8lr4nzs/6hkNFQpIxZNu96mj2h
/fDQPx0R3Wew+7CHr8EpvwBqn2xEDtI+kyKPDu134F0cyrJzsd5u39NoAsTH9Gly
xfyTWgbSGRY4MuFuYOHliqEWNdB0DIH6G/fprz1llL020x/gFnhArBBoWo3dxstm
Rcbupxu3Ir8VDlRTgw/m8ImKBzG8cJUtuSSrt7mw1rnI9Y9uEhiAPxQoCAy4VFxe
Xp2eD+S49mD4uCaqqh0OnHvtohfgu/3I4KNLux56veeZJA62qRebTS1IAMgS0uWI
oO0GLXFUJ2usgYDRAF+cFlDq4qzb2pIEL4jSw6aoHkDNsUoJdZDWetGbWjMb3/0Y
P0vVQ8zkuV8vCS83A+3rpiGxZEioGazbldZA0gt2aivZhTU6QB3KwQQD8gUpSLqM
uWbHQcIO8riOAWOTD0F1xcT9azBZeKjQ/Rn43mV8OnSUO+lXDj+R2wiJX2GiW8ZQ
hgN+pFYpUqm/0Dtz4oOnaDHni51Bf1Me/NBvpLpYh5VvH5DKm+BbcHYY8twexEci
q1B/VhLRLbLHb9mB5uiYfjU1UaHKUKQPtqyRx25dcTd9kVZfj1vLhasZcWlyBCm+
Cjuta1elyj0QZZcE37D7ZlcjirXpWFMb/nLPePu78syQsqTa171HRGt1w5gOMSom
PiE3JwPHR5hMfxOnijNQfk9qTcVcMWL3p2fVysK4i5SR/IvHBKz42+MYcZdl72r3
mCrACEfDSC/dgytsyrRIJF1Mwc9dB9ocQMlog+wB1KJCrSDLOzVWBXENokXrENiX
mZlBuNPzZGgeg9u7eRvyiViBvOd+zIEmaCVrqluAIqUqpXjt7++pd3iuu1C4ZeJo
hoc+Nqlu7uQLo8GFCjU/UFX7plBnVaeGetsZ/jSXZYQG+ZSCB85MD1kIwfJrjms3
jawcW/VgNTnI5MBr1OYl5IkpHpq/fdBPYG4RrhuWoKrn/PuuuXE6mYC+PfNV+i2R
TQ7nyH0t0WFa9KQ13acGfH6f5YBH+/kKAyGaOJP4B+r0/Uhdi7LnO6WMAW0T/UMj
WnrM8Xq/Qp6fQM7wLurbd5zTGttJwqugVrItiFCu4l8AZowPtJPlEpbI+eGO24OS
bLQUio44rNYOkNtqYefkGa/55wi09LXW4ssKEfmfjBfDU2ekIKWJoE3c+hWk+a3u
CJ4s8RFPRQU0JBWVGE8AyLd1UJNakAZQvomB3d0sDr2B3YCza+LjU2xUFtHYMdTy
jdSA0qy07vv4D69WtNCb41RSSMTyJwQdh/k9FWTCkyihluYuejD/XiZML1KGFHE2
CMo1Rs86t0d1gEmESJoE8GaHPeRNlZwTpAz6lSyRZzMwwEFj4I/jLUSbGjrus+5e
ejCKR7mf3Rz3PJof8IM8j0vvA3pkIQkJEKePvKGD5IG9Eyjcp/oX3vBjkcgIUSlU
U+y6Kn93d1AqBlezmxRLlDmB+LGm31/5o/5lea7IY+y7O6b7VDjDa68SZZGyUi5i
GYnecgilqOvwze8GDjxEgFwrjjC3w4BKxV3RxbAeEfK5IJj4NP+CJSkvKbtoJHFV
b0Ad9sohMO94rJnj/XNLiNPLQfbyo8aKsjKuIXiZPPdnQGdU//x1hj9YmDPIdOp2
NZ4emGM2QbDLVhbckZigcKStKozjWh4dJXSQ//bgflJXEvpdiIME3M5GroShQJqY
GD6V1E+2mHSJWUNXmuwuUapEOF0ZCdigAT+byENlw7gKOn2mgb/IQi3bmBL++ZX8
vn/1vCERbLuuYEi6ev4bvyAQW0q9unIaKF4eRs4H8cycIlgRPEPYvN2mStloTlkR
bmf1yqT+IIotJoAhjk0YOYSXuy/Lq62C/SANSlmGt6RvAkCMB++73wOvGCuy5lq1
QBxJY2ivXvI8OPbRMVGa6Y7ABq6XMqCoiQUBvcrfmn+x4jreyKHmbIoEaF86W2qB
936iMzpl90ol27TIR3QAtsWzlcoNQlpdrC1SuIepA9VwgYzSzPxq8Vx7M6Gdu0Hy
IjOchqxcm8WStd7yn4prMUZP5VXRxN+o3+LXBxrNzP0u7hKqQKcRL0U3yCQrfSqx
v0LsZeF+ExHr/JDqu9OsTGRRZFIIfxG/lXbmwlt7iGszDc5TqMsj1lNqf1T5WWoF
knmXxd0lTSkM0BFlxr08B3h3EjRSXqnrvBUurL7NwE3FHM1zqLC72VD7QCsPzmdh
7SxVSU59eHO4LPhXtu+7gzZUBj6Jz5148SnDyfOE6VyQ0IjmqkgDXh8/UcFtqKLC
LFHXav0UEhcD4ayOm3q5qSq1RHyQGW/IalcrugLNNP9LjKU4RYJb6QZPtaGVf/rL
4ZtCuGRjYiyBNzRyAx6PrNDNxBfuI/QUSO2vgsoDWmQFjJKOl9Fbspw8QUiHw3y1
yRctqP+BHpkEMY93g3+3+29i6FUxjNVu0yURF/fNDd20uJpClaHyXTRd51//HbLX
D6VWRAsIB06tCbz1XlVhjkaRCjrbDHSGIHwA3hL+UFudgKUwWRTkMswOuuqC1zbK
7Q3G6TNcOZRV9sMV7g0TTR/ds2m0lP6UpEKG3Do9/OxMJFQjv5b9twyWHTCgHgeY
og0P2DgPhd9IWnGiUXbL3X1E2KQiRkKNiO4B/FxC5/UwT0ut4jMrWfcouoYSw8wo
Tpa8rcd8ZsPgg0p4vanpvUe7TcvYdWLFaon45hAte9P3jwXAgTMDj7H8fQqrfs24
KAHdQtKrVGC76G25rQKrOK9L8UuyrzoXxPbC5cLqQtIRF2Oh/8IG2eIf6iZpwKSx
qX4ftM99NwrqsooufBW//O33oM6Nm+Va1rpoda1S/3Brpg5zFUs/6nzmWxAel4sD
nch7EqzdW82onO4BKJUZmHcRtaDJZmuoFUlpwXKa2OPTv1LStP3fzgoz6oGlrl1h
0X5zEwW5jiU0M/NVD4VgzY9/kWYbB/9m6N19ps3gGMJbPpn6X65SE9yvLv+UDR91
b7uz7MB/lvO7XWoeZ4kuQ2QWmaO7euKwUP9cH8JE1dhrjkI1pzM0DTk8sitPm8dU
C5Cswbi6u1/JuEFDu4IwYjOagpbGz1gvS+MEPsWUNm0eBe44VqekoBBkU2x39ofC
S+oDqxXhJYXJdANCkmzSmJxcL8nYiq/+KJmscJQ7TUjWCw4qpLSjEZGf4dtNCAOJ
n8ElYo1/W2yHT2mwr95LVZTm5SOCuLOqz7RQxaruOlm9C78uyTQbCPqfdE0q4cyK
3Ezn9oxDX3fuqqMN5h7/teZ4wyNzIGekAn6VHilkAInhN2eQKnnaZUPaOvgYX982
Sv6wWPgusAY9w7Nzei+6qqpVLvoPIB8Jk5pZl/GDqHwELVxYMPK/uKlOl/R9YQny
rnFMsMO1PKvA7aG5eS8Bz+ZKcqoj74wuCXNBwPUa66ImkGR2eCcK9+3oYXci2pVq
RcA/OvVoGVKuqCaOiPzrIj2bh6PrHBnxTz3ZN62obxPYVkrOEH8YLxkbBJI3Vz4X
jQQhZ8F6LMrnhN/FScEhAfWC3ve3vrsCo4uH/+pKCoXErKtyoFT1wckml+zWr0o0
Nr4rCeAyFtwQxVPJJH6kt4BlTDYl+m0EycEFBJ3xGfoaJ0AC8ZnAl1YlY8IERGY/
Pb+HJqnMwXOn0ld00MO4JJbqC0oKqMkROfXrpI1+Zf0GL7nKB2OETXiWyUCwiilG
wnyLG4am1WaTBuric2HK1H1pNtl+iANfZv8UJ/lUuMXvHc9DNK7/QIhOW9qHzLbB
UPBjVJv5a4M9zsOcH6JbqGJPz/1a1TqlIkCkFewCcjDx46g7bjlgEftVj8z5kDXI
5n22sduAg4isG23M4H1Tqlmrtg1wduJg+BG/xcgzzIOxtdQizYVTIlUvWFw5i+3X
IW3+Zi8q5kbpESocAFOh4qKf88kFAWBqVegtEmejuEOLU1SMzwYeYCGQRZXg8T6D
hxikI+xIwMKprMPYEHF0vZZx7/rpaAFIWxzbDQFTm8TIAVzmTBHpjNXLP9XNjvxB
pJk/DzT/o11CqTt7B/I1QtW25CiLbb39HNh9uScRtF8HRG5NwamidYb7zwkn3tu8
XBv3IaVkxP/9bqloY54hIlTXk7gCnT60wbRrZhMV4RejBANHYXMiq6cT3pIl/Uqx
Vt91NSOcUX8TdNeatWIfqgIdRKC0uSx+xhIapajNwKow+qKY7Pba0rPZ94rURJr6
FOGK7emN0/FdkiFRAuLm78CUJUl6LRqyzL0V0DPEyW3jLTtw+l8oSDUwECgEQjGZ
BezBg1vR8s7xaPSHsSqAgT4Q0LJiVn0JP8XtakgLiXuxt/j77y7my2GkyYgbwTua
nc1XXHyp77YCsONt32zA5tS/DCdNgpal2igY/1Ei5MG5/V7Z91IzXOCIoz/DZe/P
z0SrLmmtJ4ElEXNIx/Bp/p1Rly3XS6ZPmOHgF+OyT8wejmmrHrhHZw9vLuCTAyBt
+N+rR3qfHhI1hY4I9UF5ShWCct2W/8ZAQsn8WbUMtE9lA0GeMyNxOIFTfs2c2i0b
GVQRzN+PGGo+KcOy8paebpfa1JU8xKBmnZkfsRksQRZ1wWztK3hgSRRJWj4kTkDv
zJK35wZ6bjC7AdQbGc6ys0TbwMWrQ+LspjmbXpAFt6FjgbgBvWk853l/5u5MLzIx
pJwueEtVhclz9Sn2C74+Ar2bpJ4yjSKjMW+xGUBd0zHQGeRbpq5fxmRr9J6q4b70
GpX/4QEF9XCaSb/abJ8AFq7/0gkdBKPMA/RJYXFtb7PLrJ2LuIhq9I+ysvlgL0W8
OAFpEIqnPG3YazKm+TiHyerv886dadziyNdnH74D65UwkxYDy3xnrs51FufaDRas
pQSTB0u3I9wmvGCMBG3lv+YunUOPAyfWfCE76gtvW8LVWqqOIMs2jxZmIvfAnrk9
oO9N/a9DrKqgFYqTJPleHkylRASek/1n4ZcBLOoS1GbV6n/vGYi+7zF3qneJfiiB
1TDzDdhJ5yvviBtDBcmv9cTsO/40D3stUMHRs71CAL1/wk8LxkG00gUknpev+0tL
DgP/pQzTgJdsKxraC61DrqlOu0JNJWNKxjIqIhSUZwhdTptpuRxrDdsGAB+sdobg
c6MmpzwvrdOOXC1Gm83aaFTpi+TKGzMvG1eNO3Ya/MiRRlQCCxOMFaM/HofpdhN/
kd/uOYs6iJxNVMTQMoP2DN6UTTTNK1SV6LN058+ClyIdQLlkdW3Giil8q6byhov/
AQ7mjls1QWGILSooOJjEjt39z8aZG74FZGJ8dPoXMPV46EGBererzpU4uj4Qqb3E
UW85m+LunQ08wWoVi0YfQnK0bKOb6u5wYtDa3vYcW/kaohMZug1J7Zwrtl5EjXzc
3gfkevn5fYgoDAYSfP2baWDjjIb8nImJDoe501Ean8LRqOH11s0Jl+4OJVx7CjU+
KiBY+oPUWKv/Ix6M8tD16+7b25cWV+68hMMffO0G9aA+lpf271Rnh38wv5GpvTDt
+YcVTCHBm85LPppv0tXygYzNQaEJcJkFWwTBY0iAue6/Gl7y7QU2xf3tbL7tYmKq
8nVvqgZuYo9xQ9Ck818Wy9ZQwNmlRC9l+AE4pkFDlCQLCkXl7uXd18OGhhUmxf6U
xIHz/aUDbIpeRmZ7rYInJGAnZvpxKlWSmIUnu6vIZH/fW2a9LxCq/ho/mzO57nNT
t5Zw5l50oT5Wu0YycSJnb1BswOWXrm4RPq115MtyU85vmttAKwtaFpWvrkW91tlN
t+JIlXwII1Rq2AUWlBSsF8lTS4hJLa1pZ/a611QpqAB9whCs+GCzPNXdMHPX4Lkq
aYcS2RZGWMK9AF7KCIqEwb2A0r4ZSnTj/X2yPwhhSVtYpnbVW79XX/4uss+v2pD7
FPGgaRm0GDaIuysuZzATnPgK9u0SO92r9vqUIUs38N4bIZAUbhwQWc4eKv/XaYnK
dbyFVf229nxYstuy5FN4cAQQkMn3QtO1QzjHuDoZYfaWD9Z4JaLMcMeorGKEMH/L
2L9jw24cprbrkJeXqjd4A927ZRW+t6fuWT2bh8JZ1PplCSdFf+C9LmaQ2JtKWdUs
sGrnPXUoBFXU3tKGWwkHkeu/d+3Q2DKvVkl27K+orlzP95f+M8i8nVmfZoDT5mwo
dL/D8z+GZLj4srCW7rwJ5jDbi9DLIJ3/4XfqbYUL+wXbOlg9UgjIW/Dg9b8V8xWZ
3nmnBrh5W/pIvWMZsET4BP/OOXjbfHIPGnkqVJ2L3ARFC9p04O1sq4PmEbi5TVdJ
CxGmOhC6+f82tA/9lPPzfy741/CnQSmMU2R5EhBSVyab8TH3Zzm/FK8wvR2F/pqR
2d2Q+odW9SpN7a9fd7ffcd+d+KUxF1ff7YPnqCQvPh+I5AEjCKUESlF3kLNrMSAh
k1rEbDZE7RQfjA44+PrgtWtgEpE1OpI8HZqPC0ZG8kKktiSIjNNHcRFF/I1gnZV2
4bsDSHclC+Vv8zUoN1YHln5GxIuhJ/fbJZpdNFhxYhhtJB52+DUs4NicpAalKuhT
uKBXVV4HQydxav6nbEdJ4gQNbqK8NqtPMSPI/QZn+FBG5xQKrYN4IsGk7kJ1GMHy
Fo1SzO0z4fw/RK+gXDtDS477YD3qMAnGnbu7NVXoQAT/U0+Ls84iJsPI0dAW37Zw
YYK8wQ2cBTkve9nPW+S/Wt8IYiQsn/EGv7TwqzaFH23qpY1kHi/LTzlunZcBWW3X
j4Tb8sw/0QMhBT7ZpqjPXPT9v+6fDU3rQ2C+D1ToCj8VvsH4BX8wUoOvb3JNbgMR
Y0pUZfN3iyKZqnVoSfXWhT2LybeiLfSi19HW0rBaGpVCFsdlg95cmDptpIT+6GMH
UNwKh9za3AiLLObENc1BlO4RmwrMsHPQjPy4Yvp5Fx0fLWNUahDxjLEvgybI/KAb
X9cL3siNqt6k8oUPeSCpMGoP0NVwa91qbgrsWzprfpTGHVAFOCocQ+6TaS13geJK
fnQ93q8ICYz4ePW2dmEiVpPA0MHeqCZUW/RQ4Glbc2dyRHo9pE0RvmUbZlWhW5G/
zFGZwIai43jqEEoUQVptB6KeVE3PSwoTS6FkcqGduSam4VBK5GK3lZ5LfUUkAdvG
+6528JM7YrHtQH0aDHzPq4vGZAcyhpSaw1hENVn1ezyL2v7ji/2VmUKgP5S8tqOE
tJlarexzX6TjAm8WnsxkwQf53p4fsu4L35FJFK34wMW+5FRqfg1KKUNHUAwGfBcX
F1G/1vQe5FFH3S8LaI2FDo+/khNDBO2ZICW5xGN+GY8JhuR3aqyeycugYjPdEpjp
zvrCpxvbsCzN7VnXpf7mi8aP4Gbx2oMZyC0IBxMetndDgWMn9nsoyizX28rbX0YV
WzOl4gf+VT6LmKbwXKNX2hHn2E1j8K7PaAth8A6wUSGG8RPOF2I0MBRuqkVTQh0v
Lep2XH3vXj3vGTRcCEBblAGh7qVb/ynHYkwBrzDoqMUItDjNJM/7oEXfBbiI8WJn
A5qKhxlAZfE4S43xMyg8v67Zh8QdTOlRqKR+cpGZuKsqGPCoCwqe0TyALreVfZMY
H+OUs8/U0RqWEMDuN3WUy6deiT7oh795P09PeRNhPssI3dz1Xd8rmmv/7k+pG5J+
zEE91hmfSiB8BTnRKROWTlEAjsBG5AIybITWXSC3WJJS4GtQns34w+e4zGl1SvSa
TD7fyoNCtkzqd9/aQVtxqv2tXcO4dalmSUEgZ5rBJg8A1/ksufSrEFGnYAWmGI8a
RfvGb2XT5OwJyHQxFlxe3paehX2XL1MwKlqWwHcfn1Q1gTXHx9uvARVOdyjLLfml
UWze820aM89DzPfdExcSxnjuJj4xGNudVq5e/fGBylnvcGojspZyCGEFjuhGfJfi
W7Et6ILKpLSSqqbhvwUCUIYxgTWsiS/5s6NFlOAbhcA86oJmXrdhG3eDKbgyoQrW
A6j3BvPnLIqKwzYcVj/FaM05GzBXZ8nPLv2KNOl67l1WhRzyslpIHHCw3E5RqVsF
s37PGNDB4pZoWRwl+q4ARlyVP28SsWsfEMZv0biLU2d+vjvi95mCCzr0MdPnFjO9
qUqZC9UxqJ+1CDYYqIg8/rdx2s2r4hKYZPQnwHMt6N96XW/pqfwD4afqNWYOlEVn
98iAcC8ri9x+tRGYDjkPrZY6wi3CpbMO0O2ev13sUuOSpOnffLi3WC9F6ImzQ9R2
rryY9DKS/e8BjU8bM/DozEY4lun2+Y5r7xvVoAem4TaOZuoUOOulu3nYpFUd8Ng6
xQyyeI2gOgQJVgMB/4ujyApbgkeNr6Q5oROcFgR3JSqDV8v99RKbiw24VGBM1Zth
EBX2a1VGG9e5ZNQ7NobllubuGbp27TIMStVntnd42snUI1Nu3E95WEKEU/ebcERr
n1TQFIyHyIu1KKIxpJFesLHae29n/7K5Li5JyfWQC1cwE5aMGuO7dnRK3SvVs3vA
oqMGM2RUo+mEivzV1J7e6Yqe5AvRnnLMNzMXAkZOwXs280F7BO8z5gtxPna29upX
fT91maCfwMRhPTNWUYoBxlJzXSMS4Oq4tfKHtjsljogKcA7IWgK2J2/kscAQblXO
zaedW/xOu6zd7/qm9PwmlXLid6maW66vsiPKLNVa41n7yTnuBPmgTU+d3jz9vTpx
1fK7H8r2PmqfS5NvbEp+DahZ6RRJ/kqd+NGu07IUcYD5zW94fmStme9w7FU3EvN8
aW6merrBY4Ugtb27zlKAfp1OzjkO5DWyvtsT14Z/+JvCVO4WkcOT5fnZ6ZC/1PAU
r8lP1Gin4OMc0tGNLMZumPdS8PIL4Kysxz4xA3bd4NeJgsrsUwSf17d0CyQqXTbw
HPUwQ1v7p3aEt84ZZ3L0ul0bRmOYNdNg00153IJ99fgwDIWyetytKfS/rfCiR3Bj
T+Rd4eWJ9UvIT7/P3GaQ7QQ/8PnSKl67/HkWnH2t6912s7L8+o9wW75wFFWIUqxQ
uqmYpaS3KAeZjVgv/zU7t+n2v6iOADu9IGUSHdSfJZXANhpCDbvFiktYscNy97ES
kfUn2EMg7mvvfpNpsgXkMjIFhD5N+MfaVI7G25WF5mxt3AP6l9zf5JznnUkuOzaP
9VXA1BUKdpvyPLaDMwN7beTZSvNojWjGkru4N3FQz8xO7UojjDwxX2sG+rroEoyX
1Gw0wlwTqLFlUAAGd5BycZKjsEnhozCINSv3oQqJofC9teBylQTgEpOmlvtXgtJe
K2kJdsBlW43WrTmBXG+ML44coxxpqDcTyNue8myvYzVXQFIPtGJ5zmMwOja8kXuL
KeQ6pJe34pKYoX/ecNMIqS3nVH/NrdtpVfji8FF1qxx5952PCmGkWfrm0a7Mo+RY
b4Bthv6tpfUg2j3L5B/G5BXTTlEbbi+O/Xkq71BkXe6RlPhyGAPClTMJgKOzSMXQ
qSUoYygKaVNMmvfdD4Xj+ebKD+9meI/J7X61sFMwrTSGmS7nWinDu94QOTHY+GBv
oZRfaV3iIRPXlMV6e7nEBKfYh3HmoX7p6fO0l42fYCwft58k+AFZ82EXlkjip2l6
Gl2LRrEX9CIzbKxH+Y7tArOsskrcsHAbXMraQTyyw22TDR4TYJXvru5e3x0xcUQL
hjTHt34cxfiusGcy4Sm5EC81AUThL8/TFMYmwioYNiuxivmWVUu2ajKp+/lWlWqr
ZvMRXpOxTLryzgdH6nEKWB+kfVTXgdb2FAehFFKHB1s+vgXFnHZLYY6KGMp1VHnM
TAgcA1XQPLj4ZaCZHj3zFc8XTICj8gGzXp2ogPGweMtclzE3BLvPo2YVHuPnvjlO
o3YuwfBstkSqZXEJJ/CF5MxsvUD+lhTLmD3ZB0z88KVF9yWitKebopxV2eifk/rV
wm1y/8PVtVlLkSZIybmM9f3BJWV5uzehcEPd2hlFT/drU/jK9QP9hEJfXiQ2/h9y
ooYXNaqK5K6//E+9DIP+V30JfQj9rp+pcdKMhY3fR1rL/PMcqlCEJOuBCfay8nG/
g2ORcHFsVP7JQ+1r+N4AC9SA492rI0PEtcQ8Ui95/MTJ1IX1jCu9rr5pxDGy9DHp
02bMtlFNrLbWPap1Xz0Z/3Hz+sJ8S++hweEAxgN7oNI+HkQ50HdQll15IJNSKZXF
Lb3OfKimBQh6pL3C3XzEZm3iG7S8wMg5nxzCVKPmcSwz07RvlZajToCqsRcMmkwF
SlEEZtiPUff4tSK1EMfakBVyKZk/1ucXZAZHPewyiflB596Fg5FNWePPDxi97dL5
7P7gamMv0ZimmNGbXnbz9njqvLo4H940OOtR4njGu/03ZS0rlTGhNt8w1nP+AOwz
TpnyrAUSGVG+qw1oZK5L3tv6FcanfWv9+ZIKuCE7LBZEpijrHG1A2Y8Nr4CHcKTK
BS/gs+vxIJ5I3J3zPYsbDt1cwp8C7olYRWq/GGZxu+stK/mOU3AeJh+u5vkslof4
JXcmJB6AJIxRHhfDwUnz9OzVVijdfeWt0CEYkj1mdUH/BPT0sZ2QXYsjN2hyRvDA
t7UAyoVpUuxAbV4HFFb3H5uBSYBnvZ+J/uL9cfxwzBkEw9f5yUeBSkFrPKIZ/UcH
C5MT7kyVRk042jWDtW4bA4ilwNCUrqO6PTD7KjvdhyfWYjykbi12pbduTfOLZdBH
MOiqxkq6GDEHu1rO6mrhFrVgrpFB1JZ3E/un/2RKYRoftLrZVNop/uWz+QPp9o2T
Tu6lI4uZdasfoORFL5l4kXXOmzHLGZ8XretjOfPfQwO6jRGzQVA4GCBJq72hAvPR
u47xlvRURoafNgjSxw9umeG+rJqJpuGqSk1RptZTe8exZEQbftDvDoV66vhLCil2
sAv1awtUxopoYU8kQXsME+lHvNTiC7nHrUT8r3NkpQ0GCqjBE/oMOXo5tVEDUSV0
a6y2Gb5lXqZBlRouW4SQYLztc8Ql/EWYziHOJR86i/60fe+Oanl0htAlf9WsW1Sy
eDj8uKnR3i6ocmXujLthw1vDJfSzXO/GO/GIAnTMn5eRHRww3+v5mqYl1AMmq7W2
ZE8YpYyRqF8vZx3Jvd/6hJSlQGmPIXBHqaxDk5Op8WQ8G6FW5mcE/PFHcCjdpyYv
BEIJ3FIPsC6JF9ySylUDSEjGeIa+8FO2kITdWbnvq60kYh6ll9mmFcQD2VjOPIXB
MJHhrKtTjMifBYbAj2WrP22eJzeWXAlrWPcOd4sa5rylZBLyOIMFqgVB77kxlHVW
l274Xx8+KdVPP+gIYVIFQNqgvpbzP11vQYRSAH8IiE/JjiLBcVhsUzsjFgr/94aQ
0ySf7mHHQq3Ord5RIaixrpB4it87GzZesui4ceimV1vL0NdofNeFmdWaAJlQ6ddJ
pDiynL5wMUsQRe7RP/A+Jupfc/fmY2HiJ+m16WXAKJ8duhwbAYC3/GOssSz+vaa8
0xvcpS4jgcGGx9IbW36zFwiBt7ttRLV1nG6XfIiBIICZkPOPG3PLZQE5UlGCc0x5
GVKFbF9Wl3fA+wR2CaPO7sUVbRpTuE8l0XJODIzyj/6tqq7E+ruLfCnHf6slIP8p
fLJ7ulezf6PoED4tBUMrMcERSHREaSmiNPDeIXTJcflLawGAOXGUmmeEzO5bYzSJ
0xnhstL7qHOm11Sw5Q9wr6DV2QE/zPK1dItwKK4CKC+M2FYnzHxjSaW4KCOfzfj8
lT8yIWGMN/jJuMUtEMHQpxu7SY4WgyrwhVOOufgXhM4621janLHcGqRWJhsN5n/R
GoTGk/DRD0OFSqONm5N0wCi922Ks7kCrxtrawpNF849WWoLlAlw166BKU0Hs8deK
Aoxx3FMc3aEeL1/Geg5GFf41lR0u+W7ii2dT79m2+2uo7KskYoE/cIPCGJod+DWc
J4wvGSDpKCDydw+ae62IYmHY8ly80wgN8WI6w00psFPzzaANbuksqHA6d9WbB04e
kqpWNtFyEY6i7NfO8VdV/S3Sp7J8GTpemKdIpYq0U14+rHCFC4d1TfFuXOVIsLYo
nUYgHI+GEyd7dJMjyhMG0u6DcRm1oL74/AJOicI3D4e5YtcE81xKNLs0IvUYJxqS
zbJ4unllPhazRRP7W4c6/NEN5sjbfi5DfhxemmIXAlI=
`pragma protect end_protected
