// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mPGYaAB/ODGPjRLwWx8qMtnB4QDej/HmsrUXW8dh7wbAsk2i5ba7ZySAlJnCNGuI
GIx87yxLKY06986dtaZq7Zgl+AoNT+7f1XKABFe3dyCHCGbaigGA4WEuIQLCkbzv
v7oSszBqDHWB5XD60UgyHDUkdtroVK9pxVQDnJo375U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5200)
6HVdEqt0N8MGZsNGLbFnXrBNDz2U3ZGRN3a+cNfyAOdCVSo3qOFeMmoj5qfD/ECC
hL9H6hec8uYg4VCPGUX9xBwMGRxO9yGQl00wheMzYADI6FEFAIkYaMgS5fxPQGmW
Bh+ZopdjRnyzaDtOewNEHeWPUIK07oRx5BoG4ukWrvVvQ8W03jH94Vj04uSxQf6T
BSOMumVPoY52YCtbBcTAwo3L7M29Ne1Uw7STGIb+D2gaMY7mMn6C8QMWUnbvfl6F
CIRAZ6ynR+T7fRqy5B303yrFCvwRzMJJRBO6c2TEEGiAkKFNeOR2ykdkPf16NOas
RrZSy3fcaQjUpgV1P9Tr4X1iACXwQPDEMerVggCApCKkR8bpblwIVZXGGw7/CMjz
a4SPvtZb4tdQ6WKepMFvxA3jaFu80qhfY/zUKSEXZOKh/nvl+Sv/c2iH5EsXID+e
kqczDAnuuLr3K2Q0fBIxxiLghPtlWrIwGVH9hmvALfWiJ4w1BwBNLPl+HtlHyDWL
dktQr3GJtdmwYwC/KILle3fPwyacjRXrLIi7oBIotCgp/jp0sKYy9h380Dg4xjS2
mB5kC3mUOsuuugDhK6eZ7f+0r2CpRrLYCrmzo+aACIZ1nfQosr2/tQjKbdcS8hCC
7VCRxqZkyidwZyC9coJP9OO8PiElvL/IOBThsv8uO7FaoUU4/6uiPGS0IgmdpfNF
UJ4xu2ho+iQBfDKflaoI6xaWgBKpyuNHfmc6F1m7GBRGBEBaFV8jwIFSEa2JyFLu
SoXZfZ1sOuF9wgxLYbd9jTzu9OfSDT8cxjRvVuO099XVbGiS8wO02zvI/5VuLmUy
hwaVRrYtLjLYMt146fQ7TePWeFSoKa2RdyNX1pOw+ZwMjBsSCO5Z/QEVcJ2GyyQ1
Wl603SIonokqIubr+c5T/rl5XwtKsoT5GocqsJyMXd66nqNhyhSG9J9VkF6ILHKh
3WJHsbKBp18M5fzE8dy/3IIUbr9Y5OS9rlUkJYj+pP65wnVwwMKPeXrlQnNQDehS
4dBXTdPX74/oVUyf71+7Ma5b+7pJQVK5nvzBO0CrBUlKMnth3XnRjY7vZL3EhfB4
/ildDw9LCAl9u7m4BhKtWQ9NNp1IL6SAWz6ss+pcc9qcdo1d4UnK/7UXknxWNpe1
aYV7INODxvqvx4wMsN+hzKlxOkkYKoMorPJqMYXz8+ZXRckDxVrbIrXY2WmSNuW0
RdzVfsxL0DV8SxZ9A9I+5AbUfFkgd+m5IpWA3CH3SVGEEs+WpagzpHHr6pFnmb3g
38BrI1XjnLOkfyUcE65ZM3C4vz+p4wTI3EsJvQP+eq/6gNwR1kJHjjhE9kfSuyMd
r3uNdO9XjEWIVY/gBQX7u9F0I2BghN/Wf3oMJu649Hht6oXeuG/l5+bzkOqxK5X5
2peekNEXfxhYeqz4QPY2LEpzvUl/8tn2TXxLbmdE+wt/G23zqarve4K9+8wmJpJI
KUWWxSoZVSnzswPoz9XFX0BD9jmakJaVYx45rYX1ZCUtPLraIaHRlQ+pIyrbCO3s
vbpxDM2fK1sHLyoGbFOS7CDgZrVvvuuO3YfPcJorRcCXBm2YdZEpNlA53BqLVh6R
2SkEA8mjkrC3EW1lgru/LBpRcs0nwWwj73A+6OI1rsc2zSopfCgwQZKQDu92+bl0
fNFABLsX1OATYSmYgZ5C7hV5Wunnjw3H63Wvo9UAQ32KwrTz2CLBBQsK7CxyHimx
MQmg4kCqmYyKezuKupjOaNPTN9M4S4s61RUAVq681uxhqlZ0KMo5Y+cqiA1GM50G
RDomKhn3zyBJboYnWRN4+GCwV0P8iL5pUCm4IvZR2dEUGpJCeWjp3WnnmbjPC7AR
hB5YPWGJXj0sklMW3jnTe/gbv7z5UJwqCeXGcLa02ZsdSqGo1rkWfOnI+bM/VYk+
oqGvTJB5VcwQnHkLigZYcDtmCWg7T5jrMCASv5Nz1bgZiJqSIKT2IPG0ZOumddCq
W42hLCJPIecN5fm9GbFcP9sRJ/6fXT/qzDmgifSK8dm1hmaPLGvf3h4VjbvYXEY8
hV63sgvRUOsGqky06+wBfxvfuhwhVV6/k/81pEGQoj/DD5kgOwkjItLr9TTpfc02
j+EdO5JXROlgzqouY9hONrEw1kl4spibyZvnJfPtZTejR6FXzVzgdeLINnZArFcg
3InhaU6po7Aog++JToAqy0BLS38lfXaqy8vix2d9PFi4EKfdu7kCSDQU8xGMGSZK
MDnBtILsJNRkqBp3/8Tc30NyOGpoCU++0PkVuNpg2IBZwLlwe2fB6+PRu4t8Hjcg
NTdHlrz4GxNZn+SW40R1UnYXknwol/qkQeJalAQv9KSWbQnMpUBx9sYiJyKzAh2Z
je54T6x6plDjZ+I0/mRbe90fV+c7u5ApXy4OybriOAlASy2QAwnfYyyX3cehybLA
7MVTDl6V2w8cBCCnzFtvNCfvZ8DWTLfjvGwpFzDFO1ZWmT9KgxNTuvadB80uHtPL
XXKp5YjwP2UuDyokZhB5LPJOgZWE8patYSFPfNQ6CbImiKvVy+bfjYZ6rUWTAPi9
vUmH3DJd1n4l96lqJ5UBj2e1VtWEi2U/teXajADsXbqaniRzi3GOI2SraufbxWxo
TvZTV+ua0G5pRLz/o8CT+D5Njhk1s9XzSx710ws69Tq4pYqYxS1EMeCBpWS3OKHE
hTpzoCo2SOqlwHE5/GJ9/W2dLs0GLryLNavdSDFqmO7Hooz6H/l3mpbxqOYkNX5R
cSCjN0uuvA6RBsjTc4mVZZ0UKgpwyedb7fBEKGUDxlznXUYJWkX39VnlpcUE99Ap
B67RKPsnO0nohdsq3fwa7v6Esawz2F/qmljDM7/BMgnklsa0suAPrDE/gk9XnQuM
eAAa3BFiToy98RrBuMnz1gFakWCJ8CdIY+9RVznS/kWhflwS0f5GVynH4Meampni
r0EyPxNuRLh4ACKDARETHaazMzn6RoXOJJiU7ZOSITb2RHez4iaeFz5XsHqj5KNz
GMmTQDCTGlWeKHo4P16oREv4MQtoULAv1hagSYlP2XIHW7HUaVHFm9VmlEKsYKhE
7Ki8X21TQURTGwY6Wf1kwuoa8MCyGadt6GCd3CwklzK/65PrisDQBmZJFz3dEHZT
O1ssYlvTfQBkcSx4tkD9BC+SihWqdtZOJfn3UU3zcw7EVRXBDGYE3WoJnmnEVGYs
NY6MQ58HWHU8rBl8wQWKheUQF9v90OvftQzamJXocTIe2JNe4xzBnxwVJzswpCH+
bSq/D6kTYZFRbPGnXezDoCM9qpv6SuHp7stp8LDQRGMC2931zQuFHb+HYQVTnTXu
KkWhy6Czzp/XXRJhm+V/pnwIuBVkEzg26npDlCFTjsw6M1kwTSw3d66AzQIB4iy4
3ghp9UotIHYu7UQUQxBwlwOlMHyBeotbk89zLGtjmkIQX3OXEoLgxkjVCUUbmDIH
ddFFUC5K5MTVr8ckAJsdADTaMISQloK54zjHpA1rFoPM0v8geFL84W7FbXpgghag
aF9oSjOWKDOk7+O5S3q4XoUmQ1/LS7gD8bfPBrp7Zumzltg/8FSyYiRgmagLpz6F
SWxs52j7XZJuKwzM8PAqsrZNkedYD0VRqJg1GiE6FSJ+PXAXrYK2j24mRzMlsS0F
KX8uR3UL91Vb4yj6ApguebM9hldY0r2XRJ+ymNkNHCSVf9CC91JSgu7M6dg+2x8s
iJQ9dE3dF17n93425XZjy8IRdyJZDvsxHk2fi7kOqMAJtcFB+4a6sco+eJdZ/+AT
yOq3Yl8WYbbG9fQ+Q5zIV1NAT655T2vKkDT2isr+5jbi1oTUUPYBLig+UgA/Wntj
gM6IWjZDji+R2sxmj5FjVRZkOsKw1Vvb7S3eaHhyJD0J8d7uSvmiFim65KZ8GK+U
3JlfX1dGo41+c8MYHM3OEm8MzfOIpNN9gVXgq51dgbnlAB/El6UGONSO/k0ZSDvD
rnek0CFOfeyZsDdYa2AeO9V37wgIQQM4DKR0IBCsqDq+c0zG76R672ooJmh5cSAU
76BbalSL/vQA/+DvsR8CvKHZysL2RlHAgOpbcsTE5KajV+Z2r1oMN3FNaizuC259
VyDo8REObJqDr068GgcNhhs+Qp9JRgt3cSxCT1wBkevfOZfNx4g35DRsR6b8gMQo
jyh+hkfc46X4r2LpoPzu1wpAnr5nu5tOZGnmK+Y1axciexMe7silcFFSXgQzYVlZ
YQ3WOnGJkwxi5BrGX6yrpcKqDUNZFK0tD05Qc4VfR4/1s50Ep7FvvAgcV/Syxlk2
4gmbLZVBZnyx/6y1S6eRvstz75oBRZKEXw2Memv+lGrLEFRGx5t+IRlAH3VjcD9w
dlgImuMGkfeD4uFFMXVzf1Q62ZYSAIBgmMTTNz3LavrN5sIkFwnjEfiSF+Heyy35
0SPFusQtVubLSl/a1YRvKJ5MIIRnqJ5Y2jrMIgUvkAXWk15fgY6HVFYGnuTAqmtU
ScjSOBjC5IKLbnWIp5hbPuK4kVqPJyonZO2kPVlgDpYc2NfEcLPi/NhjYF/ShuCl
roTZ9NAvqnjuOVypNGEjtv632WVfLWlvCn2YfitWUqLZCIxQQ+KBFfu8fYHtOlVj
XketcwZysCK5LhP6t3nJ8l/d/VHIUDr6thfzb3CvkdaVV83WYV+AH5FTylgVJLSJ
gAxm7EQSo7pmd8/8dZ4sh4nbKv53oF71D3orCCbbN8gECHSiBBgPCWkoSCzqzFjQ
mCp/LY2mOUt5Yp3thVvcoxoS6I1hShG3UFznIvP5XH3k0aHbcwyYX6kiApEsXkd7
cmXaq+0auMm7x3i+viOORcr4kybRqFn9zZYeTnOrpZ4pmBQQX1WICNZih/i7tMz3
XHj0Ue45MBWSY/8WivnisQPsJvuTV+tbHvGgMLY4By0zlRYngNPn6X1so8cHsS3a
uvWxxUCPZQURQL8RBEXNdTLNrGxNgY08EIzTUNP0Z4LWI56RKeKhePUdz0y3/eba
OZvKGB0PoBg1GEmx+Ng//E2POXJ7MoLZZmjn1wx9St9j8E8f5owGhPYXqolEA1bw
ZRzG8L8qB1BwmxhpWQ5Vzs63LH6xaGN8rAz3S+TOVyWQtJXwctDv9+2n8nOm6tVq
JsS9IRoMfXJ7iYNlY/W35PENiETX/YcSD/m2b3LCDOlJ/cqqR5dsven/qqU8vJBk
IHIz5ueqzXlCZ39z98dwClOjEYJLUVvrOovfZ+GOCodRvbrjL1TNOWCaO8z2G2GF
01tngyNwgIH030QjBNhXuj1Wf3QbcVmvXPdFw6kTZDTcMvHBw2lBAy+TdVTqCmFD
+bxUnXcvhSROnb2cCvGnbn2Z0Ajl8imbbXep1gUIX/5GVM8b9KshyNeAoKny0GEr
z9g+7wbBAo5KA3KMoFTL+qNDhAHmZf4iyU3srWVYM0FbfXY98XiSg6LEKs5rZRn8
AjS0/3qRYA1s0Uz/Ww6JQrrMFDV3yds8cub/YvF+LculRALB7UwZVzvvLynSsEGu
7SvVg5l2n9n99XRTSOVOChvAlbbfdWGiZ/OWSfkqtHx6Dfsm40VerjMt3H0KArRJ
UYTOXUBbkcwaymHsELSDXVSMOdSQzx6qF/8w80ySHVvUTXbmvQb9UxUAP5xgIjZk
hkuSiCFUw12whugUs6zJYr1FIbjZemtE86CUpdcx95hX5t1zoaV7nye9vYxQofue
LiTDK9aSMgcIua44bcaHMGbXyg1GB7oT3PZSpgcp+I7erZha6oQm7CJFsNPgmizJ
AbZkSTgKXBYvXCPSkNVwfy5ZDPDDbDfwzWnU8FcajYVlNGOrk/DjW3o5jnOMB70E
nCQ7l1smfUF3TGis3O8HmXMkQPcnh7pA21mcd8fYUZRBK2LKWyPL5pDERPZNk0Fc
1o09BQuolN79eP3vWzVi7DdA5dTt9+cNnpdYoNn46+tXLr/8cwz2iROqDI7hLidj
zDgIYsbHw3wR94L8sHGZ/BOKmuB4VW2eElzX8LZFdkiUmUU+NQbg69X4ZjwfEFUa
ON0NWfE1Gr7SaTWw3EkGjVMtNKgtfPHzSBirEIlfSsAdCe+lbyy+kdTpyjW9bO3Z
zuP8RTgOz0HJ1pToARRwVmjEpnnHUVDn4GTNmayql5opzx3bwHABDoNYGc3pC9Vx
wvwX6HbSXzPT98JKDe5hHSu2jTy0a57zAaWJJApdR7Meu2aXAiRcv30NomSKQdom
RbU9cHLju22YruhD0D8pkfLXPnSqbV8n7/TMcjOpjp9lwNhk7sCehkSNK3XE6zI2
jvWMzCcytEKH2bqJdccW/vHMMp2o9qctuhdgaF9zGBFZ0fF586nMqFRzfUjuH4Iy
X1lkLWMR2h8Gl0YOXsE8ZsB48DBEULPdi7F6ctucmpj5L9nboD/VIG4JQmVErAs0
p5Nc7tTW/Wps4wbk6gTbZTBvdVLtaLYcDO607daoLEAu344D397MviH3dh6boFdc
S3bTgJWTeygjo1IqRE2uS5bBVqtivBVrK1rHS5JRoO2OclCmFajvBlqdQtschXr1
jX3n6fY3mWP50rKYKLCaeFOg9QroaPkb++gQlp1iU2GQDXcRfwzrTkwCPvGbURDd
OXVYOnHCoKDbEceuirBLZs0bcbLqmjJbzxzZpFbGXhMhDBDFGc1Yh3cxRNsEBAMV
ZgEoEF1wLgjpX8K3ejlkhmVBSiQ4wb/ht//QyDyczdnJ0i9wUWH6uUpi5436Ka47
G0yokW2q3XyYbl7QVIcJBieSGNOFQuAXEbjcWQuKTCU4oKWDTDprljurUED6o/2N
9ChIuFzLRaTArY0UvlNp5gVePDzX/cII9eus7+Nuz6N1OfWiF3xeMnLyVvHk6JAO
2s5LCZYZNc2PZMnlHsjCayXUgzoKc6IWIlFi+vnSR+tsQOD7ihCRZPMCakNEfNxG
Pa8P6Sv/PzDFslVJTt9bPw==
`pragma protect end_protected
