// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KSKKrXenrCnz07sl41eZbeq2BgFN4Y+6lEndKvO7yAn9c9K52e99UOvjNddGo9Xd
GuV8rRFvktRHNO/b+7NKMCleA97JZaR9pqkQIkE1tE9VCOO+CoGBE52Ov9+/WwRB
YoLPdjmcw5rBFE7SuwXhRqfi5ew3tTjcU/JupeQeI+c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4016)
fwY2LLD6HW4VXGphzdoc6I6eG90OZXu7EjfFdUzDAooWtoHDm6WIdUHwCE3Qxdgq
XE32ux/N7w1HimosZayEM8yeq+zKKLHNmfRBmMyhKV4FLYs7oz9uyVMFDmwOO/PR
9uwJbSI5cXucmVM+lk4M8e5IWvQ7KZ46MnCGwIoZYTcWeKQk3eL9MeDKx6736yjY
0PlCr2dEHjACAdBJdKEWa5cjGQ54SgReQLVp2Ay0UY3dJoq7y2H4f3UsK9hgA1Gg
O3psrTvpB/HzsYuLoN5qSTeIdn/Z2oUsBrPWHmwE7kFnpSgiCT2SZAk/Zcxq+T9+
qDu8rAESPGkcm4FmDyJAdQCoZfVYsMBRLIKWcx9SW0jcpUNrboRmCofOuTFvH249
l9F/WytWgCDlJIsiOl9Ecv+/0MRkh/v2xur1A8oBjAV8kB6ZBDpWmFrnOtgNf/zw
SE7lGN2U8GZKM5jeOrvQXHgFSTDVryKoQ0vpOs0wXhwyzTWvnV4wnUt494IFsbk5
ykSjIDQjzMVuOysAoJEUNOTz5F1286nYXgH99sd9AOZstCGUmRsoKJ9DhWgdcTbR
MqqTBsp3ZvyRPgBwlNSuYtlJNDWYRg4kjkBtd3bHLw7NxFdQTJyVrleWb/VW5eJ5
m5Zo29OAXx46jUPcp2L9OYN6ReWDnfIANJFtfNBgyeusJ1Ch/7HmkL8hcXPi+V+d
plid/PeEXd1RyXDS8pdBTG/Lk3DwFw/AbdRz/JysOYrFjeks0iQuw0BoRbrNPvyY
+mHcBlRKSHqTWED13DRG81c8peBwEoBCAAmnEvIV4rKNrdU245xNlb/K5lBuTOpl
St4lPPf/K11g9lZhBqhcUdVQ7IzpjM13Iz1+nMS9c0DSapDecNgWqfPfJUL0j6dG
tamSDGz0L1MVAJox/uKFwxVzUD1M2cUnIRFqRj4OufbIsW4kZYCcL8ZDkPAcHsgz
FxFv4Vp/y992c4GeYUL1HzDDI3MA9SD9XvbZVm1dagetMbyfo5uZp0Hc9JLEk5/J
+946G9vUsHU9pwAAxVTcZWo6egPA1+EL+BNNwCSYU9Rro6E34V2eYOoWMfy6YYT7
uw5UWgzZS9nGfexZIIAmZox8hRDOWjlyq7BXY1slql9lanyJo+9B4YV9vZ5Ifc73
L3oKIhn4MJTWNkqezTxLg8vJuKCQfUt9eFatZYExVb6Fl4B86s2YWlo/+1Le4onu
j/4BWZGdEFxmskreTQW5zGanGsbI7I1t0dF6bdtYNlEBYqvYoqWD4hlqSZXw/eZm
PYGy95ZTTZjaIqARVi5dwCyhDD1wRzgO0ut6C9Smu8PZjUIw+1h3qHOOsZUTXaTF
WQfnVVUEKbUzJ3UgmCAmVOlJOMVOb5pXNWVOijqXp0wEAwiMR1t6RnkO2ScqmY4q
RvMDHYd9mjpCW94K4T5degJg4eqJuvaCLaehICZJBnybrFJ0qFsjT2PtO4b+kc9p
p057KRJ6f+PaXUDNZKzpRCbDFJNWq6RIVW7Og6Gn1jouzGjrHv0Kz9G6AZTOcrdA
p77B60IWVs0ZSk++BtziQYevCydexuMPrtRgI+Nx1UqKaOvNbnZ43ZjBTUA4NhDC
ZhwFzKySckvoptfOPrugSjsvjvNo/fQtmmeLt66fnOTU+CicXF0AD+pGZ9o3ys1V
0l8/097iQq0uHZFlSBmHds4H1EngvlujytHty7UV1LTj0lqRJ0qdrQaUzqiwJ1OP
4PcJpod/meE6hWGBe4DSZu6eNQtzV7/E4dgZxZVeiUyb4YP3LnG4Q9qRWLVzO3/p
69y/750RRQynGxzftfVe1T6xLPMm3o+SV/Fpj0iLEfwYjCQ8cylO+Kbftg4fMf/N
dGOa3Qy/YQ/Ar3omqabdDEUsYBHovuQR5It5j6QWk3wOlFjpdWGqfn1BFNFdBbNT
rjlSq+WXB/y0oi6cVZiG/bRLi4pmT5fDJm8K35wyufeDw7ArkIHmH4cMnjT1i5zi
4IEJY1g+MRmtT/ax8F7YLjhoeQevZSMFpOT40DKRBd82gqebfmxy+BJjSv3l2X+e
y1rmOU4Tdb8XEYZDcZC3xRA1pny7gA7lJNge+zP7r6erje6nDee78YC+sM1bie5e
Huf1Hi7j+332e6qatwtew3A9JdNarR2Vnd3HCgX/j4KSnsDV7okpVDhov0NRYKbs
0Bl5SARh5g0qT7D50kElIHP9IOWRSQZp4p48UBpxSvC6gp5JVjjX5gOwGsCCYwIX
dCpNfJ4UEWKpKWwoSf7klIM1VXgKSQ/bVAB2ZxTdCW0AEAWEAxMy2UjIwTcEbKwD
UgBdg8jN1in7P4XVQJCvMebTiEcY3pNc88LeP9GDHKxWJzd44V4h5yEn+csmwYNc
7tL2zcZsxQhpMhk55WVlVfDKnqQmIzZr+nTm7Jxgp06Mpp1tHWlfTMBLwwHLlzll
+6N2BN+fgVs9wpPo3lwIlumSkhYMp73O6/cohhWFqOqdg+9w1LbG3ca7+CmHYB/C
byKHhs/O8Ue20VmeHqGPbBo2Sjza3xXAyDZae/tHuuYg5yYk6hVxBLbKTXzdWQkX
jiiYTfKmhfwYii7WmJzKLcCFAojvJ/aTKU+2CS8QwGqoAgTqRr3QRYcYa+c92wzE
4kKsB0+H7x4h5uoo05CTJlu6uAnfnsln6OgOAR+7oKcbpg0GDIAYxLSbAlzPVviE
slEGNYL78HWChXhnnzXIM14xbLxkqEiNvUYWS0zt4pzhhqfbyRBVy2EnoBvgMvak
kcvIASrgI7R98B+NBvKp1ZQlpwNoQt8eTYxch9ki+6k7za7lUZLRyCxtBLZ/X9Ja
vXjQLDTIqEOtWmY35/h6/VQ9Jl3wB7XcmJvMtUmtFUAn52oD3Jj9ooN59M5tQTH6
0CTSjHYoDQHaWXgTIHSPKK/SKb7pI1F9YT4OKbhtLWO7+r3lvVNBR3jp7ZIJl1ED
pB9MLJuprWSFjn7jQiz0nzGJE1Pe0+Jkg2PyNuwfubmLEvCzvr5EI1KVmcvmsHWA
J/oyHR8io3I+LduUHtpXf/GK+Pd+4Q70oNfseakY8ysyn4n3hEGKjaWUnSDzDQTm
5uuWnzeYyWGsqeMPcPGVgbzimgM8kBwPuwzNyTj5KfvoLuOrQJTw9uoniV9eSJ50
UOxydtPOV91tGdDi7uR0tH2iHR5lLjIZhHlbndBFATNG5TAfb5wC4lB6cC2Fp+sc
37fwGDfgaax3ZrAsQi+IQI5YO2YB+dNMPO2UFhBX0ClRV9yQuouVIZZUf5oOZITh
qqnO42CSUWu0PuBnkGPEaxEDWl/gED7/Rsjb9T36K5j092mHw3iI8eVyWMldl67f
kYiaP6+lOlMnMQFzm11gLnonLgWj3x++xAAfO+xNe91AJ6Jdq1E5tLUCf1MuhrTh
f0EFEWh8XrGKuOzbLXSncGHWT9ey8U2k10kXz9mgtuFpmFysD3uhd6JU73s8fyen
CtRThlnecRK64eesXUGbCdp+z+pAY27sCkZzKNu9ReqU32Aj2e2v0sUVC3z7T6MN
feQcSL3MRUoB0+Z2rfVN2KAzFYc2TnPCroHz/ioRK5wKb+ycVJxdjGhsKe2bZl+k
kpXUgyNdCYSP4kcCY0oinSHJfzgHIgCH9md2INXeI2fp16dwXFLw3DiikbKH5Wol
m6K2VFihQUuegPOtAOmdKXbmgh9M8wnSHGV8pPGZp507l3Y8arLoy8V1oW7yRqIi
PfZKzutQg6n0VUgpk9Z1qD5Mej8UfH734ajDxVx3zhL1qUy9XYYV/MioVDeR8pvi
OoFneq4cZnfKO21pCzUnMFfxDPY9Id7Yj2B6SSwjpzMFKl6F/MKXjsHy/C4rCmlj
9O1AWWo466ofNRrekL1+lcaDFnb/U97fy7NP+99ingK0XU/8eqw3DKyk9T9Jki89
KHtRtVZG2FkOM1hcz5Bxx4rGxLmMCOGKHzszggqW3BSfRsmaH/WtXZA9RrlTQ8L0
+NIPa5XqAnu9Nnq1c7m1y0wMYNg9JfdwwKl2Ahro5EBZecqGpV53uL9xY1yd7P0m
9EREzPfvAgX3yk7R/qMNlHly5TnnNVq1TjcsL/B7M2umcfrbXPQTJpq8k7BV7kbv
VMggUAcREEwama0nbxycqpTJmrdMmvreeMF/Dn3OMjyRrm8GlcFVhKRNjvUap7z3
VJll4bydOrG0BaWPKK8LUWfGTEn/qdP/66dbXhggVtFPqP4xCFoJxjgZB6UIpUxf
Et7geBV2egl2K+UCZezd9ja/BwrgNRLFc6C29VNKIX+HPn2OqU//+oWkeVggwa9h
KPjZZxfQOlplgtz59I1muxZhmVOFeGom/cys9NiACH/i/j37O4uXBLgqjAld4ATI
yVPemPPPbhpGBphEk36YhUWfJNWrxYeWxm3PXZEdaLdiQbmXTiYLAN4brrlvMIT+
omQzYh2VP20yy8mEFufX8pKd0XsPKx9YbCHJgwDAwOm5pkgdN+wI0N0Us6GbxNTR
0yyrgqaxcelKhUwUtG/ar2eLiX4DbfM4myiLwKALi0CHJHB3bnjKqh20LtnzVIKO
AMyu7vLlU+ovQQA7cc+ZKUj7kw8Hrt7eQ38rmBeo0bTMDTtXjHqM7tjCUhbNKY6y
uHR8VgKP73Raefdq5BIim+76itPMbjwWOtocPuzXLwgml2HnO8S01KV0cQty97RJ
dxtyb3l61Uje/JriMYcmxkAok965iPrWoNl5jvGTQmoiPnnZEwjhoIyzBxM59qVP
NenKxjAgf4FO2ZH160PLneWA9ladmgfZE2+rbejfaF6D5QG/ajZo3OqW78Ane2rs
ktR4+GHyxso938HR6rFT02JYxCR36KK8TCXTj16AAA9pMDKNVLcQW6FB+iEgJPOe
cMKM5ybOsgvFjeIbn+FnO1++391OWASrc6xQgIq69XB7rJ/1ztvcHM+vei8nTJp5
apVlK+OlCozyI75U+yzq7bZ6sk8dmGkf3TpbVso/gZCxhQjdjNzPj1X7KCywtd6P
is4L+3lMOz+GIiitLnngE27gWYM0Di5LUZl2RLMwFhK3PHo7ghWYJ9mOft+FbGgl
bLhlwotUmHk8h95d1l2Z1g+eGXmNaufzqRU4kyT9JdbMtCR7i14l3IMYCkjslRlI
BUxnciAgdps60D0cmYSwWkCIvyLvaVs6CNKX4/KB+Q7Qfs9exeiv2sIKr4VWmxWU
umLcg5/j8QcLnDYyOVNNiy9Eg8UZr1MbKIeZomD3ye7CcdSy3os+1FwjkCKx7z/O
GckvlX0m6OMU+7BmWZMq7hhTbO6Dd5B9tNeq25ohVYRuyB/fU+uTy4VCCFRkXxWp
As21gT9lvFBhLFsowwEd1V0+TZ2pLDFUomQP5rZ9qyM=
`pragma protect end_protected
