// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lV/WKybwR8fs9gCoWUylju5FHx8HdfSM0jVDeLXUBBkgzFkZ8QLoPonZYaoKOWhp
j2KVdGsipSuq6wWT+MEorGtdUVC/LAUffsfK6xmV2jp38JYqelbPqjNZUfTNR8jX
C57xBNUSUF44OfbT7ZXJQp4Uh+8iyRUH9Ti5EokNYXU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10064)
iF41bFI/I3zuDcpV7bVl+c8g3Wv9S4PhLBjoUrxL0kSquFl8L/GZN6jzE0lztv4J
SDMXrUAYr56zSgDU6uKMt2s0web00xpC3J0k4LYzlGXFPZjXWutud+rzQiBttMLC
wQHwd5R1kz9Xo70t1fvVoROwUvo9N3hRyp9xUrc8oDZTYPEE5H+TJgxwB/kM60Px
UH4DGcbNMC8ZI7MF+IH5ejjCRhC9MPLfE2OvKklMR/YAYJ+HUi1JgivSFkiDLmGQ
ZLeH7fGqSHiS1U/0HqN4aPfKVUtUBh4Dd3FRRT4kXBW92DwidiDq3zhJWD9ifTjs
t6mmNC+DVjrS3DG8IBTySHkVGVJ4DwhxWG+Xoji8H3OLo0f+7T2L1gDu81d0gXLc
/xku68Jai9pZNJEILx1JxC5O2KnB6GTHvUmvHBsXjxmNBEibewm1wT871/p8YYhp
ypfVHyMTFT/OHgNow9ahzMIT2oNFfUEM71U4Kd2IqhFkEVWCGU+2rVRLSdJmTVgM
cD1ApQw56ftosa+/71l0SpfnX4ZMm+PYxiLShD5fqsN0Vj4GBnkKubmZC5LUjjb0
g3NyyiPJZDjnFN4rgUtEiFstgph0hOVmOIpaP9g8t6pR7RANNa8WneYcmyTVJsjK
qpebydSZTtnTNNYZtW6PV8oE0cHdOEebExo0qHh9An5PqKlZaIW78ucPFS0ooa+R
p75Q+8s/yMhOOOfynPm0e5WS1FoBoSNAW0VcTwTeTma5sPd6sOGSDxrcQ9sA+pQY
zDZFIPiFrVWDoyql6dpWq+rGZ3MSDgzoHffkeLmZFFuMLJ2W80vGR8DQEV/FhZXX
JHFmdOx6R0uTLZDVAphYEBPpy0a6WzVgKjIyMby8IyFdLIIR9hfRdyb3/DvK6J7g
QVdgfFgqYT0LnMM35fIJ54kg/mmBg3bKK4dS5XvVTpSVAYo//nOWR95BM34LwVxX
P88n1Ziy/NU4LOKuw1MgRX9W0Yk+e7l3k6gI1pBrWd/KtfTv3o4A4MnqHHFReJT8
ILmUI1uRVV7gdytGrZJmT2PcZeDhsEHAD+HIhVnwpaals4TEirLTk0APqWlDNfYu
lfUeX0782KX2qPga4xvP3gS+aApEf8hQh5qgmFXsbucSFwNrFrU7SRIXXpn34YvN
VN6VEMbcVTZNR3t4GAX4Dz5aTT3U3bhpBwCs2EvAToF0fOOb7s6/DLwuKoH7eOMn
wLf9Luh0nZEa7QR0hPMqroRBBC75LmLnngnFOfDVEN605cZFc7jieE7hgIAYyXCf
YNUqSYtIXyzu1NiX9+j6NfC9/a2Z3X4A7pD4OzhY2YGTscpMm5dV1VQcMm8IPVNA
cfZ5WjyZkFdaPrDvrd1Oep40BBCvgEmFqAGT5mp0uoZ8C7h9U8sDq4GIgHu6+bLE
ZyT2LNBzCgr0hlqvbH6v63OcPwAuafQ5fBcLEspRoR6csZEp3glaUDbxss9L1t2B
bExPJcSJqUrUjVzdR+JZd2jOo5XPhTGy1WvRcxO0tRJyXOT+qKKKOzhR7hLpERmk
4dit7/jkPhYwEIV8GCslJMrq3wGSkhdvINXALLBxBklhFsh/ljRadp/GWaMTKi0l
SoViQ//911NUru9LBPUiH8Cm3dsmbg9onu4zyrXljOrHigbcNxiPio/qXGtvh3h4
D2RSG/qvzpkZu4Jj0cMXBbDUWvzXpmrTUCQDPNidu3Va4zliWtwY8vjhOLPRA8/h
hu+bYDID6SnzqspqIfFBl39VY+DIrQpy9gKveY/AKAhWVeJRmoC8s4DPrlVpAeHk
SsS6g/QJ/4VNtWyheDR5V7FzYuTzRV5E/2WDjjNv/mgoE8AGglaSMe45v7jGt7/S
DzJEFfEQUb6rSGe+MX7e2GuLO4Y0D+NJB4k5udD/o93h5blhbZoN+cj88rQP/1+G
DA8aHgoDIXWh2DPyg9AruKPizqTYZMjoVEZC+Z0MO/b3prue3tvtQZFwXSZ3ZOJU
KInsoZZufI0EemDARj4Pz5N68cwFKb9jFPr/j2m3NV6nd7MKxLN5GnhgTWd97Ep+
Pyx6/XoX/TYWMFfTbGw26Y0dzIu9mYQBZMZdKnQv8E1GJhi06SYecOozsrx8RxXA
6FOrut+ZvhD10yvrDfj9cdobhDefMiQeAeQwqt6DKBUmewQ9cgj+m7a/PmV3d9Cd
OosQlSqb0+koh+cn/+BM1arSFp9kqCYhIgad7s41T39IXotwVATBRowL2yBT8k/0
kaS3QHBmVwi5Y9btVLVjfIzQvk2VY1SCdYMQCuh6pls8Aeq11K1cShsqlZsL3FY7
t9vKpyzx4Ra/AGqlnGU8k/2HpLrr42rmv1ZV4I7NrEuVV1Jb0LBsNWS6aEVnchC8
1RUquVvpvyDnhThHvdU69a2CC3/uYbJZJ9v1YZee23TQ4OqAdlZiq5p//9/cS80u
da31WMAmAenzDwkTZY2jbJwBvhlSRh9Kc79u/hEiI166bgsKxEKGgLt8HjLQywV8
s5efmcx66QubLTITHvqGQ9b5Fk+77uKpzq6eufGQLEEJ3CFtdXAjJZz4D1q04U4O
bVAJ65nk4VVd3WPCcNRrD9ULOqFmtsC3WZNimwOsMQssIGbH9mrokEt5T5MBa36i
suIurU9WNQ5MHJsGZmqd96I4ZuO777by318Leqc1s7zVomj5QeZmX1mVH3rUx20c
IiURGJX/+GlgDTnnmoeItOpcFyxJUkOmFKjCn+XmZnZ/9liHNCG8v2LAGcAScGHd
SPzsbWesCIflImNZ8uiU9ZXN1E1d9fXkH40MGmhB4Sm86u7vgRaSBxbRhHWLGDK7
Wzs5Ev2W2S3LQOsvShkR9x1G39C7ydUYN6RWryCwHBdDGSwoKZg5cieyDtz9MM06
ZHbwWMSL56yrwlhB+cVyVfcBEa8TApp/2+fcli+8RFDWP9jhc2dX2QGilZgBmwJy
LSDMBSCZYD7mgV+24Usc77jAPs5WPyJUGVZ5+MjrhiuZiEMo/kFk/oXaGFzab0Q5
Txiku2a6B1NJaTTzOcYKaYfas6WEaYLs8sreTdb3c82LLN2pLZKWrtLru5oFN3SP
mVyMVbpzdtIu4NdrgeG/EK7r71n1tqMoOqHpjBhV93rNKD8ugLSo5FEG9a1j19HW
UZX2q6lKldxRjUZ95yDEMhMJcuVYLt+QkAWlVyAhHZj4vzFPwC/N/U1BuQH+3wcx
LLmOk2DGOLux3S/Ng3lgTtsuc6xyFoHKMLD6JiMehMfnzNr/QPmt7Pf6kKczc2NJ
ULRXJjP3oqgUlelY8rFUuWFojEdyMbSNxnk8OGwC4Q2OuApeltrH4D9QEw9RBgHy
9TW1sDXU1ICaiedWRlEiN7fcNfZPgGEaZ1OkvAJvOFGZuEOLaVuGd35yJOA6m4ND
r/IIgjleL+BO3zMzL4hpTblb/ErUWn+4elVBjtzULUeMnowbJzyGufaXcyOCRBzJ
c8mOpIhDAsnJ5lPRT7UsYt8sB+93YpO2cZxJrCzgaEpskyX0Nl/Dy3lxV0xqo6U4
gSEtrJfN4PluiiB0dMC+4/69SuiFL5X68UUM/FY1ueH91oTtXuYXwt1AALIRfl7C
1FE5dpDnODmvH2OsvzfkDUccDCEpz+c5b64yRdwwf2cz6MXFUcyephIQwpO+pQxw
CUpMnpkeOAmqpHgxKvhmCvfCrsaXVmdA+GTk+p2+S+LuVIjNPNmNMDU1uP7U2aSx
px+G3CDzeAVFN/kljmmvWS30O2Y998geQsZBy9KUU9MDs5zz1c6I3Ot9XJNHXWv0
+J6ZA58tGHe+D4eXo9vRMDm0bKdY1brWtaKB2HFXvT1v9H94iU9t1JESbqA2XXch
8jJakptrAlxGnBXnKfUX5I7IeC2W1XlgeMPzf6oiJM6WX8ftW1S8+q2RqcHuYmhQ
KUOeB/oOoUv7b7ntOB3ofcistU4a7mqNvcMK8Zx+sYpqYisWQAwebfXHmOmMyaDF
aXZ8ziZO73ALn1Y0I5i5FU0xWBTxrcuaI3yzNQ5MrbHer+DdaF5WzdlmpmixayME
q6pKu42Pz5pXF6ZKvUe494ihAPZV/ZnXhcoC5ee6yQnRHh/ateR3oRbph0IQxoec
8Sh3cvwyAoppoFwNCyXDqflnFd5uURnT+ZmUhepPOTJsoQLXK93RBiN5RVj5qCsX
ikgdj2QVej+ANyhwQtJsicBcPwEGZRCsAgEJLhIAQ8f2epbKkXeCKrk4eWtOxmhK
YwycNdL0czfK2xKp0REOR5NyqvHgz+QfHNTRnh9kn3u9z/3FWU9dIozuzjzTRG3/
ibJ0FXtGalDJ9LknAQ1aDIarDNvMsmFzaW3SkkKy7m1ZdelLQhk4uphqXMpt4bvD
ktroFtfAhtOswOt2aCdGdrDuAAwtPYlxFwKRbZOPAoYgcQ1N+Zqzgzy1gIMtn14o
vz9Hadcl2IIxsSr8iBhyzJjGTxUnm5cqzsEf1ri7alAja6EOTussCOMzqGFrc/J5
HIK/dkzoBfKUU0ZDrRcfg9kqd8n5/8s4kPByhR/6v+sTyuzdsbX7095/WsmN8wk0
mbr/LPrFwq6vALb1e/O6XcHrm+fXLNgPqiDE3ZIazB1s9ocm3cnqyDf4vt/DCG+X
3ShoQ+bCAuKqfmrfcL5Flp2SrchHM3r5eJRYshm/hm4b5GehV1Q9cC0Iq9EXucC3
uHqaoardOBxI+5fSGNIaWn5nDeuftfKu4CuZ/kU7rksGoilApiOMSzR8UxCicYCr
zsMFb62V6bxMydpuU2fu+SOP/PstpPuOIXZA02jErhiBtFt8gLuLevHhQb7dsPI5
9NPPwDKLJfyhvwOoJ/WB1KfZ4vGjqis3VP9zR5jxW3EN+gWbGsjdM/kCNE/OCkAJ
dTgHy5vQkkrxLuAIq7DsikyANHOCsDIbeP3yFzmvnxL88m4Pp6jORA9B+/DnqC7R
fSy/c6jHdi1kAFF9rxLnvMxrF8Fr5ej4oDMofpOv6E8pDkWwYkENkVP+NCE6LqLP
Nh1bN5JTqfTZXT1Ckfn273K2EGZoZgOk5R7O0Oos77f42xKzi3rmgxTg9wJDQ5Ym
/FN/8zu5oBTn591GqW0zc7R5sOs/x3lWr9AIQJevmwJaESyrapKp61H0nRQHHrJV
HF11JtxM8nzKkn+6BR9P5E2t2QWM8UPyY6USiTAoAgBxVWRQq5jwhR5oE2PRAWAQ
Hs/zNeQran6lq1rh/sevdz64dPW0yFZvIAlbT6j6bojJGBxyd/978oVwPkX+0RUI
+GpynLZWWPdLbZzZ+YqY6OAtIHAM4RAfNtt8WvL/MJxrC4kITHX2dV4zKf5IbpKl
oLtFnMIY+Mj25jQYHib5QQjyKJuThLSxh/QtBETXrwyNoa3pP7/J+YVY5kQWMDkd
lrlFwCzqXYt7lzoR9MyqNLKlIaG02vhxplzGdAW0c583smrDcgNz5uVNPtTw+0rv
bFgtjz60oLV9xALdZem0jmC10zsKZq7n7FFSbU0JjfmgpQeDnJT5VGrXcbkgS4xT
B5gowmprvniR2L8EEWXKu4s1TQsC/v8qWlM1QXDLen4HQ58H7Tui3jJ5KEyZiMlB
4kxZ07Gv519t0C4jKxIw4arxseshhvoUMI3ugv07Su8Ot64t0TM90pMXWof576Fh
IPARPebAT1ZJswm2nHIa0dx+Xov6jhDjjcP5VBHHdUwQvcOp4icmhVaMEmGIcNko
c4TlZa7FGdLEh9p+ixJBWit8qNYu48OQzCjEfOdriQMLPDxw9u0tpCW9QEZ01wk8
JpeQQrYtE1iw2BNNNRNnP5Q9w4/hg/DAK+0wMmGfoPeSPup1mT3Yhp5Eg+/8v8hL
c8WdttJ+Rv+7J4fD1LLyAgHAs/kNPGo1TTCmTx1chXgUh6ZI/t41Qz7PWz/L+ZpT
wpuj1CNP6D/tsGk3a5usg6e18QUE2RHe0dkPVtvVT9CJxsq1pIpf/QRIPWYMNzQQ
Ad7MSValvJzbG7uz6DC5eH6bNut0SuUd/mZsNbRF47WG2qGLwQTVjGUAYn0HSg0l
E8qC7wvXxXkO0Zev0sZtDlKLfPyyZEnWEagd8nxNsHiiPpspvcBv+z6XtQ1du78H
SzYuMTSEyqxkyN73ymcd/HqWYcsRxrdyWh4xauwubJixp2jPOFl0Q0JYR9ZI4IOe
F29+B0KWdNzQ/rQ3TqcV2CQneahaeYLtkeA8KBj9XZW5zCt0FUkTSmDV5MenUubn
J78R+uA+kwmcOUpMcD9k8YVBrO4t284zLp1GMxlSsGWK8U7iid9ZeAsxeJRB/rOk
NBcAOkcrYd33BE3JWFGOTYgBA9NxAFi2KL6lLLzOZguvAAQmzoL7av+iYa9Tobeg
nApmy7+ENbWOkHOPeq5nr+swdSjxRqYeaBKbxvgxkxnzGuPAS20UiKSIlniEhthi
pry13/5pqWSsKSyXTyZB6NWJUlu1s1Z2cwmBanij9zRzaq2h3ToZHA+zsaRl+0mV
1NWNS/ffqwH9+AQTMGFdwQ3TA+OcKPizjchRJ22DkTBOErx7Xg2c9K+deXJqfy4c
6nFLjAQkrcgawqUTttKbNtQ04NstaR4YdBAiajAM4e6S9ZDj0l2G5AwBo8s7rC//
c5mU6OqyeqCWg8PznerUh+GhdKdqZuFKZVQ4LSLW0MVfm2c2LbePeNLYQrVM6n2K
0IgxqDEt9d4UYTAR+ly+jkVe1iIk8Iu4ixy+q+kh/7rOceJOl3JXibtqweVBeyEL
me1yz3mC6sasIFTCIekQA4wMFRTG8M+POnarDwtB0+0lfymhpKDTwac34ccPTt9W
XVojHA+Rhm3JGyN3C7b25DkxZwL7aGbaU5AGDI64H/SkIl/apdsYSUK0B9FlBsAe
h5+Bnm2oIF0OB8cvJvdurKbFS8o0UFKdBYGViOOGw0lc4HPyp47PBFKSHxOb8Y8D
Rryadvq6LxBypmLVEMIsYISTtEWrxfWxIv72pPwZYGMUaE9cfsdg7338vIBz9Oiw
ojKT9ebxWcnCvnFDAfsqXaJe307/4IxJKtMHmn6U5dwCAKhfyCCN7GkcD5VirJKY
Hfsk0iSyez+/b/e8MRcIYpeY4CKwnFQIy5YXrM+EgdU3YytkTKoq2aKGglmUaAWE
HIbOrAaNJWUshJ238JysUG1afnSrBpNINexuH61PRuUuATMh87j8twB9gpzMw517
aRLFrzjSQKrnGlk4PiOub2Qban3R8N891s+1YA6ZbSxe68fv1ZIp6UCMOXHU9TFb
Nka6YxW9nQgi08rbVNOgUsh1GgOByFlPhuUP8XInsdQG4kBVgmq4KedsyBByYmGK
ZgM6A+p7xT4O3f6tNGuVTO/VFLHDbBwl2zimV4QV3cEpfw8ZD2hloOE1E3j2X6xV
P32DJSDJf2KV/i9hLtIEzCDh4THIMBx9Wd7v5DJhEhJlGDovdvE+iMcIpAWylmKg
lofl63xdJBlIkl07pi9c1RjKGpRdCrY86RVmvhxb8hx7h28XRwEgPzBYcJFZGoav
h6KfTbgkaAeT4jjeIBWKgtHFI2N7a2cGz/16hOydrL9UiiRqEl0g5I6AoznDCzZw
nQoBQPbZWiLVDSQGFGsgS0KMgEe2ZRkNbO0NAcLHXxix8htpTaNLmcvDJevnZ/jB
7VxfDEy2QkV14qIuWxIMtAGzD4TOyg29mJfmMIQ6D2v0ywHYkI5Fip5KY1fmqyIf
6Xol2O9R9Qu3S7GCbYGW7c5Ybfksuyq/6wTWVR27MmDzI+IQk3MzQUjki+uPrEdT
9gLLE4cGOR3vWF+btAoHowD/2/Lf/2ZHIp+GqfKZwPGEvmvgWJ8dWHxoMvz1Q6qO
AZ3h1JezPVGmqYUiWISOjVA8O0XoWMQbh9ijuqBx2gRwO0vy5Gt9790tvyUdg2r0
M9H4RDx/9fHtn2HUqezhIa3jpzK+LVwU4SDtXwcOUa2eUKahtvQp/DAOR8ovEbId
TukIGHWeTcWVmryn2AN8nZF14b4+JCdr7pA4mHuHzwMcgjbTqb0EgtNYGf93aoWM
oB0RvSh43NSN7T24a2rZAJ99vha9E7QwITwDigqk8YEyB/Oidxd17CPY+qNF1c0g
AQZ0HypT4eL+e1c9WJm/GjNZtWBYMwzyt32Fzgsh+8IFmzRqPozsYQxZ3FQsthfB
y/jg+ucC3qx1ir5R2CN93HXTA6h/dxSWz2dN+noM5CPm7Cr8MXkSSH15/AQHLaT3
NDbpwSXd7txYLo6xhf+8RP10aYtRFBia7p5OM4F5AQX2dIsz48ZNwVi4LwyeZuvk
HMlJ6aea/GxQ+vJGLj282VUmrxNMeMnbjPyoFnPoxtdKYEp7HhAM2JrxcElRzT2g
i6gK2HSr8sPQ2OzknKEGj8ZM6DbYWIBIvIY1XZieLfNafPlF9SW1TQbDJc9FmcnR
+I88+gEkIiSArvWJPO/5HuwR8HHf8Fcx23l/7TFOvzKSr0lkBaM+qe3PP2YoECzB
XabZzNAXXqpMozYBlaC/PSOnH5U8Vdg6jBQGISPmI9WHkPQZO4MVQLvRKvrpyVx/
pk7cbJ66pCmG4ALj8Ikd9IoP4yzRtwAvFtkQIUSpViVOroqqN9HTOFp2OWEmr6sP
p5Tjk5ZfxWCkgf41KlpYJQPt3OMALKfYIypuwvNB8QZCrG80POHSz6ApfdnVA+Zw
67GEJ7DidE+GjkfdI0ADZRtOr4MrTSlGmqeRmcwCPaO/14o423Q70+wk5o6RwePJ
JVoZ9W/Rf5ldjc1ERzOLKjoAyCp9cCQrfPcX5urph8fckQbZpUGzlPT4Y5IRnF9E
ceVX98j4nGSaNZza6aDbBFftyD/D1lLaIpNJyCQuDyYzUynCKXkqmx5pZu3qBvDa
CClUohHFbbF/oN5kVM8my9StxV8IYFnEGKiy4pHYaG/xXp2BPoYkWsaGOSwCdKIT
eZ8UhLaXpE0W9cgiSNClKz7i9fnL0hlYY3wsJ+Y7k6kAg/ZHFoTkP3irjPBvv1T0
2QMscp0uhve1V3R6b2+5sHfYGMx9xLzNdzfV7TuzsHEpEACcCaj9qQ7d6fRw2gSr
57nICJxh4KdI40mG2uy8q7r/VF5QJLReh80Tfvz3BIDQXhEMeoUOmBfaUsQXG5M2
FDEx3n+1adaah1yBnu8iVHPvB0hpfEsLIavoiIKcmel2pWTXBk6C+2qfQ2HusFZw
9RKgRewrkwdWxtgvq+plm0Vq64dyUduT/9qQqDy9LkzXc5cj4RIVroBEG3QT0DeJ
sZ81ah4P/KKOTkfqexchms0D6hGfEwn/BYLbtHR2nYWQB+Gx6vcxJsQ8E7hGkGPJ
1wT2ecF5YVayWfD1qxjIjswyC/Bi0a6Bls/JIm4cjgjDzojuv1msnekeecKzceIp
/HZHu/72J6dQVDj7h2Tzkl7htEv1LXLF+QlEUjt7qAJjKKdjRP59JVCdwawD1TlB
sbF4bi22QlkEk3PvcKS+yQTPBsOmoNcmbSIR//sfrB+XbdHTJ0jWYxKMreLFkhB4
SKLaZlqVf5o/t5pS9HbZRHUwUZY4N7vUyj853Um6WnK2pPYJH2zG2vJWoY1Fol2i
lCog1CKrsmpTJv0ki+iEQqhl/2tHFlh6vTuDmpkOtFO9MdCB/ZlBgzCSZxUOFg5S
h4qiUq1G26IRdnTscd5bhLETlnAx4p3wWzVIBk6IQorcODlvTPR4lHP+AC8QBW3n
iKdTA7UeaJa54FIVerGzGD1Zt6qfBHnxk7Oz1nbbtSn91aUKe1Bf+nH65v5ThGQn
HFDL8zS07aLNXaSgap2EsvS5QWy1SKC8MQVuSu5XX37wk0U+MjCuUJqiTdW7UVzM
J/yfOYcTPFYKP2YnV/vLbc23OhlpimzO39aiO7+abl/Zdw62PNFVpU6CV+jUzLYj
Z1dDsD4qEQCi/5+qRA/g7M28RrwEl0UIm2LTg2A5mmUxxH5MtTvYJJo8ZHekNf3b
GeNinmho+X0KRj51RPfU+IO6qG0UT1i1NisQ9lsUdU5bYpuwdtshub+I0P2CD/ak
zhJupsyzbLTAczCCx4JCDdNgG0RNpN1fpXU7EdC5EzBjNgO0hbWpXMLXeYgXdbjU
doghADiI+xII7YKOrEpYFZeQWpIuCoDJSnpkCckz58MUOwnio+rHf4ZQtnae5Jym
K7R07MqlFzftJn6IakbSVELTbDenbMkWaNC9CBvlRj1ZccavepYvbntn/oXdUGDK
xVg2ky2NSg0z+tFdG1lNZKBoe+N26IXAoaAV3LD+nx6x1TORAelI2QuFEV1IA6LT
AuiEhVi+BC6X5HkUefUwykPtahFszXO/g7APxjAVE2DZst1AyFXG0U4qB41OyKF1
aakI3QudUpC4G13E7c547/nTyycsWhGZkJt4tdO+seEouG+L3Mu08zpos8flLJTG
ZGX1+qkv3fRKNO7+NFgsaP7gtfCR/7ZUjwRoV0GLuk4Je+cv6Irk3kkGzyjMw792
fxE5LgpneVjdW7JX2VuIC+EhQeN9yoV12yCnSu2gjtaswtSbzskK/Xp2iSkCETb7
dSCkmSwWS8sGHc1LEWGkRpY2toVLDGDaoka8u0OgvJhWUSsU3ykq17VtR9/Q3VWe
tZqqXEueXHO1d7+i34n6FpPe5OWmWf5ruo9AHQxOfHraKjM4FrnPs8KrqJCa8ThG
AuNCLCCpXzNq+9JuRL6cVcDj378UNDMpH85TAIG6dnm41ueekjk5KyebtCUwIu4c
eB7+OKzYp//2XITrz79a9sDNMNE1iOMCyJsE3uMgDlv8r+I9gWpw3w5MnyKsH+xM
IVnA82V6FopY9w1bs9yNwJ0+LF+vzH5lA8qGS752f8mj/eTeg582LYog8fSWyYqN
RaV+DjzUAUbSq9HIM6gmnoi+9XlF7jhl5I/YXG6tMT10dEOOXQQ2AAyDfj8JmBGB
4KKIyxh0lfjjRcCJ8rORJr92lXgUpEe54wDP8q8dX+CJu4Vtkh+QTK0/tRyvl6yr
ji9FxpikK9uVMAa9GsD3/niY8mOtOcSlHzPKkkwORYziAuCnubh61V1plFZ/X2N/
0laYYsg2oPwVceQkdE9YZACaC6on6WZmbZM4C8gZi2cZXeNL92VyLtMsY18qPyr9
7xVq6L5qYzPLam4362plmZ2u6sfltqTcFGHk5DItiD/AmoRNyFBu+s2U8LW3DLQw
026ndn9tFd1v2T3XJU/bFy2VqG535B8wguBROXhFDPDF3KPQ4/MX9rhdHK9F1OYi
0nqXbzh+Vne5rsqbtR26FwGFd/WMVWrmOZoHR7IpHuiAEhS44rrjVWbEw0C9rZnq
0utgnnUyey7oHR03hR7GsEFVmtmGSKgkvwasUF25RIZyIqCUCTyCZuDZh+1sdk0C
tmFgaQeSTJI8f8zNJxFR3kyWBczyYTTh7xgVKhF67tkb+jHOv03lTi5fUa5SddQQ
cSOH5YzWtWHyBt2kh+Z9l1st493u42rKqjxwAE78Sz5Ebrpir1W4Tt7/BJPoEPmi
fybM/JDCQZCpL298wSdw5kzCPKaE7HA55lmha65IMdK44Od0vML2W0Rxztv8elyS
7CaCWoxxij2auy6gf0CIgwe+6gWFYQfQqFl1JobzlUbZt7DSGGPgqaiW21nsp0jj
tpjBs287sVvu5k1OzLvrAVavjvjVztJNMRFYfzhYdPNpKsgatS5Ymx01yZfcPD/F
3qp5CT6z7bE4X43l7AhdO+hKp27FhVHFmZF5Pi9QuT9ideHSNgbIIrkNw6hbqrjE
Q0dFGp9EUIxaAyNljkR0b9l4iC8QeAFIgv942C2J7pq89DdAiAv3cn57AXvfFORD
lWyJ8p5cn6GA2eCj9drGLGDyQ5FFeRhFsUHfbosTCF3Pnq4gkGif5M6ax0dWeoEs
hvJcB2f8Sj00i3SUACoQhM7ffTNsDgbx6x5ETEyymK4WERPPgOmrDsy5rDnfSpoi
6JWOOmZ5VQAkh0R+tzQzjg6iplbXsyIROx582zuH1B9dDEYzTaMhNsFB2NkW2doS
VP2nzKwYP3MhaYC7kPpRa5aPpRNVWkHWxpAkzarabKJujt4d7NOD3U9BkfHjjho6
49DbKCeG6zOCD2xDYmqMuKSxPTxBVIo6lsKslDR57NaGbHc+6APcVFeueMDXXbj1
MToeqPGJd5szQFW/K/Qe5gpbi6w2kHPuahGItCvrsUVCxcR76A5KfLqt8naSOgMz
QbdGEatAVL10Po62Dv1U4Q5HdANaBUYe6AgMsIhRnxbxIwWi53E4ctR0a+zBvzal
5ATLqSnmusba1vlzyTFfLjaXvbfsC8zsRy8fFryuC1T+3DBWxX6AcT+t86Dd3enA
bgrOLuczwXZ/PG8zl51Siu8apEsNA/DcI1tnFnXSBrglgNy/Cggvl4eA703SfOCL
mGewwq/KDz9f47hWt1aL2lHjNvOBTnAbSKYoy5hKITIcLemiEQy9hR8ezpuHFAla
Qxe9e76pEUctGpM6chXqrwA7TCBNiohWamoVZonDrlPxZud6SUnW+T5ShhUshQcJ
6BZ2aErjNQPoO4sHUv5sz8NT/B++65jftAX/iisE37sRPC0LADXjXfaAz638dWbJ
E+TxHB+Dh7/dg+AWvdZ4fJcuOa3wGWuqocd1G2ehYV6JfmS4EkQPXEsrPbsinL2F
UNveqNy5q3HnbrHA4d4wCPEbhQRHehAh4Wz2rITvfOkASapu9SMWnHB7qRkhxdDt
yUtpxF61H1lGzAPaHAqZ1QCObupaZkcWKidTiazLEpCRNwD+tYuRk6jKoiVVv4It
XuHTKuUN82uykR2Nc6JRvgN88XTHarjBQvsY4Ywble0imGszgSZcVYC1aSSDAb4Y
QwR3N3emeM+AMFTe2MqFL82uxP/Tnk0tB4VLuOReDFUjYceHeUUr3M4VhNwHU/BK
PZfBuwMubQduN7098Sv8aCxN229O0IJuX/uJLM/i8Qb7h1uC9l0aN/zZb9g5rETN
QYCCERHtT4vdlRrduelvZcO3GIJ6rRjA2bhA1svIQ6HY5YrmXmWb8VbLSGYKRSqa
ozmpXWw0O+N3NkfsSbmFzLTqqna8kOUkVmdEHG6uIkBJzwFebajepumCCQ1Bybhr
+PPKsH/b7opXpwqgeVKyqyydrNZgw0fMmVTIOHWNG8nbxfWTYC81RCbF6LkADmrs
MNlB4UfBCMl+czC0RZ1FKk/+yvT2R+NkVqeB3iRHU7LYaxVcC8YnkFlXfnCVWs1T
Hg12ntaVWNx/E+tPteXa21aORSbEb7T8KroKErCLUy+4pN5SwQgSrjXYkMkGhjE0
mercV/pAczhN61ZxyRrAUoCvLsDGDojFFNK/4cvYdYWhy325kRP82AFFTfyU6slB
xGlbILpkOKxSrKZ+qEnc/DSIf4CGtaotjljKJ9o3mdESUoCz6MLYMVFvJAR6PG5m
8lvu10EKdK63d/h6s942Y+H/rmLgKcxTjUypMpMtqnQ=
`pragma protect end_protected
