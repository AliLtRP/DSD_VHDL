// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n0kVLtoFtFYmdkLd9hnBmFtI+5TIf0S0vxUSd+2eVOHUqNELRCX+hlKLMHh4wQtY
yQOJWHbQgNPGgrxbgv+u3Om9Qo4EDUoJT3VnwrbyA8FyL3+IrSNXyRbkWNw5eBOn
YeqGvVEZNus7srbzwSa06/NU3ml9v8dYGlr81JL9YXw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
4lOXL+jKrZIctTeoExxg5pAsCTH1bYYS0RksC92ONBzU3kEE5pooUojWB1emRAvv
N7aZl9Hj8bYFzRthnwdcxSDraJk2SWiYRswGGu5mzY7CojAdSH5CRwokKOxtLQ0+
sB98/eivow0GI0egZPTWyhfElOvCUfZeNmkUg6O2FpOp7jd3cceP6Drfy3jS1SIY
RpPrcTckkpnA0Nq1fT1dDxLGIdKn3Ghx3IVF2K5Rns1JYDB8hENTJy7kZEcIQ2ur
YKjKdBrUU45Gp1hmNDgDduUq0NCtNodQ8dt1DDi3agEJ1FF/2Z1CEvcnTTMZ04no
SXLpaJvsvl5/YaGdu8fJ8Ve4+iqgTi7pdtR57l9LXkyiyA905cZwAAkmLRRQX0wn
/sAT5v+VHjS55p4w8yoauWmSaGpd4S9bNqmJxWexNxlfQrrJ/te/7fx2WlnUr87g
5uZJZH8D3IMKJJSZYf54JkKfh18B6fcisRywrIH0WG9g0creWZR5PnDLr3x4qI/G
0un3T047Gl7nckNHkgSFhENHwl2ghaxSo7g1kphkTjST7KAaFoZeKb5g1UsB54q+
Dj8arwxubmAuxTeWz1pvneGmM1TqCkoos9D1QjE0tx60AgQ1bpVoV4vayr9uqhMx
AFhL+h0SElydhrlKuPW2kL9mlyIYg7ta1VK3rbUlFrIl1zFMhCG3gI2DKTqowPEu
eGtndokDcscRie+dVfnFmdKYZNOD9UZvK3G2uWo6/VhYMkE0COmVls13s3RIV6a9
zhxQHhnNqyQ+wB2Lo6YS+F8qi07ONRD7W3IbppgywpT2DF0B0nyyq0JgddepWfZH
uIgnN/zK6i5IOlspDgqt3UxJiBjAS+qa0Zdl808bXwXXWlfFW2I0v2OueiQdkfwb
yqK+NE7XPBU2hOPVEXi4Ewk00/nZxuTyv1DuwcFw1Wr9GCucA7fHBbxdXJITyPdG
1V2SLOUjsRJm5gu/YgaqKGDZq+LpnRy6YQhlzL+xEOZut9mMQGrSz5XMR2h55g5e
//geyEBQn4k5JUKRwfBccDGo38UmyHlGiN58iVMDr8gRpK1nsgMqKvkEuaKh6Hha
bm5XCJ6RCLKy/Ek5uXfm4BQT9j+BImvKyBT9WciV4bup70z6X6xtKiBCxgXLEv5g
9d1XclWBB3siCKnnktq3rqOaaqOvjjivDTNu+WhVCuG7MMnF+nHMO1BAeGMdNpgK
O9nppDsv41jlqg5A1BwN61SpUm29v7MOWRpVcvhE0ZaQlgnpoPJsBg4AyV1Ix6Xf
ZyVdU81FJTOlfo1kdGdeo6nUYB85g/YtKJU5tvN610kequZ+v/2tbd2fTWOW+x5p
x9gXTv4iDftVwqXw3vl5Ua87yeXS8wp+yKVKlAsbIX53iecjaWWyWHIw76PJehcq
6vNSpZx5MFNhyHfYQhUxdwQLBYY2/3bqcC1+Coy0H7qzGSsXNEWdIVP2qyxPIB1w
FMMzCmdDkSdIg30d21tzVcJge3OIU3eFKPsKK/cVJO6lJxLstf5xjawP+mL1z3cr
uMH0ae7eU4BhrQUF3JSrv+NRsBkAkywwmLrzLWJmYgIm+2tG0ROC+7xmSUuJcCPd
Is5cqQFgkEaWbyviqTGlXqJgTGCZfQj5BHHY2mt5MoZIfWBMp0IXJVx7qpCj3zFT
7stupWUZvOHeAockxfzlc29VM7mLs4E4512xUc14pE3tmgTSlsaKJk3+AQWG8Qo5
qpzAbjEv1mXNnUXHlG+Zc2zpR1VNXEwKyTg3fR5yGdUI85JDYhvkaqJvWrklBLqj
dkqKbizVJnkf+VOaymO+GaHcwl/baBonVaMEAZxxfV/IMb+u/YpVFRlOAOwPXk+Q
ovQqGlmjwDkmblt415+x07+bzEyfwJdnC2fR+6WX01RqHFNEPa7t+FOpX/uIN1lR
6rTPcM3hdsmup4slBh6nTR6JN8AaNkdbHs8IBGGpfSja0E5qIuuU4SPJyuD9ts+X
Voeis9zpIXqqfKchqNM4Wn+5BMV7miIObtrf+/dcdKt4CX5uSVUkh4AX0ubrc/Ci
cE9xL83aFC6Smllosz6OaVpr6kGEInscDcH8DGklYBNyEppTOWWzBjw+Q5FPXA9S
GN4ix2nLD9WjuxgcEPVTsaWmsP9b2RiEIMtAGiEx2LoXxYgCODR5+Sa+ayjVSyBa
jHcv6ipMExHSoLp4TuYb+rIJZ4d6Ku1aSCpRcHbcLIrR9hsBONJiRwJP8DK0z+6+
k+bGPZGbDP9Rked1VU1Qva1hIv1/4wgNb6iyWTQ6FesglungAWc8e9nWhVo6jbLm
zry5HOC0trp7s/hy5Ft9omswypVjdvwGtHVYrGY3pth7Yz0DjKeqHBSG/hF3ksRh
vbLAtvVKim3BDWcb4guMPywjf5tfJSyCNnHJLbK8oPweJhwUYBJqB6mZK3va6IFr
6P8LGpNfrgRbYyP/p0K0dY5MV5fO6dqrPRrQKcxGNmvkLu2uQXJ0mvIcq7HD3uEL
ZPBmSe1DkMj63LBJa4ZRHc/ZvRXlH+zuH+mr5Iz06FLHnZ+kSkinTkUIo3G3JuL+
URzKBuaqOJ8PRrqP8MjL/7RiooLL+RmQ8vEcqrzNPdrCNv6YJkOdFmDvQ9KmlxV+
wTWBskQBECFPDjnpVfAXDKcBa+M6Q3aUNEDy0KUQKILKtCIuX3KXmwPQ2jbSDuJ+
2L7G/6+pQVYzJSZYJZwHEi041yax/i4VS+0R9HwwXcbR3SX6XO8FB9KZkIRItaL8
AKkeV3QHbB6SuEd56cb2B/UNQuZ3EO6HK4UDaK2RDR35UHCmxBVH8JnRyLgNaomd
jTgN5MpHf6gBTA0ZgdO5O7GjWjTIEbECKTgORBV3UjeT2EPs+mNxD0gJcyzLX+yN
XNUFTqT4dAnpyvqGbzAuty/y8K4gYc+L8WA79UavYLd5TMVYwJP45MzmwpJmT6H8
qLsMbGL1SU6sGQOeKKYQ2Jaga7IXG9bo+RXncBKd047N9j0twCIsw8I1A88ov9sS
erxoeP5s2E5PiUlND1vvqHqV3nmex+Vva4x6lF3ck5Mla1LYRvmurEXE+mJnmnMu
Wp74//W1IFVV8P95lJXFDLLQehbIUqkEjjPDhJbXo4uDoKXNlS5kGuDMdItS9mWF
c06HZX9tcqFPD7vXWxxq4sBs0cc+BhKbj7GXqg1jO5zTbMDGFwv27gzpH38BiFAE
sZtPGqOfbG1ZAQ0U5Pxzpisc3ktQZrevSTIiLAccDvlwLpw0J14iRnWIvvtb1OP5
HnZ445OquLoCbyE49pSPMZjX7LszU6PLc6yz/ZK39fpHu3t+QuvSR95d/UQzjfhv
GXW5h3WVBGnKrlQfBOqzfGsRuT6SltfAeaqOxsqMfSwkmwAgULMG8KNCcjL+sfC6
PEATP0ZylfTQ70YvHSZgKsIfO0xPq9gjQXdMHXjBrdGS3LLR3gIUb1NMumqr6srZ
2IhRzwYNSxU3fttvuDNP4TV7JB2+L+vk9O1om9Frx6IWAMuCA1vtMKOruNXDhx4G
kr5xStMiUhp0Z6vKqelvOSuXJWG+TAbTsudqk9RYyLmyvh8kkhNgFWksrDaXwhT1
CDCqdset49iMCYN9HLXvTigZqLSVFxBvtvs4nHHnNNdy7skK6STWtR5baGeGhYDk
wPoYTsrnKfCS2Zso2qkaWyLOj0KB9uNTtfRFcDG1SQ9QEO3Q8eZQNARc5gNOspXT
ADhjvR70y/nJs3ndl2npbv7Ipy/Tn3airjF1vAeS7hoCVyOfoBg29sEhV4IB7Un0
1cp20O3I3tngWLS1A3kzq5fGTjmxhyRnz8JQJ2vRs4f1ysOCkrE9J3nDrbD/TA4Z
kxvZtGIaE9CIw+Z6KpIj+PAkFHasc2Mc8/RdEZEObhJK5mTAATeUfqhAZORqppvs
YjG6dVCfoVba6bx+M3+HeQsHF0PEJ4Dl4OtgR8Zd4Ank7zRxzFleq5H+O7pvgztv
WqTgdlHREysoNXq96F7uJ4cUfjVOprmAACNBuj3Bcxljzn7uoEq2zDKpVeH0PcBX
8OVuwzSYhY2iOoZCm97rdQlP2sSh74GwCVsCX45ksKE/NVKQfD/fzM2GRxXoGRyA
K+WBnRiRY7j/61QVK8sj5JVeQ+t7AKE52ebHPyIky4zShmxLiKPjWePDKxLRiZzX
W824JBFLi2+mEB1EPko0Taex55HVZjz9myUK0BqpxrwNZDR1uaoKBBIeanaYTclb
7eD8eXVNP6Jstf1T7nOquG8o0XGENv5R66Cufto7mFxKIN4NuOmlWIsTpDlxyVNO
lmfm+/EtTpMY1BjT8Bt6W13Sj8ABtvaFB1HJXOTOqLUsSPAIVRqYDmx/E0aYiQqW
jjW7PZ2AXaJLhZGKDPCNsmHov7Vl9cZs59EMRohFa9vnRrGyoS25GOvxblR7A2sK
uc2kuzVjkhwFCRO4BeGco5lWorDmaOY80vMB2eAzqK9swThFoWISnyPDnDOQr5tn
gGltnKN/x/JqvTIi1gkdL6HafKA3hZtDBAD4Mo7y972qBt0dp4cuWvFw3+dv62eC
2wWXnYi1G6yaFALVNfMkcCaKey2mr4fxVAa5NqFf3jdfpIi/h6l19FeOY+TMEBQj
DP3D36Cth75EPGFq7N2Y0akb3N3qcERAQM+vJcYX9oMpsjfZ7xH7BXE1mBmBbsPi
6Vw1joiM37LOUzXqmyia5oF0tKGlvSNYB/hURhDK0Qp4qukYlrK7kR+47baMG8A+
1CcwH3cT4oxk7K/OCa2TwirbA5xqv/IEr5ptQBxJLdJVB1CbgrxcH51CrhfYfsxS
Z7zVy5sR356r9tMV+/3fD0g8cMJVmNYLnK+k3xtJuYRGn+rYmJCajKPOqRygaUBl
HfavV9j8Bi3UQojGYCdQT9dV892bWOqEpV5wcJoQ6VVqOoWaa68EXpBU9sRYXKJ3
mP1MuzZE2gh+VidVrsHph1nZT68NbjrVUSPGk+Q4LUB25j3W9q7dpHhDgnXe96dj
fvSzZERYz+kGx+f/W7pfUySXhZqeToLDV/s43f5eJFovdfUdjnoWgxLzme0xEqww
tMb66dmYMZ024BWssOf3+pVhA/oJKYHSUTu2piiNKOyLdsf7+nDSCCA5WX7Kxof5
W+1uOwqv3MXUgi0IrcI+mVN8IlszPre6GANNacCPKaKq7IfozonZVjEWjEC5DOXI
f4q+ZwQxXlBpQqnToD4GiLby6WBNS4mqjnjRgLAye0FAWHTPB9cDr6ZSA5s2moaq
C66/fNymregbqLvrt24CQ99PgdDmF5T8VvUkECLs2RdEtqsWhFtXFYHX7Uzsfu6F
7hHmqRrbg33iK36InxRix2uqyFcUI0TNH4BI9XmP62DoNG4uKo9WEsNZxZUclIQw
QvTApUfLxPZWWvN66uPnnJ7o4VgEdtmHgB3YT4uGsnsy9HYpw2WqCgYSPnVC6jAm
U/VVNTFGoPlMTnA+22UKsTprCNsQ3j7LErxx0JVHxIl9msvoUWce15eMgiE1A3Ks
zAzjp5PdenQJwuJFRQJw6/ox2x9bLNeUIJmzjUKuPYjJzfTD+B4jWGi0HFSE+Vld
j9Untgo/Os8NQHsftLRSOhqa0RPCro7L0oEfOeruCDKkoZu32u7GdkRLNJflAuIF
Sv3jQewMy5LA6gelOoHbFY9EHwU0XZGsSubtP1T6KjWAZwi12KZNpRdQiu+vwDeA
7fRTeyUJve6HqxY/YmAXBUbFCk7XtaHPgGQKG7saxCF0QZ1oNCqKol9/6odqtoiD
RnCWSdboMxO/Lh/l8qKG3bHEvGmG9jUKnQLQeS4eE6AFxMKILvioiuFMdLdrhslY
7Sx7NLAE4P7mRP33ff9taPp0NXmz6a98b/ZDGsYB63betuyqhqTQsIfe2+oBV/Dp
sIeU3RTgd8ipkZzg1jEsgPefZA7Fpp88ILnpltMLWXtFpAV+IIHpdjkrKZ+0adcl
40i04QAWFBJlDNIpCHqN+GUfa4QHtnyxwqbc2rkCDef04RNkLTn6jz0vYOqsB2XJ
xgBozK+mphAJAj9ExcZeF5aewN/DDy0jNtVuRdtirIgGAMmmN0G/zvjD3jFVWniH
0LD0DEmfO8ACtdUTJWJjz/6AmPRHQZJ/T2iVCSbFxsUC97gPcohYos9Y28oVu9Le
gDE0gWhOB9Cy5FMke+uDVML5nMu7eFJXvEtsfrmOCenV0xMnb9mQBJ8AYjKOQWzq
vNkXOzksP9mK4w4gqUm3Q34yQkbVDWtQQ0skFMPh7gM4QsiTFbpdhqk/8bkMoIdF
kHWpEq6CQlrbu6UdtpbVTZta6lvGxdt2iJzXepnReNe6EF+3RGAsrDa6KainH6SE
l/n0MbZy4c7BApfoJM1iCAfX2LD4m0AP6z0NMvwp2wQ1cHgvsAzsW0WUYhIWDpOI
u79rHAdh79Y6pODp8E52SO2YguhCzmk2DmKbihMGChUCB8IkQj71AhRyeFzcVJ+v
Ogx+J2pbyj9wplFP33PiK6qmUl5+3Oein6bpvpI+x4LQhS50EhefiR7OHHkTWEkt
QnWvv3qYAx8VxhEVyke96sk8kDt+f9dvlTcmbBdmyBYfFFQT/sfsE9nfQmfUTgbp
iWwRr4xfpUwu8MQYnoDD0US5Ye4FeXAI5tge2PQNLbCCmPcK4DRdrBQvej8jS8wW
pnMcmCNwODaOYM5zMfgbFfH+C/PCGFe4eI9B+FomppiEFb0mNMWpkUAbXjb+eKc+
AuFt8dcSWPIkFZhTdY6wQdFRdVRwdJhpKo7BeXywpXSihWs88KrOUcmfBzEvmlzH
yE3+1mtxSUWco5brNJKuyJaqC5+D0Buznv6YnWle5EwjZ+7zyVXe3aMkbUrPq0OJ
4nODkO2fjxj9bS94s3qfyNqCZtOp+bRC45W7/EizAjnlBCDIYUh/XvzW2eiMxadl
gxi4STz5iYI6WkTmou8KedK50pwgnjzjPEipryFtotMrFmNfCCfWfEBlRltd0PzQ
x+jLfiZOapl3eRizOQbm5sxLUxjL8AUbo9/wTgytcy5MkNBOlaqU3OXBorRe5wQr
RfEF4BjKcv6npanvdjGl2KvH083c9XwiEAZ/pQgFlvqrbL7Mp2prupkfhu9VeWkx
x0TOYK6xnjYFBx/KP3v/G/+43UeGQnDKbxyWFF5RzlMvfPLmtqCCILfbz8xXquXQ
H4E6i4a+FNN/xvpbZT4YR5xCiPzWMmSvBdVIVFszvQ4L+lMiM1fMnugFgMH9Xz6G
jtC4xtDHPSoOeL/Gn5byHvHXb1HKitk60pOJ//toOqEUv3VvGSOlEDF3cVLp+lue
JQlJaJVqD7FX48jlMgLZCXW0LPuNs85wo7L/wLmu8U8GjoznzumhCfTDZgqWX+I7
U/i5knO+bD597GMIaJqhbPs1E+IazJZJpLm4pn3BwcPCZkHYYpSPf+mPoJfuloXw
l1if5ZveYZL9T9a+dzAJI0TUetoABYWcyWcoqos0TjU=
`pragma protect end_protected
