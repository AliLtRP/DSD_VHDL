// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DGPqnIEtjlWyYQO1/3LD+cpDBozi+EFQYDGT50Xmlyj3ZjJ5KXselrLHIqpsU3fb
vGL6RopcHLRLTTS4ibvlYxtIiB8QwtQOHFpaOtuTATH74V2kPVzADbSJSSLVhPIB
WVNzvilVwdO2sCR88gBzPu1bb7NiyVszBf4eOQLfsUw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
GgG7J8ZoK3LxQ8E9ArgUWAhIHoxHOsrsA0hN+xf8h9mV25/W9rjUKbErgzKl8i8F
0jrs/0T2orA0Th4i2aaaTVsj9JdFQbT85NzUKajB2UOto9gIO9EnyqdzGm2VEOH8
ZfHGi58p8z72GBQXLWIO41UnxTg5Wfm9rmM59EIiu6DSHxTGS6TDpRD/2S1v4bhe
PA8tvXP2GLQUXKDcIwQ2BY675Zzf6WrF2jkyt9+CNd0O6mhFmIb59w0FMqarC9+p
zqtln7EyB22jP8YxRFgbhk6EHXOtQ5ZASBYcDXlhZIl2SKy5GV8zt+LCRd/abR1h
d7zuOlZPh5PV3aQDkBkBe4YojFUytbm2jq9y9zH6A58gD6UWxukay9HvFops7q3L
ZajlcMwXk7u6o/lVaZU4zGzI+OKynVUoPqk6DvSknP6M0oaXacBuFWDiwvu/aeNM
BGYblYuFA6TXHeQHbJx29XfjPyrW8K1sShdTxtf1UB4KCHvreU6gex2nsfU+T11g
vZp5RnLyqg+/Jg1lJ1HUvVKkv1eCqxp55cAqJjNLGbCtpxLcDh+/JyFHfmUu3MXc
A4CCBtytnBeHRqBwhIyTsntwdns7bM7OKQERJsJCMZNY8iBbezW/SZGTDbEyZPU3
npCD++ZkGyo57Nk6vO+wgJdxo7C73VWx7VSNku0w0XoRalwSdThURMJXyxO9PbkH
D/CT2SJhHOKT4tHFKo4JgVdn36w+Xglmt0OLoLVz1PSSxs8DPJBsXfELqIx0ouKY
7uiXiJSEJrwixgz7GKDlhGgkm+QOyv2LBpNE69lSMQjp/ckxgiEh1Yosj2+eM4Jw
PUTu89cKuicyEaQ2XRSTt+mDJSz85PuCfF/B4BT0NrufJeai9y/veofkK4u4NvDv
GmGLZsT4cX38BPhq2Neq4XGeLXJRJa9lUqwn90dvuwDfeSSuPGouBs6lGBZTXfm0
phLUhxFpql6ethx/jNgX5ISWTTks5kqyyylofcSrCii4PEHVATO812STucDUfUwX
qd3TRQG3cbocBhoVcRksG0JNA/47SP/zyXI0Ro2GpTpiaFNBG/fLI+dZqqwvkKCA
5R+iEmXX/cvJ8zRZMQZfC5iD3SWE/1gBwTWWxHcmmlN0fIESm8bCkHFbeu5Zwk09
03R2OBzuehwczWNq5zGLo7St8G6EJNBxMY9IM7jX5+rnrYSLOOWwKFLYpfWxyD67
3UrVhHIy5uhMwXCvZE39Gk1fEDXZEntYhiOfXWLSS4W6vrSmSm1jP+vB5qBuc/sy
sCx5PjvFAz4Cvs4saDn3vrfN5piaLPlMdrvf4JZI5K+fqiseBsmDENRM8lg6mcL1
bY5y5cXzqCWI3UbFUesba8OoQCghA21EDEqhhPv1lKUqWWUMki1g4TVvY7i9eR+6
sKlk3RF3N9IYnq7sSqDCeGhBamUiBTPFpUis0GX16nkPlvEbS6E73VdDE3m0+G+g
Pkx5JlnktE4C+IUyCUca8TF4vlBtkbmaX4LoMBcj4DCBQy45rPG++bbTK1MQ7cEj
5ioosFg4XDUfSEdieY+BqZa7Xf+x0NRdrfL8kHj6rgBqSdZ89NlQQOFBI1UqOkba
nreJoaG+WzOl6mjOIYM0sPLgxJdXWmigC7HcJupym0fr7l2Flr1lP56FSzctE9kR
tZ/FVD5/FZD5Nf6scS2Tz9hn0xi8oH0KyvOrlFZgpQjJRHMArNGvX7NdqtBN/rkE
AJzUco2v2lwhLlDQVCC/ElL+OJXCfb0JV7HZhC6dNrd7BkED1yh/bjOU9jZPHZw9
5/Hf9yEn3HpvqTR7epjTKF/G+FF03wFB2mOa8j5+LaM6Qh0uaQ3d9H633wh8XrKK
wk174bY8dKJF5eSm0l0EIsXrL2LcloaA3SRb4DJgEE8+RyeGs17iXvMpDmWn7PF5
ejxizRMIq0zw0S9UAu1Th9L+GWp+TAA9IIPFkE62suht7ml+ZX1pj6eRMzKQbmJC
TjePabyW7LZlDMcHTNhEFLr07Qtce4fUI0SgHSa2dmxiQJDcsds/RNEB4akUofS2
y9bG8L48dfv9hQGlAwU72eQgZh5cBdhWvKX/3v0BgdcCgAXcUzHnwobxrnSrmQ3Y
wvE5p89be+88oT7WhUKie55VTuT0W+ExBh4XTo4qvCAIf6VfpSMzcOxKm0Xfv9d9
mVadBmJNqK4YlD4tDfb4qtnu4q+HAfRIZxGQ4IKgJXr9jcDCPCgFRR5rO7fl/2DU
6sh2Bx2wJQVLVZGIAyqXZIpGnVgmvAa/60rnbIQ46AXkqITdnD0o8S4PDMtEpvko
nnyc67L9hxZLvDOuKCSrE+9FG1koLH0irNC7JUVawY0VNYFFFFwBttlWYJ9GXdgf
V+EBrmvrqXRMUkRHcQFSzn7QhewXHU5w/NSMsZNGnmmK/hx8BrKVDCc8c0kcrGhY
Fm/nlMPeX0QwOaQ47f7rc5HD5SxOToR8xYF3U2F4Tu4xsrE7sx0B9XcdimeLA0RQ
jrdXmEMIP6hQBOG0xqABoSS73Ph2CP3/8vrGL8EnzQ04JaYcbaliR/PpHEwwAALO
GFVR0KmRjLhif25diSUEWw3CguatCiAT894NNIkRPxiERFtFOBU44Gi/NlOUmyCd
eIHuUjTCxyebF6/DwWc5KfJrOU5VnC56LJseA/5hdGnoZVTlYOdwmN6+9cFuoO3o
EMsKwBFqXKnvfiHPfdhiPjR9Esb0P1PcDYhHfPRtxq0s9inUQ+mTo5Omxn9sH/as
96OKOIyfuzFJvXp+DbRLVhwqrozfOEuyLHyEMyf4aJnZ382D2p1j61hF05lQbaiZ
AxTHLQSDTxhFKGwCLGoR062379hVHYrt3XwemC1DXuwQaq/IKT8qJ3Y1LNpoXBv3
JfoZO+sVzyMkOD95xF9Z0CF4NRWQRNOrhp+vtypaOQwXi4L1GUJUud5TqY5VceR5
aJPhNDrJ88TrAjwLecHPAZPYgSJZoC2YggKP2Q2YPXrYZ3rFyDJWgtgwGUyjoogQ
rY33lX+6gHBYp6Zfqo+Fy8CI5uh/e8jJkCpez244AUkBmGT2P0W01tk5iExgoMZ3
awHdlFXE3XSf4OwJitOLx22sagsFz+rF3YBFDU9r5KOM7HrRdZb+YEYlKXNRD8uQ
joZZO471dCCH/y62x4mMzNuo746q/SAL/b3kUYyHeNzuQLE8WNZm5UC0fUUSUCUQ
cZUfuR3SNwNkO1xpFu0RBcpsC6H9tM/Qo1Zb2H1bQr1nDxIJE8OmCaFN97LF6ous
OsqldP1bnTQFcqXnyBgWQSW0x4TaV8q3LHq4RSwj9n+gvlB5uRAivFspaDEsCz+N
qFLPFzUM7Sr+VAamUKnGLjEA1k1wm4Whn/kRWDz8+fJ1ivGPgOrrWj2ymKwydGGz
bra1l7i43nuxj2+ZfiSkpXBp8XwUryo0gdvmqZrW1UrH4A/9x4XQGyBQUtOsRiRn
cwoLiYITTgkE84mVxbZcHzwosi91QV4VpuO/sC4X3wFscAGSY/I9rVmn7bSb/TG2
OQGs2rnAA2uKCh202fd9R2cbOYGc5ApGSuw9bFzuePaLhn3TJwMC0WeOI3+CbUcs
15wVc3p7HASiTtUexgRXW0MK9arCLrPIrflcaffjlzaqbVG9KyYPnn4/EhWK3A/C
gmNwu+GUO2Zk1VytdKDroAsSSIjr5VyHIlnIUnNdWSxTVO0gx7ROmjo7STOXe+Jl
v1+fOoew3oopFUOCCLmdJcK+jysJVflxjbeswaoKKKcDvFH+tuI16+S/3hMp5mF5
DFZ/sQqCSuVOpEkWxSOTYx+txr0+fUM8XdMj4SlGX9Qn/+r46zya5BIt+yQZ3JEm
JbfzilSx+b63saIKxs+nCtTuk1PNJgLGxOwCRvYFkU+OrN8jJVE42VpWc/5Zi9gj
A/cUN0wgOm4X3fHQgwieCFhPNELiudc4vruxRwF7KoFsbpLlR1yO7WwscbqVs71b
/gTlemi1GKpBvr85yn5nhdXoOj0c0kUFCAlzL7eBFgDXxjyUleqqvaQi0dRItKB5
h9/ise/qlLRbpLR3+sQiP8okak5TR9ToEJ4T7Eur/3Fp02aG6T4yWvCed0qmneEf
iDADSxL2dDoH8O4676xwLxa6bhZ17yCiL/0PXmOKoko3QEQqhj7wNpAndpEBDKuF
Mf2RA6YferHK33rc02tLpkYBQhZ5PZDa9alAQge41SCJlsJh0lABc6cAahsB2FLZ
bEAinX86hFDwM7lQpE+b5UPPqEQvyllMqxrDaxNTWlHHZ9mHj9h7uGTgxlCcrEDU
RftXZagN6n3MbrnZ9blE+9qfhOgLzw0Wfr+Xf7TmdHEO4LV9Ik8/67WZT37SrA7+
9t8yDgidBlRt/ZjOQfCYqz74xd4Pho9FNVAJNkci1owTFpeY1lPinHLnNV4QpGSJ
sRn1mUTddKIwLHw6iQe6mi6fhHHpJClYRqNd2wfrAZ68eCJ8ODhGrQV/5cuPD1v2
pOdL6n1QB6RBgGFcU4EZVdIGBx7MN5n7XKmVCWrcLRRyfNflopEuGdMClvil7Ash
6mBL5wu8LEqw8P2jdvsYNpJFboBTRU5YJv5YizrKQJuXKDvV8o1xV2hbps8k7RK7
mvuOHi5d6OUnDw4SPOstM5kic0vJAPaBDWcxM7FR9hOTjTY/eVhKhDpXTfkZTU3g
feIJt1ZLCr+N4pvSFEsodxupdHN4U3tojXHrf9rpfaIZg01GyN8BO8etWmZT02hP
mkCJ0wxQT/JiF30FPOS+kfFoBgETEen1/gnCt39yF/eZzC17oXJNihwgXO1cCwP6
KoVLsgB6JnSs16FQhZ2EiS18FiiZJNSMigm+8SLwteGKofl5XvlGQk0Y6OGDAqbF
DGlw8Sw1akyOOXEk88BrO/Mj0XiSmQK3jm3PJ1XR2RCQUt9NSm6XgzAQPbFTQOdr
Es34K4gB9oejyrpoMB08FHfRcSy9etbGHzEE5EDP70rJ322Nt4o/pjhdfkISO9v+
hcaOglBW/fYqwyh+DdvDhiBHenkUkSZFJ8B2uxaFb3tMt3zPyMpVPyr0mtS/A/ZO
MPNqbp+kYj0HC8f/2xAZzvxZziElybMux2Lop+1hyA7lUcqMjq/9Cd3G05Cnta7k
grdqV3e+kibR27Qz6RT2ll1q9ikHZBcNr9oOEdAGA/lFvo38k3hUvcItdapyzQMd
X3Phbro2U/qy2I3qrLoANWGRe0s8rDHVmtqzPj9Ijg1XXsbodfiAzNkdia80FvV1
djhW8UpnswAIKr+K4xxOS2dEtQ+AUySm179PybIX8PZ8o+VeiOqeb1WHHTEdj8XX
s8789E6+/i4VdFsbaX+6pHuqGesumgFoK1X7dFrao1smYlIYpTu5r2M5RZ6cM6Gs
zqbil04nSgD6/tN/3NpHpspRYanRvw+oEk4/RVJ55rf5PkgJwk2rLW7iorzwq5sU
W2SwK97WITQBMMvh3x7TOznMVi4pIfwcLfj64OZvmKeyucLhzdtNH79ckc6IEp1U
BWsAYE2998ZMgssxtf6lJYysRYP8hYLTRl3qNnXIbtDC8ys3L6Xd2LSWVf2mtJN1
9XHXT+PS0d6FgvqdiR2fcVoWGOHVtOqb9Uiz0K3KSVTnSO1WDjB/dHBwpffOD3xx
NTo6M2fyei4N/JDUmdCCdkctg8PKxj3HhFSwDlUpC7eEvB5IXNLhzV5fTZ/9XZw4
eV1A4VXRgyNw0yEqFJGdNoqQmV3wvLe6Xty1o8E7sX2qD6WgfUt1Dh+am5L+Pwad
qQhVEVd+nT54+AO9T+f7Ru2wKbrqQiqDdktygdAhw2vN3oRkjXw43lk5Martmh8g
FRVMdt8Fw1zIpf5jdKq/+5V23BVifm3BKpm2UFfaJwgB2t0XZMWwCuRJMPVchtva
Vrp6AVDZWNpUP1GKrS3ttw/7S8+H1936XjsNohsN9xpYmfq1h7JIGrh9/CWWXnUg
uap9mE8CCN9rarukUqQ+fR8vX0hy9xWi804Ctjdh4VraDxD1P6OdG+3y+61b+Gmi
V1HNWpYbyk1gRzwSKsWXpI+CbGJUCqO1JzENNHjLWYMYi1MaiIlmwxiyU/8dHY1E
VZBr45bG6Wjl7kgfiRNsg+ZyvLIuQW67iRLGp9aRPoF+VjlwJ6L8+wlBhKN0JHcb
GeFX3KGqgAoO1meioBhH1PWFvjJKDWabm82T0h14KvGrhURqjEpHZoGk1Ogm6hlS
gfrOBEslDBr3PCcqaZMAurgBH0a0VKmK/W5b3Q/ABs07UQSaG2YBfeIs31WP3ocK
/UW2swAdLmEu1QLQLZ8ngiKq0Kb4/XiesftYmwYN/nyHR3gnE/SJgfF2ozkGn7KP
BnXbbGnwrLcBJNs0+4BUVc3A31/FLo879gi3J0ul6r2Xiq6/TypMOBUoPKB3whK2
1Bw1QFDvtSNomXxSezT0dZnSM6SC3R5sXQx4qvNwlVD0iiuRq655e7i1JZUZdTa9
auBFW9BqUffB4CaCcACKG5GAsvud0m5V1MN0MKmMPQCXDnUJH1B1xAzXT/+KCvaL
g6MW0kYQL4rqikAP9oXM0qy8I/qMaJVgsxXtvKJHTqdWo86+6c/HyUNWbtlc+YHn
wAEHn0oKyMhLWOu6wmkPC2QFQtvAQLS9HtEZ8GzA95FY/02dUkLrHl1VIC41wN2l
Q4uq8IAHzE8t5Uc+gUbmI320eQZ2qfX2jPgIc9EmJPvgUjJc+vTxdCPMf53I4xRk
ScJDjyG1DM2GrosxFu2iX20fBviCTYOrimUluLAXV7hTuipeAgVmBCbI3DgceVvJ
G+bfZqkzVdOosB1DblaL9T0O73E5Em8mjoaUHMhgV2ojJ5zFiqlwvof0mUmaFPM9
TuIZzPG/J2X8PY+MTZKz34JumZErerknjfadijxK6rgcK1cMY6Ciucsp2GjiqWj1
EpsuC6K6/Ha2SsRdIJs+RkCDNBJH5bhqGJjVfz4+sWZGVxhB8KsBLqRBixHdqgb5
i4zuuJvqO3xSZbXjw1yUtyhkW/kGK6eoly+14We7cpmr30/x+g7LCRNRNM8AV342
ULNznay6AskpYw2DyyNKYs6cL9fWWGEkETkcRkF0253vmejf7bZWfM4xJgxrybBm
EuQ7cKXl9LnplFuJ/ARpMc9wkxf23zmgtVUH2puwvBjmoVLVhbfcgA1LhGrw/w81
MzJTc1p0t9p05HZ/T+WHjW/6wfXuUuzPf3zq6TMSvl+KndICOl8BnQh1qgv1aeHv
QxIOn+ENwtD1/OKodSSrXgmCyZX1GrESsBkYf5MScObi726uIzJFG2HhpcVX+ap9
AoIFIQ2nV/cTZm+A/WkmOhbIYXwbwS5Ktt/bfkHdbU36FuBKYe0S5L/o8fmbX/KU
lP8Tig9BlFt56ZChutTWU1hjrapvoM28/g8aTbqwiiSrzMquC5AIcEhf7VQCylNc
+bM26R7waFTzCapEG51rKWvuNPudnpajf2oQlLujAPP9HclTjsMiGjAndKHljuKy
r0qZKuBORmlhpamxzbfyCFhf8rw88+mdIEK13URelk0gqxwK85ccyT7JMaDh236d
GjRIgDUkLTdCb3I7+Ga8UpshqZJgoJHqkyqBoNabmLMcu3R4yENGmcbP0VSrhL3j
avlzI1+q7x5yoItbWbYFHJJARXmGOcHIJU1uXp4JlhCEyPVE2hnQPanh8kjtIdSL
8k/B3ekd3m6Zs5UAe2nPJsdP+48IrNsMW857++ZufUWyODoEFDbmtHArY3DuJ4aa
aSPrMww1Eo18tbEY/XuXKj9pNDXWQC5oaPOMl+gk9N4=
`pragma protect end_protected
