// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
snypXx/debboDA8DZyF8zkd0Ghw4BWRVh7P+hnJzoUgKsSUFz7dLi9KAVimGggUlWhCwVpkEdtbF
J0vomfPoAeaSwDDY81xqVpO2G5rY4hM1thtNM2HSlAH3x5Ue9UYIAXvYPF3MXgAVfIndotr/LdpG
6tlFYVQa8+qiAlHWEj20elWzpr/+/yZMjx0QnXbxCFzSLM8T/lTNR9uN0q6KS3IPQjZkx+Qs4Ur3
sRanIse6tlnmsDhod86viL2aN6uy1hpmYYuCqGRsoH0MdrrxuiXkvCZ7H8Tj4yzPsathdVKczXTD
B9AtAK4fcfA60EXGo2OCZuAHV58ixd5ZKnxT/A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
e4GnT7qIYQvFhZRczfEu5lQCX86OQdDyUhHJ13T+LQF8k1xSWOWJCm2Jw+m5S9Vli+/UyFYUO7bR
CwdK2Flc4qhJYb7wXFC1fCBrM/YRZCYbuernUd4X8n6/sYJG93DKJr9FHLJ/1bMC5PhlxdDpQv3N
nBLNOmbON0e55yCEtl4U1QYYBFyulx0rohMx+8IkiSsZR+DFD5qO1QLY8fo9IfDFmRNp7rCCcQ87
g0CFTSW9F5FPK4GuyBwnhF0E6ACM5UyHkVA0RjqYgNI/ttsLOLVEm1xrxHQblJQdSZuwmmK7uueO
y5N4mqiV8/5JMIoD90PRc5Vi/VW+KgM0aT4T89F3sVdxCYB7OTPXSPvKRUx4Vx9zohVwlTlCPn0d
wfbrz8FgiTRbl64JwwOu3Hm9f00hUVbwsCN5UMrOHhVK+2lcC5IqwBYioiZ0ETAG5/ZGk5J7TeUN
T223T6dlKoiXnP+kBfu7vkfx5+2NRrrk+K4ftGtu1NrIk3SdPrq1+fJWxkKa4LOO2b4xzWzFxi+q
uhDsC5Mh4WDYaFCFgPawBT5oZP0s42H1uPLnp8Qgqkp2TVXKLMUGBzSKlojiPdOCh8SjxBtLRibd
TYFAUmUCByi9OC7OT3iW57Q5YH1GHHCHSys5kglIp3qEQN1haZmv81D/psQHKtx2oEjmqxjU3hek
vYrS/979RRvDORQyxU92wmfdMFtXnHWjxmSMw3j0vHCCqeP9qVq5xcpkLiTNcZrOQaf62Az8x7uX
Cml8FkjP6Z49mOPFDuRFNtw8n7prHZYWDw+zp5tQuJwcRzrMqaKuZekruI48wJ5nlORYDlHfeFRM
o4yrGNgxiMs+MkSPZ2Ltc0zbgMKs8hPl+GRyXYkkwstXXGxUz41KQe3G9E/t3CUR4Id7e25flLnm
5gQH3HU9PBD7oEkUXQTZ4N9YED2B/9zNgukqMFUX0nVt/v0Mtfwp2Guh0HFFo6QDkq8Q+qWuZlTx
EunRlIbNW1x7fjJdxV4bNg0GjmcwHg2DcGQ5eOSyj5Iups4wbYstz9mGQbtdmpvyxFMwKDiAMtzp
9a305S//ZBeqqaqYeyI/2tsWI9zFa+vbconJhHjTraRxn18n/ZTfdrqP0KBuTzjZ0v69awgn9F0l
WFpO2zDEhWFN9C4J1MwMNX4qSe2RbA2gej05zT5NIj7x9JX9rcFet/B5ZK0KFIO5xaaLsCXCvIO+
+7cPZt2JrY+o1xA980zu7mSZq5tJ9AMsF/fg0z5Oz+JUw6Q74x/jbnDxRPOtRIg2PDxF9wG2Awiw
MyzLtsw+NB2kk8w4iL8NwvtX9qjsrIhGtzNc4i7ZzifUrj57epWeQQP2RRrICOirhMNgFLx4Lejs
dZ1ceOfo4dTmFQ2i7UK7Allc6YkrInt9J6VsGGr2MzeTvcdpOPUPzI8BhVUyRncXm6IR60AlqArF
m2qedcPY60ETJTTAA9td7IUFCzYrQXyovGnhTK02iN4HD1PmOBQ55+YulKcPhsykjFeFurhMRaZB
Ci/ADTEqENlb2BaeTmjZh2xW7B5j/SakZBPaS59m3heuvmC9q5xP+eK4LpiN4MbAePm2lg+2mbJu
KTV8JhvD1VULv64qcmEiaVyG7Vo+gBcyMHjbj8LOdFltDpguXWod9qqZcp4BR40lXDemTTKn179P
pZKIUbDuTqBttwZZa1WtgIri51AjPqT3hKWWaCGgHi8dOaW14JAnuXGEszjdfaBFm9x5UK/Cuq86
xLJPj0Eo5wFNDi42o4a53PYHt8fRkyZaCeeiicJSu/7Tlk8wHQUyMFlZNXGwU6Vuvc/taxga2V5h
HB6vMulpNpl8G9DAu1UZr6JZjL3suwlkdt8IGiL9e66ijwnoF+2aVHumiRe5WqyXteGUr7RTSh9f
FNgYtMDIeCWqiEkLx0BiwiG4uDfF/tBmESaYsJHfILNGDN95BbCSDOwOJ1kkB9bwL+cv3G+J/jYR
G8Ie0If1HdQFkS8YxqvQcx3DLSipBVRDbooUXW1BanA4qSfIw/F7sA5EKLw1SZiwIl+FVSeTpdUi
y0lyxm3YIyH8N1IUnJU6uEogZpOER1Riqh81mxuuid+4K4KYcvKp/kaROjHGqgsly/QnsDgCQzuc
y+dKDh6MfC9BKZsBSUMUdCPImLhx4JdD95e1MJ5b+8EUnRbCq67frRTibdswcJyfsmNp2BJbATlt
cHz0ED/qp1bdlsXbk/ZeNoeFOBpikbBEhbATWSejRhl3ppNDMasVpENNI6hBnKVfdi85GBBb2+3+
v5WajZ4EIvsT766BdijuyyVgoM1sSrnLu1TY/oIMiveex6QgE6CrdIWy0wyBKW/DVYv88hc/Q6qr
F/4voqOxZgIJSfDUTu4SSoFbyWkdj1QdRwRVGtqHiccH3yHft6ToXJGMXQ/ylw+elNyLSoHgswxh
vv0l6403dEk3wxlf1TtgstHdjcItMbb50C4qG8jMam6s49CkMyqluMwKwyIBGnQDLbOIJuqEbRk0
xKNe4avYpy1ScyoVgjONKB+o2FczjLR0kgEJBpq/0cqnj5LeLFbhS+LdGHhi9z/sbKb5VUAuzXrw
Zp4mRXWwI6q5I0A9YirXW1sREg6T3z9jA0mBBeEd4ntzFPKFHKHrq7fXpgyRa6trrtpoftOCz5Va
Ro1iebObUr+lbnWQ9J2PiUxXdbBY7AlEBX2BkbKlVn7JpWYc/TOJA3u4H4n3tP/czXr6KMvdWPcg
+R0vvgzE6LrtYb8FpXWSxLGLHpBTZybaok+74UVLA0mXk1/peO6P/Dk/uMJDpK7ELlkJYqsEtqrE
V2HtNBMDmWsFRKS++VVqhKmSMoDL3pLYBqf2nlQ+x8t0xmDn5O04mOYySoFmOUQA8Zhq5urL9rGf
o5ne5THxB6pCrwCotXJVQHPe6+PqXNBZZ+Kj+f3hTATtrPWXTW0BPyfTdlmnWEC5+7TvqOMi1apZ
u5omdzr7MKgKpBese7EjT42TiW0kwQXvzQxObEQH5uNH8C/c9hmz57nWkD5+W9nDbnJk9sBqux38
peHENxpVX6+T9GHfPAnuSBCEgR21pVc4s7hsHQwiAXEHhMmlbG/041UVYvYp4sD0qZuDr6FQ5H2Y
LCN41P1Z0eug7Sqe6k/E8DnxNDIXCOBdH+hmJgzfzZ9N1NDzkuYVkG7+zxe9lPWhlRriRwfBhdPj
IwG4UDI5SzohkberF7MOxhyBksBdrxlEobzqkvWiiPGgSZ4f3he+yMStLu80gIha6hqRwhcOGyWl
Ph1HXBRx3SZ+5bSmstcFvJyNSc0hvM+vNJh1VpdudXs9QFCiJms7N7o4nKsak9/riFFjBDje6LGN
eQRuwPcCe14keT9ilzOU5cZVUJv0YaPvNj9EcvR6mY9uahvsPfYqfZLE12JwX5ukr9e4XflCYLod
z0TOvIvD38hiQ+K9UhEpQ8s9ksJLzaCY3iCHx1SXaOG6dBuaPTyjcDIcnKlGhzCZmnY5RTzDU+hC
DkVsa9oSlGy4/a2eOHy562PC58B61fKKrPmTYG0v/gfs87Q4DiG1GZQu0Hzj1adwgL4AS5lCSlkN
GDhtkRuScvmdRv76OiR2QigZUwp/A6Za5J1P48r0HL53NwM9JEtROqx31RIgmwYW8TIFS0gB16OC
NCWT3nFKMWjmA0iKHbQH/Co9pZtKdYYd9w5fV2dB4Veime5/NPBfL0OCc8A6r1pASfYHcpzeU3lA
tEr1WDVYDCfIr3Raekv3CYNTz+H5Z8U0SZHpxSWuDkM/n4GJfR9rJEQVb/SIKp7ydAqMjnRulekB
N3ECKZfDmw3spzr6D9B+j2EzmSBVxuEkI49eRW55Rb/ff3PiOSqSKDrhsWq0eqA4uVHYbcpYu2Dd
Eh69Nk9+Ppvb2mr6v9mUiwJchD7Lzx8jBI3o/RGoYuoTL31aCZ4OQW/v8XKJY5icKsvRiPpAmH+K
ITyRvKzZX6m469wBQ5kvQCbXZfo3CtFYy5GFusVe5Na7Z2tAL2pPmAsrHrWOH/QZYVyiRW9ahnXa
vy0l10IhqvlUCfRoQ+h2xN5rjQxeDcFtTvjQ7te0Osyco6lGqLgdTJeifKs4xrfnnNpIg89i1H6G
C+PcUHq3WgrpIKvLXI+4fx2lPxbFIgbf3RBbzjxXLh3l9vKUd+uP9su8DmJ6tmXZXUEBU6UmDiA9
MfqKdIQro4nRazPCDRwLoYX+UhaKr4GNMIUr1uqB0ZA9czWMTzxmDHIH2sE5ffc4ykHmMZtS/svq
T/cgu5OCblhNgRdYrCli0l7kOckrRG3IjADdp980NZpLoxkF0YhoGJpee+uSi+5bR4ZPoWuwWG1j
hEZNutnr32cC4THYY/J6FXKtUu6QSO2AIRzzyVhXW5IugTLQsSFe6skyGiMLcwEduc88N7RPZJKf
AJp0q+/YQ61MgaUSgmzeuzrcp6ayNvuaFjAMUPvF1gh71ZZMULCcwRQaQZv7S1UUt6weM0bpc5ae
W+Zo6VsGkW61ixNz7j0uqy13e0ljLQrNXKIP6OvJ5IIRccq190QUlHejhExx9Ro4n0+zlH6uarm6
MLhj4HlcKeruLNxWiQulezfTz3vSKg3IfahXVA4GEtuHcGZf5AIFr5oue9YcY1kk63GbaW2KcgTz
MPIDyhia3cePGNUuSV75098XWwu5CDv+z5FXf5A9VHVER+G7uI8mtgafT9n5iBepdol8kmul1fC+
Prrl/3gSXwft3I4efxAMzRw1a8PAWHeqgYedgBB/WoBeMeiD8j+i6suyBix+AhymQ6ehR5Zqswx9
OzCjDKfFOvmQfM7aUFY3iorZj5lPImqMRDeWN+ecjCjzu1UaXliSswPBEf/UAnYx9qW5HnrGjrN4
g73Hy4Z07/Sctw0YIMWX9gW1YYPWZgjSaBvT6y0ei51Z4MRf/fmPJeGO4uRUJuNxfwxpaFLaNA0D
xhDTEJdux9/8h2+netjszPfH6zPck+tE6QOmuV4CS3F2HrQC84QDts99krYi8vAvdO1q+yTefcxd
D4BJYXPrqwIi9PTlGEvRwnyqzmFNbWhhqJAVGtvPYLGJ27zwBZvNfEaMEsgyd71yMz48cf+dI2zG
pqa9Q//l/lc9UC/0G3cQq1hFR+ZTSBHHx+N7cZ0ix/yildV+fWUdifmu2uoNFDjMPYlvUcfOVfAD
w5c1KWkIBiFDWvV9nYflflhKp7VQSXdhUlnhCtn4im471onSzuYl3cReOxeFZ/xhqrCims6yqk4j
QpG2/b3KtjikySzt6ES00zP/sZ3vw3nZVNtd30HYBUpn+KxnvSy37icTvNH9l9zjp6MQfOeSwc0+
GjrlkU2wMkEdVYRVu/vaHt2immwZqJPeEuAHUcS5+t1QmcFRwv/FXxTKb8uKSRBHqYCiEtno65kj
NVVUCK+eS60OvRKlztUBDHilLVHvEYWX0EeEYagxn/T0aZ9P8iNSoU/0f4ttRoji2jdMjI9HLlF8
evWKugujqYN8cFclQTWjjaVYEuVXoRalaS9ptFIWZ3BHrP9X/Qc2QtNpuH3jaK0sJb0WOR/pODtY
hrfG0x17eD1vFsgNBaGGZpOlqDJu8AmZcjLzD218liYiuH3zj0ttewjqV/5LRQ1GCdC1GQwlm4Z+
uZxVl7LxyZFvo56HnCTzKatv5VSEi1T0l6yBIZaq7psEtI+ittnkclslVCwyjjUwIBwqepT96/mS
DC8dPKgHb5Rm8WQ5B0EpbLf/MOb9KrbbTBMcvQTYkIAirfMfCvHPcSWwENank58vOcfez6HBoXgZ
2j+LvPC6zy5XvGyJzmf03s6gmufuescf2FVAZTmTrdMT+XoObniAZuiVvDurWA4EZIf4B1jHG8HR
mB4K+RDCjnc9D6nX8K5iCkTLu4qilOzhQW7Mj8Gn8JkCt6znHFPxoVJVDkfi7dk+evIhlWscZSwJ
Ru7vUCoGnpl3DsaIxtZpSOhYCaE70KzhbfXmbBypurkB5qBJOP8F6Zl2JyVpjdCAs8je9hXNV+vA
GI4sCEIooabplZ+4WeCu33a+xucGS5CoBUSURmQMtc/yqGKJyKwcx3Te62MbN3x0EIEUr2sKouiH
vv3kDa0Klgjdl7i4iRPRB2Uv9Whm+iPxLk/NwhFDHmRjGkbrLjSeKhWqrdfq134wWo8o5cezzG8m
TJQDMeAqgvUGWwiFl3Gv4Jzvy8XDH9u1mZhlvz3IE3K2/J0kEIF5VlRG1ba/nAtS2PtWwxDyAqDy
tjyejjK88ZTpqS83YfQ2gCxE5F6knkK4lB58gSDnmT581llxyCF1cISQbbnUtcGMfJdB4ZRP/1VY
I0/ZQeeTWFhxNFuPrCmi9HNzzMeVcrVBwpefkBslJbsrst0hjEcgaDYza3TBAzsNTgODThoW2YhM
pzm9YS3IvAp1QMByUSBEM9aVcV320P/Q7iyNKtijaxGpsH1I8h9WilpUg4BpzYpe1WnQP7OStCj6
i4p/RLKr+0OqDXrslJiOiwvKHLzTtEKdXwQfdhmn4or6Qe8x0YKbLtybEr/GYXIzTE/RmP/w2aQa
AkH8gPthMoDSomNLYXWlqr13N30pDQQ1JMO7Po/S0zmLmWc4z8FMyQkPGIChAfuVWsSqbiFW1ZVB
x7+s4cGRaddNzyYt3v5Rv64WUCd6ooygRi6CQHU3I5cQc9PMrMjhLh0Km5FwAS5HmbuModm7Zmkj
N0e7Zjd4PAy1xWbz77xI1CXAkRK8i5eQ
`pragma protect end_protected
