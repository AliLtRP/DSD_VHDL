// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
aUIiXlP+9YBn8ScABmwRrcFOHoyQ17H4C7DDoyaXW1YfDmyiHWYF08JyebrDinB/RM0EzSKVrCgI
mvVleyr7O1aU4Bnd/KGIgeVL0YR1HJpQN4OlMr/vAM+DkyW0vTHw25uEm7SpfpH7ruZkKceJ0K/A
/QI9+juHUHqRGtiQm+y8oQN+kScA4tf4PjEODMos/7alXEFjivngcmvMjWZ7dOUU6tnvo/6+ceiJ
vbWwJ/wNVGfPT+AvGYEPEN6tgsLAOqNZXnbJx985zePzG/Aa2BPnusJuLzw3zOX1wMOC82Bnkwb8
rQ0h/NzfVUWNed8hW6KFHeXIG/Jzkqsv8AxPrg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
V0YO90R+71jaxh1hxSUoTIliGZLuPESdwQ5GRMbWG5Z0hfjwtPomT5BAil0qsYZyvDNqNtni/dl7
1oARiKCTRO3g0k2BBlasFKD+dZ6aO8dWKPX8FQPUssThkOyIYGDklb0KRxQLk2Zzs7gocGVXcP6P
VTyKyzdXifsWX+b435gig0XjkALs5ZTzR5SW49oVOVRKedVXLoe+VxJPLfIm9s9XjDXuz7JTck05
CAQ8XJvgQW/x/mEV8kZ3WPGuvJnTPGLae1Wa1qT/Gi0XOD1lHrk6zGrQp8EfzVGAz1/D7WnOIJAP
k7oXnLf7SXm6rnH+x5iDzSAh+lNm+GKnDbS4wuNm9K16IUFjzOJEA3Ev6fyr2pNSgpHa0mfwfWXk
zQmlzBEbLuiJ8vPXMz2TZZb5DR8rn1MXDd/Gg9pX5+EIvf9CIJydsoGDCe9nMExOREaPWd/XlTXY
jT9G9u5IxanMapYG/0MAtsLav9PkgsHaxSODG2N0yhPI97jOoQpjYGqKElIX2+zL7Knte2KNYsTd
wtQjubL2d0alJWDRRsexO09pyVCNXUPxgYFSEWkOPCvPRt37MZWmHQnw52IMqba3FUgGlRwydDsM
uN/pGEDd3SG81g+74pgr0jwogNUP0Zy4EasKdoGWIQoXoCgCykSxaax9mLPNK1PeDxg2Dah94oqJ
f2c+TgQND9siA67JOQPCLJvGIEJ/LgIiNEmVGBTW9ihAwcs8PmiwBfDfwajGlskoEJlmNe1qrFNe
8pBlthcmDhHo1f8itV19eJ0edqSu9dNC7balY4DPxGNqjhtNZ5+j5cmr/4floojE4JW2R2anOwVm
Sa26lDpTy/zRrEuNaPjQd+LaZC7BddjFBaDM8y+3PKPW4b0TGi8bly0opH4C0a2Hjf/uNiNTBtO9
yFr7T2YpaHEf0ESQ0o7cf3qwfQOiZIKU/NxYp3uGmEAk8l0UPuHMEMjyokxIujkAwTziXMMWwOx9
TJAygaedc8HTiKLYeaQVoW4jyeq3hNahC0Bl1PBVQTJCWi3i59PfrXd7MIwGCKnIaHRLikHsUzpF
vwmgpEC2sA2VMs1MAa06Ot+5PnQyqHUT5x2s9cfpjUvwLux5Z7wVz3XtRv/lu7kuIVJKIPj7JvGF
EHtkj4mBF6Bxwj438dnyicv8//6HGna4MZNPpazSljI8DrUE73+EQrUn4MCKgVo3jXt5BJr3Gl+U
SUO4r8LAhKF65SShBFOleyTvXq+GISYJqrz98g81ymmh/favGqW0ZYKXSAdorZ+25j8YioDibimH
29ABg+UEHLDaoWe6SgOXkjfQ5XD9mSPIOWu/G3HIFxNVoMUNbH/9sReTK5eHfJbfxmLBz5F3Wq5T
6IfWJfyRqd9X/wfx93tP2nJZo3wZTVohvFLj4Mi1zvTrwwa4+MxYgTmy+mXfgdZewfx7T2vsByjZ
nFznc2sj/A+Y7gVGJeF3PLXGMCM6TMEu7QhB6jLeSWi/iyz95ZTZnx+tdrmeIW/X6805VtOoVFIK
kgEi1jratPu0X1yoE7QOx6rHDWQyuU2LLlxecqLbCrpkX8TBLJaG1WicVeI29rgVSdP0Vecp3Bj+
zdItg/XXpq5WQD+gTFKOOi4Mp1ckbPQVpG/ewz/czh1QI1vvea/an4rD/DOxAVt8e7fSAy/FoIpW
lAWHfP2rVI8w+gO17ytFipaXZ/hh+8DreUfumqshXkga/aY1MbQKNShuulM7WtGmsJCpROLyqD+C
3CPz6QBR85856WkkOfdKvge2wR83sZmUhbgxyvbV1f4vEACMY5Y5CCgIXPzgDTR6jwqU/YfAD0ir
rqzmrMfoWg6RbscO0YBvqPOdrpR1PzthBktWWiTHcFJDt/iO8PAf7qa2oEX0JO5uRo8B95kyYd3L
PaCzhnLgQbKFsTUAEYZbvVaraXHbqek7WYHgps8dpKPyWNVdmJiqyeJ/8B5sGMkF81OwtGjzIS2m
ZkLJebfbWfckzDFlWcvL1JlaCPJEi08MaFNo2P31SXMYWN3mVlOfw9mCHXQnGk5vfX7Flw6aV6vm
Grh/h6DhoWFIk+SSYtDSN6OCFc3jTbJCpH05W3vWgNyMBykRqBn4DfcbiPzDkHPhA5vmHKIyGnGa
N3WXFILTkiA5QXDdiMs6OwC1CqITcHemWnPc9ynAOyi2qw59fpnwiNBW1e1uwXRsyDYHlTL875au
aBwA8yHaRBEAOaTyZLix6GoTZ+kJZBcTvMKyHjBY2NHKcMI5fOlStiyvFwqFFvgNbwRop1OaWdrC
SHX3vaf+hUYdtEfY8D7BL9TRan+q6DGEJNWumnzlvL6PyRep0FFpZLF8c747HRtHIYhElyDf0brW
gBWpoQhm3/F1LeITRdCLqnjW93SNrb5lE323f3cFOUCJ++K/GwmPj+hdqTlKDjAzOHAbgCSG/lR6
ef75iJM1u5/8oSjct4Ext2s7oJ7M5fQTasXX7zRW6UXomVk3dKXQcqCMirYBfdAIpIRYzDNcke3T
ZSy+hHHqM2QYVpWc0NrXMTEAr0WhdGgSMp1mKNKxMxvKyc2JUXpZGzZ2taSSbxcgop/R0VzN4hjy
tJv3szVeXKbrAUnanCS+bi2YBbiV76gTJLdj1VhsvltC5LJGwDaNEk0CXC/IzkXrfIEDKEzECMSd
mUDGNGh+BOumJO/jt+Nh/nwSXaJgViMWD78zM7+oNTR7OJp9uTdjuc6upGwTMMPzzNLC/KSdMJ5T
TqA5M53zc8InPoe1IksMBMfTkq+wPfNSt9er5EYrsVQRm2WYR6AsBWN0cjsd+y4jyfzqJSJS+IfN
TjE//4a7ytjNAcqkrmpbM45t1Sa4Di6fVurVoZyT6JIm/4JieeIifnbnToXEq/vyzaplAlS7Dag+
uJkyQOWsto4CD0RLOm29hWNfQ3htqWduMeVZFAANnhFvEvLmryyA17m/EOAlfLwooFv8PU9vapyd
ijx7UFnYYUdVd6/0a7UdF2bZyN9xNbLzzP2LNTPwkZdW9hyG2c7VaLgS4y1ArsX0v61sgWhfjeKS
/jmlrALjGxwBxbiezKKzOYFNZYWosRPjq4dvSxDkDt05KD1fVyNhb20JDm5HC3iGWt7bapo60ufQ
nTlzCgcqGZB2J0Hxbp9rwnPlXzkuBoDeEN96Sc/+9IFsVBPfUv+OJ8zEuIyFCqY9ZgfCOP72oNL9
SO9xYTvW+sLPSPkFWPovqFsFNuEikMeYBdKYwDVxfHXkvqWp8kbKq9utkQ5oyaJzLSJrN0HiUxym
bxrhAJ/33sdZwIQdnFhOd/yr2Yv7LFnfSJCVfAJORKqYHjK1sgxJ7jSK4IWliw3lL2oIqSJ2ADQF
modgbBoO3CW8jFzvyhczS0YOJuEvWUcInWS297AOfzvgUtgoK50QZwGQOx1jj9tF8jxcZrM9koxI
0HuvtRYY4whzyHW4j6jSGTwo7Eliktp6M9ipKo2diOefwhC6ZMxO/jltE8zF06kJkr+tMXXXNdY+
efCuyNL6BTAj3WQWhFpewJU476K8MCv/IkL4oOOB14HrgThwBDMqq4dDpyEQvrL9k/F/bqSHhofV
hQpXZTyRBuI4L46SCRsH/HAYkbsvTQjSn32sFMxtWK/tgsfAqegVC4gyck9U2Kj3mK99SzE9sdZn
CXWSL0/ghj374K7NSqfeYt3VRJ8Nffohp9buxc6gzbUdLZKOFSNXBnepO0G+OCYw4L0nOrx0ZmN9
81g+mPId7Nqc2YhceJN46J4jhUhTFsGC6qQn3z+vmy92c9p1nFdMJ3ggwc9D3sp8a/GfSwEsCEfF
8Fyx1/BxpDA3qalfGcfHRzO/qDhNUF/ONUV2Bp6s6nNegJ5Ym7Dl8D8D/zGDVMG4ahdlFhkxvKpM
E9foUNSAvGPrRzIu1ZEZXT53bFeJASc7gxVAnS/0r2PEhActMrmS98de4ZgYaWRDHIQHCcgRjn5s
FWPnq/GVvuWezNyc0e0uY69ONsTGcmw81pimVIqc8BgeuZCv0nqD1Ij6Mad/2yctR+A044DTrWo0
+21or1Lbrf7yhjyJG4wEjNoO+aLKZl2o+ehwQ6xD26yJgBf9JAjxbxjbCKqo2VVN+u5Yvf3YqxID
2y0Whz0TsQETsz3/RrZsCwecQxLWNvsopS9MHugCKhitJdYu862geLmoubvEF4AYPlsXSh+CYUfO
gaPWyXZ3uooBUECt60J91W485yGfW3uBt5Sn6bZkOXIyEELq7QcvcPN1LGGNRhaufiqly60kb8ta
YT2Rj+v0RUVUfhAUMv4ZrrnJWVOKLybNFJzoojkCBz2ANTm13u9CmdNZyS8m+Rsrxs2y41dTwdQ5
ZxvONa71019IPloAbsl4v+gjNKXiMJiTVJ3ak0XrJRXpjE9Z377/gUXyDW9kXlondHF2taRHG/p+
Ga5ThV/N/5FG15CDH/8OxB9WfzYMCaJSOmc3rRcEd//l4YqzIwRQ3pzaJcxa9Ge8nVUhwnSgigsY
yKKVjzZUqioZMgpgyMkVMDequ88QtTUkKxF2httZEOErZOUn88yZg66JMGLvuQ2KK0sVf52QdYI8
NOjzH54xCZAa1dnefm35ZASTp1zhLKUqvE4pRgX2HHwwH9JbEuvTQPH7dPYo+A/Mti5y7WQiNB0c
ygaBVKkFK70YGmwuH6wJMIfJXmHTY9YMjoaDvfRf3/2cPE3Mxu0q+8RrR+s7xz96zdptO3frAy5d
z/TU9aJIyfAgVdpq6xVacOtMBHOTAdfhil5pERCCoyqG8JDK1P5+ZMP+v5aBrRr5NI5nutUOhhRj
77dVFtpn9Gjz6MkwR99yjUwk+2d4oXZ0yifNVQnrCr3oiM5NnpzV1RLOWkBzgZk/FArdalq56EQ6
GHmodDKsMm8AZpkMvWfkJ0lKeOciidhIGlWVXz52aLy8tUp/9R67dsEFn7CFYrqo9mclab7qJaCG
DstIOTBMYfWtU3UD5nneRwBfRdffPCCR2qvWs8Cur8CnSgwtUIau1JihIIba0wEfSFJCkd+dw6Zt
XwPJWvsCRBbg79VEBh4RNUAIoAZ1VO6wEJOjPhLNEV7kF57TV5gkxxzQqUrpBQa6dqjdJLHlcw1q
Ji9GPn3ZD/rHKH6LfGkwn5ItH7OcSKkdDgp6MJOGZx0Yq1rEJTHiDYe2ds+azKexI7VckMORH9uJ
KsUVnxqushLdfd/2pEVhVB2BJn9tx77HOXEeFr8HguhftzwOCm66rgtAWCiyuLSSQ3iqaEEKKGtc
oFF5YUTYFtZSg9n2rAxm6dODrRzADV9yN01lHNbUyhCJKDsX+SecgV3UscHGLBfhosRETVS/ZCzW
0EViwdIzncTCGOqCIxjwvL8W0kuOqquzhoWeY8xvAZfSHDXfLsKgCpGTj+CF7JKgvYgB1bmqXbZr
+eED9tesk9lSnOUaR63CPa+soAfBmv2cNjxd1cLjGFispojBWPeZk6lqpVxfv25cm1ANJwKRvHQf
cJIuz8kLT5nK3tJsVk1Z3piAistBxGrvrvx9avKGCMKIRphuwLHogjVJZydZ0vb54+U3A7CWNRBz
26d8EpCOb0lekn5gdxiCRXsggqGG/bmoKBMFJNYJ1+5Zqx+3HK3xiJgZU8CqDTzpvsIM8PmJMcBW
jSdgtqyqhpKKv67nrWY8mKu/0y9dvylHBvH061YPWdpFwZXWD/HoeAbn3w2VcK+1O5RNbtuQ3de8
VFh1wfeEfNTM/1YNi9XrdnZNi6gnKB6e3u07aqdg6rVzfDkW+unV6oF2AZoO7+ghQ/xPfQH5Qblc
oWq5T8vIpMtVsP/SLVX19vBi5q5C1RGMpQ6rxca2GPBhuY3ZaDiaUtGRNFpPqOK7xMs0funtq4wC
CVITwLuhqXZFEMfA4G+d9IglJsSTUgmPUgFZC9iGujwHuhp1lcu4bFV8pD8NYdBIewEim6jrXWdC
7gqMYj0GJv6PBjCneJoz6jWqsT+OM9v6Lt93QOCKeOiBE0cJWP/N4R2ywZylCPGVbATwQvQq59R7
zdcaVTF2q08Ly4vxy4IsgcdxMpY4eBISdLKTDtg4+RHK3EafuEZelqD4t4KIlh5RuFZp7pEjpAba
d0L7kBTWsFkQCD7OYd1n0LCXoyyvblpYc9PwPoRsRZCGXfLVXAhYv7VvOrNPemVHP9w6IsPCspTj
sVKowQws+GpWPK4McUA6P7OQnCCKioOP66VHjhtjtkzR/3O/w3i0VTdacfbxQA99Qn0iZHr3EU2S
36LompOgTNerBJgFJxIfcqc/AjELOrwrV8wz38FsesgH9HB0hfSrOYPaGb+smxOJbglGMrBI3LZr
or7yodqsIbJucstri971scyLk42v71BMLeZmxN+B5iQM9LtgQhQ72n8KsbG94NSUiRzHxAa5dByS
3NNbLOAHVC7E2sYvr6+abIfMJ1lNHFzWvW2OoxZBQXJNz5J6oC/6eBnrF5NMV0k7kH2zxKJfyLfR
duUK9t9GdbCaYs8sQjmt3u23FSJM35xA7eb+6tm/yBhxNnieirdCE3zM9YSVxAHoNK/w16jeQpNX
7iqJmA23FsGKYDXu1pVjk3+os5jxgaoP2uCgDVNR1lTMv2QiFeyQ6i8yoR98CzKPZtz9aj0/ulNn
x0vVDkB/dDpcWsx3lboroejzHwRtAiDNcx/qnh4IxRHvH3PlDrKsoJtqgovXw9cSJ63q3uK2uLcX
E5/2Fx7UWP2QsbIKrxyAG4ZpCvO2FIB5xtGK+378vfPkKVkhlKEvmcKf46dU3KiZTjmCZoEj7PhY
C3Avobnmv++CXmMeW2aY/ZQU+xDF+NrZqd98bv2Mqvw2i06fj4apHsRyWb3JcXhW9yMH/TUhtb5d
A9x+rVPnBbhtIY8IWLCIQk5d5kBIwZ3z8WhmJjh25lS3XBjszlAQp7zXmXOlfztPHKAcHrpclSMl
NVk9YoYaWlEEJhCayLVXHlZMtr9W0wBJETIzmv/a55fHHipCZbdpzE0ZB3zC3tGXlVOWlMawdxza
adQTSNAOo90Nhsav98AYKhh23PntnARy4Kuosqs6SviK77thqEbuyTaXy3fOffTwzjfRTFdM1sNH
cDdys0jMK9e0MOkr5ygPkw+SZ2ZNCMLQgiIEKFRLe8LP6qaWPcNdvypMZy0lwBNw1HO1n48ASKYX
d+7ek1koBwJHBBEO803hHdyJ4iVz24JnWblh+6Soq6KTM0MwOswFyIjJs2nWaRxoYYugPJlUWbdg
2wQ2N0J4S3S0szu5I06OZtux4DBMnPdqut6R3ASLRzDSd5dlVyebh4LIkMyoZuQ8KaNhEXnDwJkU
Y/O+MlDG8RG51TtGoZIjgLhkQNZ6McHT4V+69lgyE2mRSXox2YyiNCGcG64uXe3H+kw3Td/Piks8
Nf6jtayi/G/W+UN5X+VcXU1tUguw/e/TLrPA6L/A2H5B+yFbHEAtr4DORZ4YrYrv9DzPOTRucwjZ
6mHR+UT3QwG9ISP3OEKSk6BJjOvKCxI2NJegS+pslf3Hju9KXHS2dRv3LinXM/AHum/BZ49aJF+f
AcVBxVAYhSynpm/EgVfhUkt0xzbbT4Z/ei7jG1kXqwxnPFhy6PVFRjkR4QNXJjCbZ4icAFBHsY8D
4gHfLvFNm6M2msld8KgYVC12SSX+He6CJ0/wT1CrsrehPc5eq/lyxmTZWdJPPmGxVHKmYTbNsLMd
5m3mVlJHbhytiVLwoTg/6F9Iif8ncCGryAHmDyDDECSy3vZ8nFjRIKgx6B5sUJ+4/8yF5v7shv6t
Lzfr3xNwQuw9CKfCAfSh0UANWfeW1vrxF9Mx+9Hk0F61NeRld5DEijRfMXNGuV4okO8oceJIG5zC
ZVj9SiL2NZkxIfaJAArsLTlk0yR8uB6fM08YIrfd8P87eqBWaC+GrYqZWeEe8CWdyi812Bg6sPD9
lA0dGLqGqkjEeMWMh7OLc5IWunKXoOc2XkfQ3mAS5p8Kn9UcxYuJHhDTzcO9SVnvfKDKHj4Ew2A+
wif+3tiJfL+tyLpCbIUc6Zx/gdyvMrc6bTfJPPjQFq5JGERsM7TDf0ocxQwAcxPLvwGHHaMc5dL3
zZ9TIXuFSIP6uoMBA61nCKLoRJu4v4zmzgpiQQfdbW/bPfasUVAmpo0xoc5sUIVF9QEAon8/Cjgw
G8zmTQeKpiCU8AIv2mPnFYWjECWU9zq8reqnvV00Lq0dbiIXluWgR06NcuQPYS+3OoN2jul6vNuM
QeqeLrDvhtBdch0XAapP6Gf31QGj7SodnqyJcJmjoRn9fKQoQWUchGwdUJV3V+5gqnytyM+pmoJx
0zYFz8H+sJFeOQTYNINdT0gNiV13nYY+oqfiOTXie0PkCVw7OQTn1md3YgmH0GGWz9nTMq4fSRZJ
ZHSnvEsRab8xn2Z1cnz350wQgg17f5Sl307pcScmRJfDe8bmZlg8Qe7fpD9S/qB0wXjmbulDIqG1
h0XHE9B1bye5MEgc/e+1e5BCFrSviMPi3NHTK9vuvbsRzlsp+xZ8tlPmECtbxJDzyn5q6gMWXLDK
2MO7CrQzHtiiImDgjvJvk9ezYY3nnb9e2alU8T6T4uTlg0vPy/UHU82AQ0i4MckYwU7KwaqwPC3K
3M6LhzAPhT2URacE6ri1TPkDt8BIJ/H4vgnjtlIFABG7XX8Lyn6rWTJWmfH1t7g3zmxDE4huTqU5
iDSm3s1CS9daxPuuiF11R+9H+5yfl/gJeqKMgh+/79cxQYVrmdKRwhQF42x+a3V3iLNoDG15MqCt
FYIHJmxo10x2t7+83Un6zT47zR2/gcbqJXldSqsWB/XQdVX9Rmm7ZHVe0i3UgJJNsNKN+X8Lhf0s
VGrbMOXEAG0wOjpc32xaV9mMjDY3plTZ5yAtEXRIS/zkjo1pWwPvcenjpdA7Ab41lsAiKJ6zVjmH
zlODP3Ypk2qRu13KHrurjPusQOPEemTwZVBO8+p1tB87POZEJPQpSKxyRByh0iSoUPWqss57SmfB
J/F2Ila7KOEyH5vZ1JMJTVtRpkBSl6BeWVu2ge+Uyu3pruF5fKPiScn928rudk+t9JECYdLvFBwV
opAPqiT/IiHfAqtjssG5R2+ZSWWntB4gpG6+OutagUBxMrlPx5jTF/ZU1vK7iO2JHhwjR2wO/BZ6
IcbG2SxtXbxGLIlA1QSOhG+OCpl23iVXmiUx2c1PypiTRsqU7UZXWHI0jeYoLNrnRxAyZ1F0K6wS
dBeBPZFbiowLxF5El8oTJI8UVr3/7lrWm2RmxBCJSkWzBSav17nAfzYydJzSq88aayRUmEsx64pU
5VCKA0eMxIQkiO9Y1wKyt/4qS6tGzVp6YpWdzXf17RbmGpCnfrVCTdKT4EeZY3QxEg+M+yhstdpZ
4pI9WJ2EJwT9D0MYtz4bRXBib9WMc6WjluprEyzMgM6A4w7GMkPVBT3zJr00R7rzEuBLD7PgVoU4
ATEXZpq4LOH+FrYhc3qX30F6diD3DFMg0+Za6SiRW084O6uggFb+qnKER25VixYJpanA/XXERIyn
fYHVSZk3dtmLG10rXE8CG+kliYQr3kzDRwmtZVpHIIpBhdYhwD4mBpOw016McGBdbPBNJVY6GXxv
ScTJ9FLYYrON/7gNVHxbVbHslXFgXAhQuTKCAwU293/Y7/xyAI0ATwJKstD6DZ3JamZXP2eB7xYN
qcWFzbtWDmsJT8exNOjbMTarrTymIyEFqAQmnOuWENm4gRNWTxvkoALKJIIAhX27gSmmtnAj/luc
UvjM92HQI34mJIYDYqKgXRJgekGWNikLoI3X3IlBVm+uSPnsYg1+Jgx72WfKIosE3al+s3485ldh
nHyBDhvfLuOeIAC5N3awBT8ZUkY+anVnpwUhNWhvKZWLGeHsr/t60XqqtyD39DJvVzR/QU9+ddXQ
ENczXK95LVa2dnvSiRY71ilsipEHPyyphrRyKIDcaDUIeBQKDBVp29KL6AycfcRCGgKd4JoPK63L
TLdXEuFkbGvt9xu2BGKAdUxe35qcb+f5u42yM4wFP9TVoard1lP01kHSQIdYSQWeJ5oa/8rC8+5u
EKbpD5Vh7fWbkh/RGfsDOrdCf0Jle24k+FT+W/cf4+7r88p1StCP9of917Cn395IEbhPef1X2gbU
2J7xVgfKynWtCKHgkZKhHbciqhVKSWdizcReyA7i0TikHQ2/1zbZbE2iGxVJzm06Ro0bHOSyS6nc
VbdxLf6FtH77Z6Oc9zIp666f4fKF1e2WPYJEGw0YnTPRKlO/pQDEOI4pRS6ppw7fcZ2CWLyBvENp
45qOJ6+bwkLsuguh7v11SSU0AAod2O0z96hIG4xoA6sxWFXM7yo6ai1ki4R96/JdUy4udbVDkLrE
23eF9hML33cyy0q6vNWnifGhYyb4qnU2A334L/lbwL7ZXBqDllF3tHTdPmDmobaO7lNNSghGumVm
9C9LqRquEOB0UqjcxDqKRBWtFdZFNHJcjhZ+MEt5tEG+ELHTPNYBsoEIAsXXf3ok1AxM9lAuZYpD
8lBIyoM6IkQkwUUN/lpou34ddE04dkSpzF9o7eet0ik0ij429mVfdVuAxLTA62qH3dKtcLYQQv5A
swwJTCBxGNcViuPEEREVnqlR9KCFBPe2ZCQwnj1ngv0AOwANUU/udMDjCHjvhZlLTXpnLK5yERGI
c2abFQobvwSyV4kLXL+CfGBykrFyc8pqzlx3QYhHC3Cv1BdV2tDs4/X8IUOfVfnFeIDhqgqNzkei
K9T+7/IbB1ea/uJpItMdidZiejNVGj3J49FSmmNvaXw0W+7OsOpUDjJgsvhMuZkf3dMsfgYxyase
ulO0uvHn5NrKE9wi8URTd4n3yD2kwvoGoLyK5ObUswJwg3sY3Pl/uLYpaeCm6oEf3hNgDZfEl9/l
PNnyCaBg/1ro+KlKa2PKw5FmMz+N1Ngfx3XtdLyTS7jqBvLhRr9CvGeP+cCfq0Og7Ue6iIyGJQDV
/sZQtxQULgEkaUXf+0pHV2qy/LqxSk5FPrrrowp5KvhHHYkO6iSNd6/mzMVmLTl0KQ0OA/+NhoTR
Ruaoujj+7/p6/pd3DE6k9oL5ztKgKK4H5fdlazMs5s/zV1R5wkxk0NwVB3w2V3qPcKwSbIBjRCFU
FpdSNaZOfrGaVVQnuLlAJkAl2DrMNu6i7ozEQXmLFtBQtBIiBnJmP49NC9a+aGU5hlN19dFu13NJ
v/a534EZwSgK7s1T1/2rfY3/4hNn5qc7nektGRj/avRx6iw04M/SLLhIFNad3FpOWpXvVcc7QScu
hdQdrYk6HdKKkBRF7n/LFbDbk4lPKM39bun6q7vtJNiykh1KiggH2RNW+5R+pFIlJsZ0GDXwtf1V
so0+01w5O3RpUE1exkz/IdQGo+D/2im2ktVPuwulxGZXy0j4ZzKJJEhj7yNjI+JbI/eT3cLDo70Z
YWf3/bY1o2WPPpFD6HXEkVi41FAGbzLmbnjlOpGiSo5FDKA8PNc0PSFZT8oxZMOmh1v9RsuMd4Q9
EXmzWIXv/6LyJ7wFTCfdgmRDSbqJs86f71/Kne+L9+MNABfps2jHLIT5rEQ1lWpz7ssb9dxXj8up
LGxR99ycpQPnFh7iNktJ7zEK8VTXu58BG4+yk6GOz/+DmfrEYFYZKbPX1ekm817n+RzvHIawRFVo
Jc0jcGBFG1LS6ApVeMdnbUkX8ZBla6yAQ2Px5Ouf2vuCQaW1Y97scfQmGxMUp8wNspVTLW5Aylns
59Q5TUyoQmV8V1DfTlnrNmwL0Xij79gb/bc4COwq2GhFCsbXZ0vvc9Id32ydFTjFEl1zpqQkw7Kt
EiOkmUiLxO6E738RoOBhohfnwXGfsLdzOqKCK/jKInW6ypCYsIYUskAopySLiWBAj9RpLl2GXSu5
PJk2OyVVUx4QsWw+XiF3TqXeNz8bqfs+Yntps/9BmjoFTN9bQpaxA1b+E8Eh2N9pTX9eVrwzHUt8
vMDHc32F2U/cJ14fv6YA1zEBh44zLDJZh4MRREfVuge3LoUJiD+9wgyMRycdDBsXFYeU6FBS4NBm
efKyf7Z/HTEO9eqAgcWAQY1Vqzl6okArdvMKIigkBUv+ge7cbSm8CC1E3pXEXgERqF2fr0JoByPy
zNx5eldE/kQSCLAuykDyKTSKQuWCZI1ujl1oS8by4d1LjqeQmkwIAuSJMW34kCoZYvfP0B79fGaK
jIhtH0AepF0j7Zrj5X4g0tczegUveB5Ogp3Nt4m/vWukSDns4cEhrTlmw/Y+gzWZwasp5hpCxE+3
g6LTcCeR4vq6A4YhBR9zuvfaLEqxqVOlh7tIPVyZa4q5ZBVbVZRhNhs0D018wxqrwowPHxFWV4MR
NIjtGQ49urInynRaZ/S6bz+aKBjLj1UnuFM2jsQ6ZHszD5hozH4d3vvw7h+IeqPr3DRvJ+w0VjEy
T3ew7PR4YigdE4uXcu6OzmiUzqp2qCdl6umJyFetoK8jB0h+EJGHNoM0coksaKW8W6OfsiP6pRT5
Z0i8DneW+qjhnPk9
`pragma protect end_protected
