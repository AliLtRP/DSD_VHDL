// megafunction wizard: %Audio Extract v13.1%
// GENERATION: XML
// audio_extract_avalon_top.v

// Generated using ACDS version 13.0 156 at 2013.07.31.16:43:34

`timescale 1 ps / 1 ps
module audio_extract_avalon_top (
		input  wire        reg_clk,           //       register_clock.clk
		input  wire        reg_reset,         // register_clock_reset.reset
		input  wire        vid_clk,           //        conduit_video.export
		input  wire        reset,             //                     .export
		input  wire [1:0]  vid_std,           //                     .export
		input  wire        vid_datavalid,     //                     .export
		input  wire [19:0] vid_data,          //                     .export
		input  wire        vid_locked,        //                     .export
		input  wire        fix_clk,           // conduit_audio_clocks.export
		output wire        aud_clk_out,       //                     .export
		output wire        aud_clk48_out,     //                     .export
		input  wire        aud_clk,           //       aud_dout_clock.clk
		input  wire        aud_ready,         //             aud_dout.ready
		output wire        aud_valid,         //                     .valid
		output wire        aud_sop,           //                     .startofpacket
		output wire        aud_eop,           //                     .endofpacket
		output wire [7:0]  aud_channel,       //                     .channel
		output wire [23:0] aud_data,          //                     .data
		input  wire [5:0]  reg_base_addr,     // avalon_slave_control.address
		input  wire [5:0]  reg_burstcount,    //                     .burstcount
		output wire        reg_waitrequest,   //                     .waitrequest
		input  wire        reg_write,         //                     .write
		input  wire [7:0]  reg_writedata,     //                     .writedata
		input  wire        reg_read,          //                     .read
		output wire        reg_readdatavalid, //                     .readdatavalid
		output wire [7:0]  reg_readdata       //                     .readdata
	);

	audio_extract #(
		.G_AUDEXT_INCLUDE_SD_EDP    (1),
		.G_AUDEXT_INCLUDE_CSRAM     (1),
		.G_AUDEXT_INCLUDE_ERROR     (1),
		.G_AUDEXT_INCLUDE_STATUS    (1),
		.G_AUDEXT_INCLUDE_CLOCK     (1),
		.G_AUDEXT_INCLUDE_AVALON_ST (1),
		.G_AUDEXT_INCLUDE_CTRL_REG  (1)
	) audio_extract_avalon_top_inst (
		.reg_clk           (reg_clk),           //       register_clock.clk
		.reg_reset         (reg_reset),         // register_clock_reset.reset
		.vid_clk           (vid_clk),           //        conduit_video.export
		.reset             (reset),             //                     .export
		.vid_std           (vid_std),           //                     .export
		.vid_datavalid     (vid_datavalid),     //                     .export
		.vid_data          (vid_data),          //                     .export
		.vid_locked        (vid_locked),        //                     .export
		.fix_clk           (fix_clk),           // conduit_audio_clocks.export
		.aud_clk_out       (aud_clk_out),       //                     .export
		.aud_clk48_out     (aud_clk48_out),     //                     .export
		.aud_clk           (aud_clk),           //       aud_dout_clock.clk
		.aud_ready         (aud_ready),         //             aud_dout.ready
		.aud_valid         (aud_valid),         //                     .valid
		.aud_sop           (aud_sop),           //                     .startofpacket
		.aud_eop           (aud_eop),           //                     .endofpacket
		.aud_channel       (aud_channel),       //                     .channel
		.aud_data          (aud_data),          //                     .data
		.reg_base_addr     (reg_base_addr),     // avalon_slave_control.address
		.reg_burstcount    (reg_burstcount),    //                     .burstcount
		.reg_waitrequest   (reg_waitrequest),   //                     .waitrequest
		.reg_write         (reg_write),         //                     .write
		.reg_writedata     (reg_writedata),     //                     .writedata
		.reg_read          (reg_read),          //                     .read
		.reg_readdatavalid (reg_readdatavalid), //                     .readdatavalid
		.reg_readdata      (reg_readdata)       //                     .readdata
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2013 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="audio_extract" version="13.1" >
// Retrieval info: 	<generic name="FAMILY" value="Stratix" />
// Retrieval info: 	<generic name="G_AUDEXT_INCLUDE_SD_EDP" value="1" />
// Retrieval info: 	<generic name="G_AUDEXT_INCLUDE_CSRAM" value="1" />
// Retrieval info: 	<generic name="G_AUDEXT_INCLUDE_ERROR" value="1" />
// Retrieval info: 	<generic name="G_AUDEXT_INCLUDE_STATUS" value="1" />
// Retrieval info: 	<generic name="G_AUDEXT_INCLUDE_CLOCK" value="1" />
// Retrieval info: 	<generic name="G_AUDEXT_INCLUDE_AVALON_ST" value="1" />
// Retrieval info: 	<generic name="G_AUDEXT_INCLUDE_CTRL_REG" value="1" />
// Retrieval info: 	<generic name="AUTO_REGISTER_CLOCK_CLOCK_RATE" value="-1" />
// Retrieval info: </instance>
// IPFS_FILES : audio_extract_avalon_top.vo
// RELATED_FILES: audio_extract_avalon_top.v, audio_extract_clock.v, audio_extract_vid_clock.v, audio_extract_core.v, audio_extract_registers.v, altera_audext_reset_synchronizer.v, audio_extract.v, cai_avalon.v
