// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pntWVi1E+ARUEPySZ8XRkyUhSNYRe0N5kij2HPVXDfnG+KCeYDO84Rb9ampmbpYx
Y4TOY1gIrM76Kz9F9+p0n/b9RSYkJSDJhvAbguBaoXEP/XSP/oVKS900ZSw/7DA+
GvNMqa7xSBCIUr2t+6ArRhuCaFSHqNnnPwLcV1UPRpM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 72560)
21sBR/rV0EceSXsqrBLqBKxQ4cYEBPIRq0evwXg29uM9PuI19hYnLGHAjLc7EpP2
scW2quztiA43gEA50i+eIxfoOCZiap81PmVUt+FBwpuw0EtMad7xzd0vd2uIIoM0
aYVBrX1SOrReA+X5tvNy1GdL4i775JEMboOHXZLZrNd6XdugohSCwmBbmailUJBk
nwcYNW4kmO/A9SkulJ39YGb/m+o0bDyibXFdiG7G5f73MVQbXBns2cGNJTrH9WXa
WqbDW7Ua/EdconMcZBS/aSyfoVVnTtgBDUjzE67XhmNkW1OeNeBiSGhtwN9I8FBL
W0KOqkcP3Cd4kaYpw48G+kx4sAmsHjSPE2+4ddCW7ylCKIz6GQ1rlzqYKtAglE70
ncDigLBaY5n60x2Tnh3FH8B+8l/ps/eZCJC+PzPRIKpw5BNM3Z227u5aaII3i7SC
Ka6zV1a9ZzzL8ont0Mna4EbGkxqqICMpDCEXj7td+M0B8nOQc1J9mBKZOdQ2g+t+
uWFxSVQPNY4fcf48AxW4ou7qgbMkN6v5KI/IGsS5Xw9gs+PmpDrjI2GwYWDpSG7d
uFpLCRV/d42nhqkX7eQTvV7lPh7w41/cJX+joeGqUbbqQId5EAO5tZm67cwKOGKE
KEihBqrMMwmVcFaaHF8doZX0INZM51u6Jw2bJuXJLoQZmQGJVGKhLE1ml7qrw+qJ
lgv0OsVdJ99JZkpPkAMT3eWwG+oO0U+KIK/nZgNGeRYz76fENRddysvHiiGcSwB5
Xrl+2uxemGimTk6H0RUHFclGCat/KTwZXyNBOG6ztZn/PWF083GUANaWfgX+awVg
HBRYYXaPT3LttR/CyNdP7vIWXYFl+C0jFqgQY0s05w9nrJ3oUSqyptBcR2Ik66ah
st03HTQfKfE7S7PvD42PIupJDeoCJzEOqU1YqtZGllIrlS2GaGGp3A6YMTDXRnNh
qNHXpfK3YBrC3TEjU5FXiFhWQVXORphi345s+mdGkkacd1Emu77ZVNd7kHITB96P
bL4UQPMMjwfcjBMuM3joMsNYAS6r9JwbfAsgIoLDJTIP06Amsm9+ynRwIWwiTLq1
X7O9uyT6u5CSmIh6HAgwg13KzCI3g+wyGplg11ZndlLlvFHt1YIPxn7+ownebVmC
5Njs8azct68VmjVSBG+lMvnoeEVc6EEuCRQ43ycwcOskLYmB5nKd71IB3z//fXAR
cmIpWn9JZ3t9FaMYjMvbrPDQTYvO9MRkGOqZT4/TIHg9MRkKxRm0K3t1j82Woj9e
tY9x9+jlt4MXwofexng0rJjxIugZt7ZNIJ+x7gQhwHiLMm6kkQPTxlgcBrylQJaL
sMCDBgb9aVuvPvMsAkc+xeX3vXWXFGnH44N/KeZC65GS53fxEDMzw3yqdZdvdctv
eEvQg3q9D83n8+8p1NbsQwfoMM9DOYt6rRdJXFnfEYdmJiTOg8BS81RxbjVtemjM
TK6zvlOmmVepSrLHTetIGZiwgc3y/VCCIKMi9EgFDujmwQFfWDwnInKveXd5Q9HF
j4dFFdZrEQmIaojNUb6vZNWBhn5fQMjGzcUE5Cz4tbeJv/p+gwcqj9BIoKQ92OoX
7uAaLcQqLxMnaNYdKEaeXkvfIZGrB/3ot27b4rdgoE9QMBK9xCs/VSlxu2hbix3Y
+aWeZuhMR4IQDHxwvbguhaz4OigZt900yyVP6c/sFs2dBx7BFvrDB6MK02uoVkJC
rOcdVD8xhJOn14oRi5O0NDZflQLCVS6GDTHFuUg0KfoLZfbB5rfXZ+348z0zIGaQ
gmVBpZsa6FanPS41T9ym19ikuEk7qm4KaqF7Oahv05avOPiztSsAr+v4oy4IdIg1
W6jRTMaEDozvOVstYrZF71WngLfSQldRoRMAezhXazXVk4bEETEkJq60GqNKPDWv
S1OXQhEnzoKaq+D9eGEzNZUGa4OItFcAlgecjzjiCkP2wNXsGRIuZI4t1zlncols
KsAG1w7WIDpSR8yUQhMBkmxM6tjYvvLyY4ezSxEbEw3FnXFYaSA+aON9oYdOj82M
NBL5xpgp6BGNOsdHf4dBRGPIP5oTft2lv3UWaOHPU98QCEGyI8aBmA/m63S6HNdq
BdAYvBJ1HddKuUKC5xoDysrFW4nJ0LEWXBXxxtCNQ6PkqN4DIUJJBPQA4ABQDPAn
S5hHrVD4KI0LiDO43UeeA0ydfUM3+9EVCmI9LdzBwLKejzVaurHCcbh2kULkoRMX
vXa6TyAVUmO4hAFU4SKZlMWDkTDWGsy5ctj8lRW35F+H15WZyHvb79LZ/h4Pzr5j
/mfyBdVFZQcpf96oW5ZSclPmTVtwhMecbj3WQatCdRkcxr/ziCympPxkLhgfUHbc
UNmOmPe07mirg5eNGkbH61pSm2aBDpne8JFZSboAnXPUA9kFK810lsvuiz/urWP9
xTLv9BvRUw+Dhj4rnw2SrrHJiOIIMuKVz7MctuPh1PZC9srAFPYJ9h5/a3pD3LLy
sP9AzwdOzinE+AFrz3PJQ/A4Kz3aOJTXAPjf62fjD3nW8Uo3G9jEqdk1D8/3By3K
HAdqE+HRRmTIfIAHVrM8XerpHM+UlAnUNbGK8Db6feAv7yQmaTLK8p5wp2OSdFU1
JLJy/aPz6bIttNhhGnn19/KXBlknq8Z9/QMeqFKmH0+F4YP9VdrVABEDu/5TuX9n
LCsmfODMGKWWIh3OULdiD1fQt2dJOuYn5jWrIMTWPhD0IaDAuSBNfbZk7EYyuX5b
+cYSeIveRiZjOxDkun1967yHxr7X6Ukuxndu3dm5eZa4kHoFeALhVFRn1xWV+YZ4
bm4NSBdbPxVw9KOZ92TXxjd+IwnmY+XuhIvh2W9e5EWUVzv921oWr8y7p7uccAoy
21GwJFV91KAFuDXPi7PwjuOfK71wZ5agKdIRTp3jk7n8Qwx3gCsF3R7UsuX+PlvX
EqpXpDpi4yECp7eDOG05V8d693LTa0ng0L10oOcJ7iEZ8HLpP/xsNgLmpAdWTIDx
oWIZy7tFHRWHAJXpOzXlwK3KVmp/dDOC9seLa3iGK1t4UvySmcjtYvVe6Cgy0Gbs
mzaOBAoNHzJq6uUvGPiomXLaVhFJKoPQ7L20ki3BRXSQucmiRwVju6zLgrv25iuv
eZ0vpgScZ92zybtGmkJrmy9uosiKlFJgy2GGdaRy5+1ErCdUQnKU63pCuPKw85gD
k0HRRi2WSxuvisvVlt4OjWsOqdjaiTqeL+j4ZabG64FWUJ9rFH6B8QgPmb537KT1
DN+SDxnmX+GnD3B0Q/ifGxntfyzvYRLSCYpbeiB6UGRTe5mw2owxkq86ofauJ6o9
THTYfMYXzL/jVR+AnO014YgjK9ZzWsJm8zvR/Ovx+auMVnQZQVpHAl3Dh6ysQpms
NdblIWHp/SXgRX+gVxhpfrw9tlEhoQtLBy6sRkjfNCSo6I3Xb/EGheQ/I7QkTSrG
UeR17eEDEumvsgsok1+Ggh9qv4PkA5UUcDr9GjymVCEvMAZsQM4V65WDTeHMaOXe
Quraey80APhL0v0t6kogeV0u5M7UJ4urhjc9c7b4qr7+FIda0x5dUjb0/Y5QZw5y
0ne+X/uk5jFM/WaBT8q/56hSS61cYhSR1OV9Y1dRtMY9ZDejvpC+sADyH9/jTJzD
DczYeYlo606g70c9VYUfZlOuVjHopzUwHD+g6NXIx4C5ZUv6qLdKvXAs8jJ1ocM6
h1P1ycifWrXHfzOK3+N1jOexfPxp6y41v1652lO6WS3Oh5E+gmeFIz6nbWXVaGy5
zy3DqMlH+Z8XndozGVk9niyJoDEd1/7SVQ5PCECiLnhpT3cjIEJX7aQl8X79E/CQ
fhJC0lulP0gsFgCh1S9KoeqfcQMXBGPEaIQZ75ejfG1DYZT0kezve5O8RnMOHuMl
IKXj6YEiKRY1kpmtC6WJkhrRuw7rsdn2lju9C2AFnItc1Tt994kVVxGzgnFODHqG
VhoEWk3eMlk0Xf3pLHG6J1bqkuvesFJQ8Jlyg2MKazoyv+TyMGg4ekf/UeTQSFLm
0ScrrH5++IaDJyKJjAGw7zaX+7289AHay7yS1QAGzqvmZQOjEovR+zAHVIz15O2g
+kAxFJjvkIxEO4ltsRch2clG1CryVSl2sGEVykyTyLv7S8mFM7wdulM+2Jk+PFLU
AYvbDZSKELO3uxokL+dHm9Lpa/BbKmNQ5SnHgidGeHhSOUw17c8KtfdELtt9s08X
VqYZr4/87IIep6TuxUwdXXqz4v1M4rh0RGXa830ouzKgHF4ppOlT+L0Ze2nIpONl
T2TTuZ5NryO+f2Zfv6z6EPY/789yQjOf0WVrdWjH6IJpiLkeDteR9sdfQzZAWDdA
olcdPaff2Jzl0ydnvHBMiQxbrwy9zo5NzNyU+L2JoVy6kWec/oefl5rWSwp0PQa/
3HBE5aiLzF+WwKprzUU98stFTXr7hHB+UDTE/ALGCuWBqhoDB2LQgsQ9myhgF1Gx
fxseevy5yZRL7ShgEFsnRR7Eycv93r/H5b2zhaSwfR4WrGLN/qVR36TJe9hKE3Mc
5puv0gbUtCqkc+X1IrWeyvE010+XNvoWvMD4fBZYi/1hj2rb3Si86P6GUxePOUn7
9z9lrhQlHF3QSStaYH5g52T9hqrKSUCmzohCzbnjlA1o6K2O8waj4TzWwYRk0lZp
EjBNpK96ktyMWzpzF4tiIRWWncOSrUikBuyiICAPk4WBnQ45SG6RRho7mNFUWD7c
EcpyBdkdt/u3U6dofDlYIPc2D3wtMoUj2EWjeKbLWmXNFquTly9y0eBZH9A3s9uQ
IzilpRy6Xu+hJdxoJ+BgS9MVmJK8ihDRRd9j5yPnIonxxGgofpgf4TEs71k9o7dj
FAA63D1D3lLxJYzKbNiybu5Vzc9TBY+pkXWKUFn6r+vdiiTYNmQMlmF0rwva5KWX
eTtaVFS7Osvy8JAAJwcNYjm0M8C0U+LqbC4R+LwRqI7CBc8XDVrdFwZWT7DnhZDh
ITx159UB2e1J0s5p8jx2tgCveXmtA/KuhWiw9HdqNIUA8uCi5w0JqcU4TybSY3u8
F38cOn9bYFyDG1YTmtUxFoYiu5+KDVyI3Yux6gjfzScjrPbwFsZanJaw08Wb4U53
bzFVgztQ4TSm9kzxYlEhPnxBNCWfX/Z0ltf14kPWNzuVJwRjOBA2pkzBcd8ejL8I
PVQAEi9P/Z4ijOTrfevRCF8AWCVJ1brEuL2Mab04/pMq5OeD98fvYBZ4PtLOMzaD
kg3yXC6sw+0NL4T4AKWLArDNVWAPofOgGpi2DtkzZPkjyj16/KbPGpkGrEtDoAZe
LmrnOpsnv4RVoaWAApTC2kefuAKXou8wkcA2z10BUHR/BCWG4c/J0j+OVMdMkHzy
Cw2xUBwoW4CB4aaij070LnyiEIKnW2vNi7edYlqNGKakekCXkFEYmOHp1g2Ey6LB
GpJplmrA8Pfu+PgbgU+Es+sNlcy7cxaarZ3gAJ3gtpQSe93dqPKcRqzQQBfrpO2f
aJsVnCCpRnQ4n05v5/edzwlU3vyO50Fu65upjQkhJ//M/blq1no14QYUI9afM73x
iPm5XiSpPdU3OcE+4ZbHulD/fnTB830iJzMkkob+KjTq9RazXwl6wHup4LlU2Kek
eaGjkzgKVEIv4vkJDnC7DAPHCEmdmI406wIRwPIVQ2xaYCS65JtdVyP8NI7nT462
TInjWyOmEm1JMTS9grSpJJSTOnctSJzXBrovAsnb9VPevDkpOYEEC11mxBJAnPOU
LrVzxUxCV0Q0MWaO19CwzQVo/BnWX8FZcADHF4t2QAZ2cATs32sVx91zky1CSqNO
/DWgvenjWzFV3nsnaZMHroAzhhsHT7Q5+n9S3i3uo1quPygG3fZSE2E2szhyay0L
O0Y3yv6VHrdIyRt+72+86DWNR753nbyUWgBKtxUB7hSDRjz7iWtdi+7aR0dDomdb
4wwykxUjURlXz5QZl+MJtGix3bBCZgc86nUspkIP6gcwlhZcRWwuvAcyqv6urKag
5eETvF43qrWhSsv/j3njVfUYBtVLGv1PMGr2SnqPdx/JvLBODDgxjzgRsrp9kUJQ
us3SZ2JF4fzhuusaYtF68UYv1oomhFnKItwmZSuR/lPa7qBCMscv7FwfSLH1MGBi
5g/AX/ieSp+sED8n/BvmX+RNIEo4PYxv/1m8d1yuV/FocumeYsZabmF5GwxwoG6f
TuN5x/qFI4N2D/AYj1QULIH+lXVr5lx8NI9EkZ37jPsPS9A2BqrHl06YmiezOc5M
cqQ3rZ27x5Zo5vnxyWAiiY13wv0sBhKbzfwD1JiXNGd0NK06sDDQ6jByZlCSQkwo
2Nmg8DHm8xlkIJcnIWIgtkD4UKis6TW6Yviwj9/9iegzCkAt3vmeVgQP8JxPnWNX
CazvtbotFg+xvOeqObnQtXT4lU60F+DShcgw7f4OUcSnvxYpWTUUssUj3FMr+n/r
dtwAIfdO2xTOC24rgogbaUWKM5TBm/DdUVKbEKbNbB9MeWgYfmK8cSrDDM/34Bgo
2tQIpy4ECM4CUrBCwXQe2MUF16Jo2cUFmX+e/lcUT+PDQ8uTgj8SwldphFyUuw+s
z15r+tptrArz8HSi3hcLCPbiGJM9smydntb4wzEf5FDd1XMofOyaRTk5WFVi9x/C
3jz+ULZhIY8mnbssuYw9gJtEk/FS4+pPNKDgL/1QRfDtdTSMldinYwDqqzmgfwhs
8BvesQqA/tDDxZLRF8S5U87k3FhpfXfRhUuM07ETsfLluvcVlxPMxaM2Ppp0rEbn
EoerHdcuWxjKq6Fbkw2XI8ijWR0vWV+d6seMLcVcjixGuYpn2SifWsK9grBcWDAv
k9daK+YiRXPWZcyt6LlZG2Io4SpECBi1TKnQw4vfDZ+EEi9GYvfkftO6+zbQuuMh
pdJkOx1LjpfE/J7LIrF8+Dxn/1rJXpCDVcTJg57W99o8nEezL/tVIomgip90yWlq
aOzwL/5yt910EPpCEqeVnGRVF7ZftNX/tbAmTBwOJn0qlkKoN6kYxN6Xe8uwkISk
WOVtKBhNPiCpHv9yGiEEVyG4fbjlq3zXuQNNjsH8zBpBJ4glp7Om+OOv2NwfaETh
qJDEcUf2lXGHebx1O8UvGXodi1Rg5EtgUfFM/JOc7DeUjpqlXyh43TqBHETkNMLB
vLULvlS0nTP5y5ytsnFwPsFpKINmEGUX1oFFd9yr8z0KvjPGiyWlf6ymBD177PY/
q/4ctTONl5qwVzYBrmif+8fkAiFbqUi+xlwGzADBD9NfOevUY6bxLd/TqD1XNBix
37gy9CniEjLtD2u7iURykOqs/F9uI6CINj8/1m0ba680br/LRbDjvUdcX2N4KgAD
ePHSf1woUm1O1AGGjFVNZgeZEL6AzX06JF+GkTT1cwNR5wYx8hvs2R0dFOXaP7ub
p/wRY8pPl3/QkCvd+vV1BZCs3Dqsol8J3ycEOcwk9UgtUlmz/77jC00rchyv1bQY
EgSAKbI1sImSIWZtMNBGIGNaL1r7JTRjbHZm4DNJK+2DnZI9nD9sY5zuLkkMYqSH
b7Tg5aKWvVjWx72oxle+R3McdqSsEvqBMuwLmIO91/pKtVgczgZKH743GyolKCFw
pC1ltd83pIOeUd+HjqPgwCI5C58sNRHdM2lRPZfs0dO4IDJnqJ3Ka7n3M2BL2Rsq
TAeGDgXXRrZvivsQE3hrVdsn3z2uS6+fW/dJYSHtYzo+d3tRgCnj+pVQRiX+95Gb
H6wAENKROzrb3ADUm6pOQNdGcsRiTJB08Rd15Yt4ALNAkQGZpDg8xwGOP9ZLpN0I
TJ68VAhrRTVEcf4PDMIn+wAJ4AuVasqS/JQLms9N1ZjUe2z7O/Td2ZeOmLE1NEVa
HUpDGJSlhTvmJO8cJW2RVpFUf6A7b2eFVWFoNqGAw8vwJLODlTgC8vn6btqhqsAC
WOYjKffvb+u3HFm1VEOP5eZuaWDebyZ8oRIO3H+BEJj9aSYaxxt1266/bQkyl3i5
voN94RuIE2VCaGQId5m9a92RQMy755oC57l5QWFASDMFVVCSOtLlhRHzNjgdwb73
iRrwIDL0vGhTmDzbX883QXaIYWOho68tiJk2i5inU1SnypuRHxj5zEqlfb5IroKG
Kpwp1Q6dVwtjELbeY+sFJ/xvGVrZsZkJfqzwUe7g6kOACPj8r+6xi8btjXyqmvgM
1K5dyU4yyiAI5kf+ocZ8Ec5DLQlkf/tBrWm2s6vjTock7PHt2jFp/h3+7juCwJTF
DyGK8cXA60eXXitB+unNh0NZjnyuPzfbTPY3Oto0WfVosCM8EEhqQogJfYWahtMM
T443IXoWyFHNPBABfjYD1jGHgjCXRFTH41rszPZJk7xKU7M62bH9zzz7gIbWqViM
erR2xiGv6DQWo3cmzVE8r4gXtwo02RkJCWpZnqeQkF+p+xH7ce4ISC8RzVjSB0mx
x9Okv9YboPMTVU+vIbQbZU/+VlXxcC6sEl7ij86avWpdX2gJ5Oz/deKUIOtjWtDo
hzdNlBmc09JgKvDmCzN1w7yyTZYKBiojn73iyuHhNGx6drfv9vZA04QtxDfxP47K
aBK9fh2T7EBws6a4ZOi/rbvpYBVCK3aCksX1pdyQDgSvAdF3Z/ZbwQy3ZVb7etCb
KyVzkIzP/PWEbacCU9X70xgWYuGdw8nd/YXljC0UQcmqD/NVFyJUwJfA99obV7oX
L5rS9IMtRDeqjPZqsZkKZczjxJxlaZgg5RdAeqE0mu9ejf1dRPMJfM6ad7Zx/huY
F9n4xDlwW8r6JmJ5abWcV8nlQrG2bfyqp+M6e8Uu4KK1hmbWQYUdOpF2r5w7hxVg
IluIDnsx7Ix+ndAt4YpFRraDMPHN0xkRp8loIlD7nw6ekFTAkVxrkXUTEaskT0kw
nsZRxfT87vhYeJGGXBzUYZzoXYTu6WagauCbi6khHv+j9zxoiMY9DU54qzondJwQ
RtfQbb9pZ9TI+sg1CjNO3WRMfc7BrYwEl0wPdQq7eIM+4kvX2dJUDYFs0PZ/yeYt
9v0ATg9eU6jiAYntXHkvGz/lcfxvu+W/3uskSGO1jgwrGtN4gHFWDd1W27eR8VT6
N2TWpkxlYkX5asdl3aiIVCbUYYs9aHS1QZzMxwFcrPxPOdMnFmfWPlmZQUQ7170o
1jBxOf/mK32r7muHSjkZhbyfdImGDOB3YtovhXIwbkO+X9Fv4QMlYuhKD38xT345
A1+1zS/CCmPqMrb5b9otG0YJB+ktluJujFSvxerYe6sQoLN+uqH9veeGtxgy9YE7
b5uJmV2MAzE2tw7zCS4JO9Ci5tECGcW6ymdfVEVk34+e2dq1Z0/wncYr8IOg1POt
3nopZM639pSPQDVTCRl17sXCqgyDwkEvKmqBI9YhgJ4hjlywzHaaNWoz03lZ9YKX
Nn/qaUC7z9kmwvN3JQDf6rMfJ7Ns+2K6ddFGy3qshF4Hvn8Fcv9t4IGdbC2Q5FJR
cMIZgqv3fs53/Uc3CW99cy1bhas/Dq+wiUv0wy+/tet75f6HLykGrEWaaJSn1Zq8
YpwejX5gzmLpyAcyEpLoI+zf1SofIcEiBrW7aLUknLFA2TzSbqmKSBoqJvqy5MfK
gS56wuKik/vp9m2MRDPDF2aEzir1Nv2g1sZTgJqW92zMzBDmqhcLHLTUwdgUk43e
MHQDsPLcfeDcxphdpH3YzaQjVPIVOLoiV+coD0QNP0VP6R6zqN0/A/XAjaU1/R2F
gimuLg0YMQZOxrb1cP3hL9Dlx0Ng1jbtQhSpKXtUZmBOFMyxqwQt7u761Gq1M8GL
4+VlhEgFz3fVOri5L7APWWsqF4mtan3Z5N5F9rnu+qzaGN4HP2fBcWDaIYdHnjRo
LbjvLohV8AMekYcrz25WzqfEFCc4tix00jpBmrWiVEjt0emcTAukfB580Xh6JExB
cPEbcX3M+Hx+T8b5mV3AdqhSH4NbUkAf0fhlpAYl1YQPVtv/fjYpTFO34NE19GHp
WExGjR9PqzwONxPZDFI6CGVWrgASyaq63PwyTTNziQF3Z+IY3SKcEKaDIpBbrv0Q
VxVxt4MmThZKEJ/3zxjGSc7OxEWI5DHR9XXT8dET3c5bXS+iLs4FHKTsZBB5l4kr
3GFv70cZztr70LSi//Sf0/BZtWP00uiG9eMvDoP6R9IqLfNMYM4YYH1lewWA8bIn
pprWs32nzqgD3aG8GX3ktF/1Vv1jTFgwQ8b+PGpjuq9UVklsN+2TFmupgZY6eF7X
u9YZAR/UvTXH/cLHnZ4GpqQBSxpNTbzQNvQA9vIDmhI+SvBNJpB2gZ9ZwDJVy7t3
OU65d2/In/RGhbOR6GqxNOfc5r120BSEPC4//nyxJ1fsmcrPYGQivvVkhEYYNyr/
3dDDxnOAlUn9SR8Ga8l4CR6SRUMbEoK+7LfN4Y/l2IimG0NWSPLNOlS5G6Jg7V+K
6E0RFrBfpGSQASUp6pp2HHI6V1jtauQ4L8mP3YV4zHHGv2vsm28LAVzW2tHDmyuC
Tb9cgWWsUlHMEZRIQ7SLkUefzZIFZrZeiAQJSN1xL+YRuQE4QP4Es3iJScG/dAs+
ptR34ROUEqanYvVai5D1FxRYHBuWUq5LAsrzhJP2W2va8Iv/+4821ED/1V794qe9
VkdzHm0NJGSKqpbOnqfxl31QJdlFNauvZfjsJppeh/+o2If4ToNMtHqLavJ5zZNZ
3UBYU6Xdr6pdpD2CLkRNX6Bnk73Iq0IlqbYaDVkVYJhHFrGDfhGGwLP1P1bApUhs
qTi9PjAVQz0YS/0flGYBgIuokPrnz9RZ3gx116EMYM+umIBfJyJ+25mwLu5jDNXn
2fhbuapaZhdgkfSy3JQ0/UHhxTtkhOsqeVZ/7XFWeeFOP7hhWLne5xmgN1ZXeWil
fHqCDkKdyKLUPjXsfIk5iIapghY2XUiHqclIcf+aKFrLmFWqCo4TKba51K4Ej0pb
3/xM9N7ItxcpHdTxykWbk3cCQ17W5ZCLQYmw6/QdZAnu7saDp6NViP/jaBX7Omvg
VbY2mntdTXch/yt3ypxKyyZosrp5z4PTVtUMsoxHD9JEYc+GWcq0gkJOz+OWjCSc
t0Z7+AVqBP4ftHCa82xzyqwcsLXspyi5W3rka11BWGfU+niYVmauYyBSoP5iXSqC
vok/94qmYtuXr63D5MLEv2MXXkSnCkw+5mk69ywSqVbXDIQiwzQ7P/yya83eSM21
REl9SgwY6BFp47oVgzMf2bLo982UUmuva7JGmvxSb1Pu+UeLrQETgb/8cxstDCR9
xmokkoHSz1sQCZ8XMzafKFaqIEcUeRKazt9DC163EQzpr0/8P4svyMog0TLGD70S
iq6NgN77z5mnTzqHFVl7c5velMZcs94SxPllArtrgRiIVRQq1j+3KjR2VYi8765Y
yONYWJjGnzh6Chj5yxiLrMqhF6XnymAaS91aNLs5MGDWiMB7D5djLINNGRURHq4M
yM+sQL4rKBQFFh1I1Iva7CVj9PhepE4FCjDu3VnxXcGOqtizyygmvDHSH++b4Wpq
ijZmX1LJSGgR5sItWW9goVHsTgNlBzh9c1FiHtbXGQsJWpvLl4h4/4xZJU4cKOUw
tY/X+/IbVrauR44RTbwEkSL/TlpstJmWv3wXeqfl3ghR0whIXAIGud+00jM5p11H
89DD1aGhI4XQleC166L0NhFsiLfC6EeiP45He9l2kt/pu1PiLb7PpPnBYX+uSnsS
beXcDoOzCUnm++jtKy1ca0DnPOu5GguIoSLluxL6V8idEGGxxOX2d0iYDPFj23sv
Sc2kGfIKA+AvqcXPBCKPXq0s1gX2H7Z/9bvHMPx1NYZCfu3vDRkLQioGFpzrqYh/
+Z3raYppdsb8jgpO7JuiYU2wzQTe8l7Lhz/YC7F0b6ifibe4H8we0fQXYZYD9LeD
bvkO/Vvv7R9u02Leq5BpsfWAAe2UB0g0hbc34xnsam8xqm4Tw4zvKzHMQabByE9K
Y11z0QeGjbbuHcEp28tXZtEdNW+HPII73Vb3lhkIAd4tbSlYsd5V3fzTGlAV4JX3
TZHt+P3tCdHtNYSDdTGx9sJrHDbktGOgqDKx+SWA3Huf+g5PTMn5DAWh8RA1ful6
8xN4mClk3dGeL/wELlVB1P2KUIBLggFYEnTtybA/1l2r8f8aedv6p/8bOYqVbTof
HAcp8z9LgWv/jWKYuS3OIR+Vr3WJ8RtAfToPpR0ytEA0nI865j4D+2qasQCdG7WA
29P7qpDBon9YJfm2yAuzISHeJUpZmH2fAGwRte1QBytg7OSf9MCxlWjS/O2FKeIX
KK7YRnHh/bqYZPPoC5CjYFiu1h02Km0PdJpnLy403QKtdUmufF2M943T/UhhpHnG
l5K4XApdN2OT8dP0VmBuPvds7Z8HkWTwJuAG2yBMsqp746R3VrM/WW1cdBYfsQGF
R93Vc5gxVNJWO0y1O/1gBtlwZPzkmY52L9Wp+VUYPOdt+QBbTe6LqlT8Ip+pJpMq
x8XNVZJgV3Lc0hhuBd9esfHfxKEUDCXOvhFmFHcnG2ggtXaEQzXwakxYbKRv99Rb
Cr5l6JfSsV+fhUz3dLcajLZNO32VZSgwFfdp3/42DK5zg8KUN6Jxa6Wo6ayAlcKk
GCwYQpfqw1FbA9gKzBay7NjIhtO5pV2mndK/2D8leU1jAQ2ioTa7bS5dBrqHw1Iw
3Y+GzG9a3CS7HDY5ffe87yEVcduUN1gIV13ePH7nAwzD7FsalaVl0fHyBT+a756s
1LdQkl3ZlC2tdh/k6HB7zuOVQ14Y06lyKJudytuaDAEtzFQ5gSn6QEVL2SHznTCD
tFfxvWNCw98PrABWxGkZZplyetLN+CoMq57BgsBx8nG+8YzHQngPVS1S3Kgn+CiC
CEK8jLaVB4B2QePnghRgnbttusbYD2aPkwJJgUpNPl8Uman2V6cv2nJ8mSQg1n05
EoiRc6BBMzGOsJna3duqvnp6qieByU0vv9atN3l/ftUlTQZGoXMOvdnfo+JsEXfO
sTIsNy0m1sOlJi6/UoGtg+Xyn4WV+zs8mw6Mc9sEb76OhFVpbVAD7e/dtaNxJzyl
uzjBuWOOkIzPlAEMF+4ZuXhsgJdVuBJRK1rmQ+K0rlfqrY6Iub2MrS3mUFxA/ElA
JLuhE7ygrf+9GdYwaBUqiQJHfwZT94BqqqLk02NqOOpGaOrQA5yQFYplP7ozCBjN
VMpJjWVHMGGOpUrlXBVGzr945Bc+/VMqs6vw5b+Da7bcqXi8ocTh7DTvUsUw7yCi
E+FIu6GdQev/9ce69xctRJJM5OPHJAQ/W9hBiG+XmqDWbmzMwlEDZch8+N5LcFln
B4f/hCq7tveCjr7/24i8iw3LfOdx4GI2vswN0xw3cJ/1PjfxTrPR7ytS2PydLJaZ
hUZSJLtjbUYqDM6gXEt/qKugmKX2x48P8S8DeGTBZo8WVd9cVo6WOVwkiLhjx6XI
CO5gsclC6UWaIzYQLVnLve6lpucdHvzl7blSp0zRf8liKCOG3GdEQBeLkwTa732M
nOO2nGEs4bITVEm5YhFDkRmG//KAnSO8xZKiqszzx9X+z281G5CfOnmpz+HT4/hV
vFZOJXGOwLZ4q9pVKIPdWE4QYIoLmIdUCu7RVeoDpeTMgWs6yax+/kC217QYUeaR
/PnEnQwkG8RqUMeN5IeUXHstgCXzpwuxkq9NzBfWRRx7eeuW0m8UyhQK+qSltBJq
RRy31RZJ9K0Eit+z0uRSOMyE0G0FChamxO3y8aw+7I0wNIX2vJbwwFSeyk3Hj6Em
AT55CyJkeyGLN8PcL0YnaPhlaLuMsT970lOgNhEIu48S2zefZLKodMq3In+ZBXEe
bQM9DR8hLT1QGWU7Fs0XPrGkGXQSZU6z98Wk60t5uJ3D5sOpzZfpuCpN8c2HuT/Z
tSn1IwfZ1qqvY6g3xP7tgdJj4HtbANLx+grjpapn6f1U2TG2zEhiSB6wxWrfLKcZ
HPt+d8qwgV2BqS9EdIZoY9OZPUJIfEW66z8PrnslV7BdLcJF64vctkc2HKb2EqzO
ndjPGRfAp7TUBholV8bty2SqEdXy4nXYcw5VzMbVW9sxmIA/eOrsyc5LD/nPNtNG
XPVs69dfizhnHRJVXmgLWfH2xjENEnBqbAp39kUha9OTvfKxLnAXyJIrpte1CsEw
MBjHHRv2DaZ1RHdKhb4YraccK6+PvQo/DOhZTlW6qGYuDfxPxjS0CImPYy+ytTkB
FgD7hTy8kqEYLUPW2qM+RmhEcEqMDO0Gx/65K08vozI3LoJb/L/K3XQU8/A6n7im
SAnL4RTUF7MgNKTlk4E8r6Y2D7oLfiIB0Fc9gVwERaXJJ9jWfIOX30mxIdiCdYgW
PoaKcLT05Kq1gVtn5QakTTNvV4DlX779ivpbkSt2Hype5SSYl5I5tu0/xPeVPKG0
jlHFPLkclV31W0SVugOPCz17ou9Xny1h2XifR7Dk5ONEKwq2yWB6jdmRSfZKAJ2T
yF+4j9RRyw4W+GRM4xCLoWB73zXzDcRYWPHTAaqTNAL3AcpWo4Z7WyFsQbAtr64G
KQ/Psu8tcdBCbnl7fy8Fv5tAp3ESL+j+s42fJnAb01urUi+A7NXWp9p8Fn/cd9U+
fVLxyOD80ixyibgzWdNhu+boutqZ6NKS5J8wE09g4Hy6vsmPHn3wogJ0LZu1mxzP
iUWruXRU0SkoUrHt9aO4T+TF1xMqX3cusASxHgqgMF/uawtq2/EpDyGg95fX24y3
0UsnAMH0iS7+1fgwyn0LSHNieb2fUrY6sUNoFf03kr6G2q8nT0NJkOt9TVib5nze
uDaOXt5ZEvQiBSn6eHJs/ph/cQiwGhKtUwwXOIcdIf0gkg8pfDjPCp6UDxsswn3q
J59zqq4i7pcxL6Wx6ccXERz88LFWpog3VMhiukSO8byE7P8uML5WPqNcfJRIVpij
WGvL+ZrRE08s+1V1yXPODb6528osu2ok7KOyGEbjvItycbsyzfmAPHySJ89NUNz0
3gFK/C6BUUH+EH9GHRCQa1kUXpIeFnh3AjMuCS8tONYnuRZnRK82S1xPDqz7iKWQ
GFq+UcSPEoB4Tp61YWyXvc0u3qXHkNYLxvZYvb+kTQ76qsmgS1jgjpE2d0MUciIx
gNztZF259bzuRe0iIEkeGIJpKnRq11rknQJSBJBI2itWrIm/CaDp1Tu6XCP/bYJ/
4yil7lveVhTJq8Xj3P+kXL70TBGkEx4hD09Cs/5R8SPOuYSs2AwjUOBzd9QVfD9q
h1AXxTnecoNF1TbHbGIWlR1/tVDO2QSSJvTuVWXxMvdZs3oXViMB09g5kglXL/T6
WVMMUTBRFg6EJ+OFPUw5lxzbUsjkvfE0ZKSp194+IK5PANjEy7ZRLvZKhlwfeM4T
y6jVr5Tf9noSaTPIadgxndhd5NkYVLo4VQFKpS8pe3AS7Fj6jS8Eec2qLGeiGPxF
fh+D0Gf6Kv8PEdTUnsNx3H2BjSLwUbeetyAmwik3YuJJCZbH1E0FverESj9eBYmn
/9tZYtOcYNnahZYW5fg6UGHlFHlZT4GdaOxdI5C4nb0noQ48HiYgI6C+V6Vr4UZl
faMhfwE9BSYVuTIlMXWnn2VzkvXBgZ/HZGnU8Bp5oFeb7iY6d8Xo16DyF77YmohP
nZgnuJBIZYDNRLPsbJSyYY3pOU/V7FdPOwlabb1fmL8oufsG0hwthf5TpIQLgp9a
upPyNITiSrCrEevApq7FDcgOew/E3lA93Cnsm6CppWxrPbIwSxeB8meYh0e8tBRK
fWpUvHOr19VQ14dsE0Tl19VGjoAoC6ilmiZyqsa/MSRLQF+jEH4mOZNZdYk0MaNK
0CUXY6k8YSFZHeQh85QqozQ9q0nH9jHmsN9BvbvIiFavV88P5YYn0ywSpHRXl+AN
iJpec/TrN7bSgUOLZj5mx13plCtUpL1hwXkM+Fklhf2pGqUSO05EGJ5sJUxnY2QL
GdcNFhJcjq08R0zfbmRhzoU+1iL5tRDOygnTf7vDGQ0MO5zEjwmsdMlviEfJ1Xv9
UYpkaoLeEEgn7Tkj4c4nWRdTD4KSl1nJGtZFUOiItJERtD93oBsEf1cH+dm1d2IL
dCG9Ugkl9ur1X86ekMxAzckF2H0VYz9Ewm0/C5J/Hh3RvnOR7wDZ3h7+/daC8sgn
J5FsZXESrNfLpKIp9PpCAaR7dDV/Dp+I2JiTMF4qKtoZeOtZOJ4+7rS87+YPFT3x
r4HOU7X3fzEX/7O/Qmt/dutU2GiLl9H6a4xIgU7Fvx5FSXHqgClrDhkFe91L3HN2
A87oR7hc8nQUk5rPbuCb+2vjSGId2iw63h/JpPkmiEh2SZz9szGxrnRNtP9O7nHH
RoHKuJVXoHhXM+TictfQ4AnILxgIylgJwLvpJdexUGzY5kdWgxOSg7ZU7CAX7Mfk
XVx4svW0gecDoMyxf9ybpOeEYfWTxhfFGKi4m9qxv+Ehk6N9cZ4/dpcuE1Dwz3TC
LmfglesTGcEWYyhwzOK9uuUXmvxbT1ggEO+ID79jkWnKUO3cg87HSP/LnvhdDql1
5t1J9t1FahCB/vhAU0nCsiwwELk6CIPcemASDRZ+34ha+5iGgAL2tHIMmP8ittKF
4SNshuhCvnBWFYCYsygDovcoLgY8eqvKZJkAC9zDfL/CJqA8HFmXaeVgt7Aa20Dc
kT7HCPovS6DK0+2hxOxdE/lG603057pVudMmUdSDJncIey/jPyOh1JMFZIf+FLdH
58NgoxRtZMGEsPFr/0AK+E6BJnuLhSNbMiNtTi/SV3fAJ8BqJxe4rj6xkp++lCcN
BMH5/XUAF95eITQ7t84g+84UsPA3P3GyVjtZtxKIlc+o+zxILex6o20HfLqc/ohu
NeGAHefTizGMatpApDhTpvvCUGIugXThsfL5lHPhzo4MDlrJDwBq80C8ghIy5LXw
7Bzin0kezkncqTezm2afpqtnT6uyoqZn/qyTGZbR/achkvSzXXQO85ise/7GdSlk
BQmDN29m0XXAhUdYTWWSwrC+k9ocIywxY3mbj+FT+QzBHVrrqbXsA45wePxMIj91
ogt3VxmYukLcc91yKEqtvMqHnTQidtAvPonyvqHICFPKwDNlGM5WrOLmDqjsSYeq
l+kjpZjo+84m0AzkrAJ+DCSK3r3M/s/cGSqkpeirRgnPu7Vwq+CPxa7V1jQJFoxj
PGlFL9Q5tYKifLk5yPkvS0deQpVheU+rJ0NXAG8H2hfZwCYsKxkjqRbjqZrygP0L
+FqU2eE6DQBuL+ENI7fndskxDr6raYr+c70SuangO1F2Srg2fYFGhlHDD/FHHyIE
R9MEYoJFGdOBKtUt7LpY0egxAZXcLUdnAOW4jw9H8tjdvBKDZxrltVM+PvHVFZvi
cn32cKKjfaXOOFew5KE/4oG49Q4Gut9KNC5l5LwoyiRLUyoCk3vMYFMIKHawfbA1
0J6IlfrK7qYbb0QyCvBzNyDmtMx89mMC/e5En6DqiEq9c3mZi/7U4dybf3c/n4wa
WJaRvRNqzHrV6i4DjK8Ps3ddrK3RQ013ioWZ/2sgNjyp6FRcood0vqgUoUD/zF9z
fW5o7iAFiVdTo32AZsmdL4BsndV6fBljDt8z/8rTm5Ng8yRy/LRjxlqY0K/0f/Ot
/v5gg4zZ5RELb4V5m3BLt8ZgVVo8KN4HJ48JXPiWrFkh60++rTo1b42tp/3G/TM/
vg3fp80NUpIHdOwT170C+q0XIAPCR40U9aPd4bm88PbCXWnoNT5nLfKpqmuVuNxz
CrrSkhFOX03U59Yk+xSe0hsrNcau2erDegUnFAR4oXPiAR4qJmXHb9QVUITLBWgL
Cpgg/HAtbtzeJjZGygA2sNtSaqySSlNWDc+U1vMrSjJYHYgYsUrAEEonHFOmrDE2
PrhevCAdqAcKV/Yaj/uqHf+PwsNljdgjFfRN52GkMzigDznxXBXql3m8m62wVYFR
Jst/GZbn8uXqixYe6f1wUgJzEo6V7r2+vsdLE1Lx8OohSOIddxCtGRyXXBKnmlum
KzXH/9UBxxKycjsb7fzkF7XRlNSBCrfinG/ibgSngMT04lId0d7ATOCsnsK+2OOP
KroO004s6w8Z5XUKKrhDzB6QSrQ7flp6smVRBe28mA7VfXmfPb7pioW7dj+qkWaV
rjbNy1/zS0IFjzOPROojaW8zKXgfRBGsRDSvjX7EXtt1RaSLsF9clAgzXqBCf716
6KHtDq3ycBzqxUaDlTRe77kIcknTNUCdq7Yqkg2j6xzc8j0HwzkCxhieX+jOL9gk
oX2JZs8Sshc8itvSpJbvMtJvK4cjrkqkOPHIgHoLE8MAdp+LjSEtZ4cJp1k3cZ0J
sZHbwViVsV5kIcAOSivn8brocxPA/2YNjB/fBAuAsFVjDNVhFjepwJWOEYM786C7
bH71bbxudWTwaHzS5UG57Sakyk3G0fKOU9kcILuFo2w5QGhdxXDTnBkJfz6wLN7B
zB01EUr3bQ8tlx8kKrkKVErk/r3eLgZo17QRld3GWOzwjmD5krJl4/yGa0R8lG45
OE6SYCOIfkExDZrPvdmQZ88hxdQXXdyxxelP4K7azb8uXkQ5Q8OSN66kQ6Js0lyB
LPz+WoaGt0CYpVNo7TZ7nqFn5hrlQdvDLrATgBizlJ4dhNAVfWffqV1zqd1z3X5F
EHcoLRnWBqK3nyjGAQw2P50kK2h7vks3tAIpy8KaC2SkddiN47aB2g4hUmWSlQef
d9uWtmt6uU4rcRLFkl0+zTIjv3AhBK1SxIjCvxy7j0T7/31ZXB2ZCBJSn1jubJCT
6pwtBwvP+3aAQNBz8eG25fjIfE6bYM2JGIYEpt1MzJWj8WHnwZLjximare7v4ftF
B3DZxe/hi78zmaJTqVoToawBNGb5oR08eDCIDVMwP7Tb3km2SyAkpOZlaj1WdYOb
G9kub8jgAYp/suWqGFl1wug1Om3NQrXUFvKwBIwnZf2vDGNgyUoU+M2HOqnzB9h3
KxW4SGNdQPtL7GUIo1m50mcRQK84UgxzSkgS1YX39wqP731AzTSuAp49+aWDtG5g
PRjBDEmAGbCLN5fdBs4wzR8Z9F5SrzjW8gON/B0z6WErz6NCArhrV5VzmzoxChy5
zYcOq7329bBE8zfxEWQsPDMg01nhWvGbGY+w1NBuZLdVbiS6F4cLHPTNZ6hDJNfx
D5UgRmHBmqOm5+pptDC6EHrbrV9lms2eCwbaOKb5jXdXsQGrNb0C4UKiiEYSA/HM
EJXtH0Ld6GhispnGd2jR36ekpW3x/uk0XRsWaO8hQlLwNXmucrFm4WmFD24bSKkh
IEispOgjPBgQ/6cZW5KH30weOj4VPPdjjq5OCr4Po/OwB8jUAgMOXasMTJsOkEUB
GMaYSon5csdpijOp/R9LmVcJUiUCrvd5I/wMED38cZvHV1Dnn6KAA3IVf4wHmdMF
tyNxsetM7BP44FVMvhM3eGhVzTCbh9qiSjpeOH79XlhXcSjzGhE5y9d9k3+66J04
eUL8X4jyoyae5FrlR7M1VTOx/01SAL6MdhlZWv46mM38bL1pgzpOOXicL2Gg4Fyg
s/ErqEC2eBEsG/kv1Ncbzs9xthl5idzlrxJx069Wzm2uU2+z6xECmajXfZoATZsf
Lag7pfVD+/fzbFDlg2rmjSdwRvlH2QcQLtI58m0HHAtqMsv0zB89wa7uEslyJYFk
vRc/wBkh2jOylMoA3tljH+tUvGbY5o1XckixTcZcLWzF787GWSD+34myoqKchXZR
W/nI9bfP9lA25P0L1L0OGM2+1IFAa09pwV9ETpVArI4YZq66Wna2DWy3BfMGxJV6
J8wykD0MCotXWzLVQhYEgBjj2hygcHpGAj6FyJ92I1rdKTHYi10eSQpoP37eC/av
63hjXPgdD/OGnEzijlRUeeW8vU+kptpPoEq26jPFVtnhaU0VSzAIQ+flKfD7DpWP
JztjPfohXTnCT+dBHyPmjt9REtnqdlurWLK9jYfRs3EuH9xH0msXZ0cbX193TON5
DZmGjeYXOrDJOvxaJwyR5iAYglqWFBZGRe1V6wTkjBpXWmxwcPslqcwpHx/nRcuC
H/sBaWboCRXeGohgIdEO6Tugn38+DBM84FLTpNeZIgEiIujzM2bS6EpcbArP53/3
R6NGi63nIqLVWEged0L8MqiHuXT96i8ytGeME30BquAp/w5ZXHS4XUDbGUyQdFgz
u7E7HLzsYqpf6/21Ko0Nf0XN6GUQch3QIzDP6T3TLIvjGs8EnfqQbCgVslJfKK2/
sRUzNJEAtA5yt+WxEql7JUwbGxHiWefrEBSXZ3PnC1HTLLquce8OZvWxrCsdN1xg
be73zsd7xrCLLgGcfkOj5uHoUZIadjSeFc5+zuCVXDWbyGO9HmBXnG2KlJ/Zmzhz
jGZClDiJik3FZqHf6263OzskWNsU1IdjYZXaMkqKT6DJvuLf0OrLMXOW29tmA13E
hj58blQXhL1GAn41G7uYWsDBfAgJyaSQLsCDIAuhh7uMnvoS8OG0PjEdWRGB4qzD
7ClI6vMyHkzL4Lh0lBL8izq3mwAQcIvVPMkQxFc8jyQ8EMKmmYVvFfHOABuuYptY
tJM62z1y5G1Xnadf36Wq0D525jIR1U4sp5Do38D8kDktbe5iOcpRl5zr+Y2gMHde
JPdjzOFJy0UDyas6gCCCOgfIyJj7mWHosLs6zXKeHtMHhG5nGotro7yvR1khwA0P
XpC4PfpQ/0IWnStaN8d4aUphuMWkdwPdcZwhnc6qh/nhor8WOb7H5ncr/X9WCrqY
Nk+Vxb8DgPy/jBM6azpuzmCW4oWsGdnFLuraKTzTiS9fjV5BxOLKxCw2tZSvHpji
T7h4rI5x1zJCKCyp9OE8/m0uVBIpRjp9PvhEb474OtX/kNh18Sf99S3/yirnJAHm
ZUH0jaDcW94vQf/tACBfvhaQbedrUfSWlkPSRt6xc85CaV3XvoXUW6o233EdNuu8
pI40luWarSMUyI1RrMtu/eGwSI+UKW3h7B8bXkGNAkuWjDSCVZBMWSs1z/QgO9UT
IV/4eVK4HP/5puMj36GcQKyiGjAmj3YsNONnSfNOY7ZDwYpV6xQa44mMgXW2N0c1
ymMxiMZFfLPKwjZH1Emp9IiXqSECqpE0Z2igDX3Qn2ZMpMmdb9Nq24hpZVgpBx3+
MzNA1DPX2F9D5w/s62XstF4DRMP0sCZnnWanGKSDtE1BPomS1IiujjStQxEW9xXi
nqF0p5OjRiALHjwp1Q/wBZFox6um+eipgaNUgu0d5L9SJW6LFC3pkoL4KMiLCC+d
BrK2QApa2l15/kqR+if56/Mf1Nc2xjcnezLBgNg3LWGlBoY7KrfMqScdHmqH8W5G
qbZ1bE/3lVVm51+MWA8ME3p9IrWycj/vVq9Shx2NU1sHvRFqwYUvEIC97mgpywQR
cXPMBGh6tgHP6bvCRCveDdTKbxA6f+Ci6wrbrLQ/AlqGi4OQKMOibLztZxHkIio8
DAG7vhsNy6nM7PCTDanyIXjSu5x2l7SE2SKBweHfiL10w025Vqz/1HEr8M/R+KnR
qpwADc2WPZP+VP/b3VP+jrSohh0Bmo4JlwrRnvVOKwgG61SstTISevRh5HKR+dGJ
+L32eI5yscEne+6Tbv/Va8hJLAi/Yu2rgK9kZTjsG9CsO3Sj6Acbid5l63EhnlUc
kNR/bWpLUJhqbdL9NpkfEQKIZKajwD6g0XzWCrbEkIWf6EexTlVoRvi2liW/aY0y
rwDYljueVsQ55xGj8clIpZ/zqAYCkTULUk/lKKNwPrkyV5xiTv5I6/JkOiYaLThF
jXQIQq83WPwO9FSzuoPnZdZidC+78PBr92zmTMOLdy/dMw4CKjaS4AzB0yqZB7Zc
Qf4csF4suVHIfGiRfguB5ItxasmNfEbA+GvJo6fYRh7RoEh9Ox3eyeUPLIXT4BxQ
Ww9DOBYzOhP2TGcZNHel7aC+Cpo3C2uUgUQrtwbVARjZUqOghcSXyf+WJv5k3qcn
NBJ92BEByBvGX/a6gg1sY41h47mhoij+KOeRUSd0Zs02lIyTcUjVNmRhh2Ny5tG5
kuH5DRxw4Q0vpdufjtyQutUc6458n0ibuDocVmhSxH/tbZCmC2rkUmGKTSjYxNjk
3CVlwRM78Iu6TnIBZ4KXBOHGWlpAIrWzoDa3hjOm0RgbHLY1f5ghfUDzcbHNgggS
VvZ0mdCmd2yw6bVUTgl6aSXQVXdpVyHiD9a08++NAfhpARDvEC4M5HO21Lqe6Bm4
tOq+zqk0j/umXRUgFMGhh2V4wfq/JIpdSarkZLlq+cQsWWWmEk9NvbpwHgibZbq4
N+V09REtHmcCoLcsXWIIyQojUSt1a5b7l++wat0IW+RccEk/Ho35jnX+UfnXo1nc
ltjdZUcUIaNsmQT/seaCH8/oxwi6xjVlBxCu3qR9mP7l9uHseopcsjei7YRdkYc9
5YARmIk82LWAMzP7s6Zva86yz+95HQZwxExprhbrb37P5ZfcicAx3/974ko3nEk1
6st9HZb5ZKiMFC8jGtSITWRvjNI4ULLPSQR030ryV2ZX5lfBZhyFVkSzgRf4N6xA
0823Z3fSnQ58hIKZ9CGUZ8Oo2nLRf9UHcEqheGSp2778OxWEZCKe0JH7ObuEn91L
yEjACyXKerR7t963GQM9LC99k52+3Nt6OUSYv7HomsWYhaOJoVtr0lE04NGtg4Qc
bPG0lDGbcO3WUdpIJbZJb5rjSA/sm3fBytxzdA2YGnz3dAFJHnJGkq+S28BZ7hTB
BRCWs+MVvTFXzUVYKz/uMhlxGQcHcCiRmZDVJu5lt5SAGAKCC/yKSgziXKsxrxQD
7LaguhdZat0+ljlwCCVoNZp5mtlrjbES3EblMIoLvu9bTScoAWPdIoESM1d6rx5+
iYlA6PZM4Cwgtt/ceaP9xZK0NdugIWIYFFRpDH75Na4QGngWYEte8Ji9mD3r+Qk+
Tgpj9wQdOrJWOKmZ2lWf1WFy5b1fscZ/sFta50Wq5+3mxl8OienxGD20LFdGTgbq
6ELFaUM5lpAzGAK7KujQqYMnHgGyRYuAM1KS6sy8t5xR5o6pc3C6ho1LBOWSGDLd
BhOD8XtRixVWymGo0HOdWAmDIHpdyS5O/pIf34CeLF023Z5B/LT+zo7LSK8foRMk
YroWVPlhajRw27DgkXR3A0f3vjkdwmgnmh3aoQCo6lUXQYoaGi+CL3IGttPT5zri
8XJaDTJuPlrZw1iHDjngn37c09LqceEf0e9722WNLLz+028Fac9m6CuR5JTur12P
KfOH6jFG6t4KbT++WEBxMrcP5Uygvg7obQZ1yPD4IOnB7Hqe1+EIyv5/yoeeofIY
CNg5LI1RSjpq4VuS+pqgslVWxG2lWTUvwh33c65IpQ2yVHKw1gvU7TOpcKtTzi4L
1S7oIZzaYMrAKol2CGch0Yn5gD3z9TtsFEnLBv0FhTkMN1/beK5qkDWVqLPTIci5
xxKKezpWN5l9IrBlERLcOCvvzCoQ6DHGA0T9mDkI8uMhg+Rj4in1DmidO43SXYMf
M9Q6kFAM5Gdv/535cUxthu4NQKSimwMa1glGlEISARzcaWJLES1wgxLIzbJZRGBP
dxSk6QTq15GIdjAwuq2rrXv9WnVjMENg7jFEHKGGd+1nJvr1gDDJUGHxsK/8zNce
ejzOm8OXVGSNXxp54wnlnQMnicV+YRLtKiRYTmBWxyB6pevxljDAdwCNDkUeAZGL
m80BkB+SDzZlMgV5IPARkMs2nnUVC/Y0/G8z2jOd5as32FIhQoTNVZMnPtu/yNqq
Nq3YhVnHiEs5BICJNy8inxIBYvis1zwjbnmJW3frmGfq9kpnkXwcJ0hD5e7sutLj
H7Gf1vmqZE/8WqR1+IBo9UtO4UkRaxXr5dZLs4H6GrEOZNNMR0Wg57qo0lFhYkao
rrpTTdUnR1uVr5seka/KYaidzXEREVa2AVvU7nwxvFlTS5R5A0jiTFNyul1zaXXE
DzKmsTuA9CNFCKAr41Ujd+dtvbF/6Pz0w7frATqjGIlD6Y3rQgIFHBDW9OUucPiB
nrZmGRkq96iG42U6hTO/G0zDqfrLIThv+cUfoz7isfCU7gWehibcUfmSUR6B+i5F
MfBG1yC4+qBYs64+rRQx6hrTj7jhpwlflpZnR65CfplV79wZnyWKpitgc+Rn2Roa
JW13GYAN3yRoEOMpSQVOJ0VH+FKxNpUUoeRTbluHu3xVKYuzBFkVMHmWh69acLIq
uzfMIKhaNRA5szACGoxwXWljkca/bK5wbBi9zDACwtQ0P52GKBVIYvgNKhEWT5Ib
Dzcy993bvP9nTJxGHYGLGiCKrDZuVfpoZp4TUSPpSYs81VPuZh5MDcw/IEnNlNMx
Dq8E4peRzfNjb7ugQEK61GMIhCek2rg3DMS8pqiMSgGKMEkewFBI5t06au5iIH5c
1fVTkF3+JS9+UyLI7TgLmq/fuV6r7SeBQhkf1bifbZ3HK/KChxnnb4CjUWPEEb0O
MzGJqhla2HEHjx8PXc3BgezTWixFECTVjtG4fY8FGw0WOsrQBtGGlbXqORW5ScA5
jXzMIXdY0uzGobBdPkwG2wuivTquyLjRVle4U/FtBbY7GPm/BgS8e6n6vplb87Oo
r1csbEhM45qvzJjMq+H/A8b9VvZQXZpTkRBuIvFuokmOJDUPrZLHMrA/qbaswKwl
5lbVmj8kQNomDdqzKaUPnsNg4jB1PPNjiOZgwc7vW+F9+QB+nkSuFusGP2WzR8kn
nM0xwlkOaqWQhcEnRIsgXrmMutPI0qgdC4vssIMgALJoTs2u2HU3R2NDwfJOhsGG
pNmWVwOcLXrPoIH1lzT+vXrwOiOf+0us658XsJN2qIiTFYYeITuHgxmd0rr3QtpH
ErXHACqRoxI28Unm6F7LwbeiLnmbJt2rkkNDnH3EG+cH2TQQJIJLtJb8zjKXVMAz
HYh+e5RXO5nIm4eYWgOOD9srVyVyqyLT3rn7AP2NN/ZRSwAzHcY0t2QsHfZy6XaP
FaBOOmrLGOELhplLwLTpky66BzGQK1ccLvGZxjOqd2N4nsjnOH1g8YHXF/eJjV/z
DZUoViko72rFowxnmEofAauzLhr01IlDo/CcbzCXeAG2nmmz/F7cXvnVlwM0MtHD
fmnmsOT6D0kJZTaUk9NLjhPIf1qju0IAJipP5BKz7BwG7uy4JP6qaygA3+HvAgOn
9Czv8uPnfD3L0vfAD8dlQd2uwJDiWpEb0LYnuvD3/o33Ldihe0eDivrGBA2jL7G9
JfWpqYToNmTBxEGbcA2RwxFDKDE0ZpTgeBNfmiiFS1LopfjGeKdEhNpwAXa+3YO9
d1KJarqaAPQvmZqicfvQH/cWTWmq12ibOwKUeXM4iVVucM+0lSjy7PqV2G0WzCJh
if+5Y/pZ5i4uw/09ykjlwSlj/EnSPycnLmPd8bO2jkoECfCNO3Ef6b1tmeCJ7+eq
Amlu2RWPKZKW2+hSUVccSrcc93l7mW8Fp8vdKch6uQrLSgNMePb+WiW/Uz0JPgmj
Sp2bcclZ/PXhF4LGwfKwV4VvxBeF40hCISSgVJVafNxdGadKGAViPZcCw8tGKZJo
U0uG4Q4Cco7E/MEAF0Wqn4f+0+mDWjjRW290W48B2nah6H8Y2VyP0Oo8tCpeumc/
C2c+SaYhLojaPIV5369cULz9ZIeoc4kOJvVSLnr1ie2JjoKUiXvZ4S94gneio5pH
FmP/hXr8XOksO5c+UpiU6FGA+qdXFi233cV7yHdKc/Bl/Zog+J3rsccuSkMv460Z
ryFNKvtQ9n9E1Zxy6fiHMfLOv7mytTrcWtzuLrk5k7koj2DimSr5/PQkFBXk/MTx
KnjSsW317sI9LCWxIiQJazz0C3PRO3SZP6pVf6QVj8GXLhv6EnDin809V1pH9PbT
vuaIbDdm61WjCCx1hnswSCB6os02m4SB1iUhzHETm97NeF3/Wg37xZwgLWINLMRu
RG1gsp1QmSP6HjUxPcAgUpgS92FkRo5v2Av+t3ASVnLLlxC9g9d37QJGeIh5IjHq
bRP5iEO2ZZ3hTSiqqUX0tCJIBOQvqgWjcuXYVK0sVRpuLxlBPxnLs+uR4vD1IpZu
5JG0gUfYZgVQLMaoGCbdzYtol0fq/4xewZvaeyFA8jco9dcv7+k3vhhLbq2Ts6VR
0lklaEqNpP8+1uvqiQn4YcORcOUNnpAhBaDTUbIVpqgmmFUPKGxuHAabqQjotdKM
SxVPOrHFzIou6H2hzg2l/EDQv50zYvO4/iXntVEwJQBGfSe/7jkUzVQHjuDHhRq/
bD1fLdNg0tk0mWUNXLFIfxeODoA5wbS2aTgqJVpct4iLvcPVRTumtbK273GBAEcS
uVWKRcIKFDVFsMC1SbgXCF5gTNn/2Yn99utUGKS+81l7K5IlafP73S2MhBbqkWhw
dtZ0VQiOz1AVSOMeu4YGG9YdQQyoVxbHOTyxQJ1b8TxrZaAZkrST4fwxVDFuxcv0
p0iYlJdLpiRoamRBdu1HSxtOZr/wD62Z85VuZDt4VN3Hz0/JTr+O4/iUbyHN2zN2
xJDlyWZz8jYhuTG9JPrYOOYvU6704BJftHilLyD6dF7ohS9uELZ8OywS6kzmVeeN
y1S619jU+MT3psRBrtWq6NYOfADBxelu/Q0jnh/sddHR8ZfVdzKaJsJZLBzx7fem
cRR1PYHecBz6E04vb2H5BkF9hrfU6tC9WQRbfxF0VQBf9aiyNuPWnWjt4iSgpTui
Bvp/B+WloxPT5W0be4jlHabOftrLFL9neb/DErKLsbqqUqcoCUR3mGvhsNGYwYhs
OHLgnTL/T3xMgx+kJqkd7lTM6IquavkJAHsYJf/0uRJzgXYUEISX1CbIaTaYgGQ3
tdAy9VrHSn50Wz91tEpboC3VxuoJBEn1G3kZ5+IQHRz6PRF9K+7SStAJMaiHI0GC
ZOBwoU5jUXdWJfO/kZRR2Hr/4Msf6QXQv6MJGQGjrQoWsCv5mGYkcxl42RRPKv+F
tUBqTFbBF8x1UtAN/acWMCVt3ItfSDy6Gbgk05LM4sEzFdM4Szua0bSc6GeMnGcq
o1Q5r1vk1QCskMBmmtFRf3Ax853OZZ7mFKCNhJflYW8tHfzrXXZJFMUYRigDuNhp
byOeJtBXZGlX9P+ePBrA4CF8nJ2xkjdZxmC1k4GQy7lyvS0A4LFAv1dyb6cSXIXI
lsOzZfGjLBw4VJnktH4ZyeeUuWW45+DBCLDojjGiwuZgouKIzeW3CuMIFPfQVojO
cI9u/3B+SrU8Ht7XbzbBzeTXRGWeDGm52juSx2fJ8eTK9GGixRLBKJSfbGzigIdP
tbCt9EG5mJmhRflKkjGaeSpjvt4ymCbQS7jcDC66UOHD6j9dlcY/JpQYJBpdeZBJ
0XszJaG5OSHRsM+gVAGQ6hlIWpdrDL4kHhXgB6LyXzPtwNeXQSq3v0jcpHGhFEiA
7ZRUThWI9ZTyzW3bAlmFTYMbAqW1GmZfzstrRlx3ld5YL4gXtaIlZ9F8HvE/X7Jb
3jhSa3owLHlB+FqWpaot9owQea5k9j/jyvN+LfV6uT2mmFpqsaCi/yzu+KqYes4M
acVrwSDfGnBpOopwwbno9e5e1sH3DvpAlhJ6jUqkE+w9GGXN3pnKuID105eEE09a
1VhEaTa3U/HJR7NmnNOnsDTUoyDTkUYy0ksom5aVQd04BIVLQVPoLOopvZbEbseu
w6eRNsBhbrl8lx4N5Y7sC9iXqLKT/29uLChoKVbjUsysT2zNyKs5ev1Jw4dhTFr5
pGoN0yjnaz6/qECIJqQH9pYtKq8gb3EZRgfSIlF0+vPlsq7iQlrz29lWkqsDBnay
haKSicEuyHYvLpbjMWyrleYrMBN3d0U3WVbpLdPfBTbUGM/d3F2cVgdJg2dWHehb
yMyU8mEFA3zIQGqMN9PmVRFY5FgzyC4iPNcdA/UMxu+Inv1grQBk96qHVE97h7Md
KDZQnsg8WRcXyWYIpqw776vNpxPq2AnIgrEIxrFB6QOiT+3qxBKbcLaPEQ0Fil2p
L6A/BeazD2OXA23t0BofP/ps+AGGVfATfgS6msYImty0Z/2RyZtInmQ1Xn7sawrz
Fb3CqNn8e3iihqRSQHO9JKNSw2I/plVuAPmWWgCA3hzimn/RFHU/NJaF1f0mKnhB
XRmJ9OmyFxQJ6fF1wKRy65BWLudnuhED5+JRA41a+AJ1+dIDDUFQxPT4hDtkt96V
2C015vr8BsIx0vs878R9/4Ca97zKhXWZCvg2iWJvTGPBmQIrnraJD+PI0zgJ2jN6
4/i0Gg8Ocs3E3KUU9qV6fePZ3OMoeDK+xcNiA0JOuio52VwhHoTtX+JBWQvI+NfS
tXIcbYQKUQcAqOl35WD4Dn/ICB3DIgjtDvVeorGn2k5uCMJLSIOxAR335lDiXIao
LNmZN9TnJQfXHcEpQ0Ii2ckznZdaAvqwrM5KTNnEBNMupxI90MyIi7zLhfc5F8dx
w6GfvB4XgQzMKx/l2WI/nMYEuHEMp5sFLTzlw7U7rluywNiJ+JVvwurtXwI8R1VJ
l9i6SGKikoCW00RAOsGxIhgAsmcVf+NkoYgjf/GZ4ke2rvHxS8e5jcJXguLovXLR
GglpbnHZMJseMlQounuo+3FEH9FOmIu0rQStzvbqApQ77gKwuDnn1rz/u+ARFpXO
6WVGie5SPuWJH3gk084bj6K7SxFBeZ25EiLMpYs6FdcaNgK9dRvt60DRTUxtdPhj
TX1XnHUOYhCfw/y1M4sgd1lJTskssh/mji17dTZW203EhFMZd1FEHHW9n1Idc6lH
SrlDHlz3n26MASoCWjT23IkGOTjPr1FX04+4HtKohYs2d0dDWZdRQ80UF8RqND7x
3BMpw3yQQ/RYuXK1pIr70X4Aidfcdm8yhS73Vk/dWfKFB6pxOic9IxTvjgcAbeNT
gKsXjCcUWHv8IlO4uPFhmSQompHOBC1kCFT5J2wXFMpNGsX4Plpr8Wo78mNLtxDw
LMGNfopukWdYRekCxUZFQzG1fFc5t3M61vcmP+FX3ZbVV3YN9XoEDDNqe6Ktu79X
gZfzqlrc3kwT0gqbIJ9B6pP2Z9cNYHywZItyHLAqK8G38Tci2x+uzp8Pf+suQHO1
DPSOwdoE9sF+Nq7hoWqX657+YWn1nTLyQKRnbJPaFjXLw/tLqnw/pRTX+NVPODff
knVHIhnNJy3R+DI2lnuJDqC22Z1mWlSOraaVEFGdamCjbQPjdsgs+3G4qkjoS8Bx
m5CJe/LeFTFGgFQX0AV6ItYOj42l+X4CdQT3AJ+OB5d8v35/klyvSArydB9tczm+
UW0YgP2FtQW84Vk6BWFX1vm4NXmDjMSUlo+iijQXssqxUckm+bo0fPLpX74wmtDj
7WYoW/G/Fn17eDzTr+jpySM3Aijv3XL83+bpMbchvbNjK0tC2A2A1VT3xcnpEVjr
GU60WEny+hSyFaiduhMxHDL7zqNxQPJqlAarH21/o+9P84goE+GHMYEl6DgGHssZ
hGVjgpOID+LHfLGFosOiFizRkCDmIW3bp2KV0IB9HcniurvNgxLnIOGbhjSLJjAn
5gcn2fqrFlutogxy77fr4/lMcbDXCrSEUzasG+LbcptPLiPAsTYqdzE7wdWOFtV3
KkeN8ljD4H/8BW3aiezSlyJp3bR3Tndl5UcJyP02x9seZ5lHIqf+qqV2aDnlHIKO
EVIX9mtemgF6ZsgmW0PKq1OJPiTZTuuyf12gFvZeqW4bnUSbKy86frKgPagr45l8
DQnHv0/a8+uvmOU5LdERBltDNuFvmk3Xdl9t/ZxLGKRJc1Zgdj7rkEMVNpP/6w3o
DurcuX4mfOU33IybwOghwpSk5AVSnuYstV+ZXJUH/enlWG1E7rRcL8a9UcYTKTHL
E1dJc+rhday1PLsBZq9ZrVkBNT/wZiy71zW+uPn+cTks4fMNDa84zkazhQ1elv9c
cT8DCi9s6k2BkDFT0XtBHo390sQ0iPPCT5IGebZ9tRr6VWxFbnTAWWAEpQuysOD/
GplbzbVX3M5EcuA2zoppBvV2Xxhxpp1kbD+2vqrFGrbC2JrbfOFw6QqNuMUkOJrV
Cv5hv3CPo4O7rLKbtkqa8vKBuGPWcal5KHeBKCbyN56yFxp2mkX0mSCxluJO1CeE
79xMSsbjhSdRY7jc3yAP1AUPSsPMmAMDORb5UNJOcXdNiogTiqjWnCw5D1IZ/l+J
dSkwIl7SF8Oq1gknDpR6l9ecxviq+1+RKmqxpxzqwSiXm+6u9tsdb/aHjhKr2Drr
5MhWaW+dK3ocw5yDPb1jIjTuZcDj9hie+FrLvRYqBCmiK6UB1C3JUk5opQT4TekG
rOQchzb7fVIQ5rdcV4RaTp1Kxt/eJX8iUd4d6tROwxwAcMPgVDWkugI9oTvnKSYG
OEONJ7IWahb6FF66yavfhhtgYphQqeDsBEA/akLFEVAYPmVttMhmkl2Ox/TBMDEB
0y1kVupNnNiLaEffoFITVDWhVFVy8095QbpAkQQKC7ekajT3zbtyX0mxSbXcUP9A
26vB8NG8TpyIuVWtIgclOvdJH2skLi5H4KKfJRBDhVmqC+4YEXMYyURU1tNsSqtB
EaZHrkIeSWQiQICpU2Z8xr4+ecHN5Lw16btw29oplZJmW8v3b7aFHL1PvK+nLxbY
XqpNha0xHHiB/9rXTS9oU/kRs11vakNOlv0GsSqsAOjT8NusUwwJhEDHX0CVBmDl
fDXDzoRwiIgPd/zCCixvE658HyGJJ/jrQhZJZdg++6qt1RGLNONKq6y9xLw3QEdC
ujvpYubhff2Aq8cJlTNu0dmIXs21b7u/p/yXszlPST9thiOp1SCf528GCRrvkP7B
y/2GPlpzH+W64Ii8igUn4ABVDjKXrULVrGJyOR31LRlXSea0wTgV6CLfTcFjCIP7
xHvjQ/Q0OMiQW2MmodL9RSxgk0pYfLKAOu3m+63Y/FwC2VhnszmYlC6NT1ibsLmu
CjDpJ2SMYxeotsrhdEmdNYfu4qbUmMqF9aVrDHKJMKkqggkHRIFxdzwqfhQQYfRQ
w3qCL5RkV1h2VKEipjj0XNnC+gj69CyApRZKTlBaZqq+jHHlzAOF3XcLBXIpNXil
0sIZgWtxSwlewK/RrDoJnHoW8xPlG6P8vmZZ0evHJYLo+qV/E0Xhy3RHek54NgkN
CbAXl7ClxHB+h2RptFBDj3hjM9pyrLORISmvD2Xydx32HSlupg9dOaZN/7gmsGXS
VI98UyVdFGwnSp5ZHPjsERjbiKRSMdTEiLg/8tPqJpX0maZGVs1S/1C1E8WGhKj1
lq9zgHel6cyrPbiz/wR2nsRcaCKKStkLCupRnlmTSAFtqB0Ta299D3zcsPFXUCnG
iFig0a47X0YQ6h2sKNd6V6JZOVfng/ZGNkB6Nqe8QWErIbYmqnJNQYfHwFt6r9dL
qqL/p5GGum2WzQ1GAkI9DYFBBLI25O1XW8ob3nYCiaQRYQmiS9aQQQVGMeBYRjmk
oHOUy/l+3a5xX10WKroNcve8UZkg4zy21fHuaPNJju4/LwLDhsQwiwf4tUCiyvGF
Ue7GvCK8AGMfIUCEHUO0MLjhCVhO5NDxGLdBO63zruNkuoxBmQfFyJAljFrCw9Zx
USGUbND2G1TI5+q3AMJc4mS6kU0iXt0msZNFHa0JFHImQIg1MAyoTiFtSmaztZeP
YAhFfpFAapfQuThiqqSMZxeo/HS9PUN3Px/1aQpaea4UN51yZH0kYeJOx86BgVRD
G0Wz8DALWl24PMo8u1T1k5PSwXcMqoBm/4kj03bC4qC6Lh6gm4BFhXZJzLFA7z6F
4tM5R4+K5k3MG7KjBe8ybTMQIiMLzCFVMibeFnaisaJydmxfaMLnGEMYqP5zIlM7
qDca/wHSVOuUAEhFItXqLDRQEzxMvD8SiYtKcyoSuMHFzOa6uEesvYAV428TPbU6
+YE08HPpT03CEgXHdNpFDyJNapKUkpYQIsPiSEU55HGl3m2kGtSlTF5HNHcYgYje
vYgSp0hRdBVaWmMs7GxgJLjWs1D2WUgROM6IfXXUpqqTgrxr95RajVO9C3OAOTJq
yJO/K7VsGpfBI9hoQyXqPnLsyhLDh1SpT1Sa4kdoZIaMjg0l4v2PLtIhR8R5h544
3FaqY2E3jztzXveIGwLRR2DZi9L46NGOGof3ggj3RFJWuhDnZLnHzSAWs1TBsonf
O/2/9kA2TWsfhEJKxSfwJei0IInfNtXhIqYWnOppOlbc8JfU7og8qyTDnsmWNsj0
IhrmiM9OCtB+Wz9LPWMbyhzpEvOxsfItqSyTBuzFxszWkGqJOnFrxGkDJ0dweFgT
BBE6xN2BXyIK8VSeBO3qHHJOJL8prEUoNiFDQe/ZdAc0Ew4BuZxDMr1LroQh3z6j
D5hnzwYd40v9qZnsE0EWChPZ+ViI6bYOw2cBIpvA7aopmOwUiQNifTuGn67EzpFj
V+GUWObey9fGuNB8d4FV3HvRtmuR3582IyNGhDVW6sUqsuFMo2k0Q7lVWR4ADqpX
+w0nJIkuVFQ2c5q9YgfiwgRnJ9HVQqqXRDJ/QSc2uGetaLSnA2pPmSkHxt8iFfm6
f5lnmI3iJPnaO+iZvWGe3YVRbZtYue9hn/j66tHgMjdJ+mr+J2gUKbY7HXzrHBhA
CKdV+1dRZ0eYblLPNhAEo4o/nE2PUa9JaPH9ZxSDgkh3hFsJRO6bzH+PyjvRQpxF
BFbpHz5tjwIVXupkC4m7cKIVZaKLLTCv4guYBIQ1n1tFLFC/jvfge0J285b+1OXF
RRdAemIFQPL4u9U4Kd+GMIHaKFvrm3G73M0SwkgIjf1ttDUXYEGOWtRSDWd0vzOA
RhsvQ2pyW/YQUlJzegX2f3v5W73+b3L3kH+kxXUjJcuLFR+XLOZj7zZytkpGkavC
IziNp7Dgcl9Oft7PtQs23b7p9qwF3+ydbkr+uaRIva7vmj+nrV6CnwYqfJJ3SnxD
sM0IqRUioDczrxihqNCORit+NUFuCZKpUZIo4IUAGyRwssLOfIVex2AX/x2zBmev
y998gCRXsm1K70vSHvYgvvQwC1ixz4yqt+RX2Fm3zMlQ7kVUV/nxawy7OkIVoD8o
SNbvzo/vuJiTzs4psfByUFYjybnXQS8vL6BQbaTmDyumqM9SDMte49G5fhNuaakw
EAoS+CyJGX/mw8u1QDtisu3a4A5UzqeqTBh5Psy6FTawEnc42Exc+SYwEWc8Y7uk
uL1HMn5pbuz+jxcxt/Fxks92bgRAahNAGSXKnGV/Xxr9XSVMJOfmXRdxQOdoIRYr
rZz0Fi4VRIK/Mwek4UUw4onRONcerG9wkN98x4fJLHwrryZZ5wuCBCOy1VYm1Hs+
WHeBiWyFcXUd/YQ4AS9ab5vu3iVJNMY3jFjtjv0Mc/pjO72xdKE6fbv/1XGBACM/
bjfsdGUj5Kjq0fLLbMcgdYk1vNJvlWxoUHsB8QI9Ckv3ZC//D4b3GbRrsHwRcI0I
wbhzBIjYIekHZ7S8c5x569a3IHnbz8RIB6Osqh0/s3N4FYmWo8bi9twUivGk7kuP
qIl6G+dfdyONbzgsPd72Utw1CKvnBK9RxsHYi8DAorWiQHmJOB5ixe2fxD/0+Qq5
yf39CLgjjLHPgITsnFFUvojzzE+91YOqXsTDpRQQcEhV46tTtWHn0KhE3v+Gf6Xi
I2qKGg1fOzKlgKM61ObBN+Iek3kqn0FeOBKaNNvlYnP9p3edh321zLdlbcNxPNCc
DxV31lI8lVM2uWM6m2Sl16Kr9smy/JeWxwn5XuKcqfaIRXiB0ewnvqz1HDUqgHN/
o4TvpckP/4r4vMtAl8p1yjh47QCnTawkb/YW324EbyP6f64izcY94ASMHMHzGFr1
UEft1r8nUY6XaRhB+OHOUY5zgql/lx9exPCjRkTxHjQagv+kU4GJ/FIrWCIc2eKo
lKgeTUDUXBpFrjx2pRVZm0IK1LUyN5zp9l1n952uTM2JC/W16hPC2T+ysWtfKRgK
flFPY5/IJ/7l+qj+4DgFqCV+dk3vaujs2e1uWZsvKkpdys3ztEWdoyXADokMkQsT
tL0rAPORyuhdGXVX/MumrPmD1BoaaLAlNaBPutw9ixF3TU+QjpvcaCu84FH2V78x
N6PB901Id318CjubSGDtrL3ElWczEUW8ygtbr6cDB8/uSYgIYadLXElSwvOtt3BM
ICiHcTzmrWQm07Q0rg9e15EgUex3968eG2OWyba7Royo5d5Mzx+5jE0QRbIKcTYX
T9ytsaWk5eTaEKu1YbzYhj9BZThx0NLdtZOJpPlqWXmZdTzCs+g9yGnu4cIA0cU5
t61lB84eDufteZTxWEQPW7zW06wuc2Fzlf4JYY+y09IsLw62lFP+4PL9y327eNt0
Yl3+mFrKPM2SHCwkOYFXm9wQOYu9euB2J02X0rzNqV/etFjnesn/cPkJnTDgDmQv
RiS6f1gRv91uoY5ApX0xSCKPgwZLCWtbf2ohF/3bWJShlK/gYfvwU78QvuuEuLQr
aR/zr8B6hCbKl5mtAX7EYsZ6MJcVWmkuK3yExNY1eyLExNs3j3wYRbFeZsdTtQBS
5OntC+KarZFD0MjJJJObbxZBmWobXP0Gzv8d4ACAYTDxkWxlu6IquktTBTIo0Ekd
F3cJO4Hrj6J2drGp+IelrVS9zMhP0RugCj1ygKQ4J2/CS/zJ67v/vhE3l222P770
YV2hhyusPOfZStQoZExdWKoJENTq7R0PGQ65yJ7p8XsZZVLaTi60Nekl/8sXPOkw
li+wbX4xRoCEMlXp8HFS36xdiyCpUORZP813sNg3SefO4SQ8pGSZ4LqabnxR3I8d
HKZOAtg8YUO8zI1nebUnb6Ex1vqGAlz32dzXrY2kHPn5R3HjmRcfGENXfYTwgVgD
gWAdoEjGl1byPY6/VMH1m0VrP/NtD9ObYw/lDXddTr7emL7X0S5rKxM3rISF0aw0
pr6ILU9taYHIDFpqeK3B3QMCt2ZneutIahg8MG2ZGM6Icea6Upx7WOsvll1FIYIW
6UQknqboTjWuRTGV1NrKLOllzUl/lrUFpd2iwaZUs0yxhtilHOFD9yzSR8WaPAWa
Ci0Px5HhoFspLZlLRJ6TZ5obitUAXWkcev5svTSBrIa08NvFD2oGzER11QFGlK0C
+tndvDo2vi3rIZUmnTh4FE7K2kAxsjOGaOwt2ILNmqgNo+R7TRwAVs1JwC220um3
Sf/1tIayljTMTeKoAt/n3bf7tWjIu3p+l6/xqln/p0S7Ra2SvR8Z97as7dhi34G1
JJR73mEWdpXZ0aAJbNjxvayXWwWzI9pzDx/qtRGWHYh7fQFSOSrEI41gUtOYp9E2
ifsV7cDqTDMoCrCtmFhoVXWzH+lIA37OVx9e9XCz35EiUoMFUAS9JeTjC7VKCOT8
k+ux6SlwQ5yyZvQt+rGf6SXT3lpEmLW6b3B8j0A+FmnA9BoRcc05YDvnzJSToBJm
GEmKcPCBr0zFmu40Eu/AtlWEOX90DSjYrnjcGKwAGfwuPz/Zv8wrmKcfXoHQfzsq
xDw/Wwpz6LDBJ7LOa13ItuIwvOzbIaGXZCNyxSN3z4HTqgR69pxTCTvD+d0vpGpB
IHIZvthPb++6tKHWgkhcqhcmNY7POKtjMz9SpDQcAl5Dunl/oh9/CmbSObw3Htop
PRtqTOFQ+ngd99ddw5c70nDSlDPDm78f/q/PNy2hX/Osz2nFAWtgZ8XWzZrjX2Fe
KSNBh00AC9glq2+wrcIrJevmlKQOf1Za3mw2og+1PLwISD9S56RsFDnB5h4XUdnq
CUrUEjWquEDTDnud1WP8JduEnvWDavZJQmG3CrWQqWO4ibtHM/eyraezM7j+lVfS
GngJUoC+yPgPEXk6pg75waA+SBefZn8kp4qFwz8yrAAla62Q1NkfkaXYNvi6CgKN
ezCRn96GmpVsX7axxeKYZMhyI4RUH9H0cUY8BcoAslzN/pEOCD3uuIjPw3Oa87zB
+wNt5mi9qx1XH0OjD2PmP1RrCVNSokTOOXvMWniHnrc7Ky9Aapk9jj24dNZBjUrV
aH3Pzc5G08w/6wo9w5xDC2XNAxs++IcJ8Ulrvgtrv52Cev7B0rNbL5/nIRHcoA0W
AK45yc3gvWBIS+q9Lv/yDngd+Rx+/xNtARPsIL7V9fyIp7cP+gZ7bbUBqR3YvSWp
v4aAZT23mKkVSQbE+dw61d5m1c3l7jSpbJSXrVDfOU1p4OGW8WAxckubBHJFhvXR
I0yFjsViDI6a2QzGjojBoXLpSJT4+vPZxcGJukkeU1q5eHarlLE4oWNkRqceXytS
M0Hr+RAiUDJ8BTOzKarM5Lz/ngKfP719QEE9rW7fGWmMgnMzmjSO15zS0qdW/40Q
8gx5N2ywJiUO9lgQWRXTf3HK2xqGziUmHEWWCvcyrd77LIsAAUgoTk0lHNG/lEOD
lUO69htcDtrmEpzP26F+DWIFYIDqbmMW6tBMUxqkWYK2+kRec3hVoAuc4c6aeTsV
X/REi1p/QyNSTV22nl8+rTg6Nvq/Bs881K7EwrWqPSBaWSEwdbK6w9ZDWszjKtCQ
Yh1EP6TTJ58tN0ZPFD5HN4BQ9yX1MWF4GXcObzGT0Pv4xRrKbui66+BZ7m+v+K/L
NyhJwpT6qiW4HXYJVqN5ldDwNManod/EEMA+QYWijh6/haz4EoaPpzetpRKZleKJ
xW5KQv+kflVgZk3BFjtSaomYemPhIAUqy6Fir1/JxGkr/ulpWijgH1QbDCtum2uP
6N+B36bVXPZGgZeicZ8zuqBLRN83qXdQHH4DOi1PiVklMk2RPXyLiqN8MmB+HfcZ
DLVgfqhGdUlqWJUyxhbvd3PsSZoSeUUv+Upt7Jo6P6hNOUBTRyA9o4rXJjiSJdJh
jluuRsvL2s594xmSevW8v69iovMbi2NUC6XV6eK7xdkBx8FZ8WHhR2xPGQQDWpua
2QXJhQf7gvDOKZpMXTz/tHSS9FOAJe4HLLSvVnfPul7CrKzGCC7LFLCKrFVbpaUe
TSLXU0WdT5AEo4rA4uOD/AKbURrrsBzL9DFaon+naVagiJa/Gi0LHSRCM/p7/aBW
eqNRE/VATcsXQj2HU7OvNJY8zCZdWdY9WyWC4qd/H+InKgWp1puYcwxcTRJ0e698
6d8uaw5q0blaiquQXxUx5gATjFvHf8Kid0Qev0B/7szAMZalQXQ5kLfh94t1BwYi
lVlWGGAjERMkRA0OUDag9n+lr0/tZIw7FuqW+MDuaz57A0IXkmjKPR4/BHsDcU7r
oKL+nED/aP1Rebf3h4l6QD76ikY5/8JoEhN8v/PMbkee8N5T1dFV2VwH+3NlB/WM
hxqU8yYJFzDVyBzSMBQBqFhE+g7VoOmQ2I+B81iPC1+iKKYcoCjDtp1/8cKv6GKe
Z4b0ZR+a0pCGVq7pQRmjg5CrZCCMHxWxg1KvQQmOme1+N1fGlFOnx7ACwtigkqLe
Jvd9262SKwVqOfbl6aAbCXiEbALZVDmvl5/EQrFOYoKKXTrCXrMMoAjPchZ6yVB0
Z/hZs3v7RktJldtqhAy9ZXHxaLctAGZMi2nxKafIJiKcI0DTMgfB1v5gFZTjIW5g
pA6goGsco+UNZ3RzdUDzLWWFkvoA5d6ysvmupJhMgUyh5Dl4Tf2St4ohrsLLZJGk
23PG4kTXAZeziXIblaGvstnvjvmiic3UoKKMEQqpZTUAejVJ8tvw2ltFx5E2LVsT
p+7pTk8MgDc2VY7gdWy3MjdoAQ+qp0zm71XEqAxRQPJB729gI5zT2/XfZ5hGh1mF
53sf7u4Qm70fbtJp5bGhZW7FH+eRoeN8D3jkxMQd/a3+nzEW94N/7G7nqaHu9ftS
+n2suYASsSRd2i9pGLn5NnHAHd6Og93LqjNuF/603LvgAecQkYIFS+A4twITlPJx
uqDjygLr32wAU3FkpL0eAijIm0S4MKfoj8uQJA07aCjyK99c/gdyOm00DzGkYtwT
nkDSlCy32rFFyMMIbsvfibZBxVArsAdVELV+CnJ8+O3l+U90t9vXhTMf9HXZVGoC
AGswuVY2K2pq77XcdmnkZztwwE5hYHZFnI4wmWLE36bHZm5TfYHzAaHgfaCA52RP
MCLGA/L3C4mdiMuOXzfFyEd/myUDYT6KRGBV+dY5jJ3eAxsCUH9fxMUFkJpClY3R
QAE7x9L3mvSnDC4sAq/xpt56fzXGSACkjppTQ9uEVz74rj1hvVj15IXuLO4uw5qQ
7NOLRRMdXj/zfVgLFfdtN0tq3eErggpZ88VFSZnBRgSrYl/wVHbicdzUDDsslPvb
rjLYgCNrL6Ysgt5uyO7GgG7nr/PBalMf2LeU1ZHoaw/F1HhozBtcglDIgNOaskT+
HfOTqZcnSbK6LXBgNv0ftxDYH3Uyc1uxmDFrBurdzLkb3WvOwNMMKW2cJZ9vPeHu
as6efnOvaipyDgneurtZ6NOqdJwQ3+qVZgoZbZ+ekoVHzRdUub/1OU/Ao+QLQDyc
Usk2ciWFj+nkMRijIDvWlk98CUfrXTj5mOKgjqOEBjKlMWKOOJ9rYK5bd7ua+qF/
mYmbKsi2ejG6AWQw+ss8q4RdG+bY1ZX3IUSIqYll7wZVMH3Kz5b8aub3v56INNrw
z4eWO1/yerlyve7cLHMXTJJsZdVsgmyTHKjjuADwXNUny0zOZf+SNAgr3Idv+P7w
x/FHeVAu+Nf9MFvENCYTIzHID0vgkpTFtyiRStVrSFovWvIBp5cls2SRuxMjt5s3
YB0dN76gFwENmbZopmNcaq5S9DhQtVUOUEMQnYns+K6HZ+cTDA+o5gFgZD4gTKTI
/0prKtzVyONY8u+kWvx1e45mu2OaLQz64BEmLoRcUWa0hAUv3/b/NYYIAqsWCe8E
ZxeIj41kmsPVEl7NdjabRmsXcIVFJI7QMa83x0dXDASZOCJMFtXxJ8sllKojSgKx
cn0SqPy3ZElbOmt4V3zWTFw9GgTzRVvaJ7ECxj9TQcWzJX3JLW6KkRmD6W0gYBJf
ZYUn5hKvw+NTHbj5/hU/9P3RPnbl/5FSgv+io1WWbbR7pnK2zsoEjlnGgvbj5LYW
WGs5VyBwFdBSyUfF9Hxihv7TCIsCAklNiQ4qIhglF3m2odZn0LRPu3ca6esk2uC7
kk8iiatxDKcpbkyd91Q9UcsRYM1cdU8lQeLKGCPPJygd2wYZI0bSPOZpvx/DAUw9
M8WDRQ7bA32TLy9EbcCk35sPGOfEG+/t1RlB1fkKwChNdQHsEirwSVaDCnPkzok8
+KedKL24kOAMzvDttDt25BlGwrFflSdcG5rIdMkfMBQ6kZNDfjC1PO3zhNE2LCeI
jocKRG2S9D6JczhgPxm6fS4CGmQUsB+4nQRfkA/ku3/3lpE1bfNdxCfJQjTU/47a
Mcl5GfwyMx0W2fWG4alTYyZJLIBx4qKhIgeWiRS7irhdXH0pvaFH42gUaAk2UiGB
MOnVlZLwm1CeRoR2RmqxMWcJ2jZZ1jObxb7fNcNzq8Jmmst9QyRng+DerMpaoCr4
r9t/PreXHJKR/fRHZGfRUD/5ERzpIDSQWrOvTtPI0q206xKSVU7ZyEsGX2Ig88Nl
XidAKnAjtoq9IADDsDUqnWYEP+Uchob7I/1l3JfMukCzrhvtEsbD78sOeLmNHu8s
xYYHyMVYIhH8yaSRVXMw5aXrCFg2fpLdbOk+voeW3uC0BT/vxoxtVuT4tEREFWk8
PDbsuTPNyLfjm6/BNZqofYGSxc30UTZe0w5PzY/sMgqr34E+PtrYKUL5MtIqegZp
hx9jy8hBK3eGcX67CQN0zNa4mGJjuIDUwbNPcHCX0qoib34PKygvyMiEuE2bgzB+
3bAhJUVSEKW2RWWQuTKFHUeEZTc7FaoM7wqbcXZINFsp9SYkmcy0tgX0cZHFyzgp
U6OQ7McrABKkG+FSAdTacijArhT0SjuKt4DoGEnMiZyGsSfOTR+HmAFynauWe8PJ
ZrJTn2A11jnYXXiPp9OwBROqbQ5XWYLMKzJ5GIt+gCOxQTSHcDrxPva/vwCzY7xU
dGfonGvNIyxb3siStZE8GVp6rG/4DS8ExbxiycJokkJse019lqRrGGefbdqurwU+
DLQ5zpAe/3kLyQzqk+lw/xOaP4HupmZAIAFwFwSR4mYv/eDxcPS+kLCp+gJyKEG1
hQHo1TBYgX0grC9LiJIKykuBKCN7Lth99pLE8qmy9YdcBqiECd0MnMjqH73jnPHW
dXexm+oIx5XwQGm1s6vht//cvBos5ebxDwGXnILgDPr2dghLE/ea5QdsM58MqT9W
UIFYp1SduNz10IWUbRubijWfKawp4EiRmsAOyqm+7NJCGrgSBZ1xGVVbUr4ZJtNN
tV8BEtKqsM1NTo4EXJ6S0EU8p1d4NbNcytSFNAenPGZRo52qSY/m50T/fkrsr9E6
Ec66V+q79+ys1nV9rBeIlYI6zD3QqqHDzSvbCo5hG5Clr7Se1NvU8yh7DjDefypP
pd2DEBWe1xMMBOlZ+1bZXCeNq9ACx2d96z9hkRX8NclEegkC4QGaPF/zJTYDmrY0
fpBcNTKU2RVNYVeAW4UNuCWv83KSkukSh6Dt2M/HFJ+7bg3kDx4Kw6LlmZJxSogf
VIACdqdmuSyVM2+iVZSX3IReQuCxtSf+LyEk5pG9nBMJVRWxFQcMrEnoEOZYK8dj
APwHU+vECzrwAJt+yLqaXBABH8NteuH/XEStjwY0xNsAsjFPuUR0elBb9LUBaror
6gn0PVsFgH19dhLbKJV/OGlM/F8MIy9FgLD1uUlXqaeUgwnsbqa4mocsXBkx3QCI
JoNR8TAzHavRTcknkWIwdO8zDK6DF+3nMwP3WOzXo87N/d/fOeptF8V53JDvHL18
Qp/jTpcKsVE3YPJEktNweZ7xQuFIPaqVZaYZjUS0fZc2WCEqJWfA/LFU8Z9/Z4Rw
MNZQjK9jM8m6cSa9qIf103Qt3FZy1cm8I1PLxcg+3ErjJFkjzR9zFmtLreVRHUrK
tvWqQDcG2x7+TfBUg0p3SbyedivDQWg/+qDnz4zyLmbDMZtSaKmAKNMS6xQmYV2R
QmWHh+RY6OfwQloQfuZQvnjRCeiMMj2n/KZXpu4YtjGKBM5ZT/zJ2PEMiHZCYhDo
kXB0FdMapQ6bIo2VO9jbaC5fWJB/ORspNJUJU3h2/nZvraZDhzUq7rgLuqya1E8s
dQx6vw6X9LtSs0pJHjMeVajuTyh/O0do7v9YZePWZjcB7fkAyFdjzXzKCpbNH47o
RRFEhV66VBpQIYkOmp892DL2LxAVSdKtN4xmaS4BftPfH2DK3df9NVwNKgqXv0i3
Bm+Hn60rWLypafW+JzRpSGu+B2hxWA+BNMV/OId/K/GH1J6He2t9wppVdqWLePok
bUIePCLKb8K8jeok3M/NCXzhz0ICYP0/SDjDjVowuNO7j2U2Sx45gcVDYBtW4OuY
Gj2y2viFFL8lINMCkWm/ujBJLo07WJMOTXzUJrVp3eUWY7XWw2cJ8y23iGXyss2U
FCbkgeXLQAyQbQXe7zD6uxZrtrcvrHgvuANU2Q/pXUFVomGkJGJlV+auh59TZHCC
ziu+wUi4Y1iwSEKDVwAhPJhbCHhPjdUHJEH3jJ92uZgiEt9kRImEdPuxllYO2hU/
j+FKKY/lMMyM27LJAa6ITvZ0zmJlodXQDpz+24qyNNoF/clv5Jtk7LTH2BPk1hvZ
oH3pGMpRuhdryWKMmR0sFCAfaRR08CPo1tY1NJLwnjB1LfYGnMGhdLGWrCPNu+93
0+slO6dNbLgk4dbpUCUR/kxALH9Cm+scx+Qw0eEQD74QwFhELHjptGHHCaHqAVt7
44PCFU7fn6rr/KV+mnNRhyVVRvr+LzS9vwKNwvl0FDPJA2OjNCaimN4I5VrAuhJR
HvgJRlTfjNq0yy+Xgp4xzJkyK7zs4mxWlpKe0lqpNdJfAWcWGs0J+XYtS73xxrws
b8GFNz1aZlphCj2DuSEowk7vR92ToHHMqHUoZuEnOYlWu+n8CcAynYmhCNwf2yTY
2QcM8v0kFeRuAwcfyLqGXcRYC+wLgwigF1Nzy8nos9NZT3gp9gLVGJci1EvEGndU
6YkmBna/kcunpzWkbA5xfn+31JVp0D2XSvS6/zup36gm2k1y3cmBZkVDEMucjw/V
Qc86BLND7cjkPYNElCOzsJulKBoF+AtHBLwTXD1FqyzxyifV3d+HPlAp5vZygfbO
Hs61sTCY04PVRO53IIEszQGDjmYNLCrA6CZAvkypVunI6Sfsa+pHdWvzpIy3gEsF
hzFhhbLqllVe2QUrrO56H+sPk65dxcGvsx3obx6WpRi9mi+9etxgtfi6qvRTPbOc
3AI0jpAppJjtpYuKrViUWtLrdghPu30+teAs9HmSMH1kxnpZEAmz0iyLx78xJymc
83Cf+lbJXsYeShUNiNZpq488XdPsQBn1dUA8IN3t3mvy9tdpPAp4BQUdcfzBZnFg
oNs6V5WjT8024nu59dNAw97EYevqm9p1Ed4Og3t0OGUah6F//PN3oECOm02NPqXa
h0NzHNyDNjihjW0dYfOgIq1JFQyTRMWF9r/SQGk+Dy1N/pWDYny4SMOYiAAp1W2J
9UB3bqvnvh14qU+Sxpm9+rNATNb9ox+Ia+L6CT6hxSJ1gn6tftjW304fub83LDH4
NPLbWw5sKAalNKUbgJm9bvAa+98JB9lK7Bd3S8d8dIf2RB2ehGPYFfM6OF4IfQXT
MUKJHbcobJ6xbV+iPYghxedEfvn9cwvoa7JRnricKTGJzcIdckru72LwTT4uUlhR
U7anJVJp3FuICTWf/vnp74XDG/jX9EJbluvQMaMQTQ0IPGiaz6xzyxUFLCnO3shW
mw9zmcy/0DuDocLWATwxuwkfwIINuLF/yhI4Urj9wPXpIq6cDGWQt25w4ZjLo+8s
kmitpeIGWsFgJwedjLBRuw0NVy3zj9tYuOOZ4poN9M2k71hG2XOI+WeGi93vuE7x
mV+g/lZg+4lI8sdgSJHwhyuRL1XMpzK3tzESvURRDTdMEIJNKvKD8RLnO4JCkjGm
zAI2g4HmWks93rVNisUWxcR7iVYJyfBqxXXqOZXHriBQK4CoPlfaAcV6VSir2i99
G9bZGB1Hju0wuaj5G9uAecpdYMdRtcII5mdKm2kUqXHy704K6ibNxLsFy+b+ucZa
EHiWh+rlmGZyMBIkdX2/YJf1xWtwfGqvnM3ez6wvnLKYG2Ig+iqjlcE+bE68DJ86
WVFCpBCBSHDHSKVqBeTCUOo6DuANeqamI6BZfKAg1ipVo55MJsfGIrHxYiQxR4Ga
YiUsoO103Ev/aEG65EXJPVLizvLUTG3QzcXu0EdnaT2rady8/FHdvJxVa9bgasBz
JLqF53k5g0xfyIYs1YIHWBRPfI5++ujWcDgo0xMk+gfZbbdzplOtL1zhk7RqXCWf
CZ4ygWxUH8WB+kqpYlVv1QlyqNGr5Kysp288Gev+/hRLADs0NUKNAaKByVzFdm55
ADUqvdPtFgRZmt2hxSR9jntozX9KvsCnuyd6peixZ+gvZGkDrMytyFgbI6WTPqKl
2HHJ5Loi/PojekcU0WDPGx2GjhetmY6a+9EQ+LDMyzsIn1o/buPdao9FLfXAXld+
h/wCgtBWmGMjfSo+9bv+okIv5jYoVrKNTHsyqRCSlqE+UsA72VlYvwPnIEpk0AbB
Ts/Z2346EBXP6BUne9yLo9sBeVy8HjK0TP1PcHiJXv+5jJMBiSL4OnXd85a/Iiso
GeRbGMZ7Oimp93ft1q5Csnwjoxa2/JXd01bDLiB4+2Xt9fzLOaa1nOLQ/bPGliw/
xZz64Kus+SCAIb38a410DepVDIVtBZKfQhSeTT8Dvy9ijNwulgiwdC+SzeD5pLFc
oIiel/f7utToY0tLNIAwC0G8yUeKj08i1RmqXzPN7zpACG33JUytJV0le6LCBPGT
4g3kVatTMiquNtktysXZkYQeeXgi+r1deySOOTezOZqbPOPO1s17Uo46zO5HjsiR
4Utri+ArWTfZSGt5so0S9FNZs2+o7I9t398nFQkcY9iAqoSXWyjbrRPORADKeAm9
EdBGL+r6ngu7mNZz6alh6uA0Z9a2095n4TZ1slNZLGcdgFKhdisgRru0MSzdoIy+
uR+K4tRIk5pRDhcOwOMOEJOXsIDr5EFzTaZysGUrPMwawA3SPRjNxxCeAVb+S6jh
dkn+nVjPTs/YR8Lcssczq0TjMYX8+1e+dkTvBN+Tj3KaOCQzzhqjX1MC2yCi4XGd
9muC2EssaiLJDLcFiDJo/P65TmjIeSwD325QNvhv/5Bg//kyj1pl1pHzDuwL4Db5
NUOhHA6NvhUM/tGcZJAxv30jE5iSqx4hYm2Ru6ATH1BLmn8PDzU6FkQJVeMAdTpP
92ijXaLWrTBVhOYJuxatMwBj6CkXI3Fmk4FgUl7CMIKvodWKd6GIftXPUbZJz0xy
ThGUF7b2bATUyp+k5AqPZh+t8BvecewZeraeVgWIgFNGFpXfsxvKZ4gmdByJRigd
vNx6ayKpmKwXWlpCuCuMKNg3jeVmfUTvfxRLCxMRC3sJEMFEz9RZsFlQfkPM9wWJ
9jlD5s0WR8V/ad1KWxlKdpBMpMl9grsT13JfPIWvFbk4mCDXCSIjRdTkCAATW45b
No5O16+HvMiIpvOksOu9OFPi6dQs8aG02Z1YHaRbZ4U9ba0gKJBOZDuaTnBBCCI9
eTLlV7kOiEENJHHcJh3ygncEAdo1bECRgL1sVjtgx2y8IpZs3s+zn8VCzCReFGqw
ud0OC2bhh5ZcGsIhOXpBHB7Bm3C+CaL4ucN5jFS8cRqVR8wWT26RdDsmzIK3FTzX
iZ+QRVBEtkuxKVpjTd3WVYES/nncVg0/AEwfaHRMPncn5wSsw3VX2OCyFI5BxVfA
jqHCWDpZ47PEb4BBBlR1F36F8a2CrLfx607WKXyTOZLvXXGf5fe+HtZBgbb5E7vA
lkBJobYAtzC/rnfV+W2wo21vvEOK3D2xWior1VO60sqEV4NBSnV1F2vFw3sqTXKs
7Y6BvRz3Vc8Ui2ymo9jWE6t8Kf1sYoUAvlMWOjQqoQaRKuwrtSHKqml57oi+6dAQ
DHqj9VZFX3G7ThtCVzyvroXq3lGB890zHRmx7YLnhtVMZFwNftxfpU/icFL1HWxl
hnCrg+QkVte4iBylovIHQ8Ip2sVD2YJr88wRh6i5Bmf7sblfqwBCzTYNCvzL/W2j
oMwLHXpFhg7tyVHnmSqyP5C930WcxiYnU3UzBh8FCmKkkagAmW3Cmx04drTJVwVY
3NRAFujRp02f3pmJ92rVmZFO5aqJOm2rx0AatnQF4shYHbh2ZZmvRBJEGbHIXOCq
YpHxKtXSfC0MJIPtUo0GKxRVXseHjmkgu8t4ikQ2nM5KGc+vYnBYgSm8Om8ryqJN
OvWBoWO4i0tX/uU+KSGC2mRBfjh6Ehov2zKndeJ3/T3+TVM2BrG2b5Xa8vVztJMW
SqcJswCLIYXIinFOTk56q+5DIhy7Lo+ctNZJVHuBwSRM0mx/yhY77pdK32B+PNgH
vv78t+ah+7F7EuP/XbO4fitbUmTx+Dma576GSHAkHmcD3Sj83TrQoBM8aiNjRTEr
GFdB1RQJWz1SkiwAR4vPTOVI7FtymOouaBxcri8h3otH3KfSjIAILdtFTRD7cYde
/nrfj1b2vtutQk+Z/8RNfEj5UpmlvIAGpsROLbWjA52sqQA921ZWcg90HotJA/7Q
sym8oIFuPhkUtBvbtkatzRja0k+Dqaxek2LHVC+N/PtS7/+ot9/1n+XLYXxl8Hd9
lDNczBXrWDTwEUBM9dVxzo8Qzptl8Hsb1zIG1AqfC5EMX6fCjoGkeiqOpLj4Ghrz
Wh9t4KoTCAfPmZ5N5MscfMVT1qRU0mmWE7LTtvYUg/m4zkZy/34leZC/xTDUuO6r
iTLos06eV58GuKXCCrPF64e4+iz4gLM4tc1t5iFlk7xLsQ/0HDDyVKheUvfoNXgS
eIBOquFFdLtpVzW9HxVeBe6SbKHPs5hiQYYNMTrUzXqR+Ee1gCPO9oepFbCuHuqx
Odo0HcUcHVqWdW2EFBgum9qfZgbIOBzv0J06HDfnHL8o/f3CIbE0jvZuAd6JnA3D
8WeGpGzdBosVFR4wI4PrL+hmFutHm8oz8xL4WHVblrHphuQIhvBJFjvZu1Sa4i+e
ISALqXSr9mz6Ho99g420TjcjGHI6eWPE0kgifXzCkI1MjyV8mwTgZu79hLcXjZ8b
DHWIuEScBzEJPzeSmqP2f4XIrl1+5doLraUPdLEMBXnQ0uCMCkaPrD7zrLoyQjW7
FkhRqrK759gkBprk55NbdlZiigDCFwuyeJ06vOZ/uAxR49mxnyu5w5zhyVj+Usmw
TvhKnclm7oYEVcS0ddQRPbD5Y3bSU46ds14epg5uyeybXGHBdgHeNvRdKUT+q4V0
QkivlsdmGKCZTGJffUqMLUXfAC+/IEAjuZSNh1cgWGQTta8B7QPpWO9zgYxPcl9i
6ilyFEEJYlM/fSv7rr2Pt184nJ6atagtepRDSoj48VpwikGjt0Q1yeGOeZRSQXv5
E7TStz/ry7/FQbM4sc1JRhxM4jqsVIcH5DAw9YthOvZ535gsLyhK9hVltRjIRG0O
nB506y8l8V048myEe6idTojT6zY6J6H8Os/63+vgnsyx0upqOdFn+J2TVTRIQZ+z
c5ZQBmBNZBvXYgu6k3iAAd69y56rW/I564DB0F28dmEFoF/H8FlkulwEBPVDvL4i
/edJ/lBtRpi9FJf41EqgP1Z4aznzcPkH38ZLkr3yx9ynEw7fYxaDUkvVZWj74sWZ
zvPKpJcNz3dIF2V0ucczjxlcTjlRNmW6pVelSyv542s+b/iCRL5SQnhF5/AyetxM
sNVgkPl+VBst6Wi+jYnHfRsrfFL3Y6fm/wksuaTRNpAzGI+bjEtwknb5Zr3yOFfC
hR/s2QLpxHfOxtl5MuVw8rNDTZkk7z27573ZkHxieCIUl8Qz5yI8MYKjhzRcE7Gu
tKTG1yLLecploo4sDBWlF2FEya/7BruyEUyyXXwbysO+UvPxSn6PBvvwE7jzClRG
PWtL7yZBy0SoyHD05G0DMpCTweY/04XnqToHtEuZxBBhArtoeS02i0eTkc0daORz
Wx1F4ekHLWjL2iJglgFIuBvBtXiWSo6EK6kUwSS/QkVVnCNosdXi0ivcl40Fpesy
uD0fZ6JygbDxbkY/c0Lx8qBv6o9TLarF/j9XcquYZB++Gc8FIY/V/t2O5P9ODD4d
dBeqsuw3fezXoKq3L9cjdYNqKP6ZoGjM/J8o+6+bupojLq1g4j4S1OteEGplPULi
EQIHcHFGU9hA/5I3o+UDIHWBiVCdjIvFG8LHlz+3CZUYQDWKTVsZf8nVM4NcZJFU
RJJCffZt88Azllc0UozzqhYHP6VQX3LZ6j1sIhVz3DnaWb014zJ+oGSnqUE2dsgS
M17ZHtc8Y0+Kw5N/G5zvXVYu2tEyBE9nFg4PosGZGG7ZD2pXruBqhWjedQWMrqrq
wYZ+zSJGB/Dz7UwW0ncSWEBxQQWxJC+/+y6Kuy+ovmlWwolCDv0V1V/iRiTmxq+f
+E2b8GIVW+w0dVh99+8MMD6frKurvpbT3WAOTAW6L1QuFV7KHgMzGrMnIUq1uMjv
oHCcK70PW4N3SOEYBXKQ5xZoFsFYWtHcD2IyhR/5DRMQJ0cdcRi30z3lGLCzPgj4
J1Cqa4h4sD59uoJHkHwsorl/PcyzTpJonAMR2lzAPw1q/+7AL17kYii96Uz5YbYB
Gvv4N90n1EOvEYnZC1b8uY7/EOdko2bFtSjEySb8cSD6waVwZsXHzScMgqmTh3Pb
r6md5E05go36i/lakyw/egYbKYHPu6T9RsCUyYZvBs8BT7PYPs94m4AznPh6KjkQ
3HaIhC1qXaiasSWS1fIp5ibM98oZdFL6lnJtbJCEX1Ni+AX8UMi/PAnsjOtP/Bvc
kGAAJMHHrLgx1ZLvXVLSOije87hMYCApmJFkIf4wnIyZEASAjmCxNAIqgLlPMxhN
GSsv47/RAChhiv84InA3RGYXsTgcj9+YW99PD0yZAZ+5neiTDG+2jNc8Bs8d/RK7
HVClyaKB0GWBZeP+UXkm/W5UYhMidfne/nRM8z5ZU2+zISBeVQRaxOPnT3bRF3Eq
+EvVPQWyX+SZuwvloqQaZac0SB6Ztbh30h8bafBnnEE7dpYUtO+xdmya23XXuMWB
vFXB6BNAbZR1ZcS+NR5HAzml7Cs9rvYplJG09LN99e0+PU+nQSNNmuSWFS3CyO6j
doLIcEjwm5C3qmLJ/Yb3Nip2mg/k/vVPANPkJW1JK+3F4JKV13r5HHEi1D/+tk3q
Snln8rfYMTxv9AjkNcX9OHSjuut7/s+QwFSQQdOCXpiJ1Y+9mdMAAnGK9fnd1eno
2VataUW87k9mYwa58IKNoCkcvyqBMFXQfV0emxCtgDnrM/LIYgXi8G+VDorn67+K
wILNPhQKjMgwCsMgS8Xf5pDCMG54rN3MVUc97S/DiDh0ikdiTB/+ZRvxDXEORvOt
s0UvWj+mxXk4wwPkKtGDJhXvAfTHMPirJ7020dGjTm1uObtBWE/29WofQ2beEt/f
AMq1zuFlI4w0n/efwrMx2oHcPyXUhQVZ2Jb4i8THOFOHKqO6g8EvDis3Xx9+Xuw2
bhByXfIonN4KBPN43aOhtg5Y4tFWurOpMSZn2BdyCMWxEJAm/OEvnUwwZEopxJe9
SLMnHh1PXF88cSZCiYoGNL78+c8uYRpE/ReqxH2dH18nEik2FmuhdBbnnyBSp81v
rRLZre39D1WkFbv8drj0TaEGI9mW55mw0/UjO/ers6aU1dt/dPLEdWm31e5U6iUv
rwa3yAvb1H/1IYS6Q8A5U0WVkrLJDC7btyr/uB0jPS3+p/mOMUoF3XiMGHNGRdjb
2zQMxnnNG8qK2IDHYDkxWQk38mtZmAAwUZuWC/1ES5qGtR7KT5SmWVkJb4aQTogu
kKIHfgu0IDXEBsuCHu/jHM6r44KW7qXTKQeE2DMkaf8vZPyYKdfhVhPkdX7mRgTQ
iM6j723c4CZU61drqK8QosWUVC58TtOIKEEyzsnq5icsLZtCK3mXJR1Q6JLHqMGb
YVgc4jrjx1PgHtYiZUIJv/7L8x0jP7pYUVpCc7NHXuFB2Xg2BeSyr24bAp1RZpQg
Mc1YlqUgvATXncMtXiv3pGd000WNjcfrfLG+nw3wAnwud6Ea0oFUM6YpShBuV3Le
tqaCYZBMzNjaUA01L6S+s6itIEGhGKWgsgZV8ixFMfXxsuBZsX4nNU5XiSLR6dgS
QvCBhKn3vq9UlKVOqNQzRNgoW9HGy1L4nXh9+U0Le8BxeIzcDJh1EPDaL/BFbaYq
ApixVjdUV4PTsTl5wA6YzAcdYaUCESueGZtOdbwi2zTjU0pmidH8S6J6PhhGU+Ky
LEVfWfFAus8NVTSniaXpa2TH12/LfAXzAiy+LKaFCPbvvr7SiEdFp809Qp+sYONs
7EVTLxiI1XW8MqcDSEYrdw8JnifXu+/DXDLz8UZOdS39zu+TV4y+BUMbphZAo2QD
U/gN/IcI0UmMXvj91YDtZzTqnbR/U6AiY9etH2sq9+RKaxCh+pvTf1t9bDkPIVbA
HI5CrFmZshJ2R7XyS9cps1XNLDM9zr3T05D9pCzMmymLpX4WBxXdzlD4qQEpVun3
yR+JrLFGYnTiLbP+lmnE7u6kNy2ydFnR6jnGZ9kmsj/LvVHqb0kmTyLqXsTXpoIT
EfMMSXXLAA5bqz2eyYAc3kWjIPpA5EcojPFQ8dRKVt/zsXplypEFSbuX+FRsv1va
OHJqCsNqxNJ7RV4qvO4+0F3DWP6fhIHT19mqL2tFwZDsW+31xpWYLHSuPhFZP6Gi
him/J2y7T+C/nnxn/FvmCtM55z8DY5i4G1wNC4JDthdsD8uAKQoxx7vCbK4CVg54
S86BvDCST6E7kr8I6S9CVKGPm/a9QTq1bld89KtxpCVE4XNr0zQLRHNb8aWDo4Lv
I+e4Lkf4ahLop1GpNH546r52kz/3Wwe+7NneY0Xi1rtORufqQADnH17aCmlrirA2
YjgZoePNO9po384WydAj3IrxgZFpn3H7OhMb891w50wbxOjGjbNI/zbhZFQNJcDA
YfKH9WKCAqy/gwogG4cRkg1cKzzjPusQVMB1OALS8OilCjo+WuBH2f1OztSSXZUc
MoGoAsvrjeNbqUlIiOgOOAiM48xZmloyck5ZZXI3xb6HGomGFCMIiFHhCRHPKK4T
e6pf1gfa5qbHPX8bMXukUnMBAAfgD4HWvjx801gzQr1l9L+t0EW+fXMieQ8XVKtp
ElKLckUv64/C7KV9eJ9sgX8XUOq6ldAAb7i/O1UnL4LvFxPDx4cip88jOprqhSaQ
AaDnDpiB1BoY1Wt5N/g3M3FjzaxxvhsfCqyTnA2GM0lcWuQrlrXqmUJc+lBxEjFD
J7B6ZZw3TaWuFLQGyTSKENJXFCv2qDNXYk7ULJc/8hl2+aABoFoZdv5eqw1qjijV
61Y4GrsFdPbon8j3/WLSCV6qy86+AVP3+aKyQOYvS7BR2ftRA2SMWJLVR9AbpQMe
NSswyJ6kfqrn5VD6xc2KIxz+6nSqRz9RcbjYgANdMJBsVcUPZ+y+YNGAgkxJ3dhL
QW7Rji0izFkn1C8novX2oPJsKsfuwK9RRS1V5mZAezjjwQUyIk626mYFdImgzG66
0k2lBT5BNy7bK4BzD/iq4Xl9K+xlSq/292svQCAFcVe2Qh2i4nNlTaNrFYn8kge7
7JCfmYNJjJ80PLeeg+RAnIM4sixU2hwPA6wsfCbBkIlMdn8Sq1WIvbO5D1fBwrto
LLJxSns5tTKm0UlIeGHHT4lWO2DZ4jAcNEwOk7sYAoeqMThwu2OcSNrLWlBhyAyN
Om19mwTSTRYHJpmiRg0B59siU2SQ24Qto2wIiMrWuja6GHSda1v0JJcJB1+rj4I+
uey8j56eLW9MWjNS7dRcKVrZuRVksRVe0zpsp4K60q7ERVAL02ZrFVR+4vuf2Qop
jcc6c1YBMr8Xo3joIp+xCiivgVPZMRhzw7ykO36p3MqbesyI/62mCUebOjY/4cKY
09DL54CvPjiL//MmKtfwT2+k0UmayONVfKzoBax4B7oGJazc9jlQCiU2IJgDr3PZ
9LRMeuemQh91QICU767XqLgETRXCdnbTCYZ34Xo+s94Hnt7PD5Yegysg7lE0qKIV
/cjFsYFVnzxAdSuxJHHZX4a032WgD5LbD1FpyLmPQTs02mijD19j+uWpM7N0Wlzv
aEPkP7vKHuG4JzZCnTN/3CwJ3iRIQ2iLvph83rrnx2C1R2y1ynEYe79D2JB07Xw2
/d4P7dMrt6uIjxY+LsMRXo7/+YJyvIohBI2hTAhh0ZF1Vx0lvyG9EAjPyDcizPIl
+kcK1dq80alURV5Y30Qn514PhSBtkrsXdv1E9sYaLjRKRnqhKMpR5A9T6UIcWm4/
i9p5mgqzIQcHnwskrN5vkgx0jzGPwVR/fquNvJg964pJfM3EYoS140xuhJi0z/qP
urb7RnnKfPHydZbhfl2+jj+fle2SfT6QdrSQ3Ztc+UL5WcFZGyCik8KScpRgShQg
elBI7Il0ik3rOvBL56adBPpMBiLZcm2xcjuML7g1EeHBa4OTMr/QuW+R/g2ns9xp
MzOFofx+9omI/FCMikLWDu0/5qCpXfZPMzKqgb1ZmIJ8v2hEEWqvJeea6pVIImIr
TblK3oAvbqxKguCbEFdZ8nUUikdY0v2NOFPcwvHE5ZHY5En0tmmKUwIWh9pI0zWF
GpaYKcqA5+NXpTGh88PI5ybXzNn0KX95FeDvXLoddYcmoGeD/MzWIJEopbiMVOUE
aDVeEgdw5qBQCCstlOrC1vQ8GhF9zGiWzH2W57PY3IDX7tJ7wMv8ATyzZCQeuiNK
EcI5aoCm9FqoR1nQmBdFAVeMM0f2FdffVRlM2bgxlN83dkAtfnGBGgU4mwn6bSQI
OvlT/joCeV6c1lam8iMa9+BHbbamI1snJ3/GtVV8h0CH/tl75wWGJ67tIeKYz6PP
ThThCwYB+qY/QGdZLoMRh+vuVt6f5GYrTTIU4CAa4gT1uOp9wX9bywuFDVX02/IN
ddTEHS0bdfgSUdNl0i0yZ3KroL4Ad/Z5aRyBWnJzyFOWl1k+Fy9EDs4gO6ETXANd
nYWHA5WEXqvNkAtNDzhsFxGnUDT1KOB4wx2QyftSOOLCsF9mrTfl9EzoTBLaZ0BJ
H/DDcJUG/fu/QGl34cVMLFvUgDY3BWs0y1lL+TUylpiLaKm5moP7XM10u2PstG9S
8dC1tGY7audotN1LQrvAO9TPaPtzCosmLQg9iZ3CWdQWIHEdoRdHVotSf8Cy46K3
4eIMl3IV5Wlm/mf1bTFSVmYdt3EZAiyFTjtoaQq6nMJpOq6o/Yo+Mk2K0271Ero1
8QyyVt8a3Sz9B+3o2/3NC6tN/AVBOoxJv00OOqtpjMnzMNRDw4brhKCsMF40t8d1
7jf8v9eZiuior1z7ng3J9GMDCgqbLzNezqF5JaMPfvG6gNO1tA3/INUjxUYQqQNl
Ccm+MymIgwE2hwmYZjGD6sVAY/ssZ/NpEdu4DB5PAz2SoDVl1x9INHwbz0UFs9FV
G/GgRJeteG5vNjNokV5H1hg1mOAH4qmAEjzkOpPBrnjksGrIyhvg7LUYq3YcNQZr
g/WwfUjto5v97xl2XQPR7Ma0kusq/Kl2cpu91F3QdKcO6SuNqvayIvY8bGSo8uyO
YjzoPi1GiDHAkLhpPny0LaaPy3/J59esBTh1QdGWrNop3zccawuAdF6CZp4GZNjS
f3cRuxBG3KTqSKS5I9xFERcpvnmMWV/m/i0wCppvZAfNOg8L7FZLp2S1eWIH94OM
EAhJLVhK6fbHfhlqu6OM5bSvZiOSPrNULb7H8WZcR+uKbTXdlrYLBTOOHoatS0dY
oZa8dk3UjA1HBwZ2/Y7kmKFy2hd8xTj32B7owxHP/qFoM2QRJRvCNL1ubCuo/zEP
ZTWJrOYfG6rZI+xyMTYSCzj/W7Yaa2Czc1p85J+2J4E7kav1ZkM7F5hW0Nw6jvfP
thKU8GIMKC5AdDu6gUOd3rWzVi4zaJnDO5nQd0Ft748At7ey4h80SiUGkJJO4oAC
jiZ0blMIZ+IyLHuelEIy6TNTad9j9KitK/zPV8mzd8PIZhvHCRDNyDI9B2NvE3Qo
0gOHU8NBfxznqFbQD/XnU2OejzQNhTDUlgcqIKJTLPwzLL7DTzgQHSlKrPXAK1ZF
xmPOReJvW3x9XRXWo6bk2al4fzmP6UlqxF+yHd3qNRL0dn0oZrW38RBoVY21GTLo
CFictnG3k7QnFY3NvHrl1JqB/6TajHR84Pr2Yo/961rJz/BlP4vjBbDkUSNwiwPy
7VzAq+fH/vET/7+a1Z7KktFXIvVB0tJaaq+74FPeKgW+/ClHIQs6Vvjh1szHQo5v
pO5pdKzRb83kcbCRxsQZvqTDdhlW6xM2QEJdF8GyMbddmRIUNbZYZRTvi0ODr8l0
foe+vaSYtGLPkdCm5D0EMW9BkarGXcUbtjNsuzFZPIppaAJC7wDZ+hreJYgYWcWf
s+pqRT/oyY4oLpsl+Pk2BPNnVoF3dLKd8J7dRHPBrMh5pa0GHJ2WAAmP2tcbr5ao
zUkclJIFaZE6Z4pLBimXDQx2EmxI7OFtmdrRo372TibmbSH8zqYffl8i6K7sHT6F
0u3MVcTrfHoonA8baEwEUg0QTac0PgRv2PdBqjYGmX+FPKy1r9Y/nzRjqtIRYmla
QVchdUSE3c0q3lh1hmkdtUP6KvSzQBR4xbfOxmDCXtGUhE5CH+pqzoFVgDx++bu9
OwPyj4vCbRXO3wLm+d256ndyFIxdIndiNUNBWRJ7qDUc9eCXh3ndbLZTjNcHqdVv
QdlZ2uvQEwwQlkrKV7jL4FsIsFX8oEgdSIGobD67vXc3AboCvUvhY0qbFNkefLB/
eaczrO5yBTqk4U+BgzaEJCpq5blZ9SC3ROGTSA+8e+eZbI4XApqrGtiY73MYbiio
lMY0oPLcGvewnWaRXmlqk8uEzk0H1FKSRIz63oPNUZOUawlv/tMUINj9nn0qpGzn
SGRqN+RQgZX1z7agZ11NU9FRew0GlbngAWHqmHbqwng2q2GxLaELsAmtrjfB+sn/
oFMVFRpQ8SL6e0E/DNxQ/NU5o/ztUN33/dkQZr/fC7aJ1zdUqkJATh7fKOXKHm4X
P/RRDCrkq3SMDTgVKiNXu0niMT8Se8yrEkMjPMcxfSCWDZEXiTChxjADEocw0sp5
q3T3NMrYFlBGLEX/6YqkPJPoxVgJw6y4VVmH+GGW4EZekpS+4Xwe70Y3wXhadsu3
+S3yer4KZt7ZSSqk0Jnj6Ln9E4r4/OvmYLsfYM3S9KD5cF7g+Ff5T/et9tv6E3Wc
ZquO7Zn3SYxqNKI5e01RC9chXUuPnNTuVwL7YgsRoE9yNXHlf5CDxzu9jU1mTHdr
LTTQSkdWoFDURVLFm915ZyFCPPtjZcpbnZMd5HPHX9XTfWj0Oc8ZYWEuAPPUHjIQ
PPiHtO+uLqpj5AWtyhlevEwaDSpTKYe3nKyNwQ2FUgJnO3kBX+kDjxkYq+2qmphx
fy384YFaMYKZjMlmYnCKOOUCNCKMH/mnHI7nE0115WoiZdxJjg3Jo/Z9nkI731s4
Ty4wJi7giSivrR7yLTJwB8zfYlyJxV1qawVCaCkYzv4cwVbJmdweg6vZnxqcWgfu
CGF3nNsKV7QG/AzPwvrpelTnN6blhqzm2KqXEDCAdCITBGSOW3wvIm7gUashVN2P
10IKiVDt3YT4fGvhy5qt7RJ58W0OsMeVn5JaY0jZ1cNDuCalhJ7+PA37bIOP2cil
NlyzeBN+oOJzPluU652ZjyKPhUy4m0Yk4zRQMsGBLLoDuNLHYeDr1s5G0pq18pRn
EJGgronNp0sUzixv9n8TVZjXDERa6k432pqkiNRBwi8RF6xw58VPho1Ikmk6mkqj
CtUExzmxvKytqwKnt00GzxNj7xBXk6oEcCSMVYwqNBqPlJQZ8IJI0UctuOo4iC9Q
51Q6lfA/MeZUCv0O+keW5lULYC/Qo3sc4eOJeLMmTJmAoAJXzpCtWnU4olUEsar6
yquKOjLp0MT/5GhI88fJioOqOCHtBByPKpTaRMcA23UrJ2IS0qCfYtfPgWM3lBX4
rlYQEjTwUqbNTEAhuAP3ezapWoeIl+Laq966FEgTuPcDBhUCv9wHLhrZcw5ATlut
FrLAN/DcF+B0hBbTAhehCO6lWR4pRiMg/eS0D7lATQj2ajsywPXMt+14CPZ8c457
y3YmxZk4poMoouBZvtMGhX758XSWvA61WHkMRbd/3NESEQNMz/9u4BXW/M+ixydG
o1sv5pL2OTYygS+VvjpwmdH67DmFfhTVH2xYcxFCVim7FwNE8Ko4RYoDrjE6lMMH
0FJleUrlb4rtAEnKHQKSbuTyYLK+tjQP34yobjHo6qifBlnVZj1Avo5p/uUba28Y
5fclKJsrhlOtBdsaE5A84uOrEMu9M3nmBCAlSOYKDFxOMsEtSgLlpHQTqgmCgsKT
ViNKfVGTJtrL4Ii/vkqzfMeckO1OMfxEMQgOd04C5cAtrOYo9A8H22LjBM6xpfWx
PGG8vpIwApc7R1r+ULf12LeWKsaHVOKgnhTjcKv7WDVte6GsIl9cSCp20nA+otqB
DNtgxzC8AxePh3nM3/hVSBYk/bsG8bhZlC+GiWYra0pslrfMMbLLe1bvDfpSXroK
yTwfv5FUNnL1yAUJtjir5JHyp9P7YsYHZYSU3e9cDKxIymk52H732K3keKkebczD
AxLnMDwBzcgrWGHNoeLhdl1c+3QwkhMflGHHJZT8c5UTASlCgXh1qw4owflyK8Ay
aYKRrwHG4/cD1jWiVZTWhlmWVOerjf09y/hqorkXPeqSuuOZBCrTa3RldeHzAyk/
7LbxoYZP/KYwv6bVecRR+E7mrdcRiuyPNvqsK8zVqcgb4O68sVH0YnCYf2T+nS2k
tR1sUdHUta0gfmKAXnwjBKImkVRp0UgIU4pw/hpWBAiWOypDPI7upKT2agurc2bq
JWDt9NgwXP1LPtNC6H1oFAb7xOPYHMgn9Wko58dqk6Oqf87vS+/06w9N1DYd5qxc
FimdpekhhrcjHFG8Jb3JXjcR2Ng2HOBNi4m1MAJAVn78DEnHimfe366N8A5pPuNL
hHHtvglMnNkfinQmoNEg8oztMJZHpGRNYT2FMF2qKgjNvUrZxQv8NWHzNMp1FNho
CdzYY65yZFWTLNzH3nrJ3E8/dSWj67mTB0c+wqqsZU57B0HLut1PSdfwyFxGyBGM
ntDigYO17/VxhkLJ2VR9wG3Xo0+hMUTmPnbIxAl5y3b4KRD4w8eAfCJrIhWa3A/l
Ve8r/x1qfpATSIT8H9E2woDmFXyJJpSd1j932Kobt6qP14eXDW7iiNwMZp4Mgr78
dWxgxWbg+wxpIaaJOrPcT1AegtYcp+IfVP6l93Ad1sWz5tCzwl7CTS8wEHKJ+s2O
5ryfvYlnT91KMakEZWSG407XEVxx3sETgWygGUoMnAuysA/IPpPTkWxzz6NqQeDT
Cq9Nw/sWKzV4PpOz0cV9J7y+dsuoEw+srqZ/Cf6XZlRJIa7rTI0oAgXXgEjOVu3o
w/cM7/mYre1VlCXuGprd/LbqyXGZZ09h3KUhzmEa28ibOzngWvCy1bGtsMBUjwR+
+G3AHQMe175XgArQZyJvXTPR0eflWYPK941OoUAPiz+YZpLydGCPs6F279AgFaWM
eql/rr7YmTqq2wpGddQc5cgRxkMbFqu6JWrSF+5cBJyQGmTTSyNwgIosiEb4udp1
/mKf15O0oqniVmZxMFHbmxUgpuP7272/jsnholeMS0lMvpl4IaMb9UmRFgiZseHE
qlIAaC9cBu6GIlyJ6LwpWXWwtH/zhDR6ExkLS/gjHTrFuDL8amq0MoTflM5FCh1W
eM4HO9PhO4C/GGdTSbt5wzI//XAFGxMM1ETU93nEPsYNNo4Ld2ybhEtMIB6tr84B
ny6fvfpYctnMYkHlCluMuDfP4mY/5r338r2brqqqnRZKXpxH6AqZiD6xGpTiBqrj
eQ8GXoyblM/HIHIK9cRvsa7aD91BM3Bqgx9Nlzcr70+f6HgLVWG8xTw+QBbR7CUq
sgp+go82RzY8pJx3rhqZjGP1z35MuPFW9mPmdtgXfqQWz8y+JIEFTE7uEi/KGkVR
7CII8VnUbhK3E0kxJEwhdov+jvXFu2orY5OYpplAWtljQCykOMi+hZSlhFqlw3L0
+gEBMkbv1ml1nTnggif7vi72MuGRJbPn8ZmccDGdCxVX9tMVQ/h1O2ZoSJefOw8v
S3x1c0KxQ/NqIsk3K7LoRWT+Oy3P548Lfuwuje4D0ZUvR2dDdJ+Fvcptk72bA77v
2dlXUdTdB3EDith9vkRiW8pZO21S+TFCoZgoPaksuihJpou+qFB0Xu4YhCTiMvDc
YSKaCQzmQkwYR6nCp/WNytg/lqXPDsoVg+cjaxk4fb5wj5koyDD0uO7iTrZtQ3i5
9TW4w84a6lbeHUbuoSCnKdy2N6cZHpuT6qLFS7lCUg94qivxnNgsLCsn6GsdzVy6
erBpAWN7CN2VY5SsNrShwojZOknVgg8lRUQN13uXAZ27fRJeoByWcY7mqnqttCLy
lTfOVKrh+QwVxH0YyQWs0YrcM4sl28Ha0FF1txJl4yUVeyIUqD3n+I5oagDpFzty
RUj7wCZf/K0Yg6icZz4a6yZVWssyQIYaW+fe+DSSDwaap8ZXMA9/WC8mD7s3uadL
2mKbOD0xH6Uk4VoV4FXlbhcru5v7viyVrb6bHF8qdh18uwm02BLnUIvM6MWertID
VplAItk5YpmfN0SHGVrz5x3tluiezCiqfkvEhiohI6hqk7qQWuhNUUU1TwYotzIi
112BIIjEDHdnmKQhTG7KoXQhxajjyIIbxUp+Fp0GCzhbXodzOr+PRhk7ETK5ODt+
m7iEzBwb9B86CI01Y4207thw6c6GbpaJOfA8UTmh1NaPbm7pukLVZChrrDG5IQGk
gOy6yK2NkCL0lxeH0VyrQGApPif8aIQsQoCCB9aJvuZNwnOberZUe+QvcHYuMSK5
jVnov+iPzW011WyGb/eUP5yIeXQSVNgZgH/NEzx35H9u/Md4kOHc+kdtSpF1amRe
tK8mDbFhWaYNhPfC7ZITn6vZBwYf6ZyaJGP0LuIkmIjACxoKbAYpfxs8j4KRppIY
ROKEeEc17A2fJBT7DwJMXiLEpEfZsK8s2ywp0DZeOapet4eXp3yoNTFr06bxBvit
9arjuTRBrVaSZ2V72za3p0HhGXXswu7mWMQTttXDtEO4w0/2sX55/h8DiYlRCnld
3yJVJxEHIsOCO3emSFmRQUCHV/J0ncVyBHdPnR2UQIzrCXGW4Mf+unBrWkFNuCn/
+/S3JsPEbx/0yHv5LoAres63t15vDmYsdJeu5ATuKPJLKAN9xE4e2laDhx4choVV
wlUFMJmist0chAEJTwoUqb/rUi4Nga3mE+EDmf6kKQD3Gq+9/xPMXNF2KaURYWZd
t2LHfK1FuP+P5qhtBiN28k8Nn4/l6jlB27cAVqIaC8UasrLyaUnO/2iZx0a0m7Cq
IKOCPN8S7cwGWgd5EoBkr30j94+x0RFyqNcLww9+QmEcaqbHmILEY39MevduFuXy
r0CO0uRW5TLBhGiiA84CVz2C7JGIi06WuE0jVtImINhJCI9qYOE+sRYPDourQnr1
0rF/AOUcM21nwOIUGRr2O7aAcovd2pURJyK9dVpEo5VgnmkAli8yUBNsNePqze+z
9nEzN2Ei3wQP9hMyEhYtWhI5p/gBvdX0V+Yp6O6eGKj6bSNH7Ks5jUdXA1vLGCym
OOQH0XIUdezswlgaC3D5FlA1ueeBN0bxVS4RALIquMpvllxv/VmKA+Fpb7sPpQyY
L3wUvxbeoJ9JbLTBE4HgC4oDw+usDpo76fXf1IZB6k9Um7A2eUgO+4sEtHA7+2sT
Z9uivt1L0XqI7Q2EStE3Qd5JlAThDHdOK8VEXERMqjZU7iey7B3pEqyJf/+YQAv2
cyR2XkIl3sgUYMDQRtq8eHw3c6QO1FspgavNSGWBFGEi0XVb1U4MqkSo1jqn3/2L
KasbfhwPXvclHCeSHnWepVVYZFrkpy0qO4z4KgSBDmoU9b/4pu+xRl29d/TCeYR2
2J234V76CbsrDjoW/xc/aanhacF945o6raCtuC3qC1UuNwnkQC9Xy1l+LdG6EPHI
r/x6DPctjPTmk2EJUm9Y3LVBQAYjhoYziUUPLotMzNrmQ/R43oB9n8KAhIUn98h6
y+8zWYFxsarAAa/Nf2vv1InLaHxT3VKCpaHDhkQ7eNC0BNLN68N+XslgOCX25R85
42IV5qy3NvIGGI90DQesJKESoYdpiIAYeOSjNMoIdEm3VWfhjfTUIVVAlDmfxgj+
2AbZsF/qrWE/BE3YHZ/ZAijkLrqDiKNohpjj5cNjEPhEcIlJotBqMmZw0fzzqTKD
T9eFg5hGLLnA4EaLMIB9YiZ/3tqJDdtCOqfGuitd597K/3+QB7CQmRrwOL/NuDC4
devk7mxhkG+79AR1R4z9AsAQUXiqUskkjYZs0yXgAJEXFj14R8n8ZeWDR4RDulhK
WNpT0X29+BrnVVGPmKrZP+7OYfuLDq47KMPAnYH2SFFy8nm0x5nqTOxYQgnM4PrR
yOyG+up4A2Y3Dm8GVi1fFoRU9nTxpjDss53s8tR84Kt8U7nO4YG0E35dFZ0Ygosb
Tetr55Q7Jc4kXDx1pjm5e3UYMH6cTnu3jJZLUT1TthN9lzq6Suy94QpHjHh/AHAU
FqIot9j56tjKRSnb1uPGqGwgs7NSmOM4hKydnyA74/KQS9mrxvGLl3aFZ+vM102V
J4w3RHcHOK+twWEFfE4QshfDpla8IDUP0Gp8vrSJZuVNgNAGfnJyD0BwjmFYmXd1
NWmaeRJrtCfEgXVcPpzF970iioftfvADMdnAKS6Ikc75lQmCQ5w3kgM/6cqHscgx
uVTcKCeZ7HY4FLwxaSBiXt2+gssiBLSK0Tq4En/G5xEbPq3IXKlEL1xMVMysRCOU
wi0Bcv6U2SPsFldmtSqqegs4IAyU/ABzfHnNx6DtTJAI4Uy/fjjuFjIPgMsLVBtq
fENO6Qup8NCSff17Yx/9sglQ6Ei7d8zMcadk2nvAFatQ2oPGQZttdwVPQvGV1N0D
8QMj680hosasJp5rzYspdZdZXWYkKF6JwcK/FDnPPiUhQrk0AWgJB1zg18pSbWqn
y1H7lHy/AJbtKZWwiQcXQEYD/2hCgBMqmF0sWwfUqm9bBEREru6yNeauzg+sqcHA
xu3BNrAe0Ai/yVDV/cNqqTtgCpFFxGEB7CN2V4AwcqJs3IeF+peHUep3uKt6nApR
sU95jqcvTTSixMbsze2iM4p5KudTsrdr/jwQ6CWT0g4Bw5/0Dj+4KVcNAcI2R89m
Q0WBZd0GdcPoAzPSweLKOKX9Or/dd442JhlWM87VpYS9j/TrNFrfTiza8GdXD2FD
MWSHKSOD9Jc6jSDTS/2+F+l9bVOj1I66L8oWx3UbGLhLtbTQPdfWjKsu8QZoY2xH
krHNjbwZwznzaIhjBb/3LgBgWnH4UOVVOWOjXtaMTTExpsa9C0a5YjCXDrrX4N/R
GUdlRiNoTmc/v9gz4VNiBAPZMByiAUeCQ2ZuZGCXAwzCsAYfJhIjrW1//lrI4CAk
YbStQCow9D6mBtl3Ww20qL41yGcv6KGdxyCiJ4OwabgGngHb1wqSrLcXCkm6PGjg
uje9wnivOq4I+cdL2pFVupthjdWBjthjUqfLxv+ZuKoIqqFeZ/WggBk3YA9k7Is2
B1ujqWto3iHxAEJZpzPZoZkLPdkC+YaKjOZ3Nn+5cDxGa2jpa4xDa1BO9r+7cicU
vmte4g7ycGNdTuevb43qpf7JVBJ7F1HVLWiZuiYf6ZRIdeiJ7Nat0DzlDSL2cnlH
bDIos7IsHQTASpdnIK9TJy5W6wc5ipcQM1SJdsn03Nlz8UJvwIvCC55dIJoCfg3k
98gqaco5HGUByQlGG/c4WqnK4ldcyk1ayr+V2kCY1Qg9Wz2ABhRPfrTHjNtpnDk/
ncN6+z0sjg1O8LNvjzMDdNGz02W3mDHMF/yoD5RFfp5uwuBrXl41eR1vklOWXmxh
rqxKoCSzz2UGvTYOP5SxT8VShyHmKO1IdC/B/OkUz3tcGVWPOBWqzpi42ddptkOB
h18XHI315c9vBN90J/TbMof6DhF4wctIuD65wkawMPrYppoc1qbK7hkPWQ3wSHxN
davEjKWUiOb5JoKyYTthX8NQIUyIPcdAaDEq+Lu+3oY6pqcgpv2LGzgot2QqHtcz
seZhsAdfLs1IUiZhcwGzDybzxt2G//YjHEvOJ46/y3MXaGKgRL6zockpBXtDP6bt
PC4AAvo6Urhv2oY035vc5fsKSGmQhsa0WJ/pCTuXZ0x2OwnoTu97hm3+3eoWsnVO
rc3MeGQi8t4aVUFkFFewLaEsy6l0+zQeMQw91bo0ujzXzqdTVu1qNh0iWiXnoKFp
oeKDvGK8x0XZ9Uw1dM8bfR80MLuMhW7kF5lIIRaYJ8vwjaMOyxzN1a5/VzLI3DEp
Mhvv6BK+vb87E/G7kH9BzRQnW6aOq6QfHGDjPsM/ItUzi26RAh6axr+pvr2GFsQC
dYFL+bBkkONxfhpJo7Yv59hhqw1EAUKq2z6JQDI3QM0b07AALSdT27Orux3DQwd2
2Y3V7xxCh++4bdHwyWRJT6sJb7B5VzU6+5cwd7x5NRN6ZA0rx4xrjMS5GFQ1BnIb
qIPQHA7cXG5/AM56Uphbj7/OnEyaw0K2uzU8LPdw0chhyLhaMMDgvj1GoDYURtKz
cowMIkQ9Era68RihYiYTTWqoJO+NeH2EIcLEDgPw4ZF5nU05ZEv5YnudPRy/nWf/
izUTKSJl9P8jN4ke9gpnYJNUcNMP85a7AO16onF+PzkAljJ4C9MI/E29QQM0f2+O
gFSDPOmqaIYp1CVplPj5u0DLLJx1Ahy8A5TRqKrXP/fJsYgFFXh6F0jgnEsJ3jme
oOauf0aXvsgju5/IlONuUWu22goyYsoYcJ7QU8xwU+a9ARIX3dH7VUNvdjSxSPp4
Ke/hLmk/INtJPdzK/c8M7zZ5XTNjJiSq85FnTpmdDaCgfd9LZkKoAUeSPLLk+ouH
KNsQLFSH7PmdO9WDJNy0MnzXVoys3hl7j6k48vPHvnKLq/q/QsbdF1Cz6sbCO6fx
5IOx7/ONJOHHoagTSfcsNFu3KaQpKTY/FZ34bU7mqL9o4IKZmruYwq5SN8wtVg9E
pL6+GgqEL5VneNKPvj78UHvsIDAAjN9VGOE2uKR9u6kTfX2PgRYCio4aPLaC8Xrm
Y2AeXHfBg2raoaaXy6SdEmmxXiy5KhWt0ClQDINMoQ06v84lgyyYiNXqXlZyaax3
wb+UaHx/RMIkXbjNCnpUXvEC/QVdmYHXLgivdiKwUmcZBjME3FiLOtJDpJAdL2BE
1criGS7vS0v2gAxxIrcGdm1lz87cJ6f0Dm8+vsPJKIS5HPVuf8WSom655eFC7sBG
NgRDClKzaJkkET97/lYV2VGYePAGR4EoRX3VNpe/mOkJv75v/S7ysHOT7kHp7er6
VOd3ylkmQ1H4rdJn439BCMnkNfsn/yAI5igTDS8rdiNTcWcNfC0dFuY8P1x8v/jz
9OmYSZlWJuhsDgjJbH/3zeEr3LXN9Mknoev7aHlgiByCkqXh0iGLOn9TqOMO+Fio
wG0eALjJarvHE4wckKnowHnJfIVPPGZ59VeGbW5dL0aEiaPTgkeAYk6Mf5dwKwO2
o+AWNuCYhJ+XMS0S0lxMrCgzB6sYO3e9uyiNs2ZJRXE5ePrYnCJBEjCYJ8ZTSu+W
f1vfT4JMJ7AZJfSVdmVseCFFKr+GRib5LfLGVgEVGd6JaDY9t9cjTWa25hXzx3+I
0VbQEq0+MAJk1ZH7wwShlwcHtTRlQoN5UqzCrfUH43PYDjKr6+0YdfP0hYm3O5Mp
aYl5gsUnYJiPhJTm9CFbtVih1/JvvtxnwuHKoAXMtqagn/tops/OBP/E6hRgZUfV
PugpzRNpMY+j5JkkkhoEUjuKGop8m8Do9nRZEK1wZJLUpjQPgsU4eXUYH65kqmEe
xjRRPJf03jJg8ZUqC/BgVOxTUQBASgpToZpq9xwYAH3WjOR0Bhlr0HpKo7tm7Urb
RjpfWg2DaVE0Otvc2rOICArWWcLkUocag3DxwzNVKpHciiEHFf1FGGK/4zYystH9
Z4cHnZwx+JlqdnlPpovm1sinu/M95KMeTsbCyCkFlpnbudCslJE0Qdc3MfD5vv5h
IGOal34DVcCTtoeANa3nxM9jNY5leUr9scCD8udmc662wv/r0Yz4y6H+Lb6v3cyr
bItTCmi/n2O3Jdkpf4EKluRfDmG5Jf9JEPavI2Y7juMR0eXY3i95r7PfkNz3kanU
8rd9XlQPAU7uS2CREa7Yp/9CGH39t3Rbn72wJ+ecoZflOgQoEnkhvQO3LCq34FBq
CQk5fS5SQVOdA9vqSkVL3rHm3OZ/2jTFyPhcWWT1ENgKt0g3PZ3zi7Iuh2RMS0c3
psHn3lPpx/npbU8uc92e131d8Kd0hvxuWnhvXF1FyiIb24mcGQQNxMrwSZ/BiCqk
cMWIIsaAw0jb0w/rcjGI21nDXGXWK84k76gfnHJxxuaGmt5MmlXqS61hz7fZ6m2e
kYTV5IG5D2GiAQyHSYHq/Kyb+uSAZFqH+NlEWJNmTKhW1gO17in/y9idwLcp2tTi
zGO2AbWjMBT6ge6KkboVpQ/J7m7lZrYhdFYKqu/gTYQdR2i/Qpa8sGXuOX+mfZlE
0dkt0VhO9MSInSzIYQfoVo25Sx/wOzu1rDrFnnln7TkCHaEmP9xS/kCSywnvPsxH
bLz0yssp93/qcbZrD46MGQvXsafWrX986XOd25sbHioD9KIVr2kj3fVe/LexLsdR
E307i9Yj34IVeaGeGO10hOIDHdo0A9vs6hU+zQkODd6WcCXAqenO8Ju/t5vdNGBK
7/vZMl4zeO9AwC839JUIyD1R9ohPWFFSKsZW0Qr5q/ai1c5AXnUpUEWil6BqB/4/
ohW+eqyVOrOaVUWbuWywSnZNwXD4jhvDlTWF0fjRGzaNZxD6iRHvwaeQjAaKWDnF
tnyWLXwMhBnJt/AMGSnPW1SYht8Gbyd5EVMQJjqCH9tFN5XyLG6NJwJ+1Cj71Z/V
ImsZIb1I1bHC742U2MhynsIh1RBtsOE9tihBivMwpCskraTMqvaSLvSHDZZRO+zA
dHJPtSAzzMx26jBOI0TG0Jb9MpSRxd83PMFw0G1tFYVEUZ8NuKsuFAT6lvOe+IlO
VJCA6W/ZTQURH8F97B3Tz+RNkrqz9j9JaU+oGwk54ZP3GfdBUQhjjczbCuP50yll
W7fX5XRIDKIkVXHbhK40qMgzi29HtgDWZ4B61+j9BIvkA311LQHJOMuUecAvMeIt
MdMzGFrD9h/Fmp5eio47a6vicaNsHIykwPSnB/tPiN8PwE9IrEpFZ5wcd5vMYHAh
sQtMPYM4HSr37HzKeCytA9zpg/Nmp952eKb1Rt9+nAOg34ah6c4OnulXa+Bh5THC
nvPyyvvDPXWEYCRUKBCSP4Y/MRofz9N5YPkZdrrTTloPziKIsWKL9Ax75UHLGcPm
X8BndY/C9HgpqFW7YWUgJZEkSST9LcL9rPmWVKCqDWfBZbzhIO9ifWb08O6iSaRo
6jO0ZpjXo8/2fCh9DNNx4O4SzGXDV2rZRCZW9AwGJoCTh7o61s8VrK+dyuo8yBA/
tOZE0jDPPFcGsHzBjyrsqcPiPs/QoKshc+H4btVPf/30Dy+F0xkjF1AZjEw9kBHh
5vdUtDvn8meOhjjMh3GtT9zZZW2R45H5Mu04CW2JtC+axEdEfYXxrKOpyPHIQ1KB
tIYrzzpc0UCC0UVNI4ERqCzoXsa4lsj3YpJ5TCSp+eNDHV8JO6XkEkvObtEDQNYe
I85ugcbEXkYDO7x4oDiSknwEJmo77iSBrgLzw1r6+TuAzJtz0OvrERVQ5gSR0KKE
BZrGsTS7lK055Ddrt+ZX3ZwnHwJtqmH5aFsX+ZczICLxivqgGO/GyoheY7DBDix5
ZcOmTdN3DlS7GelhqsV/UEnpFFQ401zMPY9CgIXRunUMphar6JqgBSLVEJctlS4k
r50NLnrfN3t7nluXbe8qDr2G47lUXouvO/3X8R6WqIEujhReGrFSpfBqtho1Nqtr
vvJEwoohwW9WVkuQ0AVr9/CjtbBxlVDy8ZiRrvrOJurd7S9IRjB5jGg645n3llT0
yEHCTWKu5bfCHAU9e07ccod/XY16A6mjmmpI6V5W+tAEVN29iOvu84KEfhKKFWQU
q1aJjNROAht/TVBXiGTyvh7lp47HULctQngpxi2qzckmBpgTOPq1W5a47C+mrIVm
Cbih9BXZPsgjVrvhHYhMIh/6in4egetEn3oTsKgBldKcTJ0z2Y+pH0EG3sNV5O/q
fSCYuPW7ltllEewc86msxlPP/V2xBP465SWEB7gW7t1OCIr8lBFSS3igZv+MD5wO
pZuOaE857tIv9QDaOdXqb2cTEVWudTShQAUEa/7TU5OhYx8G4Hfm8bX1Wxui+eKc
ceDZvE3Kgqv+QMy33YbWBFl6RNh4qG9eh+sLjY7J/PV6i+/aZFwXI32D8NJ5xzeR
bdvrBz6HtVEfhIBtFDKp6GYFRicMFpmzm2X5NvBSK6PaPj2DxyWvyrvBJxRhr8wB
sB7fhTbmrIextHybt2k0An+GOxOY+NvZULGlgmpqx2zHqzQB/bEOTunDtjxop6Hg
WUr/WXDqyO/87AMc/uKvuc9ucZzlnlckfoAvvA9YHu03CQYiGhz3rtVC8Fs0hbDc
godut96/B3NB82K/j9Q04uAaC8go+sup12TybMO1auNQuhqXPcdNDVDV1G5xWTkX
3u6t45878MiKpmS06p7qacrr+sXB73dqBeT8GVQjHIDT10f40MEzlNVOF23kUA3Z
QsRoG8pcKpcOr54yf8bcg3FcsSW2Ub21/0Tchz1unBqeQboEe5xjpsy00uKiws2q
eMufI+b2krMBOfdhtDV8KpLhdl3SSnvXA3GZyMOeNy2mutfnD2ZW6l3HlH8XZnz+
iqeVtwOtkDXgk+0yChzdex/C4tsJyzeBpxthqD3WQavuuAfiqDksCrIaN/JCGZGp
Mg35oAG6YAzBXgTov3oyiPAFFdcX8SeRJK9nwLmEIsiTXtNIaumegmaHPrtaGc1O
DjCNekrwCOPsU3hSsBA4ViL3Pblanvyi9Nb/WIUbMizL0UTTORHwDwTn4AZOv7vP
YT6wwMlfG6EYXnckhCJ8P4MtgCQU/Pzk2nREWOdDCkFbCCbWQNeHcVM/TyHG6Bhh
m863DFG7+AkGZfjwZ0z2SLuUOf6FFw/ozBqOmW50cWHwcMIKR3Vg2N2DZ5vGvZaM
+7HHXLJgDZMJr0tF2znT9uwAfYgE6LjVCelGnN2GO38EL5lBEQa82SwLkHi4moNR
gMain6Ikcj6kcC+BbiwHQAdTysrBFsPTReQbNNa7oAzKrYCqaGGrM5cxhkRj/1fT
AhGouVhNSVxkmJ3BNxnNZ+K5Wf+iMEcdOA5jHkiKeTLDKdyqlf6xec3O5Aed6fcw
ebmeEu6UXAuFeIwHA0Ak+QCD/On+PVNjSKpLS2Un8PBQ+lRjwFpiKQUa9L03WLLg
KpiFIHqx1l/JdX5eTHQ9vYemYAAWcxtwo+o+QFv2CNX5kqIbde5dAeEMQDu2SSla
wb2RhRDPDzy+36uL3UlsJJj71nlSz2auw+/NOVOW7Q8e4P7r7d3Yv0hwN58FT+DW
0qrvH+wj3VpFzwVuA/CEPPyx1b52Z/SNxRvCtA3gfidinQHt3+Xs6QPa3h73HF41
CZpt6pOb5Xre26jKRzLAcqtwj6fzAh+y1FvWDnqQJDUOZl9xVajL5K6jkLxCYcEO
bbmOQWwsQV8abPmVGPO/4p2nMnPajrHF3Uh5YYpfsGrWHB1OwOayEMIaP3wKlH8h
Njggm7U/6/k0erEhZgVceC4YdboPMiqvIJSUY8PugUlOaUB5iVTdirVB0lqxapKJ
DCKD/m53wDyDXFsTx5BabQXTWSSVQQRUtrq+yc+GVZ6Z6tO3MQSmYGm5wXMlEmBd
g45URrNTNpN5sIESJmbFMZ+757RJTeB15rgHHR4r7t/TFyVGYKATXe+9mJ947R0b
30kBTowKBnZHnlf1fum5wGfCueEDHZsriYct/TppnAIEw3nF02X99Yy1FfuI4Ac3
TkOg1hgl1overHdVMELNfJ3E2LLYdWv+FotgvXbL9An2/hMiByfMvovp61qpe9i6
Nhr6rbNQ8qVAKXDyR0B1JZXNk9twGVLxjpV/uUUj9gwkVlVAb35K7oWF6aaMm2by
qhBI91yN5oKZ2EFSANHA7lXRzwwItz7+KL/lNakPAve43n9iRuVNgE0mDKS6ze/k
7XojZZGQi+V5D+NKs7IBh7Ix8QGQWdLmzwUE8ClvYICqUz4Hadu5z0NsxzVCiF0O
KXys+gSC8uaAdazCXdLbtIy+Lvyphy7P5D2y4WB+bkFFSG9H+hJltLHq52N4qJjQ
u0eAPX4SlyPvWvSE4JDvp0N9GQ2YRsoFVMc3n9Pn6LdHuqdlJ6bjMv8U6/T1uOaE
cF4YGokvpgsJbyvvzIMhgMj0W7lUnlWerxyt9GXnXQKwooAMj483J7yArQ4fSjgt
ZpRdVtAki3hBLhRyCdq2+zVOlcxUL6hT1e6tbWy8bsSpSCmSiOUA1gNoNd1Ax7f6
DXeEWqS8QRKiI1cWaATcTM5dMQV8Duzu21gKWs5K7f5+M39ESe7CojV10dVZZr7P
z4ehBVZUQ2Us7hyNopzKN9gmzdwZEMSt8wGRmMEHG5SZTNSsKxb7zJOTDFnYtBuY
I83NldJ2Gk2MavOj32m/LEhsNJamb2uei9gtx3sblnqP4ZEIsxrpj+xctLHKTpoe
gtktxRBo/1W1V8Mjm8M70KfZ5150ArNcOIBafOx6P34PX5P/WQtWQIq99A/bSHRJ
1+4skoVXUIneRNnPqv85PqcvCgq5ZIebqkV0ZeWWUVMXE7BfT/m4mpq7yxQKSV/Z
B8wRv50Ay6Wba/KzliWKg9TlJ4YV2RgtOtUXhuvXk0bMw68I88NdgUKiiUVhFJhT
+8EZPOF6/eYqQixoH1UeY4426MHz2ODOU18hqgSDbO4Dthtu1PBXX04cpki08+7F
PDFiJAmCDLMYA4HKwdHDYbssOvgDBq/IgW1OqRMzMUfJNouE1s88KkTd9QgTaWo1
FUuPHgsYVmY94wk9NAc7+GWfKuIUDVA9NvHCxCL6GTlvBC71Sqz2U2LenG1z5d7y
gW64x0Lh4UVLVSWl/3Bho8Ck8421uMoZ5oI1J0irC7eSNlAg/Zpx9UJ6U582EaN+
HSc73AuJIP6PEHngXrQiWZTBCHV1z2P1/p2b3aPMIsIIPL4owpZfyDt8B0EoORYg
Ruh4AGL3rFSxf6lkDFEscvViPVUzQWI0PmRify9xEry7KquckLcZmYPG4SK4Z9Wn
0BIG6fD0JwkK8cpnhIzLAEzOkUnptmw/VKXwohMq2WR2eLC1Z++fzwvcBi8Jse5c
VIGLsIf3XJALntcsAju6o/QO0i0/Uhkbo7+BnWDGQO/5r3+2aOJQWRpGxReyszBa
HLeNl2Biy0StP6oMIOFnQAjRj47XtLhWLd4FBV1mUEzbgyCd2qgqqWZjdT3zvjta
ZcEZ8YZO0ylRemJPW1ZoLOq0mTBVYKMLFLpyKmnDMFxW+KeDxirpCxxvAyWHfJNx
eFvJG1MAgoJyt10Mt+sUORkAObYX3sUfenkMYVkC+UzKaQbtM7BBHRPrcUKPBXlU
dMMBLhYfl4OCBh0/hMUBFHuKOiuW0ajyvOyPCpLOvIXb8C11yV5NZOjjgU3TUpvD
yFTiYkpwTJKEsY5KSstKZJXJsrvdf3fR9vtPF5ku3mSahvblim5/40AhG/whpI17
nCnZmzsFIxkqyUnxigQSSSR9yjC9lyBk9z7iNtVt8mrF+ZhIJoOBv0uMwcUfgejg
uJKKAYN8ryXQkuKay5zy6MxExX5i3WQnNf6Oke5YNTXsNt5X+Z72gw0CE/g6kXjX
eetAa/lfazDsKPeZ7ZnDOcIvz/ETXosGqNRo9CIHjSJZZZpAUOQZBRRYFOW1g79A
2/QtEsRU6S2y/8d6gNmNTfzS+Qtxhk/RAijGf6Pq4t9z2L3htdVNTge7kj3JeHwJ
F4euJ1B4utk2/e8/EH/XBBy8Wddd9xhG0LBuv3ljGQqtIw0WjDBOJDjx11CpIHm6
rIq7CQQl9KQW6Nmm6kFRARWpAdfgMFccoMQn+KpjzXK+U43BNUnyqv/QpseNC9S5
eiPpxscZWBaNA73E7SnexIwEZ/CWYu7unI+NtQX9QuRGc7kroFVhQHuJJFSqNfzd
bqxXL1J+5zJ920h8Rl8ugLI3/uQcwA36derHe0dWuTP3aqgw+TptFXomvOc4orzB
KSp4E0isAZo17T/je6B8YVxKmb1s0tFV5UjSFQpX9x8dL0lo/JVe/7D5cpy9Ya2y
4qPWRGy1ZOIZOBuGsY4c6FfcR4BcvkT5tmJo3etDvJCGODUg9kIretUalW4Yuhkx
N59ZE+bV0OxS/LR/C2M0dSbGeq6Si7P7qog8P8S6tZCUl1EYyUpePRmwvACdaK6O
K7k4xF5krLTAQ8enF0/yrhO/m7bhi/GQbaooZOpIIQXbOBGPUnb4A4BvXnHOHiHR
mzesLGEeeD78Zd+twuoO6OmMT52MteGrFIyGpUV+WQJkPxisTudRCi6MS8UCSa14
JJY41vFZ4SVll4XGCPV9qr1aX/fiByh4iMFiRxumtccwHloRFZB6FogC0nxLy6Hd
b8RbQ2palWLwaVn6YhQ761s30jARMLAtWeWkWEM+j8BsM4XfR8SRy0siIyC1EB0S
pHGke9dbciQ+6rbE8NycsguOBP2Me29fRcqK8uvSprd4eD1PnaFoifpE2WL5muhU
6t3odcE3sx1gE1cX7p+KLVl/1QdSXh867aOuB12pu9UCRGVG5Z2QTRpSYNAOGjPg
rn57y9trjrsMBpHTXPX6kR/SNvcvJsQDYmkcOWZR18r1qSkZY8bTyeo2AFtGjKPv
mepx8JJpYBvjlXsAoZsJWs1FtThi+jTBPM4ukPMIHSDS/i5yzl3sQZJrYSFIH7WP
Hqsiudo5i6OQXngkLXOG1fw+oqvA3XeatGncmLtKvlFXT742ZVl7qgUPngdrESDS
ju2RB+eOW9YtTj9dqwz+/OIWBjLaP5yQUC11ssoe4VVn1Pw9BW5EkMNTCkdJPvWV
yaUK/lL+Gtg6WIuMPvQzV1nWystYTGAUDUULPhsI5g+LgL27wO+Y3lmXMTRZ/btd
a2qdVKPdx0s1bElvp2CIKJzxpJOWTCad3jB8klMgma/Eu53pDRvONaFHb25FUiO5
01PKhiieaCJcJ2ue5Jjlr5cicPYfcelBDCj1XvkxjyfER20y0H7UCuTNJmf+b9NI
O7qf0G/eA9j+Q60/Znfjle3KYkaPpYqtXDfGthQjSmd8WwBiUx5mMgbKEekYDSrG
6LQNTTXvYY/0tdm3HD6FKYPYj8f1nJt+L8a8AS/UhM17/QpcVFPVtQl8VvV/0m1L
nyReEW9KtyBgUBGKlz++sSEvZ/hqhBYaMQZcirJbzMBPT3MEEjXKKOR1vQE0P6HN
ZcqzKB0Sqj+YXvve7vMELIMCrt8yxaKeYYa60ShENEA0qwf9+1IZxldvRn8r/d5s
RKTTg8wJKIUxYEpE77/9K60L/TFkz3v45rqjGK2Jm5xp5QKP0QnzTPOECyuSwW8p
mGZqOq7DHJPFdeIvFXpAMHwBaecqIPf7xTuoD63KkndbAX2rfba6D2kvY89+PPso
ew+EVtl1Ilj8g7A+Be3OJ8xfPUpKB6Fyw6BSTLO8khqIypaVZ9fh20vO8YVl1TyF
My6V87FacWKs3gOJwfmXinMALb3mkUHiy9nalsmNdJJzRKQMXs1/leYs2OSzPB0n
MKlc+lXxw99+PpGSx8gMLm0mqUmChDvyzlcmY89fe4jPiLSH7TIzx2FSzkLXLDg6
eS0UiPkr8Xmu7qwN++GWvKlTqKhe6Jg3Pvsyi9j7dztD0zzVN1PHz+lBxaDsSBbk
YGPQBEC4p679OcUFM0oXTX0odjCO9AVoeWgW+gSG/2OpZsinu0AEf2ffHULF6SGS
YQ6yH9UY7NIIZ8BqodszE7o+Gsu7BQmda+Q+7Hg9gf4oyNFNzGJv4yBXUuFe+E7b
wlqwOFcFQbJUd0dTGLO3FHZ5ijskn1U7FxaBpXrLf9fwzCj4xwsXQHudj2DDJ0hk
I6pBydRmKvfQwoZqFSYaOC16Kd/IdQo0CIAn7kAx0+00031VDI/7dltfd1Kmi9vG
Ib2kAGWFlhZU6lZguk6zc+tKQ6hBponxPxJ5YEZwVt5cfGAlbRNQtW0SRL22RQMi
mPxEv7kjYRIOfnhvFsMgqLaVX6xh8WsFhOmGJMw2N5EvFtcDFkMQ+dMuQtbyXQD9
20z2k2D5yQfXgHcQrGNqeZ6beANsZ70J/Bht9rFKNtbdyMZydM6U3mJToKS2mg2a
IUV1fWbasygHpN9FzFDwctOwq6xp+Ue0fA44xOjPWtSv9BHJd7JDYOC0jtFvVg3t
6qa+xhyJeWqt95wm3+tExaxS0VvZEt4GVZHQzPYUTitaIYcC4kyNtCefc57+BbAE
XQ75SAZL9C/l8K+QXJosFCkrtweqBecWugW31yyrhm+Lh5E6BBdIFO0TI3uD68WS
tLumlAhEl/wtlb8GHnG+p/uQIOU+NUHkmrFck78SKce2S9+qBtM0Oa5Vy7Joebhe
Zfhb4fJwBtDgtGJB3JUg39R8IXDC85sniemPxmMcTDmoYmgGvm9sr0uq715FV6kG
nrDtMFQMzUkRT48uNOmoKSIwrMtSRqjEbFBfa6N7PWMa7yPtRor48l4SuOCe/WvE
Y7o/Lqqad2wuBJmyO5qz2fkqkT9i3i74lVjviTLqn8uNgZBNMD+IF3JgdtrspxhJ
6SN9sEoI8jU14ae3LIxTjvn52m7YnkBBgkSiiay8ZuV2bkJlFtf271g3ltqvCCGI
Q0Ju6m63cvYstldyTKtZhRS+S7pqXCrywVwZgp5y/QQCmYE75uFO629ueHqqfd9T
D2Ov+gLlRjj3eIQNOZrNOQPWHZG4NngC9wryRVoP7+TdR9M/REFMsqJi4va3Q4ub
nvaee9M4XqQ2TZvaAU6u004s86vPM3plFkjyzEJ58fmmy5AtnFuEzABkXuXmhUyb
xgvD42i7xgk7+2ZjHfg1AqmxLJrLsl0krCVw0uR7sKdMaTZbjTvUPvWfJAPNOtDD
/HjbUWEvcovUMX2Um/dMWCpMcjXCzQRaCXkg/64EiJUeL/eL5Om2R8X5KXtZhfuk
WWRMGiEwhNK21pBEdk2IUjamdplh/jSMGngGBwuhQw9eHmRr0DbbqEl9ToPWm3kn
n8/OfCyHblnkeFQpD9LAgR1a7pQKzK7HEIUfnztDeSdQupEgL/UFWP7zSTE35gjP
5fPZ8jzar/n3k6BlZ7nkJTDc4fkh4IN4/5t9OI6rpQmHvY5zWZB84AyRDW7dSbCK
SAAJFqszalF4UMx+Mgwz4StFdtn9b3nzvcabwc22nAnjfiGgWjSVp/PBf5ZcF3T0
2NCMOFxmvENmcz5oyKdfPt5ILimCtoLFa9ZoHFQGT+wRvh7dnpqAHldiDuZjzmZK
jJ2sfDYrPiNE3OrMw4BB7M07m75HPdSG7SB6uqBsmLGRpnSuObgoCsKP8rVEN93C
VcSqOBxFPbdMJjGxR90rnbVOR2Qtl//Cpu2yLrTy7XZBu8DsUTH83ip2oopPh//E
nx22EjmaRBWpOxiQOzo7znilGTEK9nu2hLW+/M57hGdfUHzqNnh1FkiYx+sNXTN2
IbH5+iciUWc88CpNUZWhp3yhUvo3KZ0c+S2/jB8xXh3pAimebj3zu3YOQZhYLexL
9TVaGD67jeAZMh4+Y8BkL0NB6xYqWAcj7wZI7lib48LObrfcHW9IdayQvvfd2uDZ
sIRs19x4PAAZyJpxcrwwwVxQ0Ilk/CCFDP/cRAQeoT73W5xr7PSK/rOzFrOHQu+y
WTE1ozUu0iBmNRFzT0nd3xgsQH0eoOhB5fxD2zosL+OpYRa6uFr5kndhfOtiy+R3
5xFoicX9myasDbPW2xTIzCG5V0+R+hUAFkWAS5aSTTUE335oSg53Amr6+3Glfvr+
V7mwXMwBveicq3XAH1VTdwUhcy7IUbnhg+KZgYBSjVL9BaEoG3eo+eYDJMln8izT
frAtNUUBjXQw2dKIaFUDoLyEfaYv/6cir4AUU0yH6sDX8pRpjZ4C21FEIbtv5Q+H
DQ71ObLv47TmJfjxY+qsYkYL/GIh10P/wWkd4vezShgJadYpJ5AgFOB+8uTaosxn
/M5k1mBhq9Q71qeWVwRXiHa4NfBwD1jYbUyLb6rs4MBT7mGin1ZwtJZp43jXn4uu
78l3aMtNZKS6JyTRYR5qvhftib5xX5UGcod/O79tHNFDv0Fn5KKrtVoZSRY+kWsK
GyL+zt0opWCfOgxUaER6vuDpJcfRDixUh5VgD6ZgKmNaVXJoIcdchUMDs6DXI2bx
WapkS/mXeFWL/U1Yd0IDkfkv3rzIbsao39lObQ3rnGVach3kngxsvcJkY7R0qaZZ
X+K7H99ObzBx1KocpgLjGfAi40aUxcVnp8kIv//e8XldHX0FJb/w4u3eDbsB+f/w
bxKJgCdC/9ZsfU0bglg33LkhzdrD4mAo8VGQX+E4fiIwlKTqvixcnURdkSwBA8RT
v42dNs+YOUAoIzf44f/ywrpw5Ro+r9TMJH3SMHh4vm6LwuOllid97ytDipaolG81
jvgJVu04B1F1lGw4kuUvdVWxyjD4Ws7Lan8n4KyrjNTowKJzviNMrXTSsr3oRR9F
3whnNdNFczZqbv05HtGyUm4TD3uNrovZaC7Qu5MaC5qA7eocl+gMr6uZzfU8BvH0
6tMaeNxfijLp5rUzb2DPfb+RGwunG7rReMrSnXXZFSD31reZu03t8XwlZm2l8JWG
n1IxxoCW0xRHd0tXQ2mObZjDYH+JeaNFpelNPXnP4xYj0j9gAy5zcgqhOwp2c54D
FraD68KYGA4rQlMpLqm1wL6jMrP/dtVjJOO9FSlSvbUhqUPSA16QFnrAJRZMXZ4n
4PYVNDCBj8LnUtarbk7Cf128DZoIWxOO1sLYy1UGLpfui5gtPrnPZd5DymWdEsbN
wAzQnXSBXHyc82HsoH5rFdA+AjGIh1iBQ1D1xRPq9nIU0YQLXVpYp8vK6gKg+fZj
rTCddQRobEO5uwZt7LvrgX/yQyrpMdaWtu4WAxUnjQ1kWDnwA7Xfsjuh1NRlirJx
pGG7gDps/+xC1E8i6Pfdb/5tug6NGwtt1B0WnwPqJWqwiSKCqDzOBCZFFVJN+SUb
ZR0H/TFR7zWjMz96imaY0CFCShcAFyxPc6aFbaKXtEPuy7i0ye/XO9gMKGLzSxi5
xMkQUixI0jRiN+B9Q+XFBLVo05Vo1ZrRfOD7sWx6In2nTOgbDPKQKtB3DQvg/b5t
iH6UembfqAHZFhUOqo4tguIMggAqjEr3RG8zOByb1ZSIN9JY2tfUlHQqeLCEYqWg
FkrW8MDsa3hvWhxwgPl1vZ8aT0wjI1AL/Lp7I1DxOaaMffJ0aayj/bL1OvczJNhj
Xu3ZK6/oDNgXprUw33jiJX1rbMZiWu+nVkkkYGVaZ+1xIBJFIzsl98KgGaTYAt5o
K6BixRuyIQroncVa1dnQMrYod/dCszd5NW0xrAACa+Vg8zpbIuymQhI6lwg8JbaQ
DHrAV6FJDlNEVG48HIFZqzHHvTWXeT99SMyViCqD26BeQ0tuQOGCxhxATfFHNT1O
gIGV0I852NxjLtID+OWVYHBA5Y7PuGr8pYQzE8obqvKY/vPPu6cvmTe6addP3UKY
yvahh4yWgrcJGR7omKCVffqmiNwcuhgSz5QCfhAXzUNRw0eof2A9GPf63DApQeXg
u7XbhQEkGZWBsB4HRgP1PuGefjBl0dSqRY2oMS1lOp2Zpx0N4uvxEgWfSUs9bS+t
1DtiHaLFPg3xb12cxjqwZTHqlYJdwMxmvsCRsO+C93GabEBXZImHciUMJmLrnYns
JlLN+MC/2VwLZYGW0H/DHN1Jt6YZk2Cc9PX9eRkfT6y8OjiKH6uXZ2SvfsO5iltm
tlMtAYa55qdmCl+9lq9AYkBeTVp/lbCGNY+oWG0o27a5sRPib330UjxCfI3319hy
qH0Oiy5kQpljj7pT0P6Z/51ZfyVwvNzxS4v+wVp18PwdOxShtVaC/SXtuXR5N9Nw
9XxStntVA/8VmNUaAbdLYKzoxeIAGf6zHtBTloIfztvCxmAaYHHTM4Wdf5I43oHu
UM6Bwfb15rXoW8W11iPzHxHtIYczFr1ib2a0QPfCmLKG3QNJlPMsb8HserfSYy+S
PcvdGbIM/P1y9YgouzzoQ+C8gZargyG6PJGvg3RCh5YXvj5zo92Klg1+ILBgTwPd
TeqFqzBIzOEmBM8r002xmyqo4I24FCo5PesAPHAHpYXUD+WrDZpY/HRK06iZxTBI
mclLmMwupGNZyvVH+2tYAJkLCXCGViCmfQnjInrgdh87kIzsaVKwe1gD449ktTIj
jJ031Knl3wisGqFLkEiamc8T/emI8ANTzp/8aMcjX/r7QRbVY6DNqa3R+ciTxdyI
yBuxVnEpvyFDNbFHh8++graGPjjKTUXrJGKVh/sJTUMUJMzqKtGZPBJRqRaYmtba
ZQztK8lMfZWdYql63pIpIxnKYsVvsL80eHCPLwdd4fTb0uF0893yHf86dk9UmBia
pkn1+24kvmhuewKcWi6nzhAHXPsAYcYXkE+3mKhOzPfURGc4AqLQBLGx96QBFAxa
zrRoKDipXD949Yo76IzaZ73O98bltB6lDv4UDeK8ePQaO8AbWie4/dFHJSmjPIOy
/nXXN/HBxnccy+C88d7tiVs51rdO/YYzzSDDJs4Mrd3i3+yV6W+/vBw6Ygng+Ekh
L7v8ptzxk7Rjd47sdhO/Z5LtT2RE+WmxzcA+whQAx7sjAaM3Ew8QXqic9GqEcEu6
aceVdONh8U68epMwDnXXOwxGLutFXy67VBi9DTvSV6mslKrrZIcYZ3CVM+k21+6A
ooxn8TlGBDuQBl7vxK0IbgFuxm04urInXNT/cH4w74zHxCLcD/T9XR7a3U7aRbem
D+cD3+MtJ8OSKxxS7doEgj8MV/ZH6WCJchgQQN87ERsYT/yjiMXU6CJR3308+j0N
AORpxKzBkAGo7dm/8JJAxD0+L1w0iLbb/nXn5K6ARFsQWdZFPXiS8SSOnhnxHG5/
c8ccbF00majrWgfrbw+XRlKmMuWoWtmLVPYExIzxqNsUHgWDq4tGi0bm98hl3k9m
N+7RaLxHskDeRFuZeIEzz2klcgOGOyUZ9cVNiCvKC+yM4C8+TkKj4MFh8ptpDC+b
zPW65iM7mK2VLXfWy1QhlIVZS5zCPVcquLrxhAzuZwAGuwkdiXR/GS2ploTIdXmF
6UbJfYOxItTaz4BIgw1XVfFxUVqc6D0rvhz97gkm94dA9a0F83SZRJb9fvMzC2/E
FxLHhJIvJ6Vdm9cPIf6bZrtfowTpBiz50SOjgGgh8soA9sQE/iC3hafFSD0qJrBK
eAvkTtijmYKhSwniiK1BgU+trvTBTlPpvwYN8dYTAzwd33+XH1lpwh36W60ebmH+
Aq2QkkOJ9+hpalOIXluZHyaD/2/X8jBsII5PFy+gJjMCRBOHoSoo2pmf+cvk6lkw
4bNghQBf5tL0EbesalwuiaEzOaQxqP3ni9aiozeF1ZnMONPaGxWLKUJIBBmBE3jP
B3FDu1xSoCtd1DmQ/lvkT2jk6uGwRocUYPYyRfXCqMPkRUD55wNV+f2LN7QIqn1s
ubCPe3/MVPtMzXBO2sk9yT59D0zax++4UwMWI5YsNZZP0WTgdLGdc6m0/iyK6/VM
j75EgTXr2o8cfcq8UWkFsTv3vcnc2SY5zmsajE6Te43wAMjNZ7iy7rpkB7buOgdx
H5g9ZBTWBG0zn845dMVeAvY9axRyB+bT/ADh6XXJJhlIu29Lqx/ao2nYbbRtrsrb
zjyTGTd6ZB523ij/T2orwFLvuVbvBy9BTUyYegJpvmNUklfdZcGJcxokok46g4ET
xNsAcGtObPiqsfLKlmtVWR4B+8ZWR9fxHh+8rGkGoQdyuQp06ya3VfrhEcrxoavi
V2DdL/Gvj+7xryUAKhzNMH+AzR8YC2gOuYPjufOXM5RQo07QKLhJ9R+VFwdW4yEt
c8v+fxeoiouqgK6eg18poSowUQTnXPE5YC8/bWmTQSUgvHnF8vZ3iMyAEWdag/rD
fq5eCjiuRRytZi3tGxW2RAXMZjHx+i/IZTKmQ3ldjuiK6ebxAW77JVkLIeK4tK0n
mvPP37DMUbHa+uHEv9j246VrdknIZzEjbbACzos8ABQljifbzoYnoLOieLnoiizv
njOaV+pB4bA/UavcO8UMbeEEt/AtHwu62pIc1MTvOKiRUlm3RRe0TGijmh1U/fvR
vH2lRmwf+ileDH3hKrTGnRSLnLTCF3jEQieRl+7OyHvDy4TKiaBLBgHw/agGTwn7
WibnZJWeZdKyG0fd5vZ2h04IGgGjFSlusivRIBPpbgIR1S7dJjQrs9kUf7y1bI84
aN2EOtg7nSIwfAONDwM+jFUlSNBi4fWFNbZtdyrpLXPjMftZUehVM31WgXgrE2AC
3O3ikd3ZgfjVW54O4xEGdamZALYAWU0KPuTofzQyD7opWK07N/nGUXc/QmlHAm0w
hUYxfhEZC+moEeQuRdateUyXAorYWZbe8purU5dPCCERPc4IgtNNiN8gDZrmzJDB
Y55Lvt2GQalw0KQ5gJC0fu8KUuLrQPdrFL00OXsJq1RRNHNKI56JyaanzQHn2guq
IuCnvPPLEXutffePPNo+W3kR+GoKNRY4TzI1xEc1OG4CgyLKPTF3QKN+3ZwGTuFg
RwvNnx0YZrg37DBe7Rqvubm5QED8zt1gVPiLL2fgagKp83ZFP8bKWX3dfdw9E032
cRlVDlz3D0hnt9zIp3y2R5D4iPWilEvERl8wCb1AEDdcwEaBy4fRBP3JvxPdvt48
G/JXPJPx6qMZO+aE9/rWZYbDMmizOOdAnbeB+GLIKASB0NS1BM04/sn1a6GIrpLS
NHnMMgH9wo++Cb0RItzUnaY5anyfQPpU0taeu475QsfYN6TmvHHdqS/NtvxVBDsb
i4cLgB6HkDCIFqC3hB4VkgDLgoIk9l2VVedyIbxFdbUjXO3DvsGPQovmHjJaI0+k
y2bH6QfW9JTm6mQbdRjWYJylGRQIAn600MnSHGUrsb0bou9NQoYJpsi211T/0msI
QSKFAflttLohx3LOhg3AKHLugTYjhqGKsN3wGHloxVEq5W/FOo2QKnRx0S2okw4I
iAyz6vPSAB2E2n6eq/9z0nk5hoy6nBYnZjzK1M4z37bXAQTkwjd9FTbOKXYzrgNX
JmfWXtm6qAZY0huftbWNMmIGjURdPvelBhudhMEc9BJLiaiovlxrHl6qQEQZN1zg
08EiI7XOcP/+OOgygRKuNZ2ovE36T5JjuGvExm3k4lqAJZqzfnU0xQNp+Zh9mVtP
tyHD9IT+PsWBEb7CE4mCunFIYx9OIgPjf89kbSQideVtqAfhQiw4Ro9hVkbfR+/I
OKr4HyVe8uFOi9Mu/0DoyZ+o8Hdv6XTTnLo8FhL8Fca5Zi77Royx95TDW8NFAKNR
YLQjJKk/31Mdne050hm4zxE5i32H+MLGLzBFHNs+N78JrMPH+9oNAS2YyhZcd4h8
vzQoihNBG7FfgELgTPPi167AD9c5nePdqW0czWr9jfCHl5TiOINta9Da9FrZ2QaX
4lwClHhAz3pe2N71VmgKl0fczN6rQ9tOye0125vkW3pQhchYdruRU4CLLTcc3/tC
EKsReAHzOBjJGq5wP/MVBvreS+b0ZHoIaxIs0Dkyfyj0LjiEi9w9b/Fg0x9HT/aE
Khoq2ilvwCu73E7p1NCRc2sRrnQs4sMgs2nhVMg3ybZ31Teu+ZZ9VBACZxDc4Jjp
yvSKAzw3XQtir7MIvm9LfrrgehHSX+2hR0vrtbe1O4nR8PRe4I8LfjDOYMWA+d/t
hiKNpoJSVw792zTQ2u3j33qYVYhaKjsiJG6fksGHxQmdVdQB1Bi2TUDfQ+/zuxVn
LSygCnmLh223ekddcdEB+b5ViMWdq5zg6w7WDImKWI0qS5FQ9xvq0T+8S9g4GJM8
Ev9l1LsxxJDJzORiu+AZqdKI0F5TwSb3GeXwcDC28LLJZ0PN3sDUmETu9ZLP5u0v
vTe8HTurYFXPjB+0ovxnjajJ8NpXTpNSgslqsTZY36/7PL6n1tj/iKyweXNaR+Aq
+E+QSJP+dvznmXD0lxfY6W9NAcWn6jWzLH62AHFTNsW25eNpqM7PMRDcC9jIA4GA
IUy0szqmWg6cdoSz38rjmh8gWRaStBrxKOLL6rFrJx7eMMVqpX993QwP3SsrwpCM
3j6nwOwZSejZBSv96eXQ/Ca9iQgvtlNSlxUHllZ8NfeumLW1pci14BY4uwU8wP89
6wIPRWMOdGU/1tJIVpai5qXhA85LrkRs9fwjpKACxH5Q30jGOZGDbkjGvgstTgOq
ZwVPtQiVC1G+/cbKoWD96ENKH/ifgN4J1M9wiJ2Z3UMRYxUhfwZ2bKe4ED1ZjfHv
LSNinT7auA96S3GoVXTBRL7DJnwQtPP65JG4PexRz2xcaBusnQ+aLz5t1Kt6kQIW
ZvjbZ1JSbSbDYa7bV6y+ay4PNPoKc+uDRLQ+PIadBgxmfiEBvdWu8t+kaRvYASOv
yiDAwkuBE2AxPL0kvnhwBCnhMmTp4mpy25woRdnJq0KlXHrH4bqowk4ZJ+wzxVYS
LhHB+ms1eOxSxJ9gG473ERAtXSGsrv80z3wh/NmZEaVKLqjb0TKlKckLIkak4jSq
mjZI7fNYy9Vm7QZgf7eOJIz0xeKzKtY5vjm+J+6Nvz0YYoROh45NWQSAr7lKAWE6
fXZMsWScPKpw0cL0iluMhxbcPSWXJHkNuERWAIySrH9aYoC/3BTU3/m4IAYpfZgJ
9SYEe4OuSQS3XxQ1JGh0BHW+BzxMI6sE1lTm9UZMOvXISikeI5rjkvxzZOCPMl0u
qncKS6ywNtUWCxyty40wh9HXFIXmM+F/xykESPQ+788zmJKNJJB60/kXYyxXR5t3
kPuZBanj9Xvs5mOrKyOjLwKSmyWBkQaPu0THW5lDSNTaJJNK+szlLmrIX6JMx5u2
pWj4c2aozkiGzcFIOEvMYjByQGDz6NBhDpbK7gouUFb/AQkUUUH6I/bChvBhD92P
AlioF4SHkiXiWotSDIyOHOy8mx/kAxJQ0Bpw3T/TOdUyqkC1ea5Yxoumx8rWbHVM
s8fjP14JnB5LXbE1zL3CTwJ4XG69wHjcaH8qbe6sKOzFkGjWv4TZKR3ZmIy/5jfm
VQzg3N55rlYICthD9KNdPMGXRwwwTYDLu4vdfJ2l75PrEEj6qdohliRAGhgb68zn
Fi0mn96r8jQmJoghRpZIN4wGhncjWcaUzsqUbb0qxwM1bp2INVWRJ9ztQ7IXHbbJ
44qJfvkqSgKCUqiG2/jRnr6YE4MC8KW+Zi8dvVcoky/N0qC6Dr+U83INYMPiQk6V
Syy9CU7/w1x5meoG01NEoJqFfftccsK8B53HEliE1QSIp2b2CMbtRj8gFWDrbP2j
RYAr/v27FaCJpRCdnHrFrmfgZiwnTQt/vMROYtoS6Cf0hw0VpWggBjVjE4kviI+c
ctzCiObLpXkFLSuMhhya3wiR0ZCaWKqPx+YGyv4bX84QEjrbjNmm6z+90pOb7zne
Q/WLAmtCaLf+gAfrzs9qcnxbtsMoCleB8DoWQy00KKtnGNR3m0QXKeFD0FlPzpBI
h1Yyd/h6PIpj8RQkVlV1DEegWbpATeGisixKsXxlULweIyj0t0Eo/D8LFr/78T/t
bViuVPnnGSbq23VLI3PZMwKexs5zFQ13paGcvN3hCQFcAxJHOHusIGDmttXxcJeZ
y6cZKHVffogFI8N+bmkJo+8mbCVdKmQ2WvQ/za4HPhqIdOmBXFCJElSv84uplThu
JpmYnfJWPcxC7bMtLUPeq3oeJSx6LSiAaPUaZRCZKJeuIZYMehJSgWm0e818Y/OU
6lKqg3hocE0dU1ivlHLAvwbC7RqU7FzfePP6OnXI65yZXXJSgg3LWSzA+cMtW7iL
HG2gcrGVLjL8svdgqwX66TQoELxzlq1t4h7FY0Od6YDIcw9LvBAtVAzowKrVwxcm
WvoIqNy0m6+DYkDqZWZz7XQX8X6VujQ9JlYtRVg0yLpocpJ4+CrSnlkwNjiTH/sz
BZo7HCD4J+d0l0scX9phCaFdiRoHZwtBxHdICupNrkKAOxUP79XAD6WFK3/sTzDH
zVJfDKshQChRH7IukV9VMc1o5Y85AvhWTJL7xY8X8plW4+KmC47DQSW/YBwqAh3i
/staWawT7NC40N/LGs9hN+XuqbEpPms6e1NKFDwak9+hYlNWxUDWs1NcQZQhZ9jX
zOMAoc52Ju6dZLo77IvgtgQndm3uEc2HOdXqpFAoqPWPdHIo4KTmbO88iCtoSDGp
ppkFpR6gTBIJg+NsYhHV81ol1CMxSEQy4r3t6YyQ5w+A4tSnaz4bSd2c1ZbFD55K
oSaJU5jCuXJuIFyTmxk8KNHfcjociobDH7Cdqgpm4wBGXZ53qj5eyRhc7vO1BaT7
iKN5S/TvvwbOGV1T1NrIl6dqVGUR3tWrA+9BRm9YPwMRVf806Db+Ba53Auxl4Ien
fqNNcXfJyj6f8wp8PTa0faVrtclGg7aU5d3XKxu/35Y2sSC71gvrjv0+Ocdyx9Z/
cOFRUyn8p568RW82CBXIavnY6ItX9O780lmDTCGjbVFo+bbUyTt85MrPJpq4DBTb
HMJk+3fYxcqmAzdjAjgm/O0JXG5YHA4wuiRAZ25vmRwSQmUgRMFXsDFoMCsmGfxI
QuUrqzMgrelSyZVNZpTU4H0m/3lfzpBpuXVUzgrfo0OlTVMdn6Z8DfVjqYT9XGKm
f2YRTlgz1LLCzA9bhzsRdCSTlpZqEEqUQUz6nT5F9KAOlS69uiSHJFo+5mMUZRwo
Uzk27HHWUKi+novi3JXmnYtl+TDFiOIAvb7V5RwNFCnd4mzQW3vOnxx1nhGO/yBc
RReIfBJv5jp2cLZo0awLz35cGCAOjr1qnHi2E32crFe16FGnKBUyueuwjsR1dbO/
fru6wo5hh+OJF3FOGitODk5drzP1ihy+vwrcbEq6GWL/zWIVhyvVO9F5vrEfGzfV
XFH3V/P+uKqhsh8pNiegLdd06MOY0SLDlmrGeBV/Jhi6COfh6zeGf5LHPmhzJhoK
p696lTCWIPuBwpjU+KM96s7og/pRH2reBgADQPveydafQq2vdRcpcNWJHtiTf+ow
yu5BIT8kJJbIapqciIPKHSb9i8dlSqolqV1+qgykCAc3U3ItCbYPVe8xzri4Af5K
FtJ+7+H/Mgkgi7y1zgAtwfomsg9ZOhx48OA5w9IwJNCTVfVgGb5X6C/CxGI9ogY9
6BQseRYnxe3aIvkyCLV2cwqpsSHZqf7kSXh53YwExRQmNulqjlh20MzO/P3GG4lX
zK7VN132XF16dcIdYpRlp0MVuCcrgj53s76xXI+qarOqyz3/OtQXuGEdCMrnT4dZ
jbhH61Rgzv+ltPQJG12BBSiw4dhGLL4vXppTsQz2g0OWvTwJ09iJx8nmyqcGdEqN
GJ3L6dP8Ar2IsPE82ZQp23RukBdxo7ra88NHFFpFDTbryvyl210dv/8l4AseD7hC
hSHXhZYZ88jZizJtwvhKKv7krSbAi5HwiQZvn7C06Dn1QO4sP59EFqkyP1v5vikp
3BWvPk8SWHKM+xKlYMMV9X78sdxc0ktBTWgX3VuoQeEIJMm099AHYxmSFZKrSBHn
aQPyTlKijSsY5qlLxIwMqVv1SfjN3iH5/t3cNalOenBPwm5HWCdmu0gWfTcx7pFh
6GiZLP0HShUmJcKsxIr5bjLmv+z/O5+ZHQ9dIlEaUk1qJS8QBIvsR7EbNZx29fIw
tS1gOtYSK/69YB1OU1XjQqYTOvuItJCXwC8afugsstbkTyr+Hj06Ld5gS5EMe7TV
v/nPmMf9GeUiVeGNIJShbh0356sXYJvVhyNoWgin1XGh67lU6f7vogbRoagyL+Ei
/drZDk6U8m6CJEt1sVI61mkH0Cz5PMqgtXutEKoymK4u6fR+MMCQHjt4BvY9qIM2
UFjlJ9MuGqD7s0HTlg6+tSwt0di1liOmLZIPsDnJnsWCD0rMKSn6D+did4EqHbV0
jJTl9VwV4jaxGB8xXQuvFrbKn7UQ8bHl6krk4iJ8CWyJ/NXdlQg2FCFQbBe1uFSB
dohe/by9TdGB8jifOdmr6jbvxJMfVyahVEbXaw/12FCObcbyJNX57MiAL6+WMPPl
QVRYKRzarKQ2DuM6WiAXMOpKAH8SJ88fp39cXU+pIILoGsH5zYaJ0RhxlupDVSHd
LwWFMG8nfgdTI1jbgYRK8QN4SYsZW2wPLSvABInfPSvaDteQkyFSK63p0IB45r4T
a5nw0oMTRcRip5xXg696wCbkeCARPG6tgM78pjizZPD1kIWXYRcG61dZK6Ig7Bal
lD2P0aL8OTD4T6MJiVMXJKcxGYEsMVCndO2jb7MUb7CrxdCb7NgZUnYCSvs+7oJm
Usyxj8AJNynU54gmCJNYc9Q3e0ZJ7VpXjZU3qH14jxE7OX8wqoXiFYaAwWewTb+a
cGBx4WLX1MZcE9eOJer1d+wWqHKUsCs6IhyZRu6bLDexQXqqFvqfrGVtHMggD0aK
GjTjgvpCDVbyvCNu6qGVF7izJQyf4CrnxyHipIshb2cejhqXEJ0K7U3KoArHrlpu
uskdj4hbYc6luQtRsPtszCt0LmVsErimy9llmqCcPPeuaQHhf33mnow02KkMIeTR
p9PBOLWxJzV4+oxMdP7+65zXQd/IH5qVyjWOfZIvi/+SqBZVxTb3Qvkmwe9rqQTA
GSvacaA6MDfE+krilflu0P/cLLVUf9kTdjXBlfNjPdLDL+YmGLfq8P/Waloci22W
AVjXpxPu+BsgSY7d+nk35Lja7sHLfx1sJfciCR/BmUEGSaulVh4/TXX3FKuVVg+c
Veppqk51ctXyA9TVAkFNQb1zDVYnNtu1xUDsF4c3ZvTGTLquTBTpkbO5qVpZEUaS
KpJ+aA4hkkfoNYvdndGnN8AxFyyHlyvbGo6aWF9YALuUmmIUOJGr//RXfcla43Kf
t8E/CadKiMyp4DvZjRShsoHuGq1CA9aeSSooxIiYKcyH2wHsGyzQEHl0npIUaGBB
PSGQReZlvOGmtX6c4FbxCOTfrO+UdESp5dJFYyUWynwHWpexxpcRxv1GYkCR9055
VmCfz2gWmd19CzPi1fYRPP9+fzYeuxsfojheAb6THy72qJ3dSoSvKzi88iPB6488
ZexBO7b+g5hXDY0bovehhRbGJVZBMmD+PSkapeBO+zu65MKXdarqwRwYdd2K0U2y
rH7lhAdcVGr6jnrrRYZHe3CP+a6ttSUrjN1UBP6bgYT6b59/Za8ne3TyetEOq3Za
b0Tm1Fvf5pjn8B0incIGcpuswgI9ddDYjJ7BeKLk5kW0umCuOqWuVR7TTfo/0uZi
9Vn7XU/cRFeGq5q7yKSBNvDvuY/6bkXEgabvR+CA13rVHOJCNSwcJIL1N7ms9HEc
E8QeR/e10ewG+YiQ8J4igHH9ekW2ddmlywwNHe0zwG5SgR/HSUNcOMalIKcb0Q3r
ur09AvrQNfUlvSwWmcRTmObrKGAwB2gc7+wVNkcT+SjC5GaEtSp9Uupd9jm1YJCo
hC0k9OzbPbSzGQPmlMa7eibtQQ32A1G0ZeJ/gawNZmRRg/mvfc2bO5NEDiTQxFUQ
sTdA31C4V7N/zklqtPcf6EbHs7l0t2nhrG0+59G9O6oqzwBXyOT85gpHz+fr/8Na
nshFAmA5IdpGAMvHGJ1d0yZS6HzO0ofMnZ0BgCZn4jgEAfkPf3nN6X+JMN5D6qrc
BTAPrLaz3C8BU0XE6tcD82NE8q2F1M+h7JE5Yuh1BX0CCdG/9OP/05u2wwAYfIGK
zrHA3LaE0+55lfOwFl9hp7LTpSQJAud/ivxT8MEe3tsjuxzgevBcTSaD5CLjWdMU
IylueyCdM1lA+tyrP+grSIfwkjgsNHkSi1xE7L4HbbRKc+6zMsGkrWeekZ+z4Wiw
VWbfvo7NQWZ9b2+YQd4oQbWqP/pc2mxmtUHViOkXi5jgiDyOcVXm/pneJv+vV2f1
00ogTyCg8x6mJpMVtyW9wW6gsb5bh9L6emWVDumqalH6tmw+gkffS8X5bCm1nZkP
0etzFmCt9+EaJfNT5r1drFRp1Ir+iUMNN5iwWVi5WP70uh642PkLzGZD/vXEK5fZ
Cvc8OVBK8Q9bt4NjPYOoXsRYDsZo33MBcqxIA3+nQMgUJFQMCFIO6N8MSt2C5+7v
ZezuApnCJmyY4Nv3FFK3IOCfKT8T9p7MQF648YaRAWL52oz2fgF9JzaYQJaV7MS1
h4cGLZrxHA5eUso2INUtvePIVviQT8ANE9v5wYbW/WK1l4ZKDQI4s+nTYN6mtkCJ
xUZOhaXOfs4FzgjhOIS5xVbtQmFThVDmiBJpaX2aFqHURWBHrQmt2WScVZLp1jpu
Rs0GZgH0rG1Zf7mAT0voVUXKGcvltnyJIoaRPx7l9FF9vf0l0WDnNBJh7ZvoTyC2
kn28KbfEsUMvNANEr+5dx9DmXa7ZPLHB3tVTViM7qc/HHRj6nSZV4TAnbqFfmpbS
ShBiCh4JTnwZlZpExm6SZKhwPaWkpz9dhCseduvIpOMKzwyaQaYgXlfn9bHS606q
ktPysloZCpol3E2pvPVxvK0tqMySqRe2rKBb6+KbtV15DmxehhVHM+U5jQAi71ba
3IpOhANNTXz7lXgnHGjI4OYbkFJKyHT1V3GSORfEiuS1nPz9tzliEanBvwAZXDx7
QNveEnK1/XF61tnXCUaN7xourZ0RwtZIOiJxwq+QaT0Hmd4PPQPgyKqRDaTPt4OO
WQFK3V3g+Lf0qrS4bVcRq3S12j4C0XEIo6AMXvDIfSS3SMUO3B9HK7tlT5RPxjtM
TWEWq0YxGNuhlLEXFUqEXk3is/KrEpEqle/wLF/MyrZD1FXPDBo2vPPc47e07bQM
jxzy39SaA1VAtreUwPZMczLQE6Prf/tbIj1FFIWM/srfvnVUiIcspdYKqEezWpMC
h+PUtWSnszv24eQKYjnaLC149yJYfj7RXHUfgZ+S76QrboK6aBVgsb804FJ+M/FA
6xGPt9/3C57ZTVko0tXJGN1v1FJTPa5Z9p3snmpYu/0C3tQOGlg4CDItBeQHTmj+
jqGufbouAfNwXFnotZwyUg8O/dw+MRF3H+qVNZJye4dOVoHcZ5gz00nUHEosuDMu
0ggY0GZkyslrxGKiILiIGai2Si11Z4QpWu63w2ttet89xAKB+oTo6eO6vhU3xFVV
CTbM9DdF4qyxPv8WYH1t/KqXu4fHc0QYCQXWu1q7Mayw0poIxCjsWNsZrMTqiNqt
JOsHmrGVn54zRxk1XLst0wV8BFMQog0q3sp1S/ReKI3ILFBw5ieibNx9iZGzre/E
Xn/UlxLMF+KSMWh9Y2aaWM+5HCLmCWS070g3kMDNp7yPnxI1V1VtXXBmX6Zp7JRS
BizVSmvx5Uyms7kucIyK/YbzlifloxFEOBpsrYCSRhLaegkt/u8Ybr+wnUwM5cM5
NCWPeOUdyOj3dnGAk5DrtCWmJMm2R4+HovWLRWiaRB1OaXhaC8QsrJ9HSScfv38U
n3d7gCYravH8lMcPUAESHLehvso6KrafyfMhuc6kG4Jhxt+vvIrHKozN4XAnG74i
A37aSiR0BJXfTqXm1mWm3UAv7qmmlEGaAK3nF1qL1z9ehLZe7ZBJcmqK7w/1x3xy
iNDfHQLl70MTgONSNmtCc+lxrShoisjdvooXr+xdtjYmXYLOc0NnPDfSWDARm0Js
1TrbN2PcofIVTMX+MnyTCMJSt0rjzJmDAQzQEneRjjXGuHOcJuE81N87dD3mBOeZ
MIPgOAiz7z48jPQnF1zzRU/mLWeqVRbkIdT8U/GuL7gwbHFxTVjfXpaaW0Luo4BZ
nfcobyb9sDZavsXynOBTIoSIU45+aTMjoyzwLMM5SETBvewzwTS5ik3PzeCXiV/p
OGEbaZQMVzgBTXThxVtbLmSYeHPIt26ehHt0srtF3N4KP3kjp3NQ7MLxYCvlCRXj
8WF2HFMUVK06ad0jZ7ZnNl0NvhFJkk/lvTXSt/Pb57GazDfm6bkDQiFF+qI1AikQ
IMme6wD43df2+HOxOVdkDBiUjezWa0/zlyu6nZ6/3+8s/44Y7OCsHMk3jEptXOKl
xCsHd4Ikyg191l4DhK/APyeThpOuGYJoq5XJIF3RazjWQZ9pqfxA+TXEmd8zcy4V
7IfbWmZfdMmhOA4dhN4talRukb3AFmsEnlR0FYEYd/0mZ2QrU1wbVcerF2aSlkSN
P5x6kGGm5MvXLWJXMkrcuD5N2YyPMsmk6njipVTDvgnOW2hF/ItB7xlBlvQqgfvc
h6Ue7oXyn/eJ4CrnSmLmrpQQaY8I21pxUV/NWKelJ/xId16dIIEpFUZM8Wfcy/Z3
Ts7M1mO0hdduXlvCT+CP9T4lVaGNXTyoFtg1pL0dp/4/QB02Pil33CZiJhJDPn6s
mp7oK48F4O48Q4YPNvoiqzilWTsiFeukoJ+Vz9vaddU50IZy3/CyxXv4mvFN0SJW
7AEAo0tjB/i6mMB+loFPuRa/o38L9c/Kox2aPxMT4cBjJX+xCZnnYByST9rThmWL
qFJ2uY6TWJVm9PKkRexLtgqymHI8qx1cqcGC/XeZ3wkkKW8DMJYaE67oBvdsHgyE
EP9n6TxspEuVrdG1vJnmxjEUxMhsL6ujv05vYhLEuF5nNnlEYFlJJcmjIJ2vzT8g
KYRwc51U1XVALT99laO7FiYx5k6BDVAG3BODUoTYPiDJIkIoDmlacSHsMBsgqd8C
iKzDX5gAAOE3Gg/3Jxc72c6qJVGuY7wL398v93wdyqyoJrOIQphxRpd6nGMwh/w+
CQM72vs3t1aCPBkoRbS4S2ixthtLFNVp2MKssbp9Tum9ikoPBn4qEy8aFYhJ47Lg
7JULCiZKFVUCu9reIsREL3Kt3uirHNUbJUrhS53kGjLVzk3gSbxApxvas9h43jwu
gAX/Ec4bkCuham3miqyv/2ChHHX9c7axH5tDE2dDQAR6rZoMDnItBITTjBd7bapl
gScVRfBfJmbwxIA6d6eRcoyqvzeyoiJn5D+ABR8k57wJrtcYlG1RN7knFhDYpB2h
iW8GRRkMfbbVSZDjAFYv0xzmuVTWxi8FUiAozTThHwNfY7s+xNSpkgETcIm8XIGx
ydUxNMf2otZr6RQ6XyOcJLihEAod/lxehw2hzPGHT9m4U8sRzbkPBsajQBC2e5WU
fqKsCYxZFV+CjcV1h7GkA2Krr7UJNuyIYniGhK0xYb+tY5PNvpSohpzmYTi/KOEx
sxunn+gJf+KvKkpVClJfsq/13GQyTmbHbYSozfCscPAFpJqnSJLGjsEjksgIAQZ+
YMlBfz2TLk0lvGJjhqs9usqTQu8vVYdhLBc0I+DopceKBzdt5ms0uChvz+iyKqja
S9kbmPH39PkZTwOoUNgvK/agJpAIQGcPYnvQSsoELwrqj65pd71SpmcoMQT9EW5i
yUwSdRI/hKnQWQbS0U5Nl0IBe2CQfRFDVqkW1p2y7ZgXqXTmsXOVu5rcCtMMUsNY
xe/TgXnyM0JHmc2bJbndr62zMYftGbVoB0KEBpQkbLRZzQPsugFWhGQfSFGizvE6
rfmh2x/FEX/pvlJlpu8J8Ravt58tjjOQFSLjO/6ta0jiVEc7rg9UbNwCay1mbKyt
4o20FrEGGlYiFv3fagZeAjWL5sxW1arpmoFGlmDhiqr+vBeCol1PgnIH1EbvLCVj
HNYUFjr/mQuPhkxNGTSHvUjbd8kw91GFVNeb9hKLKGxsIVKIhT/6US0DbuO24776
nwGXFbwjpHxm1UtPrTm5h1p54aNZvXKVaP0mbhw9lSZj5SKnyk7arl7HkdwvDqgF
EwfQWI644Qd/9UbWYP5dEYMkdJr3KAL9/RUQF0frJHTub58Ux5NC546F6nYifrdA
y94t9O1M6FEOEdr8Em9ExCrsQnjVMzPdUXOvBjx1bzWUBYZLx/ZTEp6al67HYXeI
rOtBdzyx/weVIo1Z5JIetK0Q47pvC68ypOKtTe0HUrPeILy8Wo89HZT/FSbRUrV5
/R7/rsaMaSfzKtVTmyJq8GER5jvkpa8gfsp0sttfA1Lzlcgr7Qbolrv7mzJTgJ+H
6DgdBB1KkKs4blsnNJhIBac5Gwvr83ZZT8/hH2s1IhCbdVfcfZOHp2OhBu5SF0jp
pKqBr9pUqHGBVQPEjjclp5yNMrit5aeu/SrOoMCPUz3UqAOoZuy512fxeMmSPbKn
7idzakENdzxD8zebsuAibxAKuZKVemg8wMqAUNPRAUCG3blYCjzyUpOjgXMPPBVU
R+YyiDVbZ8B7xE0XoB3PMl5ZZylU42eBBkVZn8yE+3xrka9FhCr/Qplwq6P/jZTv
PCt9YZSdJVBxv/aB4x2f1ObmyC7Q87Narf5rGgqZjZVqxsv7QYK9to4fCXHZGK70
D3Sos/he1RdtCdinXZ3NH4pVCUD27GD3wOkwEm8ZhpHUNeL2WWJ1vYC8dNBIvdBx
fZBFOEvJ/UEwFaRFppGPDBjcO5kwt4JQnA8RrzBs0bPP5tBerXJrGJKcBzPK3fMD
9PsvXD0yFQShGiPfo2owQ6EWQNd5EMs+pMFan3uFQh+ph9/8CQ3M2iXhprfhCX9F
b2B0eJT9bMHx58EpOfn4cRKKww2/VgTpLM0D3mdZQyJgYU1sN2DlvlfW7Of4YKJo
1TPmEHslb1PlWNKHIKDr5zr1TylR9PoVVIOPpyizznlALslgFfYB71ALXDStKNYc
amNY2V2SfMzKkq9uraLGKPyoSYyWR2qQDTeblFDsS8fSnKRpHBSe1ixFuESN72OI
f/98NCO8rzgFyluDLOId/Gl5vSz+6Uwoif1ME2pMTKbqJ3w1NXopyq/FrICbqrqt
Qfbi7L1zU7H+7QUYGseGnxz6WExZmz4M9hlTQrLR/ZLfxpH4zjJfkNZx1+AEybgJ
eXhMG+qKpPWss7bjbaiBEnRo91pvD6JoYGrJ2nouWSltQiYCgJa0MvnSRK7iiIbN
/svXfN62151uKNTDDuhvcHxLWcRPtcOBAQzrQ99vIgkcVfSRvC4gFNofbdZHAJtt
YJ7GeCC1DVDMZacW7KTPob35INcY0NLo0+RNHDc1W1ZwH91/T4yrbzQZHGUXTP4p
f3TZtiKObzgBPLsqqteghEWCjZn+bp2/RzAdUpDj0KwjVwjv6JbzqUhMVRh2LYnu
1AXcYbFgkkdmgMW8C98ygUpOF0kca59rVfEWivOmoJB5X1qF7PbMlc0N/gwGGtbB
jHbvssf5WbaDRtG3A5+Shis3azdnRxSBNCGE3VhJSP5A10SGDfzDzm6+XEjofgJJ
2io+vYiwaeIBK2pJjK6YUwiLadYZtlrQPl72EqxZmgYBb61eVD/14ReN7+mBU5EF
zcLr9MxhUKlVz+6Xrwnqw3kJdJ1mtm5/MZ4koNc4YC+M0JYveFBhPpCzk2W1ZbSL
qOov13eX4eItXUs0oQZFaf+jaQraOjc5WRIrXK5RYMf4gZPXZ2V4LfP4RngXn7cg
I5UL4C7lL3ZgtPiq1TjeI1x6M+0GrCurLEMM1DLK9OEDvHbfkIYE3ZrxnhZ1p86L
rELaY/TlCzyiO2DiQiopMelwDxAUbFSKNfgtB0Sd8oPyhohsQ42dLWy14owa3aNs
TCONcdic06Zv2W7bND84hQxEsp7OhvKb0WAlQ7jcmcWNx/iTemVYKBFIrSp/SRIQ
82xVYNd+Cszx62mgSogi0l8umMQ1YL3T2uaUBYRo1YJWDjPwHi2TnvykkH9dUAUE
h+xS5hY2xUQH728bgQwPfd9bLRqL0F8Ldex4MKm/g9OrZEUNx2fsSwGgkzWOpy/a
Hur4n1glhR0ocMGZkbaAD/FEr945J+E1ysNTLtbS1mHc+8NPUpQSwYYOuWpC/sT5
Ie0ylmGqyocHaUNSua9cFvk+x/kilJtU1Bi3pWfQj+ibgDIKeu/KN0wYwFeAAmhp
iVT40nB4DtmOkA+ol1CJreP8LTxjtdIMnaQqhHLrDdI6N7nu7MYJUTuVglBnnvcu
9prprfCiZ9Sz4HCUpr89GUvAOLyYgHhJ8aTJqscXc0D+dpyxkmE1uroSrMZFD34G
nq2bdcHPgzkP3kTcQcD+M6NFks5TOUZnAIo3ezAH+nwW9emqSOpJMXTqXBB5u2fC
LZCW2dqbbkRjVODv9g+/5hFNRzkvBpF4Ci2gz0z3zDfeEWDiLNap0sAxLhK0FLyv
mml6Y4p3b3jWIBraN5BQlofmQGY593hPsAoI931IpWmoM7Z0FMVyOzIAQb9XcFh3
PckW3FGX6R8xMMD/+skkSnooqlckyC7klObXe9vSxz5CJhaHktE43zJIWvfFZ6oH
0ETTam852h1chcBv+gUnNbnkmRBnloQVGS+AeXtR7laVRYUDu49o3ARz5wzNXrlw
ato13dsCGIkKtCvJFh+VskecEp4M72heEAQbozRfPzFaBZKTFUvl3FzD2SEPogUe
6TRkK+5eJSFxWdpY1ItpgttGScWnc7SxLk8HyMa/xE5ZGEe3imBKKNTYoIrs7kjS
pegOvDMOVIwA50lIkPLM7xXLFr8krZQCFkTGIuPQBzbX21eE4unOxZDgx9AYat98
49xjyOQz1GWji1zMjpIxaViy0byMt+5LiLrWFThdYV2JxGaDlSdUrNfpqE242rpy
sRgJjyTrbfWkM9bNsmVllnDgwjc4fHfM8+V4nBZrB/oXBXPHUoayh47U/8BRubef
97ljALnIHivDnbVwjR+cZzFq3aSg+5WoeeMtaUzv2CP7G/8Keo5n4uDkynOVhzv6
Smn9dA5VM6RFaoFdj5NXDea3yFy2x46aAZ3nqzteeQ2SbvOEfnsqhZIe8filD7zV
sULU4t/NZfYgI5FxfBVKASm7mziTc5wnoXDYojil7yMbDC0/ND5uizOYs/GRGDuz
8WdcCuypqH965L20xiu6eyIvR3z0XE+4YF4g/Zws9Su+ZZ6whIVef2IaKEe18k4O
PQhL+9SHW56zgwPQdp8pg4MSrvLaC2NZoHe2KzbVSat+Z7tC1ukDE3ALDNLxKzp2
b7EnNVZiopQW9wBc/UeIsMA6B7iQ/tYrLmBE5LS/XlCb3SqgPRfqpnJtETnunXuf
XZ4o+L52WbM8U/ulIMFRejl9NMLS83FLuz7kBskyPONNVqzSKmujxL2/oSMAN/Vv
Plx6gWBqa3KnSeWfF8OGqghSipri5cNTNPpSnP+i98k8S5fqPn9zMWUOXJka+AZt
5CO+/ZuOXlrbQqoX4eU5LiyOSAGakQkV93hsSopFuX4NXByAuVtAGiVdTwXdHgwi
jS9935lDIEfRN4+RhiVvhbgl1l9GPSADL3WNP4fPknP9Am3sbgU6LYyNhyFjWqMn
JGBsG9YZGzHugSsREFL4FdYUFnH5AStENJY+qRWkGxD2VYbe3+oFeeA4og7PZGaB
vyQQnrTsT2gV+BVPtCNoulKj1xEFzdhk5iBTnx4amFIsCal1JCJ3tvoMMJWhDId7
kMNS4n+se5k5YCoJnrnm/xyAVesR5GgWpFyn2ayPilbhdRhBQ6XTLqci6yt62X7F
HKGkhKoOMT+4Bk3CFM7Caw2qtMTg6MOrw/y+MP89Anq/v9GkPGdWiEnL2Pk4Mlv9
Y94ZnWscRfNLfRk6pw1nKxsWXXdkbR0VaHZOp4Qedawt8CMnYyZzlnrqFgm1BKnt
z3ZGab6ghPaE7zKCoc6hspvjzXpg0EcsP0xTunFCLCJf1oKN0tUJp37Bfll0dyBo
YLdeCVxO31asJJ07tZO5mTje+Pu2ZUa0okRyLuYSLygB0Zis+h2T0l6P5kngItQo
GwYWxJo5zxQHT09MKk8BhGwwmXB0UQm+2+3Tqy5AGTZs8uagCwmTxMEr4lQmBsEX
znoYJquNw76eBqFifS6alu7ANWtp/h87q7r+4CYe8/WUpnL7UbNWDBicFa/9YlBB
jI5LTAdrMg/+K50hb+iML4cTfb/Vq1t2jIxZjq+eaiGyMNW+83IV1w13gPAGCZ3d
JUwoN91I5RXBuZwgCetW4OyocA4PtSUi7RWbIUA2vjim1fqQxc5hRema+h8mkmBq
d77vUfJMUUdOpu1RuE4w0dQMXpHd2yFk12fRpAM0CHkIPrF9SfCrTTbii4IoVIzA
Iv/dp0xwtbZkJ0f6jqJoM3HPtieYmCFhupiiTgSqq3mslViVNMuesayU3PjBPzOE
10ElLFjNPl+MS8w/gKe+XaoCkmKE4ffJP/cqWAOZnbI+JnJRzlTromijhw0rJ2g1
BXz860VbSN7SP2vO2rUshQR1k16+108NVKLBhR/x2TCiO/pM/27mHwaYuGh/1vop
GuLwKORLjX7FGXV0mtzt719lrrqwT9UyVlBkCh1MAId/kBiQT/pjSlErbm+klcX+
UelHyR9Kq+8RDzmoAd283r0NH7A0tHExOoGJY24ZMF11zTiyIbwbfIZMa9U0M87R
TiNC0UtrJUy7+NOlDUeF876NiFG18y64K0Y8406Q35D9UYQBQ8rgJOXjZsBiAUey
Wpe0NOE0MiwDNgWzxt0wFCAH1PBPhW1xXZTOMT2NFuQBi0eK3PLCkQtQjYELFOnG
KlEPZnPgT2fKa+CuFptnT/w7h0Tr/Q/ueh0yiECvJgsdZHsd4Fw50x1/YTjUz01b
4Y/U+95RjM5unT8xYkaJ5Be5WplkwX6mmXdOuWwz2gGizRjF+jG9Fb9XjeiRvQdG
Igi9JXfLz4yauTxzfT59gYOg0ctkET57T6m8MN5gYiGSb9l4fvhloCTNivV7kcZK
H3o685LQv9ELzg8CaQZQml6jqnWabpVX7rK7n+D2+022n5nGAketfCElCebxrQAc
Y1UQEqAmMKKrZHn2nE/TTRqkgBvS7h5i+wzXP6s1w721ijk0tWUicGgxPvMMupa6
UBD7sFsz5f9oVFiFzqZg1Ag4m8XaAkd9M3kC+QVYMRd17maegGejh0MmYXAtdS+G
Ods3a1o/UHs2q/v17DqWZJK1Toz/dIC5L2i+V/9e0pPZG7hzpAvjkddsD4CnvZTd
k53uDzJZAjSZZSmf4r/PV1KE+J9S1k2/0dgxTVwuV7OLNAprEnsw8++Cm0qiuiO/
BCQQ8eAWn1YpBJsxMnZkJ+UlTky9ONUR90gb+17R2ejaG3aCMKbD9vxER+DdZToP
fkVEQMFvJ1rN6JTjF7CVmQu/H1h3EkjOdlFHiXqSTAwY2QeQEVDspdtkfn4oyHml
qMsky+iUthtT4ScgkBXyUfSRtTjagXqpAR7DAA9flfdKxLvkFoy8KvU8uIRMVUF7
AP7NHKSfaIpo1ep8hEdhdKVXaJ7oRWrjUHWaKtibxf5iojFF/TqbD1X4B5EHhs5m
/1RSArt2ULJsSw78MvFMjicETjIRKEdWuu7NVhTShmCcBoyASzVm7oJtDpFnH5Ys
jz1rHZ2s26izU1TOJHO5T/4TB6EEhNFQDgwyerbPYRo3UjHcQn17yuXC+b/q4iaG
+ZKyXv/tKM0767wA8rViT3n/W5Fl+QxPiS19IcWkPU9ZfbOl1O0xS0/ovTgQlg09
PLxLgwPW3xPaa04JbDEB+XVpQ3S+BiIUq+hP+n2u796sAOuKyxx1dqw+lLAwxVXC
FzjhQK80rNdDGWJ9D63+a28moK53PWl12zvNd6E6Yzd3Qm0Kyq2lKl3OqNqBolqp
upfMYIy/cmILi4gn1sINtkDXtHtNNzRYxZG3/xSNtwKWmkxAilJsEYiRbrxy2p8C
NTnIOFb/imD6W3mCS+901KtrVQpCXkOkknR9DdjjdY2T//O6GB4MyPbrdacKF+Yp
Z+Y+6hoC5F9Evck2n2YxUKUTEIrNL2PUqrDdKVtlrT0NQkzTYB21j8kud8bzXmLT
iunx995BMom8oDI0XnzNQfTT/yTrPmwXb+TUzkZXmLxL3jBbLCklrchBOvXvsGgc
IIO1LnwXrQW4bsspi37OWkjtdG9ya3qGmd6Rh1uGdHOHRHpO668ZEwEevQHmTfRN
yLDkU2uPZiKFhaVptx1d683MMjHQGKW045p48QUg5UVZSAgnjArvHOYIW5GPKM5k
56xn1qR4NO19vVsDpv3fm5cmsgpwX+cfPYupCtzzxIPyeP9dYBlCOJ7wnn4gzEa6
HnLC02bH3iFqV6f0AYyOAWBtERc9BtgiqAoT9yevXkAh4pTjJtpuDo7XyyZumkWH
RgjkOrl3e+oWNKRdAFmj0BmRs3Vm74xIgeuZRVhbHYDfOZdMgJNsnnbURVdtKHbV
xKXLG+QLprZF6go7+t8aEkYWSKk0thbpO+Y4ptCpMKnsz38/mO1uzEjFGix1+2LG
nd5lfDe6y5rZSeTcJK/qFPOnmr1kcVL/DRUvVJ9deMV2dnmIEjviUXgvAKTDlAG8
GIYE3VEEMdfEcXPjBWOY5L0k93Yt+HghtpK0mihP3nMBfP06fIr9DDOBZonkNaF8
Ray0tszEvDgzsXOecUNh/LJexZUmpVAROMe2oQbiOdoUtWfrmvFwzkSSSmwSVFPr
8TdLnnjZFkElEtDJxMmi4HlzuA//V3wZVsuXxwJyLAW2WnY7butgtOjet3yoyxVR
iCzMI6EIIHVQGzxUXDgED58C+Q+JkeAAA2k4rau07Xp3hdqe6G25D3sh9JC6ONxY
2tQU7zVW6CUdq7LyvxJiBAkyeDoZybk0jpf8Gn6LX0qvoa3x368W0+VQREPG+SRd
0URM/sZR0+GgbvhI/BLWnCayhzg0yP9TaHIiGLmTv1zTt9GngezGvEE3IFWGJvva
//68Cb5ZRs+e4ynF6XxZlYR0O55aeiiSpb34OKhuCbr5q2erLCEWakfE8rcc2rdH
lQNh+Xng08xFjbdiV20Te5XALQxrdLCwYbHwcp+DPnf770FpnKYEvFY3Izl5W/Z7
g7qSOyWg3sqPiUUvxUTDSAPvE7wTh9a7krpSbP/Wa3NRmRC753g16z1HqmeJobxf
2V1uwulTl7krKBZvxRHCNOUPb5q98Ef/93WDRSkyzD5OFaV52mLTVHNelun8+YLG
p6cl2hXkgpAWmGfdPYOm6u6OjAVlX6u+5zZOHAm6TSb72H2PzWxVjWovgWIpD89Z
hC/hA+0+WlglGZXizV49qR5inMvFB0gSjknJzC77AQP6QbfJdeF3DLBizggTa99V
qq8cuFTLV/5BZSe0I6SO+Kq+x97AVvG5YSsnYehXsvoKdm8D3JZGavn56S1AIGvD
RL+bVxkgUHl61aS1wanbqJ+1X/djsxlu/HlmGBFYAaauF4KQ6UVv6QXocI4PYxbR
WsiT14klOcOX3siljMU+lUdxxQBQF5NxhxZnp/+SQjA=
`pragma protect end_protected
