// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ohbSC8PnpaHzt5yqcXncIRO+eB55tR/Q8Nw/gxJ9xEgcWyYbdiN8vTHSoVXx5Ll5
cv8bVqDvW5uyouSH0dMUYc/wOCbIYvfuIhVveXzVecLPEzOhUWCyfeOHnZn+rvkJ
jRNSYcH4YzkiPsdNEUf9uQdeLJE2xTd7pAog0raq5mI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 56800)
4GouKc612pjxXs7VLYgpfGQmv69o4dBwpw4E4rDT1ejvEHlNdu9PEolxFdSGkjAX
dlOK50h3hTTgOGG4bhOR6iebh3jBNZBnorTF1E+zSB4RQiLiPrYxd9kJiNvbtk4N
/Tam9FvravjJ5EkuuzYQNbP5UlaYhOTa+AN1HA9FIFrWyjBfsN13XaWChcZPtBzc
HHUdeeTecrp9kPXKJuiQtUsle5ChE3Y7GxGdex/E0gzexvJVXNjyTtXC9KAywq4q
hgE1fQGLHT+QvEiHI5kbq5a6QYqlmG0EIfKKH9JAqIqx3GxHs4YLurgn3YENWjyc
5eGzeWvOwDvhM1sc2fqhJpxzqLIR8qk46gLyCrBloKpkyZZ28jLToGT1ofmX7uYo
zisZH8jFcZm+/naVopgw+4HEU/sb6nNcds6v4zdk6c5zethuENs07PgRS5zuM4XE
mkwimmbYMY1lQY14u0GM0hcI/37RNwtlOBjI4kGrPKPgy2y+IaVgcnMGcYqyKD/j
GYogIFARp1yXVq91ZWGswmHgS6l2feL2HnEy2OXq00KXEUwRijmIu9uouhdEyTKS
PoDQtzCTohG4sIlNMWMt+HxlrJB7F9eXA3m5rHJeF+/538UvfNmMO/Zz+EZ8s5if
0OiSE5sxLZsgby2bbZKEa+VZzh86QuvzzqiO8uRFUmTA7vwV1Uly6X8LEZjxNku2
BaRLRYFUmjxjUX8aw24bQM1xtxNxJ2SQ7bTdwavTG7r8oIxx+xQplNNCmAqR4LOv
npk+Gw7/4PG8UjXt1q6aIb3W4aYrqv7pr6v6MPv2aFh9EF6rxWENtvodg9kIvEXH
MeA03FmXB3xzz/rkTOWDx0KwgraiV7BTd65SY2GUSSNT+s2+OsZcTp9eKqZC7FT8
yx7Q1LM+/ydnzvR969V+eaE9JVKV2Ls98ONwWcnPmuI9wo55SJAdOus35egWSdFk
t1L9eL9eLvAaxKGBd5UKhyXO1zgkrBmc+5wr15ehM5eYZ4koUicemGcqpJvt2+ia
hGjmGsJUAcgkRYNbnUEnBVy1l7aeWM0dUVM4HwCJ3Jjw/eeQwjarmHIKTvxsRwpK
i4RSxCnV90HgVEbSuqEt/pv6Pkf7lpepWbODz9opeuT9lYmyMkUW3YFwnKxdM8Jt
NtYVnq7gQKgEul7NNaG0i6jaj+HIYl8xfMPk5Qk+w2j07GmjwDzs2QWAafBTZcLG
jJZoojsI3f3S36UG2b9rtVWC25cUGQReGbn6Y97O/7jU6BKBYPMgmEjHv3iy0I+G
8DpgEQKPeQ8S2xlsiOmg2rZdDw0BE6BDRIg3KIGkJ1Ego8WbJ5xw5NkPj0VKKHiW
j9wrOva5B+zBWEz+NcY6sD6OLm7WYceuizQrwm9GwN1vthzN0jpOAxPfYdib3Q6B
8w4MDd+SVLIYpMVAQ8xw/B3y9k9EiLO8ndsdSp834Aa/j5pNICFVfXMvNZK/Lx3R
bsDHXZMP7Yw4Wg0ZRHs9bUokfOKcJeJx3ADK13S8hV3e1Cc28H3JkYCQGYccgbGs
5usi1hD+zCPvQ9w48nUIOVvIgO5oLAX63EdoH0GtYOsnRJLQ2iDuryn0hQcWAtA+
ghoX56xNkd32u7ZiH3TrJY+2dN4ATat/Z8CgoH8mrvP9S5wMYi15N1Ftq9n2sttN
QLvDmyqpJerRQOOkT8By9uPmTKpbyeoZFj7KItzdcmaouBDJpMikC/5qE7ohgQ7z
wIJxn1HQDcwoDHTRwMmCwW//zbGx9zMC4aPzVdcPv8VYz6gugJmVNTnetV09hdZr
7QxKYdm/CKwg+S1lvV8IDMV0OITpkRD436y8BBI6lLdJaP+vd5XprW0lR7QyfsDt
PFNg1Rtr0EHUkXcJOBEOenu4ICbFtDGCtpdm2FKkHXmDWq/2l2pbEkb3ULD7lwql
kag5NN4SAcFiwF3LryRW4eNuGAqZKU7MpAJ4Nkd8ynogyb3GYEV3fNgCQkMkAuSF
gluePlcOsS0LEpvZ0CEtqgeNezP0O3qUCKKE6i17HadroQdM7cztlVO9eMHNKgMq
ACQ1A3JRLav83jcj/YH5+7igL0GQvrtDV9Bly2GSxmhSyIO+vCYSmzdXzaWnZ9Fp
Cu28P2ny+wHZkJbzKkr+cmYtJkpgI1N3PP0rXG3gKn2M3O0p8OAdDJ1P2BEqoeL5
pi4G/8JAzzjq7RmE5Be9Ct3bPm1VOv6QnBvjaV1CWtO3CLHyunGkaVgJFcO1oMqi
SfjNw0brxl38hYesNgbF4F/SUy5l6U4z8NK11wbktYyX9hTMWK5CSgGUtw1SchzK
o3PU0ALDPB06DwLRQboy8Q2l9SgIgIeLln6Lou3Yi/VycqO7aBgxp3PvZRawqDh5
RRcKDwzDguCfgeyBMiOnQPR1R0uE6eo65MptYLW496mcdQjSB0tf0VIasxSYyPgZ
gxXdbgwM5v0Qvqaq/6vTzECEESEVGoI/Gx1K+5tNAc1fV52a1SWWjm1NBQQzijXR
EGN7AfuvVo0NGUrB6oyFagHNBX3JuL02dUPXK+NEDpVdHAz4H36GsH4pnoK2RXee
URkFOw9c07rPklFoPLvv4k2bFa7L1s/rMfcJ5MaXZVYs4rKB/BQ4CGJYYrUtqP2I
vheUEBwU3pf1WWZrEvVS+X8Tc9sJdXRWNSGowfdLTK1JI1bX9hp3By8l37m5IwGL
7yDiWkOroKgoFOB2gbpp+if+IrKvAkN3eBEDb+3URzV34QylMiTh4S72K+p0O9uv
GD54abkBQ/gUP3b1t08wV3ni5ttDfOCcVRofuQBsqA1pxd5jhH0TpWXyxsu+D90N
cRSSOHukPn71YprflvJNmRlAX7p8I/O9Tc/4PgOP/0qP7/cp6Uu5H48zfFH59XMf
HZKDXPZxYT2fL/gWrr8DlFqCnd1AgQJXT1sQyCBU8FQJhYFdM1Aptlrgt2/04Hcj
o7VHn5n1Z7yYII4enGzlows5fKWeumJSl0L9ZHrQTpSyXkaJsc+xzB+yEu4pAJTb
KS5f+lah3vlbu0PWYwEUwseiGMeRck8VM7e9+7y5dC1fyHUK4N5KFvZ1HdSl5JGS
7CsAnv2Z5rsYqGHdwTlNidOHuoD/70zzCYz5XGYdwb8ixWeK3ynWPmigIv+H7Af4
lzhFcLeRNgdfaTpS54ZyqRgewFB7Ynr0fTTCroYVXJ4n0xf/so5t2sRNggYuLjBc
yAl+e8a8TbIWxLxII0nyTmMmj76w2Zv1ITWanr5Qvo6nbJQZOAGTheBH9nbStoBJ
RXjd0gzGZNm3g6SByXFCme1H3dRnnK69EouOxiUmkX2q72wkYC3MX4WPQJuEkmkL
00xTivrMEQEoqm9Y0/qWX4XI2QIB8Nf/CE3RU+olFJas8UmWe8Z7Qa7u7mdMrDrC
6ZGTq7wOAIzmERgmksXhbZoQyTi4o6N7wS2eY7Pc4EB2Dp19nectG/SeIXTNYX05
nO2Tc4iPP6q2O3ZPYMOXDdKL5NEPZf7hf8ZNjCL64V9Jh4S9GU/GqcrLnvDCYl+n
OnIEFmfpQU/fstvc3Sg3uBuWI9iOOhsP7Uwmd7TJmp9AtX8KoMOSs7LCzqUcM6wl
I3mKymtpJYFrFHbwFq4ieqg023RoVQhxYYEpmrbUxrSwU4s5G6Xwnsnfmv8etHOL
XUwocfHDNiX6MHCmAIlQX2/KsnmaQqwJC97hodaOPg3pJYartTn4Gs+a9W9Pw6wq
GjkMP7ggbJxqrZfG4DV5IFBpekJmNb6bQLlk6do0gOHAunDKsLAx2dN9YrgJr8sB
UxUwoV1wrC4AznJZ/7Gryk4SQgAp/itafPp8W+f1f7akCFoXkwsmwT90qMkCok9m
ZhR7m3E60MrzGgSTAdW+AjMQI7mO0AEhZ7GcJxcdFK62cx/la65f/6GYeEP2k8eY
kpqwj2SFajRMhfh7vCXcBZ+gtYLwyjFazwmdNUPBQG69PVuurTR9p26aHLzDq7CV
zdwInfC92ag8DqXAImZW6hGZsOP2p7ngGx9bBhPGOtiVD2xkjcKMiN1krYFnSKpb
9ln6WixciHq/3DemFV7Vs459LSfTyUg/DIrxGNdAP8i8lZWK712P3nXtWJo8hHJk
1C4mMruGpnMT0vFM0HcAq4wLecBeOV0g7ESmvCWQWFAiH2U8s+IfMFLE07f9+Hvo
zrbJkBlluF/c/dhRWLxw/3Zt+waifAa66w6DSUzN42d4LYWxrTmpQ8BlX/Qm32TJ
0EoSCZIkR1qBtj9E93KhsWUZxBFzqO/lA/8W/4OsdajjtBE3N3BEB+SsJ5W6LlLW
3FGPaprZ6RIix+JeWGbgk3z7Li6oNkKLeJMP9k6/oY4aTvsS2SktUARL+iTcbiT4
uOPKJEQKxiANxtc+BuOltkW9J9x7W57pTBnTONYNRQ69HLRQMGtOdXncYGAsgY6B
bJkXnc3VYe3WJAhx/pFkVzHb1wRXccQCVRy02gEKaqol8kblLcbFVc7vG7ZNNyCK
yfE76k5FDo6zHehCIitIRDtexq7GdiIqzuJBFPLoq6CQJa4TfVXFQy/X4RBzf5sl
ZY755DFO+AEq96TP29ZkgdPAg71L80F+zY4aFBp+vn6We72wKXCZ40lS7mg6nTTE
XYLpjdmENadhmlEg/dQi5xjTdxQuamMUU9etEpDikYrhaK+PMK2fY3kbWrsGC2Wi
+twIt33KQNAb4HUCrFb0Kl0Vk6Et0BjfmcF4PWsKWIDyAk6MQIv0vzKb/zOFaz2N
5vkiqBuEmM3E1S0tPWCX2RzHNo8MM6eUd/358hFQ6hxOx093JcSkUW0C8wS7k8Ax
v6NB7Cq7Z+63rQo8Uk+WdS0sSJScMFZYTapmiGthBZXjVkrv2511tuBwOaeSS3hv
N4g5JGMeP388Ak1gKnf0ohZToOI/OcPZ+mAyXINam/RclZXwK3G9Nahk6I1jFRrj
QdEGx9ZQnr1N9ikFobQfg35wl9LOgLUvhdXeqQMiVpc+r6WXkCpxXvv13Ze5VQ4B
TzCAQvk/Kl4UqRNk8UUyBxy+o/GMKVC5dzwo9asTkzAdyzQKUo14PuUK2hTpVwLl
J68k7ykI/9oUvrCM4nBGJ0VbYZRXKUH3oc1WtNr40va0+TGEHwrKDurwkItujhY8
lZjSI+pjYJA57FizfiAwoInpQOy9B+W1SbVEXWcngYrQe4tcNnQp3j8KHZHJUmXm
onGXspb8GRe4UhVRD/IMz8SjUReqH0AzQSY6wdvFIjwy9NtmZK8WktOfrHNkHvL6
KgJvQ7QHoksojuHLxDDBD2N2BtsZRPk0KCMy1OU8GDRNdT80CI/7wcJkSQ4s6Cwf
I0pttkza+F106wdbDEGHso0pXDKxrs7esHYUOrpWhJACQk9zpizadCH960FHEXNX
ry7PtAO1UzKb3QoA/X0woHR18Pkb21hMzSI6qiNeYy22Y4i0c6fG8qvmc/SVLGg1
ID0iEY8UFBDXFWa8egc7ia3kzUJVFXNm60XkDjBS28+tCZlytuUmISVQu//5TnwF
XA6MV6Gg0x95Vupivg4OgQTBODQDM6nHTqiykGNb/jmI6vJCdSo+9mbPrDFUyBTX
nk/6hImO36QDXWgktrWt8txWOMuzgXOjkV8IhtJzGPljSr/BsYUqgLQT70SrlTTW
ws/mUCvBTCqc9/ZodW3CGAB9dk3k4cM5Tu15maKZ9ypnYLzlrObDoEcuQC1Ue1iW
W4Ba3hI6CsXONm8MDFBBbdAaDDHK5GqGD2+w7PtxQUsSZO4pb8Q2DBrXNvcRVq5F
MFRHiiEuYdY5AALM/G79SVOIhc0xCals75kADyzdPw+h19RHLmfVut/kXrtQK/b/
ED8A8pDgnNRfIxUZt/QLXqEUPfQWFhXP5IkYNfFaUQTu+tKs+0N7wRYl6Y/BvcTA
/+qJrC4kwmFJN5Vgh9s8Um5jVYbr45PKj3Z9zocXJDgo+imiDZ26PlDl/n2qFcV+
6n5P+YchUq5JolWW8h/EcaIMXIlDELu/zaoLQzUgwjmMRKJHKamCB3ffcHHh+1sS
dFSpcUUaEqaPKutTc4Rl7YmC7gEfNE/1qoLdrwfVTv075zJkRzDv/F5hgAzvm0Sh
8Mludi1PfaapNdteE1fykB0dpwd8JlXGxPzzsoB9U8qs0y3SHaUy76/Rv7SCfAQd
mpgxpSjbQqcdbZEroWIQNfeA+ANy/OIlD56iKy2AEFPV6/93BZS8dyUwqrrjl93K
SzVGdYGUWfipfBrW4kiEY2/PCfCAk1z6gUv+WVpjEFRvQ2a4NBWSW49Ff2JGgGuh
qpl9wDno88WTbOAie3ArJNO2WX38BrylhJkPAt23IpHY76IB8XV5muJBNiz+whF2
chhu32zziSKLrT1hnxakWTlQWWI7PXd9KrJ98z50qvJ63q1ZjKOCWPwwVcKAlkyx
sNAxY8OMryhivA0ZL3YQpXAVsGH3l8A/cnQkIgCFK2SHkjsjixEb3HUxc0RENIW7
Vh2Rirhi9OgyA6vp0LXUPZg37GovNZij0Qr/k4xb6zKi8Tibh2zFriPI+y2cCSpH
HTnhmjwA1q5Bcs/hYNPo1k9zyGfIZV4XjATx9p68ggacBZWClajm23te+tiUNDqb
JO+NPFMKUa3bK1qI+XKRI7KqS9+wN5E70orgnHapTXM2FhjWaceQG4ucfvHddoXi
EZ7KgeB7JVPQxKe/ToTfOu1ZbPruNpOsjYqkH3TO8+FhIWa4MqDaBy0nHAPlh7BZ
gs9Hgz3rzzwr/La021gdDjtSCADK+rNgP8uRK3rQ1IM+NBUTxOFtzKJ9s548TMXp
mGtupL0n+7jBrDpL/od0E0XgbJH7KoMTuKTNCU2Y/M9MDqK7465zVcMPHTQenfLi
KKwOLp4TBB7af+ojVIb2Krfy3WHi6ZkFCjIAV1JLYUHkrgd9ysAgj/OrsHFRpbHJ
DWcV/AxT6saTmW4GNZ+Qe5ZuZvzOB5+oOvUM39bH36NDf8iGIUmmzGiIQgWWrOMw
S1mk58jtw+TxohGc476OIQW+nUTlwNeFk0QvcBkdYYdMIahwAIpf7CIkpSL8vOKL
twD83akhPrHLaGYOJ//hhgrZeZe7fAelW0JmFWh89HgFA14cN1ab9WlJUmkI6LAK
OvuUxZEjzx9/KWiyuuw+bxcbL+KHa0q+2UeKFKuyCYakGeMidg99lcMS6/wpghuB
JnqJ7DHnbUs5pgRaTofJUtpKcytCG3a5ebcGMski4kGQverGaqQNGjyt8e3F28K3
Vewmo3hrJOo1+E5SH/klrb2Y9mpxOOH0kBMSSuEL59Ach2ioEnwCm3u7ons9QQHU
VzKr/DWNwwT9qEQKU18xn8BQ3o2zXxhOEO0zWY+fgjd1+lVNZUYHMEs2k2dGwrIu
mA49ximlmQSQ1azTysVo2yFZBz7llxz4N5WqH7Byf5Iqh+LMY6cQQgDRYrqLuxsG
NmLpoFqags1MLqMpbqt+CGofYDaM4kRPE07irD91Y+frzvK68PAhL0V4LDz3/92o
mjqYiEvkaAEaRsIW5LUOr/eLqEGJb5ec05aDbTXlDhXMPGXkQ+9dmD6o36kWlehh
KFwn2a2zViUYS/gF046d/eMhZka0yswcCEZ8FvxusHR5QcR12ODPAeAbxGZxxobD
+Qhh6OdXJ/lE2kdGjgUEpUl9lfg5fdW6p/to8AB+a4+OZ6b3Y9ZC9fy+CbdrlVLx
cA0mWTQzUfmZDxX4wMlFssXPVtJznd5C7YgRuErG8if+k+FXLhkTs0G55DPrvQ5j
c8L2ED+0Grt9XrCrI1UkqPW/koidSMvqoEqZ/9GpZj4z0xvoKXYrP6UqFTDVv9ua
SDOroW8nxf2UOxtE/fddYWKJ3iXpn5UVE+0OGy0ql7tHHCDbgQgooOz9Y0uNLByX
UWA/DMMiHLjCBR9qiSbZ534raaM3I9fA3TQuMBG3lQE3zrbI1BApUW+rdgRvOvct
uxSydcZWyVB5b43xkc1+cuC35wmFnTFEzJ4ucsXfuNG0YGfJY/gDDpfWg1sEYvEr
O9vpuTiQOIMAdajX/nsQpX3Ov+KZjuS/C5Os3n1xi4bqvcHYA/Yn7ciQNa08gRUu
6jBCP931mBnQIXS1OSwWoEIJj3O5hsTK3jf88pCeHBncIeTW56Ibgi/SJZxmzTNP
lEWsGc50izBqybtsIM5O4pcUUVsju/7GbMnfvfJMn/HhLlYg9+Cmgx7lLCaGTpHG
gp3o41S5SllGh/o8tV1lhgb3L5/yXjInjGW+pxg1p9i3K/RX1veQZCWGpuyudZPc
UeTh4jT0nkHrlep4Tp0guyC+DGT6BkzI6I6549wj6yFw2wSrlLdM8guB8XdJeQea
2j1PyPYqrFIjNR8+wF24zCaqq09rS04/9ote6fh/WpKt/5i0YVqMxSIvfWgix21W
6cPwk/jXVbDtv3pR7knwpQY344ZdlXGEuH8VA7FAnvS35boNtSmmAvLIV4xfaX4V
2b3oLgbbs728A5phHc3FVBO/pvM5wBrAt6fVFQAgr2vOUf8OzhjasP8lIjIZtWFe
k1xHSJCHWzMiC7Q8RvWtzcVopp3Vhe/nkx7BDaszb25itnqkym46TwhxRiPcaBra
GprcLvdvRTWLRG5/FGmMUL/8+mscoVLHH1DpcuA8HDdzjTAjIx5l5KbC62phsS+R
cgyN7ty2Sf5I10aHwSa5d7YeaJ755hepaqFAR28QePgF95Fv2a4wayK7KFarVJaH
48v33LX7rRd+ukhgqQEGGPs+JchZzXPQ6P455Lq7HfDSmWJhOTUzP5o4dL7xRxzr
5bj0en++/E//nO/mPRVWOt2MG31gMhkbZYUbIXxyfFT7Vqhg964orwOPP9BveGfl
Ycwerq/vFsifHl7LksYcj1bsqTyygoLvmp2LyHeIGMjUvdHC/OI3Gy2M2eTjfurT
oabRxN0Wnalq8cQD0kL5GX1CtZNXSDnnTIs2OatBW5ZJ8mN8EFM2oE0j2xNGc4Zb
QHJi3/QEULZlhmsE4PWLpz6c/OEhLqCGaE+qudSJGPvCSbaE28FuyyOxieslq3Jt
ewoVGEdMNbzWiXWsqgbfSenzhunRhzwWYJWf8kOCaGlaS6fMQIrLjXavE83nAn/W
z9KRSc0Ic0tW17UZSdUykksgcGaF9nwBgTSrQduYTIk23a/08Rvmpx1RLVFVQ+1r
PmY9NMJlAoasxLAVZN/GkYlg+w5jzAL+oKfp9hUGjhEA6im0X5QHmlfw6W4qCQmI
XYxF6xCTF3q5goq02KoqKIZ2osZT1MGLQ7b2OH8lomMjSUgVwoy1vQV5LcBEqdxX
5ioqCUOQAVr8f/Dh6QRm9j1G9LaLCzlKb7QB+s8+10fZCKZCxyb8ogmZ5kvZAgH3
H7rvm/3kg5KxJd+khzLd4OhPCDN2lmudm5qLtEuSoUznzKa849liJyZhYuP9qvh7
4p1tKQ5yjHuaAuL0vFRqMNTPIP4HZ/L4EgOz4HFk6uW0Ws/X9vgd1GJNUiQhCJKp
PVcQo+frA74lBvYUpU1JIfTY1rbXA5QUIfbFEF8pMgyybthpJ6MwDV6MxH0KXsPu
hNsgx/A/kqNsle148MVr7n8rh9gUb/t75NX4YBvAzKFQEwCHtUO/FqpDy1jEL6rV
D6BjEonu2nK6dNdV2y/aAG3zIfeOqmKcYgOiOM4g+z5UjROzipzUERS6r0qRGZyE
4OPw8Q6/v7yDGTt7xRjFNYIK84tO0KtQDIzDwO8yeP+cByeHx3L98t2rjFGWvXxd
GedHuCNVEKS/f1+M1311/dutySYO38b8dOn2Maw+P3ZKQQpGG/e6IXwYf8uEekV4
B5gHvcPKf72TYKazxJDfkIcbc4ZxQ4s+kIlMflK6eyVIb0OvpVgVd+SZ5U+NVVT4
KzE3TqJUf61bjfs12/fHHzF2+f2iYPmxwCFzVee/Fh4+HeI7n334H9f3V9NCHfUc
qhmCNj00UkU11/JxOHN92hmvHbPOSoypSipJmx/w4379Aae5mhH58ADfXGBu3PWS
4GKJzNnf8s6DhtUh03jBywPVO3pkcDdYb04ChUL1kSFwUQR8OEj1x1f/GaT63Afw
T/z0i8Y7NUwG2i6NtVqjVz2yjpJoV63UU5EPOCnUAFCJovpRzFyY9c9JgX7ROYcY
Kq/ryGRp3fJQYHU/HPC/D134xNBSzc8A8Hj3Wj6NLBGmnnrin9A3qinI7ONsR/Rd
Eo0O2H75mDREoP8h4pv5m9CjR8hBHOS/5Wejl/CmSofoBcIvNVNhPBmueD4yiiyu
1ls6Tyc2z+7vbSQ7OOO6Tn4iGbkzTbXNhLEo6A+Fbl//7WEphtt2vw9CJphiRONz
/0N7rf+MlFYq2DKwVa2ePgInmYMreiGwV+dF2xM7h2thb0eugsu6ZCZB3NPDxNBH
2ZA59I0A/xL1DPnBOvLeSaLh8IXrbaaeUes0s6Tt5G0Z9hvj47Rl49EWDk7PMSyj
MKdp+9qJ4zK+H0X1w/rp9w1qnEnqK+qsP04E6MHCFYiL1hZ4YjmtEBbG4znINOTB
XZOru/vhTt/IHTYetSa0lfIPbdRA5oQeA79V8qVrR5/oqHbKgaoECPCVedFhhpDT
MX6WVtUxQfUH0HGq71l7kpVKrebY/rLWc2nSKt4L76sj/bPytmGKwEqrEZHfvtr1
hiOJ4frl+56RtUR3FCDrsjpr66LOpzPe2IsdO68zZf9W9IoEB7VVdJlry3ATryLN
rTqaY0aZSA2gDyrMBr9//HDxmKbIWgUzcYADSfSxDq5MVKbFj1Px76/usp6Xvzr4
p0RRG/El3mm6gqmDxdCoLgcpVzcsGWLtv8vHikbZt0RjYnevW/LneScH3thf8hf4
hEQFra1rdalxXUSj/9B2qAlzxhCqazimtA8iA82qrJLb1mj0y3I6nFHdasYUIhc5
XQDpi9XXiD66S7HMRj60wo9CoNsijZKmfoJ5Jwj7fOuCAZ9ar0GOvKfyq8/xL8t5
r/18K1sC4Czea/exKFQTmAdd58UAFEgzS2D4W0AKdphMRsA0CdASwoqBZk+0bOtu
ZvsBDFj/NyFZI/mZsKwCX/rKXn0VmdCzzBUVe7lbHMISJTdP6xy+uPeXJDstJmsv
zmYXfRFVoi3JEuARwyJ+W6BCFUnWPOiaHkFTXcWwlVDBR0c+kvOutpIisyyaw5b+
lwdMMvcfKFUx7evq0YeaVtVd1PSpRhDS9VCnMlFUSNyKCKnaeJgeDBVYRhNVYY6k
ym/6JyBipqLDGQKB/zZqKEd/GVzyS8Acf0tD9Dxl9z5aNRj/nSUl/rWlXWPqC59W
tfEu5aGS4j8355jzgymt723p7Sy2D4XwNY8zJP3a9/Ut0n7AwBx+rtNksdACBkv/
p0u3ga0NRYKcpWTUwSQ1KO16n9xA/TjF3IcAu60/eAg88ugJBasm73t1qibMN6eK
PmHnD2tJh/a+OYyEio42+B0iNjWz/nGtD7rWWS4/sDb629NcNXpi/MF11CrteVoX
eE5XWbc/PY/slbgksbujEoBEVAh0mdPQ8A9QkC1pepYaT7DjBf/eMN17+Z96OwlU
HmIDEJgiB83FhhghcNjuuN0CdR258Vqw/3GnW+ikmztBjo8aW2WO5kDTlh6Ox1CY
7IIJaK9h6/eJc5KyD1w0rj7RMajVtbLkleIEInyKIzBVkL5QfxQsAZ+7R9a2jfm/
xja5w/319Z2cOrjx+xdXzr4lUE6NmQnp8qf0Ky/KAjda9K8XwStjbjCwTmH/4q5d
NvbUxo4lJ6o/BaZQunVDgSw3wiUuFVFtzka1WlpgM4qqfX8DFrXMMtqgmZLmab2V
OjteuERl2LhsvRJkchcHMzR3W64+epg7NjzYFn95mcMdxy/caEyhWCWSBTEuA2RR
OAMXgmDQbZJ6xHHJOgUTpWGeQRdqy6xnLdB/09siMv1NUZqwk8qffxJXHpk2NQy4
2X6cPKul5VzjreK+FPubFLjbwuBffHMU9TvnZukYhgfyQSACOee5RjL/hQwyTIt/
hkFbgkKY21jxTcb6dHRkm5eZdUWEyVhhdyn/oeNLNu6WEivLGgdDeJqzm9QXKPAr
+iOXOMXIzAk0CjqAemAKNoJ23UW+/DJWZgVuaV5e26oBoGaRTAmL9WeS5HezojYB
xJI6zeniWCgAxmbLcCAoSYiWeOyfj7Lc90FOeMvrdJjsHQ3E+3Ma4QUcSBEVbBCk
4VszaSld2Pc5GaVZRq2t1zxuMJLTVZvnEtN2racR8VTOvDC88gUDVoZwixJSYC8t
ewA7xpTnstLzLToQrZdbOhcWmJDK1aFPougDLYqlVloNmWzWmcxiSlyqW94Wm90d
trA4/ZKOHUt99bG1ZgSkAxSyXvlMcvRTeMXi0E/tGcsbpeHrHzkOuQZc7pHJW+Vm
VtGKuFH5Lhnl9Ka/ZtfeE+DRtAISbsH93GpgCVzQzFvRCwpcxAM/Wgs+I7tvodoS
xoS6WCCfejCdXlk+7yy7mMQ9PCYHTuNX0G5YARDIjyC5UiFbPpcV1XvMkyWSO34o
720ZB/28aaDnnki6RVidYJ/hPBaUjyXQsZAYCDCq81Fjwlf4d4xZrqMuUAlUg6fD
jF0iP/sjfExyikSHgTmNza97oxE51QmIaLPD7ccmmZGoqN8eUbBZCq8+2H3YW3FO
D16eGGrYGKdWwJc8+3fJWSs6aHsmRxrQYETNeEByNnpy4OIxTJTq/DJu4Ivu/i5V
bE5PElUozO6WOTlLGnZQzVwPZ1JvYsC8EWeDUBqlnhD/6UelnwpJh97Vz/i2DwBz
LmE6SqBKGgnhoP2dLAFqTS00ai6tZKWuZM5D2VjgoawS4MCgsS/xAU3GudVhiCHf
oQdJhjNJ25oyQOA8YgGgu59WPwjMy4+9MJEZOW3ARah+epG1SRGEYxHP/G2cg8O7
oS18Nv6oWgFHMNQaMTMH056lPLiIc4XXcYbN1QZRqzWd2UbeTiACiD9Yo3BioVbW
VXqlO5UyThy90tRrA/cQf/nHwPl+/JTYyVnEjuXGtzogkax2o9boAYPjXCn5Nw7i
Twq/b6xiDDTqAgfskJJooY962Wxip5i89b2X8by3dWGzdxl0FDP23iNlDXVA072c
Q974lVWs04fdUhiTeVcmPjhWf+htdcBzoEhGrXNOFeIDyzoagOlJctwgmOP2MZZ9
Xjmm1JKsKzGqvz1R9Nz8ddzTEiTAh/YdLC4QMYr54Fpa2e9ft+RSxqXTDBPG7reK
8wudvoYDS/ByUnKDG6sS9cfQtvvQUXtD+0cJEzxVf5eYoKIH5YNYTlfmzxCJthze
U/eID23HP3D5z+DRR4dvlQrcM3GezbYirK6Ao1RruvOc+u5mrvAIVplGlxItZH7q
6p1QYtrE59E8FQ4kXi1XbF8JVzxIC9Derep5/EYTqgaf0EgkXFQ+3mA/2yCvVBoD
/vqRy/RNXUd3SeYhAQuavR0bRQDCFmzWG3xp5sfvcR6NfjssMJnafv3TtxSUpui/
c812yb5jM0yXTjlIL7P6VbZNnyA+WKSMBzlGXfnBtw0+oitTRwUGvuEPWoI1U3cT
Ctk6uFeGAm9ffQY4zRcYqx6GU/MnNDeQxH9OQi+CwZ10MKezdS+uZhG0PlMW8MZW
kSYRRFfh4qN1rrd/tFfT0MrIDJDsjT6j5ikqM46Cs9vdrs89s2dmePH7dc3IHHVU
xD70IfuPtjT+8Z/JoOhHEBzofgyvYBh15GQ0UWqNfoma0gEl9pT/9BPGvOY2RFAU
zUOgWtgBaO7qyvZRzb/lDTIPP6eMt7CBu8VQNoWZm1GzhBjGlpZZCCMt0rO8LkIz
Y5dfH6PXU8bhc6LwQexlUdu+N4lzYOV+dhVniqAS+7PE8338XaLdG6bK8YTwgzlF
aYG/Tecba0GGo3oHvj1hGo+TcQAvJ4kp1s2t/wJyIEcUXEHDtylAmaaoARB+g3jy
N1ZlumY/DVOd79S9iFH2dFLTnPH1E2Btb2l0pGyqjpyQ4hmnxcgPCGaPo4IUWlOn
gBlwXV0GuS7pJmvjRE0oY9i7csi1OIaYqMxZ+L2yKD/eHQDmtd+okdXUSmVCC36V
zPwV8w+cLZZQHvbnu8pulI5bBk6WDQFIRN4lQSyj+FgEsf5HKN4yqA8r4PwJ4w+k
8bRIt7HwIfFTRBAj5AQpEfUcv4dlg5o+VCkUJOvvViiuvWOa92r/fQhjd/VvigBb
/b6psUyqkaI/p5Lxx6GPbgASxhjonEOSzMjMCJDxUDUSayiCRXpg5RPKSQbFeqBR
TwprPTvioPE6jZDmPYBQRSzdVVx5P7NO2LGV3ESjrRJboFEztindv68j3yVOFCpf
DhQ6knvOy07xODrsYi1tK3nqgdK4HzFGp0+M0EsEffN6Isth27QoTLVM7rc7nwgj
B0Uqcve3HvGr69BdTpp1rfGgXPdacf3NjPnbnym+S9gw/P8uSVlBUAXPc+ffv2KK
LR91pONFkro8cRzUK1qi0dEclkTen6PVtk3Zoj7B027SiAxdVv9h2ImTW0QCaT6m
ZsADdAHwcoDRq2sauepuYwpuogeT5B58UJP3y5HZcf5k1nkmfLsFGcITQT2rzQfO
XC6wiqPbOnnhb9o0+qdTIFugyd7pADhHT4zQoV79j1tMIy0G0Q+9MMdwZ6GqjfyM
FlRK5F6QHjFNsMgVXO10EaorQA26y859JaDa/JzzSBkcNGg+I767ngrlIrOpkrBe
UTt+9PFBU407DkZSAnG/uKOT1SOZBiJYVsqaYCm42PoLZwHXB1fgElWctkB30Wr7
h4agvnPCLYUBvGwwOvKKk+fp1m3m5/tc/Xc2Bm+l5Ok7xHEsnsCPrPSz3pOJ2Qfp
H0CRUQW+Dwk/9V4zD9vFC7jVaU3AOa5Y246peZVKYiEtxeaVdQfTL2fPut8D3V2/
ns+oGuPp5C8zaOTImn900VdNtD4LiFfSMQgDz5+K2iUq+bgM8Eg4WsnKArVjE2Wc
YifX13w1oxv/DV7cXbIqhM6d1b0DaGS1nXGg64mJrW92Cd9wOXqfoWTlnXIWvJrW
D34iivd5Uvox10gFev7A3tHc1nvRr0sTUthnPx4lXQyb1CCYuDrCxv/3Neq910FP
sMdqwUp4/x7S7MI54Dr0kdSK2ffbxTw02haSG9jBKGUy5x8ZbiSg7OHc1vlh9QUw
QToYG9o3H3rC6PbpOrK7KHccDzeZlr+R+tp9UWQ/IWdU/obt7d6sEOombytHSFjI
Y5HQV475TZ+fcBWs3JoGgTWo8pG1IgR36TzIipSECIbp1+odsae6A5ZNYTihvxxO
Fmt4iA2TBdwRKBj+2oHA5FQG8BSI//Ji8Xyll2meTFlmndSLJM3wqRD4YumJXEFV
8EIEOxLyZGwpmAD6u1kieaB0sKrCK2+DwQaPdnsaT5BszxE3Wy6j0mgsyjA4cdy+
7I+rJxAV57f/oOJ946uFHPDDYa771TjiwwdZuNjxLqrfPn8poI9HemZIvQHjePRY
dnqmlnjslWN326WcNUx63+TVDDq5xKh+k61hGbJ5I/p7DfC0FVWOQEgrShYC0sJg
3Zv++mXc9O0C8oqO/bYPs/92RUWPkMAg2SMRQaCr0kOXxyVnHXJ9Q7y5anD07wa9
VhdlSuqXNFCZE0kjivKC0jEhTxsAzsussdw0Vv1LfXyHn9o5yRJ8sarSC1Mwix/o
BfU6K5YQ5uh7UT0+klNmzwwqQ8gN/zSyaXRh5D099mZOq+cDmpi0FaBm5//0fs9q
WlIlRKpcxKKByRD5RJXPPsNxMWlMKpc9kaaJdTTEjTsMbMyFe3U6SYmKUOJv11nh
/S89oscJqd0prMd4OfsOpTTkdPM+/NOFVChXtMHzLwNxuILfoS6uaS+3naaEO7EX
j6N3yeI2lTFoY9eTbEiYsQVEf3sKCaO7tElP/EDkSFVU1/InoupMA8cYJilC7l8F
ZSOHnq66gkqY2IGp0/XsyTld6VepOAIjx7n4daDouoxNWZkJy1GufnEw5Hio8dCR
mnNp72z7KVO8B2nxUUH22NOyW+SCvKiXTf51a2KG76neuQYENUI7/ocgkq9QzvcO
AHVT3ClsDNSHjRRIy0TsQDxSsjjze/IRnvHDbjbY/YDw46cxIpeeaEi0xOgomzYu
3EWq4bL/LAVcqYgDvBEb7uQ7pJrT0Ywc4P1PHwOxEblXTEputxydx5BZWjHNe6jz
IYXbNaCsIXbh1X7Jn95qtfmWIWFwEeYoQRzqt3IlaPGgZvTER29lJR7XDvEyfJ6V
stYTk5oh/piW7yogE9TeyVytnvFRE89d3Zy0DVCpuajsoWJLcMQqOLTOv+ao2Gao
AtV82i+lm3qpuiQ3pwNnUTnhK14hFrrhYSMTnTercl24R0uV9qLDvM2UxIMSvV6D
xdHf3IqLsof5UrZAdLmHXj7lKG9CQUJZiECHtbe032fTMQyo/oTvsWesttm/wb2u
hEyszvftADjMFhcJ4I5vMuGaO3Gd1AYQnIx8SDjBMmbPO/L8BxlVzamvsqunMkQQ
mP/6TRfWL4qk5poSogDP6SF/xmEfGp1C/a2UOKJMhMW0eFlMDIUi3E63VyaNss18
Jirg+P+2lctqpjrnKsDDktqynUnTrRKP0vg4zR65FHWy/p5dYLNREngYUKZVMf27
ZZZISvrNHxnerqD59BcuRrSdtZTRAx5PZ+iaTClT79mPZh+opxOco+hEgoESC6oa
2GxcQ/wc1CIqHhyZcHRsbyagjNu8zKqnr+3BTcag3n5y0U2hylEs1I3S22kGhPHX
PR/HfykqMQbBDFzpV3WiFWYMBx9o9XqK08Skg8bvOziOIsFLSZ7sQJOvj6fKfv42
zL7oOeYTEkfoIkk2L+HVeoiMEUtnBhn8WZwo9LAERjfEiDK726FhTCPxGbudovbs
VeM0eQqQAoplqEo4ZUXnwiTqCZd0GyCfLHnSG860kyRyDo+/rZAd0ntgrm/lAtYa
ayejcdYy7uBXX16n41gn7azAOIFL2Hz0eYPuiUJv/e2j16X0R0soyMXHxK48EzI3
0+n8a1mFVASGFHQ7JHsmNvQfoUjhQCMg3cqLFWJEt4opzQWOGOuYSflUT7OZdfVF
GBJmCpaAM5WVf4O5YTlr/ehYvWbx2tviC/vIR4pdubYrRXe8mRmARQnYqcp++T6z
sczB3Y5UHHcit+Cad5nPsLVWlTjgf9iLDVXehj1ku8Ejyox54aqB1kNk5hj82m4S
0RL+NQvT8yqrPPyM6OPOPcMBYtTPToKPQfAzm+eIL/uIeGU9voaHgPjBTENLF6yU
Zi8AyPwJGCRlp15ySDW7CcrnTl32t8eKA81K+WC4lVlLfTtjNyT5ZNYxFGwsARkP
GEc1G9vWkwuGnHwiJtIyqxXxEZnFZE+t4ieTYrZ1e7jf8FYodwW9bZDPkduMFcbG
PT3XIeWp5b0cWYqZTF84i+7BdINzfllmVktfdiVsn7dg50nQU+B/+S88VONQ+3av
lO1zNwt5dNo/kulyEAvJ0Vt0NhZcOuY+lPNhMlOOOnvtlxAD78zD2+LH1ceDcZYy
+cFxYk0RfABP8DfB7N5g2QpbNjw56zXiGskxYHeFtktaQaZRlgaqMl8jt0AzRB43
ZNsUnYGr/9eMpHEpQW/s0Pw92y0Cs/wPsFtOh/HR9CbKLf0FutgWHard5yC3fHTm
Dnu12ZdwmJzjoilAsROCgGO22I/POxpdqFpnTj2CyUA+CS6A+TPSuvWy9EtDvi7j
neX0BwSCvNhWiwdHSWlLkgwSbVeLHTq5NsMnLh7WJ70SLNcqB553/sx6NFWJ6mSX
TGVRUI8NbHw5Ftx/T0gbHltgtXsgQt+7lXvTLTe8WxaJqwr51nYuXvzbBKBFwBy7
GY/LILqNpcqDi6OK+dxdqefXJAc3UtFVhiV9aHfbmC3ATgMNX+ssPlNzVrGXAhhy
8tLz+TV2TqCducPfCGk+oVjpFDNcfoIzI/VdqLSFhr1U8L8dpzPNte/+z0ZZortM
9sUHiVNmNWLlbkaK/Qe2sWXAp5g0ZckuJpgKZOY3lwLA8+XlsAWP9a5l4g23Xxoh
6zQU8GuUSPyzYNn4O6WNIJgtiSigUuNCQDl3mdLhzQX8soGwjxQxQzwqWWeYAIt0
vv1kHk7t/e0cSRaJEe+IcTYNZf4eAPJlooNXk9ytSEjwkTg5It9HbwS77lhWEtpX
8wNNV6baYlLUZXMypvy5HqmRyGzcPt3Mc3bSZdzRppxFY4OVXqxPdX//8nH/gVwD
2ECH/JTDOobqFCz9yFdQKAWMOwY+N6IEBSA/kZLfnuDU3sp/04mVoPVr3xJxmYrG
XAt5ueCY0z7yaKr76SC/Onqn2wbiI+VqjvuVWVWspPl0WNO8/ESyaCUWkBFYB3AP
pPcocOeo0pelCTgZPWUo2IVcfNXjvkhDqkVbhwfigzLnxIDOkgY6pyqTF90Cibec
S8NnoJJvcVC9xdP7ttnT10jPD0F4fNSH7S0CzEd49Myan90oP+UjfhhnxsdsJT8c
Pl1TzP/jrCvMWFjLynYkduNJO9UwmgUmb51Vs6hpjdK1bNPqI9K2GG/wI0x/5Icb
iG8YsbqFcEAc2OuAbszryLbdNyvXKSDzU1TVvvEyvVcDQWcnlcxfTw+EhTaYQLTv
35bEm4dlWLcT7rfUEVdhshr/QMekFI4pEbL9En7hUifXKeEtUSEDBHapNoDcw1Wu
y8zC81BUmUVrBdtV7BR8vPg4XP16IMgMWjCXZSnvS4XHLbIK3vKIUoKxiU1TD8UH
8VroAdY9p+p7YQh0s3icN/CkzH46vF7w2Sq5Q4e3HmkPJmcnZHgqx2Hqx7G31xBA
GP3h5db5k1oC5IFuJBZPu1ezGdpDtAcoKGyWNKxyuAw050UN8JEI1Gcv0NrFUXW8
7b16r15dlu+xeydSUC91Q6HptL7zaahRxFIzjOsBjr4hWIz8n/hWI8S5vaB5/r+Y
TRVO0OcA+ODRqlkCX1fSutbKXuIQlmT91Lix1MiZUJDUTIGNJUwYN7LE+BBcS88x
sikTgSobw8lQnET5cigt/ZaQp18e/XouV16DkjY+q++d8rOJnvvX9VEA952X/2gJ
QGoNqYurp6xQuqkGHDbNTJsSQo1v0CxST5l/2xtbm+8hxpdE6Jbc3FtkiY/KeE60
BKUOw9s+7w+/sBSq1wmAWHtN/ZiD+JyyCSywZRazcEUw6ZrvTTc9Xxj11rkSKO65
sAXgHfGV2qRTS6gCaVB6w6i6p85+jyLBsxbM3r3ef4PnDlOM9kYY9UivH+nCq5AB
iwDcchx36CPXEqvXqiEvW83NGfpSWZpWryjqL1Eqam0gM/YPLyg5MgTN1JOkm3Nl
1+lRXXUcGN80bqmiYzlOifAxwYp8F53HprJTKC0MA9AxWWrMRHeESZKeWYJf/ZXe
wnokAm4MUgmvALNXywiY4TD5b68hi5Q1xyw3nxRIGI212/EO1IXkXmAZTS4n+yZB
PnXlrJDR3c3ztcKgqPJJaoa1KD6725XlVXci88V52CO5hdQvAt0Vl4zrvRTNeaE8
TcuIALS+8kMP8W0/qiPGdNk90H4ZNsB6Uu2OPJwo28eyqzo1jif8FTki4hcoXUuE
eIfvTtpxQ+MCrR2GML0LAgb9clmlD1yuG56hFEmM8d7L3NtAoOQnzkwGvDlei0zP
sb3PnH3e7BT/jEaSiZBnL9QMGzS7Se3tcGdgTm+R3n+grrSnFRZPl4Chta3yhB0R
vG679D/8/Ljzv4hn5sdGCwKjLujJ+GQT9jYxy5tvoQwO56xKmD3Y5l25ZQcFWQ8z
rJFMUeZjoT/COqqnjx4DkEsBiJi8EyjRv5CyKdJ+mSstPcbB836PmvEbfLvyVlmL
cCeCPOtTk60KaCD1k4dPDScEV4rZW8V6V6txZHixYJepes3uP6/9Ur7HXRmPKQ5C
2H8Ygqn+c2PJyJCGNZL45aa66N8xM58OiR25ZvMqA/5d+aUEhHiHrLv3FqLLEWsn
UIk6TQ5loMkojxwcxv48WTkHObv3ccHFF2ponEd87XZKoLEHUT2TUrbLNgcPWbqG
olpWDwDAL8ONv2Ra2hbgVAqFiIyHVzzRXqHFP/yF+iPGJTjEEpUwDHEmJ6q8qe5V
BLvY/nf78z6V4SqRAx5OjYp61OVFKe2GJpo0VWcWQAXd1zs3momLGx8GwFQozbyO
3qqle73Pvqd65Dc5DHsYyiGSyCS5ieAsPs7z3cL7oUHaFyb8gFxSZHO1pgWdrzT2
Cp06vrCk/w30cviUjwXBeCi0NUPIe0xX2Aj83Y3m9G9Z1oFtuThYTHpi0BYLPZPA
6y9Th9BbccrrxRBEJ2mjrav03be/s1UKiHfT7LuseRLlTOoIy5NyE49yVcOPALsY
EMkdwi1oKegM93JPTo7o0XdmfCZJ2m6qRoGPJ9BpzBC0R+ReYy3Y0KxA/JWlrWMx
D8YRLN2wCBBX/oIeW8bBz2EqW+PHlbOb90+fA2XsL0dFtBipM/yo6CcetjozA8Wn
mKrXp+fB+++HjTeX7IPgyvOfjl16ARiRILSNakL+oRQnahCr27wR1VI4YrfKul73
nmc+UsiGLfbErRzPJ0ZHTSdNAG1YoSwstcBBIklXTzbtEVBQ4oqteOIe22a/4ovw
hD1/zC5H/budkxbaCbNwmpY6sb39wNUT4X3K2qVKFy2/OzSYP692E0WrbAN9uL3f
8YZfLMyQn4hA6pyuFeX3NBSVJQ+bxr/sOY5j0uq321HZdekEZdjQpRGYx8PewNWI
Bb4hEDRdfJUQCNYj2LZw7ff+eyvMgCk4GP27YKg0S53DRI9a6YlkIdaGbUhDjVoe
h/nxRn1OSP5NWEQXG9aOq2RP44i46ZSqzBwFTriuSQZf055RampUsBV0iYQkaDTF
tWC/ZKpLUvwtJG0S6wu2za3blMJ8C35eKenzYzb2bjJ8Wy5+K4wtFWCz8AXysiQ/
tBeovjKoe7u5kqB6idK+0mJ4PTrr9/OgwTNPXr63fNdOqooIonrnHxjgX2XOoD33
t2mnfwVA6ILM/BXLKl9h0TT93WvgajwUSCq3vp/b04gPSQMVA4V3/1TPl/T0xaGG
ut4sfqy5sKxc9XSJSWyV6UvMvLMrWkKznGcKHMn4SEavT6TGPTQilYTEQJmBZHIW
im4Iq8HeLRw7Hf3H1+0ZzQnmi63+ySnwfWH0VkGark1ENwK8Qo5W3VFl+UwMnH4q
n7B88sxe0Jfd2Gw8h9D7oI+CV1K+PxD9u6/kk69kYvfSxV29ivY2pY42mGSDYD6z
+jHDDV+9J7zh0xh/6lAst+O8RYGbyGflo3OFr/g1Wjxa74CgwzPYon+N9OL1BF6K
clyAzWfY3B7JkTLGxRn4Aia9u/TnhcuWWV+g9Q8z18EUFpIsWN/OXzI1gmqXION/
Nv+F/kPJZt+D0qN5LhNIHwL32siRI3lgBq9vKWmfd5I3VNAh4L7YLXPpkQLAOpaf
JhpWO5wiG433G57dOPzDAZu23M49pZ1KIo+OP5QZ+a1odQItZxQoWzkX1t2/xChA
+1LU4ajEBWbU+U8sDdamy4ifwk2Dqd1BFqpBEE5frNHlWLKNFOIQYuZzP6PrDR3u
smYRqHNslrWv1Okd4h9bT74WcJu4dlr9oFF0ip8MDs9veRWoe5vj4sq9XPtwP0xe
bX6lRdQommRGpPGwthVlGZEqht7QDDMa4YSzUjG63W26PbS03dM/aVX2w0s3L9tr
ICSRE4cagdzvRVgZC6buQKlOIyxBHK+fq5alYKFS6qkLz51EIuqGufnYorbGxrHl
2vKfEdrWCtgnd3PsSAtrHPNGsLc9TYBBMarRB09utY9HPvnKbt1mywuBnsJ8LrEv
/Vqkx8j/ldFEVhKn7aMWa9yKm4luVHPKRlyb/f6kn4wnbsGYsKnWVFEVvvjt0IXF
tnaUVVrC3D6QtgQRciQ1CkybxtsQi494xEUAZAPGtZ3GlFBYq1xNsgzwgixaNGrq
5FevKnp4JibiQpG4l8w/0Mo+b90oTQwNiv8/UufDThy4Z5OZrSzdzz6P0XTzzIG9
MgWlULenYUhmVjpKg2mzpUSnv0M6eSaEB1rFS615qOZV18swimgXaIyC+5WnmfAo
ReYB5z7HdA7eMLv2Qo6D6NtTaauUI9b0SwqyQUnql+JkaVjRkrKzosN4dm7wwNeC
1OxHrcUz1bcyhNckpwFlCGsRKCjAN/n3EYXqHSIZnYlwuSBThLQYiJ8qsV3AGzdj
alz++PZH1PUOijHD3/r+GMO+noyo1tduneHWtxrTgM4QnRCtE5jXPFOUh+YpHjAW
EXBEcSbePqZ051DwwWsKMIzAeTSoj7RjD6FGk4NmwCbRCGnXaMYwfRIJI+sKGd67
ks6qUXdIkN2QHQ60qTDqOpD7s9001AtwMcW1zBXopnkki8SpAfn3cMMQ47z00IQV
lr6v3vSw+iW0qtT5qJr9k64zZJVierONfsUqL1jmrLNCpjex4ZQnJn4XaajyrNfV
sbKOR12JUTZ8JvpE37aAhH4E4T8X/pVw38njDuYKJ6w71lNlZhy201mIURRBv0S8
pxfpQ93mzrjgCOI0lpnjUb4IUlu9sL5TUMEjKj5UfoobPFoEc3d0XxGsTzpWuskj
/vPzWnV3HQGTCExXPhO3796l1lw3FLchFMYedZ/gbMq7BppHoG1xuO0dfGuKQz7j
/LUtiASDoH8d9KQvyftuwcm1YB/3o1pumhI1X4mcL0ZMfte71PGXy2+4eFQlDpRO
+X6J6mYOnr3+u90qvkQDWL7YXKwio5nj6/nEkX18DOtcwXg30el/2/SzL03rIr/r
ekVQwRsyrC/Ezkf72PIDGv8dycwv42rGPumJ6meRK2O43z9rr3PH33XJgoBW8A0i
VXDg1IkI2E/55QuTRcMbvSO6GlTyXzw/v1zCrCvCTEwVne0QeqIaJv/2EuAssjDj
jEXHb8ualFCmHr71ykKBSS9o4q5IPvo2O9q5lnOQMZN2+soA5CUhgzBk4WfqlLbv
sNKYiE4AIuzZgGrq6Rz/397Y7ewnH8+yW2d37AQUFxMgVauekx69qyAOr21RpNRs
tiTEIzox1KByyu7eNNHeZDxVOAEzfekQCR9JoTHUZKm/PDKIPbJaJ1NPWMt6FJZk
ZBUWPXAjTIq4NEqGPGnM8p8cJVbUiZsnnH2Hp+gNdjyWlr+N4NhKz+qDVAw7cjEq
OwSq97/Psdy33ufFxPXl1I/SHZJz2OSwwHX9SQoXLVrYO5t7kc8FZ3UvFq24koKf
Mk/8Zju1Yc6158XHMY9D0HihOxGl+5f05LLD5VynGp/UdEl57uSu7Ao7B+PGGzMN
35plo5eIC3EUIecC/Izn5W8qGCvZj2yeDTmze/axYnVhyG5A+E5cX5qcgdqVJ8k6
XI4vTBcdA52ECw6DTsub4Q++KzIRFKuxuRovXNyTnAOPrJk1vxVym/5sWNxScLcE
jp/V2oiAxgmUHN0Ta5uQ6BVXksHCk4dpYqwynpAI+XLNL0Y1To8i9xD6eq0Bt6PK
1yuipjbk35qEuSgmo9CuURs7Kb4ydf3bSJhpoGvnBgGVJgmyp5ZzTtTSTNUiqQZo
lTVlczcUrPBoWsQ43RIUZ+gMFXsx70xKPVjHbaveH+GldRjw9LrBcib2MNrdPmaR
/vu4QMVJjl5EFcvd+PbkYxykKQTQmpWuuIgdtCHETUThfXzbMq8eeJu66+4lq+z1
XIJcURHJApUaBqNmVT0cxWstplc9POk4/gVhodtJaK9sP/BWZW1kJyjMI302Z987
Ba98MC8xPS0KA+GhQlZSlXnvhfHqgSmNPdetl8nnO09s7RBqCEDwRdngCR8AY0o9
EwTys/ldApWc2iKJotDl7C987DHDwoOpZNmQYvT3Uxex9YhpwElU70JsgFV/Chs0
+F/X4PVKfBELxXoqalhaXbCb6Q2zHyPnZH7Lc4bOH4JR78P8/FiZQ62pdXf4piG2
R2XbFG/aYpfxQ5wXg65k81UfBdnvAWsesoCLXpgl6BPnP8f3+9LhbrvZ6j5upckv
tYwKhfz9xQwISOC6RJxgzM0sAGnlsKFpcano0WzgmxJes3yXPm6tdjue3y9r0fyK
efZrEhuXgkgUn1+ch2m0VuEWJfDA0GCQtifqdsLhmlhIzOVhOI2kUEO3ezzdxhxY
3keQG5QZeT7T6HPCcwbX7sSekgyJ2m47R/zB29HvLUrPcxwIiUIda1/zQrLTWx6s
FrJEFqPQgbVDHMTMkG2zMZAlvdG2tgUhYTl69Sbj1khNHCZA/TsaWbe7cbQIhjOs
LQ0KdnGC9Lyj5Xzx7n0ZMww90APbbwpMrwzc4QSlkmh8bEvELCD3GaSlCIqcswPV
VoPi9WbWWIR+66MrB6QSS3xTZZNrC6lDwhtL2yo69KI8ktX4RdqbOByjoLCoOyLl
N8rv+StT+/nDLr8IPd5OK1XcgX7JNoDTBfqRyWsjsgeDaGra6pkab9oLg8FWke/Y
3KPvCPUHZK8JrIv8HuP4Ix3HzZ1k0C05ltmvir4SZBgySKjFJHchLblPHmOMNsNs
vEIn96m6vhkP5crVt/V5QyK33yC9gF4p+FL8YEynWUVGwukNaxE6UrsQZCAc5Nca
nOHF/CIn+f/qeqUASJXUAQn+EVP96YxBaxMoe0x6766OUuWoO+5bvRHYiUhFdt01
GAkH7rOUxR7vIvvPPsFA6zHckDf3WsOIPprFEJas/tnFtnhVjwKUKvqGY0to/rpn
h/lBLsqt5da/bQsbXGLYncQzmGvw9GgouvsdpKXnpDY21ihIPHr2ozJDOSppwrJz
anUACLeUrHuJwPdK4/RFOP1hb2vHloxtF0U/xJ4F0jlUF26qQd7oM1IijfYPNE1s
xKjFIqj1a+1Lz1SU/Jl0+RJ28cu8WEZgpdaLDrXzdrQLbYqgOaGzLeXv8f99fxr4
Utd+xENHmihrLWCkb1XkUpMS9kxcqEUAnuSw+olCYdnPGR0xYZn1WNvqZ8NEXxwz
Zb6Su9eleR8yV38/Iuf0k19N7MyGIwB+oP+bFPYQ9YD+5TQ5e6jZrWk+GPWFXeii
DZVUQG+b3BXqMpu+hefttakkaz8ocqBg5HCQ7Xq6yU3CfwBLSNI7pv+5w/O6o2yZ
5m1evQoURdf72kwkjanqQ93QhV3YcgAgC6DEuQPDwutjAr9e8QUEEftvAiBAzFlS
Zr/rpR1P6DlfTnkgaQB0qDg5d3sT5VwlqbZ263IXDe8nxKigWEDl7KznMXJIWRev
wGPtCLNWz2QYApKbsEYsBoFi1aiXfrgR8XNW/742MfUn5Nj79Pa2bCJlZgb9ddKC
Bdao3HCE8V0g1Ab/Q14FAdn4kZ/hkzAA4It3LCH3jQXqsOdSToSMGJ6c17h8e1PR
No3F04i6SY8LfRgi0NgDJadAAe24Ljc2Ro0qxGWkY/65OozqmSsDIsxhr0a5UqUw
/ITzHJTlC2Gjv0vLiOMhjWsrK0MjymbGXq7+eWsXOl0yoD4WzaFRgD5LAjuqWxDp
MshOgwsF5alvuZSMgFm01XNg1H6DMgYZWr5S5WxgFaCr5g/PQL6p2Jf2TFNAw+S9
slzMZLC+iBnscdmyGmIxFqFWWnoQRBL2FJn6BKu5Jfc5u4uN5rQTen3V2siMoR6/
mamFaSQflVXyU/5jO3+BL3RIjpIXA4RlDaWzVQpoGO32VdjaLpRziQ1x4JQ1m0q+
OXtLSKXgk1iopGl9E36ZeD1CsomBTZ+byoQ7REg4qafzy+J+47CvmKCvKO+Tlrl9
BoJNHBnaokSkaTyxvwWNToq1NOpez9U7qP4lIhiLUrsk0Z8S59xZ760NUQNoBnb4
8EECnWgRnH4xl3e0b+IFIQAFLYgn1m+mL5YTJP3ngH8ZCxF/PhYsuWuE9YyY8+xM
ENY9Mgfge932wQCrfQMQV20u3pdRUa0bdK4P5P45X+ikHmxGqGJ3EW0wwbkK3Sj1
IJ57i9FqiHQiqrjidrG30mZQzCrqpelorU606yXvk6pgawbaN85WCHulV/AQh+DF
rZL3xmzGqRs0+tFvyq44Wj2GbEfCLT7A3ITQKd/ke8MBFMSOvQ3K4bw3F3/xmQR/
8OPjkAghsXRCvyc6iE3HJRzi6P+EIfgyPBRWmiWWY57NdTCc0ordgy7DdyEXrlsu
sOy6V6MVkuYMorNl0n6puLXX4YWRLs1JlxLHuwg1zeeCsG0OUp/9JN3qXeJEPDOi
xIexU7tpdFfbK+i93bdYlbd6+rWFQGv9VGoG/+bO9Mo3e8ap2wZyMqJ1h482eBMF
v4KLssaPdCpswdu2C9UiL8mf/vGzhHjDlYxmLBnAYAu5DpeD7vwKO4bo70JB0VH4
vfQZOhaY06W5kfqTh1mZV3n/HGjnd1Wh4KtLoy8McgR5tmk5Pyv7B54dwGiqgZ4f
/Keuyhax3v+bP6EVTXN3LwEFgoenPKGbCXXCpr4HAUSiOanL2Trs2W2vDXlhWCPs
qZ5uq13ErpMygBEaZWtssOjlH19a0KhNapWLxcFAqxLztOYf2BRqVwsZCjQ071ck
fSgJiZHkwfeRLhlX8zFjujGjBophnN2PNpcE7jXS2tYIB6X7wLmdlMAN7fro0G8N
NDY2qsufNIyCr+iKE5sMVu3BwkYzGLns8bt00TEtmucUxkSOiuP4jMWveTHjVUAK
AcQ/lxQfsmqfCSiVjeumTv5RDdRw4faP/9mHHifx2qTeqfCEoaGlkmOA9lBYvpza
eZKrn9CO4HCGY7uZjvGZ4BnNeVScV8gwtNNaCFUYMfnVd35uDjxw0Gx5SqN6FNFH
QAViUORT7OmtchPDUsSrVDij3tCfKoZBqMt+tx6i8Z7X1Vv4MSt/wkbU7mNIRBAs
GsIfrJ87D1dECyFRertztyvglHX9ZdSZHI+Bp36OGORpXfU43at5P9KqLPBEKPQi
ZnFuKI8ZdXvp4kTpNW9vieXq1gJLRGvddmg9ynR4iM975HDfiG80/bLgg2NiHGAB
cB9orcTMopl5Rbdgc6lbJqyxX1fl3i///legxZZsE3xomZ4rsv9W743og1++pLpK
mwa37KLYcy708QyjDMEQ7568bsSMQ/WBCYA7/juyOujnKLvhgDst3R58RhAF8//S
ISjJ1NnUofRe0OqMjco91Fik/yN9tWpvMbeknvPDigKAIOBogXGncV+M8xy5A9hS
8ZrmjK2w19rGlEUIyD0Ni5jnyoxGMa5kAPEAYvf595cvXnIlL07ILnmbaF5tIg2c
f57UwSJyEf0ityccoFdqFnb7XlSmKUzbA8fL0kn1uAR5XPVTkQEGsn2wWvjyzve9
gVw4O0pbsVWJBpKhqr50tKEd2+j+ly1Fk4CayBVF7NNMUXqu0Yf9xNw0B/7ontLW
Z8VKNU9ziKu/Oxl/xQ0nJ3ELfGtcMJbvVLlS8g4MsNC5nHQSAqX2ly95LA8+zJE7
PdEY2YSYSMDaEr5eaarL3lsF3X2CnYtdtiLDuub9dEjCBCM52k4YCRhF3af68322
+To5ctxm3xGdW6saf7pthUEsCpyoLgfKKQBDavbN3EMSuozr2bJdSU9Bb5riZwCw
QoVhBEfZXIiTP8l4ItOOWIBx78zR+I4hXcgZHG/dJuYrvvjjRlQv6Fpl+rUE5Wpm
zNgoiigub3cyFgWQ+Y/yZof6uFj0emvdi2oR2I5J9jwQlcNX5LNLfFj1DwFRVeVl
FjN42zda6yemh/JLlIvOwU/AW+4pRr0wp/dppwKKwqLGlytmS0i9r1M93aVQA9vz
WYolsNcLohYF7soASxzoX3d1dQ4vtXB6AqqGJLM3dkEUmGBNKaAiB4awyVR9/KRH
3cdjFc/YZfLmbaK81HkCh0gP9RLusIbo1Iw8vfh22q1ndVVQDGuCvx09nYhNOKTO
d+jtAVZUKrrixA0rxQw279lT52aPKKQTDqQwXmN/5zIaOrl2POkeyxXPL3Kei08d
rggkzbtFp14mibJRoJ4m6VOLqJT+LQgeZ+o/Tk40m/D5q2u3msNqsDuwBwz6hBFh
VRnQPXeMBGVPENaXvb8uRg9QPO2MPEeeq4vl5CHZtlTeZt07eNMPxP483pdM/WgC
N1ioWdEm8ckFjo7yDV4U1HzzuyN/pay8cTVg3ZJJ+foCGtPd1KUhzGKBHuVU8+s8
6LrumPWwP+DdNVPre9AzPIsBGnP/D5LqSQ63blJM5zG5c4PM8smoWzYUgCp00tRW
+ydonXnjpw2z10pEal5BrEKyI3e7kUfDEyAuBK9pFPSoP3owEKxtUtx0i9SWZQhY
/vVvZ9oQMR1wzDYbvbRE/6Ey3nYMAiLS+ohzWVLqm8tBn2IaabbOb9U/jLBKmu9I
lihYYYTWNukAbqQHSPS9T6411HQYyXiROmBLhGjcoRicjDpO3oLpSyiox9it/5Xb
TsgL/ght2bG1gR8cf8FrZ4Yfs8hTUGAMBaRwECVclFHOTxExp7yzuIgGd/LazUur
sBCWdV8LXpXtA5qLlkIRBSnySo4lxsF4YF0jFczQ17qtPiVEqpNfboSS9UyfjtaR
/S5M2K/IXz8TqDL7SehSW4ocUsAQ527n3QJiVOfd0zw91N9T2MfERj8Q32DcECBb
MwP8d1xvUzvAZjKNJ5cPdV3RzFqHgEZcbE8cY5adKwoDn6gWzCpjodJ8f6rUNkSQ
+/zPj2aLQQkEvr2HYCfCu9oMPQhYttqojLqcdCufhEJWRSFgjlRl1TE7xxELayPH
bfqlM4LIIeYncJd4ZpnY6GBO0N//U2PU9dXCIIX4OYKdEGXgAOygU8VbkVsgBnxc
tm2SFcigZOBSXgYcF1tJJWoAUwCIRJ/PoIyaXY2jm8UQJ75Z6I+7kI8zrm3aceGz
+guGy/HvRPg2BO4G5nxBWseIlf840LTuUJ4Bp7ja0CWnvxK7VEv+JGxvxr/B9Kvc
72n6imid5YzR4Sr+ALvuqsoXkf5msJNY/4jMOWA8G4EVrzqgHRfRtaLQRAdXS+yi
ErmX1W7RXbC9t1/Hrk4hq6TMXKsLx11UX3zlJFY/QyVZZV8jBUqxJcMtfC4cX9DV
h8+KMZQQvzSl92q7CUjylyiQC9b0Q5H2hFgiloPPebSQzVmdq5XeHvtBHoS/BuKN
uSHjD6cC3VtSE2pTBXUyHRa4Q32INzitJlIu8HJ2ISNt07SWRiVToOPhxBktGPa/
JUYQOAZ4uAZiW7h4Id2sED+Bnt6icGZAm1iAW9ccHlDmNx8wz9ycRDHcg+EqxHcm
M9+ZXwk8J2Vmtjo7QeCw2yYkY9+7tFt74+1tC5UjO7HY5LJPc+6+6jjhi7EjMdCD
hRetXJM2BxVZk7hGFdS1P+GYzNQ1RAFRsyod5Vxos/9xjJzsK2BahUzOB178cFJo
+zprgThrZzrSuEJt5vJu/Lv2+6wSGxfQII8TVH36okBGed5ykpqTrDrWVI/pnmML
6RHK7NyloqhlhEIWSoyFDwIRsQMV7Kajc0OYosOilpT0FdsqgcqtpCCBbICi5Ghy
awE1IcQx+OSBv3H1SMtA564mX3Q0vnGQcaJM5tbqH6uO/Cg6zieE1F523HU/qgrL
CcOaAdTnbDwZP7EZ5eOgDzkHCSBoLOJQmxYp5p7T3AAab0drVw9tOOgHRAt7hVPJ
T9DT0FBz/G1p/siajPDwiiE1WT8KQwvuvswIJHP5jNowRN+C/wC8y1nzhAtXd2Jq
XYj9IKG1ypWoiPCD6b7QMhyynzEo5Ahtk7HPQrOrlC+FdiRx+Vd90TxTFVLX+Rjr
XFP/joOI/AAkeO2IQEnEz+4m1yiXhSRSwsslWSRlwd2bey3uopk/w58dsXTPnFp5
67E6hIj81BcHGkq3Dc5mfD6eLpx/81WssEheZiNIpNMzCWAePm+UNgZPn/VC4t6o
En2B796yqCXMFnnZAV1KgcMJ8OVpfEwD9xmblM0SBeYU23SLwyUoCvLBkHaAiCfY
+P6ZsL/lB+ChSUxEKgcCLUOCPTGl5xSiapmbEneOAQ/2WCnAiY9Fw8+j5DwYHJUR
jJWAZIYSeWua6mkZW62gWLbBTOy0c4icAEV4g1zFPPwwUvhnIx/Qr9AsWI4cmFM+
yrKiSrRcW33SIwLMW7OQ6dOoPRSeGgouNIkjbPaKWbrJinPNfWq07RisuE1+UnBq
eOSBptbJhBkvfuOUEqKdGbIQ01eht4jkXdO8ad93lv8Xo4zA7x3+LEcTp/BH6XH0
cXNHl0sJ8HyarrDRf4F4cb/3Lv2beUX1Waj42U54kaNXfJZEtY+Oq1CI8pYQDEr5
/1k/GWZFmBzrLlqDd3p2c5+l3OvEfvQLx3ndxzXKHmEyJwg2/kl62LrwmZGqB2Ie
Y4kYGM+qflx6ZBEvfXv1RrDGMuB55ubfTLfwoAhCYU4GNnyAP+dAHmSI14GnaGhN
QdKgwLstI9FAMmxAYHEMfaNgLc0Yy4N3JXZ9fn2s4kvXuR5tJAIbIkIGQLcEKu5c
IdmtxWbkzqm7ubKQJ7dwyLg/Gzt4GcltislBwhzn/O7kn8wJ8a+Hq0I6iQNb2O+e
gxjW48Vlqh8P0X9RjTnw389QXRR0AXjF+Mfs73kMyDWcx3qSLYuSYCjoDHj9dJH1
mkhiRN0QzCFtuq1zNrzaDdy3NRgrlE1ZeyPhcdxTeFwinPTxeB89QEHnS5sk8jdm
ngOqXZN+2N41L78DbdElMlOFws0hFAzrEMNmrKd9ajRP/Uhtz4sY1kl/yrw/5StB
fyDncJdxQscVb1K35ZXbuXihJ9iBWuHhhiGrtDO8+wGcqKj8iTh2Mmta2UlukXV+
NKqcxOteKX8ECUIh95U1d52fI9shvAFSr+oCu8MYtRdlXqS+BYE9nfm/h7mPkB5k
WhymO/93EAVJwSa/90OemICHP4uG3rWJtScq18bpzUfFr/aiE2hK2nPMvPnhLhSr
76LnJsrPLVlU8VDL/PdS83dhEASVJ4CzmqK4cphPf5f+ie/86eradDJoKO8hOzig
OxyCOGRQVHwcKcQ+YBjv5K6+AxxL+yjrP816NioYSl4Ll5c6/GZ21YNaDZFZA9LF
h2woAFQkcLJWGnY3njiLp1fiUPzRcD2q1qevu3QEj+Or43493FkS5aEqKvowqhqN
1nt++yBJtsxYHe4VkhBgQqO8LwLjeBLM6ZXfDw4uh8w60cNUlkP33851GPbSZzli
w59KWImNvzsYbuKwJRQ9/PMrkvDxxyOB3CvySzwvH6ZDbyGCgzDaaFbAWRh1vVcs
uYn9gv089rGByHxocXZoDi/65dPSq8g7H04uAslC3nmT3FNHC5TyDWpf5GXfmKjO
eMms1TPTF4V25FtANj+P2/M4uCrcflsh3Ce11LKzwOSqdRtM72NMBdDMBnKMcZs2
96dL34Kn8a6d6Vb4tHnwdSomgguYJ305UtzLyI60B1VycDQR98fnJCb/OIoBbYrv
vfNyljETMhvxUTADITwXSAeojP1iBRCA1m2FkqnshOopP3joaE3rpgTxtSPI5m0T
0K2y40OvFVrXwF4sSP08AFlcR7teByT9bx7YumaHXHkPLAnUGMBcT5QBQZZ0zlXK
m26/yiRf3I9pgbHNh+E9oeiBrHt8G6DBeD47kT2E7aHtr040e15VvCVU2MTsJtJr
f2MtOVPip11ETpNQoqQ5TTUXbCXz69QYBe+RNA01O0BQ/LHpfVf1ZT6GfwZys/4I
GTM+VUzikPUmQsLahFdg7jaqaQIFxxhx+HNKoW/wKRV1K1dQbG0gJwzcau2IDFRd
e1WYxlDUHck5EcjT2fhXMONUblELUNmZV0P2XwMY1820G0RYu4tqJ65HCctjwRsy
vGNMHN3/5l9EkOlHP/xco6SZFUADJSQLxrsoLuD75OVa2Rn9KdSNwhWJD6C2h6WD
seuKGk1EeJVMV0h2qRq4ogzG0XmHwN++OvC2DIf3RhF7mTxt2HbChEoNnCEGSMMM
s+UiTbe4T8qw2V5/kUaqMi5KYQEl0AKA2J+AQwSB35jVkFlaIHfGGBUu88rgmntX
zKIWwHPcczAdyBYBu88LjCwmED7eks1XNa4xBx1H1BYvZNmFODczdwKUhFvnBAe+
2rFy//xfuCUSiCU0PlhQ2LO5HOUPqYJ1RVRE8J+YWmOPLqvzsPO+tD/fGU1faVmS
XmjcTF6RaFyxhG6jyXb4vFamdzMOBotwHTqV0skMkLI/ZsjqEI35qH7goC64SATl
dy8yyOwwyi3QolfHwlx0YxipNUkxs0LwytoxG+9VJloOIPqvajB4KYLw0S9uWamt
TUGXZ56Hdgo06XZ1FwtOeSjnm9hSyFBwaWjone5VLxJZ22btPajjpcGmvkRMhPRJ
pysSG6maj+0P4dXWmLT2RO/UfNNIPzev0pCVaV/lPUETfth6gKWqNozCXmS+LIWt
stxKQhXDFcO3wyW4dhZJ0G4MoIWQwAThtl2w9UIQLrP3qiJ/ioPlyc3XICAei/RD
oUWFr4omaiXHXDQQtSPYIasCXSlm7p887GL2dDkKEcXsblqmMt9yWQiDXYnYAl1M
VyR5GlHxbdB4buQCwfcUIIPCh/AaWu7PF8NStELqKfaLmnAa1ST0uCBWrQ+wKh3k
ZoUGRQigt4zRwZ4IEjHQvAFFLQBHfjCneF5nE36f3mBFGo64FTDt3uBk9+mlnPLj
jh8pPB9HrNSd24OIpnEgMnq5FwZDD7cS21MQGu3LTVEPcQBnCwEr4fsuPjc6af1R
hvHp8foJ+f/x6ARuczmlu56nBjFYuTL2/4QBwqvmQR/CU/j994tESdDrBPkRldbP
TVmX0DycU0SXnIYV/O4cIk+u9mMqr0alTuDKIHE3pZSfeUEeuMjRKNfIRt/fvCbR
NzcNApw5e3DEq9hEZXPCOJWsF7PqaKK8cPdLEwacr+GpJ9Ewf+M2J/Lo4H/g9uU4
iRr4VNm1pjdUp7ce8tdzr2zl+9nzBvzqwh11QsPKDTq/l4Qhg/3RFs6lCWFaEVJf
EmHp0xAedMC5mqEMtbfyUXXVnhrALAd9UNQ1x36KELMRZsToghXiX1OwMVvI0RRy
mhBIIMRt753txaM4jQ1Iakx0aiBn1RUZqGHX0Qtks9HU2ZBBuhWS7zw2sJRmGjyU
HSdns1KgIEbGn+qGX5DZCW3lls1/r6C3Kce4i6S6xdVl/97MxuEXuHzcWJdTHk8C
HNphtnLQ13mUAkoiu2t22mgjW4NEMoZRy/8G+otNP0h70YTbT5QG22H2eDmzvTY7
ZELbniLTyr0N9i+txTEfhYc5ax0VNjw9ILlUVJ4D2P5CWuZ45bRkxy0Sgt0yFw2A
xRcoVFPCmUIN+zfWLiXRGkX1KbpBboIg404pi8c6/2klUcRThxnhu6ImqbsOw1HV
GrnL/QqsGXo/VA/VX7PaaCLlxwy5y00CBIPbiPLkMAVQmiZAs4IdFnQOgVpjG9uq
V56neOPf41edg3pTAsCRkPahiurluscR8VH31b0FiRyKXyBbnZ0FxrJ0PFpE1Rpy
dtCeMHTOzX2jgEkvUL4Rw1jqW5hC/EeXdbmowtS6dOrbR+FfajRdWNlolYZdlES3
r22dde3b+mTBEOb9y0897bm5HJBEJymf48ORnTV5Kd/Ev5eo6ZjO4+EG+22hhAKI
7JL2ikyVtD9X9Rc5fssmogJp2LOJPcPIiwBluU4MmHzaMLVzQj12k8oEcv4UX15K
ltcp48n4YNsnHOF5kS49KzC0ZEPNe1REKXVbKMIv3EoxnhNFzUA3UvqxoAPNhNzD
jai5bm5uwq2wxrOg0091KmJ27Aptzy5P9GIPLkmf8Sy1ElImS5OxsVawazpLFyYP
YMGBUn46O/Tw5MFV3erITD1ApyAhMI4N++CTG9eKUxyblKOngxNxrIIiI8tejA/D
88ETFaGr/T7RffH+VDeh7L8JQRs7ULP2c+R1PWcXZTg8v0N5wha78mED2xlrdOQP
VLidRvsyJFAau/Pvr5Unn3dj3XyrbnLb9gSCKjKN7Shv9n7OohP2Vjp/MHYG9NHH
XZYtBCCxoF1i89wzG0wtWpyTCSRjobZ/Bx3V7gGDLYIag7xjJzU56ouLSDQPsnEO
Y4EmZBY2veaJOsS2igwjYCEKkAcjYDuWZ5nmqV7Z9OIuS9Yb3jKZCdgoosI45IWv
wPNsiAhGgaUCbHZ6k0AaPkdFLMSox8WVg0OPsexFSECMrvTR1U3KUyle60Mtqhc3
NiEwlv9w80XjWcev498QC0/YUDnJUJJGRqjyl1BPJ/F9O4skv7RBXai+uBFeOiqi
G7ma4QsKBHai0U5qFv/nUWYDD7GjYruV9BazicA5xQ2+qv5I0cxgMTJw5DxwRVwm
yLsPiEOplngIWHPNmYe8eqWau6H27POQv/SX/IYntJMMiw1NmZJI6HnEClQwpuju
xMohnWn3vP5OVFZ2ojqi6lmGOhVT5iXTHaYZLDnLBm5DlkE60rp9IZZ+Qpgfmzo8
RZzFmqaepgNyuMafI0BXv9bNW2LachwLyfmPzkuwcb4gEUmHNCewccEHUf4KqueB
0Fi2QUidqPzWmmxlZgbNMA5EKToUeSV/T1/Wdyms3GPzpywFrkmdmH9G+zWF74Kq
7QBB8avme0cbJMB4/vWIOJW9l0B/vWfBEZg2mzATgN4MHEfACZ6WwGX+FWDo1qp7
LFWEjcuAdHmKPI3DbF2mH2zLVUZvKN6WDe8f9oZ8B46EctDAMjM4Qnj/p6E87RKv
VjVxGUcv4WrG8DOYdzEAu8SpgWSZG0ylS+oFZNW5fs32nlZObr6a/F4gnJmL0+wL
fBpUjAKUbwSFwwc6fbQuD8g5dbXkPrRf1v8wl/x4HExbMw+iKXgig00lDJdTCAGE
30G4Kqh5KqlrpWMljdvB0r+o2G0gFJE6M65TBzvcaGSWBcuzUqWz2zmBBdyc0qs6
23akZapgqQoprBoQI1KtukdiEzOtqnjawgDhhoGxtYW3BECw/BYSxFSg08gN3Wyp
MuXntwG7LfDKdhfqSfnUe1rHICS8npKV+HPfh/BoWMqkxyObq0l3rHBki07iuI9h
meXLeJHZbg3O2M2rn2AAfrpNPkOghajyqqLYdnXS+Dat6TNcz5WOEFH2h9+Pwmz/
8aqK2bMYZHq45THE2TdPw9EJSYxmauVWM+vIjX6GCZBmZVF3WF7/gFopZ6Le89i6
qW3e8mMcjmw9CGntG+3KbWQar5jbWZB01UhaoUelzPN5yodeJIcI18onMmbrsW8A
Can1D4IHXBYAEWJwzZykOAM9SV0mavvh37F34X84Oa+ZIOKvJns7BK6iaDt8Wdoj
VUNgbhCA2yDIY+dkZxOeulcr3dPvcRtt/c5inGfzgn5RIBZ7dZQApv+dtY68pSSt
shjWVDQD9cXgaD1baGZl9qwyMqqo20KQ/Sp08Unvu43U+Z/hSZGrG6ODs6Q9DzK1
E9faMc0ifoLyClU4MEQ5YcfoGYLR/CqerIKJEqbw7wtFOJtKl2hvSpPIw62GMDuh
08CTNd3I8e1C8Lrq6wgp8aKDlcvlYWVh5V7LCgepuOiVGVzBIq0nZj4H60Fq+ZO/
KNqXP4k1a8ZBqv+H0FqIgU5gDUaUyNgZ48MDlaM49sN2hvI+rnsQH+3TARAeKeM0
CnQz07x9FGcqInVfLssW27Tda1pn+i8HU3TrYfsRBVv7EiVs5bdwxyK6/yKvzzbf
MhLnzc3gSJ16AKGYFcwearo+eF6PLyU0Sl5+TT2Ap9gAk26Yey/Pec6tdymvZZxw
kmb0jJ/7cG7uxPD5nKNX7TyVv0l4lNpYNIyKeQIlyxHdkRyl5/vhWn4JQ+b7M41A
jajdaYKB5mcW1uBDE690OEslIPnIqvHOEv2PUbb95DGzV2z59APKIR+yUEalhNhF
zMPeINYxB+k/sH3Td1lur+s/YPoyjI3w1B8IIuiEHXhSG/7rrp6l1KEm/thmFSSF
viWZT21uJVxZnCti0pnMr7RK7PdmMe2TQQaRRXPmZDYTaRTCiFt7/JVhu5q+0g1h
Hi3ucrJzZjpQr723NMlTo311udqb6x3is43vPOjXXP6psZnsrXlyl1kq45nPTif4
BRUSJm/FlOInVBG26ENvFZ7zbxtFLFyMvZR6UgBHM62R0zLcdwvxzfBZv6D60imy
8uPjt9d8UoVdvi+Kmwq22ThpdChLE+U8patEr/+lwUNOKoxn/3AT8O6Wc9oxrt2L
B+E0DvgbF3mCTfswGCeqMQWexeORev7wBEaCE2ipcsvmaCIwFhANJdFwkSWWelyH
02s2GXZcgthUaghbCLttt7PPWlLeoGHAWR73nmvk/qvrUDk0syc2PuxTyIMx2wXo
GdSxA08fjHjIUm2jisk80Tw6/t6eYF67haGPXTqb4gW7vYj7IJQXSC2+0bNQCzKI
FJB/d1O3D6E/6UbI2XgyNS7P+cmKzxs0LipQYAvfMW9kEuli2HaV4SejI6qOXhW7
kU9FlJ415wJ1uxL94S7QLa29QBUv4jcIKBqp3rJZFePrfGAS07ARnIF0O7G1zVs1
EkLAcOaSeQVTMTRu0pHL7xbRPEXns4v6HB+jO7m80m8CImt4QOPHpgWQ/9w9GgVL
N44an+N/4/QaHBwEMp3M5rQbfWSjUakR8hA3tiUGmKU3Jxc3QrsOH2QF54p0WXL0
y0xEMYN7QpJ0aWmbzRIIcCvEGHtW3NLpebtH21uC4UGrVsLBECN2sWMB11wIpIjS
D4o7c9jonGTJKg+qFdz5YQ4JCZwaP/8i7JlSTYP5k9ac2X9ziLSkBvzX1oZ4xiou
A7I1gM+I1QTFa5OuiJ5CBljPRFNr7wj/FLLzjgZ2/+6ZXjwrh6ZQ1hm7QUNCCmEJ
m1e6H43XMQVASgo7pHT48Z/RUwmyh75u412hiX8zXMflrJduNfr7xS0ZeBO32mGm
WrvEg57xNdHGqIPDFhkOmlRQbNfchc5732vSQlo4HYRzJ37HsO2mzZpj4387KvLi
quMBfCwfCH6OtDDbX/Zkh4F+0KfRzaE+NR4Vi1bTOmo+9m6Dquih0SJi1VmPq42f
m2sqn0yNJuZn5bn/M6z4mZc8PMF66J28qruOlY+dsV47Cnmp80AhkItLSpJNJzYr
Axocujn+p3cw7OG3BC93OMRxYuWD+k53N/KPRpJupzgPyy5DFacggykESO5B/Jjh
7XbxaW4fU8J3NpJfdMqayfiLxATJmt1vTbLPPVxFJ8XnbaqU4r57XJKibcEsD9o+
yCyfatMj6a2Q9ICW5eMSn+WyhCONhvyuA1S6lpkOjHuOD7N6Pu3xlSbmx/0YBMUf
kVePfweWE0oUxSAq5WJ//CixANo1Hu1f8xBIFuAdc67E1BGhPp0iA4gza/5cSsbu
CbMy0yhw3gzcREcxUgJCXodws80FB63+21u2GBATaVrXCH840DLhw57K+t9ENlJp
ctPRgsiGqfyAhyFdJcnmj6ZHBgTN+tQrZx7nItob2MXJ8fLOHUBKC+sLYj7ThArO
iVdcQp0v90EDsxWiQPieULNu14Ut7+zIS+vGtYo/DmRDOgBvEy2oio7r0wXXQPjr
cjXh1KDLsPmbTAVhHeClS8QXNfjwHHkBPTB7zilYNho96G76bUJu1MUlNGNLB8pe
q5xBZHYgnkvCeWwCpE49wL0ApfYYQZVL7JaG3iExxox0PiFsCeJyGX5Ojb2cTkrL
uIrfAmcipBQ7koMC7CUxk58t4xbXlM1Gau2IikdNgJoFoSBQZKlHcWI6talixAUe
tjMxGmb1AaBW+Gk2kn5AIjgBoRz9x0jcDFfe/OjHHZ1IbvzJblpwXZbc75wjTnoZ
B4Ar4wzd8NpI4Y7FAjr7q6dNd010RSSZWuRdgs+6UYtgOj3Cq7xnPPba2B0nNrx1
9NUefu7benC13fNnefEbbxflqfk3hMOBzTvsaEzg9j9kooaS08nwqJo1p55ufb6+
YF5BTJldR4Daj04emBXE+sp9Bd6WWMNvVHOJLPe/CuarnzoDQSPYQVO6DeZ6TlxA
mWX1Go5sTotCC/eZAyR0F/MynnteKgL11Vj5nMqQDknMxmESSlqk18KEuhJMImQD
jWLmmb+j3u64F0tzf6WccU35uX+rUVhae6qUtZZuPdjcTcGMNj5ZwpF9UaOb+qij
iOCEG77rYJQ5D/zyR0eO+TXttxjFRKXmCxs4cxJ10F3bQs2XLjxq9whQ7gbYUV64
x4SSwhgZOBShnoG3vPxRqf6wRiig/dUupyL5YfqZ6PJ0yoHApWoO60IGtsFnXw+u
BZZ6B+IIYim3VR3H4tLIZI543sJiaroC/1arF1VgfMuLiw2ho48DSBeFcPfEIXez
TrWR15Z/nIClKYXqeO9kiJuDdddoM3TCkvFMBQnfIonZrnB590pHQJnXIHjQr7Ay
vw4G5JPWqm6oy1yAuOwtYvDGAxPSaXcwQNGKf2FTxT/9/68rwyVWy/UcO8k+1Pu+
SrjTJo9XGq2oxrJTR8hGEmxZ5eDBRtlE55TbJn6fqudBE6rsOiv26qvUclzPFqvD
ETEJAR1rKNq7ZWyJxqpbHl2uzbQHWUJqGCQuGSLNZj/jvCoOVWP1GQOOOVIwFy+i
SdZlc0+T9smQBvpQ0qTLS8Eqv/A3mbNGx65N3bpP3FPstaKggM4uLeDKuwMc9W4n
iU64c2DPhXmCIxM7Ca4vUEUPHqmL+e6lzmmhR8FnrTzQ/yabUUpjfvj4zZLoBj2q
8EA86fLWWPNdo1m1VZrAmfbYemjO9CQ192KTat2Xe2KG1lamqf38aHC3r5XH9y6T
qvmLJv1Ptfl+4lPsEQbzEDndxLhP9eLFDvlwdZRA4RuosxQTKp2qarejfv5kRR5O
ywrQWEA+FbFyYL1a6llDm8GV9vfndrUR/OO+ixyx7cVPPQ8/wNGjC3HMO/HCRNT+
eablh8YSreiWWumRVYliDh52BrB1LaqRO5DgJ8yfS6JbfcHqbuICQ9WQ9DstO2gH
XH6m342Br7eYd8Jl/cuHSDzA8ob/+R7EXW+i+bp/jcCS6NFZ2OYoQoEJ3DnvG6zy
LxyJcB6bkOFq0+kwRY/leoW2nVihPCUMixPSn+JOQAcZCTJCBGZg+GtUsHgUeXou
s1M76sjnx8Q/NAZVrxPcLnYKP4uuQwlT1AuUGZxg64UAzZr+LjT50fZdK/Qzw2pd
SDiv9a5LD/pspDbeDVb3jacgP5mWiliy0xgUyMQmlVsj9eoGYR5v6kuI/w0pw2ki
DAyUx4iN69OMxSHhSJos79ANqB1q0oCClZn420AiO+B7yRSQB/k2XDVRKzSTdC8I
FOXYULXx+FWZjs3WehvSECP/crW4MzzQ9nM7So/P50nTn5twJSkCKzJt4oHLCTJn
Q7enQuv3ScEKN5tcvhtBbLXyPLhks+r22Jwfgpos7Xru80OgtCuTbmdMaZMs4ndP
0W5YlPVvn9M5QJ8YI+LxsEuEn/0IHorqbACc9WSp55iHYjHW1HrEDFIICcyApyia
qBd0UVJLplorde5y7WOLUSaAOhxcMw3ShK2WtRqk+lerB14pYN5IhKP6k9xNAuHD
LHlOnuRQpUDOZ0tFJjuY23zs5SHJW1jFi1n8nmuyfOY2Hv9OvQJ4g09NQ8UMjJak
X+XAz1ly5IiWESMIO9PB2C3o4okXF1rLp4bkGuw7hyeg20ho9rDGOxt4a4W9X9pX
FZNi9nlgcsKj21G0x3qBz1sHggLVtn8UFceTSn/QUc4Li3TXzDsGmBvZHXahravz
X3cwP+l6iRZ8ASA2EvgxnQu/D2r2TjRDudRW+SYqv1w6NwjzGTpkXCvFRftx4sAZ
y4MPtXk7/JYJMsFTQsDPbyYbJL1KfZtE6MIPHGa9H3vIwwzplPyiVIP4MP7So04d
3F8luUhf5X7eI6EwZPZcxjfDbtL4Oaq77WgoVQgnffzK9pZG1tAdkFu13SRtPSv6
e6D8qDE9fPlEUXZkQIBAJdI5NKpy8DpAH9abEtGGKWfromfpbMiSOVFIdxg68sOx
tck/klYn0egBEhNlzRZCMKVvyZsSPRT2UFK55ZQJgRrmEnkXStcW9r4I208S1H/9
tMcvMUiyFErUk0OrjuWlXKZoDwju2Y+KECuDbwrAjCQZLc8pwAKM7wvOWmv8nuUJ
2Z2OQpHXTyUTjz8pUbHJsL3nxPYYlN3sQbQgHErEwI3Dy/WBn16sebuBWVUYV2Ca
ZBFgJtQM4z6ZMvI6519jfmx3myCcxYPXTZ1ovyeyw1e5enhUxIlqXAJ/HM7ptjvN
FhwIUnwKWELcxhxFYjADhWD2SM0SzMa31Fab1L6zxP9enDBbwxJ/sm8jfPb9OJhL
+hQrTR2umbc7GiLzwZCF//Ham/cQmfjT8/gTpc/18fQISakWPtuFPRTs7WTNCdYK
RIpzBIpFvVRgQWi6fHDtzHipqQqbgoJ5mbyRmOdLlAQLOeoymwtwlLk7SXh5YU/T
bYmyoeElxu+luJGMAUh4bvCVj+eKQpd4fn5P9e2bW3tO4xnTa43HInpMP2aTCBKE
cH97UdI1vE604zspw9coWIdZdugsIcPuT4/WfD2D+gyMNZ3ZQgoEnlyYnM4IQcSK
jAmk0Xt7TwW6IrNRVmgpGi66gsjnIUfxmXfY6RsWG03NIxz9rzcVF7+ycR3c4p6T
gxC5HHPqju2wvAGrg0KrOo6Vx8DngnF8yVR7n/WhRO987FzW9mtPYS4ekY7vCvu2
RCojZRdmaCuM8d1LylWR6TRRjtPphAEhE3hN+uO3tjewPhURJqrwYpvGdfEj19fv
DJ6BS5funs6ORNHMdrU20g4/gO/+HEVP7yFw68cpU3CzEX5I31LacHwryRaeO5qN
U/hVcRyndNOCMjtDxKI4ktdtyMv0uT+5y3+AAwjGq3a3H2C8dplFca5AnscZ3Mrr
TCGfMrZQiUU1akdLvdVPiR7jXMgRlKRnQgKNbNJg6xOP6yDHfVQbWDtIUBG5SqZU
yD6eZG9x1bLlphnUEZGc8p+0gMWmD+Pi0u4H/E0l2i6Qjnu2FKzHScmE05h0Cory
c14SAZvb9COBenxI4QZjlmqpxK8V+CKkhI7xmEnLGqf8tE8LZJeAzJsd5YQNhLfH
8Q7Em2532pu++ARR3QiekpJJYMFnbJw6Cv/oKlfMuoIE1212SWt7teeRUaE1Fmbn
Q5OFgZ3jrGRa0n1jFBG+r6bslAUcEemxLjJwj9aYPRCFrZU9zay0ev+CiiDIOinm
4s4XzYnLq55tviWChvRTARLpp9rxhb0evaB6EPq+MwxKfZCZmLAWV7VFTwRtv6Tq
Qw0oc54zjjyf+KT346/omVLZcLvRT/x3ZrKqoIbL8ICGnj6DMLjKWNGrpSquhsv0
jUKbMKykJ6JW3CYJUn0LSqWmz7JkUFtyOKPyKDzrWM2/J+iCNMPF+3rUDZxMSDEI
YnYsMXzcx5DK27cCpq50LtB5ykh07FnOD5q8WJlD/5UiXO2IT/Kpnkg/tYvs4vsX
jpNwTFGhWdukeJGMBAwYED0Glm9gPHx6t6xFG9I/Ok3T9sti7qc6HuglnbUeMMCI
ir1xmSLLmeJrkqhE7yU9QfBG3FdINyWIeADRnd02D7WC2Kvy2cfi4n/EZ3tN65D2
JJIaMqL6Qv+dCVCnAqyScQB+pXeipdEItxFl3pjyh2/RQ3L/n1BWFhi2xNm1BpRk
TpjoIMzRrzdBte8s51NuHoSscgSdxrvmNsy7v4vDaunrzI23Nkq3mqSzF/OW7Kfy
uMKKoInVZBKRuhNwiGhDCAR/ZEXr5mrR+L1R7NMPj8ru4Vr+yVGuJI30g/19tSWl
y2wuExx1lo5Vee0VBaL/6osp7tDvdPeeYwgYTdlR0vL6Hh9OqT6nx4yIByNnVIww
AeNgPRPyTc3Yv9OjPEmMhjzf6WNuUPZDFAnK7nMv4d7Dl+FcgJM0i1HBLN0kBgsM
rZ2qlHLLgumc29QD+PTZCxBu2ehpWY8tU93BWf2997PBIccjDWLpXIZiIVItCLHQ
kPXrg+KEnCYkWS+G1OwY/U+5Tzyv7e3fbZ54zL3Zxw0cPBaLAFw5J6uCJzT/RWvf
ogBSU5cOI1TAmV4VfeGriUCjSs6ITljfgVWLdzlzckYu5VQgc68WP38mx56lCGln
QGqyqxFVtMtAm7HQ3GUhhrY6bM9h5HOPQPXuJxCGjGF6SrCEx30dY6vfzzdy3EvH
C0amh7MKo9Z9KAjHHlNO9LvhZWtey5pxTnS43D6QHEPgTK/s/ukonLQGvbisR+SZ
skQmckB4xn0HRBw0MMHW4/h6uyzrs3NMhB+1iXBgh79WSJNKktxM9gEnRJ0jFvqH
UN0hiAfMg56IRnrpPeEKGqItksqrKorAlbTpWpQVetDaMWNBZJLNZ5WI55QlTlPy
3Rfv+cpoYlBww4+G0qBXSFbt5yVj9XH6Y9+okC/YXttd6iVM0XRObnb8qZ6v90v2
YfW+CeVY5BV6jmDIHHz/87zfbAO5I8CHWsghp5Kqr0TIshQ6clZvTdxqIpaYMGxg
sJFZ8LfNwTtiNcDako4TdYi7573h9fGAkmkVbJe1jM29xAu3qxNAnw6Z7/UaJnYg
aHIsX6nba4Ckgd7LSg1iXmtGUmGa5DGx6uYHCq+19A3aVyskc3N2RJYTIb7fGBk+
adIOKKDydN+KCWsfk8sxH68idvwuTEfWhZxu2ffnXv5HObqUtL97jbCAnqNbkLBi
LfYusPvBCt0D09+5lXNA13RCZC7lxU0hn789Cz1n54O3Udsiuodg0maDDlEwlv3r
7tO7mxv2pDSK/A6H4ET6lSOo+lfd7uPuRsU7d3twNC9CQLR92NG1aYIPTQONW5N9
904Qz37fHeqzDlV0YO+TsM7xg2yFavYAuCi+4dUvThwzGQf4oBiBwHCmt2++htDn
B0mRHUdzhzcO4HkUmt+0V7duCKusbPE325e9W3DJgqk0WhtP2RA7NL7IjPy5bMk1
DwrGbjAfGtoUNOWX+nSJF6o0Z9LrVeAL8KmQGjyH+tniKW+Eyd4ETVb11yJo9yZv
RVGZe3glHqtFnBzqioMvRZs1o8wqZi1WuW+xn0TF0wIM/0rQ0tVWV5lcZ0AkxL0n
rFd8M1jirZxu2fD5oVz80tNy4rHLerBMOFnNeGOSlDaQBrODhHfxSB262wCHyz2U
WFStVyS40blZ7McV5VWXPld7rv2uJq6PSgXzcrtfmOdvDIMEhtjxEy0Y0n5ce2Kb
Jewc5iY5OCVMA9iwSgaytojTix/kGPcHQuTTcKhH6b4MoQ8/C4woAzHtiwHkkan5
hW5KITqZwo2SVD6g7l8nghw4KFJW79BtlyHhQt7Uf9IFe3JUY0vVmvdPdVERiyhR
cGvBMR7S5+CmGg4SRQNRPfHopnBKNL53sR4VGE8ZswWThyB5dwXMVsGe+r81Rxec
J0Inxl8cFmD8/dQEOrSdzNWbxnoSNMVWGET+uJKi7RjWp/jvK+4GV8rPPcFZtnjk
F4eJ+NySqfUzb2l2MQLoPaTTQYBotCGPLIabQs0GLbLAgvGeW6Yn4euaAjkcfnQi
9ETqycxSgMn0ue/oRkCdsdPhahMUGKtasRbrLaiQ8r1NjstBhT/7rC+Yk0+u17zB
zu3BXUrizMLakKsqBvD0PSNdD4tNIMLEbPJHshT+4CTYLiQqvCu8/g4+dWPKBtmp
PzorN6BXQ97TyZdQb9gqqYCOmeU84ChZx4GYBzNaHV97w6QY+OkL6Corck93Nd3r
UGr9GRe/kG1YRg9Jng0P+siVsT4m/MW1ScSJv2L8yTAGTulW7SLWqTJmn5xc9MU7
dMfVnNmAp7+seDm0bjhRb54K60vYvNOjM/e5FTBVfXermqQwF6qwPOXL1HflDo7X
GVVu33/kNDtPvXNHAv1p6JitLy7ejv1PqweHV3W9yJF/ymQC8Mu4wTKqZapMpsRW
YanQ9gSvaNBoSNRfFip8joDvDXrsg8QqBmZC4d8XuonxkwQk/Wy2/HWsnCwOvCkf
NHiWkTrvEympWXBRcXErUtANStt6bcJfWNL2LQDsvqYlV1o9WjFIxVDSqvcXQgdM
29x58P3Eoid4Ekgq23jzPVO8uLNAPRgErtnH9Y2NCz4Vn5oyC1/ClbkcUfokRzlT
IY8KOPm2iDjYCGOjJBxoj+E860i/MT6ZSM+lFDBQxmMbnHlMrqqNxFIx81mBw6Qe
npo//IiyvkfitTb1c11MvZ1ukAnDdy/oFRKERbrv5sJeTt2uixnXdt7UMj4v7zRv
TDq88jpAhDrFYAfQY8lKAJ3HLcDzGnTBebRCGSzCqUvFCGUFUPQCPABijM2OIL2b
YhkgvNj80IcNyQIAmGMqB95fSJWlFZXz4GEZk4+H5o8jEDGEGZU0e6rf62prUs78
k5YZf9L8StPOyHu/mT2wwVXnDTGxzpfdOMlQeqWByeWbX4xkEK8WFnHzYu3xM6N8
IVinUQiw8SDKKqZSkOhL7lszfjbywVZQnaauQMQ9OG7iiBL8vn9dFPmVuO2qgEH4
acC1EU5V6ulnOt1kndN4YSNSuNAXRmvd20t1+vzuTwtSZoYcd8YLr6YpRyFy5uKt
OTGwLEjXvB0H1dbYAqRh8M0ZnZEOMIf27pkZYE/WHFO1YWM2IRMWRH09IeMUAOo3
T5/kVTiejjvextF9fm/7xM9LehXL7d55mkXLU67dV6XipQMuQXH2fV9JEBX76wMv
0GN0zWuuDQd+fXkw7cCWcDfe2NHrvoPBX1QRdTR2uOgORsbEgcDd0mcpEuvNeydP
dicgH+rnFWYjYeXSxgIerGHLgR0fZUO1lH1bBw7bhW6q39ItUL28x6/oZVq5lzZ6
HfVyXj7C1oWCKg5xtCB5x+g2MCS/wox8b99SmPT9k+la4B4KeWKVlP53MkZ/ZAVh
vWYEeJgaRveZvb71+dQLpRNo1tj0pmU+Gdr7RWL0Lnt/H44vYdCxlZ1EuVA4MjMy
eOJlAhRAsKXbhB+sCVcMsmMeVh0PW7FqXAxaSVRbtC9Acqau+0WSrzE4+td36beZ
VsPieP7J3AvGCaRfeHjH3BGQZ5iPwQMgkOuM82h55zAv0rJ/dXA+8twqSK3h6LkZ
I7r+IPCFS3CiaHezDji8OSzoURBB84FEQMzq09J3FWzpNnbA3Aii0ESE932Y4xij
XLWbw/OtG134Y3wwtWaIo/THm/fua/4iqrxTXqcSrHrMidPblw4tSndQWULyChEw
Tpb/K8qdB1EbRfpNAPvBlR88uy8Kxn3kEaWyb2Bip9D4Fl6pxfqSCK6knMPlz8zq
69z4z1pHwtK17dmh3TIYnYYS2J63XgTXcIpd/O9wVtWo1y6N4OAeulB+ehm8WzM1
N1OtcbwNXvUBSo53NvtHNL1RoByNLJscky4hLfQ+3kQ8rbgVwp/JqpRD9ovI7Sk/
iUd5JEjXCkNiQUi+G+3hMbxyZkj6BIEdsltDoGUIZCXtjzeRXpAUBFg6b6/LPoQ2
8eL4meXEUnmzMwYZQ8X18qe/tLyXCL1p9qfgHw7C/mKrxdvzeJLwGIwZrNdrjMqP
d3myZI8smYzpxlYXtVCt48a51EmjTE3odcapDQA04nvef23DSO1OzpC5NzJfIoaP
y0d9m76CVn8oTz7AJgTssKsb2uqSF1YPjtx6Grvk/xaIevf3tL7vYg9zbLvCPIL/
EKd6N8iVAH/AFHF1wWtmyapuChyaPWjsOCK1yyyPWjKg8KLHgHuhjjdAq+oFQd5v
qFo1T+yaWNIwKWvugy5OXxLiIxC4jj9Q2VInAYrEix3P3nJW8h8iezeccRUq5K5o
CrVMhy6F11KQpxBxU+/4psoVmPBUpwtrhRRN7j37saRYmHuN3zcFUXc9dI2yGfDM
4gbTVt70fniRErb7xVv9KXUSqjW4IaecAkvyvauK4NQ821ty/ZdR1IHnqqJOluQr
y2V2k0+OubSEk28DLlIVvKRUG5d5+tLZdNx6QWphFEWjK495cqaRDMbOihCLOye0
6MTbgSDXlEsRRfR9BcxaUu4gqDTXCvs2fRYQTPkWgd5DxkmWqQ4dPDxUuF6BGC3P
S6GDqPc+DPasYtgchac4XPnaLZ3sppvEZZWHCrxgJF4a0KUneQXB/EGPE/AiQeta
DzyCqlUdSbzvdqQRsvP6qkknLNJLjXgnZmILguYmN6QI8PsD+DJLPNZb81Zzc8C/
1/f6aC/K9sNCYPdN/fTEa5hkToBYJZ2QiY3/mxCy1R8A3KCB7m27Pjo/tWdZDOGc
dJ6Jggbaz5mE+TH+NzW2cG8YZASBhVUuw7XmaER1rUuu59EHsN17iFWTIcyTbX4W
HbFxBihFyWL4n5xNOvzO5crd0gzF7fcukVy2Xne94uugdmq1ayon86XQCLMK5LI6
vIaR6p1MpGw3mcrOrML/H/08bZRgJs0Zc64j1jZ8PVrD223f+p+4B+7zBKwo6uUV
DH39dBiTXh/Quw4jeK5rCbIKHp3AdglGhjJepygY3GKMwiDjfaeFF0Tun9EHTFK6
pw4JFJvgMWzlhi8o8YoWOBzyEqjqu6J3ELPR/6rJPISJunxpP1966RJh6Duc3Ae3
2bjiar6B+Xq50aS5WyvqElqesGSn5N66GPZW6kVzizwK+P8dzeAWmoVatO1/pC8B
3uniGEVTR8Rbydln3iwLH9jcBxhxLaDi0cdcIDSVLmsaqhS8dY4/hgFs1nQWnVn8
W6xeYi5gPQD6/K5E/rPWRGEsFuC8PEB4pIWRtPrXdj130c1BC8VQmNu5GA6yulOd
clWgPoYEpmVC+crj/0AyYa6fNxNkfBV5XKS5oMPpHel796BPoe3KsyqTWeOXif8X
pLNpi6V6tau/mOCBgjObToqaYJSV+Ym+Wlx2n4JezvRD/1fLzapit7Uo4aS/qalS
jWhoEV5hQ/vXcmNyx6yYBdl4Nr4ZtvGeQ8n86vREznE7DVsABv1Dy4rfz9qjgdjV
carryadrX3MzdAL/zdfsSfvnY11iomLNY/joxX9ftWpj5L5Z140iFPGJZTp/rbgB
E8CgJUOIvdXhesZxkfQ5npr4ClsJSc9PW7JGvQqy5Xwj4cTnS964EnjgX5U3CzGZ
aBzmDpa/SXS4Qn6ekkHDx4MG+MeEbmoyGBPTaHnKuaRcLZdnH2HbB9+awPTXne3P
yBCOB/1YgdOXCzDnBNTuVLmNHHIyp4cex0RD0B757xST2qZj9to5ofpXFDtz6xpy
4Bbw3bpqvIkGfuu2bpq2xiS9lvxXYzSXWKY6k1K/qgLpP1VtSHnAw3ywdjiv+GKV
pbkHzsGsUz5+/wbPc/kKTXMc3Q+eChpYw6pj6SjX+//7/s5h4gbJA2W1GzlYe3/d
7vGP8kfTLPzvlBQcKzosF432/CrX8WOPQoQiqVbJSVy1tT7syujbX+AzV0jxpzZ7
gRGKLAki60InSzy3rb+4723vfAW/gAlBDozN4ehV5uOJAWJrKAV9wxzXm3p3J2pP
81r+dDqbpnX68wGJFL6oDrE3kxNuJVyqmjCOtuzDEwVN5nJTzHOSbgFjzAKTqGL6
BSQg8E0/f0KBEDJN7tf548H7hu36KkaXImY9p8Y0Yl5EoaZ9Lg+lDxwLP10Efz/x
4+YstiTLmVVU7IEv8HqL/V6n1t3gLagHidQGMl+1in2q1ne2jo46sDJ7osWF0TQR
nn8ndMyz9C5tnFPIgB+tmhMdgSlVv97yKJXhVlHBcl7nXorhMM46bIPL3JTKGt4U
tp8Pb9a4XowmpBjuUfT6arivWyBEo0nRgVCOF0btjJyxONMxZz90P+DI8RaOT6GX
+OISojtmxuZcXK8r++qo1F/pOdEsd6B/fPGbkUAt7K9uHWv2pX2YOxj/OwFbIrYq
YJMNhdWWqdzuW0TrSlCTAWKtHXoxNTCje4Qup0zw0KxPqEIlMplWV8rVSIUg1DMd
lwL96tiKwwRXxRF5AHSQTLtDd6HMxfjSmNA2MT1nh9cJQfjCDwXDz467jeqtk/xC
0+c231XDcdcRJrBNsj4pGrQOeDvCypXki2qGP/prsbC92H+SV9dcglwSo1bl5Tgu
s9JjxEtnAj4HAowww9bK6+ecnfu8rA/5h/SSBJmymfQxxG8beAtfTFjwYacA8x2z
FBZYfd3QKMMd4m2CYygE8krybS3euvCa+nDvFUh8IYb5GIoKRzbzPMpEojsud1wW
fv8+CG9avT5/xNQZSaOsC/8fiwp6cxRrjFLcsVeymKrgIkj7i60D1uOJ4AV0Nr/y
n42km6atZ8NEg8CFDGa8y/QL2KjK8Ut8IF5J8XYClYlD4CvXJn1YRmNIluoq6QNf
1Ys/Z9BdzDTHECjELfGmhzGL1HfqnSzQ8ro+OqwGSxxDWmaSPIYnIdPcvXHk4egH
TuD+yQtg+mFjGnNBA1z6SVFaAZQnmUJi+Nmx+Beu6ygA3KbupXm2BtsP0etjEkyF
g2KSxt8PCck06F/TWsaEdzxALa9dog16b7q+OcZJ2BWZWF6LM43ckqMNwyWRf+Bz
nVIZ/VJwtA7dmJuZigkn3KRiQPFTfcQRF1k9IF0QKOPQohT6WOtDWpHppopgQRYw
RleC2ju9DbyP7eLReeGh3PONYR7Lr7tivGaLnc0P/bK3fR1GNJLlgeOqVmVHnHaq
tPZClmGCBmlTMEPUOyfd2bfgHqa8CHLRMqlcG2mH4TB/KeMAzyD+vsQJYH5i7o5X
FXmYsbigMKP0HTsk4mbxd+KTLFpAF8Xhs5dS/dml83idspguoXxatQkEb7favCNg
z5d67OQ6Cjfs0DJ4Okj7PHz+OKiRBX6kflFeJIMTFjo+uFxmlcy1j/z6ClPtnacN
q01kCC8SkA6QFpJ5z8p5ejxstvSqxP32BGdTQO11gpCovKsO8MAzd1N+Jc0gV14z
En7o52PcIVkvsndQWacPoMDLbHaGRT4+Bcrpv2PnyTIixeM1RRhOw54Xqc9SfDbS
oiFyC8qN/2Y/XneGW9fJ41GYQWr4M1yjrgt97M2ik5oah2/JKMOO5aDROtEFYVcM
LYnJtvlJPE/ScWL8znoBVcFwmo7c2QYy/T8VDS2jGrixpgqktoJBu+U/ePsJjJHq
nGHyPQP2yAKnBJPVmngJPkkVAh8zGb0H8axB74iZhfwTCyEHuucHeG8mlfMNkWRG
cjGhz+XC/k5QH+hnrf4j9S8OZ2q0mqv5NOLOdY1LmsM15Vx8xVh2hpDL4rIxuItk
hkQlsIFw4yyudTx12XDvmCO1MxG1PuDP3PFBUp9JOFv/LHmbvDaKLXb21UYg/uDU
MhOkqhY3fxRKRJ6D+Vv3oUVCVfPJMiC1857NIGnIvAv55bqBKZCGA0UFubb2pMJ9
Coa5lf+NyB+MjY2Z7cI0LxVZ0sMocdbBQRwtMF4stBEF8DuSQ8Me6Ck9nw1IzrsA
XWL1p/qCtYGDuaFn1cj5eLl2KcPVDvtiqLmRnikXu5ZXwNszqnWZRnNkry87mwD7
pDdWBeZJrZS7mkSaxy1ZUm9Y7YxommtT85G43bMlY9WiaM1XGZiE7WcG1vh0azBV
1Au9rRtWQoqQJ5xWD8CDU2zmz13pIuvr7Z/B46zgsPJRzLkGCk7td5luOAqPGfWt
j8W7KcfOGrzOvr83ZidCE7flw8hSzoEtwq2cJpb32kZm/Ml5x1vXbPyt1qjJjvt3
fP45gV/qNuDMMSI4xciREEuGeG/hvcgDzEivuofEsHnU01Yvi76zbD/BhksGTSoV
18WhYA4BSSIgKdIcE3pU5xIolEVytnh0dkufKBQKnsuPYl7cvasS9uzDnuGqtlb6
IdBIW05ytdJbfCDYOAapJ/YadnS/mzH0hZVy1FW7Xc+XRHAm0uImaslOi48wTSsJ
n6t3pyhRIxcX79G9Rx41rlJkuliOv1Eq+Rwy78GtyXIM8xK9hVsUFLb1ZOkqNdMo
g30Uh8/HgR07bm2znG3JnpDbnsikYf/qCA4WmV2NAMhMtcwLhtBgWZ/P4Z+WLDuy
Y8qktg8b3wU2jpfRdtMdqzM/ryq8y0zzcs+SEah5I33uXpQbL1nj6x/p03LOYNSr
v5OuWBTuQUPwH1NkkKHt1Eg3h2bRHMKRRxGP96Rh0HprlG31/NS19YHqrY3R2rCt
nUh9kg2W82ge1D7nPJcbEmPyvq4p1sWYUR6DUxugQmOPy3T4GK6GPfBH5edUcASK
uIupu2jiySe5yF8rAzrwShVmZrTvlNr5+ffDK5GGEI0PRp9dAFIm9ZgkWV+rw265
lq60zInSOt9lzSYsCVMGFdsz5HMU4NBFKS9vFqnAxWYePhiSP5aqDRnn82Cize4p
N3DbYE1l/5drW6EwnDxYMgFQGoVWZrkRF7HpJMaKJh62bKRM7JTnySbKznVU0HFt
AHjh/GEPUU64wR0B/9ydl5HHv13Cga4zHaxmWJy5afSXV9pFm92QyjYUuduxizEZ
ict7HjYDp2dtswpci1ud3Wu312EA7Kqb9pPNYqKupZKFMAmpv9EKuXeO5agoJgxH
wuvmqNIj6QOyqyTLidguSNDbyazxpH+CgLEDlOE3dkWkOKKwTbDHh8nfFmPR+UTt
GRKiOna/9W6Aod4qKjhmbUc3/ZTaG62lznHwocnhd/v0GLb4Jkyx96Qm5+Re7a6D
SizL/VSl3GGQ+dOavzjuEuNXfZiW30UhQ8FVTRIeu6l4BLNDkUTrKo2ZxEzO6/a2
5JxZSNnlKcIj2Tc4/ydszLoj5TFNKFL7nvYFCZoDlwsHEkoDmAlH+yfYPVE05sxj
KWk4SD2v8AnuA2q5uG6yut6fcEP4djOzbK3KAGQrUa4SkQtV3vCcqGTNDb+ribpO
KZ1dQDzTXtkT3DoAPyBHjx1fKftHNNv6MxSF3jcYOUmbJyPWvLJ/VLVrtL/8kguy
8fmqwyemLk9M4qfH16ulZ5M+rIm0VSQ0zoBltnKX6C6PdkLKT01CSoCru5SHrAmy
d5+UOpDDiabul7JAx9/c0KvOv0xGll5rMi6B3NYeO3h8B0Frx/iYnMCw/xg9mFVg
JfAPuMUFuz4YUGT6sGgp+ZvCgAYsARDfxFG4vOWw2Wpfx6feYltiDBnpsYwDNb+5
+Ci3WDGSnezkdhO88F/JidEhR+ej+3FaH/YD7hHp1WnbH0sZwKUwdh7c+49tfIER
wXnjcg2aaPqaDDDCHMTOH0QPe+csXSr9AAWNm4sCfuCV6aoqIoZSs3bdd+WgQk6C
JnFzJu9OqHn7Nxgydd3ES67KfELlwP1r2btKU58MSX1TEmtrCoQTd37SBMSx2eXf
n9CuUQRZotrj9PC+2pkLgxhClwx39/l7PxoQYUoXh7KgGDfjvFVvS7AlGAv6APvt
VOV+qFTbYdavSULpthWJls7z09rp8MwE7yQVlBlPkPov00SvDzmXaDbVD8iim0xV
ecBg2DKVFjoHrEpLAp9EpNf/GS1TjO1ojhch0XVj+QwlevBZ3cBDKOKb5/0fpzrW
ICFv8Rdo9XZIjsp1xKlTe1AwPx/fheV81bJScMvPmwKfMOFlLoTkXT3/Vm8I1YwI
rphWEF8uAPrGqWLpcJOvxv1bHtILmA9qt4XbHPBxkkYaMx4QAWSV3NMvRlJF53q/
urdFLgpDipMKlMxTYaxLYyJ8Gr3FdNG4LJUQ3P7YraBpqOAUhDT9aQjEycQfCFP2
nRCt7LyQ6Yhhyrn8S2Onvw0nvxklMqAkgZncaX/9k+f9XqBitHI6tBdD7x2Ln6PE
9ntSTq6XhuYkAY81D2iNeTryEPelkoeuYvOj73bUOUdG34ddEEBRWWz0Cml08i3n
7EA8vREwLxDW6Ne+1OsnVcMtSI8Xz3sJNNCbvTA6IO8HgJFLyPrlKQt8rZmvWY2a
b4JD3xajuyM9Z0Rzz8lPuIq919hznccE5bCL9id8bQOeuLqWzqisEe4pQs1T6L6H
Jlky66VzlzI4aq3o+d2m3wevetPdVhXMqp4JPayS1dx6uijzeGqw0I0mHWW3Qm3p
3ZMm2md8ORomF0RRWfPQS5MJRkaieln01uCzo0DCsAeAuPmNJShYK/D9SSvF3E5x
1honxRwiHMiTD5h3xCZ0S9xHdHAvRSst9N9X8HXD9ZgFreyASNgPKppSSRfwBD2A
bDpDL6Jz/9CmuOzBcRl2GbaAjdQTF/+NN3mfX3tnRo5e3br5TsTM5BFmEAfOEmFX
sDY1BGsnhBcU2o67V4vU5ppQLBrK3Wlw+0YOjyvi1M17BYjHEdQgi3lq7yZMl5dH
dhmoxlwjxIKMSZ1m7px7iXjviOHDr2vyJOGJAJ6pOTlf8i9Ydn3+1DNwQtheinfo
Xeo/8T7W+IU8o2RlJZuKJqlv4un65T097YpgZxomZTfwqsk/icbHzqfYes4FfPp3
s68SDW4OPe/F4wpeizCiuYt1ijWd76PAepMk4G7At2X/hVQqDGsAd+6ufcKv1biR
fdVxM7V1GihkxqYNhwCEyBZxilBOarbcG2WYJZhVYZlar2OPx6iOPPahKMO6L8R6
cg08M214w/SCVwh2OgGaUz5937QYnv6LbshM/0cwsTLm1rYyZaLMkTCHuSQSFFc2
FEu1OFw5sDH19e9uCN6FRWAPAMI9CkqeWgqqRHfAoB0HTUffnM6iTEkOoLUZ9iOf
oWS39GN86fZeU3HJM/QPu2kF9Swiq4ZMZ0w5iZskCvOqIkueMaw8yIOQwbyiBjSu
xiVyulo1cjc0fz+IEI/oXcfY9Uo3fy/z8xprUltIVf3KEbdAUZvdUFUR/IWRdh5z
SgUFcG28L/T0alRVdNKLEg04DpAVFkNE6go9yuIWvboOC946OrCfgGO8bKUmcBXS
uwQB4nEYGEeRuHWdNXVUFcEkj6po46YURAhKTugfaqWCG731wUxoVS2gKDFI8u+g
dhEeaWg1DZQJD3CXagv0wfo932XubF10tCAXiJK3uT2SJ47kqUHOM3fx2vryyc+w
2JfYqB6+bpNEMkOJ/CyMghTioLnCRj4sKYyAkbl70uZ8HXFQtsDe0pTy7/SOO0KU
Rmt23G1Hjtwh2/hNFesnkHYqPVTdRbBDsUgXFH4w85ejfftqzmnu2xrLIlrWFmB/
KlH8XlUcgrs3UU7DqlgjgOF6aEIyfKZKC7TRhONLj/9na78R0mB9fM1+O6RvfxfB
uHP7c7sIPyjejrKhxchIpQahpgMdaRNebDDXabO8Id87uo+1aeUPfiiYdWx2wINd
ka+CtXoTOZpC/yGAfdFds022GmpvItl3hVpGtZwUIq/CkQC+SLGfitrcI1tfmI2s
p+vCJlnzL4dbSvMh+KScxowi4hrzKJdYnQBXbEFCc7CH5fLFudEaVGyaqz9lF573
+3rfs1G1bc+9QFKF5ZAeY4ylDoIJ2JVUCyL9zFJnGwg+fvWK1OgL5LlZejloMsla
wK7kmUjHVzrQ0mtTNanfgWF3rbWFoVufJXKPsIw7HsUAGZAOF/dfmsQn3BGyE53t
YsxCaCF8UZHQPdtBeGP7ZO7lxWoU+cQyZAK+JGKcsmDDAVhH8k/BSz7vezh3yhgV
mfayqOWewH6S1M/0Q9eiTijGQtiIo0wd11kziXQPqgcYINUHqEGdvWBloVFKzN1K
2vneLOK8NPC7csZxl10TUuh5z7MGCt/5M0CL6DDwwyOE35TQlU7pLscRC9WrudRr
n8ruMKV9qCob5lO7uvp/YN7dAdcPxmn/f5nyaKE820ucWlNvYdOB+pRzO/2CY6mQ
pq1EiUIdqtHTzUKiwxS7LNaWL/Ma+sAk4qvedDrY7tITh5PWA3kDArUXneHZxGsy
ZLs3prmBYXLt3yhSXJo6tWpgU862zyoiwsvDIHGis9SBq9Szz3S4/ccvmMzrVQGv
HR8gOUKvIfkHS4ReGexJ9NCPGOD8crADsSqBw8O+PpyhiMH0plRTAXZkytP6NVTM
3KRgccd/ioPbO+yCtkuCFuzDO9Xe1LNLfd1Jo+vXciLTWyWik9X8UJ2Xv19JFZ3H
UUU9kStwLj+1NztGTKYs+yuDnkiA9ALzKt+4FX1ILmLqaydD9PSA+o+SS5IXGVy1
2k1RiW0K8vdZUKfN+keTHqfGcHQ7EHCzSyfZZgy48cyt3w2W3HIknA85NQPJp7x1
WZtgD+JFDf7Pf5eMKlICNnuXi7vxtwBc92HTNpGGXuf9QaLfsXa8MipAMUC6qkLW
Ncei64Q9UPAqbE2ZIGX1KHXHE7Y3iuYf6w6pcec2F4aOYOt1+rPx95CepnQlD3x+
CpRZ+Ui1JpIiC379WwWZq4+aXzgJas/kveMBX6atv3nEusUQ4Yn23O2OH/3icx/w
BN81c33+H/wAVl+ZwgSKzUcFSHOiNWS6/S5PjVxa3P1y6Jer+IZ6XOqXPhpRjXYa
nVE/wDorxQ+/HLnoLz/OV/H/+4Ja8ZSXNLTE3vNNASfLvDNNIe/vo1r4Qn7YV/7k
oM+rfeX1dTKinFyvJL6/LFheb2RBc1cUkzctyHHfqHJmxMkNim5zXzBYv7OP7eor
jcxmwpl8hEStMYMs5NfKuQJCfuWenHlA4odj5Wu238/+Mi5ocCjEVlQyc+w63u8C
TPofaeFBVE9yfV+s19c1Lp57GGIvZs19iZDywra2YCopqISHgS+E62gWnV2mIAkZ
1TAGnI/ykVm6ZlbZaYgAVwcCZwpBjXEPeqU4YebakYdCLp2tbFbTR88Cff93H3q3
FWPU3bn658K8fKaOozlpyzoRCgwE593b8GV4BE4t+Q9TcMwSE4Kk0cqoMOiuXrYC
zEX90VyAqUiCnH8eR83lsOJRmrHA49aqhCy0/QyqFqx/wRooXVVHpIT9wjYqLPZN
SzWSaDXSEpZkvemQAkL0ANgsQXFQ1/+qsGmdCa/gp4yypNRMxihOoub2EUiwoTmt
Qgt29fkG/xGHRX0UJe6JlAILAdbET1H9C99Af47zTeWbrbFEpT5cHF363lcn+fQa
rlepN0xO1XEO85nJTYx55GCImw+D6XYWTy/iGYIKFyMcgfZrS6M6VMgc+27PMFeb
zw/YsO2K85CL5DLGNQMJj4wVfCHlvJIUZUGEQWRwrAUp0jps8lpxKnmvVVNH1kK3
86J6JAYPGUezAmLL9ghv7ALDXSkfQi5KP841dEQwI2r+RQaEAIuIjoy0s9qQlr8k
daXYQXequoT1jwdKPodUhVbO1hTaUU/YrCjm3HM7ETHPvrKuBAhx6h0wGsudX9SZ
tRNiNVOO0txRBPqVMMY+2S033GeW5vtPsCCuC0ARqztKKPTJCmiH0Q474F11yQcs
AGNe1MSCiorjluyGtxF2Pey62f70xOhhkjA4YLUH/tYbJ9ewDuRiAh0lVb8I7Lfj
F82No1jwZFZo29FYZyaFDGB1E4UuwY9iLF2txrAaAMwMubUGwaW60hzD4Q3S+7SS
mp8UORIFwfMwm+F6RSidXFIb4mmOAYGQZkoSssQ0G57/NSaPTTTQb0IRMRwnzZ5z
zAKzB690RWzQjRAQOsGTFU3jcXrFofjA6OZwHM2jtkm6b/VRwHUbwUur21igVaOd
7l6KPkvkZ/MLwoNDmX3hLuQ31dYHFpCDpm2XXcjCO/pZYd1I4rZCU+GYqHrfQM0m
YlbVAt9mPwhVKMcP0WMZZ9eVUCoVLL/pyhygcBiPIRHIgG6ECMWblQp6C8gzgVpV
+C9Cnb5Kb3PAU6mk3v+WONilXu8A8rR+tVwSefex1o//UXUqzcRksuebauRV686S
TICmaxAlH1YyQnD+nyhABz2zwXKkQ+qcPyjB1Fkr8L6U4kXAdSjj4AuztW9/Tetu
um2PF77f7i3WQQtScTfe9hx6mYvIJWA1Kx7FFW+OvlCd+KQ/jgyZZPFlLi0TfjIg
A6GtsCbOKWgW3gQ0ny47Ee8QDYoGTKzIzSt9gPUlImIssFs6lJJjS9HK8Q9guSsM
d0J8qBPxtKVIyjbFWpdhmV0LsVh2WrrFSpflfX+OHIsX7J52il+B+bs6csHc8r30
7sAr72eChNotnJXKaTKcCWdxzixop4XqeJS5+ocYYLaEkL+ZIon+ZbkRHyt+PVnD
/w8gZz33l2PGuMAeom+Hx5cOzOWBE+0oqOqgyPcPBPP3ClAI4wq2puDu9Kw/Mief
mvolr5mlXfTOS9A62N0DQoiuhCccBWI33CRo27TRbZD5KqJ/BID5Umrb0zK//pDD
tzY4M/N8EzAb0iwOWDN+euafChR+scZMByYGJeujVLZqfB2yHmM45f5RiFtkRuz6
AQ7XOGw6U3LP69RC5lw0VbIhlUkioNopWXCSuNSAqXCYyQvowqTz9uzNDLVeGSec
QD7QXIrx0Zg9OYDri0VnXKwJw0RFSaVLed3iswm8Bv9MobDizhMzVO+ICW+YIOZv
Y7f9jIXU0HltWoEArgVGs+5csgM3UAjSuJKn2yPCAN25nKcs/USGr03YhUu4Ly4a
XpvFw3v4sm6D2pDDDGXHbBLBMCzIK02vtlRRnMakKN65o/dpTmhfxuQ2cHZK9eHZ
84DaMpXy8+cwpYYssFaIK3XeQrPHI7wxuJM4r0/FUtAoYLb41LkvwKaFM5kBHJeo
Vqp316YvDxr4dINunmzSTpqmeHGtB6RKFR+3Kev4TorLFJ9ffM/cNkhnyzdOUwV6
lQyKePQ1CaI1+bEX3tjkMM+jnREYtCbxlPv9yDH74WENDH6nrN91QkKVScQKVgfu
JgBxHrhXDXROlYOqzn1HxMDBcVZ0OWrfVFi6JfZFoF/YTG8evPOI4FmE/xWJEwOe
gM1G4H5hpDo6cuDPYh6kYsxdvtxon6Ndd0fzp3DKrpwmepogGDtFzELcRRaych7N
YQICM85i9OufV94+yc7U8QDtAf5QP17yD4XaKGJxHY6rGB0WSgR49Ec1GPGCoWtQ
zBTH5k+oMCWq82nWHiraWKT77EUp8/bXbTpKZQKfKG8i76r/ki/JC8QxDj7YCvek
2D8eCZdRKonGrqYLxsl6vHw6VxPOprNvYjKk5YLZp5rLqEzwNHCHK73YaGYQ8Hby
PEgjVw0ENfRuXPHEMbkx/Vqw8+BXSTtBMvpOhqCZwsTGc0dC0ZcLmxV+08e933qT
yeQsUWpCRyYyOlefEEwLwhCoHTBocpWTFwkrVLe1IupP8ayJjYHTcesWcxHTEADq
5o2K8CcKH+NFnKIWC4iPEATLtyp3ksvGo+gfQjgZaKlzufjMyFcBWNVgOWWYL5vZ
YqGHZ9dwLkveJXmc/16K2gTT89BKR6rGHD3gK3BLXIi7/iCVANAmYLKkxCqJUQWF
UPuXWPjuPZVkkT4lW956DM5AABxaYG/tZKlGAEHnDgnpdCdfJUSXf9pC2/OfEgzo
D3Sv5xeiIIMs9gWJ7m3OagKqAup/deG3z+Wyyz9aBuLeWXUIPV8B4mEOMbZd25QL
31ABrB0EJ9N2qHmBl1YRBifok9Kcgdl4lzBobR7NabTLTa5Myz451fgYz81kgupt
m70ksk5N6i94YgyejNF+ujWkQ8ANSWmltW/4HMB5a2tdeGwVu5oOQPBxczlVl4OR
e4dvzy2qMmByic16VqiiBQGhe7WcQkjssH4gM+p9oKAdSpr6Z/WcawA0Y3WYO6Q8
85EOIUFwSgWxaS2CMWmjucl5O6vSc4MIL6LBL01/8CLAkZ2ceNW2UpT0TCxESI0u
NQrDLtBORrRjEAHqNS2Lw8O2f06Sl5r53K4jbhHDIpB5dbxtg7dsDAoiuNYa1BUn
LAVRsSpMFMLfYZk6mTjHFB5aZ+fe35vpE3+Wfpxe0t8sR90vw/kJzutMCPXN1AUL
zusvY0FU9Q3J3o9/i2t2jXzxRLjsgopGfi9IHW/T17LGG41SpL7oxf2WnVmjFFS1
C2Snlw0HdXrryTxGXS8HbGtBcEFQruwK+eA6PyPevN7W5jmVMqvmkMEANr5Q99aN
s0MfbBxxDWQ4Q0Mkg7IEFfy0YQtY+o9AqgKcDDp31F3yWoPwKWj6ZLAP10Vk/WqT
XmUQDZ5vHhJRnJCZRKIG6GArbuO3ZF7UFn/W2bOYMcjA0bymBT80UQp1Rqjn6TKd
NENnC4vu45iVN3xXFZa3rkvsznxx+Wxn53LJr9HQ9sJvdnltraa85FfPo45UEWXD
w5/EBhYt0OhGa0jahC/oPbWpNQq1RnP4PhF62lNdD/kuIYpMCTdkCUGBtYKewlK4
A/yeEVUDkNbU0HRn4dBM8uxddSjfg15qkb5EO5YT8lBniPCR4PojTIrxQDwtuRLc
/HiKXJn18WKcM5dplaOj0tHkezAydxF8z5ZueNwIAH3KvnyCPFRU+/cxqRTghCjR
vOKD3LC7VzeKO7qLHaUFP+SRjp6WIEAxWbFI0gtNr1fuVIv+zzR2A34YF5U+Y9ww
xhwl64XvJzF9FFqlYKdPjGsjHjiGmaNRu04KEx2n5SpUcmmuidAeZbX/un8tc10y
JFTJr/Mgm9iFDJUjc6aP3HgvXraHzIrILGU6yK8d3A+mo7/i0OV78X1XXI8x29vk
3B5LdlJeXFpWxsAPscP5GS3RF3q28BUcz0hejuXN2qXuRkIEm6ehQgI1ezxeWhJW
p4bUwpsUNiXUpKXu4L8EPHrZtqYeoCniKk5cHzA77oGLeNf+rCQNFeGPSaXbIoaY
wCWKsnWTDTCW4ObFeKTVpzkkAjTOFIjoxXGF4w/1o1CoJIb2oI8gwVMXYMVsHXXp
/a3kQ1mC+8oGhQsssvOHWvqMHwBkD4oStmoIGc7LWPmoXcD2vvVmyRdTIA1Q2/1o
d86nG5By9CqYCQkTDlWEyk+u0PAWH+zA8u51ds1/aubTgx3LFXxsGC5Xd0CyuKsn
mhwZWmy6zVJKHfKcy8PiwJo5vBGT1GxeA6D0c/I2Tkp1mMXTkY6kIF2HZMgMwmVj
MEuWiL64C19Zsxh+PK8BD0Y0hqJ8xvHlOwOWKzVXFTFf76e0//dZ2WaRx6b7xJSB
p7l3uud4LlI+N5G82EqAn3Ida2ree60p80yG7QqaMYD3QaJ/h3QISCdr0YrUiFLI
Va7a+uqZLL5qq/OKjpn9Gy9opahWbAihVWwfWXEfuc25AmIeQZJLemH6eD4FDE/A
RG0u+gQE5vHn62E2mSIcDSjKhVA0wimweK6dDOPLnneBv1r2p6102CNqtLzoaIs9
T53/nLwizAhgbWIDPvRRPTlaeym5QyHfZlBWa7C2y3IV2f7kR/UG/g2r2NKIYDZU
Bw21N6Smc/EHapMVWBW2jfRQnSFWPU3ZDzEp3nnKBZnaLyAOfmxOSPh32YI8B9I+
37Ycz1e0YBwRCKKv/SBag0GA9WTuhfRQR1aVqQeUm/OwsCH35sM4J/FLU4fqSBD1
vJhE6pv158qg3cOct4VI7QDO2LIVdwImffV/riPelYiyOvZi2aZiTXjgoBNiiR9n
UpXq6rCyXPztPbGmR7iGhTxtnqqfjBOKQ7plPY7BVV+bwTpOjRxb8z6zH4WzSTgm
FqbtY9fdlxE2CUGZy/tgtm2ayFddpiO9OkeAHnv0TxUPxHjcrYvMqGblPk8xrED5
rACZjUFLs6ApOMvnE8Q5nqHXfFDQN6LlkndOVLvEZIYmKGw6Wtxw67Tydjg1SzAP
NSbk1C8Nk2Mm5XsZYrJxJ11pq8reXigL4WPPjfWe9d66PNA/FaxVS+DYzudoCk0V
Q6WOa0YClLPnxqXIcc48xSNfq7kOrM/0EWqWCOEE9/Lmunp3kbR0mfoETaBShRSk
JfgJQToZYDQR1J723/9XwzVF63MjjVC3AXsLsd5SM33ukyqzR4iOIcOQU+mlTxtA
zOkiWNmGllanG9s9rvMIb5lOX6IyrnfroFYHGlI1aDxiWh9cf67Ca2iFzmm10e0V
L91bAW7d6vUeZXUsfFPbdeX/PuhNTpplHkImrN2Jd/9B3hX+qSiMMtAtP40TXwnX
s6yzgF5oZYROG/dtozyY7hQ58vNGeBaJISAe1zi4j7G1t0ivRAVykZqFwiiiYV8Z
XAVBeWasNgSNqK9A4oJjaMr0wXj6E1fB6xZLNGNeC2Bn2yNrxzC5A0PH0sL2KD0T
gQ3zI4JHY1ccGoALb/bQ1r7mrmwSBYCvmE97vjpHb6qCjgh9eZ/IiR9g0VpV0Gcc
RP2TsJFEdOC0RO54PTE6GeYk36Mx6V/07+10PHHpSFoNqZimmn0YrFiaNp77O4qj
ka9PWsJcNnLYST7kbZcP+WlsHFzTdux/4/ouRuT//BAHs6Lg4ABrGf9UqLnBA/bO
jx5udbd+kE/s5u0Z++bEHYy2YTyg7+JcHdAJqLDEQP2NPJeKvSjFWdiPNdJAR/Nm
nawr2Tv5oGRVI94o0vYhXAC0k7Sx/X3F7LMggduJ14Wyr8qPytMGcUqE8JNJQc7L
4x33rSa2H2qbwES/RBmvRjMNddWcd3hWjdEnbi5ZIX5H8+34bXkdejG2dNVHHOQR
nnmI2XtfXp7A4w+/c8pd2iJr1Qu9Ab9oOw9JjKwpUb4gkNDpdvGpQpBbP7jMgnyZ
FUy3sYFvKhlLG3PRnAwAqckafocToilQYo1OzF4Cbo3UDtkyhle36enFId+kw/lz
a97CIzo2hYQaC17CvXU3RFRW0E7wEfr6qxo9Yr/RgeR0dN4rDVz4atAgxagnNVWo
TmR81Nixe9ZqyZ1jR/x8vV/sl9u3OWz5Fr50JOquHsd9INHy4CIy+yDrUIDMKPXM
hjhtb7QFeoVY1TnLJu8VMO8oOoAMuA/kRV7zF6h22dpkk6nayYjUDuMBJjfgmxDZ
3DIoRtBxkAItoQf+0gbJFazk2YTixRiLQAx2HoEb9UXL7tkMc297nEfEZibMcEr6
XRAkbLqzaYIQo6+h7R41MNa+n289+urTcx0hRMJGQcAibOWeGFeMy7qMBgAJm/al
uu0hmnD2YK9IzujZbIQ8qiixSjOwiG3TCOVj0BaqqthXQzw2EBw3pk+Otrl/Hys3
ByxLP5+JmaszTERtR3vrLhRJTVHnL4fWaTh4f5kUJm/AXHyMGKb/3uyF+cA5P/Pw
7A2YDrky0D2daqx69+gPPmjhE2AJC2mtDZYxCauLLmPiWUtPSPIi42UHSCxrDg53
1L/QAnOo/PLdZjpRMxwMChwHR5WEy3IAqFShtjb0CB5FOlWgHSDmDEOWeff7OISz
s4A1SLa+Vp2vEAE0QQwLmwzkzy/E91k7X55kGqCJD66oA4dYAZL+8aKkexgn0Pct
WYRxOA2yQnMerLwIEALw6z9mwNzUvFi5srK0e7/5ZBJ+nnInv600GMz3Tn2ZBWq4
3RoGen7fcXCx/Np+w27lMmsolol7SpExDi+5rhGZLuwZr+0Aj+af7Jyv3Q6P7tbk
uSDt9exRbCdwuIwjUJTmE2IUQlGP4BLl6NW3jWQU4h/5L2Q0prgMv/Jl1Rj/0FTu
RgUjTFg0JdUt73E/Npf7uPWveRlpMXTwfZqLI1sqWesk0frFJXkihX4CdLG77QOF
DCXEH4thka8fLhrmx/BzTX+uSwjKAP/m2+JXz7SizV8e2v3yTQ97NZPo8rN3CuPT
7J8hld66hwxIYZ1J4G5cuJ+GL8cklpphk5PaCCBEqS8Ulwv27wqu0yNbmzjkHYWL
tdhvc6MH7HWr21l3EEIoD2J2pEhmAV4S9ubiCIy6fIk8Mvjit9vkKQgFPFgef9gj
8/4Le+y1VDB7CAqk2vGArJtHZ9/S6s5vWG0m9qQtpg/EHBdSdekM8rnuQCUXKeS6
ur78f645mu00Wgm+hJSYJE27pmahBUbSjJkoUiBwj1by+1uSdlAe8ZBSTqMEtxnP
U614OvDnpj+huC5d2nAEWy9FNVmnn2Pa7BEeQXT3IUaoACRMkPuFwmY/B6KV5ED+
SLuMwkMa4MFO7MIT6IrOJB10I8rft+PX13ln4FkfkdGnryaoM+oNy39YY8UNDFWG
tiBu3qikMnB/LOXg7+PRqYLNOAvTSfrm+0sRL2L1zSI9hRC7FG8u0FSE+gbfVP0V
aotJ/ehZ3oMIOzgow97NUM+zkWntX5gutYQoy3U8J6fGYuo9Ezs2mx2jHnp9aWsI
67LEETLW4beAGGb3wR4fa6NTd/TyZTBHl932x3V0wcGoDxXpJm/37/OTvPTyoGAO
qsNXk2Pg/zzU5DzYwuH0WDOxQAMqaYOQ5h8ZNoHtBHT3orFT6EByyryOd7Ta4BWi
kFZTdmxPXSA0L4L7YKMFxR+a5cxeeB40V6LhPgnEE96chKVW5/MQjV2u64QdBo8q
YPDxwETOyq6YMu+JGMqobIU2a1XNrawGmj7ST3jajikZ7cZeeCycXFgCGkidCKZD
qwgZVLXYhp8tLhJj5l3U1Ui5sQmxtoBMLsJ50q9g3pXT9pIQetDatNT+7cube0fX
wg70x4IFGSttS99ej6lxvBvTr4PgE6uDMlFs2GPO3f9urKYjl3fvgJBfkdI1yZRH
gcZQVb20nH31z0r92t6tMYEKgaxplFwFCF5IuIiH0iZLQQ4IMLlKi5BaDGCVPkCy
dHLxN3AleH+mGDqPMEqlx/b/v3yNqctVIwxHNOJuGq8huXEgPMEC6WxvuG5pJxgG
FQt8JwR1inVFY4irvymcLAGU/NMTYKZQLjPxnjHdKn9SLbTjk/4l+fKPdsiNXmnv
4bt5E8M+2jgn5vkVtqjXqqKfgFHztMKA0joYwR9XCk1Nel9IfdRv0zIeJld54UUr
0WVNccA0QDrUkJKGUbIPLxdOtRxYr/1CGBGkvAKWEPtdg5bRyBT1IZBjq4N6r617
I/hyK/OQF4fHEogwIk/aL6dz39Bj4ZalxDHaOgvZAtreYOHJc0kmBBYqMf7m3bC3
RaH2USd5bzeIWkjzM+a0M4r4vURXunyGQ/Z9F5qIKcifSo1IzkefI+f5IzoBsWHe
kj6IbLr8L8oeShOraZMRL6Ie3Io+hpmnY0MWhk0Fr9rKdqz8CREXxQR9HmgyJqNA
vHkoEcXqTCk9Bt8wHXHVfn4Lb4OHcd2UngLTI/TN5yEE0ErQ0PHWMcuj4jns5dA9
0GuQC0ii4QG3qHe7ANdUBXaSX8G6jqDWZn185wrBtjV/P0tekGt71wU08YEgMEtI
R3KIU4xnHS2wKtZmTHkxWZK3hA6Z7uOuf9vTwgI64LTbyjYO3lftJWZm5Qja/GGy
7VDCJ/+EknMAG9cZ4qXcPl05Sc/fmoADfNbUdA5RGevowc08g4cW49O8zU4HsDG0
Gmdsj2aJ+TNuJWQ55FLTJTfp2UtiLzENsDFVE+GeYOROrTgrXTuahU0cYzxYYAv+
o0AlDrRVyfT2yGs+GKDLzwg1NQT+Glu4YvjBdwjunCZk9zNuCogC0f0vgMrT0oKN
X+gKZ43rw55u71VCbreKC1ROf29p1BNkSSejzyM+4PCMhALNBH5eYfpsy0gXJGt/
oR2G2leNE6OScNw7a6ugNMvZ33q8lTCbGFgNPs0bPMyblT6vlmWoV95AxF4K/DiR
xi8KsmY7jWWB2nenDyWkGssboY44c8WTlyfOXlE4xes8giE5qzrh0kaajYsbWsJG
qK9Dtf9K42QoVXHmpC5rLpuoF5FC5Gy56lNymBXiimtWSs2dgpq0dft0tIO3vfTf
enuOTIAEGaQTUwRcvCrz0f+vgO+0P8RLjlRIX2nHCJKSjV5sIx2gg45+cS8ezk0Y
dmLTINLbCF4HUIABKue06Wus0C0BbEtbNRi15LKVw882wFx47g2T1aR3RM9oPHkU
SiP/eXyMzbYzuc5JVVDix2QDIw2T4vn8GnAG3t8sZ0uMAhJAr8v8SiG/CD5cVBGa
I7fbp/ceSUHpLY7ma2wNrDSM+GKmgNnwTKRqt0eFhleJCd1xzbuSK5ZydUpw3DE8
azV/nt1HCYclGlh0g+IjrYXltOBBkTyk7XZn3fMR6cI94VRD0b37pi25BLrtAqxk
k9z4rstpuvJg7/pGYM5PB2sLiN84ml94QVDOu6PEtdyZavjReXzH9JmmwXrB+m80
pXxH5DqY551Zg/aSOZeVYIne4eMP+bNHDGhtr/BSef2s2d6+tQjT67rlIo5XVSxn
Qu9xJwJIX0b+AUrLeBYw2VE5dZcaWf6HrEDi/i3MzDQfT60IIEv3PssFNuD1OGMI
ExDGhzXKGhkIAO9zu4cP4WokXfkU4H1B+DDdTZS8HiNs5u0+BUk1dgfpHsXfObbj
Su05dU7dTZ1m2M933uXAaZhLb09NpXz2YestZeWYDI7ZTQaOvSZYogSQob+OykC/
rme7qZEmhPZoGCTUQTck+f2h+o098llkraNUciLRKJX6W6cSgJPUO7OvGN9zhGx0
dxNwRrGgRJKpUVoT4ixPodCcpRhkwrT5YCo4ZdQYrkkFqwkewChU7CXtIn1n3QUW
H8AAOVAPJ3TNxvJovNS7UynKzUw5RnQk01Gjkwu9CbU2J/K1NvRlKlx/5LYqbcwO
nTnaABtV2qBm0rTfmBxM7TtMjMsRV0c/eWgKIsxToC0V7y9Qlf3BH2OPKI1GsEYP
P202xZoho3ELTT+NgWm1KiBPuoeHPEdfXN05UWAzOuVnL97H0Bew8KHoIwgHk2zl
dj7QxeBUn8gMSqt8jzGzwRPxTDJNVcQZqW5bbzT5GnjsV3eiO1Fm/SVHzpx8HTrj
iHcptV+BzHOWgp8aMcsGoK44DA/P/LChi1mPJtU7zkN6H1kpBH/JdWcXJT+B+sVD
JXXgSgAfr2+2GCNK6M5dmrInOOkCdmAWkvr/F1e1RXzowjpNhA/dy1KW8dthWHms
efipElAPHZikxtLSuFf121M7mLrOmTgJVdyEqXTguJLMNshSJ42AW+hZOnUNzPNV
uf1ybnpRbvYp4/0Zy1I7MdSFFK8V4ZVHCPHObuuFoZiLTMTBEyzY+zJnKdWzjsA9
XmtJakTloFL15XH74kKnFYib/MyPB8AWFgq1hrDoz7iR1mPiexwQdSUpWEbVRFyV
Iuu6bdlY68EXjHbr4Qv/mbidH13ewKdpk4NSFcKNtV6Ag9Vyn1dgXCMV2jdV8FPv
yR1DrTsb4BOEpl0lQ+6tPu5iPWWHmcBMiF5b7fc3JLgsPwbvmN6Xjm3rPnvoF5nM
/JayGK1r86NpSPq5Sw+DOGcHUST/8yr/+Pszo5q4aCUtPRwMCY1dopaTfAyKQwpY
oCvmZdeDUQp+al0P2f6dUd8O9iT2NIvu/5lKXeTIdY2YaEwL+WiCnjkuyGrWOxrL
7INGeTc2VbI+AG1Sx/5OelH5I2fbeWioGmMyv8IyO5jkuTvnKtmWBB23bBPB7QXh
yABehk1rq6TFRwv2ybA+ibR10VP6syK5Hsz1U/j4q9FNUyYFQrRjlh4XQCtLK8t8
05iARWjfEBHl+x/aYXfiZkSBRsmfEusLTEox5TNwr9iOtnKooCGSvI8tKDkVDqlw
ADAK/F1IdJcOR/K93TzeArEUJVaxBDFmGi++fxotUnZj/grDH7/B+dncse+6tvAf
eFJHrCauI3ulLvAbhTAVqfgvWWgDV3JktndJb56dI3vK3uSrhp5dNj0fLFAn/PrS
F4dUWnMeZ2VoNjXvFlPLPbgz0dDEZDQt4vXKUvl56c47b9Y2CeHC8Pb3xkLD8ODZ
PP2BOOLuuPYVN2ct7QNu6BJRAYK2jVB60yoSzE4OXXUgvYXOoIVCw3hadd3IOAdH
8jCz13ujctYvjht5BBiMEC+2g+ZjSdoINcTT70K73BJso6X4qL95h67ZxbGn6MWK
rJs/wKTfGFVAEhwYWsuBrGiOv8vlVS2v3oYR0tcdrn4CmSAhPZtFcjyDLMFOnc/w
fcfkJhN8xUXyp+W3IafVeVCviLsq6jWwUzPybVHpuqn849k9l3Px+aaE9rZvFLXb
m4Izqyb/I3GDD0Xk0pfJhmUmeDWikFYg/Z8agjz76Wod5oPtPRiPxp2n7r4OckXy
GBQiEJaPHCHRAhEeV0vsRoS6WADM0/yvQZLJoZ1Pd4Ocp5JNMUlofzemNM2uRNuq
46iWWOSpPbn1WbT2f1+zNfVgTfaYERTB8LFnp4oUDarpHk8gy6LyF7mtby6l6NZS
VlgwhyYbF8NEqONXnDeEY3AP3WJm+kUAOm+PLFtpN+QXDsShT19ceFhKOHOk2x6V
73VeU1EJTUafoDqjErZ4ffwlxAXc4G9mPOnAolUIm+kgZ32QdDe5syJ7v5HTvhOX
UlYZOXtyV13wHF3h9eEVzSDEaF59Paw/F5pzF3iPGvHlsW/7cr+y6rlM5fzV0Udk
cKweVvaIQqtjUVS7xvr6+hE74PnTfTqUjGxMGwdsQSriBjqYi5W7imYCnKwyqbVX
YPfaRE43RAr9gDW4fj6b8Dgm6wnogxIvnEUrfDnMwfPEDtM6tA7vYU9ggdQ+IUpE
74ufgY99tpMREsslEbU13kaV7tQi6/UpVLDOKtOsAK7J/U+mV+jfL0tmAn3/QQWy
qD46N9w8oBqLoaMuKDp/4Yxh4go02L2mhKRVA71d7uL/Uqkm1qU7R9qalApRmIG2
Zl2MPI0UQOMgLezY2g70dH3vJU5wep+Y6H57DjkrDvHmvsHCwkSaWbUu8U3h+WkI
PHuh5UUeSVg3eqAWUHzPqy09ZemiqvmwE324h9EghyJ4eoCfH0Af8+lMjiSMBjOS
dhxz4SR03HsTU0H4e55Qs7gFSqcPd6DE7BgBUcdKW5evHjZi/Js6Cc+h5Xuw+3lG
SPckW9MJQ71POmLHsVnTdwJH1lys2xw2uGVBEGcZAenPf/C80brYR9kBCmSllncF
jC2Gg0Xe76z3WCNi/MVOtxNb/mXqyhSQMrvt5Y/6eDjbhDfaszKW5zBtvz/T1yW3
iXqQ0W+I7u+op42WmQSdKs26a6ccSMpambWrkU9KDyRyZoJXQTeJDxvtCVQjW95l
pdeJZxfjx4AOSPcxS/v/B5M/EVIUk4byZLWPAURy9due057c9N9z5jZdY+NOpNm/
lzwiRZ8dWlLqebU3WBg8hCKktSGg9LRUyaW2yZLXQjITyu4SejFDHH0ZdHtJ9mUC
ijog5tKzB6boEMP5QDXFRgUw+7c2GnztdyuTZ4AvAslOoL2h4FK8E1sDtH97rhZW
BYi2hNHV/ULlckhT5Cgt4t37iULhHYI0qmmQquL6n2cASGPqdfN4B3GBRqgxv7vL
/AhTfTl9yY79vXVW3f0/KQQnbK//Mo3pp8zZ1PiLQenEgf9qfmGO948BIYhxhAYE
fsGUdsX+g/Gk3ZqBlJ/uPJNPVLMappUn0VzzD7ikrcHeK7PINBC5nZd/3+nVtvJ0
halT7Uyb+kstgvzeU0/9dAUdnjRv8NRn+PAm6EnERa8lSC4u1/bQ9vIptZhYaP9y
PyWW8tJPHxZFeEsmR0asiwRhnitiMBrChoKQI8Ezc58K0etNQ/fcgzyw3TUlTjdi
V/HQti1oy6754b6VSZco8kQ1whCwNe/2xHns4fE/Le95CnVLOa8MlOcn3TsspSXa
Uf5xIJBC3WKVuHpeYG7VblwHqQORiwFb0iX1Uae5vhZxy0EyVl+/NyVjGrr9n7jY
gmB/7t+J7ChNky+Wk6oBi/nn3C0YSXZYm95QeN3zX8b2/SUBFWVjvt66VU77ozcA
9uhKUZT9+A23p9JchzG8G3ONsDhR/RPml8TcPgLdPNITTy/8D0Wq1LwgiBlt1Ir5
+6P1joa+WRwO0zSMnQzeeej38ULODn1XT9hAW1o2e4MnVHVXujzwkfjbY6Po9Kl8
Bd76t6436L2xZlaSO0OW2+y/s9tysg4RAu7po9s15jSX2s8Tp6kqEiMjH55BqKI1
3kp/HTljvRMZ2TtNpL+b8MDonpPuASHLXS5YExoyYxOxSLLZcPj9Xr2/9WlbWJUT
AaSIz+jyV82ezNJAcOm87Yuw3gDVq7NHt1/Oe/8jeI6RzOPUyJ81ByncY8z1gl13
Qs+FL7yOgkzdMIgJzmP51MuWhSbUBxKuY3zvxPIDUbst1ptg9vgEP0thbs4PgT+e
NYmikrgDZqYpSGr+70EneDcwprbzGjKZb4riq32AOpU/uNQHEvZHnDIHnNI0e5ex
GFFqU4NAoFNTFZxf06Ku15NLKZqcyPFO/aIJXBnPrEUw0WvAy8KBUifjgSzZ9iJa
7PNifpTmCMHira50W3mxEGIC+MMutce+NxhTsUsUQ+iaWzbfmO26+P4gkirXt41o
aRoGsaffbZlFzYgWMiTVAp86bxrjOsINiLxy4LmfJHCAedxFSaQp4eG+GCGhrqzl
tPGXKrw1JK3xOgvZVjiW24jxk6dTOqNofSa5gS+8HeeomridV6WmwJ8M5hz50LWz
dXQwT22vwF/e5KSM6BZPvyiTZDTlajva7Oz6Go5SbrktnJ2ueqsGMCQaywJ2DbvP
ZBlha227EaxnwmhepLSwH0v40bLsgzufqnhrvE9KUVxXGGWV4+kwDZe7zs5X8Xwq
VCvRtSrpuipo9QGvR7Gq1FVv3jEY+p03jgPlwS1CjNzTuI7gtLzo3Oz8fTU2cMl5
qhDHOujvD566EsPkZQ2wZ6714MW3dwiPKdSTbgFCGVYeJolrXWZs3TMsGB7qoh+0
pVmTYBU0xrXtAzp6XLuHl66r4QKL8+Oppn/h5mMykZL3f2exOLbF0CLnB2961eLV
tQzGh7XelrYjI4lvUyip9EfTlD0MmVJxo72vPxTOC1m3ObCPdov5PglobB9JO73i
9Ay/UTo58fERpXpfLDiritXDCGC+FtD5Hs706zg1IXRxnIwoRRcsAf1p+AeJU8Xa
oaGs3iR9YXCdF5pq0cM8hMqSSjNWBpKUWb4jQzU6QphdJwwiPBsTvHIHe9GSm1QM
xboW289e2yYVv0mw3Tfly69U4gHOZf7iVxZaQArqKQL0hqqq3wR17rTlJuAVWLyb
GEq+QOKV0LZf/b1Y/C1ByXD9tXdAkAe30j0PIEOivaAOjpr8MC3qZgo1DkICczmk
iyJErRuqY0ZPpXbozZJkEVyH8GmSYQ/fpKXa/DGt9LZZ/62Tz7f9uORb4SgQyxeG
afKcEu/6SeUZgYmER/uwUzrnAox3aGcce8RNQTkgmAqXhdJOl6kQ9Um/qoZ4ir0p
iD3gPYAvHliJ46zKXXO3j8tif1YMxHZaJPt0doCkTrhDLTi/9jZuiHU4wE+b6qZC
w8Di+K2l5FeqUAYMIm/3r9NzqHXqR9n4P6JVQtUHQo2f0oyGR5RAQW0ORAeHZ9/Q
jIFH4Bb2lARfrs89WLtxPHLirTpEbBGqPNRhfl6JPF2HU8TkzipFPiAF6oyPnx6h
CECfZ0kwUJ3/PzV0r9b3Ppo19aIEttd5JQhlL9FTsww+OJQN80Z6TxfLjPV5CwW9
4JtBkMAwp0/Ua/7Ot9U3Ek9r3+ADGWHj2GSpysW7n6HBuB4UKGffHEr/8VTD5KrI
106vEiR5fpBnslZqmgqBI3ipoSkqY2XS63qjIVBJFm/4jdAoz4IS+W3XWwOLmMXl
DLYB1XCf2WBRyzoizE3/2nz1BwvMsM5ktX0QMW/KjEstZL1+kkJlORTvoe0RDJW5
/olcWDRoHcfqCQ5f8/rXGY2kwpUDBZghX45+BG286yzV6S4b5VolNOpLUCmDw955
cAzwqXhTUC88bkB2dD5nmiCy0JqdyM+e6XtIUzWeefYT2Z3cuOlPKv3PO2iCtDT5
d4TBMRUynln3DbMb46oIs453Knjt+6FnR16K7b2OrspaWL/yeHnbrFg3PrZ2LXoX
sWh/gfX35mSUyJ5oUFpfzXsdGiR7w8DHp1G3flpS+Gi4JTpXrp9uML4UylC9LMkW
HR3tfZOIu87rbPTkyhxvhN+IPYM1EhXamixhnfBVdWvMxoINuFLKP4bgsofBGUmn
/sV6dxdJDaGHd8WlmM0X3tFXvYRzUCL9j70rK5GN8mMdCH85wr8T2U+TDi1XK4p8
cUjN+90zAPvNFoi4sn4PLLk4QQH8HMbtG8OLDzQ0XX2U1l3y54to3lCTjf7sLJUq
vRzAYj1/frmbeOtf9sTSkgtlyGy/slpzw2J+oKgwiC77CFdSldz1SzPfKYJjAPSd
QvzOKkPFdhchOrudSznkYtCVAM5y9XqHEbSC9pw94ZYLMlOkjnHuzQsZ54ECNzSk
NcqYHJQg7rcX+YGQROVp5iEoDjz1a4fsqbzNscsEpWLpNuq/oU82Zv2VnpPcq5gt
4cStVWP/lFPz+DrF+3FXNyqjKVKObuDPHlRwcAZ8c5cykqFyqphmhUtPTr0grYgO
hfWjn90XHlDx7x82cm+doj2/hxCL3ax0rvRXJZaBmbbt30Q57bwbN2gCioCQBtQ+
LxubSqtZpIUfGqnHnJUTSRzF7Ar2DgnHgYUy/bskWb0rilThqS83iwwo2KQ9xr96
u80uXigF5ZbqeIj+T0BShlFkyYbOxLAMPlQZkWkpMY9D/lMkq7yr9UJbZf+bKtgZ
teNYkqlyJaeDe3Wy5E+gxvULTEPT63fsgCLV4x7V9sz1+aXgP7VZXY4pBDMaeFFU
Ir+0IBMwkmEEG+eTLx7PDNpFbdzZhN/HmPZe/3Ls5RlnB8DpkMLiLLto7T4bBZqZ
yv+vpthXla7uIsdwZQGJGusrK6X4rz/zJ9pooYza7RqH3sWGLLP5vfMhAxtLwx/d
qiXt5hgl4KhgxgzIULkXL+kaccDwk/mNWYBjESunuBoFa6EDpa+w0DdGyzSvPVj3
XxRUC+dMyu+D0KmE3+QgzuO0UBxnFFsVDriKmG0VbqsKvakoboXSvAfULZXUEztQ
kWMkbhImhjyhrPTq+mg2UaAcdiVC3QjF1POKZaiHeMQsaN3ddCkxmRC7YmNDlucc
riJCYSmI1VDtbgwhRBamHp2XJPhNU16KarZIZzm/dwh5qvLwlIXMJPuAQKoApIyg
3zgp9XlGS2CwBs/ubK/RM213T2GufnvzEGrftIdTLGGUzIt8cIcdmANHSBH4ny44
e7uns8y0564OsGk+DeUqhRnsa2DUZGdjn0MAU13DT3YpbaAI7xfx0rOJaXE1v0Rc
IZCwCLpYv3Dr9VWcsuZ4aC+11X4VXzirmxTakTay/NfJ8xNynnG22no0Zvn/6mVt
F8X7Ue08ImL/0NunqK+G7WMOn/3XPq56Sq59cLqDHeoEhjdswvhyssaHN5+tUq3I
BqSkQpu+5J5gx/suCDKNSTWcsDwiq2iyab3kYtkZSeRK0kU7Uj8+MmyEer5vkfsF
gn4xTfda5001Pjj+QwiSrkdvjDsytGxElL6dfO8Sv8gBpywRGr/JhMee7dbun2lu
wAf3SLFUQDgVKK47AzsGEIn7Z+UBZ5j/ZVJcgBWlMW1u0gqpQWpIXZcPvUFTO6nK
umZvoLln0/gNGRGHrGDUrVk3EPNr+MdqQExaMVgcadEUqsHI2iEneny3Sqf6oRzp
3TwoDEOl09Qi4cm+OmRNOREB8SF7HQV3XHki8MjJPi5KfSqdijaSqP0hFC0OU6/d
w8BQBkvPzT19d7FyH8plHwojZ8BJeI/kScEcN7/QVzre52vjIUmAc2PGk32jm1sz
oPEK/I6XMUhSC429yzKqTxr7aWgIzOUCWeNZbOLk23BpHRYlHK6wnXM4Nh9n0y/9
cXYH/uO0fF/1WTJx3r+RVypo9SVWmj72h7pQicWv1/aIYWW2VQLeuJre6pzc9gSv
uzsziOaAKnqkvxqyIRH4GO5qwxiZHT0UhEOLemMYUS2++YdE6mm9RGxoFNKc2SHV
sCzoRvCk6wVxKwANi2ZTtOXOLOWzlM+qPyIlR/q3adgOCey37n6gmx7s4p2PmQl3
af2GRRcAM2ID/HwAf3/xfbCX3RIP2KnIb2cejGJuoigUNhTF82eIP0Vt6ksdHUTc
f8c0sB3C+dFOl2cFeZ0//Zmp0GiMM2NVAHAPCjxx57D2RI35D7T3vl2OCufmv98n
SMtG2vZduNQX+ENW/b5mrk1NEslhZCk6+uBNMCV7x2L+2sThrL7KPIj6ZmmY6R4q
T6/FovMpMl8bKG3PXwjcaIAW3/niMOHNrHb5fto7QA1TIez5SQRoI2yht6uZ5VE/
jmVh/z+DMR/3RsWgeCLtNn5peCXlm+rpfawEWbvXBX+YwzIx909t3XNHZ5rv7HtF
45hxrnVzlpcv0nbT7dlJsaBAaz/xePRT0nkrtl9v8mySYw2CaEATDZCJIfT3dy6k
T7mQ/sTP61i6zqkKH/p3NW91DRgu3gD05xPvyZeS0Imp9+7ih2LaHJipbOgfhDHo
xbGxFHUpkgnrzHO1oNIDNa1foM9EAw89pHBqOWoIM2OJYb+z0T7L95/9qZURSu1s
4sRnhoYfLbpxoXr4xKfAMiC8aKiF+hKwKXKw25xB57EeJgT9fY9Yho99Aip2wwTB
ALlNnMSUBWnCvA33Za3PrMM96xWRVHn2wvpiRc3kpduObxP1YIleWD7l83O28PYa
OOtOxnWmyh4K7yCpkwlgBym40PYPRDGKdILjBLOrzhZNZso9Uv/umWdE4cCfqsPm
vmttjN3HvXDT8gDBdwv7ooKUYfKx1TU1fuTFapWPvQiZEmJ9IoSZkKG5RzOB/1fW
x9+O7iWU20xC7PngcYlp+4izghM+XxLjK9PsSoaOwXaenSEmPWd1YMYvZlIn42v0
Z4Z9vWrwSjTmqyI1PQVJwXFIym+EHSdKxOSqCTakgvQBZ55Ak/nQWUjxIhVYuavm
jdiYpJ9eTHZjKZD/bOBNkYG+o/PuIGRiAWNmuWZVlThWnlQfsclcBACLUj6GKZYg
dOAPs/jHsP8vxq7Qfeewr/4gGZQzV7ym7xYeXWP8C2TBcUdk12v/Beph2nUmvPDc
hfeRRtlF0JjA5PdfDh1YLP26O0A6AQeDHP7h/5ZTJOFZixJF5Kecx+ksR5LXxFNi
cSOXRP4/me4K0Jt+O+NoOZGNWuHCg9FfyxN2TO8GWDoPnzgton4Bq+gt6P/Y3wXx
LS6uZ+O5w4d7lJXQWLf3iYYtEsU0uPaO0acG59eENwrppBgRj4itROgKPjAOFGID
qSLWvhKKE5SuMbxbCXWzSlp/ySoyqog1ahM2PWQJJgsPzQFSMrVe96+HoU6Dl8FE
x/PMjSHFnogNdj4mHQJEWudt/KnFu6VC7m5TotNK010MlKfS+LnFUyHzyyRtpepC
AhvfAwW9KB0BYgaiKhJhUPTUxpK3TPpE3GwIzMc66eNrqk5XVvk8PBLkUi4i4xtw
Lg3XS+6IaVxr+2G8x0y3VxKxWtxL1w8VYCIW1g9qY/j2nwmZMfRcuWZ6oeVVFvC9
mGyYgh0Ks2IWl++3dVpYz1vdCo8GZe1tJfJ+OqdrdDhAHHaFKqcK9ZY3t1+uq708
AIQrVIyPO/kkRrTF9kJomDi3ipw1sfYK+2l9tG+tmzwEYIrDnkxMgmsFoUVH9u8h
gieYPHtVD1KN+U6ZF0SY20cEnTqiRSVEW/JqRP0ADAhqMOFvYBGqeD8SpF2ghxBH
rzmnj9Y8lNID4xgJPwnglCGSZwE2GK4R0r9R3GcsRifOdlPHgiTS1jWbs13v6Gg+
nu+7FkKKhia1Aky4Nw82yX1QWdIM7iWhGbLGCskCCTP5Vi8EUGBGDL8BWVroJkVE
dH+wnt83xNYH31/k50/4mTZyxOwMlFsqeQxlZyIxsdzsQVnWlxZAWuadLkejfi5b
qp5WMtj2psx9zkkbEogGXxQuaEv4/VEWFsaXLRsVFE7vZL/AE4EO73dEUx9v2x1P
J3xnX4oSkmsjmCrFoc9cutdQbR+NVGn9FfvMUoTlS2om3IH9+qrpH0CsVCBW3c9z
5lp+/2akAMVHqeqAkPCIFN5DZwdqPhaFx4ZEuZtgz0ermJk3tFJujPThFbk0IzxQ
hNmNo2a+oMBpKmYe4ZN2dQMPO+sf9Ubro5rS+lZZhFWpYOAQQy7b3NrDUZm4vmus
9+BS5xBZpy6BAdGC1q0BdIPnX2McmvhRy6tECMvKnotSbfk4nTQXqAFS2Z4XCOt0
RJkUAMojBA9TmW+yihxPjc6tMTlzUzW2QuBG4hlBIVdD/a1vRnklTAA/Y239+FFB
QK1m6z34cAJ4d7hRko+pH+9GnXw36tuK0Y+8OVncjV8NFis9BpPAahKh0Y2T8QI4
8mHvi05VOYbi027MYikVsVzx2BMAHbJeNElqCg7s3QH6D4OYCBjutG12Zo+lvN2i
qzE/6jxIXkdE+7GaJL0RhpJ+dAu2irF6LazqJawaA1BM7JhPBNL0X1MO27Iv9J5T
WfU13+2YjDiWkrVRiLIJ8KRE1aJZTqVAQRlLPAwGeJzehgwKPqH+1wjc+ch0OGi7
mBydgaRmrs0o2nSrlUq0nUc64eojxqCO3eHz6ov91ICkDJ+Z8/cpK/Sf8FwZsaL0
Lw/F+eftpWy95M+dsAiOgZQ8+w509a06/+20dF/nH3qOOqwQJSZm73W3qtz6+bhP
jlgYEJ4VD6uaLNp5KZ90zsOzT/r4orS4pwX/VVupY5OlffCWxFTECWPabJIS5gAP
oVOt1gxd1ns7OZyAOzbV4LAgG6/LOSbru7FKlTrHG5KZzUKZh0Ruut0hOMspn8L4
eSUHaqdKjH7nD3uIESB1/1w4IxlDJG/IIixDJApEYGivM3XDPCkDIo1BSspgITUT
MFe017ZNBqqsu2ym/SQip7mDYxVpxpJ4x2KraNZyRQJ9Qeizt2itr7LpYFa5wY9P
ycKdZvZlKpPbaxIyvJANIM57OBuTERkWLVPzG889UCoC/MraDQvqx5xwJ/7lDkE0
m9Oww2C99wond6QtLfq3gT3PA1UPWv07uQoyhJ44npF+mbAQWORE70wzHeC3vxvi
ODgyQUoNk7BSOtUSNoBAJv8FS5k6EFtHveCLi3qG5JUrdIEJOfyoBIWMOSNNHNj6
NiMV9ga7HrmcDvoD6SlR+25hIhcP8VmUwlWVnmUKzFNOlJ+IAfyn3LgNKl7b5xlR
7aNpRpKpOhJRDwryqzIqhGg7b7Gh2FkLEK/1S6FDviJe/6NNoQGUcaff8eSvCNk5
tjsGbv6tU8BinWphi/Z43x8zGJzIUU9mkDYtEMwqSXaay6fTjsziBA2lhMW3sTYk
nGS2LG28YMPyIKBo6tTlu4BXUC9SkbuY232WKOF/bBtHtxat8rurKRZ3uXFxlYUF
HR/KWKjVFTcwxseDxyuXmoMFsTcEe45I1QvSOaunz/Y2GrYCMyO+7OI/Zct3wz0T
7MJKe6Y9Gkaouj/BT33qEjWcHMtejePI+kh4Q+P2ulD8dHt3P/7HeKcB6nl1E3Kl
0VfE/YEAe3Cj9Z66QZ2ecK0aIfMPOM/RunLt4tPHuK9roWzBZoDaVndmfDCJ4GzA
zUiV1uJ01D2QDuKhNO8HI7VZ0arNAFkeRK4FnMVRBXvCHKm4zc+iGS5vLAw+/GbY
oWE6OaSnKPLbLnRpuwXimDnxDnFgx66lXOaLz8BWwEBy/+QZi4lQMOV445UbQDnP
krmPci9Xhzv7ORGpaoxkoNCLJPAvTy7dordSdoskZY/6SCnFMQh4V2zulD4u/Dxq
bo9voLfHGsr1KxA/tqpDej1k+tvU9+FHAqdkoMLxrc2JQqUHaFxaQL2G27/T4XlX
RNSOajiFvNuhHOpkRMsqY5u5TCmAr1L4D1soxZRCVL6CZqqQdBKa7VvcpULRzprF
VmJlqDFCUy1uGuPUayKBw3VSBq9K6KvOuOJlyGDXunGVXkGmVsBp0kEkmSQIeHJn
3djeuSxflRQNm6PYFUWIqXtNlsUQd11HXi83LJxMwXbxZAEsXIRKSC/L60M4WJzd
7mqRRr34hl8xe0va2dFlR8Ond4d0d6SQcyAz1hT7yaorDcDYbVkeAyjGke3bjwac
F14AisO1hyu2v/UbiCzkQ6mq6ZahbiqCkBxFMBcgp+LQPCmfMIubgxlDxsGcqCwd
zbsv8bZ7pK9sTjTAc3cG8tgV0UwxIC8GRHALjTJ3LG06oaj0HJOFzJH3EG/4nMX2
bmcO67j0uhSoE3kMrjveNJNNEuQ4TzUgjg/eB0MU5enS71GnwOX6oy8Lm4tWkhBt
Otw5KczZ6AlhTIgwP/4EfVdTizsLeflJlD9ScBpo/zFrudDGXpHes9aLIuQqj777
/kWStH2EtUyijeRpx3UQGbi6ajHOXMfzex2cufHGdgAoVehCMfmAaamf+JwhbOMo
X4PcAbJth1TLQ5sQwG0oOg==
`pragma protect end_protected
