// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tSge0Q2w+FLfNGkMUDi/eFgpX15YC8frMGxAbxn6olgOSOsM6Jy8Q0LJJZj6jHlh
z4kTRKGoXKg+ty7bN+dWfGILDtpnWd9STwNphdGgPnjCXBA8m5vsCrCSIYPinaOs
SHyp4JdNqSFeuUTPj+HG479HvGL2reQa6UDPMVBqv3g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4912)
Z7xSfzF6AWgLTRcPRq23QsE50iqGI5Pfj+Z2/tCQpoPlrMYFjA+/ekwGPcJib9Yu
KIWr3RxUw9LwjNeAUc2TKA+FdbSvFCPA+VKwGExZc6SQe7Sn0v4jHjiktxKD47LU
OLf10CLGpjoj8f/0CAJO13XaVsZ0RUJFdLaYw6+EffKtDbKXyAfs3lHLZVMl82Ry
eJZH/kj0DR6djJ7tHk8/E8aY+3R4/j9A+iBZonQ4pwP4SzDIRPXhQ7NhFz6tbFgw
0JIDxmMuOMq1YmfE5K0Mif4E/oxlKAZxqs4DpWf7+hqb/mWUlKy0lRNxyckQGjBE
1ILytj3Oyq8CCsRY8Zn1BHGL56mzzj2QujDkEKsjjTLQcTHW7stg5RVu4UZOLGWf
oCVlcVjDZ+E5IYY9hcnvlQT84mV8zew++yStrxQS+EKrDpbjC+6V5clpe7vlTSSK
u7ouNOg0h1ne0cNyJjHd9kr7ypWDmILm5w+MJGjh0fRc5PXLpWek5A3GzG8DRzVV
OCehjsVur79fGpfXztocbFLZm2i4dS+fBFn02nPETZAszrbmkvgR6pccLZKTOVGB
oIEjB2FEF2R4CuKI3dnSTMGPG/Z3hHLRmpjoTTg7sqZl5i0ugqJSgV5oLhbIyVOf
5/Or5+Hkx+mM9nZX4y42I1XmJZenbwCvK8bTuKPuRY49e1CGI6FfHAPH3mgno9n3
IISUKUUbP9caMO2uWiMme1i5Svve+KX+yvH9fAGlNjwpcQonT0DExkx4F3wVS6rr
dXU1GNEHikE9Iu+L0mxOotAXp+FiaMjOmPX63lL4FIyaqs99stUdl86CXov4IEUE
s/o0QLLB1m4DSaXw9o794H8N2G07CYcd0tVGD3TJQbmiwSEdHUSbhTscDpsYrR1O
xU255X9RkIBbu8dEC6oSlpJjyB49L9/ASmGUGkphFsQL1GSTfQb5oVL8fRkaIro1
gvN8L9Zo2SCIL01QEN+LUa7YxJYdC+RFBFf+1yTXCgRyVZf1kU4YjE1DtMb/Z9Yg
VfudWTvkOQEtyKJlffm3/upjSOOalHEMOxuR0FZ+ta97e0XEL2AnqnFPrHHUKbQu
wgT83b9hkOiHSbby3DiEjv46SQDJ50XzMJ/6usFhkPACUdJQ1znWxk3kZYp1bG1y
YOlz9W0aL+y/liV/+lPSaUxo9ggF4SykT06+Wd2iaus3h7fj36cANKFivJIMdArD
7HCIJgelvOyYDJgoxo1TUFeIzr1Ee3Xx3eMcVU21Pw00ojYolcUhduHDwUHgY6KO
HlvicJZgFfq8jEqXTBAIdXQ3NajHJ2rwXTpg4TnzP5V+kTEKELl99aViB3ng/3wZ
oTOEBZYzvlRo2btOxFUXT8+0fSwr6L6QnKLorjBR/eL03q7wF9brSnDxt8tZN38A
GHNmqvELb9zBHUVcgACBchm1C0Z0KuC5H5mKBcXgTOggTDZmVqrbRAa9+/hWOkax
/3M5f2xp47JOw3Se9Jn/imTu18fDTRO692b7DLd03WQT4h1eOtnUIvb47OTKHj8C
a2R6+jXQK6Uuh1VdL9ok04remQC2KhXN3UG6MKW5CGTAamp0iRN8JKJB904yXO4k
x+j520vf/Pw5T6nEHNni80KEmb4T6Jki8GbH/407eqTV6L9aYd6h5AKGyKIRpsiH
rPyMk4krjNCnCEeYCtzMiCLKvxFbKZrRiLN2wKc+1XmxV9pKYI8itzDhR4eFmg1/
M+dK+Tbhc1I4j6s2WnSKHE+x6LI8grzXL2iJcVXMExSi+FxnnN9oQPBnMQNg4M8i
p9HMeqi0qMG4RkEGYZTz4zetK1j5542fQhhGWbSOy5EFQy7PCI+YWVoLbD8LZv4p
/Au36+fUUDMnF+jZ360ClWOQZUYnTX/Ap+41IiRWTtJjKBMQDtAXnODnC4VlDodL
1acvF+h6EnhlKg0xMmO7B3prB2bFHL1LuzLcE+WXNWL1+XimFevUn0DfpPttRKJA
24CSU2gQDPlZnyz9ZdjzpUxy+G0J5kLmAm+h9hFqTxLqISltvO8tmIztU4FIOHXd
mG+P9l+FkwzrPzqmM9HgqlPLIYp8E6TdVC627iqJq7LgyKzgAkKywW+/ZfEpq0xS
KEwQ6BAvic5iqtqGY89ujOCnIz+DI2y01oTzkOsQ70bH2BPvzKL56SZo0Ej8lFlw
kbVeh6KZNseA3LYiAtoWidZOSyyrJi4hYULpgJv7cBETmSzN+h4dI/Urx4EuWmDL
RRajf2XlxnMQU8DlCq1la9BWRejBwHTYab993dO+dTahcYFfoWwpPK8DV7DEkVio
WA0SBLhHVHDXaQyJUvegB9+EuPsl80E0d3wfABZnHiPSXEle9Q6ylrXQ2odL4Jyn
MR/M6EXfhcLpNjMtLlT9sf8guky+pI822kvvPVueu11xc0sTUTGvD6bjgzfrzXdZ
priW24veM9lBVmdInQTkNexoWOqYlZYelUbepvRodli/YuXTEAbVoNEWWDJ1GlPj
aezaopDjO+6UnOgov3RQmrgpDj+4Oaj/tsSj5Go2FhqiGXNa2/Jil4iNpWYA3D2V
0mz3qqjKzYaxQw4nAOkeqJxF8eUcBJq1WAVjgOTnXT+uxnechRKXJsjUXACFl1Gp
sj2UCjRro2govGeaWkEl6mBURgVDEdT2RDqc2/7scg8lIl6dUGsN/g374Gxwm8fh
1UwlseDzLEQJt+yRrF/UKCBPoy05mYPw1Rrn2raiaF5FYv9i2QPxIyRZ+m1xm+L3
fvVWgG4AUfA0UPnHRyKcCJ7Y8hL/hULb0gzK0YLnVfIFTcdfNFqAQjJ3g3Aa5Ewk
g0tlouaScKBUvfQwBm7/TjYUHU+ugx2FRfojvs6IhZSGBDBqNcV3/anY+fIdVwDj
a1+qEUh5647lOSOzdkoUoaYWcCPUwIY2xC1AnzJTkQmEpJxLXPraUq8WPIRpV8G7
9rhx0JWab1fd/YBpj8B/UBaLvmMLTxtgSGdGPT6V4czejm7daItXZWOW8acVEM2o
pyBfaiCjwfS3UPgAqj4mi83mQBIoXS8LhdrRFFl8KHXY3txwANSjKHgI3LGvDhIf
WYAwRp0+5iBLGpKylMVksMRbvutvX5bZQY5eYa0SX/WO/WzAVFQc7Vcn75N4+Srw
qP2Nd+uVwMPXe8nB1/yET2qPi0mUe39m1i2AOHJe7gPS4RODlS2mjp84OJBmfxdE
VGzWnDZGqO0fpn4DYdfutO6L1qMgOda9TbTtWMu6ncMxlcseMFHi3hud5Ak/WTOx
6OSLwAcuEpvdcjKAIk/k72o8drfxHFyWekcfI3b0S/oF+GFRW+mkSFzIAjv0tQVr
mFJMZTeP8ec1kjQ+lNRewsowm0zwcJIMAfOnO1VEe5nLYJEWeyCcQw75hnY1JRS/
3buDRf48LA8DjAJ1DY+47QmxUT47OHOWFjDH6u5q16uV1gy4Tlh8JV5494vG5E8a
VFPLnlicm9ekD8ZCYFFveVXNiJm7bV/9kraPxRFjRu2+7w6en9d+x38QKflMKd9x
UJiAMRkj32MtJis6lmq9pBqxGGDCv+b85vbNcU7qaRCDEeRp+KAVnajvpH//tKnR
Lu/ey0irob+vngxzbzx6K1Ejbp9fcY/dtESLm4b6n2Q3xJgBOc1YQPWa3kFKq4Ir
/aUuECuMKcf4DZAaZiKLw37e9FzHNRTMlRtH/Lp+kYn1h1ZzSP/U69nyZePu60/Q
40ubckr6d7y68qTHz9jSbCQUnrbHcurZz5CyHLhh5yNvRozVXGcVizBRzR7VyhBG
K7IORmcQ1derfGCGhRJRVdK8Axd3H8jtmRSaReZt7QbxsEAHB/yW77Jy0lfwIdcm
bpb90WWjVlXWC1sIv2qwSoGwYkaZUkstk2PF8y9rvvAkX/dJUY98Xz1gFhUlVxnV
FrJ0boczQ1/7mkKPuOnEboiptuDrsYCi2+eJ3WUz7bjAxLc134On689ZQQME6Wgi
qhqaDanjGUgV1PCZTvgZf9Q2+fMqlA5Ha74FvdXrDQuvQ3DIJ7FAbq6KDiIiEI1h
k43hEH6Dg2QpJe2XbbKqz1f9os0D//5WOZ6NG84pVqHywnJ5kwYwBeOgdIA+DH67
3u0X4WzlTYtKGX9kjkjo2332XqPamEvBm6uCOHJjWXqZYnLfZq4uGp7GyNZmoIOk
cm6gPl0KLJf8IHIts6XsyvSB0gaRMSd3Szi6D8BVINO7gEOjondjWzgFKm5bAiQT
LT9euQY0phB9ucGiGxyjdAUE/WmPm54ctUOMY3WtrVwwltXRoaL3xiBxbM8IkItn
yu1XTf1h6R3EiF0IB7I4TnstxcyOfdW6c8LJvlVeJHSd0/PnN7edEmQ3xq3sEEB1
epZBdLLVSdXlsbEw/O8vX9uRzrKpEnHB1fMydBCQtZa7n7GaUReOUmg94gbgl3W4
y9mr9BmzS+IDC7eIIsqOBdBanqV51cHm/nKZ3oJ7tt40S4Yj8+5ocYXLr66mkWGS
AbIfLcav9IFXpddCYAqq8JcPC4JXV3bpJGGhw0cMVIBo3Pg+mpVbBXQYJOia+cUJ
qHfJDgzOxi5A9uck8PnWyFCmOvXZdFHQU+WgyJZQUxc60WfvZn69n9tNlYVwRAmF
wlqB8HioclIjxg4UWh820qd3c4UkjvRgeUgkYP/i+8AUENeCSndoH5mwcQy/Pngg
W3ZIGOY3utE+uciS//dq4T/HyISKZKTYevKInbaKARdCzB9Gnxg0v10VtqjJM5WI
+54+T9jfC/qjC3H7wI4b0kVh6pqOp0AtVJjT5VOCIQQyEXE59Zcsfk7yppfadLL8
WE6a7nT9KKEEZ2drTIiqzzNeFgty44meu0STN3lBUDO7+wL9OJNAKbx9+vVPjZe7
wgMfXG+D+eWAcSfm4SXlFtsdK30unWKXrPWWOtKZLnWoFpeh/Wgv2VLE5dCQgUYa
WHkqxLDymqHkhb3ysFObalWMPA282IH7UDov1eMM8MAHH5ykmLjFsd9hkDm5YUTs
Ro1KDsPbwytWXoKVmWEgciqWyohsbJ83wfo+fjxWH1pbxz5MPsnp3RselKyzQDVc
7ZROcPXbBk/6yjvzrW7iRVUQfWbAH05CmybOX7RKoj38BUSkv3Crt8CeGottG658
3xksSrMo2KIRz4uUAAXN8zY9xSiXBjLQGqkRu3qVyHsJvyFXO44aG8HM63Qij8yg
jTtxgpyntK5Gr9MtkSdU5Sq6GnBw/HNBm4BVG+7/XiwVakMJqDmxM6QRhS0QonJB
HYfKo/cDVAFveR84ykmmrlvyMwsUeMkpMxlczxyP4hr2+ylpPFqlsqi1M19oZgKT
3jHBe9kqf13376b/tmI3e1m7YgsEMaXtHei60ES+M+NZSJ6Kg480qVEJMwvhkJiI
7wSq4n9D5ZcPHQllieEFC1HhyBAXtTqIeZOljyOw8bs/cTggPuZlwzENXtJz2iSH
gHIwTUryOv+9RAptabigYwmo19xiRu0jUkle/7B4NbRZ7I4UQRdaNUoGN8mdw0g5
LeKooHG92k2Xmts8CD7oAN0stnfH+ExIWHG4W+bwAxX3lFjJVQnLihNyllnn0NDM
+elmKxXnXX5mMOv7T2Ynuz97LfvPQz7lZmNbkN/tZARF14gRL99RdQz52wsuaum+
s4RB9LVTqTlqJ0v9WSkq7hshxg2/pR4Rq10PO434bT6bmg3Kbuo/ySOJ6dkildGG
7I9jP2FRWJrWQBLfDp633Ucks4uF18FN1xFZmw9sz30kqJXxYiltsMo+Kl2eGE82
+SXSvySP5VNv6DRIaUp4Pv18jUJnNvNjHlFePvsdq++YefvfHuV0hnfr6YWe+Ydh
ovCoCXUG0banLC6WvfyJ0WGOx7vvb/MuoiHSLDk9FfjQkpHeV2ZAclPdgSYIJN6T
NFTNbX25Q6xg9zDwlZWa2UDbNWd2ImipeKphcsv+b59APwfhX2BpRpAFAKMY/toY
bDArkmP/2XzE+m/Ju/ujsDhZUp48wiccsdF6qWN2ldc1Ev4e1MzK5naOKJWdrmQd
m0D7P2vnBC2eddZ7PIECH9SvNEVWbJ/X9gGpPP8HFk6lyrxG2LWC7OOPMqaqQC+z
riwaEx0baiJ8ix6oukWy8+nMHQ1fuzXsdXJtSZw2Cy9YaUecBAoKYpXjSzpfEKVo
00NkP9o6oH3Q5aykhoYZba12r11N7DB93hDdbznNFxpHtFUmYXOl9QD4IPwi7Y3j
n6pn8KJRS1QV9giO6dnEbleobg0jwm5hbaIShc1E331pcsQIc7YfjI2RXnmDgJ6u
l0Xznqj5XbulcfW7iF39j9pxGvjwsPnMMFd+dmdmA5rNUOuOZ1znP96AwtutYAVn
sw1S2aon5hqPt4Yp/ORzyibox9RYUnbUKcDnL1z9jV+rivt6SU931nfNcrSvvFfC
ABAphNs2KhxSfPnppGhre7UmhfNo/xLcM/00A6qWIEFkiPCsdTLUaPCcKCj9hWv9
E9t22i7Le1Fe7dqety9f0oj9uCrTglkj5Q9qPr/p2u3drbRo9ZJje2WQn6wwK87O
Tmvx453kHFFuJIK130x4Dw==
`pragma protect end_protected
