// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// megafunction wizard: %Arria V Transceiver Native PHY v12.1%
// GENERATION: XML
// native_phy_tx.v

// Generated using ACDS version 12.1 7 at 2012.02.22.15:06:00

`timescale 1 ps / 1 ps
module native_phy_tx (
		input  wire [0:0]   pll_powerdown,        //        pll_powerdown.pll_powerdown
		input  wire [0:0]   tx_analogreset,       //       tx_analogreset.tx_analogreset
		input  wire [0:0]   tx_digitalreset,      //      tx_digitalreset.tx_digitalreset
		input  wire [0:0]   tx_pll_refclk,        //        tx_pll_refclk.tx_pll_refclk
		output wire [0:0]   tx_pma_clkout,        //        tx_pma_clkout.tx_pma_clkout
		output wire [0:0]   tx_serial_data,       //       tx_serial_data.tx_serial_data
		input  wire [79:0]  tx_pma_parallel_data, // tx_pma_parallel_data.tx_pma_parallel_data
		output wire [0:0]   pll_locked,           //           pll_locked.pll_locked
		output wire [0:0]   tx_cal_busy,          //          tx_cal_busy.tx_cal_busy
		input  wire [139:0] reconfig_to_xcvr,     //     reconfig_to_xcvr.reconfig_to_xcvr
		output wire [91:0]  reconfig_from_xcvr    //   reconfig_from_xcvr.reconfig_from_xcvr
	);

	altera_xcvr_native_av #(
		.channels                           (1),
		.tx_enable                          (1),
		.rx_enable                          (0),
		.data_path_select                   ("pma_direct"),
		.bonded_mode                        ("non_bonded"),
		.data_rate                          ("9830.4 Mbps"),
		.pma_width                          (80),
		.tx_pma_clk_div                     (1),
		.pll_reconfig_enable                (0),
		.pll_data_rate                      ("9830.4 Mbps"),
		.pll_type                           ("CMU"),
		.plls                               (1),
		.pll_select                         (0),
		.pll_refclk_cnt                     (1),
		.pll_refclk_select                  ("0"),
		.pll_refclk_freq                    ("122.88 MHz"),
		.pll_feedback_path                  ("internal"),
		.cdr_reconfig_enable                (0),
		.cdr_refclk_cnt                     (1),
		.cdr_refclk_select                  (0),
		.cdr_refclk_freq                    ("125.0 MHz"),
		.rx_ppm_detect_threshold            ("1000"),
		.rx_clkslip_enable                  (0),
		.enable_std                         (0),
		.std_protocol_hint                  ("basic"),
		.std_pld_pcs_width                  (10),
		.std_pcs_pma_width                  (10),
		.std_tx_8b10b_enable                (0),
		.std_tx_8b10b_user_disp_ctrl_enable (0),
		.std_rx_8b10b_enable                (0),
		.std_rx_word_aligner_mode           ("bit_slip"),
		.std_rx_word_aligner_ctrl           ("gige"),
		.std_rx_word_aligner_sm_data_cnt    (3),
		.std_rx_word_aligner_sm_pattern_cnt (3),
		.std_rx_word_aligner_sm_err_cnt     (3),
		.std_rx_word_aligner_pattern        ("0000000000"),
		.std_tx_bitslip_enable              (0),
		.std_rx_run_length_en               (0),
		.std_rx_run_length_val              ("000000"),
		.std_rmfifo_enable                  (0),
		.std_rmfifo_pattern1                ("000000000000000000000"),
		.std_rmfifo_pattern2                ("000000000000000000000"),
		.std_coreclk_0ppm_enable            (1),
		.std_tx_pcfifo_mode                 ("low_latency"),
		.std_rx_pcfifo_mode                 ("low_latency"),
		.std_byte_order_enable              (0),
		.std_byte_order_mode                ("pld_8b"),
		.std_byte_order_pattern             ("0"),
		.std_byte_order_pad_pattern         ("0"),
		.std_tx_byte_ser_enable             (0),
		.std_tx_byte_ser_mode               ("div2"),
		.std_rx_byte_deser_enable           (0),
		.std_rx_byte_deser_mode             ("div2"),
		.std_tx_bitrev_enable               (0),
		.std_rx_bitrev_enable               (0),
		.std_tx_polinv_enable               (0),
		.std_rx_polinv_enable               (0)
	) native_phy_tx_inst (
		.pll_powerdown             (pll_powerdown),                                    //        pll_powerdown.pll_powerdown
		.tx_analogreset            (tx_analogreset),                                   //       tx_analogreset.tx_analogreset
		.tx_digitalreset           (tx_digitalreset),                                  //      tx_digitalreset.tx_digitalreset
		.tx_pll_refclk             (tx_pll_refclk),                                    //        tx_pll_refclk.tx_pll_refclk
		.tx_pma_clkout             (tx_pma_clkout),                                    //        tx_pma_clkout.tx_pma_clkout
		.tx_serial_data            (tx_serial_data),                                   //       tx_serial_data.tx_serial_data
		.tx_pma_parallel_data      (tx_pma_parallel_data),                             // tx_pma_parallel_data.tx_pma_parallel_data
		.pll_locked                (pll_locked),                                       //           pll_locked.pll_locked
		.tx_cal_busy               (tx_cal_busy),                                      //          tx_cal_busy.tx_cal_busy
		.reconfig_to_xcvr          (reconfig_to_xcvr),                                 //     reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (reconfig_from_xcvr),                               //   reconfig_from_xcvr.reconfig_from_xcvr
		.rx_analogreset            (1'b0),                                             //          (terminated)
		.rx_digitalreset           (1'b0),                                             //          (terminated)
		.rx_cdr_refclk             (1'b0),                                             //          (terminated)
		.rx_pma_clkout             (),                                                 //          (terminated)
		.rx_serial_data            (1'b0),                                             //          (terminated)
		.rx_seriallpbken           (1'b0),                                             //          (terminated)
		.rx_pma_parallel_data      (),                                                 //          (terminated)
		.rx_clkslip                (1'b0),                                             //          (terminated)
		.rx_clklow                 (),                                                 //          (terminated)
		.rx_fref                   (),                                                 //          (terminated)
		.rx_set_locktodata         (1'b0),                                             //          (terminated)
		.rx_set_locktoref          (1'b0),                                             //          (terminated)
		.rx_is_lockedtoref         (),                                                 //          (terminated)
		.rx_is_lockedtodata        (),                                                 //          (terminated)
		.tx_parallel_data          (44'b00000000000000000000000000000000000000000000), //          (terminated)
		.rx_parallel_data          (),                                                 //          (terminated)
		.tx_std_coreclkin          (1'b0),                                             //          (terminated)
		.rx_std_coreclkin          (1'b0),                                             //          (terminated)
		.tx_std_clkout             (),                                                 //          (terminated)
		.rx_std_clkout             (),                                                 //          (terminated)
		.tx_std_elecidle           (1'b0),                                             //          (terminated)
		.tx_std_pcfifo_full        (),                                                 //          (terminated)
		.tx_std_pcfifo_empty       (),                                                 //          (terminated)
		.rx_std_pcfifo_full        (),                                                 //          (terminated)
		.rx_std_pcfifo_empty       (),                                                 //          (terminated)
		.rx_std_byteorder_ena      (1'b0),                                             //          (terminated)
		.rx_std_byteorder_flag     (),                                                 //          (terminated)
		.rx_std_bitrev_ena         (1'b0),                                             //          (terminated)
		.rx_std_byterev_ena        (1'b0),                                             //          (terminated)
		.tx_std_polinv             (1'b0),                                             //          (terminated)
		.rx_std_polinv             (1'b0),                                             //          (terminated)
		.tx_std_bitslipboundarysel (5'b00000),                                         //          (terminated)
		.rx_std_bitslipboundarysel (),                                                 //          (terminated)
		.rx_std_bitslip            (1'b0),                                             //          (terminated)
		.rx_std_comma_det_ena      (1'b0),                                             //          (terminated)
		.rx_std_wa_a1a2size        (1'b0),                                             //          (terminated)
		.rx_std_rmfifo_full        (),                                                 //          (terminated)
		.rx_std_rmfifo_empty       (),                                                 //          (terminated)
		.rx_std_run_len_err        (),                                                 //          (terminated)
		.rx_std_prbs_cid_en        (1'b0),                                             //          (terminated)
		.rx_std_signaldetect       (),                                                 //          (terminated)
		.rx_cal_busy               ()                                                  //          (terminated)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2012 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_xcvr_native_av" version="12.1" >
// Retrieval info: 	<generic name="device_family" value="Arria V" />
// Retrieval info: 	<generic name="show_advanced_features" value="0" />
// Retrieval info: 	<generic name="channels" value="1" />
// Retrieval info: 	<generic name="tx_enable" value="1" />
// Retrieval info: 	<generic name="rx_enable" value="0" />
// Retrieval info: 	<generic name="data_path_select" value="pma_direct" />
// Retrieval info: 	<generic name="bonded_mode" value="non_bonded" />
// Retrieval info: 	<generic name="set_data_rate" value="9830.4" />
// Retrieval info: 	<generic name="pma_width" value="80" />
// Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
// Retrieval info: 	<generic name="pll_reconfig_enable" value="0" />
// Retrieval info: 	<generic name="plls" value="1" />
// Retrieval info: 	<generic name="pll_select" value="0" />
// Retrieval info: 	<generic name="pll_refclk_cnt" value="1" />
// Retrieval info: 	<generic name="cdr_reconfig_enable" value="0" />
// Retrieval info: 	<generic name="cdr_refclk_cnt" value="1" />
// Retrieval info: 	<generic name="cdr_refclk_select" value="0" />
// Retrieval info: 	<generic name="set_cdr_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
// Retrieval info: 	<generic name="rx_clkslip_enable" value="0" />
// Retrieval info: 	<generic name="set_rx_signaldetect_enable" value="0" />
// Retrieval info: 	<generic name="set_rx_seriallpbken_enable" value="0" />
// Retrieval info: 	<generic name="enable_std" value="0" />
// Retrieval info: 	<generic name="std_protocol_hint" value="basic" />
// Retrieval info: 	<generic name="std_pld_pcs_width" value="10" />
// Retrieval info: 	<generic name="std_pcs_pma_width" value="10" />
// Retrieval info: 	<generic name="std_tx_8b10b_enable" value="0" />
// Retrieval info: 	<generic name="std_tx_8b10b_user_disp_ctrl_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_8b10b_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="bit_slip" />
// Retrieval info: 	<generic name="std_rx_word_aligner_ctrl" value="gige" />
// Retrieval info: 	<generic name="std_rx_word_aligner_sm_data_cnt" value="3" />
// Retrieval info: 	<generic name="std_rx_word_aligner_sm_pattern_cnt" value="3" />
// Retrieval info: 	<generic name="std_rx_word_aligner_sm_err_cnt" value="3" />
// Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="0000000000" />
// Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="7" />
// Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_run_length_en" value="0" />
// Retrieval info: 	<generic name="std_rx_run_length_val" value="000000" />
// Retrieval info: 	<generic name="std_rmfifo_enable" value="0" />
// Retrieval info: 	<generic name="std_rmfifo_pattern1" value="000000000000000000000" />
// Retrieval info: 	<generic name="std_rmfifo_pattern2" value="000000000000000000000" />
// Retrieval info: 	<generic name="std_coreclk_0ppm_enable" value="1" />
// Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="low_latency" />
// Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="low_latency" />
// Retrieval info: 	<generic name="std_byte_order_enable" value="0" />
// Retrieval info: 	<generic name="std_byte_order_mode" value="pld_8b" />
// Retrieval info: 	<generic name="std_byte_order_pattern" value="0" />
// Retrieval info: 	<generic name="std_byte_order_pad_pattern" value="0" />
// Retrieval info: 	<generic name="std_tx_byte_ser_enable" value="0" />
// Retrieval info: 	<generic name="std_tx_byte_ser_mode" value="div2" />
// Retrieval info: 	<generic name="std_rx_byte_deser_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_byte_deser_mode" value="div2" />
// Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
// Retrieval info: 	<generic name="std_tx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="122.88 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : native_phy_tx.vo
// RELATED_FILES: native_phy_tx.v, altera_xcvr_functions.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_xcvr_avmm_dcd.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_native_av_functions_h.sv, altera_xcvr_native_av.sv, altera_xcvr_data_adapter_av.sv
