// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aptFjqL/pHm5Lintikox0wUJIXx0DuXZ4gFStS2Vc+2z2T+/zwUKLev8xRf/QNXC
/0KO8xKHgIilYehZalSkQhXFToxexkHNkHXa7HDa+TOAfvp6e+W4iYKQuAHqcJ0M
Ui25KLC0u+BjR4b0r0FprFPRGLIyr00Fi5loEJvEcGo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15088)
8fwvXbM2YZ/485fXp8kTY8WTxmQBCSrDMIT1cQYOKv2hxeN4oYHFzePoFkZc2tBQ
HU/PL3vkAF/ZdheKkVT6pXuswnVfcbGv4Tx69e7v9uoGjwLzNmqFJoTSD4SLaXFH
MtarligTqtu7G14lSYOzc1Aq+9eRAYRUgDqn7BiKBJsJ9gp3pFy1gV0ZDi3CzP3t
jQqZiOzGhSAZGoVjesayj07EOnniGB5zsa7vNPqckolc9LabiVM9Ykl6e1+GC0Di
8zKC3jxAu3S6pYWcOd/IUozfZmfS9nCFrpwUIOPmoawywOm2BrD0C/wBx7NJTpHI
mPJ4vl6oCr1+U6mgYqngNvWp2zbeMmD90APIJzN9ukBgbfBc1vZ5NeKUzNAyf11i
Yx7uwCVyF0zJbVx10uq0dt4wKPRvlgGNgyx2ukrxNKJBR2cnU2yNy924A1rvN3fm
gZunmkWDUPmbITLTkuTpo0kbZC9ZgASG/PWakTm12IbT99yUIsslCST4V7JfSg7+
CFPTKjDph+I3DmIm93FnDfnYEauWFoKWP6gzpvrDDztJQcnURE3mGU4ncQ0Qdzzg
dHk6IdPXs5FqudsyWwrfaYWEMFjRG2zeJ199Iz24ICrS5jXgh5ho+acpvL+k6h0n
Hifh3iJ7d9kQm5JQ7y7EbSHQdJan55h/kpgJdiiRUVyGCh/WvJCMMsn8ygj8slre
WDlHvYu7FO9P/yb1t+EoJuAmMloMnl5P/yhwmf/4oxNHwFNVSCG7gsTsT1fZFcC/
3FNcMLZwRTm79kircucCcH/AZWT7AjhC1iQLNWA7eoAuiluamE+uSBwjQY3Mw9Yv
S8gur1Ehpr3m/rvbX3P0oaeo2YlQrMffpMN+SKXN7BAZdb5dcDkqB6AAIklg89wV
4e9yoeTB2tOSXaxVv9fH6e9IsqbemnW21cBlvZ5fP9CNRl2UDoHi3+St0//IUBaE
wTXBmBhkHa1lJc1cHaHtLehmf0hqYiwmVnaqScr7/D0xYYEF6gX0jYpOqIcjmtWh
w2gKfhYPCe8GfeYTCHV7N4+ug0WgOxQOgPngbNIRdFR+2RTjk8GmzCkco/GDpywk
WhEHQ14yweJovE4DvRlF0oidHKklOFhZWznGPRNG19W7kIr5dRuzS8jg/q1zLTnz
0ZWz0dBGqMFSrpyPIEViqPlnjMz4gKf6rOwX+pAUghZ/X1jS1BibRKkxcgq9MSO7
hIM5BG8of8Po4brEG+ZHWcLN2Tk9RJoy/xtWERPNwlC8sZVptKzwJq4dvjQ8cE2/
8Rm5JscO9yQZ4W+jme2Cc1v0ONpeemg5l2DQfg9no9bjDmwTGNCYZ6imV1q97I2C
bwqZbgCtuoMfxr167n7DbIyayomNjAJPrhIunAkoQZnrVNQu2JKjo0R6LZ0JaKlc
tUv6t4jGAv9TkWwlhb+P7OF4QJ42DGF/6Yp+b+8t9TfDSi8zaol8hQr4yofci7qP
y9S4nMn20F+U0FjWma5y2dM0X1aALvWHzQ9JOPB+kwUnX+K2lSm3avZCJrJ6zr90
rQtoSvrq/jBIUqxcukWbdkYvE40IhuPSRNMk4QrRfKyR1p9rIBAcBCFR3AP+Hla7
jfN1otpNBuKohz1UC6md2o/GV7KQ4ZDz2eQLd7ULtiFYUcc7pvjNyfAnfzgQRpVj
Mk8Ha8OorNr5foJT69GBxdlgt7YicHkq0HxmxkCiziclTVwspXmYTPo3vp0Mq3zK
WeHCfxImZ75xXr8HeKvTLiUXIXdYYtcdN9speyg7PovndB/uooz3nx405itMCTYL
Xk2EmVCJi9UvDk2dNtbJ6MHch6xTEEEgLQKZd8jBd+JtL82dnv9xS53047rDqtuH
6O8N0mGvrCsbnWMB7j4vAt4hSpAzZsIM++jxYUq2xpjwbH9JIpXk7Lv2uuGPDfMX
lbPusWZZA5xJVsPdWHUOJBXclc1iu7jiiysPunoCwDWkhCCuAJfeqObT7kOHsAa7
6IeQ6zKWasWvRwcw05e5EYlodu55UfCaVjJLoKxnhQmwmIjt2jVumzkniQe7dcSI
Wi7whfWG3KwtXlbVXY99qKKlAgraOgDN6QLhCpqURYhDYqsMTm9z/z3BDl2kesNd
NiqTF4y2+9svKqXfjLlje/PG3KWRbFBNZekavv6hYwmc0oKVMkz3DyrBYzjSvUUw
eHQvUa35CjpuB+ZHTzp6psn+f3zAARYSFWEJoaCgVqUKIRTT2SO0P70wnjTsHzl+
HVFYLMjfcxEnL2rMQJegxzQ3o1ZvxPNbUJ8CFXTuXAFTQCJBm9V03uE2DQqmTl5a
WkDdW5N44v1BmY6VMwFc+PuKr9VE9PxbOZz+P9F+mt88/cON+THCttlUqaCN8H9M
A+m+sUI3WV3AGcaTZcDW54yFEfE49E6vEui2Y/un0HJS3jmIXLElLF5Qli56J6Jb
bEtatiYARNzHtgaXALQVTT9NCuIzVsriVDrucHIUtrr/J74AkOrkC+1llj0BkCVg
iK6E67+IqJHoAzwnSuO73TNhFntaVsyLEyVzeBzzm4g7WC1jHzD/BGyiGkLaolts
cbk0VJgtECnt/8HCZtXW21r47Uy8SWC0RoGXRUvBTH55db/p5C/IthSQ26MDXK4Q
CrtIKtLGuYMp4CtWJgddOrK3DZMrvEjBDo0MhQf7nISvwcJdiEZxwZcnUbZsJ4jh
GEDXKqawY8MJqYJW/ylZZoBYAdNP3YECDQdQ+Jx3lJVitLYxQrvjzLCg49tvqBo6
ijgq216jt0g8ymZDPFWii42zk+EYZMZ+D8QBxhWdMAIDYIVJhzdrHJUX/xhIO0rV
LtRCnDJvxXhZpwo5OU4OA/BIzcDadOE/6P2/69kzkU7cP3u+oIRWei0pV06GVFWk
R9tzO+AwEIr4lWHSZFYLJtRGsp4kmKm8sVqUSbv/16tXR2XtIehLJ4UEivz94naE
SQXYJ2iQN3itKB2fCieqIUNGMaDNjRz6J/t17fwT+jBE9ZvqofRUipDBwZ4e9Smj
lFpdUs+0dm1JPCTXkpGxvFVT7WHQcSCQt6mlIYnK1DtO3r5zTjtOFb5ZkSZ2k9bD
Xu8sExM8sDjQWeyTynVvPsfF9PgoG0C7wrdxqfSW9W5O4VrB8MTjYJiwqT0ptKql
JpS1GXUb3rvbHWYPMdzClkRF5hwXrHAg0wA1CsZwcq8y+7NP0rw8IgBa7pT9KcnY
HP1RYfoJ4B8wQqLSJvrcxewOuO/+GyAvLvoxdQo7q7NCNgxrOm+IQpFmxgtyjhIY
aJ6YOYi6a+ZE7fkH/XeRaoXzNbvoI6/d6kR9Ec8cPFb/LF+pDpuptb5ZMgirT/Qu
BvElCUGXA07WxKA4VDmkn8+rOJzKloMw/mPPqkV+1nQ7AXoCJkXQxl5lwb6TuiBj
UxHd7LOt8imObhk5qFAGtyoBP5LjRSSvbIQniPYXye5SVx467uAy3S2bPwfXTzIF
tpCQZDwYM3RuU3GUuVZYWevs7lwYl1+3BQ/5ZtWe/sIGo/LFx9lBMYvHlC/kqrrU
zORlYTR4wVIWqN3lha3tz3Yi5xrgPKJfaku13pREyzC30hv24ROrZ+fotklV6ZQm
aVOnDnP6KAEK2ZUqq7YrlbvmUFQ3DTeIZ5KQg4K0RgojkvybowY4VwoFfc9h9VMA
NIrR05HgxGdMsqhP22OMzZRSHhngvbe+DB7W9qgqeRKcYRoOLGR8d2zTV4XwrXSF
Nj4Qvo8UaP457TJmFOCCQOXte63/iL0++JJYnIrpfV7Z1nsWkK5dW44Hdbi2wbm5
6Y1HR+7PGny0H8akzof11X+6f+FyYKQMB0Q4+4kvhuDmrFbZXcpjQPfONfMh2Mq0
5CMrEkcPnCVx1FkE9FxUq4vYDaWajbCGdNnATWqzie0iG/jEThwi+R5APptipOQ5
8i2Yy/y2S4LghyG4AlQ8MnisipQEcuPB022SLN/Nmp6yRVbNLHZjrKdusRCMq+AD
Mw8dpZXcFS1g5eJcVC6ArWOgClm3XYmA5k/ULqf35aHYU5jBJgiYH29i9HN7RSXz
hWIf/YAqoIpBR8nGECy1TKyAESWq5h8hmdv/0+GuYkwvTbBpj0GaqB6Ceu93iqU/
BVSca62+xTlOv/jlSjW3MqKpScQuVBpYmhmbWOwCqHQ2hsG9wV0c7HS493QIaHtO
GWNSBII0DOOIwk4ZR/QTqyYtPyo+pvLLecLlEGziWY+4OS6pyLl5pFOSfr2cwMvz
GWb07LB9olyfaUknwBC/dtElDa9wpzubW6Zjr0jN2jlMbEx9HjGnCpx4LNLrhw+P
uUSwTrt2jURuQY9i8WvmYwS2iGqrx4Ao374w5txWQlj17Mxi3bORJs+Vz7JjqXVg
uv3vOBkdFOouoz0+B/qBS8ZK2Mi0aalfhLQlBSoWnIr/v2xzE8dzdLS1OKxJaiDo
aCcXEG1VH4HqFgMcZbCRzf2wEqri0ywQVc738SclofsgN0C9TMJib4Ivg6X/gtly
4UxrleSDYivGVn12lqKUtiGjFZ8bGUwypZcZfrzF1tksKc08KhVREYRgcyk7zGR6
HNUbuBZwJrW6Xv6Z96Tx5Jl0hTj7rQnROb3gAKF1RotqAUtKm0B7yBIv0zdC0FFJ
rWfPlkEUdP7MmyrnCZ3sgyJDbuqKBYzkfPr/m53AgOD3IyGOJdw6Ax3m40NzIBe+
MscFrE6Iz/QfiVKIuYSiAJyTF4JkmKn/t4U87Jw1I5gu53BTZT+dH4JjfFlB+PgK
muCa02qBchKk2/P40ZyWe6rNzHEvfhjBwIDg9r+F4nqIKAL/2g7EPWI0QTebJL+N
M9TLzbMCNqxG9ofmTze7qxeIEUszIJ30fFEDS8Vc721CY2y++EjXJhgRHmavxx/D
395CUzNrXfg0njvJJDO4DCmTCmTVcTplAykDikTe3M7EUXJ5ln6wvI4qhcK6hjOR
OyddJ48aMagtqeZ9NCQN4EHliD5uTSlBQSaAagrW+TVMB3OzQKPP/YbxqrqxiSqH
Q3fG02Qb5yTczan3Z/Ved83Q1i3aSPkFj2JAMS14ESH4S+xq7eMvEhcufov58MWU
1qjdYhU7Q2NAMAwZJfxTCwTbL4fKsKMesJAmsHjZ3VonKRQWNVJ9a6j6vDM3APw/
OLm0Iz0db3jINMiGZDxtsznu0pD8+wU8FCGNNA49w9xPQnQsLLWOFUgRMJPaise1
uHRWo3lb2XQcRcGBP/AoMz7vczar5oikacV8xwJb0RS7xXrroKsxkZwRcW2NHERe
QZ6B83EL82icvyohEXQomOAF2wQQqrYKbs+Dzk5ySA1mxV8v9YKd3CXy3gd8i5jT
bNg8xdJeVkV8xp0gInamgH+myXpNonc6R6Ycc8pBgDOX/i8g4a6Ve2kPmz/TFOqk
qioWurm2nL3lPmcldhbQ2cyd7WCYQWYZVp1/vTi7T9baPyQpeXypNF72BFFHHJC7
lzpeJ6oqlDuaQzhhW7xfn1QtwCucoGGaTUnbGOjEUSzyTa5ri5q1JxPaWHWn7Hpr
RFgqhI8iM+jQUedcj2pq7FR7aZEUwhf81fus+KRyVFFYGr0LCzsxFVH6JROH7Pkh
UufA5y1yFGUkM5w+WNkkDT92eXFWcPelbomEjFB1RyR3eCSg8f02ML8meD2rzJ0K
SGxRw/xYYWYmfmScIgTuajjAd485I/mIJvPKZVDbkKDKEPGZ2f4393boXn/hK+ox
dawnpBdFmoT61C98OQPs9Dud53cXvEMMCL2k6LpZji1nyQxqJ95b3qtlPJTSOKYp
dgJivmJhLZvwaPa4MmSG1AOAPj+sSK2g55coSeSBpMS8NUfEfF+OEwUMvFRSFmpe
WH2GEseUkRLJHu8Xl03t8312xmv2yOezDDHGpeNHfaSeWTloIVLd0KXaFZjJ7BM+
71Oigf4riRK9s5e49yrANvOM2RJhRZlyahRzUoltwG/s5volUZSCagI1L6f2JC5L
s7+ygLijBs78/xJ05egoiTnbMm539iGnvY4tN2gIrZTE/FcmQPQS1pUidSQk6n5r
CGIlyF9y8SVQHQ2pNNeJ1bYpIpxMRUg03A61XIAPpnT0UseVt55bTQHZisqlKo/f
vByesTA6kJI3/dzQqrg+zcpbvaLuo170jrmQX/wKxcZdWxN+lscoT8HFB+aVwFAV
KYBSvOMV9eSX+3lZJHTU3+A7rB9oVJmAsO+PxRVuZFgkFOo8U+Q8Q7N+s25R6zgV
YVBOnWcpSU6zifPKJJJv7t8lfhW5qEmSEtc6brvV2MTBxHbYhn06olXsR4iDXVth
cbEvFDXTjMPQdrhUIa4Merlfm/rS01gp+oI9TMRAKNFtMGS9hA8udCW8hnEGYTx2
QxgKXHo44tDikh0uIf7I/RjQuUN1pTl+M0arS+qzWQSdbaUcS6eBUq36N5qTq9u4
tZj2RJwl/7Hnlbc7qyeYob2clynouYd5v6ag9tmybSnRTxTOFikbKqZiN4Z+V703
LxjJnMQOJIHsp+OS6BQMyuix49AnF/mosoAuoEzCS6qXRJMhZXNkGZitULtKboF1
KBaMMD6u08ObbBvL7/FHq96q2eyBs734nC5eX3YTHS5Ilh+oFrJgLqhobdCxAEQ2
fKU8QZ6ai41NEVRdNmASzaRDg4oXwYocWLZ7Lm/C2XVW087ua8NBU/nAZQFAK45x
n9gF4n1VOEaYUyYHnJluCzvSXS3NEMVhp+NhXIDOY5Wbxnml8DNyWayRG750QX3/
Gb40ZCTr0t5cJakMQ7hAzvVDEM6iyPanEZFlvXxwjssTwfdAI6DTrK1aOE9D041x
DCboCBPz1bkkOdQbboZZM3zYi5SUEmxpbZjpsodbBdoyXm6gE+BYpyIw1fDC9U6N
T31pp08LjjKUEnTxLUb3ZC/yYzvHIqebF8lKxlDVnEZbbOooyr5H632l0L7itWGI
4OYbUXs/uQUlxjVzFsgXRnLHK3SEH7wxeYO1HkWytriCqVMmEg7lo+LXniMEIHWB
90qDe/CjfWSgsqyF+I2a5tunFOs6CwtHVXPXiRRI1S5LCpcopsKkEjhxA9B94bl0
vzaWLPB56k92jVGjjT+BDOaWiSg8i+Wn4qcNwSDEZTCIPoq5o4ODrggXjKmbvg01
2BffHSHeUz1cdaT+wnMXSgWXdfCWd+FSBksxFEQywug2XYfZ8bkKGgTCmehQhk1j
jEVZOaf5VB2oDJHlT4l4rEPGGjskp3JXbwTLrTQhWc9HZk5mG8IFl9cwuo2h+CHc
qQjJtORzvy8B9CFqJPKr7cZhOxlGZZExYtiy8OKYPWVXoR1dfqa4pmLuB+oImPxt
i6kfdSED0c91GorDo4P53bWouNdcf/wjpki9T+SFvaFCl5z4pbN4aMjNCFAiGRML
lA89bQ/5qk4mRzYZ2FSKCWxSsFcK2C1yR5dGJTBMozzRpies/IwEWO0svHh+xqE2
tq3k2LDOyRfuP78WKtLPGN6Bv0Jc8iOjDboJZDH6a18C7+RPQUM40TR1hUGj4kZj
x0qgADM8fuq7tFJnVNzVdmVc0D3BGFQLHhVv5NO4AIMj2lWlVwTUmK4NhWMLYBNf
GekWGAQxObGcTxGTamLhnKL2gVwcp2UggKms+cIvasmk54dAVGtByQcHlodDfLxN
AhX2O6fdolndlblXUVFFWko0cJH3t8+lwcxWLsBGGThrTEGa4B7BiUazmYzXfQJI
1ftpcqOiMfArj7u+YId85u6aLilFzumaEsN+zg3XLvGbJHYAzVbg+jCWHMBFkOHB
gBYWueJG2LDTqAK3ntHQJkVlgMDYksN6AogLT+E2TF9Kart4khLVx27LOtkxiW4Y
y5qN67l4U8bjvEazTRP4Rdy0xB/PqAn/FvkmoIm+9UPDCcvlfrQ2JjFb+xjlvRxm
YNIaDH09pulITBlh6TS2T4FzSRcKsdyB1Fye8TJAkreJfgvl8gdz14TRyEucr/ch
VLam09VTUfXGnB8EG2RzE2wrBjlIs2uOmkoyjkxwdwr1lWLqlaj+cOn56P9IrAFy
1pmxokOTkoX3lOhLc2PsXPcwf1jb6YT5gk4D05MYMKdHX7vZDfC1U6kKo2pMl18E
netog+JeDKSuhVAQvJ06H8aROQRdDEIa5IkS+36W1j0JMcEfojX0rnSvEkt7uImO
ST7Nxz3naiUmuNRMoY/LRNBt1qVzm77N2TFp9LtSzCm7puVgDNlGMvixsDTOl/hX
3NETrAck0ERKNmODRnpoXvE62u1bK4sp5PQoXxlkkVQME5mwDLlVjfPoaxarxtve
ezHuj5DDwSmFBGZuTBCZskICRX5R8kHeeeZwZZ56TKeJXQXb9552VCM4IyoPAZsZ
1jRN1IiNJjU5P43Ibonigzdr6pgOyGDoANmlVRsdwU9MIN9MHhqd8ygPKB6t2QZT
TY8JP7SOha1eoamqdDbu5FnBNaWT3hNXp0YosBa4St67nnYS4vrfHBwye5FNA99q
OWoQ5ZDbsMof91ItXilpBlJ1pcXvuH6EJ0etdkmSK5plH7xHhOYoor4lbAgfgBfw
RhdLHCd9C9Ryfu+98v/aSiFV3yUyL5TuSnAJA7XmC9lHPGNT0lTOG9ZN4gtN5HsA
LoPnPhsRyO6Stb+0EuPOuyaO8rNjcy+yFNhBvGwctYO2cst+TGi7FxalOeOo+zbF
9VOCs9+fd+3bUK827f7DxL7zOhAYbQst+VuGA+ravd6LtbWmYQ7V2MQZRZ7AiiZq
lGcrnvZ9tkDFjhOtNqEVnY8F0l8Kr+1Y7X01cmqBOnGopGA2+gTziZt9JBjBWaMR
BwDQvCNGym/x6j3Mk8qIw0hyQAScG7zsmqeWLWuHdJYi9HUs7rAjVeLwZTvekibs
q6jo590/4YCLloUrkZUW5a0jbyd/kTMh0dcK4Qe5sAjFAVds3Mp+mE5cSPRvGtdi
+2S+IyLGpaBJrE0tLcSwFCs+13do79lI5A57oXwY0hWE/Gr2rTGIxJCsj0rJwXe3
ADqvx3bmBM8rsagzCmfzdTDbMF6g+VYtXmH+2qbXoEo700qhCafXKGHmBU943orO
br+HDmIs5AKjCemlUUZU9YpPeyMk9UxSIdH9RHKYXKN1f1VbpUykBZB6QIoo5Mnv
EWSOvXfU6UvpT+Sk/rBsZIU9R2yvLv/V6MGJ9BvD9wGTxebGhB1zzElpHJTAmHll
1bRUyXGznhOt/uFXY2ofzGviKaIS4HZ1W6giKrGRmmy0tT2Y+U3Hfc9JDD85Vcxt
lruA2d6JPV3qUBlACCtolb4XE7Do85+ZJlveHxZA+UecpOZXH7+tkfgCdj5pEvSC
4JZufCpu+2Pfy5lLz5xd1vAe8rO92jc9oSWzAYboEmK86Vp6NaxFZkMulnpyGpVX
ZevkiQ0PhoRjwz4NGChU0p/fMPoZTAhikZ9SFtk6GGXHpDmKLcfhhZYK+Yqld1gs
ed9JO+7/LEnPvQVUp0y7wB8gWvkKq8RNtATTaFNCAQCZ8zjRMP9AC2coVsIMO2kJ
ucOhDqQ2MWOI8a3jE2vrctXds1RVGLq/cP8BbJTdaMEW5ZE8j5Gzq4hNJnMboXKz
NeHJNvdUAJNraGmamz15lCMpT9rUeqd23vcjcyIuJvxYp1B4FzoDqbdBoKIPQU/n
j7U20QHvUJumgpBrTb5RmPCwBKBFCl4RxKU33gEqet9rrA9vW2ZNAF2WZdCjjBD5
169CmcTEMdZxXzsLS9EHW5NxgiqwVzQke5Gwpzy/LsKfdalU88aIA9liZDgo6Bmt
qKmh3+4XaS8RN14HqnYkFwTx5mMsxeBajTKx35RutBADyEEomXKi6uOPLeUI3XWY
+ZQo+EObgFUdVGOZonZ8Ca/TmDwcCdLIC8VY1BdwWpGjJxAX2Ap+2cUCHz5q25k0
1+RTd5hLjEXKkfYmaYQTFDDTUEsmAIj9Neq181xWBVeUnooDjyFO+xXVsupnCfqI
Vn4mmZ7a5LGRppD1/THInl/CezqEsp1fSHENr66Fn8ja4mUaVErfaZ9E9k4l1Jcs
p88PR24BGycfWC+lRWZNZ2qiV6OoMHhIRA/ezi1kkkgTIEL4DtWXvEn09L1bUida
Idw0EJ/D6jTHEa3ckKwdwR038PYjCyPHevuRxAd5dULoS5Bg9oNWbnznpKJ97id/
uRL7KKgoafQ8Fd/+1tFmz1uinMPEX16vUAWSknmtf/fYYqz+og8wgjmkiI5sCrC8
K+C9cnhbgHWPHyqE4Pl1SW67kGzetlUe2dq4lrGTCQ6KCSCZAu9X1+Pcgz7iw7lg
2LiGWUByBFJo8/kQMfB9EW42nOi2+nPCdn7rf9HBKmGZqrPsZsv3DntZZfVgUfFt
tL82CY8YWCKiKFAcAQfgS7ajrtRTQPiVNVpV8on2DckEaEvadbmkHzNqWx0zVnFQ
dA/DJIN98FsssdCgnteFcPZ5MdDYFUURkPVB9K2TNoVnDtdB/2+MQz8E18rjOzC1
bZH7zZoMKZZweaCqVjCK8Q37FXreD93WssmJcGx7zy3E371qSmlhOkQFvH9ntoyv
zjg9SrZBHR/B7aaFbGTk/BPq8M+Yk2nAayQ9TNiyAxGUO1l62qZKLzonlpFsA/Vn
Au7K27JKbGegk08ioZAhSObAm/zPPmJ8w46C51HGpGiyWYevppPfyHu3qu2qqAeB
vm6mCSgQrcZJaju/PR0yFyubClNiitzUVlcym027lD5yu5RYsDNNNhNgm8pkM26M
RCUDhjzB3EKHdFgCwAgSVSmaMsfPj+i2rS38l/8G+MFaLhDXwz7oa/iebnkTWh6m
QqJMxE7lkp2rClQcr4+dNQBfxa909rzxF4eNopXozd3CJTuwgAbKvuHGdbVvnipt
vM/CBtdwkV9XieGioCW5fELXHH+OqPAzLU3cQZBgPXKRgF8W1uBhmnrON/DhiTTB
GOCsgMy92FeBTnlgbtqxnUaFNRb/Lu2/DPr9J/Hx3fdKEo9IAhtQQdFc/G1Awjjg
26meEeZXlR599H0NvDXsEcRDnZBBUfRJbAzSe8hh4DYlCW56QAV2vZcjzM+lvLLW
CFZElBT1U9KgJergS44t3rbWPjFwW2JksVpknCTXdqQUpa/t7nHfFalAu43BZ+01
60kj+90ph/s208rcQDC3VBx7Bwblwgpb2Eae4Q33D0MEIrBDpnVipjfhZPttGmrZ
gUfUB93UFZ1L2PaBoUWFpkRaJ1DQjVU+t6//s5GQotziffMnQEUWPZ/znITDYGfF
wId/dHCh0J9wKg8xXNmT5OrchboWD2Fs3d6Slwz5Tb4cwpW8xDflEJS9m6AwIpgu
KCxubYEFwUyPkzFDiYdWjuxVf7nh1pTEciuacIhvf5aUChb4noX+d6FF5C1fRQWO
a7HSTk3gTgJ3CFat0AhQc9Ua9jQyWR0zKZHwCTWENXcHAbUph+z0LkSEg6u8VpIU
eXr7T4jH5LAuczelpsyC5QoiBkGP8kHD+rpl5oNLGP9heW6V8VODhi7EKLNN60y4
6sI8isYUki0jCerWZ181hzDkrKksDfvK+KuyTzsjgiZvmJ8o1+O4kd3LVpQ9rN8X
EBzZ9a8szHIC6ZYFY4aRoYOruzUW694c2QoA0xNUspU1PwS1Fj1J0eDkGT+zIIBv
wxLqN2+C4lBajWzVJoc5GMcfnF1GPwjKpUz9X7gpIdmX4pXlCU8Nem+yK4iFRwAe
ZvZUoweUQ2ECWZ6Br99DxVMUu1Yorja1gqh+0Agoqd7tqVrm1/6JWJNoxcMHnaB8
Ktb1wbfzfmbYSRunewaNbVIUOLag0e2QJTGdvzy+sfAAjrYedmbyPyFNKxEsdngY
8gPEL/sX8NrlJy2ohmLU7vW8aqaNDko5aZZUFBEc03AVZgYuYzYG6OpQf8+27Ekj
LuW2X8pw5funTMOE1gild8b4c7vBkXQkRPMnoDcKfRkX5xrtyVuzry0EYnzuq9S2
qfrpMLQwZghK3VrE3dpiqdGcuu70gEXnESS3Ken8B9E30dtaTQyrr902AFCwyjII
AOMKsMPUAO4dNa/7pKpFOI2v+OQmzvRYLu76mHnJmpi5ygXdQ/GxYrOjTPAafuwj
t7UbZZQRkKDBEGqLqdGKLQHxy2n9L5wAgEuhmZrPgDfDGLc+xBXryuijFbayhbZ+
NIZAntOq2AIwveWdrwZY15cktJCSR6+lokNyKUn5mpfRCKQ+cehD9l6WtYPyUFP0
itdgJIZv+lmMvNFecXMMegFqEQb72tDaxj+H+L+1+nYYGTdTEkRUWETTwCJqxunm
GmS2+/q+QRyjAYzWvydlQHprYqPX3Sx4YTEQBUiB+mohcjisVZ+UZoXVtHAO8U+9
gUCk/vVwUZJnY1a1qqgCWJcNUb+Mtdw4/mC2QYk+jDKsVMK6rROxtWg3tAz2C2ns
1WPFp+G3/GJMcpAnjVlAAOolc5MZ9orsDHnp2jBCds7x19psJbU7BiR0CQkeDWMl
+wF5rYOHFvJHK4zY+K7z7rW27ZOEVzeikzGzwOtVnQgt313vcIUf1D5Yz44+BF3W
g0gPj8X4gS1BM/nTiOu7U/DhvjFMUfuFVD+UbjbYQnk3nvJAn1JAgQNKFsNVmo+X
Vr4uoJC5Vy9cU/qmCVaVGdD4JNfsxq3hl5mFKua/4tsY7K4njkhQiO5Nc7X2UcX+
MOoVGa4MNcxuXCJYrjIKR0XRzRRafsvITH43TUhM4J/OTXcJY4ZHWZ4w+2As/+0r
u/b8q7papOklWmVtCkbORLnWH4R5CxRprTazlBFLCefpeJEBNIXsjGMb4R2pXtWO
x0bDt91g4d2LCn3dBWx0VVchRzKO+43+b7Rfu38n/KoSLiq8ZI2B0wzau73Aehq6
3d4vlBUZELscLY2la5JBXha6N2fV2DyJehO38KGyH8Qe1wju1GiKvaCXEKtoWyaY
nbFTcFMiA5vaLjCSxDLpYILrnAZ6JBvN+sm42ydLNaTzqk3Nrq24MD9U5eLP/9lF
+hjBmZAh14HSPTmXsJu/uJu+hnhbK8Ut+7MpMBK2dQY/6KcFLNdiLKaWSH/K9asE
KS0BbOJ2cqXC47GeGcnlZhH7N/WeOdTYc0uy0gERiTU8DvhC/YPW46Ocj3w9osK4
lwRrdijVAgcwsy8kVhDm2w2247A0KMsin6yyZ9Bcczai7RQOB5xUayLN6aXenzl1
yfLovHNcitkA4ePgKCvn8d9zYTSdKQDYGBu9Ag+RZ5t5RkYxh7ZWwoWRF58PzITh
jcdL1daMsaJ6pa7MSRk9Y0txaj37bE0DOEHcczul5LU1qXI6E9fWpwEyv6NjjmuX
GlKRs6Qhi5ww/1eIb//JwyAJCGKLUfVjT9PPIb+GQDB5aLrzqP1zelVAdLChPQBM
ur6F34STx8vkU7Q/EY2UUyAQ4gd/zhgls46YbKWcJsu8N+99VTwGCaKhILZ2WyUw
sST/oXNWNLGpsLlvEpd2vh9kdgsOyAmOEhdCJmqSO/TQrRbcvu1+OhH7gecYmIdb
aD5bIjkU7TAurr/v9R6vK3WCzsNGTwbJkwWjWrgWXCoxU0yYayyHSRMKTIkjWfE1
qTfbYFILR0TAoey9JrkBZJF821Jlgj0XrTn74OHs6EZRmWFMzXWJydyjT0cWU5Uv
Ho+NqqNOiCQub9Z5wdWUQne4ljMasxdiei5ZOWJa/XTxYQ+iGemdLUWD89rbIStZ
2/es1w8yYVHIddTfa1pUxQPqSAwkzEo3i0Bx2LAZ9GkNnkUucZBc+pUmhD2QXTw4
7ncgHVSzUzsiM/DvKGhVOq/8GAMxkt6ioUVmg40MVWpnCRYil+8fsUz4Eh6NUPhz
xVnYGOMZmIoJqg/S+TLpTdixo44nffXtFjjfqoqWqoWJFO+3GmSwQQOpMmpdiNxL
+S2QMhIgm6P9oc0+H38UPG1oFMWHl1A0xrCxOJbHzPhAuOY5hKAW1w3lpJVkyBfT
kinsK1notEv4pFvsCh14qj9XYWFtsNslE+jZdzDs0z/rYGLO159IV3VB3V58guHZ
qQ3Idtpw2Ufvk8bCLP5qNIZ1EM2Z6ToxfSVBgkGgEhgupou+t0B9vp5ZSAlo4Kmg
j/juUIaYC1CQKnF/x1CxQkKvtT6cWx2M+ekAqWJRajIuD9/TC2o58SUV9MKcxtH0
3ArJg50FWkN0p3yeDTtNO6jnuoIe5/QXnzAFS/qzNAayCNE6U3xxt85RxLLKWTGR
WVASFOwm3kLKi4kynxR0JYQjclCYht8YZhTfTfYA5lCJuIEJyTvvN1j6USENJ8mY
lF9oOhilVGg46sL5Lq6jPonw/CvNBm8CtPi8aLXZRwHH7sC3LMltnXxBOtAMYpH5
pdezu4PCZwXFYNPcePc3bXRSwm4SO4hnVP4Tinc6+hmSNfFrXM020n4xX7TWnFm9
8iOfQJO7vGUE3C8uXD98hKuC7kNeUJdA1dYmv64kpPhmcHQbFu6VH8KOoLMlkLRC
OxGuuudmIqwsVHy/79k8U5mpJN1iWXaOUlS6yz/mWGigQos6p310AEoSX4YHz+AO
rm8ImjPSOmk8OYeCI1XQJOAyVsxL5axH0Lo7Kd7hE4kyaks2XVxU1+dfJvEfN6Un
jdGlWx2rPo1vXbi5Ec0T+T0fpuObt5Ani80XhdxT0ZJCc2qtYEQUg7KwrxrgK7+5
GeNe7iO5Y5rvz9t+ApbRqjWD8RY673jnt/pmeuct6NzQPCpoqFCJpeTWshfFYyUR
8kyCj0bCisAP/3I7QwckkRVac24Qmk/j0Rsy6dk9CWA1lqv9PgZU7TCo4YTbxHtU
1y5Qhg1rRqvwnJx4MGZgRkSTcdPydlbpobM1sdFEkMwDPvBIRibyrraiklftWL8Q
5Rbdx8JUAW7AjBwXJ0Kk25p2ItqVv4VKbxq+1vH6f041EZg4YMHHXlbRnehCb4vF
9e35GKLQiT6wWQA1JegONq2wqPu/kBD/NJwkPjF04caX8jlMzuqM3naav70XJy2T
zg/kuX5bnB08kNRroDDWqLKbw0M1WpAQkbZ/hwjk/TKMS4qT6HnL7jUa/txNbmFT
bxDYeAcGURzWcUV3gPuAIpCGL+PfVouTMnFu/Grarlavus5SF5TdVbuw5Z4ybJqf
pqSf/hzIdQsfbZ4BclUV/UEuRbk3UkJgq6lou9XYLVyy++3wI/wE83SJOyVCybtG
lyp7bl+ZufrN/veK0c8ghc6zmAmt9Y8J6nYEBqaflGPtyZ+NJIKeFU+fnFkk7UH3
Bl2VUGtjTEsGw+5G8+hSjvAVKLrl+XUE036DFlR8TQM4GbpOD83YV7sRiiIKS4Ys
eFsUn3sEdVsVB5EmkgPUCQPJMuVpT3Utx+RewLznIlIDcNGwOf7F2r59Ua9XEgqW
qazf5UYJYDB+/8cTk31HNzXVHK+zCctkV1vYdynilgJT0F3awNR/kvPlBwgevAR/
hLMQFDkT5wdDlr7oS/lCAnubodHyuNYha80bI9re90bGYGLuhwfQlYrQR+8GjEZa
DvIoREnFM1HfygNWTX2pQqFk3nQA0jvmOAntA5Aey+HLB4v/MsODmuNtWdhygAJA
p4CzSOL5yN2e9e1lSuO0Yane1xnnwjmoOvXW3EemuHJ0on0uiOuIFNLjWcOaxPeZ
KSdvNYWYRtOnLAoPsQHrBjuxM3R34xJ/qRdsyVh16YL3APgpYrpzJlA+oKBjZLg8
VJiJunY/kFxQCVIOW9Qd2vBNrE5hCF1DfAO3qzaDMSiY73WLUv+Z4UpdbigiAmHK
F7LduPeNjZGZ7P+TFuertW887w4prp9GHB2K3GaTHBI0mMlGGWqQHqqbplnCVRTP
e7GYZIAkBtIk8Cz4xWGXGRDyUaypxVu6wo4Kyxeuy2DeQdhGpHrKZDmt6mCQSkkW
ZZOCopYdnTySFpPY7z0GHrY0KsTz6xT0kbJiM7Yu69tVF0+LNcHMFdO8rim3ttGd
a14pp5o5jnERSK7bA03lu+zRDkI+n6dRKgt66lgtjAFQ9XEitGlxA4V5L9bsUuEA
eOHXuuBQoR7cyNU4Gtevg8AgNPoY/xfQtWyu0DjAO5zWXMzE0Gpi3/Cgck7KMkhY
QlAuwctZM6pAFHxkbj4/+ZPVErIp3RoCEJ6z3qb41UFSAT9r5efY61ZNVXDKlnNZ
3fEDUyZtEe327JT6tGlzzTHxZ6Zw8nD8lrp3p0vUWrgbSn00w5qN8IS8QK03yWlI
N5sZ+a/a3IcihhTliVJG7MCIV4dgS7O9gUf6VcODvY5OPNlDi4bsKARJFo5KALpf
9QqvuMRVsGt2G1mJ/O8dHVyW1AaYGF2DgFmVT+o5dsPtB7LlI9w9mLvK0j2k/0dB
xqSzp/ekFqipEpb/oKyoz3Vjfmt24mIwi3qinWplH/UmtI5IHG3YDog89+b5SEir
WGiO6eK3erhAsU8oLZlp/J49pNUQmwRZ8s8tmbpNizTUzMu8uW7z4/wG977E/0xo
JqQETjOtZk783Zg3WYGZF7tKH7eBkuCImWNRlpB09LgYtj5i6fZ1k/z3Jkoq7W54
j5T2abyQzWKgH1vNVV2XtAhV1nCP4AJ0xz8T/Kd7y4oSU/Z8pwglfeDuBjQ/ELuh
p5QJNueBb+WXuNcQHyxI2AlDxlfr3mf7rmbzHw1KF5ND76jCaAA+UF+ss2SKocOb
M+3K6X/PHl4BqZX6V+ZataXIF89FEEXnTiwEvTeny4fVv3HQrt/L+7IQhDPZpT7O
BfMyuspUYZaszeTI7Md3sKpf4dOXDLPYsSrw0M6eRjCOj5oRrviosgm5r63nRmUL
gr9VvZkt3qVCuNaSYDT/iMXos3sUxSzXyKdtRje9h9vhRlZrB/gQ24NwPyW583Iz
hxhal3OW0grVchRwiRb/AyECkykessR2IREWuXnXIOHxz2JLxqpQU0GGyWUkOdlX
R3Rv71+DbPzYbXSD2COwjbD0LzeoLV7XZCRHzdAOb39mCJ7fEWLIa2Lkp/EkRABn
MtDPIHWmQXoBQlXG1ybRayo4Q/FCLQO1Fr44qQyt0xKf45OCRQsQfpoZI/mqD9K/
oHS8qb/EW2A2c2MxxbCZIPQA9MuSBeJ389nUnK3aejmO9BQWb8aKHvNPBQhYZUF7
cL5VpFSsYoVCqldSrhtGwi9gMI2lX08Kuu0EVJ7DMnmNAput1+dLNZxFhLRZNYyt
fjnXZegjdlUllPLb/u0KbS4bu2tTvHnhUYsuU4CPYyaJr9YMdflYzpYw14s+oc4S
YN2/wBkKv9TyYhlUu5daAPoQ9qOTiN/59puU40brpAKcuHSE+o7+DCeuXHj/WL7/
nVCOB7o0Sgw8R3q+Gm79QfxIcZnJNlsgxz0aNCMCe2e2VAzSGgBIZxj6xEFsJ3Ve
bQNbFUUSMXGjFYEji4aksQSgPXZlYZ9uDtivSIcU+41+qu4ublPibSORhCMeJcyE
vuIPKCzKTD1j4rZ8fnH+G8EfG1l/bul40pweZLctPrLJFy8caM54TVWpAwKr0+6M
U5ckJ5C89yxW4r1GG9ljz5peq7KY5hKlFRUjFAh+3d5v1keNAIXvCsk0M2l7lYTr
TJ4GANWK4COKSwRRJzwAeLexiFRzILi3lPus9H3062HE4IbrzOsWR+YGgm4Zj1fP
vFAq5eZ/VzQYt979UEvkEybd4B3cjG5tZ0wOo3EA0DRX3+W+0fvldnPiLw6400+V
8gPSJjrWeikFGwyc3a54/jNGfMd6O1rtMt4iAPmqZl/nqkZwlxucVWIE//Rfk8mC
tlo5JtJyx2sq7E4ykp5jToA5ochadPMu/uSjmbcHppB/R/AYBNmPvATzyJuK0YuE
LFVjNkhC4hnn2vFiDXBctHYonmbIPO5S8fjXg8xa0iJPJz15zzyje4tNugsbhCYp
+zqYgafS3rqMiAMpTwsLA/Xqc8KXonGoiKquWE5FjpYeUHGVyBD1U21ksfxnn7Ld
hgRSJhvoWYUjc36HxVmhSfhBTo37pzT2KeqVlX3VPYAjkiVcySzzHxadtRXudfF0
dEQPRzi8rTs2Oj47TI51ZLQ43jZQO0sizitpM2pb7UOsMu73luhoT+Yd7kZKiwS+
VKkpvLibmoTqyr+Yq1oly1KtTrEIOQmH15+g8QLHQdPT3XDTo8pXzpf3upXhpzDp
SKR4Pi9K5G8SpvFDyUbmCr1mvccpRZXQssyQV0mO/hohMbQuqRyhL2Op+RuaxqRC
DDAz/DNNuo1oGBhPh3MBJhpwRZy9k8uxp1HJcf6Y55ggOkPxlvzSXiEd7hRoofh8
LLVwIgOEgY4ibP38wjGTE30hR0dihXxd38fYHDPrOFRUd+Pt5LRX4DIJpDA1ppcM
ash+MYsQK+KW0HwUdBOXIX4yeQx05TAERMpzlD1VX5qSdLohsPP7vAlQpuCJvYYh
n2DmUj1iY7EkuJqiD7E2dbS4azR0+L7IZVTHfACHrxs9UnVLFXTW2TF2lS8iTqoN
zu6DqCBEw2RJvECFoETv15+YjBJVOrV9i3GgFYZ6BF0RKIts/a9pNX79TCdhYFp4
VYDIwgibugfaTyKjvwI3DVrd1v6draw4hKxBOJjoSuDKyfj3I5Rl3s+qBRL6GsE4
bFArSiqUyBVakp5c1hGaj6ki7vSl23k0DzeWdpXhfUq1BiL5xJM0CARlOdljaPPZ
GRsQkuSwGpby5uWslB/eph/Ukl304ikqGtjBMRjnfpGQEWhwNkHhbG3BDrTDPqYx
3cj6bdaMaO/x/ioD2ckzSlX7WGXXdCZeZrxPkseSf19jRUDu//mc2CO/mZQ8xF96
0FUqZphMSCT5KtGw4g+wgbg8uzfB2M0Eg8sO9cXo/Y2dV/NRnWxl05puThi+Vf1Y
PCkt7w6s778lqKy2ag/VOt2s2XmJbh26C9GcbzQnwCfpXK6dYTbX1+AFbqLtr/Sq
cVxKF3cBsY1kFNe1VNDKwv2l5Fu7mOctNWGLn2SYbkRX5HqgETZLrr96JsDywpbx
65/30/FS+nlxCPfm78jmQKH/qfHxieqIeP3mM5BIzgq/m+Ujcutc4QGPkWsZEd4C
CWU7DNqBvc536fZA6TKfaR6hmtP2jgUgRlaDRzhUOJgtGrOEXId18kG2Vsg8UyHL
6A9cgqSdql4EuW3uvevCa1IdnkAcaiZ6EBUBhwHrgZ/TQ6w3Dr7YhT0X5ml86IW0
YLN9W3N5rIngr9vMkPit8uuCjTeT+ZLStIw61zWxee2JrVS396zvhmRtBFMrnWrv
j0RZHHLGfRbbcM0bmf0mQtpU61gXz4hQSDdW0I1HNwpyeZVnDvKoPZMzCJTagIXP
wn5/fMaHrvmybZrGnhybGZRGK79Pjjq/vza3W4Rt7mwq06hIuwLJ0VKKADleT6GG
vfEX3m4WduWdRLYf4zSFOelNfnnAEnbqLZOSP00ga3Ys/AnG/E38Xt4e/Ssoc1X3
ulXBuwnziRKmIKzqWH+Hcq/DdjFlBsKBoqYO6DCQ5z6JI7wgGGSUezSUO5ijkqeR
/aBlUPOnjtT7vA6QVjamCBtMe7dR/ODfoR8XREE9kEIUe9PEXww+OYUfxnCr0hkz
Dv7Vb639TdaIk1dLAl8aJq6tacTq90567lQsRt6b3TwQWQA3UypSRnTftFvQlwhn
VXu+Rw3zhc77IwGGFEDLX3uIulghvlBuV00AI3wbxikKVWW93p+eo9JhVTe2C0PN
if6TcAgajrXvEAJ+YB4EerP2I9hohk0E0OOJKkXd/kBGrZbScl9dN8IwmTqbIDsT
Pf0q7pwiIgF5l1SW/L8zKUL2aH9NSTQyTzfxiTbLHbSPeDTHH/87FkbIeRz2y5V3
vKiX/dqI9A3pr5400OX7/tSifJxbijnhCtyFYi8sSSSGzy1e07rOJhmerKiXWaCa
v2JGIvH9yA1soLysC8oTG73UUzeRnbpJgumAs+tfNnQbjy4m72xvwkQPEIvYE2YA
RFdTyHjoRenRrFkAvPu+QMFImoXJwFJmJf8ffMioHwMbOYIEN495kjTN+8DdKXVy
bK7qLKyQpPZK38v9bk40JtGtSr7N1ayakz8ba9hlQ/HsI8GupJySAeOYJYRgeCNS
ij0FWW+9aOzMgDTMxRDDqySNua86Gymoozt1Ix/t8234ixT8CCE9By9ocdsUYnT5
9eVYseLjVFztyGA85hPboCn7SgxRlti1xWWe50O+/i4/Gjawwn1eqpwpGJsNJKj7
dm/rifLzijjcBS5PLv+gvg==
`pragma protect end_protected
