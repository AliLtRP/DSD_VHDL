// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
EeZP5UYBfZHCjtgPh/nVe2weDTStZ9vtamDE3kSR6789sPPtiZZy7RNiwB8KH61HTimwtE2QEPJh
Iq/EEm+g99SbVcGQp9fkXfHvcbVV2Xu9ftupYS0OGSKHDQ3D23aLpcSSgwGCtE7kTa/akt7in/Nw
k+inOMiq2kz3fkbOt1q2GeOZ/INlW+vfP0MFQgYyS11fP4+5T2+ksUife63BjK26Oe2UOsG5ACAp
lt+5IKsZuNT3qWc3PyZModkt/K68uwwRauH4PnkijIPq+a+tdQq6piSZoJfmYHhkF/2W+5O55fj6
QHnItY45cjxrfX2C+/TlULBjipFmpjfaIm35VA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Q7UBvCwtKHu1fHAvkHXVRZibL/Gt0+HVvjuIVbqNpZBVuFcyaVaMa6D8YyTU/YTmbsj21vyVGbIG
K8jyhr5FVKO0S8nrjxDZSG2dg+OdWk2R2clfAnelyfIWqneJ+quCHNNuA925wZr6ae+7ahbO9D1V
DwkXjOQUY0c2OrwEDg3ZwI6+fp84WLqEFioyjsnqEtpSVT0OAn4DNO5c2VwYQyu3NyvXBPpB4BtE
1U9IVmvkJlnbEj1ZHccOiL66Ga7mJXivC8NuelZkQhRztncTL6UQ085AhpBhyaBxyLk2zkjxUEXk
1cJO8fMKS1fxb8Aq8iQ+hipFLn28moU4rz/2JeBitesFUkshrlr2LuAnTtUbYZY0ZhcTlbc45vyb
IHVQL3cn6PBQYlzE4JIe27qdXS4EKwEGu4uVVGlFXyu1hsc6A8DkZhMzjC4v4r1cNiEdh7LAP1ZL
7dc7T6NSrrOLl6FkA8vTQOPvKRmOKAdSvahqNPVVc6hILm5dPT2GBrzE1xc/vTy0ZiBIYu2Q0OWD
sy5R8209BhxKcJQIbFg4cR8FQUXkwW9v6FKZnhrqyY1CGSf8R2cMkVc/vTlzcYWAJl9OuYDjkQ2W
hSuiGghAczY7phWxQyZjMm2E4O9YUfElEKUKDE8lpTp+q8yze7cGYbV0uDBfzY5yX+g7AIPIs5H5
9D1LRmwGOxOTr51U2co9L39BOBSe333oHtpVBVVIuM6Y0Vmt9WNYNqW++HGcb2QGfk3ZYefMy/nw
xL2NZqJSkeBzlssvg6LnOaiSeNCFQ0flaWaSmyYITj34z8u+m738rf55gKoXQyyyCG6twV3BzUjw
fTA5d81wXCFKWgALHR33BDxa+kOC9Sn1us3oT4yQjfQ7gStOkXODu/seGdH17/xVt877O+iNLgyP
O+1KWmjh1+f6mpeh3xkbmaD0pv1Vgtai77V1fox+dehWHNtjJ0LL4V2801QDu0JGoo6Siq6EcU4w
E2P1OaLzfmFT9dZMR/OOKhOZh3Wm1daKZWGsxMd13X2m3SkvzC1qxZp5+0gu0aCvjsUDuyES5TIX
unQuXbt5OFMD493JVx5Tv2r2q8HKfNaGUMp2F49IMawHZbFMHZt32cYwKd0nyNVZSXCURuj2C1IY
GISv/O0CkAQ80aIiXszs+nZzaeWROZPZHW/Aak39AAA1+bdinwuLhyvTAVOKcDWdY6AhHuX7JiMH
W5D71cU4d+F29rbIWNI16lv4Y6dbk6AvdCZxRtSEl7QknE+yugLbfShPnIj+t8kgKKMeMxd8Frmm
PCUJK15mhMDmgSGIBvHOxidt+u4h+RvjsZmINrgh/gqLLJSHQ5AGJM5jdHCqdzsYw+C2/xnGDE1Y
LrOQ/ROYNymjjQKGkeiras1Dqw7pXB5VoxxzXhk7/M097dhQqmB4mBuCZaBxfpCo6noo7XTMLf+n
uTPRrcjbInsAhhrhdnNYkvc86Yjhkkm8I24SgKlSVfP0zhSv31W3CJhAnFNlr0l8aj3e5KXZm9R5
eNuUeJFRm2ZBhgrf1YuPlhjZnOeY8S2FoVKQ+kjskBerfNcdhyt0xUJHUTLLBOykxH6OQTbjn6f+
5yQFjI1PP5IOIioKTxhITILLml8gp4E7qjY6gtf40JRWdvDzTTij9IdSW9+vLWUywgHqSi5inUM3
5OzPOLz/p9EBQXeJRndlnSXm3RubGShTtTQtWYujpV6Sd5ntrTYC56L0dNG6HAze2fhdRzGbBvvs
0RXgE6qU3+4nB2wfSJ8Hpxkvztah1qk7StwKMqvAheQRuLEqxAczClr3YqrxRDIxM3Jkp8HFZ67P
qFQc8yauEJajV6O7u7B/xhTiiGIb/tkUKEl7G3h6JFXwyH3em97cwoMoBKQ1p1Ih1GlnYwY0zL4P
+uBWmpJwTHhA13yzOlmE0zwZx88c6Q3H/L0bsW/aTqnpAHJ/mfAFJA45yo+VYnc7ItwRuYeDuN5t
fOFDAXzrmLhWmfTyekoiwdGo6Fh+vxefmR4WHleKUml13uKJU7lkBN7xCkJok0iCzdaRmJZjy+/M
aL/P9CUyDPXQnXVFw8c3VO90JAvoMlB2o0k1knRNXpx0NwiS7rlIS8VXpTkvhPdFgNHiaOJSGmoo
LlpFxPXyWHU8/uy2QHAv6r4kl20MZ2iWH7ZQD9ybISvVaq6Yi8CIJ0DTQkPst0WQ4TwvMQhcIuZt
HU8f0xdEgsVqRl85qMib6gVYjw+0ulyFEMbhZVn1T763IBb+lD8f8yckqERIgEyg9yzMd4IEoKQC
p6uq96rwxmx8vAWqUwwJaHQthM4BSdk20Frct28ZDof55bnzfqMYdt0h29zB6cI1n+DTZEpiLhja
XFFMEehqAVWqb38Zr7EahwUELLcsDKXua5W2MEpf/1HTOKU3hsrM+28ja4iJSMSGW4bpJd0j121k
LTdaS2yXdbFNZmrfyoyqRe1vypxc76Pkydq4GFcxeD1ajZ5HfYykk4eU0pb1Qr6c8//axbAU1vYB
twS96XxThExYnCWukk/igKw6zBrlwhZ2MR4Eo9PlmE8v10142OQ4k7l4kb17CEx4HMWk/+pxgbQ8
oznJTsb5bFJvTd26xZIvezdAr5ubrkaoEB2C88YFRkAbLXrdS4DuWDPSbQT7+u8/25fgini9SQhG
YAp7gA+qQlcvTnBuh5lIVsl6UYmqiwImTSU3dP0dJKsu9P029zmBwEZM+LWrRM5QCpeJ3SwbiGQF
fu5l/hgm9jeZFLBl7P3VIeo6p7wZLy3zqrzK4wBwLv8wejl6g9jSzGnOKKAJF31a7LxezK9C55di
HfQsMgzIq744FUSQrTKs1lgC6prKuo81eN5VGoq522l8YdKI64WN5kY3TU+Y3dqowJ1yUJhIz27X
6Gem3VNnA89zhK5r2mDnx4EMqNTVA4dc3myoJJJSI4FlwmrRVu2MQN9ZDvKMRWAd0wGTW91ag03P
1/J+aQ1avzqwlhl96yBtJBcZgBUd29e/1GjaA971cCXtJyEon1i3TPAkqQ88uw+j3G4GKMO5vBSr
I2/YAqGMWEJOg3gDNEvDZO8X1SQHmoUanN/HAC8Ns5WeEV9l4oYz3zpTm1Ie+jE3ueOj1hjzU3RB
6t4vZr3KYSCdIt03fUWKjjuMJA1oaEoUw2fA1wX5MPTAWNqLknBEw7GrmLuhzxlNy0rXdEN4Xj7l
PYmURI4tPE3Eoc+MES4U/qkH0mhQLMY1866hJMISbOa1HW/2H71trWQBpZRqlxsBs3Wxsolv+ygR
ibkTqYFbRLpWOvlfxz9Wwy58+fyKetStgtkr7oWEO4Ix+uQ6AIZAzDgGgVAT4sx1I8ypJtfm8ran
oeTnzAb3ygVs+xAXG5B2JlM+JlWNqdXw9kULs3Ghv/Fmu6xfqS5Zq6yvd74YULg2UX+apf9erHGF
appkOCSMyLl5g5mJKda5xrPYMxKWyxzvWyxE02+1mtPMLnnXQdq/KkW5ujn9dPCLJe4ueBKcPl41
kZ4xr2dTzmn5JpgHnDrhBtzofnXsT+aeu7A4mo6WP/k2kvJtWxbsEGc6+2WuvFl3SSGahMMiE+AE
1gG6pA2Lc7y/MwVWKuMJIJKFcIz34eaFgTF37wEkS51RPwPiA9LrVm7byuGap+XVVjFOr4z9ExNS
7euGD1bpZrOF6O+g66lySr0PKzwkx5pqngOJbJPH0+4GRr7g0YxQHKHOe9AI7sv6ceUATvf1B0kG
W28/hadQ817RWLXVRWbS8aNRm8cLr0iBq58Afesx+jTCISWREfpj++iL0WHUZLWlLrxD0GCOZFoc
9SIJjvoCEK1kmbDaw1vai7ZJeZzESC4QLxDy8C/VwYbBGIBki7pMricmj3bonJTCuwszGU7G935l
1CDjREKjWcB8PvImZt+CF+DuPgiCtiIJtXseYA9ybvITtJC4WObSgd4YGffADz1rh0DDftoO2p9Y
7tgu7+X0GusWzB4oiSlGOGAEIlWGnKA8tsgFWkK4RSzaCY26m4ZoP8dD1Kr3kmUfVBA7C1ER5VO2
ooj8sU3DgR6e/xePdTI9qAM5wOapiIHnb6y+1a0Rqlaxo3Z/FsjjGKUK/cJDOkc5y20Cbu491aHw
oHr0zNy4KJAmxNE3c/JExSWmOAzXXQhY4pDlRtnC5ZdBcvW1qfQ4ZzHZcYuMFTnNofnv06YSkM+P
g0XyhtCHPKBA4OxjeP0mLowQzNoSnv4JqprlOn7yvBJarntyvJqYku1E6+XldVVs6ocperFecHwa
7Z/ASYVh1SU8tRJBL3RdU/2279REbK9JpUrSjJC/xGI17vXYGHllP80UQTyhIrHlXFmvnKiItiCx
1dYJvzhcRRAWxkI94TD/BT15ePhZt8DZhzxYPKy/08pvB6kGsi3hg0aO+bCphVBTm9ZwZNeBd934
znmJDnA7bkenW8+Sur6/pz0jfCEum5QgO7s9eGrCSEi2fWvdNH90BqBW6ukWs3HynhZu9i172MEd
puujQUtzdwY6tWqYNiPmgZEBdtuiFLZx4q3HOBq7OepXHyR2vlvv27W4+Wex8tUeNhMb/IuCVA2w
rbDYfHq3MVyjhWqeo3Hmqv0zF4lnloVU83z/QfGydfAefxIYrhCmJZKI5n2mAuEIJC6sXe+mcxP1
ABk7pZFJz9te6JjU1ghajrFxKTpCCGIn7p/q+QaskRi5SZU764azFMziIyIwuJ608+b/HsVIMKOE
HTx7ID4HNVOwpzwIxZzQqaKko9xh+J/5h8OZ2mEOrfTrRkNQEX63Yai0qW3z6eVQkhJreXr+t3E/
hZiYdhU/sx4bzu5frVRwFqSO3gqpC7zfqh0zmb/sKzcyN3hgzKFsCoNEa4zX/n1Kz8is70O9ztMK
lCJVDTFu5E53ODvLuoBGeNPWf69utzNwtT/CQZbMRPJoauUxQ/e7U9ax0gEOYPkdCsH+Q+HaXm9F
c9TmUjcb+ER6Hporl/Sc0iwXlyPkhiBbLcDQfZWbwQlMGD/z1BaWUxMIgyrv+Z9RJmiM0K+MdkfY
Mwexj50AGr/DQgu21uitKYzgAGBKdfW+twwaPvLpw5w+ZHBzwVaQWQ1ZNDQg5EqFhHs1DPqZP+ub
s/Fk9rn2AgpcmHntOfwxiyxNrBTmnGhSnMRk4zi+wOIr0TA18uGFodzmdJDOiFJRpGuSRvgPwrF3
0k1EbfDmhoZvWV4Le+R2odhBpcrKBuTi8hNCj5djAlCe1EsQltojPlZVDMuE8k+PHFzn4UkeU1gm
oxdNtc++bRwARykIyqA3VwpsGivNbMh9MDuFkrxrmfr/rEwwvouydqnMLUrb68pAxxWcdxZZtn9g
HCJjsEGyun4R4/mqajrIpa6oGIyvnd1Sk9r95liMjamhXJvbtw0Yi0O1MNqEEmevlHZTwzAW2AFy
YP1cN5+fz9ku8xyW7AXYlK4vvKBP9HWmY50Vd6EaE2qaESfkSsUJSS0WBCUyGBFwoMzGlTzmu5kG
BP7tcecZLPuXE1FRSxKMDQsrXWSDQLrA4aBGYFITXFvagatw14a8VMPtw461NE22FOOL/t8/QTFe
5RI+MHTJWUhGrgAD5aHjnMkYd5gFH2kEY/Zkv03hBifTev+2ewYIjTn196ONT271YQLF9gBkhJz9
rd7aCQD5zDQKVo5F029EfcGQ0anDXHMptUbkmUJ3DSXYI0ExhkU18n/D/wcG4+8Zy3cmOlAEHiPZ
XCASnRtUyAP1im9CMC+QFU5KuIPijRJD0SRPxeKf+wN2lYeGy4rF7te6Z/DaBypk6EJA4MQNQICK
BCA1TfleBR4UClYX2OEpB3mQfJlNjch2W2og2brq03YwSEOQ71b0J8OIOWzetzeMatGBldy5B7Le
v7T96RWRhusfR9ti04B1ylz/bznWeJrO7+IXeuQqmLBgoWu9sU/rdaO9w2c/lbr0q9tkvg2tqaWj
8RbhD+wApqWY375w0n883xLw/f8TH4cCkZ3fNSClR+jPIyu//PBymKbGiSWydEZ6igwW31Z5Mqm/
Vgz0VFWGxAkIdLom2Ja/4vEcKzdJxjXcjR9ntKD0qltURLBMIEm7cWwIPchI8lIprx2yNfez46o0
XZ0QqehcBjwMKhNPwNIBF3WlUf3kLet9QU/w+SWKGCOqg3kMzGNx8LCsX8kXzWvasmEz83WnqBRc
hOn8lIogJaUp8T4by5TSn2AuQXKbaLv3YqIrsMNxNcwV9kpusgF6paixdUtMTe7gDNNdxpRXS0kS
jMl9Rew00aA9qLpzXq0geqXvqxtDWOsQzIf+d0kNzS7afPBJhXeTvJfiidqjEhjO5rPjR+wy4Cb/
KXTXBdrfF8aCeMuaCu3xF/yYdtrh6BQcHjFLz8sn/cY9SYejcEDzliETErbKIL20UtRsvshGZ010
ucvoa11GyVBRNWqToLIKZ1IBNdL+/iLrg3id+/4OZZhIo8HxIIEKkEpwuuMxpVOGSi4VeEUfPKdH
Y4N99F2sPUrKLqdYugTnfvZd/QKqjpfJrwuZzT+bzCuJPiWi+bGw6aUEgzZcgldove3r/JRNrUUr
/KQMCv1352FFsxBRK1Ok/uhNSMdkFJnavQBj5VRnrYTWmON7vRbDDScUpXD3rkFN/58bh0eSkT8N
3i7DDfIJJwobZtf4rEIJ5nLYMfsLgF09EeruK86Zdk/JUWgm39xZuIcEcA5nvC2I3spAC/wEgrAA
lVBTkU08pkrzOG8y7mAzXSo0XRQ0iB99NRch5kw/B/YuABvriynXLhrNcXxr5q/duj5OD0qazaFH
Lm3kzNB8Mugs8cJab5+s/CbsO9A1ZUH7PHRgU3DSM9joICgkQRrZgbH6/D4RzsBvg26atBfW2m1V
yZVDLQ2nZFh8W7vKGhSJRcP3mAVP6FT3bAZuPWtQm9CNF3nId9jLo3vOTVgZSzBpV+K3XewzVSWY
4UecYZ48yBwbxv18yKDyaUvVjzdT84mYwHHpnTAQw4RagqwgqxXtn0WRtl5y3/cpvGCeV9dUCLe3
+QvEQYNcAkQloXCL5u87gmWQOIMwPGYyZRpTqU7DYJJFxG09txnokGkcgh5eDkYqUeiXK01nqma4
t+P9A01VMDIuZp1qwSgvcF1u/fzSftVFFLeJUXeVqWuE/0kGChNGpYn1On1CTBOhZAM/2nvK8PBZ
WSUBA4tjk3lb+JIIJKCUOnqSeAnxSYZ2BdF8lhimlqccGDwC5tesdSYwkQeMBlVOIIuu9WNBxMn5
5kdBmywf2QuFjvipjKnd8S2Y5D3A2fYXFiUgw8G2OoOKmM2hQfwaVyRDW1EDoGP21hGTb33WVnZx
BJse26xkbKDrXYLp2p9CDiYj2AzZS5P/n19b3LDDZ6i3SV91dzZBJwaNDTwQxhqvTu/c19q54rjH
z/BPvhBiL6ZK+cj63S88/3+2ui++CSNyaoIuQ8+mK7VCoMmT7jhNGIvoTztcWHyQV0lkEIULIk4d
JfwYpHUzCZg8ID2xULVF1qQLgdm1T9aD1KKHGcyOsFZYMO+ck8hf/0RZNDPsZCVJRelvadXd+g/7
l38nzcb/Pg/R3I7dDhM8OBErSwVS/YWOsoQOeIfGcOHr4465fQ8pNfRPHm76DueKnHstKqUSCeNk
8hhnwep7j1ds0NC0yvGA1xMfLfwoxrxkgfiBcX20ka6d1qqv658lq4iTgm8SSkQmPf9h6Gxy9fpk
MiF5/T6wAWWjBzNbN5ldXGAoys3+kvlLE5WrK+ZQKFu+ySCyD5XCFSRHYDLHsZn59QLfI26853ap
pLioz0066gcsQ/+/5IbJaFkybHjSn2q+XD9A7NSyvNyCPkjf6I4rjQNmQvHiNMxJGSSJPMs1AtnH
S7/P8r7SitXud47arcxe5uh5jD7zMmXmilaqqwysMcm0PBOMrtI4AHc1rUSx+XEazSBueMYDEwZS
6hfAZm9uMIsOgBmxQ55oDeY+XR+EeQgEoqQGPuTF7H5CORw8jSdKD4kjXlq54oHoNIIUi/JXtgCi
cuSooFBwqLQQrK3DQfEdNevi+x3tnJlluIdUqKpWCu6xAlkernTgWvcTOdN6OWtGjOjN6SI229QF
HWrM+wonAUExCGjbQTNQrWqyKalPgf94LBtW2w7ULHoR/5zMdOlQlCWJUXHNeHg3A97LwLb2uTFg
T8EJ7zJf3jgUTqQh9szz/NEz9nsiclmuxC+fOCFyFBgX7LNYU1TnIeR/8+C8Lo8MdjTMnOfl1t6R
o46HDaxYOCm2Nx0oWp55Ukw5X3i9js4/xIG4l9okzmNRVfUYHFe10EFGTGxX3uiZF7emNoizJGyq
LDZm5ipSitfEhXJf2QCgDZgy17PfXLLgNOZ0zNs/zYVn9nSIPBefU5R7bgwdekj48S0lTYXZLn97
i53dpdIiv7Zlk6+gv50RRRAKN0PMWquIct1Ul3+8s3WcxmSyL66wByrsfryCOIaWJAejOW2BP7qX
+3ntGOdu8cfi8NIAxoGH8JGFVTLiiGCC+zyZd20NxqBVCzjAQ2aErd0m3hULm0Pf5pX2aIUJFqkg
eXqnMXRQU5vqdUvYyOhxzyw0U472R7g51SzunBPk0mSP1gji10eExqvHcTl/+mQ64uPQRxvWHqX1
LPZGa6iqUNXH96zhkQrhSXXpPfM9UGmpqJCaHu5ZbJ3/pmtnQGS08fMpPTbin7/QT8Saj0CHmvyU
oHzkiIRx0/Vbcu56rRQZkljIfEsdG9yGLnWgKocfSDezpnvVNG6IgSYo6Go3lMZ9EXhfqYW5t5mC
RvN4ZGNEU0TwmvQKiqSoMe06CzraRsJd241n/DvaX76ydzKCsB2EFi0G8Inq/57TiC6DhZ9jsqEA
hcAcC9mR1LId2Wfti+yj0CIrtJeebEB1w0U6JWsP/4IgXYy3oALZQ/rEPOpsEZAopjzB83JWTz31
CGcMh7BnYVF0u6vw5jh0hGxZNdA+PTVsSCG1LbayGMVjhCzlbTY6FhXyDYX5NFy9T1OdIU7KbC5p
XpFuPhy4wa8X51q4MOvNMwkGvN6dBg87Mtc5zajRydcSqnPoQq7erKKDOXIUwaTABbXj4yEu5dgr
R8bJLlJmM05t/69dMPdjmDtB6E6LkedwE9G99E1szsGL889de7yh0u8fSKckSQldxS/xtRwDHfhP
H1Qgk1PYa1j9Rp9qPBbbAnUXseaky9dx78fhO22naA245fvEzlABWJ6zbGPORFtUPAFheGxWxGqm
QR9jeZrkrZD4wmGvOLo/D4Sr3oUhC919xIMC2nn9lUtEny6sU6sDleZOUxwzp5AkjPJeC2fC0xrc
bCTXmUToGY6gdD4YqS2qrzkV1GEc19W7mcfgy/29RbQzzqI3kpUxqCUIQ/H7d8gD+BXtURU5ebbb
Jw0ikr7W9btTamaumKm+mEuBJw1Hll6Ggkf0DdTs4EQ20XB9dogmldD8hwRbLlh5Q+ouQlUCGNLc
puLaQB2Kdy6cOef95JNVypbTUL6GxLUKWyrJDATb3fwjCW651dD3nSG59XSB+pEdYtmdaUNnh+6I
Yxa5ywJkDGC+s/ocR8ulR/uMfO6MhVAL9viDeog8lY1t7ZORBZlQM7IImdqj8r3TBQ4mEBp1Lq9T
UGuQcD3bimlTSmpfZmY66yX10Wa+PTLR3t2n9OguAJfNyCHqQcXNBkvkOM/Sa5dcZXGQBE9jpg6y
Cw+uNpVj+keox41Ahq19jcGTRGNyOnsVyrEn9nsMnqZ2reOBpXpLoN2uMdYuy6ogZU1tmXrmkxtJ
6u8fXY04rHrxPbfQjjojsQNRtTw8bEx5ws24U5QWv7DhxKr+5v6J7J6Jkeb9AJ59l3r0JsRy10dT
UpNHUuxglMONKEqWGPU+NcUjdUWCi62kgkDzjBSVQY4X3DQyBfl8CU3W8bv64eoqxyKficmwrLzv
eQUUINBza/2UahBCNV6PY7oo89edg57jjXX+x+ypeRRkrmGBUgSh/DDhP7NGYLDKgmDfOAijnvNB
rEYgaMuRCqMxQktVplSY5ESwz5gAx+JE8nJHQQaqYlprUU4G5yR7ZVgXuYgJg3/TdAADvO+yzNnh
TfMwDgFytRcUDFahFQcqqTZuQQn75PUxsT4ACroCE7ljfqycijF0h2hW80KEJMjnLMNx4Am8dpQG
wNeipeI8w+2wBwkycw19K9DEsgEW4fid2sy0EW2roQJ31SgBwmjVbuZM3pt0sGbB1OuHm6yH6cLt
K0hG0U0BU8J6IfWBvyjJO/OjdbxKjTrj8KV1twXafPNbbE/Cg/yubFg7VQzrQUeAC0CN+s9mTSRt
T+Au6qIl4931X9aea3XX9zyETKUu9iFKPhD/2NJvX8Drh2n5V12vRBZ5EIJQyWyQ3knohbHrk+Yt
nQHhU6J4k9B7pyZXOFO92T5McOACkc4rtTVJidRksenETTMrg4h50E2nM43GS2b2Y5R1CQQbPXqj
1LtDgQyDovueIdPbEysKsSJPb9i9c40appp2HtX4O1g+YIbkDb2nVWFWioPggyeimcAOX2a10N3V
lrfqBxpPFfTANulka8px3uIlv1+5qx9orPzZrKEpivfibmm9Kx8ClqefkZwtuY2UayCtbXuFgXNh
rRSLGeaSEkXD0ZAvqIiQKAG34zwReH3XVnnKtLu0dNN+vaIEqVNomKLxmBKqfoWOSRlVMQp5eNyu
g2nKCVTuOlsEA5LjbsB25Ne/DEu+5Xv5xc3eqfkZ5WVNS4UjoN6eNlYx3qo3xdCL8Y7J/E7AwJ/D
XmIQMnRJmGPwdoWrgJayONWXU7wmUb1giip1tpJ1q7hCx6Ra+3ueG5NPaZaAERyDg6n9GfcFQcaa
u4hmNgS++Znw7qopSiL3Th/NriYFx8pWxxlthnud1v5f/2Res8u+3L2lYiK75ww05VGF2mN+5wVk
hV5NoyKDYvi/Y8yCwRmfWeBhwqUazXfb4HD1qtKKC0gyE00p/Dmi1K3gy5Y7VxQvZ3TvwpQeP66c
5VaJNee7G/837Afhnhbad/42t0ywu1vDH7zNa01iOugNd50X+1UbyLr/lVCTY345jUAk5rve+yRt
P/xveC4StQlUPOVY/j4UDPPtWlYQhYDisQ/X0YZQRkS9+IIfFKwHXKcLCfTWxbVwAydxXzgOD5L7
ZF2q8GS4bo87HUVSCt0TmivRqmt0ONeWI5FQmkWCTIKGhKYRdlDN7sTdC2+TxpFNXfJbR+GBLfvH
bvQyr+PocszbCc/W9gVfgbuIkCNCNqDbCvDVHdllPYTL8ufgmWDP5CY5as3DBQPJrvwDnSMyRt/X
q1aUxsPnQuDqBpxzRvODZ6rwcdz2qQOJLR1SOFkx+OwcR6SjHkxQQQqEed9VGW590EM59EHLj5He
3oh4uQt3OC0Jh1XeC6zW/o4yR5bQg5ArISTTeG0B6WGapNLilSdwbKr23JjATbRx+OVJz9ScK/J1
7Vd+b1WdI1N4nvoKRwjJYNn9YRxbTnz5UiK7HDX6wht0gYfVgM5x9T+OGjHOI1x5nFQU2En54lHC
uHeQqzZBRZIn4sLVdD/9ReiTp2b1Br/CKPbPDXpSK4Xt/gRIuxCeqMCiwnVD9RLPcjtnnS6S1AbW
3ydJmN9I/XLkybVJeJImIoQV0ZBCD6mjaLoCbb3YS63KY4aosf93Yh5ERKcdXQRNyAfCFAaVC+ci
IB9lPpM9uptOoZ/iKX+7CDeSTiXcDW8Ep8xKvNP9bQO3RSVzIlg0A7gecVSjRtz4AgY5GtftTItx
WGEohqY06Yr4vh8x4VPX6G6U4RkF4EAi5JrzyBejiLF/OOmHZLdljhOFWj6008i1XPsi2vhPNIxG
tltmyNiRv5jrW6k/4L06kljRKoyrSeKm+46mh0g2cbKGqJali27GYPH6UPVhqrjZUBK0REH+VIqB
p9dKey4uWG4KfoNtajcnL9jHaVMQwOBihnxbcuE2Mj8i9DUo4WAR1xkyCcE1n4a9hsJr097oyS9P
a0t3LogAsgK7SWbAZMEuPl4FzuB54FLebrV1wUth6P7uJrTfJLR1wS+R1XL7GG3dE9llqgOapKOs
njobgFVdmC/vegC21JpXJmjRgP76qQ/P5oTMK9tqOtmY3n3xfrWxMcOSA7xEmFKZpUZlrDjGYON7
/GEfzVwzecavH3csVH7zZNhNh4ym32qXxLveuAXt6EUjFg1owbarytakZRIUDzOUrhROSFHkUim6
ZNaArW3DHmil+Fsv5H8hCrPZcz4GNcGV64a1ooiwBH5JL914I4Eh3XyuhBYcM9UZkMBapQH2tMg9
YiA+WeRBP0XwV4CF9xkksFWxdjyGMiJIKG35c0zuhRmLp6pCPH+duBsu0z7Z6Ml0Wogwaal/6MfU
7JcbUdelxyNFZLpTpVS8wwGnu8EfDczPh5wCDQj+QFnhHNtrEY7jYzymAXq4rwRZj9I67Jpd0tZ9
/SWX8cC6LRuKw204PbqoKy1/3OSA+DTPI2Z21iT+hOkxmNsT3SlnMQI4xC7Ctu2D7VA8iBACGkVI
+xjroaRuFOtLvpAKu2FcApFu1es3pIT+I8wE+AQfkM2RjCXAYEUwlnVq9fJqtNVnNx86RbOxU90m
wYarx5wh6/Ke6Mzk9kcBYs7CPJbdCAiCEAOix9kaPcX0EJJC0tVA7dH+OcwSLDQuxQYv+kFKaFj8
Fcgj6/no9hp0IUdf5yCTpJ/Q1yMBezrBDhdF+C4c9k2KcfV0utRWejjo9HnJSPQEW6XOn81Z7hqE
IY7poTFqf4im/FQCiJIZeS0QV58MyV9ub//mwXLNUdY5ADGUGRRownhIcS7GL2lkgqjkcRkAS1SS
w+tcHnypDkellbYKohNSN9Eb+xlGA6AdgT9VBd90iwwFjDZnk7/9sIk1kdwaW06MBQHJbo7yVtbV
BjDNpmBTaFUJEvlQjLRaHKRksu/zybLbDNFvUAh0uLNr4wO/bmTPkJuYj/1hWUZsXb377+AL/C9d
EfRaS5gQOP99KG5vvWpnUYOC55nS3HY700ix4H1mlKDfToiG7ZpeJosZPIvs4kfPk6Pjm3DJ0Dhl
uRdVzoDH2hLnfoae1DscD1Zv+Ui5jrtczotnCfuvlBDIUbtnMECSdK819Didm+llZw1H9/TRsC3v
cQDRophibEkDvDDaMafXfVY7GoEip66cHuByf9p00KYWIpX3AQrFFK2GRfYioN5y+4svJghZu0Aa
c2Vl4pvvDn0DXykNpvbXTprCqFbgLMhhhIQJwc4VOm6ZSEpUyHipMBzfDxsI9e+Th9LEvNjAGqim
iQ0wEk7GmrH/FVRDKPtsLoK99DU3WK5d5jC1s2lxQvDIxBFUYaXghXETuX8a2CFAINGh0cT75dAb
JBigZ4E7X5DXr21UmHcuXli9BqA7bXIKIpBgvoxJVZDpK0K7Q2hmKR40IxSu1Hnr7o8lW52+8ewt
3Ex5kaki4XBrXXP+3zNEDkF1tMnyrIcORAqLnYaLPMhXUslPCqQQUkr3gKjCCJapAodyCnu6jZgS
a3iAS632XbTeKWuf6DWT3RmA24iCcAw0/S8vOZPzpiXVUWAMR6DaM7g0cNS1VsJcX0isjo8OvuVC
GHjFyUZEZSuT26KJkMge2hMoHdW5FTadWRCGW2W2CSKSSvGD8sR10E87jv/J+8ahEW+5XSGfaHRf
/7F1EmfnOWqP1MYzyaCMAiAdViHgJqA/eLR4JLVDxJEFcFIu9VVXBMBhpGWL7F8+1dNc4OaNa2sf
j5BmmQUpsBkDLIbClb9yOoCBZWR73BmOlyo7zNXodhc7HRzMznhGnSSPEvpDTmBUiQ6eT7iABoLo
HQ9rE6xZ8ODzX4IFBtwgcoE5UwcmgKMDnqNzIkD3zY+ExpOHj7L0lYNGaWM4+4WkkBiqavofEb4S
YkYjkkXaghM9O+lt1lzwc0kN8n2jce0MRh5kTqBQYur/zZ5GrZRYLojQwXc2yMhq2ioxeF+ZXS8f
uztq30bjl5ALNTGQ+nBYKqZxaA+yhU0SUOnRW2a0nsPXXewFlYP+Joiub/c+lRHFKtfRbs6HsiN9
xGbt0rOoai7SAv8cQZD8idrp0ABMPba7X355KhcpSHk1a3h/E+wGEmH0dhd8Mw3kGyb9NM4HId3I
BVAwjcSuifNjcSJFuoVPbpC1lGWQidctX/TiMtchkFBWy78ZxoUjEZWxm0yXAHoqLtGQp8nGxSuS
qYq/RZ4IY2fNsaigzQ+QfuU7fYS0j/Y/3oEjn2GGjomhZY/zMIFGIKQxJfwGnRrTCdtQQKWcqZSd
b0P8qpQbjIaKKJKHBHGr672a8Y6etSHopkZT3pd9GfqpcIX7+JpkcYV3iqTsBDBijlYyXRYjJRvr
cGveVre70VL/8jKKNnz7Jfk5BBrBLGpQh+CUQ4g3pSZ0OdcN5tZ25Sy4s0lc+BCWfhIp1PdISLI1
59PdoPEzj3/Z5qG9aW+8nxhhb62/HkR3ueplOtcLbKgVmZ4lbp/MQKHxzW+BGBOxEVwnCjLZS3s3
Clpw34utxSBRMMKGZmlQpgiZDMNjtYSqiLHKsy1uGOlFYaRg2blDFlcPIoVy9E9bDw2xfnOinkT4
ccqxlfN3B66Xg3tKJerxbWGZ4GT9aCPMLoi0XOGXYaL3lOlDaxK7SDiJXZ7BQPRpkMSN0Qwk231q
VHldrLmUh9R686EOaTIxYHqkRHadakEQOHcDvLYoKS4eQOCWwiHvYH4jJ1bLsiT/oTyyCqpZnEmJ
0A0Jqvx1Ek5XihTQjbCNddItX7PsA8/19EWoYTHC1vPkcCAWvCD5TBgL/DslJdxdcwMdnoXAC+8f
TEiLiP6TYNI+h6mdeWODi286rqYDmx1+OGDmCSAq2lRArprLXeN0NB6gM5YL9IbrLrQYKDvT/tOT
oAb8H5/h2/lagyLCmtDHZkksV+hQocKbtFqd+kmEGj9yCh3bSGcZbfE/B94XEd7UPVNhIXCE7+hP
VF1iyVccoKLgcOna7f+c2eRlAvhYTpvcFMkWuSPFk00hRXECr/xc1iZCZF8/6azn1ubrht2//D3g
PxcKPQeLs65l+e3Qbtd/NRhTuBSM3A+Vk4tM5ff/EJ9/XZqKyp8i0BbElZxkOlHj7EuJUKN6+V6f
53JRuL0SvnajQWORKHzM1gSKJOm7Uz5HiMMFy5pi2S7qrsiMb142L1m5xQQ6R3MwYukVPk9fJxB1
EPWxh+SZ+Ga6ziKcuJG9JWgaMBFiBloVOPlGQCpm2UiZqpkY5RUTllGaRF2/Yr2BRx6cpuiRzqRg
wxiZ7QQaWefbelJWqMta7zJRt+wR4r6aVxK+QDe5l2O/dOQxFErg2qvWs/TY5pzqK9endsqM62Un
uAVmUEsoT5Bp7bSjsjLPqjJLMGGmW2Oc9BB4w/5Aes1qiNWT0Uq20yJXtJ5MW9/dNx0Q64s7nHd1
SY0XKW/sgG55hnjlFAgPJ7frjQSxLKcYS3+C6vt6q5YEAjn7+OsQxpt1/M+lvp55gPfFrTB2gDU1
RUK1AK+/zdpIcQbD32Kp7d9CF8Tov7j446nodaUH7cAOSuBaPq9Zm7sAtPdxrgW3lnlPzbanIAaS
yPUmlZZOR2tS+CRbPyjeIYKrODeOeSELUn+JT70bO6yN9qMZN3DxnPxyM7ySVXdJaKLsoHxtLToT
10xJAYf+ByWZePx8wlPvWhvCdeap/xqnw/QEYpHZHeFo1qQ1RwJhlGGfd9m3+cf1q9TD20c96kg+
1mS/TuPPHj0yGjg7wNcDOS7BySiF+2fTUBFT/pVIVJKIsVHPNTyH/qPn6Uz7N6/DIhpd/baOW365
tXNr/zL4lj+cq39nHDD85ntJf968wonNC3TimDkdPa0dTXo4lmWsmYFDSbo11sXZWmLECI9JjBwA
83uzUgwrCmh8pVRkBoCODx90aHKW7DllD80OdNKW8cy55LCUnSbccktXEdeKQoZUsdvZJbF+hwRN
KM9mxzzSi0iqAlafNwH0lKTFutbqY4yjUlMXAwlhkgnjuoixH5IEGhxM+5/pzyhLH3nLF/mt/HaX
8+4ILESj4QidKuQpIKTw7AOVp7qJpspVbKlYlK44gP5raxpZQDQHMTCFfdcNCV+OKM9FiRJ/HTvO
aQcbnejaNsOlGOoCqA/9zQRzOz7aWIOIp3iWg3Op0P/36/xjYOO61t9zrLtU2wqQ6wDXgrHNqtXx
onJmbeVFEuOYtvz8nZW0dHSYyDVqD2txyK6SxCKxn1PHtxdb682GEUJ+uFk5QOq5Ox+PHwpqY2De
pYX8EtckC3CWf2Lmi3v2rLezw0iyMso1sK8U7qa2mPQbKhfQXTMPpEaFE5OLGHb2IvAtDBREbQ/O
g7iErz1102BFxSZSIwkMvumLcPOO5ypsuDiA+3y7+6iG+Mrp6gsKzd6cjmZJ7JUOOVM4NNygtj0c
aeTD9nlHDlFme3Zb2tftMbkDdTapddG47O3f8AwOFvhrjTcmUjnRJRb49/iBegUlOWcggjA7MSpu
7wns3XOegNt8DAX/E5WZkFyijyHtF29eHXmwUyEnM6jJOqS6uhFwuA5O14te6JFFaxalsHenl+Ws
50miHWI0RLz0LsTMsRnsx68TqRZsuPqe4pfLuCr2HRwtmCh75A1JUGH3h6xgmP0H1+LRf2dSRU1r
IkEdh+UZRn/ueZAlRioLdNxEYhN3NbA2SwxSYpGz6iLMjqRKlb9ocEBcs0biZxvybbOib/gYurxg
w5azLlAvxJncjq58BiybRyQ0ARYXS96n+JqCiSuGUTIBh1KAMPh1AU0SV+sZ4al2rNXnP47T4piI
iU9l6OkBZMM8Yz/W079airk7IUQxfvS/q7UHefeiwML91KOaZEBg2a8JdrqtST6AKegXYz/L9f5z
60uyZ9V6KcUud9WHk7npcjhQypCVJs5IYjLAALPj89M3ugLavtfUJgc1AczzB5/GajFmO8Pq/1px
12xs3rWCotLA5Wfs2PZShWwv7/oBYxF3ajLJXneK1uUgMC5qzrAiQQpp0KASo0qmFnvUf2AvOfmL
Jj7dYN3Ta+waMYN2MxqCMA7tmBOgSdJJJsrIcnnA05gEF2lA/M0yn5LY0GEv4Fea96Iqcsy2mHV3
qG2JtxfXN/xmJeFGFtk+jZ58oHWqYDFByM00Jr1S8MGvYUfY4Czdl1GZtoUcRH+pxAW/VG34YS2F
zcFGDVHZlSrH0W9QmN5z8fjHrTEJKVcfmHu5YJpvUTZUHQObp6M8Mrv3kfwS37LejGch/l2yO/ND
uJZBIDyyHGVcSVz1LdYStwhNsftrWhB7uMI5jgzTXjjC46HjqLneq/HJWy0D0wi5FIiXl4gTF5nM
t8/htfjgHnTG4Agw8RWUYB3uppiX8A7f7+06VBqLOCPY4qnf/woTZJvDU7xHsSzNezQgQbISLj0o
FsasfuC64s2rrwT0wKlyS/VB7OHobLZ/UvfFnk46lzyEGtTfVIfkoa2lWNhNRx9+Ba605zZkrciZ
6dwL2G5CgwJsz/zYvPq8lbCaSiNxN2C0C5T43Tc2b8UYm07mNZEsBV/fiaYpo1tGmxKE/f7hRMxV
BIgwlNz/+x+UaFcaSityswjLJBo3a5PU3STIH2Mct20zHsEuUgfa910KLA7hK65wPvfwsG2BpY5n
mgKUYcx4gr7HFw9tAC2hxSdZateprPIge506RTHoTlEhZ/aXmkGkqAIAt8tV7XIahuSShCFeDrQ9
2FaVW18suQY6iAjEGmjEdah4FdIP869pdArhdC956tVs+jarHwRsyTWiDO0KF/Dh3eoMeDmjFBpq
zABpPgXmRNaQZbmx9T424/HFg8IctV13w2fxqtp2cS006yZpsGJfGBjMoJdWlU/rA7/guSHIhYhs
SZsW5py3uuqZe1dlTDFEIa4fHHWdGngTHDOzq4LjfA04F4FkCtlcwxrQaZBFewdDueGSwANQAb4h
zGpWymZl+ZpHex2eLtH2EDl2MWI5bMdPB5e6QIr6vlCnD1eSadKSif0R4QUr+71cLzlisXRDXtMF
D77gmzd2wK8jRVibBSeAtKIgn1HdJfr0EgL3k/IKT0JSQPHbUFzfu7Y8PmwBHByzqe1OhdP7VIAJ
l5o/0202hjGWoJIGNInsmQKhD2Ny8JQjTwFfjL1zjMXNUW2J1nyFI1ZqQO7+2+ucXbWxZwwps6dd
NnQlpYTgPURy/vq+UHUPPPhhQDf/rEsA0+4HhMQYrLziprsyIYFNINUY7kIuc2EMFxv1ACQrngjX
GNsWTwz3f55GzN10F7eK0PYyYdwHogYKbvjTD0CwW95Ed7Xgvse8Cq93FkKxlK9vgBfMr4w+ZV1q
YEZqWCkB7lDKF83rvfqRPBHbLwLqfBjFConvVR+z7btjfcUINVo8vGWMjJnI+YCBdtic/IeVoYTG
RzibKmiUjLkXgNs357zfRDiehSmS/TKwhEl8mf7v4YRe0NkSxhbg+KgPkV3A/evA+lNBpLt/fWU0
IDKCiMUo5cDZSKnU/DRJ/kWKi+u0j0jmyxC+bb6/KWls0x4lAGkLBym911Qfv1L6wDKF2TTRQW30
6YnT463n70SeFUc7bdncVniVRSgxKh4U8TPG96qX6nPN+rKB84j1QIFI5BpfYq7GyfTuclTFBQpV
7qR5RSeuVFmboPTU3mtFADg124nZQPrunUtgitIERMjZ+DCaOUNpd1tHtz7Xmb4X/2NFP64/WxK1
+czDFk3jY5/fSGgAoTGi/ja9BvhvAU3h2vOqo53dW1+ibm5R+Nk0XKDNGh+YH/mqI+HVyM9ZQp9M
+uRFtEwPIy0DaVKnbtjMytnd2ESoy5aJA5abOk0YGSbmrzQbyLteRo6ropHWiTfs+AfXwl/d+duo
TFhFB7EHF7l3AZpnlcYHKV9vP3D/rmmwduJjXMV6iky5574cPEFC/mKa7Uo30rq9wyUXgsdAu/US
PN/+qpVpTyQYW/tl5Dx/bhe9kx4+3JhvL/6PFMJCCgmUKOQuKwSCwL+SRzJT1WfB5LblnDf2E5/9
5gf0e2pB6A6AQSXACKwlzVXuLMcGW9cEUAUc4/tF/FGKGtbP1V2xRUZarA1UXM/1IkP34k7sA2O6
uAwKXtRy0S07RxB+4crU5MBIt6/fPNyNwKUEi5ECF//dFIb0/iS1BcNiJrhx43KVz+UimSRveXgf
gWLyTasqebwH3zNKaxAkHL+5MhMA+yska12Ur0BKCGqNlwtPzVrZfxVNYT6vcjy8AjCD4IYN3yba
txidVEvDVjPsCFcrNh3FiOIsA/UCcjo+kkVofPOF3CjC9Q1BYdHbzywiPckRhh5PCxKX4opC5A6e
zFFp/tQsvSd4pbYNAuBvXlSZmQh+bPzmSL0a4FMqoiKVfkyMxMZTz1OS1BMtRMe3a/nCLAbUxI0y
gXEjvUens70handoAH1vnjrT6Xje6Qxob0RmbJndNzv//vyw01pKZns6XenBWvrnJJvTYFPsYSPI
ZlH29QkLT2h45jmiMTzIWwK3vvSKRr9vhHPAlyGjUR4rIzjnBfZ2SoFmlV+JYowEmgztoONdDoV5
lY8/SvTx5D0IRt2gatuX+Z6cJJndR53n4fWhm8sI+695PhrfqLeWT7fD7TjipYTX+yesAdLqARbb
TXpNuBsvTFaakIsI+ZVi/9IkyjvVA8lstZrZI63TYwbEgVNEZUsnfnfyP3OX7PK/Oeaoxuj0o3z+
D8IMtAyz6h2xMbDjEDr0QlESRWkyguO3IbAqtx3CBqnURT43hgC3SWtDU2EHYedCj9H33bsH59F/
1s9F/SU1kQlljYuO9nn2FTL72G1qMtHPxKamt4Cv731zq5kY6kSLkKhftAYhgKIQBt8j0Plb29z8
KXO34jbmDma/XhmNRkICp4NkaIJ/NiELUv86b7xpdm+MKEHA4Db/+z108fGLhPloBgV1sYLsTp8m
/8mPYeQgptT/PSFQOR2A4de4MxWRj8V3XihYX5sSpNiThh74qbU4BZ0DccxpTJMuudLa8Xk3Hgar
/t0RrcXIlFSChtZBuIhrhFy57xMwIl4gmpN8bJmXpQ2koK9l3w0NdPFulzerpNAEaAlq7gJha3Z0
Bqx5R6jS4rRd4t7+B5dHYKdCDM0cxtktFmjo1CpsfaGjZ+Tkb5eFIkgPHXH2uad06h0gwYBGufKz
HCfNxbIhc8sKefOmiKs0Jg8HJ+UqTEeQyMO9JJO5p9YyfmqJsfydG36JY9mOkkLVYBTdMqI/f6KS
UZbo+o0e/DoZKPRwF49hhCqBBW2ldqp4fOikGozuNgzVKCs1ToGO7qRWKNZpvkDHCilGwhDmg9aC
2VDWe/EiH2PLZH3cfCs2q1AV72jpbO+97uV4nmrPj+37d6/Iy30OHca7KrK44IFHqgBz8BckzUx7
tC+MhceSLMASLWmiMIuTpxcaDG+JKZSeWbiLgY9Pth3NjkiDgp8XI+gnW/k0R0g1RVCRDAAQn4+6
/UekozTSB8saMBqzjFWHf/IltuMfuGBpi8BTbtA03iOhnUG3Nz8Z+Fl/VN+G8LPrGRJ8z8IcWzOk
bAF00gM5Gk4SoGDm/0C/lHz90lPdRnVFYTD27GeCr84yPRFYkXyGLj9Kra14Ivb2iwozQF/wfU8m
KV9Ozi3TuFZEXryBStDsmH34XZrypKsV1XVEdua14UUy8X/KK51YgyzYt9s+zIHLgfS6G1BIUicR
cQ/4GG6kkWRJXgbLJXZ08+ruar+Fo7Zb02+7a6Wa+B7UviMHBFCnOoqZhiUMbu3WHQxeoVs9N0nC
dYStvWPxKjk7aU4BpUzhPHWXzC83CcA+srH+uGZtzam0bpOQGwdDZngsnbU+jy0yTRtB7/+HBc9u
AJ4mwpVGOD0N0jHqRdhn4FY+EGS5SeZPVAILOQtAz1OZvcmfnzNAmwgLHEXnzTG2vlnmmh8WwTA5
vYYZg7/Fl+RCGToGLz0+lLFRgWaGOJ1ouZKBJtry4DzgBNmL2HKwmqLD8WL3eG2kBYlLLCqAk1Gi
WuDOYyXRD+/GLD/Vw2N04oGBEpzhaQ0mr8W4MgvTVWQpy4krkGam5AII4pRQuh2pHM2MhNNHO1kB
TGDVt8Y7Li+dutBcRgSc3LNh/+kLhW7EdruTCdhpnbQAvbbWxFpiOt0ViphSJPl28UUSYEtFXIyc
i/hXvU6s3OXotVV/647kFLvRsP73ur3NGgI8ZoFJ+7jr+IsUyRKugqmbUI4LIsRMLZp3L+q2e4F+
hPP55o1ZYDSkAAaNIOt15U5etEvoKim2z+LzWQQXd7EgUhlAdL1wgT7ejxGDhwmcMIcSwr2DvN4U
Hkt1X7sr24ikzCgcwcNSd8ziwU24LQShIm5NmVlLzbvTU7Suk00zHva1Nsa+hp+l5u/LV7U824Lj
f+9Z08+KFHs+34Ls5y4nzyoTwISb2qrMs6MbptLNKmEBjbLSjotdxnakycJOkJC/juCq8yrkiuQD
uBd9IBL/Dxw/KoyditLIXCOxXMDcX0etcD84ktH1VrYP4m5ofp4TPK5nHRlMOH6SE+og/GGrHSnf
eZJBGQq71gFMhuz0hWr+2yJlwqr7lN40k9L/MwamhJgdRyDLmGCd/UdM3naMammX0xIbMs719kC5
F1RCADF8WzUGUdYwGBvw3/dKwa2IeMmj7HcD5W/uBqM6FDoq27eHL47s40r4mKWRETZTh05ebDjw
UhQGOY81JRxz73WByoNC2tUUU6IFCU7IgWKKYQFQsIUI1VYlmjSLZC7dxwEYIsKlRyYpF8LuLnX6
kXf2bGyzvGEAUJZahiqkBkGyJsXGc/2SSCvgWIfojPbbpXLNKoqN3HmWy7ABOTecR3jfs4/8Gk9l
tktK5Xiu6H0YeCw8FBNKXOjqb7nKA4QANO/xkGSo70B7H2s1yI4wFndMtXmWdR81aviZHinb5Bpd
rc3rWxqF5KJYxORAHPfI1E3LZ0nft21E80VB3y//RsQZxdjnj0XsQwOzmMSn9zeOc6hOdNO48rMm
Yw38lkUBFDBvF7j0b3iVYRNC9nKxCG+mqrODlQkPcZuZYd1wfQxE5Oa81a1VIVTOQLWnfBuVxo1d
GnRJ8Xbz7vSqy7ynf3p++rmBe+mgj0P5n1sp8aHuDXcjHFFFGXh0IDH2aW3kpVcL4Ay1b0NTHYsw
L+3YTo/iKDlJn0Vaz9OfcDsBer/K6xLrb+upAeVrunZ0PAbCSNUFlNt0KSUtsDDYIkfVLmh4oYbr
5Y3nqryD88whP+1KFErrTMcz4s+S3mbd4qzbYPWnTajZBhUkYFeB8cmFJEpOiPPstxgCpYg0LFsj
Ed/c79VWsaP+SyHk9FkgZVAvOxKF5IXrZVKpUQ/q7NNapjqVG0xjmLCJ5tyOo4jaVXJ/l1wRI4x3
/yZuIakYrsXlBIPVqAnVy+ZtL3JvC74RInD24gJWwJ9rUiFl3Z4ZOFRYWo7fqG5XlY0VBoZx6aeb
nVOO1QSJHnh75RaX0DqLKSqZryXXR2K0YQMKcjHaJIdHnNLDC+PoHKODxLn+aq5oWECqieG4a1o0
CfZcVys7FkwEvO1SV208dlcZInlsz1sTr6m9DFDWPfAhrUTfOirBptHAogjazpD5Ix1BCQEN3vXn
OzA0bOTAeGCGY5PdZIU+Fk1PBGgCIIHzHJaBhtG08DkyhoEIiA+p608WJdHiBMewAZ7h6bfDE5H1
NVXBiO7pYZU+a3mEM/a9xkd72wohMsU+5PMhSzZ7GMWXXDAO8MvHJBSsMXRJjTtTFkqZpcWujHLs
yPTxt/DxDljPlQ8j3/ME7POxbM9bSPt9ywbDOn8j8o4RQIZnoKsFis/s91B0RQ/zjSFQtV6ccuBH
RGzGKygbV6ienOYxY3wTazfBUfEzPP/LKKnSTokz8W2hjs+UY2xwq25d86So7hM+8vdnTffP0c3n
S7/76FYlxnnjzavYUrdWU88LL9CHVP4XxJXjAUJoo3jw7gZ09Q6kw6UjsYXs62JBz6Ao7jryA/P2
pI2PVlWdtxBqVWM+OBWVn1yTsitYAFogvzTwvyoC9l/gk3gSUdlHgSQabaQl/FIj2AiEVhZYOYMg
lO7ZIlcFzNzT+lGvqMDSwW/XgReXPcdcN+RqfEIz5Hu+15ZQY4wtF289amoxVrNZhr000FDNlLAI
h4FGS4vBcRgnc7+axpD3AHL4RMxb+NwMsgIplrPDjz7QC6KZuTsw5VoJivoTp0DHLC+hGjPbeMCW
q11WE8/i7EEq5WOwwfYE0R5b3ZgCuiy86aXC4iz6LuNEVGlsWhLR9J+V3IKfMB+a0Lcq+Jm4ywKe
lhsqBTPwzqk4bUcLe8SopRBalhdmCcLa+eI6IQsrhr4t1EZFh5gJ8zyqqL6pXz8NgqHMmd8PixDM
KxpU7NKq2mlfSqIui/H8zvkwEvwtOTtxeYST9qJGkEOXGyw7VO0nYg1M7WxJEPKOV70Q++vkpgOi
9XhHrYFFRmvnwaUBaiMLwshQGBFBmJXOFWXJhQdQ7GFG+kNURPavgNbwZS3quiTsDLRQzkyxg4P5
Nba6gkgXv3Hn/hQXgC62MpRlnDpfWqeL972B2An54EVz/+Gym8c4aA6nmeEUNSEbsnapAH9Lu5hI
/Wnkrh3LVHsWPEAqEHPHuyyYKCvnZ+E388lvy3sueqkEWMprQ1vpCs1q8hAX/n9q63pxSclYAjMd
e4et0IjRQWQHXvvIHZlMK4LILXBvp6YxsToM2hgX3SHGsSOKXX4H4usBJOhoWEipKEbEInyo3HmQ
BFZjLwRz49OVirj9ABhkHYnLObA9MTz7fzqu6tIQEWPwtE7gVgvG623meDnyTAE9cjbhMcmfNfPK
r6u0BaN4zJOInPDeqM9QA4Oy+HG6hzZ2OoHOnlF3jzTtoFo1Hs9mRLLBSo7ivIfV+dLigdnd8Hmj
QilBZoUThSzuU779ExaM1of3Pj2XlRAfChuwobBzuTmBQ5RrmARHF80agvk6Ly/K5ZlPGfwAx915
b7vcDvRzQmesc87RW3bIvDDX16Ac61sdunVvVnVdMhIUb2tHQ675ul4a2Z+BRGzhOKolJyIO23sn
YAYLIyut1ubwnipI2f3s34Neog6kgwpN5SEcB3K5FUE2S9/tlvjxKYLRBUQbPfU1bjNJ03islmbG
mqLrrzZbsoMbtTTMZ/fU5staEvuTUYfUvroJwIM0N7M9T3VXgiTi4RXAfoiIQVxaG7c2NZTgUVC2
g7cIv0EapctlmOMXQRX4ccCKd7wnYOUJImhlOLKoMvruqA/d8ja/4EJtVSa1CHxb9TTRy0uKRn7b
Ju5w5NdvMO9TcMisy5OoOVmogXWkZfRjjGgNvE9cYXE2njzxffpGIldk5ePrmbjf7GvB2m2Nj0ji
+uJEnksylXOz1Z7UH+6oCagesbnbvUnDM23NdsWhb5D3FMYOxTLk29v8K2MLz9VF7Oo55bRxl0jn
UF4bqBLHE3qghHTD3fQXYgPl7Q6G3CXtaGVUUDFCRBivK6hNOXHHaI22SIwWwBRJlA+oR+10FhcA
DBQL004l8BFfYKw42c8PNbil9KRR8H9GljWdTb3FSvIcA0xsqNxK0ts42HjdOb/iGyQKlvYD5v+M
58mr3BOlTIaRBOh5IYzratV1jkl90T+dueDYOUSrgmLkSbykrkblzP0jdLXfAXvPjAg607Uah5bh
MUvzEupebcBAcwiNVoxhVF67JhkNaxnd72BFAPRS9c/QbZVfGq7qEB6gYO3lljP5YUhUAMJXHljs
URzMo955EBqoUQAmWehXTf+oLdbW5O7Dwj5HcHPWRWH6vOgw8uQZNCxqr4oN0BeeMLnVfrYRWJo5
c10tgnxMNP+dnjX3DI7I1nGvf/FQ3cI4wq5eU9YiYYq9Haq4xxe/fn5ZdCjR4mg/jUsoYK/7KbXE
1dFzYzGoRDfneqYuZ1rfclQ24iOfCopFPN209/MlLWewZpBSiJEL9E8F89N5OlQdfcCzpsBsazHB
e201MI9RTNdAlo2kK9bNOYgpjuqeJMqJrTN5NzXZKgCzKiyAl88md3xPbNtS8fswbBj6aoA+2KOn
9b+coQD8+q510t2yHofKMgYj39DHFp4Rr8J6ze/gZPxJHLXEL/EFajArqMnaZTf4N49kRIDGp0pB
9pwSsFg72MU6hrH1AYNI0sB2v3OEfirKwRs9OLk4UzLh3ieHDjeNuwxlpJU4aaljqIr1Coxjh8ly
7S2ETmNiKCliFXJXaXVQ2sRdQeRBtJ+JyBEeOMaZthuPezSxIntIWSQncMOZa/pj0KibTi9TFZJM
pWTJiale1ydDo3b8cXfIfrxSCRkE0QmrjYSLCzRO47dVQFtrqW4ktbh80iGcqxPLuS2ZzBXSOO0D
vlB1UWmpfOd3+8LD6gNtodPCBGniO1ueT8NvJkZFEJx5Sfu8d57XLGPPtOgNvL83/PjgxeYo5JIV
tBlrIt5AUI/FwYdE7QEPuPEFllwKOixPPQP4QwbQnykY/Jp0HxKL9g0obs011QE4ZY3x0vUIUQnp
MQc45z7YwXm8zMh+/Xgbcd8zFqThswjOspKhsE/lwfh0vE86oYxPf0Snmjj6d4ItGTuen621BybQ
umAQR7dUwklIVCYA/4EzfNL/getpoOKqGa/6KyK/QWlMuxeRh9N1bzx0SS/nIzUfhYSyt/Xja8VL
dagq+OVekezDHn2zwORQHY+IXs1Il9BtRufnK6MRast31IMImK6t1N+XXTPmIUjkZNkEQE6oCF/8
pXAubtGhgcuDk5pu1ayIt/miuqv61EtS40C7HpGQ1vQC6ng918opwgNhMMBcVovSSBBDkPJ4ty6Y
3w/mszhlbyy57H3mIVCddP8p0ktu7EP6imlruOCYUojcNJV6CAnkGh8VYi99vjR4vozS4EHyRNqW
Skm8Cy8MvznKqK5/DfKZiyEmzH2n9W9/FPfGQvDRlWvsSu/nVrbRMrF7o6wKZ1U2yXQBYQrQg4Vl
XMVe8Ijz7zMy6Rd+ECrAh//LV9M7mYFkcn0TGOdOuiWHYt3DuyyIJ87u6CA11F0PtyDlwxCzrrcE
Itsp8Wo64Mx/fVYO3zAr6pk66fvGRZ2xjwzGAhpqxFU3ztUm9ivkWmMnSY12mnXyiJ0GoCfxg6lR
ALiQ+n9JYd64A2Ss4D9O1hujQvN/GLCbKpstt5qYAK3/sSriXea2UQbFAnIbgnh5X7UQ41aZJs/m
h5gqvXfmd7hJOeqCe9e1e7AWBFqi4DQwewHgaU8Etu9pg/cSlTC566G2h/i10JGmKV3M5IpXy9lz
1O7Am19j784OBDgg2Fan9TaLPI4veb0+sM/Ovt9ArC7WE5yxd/TyNxFLmTKTVbV397IhKEqk5qdn
2qmWC+WcGSxtzHF4Bq7x57Rt9p3SPIYezulfRg9/HB5Sf9Vitxov/k1KKBBclMZSpKTvceOgSTpt
mzogy9BlfVN3vZZOsN8jtk/TZR0eap7TkXFkPWoO/kyYXBAY2RJx5UlQ1VCoAdcfxPkCwjOwGFas
N4KxfqJb1XAotpoJYTS/X2abADMz3jafGZX6M2d51BXpfwlI6wlVHkrnzKpFY5Zr9gLmtr5GUtEl
FoB3CY6lT1ib8PHe88bgYLA5y8g1oOSJp8otw3KjQkWPz/YSOGKzadBL+jPoTVoOkmeDbNkfG/Yg
wMbgwCqpMkA7rmPkVhexUa4HEus3OrOHSRSj6Khc4PLwNwY1uhbEmne69VPW9+PpkPmYXzmCvMX4
5lvcb/O9YrQSoJLmYKgPPAitETsVTYju095POhHddb3pnaTDnpFoTmCdvj1O1IkUWeTjt44fMwyY
ffyY69kAwerPWNYdMZoY1A4ExkE80gTf1bTwNX3CHEepPntw7rgmWN/ffWzNwqCIS3o/I9ZAAf/X
Otg4wdMe4P45LbZYyyJQ3RBdkvoaSEmUnsC/yyaeNTbsr83a85aHiIjtpCz9P8LVTNhG1o6T3Ah9
wdMn1WrWodkmzULQZCE/B1Yb4qH2eZj7iTJ9KDfLlX/dPGHb1A32p1AZ+zi9recQGoCUmYTSbIGS
e5+yT+0oVDhz43J0gXetJVF8vjMyDtUD69sasEVwbo2jQdwOeg7PTElfxnGWSuzKIScRX3/5Jitr
XWGNtClR+SPSINo2By2XqJqEu4pk4yG70b/Gy52tt49Nj+s20bb+7cPchqBklFeTR9ulwqxMzEzq
2kegCYkXbIP1lBEc/eFE7PMYLOEOQE7SoGZl5jLDzvgKxnYvX+YNNoBRJIyUu+FexzZLdj8c+Ogp
T3Bdp5kJHgv/EauywsCTmPtaMwSHEZxMqbPplpnnM7GAVN6LIqnd9ZwRo1irJ4PkhHovx3JRSWlh
94t+NWcNL5InUddtJIkcJlCb2dV0QUYq7ttOoCZqExCFsqDxGprMJXnUPnQcj8VtAr+Qwi+vaZ5B
VEzFHV6yybTi+tIwzszNeRpmi61Lzsam7wibQVLczgEfxXmtUA39sxjYgR7jh6L2tk7Bh5WJuo6A
0xTN/CAoFatLquW509LRHLFdKwR0p+dX4UuwDnOYbwIWHtaWBtZZCnQwIX+g6vMOyRUVzquCkOQb
cwFwrzJklsT3istx2IpDqhjpy1acwk6zRWS9hXz7q4W4orgZLVxAYSGuU4FCWMFCdxDQpKZV9nKT
cw0PUdoLGx7QVReZLcLGQXiFX4z8TrfBKOwk+5JyGMED5iBo1VictK1KE/jp4gs+G82hEzSmX+Af
8BzgYnIURmLsqqC4wLqhox3GNwtGiYkDJ+zAN/UOnTSfRHL8zLT7al5o9Oly+aU4S9ikAHKsy3pz
6VVZWPv1SJy7Rj2QXHr5A9fVrOCzEzt1hH4exhUczyv7tEXz6HEAq3iBsQiU3L2KX7Ga51w2ilhv
ARbsSC6cL+nNerUeVxrV75O2Qn1Ay471XEqk2DFbKDut2nvznZv1FNT7hnsd3gfIocr7sUCdTz8C
9e7EnDBfv6rPO4i8ioq1B+Tp3St8KmanhAXOZ8Nc/SQ+mWrbMfgAbTKbdorhQIlWhZbghX7efTR0
SN8yCgtoe7UcHjZMSF5xPO+++PCux/YkHohSvxXw0OOHv4+awct/I5mfgsh9qihu1qPCJIvH1VRW
yMsUOrd3e/3hPKF4ljp+OfnPgHhHdQ14FGbCzsAwZKvjwhylCMkSHLL4DGZBlwc6a1ZptxKbFnC0
ueHPBKf+MBGtC6tRQhGHxwtEtwnlQJgmxLCFy8PgRaeWAXSEz4W9HHBhO1cdYnoWdt/zeMsyaDyT
neeJ9preW5rA/412hlyu2DSENR8hHqGOClrRn7O2Go3xyi8Vwq98TDf9BggjRd0wGVGi4tcFi+mB
8Bdjr9QWDlF3kIf2sndbkFgj1tn+Eloaej2ZXqHJkVxU0cVQHZN8n5uQdj/iNj+cTlCZ+QQIzGTy
f4x/DE8r2ljpKs9gsrkFT0cDAuvdDLR5s0oyr8yISTrQxdP2SmRaGK/AM3PEJPTA1z+euJ6s8r22
M1qexP5Dr/5NbT6b18jTi2VgpleHHbqRrInfox2V8igSE+lw2Yx6VRDVoDAG+M3d5VLxUAMbbYH2
AoG2GsGFO04C6KOfPmaJDFGjvwRHetRcGQNJfFWrvGN5h7VxYAacdthDg9d2WgtOB7C1mbzGJkIK
U7dyj3FKAjNItT9okNl/4hj2uQr8h7n7/mNe6nPDJeJWvSQUqttKDR/uap4VFUKeLzOMemhaUdfm
u++oFoo/WATck3ylhzmmYiq3TosLsNQlPR5bTrawRjk3qCBVYrUzifevWf7Ii4aTOP5xcFZ6+FIw
ajzkhc1Iigik1/2Q077mSvmqdUzI37Pcgcgjv7seMgzn7RY4/h6FEQyHF00QxiudzqVseksYT+nS
gKtmnGDdAoWJLTlyXH0xXNGPHNn/U51UzjYgDmSDFncXVZximFl3RymD4l34SrzNSGSb7P03A2Ix
JW7pkDDaB+2ummQElzTqLxgO7Oguocx9IsYi+/ZBUbS/JPPwaUiGIqcUDZeDDZT1rAfYe08a2LjS
2sPikMhlIThtKRzHwZBLdBUypatJlLVfz655aS4dJoAhCyk4e5qtFzZdxOX8Wi+R64a7PA15xHe8
qfIs95CznVy1GjnRZ3bKqgOEd+OZ2rnYS5m6hyFxHW7I7ZR/5AFb6vCDxumtt739xwfju/x4FvEq
y3XkMMJ2a45sPy0Pm5sETTsxi/0bN6B8LBp2afgOBxuOoRGprYhbBZH27Y4mvEYt1YCdTCy00+CL
/XtLmif2zgDEzI5GXHQc+3sJ0+tAt2OupIZO0rx5T99HjDKPYHALKcIXDY3xlCX4TtWOj7i+sqcM
2c31uRAf0TRJZYVsKLOMeMR97g/30sugqmYoJYsKikHXQVuY0walKHaQmT01+L8Yal2wdQTWlsho
9stJnajOpcSKDJGKPh0cKtY/kbKQluhdOWWd1Uc0QPEK0z4rtKAMHU33rBDJ7fTFQwFRUYDe/kam
EKAVvF5DXwdoCHs+YRH1P1FlRuxmmFICvRZlTf0R2hLS+HczRONqC5ybKqr+yLYcFKCgZwx9SjrX
nZWxfXaqNYfTvSj7Ga9+wcRRZ/TzjPrCjrdvi3Celn9x414xPk41DaowZJCZCC9C3Dd+IoVOn4g/
izt0hQIZQL+rF9dpuv5Qa5YARJhglO4UNkIOQKthxtCOuyahX9RUKx2r8ohwVgBPq5o70yqAGXyC
mM1tnOZKjYtQpYLgMBEgdyy7VcZ8Qatj0ZB6wlZR4Dfk9ErMr3S47cBS/mqEeiFWDRImJJIKtmSS
gVXJiSkO7tnELkdB8pYH45RCp0a9yUHUu1V+bsqcxP6CIGCfhzSpsEbrxGqdOh9WCMJaLSIDsG91
vInV+ihio9AHoBAMzagCsomUO0X5gyUyW1vcw1mOCMY1xbQ4Id9pPXjcvs7Hcb4IHqdIEU0VuhoB
+aMLlWZ9q9wD8NwUGaEMwJYdj6VBJTYfzlFQtfP5eta160LbT+lifiYqSzYWZMAgG5LZUm7T+JI/
jqGP0XfcFLzTZHZoYjwkAKqfvuZgh3oGb+FGs68NihkanYvXVNByMtf++2t02C2lmD8icCYkgLbW
ybgxyMKruA6qc6VVulzq46j6VzAL9lv7bRJUwe9z4e7RlT5czlyRxclMoR3CC36xIlrRn62ksQrA
rNzMhWBq141Z4Xwut6hQHRKdHwY4tdzV9ZgGkUWTTbqCiIlrF2wJ/3NKf79SILFC2tFPuAo5nRyH
4z0KIwk7emO4bAq5TVOIxkM9kXExvUG6cOS8eaIoSrWelnNEcsdpV7qAd1d58SKkZhlerDhTkCat
N+3nwRB1IhiD6YCiBWQVvHUmJJHBWl/gFW2OQWGEdxp6zITsSZY5kyoAcBlqxZ3kcGyPHuUYrWui
5Am1xZ3GwzXcmQKXO2+vgRF5V4mN+dwkxEDUUAuYVfRrszPKPQmcY4LBTHr6m+VNFXAo3bh5QZGN
M21FjUS/uiTpYEqdmfHD6ZzKwB97w35qVqOTiMmKYjRSIMwF2MZ2zodjcbHnnNXGEyRlhpMUgFvV
xQcKzU7qM1g1OwT0390EmGRAyIeN6VWC1UaN7OOt/79ZL12+vi04RICcW4S1+8Lz090LX13F73VD
Den9RJGYwaZ9j2Sgyr0Pb+uQTGsskRqJqJ9ZIcp3ZzetC8GOvY+Mtl7qS2S3SrriFbX8B/zuKaQZ
0eRFkltIKdMcurDxBrWS+k3dqk4/sKlhXElPrlnCPZcfEG0HdHLm5LljtCH3A1AuC9ASHm4mZBUQ
WZ89iyJeJk/MDxYl46xuNSwtRKJ5bUJRV8MuSj7eSCCNcVRTpftoeYxOqhT+RU/wMHczPc1reiB3
PdO/q9bAPjOs/fk9lokMNjUOLyPYtE29xyg7+/ZV1cgEf7bnuqa1wj66z7dopjAohMOxWZYNB3oq
P/IQ+KcMuKtSXOvfos/W5esM8aND3yfWZLpy7FfSzpYL0iYYG/rJRmRuAc2p1PIGI5qf+N/Wn96S
UB7dIFjfFU87Gcw7mdMOEwOzsZiuj2MAc/GCe0c7P8K+lHq/NzdxLncEL4CWok8rllceJHzABvwS
ux3UKr1xKyZmC2+9gyQsfKfauXQAPV7fMRt9Sq+7+xN3rrmdbVZJswNxTMvgqOcrGyMvbS4vWwKq
wFn4mo+5IzIBVEnZhkmHo4XHqzA3Rk29nZQnh0w3BJO+IXQoQUJOKUNcxyor2Kjl7SvOZWDyEWv3
/0P7jVt/lMWpSoktyUgT6U2zrlvd0qXPyfQg4K84R3bjAEU63+qA859G1hVXBjroj+6xihdxIZ9s
EteJZcJNP4yKzzKi6zLaLbYYOFImW7jvEznlPSMYy2N1RFBzfuWzhA491tQ9TaAzRo4caHxv6yAV
44HZD6S+hy8LmNbuGuevw04+HqQ4kRehcgC0cEsQDv0phcTGDJ15hYcCQRyO232F+98IFyN8YhrO
EaNVn2tlJJ24u0V49RO0382J9M4AiferxtVzK8lgLNGepM+MdrtOLUU+35BE0wN+2U49Kx6BwIaB
lWsXNxqRb4nySpys8jAT2umaA0fN9lz4SiCp+ZPVHubuv829IqpPaX1jpT9EHHr7Iti/pw5QIC50
MAFONHGjL2oMMO5T5rKYjBNZiCPDdGHxbHRm1r8Sm2Xct1iYdEt8JI4HCOXmX3vgIXAIzoCTKkeV
UfOvgxppn7by1Wz9ANDWInSK6wOwROTR53IerVH+7WSHCmCCfPExbwZXf3WNqE+KkWFGjq/6UFV7
Mwk4AkopLphlXH7Mx4MZt/IRoKfNLG+3ftrrVS+eZEkecxTHKJnMeOc7ZLVpFBhAc9ZYVzDmS5lm
m2d6Rs+dZv32KQqJr6+aOCHRo9Y8kEJ//ecesPYRYqZFZCSfAsJnpp6Os47qeYrPhdJ7EzuMwcHB
55nsqmXnRoVdF/BOLaYgSu4DmNcnCvPGdZAgdgyM/xfeRKOEnsf+gcPYYEwLGhEbHwjdx/J1vssn
t9JpKomkwHVyZgVSr2GLoPwAvj85y2yzR7fnzpaIgMQSGO3stt1BEXl2rbcQt+jmDdDkJfFxCw2f
Fme9cq/lA7pHrC+qjOxm3cEy8CrmyMjQe6cPHlSgmjxcHCFraacnDFmJRjYMi+chBbQq1nbc6vCi
diEd6eEyzKqJnBNhHyR6NPIwHbmkrkOF4P3KB1BTPHMQ8tCZ7beplbvUtDZ2OgwnM+ZP16JM4yZw
yhoyz6HdXYruGcrkZuAAfjSimU0B6Ji/A3sL+kdXFWRG9JebTz/b2wrnUu9pzQxTypu2kPMwYFAG
2YPY+JRlFvVf4VPoVs2dLOYv4JW5BZy/zHAOhMKts8k5htz51TFmkkPf0i2V2n9XcwGokAFqzryB
ukCvpvB5su3uzQulYiaDNr6zF0PST4ippGzeCb05C4b1kAmbtED09+c6ykCGgBTAbSiCeZUKthrT
ByJqyYpTQ3LDWb5v3FUh3AXUCh1CLsayMejtnMQ9xJLDZdGrQEHhO12m0ajtLbXH6r9W56yS0v54
cIAG+zR4TqRt6kToYWCgYLGZN1dBGSaECU0eltVNfDvx3DYG6b347ERbiUT+2j/tbkgYvP6NJxwG
1XhAB/XXjhCseHjitVxG5lFjwqttZLjU8m6Xxd/7n7zarbhTuKcrAH5E85COKClsR0V595pBK8T2
YknxLv9pOuAb1ZH7/Xl72nO2L+adHE5hNM2BTGiZc65x0vjUFvtFLvZpXwQaH64kxHuzyVRGpDGr
E2q8rgtqbNLW9ICj5mcmbnWcusssJ9LoQZbcw5e6JDSIjUwvb3s9lDNeFBKdel8a+m4hquSgp5GP
d1vvShw7PlsYkMbRsNWXgGTF9KnufysI4K7tR4KWopBXlhX3gdtKjvau0T0THgUjBilgZODLa0R/
IvjAaBFlltXjAbW+hog2LPMI4xd+DBhdoLddbk96LWOj80+ShWtMdhVAbraW9Z0BbZS0O2TDECXE
ht1WoXmb6faLYFCBZABRNyOkEE0QxJjEOBR1BOMSr4k9SXLatNhW1a9cjh8nKFp+LYzsTKlU6ASw
P5sfxJZSVD+aObQO6JXH4nmzP+Xn1eRisSjk5sfRGrZRkykMCiMl01LgI35bcrmb7YKVxJSjjyA0
rIzxFTplM4ERaIEZCiEzI2QN1nNEiha3bjLvnaDowr2pUqV2u5sRYSJ5TIJ5j0+TzjMbktKFzk6T
uuMZttJ593IQ3CvjuwBFmAzRlLpedyyAqW18sKcih4kcE8hjOXzDG5s0mved2TvEREmohzzNxGFO
Pt93bH8gflb3VF+EhQfdhjsssHTEokCHf0odJI6s3naOzvFeJ/8/A/Gz9LFjG+z/AqgXoz9jDiIr
b3BtWl64EIXGIXjw/4J/tciRlDY8pdgrPYOSfP72Wlqq+mG7YFoTDCvZ9mnnSPK3QbbyAOI1WCYg
HT31TMPK7n+GAd6Y7hhmBU0MtZbGUAcQEHwCw5EJ0Y6r/k/KHYLQaEUztSSoblkD4RqFAzS8O+eU
zPUa7mHtN3Y6+TC/8csMtcQGcZYQDrIBErqpOGra7fCxghOFCQ3u+/MfothZfJT0Kpzv4/7lQMeB
v3VhYFePPsb5vNNRcR7pyF1VJFA8NcQoy7i0oBLge0LeMFgPfItE32pYrSWMvA7lFjDazHL4tyyq
iimLvuBMdwx87HNV9zFkPSKezpuc38m3NMNUBYYdoCRT/hXlyETM2m6qqIa1cXtuCDnHclePe5JC
VXHN2FSPk9+j9hSP+JKeQYZCRSpqdRZfd1788ih3nspXOu34z5lfKwJT/qlEta43oynBnl6OIfBl
taqQQp7ldDzXF95oC0S+uEqrGgtVSOneCy7QQ+mKVVYNUEbFk788ei4JhPUIM85XfU6Zi2G+fdm5
g1C9h4pDVpuxz3ZGYdlfYnBmwg63WLzPnTnFbQifi97MYn7sNQfW2K6iceObrZzcWeZ+nbQSmxlU
1i8C0YYZKvXCf9TzRuZw/CEJumUJ6s3kJmLI7s6LunUQYDlZEd77M/MVBF2XZ9v8rAkESORyODLc
BtKrVIpD1UCcZ0T641bSuoYvMXNNxMDJDnqHjWwSGtqB5ndTMGf1KAnz9NSG7ovjxSO/BP/Nk7oU
7/v/fsZHeOJSM9Q2girMN61cp7FHVWRKVww6J5TgW9kCGEsxopl/5IPgK3ystLIe7Gy3qzaJpJAA
6QQQJ68grFutpJZy3MIybBHibcVX+zLbrfcUcUQnljhKHIKiDjJGb9n0hGDrn3N218bUSJCZfw41
wGaTt5Cf5YXOrqIcrlZ4iYxo42mdqAiHpRJCIbH0oLZBuRCdkCmArgrYYpfRqiFxZpjJcNNzopTd
aB+8AUAZM4/utK7A/KXZuZdTYQe3Ilob2+J7MQpz1cfJr+69DNDML/U3+2G2U/IoGrrFoRoPZ2xC
ON76da+EBLNUm78dazBSKYPDmMXzLuDTUTMo3xoIe7oq0jC0jN41DVHZCW+QxmdVOcGgHxnf/bUk
wdjmeMTjEgYUK5lUsA4NAyTNF3/RfMCcnnT7jJRQrZMe9GuxixXEvh+gn0leU4oV3xz6mUHu52Kc
UBWwoRum9NquKOJvQywm32mknXXCj+RDDGUlH+Ot1XoLCwCtmbwXM2EHUP7dIk+cyeKuQMFKEwUr
d1xi/w7b9bi6Xn/8egaXpqjKkHDvgx2xx36uHlRyIRdnHr8ze+X4yrCScDdYlQe95g4VLzFv7ThW
Fdi+VaKw0/QEHNEAaC62D3gF6fEve2v9d6+ik+1mcJigizWYDNyALruHYQ9b/q3NACiSInwBRDXw
LgEZQruK/2NQsKaGKRM+l6GE0FehDvpg6jzKSr1DYC6Z7/VoK5ob/MABuBOXzfDSnFYow51OC/0A
7lmVNCB8wmIwPnHyD1Pd5g2DDljn00pSZmrndIPil8fbYyRM8ADmMpKSbrmy4LMzvjbihLDSSbbC
DmgXCaMYncbcHY1CtNRUb9dgQTbYIfCAYUGmJzbRT4iNZ04SseDVPq+Fjn2sUfzlecLRPFr2MtOl
Fs7IM9KEwMSv9dmcewrvrRD37/Hk31bbQuEjtr9+T/JUWQNewrHlsZGXsJV0I+kDvc4GdjMbfl9L
8aTKQLGp1/DijWJP9FT/GYcwc5P+1UvW3iOcv6hZ1RkyV3vMra/PaKa2iDgpxXVusI29KAkWvA73
tp76PppqOMgNMbJw5831DFid1S3CtbNCExDK7I9XEgfNVIfTN1tjA4raFCH8rE1OxJExkUM2c90G
3u+OaBv/Oxbb6U88yXgTK68J74Z0WztGyWIDDVZPiD4OVXUSrV2aZkUCHZUPPIhXELxiEb3DOVDO
ER0um+Toy4KiqC9pYObiMbdN4ad0uQxe1RBhCchmbSR/Wz107pZKP2gxV18yAgWzIfxQ++jx6GAW
Zas446X4lCVeOgCmz70E0MN8WJKKBpjhqab/jTdvy6LtH7G7u0CjifSt3gAJDkq7ytqmEiLzLqZc
hRe8vYADFXvSIrRlDhHhgH55ueMcMpdbHvfybebOaLSP39utEeCxQFZWAS3Nt9165XNS1myam2ME
tbltDUrKFLoOu+3ThVSKUZXikOBCUtXhxqfHQ4CouwaAZzI4jTkWcTEW+2O1vWPkjCmudftCqCMg
u9BD91WtnGXEm4sLF9JqUls1VAQtFpnh8aAh3ZsjmFoPQ+tKKVWTGpHf7QJ8jFoCYM8AgcbyJKPq
AYtq0ynz/RSErBOtMUhLrB3jfzJgKCnpuJ+Sz0E2/DKoyBbzsV280UOcZnrADXNtaSBK1eieb3p/
RrEbi7eAlXENLFRlq3Lwe1vjlX+DJKUpYIETXXz4IykA9L8gOAVi6F0IYS+rmwWzgt1vsMaF2EdA
mBzhF7QyUkq7knAdobUbvnZHAUoTBTnWbNJFKJRhc/kHEvoVLZN1cDRpi6ntL/vD6Ks/X00673L6
MIAMXZ1aKnpoRZ6SxVrS8WZ6rO6GKE+VUSomjbZqOmvwgauS/ylCne5hbbO6NOJqRwheH/ADR0kO
7Wtg2KC1n78Clk16bxMMAvdgBs3QJvKHIlwVRHTRIfLEIUY34S4F0HGGuTESonlF2h0rbej+10BY
91K8YoijLTacaglIWEjyc5EBKfA5Pz0PGGkxFPfyw9UynfAxKtJZCN4Onu/Q61tBT5hF1s8/rcjX
l0v+82ALCmB2aBvYYpCHtvqJJOhIKLbSha1X2Atn3p5oe98pHD6lRQjEpulCZYjFqKqQRl7xhWYd
arCEhl1Ai6ZByy3G9XItlyAkvOd63P5I47+aN7izDdKARzfqSNWe9CgyHOge1721UMGVvi/AbUmz
/TxOlNTfq4/VRVf2iFajIZmqirSD5cOSLNpqMRzXjjeF1Y6u7NqGbtlbu9mIfgl3Krav68SqzFhv
XKPdVdjU6DV6tL6IRVEA4hp4lXLAJ3YO+U6RoxVBoeE/EhwQYd8UECy6rwXNX6aHwIpz63vtUso9
AgjLttTfcKLYmPFbWISMqey80PhRC38+002EdEu4npbmYWINY3J9ZJeaVwE+NACYwJgVBfz5B9WV
IUOzpvrifGJzkqKdqxHtUmBgVS/V8jCIPuhW0scfl1HOjaCGqrXk+1XrsMbeGo5taDuUJAhKmJI+
EZQ4EQznjrZwdSu1ipVRfxNncGs7KyZVlclO3cwR04ZZuKMdGc4A9AMswaaFVf7CZKy5AbVFQwBX
qc0mdLttqHedz+sz1ZO2sKpOvydYnN+DwL9/OpvTVb8Hg5DKAHvmvKCyCIx7bOpst9BFrdw36tYi
IZjizGdSCm2HAomFzJPjF2BjZ6LV0XS8SPGqg4YVUIA9hqj24tFY3ao7X3tZKR+UBNdMBCt1bNZf
7gZUKejV3B16me+z/MXApX4/bVEgAgwpGhxNvSDnAZyDwol+vmC6h1hVgaFw+deIp2faRO0yMJH1
Gbp6ncgIuaNCnAWWmCGBuFgOQ/WE9EuO3+B5k04t6VaZIgFeSMVh9LNJ6T7gF2Nwkmyrif/nHRkR
6tDizcm8jgo61kO4Cs5Hb0CURgc3gXOUtAB7BWQQYclq1bezt2l8booW+nNAZNCuwHE5EhOcM5y1
neLbn8JCXBVVsF3FVvmjkn1xrFrGP2fH2GRs0dmOdCmqRWi5+QV1Mkfra0/YwJAdgItq3TozOYsz
B5Xx4PsE6BxQelRs7UuPvxw2/DBsxM9NlTIStNhw3KttGfJAShI+ZTQOj2BZ2OF26VXkPbzCfwp6
Rd1FqfJCcBWTFZ9QD5fYgFzE7BPzh+vC0krTRwdDMughjdk389MvuMDxGHgSu0UMDnDco2UtAZxY
Go/9nn5piJlQgMqgk0IPlsV8g3k7z+K1AXZNncWneL49Eole2P2J7JdtXj+9HT09/rENc08nCDey
0LCFta1Zer7pfaOQWFP318j8EcTekZ9+3h16hWCOUMYiu2Gt407x0iX0sfMZTPMbTkmD8SxypN74
wDWBAzIIJYyTQGKCPkx+y5qeLhoTe6s7ssTJs9sFJ+LznAblAWALzPhysk4ZNeSHv77B1pQxqDMD
9IUNUDjHFb0lsm5Uiw/AQpUhGo+qqXHm+CRqafN3Pw3X7y+ji4fzyzu+lG/YsayrSXVvE3/zpAjM
PS/NH9ehViwOrwP7Z7H4w0JMmtjs7/+wCoIsWaF+pqn2O2GQKa9e+B1xIijQVJz7d+e7XTk/2fKf
ids4QHeSOeY1WPxccN4jsTBw5sIHvHErOLN9jVnpiGvvJ1TVrG1PKiN/42ytRih+2b816tfWSG+X
WbfRPDsZapHA8f5kGDRfTkW5J2Id1nFCwotwVW1DdWEDXQngQxuI17xgSonRYg1jW1ZcOb7ZvEe5
R2/GzRjcal3FKSIzNC6tMcC2+Nr/t34azoFnZ3mG/36bglCuSX+I+If0cTfUpoBvayGXajiso9PZ
f4UIKP7zWOiAbpzOQCB3y7zNBwo28nexRVNOKXE6+xpUHEH2gpiUZJ9+NsTNb/Q6RlMI2XIh2MS0
a4RQ8bvuG3/V6Klvuu2BXkt3YeaimWIs5ablP7FJfCwAhBLUK2yOMd8/WXd02F6yzI+LeBBKHtmy
J4s49kijRjlyKfHbHaIF7JVP/7ikAbDvaoDwmY5f2DYkwMOpfH3Vcf2qg5/qmPmMj+CnDtYwqAr3
/tFzNB7rp+xNUz5BU8Q1cWv/KRLYNpIlFcc6ZgS1qfSS4P/pGr2pweNENfIAob+y3n0FUX6YKIO7
AKwmy3HzRlTZkcsFzLuVX6N1IX+VG75Plxb7sq3JAUNrBDtF4b+8nmHAugRKRZRLlx2DqrdsNDAT
I9EllzG0ihxRl26Z7Cxyyx/OYLfnB23SVIK025lRBIJ9kAqZIhjEsoKV6nyvwrVn8/uFIdiJVPHE
gSP+wn8ynziTGC4kmGidiZbh64KcFOoEC9l6dcVjQrgyNeE1gBkfzKdic72uy36ZkmzaGDIN686V
L/Yy+/GIiAlR5gGNlvbHrpjydB9A2bv2+nt4M3N8d2JE6j5Z4vu6HGyRgE7t1dtDwhoj4ZIEhdqM
beugOkiycqak2unf0Zd+TNObIb4afH57wLe8Dh90KOWGo5uJd+lsFtpCGzysfD01mVZTVr/aL1hv
Rly6Y6KXhGcG6ffOXslft24Tncgk48Qn1QCzbpRmic3BM2vZ7Kx+lbyf5E7H2ZnyB7utGa+34nt8
k2PYacxb2CDvlY97zdtjPt6msV/14OmO5jFepwXU+JhIs23pGBuuqyBsalCtgQnt1J16HvRexSld
LUHNCeJ1GHp4RL6k7GZjGEWnmsFeiSurqrZXGWg+vrV+yqeiRrHdiGW8/RBszZUlfyZ9jYS7oCJK
08tPMimd4v6yX/swYoheXVOk57SDjVO5L3rb9XEaeQ0TYsyImisokVnGLY1TvQ9DOCGSi+aLZ7am
YjSLMAMDl+lVXigPcCVt33sUuhAS9ZQ4U0Ea6rhmyLy6Bq+oDRrCu15r3olFbCwAHTAiqCeo3Z1F
USGukSqe0ENRcBWEp7DcM7U6pZac1XgkYUvVbVWS1Q2AQgZuC48q55cc+a8DRCAGRz11hcPG/NIu
TkU5p7x0NPKNxv+aVYNMLLjOelhm8BZVhHDF4vb4NaNQLe85ambZOm+5mRAhsKGmF9uyYC7CcS3m
pNgMTuvuDYG3EAYKgnHKGGoIgaJo4s0TAMI7xHeT+b9KE3Kys0AyTd2dSeTZV3a/+fq0e3oFg8df
6010iVLXVrIuklUuUmBlJLmNifcz0Qx3R/71KhRAGkUWtr+E/yoqpH0YRENzQ/DU7EeSlW8OnMmP
a6RP4TdMd9GZy0IaBjW/Pa2Xmz1IkM1jE3sH+qBsYIf25Su3rX0rn9fWuY2J5n3VyxsaVNDqbMoj
7pQmxiZTEH8fPRglPNu7TAfFlv1qRr8m996rUZuQN+qjym9R7SbBIWdgbywrHXqkYEceuQcOPZfb
12YVkS08X8BToamxiJA/L0lAfdf98Rn64isLE+SmqX89kpOGRJFflUNXjPOxgt+dGglkLJmHyNhj
S60U1np2qyIrFGHHKBU8tFtZVGkzSY90lrKurdoRb4oLG/vB4liKrUTSQcq0hSrBiNU6Gm5O90or
41rUW4n0n8PcGWsI54I9iK5iAA7Ei3H1W/04r4SinAN/SRqhUB56bMPtxi8dnj7V4b3PKrvqZo/C
YXZAHr+FgooUX9HDUJ/bsV8yq8khKbs8LtXNs1wddYQAowmZ1gBBN+8DSr1EdehxIYWnYi599hBy
QrPrDtFjwg5CsYA74dvZZ1TQnXWgaTHj9GQLxQyCZgceXPap+9dlYXgmHvN36AVI86CO5nix4Rjr
eSpErxEGy1ySNvbTGe0+7H9QPXU8sa/hAp+zhnxMJ7cJIOxKVwgNYKna69Am77ycoqurBvIA11uV
W+MJE5QWhdpjL+1JLcoyhkGYsCFn1C2zVqc2tlVlPDoX09nLGjjzGr8tjY0JIn8xiWQHxreTvjIA
mtg5AC/vhYjAk6eMnkHQ+kqN0TatFW4Xa9IbrFYozr3QS6hdo8CRzVdT+p3UzkreaU1i44nRqxMQ
iDVAxBiMoZk8oqtdpTBdUAgTXCdRuxm9zK4p6k0XTC5OrE6QXsIqQovw7Nwn4qZo+X8ZQhbfOoez
t6RwZsQhzG0OvCsZi0tQUnMhwp3s//IXaFxJt5G995ZMxevtlhpz5sWRwaBoHxm/h9AOxsxkzANJ
PETYqDbliyA2kuvmg7Rep/+r2dpqpCVmlPA0eYFZqQtL52KVANjqYHZSxJqjXuC2oomBkpAcTrUE
/WlBoPGPeC4313rGVYpQ9yzITg2jY61vk+hRYJDciFMNsSpeip6g88Y21DRWMktuw54kIkJaQdoe
T7gLj05Loio6TPbYwo18umAKJ7yEoNXz+LNZbEIJyK3niR7nhu/n17b8EMTTHW2gFmkACNxIGPOl
Q1q1pQgj6FufLv+yfNMUq2bn4aejQ76BUqoa9V7fx+vnYMYJXG+2OyaDy/1keDduQNEDLvMdI8xn
J/sJdQkLEPrVwBgejSUN/8wAxLBWJolovZdrsTQlaYCz4UHnB1Esit2NNwAd/hlsbuQ0JlD8dKHo
84o6AWJ/TBp3x0bFiKMwoyx6bpkpPpiQVnvabxBs9GRbFKngj8Heh6WiCMH0sDoNDTCAk2s7Lg5F
p3YZxiOyUGL60JvYXO9WmoiP8dKcgX+XbCJKvCWsR/rMQ9wDeqX7nnoCzglR6pYFYy/c27BYscto
W4aSuczJxDpk/UOW1UlrEYO4PQ+Egj/PTkYWckYbLBLvpgDTlfqwJ/QszElMoruzp1QUMhgkFJLg
6CdOC6n+oQD3RXLQBM1yYaAVKz8x9qBnSdz6AK+x5RkiZ4IiXJ0WokhhqMvBg1oWBqpjyi/lT9II
OH7e4uxLEF0sXSESfHMtZsiXVds2l0D8IUaKLd9BtkIpAtPtbiiJoPzLeTZV/qnspT6u+jMfMgFo
r2fYeRgvjRnmwuUX19N9588D6Y1AGKOlcktQJG/HERbY1Hnc04aycSUKwfQlqpu6LCVLX9mZjXR0
UB/gkI4AZ1kmy9KxU5jTTSoKEvxKndvCW5vPvCJnBM6vM2X1rqXyFN3DAa8wki45o+xn5/xuoMLd
5S4Sauh44xSNyH+fiYDXNCDml7A1xBelad6yYA7xdorWIQL9t4xnfIL0808BWfj73pnPyRJnBh2c
bRlZhtD+gp4QQ7AAZOZHy+icGXaXyNt85We6HwWvGacnzNyrXyVbO/isnqFenwv8qrXXQfGSr9Uv
jH/e4U+s9JtY/ezMZkEZigaDvRfZPycv/rF0J5P0KBmcsFzhZ2WK9XT8ExVqb/dPDZBcI/4ThJbS
nB9CWKA9u+kqmk1QWjPCmEjfen2vNmOTau59mYvrYEQ+VQl7hX7HG9yJAeoXZA65yUoFm/vCX4jF
BmSodcGubw0ug1V38ClkZnsSJYrX2k20GeQBG7a/T6qGfiHMphu69k1MnOTcFkZMHYSLw5D+N+i+
5ZrLJHOaNfxOuA2INKjJ2ZnvrDzAcrcs1NEWG4mBdiR/xoUeoqGHzE0598W4Jes5fsMX7BuNbQ7c
IWGmjBVpXUK2lyzDdTEneX78cUhN3AtYhy7XwS73YZLLRRdWOMkrOW5k0ixirr2v7Eivqxml/6RJ
H0zWDpCLq00fYS171wyQZhCQC4L3H6JRhUARH+dX1Opv76OCYbzm8RSiDXdB9aynjOarSKkqZofs
YhbXLUm3aa5Kq0x5UQvhtm9HJ5yLwprGLV0RU4J6Xq5iu6nkwZ8/0hlNcJhV1+szSGc0bTejgeD7
r4mWjyzjw4jU/WVoF/RRDPyWHcUBofcXX8kZyFGbBUAVW5R5XpgZfHS8GAbJYQKd7zSswmbzCsr/
waAoiWDN7zbQA3/bjlCDYcPClT35O0t/5A8RiC62IxWAsgWt/7Zok9PaFkZfw1mQFYpK/iVkhk7C
pwB1SLRebBOzbdv7zpDfpN9aCTeF+HP/aWbs4C89wWLPkT+fHpAuqI2p8lhhieIW1RwnifpJTvV6
0OKi0rSJEuoxAPk6wqM9dkjoAfY3NhgYQntglrZ7D/zSieEc169F4oyYtFOcUthzdR3BNx+E6FMR
x0n8F9myYSmZwkc1SoX2/8KX/N18caK1ht/OHjYKr+MY5oLJvgKG5Rm+wQefF77/wLxNu+R1x70o
v7QBnmZWR04D2nZCLi0bNUI9dI0Rc2y5C2OQ4ADkta8HpdGKH0jCrqSrAInxm8P44Tc6XGfb+4jE
1KPJcad6dCGmxWOSbr4l6zSeOCEhqfm472J5VCce2rIBNIyaZCoMZecC8JP9+/i5f13FbMREtWqL
x51f6zvGXpNSx+gnU7arQceEB8zMpxNKlrUnZliLmNXjmhJNBBAur9MdH8Te0IAS2JbKaPCuuQVq
ds62GjV/nUY2DMAHfRZXqEMPIVGRhgiKTFlALpM8QkusSNOJCNFSwj6/yjd+VQPWy4zd+uZhhOtp
zWeHHP21Di5HRE+CV6ImhWCl73ZXUpPvDFJ4kbuSQLsiIulvr78GlNlnolfw140Su/10I5GRlEfS
ValRWjEZPBh1znz0aSZR9NUsHGsEwnB/B1pTF3fqr3m/7pXCvq9nySw/RZcbNE4dHOW/qbqSVrnt
s4Gcsl3gi9Kq/v4+c/hhfUj80GAPmOSV/Ryeu7wyBQzTqzfBMe1FJ78C0CFY38iFMHYDRLkAOfiG
xVbLjMnenrCPqPqp5STxv6Am0nVFYx7TAXzm15fgcSlZtyvu7U+9lwqJRvfUKyG9JPpejSKxc0c8
GIgQ1LDhVsyd57p5FGtGs6TJ4uRuaNNh6bhwpTOrSPgnR3kvP/VOh0KpbshKzAbCIQtXqSJW75YP
Td8vdJNAmVFqiMgQo8EHHZfy3g66I76r+FThZTzloJQAJ39NMCsTBMfzTi0ZM6ui9HSetnjxjE2x
xnTCJBIryA670MJHbevd7CBy2jvLZ18snkWpi6QTWfdZAZMQjkMLS7xqKjlI0KFAVF08/8JnG4KE
5dcOU4S4BPUNd/WuCqtxnPOItGOEieddrGoRMFyJcl7Rxf1d3hzKyK5+Ns/253KT+twWk/hvpT6o
jrsel1eoty4/g6/Luv6p5eSdyJL9vg6hOCU8HZ1mDyydNigTYuMmwW5jpzQTevtJczassx7fcXfF
xUrnTpSdv4jMwaSrTOnnO0mJ9Px87K9OUxtbQcTUV0fHvvWSFB323Kx32hOSu3mtjKW2v3gWzF3A
XxbZDfG/Eu9PxK5X967RPXHleDk6tUjFmQKiyewZ7eZipv659eYm2GY+MDhwpvW+wivD9k+PFwOy
UcTvNVv7VKT1QRTSmjDsBYEyy9a/gEWoq7jG90gYTdVjED+t+Qf7in348wdruQtKN6+AJptRgBWg
kxhfvOydZ53AMwCBXNnril8kyL936a8A06RTcxOQ5ngSOZG1vEVU44XM8O4U0kpemb0vWiHrEVFv
NE8WGLI7kwrJi0EoHMTSwhJOVs325KZJOo7PvoaVeQxP8AT0qOksesxc+TnNgHfnvXnfaIow063R
a9DMPN5bqAqOUFKbaD7FAQQ8BlGh30n58lINAbdNAFxIrTEW+HH3X6arkdbthawOnkdKJdYjLt6b
+Ghvr1eHTEP260zpq+mm32iwuVJUx1Ate9HrWybJ22cbXiyR1NR+No4O4V7IKTu2QTAXpXC8GYp9
j7CzPpanyW2hnOS38be9Owk/dwcsX0OM5NH+lANAZyS1Y36u4POfOWYr3JWkya4jaGRwHSz8lzkE
xGu7h/XX9VumasY3JXISQvm9iZ+iZ1vYtgpV886xM5jY70SoSD9ECAQHTkpD9gTfznD9D8bYKw04
+klMae07Ss2lXnmJXFRQ5V48auNmGL4lIVnE4BdclZotvGfFqw19rmVo/gMf01AtqPR//FiAVS0U
dqA2lFeD2d9nJcqWUOBc14CVvG1LaH07QczOcoEUmMntZimavZSHVI+6aDNUp6ti/Tc74op5BNgS
aqMebz/8VmMRWL2kJK/91mCLmjVkUD/ErO2w2M6BiiHmIlIXjolKt2CzZImDGQcfbuwtYpKLmUiF
q8i5EO+ogrOkz6F8pI1GcRmCAUzMnStk0Y0/Z5TrYqHdAENy4xVkRhbJOU1xycsPCg+/Y54zgD5F
T0K/4XnUnPpMGarF0oOj+zpz0TkL72HxRbeskOHwn3Ye/lehpxLfbLHkolcK8WSveg13cHhiwpMz
oTeU4SbcX5je8nfTvUMbnUymboGsAAJux6YUWQ4Y2ML7KFsDLtheHVsoyxrL0Zb7/HEIQ8zMEweu
ePSngBC+85iATeLxgB6CGAEYXI+x4bSWa0+Brq9LYKnBMShKdq3xRbdj4tqRo3ZItyBDb9SUXmex
gjhCNrX/0TMzDQ1VUPpTfX9sIiXOR7fKlKml5mR81svEyzJV/J2wMfr5AuBsswBUPWvDDl1Q8Idp
P74XDn51ReZ1Qpj6cbArfyfwokx4z4u30Ec2j/JC7RbDBjWb+XzkihUOLNXkiYwsUZfcYzqZRgfh
6gzXZo2ocdv6BIpAcHXA72qwpHkrK7llSos/d1utS4RST3YQDOIwQiyUVYS+QbFfMdx17belclmD
ZfhrU3YgsmQ21qSRIfDzryQzt9jqPQ8dg+0a1oTpBvx/Tajm7IS9DADpjCtdjUJqeu/TIMTBGxnM
EYg08OwAJbHmtm0ApNcU+yyew/JUmW3OU3h/x/WSkWt3qprW5NDbqAE3nq2iGnlBQWm7W0jua8dI
B9FVliYFeAdP+z9suOZ/lZe6ParFdj7w2BYMFblznYJLNS0SMVnGexmpjO9B12qznNxUZVRZw6NQ
MEg42Go30TBPEIq59uz7IZjGoEUXUqoD3eBkIUy/Qm2xfyNZyFPcipRrebpDXSQoECKb86QV4bsZ
dvEbwpTsKBb7OaIZDMfDddx3PLoEYRoYEMWFl8Hsidupi2xkJFgd6rZu2JGeU/kns4MiHxUluImZ
hQfFdSrRpBei7DA5gTE2GioIeizwgkWHg6XqK9QOA8v6x8I97LeBJXwe79M7mSr7bIx90z6q3lpQ
/25fAaBUC2ZfYgyNnRkrJw+8HxVQu7R1lAYWcohsOiEYh7qZeq5roEkyejsS3Q07di2MEpfPNEUL
7/CKMa8HsAOmEDjM0VPVI+2SGfU701cwe0VSBZrjN6HSjZTJzFhehKycVG/JGZtxKULkTknBBnaw
LmWVsNQXgH1O6NUVPWaOf6WWFLIOGKoWB3LJmB/YRj2CZzxa3JrEANFLCKG5Ktuw4FprPYx8d5HN
nJidKupF1MzOBsxvGf0SmTV7uOj97b32l6F+p1EsQM6DL89Bl/KXdgTonUNGztb+n9afT9PfBfD2
5kn6ZDysLWfxDsHo0E1mTOSkQZpdjhl/+1yr6AOLq+G8n26dpwQu+8bDLCMVSQolJyji8nmFGLcz
QiDFsdRCRtXbXEAYn6zdm3SMxUtQPxJ61Yp5gkRdkO4F2vqZ9vfdMwezl4CHygqGvS7MySrAhz7+
NG4TPGzui7k6oJ3e3GiUAIyF65EEbDLhfvETxf+ghKTqUdZuJEpcFbkD9KSJ2BI7xcWb7eT0pxlk
/w3hPzRY95wXeDMSICw/aOpBzbDnn0NJy5FHV6oMBPfI4sGGe/ozP4eUlx0qf+E1BLsQVrtcXLR5
0MtGg1tqsBNEDwRy2ARl1WZUMtcFTRSykVMJYSpuVABBgTaUYHNOEBimHckwsy0Rvz7/dV/7zZ7m
wiEsZT9gdaCeA8z35lv9FSWM4Y3ZhcUTvcfuCOJicu22vyPHyLrRAMQqiyFs9HhUpnvQ7wv9wCiT
5Kk6RMmUH+sziiU9xKrVzuQgqHU2N4FVZ0gMRl4V5wk+7wsxY1jOuWnrvc4FAtIxG9h3Zke9wVBD
NgWEQ+OOVBpsbIwgCb8yKzym2EAzdLiOtsiIa2hI1VQqsZkXFRr8xFNFBq4rKajep5Hv/QR7iLim
jszdx4fDQUso29EKMlHHvR9GyE1BABd3LFaLpoFXU2PR9ZL/KRo0pFQWA9ybC5l78sVek8sYUg0d
mMnBqg0yTMzJlBKnJLIl1orIT9FxzXVtqfX1FGcJLuzuw0FhGPU/9qILG3rQ+LMh++A69f4se4BP
wQYjpRqkw6g6Rwkwx7H3NhdAX+YvNR0rCZ5Q4RRs8wjhecIZA28uopfsy8Ds2YHZF117QvQo0U4Y
w+iCfcNsT0zgq09ZZdfUg2ECU8cCxokdmyReEdYKs06zZkK8gSiV/fe6+uEpsVfem3eFPmUhRucg
EqRAtsnYicon6ShjZDrk1rkHUKvJBBtFR9IceAo691zSBj+ZtkKvzlDGB8mto07vCMUBquoqyYtK
JHDVnZJYPFA9GeVfO+XGx2Bmibi3LypAkpYH+nYC82uvf9kf+N7Rp1iVi0qrsZ6zXFSBqAjPG3Zp
K4WtxGwua5T3zBv1ZgW9SOYA2+9cZFGLjcIQoN4ji2XjKulPTgWTx9RZOfiRuNY+9uXHL2hzKYZh
tHosBdzB+ekq//htLgqpoPpLr3b2bXLjl8NOl7jm+kSU8u6Oim3Wqno3EW6R6dpgl2eWlD3FaF7G
afuLJT5HtHMi0DCVqxjDMqFkMut/4GQGCR961jCJcup1ZTXbcwNneGNRB3tALNh48SwZL9+SrAKy
VaKQvpmNCvNL+Nm4++d9xlUXvHgZ8UFyIG1djmm4f42VSR0q/jvO1dR7hXzQ+8Q87k37leoDO5IA
5foXO6/GtGmLITuCIZM3YKel0yVaeH7MPfPIBxCA6KrmIveg3470Azl457DvVQliJfS+zJCwIlTu
e8mleno4+EL14ypKJl4lNm1pJJHHlx3XiL4T/4vomiAVZ3nZfFMWWx+Q3JyJrCKjStlAr+bISB1t
8J/6r9G0p2EL0TFkQe2cHVGyFrOaWtEm7O0C4I63ew2uzzP0iW4o6n3ZWrlckoglEqEZlF95FQ8L
kiQ0jPAZnCDk3Bwf+bDJ+tQkYtSPGYKZ4BT+S4QF3DFEgdhHv/b+ghoB3kGY80/esyaV+PzKHrVf
lDlz0fyb8xeHH0UXW6yn3LMMlr6Tg82I0RPKn3Ecju2iAINTyg8b5mau53ucv8PPrimSib2e2LUD
/9MSTs0Teeq0QytZ+rB2OLOOqIiPYPCDBYGuBae8HcrERmnrwVWjmPFcvIwSCobCwdPLZSb1Ucjc
QvcrhRSWo8YzK0dgMiAZ4HrZ6D9N3bhMyq4Un6mbHZMOBx+CacW1DP8RcmKBRKXMC36YFsCFxuZ3
4nMWm6U0b3oX+uuULwpggm93f+0iypSK+u4tMv4tWNwpqJ9lM9QcjVXfmAhAUeOTG1Kg36TX0IKG
c/9oVKu3DUQiASBm7zjB9G1muCdn3ntTWKv9bvemIGlIr0h2g255R+EejZPGepaElZZSxlrXBbCj
OBdGKt50glJTatXDlyUMrtVNa7SS7nzS90dL8bL0Si7GJZt4bWIDCFW/IysVNqB+e39DK8/a3na3
f89FfHj5yPZT2b4PScnquiWCZkbZy3X41+Pkp3i2c9vtYgsLms9QXm8aYZLYKy3NuRx7lqecLHEz
obd20nVGRX3Y4/+7/IOsvngIFmrtWIwnwGTflB8APmVKYxPUiWGILeN0PE+Pa8EXdwmW7z5Xpf49
laGEBK4IahqsALlhG1EXYlj2GBPcUpDi9Xc6tg+QK/SZ0wpxdEaJ3dS8agKiMWm3L+Ef06XPkkrx
u1HmvjmU5ZffLoI0I2QcCnEe9FdzjA6ukbnaitWCIRq99LXMdeeIX0Kppe9S8ql+SyN3S50y+EAk
yPr6ybqDeGtfgO2H5GdOYtTznCzXiG2qz9rLlNMBiCB+hV0aeoBP0Lhcg1ws1NZpKb3VxJPuvKU1
5luMem+gC8M9pEYZaef7zKyFZ8b40dq1psSW8Vu3iBkQI2UbDgkSdld7MtJX4PB6ljVsdsC+vnvg
oqcWrhzGB5TSiApGvtN+w+7IYtkfJGlbDy+HOrDQoCluNwdxm4eSYUj9D1HtClmVULHU6pGFK7xp
iP46OzfEuJ3xTCnLUq1h7rsDEFwLAKqyk7in7fO1KivfDevdYeEiMiRUcbCQANkwq6JwMxBYv/cr
6IgUKsncaTOPUfUZM7tTpEhwiJN1KOKHjOUUVUvDbAwr/QZh1q3m2zappVIDszzsXVKt0L7fj/6F
4MRdtMqm6BnMhNWspt3FaSOEX76PSTa9HFOy7HttL85liCOQaJs3NsHwx4hNjKAGyqbVRzm2t/84
mpxfGFJ51NzG1auYtCWpMRUWgJKceM7gV3mPGrzkN0mbRqKITWBFvUmm+pKmFrNAysmpgsX/Dqkn
MRscugMXQC8qUZ/E14rOzoxxdEiRHRpLn/CfLMPXajsK6Aq+F6Fhy36OcDpoDDMXd7LGCAKzEBgy
gyW9ERirb6F2RVwDTnXGy81afhN+KHvtJIqKlUp90B323Te9ltm6SQvITg0yvaQMGkUOn8dDWcsJ
27maqSXYVlTXnwsL4C6uv80agz4oG31M8b4avH7CM7bLIFBOmYO79Pa0XtgHH4saFvxswqgvl4Zz
UAS5Eh8GqDylfRiJZF4MsN4fwII33RPCkrUOkhJD2Kleu0pnLtvb7d7PMXQa/aiaGuytWAkkPj5r
nbTODlSbN4BLOBGq4aI0RLcORyUqVR8APNV66QjcXKopvJvGbiIgpp9Ekp3I4DS9UKvciKguyN7X
doBzaMX565IdFHPJrvrm1KpuAmugnaXE+b60qD491tWTKJO0zqhBS7FuzfnsfKr1iihaL4nK9rVs
QhzgbcoUO4xo8f2FfJfarzLYSTmXIRqTfF3ieqW739sy8EBrEo7T0X+LKHNyy4jyzkHetv9p4eK5
b4t3lxXKGRKr/wlsSjA2jPn9mLwC6VSU0kqrnImLYlfbcW9g4zWGs+hyofrI47lpmOyigjnL9GDj
r+J0Ltt6a5KhfTPODTSkr0ZaMpSjnc4IZcHTQmc1SnvS0dY8TeAbvE/bGxfr4d1irZJ2t17OJdOF
IEpjVgOlAcgL9LL4x7HVBYEho5iN8BGzcjBLxBqopkWPAMj5CTSA/LQwMjIqdVYwjCeDyc1NZcf6
dxCJQfy+OEHPNVPZBi9/EZhpodEuoGrgZDKA+bovCoNeHXiL77JBTS5m2TmTCVFhBtf6X5/iEiXW
eHnJscHn3/WvDJwoVuE7lp+0A4sRR3m5vqvUG45AopudMiF6H6SlH2s4DF9H2WHF2pK0qRpdJ3DX
8cDlGatSYiVsANM5du8f8HlKae0m6fTJz97EFzW5tiGHb5ZDm2MMI2OS7Rxr2rg9S43/4t/L5dcs
W771L+5Ig1hJA7OgO7TWjV6XOOMd/Ce8s8nYEmLuM24orKjC/+QJD0kOcU4i09Vy+ccufiHnVRTp
qG8pBg4toD8HdgThpEFdmsoS8af0NO+AxS7CYsoWyCfgouhSuaMJht7dZ3zUJchnBTHPLGEgHp0i
2SVkOKod7s4vPJ/KOYq+PRlXzl8X5M3WKae1CSCBgCcN9TOQ2E4kbyySWv1nVNByC7qPQuz0km7e
zRcjSq8dmYQ+W38EzNipH3uAsNI1hyEYid0ks1LNr9oVKvGNAIpaJmjYXfbYPol+1U8rTyJ8G6Hw
Gt7OeByEkPVPzT8+ElJxRd0iaYGCKNWlgBP71bbblayZ1ywu/rcycoRgiTJkMHyA/aREuwcIPgEN
IzYdLcSkGzMLkYkSqF7HI8nK/yIKf6IZ33rNSmW6/8ItPCWXdjYVJBNTX/fEjPfgHIlFCjnhqv0p
BzA8zNdISggeeWT0fUnkOUmOsTgXk9fG3KRGS/M4sA+9CkG6/+OIeX7ETTEUzn0p7hd/U6IlOt4C
rEZS4ftzr4Ptg0gEe2JNP27kUMod2cIGugHswNm56a2Hcid3tYa8f0Pm4jFLvehgO8a0RfmyVyYe
6PhJvXOb1OzenBHpC/x1w9H6y5SW5oR7nx8FU+8JT8MgHRJhpO5fK7kAC2bBgW8iP/EGRo8R1OQR
3hw44epzHQiC1asJQ5LKPmnOm4HcU8AT0pHkKkQi8Nk57iLI1hWPBfA2caUID1WyE8Ax+ZuLgCsI
xYbh3a2wFa4DSLLuZo8UdEg+NfRRQ7VbrOU+ZHG2mj4S6Vc1rfYb9xJEjVp11OztcT6qD3QT+BSt
CaKurLHez99/skf1gEF8q1YK0Y+MbPNiIxjbQd2Bs0cD131DSOjNgDSz76KFvdxqFw2kRKc1orp2
4BUw7Lrmk5PL1aZO/kJ6ag0wl0v1NMLB8vLx4YIyJcFP3kRse/PzAxDEbdVgzeVsrJumIffp5M2N
UrKlHdGnd8uYSx5MjELyHhSulGmlkOpmr73FwpB7OdNotTNLmYHSgE40iO1eytBhWhLUQpl/9yNp
6uThUmlen9eM5DDlVzkNkPf0Ztif6KeppYmmd4XaOFiQKAZAX6AuuTnpWCzWm8Z0lvpmgEJJLnJv
8EDYB1HOkE5hwtkPDxrfEMBbk57MZOJrJV1gk1OC5eZBCnfGS1J8V/1UZCVOFtGRoonuRi4NTStx
e1iVNj2Hkm3nog7NcNAEnSoRXKeL0EipwAM+R0vZA3TwPqCO0Okl3sQYlt4pJFanOiZYwYLNkYCS
IUOWj72nW2CUc1oDIZ+2Oei7ggV/Cf199uuld1ZOK4PIC+E4ivTS3VyhYWUdMTC6uVdmlFvq2XIU
l3q05ZwCC+3SwAcA0NPQHdL1zxlwA3vGfUAZwyrJmFPvtBZvaP+hGTHIpQXniK3kCzXzoUsrZTE8
+wnIr+oj1VAnLgwjpNTAUc83fIPdhl7v2x2VHMnj/Pr4bm8vOo/viT0tiZLt/GUvcWg4CFl7Y6Tv
EgsD5R+MyAs9t88X3Ym8kkDZdcMPCKVGEYojMbmYhRh2K1FrKgAA8JjbWF2HrIeCmWwK6VLuSwQT
uuxwbilyzu8vB6klfQ4LQ2Go+sQWRlZKO5slPI8lj0YfEBYg5lfJ2ROjcUfiPlZwbgwAJXVRbjYO
bxnUINz+NBU232wGrxPEENOTZ3rZihqjIZoz6N/Rtz7YfwrgqWzg+7M0jiQmGqPTSnuCLfyyUntG
6i3LfC+SmGlNznUqlqyt0SwILAIdG3no5ITOgkoG7LqZ9I/fSE1R1dSyf+rMvzsoSgTrfaZRYgZP
wLmLn/L3EUkwWLECTC7lZnuaoFnn/PvqH+vqHdXyvxmOBjgmftZv2DnniOYF5wjoQWpPL7GSF/eD
ByB9fCymt/+rPy38ezMEn0x1XxagZihgs7bbloPWbFX1npYpxQactYl3KAYY6lERLw/0zXElz4WO
NC3//RoEebN4mxIMTb7/atL4II6wea2H9A4/z4E2ygQFB7EhD2rNiISOiCTlKjF4MQIdiiPufiqA
krV19ttYtuMuwFiaH3blQPd8KdbDWnRrU5pHhNXuYUSkHHQaPcEvqVlPfOHs7KxCGM6WSb5cj489
MvamQ2aomEx1R5oxPDPNiBwj89uUGvILXRPiL9gOEdklNe+L5i27u8ppBaBqR8Rt13HN0WpD33b3
BLNIhBVxUPAiNRPwqu0wRLtCF/upy6irMoYFVWSx1Kyh2c+gCpLgYc9wMiEB5kbHWNKhxnUggR/u
Fu/Uicj4FoMUpoZwUQvFGX+3p/GNiAl8YRUyXBq88zQGJ8zhYRWgOwijN+nMZ+9kDdBYoWX1rP7y
+YUaeGi3wx5SDmYJyaalAzs/3uU++/I5nX3cBRPWNjLK8kGiQKVvzl2ukyeKE5cBwTdSCJfwORBS
6mZ6dnL9NmavmaCOX5BfApOIc1jrQa+vfZF33c95Tzn/
`pragma protect end_protected
