// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aOkHDIeuHdabtFqwCVGIJlFTA7ysIi7OwinedWWZbVAdGYBmXxF+uNzHLRvA8qpq
vm0U9kHME+jZekX1YpRKbfI6XNsUyj93THTO94jvsTssQkg2FvIy4mwwQHpEQCRI
wS4kS9bYky3Wefnu3VWcx6h8tdLn8h1t0jfAOGw+zbg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9424)
XYpwQQ1msj9NBbfejw6GMDeclK3+cfr4mZiePa5xY6cgTUSfA2wnxBhC8zsM6SMa
Ejsk0dLnK4mHJyglvcicTacNdBld6vk/G+ANiA8PpF/0vXim1YMvvqFDKU9zIUv0
81fP1Y00DHeeuTJoZjEneQUUOqTW31h7En0599icvNRzHqARo0V7XbGdD/pJYtS6
1jk3ZJZ7bliNO+GO2aBRkKz7O/RtVBRY9E10A/cSxfht3+luZzluoVHNqgBgvIOO
pM81om5vvN9DBBjGpYBq86n20d/PJgy/naJGPcpb2EpQ7FU+6CZ/2y2k1Y9Jmvpk
ysMzofabFA0LwFgf4+5wEyzBE9I7d02BNLSQURKC0y+F7TiI4la8y87vtEhSRHoz
pS5sIzJAnVH5iN1pSa2j2oxVpmc0QN76vslIPZbyiyJ7YSePgJ2KTo7eY8w8/sx5
bXLyVzvzumlK3MB+cPoL4UNdfapEIuX0lavFN19BdFjH9TxGyng4hKETjZg6DK6X
4ACSiHAsLH6dMjAySA19qi3LLGHdl/MOLewKGG2FB3XN7/giRbT56xTIZbcAwMWO
PAgf3/ype1pKSA4wBvKyXvloxdXQIQOg6TCHlA5c1WlVexLvyJZEG4znoWBJikAI
YSler7n45Q70FNin0jvVfTTVnpvXTJ8ZMI23tU963o6ybA1GvmuWcK/IX6VC404c
wYrqlwv8iV9b+v2h/qzlqawejpwaEzDPB9MZI47h0mV0r3N5mPGPCHrTnvlCK33M
Xj8aCIWdA5geqg5tliDU+tKI9F5I/XBRsDTGdvM21ShDDV2iLBnTTtUW/vPsFGtJ
9DAbdhio2YlNb9rgHB0iE+lPHMHDPMaS31Q0iWALvBnbL5AUOr4pjiVlDK4EEHTX
aZEY5iPVONvq6D0JA8OrX2lA53XEKx33VRCfxUxh7zWTQ79L7Myzph9Nd1vxOYx4
wJJ7EnlKyML/oEPCMIhkldXJRuqi0YSunQ/N3EaJZ/vBXFkyp5VNWo40dYMR5j0S
Oqg6LFrrCWnK8ykqGhG7UjO5aR0bkdxzaqr0j/0RFIod8rxWNEAZrI3maSMTZBHl
XxgvLRoSV7yBoXTQ8rUTdvZO6mCTm/GkeBCzKXgLzGMap1a2AIkq50+fkNmqrF4y
VMd173Y5r2ZTwAdYgMNqwYvmibZN3XgdlcuEPqa5uGyxMITVncSbzz486DjSrMKs
tnFej+l9X/7Sx5VWdiAu5hRYoep//FP63QTPcTTwkxqTkApvitKsKQlsUCr2OhX6
sC1k3mjOd/EdlSO7PL7o3ze7mFb2tQ7v9hjkKlyZ6oDECOFaheGGuZRikawa3kZU
Xdq5cNEUeX5uWYH1oHWyB/Qo3f/CHwIfSpVVHdZ+XcbZVpycwecz1KQMiVpt3iPm
Ub/frKVDZ3HhiXoPtjms0q8Wg3pKMi4pGHROqp8leJZT5uawTyVF+yWx8b+o779k
Yv0PHu3aEtxMYZgUjglJKjeR8L2J3nTj/dCDRp7H3dHNYpQezQ313jI3qILXHdk3
7eu4xn4vyWmYoss0O1kjIdg9odzUBhZdyAqCoDxxoX+9mdtzA5EyMsRQ9SWMEMRe
vIf1vXdh025WGpjHPrNlJUikJVrgVIiatvhdQu0O7BAkM4upYfByVuDR3Fx9oYwP
Zuis0HIO5R6KF5ZFT6izm9uCeuc2iybDvdUBK5uhB15Db4hQ0a3AsILj3oFNF5fz
6Jkf5nokiizJ3OciXxu8UgDivjAbgHFUzgnElRpE1xYukuahBw92IdQSoqRd6PDH
SiHNzqR/epjpmInY0aZQRkwVbYBvU/UJvUC5azq9J3CagaC6Hb/MjoJ47x1isGFG
bHUkqTBjZACx98488MRH6oe/Q+tgcBVBXGcrLOQhk5jDE01ij+1xfaLufV32wzEu
V+GGMwHsw7jYIieCK2rj/+b2IrkUh4K55Xdb44SvaDKp0nsoSxHzhNtmxZjNi7EA
qfmou/+cSHmFxw6gWtxCf8xAg7TMbGQlNi2PyZEryWphU6joWPs7jk0mb/ECLneE
fWvkONWirfjBge9uOlV4v7302X0YrhpEWxn8gW9dGUQq0ppxXWeNQNlLQ7ppz9xB
WqfwmkNokg7koO1JdQQKsq/VvqHXE4OPdeqGpCBm1+mZgdCAuLeswSRiuzJ6ZXQ8
nSBWhTx1hlF6Gof9c5NH3vWB6FxXBZUKAcHKqDVogJJmWEwDrUqXWvSJGDJ8oEch
KKpbqHPivn7W9oNf6sDX5VbccYaGRP746yW8Xdwre2m6ujEttj9daA7htdSbcDgc
RQqsJPs5W7ZyMPkAiXFeObHHMLt6kLVOBAytubSr4D3bN6m5MztHFYkIYjOWOvUF
dvKrKJjYuy/VBdhVPgYRh9IJ2trlHVdOoLxXhqTG5EYqju0Eh+BCGHRPfgA1zKlu
InYyTxcHOad6s0UVwf0FHRZkrS/X9msPsC/6lwJhLuXph4m+rPLs0kt9XfG1tH7o
U1TvPXVPvCEUIM8onW6ERlDP9Q3hhrqnqyZzjXsaTGuPth0T6Y3xQoV24zcK2gPq
pzpsCPw0a3UhzWRgBhy6NJNzAQoNHyk923DK1PZA2+qU2xiL4SuwUgRzb72PNtUp
2e5hjPlvzSBG4MlNW5snDyWTddjTwAYVPd5I1wqvOje/llfHS5lK714yHaMV0hrf
c1KAUiL4aJUEz9eSHqM8zmKm81A7MoM0AbedgyPIMvUKjWtrIEL3d9cqs/Y4LGX7
/NIluVw8biRHdEc30WbRyYVzTAY/cg+JcUihyjZehYnTdJlvMDm0TTjfEvGjmsJu
p+twlLEBvIRBqI7ir3kCPoSKEcNZIGOOFnmwvCvD9yyYihD786WwEHiPw2fsiSm3
AGUyLFjc+6ht5FmRQTTXIkC7rFZqvO1L9C3NDJ8HB1liTvnW6hDT85X/q5JkMav9
zUmqSUnCkKY1S5eccmWUtRrxzfRvGaLZaqbdiwZ6A8QrNTHfEdruzaTrjsc7YnXS
XuVKM5qSXtQ6yMhBd4ajtRnPYUPvvtNbgqSD89UXJs2XR+6GNX3gJt2oBDTyhpBI
mtPXteR9ZOLuyV0pkd5UISImgll/FBBzqzqvQsJqcH/fNiyiO8mSnGyY0vAjnotx
yHh3JOKxU2wGNKfFQjhvyQ2Q8Dbq/VP3KMxM63/VdMYDiNZh1wYpySI//9yt2Qpp
KwRn2mOD0V5Ix9B2KUASmQVANwprt7Tlyw856WmyBxfF5EOriRwjmgSi90Nrb+ah
cfvhtCVdgP0rqtyTlQlhCrFAwK2BpBNX8F88X4junCtYGL8kX5URY+K1edxLx979
ZZElnNTR+Zg+vpkeifeGkrqAqo78paHze+cIdpGVmpH8IOfwGzFRZMFyZ7KjcTwt
Lv5LLOTRo8cs1Q6sTsyXc7aUeTX3bhbP0JslX7IT4ff4qqJPHdb/KaBKPZ6J9a95
GJw/wOBAikBNQPhl+VTQUXxYxRbDMVwPNbXrg4ZGvsvcjC5JuSa7Hm0vpPrMk6eh
qYCp0GsK7979TLJ4YA1QKaJun3vAIdEdQDD69e+jiJt3NtkL8M09aqnx5z+7a683
tDdpbC/XaHXDMY7R4tR7IeDrStaqkS3UjqguSun+qjnXzSQrv7mt2bwaKT2rV+H+
JVejUTGuwx1S4HQNWCSugOIx9J3jFynrf+xojCNY0UAfFX8GjTDPCXhU3IDmu/M8
xRjmcmPo96jzqH8oSjsHgG4K5d44etCTZpw0O/eNNhvU1o1kWNoYaRxZHinK3zuV
Dr06ejlyr8ja4kXqb1XfuC3uGjgFMpiiLU1zITET4/lweycdqJGZ8WmLC3lr1aZk
h8it7jhdlllgDacmosH8lUESIf5xxYTXQSMVU9p4DxcVabbm9jXKNSGDcLsh+luJ
tKBwrtl4kvPhHX+VZY9Sw79G7AX36xETh5HhhnPMpyZwrfm/AltBO6hRRsRzOqk/
rAuCHIbS2tRXIZfkdl+WzjTS8XNOIiaKU0cX2YRBifp7hsIe6vkfwNoSnOS73qYF
4QC8VSY79oBWMM/zG5qqC6W/notay3ExNeN3Kv8RDbcJJVTuoEFH1x04YRiCNFuM
OKqcV8TlnTZwn7kXdi68V6qFFvyAh5AoxftSIbETQge9znIZq7Z51RH/YButg9kG
RFkBYcsMaqvUW2w7O1wHAI/iMbAgK0zPCBMOieArhWp2HEGJ0jFgFGdlK/Eh8qEx
cvxnxGZNK75uShnsRvSKGiV1DczjY3ZgcgjHgFZdadztIvq3HA7NyGNzdlcX2WP5
X03J3pKmcfRe3+Rv2E5Rc4ZZkn5hHgjdq5xVAtNGpgglcj1us7xIub+sZNoi53yy
AoEVMaHr/Ojgzm7Xql6OCOH0CWlgFXPlzCQs+1uqs2n8Eb1QGDt+shKD5heRwGSm
dxD7pRbF4+/6elLzCtIQWGthq3IWUaCO0+cxcFi7OzG1+eZIcg6GslTtU9zw6Grx
nvOl9BTzJ7UBmLzjBD+jx+alLD9Z0rFZsaV3fjMex2NMxJLTmamaMZ2spO4YGsQb
6gGwAVhREUs62r1wD0aqWB1oE+rp95fsZF33Ip4jSqO5/Eg7eTDvIiFT89QocEaL
94aHmF4XDrra2QSn3fKsXEZVd1Q001giXCcDu91Uc7CcougVjpqQnNuBmuT5u9l1
1fFlkf1wpmIb/GmBlD3oYlzpww25Nlc0suQi86L5S5h26Iq8gvx9g9dbG3nj6Rik
2xrvl/0VI9EAfK+wkFIxYAPLVxNJpHc9LrbF2WeXfakyqqVJwCGeEFO47MAm4fhN
xMRUXoZiCrUm4pjwX0GYrTtutQfuwzEfwSMonkTDpUdfAD3n7KBgfO9RasjIlm/x
IlAT04tqd9Ajmlh2YjnCa/04KbyZVHG+yy8a5i2lS60o7kAFMD1/aLonmk8K3pCE
+aYpv4QHa3g1MIbHDxQj5AViEhwh86emQsOIhraG4mggdk27VGzYBTfwWBQtaltb
MAUPSj3GRKJyTM1G2t3h2Y9TA4ScYgTcG5YPL4TvUk0PRmDMMzBbLtKrVti507Nb
xd2mZAzzVZBqrdCBS7w36hMG77/gSqdraJ8pjMj40Q5mPPjmm0fJSg+S/X3nyPrG
ZtJXV+Dc1H/+3WQWtCUgRhfBAcM/HrCzhJvlTvSsZnsRFOJ6vFXfujkobEZRaREM
HYiYU7MH2bvfbkVYY6gB19nMyWJfyXhRX9RT26/VZLYKCXsm1C9/G5Bq4owdRFN1
AKO1dgdXZ5YhVdTz55i+J02SHNio0BA7pZv5lq8VB6ZK5eRKkumxjNXGYurpeRry
2yZMUfYVGW3NzrpdgFhQRjMdiuial0mZVCubRYImoeLxt1DxfZKoAkQMskKt6fLn
2v7gpZhIwHYQW/F5h3oSbtpEmmOCDT/putmZtLb6xc/xe3IKqlbwPAEA1xkQuDp/
GVRqFxMMevRhtNR8qfxWvCychPaHO3us7m2peEBtqzHfN5iFiiN8qmGkEOGeE1iF
CYV5RjJ5twuEoLTNQEBz+ROld/5U2f2gxZkTsMq/8Y9wOuCvcf4QGNeutJKCt7bK
s4L437ZVpLkqeWP7nfbcmVvxudFOTgiPal5TQbmdrSVulbfNg95IBB4ChGRsS8Ns
4XaTimakYAmbxG1NW5UqiZiMeMf6v5EXaIL/so1nAwcemI/RK3IOicQnMhoMD85e
SPjiQv3WDegjPi3B7zI+w0nGIEp6Wrxux9p9jZI/nhVul2RQl2ESqCvBasgRSZ3m
PgoymTkanAplgZH6Ci2S9r1PY2okn90J5pAVN8UKF/WhePneAKWgx66xg8oXY/JT
WSkqHJ0WeNclxZTfjhheWLzpLkS7cPzKXauQ+i08w40H0aBEHbxsgPZBMMK8FZJG
N70CTkHvevl3bZt0Ht6S35u73yAXMc/KvuRotJFYMZ2/qHo9M19oGp22ccxFj8Vq
TzTooxquZHgI/Nm0Of02CqCPAaM4FLq3mhpysEuwzv0m+8cGjNF3Z4RvMqW82GgK
aNTDICaIea8+UPu2lQ2Hw2GXKnyFQn1UEOHuJ6/cb78zx4sAg9udR23a1e7d54/R
3mWMI/7CD1gZ16WE1qTgqfA3LoOWDW7DIM0bk/2MbZoDHZopubQhHiHuHRvqpMnT
4ULMMwasEdTLvWgNvN+UG91Q5M92sJDrPqyzQ3IXK5GGA5w/FiNII+ovvjP15TkC
kAvWyv1gb6luzC0SBgoGIrmasn1e+F4NL3ACZF7ALlkitvFajn3g3uU6JwHAhgyv
nBprcC96jTndjRRIaNEa8zLH1ZC4EBNMHjDwK54Ja5Yq4f0W8r3gp5nZRW7ABPoz
Kfjxa35Thkm9DEjQZ67SsOUnRLrmu21/KzTRbzBOolyH44StlIGYCP9+AkDR5gkC
W0B7HtqJRO44zqh/auFvqoiOJPJV/IF0YuOIL6tdztA8lvxmL1BOn1ndT+KCNmuS
nnCEmnHeuRGt2vSiMccv/dYiHWWwc3zKUxj5a6Q6WX4g9K+YH6ycPtNgIiOuyW2Q
WN/JCr3Qxw9b6qoKD42R8RRYVQyMlM/l/UN/n4q9mAAze0JhGqz6Zy+5gMps6g75
wboXFoigjyFAGeUg50eAFKvgtGusAMYTezEey17KiibU13ousLL80xwJpBTDYutJ
gFCCrMGnYf+15JREknhEhY6YI45H0wxnt8wIWXgRazVXJQNapFj/swrGG2nvkUTS
pXpKfC/h1G8P9/qriSOW8WbGA2GpTJOryYjLi/qNCP+rgcVdxNsuJ1xY83epNfA/
R4gdGE+5pFcGDmqXK9I4CcDP9GaybgLmXNntCNbO/mFaSXuIt4mC/OUW8q4d5Ujy
FW0TOPUJwQ/H7yrUPWC/24cf+KUnCvvNiXm5WWafBjFtoYsFLAZNAebHsC6veDi3
U7nYRCLiCrvDG7eWHWxNm+GYrHSKYC3O3absffysC64GyOt7CIoKZ+IXicR+Lmt+
a5LsBB18ljP3Fu1bGYcrLBxqoY17NBQEV7tHbTz/6H9mOstmB6Cuer5JvXYZ8M3t
UV4+6WL8eITTERHTvc2qCoFBnTU+KD1fUglm2/V5nseVD2skJRg2fBdYqvCw3kfn
y3VUr/bUEXSXo14wqm6cE6VfsmWn31kKqdednxXx70WmpFjBcWub8RiGWBbSQOJL
PxCxNeHNil4C4FC075VLfptVchwqrjaSqL2rvYSVhSTaEBxhE1CsC/NuWiAZ/1O8
QlJ65DOTvIbvphYaEPkTTpLb7OfEIWVKh5USkCFdOlmbPHQtoFcUOBhY61h5nQ5f
0bXNrhfPV78Wezn65A3LSdyfDBKEfv8q7Mzd+Wb4eA3cjqfVXujIG97oMwPy6+9v
2CYv9Xwh4PkN9PvAvbotG+w7xnXmHRw3RSCiWGmkQescbr1atxbY6yxWRgAUIXXi
Tv5oJ2Io2QN/gqy5mwOwHHCSMTK+0Go+7/iUxj52i5sM6ujG/S4qrlKxjKs5AQTS
h1JoAsaWmWkwYmDD1zM5A/9SfDEbjh2fslc5joL6qs33lVq6ul5EsCdo24NLO/X1
Fi0BNWW/Hu9XXuW0uKxqx/fVwTvG9R9RtoEz/ZaBrdMPETjySuClzujBmJXy++y6
Ek9GLwxhdHPoZT0TKKF+4pru1CGQNBKTzmbrRf8z2d8b6AdunLXg8suTdMX2L24I
Uwl/F6e8Vy+48embfg345Lk9HQX8+GRge6CnQRQk44x39lE//d4iC/8A6klfSVyc
CsXn5sOA7UdPFayt5vz9MhnhM9XvHl0TNqbQsGF6chfLk6Y4WAb+W2Tx//K7PAAo
BUUQELXwLL8H+AGndNiseOyiPLO4XqmKGT6oVkzXrmId4hYjKAG2/Jp9keib9s5H
mTph8dP1H2wyDw6DuoEPb1Ec7cSFIol8s88Iu/U/SZWJ4QW5pZ+dEA2c27oDasrH
qYanyQb+sd57xgC6/IWSd4zGZfcQ6ev/OBiMGayl5lNrWBw8vSZk+4GHCQP5gfsa
YJ4DjR1zjssIzdCAaBg0id/qWlS8/OkgXfDcYLPE5WYGPYvgh8PJWgpwpG7DhTQs
x+xQTXuSXXFcYVXJ6lxmKi/SQqizn4Qlo9wHV06N+KowjfHf6F+l1U0pPLMNdEOh
rqzHoflxZFU7s+mpJylw/HNkOxSTYoZKCpMss94PoLM4SD4rUJTir6mt9Sjaitz5
YteXM4sCtnGFJhZc2atGxtHoGQckP6WR2rvjWmhhMs0w5NFZ5oJ/HATYtOUztvAC
f7ZsC3xS8Z9TNmDAN8NxSW3QRcA83/SSE9QhOvV+G3CvHChx3K2HKweDeO/K2IZG
DP9W1kuX5bXpW+lKvN9hhRKK1UrlXUnJ8h8EY4L2OjKm8Dh7NonkX4olihXdy2Xo
UUeR3WGNo2MX7vyFlP0OcaMbWc3nSFYPK1EIEobB1fJig6+gVEVktEDZNZVCQ+f1
OtUniozhBiFLU+1neWdFHJ9/CDJalHDMREKN9w8siUwHTgCdvE+GrTtzFStds4We
w3lHfPjtoI3Gq+vkGr0zCwLUheRsxsBeXcSJWTIwdMQAhp2aWdgizuLcFaY9xcaw
E1vczCRUQJZyIlwyVMn2c8U/7PPd36XGzoTU7lggM9c760MnsCRd953cDUuYjotF
WA2juP1yFxIm/6nZGP5uAjbBsWwdytR0BfQ6QBGBjdF7Zxz9kwrC9JxNbyHvhqaw
HaGD2XxBquTCWeWBYcv8UX3w59ihF/ed7M0CZ9HZaj8ZB2JMvEYc/oSZR9t2pqqP
J6SPPHtgy4L5YdCYLDWZYQrLvKVBo5H1Fg29LC/RHcUzEXMuxrHPKrPqTmp69zjs
NvBHudJCUlj6f7DLuS7+b+Ulj2bojH9VCkFML/9ycqPpddUMpnk0pzgzRwGOyUQ6
V5/YkEr7U9wZytMrGSL3Ns+U4NzO9VT/QLI2ISn8fEAaFEQR9Im0jhGYi9HAMG4F
OV6CxFDFPVhixYtR5ra0DCzdEVA+kC36n3WJuyRE9qDB505zorle/gUGoI/mk0pb
RKdht+bRW42HloPc3g2tH36UkPEtXr+ktw18wq3kmJ4ghFEZk4Nlu5xA/4Hpw4kt
vSoeJgjjca47KvcpPYv35/pmtKF2L9KIA/OP/8hcOco3wY0bLfUzNN8EgZbj7xP7
x580MKY1iknTKw30PYkkw79FSLyT5tOfypVwRBr3kYV3W0Ks7B9Ef0SgIYwrgkLz
uPbdtyaLmdWeeOF0jV+WFLIJVL9d4njLzXgbOe48K93/MVqNKr86Fl5DNJIsLM1o
NigQBVlnbY1JziDW5nRBfIyf/9poHD7DtOThBqB4SoSy5CWN9XcMmw3u0ttPJ6bu
RJU7XzqOOPFE7ZclLomztT/Qyt72uWW+ySw5xL7QE7j0gwQS2eShT5WNHHNsqvLS
s5WXFUyvV8KyWCsfnRvs8yonkCNVobyoWsDiQ0q5/8WxCQ/MIoeE8GIrTmrPBtl6
Ez8K9bfWHZCOUxJTWD0Q8FJVJf+gD90BucHqjU86Q0z6kRHA3pPw3KK4j/uUhCDc
eTSTnEhAo/53RyLFccV53LZL3mZthjoVpKBss1qe2fQVUYTkXqIsBeJOsuYCLtEn
pNYt3dj3r1IsuFXiOCCCv41Vg1TAgUYdMRtUA1JlEP4QoDpWeAmCyJNLGO8oIl7w
pBXwk9jriFSwkFV0SKg5P6uJZ2bF8sJPd51LX3wkPZyNhvJKQTifdzE1lu05F3Kn
VmU0IKVk0JMmmvw8ijaSA3fVA9TsUqtrrWPuUNw4iDNiUpBA2Rs9NF/8hafgd9eB
sOx3jXYT9deTyKExtlWqTtlyUhyp+tlxmrmk8RQl6FUsSZijeLzNiPLoQwAVHbjz
76OIl6QbK7n2XWPkMQpE6FVWVYt6ZqDtNiIKqHwMLldlIWH6G/alCF+9AHDrD0J5
l9Jci05SNyjJxK2IWRQul70Hn7hpw17/UF6BtpE251uqYAxU8wbLJTuwcyDvy9e7
NJlLCdA0grXZ7QJAeZHOsQLY+VlfHLmaSRqk6W1V7JDnQnu6xLkHKMbp5vqHTAbB
DSk+rfZ3jDoWpTMQZuj+x1bc1LKgHBnq7eDBSbkHW7iye1ua4Lr47uiGXIZ9IFsT
5m2JS7qh88yZW+LTIZNgQ+4va/naN34tLBIuVz7mSwLYQzlgPdGK22yeMeq2caRP
/EqirXdbXgUizIOaQtABkzOab6FFUGIk84b0BX3SZT+3OSb8Iv/YyuD1LDJUGaZa
+l4+IMaavhV6MHmHGInDpGGCyplk8+GPTouKY06805Jnabixdds4eZyhtqNAMBg4
pHnwNe1pc8ftvxNBlEVCmaIFp+Vf7sAb2mGwf9I5atgrMtb+11AXIy6cbe5QTzUp
VyUUKadTXJUDrvNXXMShj67em2+GEkDV2t/M/aemXOfqWM758QeRb3UHWKmspuZU
kOC8P06uoUAQq7nRr/nVvFvNNzPjcDd0EzixCaTWXn0BTouCIPhOs/yUBKkEQoOw
tPRBxA/slQxHp4hoEyviEWJR6V+4hdgHd8rF+1HrhR3/ydjKbJM5EUeEN58WT2qo
Qsph9Qq6LB+2EQmUieVzla/lmO1biqj98fkUGS/a7iCXLEIgfdIH1+xQZvav6HEG
HLdgkg801p2nvIV+1OXyDHkqwf6t+tiKiX1MOpiYNKHT0LUZgFPBBRHQJ3xFLT6B
0IeiscbBfoCnWnBK8Ax5GdBhp84HJEGCJd/VsN6WXgWaVQOTBPjLTn/sZJk3dkGc
IzLzcIB6Mnxdbw1rm/TXnJG1UETP9+bbAlBtYG96RTulG21ZVHKKIzK1afeedWgt
OIxJQvzsTnAYzQjT/hcEdvNc3svE/i/4zn3/sELjYC0vSAMTS3SKXZeJNFooHHzC
CkgyOL07AgGHAWHJHrmGP4ZvdswKPZc9aLnBbeJjxjSsehd5RU/LwgXHeW6ZVZOj
1JuAvnhSfTJk9UzSpHLg5Sxpt/ohPuLQtucP8sDz3rYDusck5mOrrerxIf61hXxc
P0lvlAEmHtQ+MWEIL3NtYXSnO5iZyXxADm7IDPbPcTvdQfs6R6zNQpqYODuvNzG2
rnRPkUuw48yz9MZHDPnIy6/2/+LSRnIGxpLTKKNqxyYD8gKP22Su6xDETgA/X7ju
exVtIlatumeoZg1sYIhHfu9IGHbtoxHej5A60vC7RZRI/n6464JlqChpsy/Hd23W
LKAFjseUmLZnwIZIMed+8IK3nG6jFxvpXVWMqriyIdiouqvhYVWUYE7kQZs4bN6b
SPp+l504cQTc+LuGDZtcaDGEcr47lPH/HSuZz5MlOODu3GsmCm79lnIzKu1pjsoI
RF3jbCKcUWQYyGRk2wOBzESOo73M267sH885Fl5kF7cIJ126TTBbWOmbQ3KYwKRd
Q89eKxiCYPDDIgPBfhjA8OMxd9DB7QD9CvnlVhfAEWges7Jrov8nMha4CrS/39d5
fZ9eRElGT8TiOppqp6CpJ5xwX2/gmn879O7d0qU8pI11DZvWcWTVcuP0cIUrHJYz
zJ+f/4H6wjiNmxCaquO1e7IXaqCeqUW4q+XBhyCScn5Desto7YmE1J4ZKyV2Yy/R
AFociTxMidoawDHs+t/hdapzGp/atfjgs1ed5E8+Ow0V+jOFgGU/OCaLelwMs35K
nZpmVR1zP4WII7vGTZ5i7yM35nrCA3gWKYv96g5yLoAEST3f5EHwH36IJQgAzlwA
zsH2HeIRitXyO291e0BFwaaTaHSwoD0+ZJ6cIdRDL089gV05iXceAbQq9HO9zKye
KJdMSHkxXWv75peuZJOeREtCyE0AqwMxT/nvy1u6DqkF6OniAEhVFL3sRkyNBMfH
KzCsUGslN/6mj7cRSwMuOT6bLrivsoQT2ngVp1aLS51s7ST8jFxkWow1Q+sVFHoo
GVtOreUMjEa1KjsHH6kJiS3aftRYvFqOMnq7QkL68LobP0QYeFRjFjXUaL7IxTbU
dmm8FTDpQSO4Ai8woX8zEVeJ0fjv4otnwQCEVdtKXhncUtyCbRq3aRAPKoWNVpcL
wH6yNJhyzx9M3P1FfW9V51NEOF6vmHypISPtXfEEmDr9m2vcZPYqbU+JOcsB/0mz
Ty7wR3n6gZqClvrhftmK/dcP1EJjZ992I5GRI/HZUzPgLFrkC6lKn63KVVoeaKBI
PlGRakFClDjGSTqKDswbCFqhCaZbIb2oFDMwI6RGBoRB3JTUhzXIymiHxb+SzCBU
hzl3WJDWF/rKifJrFZUHNqmrA+Kkj9IYwjFe95Wynd9pxRZ44m+p75TjUBJWTa8F
6snp6KEX/rsgJ3OcvCqZaM1h4rFmk9BcMSEMjjZV+xGhAMyCeM/bL7W4Qei4tqB/
H8bw02Brd+csi0B8APmuwH6KvPYD8z/hXKNrZAJ9zMZaovp5EnXkthWw0P1fF5Kz
x3V4L7n5aPxHu0bO40PTHjicgm7MiLqAxC8LwMPRuWTJXrnWLm660Z2MU5gRBbNp
bv09WTN4rFWBOz8QC71tUk78H38qGRcOUOqGHQ8OqE/v0d5PyXT01m3rtAv5BIMO
TOwngSxjNMvdoC8oaqv6NA==
`pragma protect end_protected
