// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YsNfSdgPtK0E1m2UTCo9Tfm+zOz7EVLZ4knacTFGJDl2/RRUh6Jt7cI/Z063+I8h
NssL2Q8ZWRasV2+IktodBgoO2I7vTX8ylY/W7ZvK2EsqPpQqmUfux+i2bnqhK7Y2
LqddBDDk+NKzJamHOKbUwDip4MEiViUPd5w4CzhapF0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19648)
NgWDtlekYHSXR1VGQg9SHRFVIKX7NEK++ysi1wZE307BMwFvXCg//3fTaL0T9FKr
Hhmv+tYhqknf/WY/xfEDWIjk8Lh0ZXbRiEenJ+V0uhDGF1Zo2+9g4Bm41IgjWOIy
NJWQhEZijZY7E8/CiagR1gla0mNR/ko9VKJu2dMXjSAaKN2EkE99k4cLRYZvMufP
VI/TdQxYgauizrxjJddNbmnGKQR9vNrhNeAgeIbZV3i2wKi8JVHnjPcvM97tppRF
uK4qd4xVhsaiK/454yCMTaWrOw12gF0nYIEgA3PKx8fKhSDYmTnx6uNOahm2qt28
foNcYBXnQusaGOt6ffY+bczahpTg+225QcwqXfeMb6JttHRMflYIygVFwAZzWWuq
gHraXjrsFX2/fDC/wUM5WlGiAArLZS60HosNCHDIn8ARHMxebkDm74va9lhmeSLY
kFZ0OLdjXKb5XPej+tlV4S6bbBgKmoIVk5UQMYRD7O1keDUuxEdgYlJ8wHmHnxUI
W8/x23Vj1tBO2JJij8tMBmI/d8zKTLCXX/1ThxXvMlTmhSkNtdtqr9KGgjVPXHrp
8NHsM+qixvvJOcKt79Zq93DT50QgLefz86ZWlv4AXYqGxHiLm/8Txtrf918QiIa1
7QWHrDntKsYAI0fTkq+zLH8gi4JVbw5x66/e0r8eJFotB08mw5WKMnOP2hA9Vi9W
Obctbv81KSCaZVqCA+gbpqFHV+66coldrrMIgczVKRu7iLGuREAOMEz++5yPHriW
kv9ALKISWAyIA+Y7ZCa54UbQT4GIDWwFeQ8o+woJL0FRPDkpPecO671z5idTfzog
Xvc8CDh9cjUWG+PdtvaWuXhToDI9+6Ehhbgi+OmDQ4OeVhNsdYsJs4VM72NOI8jt
ZCrHalMN+7EO1eWUB5fsaoG2jmJNnuS6BJxx6DQXiho9hJHpFC+ThpvZH2PQD4jJ
gLzyp9Il/bBtzocNWT6jgKtIjyMLvRv+AEABJ+LILTpciNV3KAvo0yqwy4gAS5+S
Ud6wcxvq1oaOPmGz8aquZzmbGhn/kRUC2jAU7EHysl6lMbZIxtGpzrJPGSiz/L9t
3817Cy79AHuREM+IpXZfZ+FX1Zbug9zfD863sDc3IVmfnmf51BtI49Z4XNPeEDDj
EPQqN6J1jw78bAqfkbxizvmTQfFUYQxdJ5CIUsc8X25JWotBxrZGsfUc84Zyq8uc
rR/y4Yk/ZBeyeac4WImfGSvXop1R6RRIzbzwjrvelNI/38N5W5DEUblTiA2bHeSq
7zweoMGaWRvFsJJJnZmhwT1rtbWPyTFBm/PuxBuDbjiyabnP2RpO5kFs3ocEJUfA
jBdwuWR8dj7hNQB6B/sqRfwQfNvS17v9CkeNyZz71nPUgfFjjBLeXT3k2/XZhFFo
p0L/2bbMsvFuZQz5ZMrOzpHS0LvwtKkfisROCrtpbzYRId+hhmFUEs/XzpbuRkS5
mu06IFgG2MEJTL83qltOei+5j4ODgT3tExt8DHZB316OA2gzfr7ANQM4XlW8ojza
jgJr35xPCpyXt6e8SHfVaCyiIi9Es/VgwAIk0qIywcB5xXGub/lwV1VEO9LWxne2
q201Q+zMO6Ul1RUYjfA677Cqt0RWBiZc9xTnl79g2vvWBlq6v/I5nHQOoBcGBgc8
5OUteYsS3NmwYSr0SNiiUT8J7HhBcTAqW+QFlOidJxIc3ydT10hxKIUKtc9/o+J/
Scvp2h+GiGaplN/d5WKYjlZJh3xVSZtP1kj4DEm2clnwB0TunQJRozFyCuVRrR/X
S6osJZizqHA37UmCQGF2HtLcpQXMJYx52VPFtUsFbD3tS6z/7v/r07l192lKP9sS
wjentN9U7/IS/rFpH1XyouyqHQbH35KR+XvM/fNLvB27s+zmZbKUB+cee3PqdsOv
do+vZOvi1qGM2Kq9rSYb3s+Q2wnt7NLrQhhFN5Yhu1q2q/FeA/0SBc6XCV0zZqAE
QoaaHmEh1viJ1fSLJQZjLyhZlN42B5cXGlRr+HC9dxAqqUeyQCgfFpPDIRdLFNxT
sQeW3OuXeBm8Emxs3GaoWuQkcHNawbLDCSyTgp6cDkfFZZFVpTl0kUk/6l2w5sih
qz1E3wfFBiMlsmQExH7TC6b09Z2KQ701Q6ev0+YurBdar+12/i2kAV/nwVIVvuh3
R+/O/Iq2xvclEe/SqUra3dA+biVx+MlsuSTf0Yg4FhCgGnM/87fazAb3axsUD+dB
yNyTW6gmC4muGZmHv3oLTjr/1WffJcq6Lifv5vwhtEtpydSp8ViqeM+0BNjwS6OE
fPIIVyY5mhc0c6/MG2n5DswCnRPFQ6ZsgNLgp/kYfbbtF0gRphdEVdh30F4vGrha
pMCHV0oQoSBpvEd4B+Xprdradzw2DJnA4DrSlO/8eMcr9VrTDh48cxi572/4yYDm
1PqMNh2XAf8sySxGz2UkWxnFnb2EpsqYXL2g9MwUDr9jUAHwHGYMc8K2rugQxnWy
qLlM2GJ/J1PPDk3PaiDY3te2VFzcZj45za+AvBRt+/UgTgyZVc9JcvP1f6OlTCzo
1gHsYb/EuqgwWVPnOFefxgsUHlU12qgzxftK5ijG2KmtG2ESN8SP62qkvckyGBmU
BnMAnAstetO9XCxNKm41BJZHG067csbpE7g1usKjJkEZVJzDgf8EDS8cRosDw7XK
X45N0aGSGL4LeBBhHFDFwngC3zhDdy/bPxgrhhpNHs9lVXCpEKgPYcaR1Nxy6gGE
zoGQdD14Lf0WdK5YlJbYX2fPeZqEuui3yJX6nWKktNfIAybC/cMrjeneH0bS++LJ
CjEUoDyjEqvIhzEdoRTLh9wbGGuMY0g7+irlEAux55OFMuHFPFNAZWbV5QO9lMLb
fXJDHHKCdWpta16hSVSWzbRSoIbE+DsZPkBWhLbESOuhIM3w4IrgJEIFeLT98ZvJ
dx7X9Thu792Q3Hpr/pLOd14APRzku036GFXNRJCAZ3VSaljEXgHeDDjToPtOXsl9
NZj9uIl77Fp5WQRCYafqouTEdR9QPjESoMggzTMPAv/IQQuM4uUnjph7V/hs7ici
g9sZWecW/zOy4sxgtHXP3GRgX/n2gfgRY9+FQnIi51z80rjSPfbdFbAANpEA4KRO
9hSFOuSZuqcp5wYLhthFSu+n6gICJ7Yqi/6RkM3pTh0xCY7GUddvQdcCw4DVWapM
82MrAuPWxq4GZ0BEO9KAKX8cl8UXrt31v9dtztqC1F7bjsLY4kZujiAmMiZb1EYo
9p4TvLOoT8V8cHrCS00ggow3yNylgWQSGn7sH0Lxr4o+rciexeq2jZIcE8ZEM5IC
IGyjcBR2GzbxwlAeyz1dabohFhM+aExRsUWgI9kS9UOoiDkmTXB8pcdpE51BWXfI
bQm8ffStImT30cq/Q8NeMivBYWKYWkrqDXGUbDqbN9qT0CrdicFFOaLlJEENA83T
VG9/HRlJbccXZHQsJGAkDg7KZZO81UwYppSI4M3fvRB8fgSgYICH6djA83MngoZl
NAWQKQTrv9qhtyk1ZRIyTfEz1KIFOU2e77ebONfFcnckBYXcFI0fFDDok0u0nO0C
WNxtPtCS8BBbniAHR1BGWT8Ek//LVhVOU0YB5QmwHtmwbxla3B46O4iH5920Umky
zR2eOqlyPtAnRZCR+FvC59krVf/vmunbK2FlabNU+3DS0xTEUPDyCOudhGqE3cCB
5hAnHXB5x91SoZX5+KWN69JV2ddmvKFIYFRcYQsrr4l23StcuUHAC4/2mGh4RsOm
7utftsI1lC+zSJIYSbAtxrCRnAtXzAYFSpjL4OGUr1QLRwMdx+8K3VcQRHyOQh4u
IMKMsSz3fl0I0qgFjkivg205rYZ8S6lkvTPU3oJYSF4N8W3kbF0vKb0Yth3ajM5g
mz+RyoZpt5yTCpYPxxkLThLcqSysPoecXm5qg/oQLsmsYjfevI81cFyaanA1VIWb
jJ5NFSxHx/TQOiUzIGYLp5/LDYCXLB9ubqfcYFgu48nnavqQnj5T0iSdLhxDZzsj
4Mw1gdtH9XdShS9EtlKxFWnRZGSdUEi4bFxuL/dIw4SCWdfTM9lDiNjAzHi0ZF8F
+Jy3hr4NltNHldttz/40NcA5pH1VMcAUcrr7OMay4vrDtOJrFWboe6SIDJ5aySSu
UPZ6exebyvmKPs4z1LpRUeOA9pLfMpKSPhZHNUkgae3UoK4b1U7aZAM6nmWDwF7X
3Bn0dKBH2ZnqIxqEuUR8/9y3UWFOUuln6XC8Ll8O2hjdbsGTLcCuQYVn763vLVJo
/eEQadXuYOYJkkYHLtN92ZRAdBr6htxWJb5uTt9PeGs2FmzyPcL1H24m3awM34me
JByv0S71/mNSUddHa+jA70JUT2dh2GP4VeFt2jh1U6dXhlTPYWJodZpwfsFXidcW
KV778EHPKEXda96wbGSnWjqed9Kfsd/RWuZx7CRWLUWD+hBzICO79GT72467HTYo
oMk+fK+QuZhv+q+3jitQrpEePk2zVtto7LdM1LSDVKc+kVkJCVTmlEHQKmbT0N4c
1e3j+dX41VTqOvhN6/u4cWR8+ct5UqNsEuT02tgQ+W/eyO9tgrQIY4/K8SbDOKH9
gvknGG9xL5wl/mr0wxAmtHYsF50+aEblazz83zpfotENpr9xMr+MpYEx6KQcfMN+
7s0DaARbTJJcRXiPkL8yTHZ+JmF01F9n8H+JrIliQM6FE0UkKH10otYHIAxR9Z1s
v10i52xoQEJJVz9aaQce3T4+hQtDG6xBjcdIRMRnkELmRScaZG2hZSjCpBdiSSx/
4trFYeYdeG6ngoEFRHYVZ0/jRxnK3oVZb52BCZwB5ChMm/L7utDkirRwT2dsuinT
tCj8JIhuU6jrst4VtnQfvX1NhZ2PyjuCKPyfGLgOl5Ab2OQMxqiKoWgiJDvjGPQ5
Rx0grCOq+N9omLJaWVPUuuiBY76ybE50bhlG3HDCaFa6H68O9RuhyYqyptshS1KP
RDQk4WvpTJobOws2JZIaBuSa7Ad0Tj8+zAFprN8vXKHmFh5ueM0Tl2cEvPaG+CFu
gUWSwwnMidLrumtyVXZ5xB3wc3THCd1zVBTBPn7c6h/LTyHuMLx6+C8edg67LPzW
QemH412VdhuFOzbajBtKobbyZsljZM5dYqOasCHpRjGjGfL91tz6JqajYcTdm/9p
ys704hOxBIQcQy5fV5/9XPGonM+NuOWU38wuEYKrKNyR7UNXWlNo29gbbiCYmTv7
Wp6KtVvJG68469Z03AOse8xQaA7ahXaA+vVY7uZrd3DGFd4MmP/YImMDmomzJSEN
6/Omrlxq4ol6OvQbp0MWt2s+o8IoTSG2ZU4lAfgjZ8l8na+aagjVvqGrNAPl2KgQ
kJaqbYnYt8yskAOPXjoboXV2Y5Srzgl52kfRjeL7byaMLJUCE9GTTZ1Dw/QooXq0
pZDagB1bS3vjc8LtNFYlRw47+jxumJiu8kM8cndGfmkPx1OmLoMVEcEcbupZUqYy
8YwVqKDYKzYSVTfUV+LANeByjzyU0vox1wfGKXO1ijRZYbRC1v08lAOZdlJWdpUM
1XxWtEbBgxRlDcuC+NdmEZAvIXPiFwKwVdkz75+FPIV/KMUWcq0skagszpOEuopd
O7HpsaqMuBab25LDN+84hXSCPB6OWDhyKMYOveOUAYHy3RzBRw1an4R8wjhU7X8F
wQfnHpffacfBVQfsA/BPzAZezcbClIsBVBIHtapAdTkWaadqcnyXP6EabtO0AtUK
PSU3rWnqmZvNtJ1GLkLq2JhkFr6cZNsUEgQWbD0sBz0/s5ret5CAFv7lwi6rTKpb
7N2yXHmmTcHxwegcMRrbZle9QYhw0ysHd+XYxBORUQ+0VuUmbmW1R+vpSOpq4wAW
6bC7XHDuVEX7ZGMIHBZzopKzZ05jGo/T4effMGmQwez8SOAXP9++gGoHJcnuEakb
SD00umECN+uUhYGq7sw16Z+dTVLpu/GTh5rs3rehA8Dn+xi32h/GbU08+zvp4Y5f
ANDrWbVuXio6qru5nKggOzGM8cPS1jzfXPHaxqBhz+3jP4LTTS6w7ooKdIihtJC1
ZUNS0ACeUogC+SqQ0G6n/hnzgzelsRsMPVsM/vUGIvNDCXVHmFHkbnHM8PkbdOTZ
DS9TXc5n4zU7geEvN01sV8LffCkKG8yro+BdiDJa58S32ypOuD5W/UWHmarZVpEC
agIxBYy/2fyHPpoepghV4C/saVlEd19DzcySIdLPI1Zqfy5ToisedodHDcNi0IYz
gz/qyOS7s1duX1dyNqD5tXhDcyEhrDUCrr6TdC5n192axGeWCliMtvv5BSo9P+Ws
yqxBXVX1VCe8b8rRtrSmUDr2CVmccHOailGDmESNpcuQ+IO9fo300aJTADwuHABP
eoD06FXw8vFeyB/2LsRhBHHQ9SMJ9vSzRK27wHGYlYpIZ2wNZ+OzdKfBJ12UT3RE
WXQ/NQU9Q1q7UIfinHZLE2kyweGd8ieNktpAWU72MPo4Ci/ZmA+CgJEftu+m2siy
AyBIO/iiRzZxXveEVwa7Lkzpu0eGFjB/6C/eJTsm3zV5Zk47bLYnbMMUnXl7dh3B
S1TPnQ/CotO4q3K1q+wZlpaqFzdOYH1tFj+mRkNs7YpeezgQSaV4i4E3ij5bhGhP
9eNz0qVmp5I9/jBdc4vXVA6eTCec4cwRdlsttTNztQPF3i1czPvk4NLloqmlNegF
w4rh4lDiwEdXhkZ+MtS4x5DtnHovPjUDbNr63N20a+fk+Ks4sh12/7ILlvO1I7Go
umAJkZOmQiQrwJAVnSpbpD+zBnGN6DYXF8A0SUyOI4M8YXA4ldlNOKhXkp57BDtG
nhQxDtb+10tNU8mxGwmsu5jeW21YBZ4Pvlfs2cOMPhFt/dJ+QKOYGBG7msugohcg
7DNL4EDze5+y35F0TByk71KqgJ1Bhm7CIO2KOpDBPDNBrKsXQVSQbVVeKOrqugS/
reRc+lm/cuoR6e2KuaOdZigWk9RPwZPPtUv3giahqXusJUHG/LQS7PHMhwzwz1Lk
8zINvMOCHejABbqYqBL6pOKg/dYyAdun53tRZgLTOuH5EnFr07MiqajlYethbIua
51pjA95ZoorZjfi+HnW8EHbfux5tlyItFJk/38eZegySRXx2MEPos7lkKkfNJutj
wQRsFZWd5cWZVffPZXjn+IoD3EOUeA78/NRqlaMBQIQQeFpruvZW9aFAv7oYDhWq
0K4QALoM1NQQHQJFXZhKb6I++s47fuO6CuW2AwaKyVh3xo/Jlm4SyQb3TMDyAGHO
ifvjVXS6kskksdbjxtWVW3Qz50PDBJMkFsrUGsRrnykaTUlz3yxJAn3ALgENriU2
H90I2zpKt9nqIxEOLWwsf3cZZ/F9rKbMO2ba97wUa0IETsB/zYnorMofCbD0eZRA
uym8cvk4tigY7+NyI0motfiPYp5rojlv3JZ65QgUBAmqPKyxma8P+Ce7DwnVh5Gv
+CZ5pQU3IIbnoSS6PacF4hw36f6eGvThHpGlM1I4vGLsYhQT8MJbive7bFAUo3EE
NvbNqUPM0xLOVS7VCAhjJEmg8dz2Qy01ZVb6tfojv2v7Vyi8OT7/O0lxAkR6Cy7x
WeDqP84GNQZ7XjLSXJoKQtkI5LU4l6rRwML8tBzf1VaB8SuawHrTEzSZpiNx0Iel
Uhq3iATnQm1+4Wxnfq1kY3RUYkfRkcX07sQiJWtOI0uxag5uFmI1ZmKUm3UrjX9H
DHOwcmrGdigM8niWAFo6kJ5Pw/PhjFl03s543D+QWs9zvy0huQg+4KFnJz1jC7W7
sRo4tjlCkIsu20pvxejkbi45p3T1g/4Upkq5s37j9Qcnqi+Z4VCt5+F0ASERf91i
e7zCECLHOr1yTu4Dj8DcNIK1vDgdzYBDZ/4XcoXDP2u3HaI/sPFLwo51OOX50Udc
NlKihRILq8K9jo1T6R9zfwvKDFo+hhIaeTAhQaIXvWER33n0wEhJrom80hdEIH7R
JCPXv9KE1pD3Xoj0EDlTWGdomqsxjEaWOOtUp6A9NSlDPKKK/E2xeqriPHzwPUlj
C7Cf0LfHLhvRHTka/4Qte78Ts02Feunc3WU+kLNvQpuHvpTq6OOoIHOq8DmwDe40
XQrnahbueTXx59tZqHwcDroE0+gUVzqA5tDzEi9bpxB+p8iPbgcXhuKoS7Ka0LHJ
S9z3jPxg529cHkvipoFAw4m36n8zod1+eikeGe9vNXRj4w5BhpS0VXOfcrqzzxDw
pp/wnZJJKb4GTHnZQWDWuq0SYweoBUtOD7JHvcOdQddd5Z3cjtLQpBN37fg7wXj0
pkjJ/guNA5C9N2F1okfB3Sr5Gu9bKZPmtj+qWh5xgJ2aGo2X3BLgnh3hxnqmQlOm
/wVAg6OgsisXb5PEeIclaKm+agrg8hV0Yz/WpJNS7K7zp0txYjQqvH5Y3BvS5DKy
a9aOrd6MjgdaSoWI/5qs4Qb+14ccam96hRLd9CQMfn7dwkDzoF7QHXCFf66vg1bF
EH5Da6+l7V5ow+RRpP5+paizvuoIZbdn/ooOTtN8ctBGQ6FCE5Hs4aAzzj0bgS+d
p/rj+bD2LLVMuH1XvJmz+STlKSkS4O1IXhK2nbfzSIw4/cxv3Me14bpA5BSlUpoN
5HUDHNQb0/HyzFRO/Hn06kSIgfDvY4LkxQk8gpsSKoHCoozw4rmzPRdDEY8AtS6p
I6T7S7uo0hcPzqHZ/QmtMyLGOUDepRyFn4TxjrE3lhHtptL2Br7ZN+vyv2EIrz+u
FWFbSEMvHU/r7KTOxhVTUJ6v8ANnFONLpX6j7WuV41crYz5p9CDz/u4h3fmsVBL2
NFCX9fVGxsOIrFkrrlbWzMid0rEA5sVG/IPsGmxoSuKpGssMO1M9vUDIYLiD7s1N
yerJOXEvUU+tpM2lfu90E/rLRxvT/uf6hPWir/JEjjYAqkKbsXoW29NXiDEnPq8t
z6Np0iKXwHbYciDIZ5/jGmAk72auABQFsfST1oTGlg9B1Uy9XrLBT1xG0lScGp/w
MFN3dJ6Cx8YyJdORfDME+++w+7Kwww5MkrKrPBI7618BlEUftYavEdeV6J3fTc8k
uyAN2u/iUoI/EsdBGWdBkInsKIK25VO75jLIz116k9jdSSffxYyk4pMOFNnZB3+L
Fi/LO2xaiSAT8ITKFmhjRvEgDEXWyf72UUtVHbZKY7urT+i7nyB+HlAFvkYR5sQl
n3/FxGPblYcPtbFs6vSywW7oU2pyCQ55C2qBLcAajTkRA6biJ7x0jCToA2dhKgdG
z/43jSZpMeA6UXPEJMUt/ITA63NmsmlWG8ZoCQzQPOTZ9XnhJuqNcGXBqsOSwbeD
LqMZ5NyMxFyPFDow2Ov7gPkHuWRWh8Uy/KDT1Q2w9SQS7HpD9F3easXG1yH3ZEXc
ULcz0FdeetDGe8d6BfMGaCL1tfWWTyic4L3EbF/YQi2iijiVbIoN6g913AutLvdK
PWVJE7WUhpHEyoTo1C7VC8mjnrZwtYhj2tadSWeSkk0tSzRzQq1gjMp21+EAPIVD
Gwc6jXX3BPeHhAKXpWX1s7mjYotft/zVH8WkIKJv+XpLs6nNAe91QnCMhOCWcdKs
B2VaqFqX5KaqVJQfpKu8yCQSD+xuMmJ08yVdpJaZhncCtVOgPGEiHIv4hesRbSIP
PLyEot3vUIYKLAFUuhGC/v8fyjlqbpI73r9XiaCrCgE4ImpR1HcDxbrtzHC8BEj5
Nt+7JihNwQ4RuTsTtB0nELbLv8Hp2CZnb+4SSKVW7w4o7a8z0SfDvItr22E77Dmr
GHy3LBAe0Gno/LfPdMlzx+idNzH6ZYvZxg7chKjF/eo8Ua9q9GkBEYaQItq7+SPk
sU8N8HoEVVPyX1TZAxHRGzT+ZUuwF16LEUXPPSYRAPGi3AK/wI4IYGt3EDbILOj5
zlV50ucOy7kS9tH0hO58WCe7EN0IykQFbGfc3HInmd0ZNRzPQQH1uWGt4Ln8VAuI
znDhoUvXI2rVZ9bcz7B8kqA0icX7CqGgR7NwP8jsZY8kP4c1FX+/i+qaOQ22GBjZ
kaUup7MHF3RBdkd7Lb1wLba/XLf86j39HQxWN4VvxJxiVzTKO32gjqxMrrRkWZhj
knioblr8uCZ5NYbhWWHEiSf+00C8Yd53ZQwWpeF2q4pRfvYmIg2PpJULJBqSWYvv
OlaDGNa5pGjlF1Xz59tDwfdXC5baP0rhcAEc+Sc6gV2RTOUQtkTVZYucgq6uuT43
iNUfiq0R0GYCP5aAEviYc6Tox3phHWEi3cWt9OP1AXFtTtJ1dMwbJepG82RjK/t9
1DgPqwTfPVTZ/lj3twrqohCy/cCpvc4W1LJQai3WdkY61AjpHewrZ260alAZxk7c
Qyn5hw6Icwk/i6Xk5+rCrrzOrhZjT1WsuBREWGxfLXjnWjoQceQd3+6BvLFpfhVE
YQSQMWtHAs9yxV3mwbbsRAFKEJVqYbivoZPBsnwerwelH1V8EjZMFn2Q1Skh80s+
wq7400g/cM1WeRszuZ7cVSgKagnH6znv06yKKImxzADTpPw/bGQ7QZldVqBpZKz+
ndb5DrbQfko2BvJhYsiUY23s7++z2803kpagu33KgI2BqpNiu1gUTtVQ4IVvc5Cp
p9uNePc3M87kinDJW+Qb/jkN7xxnz4AxFj2NOfhg3qKZh/L6zJSnPZybw87BvGUt
mUroMMspTsQ+Ei2WthM3KTMkBsvY2XttNpeTBmHqJekwchInK8K10Fwr5PQz8cY3
9HXOtR7MuythrAKfIU6H0gSBkj1JOGkQ3wPS43d6/kM6jJtiRdPucZhQ0RzXd+l3
6fN9d9RzNGWYhRXkvsfiRG1dp8/Fz0HAX1LEsOqs2xKr3WLMDpa4uaNnIvSRgJYg
L6Ab8o/fCqm3tOor7pAThAFiJf5Lg2tZLLN300lXg+tIaeoXc2UJnU/aNqFTqMwo
UbG3e5Jappht6eoqxQuQos0b93Zn4KpqLHN+CYFrOuHBdL1LQ/1PQVb+dbueYG7w
1cEMwjFNdisCV/LzrcWgzu+K/wlhyG0EycF538BHi5YS3pu8TGUGDPNYk10w80XM
TaS3Cc1F0UiMmz0voql+RBdG3/Wx4Emjp1JRYMOnnNIuH6fxvt32jiOxQTylZLxm
RuS8WP5ZgKOpmCYY8O23w1XVHj68soJgEO3l5kevZQiYKYZqqBgVAENLVzxa27pZ
tsIAfZykP3TFzPcbcUzvu6K6m8v90oxdGBkWcja0Ycj8rR6QBSOetBsMlFIxIAPm
LglAnG2K0MuqD7nSuBVSzsqEW/nd9ApKrPzm0i8dRzDJ/1PoMqk+2XPLFfJmQLIx
w9/P/GhNiQY9p0gaohPLEfrHB/3S/jhRNcr+HSp58QBiaiOhNOpV0EtZgVQ/naWW
iU5qdiXEVTrWYqcXrmCUGQmSqXrrjuz33Empu46Z/sA3rXUh4UYRB+7UN21N+o/8
jRWceHLuPW84nc9VmnkkPJgkDBCH79LSeohCm6uXro/PbTcHcPo1hpF89WPcLiZt
JyZy3o6NvTk13zaJ8q8cFkHSmWC7P/METixZLw/0TVLE4zcjec5mjTWh08afL4xZ
4qqNcPVB0RRX//bO3WijJTQaQuuS0S0CALKFGd4PQbwM4h30/4RsUVHP5ZsE4c+x
AiJYGMCshqX+KYHnWqS7F6Ww7Nl6l1vP+e/Ep5Wh/4djP1hQycRc0Chjw2YPbvPQ
YHrtnXYhQV18Kozl1yv7u/a4eTvw7Kn2yQRFk33cf3o/Nn2kGFTe/0BvgHxTaL4Y
E6BOnclK5n//8xgllXX2OvZINdTmfWuxVEX6wNnDz+ABOUqo/w4y7XSoNUwPIXcZ
Fqg7uwS0D13CnR/42UhXg8pyiYfNrIWLlJ41nU6jGuWyzZI1mgnUQztRmDwH7zN5
RnhIiJnOY/lzigJcPAChnycfBr+y4Jx35UsbbEghLQS49w0nxQKTqViGcAiDaHY4
+bdHFM6C78ny0SUMzg1Dh+wzVjPSreCkBcRwZQkY2ZpAt2Tze7zvqoTIf5qUgh4z
8u8ek5zxG+UGFhgswPfnHmJYginJmxzTJ08GrhEVwVAR85gg/gejCQ5n3s0kyEzc
laTV9ykPKvOKnGca3echXtx6kX2EwMMytus8HSBZ7QLalOmBE8E7CUK14at0QKdJ
WM9FkH0p8vZcdommib9RaHAmYuVVwmXBDf3GMvjenzsVpYC6GbM0baZ5U2iJzDLQ
JJUjGpjJ8p50u8OU60Y2EFAk5d32VEPOBLDILt3VIyW9/499rtfO9Jll2eRhPbyb
n8+0z+WH603pNWer1EObhltTPwcr7elXRD4KODnsJlUSi9H7i9N3rE+M6Pwi6tvb
972UafAQicc+iXuNolO6ZQS5sDS/NueW9rHGqc5QTOF74a5rVHQif2iOnET3tD4b
cgkXwQQ2aaJjIjOq1TynOXr8tByPFNu1LuAnhUlHL5fTK48eFR4EFraA5XIgR54I
+aTyfYZ0wof9vGTT5Dv+0a46T2RkKxXxogPnfxI5vAzgSLqqvE2ab68ukZh5Yu1D
aboES9QFEtg8haeNSRj4VHMqKYs/+zfDVwOHi4AizzZBCg0pbA3y6UOxMI0narCU
1BJvMUPxMwGiyRm1+vH7L62ba30nj+acJ2dwrmgpbd5RH7iMjYtxS1ZMAoZFx7N9
TCviILbvkH4RKVOtCmja/flOX6clQ538+DT/P7nv7AiTRIv8b0ldD1DM8bxH0pOk
s/0HsgDqqOEqHJ/rL1iPx39Fcd+DHfmL/gaC7YX+na7a+LjNeuYcsYJL1J8joaVm
PkS616zlOPnm6DAORkTesD4WoSGenqQpYY79zRpVmfagG/KFUuLpgMZpn3Q8/Bnq
c/cVpthAB8aG+OoYRm1AAkJdEdI47DFKx/KiljYhinpqyWqXpwgfI+MDWl+xZpwT
T0rkwg/8aUsVFDB5SeZ0YBPPu4LEvI8ZI0AqqecTScTSXIQQes2rnd4D0IqEkfPs
VMBKk4PsDQQONDK6bpeK/vcFJXFEbGeSAd9V+zFKA8PfnxbGiOX+NNMj7LlrFkxe
dQgK/t7jqvZP/FTRlqBAxhy9oo+jfebUoXzj8q6ODRCurG+DO+Vv0UrCxwfXWGIa
bRfbwrw1E6L1csWebY+CR4mptJT9JICve5x4EWMmsKicDJHUUsonQ4hEZjwhmANv
AMMbySMAso1D190j0zgOGEjiKH9+r96rYSth1YL7TrA5Tu//qN3FSjccN6tar17r
nnWOdxi2jgKYLWeMojjm0GfqC+GoClqZUL4iQB/V60BXZuU5HxcQWnIYjxllZ1dN
qh68NDmvFgu/rZLIHTJPuo3rdRXzJTL3IyqMCYXQQZUxmBKRqwfiGjrg6ON4yTcL
NVY+/cbvCuagOQOTP9BbtqhUAAiVHISGjdVn23/u4qADYEozwcOpDMbA9q4c+86Q
6wn5bM6VDSBCD/zAVIDH2lPj/305WhsIuAtCdt+gPWBv4tHQ9fnEcAEGclvpxZOc
E4tqOtCcBdRjz2yqXILuYTeOe0uNqZZOdhHwufSwBcvZiBR9pK/MdRPuzTkXnEWo
rfzIipaAErc4aswrKPCmXAdvXVaQqFzqokc33l2BrmgHIcBwIZ344AovSQs2TlQY
wFORgd/R0qlMaLrEBseJkquXFnss4VXxvIeT+3bcdRBr5pU89dzvdra5FD/Fhq3a
EIvAQLW0JXllqtNYQ3z9wNc2JLuHFWEDXiLYvgwL7QmjsRhfEsftqgx1ACn2bzV8
aSArkBUj9t0fUJ/wSNW8D9krOkMQHo+v02fopJykZ62ARJlg0fgAyeCSmyRRDnjl
AzEIyLOUdxDJmt9PvpYMUW4UwW+bF0S+gLc2y2OnNg34iDs2y4HAJiIjc7z1RgKc
s73GIGKpZBY5iZ5YEVPsiS7nGQo7YN6KbgJ/cLPEjaMj9Wz5u9aobtuIRnIA20nu
wgBNCEVPySjRlxWwHorxLxjcssimOcrhpd27FnGgy6OevY+4SQhhYgHbNS4gyUSJ
6TcLMQjHyNc3PQt6lvUKWfSFdL0lZLa37g0u2R/T8xEIGLTWcMiih47vLWwXUQdc
IxXTfq4vycvFLO7xEBhQ8aS9k/W2q1uTxHo1Tzn9xEQeCCC8KkJ+yVfT5wJhcgfY
PKg+mMEpW3jLTs+v5M+veGrPHli4dpwcdHHAIV6CD3Ov+QPfOCq4kSNMSkkvdaFp
w9+7F+FqIHrfR/kauIsgMVY6pbvKHGIwC6WbyFzuknk3akNdxwjjRR540WtUmesH
5CEqVwOMl6Oouh4gWZli5vHG0locNvPuaUNAseaDJvtISDypPjQGR4xS9lIUQXut
PHR+h4p2YjIpyv/7h0tkCrMG6jqRPJU6BZlOJQEdObrvio/7X1UzkmBV6vQYopRU
vL6qZdozimmMd+LczxnNvE7bUkaJGaHSx+ksOUfCqsyffPEHxAzDKcCM6/N3KiMS
SZNe4PL+Cks09SStgE0JsTenzWAwoG9WciKSZCkOX9mDVtQM67OSoNtm9plYDeCh
GJBu/zQRLHWmHh6uA9Ea2EGi0cY1GETnWeblEPDDOXSn81Nuw+mvGHjqWJlZgFGP
Cexf+8Ape45tc317GuXbCNTe5BMPWA/eOAXEszvRXt9LTGQR70zE90FplEaIkUcE
rkWDdOqER6Oo40ZB+6YmIji/jEJgKCS6QmdjlQm2QpOZL1vTBhGn2QOfi6wgg/0z
psk/3mVbylRYscSaUYFOVT1QjmsIYvs8xLJ6OJ+ofzldw1VQ3dTP+8GOJvkRwgGk
tMHTn8fAhLCxa97haeYQOnGdM7Xr3mGsqWonnNTghRzhVWj1xmFo9+aXF+Nj/u3p
jXeuDpNIIyQXv6brwf7CtQKlgBn3N0rn6ZFN62dhJ+s1pVsj2xxDNpA8VXooh4+3
uMPGwzZisnUwhu23U4VXy7FUb3aQhDhWBRFecV4m9vZ82cIBYaGvH27JFnr8axCO
owDn0z+IFsj/U7vA/q2x0BhLyHR6wgevKP9UqHCyN9FRzamCMN4+SoIUu/xT7E/t
GU2buAMmoxa9vv1vFjpMcGIVB7jWym5Pe2TL29XVEHXZIM6/LZibmga6xesADbIv
CdedLfxLTW9wokN+/LK8T7CkUxuVr7BIhYgljR3g9avtnI0051IRpO+/fL4EIDi+
yV1rdztrIdURFSGQEfMbdS3Cck3O3XNwcDDH703b9S323DVYi28tr4VzAWl2zciU
N4uxsS2r8AqGe0MrEIbc/LsP0yzcMftAFuYY6+JVuFxWJXndATgZiwDVgyfqU7wb
kTQ6q50yo4cu+JHc96RzaWPCXpcgGnj3lTDXCk8tbtdAXwz2AQzUhWNm8GoIVAgy
o0ho5vSIKOmIYb401MkvprjwxBHp9VOLPgCyQ90YMZWzeb/89shty8Y28RDX008q
CuVXUN6lejXkpOTOlYjQWt0z8B4kRQbYVUeE/7Z9x5GcoIahsysoLlGCBuHj/3LN
caUK3liegEhHgr67jSzz4ZBLCRnmuavUkodRzaAeR22nWRSDz1nmB7D6bJoKaRMX
HruFuUO0CVPhS06gv4NpOQ9Dm5NSHZd90Xdj+SH51CnfZhk/uQIdkru0WfYAUNNN
fJ5x1UZqD9CSXlphBKLxxkZYyM6xxGR6nUt+ZoBrBYt+RPPQEipVU+q0Mts+/Lpg
YikAR8ZxxYoBqu8ihPPyJH5HQg0t74ZSxpru4v7cmk5zg18nHhPcHbBkShoXzsyF
M73Uhx4Nu6vKxB/NVISzgNesOb8rRMr5Fy1HRhXhyhwTfTom7ifx7UOi8oExoVcQ
0WEbS3dIfu7Pqy89Ntb9YbXA/+8dPiWe5/F+4pjM731EcCDmkUcz+zcyWMELYFkk
mTMdl6uWCkIkt5sv7khMXxVFIW9/bsTqnfH7fko+BadnVdfYjIiUPdlu5YH8+L2F
Xqxlk7HxmkiCafiKQNJtVB0QzmlPNAXjrzzsLq5j2fDlfiyzI0c5YaJtfMA5bpa7
dc4CZX+rqAmhWImIo492yAHFnTQbIWWoTWZVwQ2NvE1ZCcynOztfc5jPjyOKXHPK
W+slDbDK4G1Z9oqgi6V+jRtEEbJLdtdxHnvg80zHhfc/DyR+uYdKWDsiZMpwY7Jl
ZsTbcOWpncF0UC44g+MI21LOLl1M1qcxRyGby5h4tSFG3y9RjEnriMJQ/d15tTvB
xEYMR2r77uVYkW+I97y0XgeT6G9OUxtPm1PxBjAymxn1AtYtRe8U3uJ+kSPQECkF
yv5jMg6mCfi6A5XKbtCpkLkZ69GdBeQ3SMpMzvt9uhoFDw7vqnFTg0sL4YmYSdIr
bIQQpoTROBb3WmMzajtNLpfCjJMUY0rZnDDz/VhjdTUq0Uthrp5d7sXvra6mzpx9
/w+DGhVeqjgoz7aAdI5Q0py1jpOuARwumAibC3VzaZKHMg3xQMF+YwT2Xrdjitet
qfmNIiNmptghDa/gAJQqNWW5a4hZR8eoxSsTIy3strlxa1U1b+U2Ubb14sWFHw7l
q0OF06NqG5Bc+X2fdLZ47DX5UBB/FCfWq2TO36JiWhLxIZ/r0i4tMiyRkisova/F
Dsvj0JgwWVv9VwmdTZxx9S0m36RrJnTfWDiNdMCOU1thXUQfh2FLbZR9dQwV0rQJ
jo2BAQHrNXLs/PvQePQanyDMJsgqaC3T8NGBeDOV4qv0lHk/q20Xbsg6u2RTMJDx
fMOPm7t7Cf6Yj2dnsAKL6dmKSJSKxH1pjW/gK1wVp/0SeQJ4BNDjtc6h3bSybp3n
vN13tnR7zCwFLfdYtU8Uj6Q5g2M8w3ULiDCuaMQJUtI88ApXmQoF8ajqTkxPh9ki
PV5XDzn0LnnCsEI1wSWnNPd6Rg1+dmNFtHTgiU1+qYTIR52JzxNP9scpwf4ZajJR
KykGe+VroTx92OGuAQ0ieA8L3AoHHp4n2M7p33WKHOtbmakUl/BLtdFdV1rn/6W6
Ln41EeXGaLozkgMqaAx9i2qPgq0Ijm0YqoOYwJitCDkEyeJOliUWsewxX7t7e4Rw
wUM1ROfklljKo7iBDENc91NneKjnJPaZ8gRWboNF5rRunUdu+Z8FQuqxErteiZW6
FbPyFPc5//3JrgNBE7Ut/ULDPulkAWff5968p7N6D4wzYpzk4oZGTm1ChcvWLH+t
xYQUV3HBGIDvrDHmiYCOtcxiNMvxVUF8yjmq3S34ANK9VLVmfi2mPXJZsHu58dVB
H9awgwoq3yAsN98Fd+nKCOOS6f5XhVeJMT8E+xNkbOxsuq/W4zvi3VgXff5gq46R
KbXfViZQH21h7vnF9//WFmIALzBH4Xoyw8dNWwbqYjjCz4zteq3B6LB/zclnyykk
0m5OmVONKIla0qO0IGiAX732DEDUk8i2RAra3t5dDWOPuu50FscpPpHpO4I0Qew6
WDhfsNgS16b3OHJ6ETPCQkNfec9WXEXLIOWBt6acCpyRx56Lr+2+UCTuzHRoRVyc
wlLAhFfbfzVjVFfoTlIUpKI39i6B02yp2p+jisp2btxiwvohTDcrq6X7WittN6Ap
A1NNZ2dmmoDY8x9tiRxlhEIxeHeId54nYgBSZ0K207VLQoERhYuUTQtGcu0QJ+3m
NbH1N4waNy4Ou1qDSiHz2wE4+jHFJFEnWFPSYa+RiLyhpgDNS6IoUEjl1Xqqw6+P
u92ulSYIrlhj4ts5hJ71ThqotA//pg2JLmRjdXdc14vzQupkzCDxqreP4nra1IsY
H2FHJdQP63XtmWCiA787wS0XjCa66TVHnvH6m4hFFML7I+LsFZQ54dqk//5Ua28P
KtmAwl3PFeoAIPL+a6pP2LyRDWZ0+1nKLGHytmTxnOa2eJn5gAz+wxAq7mwKxfby
6FzGoL9cvdiJOhPVnjBDZWZGkpS1yb0Nn6TcRANraVl8YQ/qoszeB4z8y7hzx9dz
ghecSuXqNHSb8UwnWN23dD0xwjntGOxIIal6r9usdfxK59bR+CzD+RZvcmSl+pSA
5w05eTDBzUMfYcDTZFwz/ri4aPHyxdi9CTSLM6rHhsTY69tYgKmUi2QQI2a1JLTn
RyNIOkb1aA2oBLFs3bqlP1iM8jEJ6Gr8W4WvWJ9qqqLibSfpYYgkbXEYheuvfr1Y
qJSNhmlE+m1xWHkJpKgqx6vFw2yu01q7vqCKdsb7OkuTQONKFT+DJgKbniD53TTk
HSrykImKtyT4mb+nmNajQeoJ9KJ3E1uGU0DDVgywLIowAEofdmJvvGWNUGJ+H0bo
Ju8iVC/WvvnAr3gSX22yyoopDWJBCAsjFEwL1hw7XRHxtMz4QhmkXk11vg6XrKX3
46bby68zXHu5vlPbLHCd2X2AAbDBV0U5E3M2vqWsUlppg3pp3e/SkFh7bKtuMqZF
1MY1KlVecBuPgQNktiW67y5/27i9nHmxXL1RYmmJPajWb+W47tmZSKbYJChYFrm3
EGro68Jy/md50/tkdnbyOe9Gec4WxDq6WWcIjhYnhVYxuSZnkEeIN2PU4limv3uG
K2A+TPUtCvJUYMZo+hzowSWAuZlJn/ULb+aemvq38+w4LYx2+tVlzVbL5ZPRhhv2
05nfrxAjoOrjPskW8M+9OJFYFz+hWuDDfEW3va6qGGH+918TGi0mkbfUhaob0uDl
EXgojXz7Lsnu8X4CGvhkV6mscdyEKgG14OPTTvOLMY/e/vyJSgXTxatpSVgZ+mjk
8cCEmolBLw/Nfoc2lAOakecUMgAX67I5XUwfvWcAMKGEWFUHcTVnaQaEK/62usJG
S9BNIZy2ZUEn+7HUNH9jP6ORp3CwOqlbAMNilHP9SXTl96AcJgBULIgIq0Yw5pyE
obu/Rv8c8jVMmig2dIVNrMFSBsqm08FwjLtEfeZuzkvS/xUCrFjGjceBIH7iWpnE
zRp6PAW3axX5yl/jGqUlJbdtKiCz2+AYveCs+at1W/NtRu1BhYgodEixo8m44yEB
RG6dwAMzmRjfTDHQj74m+TMwCbtxXKNho5vINepoEarmF2hl3grmvW9SHDeb69pn
/gcOxpHn7E9wU8DThf+9gUMfzSK0fI3ovUs1RlOPRIg2sZFcekT8R/d+0BM9EHTv
RSsSAJG9JIEe34ODPSeQbmGyrV8cKa3yr4xjCWBbt811BmiNsB9Khk+0Sp3cZggi
wJup+iRKWxypktpooxYVAIH8ZzEIOVyTs4OXZ+5WnKT3jHyGC3oMgvXzLHWUOi1j
CvJcUrFLxerHibLR0vKfT+kNXHwPAV3UeNQQ9Erofy1xL0jOc10E8S2YAaheTGlR
agfd/6vyyzeSSiv3xWsu+aXD8fMFQSOQhRb5xnOv39/AjvQiXs/Va95HMiIYneSH
PHW3zMjlhYYkJ0LWH74FzN1Y0BSBsp3bt12JVew+/cpoMG/nsJbRDvqfbqNMJvtT
EUV7TbAehUdejxOfrob1DhI8rQcyInIOXgWNaWb5OrtUJKVIrcZy6Hl27KKsaWlM
vmE5chx/fGkum28E0YxskHh9fcUZdt7iaROfHQlKTcGTFjsZYULbo6EXEZASNbri
Inq4HdbuwHeWLrJLj7V5EqwV9Ms0eUYxIUT/9nd1yhJ9p8rKZsa6sCFrGnxXLrzu
46lvIqXdnvfw+RjKx+wszm/zPnIozX7ukHRJTSLNeDkfVm8qXpPIWlYuOJ5YThZ4
S670maJo1l7Bkdg9sCXrLSES6Q3BXMauIHHbdZD9+ZVmuv6F/dYQlODuNlSLZcG/
vAKRC+1yQd4wDkGxNAgGiaAa3VgvH+ZoI//i4/sSEIESHBDbbK1poG1n61ifMbg6
l/HVtkOltknlrGiBr9ALqZdYcpvScPCA8TZDtFD+3Phi/JxLLNfnUxsTjiKmbome
EqTzouGl537epmdD1rwK8QQghvo1GOCX2k1SKMFEiQr9SBOYf+OoQq9oIFLejBp6
ajxyAGjZd4xVMy8yKpAHBjMns1kcBk/Ef/NBNdfcD0hrc60AHbagXeERts8MydAB
xHokynl2Yd5sj0EgmMcTv/04SEzYZym5jieGAeg5E+ehAuszTBTG9kW0q2I6TDah
ePNShYn1kWG5dX87awjPzbuMQ+O6GIVqQwbl6b1eP0YmDV3mpcbYkHA7v2Xjf0Pt
adGyQnOlxEJX6Mly6Axx4Imn0B5mE7ZTQi8tYIQv6C1KYHVt/P1wyJgG1TrYrvis
c6ul+7P0wz1fDIFREYAlViZoIE5aZ7X1AgLph+9BE1lt1YuBqNqhCnAK49LOKFVZ
Go7VEOvB3ikUOp8aH6o8fGIXZH8i/Z1jaK1U9zUtaURnJbvVl11Ly7ZzymTnLAvd
IQ0hoCYwq40ZEpy02Yk3/8YVAQESqLpl8mbRR6oQei9dkobIDlXtcd4CyaqJ1UcN
u/EL0WdIe35EaWTFoCybzCl/MvJ6PD2ODHD62RXGRCDrnMdMdOupnZjfFKtS3iLH
aw5I9UsfIDTdhh0HJ3mlMSI2CkcPHJPSqW+myxyhUVjyXEabdCQ5NYKcMierihQP
Ix+vHnnNVsutUBLodAC6ZlMPdhd9aKwbU4aKcsS+cPRQXxVr3+NaZn+wxoHisV8d
xQNXXGZJ/nFxkecSfMj0LV/xKlxJEOVO8km1YFNKEJcOmjhAFsoLtDHOenamCWlJ
+Xia4qu5is0pwOmjHwDF3OoHmXUyvdHmDyk5QOjCt+8/eZcQaszEdcpeTsOY3b8v
nztXWY1frAjhkGIDqKD4etWsaYHnHvxWwWAbN57Pnjb9tAYrcvryUoNddrLmOgLO
DUwwQ5ZGCQ37nAqF/+jatUcIJxm68zzyyZUBnPmcCLytRJSedAlmdwKnwgo8sgfv
2UppH7Jv5odfAWzHN/+4Ip9QRvMM2ynHvq4PfUIUfIx5r75AUxioRbzDPmCS5edr
HKu8/4IU3b/9QxBivOmSVVMrWmhNohBuWi45Gd7FoHMN472E5Pjh0Jhz8QKC3Psb
+HSs1I5n6jo2+z+83N0xJM9BwfMMrgoFZgoghGIagcm26+mTdA3ncKbH8ULIiTMZ
7IU0fCvZm8kyfoWmVD752ZRCXGVJVJTRhe7TuW9bmZUD3RKHxOFgJZunAzjRAUZp
Z/b1Z6wYH2tNYxv2a6brU2mfkrO56iczoYqKhLxABTDavyYCyJs+YxDgQcIBqaKL
NKEkQ7zk0PRcbNhP+EcoSZ2KyOUCCON+WYk4eqOGH+7WUEo6LGX7z7XP2W5FoOiF
yWdyUT3FUXEt5DwESQZXsrFs2Sb15HFsisIWf4Hd+HJhJNvPoGwLn9V8Pt76FqT5
yblfOX+fMjPf6fSAXJwWgUPiJqxHCu/42lDY9DXiQwXf+qwsRiWNGNXjdqDY27cK
XYfo5iJGXAkrkeXYJ01scacZurg0ifGJn8FIV/k0qoe4VBJxJJnnBzu4P9UeacjZ
r8zt3sV2j13Aladd5wFACLmqmFST0IPVr5lgxuO+sh6GCacvdAI6m3Xfny7GFpUa
VP7Lc0zQKoeL7YAQpiu5NLWWnNgTJLXfVyIfycgDy5jcRNCoxwygsakH845qhW3p
Tww3OtefnuCno643fwA73CGbr5Gu7uHUUjbrSheOelmcP2PJwvTGGo4yDK6yo4JH
0UPS05oUINL9PvMYcgb1F2xfXf7wL1qlRvM3+fef3W6Es+FS/0P3/Ll/YgQ4Dn9Z
c6P/JN4OT1xIHN0jQbbL06t7sakRpOfW5TSDMuQFpkoNx06Ir0otBqV8fZf0NVxP
ZNxPD6HzoWGofiDop52dwfBSMge6egSEBzLJLJBGq3jUH7RM86+F8lmhBEGQAOPf
NDaWpTfA3FkJZc/1cZY+cEG37bnJCrAhQbVcgZPU6qsG5Y/BQ2JiMoGlZbD0yAJo
2ywLa74JthZBfHEGuk8dzy4RusE/QbjlK71LN49QqC5qLkEHFcqYs+Lu9HbtoOK+
hRPkW6J4EZ+ADIvwbjuT1TjRXqegF3ePNRjt3TfDxIE6qoC6yWJDbtAff+p58pdz
OXphwqsBnBQ9p3OVOVwKKgwKSu1nF+omevrWTKIwvgJcYsIFMiAQ45sf9wUS3/+k
ZtGJB7THlCPszp+vP4aDIPaRRm4Txs/BkJKU3BRxT6zqBlhnizhtJWrW0A+phyOp
ROlY2p4PRXLsQnPLJEpHwxKdFCW/hFnwoUcf4vDE1jZYwwA77XkXQ9oAOX/YOoRC
GjEuC9arcml2A6Q//GHQZ3Lm8SEASetYdr121BfJmnoVmg1jHu0OMY8imC+m2UqQ
rpnYlgmBrw+kRtI1y1ZGzd9xo6c1PDA9pjUXsr0/7r+vTKFGJXP3flEVL3/Cx5rr
9mc5c8hy0zA81eUzkzPhreLMAj7zwCn1o8S5M3VSH13FEWpnwiSXAP5Uo17TLx/m
lln6sn4dzwWhUJHS7kxBn2hMTlMbEGOAuTEJUJCifsGtjVBkAw/XMMSHFUbDYzFp
xvXUBK//iBUoE2YheKoPX6iecCBy1+m3tisUjbQTvYL1srGLShF0ryDYR9VRCGe0
bN/nMkyKyPR+XlOqE8nIOK2Ohj64f0w0Ekf6D5RNVDoVyuRdVmzk+8k7HU2nK2hc
CoHKzZzRay1irVlxzTePutgalTBjNP+l8AI2CaRaA+Hkb1ZZFFYMO1o1T+FBawDT
pL2GqOnbCzOBDI1VeKmcnmU/y1BbixDpurX9uiEIJQ80uMX8CdJJ6kBMrg0VPp7v
sxmaAOTO+rg/63/T2STN0Ph9ZWCLQd9fmYts8Y1XYSvc/GPg8/hLF+09+3wT3B++
yDLkYm8RyGdGi+okF2UUCcMGkogSePJBpINdC5B5qe0q1WILBVQihiI+cmaahi9D
U+AeDKP/Zbkra0Hz4+1DPS1bzoI52Dc/AMfEiRTbW2SuEnu0dO8RnSmPmxefTWUK
enwL47ZXY6QmeXfFbJHdQWlCYMCog6JqNj0RZZh2DBZRldUq7RVweo0JsCCKKZfK
TCamBN0y+Gz7St7BcW7HwoHHl/E3SvOrRTjTtsLCAAg+CQP+XutE00DMU8/ymJTq
qECcIg7y1tgybjVWXUntU1g8G/b7jKu7KOAVXv0vJaZioExsc4DE0T6bmtmn+Zfs
Ztu32ENbOqpjGM1HKcSDI3q/EWGlFjuDfgOI1eBTUPwvD8Vp/iN0ZUqj+p+5N00i
ZDw23jFUA72f/pensGT8v0wmzrvoYVxSVEH8lbOuP+3RYo7sPwX4+N1tf1O1YZZX
QrkQj0Efk9PQNsPzODt15zWPfKX3iibG9zGx51W/polHG/wOhLDu0zLRisiVEly0
TCS1vL5bSFejIYMkWqVlI4zQ4zoOQTXiC8SlPFHtWrZrqC0t8laaMqK8nhSoyB5M
JIt5Mb3cZ3kMd0PgLFXJyVY7rjZiRncrrmG+q1yw+P2s9/6e1sWNAgLPioLksw1K
XF6yDuD7gmdY6VacF81OhsUMksZe3IPe5g/2dAT9PgnL1l8XKqBo7c7k+tJMUj8L
wQoKFCw2IVpmaKwfX+jGhHluyqxxU/evWqasbdsQI50eeRpv9w6V7m0L3mawSX9a
FuFP8lqg0QzYNaqJoYWmpmKtsvC2Ew8gjV4NKrCmQjlbGjHpxMLmS8mTx9HksXyA
9iA8kWL/UsTjI2P7+DiratnkaQQ1HYAifevQzcp2x8d1SjH6fEOV01m4sR62awAc
d58p9MLtXwHirdM1AkFOJUU80m+XF3xwrdN8N8CRkg9AUTGsDmFTBqmjBQdGrN3C
S0h+kL3OpCo6j0vuwSfHgrzAuApqom2Ys6z+Ygb8lTLU+KPxxNN2yV2GR3suPDei
WJQ0b8VWHHW6KeZwrGAMpF+MASchYQCzXcdpZAWRREz90feCgEuEaSiT83GERUcX
ZBZKcltfQ8URkH4nfm5/Xwh3rN9+492uN23Sz1tX3E0HeMtEgO9zy83a3TKHEt1z
k0rRKVAUqHYXvLxvb8XsywHQRzvAHKJTybSf99biWe6sj9lf6LQ+Rc5i3SXd1OzJ
+z2K5qaoMtnl44dPMrkR/rUsFvpNjUWVs8P3IXGtQYBQFMq7TI1CNZjdj+Me+kUq
rZFw+QlfnIlBhy/hcOl39CDL9+78AKghCNEQCJYcuea4NG4XNau0v5hpNxxzMIN9
dIoRLyGREOny4Dip41qJEAUT0QveFVwwtLVhcxBkS2EX8f1YUwp0EC0DYOKVUerB
AQIrNlNczPyuQTblsNbrkI8LXwuyJAvOmNAU1dxGL3YBtnToopnB9PbJgfeAVpw1
N4mk9LjpXfPpi6ODjmxxiUAtfdjt15PyBIERaq4jmahi79OITxkai+iNvvlzZ7B5
8LIzLYOBZbBh0Qh3i5ryiPGppSlYFV51dSmtqj8xqXAQeg4ccM8AYUi2mtSHtCjT
iN9F7RuSEQfPf9RVuHQmjyg8ynIjTCeI7uEBwJZp0JO5W76IJ62096mowv079ZR6
VewDOrYSKmtN/5UdfaMJg3IKSHQUJ5TAdgeuI2DUm/Hc0eAWEAqHDwIpwpFljJj3
8ZJJfLrmSvh0CU5q/VvTFhSe4OHrzeylAuLmjiZOLLnIlydDmNpjnoL1auJw2vBh
ywzHbOveBVJYHNNvDZ1NGr4fw09lNphFpT7JF7NuzI/UriiORB+dMt2VM42dZeg1
zAVM/26NPoPNCobGntq/q3JNtWgFdj5pTlIfBRuQMTB44ChILzt3BQITW5RxAEj0
WCzHMIXVRf3EBUm/SaoHL0Z5CaHu+K+uGaItFrs/A4fyUCnAV0/3Dsu7q17HzUEH
BiSvjE2JoE1yA/x11UcM/8vOE96cdGo++wab1PTnaktNFXU3YKTmmqovF3Nhg8kc
/K90arBTjcfED9zOjKnhXjfxM37TpOjhx8tZIOYHEsJ+FqjC5V7TwE9zDAsCKj4r
q5k/iSpWWvekaOzJewm1TjLTXcITGSFHZK42jF4D1x+KufIZ8An0fRqFN5ranQ4a
dA5Fxue/8dpQw7hGDePA9Mnfz7v8MRVGhHXNbzLbu1yqjcwFqZRE1adrFvSFjXpE
JHDvxaHsMS8Rya9DoCaL0JEIqQRbIljAw/3q+QxFn9VwXiTQcEDC7SwWx49+FRP5
io9tM9IP/8By4VxnGZ70SOALYbyPAAbA6CmwzzNNBIDbMOSPbUGafjXSpzIt+JM/
KJLgWZVNpAXq6nblSS5QkdVAyzvvO4e1MhlQkbVSmTMfYHEn6cZrCN4zrkUQJ2jY
yXjnScoX8fEdcD5dycTkEivgehxfro1/xVb/PX9Cm05VkPe4A97Y8ECiPlJnUnTn
XxFkzGlisM1dxZi/UcAc1ZEOUIZ+eYZsKmlJpUQ9vAo1hExPUJSrDzDldUiVWMcp
X6pttsCOGIlbUvKxoSjuFShN19V255qlQQ0QxvHiRw1VK8s5Yq5oesPM/EvgtWLT
Iw8CMc2rT5JwNZ2NAuT4kppgpCuBw5qnnHIAKWI+bYWud99Mu4oaGhGzytmlD8HU
uJvaAscR7oWXXYz4W4Wmcz6vE155mtm5UZ6LP5Gttsu/TVya0k94+zjMS06vDN76
lvuD2r2JyE6/1zAqdrapXoqgpC6BaeqKIISH41pEPNnVl1xOhCZKH49qbTXMNtw4
IK9fw7Hh3hsS9mdtiddpoxbX6wL37MjGK4W1X5qv4ngZJNoOIpSMwIpQbNNKxR9T
I/itePs3ivA04G8cnaksE5VN5gBLPAWvYwMdfh12lFF3cLdMH3Vw8w8NiMSkQUNN
cJ5+COkqK2STU3FN3ARfHY5ma9mNK8FQce10DbYtKok4H98IABQAsdvp1Czu/Twj
TmZ2f/0BnCRiBpQ/MK15mgafZNtLtAhpa8HzHlGuBB/fPbKw2W93jbDiM7Gqy2tJ
2Ipy0n8zfRimNLDghxkASAOtxC3aw2iyb7hVa9W9WF171vkEOhaSHDh8V6Pg7+hG
F73IVKBTqPiZBed9k6EX6pX3kS3JXR9RMcatiMUU+sxS1Xen55HYUuOOaDX6P+sV
IW7Uxj5QduoYc3Ek5FKpgo7VN2w9pgjhv/fwTEokotV5G62c99i+IFl/LTgxN5Pm
Rv0cchPbu6rULg7MzgVZann4ef4/MujOwhTQLKs8oibUrEHs0Ikij6nH6dk5iaF7
JKTHxLukKryxYofXB97wVjHtc1GJ54FR5mVB6EyVMhF8JpedkIShd92Q0g1smXld
hlxzJqH9N/MWQW4WSNLjkMLPFeg1vqlZYgKrMXmyOpm6XJ7Udt3wdyL6g/HnzzZS
wJYx0CxBpMBsgUp4fs6Mbg==
`pragma protect end_protected
