// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
WhJSOmywPNoQOHQhh3Qen4wWPIDJi/zShGspYBpGHCIHeWyFuTRj5iftVz5Wd6P2UHrWn9RZBEky
Ed54IKu356tMSrAI9G33UgbiZmTrkORWdzrnViYguYjPhY7HLdlymI9UCER3cPLr/otl5yj9Bhlx
I9iePG9W2nywGCV8TA0cuNFCpUDFoSaBP6Smz0rznMKMBF/hIK7XP1hqOgqaKw4LKH+DcGhDvvom
WglT/Sy+esK21b8eV5Lr+oaw2EpT9Eu+6kkJKr5yYSPzH5fFY3T0X6Exm48zQHvXFkR2/7+Zx9sQ
RVxeudPNyLdnJSdfulQudnU66qODDJ6nMFAxkw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
7aQNK8CDrQw93KwQ37kI8hOscKC/mYW6a8zSaJrDGrwbm+bG/zOjf9WDAlQS8CdJX4HasfQ9weHi
8uYz2UUIktdtORKU7BEgEZPHPOos0IYU4q25dxmmzMzobhXdWZcNyWno0wBPO97+SrMfrVNcBSJm
yBR4FIsXHmgtxUfZNOwIFqBpfH2JuorcobHz0uZ1nErz3HMoSBcU1BZExGeGLB7xRo1RgNCf5wIg
cSOAaQTecbPd/dddWdn08d+VX238KMMXQ4yZzqcHkMW1GhGQ12TiBj826cVnAxfPJyecm/dSmWTO
/VtbrGR1JnABNgAVshuwpB0635x8mvKM8aFXcWKtMlN8Ziz05Y9LkJ03Xw3d4RFYKJN0hiQgPrcE
SicaRNwh2NWMOWqRtKP2gBvmAcXjp7+7wg6D/R76toZTB9Y3HgxZ5K9WJa7uZVuSoXADrsCJ7OLe
243KaPpvM9jkqqkHzlVobI9OCYsvabZESwN98++NgFdbj6cuH2jurD30BFSuIReAMBM4lznnOS2/
o5w/Q0vDvf1tFb01HdwwUVKEPueKJeBL5USRZDIgM7lOfGYgq2D2b9MCJAQ06qRG9Ve+rCm3rGAK
k6bB3f0QIFyVGvH8yg2qc+FQN2BHviNWOCbMt/PzkeGBedRvBW1FDwqMP3NU7JO34/ct9U1O+e6D
vjp5pDcvXXqYeMjpjQ09HtZRGSidYf49O8PLKzFCTRKZjbxDHPTdLrJ13Fgx4bjL14Sqei3ufb44
bgwe5VFYEmfDBElzkig+W1I/QhHpZUf7KQT1WvYKoP8ZwOl4YbeNlUXftj7K6Bd6ttatNQl9a/tw
fnkE87jV90GSrZ69R1xdoziuUzojFfvbn/FwVk9PUYtGoGkVU+NUXFdjWNvdZL3tHnNTXGpQC+Xo
zxLIIPfQuqhs93/wQAh1d2JozRAUKzmYJR5PyHZDTDiWp14/016OfO/0/Wnyv287Yif7Hvi0fteN
iFU6fxzu2QHpdMWygMokOh3rykCeHj8w40+MgBF0bPVVp22+F6mD6HIbKDqKl9E7WLNWCiqypxCQ
n++QtVbqgEvAk4y4rihbfRcY/qh056B3UkPRZBYQAh2mwzEBoL90XQD2P/lgZeU0MtY9oT/dfAEQ
+FHVJzDa+zFQzVAxK7uposffK6z9wnS3bOSuuGlAty4gsaMDk89onzUAiX5pDxbBQ3ZojhILmbk2
YGqTc3feO9i8ITnIVnzwJAKluz9+HO3MMYVhkAn3fGatS/Og+POjZuvzyCNnEKWt3CNxXfkMf528
ugco+rmFIYAbRhpKV9blukLAL8cYHEAWIQ92CnQGtANfZupsziBTDxUkk7pWEVFAEJZQnpB7d/5A
dqy+TtWKPjS+GtXFROXj1sY4dpTkVtcJEJXaQhBN3Igii6Pd6Ek/Lq5e4dIMONlts8Igtgt5BZG+
mISVQdVTR9we9oIwHA7GfFREslLk8n94YQuj7chQ0BrVfcn5X35KlJ91yKk/eGcmVTcQFv+4z9F7
3wu/1sxaldYUQm1Q542NaclHBnuinmdwuO1Y03TC7QIwaSRM7wJZpg8QhP9W+S8wUdTx2WicjROR
j7iiyusnUDPJUKWZGvnQ6dC/NuNu9gxriPN+f7mTLtiVAcX6HJBetlnyT+kXJkFzBKX2XLylrrfs
84xmDBtbUORBAoDE1gnL6mNpCuZwYhX0ZGijK6rku6aV64excWpauqC76D0Vje7Iu4y+f1jKo6Fw
73Se3snmLA+AkzCfZpppogGXuyDwgU2Q/9GzvuaMAYU5SB7t84I44eyWAUyf0QsRkYLv7+pu3QBj
aaTdDA75ObkvKw11EVBS+58dZE5XiyMBMOdW5xVVvRVRDcQtC1gIq2eDYtiqQQc28MUbuqpneVOJ
aJXufeNRCNhUxWej7ddjjJUyaZFBl5KsrTwvCWLJWdXKH1tYKj2pJQcfBrcp/G5Uh90t5rKnouEV
MCXoq5ItqDQy1ENgICJiso/km17XCGO0M5iE8ckkNR3fEKIV26ScSlbsqgxqGQS00R7o/F8r9N73
ynxVXWFwV2lLqEeeZ1RXXH6fY5+KI9WGC1QzaeZ+o2VVcLtdmbXNsypNbRe12Fv5kk6aKqPjKLUu
31GYjideuBvyJapYKNvJVLiMO5iLHJ4OdyNyrpNGRpT8/X6qCpuJFFc1V+JZaGFSnCHQVyZHbHqN
ggmFpcrNLFMbhsId3qNocmAjfgkmxVI8PyB3nAqaEBsKabOM48i6JPzZ+sk7BrzFEIvs2+7edYJm
YADJyta+OlcrHv54zPSRkJTpLCYbZaCEIuxbF29ZS2oOzlulouhaIrAjIQJo2qR7U8rnOxZIBXxP
z/jJqZF6kkqbeRiybzSGpjcX7wizZNNj+Caum1fZB16uhROILW5EcyeisOpNY0BGPhWSGJYlPFSu
uZ67RafzpjmP8H4mdmh+Ec8VnlXLaSEEL5l63fp8/u/8CTPkyZEmv7TTh8PKrp0qpgWzngicGqAM
tng0W2yiZa2gki8tEJMkfVfh3mFkZEIwv7NptWbyYa0mX1jXxYMKvI+DS07glXq7Kw2Lehzeq3Ru
Utw89n1OtpBdeCy1EneGGouVyqgCNzEr9dsOBxY+RNWWWJsmH3tE5GKqbICHWWwDqLbD9zaPvegv
LfFOa82W3pDtoxwI++JX1XVAdV9gVSYd5KyrEIOSzdpUCnMhF19Kvdl4Wg0VyPHbp3C2tirDYscD
RpnB5LFyoB8VSgSJR6e7QDBjH1U0/aYnDknNIVxRZ3McF6OV+1xoJjwmy52G8QprmRD34zaZztuG
pouTbdv/INA1l0XsWoZGPPgtrBVhjnKewvMW1n2XBQ4ZStJGkAxLIYv/ObXSTi9o9Sg0KDgv3KQe
zCbCjMyVRMld/IcW8DN6238QojqLtRX3Mgkj/u5Vrmq4lhQDQjJOaOKoatAPExMM12mZrrvvwM9B
XSAp0DaRU+tO1Xtu15+De1LBe1VQWl+vQHYOThfeWnVZu3NtvPFoGsbLQHPmSFSuzM1jSrxxFBhy
CMzS6ilG+v1CJmX8aozEAUzFHxjwDDKYuBk/dytrN/5r2rmeXULMSSDfAFL5UqMNpv7PrcvehOk4
oImD1MeO8zfjzuMf6GBvMGEiKfFjvvTS5o6tItiiJnKbfdluBuhs0WVIPU8e02SK503inpRVghWs
zJz8JGtylunQmNpXpBBZdqJgk4kQJG6TCWlfLn0OZxG5uxVPXM2EOpg1UN/ZgryQn0ykFkt9yveS
eDYi9saMCo394udo5EPpKnk6Utt2pleRC2pmLZtOynDX36bpTTiKyz8NMl5hu08N+OmAjyR4N6Bq
ZngKL98HQSlO9E+jBkdXOyMbCBJjf1nlRkSNj7Fu/1scI2T50AKN82RDTSN4kNoVW7rMTJNc0COE
h0q42dmDNF55Si5XAURPrUa0ZpMF5b47vtoBAxtFcxNzW9/i/7zjowaYZOZtVBrZwiQLCd4hdvQn
fNS8Ta+N6LH9dXrPwxh5016It8aBghS335nqyvZQgQsZxpOoZvdGHT7T9xIHlmDO/fm3/gb59oJu
oVRMAxyoYDE7ogzlYeHQxsu/TEBq/a73/pazPbbmdLzEcYmTIFe3R+rzMoMOjmOydoZjqVOfu7ic
ObN0H0TTwYT76tBKfAHwm01KgrC9LSMmcF0fuuNyRuYY8E0T57tGKAeF4/V0dANQDSTM7xAfpf4Y
b7xepyMoUKKnvwiSuz591oy5Qn1luOBoHiHUg6QxjnpxH4XOVcWExCvmzn2qAUF1wOZtfOgCOch6
vm36K9eSSLD2EZ8mpxfCStHeqTvUBu4hoMhhyvWN7Snq0YVSbUnoxa9QsyCRUMWKmD8Cjst6E/oJ
25ZCwuuNKd3qEYbh46ywHcKO4RpYo84wTIUgTjwi2z70jFvt5jrhHEijKPa4zgTG0ZZ9HZcSWsed
hJATNB6b+B+u07k1rqZKrHqEbxxZYSBXQwILfyCcJvRaQLigsGdEBJkPucSZv0M4R8pnNaZg2/fQ
VYVOzpt6Hrel0NPDGrhM69AxA9RHF85hF86PjCUyapAHbypNUFwDEfvTKeYCuf+dJmRNGILUss+5
0nA39Od9pJAWCrhzEzsNA0lEBoCFjIG6CJz4N7tom/TumQJ1wEHIeL/dTdn/VZ9qMWBHVy/cz/RW
teQK7qiBH9eHJCElqO0LzlktkEo0bTYDx1lFI+ybkSJIsXEep6luwvmIvNlvlwyaQACevy3xiStH
Fy/n2lkPhz+QtqwxQNs9EYKlFOMxI3nfVDJuRm5HAueCQr8pIt2hc5N+kJCaPjmRp6bK163YYXOx
g3VLw5TuTKF2C0jc2A3b50TCGhsgZZJirmygAosVMhde6qBrhD4aYjYm97YL6sIr+wVyC1FmrprL
RD4Dl+sBFNbbSvFfq2AeorU+zusnX6R6tMsnSrQy/rpY9Dt73Ya6Ruxo+wHjGmXOflVwDoFlIk40
/LPUG9EekE6zjl0FO786YjJnBeznmipksKiALLMbs2W/68qcMGPZHWTKK9iOYdZJbDcBTDgquxAS
raWdQJVl/gFCsEN2+jsvCixjhJY+THDW3qDHubCG6RjMndTsiRHNvc3yRutx5LRIGh3Kv1qoQo9D
7zQWHEklHtt/GjXl6RDzTCfjQkB1yDZjVtmbp2Wh7dIrqFC8jow9COk2rkkcbU+veubbA3NzvdZM
uNvzy2QZtsEVA5+UAb6I+hhXY3y5S+ODeuWTgRhKMi7avLbF/YxWtZ6pQrkSuQzkGIBVuVKfFtxD
oH1h/O56nk9ENfJmDWdL2kumhoOQiCV1YpZ+kGqW+e4BBgZq2Zs50hLKHC1kIUzpwesPBGHNp2YM
hYAj+4IfghalwwWqIzkDm13CuprEpkHFYMinKSqz8bSyyKnSrUTDbygkpI5vdn2PLcEBVQweXdQv
nY37Qe856xle5gV5KJTB+krDMEOKoMOstmb8HwUafmgMr2AGu0UA61tbnI2kTMGsx4G90dFktzZ2
aWMYlLT3Z++hb67ZJ4N+wStqacdPauGJXZlNe9v/5iv0024JLnHDeW9hoYflc5fqX6qxRpE2BwC7
VBOCz0SyitAL/Y6R/LEBLowXFecDE9EbsvWQdnpcq2K2/Y/DbgQTYZ6gnaqW+I4G2/SulSlHMaHt
f2BOyRClaxfDLHHNDLmq5Dyn802t872AqJ6v/UO00wCbhytxXxdaL/CubtTH/ewkWROW9IGHST+Y
90O5jux3NtiF5civK+ochMnpK7QfP9axMt4QalW+UQKg7rH+3t05PigcHJT62ftO+OnYoVQZzw6e
dV+ioe5TuKQ3r2iYmcXmgeHoIyvJMmvMdCXBLT+ubofBglaLZlrBvxSipcKLTsnT5YxrEemsJWrJ
09AcJh8gkaCWtnwPc0ShtQFXsi/uuYQWlUJcp2mhUoVppGarPKYj+pwVrtwRAN778IRRV+Sebhi3
nEi8dncORUtziNe9P48lQ/Ely3uhUZv3AqvnwISdJQVX6IM+LXbLgWXA5/QUpJowjhZi0wDwzvrS
rXpKUFlOmNQQEuuJmYVP6o35mhsbPg89n8jTWXIRgEeWDTjfhyvLOpgZjHViXDbcOdxyIsN4oUKD
4wnepnhKKnSXFZIm4FKkHqorsmEubOxNJ5jny9+ovwDyKi+ch/Rv2bmZ0j/etmCRjGIB7GqGB7ZW
YLNWF6zDMeOGgmgwH3GupWWZTlH5r+zj3cqCwnoxVFWJsLzbz6Q8P6+MFOd1s6+Kwp9qHwG/1wzx
u71sziubLyOlcN69UG7u7scIVZS7ML8wBTfgobgkdzblMtmN4OIPMN4xy3pPqQq5gQEQG0ip3Lch
+laKKfduH3jabgMsloCSai04R6UXaezqyZNYjd97o9kIsJVj5119bTKAzWYnb1eui7Ug35g86T0E
Oi0CqvMiQf2jIQIGJpikiK0gg9KDBHcOyit7M8/PhodKAY+/3BFNM2XEE4SH+OLx0sxuhUySzAev
cykVLqK4w4HYAEYMjk6diY/bsm8LhGJ9wcuFdcfe4Gm60SVMfQCh2gPdq75TEXNvJbC26+VdsBOe
5wgRXYxd+viYEpOl/X/Z/M4i7aRsqEemZh3OKFwQDRkLOL8m2OaVBGZZ0kp12cip0ntE7TdzQ+JS
+JNOrKTF0Pazoqz7kXMuQQltq++6hO3e3KSKAwz8FTT9++Ugip+yGpb/PuqqjNOPNxfS/BGZ89aU
Q+cD6tLFLS4soucxAAw1jNIKeDScULoWJdlFg+eLX3zmC+16+EE/ILuUbfbgJX5J39HeSzzfxx51
U+uugqv1owCC28HxehBMc5Cc6j+B8e2IMOpu7gClrY1lD5ZUF3dnbMk1d3MCfclRATlK+9nriHmD
rpl1YbIgpHGPvNKlJanvkf4SaMY1RUDdj8FCL5RmdvSZuR+FI/fMgvkrQexOGPp7YZsTCPIKGuSL
D07xAnPL7aR3qEy4mhT+BOgeizzyL08BAa3latmJMTRKDe/MepY9bMcrUFDcJrO2+jzStmWhGC41
YrciBuPNPtdGGkMDDWai+Ee4aTWV2IJLtmq5/7+scg2LO0521Gsnw04bBUG3Jz3bc6EPLVgqKZmu
sP9qKZRf6M+kE+EQTVBc56GCv/o+rSesGHc4Emx1w8JTroNJiTbCqNUqtYCjvOxYQ5zQQx8a82+1
R0OEe2/wa/ODgcue0l3COVZ717Kf5VItS/WeCLgNwdqNlDvgAcT5mOqT2K4mVJ4GwtTB5Toi3DFx
zs3lOiRtjo6rsQb83yhgRbP/vWDedqpdOmKSkVhCgBkUNUuaApqq/yt2Lct8HMJSrbC53aDa6jhD
RnycT489Q12hYc3iPw13V9EhCdZ2b247E6aPzbYfA+eRVP8A5LO5+mSFEw3a4M5Fk7uGmxhl9Wqb
uuc/yhsKVAOu4YjGoyHQVCK7KeZDK5R0ymkMOTLE85FeCzAdP8Li3bECn/XuUyO8W8f4bR+eXkk+
c8HQYL0LtiyT3rRM8kNWUfUJz3d6RW+bqkBz1pcz063Gh/rLB3Sts1IEUth1yC0sWREQCvzD0ebu
Hvg/In12PmsXq0Yw0DfD6PtM9s9Qw8HZOLmNnb8MqJ3PGVdVRV/td6FB9tDj//YkYGTTX2qLzzlG
uSyObqOBMl+qGjksOsa5NqzfFJd22+dQcGJSfmH2SCed83bA68xXj/xN7T5XsXMdOcOU2fhGruCZ
+sGW9GUyp4PasGQ7VrxSdYLNREKpu3y3diRk5oGjhTDQU/v8GNXWBFRWFlt8LNm31Xr0krsDoBqR
H/vjrRQbW68sRwJsWlW4i9xhEpqE2wnStsZtGlrPI1C0Qyh8a0HSp3Iddg/9AmWvz+I9Eep8+53F
tKxp19zfGcJOJKyEAchXzRezU4cSeK2IOslb711uLgVgRYs/6+j/Lbl+VpcrMROt84jaXGn7Igdu
grlY98nHqvsWlA2yDVcZqWObnRzOQ0ScLKdUW7XMUXqEAm2/IIL8t0LZICqYxdN0BQOnzph030J0
10P3JCo0QrecxCYA25yAUuOq0+EeOrQ22VNTRG2esk3XP+YHCMIISsY/RGSjFhtQPm7IUQ0thnnN
Oj1QfD7mT4pV5D4YWP7P2rol6gDTlMGUQ9X5YtJe32rS46W72MBKpxFsKA3dbv//E3St1tJ/fmJk
vopvpy/g9hgId8atL2d6PsD10Rrra14BN4INXn460Y5ypV9qfNYUlAigkn9D6PsbJzP1lf0/XkfJ
StiImJF80Q9AoC+hguAOJknOuJSrteygWH04gD42Nq0pzYaEfJ/b/gU0deD/MDI+jrz4+XkJbiiu
0r0OfL77vPXdo+DUHvH+nFyJwIaBk6scGA+RXgcetYWeXc6cqCrIVmM/wklA0fkoAb8Ie7V6/TWY
y9P7JrRHvcbZjThZT1BrBIC/5sE4rlZbICFHC4sTyXupT3S0rV8wfXV/5phKY+XjFurDmQcjW2es
7TwkYD+1gjtyB03b15jNM3dLHC78Wsg3LVRppUfjmjO8UEqyfna+/9S52O791eEvdF2zOjk38Mhm
w/XtSGCdz32Jg1a0hkV3Acl6YV8Hk+16V1fm8ztnSc8+i78U2sPcYsN1jshibE1n9h/zm5663C7v
NOeekuOlr/uP5uu2URx+TPoIEppR/HAHkzzB6wB8uYsBYmmcoysL6gnm6vYv6f3z11rM1YneWNod
sgjJ7ljH8VyIXKlie3gO1nfaGHqC48Edx4C9dkCJ602Zf5BGhHxT4G3PDq6FCcfrumapfvk46KSI
gphjT1HzLt69G9VwE7JZyPrRtfi/WtiWKnc68SHF+DkATBsZPfXcSdjM1cJyKP2I3PYy0KP4zgOu
6lmjqvfJqzjj+BU/GnqOfsmiFLhJfQjACYb4IojOFuz2cA9Jp78SG1DveTk6GVTjZSoGOFdxw6qb
aRfSPM5DGDshJ790KNtD4cp718bExrHHNl5IgVWM5yF3sYASqXrr0GygN4qWNKrPfEEND336MTMn
/8+7kZDeGAlFItawrC9cJfWigaD5WeoSjG4YIGpoiXXLSCVwwxbPhGqh+PV/78ovoTUjLZ5GXLeo
UjrVCeIXkFs771Ll2jOPFmOUgnaaglE1CyRfZr9q88Ro9VaoULxtEZwW9/prKH3vcbJW+VLaL1PO
+EzvNwo6iBUjAxhSL6v0pyww43NrQCcqqOYeXMzdil4Mu2Aq5Hk++8K16vubEW7ZdOaHUSulMvUQ
PDrfuEydz18LZib9FEHHNi4uoQqRQIYobZeeiT1YQV4hcFMVd2GFQSLNTT8Bb4AdVDdHQutitmGy
CzyvLgueAJYf1Lmg3srNwM04UeeIMCDYFnKblvf14RmUMp1UP93O5+TD+Ct87FK84FirxQAujMxa
2v2Z5zA+Zv2oY+pkFHIpgalGYbciFedeo7IKkBm5/9oo/vIDsEnOgmKbAXWtuCXGCTkbdjxqHENK
GMD3SWKw0FPIO24ZZ0LTndr9iGIV8gpyTy5ad7ZdMc6NmcrarQU5dcVPAuiIPZ1IygMOB98iR7sx
F+zeikObMgJJy2jyUrHOdr6WAXpey0Ujd+5xWCiGi8GQ4xw9RniKSX5rJf+xgLb4B6iRkk5jlOEn
zmJh8ywdcJ0BZKRlFTqoSQfuq4r8ZkgWIyx43EblhF1NXLN8t9FmP2aLbvUmfEKz24tDmJJBDXyj
j2uGGKz0zkOmmFncNR6XYUdBO6sYRT1UCLqf4ItdTXW0hHSGgs2pOJ27mMvrx4o3XIX3fF0OrpqH
g6KMtO9twovkdy8ToHOroE7vxBnwv99jUxvcWFitkwZTXXnROJTxDWWq3PqekHiq53RIMMOy9vxP
9/ivZrhCcJqREm5pB+D1BOWMbwLYy6enrM6kd3JI+IbCZQevA2+Z6vzBM29PAHtMUJVnfy8KobKz
LZluQ3j5QHXCoXfOPXL/6fqCaBx9yoPhsam3WLmNjtuhGCeG04UaOgpQrptj71VwKS/LT34k+c+O
lbY+llyUeNuYoHhYCtb2oLqGP9qJeFuJxWx88LxB1/rK9yo9pFWl4jQScO1Qvn2cUSm2FjPqDyYs
MXoFIAU+cevlxiP/E8DeYk7pGWLT2KyZ5ooZcq74X3o37IYo4HEKkou4D6hZmEq36z8RTnPJn3lK
11cVSdbAEqW+3x0K1kpYjNkh4XxBe5JdymvMKbhiOFnPBdODA0ZYZndLJqNvuu4zhFCCvUb4NxrO
oPgN5Wg2xruPhcAMk+A/vD0ewmrqoDDEQXDvDfpXXjrcL9XH+GTCsbui9xsADW83wCG1otbISYS/
FR8YGOaos81mBUEqYmG9U98pghR2sY5O3pBv385Hr3r2yIM+xc8bXuEAV8heaRuJakSGmW8TXhiL
ysQQFwxraSF6jI2VRN5Pp2S8HLu9U1oprsFjRe2+3ywpxEA98f1J3K9eWvRtnjZ+5mkxgPYDcUNo
vTYtFUsW4YUulTd0NZKk4czGk7b8EmQ5iolqTjMBLFcFLhdgI8fBjsfXQg6hM7BkL+LjlB5DE3Cr
mYrPexhHtPDfhPRJe5uWGJTaHH6U0THTqnXvXDWZ8gx1LI37i6iwjvE8wAJolBh0eSOdT5zoHsYk
VSFZx0mZKtVSorBjA+OzsV5offDJpudS93gQ41YyxNo3xGaiGTOYx+NgNHD6yh0/z0BfIPJiZSA2
sR7CNkEK2+9esWimOiyxCsBaHbdmkFXeG1RmoJmQ8s5TRq66YEo4OtEa9xOe6XOZHCNH6F7CWBgy
788Or2PLXRMZCk0EIYKwJuxp63zt64Z72C7KHfLnpvRJ76xnqZ3gkSViSTLcV+o6l74gdJDg2m3q
gjTTVuPPccUjkgzlgNur0bUrgCvuWY0YR8pOLTKBwPIoEaGCKcR7xIUPgetncdpDJvXmyOUZxrks
NpoHiKXIKKbPf92AxVkDpuxIP7YRkPzBFORLkDJ2QYtGMl3ZzVk150Bsd5VIDVZtUucMT8z4GvZn
zTlGEzmlR9+I8kJomqAE8f0bLteskGm33w/6ZIvFvH91Gq4W9Fp78qUSV/citcZOaaJWV2UNwmUr
HBWzZPPy6yApLRD+G/zvcZLVNHjc275wuV0FSXYh3Ve+a7Rdc9pr8WDUGBEI7gx+XvbUEHauh5G4
5eNkXg0e/hdCMQpu2RqxpZhg80PG0qmGJBd5bRsbTt/LFg7fwu63z76pJm9f+YJg0xR62AKPwSQh
qPzAORem7Y088QGc/WgCb4WCgLZhUJ6xGy74kQG4QtvSyx9Z1Vau+gIb7J40gS9Yplm/C3Qc0Nhv
1+a90eKaYprLnEtQmK4o2SOFsLPzRlWb54yyWqSM6IBK4Ko6cAaOlaA2MEkl3LvGUvZGIVQl8Tj0
BGZ+v7dmT5JxTG9aLVA0Kd6fyq/uip9f8yBP4wSYaFdB4Rv9gdixtrQnIMxcbQ3LQ20y3/nWPw/X
orVZGiF3Ly+HcSHiUeY7mARP/v93swysn1YM8p4IXUBrOFylxy39ZUbuwYiRL/J7QizLj2ep2YbK
1Fu5J/i/Ny+aE+d9Bu38Ye9LY48TqFviT5tebBJz3uRuRpH7rEuVo/GGtMjwSYH1+VtwSkAXB0Mk
vF9Wk1XfTAaXZmbvvNtbOmcDlvapFNZm3T7rMPJHXSwZ7MM497xLGXgNr0D7VkH387YSq/nmSSeL
M/aktDk7QLh9daEJRkYLpgUfUJe3ex62o12lIujuvlxO0hhmMczBfUMuVXXmAPG6aLN+qY3Re1YO
hXTcqJeqB6hvPMUcolimfvF4V6uq7P5U4Ka3Q7OhYPON7g0Z1GgqQLsh/chJEWVApUV2yA2w89B8
8QjCRoxEueXDXruQai+N2iZi8JAKucE+Z8Oa2zROU1RhJUMY9cxB4AreusfQifMhRrY96qLCvWR+
CJ41Zrbtu0adrM6pO5tuOmAdRz8705dZ8bs0XuS2b/9/n3C1pOgyFNyc50irOgtZvvSyjI76aKBU
dNqEjFnE7XdaX2j+5isc5KbFRAOa1ior83RRjuUfaPgU5AuHss6POYtN9u2ivJgtPKy7/nelarJ5
ds8ErUTczx2X9T8oS0ax2RDnY2ZO+vSVuzNujuAbRtyRUN5p5+MpPvF3bVsbDEP5XnlHEIz7L4Vq
wFsyyL8RifP5eD6yiHKklV08Ypzfc2s9koebGZXsnkbiFXTMrh+1YYPsm4JLaPnIZq942kQg0IC3
TZ7RhcBZqqAml0Fyka91jkiiwMzdYycWy+tgYrZRuxyLUpLqeY7R7D+IWiV2aBA/2YhDWdAOlRs+
wpP1rasXltLAPhKmmkHtTQJwvJIAygeU9nUqU9XloLxBWYixsVLuqjuIjnTcLRHHdyJBny2YJyF+
EHgCg7SNTK2TBZvkrt9UbwDwbAoGhWYc4yRwv22UvapBcel7XN6BzqASH+DSo6V0RBpUxgrfDIRq
jyRPHz9IexMWEsYJ11T3h4/0XVJEjprD2dD/x0SNpDYMPWZVOJg7Xxn+JFx3VI1Z5fj74E7O2NDz
MDgEQEr44ui+eYb1xXZbuF6a311PjrxHSWjgkto0M6bQR8Pb/wPeXf8S+MWxaOPY0IXDK3SEuBIG
16xxeio1AWBMqU3ldH5Uv8uU57oDVFg9Ab82jw+Fdzn0pgexr9tDq1UFZsOtzxvjto/ivnIkEAEw
EL03Mp4RmUKEVaNdI2rIVAForbqOcXzLU36SqGpSkS/XvYIqf7IB49lNV4vD4RrtpsZhj5KtGHUV
cJSL3DITaJkxQr3jNPyFj/ErdYBH59go7C2GWAHWsbd+XcSLE7LxgcDW5AREhcLHuJm9u6r2hR3r
mt2FXTnQryq6xqC5yPNlrObASREVjyFWI5Flar7LR1QkBtr9G3sM31THKsi7KgPkIX6jmU+Z7iGN
vNjnosKL5uNLF6zwOUYyRF7MWbchHR5jUIxlQtVSi1K8jtcnfJNbGr0HlVJaeXmsMAVutgLkCiER
qGeAnSx0I14GFOquobPWs3Qv3DDYgSlI6dMwE9k7G0Tl72k0r2qzZv5jG3jeTi0YFYYgmD+LaUTj
K8/dEZpDevAM6qOMtYLC8ZVwW4Rv4qdZgIG6zyLj1Diehr5zFRDfZjumgdt6lPoRLKqT2aDrtjHc
Mghh2cBzlvQoRgZXoKolgmCR1qYSGdMCyFoirAGGMDKgYfORWittX0/n1LgwaDW9qR9/krJ+h4AH
ytrBICW3+S8kZ25It5iBeGgITrOsWcQ0p0Rk+tHm2s3lkhaRJjAxJZXPW2TokENZ2i+Ye/vwbayt
DxBOmns6jKSXlwQyRTxrIl2VLaHwCDcxqrkc/wpOJtaG3YK7Xl+V3Qv0DO0eWIOiD5F48oYpHrYa
hGEoq8YjgMUGnsxXaJeSofVMBGg9m44VOcZQ/yVYST8IIdI2HTbv/uDz3hoRJU0PxfGZLvmlOGd5
7JPbX8dRGdM64cgmGnd6zGSlwu14ret72ge+Xp00VYrEOZDNiycmeucI+yS6o5vJssCH3yL+T9IP
4zvBkf0zUt+0GAfBaYGFITHmMysBMYfeiFe1oGzi2nA1TNJPhgcLFhUZQk9ju7hRikZDGr+6Hx/8
rZh5U/E7KzeDO2q5/mxCwvWbAqzHWgs/E+h8f3fxpSHkwCGe2lsSHylcTGUiKlivEy/D6ZEbdVmO
ODwFy4xawHpoW+RYOEKgBfMkO2yb8RyzBs8Cs9kGQdtmgplar8iicazRnaFuItpWWUqVxoNXwVtT
Kg2Jc1LdfalHARWIYQfiJjF00nzYkTo980qgo6rvO5q3wGdTgqP+YDea4doqQM1AjJF61v3i/iyO
2FRNim5tDiXH2hCtWLHplW+gbHaJpj1qqpHPnoEIePGKbyjJSiqT0QYXLdcU5GPzSlwY1hfufASg
VuvZTnUj2+VEjwTulo8tqzoLVI3VIW3MfybeI/sZPTZW5Y6LSLl5pdh7r+0SesIlEEdb8t5041ya
/hyWVyymAAFyg6YG2hBmpqXyLXqmEEPtH0IHWc31Kv3qRuaL7kqywXHBAu7WSfErKWczod9eUkMi
k1gNczxOl9YqEiStGvbXbNdl59ZeLGwvNPtyrIDjS6PEvnrie132fbqsTrz1mDRz+l8oMyQIjiDJ
9CGSVZh0bef4taS6F1cAnVfVrwjTjgbq8tVKS2FqmeBRidwvRjCCm0uG7zCdrHE/xvA+updiWADR
gxVJEOZFtr2BGDtVvJEi6X2FJxOAM4aa+X2dT+oSrXPw/qs47m+thX97bxdGD2OjOQ7w5cExVbwg
v/11+3oY3XoEN77CtMNao0iaKOsPs3Ccmw+v8I4m//84ojcR0LQH1wOEeCgdI76cVorg9Oydqz4G
9rwEwjfg7NJwSTs+K3yooKq6gPoCgs9m6IwYMvSzKX3ehabs44xlbnbYwsgW2hOz9Ljrrb0NiHvu
LBeCseWMuvzE42VhyCRUUfZO9dDXVx1LMbVdEoT3VLuuvdyPLXmWOjlqJ3W+rWY0yAwE5ndEiFYn
k0Mq9cEAkBwVYRbAIwqyrYZ3A3ytHVaUf5znYwc6sjOaFgdulUiZV3kjEzJD38lu/k9AAkY3E7Ja
UiSFcuggGp4aW/iaiITBHb8s29lS9RPnQUlipfaLk1RJT3loYJF0BvQiU5OjWBTxOOVj8SR5agJZ
NKydvqfPkT/K4CwiBu9bP8wnAUlZSE9PV2oXaPbYuWZ08jPYBXY6cGtOpFw370X9zlK9daH15m8f
JGF7IuAqm6Lqp16Ulfz4pvvnTEc/O8ePrHV7lw2f9gQ7K1HlXkABefcM4rCiFb+QslvNA2+n+EXv
85STNRusuXhm2pclyJUVWl7B2+aIVvOAJNFf5McxSEWcsAU4Ublpks5TUYCMxuaf+NaNNO2neqOP
Pw30JzdgsaU7MdoahY1ifr7lU4dysBAG/Q3S8lVS/sC8pGNV5miDBmURrduXHfLNkZIrZx+f5UES
LSuHisl7ggbtlnBdQCeLBFVCDQywMvE2KPMpedXNp/sBEd4pH6ayeHK5LcVnpU7uV9DrGRW4BMdG
zlAOYlTqelou5e47miXkJgiDHt6iUWf36D5oUrCb0Wrqf4iDkW+KOrqiFaIg00Zmf90ARupk+Y2V
WvVFdARKT3Etwrb4iQR2VmC1xudfP9sxn36sxUI4DxmOt0zIAX8HTwTB4O7mQa4YzQPy+93UK58w
kSb5QE4JiTQ7I+HFd/DKVtwzmb0+x8X/VMwc2xXVbrrBTPl+BRI9lZ3d4ehYa72sw7EE7wKeYzY0
d6dLhk1/CubXY4/kQhzRmhWqgaPr8t+tCJZNoo0QO0Krlx1MGFSYy9VWz9e4p5/RDrPXemRskiHj
URTkxr6v8zpR/iDPdZHJ+dwIEP4Kri1FpIfVtQiiCuWeVU/ukOPJlQkbbzP23E9SP7hx5k//6Ghq
GwkO6PNSBGIMoTY518mbnFCkPEuRG4QOE7+3NN0aiJkndR2qt90Er/rhvRaXLqSzUzpEqpaA3gNK
ZMkjIxUkHxXkxNEJMf37oW8KjeIGM0EB6lZb71PqmeNEZ+gd1Tu8MniPnNnNHlDc3/XFCarebQnr
DEQdhTIjRiN1FYb+ZNAqNZ5cUF+jIIcdJ1Eqsk6CLwWEPpso+fAxYG6yWLF/x8h+NggpQMn99/qt
1fYEh1WyZ9U16rQRUojizqTlPbnhYGNZZQkDZ5XawQ1EmKQgzZSht2iEZ53fzXM+JFGMIvwx5FND
6SoXHLpWWa9+rubSTuyGsVb5QtpStyujtGegGGtA+JLSs7jNOqEHhwurnL9fIiVrsnsjbNDGn0eP
CrQoULdJ3uFZO4Y73gZ9mk5tZ6YXe4MraXHAt5SQMlbp8lAsSJEBmL5y3Awy3fBoyPhBSDlosjf7
vZBTtda56Oq+VJ3WhDtKf0ISnxyfEprAhB7n/4/issl643pgn6D6NT4Cf+dMBIueNEjOEU82KZJJ
jnBqsy0Gi4l+6YqoIq7GnuZp+sWXZyHnBT9Qa8kxtm0rQl2zI+zKWaLpfmxPU+LLDw5NuK9ybRZK
DrCSC6fp/syzURSX4RoI7ghe3iUAj/yyNuZ4tY3SXoFBvlOFqJmU4oI1A2HmSiHYDvjwJ53AjD+K
Ou4eL26rXZlsc9eoOjzHFmPuHavw5NiA4Y5JIyQwXQF01n0wFAHzhrBkGxNoWRGaId2Hq+OtI6dh
udIzeCdwtkjRFh+ESrtwSNKS1YNav496fl/VBClarHCBVd02dQB+Sdr60/iWTyaLlgm+WxhK6dFj
3qcNNsmTbeIj62U/j0M2nOZdlxUp8eBDWiI8sVRLJ6wgDlICTa+Qqtu0lmkOV4AwexjhwqVsDSeP
/3AJ37ybYKilJ98enSXPQzhbkV+jc63mkWwr6cDC7fOBpcUQpTtWjzetEVZ7Le3z3Lfkq+kHuwZx
oOueKFdpytO7b5DQo1JTKuIusAzD+BiMHmyVbma7UG8jRU/qeJ0IvFCOC0hUDKOmBdDonPOGxKD5
nBp904/X9xLAnfCT/MbSCIRb2mXZ6g3kexPntEcJjVSiSOEWrcJGbPBqxVZLQc6iGmX5pp9PE2g9
a7NQazbDc2R5sJAMlViYjxLzagCj9vxly20eIBWQUSGhw7dfEWBECNMp8e2MPw79H/WB2Ek7M3wI
aPvJkflUlTQ6OyprLC0k2NygAgaH5qaf5TEkdT5OFdMxR0nh5Yj3GP67w0+c9uPW9eBf/4QGueXF
Pj8AVRJttALGb3W7HqL5nIKnLqNdOKUjBR0bOI+AM7IWQRf2TLSbLahSm18XUH6zC620oq4fMwF1
/mVP5ezePGqE/bi1oSkvKFG3n+gagsRyFhu3izykQamYaABPmB6zgaC3mFtudukebQlTX9UmzTKU
nLMvW2c2Pbmp6wyY04cR5slBsYohMJz/LezAqWg/3nUEWhb5oZLVgr0IWfnXouFC8f3HzcDnNmHG
ucVT0E8RXQN4KreBBz5bzLs8mpiyxJgA9TGw6KXYx44ZteHgwteVoR4uzfO0b3kWQSVkaRbCO8YX
iDK3/ZwBeCex771WuT4GMQe43xM89pLLIMwTqomelIpW2lkbcEiEzZvZbeREvLi8KWOCkZfWXo64
KBIhN22Kaz3XDq1GOB0vfvm3Qj6Ssqf83Cs/bGNsjE46EQg81lwZ/HeIee/sjBdZCJ/7gdzI51x2
QTBnZDSx31HxccD/mw0n6dKgFP+0igsvQ7P1tMSxT6dl0yTtfLZpEB5zUGJbhyLgsNQ4F2qnlTea
ryIgVc7/vXGps2d3juUX0xrKph7ZhQcy5NfBboKK4EnQ+xa591tUHuCNmNTix2RSZaa9zMEsGeZ4
S/oRm84dFZUvYNxDgU+OJwWyG9zrVa6s4keK8MaVvvLzKDT6a7gLOHt1Bv5wftI6ae59tYDMblNg
mJ7tzy2oSfx9gP4uy/QFsXDpd6BH5m6CCbKQvp8BhhA7y+tizfXXUqdVSDcf52EFmeocC2RIwGA4
atH/izqdroequ/1G9uUPPsLRa4OV7KaY1Pb8lHLLk7BhBVUKB3MZeNFSKM4Bq5I7Z6QXElg5z7FA
TtoOpT2+2Vk4s4lbrJzEASyQwI4dwhk5SzraVxfKv3pCvqLzVn4wvUOoisOsIpWNsTaksM6zbW0x
yyqOnqNuFFHq4BC9wMoxiYSpR+QCWurVAoAiGhvv030NwmDExq2TMPO4DF6jbIIsdkwUTZMrRZcK
dCQs8RPR4ImGv4R/lIQ=
`pragma protect end_protected
