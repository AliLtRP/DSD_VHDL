// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Q1wuXCSBUG0TfGFNMH6mHW8pNoovwD5cq9PsRh2JApjCVo6CbOyE2Ft6tHFem/x9IAxoW/zXLOrk
/jicoL7xV9hQsSADmKYDEPBxSiW1+rV2O/BAjLBzHrEYyDiVaiTTSBSC8pAnFLyD1kA+exfkOHq2
Qs9kDDNVVNUPS9EPEJ6LSh1dsPZYURL9NykPD1ZlW6S7zxJF5ppHOLVQqOkKVKeMnTOa2X+VLYVb
BmOuLPZaIWzBJFBrejx23lzBnQRAN3Bu6Vuc9JbdmJqZHX+U8msuA7N95vQtSv2MgHUplPcJCIkm
vFXffB84pzJACo/yj5+hL1rWWkOLGW7VPqvrKw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
YUEEQB8yFRByiVs75r85KROsG3ilaf+5NePkW8q4ATnZi+ZgRjaL39v22ur9Utuso3nnRlMONWMj
QqxU6vQSZo5jraYmFcPYxxNs76XRnA+Pd7i26yRM/65eTcFD45jx0CFvrQ8AkpGKozZuOHRhITaq
zajoZefXIDNIrlotn7dm64VzZAoll8F36jK4xoxssvUxnjA/NPO3jzuf1bQotdt9g6ZYSlj3SzZL
c9Olq5YUy89MY/FMco9rC3QJsZuzmC+WR99VzsczFX8AIn0NAnT85/A5zRCBesdkNOD8ShEPY/CB
VZ/+kGgsP4fAOQhVgY3z5XUXFWgnt1QACbyicu9AMKxPKF8hB9tPiqcqw6dUKDpGwwEIOpM4awxt
pFwn5E3DWUi2WRJM541Tlnp+mjS549oOK8VfenzOwcwrlVvlkjbfP4jj0AQ6seH6523IJhpep3J7
roOV1o6cMm/XG2NNWc6UILsbQk7TwP2wKZpV9eGCZ0vLL1/jgBqWi8N9juFhqjcNSQ2pGWS/XsQV
i6vFG3nRriLzK0kc+MC8RsXSLbftz70CQNkegWfdr1/QLnJLwWEj6UotUxfjoZZPCXDAB9ZP3BEi
08hNnoYgXsSWklA10F/TvlkS+BNNTAISaEDxbV4yuyhFPTR6VAi9jXtkMJJK8HsPkTqD9Dg/6kzA
24kUCXVgeFtCl0eHnwLgD0Lap+spXf2kslWEWcBhI+IyIpu3AE/DOVJPynOcpOylF2sQkFQEW9SW
gutyy/qlXIs6UMeXdejy4y6/7/wgINZ+J0YAND+zNEJl8gyN6ND+F3occKDritnECSj231GzIyiX
4yJcWXMbJX7HDqoCx/xLHDDGsKIUT3k3FElmJv0iQuCVvwmlUI1hc2zuapTDOAq7OAr2AvclMhlc
HKylH2RG+8NQcShISscC8D6q5RfwUKio96/adSjZ/tY99q+SgF7gEC+8lJ1vnenn/zUhjd/BHK6W
G3AKwLhhPwMrvAPJQkvJNL/3fMi7KtxCfGiEDZiLyfvJR7ed40ipZG+Dly4qogiVv7zXPGNo/IMv
YN1Xb5yAA37bEcVUO/OtDzmvgile4SlS5GLV+mxySm+8iqXRdqyaOFCTyuQ6R/QPHPz8nQ3sAEy7
9oDd+N6NqjJi1tJ/yXibcQSuwACjjCb1szg7gf+lISqaikFFI/oP0wESEbLkBjgA5KwqcPyM8iOz
ESIsacoHZzF8XiTVVw3lGu8x2hLccLxa5Oe/d366T2qDLhJ1/HtsZC25X6szrua87CFV7ODCHHz1
4tvaVFM1q4IOh32DOOoS4+c9Pi0TX8l7PNV7373UJqPMy3pDQ61GOGyI4FdFq1IAyB5kM49GTXv1
1SVwbo3K1ybqEfD5Qq7ICd3vfuhJeZDqWrumbEdVmZec/ShnyWkCDidRwQhOMNU/tvw9oFDeNq8e
QtBL26fL2qz51vK+yYuz+QrB8bVXFtX+eSwzcncfiHc9B9GKItY8y8A9itnfaWvmiJ7Iq5JDZVfd
20SD1co5ajfAbY5M65TiFjqqs8HbDaSJyQZfh3XLP31l0YI2y36UtLqi+ezp9C7ZQqptXgJrUPXn
rbyRLhUXK8WvQkYZrMWDDz8TEDauEQ6UPkDyR2EwTtdB9m4iRza0VYEcf8sJ/lnUXArRFRrtFVbs
zwRF3BnYa+aSUxM1tAWphkYtKN5zL1V36NJnlqHrN8gG/6LS928cxt5hya7eUHb1Lc6PJZ5GmW1f
0V0+C0Sdyv6LKrja/M6qlj2bkBzo72FO7n2zsep1FjRfWlOixn4aZ1CniWuzPRu2i7JOTGalz5kG
IIFsoiaHhHzwF7VFb8E3zMxUE+f0KGZnGxdaeDTC8h+bEYB9jRFDOp/rwFgsMG4X6Em4uZOBMz6K
nAezJ69wdYJxwfS48TK0WDfe1QzlSNoiY4fw2DXov74O8fP98mY2PsZiPpjD5Qp0+6XAr+ukrLSg
3duW+ZSAbKBWaehq87RaTK/8ZkXARn8Tly6NQUYV5KPL7Y/vcLBgws4uG+5kju0Obt10yL/kxpol
OMhOuoGp8FX2YEOepeSJ3tzZK+0uhF/CDSAjN2f44Pldzd2LJBpXTlzTwzaH7SqXktqOKnwXWrXj
krV72qP9wkvJpV6p5kMXgnjsrZ5EO/6uxnx68OUKWPK0CTC16PSu21Y9aLd4dbC8eD4w08OY4fUr
RUa3T3QXID3gX0shBoqbtwKC3afVFM5++TnHjedH+IYZS8MO61OEaIJC1Jq5yvYieqq0lCoMoJ4D
a3g4LQcNKSWHF6hsGChfoGS7U7tW/Rn5hD/O318x/hnldWGQsIvADjDv0NA/tcyhexW08jFxAM/T
ncVb79/dkd07jbr+fYqw1m1z5Q/OZ56K5+8yQ0aoDXHxKxq7OF8Hl4ntEbnYzgm7bcQNMcp0jNdu
VKdIXmoAkEbNaWs0nHWdN65xQXw3A2izsx8CK1cb5v/bjEsW9wz7ETI/aL0KX7wheH8qI9xkO/pq
Nu7zKN8QSPtNX7NVOw4/M+N5SVh8O10yUFUT/n/T2sK+RrymQCn03A87i9vijvSMZaCN30sfbKjj
cV0QXC56KuCK1wStVQt+85wOzZMOUOgi1IaLwkbN6ORxQ4d63Go1lVeh4tZazxqEhyl9PBGoIVXn
wc4yQhKVSPHMBM7tZQaj5gjkifCwRJSC11v+usfTfIcNeKskAQ9hXHs1Smw0dk72ZBbfQrpQh+v8
XdXyMooEo8vtiuWDvrLY8gd3GBbwNlw6t46imMLJa7fGOi93e/8kLAmyp6z+fqGKNKgrNjr4Pq+C
5iv6BtqSVDz93MccgJdyjdkk9MJU4EOLD0S8hrRmqFoG6YCmrTqif8bY7MFjD2o0mry671HvzKtL
35NLLjQGFjpSJd146Hakp/BQHEePKxtvs34EML/qoaHG2rsRax9unx18/eZRusk73ppVoRFeUsZ4
hHhvd4EmGbKeJRP7rW/Vgi9wJgu4Ibo6zN0GkNKI0qDuYIOrrN5n7Q7Dz22cTeNJRzMHAglGvob/
zzpXkQuQJMvsZiY3FmS6qLjU3vTHIZL/6VSBwd4tDtr/mgpUGueRqAD2sjXh9RKY5++azxKN3QSg
GsSdrwx/uH7E5BYeuWy1k0ZvUoGRhLOdLRFJutz5vHZ0dW+1UF4G/aJTMjo2dqHBcZy8Lp3oMfEE
QclcSMxQbkNtYF++kMMzZ+sgCHVkMm/M+LjpR009QjVASSdvuav4itUHeApVvLq7QB42ReiXGtkZ
glk+zyweQhUU3iur6DnC0+SejrqSk4BO4XYadse8Xazx2outNE/6s73lKUPKtBI8njYvtKwhJYqi
rFoFVDixbQ3Q7zS2984mIAJF+nbs5L2RiI0U77pmdmCQMEQSa1DNhsvUDxKZK+3ahSaiCpUIoO4j
wGzsML7s40QzMlJfaMrwZ/98TAIji6oAbDUbXjecSfjPT6k3OFkq0wVLNFIPbqZ5n1aBvoU39MVF
ZwdtaJXwRe337LoP229pTyvMsCIYy+nPHT7aauJvOXR5WB865scyoX6nEpSzKniY6THLJnUu4J/n
n4XeeLHI9JaKx77KLUnsTDWAt0C27qtwh3fj4taOUseyj1pzDE3yvtEVHjypWZadbMyz3GgG+nIG
ERRkXqwZSX3V/khLqJc8GaJIFGXE4vROYgrnda+V0fA/JNB+H8GsyRfyBX8b2WS3yVgmeLqRkfUg
QwXQVqgLSPPEWQjk+tYc13b1CbPdo01N3zPQdmbZ8uYYJZOQwjCd4VSJNCeaQ9UXqkWhI56hiNIN
FXYSdaxEXNq7ec89RGckYzSR5mLBroEBbnJSIQEwN47oYT9ci/attsM8a+ZMOFLPUk+r8U3REMM0
/Nq1sF2D6/RLB03BvsGmF1Tt7/50IQx7NeNcL8vYnVWdGQBow+vw5FokIS6avykJc0tyvx7ZUT4Z
GUHNfVnaQQUBLfmwZW3xLA5hvW6s5aLY4w+XqO7L57AIX50Bhdw9eUYfpYhKIaXRPJy/nKjLuCsa
wnxGur0CrnEmeJpgDllQDXyRVZK+bKRN69m/HI1gYk39g9ybTZrB2SKyxnGqjVNtTQxfQ+TppIZs
VrTNtT+9sKFzaZdhhL8j9+1rCjkZMB+cgHAFjj58+fsnjJVoXaxe5FYrUMkBwG8B3RxYpQp9Bsv6
ixsd02eqLWfMPpvJodL99JGQwGySQ2ifitkYmZN2Z89wbr1+42AQ+aQ6v6GQtCkQpvaJGgPhDZYZ
cgop04k/4iyxsyrghbSwV5ZYlks5VrnIaB4sqERusZh6yDFVplh8uip69PsgFxYrUt+Oz2iDE7P1
TUhiadJLQBCQ/K+AmXL2ptLkIAAjQFgEQmnbgFkqxTP1YXPpp0LCxCB5rH9lFYJ1A3g5fQJ5jnfG
ueH52/B4j56yeRitkwnWbbJdSmE5EXiKCgX+IrGuehFcBWVr+pZOAV0laDYBj1RpUtzAakI9pYs/
3kiEa6oDvns+7ui3TjIqIIExGZS87kX7B6DOTX9Fc8HIBZwnfcRzis74iNXpBspru5tEobkkEYsV
5Jyc7O1yK1rMkDFng+CEvfC0NpdrGq1srqYDox5JPA/csFEBtGcChyIDrp7UiTCC2I6yT37DlZ4p
6ekGdubfmh9kXEet9zeSZMRjQlYIxTHEYdvyYNIVDRg9bfgbI5QaxC7Va+LLu+eMecXQjSMrIqnB
ouzrigjFETQhB11DkQmyAi5eyOWe0JS8RIvJRrCaNFIj0mpRrSz9IQbfNozduLb7DYfPP2DbBdOT
b1yClfUr3/Mmmr7b4/3wU+icRp9SQBce1GSjU2X/eXKK4/ZhNUnBxhMLsUuSmvIEFcB4PijMY9RH
RCZd3E7LWvmmtohnN3OjTnIqWJMcsk2DnGCwgtqGRCE60CNv4AWyQ7605AE5TUhN1KlePNGksi0i
s32CHTQWVEmPDs+WMNXY2DJtnszysmREJP1X1LxEbx2b6iTmFl4NhRKzdjhX9dhNpt9iL9fTd3Mj
ET8hbSWX51wEt2m/E/Xg3uogxFnRaYMLPrNsfTivs/A4akPUx7A3mtSjFMApbplEKWalSqOCt2rA
kAIzTw32xeDeHl6tO8tJ2InL4cDxg278UtABU8xujR39R/1oDoJeL7sEUQ+2Kk+YyQd3xuLYlmlT
LaiCQAN/gAvtMUcmLI4+BbL1KjXs92u/DLfi9D88T43F6xFRgKkZOJuJga6Nhk2XO717aRzYCIdE
iK7u7qbd5hC69ZatFREx4JQJ08COcU3STBb6RHWGvoAkcP+V1uyYxgi4jayLPdAVhOEDrb2CBI6v
J5L/t1KDWD7Ma8EmC29yM9uB7kVZiBwLw0Me0gFZsKjWGS43LPDYvgFET7EEs3PfcretdaDXFOxJ
Akmh6U34kLK834f7Dzmar1JAetu72+mdJm1eLLBvY6OtBpAJClMj6tTxXz8S7ZIos5TwZXcoZuNV
KcsSLZ4LnKa+F1NiGXG+h+UKGj3nS1E7Jmirk/MHePyX7ROUBs/t8GqkJaIuuSRcM9VfuzekSVVG
wyIPF5J6ucYVYKxHuSuatn5QDr3EypeozL04k9f6UN9ZeiGHwZNBsxwfCmkg5xrlu16cVTY1auXP
xUuCstthk8+8NStJ4RDQ3Ah1tUUet4Qj7S3xQFDPWgpS7/jIbXNXlyhv7wVkT3eSJpskzplS1U2z
l4usLUSxltD5NiMku0oVkMTkvRmf6G4Y00+zY7j81gF0t6hXFRqDe1UEauv3y0btj6uZvDrWtQFL
hz2SZ9QiOHsDBcRMBk7VGckVtia5QGEifa1AwExeOFm43Z9G0Msj/JwgTzitfKc4rQfP7oCDP49D
jR5L3Nx8z1YRlm/8kC9Q9/IwAryYo6QD51OHCYwD9iwmXe7lLPdd7gRH4njBt4Pe1yIkGIPUyiyc
x7G7SQ/fRxNDd0qihNRhdHJBNU8qZcTZsyM5MnjzsnILcY6LW3q83d6N7F1aBX1QD7W/YM0gdJuo
9sO2+18QRQxUXgCCRp121USb3hUhx7NbapLp/9IUCY0pExnlQ6BNLTPpD4nzKER9ayAmH+fxI5rk
OyWPcVN64y/J7/BaarqxHb+zGkqnGy0A+ccirgu0CvgcTFr7papiS9aL1PpKKgPxtCiJ4FW+iVQP
kfKaYLh/p6TCFiOFNpn3xbOz384NJnGsCTxk/JAtsM+EPkrkNcMfKHdFl/4kQINo15W7G+QjdJx2
5Lf9Q6Kd8peHzdgiB1q3FRX0zGWMcXMNELs97Mqch/z3YrNNOgF4TzcMEDn8mNoiD1PKEIZPflez
q9e7PzXB5YTUkKPynQiCeoen4ueQrB+fv3JbzcNdxB8wf6e86JEZ78X1AgvPpf6HQ8fYJqjCkDwL
PMswAvrZnDfQHFTijrcX5LG2Ifd5GBoBluxM2EgVH8kr25CZs/xh7ZZoD7hc5Wlp9Su3gmVgbz4+
GbaHYCmdZW1ysMoLB1+7YzA3jRRrcW4EavLScLR9Cs3mJto+oLf5XD6P5gL/wFcJZzVb0TJW6zix
+ZlBbwC9aPUTYkUv2vk/kk4Jc1zWyLiRhPZZesN+RJzpQQD6jcN5ip2QluPdQ9PJ336kXibpJs6o
im6vYWy1OtCXqloow1dr3s/Ullmgyc6UXMP6NedLidpkrS6WxK7M7VodoSYsTOGA+Ysqb6VJ7t5+
1wXUNKTFT8LDQL4XgQSIgasII0R2Cj3MrrUtoQwwCM+sxwwKoNaiodNFPM3PgvLvaBwQf5hRVvrx
iz+1jVKOqfC45tLJDv/VbVel/6qxxugRLJkGGkGFgaSHeIWEJSjQuJK/XnGEjapFlaBr7pk9IRcC
IPNGScTpf3cOQ8kt0mx9tQApH9Bq03dZs76n4lPguxleIVm3n8+2v+vfd++dzqNKCLAmXsvRN3Yl
QmcMK3wGMvxe1vG8KR2et17NhKTk+blsSYRG5mIW7GdEbkFHBqISAJN/mBXVp+o4kVZ9t20RLd/3
TqHCUwrW86Z/phQ9xD8PXCKNwonqtzlKZ27rsdCBash0PsIcYS2NSs2+31gR4JOlSU3bLSRznskR
RERvroYFM5rpIUJX16n+VB8nRhSR5iuXmaM3rHAyaeJtvOERru1hg0xk7eJkcy8/GvYN1tuFdZwJ
b+sek/xRHSBMlUtfUTT3Ha4iLj9GZ5u9Ax1Qjdwxd9VHTlN8C2e2uwxrYnHQ+fY+4erNpFv8QdsB
raemyZ55RLwP5Ve+WbFuCYP/p7ufYvwNrT8W3o7U/rpVEMtXU/8lkxa07z1NYMvSxa/XxrD/2rTe
fmCJ5K+N9Hs4FGX+KK3O49gBHXyr2N1tNfPPkaytgbWstwP1uAXyD0mGYkLcDgbrPyhrniOqMJ3S
ittVn7eccIAcTnkaiKbbvbiigJN0BeSVnAR9CjMBqA9CH54zude7a0KSOxgjhuJMtx6B3mOD/TiZ
7Tk4DktlYixQrd7zdVn7kLiFtmemUFgXsgrC9C5cXEMfneeSE+4kn0vypAQNQHuFsLCP38JdT5Di
E4SNUDBGcIRoCKhvsLLGD3kQvP+dZQfdDMKwHDN1T4H6G2KYXTjwRxPidaG2D1OAt8Ph9D7gFjDV
P/3KJjGG/Px98R57d6fyfjtREHf2zkAi2hCNsIX3belHFxzr7iXKbVwxakkC2AT2Co7GiAAX8aGW
uoxZjaHJrOO38NR98O9iQ6qsJs40CoL4rmcygbOYHPbycQoDqWbyCQGWFHC0Kzb4LlenBbTTBfOG
9ByftOcGbS3A+qYuptDNqSwi8H6+zEEuAWK23W3PdeHNsFZzd+02tVh6kky+kjYtKKEJM0WhncWp
BzNVULstOpASGLUvElVVvdlD1gSO+M1WHVIGKtohrVHtC6ACEc05sAadZRIf4yHCi1ku2SPyU2nb
eu+DDbHJgoSwN4lyTDnbYd7d11Bvt6d0vUMKw0vqmy5ckWcWJCLQCIkYrZEvRCt5m4WSo3LjXxWm
0hxZIr2H2BQOVE69FT/PVysE7K2Z7LP9NOo+WD0vF8Sps66azan8f58c2Vjfz7o41Bh737EHXuf7
Qh0P6+JOMmFhCe0rwDLYfGZM/iXcQDw6BUgMrPvf5HX2Ly0tqx1VlvT887KyOsDhOXL0pmmLZ5lU
9/NRfH6MNNFW4HXlLKEKuSFaL/48jZa9q6z89TeWQ2ES4gFCmTjepxwOQ2t0j0dkk/1Vs9m6/Rw8
SbvPn6EolZNBmrUf1kpWeqHi4+KE+qp/ErQwR2uMnHSedylFhBNEUhNGL2qC01uTkfUEy6+0ZrLd
2OS806nSHxgnL7d7bsb+Q22zwPOL/m+A3dhNpf1To5yDfzGcfoQ+G0PU54RauXQ8+HU380x9zsD/
NGRt3X6CS53l0KuvYvhxSc3TPba/Tjjo0F4RHFWKeqGikEA+WF6GWFQ599znwKU1H1mvGtaR6Gf2
uAcoNm1QqHDgC0Fr8q+l8ByAMYzGbRIXhVPFD3n2+RLAatMRum5ZqkLUEsDtzQn3uKF/OB9kxklp
HPuYN8SF6V9OzKlVyRnfGDHLcEFummhY1Z+Q7KeQOogubdIMyph3UE2SNAG3TL7OaaFZzNZu9UmA
q2AdBMQ8U5POBtW4RIZqGHOYS3Abx3W5a2CFG4qMPknqN1IbY6Cteky5RV+haTAFN39Umq7YsVSj
fbA8sA90aQP29QrBdwFprchOvulWBAPfMOErHAN75MAQY6UvfAeibJ59GwY/nepJKKOwYjW9cq6z
kA4qubo9Xqt9VAGIqBU8Spd8nIIFUG/yYRhc7ferhu0UOD38Ieb0Qr4KzTuFF8fQ3etQL0TXhx5Y
IYQtqIYy4T43dnRusimljUU63KxBCPelA9zi4LN4s/3wQJ5+x0hMlCgWyPpp8ZtDe7bV2FP44B/+
R5TtKrTwJqKT020zHsz/+TjOit4TuiEPYod4BzDOzGYqvaa4Q3pbIm1+EgBS02x/w+IZk/403EAx
b9C1fkNbuBTvvaPJbIy46Fhrf3ldwJ74h/CHZn2W2yk81NKSVrjWWgQ6qcWsEqAtTj2nzzv9EQSi
+5hLEfuB0pqj24OCtiCNue1WUhCE6ZQ1UndfH3VkxsY1L2VkGzxatYN2ZxpD6nzwmR7+Wieq7RAj
UDB8Blt47c8DhYTWR7D99iMDcbwFjTsv4CW9Bdtn+ccSKKFC3LjMpkCszdPqOG8ucE0IrnqFLOpl
qUy6nZunhowNwmUxgzXFkB8B0QYwIZ80oY3XPqk3L3L9Mc+C29A4imPd/fM3jXJkj3tXQxC1MzUF
RgI7W/nixMDl1kLnXy2iZVZJJOaYxWDmrx9YVkffermSP23E27C3qJzAZLdWvkHXux6G0Bn42BOs
TP679+waCtfXYP3sNVIqK9mxzmrWgjQkOhfjO4drJCoGHto/kuoTRw05uQB62M3RNcxxyRQPIEQv
22K/dUmv7sSEFbsHwKlqfP0FYDXaQyvi5kdY9M+Kbu3njqgrCK8bfNs4sA/rkMPsQBI/0seheNzf
sn5s1c3tnApFd/um1NTcDGDvrmrcb/N+CTGqiXhMZ8NfVnI+NpkhA758vzFFU+XikOktxPX3W8F3
Wba0zakb7y2YK7hK9TrHfUKGQER1Ldd/YhGQ/fY5TWAA004dJUA96ifMEhP6u0ZosRUMRsGDJxGm
TQaKjqhYLdlIjozhe9axnrHzNNUpKwi05upKZylAC/oyfTIbBI1hfmsYxjIE1yPSkqDVGXMOnGe5
U0nOP8JPCjWIMoTtgQ9jZDn+jnPURACqOUOh0EwCEYmxnlCHmt8iHBMX4reL0ORnS+//7lGekH/S
QYzzeehPCB7uhbjLgfXp8YL1PJCY630dH0EzDIiYS5ehSOkJlXQC54riSjWCmUjp1Gy+hNAzdvkN
rluXqTr3UKxrsRLmRY6SaM/NO2g2vHuqtuXsx1swcfTNTTtULrCxVMr4moWBQ/TNMLi+rmh/O1PL
U7g+dFeuiaep0CT2flfTXrdX4FukHweYSBkJE/8x0vZXEda1/JhZO6c2za3ZCnZ47cjUnLHqnmst
NGUyUohrPvK3yTRRYfl5l8XPN5fEGQPTTrg4Db58QfhxzJVZGoLWH7IDBhbxafCCyS7mQaOCP5gw
aCyI9YOg2B+pcZer29DrPohKhz7DXGdmrfVdD69fkR+qUZar0F+0ND5hKUjxH3aNYQzn25oRUNKB
O1bKsH+aIJvCPhmFVQRT71E98RfJ2Wg53OHk5HTkUyamT89OjfK56s+RC6jBNyUSKEOfKtwzsewp
/vtzi+zYLODmTIZVw6Q0Nk6RqiRIpJb15uE2sH2Wbt3xzXE4SbvJ4Ey/lndC1bi341kLdmFZKL3H
S/PDRJ5SwDnC9vIbYvRtG+ASL156XnSzxWREf5G8O/ra2QHWeBn6PxS+jbZPOPpTTNkQvZP2KDls
IuFuE/ZfI1hvqooFO4HNsrDPsQdk/TI2gCvDbU2fMwk9IiNmpcekvot1h3Cys+aDQcLBZHNMpfbE
MbWhjenODt0MIrOoACaS4rwz3ZObQTHOVqtpjXR7vnjlESBdEz3ldbJ24nTpLkJHA+rqk1S3X1Vh
7biJwN7kjGAC8wwd4PxQ3put1K87oBJzGmA8rbzabELs5t4qVoTf+Dfl11IfLFJG9OhkG0EGLfkc
kqCRAp6QDxsjwdHhlw52R59cuF9eFphaPxmPo+BKg7VB6nLLZdylF9DiPNOQUbat5soDB9Wttyt6
T8QUpIn0yyAdFDKf1s0FDhyU+ASwqIY+a+lw6i0c70HPdXV/xzL4wknvimYyMMgvaQ/D4yIKJW0H
1i61gqVXXtYQGsax63eGLV8aEKtFbISI2dsvw+ijZ2LZ92uq35ZMo9IzcFYhGWHbVP7Wl/7rOKz/
7m2Vp25z1837J69g1UnMq45vUbAgCoQwt+36CkRbwxy9BdwjrAD1UK8KwxueX5nrXaMT+1+aFeWA
mQwkneFGqyFjGaPudaujRpWvR2QO5LBgPCJSuRQfkJTu2mNbDZjpV/+DUUKpEQBGG//rQ2+hroCn
iucsLy5Y/Lb8pRlWD4bdtM0KfOvRnK/Q3L85IGn/slYhKMoDdBf3Rzl7Lmm0rQqbIp6m+sCJ3dYa
Hekq2ajM5ZC5w55ybgn/PRuzs8ukFJbFHMFUr4bKntLIPqt2DUcmG+l2LbIaDQseAXDoeCPEokgC
GtzYtWl1/4P3rUnT72DTPrayufT9j9iivsGeknbloNdiEmO3HxNnF+hDn12UguW9bzZeUHUF9AEV
6YPb2OCX4eoMn2A+WxvAuq+MUtbdNtzghwLHpi6logkDUcMSo58hWZigBY+LWxJORnyBkYt/70dJ
DLS0hLytnHyagZ3a1Pz7HSYVgfa7KxasEPDanlcTYl1UaHiz6Cz3pkgltHMaZY0HUyeBZgx8RztK
gX9GF66/E65/vd9Qv5IpeDDoBf2LPpGP7lIbwC0uSByPhlZdqHkt6l0+iQc3Sw4neYlQ9BCAuyx5
wMDiAULrXKyqBLnp8VhQFAjxNYBXjbteeCLjGM1URER4fHweWaKEZCvwYgad3iSUdD7Jnb1wBsLa
cKMHlgLb4C828iUNomqFqqIN7S8NDm0aG2avdUqw9LYHNOVzGCAYPEJUHqHyiNidBydxXZjzAjS7
q9pvAX0OEmYHyVe3DSu1dYgEEuuFnW7+9imDlXvziBpqHPIcgKyI+o2GFwdL3qksaqpH3GVUthUP
XzfCJqFWhqPAUYPhTD7WB8NTUKfoWeTWTsXyKzH6ssvujh9ldhlVs1E+W5eXZ2pKI5QP214ePJoL
3bExEXTN2/pipA/pdDvtA+UNOlLm125VyHiVp1HRYpOfvC33kUgYouF/pP57Fpev4geTigIZD77V
Ww3rIxGgMBpSVut2wUmxskQEfR9oIbUPjQ9OUkXow6r/tN8K7t4P8xVkciZnxNmXB2is4cSa34cq
MyXJvCot/Y+Q8zCnkaW+yHaXhK/1KBlmV046ys6W4QvZilYKTCVeobdRPIaJ0S5StME8ZkcM3Dgx
zWas7Wb2cASHVQNZg59eS1d31mnI/oSRJ25OqlVutwJ4mqkoy1KguaaqQC+ooi91oSVaxBP1HhJZ
5fQib7DZBniTCrjZ5kTcvqQX7GDWmZ5IE8OcAUdjDw/+DewTLZr0nkT+QozsV5IB3drueCr+Q8Cm
FWED0puLyqVbvW3G/qolT/IAmfT1uz6bFO+SaJp+w4KKnm8HTFa9Ip7p7Yac+hfOpn+SaT6NNuFz
Ycg41x1qIkRJr4gzIVLb8+7w4428tpp8pwyDdapa4ldQZj+el+3K2uWr4BwQ9CaOTgYM/6sWMhzG
3ET/6LavyYM3VCf1wcZy/iAnTXuV1wJrekPmyzr3YqoNCs/CywlNwm7HWI/Bba8r2wtEk2776gm4
sJ9L0tOlHT73t2+cR+6RkGVAiaYjphGp3Yt8Kgi/bh3diktKTspWbv2m/ohTpKwXL69827KrPHg4
5QJ5jrvUsgNsNk/m6/B3p2UozbiCV677aix476pXKrCbJN4G/rdKWT1/mK1pi0DxhpZ/H+DQg8O4
tyjSqo4GSTygcrEHlVN4aPi8ojfn7GSzkEIIB3ZZHDFFXyB5c2My0HInCgVfWYYHeqUj8RsNldnd
prm22JTloblgLyHDhObs+t3Mrc/bjzXohLqcPcUawbxFtgxT3FjDAP2KplGZor+ILdZv5PgJ7q6g
81w3PPb/zGj8pdh8cvfO6eGvF/rNiZFw8h5B55PVUG/S24loZm6AkmHJaQYqEeMG1V2MirKCe7e7
ddmW0JSkwbpWhPpD9kwCqwZAnrGrUGdO6DQmoveCaXWsWao6SfDli6OjQrFq5wZSe3PDWGjKKdXp
98pT+OYbhZxZtSzpVz5BCYglJS7sOojJDkj+Te3gpTEUoIq0N4zKveUf54ARi4/FZ+u5Wv1Ah9/S
VvKagY/a7f72OHIqzB+NNxas6HnBh899iwmD4AsvBFv9EZQg6uCUBc1usq6vj0MCq0iBbnOqVGjF
CAkF8FoxHTxs9YSGl+oDcsOhS7xwGjWcGFIjFoZaBZisb0ZhiJakZNcV8BuJZkewaORrT+cUE4g+
xeqMshiWDMV2KxR0GOHWKmO6dDdSADpkULzm7hVC/BF1+pKlZyYsAoP0E7R5WP0aNlyuwsuFcxn+
4insj8REIZHOCP9n9WI+VCeSNrB1zLeDU3P4zqf2vdfn8jrP/djZYmNkrgPxyOsUAGsca69Jn9cd
EwbIMpGjzFv1ZxMM2dIFOVMnz7RkpsbXFNnBMdkD0pdSWqc7CX/YHGc31s5R42MPc87aEkXxt7HT
n5148Gi97o/t98lwKT/I93Dn2TAhYMzAnGvphHuX2o5sdXsq4zpit1Xs2RYl+bguFTL0GTgMheuD
lVEgcLwxtWw6zo0pNzy1Pwbm3p7sNMA8bc7cKYAKEFjc29rB1rPfT6oUm7Z5jmzUNYOzN7kQkFQG
N09PuKQbXEbKers/qd5vbxwD2pyuJVku+HrylS4AyAFTXep0tnCXiJHeZgF2F0r6pPC3hRw4oWUu
9om/70L9eyzYucfo7iqIi7WPmh18H7HxfCmrLPp+42K8xqi2QkOVwAa8v/Cn2PUXYFfMtgx1zXwB
rj46gsclIe8u0CJbvJI9P21knkBEjDTkIfJp6fuWmLYq5Bd7LQrL38o1vSxvmVqN/BdqIUuSF+AO
ATLa33PEjfLVhf4RobFK8dhSCpDUu/x++m4rVqmOluDRyVsfiuO1fNEPe/lTaGzWlTmkBzGZuk9i
y0M5fv71wjll6sfC1LakCtSlwMMdstC6pLY5Vfq7/kfPIuunPzIC1bHHkzVxk5W8EYlA6IynPLVi
tT2P0Kewx4fQnYllWT9gi6Jd7XqjqTjFf4HaE4Z7F8IbrFp5NVl7XYUy4k4dkBgclbRDZrJ5DrV4
s+luo097l7gQi9t8l/nbWQoz88lxmgRx3gQCka9nZj/d6l5QpqmgnK+DpcdwMZRqKESvG/VY49vq
nYRt4Ml2X86nyi5NxSSfQqEeXEelv3mwBONPnmu9AqaFhOjsMxSWxDYV2X7woIVeK0M5gQQoolBU
ltY/WG8+yAErUksyaTwRB47eMQaXYrJ9rvhDoZnU8W/nEsyniL52IQ9yKq/RyZG63X2Ym3En7oIq
GVtCPrDL7Y1XIb2NfrxBKgVm27ZUOpZd/1KgwcvtTywfNgn71XbYbdODbkGZwdWn2C2cx8xzv/xd
KVz2O6RPUzr5xK+xVW3FDHKH9dIE2eUQjc6gnS09i+CLXsZu+EDnpKl0TVX3iVn2HT7rTDZJDa66
LfZAGJ+9fYQJQ5jK2usVClPaoZ/q7uh285PzumzRZPrxcDoBtCzvqpndnvs3Y6YbxAvhRWtx05iU
6TqhtmVAUA3YKaPSsxf1CaSgG6nu8NPD8MLu0FlLZlAbU57UFik+zaWHdYJ39MIb8LfpRED2dgsf
uzQabAnGPte4n9heXcHkdHKHbh6K+M3S1GBzW/E+bmn14E5QL6YmuPfN6iV94HWljNafmZxgiEhZ
jM5WKdN55Qu5yEw/0Amj3N+rN6zf6gVyLo1ESk7a18VtTiMxF9jotGj8I0yAQ2bJE2LldA2xQeyp
h/hq/aPlLnWA5dZCJPqEA+MbbyUmDMonkkFiohQtQHpDCOGjM2EwghcSu/0xQxF94srK107LNd2a
KFvN97OJ0v98rVrp7kdNI6TxmFR0sVq3smI3VB1xXLGP88/XJWdwvr6PI9Iyc1RsXQ7XAfxWydp5
QupDxDLFuQm5Z9pH944gQK8+mLu0w4ADGL9tGIvWtzLJ4uWH9c/xTp9zwOt4v2r0bTQFMSLfcUDV
iU5li0qeCqhncgYj/1TvmcOtQ7zc/EkGI2aulPLKtFm5f40UF1N/2H+LUg8s09hPElEZ1QZ4gP1/
p/7wN9M56x+4fgTylRRkbMTfd+zLpLXuqJHGvQg7mhFK5cAl4+gAQWmrOPh2MRrCJb3/DpLL/jJ1
EKAoHitZ/7wdyA5XA/5QXXmJsF5Y8pSN/HLRxbC05OaWJCimn3QLFGaLDeYcRBfxIHaOIbGe4y9a
+OCsvU7CXzEMu6iqHTZpAiay52DLIlYS2H5goEmKT+yaDHs5igJyUneDrsjZHRlRpkGMjk83gfq7
XtgkGjA38G1/SbjufcDiQxX/0jgMQtoFjs4Qxb8dfA8Pzt+sVst+XhgNWoc8nwdn5S7Kvoqs/cYT
vEr91oFuLct1Dscy4un18E4ZJbP5Hm1lHDQNfsi6vV9pD3FVwggVvjn3VOduhhEllgulPnhK6jsK
SEgh7duBOlIBhW1Bwipv3tHEYYVVQJVbevLtUYe8NtVJI+TDboA5TK28yAznrLH1YdavttmjnQVS
fmS/xE8cZRILT08BEKYVHxZxibdxI5VkW4N7lLLLmmKPT8VGSoNOZ7S9ls9Ljm8XSTHSwYtFF9YC
3du0CRtsK4T5GuhAQUnfk6LwzShpt/7I6pmyU02WtV9IFv3wFvZqoG280UtXCA4RhBdTx+7PuMMQ
sw0YDtGSwYB2Cx4KMRN51BXiIlRz9PS25zfGkb/LIV3CY+H0hLiN4IvJ8yPKmpnVgmjIGdeXP2Rs
xEWdyMsUSAdMdw2cZ5dBXuwx9LK164HBm/lq8AIWDfsT85//XQmckcGL+zmhcfIrmsoxT/AyUsaa
9xw6j20UBxu4RmrLPXOvxS0sm3rkn9X5C8Pnr+j88AQok+ZELI68eLrdgjb0/J8+uloIfTw5IUKB
fzqHsj5+nqeHab+Ke1EF6KzYyTSwRnJqKMVnMNtkKx3rVggnNNhnmyeCGNAnkXMtC5rKj5N6/Dmg
mpB+AOqHWUCi43nRCK5HxKY8HoTI07vMkb4223zwtror56PECfv+2IzU3EJM4lGMcYm+FxnhlvFh
P4rD5nUDMIkM9M1+xaRhjC5laLSUg7kWwNabcUgyX7moUEX7xTBNJ5m/V9udt8eH4GFhl7+/Uw1R
dcOuS+s54Ad+YFO8kayiXalNn1m/hZLK93e18qCsmRjhIhx0kR+V7x4UMhfV/xN5VDl+M3lRuQrw
0jj+5Gn+vR64on3xjlmaamwC+3flMflSUR4vGv19AO0lhKWxdyMnXO+r235hpt3K3u2eFrXDQqm1
WvL8g6HnomvY3Qq3FZTTlAMYijB3yl63JZIngbk6DBwieqtEoClOr5tTIEwG+2/2OjAOgSqOHHxr
15N8smyBV9UGiNPe3EmSxlatFCEROgbKN5U7AVM2EI63hXorgda9frAwd31ueStZumxFQHjtSwdo
nQFA44cGLje07cdB2PrJrxcdcSDU+gHh5Qb2mXmkmnQ0pbx+gTcBNF4kcvjAlVeWKvW2kgNEfSWl
m0fCRNjFXmxFEz4viyC5jhH981HOnSNFC0cxvHVwA9E8zvwIzis5Q8rZkKVaQCZ16DRDcbgLFqIi
qtXXwsCtl//QeDHiSXP1z/x8KQcjVgyxlz0NcbAS7BRDrsg6wZi2cE2EXsKQ427UkSzeT5ssW7bY
YP53q0Nh+0sLly3k6y99YPrNILan6FE/afE28c1gzlJXqS86EOWOj9N4pneO2w+4jkbTsW9AfDrp
8+TW4zryriW+OmIG9WImc3EG87F1Yjvd7ryYQUW5Tg2TTFXHfKdN6H4VJXGoUPlj5eJWcYfZL+vF
hXplVzpdGlpdWc9DkxXvabun4zmO951ygHKcMvZmEoEJtGIZxvFmYyNXINye0wFt64MTq7PBV8S3
1/B7m/LweMV3UA14B8i/GYF51805F5UVuS/iGcpOr/tHpLG2Yn22DjqR6FE7+l88yFu8scnzNXwO
URgRhTiobacoUJrOIAgDQmzWrZIhXG8rd0KPycyA7nFKyJlQqkwhr7C4fxE8IJpsaYcmbr4DDD6o
hB+f51n5w1bE3oV8UR2YDXtaDbdQOwtMCfmpixaPZR+orkph3QteYC/gOcQB1hgWf1vyX2KPcwG3
RbmSOLwWVKrqcb7FRKsIuC8d6lnnmxddeYUkV9cIEiGK368yIRnVvoBgAZKrxFmNEirA/ne8v2DR
Fj5l30MPbXEEuUCdhfVhO4xZU7TzWfTLn87VI68U9Euve22e9BpsIjrj4nt/kDlJeJBLz3T8FhWo
2zlR9107fxk8ppXzcUVYEZ2lWRrQjpewMZr1hxCMnhoYS1hG/QFiFjVMJPKKyGibP5gDUuqsxN0+
6Fi7A+4++vYZvxKx49bM/kUa4VLhh7PvVZsPafOJTITyrjl8E8ElQtQ/ABh1hQTsbkj6SjjfDE5v
TLSR2sqWlx9NYosJeVB83XVNU+rJPDpmZQDInmscCZV0N7rC54UXyO6LxAK2f6J/yib7DAGEhtDX
eIyoH8sldpBHydLhgjr0qARJg4kHskqT6iRwQS6m1LMlJMHxAgvBcsnqF97BqJ0mbQunfdi7rMlw
ija/BiWGL50IfZQKQOaQtd3B7LKnCZ7u1c/A7hY7WWbG4WX8bq7ftTMjWQhGro37Doqotw3BBpoy
CGeOuhDObiVUCZTy5GbWvtZXIuKWQOr+5sUwtpAcXct6tzjIWW/9Xmr4hHXlIy2IjxceeLnx0pwQ
j2A9/C7o6oRUT/m6OHrwsfGGIekSA4ZYVeoAo6Exu9/vCC8oM5w4YaS43PBJo84Gb8Gr4YcqlqmP
7OqoBher1QEcIHFTFcssTu0gax7vpusy6Vm0cemlpvgcdqydJ+dkR0DCzsuXioT97o73e/7RFCXI
9GMWwzzvseTz7FTe6D4AG5kUOb3pQHU5X1FQSNw4bJMbZRXIM6RM2vOtrXPn/t0XFjFsucGYaa3A
jxTRoSzNO0+ZS/QzK/BN95XUucneQLW8bSfhKfZw8IKhxm/SbVIAZq4/WEQR/0cbBKAdA7/5Ldqv
85PwGUqqYmDt5esW3N2K06VcNiBWicsh9Kobjz08fxLo0yhxIiH7aRkd3Th8Z4pTtLGST4USeQTa
IImA+YxbGOQTHlZxh9C2qsT35MIbLxjuMKsOpSt4JFHMvv8yvmu4szxju7QsaXIctbg1Hu5+3fSC
fo9BczrGxgFm4R/mdfd2wCdCXM6nXnHYvLvKXcmbcWfcFSt3LxXcwQ0amZeAEZPiPwZK8wmfWrQX
9GQLrCsAUZCMQoeCY9pR6bV5QQOm1Nk0+W2YyzX3y6n/bONGOmLqWTnHJPqTjekfBtvND4zdwLt/
CvZTGonxGPTUUCMYNZiNsDkBZsbspQMeO1WfqUvAdzSW4TJxxy8UNh5aQoiYlbVr7FLjhD9NxJTQ
j0SnoAwWUJ1xbzc/i5qGm0ETsRl2yKx6pddH5ytKsqW3d1Q8h3kkEOsW/quZTS3AViRtaQ5ZgMul
/F94tg6v+piYKsocXOpvMXDS9Ht9rnkrbT7N0mFt+IDURJwspCUHOI6D8wmHeNNPtDbIKW/yLtM9
5um2YMbfTmiRQhLR+LXmvcd+LHOt+8PQlIJb0ZFotY2q95IpzE/mXhNL0AEclbBHiglkMARmGsrQ
HuXpY2KOarAz5xnxVW4VKgJztC3DsTZ9keofa31S20LrUnhZIVl5ka6xPEHJ5CwYCKzJr211JQh5
U1xzWZxWyX0OccgbTbAMSFNAz6/JEjDg/bwuIFlAk7Snk3FDzUTa2UOa8lEoK1HgCXEewlvHtRWv
3SoBauDOqPqHJj580nj9tMrQ+MzeCf2aoudpifDis/eQFcpAjLaU93wkaXhH0hk4Wer6GHk8ULcp
OoNzDVBNjS/0o9NMaxV/f/4mv/qIW0wVq+GgbTjWN/znIa+aduznxD6UJOCI12ngBVRcyPiP36pZ
Y1t/s/MFyrOJ+bhVIOvf6OiLQWHLqEsqK3X5dbmeYvNSxPslP9xn9xnFxJeCWdR1kW+w6pLYXW30
28p2JqwSySL1vdSv0nQQ1efvYr7jrJkSgeE9Ix8mkAZWUx9I+3nq3dRpGz8t+TwDEBwGLAHqfTIW
eLX0mHvDU8umPvI58ge5y3Dbbp2KbORXl6FDKqbGba9WnssQPChW51Gr3ETVNMwDS64tHSBxaGvL
3UEKzm0dABqJdF4tBozBxLoKp+PjwUWMP6qMbjt8ppa137KGjRTw8fRKcoZ521t1tTJaW+wGNp7u
tXVm/6g/6uP6EAZFmFgo2oGNiD+3O/K0ZKuNQIi8Z0eGCHzkZbp+M7vzO6R+VlGtL/a9LdOFAc7f
o7Y5bFgmiEsHXXmDeD5c1yIlIxrtiqr+CLqP9GfTtMlSx7UcCukXWWGZCRah5sYoQaNc3f/cEEM+
36o6RKDve6u+WyblGpGPN90LDsHGjGv23CT6PF6ztbEJdGsZ+Wetz2UVwWkDrQ26mcEPphCJLm0A
5kdLfY+6Srluj5opG9IqjMo2F22FiGlanOwtIx3T09I8JO9f5GpBbNgi0FRD3u82jty0YqV5yaZ0
J1mv9LT02Rvx09t9U5c5sV5+bbAzKWfNJI/gjaBotByUCsdpEqmMGkdoFBC4+ypmWRjlgExQYitd
DaQ/noA29k8mzAwRXbwnA5M3PQSavk3jEAM5AdElVLCtYyf+0+K6fF6obxyOyeSVTNzxozDIQkDT
TYaV3mVfkAc+WR6e262ztqp/jJCkwxq1ku70eLNa/F3GfeWVzPqgdR5I2jtGCObgJJhf8TaNkfie
vILdYPK65BnzWv+6VPP0g2HQiVFfNrYi0Ia23W4VYpGGJz6lQBn7C/K3MOo0zbf1FsQs/DMCSziw
wHwWqXUZyhdsfPmm8wGA7ZrPgyECNIpXUTCecXemI16IJMUZx8jqRM+bFNadAfPkvCJPKJ/j5DkV
KaacOsaDmaAOtPQ0XGsUyBPhtGtcFfuSrm7pjBt0Vfzu/uzr7fhoncgtSxoxBwxluLtHWDjV7UWb
qGacdxO9ImRR33eCUV64iXfC75souhy3X7odsVlo0NhA1CTK2BkaBzarCzwjju2gv7xtq2GEhRW6
JST3+Gw4UOJTcccIKxQM2rx4BuUKLke4IdpJ0OULGyOrcXesKTzFl1ZHuRyLSBWCe3iWO6msQzPj
nlwqE1n4AbEm8YHpQpF8pIUf5GA7M0TajfQAL06iHoV9LGMwd8ikZ0SZxw6uz2D7JFJiLZPXFHU7
3C+U5yJ3q32R8Ecf9URpFfXLzapNyLG/Il5IKGLmGGnJBbrDsBhGU6FsDlFaIxTZbpmLUty1sHhD
f0njaRDWCBvGx8wNyizVT3c0CBgFI2WJ/egEZySeCj4Ci9C8peVqTjigB2I0xfApZEJQT5VMT4rY
eqI6+FHzaQFlF7jeuSXNwlTmebwZ2AqV4Sng4C3wgamMOC5n0DvMTQ+bmDqQaix+4mtMIW+lVKuT
5/yjbnl/fXRQ1Ih8lrotoXwPtUv2yq2aMXBOWMofIZB0qmS7uQtSRpFcb1PnJaU6+XZEM5eYZEJ0
U1p07bmYiKT831g6WjNsmkTtnebDsRkknv5HdIZLeGdNNfrla7jqyZP5Zt80q79kDotd8j2PoFpG
mGID95KYKbD2kr6EVFZ1hbgz27OYU0UpV7PkTSnZjD2Y/SE5+1WHWZ60UZSy4021N9lfm8+ZtZf9
BTmOFHqgZT/86J8xoLBr+sgrpjMSQe7o0UVHfY+7yuPKsWAE5nZNPMqo76IPwZdqR2imZsEc6mId
GizTt3aYGrX1hICEfeaGfHfEwkICHnTk+1UFQmQtsbjhv8Kcr2C2bwrSOiXOV3r47W+L20RliCg7
CiUoge8ZhON+yri0OA31hBDEzkH9F3qydJsoTTb9ygA+HRKnbdKQyBHFNgyWC3S4AFM1dVDKUFit
ZVTuxX4aHnsSNSMxAPG5SmdKhNoAbeU50GO0IKF8U51c5wlWFMHWnx/iYr0svQf2FUhYteu58c4k
jxgU4ZgwulaOo0ntE7te8Ab34jrmWZcLS/idbfWTefc7p8AuV9qjNkdgqXp/KzUJsEoCDo7fuy9t
JhvH1WS4FSdBo81yAGUU5/4NhfGLqZs9mFfL+6emOO7H6W1rUxqpx+RAQbNOX8cR1KqRY/F6uzu6
SMMkfJSkc4Fj83azlCNT/Qy0WbJa1fCsjd1DMKWn852JDLfwbscMdGuCCDfOwmm5vJ9DQZmgKUCe
cAS8bGl4t3G9dTtl1bJ4mlz9WzX1TOX1ZBO/18Pv/kKxnzN1FtFJnw1Pzk4QTxD+h2QrwZuwd/6w
Sqi+ydJ4rMsWOoGxkveCnpmbEm5TdsbuSx8sXuovuPdn5lGmGKfJqb5IYHfwRFS7+WBcJocP0gqW
Adtxpu3JGyfWCYjmVlbjw2qHIgnG40TzWWk64NswsjDXkmFd3NCJpzzOu8kW3vGmqglsSPNXo1qE
Ahk8Dit0zPduC50UvEodT6DabBdg4E0NFIRSa4W7+aHxw1zovlNQvyxvo3CAfh7aTEZ1G1lMSsGY
Q+2kydrXtEGadQI/669hPvqr0wT+YpLSds/eFNWnvXBepDdG9Xp/Z3s0P93DQQrd7Gf4Sy6mYy3I
urNR6VgNrZcrcejMs5Ois9CV56sIpw8QHO5zOmkaHT/vBexm8awGOi9cS1al6rVJDRgPWzSum3Mi
xBZ9/qGiQhP9AoUajEMXhSbP2BrNWyaI7X9G+f2rh8mXbB0rXe3oVYCHWZx5+FoYDjQJ8iXm8L6V
y7377BX7Q7l0YJt3syuLldUW41JLFdqay13bqxjtQ+JtioLgy+uE+H2EAtXssOsYxP1wqBKDV0PN
I5pnvldH7AHCRttceD2eueEbYduZ/2KbJy2fpXj0WZ0ypDmabL7TgWFEkZpyrKFNYnjzi/LlCH5N
HyFjwOPw95/rVRb6ViHNCNhPKrdKjSMHgP6D2RM5KV7drXSo/eLz8qRzkxLJgk5c7IVHOGNxzVQp
XT53NF/sUg7mf5pKC26Zvxw3KVFphuf5GhRx7cGMa08kH1dE+2SWScmDqS5HFmsCCoRB+8URyWcQ
YxlJSZSdxOFGu1NkuKVcTftn9LGHBkR1a06LdG2VSJBE+wQEeURVcSCCkdbTBHklRsT/RQSCuQxQ
QdiGCljLob4DiACycwu4SL1f9bWltTYg2sx9JWXDa4omPAIjuF4SPa+YDOPVaWAJq/NcWOZibuS2
hMA3yswfaPw/H3GJThzErW4/kJYP3xdFyoXCezC3rr51IO/XG5T8O7oK8TPYN7wlI9+lt4iwOxqG
H6i34aau7B7WjTgtwklKJZ/tv06bctgZsctH/484fR5PqSB9yh7tRxkxN5DTXXSWeglmhmCsG5Od
paZScGX3qKEr9l7WU81amaYeCYv4IX64f06kX4wnZazp1GyMdZOXt3V8+fjewgBOg0MRKr3Ln2Am
hqJ4PJSOkCiaoxQ7eZ6qse4lYcT0ANvvm0R5NiSgsCttDJDa3nP3uuzg15qQeODPI4PGUGVDojst
ylv7+0wwDSn5/FSilYbeFAcF0+fXxCFnSeByxze4F9ErRIyc1hHdQVJoFadYNZk7RyvrHL48Ufu/
Vqu9qxYap6F1SzkpVTjI/c/TRj2GtbEuGWESwcW5INMiD5FIaeBWppyOxIjz5VqlAhO9XY9/OdOW
TxmOgcePNYp9EAQSlFMJM/TRDeZa+GUl5amhC9oGNhAC9v6+gVXzc63B/CxADQ+heP31meYjsJKH
P05nqc6Eb55urq83cdYdSNt7uWnRdcAs9HP/NWROT8bDtR+ujXdBoetiVx2rYsi0mE3EALM7AfBG
xsZRpAtk28ohH1/gEmATapWlXjr5XpdWlMDIdjkrYZsBFtDGBW31KebX3QP9bUfz0nNYc65WCPNX
d/VoPpvjjDiyvh8fuseFJBOlfq3bMbBSGoVdPF3CySBSlCq256dGa9QEH4+misqZp37rK5gl6kJU
FbxAXJHDR2lpKOhK1O0Ge80dw8uWD+GEo21+NYrf6aKgJfCCeWvWTKq09DawdrReiR/2pUVyhH1N
YyLTz/AuNxnCKXFaS8kfDrJ+DCSWTj0+oZzXn3/qHCN/+sLW57xIveZHhmGFnkg3HdG8lazu9R0K
tCIspi0JIAnHurJNF4lpshs5InvzO8cnAnemGeftkzx1+oBqHDJOWMYvKcUTLsQqVimt1yW90W7H
jeOchKjrFHKtl4cI/zxeBcWZgZMXaZ9ftM2emAGvVwa2OVX9M1m80xrIX7BX1Vy3h3Tw8XK0JLlQ
zF1RIPIR6TC3tyX64Ov1wM2rjLrC2kZkvqQ+0eYGPYsmTicGajXD3WILnxU4dvF2cGpchDajN/SA
7Xy5T6SFNGUMq8/i2kdMNCSd0lWHMLhvIdbhspzvPo7V+jEIM2RdaaEBkWecMSwdvXswEDaN8oJ2
Fm+d+peyKoazh3WCwMIhx2Mb0Q7CYPgDdRCLmnA57X24N1CqMq5kY4dgshC9AqhWFZXX4soohEGA
/Em4pyxOUYnXxokJp6X3pZROR0sT6aKUB1HHogmBhs68DTWF0HDxIuH6weci5uAPwAk0ZnbXOJaA
lJwYAEnJMQBlwSlvJUdZJjwnbYhX+lkjZ+O/U4EKUf6U8OJDk+m37T/M/mpRuI9m0s+zR1lDnzth
RSjxkezUIpLmVZDSFxUGPiT7ycx6j18o86Yw1q4Uj+CxAiHUtWTgukJRjVFWm277roEGlof0i1BG
TBuNmCQJz6Vy71LW2K3OVKm27beco9xSuGbgSp6jz9TeS0gs/6HwYL6t8d9JCCg3BRxNZh/cK3DN
rlx26yDTrxV83i6+5U9y+5qXZve/BN+X8K/r6ZipQbNFGlLiQxrcWToT6/nR0x9vQ4mqjbCtMMYG
enaGiK3Fa0VOI59Rjpua4635cG03ynvTHNlTpc0hVyvWJQefascIYLhu+KxwbDh+PvZ9zG2NfPK5
BYP1CwmEMT9OFVwd6HYSxrcokj1k6sPf2xeQNRqBe/Jr5LJf+FtKb9ltuzlcWcJjCbGfDvi7CYGe
MlU8ei5EC72NjTF7FOGZNHs6vSjIAM9NoiRw9E8egg8x1K+jdNumx9ku2+6vj11Eg3pv8KWjW40c
0cKAwX3W4CXmBxtLMmFuClTUGBWpjaIe4i9+cyRXcigVbGPVAy2CO114r5ZwuCrRN7D1aoC7Flg5
/o4YYkUCt8G8Z4Tk6oyD5UXJubOjEFosFLf9XIX4ZwuIN+JirWMTpockJZZYL8FW2Cy1xuR2YMFy
pBrzFytXD9nt4Yd/leVYYFX+Wdz7BPR2YkZngKuHLoPKGWIYqtZCLRaJsoUnXgf0LvU/fg6otldQ
D/YLunrNZf2xEILPwuVgdHLV+YUsdf2Hq4IPUnb2Eg+c8Wp9LfOekTsbmpBFyzzZFjRRzNV9TaHe
qPOOjEdwJ0d0pyKzf3NBJmjSHo0A1H4ntcL11hYLed4auByQuRkktc7OqsNsWtrv5o9N0g+s5Zry
LMX6zbvVZFSheDV7vdovi8U+W/0MdCmtbrl7DrM96EHiFRDP1An3xaisHrZVCRPb1qB/x1fgjn+1
t5xTkucyCpY7Y3mSKLtn25ty5Nv28fCfequqQdyooi0dnxBBPNE0LTO59v1XG95FU0P/WQ2JPaVs
Ixf73Xy/K5JaL6+N0rM4JQJO7IgpyVdVysF5v5J7PJp2/iuWiJfT3bIjJwDSR/Mbs/fUJwiSCjBQ
tWe4k1CNrOrx8n6cUMgHqc6nBOfbGIhJpDWJyndFvzTf0QeTdB07UeeLbFqQIPUG/h+zRizApR9O
Aj1/4X2UDgUjtUxhQEHoOTA736jTufvGWjOJl9/E7nM1Q8o+TVv55MEb29BPV8XJJNJ8FFLrXbiL
RDrzaonK++qF+oFFZ3jm1oqGpEY0K6YqfIaZ5oVYNqDVvQ0dJFkAAXlu4JUvBHbh+kJVHkYbjRHs
SHurO3wL4yaX+yNOrht/OVJzOxWi0nOC52AFaI0tcAcBwizc58D+HUs5kvbz9a82LzJtRC2NsCpL
sxgpUifmB4LQP8BU984K7taeVdmQH1pokV+LEekuaZIvl+t5LVtBVQG8qpWgxN3KTHHO8UFLMqBr
4SW6lxBPieSdt7itDi8hgwq7sWRiUDthEECZLzowN9s0a6OWc0yRfUV7JFX8FCxYXAspxihWC+9r
hZLtax5xCsBARhw/928D6pFizozOLE67JMb7O1Cu0U1Vg/JuUvYHlgp6PkOlDcUM3jb58t+Wr2Wq
+toH+JFTcgBt3SSL/0dOn514Lx2hxEL8Sj0Xd+jB0ixnHhkQn5X0P1RhHV+Nkgc6K/PD9l198tip
9FXuWfj65jDOq+a8byhLkolxS2IBDcNlAe1S+GOGlji0slVf5LBqJEYotQY9Asva0stvOkcoJJcu
PS4IGTjwy57X+QlMfkXuOfqdSW3WWoca4sih6v/gtZb5zz/2o3DqTGm6IUcJd/EJDlx22khkpGa+
zn3dmO3yTgCZGlrjjvdtWzNpicdgwEx3x/yAgEDNUjXKlfxgmgavEHZ3EVkTQfeRvjDH9fI/EiFS
SeeXwgXXZJ7kozR6YW5a0jcfcLOVKiVE1/HrTV28ND6dKhPTrxqFctGUGMTcpAq5e32FrOtVRRaj
The9U3DMwZQ9qwPCwkAT4WBCojxget2OPxscIvywRV/hWAm+6QUKV7/1VOeZ7vDM2vlloFv25zEK
6+HEWGQ/ubAGkdcgmf0Kqjk04k2qLPipv3RkXl9TB8RKPj8weYBnveT3FSQ/1c0zx46MD0Vqb6Xl
qHhrYmA5EPhcIBEYl5HuPhCrcvaBs52sDKOT3c8EcqdsCrrCyz/oxafNm9Hby5Dz4SstvyCgITHP
ztAjjUEapcdcQ9OFJWWCuLDQKzt6NYBWf7kCOWfjoFlcqLgH+YHE8VI87n47ztG5WoGsF9r1lKUa
o8J1rKVsXBQ+0RYPXN+yVvXBNHyYbODXtdfaxj3iTh2dMW4GVNX1GjEZ48YjYvGy62sOxTP6NE5i
l3M/5DXAOr5uzqGZDEtJxlkAR8WfC6ZN/3mZMYwhV6B9cYMnQZGPcXaciYrOa8eJcdR+Z3Pm/NGG
Msv7qWuxZAA/78UdO9xvLeVmWa2VO7ELZ+Nh3iR8rBf6jtyzlDgr0lhPphpebuqH/uN9cQDViXBn
LCDD3XNORuprFnMUvMYyfDH0u75ycMHwy7Qic//zLDBZNalDLQgejsPGD0lRmcYwFCcoYeKgujGm
nMsTerw+2KoN3/Hcu6RB+RNoQ3Xt4J01TCMvDudzkSC2EGcDsXibXlgegcMxknYQS2+d6KSI+pKS
ACRfxs5+1WjOKnqVtxx2SBK+DGLVBtG4dc7qZWzrq/RG3wzz/ntqTq4FTqfQ4taFazIE/j4MT5td
OCMa6ofq+/2L02VlG6CuAYGwngoI7QBmnTZgSpCZfDHy+H6RzFeTHg3X9B0nTEyXEV2PjdHQ9gB7
HLMuJmV0zdE+r3W9ALz/6xUwrOJQz0RlaehWrGx/Xd2gUPR3Z6X30eVlnyatH4stpEusCqGXU+hj
qYJpiweBbC8yZvZvRVcP66R5O25VdjGgWJPpBSuL+NeIs8d81x0a4Rdr5x7DKDNsBS/3NBI49run
lNEq/no3Aa65JDUEceQUtgf/efIEg8zNlhEsnqWSk7wWHz9OZQaLsBKYiQscYJ+0AQUdVlxI9Ezi
Bp52nz9szWispU9KqIHQmXehB2Jrm+ntaTdO8d32pfgDMbp7NJO9UYQA6WBSH5XEwueDFukmR/7p
ShvEnZnKL7hTyc7NjFsWK4dUD6xA7Q3CCvoG78QZRNaKKBh6+QFGjBqVeH79ocg7FPwDOOBfFANA
A/G89Px1Ic/4b7Wk8OfHQvOVXvk1A3ync4Kciqk9F0nBwXRYexv1vIg1zzHlukb+UVH74rbVXoXE
IpdgU8Y6yiZSbLGwzjWNEQLK0RkPsKOG5yPP7+fR4B0Admf8+PxS7WRiifaSKHqQ1W+GgWT0Bhng
vaAuizMwaus/bqlfE5O6XnMWEABoUafazx5/fDXyZCWG7TuLpVr3jviJLwuDD+waxp8r4hT581KE
lDU9xmYiLH01d4MfVbd09WNsGILN0tmjw1CMNeUMAwEzeSEI12z/TvSjAsbQKYbDZ32SpIG9Vc7y
Rd9VM/AUcxczgR+8op8OoL9nUmNFbHyx6xA7E6erRtDqn6g7Uo03U36TP+l33+N/60r0fbU4DhSI
Xy6bqdNS1UdQufdZ9WbcmqWjJTnsb+teQYt6Ovbr9FwwMmGuT5Jx7BoimhlHZqQCChgN4TlsrYEt
qcl/ktVGp5eyCwdTmysUgaaVbZyX7C0RYLGUfGY7/bSnwK41JpwuwSqZ/pBhkFtW1WHu8hfXzENM
soDSqDYpbwB1aHKK38wspWaU+7XzNatrscW+M1Ye9R6kJtM6k9E327c/VwRafmTMPb029jbM2Fzr
0MIY/Y7mSSDczbNMpxZf/RVA7yqXYcm04WFnR87dtmwxCt7r0Pqxzja2fi+JEA1e2eoIz1Cj+yqc
LRxXenaHR/YvVYP08Wgg5iLnnDxkYrGHjc3NrGRa+sAlMCFX9e9VY1JyBVaIbEhT3Muf4VaztmZT
yDSxZn+TAdZu/ei2w+Rl1NjNC5Ag7hLtSRzIT3K0/bUbaR90ouapAUAJcKenDegXUJP5N3g2ik/K
qQvdFnQbDLlmKgkPW5h1h9N5FwquXBZRUjRnt/NZRnlt93w+9yhk8XlLWgjgZHJVndSbuGSdY6LP
X30tutiO0Nu9I0xIeWEcfjCEL6OaGMPxGnYVDqvkUafIeV+4GO20DMpztaf4oyqfmDYW9eX7Hx+k
iOdBneBuN5gvQShZBYG9mHJBXNDQDUtnjPG+F7IdvG9aOut6XFF8hs+mXGx2JWR7nUtZdgHJnKLT
H5l26wqKIgC/Bo72GxjxdOyviCtwFkvcPTdYrPFCNP58qy8w8B80ZlePKUbgHjaBgobuNT1X1YPg
vDipP0fyUeCMYlpNjNBS4Uyt76OzWwgmN4FowKC1ny+pf5Q3SaGHmQ3d0fcplO9SAnNsFc4c4/wD
3cvP3gM16jhy9WEzE9kOLBbS3T5k8/kiRcqBdNT+p4dkxOE0BJPvudTLhVfc5buP1uD3JfVixLwj
pGylGK9x8iHcQ7xKeM1DujC7tZTKa8Akpp5cJ9re7aW1B1aAh8DarXuah6Ei7UOY8IRV0vZ6BDv2
2NaucbHfqtp2ri9kcqYyEZOGIO0PS1GKptfMWZZ5bmT28nl4bl2pWscD8KxqFOJwNUTTfqihEfT7
y1ga1U/Nshud3DwONK8GGRDmnrGhcsX/adJ99FqFpIo0jtCVFkzesDlU+l4s+uySFE9p/qyNaj2q
Gd2MklETysiskyYT7aTx014mdj+cHU7UBvsqKUdObOEEmmAeXI/TZ8f7RTEMlZifSQORRCXhDK5C
tnwhifXfHRxkUuXhdkvThtt6pgV4UDAPOODNBHgH6nh1J5iLblP3GSB6SeKUJ/3JQdhh21iJSYSP
AicLaGHZeKpSmyAdFY/evQIsbqgJFHjbrM4OEdTNF/OG09OihMcdnYSJRPmREItcXV5pJKT1bLyY
qmF0IFM3oMLsQfeFB8rO3QnKMC+xv9NEvh7NkfNqUKbOX6r8mqjFAuuEOwWg3Lo8PMsOMYwAuBRJ
eRCUSH/nBV1ZoGKMGf5hHIXfp1sdx3A7wHbKcZPoRs7Ri+MK9PRZL4moImh0rBjswns1I5jxPukn
f8fzZADG6oXZ3t8IACEFW/j4GmeEwkO3BdILKdDZBszQmO96AA8bi2JP6uSwyvWCZOOS7LwPXS9t
GWblzDEuhE1v5S9skPOdDM9RbWfK9KZl4tVfPa41OIG8rkTLk75XyL1JiKpqVZlSfwoqM6zcKDdQ
P+Ow6o9q7lzfpjnOiXNxSrLjcZJFnjlQyNH6NKA9SiiYg2n4p2rZgkDT8EFZXxAjBcxhl/PbzT8Q
bLOzlKz7x1qXemFHwA1EYyWYpB0scmXhDtib0iRIavVJJue1uiBZs0h7ST8HB0r/IjQipKlKr5ZN
sBanTLx5Fztcp3Hd8MBOrpRyCO1JskQJkIIb37RWERNzm1/sI8YpY+xBGB3VfmB2y61izjX0y9bf
B/Za1cyCvWgr8p6lLLzmerme6Q97IxhypxYtFhnKn/LLQwmZbPjxIM8jXb5kufD/3lHRDQsD3uVR
xla/kDrfaAjIGb+ofzWXzaDDj7tRbpFcA6Fztr0x/hehPE+XraV5asPW1fQAYrG+B0+WnXikTQvr
1c/xh30Lh8iQeyQgrFfyq1w1i/UQfjvvQo67kXhn0dMBUjBIOqFWMqkRX6Z5fyuEq010EEqHgKiF
ceVLrHzWPIG84RfS6DYE6uXQ3DkE6N7UBc4WMJYYX71OWXfEf/kCAcGOnXYX1CWT3SYuLPLHViSu
kUKmFxWE4TlBkhGJqNhmRSe6yWVUAgbziscndi8k80zjW5B7OobFaB6yWjThBXMc3bhBBy4KNh9H
jdKu2gIPLiV9buTrIW0EoF1yEgo2ijdYrKIbfHUG8+MJsg5LYZ/0D1d237boR83vCakz/ncjaZ4t
N54nrHYZuPyD8ywCEdYjCkktEYLOdMSgPzfP5oB5q2tphF4AgvbWyU7xU4m7+sMzOFiqbYt5ovts
LHbrvxyGl8sfJfy3VuMANf6bdtEFUajriuMqgVuMY9MViDslSHMYMPvpCC6XHy5/e+ON4eRcOlQE
P3PEeSXGifmmcol7ufwUNlVlE3NfqkI7RGixB86ZH9diVpjJuWAAaNioarbquBOCKzD6J3yBkQfM
pUIVGi+DlxYcKj817NL8EDU3WQG6zFudNG8hlhPLxcsSVgX3zrCQwIP9/TycRuhlTI0B1BcJc4kI
hya/iIPc+xoN4MnX548D8yYsUV8n3PRHMkQGVNAn0VMIY+y2yKE3KNAKn09Grkw3Ph15prPbH4FB
bIl0z1OWAe22dvLwHAVtphRNpnTKyy1+MVmXmHm2nSR/yRH2gUmdXofm+AVcHXA5kjGFV0bKkQ3P
7N4uSxMLZV/5wcwq3xasAzfqFBJSk5unAJZmO40vTSjB5OgNnKFBqMvggvYhc3KVx6mhU2c0k4Xe
QK+jsC5qg15DTNXl3xfo8/sd1/FDFRalNPaMj5LXV4LCRkTQapbZiJKLC/Bw0nHI9uozCLEQRRoK
P/uT8HoCKytNe81kRPUKI6gixpcckK//Tt+GF87/RAXpkHrHhaCiuBQV9b0nzOJCksWievUh9VvQ
p6QLThrdr+/lPHnFdbun+zo/6PJ0bdBDgy7++UWl7pRp1WRsZe4/uTjnaSskVN2pN2wOG6r7Iqhx
r8fHer1LTHGnb5VDI7LqRpuMOTN4Uwg5q77vcr5mzglxBHIgyg1Ui8r9ZVj7gzvTpDnqTdwb8y60
GCg9E+fGgVaOHrtuswjh9JpaTgHzRSg90WiF7JIhCZd58O11vNvRPuyVqGfBVio6DAV3L1He05Ui
UkOT6qreac/n1unro4RXM6vo0Fe1TC8Gkl80VkB7zFZnZrCyYvX7XYWLpG70MJF8frw8QMs0l3/h
15KPySU2dbTeFq4+IkYAzcf1jl/HBfQ5A1LLL2AHn1tGuU/9N1RF1oF6Y+ujh6fivCWxy37sV1FJ
R9iQ3MLFvXzKPwoVdjsIh1rZk2qSqGYpmiIr6yflid1FATMK5lcuk5mnXbjwiaXtzpPasPPWbyXW
ETUUxC/c1ssnv242LbB1G5OxEDOV055ba3zHPAAk2mVpsK8M+MFs2rtIakgDcH5aeSZ89xvk1SfB
E4XfbGD5dkqb9+6o2xWKiVDmZUO7dc2KbfxcFz2No6SUMUIR0WUCLf3QZIdmkG9WSq/Em4tG2z3w
sn/rxzf/49KAkGBbsjgpNFB9PjhJSJYkpIrQ2iAT9JlUDaTz64uq9m0KtmiccrKvUOCUgopJ5Bid
xAWUDZujDAZgK/GyKraCAD0UxEqlyZmRECW305hCyjF+RRLlVYhEiDxu4UvhoyGhvonTGCyUO/VS
grLD4MtNYUUBsAe2XbdvHTsDA8vbbYwoJ28pqSvvubBLsjpE+Y/0KmCbtpwq2oEjeNyn86+6lFfG
kku+UxuQPWhIatzpLLtBDZZYUkhDyDGNUOJ11c00p8Xmupu2fFOVDwrroexr9aqZLc8mYFl/xnxu
u6399u8gHDnprzKmRDYIQmpTHWeXLdhIKGbqxzh50LWlZgulEc2F6WylsHqLj2Zt0wfif3oMrAVh
1qAzFK1IQ7POeXdvBeBaCkEp64Bl/vADCLtyzsOqSANJJiioWR5PaJI1fMl0hqO7KOT5H3YsyLux
hidFBnNMnTy9ZsL3s7R2Hm81jVrkT3SeiHztqOZz1TISAjoeop7TDip1akttRs+0XcB9tMDuFAys
06vJaYkmrdXs4JUpwE41+TBKamdFeMEcSHXdG2fTG077TIeb0hrGyfw24FcpOjzzsqLGn+7Vvj4s
fPBmofYgKESouYibXPYiFOFSJW01Ke4pml3otefVt/1iMWRtP6zbC8c6wx0bBclrjO3m4mzCv17s
cI8fCuq09crBnfJygK//wo131lJYyC5KJyrBtFnZupRQD7pyUVWkmT6n46gehB0+siYglgY6kT3w
rv0tSJK6hTDoQxWOszYTejXZKLC9akTBTmCQ12vfuoP1s/Ofveud9nhWVmBmb8Lr3iRPtnQEJzX+
MH7TwmdVS6PwoJY+aumBP6GXHkO53psHefEvDcXf0wgqegZUoqItVLl++4MfCOiVTmfdFjhV0Odp
yqTzdLZO7JbHvUBrGcBiqy697VlpQTz/RP17Oz6nAKa8nN6gNzZlzdHVn0WnWVALjsZMO/pGwLM+
Ab89IPeKPvoLEGpqo7xfSCCzdax42gYMxc+cEikG3/wyVhAQB+9LOJ+8ZEaJPc1pLV98aNxYxSJC
10mFg11F4bDL929lCd8FccGEKy3+Um4n2DuaxEq0XnwLpejOCN4XBDxp3mNxNvX5KXa2DIQ5XAJC
q5tcgMBb9Ju7OK9oUcroNek+Rde81RFbpmm4pMd5Zu3vn/SmR9Obzft3r4mqbhKmExIzjIATrn3J
xJxiDVGosC4MOLsIuuYKNRv5xyK0evkrTNWQ4yzQvVNI8465q8CCrhRTn8cEkiCMl4bsIVT34+db
JxG0akihxgBEOe5ySv+1xx/SXqdE9ceHqj4RLO5KANY6dI1MQ+VLYnLYTzjCvlHfQKPuAy91xttk
7INiFLf0uVAzXvewUz4QUW8WE8inQ9ITV9Pvl03/DFJMs4P6hZSVYtyPil3lX4taZ0pWKIlAn1Wp
oc0ZnLycBi+Mu/0laQJWT3rrM7bQMYIf81MmgJ14bjV7EmYeNA4pAPbkhMi2UHhiFfw4E1+Xqpqm
Xhi/haK8Rbf0pW4htj4gbSB94G2pU4HhCVl0w08eZIklvTtFUWjQUSbhuisoMEWuD4UDQ6xEGG+8
K5nhxMteC79ySSoSbF7mwLrkeH5X1bj7NyS1ohT7HEhL89jheSF0+ILS9bUgAlEX4369aDOrEpMY
hiEBPdVj7dg4igc96oo3oczoKSS8wU+y/p5x3DcnOsxr1+yxBRNhh3BJ4wBT1VE1t3QsTw4tCqsD
877ytymDa/9lGfC3yaR2Ysp8WKyw7+NTVG8dNjAFxNqAIQ84zis2IujpXwp6jntkydTxEUfbJr+9
08V9GgMRPuwQc9DlrPdM8OcNygGKePGZ5jYMUXWQ7drc6n8f1txJwXm9moQVsL312t5y1X0D34PI
kcsusS9l5sMkRTbCpW9OuPydM6Q0QhiCfUGhHuyljYI7QtB0T+yQ1l6oXMtyfNP/rRIvblh3/xCU
X2N+E980LEHl4ehnZVrU3qCBDbnfvz8pckaq9+bQtcv57tdi2GoWp/jI8TOYCABan4mfF7F3dvEu
sWEmiwJ4jnd2ae6v1ntTxNVhYXznNONbMfzxKv9r5zO4KYYjOSNei8g+NeaZRTRrCERYorw2HKGw
xiGAIpxs209U61YAlJycvxBh6trf52j3W7RDCld44gN6+j8firqCTdINNqTArh5u+6XavEWnt1I1
cOMwmr7Hi61AqeucNlCLz08FXWWKGL8EuNTgAnm6bN+Dq4tWIZy5+R8CIP/L9MFxxbmb3NcTbJnL
5bKvdkoGMXa9Hvq+f3OZyZOK7GSAGMXvJ4pBehMC2wvEA67tdwvLxDrQ9aMRcawPdUvK2FKDDe/+
0hHw6iMmkzaxMmelHrRagc8JnuvMiz8htv2UlthwzPzHfAfSB8UkPTXjJ4MjEP1HsVGzTOlvOfBg
aXZ2uG3vTjpnz6YvWT/pGnpelBOZocsrb7fnFWioNP1AWi3FqGpr199nJnygXXOhMg9LKtMs6vud
quzxta2r3VzsUIneU1VJs3/szzt5vNXnn3sfO02EV1YbBGrp2gkY5WmjSwkozsLmRZlgwIlT9uAd
/Yhgr2ih3JBgV5o28kdMTMkT6Br7DqGBAUp1ukDJQJlRogydLACcxpE3BPCdZ4AFyjSKZpVIDair
qsY0ynI/74Bij2U5ih2MSrwZDKT8wmAgWu+bR+59iqn9TsjPa2kmr4P+MrQEHLpJ4cyl1N3s0C75
e4KFa/e8tmIpW/xvtC4I9FObXHs63C83sh5L/ct7e5dlaulMASliLwjYTjDAEMdc+7GXHqAJJBBG
6IhPE/k3hV5+2Hx7WgqnIePHfNbxR619OTGxyGmOa/OkIx2Zy70PANDJojtQGgdJk8fcf5vlYKZO
S7mPAnmBMmUdEv0Vz3TC2inr8LN56Rpe30kxC9FkKsQgdpuy4B0Sf+q0HEBYCTMcVn1yyiQUO0/I
4Kt+iK+aVT+nnCmbMJY7mTaL0yF13H+iwNytsLI4yOCRr277xz22J3H3pyXuO0G3iTL9twIWG6bq
AQcOjnYJ6KNq1Qx9YivqyZxTA9VIbDM9KcHLy78QPOyDOrprQJDSTkqPt+0nkaj4bYzD21f0SFAz
Xf9eJF+Tgll/jAqrZm2TGi+Nf+jYCq1q5ZHx8lq7AKXj5wVcXYEYNcv5hbiYxvw0ZrndJDTAwxPL
ClF3/g5nBg3gPVNCY3FMeDzqK9O86j7cYA/MYeSikbnM/fxEu3KZOw/Gqj/6ptU/KrCe85vR26as
i8UBwd6nudnR1QPnho1cGO1WZCtHMjbRLRwXaorp21WaJYUec8xTIT9f1GXfGEbtE4FCrvVjEZV8
RFlA0ZvAdShy2UBPGJx6Ay2UnFnrRfs/q4Xv/ZF7hv854wfPvU2AhH/XouHZj3JgkxCPyASs0mEQ
yl53NeAWd7j2zZr2DeyOXAEsW4VQyivn400aYV1gxK0QZDdSM3tFEV++m0ePFXzyfLnvVFyRD13G
alnuG0E0X7ZHtuv5dbA4jxxiQhAhBwSOeM4xiykRCmYxw4WdBC78J9kzd+Yt4BvIym+9I7hmXTRr
+Ei+GiDcw8gddQBAnebBUvS3wsgKfuztO/x3q6Rc+gPLvf6cSF1vayr/vp6cenGv3AF4tDmWg0EW
JGTtTJ4te0QGAC2U6PI3tiRA64LaS1Y7qtiX2MufA042EE/bRL+3iIv97CPCXgFtqCKoqs/ymmvQ
ic6dLxwE1fEKQQp+A2f1oU3YzWI/WFGALpeIw5AxgIOM9t7sRvcvnXIDjxfiC3eyo3cJta97ChzO
TtLOEDyUHMnYeSuulCraf8A7Pxq/DfliSST16VlL5voEkvEuhta+Zc6xxCnWNtcGL/zmjiTCYHbS
knH6lrZwx4FzQfOz8bcv2QTn+9L8A78pcfkiAdAmChcDqhx+DUjtYsPST0dE95dF9F1/Df2RP030
tHiQvFA+JrCxTGMP8QDsvlzJmhFQrLo5iET2fyyqXYGyj0w9YSIRP+V1qaJNkfg9F0SdvQECvw9v
BqAS00AJKbv72uSlxR0IJjv3p6kyzqwGrFhaB3NOHBzA6f9EnNrVOn8L12XyBbo6DK8/ynn0PXgc
kQsga82CyafU0tiCLoOaouC9ZxncRrzzLxRi1mk/9pUjOM2Vm+fnA4z1Pv+4S+mzBD8e8DHgF4RN
XdkADUIZYlb3fy7+J2vf5DpcfgwU7p8VZWaG1a7CkzvTbcG9hFcs/ygBCNJKk4PekUNBcr0TimwA
olTNW5ROb6bOklf1d+eqPJi/NIp/5r2/zVSWZ5PpU4cI5EjlZ2QAYSyh6saZZSe0MtL3jiO2ALBd
Ozj6atqPsGjj4tVpa4m227rQhZZFLRdquy0D/l44JTqt2mmp46P2MpkDn3B9hGQ2VJRyxiUTvNPe
3f3Q5qqlhDHJhYMHSB+eyR0SbH8aTbgz66MXO90wuWuTeZ83ChhP8RPvySfyiqmKT6HaG/4pN5t9
jiiWgvzAbnghOlw4PLEdzO1AYtZ0JIAkGKWpLLGOq70jC7mtpqEdI9MakyVf982YbST3dNsHWkfd
vQNWyhCSKgfquJoprZUsVKxnQwrvo+ZUDFRohmhkRD+npG/QOmSs1iZMHo84Xffc+HLk6fC0yohE
/1wKNaXXqq/UQ9RYsWy974tHRDTzsLCtN49GgcBtFXfVm0ag0ynK4GMv3pAWz4xZlw/8OtpUk0ag
vIsYA6vcBPIU5453TukaOGJucr9BVoMFWVFC5e43L2gigPOyo2F54wW3xsB+UB6z0VQgFML7q+Z9
ZCSg8VAk2ltzp39wlsrbxMpCkeSpkMzikzFwbc16T/GWN6KFZvYVl22MyYj8KywVhwggD2VB5out
hCwHItrnGi6pzlyfzbNvcwur/Z8SQozrBqyWlRa8CWyiw4R0eYqaLrT6X30Z2lFd6V2WQYJ4QD6v
0Xmpi4U7NkR04n5eHzkGxKFp/N6DeJhnkmzcpL7ypEMP5sZV6FWse6PmSg2EYrkBJitgpOnEXbtD
n1INcA3DyXib2QdnCj9/iDIMfGYeuSHAm1eX+BLOrAeqUpbart/VEDX3TSjyFqx4GdyXjZwlPiw1
2OKxktQJjWiIyancnlrCDK69d8bhyGf6/SKmEEdhS2D8eQ0tC8P8yCCTXrRZXKZdHizHISbfDWzb
iIJAgJn7T0DX60SwcqD3NaPW1ikrpK5g17IVdYSDKpRWb34b5zrtJ3/Z5dX2A2Wswy+gnh9TCWnM
3gh41XRUrpXxwX9LmTB4ibJ/aSPcvZ6K0S71t2rqxUrNo1Ipnlc5bHaYqwlh3QuI6TdetFlyaE8c
2FMx+UfiiLkNdxcrbJZX6ZW5UhAE5C7yseDhkdB7P+6k51GB9aLEziFp/L7iGZjyELFsddYpm4/c
T8M+YpZdQHkWZariQbXMRv2cVcZoK4Y5PxmosJW28px0/LnbLb7/X8D4po1aI9ihyPzo13TqWT93
kRnsL4ljWZkGs8hL7ukEDI4CWNiN1MWm2xaX1dY7KIbl84gxZ3KkHxcjH+8SEvWEnvQXPhRc830r
PxPZCjvKHYmFFePMpVN3R7cvArxfB2wH2NLchmod6V4OgJRovZyoaPnoqtFbzhbgBDIWcqvkPFID
Ci5p/BmfhaM55XLdcXgrWtAteQoB/ZtDQo8iNnZdRQdmOlwchs/jM39bDoYeJtTJZzHeM8ikBYd4
TzJaboecuhf/e8t3/B/8KqrmMHifQWvaFIP+VHKweoTg/n79qlzV1KpjR+6/u3XOLWDyXXH4kuxu
UW+xwLW47T3C7ecGPFAo7oHrWPvYcGv56UzIMnDHE4K+9K729Ze0MegG107QHJY1neGBpOIPUCgO
ZRwacUpjxar1ncW+vljJKHogaWdpz6jpxKAI2vdd+13peuniSSVpD97rGlZ6195yUA4tmZH7zhQQ
KivLE5XLh32ZUzxE/U9NPs89j8bcsAmm4NqlVZ/nkGGioAjFuntU0Lt3vEVPpye9K/msGxpFlBK8
/wOCgScohtxBWqxhNdfNh8BcwkpR2HllgpBB/xqui6P5H5/f9lgbQWA1xUmGF4Ya07WC1QFvlmux
VINfYiqC7VyYbp9Kt4KhP86srmUlrwgmwsBKAoT3QR0kmgypcKO834LzVD0JbJ3elqmUMXFjksqO
Xx8qaFDHdGRpHXYjwXYANquErIlAgcd2ug5JwFcfYeZWyprzTcxc7jw7FkSqnEWIN8hRs4DkhQ5j
ca5qx7rQke4xGkdfvS8nZ5vUr2flQElXNqESlIfHOaztVbY302srmUAA6QDLiRQRlCzcqoH9l6H6
qPF4LbeFqXWmIONnBuocoR+znZJu0e9RoA6Pa7RkmIDxx3rlno9FptyGlwuhcpc3tygqeZyoKa/c
RO6Btq558eEPi5GeOBr3cVo+GgkvKslg8jhyzPM7iBCbP4e7nh8USsy3AKHSth3eq4wYjARVFhPs
JWdUTvh4jnywT9KIpPGGApCHNklqvpgcg9mnmdvmquvjTYb1WfKBt8aEQT9mIOeJwRbjqPQ3esje
mzUTlXmjRAK2ulnebX2ZAVON5x3/6k/LmO+Dh6Jq//m7ZguA9Jbd8rlQCW6CYrR2/uaCpDzFDltX
+ECIZMFE9/IHWyopiJgv0q8BCIAl5JfvoNzzXcAVedGcyEWlRxQ03aauoDKo7JtJC5+PM+9fUI9q
AKIPkys6WS/ifMWFjHE0y/rX5ycXlmLSLTBWaz4WqLwI9Zt53FTElJILxLdoQFYI/EHCfOjxOKeC
gQrW0nZKPGDfNOnfDPHVbPRzzNcyeCih1vwJC1wEYFPqPxgGMzgf7LAoIPcovmSVNwewie8qzgZR
QgUTvoIiChjRO1VRZMrsG4DtDIsen/4cCVyuYcMnTUsURmYT+TXtj3uONNmKxBGkefcX+hAymRTY
An/LqeTmxxc7ARtt1lfJSICKVRCOmDdW7Hjx38W0M+VJ3AvbvzrvtsJJy3Mh2j2HTrGvFq6523vm
vQiZ6BCxHJJ84YuQZnk0Hvh4yf6tbY1361fGGVu8DnW629MmGOoHrAhtGc8RvTc5G3Uf3Bi1ltSB
B6ZmsTJ/Zj7k+/vkUyXu6SqfhBY932gtkBz/UiYdLSbZC5ROU+ec7cOr7HuDS2FbzAKSlHNO0v8u
3fN9CXdjGqH4o9fdGZ3lekN0Qr9bx5ZR0PXVRfS0L+m9SUD8rP6CUxFRWVE/oguPyKilwvRk2QN1
TVASZiFM7ge5s8USzg7a/71Hx1dTCQ8gMVO3ivE7fvn3fFIeB3TalXAFPGyr4HfS5+bAapRI3EJ2
zPPkm5MGj4dDsmbAwys7F4J7i2ZN5jT9PhMq92F5Gfp/1hmIg857+bsFdC3KhXWHBNVLxNCMKhRW
vGXy9uoLhTCYHQKXGYy9hrTENZ4Th1xSlDa2T3K27AWu4VO8bo6AWc+yL03kTbqVl+udlz6fZviC
ld1hAILew9mf6zR1ovD0zj1unG+l7+F97XApfItJ/qQL5s/BFfWxlsg8G6cErGakuPA2F5fk4Oc5
3Eu1dkBoHrmB2nLZb7NrrNMPp9trYF9YTRmMluBMYtwX2B5WR8SMWdceDScYTb/R/MbnalB1m4zc
yZxiIKAHchnPn1ZcmJVK18srUq3UzEVGaUGhMBCnyp+SHkCWJf7OQhwXgNvtn8VH8wtxJ7K4AJpE
K1PC2D+W6n+CKrN2ATpBS9HU6vdezob/Y3Bid5K2L3sf5hbO8SPEEVw5kUJIPFHKD5u2aM1rhRXt
gBvYEj7avtXMqVc7uYwlRELh4Y6a3P+fXL4q8STY6sjrstR3NGbeeB/W5a+LF8rLS/9xRj1kki/+
uHlPsM1wpgvdbnyWS90a7U8zap+bgJ6PJxL2jmawLvQcpAfyKZMZix3TmajeSdyznsFJAR2o8/yT
Tud8zXDadvJX4K2SD6SrRoYv9hQ79up07UTshdS/hQnx+7wZXyEnixDC9Ld7i7ZRaZIxVXbbkrdG
Q8U01zyIMB54d+R+aIl5/Hji/Z7eHeI9UQYnenhjL5lTQP3uRc1wF/lGMkYTME7igFEnHJxsQD5n
oocpMSCEFEwxNjFtCojo0ujT0yoHEWGTZfm/ZXaWCHVuSV9OxqwTTpZyg8CNPXIt7ElIY8Ik39Yy
ZcD8K2VR/zy+Te8yTHuibL9EcD6uRZZFTseKRYGL5vNVw5JsV2bjwUw2Pq5tbNDxoNae57HIn5GX
fZd+tuTVg1egZ+G5w2JhJAy7ww8OWpuDXuYSfPuDz5ZGTqgQ4DYcfMprS2dqqdFeVXodvrCp3AYR
8uSD4wBZxvzJsxMKaxSuu9qPMV1crd7ZayOIcjA+cFWRQHS0G1R6pMYqP+wfRY35HMjC6C90GceK
PNsD4FZ/KtRNktDGQhdW4CkpHj5TkGYCD39rjhIGBivr7+x5G6bbClskwbdu0FeGK70A+0pnDKbY
gzY3dDmESXsl8yVVkzcFMv6f3gTObnl2ihFGuGxHLcks1SiD6IysqQXpIcJXSskCbmadkjmnYt4M
GrywaQsz07j2MRn+c2pyCnYNsdppGDgXAMXkVFU3Esl4fH1Y31L70BgPM2t3i/zjQFCdQGSt+XQE
J7vIyhg9xfyHYBMQHGv33LodZSgxmhOkrUcuFanFDtTF1Dkp7jE2++sXNUIyfhjVNDnRPvl3On1Q
MYEXnmSxGj0n/UbdvhZWna2ncpU6dmnEZzF1bxt5nGzeRDxvab/ceWQ8/Vw4NOlkNzvVykEPgEdu
7KNrPg8Rw1t0hHXQnlbiRVWuciCx2YA7HbrrlzbPDWyciKHl5mnAoBzG6jJL6gDDmqGxVJJjqtn6
57BHs445mLp8rE1FOG8xyvrtMLT25fTR4jVnsYdvY7rv7wh5Ff+2GqGTuuiMjO0ZkJQeUvGWhW3m
aSPx+N0J3VuVOccN/MvlyNWzbQ/8rYJOVpdKjdMcJHoJVIHgrfR1p3Kd+qSAyef7lVTnR3kyHQRV
GEjgFtFwrh5/286YL/U7K1lCwIht1YRgNeRFYVwudagBoehLJLKUtrehr9WzCKrApiTH7cPFx9MD
6u5MDgofIk+6UgseF2kM2AOF9uciiu7iLalzXRviac2JKcfPcdMRXb7Wf9wpxGqEIvRR58wROLX4
ohlDptwtPVtoxJILVNFBSzxdZDZ086FAlvJWDP3AoHLbDJZw7+apssJ9gnMi8sruTHhVWH6HcD2p
8uaPDY3RwMpsu/AFerjBRZPpejC1j4k6XuJyoK/NH8xLhovrS3H4jgWtwU45MfrAldKHQ6lHCS+8
i/VvYJInVJNmpTfmKcpRtEGDdhyCbCWqNxshZzWlNZKpLNlFx3cB9EjJqBLguToT36V+HWZzihzq
pnUgEUfbVOFbczPo80EQ8VEzlrKr4eDd1JxmQx6L/kQs9Jpn+rsKW/VTACaC072VbVWakUcAjSAq
2dSPKsZyQnBDiL6LYlvJ2+OI5wed9aHH+DhcZo1xcYEfTVv5iiwzTRHamC6qFmgvsAxf+TE9Rtbu
HxFzhVHFkksJdQ8pSA/La+8QRed7g7HwSKcZsnSfFxbZlxGonnHcB6Ar8vYh5WstIrZKjB4Im6eV
q4H47BP1PJzS1nJolELhMEFWEJMpkuqpf1nQM7p7uenymvbez9PeBpCUpRPKvyo8LNKKlRsplsAw
fFLzJub1xYQJU06ovD75fvzEb12oIUfyF8KCWrRZcwsh8DB7yFoVDWH1k9oGKWEy8Wax8SDLSQcy
VaiPlTWhm1uno0yba9CAwv3H5MMAPNLb+OE49ZgD+s/cpvmVlvx/Xyqi9PYh+TBCIjvhvD0Nlbbb
uFE7n0gXLdVjaTTLRfgqxz8/MfqgvDpiHgr1ezfDQKzc2dixh+woaL29MzQpFQNF7nxhM0+YQtzB
0VlEsgBqonnunNHoB+6Yl7QCEtQ3By3HPPSQie718gwNsgmWFsBn1QB8N545D7Kk3jmDpCRF2S5v
Ofb7r6F6qEM5MMgAX+hMlBIHjHpCebKxLSoj2zAOW3I26MwGvmtR7JOmZnIfI0Nb872YDxp0JqDT
sI7ZXNBdzInGivTnTEsuloF9hvWYNJf0Q+XYdTwYP/FU+c/mgjrcnZpO5IXdgADpQ0I/gOnfMW8H
mpv/iVhNdoZzbXwRN8oJIs1I+4etL2CGASvvRbDeP2cLv3r6pVbMB6Fed7qjkmEsJug2T46mYUn+
djCNnJCMS7GM2pjFbDWNPh+TE+WV11Lfs7SeDqb8/CmmM/dlobNPhsoRq37Igge9GpYUurtYMj1G
A+P2KDSxOQftBHnDhwYtsu86bV66vnYon/kVVBCVroby1MiW1ZEXFkDXeiXjtk0Ed9CZmKQkb2y1
G/G5F7fPw6QOaX16J5HtBWTF1CKl3+HH+54NO/qRrux9+6lrAvkRcJUyoD1rGQ0jrHLbgKRHUAkc
fBTQiw1tCjHutc3tuX4DXA8MLj72pwJbokQiRSgPD0crFRwjGiRMgBTAV9gzAsI/mlBdBE41rAD+
EcclmgJDIcLn0WHikWYAWl6/GbPgvWGwOEUaVjhN6HWyNO71AnNdGs0Gzo6mHY2aVSiGgNLKPg3z
/uaXzvPDF9E/57Nr8gPMspVaAjILf+tNnwe7uQlJJIM0UAw4zyN7twsb4lpARrZ3AQFC3jtlVqA2
sRHZv6K4Dubozg89AscJfqIFVL3+Ajy8YmvUlj4rW6n3cyN1Itq2mbX51MaVn7cYyqK2f9e7MbLj
diZCR1OEIvFyBzXj1zywd8qP9pOL41N+JSnaNub3A4DDQHRvIVGYRW0Kmrj0v2JF3roq0rSyiOly
h6hjk6miBvqUkYx+2iGsdpfwh83EnXXgIuPJEg7ItLYIs6cqGc43cXFwUMxQFqXtu+J9EG8sO8QJ
BXYSzIUmah0hk/fuIoVVQi2XWg4xq++AHZ95FQEq34sXgsQ3HcT+CYKw/mvSIPr6uN8lEg+QJbsT
Iv+YBZDUY0EgEgJwlt4TKQs9AELKmLh5mXIs6PL66lYRC8/vL228KsOLzoRnTgi/fC+rrrokwCLa
Dpu/cWGRzBty3LmezcvXNzprLoYbCLQcRyxDSbWTJ5Qm50YGw1jG3oFQ3ACVgjKeKttjpJv0slfk
qO9t9NE5vSmVBOc/LfJ9+F3HFWVxd5JXyoSJ9N2J3JR4YCF0OXAw7u28QyDJUgxMX+BDPXJudNWq
tJKv+63yB2JH3+zPRN260ElNSETY/WnXO/VtJa0Q8UnzIBr2WID1N5ev9Dr8WbDZSBWl5Dp3KIgs
rI+vOv4t3VTtxuEGrwcvuy1Z5puPqzyORhq6hCnEYFybToa7BN/07yKaMJ28P8UT84aktBr9Sq8O
n5F6uZRtNUAssR7NjtwOF/7basxkUH/ofBGoBB7Gh6ThAqzvR/77MEAAx2gTMvfqCtmtVNafFy/S
ec8yEgQ6vu+NpWcMVfMPm3SP39w6NCL/VSPBaRubBnpNSXLEDBJ3L1FJfvFyFu/A46IMa9jieR+r
R5Ltzh5u4NjX2PSX/cbepRJqcqKuqPtcz5I0v8v3cVDuKCeuN6tve/83jBPDoljG2nhzuMDQh9b5
bPrP0dmZ8fSCIkEUcHKYkdnO+Mt0WrDJgXfinC+LSabkrNvpEMcRs/880hjn8ZQ0QYa0CFyCGUTg
toZ09Cnsj7eIELGX6laedMKYrnwPs5BmRzEoFMbrOvfiFuXH8lXuQOiHcjpUGdLfBOIvmaG9g0h7
XaqVJrpcnBR5ViQgTSyvhUQkZAAGhREZFxtAypIgZJQChjxe8CQexrNkayFLZ7MOi+7M/Hk0+vcg
yRMQhvLoZcraoodqrwOLfToTkDTPdKjq2QTQ4BqqZyJsr56XvwY45OXH23sHSvodweHroQ/RazEN
D0/my3WTT/246rsAuZB6rI+1PFbawwHEoMdCoEJof0dNOPj5EDzQog33y276YjChSJemzcaP2tlt
h+TMqw7vMiakAlSlN1pHv7cV9usllZzPLnT01Qw4T9l2CHiCDFJgjQQxyTDika6EiU/6s3U/FfaM
47CeUh4MgYd2o6yzKJBsJKPWuQ1VbzmEEZfxw+UHJaoQaxhqW+kS+UINvEne7k4R7e/mWAYALkvv
NyXZzq9pTyXUZ7XrChdDsyVAQZNHoNEC1t0Je+miDEnCwy58IVHz4jCLTd/aACMVDFWVHIMacvYk
FYrBABQZe/OGQYWP308fUEvxhNowVZNudF4xKlwL4NFkluqXeKgd9t2bHjGmD8A+g2juAqXF4wyd
K1muEFb4c7OmaUoIGHwFQ/VfskMUcS9X1yn4zGc9y6cCHkkEalC8SApCqE6jXFh2if5kabhsKZe4
s+OKRACsvyPLCqMDcJPlNRBMicRIMfBc/gwykI0TNBNvtzZLdpsG0UEx7wyLofuFlRThndxtQ7Fh
l8jnzXUexK6tLuMMyjytUOrgnvWR/v5AslQCP+9hjCB1IeHwQhcO2bJdRihzZdNQK3nZ/5E6YjTC
O5Xkhlg5mWOKHH2BjdynLruBdewR8hEUDFnnu7BuLNZAy6JHdqKxdySa6gCIDG439ZuCKmqesadp
nhcJxU8yhZ32GX+HiqLKbWa8K8IjmN7EhpbjZJjVL+C+hBbWPeq5+q08/z6IsXMqbEfVXKD9pb8X
zdAsNyKQeW0g3/LZdFXTHdXQ4eLXqJPeDUeCXCtMhG3aLF03KUH8L9B7yMQs/KWgpWcFZ4fpz/TQ
jMLmQ2aw9BW3DttDXWWKwRiVj/bKnZMIs/syVBhHHfnku5t25z0cNU9xjDmz0RcSzQkZXOUniX2p
Fh543h76PXG7N9mpV1+xejQVaq4vEB1jGBgpKo3vzkXiPjNvTkYD8MezNljqVbJJTeWV3LUYSxlt
nE/IVTtgTVZNTVgx4UolcddkdjAkCoEtF0I/XBSc2dcohIIZojETTKd6swYV/SRRHy8Jhha9LLOi
KLV2PopYXEUie0VVLUGYSDu1+H6xA8oM5xz6BA9SsAdh+8VdjP+Z6tVIFBtlGuX+wuX+9NkU95bz
Ub26ooxq0SNHohqDow5ynGIqx2+6jlz/32Mn4R1hty9bfH+6YoJQm42JoA34q6T7JEL6dY4XihRe
UbAcededCygZ6OAZKdThlDFs9vStJDeePiFcmuoOuiqDGRufiV8BNtD9XPRpG2qJkooC+PBU5fnZ
zEm1ykjfPmsVch34BBeROzXE0TbcohBynpuLME5Wt7x05qhBx+yYRGY2khHNGzGwSM2RRCGXxChi
pCFibSuvD3Zvr7if51ryYGTHXJedcAnEe/wTOpHNR6RBhz/t8n31laGCei37hOYerILDUnJ8WwfE
+/Bby5/sBsSe8qw+pkM7p6C/2QOn6XaNsOfIMpLmmg69wYbqWH/su3mfVBd6wtoDshXD8T/RvGCv
ZSP2CHRPMFjOphemafcriaTgy14LGxGNsWjUVKVrpm4r6NEGjw9cRwwmMfzOinhg3d3QH1MieoIw
8jZDdhG5GTC7dKKr46F0xPrA4c/KwqI7GZX0eKMh/zxuQ+5MC10vRMk4+Jow7tyRu75AjW0OxOab
8OzyyjCK2iIfLC7WLBCo3AZc2iiduXGbvTLQnwQ+rK4WNhcjw05oqVcBI8lP3gwPNqvbF4wahJeh
d5po3o9ZwEGTzXVdYWT6DJYvmarla4+utq0fCiouHh4cIDB/2ugVyUcjeegqWUg1lBYLLMs7SJ3i
52cDwE9dh9cP3nKfgKqmaew6klBUqADE6Tz2JPUzsWDxy+B1SI1Sx3b68cloWn3bFaJFRa5WNVoh
cYzwtnQIo+ed5zsZ9Ze3dSfMtZommFxP1NCZ6xZFrFv9+FfzAY7K+KKVE/6aGCRvu+zgXBDOAIUp
cgkSBd0s8cZQj9v+0lhEpAdLEKr57EHZGpcfzhCAcXLoT+rNxcpTSzavB6umw1arfP9JoaQQ0h2m
bVEhUjvidIa/cVwPC3AbjFJpRlvszelX+wwrWTgibhFbg+GMf9MrHNy2DhfWvgKAYZHjV+sO93f+
up6fKq/mZS0Hqh+YZrpI60RZheX63ee7jAF/B0NkjcD9vBttiMxygCz4sqyRX7mJI4FVvNjffKal
x2h6DwOUkG8ZA5EdwUKycozT+U82F2hLEEgjzeYgCgJlQ3UhKIGgodeM4oA0XCWCVRGq8yVMnuBP
qm9I7NIbz/XXgJF7tX60PmigVviNMG11Ykx+SFRFdEuDYcoouDZvuOXNHyjo4/JXkwma2d4j0UFC
2NA3cZ3I1nLYl4qRVBKhsuBQSnYWRCLwJTFlzlc7J2I3Q+49fHs/6n25VSkm4AXSzYv8i5jwyBvc
17+viclmFcIE/vEhefF9Ivd5S5IMGDLy4p5NzK0WK8I9fQtcqg4qcRUU0upCKg/bBrOAVozrOs6p
EjJqxujkJ9WRtndVyzugm49hXMgEhMhaRSnF5w+lOStmKUY0fnKLuwA4ImDcrie3jXpETKBMJ+aP
BdkCGrg4N9Pj3MacoYpzNB77pb4SfED9S8SOyIrMApAprHdVwFx8Ovbt1hkUOzjWjIlXp0xGYLrd
ymRjJWDwfG1BNJMM6XOidijW2hbCxMyknts9e7AMJdgTv5IStjCR8oZuCn+PAXtJcu3kupYU3NRi
pFEZBozz0Yveab19pyAA0KL9kNWsn3j45lJi8cvbxqEm7ZqeSiK0b63n2AcuOYN6wTAdTN8/wOJ9
8qRJui2UsmXwf9tjr4tLbymeYd+LoLMEiOdNj9qx7Dv2NxrLjmE9a21+mkVm7Q8jPP56+EV04jub
AWS1e4CqcEy41UhlC1Q8mcYWNXcjrR66/833HeKUOXpvvskkIWR9ujJ9g/RaIj/JOYnKbTiwuH0q
lFLVGs8zUFxxkg5vTElMMR7mcLgKNqYxHwtHfNI3huhX1UGrhQDvKqr/HDIgkkasXJNwbheQNSrX
j5HZYaM07tPoUOGyB0QdU2dv0KtfQ685/pOI+KfwYlm+l9yqSKXHStSlv22hKB7yO8nQmpeSHUFn
c9imzH0IllnnHh1f+Hr61VUwpeMO64vXizdPkYIdKPH23kC+REMl2NnHMyO1jYzoMY3Y3ZFZU6Wx
/XoYoy+n2nyVJQgQQM6W08a1kxMndf6Bz93Sq+GcOJZZSqNopCoLfp09ZaCOoaOjNjcqilo44htR
VulBlXwFQjbIWEa+1owKL8ASL3VMlN4ipyK2IJGLLn2IOVHKnqiXmgYB58U0/3b/MC+oLM4auu7y
OSlDceOdB39DTHD0VveMZkhIib1D9gwmyL6SiI21fbmgKu7wSvGVx3zMPvps5dtLuBj2g0tTJfBW
PQWYqyWLh489eif6kYZa4wQN3FlfEtlmoK+ddb/H9RdcGUyvCyCIeBEpmeQRbBCF9dhPQY4iDrBu
+nOeegQYqCbhJ5cgOZO8L+PtUPd/9BZSIZ+mOfZXqoTuHkZr+Qth8uGft+7AetAwQe+3cElnDPQl
ZXAb2rmxH2h9kaSzf0yMmkVavn8nFMb2OQy5AGbko8IJr2QPcmUbd9FOvtVfqHbEqGT2HHaYAuaS
nN4EDDCb47Qx1gRK2WdmSRd/8DPznW8ohVeOpreUoa7g+cY2J0v46zFFwiommtMfQ4MoIYUdeq+s
1yeaM6hKbPfXYidI1wbgTyBEodL1AxxTtbxm0aKwasmPZDiumYgas6GX8RmUFixbdLV6tGiRACL2
3P8b7yqh4rufw7/KHeoHptQv96Rt36o7ivjlAtd4aoryhPpIzfEdqQvqqp9ul2/QuirxCrU1ATsN
KrhiGlUzmwHCyGjyufa/My1hAvove2TfeRNZSBmqYOrlx2VqdfknxkJl+EJsY9+7L7GI9Olo1Nvc
c/qHgLnIUZ4NCEkcuEGo0YwCvsoGnl6YI0YLGLT9xFsDjBK5pix4WQs/djkHgRv1LNDXn1FGrf+y
TxJ3tKmsY2gLBA+wyL4/PFKn0Wd/CZIC1PUCB9+sQE/cAsxeCDiGWb5uWFjZ0V+Sq8BilU41cGBK
0mG08ON6acprHcbDOdpYYz3Oid1qu+pXnFoW9Xbs0k06SbjKRKYFMFRDBsGqeaa4T0DaJd34ql4h
dvOS4vuyo3nfL5JeU4PIGeViT2P7suK7kcrQ3ev8opFSdfH5byRWNaD+1Mr607HSlb1DZXrFW+hp
dgaQCNOd68dAc49NEDJdmCIw1fpOMDASwYcMVbIINM7gUl1XaIAIyQTGUF8IiFqmtSuG2NPyWyVN
/xmMlm+r/jdNa2GwXS4ouDFJIcHEmZC7hk7lb7Np08QHV5nA40tdwNUvvJnL9W5faTs6v19hCxtT
hd1EpNn2l/UIcRfpJqpJHw27K0DouTBFXSL7FwjZxHzaLPQ9mo6Hm02Z/9zsqgzwflrKsgnFlJga
PfQ0WzJp843nWSYSCjQ4rxOyi8pzuBpNd8p8sQFo8tBvc+dRzc4J8++MIhjJBPVVl0BjuHJx4Zbw
U6jPicCcc48cwN22YzF4kfOTx5u3LirCW3ngyuQEs9f7sjaFSJ2i5Z/fzb/QNIwMVefKBJE9lQ8D
RkfULxHAq2zxTeEPkNyj7y/cWZv7IFq0mvJsJqRL4eU1rJYyCIvbeJqend8fUJNHD4UOXgt9nJ3z
Yx8R2R1Rb/BJKTVStM9LMXqLmEMfu28toHjYMjMmOhQsNuQKSm8vS69jQiPFr57ATKKd9cbBFiVv
K41ywQyLJlAQkXftYFyOuBSV+DvZvwPmLcbCyq87pIweURptXzC9CUauhgB2e3FCm67VC1M7xZIH
sHG29oMQv2rWRQkf7/IHjVfCFbidxDAjGmXbjB85Mhk9jnOQGy58Kn/WbpswuP13pHIsplV5oYIE
Er5L3gIfrXgF2SyI+FTFwsWWF2V0fLkTfIdpMjqh4ox5Pe55zvHTluwAtvV2LqOzVPHkSwq4YmYn
dErYsryE37E1d4EZer1621HFKAjRz+WTPNSvX8zckgUkjJetvOsQSZ3zkRA/dIamWBAf91w1hIvT
mrCIiL1tZc1KWcbh2XE1odC6kkGK/jZkLGcHeE2fFJZbNa5g4nfRyJYTGd0EDRQeSLEwQECbxDrT
9/9qzoWaFZOlAwQhqalpO8SwP/RuyEkGjG//xWfGeTqlqFT5ng3WegACpWUx1hCoc136OitIiZHt
cL16n0Bwy3KN+X7gkq4oW3yOBI5pD/mDUd06Op+FZk1jibvU8OTWJW09HLjjPPKSGSek/xgcGDYn
agD6PozyEEeasqRqNM/vcX46TdHwCa8m1fcfZMiwx/k1bq6T2P2RJ92ToM/yD52Piso1U0b4Lt1z
iJa5McHbo7kjIin+XGHOhMWLGee1Rd89Jux5RmrnEPWi32p/cmOKxHGgQo14QMD3zB25kQXRKuB+
atGwMGAZw/X+8fyU+uXIpfz0XO7xEzqKcyzlxYf7u6mf+n7POTRJvPtA1a1MyMGJoMqgCqirGUqp
sXu+sgYWODFHuty+kXPh7CQPCycn8ORTL+uBeq/sPE2sLTHqI+qxQuYjEY5eEg7BhpsRVogPJ5Wl
KYlAzE0qq0YdtJg+T/RfsHr/nTN0reSLEznVQ4abdhqgiSvcbjPJ78icLfXbxcgTGu27Eb3hQmJQ
kFsuiuHsCFLAHQ7qXPiBBkAvxI4PeBW99mUOCwnmu7atGPXJvOftQitYHM6OOI+Jn9RilA0MuCsw
vKJX3Osf8pmm/v/b5aT8jxw08eMUbYsFs+F46jSECedzbcmjjiB+g93dEXUAlqmjyoPtCVPihMRi
TfknxUl7gblri1EFJuANrLFAY26L7X+W0vqnkwN5EHO731jou69bXLVTjG70Jl7G0D2zw+79Jlow
xb4xzSfufhHuRAKt2pvBXohBK0NoZf30B1dzK+loFQBzLfyK/FA5E1B2SAOfbU8fOCADb/Wx97dW
Orn/q3Rx4hdxXGB4XgNiFEhoDMfon7Xwa7kUqs57uesCgvybPgOYiudaamkT5xAo2Kv6aBftxCvn
kXpOyEnMbdANyqt6S+LiPOK+Fm6yrDi8ixpgR8kQou2m5COy+4pioCCo+dtBU6XQfF3WEKsLTkyQ
uCegtAY3W0tWOcKwmFkYyE3FRWVrXVlYR+s53+5Rbf+MWTM9a67fOTn5XyqcOPmzNxsEFqFVTXWG
7P3AQ+0ETtPl1F0VxttWc6rlzavn5mvV34sGfmbquPAQ8cR1LlTUpedbp9vyY4wB7bGbG4P0Fxau
/W2JjK7T+EIdwX7ZvWMFscoCrCmrSG625G+jAoG+3XEpW1HHONdmb2XK2gjEHH3LmO/2DkOgCv4F
ExsJ3EWPb9GqMXPb9uhprE0WO8Mc97mNiKA2YnUimq8H28FfXlc6JocM3BWfzaFLlSMYa0jmTYrL
GXq20Rjrfisq27bcjjOjdFHvEfmSuWG9k0IrEbdF54ykpkgBmhFPSL4OEH6bOL1M4y8TAQKHBXXo
o0RjXEBCb8LfrPIjXCYd86223khEvv+NNLT3SYnneGiIYOhwyzINnkSpMtTkI6h3DMpW1zC+uzzH
1r56Duql+1/8MebcCcebTJ4crfQyXfXVXAtgxNBavW6G/x4fPXwmVhKS38lcMCBzCfnT9V8bm2Ya
FV7Mk9eXmNKy/qQVlLEDVTtaxfGYhtESK5lyQfj6H+64uU+T6U/P++VJf6em72aVXzEgHmF1Bcij
+i5z/RXFYWjfZJXUOIQHNO95LAzFt/L+EJwq30tv/eyUNB1D1cwYnHetR12xNVkGbqB+c0MxjVz0
hKvvG/XO+JArV8RdTM9GGO5M1por0uHX8gmYclpcn2Ui64LKAGzy/6HN2eD+7E1C6KaEWxeq/WrR
aKc6CR0hbmYwb5tg6XxqkYIDSc/Tn4QbsPvt1WVspBt6UEQwEkLuOVsjIqDX1NpBj/4J833WAp/t
rYVjURp+1J5A5NlYalI0VgYJOqGG6u3JOUdeEr2bekyECR7HetBXCCSACNl/9CgeFzyyLvAOwZDd
3Py4IvAX1ZCvC6KKwjnzU34GJgzVZfB6gqKzGLnJrUs/UZAnBr2w3Zjb9sbfx6oUpvOBvz0MOeEV
JPQqstFMkvW8EWeTBugLKPga716VywB1NeqOPpwIu0s4ChZWfWvIA90O2HbLEyqYOobkyG58RHfa
5pXmBriryANpXJ4De5R/JJqqgB4mBf1vk4/GrlDUJbgl2ub8itu6jalAHcyl9z8I/gfbW4HSUsZ0
4k38ZVtKudfUhQK0qMnuQSv84H87qjTHltrh6Y8+Le3oCFMnYPDzaCo7YASIptbM0bhDlfeBm57b
qQvz7lNrg7x0nft7eMRuuxMv0CKHPxgmgN6XNjTn4gbdEYWS3zN4HTdXAh/76NMPK63dYR7es+Ps
pWt4SRmMw+BlLMhw9BRWKnpCLgLaHJYdmB4o867knrywsD+t79pBJEGQBmFK332UF96/ekh64Liq
64vHV8Cnf3ZC8ik7PrwQM+TifzeXTdJDnWunh/qinhWA6dMbWFUmsC1VrCgAH7Np6hBO8zCVTUAH
qK5c3HC5au3Fv3vUla6N7eWF+0cshrGiJnSKsUdfybGEBsXNavxJh5Zi+61BrUFIAFTkYzeXra3n
7H6VIGybQNFWLq4hG0WsImfIGm7cQW9MtI9xePFNhhWiV3Zas3+04MpZ1A19ArUr42jJhuhbaouU
k0kf/qC9M13I68JKjlkCb4iRCQqz9jivsaxYUn5F+kKxnvTs7TryRtJTUpVOh1p6jQAIPV0y8Qps
z6KiI9nB0Q3jOmvEL172b7RP/izFgv3Vgh/6VguS2Evi9h0rVTaTR5wEZENf2cbcFaau64uQVqiL
AAV0MF+VbUNp2/r1z82+eX9tBab4A7OtajUjthxXzsrt9/cbdVDU4h3mGNBg4AjZkRnv/InmAhqB
ZsYkqcF6dIMZfS1gsxAMwYcoW+seRnerEodiI+HdGyZ0UZV0DfEn/fmwrayv9oBgIsp59i/47MhK
1cvWDjF5yPg39klUw4JvYF1lYc4m2/ghVLmoQi5WKSv8WqPqKnSDKbnUApCn/YT47+s9bkzfsHBh
Q1hqi4V3A1QAt+sCkjf38fkydoQHHlCS58PST+7LsSGjsVL2J15Hyd2SDp31kUVDwwVRLgvSZrrd
ftK6r+l4kJigMMs9lh+dyPPtQ6alccQ4GQuD4vcqx8bxH+TXHjbKMEE9jHadOdYrW6PGCyW0UR43
bkVNODPdOpZVGpBb4FWe3qN7ZWJ+phfJRv2QkCfjdwwNQFng2h1Sem3KB3LbPUg+TqkI6rh1A7jZ
DbghEB24yZl8ZdAe9s083QsJab0vcGcMzWcYtVQHo71TvMoGGTgs72KWihq7tq9z+PawhIDGR18t
Kb64aY0fybKE+l3i+G+5Iek9W1NGpeAao8BarZeEsEcI67UsVT0uSV09lsQvvlY3T5/FfBMF4rL8
1QKcq2DkYY4qUftDDtTfu/IZZEBdPJw9Mi5kHIpEyrNULS8mHp2BM4uydmngaD74XMyf2fG2EOc0
G+jio1OxzEJhpS58OUQq53JjWt2BilskjOYk0VYCrGun87CC8QchfSPbUTj7XEZzVDbRZu1zo/wk
YkRBFRQ1XfBAbqzvvp6cH3SUcJQhEjACBfomM+MHmj7b0R+zyZwocYLEvDzMIAoLX5MGcsp8E6hl
RjLdKPejou8RiTWckksjduTrPSr1Ggiu7OwkFFaD/FNx/16a82tlcYY3Vv5MoNJRVhzNSo+9uliq
tGz8um0rB+MIdJjOC7ZUijqebRKAvpOgazJk2ElHg9s0s1DxJ9/gKWXJH8wWwF24SiP3aBysmo0Z
eydw8v39LKKh6qF6ktxzAojlRQnkGWmCXST/mPGIbyIvEtfxtyhlFnWKOmarVEjRrWlx3UL/qGWO
XNG9ZqjQTb+wOQdRh+v52+3tkETM4Ruzpt/h7Qg0pxsW29SVydwUH3qiqv08h0cAR0pG9rL11WY+
DzUi5np6xSA/PpStO9dPaow3AwoLlkMESlHkyelB7zm8J2bfZyTLd6Vfb+MYNlaImDnqmX5O2nYW
f0ZqqSGP/7JyXfjKR/uyIZweMs8CATMBG6cI8LK9sPcxYGTjPGGU9izBQ30RJP9r0jMG19uFd1eW
aQjoseK7nWo0Uh0Hw2ekv3uYdhUye9KDwdWUKuClTV9bICWF4uBC0PanQVUkpVjzjTtxw/fvgN/S
AKX1cItV4gy0hJ95gasqNjxP/I1V2RGlMXlL+sSA7HqOJbqQU7jh4svZs9VDifiX7qTYmzydikFx
Lf9jty9xHPVrdSCnENf79RI3i+WARoMPSfunIHjCnh0m2NPBMR3ripHHLkztWZe/W/U3/mt8zyQc
/fNxrqN3PgYAkX7S2ApmY9j43ygQ5yIv0AwUrylk2um8XGo6yGnIoK0feAc9HbKu4e4rBGh0Vo0z
Z8M8BU/RVSqP117SC7xT6QW62RdLbim49KfsFYMkEey0b+Q21+EHaBGQq2Win1uHnGPZMC0IPUhp
I3Zdx0Ip0fZQd0Udp/N/79bbjab/NgaDtY0TaG2Dus64+xg8cFiFR4oy/S6oXG0PCV5gXqdBUGbX
fIk7dJoRI9FiaJDdsTJMZdQ9TQm4kGCt2TVEz4aJpCy0bpRTUF5RPm4pEpY3GJ0HJWiSR+lfY4rj
pJz26cWB6Ms/w++0u870UtyQPQCmUErYpRjJdQBES6w5Jy9RnePDkjWXuBGWfQPwO/5OCVG9+4KW
butNt8Gax3EExnGbXASG8v07zz5GLmIGVmZ7xFOtlxDO7H8flIZzztpZHVFaSZPhzug91p/1pDyw
Ens/9EVzbilKo3l9T5klczWYitHsrAKOnFJvYtx0gckFcq7AyRRfIs+oxCl7aaWhbgfTPRzTSDCn
78aOtSuJDhCsrWNSraIquk7yf6yovoSuOVbknwvl8M+caiqw1pc5B5WAK+NC2lokRlc3fUjoJ+W9
Mquhld2WfDlefhzRmDA+xAlM+FEDPYCefK4AadJNhwUIJi+mPStmhZf+ToVSKvCnt3z6M87RjiNS
arZy411knmk84qLPv7+QCsuLbxHcS0ytfnJs5KwXdcjYvtKeC1XDvjQTDokKx69qO6IpbKxrsCO2
Ml+GpE4+Ri8IYURXjg8OsC+MvH0okx89Oz9RJ1VBkQHDleT1w6j62srWzhhoKqccXHwz8KEd1A1+
KQcyoAKcKd86cMm2WT2HbOTwH+0ajXaxIgfAIWHEOAr1lHm4N3bOYfyMeKV0X6ZgsmLX/wbVulHm
yjyv7KqREEtRUqSMU5d+Ceh1B3XELrp0+z9s2+p+cb9ZFwE3WjPgvHfUQR/NR8UIyhqEVSj7VKZ6
3aEKJt4SjK0UMvII66tVKO9hZqETHFih0L8nZNCi2+6I23hypCGnLbrexKbo9kA1lJy9R4vUfr7V
yki3Z3lNOlA3iqUQ00Z0EhXJ7La3De/UA9xX4dh5Ft/h3WTBxaN4umafGSmZBriutF+reaMY93L1
oLCywlNi+Gb1G6eo74pZgFiPvmdwu3BQGkg0YdCuV/hkrJbv420+d5rz72WFkgCTwdQTqZCVysnl
1MxqYVnKfsVekRGkEOEWY//fKqyQ4GXRR6+cZ0rg6kufSZOfVFbuCJslV1Ixl7q8o+1FK2zSQ0Dc
sOl7Y2OjMZUOmkffH35r2PTVgBCzL/j2Xip/uyOGDVdAnL1rZfNwumUpR7s03rZOe4RKh27Rj6VY
e6eXSl6yy1N9T2r3pH7w1gRiR4FPK8qMuuR5b+RaDLigLD09JKzV/I1JDtCtSPfz9ugbqggvx/Vp
eBxWj3aYfUkSIPUZ9RsSvCkrO16DGd+qvdYzSGOc3sPWqtp9MC0YvSykIkjAzKnH/K8gQe3XKB2v
GWV68fvTu3C1MDbbRHMg7oZedUpjhALHW4n14ZrJK7HKn/mFh9cF89u3rwXrNFPS+bws6mr12TxV
azuUTwk4Wo/ah6oG8i5Wk0p7FiEjycyinlrO84zOHnFR2oMIH7b/1aMVWBk7R5Hji7hBl+HSN1f3
rK35cRJRIQr0H8/FkzxyAiv4iLcFISz4fGbh2zWfs2hXq8RGnSTmZ3gbDr9VN7ULAVUOyGElryOQ
ZoF2HJEYPX0d/Xs/RzzsWz0U5YFSVg0nhJSbhmD3AdoUsUMYd/4w7ab2UOcsWtI2ybcYa3vTnNA/
6a1/oTVl1eYYSvoJo+WAriyo5gSrDeh/IbrVjz+pZp9N9Dqb3SUj4dJmfm9lE3wToUXAHSt2pFbU
3MHZbcuO4fk4u4OLd5TXXpKOe4Oh7XYwu+8ivRIpx0xnM4amjCsT1o2oLnsici6OFS78ELqrfWcz
KN2uVzSyPZ2xvYUjZqa3JoDK2tXz5xtN1DNk1h2tYYf9Zjp1DuINAyM+G3ReQYKZUuobfa2GA9oi
cJNwx6utwD2bTZpSeGCE6yfqQNwSmWS0IAGSdnZikd955d+7CJLs976tTQ4ujAeaqy36QBaUljxA
hMe2Ypzu1oCWost4cSKedxa/xvxnywXWEe0W4GmlN7Y30/bkvO9gFZf+CmiWgHakERQ/XZWsQ/aQ
7rmrei1SQXjmg0RdFLCKRwz4LRGQKVFOpTCViNxh72S8YIBvDFxm0i5UL/2hCMEflIXkiFkbBys4
MQ3SFGdx6rffFr0wt9VBmLYAN7yfMKVFxnlcEkgHspxIpIlwb0AYySd36f/tXuQ4qgZcXYEfeaZC
Ofi9wU+htTtPucM68J93A7/tCwQk8EJLJSX+HzvjEUkRBJ0nGTe0Q3EapWYdkY0TcPphmHFapo0M
t+wdjreBwOablfGT4kkL/WDt3uLm9ovVUxRS69LMHN+wewmF5RDNZm8HREm6Jv6QandKVHfY30Xl
IHsxfdcALaJjAzOyJSm30uU/ZwzTOeFTlTwsschvpSyR2cJdv4VBuLogj1MtLAn/22Js2699DVvg
2DzyzxYjHFfX/OHWVSLHSZ6vCVidI67HGFYNc+tWeYGPyY3Tz5Mgpe8KgXGJG8llEWzulN7FQBcW
k045+TJc8yQh1WZEcGOMrJzS1FFk2mB2HOV63ELXXX4VSNml4WBTvybWQFRrJlGRIkpCuHqM8Mii
tooCmtezn/1sw6CaWewub0Zg18LfX6spdeG+E8ekNxGzRrIfhE3XbYMxqm+On9oj0S05Pv8jzCFj
uC9QfziaGgk+TkGXpownXI70cG6J4Hvxs0zTZm4fXDTLdFKzE1izo+igcxpNDA1mMR51yQXXTXwJ
4N65xXlfCLb7xPGSh1te4c7pSj/FhbUclLo33jzhwZ/t0dN/TscodrFoWm6gQoBgqZ75mI+wlVKN
ZmfPldyPpKMv7kg7w5NVZSfhCUSAJwhUfyTBvZO6FpJSrOBN4ArDCxtYIL9zI8Uck3dw7jqNSDmT
oYKFJapNRhOH64Ut+lWzoh4BMzI8dN9KdLjtYKbzXr4gaFyfnAqE+FXRCdiWqvBp/yDyyyKdJd96
MKhI0QoVCVT5LFqkrP+qL+MLveKEgdVTSGh6Qbt4hB8uc6QueSDf7DZNEPe2YmHFOTa3bMqjg2A9
95hV6Un8MvfGaxtHR1r3ESrBH+cOLUJfqBblJRjHtnzm4JRvIyruUFSOC6qfIt1rZRkbQUCZT8Jr
y9N5XMjdAwBCOb6tfIdXD7KOBXp2aTTISZ6YIAz015li1EvX2OlmeUJoAuz8YLljAyyGGcl2KVax
g5GTBahp0+fwScCcCf4+CuldcQIQcrw0oE8t8PqQPjl7wMJO27WCppol1MADA74f1ZdZpoQQYTGx
96LuOak6bwIDrYIW1XZokuHMGpm2zlO/QbZyzFFGiP/GOAs9+kFRC+3Cn8rCzr6/JyXGjdLN9Brp
mDs/mLBh76VVkSgEYx4Eo2w2aS1svBBvUYTwdp6Kp1sNvybxMjEe/UIlV0HXo3Kpmzhu+arQmaAD
mQ98v2e/EWVRztAFjr3zpmKXL4jx7qVIIOC/dl7PbgCUmJItM30qKtE9c/AGFLvuR4Tw1AOOMrMY
6OBUIAQ1FHoLvYyCohAfFy39xwgw7BOakGaqx/WxOgAYFHxZBhoG6Rs1ZaSQb5uzBKrS6BANvgVG
DxtNhD70mNu9chWEbyKIsL/V3kV9PTVpJMSGK2paLBLWrzXGJMjvhRXWz9Zte9BEBJ7UJQYmpB1s
EfssfM9i+MJ/e+w/2b9thWg6sT5/XAyO7R28peASxEHmPDahb3bomFH0KIkrjFhwHaWxHReZms2W
QJo2uRfkzpiZckWKAvm2JhkMSeeRWjSf45dMLXK3l1zvYr5QdPWbE6JkPdCdCgxniGNRjjDjCIif
e3pu5gQaj19SOiKjngVwYYlDtHf1rZyiCNOs+Bgmwal6bx4Qr/9F4mC4ex51Hqf6bxGaBW6hlhdl
ytz6ez+BeSZrYQ2ER1SaJUqmE1zf9woYqkuF6EFc4R6XSgEj4VgvSvMj/HDj/c9P2v84yham98N9
29iwzMrip0Hc0Tb+iqWvryNpntZ758oJ61L3VUGk4ADM78Pj3W4Z8Eu0f2Pkzk9lEaHCPqwCcyHx
m/QbaGNlp8xsoju3jUitfX2DR2fAXNBBSrxxG9tmlv2EqGdoSpkvO2SO3mhY+GcWogOlKCBPDsyb
7fyJjvZtsQScsIzPRNw8cWqR+xKiZFablzBAuruczh/u31dvLmKTnXH3G19ZpbkzGnBv6AAZsf28
J3Jaq2FkXM59R5SS6Kon54yj8BeMyxcpyIWPyt7JtofzUu+1ujELaHL8VyyQy1Rx1KeejajXJPNT
lrEMT0/wJ53vDCqYbHYJC+CX+MLNlk1myzN9EPbegLggARc4+pPOCck1PwKKXKAa0S9blIi6ozop
FKQE6ODkHz1BZCgZjVCS5WqHb0f/9t51+xX5W0S50KIR5Z+exd7s660glKBAG4yz2psJeclAGEdM
DxdSal1keyDNXbBCH8pD2wChB4CB32YomFKkeRvDSht5NDJ4gDTnwJmXX2B0AIimnBezZE0C5qcw
qzQo1LQeeL8YOWV6ikDtv9lN6484Yyu6r9+kxCwxzI3+Mwo+p3XMKYuAX/05FjHUuHXpfVyEc1/G
LByjzKDi+lvSPHiMAYzFiyzGGED6IOf5QPae/gWPXV1iCQV7FBbX47ENDlpoLluwbg65DmsgNPjv
XZMtM7shWEp1M00DQT1SxbD4gvC4cCtm/DuGXjflqM03+q4iEnA37IK0opUEdXlfVluZ4qYOHpgF
QuMdzqum+mhyraoGVMI7MzgNScq35GRUllnDn/LLhuJIfkOABbuxFwaLh+d928qApGmSr4X2LIr/
9zuzhlaXrtcEvepe31cYdoQ4+LVq8F56Zf9Hz6Y7eCV6jb/1vobUPvAt0xcMN8SIsTKiDcxtznrl
ttjYPHec9mVXT8OaqO7xP+vUffoc2miHHnlj+ZbBcBqV/sfsQLR8u7CJjapYusWtumtq/ZiT3q+h
ZLM7iTK/QXdAB3WP09j3iKeXkgIMJtbvFXVn4NSOkWgYFyoAeCjJmV8hy+hpiTrkQ/VTj2lx5DOT
MC0kT5UMPanpuax8PkcDIg8Ef1QliSqSV9zAeeGIfaLY1WT8S6cZsUiqn+XVBHsIjci1IOiTomWF
x9L4HDmEiJEo8syOmL4V/wLqaDiP92X8RhcdggVJfA3A7bZeO/mwQUvPe7INqHtmxmaM9b4bGtzD
d4OyZiUENU0VfEaPuaoh4/vQyzH6i66ubD2CgYMJf/IVquvEO6Wy5sGH9iEZZN/xnlc306bi9wdM
3q1k+bMaKdTd+vAIktzoD9kSC6GQJkDsm7mbIy0HcQFZIpe+voZ8IXwrLpZrqQ39XUzd8XzzkLpW
rUs4L5832Ctnf54jE7Sk0VWeF3c8KHPF1EqUcP0gTUjR7o3bctPKYCPdPWRpQfQWCUXvPJO6uOsj
GrUVlerWf0lLJtcLds3IbONnCKPxIe/WLphTSl+MX3Pr8mfHNUlmkBqSe7GFvjmU3YI+/HfjeM+Z
C1PzPwlEE4D6ngCokiqJmRbKwjMl7A+aJLZPZLNMeLDDF5Zh9hLRm7gXe3iPNOfInl232tzPRZVO
FY/t6e8YOa3yv3cBysNIrL6MtkZoJqUHWthF8wopVZ/w9e2HzVYuvAlg8htIjf3exly24HPH28KA
Vd+UQvUzfSm7oMpaCYV3OywBpk6J4BHhVQk23JiJXjjNakqoFS8A4JTpgkDvJ9d7sXpT/cyulxpf
FNTJ2vxWBGpkOrE6LFYryCjmNJoe04TLNNARYH/CX9EWKGQnywqlClY/SRxa767PqLHMQLvlYLLo
qmRtIAkXgHAwmDZO0zTPUAyKQkHl82hBnD6Z4SCgwZEqSwPP6ZAeUvXSksJBfYnsylIaQ7RsXqgu
0FFAp2tXHNwlmqHa69uUC7ZQVEQmOBb68eClUXD1A+IeFnODyfxVQVfFfAajMNDrjp6/S4aZkDbk
ElXGljnKqGeScm7o7+gdMW1PMhKLlO7udgwW5ce+QiMtkkxVHS1O6q9+dHdap0bG46tLSDxYBR3D
oH/onT9FmoaCOfndqx/5g8/LwuS7huKd5UBwOj14+RVxGwnKkyjiXDlCntg8uY00KRkUs5vvuXHQ
RVGreWMH3+cSat4oDy78vWAZSQGBT8cT2uEHxweXOc5TlkbxoP7fEottJKNPV4ET2zetc6wWRAKb
1sO9rdYRY6zGJUC6etgtL/C0vXwWqjianCyb9krjYLKVqZJxgGxYi1aN1wiLU1ynQWNw9i31/mQ+
w1ljosYI/H3Nu5iljBFDBlDoNkXTlGWNXI0T4CE7NrMDF3tj177vn7ZLhbwK4Wv+H3aQnV7+yCJo
sPdTLEcO8I5ZxbsP/py6CQCRbvzMJJodSCuWnyxzsZlz0RU2Ckf4VTaGEOsPUseNedr5m2G2yu+e
s9ZQt3yz1gMvBx3jR4Hva1DVipTYpNS0fpIe4hg4ZzUjI8Y+P4XZPctr562hjAPp04s1rtUueG6A
VdZc3pjfKLdRvMZtJy9zIJcAoo5uFd/BNitz205kS+6U/BOMiEopsTodMb8vMjpIf3KCVY5ut9QK
pHewFx94a4RF9jaGULQ9l4tVgkZLNj1V3Yfapj+yykHMDJUWhJzrQWiY8Rdk5CETzzxGdP7ZX6u2
2co7CBSvd/XyXl1v3qcDXg2XNomjJq/ieSMV3//gTPJi89RBwwdmNfxesDVCLvjjcLa844SSxppn
Ah+4v2r9d/XbNNA7w8FDHQVfyXHrzsVV5jPEJfDBDGQx2xo1c94Wg6cI2BNkxKeV3oOI0xMukr84
ThJl2QfBkh2tOb2egX75Lp9pJepw+gGmakMvWRiXrkFUs6Uq8BlKMeGSvVcBvNQIUYloRGqC8Boa
7BgEsOSDe1sD+SGULSOCTsruLvxRVQEFJV5O3KwZDlOCnEC/oHVWW13Ctp5v6YRse7nyie8q9M/Z
n5nRQKKoilTAtNa/dDDF2fklFXN9uVbeJ6iHUaZZY6vO+BYtO+kHGsMJqknUhJiqeRpO9bgicnc5
+jw912GRmGMU1DwBmoHQnwmCf6GUMvgCAlqRlynyaSvHrM/GQ2uPIkIrILgGgh1C5dMMoznaCt0S
iuopn5YUwYRDEwbGm/fv+9x/5VjuO3SO3sP9m7gG6HYgi2WoRvMhq6V+lkGtnVKJw9O0O6ffgcxc
iwJRf2bPmp7CoWvGyZc/4eTojHrG2Piwjh6S/74diM77yeColh5HUbiJAI7O4Z9g5qRXYMVzvnZv
C2Qm9fPtW0B+XHrO+zUoMvbsyozAwJSJKv3SbeIqzWDk2KzBgHYEffnZZ9+8GJf3OP0t8X9FNNDi
O6mkxuqobU0bHWIaffmp+RiCMXBkC+voJ9s68oG+f/tWskUlJMC0EAasId/9otz8s1oe65ec0Kid
WBcGnTe5/I6txniqloNeCzQ++j5JP0MoIvTKrmhJeuc1QdGbyqDkiX8q7cqGGWWFC99Em+Z7RQaa
c2DbYHvwlWPtINI81vxvpaBUaxe2KqBKORMTXRW1jq6mSULXqIk5OMBohNxfQcb2jPHu9zAxTMfa
aM5a46Q1OKdX9YVmYMbRmRQUxfq87u7ygF0UcY1x+kSZn891qz8Axy4tm48+yUWBKzW+9H5ZUcCB
sCU1kZoAow/AIS63KzrfG5Y61qqn6jCoor8iQk7GOnvKEfRLhhgdaQSQC251g/R4V+H7SLHoFoTZ
GsCAb6Ywl2DwzOA8YUbFj77B6uxzeIvxAB3ILYzVZkmHUOiF9XrkWbmblbxpn9DHv/tEvZXWLRqc
nj8Rh2bWz0ZOAgPEN+fIbRTSmYZHthHusBDE8j4jgDSbBWNZHOvrMApQgBF+qcz9s8IrbsD67yRb
gElylWZwaYuTGd7UzZKaQPUJYkJftZKvN+/iT7q0VRB0pcAhN7B8kBmtRmsZ8kF4Z2He4XVN/ZIX
Vs87JcMOw4MQ0dP26GbIlufbVGiv78vnvlbbXhjzKxdcKIe54w1KgFQrWylQa6s2pvBwcv+caxKD
Eybv4JDJ6RLX0RJziG9fWq698eSBW+v2Wxd74xnDw+1PC7wT0H7VvoysWBFfmR1PVTuhnssXaiv8
Vl3Ta9hDNBRAyN5DQvtyQH7oeizfTXc5XZFWlVljymyW28sKVxBxdcfW5DWiU7jIi58ZkDek2PRT
fKx6OOyLWmE6KF2D2XkGsKPHtiC6Sq+66sBbUS9hHVV7NZiaRKCr9X8uJBKFVEwsk/JBDpUlhL/1
veeqrXUPIAnTNtfl2qq0TLGjjttI2WPzUf16QhcnTUftPEcOSZ4NCrjhmasJpCF0CEI/A+PQuuhl
JdPRb2QIkq/kzvnH1Rl+41VBS12it+oJaE1J+aXuMODOOtSp4ocp2c6FS8pUBIyCZLyS1ERHCDV/
bsKZcgDJwhCFJFITC+1aBB0xVYd3R4eson7KnHLUYhfx25KeNBBZOQ+GOtuPAE9wlIMK7RuxGbfg
iQS3TdLjDBcb5c22GGmjFj6WOAvxZ442ZcTYyxIffEg8PKPZWPVo9E6HO41hIWwfxAfevgKJJYQk
aStqx1LOCysuShROoTx0Yq2hgkXVhqxPElr+TxQV+QrRBqPV82IzUwy+aabZOGUGZtFc9bv2QV27
8Zt91qWU/UCjUsiJ1qidwaoFuNBDlKZfPbnFPYnOX84MRzC7dfPeZniqNg4WALiTHsf4cwABNO4G
cCe0j6xy/WJrtkmgR+oLyK65t0bc1BRxHg6pvXX/ug2daCfPXl6fz9GZYTjzvO+MmuR7ktJr1oK+
E0eo0Di73bo0sgoeVusM/2LJEyZUcMl8YuatW/zlrSCKf7dOcqLwb5tTDbiajN0tzXZS14EzR6kQ
gEp3rx4tj63W23nLYFsNUJtZQEm2jEXyeBzx+V8aQbEtiKjW/R3ratqjs3eZrMT6GBnGNn4avh8d
WdQuQCOhx18Rcj9rt1jEDodeNN0o+0GFKdaujMyke5JPcxhcuGRkjS5kjR982CfCEB4fweIPOQNG
o7EWiEF9lY0Kv3yW6FBEOoIG83q2jsf8sa1KZETfNhuKTpfrJOzH7DvchHijhfFWLX/1lYKm8LXg
vPcjGU81wRlYZZAEftuFNGe54qkEfv8XKaOBU2K0vrjxzX9ip8JhF7NLctfVlDZrrniinRM+XQ/C
VxslFDdFX/gayjCQLmug2RwE40vjvCp1kUb+Hinaesz3PNwc4D/x4fzhCmkzxEouEP3FMQdW+saC
TwqHKhpG5wqN9Dheff3Igcn0F3cjjolWL4eOgew97iNEsbsBfBlh9qQAUHL3hztWXiNrZ/C6BcIp
x//r6no1r/5PX1zyEoVHZImyk1k5yjshQ59W3iknb5IVwqTLWr24dSe5bcY67F34tkX9LgvhBne2
u4MdIj2efXaDQ9Prq+KKNN7H6JRE3s200458XKN1ylBx0oCjp04Kj5ANAnKBYhCAgO9gxWbgGbDj
70X5fYxgWcmR1Bi6ATSOQX4t7lbmRZo5HtOL3/Vx4mMZjDUU665RnbqWpzVzImwYLgLtjn0LMlBR
3xaTky8/E3vyiYqBaopC24w7SZ4WoHGTR5WeBdj8LWHUJfIMxvG9UxDtXqMI3W4sn+XZ9CxSlqH6
aCiaCFUyZ1gvJa/d5ZDYKE/dJQv8byaeT+OaDHWPUKpL7zyXoScsrTOscKY4Z1Wpjy48hCmLQ1Fo
n0VZOiGdDvBKfsNPSC9ZdHfu/gjFbbW2jImbBRbwfUn93w2bkZJDzZRkSw13XdceG8J+BCv5q+2k
Sl78oLuJKcMirqLO0iNr56H2n7Yg2XfxdnaktYdd17fYgL8LYbRzXQAyJsB+OdqfLN2k9JeZD6uG
gQjlOM88dM5+/1pFf5qDzVTM2YMc2xFwn/0oxtC5/b7sKa3apBJsA7O0kNF2HNZC6Frbk8g7xbZu
Ia1FfG1O3k6HdHSHhuIjpMM6YR+fdBuPa6uEbQNMj+x99C+K7iJ0rRR25w0LBHZS7UAeHnY9kBi3
VEOq+91d6z/dUMF5F8+USV7uFZHJCjRwO4YDvGhIuflU83WwaHR5xTYBP8P9CZB9Dn0seNCssLTY
MnPI6tTieixVDS8/WUIuo1Mzn1eeREs7yHbxcj/We9gxYfNLP2C1V/kd+mb7/aOCt/Cc9Z9Po613
td7qWCjoonMmWa5xuiEYI7oNpM0OxqcCLifRKMucjT7zjC6B1Tf5ci4IFqNiSNdPi8lo259ZiXF1
jI62ejMH+PuGhXQ13p+9ZdelC9fNButLgjUqAkDySp0Wbbsrj8JDxDIB//f29N9b3KWoctNwEY2/
doeP4TRxLmH9cbPkEh5uTt34f+7zb2Xn6bNmVcKAURJ+S6Ie5aCRfiUJJy4XhifM4NlXKshp9xAc
1zeQ+Tu04QbRqdTEoSkoLs5UofjJam+4i5+GpOg9EPTcMeL32tTmNIzmFG21+D81aS4P1PnmhXc5
gbChD3W16VUdLG6JlJzRH2k7jA8zPct9EFzqxZe7dWd47pwIi7DMqd8bj4BKFQqoAMBV+i6kXLSt
yI4wbfWBAJaWpshEBgn1ibVFmADkkAw01exuFqxfr0f7W4dbl8wKvWz/6HSe5HW/onZ2yJPPiDmg
86S3QdI/hrpYZMbFyKoW/qUpawrHLTbtbRvJTNx9+3gY8xMsMVAiMKMuBSj9r2NHfZEhL2BMwwzI
cwaZO1O0wFCuMSBSyJMmLq8YS6gtLX8xBN0dA7V/teV9SqN3e3KBO9dNzEiCTXYiXB1lQUGMoP5s
ZZp3tEkJJFJ1q0xRGgcLXriXNHg9DjegZ24Lg/I5wGfZmORhd9IIzswDlXHWhRpSv5AFToh/7+3O
LUwtJVFQQehePsJwqEjCtqj/SylZRglafXd6skJH/Z4AWOFBwSZ0Duog1oo7FNBznmuPJFuLgdVD
VgvMfbIWY2Y3R3v+2TJDLHiAwGJbuN+LR4W1v1FWyoPy2XmadZ8t86w+2h4r34v5ZXxW8OcHYNTL
BpHoiSIvJb+NxkmDJ8+G+GMDalmJqmnoqMptmjhBWd/FokL9zbZfXvAN07Z7BXKdo5/lK6vSK+Lx
LnayzeXQFZNJWw190+vPkyQSCTV23VUOEw2dyz3MP2pEOdIW80MWObNG5z3MHnJlzPGZpy6sv6w8
aofcKXjT35bsbacbDtFE8JFp01ye1ILty7fLgest1dyM7Q17VfyFx89n3yrXZfx12ks9Z4Er5SHW
Xj5Ixrovp2F/5zAymmv5QPWc4QGfshfCAk0xJDu9UVX8bzCLSiprHN/oZHHCQd5RiDzE9vC1eRLw
gL97h6KXQGMdpP22Qvu/1iy+bec/pq5oEbgZ3OKuG5h/h/mpu1W3UB0ifLzweGgy33fsLOgseNe5
I16iYbv9GB/YX1QKqZ2uUHbvaarLjyR9wWiAJt4p1zG92VJV0/7ovElp8wugoxJEYw3ElASJ9t7r
FIRh79zkQr0IM8tWQdF38OZK7wTs05vVzalzUNNKMO03egL3CknfKck+AJ/lryyjiD3gBxbK8032
8z4YSyxCeXa7eMmgDkVZxUP4KJrHepZbMthOV2ZXOB4vfbpK88vlq+wppLFaZH5H7+DY7qeU325U
QQSkRVABTvq8eYiGmNbRS1o4JAFF/pRmw6erzJNsl/7/mfDZRjKZiWfJZZkdPqvCUsXC4uMbONNM
e9Qs1qB7V72AHBuAFsHtvmMhDXnWCJ46G7E5Lt8nWawCVcOeO8/5AB2rEyyfNxnPdclB7h/FQ/GF
it9Qzt8eau9reSQGpJGvd5fldVhS51wfs76vZ11Pk1/Wik4hXdPYcojVWDC5DeHFN34+tiYcCiFk
sWiJ+Ourm+l6Sw/c2rH/ZVXllpTLzXj+QzoWZ4VjZAsfZj1M4kKkzAu1/HD5z8PNVqUmAZcEyKgA
PtVkLWQ+tz6V+lgajQChZ8Kd0ihDde+WcAVMuwYcQtkiDQxNyitPEiUXu/SPOz+SiqXDaowYRScI
nr1TBfNq3uH9OyvFoJCZ4OknmiEMkRYi50aAgz1B2ZwLMxRfRDA6Ju7cMOjsziYokqta07fc86Xt
J87Sbk8Be/ZjLyYjimjLs5eYOCxMUBesIXL73gqa9kkzopEACKA1EnOSeIQ+Rii82h2TsDDzWXeb
cdozdomUTj1vsEUrJd0/QmilDuNFYPlJa/ATSkNRyaAsrnz7DMQvvNm6FaiQTlZkDAv+kQSWD7Tg
4fsUYu+qhk/anFHd27eZysEg7Omm4/UIxhAWCT9NPVeB64UX+7xu0TXkUqSs4t9s8ZMwDWJh1KKw
oDoyLZH+iuq6GmWFEBOIGaYrmZeJs4//1OH46WjWFAtusH/7x1WWSFelUEX/o0NDOcalSQ5SaRUN
pOp+VK06FQjkMO6hN8ePyMTbVtcvvSknAfJ0q95Ae2EW86AH+icfVwoYg2aQdTg7K1UbZiqE8pDC
4c60lEo9MiNhsSuOcwlYyCpZYv4JQ0QuhG0co740h5kkKQvXmT7VhK24SD3RBYT4HarpkYLcAwtl
5TEzpCgPfUDrdpS0FLu2I4oN+7p9qmsPm0VZCQ8df7IGvBdGWNwygCyKREE3/7gledryWlHBXTeU
1IKbE2P0D1VMlKjU33K+Fzu2z3QtQZR1Egm1XrMyHV6Kl64gWJDAoVlBHOSaVXyKd+fL3+CR/3Vs
LxVslaV4IW1qVihB7fQzVTb1XkNBnhQMeRiZySmtOySvGM2GzckcWRQ6M4l/8CqxaRPSuH587jvD
r4d1fkHj73KukL/Qcgh2UAM/74J7MbCeh4l4lF8rMGrKc3KvHZ9mNw0EggNRMjBTRmgwIYbYzbB8
nZC8sBq6Np0s2C5Jy9CbVf8oi477GAeQhZGhUUAcTSBzyha4dIGAtGCS+pPmAL9URfC9HATcVHm7
OpB5fKJWb+cbQFzxQJsa0caP+9gphdG11puT0W9gOJ3/YNz/a8qdsvb+9Ty4qK+3bXwVFUJghWeE
0Xo727grLHglW1uUXd5g5MOhQbe9DBlD0Al1WWAQsl2xKFLOfYSLo3dMiOYunHIq8DuHFMEinKUv
/t5ZB+cHnsFKkCH9yL9hYB4hVEYQdoi5we6h+tR9lolEDD8lA/HV/i/0dGcG6rIU7jYbgCnYwjVL
UQ5hXPNf9XNtv3mVrPmYtUKIoA3yzkGay9gzxteu+dHm86rOqgDGRhrHYOc7rsTgUq2xgsarsdFU
wl03iLQ6R9FrYnsEVg/hXrACfAj76Lc6uvOZyTXv+JpvHbbI9wj6+Nv4TWemWGZ3oBDHrvHoqX7u
NDAZAtougGz3Oj+M8lSxK5zExoS2Q5UEk37Ao01a+4MuhT/iE+C6itBrkBNfulZYwErqujK0ZRwI
tKLEhhSC91mFujoN46sjIqwchDMbTAWuIvfiAZzw7tUEaMIq24fv4RaLbX0FDzKek+rj9iClS5jU
xE19gWQMwyQg2/fPwKeOCQEtbMPl6jZNpA/IM2I18isO9+ums+KJWA/FYKyfSxtCkWJBdMX9oks3
2ZUgVvZLXoG3iMyx1FYLnU02RWeFQHPym4bLfnpWaMXNNoiF15FHqWnmW1fxxmwyc89CPUxNZs5p
mVR5V8A3Mozk3f638eXYYguj4FcHscJre93LiCuMRGyA7V5vNuw2Vv7eJpt07yyXqdXJr/1V5fKs
eB8/MDv8r5eKuLT4RItztL4E52xar6rRZeQUOcg4utqrq8F1LDc28rLGVLWm4mG1Uv7yIFEaaiL3
xjtgAKRwUSAjdJYzaZj6Cy4QQkqg9FRVG2SPrRJHRfAzkUDZTRFU9zQXN8i+eMk7rxuP+Fn8EgSe
zPHRIbuK0aKW7kEjz/8Kr0mgCpkVI0N8MYH93iVQYp45K6Oz0CbKzf3phkVZ7nsiDy4d9rvFf9ws
fGBDM99h8hw7E+SY3WJ1yktHybcZBUtyKBVRGPAR5IDyu+8N88muSJYri7KbLlUq3vtA824/HDaF
6jr5ZuNBjpcvIIuQXtReB4iipQiLcTK0UWIEPz7RwS5B0bjgCFik6KD6zxcWtxTUTZwI3gNZ04ld
j3Lc/8l0k5NjvE9HsNPVqPMGqP2oBXL1JTk3/DqtZ8ElhomJ3/O6S05pPFkCH605rync0CYiOYpv
rckwP1xXkFeXuPRLXxs142DKjAfWm/eb1+rf3gA8r4Skh7XPA72iWikVYNF0HbC3CULD3fkUMUDH
a0LXYnGX2GWUEFxsH1/Yx2DH68spFVeYz1W9Hoxp+hrX23x/LWiHmW+nrZ80OfZ7WSzCAIRS7uG/
rr9PLErElEKMkBMX5jpeWBQ7zj+LQt2xAa3MMO73wVE/l2Ue4Ko+KMbHOtQHY2hOP5uJZRMytZMh
d3APiW+WtZ0LWR0aSxIZfW7P0pzVIs4dN/dnyLFrTtM3gGfzaaQD9Tw+fLXb4HhezlhbZtojf0Vl
uVhMUIUj8AJtTPfjah+pSyWt4N0ZZrsKZu5TaOYVEWNcqYC73NxemHYl32ToEYHq+8Erwlu+rR4O
xRyhjr+kmCuonTuV51SCQ9Aocm9mpMdCWmnEAJ5cww+v5tfEniE5V3kgIrN+Zo1f0LRbMvHNOALH
EhgkofT27UCzhYLUCL08J/n/R0MMrxcRHNLaGyO7aeQvylKdv1BlY2wl6MwW0GShRtyOBrf8zMrr
vMkqQv/F8M6BsJW7Uwgd7/k7szDAppzrD1orjWbH9tz5UExu7FS6w8YyObWMOXP8NWiKZR7kvOVD
xpbf9Y1aoElpAZbxAmEJhm0/ob/VBm6VVpdF3kY2LnFOJsGAar9VDfh3cKUgXV8E+0KPM9VsdwCs
GpmRSB+U8IXPs1XrZ43BqeZLXiAptDqKPwugnReLoejga3H5W7lgtiLX+kFgGmq6/yYrK17drcpB
l9L8MEKxHrNmjaazGIGzSJHYQA8kUt3kxsYIj6Fv3JOZsPW9RQZTM9N9cjBC/+3E9iY/8Qj+Iwji
1r4WXkw0ib3BuHV62YNMaRg4ZjENlI2WZnacmmfh9j6zrWdVEKbpbp9Objbt2enZx6bsyazehzVt
lo96VjcOGa48sSyFjllOVXCZbDJkWEiPEsd3eL7iwHGiq17GbT4YZbLiIFSCH2YkVBNREXl1EElC
yOeCdo7o5GNsQNBMoc8Vi8rHSgdbrhYigAX5p3vBGX9OW51+TAOxH7PtogqXtnPA4AvpAo7jGf7A
FDslOt0Ujj9hhdfx0TRnP2tjRF3e2n4jhXyRJlUFn+wqJ/aPNwsJQ0sQgZKPAxSyEZs/HFlndINp
/aW0EiHmQWy7UJXaQ8VHkgm/xnhuT3tJxQ1U/kOeXbAs1jacTVcgKdybVKbj5XM+6026eUm0MdmA
slLv4OPX31/ULdTuzclYdGDyQO2na1ll+712vTNaCyDNB70De33tLuqWrJpq7hVQqUch+d77slYY
EkozYQIbJoFRkTVGfjywzRaZg1Kmb4uK51k/PbdFXIOhRxGsxwP3JDDTl2gnNJ4NXeSvHXIehP8W
hzEe0HDhR+NoBTdFFoUt5nhosHLs4QE3ljfa6sJ/gJAxVIsKta1LGO3vKjiFtyR1JY1IkA5Me3pK
oot6FwusyaAX0LLNYTC3JC/rw7B2AEp9xSFaAODMdki0+vUyHt9VemVYwNs3+DtU2LceZl8XGchq
TyNdFE3DLBfeWjD0NJ7VKozsG53aK7GGGahe2+TTWB2QpeGbL6iiS5+b6qG2k6t+F724O4uLJyhq
emVE+ad10jTjE4vLwqAWRV7kKEsFHTojjPUhA5a/5NotM2ef1Lp6zKJBUcVXnndF/v5GYw5kcdHh
eBgsNNlkXC6tHUqsMKtXs1DcNTi9t8xJgfj/rIijg6/g0FPvlwi3QRbRVejzVmBP5kzEK3I2vOJC
ZFdlQWHcp1ZgFXhC0M38C0773vvBi0O3+Y9kDQRGYBvHdd2alZo4Ck4PYSvjB+uBMmzU6Dvuxees
DmlaWjRT0NeJv08590OWP/+knB8XYnZH3NNaDJIjHzL+kv86cZDoGSTOGjRutPy09KJVHd/6pbUw
Wik6UKPeJ2fXTYaT4lB3PF6xBKXTha3lyXUBY895Eq86wa9DCvItjfdRDYnIFRKKLEfM83FbFxP7
lUr4fzxmtMx7VFxGOJfyOjfSXQ8ye/SuIBt4vzjsU1SGAu7NadubATdetT6MF5cn6pwPX4ab7gCM
XE0awP38HnIcLm9aJxmTg+4JWg2Ehbjl36tYzgJhhOdWAXPs7SFuUs8OlvH5EyTVThuAOn6ts6QK
6f1dm5n8zCUGgnpsJmXvlC5NDNWsbfmBaV/SICStgXcDdI1v95HaY7y6K2lNK24fKCKFcI/6DzOC
Y3XPe1TMYdoj4DD39LyoC/cHJxAzmB1x4t304N4kiQjduLmp7XpAxJxQrufOi7skX0gjoFUO5u2J
w6sGshLVS8NZhGn0oRZlrUlk2vsfJMPGVlO4pItHb5P+HVFXD2xhPOZ+AhanLqRXJ1r5u2OxHAOM
l0xxsZAIUTvcYH5r6NYx9L79NhtEpSU1KXt8PYnyVtAq9vB6PrcC54r6TMqNUW5/hro23ZhH83Sj
55moS7zMkUY9wZ2VlmcFrKoxUsVPJIL6fCPf7odgqWXLpAM5bY4hnBIzUOxkCx3me6XC6OLakOIx
Czdet6mvGxgH6NtHs4cSkbkrFjACJhw4c2GapiqaiVjaX/vjNMLbn6/T/JxsBUIIDfr0pNjHdQU1
f7xq2Pr0g9P1Dm4gOHGeEjR759AVmqlcb6URbCm2YQbD0E+hQFCLgzfbJup3z0E6Fq4Fq8sUyyOR
31W3KXBx5NwpxcDRPXFNaF+nmzBkw1HSmjeUYvdE+DN0C3rnC8Q5p/hVv0joIq//rEzKNRjlCXjM
TI0oaqPj1+TcQbscvXYvDihbHHcTSAkX+h5bzYQKAQz4vhNsJxdvsmvVzAsxUniUj0TZgiHSYkce
xsId0Avwumjlu8RANsRYqfE1Y9FE9uNfsi73a/g0SioCADH7TPgVUitkHawpgILMZYHKqbEfsUJd
+ABADaaqVVUrhCixuXtBlryoZwcY4PFNkmCSa1s5yjAUsrmldAa5txy4AGmoWtKEVu4tkvdod1ey
863Pk+gPsYoCBuThB/lWvGy8mIZvsfXeQ1htev5kbKj+t4QDyrIpjNDVHbafYPMm9tPYJewB1hAL
A+6qmKXDze2/tQUGNCZfijTwVHKCWSH931udeIew1Ki9iXcglIW5wiv2vqH/zm0Gy2yWupDWlMrX
BbtKCPu4J8DEBz8XzyJlxYjKHN+PxND0ubB2ftIyPBCmSGcbaHvf7mbIX+HJaVXvnJfTeUrRi6gE
TqW5tAmfwqd2IWq+OijSUh4dopPkuovZ0kK3tLkdbdAo53OWoUzgCQAc1Biz7tCZWB80PQrO8OaT
HR7mWgQR5hPPvRd8fTycJd2WrzYcrBf6yciU1ypmiZuun+oTRD2j776umhKHVI7H3O0/Hjk2M9Eq
NZXBEwIE8qKVuFnc5jBAQGlXtaKl11fIAxqWQTuqsUldhAhwihmoyzsfPGFsDvld5unBWz0AGwHh
MRf1yR5Iel7TJ2uO+vjiHOlaZASBLReWoJP2eVWWXLzvKzNveN73nPizv7AmuQqxIqhft7Vw0wqb
SQlmrHSZpEM+XeTn7eRs54g/lAoqHLkN0fq8izW55ZXTDGK7jk4fqaf2X5pbsIEBnB6PW+ZCFMVq
gzpsMyj+Jqwvrd+NQKqmxC4ae/+qU3JZoCAlsLsmFIJTnzMi4XpziEtJCpp/n/dSpV9cEbuDbJMM
wuP2/4EmJhZQnPSPTgQaBhkdxg59G2dBXEtAbDbi+eZLX8KR+Y/xPvqr0gahQwy7k2ZrPULGmul7
8DaK6HdHvf9YdcK5+RvcdG+elHVU/LXO1TEF66nAsK4b0IXVYolu5QnqcQZIjOp9MsBsCHAnXt9c
vbhdJG2lCMbYn2NuqUlDZJzd2MGPq8fV6CWcsFPezlm678hrtmX+nGC/oQzh787OVXIxmbgTGpP/
MkTDf/eFq5I8HxSMHNnl5T1JHtyKQ1mYXe9Gj8rX+ke0SYgnkvT9aGrWw17l1v+IUQg1IjODaPWm
snWmgRZzGpv+6O08V9tTJYGS7f87pqQBjoj01+Xnror/Iy5m5+hqKCxvjEBqplo4Nd3SzUHPZy1z
DezlI2EuweB3hytgBeccOe1WA/RBQGIl8b5ouzGx5TGfl9OoWvwo39QhpEqqbFUKktFDDi4jt7vy
5+V/O69DhspU5PtqjOXE9x4msJT1zaOxtKJxmeo4ZXNWnjFNqKaySWoywlpwSiKdBjXgcMPOUXlp
pmVmAQ6+efVUwmulhPtOm1a5YxqrMGzj06z3+UQrs/UCx7t3UglVteH2Ic/i7L57b3n+1yheAp7l
D3xzr4qn2xgUFTLh67DAhOMdnCnjVL6MB769gh07TAxzHdcad564cDyvqD4jkskBN9GUV4HsgoGB
FU3epEhDZtZ3rFRHpEVirKckhwmu/7f4kSldmIY/hJ6sFgxfIxWFTBLFGGz9r6wjjCNs7/8vYu0U
RygJYShz4oThREvQ/QjRvc6rIwRIOm28EOHqC9RKE+4qFbKRyicGr0T9rwfa9lspmNTjEusoWWWz
CTAAjqPzxntnSkYU15gcwjgDLt1a+Fy1avhBzYDgJdO/9Cr+a4O/ybDUcNNZURdZXWiYSM4Baq/Q
VL4XCPP3sZ4z7Wlme8efXrH7ahPon9PwILUdGxC1KhsxHrV2mcZnqm8Z/ci1YplU+oWOnMUtQVWm
wrRe7M6D0w1kd60L5lH7MTR7eHE+yDyxxg9QmI4f9VAcy5W7LWFIm4QYliA+nWqWTN7bHBCPfizL
/fhLAImwKeetqizuDXfNKtg0lDNDtOwtcBNZ7XHVpGc3lGPQkMIUydpAjR9h+L6LFHrTODMTQAbF
RktY4LXc/QJxx2ZVJgzn8HmIcrwb9iqa96uBnGkJ4n6a4K5+8SvPs+GQmnnlIaVjZ/MR/Y2o5+H7
eGQVC736e1/8QdRm49QwJZNe+kKQwro2x/3BwNv9v0guAKDtLSssV27Fvx6VtJfYdBJM8iZATAar
IhsXNc6g3HlCKAjTndzxWEsha3uE+uZDxkSJMyHwPjgbeKrf2DX6Q8nIvvTCXv0tBbDR+bDUqips
ohfpLwuv0dI9DMqwYwEE8Zw4rBLpZvI7+mimesoVNw2rHU2+Gsr/wYcNyeTpkZmjTSZ8XjMgjrYG
WMM2wrWKPt3DEakeYmzJN7dwl/QiIGelgllB7iNX7lat6aGVl3DJ06ibJX5BzN6Ys5uYKcBHOZyw
VHnvUkljMWY7+/m+WxI75uvEDUVSCG5hLH29/ExsyjGUktQmLTUGcYHT2100UY7NSzIz+lHvTm6l
8wdQvQZuVKWHKMojb2tpyIm+x1FmJfsUixLu8ZE6DIMYYePW/TtYo5YILrixs1k2HH3VNKPjkLiS
ohy2+1FBrAefIK4k/TCUQDmJtcF3gR0VNd6LROKkMuasy1p1pbFVLXQ17Iv2f8MSd1jcM1qYpCS9
MdawSFwtyDEUiIKEfv49nOpDXk+GtyhXA4w8k7JVJz36G9cRLL0lWkXR+chUQ9OZFCmIsE0tmnAp
F4BCeGY11bxaIBOSKss2zC0BDlISF3k6DbmpctHU6SJfltLM+o/MX3yd7qvV8kP54nkUXkswxNdn
ccJoL2e6Q6QgYltoAtBXkki5ewVlOQxBsfKyz7JdvvwP0OOaE1W0K85eGc7qvk915GjmDbK5BPFg
RP68s+oqp7KLrr2GF9x7TFbETFTdKsOf76/6f0qdsxCGw5tMIte3GTKKtTpkJgXD2Z2LBPSqpad8
MgFsj2uZ53En9uVD9TIlKI38iwJA68MMGC4amua4MOjhER4OV9nfRXLqAnmdNgjZgzf0IGSwd2MD
xyztyJ+xkIKs4owpm5YfYXTHlF9jP2DRvkr+UhTCb1VLZ8EEgIkwGPWQVLNgjGZDyH+mHnvoH3Rf
dtjPu7DX1XvqppiCR+gNnihP2J9OqODjmpAzKanfFgz4QpLT9GjKjvWjrkU1G0J78tDUiBRNa5xy
i16/v6gzIP1Xaw5R8SjNdoT/AVyNvExeY9W/9K1bTmAs35OQz5NcchNH3uqWi22HSMWWC7+DBjg+
8/HrLWeMHtYU3oy2hrWQC93V379+gWhhkw7j553vM1soiDPe960cFXkUYrvOi6z3ANPFl5oHmuNE
LhXJ/NxqyYYX5SYpwOjQWucV5tO3DZcRjCgPIpICY2IwegWrxa5wBnkfnGt5xZTQVHWtf3TyZvay
iYKoDbXBKg1iP2IjH/p9BZCLr8Z5jLQ5/aQjKdp/tVnmu64yjm9Nro7eDIFufGz4Lsomol/f+1G8
ztJpPgnMt9VPrvtfPumJTxcPAALo/HdKPfqE49uJbSYMqdPsDGGXYTIBGlmE5b6RXVqqW4QHRT0s
ObCNy/H8bBIzaooGQFpQ/7qBfdw1C+0JbkSrNF5Arrz2ELI8tfdpsk6aqR2ZO7ecVq4oGIIunlSv
8OZIxDKKXiUQkFvTMcbvepMAanKDsfBpbVEDxbzooHh6AEDGH33en0fue7Cg5WPnoH+MgUQb+D87
s3/l4M0fKf33Uysw4VXF3BQ6+4nVIADAXiA0br098gXa9Ju+qdtz8wcQI2RbjCtmOaKpWF2GOe/R
PAjTm57M/JNtycEue+cWglT/lWABuB5f0SC2r7XptzX4wLAAbqHxox5+pi3M4JcpCfJ0u2KmjM5B
YFLP7QexI50waKPrqb/9+hROIYKacZl3OAAfQnpESquiAYir2bKYb25ocW1OZjKQVB/XiXN2OVkd
QaqWsTycP0DAH7ixyQvwq1MdmKLrRf6nK1WLEF64dY3oKz6r2IyHPFhEq14ivvt8InoEXa3ivA17
hM/wAPcCwnfeKwoi2CZ6oo0ejt1tnuXpdPT9IJZZhORhPqoyECF+avdXlxHdWVTVG1Gcl0+Bgu4O
YW3opyBoRtBCpyfLjWzRTbUW1/wcbkNh/lUEkPNpm3jhi3Jt7hQuCo5aGEKw6h7IcZHEE8lj+Vcp
d9+ejIIDUjMfQPy81lN9WbsESFBzpX30C1HoThs8V9NeYPKKykM9+obLqr2H8SzSqKM60qyEC0Lc
xKsJmt9K8SAXEl4C2WCEXhUIdtPT2CL5q3J4AGh3L84l3WhVRud6Jn8ma8dVbwz7HsgaIo6VyGnk
na7rF7SUrPyCZoGnaPPI681qB3AcDTGsNSetljYALbqrQk+5IhGVAvSd8/grlD61ZctJYs6+Qyrs
dGCTHMZhoqtOUTWp5Ke8Y7u1ci52ivcfWctZv2QgpEUwJuo61dWgjhBaRpcnKIkDhZ+q5wcS8Jvi
kFJ8HaeVeKF8LgIF3ndqTmyP58cT6p1f3Cga2jgWgS35wUD1M6hKEzdsk1AyFk0pMVBkW0s5Od2s
BXpVKU15ocuWVUlHd3Obml1D4Yk/g5MLAbByxsmFRxwNYnitIMQlqyDBPOBRlGdb52rXcitWEyl1
Wy1kjb42K86uh9Dj+SvBh98bQiyohOdS58pHE8C7RW0eITU2QbLVaWkJRKsVI/6iFFIOlKUNUgTm
YI/N5O4N1ElFBCgq+qP7qorjUZfkTMbi2VrgViHQdWBJms+f51520izDCXQhIBvi8JmcDYgzgaRu
qm5R2hPsJWGBAAqJDRF9Cl6/hr0eN4K7w3Y66pvoRJlFATfzEfYzON4Yv0/F5CbUah3LGHDkhPdS
aDdFPM/hC9bTOgRaknOuvtVHWnH1ipeM4svSPy6UsFkCFgOFBUoXbSClB8Gg6Y0baSk0ocfkSaU7
e2DaPUkGdEouIrMhopiooPGDQOxh6HiQBdu5JJc1n4rHMmJLZvkvKID6EW6cqqmIel8qSBB0wKJ/
7rGFu1wszQl8WYxb1RlCBjFhhERSyiV2ukfU0GsP2DhZouOWpI4+q/20VAztO4zNrfr5tZniAIF1
ZFRo7k9G2KqzI4nnfsuOl6w051SmqnNUzlOZhnAZ7QHOYvTtiB02NEtpIDZCldDUkrZhU4a6wtNQ
Mq6UzekBXSOT0J4SCuDQWCddd6zx3E2JaLviMwrfQakSGBhc95NcZixJAk1TipCgLR7z8g87pQiK
blrJFNsUT3n/FMtgOsyWPpD3qTYWu20KQYKk9fFoLyeYKKnZ/uA4Cywpn0qv7bvsKBOEdSOmeSEl
j/kAMiUQY77w1UnNrr0UuK5jL33VZjiXJe9qq8aF6IFbePrRakpw2YMwvwS9gtE6LZ2pTHuofVe5
m3RSn1t4+Woixe1ldNUNQakfsehr714Wj7NqA5uG5hALZ1diGKzSzecqsmyVp/cATS8rXJXmQhOd
vaodJyP9KFoh3EHQBNFWlztickGzwE4j7Puk1IReZPH20pkOFN+2cghUsl0EYA3sNZkwEVsYiG2/
eQssf8r3xckNh4E/aNZJUAICnLkl4JqsMihryMn9NW8nHpztJ1pPGwl8yewGbtPWUqaP5M+/pZJZ
BEdEs++GCFWFP+q5hNQSGHTQkVRkQQDOf3B8/y2YH6xjGoLsIJ99CYE0+31pxlEkq3pdni2LB+7S
b72Gf5baQHoro4MOP0REMlO0m1oFS/bwyuhbYewnNPmAEBEPpgf1Nbh+xrjBFJlG2XrjFMbR7nsY
285Dp1tzAbYa4AT/xccFsibfyVcqXIgQvMbeO0E13fk9hJBOuTvjVkG0C1WaQEsLKD0nyxhkYBiO
SKttkshSIQ+/8FPQpMZyoLbxLg5STIiYKd23yqAJ4ssAdWl5Ex/wj+hknegOCOO17e8mbJWpob+H
XEpcfJ30QK6P3YIX35apR1EOAIs7B7j3Yc67YSfs7RFe6UkamBo1k6HbOP5O1SwxdHDZ4A2Td0YX
Bn0QAvTbwMbdrO8AqBV/7eFDHx0oBMkJnCe6qi5QtWuXMxHO0Trvrv3kDfNOT50YjODhdCgyQgYN
sPLfDYvlkKX2FMBzU05ayEZ2cRit3jWUNrOGtZ1Idy/J+iJwB3Q9RYVuYUQr7saXOUSXBP4c8GaM
QPlLERGPOH0HLk9Z95Ttvuj08yN2eBBg23gAdv/NN7wMH5mWSRKsvMJEParGpMAy+82p0SXhlW0c
JKQVhOQBj0F/tp2f6dbh94ZUQG8fW1K40T/hz8ZhqoYgSf9wI25h52YxSATW2M8Avrt1m7bop66G
kooUFU5RYcxcfe4GxyaodZorPcrzBwXQAd4pHKXPzjw+9JdxFTxz4tv1D0k8u6aAuC5ieEHSHqfk
E07xH6DcvtlHNc8hP61KwiqFyYVq0VqHc8CYymfHiUSZfx0ZDQRITPECsfn1IAG7PMyDL6kcqlWZ
usGKTCl5u07B61q/RbV3GknrIUPjCB5PJ950QYXnGJPdIgQUq20K1TqIQIE1ESRQ7dITeptX9tJq
HJ55TrxwR5o9n1GSEGOmMpkuuEpgvDXS1CVeUlZBQBDaqA3H/sVOq5ggTv0sd0gcp+CwC+YdjCuv
kw2URw4RlpDMpTm6o+3BCzbNFnIOCKBn5c08t5gY0NS+oy3leMaHu9PvH7fjM7MknguuSKVVKuNa
tkqA3xQygsZvN46GuhReBoiTCv2MV7F3ig2odif1ztLBf6cMNNdPL3n0r+P8nf+R32AmjTNqaErW
b5uzQ5IXwfRVHDQEBj301xLjqegER2/NBQZz/VkLy/YOhWWY6GnzHQXn+bi9AlfoNCzynOwGx568
u6kCVRH30x9cvFnBD08p8J8BQ43D6pB+h/vh6Aq9xpx+O3jJOWsrza4ekxTms0K8Esob204/jFsK
qUHg9E84mbrma09lGZ9J5MEa/ZJdQIA8ixVCbdrw97qrn349ARjWWpdwdNcoTxIoF2hAkyRuyqxu
v75aNilcCJWEadierarBJKiCbOANBN+eq/ngRhDi5cWWmAaWgu+7+va4MxqSEe4BmEPmKpikFSZm
TZoRyQ7DDRfAenFMaFoZg0FZZDZ4son03StSc/Wha32Kfu3LGzJrISxxpnct/V4zELMUdg9EIQ8D
Mq/ALd5PusoIrPRL/4qq1erEa6uZNxiD6madZWR66CJ5Epw2lkfGYlcUgzZqMoJt6sNkZ/a1oh81
NFfIJM8dEqjLShmRrFZOrC0z0JsaYuNwpk3h802n2O5fd9QpPtQQDKPsHDSDAc71VYVSpE+S6mfT
+FHApQks7KiYxmnsaI5bypQdQ550r37EB+Z1HzPcsJpStA/rsatNxIn5UB7bhI1uxEUOAHBFxz5B
cTaWZ/+45Ns/S4rWqcg+EgDGw54AWUmJfwITMxlLLHGmcgTK5lc9mmzg+3BjUTXZB2bKwHM2qHmw
1iUFYorpuQ3PPHWB/CroWzAV/xQaU8osPk7YHOprT+iShPg5TKeijnHu1OBZ4GAOXATRvnNZBRZ9
5YrU3svP92O0oHS9bEFhVw8T8okDdS8/7vrpH58jGX4Cm3tkbZaVcER5C2rS9uvmkRzGRaqv5DNU
zefXKM/6zHdC1ep4fpQLgeuziEcv+RszC5QA6mc0lPsVeulw3sIQkt0vEvi/HmKDmmJGNWSj9yhs
eSR/kNS9Vim4WllXvwYZkAiR8db6XKr2LdG1j+iCuzKn8jvkpWZK3OGI7TvANqTHf094N30NqFId
NBZeAzahm6ns01XERnBuZup4Pks35vAHLJA5UldK0VFQaiOxo/J48FEMWOkil2QOQ5z2xE/tNMEC
q2DAMISyHd24RBDFk7ajytMa6uDkqHLVs9Fi0edvmC6/kzxW0AsAPi713QdWhNGL4POis6n2+TZ9
PbQBKwBFSe6/huOoOxIk5cAMiynSnxbOdGpW0nLKpADC2DvTqVjMTEl3lWh6I2aJseHq105XTSVh
gcP3pdTsTr+Klm5jTJ3E5lQ/x+Tvucn6My6LuPYRPNbgj4L6446IpJnM/4YLBfzW+DcrwJPTxQhk
PW2qob6XnKJ7K0f99mkDO7Rb+Z9kornqRr1lmTOdvUiHI5M4/NAruXnJzRZWc3H13azKuUv+H7LB
YCan96BvnQQw1lS5qQa575EQlH3Wi5DZki+uU9vuRMU46n6zlZiUGK775VNxApgZhvZ0w4nDfYuI
Aq7GM1p2DtZhLSl+1vKbZVTUUSa2ZBofG+b/foFwVJrx4rJXRK4RSbg1RneNYFJTqGVE5/2/beHD
51P1MOtMGblj8te+GCmZD6p/zrRbj43Z90VHwS7iOQZCwANVAECHHG3zAub1b5QXV+NLA5dX4vGu
mmcKxzPXi2pt+v0bvI4+lHq6E1iQQZl74h/DSo5qAhIdUtx9TOmoYIUuaqgeNBBO1+81jFnz+p68
S0NWAg6RBxbu+2XNsPgjj5L5rQol82KLriZ71cRxovV3T4FwJsKUL3GFdUkXDtn+dQAd7c08syBC
avWxzi5mJwy0zQ5Ii+i+moTBQt68V453NQMcLAgVnzsh8TAHhMlfGaCR9hNE4ans2P+maCmbF+VF
d6tU5s0tpvbiOXSoBR1MSAKmmsS/kXoHA1Lc1Ula2/RTSpmGnZqSNxPEtFGLKZ1WhT6PVfSl4umL
eAZFXO5mqFLx8D0che8O282RARyGDrtQfIg6WYdJRkypcW41J5LRhdqMrhhNZsph/UkYU0k3+ioG
BaAUvuk7PAQgVxkjsNR1zJ4vwI+dd6KF2gTIlxqnll9iPdhwxcXpBfNo88mqww17kzcsgv/eBKPu
dXBd0uTn5NQ9w/jOvypRizX01sECKCLyy0/ANidpeGph3wiCwJGRh/zbYRb4xO4MKa/0RMyreP3C
8ma7k+WCPWv7JUxY9tNN4IGwJmwShvcowH0+o+reAemPRaiLHtGej3EmywrmqfwDY7zMxZswXnIU
VHc9YjfHxvZOtlE21fWmGV+XFyqQfcRDG8e31rSqDLPN5D/6mldj7pwnvnA7eFnBKUV0RhO+t0+T
7kSQ+5QKwVGKdYJj7loorOV3YD7F7EhMN/Bwp+rOInojlqdcc5wEezhKWxl+rqQYXCuDP5MTH5l1
I4htxoFS0xQnK+atpVzyxHk3/sPQNBx/6Kchbg1dIgLNGg7fgPsSt1T9jTOr+OKzSw8ZwurYlg/e
uKlPDodyrtjK5xPBmpHik2lvbu5MiKgl4UgQsiLE+lVgXu2C7nP1xvcJYxyTsAKq7sNCip+jY7a5
gML21FLswmwyRZblvE/gtMuMRjGm/gZpInIkke7PzHWfMqeYwJVZaqUdLmoZwDhGzvpBKt4D5JQa
mymw1kJFdGi//FGvCcYjrKSUpJBCGBCJ7JZwJb8KMPGbiyipGpVw6Z006v/yw9e70hd5claiqaOJ
ultmRE73JrocSRPqPrY/vy0KntQOhRCfHhyJJM8D0cPNqpm4Hb9xiDycZDgU22pZDydDxabqslFo
2x57KWdEPQHHDm13cOABMGCBhJvlYmsCahIXJdNUcRWG3zvl1iExfm73laSOwTJzOEpq612yJ8En
yP/tTJiEObgXYaHXUXVLkVhSVADinD2BrG07+mDR5BzkDzm4xBczy+J2SnJxl/rY6lgwOBuKRlkt
xRm2jekDkLLiMh87daS5Bl4hqpFxmd2sUDiaunam+VP1q3CMvxwRyLh2XKTCMVpR2OLA4ZME40Um
ab1LTCuBrKiEtA54V95YpPsQ+ddPV8IH3ob7dWRnPQqObklcaEK8LEoklz0S6X0AjhM1xFe62JkJ
03BG3A64+SpnbFR5TxhC4UDN0Q0unM83wdAkpwOCTKgq0WI8kXBv4Hr+f9/aI+x3EIH6UuhCfRpy
X9Yo2DZxGHHVq6r4L1O9RaxexDnsXJ13MEmDnk4So4O6U9W2AvRsqTNWREbQdw4upNjI1BrUcmCZ
ARY4gMn+cqQSOvF3yywhmBPLZsurIe1bYWwRgnAZ7FElSAA0K1BhxBXu7obAFoRw90ygWnXoU7E3
zyXetfhPxjHqjVVQMG04YZd1SPAH8U/cBz29YFCvcJRwtxYQ9EJoVxHE1MBBzqE4v/5yRR3OPZkG
bFeaDkthTykx/5R3uO+9jVRQTBdYYU6E/qm5fNrib5IShMjELbWKEnLYR2QyAh8ZH9AprRGQSgyj
1dxHmfa3Wv8nSOMBLF+Gu8WUSunz0FwjFrwxof+bq3xTMWzmpGwTYkfLCuiOEB5C8y2RzrIOrUBl
/RXkqWAC2qILjja3frnxJ7w47MMgehThfmkkzoo/iGPhZewqSGqDRgxwY4giEd2rsODOv1aTV3mN
pFFtQ0QtYS+iDxNIilGSffhFm4rYn6oVC55lcWlT2Q1Q+Br6tcWGNKY5k5ggi75poBPMhkFooXEG
DMPAr6ZQsivvnIP3CZ/WYigqMCJpk2/DzOfmbSLFED+9oX9+wumHIDrAAKISbudZsgZ4Ju/B8kSi
7cbNRNnn5sAjZ77Xu8PRCeMRhBNvqxlm1cWNFnrT1sUy3CNK2NXyieAzsMYCuGylzlw4toV4Sawo
d63H2zp3o+uOdlHiiERQZIDc1eVJWGwki4wxY004yaQjkfl3dm+P5xhEHg4C7wGVfbKf95nrJc9F
trmlm1Z+b16Y0I27gcHA012N3ImAtGB3sQThCm5a/kzOFC39N5qML9eMxpsnZ0nntav6iVIsDT8E
9ibR6UhKwrrReKp8LpcqSWQGT3ziLX9D4zVpmL9LPe3fMyevI46n18zruYPbiEM9zc/99zmWI3gw
qyut9D3VRPflfkyN8jMwAcqj4La2s1RkG8W4icu+N51RNecuwkEK/sWIu7Of6ZuyjM1l5mnUe2vR
qagAwjvQLoVg2Xb1VoKZNTkWOIGgat9PkUJ/5IhbNvNujOHnZ+u6ENYBt9Ojowkl7v107lgrbmas
kfo1Tc5bg++m1k0+x4zGiLpTuc1/c7KVfFOHtiWS4wY+rtDBmwzlce0tRVOW8wSrAhE95Fw7DZgD
pVBdxp4nHsgQqOTbDUiLuJaKK+FCSU8ENUFkTFmiXPBZo7q8AgV9TC6CglUYBJ48mgvHdq8C0BH0
ILNSnY+Xw5Uoz/rWn5DFbVFEsqXs/u6vHgd/Qr5WH0oqEPKDtuZ06tZgOOaKnIPgFu/a6gcqsHh2
SIzLPtuHhTBr+snQS/vHHG5MBYQadvAMvIqJXh4WmDxy//KuwoKWp9ptt9jbap7Raq8LK6c3ezR8
sADVOHjfw5UAjKNMDitKk4qHxZ5QjEGrFBnCesxtz/3DN7GIm/hwvhE8L18lSqPSaBfh8Pk+27Mg
4DbIjKnvC3GeWufSSF9aHk31M/Dd3DhhJ1bxpVtr7AZ0O9z4tfg2bh23V90b5/3/tmCRUwMUbqyM
Xxg/rXm16MnekgRmPOEgTpdu/HF44LEcKNgvFFmLaxJ0KTVqtz3b/9pxeRCo9wrIu0dG3XWiJjEl
0T4FcYLgl2aMO+9W1CXd4BNKaSBQLkaVxdaz4Ix5ilb48tiqK96jVJHNfEyY3+97gNkjpIhKJsV+
hcQWaL7srjBa4K3l4H3ZyvL6S4hjuaMnP/IQQcsZlyZmPju5X4TahTYkbeBMhQGXdTtO9WVGxJq0
WKCkX5bfS0UxX/5wv17448o3gtvdKaxCJBI9c4ejz8dh7hvOs1AX1hVTs+Zf+uW3fIjWgzYdNf4+
6f1u0QEGd2IFJgpF8923K5n2VvnsWpRw4eGLWwAeL+7ark1UF8xow0iXski7jbB3DH5PolvGG4W9
xNCWysS5nvc0ujXY96FNXZWRJ67iqehhzlRBXi9SmDH8d0shoUM37sK6GgE86WOHpy01pBhecVsf
wOtGYp/wvKqcuqqmlF6clUidOt5AuSJZ27KUA2J+ZMXEZBf1o159sNSDOIHLrB1UY8MOTiIAGxLA
Q6HyBcaIGxnhG3KA1UOS4J8e5iLbgPOYXJmPwsqaH2fmmGxCsWrxVQJhbVsbNOqu5mevmSHkhE0c
JhwdVihA+TgPLPKPT09dTlYNlkEcrlkHS8Y+Do1VokmrXWhboXUlnnpbVlS8eFNPdfHb0TCaSuSv
yKmdQsGo02h5eB8JW/cyxA837R4aifK/PHVDn29D+pfVpV0qLEPHgzdOeDmpqRiZycPj8lmey7vf
v8foEfeuVES2+Ip6zH7CX/qV0CD9XS0QXuhiKYjak1I6QA8+Y03tsuX44IahG62/1eS/JnBaWL0p
y8Zo1ytyCWPnPI0vQths2JxFmqv6yAjlnt7ghcwFRtgj4bF+VdLTBnvBY0veWLOou0r+qtXivvA6
i5eSOUNORJ25+zhUpRkB3fYfZWMq/1tieLEhEae06/AK/UiSU9UEzzEwvEWp8xEl62ITkBarPAc1
zmtRxVn9Gqca47FCGYJhyxT8J/8y6hNxIigjBOYutoLePTGzNT7JG+orYiTEEtFIgdmNin8TGmwA
7lbDGUVL3NzpJ0IopTOyVbAc0RFc42qOVptF1jlU9fnrXBcIw6jPBn7pwvvCV/R0f7U9hPeyWbCu
KS5NM+37nHlKwZdsspVCSAxF29D8LfKuialdXj0FnHJpyPI10Djf09A8vQvV9giiYZPbem0NXzRy
ZRo8aO5rSvhuaN+VS0q5WXUoPyphZzhnvvdUG66QrMVVtzqu0N7vwSJ0wPenBvMUzXmIx+ghapFI
nSYrl0wuehgukNE2Y01pqMoUSfyCY4hUb32ZnQvjgVASAzvDApyQWr2pbLqzgjp5KFa45WMBMY79
uoh0VjjAc9OY6TjHfCh8oqDFQMrNKHIsOjdDtdgxPPjmizl7RD47fLWTiLwAnrohRTzwSVtsMvNb
7lRQO+gaOZ85VLqN8Z2m/k3UBlFo3Ku6Zrkmck7xIjfQaKv/8umP0gB5rXch+GXGOk5jmjrTcjAm
c1W2KQtIu2az2cmQYVREJ0jKHmbhPq7rnKtafzHIiiFWcIhx3XGMuvWaYRpD7iTfWY7czJ19igac
tZEjNJUmiMBGP1sya6qwr+SADxKLQWwgZJwlzBUWXJWJ0xQufsR4lr5k8izehCIYvqRpSdG9EmVB
yMl+qNTzJMRwaz4QhTf0DUH89S/98blcG8js2x5P2+AgSaxHL7Be4TJK54+5fmote65SkCCE+fz6
oqGsgZxDfwRsfznE5SESABSWntdkw6ReljWdYsXakYbB/GBWikT79ivAXvv2deSB/xOokEHUqfTn
vx2wICLi9oqMye7B8+EBJCIKlZ7PnfKgLFQ96X30y6MUZKLBnDrSvIUAQ4/R4onLV6DTPY42gGAl
Jjn3jTO2PGs3PKmcblCW0Lxx6FhQwnEdqvk0YsJPntb8Y0w4+wydGhiIlP62iCFgrQUI/ZWrkfHt
zm98zGsJrTJgDoWj9HYwf0UMGgijqPpc8byOKzzZb0RE8reFlrvvvXXOkMhH9jjfrR+VYp/3jHXr
rQu+x3/An0ekdeX5/OUcIF14MWCS9NzVciYVli+2VHF7RkpWKxjI/HUSdCg7b3YbY1SJjrO8P6sk
adE75e6M6EVsRbdR3B6ZIUtFXqx1pbS11WbXXSvVri7Vy5qHTXZ0CWUauZvHRXSLq7aiqmLzfWTI
jnBJ+gdXQXyh8YXl0pNORrL/sMsYr7QRrRpONlW1L64+sT+KWeFAEgUPcIgTW1GwHisOWRLgsIQK
VUxJDgkg4pL7ZQKtwOgA/lqqLCfVOnLBl3aJK6R2j/Sj6GYJkd3bKnQ42qUua3Czu40Z38jAcJ7y
aN67rzBuuVURcKx2rxrDuo2vsMQI38a917UvCq8BeCzX6ro8Ql4Mq4MwVhkiSsYn1SXdSXrsp/Z0
5AJeF7O/sBD0SCOcrk3d+xE4QZO7AwuTZtXBa6nQTwpx5JCevU9Y8DY5DfwJa56hwdVVYPID3nRj
gxHj62hanua9EP7NcYt55mvAdAvXGP7Lm9OwSzJQ0xa2URMWx8SBu3sn3oNZEAwkKNlU8KzvyzaR
a6kJL4998/RlMzQse2J3Yxr6bq84kLpImugvt3pGLwZFcHJgHBMhmHynzA4hHQlJ8w6v6KzWHgLZ
e+FrV1U5YMnSvIXo7f50A/k1nXMoDL0jr/F3FwS1+rM7qRMS1w0PXrSYsIYkJj/ax+ctqZeotn50
3c/48G07nfUZtHLuzHuCspt9PjSzT51GAVWkhpvFCkJJni9t/iXGOZHjaaNDSPHMaXpDMrUrYIqJ
/kfMev2xaPDqLgX4JPw/iNpJzOHeovTIP0+jbiKDeTbe4d/F2GFdiu1q3kaCJY7a75z2IM7kvZ9D
b/uwKHh+omw00DQT1pUY6TUxOEmKI1Kyy3EemaBF7uGrUEGcjhL9sU/yeVwNKKfj+xOxnulGm9mF
LasX0tdiym2O3WTtwIEDkfXyJGmhzoxoLo0LRnSdXNAWXybJluEiPC0P8wM3Gh21XwRLZ3+jfNLB
cWiEQZCohjkXYsadZO2/Us+stwOivnSJAFomAQuxOhYSk0eCBoo/1/5XaXfcExUJtPVWTlDsZPlG
gLZgpcQcFMYdWM0ZkvGt6PDH4KQxoTOSRbxkApTUGJWu//vLqt1zxG2u/nx6t853fiPc2+8zKit8
ZhcEAW6iv2QXoxSLRiphuVtm7PKXH1m8ZBhgi11yH2/ZTYU3944FXp3Kr8vAs1u41nYRmJ1C7sMN
aYKC4DuPD7HKNCf1K8egZNJIHBNkitnFPG/kY/UXS7K+xD6c7i/aNx1czcpqbeIk2A3Au0s5TcH5
2gtU46uSwS5zRXks5uYaTGLAymClT8kaJ3SIgdBvgGLjXNcW8VNFRSCFzxKSSmvNRjvSPc+0y7I9
JaRODlO6oSV31W+NyG7E2TG7xWO5MPfAP+adiM1pbqB/hRPsyIkXbH+VlPCWGt+94we4j0hbjF96
vBNBIw8H9IgWnAqRzFMc/3d0GvPvuEjOa4dmgDRVbX9OVldrkQreAV5GLwK+EAc1Q2lLar+zekIS
CQQcRSO0S7ZrqFAh9/xthAx0E5DInLeb3hNUDpCL94WjZlit7zjU5GqEG41k5vz8JKAd5JSb+ycC
muZQDyJvc2k+73JEUA/jv2h3HSvdZZTVJg4sgSeL/MemB3E8pcalhb3zHfYqmK/GEJgSym5Bx30k
356R+AW6xX2i3IpKsrqVBI96dPl4N4lIJfMikYQOEqm4B9U8Fi6c8g4VfCVQdZXQKDBawAuhLuj8
+4QDOtDVU4xU9Dj9fHZGMVrPnRTS2+9vRa+Ya/A4lIdcZiAtrm3GK51ruVvW1tAPsNPNTmshB4Mm
4Ht/fWReuzjCF1GbVROjWdrFE03i6YMwXWsaFBBPPcGOM7+bh1Cf7SoCZ1cNmRfWIFSkJVg7jVOD
oV1qKVvHFPFZ92kVuG70RtukMoQjSdG8kTdpYBdynD/Sa44ugSJaRgOcSOuUBgHGl1rVQsPS4ieU
te+WGOucoibVvLemn8vh2xW9Efln4EVIAmG5M93TAJqSXy3jyTJcqftXBnHscD/PLrkvBooTQv19
nvQ5K6pSTIntpPhn79gsKjil3wp4oa8lgT92VATLWcAktvFqzTVQoIpnNE0SBXtl2TaOa0NoYLWt
wFhJ4fygA873APXTQ+V+2BdcdW/vT73a1M0HhaGDk7EtGy1W4uv72TfzhCb9NTtKplazCxgxVfvO
b6HO1QtfxnmnJBdW/2sRYlkyiS8GH00934qMRbxiZjpSeMZiEfZoFmTSlWOO2zjrs2Hy8Hpnx6H9
uPUeznz5eNXe0R3naWWKNeJvJGcQquDkufhvmuDGiDZfnZsi2FEgN6RN1JSuu4rdwcsVSjANp4lH
yQUEwCHosQNcgDnIjQxJOMEp+ZKNju42IxZ3rbwXP8aRadoR3+ZGzaxPUnPiMNRxK9FQT+/PBvxn
X9Lws+RBd53KoadUyQI1of3tlg3PFOPh6EYmVnWwv0qsHRnSVOD5X+XshOfzSPk4Wzqa9oSyyWbn
0YmpO4G/vwTnkk3/LLmcjkSr7fALF54XBIZPuFXq/UcsjsJKZgNEFPn1ZMtS7AFwdQVIWZ2+pbl5
jXrOl+n2kLwCxBUzf+6emqjSQu1ckfPgE4tK1wexUyi7ytV+16wuFqy7rpMLvfHqff4MEk0CWaQW
HAjkX9sGxYwPp2LkGrt+xcwmr2bPMWguTuEYwPBnkVY+MThOF8XcZqgC5lrykLmBv5U2mI8FA3YF
8ACC5nEfZdTKGO6Pbc4Q2UpYy2ylNsDdLYoGKRGC/ilZ+2MaUSt4YvXbchP6I5XM3QwiVxcaCIdj
dzLkQTsbk64Y05aNyT9Vl8O6t52f9r4/kcnPNDpxpmWaC3iRsorc8oPZO4SkrkQesTmZzZ/ssLS4
d+NSNNmsX4dT90VqWyuQ4BWhxIHwPONbUv0vdsVFbFSU5u8Gn060o9vQ8CyJ60liQIA7T7BxdBnH
Xvm5+lFY6PkkUE8P9Wf7FiLvBqrF8DADJWp+QHGSIJsnujHcRUgwMBc8smYtleoxNYIgA7slbby1
0xoTsWSagn5wHQqtWH76gSVUk6ZhjVrbkJPe7GXtcjibBuqONevuEPiNVv9n37SNtcMbk2zGoYSx
0FJkXP2zoouispcQIyLlybEdmytVXWBmrDMUTnBQQHQCkTYrTVFUffQx6U0j/g8+I2AbeRfixztQ
utXaGtsQWgkWYjoL3HomjNgfMrp+YTXSJXb/IHIwsUvsWXrJGHaaL6BJ32odOhtkxSMuGm2lqeQ2
R3luwBU9hU0IhUbECcdr3IipNy8l1oXOuO2Q3bUmyBrpJc8vEWmHnEJvhUG2wGJ20EzC/wpiX53V
mLwI8AgGyBQEiNhExJa66u0vqm7zT7ZSdK1ar0O2QjQ1wf4vynvplxHJJ34rmBG5NGg0T3IUOEQ6
gime/wL/E8rCcD4AbK5Zd6JiF6UsVxt0m7l6ZtCXGtiRh7Ccg/JcqRZ7e+pUGEIpA4DzEZ9bWqyT
SUYRGG1EtGSYiQ9ukErWyD7dbSEhRs/1EJnIVnPjPSlkosmLWfffv/012P6OjMY0f6tvICb1NsgC
+VPh4VPzPLtTVZWDE5ti6t9B0ltbbwvjmFGPTP+Rh2n8Xc4gs/xyckA4HBYYL7tBp/qFG694kAk9
tImAhqz4beZnbMtwcuZCIg7DJjAs5AxhXx0L6vOFEiwHHeHjGitP1sLBYrCxM3Dr8OpA7CQffZ/Z
hcQqjeRYg32ZInvwjaFMLb3ZXpj086GSs040iqRNmk77fbgg4NoD0UNc2Y/jjfnUv54Lr7zpyfYJ
DU5gos+P7UjxGNk8GU3wettpcZLn6Jssh/JKcsbIkcNMPiGzwml+QslOqdIQhsIc9/DbXFGQl3aa
ZZQ6QoScVxv0xBvlVuY4oRCDzp6QctaEcZ74YjQW2UAXuO+WhVkyHblg6EoQmm2H+4Q366GZPH6V
LgB7Dq//3UTpZ9S3jNTUciXZr05FL6H7uzqwsnW6zr9Uu+w2MYkVi4gsFvGCvSyStaQO5PwsNgA7
mMKrYltB0R9F2kZoTwiuIKnX1vena18Lm5SPCvXZt+diMugvV3hTg0wJKVqe0SNoFv972OdjgMFg
P1AHsnlx/oRWKBPN3AztEEGbsVhE15ZWkqX3SdzsKqZhxNAuIml87XBK0EOM7gGFxFzTloFq4a0k
etPhUE15VidMIOYBS7PxHzG98Ynvz8F7TET3bEw5pnXM4ow5UyX3A0UFnQJeVUsqTyoU8HxZ0Oc5
C50RhFM+4cIYTb1HzeK2jA5ZElAKaPUuI7AVICSukDPuk2cCqQyZAxLomQxD8b7ZDR3rFXMMZDQV
879ceNzxpxab4nFMehBAkmTolcHQXSStSsy+8RAIRgMhynZ+cqHFsu2g6jcfrFlnZOtJ3HtC+YxK
+skhhEJdUWvAvUypcAYb2QS/NlDRhdvCaH4elSUTzoU+jndLg4aGA6O6hAhsE3bjjGaj0x57yFUL
wewRXqMOrpellb06NjUqmE1pEIpg0Fm3CnXvIXfQRYWWrh1CfC8krrqo/q/+hh0E2G5sUbWj180v
QzzdxjsXI9O+HvBFwyvb82vjf6QkuZ6GL5ibvFGI+81cFrVJ83X1AZXizxaMD9oyfuBirblTig/A
hFf+nT2Q7ZgLXGl1CI5QcnIOuRTCNoSuPTyAZ2OjveIlmSW7FFhgWasMDmgMtU/lL4lE7CbGvh0l
PxuegiArQDYIIUIn4qJFBEqp2KmvIe2j1ajXfnY9FiTPA8EIL1jNm/f+Ye6+vpsPzbanPRSCTd0q
jGv9KZuOMHbT4ngkivBGiSRrRUcMYigbLJ0oGFshgJWMQ6qcEThfY97HGksW4mVroHgSrKYZthXX
hPY7sLe5zc29NT/kHZ6i9gauT3kONCzBoxl5p5H2wq9KT5Xi7H2yF+wdH/Erc7CqEgcT2KFjDyNa
TuvZeYPQ1xRpdszSSGaP6SZ1O+QvDytIMtpmLsGVJ46OwooyZDZMwooTb14WAQWX5jDlwm6yllfA
misE8PhCwUvFXVtxsO/He7Eu8+EgS1w6CktzFuGa2zfE4broL+rq6Pabj1k0csdTNLemSvxd8Ak7
VNyWu7vFWCynNTDGrtorLQ1EL2EzR7Y1IRTyaTA78afJvefTzCBNrwVrZyvWM4cNYWi66ZdRTW7f
wNr4YZSR6NMVDDMis2OQQ7RKiLYaXo6uMtfE5yT83c9u2f8UL3U9DOXabZXsNFKa/YQoYEfg7ECL
JeRXLbmkzXRV42poCv7djiGwUDcsSJq8Oz4ZiPps7+11kAxZ3zMgbDO+16lp6q7pGcwg8X+Fdd4+
qlh8Zw4S9Ry95W3W4MGjBfWLoD9kjRFymcwG72x6jSWer2jr86AfCXfK6tiXBEUazVlh51W3aCgw
4wTU6lNrFEKriTIvHyq0IhwWKrbR/oNCYRSUiFL8L4C07zVYX5W66w1+ocSUQY3Zi1ivMcqJD8sm
pMZ+xf/7cBb1mIHLu5X2GSapChItOplVFnl3BJSp668NoiRBWky2LznDWqNCEnb+gKsEp98Z0/pe
Y8xlR+LvcJIJ/DC9GtcrwXEM3K87CQHzG+Jsl61T0xLvhRhBFlUoVnKHe/U2FCHulv87yvSs2aqX
LbBbfyINK2WLz6VjFHASd11fVtjcYYBIzeNlVULToLThJMC21hE40P0z9dar/mlWxXoT3TMP15JP
4U3RvhuHeAKwOd/NeUcFn/Lzvr0l70Ff2f8aA2+KbrE/waWCAd8cLbenUdcP5g2Yzr/maY3LxFtJ
8/gFyix3IPt9g4m/+pWnGtZy9n0iKtDCXwlN+V/cuiQbyw2yGTc5aJ6mx1FaH8KYU2Y6LrMqRY8m
4P6fXOID1irFm5bmZKLtDn7jev5+IRxD1CDxbZo0ane1LErQT/xF3EUiPp5r5z48NzexBa9qapf/
9OjsaqHbcyuER09LB/ATGRuIzvPZ7lLko3I8uMUxVPUeyXtaFReimUl8If8NRu7AmYaMaJc3QONg
YZJQfGGvlTHhVvStT7OBp0DlFYxQZ81hxBFsthrSTEEn0bSSQMicr0LdFOdAJhVTZvw+3H01Pee0
8TzUC1nXmep8TbJ7hQaY6lxfW2CTgDKPWtGmSwkqqFnObhPhNTPlJ1/+q0i8I2rkIfH//azChoDN
ezj6vDMdrSAFXg2R+zEb2Qu6DSAFZyyLzaA3lREoiNxKD68Sv1oSW337TYINfqSphY9Co90nlmBj
Iuh2Zq/unzNqKsvuPx2wD7JUg0Mhke8f2KxRley+/jSJewxUo0sVczPqReytFgPZzyY7kQQJQySt
CcQJ+HwVmDyUB+Ul49lBMiW/g+6rC3VYjO0COFPNindQ4Rhh0tcO+WBhpMf82oIyRGUlrSjlhrgf
vd+yc0EPUBRj9y6dZw10gMwRgNM/KqFo9/p+rU34DsTWZDP+IKAW+4rp7CM+9iqF/4ryKgx87DlR
FT/8fMMvs6PX/XzNhV7wV3V1U0kzf5OBejQtIqcN2P4IO9KB5uyyBXGI2lX1txiJVLOHLzxDlukX
FfF+ERsXlMK0Z8OqUFEFcAyFLFxZK8/nX9THQ3mQfb0LoktOLfBSKlkiFJgLQzGjZtSsEJh0yle6
9kcnDXYc3S/itDXWMZbPvkoHW7CaUyME5YpMA9KXAXoSWP9JfLsMCYVzqwkHYPSr881w6hpuqTfQ
dydx/dlLoafHsJ/Z6RNoHCcKV36gRI4B4WkM9UtFmMqa7y5KE9/UV7FHoj7M0woG4zjYBXYnjWrw
3MgI1GyVDfI7wCPImraVj7QdEWuYxHOYLgJTPK/k7i77LQRAl0ZKyuLIEQjcK+4eKTg3qip/If6Z
25LNk/SundY6Di61j1Pi6rmHdYpExvgLFIxlDOGrkP4lQJmi8sTJzs6lnkgjrCe71lvnu5My5v9v
4A0I5LQ1qpEzHfwGdD7VQNIxls+AxRFVO3PyW738+4HyFAkdgekRifk+7205mUNy03rF43bOmQkV
GIElZCS2qecWU+EW2Uhi+6xwoNqeqELPx8WS+SPzjBpwX6pgBPfzeoboS8JVQ0pVZ97Cub1FOclZ
v9OtKxjPNPHWDK+RJtMFtnSDXyvCzPhbUe0XAWBpZKB2Q5+epi3b2hLXW2TMaMJEp3yx+G/WsxdU
yB+wqGHeCi5Og/+hNAleJORIvUZMtJw4E45bFFJLmJrCoJ4TC/HBvhwAGKm3RZorhVXTAVaCZVVt
nZqIlMTQ0JV/fJz0P2gASxUAW2w0kho46eJkPRRQR7QLgv6MPlbjcOv3jo0jXmZabduANaIHCmXV
9OtXUN9Y/8m4coiVym4zRDe0oeiOlQgBrdslkrv4F8UpRklcliDo3RHYbY25MHbHI/sLnyOlIJ/V
dtz8QacWUqHHyBzZGLAdhyX5fFpGykLIVg8WP39RUqlEVpoGJgFY3+8b/a23TDZLR82rb2y2sH9w
lmwHoeLhjolLBuYQJq1mjvCtAZVYsoDYQ8hvVnYrC+vX3KS3KRzme3hjMzQBm0rWerCrNR49JThx
sl4wQlVWgkhu1/Uh9/8MMDTjus0m5kspXGkH4y16jxin7fHT4NMtmoGEQ2WP4HE7Th85fVGmQ25/
2TsaC5tgLeajUwywCb7ptHfbSWJ51gyi3UnaN8H0RfyJ6RxdDLxe20dC0aT6y+RSDASpmj30zGH1
fPiHLon03/Eov9hxWi7LB9+jurHKTShYQUdGCdpgRbF2eF3ejPKlEjmLE7c4I7tpbqOMOfAXAerk
kPAWHKJ6NTOO65v/xwK1Lu+q06+lq/bBsEgwBIyTC5/OL51FE8VqY58K5syJTkbRPt+bW2Yl6Flp
Rv+9ILBoRKFTZOhUhvRxX9qhA3wZ50EcS42R/pcmxEmySBDt84Asjyn392kcouUShKMEfQV9N7sf
3LDe5Hrxa/FfN7Vyx+HTEOhPcnf3/7ajcGFKcY0k4x7j1WL8DUkg1TDZWYwpwhK1TtOEOc4fxi9t
jplXx396mH0esHJL5RoKIwgMpPKcoOwvoUXMBxfHNyY3aD8m8h/TRSBqgbWDcZyiI+2rqsFQhGjn
Tv/f72FIpfDn35sVFH1DfM87UJeLkHWxrv9C2fMq6esy77prU+gFNm6gVbHcsGisvCtd+utlIw5X
MU5wAJ+8xcMX++qMfWjFl6W/sBDl05PPbTnmAkQsfSeK3nRljtr+PL1jbCczppwEtIxw9e6AZKy0
2z57WR3xjl3fhLAqrjpLlIen/VTC3HvWUJ7j8Y5ERa/IFJ69zi7WSmF147wMa4CHfFimI2k3afCw
GyI8m82kP/sWOsxVw/uymZiKfuuye9t34HoUMi6qdG3d4KHq/kOmHDQM/pwm6WIeda3l0niewbkL
vRdG3m7Iq430MO5wWvAOLugGI9G2wBEK3xOBf5zxc6Mz9Uy1BykbpVd4/BiRlux5XOjFjWHl9GAP
dAmm5h5rpaXpcKJjf4kJAgZr2LO80hTcZQ1JRyLQmnj2B5H+/G5LPZ0pYJu9eWW2nphBQ8Y46so3
YuGHD6fi5SKVG50rgosMnRuBxlcMtdrGIzCcUSX1UBvrRYJYtf0CDz9eQiGlGuR3BVEH5V5R7i7w
l9Um59dDD+/jO+U0ozJR5rMUVqu6rQ/AMwIFGLDgKJJolhhv8GRgMz0Ffe3MsxYBzI0eD0/2HXCL
RWp+HtUpzCDeNyytvguAzAfcRBMHgnlWo2x8vo0+bmlmT7NIcJjdYEnk4imBen8j/X0/UOv7YEqC
tCgORD90UhfiStRgkDlvJmMu9FBHInSUvTn/M1dIsMT1pNnsUg4xj7kE4LCOI9K2DrCzJz/EE5dS
yL6DOh60+XpcozSivpWfsUwPti12XXmDl13Jw97tFVWWCGjPwq2pOeGlfrjpc3lnGYcw7c6fN5IH
hRcE4IBmAdRBPxDi9Dd5kWjvy7NFZ9fFYD8O/G9PXhG/NMtDFn3YrimiBartOq7OaXk7r0iyXvKT
73+cKVVVVDLtqFu9hynRIcbbinTHA+tzKtQqXtkf+UX+2B5e2zQM+CZYdLMn+gkzXddHnrLhXkUe
UVeCjtY6qTYjBfyuWmJJ1Zx1xrB/Bu9lzbDMF7sn7RGRm64tDIvkH21WfzPhqzyDGz2T8gK/CHrD
IWjzDsjDQ9WSEa2zscCOzXgy0YE8+OlHrAisys8+rPXBonKlPif/nGDLk3s3seVCEL6l0xtgMPgp
KpsgLc28y78jAO66AxCCAC+AzAYB9q+5OMsYIVeeUuTkgFcwCfV5ACzr15/IlI5v2umin4HIfLST
6RtAg28C0NK0W/8tQsgF9it+Byu3UiMOmXUyVM8Hyb/6LvCcMrAvzJBdtG5m67U2bm8624w5IaWc
qZ5XDOadj6W5Q3XZKpuqqox6JY5YeDL4yZU2OXLv2ed7UFak3aUVVfYy4TTL3KiB5JvaT20Lam+O
45FKAJQN5LfvwUvUnVHg7UaTCrMMRZWP/gLgM4PUrWappnDz4ht73pToPi3CllHtEsb0UqRIygOj
dQdvO2Yd2PXQt4B49FuhxG5kt+vnu63GI46YlMpKCahBjvM6R1OK9+PRh471tO4kv10bi5aP1QQT
C7b1x8TD6fWuOxo5BGzbopRJFK4OLuBYXP956wkFX8bzoK1moZqAJZEbPAo272mY15Rl+KUHnGnl
3W+JzXpRYvSI5vasCI4rF6/i2makcd8iBiPZrZoOWTAA0hQRDpvX/sUVd3/5uJhGue2YYXHsTEnI
XJIlzpObaT5+lyTlZWlEKgSNu8mOuAuTeLj6blCTPlJ99t1ZuKivu3USbq62kxZ6y6KGszNlvbI7
Iy3qk7BoO2n3s0j5G27uRt/SNiv5CNumhclIBk0DUcSt5vQegNuO0FLOP3I0Qfx6YjcmhMQXlvzz
Rkh6syYX/766nwEgmJ/Wd2CmPgk6EZu7P2ylNgGkzIEWw36doYkTyNhm8cM4qfpyPutTmSYYnj1+
PVHHyj0xfY0f6Sdmg5/sVkm9p0ReKYqYGeBQcm+epQ05PMIv9MDeC6Ez4GFv0JmKnUJrzG2fzRzm
4dT+xZ6koML76Otm/maDecFEkb/lh24ZoD8sTO3D+wWx35yQCck/nFM05hP1SPp1fz8XLnEiRW6L
uq+LUDfM7CP7DS8pb9Jjp/E9VyfUdAzyLTzWnjoPo/7/AJErUjX1nyMIKwC5J6TxmcxMiug5WgLd
LYYW5dGFNw4ar7fJ0FdRcWrmMJqo56B69kmq323eiS5qU7wnWQJ0ZTWiorMKIOPu+lHO6FOKHxfe
c2DEm+FUCx716c+effzx0M3WqfJSQjlupd0GfntQw16TJD9ZOunKBl4sbS8Vs34L/8qRMS1/R3t9
VS9yojaQEPG3YXw9iGIGh/V0wUwEKtFW0Cu6KiokLA6NWTwxwzqPZL1oql1eg3gUBwLhqCvKw3up
Cz8+78u6YLuH3kx4B8j0g7UehEzGS4HFd61Xgw2BEO9/EI0tQ5iBv0NHEE97O8YakllP0G3Ii+os
1QkqZwKAQpv7heE1QjIoPbuQTTv/fex8T6yqzYaLq8wlcfe/9n6Oerz9Ht0bBiPptWzYisRfrZqr
ipeu018yJ2a15Dt7JRz9rjwH9hejzGP3No84MqTWsAQEKJZ0Z1jKjsnUeWrosPBAraQYZVTxvNqp
tFoQYVx8YCo1lzEESPkjuenOC3/tBWu9riBlSb7HyK7mg/su1BrBfHht0e9I2jio3ysN2m+W+MZs
g/mlM1bik7RY4gZV0/fX9EVi2fwRAZ7oERJzCNKBXEhSbVSfOBLEJbOkms/f37mkdU8AZXaLl9VQ
C3rJ5NJn+T0rjIB145w6ALci3XHg+l4+Vt6b5/bF12uFC1JCem9gjNp2YPBF5/pUMqOTy9vlRVlI
TguNrDWSeadX0K2+aB6J1EIOjhBSN0oE9bUWilczeDSVr/VZld5VphspTtZ9+37cfgSWAHURCCtv
Xw+roUQtdQF5Jtgylko3Dd5H0SKoa9K2EJOOaEMfo89yFN8B8Sm+pR2+JrEzHE0c3VpGOQSN6G5E
btlCcA1/fD8UXNyAA16BiQB+LekTQFk6YVhKS6gnPNRYQSnQmV8Wpa5BwYuCN0E5OxsbfEa6NteZ
qX2V7oAoLYqX7PC+GISmVpYA88iau/9tXzwUdgVD2y+vrcgFAO+OohAmShlzBDjznHskgonJwx20
tueRTpqCN4mJImuCkkjDSe387UOHYxCULUz6MUMSjt/d3SLiJHvVM3D4uHk2Rbs+SQ/v6DCR/oJ0
frytT26b9sw96Mnd1rgf7G5aXyZmx5IRB/DguExPtC8fQUi9p5DtaRZ9fxbYOZ/GTMfgPdt+Wuk3
n07vGBnkz9DXKWsyySLHnsJ29rjNnK4UxXDhy1+SxXmdKFAT18ZojAZjeFP98FT/v3WNjBY11+xl
Fovxo04Qsbq3KqD+7JgBPbnsSlMoCwrGjBPVJaLe26E4w8aeQl7MxQG5HqmuDDrInZSPtuqZTZGW
ysvsRveDGdsIE8+ez4+QbdsyBkUFAAUzGm5ZbEeFg2JMHDX4S+P95WikmWZzZ20iRQEotgJ5qPVM
YpsKgdyR5mvXokxyp3eIgADNRCyWUpSfwjxkkV79ujF0RABN2m3RU2DzNBxyLKO7qnrTqdl5Uijp
b2MzTEiosFHCWI00p8Ux8kDF3MoLN+cH47pI8LxkIe5PKOfwMJf0bfUXbwv5jAkRI/VVarK/6tIQ
snJro7lnG6AzXm3zZzxiP3EuqK8O0zJaWgqlSpvrtBw+1f/A5qgULRbGyenrD8vDfHphLEsu1/+4
jO9KshW4RnMlm/p5YCFappQnB5Zl5V7SzqDOlwBL9idyx1aCuCz3e9VTswTuiA340n6U3aFaUCkH
hooY/+2/IivMclcqyNJ2hptW8YbZgYRflgayQBZf17o3bvPGKuMHCZZYuPZ9VnerDZX/3X/w6jFW
C+POpNy2umabdqp1nEsBiTtF31v43WIl9lAKo5IwrF2PIWcPkX/TQFQx4N8EHnkCym4uIK3PAP0j
PMOFy0PGRETH1W+wkITUoVe7M065Md4/AmjPl2DFwwzmGk8f2Kw5zIrCMMdsb5Z1/Dwue1KReImf
dk7RLvOJOIIROWB5jfLG9bkhICXr5Xy5ztwPGm0UMez4ycfcbaiBzqWTwbgcD1K519+xby4ZmWia
C++nTNIrSfU8MX9pzA59Fqmf74I1UYwf1bCfuwPEGVJl/zl7G8zlaEtu2welogtr85KNhPOYtaaH
SpnpYfSPNV/6UUTIXEOGiQIDV4mqCa0PdrBiOmXZBaUXQ+VQuOGrPOnNo2vIuyOpBMZPI0aVoyj4
/uTedgNPNY0sbQuEjWIO/M+N0LS8E0lFGBiqfT9GOnAnSO3/ojQhuouQIm/dmxB7FRxZHY1R4ca6
MQJk8QeHw5KTVha5RFJHBMGByB/PHaPVVJS8Rvc/+LAlcgfNxNGfWYiLmuaPebiBYeVeAroW2kxi
+LPXijNhHgKqsX8zoAQ+269MN4xXH+eE0bIdiEyuBRwgxb0yZtKyHrc+9FthKDggLoUE55klt0ho
TkNRIuwrIXP4qKGlLQ+hFYyFJ/Q4PfvviaRrzKbRubOVEVDKW1qNltbscueiwRBVO+rYQ0tFYOJY
5yEbcbbFJvlYIjc70IH6PqQbVaNtu2E5dOjiWAivDlB9TjScAmX3XCtwseCIxREeou1RnyW94w0S
RonhB5LdYsSjv3KyPH76vTihN0aepBwsDJ9DNzURaVNNyX83JdV5qLSccuGKIV2SZjQUJDIXk8Ew
Cd82cZ09PVy7ghOIg2Ybrt5vc8QtqV/Wro60Xm8XVSS7Tk6xv98N/dcXu9CgI+QIRR6lN0mhOXPG
Dt+znQ7oRxRFzPWCM0+VfLXJfnn/iB+1f9eGq8gqEQNv6D9WOWUnLt0yb5tJwDzO4ChQl4rMGSsg
5amEKf0BpCT6FcTdjGCofGkO2AXVYoOaRKrsNLBBNacS7Dtd+LVz7EXxlh/VnOovq7swkE2rZEi3
U4AwlgBeonmTOe417ErKf5VyOpRtSCxoGgph+3+aDYfJ/sKZxgZre54VKgWs26hF2Ex/vTYcKrRR
QawMYiyOCH0BZBEhNxZH7WAjjYCIHF74CtxNAFwYwppnVAGj1FpfhE8s4z8aeM2MaHQlcJhm13mH
EafnpwjoFd9W2WDwm1wz3yeEBFQxoLGWpnMkeoC5Kz/7DMEQEXeBS1OkmjLhgDn1Q3Rb7J7Olhpj
mb57xOHXi3NRTyIoTnrZG3P8zP0wZ2K1EY6R51WALu4hh3w+Udk19pI3z2h8L6bNtWn58FnBG3mN
DLm3JVM15I0pR4tHtX44GaJagt0ngq2blHFmgoeuCnDZ09dgwsqfVezyZ297B/X+/61LqdzalE4g
PJK0TOkCXHPQaQ8LfOIdTk5oxQ1Q7obV/58yXK9XG9re/r3QY71xVKA25PwVcoXHhQrOCEc9mbqy
5C5K92BgZ7kg9uH8k47EbqXnbno4UIqMqHiNLwoEkHKj4m7HgCs5NyKo/s11gimJ5VGQxLy9rSMb
ChJa4x7fcgS2S4bMFVSQLWaeRQaDrMhLdDgA8/CpBhRuMN6NE8PYCnf2NY+NIpNfDlpokQ6IiQjA
mT+Udyhhz8aTppoTyf6uTEnTaQcTgXA2rOi1ePiSbssezuO1JIC0W29NRnI57fKC1ySPfU64lPnA
FRZ9td6NIqSjjsBi1wRuenwyeAncpza3c9y70xZG2PRjKpl6t78th0Npt+Lv+XM1o63ANORzyAlS
1v4HN+3bb0SozpkMzmRpyg7TA/6QvQ6KbRmi2ePpdHLb/hfa64yCy2Wrs+RpBOKTrDJw5+lyyrRl
ypJzkV3rkx2OIXq9juSH+64a5OnMW4SxbvSgkSz+3EecwUoFUeVbIKlzYlMBB1Ae1yEWEAJ0cBd/
3GT35jzlJGwFZ9sfiOkKinsprYwvUNh9fqVus6bF0s6KWgOFZbBQJc6NxXMtBlEHWIwFvlN6avzj
MFIDsqOBC2ye5p3ODdh4mN7jzOpc4yuWLCGawLq+mcdL+3QikwQZe5tMp6yhYQ+D36R5xkGh3aEw
WFUMLHGkC1RKR46KU8nqjHMxSgTZqyq/YrAJtF5ZxCsNHUJAoD3F3tXYwLJ8OrfQaGpsaqYBp0Yq
TDnZ+vV4zegDaK9dkzORCtl/v5dLn+PPu+eTB075RjvpRaiLkTL1COLWzl3iJ5Rk4YHOfUh6VXuQ
khLjkRQurqZzwbvrI/KJl0GjBRXAnxwQBkhKt6K/Y2SI08ujbzp7RBA919eKDjViDudWDEnqaWvu
HNQXchnLXbDK6q1WaTweRrQwXtvngCjaqHgyfLTkrGHBug87nUopYdINufZioAHeleyx6GLIaDll
tv052tTonYHaYsccgCijkRNSgBGBph0TajCCvp0nfmX9v1mTOF/v44gv3tHEhg4EMurM3Yj4O7vK
fRmVt0ekAqyZR8yGOt0rZI600Y8tSKEL/APRmw8t+BRHzYzCf6eUMUJl8fYKBNt4vEbyKaZRk79U
lCxJcqKIWGydXg6kYjkNGjvwXxxn1Z0ZvuevYL/nblP0ZzL6pBLuFFx2+bQD86sVLLT5wmafH2GT
eMij3xaeDkBDtQ+Er4wDVi24OzsS7YHFR3FReVMYHYPB5fB4j777wGiKzgCLxshGY5551dWYMBz0
7q6AcWnXJ4c467cre79uKK/91yeeUS4yd8hYaGb6xjhYxnjnBP7BF4CXg6zPkXpRj4Z0TJ9P4nvm
RGGF7K+khk7P66HkBEobWgfLKvg5wCDWBredmY4u1GrNAZ+MPh7t3cI4i8LOuWXEwTwxK4S7UV9w
axT1tOrZ+0Nx3XikvSrb/g5Rdz2zTCre72jIRbdiRp7K6NJOQzXkosirsfd8djGszA7+5j2kMRyh
6ZuGCtULmUFpvJ9HbaBp3NmXVkoztVznTzvAUf1yMtXOULLRNWV1HNjIXTdAAnro/wkUzFBCdHQB
+SNsDpOFj3oemicTTl/vhpgxabLD/InOATHn/s1W7LfvK4Ja6Xpz2BydZAQ/YIKM2doiNMYYerWw
/QgnaX33GAPC6QXbmexsxUH7jLq8DhyuiAHE265xRI6CYedtt2B3DiC6hwPEKAEaPYqFXPRkzz3z
fkDqaBMDxvhZoE6MdNgEjASISNE4EvV/q/DydCTlmAec81k8BtiF3ZsmgvgUNc/Wwu6SR1Z1KFsB
VO3GvbQuPxtpw4Mpk9/IJHkgr/tQq9f5c2FbIFImfuLTHqDM0Kfw+W7DAc782eynGhRBb/ejkHM8
Ws+r6Bn2g4NzI8rLFYmD8gmBZZ42tECK+Q1JMKKw69HhV+jj7ev6joAKwKK9ca8qPzE+hSwmdz6I
9qP3u5PvPFjEdtf6DGMwkEfUQjfEQZqm38203U4y5kRv4rO+Wc9naEDLuOFlTtl1KSFZxQQXqUV8
qq8RQNnfchiTLGCYLdYovzMe8nTvqTYQU4i8sLUTbz26IxEwOj5HeEH/eSRHUooSwWIWo2DNDqzr
dia6KiKUfAgO0pPfWJ1cg8uuMf0awjGYA3/ohLOzMLHr171eqvQhffr4XFOOAxpdsfmSr9AV9uit
DsXDK4lmCk/hXOfSeDtQnVoMFpEIgW+6tbhHdvp5SyCHnlKRg+Z1qjvGFMYTHrPiJmsIdkCzbTtD
FlVCaViTApmQlm55Hgm/mfTD+yrT7AIDiAY5mcZv5MykAI3XtBcfhKB+0MYtk5jM483XvXxb95Jl
u321EdkcQjYB7tqSXnQRq3r9eq9x5To6+dSI70ANXYdcRUnz5KtQyyBQi2XW+qXe8fh7R0Kr7JqC
RMNkYi0jUZdOvPKGF6mLESvD+W0poPIfWiJOe+MT0BF8ntv8sMMwuLcRknryWCnZiNAmsJtcetX6
LHf8P2KJvkTH68L2YJuCEByz73Ez6OcSS7m8J4/6nrVaDy9nul7h0wsjr6n4wilT0y3Bk9AK9e01
qItpsGDFcJ8z2o20xiyOhZfQzMK9MtjDnOeswHzI8fOgLTRlmpJueZMckVawk088JoM38IL6xXE7
oHovGkyfKDiqeze7Ud8FdVFCLt/B1VMUJmgVS44oH3mllma1sV6Q5NFSuNqk8MPzKmkA9c9iY4rk
Rm3aJM1Oe4KrpObaSK27WXbF4EWXEQAbBPBggjoYFX2mAOzmUS53+rG4WCqFMLPYKjXPhzEbUYQG
7n/xV02KOluCO/PybJ4qjNKqgiBGo5m0HZsDbbA6Mef7gIykHlF8e7QXesHXfEA7vsfLcMoaBx3u
P62/t9u+lsHTYwlmuY+S6UPDDwm1baJ2sS5zWrfg0OxsXFGx36bC+68VIFdeA9PVXDOlEQiBK2IF
XlNT2FUt9YneRpRSRxzS54Mu6lXH/QUAQKATcUZYuGxzzIKIj07x0iF/fufT2NIhi+OtCzm8eoo5
OQhsEAmKIeAqg84SISAnaL5j5lDvnc+Qeh0p9mzJu+9W4d9C5dBN54xRKuos8lNjVQKEBG9PMj7A
HxGz7Co67d88ybN3ujVWv9evA7ZyuzloDONb99For5dkxRkMm+EOM4LQAL9JuZ+RI/5ZokJdwCbT
qUmxbCwQEqnyg5wZBCXXP+G/BJCaPz6S+nPGVM3aG7cGEueYeJV2vNbReHMvSswGYMz2+5IDU/X1
hT7thlJwpbFpJn9/PW5r1yUu0hxfaL9zHZdGb4IBUO+aSdcpcr0IGhs5UYiC+NPBoRXZ6/hyYefo
hVbd78An5n3rKkPi3N2Y4OfLjsynVmykxbwHKZi9KGZ6GMvS8IuvlOPAT8idHAH/Y2Xiksz1xOMW
YsUm1t9dvKS6HDLXqruuuTrLLh6NHRxg8Yp3q6CK3iJ9zlhz0wiYWGFkN165dIAnbEVTrkKQrp7S
Uf2ww88C1V5X1T8QPAxOGyOdDkTMwPaEeczGvUdLXfNZ/IHDetWThVET3ejZv5yXkTSHErtRXSgA
hCQk0XVU8ZIM7JvZiqQSuVpr2yuCc/l0eCuf5Ksl58bPohC731QwjZzJNlG4H2bTj3BOYbAFmSO+
ceuJ7Q62/HjPzzkiU0ysRFdGDTQkzpa3GIQIOixLS0xxMEYMLIjZB0zcvYaqdL3MNmv2Xd2ImX6N
zYXkXzoDrheqTy0kQX1vWd2PaIm6qiz+iiJnxSPGKpfGJKo572rxIF6Juc+kqCIwWXRPKL5eXrHA
T3sRAqTnlnbSaPx/vXGG+96lMXlP4QYpP/sG1EWKZ14ihibWHTctOC9LBW15xbOC5AuqkHMUio/X
ALF7qdCkhHxl3v7ahZAuSRKLnmAnmiLVzDW82nsbY1ifVwpNGho5Ngjj/GORGM6kfB9BSWBqbm6Q
q20EWdwVm3UzaLvkVIrQnQvNY5spq6nrNAkw8MmmMyZfAxNR6k7Xj9FVpWeXPwsm0tTLWpwSU89P
pJkfnD4fA+tfbWk4lQZC7GG1Um+likAUZcz2/JdZvsTv8whh1DpewnR1OLVvhYtvouBJypbOy7P6
oNIYDTI15r+/QIZXDx0rC1rwIDBJdux+O+j7/7QiEitDRcz5/Ylm5tWMYaYcstyfzlBmE3pIp7sI
IPUDuHwyiUUrTCt4rvn8hz7G91c29S2IMOEX0ysRl02SfHWyh0iLo0JST3FwGnRbD4VgXgaTFwJc
SK16hqe4sg4GYP81TXCR/Q/CcVYn55jAqpOWYeTGb3nihMpwgCVdoVg9nfxzAQeoOrN34EkOBxHk
XT3h3LNrc5BgNxvZl74631qNiIq9MpEKM1dUkA5Ow8Rz6KcPYB8tonKwzythF3w4qaOVg7J92+q9
WqXkhe2HajlKXHyVRypX0d/4SB65vBZSbwDxJBfWzipC7XjxUX3bmu1zKG0Enj8ndUlnysIAbh5K
I2VV9pYY9rQRJUe2Qk65UEbLTFzaW6YOGJzbwMHjUVF0XkDbp+Hy3sbFdGth3asXk7ZtlWFxHpUS
HekCOdnHCFyvGbTZyDd+rpM6YB9cCaegu5p+uiIGtUpgvmngnLLh6Z00XSNt8ojImc4HYi12WNak
orOnkknV87rUYQnjv77Ut+QLdRScJiVFe4p7su46xMCsIkpCwKprA/YpZGgE7DiUhQUD6Cbtzi77
d8jdGX1GG6jNC+oEGMpLHNO8Hq8wXCBM8VbapGwqTOTUIZBQ62NEDNXLDG7Y8J171+pBlZkBVN0g
4s8ouQNMTZZpr4a0+9ubv1qsyguAM/eieyYK5j0015+zsE4jVa0o19NGEDEIBpWwhbSECuGOfDXc
UNjdOknl+WYAo1tanReYnt/5SmInpkc7Gqp4c1l923QkM4eypXv+7tEvUKLgpv/xEd2qusidhUN0
DMfaeD6zNAG5S3sSYeZuGztXP2qJUHNJZSC5cPo5RVpsngYD25xbxGcMyjqqKPmQRhco82A55gCL
zUlSn2QEGsok9ek53jq/noT2kNWd0JNBNnwJX1henTFstqqHKVuuBMGVuJrFU9wuAuN3uPzezsDr
kXNlUw4u6fdCBJCcvVHBXF79jA513yGkcZ+C7tu73f5RYbCN/zZuSJNkclL6tiwdT829HydiU9LQ
B+yetd3SH/ApEcuSO4XNVboGX3LHH0clmqULbM/gVQXpmzSC8oDFKi6ld+LDfM5IDfM3zjTABvA6
/BOcgTiMJcqepSfXGS6UReG9isN0xy6OUog86tGNKUG9w5tZYNSo5pc/CQ94iAOTVOGgaIdq2VTX
UfymuLeXI8+CXNtniRiGvJpeptqg7uc9dIvpZgJxgD+yVYSAMOIjXs+B26Zqlj4tv1eVVWIrJ9Al
1f85DCtuiCXA4cwYAeTr2L7qx499gdN16IyoK32B0iv4y76XEPxQD6mkK1JsVaaIIo9Oqot3gcmB
NkSbWzViUN4cSYNU3/aM+rhnNJz6PchKQTZOUUOMsXCWVmJwTD9dKIbiFpRDTNBRnxOaAl8YS5zj
bvDfnBqN9X4z3A7Ij9D7C3jgVxVt86ZijyltHrOC7sa8YvCDEGrrgaDmt06qevasne9BnDCH+E1q
mI04GAX7AW4G9fgjuiUQlv9Wjg+c3WVJS1D/HkN37IEjMVfP3IbaifNDu/gK/Vz0UXUh6UQ2chPP
n+fzwZ1Do9fmoZ1rwrGEStQbNPvo16VnDYradZo09ch48P1ioxVzb1MgYifgHXoT8ErDgvZIekb1
pqnNOQo3XV3Z5QlnJ9VvSWcRdLsqFlsTlGu4aR/eW1kD0kkC0K4eFZ67JpbBt/uDGSjGwUmrUSAQ
N2G4GRfp11rzXfKhXmUntF9ig3b35S6We1IN4xX91bR364MJ8/3m/ORqvmeejjN5E9gmzqbJGh8k
Nfr0y9X+nACArc+mFXcwiLp3MiqAjNlOBUF5VSE9vtwdmFWVhqKRxtL1Q/FLdDeOSsWEUGrpYfn/
3qIs/xYIdL57dnifLNl4yHa+67TWtkhfzA38dCKqhGt2EVdNHjfqeOADZjm1lUjAEQfnBb1PLtg3
G7BtdokvP7l+QRRlQ/TWmwQtGg79V9V9HsbylN2+UCRVndM287eiPnKTDSdFTKq5LzmX0B835GKo
VPo4f6l41zJb8UYL7MesQZnJwH9jXjaG1tzVluzt7fWLF4zMCDKbCVuS2X3GzFTh9QQueGHF/ra5
gaOFgdjbLK6UT8ECFmHyOm44DKkfxXi9ksBZPt9Do1dSw9XV1QacgwVDiVDBKbaP7OuGjrKQtlBz
mR7dmr+eLR2QiZfiuMmHNzwyDjXzNp/6QElmT1IJjjQA837PrSdgP5wyKpesIxYo4eFDLKPQbPwm
J9lrlEWQ9RwO6s1I/1iNGiFhhnYv91rc8pdLPXFhEi1ErH4B9jzwIJj8Op9vJHKHar2gRwkibe+6
lgMzb49WevRqQnHUmWZHNzFKVp+oM2/dwQcI7RAoUOz1WPxKs6Ug90iz+9R1YvDuJXBfrXJMt0rq
wC017z69e3BJSCmSyBSJC6EMiwY+/DGSNIhrPf9wbJNKFt4UQkAKRm8DjnPORw7NZ98tzEtLiz49
flIxkZ33XUWz+dmvgIimFYqJU/yJDU7UdScZOGHs4DfyiBGHG5gCgZr04rHUa4Yj2ooGrOhtiE3U
Fkmh/DFn5LW4fNkJ3qxXoD7dj8O5PRuuqR8UrD9sPN4OTYe+wywM4I5Su7BFatlh5F3+zQiYGy4a
WoTnMoWytq4t9WYyrxBF7hAWhg6ocq8OpxKrs7C/gYZcBYV5cGXB3uVIWmaRSa4FqnH29bzDzjRz
/ZJmDlZrp3Y3ZeOTnY1hsjkgN9Rna+Jp2OcidYywJuvdarjvim7yG1tG5K/e1AjwVLqYsPMrAkbA
pMQa1P5y7g/1wIDdVU9P5+4hUANWZw96bM0gqTyTj0DLNGTmMuuzdFmpQUJan/OrZqDyd9Ce2K77
jA9AscGNqwnHrlVfH/bG319mdy6kdbjKp9EEZ8oE1zl7AVO11Q1OQiWBAK0QReL5oTXrYppWpkKD
VsmIMG5vdCr4CW6O5xLD2fCHlMTWHgqjbqLiPa8rLhGHxZs7L3gOPVeBJMAZsVLtaOxREKZKaES6
pz2lEZ8MRLFYgysEup9lURZ1Jsl+Xpy5RPlt0Q87i+zdgxzABGZHR3Z+/Ubv/PyjFh4HiYLTzrca
qlOH61a19Gy+WlUBskL+OXVBW07UDsrYXt8NWwGSu4Ai6ED5Ix4BDRXzv3E7Q1CXbTyg0UyUG+BN
emqk0mR38a05nW2XNw3oSqqvERw8T0VY03hpXDDqjO9nBHG6WIUPYyEGd0tbSMJvIP2r6+cCXEI6
ORGcds1u3HfcmjSOdE3N+2VlxEQbs9WXRLQi6hUGcvRFxqib4wPVC9QVKGykG5F/YGdwLOKkeHJB
NwpB/CUC86PcaZJVICi74BPccrw1oY2KeeUcXVkjpPkF1MaU17gU81BU/cpDKQtsU3KKrbgMMkfr
Spwqjz7hCoU3e1K9fD2R0+ohBwl6EbX97HXFofwC2hOhTYxjvbj/+uLNN3pY40Uu/ViZh7Lccie3
R6aniXN4lUkYxRy9gRokne3n2kWezdhTaQbBJyY1bRyM+O/BPyAngZvkK6rlNchKpFodggqlfmlv
SNm+s+1g0CuH0f+7BT6qEtDkjku/NbYmrv3IOgK4QeUV7BymrzpeQeaAgPt1FkSoN7ECWiix1wNM
TTVukvEDf19uQd1t948g6t/1sFSTojL/39d5TeDyjg6VSyslVkTupwUP73xgr6YMnxL+I0A4CeHE
iJESmorCzcNc1ea7nHafXoxVY02Q6p7a6yzbdk/VqV2KcZKpVaMxhDBYrMZgJp/YEX83Kfql5VYo
rn6AJ1CJdgDZ2jtqmYTxXnE07P5jmdXQt1h9ThaYOFGPQ/3k332cLLxB2LtaQ0yjG/+i55igriax
afxSixYXTv/cqDG+OOmrksTq5ShC4cuj3Yt/2A7JTjiScCwDZ8CW0ZwVE0fFDrR17vbh8sS6kVrV
5HGV0KljYO98Oq1tsnqftGRQYuLHZFtNdZADSMroMjd4Ba8wOzOKw/tCxh5djJxUcMghYB4PGo2y
6AvgDWRy0QMdmUpoHiwyThpy1HMPtnCRqlypu7ZWviSGdSZtOaIaTt38klvdpIrCnXouBdYvlZrk
qBxcOMUHjyivQmiKl5RtP+dGvfZ2yzxgvpU+mUrW6KU1pbX5+Y0HXuMwtMoZWhPFHZnIZ00o56Op
ExmR3PaMJXtPFjmIHBMEsdy+AyLXgafdWeRljG1szKGkwXfRQmHdkQQJ52B5xcodOfYV9Lnaldgj
hq+L3bRcFPIbm3Gg+fFz4YVlwIrWy72z08XUpPh3oVXjY3q4R56N4dMhwWIAYJ+tbOw768qD92+u
2ISWP8C2UsWXUBDDlmFzGk0k3Ar833qrfKi1l7p+04sATIVI6zlHDiBFGbPK2RkCOkzXQxMXBw5g
J3KuMBSaQd0NG4TpMaxMskQUXZyhJOb6m9vx/6S/6srzFy4rhjUpFCgEBEIGZ2O8sEwP08RdqDpE
rMKz+nVbSSrGV0EKtGv+6VAgU7qWb5nInrVaQHbLTG9F8RHpGzZ+XqhvQfvWndtiOlVem+qzahnr
G0vwrc7cXNEgRjrb0xy7jga1lZXas/xIArf/lIUvJOqo5w5RV7bEHHypv72QA1GPLCAvPeuTn+GA
YzuSsnwm7T1RKqABxL5SSvzuVbdL9lo7oBkHsQeClIaJqffNGYly59lZKAhYp1+wOwJw7P67K8nI
QkWSGWvB7MKMCiocwMyq7E+ijah4+6Db6kgd1syI0dRyDLpvLdFUTbGt+7cVygSrK8Aol/yeJbze
VL09MQDQu6b2Fiudp8ZzWXXzwSFrzqb3MShT3c599aQv1CHNKp9jQ6jmswmh5jXYsGvCXV62y04L
tYlHs6H4bn+Yqz+zqmBi6TfxLDz5QqZ8347zAOdC07odMYleD4CPAWnVtHtLnxknkCp4Vsj0nIhv
1nluuKkbgy7+/qJpAXDHV8oo6mA5dOfOrNYFiUh0PcqYM4mxe3czEG0gGZmx9KULdrWkATu3ZDw9
xTBErbvd+LmfUpmo/3Wh4ZArXVu3VOGAsC27Vp0RuMEyCs9v3h6lhR532Jov6B1ZAkzPR932SMPK
43ChzSzO+xhes0XCrkqecejOeSf1p3Pn3uG+uoMqzgu2Y7Iyb6VnTlvKm64aA9nLPkY06iP3imBF
DcQTNAjEBC0PZwLnNWAMq2dEIumsJcTEPPU7HuUUCpvtQA9ZW1Apv4QKVR/OYM1WV7hQ9/VZgEeF
v6h/f5Orm0KFSoMPoecswox6xxNFsV83fk3eCDgedyXMcDv4X4t3K/OkcPEH5roNzmkkcqb2lQdD
Z7iO/nci9eNbLzIRI3CU/OHVdAG7QsTRBj1GaTeg/QItzB3IcBNvR8H7rxCKZ7lWXW++Zx+Gs/Tm
YzLmr4EUHRCqED5KUuLGTnVKz3UoZUYVJd4ymlJlOXZrJ8Ez48bqdTuNKPv/solF8j785Cd414CE
40RMlXlx2tl2xf3jH+wUCy2oPoAE9IJu0BUcihcFcuANdmvB4k2x5FVAV0WbE3gBcIAhTY3s9D0d
9G/EnBG29Xt+/HppNT4aMB5VlJXJBLijncytblbTJGRg5edugiFA31Mbz0QVqkkbBwpCoVx0Weso
JLP0zomG2z7tMonh3cnb3QbxUBlFP+AGCq9haGtAu285fTlT8nluxigl5YOnqF7YaqBrFkIBjc9X
L5rx/zgbinhbjKiZvdb8HohOzkQGOnedRCKCLh2d0qkk80YKyx522gxebTdigvbip1OneyYVWyAG
QXavk2QLqgrD3fs5C4sI0bPos7NSvwp/xuZ0Q44Pek4z6zDanbhGdh83rtL1x5VzaGFPtTFcaRXB
2u5Vd0AklUbaVkt6DolFb5B2WC6+Rgfg9OYb2k32DjLPmaU+K+o5dwGfLxzhCofDD7Igza+aQMbb
Y7huZJOdfq892BCSz4LaSQafColnO9tLESwbHfhZ/xUq1tRdxM3ZS+/rkiWVl1yhtQM1kiDdGJ8R
/jKTLXBy3HBQG11L+lprB2oZMK4VaKelPpaqYhyTLHIa9s3TGxmOH0PckuqzH/gTaKLKelbtdMjC
v8bHTSjmKrQdgJ0lSk+fO47plhZBL5klSCg6nOheAta9ITPKTzU/CvuVTbJCtbRSW4spcFbTAQ5Z
BKfowY1x1fKlz07hAcbbmlw8Q+02cIj0GuNAYk/dssITGbfVczu5TJHr7YEX3J1EAbNJavYjYJbc
uOh3nLvL7sM106avxPnz49mV//rCSZBcoY2UFSdnmKiImX2pCav3P66Fi4WkR9jO3lM8sAX2XKCL
LdiItXjRADW6CCdE7ZXB5rLWvYmpWuKfv6kwrQ7xjfNBs1H6aBJTUTgYyfCyiJ1AOgx6pU4Ov4Dm
Zm07eqggyzEKOP3iC7gWmxE3CxcGfWZvOP+TfjvMbY8o0YnHCevc5yUYQQCxtKg9JvMjlUaKwKni
IeLnp4bzOCmCarAgF6lDxSWUdXOVebFlrotWLBXNbnb0JgockVGzaqiOwxUhg9sr76TlLsoz1zrN
DKsudgirJlk6h0GsJiwvLQ85FROA1SuLlqnZqvBRRjceiZvBd1xSbk+YLw29UbhsyI6nUVMvVoqA
Yr6vSIoCqisNRsnNlwAhg1CaUQ0d2ZlOzKOgZNPNQc7OfXUZ/DsQrNjiA8gbDDqGeSh393NhOVSf
JRyIS6m4IvflmXAsZOSrwPlHIFynnaRkYsRtFYOIDiyZb+xcDxlBbZlzxlmSayw9Ygq9CexircVw
4RhwkTvbqTYBffrME3pFYRx4QOMcd+4AAHwBxkW8qeyPqLqYGJ0L05wvSXTDUggDGW9xGyYGOU2C
Q0kTigw7sVXE479m7CvHl2es1VNdnZqLkQzWyKOohtKf4zlCoqbdWw5k6s7WAbufhFzA1G9QZ1In
qyl5+RKRqJmV0nLFDQsM9Er6U7QrdWD/RlUG/R4LmvQSia2Qff5ynKh3rBhxeee2BO8pGJJ2FozD
hT0PxnpEuEH6cAbi5NhQ/xbPt4Be1RwVfVdYhIGdOtVjtp8TAqkwSmPuR1IOQ8jPGI0r4iICSeM1
MRGYYPdt0tP0nplTu7IhXsh8BQ0dspdnKZMmK1Qmm1HjsP93ba5FRRK8OR8NpICQDR+TyKOuzy3R
wlvSCTXhcDCAbxVYxDya247JUAsFSanksK6Y52D59EEYrWwRFCl0xqNEEte+zXRXcaG3akwRs2nf
/ynu7j1QiedkiQ82VQPQZfZHk6hfDa/RA/O0toOBJ+uApKRor9oXOSiefrJexXlR7W8lKzOWFijv
WwDvNpmPROv/Vbdz1DZF01jcZlwnfWBuyra7D7eglJrRdoJN0G9CIYbGrIqtNJAUREGEIMDK1zAU
k7082b7WnsBLJC5/xfGLtMqwU2xX/8smLlJaZ/pdGg8rddWtFi0WnOqjFrc5K0h+B0y1LYPrd3t4
lkAnuQKClpa9rkZDECHJXxD5xziCX/76F/Ah3bItvE9MLI0JQwmP0b5/waM+G4sZo0OVTKbDO9pQ
cefJghkOh5w8TWs7ckAuIbUGqA9GprvVtDkU2flprp32uIhHD4864LbVaIpeT5a83ZKgINx5bs+K
gXstUu19gzLXL8uF2V14g6CE5mX+2JaMklpzejZ8cBnutAThPrR952WGqzUHydiRCzzlIruwjau6
Gpb7bvXuux/S1h5ZcWKp6xFBSn/HM5T/h907v2DVIjUDHuvd9M1EXVmGPwcScTr6pqI6Am1tzaj3
4lCip0mKC8vXoGjrMlLAchO1SrF2YwIqdZHQ0NoFpG+JIIGfbOXbqOzWbMvH6USpEPLjGw7rNytE
lCjDUXn62t4vF/3cBcgAi3J9D6LXO52CT3h9MQzCWKHTUB4hllddsQT3ITcayohj0+bhObynznUD
+iePV2mrHxgZQdUHmRVgr0lMWfgmI5xN5lM8ewqnzgaFlsVmRbt6fXamyARgPxPTY6bYCI9KuZKf
z607kXjBh/AbzBxd/e1Y+HYZ1c8iNAb6A6miSQV9Tzt0EQzzPxmvUl0A0hd3N6bXXcsFkzf+FmX3
BiqpFqm1ovDHXVO9Un3qpdLBJjumV8w0acYkG25FdPMvhxd7qwZHb7ysjzE7FMttCiuHvt94cFEp
xZ53KNLSTqHHqG0d7NdbY7qJUcWbhg8/LpwqS00SoMk/AgMmTj0eijmoC+V2/EDkO2upCFmsbNcz
Lay8Kl7/qApQ/XxMSTDvCrdbuTmhNacfiMq21KRMCi2KDXDl9AvylNiGEXTNYEXBbjea45zVO9sq
ucsG57cK5DYkeXVOs4CR6olUKtCM5xaF5sN/Po8j43QyVtDV/KIZwoGklxVYLYul8J1UqLZNpp6m
nhx730G6NWUpBCYC9H2AZhdoJ6X8ck4uP+SskLHYTEYWOzTfeO2G9NgWnFbAk7cISzu7ejsGZQ2x
v2S1eEK9XJ2aF7AsrkIzfBmK6W9KUIDPUGrZ2zKuVApB3LSOaZNmkRoI4YtZcTTIM66ihwDBqFnQ
NP4eMuFeuAEKT2Zi8ySKQUffoiO4biQtHjUV3z1kuQJat2zPb5bTCxT/ZbJXCB9TVzj3wBXgAEod
O3V5CxQz9XWleke7H0MusmXYjcvlN/S16pTiWRa6AkACOq7sgSdnbEK9QUFfR56MYDeszWEdlnPx
emStxqT8uSDFZQ3jqZtHVFblbTtR+aQct0BGTpbshtObhZfyeZa1p4MTPdWmgBlM1JG4av+0YzyU
GTC6T6FlZvczVUg7Bzf+IH228aCzJrz/V1GeVwa7eV+TZxy8p3Y4fi3Od+jJEICi+Ms0KPet7/KM
HDWpPE7LQF/X06L7FTgzaux1krrjkUYwYE3fcK9LunisAfqxszRlWEbkSUdcU8jdpGBvqBmDF8bf
eog59jNBWlNa59muK9QzO+1M939T0kcwZkvVG70ArpPEl5znX++y953hwk0WJ2CYA6Tfp4kQ05u5
WZfEsgO36naX9msZs92Wgbg7/L4coewo8jtuLkQLeJDCUxlj/I1SoKITcJU+gXjBcSGB4FMGldb/
z37p+huC9jMIN47XIcfYhkt5gznoKmxjYXb9m4jxC80dJYjybkFSIbgQDwHsBbd7fdb5Ib9LzOWR
0mNi+2u94som6sEcCW2AQ3DEyKCM2DfyTZDzsOvEQxUpvdNF59+v+tBIWa66DnfZrvPjuFSO0Uoe
dP0OfF66a6VvHSShMO8ZPn8TIqtrDqqJ4IzHkRFdE173zbd1LW+XlzevvYD0ks4wrJd97bMcavh3
bD+MigIPZd94fLDIJ9lQM0JIVcTfoCypSAixFVrMpYyg/IJoYtjWESy4ZfobsvVyo2v4Y7AqfyRD
yyO1C3baySryL9mdPwXr9dUgeqOyo3DRN2ZbxjYB0qXtcLey3fX5LRj7PdHY3Q05i55Ha6XKdp2a
WfwtdvOHQZzNJY4eHd8KQfFQVdF3uz5rjkCGQGQaXAYHk8BVw3lKEGbvcGhorrHHLAwA7QddBFr4
OOV0zV7xQoKEvFAwKbyfkTS/5EP32exaLjCxCdGEdlx7bL9qhDwpbLDNZmSH8b5dqAjviQbkRNy8
RgHwUR5iRa4j86PuRA4RMl31HMiwNhEAWWydPZKssmaJttZtwsodT5tzNaU/pVUwPMEVJNTl2qt2
09Jg5aENY9+gleEnepXm08uVuO7T9U8+WLN2B57jFpI0o6W1n7/3pBDTxitJLPTMVGVELucLKuxN
dqS9HSOLX/gNEl752SgmG8Oi40egw1IWXIXh9IzK6+Fd9NDFZBSn95O4oZvMpSkT7iRkDzI+JvvD
Mw84AdMJklewkZCi1921UrOoRqD4ErVoUPnBESsIrMGUQboksINxuTQZznu0yK1PfImubuyxy9DN
p/pyML9ICq/xCmzJfl5CT1ktvB3uM+2mhU/2i9nZrBDwo9lLS5hNWipgTLzpsox7mrySwA5g/QrU
bpSd29PjtCgv8mf6CW+McF/63sxn4oxo69HecGkZiETYyl+k5mO4P2VLzDnQ3SwG0P/P5+qK9zJy
S0lGSSQOl4paM2d2Mvi1eZtzTGpRkLcsKucDHOcdrW8WBSBTii8kr4MSDokVNShbfxZaZrxmPscF
0Ls/s6T19kbiX39dHW4oc+IPu1zR3fMsNlKifMTfQzIQpD2EkvwwK1XzfP/l8L4VGmjblZJPOMZ7
G4LGuotQFqNqyjGi0KL5cwFdYHO20uiknC4M3aR1Xe6fQM8avdgOMd5yxXRQ2z4c38HyKpaDZoDY
oHp6UQlgP/JzSKnRlm1ZCHOBlwbzfhUPyOH5wq/Acy6mnwiy2JChEGrptsZkZYyPMO2ISJMSh/+C
PUrsVVCeYWXRsiCYwUp30rEb1NMUK3Njxb5uR5pRlCdST8opjy8xFgsc5kZXhY4RGQ68cMtLrHml
7HdtIRLOKzVfekPa+gScUaiFjBOOYAK6gW13SPSpmz/rjObykKbWZL+M7WcS7j65gAZ3v7L/2Za6
W/7bWAPNn9leoPtjJ8IhjG+c+gIKN1Gb+Ep/IzzehNfrMmkFgHk2QZiVmPNm7Yf9Unhzzmm0jY37
zB9WojE4EC1RI1tH0ZL5Qg6YnjqGrWDlSHnhxjwiY+2GPJPjbt7ozELhxdw72P7P5wPWniuW5pnx
MYKUT060UZ0RSGQ2Oab09UMNYpN7H/2JcDQzRd62Tsqjd/TqIPmq2qwTTvU5iubJGO/J5xeSeVRw
g/Es6t09rwHT7JBm7uzYOJlcb7qzJicHoyu4EcA9Q9aBKdBoJw72VAuVuHvxMmeLt0YlQkeAmnu9
jrXqp/aoWF6QLLC6XLyEdDgxzBvPpTUMGK/WbDdY/W85QBCpunYVOXiG7nwb1C4kBnWOjqQXkRkZ
dV8Ap5SSxF5BOiLeRi4X6QZYjO0yRV9nqdikYynRYydjvQtkihTVUsSBMC7TyWUurI17FbcgEjii
3tNxJNRwmD3emmLQQ3+c7cI6H395jGzTf5zcnfTM2r5vTEJB2pB3lxlwzYUjpKZrXCo9mxGf+w1Y
nlRs4/rN4aeIcfXBK+yatcxeiwiX8lkiymedpFTHya1hVOwWCDqEey8TMVAAltvLykicFtMLKJiS
iOQech/Ndx8AASuqXuXKgyUfgAtZzacz/JJh8VEZAz19vMmFEcjoGhWzet12HFDxCeVgSWZAVGAM
rRN9zdPPAvYQiizM0s9qnlACh8ZS0wsqflJc0J6eVu/wCKOiQCUbUClhJEPofyoZ6Akq0CPADezG
rnR3MFaFNiSefu0hhKKSraPZriBvyXWlirv8Hf6jJ0HEV65QYDtzPKA/+D9xiyR4BW+LaCN98Ia/
ZuRTjw+TzWYrvMvgbAX1ZS0SDplHNdCIrEIbWeKccjK5BTOo98Psyt1BYLZK/xSMzkLoIMK9zTsg
wL0En5cAavaItU/lhn3DjNUoDda10HBD8DRQGxq1KW3QHOy6e0JYKyQT8dWFWLUYP/bm0BrNYkWI
MWntLb+vSeHKdQnVFE0WtBI28ilHriAuETcXF16XdwTNHopwC43ooU8CLf7FClrcOk6VHbHzXyDD
YhxPwiS9jB+hBoqmqMzsKYMJuBbTUUBnPTRR9BIcbs1dlhjjJRbGtDmsF2GUxToSyfIy+8tVuLqN
I9O/jnQlQuzmcVK2Ps3JTJB3+9Up/5YxPWm/LHFc/puHxEuRI7TueFIvTOHMndejMIfXvrZDk9Dj
mCrMs4H63xnwpf970xQ9TKrC3kFwLrK47Zd+RKEBOkuTDiRXsToAi2KhprtXGXC39WSJ7GGbC3yF
oI61eGcaNXz0qH/lkjPhpV4eGv0FujQFiY1LdrH3TvFBHEcuJ7E1vzpmplMFUcpf8DmjcY9cXkA+
W29WUQmpZ/SO1xe3dCtYv6GjL2auzd1OaBiRSzjQj6iCPjMdWt9k/4T0vvbjKczW3u5vtr8PPQ3C
uxDENj9WI2NPezkQ4Z10jo/tQtMda2IlvtFYgTfvpxMVYlqFuwtdik8C7jPnHuWpdfcknQiwfXxQ
BVwf7huJX4xGyPdgokeOXDKhISKBf36iQEMnX8XtshHnJl4Se2S61kNox1UI2GplU3bmBIX1yIvs
29eIpIVPrufoVasdgxmJxu6SmZS4v0qAPHWtVSdYhjZHyTbi4m2HpxNfnN0xFvbuiq60Ety8n+JF
jinYEdM2246X7h8/gsvVerzNAean26mP3QBLFzQoZ37ERLVWAmIioHsqV8cCn6KNC2TKyRCj4N3M
b8xi/JL+yYNZOoDd4c+3k+ZznbOPE7Xu1NMF8RtqSk6kg8TfGpfgCBcsfOTBb5UGpnqigvY6D4vF
KJLgYGlyoZShFGqRdlnjoynak4XuZaykzh6mSC9mn3cJzusQaADNm5KD/23+hzCN8nMCkLJhrgc6
GgGWK0FsWntNpdlVYi0vys9/JSe6Nlg1voq9o/JFr+8s2v4xcSLG9w1riDrb0DEgtgx+mv3v9qO6
EQJq3YdMqqdSxBJXM2qeDxe8UeVR0Qz5f2qKK+KPYItjbyZ2zN8jOUC40b/V1F6wkCO+nqTAVjH9
yRwQ32ZeqVFzFGIrlNWj7DqImAsAL/8p8yWSqKBTa3lS5tobfYrYHNxFgK5CBfaV5pJBtjH3CZIl
BONimmC2s+L9eYDrSyw7+tQKHgnqrWAKaYFCZNTbaoqnonvQtwwSefQcdaWuMZDxZ0ge4LkZ8+6q
Ijtx37YMF20K71o/AFw5ep63/TvGsPLhLwMRlIQIWlbI1vL6bbAtOY3IYN19CCi07X1mnEH0cqET
6yrSaj0JUpN6LIOSyDFV+1x1+TQZYeAGU24r3PNLovaKpsJbf5SyB7XGpj2cDD9cK9QCoTgalElz
cwIDiAV468tl1ZvOgnkFhXCaQMGPA6Fnuyy6vCuiYuTWMQAtiD/w7J5qVoTfdZQSkZCKi1N1Vali
0kd06kH8JBFPeuhPKxoidFDSjcyq6nhu1RJYckLjITIk6OhhQNpXGEaqRz91fxL035h/Pj4E0JR1
8ND0WKgwYAWbRfCLQHzKS8yVNhyWW0CLo7VXft7VClh9FNJ7y+WF+u9VYgkRd+6eJkVFZMUBfNap
5PCWC4H1OZXzvMkhSGDDcaEUuJlteWfD3Gj60ockiBuTPXLkNBHeZn9b+uLN90BL9XBXWRXQuvar
C1z8sUJXrEF9AtRMbg5eAsUv3sgYxdP7vP1PqKxmcew9xslobYX2lU2kHPeSXGtzOIrBfNHwbSpe
LE1DhH2HlxyJx4q6SGxm/UCpyZ+yR7T6OvQlWmjbzaeF6glePJ1Wv7SfOTBHnGzl4U4phtF7IS4e
mq2p0nv3YwUUpT0bVqbYm5WWaseeYCEeEOoaQyKUSCQrTTGGD+gN8xnhFpMh3NjL/Qnm5e5NOi+7
I7GbH20rEATanJWhMSFnZ2K0SvdpRhmGNaBlsC2rQVstMkf3QoVbAPLALn3wXXi7Jx7OsNeDzy2r
WkgNPLWpCayFY0OiQIanzr4n15bZvXldZ06OE/v+NKtmtDVRbhGXCftdQ46lmt3Hw+BL3kOm6u2E
97uNXphNVJyze7WIf6Pfn0d8k1D0yOE0Q0N4CGm5Qaed4mRBzgCQ+bi3Gu8ZFPdBHRPEwmJrIqa/
fxiYTlH6nqzLzdGUtlG7/ESWR9m8dFcUuGC3xAAnLeBjCL4TcrGDkjSVkfc7Bu+CD7BDwHUuC8rG
ER9yLJpvfQACJHvihP2zcsb0RGCyE2AAi+DlqHS0uQbA1XoJMhM9pkK+mWbaYiq95iU66NWQCv3o
BbVKvMJ4dNfmgHHLfSa595E97yuhrVmyqhRZBX3rW4rmz3/EBLrVJWgK8XXDjkG3Z1wvUIdaa/9t
2GqjVPOsaEu/5T0hsVfdnv2htzehXWP/zNr3OoiiRz2HpcC3nA8ijxmJkBsoRF6JYSxS2ujGOKa+
EpDbkMtVtqYaUiabbyvg6KtJb3repvs4zhl7+HZLs81btwjrTFYiliLpVf0RePErl9CQr/cA76QD
Yyynl1Y1oI9jFKLEnVOk+lImikfVN9A4WPSDN5PmO7S0UJsTAsMgUzpDOCBpmc+A7N1SwP5sN0B8
9iVYVexfL6eA4v8PM5PNDEcn+YHNNI/G4iQQRiiDmdO0CEtxr7CEWwX1InIB6K0cswdJQIu1l0+G
lVvtppYkvGE6dywdNHyjrqJ6E13avjKBGVPcYmFKRTJzgJHPTf540pZMhPFG8FpE7TMwdZxEn2cq
iBS6vPSKiaX4sKvpBr0ahKQRPoSqvHA3h4TYQ+5gDwp6D76vdP2Vn0INruG8A5fj0ytpAYtFSR5g
eEO7iUUP1aHrCyU+tL5Dbg/w/IM+l33lpp7qJ+RLj4kW8mqZ4RhwyGM4yaf0SNDNPSPbI+yiAkFb
MzN78arJcz0UyDcLi0njAQFcjgyHWRwrw3gTR9JVquame/bILJ+c+uLLu0J/XKyQMXUMFumrF+em
eci43ya9KiTzXCK0ix2i+WkhSgGZq1CVMVBAKZ5CAUxYOcIDlw6C/GfYuJL7tgo2Iex8PkfSpcVW
Y85ZkoCELQ2gk/05y69mKVreJJmAeh9zajMdCBOV9FZYp1wouWBNiTfNeUYTd7MUNbIyax8FV9Xy
BoMCq0IC029tOMBQWT2EWCLfAeUI9h9vao8OpW9d1dPBQDbNs883VtV7QEPV8iENGR31XFpJkD6I
0xw3RADPkNquLTHLLdA3rLxxfd5iYqwHYhM1iCEI20U4F3Jy+n39F5yGCeZj/UuTXUSqyUWwg1Hw
IVtBiDwOWvwr2WMhJ1ieRhRN90cfKoPxJwvjnCBqRx599DiLFYSpEPbi5c/oWtlMwXMtBQueDO8t
5vYP1XfKPZy/11Fa7DgK8vKC0IUGKz7hFHKi31cklGuEBYsGmQGkElcDKzJnqYlmfYjbxnzjN58b
+Tnlk40GKTy/DvXBQJYcxR4/ksurkvFQ2kN3B5bPEy+YzsjMEZS13fo9QYBdCZuL2o1vOjtYjDpF
u+ZQMyqAqFiHmC4AdNig9n5/RDV2OPftrS0liRlpt+YU0lJQRvH8yBpSMui8IDjJWCxEf2s0/KBn
3U+kvyxM39WcbMaz+ksF0gqkbRklV4HWU+1EM+pF+bBwV45y4PTYqd3VpvgdV5ejpk2ibNDoGviD
0K0GJ13lmNOSV0+fAx44OYpFOVlAauOYlsQ4jDckFvsMS02WQjCKGDdjG1hAWrp0wnhSk6XdMZXA
C+ZTeM55LBci4rA8318bpTzCxt9kwnc3pkrjVQAFVCe+xiyhIBOGoQUbo4sb5P/5vdsYrhzdr1bH
WsoHv1vx4GrgmxXY81qprrnmQQOSSJdWH0i1uyiUEkFSRbAfjTdvEy5CZt92bcL+3C7Zdy8pAOuy
ZQbg46pKVIT8+NfHrx0JolkPgNKWpmD3f6SVeB27aGgslutdhY2Il4n3Jzeinh8MSpFSW+3g7lRA
OlEi/6Q0bFZuRI55GQxi5nZlrqwFAuxSoXCVDJssqtavLgy3WY66RmoaQBdFfqWO32JBLbsvFPHI
I2yiPqWE59oQATuNFIfRT6r73rDl/dlrTUJsKZGAiaK8OUkNkVybq63DyOLC0FgAQYWFFSL1pSjz
THdHgpIFCB7TfnJuGdVh4ApiGU8aX6oSp7GfFtPD6l1sS/6PlErLU24A6pCLoRyUsGGuCToibzBd
YP+sIt92A/Wn2/a0BEpVCe/40lLLtUYBZG6TFbTUjWFQwpNG9iL4rKJ7k2MWqcALW+iKGuZQ/msT
q0v+oqSA6uuTJ7VD7AcMT6J8h7CoO5rqrAFdgX28cwrnZThTrDAdw3IF6CVJWn+TzrYEr5Xzy/jo
6LbiNiF2S3LfVXmxD+BEY6n1ArkJ9bqlgtyB9nuqL14fEYVrkdbLn64hDdYIyIM9QZCKlh7yyGWW
YBsxQxy0M4DSQaEYCS+e98EF/kT4Uxxb+ZKA9g+uQYOI6FlzJA2c9fGzdjU0wLwPc4gcPWDDlYXU
uD8ACE0U2H6xAVWAgrQVYqfJkHn6dUfBEyQGYmN8mJwONXUxdZSZJ8UuNEl67q/z9LQEarNsGrT4
hY/pQopytC04Jw+uO8+4WPK2xFgFhAXxQ7tKjsFeUbdyTbvgqVVAMFYYQqj5WrjKMSl/SPoKsQ5Z
hE8JLTswWYoF5WmTih7V0uZeDuaMlkJSWJYPmLkuk/IgQgoHMY8x/UlV8Je6R0o40GN6at4XHD2R
FuNz2YtlPdoBV7m1ceg6Ddl5Kb0BnnMllePfEuG5u6c9JIoIRUF5e4DqhX7/zR7s/Lzcys+/145N
deI+YKC6FjURhG03jH5mMPL5RTmwyUi8Yikv39sWPehuLWEyRDVnqKkVYWQ/+whh4VAiToKofm8a
kgTuqA5YiF2RvCuMGiGtBnCjLQnahyMgCbBlc4RjDHheKdnBZ6yo8oZtkTQHWlnnwLsvM1Fsqg0s
pCYf2LGik4CfaQwXmbjKRspOp1ybWswzgm9qM60WiqpsC4dbskkqrwNH2mMxBXuBGFpkJQen2jNP
8my5Ua1dNiS9mkrN+Y7lu8xiD9jV20nJKid/gIqOoXN0D0RryDPQzbTFks3hsdUSnbrGgfRdDnS1
Wu6zv028ozrcgwRq1t3BgiseMAC/usikUc7eyq4zedtZ8sPmVbdG0X8v5XpUHiJpIBc/0rhaZwc8
DJ/CQvelyraSerp1kxx5spbEquf+3iQ39+VyX6t8tBbV6YFjI+jt4g4gERKnRwoROKJ805zJXYp/
izgUrAmtGhliom73FZBSjUGhDC5ymJdbFErSW7rSktarLZicemzDJWkdUKTuYQ8YXYkWQxaJ3lp+
5v0ss7wDWixLiU/CdV/UgYX7OhKD2ENgZDxCHoSS2b0TDCaRYVOf7waplc2cG0sXuCw73ry0ZrjQ
+ymiDh20maT0iEyxw/k3OOVlYUmP6PHDrPk3+k8kXgBMgKAqeQXnDWEoO8vxu2y6fUkykKhd02sa
96xINnDrmm/bCoSfRWJkd+TJQr//jf+L+Bg0sMgZfQQeW8KxK23fzE6ZOaHQLtMeV50d4rAC4XAb
Y1HSmqpHN52N0lX1pdVRKKMbQVeNo003epenD3PmAuPzzddIX4St/zzMt40MWntQPeM4AlDHzwTd
4fjK2JRKJEirr66VRrjtbzEtL2jQuZCbKCe1WqhURJxqjHezovnIqGLNiu91c2WAOrCtvx40huMo
/B9nayOiYXwI3g1siFhdznFYrKIc7r8gmUtWaxS2Hkqt8UhXJ6LoWtBXjhNY7pbyol6oJc9MJq5s
gN+lOys1lynqvE11XUQsVStyHAWPdjwJCQM3mR2uyVP1IAa4g2y7JvMRvsGy5FCZXzNUHu1o0UVO
ehEZkvIWCRXHuT6ew5WmqoZSsYzQlJZTvyEq9kp8R0RGyo+UFbVzJDoRmi/t/H00+1Nn5d9Vh1rA
bix4mlQsaGyjq7xbeQDKd/oF+w3PIZZwF76QAGWb+MaUtiFw+AJwIp3yRnEOwehk6TB/wyRuk/vB
rNT6tEBGIczYw9ZZV/Zxfj+szkfw2eP9zupJ/6U+zWR+LMAZ68+f+Cp2U9JuFKhfD+WCg+WCB3Vl
KNEY/0MIfsT44RoGQ97tLKiLMFrKLrMuiQr+P2YwCbx/GY6ExnvK/20S+zzP843af+BeHyAujxgL
tkMIYVpOra0ihUfLQSDvRqf9sqMgJSXLTFdFcdEI6yeO/RQuY0IZYgBevvsKXDJPL9R4CkSJYzyV
cvylp7yWoOHsmCnb6E2RgOErlSqI1Ag6Ip4yPA2U6bA3FEvbmN87cWJ8R+IhhUf2zBW63J0K2K8w
S88JwwTxw9YMZHEBYaoE8fSuDUQ2XzvbisllywYnhLzbPYbviVOvykw4NEyK0wd2r7s1o76Nsem/
PpI85u7kpUL0SHoGFgF8YvfYschAugB6qjp7uh2aQNRSjoLjBeLST14mj87oIVS+ltSQWc7k/WXt
KezoHXMsY33mAwNnmSITWk3iRZ1IogDs0uIeeJJxKY95ko02GHC0/bwoo9fQALsUbTSSrz4vU/Kx
ToMtPMUFg31U6kSKW1Vj0pup3ITiHJmxFSF2tq2vo7JAa3tnHvWSmT3a4nOpzhXUk9YeqxeHPRBe
ZXHC3c+eclh+0peh5QcF1uoAnuWPr0ClqVRdlP2FkokU4ebrM/5Aiit4xL+sUIx+QonNK0y6hD9E
Dp4HPhNGt3PLoPeoap1JAjE9m5/k/QKrohcqY+I3nuF66z+3TlHzHYdeq/H1DqyeyM5XbD5SJpxr
lNTxUsmHnuex4axXLY8ew4mABT6dD3eI8oVWLI/PTDFmNmsqLpc3KWyb1okj3CpYjVfMMxfsgXUR
vsuRnDTmYuoTrsVbVYpCO/R5bMO+EtuuR9j0UvjI9ONZENs7NGezskpCD0oICVS+H0GeEs30KHFX
i5EN13Vggn3HRlomchXQj3pK3GJOW9o5k0WHM9w6y/t7Xvcg5F6Hu02e1FWXqx1OBSiJmiKG3p3N
cRtOxms0oWB6UxN7rOIGNrMP50mQGHqRHGyIFkNRU+2hP5XGdpMvXh2RbPeJPhRTBgoIrtRh5UHv
7JbTOmLl+lrsnvyN5/7y/ryCEyJHEfFdGZmo96/pIRlnPb1icKcuJMw6iGmkL5wfCRaLC8W7mSHq
9SyBcC0SFEGYnJbxlhsjBpMBrNGWF+sn034bWgRJHvnKeqhBA7Lz/0iMqyuA/9ETAI0QGPs64CES
ku/fgyESTCOY1R8ucfzqdNwP3DrYCk5giuq9eSoGFBLAESUFumRY25P7S6Fp4o2KRbwjxK05fUtk
5ZqZx5hkQ7jN0P6hCajx5wp89A1HcMxBZDRkVvTwQeEcpEYvcc17ohthK02yMtIY+RWXjbIWtqwJ
We0MhA5st6FuI12v21ZGRNH7P9E+u4zUrnMCr1biwRkNTIGvxGmx8A/sZl+/WjbPJB+ndRGEGpuH
USaEwETJ6P4WbtuQ6CFMkhB/npDLb6fzotNNE8DD+g5xHxZ/05PiU+cTEH8g+Q+bMjIXGXoB/ewO
Iyin6HPzsoku3GAXOw2SCGKB+y7UoVT5PvJVx5FaTot0RFG4ZxWsQxc/bGurittqvSkq7/LbQzGZ
3h2a+5s87s+uZWGS5JBLSMU/H+Idmtd1zGKMkepPX+QL8UnRdx4oImO2cVAl50w0Vhg3vnQIwX8V
HwupH+czDgPy2GDYLDhz9+gu9VSPP9AMDmlXFRNLp0Ld8VyEG+VgOAOQG6vd394htYFDeBrdcAdP
8HFKmQEPyEz776FjTTRhl+sm/gp+pEMCrcdqg9i6i1co1tVpzQKLcKAudsdfw6zFmXInFok+pUqT
GSDnSlNzLVAi/nIoFQpCOkgBp3lMbvtj8QXkZlbJdD8859g/BHcOzYywVKE/Kwvp2n95LHejaABK
WOlN88IBIgHZQ0RSCRp+F2nrcNpC6OrWfbxXO+v2kjNySHpcLLG3R4ff4BOSmQKROZfhhT7SzC2M
mqOJn7rTaxFqSx1bjh2GlrBSmFuU9DX2ipCIWDogemxbsn3VzQx9/oWT4mpI4AxNJTcRzdVIsDtg
EQrc3u7pB1/P4or/+c5AezCgiGtzU1e3F+BckrDTg27Cl02jKp6nNEeL4bKaSFBESROn/o8SA9zQ
CZ69oL87AeLATvXNNLa4Nv4SiEr7wHQSXolT2einsKZ+Jiqm7LyR2ambn9XOeVSy+lRsVkX/DD7X
bqm57wrEVLOmO5068Jbw/c093qzgwt80uifY2q5ofq2xTrNynFgZUdTi6qNu6kQ1ZW3p7tX/V1AS
5k/fbgYbKxqaCf8sxJe8jUuYG3tbMD8DL/jPczYJWQmWnrGyLQncVrLsxyVRcyhuXjQJpmo5BrDL
CgGPNSebUzLeotC1Y7/BE/aRvw2GGCSMg2KPFLFuEgQB9MhZ8ipSFfWnCFHxJTBjcSwsaFds4JxX
0OucIANX7tKP8aEe/WRcJ2mZMy3sOVKU3YkA2k5dmhyd3krkukGeLxEKi5r6AKelE+BtZ4e8aUwV
YzvXug/dq+ySHSUNtpqdPAzWIAyg9zWni/E8XZ6K+0eS6XoSGrlsH/8xDA73cTr9x9sKLI5pWuaq
4uX5W37xB1aLNSDuPjydY4g3QdqKDYMyuAohjb8pP83ANQfeNGWTLBPiNpGL0O9SK2RnoRnlKD1A
98Xzh9GKEv2pRqJO/zEqzNHdAlMNsRUiu+QfCHvTQdNu+BMwc/qxn0b2pkKa8/xdds6myC/CBmFI
OUTq6KcK1Jrrh64+/fafQC0T6mdYhsa7R518B/z6iW0DK1PO88hEOmQyhelkHYK2BqiJ+HB0SM7n
u2F2ctHcdWf4ATDoRfPc+0fDTse047Bnml34lS1J9iWkJUIvjpz0aeua1kdOwyCpu4ERURm3K5zk
uS41E7xs5NQ43VHqXZz9/+1Ypl6S2Bh2D2T02uJFMT9ZRF81xDYrt4MiAOXioIGPB5f3I34CdjOo
3YlTYyHStTOLQt7A0nSwkncOg67E1cNBGlmz+c3DPwI1h9iY8FrmOeM/2Srk99k5z6qKJdnFevF0
lizxR3efIB8PSsUvg3xPxp78oXFiPskgM6lyEL48AmwtZIP3SqNi6IqIM7orD9VzfI/16vY4aOZN
v4C8kT/1dwSGU+KPrQdN+1wXmy1gWxxKHtnz8Lrh6xu6+mmUMp/xCTatBLr8/NrPCGQ5jv9NCKOz
rNZG6M05NDvBX63+qPkT82u2YmoitUEviQvjAm7FsTG0gw6aN93XQ6LdogZO8nnDTApJD50gwb5i
2WzTsFe9laVliTdWR2iWZOdMpuH+NHH/21+OieHxTwm3BIZV7wvXEggVwnvbSYBn9qA0Q6x9nsF2
kqZqoE9ChTZ9bHNn/ck1mR/6dksmomfjEIhv6+ZaMzNFdfKuwO4llAPPHq672HdR2oTq41Yrtw0n
5hui5Cg1c1r95e1Kth+q20cBlhOOXETIXOE/fqZo43IyNQdJ7/ptXBVS1QzyOl5HMpdSNjYOqBKX
LEnDhKFXDY0h72SRVbjr8/MMz6r/UkbwdLoP1Fg/AShxgpAOKuSFJ1vUJlUg9Hxjl6Kmxy0S/7Hl
cjDVKfByT1f2cZpEWvSQ9eh5XoHN6oQgaCMPNKPRHxc32kc7qXnwIksBw6qfGi1LvsM2YCgb8WI7
kc8WWvN7D89ErNPtP4IWROHPAa2orlusatmkJy0g10GWtK/3KQSYHhQcw8Z8rDQLR0tcmZCjMl+T
0mlYs13KyrFt7jFL3KkYtA7A06uWGStGWgqrkYdLfZdB76MPgK0LRq6QtFlqLQkLUgUDGP0Q6LVA
pvK7wSgsV5A77MlwSea2aWUC7T3gnISAECDJh01MPWeRcMt/aerXNiqgbUfij4Z1IxK7tmvSo3Vq
ceta+6hdHnaPU0XPTY+D3vB/IcYoFFrtEYZNtgubkYKs/vWSZ7zkXaWwR9Nj65Ws7xOr/6+ELP0z
QBBuotnQuYbXYjln3npo1ISQpBQQBQDhsLfSgdFmgpDQPBvuLDcJzeKIiWpa09WPG/Y0r3JHUHsN
CXeOEGMil/oGXVZNV+7x8aGXIXsXkQSUw5r/b5h710q/MvzrNkdzoOQWl4kum6B85gFZG/sSvUus
Q6ihuAeY1KD3pXrHWCG9JLqozhXYaYpHI/wNtY69jT5OPreeDh5NGM7IewMNM8QXzk/fH9bfur4S
SH7NHnXq8rD4Yyicy6CO9NtvNpzfLDiNB7ggY6suRclgpNywkrFWC82+sDMwYT6P6KkbpuuUyw0l
pCwuvkUZB59OiOC1XlkVvZv3sBoV/UmJTBUlaxPis69PEOPcu9zY8SsNMYktSiRygiwTMxQ5oIVt
sfym7pZvA1kgsu/bvCsGqmDC4kxOLsmgLgdZzUVJEnMy/91BGbP7RPEYruQWM0QRs+rE9jCAdSpQ
qKGjq3u66aUk8y1P58HIJIOWLp9WcWDzWAyCEUJ45I9bNu84lboQ0B90m0O9BpyRZqXl6xnc/io1
6D7q3X594uOPNf9UNy2mOfE2xWn2pYlWau12fTnTL77dzDc/eQJM92SYarvBNlRDef1TGONIIBxG
vqrEZBuRN4VMzY5DnzjBSfJ36SooWPTjiIo5A7NAAKlCHIOIhobc+odsP9tGiGx7sPO3SC0r37Mn
qqxakjDuHT7FLMU8HGLcEPOGxYiqK/BnTFU/WXpCCE8E15I9L+y+dzz1fKMLLPqyxMvDxn1VR/hl
Rnns4Av+h0+c+IRtt9oFRQemxUzH25eY2o0nEW9fyU5DiZoCeDHW86c/iBewiCSCocLEWY5PEGPJ
LUrB6HxUQQZG+lBRuNBjj60T8mC7ETS5Cj/ZuZ5R/1fsyc3otRGCGYx9jsl7fjTOFUh5iiqdqDhM
gNFxv98Xficg0rZkvt3O5GrKKRGmQtZrt2IYa482TO27lNsn8w3AfY5MonGY2JC//fOqV5eLtoAF
sldZtDYmJASJcKaC1DvJsGXMswKz1WBG8MScW7atyPDTixjCH28w+FZSBnNrOYe7gpHA1vTM+n25
wZqeOEzjPsygnV9mYyxgDGlFXeczuha9OomsY5W1oIIfhcUAWR5ciFDEDsjocBHQuZPqY/NaFmLa
oFzSLa8X5ioW6oCWa5KckxHUCPIMTrV/CWngjn/3Qmgej9os/ksAZ2zV/29L4LEe0gj9Frz8cDP/
Lqb9fdjugmbzMfVmsgL0ZeV00PgldJi6W//VvoK7n8UxwIwdICLaWM/qyBAo3KKCJ6C8/MNde9gV
VY1l2B+KkipstcRyJROcIJvmZUwGU2oBIUXOt5zMYimDFgq5kJxKLo5hRQ==
`pragma protect end_protected
