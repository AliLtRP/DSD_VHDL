// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dT/T2aAm2qVwDcVj5skenf3qr06RbsyuuOT7dWlqfmZ0EjtqFKySKKaAaNZ5VpXr
MAwArvBK0Rjmc4UqefsSvRUkZElsKCfGGW2Ii+HJvh/T0sA4FsP78iTlq5DnfgWU
qmaWqgG8L+D/A5brwX4f+YY+ncpuhGU1aRpNDytWCVQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16560)
aY18+jikitb3hkOE783CL8RJJfZJL2ZGpaWUbTaAMgA0mQjig0h+stG531y1p09n
u0boy1qTTMG6U1sGYZ9bpbDeb9DoFH0T3aKLUpug/vTKZ3O/dphy3rmhXrxCbseW
jjYktmU63w3pWkB72aryP2tu/IH46H+em9KJ8jvjrcc6PSoqc0gq4ukxpiQRGfgO
Vnv481QjY6XTyLV27KQzo8Il1TI6sr+H9aajturLCNaCN5WcY+Hk7btPTC/d+Tb1
pvuMeTcfudtKneH3PbWwF5IrPJ4kfz7GOsn4vgGa4CFl862lafQ5FB82etCWzHdY
Euovr6QSrJ+ShKh0kUNGp+yxdzl6xUOPO5OONYufBg+A3DLsWRnsA5vtDvHWiJJw
mdEFvPx36CK9LnTi1cGp7k3lyTDyETfDSZb8MkN5txs+epDhw+zQbw0s0LIYHf/j
zUxkAqfN5djQp3r0XmVzmZ4OAnUXX+BOx4guqBqwFCOrFMH//UGxmXxi/S8UhCSw
nDcasIjV2X0womfrwsufsutBxV0sbNXEbiId6KUo4uXpaoT3TS0Q1udRAMcdG8GV
3i4ykDwiM+sCFV8VuYll+SDr1X8llbYtef5mZwhFb0AC0elJdiEhNbKL361T0Drm
98kdCZ3Irej1W4aCXgqRYzfgpgOfSSEHBR3BHcwfwVqh/nNZY+gY0cdqytVNOOXE
oQMkt5KkW+xkvfRvq8andjcOE62Z9jtTsHmIf6hi0H0wgz4oCeDlEWPU7kK5M1Gu
+F2lIO9ZvYpOHJrTmYm8voHXInqouRIP2beMRv6bUbC6GNXSVbq9sxHsY7VGOjFx
o3/8cntioSfmUBlzZjyvR+MEs/5zAZrLAvEeKxIqK5RZnQa6zHp6OhTzhPbfeDsv
qIBHB5Xle2tKXreAGmAv6CLDl8w3WsQW71HZU1XzJGO/Aq98Of1jC5DCdjTiRh3j
O9k+gxYdxaBwyFCv6vO7xoqiAK5ybQwrEwZTy6UVOZH1hi+sugYfytVl6wYWOQkd
ZOq4jwOx4iLIZIR1AIYcsBg+RTkKC8RzkDJNpsx8WOYcAbkneGw3KjYXPw3YiNEA
RVyHjtQ4mzyo/PYsYdOqG1ZCjglrSkWtpKey9p0jGKCkjJZUVRIlrDdhsPM9a0bB
8BXwQioktAz4Urm8zhyGjtoamRu6jj6QvDHnFsGnIcaGEbaUuUdfkC/dUHauw9bD
R7MOKM1FXRAazBHL9oINtHXoD1GyCOOyeLNjjPiFNLotjD0QAmELtax3WzUpTxzC
XOit5PFCPhRZmuJx7fU5tUsODucBjXk4s0ykrBvk7dZUPFpmVpFN4dPVZ7kP9ymJ
2uEFrHsjvmDmepGy6N0JSdXErgX2x83X45S4Oukkq578hzr/E3Hm0SsZlQgQ0Pdd
n0nMs66LVNIvCVPqs8L4RPIRhZLykCoh7SFrL+zvDBAMMyxLfwv+lFmwMN2PE16O
ZWgogcFxXKJaHNsgDjFDLK44Vev4vnzBNC4ziOo1pl0XcsGu9RZkR/fTl2S37Eu+
sZJjw5hYZiuM6pDHw3VZRuoBk3jjAMF6qvSlMeO40DH2dBxq07tINOZ3SPjHCz9z
5awNOj7U0l7LAHf/LIg5bzqcKyUPQ1RPObzMjdeVCTEBoPGrlWUfdu+Ji+L8AlE3
KSUBUiYOBDwL0bqQYWkO6qy2AFKlIwvWUG7MvSRumuhJPfQ3hpfOTzBUjKiF42Te
ixwgY/MFkQtU7i61MOHCG0Eu00olhSN3sB5Tm5aQmpEEc7g7CSpA1W6LJpHgOAtD
IJhdJjac/De35NoY+1rEn6rHs7Kn4oRTA2UoT378rKnGVyO7zO+X43HerV5mDcBk
JzuN0eUGjpBzPJwynHx/F4UfnP9eTSlOntutjc9anSWJSXVOadLzaxCEwZT8KnzQ
pbtg7RLvft4r1mfRh+jV03aAzZwHW401ZlUJ5bUJGv/i9mLsPwVI8uZJd9YBc9GO
vxnpuhrAbN68Suz/WtskwZqX5gVJrXs6/McqloouP9FjaL7/l5JRnq/fDhdRlDxR
RnGmf37vz/dVhQCJnyvTQH3bAi9Ns863igniq2Papw9jZvYp0bEmDSHpwyXZE97+
Y1WX5utPhEH86EVxNS7lXwJRr6oUFe0OjMJsoOu9CFy/m1dLwKWvwC0MInGGOp2r
NMsHlYGuQ4wiOQhpgc5BbeqK16hoVTy3969GfvLAaV4It+Ly1IuWulEMAFbTVaNs
5MiVoQwbLYKd4DpQuGfQ9xMMn6Pqut2MOeONs9PoaqEykCXFkQwlikj5WuYzQLz6
KBp/h1jidSFEcgA/wh/4Jg2I3w9pkdE/VrxyJJM8mUuExmS6Z6ujE1VOmjL9lb/P
w0NafUS3o3+3b1mK0jhsndtDE8DpL4QTuEigbZtxykTRMvt2hTDd4n7sduJQ4Rqj
X0G03kCZ8PYU6NLhGdDlLorPmYWt3uCWzhoxLsepMmCRhCMfHs3tqsuohw76hqXM
FFp9OJtbVbRiLVFzqZlqiNRXf9NG9HUhDw1z2a79asG6UPQza4G3/9RiUlPkjBsJ
s+Q0Wi8+RN2SHBc1gFi80TbTdRklIlLguT0AcDg4iXdeFoWVHlyFyMJZzpKjSWLF
axo4TdvbGo8ldoYWe7qJGrER4NoEJeYBKLY5WaWksThE5uT2nK3zxG54XNBj0hyL
TlOa9tNk/aAlvfXnF1s3TY++QReIMJkBCJezxTiBvxxTC2WpaPDOn8F0gBwbQFZg
vCR4PKJL5fYWpuPI70RlUXf9nRrXBlcvBjY7O0tbfbfFB1CUOJbPlIELJ5sc4H6+
Y9N3IcHNqy3mf9ho6AtiRpD6zGu1S/SU3SN/v3E9kEEP4Z+qU93oYt63hUDACuHG
nQSeFibb/eVk/77uxY0VnFEvDeO0xwItoLKUGMsAjQ9G/Ky7N77UhdEonKC4u6gq
Pejh6vFiAC17MM2BaqkZ87PUHZJ9kGKo0zgmx9lvHDSWji725v9E5UBukZ+tgxcj
rPkytHLkgxf71IhmOc1Ai/Z0Hbumtre/n6E9WoK+Zm32WDBozMZftR2HB+l6aUKu
nr7tFg8otuGhhkDhjYKWpJI23aaqQoxoJShZ4/ZWYk5BLTWgXmexgfSn06B+oPCL
iBfhleY4iHmpou7zg4plvV5pvWFuq0NSlw0R9R7sL2/uGxE4GgspJQSOIawrAVtQ
V8XkO1wmnUnQZldHq0c4oPysViCT2yaFsI2pdVkMt3GWAf5n0b6vGuGSwVXNn68A
e7mohfjiP3RfTtVLXmqitK1l1pjnqSMKM6KfSx9iGbbjrkE9pOBEZx5mlWr1oySS
rCf23NmlP5HuLpI/MuswmbqaUE+9Ip7MJTWGtGS5LHVvXrE3kUGkjZ5JaQXwqqj/
CvqXNfYyQ7MctzctY3fkGw3KDWXPWiBMhlZ+vxtTZRrYl/+ebACUECDaIlmQdvF+
rTuQ6vj1hsdH8RTRcNjEaRB/9qUBxaRJm8Rmd0EIwxEtq0x/DpMdQpwkYhIJMcjc
lS47/q2r+VAwQDn5oBzgeIRDabyNNB+iCs0F4WfvGrb6EQjtEV8pNV317cVId+d8
hRcPIvnFJEcPigCjX+L9z7GcTeFZR47WtQz13vP/8YAmVTzVYJmjpClup3Y8QRcd
CbNzN3fLfjfwd5YE3q//0NfU21aAiyAxuzDOHXSlzPZMmDHlcEZubanQxVlDCCJp
Y827EC/xGq003nbbkORy3vp+NzPYJGcWz/meAfmjLGFvsqBokmgMVj5Wmg7mSoff
V18KR5kGUUj69dQc5uXac4j/8xVIp1yDYh3t5usHw0MCI6e99l0trzWUlTxjds5O
UJtA8iryTxplAKU3335h3JbNRcNkXWl/vLJy2GEp8ftaxwKRbt3Ri1mAY2SaGXMt
3SjmrJDugvT1e3pfzNkwjgY+2As6r7DMYplZBt/Wigkt0g1ftWLTR0Mp3JBx7PVE
6k2mb8oYP/f765Wx+aG3YJEirGiFOp2f4rBbD3nVP9aFrZDkaPgTBaAOsYHA7LP2
nctLpgsDWNfs6iRNeg4EvqDC+8dCe5l0VB1SRAn181uA+txRCbI8QlCuRx2l1Jku
c7txFFpP5hWaoKODbB4FHW1P2mC2s8q+tjU43o5b+UOCu77NAFSudxpb6Qkyzb9j
55IPQpW7Ot5i6VhB9g+Y87E73MpmH18xuKGCzhv0USi+lOda4vMVrqNgioiy4zIT
z1t0pi9RZYpeHnZ9Ef/Dr0YR1Pg1HCPQVpKSIaKs1SBKkwWgrXiraFizbRPG6eoQ
xV+vxfFYb5zvSf0BXSgP5Tqm/1zWyAKS08jmV9NCA9OIrFaXkOmKeW+ddKbZbmrL
PTTR/YTj7ebva00CAn+h3zTmUmx/MRvva3fw0S+GtMU7chXzcEOYh2vuneZqHpFx
3OiDhHgr/HtYX6EYYKGLGuCzG3RbqItFl7W6Hwcm7c91iXfPjXNm52hxw0HEkV/D
f2G41Rc7Ry6W0tpA22cRXNXI0zaDRWicnLucENzDwYcyJYiPj6pLZlHIc/+6eTym
gUqVCiMbkfsUNElUC/uiD3fBCgjheragUmw6ZhQi/igeFXcY77LACjJaW/wBCRP0
brCPbw+/7OTTpGWzJkKInqFfTgDY7vvUGK8mMP2MMHqpnXw/PRkPchvDtloGFo0g
5/AHhxpLtAiIxhDPaLs3rmSxPR+SNKNYpdjYE+6B2JtXUFZLXee1ok7v8URu9xOz
bgdx6kuFuEcy0auoXXpVg+XMEWbfmhOSXCR8N1wbQwtTpdClQdfTHMRUmzp2awl5
FVLnV7kf2ta2H8dXQFK/364s2+yilOe/mde9p+SdRv7E+a9RK9CURzw50qb2oCev
+hTuoRlO7jSU0RUjKGn9cIAeBGHn8zV0MCI/xS5YgRraWZZj2BttIRikI9+2/Umz
xjOE8gxT9ZqEmQhVwxoHSauHmIC+CcbSMf0kj2S1VPm2CEPwxcfVzaWV2fHTLZ1s
hoTKUhzKGaJarDrpNl7ceMhoEGB+X9X1fBF+3Ex0Q6cnNjz+GApgDrCWrvJbG9/U
SHruMaIg9qNuVm+XTrxqX+46XdVIYTL1NcsbssGgC9kwQqElWoavcd5+4QNs+t9B
ruFdncqo6ysNmqH7l1PPGsWJ1IGvhMgW2DaWwjZGJVnBVKQq4FUuPaBBllKvRLR0
+TBaDO+FDf9hv54EVRc6RfHRu/FM5sQTVK54Clb/X5pMSRVCkrIjd69kQZVOan5V
8Dw2UTNcYgI8490aDFvLOX1GYRljZexBEwebnKTVqrpeDBkLaBPOLd7X2yk+OxmP
4tOoV42HKkgNGzciaAS/xXc2M//q6BfqaQc6TFRvGzk452fkF00amahvLKWl39+e
E2VgJ9hEE90TeeqFxoCp0MlMuJkik3qujLIJ0tCQkKkJBX1AXO2xjTrgZ619Q6rv
dvm+ugHPzcRSwYdq769N2+m1KPtmn21v6bKEa7jp12ehPJxe2qoZpyLa5/+CAo33
wYlFqXtzTzcKHv2VcC/5ASiaQ0WAZO2liThNREyh6/oJYBIcu3C3gckH5NLiI1mT
TMkbDbZ7FFnsxFQJMjIxidx65klI/neoMHTLmDz3g+vLl4oor1+snzXlf1fTEJSH
rYYNpZMWMlMUngBcgMb0z9dNjfw0vDwEBTHxTMKnsgxvDmiZTUVuOuGTihjmCDyA
BgEERLkGaTulPoHfEE3MI/+3ydh/hnxqQ9nD8W6KvoAOGcEsW8msLDYDIfiU5H8Z
mCMwu26t25WrGHpyoQPi4C6gCFOBKA67ZBUYpNwHHXAOPTLbIpCfoMcdNe6Ot6q1
fhvUkmb8aJd6s9A7ilgXSnIsA8EfgD207gk/ifaD8VZAJ2AjIvZxUmUwDPi3AjY9
DV1vPVP4f6ZxDyS6VN+n4G8XPFIY5Z/MqaGjzhDaxr9Zk4eR6YBFUNYVwB476wxb
zByZFnKJNPrpoKnk6lHQhdhjb22G2v48Mjn/A3T2O1lTk6divWS6V59/NMdCokgn
NvoVMslJrp4rKSQiXOE5Xul6r9k06gYGbcF0vU5BGAq14wOFEN/L22IS7Laz8pIc
lc7FljyBtmxWacKQaib5kXWoQllE5iLkn3GPCwKNbIk7/Glsr7zgK2rLWpsYhB6e
hNqc9/GVz/ADE9rkrvJRz/anWUYXXv1AJapSip+x3BA1h78y9SnmqvcJT6e49s0R
h0Bq1RxRhNjgpSO7dXIk3S3tbmwfMq3F7ajESsdJF2lFSpmCV9y5UL1qrM6WjQza
W7UTzh0eWYEmxqFikAx2BwgqEr7+0i8a5/catGDyX0iU/tM+FlKZhBizlTMOgTJv
LljrR7qB5NAcdFHFEC1EkFRHV+jKag7W9Sykne6C7PMh9yinAEC0uCQIfrq6dBMS
LLEol2xycDXPE886Esajlm67ILkfhmtBiP8gaBE/MR3r84DYQ71dbdSjy16SHnXu
PIDUv3UCHTHuO38+Uj+Fhjv97/xLsz7x63DL5Vt0OixNrsu2s4browVABhrVTBZK
Y94BhCsNG6Kcn8TQobr7RrPDscjwY3uXXj2zO7Jq8ifuMSJuUr4ixQQTqjN4oszn
hCCMwgrTp2hTRrZMc7aK2xvNtf1oaLFv7i71QH0Rn+CFFtVP76KW6xLGyXPg7eq9
lKlZrzikeDdkBCMTU6Yv2t7Qmm7qQvRnSNofG/B+wdAsv3OQQKdZ395C309Xv99O
6qey4Y2eMS7gycbHwhqs9I2CzqzfZ+seDyNkgPBAgKTn0d5nYqrBOcw2RHdQz8Dv
q8J3yYiSgihK5ThVG83w7BJvM+H4/vokV5Smf5SWb3NouaIjBs4QeqrPZXL9b/7P
I8fZig9xnivOnD+uIxeAaflmukrel4OwQkCf17u2kkCiywv7K45hYvuz6fzAYDP5
OyByqdsUtTFhfI0tiDZ2LcWV+BkWLGGB88uj06nYyqt9ZHzfvM1uo/0iseEsCwf3
Gi3L8QUXPp6b9eIdm+5/dNBb7T6KMFkB3FjEbJWs2Km1dHaXAV5wnubDdYV9YkM/
Pq0ZkyOoOXNGvK8TW7csAU47rKMfWR+4dou0pdogUCRwlSLxkEUDqarde/XI0HiW
jV8hhHuymPzxCDBjqPde3GrJjxqHOzYEcHGr8ZJOYAhT7bqtBIEHNnPr/Xy6Zy5h
ZAf0atZzlbKMocLqJ3Kv4eJO5fJqw3ba47r44XlCAu8Zth2k73Wk8Ngvw3QHnQi1
x8Ua/VJRuojE7cV3Q8UlD+bl54+wfIBaNpCC4eC8MbibGPL3uU+44OZS54Fu53FK
DmpoDnnyrrAZq/m555YK1SpSE07kmCbEciyhaC+zN27dzi1QOH5tD05VDgOUN9tl
2Qh75RUVRlxmzkwM+UT+Ba1Fvzhi+YwzyKgs3DOqp95y/0m/c6Fiwh47Q/Ablxmz
uDhPVmVpy77ikCAuEKdrRsOcjkR92Kqx1m6b2uLpahLMoigdFN7Y8ebVfv03gEsk
OyQTQoyPlir1HF+d/2djP1JN5peBBAYWc7XqcgMw9Nh+A2Pd2ObHdCSTDPQgwsVQ
8giGD0pn4IKIvGO9LsLaphgMkhLwI3kfM4Ue2w0o7D9HUg4XXzdVrg91YQY1nIfk
IWtmIIg9W/NQzgmsNvYmOkeQz44OXl1JbsxGPM00NKPe6cM9ULGj0qGkSjph9+zp
9GHNCzimyyYsmZyGd9uSwtf97AFMz8N59tVuPxcjYrtdZgP3AzfZrHoI/QuZTfPr
Zjkdy21zi2TkLdisrWCY2oEhmyBH/fJPC1iYky4AJImWxURztcSMYAhI5vDRJSBv
9efDJ5zcl2B+cUJ7F8hSObngqXH2p6gJ0c0jt55wAZjOEg6w9YfnE6e2PTJAw5ZZ
mh1LcTslK4CFBpwbNXSdiWMeHIODSv5Vm8HMiH7y+EoDDZR9aSIuyRoiJPkar6N4
3Zm+WvO0ZQSWBm82L7E/Wb5TOED6Z13rsRFrirjSzCUMzb/w5Bw2sneHHj2blORS
gQXD6xwUS3M4r2iyjHMALAeP69fVMl30xcjZXc6RbQv1WkL+iVXQtX26Hq9Gnew4
68cPE3qwnooZ2ba41ehQx2OPneSP05tTtkCNUAT+FQKE4PNGxmmZ4Vl5fX8vKuwV
vtj8Hd7ux4sOOIG3+rnYfYXdnbN83z+RHL3yHb+MeJLevaRYhP64Y4d3s5xkkwXP
/aszIVL7C/78DXNfVPN+3+mttiXTxxASzrdkbuKtVFUZgrEqO8LLIA2KigzGbQqy
GKhwk9vamAsetVkKjkO5dS7i0S2WginSFOffDU/BmcHD+JH8xWg3H3AHzZ6FtLPU
bAap6glHVWhdgpETBR2cVUVu8vJrzi6/hiXLBEXTBJr34t6/n1D1HdxEmoioNOg4
na7+9Qu24HJgItjdn7HyPnJf9cKUAaY4dIpcNnh2UG6nTKryaZ031v1t1KZtWFkX
NQVP1jaZbZ6CQldFtJn5ENxtjPo+mELibSD7hbmPqJWFo8LGmthAU4UWT8g8kOAy
d+Xh2XVmp/eqCZZdD+YVuKgzzOKCFN+fyUXHU6FshkIl2FI71AtcaAjCUZDuqQz9
3amko4fHpoL5ZtPaMrHW1tCfu14x37mTT4RJYETcUmlYMYoqd3+lRICKz3aOFV+T
9cQHYR8DJQX2PxGasS1dWAtj0gnQaLbuxVCV2RnW/A3soE1AvpFpcQV+teNRj3ot
QvPGnqhAVxaHWCG7NglV9uRJDXw1H/IanhXiFdno2LNPJglOSPzzLKKHUCdoQmWW
0bfj/6H5Ak/wu3lkgRs1xy/GPFzVkg4/yaZFv123ij8wQXyy4s3uiyyIN0sJsuzq
urMrrkV8e8Ld8ae2+Rx6d9RJ4+wSpRMSwa+wTPOLs2KBwQS7tABfmDf3QvIOjtHo
KsdbUu0SIC9sULSBvOyKXD/sEMhs6a0yuKP2cCU/PZ9C5LA7GMtnAF4bitL4RApX
tuz/LmCaanbv3L9w62mC1SfdgVd5xfvHsywP4sAGljx1rd8h8k/7DZLiDuW7xgbE
+EEJnAqmQc5PZ5AiBv2Dzv1Ad1hUVIYezD3xvW7vv9NF7LH0Fgyi2n9Mx2/1SyDP
KiUEmvanfuX4+GMaDvlCITgX/Utpozs3fF8MOBQ5f+6YnY1EuuLp0ZIZZvxzXDgS
n07UG+6lAyhTdRECbSIRAhp8kzda1EQR8Y4P2emuBkOOFHRvbuU0TMQtMHWYUQ2o
us68wBgYS/B3ioisHAsz6IJF/ui0EFpOlTsfuyBZK57aAb3YDoLw5S+VEIidojwp
RYTsLP2qcYB3a1NqlqPVrBwQqb9TEa0pqzpsRwaQHUMMQuziEyEmp0w/c695+Jmh
9AFdoFG7MLi73jahQfMGJ5cBOAJoCswNaPpOQBTuoWmAySPz1y/1YYBU3WyNtiR4
ATfHxwfbhqZ0777IEk2m3AV7moG8Vpi+mZuNaN0lNLR+0WKflPOfTrdHIvZS6dex
TNIECcQtSfV3UcaCLUAie+nB8YufEbLbTwto/Jk0j+noxHdiTn151YJhNtKYUWoE
F0Yhj+FtKckcIG+mo6jOD9Eo9H/Nvs8OtRNsd2AEa3IMY//0Lgf0PR+idLEkFtjC
vXjkRO+/AC2cCQjAfsxduwqSNYMVkETfo9q71m1sambw722YYMeLZtI/9z0oqxUR
rFY1x+1yKQDsa3H2SXoR8fupTQ9igkrh+HaeuzSbs6t8t/8g0WEJNICERjOSEvHQ
hKMEOu8/wLTKG8Buk9+mA6TgZQZ8I2Yu2TE8nINAozYWwvKJTJOPXaBHH08wcft2
t0BzQM+pYzBXIV7JkEcLpSedo7A+1kElSTxfrmVmjFlI70uW37hjieP7yPjH5v8c
0xnteGeXUEr7g4b12uO6xk0S2IZHe2pjEVUbYHiDVemjjK0LZBg7l7cJkTgT4Mw7
NdSKtB/8mLK6xKLHgu+jkmGNuvf5z7UUSeEBUsaomBVgIBEXsYKraFaGCQnzGb79
nY4zMlTm358EZ9rluOLzYgrRfOJt5Q9WjFyht4/1HDyORtKbC6jUBeYWhBKKYcXa
TxftS69UrwEr9DScoODx10+9DQnbmh0huIHjGSpouw0drJ7CsOz+Eg57nc0bmF9A
PWdJIIhIxmcktAOg7IkWCENp6pcd9071O6bQO3uObz2ypjIQjCC1qG+45PiYDfp/
beQq0OHhfvjsL5O4YQ3ncovgJ9uIWVUxEZrNhjlLvpXH17pKIGgY09jqZrCPi2I9
an+QtIyYAzjGVMAazhqxnMWIFMlwNWtXvvo+G34aHh4uhn50Nd+G0CzUKOT4rS/2
in5KfJ2GNePFSjH6fWIjZzgPrWEl0axwedua1pfANIHitqw8GmZ0y+ndKfI2qgci
usfBKwCPUeimcvgP1iXR0lt3zXGTYvzQLMRqR3MNTQAG2/urFJHGnMjr+d4+aspc
kU1sXaRLSPAZClBELHoEeedQIAl1DTSrVJpqGcMhBY/aRZd4+W27y+ADrcPYqSHM
MvWkO+R3B9QgmHY/uQeq/bXP0e67KjatOOa8vN1plasFQNQxoMx8pDbzOQgWmJfH
mlOuo9tdBTPKuad95FWDid78N+bKvr7W08/6G3Il46Gkl7nXuxkvKWg7u7beVszx
GaXKWl0NzoKqj1RHvTSq8AqtfgnHPiz4aFcHdNG8/92kM8lxpIHPsLltx5yxxNhg
eei7g754GmSZl5CXJhIjrP9wlBxLiV7ZzWhsgg7aeNgotZyCs2l4GW6NlHJsHWkK
YuYbyidDXSggcT53vgXhEYILdc0W5v3vK5TQyyS2iToaryJNzk9LlH0LL783y9kP
KnKDdExFiZJZFKLffVq49iYu5KEOtJH2eZitxaaGYD0t2/xXus6XlCLf3iW19qwX
oYLeo/Kl1z3yklE7SQm3tApiZk5z7TELnlXUeN3w1LkaMHgVgPh92rgoi972p5fu
60vuq+dHnLttGwXJRmrxYFJw4956UhoQgrIN3TJfvNXkGpS8d+m0s8c2JtQpvRAU
F/nMT4EsCjxKf3DgweyDWPwMehPFmbtb5a9mGqzMHQ8E/StwKalC522U8UbVh467
ye/HewjQTjvAf20U/OaYkjcYHSW0/Wu1w7OyI+6nA9batUxU8yv7jntpL2yb7p9t
Cf/bsEgf72MjhztPsDC2YmTB9o2G08o+kB+lmqTKeFN68XB2BzkhWa2udcKwffBV
GHXANMVHg6O+3cx8JASNwWNbdUOuXbZBk8PB/x7ulhGA5EKB2WAp40F/thS0j9li
Vx8FwCVU2JG6YMaY4T6QHdP5IPM4ogoDv9bVvaZUwnuyTTgqjhhKAr9t/qMq3s+9
zpVWUU5uIdJpz4bOmhqO+CrkkmfdzEDo5eOF6Q9gXJ4F4GpopIv9shXZRYnrQEXB
OgA2efC9SH0oROUADfDPLZRF1Z4Q9i7mRy2krvHOgtrNXJ868/fvT1GP35w85lLP
QhsFpLEOrUP3P3hPy73UyHEFEDW86jt+FONSSbxFK8AytenTxUCaMowfVXF73BE2
JHkZLjb9Hd1hjd8mLbFyGYsApDmj8mF8MfdS76AvmKTo2ybVsR4DkAYn0rx6jaZV
5eTKEJFdTIHfoTpnPHARY/+N40OJNxMPNljqEsnRTdwiC07C1wGzvcseyfOEKyln
c0cInOSJ56cWRUo7ZgsQ7Q8afMOTturFwCxRLNwLwvrpUXUBWC+esIvY17Ys9SX2
Nec+m5V9fyPe4lxWfGIOSeNl9Q6F5cTLvTXcyu2XwzkUWfe7F02FGc4WiBU/Y/Um
/Z4me7iXwcfXsVqP6XqBXweVVKWz6zUinJutocjGpAjP/pm8zCBw9J25cvxHChuF
jax9E4xwAfLScvfsugv+XgaoapA196JYPKTix/Q1ugRN4YTMUPfHXnUkQuYp6fF/
smmXLuMgn2CACKsq2hRPU33bxfbj+F6gzDC8Uby7+PsmvBpUilMOifOSL5OTb9X/
lsy40MEC9WU9L+oOgY4z9jzGXNlT/fzG1sBFA2IOq5Hevhd2Wq5c2zVMYqB/e60T
W6TkPHkMQeAb0BR7ucltEXd3tvWJEGeSK+RGhS6oI1YQNGR33PfAtqZ8q5hfzOlF
LY+xpW195A6VU0nX+3ZtlhFJCdcXOj87nGZZOvuegfHejEJYMnaQAilI+wK8SYt9
3dyQvIgXGG12o7K8Wzs4ydBhZSIzn+o3C292wozX+PtqvWbnQiqcuYy47n6ru3CH
pi//bAgUq9GlhyBApZgR/HCodDeVr5901wpgGewTafzTGdWifVmkNCBRxRbk2aFw
1X6GibuyG5lRoM2J+AGfVOevRzRRRh17XZXqkQeLZkEF+GOcEuzaCLHAF3yyY8S/
z3sjUSiN8/NI2mbkkvjhdPcQNi1HXaR9diHvm/KRvz8k5c7DQlzULv33oJixUaLO
K205M195D6hYW3mCe3CzP3ySH+jgz68ASlGOy7vFkEUbR0pseMscTRHWgeqg2hUO
mIqxSoxDCPDrqN3VhY49j2Gk0pz2dJPY/rnIuERerlNiJxkzFxrDHenV1kKIVxZ+
1n++8ukuN0+YKt+Al5alvnLD/OEiMMbWWA7HHub6kyRpI5a2RvY2L/yeajeJplC5
fThcb66ZeX16va2zzneoxssSMufviZ6tGRCwiiw+yoKTyzFEHoPShVCU/Djr3MYi
W6cQERt1h9CaV+x+t3DJ2sDvbtpivsFE6SJYMOGPJCvs1LvJfRUo4SN0SJwW2t06
W2W8gGYuqMwEqZp8/IzWjpgEDJTdRatg5tOc/Y1C14FYDpOnagbTqW+VTKQ4S5JY
6ZS18AKNALjjQ/q7HA8gs4KWU4f3kc6kaZATEzFsvbdF/2Zi9E5MJHkN//D6pac7
q4+fv2Eipd+j4993XoShdXTchxyXe2IVfzCCrZ+1R/jk/KB/sYltMD7EivJquEsP
tCcNY7uYeDAxVc0rrMkmSsJLfSDcjqqi4NSfvJUZ+w9GEwM5AirEP/jQeJV+2xap
VFFnBwAIwhiNqHHtISf5yFwJ2OPniVSqWUl3CFAG01uKqFNxIfGXL6jrQNVBAFMf
p21H2DXv7nFAwx3FIW47lk0cgJZ8lH6a4RyMOI8jfSjTTJgx9sN4TAjN5WTZHYb1
es4u7E2n5c4Hvi6QcIMaPgJkAooknUqTHI+2veVjf1VToB4dCsxl0hLQLXmNrZE1
ZKFge4RJ3qMBoNTE1Gp7ZApxjpYL6VrnG4OitySHLsAqwcjwGAtzLEh0U3png43o
43bbBDL9FMn1gGCs2VlIWe+NdG9tZxYTKk4aONDGyFRnT0uTVX1aEEvinrrILMRY
L0Fl0CMg3MK+OcypZSYQndGaxdk9BK4glRNEWSZmiCx0JnavRlNo7mc5DJeGyJ5Y
xBjAhbmGofWVPiyx+Pe1aBO0jA+UTXcrasLXdyVTU9UDfsjnvSJJh7FnYW452x9s
RUkn8IURx52DRQL1hk8sE2YbpbZpQkxLglqWwA4VKWzoYnFOwJJKI3XJeIV+4HrH
5aOi6284K38tMFW2r//FREp1pvDyystJXpFM464HQAQizBJOhgzLv2pqltMxXnt1
73XmlTVAIAy0AedaXkW6enRUl1v8gp0n0WELjvVc7MpwNU3PVSD50YdPTtRNVM04
QmUGMTmPr4xX3oTnd4vk69dyz0CNEGWJkCfvc6qX7DEjZQBy4XFi98gkHEqhAyp2
29ujkxgEO+0j+R3r7up9ADTr1h67q7LQhnDbhcu/U6eyTiXu9xigH32uLcaXyg1Z
6G2VarbTfGHKO/cW7NVIRlf7bqzZ9pMyIkvAVQ2FHa0oO8hBlyT+/NQX8zlGw6OX
9WHd4yOiU/o34cyw+kRGdii3/oZ0o+8MAQHeotGBOGou4b7ZUGcld8ZRYyGudNXA
SGIgKjuQa2VNrpvXY3x2vHXZ38yKSABw4/ULaPY5jKJIGnRwt3Ui14Z4fx5fogPr
5rfhg3DGf0ITI+U/QhBsLfjz8WVj/kGi8Lag9p9mYNt386GDgL5etI1AFB9tBTA4
YgR+xArTS3O3qsYxLxhGVNJRp5ydYM0gHjaP/3KSoM8p3F3xuYsdpcpN4ttm+Ipa
smD4NaiL5a98HfDAqn8sJ6mWf+zXMzZVAG0MdRBYrveSCmAqEhgEGl8T5HcmCOmv
YwEkrgjH9ChmuVDIdCeitKq87xKLrfhmrBeWNLTCLzcE4Yx+2woOtFSaQNTZF2uO
jEKRT9/Y/zkt8MrFJytj1jgeZ3Vaf5EXj7yb1RJ25mTTtzVKi0YpJxDUPLijMxnk
05j01Aco9WL0v9zKowsR/tuuQT8oND2x1qcmoBeDiRho3DKjKQXFRN9SDMmozDaC
3jIlF7J0c6iEAs4fQsfBEUwkef2b9oMfFKx1+HTejPyyYol62wlV2TEordOl4G78
HjFdE6rD1Dg0E/9RvZLkyAjc4H/0ORo0BviFIUxZ7G/sCIA1duQnnDoPXLic2Xr7
5RMbxL8fulAQo3E7MiaMQdfjWKHhLf3/w5hREpr84bGxVmieyY/LvgwLP+TXTxve
tE8m64SdMbGNJk3LR7jI2epnAKU4AwCs/FwWdinYb/u573O9sezcjg+JOeUGTxw+
CjcEsDbQsBp7j14XlsQ50J5ee+4nVhnl8GlWhrOY25kto7vQGDTkRuZuVW+uAYXb
FA9Gd6vxLS/NRG8oCAOy2107s+PNwvqKTYpd/y23rxCLI9Tdqj3ND0C8u3tZqk5G
HOKPyYcN8JhIRfOrqS9uvqGL56QwHUkgKKJulJ2KvRLDRadM4S3q9n34xAA9U/sA
Sz/rymT6tawgq5LxBq9jRzBoImpe5UBDq7dvuFuYRPyEZsuzTZG+gU59EB+X2RnT
7Blv6TD7s6hl0H7E0Z29gWy5tBaHwj98BEJHfAhbJknhZiRh+wVngU3VlamJnt89
WalJTjp15yZwBHXfo1ArZx439Nud8+8Fk6bvNle195SSzuTj87M8HYcsaGEpwZ1E
my1K0+hdkF8dgbADIJppwJAo8gW5hS7OnC1aHHA5ZU5IhmRXmK61QxoxeaVSHotc
Pl+2x0M6wkujFIWtE36MJw4PwFyEjTSIGgW5YgIyTFgPyn1yE8bkn91YE6fgmYMu
F4cYGEjAczFoJNWx0EedE+mbvTigCc/2UH/Si7e3c9DzjJ8+uMxBX0kDdGnHsQ2f
RUI3xA7k0FcEU7g/xku+jNwjYeIOg/lHPqLw27NmOJyqkYWVrOuRJYan0NvjCYC9
ou9uCIykE9i9Ab2Q1MnMzv5yPHkcc9HMbMJldjAt9tYwaaDtx1BYmn2rslhquNbb
xjKSttuW/we6D4pDWnaV+XXQZ9ovptIdPHCok0vTS39/psBkUodtKmV3CfjmrHuq
vWBLFeHHm6c3U+w7LAq8jmuEiQrPYGRYC7uHXR9RRLFEorjVZ/mHrEIQ1O4Ktla0
7ABROWb87JpFJWZ/bryeJus5ywrkYAshAVmw6sHgU+Rbkp1Vi1jN08tJMCQq1ojo
QK9OqZMdwqoXJITZL+V8kWZtobrITsSy/OJ9v5SEF/QU9W0fVZhLDIAKtVhfm5UM
gcprebjsAKKdWjkFPT0LYni7HhA+tqzavMKr+ezjcjhFs8s2DArMCCqgOW7nO32N
75oTpR6MgXrm7OxreYwVC3f0yjW5zNk1IKAKduyEvSfu9lgZDWwxA9jkaqOBKljr
p6G/ekFIX5OlVCUeYplj+hEPWhyldiiG83qsXD9SBtUJqy+g5o5VcO98VY3LGx4u
qNnBH5r6jVx2sKOJ10SN6O9QBvK3ZTvgOSjtDu9dtPdNxZJkZ19qCi6FEXtzK/Ij
Fbo/JlxQp2frRVNpPC4NIVQf5SCSrSqdAPODodx5CXXaO/4m7o4T75RpVk1am5QN
tt6lq0WbrbBw+Dz9JHsrWuTFqpvTze6ac7AqoYIVkMduyAjOFRVp0jmz9JF+zTu+
zIs/A4FIoSCteK8eDfCLGuFwpjUBcgW99NZM7VhmYbWbWVwLfYDnu85yDRof6LGT
bfBlbRlv4k7mfh0XiI76+6zRGHXcTRlODbx/cl+YWy5RcFLx3xuJDie+JVcar7d9
PWT59gII4kWrNxJfAXXVJpiz17DaRQ3GntcVIAevMr0zJFxKaoppF+R3tVLZbBlH
5dejHUAR6AWayYwSUozBLqLJNTRLYdHL3A2zVQwxBiTS8H5Oe2U4T+O0m5MdrFch
UYwE99G7wL5xo6wdcRNZZ5NrdlkxEi7Qtsj/6OXamEZXuLr2qUEOwyxKWFNAYUNR
7OUNu4LGEOl4BtFONbYEdNz7tqWUrq07TVdp0gjUhQx1Z12sS1b9C50sm6zjEtcT
JCtXrXvCnybAo0VWFzfnONbC1CHb56idrotG5vf1PoUuw09Xm/VbkBv9Y2Hf/nBk
bXH21kvc3Iu46ZpX3dczD0RRL9cZYfNm7/OV/mBSWGO2bvyjW5XnSxbCpaFfHQvK
e3w11s+Veo4REfmzJvmzJq9t62cdlir195b6G6iUUmtyXbzl1L6/4j5S6s44Oy/Y
dAixrNH3Szb+T5gW1Anemjos5QbbnSsz+J2+tn0SxDPGn73Yiuuejos1n/3d8HV4
aMA/Ygcc1nKZJikQW05Oxutwz0S9r4l/vBU/7XFT9X7GiBWW0gOChHebA/Nikyy2
bDqNesTZsN5HDKebVrVDxqLMTzLaskko4ZN54G0YKuO1kN67lnztsHr4KPpGYr6D
xk5pS5Tg4HPnASi40e87lnhkQDvYsvInEw3rseurUikUnyDv6jEYNESdu39QRIcc
q5DozOvs6Mf75Lzl11vP0V3lQo3bVe+FOI6q4KoCqvLvdQJa7kSJfVJq5iNVa77a
InbXAH0TYOa03ehyMM3wHm7fJzly93O1GAqS3xtgspCesCZ2Igrvitdz5Ev5issy
gN7Hqva2sVoZoOp2UM8T8cIgPefV1t0AbNg2oKFCgTtA0jH3A5sQKatPAzXAqIkr
eQIWlIYTLYs1bvLsxrYKBJMJ9IP1R8TazmaxLmY/QlSohVFUi8TFYLduYMSW9DTy
UN+J8zE+6WRAhBcVypEICkk2zjXd+3aWrjtpJt9WU0obolARvjQA1KQabyxiy2TE
g7n/RAg/+tlKPqc87lB68tA1ienkvXtbU1WOPUCEuADIVAoCdn8bV7rm3rlTN6NF
qhuUgGrvuiW+53HC6dEtnktW7RhoXaaCUqz4nsLxjOICMzZbT9s3kBhTwQYPuVJw
ADx4DfgwFV7NOAAwLsily5ZgyLDuTxOq49mMYE7JGT9KocTkh5gxUrEP43HzGWoJ
zXO6IvFORXrbjAczBPUEj9q5uqmy9WRAC3VV+s3SaZMjeGe6Nv2eRngUCXRfsqTK
/QBbV2lQxoGvK+SoJQSxhqIhFqoJZEUosOoLAF0gvX61BXZRf8bx89+2C5HSYGvk
MDARxVkxUNqH/ghgdJcwvNuUXgCJX0XLcZmP/18aqkmdrMJjPY2Qo9J/omJNWkmF
qSrZMQe9Dg4O7cbZQiKStNarr0/530KNUWOGNqC8/+XPGmkSy7t7QSlv+UrCEfi3
ThvDujM/9dA5w/GF87wyz9y08eAKj9LzKBstoRvVDTDXsaAhJ6ZwOag5NBCJDcBB
4d1UgBOM34I5VHndUoMVwkIVSXbjAogD+a62kYrCUzoBsKbCJ7fmUVFsM6MbzAUk
tv2T7Lptz8JEb4Mt1R0ErBrmOjasCflwKchXUPFRlo0hP0+eJgrHUk4LxRb3v4Lz
jMwMK+hdGJC74e2RiT5rcz4uiK/1wIvIve2kfYiHAcNbhrH8toGkRHk5KchquQlH
VxuFnz3q+lpXTQ0cOt2juuPBbH2gIcNSDZ2AatLRHNJkXOPyK37DYJzjLoUQgzWJ
W9C6NeDajsnKhp+qwaY4XOESpSeRzoAHyc3UcD/Tr7OXkD8zZ0Xt3T07lEyS25oM
38y/n0zKNlIhbCeZW+o4i2MygZNwmW4ofxTc5xfUzebeuv/wPITr9JMw+EE8sppR
SgnJ+xUImWqfOz2EV8Dz5mh0XqjR4wJQmzJLGkAcnsPuej6doZ8fSUb5UaFHhBm3
QhPWQOtwmecnoaunNbD+Kk1rWttFJ84cxTfqx7OmpcIXNqRRaaLF5w9wx0s0En1d
mhpBo+/FA8vaJ97eGu/9rOUFZ5q7zTnPhwbO5pAoJfdRgAvqeSfnpI+RIoVc5vvx
KVXavQhmPPood5cRUVz4rGYhj7IlPJJjDUqEMyVd4xFAqCnIqC3mC6KP4nEmpasK
NFekN8JKcDIfaRjD217yuGNBTmKWQnPwkMe0Rw+cN2vn20BOC6YFGxH5hZNqOciC
EgV9FzrbkX8PpGReaxIvoYSoac1BwAnb7ANKmJpJCwJiFF/4l13bnBb/BC2pu1nD
dCXPzkxJSfJLJNezvuKadweJi2ehxhJl1SVRtZojZWkR2cCF2mMzYlQyH3daR6zf
XMZUfr/Egzxer+Wx+kPdCRIulFuQvsg8Mm8S43zDgjcAHikcjSLicUKXvNfm4A+K
eSUAqVQavoclZZHVPJROoO2y9ZX3tbcgQUZll6JXtgyoSjTlLkMeq+s6h8LbBp2u
WYMshtTnAZC1mE+jkGUjerODJ3Hxs5uP4bhbwlw0R24RY/hJ7eeuRbHLQqOO8VQ/
5/vv//W0GaySGouePgToYbeIy0PjlVdeQPKnoYyVJW0lkLP694eWrjIuWlPt62Sx
wXaRr1sXX6UeEmEakuGS7gOuWKIG7UP3Fd0kJ/1n43Hi208YwwrNOb83K8rVKjS+
w6iEyPzqA+ZZNZeWTfpalYnfQ7yw8MGBzykmkPjrFI3MrdzoyJ6Rr/VUWs92V7uE
eNpLtSv/rf15oEzBH7zPFwcwifSCGk0Ho88XRZ9adWaMR/KrhHjEz7PbMuyHZZ1W
Ax6VU3LWp6D81ThjVcWfuEScRL4iemGFciLSJI5yoWX7BPuSqjAykFyGWyeFt/1U
zX2dQWvs83kGC/A8O+Ef+8ixrYGNy8sDvOIf3SMshv/YnO5jukNmFpNFf0dAewaw
s+iGgrAW3ercZxJqAhe+3J+/hEu59gqAJSz2brOD5q3pOZfC74ePLOMyKZyPtCW0
WJsfrAKTGrPMxX0ua3gtKCwBHWS4g1EphVwIYjYg4KojS6GAWM1nIolR3O81wuwQ
KGz9UGLlQLxbGG/cbVhNDxUguows0fSZHVrQ58eFpLfDq9212FLmrVhYtt8ov+UF
LnHVzmMUEd6dQfC76sbJsVp/WZzWiy/w+W9IcCuw5wn9s3HNtJcbEvnJGsTdMdas
KqybXJ+UjB1lEBUcnp0i1bFZ6VuL5qZ459WYA8KlpyvF8KL3DYvRLyrP2qqsOKmI
T9OOf6n7SxSgwziTtv456ZisohCcOLw72arh6pph2sHeyuE9JNdrwllbDhYnXTSP
kVMPuQ5/Xn/XSTjSjyVjukpYfCi28K7VbliBLkDPoI9b2Dp7zbd8K++ij07CVwFW
LP7TjU2VyogvMG5Qtpj5xPSL96WodvlAsftk5IvWRdWArYxc8gglUCbV4XTq8NBT
//qF8LkBDbo/+VjXo6WxweWabbTU3JWPuxkq25jynzWDXOW1vAiUZj7qGOZ7NIAQ
2RffGZeZOs76cDftBQdRvtDwiw1cWZImrN7vlWVeoNiSNwOoQvqkiXz5FqUtCMTq
6G11Pn+w3TfIK0/sW+VYHBBKQ7q79CwhQwpDNDg9ZAckME2NKpULP12o9mC3Cpkh
RcZrmp1sxx19Vdk974LLtVtPu0luv5/jrHigok2oFDHljbV+AFxr9TpKkWeV5x57
BA+SLhkgn2yRTnHn+jopxJDw9q+U+0aQ4cpnUr1xme0HmxvxhjmtR2WI3ZghBDnI
4uCGGR4jXndHT55d2cxTw76nLBh4WVIPlAeXdikG9nn2S/pL5PMdrvXq+dV5gq6v
HnHVghyE/n7aHZc912L1+6ft4dMb1aUNixrZL4e7f1kHOtNxEje/uk7fRMixZ1AH
RVdH9OuHpLgF1yQakNQkyJwWLIv/inKZTUN2cGZaIpUwplCmYLWfHiWQ7pA6q1Xs
nXAVLj9WiAjyaPBHzRg/ZEjAy/NWVN0eDNCXwXark8+wpcCgT/oXAZ5QFOUt6PJP
yCd9tQnN0mip7jOEjEm7hgSUgNuzVFsly/lZOD8r/JolhMIJx5wJOOb333jxZKQa
Z7jnpJGJ/uoKE30p0PdgyXme1tSIobwVmFkQ86QiknJKRMSv5mxvFkSNuFiGMkJw
guzM3jR9IlKDdiOSSUlsf6EALGF+1CFSdUM54yoAaituQKbmHJcqCTC5VY13tEK2
kwPwPhBdItpGNddbWr1LhP4XHtbNIxAMATfyA0qpLwY3i52Vy9Vp+9pRYEM4MNGI
SXSK6koQeceeQFv+J58rL9OgcVRimJTkuwywFeZSNiy9hP9njq50uL3AJ97uqmtl
q831n5Ad1anboq8JhGZTts5mJO4lN6YSN64TE2+ukzAT9/p9FnFbXr2rGDEpvgXE
DeA5DtnIabSsdHQnnsl9Hx/UFhyJAFOduimI/XHE0VLDrgQ2jE+CZ7w8XfC3Qatu
FV7bFYACo5U1TVBsq0rhiNHa61mIDY63X6QY0IeWCBJIlbE4IEYpKKNa82t5TUFV
pjFx79IaC0mtZntzmU9nfTBUBO61mREgwWWDPFh0IqufYmVeL740MuaFiVegGA4C
ER3V/vkTQVbBqSi7q5wnAgeEaz+FqYL2Jb+HdkrVszezjmdItjas0CfypXu3BBLP
kpsSJv8jFZr4aodxnQRMnoDTUgnEDLGY3ZIwA/ENpmkvRbZ8Q0LdkYeVarH9Tzbf
W3YQhK40t5z36uZZn+zzWVL+fe03EJ5Q44hDcvKic4G3g1dd0gNYYGq4Qw5i6NSK
NiaDjqEqW7bkwqAmIPF5fCZWrwrRvs+A8Misx3xTLbz/b5mcVylVRdum57rg8jVB
9tERNpNjUTekLFfjWaqv2xJS4yuny81tOnYzPqZ1PWCFdunnbh9I8efwpOR8tN8n
86ycG0bGN7SlJ12j5Sy1OnU90TTCmAuqUoA6rXOMNcLAV76fRLqCxiAN4KPtvyrc
SZzM9GeBu81C0hYKv5HEN2jIBoE9VvUo1gWckVL8duL0Zbi6M8ogHqvIlvbJNr1m
mV69iqnfPS5oXpIMIMucOIyH/y+VP4a0Ynnm2lIhuALMBENWi6UNJUHuMZr87P01
WErxgtPJfJi3uNtqana0ITIV8xmP/V2iXxEIOWJ9g+/CKQQwKK/MH8ZNDu9h0ESk
O5YNcFy2/qq19EDIxoHfSoX8D4Hokwa7Wl81gPrRB9Yft4AJI9/5yfen8Ble1SXD
lmutwFqpSj5ZIsbpPVKYE093jYDIG6gcS4ix8vYJd7LzqrasWMxcCMWSBxJj8IMS
zVvMgzhRlIkBZR4Jigi9kR7U2Yb+mA/wZF8iMy6rNKMDFeDGtgtCQ4LKw0z7FCm3
EN6LNCFZlLCYFbkpsvi2tryxD/TLlHD8iH6ePI9p+fHbxojydbKfhT4Nkp8FECZw
iYdpdkuQPsWCt7PEgkAN763LGxBgBNHlqWpbcDSnoW3BJYNwK5hlxaDdghRQhNGR
Ec56w9Xh7l2aSiCvlQnxfl6He+E1+YcmIWGc/15LMhwGeteqwb21LTtuNGYpFI3F
L9TMQQkYILrSSruFZ52VYoW/HcTOtz6fT5pWxMUSm3GNaJJw3em31Tj65PWGVWi7
31z9PAZSZaJRVeatk9uupBufrs8cbOahAaE14dMsodFrs7QB7a06VGu7CDKi7XEW
fOPgZ922OiayZBaQKM0/8HsrJPB/S6EYBtS9s5AzEnKaqSgjVvmGizTpcQKH4Xn1
vvG8+8tMXm7J0vYZheamVBPij/U+roCA8SIGG2Xc2RzfHJhLHDy3kIOOZXJv65qc
QsjTlosQDWTwPRxztOP2xyKyB0sYdzGv8/T+NMfWgL2eNajWpCYfhbYlOloSz48M
gEWftPu8w2vxAfPXUDJ7KyCHsDAqiab8eE2D4oZMQHB68f/iF9tIFi7Zrwyau/S1
2T3Xdlt3yGRg84W0dASEAb4FkyUdZLYuuHF9Va0B1SFdgPt+YBQeMxVbKBH91pCe
`pragma protect end_protected
