// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
b0PVwoO2jbbfUau8sExgfb2M3Di1SbceE3t6ol6TG9LcNAVF91RbWJ/N917knh2XvMvSxy3oeTWB
GLOYO+fxtyiToRkvmPms7tdGpcK2zDvzUSZF8ulUX1RZ3NRHGt8e+bE00l+w/t7OsgcyusIFgbIi
R9Ul/BVpXmedcyaPvJF2VeqVee7ZxdfOuJnBQel1MYrKVnLnyQspZuQiNp0JfWBrF6yS3rKuPp3F
VD7BevawQa4ed2vnpXnSik33KqjshHQgNKJoAKaAefYKESSIOm6PmefpBE7q3O6yAAJ1BJzOBHQb
KM/PCs8qQw+sQCrk4wGu6P+w8i/9CL0H1kO1eA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ZVKEvOOsqlX9o/bqx6H47k1ER6zivXsZDEnW+qWVW2G3gmPsucrx7RfbEB3AxQsOlkHfo349pW30
Nt1t7pTRwHk/fYIVLom/x90ZTlVWqw+c7SxPtI0ErOpgzjSX+kje5X8HavAHsJ+CyRrA0dgiAE91
CramO5A4hXcbQnTzWzroD3UUFYomUc8hiWpaW+s8YL5m+KdIlTLutxqbW0Jkkn6HKXYY1qlQXYOR
njfRoRC9W9tBoh+CK4WSUsbnlf4FsnUD5PlwCYsFMV3E0ie+qGPC51Vz/E8D/9pgpA1s5/4OwcJX
aVDXKEXRVWVnmtiqZAtV2TdJ4SQdRBfy2N35OaCVpFEnUQvHlVW3Z+hoGFMLhXY71RiWTWFV6Apz
jpYljixVoQJIkyfXJPotjMSJNbkrwXC26X52nqJgT73mSu7udVRDJq7eIard2IeIvLAbG8mCQ3/z
COQwoONfBxxnpQjAVAN6hOeemscr8/gjST88MDUOyhqz04zRvIJiPiV/eQMnf3YyiphAyNABDnc3
ibwrFNypd8EMzUelhSu8gu3rIZdyHhRurJOkmXonn7IB8pP5Ry3AiIy83ZCQ8SwCf+kcVAUVk55j
1V6sI0BCxOgSakm0ytiwkBComxDKle9EQI5FoRlKpjdCSGWhkIEoZzSneZwNIrTTcFkWUbtkeqfU
PDri96saRArwTRrAlhzk8n+vJ+Sg5nYcO8FKokLUlcRtkzeaTWB+3RGJNiOorb/eWgSWUJC/R2DV
IyZqxdILZ1LrS5YqCYit23Q4estNoQoqErv1tyF+l8obJwNM7qfSVd9lsfZBgSRJNpMC5phMxEZ0
YFXHHD5YAgThW+E9PkYQt02/pxv3z4a/i08zwT8Fsi+zveE6Nms5pCbQtQQ1m3AGET/7VfSH9bMs
XkIu+PdTuleKDYk1Nu/8f8zif0Id/W0xZm4dVJSkdtgU/HLjw9OjyWV/VVD1PMBTtLQbFaTgFe9Q
SwEFXx+xyJhVG/REGVytD/fdny4jSJGq65Qhv7pKRZwXDawfLYp7LJ7vKbLHRSp8sHUYZ+wrTKQ4
aP3TaAvm6g1/p4i7f8mU/SFeFdTWCdmzbpAFQ+V4ldzTmT7wh79Po6808qvKtA4/xtoaE+PqA5MQ
zH4btx2llJdBIjxeazwQAoi242bILc1nSAQ7IcchexX5WE5kT3SIqmDYGtCjfih4/NsUw1CnmRM1
nFCEqWEqee7MwlVseodiZaYjQ49Vu5TeUTBs2AHeYRLpQForw2F6LHUo4o4obwQ+6nd+yNUpXYfT
bKPjdb8gxUv5DQiAlnqY98Fww4SNM0YREVUMfxV33pyQFpZ62MbeOO4OqKAgZBSbg1U6207vDw4/
rS8+9ie3re5DPhKjflOhtCvqgz+wpSQN7V6OB/wmsBWXGJmRSdX7U8GXAgV7j98Z58NIvgHR1awG
zM6JkjamRB5eADdCKcIxcGMUcsAnvUkx+uGC12x3DNEDHrTrFZgsm2Ts4xv0gNVfchXMaZ5AgStF
hGLHYbSxS8uXUUBEX2xiEVkN0pXQfskEdWIsHedI1MUiTCn6NSDeIPNQ7rNNqKyqHdPOWV16NF5X
Z8ZGDNcA77ajjpbf9txKQG7Nw/n9pi5cMv4cZ0t0LwKmnTd35ej/TGnS2lknbYcKBGMzOT8zGzh9
PkURyjxa/4XAjk/2kyN4E+kWZkhN7po8Bzk28nrh7/Z0sfsMuLis6vI/USaEYi3HF8L97602AIjg
eJi+RFJof8S52pI9WVWGD3TsKZ7fyAC0Y/s1TYsKKoAWRi+5ejOUuo35ZjEQnEArjKLAFsb92rgu
R28pd9lT3KTX4JcSoOLjErlehH/5k7Pxr2nequ6uQynGu+gQyvXbEV5h3G+xR0dyIjJdeL0BUh8C
PmFuDYuUAn9+qXw2aLnc81+uK2uUfYn4XX/OnZNZrZeyPFpNsQ9csQ/ISz8UFMmE/8nh22iT3V3A
TTlyZkfYY6P/KJuVfebDkCLtOkWlN0u7Kfli0XW/VdxtWTNgYGjeNLbeM8iWPVtY+0gd+wpALQtl
HKd8QcRkBU0waZFtYp8K0h5+IxQabJm13qHa7HWU450R1b63eFV0JKxdVeSU4lO80Fx9ObYKgT/t
mcGsNE2jorCWK5Oo4eYkK8kTBoHYH349F+3pu6bIaeySxDmBI0CAsbSScqZJ/lTJEwfNb6Hrisku
+GAe/L0BJe47yeU68dDv17lv7wz4rLAUnWriMWxISI9X4sEKE5DktiOdRC3Tx7zwDR1CN/gT9dea
+8BQdUa1rZUheHvi4FAxsZbPT12TiTzvZzcW4krEG0IInaY+pltTsSjOxSGFuW0NLtvqNaiFtxEU
L2ewG9G9C6WxtgB+Z/1e4qZg/SPJq7VznUfVJFACQ29ktV8+nzFFflZ5jE33EgfcOMKVDg0J1qjA
zwLewNfboAGM/FWWNubknMR2IW1gThn7U5srOHPZiMNS+S+iFStc6ytyHx5+/oyLTigqQT0cWqiU
Mj5hjUhowmBi6aZL9zyIw9cpi9HO+u1NXMmzWNcNiTWieR3GRrVlHjmY5kPeCD9vUj32mI6IUVdH
ka1C3PXzxpUFpFgeszd8zx+ceLF4JmJnpwlUT6LXWWocejZeWYOajWiUaiUW8dPHS88j1k99Qcmu
PYLEZ7IyT99HU9VnKJSRJaR1MwTo7rS7J2KYJ5bhVLQplYtJXW5tr5nTNmnIN410D1SjSZAKRJcY
gyf8UfVFQoYIpOSLhhjtR40np5iPnu32kyNaSyE9Gf/8pgCpGTXFXJi/A4bPjjd9RpdGhwIYxutK
3ZGHqx64regT2TCMXg9MVnSqCoi+JrElGHTMOEFsxKM8roCb4gvxfgbJzHij+ddZm5pKC5Jwnc+D
yF5xfvrfAvVi6lYCieszrpDNYAqOfNpfMgmJvHT8yiXE/1TDrnl9/ceVLqIiT6akwTpbjwBBnYik
yFtwhIQHL0cORK2+V+wGXRs9lkKZckxhekR7yIL8LmzZeYMsEHRVBdgLTC529upzR4x1SAmr43Fc
Rt1MbRBijtWCerFp1f178gvg8G4wLvYcmXK5DsD4zgxFyd+WW5IELjy92zNH9IBf3ifl+vCDrbeA
952VNgEGeHJHehx4zlRzi29wyPYrZG7L66269N7ge6H7wydF2SoXI40uI4Ef8f/X31eo2mOBxBbe
dDsbiB8f2/2LlOGYcYENDCu849pIeqg2Ow5tDf7zv/Vk+XRhe2AGw1/wBnB4bPdsu3qNaxEBEstf
LgEHT1AncPqzBExHptePhUPRI2kAZE+4JW1wMySzeOjspLGYi1VJAqrsPvHzBqo5ajz3wT19RvSe
n4YD3jxH4O9VKNI90XH4VICJDg6iO5ii/lK1ayPRNUXgo88mUeAxzTzYjAFdRUP3mkca08st4BMu
5wgsoIOmMhmjC3fLpakQW3IFdc2C4qeTmpW4rf9H5aI2w1SIUnX4cCwXNxiozb6yE5f2WnitjJ/e
ezTu5ybjbzLHv0wZNy7uKo6oimFatgEch8nri9Gqy5151hmwQVokiHh6qQZjG3a6GG0E2+4iAqCB
O20+1WfL+VBCCw83zGZnkdvh8zOILmWWrMsdNqSyf+Xr6l6UbRtyBnvFgRcGBoQFGV6NcYzI5B4M
LdYQMYf0mRFpCHh+IKFb1Mk32x98sNmxwg8cQ0N6BzOcfQGbf6Onrn6oyZ5U4E+MA4ze9rYHfk+n
Ka1qNBBYVNsKIR2E53ZQsC0w2EH18weOvLIBGDKqwoRWZEkoFYR/JRgChrac1vF69xZHskde4k3Q
BL46P+5GsxHRllwXOQA=
`pragma protect end_protected
