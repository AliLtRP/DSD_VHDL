// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N8zuL3brYd9NKvodm8SEKQYmhETWlQjIBuMOu89647Q9sTYmUmqJx7CMlGzNSRe2
zcdUORDUl6xb9rPvuM2dupSJeqlNSMoX7S2sTZ5W/6xMDOEngCDYO0Hnu5S0n7uJ
r3q0YW6A9bSdUBYLmsmzTCIL3CEP66zq+/s8G3G8RwA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6368)
VxkS8ldbAmZPicu8hMtNgJI+vjvV9JKRwgU86eJeQRNZ8ghkd9vOcUryedTIc+pB
d9VKVvKoZfU1qMxAxxkQOpq0tl3QrRnquCIfKMr0LseORfHWwDguNqzvr+8H9Lli
BcE3keZocCX3sjSvXIE8iwmdckl5KvetDryzAVA6nXLR1RB4j/5NXKGVYEfPwVM4
xytO6AyyGDjj2JRwqpgNohtoHBPvY3ruz9vgLThFc2tnT7wL0i8v64e4RQbxtfbK
5t6oRhZRbnk6MyvNz2xJT+wBVjrnP4z9txsNPH01kuPk8RXoBMSHgYBj6Gmfs7tH
EnDFUfRrgiGoXfu2IzffUuC6CWAb4zBFUDAwXsG/lb9JKNBnABAOZXP2u2MaKkCL
zKNHrqEBtdUrBR9+ANWJIgWq91eO2WsTLa/iAkFyrXp28jlVIY4jq/8CHld8LOuu
+G1VFBWxiSYX38Csr7+1UiU+seSEcVgs9UHkQsvrfQeB1uiHlacD8CGU56hRxd1g
XYcohwk9N5lnF3bhMVFLTg5Dcus/wwCw85Bm+zpj1UTGwF+zpH0AJTWxJ0gwK2Xv
lsYZyY1YywqWr9wrjYhC97XZEDu1SPXqxqz6VTF3EOhOM1wNNBL+hWBAuRIYRbBZ
wE14zrUO5/kWMQHF8yqGnMflIA4yE2l9bqd81iNdF+JtK1BisiwLNJEisocRXWxn
IWm0tfKj2VrZx42Ri02Qal0DAwZTga8sNWAD/ZQXWeCje2G5nZBNSKof/RCh7fGE
AGzEXw1wiXQYqUABaB6p5vt8PWQOhdODTC7B3scaPsLYGAp7Wc7ZOhLvCfkfJsNs
BD6s8tmLOGME1g3qSVx2SZN6gChb1VESbxSNcprU6EO/Jov64EsR4sa8KuygMrL2
rTqKyCwklc4LhK1UpZGyFuR65+ADIGNVb4dSxnJCmn0wSK1YCOcbxqLejFil7HFR
ffIhjuU41IOUr0bWSmTCvpmztPQJBTmnVQvOf3bOOQBsv1zyHZzeivYcOGIQ2Cru
knXCuknD1mVy8hxMC6zs2uaimN4F84PtBn9lPycMvIm1maK/L+PNSnC2qxazIowY
8qvybD8+uNd7sdlCNCavUQcf56vuVROuU2X95vWMZ8Ij4joTYTGcWLbvdcq+n/s/
2jD5T5i11rXYROD5GlWgcJuvNPvFlAPfROYpF9DYQnqsd54Gblv5nG2CzsgctDor
CfU4RbaEdIewGIRemmNHV7JuuUj1UM+9w13SVybtPxiFrH6lsCePwbWP6rPdlSdA
TXrVmvru/TyGY3HysvHEzIuck1V+Y1LymjqX3RJ9WvNDYxT3oeZsPWq1oqPGOy7W
Eqtl7xtkxHTB4VRsKsBo3EUvV3CgUWKFN0NUMweRQ8PWwJNasaEQx98EmGjkyGUp
a1IMqjYTo+OXCmtOm34zekp5oLfrkooCaZMB3fy4RAu4ShJGhbqXTUzWM/R7koEX
8T8Shwrw2O24E5LQ+lTthquxwae/8OuLCkTP5eGLKP5Yp57Py+fA7DzNhPWPxvqg
BikI0fDfUGH1aUDo5E20anzPRJyy6nvthus1qXSF9HDS+aKaDFplYG/PjXwHkJIA
rCX22WsIBsfWEcPm4yMQai9gHeHf37OOoHzz4vdKDT7GamTqAs6fTYwLnDW/gkKi
d6u4runzVQYYxksAgAt5n0/cSrUv/nKRXjCFbJPjUxMvqcts+u2Km+O23N+ccV8x
5+HnfgKQOw8M9/e+XXjtYcxLZpj9s/VfRawwLbxhgVCZHwOgPVUw5a0R/ejHj9yk
SBVHN9CQZAy8xapLWWESL76bgqRzrivf9BzyzjLknuYniu2vT5nMrJNFtb16H0jQ
euwkjVnDUq8+QMmK+RYvKWtDaEFYju+UMyET7rYPl6LleVU+13NQs0nDLqbPZMEJ
zWGAn75aPF0uNSeESuDPrUgGbsHPjCxk3ZiAgR+iiNmnsrjVdZTJMIBVda8vQWjz
u7RXpqAyNc81hRMkMc6FDtCG0TBjmXuDezO9sWiqPlFK4sPJdsRQIVIQfIErqtTM
fhY7zOqNorFdF1HgngVhBZaAGXtjCya+H1dBO60qjFUQskSGSjnYaxOH2R8AJh3o
zPBohcHHMWjxKszVX5jgkJGza0YmZK2IIABdrEnWAkgKcBM2aYVjM0hNlN/I446s
1lbqbLc2K6cxufNWBN9EjJkdpe2VIBIKSy7T81Ce4dzhlPqkpnM7X0F0h+DeiBi2
V+s2NXZue7PJwoGzqVhpyVUXQz7fuL4TpPbH5T2I95wvd6mWXEGIEAGrVQh1WhpS
CJcyBBQdQI84vKS6/gAfbhUt99xgicLOmF5OMJyB8icjVixUhHo0nk8Abucwqp25
BQMcXRxk1RiWSMarnTBVpEGoszCHCBaB+stB823BKILY2PjSyPeP6C1vbS+LksqG
GiiNaMGJsi8RwWz7pKkjdP0r8wnaz1+KHKoAsbGN/40d+ijpBSyeWkjtqsoxrC6L
YbrTMfsPGs1LuYEn51jZclwDIjRG/nj92JPAqda1W8MwPNhItsCI8uqaXmb5ddw2
RzwJi630XlUQPphmtG9Cmw9K+Q4Gs5MOiCDL/oc/yzWsCtzmw8lF9mLF5OGa0L+c
awG4ibS60TxTLTX1Qj8O0h7ieMSNKvKCab4r/t4XCICoZ/jF1YDGYhySIE+KwCrG
SqeEZ/pzPFkAFFX7U2csbkAW+U+yWjH3qa42QkVgeQs5ySVtqWTlfFQiTFVDlyqH
JXF91FDrHiR6qUfNOItPLjvWWsbS7k9Pels1igPBt46+EUG0Gr0xUULmdAxYx+qC
H0dVOYt/NTfvbls2Tdqp/lAn5QzKyeoSveyyvcMbVvClQAmCspXHByHtf6/128S+
nPl0eX0yQMKeZiXmg+6zgFMQ9jjK3fLzTeDMUYchm4kGi0+GZsTITqbVbQXH1orP
ZeNLfKS+rbVh4UxX4cruHiOMqyQPMskMItm9Y5nX3BsAMc6QFzbq173ISx1Mabv6
XPJrCxN+tuc+zL5iJYyTCl5dc7+vGCxPQEeWFhzppgI9lgxFD6JKDaIVZ7bt7cxp
8BiUzzBGRGKFxrC4IuhQB5rQZjK5DpRvXTsHaRIhORRQh+09jokSR7LuxFG5jqNc
L/MbhB8dOkJvtXNm11g/pjNmNx9CAhuGLmTtO5NiLDaLRUXALaesDUxKi0VAeoPD
7x8mchoFl97snUviUron3/QzzcQoVfIM0bGeyLRxWPQ/P/YXgaUR8VLespBKOX94
QcP7Flk74+nX5rZuUqHkZzSHyiqlezJuXa+AVKO5zgld5jNyGsQaHqmT01+IK5SD
b3UjrxcbfZ7GqrgarP3TPOhl2htcHeGCBO8fhUVHW0geDQRHNJH8JwOPWehTJJxL
B4W0vCUSajVEvAndsMTlcO1nzJiDoV6JSh/HJPvor5CBO4SGYSdS/6JrdR+JbNB+
lVN1gz3Kunivxt+dDgmeZo0Ne8yppClBoa7++DjP+kJ+OOhJrJpwK/MKDuDYPiHe
R+BYAx+2VBHljo93Lx86/6IaHiDMNRUxpyelx2fXaNB6yqHC0LQ10H7Hya6ch5lP
+rvS0tnk+zivqIZAc+BQyP/XmVUjGx5OvQ2T4VsgMAt7zyU0Hp37MSoLnOj/awDl
EPMBsoo+3fZw3L97q+pm4/s5yk8EyuiGYM5ipj2yb0vPHHuSXlTj5R6yTh3Oxcme
UxNbidy6RPwUNPonnCTm7G12Ciy4SFewTrm7ibEfqPovv3+o6aQbDhg0gAU0x9WY
h8XlVv86u5JO866kQR+IS1jvVu4m8cBQf+L+kZAorulF1cWfAHCJ5gMSnre2eScV
FBOiPePAolHwJfwDQPyqaML8t65+kDbEm4rByQg/H6jKugaaM288/Am+Pzsa4nAL
n3P0ThXNGqkqlEF24T0Kaa3BJd1Ob/B9rNbkMlm/6djRyecjmBSP4sSFeHCSpmvB
dzlDTIdj/ara+teONQ7H5TVp+T6FFkMkgtsDJAH8TXfjXoqE06kpa5mL3CfkOxqQ
11HXC4ROKICAYomghZjWGCaE8D4Sj799WkSigQ2zXFtTNuSus33BoxxuNRN0mOOj
FlEWwDHppCILLb5w0jpcNFj+EjRyfKAr24cmUPz/RWSwGgNEbk9pyqUtxFJAzui/
iVPAl5dKs40fWhGRt1WlzgThbU1idqsYN4EbBYANg8ptnI1RQaDoegvDVxXMoOGx
oteehSDia1nCSkoJeySEhlTV4psAtaQh5JPA2mF2B+Q/5rdQXAilXgY/fBStR68Z
XDluj5Ofg+//YwPVMj8dvnJFlTbe5dRMrGp6FUBdF47qU8AdZVy7Z0ykFvNm/tfA
EGVnaCa301LgwqvvSmgXhkvqyC+clyNJuUdlzB7GTkeowbYm660qyYkqMiVW0eEQ
r8HDd2W4imOHwuSU2DqflqWIbGY7io6e4g7b6x1CQBXGXrj/G7LEKB+4XeztFuVU
EyGzAxF7qnx6AaMNaw8YbvUHaIog5LworwSfuw0shfTe9ID8lcNZSr/dIMU02pFe
ljCfNA5VXA6tPvNn9qIQaFBNtYLdAPs8vzfH0AaJtj1x0JV6Zuz1/0D6WDlby352
hINeULiYA9p+k25tf/pm8DsFgg1LYD1uXHAdwN+vP/3OA9a80qNT0CWtV67+dHok
vLz+K7rd9cNMGvJNYu5AzVw1SoSIiWb6nRMSrNqc0pCZbUgHRGLCZyMwcYjUL04x
Aq9IOxcI7grsNXu9rr9i5Ds5QfzhfIyEq4x93rx4gISc4VMy5ba4NZcjc9VI3C12
TE9lQm6gR/12Z+HSFNBESk+fqf6HcD/g455qsMfa4RQtwibgvvnpW7RFmikU2iZY
jDmpihxYQ2FfOL+y6wSgT7sV/zL0kbf7hAGx/onZo2bSJVkiZHKY59mB0KhxCCLe
y6lanYoJO1JAU8XLiCI0OI1jXHj5bJMXnP8vuOBy/m0dTaI6WwKyO/DuCv7cKNkI
xTohu2qHgnrXW3SvAODxb7h8LQZqPVt0JHtDjWGME64WoNV3Qbk2odBuRr1ISMHu
ckCBaOTwNzUcpjVQNcjHgSLwQ3frDPn2jKDIIWy7w/1fYVoHjQYP+jcnjJks+B30
rcLDU9QLbyimLCzoevUZLNkst0H0zio/UU1iYkHuzrtlUqV0BX35/v1S1fygA/yA
Yg6fblsbZ8MVMGMpx2v7cxcYoXXXV8zWI5WwfZnRQkKL2IzzW6N5XQ2bbbKtklCO
51TGP8qOireqecfHGIYU9/rVpY0d2Acz9pO0R8LsqhUSM2PrAdopEDx14NBXiicx
lLm12K2Yv8ONz0Xe9c1xkIkBAFQ18T0w1i8zSdCOVT5E78xxOX2fZy3lI0HubjbR
etjfe+cC16fJR3EwOZW5S/A9SNdkLxy/cMBHnsXl1gyOSFYOMAEfR/lGAikkkuVO
+Ab81Ih6yOK2dQdv5xrpTHCOa8IbOELaSKJCbvQav83XQYe4ciPmEyrCsbhRrh1A
7BrDXSb3aORnanV+33Ry/ym4U2PHeebTWxEJvNmOMAd4aWOWveGwhRCJdlk8bGac
3LGXOI8HYdGjZdywJJ/u+NAEx6kTSKJNXDOwPlnSBiV6UCam8r4Rft+hzvnBOtxB
Ws7SyDh4q/9cGPbAa/5pbsnueDPACuCESuC2ISkrfOo96tWDwwYrzvBfX0uhwjto
bgWaDfUFYR3ANp9gfdcDxru958TNF6S8vVOSd4L4FXjeXEo7piBzv9IL4u7nPjp6
PhSSiw0WvDE0l++CraaOoAQZlHODKKpZ17ft+tnEXemvHGubtfZhYoKSDVIhIZsb
P4wvq2G6NsuOLePL2xjhVLq2eXYnUTSzij5tsz10HWNbYOZe1CWbm1giFViBWJgO
0mLK1olWS+T1xsfpbZtki/dJ8SYFw45Z58ig9q8FWudLCyYA6pvtF225WAf4fy53
eY4Vh2wfmb0EPHIdOr288N+Eu3zL7sf1pFdRl9PYI6mTafkApQhRYaksJvD7mHTO
32NmF4lak+Jf7wYhhoTwEOyTM5UTczNpQJgAQKCcKd1d7OFJ3Mjdi3Qpg0+67RxX
ehIKNDN3M7lLN3z9Wa/Kjn8oxBSIWbIl5+y/r2VqpuynRC8jjUr62yw8VkBnA14i
7OwmQgsiHBX3ZMzY0D3etHvOP1qFeC0F/YeDYoIL19xivrgDevl227knH773upjH
5XgIczte91lz28ijJfDjRVxu7z5DEZ5Ecj5gi29gkpLZ1jGjvnyekXgAdbiJPC7u
C27LIDsTEoiQPZWhUSc3beX2LaiGPabXV9wtTh8HxcBrrgggSEdHWctSm3v8pr4z
WXx31B94pL0N3+Ck3wJn+wvXhSMyXWKACm2xwgHqFqYCNcb8oFyz3OwTE7VTPlt9
Ya0oQedJIpAc/QcaGKQdQ/4iDeewut91/PxNKdBszfQJMr6aXQnffbGg/pbeYvh3
YdTb2w/nKWz9W3oM6i2IiLEGQEDMX1nbYRDraIty3/eTvPAyGbm2kMq68zRgRhVq
SMgjntXiZByg074GLgiNo1RhAMFGk0B61hZb6v+CLsmRoIdP4bymhZGrqE4F1cIT
iy6gSkgkcBtCbyWoMViH+YXJAcLLLFJRl2nrrEIWRgxqTVw9h3QqX09Rj2viSLhW
Omm3/kJE8KTzo71D96jiIVG1q+M3HPxtSQYrclmUVDx/6dGDk9yN0ffbMNxfVW0L
/58+xOUWD2SrssaGB52L4uz3QghwlKiIJzLs/VYNmI0JVDRQPgkcy/cikbUQfSBH
zn/ewWjTUY1UX25y4mVKyoCTXXE6+lyoYhBw5UrfaBKHAHP5uFwWsts7i9fDqVoU
Jr3GEDdR7IKoswp5TQuTwOmBWXqBHcgeiZIYl/hF4zukuOBBa2m9ECoqu/QrbKIx
EEGHiY+hKQWX8gs38Avy+ZspX8z9u4LBOnz+AMGIpNdV6LjxsnQuZ2XdRsXoMaiM
2vtqdiINfKQ5P7mjnKa85rkID4KAqVv9PtqojNdDw3P0bYIdtYfcl1FNn+1MnUjq
ArZlMI0r4XkBhlXFSRdB7mpah7uo3XBeFgRLDnOviYAZ20UQuQVTyBd9qz72sv4v
dRWwhlT+axrl8ZGdFJpfBtFQkMFLvU7PadzIJGz7s1R2MsPdbiXZ0rWBkbKrVjs3
I91X3UHV2hIHhB4VlcIiaByStcSi+l55GVp8tLjgBCci1nnAo/dZ6jnZtk+kN8mg
VGjW3QPpDDzNw0w3RQffbY05hQVOU0wGXCy7+7Wdbwf44LeObqZ9w3xr33B9Z0T6
Mjvcjwx8i5Lvx4nQawXL7DlfpTRIenBsv7aJlp3mlbZiRx6mbuh75kU4c3pkozSE
9/Lcox02JHR0pn57coI849X2ED63QfkdcAyJI1pno3UpN+KOaz+YMKpcNbgNKC2F
bcvcGsw6GM4QITWUu+3G2qVT0SGJlFKfB5e8KklTlYeE0v9kgELcpupLzkmqORFv
4uiPCdEsI9n0cJFQNR74OmYacy5T2VN/a9ikw3EfH5SRrsudRsSKxD9yGpsQ51mc
4Nh14K5OU+/LYrUeJcr/Gtonw3XftU9DUOVBJGdGcxn5xdDA0xwga9PKKLFIwEAe
UhIYWl+yYs7xATs+8Dv3RBWWBI2syZQK6B73ekmjF7vOuzfOmT9MNPe0Z0sVcYGS
4NuKX+E4yDhGO6E6gNRxlLnWxd312OfUC4zPxLgrFs3S5AQ0NB6fOUk9eDTWhWPC
Od4SBZ1bALWD3czBX/Gu8/jh9wEXgA0T5VFdUZfRCkamwn+EQnD7xoU+fjLW0uJj
97B/iiBSCwWyiaIHzuSqswkxvMxqwsP5U6WlJtLeFh7UC51vVHSP/1m4GUheaTHl
QZ0olrfnrSrewcnpe8CggS09n70sldNCswL/lUSrEiDY6CxB3mP7BGTKgbTfXQOH
mWOBnvPxvRIkBZWht2h4fY/qxtWHYOG4nO8FrULWBahmoVOgyHsQzTdIe0HA9dH6
YftYljK6oDobJYq0AKsW6/jkV4+J51zEtr8g621oP+USfPIhwIxARiKd9pFGnne8
pI47CdR7r6JFtxXZ+IJuHrJ5g1oI4PyaJyu8S4Bz540DmjssxVWVcjXnx85cs2l6
Ablu3BTXai9HjexQDBdW6QeEl7rRMyyMt2Uh07XnQbGdStK6V6r35zK0jqbzsxmX
2j5OujnAVCqJajuHhviK4P+mYq77XK0GF0r5OduadISmq0MvwKNvELGsMtmjEWSt
EhvZeyC2xziADm3KmaBfvw1MCP9SMXrngSEIzEGicpdirugcsrd7zluiBLEBlrkM
Rg31zfTZ+BDU4zhn3mr7grUqNRf66xxRJhD6QBhgKMbhTpbFd2p19Xh3OhuWQigy
rRGY3Y+b0kzNeyPqzVy18GIgUTu6gLig9wU07hCSZjpwfN4goeaoobzCrMXXnOAI
GVbP8sqXZXJ5KtyGFYltFCl6XpYPFzeP5p+ftw4Lq94=
`pragma protect end_protected
