// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sUaLEzlAVSGrRQeH/WH65qL0ayeijl75yWylIqixOzxzNWgxZEv5S3KfrOOSI2dG
rcP8hqfy/MeiRsP3GvHI3oQda5pbh6GIXpuGSplzxOGRWkh97HOwwH4BNHoQg4qQ
10wW4vNEMvxBY/J9nCqbVXaCJ8xJErk4WujGD1mg+1Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61984)
wGWBnzmjiCmKLhgqyczCYCKWkxMbr3JYc+tKFV8SRcrEd8o3SmYXP/UJmveLZLYD
omEEAQqEQBPUAFoDU2rnGdEJufXboXn1HztP0YH+7vUUY6mVtzA5yTmTRYKIItfC
SAUqW9KfqHZwGsvhXT879MRIoJZjZ1nKeE6MT8NvgeoBIZ6KsiX3esDBwkqWboL5
K8pK/SdBosPYBRNig3qLNlokORGnorvNqgOLYD+u39Q5B1t4CjPpT4NShmGfQ34s
UMUmcb7d3+tfBC6bqvARAk4iFsmr44Yqb8N4s0XWknRBXZ7Rv76MQ8FCtHNp2PGv
igi3GxDSI2voPJ/tTUroEYBeVaNmToS9jpeNRlSdbKesYyydtJmg8BBS//yvM0g+
fsUFGyutxnkZz3x8r//WtzKnBpbCtdo/AvetP2+l3v/7l1aWWJR2tsFAYHK9Fpcq
KreSzDDZodVWmwAmENaqK7PIQnsS7UmKm13OSZ0yx5ChExWEYp4hz4cOH1Ehjj6F
QYNwqCrYs410uZetvjBKtGKPPw2xvXgDCcbjzPPfp1dmvPotvu3y04Eh2+DM7PYl
bazwzGpolNqS0Z3R9WMX0jiClr+pxpqRibU3n+WEt3APNJPzW8kQQ9D7qQs1ZLr4
ZtF4cK1s//KqFNv5L3cLMk6R6dpUIb5rc4rz8bn4LVOUyd+yUtymQExJf5dGeKzI
vZtWdw/saLRiIuaKO4+xgri0Pmv/aQ9X6nWSMQgrTL85rwd+q/i7s9wstXgYs2A5
aZOhYnosx8GXgFx8LPYIwOBmU6n01bS6zsj+tGOgCS9cTlTqB71Zbo4anDj0n7QK
a0IPauV0+jQao5ZuCIw58oEyZyzkAVZCi7J5B9qJobdYy9LA8z1654SXO80Ifhs1
eJNG+zA4NRfS2Qum9WpKPdX1Xvg1fjyFwYxzgaqL/PdTd54YWeCy5FAbBfSlJqqr
W3H0ZNwyrCGOuR78oe/dNn1PSQQhZ9o8LUO/D1d0465JoeDg1A5FlVyXqgBfxRBi
XQK7fvG2GMpMR3VMI7t5i4XXR3GEx4uwSd97D4gZjNViAWXma+R75GZCniSyDxK4
cwmRAfnfR9UBUr6OLGEzWXynW5CFCHGQE0BdREXWCQkj4RgsWYckJ9XHWI4zG+nv
wNEqVf3heqCGUZfeW2CQN5g/hUG64Dm0lCa4udyqGPVOMbyqju6PTeYM54aJ57Uk
NIlIKTDssxR62tyUIH0bf0VL4xI48EnPrcg0dJMcH4+NZMxMsXc8ZeHD5I4lg9/A
h5dKnkBhLoiXN4a2rMC7tqMXucLNRgtRFT9fPg8N24vkGBF6zgDC4BAmMo9sVmgO
/2Haz0N5fphqGoudrwZ38YbH5dC0GS9xmWaFN7Z+ILthfdJxurUhk209W6vWQM8j
kwjnpGIDioOs3rzrLOmzuMnlxdecSi8q9LEJRI5zoawNDraiO+5tS1fK8Sx5sp+M
zSSPPDmCF9XheyJ6PyXtZ5kgFjE4ycpCFlsDdYfPlSF0404Q5YmDKVmXTfchwvnw
0D8sViLYDliyA3BFOGqSTASbNv8P/rZElM6d2Wpe7WZvT/3acPdbPgAnwYOmRHqJ
xecCuhZFEq/h9CeNlGjrW/AcVSoRlmsl0S16VoDZcg90EeVzs6yr+AGMkn43S7ZS
sSbrfy82Oj3QYDRrkmo+w9RvVkXyh2HYOVXgbJAMtA6Y/J57NLeO4SOC7cZljBfa
VFHdF1J+CET1gW+zTzR2dxkzmCEW9jxCcVM9IO4GW+QoALQek2SA7j6Gfo1g0Dh6
YbHJkCYPRQWWa101F6U/43mhjg9onHy+zdolXR4Mf8KUVxmKhBI5yf0JcVVjpQWu
r4gm9ZauYn/uf21+8wjNysFjT/JhPqNNf6EQw7RN1vOGA0lSvAiVsJbFb+QQBoWq
qDXMmIJHkM5fJshszOlo/tMGuekW0/7Z7ww3AU9qJ2cpMHgYZcUgvF1XR6OJ3VYr
luIsXZjrq0ReaDNqqLU6dwU1mplWd0LEGp7Fpvt8DE47vuzyTd5S8/pYXFHUSeFh
UKaLH1kgpKTAuLAvI1DNkt4mdbMf8ULg3LqDy8XyPUqBZ3ccYlTzwk7T2nPRZzxx
gg7lhntwOe8ahhskQPSuXvF4+BLe6Axoa8rdlb+Iou+MccaOAuPG4qIY9jSIFA1y
t4lsE7Z6nt/IZTjkaicgFq/gAAGRjRKNrj5fw5Gq8BQLPJlsRrOa9vmpZKyQk48b
3ah8aBjX9Ot/18atfv5spcatJhOBHeqGigF3KfGBssfZ50LEVXZOfj7hqCwMXW1w
cAjoHKf99FwC9OCOOqwxZQ2wH5c2Qsb0QqJwenMlEYh9ZT1vOejENNTjz62TmboK
yHNqzzf9y2oA6TINXDADOWDDxIOJPzf934rhX7JIT6et3KvpoF57Eh8px/iDPWP4
69+AiVhQ6qcNJokRrriiLsvAjwjHHnjhgBGXTMylHvOqXOVG9k2YMEsiF2R4E2g+
igJQcgljau+CF8SFhavZ6zcr7lIdnP/1xVKdtHJ335a/LhRS5vdQC2A8jFWk8VSd
yNJrUKCodNep/VOeBuYpsvsoM6cie4urN4x4jPFgc0a3YHu6tOf9nuoNRMMKCTqv
kQcwlQBWnMLkmbHrUxE8h28VRH4Ajwtmkvt+IiRZVIqHONpD8rDyLqWOYrlglxkN
lPnGaMTxtbf2wLAqSFhBxkaIJqqcuwyUWoXNR+G5GdxEMD//FPlJXl4kX0bQZ8gF
mXOaoPmYoEiiMIsNAHqaBqOa3bPahOry2Dn8Aiy7uX2QePbJxqk3aqdR/TvLsF2S
ICVhWFIk46EF5/ho0+tmeh29cx/CoU4iELMrupw5C/9EaXv69YO9K7znZUOGb7gd
eikO+91IamuyC9UcRpPlA8pwq5MsgswxmtBEyKofJxlfeWUuy368XQVuobPWMe1X
K1Ryeph9EzAGuXONUGB3EOsBllOyjPI3QECVOlJS6ynCYj0YpERWKr2JjVAIf1u3
V1lLzaWZguZMGIItaEE+iRwF/6tcScwjoDaEgN6xczLcM1x1q0Xiwr2ryaPFm7gn
ePgOmrbFWX0retYXDO9b0fAQRwZWPN3hUlnRUmeMejqNF93qCWm8+T8W4YZv9vAk
+6iGcp6PnBR4eR2ogfhV1tB2i3k17DLuTbYkrJKIa0AXfFwM+Q+kbN4WlrQLVdWc
qzyW4lhXuorYbpO5rnD4bJkfEi8t52BLXQawybX01c7lEFk1h8IKz8cqs8Wckv/j
Rn/P4cFmdT/GFjHx1QfD9prswYYu9sGqdC9UGeJ7xBBieEU3w9ol2mRYfSg2Yb8w
2BXjqcq223Q63Fwutj40PNKWUfRnE2Xrz7XKx5y0fD29uBvURT2KINw/Gol4ObXL
HCcKAWfXuri6DpbJrDnQ++NJQT3wBQQl4/l90AXJDg6cE6L/fX2ofF0BgcQHXrTr
SGZtYguhw0vy7Kp4enx75ydvZB97vgconNjK5hby7pXJflvThVTpfhVfNMYKOKCb
xTk4sqNghWXIyWPGLCo2cItTJ2ru1ZtMCjftd1Gcs5t6h7ubbvzcRPHLT7eofLOw
NCKshBvEviwg5o8SPQ2Rxt/HrTR+XA1pDZGJgF7Cd1ZHGcIHEb7Ol+JY95Hpq6JS
xr81KkI2J+8uoqS2WPDuHAqfHaj5M2PeATNdkvPkdu+tszclaraYpoLlD77A2IgG
QHpboGEU57+VYu9BIdKcZT7eEH6+SfqYTEo+XvgZaY8vYzHQVB7jhRmXOaIpGU/Y
tionU/haUEBCecGofxD2tS2BSYoNRDnRKzmI4L2cE3CNSkfJLQj628nssOllkS8K
XqI0dh1CuS3Mz4cIxZ7u50JLixzyA3FjDNMyaGvaAHU/F/Klp0iN1OPS2hpD5X38
PHLRGLT9I2PTo3MLSb8PdiWy1MBZ7IgNC94bQpQ++xAnzylS87yplNBh92RazSQu
WqUp59NxBuZSuu70ac49+U15wWWSibRYsk8HNht0qCyaci3IUM31/L1eiKLTzoeP
le00bTHjk46GrQu42GWYmhs116ow6ZthR4jRo6xX0u5zIrHhY8DxBC1v93X1WEvp
QrMoe4ZaknprPkNm7jxEHV1sCJsTg7vJRSgx2NyTbDrKhtZAS0MwRPIdtHGEYJ9j
VhfaI33oJp3RPRDMSLx4LjT8uTUpWeoCFiGHrmWM99eJA2pfwqMYnqZK3RKQH2aM
uuj28R0zkq8Zs1kFi6Xe4QHw2GaFhwm2VUV7hASXV6XyhDXcrVPLau46gNC/DRbV
jVa6EQX8KdaltbN/cSbbye3eg8yj/TPYCiN3Ym6ZgrY3sm+X4Mjl5AMJ7bZYn58D
Z6rM0z1MX5vZBEdSiUXAYkuNYUYuxsVhdpewz3HALpGWI2IU/FUyCTN3zFtyNXlj
jxWlhEdyAP1fBgrYc7MzWjmnqCJe9wGpeIMkPeperWw5AVI8JZiqs5WxlMiXccGU
K9XIl1xSXEhxPOyBt8KvAzUJORzHTL1jQdVNiLkndqhnhP+Wxa+96nrneY2SN8wj
c4hLlurBoLI1qLltFCx2/VMsc3lT0S40HzsrdWvSgwwB72A8MJHejH7t7LQ3zwrc
LgxbTt2FwY16enE4KXy8OXrw72IaSSuXsbGASKkZTEyg0VmL5PMvDoh2fAumhb+N
8XWWW6eolmWTXB5dqfUSDF56Y1wlLq9pH0Fb+zptCTJD4u5yp07h70ikDbuDfOgC
HPybGS+mWo5/EUMh3FNt+rZVB/kWORdM28iIuUUsilZyWmx2Aa44Ik7/BYNm+RXK
cdTgO5lMprUPhK7mwjbq58Xc23n2Ug7LQu9trlsxkQuUnTjjGSuams12gNcH3+fh
7T8sfcdGwRknzc6yCRRE2a5UTuUzdVcw13l3sgCFHM+AOJHDFxlh9PY7L8XMVo1s
+5A3kodlKXAiNIgkfmBwOAJnfXFDaGnV8CdDRhYs6m64JSAU0xvnFa4S5/9e8ZVV
gg1/qe+dmjcUUYFu1KjDFukrH+H42ks9sYuovgGkik5J9T5F7vETYsFZefq1eVZj
/0EjzNwUb2UsKYdRqFkMC6qp4OgpyKXmCXQgmIRL5b0+lKUNxCpIrsdRLKPuJKok
5O7K/CR38DXR3r3eWpRIulEq6WOMje89cDmtmdcEbS0Ac+jU5fdeDxFiKq9kfITR
r2u7IJWEiayJkMZEd5TGsncDqNA81lgah64V8sPXE2/c4+J29OVmECwRWaBewuVM
U+wlgydgsjRDMhwZkQ3e2DQMUnLzaBtN/myJZEmgRjkxs8khP0GiKRznwhasYXHU
9MlFZ1ddhDOVa/n0pA+0TT9tK8As+4lKbg4hHwB9DXo819ucwr38v4Riv9JBhOV/
8JKKGf5cSPj8pJHvGa3I64PUyfHAoov2ZYAlPnIizfZhkDeZHr5NNjdubfhQ8WFA
in2s6WCCOrxC29fzMJLAJw5yKKvZmCf0vlxzBmel4L5iN/SaFaUTgGVws0eeWcJb
0Rl4lnQ48HzYagsxM2Z9m2Gl/AkZgxhMQzW4o2oKE6VAWiKjsx+fXyB1N9CgmptV
7ApkQ1sFmWVzJWGEaJQuWpuJmYo3LBcnIy9dM4LBLtxKfGzlFf/AcycCy7drlLtT
OFjiVcuIhup0E/1LtOpUvYNGJHlq0M0nvGJCokJguCxEcpY+u1JWHWOehpnJP3gJ
YHodEa6ylVZVcK9iJuSEFvd22EeP4QOwulotrLRScBndhVSAvv7HGRBeHuFki9qs
lhqj6F9Vky1ksuaaITkeKjN0oIuLfOTZpQaVwcs6nyBZ7Ug5+UUnr80WpeQORtUF
Yz0pOCcGqcGP0VmBtmt9v4JiWW+8z91a4eEin/EmC6d2OR2Lr5fjGoAFZYGHffel
axoBNXqgM27fl01QducAyHGzAVkHxTyv1h7lXS6yjSRcktJ21ACbk8Hr9bCcFCw2
lp527dXWDdMrbOgRApvNjzc0POw10fkBr+iXSQJ9V2HmYu+MgK60XCn/MYfNocUX
kgDw1tBIuW2HKqu+05HXQzbIk5nx4vM8FkWZ73DaphBpaa7MZ1E+G6xjyAuP40wi
sPV05itRFBQQiRTsEdst63JfotiNdxMci8NeixjBnA2BBHbPYAudKJMM2gmz87kO
70SjS+68ra9paKuOqLQsMtL0fVMfj+x9L4Fr/nDuu1VDgqKVq4oxOUXfs9/iLhdi
eUpGsAz+Oer9d30xHnUl5PL7Pwq9ss1mDYR1QX4wWVHzdrhPrkgDUDBvGdScjdn6
DMOF/ugdJAxg1iV8WBRVuhBLpnqPnrUeoT69lrC0BPbIje87NnYAY7hx3SIYfKgo
sz6Pa0pXZ1chD6GV3Xxu5kUC8TLK4uuBKGUmXRg7wJuCwBSYtKIOEnSDECZ36opV
5B/Yn651H+Q8ILv0evRduD77hWT+Whk2BeaJawGcFBLbqiehQZ4fcp8d0+9cXMc/
mzcIlAuevLbFcH0PT3F922aKXK6494nj2x//vg9wmlIrSHiut3VydLoLsknDO+k/
1KFhj9VNZ14pcQlTmxlZVHNJaPGPGzc9THZXRtT3bJHiOxe9buVMTPTcQXXEH8pJ
owZyS4Ef5277SlFFCsKh5Ij2/rMPd1he5KJTbvjnQQB7axA2lhT/wM1IdVCJ2SHf
cZrWCXh1OCRAtmtDbzrRdPDncUhE9Jsrma2hqkVV6NJ/0GL0pUaWuV+8lMaARdFa
wvu6X6fRbY3AWVa+VvD/eb87PkWV9fhZ0BJQ93vXwSy2IP+uagUxSvv6EeXwzyup
e3TMxDpp5zcn4zRx86kiIW8zPXixXIhF2jj+Zd7jBaSCaHiQQ/3CtvuT3T/t3yp7
cFxXaSqpjZ+/XubxP626XMTqVhhEEx2cyN5ww3yGMicQzxi1gDrQ0p9K5oHptKp2
t8EnbkGACD32LIU4akCQWxarCGROuZako3UU4THI5HmCP89f7qgbc6jq9nY9ksN2
pwFFx3CeVUb9Vd4wrmvqYatdZMHCfCs3m0M4sZmSRaqMnU9YPqxVvGXzxOwGhGdv
9vdfFtgO6IF2M3jxmDLQNdk8LAQeHto3DlqgcgruQG/ILITbsnY4GGLzquSEWQyt
GlC+RdFmgPWXf+lpZf0On/fVFuOJEUQ2FpsrFbfNa+fzdXJNuLl7U2Q4qtvob3lJ
vwCETNiDYV4NbsLZRRBBdn39bGAcCkKAGtVfguun9xglWsVJRcMvr2XKogasL7d8
bZsJ8DDv2cdItvMAmEzO69kp3/vu5G/aQz37t3dkPM3qaJB+ykhug+auQyYGSr+p
9mq/OrAtP1nlr3E2rAEagzxcMD0WA4auNQzVOWpZplBIPQFNepsuWZULh4JVdwzJ
lLG3j9LBQ0t5bIziLZaX3+iW6qZspc4aZVgnM3WFWNd4SFLLZBrIDMj7NppMB83i
vHcP88Fjo8BnNj1FhdhGtDADhGRbRkQmqX1/zix2XE/5sGFxlclF37RDa3hCUmAE
9RWM6yebQQJRIyGJ+rJO19gKaLRtOPbXSlVtGXW6Th8m2C5tniri4SfPDrYrNs6z
4D6NZ39DH2c9XRZLiyZPuqKBfUptlNSUbsGBoXJ5dHr2C87mOVTw3XEW/8Cfi+Zu
eKgo2gyHgKPY2Qg6U2BPKwxw30NUWv3NkAVIBiPipURbcslxzCf0fNH+lNkwLuWG
AONLM8HZe+NT5XIL5Xg5wq+Ynu6pc8VLm4xiL7fyOO8er/6z5RNLjDNENElgIuAD
Fni97m+t4reN6Xg7ArdPYiFyvA5C5AkEnW5aWywq1WiNrDZRAuestjoyoFV8lsfO
H5bmM73t/xeO/EfQcHgIUIoa1YUk6F69wR7ro6iodZAF2NXgFqDPVMeOt3Bn6zNS
s6eGldd/fwe7pcq8snLhPoQtOO/ThywR6vXVwGK9izLPkYetMaxzLCOvAGj7IUgy
tDdqg+e9byyN6hxfDo0O7VX6t2PqIJu3K6O/FPo2pRtpG5euzb0p7hz8eBTfIXVC
aAXGyP+fBGhVjK4QNVzK3PKOYpNXVR0iGnM1C1A1dEup8xz1j7z1TCsE2GIXTarn
TgjOd/S1Xo04iZT6rZO8dX1o91iEaVY8D+foa7SdE+Ne5P44ZhQiCYDmSfhJ4++l
GH/2U05k3fm1j3WpDRDxyNw7rpMhNeflnS9B0YyFixNRB7a988GOA0vBWPHkEN1V
Qx6oj7YC9mRxm6xUKnnFqzIXDb6zbbqhzZxJfQhrW8RsSu6CQ99Bp9Rpguy+FLoJ
nbH+83bIosfIroHpFA0yCiz2z5hPC8xvgAPiVBZ0xY87rAKawad0jfQzrYPlfZYv
gpZ+e0AhKhyo0RUy4LzGF3tJ2c2jpMorUdPZzDBXswcw7hWMJS33SuMHi4wN2sZ2
j6nIfx9N+Kv9iVCP2TkC6LWbOdaULRZRF3dwI2/upMYxkfG6zgqpDVsN+/bTupbF
5/O6B7oDwwEhx3uhzn4TH8g0aXxUz1OoPPXhq7pxAr4ub23t1TXNq7lxJDGTCLlY
Oj7tXlrAKFQ0orzjwcWYgID1X7yY4IRpzl5tKn8E6JzRqReS7JM3PyKobutMsY1q
Vip+r2VDcoxKYvPhmk4tUd5b276fkayJvDyaRaXvsS82f/xpS6Zdeak/Kve5l1LU
shM8Pyj72ciiorR8PyeeI59zpuJFOATq5nwr4K5NWKdMjXwlGOPxNkq1nBdeOqiM
/0HI0Y711Zcb8gCUVenYTlmFwL0R6rtklVjr1B7V/wyTwSuCmqECyV/pmM4R6Gvl
+6rriQdgBj4Tcg+mDpKIX+Lt14KBWt2/SjWlIzxr/kXWCv5U0x7/xLZhkkq4PsbR
BvSK09ze2ppK/5h+jf5l+c2Xdx00ImU1lyWSXOpDNw3RN/+XYRlz9lwdJ4tC70SH
DZmbyLxgfZprZgU31kcSJnNzzQEaPXjw7alx4461+4J8fjuzl7GQW3XWos1uERzF
bppWlH5EmF+JKGhOvwQfabKWD9nfyk/lM4kpVWFgHe9UX05arQN1KW77RVmAEGvA
I26p58RjtaqBEmqu72JmarrF4BRQM6BydR5VSraOMvm5vNKQiK4ihR9WUa98jif3
mAlV5CAyHB5lZ/GXJJaej88kQ2m3Pmssh99vlx3VmpDW8y8fNzfQVeWFVKp8jrRL
ZHRo+J4t38DXqICctjzXM9wyj0cRaDYxQZUEzap5Rt3fd7WYYFtK+Xygfv76Ya2k
tE0uTaVHZeyc6/i9lrVnxBAWt4Gk2+tZ+k9LW6J33hN/Q7Oyf39AMsRCC0qVVkBw
RZYenG3JI5hNB+yZueGz8T1d5PmpeoBNbRU35k2ogx6WkL07rN4tUl3mR2cmkkVJ
MOBDIJfztAdKS6OJyqwH0KEoBwf4H3ifTHDNL+jkWWuVKFUpi5gjXMG1zx88pFCp
ZNPOwKdJu+OIlApWFM184oQIgdZwLRo0pbbMGLPOwZtDv07i5Qi0MQyeLT63t8UL
XgdYxvq4sxwsXMdMJpcMXT0kmTykMzoe3oJ1uDuG3PGVzHEZnBRQd7+pH41SV+Cb
SjvRF+eRWQzlmTnLs/ND0DAliwAMUZXJOP6nIMG7SulD1hvLoTBjC3atUQOm5KMS
O+wfVO8rXUT3436fxwRkjKKDwQJvjnns/8Ph7CKQCAtDoOS4zcu5uT9qpmtc24ry
JkBBCpmCLvwZX0IZBn1MbELT7YM4phN/FE/P9G4yq56M7kT6arBGe6ozen6Ipnty
O6gPX9U8LFGgcWDyc/dJcf+ItkUR0Zv9Cur9N7hOs5GDI9yQSTYQLBK8++mbazeg
LCTtBvikoDTB+MHyCgG8yPk1aJbpjg43rnz//h9FzuaQopeEzEdOP1NWgvoz9U9W
kGondmmsd0KmtaDUZUlp2Q+fUaMfZ9eQVp+UTNtlleOxNfpiSr7b82zez6ZjRCkP
GvpLzYb4iMnNKwXP/k4+TMQIp+HHHqiUNUlSl8HXyn1KfkI0tcUWGo9+qz9YbSRX
RZw4ICo/AIVfNB9Ha2yhLN217A5OBjaa3MNU8QCqzUPsnWnPHSkPnfvt2hL6lZAh
ahyluE4jDN5+oKAopfU/52na3klyYp44cPUh+fJz2CAHcWIwtZkE3T6vEaS15zw4
wW/+U3ZbpbCNG/017o41GI9Rzng0ybagJXiBaQen/WFD0PYTHkLZ7f6xktzbcXXP
3LmQ1UZKVkR9iyuQALgNmNa8VEUE8kSdlZ+StqmeMmorPyP0PYrqjbOMXzE4/ZuQ
h+fhQ/iz+KK+Hrww5Okk8mk/FICPrFlxuAzEkyuODodu9nzvIxvxLIXO/F8RSXBq
/AmZpBxfJs31kmEl8U5Be9VK11F4MWtvQ9ya4CBREdAUz+dzf68WlIyzLh2xreCN
4nQzecWhLJn3m6KOAuDxQ4ER/rgFP7wYSPGDzxoqioXYUKgyNWbaU+rGie5HVO9p
xt5WSzw9on3rBvJs8mHECtrSJJ1Ond3XAZdwyEnyYtyN4T71SvM2RTln/g9PfM8C
e7xJFiuRjqzrMzfogRvaqWYUiDMMDAVbXVHriopWQ6sjK/f4LKs6xjBVjwusy5tt
+Ij1MVvRz/W2xPAQeiAzuc/ci5xhTI3TXXnQ7U0jp2o49bzZ+YlourDuxtbLiS8W
BtxyIN1l0F8vPeDymsv07xn1qiAQOonQje//sowqMXR3CLfq13anKc4woigEXS3B
h9bt2kEvs18Min0L+acAEIz+IPc1xcUPB8aW5tFU9UdPY7uVb1LSd0BJbpClOMgA
UH8jbRVKDmiRPYDE4oEzCH0IiNTnstekoMHdZXiungvvQRxfhDPcSfU73ZsO49+a
nHBrtV406DMaVs4ffYfAUvif19MkNC5TBjtVXP6Lo2omkziSFtkpaWhRH8gSCm3M
1Ud8Of7OW5EOlm0UZpO0v3Le503LubE7dZ+osqLG9GBI6eLWQ4tfgqJE1bcxQl4S
Rk6LOzwtBUYPLK9p3jlqdK35pwYlSKYjnbWwxq+bwe3fyWBdo9G6y4PeA1TRZnqH
s/bHGiYg1gNPSoP2tPMDXmRTmaTD5uA3VExJ56rIe1A9qoaJG9+SXx8dILMBXq4A
SVs6OemBlXXlm8s/8C2RUroKunMqBgwObfj02+Nev2meRrA+7AE72WQ403FWVqBH
FIOItyazTib/7Dvnlcb3Yz5gLMuAO7u/M492eN+9WMwJbmiD0ef4O6HZOrwuKO/6
nvppk9lg9xgXejytChulcAw7rbNe6m4wTB/k0AKtPN/t2ori45WA104Zi0JSDGNL
aq4alhSb7+zoJg9CMhMrhXUkJQyqibnJSX+0whQncbilDf162lCdwDi0VSdABZMb
0DavvfpkKl7eieClVACi596f0rBohsvvyIjxMoeSXc8115ibKrU+ffAn7DEF3n97
aMw4BCkYDUV+kalVmWsZA7e64ZoUAKmPK9hsJq19p50/JqTTgaQJ9/40UWN3N1KM
e8ocyMXt6GXy/FoU1zHU5g8mxNILK86mVTppJWxJHLd/1SQXMokHY+X0kYglP1eb
AabTItd3B7CS9Gi4atV4b4s5NgcrA1ivl2JIjZYgMJsnHDNIG4KIgUJO1mVrwvRO
xxjzvZfOApU7XcX/y8BLvmBigNSWecEihljp0qReu4SkYnAdt7Oh3bR2VfjY3vi/
GnXcM3w3K8MaoiEG1vrd7dfGuxpgxzauXvGGZr7jbvx0J3Yt2kM9ldv3NxBnwcpJ
DWdDd1OqiiT81WkqPD+URz2dybUHSStiDx0Xb7CiecWJ7apaWfU+w13il4iVsMms
Xu9qPMt58clwReDrlBaHh7qJekWM17Nlrs9X/lX697cF+wqshyS8BD6Qg3Mtuwla
rRFT/vJLE8ZLwGgEKUvnBj8zkBk8fARB+it7O3+VHib2fnmlqqPYCLn3fqbjbRDU
R71eY+PJM/WKbBoIoLGMCUJM24vtdQKWy7wHQzmuqZa3jbAgqDN57ps3KYAWuepV
W72orL61R1y3yPvV3/la911sheLLngki53BG0WhkYdd4+ieL7111lrETjTAyKdXa
RoUFrWSNZ8EL2VnoVj3tUZGfcQvFV/ynPcHTkVOONTOP5QE/BW5qBhN7AcMVo/6F
9ZCtBPogEDlkXJ1ZIQltaFO+2MMG1/3KGa1P1dZ9RtwF8EymVxzU9RLLdu2r3M2O
ekxNE6Vnch2VXRy/jONT+oWyxYZFJ84yjINcmY7oUKhfAct6o+AsJYb0qlXhx6fc
7+c2ogCZ1aW3bldDTOpQ84v8HwPzUIdi2epZ5kEJXkdk5gnwJA4uwK0COxLZTfag
V+WxJULpb5HKxT/4DgTcyYl8QPbjZ69lbTaYr7iM4nIGK1ynSpN7uDch/pHu/alC
ZlNJTIfwDR+/AW6HoteWa+5H2qbQcLUFNgC/PUOlvQWRjJLshA25X1LyKaQq2KJN
qPfq1wL8y0iUaphN6biQNuVo6H0mfOjLQ8WbTAeMvzZNm4aoqYki6+LTF5sXUQ1I
qAV+OSLgWozS6vGU8+IdI3t0BMVukXIlBs6Nky84Tz3YmyhHx6yDAWWUsQZBXqPm
TgkmM0sI4PlyU9CsRB2NVvaiPu17bQOLJQaeSQKEyLTmCHi6QGWZKlZWfd50PM0t
Xd3YV3Z+RL6zJt8qxDf5M/briUlO+QQaB4yj8Pg0jK9aLSXqJxP5qU3zKnFW/jvr
h+r+NR5tYHzxfNUtlgHhbLFk8gbYxSkNX4KQiccer/WVedirBQcnsfYqwhEWvob8
KDheY0i8a2RJ8OWpN301XF9fG73uscAT8A00m3sS4m7EW2omKDtXUggeBrw4Fg3E
USv7z8kIlSZL4KX+yDGZRUjBV3D+L4+PEBjZ3rSGkTAwe+bNtht7LBKY0WTVWBzl
efuHKuticu5jSxKr/0rYlGgIFXttZ/T8aGSfq47dtylRzCiCTe8nr0ALmZnC17Bs
XsFD+8CtiqqgO7OczXn8MXKusgZHFGAr3hyqX+4ZaE6EB4YJzvM5n/Zmj9BBECSs
qvf4m7xhOnslKQI/vBqSWs9YYYnxju3soxrsnNY71hcyqxwYlOHsTSA0zHELqvNH
VKQELewI0d7BcMtgzneBa9DJHO6o3J/gV2FW424hGGHm0Do4LDjccNEkoqfCfGnv
10zi70zzkTiHRRL9ots/nknpberRoT56JAU0RXxFE+acqnzPHKVQf2FZsTHHcQVM
DZA1I73/DDiaLpFx22KXvKBbnrDoeF3X7zNxOhxSz09hZyUztWpDU0EVMvfUf7VD
4JWBd/64E1i2ihde0V6CrHCzSHoIIwDk5kxbCaIkhMlqkjA6J5ACgkvHdt783cp3
8LzfIQaj/RcrQIRevwVi1f1m2zfqgEvFi4Jf2phEvE7i/1AVZSHqyGFzFFJSt25H
hmnKIHfckzT30P6b/NP7rqAwcdtsN0QzVukfQOt4WwiMDLm3Uf+q2ZRPzwq5HlvE
rBc3xW1IlD5Z3xUNM57NhhvvdrQxYr64HcQkV64ceaJOzm+OK2bjDxq7lsKIuVKn
HXdKaGxMblbL4VCPDVf1gezddQPBjjyyftEaAeAWiwgCLcsB/iJHvFiNJ/zH1pWx
5iP3REeZ54ERr0sww4bxscE67tVcm3jdzAH1IsKcl8oJYeORd+6lXnIv490Wv7zJ
TY86XouBnTkYOkkgCib6CxHp/DvaX9uvAhmq2rRB5vRTA+7canJmOs+liq/dmO/F
Qq3f6AKxWwZJrvWpQf8Of/uum3gF7Ou28E4aiVHoFRXAIxXjy56O5h+u7eRDB/6h
AbyrbGMVglJ8MZ/8iqXvP/13HPytlmBZmsjfj7qDCAceni9Xd16uoWPVbjRb10t6
dZGOyKwtURbcFBdUzz/xVVJgKWLYe2nsNJWRT6cStxJ67F61Bl6lHhXr/c3LIPQ1
DGTW1VNpXR9l1KeB1svTBG+d99qhN1BEqa92nBW2WzDyj1LdpYdixXLqcELqOTZl
cMHg/+nB5lcKVW9qTsb0yrnzeTjo66XORDgqGevsEIftHsFPj8vXHFDzPWPY0XKG
gW3tzLBH9vOTZFqo27Xvv6yBga2Uz1BRNoMC/9Mjp/OADDB9nNM/+v454SrPdZ6A
lUElMHQYJ6S92X+dIudvsNtF/CFYcSK0AuoZiCdr6xx2w1ND8a3EZUQraThqHjzG
pK8uRhdFs1f/xLWvMW7466Dw3QOa44OTZus7ZP/fHufTxoCwgGm6d8+CjPM1PKWM
r1CNnHxau6ArQQnVYQUjvHsasOiOjSyISO1BFp/nZLDL5tb5kV+IqxSWmD7WAncD
16YEGLSBhlgLXidH34AQ9RKdjq//7RISfiKh6+bRk42oXj2YIK5b6MryziSExGe0
u9Kb2R9v4SsxItkwtYkew4hR4fdZFVWOTXp1ehtgTBi3vB+9kEoUn4glsag2gBPR
IJgGppDnxp97pWwg03lIyJvyPH9lQ7tcgRsg3tPUjxg9O++rfGlFTByRXXu0V1ov
IqlByEda/HRc7NbRunNkkHKfR7KcquQxGrWTm7wOR9pu7bujSPcMr548VtcvVx1d
Oahdy23uake0YsBlLuVGjwFSCmE0gTXXXHnUtjJlV+/SlDta49KXG+g18ryIXbUC
iT4zsuBmrvg62D03ixYgD8IeyuGuYJ088kXzyOxUf31uaki7UzN4zg4fIEOY9sO/
NK6PciKph3/tTRqDmNigfWCq+1Ygj3sn3dq9/hnP95oHD7RBkm1D/Prra210lJ2J
bp+ZiXPxdCne83rwBc6vf00gnPI9ilUwhbuJsQF41WMPyGGMA3z7SKFm8W/Enl/e
scDH40YJ1wIZsFsJeT0Wm/Ezu/911WLSJJ28oOY594c/4kDf39Bn1AmbPuSdIKlz
WZ3tRXEap5YIzPlwXYWflaEESQSyGMz/wqZ33zawJqipRunxmJYXLlXlSturkti2
k6MP5Znsc4DLoNgkfPyMWdjpZbpvLynWWfF3pIMzDcEXBe7MCKlH4kJpW+Xvko3B
qg0xkgyIevmr5YnHmJcMLdGUl+vWslz9VMz2vQ5QI3q+G4YKGBH38P5A1SgZYnIg
ldN8s7OLbReIFFkUJn19gUTRzOo68pegbYtrdaTb3mNynHW0S7KFcaxxZdQLtBb9
f7Y6B5ocwpIUL3ANYvBsGKfk/VmYvCMwE79uTHd0nDhzW/DKJlQfhdhLvyN00d9n
RHhW8HCsmLBS5u3P3RmUJ0mOkoishokhXeE6VWbEcW7Gb6pjZj4jAQkFlOLYsHUY
vVc+xe2vPyjvVNKvm/6mxcX4J12tevJLTxXEbCbgGqENdiDTz6ijMO/ddmbFI4dd
IV9B0lN3IglYJkYpc8nUX6WQDs2VjkY39vXtovrum7ioZlB653h+fySSyVn57q2K
weEI+JsfcYZ9gXKYnebQJ6VnkwIeEmDWlRI7vzdt1p+pxt6y6Pm0+8nl8ftSc9Xt
7AHWu9q8WYebhqJPhOGmuuG/1trSK+NioI7KVrP3u/yEug106PSdCpx/+TfZIG4Q
JODxBoKvesmZEGzAcyvbCblVqLsGgEId63miNRzsUx/0gANWGWF7lIlxQdDadIqQ
hyRxopcBitI2EMyxQVuUGiMoita97fFFpB+JL5NIqO/pOcEYQxP6tQ/PFZF6GS1p
3z86neKO9km1iLJgSQGHe/+lKDNp2XY1DqvcmzYjF+EagKyF3j4CL2fg8U9EWQB0
Cq4j6hZlSQIeYFo6qex1u92Kz0Fe/4Odu6Lry99c5iVsXmMUiSP4FVLgWKugwORh
Ps64mfoCpm0m0XWc8DgiV8pAtHU/cfjO/dHYU89tGMoipAVqakJPN14kjRbMTzfR
uSHtAr8POGqw4/OKSDEBxfAghWsJDHLJIONlPJ6RXMZn6/Py8nyfPrAh6l0Ugz9R
03UafCoYM0HoyZN1qOMNO9SpYjMC95k+wdfk489U53TssFsFBbUKvnQuTuJ/eW60
gnuqsx7ui8oFm3nnyhJn6RjkS1iumy2HnvH6WebSad98l5CbPraJ8UHw/7Ko1RZx
q4QFfRhF1Ihkv8KLRHYcXWThQC8NXMzS1SQlh4ACY8zA15nx7uv0bVxoEWZYr24h
xOu2XXy+EPZCjbClbUoUq6xDmx1dPen7USA8HJFASpIn/i348BcJLPNTdeawkg+K
/YtiVSN1IbzjzIGW3Nbgy64dgj9YtTCW99el5fTgWdiXZCyd0NnpojZX44yH/W/A
+WPv/DVDdWrPW3duUbGxbiz8ZAbEMoxy9RtZLrXd+ib6ju4IYbfNjF/6JtZvebwr
bSMm4THaQIY2w1DlwBNoZ42nL50ZgyFNFW01w6vUOpql1l1Zo4QTc1ANDgMP/uHB
S+1tu/QS23v0dYTyfPi+WmllLKcKoLaBZo/HrrNqkddLkKz6o6XcYx9vX7pRX2Ew
SRQkR1N7u48dn1MDLv2jmEuSmJ/3X+JOEC8Lm+0kjhkGDaWSfiRe3HKoGcVw780r
LWHD0UUODJigtU7WpYcq0Al+5RniZ5g5esG+T1WFJVLNa03/gZOv+vcza5jJBR00
eih7GL+9AQvJ0GClhgJ9VnxyA3xydb9+ZmQR6Dbrx29up4e7vAnJ7PJS+ktn8eH3
jC9WgRvFsUiRTUORh5TnNFOB+aMW9AYzgacZ/EUgsAgQ5xiVBfJZDWaywYhmZeTw
wh7JeGbPrtc1kemc3GNXIHj7jH7m6CGuZr/OhVI+gLy2Oc5lvD+wdGuZyqqnFaSP
8JZXv0vIRA1j3rhTydRxymDsagI51bGBoGAz2veyRf8YAypEO6I0C1qY5Xy2WAk7
unvZ9n2ynp7xKji1PjtJEDWiw8XJ2ZvIoJx8zELqf4C4lRpxHrOqlniLafheQAmV
CjVs9xOA/QHjH3byU6spMjhIODLhZyUTToiDVhJU8dQEoQ2N5tZSMR6jDmricKzV
BUi8ekbS6Cyqbx8igAvZrk7l2Psb6XOUFFYzjdwBruM7zC3/X4Hr5qp9SBhkU4lB
KYhsJ4FbaFvM2Lo7eIkqketerQP/7cTBBZr9kTEJrjP79hhokSReK1d8nf/DzPpN
q44He5UWDY1EgAzKQwCyS0J3fJzL77rRUs3/JHx2w+BiQoI2XHbNw5kVzP7Q0cJP
9bM2cASB1K2UdYI4jx3Yu8MWer5VGCaMvF/E4ROYBRj+8VAXYCeJxEChfhFncF3Y
VVviFegYKLB13YYAHnKO/pw5wtFjYU02bD+6kyF3rPT7MjTkhYiJcUQeYTAB2/Ey
LhaDxHFr+yBNyVEdMbS51G1IdFfnnNs3pvyJy42iHJJzK5Qt8MOfl+PDGdwWI+++
JmdZ3KPdLDLVN7igYSWIlNZBJO0/iq3B1anhWEPOuLZ3e5duLgG1pzpfUpyVXSYh
BlixcRK2GN3iXMixR+8sskg1qml7OcuZx/qVyypI+/4hjddmLcdfR3yWobEmgT9e
bxuTiTFPrYDcOmYPMAgGXYhytkGJIMAVc5LTZ24jJHmba6XUdHdxqPNRXbALyn8h
X9ANUgsVXaF0SIB+JFMr6lhi5Z7ynv8bc8AfLlRkWfpobqb5l2gJ7my5ZnXH2uNW
ON3eRpxhmHdDz/M+9GqbnmXdCeoHnXYOZC25THXaVsVVAV9gAtfi2I9Z+RsWLy//
xtEk6gS4N+495cjC+Jxie/mf9c/4x6VeydphbnQGUqpYqTEq0WniOYR+N5lYYlUq
Rk0O5pb92cmv6DzKXUNnqrW30lup6AmsDB7qDtq+t9BSylgYVvONmn3lJuJAALt3
+VO25zlODBwCCmQpDLorlzns+mB33P8GFIClHWJkykHZVQaSHPIiOR5N4FUeFCst
+vlQ8sp1JTm+XefLTltTN5sorILTqyBSjTzHxgrnLKhrnvLRbRSWIlZb/hhXfLzR
gYHhiJJ+peNrW8COhwIsXYV/VhqAZTsZo9KmpU/J8EJrvjNtuVrjadl/RJRdxeT0
SfpRI6fBacMKwVlP/0Qky8+aNAJf26+fY+xQBylsYmI+2aHUnylCH55ju84FPV4H
mFIyANVARQvMSLbDaQDrIBmEPidmB6q6MGi8kqbKbnlD/WTJnaiqkz6WUjxoSEtp
RtDIrQbiBtZ5K8LmoEOXALKLsWiUvbEhCpr01VG8DXJj5RGplr0ddifU8qb3mnES
mqhmaN/4GnKTXc+SfWbrMZnNxgeGHj9UUxYldYu8sKBJ4JBm1Q7aX0rm06QwJDA7
ajg+HqNFJ4dlqvPMUMNa1GB2edELpmULqbPhk2sUxQdsD7X41eJZY1ImfGhQ8Us3
/pQWZKMm+fy04epZLHOF+ZurnZ3MB47vleU7WI4XHEPTDW/0d/wUod3LGp+f7l1f
qhUbkQWO9Ampu723mNQjI424V/ynTKxXdhpLIif1qtiIoPE/ONAeyVunyGuzfInJ
jK2UPNcaznoEVcgwLe0C5XfEGi7DtU1klf/MptykuAV0F1XgIeoBI+/dsNbd4cqc
jLJJCLXq5LQiMsZDeIs+ULmovPYffrCk3aR5xfwHmcLzHmwSw4aIKa8HDI4sOOMs
zoBV4nMh2gp04Tqof2VmtBXLptFtpZVf6RbtPQehulDevUMRuoRnAaLa2PY1ufCm
HrwrCHQUpXq7AUWzFWh3PgGa3OdmjoRi3/sE0UWtmXDyUEkKshV6kjyvKiHaVdMZ
jbfSTKAfRP21JhDnSjXDad7lOncryEFxBxruuSz+OeK4jfVVTUg3t6cOVPgTqFh0
SyN3fQwDY/brm+4zJUXhF0Kd2nlg1TrrO09rIYmDLWU4bL8EDsjSa0HecrZb31dc
ygXafYwOXioGS4BYvtMJYInvz14lTPoQ49ZY7q+A7+ncEpr0msLh0rXt9V1hEi41
pXkL2510m1JZjAtb7G1e0yDdvhN9uKcMg2afqO6Kyjr1CILXwRkBEhm34aWwcnmQ
Gg7+Hzu6l4n8NwelloarIBkRlkaSTHqMJzMn64ek0TBZarMGEVlpm+XCiU4nJhFt
bKsrcecw6sYkgTTnEUoH+6xFcAAFxAQJtjoHiC6arahfpwsSQ8ldv5cXwC460hGb
xN7eJYXKq1LGDmzUsQhQSJ/VRHIjeYgPpGfJ9dUtTJMZ/wrRAqyuFc0Fi6BQIsGX
5w2kgz7E819LbGSyDxuMoCNixI//aacTY0zb3oscj0g1uUGDz93cr9pYtU4z45D2
HHtWmHGDxnskPdyeIPqSuVQ4TrAqhchARvg9v3K/Df99y3zfUkBJFbKoeko9F1P/
rZhkvLcTxxJU3LT+fo7E8bZAT18upKnIwyOkqZhgKl5LBa70MvGwt3q8VZUWayCk
oKQqr1U7A7TSi/ijRDT6i7+pYoaoFZ4453tRHcPxJONDk1DyiGymFECvh4wKlMm6
A9EG1+yifsCW2z6ZpaNsjKFgk7QuFmvFBfJLvy3wQLrAVkuJ4mGkS+kMuElhx5Y7
mI1Qutysq8uL4ZGBxHcpCYjhKnPhX2XCbU7AKr3AhcL8fr6vKgWaS0Dbm8IkfIks
a5IEbRxKkMi/BDQ9in3vGswr8dRTjwuYNd9USBC5IF/dX/JG3mInPAj9hplZD6G+
GLHzOm7A1bUT5GQg7LntA93HOCUujM8w17SkAtd0KX1CUFwqDhfrgEh+Z8SzOvyR
x0NK+jmVFo8rbtcFmI5aMzkpVJpPd6ShBGCIy+37UrHVYYPaxkCMvJuO5snj25h7
07ZSuYK3qNbV96IvOpTm06pnddaUmrCo7xLmr0dTigIpT+eSAl1M8rFpBIibPtN7
3xem07yTOVhurMuZCMWOYujtkH/KLgzhrEZfy53gbHrJ4mB8Z7mt4IIdAVM900Lz
wjeZJiyqftu38B1MVn1y8Q6DWjyqS8YDxFBLxuNZZ2+0jh9+ljyzgvFN1MQmuKG4
98b/DV2ApK1/W5pnkHyG5qOJkRhbONeoch4S+lxMemi5Nt7e358QRnWkoS/lWuVF
d1XaifakRU94sg/kgQQri2B346kfVp8njSl6Svgz2GHpvIRSSce8ysPB2TkCpo8n
dRzyJeLTfas/l8s4XN9dQDuBq/GosW7VxUD8ijhU3B0+4ptihcFt/hHkAEm4XWmB
6tl23SjngCjBAIXA4/l21uBcZtW9hQQabwf61Hr7W7c5gF/P9qZb4WKdgPtsUmQR
i2UZTDQZws2fe0sKSEpnMFELbhS2EF6aKVI0KYbiSp++dT+dTwJWfyzNQtSeMq9O
o+w3O9jP5vCs64HKmu/AKuBbMjDQ/dukxMP1jHOtGF3j5lJvsBwYdWaiQ4c+dS+P
fz6jZ8RXiZwQRchD4ve/MDvn/sUL1jKKKuCfMP10/0iE+5bUFFVuoEIi30CSJqLg
7sJw5la+np/YyAQfAPMKfMygKMSNPBre5zsrCWggeUA5n+w5HP4thH2LJwZimvP4
ndBSNBF/YHoQTckNYr21PcRP8y5XFpQDh4zTSITjIWsS9iqWcXCnZsGxOh5eq5wR
1hNvCpoSFosuF8wX12ebyFPgm/vqQCDcD85d4MEM7BKc4CBdX3taJj2LpoNPkHO6
HFvqWALtk83M8iolMRqSx4kLe2ckUF8xa3inkIFnVkJfy4mLsP70fgk1TK2Z393M
hFbpdRWq/5DLnBmeNac06bphcY24hapnZ0N9pJnHBUvSiWpXwdX5UcI9ESPSycxZ
b4HPYfNZZ5TnC3tPDqyPHa5B7k2NSfpRf46FHSqvC1Lky7/GdYt+sP4jxeR/gFSu
9CsIrtlGi5hj6Yok8Tg8MkT5S15aX9mttNZDsqqcGYVKVva+e89E+UrZJs2DTxC5
zhearHnwLZydfoMYIQIBBRswOTDl2L2Q/o4Z8dDPuAebnD0BC5jwTC1FmAmggaCQ
IkKkU/NSjlLkN4weVciGRyquaEpQ1qKYtqVAtxahHLwi+8PsBDriemNsGiUKWi+X
oj3GnPVHDQXkkO1YYIrqiX/Ph4jaTmGhn/J3CC0medi/0Mj7R0BCOXBMg8hL47uv
x1v79fvN9eWVTR7wzuPg6n7T6Nl0BNBRyXpDZ2U38p88atvPDZG+qIW92tvnWEEB
M0DQJW/VQM7d6PSaSISd/+UafI3Ux4o4S7ch4/llK7m6vINZVV+fBZmRf/WsdtlH
5dLdbYcKSZY69Q/LI0t+OlHmR6wkYPsAiQsdtXOcb0LYwoOonckJq9BEtGL9R/p2
XJM00R9ixVz5YDe3TDiCx/LTg8HsW1lqQ1g3qfc1ay6IYCV0XRGi73PRC6n7qYZy
NIX0n5xMg+kc6oXWnWR0pLZBYBrAhHQ3vhSXLDXX3fFk7K3TpplAW86SdZN9V2nJ
887n6L/LhpI7SD9Z6ts2y+gqkP0PAKMy0fwp8x2mj3OdQ36+cgIGAPlKWxa3qowq
GEiSLXLU8FwLQVA6yIcz4thNGsNlEU3b1jPfJxb9NfRrDmXrC7maEPR9qNdpxoOh
gZqk9C43tjqtDZfxT5SyVhSyT4Dtu2vxk36dIWYp4wv+psI8jKQVqdOfCQoOIQ0y
i3xQynlgG5NVwZoHwWuVy7kLKeCUa6LmnSbm+1AoAJ3O8OVKwdFlh+JBeMqjZjFm
erqT31TKLOyGbpLsFZYY+CQIhR0ifwEO904tIqz7qgEcbFCiRfVEcPDcE/yrEXAG
UL5WAC5Jl98NEV5AQc/pGO/T2w7cealMqucCF8pzvAqMdKH/5Er4BRKVkgEXGRmD
uaYVBreNfpY4q5ar4D97hmjm0n2poGOqEXW+ll9HdMa0+AhiYTxj6dG7TrjRdJt1
3N0GzvrKrPN2pQQECxBU5ooxkqIRYEnxNXivYw6awwMbDxETtGnE+AYGtbzD+hQf
/1R3tGDZCJTt1chssv+9XQWD/9+CSaJBXUkFJlTCmNGKh1jHCqqeuuzOG59Nqc4i
9b2+ALCxwt8eK6YqWT6pqnEJhyoaF+DTBtC/xUXswiIhN5wGyMg49AI2SPF6rhv9
dcLuDg1CV381fQE/NMC/QKnLgvkw+Dvr0YFLmuq4WiWJAunfBiK74r94sW0fWN7C
1j/bXTaVShAIADcbevd1p48KLv96os3xSeD7AAnbIrULgT5eDNpkbj+Kf5V856uX
wAa+Y4gnIMMBEHc42d2w7X9b2Na7XpRy5k5VIwG9s3K+uEOVsvbXDbmIS/1uQF5j
GheoU8NuGX4jP7wFwp5eJYyju3P5D0bM9oNQzXUnbeZJlE8qpBLYtmeXk7xQvAvI
e8Ck47Zs6VJMEzWnEw2HOoF9AIYCR5jVxFYT4r51ajCBczS+b/wvPFFtj2lECmof
S4koYvaWRkRrqV0Nm55tTLFtMYEOx91F96su/UiMj9tcGfXYBw9dQmsTDNcNMwgx
O7dmcd9KyDgTlvPJkxVrURp4Rl5Qm53CiziTi3IMiOxCOYJeL+bMeKQ3g3k7WeyU
u5dqYdL6FzHY9mPq507gPqR++FBk1CTcU9NxKOflflEw8hzXPkPXkjH1Tx1LVeKp
WTn/W8gP0l68mzWI2iD2uL1cdfF9aOi7cLj3B5674O8Mr32mOQNE05tj01dKgJz5
p8IbdNlJdsnrbMghWDwxdWK2ssi01luRiYgJq7sGhjkSv6xsKjz3i036unaJFiJt
IxLn9vWvVLHJ0gqCVtDyiml1zR++PzCZ+URn+0G5xBKTS3UGht1mN3nmN+goe8mA
ptZnq8Tk/+HJkrCWjUWr5eLz6xGbs8rv2DB1Y8NyNsNHcb+59VEoWJYCudjzPk7a
R2NERCO13+7qgS0frVfGFyT3mDrieZWQPKSrj6P30ctxdXcY/XuH5rEI9FL987v9
bKTqAchF3sEkNxxpeXiQDZ92W8Itx9/mkhvacgKL6NjEDLS0upN/Fk6+cHNE1QFm
9E2xLqEix+XDzIQobqbztlljIaFgm7X7cb9rNs5oHaYnmWBM57kMIBdENoMwL2Vd
1TWlgM1nQuCXEtZwBPwJEMMWaYLdGfZLkpH1i+DnveJiTJXOwiR/RB/IFlWrEeFD
pZ9pl3D9Lb6B2z6Ue2S+7Ns5ANR60XwoskNR/5I/EcuYokGmzqyid0nwMfhLPKaH
LNXD0tvdDEiiot94vJPHYXZ1gPyvHwuavddoickUQ93dnkcg/k2avzLhnN3ipQZM
QbYPYqYUtodC4Kbe8PzIsOKKGQS+ixcVez+kdc7uAwlTgFSUhMUQEcrCSzf8IMVr
6pmTwObFcNhMrYhRcu9jMhf2iAf2wqCXeFn2uP7VLqDI0YfbMFnTzdCVwVfyFIAm
yVHBf9RBfe18ty8DDHuAz4odkepWOKwc4T2wDxbcDMRPx1hll3pXW/JKwjDSuNgA
LWGfogSkWsuRddAl8MWRin2dvkID5RLxLitImqCl9fh5HOexfXqjwndxi+FokTPb
qAM7PYUWgegeOU7kjvypGwpxuwnYXObMWgmQlo5RM47Qy3BZnJXCor3aaPLW1fQs
AMe8RPMsmkjcdv64Ak5Vg4x4mJzXQg30YR2kW4977huDUK2zndMXgb5L4Ch9ln/A
87Ow30b7cKVnib5TP8i/UtKsgzLt22ELhiNp+U9BU2ZtGMiIs0SeXA3aX3xJDnKd
QaGTsMYypzPRh77a5/aq6wKtpPquXPDOGWCS7nFudJhbPm9GI8kloJd0KI5m1fxI
D6TGmqErmhxrNH1KW7SdGhh5N6VyBwkRtHyf2TWfXKOzbt2Sxf+JhPP7GMap7IYr
La2fZXdgvn3lb/F/Hq70V8lGZ/xHUfWscvOgnM+kQawJnkr2QO/zxSeL+0rj7Mwh
izqv/21H8nhAf367CsuNdDIRAYsDPFfjdaEQAjWR6ocxwjZPBq+I+02IFflWehD9
5drPTaHxtSQrOgPspSSDkTAIIdis1V6Qb4cr96Yei19omW+YrnGGEam+kkRn7S8L
N1C0l3dYXBxAqDNJ8i5L/ELCGfGaB9EQggkPSys4zzU7Q2CSbq5B9Sd/d6ATQqG4
yV2w/jYK3rvQD7WL/GIFz9YzAyNeHCC2eF9IaIeDuEaXQqFla11uqgo5hbtl5AGx
byPBhkuCZp4uIxjFzGy/IZ2+C2AStbj7YFjFrX8qCyj1lHc4CfKQmkmtH0KuToES
x6oqlbIGnZkF02zPxZkAY2KMz8/eDce+EY97RT0uS2BpNUgpeTqFR6nknpZHX6HV
wjdSGSKwfHZV4xajpdMp66eoR23g3Zy76ogs6NFc5gG7w+T8yej8k30aMyOZLHRM
DFP9lP/KIIGyHeQMMbnxRbawrHalUnlGBcDy9ZBAkVBymyjmfPuhCqHQww9vUzFf
3d1l/T+l8HuRhgn/F/cOuf0CMmMssRhwG1/TvXa6UTTWEUi9AZqW1cewSqhaP0AI
ocq6eHsuL3BPNCC6kzSM055N8Rvqk10MVzBv7KoM4OxYT5XjeWx27yjKmK5M71IV
xo06y/GTbC9mSEhNRlcHkIm4KFD2TQmcvD+EK8tdyC3et4BM/c2YDtgplzSeeDr8
0tkMdVNWp+FfmF2KlaDc/boWcd4KaoJMIWKUsL0ShcDlLhPvlMbkhofwj67uArhK
xTfIUuNQsi3BxfxqXgLYBZCvvu7zEWD0wDqNKhzXZYMdsxWOpZtguAD55lerKOwQ
mByTnMylAE+LSK+FG+ZxXXwuPCVDADVAEmHxQgLVhiW1jepKdMUcF3YiCfq6IAok
sUZyJFOLGboKhAtApAghHfFULjtf28f1oKxU5ELKuXCWzsbwn9XXGbGCpewrHhoO
F7yztSsdLWw9s6ZFQ0rGTfPvn2+a034UNfTBEK46mjHflCTY2KNuFuUJWj02H4Zk
GEaLPvMrpUb3JgdBNsOqJqb5ETV9hjc4UEnKh/Go8kbEWjJeTj20GiPk9HTPQoet
nqwzVMoflHJlHVwGsrykFhvOmTr1nwmBZ1TRBH3tLhdjxU5LHubjUlh0tU8PhMdr
iv24myw20pp1ghSrVcevCwnH/H8Q1sMAKygqjWuD4HuiL+H+XRZMt9eh4vayFDXv
GAJQx9bCm4p13vCBCDv/9woRsBrXIE/0AE0sLGYIBeQMzswiHmZRdEpeLvmt/zeH
/eKpI2v6N0fTY+7Ntv9S6y8c1dkPEKbJ7g7U7vzGdl9Y5qU6wHye4TI+NrJMp5AZ
vfe9ZCguBC4BsC08BfBvyHw/HEz844g4OoocSk8BRWyEpQq3X6OV/JCuF/tKP765
RLvi9G3pK6bwSCruRtexkz0h3OZasdo7Y+x/hsifG/dVHPvHk9u6/gFV6wgd1NeP
PiXLyeb3zZYEhorKBV+0eD6MMS/26jfdO3Kht7glMgwDCudMpnR5pGPVml5F2wrA
ZF5/NaxIvs0RY8UeyXONKnNXHuELxHZx6swQjcZIk2lmAXXfzlx0TxzaVbzMM9vO
uO55F0FcknV/WzgOCuTpygGDSKwA+A2SAO/J1bqIXf6V+4yfm4D9iz/h1tp7/sCO
TgIrRdMGymQ3onj45keGe5wa6Us6PPRU5W5TQ2wEn7UGqeKZeL8fSOe6hSwaLIz1
27Ward4t99BOPbbj6SplL/nfx/V03nx7cBT0BEAsNVxE/+iJxSWjNpIBmUAWsWAt
gvhRIvqT2Fo7umM4LTAskrZmcfx79se6lv0anB0QrBWhok1BkozeOxcXUy5sOET2
D+f8gZKomnT64RCMctN+jZzLO9UyqlVyKhFc4RFeoGVzOXVyvv67WcMatul/t6MK
6CmKeNJYkSHhkb3oFtSK3j8o243RhNWsapNHZdZhtl+CR5vg96F0pLTnHyCrDTbw
L06RlDKzM4dHr6s78/TcNgCyCJJC0AwATsicWMBEa2enrrOsGvCnnKQx8ZS5q/Og
TlOB7H0lUz9vH/F7vduGh2X6cM5zqfT5H95i8dzIFyK+T+MImcb1GgsnE0bPXCBL
bfx5paOSxGphFPFQQVOhrYLVl9FCYnD6M3qeeRjIQ7JfoPuS4vI+ViH6v0SBxJwv
RdXYSCLiWAHNt7B+pzzkynqLuJzJNlaYrPJ+wT5yXX+fVgfj0HHkdRCgPYbAiaqz
ILLUrw66ZUQYyseuMcm2cPepj9LPIaQgR8k6dMFUOoh4UNqzIzDFc5AywHqipBoH
0ATuwHZVO5A7D1YvtcwNZaKaAVhEb4CYFNPM2VYcYZy1mqh+zum0lP25RvxYiPVL
ZGUIvJkoj6xkjbioKea/bfzU+FB/Ngk348gli6qNBhu6GlpIKfbVLiQtL2BU/0Wh
UspVpr2XmaIbap+Jiw6dWFeCBvzg+DQcNo/yc6KpwG44FUnrzdLhFhxKqO+aK7XH
QSYC9v0/DXqgYAIS7LMIk5cOKBbibRFgD96fDVEORsbQLXiCCw5osUXDGG18PUVR
XoFAk93mqFpn1IxCNbEJNLGlQLju3dsfPsPdjTooflevkxyd0LFKE87iAXdOgOM3
hreXKOKtOKp0Ydvk1h1if9vB1zlRnuxc9tJ11rRhuhYdfcUDSdR4xqXllBD3lN+z
R/Hpf3GrDvfL7xyoX0UzctGgF7lQXBDhU5DyNhA6nz2yKSPVKAd9bkI43Rbjkr+4
Nz8igLw0xOdBN7iU+bOkkrJPFIAp9UkvCOwdgXHlhs3+7igB+USPyvBij0iDCHea
+N67cYZUz4MB4EL9tP9cdQmQO4b0QptRWUQJC5B5MpebGjqRzE9H+7bcHkJ+ewgr
ywl/fvqSdUC4ulsIvsmIX8liZmXA2eRkoH7QqO/k9TXc60rA9Qni1npcDYj3RC1D
hYN85vc1enQsinvIoCFObVZrIyFxfhtBUGHdpfOL+wpsYtu6v5Nm0NzeBMxvkMj1
gJGkBGjxE5+BCk6X02Kq6tLZKmUxhT29YdBvVvPd8dyNsRoquHkMe52JDga9VsT6
phFkNtfesvLVi+kbQhCd4c/tk4SerjuWFucF1V8QfByE9ziV6XqD1s7iy4KFIWIH
/cYQlXwD6+W87FeLLFzxC+L0pgcRYVatQUZ7M5PvNe7Vj0fFTadLwciUCRnacLvJ
9Ah/8/UgnEg9rb1inbfVG0kH+qBgLANbkHZ3YUM7jxKNz3ME93A38rmjRJ/+VrwX
QmiJL36Nfy5JC6/Om+wql2y3qYQ9lfvH4hHy4C/rEbyekgAjW5gKP8vqW/AEs9BO
7IOB9GmLGrWIKAJ2PmTtuAuVEyQ0TakU6WwHyZ/5EKIyGo/2D49G9O31kq72JUQE
MJdZAAmZV8NIhFzEpzB7WWDngtG/oMMC0Ei6Q5O8bt+bmg3aN5afkvfjVA6lI61S
NxGiFBGC6u1mKxUL56TdD/rNq2pmpgnJ7sBHjcuDloS3XxaNMmGsSHp45xnzZjNJ
EGZU81BpMTN4x/nVPIQYARGnoA3V1d4xiYHkdJ2TTSHnBalZV8J87mmdQUW3JtKd
nNb8gR0hzfrKIctaKxkisd69w5iNXE2IkV69+oEx4/qvCMqk46dHm7hD5+2LvCbf
sLK15WFB3LC7dH23368NA1lfswOClmc4eK44sTVzSG4aWynpEjJx4n6mZIQUeyyC
u7Jr8F2OrmP50vDot9AH90QyoARDwrdAkahBBB3WVb58YAXjrtuP96FZSQ6V1GCp
GbIVw6a6Op4jX/o5emCqXjucpP4HbUviUTYerNRt5Ijf+izxfThvEHb4MVtQbGrk
OfC+napATXelMLXfy6mpIFbDSNAqzUzA2eK8E/mCiDTVxIdfTZ7xNQB0RX1k8Iih
TIjCvYDDuRstIEKRx9yj4d4ZPP62R3Dzq3gYI1w1a4IYam+JUHkmiqI3hSH45tth
ClX2MdnrRfkA8CX6d6bTv+hz9MCUbD3kNgjC6MJqIutVtPt9tQ11xTniSULstgm5
HWjGOc7sYpsNI9jpnef/2qMYV3wLGtf7p3UmolNmVGlZ+kCRgOn223I2g67CuJsk
ty4zqOON6yg93nGwxajRtQat8Gulvi14ASFNaGpcNCVvfP5x169ftkKjoE4DswG6
GWsGWmwu7ZqRTWC7Ud6ztfaUzQPoYRFAAu82G7sOxHAtxL8D3CEGQQvtHLBv/XG1
jSr9T5AgDO+gRAEgfbM6hgbQR0fjDycx+1atY7ZzFcd01znYVBFBk9ZcQaiu8PFN
bbtSUB0DdvrdFeqvmY2q/FyWQCQY7JvSilp5wIXvCn3Rw2SioBhIYGk2lkwuyqGp
oBMtpE/331Csjt31ICCu7fiO0bGrGCXY8lF83fnIqCrqF4sceyg9BhZjbIMGWXES
ULPlhPMCnE3OVaz/Cj8O4jdsOHheOh5Q4aM2AWmoyJsYnGTDBBCAVtpMiVNS1JR5
15K2jep2pXWsrmXek45xFgmfWdkZkCy3JN5yKA2ytCSAS14kP5HpCCdUjBtTIW6F
xidSUVe+1+7sWqait73XYuZIyzSlT+fYYyzToB3sCFplgZ2ph0K6TMRck+ivw8GZ
iIMxKaUaDugwle81xn2x760DXOpcGWTm6IjTTIV40kyrlPXYQZwpFiVPQapJxhXq
shVVjsvy/GZDKYRjqhczCQE0ALg4bFLFJ79/BYb6D+KQz1zctiyiVVp6/YA0fKtF
EenzErqE79eSsvzSY3XCrnbWaTexMT7gQ3WjE0aU8JjiEYJM6ZMAen6fmq1E5JFe
9HrSRbP6RViS7bDdrsaPuQO369dPpfuPAsp17vjV3jKRGbblrlDZ4EZ2TsVWnnp7
0nTmltQpMiVHRma+XjHWickcKbW8WMDnCQzoOgtiwt6jpEr4mg4J/JbNuumrBZMC
PwAWNZILQ5ftn8eSkQwdO/z62hQeFz4t+yv0aTmx4FJf4XtL35dLiLya5OybWloa
+drEqL15hG2V0fkYZRBBylXxGPvGOwIWosdM3i3Jfs8OtoVw8ZE2leTHr8vRNzSe
N/V5y4aCqC7qE411qM+oKDIT+V/Jme77UY4a+wkOEKmaUp0r51ZLnn6AV2IukwdN
mxmtsyir2+JCYiluX1lysDpuBF5hUQTKXRC4szRSNvId+Wncf1EoHT/hNu/pEXft
M+atZ9/Q80dAjAHutUkFfRiM2bVf1v8Xf3nmXAt8gKj5vDkmT9Wnyp+qaHplC//a
aO/1S25OPQG4RXicxEWgY8Mfe9lADMmNcgWXXtgDsPiiZQAbq2mwcLZ4w/twAt8F
Ynce7k1Vck0i6JQaGY1GBCp19zdg3Evvg2gpaDYnPNiN2E+V9lhqD2dJ9RFeyIda
aHtMfdB4xWiru7YRBq2+AWVpSMAiufyd886iS89Xl9OMr8vBi8zkPlETKw3TpkHq
jiPcQjPhXfYBKPH8xm7MpQKgqod5fbMGitsev9iI4lTILmauootvCO6KysP8CnRv
Qv5CII4fnxVzuhP8HW9HNtv2nWmZXNBO7+owTdwbtM5Mt9p2KpEGuU9tM3CRdJoz
8tDi/A31gdvYRM6zVKM0xvtpOkhF+gFj3JU6oaP1aKGvL8KOisNEmaei8NN8XEya
V/W37Y+o5JZN8BnQpUfwrak9DvvAjvmMmD5nzMtNBrhuJLCMErX/yY4Mv09mnij5
+hZextj7CTvWNodeyQnteVLMZVXPOChzNL7Nnaof+h21bD3txugMl6rEM7sAj6PD
tvj1yy54teDAkJfwQK0yIv6DjSgTkvZKsGMTT/Dt8B6CQiZ/I+wgZSdJ9ESrR3UF
CWCO4kWLFh393uyAUvLx0Xn7W4SkT/+n/qQR/Q2JVl5K2DNYiSDIGFdjdXEp2XGq
cBaqGtnEyOw03sYlRR+R7gUuQdqYNYdIcrueNG9kwXQ3TOGYqJhuBIq9PeYr/YJz
DHJaywsfAkhg0CoPotcafi1j+FWmocdlsoLV3pxP8wbZ4gbM1xJ1fVotf+CdUn9s
xmLdMf2X3zW6RJfdEM2bDtFYl/onpAEiN7HypaQOnuUdzSZwcacywusTyu0tJgsh
Otndvg9l2i46hIp/1e3NtXCEYIypVSQB/jtfFLxPFGX/g6YOFyuwsgk8rVaXsTTn
VIiCXH9gRf3ymORXpjCIhUVGubQ/9p/c4rF1u8xbcn+KzSkELzj+KoXR301ZbknJ
iHSA8+MilX1M0IGgi8DsjNz8pJ5A8N48hKpB78kjgbQSzNDljFo72EWaslAhnmzt
07iqyPaR0wLuv1q3MAmoN4ur1XdPvTbpjyNUVaYCTL2QaCmbB199VdPnSgTUNyQ3
BpfI5XnW5F9oi8eVQKV8JHqkHZTNouiEfgIs+XT2PjRJwYu5C6cJ/xEbINcogq3C
nkLBVi29x/6XjlHw01TwPzAF6s3nFbbHrLl/WMFkAo+LnoyrGYaZKBFbmTbQfKCW
R4834NhkxM0jfskPC4hKNYq19UiIb9kmVvs0AeLXqe+1A0BuO9IGOzgmERF/3jUP
mi44Ytc/xRhciv2QuerZT2ZlyzTW8uxoBidUWr/jnH1xMSeq6N+n5iLg7wdOPTiq
8rmbc7CGSACHjMsc/k/wTCQdV6VdUAPqdGs+OmdMwC47Vb8omUV1N/AZsQaWrjcR
GOHWbO5RfPbgw4H15hrO8iyC6gjgizEzoJnmz24V1kSCe2YorDB6j1KTH2poA8vE
7kfmwJCcEgcA7f07bfZV92s6AURA5kOpI3pXkru0w52p+4m7adGj7ivzSQTkqOSY
UThDC8qdaBohyEIumDLjFTPfeL6HYo9gXhbFdyMoN2X4gZqc3gSKePlabGBZMc3W
Id3Ymsv767cUKaaiC0+S1fUiP1hrio6pmgYjCtLfjqd+D9aYPXkmceQgjI+6LlpN
gtrUdujxWUqkXohzz2Y+vf0UHlUa3Wug5RIr4S/hOStTwVz+p+jlcBb6HnfRKc5J
UZel1iEJZmfTgxyhtQofKoAQHYlAAAVF8gi/uoBJeOI3pYLxAOEVkOIsgwkVbBbF
OEpQaDIDrVPFBmgCyBukujtMBupi9bQ+z34aMH4nys+PMzO7EzCmqYxJjmltsIMG
qyOpnKg2u6HcMJjLXIIQpYpbUsgOQULSEaRFJy9bmFu1cSesi79sgBWuyZqRpDIc
RRJc3297ijIL831TcioVD7JONzMLqx7T2qLqHaq4S4RUu8z+H8cz6r4URujEr0Il
apn9D2pGKmE7tNyTLgyZ79rA+HmEHe1ZG6iUf6XsXnRaU8jGuRDck3hPpfKstF61
lNSo3BXbRx2B8898Uum0tgKBJAm5MohvQOzLav3ZxSYwl8Oxm+NC+E34AFWPAihc
OZH/DgSdG4AAi9FL0c3xgIewKsCEKuLpt7xAuj4J8lJ7PIAAhHG4qhR/HOsG9nsC
OtiOYAnOgtHaxt5iiClmkOSavaY5BLXDkP9VRuVoHxc7f8wHv1ZM+QlHRvTogWoX
zV05jpaTXtABrY6rj7CMuCkEebd9EsbO3WVBKKGnxfMtCNLGBx7ya7tf9qlEMCza
TXXFajWPqTEE04molTkhXnzKJuUn1sC7qV/DruaGmGYfbHc4sLuypWROX5ThECGi
PU/8CwC9mUH3W656S4lQU/H65zAHwgPnokvDHkd0Eb5/z5V7kLLTpszN2cJ1FPAS
QDhcBX0qPYBPx5dBGpdjegB1Em4RtKNy0+ullOEi/UUORW969FRzOsvHvRrOftMC
7XDVXqPihbCNiIf9WyX2ojGeCEyK6q8rAgxnbAzqGa8pb5kltu5Ga/prB1lFS1lR
/vsLmC4phaUTz4PWcFWimxPqUoSnGxIwNibgnWk5qK1s3ZniqGr+4VVRp8WoI9Dm
b7OmJ5ex4CUPSrr6amJEMR3TMyECkAB3nx7P0OwqXUewjguvCNaApAWHdjB6iq/W
kzAaDro8BHzIEnmI3sbultwP27SlaZuOpm+wJxUgIupRL0Uf8dAoNTKszceR9Thc
9VRR3tWgicI06xnTxq70NKbezZ0r7qyH0FtwNExgeFPzJOOZ5itKHfpkDk+4sNqN
8zI/ENH3GsQbovS/DZpXnNfWhBhCwnNSIatl4iizm1sr9jofCJR27PZarUiOjwfs
Jm+7qF6iDCga6OwGMMlriau0jIgKjq32Nsf5/gifjAXpUiGJoLgWWiE15vi/JRGf
sjouiRhFzWiVVHQYCUV0yePZOCkvOqga2YagP3H9YdnS3d0GWWeA+GGAyFUXc6+R
WkZpsgIIALEWsiTbvVznU6cXis1XX99TiD93DpS2NRyX8Dafsw820FREJuEJ0Jbi
4QifrknPR8cNPPv9nFsz54juTy9d6NSup0naZbx/43xdYTz6Jt8OiDJZ2QUquKJ2
ic5AJvfuEkd/DLXUdzst7epoIi7zoTAG7n5amd4fS+Iqa/WUFmgYrhvYvAxofpjh
077Krr03GbMfVu68mkgf2jMuJedQah2O9TlZWSjkxgOJJAc1y8Kkv3zTrqx6PERA
dns1TpJIpOszemE20Pg9KXxGny4bYjUlA0nVfGDuIOhYy8tmg76zEkQMCmQRZcmR
jqP66z4oOlYmCdQvEU/vOF3EJL+mzdWe4WUCar9HzHhIBYYKTgIrcjd2YVoKc+vH
adPGKGf1LKtKbTuLUlg2b49bRmrBR6d0LEfVZrisH35o2xEEevE3hWtMw3od/2VC
1go7jO5HN8dEyEKsmKG8Aoiidol9Dlisciq8pxB85Eo6Rgx5sgMX0fERRBezh6Fn
NcWbLB4T29ZCopIuiKjOtWA12O3LrvrgarTetkMO8lmehTsIg0yTa4jQgUS/lhjw
ZKH1yDcKyKHDQdMR5rpIpfPVwujgiew6/tfN/JFumYaupIOZMBAr+hzxtRURr/Q5
XolNJ4DqPeJ1xCX2P5JKzKe4BjZoRlqRMXIk8DFYAEPeWm6eMyGf9mHSDZMlT11Y
zewRf0TdBKWb31bssSOYymLBgLxL/+y7oIEfv52Vw8eTYSLcH50qXMjQgdkGnM/d
jAwfmZSNx86msGhuptVwOwMh8ntXTcT9sj8VEu1AjlYveNdZRHqTBZv1ctQg30Bx
3puFEqcxAaHiz1EF9Rb3/GwNucIsr+pm/dPnfrf+5hcB8gWLIfWn3WVtDSrcM8mT
CutE49yvKT+/jZsJeO0KrFxYQumT7SOj0znZp/R3PpHcDK9fPCYG3Q/DEtaFFZFs
I9AaxbRa/DYXqSGZbRuVV51kuulC0lMin+CnnVYFahps+Cah1zkdPffuKflRlDFn
G07Qmb/qGS9fNPmPBDTYfuyDai4rHZLakQIer5Ewcl44Wl6Rz+w/4fwNrzLrqH/z
thaZ0gLKdfIUl1hAMyK6t9rkQGsXqKsWYEEFw6DqPGNiDyQm0Mg+Ya54f8BqiEfi
BbnPB+8XcmRiVyJTWYNHfDs5IDUfZ7ByMuNdLNoHKkEf0z3/vgziesdJP0JInaWm
damnpfJ1AteZpT0+oG137c7sw6uHhuu4zEe9T4uHbGZMNdr+SB05EGFdOndZtJ+g
5ex07wuzx0za2VNKBQj8JseR8J0V9pTKPrrjBtWuUUgEBiWqs7ekndmH8T27NVGm
mgi5QWFsi8sNh70kJnQri0EZ5HITWAmFfkVTs2MnmLICGj1nMqCrgcC1Mjvr7WMi
p6yNYQiDsN32INRWUHgkJoj0iy5PN4IS5NkXhQE8QnHqak6rnPNDch7Vn0TGWAmg
sD717VkMZSo+WBkSK2BQZ08iLBvIwEfaKN1VogOyZ/R/Fpk0M3ECUUNcWcChBFKO
abuSVAk/hp6xzlekKfFFcz7bUTQPJjSGt8OwDBkKMOn0n5cF8301jIfdNUHX0XEV
S8mxc7to7ZsHka1TTYlbGJMTxa1jQptQxE1Tu2LQJesxoo3SosAF2HjMjT5xpNjV
JMe+NIvscQhsGkyrGS01AexG/u+8Dyq1HWGTRfVrIZhq+6LctD1wKy53sdubWOGg
KX4Z4HJXFuj90ylmHd6TltGrXyhzZkd41rwIcQgFCYQNARvjk2W8LTLZ9bYPTdoz
wNmYpqeu2ehy2TwUlbkjPqPwOL71qMh+TAEXocpqnGhynCqGYlXK6wJLKvX0gTWc
+qhd//6WbmO2LOfMxZR37+M1a9lgubv8apn6lniJtjobnFnVqbJ9sWDDN6YQxvS9
z4OVm9z0McVbip6kDZtsKK7HfMUfPVB3xf5G3aZAuIpQWE4a2fGNMtMb7iG/6chn
LJclA4RSU8EEw6vprrsIAqlbsJdJjRriesZrKWaqLERLVGr0sx5CfXsz7hR52cXN
3pWgY3FcISe53WaVaCikdoSAXVpi6tfMJdyMMHz8v8QP9QofsEGssE3RbTiN15S1
yDkZR6F4Fls2AWl9SMSBTeMB24rMFHn9Msrtp9cVpsbo8oa6txUt5m+YW48HyTct
0MfJ82OYnqrfWbU8vJE9rWoecx8eFFOJJ3TgQne0jvEZ9Q5z1MkZO7B7W9eyWDvv
VPotB78XC7cxJsco6wuXdbAt7AfolS2T2JaeBXvTmWH4nKMpFbTGSaMewo5nGV2N
bd1ss0s/phpboCp3+g2bhFKw5jjrasot5YgQGARoZ8iYRBQXq1tKAF3G/5Flykmw
QLtcvb5jD4GaXQWjOPHlkn5xgrTt9e+DI7hNydtf5+jIaPC7B47abzrbu2eefxF5
EpvZxVUND32M3gSV/AMY0vmg0xwJ65gzIqG3JE/zyTrUziy1hJAgks2j2iOr8CjF
BjUl00VNqnCAenScXrKpWYH4/LTeHeaHRcIpr5Lr0MAnTJIN0H9QQY9u1RIZqCDq
PeFqldcsHUlqc1jVqIuOQ0PUfufvjivHGlzGBgnN4eBTk3tTmHp3sbcOM/kElSuP
ncs/hTp1Uctm9oYzpYG/0jZS6M/aPRU78n9RADjHcx6Z2ioKtEjcGOCAh9vkW3hH
kfMAWLpsxUhUJpegwxfnEHKHuvI8qPxM8iV9Dr3Mju1K6gK7UvbZ//0jCuwvtDeS
fs1Ns/SNfBTdwtmr670z2Eq5EV3kM8Ef/WGUUAGi3xEZ2wpi6nl2bTRD6iGHpdUg
dpfeaHOX80O/mpPIkCQjVrfowJdIqi5C69VkYSUNi0ysYcz1b8EyPg9c/h8P5sW9
Mpg3fi70EpuXIqXPpdI2qmbdyqOr6bR4NXKsK1K8K2TxTztpwnpb7O6GzSCv8BaW
lGEFzcEsciYhBHbDuZ74h4A/b2IQAPUWqiPW5Bw00XhGCKvsUQj18Q1MU2zxmXp1
/jxKy/XK/4Yt7PufY1cEG9gsygxlN7AoKt2WtYg9a6qMWjyDyQoEu6O0UV5p0Ynm
6sfEa0d5Cl2Ka2bGQQT3BAz4WKgxvCcELwonG8eskTofYeuSUgS/S54mgzu1lrZO
j/fpv+TsyBRrreUzumSCyF4N9zeMiWUZk6TNLc42ugsJYyJfltFBG/EKHvSYpuVa
kppWzY2NsSSzNjZKZ0viQKvnLpFhwRa/QZeEnqGbsGpaYUnAg1yD609nVMvn5nVT
w28ep4KbYcGiPBgwEeGjn12txcSJNckH0dEIFRh9gCJO97UVQ7qqik2KxL7Ml4NY
YMW/ZtZ4ykjVxj4cFSGaHAJb9SDd99mdNN0Jujk3UH0NOmm51R1AiChARYotLkMN
xhlNlVMSYkBj7bGPOoQrgegqTSYKdGALs9vq1zvKBoSPIL4n2soN3hu99+MlVY1o
hcIUVWleJ8hf7kObE4uMfvbAOUhE5tER+sVRzYdtXpU67IYm5pdfDYoUKMdXLjve
1F0T6nneIrycGb0/a7ySMPyONNZkIx7bL9a/tNYaReGLOg2ozXjKXVLYiG5fLBZt
SjMnJN0ZWBEw4SyImk6CbizbwwVxxQBUrifbqmw9WhFKICEwbqSdRuiGLt+B+mSZ
+l7ZsXE1euJ0KXLIvJonS7gIsF7iAgblqH+lGas7z6dCoZMemrVt0KyAseWgzLP6
3WmcEN7dr2mtlIDqUDd6UNHbaeyNALsrN1vDurIpLdr92+wGHMo3JEPfM0nhLDGY
n8igbln86lpEDALMWOhQ85YxDjcD7fudlRXtt3pCG9RAgm2AFOJ7BbKzd47AfMI8
BfowOMrr7BiuYjfvkU+EBBhm1xjQt3DleoRyer0TWRSm5G+BIBoHxzSO5q59vheD
vm1O2/381/nhweL/JRhkJR6fvMklD09L/Jy5o54mTFEJfeDcmbh6hXq3VjWnh//F
PRnmLXq78iet6iWMIs37pWnUD8T87lPN4KXI3Q/bFUL3Ob+YmuCFSFlvrEt2eMCa
HuJku0EskLlAArauIiFsprd3jq/emxsMhsBpyiFFSigWgNTSV3GMKbogaV6g1z5x
ERa8MAWCbRsfiXejxe1xMimh3ffIunZsx02n+fatw6TjNOjlbZvIhP1jOpj7I0uz
X0sz/XNeD6xgA8bdnUyh2sX2itY3u7OrpnwYWjcvxsVFT4QQfnX3pl2konQ8Giey
9YPOw2+K+O7OrY1/0dMcx36INNbbV2ozGCnlLLPzKzmBO0X8nkDvWK52OJqomhv4
rwrkYSw/Ckuq7HBI3ZNZODzJoS37w7OoMPZP9ieEQCwFAajJQLD/4tuUqgJSXZjt
MOnzfaNiYO3DmqXocGz6SVs2XBEbTVBP84B0Q7JMZyspKPaUZDXBxUDkJA2yIPGL
Xwinh4+Lr+TH6jyb0ECGBsBbNlet1ws7wmmUTZ24oAXxehMAhRzjBA2ExrxgmGWi
2spI43UaG2wDC4OOMLYh4QAM+89VVpr+iwESzGaXewdUsD5sx+YxkuWfWhRbuweV
nkP8w4aq+hPlIj+Y80PHo8A01s0Z5l2kT3xSclxtvEW14MsPCY5n1UXuteTVAMlA
LeYoEdo75ffgp2/0aES//1Pauc3QRtCJzDOas85ox7QzY1HLvTAsQbAYEG0MVepo
SGSyhEwSunozf6LWtpAF2aodvS6IYB+c/kCcdaageney6WWNhL3zkskNP/Ag+bKU
XedEwD4hlsVngwF5THN+05jcKlCu8mf0FOIcp9cucZIxGMxiYOM9kxTeatUBajhU
tbkIReM60Xs/phlAl1sQePPrzk/Ninkt0d+coUsIwO4J12Tda6Sk5huCj+awOBno
eymsDynth8JMVpXDdkaQdzB94wyjtLizh+po4xZ9pnMZrPyRmv7MOMiE1DCa/Kny
9l7hKUwpRvje4bonT3r09Lcx+nb4zABlKUKXodH0SqxB6cd0AGrnCVuA05TMLeDu
q14wMkJuISdCWGAxMdnhQ17tHM1ZM/KXE/xw6QV/J+WJ+c77DM/6gNkaXJdxBjhw
4HCGtbTp96q6pX9bkHlaQigklfQYotRUaWj/8FZ1M/uxz6at/SdgUUEnnTvJ53S3
SmS9QuEdZsmnvwv7Bz7RYj8iGiA8SwZcwgyOPRaQp2ofCNEGvg+2kBc2b1xBWyxi
5uGUvfm0eHvLneCBj85+HcNxPVpLTBSbK5P5Q2gi45nuPw1JWuSOL7v9N+B1rtDC
BcSz67+sEicWcdE6oBk6cfN+jS846j4AwSejLGRAOdGNgHMnXpHFOHeC+4z1NBlB
EPa3QtsNqt+8Ldpiv/S9Ebm8FOoUPSReRwAyA5aoyEMhpg5bBFzeM5A6m2sy9bbE
eO1tYhTt6ooImrKoykUmtyiYuOADU4HDlK+pSanDEy9Hq65TfKZxVVT9OfCnXw8S
7upZ9/b+/iYBg8obPy/P1Q7xOL5+OrSYErwh/oWiv3c6SNyZKB/G+noyXN96L9UM
qSxki9eqYBgdTv2Pb4cWqFyZ6rDP2aoPImApZR/DVq5x5hENmssMt168KkmelEmG
PpY+VitWCZCgwL5OdtmLLWFcuX4OYi5/CPdoifIdJp7OhmpdrlqejVMi1XEz1KZV
KNWzfjmODd4mKdKRmPr7/3dHKwu9HpYvOz9sX0be+u0NyMJRPB7ZK0kd408Lunok
P0u69RrcPSDJN7NzfBldnbdqsPPT7KjGI+OlLKBtrJ8lbLapJcP+bitiSBPrc0Ub
48ybtrf84k2OKxbwVGYZiZelx2NWG3FhPEi6rvV77QOTocD0Ip1R0HYcW+NLXwUt
z3V6dYSFsZ6AXdxkoElltox3Y/Zj39rwBNwxvkDAghhCUk7zL3vTYZ+nHBVodVE6
c1Qz0cZJGh9OENLESISKzqeYa6ijTQbx6HZohgBCaBl5vbEZmJmBFQXlP3v1a06J
uUIoKiV33oG+AQgwxmU7Im8qkD/xd4XKV/u/IhBSrfy7dDkKObx6vJR+57+lxXkU
yvgs27ixlTCz55p+xxZf55elQqWKMRMHQ2AtNg4SKFaAoXlgqfHup6ThV30yTW2+
ETUm1Axi1f9jYIz9xJqA5oAVHkQh4Aj6l6Q/p7pIKVsB0IYQ+WGEnQKH78uehLVn
KEs/MDafKjSFZSx0RL3jWVCpZ/fmrxdHx7stjHTbRD7A1wZ6tKbd925pNCWDpYJ6
DSOwsm2tGg01si6s89bTJ9DtvX/0xOXAMOk8FJcvJR7GJWXujVWuOOv5MyfYkqeX
VqwtDWJuVz4Zjd9bdBkM7HzKjwPfTs4XBpSYG/2/NlCOfFo4zOBOnPdy/fhl9o5K
Vl1yr8tETvHwYMaBMRoW9/6VhT+BFHVC82erSsE0gzo/b9rq1f4+n2+N6MqVXCKH
BC7EdojJRT2AVL56k4whRWQG01vU9a3Nb6Fw/k0EGZ1nVrKD8dM2g2pe3PiBBmQj
xP4/9kEDneEjDt9JuzDQOu5M8RqlsZY64PFNtR9R0Dqa8aHWHr+EwO3KX2J1GUZa
sWSRZHjYgQc8BEs6Do8oiNF/PZvsgBtF7JlH4xYdwCZWlV7+LCrExoWHKQjHY4PV
cAknP3SetEMilGnKyauEi2eApWlFrtXgKPYNDHFcm8kL6xl+0gehrGgj55YhiFd2
RsZBBwskrG6PJwizUQ4cTdqoO3lLEOnmg6Q2FxMj3YQyVpUG5iTK8YDgdUcMe6tq
DgXFXCeKee7XsYzOTu8hZZLf6tqQloNwIqKg2WVDxQCfAWujAIpPilJVgAKk9XWB
7R78c71chi/t74A6W4R5i06/3VzqNTXSE0MOyLs5E6WNBTt4s9UvD5cQqU2uzFXo
Pcna6ABXxaV+WlX2vmvHM2EVymuggW38N90x7eMJWyuy/8e7OoNeQUv7R8nJvBNf
uN4/esCmHOWPEIs85oHL3S/rxlX/SHQ1TkWCZL+QqSS4aAf96dK15PscjTSEIRb9
DKKqdInmaSYp0pzx9RGv4YR4osFfe2UlmxOAeWJmzDPRQPVQ2WQzS+In+H0Xd5Iw
I/eZJDaVbFp60bCl15886rjDAZGg4TxL8lRBg3IWBnC0GgOFdfOPVjx2h+MBeKvs
dmeNuhdd5iWGXmgCOTAgKjlC3BUGbXy0HUOyaF5d+VcVxLwSF7Yf40wfTtsaq4Mv
0+/r8P5nLYwOIb+VD+x9THVsD9NdmYd7+9yG6PflMxRdWciQBIQ0vcit28WQsruJ
lumODT0caQS5gULGLgLyTup7AF8lDMuIXhxNK6v1zWRRxjRaOu/FqoY9tngektXT
MbKOjTVpWc82YuwCJ+kDbzF60qsAswvRbGdeNIlp621HYBPmDTqBnyYg8jdL+yRR
dAZzT7XJfbrx38AeWXi7i7/OVzZswMixiJKhoN6x5YDSbRalyXpK9MN/0m4XTwfH
d7v1ZWCh9whd0m1ZN4L2yDAwoKIM0FsmzYTJGEz8GUe3N1e4D8g1gv8LkT4H8E3o
RLrSv6uRZCHlD5+ZaNITw93dhIlN1+ZtocWJCGX9HY/sd8NE82wL6Br6zYMFa5Qs
SUrzTsVKO+fVCflkbLrHOC88YLUPvaoJ26b0NTYNjgZ1D3jvxFh9hY6Z+oualy4E
6LiTMA2RTjU3CfgJIeavd4Wjou5fH0lNjl3ag+bW28fOO35M7bH0ONy4F6ANGz7K
Es3DDJYGKB8Ihh4DPYWVaZYWLh4VnA5L5B8RGz5m3TdewMQ9QWWmad5IvCh7JKOO
cfQLmiXKbsJ1iDMdWViB6LnarHl0dlozonW9SdHvVGCaZY5UMACDINSI1tl4Up4q
11NaVxsyXfOH0bvXQCwa/gUXmN9w2tkuR8+rLyjjzQ5gQwA0f5GqV65b0/SE7viH
vbaZOnq+Dy51WCJzvWgno5chUsZDst2pw6ICT+g+25f9ptsq6O3bBviTAUh9Fy+j
cmoUl4tdgooVM/X6oJYnMi3O4IVz8ldldo/bZgV+ap82SQoq174ot0unJ8fjCpmV
WZPOcmppuS7Gf0jx7m+/TeAIO483CwVeJvMSdt8XBu+jZG6a0L6NeKDQNm6jdI0d
tCCXZ3kszsG6zUhURoMOzxFG4efmKpTjnbKqKFeDCuFG1a4l81vqaTHoCNBSolNp
6fGdbUB9xa+CGa1F56cnFPPM2eIA4mgOpWEJjMitdQlP4Zkv3r6n9qvPX3gWYg5v
mmpE4t9MMosG4rjhd1YTaRzywGzDi18Uj1CZJrjfqe68IqHbAtuAcjM65AZuWQpd
W6CqgnCYFie+WLfI9ziifyzm0TcwoouwcgwyEJ/Ul3cAUMBuaPGV5Jl3iInwgFSN
UIiBsTYGXcP6W3u164t5ualD+RDfzJtC1ff2TMpjuyfVanD3CSlPFTpGCr9cQZ5y
PCfRcYa1QtBil3XU2UwhHeYzDkecNHFTcO/kYuzrhvDbcXowLRKC3Xq0WAQndHq1
qEm64ei8coL4ZaFJmWaj/u7XSMT2aa/rJPrI4SLJ5U0P9wnqWRVWJOOhcvUq0gEs
nmibr6LtFIVdy8ENcJEJttCxINY1ZNYmzGv3Sg67DsEeO8LQM0wd/G+zEnaRblHK
NAqoqAzTm0J/Ukm317d8gNAODm6IlwYIKZJCGfi7pW/SR7x2NKtxjdevWSVNDdAU
ygoD9aZfWDHRCAs0q3TTkARRQgToX0EGbPlAvbHc5Oxl+1ghoKRWg0R1zFL8undK
o3nQnY7YSZmOV43UVsxWRlm9JgqPzgts+ElYu/xJB4YQJujg+0Xr0vsZVIVd60nR
wSLdlJ8FBw/cUTOfSlJ3P6B+ZQVI7yt06DcjITsxW9S8tjkM1sREUaqZEzpO5QBA
MhuNh3UUXpvnFcsEPvkQHRvNGmX3Gb7WhD9HuHyv3grJ8k7Aerz5PILWA4sJfF2g
3a/bitFm9hdssXMupumiis7rtxN/Rqc6iNrD6foobueHJFoS8DVLF/gxqG0aJEAy
GTS5R2pQki6KKQmOVCDWW/2fKatsL4SYFX3VggQLRObdICAlTaaaa9royyw1NFaA
ha6h1+GPm5exKVHrZDCKCRYoO8IwId4I2aMDXUpEpa5ywgnvPOfLUqlNQBb/CQBy
DADmiJ1cck649urnk6oHEJk9gZ2MNSPxwmQ2D2zQtB0VKQ8YMt9rUqWv0FXg9otx
DDEfA+k45h4VEZ4xinvYVKprCXjfpgrfPhC1wbYi9xF3XHIpBs42UDPu3kkDi/6K
VY+M6I38u3/ya7SkoFonHSl/xfAY3kl06Sf8X+oMxDY+N7opuPQMXIk4Sj9P6/Om
svwdpllBVtiLSaTCgoRsd7S/eH/HVNTBdCKjhLgoIDfpY1W+A9XfxxZw5yIwY6TH
MKGiCfieRCEdSe84kDcssm2WNgxGwhSdbrvzCUvKuVmAe6BFV8KdNqhHlMhSR9GJ
GKQy3QOXpnNGvg1ycjUjatQBN6ytP7vgoLi3Vw1Kju7dtseLoVZFAHSFKAQeSPEL
duagW3PmSIG3CzBIkwK7Wii/pCcyckpJ7pE1gmZBt22lF0xqaU92b8+at9mxcXEl
plZEjrO3itdbUnpck/KwyQNAXpHovCE1kTeIiydGOFlbAEe60+Oc69hAH9z5dBH1
l8KtAon57+5btyHq1xBGBXBR/rN97PAVHA6Jk+KNjEXVz05gtu3OQEAsInPxlYyU
Wyno/SYPlTAQPOLNWgGY6/mKDfqQk6h0hpqP4L5e9s+/jXSAPtNF7pjRkOfmK6+B
/jgo4jdF8uefCttOu5nlYfsNZhk2ofhP+VyrSH1Uffyo/cTxrPFc+4TqHuYJo6Uh
pQMXov0vgInvdxZPtnqiwBxgfuui8QBOVY+SYWJwMoxyJHWljoZGw34gYmcxvZiL
svkQ5BG92qvxr2his5PB1L/Yot8/8oEGSc4BevpiDaxmfNcx9r3f9kYQpdzbOVwl
cSV68MqZOsy6dgBGnW/AIMmRUGKVX1WJYSU5yTfcUqiV0dod919wO5RCZV0bPxao
fVyTV/E0EbUCMW67wwqAl+JdWiZQn4enooerv75iMQnmC0JwmpBPXAqnxY5rnNZe
RBx7ra5STjrKQNxEHxtzcnyPD43ZHrL7DJmppWDzeb7Hn3AXlcpCyDRIKYFnpUkl
uFeRjZqfhIoAojtK2RpT5vq/SOjH3JT/O33ePJ3tfHkksel+yJpNyQ3aww6hcKmb
HHbOIcSbi6nM2+2qSq++lpkBNU0v/9uvix/wPuf+K3Je45aEi9EEC/dBfGNGC9a4
hlnj0h0eNvW178hA37v+H7FNVEZhzBjqp/NaxhuLuP8pvXchdQCY/TgYKexShRe5
O6ogy3e76RQtBhg5jZs/a0jQ4TX6QquuFCVoq4F/pmYA4VL/YzrN5yauNv56fw/V
lNBHXvPGLcPOUmiqFFg9iS+vZ/p59+kjGGjkbHICvafTs139m8bNGh0eecZ6PLxT
iq3fLkVRRP3c48mrN/d4CmQefApr5SIshmBys+0RBWbhk3L1GxoMC8SGFR0GfbLa
DM4bKraVOhApYJfMM1eLe0H8Gq513hGdIOb0pdiFxIy2FMzaMYkszKXl8Dx1HX4M
9N+01I6YSThKcQdooK8Ik1FqvuLKyFz6I98u1Fwi7KdgXGh530Jt1WN+bwTjX3h6
GWDoYrIa0Kx2fsqMsXhcsEbNDYlrVWwL6CL7u2O+o9u1DKrATdQ44i4r7ucmeAiH
eazATzYq8Vh0n31fJp2eMsLR7pD+E3ywuQAcc+QNoL6bdVWCsXd9Meq2Qxk1pXrr
pzHvnp+ow3+g8RrCLYBWzK2U/ZQNB2miNJdgx9s88D/KBKSiXxOW5sn5b6W5c25f
diA0mPBJJUEvByKnWLIxe3v26fRcOowqyABQPJzpu1sH5k0VPaTvJOeh17zgdNVW
R5M7VZb9tq4gcERpUwW4/ccZKCWRPlJ28A+TL/KaQjDuGnTycI539n/yHqOy5BsZ
aTkxtuDSM6kTQX9+FS7vicH3+MvWy68F/kN9aP2/Ou4SpUoJnG54BSLhPXv8+l+2
n5TUs/0vxv1oPkf78+1OYw/QK/XZy6oPSBfy5UfQ/844czJj63Jq4XD2hLLwOuru
jmWsQ+JwA4iE5zwQj2zMhZOxsPTaYJKtOLiTOjrFbih8LaR8lQW57W27u+gp+UDR
/DoliWg2QxYXSxivaQqy2FrdeYHq4KRyLKYvxf5h74ZBKPd041Sf/dt31IUpGQhB
b1xx2XcgKUST9YXfIc5qdm97zjmyKKLITFFcxB6rwqdtZqWwnKWC43r4BznweFUX
48+rcWnVw15ace8tFoeALRmYMEg16XbBSAKGzwp7IjmZyksKp8Ha8cNmERJkHjU0
FzoblsF6aqWo4iV7WzsEv+nf3sFHFMOfUkRdM1101UwpXshXO6mG6ARQQ/jBJ89+
iQGM7rZf51Nkou8/eGf1GCtkqIhWtOe3NXTdPMuBP62Qll8duio2oPVix4TRu2b3
0K/sqi4cUA3QIZiK2s3DyKZ9SYvBdcUCxS3X5pvwxyfsxsXVZM3jX9u935HxuXRP
zfHTKjOC9ReEfH5OcyqFzbgmfTMThmwQi25Lax0RpmIMogvtHjoq5NDr8FSQe5wC
ieaavp1E5fsp5dZ9Lgh8AJ/tePu3xDe0bcssbM8Hx7n61sZbbtdjhnnmn4lG3Xw2
2vn/Fzpo/+8ITeEqYLrgnFz93VW3z782ITqEJZEV9hpueKl0Kt6QJrGJgJzG2sIq
Jz99ThboTd09z+HkFTYl304MD//O1TLDLemBZZZIruSn9oXTVc+fteMQHp0yN64K
+iWGDh5D1pCNolg+DTpl3MJwY/jhLBpJR6QuteC89KJ5cPAiPp+qhZYFfIEGXfcH
XsDXI/UNVEILuFU4EXGJ4u1JDX2AUuB9hM9jtrMIosdhiIiG/y2wDpU7HOm+Lbpo
dcSA1lM24iTXze2NH6CmSvh0elBLr5TFEjXzB2fvKjM/eyRsF1S9CPt+i3mB4zR2
eD3d7mtPongmFP1TgdYpdJkduNSPLJIaJResmcOCL0lvVr2nMMVh6c4CbxhoYWcV
ke8+EyKlomJPzdvyDD2bs/2lGDW52RORYxIMKaedJ+EgfG+xTAyUj4zv8X9QXu3t
TTHN46Y3nNcLn/NsZtkMfcLdfR1ZTv8a2fO4G9piEsdXuIUaSMnjEc9sUAjXsNzU
KBBtxAtfCNozsVG9RxIdkGhT/X/MNUxfkr3TcpzYb7y3YAhNxGeGFZ1+LzKxl3lb
xvLpZwbkz0ltDUZ0c2GaJ3rNPmmxFe6vAhkfpw7EPXmVb2gQCaGG3dmtHTKmIMFB
SeBLqmMdyfRpKlQj3tB/iUweK7kLO5+T2+KV+NsdtiLr+iuxSSwFo9eJ+/eeM13o
9zczP2nUv78aRnDyhj+L4b1dKIqWP5M1Bv/PQygM2iakLLSbBF+Q9ei3+1KonST/
04rfCiD/RU/Fw6ynuyxZ5EXc0jhfrKl1pF18RcbI+aUbPlMl+UV1+FGLafEOgZtZ
nBchpP096YDpE0swU5RLTMPu/dz5GA55vFtxXoOlsEPkmkzEvaC+6mhhfjdeX1NY
6hox/GAYj72E8ZNMeiR4RV7yH9SNydp1IcRcrEQdiZK5qEK1oezyk1GlMeMxhDWj
TfWQZSduhk+BJ6dJ7u81tE326r8C80h2W+f3+qTCN9IDv3huP5BTGLqWar+KMmsh
4futHzdZ8ms5pnWcXnBTYxchDenrNS4jcDeHHcniFI7N6g+LCQiSfdYhbHmPb2KS
RSu/IehbaRyUbuAbbNkkwdUcn1Ns2Xaok+ydqD76XoTOq75FC7HBIwo/ubRJQsBM
ngykBKES8b28JC0ZEgPOtlHUYkTSAweQsZgLs0pbRkJ7T2zcZFwX/kOsaak/X9IV
xod0fejJJ/3kNoD6yrJY+8sfbjp2x/e1V2ub5ClAPK9Tz/CEH6bYB5rXVqs2D2Tx
vnj0gmvdJ/oNKu9wpVBc1OBARaxJgeVpooifIVxSVpsJIhHjh2JlM6d8SM0QlSK5
v61Csk2471C2c4yus1wm4e2tysUb8yhVhRiFYT0uIBCYmyUtFcs8gibx2951z/z5
YqrDbZl4ywaq7kRBoz7J5bVHTSqGNol1J8jDwkrexJEMgYEzq1ZBptqpnUChI8ys
sjXvVd77nS1QzCNmD4a1B7KGd+Pj2XNvVUHMcA2+qz25AsQ36bQFDLGFnM6aKzBJ
xBM9p9cdWaY/UuWNuOvoquI1yciIQGsciprVwWF90hqQkCWGPB6+8fbFrcE36JJp
EST/M3c5nqxLgcklC6rx/xFCXoOqURwO1BqebPtuJVTzmRIEzQcuF40KK+uLZl2u
v3NSHdQMIc68mluXmfjTYL67vLtsaJz9X6XcNA8hU1jXjb8CeGpApZfcPEGTvLVD
1g8FPE2La7YI21IRStIrO0OZlJHNQt7oA+Ezi7tWC9Ga3YJRTlR1NB06oBYDZRrU
g6r4CIGRp5VBui3SJR2Le2+CmL33tk9loI/d4zNwa39lrKdG4t5KMXwhi2VmxrVv
mc4mrTeXhYCSKoxtNOapbzcQNQQn4BAZ74NZqLEyi3xhwq5SbJfC3aRswea1VfhJ
+w5ej6juxCsotr/+1gpG5HHBFzIicE+6Cw81rc+0QO9H9RhIwHj4ZHEMEJ3RrY4l
kDzHkg5f3FZ7RqiConAbBv6BQBV9UjrjsB9fbY+FSjkV/4MFSctmUJY+BkpYvlM0
IcZAbsStW9O09q59pvOsAIqB2Wwn4U8WsJghn/oJ3xqDOUrrvvODpbJ2QlZ82b6A
89LyPMNyBLRno0xUz4c866ms3UmmhKbqtGMtDB9j5UcT7mXzDN4Gj7R/RiwzSD7x
Br1ofJ7Cc2Z3U602SSHQtAAVe/onbTPp1/bzMm7u3O2QbdapY0UdZHpg5UO8Y7MH
lcM10nAeuIHlIiB5H+KZJaVfRwvy+kAwNF9zqB4fow3KRULTbbzt9iL899+43O4+
ACeu1dJf7hRleC1Gr3ySqVkThmCzW8wRfemeJ6Eg5iRdP5Y5p4gGRudP6xoHHSUs
G4FF1P9ar16ZtjDyFR7z/AW2tDzvMiVBHIBvSR2UnPPVOrVAnEVnmPM5wM5lsvc2
BIRevsW6c2i5/SFmoetguyQsWe7Yq3Wd2FIhWS8crCKlhq31K0Ri/oyjAD2cCkNN
dQGsXWurCe9sW2dEwD40cAZW1l3yr6IHqO9g3iMA+G3IFbG3k+RTOUembYhhbbya
RxVeSytIrqK8jytnG7PB5NYbfYzSnfWTcWEe2iD4v9gugP6Tl++2I+LG1d3d079e
kpfqjvn8K22ttFI0pMA+2wl6BmelURc85dB52MClpI6hXsswz/byzKsUQFYUnxGE
iZKbxnx0S+TanEkGdJWzvoPEooHDbbXtWu9lFxPQTCZGJbabNlG3liZiCzsZnshH
/QIne/viiUrxK80FcEBDuzfKoJYxOyJnTMtnKtrW6yHL/MlMxr/TRsi756qht2Rg
Kv0KGpMSSF5tCfeTxUMt8Brq8Z8TsuTsiiitP7Mh3pJZwv+0Fjv34zrKYiT1EJvm
o0r/8WjRt3wjkhdgnVlRC0i8WV+u+5BjwHpqM0boR1PXa/e5wBG9IoICQQ7B2IEM
T7JA6KvDED8cpJR9xbF0QJYqdudmalPIFwwS/U3t83y3WQcEqbEaY+smoqyKknVs
IX/tb6N1IHTVLC6kF6d+eCvyTV0EYpb/RZziGxLdUIAzDL0NOgEJPJIaiipNFD6L
RTA5tA9mxcGfWnFupZhQQwoRXvgYe+y2dNbOzZp+VbwVXQf+IcQcHiEcuEanoYaA
eL0FpUSVxgZ0zySMSuD/qY7utRwZ1CqlrVt6x8VHofq6DGwWvl+jB3nKHagL1RPJ
DmY9+s35laidXt/8x4fjNUZU3dpHQSofNbb3iUU8GTlQCWFvk7Uf8pmigS8Yew5E
yS2hAg2R/FazpeZCUxNGFnL8nRg49H309d7Li8sKfE4gOZqdCdnkQLK1y8TuQPp5
F1hItL9KqOeXkiEp9JKNnH+xjSm8LhVlvzB+92DdvambXeAjDLJuVwByfPVNZUzl
rW33VFs8y3bRn+K4j/3zwADL5dxdf1o97qofb8aTBiwm5Gq+Zf7iQtmtdbvtNQHR
O1bEEtG2S41vVOSsh6mep1jHLliD7RhHJpu4fIRHm5s7JlVYAoTauim9ufj6p1xS
z9HnRoyBN9CUP4BnPg/IAFpOFwcTjMFGkb4evzSR6hcPmSPQrhBfvijglHgpW6In
c7+sUCEECTxzq5uq+B10sAQ8ILVe8GwkcFn8s1zNYSHkP3+Z6Osah0T/dkfjqLIR
EbwWXe2UZHSdkUCMIWpxkcfBOwfXKnc9IQmYZJVfGT8043zvSZmkJuWmbhKyGLFd
hJFEXReWduittxx/zUknEVrpRRe1EjwreABcKR0qWOS53Ub17Oq7hQkrWjs4D9tZ
AI5rGEIeQ1qmSQa7hjuQOXT4Dy8uwhJxOSIxMr+WdaUj1hPsemKVZjmOS7i+idVF
MP1xWkGz4EWOrM3OFOlcvWfNiabshyGEMnBATy1QaftnOQUWOmdwk2fC3cKiLKIs
pHgrFdT5+rl2ftPgrxYOcJmEA6nkd5LSmM1fl6jCdoSz+KhBCGufTtGTIJVwdv7V
dgXf/etIKOpTfowswWG3XV7vuJAu7nn+WH4aqYiMhJnvpLmRpqqIIsxRENXsIJ4t
A2lVK+4KMahyvSlNgwYNz5IB1EXJTmOVCLP2zCIT9EcCKbjvXOBjYoOUjHTz+Gdj
/6cludG0dWUtKivAKlK2YMQDDK9SmIcsSoWtd5Rw6v+SjL5ZOJhedSWNU6XCUsxz
FgSUSFiF73zomzQ7dq1ea6OwTVcJbxln+Pzom6E27DJJsW0E/ki+Iy2r5zw5Z/QH
aX6YB1hH3hiGjzVocXfay2WQPpoGnqkjjNoN7Ivk7Go0kTURGOKE6kzlO0/ZAymN
+GWxE9NBjxqXx3sOdYzdXUTMQ9jjxMOxnYaHBGDExZDpfVyfHzvnjBGgGHXjterH
U6/TB25+Av/EzOLUSZ8F/tyZ4LYBaiHxjiKGfSn956AwMOyyRj9k+QHXOxMUKGZ1
1jAHgmQjADkDaXMa/MjoRSmlNwaMvf+9vzIb9GtUz3iPRHoZpxHlPe0Bh8bO6kb0
VfLjp7nbyDudN17c93ATA6jvQYXPaiNZKdEUqQPq6hiSHZW9JIjymvx7HtmRe0ZL
kO1XB4ZB7RIh/7FehDQdijchpdZ0jj5TzbRrBOE6IeGlMgUWNJlzLEaZcFkRY2GX
Viuylf8f4b2iikev/c+AIvqLaz5sceN7KAFqrD3ZZ+rhgZqsj16PS/5xXU2d1v2A
wVpN/Z2P66PfvQOaLkqRiG9V3GQ4bw1t98XTbcYgrpqguMDivKhvHU26f6KUco9M
JNS/qo79RlQzpQptT2F7yeU+FSn0BU8u4Bca+c7TymC1NC27sxqg4S3ktLPW4QSZ
E2zsjss5UV43hiq9IDEGxs1NkanF/lxBzm/B0G3I6YS2PfDCuNZg9Gr+svue3R1d
lJtTdRe7jOR+2Am8r84x+QrUcZE9iJyFcINORaKThN2zi/fXjcdQxOOHbd3Xbuyu
UYrRNYuV/GzGX0QQORI/84s5ug7ibBj/85Xm9clvMalazrr0HW4vvjdcj1HGizwY
6Tvx3yAJp/oa0wwu8IoekE+ItcxPhRd5kEEiJgftyJ5lt6fF1AQECl0yIjIAFs/g
CmkGf+lSD6EA96+PKOhBUY/D7j5lENkEP/P1OvBipqlLymf7ZYJeHN5HFRC3Zj//
jBtv1N/RciGOh+CvwG8F65FAkDCHQCLuGbosk3W6Uz4m4t1pTrfBSxIN4ULCypA3
C4tNld4zstd9ES1/cMqRjeyFbCnCyFQNiYE3BYa94caebL6TCI+pYmuSqKGsq2R/
UjQ+CLbgJS0c/9vDBToUd+XSDgSHg+Lq8n22E6QCxYMz6AKSMD9HoB0G9wDPYPjl
3xkLxoVAdIdAROBW1n64oRsQ8YDFfsfM12qjasEXdo2bfPk6ht0TwpmDEm6GLlaI
gmf7BmLPDMH+7qr9/eKru8iQytgLC5Rxa7H4EoC1KV90MSExO6LaUEXnoXZVogwA
7q7kRvt+kmt8FudqUgHPHRQVnXqJPOmee63GYfzoj/KIaEohWTrtiiUwR6g/1N2I
VLmDFJ1hZbFXjb4cKcqgVrYYJgKVGBfhYRaa+PHCcj8Co1y8dfF19KHMDPPpZEU3
1KFuv5zsh1GYCG4X35uPYjlqQxTsYIHGxfg8p/cc2a0Ghz2Gg0jlVkpbfI+zxZvT
Nfl9yUvfUjS6HHkucQottvlkJxteRnnd6HEoYlJxSMYu4SfrQY5s+Ish0lUV+iec
XgJDl293HGVJJrPuUhu4e6ib6m8O6bYF+6f/8goLrDVqHsfz5Zw7Qei17uEhY09b
CnxpYvqx0tYilNeJ04/2PGjUji8QQzgnAimiNqTCITM7faqYF9PpIuQwmwrX8jq1
GQVgoL366wWA/QO4yqtpPrHFgzNAb0iLR0iYeN3rkZhMdJgoIgiBkVzCYfjzS49w
9KhI8YhVF9+ZM6L58+zuF1U0GvFjToZFGl+7L6UBI0vFTtBRB0KVOy76MnfatROs
Fq7ssxRV05iz5ukx2DqIo0B11JLjOpVGA3xh52bNxywCPqFBs/R9um/xyh9JTAXR
GgEQ0AePLFFmNNUxU/MwBpmOMcS1bpXmoShavLF7CyFYRcPo+ge6h4PpeBYJ1DaS
f+CPH/aXsl6HHwjBggdLelGg7Y/KT62+XLLFzgWFW89i7ANnVBbqMN/SneMBSF28
ciFs2yguAgoUu0l8NYZNEpA59WqICwIPcxfRrzw7p9EBQW4sRNJZ5YTIPNhEIST8
TUSY/pgj5zpluU7KX2u+ypFekaBzIWJsQjCxi3O+ruIe8/nCHzTq4UWKsxut+0du
zE1681JQ8FysfhAGxyXpRQ4p8T10c2Oaug3duVkOI+2cFjJEKXRsdV998NfiAn9U
iGHpdyL/j40EurBB6RcpQVCkgV6fiZaPBlDPPi6qDWiB3mm7ngdKGeULqWr2abBp
yhfKjCq6bpeF82re8j6b/mfoxvSB40+g1uTTHpSOf/eqckWVKekGDbLXiuuw7tF6
XwBV6SXKfohH9drd1BApCI9S66EHF9F8JaMz9r8zZj+4067U2+GQvPfnxueeIgjq
vpkFUBh79Yu9BpbIrBNtTnj1fPy+lmxMpSzyuC1vRXYQk7UpBgV523Caacha8qIH
bk4RDo9SKl8t2OgM5ApY++cIFwB9Tl1yRa01oA/ZoR6Slcg67xWl6cljVQGyIzL1
XRj/wU3ArBk+Y9vUBuFfC/AY+33KmpkSXCKjtBwyv3NCeX7ZGMMdLxZeKT05AEHH
t5tHmu9lFT5nF5q3KCebr6q7+DQWGHJA5nPCa6BalStYf0hbGq/AwXQUusi3SGaG
DG7Hdu4TLjenJzhjpz5nEYU/+0i90bd9kP1qY8yTiPkoCRE6Z5Wh0HjAgf6gGoEN
k5CHeRtdNRae2HCpQjBhrXjaWX1iEA70T3j048T/180iJcpdc/KAkDmnamvC9iLh
DxZHFGwqG2Rhi/093GLsvBOm1wxeEeR08r3QSzM8KTtLNJ9C4Yf2gMm7roi4z/MW
a/2wLgBO/Rd18VVbureA6opiqjShj0iQIjm12LQCRJvSx+rw3Jes2UCoaHcX6HXZ
uV6XqWK8NOBfT39P4dkoUnyNzFxvLP6r6xHOQQ3ahmLvb+qE9j2N2jfMcTZ5Az8K
tzECK41se5FYQj0/D9u8Y79pyjo3/G48Bpt9KV8z3sGdSL8fXpWuCl+HfdD+ubwW
v5Rv62ESIEEGA5Xa5e4MGGJTHAeKgPC/VL3ULWcrGEtTrawFOJeMsXP0VRXIpKnA
opMmtrZqJ8Uc8/eYZtEnjk6jLvrPGTywrJPMuUtHBuzu5+gBGqteDstDI9Ji1t4h
I87TvBUr456i4O5y8wyTTfO7mKQbKPDe8bLeVaJeAJ8XE1USyEn+V/E7//nY3MKF
h1rIzjlXcInjVFudA24GMRJh8GFcvIJRBxeeos/0K34e/FZEIA30Rz7wX9HCY+4P
aIPQQS8a6SkLROeQORHJDL3Gintl0NrJXdeVtnbXnRKQoaT0NXlMKFWq3u5MZtAp
YF2587pVHSMII6gk241XBCU4WDZpmcerYYz4ZMuv+Xr0ePvHYp5KNlKjvtwQ9XKz
qlY+Y7lBaUleCDAnkqH9JyhgjrX6bdg/qZQkyuv7IsubhQtRFv4GNYUenu8NcNmR
AdHCIGDoBY0IaclamcUJEMDPPfsMFTeWhdB9lq3W8phHLVjBgNNbk2ZOYbUdyPYA
fYkUQIO5BK4/7UpDCTbceX/vXdaP06ibfnKiAWUkiTko+ewul5NeFvDnFzoAt/1D
NHv09Mvyl6J9POcnzy7Of2BmsaQja6IeiKaRYF3wRxgX+9GfvgzVb8vyb/LUFERu
7jLeA8JyfX3mEx8wfWCcWy3VYV5geuvJzpGA5YDvNg5RMD+Skgn8JTMlx3DzTsyo
J2qrTkB1vbr69CPH7uZRZffXO/PTD57AlI8RJeEG50Q5G3vKywWPhom7GAns0p6R
Zjv7UCYP6dRlBcQCPzxQvatP1jQpMNwLNJSaecbk1TIRxcGjqmwxQP7g0C8ssAaw
eEpBcMtcrl78rwxSgU92UlJWAAed9FCQZWGB3uM57DqTzs58oCZ/mDTueOYgvKDG
2IWcLllARz79ROIrhd2449T2fgUTNvqP8m+ApanxVh3l08h/LJhq8hGwIJxMImcw
GCOt+XYDAFRxDmpPxmrTdmpOwfxfqnrUYN8kpbuK/icIUjogGV16n+PpIiRLeFn5
k7BqLheSNxOY5f12rf+MrGtVJVBO0sfcyGLGs8gSjv2AKRARqz8j+TOw2RoQfjdz
vwlDeGnpRPrppyzQzIJ24ecI8GUHW0RMaB4lzVRepg/JCvAZSh/MDLG0ARSba8PM
jvC44xetHn9eLE4fyromEKaCYopeuq3rL1dB/biMAvSnS+viNMTrB1BTPRjm53Dq
LDW5Bi8VzHV4H6uBSUM4WbBxdsvhZ0n0UN3zovup1Z7O+8rejPCurMgpoQFzR7Ah
UQGBIAEzeXqTXbQBPsBk3T499sGIrsEvhTGW/jjuz5BxDqU3rpzheEnlPnP4/etq
TDoczUk3/JruOt/h+npp7+Eorfk7GO2WUwRd8WWqq7lVBeIBtRYkDygqNPj/tZF6
0DA4AAIcDSCNtrcDCu7OqthLKZy0m4WwA9+eqS4vCXsaF/6bIcY58Tsr5Sp8s/nC
6HWPL9XfRQE1tYJh3BoYIice8PIf8VYWnV3cI5XmiLLOR9sLHlW0ki8BExlIFOZK
IOjaPrR/NE31GbpmX2W9V5o3tACNz+tbgp38zsUMdvNDGr3HZRw+H2F+fFawhjqB
J8PSHI8puXXqrkFhrm3RbX9bCngAWQM8qnmc8nAr4q3mi0GRCEUHkWOHU+IqZKoH
AP/h0s7uy75rQXXRzZz7LV5uuzJpMVKznzJb/ku2swFQ2+PqHYuI3b5mbvDiu8i3
LQaYSf9IYkB+YlRuyu9V+YdWCnQjwaeyscZcjqlvpbFnBL0e2e2YyVCuj61ikr67
LCjIeHG7RdPemwY+5GoK0owbfZX4QlGd5cRqBtj0aZiGpAZiqbKq2AmLZjQJQXry
Dka45evSF9Gn5kwSZ9MlyZOplNQ1X4mJ4WbW3w76FmTwbRjO5H+wpiO1va3vxaTG
MBTxWbPnQFiqVxjn6Jg4L/UwlxkkeAV0MthhN4/q0UpLUK7N98WKU6xLFt2tOGUr
sCKUe5SUGihuoets2NTfXbsIpaWVyDv6KM1wXfMXFxlPfj8Da5fdpTVtpzM3znkf
tinpZagEBB0Z9zg9lNd1B+/KV24dnrCfvzeCVkrn7QK98gvDet8vR3CRyDXA8Yqc
q81CifaJ4k86sZvpgGviLVqJUev4T4t5fcfnXI2TCgi770iNXe66papzETQ3zkJU
dhW11lNEqTO+3lTjgf+PJxFbAIsF3pn9vZL40qZCmiGvZ+fwCahBzL9kYFTMobgS
Fb5wPemsloHmiLrSVL8/flFJU9T3qHUVnqeCnrTalzVMO01Gkyjnxdq/SvkLpOCZ
f3LB4/RT5LE1s0dX3CblKxOiMCOkk4dPObxamV+g1uuMloJGjufptzvVVrtSn58v
2EKaE5TPLi8jaEV+GDRUJFU934yb4ALcW30MAOmLKI89gH0LIK0W/GIttLp97ll6
5APa1geVXTOm4FcrMa+wjrcJOGH9VEOCNaNlsepViSfRjZiYPQjniXjXuckGbPE+
2Bh4j5FhdMX4kL6hr+uggurctrFaDbq3Em1+fpJGOEJU+BmfwU2HU2EGfhwc1VuE
jccQsLdCEfW37NjKtYuCgrmhQuz4QdjEYe1KRy8TJunAtoe2dmTszvVOCAkXJjfY
LH3SN9VvQRTWqR03mDa6gK+06qMQZHOLnoQmQ1W7DCO8OGep6GmGFYM34YlbfNiq
rs4Dw39nXtgkamwjCe/NWyvyH8tfIc7KdxCaIP3yZzAue0FK8LdJtyJTx/CJ3EGA
2zb8gANrXpmncQyXS0EeOpfUDzDLoPiOpbJroB3WyhRtliQIJ+pPlpYfPFjnWmfz
SqdYtZJhPjdMe1i8VUBFzjXM9Iypoa1ZEvqqmNURUEEj4o661zPv4iPeu0JANIGA
AjKalhbT+pqF3+gtP6uUpEeavX5ewjdzjuJ/XNu4h5exbx+8f2g5EZugIM+MpSjt
MZUKE1aFQ/zZiMq8OgFKeWCBSnnvrGYnxt4lr1antUacfIY4fT+jVGDYvW2OAu1u
uI9jlToo44MfbCDDe30/HMq+n2Dq2a4FQQGhqw6LW6EiPybIo9/Yi/+sNdWE+2JG
uufWePNdtws3qjPQt8cqXh9OJ3mMR0jyot38hQSbpkjdlaIxqo5ImeWJEpm9re1F
Dhfl+OuB81mVSI5q/TuLrcdw8L1fTIbRa1ZIDydpzUhV/RUNB8nQZJmS7KosaWgC
LtPTDoQ6dndg7B6jAGL+hor0p8VFBKQJhpxu3L4ETNfsDLRNDTwvj+QPAABYwhJ4
3yTpDu0tNmlHmTAh22dg0vs8fOATRqDp/3XSzw+MeC4DpZQdTKZHib6fkwunLl1R
O+x1k56+KT8dVNWs3xq1WzKEFJfGEgHqa6y496/CcvyKSkx4AFWjIFDw2lD+PPDb
FiSLLoyWA2QtgbL2fe0LcjzzWeHc645RDwuvbduH157f5rSmuTAv/pIOxJOkJFPr
ZcTZkhDx4DEQWtFl7ZkB9AvIMPvbYJk5oRWf3CzpzC/hnzB8Y9RNvzNnpf6ki3L3
MZWWecBJ/NYhfZR8qmRjf9k59/vTOyI8S8j0CUAkFDSot2AzJp+g++ucGUpuNqRb
O85tfsxoYSRbnfhyqGdlirh2QTJMonOTp0eJFPPzrJtQSInPaEDYMuuLXSLhCriv
vTLG+Vj1pwWL2pJsrZ16wYj8GV79Gj3/fJadhhs+XaNSjSqwyjk4lweLJz9z2eR1
TPP6pkEPr1YY0nzj/3mjTrPJMInNMdirQKxtt+LgfxtyX5DZJHDWVudhzTMz2PZk
HOL0etSGvDgQavfdA0rosE+/i9jBfBOs/oWhphqYl6LcIkNL7Qoa8DECgVOSrYSZ
zmJgD6hcJmA3yICfmMB69TIH3qq/+pDdkpmYDFu97jGBAwyWANr8IAl1KECJO9Xh
Agtk3yLP/oRTVA/7cWmvqC9X2xauuHZTiOF/Ue7Y7n+FWXkYu383HKLGZBg0OP86
kwDZEwpRJbPON+MN1sD324jZPPkRMkKKEmgaReX3nEPfUF0I7nxNHv/C4D7etzFu
Ilv9f4o3XxnjWTaSBOkQWqPE2dlVFXUR7cio8tbw/A2Gv1EPVVdBjC2J3E0xMwDz
63aEtExBYAlAkQbvrwxH6HgxaWFELkkcJq7pxSNrJgY6suNq2EL718l6jaMn59iX
wWGqPiZKZSUWICmLzrjgQOg7XdD19RfrffSQ4nTfPO9ySrAAIai4hKIeASXVI9g1
3z/QJytCx+79vQEzAnslUldSxhNxafHrpH860PJQcxaUY0zp2/hodx8Ft/khHi6s
o0DM3FVlGggHrOS30v1yE5d+TkvuK8gEKX2ESufeA94te6d22DIim8JGrj++nUx5
8XoP3sjQwAH/WZP/H/jv2RamHaWosvELLaJtYGPc/JJEnQfoo4D1Eg7ekW+9BGIK
/+qKm0Ad0r+FqTNpZjJCStSLenQEzA/9crpStXI1/tt6xEoTES1pmIR4zCsxOT9f
CJ7myEmYVPdCjCfHBg5meUV/pmGJklOmbnBHkTcE11zCb/7Omkb8FbWyrzfk/o2M
pQLMjLBOB6xiNu+LI0Ep0elbOjAn4/yPqmdmOzVB25FzTOzjWGID20FW/UF2zRns
0LPBkrhyWYm28ULb2PN5vg9QQiqd1p74TlOJwUoFo0+ZGCstkUbfrZMvEr91b37J
WkpIullW0CABYzhNlYdf3ii6sdR4UWhgUxOAR9KWEmaMjcvOeT24w8c+DjePlBq0
jTWkhv4sGcfGl4E6JOrJsCmwvyH83qvNlBCkfZlxJvfxWJUa40jF99QenokZO5kX
6J0ZzzRX/Dha1wO7MNtGcIMwhcMhCNFpvfSOa080N+EaOrGeArssTbpyMApEnGRn
2je6reqEygfBCMP/Am0cBZQ2L6eF121y0trlyxtpUb+G+Vj71vJ/ejCugtzNfV2c
SCefncRyrXzI6P/go1mPqkI4BRsHbiP392nPxO1CqHAEzI8kltz01qWPk4bSgkTN
jfWTnUrvKdpGpqIf7HgVIXUg4fYXZ9pSULUHEMHgSmiQHewI5jHLGHy6mvR0H89O
D//cL+XAvodt9kn69n5XlwjxkLJk8JPaSiOXlP1VCwhGuIfyN/mmgqgN66pmRm5y
uM/jAhIDxvV4iyHWhfufbvHjovirm8U68WRCsp3FgyI9LPZKo9/eBwHtuZypTpF9
/MZOIeAL4IKHeVvCyvCviTJhDUmnLtHt6X8rLGpo5Dul4jJPLxnWqOtbeztnR0l6
wfEYlt+siTHZTUzmul4bPPtJ8wZS7NRZLTQtC4FdiZRTYBxkFHtd5htClf9weSrW
3HlDQ71Ahd0/rVZqZgT2lRBdCT860qH6ekiiZGKIRj4va6ZBBoeEAkp/R8j45IY0
IV3mYDnwzE76OykH+ramKuP2ohet2y568H4zt3egYKTJk8oYrkn4tx9dU2cxM8Pf
dmVKqOmVlAdkqV2vUZGb8N25HZxEyeZVeKSZ5zohJXI1c9nmNR9cYYqVtitrHMED
GHfSIuNNunjZl+0Jl28a779JtcZ6zDmToDXJsnsW9ZlMHzRc3P3nYqdIda6MYtxR
OOyj3w4lsLlhcweVPFpKSS+AA9yRWkoT+mJ02qV6EGZSZ/h9dcLgflRagc6cVgm+
mWiwPgmGx87Dnc5WaG3kt6yPqPgMiW1YbKUhXQTTLtMQ9tLzwiuaQ4d5MEWLgKUf
xtsssrx+R5gAXYTasl2lFqnzb/o3nx9l76LIVT6ocC4NIwkj33AHemWrKFrGKYo2
U4X2w1xso0IoLvm4C9SoMVhamGt79yeT7jGnE7BiJek5TfkPNizP784f+ERl6rxN
2pP4wjdAGxXY5b1W2glm2FrMtUpNt00LM8diGEXBvbbKEfb8asJMehVHhLdIZa9i
r5Ag38ZbfYwJ+b7prkOfjN3IXMrvhl+8sNTSdUO0V+NVtJsPCKvxcoS+IMC7tBgX
DvyqC72nd4i9lfkaw+SZTZ5dCrRnQG/I9GdVk1Iq96ieqiWHuFNcQp6dIfgyUfuT
MP3slpLioXbC72Ytx1w5gS+H5y9KNFXI7nOCOjxkQGT8qQ/tKxHa/gJHxgGNYFUs
8V9jPVdFMH2p6+IeataX2nacbX0x2XvoRq8bhce/JN86dnkriS3dZqBIpbM7EwIy
ilWNYPZsfXu/kye4giqTuDkNoDG0y71y6I4etg5wJblDKnlvHpdAVgn4A/vgAtGk
/2/zkJvRjoE4fbQFtN3j9PN/AZUcIxiR66oWCXxancziX3wkQcxT443a4HYxGF8a
u+3vTeWEjrcP4Nu9KqwK988r5Ki90btMUK/oFCd6yrZ7CSCZ2ZkqvDu1O8LdvwLT
6HfeDgxcfwH1BzBxAxH1/FgOWHSSwj3MfkpBmhLU8/BfgkAP2GG1ky4Uh9Ddy2oW
d4sPyKOcYkgGikuplpS3WGvq/lUJirbuZsv7RrffQec0+xgza7JP5oHvzT0XRMlZ
T5R5g6ltZxLr7oDk//WuhaALYfe4915pinazi9tzihIOTM8sSg3SpTFupLwXLuIo
ce6sr0idn/Q9CQi10STBQYFkOSHb3s4tOwm9zOv0H7pwxIjwIz8V2NhYapojBeE4
58TW6D3upwtPbFT3fKTrC6ab/ahv6c/rykTPG9pH2/yEvMp+LU8cj+AzXQU/Ci7m
ecF224FCfwN2vayGgQfhOL8dKNSJ7FGughEqoNvjutMMVtsb4qs5iu5q4915jBBF
sqjZSpyFxTkoYarotRz0qa+d672kfloIpSKyKYfa62LIiaVLOAGXCR97B0PjAEWt
VndlHY6cCsmLghDwHPCkIjc27V0Hjy95Au53FKBAc6YKXMlMrnrsKQ7Ax/ihEvaV
w7DyAZTQ44WXL60TFDSiQNbyTnhZ5oZct2Bu6MQhHAD/Vzyh9uBW7BHsdepw1iDT
fMaKPcFHjwlJWJrUw0SsFDgO5vBuxNKALFnVWia+eSfKpDIFKOE8+kgJ+D6J6boO
qACg0djmTcKYh/wX8cgXFF/SpReh83vCyzOTxov9nGuuuCowYXVhjvA4/vd/Mcnt
BZV5O0L0vE44yD8W4UNefSNyMn37hBogb4In2S8gwnMkgHF+oNWttFZ5emge1pAq
BVqaXGq3xujn4E4z+2bkFNDNczPL1o8bJFNwqnxUPwLZsOASiym+puHrd/Y6iRIj
A3NV5XTgyzaIBZ/vu62epXH2JhLos+npYAvPmFkDFzszKdig6zR3Vs3bGB8gJGUa
VqZEiGGsIL17PJdBkKs/zA0ybdkX+M6jbferZ/Oe0XodUJmtdyZR+Yncg6V2R1TC
NwYw1RclC++IHGy1CUS2UgaQQJ49rCo1LN4AG5qOm0VU7G8FnkLzsVYcQONxm8tz
nLz08+v1XEollJhgQ3HOdIVGrZ5SiaepAw3N6K88VYwzY5x2GeOaKLJsPtUy8e9T
ZRrfPb2OUl+Z3R2derYzT0ip3cFHtHaE5oVe2imLHkJBMzqTpBSX8wVnXQOAiPmf
C0LiBsGM9tJAPj2aWjzSty8fFei7uIhn+F1nE2OvcpARc2/LgFjKHZfLMX/QFVAR
aTYQLxFvlkMxAC8xvvc5+Zxlk/TJ82xAIZUdrHSXLGDIUqW1UxHP49zqEzphtuBA
OUrCUVXcAJWhsVtCVjtfJcpUTDfGh8z1ISeXdbgIiA1O/VpenzPZNECMfzCTZOc2
oIa8IZ+TQzmOUlE5QyW+5SYZRoK0k+d4S3whhaNGoeDiN+QPnQV+VQPliWVAd+Kv
aJV0MdqMsCH019w9Enw35047pDbFkjZ/aMNP+8xcfMRDewhVW5bC0kAXtEIhCO9J
1e9wNxSg2w5BDC3K6bxDIJwOA8/lqWvkcOlAPeSQnyiZy2TNXNOPNlKhqzslUfew
Rvc9DWNeZzgNcEda17Yh6QgrvtR58yI6SFFqp+qAGiMqOiDIgrP1bz+CoBh0iUV5
T1Ar0gK4M54PlpY3AtLE5fwt7BFJxMG0B6HTCLvQ2sBXt/Y+y0Qs1Ce8uvk9FjjP
+juFWC2V0jGqFc1ZmKGL0zsgRx0Rsn0yCcr4tdhQLCH5TN7Z/2S6kcb9TF3sMQJy
PWMiRHkRKBLCDLeBTzY9qEn/OlZVj360yeBv+6HupCOcDib7aQHVbAAmb+lA2QCD
VCGbm18alIMb14cucmMgHdCxJO848HN61fdMFVJ/R6Ilk1WzDjRvJ5ZWTyY20XiB
a2iYk2N1GhGCbZazRfRd43z5YEk6e8lVn19K+YZX7DJ84JsSK4dK6HqtX4PwJJU9
OeymS9XuLzkWi2Vu8Dnd0+futy5eaf2fipGwlsretK7QG+yX9Rl4VBqLA5fh40xg
++MZpCL+CF5Rq9Y+zptoWiuolUure7ZMUhsYHv4Q/ycHavnOqpkfI6NoRoLHpwmW
xeDsLJv4O4yRm62m1ne1BKlHDatXMupk+/wgBEvUKUPZGss7EWFJde0AjKWYS8Iv
rlihDcjHeSBisZoIMnsNG8RwR9nMVVfbOPuLkyyquYfbii6mnIHGZ06hQBlBgHAE
luld3GVCzIsl7DzGW1fHdTxIzD3IorAi17DUC7PK1lNhwVywlA4d2KylB+CXqZo6
8xdd+ARKw/hT0YFNYrCW+2PCwYW862E5E5KjVExmcuOW5otCQAr6AIHTKO4meK7d
iCpKDLV3fNr0qk5R8LvKkMv9zRaBjdxpOGX4hWPmDjW7qmsZCItUilDa2K7sdTeC
3aFvdLFauBeXAW+OJGXzMd56GGDZJFZd6sSP1zf9Vb2g54xO0lbxJQPKisEkY+uv
5o1qHlv9k+uiWDaUBQfijclQkvQsh+8SoTv6J9UKwv84VyV6J+/0eEL9Mk84df2n
p9DJeZpqSz2yuatVcj5ahnep5gNH6oukGfoKiLiJB/8x1VkBc3y5bLM3ZUD4CNjQ
uJ5bZgbbrYgUBU4ihTLkGU0RotzpIyC0ro2ateBV8xf+llpM8UeaRmbp0f21COty
g784FmbaswEGz3l/VKgfWl6GRUjgC8ZNv/4Jg37I7rbM4djagHL/+Rb0uK0ozF5x
Gp5C2nZkZDVXBSu9v/J2CVw03a3YeRuxiELYl5AND592s6vOda5TQf/1RvGscNY7
utNw7bEJ9t7LfAGnoDvCJdNR4I+63B1bQi3TYtwOhEsGmJgnBYPLX1n9Dw7Q52zq
keyvl1bT94Igq2LPsGFRsiJ81rlrIxvI5/QL658ZAMEWzIshkhbvIfV1lWDHr+Vm
8sZ2RpxcvZJwFmjuIt5daLNP6EVXJdgscgVa35QWn8AYl6qCuQbGWQc8uGQ3a+qf
ZTNjbKWqLy8nBha2AUzWfRRI+ftEYQiRBz6WWmfYFag4xCZslXZFCu8wceLI8b1c
2wJs33CKcITf4IdaUANK/68TociUtxGv/EwEfg5BXJ2maqqtsOHzJwNhIA03LZge
l1H1ajFyCsN6f1XOyBknic3AE6c+ApEQ8aHWR6bGnPdLPvsYfhs/QCqsYFKyaKw/
bK1ymUTE6C1PVoGhfyBix+qRZeZoWaBxZSFi0KcH1gfwZcOABnoIdfodCW3qetqK
7blqaHJTYvtLMKOcikJuAjjq6tQw8L5SS9rfV31oM1yAv6p0BbDr0+Qtd6qfpLwa
R2sIjOdK73EqM6o5i+s/M1C25F/wxCWiSRKExTdV47y5ps5DPAd80ILas8+OJSq8
79tipuTuI22xH7m5UwGPvnfMvMtelB5kM5/E5X6uajIeUnLLYDU/XCzV3fdp1M9k
o8XfRghgWBUkfBVhx6kby7dInHbiRwoTBdgw3Zn3RRmNzt2JRza9QxmbYMQiHs9c
BwrMrzNIpVMxJ2fUdAMAUSPcJbvjPoJwXZ+Vz/LUItI3AvtD4F4e4QLaMUpMq08X
tactdYjSxuq+/cHAKZAWbfme3eZx7ixZ6JkjZGcswN7wVIiFfhpwJdKYMHhusgH/
4PfdYE3GR4xIltp3lPpLbr2nRRkx6573zUoSlrYkxbIVTIRdnukLXb5u2qRxDta+
4O7S67liiZFBLggdTAFEYp19/nhJHlCHrhpWeQ8TEDqUEf+3WOVtGmSLoGz8ef/L
hQmImmYxCSG1L4VoRdLvSxZ7nevTpI9CeLMpXNVAEP+5M/F2awiuu3rC3p+Pv7UF
tNJB7Hd3rsvPQLqCX7wOWpor/YTHctygnjb9t26idjwaKuAiyshVzh2Ej+l++24w
0GFtja0ygJIQjGCVReL9cIwExwfNkd/okQIg00PNfZGGhZke553+HuxOdpS3Re87
LacWdZ5M3/gqI3QRLpL4nWY5hFin5mNx5mn43oV2+Z3MlbhEvSWBi27Z7ritJK5M
Mlvd/+uIx64+GP61T+UxVZyWrbohA7DBS5lVOjTeu4xUEOEyoik+ncTrNV1AO30m
wbPFrCGMNHQ8fdrJTIuOLHfeMo8ACoEWwuT0ilBMYeGf/cbB2uon2MF+ckFs4o/r
dxQ3qeCOdhLdYflY2h42G2ssFaRlHTYBrDl+GGNgvBRtai28ySX7P5C3jYw1guZN
O0+wexC2aq8S7Ew7kt+Kyhz1XW9W90FCCN1pnAyX0yP6EaRD9PNxb/P+HNdfXfLI
ZU5c/zal5MAgmwoMbO+pWj9VZtgAqMQpWZR7hUCBe/ARZBuhWqNg0F0V9FnumNvK
S8fZs3eqU2lR+UYqfi/v80w9Is3+WCJMOS6enjnHfO28d32oodoZdalSBL2xGQdU
q2xdcH9vtWDYBVClqrve1H/gD/xcw/0O7DRTz6o8luPIvAaId0xWSQEm3CiDz+Oe
B0FnYLKZnrT4V0cyVPByoispbh91E6LQDvbIy3wdQa7Ei9SSCsA9Hr05lIwxzOOP
26AfNRNCQHdKiPV8TLf3E34W1RAojgp32mEH3LoM0oarhrrlmYIsjYE05A/hJ6fK
EJEauXE5UO/zrCnQItynHQMXEvibHX5QhUvvYmdtBPS+8QdzFwlvEz/Wpk7jCJCR
ao8BfxQjINEZm0zGUR45gfa7b53BsetMXl6F4bhL7ju/YZ2nTRpCgWSt0MmqM+qe
wLRH15+VrsRHqxLgygkeXN80w1a70WrItwjDfDEoBkK+nKQw1hTUAsrWrPM2F27z
vnSyDvE/Fz+rBWTZskqV7R2WaeJN5h9wHG0hVRuLzuz7QQarGI2q82dvOI+B+DpX
2qZcs8NPYGxFF37o9Cfy7phQpjo/lO4+EtaqM8aTIutgzWLIccnaXtICNJ+F8ep5
yF8s5XsntP+oGxEOphCSCGLbm4KKJ5kzK7UVbs35AngQAuQm8oWC7gLcsKJZZTCY
pT4/0MZZzTU1QRC756hnQ4TzPJt91lj3RlugxI+KkmYBxHhAek6d8XcUoJJhMvCH
gde6ZPoGBs8ET/FdFCd97I4TC4ew/LnNDS5ywgLA9WpfjPInO6t0eWT9kxFjtz8f
E0aThPu6S01uXk3rjj1hL4akXWr/M7RFf7vRppcGLbfAj0oBJsFeyKayweEezTOG
5oWPIHJYzeZWkJ7GluMyj8Rzj1XxW2mwvXRyR2Qf0psIOXp6ssYYZ2RxWVT16fMo
BdEuAAa4NfDDENaTxkLB5aud63hXQf0aZyWKBhCqiA+MlRNOs965leF7k22LsWYC
sPMxh0EssrSwl4J5swBgPgDfzjBuj9QfwsaYtn5WxldgrPv0gSx4UtgdmbqzEV/4
iRQHLC3bOJquH0jiDPmuNLVGHkFD94mL4w4Nr1c23xVDfLxMCDhLqzeuCf9JUIgA
wZ8iySWcsOBtZYVg4JCVcFlzLlQLMOK1tZjPASNE1e4TBuGmI9IpNkBFkapLnie2
MqVJPzvcHpVtckXXYuwb1ybx2A1KAv1HiEnLRuvcEcbEuXBqn51eynOaJbb97Jha
E6pDvxCjNg/PS6a+dxhogCjUlLwLcxKRyATFsN0leYlh6FEsU+0SIFp44sOC/YIh
/k1JKk9KJcIFfOSHuXE/KvUX3KI268PHwhupIXMZbGZmiyjGJ+PG08sRh0O1APUS
NjckRGHgoUG58unQn4FvWHxwnpxbmHZzCZYCCtFiqeGfLYlYUGehILZkxBmJYbnb
IcwTLwij5PaPm7MzNmXi5jwe2cf9Tlf319shHhDmFWDAQtMlnTES4rKsRt0z9vsa
eyk3qvIJIlrXL5VzfSd4hWOLrlXix5Ci2n5NGk83Qg3Pr6WXiBbSiL5x4zL+9m+b
8iUfetmkpQm6fuEhUvqGZTKG/OvJYjPbK3mgSiF6mkDhQGjoixjo0yVnh2gY6J4L
5nXgtj9on/95wCTbw8FyNChDwb1cnfXejFMOK86yjpalZzA/5JxCKU8+5H3FbANM
sajVxYu0lCXbZUNFvyeta5OGNs+PVQ6X7qSAOgOwGFYL0fuUo4nTLMV5hle7w/8R
6tIdjKYAZw8pGNiIdsBINqF5WKk7yVMgbH2J30DqHZu6BAlqKzY2KfkUURwrzvuo
ywGNW5/t3DjK/ug/AmUwJpyBnXBUBVRHbPLkirv3fDbUzYE+j8kbEkT3UCPmRXlf
rlvVYZQO6a3+8OPHql0mTxT/++8Y1tnGE401IG8zC+/xJNqbMyGzj4bl9XqtBaTg
xF0I+zQjKN9DtbrKqfnaNGdz74lzjErpHyqxC8EnpRFVyCEHvuPiLacBwrik+lQW
62zoN3BMpUKOnPJeCH1vNHUH/0sqTdOneu+eK1zkJD71vO5ioyEF5UVnprxUD/13
AxleosSRiCxbS+hK6EWYFlmhKcsvhY6PfrquI5NnXWTWPblOXJLHyrzS5iz6SAlN
32v1qIL6Icah5uOlPmv25Y78gHFpXeUAcGTjVUcjt/YZYil9FSwYkY0rkaa93Lxa
zFri0TvtOX9MmjXha4zTYtw4MmJ0y5fLbdp1tvqMafPKQW89k0riToJuzTRQZJzf
hEOUkoVtP2PC1MteclcDeQyph1RJ16Ns+F1A3Fy9r5shwX0p/OjJhMPqnLMaGVcz
SFzbLfF/upwh8dxx9ndY1+PsNpY76tVhBEW5wunmVcooN6IMak3cQfhYTPH02Yv7
GRHPVxCFUjzIXeEDlcETAgxiZVj++tGERZ1I7e27bJSuKE/BqHOfsSFndeb3Q8Zk
ezPjVaYFjTOHyLRwS9nsbr2R1eGqwthZ/cnCYA3khpCO6wN70cbxuZ9VMs+O92UD
dpt6/cEOxReTGqOz9RgAWihlK7huCyzz/2i/aR9gkyA2u7N/ppS2ajFaD+omhsKg
3v4IrnDR4ykBIgrqsP9BP+tlm/kT3fxpBvtAMMJBOfUZ+Yx6qJuYi24hAYGrOg1x
Mvn2VM7DWlomVzW4hp5oIJ//HOoilCmKYK1LKxM+unwJtI8DlR8G4iMvQra2BVQv
GZZYilrsWWES48yLJt2HDuz57TtnPVCo9CaVl0BWfEB1McsFY7CAnWkHm2B9Kkqs
Jl+rGT3WpUhKGGwurHNsl3Kss6oc9OPgv8BvD6K+ODyhidnfSAhPxAtTeuY06xMb
xxzeZNPzQ9YbY9N6CWH6EIHSasSv+orYmo5AO6okM7QpS+8FOlw3shV7+ALJ2v5W
DNlZ8LuZh/O44cnW8zdNbYl6p6QPhoDBh8igXnfPrvdu4FNvbd20rPchBtmDf0Jq
Kh2zoCphLZkNmYt/h0cY93mxvQYEWfX+S1u9vBkZiCSCN3pvu36llIkExNUDoPNo
H54o/Y6QrrF4IfCqfRUkwvxAc+rK21v98lR23qzl0dJD0vSg8WwOCt69+G/AcLV9
p5OX5UVwu9HyFvSoOJTwTI9R/4sQ+wxrLCwY+EqRGKdOlBo07ECL9Qe5pxlV38lt
1/9blIWaLD5k4fQzbdpIcRLi0NkEGH9nWuLeZQ8mMpIJXFBA+ODmkuS0n+INUfZX
ZxyQ/xqQkTkF8xs/fj8XMlJeiwDLz0zD4l9ohLQOf/TwGt1WEHsiHEioZE2LX8nc
vc6nhBim1NwgB7UgD8AalaVtmSLjYaai2Ei/OBSywapShYQZJ4iz9N++AhIG69AK
ePhPFizTC069V1fam4IqDnlHB/N/2j2qEtNM7D6Bym5JrIZo9QcgOOzT6tXMhMgQ
sHmWB4U5+ccgMy0DgmJ0gB8i3wTItP2dACDt66G01RTIftst/b1Ml1FGq44cnsy3
uq25fGTmpLS1skZOqCwCghv9aebMmnQn9oJo0w2ZenmsKSHaTJys/JagiYuBHaEZ
WS+HTYhZ9xPleA3pDgtCtZOh//9q0eGtHkZ+JEz5RVKBi47mLyCJRp0srpDkz/8u
1G5C0HHcjQG2C/cAkHlxj4cFkxyxJrI96Zz8k+KQT8oUb0deg1Kvi2d5fAbE7Qz0
gzK2HCOCjwOmQ6q7VpFNMAXHqSXALUzsKITHHS18+OUwicndpVquX7aPxJcAiTj6
D8g/ruc1oMZrrySnn0X7SCL4qf4C81331VcfXdL3/oQ1KTFfwmLCujGrL5Ajzf2A
M18yR5nOTmNEE08cfuogxfF/8mjZ4P0t6hN0zi2gfp/YwTjaZDaO/OVwe7eqAm2u
+vaL2xg9oUsBzrVJIvesyxye6gWxHlhp8osD6JeQBT8kj2N4kfEqNe8k6GFcWfL3
ar/kNj0xVB46fBc27H1zU2G2UM7IoVTeCYiyMPaR2ejWdXiLniQII3sMSBqpNmLl
1Xnf7vF4aKmL4hfZ4QYC1PNXd576xhH4lmx+cp1+DjlWg4IP1RvD9b2PZMyiDI4X
o0t5OVoo8h3d4i/GcRc8aI8VXN4euJiJTrcSgb17mPm4oztpYU7L9ZfwsCcn4CUg
P+AaIicBVbAieUsWO2hypuvl60hnah0SXANKSRkNlDC+ExYD262Zns5vWfTkeZTI
SA0n1/ZeM8ImcIBhzI8HMwg7dx/kB6tuMNhWrxtBq/kzIivftUgNvTjW71M2Yy7h
qputnNpFITBIRi/fsVTjOAZIDIooH0AccfwpW+sVgYZ4Cenh2auvHVZaOdANS8ZI
Crb1jFg07ROfcPuLC/9CUFh+PGR8q2dDSuzHtOHdqJnJkDAXx1oj4l4ASiu3gLYF
yme4UV4HazeAdc71dE4HZEuV8DS49scc3CDHPu/K2FNqFq2SpDnBIn5mOSwkrqbD
T6J8CvrYxw9PHsGZMZzb+D40f4sads1kkKSqDR4lD0CXn9Ze0QENPmsDq1Ma+1Hs
368UfMwAr+ODteWZmwLbgiEVG8ZpOhy4jtCWM5OXTKSDPpgLTWmoGSGKMW/oLvFn
bhrBgYKRg1Yx065dzfjYiccud+fvEms2oLoeQlyFL1FQ/+thR7uBzRBGe93YdbqK
Fk051CgVs/hpLE0R2hVLy9ASqwIAs/IWCxXMQp1LejFXTY5o709PwCt8zcpjDeIL
aFZ39Kd5h4VVq7OB+2jYWaFL7sHalcIXRuePmUvPYGwk3rNl86b4BiHIFE0PM4Ii
a5Mz+av/tIwfLBRuM0eychTpY+h4xBmam0QuG9CX9e6dI6W61hHUBQf338MunsmH
vC+BK4tjtU4WzOvU7tP+CoKsZ/z+xlsWHYeb6ptoi6cOb1sGt73s37vk8AMmN8fb
7iroAkH/9hTupPGb1Vuarj47/1/4OR+QqGE22i+bOl5afo1QeDLY91B8dRaB9xmv
KCRyUMwvUuFCIOkn8TKH5iPqRu7sFRHZc5Z3CJry7rWwmqfTgV3Lql/dmWJuIqy5
NqWtnJQ0Y1UKFLsYwqPDOiJAnLJF86LQM4JkcQ61PJi5uyEj+WLuGVdrNNjuXHPM
n1cHWOFa3lFkEs/dGo10iDlyxpwLgjDjJlaSabkN+yTpD2Xf+vcYxv7uWyTaO32+
E1ndZtxDvfZUhGuAXjg4IEv87QMFI2alNRRLFrDXsHODc0LxIE8sseP8j+lJ+IKp
PANE3kbDsxcOQ+ORGhDlqPzzSvyfRixzn8RszHtiS2C0rzuLxK0EAdQ5+BGX6AYa
krKAbfXIF4VUcuDZqgGRrULdY1cSwZYanQwoGD8bXPdVaU4zvDzaz48kyFWRG2n2
PHRU0bhQs+vKAeP+NyOVVKLUyPvn4D8PgaAYWcEIjH914KIGCZ6PM2yULVEY8949
gwH5mfm0ReYEzlD3BfUcnzJn3GX9EpKTXvXcJoclV0X7yza6Rn2yZzo35TGPj//N
zp2iN5OsqiT61E3135HWAj/IY5yrdbnCLHX/3xPpXNutSaFa2fErAD9+y5nab5eL
9xtNzV9/++RFhox6XisFRoA+Z+RV7XABUGxi+iGn7k5g1KmP//7MjCjw6zs3SFbi
U90tv0UN2Zhug14dxjMgqkTtupoKo0TFsDeh5xkCy5fwEemHlfAYFeQnmT38fHEs
zIp5QIp55/ROAgI1OyTNM0+MLJjD6rQTgET03wgbIu8iDg+D8gYC0/Sw38F6s1xJ
WM1c+VZN5TFaX+sL+wypHgiqG04577corjOTVQVaUjAjIu8icIlvmwZuCqAHnPTx
sixK1NcPOV8Vhbdh5UljEN32meGbg8sQgob1UeldcwZEj611rsift4uqZk40xmgq
9fuO0Jf+sQTr3UeyeYCQD9gYnc6BcxvxLguBsAfiQZxIXKOU6i47fQEeFmgIEQiS
FGfQrDaxSyNpxmsPgOwtF1mFuJ3M6jcyyOMN6Meg0anQg6Gp0RKL8z/suAhZFWU3
D39hG8O6K8t1uMXyPS6xncYdLQZE2+RXs/DuWqfG9wtNfmIj2/iO6Ok4VkhVEyKQ
XB/Wr3H2Key1oemDegPkpvHYwIhaIyLOzsh0Ay1A4HtVRpCgMhpzBxq0MMXLy9bd
5Ulx9ynZttf6nDbJfnI9LtLVMYS9rxv6T+Lk4ervdiZIZBGnFMN+DsW0Ehxwq8i1
0aKrXADd6/lto6+l0m1dXp0YURZbssBTvezZnAV0Vv+B+T43MCURoXz+WzWXl6NK
T5MGcRE/tZ1bylW7+JS48q2Eot3FNf2/RCZvBAVNgrCg3k8pa0UmEGVcxdvxRhPT
JA5o17pYNW9PFGLgAmS6Ik4dMUXDIBH3NgS090ClFYrLVctMqShrc0ozG3f+HsxU
u8ZgZdFl3FX5sfKfy+gL1Y7okbpVflvCMAnErPENEMRryPEXah/TxS7voq1IXJia
oMS3HkxLtHRAQVYrBGWcelWgib9RMgLxk6RIYWwNZ3BqbUzYPPTXeGeOuOjSZeog
Aterac9xBbiEcB/MwUGWYJJmB+YF+jgdGL/Y+D9HWKpbohq5z6qAM49XCA/1Adnq
79rzA4SZHO4bgtuj3sl0BZc0PF4Dzco8qlFeVCRbpwjRnUSQUiZbemtxZxQPYEpt
uyPYPoBHUO2Jod34+csozNAvy7WL1Mlja6y6173J2yu8swabqIjKyN+3FBRYGy3z
qqAZTV9/lYfLzZ6SxniVh8GcpTfAyNRoesR2rXKYTWWOwlPdrBIvCqJEykQ2KVF7
XElPhK3TKjZw2qG6vgwHOoie8/6RCpGEsD1YEKdLgUlnBA54hae7mF7ZaqmWUD9g
WrJaRHD4laGTWlq1wpqAegBdJ2r4dT+cR1k2+nUB/Uy0rk/Ze80oUqZ9C0bg7tkB
I7IwQn0On2+SRuk0yR0LCPXvqZYA1eV/QE3ayhCJ7IAXNkXOj6uaTutffqss2HMY
PEDe8il2JM/WA9LuztyaQntkSOihhggzEguIVt1rM9axpKC4QkGMIXiJxGlwdC0c
CevkEqOYNbApYCOYU2Ks45LqDXaSDyY1QdMfy+I4EhobT2gPbx+aaCn/3dhoUSDZ
tc2gsLQjia95iybt2U88WDCeYRS/oHErt7W8P5YVUQKVpDXlCSdZoHOD1VDMewYw
+GY5BaxocMzpfvIae/WmTv8toc93weRA67uyu0iAgI6y7v/K0UKZJd9QV12HdSjD
pJyWq7D+p/5BKS1yYLXd6vKmnWLjUZvjKRuD3wwqec0ipCQ+4THtJXxGDWWModkg
b9JKlIbFNC189Z85rfKHACzWKf4WxehH2pR8HnmUOn8Y/RM4ZHUCwdVYGBO7tugM
TMZI4wPmNrnFfVjI0ZhXH9WC/CQrIXXf3EsSBdnXnMnOs7k2qXL7bs8ClwbAgpjv
DaiQo3RWxvGmfpuXjYgN8uyUWM+kidxT4yhFmECafdRwX4mlRgQKp2NZtdVcM56p
5b/E9bSE6ycg69cvtYWkwGZO6zE5onf0WMfppO4EJMyODtk2zXYJMKiP5pWqDlpB
DO8yXAVEzD8TOS6X1zSOPrB5moIYBIbyN+oYnYOVDAlGMeKaNFhROeeY3gjUVTiJ
4bGTlbLAuw4D6CQBDtj/riL9Oyyfbf6gT3F77FOgixo9DptM4vDClEFrrGybuPPd
qJtxY7C6z/11sX/wmTIgXNK3vghldVQ5aL1CqTpaP7kn7jgwPQE1w2VGCaSnV690
KOy9dhml/hKjTS1KFKRZ2RvCoq26DemUF5jHnuKpWKvVSvEh/r177G7elMEtxRPP
4ciGgwjncySqPLcX7xj7xnwTekeeNv4zsJFAyRNSs9QuFe2wkOhJi20kBNkRnV17
94N4LGPSBQBzcmXfNJb7rVbG9F21u0Cz5rF0iZmfQLB7RyUEqwKcK2F4cGBJ8tmo
N2rroyZ4r+nyVjHpelCfa/9CBb/ALEIuHJjkpJxQKILhcf8T8kd9v0voSpi6xgsX
GdmOfs32+NnLddfMY/7SH/y0rHnIU8aOSfhY+kjg0ju25LPlzM10h8/FRmr6slHZ
2uoHKApp4ig6jHFuxSaruMccGpONA7RR+QLQ7bA4IZiCpAFocLthx3ASvBuMGuL4
yqblTZw3laN0o/ZQmXHyVm0k60SvxSt8BjZVfBSQEVenINSshES+I/RnD63pfS30
pse7GXheb1dMKYqubVCoJHTkIFclTN12wrKLj3SKqmAN2GjGPxVKT+72ZFMBJaTX
OWi9SB8cqYdRHTOXeR/9YY4pMlNkaQ787jIIJZx/NUbdYRCg4QWUDwWJOp5b5a3I
SA3t2OfvR+AWfKrIhazCA1S8X4LN2QlUGVELGuJFRpQ5/fuyPU4BK0axdqylP8Zh
29kF2jsxKirNTp4IeWzT+I0jKoRdKkrWylTabz9oavYHhZ8Xl8hlMpTLmwH0dIE4
6IIOCgmbLaiPDxluyBIFqUHbGaj9AW6fkl8ErYI57jMKt/dYuh2QlRiT/y8Ovm9g
oUJdP6vZAlLDMGre4MdOoWvzRVvJ1P/AGXPSXXnaQXvrUBNre8+xRNcxTqgJYImC
+YZlAFP2qRpLJp/1clj3UyKr+d/3LmNz8wZw++Kcubf6IbHkx5cos5ZzxmM2+xUg
Muxpjs36VV9JC4obSb2nKMpKR8e5sqBRQC1rgpQfNMsftMRXVgjIZce37ymlSFYk
RRM7Ql9uS/BJUT1liXGc0cFQaTcUsPmhWegoRxNkewYzUupjZiBEz7O1N7zJd3oC
3ueAxmGdAlyNlgOBdAUeU5u0BLD8U7B2ICA6ZhfwuJmuoAXF9OOW0pchPyqwQX7s
s5WrUzA9NlVDgAFBnWXnhn5Pp4bG60QTBIKIoN3rFc+WQPQxI1AgttehnVh6xbVr
asN8O+zdAnrhW9VYCGjc3FCGsfZbGMHYnE83RiN2ejDV/weLwoFLEM0bfJM/q8hi
06ISEGKhB7o3lzkSO/BEkQpnT30K1KiUO/lFuePB7EUswTRey9qUv7ZtxVOXJ3UQ
ZIujeo05svCvKB/CLXMjNUUvKY5YvjhVjLAdxe2+Gn4SoaF5ZfS7rYLV57dUux/y
OnCIjQRrC+I43vpUxakmIwlkWC+9CbEbdGj1THAoSGUFjoaadVBXAAvxVt94O4Ir
Q8stX9GQ9zC9t/qyd7c4j0kwU6aSQQFh9XcxIXTh5DPmCulzUgaha71Tf9BTTeG0
PcM0IBCm7GASWXx9ldLt4oWhJbMcaxVafUeh5aB7RrbtG154xxMj9NXJjHRliOm1
SM8CXZkC3rs1/JNZeIZ+F0RurLiE6iG90Iv+1ocXnVbbC+euVeO4/dYdOmeTcpXO
yYWjLP7tKYSVY+J4Qn8zZKECKe7jC+BWaq38aT3nOpwHKqsEj4T2RCuaGBoT/QWa
ZqFY/xeuNuvsMdtl+7v7aksbfu/AEzN5RM4NHT/jWVLDn55Jb5245ius6e9Y34lM
yyoftkmwM3OsrPdpyZDvETr3cXDD/j7YC/bKVTTqsnR2RjjNqmIcWvjtBlvFc0++
33a8EYbeBgn7jjCn4sbmwSrriU8/hHxOq9JbwwoxJiHCmdgVr72ElBeYKMH7rot3
c8hyZHSFdx3oschsEJYfWXjF0hONUdXliQW0fIf6XrvnkgXVeNX0J5AWtEvxQTZJ
y9Ui9uCPiLNwurWNIpbM2ZyZcBYwfmznWBqc32rK5iIAUc6D0SLHQ5sT0Xglg61T
bt9XkaznZQnTssnSaQdqA4jbdFTEUZLbmuIzpiSv61wOpHmDJ0Ezvm6f5ARA0t8O
DZ7a7cutuD7MgtPCnF2kieGGJrzZDuvaDgd3hT/IfTXePeE8zoxSyhXBwcr2N9q3
GJpnQ2pjoCS0q+6YV7que3UqAe7ittVPZEushhaQfVAyu1ItpP3l6ufyhrXpvr+N
3lohsFzADHFszkR38K7bWH4KD1yWZ9YtjJKEXrNWygy6Tgasnzca+6G0CTx+Oy9e
Pl1UI8zsXZuJoCPIYXRhUBi86YzeJNCj0d9v5ixtJRRzypNMmhylNTrdSJ1K1gKU
XB3pKGMDWZvIMwg1UrzKG9phxEH9g2cAJ5sbqkrduKlpIy83+98YuAduuPyiUeGe
ee2Ku+ejfdjetjyg83iK9lZURnLquz2A5uC3hyEYt6inIPYMjsI9hGkPnkkpaxts
2vfJnftW0ieCIDlpEsNnyPjTUA0J4GiBQnT/ec6nGKJmpVys03VUfq/VL9S5259F
JeJfO2ZzOMbF/wxubOeAS23VHMnWPfBaYdlYsvmtU2P/haVt/HoOA9lfS7r2nILJ
UTyvs8HiWjVPyDIAMC0XDZGx/EPXlcDMJ49WAisFm5WFSA6I1ZDurup2AdA0Ef6C
hUdQU5gRupKi7lRdmOIvu71UaHd2jhHLFK/oc0+eC6VwZIZRXaaP4BiPV/faHXPg
ChCYjM2bPI0ZMMpHH0zsB7jgD2RNWFqLK0Fig72QChgcdyX2emhFerkVOoWlZm9B
dlCXsXx58Yrr4x5/7uXyD8tIOmUNOhKdzad2stDdjv/3zxmWvwnaV3wlaHbXO4rY
3uQGjlFeaYL7qPDzAkmUjm4TtXw3nVZH0xihdv6Sf4ea/fmuTm4cziQ4SSQ+ldQk
BW7pNkkLc/GQtAUV2Ojofvv70badin9L7GwUKq2VD0FZfw5H2ifVBETA4d0LNtpW
1TrpthsAPSeRS9LBEJE7jlg4BWVYo9qZi+/oR4wHYK70RiJRMpMcfAK5gmP3hYM9
pCDmvHrcPJC1Ca97jEwY0BzU1nk2XnnvZebTNwJPBrWP6SJb6qDaCS6Bny/trGCG
Laif61tjfaqVV14XKb8nd6tIYfTPPuVpIViSoRcKTm5lHv492A5TPWyORC2Tyd82
XaOsTdECcoU9cKf90B/77C0Ia/LVycrJ1HWj22S7VkwemBctLbTlJsYCfbABvbAR
sn/PTx6jlNBs7BHZf7x7arVpWh/MK+5b9y+5DMZm5JVcr8XVMe+p1QLxqsPyUq/4
mKI8ruLyuX7siUxKjkY57TLZyxoeFE78KkcDvwYjI3H4EcO+N7sr4nAxG+aeG3lR
7loCJbcchyBUf6/La8+KikzxCbMXw/PIZNWZaUAkLc0bkOJBByXjjuwaZV0uI7Ox
9iUzxzyULoybgvEkkuNPn8yrkKGmPyw8p1qPrOanfhxom7D9fRB43Zf3E5q422xU
Ahsuhw9oaS481Qvuhf1rDcJjZdazUVYobDhUYheuiHdKS9iQ+YEHfY3d4rqaryEY
iDUTiCkRHzAv7pkIEsUVmP+mbu5A8/dLEKoerEtn/PjfoeiR+/hD+7o3bAA/j6Jn
pIm1gZVegWn763La3KwNUJiIHZM+SciPE/0ajyJlHLqfKBeJKQJ9bae9y0Vo3tRw
JF9VKYjWp4uOH8ym5reysHYjPzfnVCJLGA4RG/MMngp4oJLIDR0GezJI5pZ0zEaC
ZuOc0s8CloDhvd+YL7vYMfIudL07mpwZZSexz9DEnVk5/91BO+6u2yNOmpwdHyjO
C4ixr3xbRpkjFV+Z8AVzLJ2GaiylP0d5WbZA+ypqXTs+69blRPTXiYr4TeU+IKJQ
pnJnnQlJ2o04b3zA4HtJCHt6AM+7iAF8aWG94ohd6IkqaRZx5cQfIxKpLJCvGI71
FqQ0H/5EIn4Px1VRUpWYId7kiwlzl4M0v+VHdiVx9laivL7r+fEifIkdEHHBXpsw
zNrJRriFW1piuQt2vhP5G7oQGxiR1XnkwYtOFpMSWaGI42f6ClsWMOlZAAD/iMPN
V+s+be4gTiZX+APU9llmziuZAU0AP8XQLaF1USzPk7mpPdsAjLr9NkXwp3KeUIuE
73gE0KRVBDY14CVbM1msAAkG0s70jOCkfLYSc5XzfqE0W+z1ZAtD9LWDOznSNB7R
hY8nxL0tOLG0i8qjkF2e7h0wcc/ncXd+XbnlalGMzffhOPNAt2ZDq+jthm1mQ6bv
ILyODyMTQ1J+5kuoHOGIh/QD/F2VURE0lPtYB6NDtc3T1Pp7TVtI7zlFPMdwnPNM
uUJaeV7LUy1UiRzb4aNVTFXqO3MNcprhrmxzpC0bxD4RHqpoL5pyUzhiSnd9O+Qd
JLsxoTPkf1GbagL8WW8zF/9qDBRyPOKU7EzjBHh9WStYidTkT0lr/dOQxrEQqDKU
8MNTcrw41clwjQ4slmOnU88rkMvoS+3Cf02YILcS4Cu1lZYqO3N3al2wyW33UiXa
wNocvCQM7qdL3SnrPibkZKSiByV+7ph+mvxeWBpezvTJ9MHMLTkxmU+lNuv99Rwa
kMv+3rArYB1JkTKicjgmUCyQ8k2IrYaT0ut+cCsVCf9XKpgyRAr/OZY+qf7c97EO
u1sW22eSk1UHp7JSTh6A4VH6hC1d9HcD7VPRaeSknsQ3Zwi/9q4fKE8OqZgzT4yr
ttdODtxgjh7N8kmJKTEBpNJV8P0vJbz5DAmJa5CxRaURBDfAB2LmatmRELDn15mu
9qKdKIEGG/TzCzudZ+v6BoSrsO8UAxStdIgk22LCLbhRMcRZBoyNBkwHmS63mlTc
iFwYBhFsp1YNI7uXJdpa1pTaydvQVDfCrMLNSYJOOq58gXAzM/RCg/cbxd7gKfAl
MZ+FBSUY39XA84Px5/1/l1+ytW/TzrZ0ePem7OKdF9atsZqPjHMnY1U7zJm4TBCq
1fViwLwL12m8Z+Viq9ae/KQFzprHQSNfa3bsNzD3kWAVRjt4C1g9wqo7QD2kpCrb
5zMTYo7YHtADp3E5rI6zesoNFiene0dm2KVV864MYzIfoP/tuSS2KvYTThQYSlUT
UkeqhgnM4CEJBCmJ/wFF7ipBw5VZfB/FqGn7ch1WM3hLUsRb4xMbLLN2dvXvf0CA
573YI8oeT05/zr0eiLXgdCCqNTFg5mpLD5yBe2dvdN2y2GyPQV9PyDiF6x5mIVCE
uTpcvTAbm1J0wJ/4madLdJQv5BjF02CP8xwvC8pMVxFENkp422bcFbZ65RlfpKhi
ZAj9bhcdZtSMhQRv5fdxlmxzaqNYZPuE6AciJF+veSxBRonJ7BtnZFa1xA2/cOQG
/xVkYOvXtSz5RkDL2Ux5se5nCnqRqnkHde6fLfoHGzqfY5uELbXgd7C0hvFvSH2+
wSnobn+LTVsG6A5Z6JmYRNHzJ2NC/7Bcqbd81rd30ItrardkMqBq6qtGWdYWdEwU
qjRSscFBvYwMcmtoHTkPrssL2Ir4nOGsWF+umJINcvtrSHXNvHqKRBynCSq5vXHp
zq5s4Ezx9caV3PEJt1o9UNVDnz48gSk6+1J/I7pTL90V1oRKfo5poBQFqnLuPBFv
JdZFUXslwD7YnL5t9AfWrX9sVD48Hi8/6BSKTr39HECDStLbtLsdnJEWmnVwaUcS
1bGpSkjnnVBrFp4XzfPZnc7ALDclPniE6gelRSvUuuVjHaP/rRwwqp5TZY478N3a
BEw0+HZHUvf/rBPoA3f9iituV7HuCOnlTb/keW4pCwrcrFTzRPc3iyYWJRxMlU8h
zXO3/jNmNNgbAyMGIMDYPqgw+N4wvIb5XZdKSUMykfOBRKqSnJzfaOqTzMtWl07P
hARrZv4xDDpXutdMr+dm0uaR1ThVA/PebskiLu3oyHj8EdO0QCnMJRhTzJE7OZ+c
gxEGRItzB33InKcAz10bhbszWjSHJf/aU1xC4yCErY9E/dzeiAR3dj0Mxhcr3ZxZ
CYc4lAVrFUk69Ur6EyFi1AeDMCl+h7CJnqZA4qxqrWGLDbVbelHuWrR9lpCaKOwq
0wsAe5/gJH7Yi4WXGoNZ5yQIV+TAQbwa69m9pIMsWmag3oGA+uQFAIfBafgX5U7z
Tag+59L7PSAlHvHK/Yht4pDTl2caww8P5zUAAm4EPuC7bvGZO1QWgNzwgiiTRaQH
UfBCEkHKt3yD9Gcf9KFx+bt4sD3DFskQYDWL+uO/Bmdz9cYxHMoDEzj0jpSr7Rcl
zs36HblJlE7Ji+tRA6vB/IkYO/9SpU2UCVD41Xqbgx/b/epFhSO0+n/XvCVoMWCH
ChpsDSrOBl1lLVNywA/30HaxrE6Ug+2uaZs7I2SkXd4Z0c0vx/3gQcLEckyUJg28
WCso2OKNyvaWhhBb/bOvoAVr4zfYJdL6QFex8uaOmxYGhQ93gNmDOZ2FU5zJshQP
ZBFeuK0MUgK13XnMUXT2Eo6NHRReSGSvRBxLYtuuJRdNfEFDwG1ekfM0zPk3QH8o
wSQwe7sumgpqdUEk86jjULZ3IYDgyHTCdK72jdUcz1W16Oq1+BCKJkyFh8q7LU0o
8TvJSE1weQRIlLl3uqvNktgHEhLnPiTqb+FRBZV5kLjGGMG+Bera0NnEN48PsPiR
/Ock8V0ppxk/PoKBDLMcYcExohSuCnaWDnzXL+hW5zp4G2P2uUAgikiRSTEjOYGO
0tNEXFTWBFgdZlrzCqsdkXluoeQNG8WVnZYfSAEhoMt8SBGMcQSxcabqGUbN/Htp
Wxy9jQsw6zqsl7a4jcg2DI7lo0xAjArlJJhWyc1uzarPvXh8bP4W1TBZjxByxsRQ
yPLoUgw9EHBD+Vj25WZpTMSrGm46Hxtth5MkHG6ezu50c1MwjtZkvPWsL2XFRKRs
nJkOQjdPemyqTHuyNRb5DiiiUEvmdO629TAjEjKuP/x5/duFhABoyX0wPm8T3g+s
jf1fDvhnpinDZAHxY93u1MIKwYDbMMoA4wHRb+ejSmy/gep+RwPuR89Sc78tY7Vh
nsRn4cWf78yHxVEb2/46DPNOsR+zvLAR/nY01bgdfgrE6/RKAVNbe4osAk5A76Ci
8RH9FlxR0vdu1O0SmUrwzrR9csf5eZR4LpoadeeGH8GARRf+04JyhT8c7XyNPsLz
IC7sC0hOMllxdGlzNCXiFYKgbblrpFfgtmYtOrIUXJEf7rlAXzPlthdclwhNrax1
5P6AcjP9oLnuqjXg8QJNoahG/K9FIfHHKLvq69oEkK1xgnMT+uEh0gib3h1tkqDV
Sr7AIE2M46bPV+y1QDB5bVU7juwjmfoKvM7j2WAdfmVD/PJNX7s3HySacaKXhAoI
S/6/4RdvS4rvTsk3hDUVkJbH55XRs7hocuGnqTrt5uKu5qO0T4xpFhQhefbOeLEk
nBOSYzP6eXoZcBlOb09gdo6Jvg2tFEZpHuN15m4rlK5w21oh/V1dOD2TznGAgjYt
A5V4WRAjVXOy6BR7SehdidN3PFandW2bnaxdK1QPzSQcgXEQ3VNTpJi2HXWQ+hTA
STNGgqDUzIBB/OfNwwpSED02rXkDRjzmJeZVxKa2cAXbvYjPnJ3/3qduAbMEjhkR
LO1w2u2WveNT1MLOW1ugKcQGbqeYXP9Q+Af1A2HaVKK/my24rMWasuN5+NbSRA/V
MUBWC6oLza4O0P9rYISCJfa6dL3Q8nDsl1Hf5dxypKeP/WzonBvRmhqOjn+iXAOC
+JjILTmGZMcKrC5rp6afu73PhhGVMV6oKI/jEm9E9QlTyxlE9DypVqLHNDvZcFui
9+HIUGMK6VqmCDMgDt+bdqLcI5ibsCs62uxVplCdQar+HuGe4ficNEzS2gKEllly
yF+aC8DEINc8apVAVG/b9VxC5ufQBGY3B/9tOEYOA82GMbzyGnJVpRes4kEi88VL
LtR63tqWYIbfCZPApr/VB8NRBzl+wYBhTjmQ2Mla99cq/bySrqq3Y+LiA/N2tP+s
LywSsSty4gMtw0AtDYhzfNP32YBbGxC9sSaIRbnSiHpqDYS+PoNIpMUWAcY8oxrP
8xu9t+mOjTN7/YjaMOXK7S7RXHadmUCb5RmZ2d5L57LC8Um280GmKCbNQGGwO13v
aciArpwzLUvbddweyXEef2bCCGEw9auPc84f3I9ZCLq9MRj3r2zfx1MKWkq0NG+Z
tWWdnGLjYxH3IgWWTPxjyP1Sz1SvkySVM/AgA4X9BdFjzu5Js1nEgHuN0uGTpT+L
7q03LF1USHi7k8m6pSkxZes1jA7UxXjE4HLYKrV6qVCdfl7/UxxwiuuJs3zxjwCy
63nvZU3N1HmBJsCroXKNtM4c1o/Rdk7vGiRlFTclYoh3F5L2+ddwMKf/++0VXTs7
I5aFfigkomPJzs9DJeX5tBqJ7Kzk+T0YHhBK0jDiCcNNIvU0v6RG1P8fiabzyi5r
RWlyfbqlcSCGg6+08FD/rrYzONfvj+6kJxp3Z+YQ6wv79hab0iP7KMrCKBRmii53
gsxOJGg7v8qJ+/TwUtxZVU6uHrzWnrGUvVm6HAURCKcnQmOpby4RAqaJlj+3Kjqt
hyvZ7DnX54o/6X3P4nfQSV3yR1LXqr+i0el11UqHz05Y6CGtDxI/jXD7y4P92YLw
B7jRDkMUahX5sukQCulfexZ/4/YWuHy9ssqajqh2w2BQj4RD/q7IQjR7pwKPqOb6
F/vYeQBdZjO6C4eRv6aoZx6glPCG0JFAtrW8yeIQ+1VKwdwN+qwq9L3cerJqUujn
BWIZGTumHXfpV7yhx60/T4UYNNLXahtS0dX5vZIiSrgC4WSJZ6O1Ag0Os6PBDXed
Dw+ULpJHjT/58aCR+qrHmOWIMppottShssUHQGLAEZsgw2LvhNl30jnyKjJVw9CV
EHMjVi7CiRu7ZKHXvO9MDVC656zTQiNIRFvuQi4N/cM82de5nvWKV4UMUF9y/+N0
uM9L/tWS836Yb0BUSURqxhjwW4kvj5v2P5kVdgnIMN+fi20XFUaFZCBq92kI3l1q
/4VWXGUO5SuZ4eIibhI36hyODQ6q4Vkv4f7L/r5gshN4Z1T4XJZxkeXNsU8bOflL
8zJYj7/ycuBeM8dr5zPnXcP6uBJ9sE5WWiaOSHLZpieAQgD5cuS+aQbfX6qbJVp3
PsicxG9lK/5x4uXy8VGBxxfMnVD2LfAYSjLij5I7OGJMgO/1kBvsFPZAfqKbdxMt
/lnzl4o3Ccj4hTK4hwxLMlBCYDZEhUB+w8eFWqJu/6g2gx6bd6YLdXeKvMZ219ut
veLZ7nvhI9JrLp90bwcdoMmAOXXSec01tN+80K9Q5v4VNHHW3Gg7YgOnTHoNzSjB
J4rhuJnLqfyBhVogPPS9uWuuYdCa7Cpuvcw1kGkBiJdRMsrSwVOkSyzzWznDNBsm
FKaZJ8/Gb44uqF3Db+D25Y6bmq8DGD3bxN05dt0bZKmkn7aoCmp7H23VUvz78UJ6
t7tt9MpXfZZ0VeO50YXvk5jnZJPdRitEw6rQURtFmvC9BNcZahSc6ccTab4VVj6S
67uEM+yA40AwUzPqw1gp4+b4lTWGxFd0ERxX6mZLPqMFAaGXID5svcPjGIaK4Saz
P80JAjAKuLM9xSt6hiyBPxE88juIgdp0O5u58DbD5XCl2C/sdMvfy0VoPX+ew7h9
4VzK77qkjil+eWlGsV2q0NCepfnnpSpQWhQe9JoI6jf9vZf5nflXn19vhx+E52vB
pdSEaXnVtysv6f00JED0YOAxqNoGqEHurVhfioKq5Pxt5GqS5OBkx3dnu16Lxput
H/2n7Wxyif6ow9bArQ6p53/EYNI4C5WxFWarA/AGl63qCxECsZ4DA5Ihxx39Vx/t
14Vopb8iZH5NV2C4/upZgdeGIJU6c6/zNbmYsSIJMkkLVn7IhY38b7WoCPfkQ8h0
V3SPhxWkToRGTR9paObbttLKIxx41KwcCxjbdGbKyyMYcMAD1pKgfg0rp+VmJUjP
09cTlAFCQV4tLJeTwJ6WZO3p1Zmz4MMQnF51+CpiMEIuYGPtmU1yiYq4Ug5S6QCF
e4dc5V42o9sANWJ2VoI3xtqRX3MmgZS0w6VLWyLNZGxeN7uHSmbXFvNDa/UnoFAb
8GJVxi/iRkQuFkuvObnAFzOXeenic4Zvq1+MddUf4bdxF0XDvvL6wc2gSy6OLUtd
ASKq758dHIVkOGFbfJ5wM5kHi66+OotUTSkP9F2SkSjaUXx4n7xflAgvbCggHWq8
pNeMjS4vxBlIfEeo036g9STO2iZ2k5ZOJkzfTbk2umI39YeVQBocObkCoTs8J1Bo
t3EhNBpaBv8s3eG5056NBTBpDbSYCJkybVTv60nMtO/SM4/uT7ZYYiBbqWP6shYO
oni5XF/wdyE5kudKAYRz1HvSssrdXb/OkwT4bgiIR4NX2GG/0PrNcyjEpkS2TjhO
G74kOdtBW76Exhva5sb5PpgYwfLHlMXMYvWO62CSJiqKtIXPBAZV4yCC9tC0zHW6
xtKWoo9VRhsJWdov7SBqeOA5aIELqAsHm3UX05A36rOnL4Gw4NvgKnUW2l2u3BFo
vmR+VLSHoVOXtFmbjTnfCcbE/WnSpCKd+ayrn+CDk9giDjkDMCMGtnd0y0pA+Rm6
3JgtJVsnbQWDxVBE1N1+JQG3fg//K4VZ9YBGrf2av5xC2+UtbiOzC6gjMiexLpEa
PGJVsyAPcwQ87U1g3M5YzBzBd7+o41waq6ifcjwR4hBFrdtX+pf1aW0u0VT9xArn
M78rDuWKO/mqvo3bT69tQJbtUbgYVYJijyGXx/aIYbPyJQIgSD5Fm/kel+KutNKZ
r6nibGrP6O3j1FnKC8zK+LT5TfgbcFIPeYdc5a7kAQ3MF6ZgFDDHJAqF+mev9fQ6
Pcnt4P3HgAggewpzithzChLXTi8PFpz1ljX0/kYPnhYRHM6ctIp3KWBYVBMT7vUO
TTGlhf7bYMS/X6/DAA5sHmmJHL9YUrZx0X+fBNpffyfJ/LUJJpH+iPk3Zh4EKN0J
vcARf7FGH8KOqDrASwWwLjcBHiQux+t8MlG1HfZRz9NiDlVK0Hzt9G30KLBvbAc2
uhg/8vnzkcRZW44R8+GhUdwuGAChcOA82iCxAdKEgm/N9GjdvO+XRW9gQcylG5FQ
6uEHEhZB4E71Ph9VN7gnrpDekD9ghkQCM/sBw+6B7wSMAEodtszVdjiqyRMFERnW
9vBBjFXIz4jwaLXYMK6qDP4veYtp06z68JBUMcOWmNJZ8IbqVycnhmI4clb3JlUP
1w9C1OJu5t/Fj8eyS5VkZOKun8CiVgcXS3P9lo7//Mtx+S91WDNJbQSiWTXgj8RS
oWCY5MxjHwmtjZPSG6/Ks4mYT+k8oLrxwNXd/RywfA5Nnp8y/HdAAa+oU2Fgsofb
3kK0s0H5bS/HypF3l3KQCykAx4e1BtbfNAiYWNvEKYL5MoY1mz1zCdra9/bjmPO9
qy/0TpKtdWxIaolwrlt724Jz+up4Vfmz+XJ4tD7XwlhZlnXnH7TP69TXO3ryVn0I
NITTK72wWf6OZfNNhBJV1hu1EPSw3xu8hI/uDI9RfmqodBuRpppL6Be7WMMt+DCl
brVM+XHIDVFjx6B9FiuhEgijuF1l93rsNDOIHZDIGD9g21O/7zKpFKQmZKikj2h1
e/20aLUCf5rhIJlQWRRJPCVgjQVl/lphOl4LPpIuYbEOTsiaStaS6Vi1NRMbI2t2
PAAPlyE2XOVOg6cBEthg8b0xRjPz10UvncFYPPJoxe2s+HVz4G+L8kymMRJfQbGL
HBR1btTJyIIkHZJ1DsXoj8nTkY6db/wq2xTKI3+S9qhbg8/6vMIInYZIPgYQ5sqt
Nv0cyMfVfTfYOuhLIC24Ecmqqz7DxGK4sNJLZ4+UzySadg6PHBDLc9M01BFUJX81
YnUJA5MGDehfcn0kuQY/fvPgMTNjy2TcQtuNqBxQvJEDeBGYHfHpY174vz1r5m4k
l0eKRSe4MB3fimdcZ4R6fcefHez80WXSNHVvPPF0JkY08tu6gZpSYIBuSwkt072V
/PWlkS0hR+jcVjO+LIr8tPgY6Psqah3tC9Zd8IKvzsxf3u08Mfdc46bKOi20Fw5E
t5qJEokqC0fdrsSbGsBp+209ViYFlfi9DCxO/LY0nUndaaPkInsvWYou+wrUqIbi
f547g1dbFmmcmvuDYBvSBM3Y29pnYfQT6+fReatWqbieXb9LXpdTAj6IhK3UNMo2
5dDgPjbB79BTrMUfmFajM0JNkSmj7SqVr9+msdLzE5NuZDOjqp/RCMUB/Hs47QKY
CyftTrTfSEROJeZvUig0XvhAEY7arEfUb/6ggLyXjJcodbnbJ+CbspA6otNeJ5lm
O2FEqhVForQHh3oRzUoVsmJ2ifLeP1ThihBDUUmil4ghOC04uq6snMeFPQ7LW41x
VbXExrn+XuEYQRLmKBZ+xRCzEXKudZr+RGgWBH8lp5GcSZ5MIuyw+Cp7rQUm5f92
zkysfW0zfs3WLTIjqupZ9K+ZD6GcEVUtgSV5lW5lzN/yrRqPK2Nr++oJ41sEV1vp
sVQc8LBv/e0m7hdF15471/zbAgLdJBDMYfirq3zGuYcbBGv1JiLuBjQMgUl5McqD
A64UZLBn8SzXNSpRCIgRDaJu2Rq5Jc5xGK6QvdAeWjPA4e5tSQI3jV2E9dv425PG
mRihkDf4qVYtKbGxl2C1RFwQucDYldvb/2CjPjKF48kDn1pzyaKuSpMAnu40PaM6
9aG5p4ne4ZyZ1NWg/BfUEu/ET6SoeKSI/5qIq3mtBuJzHVOZri8Y0ikqjm/jdMzn
F7fCWUw+LPkA/BiQcu28zI/R8VkR36/DjYJYMXS65NQj+aVTOnTVUB3QyMyGTNrd
Ne4AGi3AoCvwq1WVjAbPkuhqD0DM2s3V0U0N+7VB+BOoi6qcEvAv2bOEMRzkcIvE
Ip1e1uzbivFCp9eBtP97kV6N0vnKeC/UqY9MRk8mFKXCuoHekbNFDomcYeZEMukc
45jD0kf6Vvgb5JWlzSP1qDS6szweKBeWbc3OhZQ2bIRFLWhSZrF4fnwG27+o1hxH
7dW40VUrVoLsYi1uq3W1IydsQxSyF6rPpvBMxb7o3ASf267CwdqMr7Qe0zRyVt+W
CnYQI+UaAhn5TRPu3x0eYKqwfJ/2cXgU1n3YirkMDmYzC52UyN2msQCkV2sotoq9
rsbRIw7QiRmRbXo6E9TApdT+A1lgN4MjqQcWkMgKveM5OwBYWl92esNObexcZifO
bJRO/AwF0x+qcDXSS8w6HBpAANaqHyYfdA68EY5eu2JRdlsvOJ94A67hEmG3F55g
+Igi+8MYP+3Tza0CBpErbW+u2L/Wxqli3imsLPsO//H5UdlxPkgGItvZKhN71MFw
nTjiZxDBJkAbu1I0MaU/8O0S5Ps984C64vEyk3LxqaEJypcIB5RRnED46bPeTYL8
/PMLlq0yRFgYWajU3mhn8/W5WTQHRd8614pFQVFwQvu3vRzmU9hpnhpmAGTc7VBL
X42utUq2sUkZTl3+H8Pl/hWGLK1eswXkFB1n4uDBFBYSibM0vyRMQlWOEGLkKT1g
mcHiV46GKx2biXwZyMrY+I7Nf1hxd5LPlZa8ZLIqyARtYe1ZtpSHg1OECLOCp3AG
9w5LZ1LN1tkov9RxXmM05A==
`pragma protect end_protected
