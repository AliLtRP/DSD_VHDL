// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QDzw0GeEp8EDQPKm0MICAbI350TYw/KU7ou2NBkrc98JTa8OhUkQXzjqXDAo+jF1
ap6NIbst1loY3P1Oyt/1FMHCO5cL3+CRsHcMdPUshw0z80HyThqXRjhq1xhIlOvV
5+EW/lEEGCf3zTTB8wXoptg9dOZSxryQDWIn8Ym88w0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29056)
XylCcMMYvOHhDpL/1LQmNrUcBqEQz48wUqv0o+tjxk2aLo+W3uOuX5PVnFaJ4r+T
Xh96YTvtby9xsr5DuHBcIzS1ew8uZBmoPpmBrK7KrlaDykUt3vUFywiciyQ0J3Kb
mfvSVaOe8Q7fVTWVQAnAm/14qMNBMlF8kghEk0pfqK9YN9DxHNvgpEEqGKD3N22O
vIO9QVN6iQSpSbESCFq7pziKds0BQDWXsf1E18PEnNru//sFeY/4HezLGjRdvgC6
ScGUxmlR8ouW/SybnLJoGIIBB7cylGmEwjAPnbC0Ioia6CprKuL62E35iLvAcndX
bjjOI7UaX5t2EZsrLXjSTw3brxF51XJt5on1UNgVHfnauKuIh+i65Y4JOj90vjTF
JppxupaoCjTPkBC515TMPbT8XuQmW7zIVhrluQA2tZMBFFtN+tF7zFmw5yVGMlYm
90BIV6LZNT7dtqq3/0G9D9KNscrtNSKKCFUN6WElavFMC/Kx7bSf6r+CJqEvaMs5
hnDVlPN1FsuWROq/7sEcD3UOGtk8CS9T2VsXifZPk29gHzz7y2s3LRHRSyJWSxcL
T73115lOWWiDW/0IBBn9iHACe5HZPlc2C7uFpOMqqNJxPmBv9CQub/GrWmiUkulB
1CMh34IzE2+2j114CUoVsrihbO2+XN2qJfsEBtZamRtglYodMLCNcXo+psWeiTt7
aLC4WINklggaAKgupHanlVhcArdmW/py+Q+m/qmWFIjYA1GKR4PmYTcAInI12eBc
B2Bu+7qm5y6FdJZH2GqpTJA+Fr6PJgN0mXXJKJcIF7Q/sWqPVCqZl2h9lpalRIQR
lQhlMxnP+nrX4qCXEZbl5uFT4et0Ke9bnJDkVA3FibO/LEeg3qvFcgY8wNouCJJP
qCaysJog5bMyUrg8jvs+I6JmPvuN3cNaQ8sGKL7h2cw1N5EtmWvT0GPLwVuPj5JK
cdOBLrqeWEWtGLtaqAs4Fh2AqA6f9w+c9IgUIwF8qh6/pT0RO43Ca/05Duamu3Pv
A+DW1dewOhDahgNSofhSE/FhiPZaH8vV/BLL0Xy0gfTMCfbDI5o5WiQIWtOeXZqe
UdMrs9YqKRjNxxtNeM0hDbgkB83G6nLlUOVBlrgZvM5ORlQzqiEenis8Py0FkAjP
ZxVkzpKUp1lNdTAMkG8Lp5AhMDV07lxZXyvPRasidTxxI7saTNXhYiXdv0vh9LHa
w0h+n8ZAXwWS7s8PLy5WW+t557PgJQq4zg5/9e+vyrBGfZn94QYtCv/s+hiCSMqN
JG9X1GU1KmngLmod7EfCKRj+OLIUOV/NBDJC3HSW+bf+WInwj5ZaHjPaKESxYjql
aKVTBXJKDzSwTThux+kdO2BzJj4gN0nett+7VMevZkPcLTDbwTJCdxFmkndqUvLD
NTXtn8W6tuxNEXKBCMP1vAf4VIG/M/QqAC2D4VxYtKc/85w/e45pKwzmKnAqj9eP
GNHbXmlBUdNL2ySOiLc+15oG1tqzhzlj2XC3WaD7coRsD6x6lo0go1kXGBH5uleo
J5Z6QhJk70bHAZTaLoJ1JK5uY5sHNSi/RaeYx0CbyfxaUz12KjAyLtF2UJQx+mxV
6MrWMeh1ii4n0oJdhNEaApdzPezZz1zMifu19P3gVdXlUKqcbCKlDkSU1pXNfOvu
DZBVrCx1l1UnMxX4uBYHGRWtWeL0YBjWPaFngrjFYwCjPPc5fLlC8fvt7kmDwV/r
eyOrsrIBRo5UkA4E8uHHVOcZ+DMqkrZlzDZBDydRq9NYILNpt/bt8ybiKuMGk4BQ
7eG8hcKlKVY14EZvxhiyjI3o50VoouZpgOHBIOc0S/7V0AIWEGvD+RjXCWeumQ1J
+PG0Hv/cBODiPmAhVTol/2uK/dwHISFu4GfBaAbuszYClg3i0CeXhcQ8jc9PgCEG
4nGU3i5Ne76gysAmWupvFwAKZoai/7doaFGCsgZ29iVK0W2fZG532GxxUeZb059q
QbaCZKPBsG2u+EJP9e0deQMns9x5NhEUWnknxKAfUzVvvoJbPDGvjspODV8V1aPN
kUpqUI+EqTCYF1P5fc+5ldo1mPCFz5V7cZPiqlbNUbQHMFWIuWMB2LVXnlQkrZTc
zh0sLhJoU8ArZGD/VByoM8YAmGiWs4HJGIuZ4OsGAlEOtWU7Zruai8ulCmmIs9kA
ayEU1i3DlSbAjuSaruFx0Ez01aUXslaUMpTKES8dCR0qkkJRmoagtUyJfm/QdyvT
HHYzKVwkC9xRpzED4wepOle/Q3qkXgMI5JQ7bowyrSuY9VqYEhgGIWgEVLggTrA9
nqIl+uOtT5QMVLIAv32j03q/Dn6BtBZrYX6cf8Qdi1OO1QbuoqI9u9Cb8jedDWWa
IEhVRVl/tc7e/f1PHXlZ/uE0XxZidTPsmvLeg+RtLRfZNce43vMg4uMjnspNM6XY
RW0P3LcnZDnFlDYGL7x39qDTszLfNFxiV4/tj9Z32qLIl958EbqdrIGvOaJBzPzF
c+WARd3MW9kz3vKS3dlbj1QIJguUT/D6QscR0Ps3oW99R4bssRpqB2n/K7SmoeZE
xjEWpL/1Gs3ZtHSLeaJ93CryqjXyC1njXCmYAuifkDNEnD/B1nCDZzCQ9ROy+ZdJ
ETWdcFpOMa86QWZABiuKF1SK7ctkSyDS0wHIBJeQOx05KJeBNoBx2H/mAXn/Np0C
LFp7DcLVKt/krvAprxbtEznv2gWTiktuDtIq4DVuT+fzxwFGPdWNVVG6ErkuQMRI
A2zvoIy18nTmz07JM60bDNmWiaWToPRT2cPZ39SuabsEzwrxIvdsfuiz+DodOFT2
QEN6qb+ApemRwbpmW6rVUTJQRll9O0wB4lFPcfKXkiFcPIZ65dmsT6ADuDwv4Hxz
1ZNM+mIRjiwNaOppprNvtfmKlztxxGFJTMmiUcI4fCq+p0nUe3Xc8UmO/qT79zfs
gZloRJixYpXDt7wmu4j75MYmOuMoZMxuqufBxLwX5AvTH6mXgEmUWFyl28A3ASu0
x/zWQxYSAVQghI6O6FhSzByVpps9bQ8s4ZBd3PKUb1eAGbgnZW6a1B/zSyHvCTVA
sd+mwT6GctnXLwyJuD9wZ+v7mUEflrA0Ib1DFT/irvm8djVqQz0/mV/3wV28R1M/
XF0l9JDlKefHCrJG3/qMgVJJHLK88U2ICV552hop8+tG7C/tp3yTGRiOqHY4rzTV
JpH9Vjn4V6rI5nbqktxjTkHCGfv+6SkUJMrfT0g99je0jm7yvuWBM+uAWIOS/cqr
7F+WTjNpkVUIr1D03W8E++MUV5OpKfaBXQL/CZwWi6wNnOIP5xGKtd+UsZruGrUp
RgPRtU/ka3lkhbPauPTNV7nNL8MgPqVRKj6GrIipOHTkuQncxgYtl9gzfPxl6Vhu
kn4xGzW/zZ1p4KtLt/LOcxeL45RgRqD9JyPn+j/i07VZbXoIUZ+aHvKqQThXywYB
u4CQDC+GXSqtyMENDmACbBW24Ukca0o2UY/iiB0ytANzaQjCtPutEUw+Fb4e+uGs
LB7+v9ZjbG/f9pPJbEtqnEBjLx9IT2QBpurrS3iDzfdDVbqDZmiu3o7Tw+ZoYWVR
EKmfS/JjNPwZVe7p6du/DzWDK1rMk/cEbte0jfta2yth3ZYuy9H547aRmetHv2Oz
XBGFWtzQyV8U/2JvLHJ1OzYGzKgwK++DBc26DX11JXNaBCf1GXNHy0XpeicLfrvw
Rpvmn+Kh++i6bD3YZCGo8EdTVDcNzCvUdNwm2bvUI/FP8u6eUTncMmy7rlOPJzct
jiLYadZXamNlMnyFQOp1PrXYKDts4ZnJCR3urWg60Xbla+TFuNArNt7CyEQYQH0m
Cb/y5BdtqDMyYpXT4V3sna3Oe7wZD5HRkkSfYnP6mRXVx26xz7cia8WUWhGv46mJ
p9/BKBin5gJlRw/frsq9rF1s3TPB0F9qHIBB7O8SMxKwLpVUxArOPIoI35ims0gl
TQG7wpNd0RDIMECP/cwtAujlPyy0myXm7p6zMrgcZyGqOeVTf19RwV5yQxGA4YC3
7QOz5stwazBWAv89jR4jtrgVEaxz+qW/l3iQNmeJX7kiOmr8AvLPvCrr05k2Vb/x
LpLfK3QdSWY3PgPfx5cMq6KYrfcKsma+IgiPTgNTlpk9tIQdsjJRicxWmfOVN6dv
kzFw5KhrnIJblN4hBa9lB8FcrVA8ffprHUfhqY2QvoBNtaGskYnpOu4+D1xgn3WW
amZcbItfM7dzdvpJPTdmGOJ5/7K4gU0mZUiVeBamuflPTbvM9/7d2W4GBTVw0Hqy
RSOzQw9N3ZBfJl4Tv/cjHRBRquB1oa8MponpB4r9x4ogyAKp+O1NcwEhBf1I3uzr
15IuF5WYPxbfkBkMG91XA+3FUKZXMi/GQqZGC6uyZG9CkqgpzLiFHbZEnlm69DY0
KpSvrbxxZuaSS2nWkOxl/Xe08fGB+EO+TBqtNHV9Xy9uGFk/RZGwjrLopbuwyBI9
AXYSwMhHcqyV55GPoI5cYCFN+JvUMjQymWEL6n7jyWsfZn0CXLE/nA7UetVFOIWZ
Jwqlf1JX1+neUWFeSFlb2afc/8Fa6cd25le1x7ybcePS+dpEyORlbycoSV8+EQuG
IaHc3sk6Kc4/ow6L5kFjm50ajlpbJbX7rTmhXALCJetzZoUofEOCht7V+MB79ehM
ToAcHr9R6WsXSztYO7Eq83Fvxo/XPp78BhAqoiEqXxFav0KSi+IEqRa3XPU7K06N
V8JnMX+LsxXqbZOaMzQTRr7fj3Ai4jGgTZVgoHLMj90AyuT4KHHUN0OBF3IFltWP
3XcWEZKay2ldshQetCiFnKof7rWeLG02BHS7L7pz8oEud+vtyO6Os/YzYqvxc7w2
ONt6De87yM8Pho1TThMz+ZgLT5wvAMIVAHiUHViwTYwOcCZvG78PX/jzmpndwXuf
kZSBp2gOqglgOjxSiaTdiz2ZAoGTkZnW2L/meYCZ32eSKna9FRkbO8dENpTM4xTA
BY3BAJacKPyytKIaA2cnrmk56/j1big/+ln3VIAnDuCWrLwUCRS2tUj3zNU041SX
vq5PlL1YK0yaykZ5F1GcY2tUXSxaa0LcpxlF3HMPAiwG/nBVF0b8j2jz4M7+h1no
6/6KJHGkgxD92k2LAXSi+y3kNvVSzOEXKQrpKIvtzOIlmJ9gukwEVEU7Gv7JungL
yaw4xfN/++Z6BHZRlOYF/L9tU8JGjOUcw9pvJKmvrt9Q50Z55oHcIibZl50qrFnD
ZepQGg5CDU6zwpH0q9szvKlI56U99WEN1I1R7irXbKhRY4TMtdfYD1zLDA+ug5tz
ain9q8dylzz4E09ymt7oSQogvvZovvBKp4+wJCvGt2hg2thyaMCQOs03HA9EvZVx
ILJGQMgcHMKwX/HW9uTDn2uhEUVHLKh+7pGck12TJOBUO8j/VBwJNfj0nW6W3iCl
21lpeCuMICdgC+6T4xTQTRvOYajmHZDu34lqV8qgMXr/fSnPDX4+py2/4CxmRAjy
VzQggPDobDrjvl2t4TRz0PHQHxqL8CxQJoVDdptBOBLNsunO5HByWWiBhyGPCRvf
3jfS0HiGyWeXwYelEcv3+n2ws1VZDpWCsssO0MBhFf7riTFumEht6w6Vzd3kfiVg
7E770t4LjJ8kb1NLYGL3UNNkFwrnvfMc8vF33Kj+LfXvb3virMk29JWIEW5kz/4r
MbaBXZ08lKW3KQUKnNekcuNYRF39BRCFfBOuWALu7y1k+/3kdaOUwsdElJJ86afB
7NrkCovK8m5M2tu/V0w9zxaPDWBg0I5N+A/HAal4wRUybCRUp6KWliAZZ2YtLzKi
QJMbmM27HEAufq7f6tC5+Q/qQYX5JDNfziX9ZQhGNyi7XAhRdnweQMMug8bEci/q
CKxMXnJG2RL8JkxwpqiXDsMJrWzIL0kLbrP4bYPutMu36OrDLw+EySzJpv3qn1Sc
va/ZssCqxihhWZfpiJ+xv8fLiRJctoB7dBkCDnHMBQWh98fhLOzHgrDhs6zCWhkB
u2u/Sy42C6Uuzou/V7Pbie9j5FyswL/WEEJ8/H4BzTaOHRkeNivLKuBl7Eil1y1F
PNrVhShftxE21b2tokSfqwf+u3xuyL1UzabCpSh3yMsjXaS2hxdKrGc9M3ucfq3y
WlekCkteuUuZPWxFmCj8aSv5vIQdQNU0i8p1skMNZry7EZo/aqj5g1BENqVlwBT1
YZDWJzPQWWzWd5uXSrn3lTstDV8qpBo0u7kZMBu28BWwdtQxhf4IJydIifz8tCk4
4UkQ4gd5Tmat/mAF9iwEHlEQPM+r+K/9iTJlYiNdRSfNPGWLL28qWo9H9fVor//w
2Klw/W7MvCMXEUxBj+OFakia/eG2BrxTToj5LGfEhGkL6DFZ82ztE4aNt47b1/YB
VSBz3rGkbqO4KzbxiyBOxAkwt4wvQk8EvnK9Lvvm38j65LZF3SfrxQpDV3PNmIAP
nzqH458ygRjN5J0wnuKhK0h/POSRH8HQR8VUcF7kgE2QZJ2mU9AZRfEu7H6y+fqT
79VO1POh1u5loThETXUl5ZpQi77pQBfMOmoCWt6w//17iWczJy+m7Lyb5dJbTWah
W3jRMv/L15KPK2XtMKwRl2ZyVWoqjTSs89FtrmiY4yZuhdIy6Gn4TeUD/0fKKo6k
odM3yrhtWM3yNL4FwQlTyPpWM4Jz8074M8Ih5T4aY5ckMjAymCoccK8kWBXukZm3
o5NPr2Cctvw09DU4KnRj51Oip8PzXnCGOp+rPepHgFah/R0vGZpoxiZuk5j+/mNR
1ug59pJkrubI6SJzdrc92V65wBRFE1glsCVKUH3Z2Gz19FYc/XpXTXZZR9oNfsfW
KB3Dtu8XX0TF+n///SalT/Ferkgx4TkaxJrBgzV4VTMozScPL5RDbfagUbR0MfgK
lU8RE5eD4QaMh9Wyw5cQSYLNDTAEwAA4XVCW4xLBgmhGAtfrAzeT9bBj6y8SQDH1
r/sG+tlmImJmgwnVzb99frDkCIT4fsQufOA+MI+9ydaeoaME6jCzC/x9+9dGVnQn
fZa5d005307ZwD+epKixP7K67PzRcUBD6TPbBQGOh2vnLmcUdrYFz1t3tIGFasD2
8bw1vd7fpdhXZsJvTYRNl9NoRb8lsJ1MRGsCPlwi4u/7SiXk9HGCBCdnjtaHIOtU
4JBJBdU2D7QOq190ndDtpv02dDnj6eiLqka7gWz9+v8ITU+Rs/HLbwEw9Lr57j+m
qCfOtwzxQwAy8AjiqTMUpMgxqlerI/e3G+9+K6muFX4fAy2LurLQvwI6H/7pNyEr
Te11DQjeUIffk7Lh59lsDYELiV8/MOd0OlEruIV4/7RFWt9nA3sgROLG8j7oXZfV
+9Dd7AAxPsfbiC9EU1cLLtadBcjh5jvknzw12TlSx8buebMkY/uzMrQY2YgaygTI
R2THV7uDucDM5hEAbhnEmtJid+ZvpOrj8hQgl99f16RxNQLKVQkqfa+PEYMq/8oP
MMnrU5AKADh8uqYj2RIknNzA6CmZoDjFZv3CnCCdKDSJmvNXJLDVtdwXpgkBjMwD
pNupsyV21hB5kX0nZN1BDf/F0+ShZVXTGSB8LvalRY0tFpX4006IWKjlscljfVe8
i6sFDmPW3I9A0pu8rVFSIPeCHfczfZjlEmrYtPpSi5HGgSm2oSH7Iuil5xU0Yog7
ZRKWo80rtyXgZaQLwks1tl68ilvNX4jMnd184Gql43osjvpe4GWz4FKKhhSDIHUD
g4OJVOLEtEfnoTRxZ+yY/5weNAB8/Vdv1VGgNW0qtl5namuvpf6ZXcByhAh5uw7E
eYxqHOQeWcFum21I+KfdBJpfQ+xJEcgBImjtuE/uxniAKkYeAAgRwFTv5iZCenMS
i0KZbvKM4YGzUxYUEDpT7S1ZmnM1TIoVYZi6m+Es5Hck26g0cSRMrk37ie1vJ71k
5JrRDsofIhjXMw94BBz1X+v5joIFaOJe25YPKDtfaEbnhS237XaSCOWGckV6EjEW
Nu2p6A8xHVeAyLNC7vLeNvBMsLZ7djm3YgXjIdI00XWvRIu98hCm4AVRpoJ7H66E
8UmSEsmh3X5piqYVbz3GfUULTjxyn0oPCdWAFl2/QdNBlbkBsbD+TfS/+YYzjG4M
E7KSW4ybAPi1Mp5BMfCm30nMW1aVu2K8KorngobYtx8sT7qclLNP3wr64k2ThBjS
utK6ed89/SXUt4zwa9dqCmfz1NKNeEqEk0kOPZmuceL8cRbBgX7eXcRXo+0L4Qp+
WUJc+xeEBuyqpRhFBFSqydUqgyu2p6YRonUDUlPHRJ5VJp1OkG22R+l91BUMQ1G/
qJb3Ojjh8Ys1hotAgqAg3zAH6NXpr9Q07cvhAKim7H4w2fbzkJ03NnIXOG+FEdnW
yw+MIxRCBoW2PpHGgaUNXKKBqQt7M7AzgOfD4W0yt96zuUFxu3D8i6RXl7b/7oGY
rp93BhcSbrb2VIbjbcFjaoQ/gESI9mJLdEwh+LgQBJpTG/9Ie78V5kWPvxImEKwB
2FwLkE9IX/FDtbWARrgEwnuMLbUw45J/nMe7higYafORg2DxZUGaTH0UT7r0oc7j
WFzdZWAHLEAK0avZyV8YE0m1RZNrhRCStrwGajNS7mL/V1WauztP4EkA6glrjtXJ
awDYketelhJzVES+XiXp3gzS5Ymmc6Djy5fOdkKbWbKb92I4lABdoCa3Otm1RlgW
FiNZIbbKzYugjnQJITNYN0N6SgiiUlc+rK+detmOLSv6mJJ1PVpSyyFKIZM0AxfX
1yMmbFVBCBVkzHIkHiYXnRP4Hb/p1cfUQWSO7e1P45RgwRy9G2Q7oc0J+M8Hq4b1
NZFrF+/jdfedUA7cFf3P4RHkYpK5ILi+PSUeAFzdozunv9KJsNleYdaCppTVmuyy
Eq/x8J0ehX0yVlH6OKKKZ20IcHQUCEyKD2EwAyGSutLB5ZhTnsJ3Un967Ktvc05o
R/IbqtiyD+L5piWzUTGOcD0B8yziGSWxjniCNsnPI+g+HdYLnOycqSJ8Sw2c9W06
wR10qCu6zJt65tBwyV9FyJKqhY+G+0BTFkELjIijEm1NAUIZ73qGeEhxl1DI61E2
xDTadXT578U94ypSIapy/QYqaeeXvTxo8vBty/B4VUcMVcMefhYUI3mm8nvcqQZ7
bp/BIX0rlw+SwpIqHJWyogg4gROeGlyyozin1kFeE+OcNZ0xGHWULHEBRgQULRNz
VOfwe/7zeGbRAhyvxhAM9/8eMSzI81j5Ug8PnKbsrMw9Tjzz9FqG74qUnyIxZSEG
rDKjmlpAjsH/y740IgEWYWa3XvHKwHxpj8rpYHb3QOvMbwm+Lc7JW6HQ4axFsEKb
F5fhWP5+2ktoiKIaa/tEEYAtEfHPAawIrlu64z7bgu1tU4h1zwcsYma1S7GewnWL
2gA54sgS6zKX7ZYUttbx+hgYnACJNaoUJwyPMUmL2pMp4ZrR3kzezuNqdIflgICH
KdZr7I6XzD4btpY/LwLBgI5JpB7Psum1+c1cY6sx2KzMPz9nxOd49Z+/8Q3pOm8A
boy8ArDv9e8VCFcBkJkjMctqPZHt74OmUCMwRfPKpk/D9YulS9oCgj2ejxm46/Uy
XuNgI+YOFBddnvpoDvne38/fkncKloQZZGKQUiTpQBmioxqPq5nTvkilUguARLyM
URwV0XEEMmrJCFZmo1aYVCPaI1SXgc9ruVGU4lvvqc9s37qRqGVCHOvaOYW7bJFL
l5BQNtcRGfccPpybm7ZvwS0TEbj8/18wKVxEBvyWbqa3alyLc2CBzrzY2ZNrUm1l
neuYESj9n9PryYC9E/+xcKC+koNJg+S1nxZBSQXcgsbwRkyYh9e0fXY+qYH1LijJ
W5liMQxI3gll9SrMm0iR/rbaRYE1bvFuedF7k1E50ZQ3pZ8hQ2/Q+ghUzmJB0kqn
/hgQCz/m3dSkrnkU5T4ZokHiWhyDp+GruSXSlDRumlF35GmUzz8ulxECn3oELUne
XKwPcaAn5jr0qpYzFiWVjWuvjdzlM/XvvrtTQQ5Mm9MxGrBwccldEfbpy0Hb1uCb
+sT1HIivL06qLKqJFDM+oMNgfo9KONNCgNOZRyYADgnzx6fH3VfhwPgQpJ1xe7nU
XR400CtuzGaKRd5jIgEzaHiLyncg5q65jobK5KO017zi3EwSI9/R952zm6lZuaHH
RQwFr946DXUY9xbqQs5OHQVC13ouG3tXQOMMrl6+nmYC0kiQNvbvry+8KKo4N1V1
c4D7B7zWWwo2r8YN4uZ02KCqsvLlr98t5ASX73/sphLP+ySbueA2pT+HnejgumoV
Du8bMGrH5KJtAIn9+Wj4WWlrvGuSuAjhqC+RWThgpYNdwndmUKaxL8IOZSJhMIlB
9jKlXBkAC8qEKy/Yz7IyTKaWdU61rgqjRKC0YRVe0jVERRQnoeSENEz5r4ElVX73
OmA4buCWTKN6cXnQyLEkvYsydj3tnvAUX8V0PZ/GamxBFH+XS/JdEbsjkkE28D5z
/LDFXa8NbwM1jw7trmJxkDGHd2e1VWpnUuOW4ZViG7cpgDUVF4l8oKu5FMuc5a8P
M28rY4dpWxoQB2d83nEexXTXms149zdR3yNDVtP7qr4qdqinfMIP4jsSRBlUL+Vw
PAep3NHD+EcwutQalnalbvx1Oeafk9qHFHx/a8X7eic00K5YjoIxdstf5VSVGKiH
in96SSu4/tPlgH8SAT+E7W15wdoPPpIySJlQOz6q4K3IRJtdGTKkZxa2EYpsWm/U
m2kazFLiIjQ73l1y7nlYzsd32LPsS1WZHQndLOA3fR0kHOoKn/+Yk2VLNmb9sTKm
jDY8bWPhsGAInDGW9CwE1U+vnBhFfaCCw7LSuCw2TtmpnkYtl/Sdsya9WjU3oYDZ
8HpVVPYyyhScyQX6qyasq6DzR2MrpgYcjmdY7ZupgUivzaqTjOhWhP9CJtJGGcjj
XmthbWYkxoWIlImCynL01Zzcbz8LM8rB/Lj8pBOAZ910eOmbWt7ucg6uAq1N7owd
YMEvjfnzohP/dPzbVgvnodNI+EgzJy6TeHgz/w3yOFaqEFCmt/iC8GW9iFgZz6ez
UnEKvXNjlad3Nhr+69tcjVavtN9jSjjomz5dopXde/35sBxBGy1hP1X9EG5HLXla
O+oZbtTy8Buoafi2FM60GbOl9rEVpZivz/fKng2aQF5g5RnQjx18x403hcfzG8tp
CcfF7BXfgf+n4bGnicjx/0vaOff1Ohe0adYxbQ5O+Zp3bV6LVYIoP/SfgjXpvnhw
sE1JI9UQwaFgG4Kdt+iLohLIB4wNAoBajDoD882w5GzqRnDuDqvyUZosEDmxsx5v
TiM6/WpUPIl17N3dPmj7PrOSmoRHv/kx76HcmIPZUk73dQOinHKuHLJf27VLR+Gc
wydBCJCIfDwf/o1UcKnu8c4tFPRw9Tyvas2ZY1mQBnHnJx2GMhyHOVFK71U6vu7M
tIa6QZWbQltJGF5PjKzW4Y3G/aXRKnnvg/ttRmXboJKTC1oMbx2I1CdKvjwz2wum
2bC1cwpTMeaN1vDw+dqKriH6+97zqY6IHRS7wgvueaclXtaLqLi8cpob/3BEoQjK
c6cwDVkB7iA0VP0xfv7kqekrbjedYtMxitqcsMbalV9ASEm03lqRyNeLEuVGaVRC
s0GJ0thK4gYLXBYbFZ5ETNev/uKEx2/xMksLiS+ZphMUrUOuqfCiqwj3jpOTWueG
hqfkuf4kxmAcbI3htLASwYOQJLavEnAyttlduKyEJKiY0DbbaMYQi4lHdsZJTBzE
GXkS5XwUttMmwpzgDmCvXKgThvVxW3oy/Rwq0j4GDPNE0Bel9lPMMjt2nxBkOLyX
GZdtOkE0GLMuS3LL43gvMq3JyBTGpvcduTJfBeJ6fD0B6ly+WivaM1QIHnutjj0n
D7BGRTipN76mEkDc/OCOtkmc3PPmJG4IMnvtK9Ra3Y+x8bAneiedcDY1LcbCIyxg
NH5XDm/122VwGkOucH0P8LGDydH4eeTaoQs2+3HhI1M8gCE528zhw7XuaNQ68/VM
HsLWbhdgeueyBxbIngX8JvariyoPEVJCBg5ce107WHEpEIbwQ2/+CgV7dir/KJzl
OWAY0jimxqmkpeCx29M8mMIKV+YM8jIF93g/9JRADUQ0GKce32E13zyaZbdlIVtl
DsmPO6vvZTRFS3kQ+W2aN+ODVoYYE+5BnN9Ebqhi8a163f3gEkR/GjbIKuB7HNX4
DQzYS2FLvAHCJVe3vblsSxnicqkXpiMcr2C4WoKOq0R2xpXZ4wQmWZHKDwe6YUPU
SVJHfxasWsUyfDI2IcvpowYUzMsSoda35wzL1OpTxkax5M24Ro5cN35nc0znvZZ+
g2nSNsBD98vq39T+eSdsMlwz4mNq1SfYzo83d02JLODhupGiSAlWV5gXVcwVNDrX
kkiXwxe0OCJPRP5MmQbGb/KhAt3cq50282nIkelVDoTZ9xjMz+cFTZ7c787TIUg7
A5yKn7NPeVbcVG2yFlH5ybEhHGqLSORLPA9gR9oV+0IHPr7u9N1uLSi7X5fsjJwo
kWxmtdiFY2pMoy1in8iW/HywMo7E2wdpC4oLLjl8W8sTIuGnQ6zi/FMIdbcTSK1Z
f+OJjR6giw2Mji9Z5FUN7bPZdH3dtnsMc6t3bCuyiKxoQaBwnW8YKdvGUZy54bWR
RAQAj+/XkpSDGgDMd9dSz7Axyo0AVGQtygCUAiTJ+oMOF+eo9emyuYd0aXASiat6
3ip/bF/l8ljDR3nhhQ4OhZjGOFpYB3liHbcrvqLlXeWNmNPawV86CtnS9woE2HC4
XgydhKEOfVQaoHmOr/KSwCh7mUwIK5/2FNyeuafqDQsIPd1f4pTSbvXNinVFJE3h
Gh33TfuLnvKVNZrmij2iIkssJs9OxdCdJv+lrKc0atCoG9Pzl+qSCBb/bAW2vLcO
Pt1cY10tFK+wKkPPLxQInxvztOOgE2okNvtxtaaLMRYm3f145MCX1FCm/5O0ZSM9
BOvMlzyuN8CK140T6y4JiaQH2038fpXn95UCelqZ7jWSI/ML7iSPsZXH58JsBOJi
GOC4A4mt/lcK7azecBE0C3XaE8DkvWEQmC5QwFWY+jGm5sU0OYfZFRu76mB+0BWN
1CfVCH7LGNJ5xpwtX6xNoqc41EkbKKIqxTDaQodzIhEn1FGHeJ05Na1LsO9vjBJJ
7McRc/ZdX9R4uxyTYWoRArVwsDk4SHeKu9HT+J4Z0U4k1X8tPBW8ozI+R0b/5rh1
YGCpKR14CFbKaUl+uZ1+Hs4YEvJ95peE5PaBzNG0ym21HLbK1ZiMwq+ThSTp61eR
SLQM60tSmrRL9s3wMxRiCwKw24RbqYlVMoklqNpMW8G7N7jsEvNTAcTXcc6k5r7O
yV3YW020Cmq/yewV86jwY44G1FZVlgHKa34NUL7pM/99QcyzEPqIMmjmStkclU8S
UB7RUxfMAHn69LpWHRrjl7SFxGaOx7KFF0DSf+tRDiCVfLa+54o1jdin2E6ft5n7
3hHa3Sm+DGjwj+vOBsO/vbqh9T5d14O/qixg3GS8zpTzODGOuNnmSaCK7Pg3ONlO
iYpfCvdL0uq4VLKoSLelqWjPbtMVLozzVsJms+Kf+n/jafOkTSigApWAiYnjBGD3
Ykab8FtCsOTY4Omo9s/ptCwyyypAcM80KmWEPEL4LehIgFRXg33dSjfFrfXu32Jy
V+zpJ9rJ2SvaBfL9gtS3bCnjb5YgFT5hdNCxPrCvQxFtnGQAjUMxd5oqrk+tX0sd
ZMBPW0+WFKb6s24628kv3IC0zrlmNK8EPRgELMFhNN3G/AXqfkZa2aRdnT9Jlt7r
JbAMLXXmamY5wWrJc5Ylr20Vl31JAPxwYpD/7gZKVdckLIrm7DF3B9Ye3ejXrmcO
v1dqoO5up8cc1LhYjcgZxfpA52rMtcEqfk+ZQ3kdJrnFYeKaETFiIL2LpvCB0t9F
dWoIFLlw1tcqNAiFr6kAkTunLaZBdM/FnXLUHtbdjzMtIr+bqzsOvL0EcG/N2YxW
pth5GzEqdNMz8uDD4P3B3aqiEWkTEijWAvQFmz4yUidekTBy2Sx6J+6JZqc3961m
BAEI7N5a5E4Obslhmw3fG3yzylSsG7uDWbzTRCYD0BTWbQ/M0tRtn9jIZ+bWh5T0
u5m8JIo5/c3ivHpLnDuF0zvMZtF4Hm7wz60kNwxpFlRarM9l5Dhtx8/pg2DbdUVj
rtnDKbIwaKY5kP3AwfLmrXXrbTq8lqm5Dl23tkX+LnuzaVq1wg14LMRkVrwVal5q
NPgMpXMZyuo7GojueUJXGW34w9O9MevUno3wMKteh5QJ2EI2Q1TjgvWqW30fet4E
ZDIpfAizcuxf8E6fdSt3SJJHUCoDNkB2lHWJTXOcKXlf5BZvLPw197R4HnWJWSIN
lHGryAalMrsUdZipMUMwWQxpkr/oDCNERS9LUfId4TuWd6jzF72abKOT30ltMcWo
uzSQmPwxdheP4iUVcwftTYBlRP36KbblbtwzevrX8/rsGRKov+GqyvM/xibepgwN
KAiwcSVfibiMxqCYAprSMidD6cbrLBSDwgTYnsyvG0UH84EzpUlmC7aUwnBj6f3s
O76x+WC3dtwwdkuaMkWTw24MHhaH4gECKc8/srzbF9Lmel1fGD2FQs9VxUwksfAT
kzWpsjRpdrr6BdYQa4B/gyPG1y45l1o7H30rg5pdwNUaJlgYInj2tLV9DJBxuoqE
5i9DefkZ6p+9gAWfkXAziClbDfJytzBBVnFa0mIm9eJNv93wyuJWIFlDT+pPij8k
Jvey3HtfrVABEUvvREr5JMZKYF/yRQ3QqnFWwgAZYyZ6Kq22nllKlERuc8qu80zE
5/5haE1WNrGhNhI4iDLw1nKYKvVzJypbj3YCDKDE/6521x0ukLTwi0IiY5cxQBCW
7da0gQ3B4TCTSB3n7il1MQ6wzHYE2eckwEdBPLJoF1cvmuAJ9/PocUHiIm5tGRJs
2BbsQM9Tj2/otLIU2OSdbu8J0HPRjCaYWlwnI297lxIFtX54ArHv4a6Cg9MTeCyz
6OEzpoYaoGY7BzK2O1ycr1asuPfmRITUO+0Jla54hor8LbAXT6Wl86czPUJfpVhM
+tpmrWYwdzf1BUeai0+blX8NsAMCL+gDZnsZuDHaOV5AwKZxL+B9+n2c6cSvaBzI
ji09KUnfohS671rBDAkT+uSnc5Q1fg1lwZ74MLTarEC+dCW6jGVebn32mfWfc2SG
9tuEdfeAv9DIfe3nV2BEdKo+Dozv5cPOQcGDvYiHE+2qofv2f3JKM0Se6XssEr/n
KCCyW9hz3QvCDg7sGuXdtg8JafX6GCsQdItGrPZiLe1S3KF7KjmxN5XtZYLrafpO
PXBUSw8Wg9cp03stQYA6QwG2VgJSeSZnhYmoDSy9qYiUzZo7ERfyrr6/1fRJT8md
NOVUEztL3VNEFrMCORm0JEvfXWf5uCIpWj0RWSsGJ1551qBR0WLX5eWa2fJROqaP
kLni1QJSX0zDDNbVndDMX5ee0ujTTuAJivBkc73ODT+7BzSQUBHwxfgfTBfxbLRE
HpbBsb9SdsA39Do8n48nr97vIesoMUur/62ZChudbjDTnjp1Ub/k1Bvqrci7N+Vo
9lU5+gt/iovPANzsEX8G2gFD5SLdpLs2n5FGCEIYBK+DK3H55fLXF9DUbYV+8121
Ol0fp9s8n7FH/4iI06UwZM+ln/DdpMFYpOmf+4CLsD3lTNp9tuZbA8w9FLcadVIq
ePH8sKKS8RZyMbg1yr15iBJStmiru2XIKRkDi/Cda18FlmvgAaX4yDWomAefVBd3
rWLWPjrKYkqhpe7e/yslSYg9KPEVua10fYD5q7h/szbve4RvrFTq1JfdMVKbkuW0
Lzcg0Ws0aCINinfTAToplKBT1eygLsK0rYVpo4EN6z72f4RZ+jW3q3kVYrklflqd
x4stLOnRrvW9SQj51nUaz0FDKRDfby6Zw2JfWEcao9RyRlI6wpdSxj731LUbWpY/
5ta3hnHarBrfl3IbwKmH3jJbHX7rHKLYE3n5q0pABcy36MX8vobi7hN4e0tqdAkK
nxHi+2yKoswQyFLQ7zMzkCdb0NzpD1hdvMFuxPuTUhlpJHTKP0tC59QfqKu8KEeW
Scw/PbDIXe47IZG1u3w9hD0ivAl/t9NqM5CsEUgMOKMR5fT6EJa7nJ+ZpTwbYYv9
9D3xqOMbwKX6sPM3pQV31ffSVqL0R7Ucurnx5020gapLHy7qZSRNEYkYT5wYd8Lk
0neyDoerqzY3kDRVa9yE+87eh6P4uuAF/WrRsubSdbRscuhuzMUUSLVOPUM9KkKI
0WgMRemgvo7QD3XrI4/Kc8h8CRETESucL5YfCx4aQcPcexH15YDBu34qIKvuCy55
1eBN5ftvJ9FvP9NMCLk5Q18wg6JH+8IUD/5hr5HjM0gYNDtLj/0AjPx7bybcEkgE
WtWkJv3PqjWhQsdV8SOjdEdnNdvyk66blJTUJqXDBeWWgmg69QRtJ7DpbdnJ9ABg
Bam196wE5PSbeMyl+QATsssu7oylxnvoi2Eng4oOLGD4JK8a1Xjlbx1iPUFe4dCv
uRV2BYmCq+hKlN8lBE/OHE0A1XZUZP5Ywo+ksqVYBnTRAq/10GA1r/hgi7TK3RvR
Wse7hdv/ZB7V3sKqVfBb/ZThAudjc9WtU0c6C4sL+ZqvxFfVbS+K91GEWdqlHnIw
Yb9IonsTlhow1JnQGbP2/MqrlDJvlShy3JLPTxGrwE3758hwDli/BrNdI5ZTP1j0
6Nj7CkyyvxM45vy++DDUPrjPVLt1IL5ncFS0mGtnMYvy5JuIIfSBVsnpYZXD5vBV
WFJsEdDFnV+ZUG7bXtbQ7CKU/kHaOQmYlYuXrNeiF2g45uwLxtcurWVDGqZ38S9j
M+9jCHQ9Vl+ZswwjyN74Jbh701mIDJQd+Mj110/Bh7GZL3gNRwlosQtZZiZ7AEYX
kzzQ/2B6XzDOguGe8Y9arm/nWzGqB3wKlJ2OKz51LjHtwqUAtrYDo8LMO5MaRNyA
eg8HUQPmw9q8hOmJzWVApt6w1xP1C8r2SOd6h5UG5c16HUYl3xQUCIr7ABbe5uzt
emy/f/vNBhCnM/CfreAjkaWgi33rkrLcbmzsUZDHLMvIORfDoQyoJ+B7sTQoF1SX
LOLdaUc9LG3lLs57r+Yz42UduSCZbj0cBKX8rpnzwetF1/3jTN9Oz0enj61nqJjX
6+vkZdOmE3pFZtqzPpR/DGFcHXMU2oEeoI8/Zc5eTPi3gNyIQBRnPcTAUb0I9YQH
NxlVB1p34XjSWDlByh7jXdK9WJ9toK98Y9iOGCFuvAMvrJSoVmOL785vMR6+6MUn
CNR/AYAbTW6eB8Uht50eeWfowA20DrRa4A9tBQo8zLzLqUNwJzxrhw662iRRKqKf
sG/WDxzAUKOgqWM3m9APKnJVK7wNhjv2LmahBLLmI0NOgwFOQC4hGrq6HbzGcgva
RN28Ze8fgTd83lsGWMg/BCiOCAKh0pyJxC7Dy5qvF1oUINPxIllqTpLJ7f0a0mOU
gGDes5+vR6f2Fg07ryt4u3z08ojCYebn3q7uCpqcJnu0PH8n2+F9B9po8diZm8P6
ukU8cvHpNEImBva3lw8nKeCUH/OciUXZ1O2m6a27zew7I3vv05yP8MJGqUcp55uH
tPm/dIaIXcybsHH5qompFxjgHYc3WeUq2HDtzXarj+5dHrGyiU2AiJN5JTR3+O4G
II7qgDx1sl+aQe3qWSPeCID5dAvHH7e7b5j1STRqqu09wQF5cQMKtFSKX/1EgUl9
N37NK0OXygEZQqc/p/psH38hrdyx3n38gYN0t1vHqPNvX6P1WYpvrHI2Da5lOzWh
gUQe2pxngPgkXa23c9THNlWig6kL6AHs3wtr22/9DdrF+pKNE52F5yGY2HZT4PSV
R8q6Qa5HuBFffsdRJImgNeA3n4IWmvnAjbX77HAKjgU6N/lU6C5Xs/fahcaElbAH
yAYp62VXrkqCI1CxTxQGSP6Xw/9c10ubViHo6foai2H+QuWBzInbfRY1x1go4y2/
edGKnu5XItH/ZSuJ4Rjd3hpf6YomtC+kX3QMzfOAghsQiY6yzTOeYDywqbjG7hIe
dVWyzjJjU+3tPCjoh7vA+5m3yJNAznZwzNpECOCS12k07y5gIOKA/aouIFNxxyH9
Bp2ztYT+zyBNLjSuC8GVHN2byfhNPAf+FV3vVPA9a/TMP30DXmWxIVa6nsku0O1y
zqGM0acszSzFTdr/j7vEAIABpaPuDNcpGGbL6UoFL+TsC4Pkr2LiFMDkzDfmNprl
Wh+9Oi+GxdUP9y0MJE2rmDHXA2J2LLLUA8sHCqeZPxmhGRxwWhPyadYeLU91b5PQ
mD+FIC37+Ix4gxrVdSVnHxfqNDaGKqP2RWxsiTj087rDx4TMHolt8fuPUAVSU7/O
8zpLuioEca6MuBp9Or1aT8qHm/RLIQcN0OMw2G2sAxRWHqDLpiXSjgyDdXnHMvfu
gDPnuzu95A2QuKxN4mLp13QeyAVceQPIlqvYNitkSGFl+vw3QmODkrAaywFJK1oX
XUrdZxCWcOQ0kbSenaVL7O2ZAZq97yX9axSdmfrdeyu3gDD3cCL6vSPcXMHL52g3
DuwFgvXE9BftN4bePf4EOpAJESo0pLODEyocmj08zcGmeMtQ5+BX+QY5bvkYWpIV
8xw36sRaFfThH0Akz5SqzE2ESerCSxvTM2n//bMewzkj5VENp7rt83B+dMZXuHWn
gKoKQCXgrlLMl2PHSM9AJqFGgUmwnIsUNnBmPvfNl7RsZmAv8R5cwQox//cqb+vQ
TEWm0nsevX0oaZkgNycD6owC2p4xrrJbLp53U50Yo5bq0jeF8xTbkoWeiejuGcv5
EbhqdaznT2pnBmAJ6bVW5jHd0htncPiy1zF2puFJ9mPrpU5ItaRnodi4U1zRN1K9
Ca3dZSEELlwN4jIPxnOPZaUDx3H8U91Vc39LfgjGHaLL6WZQlJMkFMlPlWhkbqgi
Ie7Kj1d1Swq75YxFm6Nq4w1rV73fXTttRMs381AJBXgJ2s46IXmAnQcr49DDhJ6J
R+zy2bQmyoOe3vEV/DvrflxuZG+/5PjWpaFDfthjhHXq4/mfcW0RF1UXQJz3t0Jd
zKcS7N9xsuyApElJ+hIpLy3Xx3gUzNg3YhXt8HHxwzOzITXaXEx1hiRbHMO5MFqv
0oUBJ3Rm2lEVLSbNiuf9xM6oF6Rmwug/MWMIqn+SwYVq1fygwlvJqZM3egzJRTcV
3Fq/YHb5iCT0eU2kWFemI6yfksgGSULqT+SbNJWj7uajlRhVhUg+gY7dbtHMIQnC
EyO+5GWkVI5zyYLiHNDn2isMIp0/EHGfnv519yzssDJGJwR4Ru7HnV7qUHykttnS
VOOc1Lx9aoeX6diXhkiSjEJsf2UK0pEgkmbcMq2ZXqvB48rdEBqSChQN/sFrPEhp
IDrIf6sCMj2qB/KRsXIKbw+GlILCLJ37As/ZTYvsXTIR8kQEV2WidpT0oyHqHzmU
XEI7PasY6ZKDDTX9KBJ4+9+5IaU9fMls2cG+ibXbdr4fKdw+GYqmM6630xvYpyn8
p6RLKbNIY9nmuNSIlW59mTsOhzPyIOEtZw7wnA0iC15sUd5cattTK/Lozm672jak
2FBCLM1HVgzjYNzI3wEcGQiQeijyYNQ/6IPvScXagaC621ORum2d7LyA2Qx7QrV+
GWmER6WEWr6/BtajOJ2VgKfyua18InvARgrJLq0ZTn+K60RnVw4gOJ4NLwByAGli
M+Spp1P/3N4wNzqkLaY9YDQ0V96FTVLrYKfWmyO0MsntBvh3p5i2Inj95iy8ozMO
CYcfS6BvSinXs0WtuHujjxsJWUJaY1y/B40AVt7QhAOg/pDlt5K33rSgt86AM0dV
4dK3xRuNARcJy2KGNG/c3TlQqvO6WlrfFLFi8ERS9CtpR+yrWHck+btNcvfxFdC2
639QfCRcnfeQPGC9J5TK4h+dK0T6PO3+5UK/SnY+U8NDQkc2ggdZDQ8dwTFo5NeQ
Ipv+Ye/0zutse+qOwiCaOEaHko7iLXraP9S1DqOD3AoBvE3BOl9iaHEpMC3qyMyE
gadxEhoan+kpW9TOkE4TORZAyHV88ffgjggyfsZNefpD4woNhi2Ic0AxG0QK7Rmc
tnaY2KdT3w7tBiXYysu7OxnleeJOjgnIancIC9kqPLBdRkHPGPh8ewOs1nyG5vlB
rOVelC48f6Bg8DXz6oBVaaPA3zEfvqxIqPJiH0Jw8G7EeTTKsOpjQ6Z3SGP7KFRZ
6OxVAT736QAkPt9wi/b/HqgO/jzWhJObGLn9nofddMZ9s4E6lanZfiTCtqaur9oO
OHHHdPVbKmwMnzrOIbkizPbz/ptaGTMB8EWk573WDweD4AMS31pnjxoxT9nztuoz
Kdd6Ho1yNfHqKlbBmmCTcgxnqL+zzG1tcfHamk3no2tcvqFnpbb0t75AD41RvXw6
TJUJECkWrJsxHaNSZRqnrrtA8usudJO7CIzl2oMdpcZnYjP9xQbrC/CqlcborxAF
O/PsgKFV+HQM6VQS6N1zZtr/oODxUi7S5LJwZDatNY69dqXbuWB5pdJL326HvxpY
ufIpZEMZaERnfQCTD42IZYhLK0QLJ/+UAVCASWo85QDrmVMU+ylogWoHdNRoHg6t
aJbJOhnKn1cEk8g+LBZjx1qkGmf4UPMIu3cqyxOF5iAnJsE5QFG4KIo6l1SqL6kA
a3toQZwQ4tD4fsL7tbOh3FH6d6YFqYlaTn0YmmssMM1/zYXo7oX90QJN8uhQW6PJ
nGK4KiC9d6Mty/ZEHtyJp2hf9KxRSNlofrsHJOhuMDEF7lWdhaMY4/mpNIPjwI1c
mtggV2PjfHrtdw3/Ych4tYDzg0Jn7f+99PqHVRPJ/LtdjYEWaky14uF3hcSXb1uf
psM5LZBJxnRL3rwQErAX8+t8gRajRPjumtfQ1PaLj7vEkd/PE2j5aIEHypRXhkWH
NiJwT2ql6UnpwLrTGgRoAib7bEn1qU3wQAgzENxbiHxc4O2hqFujMg5sIkut1zHD
haFKurgougYgpyAh8DJs4Pj62QQkZ1ilrMAR1MhyQ2GAOuC4p1rIX8Yq0FcPca1V
Cw1jK2mhbrYOKrvaQU85o+XlBC0bpA/RjcaQlefX7eESU5UsFXRNVhE5iid5iBux
jjYKoAdqmA+kG8MuGh8JWuj6+qQ30zt6lry7osNGnL4Ad6GvMLMm7SUjfTERGMDQ
4tqvFqx7WZNfoZucWXXfj0MLMgPidtiwTUtwpCQkL9DW41A0TnFcygwfa4yoj5N1
WWWjEIBTnbktdKRvylmwOmiJdJ/Y38sfnA4Bc3Oic1pVApkogCCYJxu4ZnYXRKRo
btAQVW0d7abtegYuOzjdEDLIvf2kjfphDSlHxzlw0zVdJx/xOEa+TIzZWdx163V8
sqA9C/RN4j3CsoRdNsnjplEety7UePw7GAWetoqtER8tJAJ0xMtiL8tNkqAkwQWC
nDvCtleCHbJX4FkEL7DDdl1ajZYMf5rCXHFGvVPpyME6lJzsgwKPpWmktHP/qGMQ
d48xnhHvgTDrrSjTUu7BBc6Ipx/u0KPQ4EFJkZqC7nPAMEwmF6eGONkhRXeSezXD
stKWARSlTuMzVVDUKdwnIwWd8wNnoYwojoDh9D1U3YcASQP0qVw/D0wF1NYwvHYN
SF4d/QpKBks4gKnzqiSPfU7gVMuj7xHiQlrBWBH8gElHD6ESd/9WM6kbEoEswg3C
Qe9UumxQJkmdnOyRcEcCPHQM9Q1cudfEdv35VL2NNN/ThrEKRiJbZ5/5Sxs+U0/L
YDw2yPLF5iyZd2gJREwUR3jYSwyNNIBBpPxzRyFd0vHgX2M15wDT9vW+MYa4dfFf
dHh+NBzs4oYhjz42guqT3Ihgf+Vj65v7ufCE+z1CGTsLqio9QpxjqpPpennAG3iN
KDP1iml/cUePMS3cin+avnSYX0+KW0jxQw+d/ik5v2+fgnNaq0aGI2J5SNN4e6Pl
gKAe0JhWTRN1QbXmJcuMbgmjoxIotHyPpHGUiVcw2ks7JaxbcW/7g0q3hZXJDiX/
3oc4dYxGXAP7VsepVkvhGgkDskMD7+SC20nzUjGmuE8Yt4Vu6M6L+WIwtzYrz4u2
dM0Ddc7tnJ1O5xaUiWLO0FFBT1ptP7KqLi1GOH9sNPP1HtvGzzIGElIUDviYY36y
DZ3iCR0HNWClsY1kz19CyRCFA2O4dFkVjeZPoLy1SDsVl5cl3CPflL5DCKx4QI3X
C3sZNVzOMRC8UfDcCasj1AH2C6jP4Sqnivt/FvFtKfxCDvj0jIhg5nJhaKv9RUE+
xK3FSX2/UfsIaHvPVBpJfd36UQiR60eZqUIm1mYciPs6PZRP9+g4Ozf9V16U/dqx
p13vDzT/JiD61SktVhqQIM8+xVbOuxhZgoQQVj8QwJFlT7lwnVvaEjSl3ilBrhPI
/cjbSaa3jprjUJKaarkpNioq/kVVpIE+4t5sHHwa+WLpNNQ6UJDBBAmxXh/2e13K
M1xpb8UUQ4Ya3HzqMwbm3W9nPvHvxrQyMCllYf7twpIIitvKhkH7AAQW3bRNr51Y
BhrTwK0A+tHCk1LYpNMqFsH9dIJLZy7Sxe4ca8++QU2DCewW44oaW0ysW4WHZoL1
6LQ5WbS3M2jqDGW+4A0ZjF5MXWwDIqXNg6jPbGUuj5y9tfo1L9WSVSVK9wYrmESw
xCrW2iVV6QstJoKZHRXIhVMpk0PCk5On8lchVL9Hh/x04a8ne/SXAN9e+TowO+D0
ShN48WyKZOD9OpvHnjZKMW6OEUXQ2xDIu1rRwSiCBBsnzudnIcUV16/T3E28g+kv
yvfaENQbcT2p1yG8ePoa+kW1VPjvYNFXr9LV7Y16kSaMkQxLLSsKm09MWZS0zjaC
gAGbRXCPNVkHVYia8zkUoGgit0RWq8MkFbbUhXIGqWGKF5t4os4CNqR5WZx/e7nD
KWM/58IfnRZMm1tC0qQPZRZnA/YHe0uh2W1MPPcmbwmGuqOd06vge0vfKfehMYNO
h/PsAucsxSZXUy9HlQLzz3+60DqXemm7LuwALXN4++DvBUfUaGgyVLy71oflsgpz
tFsp/QBF0+1xWFOh1DW+nd2N4etOTjqkzS2xil6ls6e8etP4lI+qi/i4ClZCI5Wg
XvZTDiMJHhWHdUQKkew5C3tRwo/eGUo6DlYWw5Oo+NP9qr/s1I9PWl1o96azm7A/
Bp0gcNEa+90G54YoJk5IjqvIvzukLcg0BoQkLKsvod/RdeZzD4GAtAnw2///hJjH
Yde0eQ/ovjA2uxdQb1Wmvg5FwuPLdUlcTh9zBCSUebam3mM3sAwRuOGbT0uqFoNx
ZiOKYlONE4Ee4u5JZvrkhFNpAx8Z7+1xRQlKIHk2fIzaaFHYVMwktBqzfTZ4M3OH
AXV5pkL+pyI7Ay80Ma2AAns5N649uUy1p7q/6UKSssaNbhV6sqYLnM8TOS3R3vIe
UzQRxf6rBEgGWiLSj+Ibjs2SvYSYPL7jxWBfH6eTH/w9gnVZn8DIyfOZx4bNeWmz
l2Q4x6hK8QI5ZZSFO2mrn20POnmsINBzWWhGeiombjEGY3QPiSHhpIWOOjg6Qq2p
EfPVOHManFJLmOjt2LTqWvSMfUPt0tiNAWqOP92/GygxS7J6QTO6KZXqhR+Oh99s
NvyBW56A9wRjzr9LM9tz71dgnt88E1bFP+OwyJLoGeft0AxTnkAKUJ1DYTuhZfRI
IykA+aKrVqO00Mz1htyceDhMkcrKxSX0g7dn3owIDSEgP8coH2Bx6rZqGXpr0ysA
oa5/56gRVikdSvuwWiKlxLb0yagjjoe0jDHxobwt2T4580ZR4i72TlAbiVQPdlB7
LnbuvuZEYOfWtTazKgrA6ORKwyxwv30cDRNZ0UKjCwvOwUMRv+SRtCCgA4xKmYc6
fI9q+xWkJEB+6+I7rMcQgsu1Y3rvl9wUeeY6UG7eEAqhk+WJrGDgP9MCUJd4Djmt
eiBwptKYy9yBFWlpewz27CFd/KkavFtDiE7VDn0JxFBle1TC1E7cwfK0MzR0ov+F
e9SqlgCeved1YAUmxApm4Z3QFnCJOvp6UmEWMpxQV0V4mZFH8IKFQyiBT6Z6LI2h
e0Ln+8uCYUnJ5GH8WZO5q0FQLaU6yR5xZHA4opukGUGapAURHhnKl757r/5ZEnBb
gQV1Q6NWbtUr19z4qFs2hqE5sgF/eZBo94by5ki1i1fsDaZTcqIoFvoZSQfaRyg1
nn+BzIazD+M7BRlKy0cQK7OmCUePIHo37Qt1By+ng4egqnu/F22j5NE/vaM9Yl6u
DrGhzHPlciOL/KBqhcb75KqR3+QGBQNVSrM4Vt9ajT6i9LzP24qPYRcLll/qyiRs
YdSAaZWGGmbG52BYmXDaJz8rSpRZu6GaL9mfmOOQ9tDGwCjGBBu5uIKc/eb6ZYdU
QYA4r3qto6rhdHa8siz19c8tLl91N3wSUXSgARDnhKddiypIoqvRq9uJTIUQjYkr
G0YfaRqxgfmHfK23n2g0bNtEJsP7nWbo1R2/mPoFc3osFeBYLtMwEUT1ej2Xc5Wl
+pOoBqmaxrfcZObaIbXV++wpqIdRShDKdXy9pP678i2Fbi8KlMXYWbi0pV7VEC7O
R3gCjF4Qej6CVrODvh7PQDbO8Z5/e7JzXQjo0r4fnkGPizai/sYmL66fAaQcMUTn
BE9L90VsPzNCUoDSBizQjpxcmbNTnzTcbwAzJsekwaOFHQEZ9FyXKgMWaqegq6QH
OJ7Kr120L1/Hfnds11reouktV8eXKSSKqyvaJor2Nnl3SXmWXaBjtnNsViheZMQD
uL/eFSv8RkPoJ+czXkgzVNyjhtVW6oXXXLOeJxxaH1j/CuokkArHQmgOaWqF1Efj
8PHQnmW49dxDUNcxrknqDOtnffRHrrhEDsS1E0NI3v/0uExzaAeLX4cLZEyQS6qy
1opaoVKK0BBc4OgY3LuAUALhF8jV+GE+aCqV63XHHcDIGkulMa+Frep5B3cZe78d
Qz4jrZcsQ0UAxjnKt5j7r/RaMaWhIM7ovMRbEkKTZbnm8ilJsigmY1tCDnP9LD63
tPvu1+3mGq9EMyHBsK38PwGA0xFHFHDf2p9ddaJkO32ORT09zzKigVNwlbSSevcY
07It/uXkhuwA7kdGUYpbmeVjsgWfbRCrYTMlVMe25iln1BaSmMn/FKI9DRKKL3q7
LUgaSxavB3AvTDeJR/lFbGHmBKk10vmcgr59uyXnCptjUY2eiuEboQbLbwrBu3TJ
wlY2rlgLFtZBMksij+83NR2wvfRE0bS/nNZ1zWp/mKnzU/Coh4ovfUp1jo65k8y9
bZGh0VgZc2M+vEOX4jC6ssnjy87X7DD5sD6NwKRTG+nNteadkjOMevktbM7K6UJY
43Fl6psYPY0OMqtirrrX0y//ibnSxOqzim2VAiQr9PwDCENjw5j5AEgLDZanYSi7
G6PfpezUWaZqais+nQO6T1hIadybjXmxtzyTacuXJPCC2tknH2cCxpTriHJbaxVQ
azWWTycBZIlYdQyLY0TcQBHfwMr58vQVSFYiptgld920hk/BUQKyOqbcWVHaQul0
TgrGEXDETQngs1rKGDfk2Qla9lgMCv58d/c5dC/jMyAUCItwafDp55aeqq/D65b3
DV42YyhtzRyhAGN5Y4G19PndMw21d84rqfT+saMcaXCL94wuNL15sFUAObv8lbil
Rss67taqO3L5WebWlA2UTbExjYZRpSAd97X8EPCbSJXV+5jITszjNWaodbB4j0jg
bmDGtGHK1Ur4Jqo0GfeIyNiO50dUUR+DiGW+8rV5AXH2C601ubJ32CxQvJzs5SsO
Nvru/1IohXiEligOQAWLvTiD8Nxccf3hexngfvs+saSU0IhJcL+frsNduc8Hox2h
LsEBeb0PYQqtmElQfFsm7kq6EfDclVsWS/TtycLqkUanA1Ha0rtrfmCkFrqCn7l+
cYUgKxGhf4s7u9+ARijNZf1tWJFaw8ma0RkfOwNj9Chx8FGoBdoQfJTM5qo+s5Sn
RzU+zxISS6r+CVuhnF2QmnA9ZpmKttlx8aUdMKVhTjlZosiDq/8kotXnSgx7fdCE
f9N4+1zV4PCM2ezdDvXk8aq/0g+LYOyvj0I42IDaXEajNbN/d4lERVBhWUUZzGh9
uvLefdEC60q8y/jjMRaSRc++oJ7Wv7ctSZptHHAXU2m4NBYW+X9/peUW8OBno2n9
lGLHdjuXozxVfgrmo2eG9MuilyoMSZ9VZphqXu5oVvVmeHhaUkCkllYv9XLpPW2P
hCwfrZ79jnjSoj7Gws4SNf6KsShu9SvoY2lOzeNToY7fG5a0SWAgUyWXJfBcjbf5
Yx7AnnUejlsWsemD4qlaq597ReIlFZtEbHL9lLO89NSSJQuT/l5G/blfQLJCO4IC
wWMbT1TEptq1sk8gHaC9DPyEbdcTLlvZKxRUADYx9o3nkgbi3zTTKsG4SHkCfhA8
gRmt9oTeBQ6ZRPddWSaYN5HU32bcMLaHbztphJLNzO8iv0orPB5hgGvKHoT7yRFA
HvfoocogD1/uebcle58mCde4N8SDltNuh3jy56z26FTALX1bYhAkqldEOMUrYaLy
utNOtvhwO1nUtKPe0uoMlcr2iu+4p4yiXPZBNoJWh9v3B8hamwXrRN7oQf1Tdbib
rIU7DMBAjaChgwNAAn/JNQUfg9J8YZTTh3okItPaIzVv2eFQYJc2n59U6JfD0kMQ
pQYJMCQIUGrdf4I/4T8pv0qILWnQ6n5r1gqYA10PHUapi0rsEM5BHXnBGDojXz7j
rmxInJ8dS+ZtenouoVTdQvfzQv456WfrdkT3fiYH3e0D0Qo+qMV0cCLvhH0cZwvQ
FueNwqaOJa5wvqWvrMDj0U6Al7jU/vgON0zce//F5Uj7T2ZhtSOWa0C1UvVm+JTp
MU6YQ8qESkmQxqm4Z8cEAAg9swbnSgyaCf8h/wtVxxjPYnawWeA3lpYyBxF/+hjV
UAzMVUsvnR7ACagH+LX2fygpp2hNVh3RZx4Y5wPdZEahVJGUmrckqPoArq8evD+5
avTEL4BbBQn+DohVMTUL+R2QjghLKz2Cj9/sdGNnNPf6oKgzTCg/QqL8gjDo9E41
Wb3yRYTzMcvZh89m58jyarBNX6860wjngkJgsQItou3xgZTnCJysCM5wATwvQ53c
RehbNn//4PM1ga109maVGJDbxlut8m1XBmqlDopbhUXT3j+j6o4ODD6bXB0KgS5L
Bckat8setKX+X2gZncHKTy5aFYy5wj0pWOKJU3vLfJhjR4tmaEp0ya+jQqRWqebj
V3RycAGhyox7feamDYLhZKBEyceO78uyC+b4tBdGn1HBoBxtMyArn28ebJtrri2s
r4fvRUM3FJLRI4xbYqLXFwl6KRMMFznqLfal4xSXqXVlKtouEE7+Tkrk4U8vVIf8
KMHnYkyNseEat1ENEU/dsWUiViOIiIV34ezHJm6oIyM+mK8nbhW0/Y7SFEZ2f+2j
lL3dNPaUZgkohHXYfHB2JqhuwKbK/w9ajWdKNVsljcXLBJ9cCQCPiADyCw14Co88
nZyXaNYcatdNYxv2CC+85VkjngozKtxBgdnc7k3mUypHkDzi8F0hmyAyRpAtkpw9
p4OQMBJ9Yu/cWKUITc6QkrDJHYJ9EwEWriEY8ljQ5OtP7CTi1sOcMT2lcI5emuH4
6P1wWBDc3NLDjwi9174fH67KN8E00w3k6/cQga8S37qudGUjMrXy0W/R9pmkAWRF
eI01S+RskUUtwCq3Th1C8/Gqw0oqb/I3+etUb6CYCxY9Txz19U5mNSO2SFzYloxn
cTzP7L1P9C2sLGEQE4gLPea56X5EfOm1dTmkpsvXTuo+icPGkdU0RKe0TkZJZSgZ
kzYd56c8jQapl0T9ATr2K6HWKRBH7/f0VAjXS5bCiDiO9qhrtcUzPWxmEekKfky9
m+/f2vGySSOm/PfYMdoqPMybXRtoHO+WVvaFwf4RGipq1nEIN3zaU3lGKuyXTdZi
DJXa1OG6kT5BLC3MwS/gbeaUDV6i+R4fOGU10qsFzR0+r0vCIsgj4P+vQsptQwfM
6i1lSmN2KvbMPYWr05BEcEU3idhwcqLQ3YlfLIH9RuZYCeKfykjYm1p/4SF9GWJ7
5LLnwZjY1nMJsiJfZ/V/0H88mzsrq28ueOwuBjkFgHggGyPauYIcHGJUD9nEei62
eFQg1zgLfOC3gkGydj1H3L5HnGsvIWuTTwtg0cpV3vCPwwUUmS9+Zbu8JULAGo41
yyuiwc6c6XXRHrG8kV7qAElBbOwBcq8VSjKk8u+Rv9IEVcpPFvTc85TU/AGKjYm7
BSrXs4tBJLq4DKP+qYgrLzRfvEZ6N/9RwMln3uOjRDfdK8E+uKU7uouEglnpIL8s
ginCgzTp0mM59vKhuP3+EP+Mzn8y2xdpcs84OLhHjF2vznk2zrqE1ILEyiEPJsPJ
QgAn0p3Ir6iTYNSrC51u5OLsckDA1YYepPCOSdJMVXT/Bedi6NdmzY+0DtMNU+5s
5S3WZEqEJEJkJMagwa52NcB/8YKhFmHSPweGEdlBV/csHaJyX1BmVyqTyst4KBWD
B2zjQnGg14y+l+ypnptnBp+7H8VIMu5TA/Yd4gNa3nanhtQf0zPVLvl35qcgf1KG
Ultr6Vpk/digsEI1i8KQLAz5Qa8lnvQVYo/TY8xqWkDHHYNKxLFIeiN7vLwwYY8v
EGmFsbGtMDWzZDaMsjAlGnIPMVANAGgO2gK8Ouyab3fQkoPvyxQrp3X4Fynoaou+
jGbTmK1HSL1M0Q1T8z9HqJ1uFbqjLvHfH9PT5iBaFo0cfGcqPy33zu+88tSw2wiw
pmlHRi0yUUw4L2lMUaiyJmQucjidVIIzZlLNgyHh36q9jZ3p/6yE9GeMWkIUrNHk
LI+MjmUZjhcSVXeL4wV3RKDYSXt0Gs1Cti8emeXbuj2w5reRM9o1qd7n0uzSMnp5
dT6tVXVF63Smfak0CVBnzmsuNyLNAkBiEO+sfPu6fTlvQfWe5fjNUfsPMTGuEYI0
0N8pW1yPu7hCJrnkZUqDs2RRW2gd66xiUMLa698iqqgBzoqTjPSUMIMYLb2DCcCZ
qeKUNm0NKuahIFkzX2X7Egj5FDRfRR0SxQFROHCZ8xuMZCcYuiG1ovHQdw+FX+Ga
EhtiGDQkIuGvIz2YNDB+sKLAyw0bZIfdm/ND5GEGS75wz6x/FswubUM1CJTUGfRp
OzAP379FZYC0c9XzH7aahh1tnSTHRSL1v1fPOhFxJww7v68CpEHQY/+VFOJbx8VP
soF8XQgcieyfKkogdRiR078McteUBj1gjLsl22JuywbsZradBFV5gD9aMO16wpea
U9GUeDH6RhHM5fnxwU/KoFv/zppb8Y0Z0SyfWsFRgTQLhUcVgo25pEB5h5kWu/IC
3VxBCi6gtloe9PHLHq1R2JR9paFNBJlCpWE6JmqICgluEIIFTn5yN9yXcnDofPl7
QevkO9YKNSs+2kPc7weUzMEY52CW0zVpIElMxgUokVf2nx3/JBzL33ZFgyA9oa2z
YDv+qTLOwXag+In+kFUtFYXilSva0xNRFYTMhvNP2c/DiNoMfjiPf1jPumhxQ6Gb
PEbKv4H3sPlJ5gMaErQYubqXBfZ0HBGiXWmVGuRXUPEpJXo7CCGNXl6dGewuFf0R
RvBw+a5pnJICgXTslHXWEvJegy0id+o0EOIURjZV0j4R1wCM7kA68YTdZlCUd1VL
MZRgCkOf0hw3sdOAOn8npzHpmoA9yi5Axu2qKniLosKgs1f+1Zu9M7iiem3rg0fZ
VO3ALTadfzlgixlHHuXA7aSaxr9tvL8lmwew1RdjbzdsyYlAAk4eABZO7VX4tKvm
3FrWrjPiLrsSa8JItAehanMDob2HsOS2wAMWe7JmRJtldwKSO/zwBz9xm+D7lm/V
l2PWtn+MtTOHsxILyrMri44mRbmj1onHuDubfoVHuWPyuXatiqeMhUQbtZz55Kdg
wm4nBZc+EhWnVvj2iu10QTneFjR74ejVl2PKz41H0xY76vRRwybMWxoHVXv76BAG
RT8IReXxrHF77iUZNLIaNIXfH0yAGY2iBz/a9yEIHVxQ5vSoW3lkdquEUym3us4m
xJqAVduluV7LirfA3WYLPYZWIrlpODPTdYM7wEoT0q3AX+8RUXtm9Cd+Gtj+Q5qT
fcfIik32kwR/87GAf2+5WejADmOep8Ogb7oCDxITPtKqdCpXZQZe7e9sgmyg1q/m
ZYuSv3YH/32VUDUo2r/YwMUukgmA2UnUkiwLu5lbIEXciwc069kpFNUzAldeQFfq
AfQPLVnSkxs2XUauRAVcs+yBUwov79TWNb78ewR6GQ/h81aM9yweEp4P51a3Zf5T
P7DK0ebFoQMq8/Ll/nlHUF40kF9aCQJw5KuHxgHAaKQPVHQPCvX3Bo/gwSnNBSTk
/q8bcHtUD0tE6O/U0zn/AFDEdGBAcBg4PGuqicdbRJRiu+VLp69rolYa/2N8eQ0B
UJxmhTrSQzkv6nDJxxtLfF/Ht/b4eizJQNbSKYe1I/NGOyTlk23UiZslTpZtP9aN
0455cL1LKwUcwZAH0IPYsmLzSSUP6hN26Ktp4jgeKI8HLZlzou3zU3Ev1l100SE2
auj+uDarxX4JaBYWfTodJhpxD+GwHE3a7jrL+3KV791AFyMr5HvTFlXKjlOAe8QI
wD6r22Q+0sp4XgXzyICvlWE0E8RnJUOazfRIGSKcnPglRHvE1m5ZRTs3ksASiI8O
sR7Ni1VvYqOTVqZrmSmnjHAixCrCKr1LRImKTmQZpi7u6GcpZx9A9HLmNMk3uMF3
yn9exnynD2vDLoWd+RoCNe5X/fFoCeFkCppGM+MAd5dq4sFSUndcPQSYhNWMcY1Z
lQCf5as88itxFhQFrYJP5lJKlHK/EWVZ2+QluQvFC4sKeIs1zUH3BZtGsXKpW+zR
4iu/Haq3h6RatKpIvR4+b8csZueFUUyMwRa8plld0PSIkozqmyATXGhKCyd6ELkK
ZgtWr7os7OTcVDBgVMplUmTOSvTPf5bpm4WDL3JRU0hlv26k2nvCNbCo2IoySQ8W
jfQm1GmNfRXGET2n4WDOkI9WwS0N+ofsuALkK10mXqV5PDfbMN+kR9nGULGb78gw
ZLqdrrcO8plcInbK1NNuk1uvO8gh9xEO4cEeDxfgMu8JtNfKhChePrfkTe4v4L3K
/iMJWGdBtQofi1gxKRzQR97v+eTOBql6uaXXuHuyWUmdQ2bzXCJ3FZCstLhqUj0g
PuzxZXW8SB2yPTT0/PltQ3qQBA8zunz7sCTcHD/z8/xmtgDsCRlztCA/e5zgl5GD
e+sGqGDxi4fuI3V9jVhqwXqHktTf0RDNAyXDQhzclB7X/2GkWwIS6fjWUltHNeWA
212BpT+hAq/iYvoDBnZCRTpUyQyTGRLOydZPaDuK4AJGU7WpfFzoQsMy4qOTWIPW
feEeFWiu7fkHNbtuDK19FCZeNhfLmXS3ZSyCx2CdZbSVdyrnlM9VwpKK5fpNed1y
AoLLpawc6HGcSqAi30IF8MQEyQVjGvAkOQepeuo+YqAicDRI4r82qaIVordLP+As
mPp+mDHzq7BJNfaiTx89l3py/JCFXPEjxhN9ZkaWMfnSL6Zs+wIHG0JbsA6MZsYY
4EwpAfIjPQKFmvn8h8PVwfAgefS9+uHpx91yD0nYc05O86VK9UUpfAUUuTJ3aKQu
2YmPKyZUaZnP2HSIo94YkL+SWM4pfPlPjD4YextkRdjEKlR6BYhRdO8lAEXXig03
ZLDhb4YRsz8kgXcd3C8Aeb1QOtKXIXSMIIvB5u7/YJxJvkwQpA8NzwHYlG9lUSeq
OM086B99pYy2H2zK0057SmEklUeTXyJUj7/YPDFyc9TO72TVoBXhaNDLwZzFihbZ
rAHqeQJjPNnKoq1QvmBnolk+wWRVO3vrpxVLhbmjRsSexw0GBBG9wqAj5cufrF43
Zvg8Ax2yXM47VE0Hsl6E99i2eSWZCyJuOK/SomP+BNI73dGDozr4rpgdlyILFZj2
c1+Rt+tOhQ67wepvXJEaCNnY85Cuu7EgL0e30+esO5Rj6oauEHubG3FlYOe5hogx
3p4ZTQhR+aTz1I3dx9kfLIOqX5um28mqPRqd4+e0ShOlm7j6QC7hW65jGXbY9evy
nT2zNOKpVf2FyJJDeuPmJAnaUOHLLxx/STyA1hNWZzN3MqHZnuubApAAHBhkrioD
ajq7r1v9rgHi5QQsQupj05RfccA3ku28lwfzvDgrxNDUw0N993F5N6BseK+Ix5fD
V8fJGyMervKa2mGHehNK98qTX+IcQRT/v2dxY6pXBnm6633qMW/1QTeV41hrZLFA
4uog3gX0BD2IA57a3TadJb63si2jGRG/Jd7ELT12XRfEU5VJcfDxq6rvL42QKMxv
ovsy9NVBo159LAed2veck9p8UnPGV/Kt5cBC/N1nWV3Nm0gygNGNtXl3HkhVHveR
2uPG0dDun8T9nGwvI2FM1i86561ko+Tx2ta6NB2M8cQ0S6QsmDTgN2mUhqnphrWH
d+YhdDbFk1rbCDVzr+XMsoK0DxYBDKKQhDC68254Ox3ZRDrDP3mgfu+fECoQ05e8
fIK+8pcu59w4EZgMVOKr7zXpjy7ekD5qRbe9h717GjbxoyMywTpOa0Asadn/gTVY
tuS9aCLQgZJIsF1SbdrKiNhWziQ74+vWUPqVYFOugFpzr9Bp6byR6UGFvfQsWRJP
NfetlKkQ3I3GrjGaZfXAL7Vuvno5NPfVUOdAUGWlVuerrC86IZr9OM/o1/DE3orA
I1trZFS5mQjJsnjXN0htVELrvRZFWn4C8TcIAXZzWsTpzeGnjsqB+RY0mVSr02sk
wRw9eOXMUtt/uqQAOfMzNN0JfrXosBjtMHzFBP1Tjev4Rzt6+fgX9ije9Xy1/GpC
Xv/8CnO68Uzna6IotdjXgmVZQ8R2U4vxKMBeg9QvBMgBRWx0qjfGvnFuGJlw7kqr
DGYYyp8JdsRh66eBn+6MOBLxqsLNdyROWQBYsJMpBhgf/Yf/Qtq4U/QaTYRyWEFw
oRWonxwYsiIswnUmQvb9rH0wYlyBVYDWwK1f9sI8g8Yzrv4PrQpOKE8u0z1kcq82
uapPCVnurR/hwE0iIlH3pIZ+8uwJunpTjRBbCnjD5Wwjvsokr7c3cxBJWsTR1Fvy
ekHhnX3Q0ndSA/8lhQumWUKo7QC0m9zOeq71HUv822I9tbhzeFXXi3yeH/45od4h
lFofIUjWTZJQ5k4Iwh/GLrNKZLk2s3mt43AfOG/oHGxUReiuW2ABi+OcYZMvTkWV
se2xA+8BU2+XutZePzBCMmldnn+a9DNMFbenFl/VWHTcMeuJ78kfEkowW3kbYBng
ZfJ7Syqy4MZyOo0JiEQz+daMx+IQqMRle12nnThbtfTnvg4dv3EIzspdGtNLmR2+
KwbfqrPZRFc+pp3LRj/KwemHsGZJbaoPJJRedWRuU0z2sV7KpWQWJk/Ln+h0zUOH
CzOOZxr6pr72j3A4UwTTLhgQu05FLbtR7ppUSCpXiMJloT2C2ldnmPvl/0MDhvBz
SwZOfPR5I0A8gN8939lqksfffALxQEfRZP1DXueH1mfZEDS1lamFk8XAoBJahtQ/
SnXzh2KdQr7gQwobyVsq0hXpMvIzvk77M7+JaYE39pNT86iKWUqf9RxLVLhf9WkK
wUDKPzy7CFGeBOMZ/mi+PQjiB9XmSlyhbeZ1A3rZ295MmfyAE7ABiYMVbCeT4oRR
j+DpKN2lzfPF0P13KdBzNNkJ9/XdQGdp/Zo38OGqgBhyVQYIXSPf0dkH+FfCoHbF
Hs5K8EylF6sDhNAs12J/lpE0rB4UQpuTNncqoOYsK1yYFckRndR5EcwvBc6SVq7w
7DdIU0Mj9gesoKkYiXW4Dpevv7erdl301cOgErf66e+nvcLiUDJUSRwckUVWoiKv
BNow7a8nxm0k+JpsUTEc2Lxn4Ea0u7WMcSOKpxCtxHTNJ7Zeez23gfQyYk+ii0MX
hSO0gwFSrxusutSEmPub0QCg4aA3g9WiiWhRdpQgaS/bRP+ERNV3I2sO9yo9YUBZ
4uC9P3dalOZvo2mdsSBHOOTY7I72FKc9KU3vbPf9KbEMda+1e0zAqoPh0SrPBLHp
SvRZgKasGAJViLoHuvSlPIkSC8G2VpL2lhnugLTrWxgK2EdDhz2ptiQ2UgGPADR6
FictX4OGi0Db/rgr4dn9IslSAXaLNglWr5dD5tE2dmiejZ8XuwwGfkt5MX4LN9xW
7UKfWl2OZcjlYHgM+hpNLYkfM0ZPeSusESeCmQ2EqTIH5v+Gmmtt+URaXymMDLvW
eKyXngbMmVEB1LeikXG7q/D4jtObyZb9i06nRaPUmByl7bAvk7kptQbg/IULpH9F
Bk39W+4h6/p3QnWUB8bcAXjXAUjWpa/5H6qsTpBLaXmTBuyPf/6hvcs2olTlvWxw
SLJqsNKPdQuYDwy6mnz/2mZEMVN/2/fO1hI0/2OvE/fRWUYkjlcnP6xAtpPbXc2T
H0X7dAmjjUjQkdm58cmrC92TcZQnoWE6G5yasj4pfkLvgBsu7jLduvjOOh8o8Ddh
98zfPN3XoXsruxCF6fynZR+gPkmE/rxEadpoACh1yJqd8RqSNkz3qbOlgn7rIo9P
Fi8pqHmKtgaVOV0kvtQv1F5zGLyZK+aEPXOQSuHOfG7/GMhDt3erTWsPCg0v6BXp
69eXGc4wYfiQ5x3/38ZYkZvMq+XS8oeAIoANzWHC8d2b3InrGRFXNRqADE5b6u0K
VHG1/By33o0jTH6aQ10/CaHWijRbUJ26Ks3jQHl+JYaIlA8CrCpieY4cvJKrexY6
jVcHO3cJRCQmCzCVxdhiVUN/9E0sYI3U1WnRjwJ38DysaUwtwc0ewAdq56da5UW/
pJFhWwfI6rG6Yn41MXUWLHdQKuOUZKttQ8gUzGvUSNji6bvBfmRlchfdiixGUU4H
WJNXGdz47QAqLRele7A7UJUAUdwUKcjzo7ZidiR5w83aOq7U89cGLr//MeHYnJNf
MRrvBTZGWbh2Ozg/CYBcR2LjDLew0OsVDwWD4kGcaCiKnnD9UQQ0R3ZuD5iF79Uw
8VV3yNER6sQbOf0gEnHfae25v1pGpJdNOb6KsBuy3jccVAThaCZBA2dRG1Uwo0XA
gxJy+gBnmAE4QicW+aDGoSmHiNo7bbj7/V8P1txQd+Lzi+xSi7rSSkA6aPlQoBBv
fyPjBfim6VpSQ5Zo1JPZxJHSYnhoEevAezPxV/vNA0Kp1sbSx5KSdGdxCPhTKELp
p/1/oyWf2RZG2rH4ibtxPFgT5/gM5EbG2uMreUfrTUpBCG8gEJNZ0piBk7MGyYWr
ALiXSBN3Mjpw3bnE7HxRS0ASsN9BorQFOHxqbh0/C/zeato+Md4nH3k1viSfGs+/
5Ln6ml/iNnEyZsN1pPxNdomyYf2wym6wg5+IsoIjLdJt1+l2aBq+SFYbblw5Y7Ht
Tiy0JMwgTsb0i0LrfLHynqh6SJbXzH66hLyC5Ok+KTKzWcQYOlztqnfEe+lcxOty
hrm+2p1KoeWBHrXgdzolV4I6ZaRFznN+FTbV/74vs0cPpOSP3K5NzHqqxcJXz8EP
ynEMVEGELrGavHs6vzU/RVgKdUyICVBu7RtUM6olmItT5GS6YeJ3DTzoBVYbFknV
1T4zAAmbMY6qCiqINLZuL7XwIK+VIBqZOG/1Fpq4hcgLlfbQM/ANpcEGENwR4M4t
mIeR7GZuoXdeVapjxBIEXbuofQ+SOrp7azhcXhHOBlXwch4H2XpauJim0NuI3HDw
TLUZHWFgWAfQ7jQbFR7J1P8t2U3k9orKVUgbOkXC1J/5csey/1PsKJtN+LTDBkcj
HiHeHN++0pzVflWbslilwtPkm8eFwkz0EXdFby/NRElR64iz21IzpjobxV0QBMhH
NtVPyknAspHBY6tFVwKTnYDdND4d1FwFfjYAHyU7lrjHnqhNlA+XuJb08Y37r7Sp
zOosekQFXNE9NPf5k3SSVcZSmtkHvVkBD7hcF0R9V/SU+Sh/My6U0cyECTKvWkFo
k5QnH5DGqoSGJ5Q+sV0l2lJCKgfJE2pGXQmJO2ArJwVapExpDVENsmCJgw03aYnx
8QbVmizkM9EFN3kTHBNjCO6Ad63G4voVag6RKsxaNWzKT/lS3kNB9b0vcAyFu7yv
RJQVvp0ZIS5vjfvhevr76xxrCbP0x7WGGLGIXStE/OrRA6SEtZuT4loFprxU/KcO
RXbORKsnliEtLiy+tA5bSAd33DavNHiQUvkUFc1qGd6w649E1nSwl5OR26Y6j5sN
nE8oEknQ99wyAT0Mb2nT6zZKxLuGTnl6sdq+UMqWY3mymDo5yOLUtqVsZ0A4PBXz
OoxI+6Lh1ThdMQEWLtDeaXBtSIh6hamF3HuzKVESsBAGzR2Rhjz0cPeq+s6Q/anQ
tVlbh6w5RZ1e9iRHZlS37WTBP+W43bu7wTB6rkjWBSyHUv5ZuZZa5LIj0NjReor4
vCd1yJmStpMJrLR1Tb0X1sNfhHszaBdDN1WfPahABLTKUwGdIGioesdgSv7biUiU
idYUZhDky/F5Wf6oqDlWov7Pq863h+qSra/WXn7iGMBZMHhInU5FXOjOtGwVQApN
EhNSzpII8FJwT34jFUda/rfu1tZwl/H3Dp925jc0LelB4JlWhMvC0cwoihC3bXj9
RjWWXHEp+GGJMRC53GpMyKrI/W8vzGn5bjLE2JRwQ0Qu/E/kV3QuLXZmFybg3mF/
KKiU4DWdsRqYmdjUe2zLP5CErOR9hTBpa3OvS6GRhgqvm39/8DQ864lMCXo08+Bz
Pp12qExQfXxf3CAkESDqArSIfu8bI9i5iwPrvmIC3M4YqXGHFCtF0S0WTNNxaVGP
aIFLVV5GGWMr5YWVoPcZivJxZWLCtgj0D7AQF2rswFHIamMArCHkr4aPa50CqSlO
/3OrQ8T93/TLEqNDWw0VbrAwacg8ZwPR4N2zskJwBsm4y5wpQgMzkaG5RokkhESh
FEZeEQkAUXRazkmcM1OIx+MfnMJwi9iSifQrVvRA9sdjdVQrMH+zd+IOvNFEd7/N
qBI5qO6VYPAuvZxRPGi9cHMIwV0oXqMiHOsedFH/9AsW1B1pHisC6jWzq8qNKUFM
pqBszEH6+NHW+z264gVmDeRVBHTtwXJdJTOrjcMvk54OxhQotoNhRRWXmKl4shjM
Au0TdRqYr3D2xBN6kEjVFIJkXTXfBoRZ+IuU/RIkmFNG+sXwnoYAlNEB6ifC66Gc
0rIlCgBjU3Ns8UuM9X4blYHyM3GgbOS4jzGO6+G9ItbOy8CNTNpV0CuOf68aBDPf
WymXk2PeF5qcxTpiGZgOtxSrTBuQU1ze5BtiTb/m1ulqcsOJuJQ6C6F72MmO5qLY
N+sOmBGV2xfC+TwIHgGuNWdHCBuvWt+OWBvssFczG0VJ92RwNuKT7NqlZ6HuPQwu
Ltg8nCQeZOSjatg5wLgZa7QOx7H0F3RunrHAn1rWP0VJMmYlisZEPKQEv7xNN3Th
cB87+50d/i5CU9Wb6GpIFRXgtXqU+vC9xlN19QQM/qUbuFHnkk0zZUnvoH7Y6v+U
kblAqiM1zi9RD0tDEb9WZhguwdp3gH2qSgW+3fWc/m76jrD0sIb/CXXJrNhgKNih
MCysKRWJc6eJCfxUQclf+7KDb143//mjJubifoU4zRJuurUNz6qFMCnUyXgUT55n
26FE1OvhayD8VykzHxcj3wEmUzVfRc3NvtfxbMATsOColNxN7EDn8WU3VSxcYYTt
384GfRZukIEIysAQaDk21/j4sA1PrjjfuOTXQEteQnZF3oWtQY8Cvmca6uHD1H1I
YlltaTfbo+UKu7MprQSQAgZ63Aum39FqujlLhtFc7OZj6RS7cIxcpFNtDKOsrvDf
W24fvYBPOcMIzBbv0EN+xlBJ6XZkQksKrz37uHYBla+8j2CHLnIOIPUYG2OCEf/5
rD4+Jx7Zyen+TqYrGIrFkqe2zcD0gjfw4jyANn1+ZL/CWY1xSJUlraCTOPeIPYwZ
sz03Ov7L1S1GNgxQATOvqnVt7/IuUkOalOfNnkCX7DO395HE+oVzANh+fmdRE27f
D+6pDV9iKYJ9t/1nz1Dn34pmmQ9mFt4r6Xwjfr6lDd66OpI9ZOwov3lDU6bDhWn5
8YZ6jXBxJqJcGRiWqTHBmh4UQ6hIDSodygw4hU75z2yF51MsL2dEB2r/VC9A7/AU
VA3MV1LczbwQo57Q5Yfdl5oHsTL7c4Zl+1n+XYX64vTk3CX86a0uAfKkjgwrWzFW
rc6lrSNB2vMc1Dcpr5qyxD5cagYERfy8G3Op2kTypUgP+mzUVTUs/+CmYF/XzA+C
pVoY0vHbGuKRbENQKePaGjKz9y5HTxHB5UqR0kCEZQfH7tgwxwJ2K8GwSZLCwOUm
f6ogdCdSxuR1yNrfBQt0rE+8MfeyuuBkMjeQ/cUXHPldxIFfSAbToBT7gxdFcOUK
dJbH2FC5uFFPUmQuwXa3lfCzVr2KXSIYA08A1Pz9pGfMbPA6O3bLTIYWTTdw6o8x
ExVP1lpvyItznhEuNQ1vWtWS+n7xCP7MRtmZzALVZ/PbYK0ZwOBcC0W64cKecbKC
1j5eCMP52RGn1YKYe4kZIf78Vo5UN/Gpn1jAchrSg/A7DaroLFfho4DOy+OFeqyb
2iZeSBCBmQI0sUBNpeXnGw==
`pragma protect end_protected
