// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
IymIG70IXzpgBYkCvlQwg7UL7PwF6BJbvNc1hnB3IHErGw2hnR+AchKLjqDgys/9XNMkn3/VsdGL
JQ9pn30/kBS2imaQ3YtnfNPyp55dV4RuvdXftKUA1VHIWiiK1TBq31JeYADD5qewn6qa2JJn0a62
1MIfFhhNJ56eI2308Xv6JswgG/WrZ+jyAt5s0UZKPnLrtv2DQQZV+Q/XSnBZZ8Qu/REe/kvXxcLp
+kFPmYGgGjfNFbWGIV34S4VJQceSi7D2XU+FQa4RHZf10gjQNJT1mUnGXFLJaB0BPqXhUPP4qf/y
mcNNvCuHapZhpHVxEaKhHw5+COv6Pr9XcKmeHw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
n12eqefYdIrBUkWcozktKxp0q5Lq+bkxMv2GIFd9O9MP2FqM2GvEtL8kxHSmqQmeyXAXElWdGLKA
AgvcVFmbV//GM6vJ0S0QYU6a1RsuSIARMRg87jhmpXnINuPmZzddMzub8/tG1YRpwh2NQKlbSdk1
DBdu0NO49x1fot+WQNpo8UZkKUrusl92PaegUnHi8i/6vK8aBJLMk0aHZDUWCUydFm6CASp7PL2g
ea1HLydopjcfe5TbXMvlnxPMf44iLJBCq5p6Ypeg6GMaAQMcS3BsT6Ymekcf4NBNLGl4MpsY+uLE
wwsBR50s291XGHekVeYWbBcpf+mWwkfEYD51v8ei79rNvtGWK07JKQQ32z2rLEiygZ1CDFpBkH8F
qtMwTwEriL55jzoB3D2/D7VXTzTUmyhMzwpybmZ9Zh3YRIHGTH75Yblki6v3dxB9aFSQt7/CGd3l
NwpZcVZPCRJeDESD1bUmRriZPgqI56bqNJ4QDJy8WDBiYGfBrTm85Tiwm4fKbUz9H62lU3oq6hHh
3q2JpqT4tRLks4jf9WDpNiHuPKjgsiXvPX97bMcr81/uMEfI3OG35KJhzL0swEptlSNrVZxdu15J
VYSVDFIQYNfCnA7O389MALj9hWpoaJOhh7CcwLirdNiwWlz69WCEimxwGOjgGzt1/3RYJaFI0uHW
fGqyqUYTjXP7/YRm7OAG4nhI7nhSOUVnyHXLUSXJOxavIuTkhLRSh+fD/zYbEh7hLiNeH0UFY5p8
mZ9GfXeKGF6EJMnqxR7XX4YbwfxNfSBGd+39btuKjnrzbAP77NAekKcZ6O6AvBj2xtYzZEFQjmux
aIKL2Wn1LcY1ZpfEbgOudwXkni36h10yPxeh4EtaeC6UuT2eozDZxLmVeJvPXY/pmpbFJlCb73l1
BWfx7uleb0CTHuPfTv1pXuHp3/L+e0TE1VcntHS/18Hstrpk95EtXFd5sT6yWiW+y4fvLTVVfAeV
ot7+GugLpqEy3WidTZhnd57IRBfe6F0w0r7+AnYsT1bCXQ4Vl2j691TomaHW+p7jN5CJXyNdrbFL
T3rn5DU032TSpP+nio4spHjg9h20nfqXk6Gde7B/VrTHKv56NbBycK+JGI0ufFZT/PyNGFTzOpwy
xPmFF/stJIU74obF78VMTAwqTg15W7XxXH/8sA6B05sulvVSYCokIwgsV4neiksUkeVBRj+HcvGx
VRVK89x6VpylMGYuY6vZiz6mhVUrGTiTi25SOqqL5tUxTpC9ydzZsAFHQjRhmiN6NXjJduDqzMWH
FETGezkL9zvl6DuusgeLHTrkzJJ8dEdFsl90TKMKUQwFCIqJHvzwJVbFpurRbRoHy6DFUkbLmSG6
GRHD+79xEtgmp1HQdGT4qS5q37K3VjdpJ6i65Wh/rRKXbQ44pC8FK4p1HyJDfl0FC4iZe6F+ufn4
sh7fCXstMAEamwStJ04w+XeHkfyVWO6MWXIJ9RWYgS+DDJNnY6vpO6YPxHnExmxPxfwSQw0FqeVf
XIHN9KAVIGmGfW+xbR3Ud2iSX2cYzL3I7Loluui5VBWe7FWk4wyMY9+luLPX0DEBHMfMquXr7/8D
ARTsWQrzOzhM537DuwLj/tO54H2wown/GY/2QBueoUOi+WdIly4hAHl+FQewBId7ccpq8AGi2x1O
IOkDMTDHmF7X88VNIUtjHsTWl/2wrF0ir7yyYsoucsR1gXuV1QF1xPcriL0JcScgRBqVwPdpzxrr
KuzyGHCAGLRrB7v1VecWSIs0F7KnRDeBaiSMn5FbfCLV0BCAoG2s0qpsBX9fQea/zR/LyRiuhDCD
WkIDMF7+6vbRSZB4Q22QMnBcXAfP4dX0UVwZg9r3j5VwhrT4gTx/hSmm6YZpVHeH2fVG1nXqb297
waL4VZ5u67RvYm6BeiBXPH3WEHnzKjP3hfHYMAqIpZ9IpKOvWmxCJC//UsjaFusJi3CqakA6c3Qs
N93xxqbXbzAmQMjCodKZuX481j+CMojnD12HUZGPTG2F4g0dRWh89NqFH5SnGd8Eq1k+5A1IKeZ4
7MfEPp5k+eei0Qo3pVHklEBUVECgqy1ESRw17fiPQPnCWz6PveUg0L5uI8F6IFnFujSF6q+KZAK8
EGROWnszdcPQluWDoSLBRfbKS15iilGubOfptaYtLvZmmNKkRpmEtC6UbSZS3VUB2HeZVZYOst4X
erz+kTYQVWOVZpBQc7WTDed/ox5oaSPrutKLVIV0+5N8QjYCoY6J63oKFNQGhv6ohL87y9ZFS3ol
I5fWFcVUQuRdgNp7exAGE+dOJ5zgKn0DH/taqeXBZADozV2eiL8xSdRdfGMG1HMrlklb1scUXkgl
aNH1sJeSzDnrfyV3h5peL/CNuw3q5T25k9ktpJqhtHXpXDwHmqPBokcKyMQxRP52pCfq6tzwcCCR
AWVuBwy+hAorjKJdGF6KMwRxaDChgBf0prDgjrNVEBSd2S5nwvpKF/XBKo3v2KU9hHnbDDdU6dI7
s7rVqffI79vF4kYHB614HHKLLT3OV+FBXpA9tDEN0ABDTGcdc5iREiUrXISw409V6JX6uwy25v4x
UcebGJgE4O19fvcOnbwxGT45ATOqEMpa3fVxADaxGTZ+8Dr2vgCqHusDpK31jrDwIVIX3paCdGeX
PjfBd1eHbIqbKQ7WSZMbo/lcE69T6CNQnxPbN0DtBi1QIfW2k/oiTpM6I8kMrn+Wa4bLrjyO2ZTi
8o4wTDeU4TD68QpnJbPcUSDWyVnB/2ig6zvP0ICdDTXzaTXBWZ/otv7UMnwtNpOOJJTI/9k4EM6d
UWd8UKrlJoU3zHpsGmtYrOazpunW9DH28GIawyOO1ygg1Vp7tkmULEDwuxc6MGbVOEEdiNj3vRFp
ZHb1gUrLcNuISO/i/C8l5A3MajsvAFtrB5H3PyDTXfPjwehogL3s1IG2TuMP+t7k++DUuGSvwWKw
bRBmhGGq/8Sw+Hsg1C8Cvvl7AB/fZLgLTWyP7KSz44HNtIjotdFy3fKwU0HU/2RYpCZSw1fU3c7O
8p1htqoIeLwXFTzoR86KpIBalSspfap22w7Ndalw6RUrlZV5+57BpzBeO0rWEPpUfEZWVBQVeKlm
ug/kXp0asitxm6hELVHRlnRYfshRaxbklUxZfUfFXh5zDMylgLBYPiDwjFPJpcCIdnvkJdG8ukT8
f4x4AdvRYKH4ppeeQeyDWDgOrwZ5AkcBzw9L4hSFXqG1nFa9NvvEuZ1qGuTMLtMJyubWp+wT/WA1
rWymadVrcJ8TD2H7xEjMFzRd5d9wFh2NnME7FNFLXlE3+kUvBf1xCjuP5J8MMScPit/hrZHs1bqr
wGRN/8kh3rj83DPX2DGd4cVLHsR9lKBYAhoRQR6jxYph4O3aFm5drUs/MVxCM2B54APDYA6siOpl
P8PzVTlqNKDfsIVC/kEhX4uJY9ylMZ6qLQtif71L8SYp+fz2wmbYn8KyHTrqOy3FzcL9SoT28lCZ
C0Rl56yehgVczkzsYIX9HdlbyvE7MqqJl0WCaHK7CDZLMxHZtc9WXCP68k2M77ngxd2ZwuWgQMmc
dFw67++SDacqUSX2s0UYSACSBHrB6wjqvJfM/E2hIYdy2MTFiFcgHb/UocYr3ZgZEclMJXe8qWNa
nBuy1L+37oI8gjtg/jFd6oTxa2iI/61yEhARmmTn09bn2rfX+5EE6SpMYhcw1xtJewPsMRCKLKif
cjlboZfZeo8xJOROVxJjFgiYiXjqen1sLOITTDehbUyUluAlmN2qjcVywWVTndcltpVMRefDdf4q
F6r5B+UtpeIktgldUgXMyRV2GEbQx17Xs9pdC+UjFgC+G2IdHH3ilSbHt9t232hlx/DeuiITM+Ak
p9chVnqW129954INXKaf0+m4iQwcmYxDiPF44LTdIlls/KY2Ld4Lk6v4l+OlqUQgoQCy88mfAew3
4PvI59mDewhtgEtyLegIYiQ0OIgHTXVgzYFos3lczhDON+T7oPHIOOt5TRGv6QEOgpnzP9S2YON9
2LLyXK9abbRdWovXi7gtxc+P2Rsj3UdQvH8vBewIkxMGlfgMFCk5p6eDTy5LMh4aYdW4T+/jrNTp
dZOFEdZwf4h/VGtFoFYbKyNX073MpzvyfhLyTfVTaNfkSK7nq2E6tC/Dz4oFMYSdk38Yj906S34m
Bnuxd1tiYK8bWvMZb7IR+nG0+RS93xsT4lNuYZEGHPB56kkXWTSb3AZefPUTINIwoezh6ZZW79qo
hmwNTOJIt6P9RYwAa+wiQDDqlZrIW0MpqRb4qpo+EBu7N//5dhcMxafhTy/+8vEPJZxb20JkDF8p
JvSgeCqjD0GhYt1hJEqaeffZu2xeaSZt/Lk1LBLEXGLXpHozOa5i9FgqwSjMygMafdbVinQ61UmE
TS0aNNB1HXc1CgBChfuFGqeDQjWSSzLGRDaQK7kLkZBoV0suMTbWgIUOpmlUQfRG8cRRBA9bsNcV
1d1vsLog+fPnzhrVZ3/LCyYZNKfw6j8qlnIXZG5LD4wvrqbg5NLZfwbfAiCAGDTQLsFIzBeIzIAm
1V0rMHYFqRE8p0FgLfFRBUgK5H4rQvMSXZeNnYBXlr0jX+CKmOmobEAArVDlYxJt3XH26/ih9xGJ
uS4x+/YO3D9hk/XirhcP7t9ZFT1bkHz6yWlbPlDiXiKpUtuWNVRdDgQGtdxya6p7JJ/uo2WbkXi7
r3U7kIA1yMK+K2CivjTGwtwewbbaRGWoGwzDfSkRELbucSxTusAT/6XuvK1T6jrheX1Z/7Z+zB98
B8H6vKzY5ymc0f6HkV9yZ4eapx3LiTVTbT7AJtCWc1wT8rt+uFAMM8ALBbRd2rDn4gjPjAsgzRXI
zUT7pYrhIU+XouorDdAll1jXLT5mQP0qjjinZ7T5mEaYTclyrNHUcCgoXpMCgJHnKTTPRqwSl5eS
B4gs0uYohp39y8IN1PUGlx1pYUmRJsgLgWFDqFrqaiR/yThOKti2idbJmFt6K/HXNebe1revsZZH
qiV+CKz+Lh6AC68OhQru41ozH5c6gxeTW4VuFWg6lTL+B47/7n0SFVBRC/SunRmh64HoJzVDIEp0
DJBCcm2FrfI6hqKIEjLJoi2PMiLoCEsyAdcE18Rg77dpmzGfbJ3u2GuElwNuFPkxDQ3y2NJGTn5k
JavIm+sdt4c8VnadLlDdRttwL4Nin72Fd8jW0c6X+bc1EJZJUBToexehmzIx0OtQnGtid83Rxeo1
a5GW1ZJFM94afAUz8R65Tmg2sFmDhLM70u1IaW25Cu8YHSsZqRgpRzHF5WVIV7GwRRei3JrAyz8H
YL+Tuf5pGxWsDcVres9AQSo8dJp7ZnTPZruBBWzU/T9oE/EWFP/AF4zF6pvQR+OCI94rTnw5H1I6
xx1ujQV4YPsQmx5cOsKz5fpjoOkheQsNgDxYVRlQm1eWPJEUHSOo+5tEve35HxqDHie5HRCkM6vo
ES/0ezIo7yoAbvJ/xX/aR1DBhkvSX5ONtpAr11gbLtDi006OBnNisQM5enQy08XvRY+QdnlKnT39
alp2fbhS9JUcgxJCGDm3JQZJaU9wy+cR/mGk+SPQNy3wzGBUBXNsxe612MhoCUcMfYI1N9aOzs4g
nyg5u52xqkssKQjNBYWa8ZLH8BHd8zspW+IfCRxADQGE8pzNdr1JUs+RYBVaD/zx9kLIiB3VjEEQ
IRWcfnOi1JTtk467gCJdICCPkDgTSCLZJdbgx4cQ8UuPycBTlzTxz9kw7gSQFy/VjprWhiqflmpo
aGmMXOHO3EWxQtLcSHeM0R0TkZOMjnpc/nx/HVpXvXHgmijWAnvEUPu0P3Ay1N9WdQDTOISSqPx+
IMCuJFUtQbyK/YtlLJeFtfCRUA6q/6dXKhihoLPmrPvL/hbNhFF6Gxb4coHz+T27fgJx1CbtOeoJ
1G9PgA/U+VWT5yorgi0r3XNn3m61YCQYFy2DyJcCwgQV4EqF9EiTmHg7TUz3XS86Zf6gGmFJC6vX
oP0UraVeOLJLJAKQ+dAZgrDMdMBkoftT6o0QkXAf6a+gyOR9Aam864DFTFtotFAEcIUQuQHsgddj
u26Ud5fqEHrfIQyQLUriWxb0IHOwWqWfFRbSWT6jbAtlBsBnwI+Koi+jQW03JsKtw3m4Bv8gRX4F
7FSOS/T+urZtS2LP4bLXEpRgMa11u6iQqEAZIpYib0b07auP/yFda+x5jj2j+g6i/5L+I39vRSoF
IAhJZIiVp7FvAIqahzhep7qunRrWK0K+A4aKFe8Tu2QKQf8WKlnFX4fypwbpUG1RUJ6+6Nl3CXHh
LoMiFXvnsyvq9vnKvA3OMlPUqk69LKtiGsAHYL/XTIoQGZQ7btuuyEMqoRuLhubLaL1nDAkTLpVu
IsA+KghXxNizDUNFHXA6M2XRnH1SPa0JpU+pqpUgqqIz0/GQiwETvYQyquS8Yb3FMZg1eXP1HmRH
btUe4SeUPxQXHU9+bqk120RbSb86m3MHcj3o9Sc6zUV6pvrvBk3rtzU7VwKfvOHXpx+VOq/E6Y1/
3UjhZJ/OpK15tQ9u3Q0kz6yYMp3yuqRsTkNlo4YIlEG/DyKSgeO6uD2wx6Lrh8ipRtu9s8ZkfcXS
OxFJFm9313X4zSW0vlIt7Ep2QZlzVL/EnRdK8fYjk7O8ELhSIrmTCKBI51WpSZJGXALKOaJGClak
I4jk9U5dMzIV8yUtvbZ8bzoUOFgth6BvI95N76mlWMoq2q/hGnMJT3jw3L/OM6SdVNYhwJfMRfWJ
VTf6O1xE0BtiZnousujb0JKklsQzRaCduNHjRAD7GmI8tlc2Y8TskiCTjJ/pHNcdx85IsSunHxsT
CHJ8Bd2XFeGmYrxWac3EGUR+0J34hsEJT+r1kAxi7jdmmEcZayqfuQNWncL8mmULaZtbxeklACpn
d4Oe1z5ZgM8vmsc9S0ImhShzBATFBs0xAqOLEMFFbKxXEWSIW5wUucKiouX27Fd+iT9BmW+BQvxe
cgRbMFoNYJWLHVBQnJg+J60TbYifXucFBmexyIKBACOM/yqZRvHwq5lxnuD7pHg9yDzAiyWpRs7B
ft0VoD1hUbZnrbrIm0Ls+zNd3aid1EAfk3umrZaVyapZQ5qRZx4TBwRykgSV3DBETrcAFLy4Qf1Z
gsXTLD6nfQ1xvsx1qe0n+RYEXrqmepW49B7OYaHRzzB+OO35qegvnhTUrJY08a8KuMBNzV1ECCnZ
JSJc1AwtNwT3PviKu/NYyOMOCz0VwXjy3RJ6rmkoWrs7szpkqEMIGWTLGfLXfvcWvXxIc4eK8WZc
VrVSqqSYIyo4xFCApwwVjHKchVaLPKleecc3OQNVUTBCurvzskinJGQwXpxmBHbIKzFs1Zn6jhBb
DXFllf3FxkGPQWEGw6E+sBFtGGUzPGrVJNh/mxMb5L3mnmXwMzz6vc8uGcs6nCzprHaH5+eM9TR4
4kRqKlw8mWk3UnabPiqtWTzozB5bBtT0VNDVq3PzkbZ3mcL4usiZ3CFlgX1nluAbc52IUUgw3vKL
kQZWXOnWf+aGmkrPoOxUOAzqPqM9XmbyJDS22dRfhnySHm2Ul5Rd2GI9N/uAMjhRd9O0KiqCaa0V
cHcp/gM5sODBQMSX53PcYxN+MaEeS8w0ma/k/ksSwDfd6v1AN7+uy5Um/AIcFWwS5ZfcKuX2UzOF
hj9CR6CdtMXMmz9wQeXZUBFfMw87h8GzkOlUTmEV6r4qCQ3T+LP9Nx9dSpSzMwqa/aIo6vfMxSMw
ka3qJ5BLB/R1garC5r3OhUkNk9sg03NRvgo96timhVrI6AHSQMtjK+7M64VvXWS2wsgmXZ0Um74g
djq/ioM25jBhQQib5R8od+B7O7IJOsc7+4dWQaxAYugZVgT5jlLqsyv24stjv4RMV6mStuR8A5+o
Rtdk4ETafx2PCK2WmHVtTySQsn35PPSJiRbyEuLtUnS4zuH+iH71ZONJ2epz2hZJjMuFpZXrqL6J
Xr26BQoLv0ODZVZcWo6w1OU2tcO+JalhYsk4ymX18AHV/TRDn/LlkpS/jac13d2aOCGN+HD8WVF1
AaFjkZEHelowMNas3wEGXTPPBDQZnreysftcNR5QJ/TTl8uBeh2YQsRfO9i2cf8sRCc6EI1LepC4
/Dwn5xS6kZscdFr8/Ct0WpykuYrtiYBuUqHmakxRPfunMlZviEyHN9PX9USlzmWKOZCFJb5bE3Qv
GtrOiflXCofA/bbDvnw1Z1+7EtEvwnrgYsuPBm5KvjpnsgKXoqeOkzOKsi0vBU9ad9nLWEI0Fvha
bMYL6rBD7OpXleBDE2nA0bA7XFDZBcQsdFsijgQ+nwcOWjpO7wZOnlafWhS4SoS8LVtsq9hiqBi5
+GP7NuF2joY58Igmv2gTO6wTIDaJTrB2U+F/jpqi3hn2Ep9uLTjO+IcWHpK2WKyriEDseWCcG33t
vBGGViz+cywyHGawmNUDiksHacc4msa+vyjAo3Oi46svyyLMKXuPXTSiWkyp/puhhNHCfhJ4Cona
23QTefARGT9/kAV7dMICoKnqcur8tSU0cvLX/Zl6MjUtsBkFOrGEQD0JrY+c4FZ0ToJn4Fr7aMgy
4lg4Y3rhA7mafHxIgVdCgjzhGUkTF8/Xt+Tx2eAWYQrcEc+yQVipbA2UBY3QYj4rB5IodFy13qnq
Wj5l6Y21kxT0pAIc9yLc73Dlg1bfVV90zx427lTmIEjHygYVGh41+q7SAGanZ7m6nDRrmKRcAhpw
kxfzpbOjbvdAimaaHz+k4+ls847jBE6ecPYVF4Cv9hz47pSqRrsPWVZecQn3HJo9Wza+LbIppRj6
ZvWU54LQrUNneroVDdy7GwVwkFz6JrTYknf0CJC5w/1OJaouzQ+vXGb+nPXJyFZQ/Bzq8xgjlIC8
5r06cGhU8IeVoJNFx/U9ZsX2p9F0sVGRKhLu4I3ZLd63S12YS+sH3YxHkM7VCFBYBmd8+ApDGugn
eqwlM0P3Q2DiVcXEfdboJ2tvaecoDn86jWRnR8hQzAiMFi5eSsXaU8DEcKX3PdAFsrA0a4pcRDrZ
Lr9IjWBxfbPgQalML8xtGWv2BSnogZQr2ETH29UYdBDNJOU7ahhxM3yAu2+PqkNfGYDoemJnDOZr
36X3GzAEMW1pr2RvVUj0Wye+l2kpfvZXc6YGVkS51sPpV9A6Ix8yNpdJ0WC21WGbnbl8+Ik5wsdm
duqTCjt2WIQxBM8M+lwxx0hyDTMFQtdWEPQJb6oSKiqgtl/wk8s71p0MIEo09mcyGOr5RdAk0F2N
ARJDVnH9iz5genvRbrQ6zFTFHji7X26wO0QO2l699qHQU2kDphSZqZiNicAxKhIwPM8tAD2yLpX6
mPEXcpS+goDXehqig59ysLSMwPOAn9wQfg6ly5aBauS9ZOS/8znCAXKCRNfN0Md4wYYfcKsw2GCS
Ysggbs3LkkYVuRepnGrgmlD/LcET8bhS0i3JUxUcx6OPIXdSKrBAHmEp4CrpgrNfjy1ssXgwBhVl
kVp2kzjtmWa/g52pEzeelExQi3G7P6E044Tzifawk1nigG9yeLjK9sZOEtjbq0wdn33g/sKRjdbB
c+lyJLg/G6G4FqBngEmfCMgcQQG9ZHEivxP4saLsaDW2upbS1gr+dfX0D3M9+Krc939v5wcz32gU
P61atysy8db635dPO511udNncY8P8RUeLZBY1V6OKu42DdlWn92lhho/jKo/ZAPHvWkej5WaWJa0
1I1exNDnYMzxdK/99N75tcrbYKiBalxMtyrkhNBreeEXnCdrxTVLxDsqGyypNF+uMySTE0e2yR/T
9JOJldfu0w==
`pragma protect end_protected
