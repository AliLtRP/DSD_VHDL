// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ru9W6jLuLhmWedJmN/N9zPYCqRmmplZhHJ3i1y7s9756w3tlA9sGIux4XV/ZdxaF
vpryVFpHvHsn5dOg1ILYnAFKxKtKY4aCSiATSI3G0gMuhX9kcgITp2QJ6KCc7dIw
tMOksf63r5anAvMyUU4fh/2alA2/YADHRZE33z0Pid4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6608)
fdT3vsvovKeJCe4UphoxZF3wfT3gyaY2jEQW9WWtApRs0+73P+BYF/iE2mYGIURu
Ao6x6UOIajkPhrAcba1xplrKmJu1S0gX+qz6Szhm/tHU9XD3Bk0+auCCwdWkAYzl
SypIG8QD41/z5UlwjSFjc4us0J68SGJYzdiYsMzR+uzbz4Sy01N4/cgPZo/NzQ3U
VT72EbdTyRvqqhCyhpXgNbYldMaSlzQs5Iy3PWxvpJ07bfg+aGU6M+VLZ1gWNDxi
ft9kDA0nmzXZyDrc9MplaCynSXsdtGJ802fRJyxTQj832QWDP92ru2tEsl9NjWrx
5RH+fvNaX+eYpsDDgjWjA2lii+IZh0OkwNDtuaxut/FPiSeRIVJ5hG1EFikICfyr
l5xK/R0+ECiMiSdVhNwN6nGrbP8YjCZSYy9YDjNqfIzjW2mfPU8bpCLeYMCVeuSP
JF2OAeW3gy6z0AD3ximSTecDVkN/ROlUQEtEMCUiGCc4qXDgHrrVyacZqI6z+6S6
xErMDCWC3UKwihLmNgN9rMGcyHGsz2W23CESljQoh5E1XMR9QbUH1RrAygARWB//
I/2LApzJbZAfvvlxu+CmbbuOrrVQEj2PT2D+uJByEyiKnkjgcPX0P3BKKy4elLGq
41U0vzaZY3yBM1RK3D8PuMNsbMuJh2GdtbTyaOJgUnDSbfnwCQYDYHa2tk343hCY
tBJAMicj8+lKlsMV8t8fXz3wlSKUpz345+X5QDEKU8MQrDnMxm/COELjKVi2nLBV
N5nC4TT9iZvKd5TLe/gPcrRicsouJM3wNMSLFGpdTgfnCHSX/W8iLqj+93ULEwGk
xurgUHCWkXx/P23mg7a33MJs2hhXxU1DU1J9EYHGJ4pzpUXr6YnF0hv8DZcBTasc
fV6H2i0QGh8bK8fRlNmzSr9/tBDqFSFwQkhye1RWPXByy2XPdlQohYlXPp+tSyYn
v8mktG07clmSYiQGPHZO496zyTShhBtWXjhXMaZVZdWcaTIWg40UwPdBNoR51CNQ
l3XTKJ/NeR4D2nHPAbbPvmNkQ9VxFvoW7QLUFK5BgYQNpszIpN74DBJWpLAGlgWi
Q/UNFfJgxKs1ziNRrQ9fcSmZHajBobML6a4gSdAIbG5HbNyO1U0KNZ+35emDstqt
H+D6t282NdGXGYmZ5QkGcCzmBChdASNdRG2WtAUQ5wjmmV3LC0iCQbWtVg9Nmsx6
MDZInEZNmQF1QTNYyIBxXhxH2BXoXHlecB+dkLkIlw5bBV/HbdUJwk5RpfyK9Tj3
RZ2o0aFQERZZ/LNxUlDvorOBja7TxoO+5qXnBX5oZ55/KmQETxRv+MRG1txhogb+
+MaqztOXdOAy09vzsBCJESOl6oBAOFJXo9A2gSoKN0tZqdgFkPHBwHDFiDyRzpCR
KwiR+et7Mgue9PQ1YFitcWruvtI/UyrYdtb1pS3YvFhMPPT0uPG+TFUp9Zk2kGWs
nqS+Z3TLJlMTTb/xXrVAnJi2J+pM21k8leojxx0hJYF1V9MvScz7OQxMRHtrQegf
Tv23UbsZrtUo/cW12NTaZ8SwkvJQ7s4cNUs3dsIbbN77sk7L7ERjDywt9AEBAQf/
sBmxHXKHoWraPxg4bmlwbf1pmbpJs4Ql/6KyJ1GqPPClRzBk4gfn5AH/2iUW7AP9
yDc2eKUj53LmEzFxeH7jYdVFAxBoAxxEGk17ICF12+qEKgrGp9s2GnMA5uJvq/3B
5TwZll/rrD8fom8t/EaBezp35O2UPagg3ldg+2GPhP8vlG7rbAy7pJDJZ/htPngT
+HQoIN39gfH1AlO1ZTNHDNBssieNfHuFFanyLNgk9XqHE1T4HnvJQqQV8T2a/kZF
CKa9YvKL2SQNK6j4U5g3ji/tMlv18xF6TqmzT5v9UD22xWJgHywneuw56q6DraG3
LhQOVx6Y+0x4FHPePJMCs/dNDh/cI8b2VKe627UwZ1UoW/s+Ac5LXHzz7akLgJa4
37V8JiO+2wj62CAOkM+/e1GoeDd2N8e9OTsMyiOWr4h84JL8VtQRXsDHAvgRaZ1v
YMC+ivywNeivj0B2MyRHApKUcShMdV+ucdUn0do6t8ZucFiUkNZK0cjQEhabhn41
96n8gAV7wNyXOQ6ChWja1OMbJCZ03Ld0Gt/WjqgDVZufV6o2FFkzl/ALLVbIsfAt
+RF3FGsWG0yu4079wONZJZcU9nLzdo1TTSTyKMHpDY/5lBV7xEfbMRa9y9j1kTry
6OuSSlpMIStaCES8ZHv1zDKAX0lXzl6GOzRHbHVF90K/p4+87Z+VWhMZYoPSJ0Dn
Y11l7e71OJocpFzIa7gmamfIbqajIl/grwkaei25eRgYdjANiaQkYLztRWpQ4/HO
JODgIYI+MiGS7Vmmg6pLtiIpZSuaMlrDOilR4j+B17RMtgLnXG3Z1lLVYtInELit
C+LkPN0saOhxbCluWzF9hi7HFL/kDvyDIcPE1wtB62sdojDdNMbnhZt0K5h+aPsM
V4vSzU4t5XEyGrtdL84W1APQPZ+YhBfeS/2eeC6Dmche0SDHR+aKZrhWLjIDUGIC
70ENiJw8gY9NtEcIM8DZyH+G0Rc4IzpWm9QQVDe7IFDFUUr7ZDi4LcT8V6XOUpO6
9B54Lbf9afQLF6+S5GQERmHmLimqo6fDXlxwm7T3iT3+Tzp1Ry7PziqEcWm7DlVo
ALmczFPYYAVspFgXvaVvTUGin9pwC7jjN701rQ4VlpHsdG30ygVa+Bp+x1vWLFKB
v9ph17HzKGBDeD2iU8Xb2+wFzQ3IqJPLZ/MMs4vmoT8DZndjY8czRIw4c+0yqYJp
ecK33WRNNIVQPP+Smqbu39MaBIOF54VDqND9vzPgZNsQdyogM4PBUD8UG5kYDw1f
bQFo6Z2HbxS2/X31qS5lTC1qJk7Co2glTs6gJcBecjrIUl8rVE8ebeNWEiMU625W
NLHI979Dv29n05ecbHKL26Zq1+C2FF01J7FAGqnxjUwr3vNMeBvfPQ0on2MUM4Eq
kzA7ony3Cb9D/gv7TZocWO6h3ZIG4S0oTefMzSOvjRJHzWi9Dsv3WKzwEJCwvHYn
On/sM1bAknxvioyw10JL/noXpyHi4OuiLdAcjWgEmgbHOXFp+orQ1Ix5Jr2Rx6qv
MBkMQtizmZBxrbi+sHJ9PRV1+0RpzTbiCXnyer3KJsdJFGZDQIeKWIw9Ny+fER6M
CTL39jI+wgD0Q5zK8xj9VSWpoJBPS+VZ1KMKmX2e7HZuOp1RTyU3cS+2t/1S8VSZ
wUnGYQP8EUfB4unHa4WJocf31Zx3Z5lF0z/pg3PRevELIto45jQ92uamEZsL/C7k
om+X6nCZDCgDRyZgyUv3O65jNJkqz/09hFWYA9k1gkV1qwq+Gj9i9auRDWDwmtA5
fSG1FQZxFgtLr2WPdXy59N/YTJ8Va0UQer6ASNcYbMYbLUcfdF1wSgmSKF9EpztM
vJYaBesV+9E+jYJMc/5FGzavYaGOTBGQo9nqEs2J0i3XOV5QDejHsZC3t8dfSgZ3
MrdAJTgyLKb/1a82fx4ZdcgH5avnPVARGA8KKIro0v8cEZjtyd8M2hvJv5QnuEim
GKxwN4m0HbiYIJ5/xkarLrAiYpRilWFjPiXnFyPgAG7OmW6mb4Zd3yTE0FqWR+Mo
05u1flgFuWifMP9Gdbi+6f9qxh9J744FRKqfPeDUUzjfchlYEpqFzOqF4a6n2kZb
XkHw+wFDOUfxvMZV9tZ05iHcxVzzr6re8Nh+V0we1sRyFaxKU7/322zZKMV0odBk
ADqPBd9cM/msNlA+/vFjVXaB/tygvbSlf4DkKt+5Gb8SpFpTG8fJrH+xT/fzaOh2
WW1nIezE41MFKqU6WBZQg79JSZbcLxBYkbBlX/t1IXhKrpIhxLEi0Bycb6HNrJ0p
uifggNx0UV7jig554lAMEH6dE8+vSHdgpLhvy3Tk1JrQ9Syp+9mYfukAPXq9Mi3y
gvcv1P/SEFAKMJTkq1yT5whxPJkc3Q4ITbXG3ubxYxLdceYTlgbofFdXd9tygF/2
2sEt1REhChTcjH58pSDTLU31JabKbi5+65yyUKMaASxFQFFORw3UQU7+Ke19ZJT8
Hb+pf1ontfE1LkvnyRvW5eksi2tlMVC50D5Mgmm+eU77M5CeW11PjG6rnP+7U6gD
AO4YZoAFYm1Up9TizBa0/p3Z4Dr1Nn3g87ijYoyTZE5ICeLNEm5jeOn4kuaV1tS9
3bnH75956R77sm6MWBp9GDwfsiYwYL5Bj7NSn6MHsag1Ef/euSVWlvSTu/Gmgbar
e/dQ4lM5poun8EXrqBirqL3PeDSYBgVLgAnsD1TfjJznh4BZTq+WLNZDjeMUw1d9
UJdKadP8By8IVH/CYWR6d3O/hONcr9xD84hnpgbaL8S0CcrJEdFZUA9UbWqomH6i
THw7Sin/rpsc64lUki3epVAhiKkuXZOiaboGWDH0mA2vp2Qs2Ak75tVYONuFK6bP
xhASq/SfrOuT5E6FXeiTSI+OrpO5CJhPXHH2GHlFJSFynyyKw74tGrwsnRcRUmHa
7Ga4x8cZmxkOJ/8jTtLFPVcAqzC0DQJwOkjesad7hqUYVx2MHYvMbyHTnPLICX8H
uyA9nCKEg3q0VfctSx++wzEFdb/jfp10SK6y/D7PZChAc5KC5CSun3Q6c3/u/F8z
VxxTEd50UQCZSwty0poIWZCkAdw6Ab89FD8Uo+julIpaOHUmHPHV83nMX56LVV1K
y1RfOogMceTZtqiDHekjK/IR1akW67q9vlMtu3rYAj3wbHQA7tjKEmNaKjfvQpt/
v3wJoTxivkrEhDpt4Z2XCzG6DPhjxIYIwugjuXkxvdwFSAn/KQuRag/TIEmeuoYd
3lVqt71kmYVTwLeMnShIJuKkujVtmVqr7jLbsLImx/TKu6abGCELFe5uLLxzfXx7
wRv4lwAOTpnMSXNvWZOjSs7wt+Mkjl+zcJwPQ27BkB7nn20OUa1IEkoT8nYBfJCz
UFW3e+pt9cTC8Ojy9p5wYH6a3zuRU/pHdy+Q+p7/kNeJblATgi+gHgjd8MWPgHY+
Jpz6i/7KIfBlSCzJ4ije8lub8IIwAF3Ee/VGH3S99Ukv09pipLM1/uKitOXw4Lqe
EL1Qo2qYzs4xy5CwKQhaG2fcSlXfu+ULQieXJmxqxUsVpM/qdZAmsszNhOzi+thG
zzubVX3JlxfUyGgLrHHyjKQKv7JgaRfLVnC0Y2zIz2tovEzuBC9Q20zpRPuuXgB7
/sOgXdDl70EdPNW8l7JbmY4svpVjZx4jPRrpPRFMg5X2isII0R+JOLihxmQSPjUw
VzxINr/PUEBPptLZWyfDd34xWKRvPdNkU3avi9GdMmf5jlkRFDSmltOrgtd70/Gn
+Od/SMjuVhgsX/PR8tVYIKRhbLLz4VOecK/ElfVQN9pvYpNIqgt+E2147XZ0Rhux
DbKaBwFERwNFcO6uWeBLyuazHsEw3vQqk/3CWWKqfc5Bze0nW1Z9OYuX/OF6T30U
Jo41jdP+x2l04FiJyJJVWKKKPDuXH1PTVKS/qC1BeSEuHhLWXJBmSlau+MPGhkXY
d2FxKSqljIIHR7Rp0HEBNwaUFv9KGnpQlT4PkLhU0i4AazuqJaNYQYAXdy8hZiON
x3hO8+FuzAXujeh6e2dRwYzQpoozz+SziViWXQEK0w5oNRchcwrdXWNJBWyHiXWr
VTARCpLr7ZS0hQb1lIIa8KfBoPk0w9ZX+XoX62rIUy2Oc8F6G2yqirW6p7bBPVug
ezEZoIWNV//T9CZQfstljpqVEPJYX6WNcizdjZZCm0K0w0BlkSlV8LpBomix7Ifk
/FdjkQmZXoR+VtC31/8wWyNdeBcQ03tQyjK4EzB/oZshwbfsDU0iTFMLfbqYe0/n
U+Wgx4LE86dCcahYjv8696I3Q8IVvjQ8txmUhO9jsTep4W4UaUin70soeTgU9KbY
nK5XlxN2en+OYNOpxnQ6BMgV3YF9QbUXkAODNvyy64dDe7WpMqjw2jD5vi7nY3im
26tsGDG9XERh6VxeLeElwWttOGUTnMc3D1h8CsT6G4dDRBnUMTh2LVOKpZRrHpLg
0Zy1SrVMIAc8hZ6RqGCN0YwI3TFk3ju7AuyjLlWu8Ga12GM17pGRdj3bLV6sbadW
Pb3QC8OmOtK8gHsLNy/d3o6cDbjJavYpezCHsRFqFViA690GwK/01a/Da6YHVISE
daAE00CNvqbBueLqfSZIeeRHWnPkJHXCKe0pD5OPXhJ68Io+NS6icFFJ1wNFQ2HT
hM1Y/J2SxZTX+gS89MT5zSQpGlRxXbcR1+HrmFC4x8biutYsHh2p+jY/Z8AuzHSE
MxA3RDnnUE4eN7RRLR8ukQ0OMbssvwEbe/SiT6aNb+n5GkmFH6u71++n5UHcwIfI
Ht9P8DZdca6QGCqdBw98Sxmcor6rJYKNZWBCW8NnG/tRJBJLWN2SWnoDO5pfTUJK
+H2SP38itGkcjCoDpKbaO9bHVvgbOh8wyhfgb++MuyY/3YQ4nYTzk43Gs9Lj0lIN
yY0Jm1OQDDmJWQzfl7rnzO7vzTlv4mxjNORGb6W4R6WJuqaQIQ73OJ7EllZD4HuV
Bdit1UnIW0KXGerVXfOm8TCjqGcKkqKM0tj/bgmM7+9qraldoZ0eRe539mBGyxAw
7f5O0vT4s80qnD8w5b8VCF9k7aCTReuSC6N6L32JeA45R6+9nIX8GC8QO0BtIG8A
6oxT3D9PW72/jGYinvNG5zkmpxSWP3ca7pswEdTOe+NAK4OtMcBQLtbiIIsMhSP0
k8/DBtKxlSOEV1cBS45wBZ7QnUZIUl+cdeT7YhRy1f7F3rqvHlaP7OjzaXbVIHM1
pxJVmJp9w+TLTbIFbby2oxhUbheeJTIiyoUH+Zt7AkSwwK9Au7eS3egCIIBhpm2m
/LY/vMSZ4M3f+lBSzHYhPw8d6gLKWz2tk/vR/gqe6uMO+aWQ9qulb6iVetw4OFyX
cFUZKh/27CU/ke0PP81J30QPAiCrRJNQvd/al0kb7SFkqNBdpOqZtW4OYmjmLkUe
01YtuSw5sGeg3pEVkeITRJNcz67S8RSMrgKRxM4taIVXvoSnS7OQ9D9WJkulUW3b
y+7ss1lKJb4VDuCJb+ne6wzOzuz7GGjmVlrWwXCkSpQ9aeK5IROdxzEsyUX4yxmv
oEmDIoJrwCXfmyk4Fd1d4KQFNLMWShO73oqYTRW6u7yM6ISLZlcIULcpwe40qTgQ
XU64oup6o2x3rTsJw3zYy+Me5eUf202XKjW04So0gCHQkx+qm7qbgYeWDal+23V4
QBbzaTcYuJ3JVCsUCggieeyw/QoVFTMyVQTYbxyxKeysopscupjWZUj6q/FCUeDj
twenXuhEeT7vlZHPPg2mzl/VT3KPoK3GCl1ubf5kGuD/RrNaQVWeRZmM02lF/v16
nzX2X7+7N5KFeP335saZ5MaCaDWpk7ye1ELQG8fWPWyZkMQafPa5E+ALttk52DqC
KaNbEtJ5o5nIvRWtkUxRURmgCfuWobG711/rRZzKCD6gbf74izB75J+iq/q7wbZv
udORqnhXUwfDY4VAoeKUHQmg0HY2bBfSP/zD1crD84A8x3QOt6Nrn+bzW7D7SUZr
azy+8eJQrR6HcDuyHVevIxVbc67ksU1ZpVaR1XsxICn0SzURUbf7ZgRrlH79lCWI
nkM3U6g9kuLInyEIAVLDKnlZqWDT2O09CQZNfsikygXTecqcr58PF1CmkLP8OnNr
hcwSFMfqiOhVrtI7oibahElMsZxlPzzZ0x7iOh2/M61lDNii3CtFqGeXXgcHm7J6
CF57xs46gHwKFrYj9RNMXVUzpd/QqQRK8mKRkSel83gXibYLp45ihbSQFJsYecR2
lnwcqomnf6TIkj2Ey7DQqy1EPvc2ZnEuMJnFpEGl1t95CiBI23aDrAXAxEZwcmVY
pLfhGys0wHi1FpL8yUo+ojmFCBrdPDw1Sf+s6qZNttKlf7BWCx3xBeUOoGgE3eyI
/3GoPT5ZgqbHqcyTA4J/aUqmaXZdPjE1f93IF64d2JZAl61ZCnTq98PzMfuTuDJN
P/HMaHYqbygZiEc58JOH2eKmbSNqgI1fBcjmLUf163q7LddT5Vsv6SuJDwSNCewa
QnU9QciHCmDJosfkdjRuHi6L1fF4mSNo7JuqvcJsVR4FxVvCP2GDHKP1+ZoGrVXA
NgGLRUnt4eDML6J8VFxlaB0Lnj3Egk+g7RZvSd7UJT5X5E5+ZjD9AXMO+jGYells
t4pkYC1sTx4aiqcLBkfCXpAzrrfczMw3ASEIsBGARnqYZMlLgnHuiikbFxYK/uB5
jphigvgzD63gmsdOa74R+oeM0bqtA8u7xtcYMCFTOQlEzyGcu7CMRwv0TaYPNe80
sdxNLaig71dBkWVYGY3vpqqpaoLgY4hrUBJ2Bu1eqjyQVXiSmQxKPNCL4jevjdWY
QHE6MhXglJ73rVdzANGDAdAA52SPkfn/6BrOmYk9z8CHZy89lqNr+FHkSNztqEEI
6SNyr2aua28J5+95Nwv5ImVOSGBNANChpBJi1vJp6+yfvanqU1EyU5CaR+89am2/
oIaHnIU0DuLAJszAHIXnW1vs2fnS3fzunyT750WyQDQ95RPfT93S+HBYRvX0slTt
fBzitgL4PFDaUKAmiO/rGBxeqvspCKT2QXWZUEtX4hijPqKgpny8NsjfDYOALGUk
CJSttdcvR/QMInhsvxIEGBvJf7md2R7D/aKPJ4wMgHsIp1Ro8COIZ4seOSqrX7Wi
0YFAkwj1VHbFm4c4/kSukYXtBDC2som1RI9E0nxFduY=
`pragma protect end_protected
