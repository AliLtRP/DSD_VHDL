// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T5f2610arXddiU2RMIGJrud/qSpMB6/2GqJvO8Y3TFgpCX+twW2NXu2aqu05eeeh
1uqSkmJgXUolGdd/OFaozSbvpaW5+f4t701v28blGQMnyEpYmXMlc9a0OG5wDCT0
eUDjC4AdW3a22RkHSERpVbxS/HLDkQmTHi9Y7Zr6tsw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28176)
DqwOJ141udw3w0eRYqgOxwws9BTaXkRNC8TYvueBlR51zwd2L7IvufZiCqG97nYK
PxP/8xpJVDxdqqmCoLMXBejw2X1HDWPm9ICI9PrUWVFCdgQxdqbOUffFxvyZQCcH
P6Gnm7TgpWcbCMGkHmV54rUIBWGYfABASOnfKNJSOcNcI6ntud2+c+OyW6NG7ZBJ
t+Zx04s7B7x6mBumBfNn7NDZlo80L5KyGNNg6wpiTqKqb/fAwEYeGz8Jh8pkFw1k
HPVmwfG+JK6Qerel0VYU6Gz2cPFPQbx3kkpVfQl6n1U2SvK8cxHcBV8N+o/MxDWA
S+EUz6fWMv1L00GlzWYz6mwGISQI0Ze3fPjeXLPsdhx5Mgi82CzojuzrS+2AMJfk
uAzVDTdJ4TnwWWo9TbE7O3Px5vQbZUcOrPi5XoBbKgAeV9wLHEeW6MbjJCTs3wFB
PfQL/UQ22eippwYRxJMtlgcoj/flctJgzVEMD/huKSYkP1GVENgeqrZ1Hht97djS
0vmr9riskRI1HcauHuh7e0n9X11UBP5Vg2fkj+yb1e33tU2HQFYmZgwmmn4Kaupr
hXh3pxk4UJ4j8SYqEcQ7XEunHKT59ZPee49uVReRGSoHv94cPXgebqJ2f6YW6tbq
+0wzZ95vg6UWc+XlJcZR6iUJ4JB+Eu228ueiA1rWhkjfKE+iTERMk6ASfbrdRB2t
r91fWA3QZfZh41ZtOD4vs6yiz2S2Qap64EvKIMbuz2ufs4xRWzt/+pVoRKDUgJ+R
nw2i41XGJ6f+W4JSxZ1FY5EYGTaBQ+c+Gktv20ic/pRHrTqGYt7KHuanBcCeHaqT
tsMZZdadaVutSxCdiBuVDpqqwlBV0MxsE5l15fnqLVsQw0Kr5rU1ssBHNdKmBbOv
pzXRt2ICC3Gs1RD/lp6/Pr6tyJ01b+ync9c37W4jSQ5H/3mUOgRa9QL8xYYHOiIb
QXWtmvL038gF2SF71qpAFpW6X94X3eWiy2FZz8EJmlx4xMMetCNvrRCfeeNsYtqg
j/+u9I0ASSraYkX69gKtqPZXTW8vb5dkB83EK/+eJPVOuzVHSccBHFgb0gopWSfX
qmUo3+y2c8YzjjcQ0cXacA7FOu7vieighc/yI9rG/TO6wiHI8YpB4IHrit0DnGfx
jKCBhWvIuEPVYTMSnHuQLMV9u0vQepcXzmXA2lcV9z8w7yyjmEjfiLlePBfEgfWS
CGsIbQ/5XLWsIm0xFgftGywUiNJOwwZoISaW7LL5pvZ/Qt4T12ij5EL/JXwSUheK
d6TzTZB/1PiSn7gnahpNzhSua64JHoJe0wrRbdxhfqXdQKwLNr1lrLhYN/2Y03ov
WHiXngd/tl4009IbsT2vkHjzNKwMvZLv0GLpA7TXFbRArQ7KF8moO4mpjbocVRS+
F51V4wQElcQHfF/iNtlzJOZQY2VrKToecU1t7VttnreD6+YQ9cUaNfgIbMeQcw6c
RoScCM8HoqBOG8X1Q9vyJgi0kx+zslhKw1HFch1C4qrjU6rOycp9+q1A5EYEIsiA
7asuxa61tQkZ3CGy8qRqYx0mB+8zzge9dYkQOu+bz5M6+y/RdTvnZf3EedN1giqA
EgOSXF9W7qgMSBW0K88mSt6uwaPb+V+RUFz0deBDv4naI6QUrUkD1+PU+6uikrkt
OcFIcC4Wvj+bQkLnKtckNUA49nxDtSwaWVJxtU+0No9ACtjd/1VmaxZY7lY9CGrG
ABbJ+z2FkZkGuA1bGRzum8dwoaKqJllQ15f6Me0GEyaP7rtEMtj96Ku6yN3bhe4x
toCpGTFKJ2jG0lo2tyvXFp+APfjmagzQEaAvQTyOmBiCz4Rvz+/SM/9+BGkLX4HP
49uW2UAaEeQ8O++Cf1BcukVb3rfN3VlIwikXwXHnOePWvtJIkZmNCsBe8toHAMSX
NjE7NYVUIblWwOKq2kpIvGj2BxvJKnRrm4RpXEU2KKGxCFZIARAFXH330Rzjx/nJ
wnEborJh/qKrOpaoNTjQ4+FXLaVe4eNP581YP7Nn1+Ysdn+2IH40DpZUaS+tUiC+
WvQVoKT/g5KOLTHjw9Yb4ZHvckrw7SRhowGotymxWwk4BIjDSwOkQ3snBhzehMU0
qQ06DRLBIQpSV0J9YORp95B6yRZbVTld3aase4WvyifPAZZOqXcUhvRB84cggO5G
1qHzfJY4lMJCXe4G+ItO2se36Q5tenilO3PdOe8iij+aoEqV29gO+z7mqoQuHZ0Q
rhp/byONWUcta96CGZt7BiHLN2bIBYEGDcRHZJhh0pE1SMjyotbrsCnRSYLEWq0I
wuV60HS6ul+LklZyPBYrbls5MLjUF105+kV9V2V6p7Ve8GUcHH8gnWQYAGDJAf4j
ywG4WI2Svr4o+WvL8G/eZEzbshBCAyJWf5n9W8qfm91a3UhNtRZFEDO/TCsWOMV8
4dn49Co4ofTBift0JlxOFg3UpO1kVycqar3v8EpRWeJTxAw+uyQOA6ePYvWUxIOQ
V4+lkAAGYsY/s1c2+G98rlc0FjQC3VfUMVcOLvVtHfspyo+d6Z40l8KLColu+4QK
I7RDRpUu98z8WDbbNB/LCSZ+tYMuIqDykFZAWGnuSPYRtadJ44AQ3B30Uv5gQ+/Y
ZwrGhkTFtjIAI0E14SOWsFtB3V/jYz1NVDobeD1Klyiqy67RuL2B3w2PkWNC8AiZ
WLa/QKnwwd27PaOLlcEtJpIQ9FB1FypI6WcAPxTtHmnPUtnuAgoTxvE3g99IOEPu
W+BT49yjpVVfONlucgxdNcsYrz1VSh5kxzVTmXFCulrkHkuKyKqf4/1NPm0blkQ2
dQRySxufeQ0Wsu+mcS1uujzXU5aTFf0n79OdifBqyvTKghFCrWOpMjPxmi9Ebv8/
moHFaOOhoUvCf5CeHDCQbdiXVys8XdJ7Jw4/RtUjNCYGY2VwSaw+Hzte0m3g02Na
r9cj4aO5LZ0sT2+paMDoYh5XX8uYwyBEeoVE1oeDB3Jq0mWHhLRq/2gwKy5g7NMW
iqdzQDSQJ0m7javh0Tl++xV8I7YGqyrS1LkvTNMHqlZFzUwqXkJ4qBWYjxWmYdMV
x2MNKNvLvQrgxUnYnwv/Jmp4IdlYZMGspBo+e0Sr/5TmQN/IM7BI6Fi70n/Hy8rT
tmprV9zj3K+A8n2cgwIAvAstxkSUCWDyFS2ataczh23KauTJE+zPkPZ4KRau+/sf
32JIuAMvGh3MAFZrACKdJnUo8hd7QsB6cNDX0nO+GulfBDCzzh1iB4cthEpKW3hr
eMNveNJeRU6le2oe39qJZ5rP1Lc6tupL05ZP+sQ2JLTcJOzvqUIGJksgu1v9PUUr
gX51GpjEn21oD4w1JZq0izswwYIfelduylMiTWs6+zMUvU+VnLh9DHxujEoELG8C
e8YCwzhkdDBmOUMH/XYmMmLmi9PxPjdQcIJN6w7lVSNNKhXJ3+W8Ls2qXHVjyJVr
br24m1nhduZEED2N8W4O2yk1QZQcIv/dna1s3+yAbeJKgpvGmFkETuqrX+sl071n
Bk27JOyJ251H8OVI5Wq9HEi+/zCZXRmwB5tzgHzgvATbzqqBlt4lW0WHHER7r9HO
Qg3eWgiSv3zcJvyCKbbVPksPamSVDahg7QwqyOEdHqx3EA6aesI5e3r9lf98iLpm
yFGqC+kZagaRY+nahDTdTLZNvnGtnzDJLz12U6h8LknyLz81jZT43gAlWTsWViVo
vQ5X6KDM0+A35XM0KK/wWxkbiGxTUwo30yr/xr8mVsgzAcpSK38SQuAIOJrOqNv+
Y9EAf8rjxiEQBklWREcNvrP2tazWZM0A67mGu2Il2eEOVK/xioeEPce9RRazQdyk
72YROUYwcb2t9prqYWu2hlCp9JEWIGwn4cVsNl3SaLIOA7qJC87FWxlMooL0YQxM
G/3gPUVFNNKn5pNzAjs6htbWhmlL+PuBTTbxagRNPXy8Ovwea/hViRNH+tfQLXLa
7HhZBCkUkYxpGEVICBmZ61W+kRyBSO1gV+wwDIeQMI7tKH6u0B945Fgzt/p7B73j
p7oC/qJdYs5m26BOr8R3rXwNVOFP59Y/Mgsbpt5JDeJP5WYHD/8tg4J2oq6Qpe7S
m8IIZWSJDBIIDUeNrBq31MQs6tuy1faW8E8858IiZCsKlabvcLc7i/2UNHp5Q1cr
zZZZOJigfnyt/64vtsun+o8vRuaBXgk9j3Na3UQLnGxrWw+jGgeCGgf53QAXecpw
QE88eUIPC2k0Z+2ySVhwh5GP+AN3AMC/kdN0d0RN92bjdbozEJB0yymkxlzwbRc3
ToVdxWvDUBH2HTmdTBNur29TkqG3qBDc8eB3VO++fx+nqxwK13Sft6pUL66ttb6o
osXUx4jQ5EJPNO4z2+owvU6Mu9I6mMLncc3yKoVlzrrjEFC8c4OIbeP0lqnB2sRO
C+BYoPvMnYcBmxcc1Ik9+r0we3JrRJnim17Sj9cBstuDJhdUiMFfFym3qqc0gNIn
WsZXx04rlC6hAsvwFtjYXuvT+kd0THrpkFBWAi/MUKH6eTiUd5rLKQH36UluKE0c
/3tx849hD1ITSjeBow5IIcOPJdikCPNksXgttompKxxFJ0RRsI+5Rrdsa9fRqMy7
COatiPolJUrFWkQ35PDTOFQzF451XQmIJ7deOtmLqt8MRJJUuX8CeC5V0W7K4ZtN
VVdoDmYRRH5vFB4XcrW2tU9c3IL+/Uq6pLQ9kr4/3+3/g8mBDhHTb4ndyltWxWcQ
6vbbpN3/DPA1yvleRGP0acII0MxvE/r4oTI7pnnm6N58NPKpd3GTvsPzFNwsxFR1
6dBd/Rf1HfGg6eSynoc5acQPHfXC6QLNELWfZXh0NbI9mMDdYH6VPd5xdfvIP20x
eTV4ipnHzfKQQxzwTgzZE11kA+IuKkxhoWQGk3Wx8sb/uD3UnYbyyTdE42wRHAV9
LJryWHR33h1yvBJlV0n2A08Ta7Q0n1/fKSGycKzpztIwKhjoQ+1Q1FO2KWXcCBzc
AhAR4iTOPlus1yvq4ghrw8DXaWErNPu7mR9AQXlthcX4R+1oRBSrUcPzVIrOZDN7
RaeSJzfwuC9LX3xTrrFwDOUQKlnEsYLHa5FqpvENeIoU4Sa7g38Zc0ZC7vWSun99
RqXbCN1q0U/1GF0geGoKor5bIiTLC8ZIqM7rAZr54OAJjo4bIBdtyYCLs3OcsF9Y
tF/ALREy3Otmh2STBOfVJPIovn6gDGEwJYcJjAk5lNK0rWQy6rjwvWVQtIKPrIpM
Msmg8+DkzYQU6rZ/RQB5KMOozlUliL6x1yCB/6DUwhUN5cmNey+rKzT22i0jTZB+
MjnsdwtxqlTEkcmxjmsxCkB1iuplcy3tBoJWPKI3YeIHuy+ruMRX2jwWmdnanqj3
deSfxi+3/2ls5SgWOKvEz/YwVS3Lp8sYvPogHkKWdrwnPtLxE3D+o8eHECz3k1SB
m0pd+xp2sVpbc56wi3eg9nGxBjJu6NbxS39jsHmhBHBLX3GEc6L2ugP5kkL3Hy0f
qoFcRPYyLqtmDuKQu1KJncm+tIMW36onLhYMqdBfXyf8gsq4RLg2+BpbrWEThYs+
ZD41ei5WrPmAfpTBlWG7CNLYCQm9EJgmneWR+USpE5YbR6bmRZL1/U8M7ADn6sKI
AJMz40IGI3ebfTW/2sW2qi9i5iA5KqxgQeVrmAYiMPsCBsSRjd38/HWzevqnos04
ZW/wbwjqkH/1GoWOdzKcChDMkHuJP/h/yvQSKQnRxClRjvQEQOS+2HH80ExZGSxZ
9rtW2z250xhahJPEtlbixMW9st9oLHOc0LZnPI2VT5gOKKQ96x6T6Q437K0xCzLo
t2T7gp6uksSH/8fNMXNakaWEwFAJdNO/V7OJtFmtlsbvh01LD8yOFWjakrgs6zqz
QaqJWE3K7iqIIA5EmDjbYzIv+YsYsFirNn2N94YLDSrDElxgBqwtxtlLK1RnZnxw
I4VHq5GzuqxfuTpmBMvUttzuq6y57BPVmOIJ5qRWl4C8l7HR10qjrthpCEXzAsTl
gde+aTHOGBL9dffJvj/v5GiEAcdmpE+wpSw8m4pCWp8H/toVPZ6BucvDPuHlLx1i
yWWCn86YKKQbtHUUa8JMLM/j7DjyM8OiW1A/r+GOOFlQgCZk8mJW9m9DwZZYoS2s
YwW8gIpReKu+nGhSFc/6cismOPUDqVJfHfkkDHDpiDLTE+zNvrKKcPsdwjdCLN0P
9VBnBo1o7y2D6lrZiN187uz+BRaygwm9J8mBzF4rsNK+8gEymV60BrCF+IomeNS6
QMlxHZCjO3bdw/rbBMk0rb6gGxkKdvSJ/TMQaCmTbSfgsBOxZlTK3jYzRUZ3fowd
KWSG+m6Er+NopVvnFOkdkytUPPSfnPARuEly9KDSNs1Jc6ZqD8cabrDf2R6rut8h
XOaedy5vL0mDPq4oRXG/v9jlNAiXIu6+xWOojRkv6s1TQrLHZiLJ69LKyNNfXu9C
3udEBGxMaeFtj5ZxDP03X0AKiKHcHoF+JiGXIKfyEfYH5YCLG208ycJf4q873CtV
xPA8sQNHB0IA2ypzFllXRuM65gFFMn+mzvHbtH6UPN0iPP3ywAHeoW3uwx05XGSg
/E3y7/8ZKgIGUn5U+DmkeoH4sn7+j8TX5OwC8NEuGr1Lzv82HNSaNWlmCkfH4jVB
3fJTPWBWOyS+xcS52BeS1GgY3xhSjYxaXXsHuDQT01uLhU+d5ywTdAVdc1JGil05
QLPvvaOPTri9HOzOdAxzVqF+a1BELU2MN5URDqnVgxz/gVMYwfkA3aQSPWcz38y9
nJjJim23wR7Vpaqf2dvgdqcrB7ZvA8uSVSrineSsMVRXz+gWovEfpa70LrHMeWSL
3WifZ9utQQZHUO2tnFoUdJnnC95f6a4W9nVmaTpS6O+YjNPAKxlbeLVxu4P/PTL1
/JFLIw6XQzrlcBEPqXTp5YY8rRvbkeT7/Z1ZgCztxwJjisTBNHY/K1GWqGDu07m0
aQLg6yje7EMfRPAfWHUXMiQFpSqhq1m/eCVcfUSbg87EwdXXfnGXexIe0o6T1Dwv
z4CxhDqbS9hMXEgEbj64No535kRYu/St2scEnuiCW+FlpTYPdl59eYMSommTEC+1
Dm/XCVLI7s3dSknEs+C9uiDYKAzUJw3XiwzP+mHN34fTiUOUPV+7XxuGtaYukIPV
nqK+2Qhlm+iRlLQnoU194956+1cHMDBssaafsohBHFEs4lI2RzYRhk1GxiK/UWR+
jN/Hv9dFjDKwwxNXVZzGADhbZrHmQ9BrCROXIgg+T0VsKzlViM+/hQOU59yD/xsx
+E/dsGKzF3Pg1MVoOXU+8r89/Pxjzmfmjt7MKj1osuvw38yPo4mfrQhU3uHF9Ldf
IxvrSh/ToQGyYv1kqTuQN+EPAoBMFUEfqLaGUA8E1q1MCeHoMQppj3LCwPbA0xg/
+lDEdNVXDAc0BqCQt82ursqu79XdrzVfRytdYaq7x+PhgPn/lIDpbjTP7Ly492Eb
/r3i5pACkQKe32uxBvPCV8HspLaVtnBH8uUG0Rc9Yy9QM7VZtsEVOStInMkDfp2r
FlMumpv/ctidctLEv4801L/m2Aqi+4SeahKlL4bjGZW6RkwLCvqYklARjUOYeQzy
H8IIavllOTMry5+uJIZjjFomlA88S9JyxzB4YswS2+akkBCD0uLJGsIzTVt34JwA
0YX1RiceRBcXwSvHk6DsIxQ6EkD37/SfQ2JYnUZ8P4vhwR9Mq9BLls+OMoXHIqMr
r6cKqr94aXKgXyinUsQHYSbnXQhsgV+sAR+/HPppifrjV+DPg2d8wXClduwOYhPi
ovo+fREtnw2fvSj1C7IGR/S1n6N8OIgOHBs7ww6jcK6pIIeqU14rggrar9m83xgk
vy7zgA2/by4akx9Qr9Vj5jAstctla12lxw4rLlydWrSj+246/Yzu2z6YYBK4Zvp9
CdAq/HF9fScQ2hRyxs2vks5jY++KwAzPXKT5vgs/YJdvKoZmegAUyVroS7LDb20/
TRTgxsgPl0QUk1jXTFNnEKS4fanA37a2IvKmEQAD08Y+N65GiOMdWRw5mNHaHH2E
Ssi/PRkUx/D/ZUDowJX3czIjyIfFkzGYjBxxKHkIFj1luQLwWnL4Y2aDciNXkZeb
grHYNPYo4/jaVsmhtEYPJUxYFsT5G/9Tx8XE6V39erkzzkRUc4NTXV1UY42KIisI
MBWx5ScUEI9JcuSbwhIW49FdGvdceoxpNAMYbbZsQmLHrKfLj/5bsJY1I6PNcQJk
+Fk5JLBIypnjP/QTXZS4WERnZSwsCK4sucLIwrEdc+elxDc8FhwdqNiDnKKayq4X
9mjt8YtSkCRF5i7ba5Dfimiec1cSU93v3BS051KgNXzk/IRUphB+b9qIaRD+VLMo
fLynNZ/j9a9hTlrWhCKlRr+fJEGiQOJp28qmfDndsWvmyIUwCMbwp/IDBWMRK02n
G2O8tK/QKGLoDZfJvYsO7BJschJ6kMV0yxadOmHWmgiXc31BmjPdbjJsN7OYz3g/
Hu49Q30h8hRODmg1Tagt7JW3F6ipL589zXr+/yyAQWs5lyDOKFnNFXK5oTEUC8dM
ZJy1zG0nDSeetKckoraK5IUeV7soM01VqihO2WBPeHsqsyCug4Jh9oVXRuLHTY17
dtjK84HHCvpER9R5Y0UpVuVKFaZ3qvOYdv5c0iLah7lNH0pUscjdXX+qqzholyYA
kgImsp7h0954YfdxP0nfM04p+Qujxb////UxF9SLJuNRSFLm+UcETrhV6ydBOm6R
Is6sodVOxKibOEHaXMu8SLzMNbcvGlsdRT9FvdQg4rXlwxBd/NkbwYqjOmGWch3f
LZI///LlpLdFT9yGFcHj2gf9MjqmacgUoDVeJOu2FvGytWpUID44yWbqp+YQpIP+
yhjGTeFvhAuwTwYvDR0QOyv9hRQOIrTpSQS3rCEbe/WCgiyyePQr0s+TMmwViIc4
7uF/7+fsLSRslOTL/dbozR+FIfAaCFwP0G1OatYIP81KnMcvglGTOeY0Ik3RBWKk
sgAcs6oIQcA0lojoP2nIiPCbGg6tfqwLToaurAbdOieZ1wI1DCOC22Qa+3WLvgjB
MBy5PRvBq7efBBzlJh1WihMXAZbQ8sfz/eFXNAdJZ1HWGSYyNw/8WVR3ANnfc2G5
ZbgRGlBEJCQOOL8kTkm4z09IZRnSpiDtP71adlMk/2dbb+iPqox3A9kCsmS/T2kC
gZW0L3pxvm1o/N9wyEuGia7N8sVFI+r8uFRIu7Ul9ODB62W6cu6XipZLkcnCXbGa
oxMSWYidOhIRJx8RP2gdsRTkNz4kQ5BSLqtl6fjYhyJFEGxapOpD7ENo6UtzMGwV
X8CcFylQHa0ziBLOR0f4alSSs/bXJZkjG4KxYhLS1Zu/QgIl3yHiWgmm+SAXnjX4
CtufF9YTaoFGxKPF3+fgEyYZeJQK9hegXLV40Was083cRUg35iPlhlYeNVZr+gPE
VBQPChSwlHw6HRDYDrG95H0otDYJzWFoZ2yvu48GY472fAYeXM6r7dQwabetHGh7
oP2I5Td1RswU/nJDqgDHhQceAUTvnGuCjlZWtsWgkxXHA8R2Ic3ofz6FzEEkD8hL
FOwRGZfOn6OJTpRbkq5jJNquLTp2C6yDHu6TuTcgSXBPajhOILOnWRe7Y5NdVXd4
xtewpKA7QLqIKtDjy8Hi5UwHmiSEQBg+NoPyE3MPz5k31jwZ9jYpH/Y15eYvtN6L
Vdf92akB/6X9emrBuRWhKOwa3NRY9qW1vN2Fbtcm3pPjBzKY+9VGMyblpzz1o8nN
YpbpoT3iXy43CE4xmkO4q6OUcPsKz5FfJPwCcBeeCP92O4/S2a8garMPGpxQPVH8
XSCYkW4TL/B03NM5amUiw1cjoqOPi4KuxyuUOch3bKPPGx3HkG63dpIjTNU01ihH
mE5Rz6+fqjkMkslS5ak+NUTye5Tg45WqJgQun5xEId4xYLVt0OOgBOG72YleBCHz
/gQ2J/EhC9onFC40V8veZDzsGPTtqahcZpfhSTIBbOjAFP4aGIiwpSX7svYYHi+s
ES2bXBFWHvVjgEbhu/EYRhUy39NiawDe6Z7JzuaWviauwQ5W7k6MW3XO06uHraGz
vIWxTCeunFlA5sHe/P8BLAh0ZLX8UkrJbWw5HWQEx9cvj0xpFMQ6JGsli9HOs0ei
qom+UnkK/PQaojM+W2Q60uqLKlfwakM+qhpyxU44dcBdmB3iEbZaeZX87sbGj8G4
sokG9CqOgBjdeECkucYMbjWb0bo9CsmleE3ecBQAaZoaGkMdH8LDqJDW4QNceiLC
VfDhSF8touGLVly04I5Nxtovga929aeAMnNYSwdHJPa6GPU40fj1sbuVPWewXty2
XtkeAVwq5TrcCzwcX1Gb33Tigby7bFOW2NQtV59Bq1tPQk520HHChc9mXEhF7NBr
gq7S6FUqTV96G7Yr+hCNItMDIdUOf5SvtXdd4PBYtKBhD1ZQTJ82mvZv70671w4f
rduRXCYXRZf0vN4QANi+W+08BbbU1Fark0TQ+yf4FPH/+XC/t+SF4jGeo6MMaroO
sMAHcxCNrhuG68TrGZmgexx6UxGpeU7QHL2EUFYjQZ1TbItcrW50lWVVgYgckWFR
K7+JNlzmxl+5g1valQRS/zLX2Tn96GGyQ3H9CcIhQNdpoZYR3mWXn67B1YjTO4FK
dEmZYBoZxOK9XDxFWe6qNnj+lzp0PPmgJ4orRIbuLeniz0ryFDH6vhpIYvIfvtvF
R0iUSdsLptv4Z7bW67JLW3bYSyms2HdQY6QapBI4qHQteZoM0H55j0Y/ijDpnJ26
DSBuXZGxB3FUH8ElmMCmO6S08QviXVCk68psZVK4hu/C+FM3jON443d4/bLwij46
DQXa0gxXeeKX7kF9uCzaUPtaZHc6ZomPMfd7dKI8OdXBalnYSrvq1RyxKPuMJu9X
9IlSwX1AQvplzK9p7Qk6i6KqGQSfc2G8s1HmXspET/DxeqDGeAV294sej2LH2PPz
ssC5CQIS1GX6yqIUk54qrDqw5RMMItIpHa2/KeTKHWYC50A+gkDiA/ZsO5LDcRpO
5SdCJ9TKlYO1es6N8B8Y0ZS+2xDYH5jeiAeyHXAKX3khD+E6gycCBxKuohU0MO95
KCtovwih+NaJ9cKqH9RL/39+Eui0vj/UI2/sfV63Znm1bN4m3pclWMml4KyXOytx
4igxBda6UTdjBZquTdWS/npesj+NV77M4ApBuhaJ5xUtC9iBSazEyappUdNt7CFX
JfDiNB+nOWBKJrqHdsGAADhxy+ssho4YLj+5j8BHNsAizmkRVQuuS8SpSt8PXAR1
Mt1FEBdn4uokwIyZpfappR7gZv2WvAA7H3sQbww8Kt842HEtfKb7hT/fWBv0dTZ3
I4uM2mFYcWzBt5p+frnc9bx1y80kTLUnK+dJW2ly/ejqQJWdhDS+g0fxH2yNoUxO
Fs0uJFOfkUm6EEHeg3wqkg80meLOWRU5JF4MgewFUtY2iq6X5zEKmUtDb7KTBueR
pKRnMPzF00p8kMbHWL8SNj2ODZRZ9aphgBa4qLvVDa8/NwIpyz9C//9W/uLSZY6i
iCYOWogWZx04adpC+2cmH7b3I4YkIA9iq6x7Av3CiWtDh6MQS6Q03DfdXEtuY/UG
bEh+ZixXRXr7jghpECfQy2HFD2QZVjlXqS4fFgvPM6nmL1HXXUPHkGagJoEf9KPH
R/sCLc/FyxnnrkKqvDTjjnN52WYTjVVBDNfkPm05ZxzdfAAXHxmyBEA0yRa9sSj6
2BxZiRS8hJQfc20gFeDQYbs93yb3OGFnc3u4SkbDOh71zXJ7vVgp8ojZHXfutuZ6
qqC21KSxbyR9wWmNhPdjzAJv5R6knav5B8oWxXrIZ9s82FSOQ1WGlToqzdGsAg/0
PMAMPW/mxhaRNQY228xDKbHiUKCYOgrfdqtfUjKPe53mAqKIA+zQBN9D+fK0YN2I
y/E1W1oAkfYOMCzeYrMhcpLeVNB43CAJTnkcKG2Spk2S/gPhgjNB3vJieij146Yv
rKQqPuzBS4Uldso3MYcHannOUM34R5NjX7TxBsY4IxaNSJ3mAvQhPS9K/kYuT9GX
LdIRDAQ8QVRY5w7LipXZ78LwHtyD7kKpMqmXaJJ4gZSCoQbJeUJ/wYsFG90xngAU
It2nrmSdNcgjbp75Ytnc4JZCpJThTa0hAIh9CVlbXKCV9lyeXbXwBoKy+nDu8oat
Gi8L3CroRSbg4OvwpQ0GQzlLF+xXfAfxspeVzn3pwyuzh37FWAf2Nr9qGW25XW7u
VeUSO5KeuTifyt7C+ax0mN4f730sUeY8gX/feffNRZK8s2non2nmDZBPaD6UO35d
5EETTpwYvBIREKYjzx9ZPrLSygO+/3nFZ2vSJMKP99flcyyRIS+5k6MLZtxssmsk
32owodOLGXXsV5OhWhhndJXJhuy7tZKxHRm07cJ6g8YIQgihfO3kwBGms/+wt/s2
54/ik5M+w3uUGXnM4U2eonh7DwXNrFsef7P7//rV8WTFzBpwFPETNxSPXuaujpMN
63bjjKHh2/hqi7iUmIlUB2W5Py1bpYMYktSmLxspMzxI/yhxJpCV6AAzefmMoqsg
HB+bZ9XiAoeG9OZRF+9io/yOdhesQ9JRVf/TQghUUvu5KVl94mQlTLNnnPuMPBNK
xcBZd+SDNF+BInwNVNsdhKKLQXNxuXjSsCTvIcqZ/ET5UIlc8DQruJmERh3g7uzl
v1TD+onQUnoIinY8f1iCvIscuyUka4RJtHVBtYHp0X67CJQkaXHMuLhTgFOqqSXt
g36IVXLt49oS6wAFt6k/zn00sek7jD9OOz7tNgKgKpMEskfN8+SjWpDGupYodXla
Kel4cQqrihdTN3rsvE5RCVPDg/lUEc9QBEtl4DzWknXZbHcuGS6oQQ6NHr+V09Ol
/lBSCjWYcOtoB7MUg1Hf9lU0NZqZ+KEjkENgkCP55clBgL6LtbdIGriiFoTnDgTh
M4s/N3e65J/AUXRK8OuFmQnR3F55SJKaKkwSr0mAmarjzyEF5KyimC0d6osfCDIp
+v0mBDEjjuAiP33cWbbMWf21/5AMSvsN5s6eP9gLL0MG+Z4Ua3dKQsAzcCpFYNFS
sST8hSRcFgcOlLsNmmOtQrxGXHbszwV7scdIG8iDN4RYvRHJDnoirAmdpQ7om4Pg
tJFLBz1Gdo/S6JW99ElaeuMqajhKIwwZM6d++PEsF5cj8HS5i0ELHKqvlBWLS6Ni
55xpJd4pjifML39OHstCvWYCJlL9LVHybSwkjzT6b4M0erdeYc32+AXTBwbbMLJI
tA/CbhS0l8Lb86CqnjvrV5VsHlWIvFEUat6hyG1aWeWYpPKDuOc0yQputTYyDQ+J
vp4GaSaZxnXkppRVSsADhsWCPiShqWdeBNoR0bj8FEII5YZx969gyJODAUQW9key
6NS/U8bcPoSDFN3O8iy5o3O2bIp4Mm0xUHp2J3/xwWq+TinNbc8E/zI/ktRhAdFY
7R7khhi3pMco9BP3Nb7EGEZQS1LI0jF7hBW+eGcX/ypfiW8jTJ1Yj0rS2KGKleA0
6zrRYLc1PvlbEv2yPwk6F3v1A0Y+9wvnsViOzCp7yMKasmBUxQkkXcnmzaIxKgKn
dmH1sy/8YrQCXOvO2yArKtlsSZ71FVsuYBr+JoYg5TOAaBUBovV5OLaCKuzidAdA
+KikmLWklfq2GwjE5vcCKZAfMuNRRyfEGvbgaBYu6tYsGvvVlwdpcwQLPyjduVBu
coZsNmFwaWZ7JKL65eKRxK+yhkIpHZ4c7rRvEMtpIQyLd1p0i0nYRH8Zx9aK7HKg
u2U8iqLgIDJm4/fpIh7YhU5TE/wkzxB0rsjENz5UZI+O658IMLCZL/jtFui4WMRi
I2EumueOfdvtOiLiL2qur1+mdb0B2k6NDrLh9HtiU0BnyvJbNetQPCEUeaMzuON+
NzcdzsRqrrSPCYldOIZfx91z0NVK3p4NGyaFtFOhRTzTR5ymgWGyORhXlrOMTsoH
39y2sZnodS15VCdIIFfXryP7U7ExOR2E15DR9BYUDCd+HGoPHVpppcvnhxiuxlO8
304SdlGFbi4/S7BoRh27UtgklrkRoaSHUEGMje07HpyTRAxvkfWB0OZ8IZjYc/Yt
t2hEeqyMSVqrz/QXQ1oC8hPm6w3Ge0w7rlf2/LVbTIDo4kAN9LRnohz8mEzGvGQl
mT/IaTelbXamrl76/yeCYHvO3nyetCrgMCj2nfCIuAAtR+f4BiS7M2QBTfaBUI5Y
Mi+0FbixPTMjUyQeNfxGYmq+JAosr0BTKY1sqwkAxMP+xNaC2SblgRI2cyd7mxRy
natgdUVP9rL7WEHLHbmCkgj5TzMHXomAK+Mukk9JHjU5amoEtqXOzbMIwd993209
pbI06o+7aSxrfoaYp4s7NCyMXT0cQDLUiTDlELlQ4noHICvnqdsT0jgBVyWgEvT1
nZ4JjnGTn0xXqqHHs5dblAuLCLN0A/LBHPrej1pm5ah+WlQG61TvJSIm0u37jaRA
EjYWzUFwVMGyUwWAyIDXknLl/EwfK/uB54vDQG4B+FtuicLAls4P9ifDM80pqgyt
WsFLiqYRN0FxP7yYV7RzIbmMSrDy/IuKNRK0OR0U/LnvDr4/+fPHoFvofH8LYo2I
EnJ1svQ8uHAry+dWz8VVGnkSal9/CSnjMHH6x8QHQIdkBUq14efzxwd/VH5s48Cx
9lnF1CjomW8SeIg1rA6FjCF8VS6dhNUmNdXe9tMJg0FUnju3+rW85Ra7N4bXAH2Y
TSMs5I8m85+RkbSl9rcwtxpGg5bYIGn1RoMcPKkqpj3LbF/NPwWs3M7LQ3S2+x+x
puuPKU2Wk630pV4OMesMFXwWX6HIka/0jretDMHJAy1y7a+zLe4ZH/5FCuQ4Kd+W
HJ2SMPRXNvKroBkySOqL19meU1AJo+Ivtl0HJH2wnQ7o+zTw+jRkktj6Cv3BER1q
2KVQ47c5D9mxVsRLad5uTXlenopOmuVdalZU5c+/iJkFCRA7V3bnslypdweUdjSq
0dnP3chMdfXT8aShb+tzl5dguhoiA1zfrU9WFdhQWtiYEwwHVfE7pna2D7QHSlHL
SH4UR6F2ch8jAFvnVY+gdxjcnikoYRbLpAhxrxLQF4mkXPKhSS4jq/K72QKMPArN
+bVOGYWgqcenGdtYC8yUeWhWuExbxm5XYB2X7NiDM/UeS6vbUdH20we/fEBCcRSf
7J2S9NmKilGl7ucD8Ged8ZKHzMHQyoIsx0tHKuOP1T+a8ubvCrULTKjWPkUsRv0y
Dkp4DeTQlNpHhGTzRtARc33Y03nihAmYr4/MXDx/7aqjpMXYnSupyAxch5oDqa7x
oOrYyMMpxobm0Bre6wTuNHktas1MW3LolgBDr47Gtu1pv8CMWoRrvwhmtrVzMxhV
UzS/9AxxGo1wf3mepgH03NWRVGUXl1cx8PYNtNPtEYqArMx8yYOaToQnqv9PEmyy
FyZnf35FUc3cob/QcTkZRJBPeuYNA1xIE5yk6/M13K2Ens7C5tdarBL/VeMT/SL1
HIDG3D1q2s+8MMRqNELuc74DTbum/HrsAyS+Eap81sGIWj66sj1ovSRtt74sjVR0
VpVg+3bxEtxykL07BqFWW0dVVmewcKk4Fl8bcXde1IH7nD/tTG9nKIJ3kX1u11eV
UG928wMrCLO4+j87c3JpU51TFluKapZ2MfetyRcqtmej0ndmqNVgoa8sEsk2y0Um
a1o8+RXnlbuonRFwSUiJ5SC59z1EERBmkGX2Od8HTYzmqKFEw5q5LC1SU+6B0OhZ
DgpwFIrpqs5xxjbURcsWAh3+YjM4L3GD4i0omyXx8cEjGkuCO3QzgjW1lCK38RJU
u7cXx6xyyPj4iEA/QNjz4I8m4MXvcwUUqLpFRV8+oOb/8Ad7+YV+HOyWYED0PYWh
0jWOm565DkAJU1u07kPnQ0hl/+td9A4kBJsHvmM9EgOrztDOQTgSLwSFHXiL0dNg
lsGRPSPcjf5Uu7m7C6oWMLe9qZ4QdBvx1zBaR9alyTBu5bNPi3ZqtkBrEzA9wt4D
OVOc1Weh5Y7LSsRts5SL+E1zCcuZez64STeDAC85dhZDeqlc2h1oGDgxPHW/i2SV
l2ruOAl7/803TnGn1aADfHepsoJjTDBe0Xa0ygPJsA7xdlV0k+olsO152j7pDTnL
qnDIcU91U+W6dHt0A0QSx118RoJV77xg1mXDPoGlqTi28VMjpHxS7smtQr4Fvd3A
0fBYtLyKdNer208CpdlzOskFFUfZF+0pBFVlrOESN4JgtMiDzKJwxtxZSHmg65fR
p8KltiMBDIJNIT6rJQqyRZuc370KvMaHgD8CkowCaVMrrkPQri11BxyXr1JuYsSf
W4KmO5RxVaVKblmyEu5TI5LYAyLrTVsvU0XdU5U1FMxRxN8tCRu7CAW0v7ubJrsJ
rDs/zuKg5yu/PgQOLcTppSqG/mcNAKexMv79jxMPkK9hB6XguxjZ26D37yIQmrTK
Hq661UWWk3vwt7NTZ6F7XGCpeIGx0nco83vSNw/Us+yq+rnM8XcZi5XK6o0/bHwQ
Ez0VAbXERoyu5/niWmLqUf8B14PH7JuJzDd8HMFguJ3b5sO+3bEc7UIF8TSEZ5KU
SddTMNRpQzauHp0AXyzFw8JhvWYp+jgVEay/TE5gq24QHfqJtUGrr72fzteeSxYF
0sPibrcKzeg0edBMSWNILVwvAf/5aYh8GOHX6mDu165A+c76VGIu3Vw4wrKeh1Z/
+gnUZ5ccknwnGNwCxEb9VzbEJCzKFmdwXEeFIj5QgE4AAzRL6vhfrRl94UTFzMhB
MS05/wdysVeGvBRB1RSNjkLr0KZzw0XCB3HQvjusO2zEk5jFdmoeAvniMXtR02EN
KjQWqnoVZqVAjvn6/mguwAbyTBQAcDuPAeu9ypZoE9FVaWBVumNdl+rSjehtpt2J
aq9JRuB1BHHd2tu5BDMdV2LVgPFeLScn4I3T0S4UVenfWcDjGedbJK6sCEECuvyr
jc3WVIVYX7N1oU75/eQRyHWaluApStTTDA+ms6UMBTzXRCc5Ch30tuQ91Y85o9M+
pcgIxXgcPGSWvkKhqMTtMprlaav8tshTXIaCLrVC4uJMXKzsaOm9/AEp5x/WwjPk
079e+9Rnm0jG1a/n67aHaixZ1teQCrRhPQVOxEsYSqazzlosaw/n/AmfR2/R0fA/
l4sCQP5HJDvK1D0AI8KEnf6hYHzmzvKuHnLqtOowkacOM5KM16JPB5v1OtV1V9Ob
12Bi8W5N/+L3JAi0Tf7mGngeaS9UIDjcdMKKMs/z+9IEb6PQKLWlb98f3QoXSEDx
jZs1SGNhb0p0ahjO7Czqsz8unRReWTjWVChfimZxjfhPkv67ncJBMW56B7rcLeqN
vEwuFzPWVLs6/+IVJQcDHUY9ZSDxUAdIXXdKFexYLX+dYDq/RjxXwqHFY22q0Yu8
fez8kYi1G/LBcc+83T4DdxFYp8vtXYQQLpREk44eNEWuQvScF+gp+CtHSZfMgRpR
EnsnmuN1/VJii20DbCiat+Y9XXibTe1ckHo96iOOPeex0U3S/JpZWW2D6/Y4I47U
C+SVjah8k+qlLYKVp7OFTVhhAchyiKkbyGf8tUT8qpFwhEw5ahVmw0Z4MsIHpA/u
TJLXwBMsGgsXj1fdPI6iOdFrKRZst6TywyOAwnxSwbEky22YYT0VC4jTpNeqsfqG
m0SdC+EiVNeC0QMiwRgnMRPaCgziYj1nlD0BSLF0nERnvNuUk4lvAa3F6zRIXTDr
XyRII4wX2kNGo71l6J1QfGhktjGlZsld4gWbEu95lnrhlxlukatLlWMp6KqiUq+b
VYic1+Ez7+M08SfIBJ/uBVlgKwX3LQQ7E0WlSpODhRjxIyzzlvqquyIvoYivGU7i
wtavtvsO0oM29XtS1pXFHMSjB4deSQf5TJwGh4ju26V1Ugu/3H1h9Rgo6YjYLaKn
IF7H43/gazwA6yo5pB4W/2RUei9XR65SoXFtkcETxJnjnE3GecH0wC/hI1gnMA5o
yrBg10AKqD/mSXQqAjyTy46bKlOX5qOcBEOitdTrOJ4N87NrEY5Hyx9NGapJfWCC
W39dxAAG2MA1A8v29qAtHC+ll00yI8S+0kxpFxvWIcKEtLXWQahcKT2IH+x2DTXd
0ur6W/FHLb8+qaJjj2HN9fer6V0/NQIH/fsKF8ruCAlgOEpu9HnJJZJLd7ZQMkti
Fn57U1snfkusNl+C+jNZguc8e3xGmDxFuB9VvrSVdSSEyMeV2A9S9cVoAaqIbJ5o
WcHNsPU44fHmruE5LBJb2nbE09YkJXrJWh7tO9C0tlL/VDPmNrnW3bM/d8X22sUO
krjcOl6KCnnBe+4IcBOXkfwzhGvjeGcQb5J7oqy+UHfZAxuRedGzcaFHtT9AIuz6
tIo/lyWSxoYuRMBeTuZQU+qJDWLPskuTBleKk4F5h2d3uIC6sx84pC9hV/b7LvGm
tXm6U7eKKbgHDOhYm8g+uP5a2GU/cvMHyP42aGP9oz7cA1gLWgXZXYXd1Pq/o/yC
KfnKuHfYHFWaL2BUC0U+v4PZd5yP1N074ltTbEU+73/GST8OGM6urAFPGuyd1vEP
FXPB4gtuQ7sROX8TuzO7uVjukTEgwFMlHd8/9fiqC1rN2+XJoGPfo6ySdLFdVrTQ
SMJStWcWInUw486Y819BRC1h7lv8fUvP7BoC6BF1U5NHxxj0ahYPey+pv3m5g4K6
3At2ILxDm1SsPd/1e72Bun1yg6ht6wxqU+mv1x2m87mGmBLzAA/g1+WpfgVMhtBt
fjSpo1KdV51KwpESdK4mr6iKrKG90yOn7SfBlcJGz5kG3EBsYXF+4fIXkZNNyy9U
eyUeZpSk9LFzCkXWqkXaEDNiyQvGFriU5VEqc0Yekue+JiG3Wwe8Ud0H+pK+mmpf
xbE73U9svYoV226vcBZklaytjrveyPXZWg2PGsIHVvFT9e8+Mo9nI3Z3uMvI5HAq
gOQVHW6dL+hcSFoU6qntMce7vccEquHOExDWJav/kV+98cVfDFXjLEg4yIPBJECM
VZNacVNKehZrMA/audQ9Bc5nzxEid30ozfZfz53PJEDZEgu0WkD9cRHBlf+GEp2a
1AO8YxhOdSArIeJUxstAz7iTqkdwaIw7UI+fw+jFU6Ft2JeNP6KiGgbjxsc6dJk6
3uuZ+TjJ2SVi1ArDZ/rQQE8gFv1y/KkGcfY31iCN0ymU9QI7vXaO+GnD5Ms3DDua
jvdWIvNzueNLDhMNy6GQuCwo/23sqeKJCuBmYfc9mhyDCaZ68o2CSZRzsvVd2u4o
gqKUYHrdDJzB+6wCe2xKihon7jVKyI0wTT1AINPsZbGs2qrb6BBjqM7sdG3N7Jzy
oPFWGl8eq2vjhSaF7mpVJZq1VAenhHaWvZU4fDgDYi3z71unHoEEv7mnKVxROSKk
B+cKaZLj01I/ZKFE7WNRIz+gF5A7xNcPcDoY5rbaydglen2yeQyqD5cMswKcq2EL
8owhgEJ9bTyI0CZE9re1C6yZBERsDwDQCcoMrZBeMQrvHQ2RA6rR6kHfWYmJxdr5
1AwWqeCkLd0rYW22I4M0bXKapwujaNsxC4QpWJno5kQLbMhlHR/UPwp5ROxwVLBm
u9SbyivFKPlNXOOHfpPY0ESIyUTJzObgW74+8vdTb4AbmAkcaN1fa1IyjhHi+pqE
sV/kkh6PakaEQZ88SCoPlbNXIRQY213bF0NLdTYtKNif/9MWXf8YAYYD/sDSeygL
pHD+baQtQevu5R4gfRVAPAqTqmeaShR//JSdkCZ8tCG/xwG9DLBf5fz6YezJ/gCt
tznw5D3Qm3BII4DSW05/gnU7RpyeAozXSu5c3tpq/U/Z3eaC7GiKl/ExPzXMYqG9
S8d4NT7d3pqICAgFK91Q/rI8ZGEOSC8a/vrM54HisDhrQrvIgjFNhLmHYBG6orwJ
k1iKo0K+Z7UUKdH4u/wZ2Hg14UR9wSOwA1H85Mso7Cxr437Rsmy27kU1xlUkBIXx
qe5CDYbTiczCRp3qlEfdNKTsPe6ScnIDI6idRn/Ktuj8A+j4qcDjO2LTczFUTbVM
QQUPnf7uCI0NgWza9e5SfXIoVX0Eau2yExRNft/AtiMQMxFU95tWIIddn6K2MHHw
UNN5bGFbKZ4kLfXvTz/w9bRRY0RVXWQPlPUZG//2uoOPjrF6MI8d5HNXLV8/Nasz
R/V10Q7cawvlEVUBNNwVW6PAaDgBOKXzYrS5ixRphyUVc0iDUHYJ/S/mD++psvK1
UFx3bH1LVBLGyDZMoJA4QRyTsBhNqzPiAbGrKJcnmQAYDISD+GFaOQJgoeWafu5G
I78s9XtgsIfSk4xsWSLk4EGDEbz/KNqHxZ8b1bJOEwu31YrQqzFDdQLlXbHwkEXV
ZzeJewUEeLclH453Kf/kpsKxN/yxqm/yfOhwU8ePgwTC0uplPuSCQ6fqeAsiz9dx
QQ/JnPfTz8Ws6XrjDzNEqhh1Gc5S7tNY/iHnr7fMPacWp/nvz52JewIv4wybQX43
oyTxF+md7SvQiLLt7Z7CP6BtcPbs9aoLLw50CGfAuSx2gXD4tKhxJ+qxnKoVtzol
iT/nY5MFCk6Gl8ojOUoVgxJy8/n0/mcnF44Y81I++IFHpOBlDsvbO0/ieLDgFYuW
InCvlGHiYetBl7Rt+TtopTCLWMIBYBt4liEIr9XQ2bsWsBrdYABpVamw1MgBvy13
eBW5rZbqpZzu2ShDyarqyj+YRC/RkHUj9qsBkyF2kr1jurHr/HDJK8kvZ0jRi5Sp
b3wKvKYkoO+tKo8hlmWXtDgkG3FWkPc2LWehhnneYLuHoFhKf5vrOy4OCvQsUdKi
NSiSRGDxrdXTmC07ph6F06E3A1hHtgHWe2d8Pt6fpWPT2QM4iuGWcXzL+X3bHGkq
nqulp/g2DrDhQcn3Fea20EAta6CvN+sA3R6V0htRO4KBueGgvGQIkSJnoKATDwcE
28/w5egMcZmfApOy5U8YTh+pUtDET01YebUWr9O54f213sxkGFrFDYRy4yRrJ0dg
3aPceiBP4WslByXiD518fMAG6eBGAWPGtEcm/LALRsStTEGS18DtPgnNAyT4cJ+T
A+nwmQRTGWGAf4uO7QgOHJOB5YWAkMYBbDktH8//LjFKcH1A4kjFiULNG3RorV9I
VvsGGyM4eBxMj0I8PXW7r/MSYZw1iHHyDrgHPd5ALZaJUDX7dxr/NNdPYV5n830J
nKhLQOe9Aib04Z4hJdMTY0xdX13pTlqZZ/KyCfj6eaBIY9jo1Xi2xEjqlkzCpEJo
r+VOa2v7sD9iqOYQ3ljrYQtXKc8khQj2/JneZtnwnyuTvKU+xmdJZ/hxJyBL6lyG
co8+WD2pQ80JmWmqL4uzKgOPqUZCRm2eabwHCfFj1AArD5qnpR4dq52IAdrC/Rhu
zOqIzlZchVaFP4dA8VVdK63cydSqA+JQBl2W5h5QGxd+DQE4/C/yzrPsFnNL8J0L
MK6yRfzMv6AqFIbtapsJ1davQizRFNGVWFzJxVaqWIM8evSw0OP5H9tBRfGC7PGY
IsWHKIpMdOa08YtBy8K8O8MVkm1fdRm/DJW+oQyhmZ24iNAalRrW/pcVqMod0EM/
+D2L1mqUWmhH7JSfzd7zrTVfF1TUxMUwDkOTbqEfkLN0PNOqQhmX9+0P26xjwN0e
HrWcFfmpqfSLCF4h2IlGsIJ2ciovfhb4h7Wylssi0xdysyXBvHd/abCWCCQfux2Y
vem04hL4bWZTXv5QLblzhzMz0ybaOHLWy5o3reBq8A36hXkZItHRT7CLKcAcn+FM
d/AO0PNeE5FY5KhBULDhAY8Zrj0G90blZtd3vyB2xpJIQyvbqrwbgF3wYelrjQtZ
7/bm2a4mx+ZPt2YZalAqsuaz+y73dHRof/Bd8d0EDg14c94zZtRZ4ojRTwNhSFPj
4RyUxEq91jOgr07gqx6gVCa3O7N4wRctUAw87NF9nSk9F8qIVpL+S5wvbG3fEX9p
gRud4/9jrPUeOFQGv2UV8OQUOOIUiQiN1yac6G9bBxnevTUopf9pZgSxofDsngOk
RsZXA+gDnl9b0RI6NncYzR1Q31pFSudOJuW5JIMHN2kEhGHr9WfLqbxS/eNINYWM
3vGbjgW401H/YCGJGZ8ryn1EDQmAEDcyfkoglhAxE7Kr5BVaJreddIk4jjpA9Xnn
M1N3snwQuM2FgIv/0qCj5RPlLpqz0hwXLfMVS2wTMzJ8LZs80ftY6fofGOO6+0tt
79wtyMAOKeoVnIf2lR+G8J3+hdpNEE28oDwctTQnMVn10h4rYbkp7yLKkne6xwQU
YoTUxwsjXnfaAVt3VFeAyLI3qHLXwFtgf4StvEcvESm6LBHcEw2UJV4d6c2X7B0f
shYMnLRV8BRFCt8jojLR7qhOkX7QjEhArCUxb5WV28aZUoip+RGRav4DWyKtiKuz
v4Yo8tG1jHWB1NRk5b8gUCwI3Am9t7eDZH8gwyiV0BsEgFdVwHjnGYGEduFynImA
cXc/R53oKv/ilzCqstwMhibmxPELfQXzZYzkY02pC6iHhXzV1xtKgE3GLHjh/dxT
gXGevvE7Y2CRYTmIusEYJHKAHfNNCgRDE6OYTWqxypAuikJq0ZRdDZjVZ/moywAe
uJlZKgcBUK1VBjDO0BYa0bPL+vAmia5WDfBkN5wyRVmC9zpK6x4ES2vcMZOSiVwB
8fNQPnE91gygwDZo88DAH+DjNPSWmNa/8yhcbOSkVjvFMMtJqwvlVBr/2uZ7WFlr
pK0/2hIgFLPRdlbVipVv5D6niLzbp46OVmCMbPgjAx+sIqb8UuQ2noHWTiAUkt4h
6v1UiwdabMfhdHZ9P/MdLafmJvhLYHZRck3nbS9iaF/FDVMeEP9NlOqQStyRjRNh
ffIFeLCEdXXt+tYnpVF/pZ3o/7OIz181LDS25x8OKDCb0UrJ2iZ7Xe3PehwdjirJ
I5TQl+Sm+MF3JITNgJgV9hAr8XvWhYz/eDUzx+HlF/CMsFJZKb8/KxuV+NxhU3Gb
m7+lt+jy823OvepF8m4vDhP+A7mGxchIWcLKu2deT5TGVWd+T8noD+18pWwXECm5
tvK2/8OCIZ/9gLBsKFV2xZFbeEf3QYnFNXBRL1Q5+4ArdyXuUojv7XT/58b/1IgX
OBT9+9K/xXS5/D/1fnYaVvK0MjGlfNdjGgQ7F6m/S9wFBZ3JVCsfhXB6zPEW7bJa
BC2o7NgGLLbjA9cXDaZsK9GMKaUx48uEkUGxaNTOECrC7F8Hg/icF57L/t+G1MYt
xyLQFLMtBiW7d9VWndTYPts9gdpFotwy8Lwpd5CGiyaB1TsfwaSTu13dsEWoW0GP
GRb+htnGLx71EYouJfE7qUpcl9DuUW4Ry+fI85spUWFHXqkQzPSe40QPeRuRgNv2
KFORnszwTuBV0vHJ6MPpzIp7EOQ7mkWEvjhySM6aIs+oUA4icoNEqxNCQSFTxwLO
IrWEOUy/au48ggXoULvfY7BV4mEE2nESozwqBruGHe9x7NtL/7zlUSjd51CuqhOz
hHfdtLr7rFfreflWNJsWxQBsrzkHB7e8cAdISEZguVses/8EEFMxqukcKgHgYGre
2rj2W0XWiB6jsetF1wt2/aEWeFJtRsmOpraWtCIH1AY/wY0iYHRMxJS9yUNBUYSC
M3a+nHPVdyxWb+Yi9gI7lgYwNZbMn+4S6coOvnasovRbOqeEdw1Ye/p5SFQkZsLD
MCiG+PGdPv8QNTIHCaaX/tuw5T9eE8wkTfCBYhPeh9m9Q/m8By+Rxszg7E8iR0Mi
HvF1TS7goVJ2mMFmbDeJJ0KglFAhKUKdXmE9TN6U2vJwktDja91w6GPhJXtqSvfW
ZC2uZjzmuJp/dGiqRjrKvMU0Z8ljRH9DOIkmKIqEgl3Y4XgVrVCHiEMe+81ufYIB
e9BlNTcftJd1DEr9Zx4LE+YjjLjyORCIugOVdtq4UTrocmzon4UbrbxImUJp1CEB
FoHuhTm2FkTaVvr01zjyLc9EGtOXqfyQ8097E5xdcXe9mFPkEnu037uoWik4BiFZ
WKHX/XAkpVyh7innKvNW3KnKONGBze2PmTQTBPvXcUgmXaV//7mjjf2Yiixg6BoC
Ybi37fXtnwji7uH2M07N6yMej/bOdndiQwXzgSuzCmdYzPeA4+nIK3HWTwELOPtE
2HhOAIOPACMoULo58u5y6swxGg0MTGmbA0K0PnxcOhbaRdFM8k0lfrlZgzIdAVBO
L6mijjgmdIWRgl1FaB2WQStViGWam3zs+y92nvim//iMab6mCKCp/SAN1wOydnXf
HM+t68G56Wkg293aOoutLmrZ23iejiFAAviTw6JowwSURmii9XFUyUPzVlW2mll3
aThrom8gYd169arE4JSOBXU9i7gnaJ6c/vFyalikAE1g+cKR2an6oWTpAJ2tlGoI
OfoR79PfyLZG8b60MNkW7JVcibydQ2Ps8SRaWLr5zmbHUAqn73aoWeGBlKaKZeW/
SpxG8fLFeNdzqWOn6lJGy5pf3cblquEAHArav5PnzE93z2dPUJBtOh2LUrxVmHbg
bTQfWnpZ36oHRiXudpFcxrS4zr4Wct4K3j5en9Pb8Hv3D7LY+dHs6wOVqXekkSoN
rnn2Ct7h0U8v0/EkL2RD9KP9T+9Kl6t9UEdVbGxEKYFs7LxLdJBl6qf1aT2JSXbv
QgEtNn1U4vdI6lezsdADvaW18kCDNLg6zXMyHCma9kj3mrlyI8nFmXX3zGwvaPY0
eKBtSUxLwyxkuxNPYVKd76QCaecZocO1dNlw7/cY1OpBlGc8i0TpEw+Oq5RQkibt
YeZs5ZgmRJRzCzJnAEKqRRd1lviokCmnaoMvZCiVf3+girUAR5mhmkCqsaFxeY7v
xULfRJ/LP6Q20f88lim9bqxZr9vhG1QYBol7XnnWKx4+RTfw6fJhAFDbUW6D5PKx
19SoTQnQ65CJYx1qrkc+2h2TZ7zI2UjrJDQvg8ZI5JmmsJBYm36M190Y9Da3u11Z
VXc+OagKt1STK4K77OWCpIetzDYnz++x/UWxyOtOTGANHSddJyMW+MR3dbPtR8FE
6xHYPrAQ/KP0/1p7ecB0CHqbn2pwecBH91KtTAlS8DYPmgKs7/5KhTOX6Yp20T8t
H75kqdTWAMKrVIh+/ZdyEedyIvZoqXJ/QiF7gqjfi4AkypCUC5HhzsOqBQfWsLSN
z5dZVbke77L1IR0pd3IziwDyPJ92hnHqxKyawn0uujfWjPm4wpelXbAvDmGpnjgd
kEdFakQSduEVmnsF+AZi3Rdd6p88YqYPBKfoa9WO59/IQMsdQRYvTQ8Xnzj8mZmM
D6aSsQ+HSy8U8VhcmP0ghgDWjnIeow6ccxXX1vOXAcN2JgzMOWRMPHI7qPPa9PS/
VIh8MT16Ir97IyI3HAtJsNMMx+DFEozEZEe3p0CSMa9gGjGBXXL4ecp0xsWROVUU
0yOSmxYfnvv3nkL4bJPiBslT6/WOHJxIeI3URa9T2NP4EB6c3hPp7iv0X5OoIcpg
FTlkJsy1BbK63qi7GktDiaVKo0FfY74WCP2GTY/QYNjNT0YMZV3RDCDgKCj/UdRZ
lzNgw72Fibcfzr3MHSRagrYk/XH4fARjI32F5oxPaVFbo2Y5oQNtR5mjWppUoND7
ljzHaiPNH1DhpeEJh3ByU3BLi6KFK2fYvDHEcLDokD6fBtjxOkGGWiIqB1egba/k
Vx+j2tJnR4EMC/HRCFpERr+RA7+THaNXIcgwZyIKgLvk2iBi+J8JisViUreLhCWX
B33M1JSooASZJF4w+DGPT0FToBQIGMZNpynuNsIhd0D5TDLO+hrncwF4axPgyWud
1faHXxp/vPGZGCKG/3WVVv5jB8rA6HPOoIZ6YqIqm4bs/wx8PY2vJvUvhxEPPfRd
tL40XTR2Zr1XMgHaWr+2mJoY+e0GSVE+0w/Zt7Jz4e+sUhzDVpD1ff9sfUx58mhP
fqC17Nqp5GJKeFK6T/HFyLRdUhndQMnpCJXGcOoaU3t6AZsqGLFac8rDt5MWWGDv
Bmz8Py47eW0yEyvray+vUzXh1DTBrPujkIc2oh/263ahyRcwcpGfBd6RmI2ntM92
fxlDDqUaPko8WZr5zjNRUCxFTtcfL63gWjYCJClc3Lsdqqa28Va2f6HAsTeJ8nKj
YyWAD3dCOFZ37RCSbGAHGVAFuKwEev3bP6hi0EQ9Iw9olueLUTI1D6AKKzGkc2oO
7GaqQvZTWWNsb5kxkZl5RdtepyD3hvd0avaQtWpUXintX9dHU7uDcqkKtU96KvO8
x3tdfdYuXMzDn3haaOINlGKCbYCkRt65y3Me6P/y3APLTEkDGu+M1f0qaik2SD0u
12doiP8yxkvAns9RzY2MKFmMS8vPYuCVwMAdD9iW652qOXk/1pfgrbNeFd44Ul6y
6Eq/wsSbhwM12Y3GEOPDZW/2mIMH7GtLoLWjzNb5hpik8PM+8BBetzQtw9lV4yBB
XFzXoGSKaKExSH7WhfmD503gxuNfy+Is6BMs5r2tH1SE6X18M3DSZ8aOK4+v3u4V
MfNCQUifb+Ft15QwYHPQTIz9JmkWIrc1FwQ8UfKPTVrV2VU723jkHK5tuNTyYjDR
iNkjl3+SVdyqQ69ds7qSxWwzJkXPGdj9R/1bQrGobYCtv/i8tIpE9G5j5IjH+3la
frbJmcdumjm15iN4jzQgXSq8jeES0JNo05mos9E6hh4TcUCwykl50BPTNTqNMRIi
FLnCrRVjySHMx2iJPfjclYidRcTDj49F/AD5tp/mJcqo/xCvqWGsNlRL66Q6W82T
s2FZFJl/mdEHISafjWI/j14CK3W/6SSci+NrF7z36Fy01q/Ph889I7Rd//qYKIRj
oejI23nQHwF/kuYfkojNnkTE2MXxKp7LUh3HmycHZkfBPkQlr+eK2T4Z5w1iI1mj
mwbXnrFZokS611BWoVOHo49W0fjoDgTIbBkfsYXkxbQov0i6NpqHiBPFuWwTAKaP
ofO2obd7JIZXN79pxQd2u2G/6XWnY39YVxSg8S6Vz8oAqAygm3Z6fCgNpKl7Torn
CTz9+46YloINjC7Jb7/7NwivrFs8GaY92lOVjP7wMyCgqfgu1g8kt5vlDFN204ay
dAE0V/rBkv28nTs8dUGuvu2dIP8RtKBOcrA39qJNGPwFQD3OuiddvPkpNZwR7iEZ
KBOkj0vCVdN0eVCZF1ooeoWlBNILg/MX0N89gG1cxUhr7mRwdXiXJ8rInL23+dq5
/MPH6hAqc19crlzkfeGIguUKJKGg6N/G3TMYb4yhifU37kjlIHMZanj8vdIjqgzy
qBUUKfkZi0+hVAOry+MlmyNNCn9QuMfJ9POUJwEOoYiTaLug7tGOhprnpU4fwLdN
dS7w4vbMjO5xKeaQl+s8siSka+BBbDegq5wGC/kmFmCGqScPPoehyS0FZZ9qf5sK
DGROuxj7TlqPwv652SBJj+04bfPVHvOLBZVpWhfGw4DxoVuIsbSBOuspg0hlhrTu
Xa4zc8PBcUnXJD8o2PBOvqWiObod+KfjXi0VMIXkYrKxR0f3ODUFlsO10dgLnBTd
cvVzvwIKVHTzLl/wRJYyCz4XhmqMcVdwlsJJAldI2NWhJhqaC455lXQ4hcU/KzqM
IM/AiU+3oAsZxAX25OmoGhGkZTe8ZoLE4P484JvvMeXzGXELTMgsEvF1y7eLvwa1
/z8z7klAPAt6Cm9cHOg+x84OL7tKjgxpH2W9b9xGYeEZWvoXrosDxRRR105XEt28
UyeLp4saeoUQGBj5FuPzemSgIQ2VQs8rPNkyIcXSjObH6EoQrdWmyJcZIKxer0Oc
myngkfZ8ljCvPAnRZcLxlB+ObzLE2D2pz14pDD3YPS3fOZ72zUHrh9YNzOBzDbu3
hRoFxqR1l6fdIFl4BXIGt2ab+o3R0DjrAuqIWX+hyTIQca2mbXfz9TRJejvTPxow
EZ3SH5vREaOIrj+bf7G1WLKpEUVEnTeTsVlX6qot9BYzQ/bFIFr3Tm9WqMXSEdDB
aZl735MjIWUA8QBSMickQG+NtZAa1Ay09hv4SvEd/xdtcbeJzCxaty2s9WvEexHa
Jf2MX9JekJHU4yEghuSo0HbugX4VW8YwnthPnEVXlHWogVM6soOwjvP+JifpKGZo
A08j0hyzi2y+BJwT5c/nBiv6DeNhGPypv0XGuMZPVszjGhMKX4AvD6sCGE8hZPpx
oHyu0JSVxwnUfRWuI0M2K5QQRQJWGKIBqiDZIzgba8jScLM9Z6lewjWVMDWNaOCl
p14Nril12jVxnhvvnJ0EqGrv8xNK29pfzYh9xXEt/JwdTuiEqE65vwPk5SBMvzXz
v4L3FsBgigQ71IezvnGp3F/AsrVTfgcV64fKKlhrjkU/6PqcEe4hOnjkWX+XUU1T
sdWSNzqr801G4+ARbiaBFJyfo0c2jeXuKV9j5pMV52ltqqAT04W7HLdA3NTXwFSn
mn+Y7dbv4/HVJdIl156x2MtZMQglPyhqw2zQGaPrtts5hU6AyX4KvYjAWJ7Bbf+W
uu+zul859Pz7sptjHoKTocf2kVt3wkmge4oeRVNAPAjHzF1QtP837v7bIq3pPAJR
LxzUuTGyExIC5xdkphtA1J7qgmHfhTxB2no9NH34oeHraWPa72IcSwvHcy9seFuD
T7E8CID7J33NQxxX1YsirGW6VmwC5GR32zsrIkM9pMGIFSmPZFCj6NOyRm5FXurh
qb1hW/tVrRkKarD+9BGHxByfP+EOLob7d3x4f2cRGwTeDMZO9zwyNhfD/wkCo979
wjVG2fFgkXLFZSbwGBJNI9bRHvMIKLUtrrkfyjYyVZ/dDiI9Ql2zAmaPHKIIPbTb
6Z4AqxdUoT/Ui463z+aqtwuQi+xnOJPv9mnX1U4kIlPKF/WHxu+HkKrDVJl8j16W
2VFx3FMuoaIprioDWIEPQk3+2mBEzMSQc/Bi4iA9U2bxz60MIwCOntlg0rkpB6Gv
NG8mugpyKWdL0/brGCtPjX+bQhHIyEuhE7u3KWrAD/Y//dEwMsfqeDYpjDb2rz/8
EoI0Y/4umzUgOiQRxfsDsHbsR2wYmcniWtM0+WsH/JSuKFnFFY+9MppBbyO+ERaR
uFcTViv8MyRMHLZb+RjA2k508zqPEcE4rlGcJFu1yhGXtfJES/SkdyWl5Rr8+Rao
mnGZayJklvZeBm5BaLavZbeTxP5tARz8bTfvbA39ROgr9yUKuCjdcF79EmCu3iyn
TpCoGDcIM4M2Q81MpkSR4idVGLmjrDoKUNn5yYHh6ideCGEVZ9D/R3PnVK8N2ql4
/3EpTCkSKDGdHw6k58YdyE8Vg2/ksJrjyOgz3TypanUN72OW+dL2K6pv//2bhm17
LfGG3oTR8U1oF9gJVQVrjN4GnQax3N6ViHhUqlo8GnUWnkRaeNK7ibpo+bygw1Ca
lp8LTsRVePrTSv4oyo5dcNnaTlsLMYaF0ToCmI+Smv6M7cAINBj+rrPSwMn1YURT
G2snAvndaOyrXVMB8Q7Mm86Xx1eStQu7TIH1Lxkk+HKiQkb62Byjkz0+s+X1w/Jx
0fjyRPVjQSF4C+ECu52N4LJkBhuSdX7SoYjvkm8g5aKKwFtK9v+lgciIGzu4frCQ
NxdeadzVguohNvqbP/l9ev1rtx+KAhqnWLjqq0XYW/+1D0SBVwGtoX4gHmkQECwL
8+fSQDLR+kRsijpZZzNfa93haaYseGpYbUGtnFvlr45ukr2YanOsOgXEtu9nTXLl
966wzKi3rog5aIIkwgig0gvP9Oq5BMdcAVWkkaXjejJtTMS2PNjW7jodITo8in/J
cVP+xbdRH2btD+qeSec6c/TBg71FDhnxxKHPfgjkVPZpmhLO7VdcibkppFZTTk0o
rogALnKjfrrefU4w5nrPe14If+qiiAnpKVAC0ibI0V+GSwBS8R26C+hj+1+fwxNz
s7tU8q4Ixi0tYKDfIOioq9nXyDBBHOcLu+ehzbnA92uJuSArfGLDjLBRhy4H0kp9
5+kJoE2lmGyh/VaszmLVSgXVbQ4YlHilrguNPHahDhOmkNmn7OmNwBr1r30mfQQJ
9U6ByJeG0zEZKfQ2PFP1WWgduYvxceRhyYE70VERXaIJvB+exwDyUVW3H/vVSo2u
7zH70gUJYuI4MvL4Q3UJBQEf3FXrmmvXL2/js71X7zFCIAeomcwePQCT2THFat/7
vgoB3VNjMz8vf404v5SDkmjA+s1IqDas248EhL0IRDb6BFMD30iH0Ap0n4tBTjzf
hpTDoUOIkSuI1CpWs/eW0u14QkAhVZSeZnBkhfX20CRA56wjiR5RSNqlh/SH0P17
4x4ym8Os1xo/1wxJ5pcTblM4zX6uCM2EUJ0NVJKbf97+Ib5A7ApRA0QwhuBVmntf
QurYLStI6Q8hqkjFWBZV6Y14Hb+hc53W1wQHUaS0HhfzL6WkEQibxzrZ2S6bwKgk
pbjptmj2CUV9wOBpox/2zM3K8tOyLlLv+ExeS/nzYXQmvBLzzEXEUIe+oQtGosg+
sqQD8U5G0OJJ4plYmgQcrNzbYuKWHhuhQdKLiIt/T9YFjzqe5nQ+Zxi8kc3tCQrK
35fex76mVJDsGwqVf9E34IsRvxrbrn+xfLM+J/6TScgsRzTfFHNbEozsi6R+r1lX
xr5/Y/PAX72TXf6mtD4nlk6PeJgBrrhSMZGh+wHZ5Tqkx6RO5tPxTLNYfYnfnAnn
mwzR2BOUotRSOYXJvycx1JMv6DzdJgOErlIA3rAfaaRidA931EMeGTnDelAL3gT2
uSKqaDDENKrP9ENGDmA3pvEOodZSwudIhWiD9cHltoSQLVXUP0pvsgYt6ajGI5dD
bduM3sA6B/A6MJlDjO1XaBqV3wvORsZe3AGcdrOhbDKZdL8nU72FEI86HE9mV3oB
j4MfX7Uz6Yz32DfcECyEONZiEHrUGbCgu5zH8PdqiJnmh4kmzPCZUsfXyfFvlwMy
zKFaX4B/+GAlXSEWs4ipJqQCbNX7CAUMDeeDNGjsxrKmn3SKoUUNOgfj63fUCW+t
ozL8PU+pgN/k0RuMTwkB50mJgznoRUoX+l0YkZ4KCj/ipKIMmvlF+CQacOdrPQTl
3t1Ej5dxcQFg8/S1DKfvC06SkjCJaVfzQ0QipmKLWIPQbcqGRM0OldUorg4AM94W
FO/bvHwbIRCeGTK5PczZhcijtolcDbD+EyighZ6sEeyUuOcBuhq5gaLyTReCyQf3
v8y/DHDfNofl+/uCCNAgWFf/sKcVsHnxoIphS7X/bv+EfWb67Gd8hH/bGQQ3DvT5
oepgcMwsdVInaPJNsaoetbLGDwOb3j42hy/k//QNTgppQQMmahMTLJ7u96d+tECg
Ib1rM4+YcZRyuqANQ/ZcKSA0fKIERyUbXnc6mOnxkzsiOceC8N3CCf68E36WqJ2C
hZLS3AG9NVwzZFvxXDUlfUm0KOgPB5J7jWk5p8vmdGu+jAI5g0JRVm6H60zlDxd3
L5oRlsYLtsHQ3Uys3oTulrLH5M/eiUnHbbRVRLaQhWQErzQbk5Ml43apb9+ocOfa
83lSqpm+7lhrlRdbqkkjw+ilitjwxb5ggRZ79fJBqCA7Mw4ohQqoiQDFTLFi+LuL
hWtQ3FxisJ7T+4n10AO9Yh/0HTgcOtQmpGTeyVfMsXZjs4/e1ocau4tQu4RRuPiD
WLEwANsy04c3G7yDUfw26k5Sbxi1462igg2sPoyywzA85t1NDCy/4NuQ+/XOn08j
XycJd3v8SR59r1P5mG253voulPqZPIOMot1/RujeZPKUg7bNOX8fbb02wWod/3hl
kTqTUscypbqasLT9Bb/ZEuiSXTC2q+X+xV7SDwWR1e4tU/xQvhkhExsZzjsmG42m
M2Ojx+uMS2L6wiBI54hnN8vdG7qJyAdq2dhnn9dX9Xcb36jW4odYR7mhuRr+aqB/
q2IDSCNjC99ahAnx3mrFO0jRBglsAL7jZ6LkmXj3cx7Yjdh0moKXxLy7Xj41lQTB
J8KhXNAIiUlthHjM9sVSmbRCGGElzrJkmEr6uhZIr7FozLUkPgLQCDAC2Rbr1qHw
ZyFWtdvGDoAH/YYDS7ccTlEXMqLBpAOj5PMKoZufc+s3jmAqRrToWH84kDhT5Cs0
Lg34CMxedO4QTxk8ZGziJfAU9k5SleYMN5+cYKgMPMkSmmK5ZKjdm4aWD/4eQYwZ
ofehFO/eZF0TZBRn1NT6SnJzkuDHBd4QyG7eh2+nji5l2Cx2Qu3qz6o/gWw+h1GD
r//XmIBLyoz7fjX/4x4V9Ee739iOi/KvWauqzO+OPPSVuwBXaOAcI2+S3nLMd7Nw
Q8zcmlAHmy6h4bUkoZaM4rzo+MfHK3TCAkMBO9HzMzVzVuEnqwQFqo0+bU2STUJK
C80fijoIDzNcZ2U8s20+Akvd0JGl3rF3vq2+J7TO5cY6TlaYseBkMq/T3wK96pFq
z1Ny3L4ClvRIJCuhHBILWhOfvJLJjC+lR0zirIRaxuYFbAedLcgfI+JDAJiAY+bM
0FiPLrD/xlnBwSnD02M0gJyqdHQk5z63x8kCJETP3iVbL6B0/ktB4sM4KuZS8iDQ
pFG4Hsl9D6xqttN69T6K5XGym4bfffQPqDZXB5cT0GHjJpd2Wxxl8AiKr5PFBfW9
BdIiVIhdmtlqTs4l/0SBJtMrqYK925IsNxNtjbzriatdhzCB8m3DSa6taJeYn9lU
rcgHCP3RkgQBBahScMoruxPXxXGzF5x/6bo7V2pcsfRcizIsifSrWEKDWu1xjU1G
7Jt0sJHyepbWbOnS9Hx0pcFLSZAvHiVZckolMUZu4NN5jXoR24VaFSEcHmAWdUwx
PiNiFcau2eo8WMl5B9gRdr1dU2sExynwzHRFx9LpNRWbXy/WGS+bMVwSyVXeteTJ
58LqxRIlbg1XO4l5cgHBBi9O/fqhiQ5M/nGt8P2zt+vwy3WYYQISI8dWB46j8v4f
JsOQZOgFjz1apJYyOK7koVHO9M4MINu05Cw9CghI/qamH6NEOUNz4BJwFGnRXBif
smuz50DzroI1is2dOiR/GSnVBZAy2fWlACCpjQBQ/nGO4PyIErbS2HBlif2fY3nu
TVm4nQvuR/fJrOkGvaoW0wZA4wkNW8HTzXB2zAVXwB/52cVUZiH0iUeVU5hHvRM8
CPRJsXIgEvA5ADKEaV5RMWfpo3XzoG9K/pU5x/4sSFUfDxvJY6PBM5YutAQ3PunD
D+NgfW2N/IWPQ4yPVnHWQ2R5WLXkiC08sXg6RGdP2M2vTcBy2dJsUC54Ks4BdGY+
yMUdWsG46GzBeL+U1CIQqei7ySiMcZox9p6F/x6W6wQPt0NgURcItzv/TRQXNber
MSqICJK+ziWoJV1MGZfLAfXEe8GlDsh+6hi/w0qzJK6h2jUc64Z4Nvxa7k2m5ft0
kKLKk1z+OB6Z+BQw6GqRCbV7sdK57IKzrmSc25W9Z4ZQ8QrVwe/f88WfWpgbafwt
3IUNx2BAgjN92/PgFdGC6HwfY1IdMvqXfI8bev2T1P0SPGyOAVnfbzBGDyh0hgzN
NY/ECpxgl5PZzjhD+K+TxDYLJ6E3W59zZ+5P3lYrKik2y/oXZ9SlHmye7gqI8j35
bEu3ad/loqsIs/P/xFiJlmmGvF0QoGXxzZXgKpCqA+eh6sPRZmbtO0NjLmQleUZl
UnMt18L2BnEXdDcEOQSOdhRxzZcT7uuMibsDYzy/fiT+ArWC6MC33ndEa1btjnD2
RRfGmoDambZb4+lArKy50GZobdbrLl7Nd2koYSw5fBLOBDR8Ipc61Krz9kIfeTat
0l60eHu9AyKglPvwhFFappN9XU6TQ7G0zKLH7mGL4l6DYWz2oS8hyYr7dyXFVNyf
ygVpNXQ58TCtGDD1pxd9FHbrFd2Pw8sqfrAfblROslOznoVqj2biBZVVgtX4JyRl
wQwQZfIZDAKiECXF+jEjXLpUnyLp42QCMLqUxKbjdXj041ZfGPskMTceDvinKjui
t9kBjenPS+vHTRcQRM7Hy3MVSX6pySFIgLllFVy34KtmJxyWmJeRIS3eM5Xnk59/
QeX3/nyQnaALwe5oYtBhfwBgGNSNna6b6ZfdsRnTeWT82KfMkdbaNT2fsnSiOQds
5cXfHYchkbatNuLoHg7Soo+BeZBHUjS5vgDKSFqAjOXWfWn6mCm8ARtC/gj6xTZL
MmT1OV9oxx8YSx0qru9B8s6W/o2JgKeeKwauVE7937/WwP0KzQba+OYpcpcaArrT
IYWSG8LGEh4pbbzraxJSYp6jS5MWLZLqVzHkdQkmr9J5CiCUyJXASRhSav758eHF
hSoV3cXTv2rjDNY/uT4hWEftX7l8/+EeBi/ILe/Q6UnnKrdGx4Kq+QegJhEjk84h
/8IAGOvz1fYdOa3tkyqA6EiOWPBkbSnWF94w7AFM7dY8iR1aIw6lQyfjaUAGD6KR
yGQgWG+MYyX5c/41h8e/wvxgawJupruxlwmfdfG7pCCZBGlEi8erKGiv1j/4QsXL
jkpfa+NTj6hrJiXiTirIpPIUOylR/9xW1acZ6jtOf9Ela15SYT+shpmJB6FuPQad
WJ37TFpLbHbFzJA4IGiQJ5yFM96hBaPn6rcxJy6c9aQG+HhdG/aboLHyyNp9SmDk
LfN0uoEOiCTT1OJkPNabFjuRltM7dCGxVNdB3TSoW4rlzGKwaSAn/ZtKprJhdXK6
awdWYDWowafcf7kuq9X+/Wc4LdqdgCfNoN1hNtT5dpqeBA8YPc0UPRwjr15FDPqI
sn0Q/HfnuggQfjrxZWbR5wt6lCPbIUdsW1Wy4PombjuG2Gk0xf6r/eGiNp6L/fx/
nIeSENRw5iD8MHkV4tT8SNDIuOI9ckrTOGrmdIB5Ftw8NRHx8x/UvmwlFNZzSTpL
mScyG6WDBUAZgIvC9rNJxAKXiYEHn2AZ6NAygw2I8QK7hIHbQFhHPcqU+pjfqLAb
Pt5A+5YCR4rsD8fmLeof/FC57IwQsG54GNqpPmcPdgv8Qs1n17YVOm11tjFhL9fk
DzTO8aPF55ZmgLVKIVkMCvoj2sjfmiw4LqAKe8OO1ay6EGBs9rcL+LS0YXnFo4KW
HJkEIjSpw62o7SGKd06klOAheqG6aQJz6VpMEKYW5V+vHnTZyzMNdXvPw7K4PQq1
7M6l51bFtD63MlGzh8GjlE9Y+LLyeIMCMayA8NgSbOL+HyirW74YcZrAkW+zEoe6
ciqT5Wj8vLMcyRBw3FD2Daxmnpd5BI1yskl5NErHuC7HZ/RwPJMrCJqNSOkrm6D1
fTlEQ/fhjJUIfSs4DudM4X8p84cNqVUrW6Tj1qZMeh2oupNU+i/VB3PyFqKElN0V
LXn/e1QPt8TGxcXRB8NQEwuA5CrrIB8wGv8yCx+nwMr2U1W/yaTGwb2ZWRRcCu1H
JfWU/1xt7nDk2oft1j3EkvnHAqN1l8nGS8XplUSmLoVAGnLgQiYdbVPa8ALvGTh6
84kBvV7bfdWEVTOXy/jjlOIkc2uecOHF6ufNAN7Uhldw3oTWuklJofmOs5qOXP9B
vKbrPkOXUmi6zMYV1e48CGWUVxbDtcsNCRa+M/N0ewM95NgPfnK1LAwvzF6uMkuQ
z88kWWD8OvLPNZlHgAwKa/qoQeeRrTW+sN9+d75ZVDQ7j/FqE38HK0giPPV1SZTG
JEG7qWoZ2f506X/m08S9kjyF02590d3EewlQa9+BS6IRsxY+pVZVJsaWDpseM3S9
J9x//fZJ8UVx5EvBcajxm2Qs1mvLeqQXO358sn3sH7tUuUxBbInhnT+ykrz33Sjd
5jPAC5T8Df+kCAlzz2ROpEdkU2xP6/d3aIwTITbs8nScZeZ7dVw+YyTzQLPthVij
hBTyJV8aaO8EnYykO+zrcH3FuTZDzHoGQw4U+ECDMrczvxiUnZfYLpClb2UCdB4k
sLjZlaW0zFP/a6nsEmwUb7g0w/81iD0pqs0pMNm6ZEn3R0USBhw02E0YG3a77+Ng
vcPYZ1eTdSsdAoVk8Ir5m9dL356AX9Cp5dMCRR+dT1poi58RHEdjmnXW0BwVufva
FJyb5vrAOjVrCYHUJQqun78tlvfkizBzYrWypHN7tPGeOxepQ/iOZR5igQtK1cuC
p+8GgGbhV0wThZyBGMAH8XnUrTQbxFMsGXtemErrD+bvVFiwToTnzi4+oJ3GGUeI
C3SKYL5PU+bLNEbO5YHXMRn73G7OenFLvMTdLFt0mQDkXZRoXd1P5A0rxGtNgEXe
ke8IoIJGEDC4rjVul9eRPUzwzVcfkqdv9adOUk1M7ioCgy9O6vZoRDiFqOKdCK+X
HAFvAEE1JLGYBFNKe5HOameJwXsePY7rkIbLA7s5554gcUMbOlnQxWpYGQSOiwjk
+7jTLKjpXOaLcvwTviuPnXKQKpUaCrRG6ymmY4VwsE2TQdG47PPoUtoyuorLwFiG
2P/ED3ncZr7sh34ncXMMHa3jzYQrz+2huMSyxe3fwB1kvnT5bHQ7c5Ae7k7t/coN
TbjZPY3g0H9oq46rAUyqNrihpaS17b5yiJd/nQpV8HAHiyXJxtSiDRRZHBva8NG4
adcJdrUO0k+vtImQfe4zNTJKPFm/HSYTT0aT9m/cp8UQ0vHU78EW/Q+6Bjo1hElx
MfocDFs6vVHwgJ8X1NXxwOHYLY3I9SjLnlDxdnASoKbArx8Q/qpl9vvZewug0vJ+
oZQiOCHribfefNzoKY91RybkX5glYHpAuPo7Rgjqe5bFZ/ZbLySeyKbOHMWnzp0J
HcU+RT0ugz0HFWpG+6faAVXW/UIujxYMbv88qzIZvxQTHzLgc7ztC1b5fx8gv1qt
CgxtApgPKeLz5PQAolawMzokeu6hgUPtvdEidX0EpSbbW5Z2yGRmQqHi72a5F3M+
REPpAkakHF/2hdQfS+b/pZt4ntrDCPer0g8A4C4LO5SJFN9VGFsWVivlMwHSvLyr
c3v1OWV7tHJNFrGclb3Ts5xtM4s8dAp+N62ZNhAUvpHOg6sXT3RQx2H/wQURXiAw
1oTxhNBYLfQ5OZxrMMEOjoK61Fksm/u8fmpQC24nqcGwQRzkYfNuQev2ulop95nG
dMN68aOdRzBYeysoTstwvYNLDwFMo30dP8obnlaF+iCgVlloLRBax1UpyGtQ6NRj
XTlkc4wcB3Zx+vbu+GaQRNfd6g6Plx11ykkeid42o0G2CBnaHVn+eEZvliDiUE2O
Y4zIqy21qc3Sk5qU8hRGTHjnY9zgD/Q7dDyVTq/JVJO4yCi+TXoDf3XvH/YjsnxZ
TTYJl9JTG52EdRU0pWLnvnT25Az+H4nHIJen1RcySF/ZHspQevg8gJ/1k9rtLbZ3
yp6fIp0r5zw8sYFsVGn8eRNNX3WrOeOmGHCuSKKAo+T7QQB8hdABAUZxyIB/HFPp
vtW7v+vgVN8t+lh09vJzQOSnXfhq3KiyofKreQTZhw5cseXiTquH0lbh+m1QBrC6
kuXjqnmRgwrRbqB7d6Rg+XQ8dSbnLnn2Q+eLkRU3ISLARJ+FmIG7noVUg021jDGo
z0p8CR28TJ8YUEx9t+rYteyK8tgUjcYTejqJkMxIW+yNSy9Z/WoBtuqsFZ/NMO7w
`pragma protect end_protected
