// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hX4Npj16Ar2VVqTn5vf28DB+NCAmqrVA5GMaRa5QHgQBPFBzmkT0DQn3SxaceWnZ
b6Qo3TyR0ZoMb/1QtOGYmfoTVEP5KkA/8pf/zM6GS5otF5fUHNKvc4DsJD945zHN
uLZYzCQ+1Zh5klnUKj+A10DPchrQERWkBwtQyEr7E6k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43248)
KiDSfDE7TVxazM1zF5KpRBtaAMk0I502Lu36XZ450pmToDpKNf2yKAaKYKVXXqRV
YMTF0yRgNpRjk7KWLkN7+9hJ1VtEwscba6Pemz5JS5jPwpqp9AWeqfU908Z9tYWR
mJ7o3OOtU1jlSfN7CvQdQcH/1QuDkoIqH0kHE6o8cFFAiyLcPHi1hys6tt+KSzwn
g8Qaha74zTV0SoMnNMulsZ/4yzizfNrzfT4jxYPYTMREplmttmDWDM8/FWsjMoOD
mlixccn/eEkDkaaCd7yXpM/YvwFJsTNAUArGesvmldFXWRe/bb2TySEWwpOQ5oGW
2IOd2MROtenXaURrL8n/FiLtvI508RXP1VwvVgL2NsyZKQ4DWCD6ehn1i7zMwXk/
V164YMFTjExGDoLjoQ9l8X/BvtSqQDDdDjBIY3I7A2oskOtMF1fMg5Lv5Phb0KdF
kJiwkOWvNivyRmfchiq/OJPKv8Kl/rhDU+Sq95lYQoyB5777+IWse8ydVR5GZDBG
eUnSEt7CglFA7/nnyIU4zd7eSXLVHRyamk6YK3AJRp8TlNKKQohtE6Z9Do7ZNbuL
U6rr+o9R9pN0i+Ui5/4Ftj8GRaRRhE4ErPvQ6aVI4BelLQkZsGpeSzxDj3rIWLxa
jOMGYBvwV0umt/l+f70zjR7h5ZJfO6Fa/zTorQthwL2O+FmKwkUZIjkA5eOPTycr
D5tQ3Hot0LPdU0/SQN3b+YLPdr1OjAwTzrMuqT4s6A6TeQ5lmmDCTyqxhjOvESdl
kulFHCn7+S35gOU0q3YfAT6NCON/6x3NRbCOSasPU5u5ZD8A0ZRIWf6BeoXxkdFa
t57MmVuVCRP3u4/4LpPjs5Obh/9iuYPxtiHo3vkrxvsN47CFWKLcd/SNIutwTwL1
sTMBGVQLMWTCuxxPQTsrCVk+RtP+58ArUAleH6+LM5UxPV0DZoqja0TK+yq8oA7E
gfGvPRA0yFAbaUfojgXxWzm0OY5nXYsCBAjgDoEu3ZO9/1n1M+a87LPjvBu8KHEe
bCddsox5HCPAgq0Zw473o5AZiPlO1rrXNQpbcCBFH4nW5YVznNAbDwZAU0BxiYdP
BpJG2GSD30hn+QVEwQuxx19OCNAZnacG+BcF4XIhYAXsObFPv9pI+te7J8GfQOdO
8pCHh0nrqyH32QDc7AjMCTA5XEqsHt5nbtpV0nm67HxlWMpikap06XIz1vhb1ZbO
OsS+PIPY1SRvo7UCknPz0LPyd6ICJhJdTzvJyH2RF8VF2y9Rw3KeqZEm6w/SWIvR
b8bRFEceK1KUoBNGg6ro8gMIHEVti4pd+TkhqgPOGHeS8prMfyQUnkQQ/XmF385x
BB14Xdjmv4aiiPz0IhVGfBlpTTX0ROfVl7zJ1HRyjtJEKMdwrfawNU6srTpUR72P
iBM1siFPGkonmn60WU5QP7PKrbi5aS4zMif0yiRZFWoU5t/gA51j3tR9kiT3xbVk
CCxfvM+oht8UZt20JVKGpv7lsvjWU8AbgotIn6LoQ720/cGehGrAQW6YJqIbxhh/
SJ2PNsvVoZsnlqLxOYrrJtbOrbsJmUF8EG4uPfc33O7FzoGSXrvihfmCuBfAjjsR
pb7eVJ9jEaDjhwZUiR3NYIwdnzQHh7wIZjnwDDFoaNl8BX4haAx3XTkkKKEJJiRF
KWsRcCY1i02qXhA1HrU3BySbDIek+SJ7DJeE/QSDkdfzbXADm7JMwz9OEXk+VlQR
/ScHCxo9ig6Enz2C/IPVX4GUeX+S3qEdFVq/rSG4MPptnU1/0E8Xb52gD5988/jn
3Uu5QSrwhj8l+GoKb9MBYn50qHldiQz4pKyL68c914h1dl0d4kGtrMFfURlHAZTF
No3G8YhhoX2dgaBcsmmZ9AR7yvJfcwoviu9eZdrekQuPaL93IP44wlHhLp78zRHX
u3OMfDWKpd3AeE368AvimdxJYp/wrfl8sDXygC0jq9fWYKCpCx1mVDrQAlkQHXxC
9m62ouSxMvxHGimz2LLP89ueljiIshcF+3AGK8dh6KTSt/QZF9fBUyuXI5P/V8VN
VuQPN063Gl+/aSRpdmd9tpYxXDji9M1GWSCMT3KsPFN4puV5P/fPweYtcbZHQet6
/vwiLF0jLzfuKJJYLUy/ocRaWhgmeYqJbV5SOrynBfHJ4NFrwNDjfs9jQf0nHtq6
N/8CfMjeZJfevZktcGhAg6vhr+6o+re7GlFxpwZGTCg4dEDPIWf+7cmBmK1nYNX7
7jHM6EYRsT9HRoRDImt+1B8X1bsXmds94t/KDUtDNv2wAlh6uObnbxg3YKTaHELj
/rgJ+k361BQyXTl3y5ZL1issyahec4Wy4CshXusTHqRKvgdE/0ZYCCNupnT96Ex4
OaV2ikSIdmNA/VWdPph0bt9bhhtaIzz38YXlHH7cEdRc8gKuB401ODbBW3TUdWpj
HHyvzdcyGJDwNvsT5W6soiLK95g7QQnOEzAx1sxaxMcKotCxhroQmxh/Lnuqy3vT
XU/o9vYA/mmXfbXJRvPonT/CKNSLs2dI/eakvHbxkhYCRhzg6KwfcDnR3Dsn3Rdo
5No6BO2K6qGAHMLGTL/CIgGiqGCxBh9HXSyvwTN+cHyunLy4ygOTkjLmbv+ZPI7X
kw48uH8TBS6n/PXEXSkTZ9HzZG7EtLvf0g/lbCpiQxwrtky+TVPyRqMcTJrk1D6q
gHDQ12vp4y4Me7UnOvWX4VkOk18RcY/425OZ4aqLHzeQsv5/jjIqLVjAJHZI2rUR
c8hXR9a+b70IJtLsz7QemzVVyv4OI8bMYkoEHRBNNRBDmwUbZoLp/gNCdCCfIdry
a2zX37EM71cVWcHhAZlCYQ7o+CdWxdIZBN86SnkURUWHS81JGE5Tvqti0UVmkn9V
HeIU72GNd1mILBDfAOMzn/y6sSu9krmL1hsN4gsAmcRRhdSH2WHSTzxakdEfJ9mu
LeXyLdE46U396CC6wQKdGubXhfV3i335hOiZsr9l6GLyXAp50JW/+nTSVKuXE6JT
W2GvUPsjOsweJJwnzrLDI59X5/WG3FE5Y0iKbFND6VMD8NA+WLDyorEpubzKlMKa
XJ2rEX5z3+MWreyBYwz6NOwqOq8yQwWDHubMOYEn31oI1gCMtx70nccZVMFiaElV
Dsfhtni0aIufxgitRk7Oc42b8m4NmQpi4CtYIw6gK+iF751SGiqpYj3Ab8MVRTF5
/D2rjwrSbinDIAPKEWM/1/LNnvSZMuNGEJM9M+BcVmlNYykhIx88U8Egnj/+Qzk3
gDPqw5m7bjnhzpsxvgABu907npUgj/orjiKrULoLKKZtPE0Lbq0+FIPi5CKRt7WR
EEeYst7SXBGVuP/QrtMklO1dLWbVXozvmLkvuC6uYbRaZ2RYdfkHEdutQupXIZ4E
saiWsEBhXTyK3FCyb/OJ8z+mi4hUcRzb2PrrK62g3c8kkRe13pQDrzuYPvyai9HY
LEkjwEoLfxGkqkbeqsUdJa/EpMNxqQ6iBLvuBKUT6eaWzRXxdnHipC/gogbIB6LE
To3MkFV6fNReH6pDZw844YophE7Yyp9u2mi4cJIz9XNuMsK86VWvGRNvRWPd9gry
GSzLYNz8oSyKHlI/J50I2xhpvOu5FLghjBST+MQPYzHiTROg9qCI+SZkimU4v8XM
ps/OzKxbLQ8doR4I6kSSYa3QNohc37ZePtVaFrFHVlRfIDfhW4OM6JqtBDEwqAdS
c9Rc4bq9cUoR589vy7crZkwgdwh2iZ89LEvPprGbTIenHQgEjvMc9Xcbio3YrDqk
OX6i3ZeJlyVWnfX3Z9SO6mh8rvfSiZChFpdGdzD57nBYVBtKwfVCKpiReQv6Xz7C
h7KeXoLf+PYo97tZSw832E8XWS3DYxRl4RbDaPY+SsGAyMfazpNrg9K55kza+XdK
gF7xDa0ILsBmbt7VudUZpCRrEPP+e7Rqa554GwZcDeJUy5LXa+mnYNOzmb5shqOk
+Lt6adfmbl9XuUZppeYBuLG3amQ0m23WXqbBu3nuA/Dkm0l6c4MyDZWQC66eITT3
lxcNxF8XhrJeXheskoqdDTy2pCDx9PiWjkToAntiZ3ExaQzXZdww9+Gqxgpfpxlx
wUfr6W/e6VtIhLXGtHrpsjfrElx2CttDgI04K7PZ6rFQHLfmITR/0O+DB6IMG3Rs
5hZebhsU8ngXBMZOv6GmuS/G21DGEYvXPFZsCKLbU1sF6lV2JXfZgN4e4dxOdhPA
bVWZoq+YcARbPRbJZo56UwkGN07V4mFakT2KYuD9xNEpOr2/S32H/7cqw8EhefUq
20MUje6szIs6yEyzdZyZzP5L6qv2Kgr0rYB4uK4ctZm3Kr9HZ7LgRfV6lc1hj7cB
OcuAZ1LCuZjh9hpFDcA9/bxmStoX7Wx8t+tgFTp2K4s8rt/ICOMGPKgXDzfRm6BJ
kRmALlmJagGCHS2FskqbomsTvqXuOLqC6KZFSqz3Sd+HvhKqMHQKaPRb2y87x3r/
/xYoN2Z/dAClSQ1ALWu2qpVO08o7759J+ZBApEDx2obd9QI0CPn0qkSze3Eb0ZCI
K+1npNYr8O4HbBK29c5J3Sh1QLy7iwb4bmAqP0h2CUvMpeHz/OVltWcymoYusePo
+bEJDxCERyo/hR9mJkBbWk9VXEzu0a2G2gUunPmnxYjJy8n/QpQGePICYBfgo6oY
X35vZ+bsWP7T21JSS/uFYPLPHWgzqO3lHC3LjzMzpLWFkqsh60MuQ8tAhTK46CxP
b1870depuvTnAhO8sHcAdswe+j3F185Nf8xpyK3KCbx7YhwSonM9fCUT/hCE3HKI
IVdNIaNDo4EFBUBlhe8YRiLhTiqORkwsRF2Pe02ncxYX3W+a27xMWheLJ+iQH/ZB
7R/JKLlx2OMY/3yqY5ZBL4v44btTiKNfKZlifKcd8XUvUyhxNUlGbqn1JLWHDGdk
WeYpeWY29bhflrk4YPUNI4CJxtWUk3N94hHtqEf8O9AFW8GB/ksF0cqUfl90UFol
g9A9LcIYL9UggXRWrC76q8EmZBW41gGyQiSJhCrqLgHp561TmfkEWyt0wGGE09gS
8ZbUWkQz/1co9XyZC9Hj0jdIPAGmllekPjg9I7aI5VizmMUPAVeZiKDzxMVM7T4q
TBsPCUQkityxHXsBcGXuEH5zWTrp1SXd0nkiWU+S1MPW4nvv4mkOiJjZr0c4RRPM
RLKmoKv28ePqzXcGkQ3pTi4885B5Zjsn+WNIG6sJ18ICM1r1ZkS0VmDvn0m+jnsR
LSuG3hTBhqw6u9Ot4rY7vsakf7Bjoo3GBzFp6E5Hah5buV/mXzpCV/HD8STbXXCT
rbqjE1LPCUXCl22zVUwfvHbac2rxvZ6XTzDChgRpdYPIaq/senAwM79P/GdTMoMx
U/o+G4fvT2afOCartwK4KXSekixxiqwnaT1cwOXVV/OhWGtv7OsOafxPqT0Ulbra
f/ajz1J/H9zB2/ELjMAeKIrbpptvDI4KeHTi0kcb/0Y3x3/SllDm4pA+6jeEDqbf
KSvpIaJLUsZsIOy0hc01GPJLfIx14ZBFWho1KQ8RYcWkjdef/fryd22yTHiLEjdd
ZGsXymXSzZbx3n3hWXC7HdJdQzZskLRDWXW9T+4LuHJgmqdmZDWMphCFsqzfA1j8
3yxHgC/scenmTy8Fw9c7sj4zz+CyA1px1edBa9kH3ttYXq5r9Eu5FojgRulttVuS
yIPPI7k/9vCx5fEfZZug39NeHMiZMMPp4L2qRk/aE0aID+2laW21nbYB7li475ec
HcOw3ri/qhcge4P8R3c8xe3RuiEFKdYcV8Xwr6cj7g2twL6c2tZtlNKgy7h8uiZK
ZkVY8SlL5+NfAkPuMHUGwso0vz8zKVj1Sf6eCLw12q2SFWCE28wi4Q2f1ihvFOMi
CaBjCg28+z031OGUQVzmxlqg1KS02VgzJOuiHjnKNQxyePCtW3iw5bA+9MdpqbEY
R9NHhxAzrS1atYrKZBcZwZW0Xh+cnwjCjCfwEQLAzFHMZ5AzQ2QbXz5kZp/clb8x
Zi6hCa2ysX3C3ohQBsNIELDG1dfFCJC/NF3bJ1jpTxDPeuLAfaqUGrqJTc/tHcLr
P8lZTt7NYylGCZ2+gpPeGMAyPRjDbvMp6HGYpIQ7s2Hw5HMr+0PnAqxOnvkyKZsU
I1jYoyCfhnyu53luVKYPxpWxTmKfbQTREyGu240bu5vb1L6SYvl/Z+yEVhTOSK0r
A1+WQVg+4B6Wg7du30G5OqN0wfL/HgYP/kLUDR9+yw4VEHEKal9nRX7DMFq7kOPK
7Tyyn5pcCdejvggChAI2aqi9XfQMRVZBkeIWFeZRWx0J5xSTHZmXRHniWjAapd6N
uapIchuYh5lDAFZXw+2A8uPHuXyx6KxZz6+eO+4oGKF9pPMhWnRmjtmZ2moVwbnL
s3FqHoITPMKs7gQFY+bMiGRL1v6FrPYVnWK+uoOqbq34x/ZSiZz8VXUZ00nXNe9e
QJmLpSyR+tujcv2TJ1XNlctTRKkueZ8eoBFZPEFYNlTI+m/J1CE2Gtmj4KrT17ZX
t0Ic+FgF1N5FTyvMkBJoLP73sWMTKbd9x/ACuLTX9U3/0RuLCldfrzYWJ7zbws2X
CyDbMll3fTFuCBQYXIc7nlk2HePFQutAkwHNjr2m8wTmxYylhIVXUGzKEMkdAKW9
7kLU9EiAS3qmJst+1GX3kKOED8UaFznh3SNfA45pzAJV5jeEYt+wI6mJxpyjCDP2
VvUNdkoV0zZfnueR2ZBAtRb3wni4EQVVtjYnQK2VIkHi63/jHBMDknMhvEuAl2Dp
yGKxmoLZmS4wdadldcqpmy9MpiILZ5ezHbgcyRoogYK7CnBS5W1JDGglU6Ik+jgS
MrF/N+XaCpLjJ+lvHol988lPDVId77mrbua26GA06XT7AfzmqQQlLAtszn71v4H+
mDMnSDJrl+fBdtQu4PIMJ6OMfKU8/GiXLzFRrWSF0a+snBJ/WmMu09ppHrmH0OEu
5Zd9+XhMXrhMSkEczMqQpI860HvBxl7DS0+jcYscWCngGdvdxC45fWnF+bd7Ndpk
wKYAVhQw7LwJDKFxBLvNp0CQHiROhFPA5SDj6XH0QOLMPKYgHr6VMD3bD1VNhz44
1xs7t601VHwUxExlqufaLrEpcSXASsbK4eoo/oU7rE2p7dh1EYrcDmIBMtixH1YZ
9Zszgv7ByFCq41Yz8/EIGPFixiXzN/E00SCGmtRtj/Bh3ETE3khxtnUv0zCfzl0c
Iilwy+CiWE2sGlQx6kKknYne1euvgLws3vA2jWjXVLyJ8gqdLq6qBCT8d0Acvq5Z
3wMpxQLyglMxvoXSIvQK3s/Ez1SLlO2vDb052XLowH4aWEyJFfoh3Tbm34n3ibb3
1EaoQvdKg1ka2w8wso5YHcCDfeHDuyKnPQ8gV8iTn9QK4pbyveNnKphl8IQhRWlP
4mqubkxPo9v1/RGdkytJxXSaWPnoMiNe4TKu3fL1le/SgTaEiIyHZp4+JtM2T0si
C7X+KM1ZNnuRK8Als5QfK7kJf1uEulRy+FeSHSX/xDfoiOeEBnxtnQr+Zj5AS8M2
3gbSRHeKKD+BhsRXiTDAEro5X4WpvWl6cxSVn3sdCswEQJMGGMH3ibrvudVegyv6
rp9dOtI20p6fh6UQbiZwtJnIaBaY1UumTPGRBzRC99uFxXclC9gHSqexqjDBrsqY
KGMTWSJ82M/38RErJxTuilfiHWdkRzkxZWgjR+kccA0VRax9FGK64zankobQPULs
MokQqyIU+SuDZZj892QjfHI5b1roUIYmpGL6Hwpy52JCBAW+VEKeokB8I/t4eqkU
PGgC3fVRGQKzjvr8YUTTyiM8+/0+Bz1iI2lB6kILY27YilcOMCs42N06FRq5+Btc
Wwgnli5GTERSAjaGEv4fzindB0z9iirvxDtjhBbxhyAv3ZGQQT04DRguxdxPtVqs
G8IsMhhItX1uTB8q1NGYbSccpYAAQPHa2K4or0S3zQVSwZ6h4y7FiOeoqAAp9L2u
YEbEURnohC7zS9SQlZ8vQJOCO6r1hJLQttLkvOdGMKIEEmIwE/bFEW9fSqfC6g4T
oMOWx3wVdwinFRSGtG4lYuHN97D/0L/BiJRxaiY84abZfIBJmqo96AAqstJZI7hw
4dHVlZDNlXl8dTJFGFrTbV08INGaJEIjGvxmYhR0zrIvASp0LuG7e3Z+9Bf4xlsr
+iBLxh5Zmf5VNTNAjyRKpu0SpzUpa5f63uFZhuu9NNHGINvP4LNzeZU6DkYaAc7F
5prQG5T0qaq03TAwS/X0yLmCq/8Rt6X0eM5m7qqqwG2HDrREIDpAuSeskCTTBZFK
jUIy8cw51GzRi0Q4QdNisqmLe9SZwaea0eFIAOBY7gGP3UpXAYcN6giB+UuwqHi4
SV0wL1pbSplMFTHaFWDn5BdfqTkC1/EWgd8PqulEgHNtMh5Gnygz231Kdh37VQ60
hxDL/fd4j0NFmZ2tSaB41EaPk73crCwTUMaggG9rQgNn4pWPrfZYcK/Rxl3Pg2U+
sK/XPCFsIrsQs1jmxnKO2isKNBe019m9XMbOL/dGS5YvfAgwFEBJRTw/oEcEBhgm
72peq+a5dMbBnCqC7h8skAlQ8HhdbQ1RJ5g9zztPa6vzrXEvkXxYayS3ksE5V7qh
+W7dKnNYLTHl/uaTcotexL5Fo1g4HFoO6uMQpkZTq9DfEBNh2DXkssoLEU6Zww+6
Eyb31YooB7JNjyWjWSjx09QQW7vInSLwvnZnlta/WgUmmldhpU8yP4NB+/I11ViS
T21s9Z3vK+QN6RAEGS7KYyGQ/NHrhCh59UiNypN4f1uplmbQ1/y6A3CQ+B2ffMc+
Z32CAzSOorpybmkSgxbn2esOC+zW5Agch0onBUI1z7/C7l6e3nqcYnL2K/eIZSF6
sn9Wrj+8v9cHpiUcNw14k4yrm4sxiAZCD1p5MVS2Kyoj9lo4DTpTdhxQPW2eow4d
WCk94ZWz3OvegBv658jdXf+1FBAIwCPX+VLerfpPRit81beZkm9Dmn5M3b27fq0Y
ev/aDYHEg4meb/ZV2J65Ox/XVQPMmN3GGn2shmyh2UCV88BaZCIL8Y/uHRvurNBF
tVnCHTh+ipybTCBdP/ngd+czxYgA4rtcx3+fLSeKLFVH5pXXAtWhcX5NqakAgPY4
eq+w/rwUorjhrGxc4TyaXIqLsisqStSu6sZCaHVF4gAAfc4ycrssFfXcgvYtN9uX
SksdUkyQFjQsSWH5gMxk5sQDH/6Ns8Gb0EpfcqcNQvKsXaHt5Obu+o5VcxRTSbnI
DGQSuTzRoyWtIVinr7U0ZK4VPOTsolmNN6x0ajqJNrgI14/cG7TGS3cOE3KcOtYx
a4uSiTabGlcdobPBGEeOkBZJtnkuoEO90zsYXYWdyG7hXFR8C6a+9jbWCV49gNyu
yYlsmzqptUgXaChZM1+ke3qZ/rELVWkNs2+vCMFHgWA53GmzgD3cp/o6AaB8I1f+
9EQy3XBGe5e8QeUJ+pTJPmJbVCLq6orIQDm0D0IZ3+kF7HqwoxTJ6TD+0wa24EJa
Uxd/KuIcdh/3icLvya1tdyrJWOtmazTSuYxs7XVEwNgrnWVSfejkSydSdU9c/T6t
pZuF5bYDXLmy0mx3GupQbF6N0QGdi0bAt6CgNHVhSnBjccZMXl6haGi21l5O5EBD
THR6VEeDno+EDXNoc3Vm3HQi7GkHumrSpM1hP9204ded8a9R07R8o+BfDG4/dF10
J8DqddVcptqXjSV2YHv2J00mVT6hG76YdhWrjh8nEDDPBi+k0dbJm7+mL1Pss6Gv
9A2rDWRNKeVt05MQbLuPJ4RsY4EsLvhr7cxa9qH3f7pCVMals5C9E1cGgU1ha7c1
WRsLcNp2jGzZLbtEDxD9fQd1Mk4MnEs7zpIdgITubuD9MLWJtO78pUFGqECJJ85C
WnpDzf19dySNXQYfSjKPwxWf5aZLFhGo++D2fuQ8d9yKcZcffXu1Onv91tlS4SRY
BjEkAc1ARnBhuB9cIziNs7n2jcrw7H7OLaa6cW8cPeCiiq9/5c44bfMA08i5/zMF
b2IEQ4rOYS1D7YfXcSDgvcZ4wOcBkguyDID/ZnsFZ9LDk65DfWKTUKTcJf/XW6j2
tSSiFZow93JpGW9Rgk0fEmAo7Z7CyMug9TSjfQr8HYWMCZLXdc45ub+uCYQ8cvGX
V69D6AEWFSWh6CWSOuCAzV13HnSbPXsOwjdpd8U04oPKDb1RDEHkBzT0V18oJCuy
L+6SOU9vpewDF/rLooYkWlylPZPcSuqy9v131FIh9l1QBL67Lymiq5RfARr00m0G
3Gz3Ux0uMYS20VMdTkkE1x6N8C5AxVGcDwFV7Pwlq6fklxzpsfxiHun0+6K0iDsK
NJW5bQ8sedBK7nCK8Z6dF2LqhwSKjHgIiJ2OQLZxww7K7+r8IqRJp1PRuRN3Av3W
Qsk0bYAkO/1/yfiU8W9LzRclPRJKuuWhcuMezi7mI63EeNuYPMR1MFrjQ+zRqMyO
KUa75cAStm5jWfe30AJBvpbC3gGDFT4kFyQl5FQ3RQbT7XvRnAQ2o0HEGTK7Zjpf
IzAIavOpTBFIEaz1zHQgyjhMnvZH5E7AmOMQq+ByoBEDW2XK5XqCXo28qWsQCEf4
C0Desoj1w5UQ9141ag6fdB+//kA7nKjHHMAI2fFc8M+pInqWjaaXd34L/JQi6HZg
Xq1x6ywkt9GnLYvB+6r1cZHPSc9M89tTFFTSNmeJiKzQDSr35XLCT1Q0tAWYpGbb
Vk728BUJaZQHVEMITmWiSkpjJFHM+4+SJhecw9PraumrL6zP+V85kaoRK/ZIkP2V
buMPUxYOkikg27/MgzD0rSHQAfyx6qH2JFus38F+c7s8C8YjbTaKgu/kn+APUNZe
VDAKAmZ7nmpzE7VQ2+Waqrn0Ksnyhk2scxnQTAioKI1+vzri3Mr+g89aYMXy19GY
SXwCFlifD2kB06nCd7X70zVhUqu5o3i+YQFmaWRFSd+XJxvEoybh6KuSCXGAAp70
Z8e5dtGj4GePaADEH374NYHcYTZAjwtjH9Bb2Ty0XcsOYOMm+siVinsOc2u/kEbv
4GOsAeiBU7TXI7N77C2wnJ7lA7n4xcHpY89PBobG+l6GdKOaGRVc2Sfx3uGhGfYn
NxFxiteQKBUfWVedOZWfh03mU7wc5X83viMsYG8vcL1EySZhFBHaUBZNMF+dCHIK
ZYGUP3lInIBYXnXRBFZwZozmK+ML4B1chDLBj5lV3hB85Cl3wGY+odKXpXHgFNhz
AdnzJz/oa4eGe0WSw+PteiRzO2hS9F+LRXynsd1nBJKWTNxkKWmp8TpwH3FgpgH/
b1XY8j/rTgJcD720ho7zob2jkltb6jSIjz/lnI8MGmzaA6B7YY8Np6oizsp+8vTt
4SemX0YvGXyJvc6FePiAVNyZv0AYZgJx7Ylo3m0nohPe/+FM/Cflwo1KA3l4gDxU
1sfRaB+qxvHvq3VHmEjSXHFcJ1nCrkvBfsCq1rR2+cKxemB/ELrNLNEcqd7rAwcv
mtrDTmj2xeEOxi1d+ok1Hd2wLNaIMFyfgoEA6PLxb2YZEn/Dw8Ki9fmRvAIVGAgG
nUXIQ3WYo5cmb2sPo6Xjo2d+aCJh+W/WL9Oi0frS05TswBK2yoPVXje7e9+CeRjk
bmRXtjLQ/fGKhdZ9AxnEpiWkeNF59rC5HXH3BXlFyKJTCLzK02em3tk3qtHJ2Ppy
Vp0+MCog1OoO4wXCPgj727bLcRznt5ZqRLnT4n9h9AMK4ugSoRa0FshdRsAentJt
QezQSjXMD06pZnbiv99DNJf8LvR3agbaJk39T/N2CTxOJyp/01P+KFG7l+bwWQX+
NUQfu8G/ZW2SGxhCykv2NsR4Ltx5GUlSuYGTuPi2xJLvxNwU7AprQxV0rdc9oJ+z
JGPda8D0K7PM0xxzNvIjoz1HQiysRsomOjtdRa9quEKsZVevERmExpRa/+l4zCQm
xskPyNkVqqudU9YsIZj7tk6UviW8Y9vQLdgSQimSjjVNe1bJwDZ0VyYcq8DDV/Sc
LxtqT6swR86nBbPbjacPtUIldMCig6CPvNWHc8EapGELAaWPn9Mu9a746UMfmNsW
HZ37FgqjeAmnEGeOKJT45bHkE2CszImCRju2OtgrOBdhndwSNMmGKNcQUCZD1qN+
sGiWkdCpmk4132nPFkH7UnDaW9eZNDRCqPoojQyTMv6hl9U0CnANqTJPqZpSmy7+
Sr1girO8A7SHdiYhKZDY7Uzd2omJmYvHuCsBxARu357zxasgWM6I7eqBlYxKDfET
jku+TPYfYPR3cTfpaU0YtDtfrHeLzy+73CgL02e7UExg05JPZp5VgX6aU2J94ilz
Pen6nLeMBstkcG2oDtkhHadILqaTSdwul+j6OHbJv6hCNgnIwghOfPsJlmMTLMVe
MwUQTC5wb2oZUNVXS0G0tc2y0aS+QXny53QMRC3iAqBYIWPX5c33jwf1jgIxs/zy
uw+yy34P+kIW+II8CzKMDutvWDycsXZVjWJI6FU/erE31w09ecFvUoIxecOHIIn+
eroeYKq7fjNKPvsmoeUcmb/Nu2uuFRQSKNAk58Ko2MYQVj1c0+/3m/JSzDdApFqY
Y9VkhmgkIDV7B4Bgkk3FQHzue4uhnYGw62+aTzhkqmbk7sCJ1p/WNF1ygR1Mqst9
pW78LVromn/oQAHilK2nIAnu72XbDkt37Pf+OP6sWkasvaYAkJtzzimgNlw2Alry
3JfaNRIXgpY78/N6cl9lD9U30WB15gjg42zF+Ku9n6EytlnU+jsHw+09YyO8iFvZ
chiICu8uqhrjZ2wcJjVsBRxmnANNNj+flAq7tX4nJGH1nGybsNixg7FDF2O9eN5q
xv9Oz88UH/3fjM4YAaLWh1xW5ZeMoUemNzNNCxEquvnT1BsXtK2Up+4wOILuwsAM
ncEFSnVI5O3/VyKB+AKEMEM65cbgLHB+0BS3lb0UrL9qGGLXMLsWPMdBbtzkEH8w
NWyVA2wR82NfUt5g04+ZphM0CceCeniUucXveYjH7Xo8RChrwXIvavlpWKjqZ2fI
4BllYuY/YBts/oFE34Lqdc6PgbAb3Jeco+PpjlA44S02ycxn7DxrWBLV86oo1RZA
vFjBIeGrfd7E31zH8k7MuSSAOkH31o0yE4mePhKTX7jB7deZzFxqPyJ+vZSaNhvQ
2gsothHnH0UWbQaj48ddxUImXpg4rGR8rb7mOMxqlZnvmJ6k7hwnoSaJ/bsrwYW2
vtG9ZkWDYeGHvglpMRcqdpCdVxIjHe5Qw3aVvdNxEqC5BkGR4yS8BKMl5NFU5Swl
UQ7Ik3mV1C7V2PfHB4UxDcfcxbV/vFKBuJzh4Gr6qxZUVNaMTuqSgiXbvHOiQpdf
EWOoDsYwB+UV/+rSEMPSSfuSEkZP2emZNvcLTGCU+TFHGG+OqsK3XSouOfgk7ZM/
+l69hRsCNt+hmyo2ontbmOSAP0HQ6PxGgk8kJksZgNHiOAq8wQvCXG/lHwZdvv9d
/pfVplSpyNST3jhZ1lMf7nJFwAubivZnFSRlnhMRVWCVG2XQ64JLEHOR3cdgLxO2
oaOLw6WzsHkDpG8zJp4y7DWemsqjyzpH6VVoD7ad2W9ApxoDtZ2b5VR/1sY9W4gU
hkC3yP6HzISqIwNsO966Df08Kjh9TfTVicwOKONAdPqJTekRdBaohwmLHmtk/eL5
ftvruDrTZvpuOvG16qQOkKW/05sC8HijJtLazBlXidli0RjSd1kYIe8/ZAnJP9d2
J4sG73S6K9WJdYdywhBpoGpEZSgjCGSyAjTNVtVQgz5I1p4Z3CWEwbws7skulyIc
RBRvQLHPe2cxLy7TtHawCE5dYuB4XEBQ+06rzYapP99DxvDJonoBucpul3wGJV4D
EIwlnTRsyxpuUhjSKqKZqqoo4gX4BM20iT9XG/c5zES+YVbbPVhcFPF4/M02fDOM
JeztOn0qqW/q472dJK3XG6Dn6VSV8+atUJDKRcy8QSnX1D8haYYNRwfXPl0dJ+Gl
5mYN0py+EMqqTnyGvXzQNZRS7/TTVeXei9GZSoiIuJO0NHLk40eH+mzJDi540ujQ
P2d4ZUBF0c439SHMXzvamlcgMdLS7SgfAcEsJFQ4voWGi9EL/9gc+YeBp14axz8H
bi4gJ/4LbUEjx/17DSr18ZmH7xRKSXcw62eA0Bp9ge93nVzhlrcT+WwAEdHYCQxh
llKRlIsd8F1c8ws45pJ1vD78RW9rjnn+LYlz9fMTm0L4iZA3XlHLaH9uNjlzHJsr
pA3K+Uv/okiK/vaDleSoTOglezjoZ2sR/8s1nN7vRJ34f/YhWZQSB46MN24werMc
E7Qwm9Pd25UjLueJod3Si6upZIO3JgJIs7J5Nh/VQ+U8o6+YrSUE2hpShXjiOquB
fb+TnqghQi0KuRde12DvumWA6IRwjVpxoY6JV7hV9VUWZ3DgMwDJTaj7NfG+ph6Q
w+Qb4HMhmPW2RlHTpqq2u2uEe2w7gBCXel1Kcs3KLCwy2I158Qxip+Y695FvF6q9
07yQI41oxcZiagPXPFYHSi5CSSNGXkte34hhO0P6oYFvxHcA8n2D5WIK0O/StQFL
o8ofnZ8i/k8MYiToZH4DmuXGNWNGNGubw30s1cCC1xESaH6acXnNU58NEOze5gzQ
oN6+4/EFkf/56YG/8ZmqEl7mWZ2+tfL0YCk2WW2jyXdqRgSiR7kOUmi9PRyDXtRt
ionTWRLbiiJn4fMDZDmvgCTG6GrVatvr2Ce7SsObzJAuZZfpufUyRHADVaek1/2A
ZRGPek+kbbAP2N7dZapjkc5fKC2jyvD2Ip349Nw8mY1dayhmcBw8/zoDhcBPkFeS
4nXsC72Wx7gZII6yKGfqtbW2J4F//8olxI868BQCCNufhjy/BdoonzRv30rh/tIG
sc7eSKuNyJjKYs0q6umFSDQv3wHXkr8ag9SdWdgGeTdYvoSMblOC0f6f93n5WPA/
nTVDl9kNCydilukWSUXnkzNHeEB8xXVkR547C86xZQLwF3mh41qqhaBVWhT0qiTr
2poso6XdcwUgFs+ngD3rBIlNqkuHn5Yk16QzQaRP5YdzdjYH/2HZXOHqy9kYT5lc
YxexKlCgswJ+qLHqggzYhsPxC4A+E02wDRiqLpZT4X8Df/2tjjbbiXJWdiZtAVcn
r6yQAR6ucTf8CvEd4GI80dUBY8WL9Udfbc+g9DfzEG6SEGHeiIv7plpVf6dHYQLm
iD1YGvAMqYK1U7DOk52BhdqGHoGHPZrc5z17w0tmvB2U2G6n54grnGcV7W9VLiKI
a6PLnhgp1L5nVZRlf6MV/miXMNKpYjyEioQ9NB5lHDFvTc3E2OLFrTE4LpYOzL3Y
+XzAvnwFrztZ4LvSlyHJGBAVCU5+av6k/Gd0gk6qrI6IJKPqRo3CAHojt3iH7nkM
vguZRnxcmsmhfREOtKpDTRSyJBvFf7RV7uDaOhUDrFIWd0DHZiWP1z0cD39+kJR1
0ct8WmxgA95LSA44iwrt/d/ALmgMRl/x21NRckScZzGO/dznfA3RtX5+PwYubvEZ
QQ9WDUQSHsw3r3NGYbu0xnQF51w9NP7GfLydWzgKk4770s6TRcV2TEYCmIjEA5Xk
yti5WEEeB6WuUoHd3mx7Pntjx1DByGzXAVZLAVlGTtEt2JxJTjMKvIkFJaF3BLwi
U7B28WKxWhbQYlI0jmgIWpn8dyiASe+mj3j79FPg/PdH7JRt9tI5nLHiVBjjvZ8D
8v8Jr96AMG1VE2b3VMJHompeokoL1wOnCHXH0682IrwJE5z9H8y3cXnSa0FSxB/2
CqLh9v61fT8otDvvD+bgRmJIJ0CrdyDqftHNDkyf/kwnfOni3E+mdRSoa6796yl5
gcXhuCMzsgr/obxG+cLcQvCKxSaIoCDnNYDRtXzQJyMIL0e0PiMz0GYoxRCMz9d+
YdzmajKoJIVjpMsHxCEQPld4NypIgpFsGXvJ8QjZ/T1/aC6a8+YX8bt2mGw3Dce5
OZtmhokQZs9H3yysvPFdYgsuuentCR/8M42VPUzwX8XfSdqAoRVv1aY650+kVAy8
ousPNdEDkwohHXJtTk5F36ERKAYJBMMH1vUrgo1Z4KHLCbVq1JJU38t2J2L6cHWF
FUfQ1ramNo5ox9tXH1QzKsBVhxwRLU0SIQV651bVnZhPbrGCZB3y7/Jk71aXL55m
0F8czxOHLBJF46fER+3B8SvLaOV7lw7aX3bpiUekjK+Gxzui7tl50fe+JzCD2cK/
QqBh3Yny4cb8Io1qoNOpPgyHDL92jfwZMUySFpcFvPBkYmPyQ4qKv03KqaXcH9pi
dD/l15aBrPJgTrXVRkfRUEbXmRfwfipn6Uez+TTZa4JH2pCeW2vKrZQCM3Jo8m/I
A4k842rgc4h/SdcxsVr/2ZLNwA/4S6f8jWFZs459AlLa01gUj4OGmS0ZfmlefbWG
kyL9lOPKRjynSUSXAyxD9a/RBnxTPXBfPobFhyme1IPOBoierPZ0vP2nV1RHVLJj
JzkQAvSDm2tNYgheaZI1wTq455dEwUXRcCHXtlW1WPkVmXZn07bmmCrswdUpzB9y
UrS8c1NbSDGfTX1Yq9XqVdQKtcuGoUfKrHjhdL3hdOMkOmz0vb40ggtbkIoDtzs2
200NDfONlJXmJLNe9EtfN73mA40qLeDtwh9kzokU5E6fTZyDUEszheLv7W18QPH6
OV4bfc2euYQHuiyWoJV7xHaqqNLq75ok+vsUVPvJ6/yJhnMvcg10vqNi3lMqkecn
Gy+PBOoktLGWp7BRQr9MXr6iNilGvEiO3bMoP7KNgamsQ2lJqpYS0Uwy/+jQMYf5
RQmx8k354VqzRLA+hLao6AJ66tFZUwvzX6r3p58Mhg7qrgIbwVtISy73+0nLbfbK
CdABSb/ZIS3bwKrpI9AfqBje+Q+5qk59YR1Re0o1/TC8AlTZKNIfbqQoLZqR3+Gq
AdxowN6i8gkFJBJp1THotlWXupivHMCRqxNORZdLjKBe4cGSUl2cxYP1exC33Ppg
K5Fk874tTTL0IkubRLYEr5zZ2h5HBf/BmqpXpVbTLvPwoXNUCRFCjJ59mLwC0Nhh
QZP4yUh9/i8m4HxQDr0hBHF/+8co7fA82oc+X3HYeNmA9hsBv5g1U+ufKA1gcsXz
/VtcK7gRT5uFfEoeR4LmHnpMAkJT3oNo7dbg5waJfgh77zVdFAyjx7boCLy780ck
zFCOaLqM3Dbgo4d4GCaATsJHzpJebDN4+T00jtRru9tcTOTxLKc6nmCFr92v+7aD
epuZi73JEFsX+x/uf5AjkqfxR3xPEmlrIQZ0dT8U67U/1njdICSFQMKlOUwR/CtR
rXQ8+Osc8rbMDsNtW0YiwxXTl1dlBJonOTnOpS4rVs0FRP61AEzoJap6MKj9Q6yH
9tEhqai4zqjToJtPlV8UIrFCTKfeUOhrV/rwly/YOROFdQ+XBDxaMNxGHNjzUeE2
RwsTO/aRs72hja9GiatCXwnZWuFrF5tn0wOLScULatlOpR+eqfavcNV5GVO6StdR
BqFVbbPfeojiZKRG9IacPNNEzVMUJY4TPXz4xC3s3O1PgT/segch2BfP7U6XdlxY
SQlWVvsv9JWMHp83nlojbGrnlXvWfwAq986EENCGKWrHLRHaD6r5QGgzGVPD4VWy
QjB+OkY6yvy4Oxkm78ZivFZaY1VPxB5pM1Jjf6VlAqOb9fBX2k8CJEgbQJwbvmBQ
rzzEGXQIefPu9J28JY6Y6Qs8fWtCehae05MVXUYGZI7GDlwf67hhLAyCzFF7Ol3r
bqgUhTaTwpQrpmuSyK2OhXePgsDlvfAoLRQv+J8FrV/BnIeJ+jVTaUGb3FWOLEVd
EhbL7GYPDT3FRGfZHbPRTs2BylxsFov0XVIyX8+UAzEyTClAsulL78zRwJQziXoy
WMuSJiYxb2bnbjctpLsD7c8+9IKigs0dXBpi3IDZJHU/kFvoMqWhqp0jKwQ03ukL
eAd4UR8qH07fzMbYFV+kUSrwLYlcmn0QfpOPB9LTtYNFlrDtR02l++O5P09nFvtu
G2jJi+UXUVGUUpwIt7WSOwdUsIFNz0X55PpStm3VCmLubDQzAxE4MQanLB/WVA/s
jJJQumIt5mPWyzH9Lyc9x0Dys9yh+fVf227NjQk3sjOfhJsqO+xpK9Ohqte+RkDU
4rlUkHTSYLCsX/0OckkmyEJiiADez+dov2LWaOufA+7icebXm3D7OfPPKCt/WD/z
GNY0I5lBpkLkedcRdxybfekZnYsAyNU4Wl4lmZWt8glKbJ+hHGCVHhCRPFDCutsd
Osn/X0q/VTjStMloVhEOWYdFsWVJBMoIQLLrVL8WPsr7+O5qT/VtjpEUq2xWU/Xu
3x8Sj116FvYmTaUSACSszI+t4mCF1Qtknt9E56bvm2F4U9PCdUG0sQ1sfJ2Wu2ya
dtEyGjjxWwYUbHyeP2dlw+cTGtTMvnI7YOCyXSki9+xX3yRbwmL5D/EpKgZWAZZh
j/7RmfWxVUUl5DhAbfwEwD6STirdUBBrGmuZ4TCwj2kC/P3fQn5e2nnAVDbUHMAJ
H++wCM3BjjdPijN8aC26Bb18NfheLxxxhDf6chwCTXfndLWggFNUGSrbLvcI5SeZ
ydRnBU0Y/ntj17MDEFNapxSDyvyT5joNmYXkIUGvrt41XJBO/rg2wFwobXLg49tl
VqMpCZ7PQoCAbOYv6C6qJTebISPlK0aZi3DDbGlMSXGx1CBA10a4q/ObmuIavQcN
h/xsIrQvboVUOL/I5KSIh76I7efeaJD5X7BqhKdpm+HagHKAqa4KgCRXRBhr9iL7
mA8y2faTozkjCYbTI/16aFn/LaS7IdCVpRnevgBofEkFpYDCHf3hYIT2J8mMqvwb
LjBA4TtxVm7vBNjCipa6gAiuzGOtZLY3JCHdxyWWIhASEbCFFS1gnX7UrZ8yxA5U
CWEzWDs6FMAylqU+Ulb+B0/brNOhZ1kwjxnWbiUagKV1koo4Mu9+uNCuBdVAdGnL
wpV0HtqKURNAAHOtjaXZYgnAGAySemhc7KaCSmwEta+J678RMhxYMrFmbTjAd56O
xG9JpFKjnJKvewWhwqikQS96cfTay4Px+d3MUcPFYfoqerBVGPCPLPurrNnW1Mnx
fkfP9c5hmUTXuyh/qJGHdRhaAud5fZkTL+kii8BgDAcwyrr/abkywrZKRtt+haxs
/nDXm72iVxkf+e9O7IW3YiO/kjaH3UwwvCvHK0SmBFyFh4SeDVvPanNy95GJwOuI
/SCM1l+9+69HDdSVTdrn1085tpnQiye3nbkTj9BuQKroSkQ/IDpVexUQELoTuJtB
q4LJ+w7jWrCvfA/D6Uvqiu78vCDtR2pMI4DBmrKyM90Smcryi3VA2B/fJwpTQtM2
KQw4CXHF45Ri+h+/gzaEF60QuTryi2th8tREkKhrpykOhTMSJQ+u8p/EcqRkDljQ
xoxuDi+h/un0v1Y+8xb32fsQS9GhGxfzM1jn8W/AeVKS9UkBkrR8JOfk+cQ4QV+W
pGvIxkPGauXJ1tdkN2ivh/CyqzF23IaWjY2WS5E1nZnjbymmHYHXjc0EWM3WEfaa
zUmyR+KavvtZsBeYV4MM/LA8OpNRGLxRtDkUn+WRoI4fAxtDtLBEMI38nuUQN/4Z
Ct3wsbvC3YrTcEL4hnJ97u9bt0iHe5iczJGvXbpWL+99BQhrRUg9P+XNcogSyJiD
x9OmVjwq2SO/OzcUfd8+8NYxmfu1o9JaeiWHRxQGOzQWZsGs8rbqJa/oi4sN+Mme
0MQWAbCPLcGenVhYuWU+3dou7DK4NwlbWnsjwZXoVWKTOep8riXE59Z9V9ytGIeV
lLbrJ0uJHyxoOYvGVpuWHJCWBzqgP0xtPeu99u2i98Ce1Wr9t2kZHdjrxOQFv5d6
rrhjLGdW5h/kZa1G2IcSjd/cqCTAfPjHulIosk1yVGnUKmjNHGQR1h1xVOi9BQzi
szbJ7qMiihcms6w9w/4U1jg6U6//bmkeM95qvsehG4xB++QO1S+zFMN/98kMlAaN
rXpalu08EqeEmFRCsjfMgApZfneLzvmT28XhxYPCryITTgJhMlsvT84HApWKHEIh
2QBHBGCrmw7FZcXJAo+nGAbNenpBTKUIFeT5faPHzj/+lpDlsfmUXXKhbd4NLINR
qV6n1s2fNT5f04cE9eXjKl8EZnTki+fHdG0rW3Svu4R3VIEoIvGouw/CP+14k06l
4r4t6hLgfsekywXKQIjRFTbzHmuezpp/rf1IvBuneUY6V79Yt0OThAGNzI25WlzE
NaQTPrF/1kj8IXOeiOhVmbbOjVKnXRPMomvgf++Cjvn2Mm0/9C9LJDfjWE3rd4D7
Uzgpti3THKRuyQlKZ22+zEzS1bEsWQ+orRJZ/9kyMoJqytv51v1Af1i5rvhA4fal
Od70nvNWAKrz8JTEEfqxAF0j7x6JzbBWS42awzzWwQY/90nU9wfYGvHXfHP4kXwJ
HEy2Mhly8IpeQ2WcKo+gkV0AqxPUeCwFwBHxgQq5hYIxjwgvXW6qvQgx18jSsJMx
v7a6cr+OF0nWUsNThznjyBZSx0kawobE86hkT6aDamQ5mq36qEWS5N7LaG7Q1a+s
EBCTkPU1sHBVCEwKNzrwxV+jee30tu9qF2L0sqPuo7WFFrsCVYQva9DHC/8qoQCq
oYjTjjGlhDgH73u5N3B2wDkhl0eESDdAuBSsj6XHcNPDzqJnLRCicqwMkqp/YjmG
pcnW2a05meeU+T9Pl4gzymG1DtkWjJXe3DTBVUfKfxr0841C0IcJve5t7U+oKW7y
Kilk3O7LEK31F0KTFmNG9oylmkECKgNNT2HBFDYAYEF0to41qf+kL3+ekagFy587
yXi5Vsq9PIdjfZ9lUOrPGPSrTcq+UmUbzoh1Xe0LL+Uihfo07EmBCCjpOjHhULLs
B9O5xU69b4DVbNMvl/hbV4lfSFL45/jgGuP0oTtjtgF5aYL0i2AXDitJJT6cTmCE
bq3CpGLToKH4oYGfl9kz4nU7gCxMOd3h8KRKYIP07BPy6fED2zy4A2t2/rOqU2Xa
wHMADzynd7TVPjS7NbH9slw8SfcKak6L2wtO81ysutoOG7udDZQ9N57QygU8zcyn
f6yhq+FCNKpYqS0WcVhKCgV3FEZ3rnlG1Ri7HNZb/ROCS3faKECGt+imO9scutJb
MAuobXZeFI+5tD/ENZQkVE2OzZTIjPLVmtaZ7m8Hf+l4lyWWR3VIdx7MSpiEgrFu
4I80bvCyVi+KS1LHKt/ADTwtU0hEHq5qWYlZpTCVB90p09jXlW1XRIjPNesLsLaY
3y4SCPAep4TfthKGl/qJGCmaOPSp+6a/rojy5dEuWSifdLPhrd0Xx6kB3GvSPHp3
ZRqi5Npg+6x6GowhgFvEJXO5RpdymZ2yjdqEtnyes/Ztru0+2Mdhq/cR3V3y+oOM
632zOYHV6iyUmvxZcvshxwCZPEXinAAJT5H2nmqtZu2s68eZFDRCuGpbbBvDesko
VqHdD3Vm1vt5e6/chQDYQ5HU27I1u8FuAWkpshWQ85uVcCCpa02o3K4q+nGkU4AX
/ZYnLo1GuxB/9+Xj+IkP+aCc8ocxQvtVxNcdR5jq6hcsz4ePnBMqbWqP9YI2PHe0
NN9o720Pg2K08ec/dMyUYNdimyC0ZOIk5XCW3oPlpcY1grpg/BPdTCLJf2bXxvRt
KPMx7nGcZ7uqbwNzhWqnqTunzPvB9pUEi/PQTuop/MostzgRKhlAD6ynYEMwUFgv
PRj0Id+2ESl6Ge6upq5zc2lkwPa36JoaKETaqg8Pcq/Zw5BfRQ6t8vYYwu5ZOGSU
7naDOCCRxQeskh0W4orXzFaFTzGYsoyqxV5qgv2FWG8960t9w0wJtFz6I3b0eb8a
apA7/PKqgMKGwJsLHT3GV+o7fBlOm+ASQ3LYdaLF9elGGclpeB5Q0b5Geo0T0a2t
hPHnIi+jH7KmG9mvu40OF2lInpbwN8AExRMXZr9gJZYGHyJGKjpWRqfmxzKmhapW
KTaTy3hYIxOILVhJ11f98Qd2p4UMN0pSOGwRBjfUnGcZREVKKCNdanDIUXD26Mlt
+xGaFrpX66cSyRifs+Iw4NpmmPpONgMdXZvGBYONUyYKjsER8H5l7Th7NiWYFgrm
Pen1usRWK3NrGY922FlThr+HfxgrPBcyulnlSTUHNO2PUmcx6we0B2dtHO6wE7q0
G4A1VyoJ4Q1XWYbDVqP5zEkwREpzak8PbtvOtpbBsN9Qg45qENsBC0lWPY60wMNP
+HyVTqFbmuE/tm3Mmv3SPJ5hNohCNkoWAVba4fAzSSscydlKW5NPgM1czuCRuVx3
0pogJuhhOtWnskL5DmVII2UBuMaMd1gJdkarWNocStBd1EjqmzKF+xw6N187By1J
C2LI0G7BsliXVFz27AdHXzvcmkRqeEZiB9IktDgzkFf3l6fRRmXqawNltvvJHM5Y
cOvyTDhgihrPIAHycqVnzQ7a45LvoZ1mLwvdYJUciNvE37eiqcGo0CkXmXkDW/Bh
vsbpYxAx7HANfKAK8orBqj09o6QTaqKfxM0KXASCg/JdLnjmCsJOY2XPLL7H0t6z
/ISYwrTohd2msuRwmJjLNT1HF/P5ud1EmimTybWdQbSS/6sxDRrWrnsw50N/Z8Xo
j2tjLiqPuhZLuFCy1wF8teQ2rPJ2/YwgvwazyPsNLPffIBcfTA734dzP7iOvsqiY
C8ukW7sxp6Zo6UZHhBwZHtfDRvmfwyBjPlZ60L7HLzpCcfSiWw2HImnByQ+EEbDL
fwYl9kse7JXGiCKZ3tgOSf+8geOI81dxQL/FTuBBLU7loxvbC0vZNKHEIX5qjGM6
JDM2AzuR9Yv26bewuocTvLkpAlcbFAzIaNWPGbfXfBePKm/GitEkY7i4Z7REazO+
QKctwCMe76TTbN+tQkEnNwrQ8HpbOa5JY6z8bOmsLdAz8XAutfRD0FKZpsuq9V0g
TzHCoy3MSwfPt5jgzlC0UWtxAho6hAz8T8PIeiMCnOsvgbs6ieSmtNVQBo+hqwUB
o6KXmXK8qtS+J4AZw9h+4ElBFdR2EKP7InA98U7N/Bh6i2FpDzokKTjUTt0+CTQU
HpHJz/DjBgx2sGuJnr/zZ8Xi9T/2vkHucfGvSNlTt0MIKTv0qzuixwg6AZQZ9uuO
F1pbVUrf3Z4apFk/LuK2e+kBb9+UyB0gZH/HnK7yz8Ze/s/ocaxxRnHNrzdoYqqv
AKElR18XBkgcUkYGOauwUKU6w/Fuc2BE+Jkh6RyrAoAuNhaABkVEpNljZOyuhpur
+fHAnOguDj4mX7RRVcQgvifOQUjWY5g+PCsIb3vgzAZJykjJfXlO+FcNhd9iycY5
EuZRvr9pBJ/Mvq7AqxxtqfPF7G1B9hdvb+K3m4EuSfV05ILqKVbZJ/hd3l84wYdb
owNbW3K/gZ5/a0PfSyHxMO337MoFNYj1kK/PqckO7fwFLr/uskbcZ0RACKsSymbO
a5H01tse7W7aFsKvK0EiQ5nzrwb3r88jGKFT2pqKse6S5Ms6So+1/TOwSn9wfupV
TXhi+cbBmChRfiTiGglrXxN5Y563wOTcnjEp99ToMD3Q7TZYencMCD4PPpvUbWgZ
U8+BizRsL0GfVNRD4YVlJoOYWLyDfzpbCbles7qLVzXo7X1d8ttDKzKn7E1OZiMl
yqnZys1TMBoqFYKRm/nM55rYhlfr+8LCGpAq96IA6M2AWluhJaFDTnuBaU/ybPrC
3w22TfvmFdlWJXxAsbAoKA3mYMsDthbnskrikerbbZkULkY1RxP/iOOsaEnWqCrw
GtH5BJjzON4eDNziqNekG2Ma/4qMbE2IlBvtJteFBhpQH9Ri1cOQ333eFmkpHPEo
QxrosfDlOpkDSx+ciYkegNGUCTSyHLFqjFu32HqNE/IULiHM2Rhj3xbTfHPGd1pT
i0dWTVvR9KRrZrUQXnuTqpHYNLc+yqxJo0OvM+8oSYe+ujA15WYdA7lvlMHX5XGy
oIDsvNdlxKMiitMLKLYMMuwvZIGD0RGHALb9GLrbj9DoMtN2beZEwffiSHf098Qb
LkNqJMYnlBNx+Sc7OaOA99616p7/p8mW6uY3i8VkeCQ7CxANtHACi0i5dMP0kBTy
jB8SkEHYtvWIVl4HlfWTv4iJxu0vXblYQbwgL9BKD7bDmVKIJVeGoPj8hE3mRbHy
EsZBYb0gHyxYL4Mf1Bc1ZgP+f94gNg+VKPMx+8YoJvvm+sABeGc35YU6ryUpP4IR
2ct9cPPCTmeyUew+jTomt7G0mwGBrXyNQpVIz0FjaGMPE9OZdkW+/PIMmgpNTChu
zKBf4zspzJP9hrs3hHOOa2XtVJrjzw8rpsRO1bD6OL6fWP6xPRmt8omtlunRu4Hs
ubh51TIPMmDCL9hrmq0bCwn9ubBajWOaIeglEMqU9xt3ZMeCD1VOZi6Y9vsbLQtm
R3q8MAQkx5b4PBwOfXPkaLGbGW9Puq59dYAgU6xVcfCc9GXaPm6B+t1opCe9dAhG
RS+OyuLys6ZRYPXZdoK8URj9g46dGAIxf/QrezuwEYVewwOuS5PNgCzfP2dbuao7
t1aBe1bmQhCObpdRrpc15GKSPw42hz9KCywaq9KtYyy9QeyknxnAgExHmz2HeroC
4Rvb7K3HawAKUClxk+wLkETUsQaFa2MNzNekdg3g15kIUIXfL0TO9A5x+k//wCdf
ghYQYiObG7ksiSaOuJ1SFOBG5vY0qkbmDB4DzTAX9UMLiN9AYH2AYwwTfJT/b2I7
JcwImiW6GNMas9KUyILAV7U1Pjo6NIbvse4bJziJOVXRtAfuCymXRH1qDYODyFs+
gspuZxd0mbjaQPiq5zjVBYhY5bCysmLexe1LhdAz4sOHmllYKY+udip8N2VtJG+K
sIz9fR25/ycj5LlgAVq195RmULuI45eeDIGuxT1UxKgVnfLZe79DKYMFn0vDjEXf
SuiZXA6q3UcO/DOB+Ilm9lPl609qFP2WmKL9nFp2cNN/tI66FQfA9ZHoT0HyWr2l
X/Za14a7EVol/rlxnI9cHqxHmoNOPomvx6m/GaaI+97Eblr21RCcFg7xoQXoDfoF
jS2TtEbwiInTYCtubf5F2X8/cOqmatMx3gybYubv1Sc6S4Q3WeY7KPwKxd4geVun
i992Ag7SCq9HAaGJaTEHtr5ciQ8VL1isTbK+OnpmvjyV0rh35yHl8CXdJq0rkn+Z
DBI8J4UrRzfKCMq1Gp4vXEoMDjuQ3lRwXF3vM6FrEuHudd8rml3ZXpxv2kUqfM6J
IdDzxvtzifFHvYkjVg0Xu/KuzinUsUn04m1j1jXMt5eEu0ADusvAYurQlIxWYiZz
gsQs5vFlKYbQ1aPbZeGtI4InKZzWHKuFzjOr0HINz804eUGtMwToFi8wyqAxNKyd
94HCPHcaqEHMXM3eJTfiKa4s7oR2MQ6vjPS+epg/XejbrIKd5XWJSAEfmsRkkCrr
R2AQm+f17CVgoJx47EFTA/+3swSjrf/7eiaw0Q80+fc/N0gYMyTSbQyiQctP1Bci
hyqRAK7PtVnXXYLY//KN3Wl0vpnfyd8xNFqF1Mm7q1ZUu+7/Dx5IamLhlUhtEgwJ
V0FxwZshGr6jafUZGZUgalkARbiqZ2tJBL+eazInXPX5PGcjBD1OPZvAQvanYE/z
Y+5k9d8q90nzNsgh/FULdv3CRejOf/FDIK6LH2vx1LieKnCIfJzIvAAqO6Ha1k2W
G2VZev7tUvu7kzJShlyJ7MRGvYo58ADBhFfXVsuPUgp+0hTm3Sly5Z8lC3I1qrQP
EcOGt2ail9MSYo9bH4n2lATy8zIpGxKNuZtSOZ+rFh5aeAHXuA6xrNi8eG26eDiz
h9ZNZdgGK/hzrcBDk1j8jlpRWF43GXtd340JiK9S65GZiNrb1qbFU/80ySuotkbV
gF3ec6zI3vLEJE5tvZfOAzS2fMnb/wMOBFdOKKx3nLqJQAMJZFRJQkED6Me5gBdf
tj9OFbUwpMlZgFw4lM7Twk56W5QrcyVBJ2MTd0YcmYxAncRumLASAMzX4DQAh382
WY/7vTS13WmjPBZvhHsQr8Ms6GvnGpITmM1peDFh04D2VAFouwvnWQh5NOqMOB9l
IDmJR0WWXElBCuvVtRKSwBhPQv1yhg7EAgtdndiwR7Q6impN6EAdFiPoNM0U+TBL
X2/6bHoG2LNSK+aP5LqJGW/vt+t0qXr+aKYRoEDTycG328nBHAzaok/txrj3lvFm
/dB1CeMcW8BbRrr/B3nLq6T/obzd7+IRg4m/mLZMem91UAoILUi0R62RipKkYwq+
mh0DdmeIlWfmVQJGWNh+FOIi1Cez5CaPeSvVdrJLQ9dRxCNq1/hqjjcF9VyME/Jy
9m74z3b9aUza9zKDbHtjgmFmUr8HZ5VOD52ejNadlKzQxuJPOI13O8EZ6pvziNAC
qePCvlOFcIGZApuBvQIosDyhDM85AmKOsp5+6gxBre0jAGr8w5Kh3+DjCyCj2vle
q7yJD+FKARz0TcSDXp8bWZl9Sz8DG1yKjWv9tIk8IdR5PMpNrDl1+QpuvBAQm5mM
kgK9y+beoss+D8aMO/yIlh4DZMSwfD9kaqmOlIY0Fer5ICDgEF++p3izGzf/Kh8E
ipA/xwOV5j6DIIkwNf199grKsxWJpUVHlXP8CNnJBv8RyUA88KN6AuwmM9oIQ6rl
yqfSt+DSSrZ2q6sTs/7/BS2hBcqzIYQHInIW4RJLZNJFkzfzB82ZJxEt8zrJnGMn
yn1RyZRv6bxmtV3N/V7cRkVC0JKwcOpWjG0bTF9fGT0Ky6eO5nnEct3jySmfS2Hl
9MvVObZJk3xcNU/Hmq4qksWQul37Hwa8HTE+0ku/1e+l+CMf2LExXiXXjyL92Krr
4zrZbdsBWN+i7oWTIMMFzD7W9W+BEgdRmDTVIVP4WOqrrkMSF5veAlpHY6yAmfLS
PmYYNCbg4OYxP6L5hZrgmANcsc4PF1bqYCnxru8wt0EZLxViB3AcqoYi8ivZgoPW
0NVx7Jixg0I4sElpjc4aJudFWTv6FCESDZ2Z1UWbkXrHXogu0LdVxY0OqHJbFlG6
969stbedlEMan/kCgIWaruHgpl//gBVH732vke9kx/T2+RvTsVUvXinLO3Zwf+kd
Wla3m+iZ0tyQdruNkHPhd01KdcM+hJyV9bF8faSG9lsm646AwDEa0Y/lbOwLCrrO
4YFbzBmZhSP27tXVbLLvUsJVctaDa3juCTtmAlEjU0Hd6/cVjbr2Kng5n8weqxjm
s1EBNzGOik+SDtWiVbB0tD9lN9krPln/jA6HxpIKv/4nD/PfbfNDBhMhpr9o6/hX
HP4dYse/r0IeVHStJDg7lsc/tTr4UXiqDAN3VBzsjxSICAC/cvCTxFPTBZUqNUR2
aFlnrEj3iStgN4h6xEjwMP/GHezuzX4a38F/wb3342WQ0BT2d4o1+MJ4ocnO4IFo
Nt921DlSIP+2WZyA6zLDMWmklATpLnjPe8ROr3jA3/I4+Bkh8/NZS28YdPVAKSj8
grcBIQGfeunokFrK0r5g3NcxhK7UP/pQkbYkwcwgfD2Oq1My2xNcD3xXoLwY2c1D
0EwJOswdD04lV4wznPG0Hip3A+RjUaE38ufkk9/O6udaBrH5byuEKRBviAMzMfsn
Xwr58OQX8HN/QQAGVZcJHHZVe99qAihznKnOaJ/oYXDaOpc3at4H1vNnbEc77Svl
RpZjjGTLIu7NJ3qvtEHYIUR0n/SYV8qoAj2Q3/C+jlYdvIqO/EroFYNMSt9U8q5b
CWQNqpSO/hc9P1K6wvV4tHaVoxhqCH8Jep5fiY0fhM0C1pEJLC/49cp+Sp/JooH1
6jEy7MReevAkgW1l0agz87IkksGs5NsgQE3CMoy1sgmTpaJoJTJHd5ym2E+mmdkv
HTTjVq0s5R7I0k4ZHuiofp4YZgIPP6EFiiGHOCKiW0/NpXh7vGOxKiw3nkEd1kXr
3vOK3Vts4JyVRZgfuI6/tJtVsmqr8qAvJKZXzgAcKPwtt7IzVO4XcKncCxlHgdAi
fzP5CEqTmKJLcAI2wq0MRYp3ObvIKjsRAr1JhfofjQNmEiWZsyAVvLiMk8Uhe5Z7
jvC4jZXnAQUSVTQBMxbJqY1LitwFdj8r6b7GmbO8PaCpe6ShxmW4RMPTzNA1o8+L
A1C73nSrWAzgjCavaxLMfkFZ5slPizdMICifegVnONf8zxXXJWTOIaZjmRU5xgYf
QNAQTZimw7q4EvlZ8kAP2v1miSsd26QkCqVkoIPKiB9uW2DcW43rl/Yh6SEGyWmr
Iqhc168A6dNIhXSwG7M30z+NlN7/Rt6bsM5QcCMvCeuMAoEq81cMVhjN2xvly+IA
P7yp7hqz1n6XtKCAe3VXRUCqFXYHzJ/URn4ZPfOwA2sjUnKz5ZGfz8YDRCwXjjAH
9axrQqc+wwkqaGLAap4hJx/ERZGwzAwuBQWQTcg9PMVXk0In1WS4GqNjT7wgG/vM
0JUoMhCHZXBmfO/zlmPtXRZWLn5pKfs0+YwquQvOvL8mfEekPh76IiB82RyopwRM
GQzJP74R6hY6383924jszTiaSSSKGFTCXXCDgxdl1+Wc5rx8PpTWyNthY3W3KZXH
jAMKYBDNlzzMV+6yUOhPsb0hSSoVtb6Nq0Nfyr6JSVS9trf9ObGIO98W9T4hfj8u
i5VuGESt86y16bjqS/L2pyThrpo9+jgL4kDqFGpaWJb058QzGZRnepROPjyddBg1
6WuM7roCuWTnk8nejVZKupbLNgDZyWe+spljXFb5rjh0i9VcQ8gQnADBozgZphcq
4oQglSjlDKeMhWmjRK7EfaJ+uhhk99EN8uwSZJy3G05ZHzOxHWDVJg8u5i/CQO5C
7ZhnDCcHu2flWSXrJcvCn/BXJ5OCs6KZE3kp0FtEA59eHrnDQQ0n1itUwoJmpmIX
MuY+kZHgpuHXD2RxK07DYwaQUyg3Vtubz64GDRln+wUw/cM2kNJIUIZn4zHIRUOL
53yQZ9QAvYqTtmYOO5qsuLuZ6g19/Y8hMcZCrOPgBFZMCDXvIlYEhMGZjLX3th7Q
6goiHCQmgVazBG682DA4Z3pdpiWYCftGJgSs/v0IgYqO0/7Z3A2jqdzshIkMmdpJ
1WrYpeAzNAvLA0fGXkH8Er98GjPluMsHGP6lh+VAGdVnABxU8O3Z7DQOvYawp9pz
EuacX6EyplYufqwWOYC4M44KgF5vwicNGi0Fp1Wsi4rZ0wIk577nvMxbmKCpXI8L
aJiBWdueGKfV3FQ9rBnrGj04j+CoHaX3glJ++1QIvEkzICY88GwLE7mqIFUcNihN
UnByQnF8zvaTI0VIwQ2GaWZmUtKN3oH2HUw/OO2X2M/5zhNjOpo5y0oeeIMJuqOj
TwlrDdeYstF+CUCgM0Dm7xE551fxyX6GIin7UPftUS4Ml8bCm25PqXsErklB1Opn
SVVST4fnljI+5X4AdzxCA1mjtz+5wfaw7P7p9hDLV5QkRY88HrcjbOnxFEJlP1w/
Ox1xDy/Hz1jb3MySRLwLsMzvxxahYrfml8w3t6jY0DJWUC0eDFLefuHqOL/gkByX
BM55Hk9nFjZuGB6LkNT9Omsq9tN43lw/ouMaXgKm2OtFaw4UwH8QUv/o7n3E4S8W
fggBjkDh/S30bzdTKZHZyMg/CyRMDnmAeO1X+lGiUzxqUc+//sBKZVSieMJ2TFhW
7uI076De5EpKD480ec9AiXAc8qc/V1cQl63S+8tqYNU7e3unl08fMEtBPTJTde20
5qyGCPl4a53mU1Rllm/qrj1VKOL9a7Ihfts+lAWKHSQI6HVLQ4kwYiTcTi56OO4h
9LXXCG706+VZHh1uCyYcE5upHPOfN7x/Eu1xObJkHryiWP0R09YRSlW20LyswOGo
OKV0hCuxwM6ZiJdYfLPQ/l24k0ktkU5eI7f3M5yPiv70NjPfzTu9zMbp81idgSHz
675SIiq7PL1GSc40QvWpWImDGPPrZD8wQdo1HqyrYbl7wFDI8/fHWRxQVVfNTaWl
jXOWAY8xTkfQy5QRaLerxoj1dUifzBNKvBOEFqMUSTHc7a7HPAgDgPeJnIhJcAec
wo6GCYMnA1JvoyonIy+nUfcG8Xq5ePFnTSPmtceupAXtDu1tbswAJiiLSAoQfgy1
sHOU2ozteNE4D5sG+rFrvXUTxqSzleefXrbZIrQ0MuM+9WB2TaA58TQMkg1TD188
9dnLH0bRidJoE1uAm8cIEncr6Euo7llGcNVKWIUBgiNxjoVy+2t0Cxu8pzmsxPOv
FoRnCtliaS2+7ZRYB7nAZh5IBMMn2LXjTpkZUkez/6EWpVy5U5OdZAz4oZauPFTo
KlI/uWqLGIkDNDRoaPc7XcE2+2gox9CNlL/0eK00HNrM9vyKtmrNeHBMB+aDatO6
Ub+LVpWp4dQ3XvaqWjOQJ/cTk6pbECySQ+t/iJyDyv284z9fM/V7GfHAJ93TlYke
ywrr6/0wz3Z9IfP9P9saUbV2Gr886dtW/YK0mBCh5ejAhYj6X7Vji5p/WxtaeLLR
gbzwOVEssfc1BW8G4VeWo2Ip9GBHfHbR+AdB756p/EvGmTqoRxzbsqi0e8cgiHQI
30O4GSeQbXHQobTj5WVIt39lr49ZJkScVRTKhtb1Hw/X/ZwRPtWsJiInwvwnLMT/
usa4EnzHkd2/lacYlBV+9AHGpqKCMRSsSAY2KwCB6IDB9ciGcw5dx7Fv07/FgBZJ
x1u6gc/smprn37Y6+sVHZx145c9Ir+U92R3MRp2ZfyUAeZOnAQmtUAArIyRiKX9G
YZbWPoI9NC789tXjS2Rxm+z95Th5CpiUsGbpuIp/pybAJXQZXqihzkrnQLPxAVmN
XSqxHlNgMLYOa34Ln5ZK5foipSYiIIIQzKA6apeYdzTlB8aQb1BvOGsG3nXpzRk3
EwQvjcmkJNyVy+0FnH3NlkXr8zfffTIqcvRhk8SID+y3bYzvya8/GvyRPIt5C/+j
OpbUfA+tF8LPMKkIvOWkM54rV5w4tzqtzc4lGZygF5I7KHVxX7UBnkHX3dJTJPOh
gWmOeYjDzXLEQUa/zxZB17N3MWBFKP4G8k1nH8yJXpIkKQy3ndq+5wSzvaVzbyoq
LqsMunonrs4FVsc2zz3Xnzos/oTQ6dseX2zWGQMsOt6XpXrxv+QNNV9fGc5aAKya
CG5pOeXELt81KN7VyEdjDMvajd4BpoOhHwSou2qri22Dt6rk6WlL1MuQw9cLN9nd
VVGl+TTeZ4ClJsEL61rHZSIroZzLEIwyT3cLT7tz0krQ3Qy1EF3DwKa6xMwXwzJp
L4Ida9/4qqfB/b5lccTW9E6ApoIDdAD6ZCvULdJVu/w/moW/4ivClBbTbCAZeCHx
AtyEICf2J6MsJSXPJAtU0fYV7LpaW7GIsYqMKL9JzCiw5eYRxE9sKswP/lJ+pLcD
vitSVl/DEgjs0/y5uKDZ8Fhkq5s6W5xrGI4CyQ7Ecp7KIwvSZ8K5Y7cDWkTIsUC3
jr8SLv/M50zLscfoRsJimVlof9dVWEU0JooHGPi+g83i+WdidlutNGKiu2JFV9sA
0mPSleYmoZA/xk0LWQzp8x8VMP+kyS/OZg6HrE3Ar3sJcYZfNtBMMl17Z1SOTVxU
H0qMBgSoc3vVqA9ZwVzUJpc0bgptWag4fTT8gK2Wkzi0qXpS4F7szj6pRFo+4VBR
bTDm5EFalp5VvbzRPKBBqh8gfUXbpFNvkT7Xm+yPBRzV1uG2tr+VkWaBNyW4vh0D
IuZPvNcA9dOo7MTjcYHP3UP3kFKNowagmT2o5qvDuvA6kFm7mSN0EEFRiE71Ll6t
LseQ7gsVv5BCKnpMoFc7T/09oPuu5k1VOm7XEFoVx9ea2gD2HYvkHoFaQrTvXGvC
6W9bLEOy/ZU++Hcsfxxg+I7nVAp6uUWR3OxuUEhpQ5Y8EED7ogFW+UFDh8i6WM9c
2/B+CYqWZpeJX27+fGmvBLxtGf28fd2G9rciC5eYD/zET1xeibr+iYaiHn2+o1To
E6HSRd+RBkk9clq/ZhOQ0Ja8yT+Quiw+EuNIPAkiH0AzSSFfow6UrGDU4xln8CgU
UxPC/udL2ZULDVlMKO3d2rYVJJvZ8dXaQ8oV3emOzSWPxzfHNaHtvcTD2lfn6/fG
fIlxcF/KghzJ0i0FrC1JJe8+zTTxNcaTqCS/+F90OzA/oEyA6zK5xY1Q54j1p/ER
13ywP+BFLPnR1GWwgmrKtBPY5N95UafDcdgBl6zF4d/NIIu42NQu2UrkXPlt7mrX
M5vkkTuORpJbNms1ZgPLK3f4OHE4hmmxKyfTrYkYo+CSKSyXXHAmzVt13f8+o3yn
7wgWGjJzoOBPkc0BNLTvyxuuw1LKal1l1VTxNsu41kdsjfM96FbCNb3Zg80W3i9Y
//gG68v5oMI92fOIRNagN9MhhRggc7F2bZsxtFqUgS7PpshDRuEjB9Nw4AOFoo87
y6MccCUPD/Nq7hVNgtTiCL6joEGqIIja6gmYhQqx4bS6KlL94kL0293A9N3v8CkH
DBJtmDxgKXWhl8eYqIyiTrvna0xZBoFeahjE4RuGMA0M46LPNbm+24wBMMbXdfkN
Lbpi+9SvZsKvzk8u/1MRRJzEk77bTlLc3R/CjA/+F7tAQs2PXzgpsj3ot82FnjxV
zOErNdH+PEJUmDrtEtqDrnRxtZlJfPuMPrvSLtf0ngy4EhgwNvn7sLlr2v2Xr+l1
eUDEvG5X/4mgbDZ72yLEw4ORuLXC0P4CyGs0v6AWL0UYPpQN3GP0Dg4Up7QYt2Xh
dH5XB6c6hd0+7afK98bseU5F/hM2XTnX+9DZaV5TF0UnlblP68Xs3Sh7+Kole5Dw
qXFqqHmkpgki3cqxDcDKtr2LkHVssgaAnuunpyjB+98a8FchgEHqB9Mu6CeqUYSF
f5W1dtY/8uxe5YteM5dnq8J3MGZHImld9VHUX9YEooHM8y1N67iBaLd/d3NB6Kcv
urWJpibILKKKW6WgGZ9O3WdEoEGRN/2r3wLIiwI/XYCIN3K50F17uKuLzZ0P8kvn
SfUj835hY+kjfGmfrCDwsOy2iwretxA97vYgVcLYltzBDkEeFr/Ac2+U3L20KIxB
sf7riMwhDhjc5ObgLkZ71rLOstC6DYZaUORe5T/jzBwFjTIgUhEbT6tyxl4768cq
FtHu9LJpwuY7t/7kpgpiV8TgIKWVlqB2jLQ5P5YU4SsbCzesQRvJABGtl6wUXlFQ
NjZUX+Tq/SJJtT4aAxsmfiY6Xu78fRRse7mf5rdJi+heKSmWnPBQsfZYgoagMFd7
izZirAdJpew/4wx/C7gddr3PbyagyfAWq7tEPUBoDKlRr/axtYvw7iEjoKVIhcXD
pVQNuY6igGNPU4A84vkZk/uVipSdXalpu+v1eg9gF49BXbml/uTzS6C0aVyNWP3H
PfbgM54u3ogK314Lij4r+ZWXNclVeSmHJpyAHu+nxZ3RhlsNUWlY4wt9bhP2ylsM
6hSZdNaPrviy9ARRqjS+6SUM4b/UqE/GlarKUErYi01wIxpscaPil+4d7iYnBjHd
aY5kbUtd1740BPyayDM9sWxDZrFk95SadCkB2FwFow5ZVeNJJKPI2Ziwcsw9m0hr
zcGE4w90fFNkTyPyzksclPZGGwBBT0qknuLTu72NifbpHGxg1tl+JOQkc6fYAHcZ
qXCrjRvSlgjDLEMHJJwBXC6KPB0MKGT8qxGZIjBJxQoyNjoAFu6TdkPejUUg+ft/
AcmIi7799Y6/vhRzPEYf8sY8SJcxBSmeICNR2UpTKQ5YWJ3ivuK4WIJVfQp8wpcj
2jASM0RuMFvC5n3nVs5DKCDirxWxYkiFTWrmW5WNGAY63+g39uML9W4YDZwIIE2h
I4y0TsHsh8++h2DfG2X2KlR78OIZEc3Sxx8Rkb6OVJzLdcThS629zh+5dhD07HLi
ivnO+whMZCo6cYSaSogxJj7tVkMo0O4w6fiAi+kvnwrmsXT+N8zZEKxW44Ahmiif
xNKMYMavQPgS8dcT8knOR8kihhfDDcRanCpjc25gA9pv4gwQd3Vsfrg8l/iH6Rcg
CNa2a50mohh1FTOjph3opLub8DXDqur9Z4Y+HTBN7suN7Nott1sg63ZsihS+FAJk
cET+68hUHf++2hYSwx9eCXIAXFpgrdPRQRcMvuNmUtuR3UM4LJ2rvAt0jFLBVQ1U
eo04Jl27ZoQmtMZcUcuU40DLnY2hupiQslo6axcfvPNWWn/nzvANLon/ZYTuPMgP
rMltfLEvfVKcJ7tkj0hcDMKRNAbT5IsBfOh62Res831sRmgAzF1FM0YRvA15tltl
NK/rcklmrgnsujfYRGRpCV9BU1/57woJMwQ9JBgW/lTtxsjsy9TkK4L4UNMHnygT
2BEgYOUnpdmtoVCgW3gglrveYgy9wUjr9UvdTRoSdmKrvUHRe9rr4DFmJlHxiJE8
VrwcPfi8jXHH18wuoKSoTqjANP18XXC+nSlyixgmbkAbyiaQg4SOmoDeUuqqgUqL
OsleG8cU7VM4BClXIUoUCFYXdOOkGV2XHyJXrrvVNx8EfHZ1alX/woPUe+Egpukb
kXBPZ4kNJMyjTPtz2bGKiSYwBfVPIpLRu5jxOEdC8zKBsUv4XkSMXBKtoRWhcS98
TEVOTFlRjayEkAr61KMkLXX4RPGu5ACW74l+0d+8TE/uMy8G3b28FxTSeCF0fRu+
zp84udj2sYOLvTSp5NY8N75uwfmJenHGhf8N6hHeXs0XKI4z78yiBHvXNuohqS2c
XJfrCecKzZ0fAK4g2mewmBUXYTZIJFK36gjYDh4+iLDhE39d5um6VyWQ7VJx1cs2
vzG+HraPFsLM4ZVRmetU/+grFmGku98noQZPmyWUsrWoyn+bK7R9NKJkLCbdaKKH
bx3wqHX1V2SYjlPVD8tLO6E5tZErEKl69n7FGA0CrLYJOrB8E7TPDpKsNwrFxQNz
cD2BK4wuD/AJEhaGudTy1rKe3Ibz4BPrN/BUPN49oPZVPSsTFjBl2IP/YpSeL53Q
7RCve1UEmcgYJ/BI1imYLe2T7amTTEeqTzQ7YlRDZuWeX0io3618nCXCKLonoavN
6UmtRYh39oi+7q1xf/h36OHVyL3KGQ/RqY7/vn22deMIIocMhMCmgsD4pG+5o4Sw
p6+EAMPAgsfkoJSTH2tf22RFsp6nlLb5WEdsXsd4hQBqiXrlX29BNYA/NuZjrdOZ
sjz86x8M/GfNEr+ntuE1nIwEQvE/dp/jcBttNHdIxeLkO/lGHQHg3qvqubso15Mp
EUFobU3eDfZL2/7giDo7gDL4jTEXMBlUDG2CXGqsQ4DKBXWa/zUBVBrcI1MuVG9m
m+6FVCXFoNb1+H4rtl9Vtg+dOJhDirt3jKIP0H3vaxzI16E9vzJ3oNdysE34a6iO
NEtpzAA4UIEaZdrdUkvBEmAvbSfQLZNsH6WsfDOzorGHdTIExNcYaY9g+mbrT4ch
5G/NuzG4oeU5uNNAy9n1lTPKFwMh8IN3GJ9d9Xh6/vzZA5kantxeHMQ5pC07Vs6L
oInUjSKmOoHqSayX9HJm85OCd5QqqWyogRSc5wszn0AidPk4OqDIBJlYCXCGGBWw
i1dsTtr22kTvSLYxT59JTiTBEev+EzK0eldmLFzE2eAoTo98UdNYDGiCERS4tD6d
4Xyz9KbpZ/Qzh1Ud/HaaHHOAFD8u0vAQJnqo85xSJPQZnmkK2bpR1lbHNDKSievC
VCMsJyyBP/BXZ2APXyLWyEB1eT1oecGLnIgY0UqYAR+A5B89QNo2VVvJ8gTZSxSQ
O9UtyVzb/rFJ0Kf/bYS0mlayFVgrZ0v0PKcWtxgS5eQ4yHNBGnf7qXqp4mmkH6c6
dOsLprdgli6tfZQYcoyI8CMe3kxufYG/rAWqtsk4kT05G93c5O71NQQkjC7CyRZU
gQ/uQHBbLVpmoSFEUyX0PV8eWnFV/3CCBN/QCG7HWZe7V2ljjbthnjetWB0AOri0
x8TGm6XOm4PKCuZdshCc1kugAoFZP5qPko8g4wdKtxQSulVqhRtnhfPL3tPQplpi
lnwyXtPeMXhI8qRGCw55lpriGRalINH03ylMUBPsHAR9wyKBNayYRLwZVadXGSZO
GVFJVKvBkosTdpgiJ+4VockA5Rb/0w3uIP1lGNE1DOhMqnYgGbJD+GUClBPnOm3Y
ziaXf4xolJWXaYUaHfjQfDFeqXqFZjB7N94Cinh4LkQeUfLtwFZDzT5bf9Cywx5Z
Fk8GnjW76zOYVPW9QthZEn5jb/tnHwNBmzoWj7umulnfgUe5AMFDSGvjPPjgRiZK
LeoWhgUMlG582dMo2RNfT2X6LFpcQHFku3h9WbvJG+Yq4MdtLGVJvJVXuiAK36at
7nL4BnLzGjLlRLq2IndDocDw2gJLM0fo4B1CG3JehuBUqWg2kHe15B9grH2dXtoi
Ahhc8r+HpsMsQ9dHMrxkF+qSqYff7fX4HPVUn2zMKl8yb+tPQamztbyrCKx8dhoF
1budf+ewe7ukAo505Wlw52lE4S2aqrIoPZDDVUhGtRI1jdTI3236o1CBUX8xadaK
B7pg1SKX3WVt5OjP2C1NXmJyV3HD8A97WTYLO1Q6LPfdt47aGtS0iFacdrEB7v24
IAXwU4w9ZLz8pELj1QTJELDX1UXRp/Zo5qFoIRjfcs3rgjmz1XtqBIkHpdOK+EWs
2mJZXRwtZ54Tjk/5fyp3fKkt1/A/7cm13fHIaKVgwZaaKj2IOihYJx+7bdrdlRXf
ENoE6PwcL55/80HuJJMTAPuoyFw3J5K9JB1hIsYFNYMZUs0Ax292Cmi8+MDH0au2
t+eTWe9CQBpNHByXbrmg6m/Ca6JEf2JOX2TguYLPzCr9/31IlAndX8MN66s0FSxj
Feq34gRpLwF7GauumqJ8wnGz8mgb9KxBZolWEoOpw/qan/28qSMcutv/SEOL5l5R
Tx2uItr4C2wtn5rm2zU4q0Ofu7KqbQY3dZEnLHKmqKiscMqCuc5rnmk47E6Ao++d
kRyZBOkp5lQfrpNh87EkEhpBfNqJpgkY0sL0x7K3byM8pn+Id9nah5jwIQc5V8Uj
I+GXVTsWcdFO4WQfml1QmMaYDMUpox5ZTRWTKpZvH8IuxEj9KrG2BUspG+38Nte7
FrfY9xPFjYxI5bdas+dIEM1QqQNcAcJsbOD070Ne99fGx5IJttJsPP1oDJCrXNGX
Cd94nA0joBzMuU8iSw5g7IydIgeCyGXZ1Z4gsljFNCt1kICcfyu9qCNkNOzm91+p
R5AXqufupCh0FRBdps+wsCEh+CMgMocvB+VOea81tfxFFcHxJBlWiUpLC+GqbG7h
lp9N0R3OttV3TbKRrbgv+ri0BGeTC/kfSZ46B13/OO38Ui6lNOXhNlZ+P5IhV6bW
lUYl6bjYHRG72tB9mzlktBFR5d2/4x/hz1A5ozMDxOHROwrzZWrODZK4aZOztVJd
3pBged6KOvjdB03D1SkUqSTOZ8RnKgzgJfQmwPlRIhnpcM5P5YmcXiO280lnaE/u
EyBbnUfBXCvIkwVS5nIG4xBwATTTaO6rOAIFE0yP/9cLrXnVgTXfEWEBLUSoGdH7
pWz8RpYQPOOZ0JQdbNLBaa/3ceUvgfsag3lIuKcMnB7PzGVnKrN7zeCy+QNEUoEZ
xN+k2c6SoTYXy/zwhLBrnVO39lZtfBrJFxaUSwDydXtxpXZF91vS9Tstu9NorzeZ
3O1k87cwcLWvAabt+zk+fU6ujPZ66C6H18dKdhBPogofR5uHVpnwJ4j0ktvoqkE4
kGzCgv/VWwLwoYin2GnKjuHHHfvHUfYWZM/1RcqDOAumze9mE1W6tYbUb2m5Pq85
Uaa7HgNmIrQckKx/mBTwIVTZ4eEZhBRF1RIdfW5Vbbb+sotd7oy3AwK6czhICpGj
gcDX7pVKLz2qquxFncSmZJhXxq+EoK1ci86XAdIcg/+YWBcGNjW9Ouy4k/oDBmz6
N2KpY/EUzLGiWaPXEaV/bnxg0eqaFSMy3ErdGgz0+MRAE+V1s9urlb1vmnUqwCgZ
0VaooaFsK9L3cPGCh70tYKKK5s9gQE++QfBoot2v2yHpYBn1dpLNkw0OUm8SriQF
gaAfbjvxzWuO1Y893gEMzH68EzXb5mZyj17D7YTlNeuKN8dcSUzIHm0UDKl9vRzJ
QT8Dh6Yqeay6BNIHVUo6V8KcPzxFcl+SwrO3nXjQDu/aJqh+v2mF6u7CIR5UZei0
9bN4tSK9ACkme911XKk8BVA2k1HpbKgSwk6dIA4Vbj1EtShqL25WoDh4TXD2YsnY
rxj+0HRy5BTdGw6V0QeCwnaJiH60WQ6F8vGkFi1E6pVHLnBKO5+5lQiU8NvAUwv/
NBzhpsJ+/fI+J5HcJ7BBXx/1udlyOOy2uOZ4TOcGbDXufCv3aVVP55NaJ5GeI3/J
wGDLmz/kFiaDp/8r2IWUNzzZhVMnyJEcjv2E90BWWdBPwcQsIndDKu1dxQCSS3G7
8zcBETGh5UGw4mFjuxl0JeFvVPCoiCkfRhWpPe3LL/s+GhVXTwdwYPn6L8fJZv47
91c1cWreypLJfzN2AITMpT42SDM+Rf1+n/nifg/BxBv1ueqWKVYbXBS8wl1OBwnw
hnsEvvBLNdjfIzN7nlXBHE7WVqFLUD+LVOEnJGakcOMSS+lSvDBJ8+2XNtKm1qer
b+PBEOn6bltGTusclpAZe0gnawwQR2TZGzGw1hmZEnEmRpkgEloCMqtar99cYRL7
BCaTbL7SuQadfqgyvOPq3Nr/CPN3Msz/zfdmGiSvUM+3hDFS4oNKklVDlbVdBZgO
SE7EbvWRtzJtlXzFJtC7XWUtSnjTzEEeEnI0mUPf28EpA7PguJhIZTY2PXRekRmf
sL9640htz3fNjWPmZsyu13QFEbl77VZoptC2GkP4Y4l7xVtpdA0ijTR1GEqe6Qxv
NMWzGIo2B8CkZWmU8BSm1omMFHRfp+1o5Vz4u5Uqqosv4bp17bsPRSkTxTGPeVIt
AD+oa92J5ox0pIdSd2VMRFlsUtX8jPsE999hZq1w0WJiL2SveaauRCAYsPTIPqKe
nBslkC/72WAuWEj3/YbKy+qMQXIXAAn9qL2cwXOFLES2p4S5mGiFfkxeiF13RuB2
UfpEDQaw4ovclcfqsbpSWQBnbbqGc5B9hMZbvDS4Ke/zk2HrFhjYnm4pCYCknmyR
DQaQGoB+r0gmimY3yb4IxKy0TGADEgfL4tVttYsCcvj6jdXP+cuJGPy4TeNbwR9v
zezDqKp7q/92vd1+Ie9uGtbJEkwXQb4LlCc6FR4hm+qpkS0ayt+DCWlXFCHfGyyW
/kcCZmUkEslq6yv7kt1TFgjL4YxJz6RwBW3PYUpIriwHp0+uX3ZTDhAcG6MN5REY
lDX/P3sV0a9Q0Lf2MfjfdH6UP5t1Y8JHoisqBiJeCerWYXZnaFG/RJer3tMLLwIY
N0BSOb1h4ZpFTA9tG7mszFOKrY/G1Seh71FbX1eDGmKzG26c3FV7pkkL6a9+WBgu
BFNS32jOWQ/z1ZFoSJrk8ZTZ6TU/Y/Zwbv9QjBjMhFb6EKK+csn4FawTEg9FwUnn
PrfUnzTH0U1MEnYu1t7N0Kw7U2Hm8Ly1oSpBvt1rgmOYhPgA1/W8a1x8p1BJA6fH
2uSxP5uccgukQhHe6qwqRh3axInc5/znZAOBfWrkuvGeeXws9SJgy1t8PXe1I9TK
ABnIiQ5/he4sM7VBVnPR0VJYLhYPz7sp2r24v9beMVOG2uRKyjw1yYaf6LhQV/lj
2Wfq08DP7YxeSIsyrkrVKoov2J0e6HdrbHzxgIhgmkmGk2CF+BIS0JPJ7IMnoiM4
g3qVcwdmKHsAyeYdrkgtQ1VMJ759D/EVfDk7UF/B78f0rICu6QN4F0lfZbsR+Mcq
HO65HkLu6jxVyI0PsVOE7/dwdg4ze4tqkiEI2poAc092nVwg4R8Rv0WWIRlxo3Mq
ccPQxQ67EZxstgfYlPHj7ICFUr6YyeGP3+CPr9TiBnVQG/rQuqNmdODwtgmrPUbG
D2fQZzlco1atlf9OgcRDv1DuEb5fz93ORAiWEjDR67MeSshA06XSDotp55jEGotM
VU9Hgp/kNW8Zptf+dyzh/5Xj/06kLuos/hckIuDqsWtTwMVMObv3ggQs9WLWwmGh
m6uZwaOdceKB36C4qse6z4HtYRf1SwS3NY7SAmNCbQp3HOrWnmCy34UeaPkkqgpb
cjIdBoPe3KMJc67owqdGkmMNcvZcySNjCwflzFTnQ9/X/YSfN8tkE7LtjsBLxgS/
eEY2tgq5c3356zAhZw8vRv89c0z1zlwWJC8q2qg1NOYZXjkM8/8577mhuyeqeUzJ
3GT5dJGuDMbbEpodGGgP0+YXoiX4JwrRuMMi6MOog5oSOOUzAVyckEEtl9gGhazd
mYMhYvs1k8LCLFbxzdUkvZ74TogDrDXZJbx6JyDcwIyMspudLjCyGXmZ7iNzLWxU
NCUakzKBP0HAbnPdmh+bqe4Z4f9HydH0zjLviijTJKcTTc/9sCnOp3sLPLjXDllY
o9+HNW+k2qq+wYoGLioXsjd2UwWmvtMRvSaSloaqsZlpMuFlEw/gkZeCBQdGLVVB
167iaj3teBEY1bQ+2Kf/CWIGaj1XKHmSO3yn1ys81H7utCdvJh/7kY6hZ/0AYfAY
2Jw8DMMNguQ8XbM1PiFLkAXXInxJGfJvRwjbjriO7Fl+ZdWkGARoK+S7OH2GpOxj
7PLOydJyumn2y9dVcSMxhiKl2IsZs1fR3qjV45P24s5nrrgenPU+FBImQxC+U4T+
aY0oriURnA6ng6z6N4qipj3RnKz/Jg5fQb29zqH8wlgbTCid2SfSXno2DBjtvpGX
KxrzYWbTVfwIFjbhNaHsOjebJiqFKwFoQwZHGKshtYhnYUpp48YS/W936CDrJbmb
ovgecDr4Lz+SX4bg3ucos5xKs62Wz/y05/NsxD7s0ln2gDRVA9Kjle7M7zz2zb1u
z5ZOU1J4hxjetNM4URVycXkCkcn6vnm3UyssyA5UXbMEt1bSDZY4rI7cy9eTMqxt
sWfAoPdmGAQX0apgT6WJh/ta1oelnIc4WJBDdJ4eTNwkECx9UyYfUpeOKO+en1Pw
OkAiLByDxc9P+et8RNwZWpKNAB7genlRIba2q3sEV8yVk4F5Ykl888mAOnmQ5Jm5
PLbRT3H97P7nHfJ4/jxUiiKOvgZ2aey2woTST5BOKcqP3jvc0NrG2YUz1D9Ja2Dm
uZL1KP4Nhmj9UYIQHaaC87E+kQkS8BbdcpB1UDQeB+B/wdMP7YK5qqIOJoJ0YZGK
emVzimvU3H4YCxrwAhLt6gJz05tGTdrg3MEupbkY0rK3bBXTrCSsxBSdqyTRGC77
/LTgwEgk/K0V9pIYjYnWoz2+gCey2b6BYga7K4AH9FMRDsnT87YhSe2mkGXhR5Hh
mdoTEEBkG+uvevRjJ7ELMN5xutuULNtE5MmP/jOydy3T8b8QMoSgK8M4ksUStbKV
A+HXsP5YLGrRq/3P/lodNj3ZUzDMxtVGUwTKDrLkeZ+EIuXzEAeJuMOrg1edczQ9
sfra4VmqxnQdO2XBbUTE/i6xJrPwjsc3sib2cit5AbpRKf3r7+iTRa8ssAWNTkvL
cAlt91F8CeGnJR279hqpW1WUp1/O6hcBvtj98rH/fYVHd+qbW1gZjlR589yHw6Yx
mX/FtQFPoaJG9iMjzV33Gsh4vVF7lZTUi+lZs92F2RXl+MOXKpsOyWjeOkTjYfyj
HU4s1wz5B04nneOjh//pHHFDTh2rIyYlGd1aqT2ktQsvS63Yl1eBoSiX0msqjqog
PhHJ1NMn987ZNjQrQQBWStPZ6Lygp86nShh0QXxCkvG9TQK0BTd21xEzNO4qdshf
laScoHxQ9XF1lM4W7sljMlv542jlQrfFvreN3coHR+saC7u88uvGTHNqnL2H7xLr
PGEdrWKeTb9NYW72vi46BvKIx5cENeaEnBe8kPJ1yWMqWVc8L0/WcKpVTEoespFo
NxzHnRMpPzUiX55+utPv13YmzcQ2N3bGVk4WWbvzy7MbS/pyIcbhO7GgMaCOC9aD
h3JP9yNz/rJv9ARScHW90rk+mHZHxOb0RkhLI0E7nQsMmt/sYKNlLVhEZcVJjUvU
WFMN118L+QCDnIHce44o6oUNMDZPV4hijfXlj8utKBNbg9C+GlB3y4UieSrxEuAt
Q3X3bqxM7v7ehXIvgkuid2oVEZH0gYKFgR+o+gvKWT82YqMFWBVcv4WcuJ+Sg9FK
uUY0G0BbGXggow7b4fWk9tIvwOMKyq2mXAZK8Ojj2ZRvpUDfi+tdrzH6nHg3gAeA
MrGD6PvZNO4PSvFoeIRcmPxUaFP7sFar4Y5s5WiC4CyAb3DwRkRTWRKKIUIDpNrS
cAR5TA3mTYEJDc4wzoVrFMGw3NkU1GimVXqTN5/cyoYvYXXXdF5uW59stzSZYszi
I6eIK7QnYUOe2PtoRJ8RmdnTXcokkM312NatltQijFVz452dV7JmdJ+lo3/omJe3
zi38q/vLYf/LvMqQWgbjN2ND/HKs9v8MEczSt1uPP9YebMPuTpF0i6td0sdNreBO
jGQpyDgu9NarTz6FgNB5LGq7+otX2LQeut5Q8QBdCgaZ6wCKfyFievdWsgx8o9dk
qCZ7IPYKPcOWEmxH/mVlLmm4QB7wZEYYxqBWmpSjauCSCWE5qnq9ff3ourRXtA0b
ugZfiLyAoauyn2pmmM08IggVl5Oj5QkOS/fme35oWE9jZ81LDNrBXk/zvaL4jPlB
lFf4evvm4kqg3qLq0udO5uv0tbNDpHXwOMZamx5mm+OmB71cStowPM9TtAIv+U+7
5q3sV+/ZBfHkZIo+ADfGMurWEJVPSPqdtpvQhogrxfplL6+xAlk3GlgvXcndlq8a
tI4uNht59THNyDXiy6tefw8PqfuvY1yicOVSuHlINEdEG97relh6YLvpUcxKog59
y4iJyZjxqfyWwy2rrIH2roaTRPy4MABi7I4FEhhNwVHLRppYQNaoZTosdrbtj5t4
QGmm54BxNvCqwPysc/ywikHincpYxCztBOBkMMBjJyryu7Z2U7ayDxmySP/NMTmw
cCTOdzhQjYgf4pAAGSrh9KkwaluZCEtbO0at0uuNR3VhE+bd+91JVZpDzStvYb8h
VkKMFTI6J4mOU9Ca/5eTSsbf9IKPIdU2TuFs/ROsHZVGz9S+BqR8tXnG1hGkS+k6
6n2g7JLAtetwyNaQ1EOs0y71VzwOn1gVwyvSPSsc0RqF0LV3a7JVuHdIrl0M6DCB
NUP+4qyfbibZFXwrz8u/eXLMifpG/txC4Un+ZS396KvBLnc4uP8QSIs8qtyq8znx
z6aifCOZib3loo1R9X7NF164Owu7XeKBzNQ/l+46eVTh3PHfOnwfmLs5YktP01Z5
hg+txkLi5w/e7FXroOgLHa+qcc3x0i+5hOiaA/ELY0dIm/n15zFfltE24HJMsefQ
tCWzhls1epkluHxaAzXcfWoCShkW+ehn8FPW3GmVdKpsEC+4dqXFV3AD52exvnyW
jSjilBlaMSU9oebwPlnhjSm9bZ8GZYUIYQS1uRuM1H70fR2hVbw1fR//LlofhXWM
da1wH7vWVC2Xu7RAB/kknf0U9NxDcMINc5OhYrTNeyRB1yQrE9YRHDRzcNpmVhTH
fYZSUn2wCzDxfuZQuMmhUj41ifXH9aS+nAeEryJm9VxGOisH6zke3VuVFHothwKK
G3IZ4tAj3AUmjKeUD5UcPX98xW1Nh/nL8WecRTmbEXKbMB8I5+hptBlSmaezN+Zd
6jZcwEjjLpFVwNWXcX7yM04KTj/cBlSfnPTD4IIfAW4/Sb9h1zuM57U11dOReEME
+d3bhq5nfbWVw9QsoyGSSq3yc3VPJnDCUQtw+ommMHT9huu92fqy+dguaK7AOE+I
pUT2JrkqD/ECiC0A2qiaAE2udfP2zOMVqkPh1wmavEKu8qk/lQq7HQBJHQsH3dbQ
SCtgSFhR2Fx1S2ba8LgTgb4e62r4A5USubuVb+aaFWEBoPcwrOolcc9iVox8Rjp0
H8F4mChSDKPCZG+d/aBy3lL/jx/mjnI0PaLzOdZwBlAXIZHJNo0dNpkaMhz7dArc
124f8FlxogqGGSUuJP+cCXDYX2uobZ++I2SB5oswPMeqLJtm7Q3vDk/sfaHDhjbL
lztFkkHiOysQC2wh1fLnTKGdS4kVAD7V9FNTWOJ/GwKHX7pT8l3Zsk3DxFjTZ+pS
t8Uh9U3H60riZ+unXedrHF8Oy5OoDmzNEZHbbukgQzOZly1TdQg2THnC/eDmpUB5
XLOTiBVMgTZVJMrlKOrkmdirfTGj/a50zoc582CM5EF2qs2KQhITFHZQ0ESKmI7M
DYn+U4X63+Pdv4QFU/JQEX0XXRWgZn9HdWZESd/MvqlwWbAVgm6X+MkdIiiZlBVL
N9wKKE3l30yi4IAdg9k/qg+/JBBJ8qtdrjZJc0pMhtL1FwYHAkFZGuiOc6L1FsQc
NNC/Ju5xU5zZHzMjzS4TkIf4x7TwIk8b+r9KH9PWaFC301u0JAG5jy+cYUGKKVXP
xVoripvt5TtdWgVDvq6B2f0mHsWcHeZ6O0Kpfg3D6iLCA6Qnlu+ZZfQrdHRLQPP3
2IqT9hKIICs0DxqXDnLoGvEaNx8SMRAfHq/0m7+zdzRJu4HCZBATBhhOdnYOvdMU
jAGCcqpVIpYxe3wXZjlES6wrc5+nuf2kLYUX9OPpyuZiZ4bwfKFZwlmbJQHRfSw/
BIg22aOBCMPym03P5It11F6vMfgTTCqezZP/fJZp8l+aNZfKq/1aTYgMWRILXrnJ
w9z9jOLMj1Vx/UAixjG6hTksH8laM0XtXH/YUBwShGuPX44gGZjQ0ygtxLKmI7eX
7Tk31YuB6UdYmEhRcMu2A6pUP+UaHR5+tFyOtV2ZggOQtrWJ53hnF4q8SU/FDx+b
voC4dF6tyBMrht/TsH90t79FUXJx66BbdEltPFh3gAhVUV4X128idFLMSGdMi/ys
fcDc0eEqlqyVR1JirvSOQot1L4SMoowb0vr/4YXJNLP84ccW5V9SiSmJu7vn4UuQ
RFEPBANjX6fDZ4e/wo/P9nhphFbgG41L6SKGQCEvtFwarXBYZL7Zbr4QhtwU7L+3
KFow9s9M8ujKplWgYSzQUjsDsAXFY9O8Vv10YsMx+txcjrp0GEGuOFB03cKOidid
kFysZFks4wbr5N1+nTZI73uvamVwuuhRUcRbQux0XEZA5/6RH9W2kq7/YjcqeFP9
bmBl18tP7zQxqWQpob4PLTcYg2Zfd5cfl6RSaaHTS0Bh6FkN9hcSOFcl6WgXyLc3
sYWRUBf8XY4acdi0/JW7EjmwmCFWnSnPub8zb0QTPpE2jWgm1EipkVBVYiJN7Xaw
X2Tt7GJgLC7bmQ8RrGBh/3wdsYNDju7Zcwc+JluJaxB6IZOmXrErMo7vleDL3X29
lpRWfIDF2q0vn3uCiTmiiOU+J8n3POWBj+dlX1brYhUY8IEuoysrs/f+gyFpZzBx
wG2ySYD0x+wom0ivYgYQyZrUuzOwFSU1XWy+UDUBn9d228Ba/GQGDDXSsVbVKUvr
EBcefaRd0iNP/ugEHQEodZePSNa70ubTdt8WT/jzKb6K6MPMCedvT5S5RT5nYhNK
PpIkdI7hRSGEtQ85BuwTy/f0Y3wJQb4J9F2omN6GGgtOurDHAqld4kn+mFONpMD2
Asq6f8gZ1B7pkUq6YxjnXUmNoZmmDKaZJp+0lSoe9cMXUEl3j4UyM6XsDHii0aJR
TKzOK+b7WT1koo7AcZ2XexdZEaVLsFtN79OOBuwaC7yxqQnXNZHKHKr+zWtE+Ib1
UecGjTnigeS3yjaE7Ysn1AH1Htmp0DOVeAdTjhuHQNlpZ72SlFMTm1sLPogZu+W1
aMukMnDWYycBfwgY+GTZRX2n2WmzPhX0dqC9S8jFPyJEHsDtFyvOW+T1sXsgxgLc
2+fQ+7SXXgnl2rSNYOga0nv1U6IC8d1wiT6yXIu49yF1edDbTIq+EkrUSPN72Fz/
zO9Br4lwRovp/U0o14TUl0HLMQuZ5zUARwQ+HQ15f0kyCX3zuKS6ACuHZxKCRtXv
7HnQ/kYNGIVxBifxJvlgigOPgYhEyKy3DMBF6Xe9Ndp8CLGC4l1ZA++S1ScyLiya
BxyLqPXYlu1hZkSv59zZGZNW1pmxn6JNJYIXKjWUsNiVZlL3B7/CLk8zkJWT4nWE
Yp9N8Z+Yq5cIe59FUsLbeOImkxp/nzN3/udW11Vsj+XQqRGdSpDayrc/Nt3vJ5fu
ZhpzDCe3Xnrv01FlE0zU1hzSDFBQX5uu6LNd/8c6mvky0Lvc0vgijS+ca73jI6Eh
Bnne50e3C/UFgytjp88UQbyQGLJF5SOGEQ8oT378IhBQTc83LS+7Zgs/nCUsPut1
VEVpdB/w+smPZM1rjpdbUT5XIPV+YVdKXc6JUMx5lh1BKGnhFDF0JdLLxQKVGzqu
ugWSSV+tpbozDYb5RGPvRi2AZ/nOql29KkhRvkhocFYDgs0cHnDbBU5xrfLdNsa9
6nZpGDS6jgsiXHfKFsSAIWgqHPmnaOZXCKSnbgY87BbfnL1Rn+wxgCG5I8F5rKYx
0eYzvKZEkWc7ZvOmnhCE55qVRYFn9tG7xTSJ1Bs2ZbU+85KL0k+89oyHQstP1kXB
Rk3anL9Cyrokl1eQ6GfHuA0pztWu8pWA2Q/p60419PMx9UraVVlpdxfG4cvfxiot
K93eW0JrfJQS3cq1tbFZLfkupF6HSueXux5BY00UtIQsBNmntOhBRzCqad+VjCyL
9z0pdqwyOUDdslnHsdHrrapWjZ4toM2G0pf3qV24buYAWT78BjwLR1dWbxFy8xpT
aNH909fRpNp9OJJKs8QYgXqPK3Bz/kJ9hoMW4NzJ14r03R6wcqgUFFeFROS7AdjV
iKRpBkrdNSdFDkBFIcR/xUOYiyPbRbqS3Xlh+AD78K5s0tSCUnku6JKx7VSJTvDz
x23a+jnVBFJM0y0+BmECuIuXwI7bRkIVcsjJLD32hW0YAp8jXhzsBbfh6KciNNXJ
9s7qnTc4uBX/GiOJ1dJ0qO+nU5ATGT8t0uNYUSvqKAJ6eBNfSalvP4WDmgXAJR7P
iD90Ne9KKmkgozY3o7XSQcU9iBCE7TG38FoeyEPi02pnlquHPPEkjcY2YyzGvnT7
Qj2hSF8PX2V8tXkKn79mkBeJYGqGyGyJeiWsleZhTo1HTZZAtd5Z9jqeNLHaVnwt
zV/QSAs5pdR0PCGoJQOy9zie7EbVOIur/dTSJgaqQSB59WVlBpk10HQIBEgxCIfL
f+kraMWF5UCW/uQvS+Wd4+J/IaduyL3PHmq9tJ4uXs52zimZIHGAsQBmMdBoSv5U
Aq0FY/usns68j2+eDMGBOdIGOFkHv0+/AUpjLkmj4qIgpQ1YVMtNK+xrDkFp0P5D
5tcD4Cqc5X826YbZNZw7mbQNJbFqjqUPdrrcYoSj3q1F9Brwh+qiwkLcNUIkD1jD
0Haz3NMhakGrnfjnj136lsYBH9OowE9JagcptMif0n4vdh+HiKzYr1S46/x8ktFo
Nko7T1310QWkp2jE3pCjX1qRqAFINz7tHYPvRckFpKUERLca+kVJejt67Pt1kAMa
YPL1Y9ODcyhyL46fUCqQkMeqywPTAxbR5KkEmT7IWKo7GTlb8pG4uL/umqNKpose
YFnKnuzbPv9rODt+u90PdryTUBd60Sn4oNawxajg/9ZPlFjWTUbHQkvkiPxCxoC8
MIuWTn11P9Z876hw/jHr/z9/4AFZrE7jMIBBhF8ZUoqDzXDC3vCrsPDwnaa5Pxky
pi4aA4sHK0enWoZPFrSVOWw2z+t5tiqAjFz/c1LPDfsBvKG/5Q0UaWcKhnssSXWi
PbmF1wQ1QJSk+SQLczU2mk+gCtleCYXlkSsMVjKZKzQSLjDVSEZWjciEmdDusNkk
oPtzYMkzc2qVI2mOPERrLobMF8svNrseHBeWNzRWyrIPPpbOmWRN2eEvaxBLD3Xg
kAL/W/VWxeHP5vr9IhvFewCAzJtpk7eVq3QTquH+hQy9aokDA/rFscNqgOy1D400
vzYzLo4g/5JhLrTXYEuW7dUHkNqrHgKSfCrLAqyOkaSVxfQw4G1krZLwhC8lOw8a
e3SDlbWPA8FsR4jhlINywqLcd5IHlIMDyCsZQtfJ/Zlwnr6CRtss7DZwmaIXQcYH
aqnojzOcImeM3FeySLn5H7PcyEVsZMYydROStla3CamxzWHys5k+rluwn0sKitep
wy51lI5Is8Ofxv5L07rnisEkH3TQDgojMHnpzNTgj9THVn35I8vlyr8Eo8F12DWk
lTNJljIAtE7kyguIotb8G6ZjsKOwX4z38vFPGA8IWM10geinlYzOYMtqyOZLU0Ec
m2SbCB4TjtOgGOJObCovPMz8+MRKhnIEoMKqbXiMrX9aUWeZKMxayumYxGDvVPP0
vCjrpb4Mo0iQeaIN7RzawxPKFUVr6ehbYmQGCKigpzUG9aVQ4nwCT5wRaWJhWtd8
b8tpfrvXXw/actDaSf/nXkFhnfMT9lWxEVXuI/Rc/4NfOGDYmpK7apV7QfwHJEED
6y4M0N9Xa9C0/51NSuXG8lXwVkMFmlcqQcds84acMMkVhRL0Q3qKigft5Vh8bOR0
86ppFQZizBTS+SJ+/WzOpTq65H/LlIFtGglc/D4MlOqjRKnPEkDae3LOi1PmDO4z
HhNqPc/xv1qFBY30kCTc99kiQRNqlJDC0nlhmVTXbKdjEWgsPP9/eEkvZWVedKQs
DWfwxuy7GEDy7WlEjDYhNTDSQ3tzs76oUDQLXPgbjdM6LR8NPC9H9I6uE24BvhoN
q7hO6zbM6196OcooxZMI5agnmNYnzwxoSbkwCOLrSHcCnysA36Q8jAJ0r+ftb0EP
SMlFpyo6PNlKtrfsySwRA4DDjVNC/oSFRgPunu+0RzKbD+Zcnq5fY1irSmHB7AWR
MC/ORGkMusbcYLkq40sx1UhbiZOFhu8OIOkleD9FjIKD/BuTRXKQc4W7D12N8aBl
GCcrk0wY07cFAwXwmmCPVSxd3aB1xLOlAQ7DIhjuZ4sCdAHtpK1iC4ZrfvONuVMX
QN/wiLahj15OAGJPv82T2ChRQ8yPWRpanltQajM1PKRcBvY7xKTjrBSdJiABOyY1
YFhxccFxuTvCKqTbln3GEDJaBGBBq9o7p7k2Ayt0UBKwE5gkEfftiltFEccG53oq
GDbX1l+W5Tv5X9EGmRA/ozbJmFxFpEPEk8mueR0RPBQsn5hcLhgJljaoLq1Y4DZu
5zpyDtwL6aLUBRfYtsv48+hNVUWugnL5xireKwV8bBuwt8bjlytiSnVAlFNjflej
Zi1oCBRLE3ZeyGwJTUI/9QMPoMzFZxH2VELSnGW026fPqXxf+y8O9eABPhczhH0P
bN67PJEheQNd+ZTRfPuCCcGRwUawwOOptfLHCpyLSULXLtoPSp3P4VxJ1sAczPNv
ICrCNrJn9RVEBO62ZsCqQ/+khof46ah0THq+9sz2CJfQSTX5KwI2FFoVIVTkazho
czbmmxlMfgIIdlVRjw7aJ8gN/av/GxzEvkW6gYqpPdFgLZuchFoqFZBgC5K7JsEK
50+OnhzCBdyDi2GZNHGiAitVwml4fCzuejNHJtnh0rd5rTQ81kE9s6dVtJyip2ab
IUiq8cTwTBYI58/qdQd+ITTc6wbf5HblBKzDMnJq4XRKy+DIqc3lqWfshGFNlw0H
rp2Xt7qVZ3SX1L2Pzr9mrkVd4HV068LL7Cc+4ljFYmEipNU4pjilesL2dEq2fN0x
V1+e1WHDOqV7W5E/YetyJ5IaC1f+Sfo97ZcKmaTvA7SnnpXPi00gvBDzvEKvP42F
9WJUFLnmbpNRX7yPXOpvjrGc5EFmDosUcpSW7bxE2NXQLqCHnmnANquFlXjzg/xY
23MV3DjWqVpmrE1PFSnoXBkreS1NI0TUnArjLDEhFx+YIk7y/ALD44iDBIF2xOnM
1QUtmuQfxMYMOFDT+BRVQAlZ8Gl+Y8aeJBNWtM6ap01vRPjLBrcnJG3ARPgvsWhS
zXQKeVcpJImkjSQBT3jLLXSDcoQ1dvuaJiM2rUdr8as9Eo8kb0IV56oyfImZ2J9t
N/mJTz/8lBFP26ImLoKlC5Ls1xfGEisju5bMEEIrS7jjsrRTDV6YEI7ZxUFUQPCG
+5XmHKx0ACFeR/kGPc5w9RJVRQxKxRK3dEIysg4aGBkhSdiRfHVlWpM6i0d0+D0S
vhpA+1H4W7CJyHzV3qJ+9zgxVYdMMzRgV1tXt2N+wveVeJGAp3Jmz0k2dgZRNJb7
Tg3DrAKy3H+z1ikQAsMEX2kzfyO590vCd7i0yechUtTK8vFCM3rf+0m/tIB3E47X
6iqa+guQIRL4ZwrC3AHvd4lpWPNQFQLrfL7CCQ1K+lWhcC3UbvTCeDCb4w9aE3GU
qWtk1+qv6EsA2F/KWJmCaKYw60BwTQLQiFogXJ0lVhrdARb6bCXl8UE0mqmAzesA
+SZURct9pzb9SayyYttwaXBpV600wjcSB7UAo6Tah2prb0FBk11vjxzMru5JKq1v
GTSghzisyupCXk5OkbbmPHVkI9E6zZ33ZDdGZgAXOXO2IkpxuQAQKH7aPapr7/NE
QmWhuODSFCxtTXoyPyXiY+uuhyhteuXIeLhxpC5DJTaDIo6OQG5xVdK/AlkOvfoI
2/Tgxru2fPgD8RejjPqqig8S2DsCUgKyWS8Jxdu/sbT8FEwOR3ejphAW3UfFG3Kv
Feq4YKbDglGJ0+dBQkivPm19AZ581ZjIwI+VPDqqHjbA0nxzHDUa+llV4IUAAYT5
w5iV7KdQVVQ2KkP8crGhuP9ZEhUuPBcf8quiEy3YMYlgwRNTIOacjPzkYGJlDwt1
TOrL1GVTTZ9z4XxHZTr3D67USTiqLrFJCf2z5sUSpIfEDBkSpfgyVq2l6zOc459v
sVDold0W6C209e5O/or4mOFrbG/+PZrFmkmU6VWeIfC6JyFPt7/zHcI/oJDBOfNl
9WeDXTcUd60ASm1R323VlYR4nOvbi8samDmtOdAIgkfiv97Ap610q6g2RqFLwBlu
FWNb4tRGuRR+EL/94wF6jxH2vZU63jE89NppyDpHpAaYRHAbM6cdvfQjeGgdzBxm
DZC80TQMXLE5yp/m5rRC+JYdzZ+Bq3uKuMvud0Zm5hgmeSMOwItibTwGRslYXQSQ
EqJ/DWBmI9MrRge98vIpjtcXudbtqT/zyq7uFx/xk9GMt77wyEHKnBAExkZGF2A/
+IpFpIZ+e1A3COp1ih0zjr3k7lEiya0lfxR6qK51JOAJYXFzRnL8VMeY/k0WJ2Sc
P4qTgTrshgaXvQwCQbBWhNIk5U+j1g/DpBCTvXVk1SHBWSH1buVPdruE1n0sntps
oKY5xiHIcOD36+8pj99DZlu1GUrwa+bj/2InTkuVKchqEHvVRMdQsq+zifdBHtNy
d9mvnmI0yMpfJXX7QpF1NhJqyx2IpZCSCpL0VmyolWevvlnsP9BP08C43GJ4z7dE
y3hmdM/iguHyAH8a5GTA22V4ThCJ24W7qzlquEVwl0m5Y3zyqTrcZ8ZO+jfLzNfF
VAjDosW9F8kiNePj0Y3sqXB/YHCw8AWlA898xGDlnHZ2WopePG433mSiFsulRzgt
ES8MNv4L7/O44pWG4HYJdcIhZk0C60WMgk5gFa8cyNLvE3jttEfK0lca/x/X3n7S
pHXTfx2z2ekGstQInDLsH+N6GC5v7CvpHHFzXnZsp2uKLr1mEd5Jg+Ebv149evVA
TJ9meG+kMMdbHmdOhOIQw34rFdTS78sKeT+8ACnbjMLhxLcq26yFbLlXxpdA16IY
sRecIQ4fSpkBnL48OxeWUoBNYtznPqeCDEriO8gc/1oFPZBA8R8G8MphzgQpWOol
FHMmi8IjahAdNuk7hUS44U7qcwcWcjgpSOR67EXIdZCB7LPqJstRWyGpl0PuevIT
ipWSYVmoB9EOD4YYrjVPqeGG5XTiC5CYBxTAVcBpGq10vAHrp5DQFR/SfiYKBPZz
qbDgxfvyFuf9/eUh6IOLioqeWcu4lD4F/dJ8jlwjENVNQGHhdNyjtFFSnhZSJxbz
JdJSKX5NlJnfaA27gLZyTu9Gw3Nl6t2U1Gip58OhmQ6DB7RQtnt30VlLIq7i0vUU
1iBykH7/Q38j/8nruQY49FxR1RlCq0Ll2I+RG/dMSjOqVDQRNyMH7Zl3+xGRIJQo
prXakMjjf+rbNVJu08E4kenoAXKMc/yVycsL8ULYls2XqzgUmUND37ixYg8Mc0vk
Me0ubmU62P0IOnPWhLRli0fzRk6ve1pp0A1HnanqHSEvIxubyGmQsi7I6AOp4O4Z
MTRhXgUIdyJuUhYSsQxV26owp252vJ4kG8SXzyi57tRpI2fgaFm4vafuh0QEm/pu
oymF2fwfGlf7+Zyre2WDR3V1260AEOqZFDwDKjln68hbG3UexR44QReEzsDGyAzk
2DTTerR90XGZpya30cYOQMs6eyYAfRqyI9Lrqt8VS4JsmOPaVwKc5BdFT9wi59vO
Rrantwp+CzxAsoe0TpnVP5QTKhdgccVz/KFt5DnSKLSYQyTu+QuJNx01rMyXO4Xv
WSgEU1ke4OXshGqXSKYmJDV3BA0pEavjI01upigzMNAlggnk2dgk3rb6vtfq0e+s
1+4efQi4UBd+YUVDNuj4fRYmo24i9BtVz6rkS+bxQtpMPvB0LoiTaCZgzwJoMoim
lxKyy6eyZk2As2KSWMY0JXQmKW3HW6cIH20pSnoPnGf46kIMOv12vDvj3IkVZ4/k
/jXjV6dTWBtH/iB8IZOMXafDBtyOq6jsLFoCTP7Pfr8RDNV0Q2ul9THI44/+8OTG
xEyHfShrhrHvi2tr0twMYveeKV4GdMNrZ13zVALoYPL5J7hNHzJqf3cCAOhdP4Ki
tDKQpr3Mm/GssXzTLklVHRe/RoBeGcSs49t2sifo9m/CUWkgoT9XwGf2xaku7Q5Q
epmqez1wS5xUFWap/Jc2qTyDxzD3syqFv7rxpJui7lA1qzc5fP817gExWmyVBXjh
J/yYMY/aa0zPgVSZv9bBG58A9pvAcwi1vs2ux0Wc+Bj+I02kr9A4NQhlaSeszcnb
Q4Mgm4WnbUYJ2BMdmjAqLgYR8PJavED+KjQH12+gHYT0Ox4u7aTCCqxNBFX3YZrK
JD7OALkqc9jMOfNISfV6d2dvPc756d3mhuieaTDadK3jH3mWRhYPPMeEYcLsru4g
n8qK9Fhk5Fj4dJWFGHodhTt2y+TtsatjeePYf20tqIlJZcsOaVeiVBYQo6p4dQw7
9M2v7FF4FBCQsur8P3AEMUCuZxX7a/t+RGJKoaZDX9HQq4UnzxzyE9wjjB2lMMNv
yTv2lFXAlR1qHQkvEEndMhwqB+IobpgWyat3XWHYkbrZeMY6S163yTwYNPit7iQ3
oVSvUjG/Aw7kDEAXAwqBfCXv6t9bi5noh0ZncZXpIFQGQUp7yZtdV7PjHiMlwsNY
tTZbdhNYwzLEJTU79/xIGJjyO60vwCPkh9FlC9mUebPvrjfyUAIbQ4T/OhO9lCV6
lu8pN5QTeGKTdY1oBMsAkJltKkpV2DASlLTLqdtYetFNkkqw+sdipbAjlrRn7QHm
RhIdfF1f21OzcA84EvJ7xUqxROLJTQ8A0V+7D35jovq1US3JCG707ObEsUpiHQcz
JJ5FaBzVAt8kfe9wXQvMH93nTMH79iuTXo6DAquYKUdDnH2K2LNbdrnz6h5DbNGu
OCWjksaiCHLnGJlD6IjyrKoVdHbUAtIVeZl2xB02L8GllDEVyWdExMmcBCj1IRYr
rLtjk6Z13r8NFOfZtk75buaF9DfTFMiVuKyMOYGxcrJRcasbMejiuUbkCZw4qlPl
UKTWImh6Iknh1+aLaPgdmITxiUv+ibMs+V0rE8OyMcja5oo9yEGcRdUICD5yf2uJ
neCQcXZ2xiGedBkIgl75RJsrl4mHuPyCqmVKyRt6bggGHu2dGAcXp8etJxvZJUfJ
zsLOH6+jLVySbhdhkpSeT5jSpyXv4pV2CheRPtv9XPD9t8nZuYdD3Q/U1OMSu8SG
IxcHWtRu+Revz7RVrUGqp4+Gmoj5dGmRZwnlGFaeiTxHscvKa7u5BKMhb0HxcZ5S
zB1Qi0rf5Zd5I24EKr7PNagz1iAML+sBPYghrqwAl3VZjESeMrZZM9dKNjAGEQBS
wU/eGNA8/M+PzGdaEBD6RTrbLS0wWh23VShHcdrr7n/7OiuSjBdYroxo4LrL8Phv
QWDGnQvO1sN1zBT+9Sep4nt7yhicaZadAgoR1J03LsXNjPcN/DFR1u61ZzUMXXPD
arURX8v4vs4/6IQHfI8mkuJtGeoEqHXA12SDMlDHjqR5Go10PCygevwv2LPO8eZB
buGNQekKc6ymfeTgQ0N3RHnNpYgeBqT/EXlVDesmpilj0Y1EGTvwPmvjZzPUd2R+
i6sKcVh/HguOeoYYcvHAycbgUB1l8QFDHup0Rvox9wTNZd2eFMuY7eNS2R0JkqD8
d3r8ZflU1TZZhLPxXVGvdvoicTzIGVuCYxJEGvSk8beS7mzXIXiYZfBtZjtCZiqK
QuirzL8/NGSRfkMqGFsUpfPi9qGeLl2va9LxPtHrCaoDHGLKuN37AbH/LJGDx5Ge
UNy5XZhbXAm5nxsvPHZnJwAGzZn3csNcHL1NKv+9d1XjT+KqPNF7H3yJQTgHSaCx
K+y4KKRfeqWWgNwAXhwA4K6ugP93WUMPZ0P4VCfdequKNcjsNMoOQTMZx+e/7HPL
H1CjWydZZPV6iOdHT3VTCfh9vDDIbGrMk6bcvey6OWWuNg23StAHOBoIE0+AY2U1
o1NdehkakjhNzRUEuiVBjPv8QVB7CuRWr+aqIDiR0UjTJG3fy98J5Rd30zF/ciXa
ufLluZH1LGVHGVBhfxecd4fqUiIeO7UOpmY2tUapVkWWpUU75vYjK/SL5jCe2z17
qfYpbvkFKyalRZ67+FMsW4cVfeQ9MZZejlzIfpZawMaNS7iyAqEnM4la2cK+wy41
RRkBFWc/ZFAlo/GJby1uJE4F+7s7j/74aZaI8QJOIaEXetxYepv49/lSRxgLndS7
539Yj4Wht1k6/uOEG4JtH6K/4+A8JYY/9Se1178qx/idOnWOu/B31kuSr0x8jpHM
WQzTJZfOh+YibV8Dhp81r/2KmrH+fXRrMCmxy743gJwr7sKexZ2jzZw2jZpgB7VA
FDhkPUSlqd1Dr9kOUDaRZlJlCB5kNetL5wEcaVqwZaKyamYKas+rj2AlM04LFxVX
+MIzxJ36u8fodH7mFayIUt3ACjjPIk1ydqN6yY3B1wrFxn/PzxFWjb4NdNVpIqzq
L8OB6irkstJs/8YRjYUCT3Oy4HkmFPr5wOTiaKRWl5TROMtK+ALswtyKiH20Dc+o
7fck4jgsY277nt2RYQsntqQn2iCzT8wKIqnH9abfagQ1ztrd3bVYwmqLYY+YHxpe
HbexpWDljX+R+dQJjL7MyVjBqPUr5rNfHzqqWk1qccG+Tbn6ZeoFXWyJzQkK9oJa
nGEwNkfjYJ01uhWHh2QDjSwO/lmvwHI6cpYwhsHZ88J9on2h2skX3fDzPnX6svxx
PNCy9nH1+OkmqsTQzz+wTRfj8narooBC5wBYiaYKQy+L30eLB0pxmR/5GaqsdA4u
Gf6h3zYygm6V2ZwiKOiCdedV2ScUSDNBmPixefTKKgRA2MJaQW6zMwYy9xlgvSl8
5xEF/gMF1GPKa3U1WtAz+9ROZRbLwlVzP/4kVCoElt4MnMejEO/fcsMPuJK/ABQ0
8bMg8PpyEtVTqMCxkdpEWdIeZ3GxsWJBnBttFt4TNIf9Wr4y92OXj0gmhZUis9Qc
JfJZ79T2P5tds799Xkx/7BI7uN1isBwZgAZhlVISFSFH4mOWiXcsyvGI6+mIrqS8
lK45cZSC6VcWEsZcwRK3PJTk0Bsk3tIDloEF/TSkHC9oOBh+7xyx3VOhk6Wh3aq/
8olYZHa4vd2FxfFmBd1o1XOhamfhikDu0ZL6Nyl5I1qhWXEbVBvrtETlakQ61U5T
TenK/VHmM2p10zQuJq3rBUp1i1w0PxnqXZlZnDiP11Pwr6VnSUtP3GnrUZxRnnsi
MZIX+ST7vtMz8DvEFWYcLZILueKhBuvmSCPG+Dq1BRySjfvm+PxpkyBK3zMfWd0U
TaJIyj328K9J9trYP62tWAiigJyibdI6jR5SHOkJl4kaqG/fkXqEzYR0/qgnWjG8
h5+NDQVyEzuoVqWeiLgTs3eUwsUnv6Kxn4WcOR21P+lZaQtOBfhbJs+VK5n8eYIB
UY2H7xrcaqSiNjLWVYXV96FngLhdhINm4kXt5EH9mkxWTbxoHrfmspExEuINhzsY
Kt2QL9ICaTHJrm/y+wNngWKOEH1x8CbD9MndhAclPcUwaUbFSo11m5mhtrg+ZchD
IOyLjRtfYFZs+ystcZexvcQbeTo+J3xRpcEXYpYB+eq+JZBfu+zuzvwQi7SftYJE
/SSfVS5unsX2b9jeRBgvXRK/9evoWAlG1QBU++JiGtjFcK+6eiVYxGipMzZRQamW
bTdchkkPPb7kClHnae0aRBw0KbGUl54vk3EtunzKix7P61/7O7Z/Zw99F94tvc3X
2sLJKIEEjPuPYoJcqNmfVk+on7+ctlo0Oh6WllNKF0qf5jSPGK6OKcTDL4nTwx0E
+8GVjC57iiLn6aaXQgwqkCfMGxz+ORjogLyBZb3BwCEP8X0H5rWIrT29F+1sUTW8
8kUHla+w4ytUJC9e05iW3DuDXBmyDu/WQRft7eJZhm0ecnu/FgrlIze04RA3qLDs
GYVLkSC10f0mV5K1dcYmKjXAxbLuleS2QwUybagzbfUliXAYOZ8LmxH7uFKHfWA0
ZTVov5ulCOWNd3zI3Iv8J8BazzzI/UOOKXIPDnRa/KPL+yk47CzgfHrlcIIm1riJ
TpnoXMi8gEgNmymEeDBOfnNx7i807bZvu3Z+iXK2xcMPGkeDIPxD9oZzJzWYT/tm
EGeTOHu+4HT5DLTtWYYoRBH/bdI34TLTUo7UOn2IidJl+o8slMqS2BmhBjsO2ZcJ
Kn1uhbsEIZa+zCZs+rLONA7Y5wW+G+nzUn6mliVN2lZ2dpp2MYIQZTArYwS1Ey4j
hq/59RL75T0fBOU7JVwP0DxBIOR5AZDrLI/8nctQQYLekMrNaznJ8V5XRax2ebTx
pvbOZ8kJymmCFwC4Zf2JuxzQLiB1zFnbNys4hRXk9zsF9u0ZP46AWTxK3XMIC1Rz
27Qz0fu/PJo5gJlJV5VcC1ef4qFrDYtY8+W1G2WbU5NQyA4UK0iSa+6QZBLvRmBu
pUAVpy8m7YJB8tb1ylFgX7fVUBcoYPnzAI4jm0Ny856CS/ddYg83MKmJPi557Y3c
FT2C4M3yEhuBJ0S0Qd05IRTfjpBNg+7EOqm8A4k9K5UE3nVjAjtHBG3zuwwG+FRK
+hM1jZu5WrtCELZTyT4gO3ylbzXe+AHp87slodKOK4sgf9p4QVu60COD293Kphtk
cjhRDMnMVMgI1qWvaF3ra132iXUA/NXNkudymXLVWrsdEEZluYTxsdatcj9szQqH
443g27/Y1D/haOKee2Jegzx+89+KyiGGD7eeusmsx5Wj0BQ0/yKSFSLZVE5IykIG
`pragma protect end_protected
