// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:10 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hlcf52o5K46t8BD4EfQkNiDzc7WF944eOqNbM++ANwSaP8O9qg7nXQifJKNPP0Kr
y+4vJx1yRYiMo6Vz7nCpG3Wd5lbCAClpqxgVlAdzVxdjwj236GzcfzCvQ0OTdZgz
H1P3hrwJzp8g0PGhCrWtEUuC75yV+HkKL6TQa7T/Pe8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 98368)
yChkUDc3TyY1VBr6l6TBy5SRa4EJUjopig7qxmag+SMYvqaR9iCNgRXdJK0HGowc
f5YU9Cs82fda5kFU/NO/6OqEqfQ+xCcX50LvpgIRvmaAOxAgjNEYV50Vt+z8tNiH
znXDo60VG77b2ENg/YtWz2mwgJsfUlOUkj9oL3VUu4ElgW7VokyH11DtBFhMuHiD
o2BsCuTGU8vZ9/8WjXRdclXTTLUCFwuudV1W927010OqfJvkoUEMgNFjHlAjyb7h
joRNJkbmBA5ZVUioWOLCpopdatTJLyoTJk4F88CyhRsPnuLt5N+Hwz48L03/qZrU
o5NfvzhZRVJujJhQL6IOdrIfWlc8D72pNsMQLSxFW1LcWcnCzxtXseRk4vaweswf
+pHk2nwvrygQME5MfE0uocpkIQrK5t2LsZn5seZUHhcn6QmnMd8Ko7Xqt5VoXY4g
XL3WQWyveUt6SX5g8VG2KwRtlgIeO6oxLMhtnJ1Y1YaR+WxLe8mYiYdu3LalXYDq
J84Q7voXXXe02ZBC4oe3oc8DvT5bEoatFMBNYyFlsbPlQd00PsbvByUNtLmUbjNI
rs3o7Vr58tQ/IARTkEzOyD8ACUa24p80Za66iFUsb8WgC/OkkhgbmwJUq55MdSyg
F15NyA0yXlT1ElgGM17n7mOTiSAnNadqoA0/mcwnW5A/YYCVXV/VMKnnCuUIQ6EP
ZHN0EXPSZNUuBoCF64y2UwM2PKqwc8IV0Aop+63fZjcVEx/H4LKpPdiPoLgLXDyf
3k8UJOkcDzRDixq3FgLWXQ7X5sgGaICsQiuec8f1ueI1GFDlCKgj86KLz4NnC0Mf
NvoOpLY66rZ/0zHCK1Qrk/zQSvcl120fqL+4Tqr0HFq7fOfZtxuVVrrjzFd9Jev1
qEJvDcO1K2vficKEWFQRxcGP5VvbaRXwBtnuhX5dckMNYFNE3E3RreZGo/VP0CsI
qemBFgdPeI+d7QcEUuGdcrdMBnv4Q799HMV8kgyNy8fh+ohSi7GgY3IqgGD5YFwf
4+oo+9a2m6vRvJO1fPHbfEiQXpeI/ZPjNhg/KPJF5kGvtAWaPO7Bw5FLie4ce/wS
9f9hCmtcAsGfV9HtKX10WeCk8AGU8Tmom/ClXIWA0rOSa3xnJ++ly5+toWVUxQjp
VtsuBIDArnXlXi4mw73cv1Sj5cqlIUJkmEMBg5AWGyj4k5MWqzclDX02eI4ItJm/
szI0RtKMQK6xJtl9C1ejRl4RTNcVjc6qJjln0PWBdj4QYqtm/sEE7J7cu2rOHT9k
Uea1spLchS0EhbsdFFVEwhlKVoRFfx6rsNFK1hgN6A6Auw0mS0o7b9wkeOjOVBUN
MMMemjYl23hjpWaXvCSKmC2KI8S6QCAp0k4BExjfnZ9wDe0jtGzF0hGawVw8s0dk
Lpv52q0VtLjTRDiO+T7DKBNFb/llt4/Oro6bNMH7ZiM8szyEixhF2QJ80Xj06ot8
MZ3RPzXOPXzyrK2kot3FUChz4Dksq2cyShgWSNzEqvbf154m9L9EQ4+tk7AO0V37
zP6ABr5OApPBA0f97dNeiVPWhiS3Ukl7+qZHBCMWXNh1s4B1PnSKrRSjlB/ywthu
9fybHzqMxPY3vF/NW4ZjZrGUII8xvb5jOE/8bsoEnPET6/w2W0NsUgvGO9pwtr5z
kDGOoHpUI5jyBi9+dz1A64oVwEA+irzjVyZ9Y4tOid1t2bQFw86Xrt4/e8zcQWoY
hpZp1UKwjUvKD6zXJnZtb0gRFUBtUbmv5XwD0cMZh+46nU0o4U5OveadAuuCZUph
p+fp+kHzUsbjdyzi5qW4BYm0TLr5f6wwFlZwVZdFatPCezbvYdYO4+uwXaNmRs2C
qp3PYqjCsBtKMWR0S9IN7D8kcwDFiRJiNhqAECckPq+xtjwKZVKX6whu++j3pE2P
CtqH8i1EizICZaqUiAS6oZb9J69rYZHxtcyCVB/KJ1+X070Bfq9OQVe9U/xfzyAO
iwhBz6+WL6pVckcoIlLFjlvk4VtKFX0m9Pin846/G0ZxC4mvBc+blpyadpFCmDh9
OqFsPnGTHhQWJwW8aC+jDH6uY7ckxjRjPV7Eh2fGcOrVY3gg5tZvdErNi5Yp9KM7
CKtyuvkowHxV/rSf5WV8GERfCpwTrJgX3po36jeK/C8+hTrstUE6iIR6VqG0DXZZ
oN0Mwo+Skke7RHxQKiZ2LhTOchjYYA+nMnWkO2M5jB6n2m68bZSaPz0LNWy6RKuM
s7rgJhEstUKmDx/Z+BfgttiSwr2Uwj3CT8EHm6cERXRZDnw6RJoZYMpbdoE5tbHr
QQWcA3T/74yboQQNp2TadynnbZHxQJDIo0tLchzSmFm/afHaVfr3YbiGZ9QgPSMS
1LO3RP3fyVYn1Y/pJTtI4qsr7ku6dAoUdOZ5y9h+GbLmEvIcMIdCERtdW519JraW
6nSCWB+CkQzookSPFO8CPQzcHchtU57W1ocgOOO77shIlBTtHjspDr5GeyZzaTdV
zfAaoc3zmurJZYQxZOIzwUI7+KMn902aIRb9yGZYHmQw8ujkOSd7wGfnT3AMXiAc
dDV1uDNwEmpxVdvh0wVX81/nFqldaJFLMjWLZZTPbxC1MPJg3Lr0Zc6NN8zbXHoj
cl9qyoNuVkR+Ya54Kyo9HNu/ZDnrTW93MDtFmN2WVxr2as3ns2pZHxYIFGJb/XHP
D3GjKRT5ja3d6cbvcQviM1rWiR2pCngfhJ6E1ZwomIAkHJbZGysM2v/dGKqD9ypd
JDEcX2G64GiCuM/7Jrxo0NrN+airU8kPUr+OY7I4KKimG1L8tVVybUav7PAnD8sP
xi16vTvg8sV5EJpt3To0nNEhwVtqgYPZeVYoLffRzACLot9oqE/aMlTUNxCUkB9s
tZpaT6TR+rm5jZswueAO7OZUFhHZVjUSnnA3y86t+4M1draWACqmNGQP2ZWwbJsR
esFmm3gYZhMeyrYbwRD2VdFrBTHcB4dQotfcKtzu5Hwb7J6cf2s52Goq52zY8RdH
Uy/mFF6EYb6+pLceCtUTy0HLfF7U5Ha/LVcguMLiNpwTZye522XaxS/9bTP0CjMR
Ykf9MLjbeDP2nI2enpMpWCp1s94KZZ7UX+2Q+usLxOHyBrk1JjblE39iqXKKuRBH
qQM7ReoFOHshK0clJYN2Zm5qsz4NOsRfpGSVdi/dxAMMKW9NAy5fGyJcEHQxQfLm
0sa7sJljB69Ck6vXFIBbRsoL96jDYszBs9OD1GVgBxPKoIrcBSEcHqjLcsrh4m57
IbA/M1NxP5ZOsfnLRZufsZ8o6cU/6ImaILI/BwNf9i8hgsVDwOZoVqBC9IV2eKk5
zceS9Qei+DPZ8pnxytyzBXDqpBM/2lTLwLrRFcdgSluGa5v5R62aMeh8AgL2GDxD
KV48hcifX0DXir5pV5GYbVi+/8a+Pa24/ytheqmb2gJllG3K+cDCRMKum3Mw8pT2
A1sXz7ZeG1g4XTw5EyQh9Il6uFevdP2q5a/zlNEbqzm1mmVcVFFmm/nmZYJR5s8D
XX3poYVJUWZc03c2CSxCq5ItbbdKmbUjQ5juLgIPCpE8HHDSwZWZH3ak20tMxodV
4IMqLz+j6ovh67XOv1Y+C7hL506L11oB6MeAYkDzGHjumypFs5nmtUj14Lh7BbNq
wTPAnZzQg5W1bhj6VXnMAUlYNspAdkpbVHOv5D0MSwQJP1oVpiETAC1Kddg9YQNh
fARDm5PojAWW1UH4nP3DoXVtBnJtK8Dd1KdxCD8EU2W/k1E6lDkZyTtVRijUJ9qF
r2Owpl435Str1jJdze93frJuiUKzS4U5zn8RQUslT66JwetReixOyuHUQXFvb5Yn
6FSLYn++OJBqAZHiMAt5zC3GDEB5nxatUTmyJSixWQn+/mCH42vx8OjVFRSuyd5n
CSYdUKTuE5TStBqUpVgbHONIPLMI9f8UGdLEEKNZC8k3Gg5UmB+VzT8hbDF4xRsV
CPdTKplAr03VrqHHlN2aH3QUKQVvtnDM02PJrW/VQQLSoLJIiKXIBDZCwI7ReFpn
WAb4T8NYi/i0PQ1o/IbvA4XxAofZC+6nY1IL2GtalVD+eiZ9tenXOkrUmznvMGQQ
kmIropBZ7FykE7DG7xmu1iI4rIZo4eW/BeoUwPJiPuE7Zz5ZeaAiWNbLSmpv1O0Z
2dzpqH6jURXuswOfSzmvNWN+6r+uwjAXzVCr5IMBF5X8bsmaWR2UTv/WZkZVE0tm
m4lyHOdDKoatZqjy1YQSDMcUU8luRmAoQdEMxOA77zNLqMWrYbQMQW/SbqRYIK6l
Nk//Yx8NwXRqskT7mAd+66yIliMejJ77l30m7bPekUvBRNtehnEQKxx8vtNBeycC
uHq3Azxp/Zdya2kGw8KPFfovzU4mcpeu5G8DiGG5C9coUk/X254QPr0tMBkkfRz1
zMygZP++hlQAilqro5ih4FhSdufr2Us9j7aEISIOkDFiSZdL1cEa0lap4BHdwQ/R
RvidSRSkhjTNOAew5L7lbiWYIgtUbDZhkySHZGUlwwlNTUAvDEHvCJW3lbhFbXbp
xHKNYrYbnna4W3iu8wTt5L8ipfg/rjIql/lP64+acZE5EyBX7MracuGtiPZWFhXH
f1AdJAfqCZobDcylm3kQjyQesu28wH6K+wA+mnzcdcjywgz+S1Eq1PnMYV6R9KZn
zTQ90ZZkmzedNEAsFjR8Z6a8yW6YmAGkPTIXhVUIM1RcMIhVjSX+eX98hgD3aZbZ
iTKjnunNOevVi7XIOEDzMR2rO8uRv1Sp7QXhyUP42zxL56LdcTogXglW54joiv70
kev/YpAz7JBLuzhVTnOTovjR7EFvedRjY4uf+CmtvaAk/Ewnvp5kxgbm0hGxbvHP
shLM8ObXRcFvL4cCIq1KbJeDwWFTTp5qhCEhfJ3+XybFoMSoKdklCbxTCYdiG7cc
Rt+aOpPMAmouUykAyD0G1DcArRwLAY8onIj4ngxwtwjH5Mh/t1UYWzd1qkz5uJLC
ZGYIzD2GTmi+irbFF8s3tR3VKeusYAN27Vq+QEv2x0PT3QIe2IVDTtTE9eeFSjzm
ckG5l9/ohCeU+LAqboPt4CGG1q/+5SO+MI2kum9gPOBlIH5ZRrwLqPNxQzXr/+v8
3GeIHhnEaKPBwCxb7S2zRx4kN0wju1tjp6KzxmMT/1X2Mfa5bWxxaZ8gQFvE7DNG
OPcVuNFZX5VHLHvpLoAhuwy4dPH+FjzDtc9UHpCw//rICfQ6b+vFoEgspUwddwf1
qPVtnHJAbW1iXfMApA0zf/5KCFNBDi3KtCg837P3qQ3X1yxIrPixAHqtHMhdRRNL
SSVpWLXLVwJoDIy/OY2qXSuCV3PdTLJrOlT/9UiSefvgqKqhlOvyJDDwvvB565bu
obOlMrx99bf4pkHTR96iG9c/UYsUHAM5Fe0SZAwW4kGoq5bdsSKCziaW4JInQEzm
C1ImhFwowjvmgqWkNSm51wYBWO6VdOFkYpLIpsby3Ti8n2eIy0dgxInmHKGgyz3D
XRO8nVO5QDhkkpb67bR+vrFjXcqngRYpRZ6/8l+4R/lkn3/6296kS+IKOpgZefN7
IpMGWINKOsJr4g11ut/QDODftxhRqrmLP3J0NgQgvXkUbP/H9NJX490K+2Wm88N4
kZ6uCdVXMMmV2DrAlF7otJzXF1SyBX43pxuRTEblV0Bk1u+sn1mJ7+UHl2AnR1KT
54mmp4a8SYSjkxVx2gdEF2zdRcoiA+E+wBjY3YbR6vNxhoDAjj7cBFH3d/DKGh/a
IZSwUFRt8C0tH6qEOqecIUJ26Pk1p1v005DE/kJE7GxwKu4EWO2NLMlxqVh+jPng
hIvg8/XJ76+5C01arWangjOd8MN7lfwe3aztQTmKy6ddMbpYZC1qNwqBIgiIoArm
9EmiXK7EGq/fCLv4jzzPb+Oz/7ifUEH6RLPzJiAGPAL4PbpnrQwduFU+nhM0ieUD
K8xDdJwgC+DQFo76XFfmnnyAksZJBluO34g69P/jj7ZVMAUd+UWGD4jRj8tCnKMW
68oQaEpXPfZ6U/kTe9WfnyNJ10mkW1TrA6xia5waZFgvxAFnBoe/0Fxlf240q8PW
WiPjHhraPp8mVWNk1jwX+/mry54NXF6hU4TpE5ZgixjcTaSt0LpUSr8KsE62FFDo
3TJYyl2aK+s+LVaCDLe5CFo9EqSbUJ/SNQ7UgnIqkWgLXkakl6uGZ+x9d1n901Yn
1vyg32JJqDtnw4WydE6lov7iA1I9MwEX3mUf/QT4I/ARaPRDlTPetaZ2L+YXf9Ih
4l6IBix0g+h5mE/jtkJoqT2o97k5x42VJX3STlZtRm3z0WSxoheJNlHr4FnoE1om
cfAD5Jk7B1agBdOToIJ/6nK18nFEE8Z1yQUFp8dAK7yQQ1CnSKUQOK+zMbpWEiPf
BkerU6OcVi627SZ1I0shouf3SX2t4Ip19xJkkNAPUNpJ+gRpHMk1eDk3LYwnEKK6
7k7OSy84KhSOp2i0RCXYHDgIPj7YQkKj+icfIWyFtGPKK3SvBQo7ZDCVhWeS4rtH
5d3LmA6RjkejunN6iYyXmmm+erqfpaNhajVVnk7q/Xx9OZVmdTKfQY11vooivFyD
JlXfPYvx1eOhWymhCDBtxQW4c9tGHzAfCsa6Sgpzh2PM50VhNilh2Yv+APhTUrTV
Hux8LNJ/NcGioWG4px3hN5jmhTuIhdm5CZmdtPuLJxTKqECIToFBGWicOmfloaEL
zkSwp5xC0e9eNWtacpJxe52B0yqdTyUP4IRYy2gCv7eCW5t3DvFGd1S3OtHUvAse
iBz37FEc8jSp4Ct91tDfNcCN43w7jBEWMzCcz0CZAvXSn1PDnxEqhhbT0/j/NPqR
dj+sZuuhHwg6zr4x+S8EwcsTTZCyFy3xk8w+VO6tNz1HI3XaxqAwYJEpe8RlL9iC
bvrLsrC8VlxuGOWHkr+QweZD+mVChuW3m6PJ4hBHmDRXfgba7apPAiUWdTDAkj9c
X3yHf3h7NgSm4OdE9A3yMZrxaw0MWgMv+LwOmssHpQ1nLDiAIzPQdtp6vouxUPDc
aeYifFYtbWX+YaR7L85JW9Rrn1MARhvM78x76cPx1bGsAcOZTTBAJPlVDQMqcoq3
Z3x1Ntpx4H9RLTcJMdq0lVq7v4Pp6ZpWe/j0DgsnaWoe+79QPFyoV3V7DJbKH/Wa
JnAVOB9kdsQETPBEs2Ac2AxfbjF/5JL7Q0hgJXywu8ubNZIEXyKCRqfnsyWO7enT
kGeuzw3rSF8bkf7EShSn6xO/JsIlZ9TtYW4Wo9WxYOlLVvXRywh88/+sPqoKbL7o
x9vfif4MfzZ22zKbizWD9g/t7QdzWT5Qfxi05euujblNLFcMn63pXGZljOdE6S6N
tARhAchNqjFb/o8DerR6WpEqfkYFQrs9tlpMDNZS/oo3E5rgtQAo3ULGw7YyYVHB
xfz+A4+dJ32S7+CDgnRd4tnhlNM71/zbfViw8mRoeeHMxGbqyVe8pAExbJAr6OB4
maQJ0en0hgxA8nh4WRaU3uSrXEfeFtFm5lOelGfql7CU/MFUFocgQ3pm3fu3OShr
59W4nIUEazy3CjcYRTipD4cKSBNj5Osjn5xL9kEzvBdGYvisjLdFBpjOSL0O6LPP
01q9u1RWSC+uhLqZJQQ1Hm54ZdkFWV8lgyp03mMoHTMlDNGSl0mWF9oX0sLAgkQn
Tj8Pt+/uC5enQeQipPtISUFqb+CsXqjOvTPx7SJMegmlrnVrou8OZ695PZ+m39hw
RYmtKlQP3OQVlLsw7Futo2uJhlQqSzZ0GZ84lZu+PFrKfLrtq4IwpufUNloVvCJ6
+oQnTjUJSJJJQnET+z7HNDkhodzfdGpeNnq7CCT5kFwT5FEDjsISXzP0pfWHYl3A
jL/ghyZqY81jk1gqhmI9vLBtTOj1GLTmcm6JvHewvhgMY0Mrp2iskrVWChFLhvOQ
M8K6RD1v5CGN7KGKabKUCeoL4UiPLxGHqL9ggX8rY5xUlidAXNeXefX5GLMHUuRp
5mF5u7Jz+FLaqJULhJRSou2rBE71k2tG1c4OZC3dFWouGiyrJW5guU0OxyLziXUi
iGecsBIafM8znUg2C2wFNDxAPN1fZW0Ar+SgcWHr3JFrzAoJrfh9jO+12CK/ihKI
eNYr16rcMoOmVNkftezahn+MRcV+Mspa+TNfJ+CHFkQ3UWzQ7Ls9WPbcVfM9gknE
RL6IllhIBE0xmnydr8mL7h3WkxU1UrNRtky6oCOte1lvBBwjmgjearYNZQA9fFHb
FWVUETN8HWaAxAZR7HYxoZD0HcBtRyS52kRRDF3VFUAaDlFogvPBXe2hOwe3gJUq
eMKFVDtG0MU/lfATqHNV6psL0UPTundWGbCo4y/ukPXQGSI7gvm+qdVWBz8LJ+oA
ZMQdVGkynmHieoKbAQzs3p+iWDg7gGJ5mRhYduSsR5x4cxFCs9e9MR4GbMoySHNz
GgmIK845sjvFWYBXdk6A7kc0TeMIEY1SVtbdJ77S2hWYeCEpuDHAr4MuhgSOhd08
m4J0B9yZQaDiePBkEccxOH5LgnqopYYOMt5jPZy1wCN3N8GAd+0dF9Shnrki6v3b
XghtosyI05tMv0PCyyRwFgUycBK9hPiyqefDqPZpZjq6NPX/6RhPuNbre17ypOZ5
2An8GWFVVdjF+HC4hyJYv1yfJa5K7rhQVo5aNSAZrQMjeyCiz6F4BB6nk7279wnI
hlghw1Ty4PCxZcNZXV1wbzmeFeV/hjwU8+kFhHFittxtTDHdQAe1tcaKWMBVhZRZ
I1mwRThVPRM77iW9o9rRBUCZuA86U8xHFJzfhxs28kOJ2uKGLvxJdyuOBvpt4d9G
jWwXhiYkmir+ugwufLDdzRiBuXiGIe6OpPGM0PDX2kOLQMy0pDH+HT4VYakI9WMs
150Y9ye24Jsvy/hadc2/kw/ZvVctUzK8QI0nJbupEA0jjnf/d1axrcO5omNFLVjA
R1HM72C0k3fvJR8r2GH+dRX60Z0MaWDXCGEVA6VBoNF5ciJ3TYHzfEK++CZxfpPk
HFQ9S6RlJdmq4P6SaCZShBIkFZCKKuX6A4HxYLtYZaCJVmqZWR3FWs5JvtD4MJRq
yHhlB8FLgjxbNqZSfwitpmCHILLADYrIUM52Bq+cPIShfiHArTIXUJVlVcPrrYTa
6GCs5NhRid6nODkBJo+Gx7DpNUz404Lj7mYKQr3I+BJ/6Z/UtVGFD6ZvD7uZmolW
3f/6fu7kBeZDUfB1/r19Cjdc/p/JKi/xJjt5912EkGbvHijyAHD1Fo+ShgAkd7tM
l+/Aw8wxCXX2hpHqUTkCY7MOl9GgfQZPwE/i4ajNAFAuHrywAG3QMhjlGH7bSPfN
iHuNTVyEj53XnkOVwiHLW2+LBA8rviRya+tAQEuX1zhygPaQ0TNUqeq+TL9c0GMZ
uz9BOl2vj34Km/slurFMBcn1U/kGsLBdQy+H/ti8+MKCKnmbyIiMg+fjkfw9Qid0
5mwZBdwEzzhmGPOffm8hxX9nVUiV2HN7cViXQcEEOXj01mQUIaqlQ39SLTjxG3Rk
xTA3pwjvVa+uCOcHTH0zjfB6m2trSyRZDbubphiWrJplL9u+/ayQd9rK/o8uoqYk
dxKEtNH14QO5yACyTqFB/V5mXk1sHUzp9UpnXx6rcYnQwSOUZKWohVk+aau+bPnl
0DitvSzWLYeEirjliqV3Kqsq+TxA7DNqWonRk8pBSxirM8EezCfl+t4oWukpBZyu
K8QKxFsIU0I5cpQwC1TWM0e5qPouaubE3adMdWJzO2EwfjlKo5tGiX3GBq/AFam2
wt9nTMrUlIcD9A9vcZmkyymX5NXkU1Ye2SDykHrVHWtL8Ra1c47Zbr5y9H0zhK/a
Tx4tLueZjFF05r/gjnn+4JcrndRp7I51MIRZetZ621qRMVy5H7BnXuT0ud4P4nlK
pd2Inzjysn2fHVd2It/sZC6Q6LEbpjnYGAG/tMcSKi0JuligKRjzmfXRkMSFcqOi
1D42Edn4h6fk5XToOURdROMolMdSMrD+ghmZpL9dDuXX87UAmHUTr7paIaHd5QDK
JgNzv6xZk1HX9l/JMenZdbI8PciaVlfRnLlPLazbASlacQGnbbczDGSZfMO6ZbRa
ebuSF9MDWMg4gRt+hn0b+V0br5qO05AalMY6+LntxMrjt4BRSNm9tqvol4tLXQni
B1kKGr2WtPUZa/Vbq0SseodaXPehJVZZUSAihMED9LGkSIUP8wZCB8aMoAVO0OY6
R1vBdDB/uguhtaU/FnNyEdBZpAjBzVJrz2xk/Qd7EBhtsBEeAxB3fE4gPcDh1MGp
QoQhmZNW1GzRzX7x3P2j2tAl06cPEwd7AUu8Zje5PxTTlLDHp5HHUxX15TwDvQF9
bIpJo/UJ5iUvjssaPcIxow9yofKQNEOLhmpVNOErGAzM1nM1pg1KYzFrF/AvSyTp
AoFpIq4pQyeSOAgRGkxUbnt4a97oDofUyjPHUGp5jAT4oiLxIy/ikpF2tXpRzia5
ou8qNdycS/3C490lvsJWEBlwQKuJJt6ZeBcKspElDKHk1vjBLAKMgcbcSay62Pzc
00kbekU5vVimWyHJmF2NeOZEMwUD1gIPajrIWl8YXotFcjiKlXo/zWzxZiQUpnJn
ZGbKOudWEDDQDyQa/KrDLr3NgONC8GhDR6op9JAtW/MdNKSsrOWaZ7sGgb5YwEt2
eBQzbpLmA6Wqk4q8MsicuVdzzWpjrCN4cWgMsuCQ/qhxgW+/3KcGClZudDHeEv6e
7/lTp85D+AXSxa3/qyzjlZCmuMs500espznPhi71YSVGJC+4T+fYJ2ycNEA/HsNO
wC37mq8HNC1U0nE1jLJXBubh6v7sdq9AIZjrkjSaPLkurLTxgfAnERle8VddhceM
LsLlP+/ZBIP8XrwGxnXgOflsKk49SxV1C2QA6nGX0OgvTZYajWzkR/HiAyJZTI7R
6QO98K17wcnjJjzlbxBBhJG6Ycj6yzZ0NJRjUrubuxcths3d0k1YigSuJz8U0LFU
iF9FAbLxzeFDYbJO43xE2x1vwMqmkJRvMGFosyhDcY6M5pDRAN28BqqA6heBcy+S
Dqv+sVvDxxunizRqz1kud3mNFKL1ZDZiddGdCOoWBWuQ6Sx8nYhLHdg0TJo/bKPR
XehxWzs5huClPdD+MD3FT5Rjq/3qmhPWjMN2OwfQukhWXYKCqzVz7o9psgZdjO8x
pRhJFcU11GUhwn0fG/q2VGX8Amc1IfddTcwjr+jTZWIc2BeIWw0EfevZEEVqyaMC
3uPxxk2+pyKH97z73B1IIhUiW0iFNyfp6SzKCh2mYFPHWRzGVD9PDTwgnfK5FMS6
yfTo692JeNeyVgOYQ8Mf7GwLPnkXQ7ufEeK56a9ndM+2P17YUJWF9D73MY63GXGl
VbXhbGgaer2u5XjEbRq0v82jPrW+acJplUnsFDDKnLga60C/kH2wnQIwYnBqulbs
pkcGQNMCNqkyNIxtI5Hw3zGbZHN2Lwc526aP0Leip4rHAf/tElVxHPcPL7z6pDdP
Gr1wna2xvRObtPXTVFsix7v5NALtNOlMwTvRcZqdnDCNXaimUOfwaa0omfEh9wHO
8PgAi1B50clFC1/N2lvMlFp49nP2XlexuePVO8xU/7bPPvMEhO+PYBav5ctYLj2z
65Et5iMhvfGm9Yw8XnABHYPMaTY6kTt3yh8o5i55R4B4OUgWn2tL8VtncQb51bwS
jRLfIGUejv/apEnpTFoGBA2UZVc1FCELyS5OO4CWxU/Rg1i+JPlOVSMNc9TZlKqd
GTzTq5eTm8bqTxNhL2fhIlbGYuKlQCeVM7Xv0lthEywKfGK2cCcaDWTizNSa4kmK
ajzjyzZQ8Lexb58eTuj8aEH2PBbIlSB88cltIq89Q580uxrBtTd/W076fKmidgji
ZLqlKB/rdLE1f5Y36JQbvGf74lybS55c0H/GMEGJ0CLv8UVk+rk0f0ucBCRZVJDI
gXbLBG8ppfsFGMrAgetV8U21eR6XmT8SzC6dtuC+/4jamiEIGQTdRy034GyhEvVh
HvsEyqueDsouBbdcjdIHTztO1mv1VbdKS9JbTxyXhvPjs+T2R50BY+AnZBI/PjG7
tATBxJwTDPqJ7D0eKPBzVcULjsxyGYRwrBunfrc4BfNkdIxSdtdgitYSIz4LcxaT
RYlL4xpkV4DGcLyAF6StA3hluChpkPO+g+qFTy98YwCXKMFy0R75Zkkj6iazvI4D
gmgg6TV7ipwvOCymcYBIeP2sP5PC32m1WXHJMqdjkutBbR1Nq1UbvKJL/AJ4SXdM
l1p57AisUZ/+PHwPnvagpQGVd3obiVNNVDx/yE61hjZ+jhS0IrtPIr9UzNc933BZ
YFR4og6vCR01RipXqrMivaRDCL2yhqUvh+eDrDjeyd8xazf1kCVu1xW3T3ftfC/y
geSJeYoayDbGKk2xX89qaqUdZxVd3pBkjVH1LPh67vavhbnUKy3oJPRKRg7Lm4tR
5DipCM6JZUJq9CemIIgt9QK8wSMXL+7ymdlQNmfPrkpNEA7EzAufJ30hey0hVh8g
bQOdNwg4W4gAgrgtV4AF5xta7iBMr5VfaatAfUCfZx9PK9QpUhvAuYtbK08u3Glv
EaOeEGd85yr7x/VhExlWOOpEIwCNqgcc150tM4Uz5mEAVMZhBz0PXLdJc4dQyxC/
QrH13KAZdTgaKTjl4su+fAzZPMLmd7fuvYzY3DTjzFc5CDEYG2DBYs7YRpVi5uZF
zYVYgAHaEplsACnlg2xXH2/T37QQ5wYJYo9lmXbDfqiDXf3aNJEl17Vx/LVMCBPp
M2PPz4aZTkkOfTq2yxpdTxvZ73W4DwKpauDC+mJBUEhMP2oU2+mJoIDpEydI7qMY
8lk5rE2AuFx+JpVJoe4vGMqEYPYcd9d0ITdRQb8EKvt3w9kR7Cxk8omhqVToq9zw
y4lebZTvmcWbEP/dnpzwRmg5H1kgFFk+cT9wUwHmXPO6AQaNB+jIZImFVvc+KURi
Kk5c2rgZH47ED9pgTu90McSUFrbeePNevq2c4Vfp/vbWFxNMUqNzbC2cPIu+Wr4p
HE51mMa8aC/SSC8/8QkgasCN1vb83Pxv8NVzU+GUAmf3OpdrWa+8u8CKNBfACFWa
3irpzBgnQsgJ1sd3l2ThWOPBGLQAOkTgYQeyQ6FhuJ2HXUBPdrparSEQ080hwl4S
oCmX5GI9Ltk86qLtbe0Ri0/20Xo5dsyj7l/DhBhW3/zMgFmIvhMyi9MrIWVDvaKx
ZtpglNo5XWrgadWZ1HYZQtNxSrIqpFa5qU09zJghbP2fLukZzh84u9eExtXFv+hf
TRsp7WYuCDWeS9pDufIdzhDQXXqsHst+XnpI/C8/dca0Gsn3tZVwv//5WA49SoR0
KJ26TPnw9tlulj72wkUfibORvUM1tcgJy/6SeDdhHzF+B7BrGM9dXe7cGc+22e+C
GZC5rpsFcOcnuQcIq/9FXfORilhn0ryi7qBRBj/LDTerG+5raQSvOqcTYtHsZ4EO
iLaPqCk2SagoWbT4RSbJvbnMCCNZlZvFjMXB5EA0UW6+H4xpE1uUX2XQmQXadI3L
Uc1oZqvGYrn8jCyvYyKzXibTy7HtLzuOa6LJwxQzy35BWk60s3s2QdnZxrxL2Shm
imz28cTxtv04fxAhRGr7h7j3VIM3tytvwAUmeohBbIMGyihGIe+8lyKhdTPm8x1A
Bmw+0aQ0p9kCzkMkiQRJyvdPqN9SmuqqROi6gOOGKBvfI4xf2H+csNKktFioNkyO
MImD5/S/UJualhCHvddPDDRyq9uKHfVXReaAwgUgd3QKnvXW1H1ka+lS2zngk2L2
m+JmAqirie/I5YRjJeAM+fbvBhiYDgR46xqptOCOssq71g4Jrcemkqilxehk3ur0
rvy/LVd1QavcWKNicPhATnuUHKPotAEgq70Y5N4VOnt/KBxcXH4EnnhpivFepo0s
vqYbIZtGpNklEFqjglhLZZKoSYOfFDKdtRYHSoZ/2I22YpZeB7KsqDX+uxQBtbsF
XxteeF5Z2zvOrB1oDSbYEha7kTSnk0uA2LiX3wRIYyaBdi8dV9f6bcwAJrNv+QFs
6JLKN0pjvbg43EQL4SAS0fE0zor+Bk0/Rl/bO1DHKH5tgbzp1e/jFaxzsmikz5LK
ljzSzRIfSR1YEWb1GET10oT3PlmHCg4dqV6iYvD2KTJIqNSZwuwGZ5PKV3SI7mYb
COZU99tkBHNX7cWJMzjUbzb0DDWtYyRQ4339AWEz6c1xG9NvKbLajkDUX4GU+mZA
KJOYI2+DK5QoI33d3lJsoJmTesvnbaNYJwikEUpDXn9RpLVgMRJHPhnsFZ5z2O7p
uVLB3zO/yrPZpYadV5cdOHQHMjJdfteG1kpZAxYI9xmEmoNHp44rfrKLHSKjj0IK
TafSp6QYzJWZi2kJ2lxNtT5yCiKMhG44jmR5pVj1RSJ6wYkxMhByc8TQI3oteA6V
mqh/c+5OPv+34l1J2AeoTySiRJKKAiaHsCCfgiZEmZ/X4w1sDKrK/1Lr5Z8uuHP0
8yYmzHlUWm9NlcRDPcLYNCb7kO9DSVIGdFeocP6b/BqcwMb0yLV3Uc9E8Ii7r54N
OjnGcMvSOB7bFVOa4rz2NvhH80n36a0nTIiuKN8TVg9lD/alym9uNAC1ZID8c9/D
23cA3X5jqbqVJIhIoeewsm0X0mrWhVtciv8wj399rdUqhjnXSnwoGmu6+x5zeUuF
a37Q4Ln+lge/3P4P58ESvT99MAk7+9lcuQk4WPb8YiNuw/geJ0cYs5c+05bhGHAK
syro0vYaVcpYYolz2QbOTTHxkkMfF61WHzVWoZi4cZYVUBSQtR96cAeAbLc3YxxP
WWLL71kk3HfG5B7whdle4erOPoOkWVs6YR/fTazn305EPxDSpEjCUcvdRgEZGEmL
qdBr6WI2VHdfEh23nj5PhbfqsAFZr1NY7jvNtzoOroLkg2TVieJ+Hwn1lsYUu/ia
pu1MO6ousU2OsNnvJWkNtMaKVLprA6pEg8OmnULKZFmnNuFzrLZbozoVSFikLwWK
BxZCbTq1MOsQ/uLr8Zr004ScLBAUy33adhtPGH3C5IL5vqAQwfWtLF5ChSWdXQfY
iVsHUA7aOBbiAL8mIHtXXWLDWsCpqoHyJdaj8+iLaa3tBEc7lk+5H6lWGSMHfCtT
/ma8sHVzNlZNQrjdaD9PiNfMXIMXWc2m+96mDowPeBplSodfv6dUb/Z7WwlABWne
yWfEkSR2wHH5VOaaZ1uh/3KQi6ldyGZk3vm3FnN2d54/EakLqJleODov3sgTULvK
3NqW4xL9N7tvSzTHLS7S109/K2By7/p97m3mEu48pmj/aZAmLStQgOAdS5dscsys
eTKQDmZ2OviPgqPbxF6R3mM6BmCcQxdQJE7R+4w3L9uBjQL5X+DVWYPV3nUE781n
aPTym3r6yYh82TF5X/D56h2AAiTu35mbQFcplKuXAp1UqITHYBomnX4zlQ5fB22l
a1w0uxmScJp9bUQ3fQoDdDAmPsrIZFsTeP0MaqPGcfWfOuejQVYolpT/aVPBtoz2
svPoK7tHZDDb6xMf5oklv2QqquYVkb36GeXzhjn9OU8SjkWSOgtBpQ+EyKF1RxSm
7DfT1gTxqgbqd0k2tzia4V6To0uStrF7cb47yUzb53Ff94Mehb/t0mKHJyi2ps+a
jFyiC0aTEiMSX/1dm4s+Q46xjR9f11R4K5TBV38B/IxpfTi+8TfI7ilqz0a92Uoy
qSbzS1roeYu8XiU4EVN/dj9yCwh+sx1BstbZSwhRc7nLVaVvBnROeKf/emze9Eer
Hmwm5XekBkCFhGC3HfxxGJjLIW3Lcj5azH5hs+8x6tIk4ifDKSerAlCuyj5iiq7r
PPgl9RYonQrsSYrzS2Bf8aFR2Ek1ykdtp7hezvN4DcErEGdCxzYNl+s2AZNotyFf
M72lq0T/mrPEc74LkMN1AXAsZKGGTi4Tg+SP+/nQIHerjaVcTMC/hu1Ff3+3oY5Y
Pb2Fa9Zi+dZ5hkUinjlj4G643j3FMPNk66H5rtiCmsopbzM6BvEEnw6I46Ull/FP
yiq6pW4L9fp9KeOdKP0p4U++nM+kMLUk9x/p8dkKGw/9g2YW7DPjA2HcKIwB6OAJ
DTGgjXovOUvDfIu0pjWmgcKw0Hp8hMDtkyBTndc3MIRgEFnuATLJA2dHcRQvz6uO
X20M3wzT7BNqQ/bYUjbfGZ5FIrbjifx5RgrmOfR5/cQAtLhdUTX1mjT8IHW0j8U7
3jYlgbHUuCvpBCcu+cgq/QmA1kkDBDJWY3vCoZTUzj8atlJg68XZdDHEuCwbfZfR
XuMKREzuqOTL3k7F4ZT+1i0Z7vBWMhoaODiiZqpnNHuelwXc7m703SIEJoPRXzNb
Zr65OV6rWKShL/59hgAZn10Hp4vb3UKVoGfrJUbjKNlWntYjmBf90UCrc86p5n3n
kiBFqCFZunRmE0UMIZiWIJ6vKru7v/gxSqSnMbmxMhNtAkV5VNVYDcmQZ3+hlgk7
toFyQgZ4xlK3sMOEYrw86BRGnkEnv3gh9wAtezSyf9wiB+AK0FYVvLKO1ATvydjP
R32fG7Afvs31WmEygR+QLRhE6NZlhfCDxgXqsm7fA6DKoISxYL+78TBGRBvp6ZfC
5jd/L/IpdAsfHbUItSj88r689Q1f5vt49vX3ahnEsek84sukpy1f872p+R37kKhF
iU6EYtjMKJL6KirihsfAgLW5Xx7lUOA35WkwCv2XopPrqVS14osNd6LMMCwwIVOa
AuFPMzHIja3fCOKxERGZwx/8nn3Wz3UeEgjVI13hZBT8VnPetMC0Nv9tLTzFIYsN
1iK9kI9tDBQ2mnXg6deJ+WwEgmuyxMe21WPtbESgPLwNtReNtnPSmwtTW04sEzHs
UjXTLCgRjyqDhYT8O+NkJT6CYfyYpsgkCo1EQxMcwskpNyDpSw9LJDYKFr0/zm5u
L1mHhZZYn6O97kd4+5/tYirOCqJFHn/Di5cUNAQ+5H7JeXTrlk8hoqKiaZqRoRQ/
/DlnYHE+CRQcv4Q7/tPhQx7P+9j4e5H8bl/eRlPjj3nrbDq7PK//dk2mD2ABDDZa
g+TIFTH+H0tTVz2SQepYW7HjQRIb4Y+dEzbtXAS08MDSVU9aQbaFJHM77VBlCJO0
HugrmmnJaiWYZoHCZQPX4ybtThahfNqXGWx0i6Q1P3TPHu1/OhrlMOyEemrv8XWl
YP1XHSkYOdEwx+5GmiK7FZxY+8/3f9AS/AEJKR856PtzHAFWmhWLRdHEhrFHGnHB
k2UAVqtfmwG8xmP6QB6nzYcIFFhERExnT5Pu/15DK5GN0diHtw6neCa7M8ehUVFh
kMzok/0ZR0vWCTePK96vI+aiuoP682A4vKp/5Yue1pZ2ELTb7We3Sh0Uf+KdU6L/
/Ba2aOmnEuYxDsHK4NZE9T7zyMSDlpGY9LpV812L9xwGhJblLZ4Xw+bcjQhWa2+s
Hh659bCMlJUvz6FhmFRR7Q8M8IA5M+4S5+XevcvQDkaAKIttYJf2Fp63S661BXC2
bKZg/LXKR4Wq35znvf7L17LSGJDu95D9WT0kCojHreC9dpxBZGJkQbpTz0x09C33
o6+mT3kSlHZZvM2ep/kvpPhw2PM37OlfJck7kxzF56EF5c9iS2Y7+h+2Ho53LkXz
sfo/fKHRDQ+ouhiUfKXC96nOz2HGbZ4NPLYM1yVDrwq7JukrRoRYSpTrKgKggIWs
W1YbgFvrtBq6+SzF3oAOwLKGhSVwZHqun3ucdQZ7n0/7VHa90NrxTBDmArhfcVoU
8T2LeK2NXtypa9vAS2gI8qCLB47BKpcuANtbPQJSFxDn7ZNSgSxHkRq0YBD/GnB8
pE3Z5SILNM1mN8X4vbHp6n9nrdX8P9sEf97XjZ/muqg2R5T7GWGk88nBqtkmWQ+V
3pXWdg+LNVRiecILCzLGPZAT5WsO5j4CueB603CRDzUDUPgNOmsJ3AzZwgOSPnS0
wpxvk8oL9K+3wOr1jY+4FDcVX4IDvPB7DXddR/2vQKCnO3Tv1I8Fc6N15Q5T774I
mNIclPA/7qQqBwdc2CFimO/8X2LkJxOiTu+3rrKWw/l9e0JOpc8xznYPT/EV7jZ+
FiYSUhoxprxdSmFoiCbHeWSz2R807zzm8ZhIQyNfpvBXrFJ+luv6I2v8cauOq8+y
Q8hARPe2bNP6yrqZxCZfZHcanxoZZw1lHnK0P2WYJkyPsd01Fxt8VJKdJ/d/S8XB
qpews1CAM6K/09KuyfD3gx2AjnZn/HVSOy3GP1W37V1o1F0kBB5v+qMHV3pn5c6X
Uv19XDdI5q9H+NgQREpQUTZTgwewCgpdlWxuVNALA3p2Y8oQkM2tmvcrjOrZJopg
/EGsXHcQABJ68DzBpQiFwWjtrk9TMZtkHiloqRW++LVAH6AQIvf7LQNy/eNIYeFA
aEcJWA6pcErF2wxghmQ28X+bkKXLghrn9ZCUAGUKROmeavKI4w0j0+WWAvEx99CD
UU4AhdP2QdKqO9unwjGmgE4SaStW7/0QnyPb60DQ3NGzl7qPXCNUmlxYyFqlGiSA
6SHbh2oEgkGcWvm3c/7yHoeC4JlviECwGwyvGPxOU1hJ7uA24jltutwJCEQ2aQhl
XaY7LI1c5zTZJrrReFoBOUYeOhHkmmPVJqIdZdG31Hv1HHYi42sOApLE4eaq79g3
Fowvye/bUEfyYF2kCNCr+AO+8/P8uNT17zxfY9XbfutKveX0dtXS9EEk+IUVDmcR
HlwDfni9WNhZskIvHAuJqMgS9Q+Ing5CQQTb0gc0lrE2lq6jj1cRZwrsF3Y07wye
qviqDUNVjCLxBArCCSgpIqTKDR+b7e1gT5O3MBGxpsMgiXTm6bOBRc5RFhijmccK
DaHdSB94vNwP72gV4yKXiQImDzTpcsEhCN5WtU8iXzwB+youuEjPYtXyY8gFGHXz
SRzC6TEVBCfTpOOzyaIaOeHx7nOWwxsYI5vwgw3M+Dd650Ga2pW0y1yPbYeDn3UP
+5qLTYFSOnHPhwmZEK/Cx1BrGRTyt2tMI8JNn/SwbQoU1h19qpmx6pKlPf4M3+e0
FBky1Bg+bgFi9K4NePGM/czGbvTa0PtS6/4EeiN+Wl08vaXMUtDDqpSlPkh0J5b2
KN1jjfuQZutk3xGg8IZ8ryLQJMhK9U/+h1O8Or9EWIcax8uQOoiVQ/H3Gt8ZLjl8
8IQBcRo3A9Q2Au4hWZgaLjYDtEUdgmxWsPkZlX5LxYwBViLilJLXALXhkjgYY4JQ
xJ5141xCtM9r/fMRPzVGxGJ/UwQxlUrhGVgJosx7JXwoJ6A+6stiQ0FAezcRW5EG
obnElFWVeVZvu8XZLpgKsqP9EpPWEV9mKn6uMkNUxH/0wR4VpmttYpTuE6mSOPvl
pYELdRxQThB1Q7SCr6TDBiB4c8XsCiN1R+SxOxBVENP+2Wu/yTE5CnNbpQTRlZNE
JkmYPnVYMR/D0hfOG6zw+3ef7npwzyeguEIEGU1TMAHjYyyNVdLfTifYnVchGnzi
HZo2XSSJ/GKgFsUSXefogCsLhuPpKi7FfGSe/hM5MSfKHy4EvnM3OBTzc/SSR08F
KuD4zgdWDBT8ePDYW6ZAerVN7fqRo5yupSee0wQk6E8lp+o6hBKScV+aP6vb06jH
qsM/5sSwx2wMdOa6LrFxrPkfmnwNhNt6Q4FxNd6ca0wAdnPFREq2QwHpHEeKh6rz
uSonvDr94fvrrXnEBiNadOiWP8GRAOjM8T7b/O0p03dTkh2hTql8XyamQCJ2htG7
uZYEBKCXmuA2tdF5NpsE2ogk/VuUw/W4iGBIyh+jsApnrr0y5jpWzQJrCna7D2qD
+qyXT6ntR5sa8Q3RoS6LaBp01ACm3h4pXzDzhXZYBVv9d0ed0Clqz8Aqrrozrcab
8QVqLGccL0nm1TMixGxJ4Gano04Sw9WBDtQDSOTry8JyFkI6mFg4WpozTrM+qaCR
AbdVqVgZ4NqL688Y3MnvqtHpunAOt5pVh4oT4HXuMLI/5kILtcktVhr16fzaXESS
OASoiQXV1dRr0fM7POjZvBlzDD/6BjXieV2zIN195evwnrRYPjbYIHvnU0fZ20PE
kh9oEn3ZyXQqEZuldN94H+BY3dUFuyWgqFERmD+lu0ykfiIe6CuvY1POfNJtBlyS
aSUtKlS77Dm4Xne7ecnes5JFrxs6DhU9y48IRiG55JencOA4J4yIIF/qLD9LPTQ6
1wSJoCv9vgbvv7R5rZApn6OlXMIaBiEsGcr+miGfXwYrZmF8lhMmFvxDlFBJXcKo
7YwOAa7obJyllN4tUVXCZO1+w60vCoUPLaTvFMZzJtkvCtbiWlSLdZ+9GJaa1eU1
mY/1vviYtgVWbP3UStSylTWUffiW5N/x3nJ4p+cgPg5gJ0X4ZWPX6sp3XAeJleMK
fKwnR45GEOlw/phy8DZMY60gx2SnyPMnTIQ0klCTOX3nGDzvONwzRsrP/5CtIwQl
QM7bojwsQZjGSvWjiwUoYtUHywgPEVcYpR7IpRewcoEWjTXUORRfTZE43t/6HIp8
frb9Y1y4dcFNwpGwL+NGN5B/ELl21VFjM/w8g3wPvEuDlWG/ukX9QncEfTWvFhQg
Vlweva1ky92dC8CRL1Dxvoa9Btc0IGT+Y0BPPzljUpwREFGKkHPVB+gRjx4qidm1
3z9542ie7g6piKQxDFLpwQKq8HCap4ci64cAO34O9eSorN+DxpgH2Mjl6XrMFcWT
8RPyQCGx4vNQ+oBDidBnjmmYtUwc8ovFhRnLb5UMc9hBi76wHhi8w5Ifi8jzpEoG
If9pRmhyaM+yJNpXHIlMxD7OwHg2Fkax3o72pQQAx2QPOqtlJbVpZ17eWbO34Xav
bcUNz5/aVi+f6ZzXBjgPU7DHtOY7REp6x0jS7B5g9wc2N+XIWtoDBM6SGUk8lwpW
yCU96Kp/9MnoB4om6C+HGJmRnrfVrlzrJcz9wdWhm5vc4sLZO7uJupSN73547vMl
wUX65VkvSIih/3tTzDFK3u6RP2HVhbQLUo9PKg6UvveCQ1qrQqzUS1WDS6YauAIY
NzIejF1zjNu3fPyAz/hpPFJ9Kra0yl6pdrMxxELWLFNxM0PsQrXNXJQsBi8EU6E0
BSZQNtl01FFSHFcuSAOYTLYLGegwxUgjkZjwU75p/Gi20Gs1lDEDN6yYfOsMfEji
BQI+ke4oauao8YE0IrIvD0lUEeR7B1fty4ObnFsv97xU0P17dX5M9FTmhvmFa00y
2xRe1jJevwG2KAIwBY/ce0qJl7keaQv/POHE5hFsgcUZm70SQkChLLCrQAjZElwU
Zw0KsI3v/j3JoBdgUFhp1qZXLE4fWivJPTfdS0FIkENWPJJi8CIDPcVqhjNp40vy
Tq2MlG3QDndzOpDc2mO3j0XlhKd0athCVL5L2rffGB55q73hk27/vZ6yNZ5unthD
i5naWvLKGeW0B1MFMLl606bo55v7w6EKB9xg5bjVWQlS43sagUJPa8DXshwv2AXj
fU7HokEs+J469hyQtAbn4gvjwNGphCq7w+pRkQkopxztDdPVt+8XGNBglmIs7kqS
M+X4RHd+aOJzoa1dUVRPaVPl/DVX7OydDKXKlpuOhhcLHQoft+7cowl1l9sTQ00H
wCPmbONg5jzTY8ZfOZZ6bI87LXa+ynysXXmQ8jCXFJ8rnp2k8GfnQJLE8YGCI4/L
r9a7n1L/ePdNgLDibKdBeLF2OR/g3ejjK5F8JTS7sHyWn3aFsc3EjIDLV6Fu1nTi
hGRJ6qZ8rtvSVwYmy4XycYU3EfAUwIPpRjxIynXP3kH1R8NsK2//Fj4rfthp5W/t
6AM6keZ8rlMzJtfm45z1FQt48II6RE0Xss9CoVA/A/o3B6BLgHgiSfs2QxBmzNX1
kwM0CsN0c9EJMwmlfSa2bz7wGhCtkPpD+pFVNEOuL3b5eoyPBbvweuVCU2SW8RTk
5ToJ9wJLwr7wU8eZ90zYbr8HyODYj9a4nRnGCDNL+AK9/WZ0cEEz2U4OEjRtFkjC
vci0AxbPMQuI+J+UbofwL9zyTDtpdYB/sU8ZN0JqsS1vmdXedx38e4wBv35cO+Sy
5hsrsRgD9adMT+tOTmc6BzniPl026B+yIVapGfCVW/nTH9jf/5zjEgATdRlu/xCj
7KijH7Vmyb5r/XVK/c1s0fdwadDEhrIX6/IzE3saN7M1LfqBC2NqhUJI4vcnwWia
spQCo4t5aOKdDzCCQGr7bl6b9lGi6XtA93IO9FHxZ9unQHgyOc9mqQUe62a0DFq2
Yzl1R5XAI+CbV4cile/f1AlZEqMKolGR7WZuapy61IJd4Xg+d9401TswdXAHupDc
d2XtdLNEs2fiTTKoCgDjBtieku2+Kd0sUcoxokFHQPXB1alukwCIr/I9M11TI+ZI
pWLMKG+Hi6s10LE0VnMwyTv+T+RJhp00o2d5r04xP0PLaOXYHcf3aorwp4jAW4nr
zyLMJijiOdzbJy9KVaIa1tvwk4ck0A6v5QvGV3ZaSajjGsP4XbaZ8Q7zDaggO/d7
yN5fOaUjxP9C0FGR9hcMAUG/iUVorMKnUOZyB3CvgrnWF2BwajoKFMbl6rsjHC8R
OyADVHGRCqKtEkhpQ8ondd3QNy1qcPGp6goAAK4AWLpukyNEyhA2diKMoz0hA85i
UkA0RWsZ4wN2kt8XAA25vfqHZUYSu3/ag5hLrFEhMNczgRzWOrR639GKlGwAKnx+
vPTRikidsSkk5zySwM3GNnvCApDBDyAjWTYlXEbrqFPXns6/YBHVdyiO/Otd7j/E
3pSIvo8/O667Hk5dTSOys5w6Yt4tOpkloIm+oSDeYFUQlxsVKWhYC34P7nB1Ycoc
0bws+t+hJpMGgN47EZpE11E2dnL0KsqAk5VliwBHRlgdU6xy/d38LXrIENAMrNGy
esGfrwFOoHue1XlusZAhyuE6eLUZIfXlAiR31Mi9E3M2+UBH/wollL7DdftZVfdl
pOyEtYyCMW1HrWSlkVK1GeTdsfml5loUhf5dqL/Zry5Fab74xap5ClcaLZ2mqCd6
fZoTzWuVxv95cZe/Xhiy+Wp2tGICAfpb3mvi/g7qWRXUMvnVMvWJfiKNV5vPGhn2
JCcg6TjkiIgO/wnE7zVsUUwkQVBjmE4K8rJ6zkm81U8cRx5KwrzJZjiclwY4mKs4
FD7snVBl6kc3k3xWTV1cQs71gyTO4ArNMJAQayTrKSG8yT7Vgzli1idSm9qKMmd4
4iIi3zU1RpOc7RPi62w8S1Z9rVbQZN4mEy/sXIAYhMYimjVnOuIKaunFexXaeHiZ
0EFMmbxFYWHXvinad0upwQvOzCcbw5mlvrRVdCcmnGKFGIEbIaG7gOgcxAYnhfuV
vLIQqBkc8sHLREcq76uKnO5yLeYXRyNXFc8yNVmn5yJMq084UEKtziKGqJaWLsqv
Rj5C0EyivD6wMmhXRAWZC54RUiFrPwjjTJspJlapPf2rElQH+u8+a4NfgcSOatAe
KRLeVGr6fHVitHmqpfaQIG33Yt3BADwdTBbBm/FwwXZGw0sgp7e2x7n1su+sjjP5
vsSyOUoypO1VbWP42AhgnhPv904GCt2ZTG7Xh7PtgxfvfvRNvYDalyrVfXislpro
+JdFAjTx/DiXcvjew3tNRrsJhkhs4oC8QKTOW4N/vpc9zuPLsaJJwqkbiiqJHo46
MSHZZX1dQwAcvDLYJo0sHSKitDSMzb927/RCLdFSSps8I1qygMTc2HWlpASCGYGv
R7DnSaS3oqdXZwqAlLf3EQERxdfjZ6u1ggEstDom1FOY/BavjG14W3q0Tdv4Xijm
Nu1y9v2nX95DjzDtCooRqXVSUn8p3dwQ5uRPD39uIq3BCc8MWAoQha6/cSvJPbJW
P7ZtVrC7HNQe13ogDdqyE2a+soDiJBUBl9c3YSSvpmfNk37GqPLkfAESjSXi8Qhi
UF01VeK37WC2ieJayq3vo3se/5P6ltGYYUKuMbGlRF0omTrHa6zbVPQ6kIKc1A1T
ncTxuD5ALzDf5v049nui4F+vaDN06pmcHOlDoElJdJ5YE+kW0pFj0KOfRIpb6CVe
+eZwKPSQMRS4Vw9U1zEnJPEAhJli1a+CngkNzAIfJuBCItkLSolgZt0bsA4g96tJ
HvWAUIu4d++KywAjcHGl0TOuCK6ORu5AZs948vJabQYsYbdqCBZEgkJCNlRFcYPu
djQxdIy0Pu/ZvsWQORfN7FhPzed/YM2V+7GFkAOfIruAAGfuYVWjlcO7mqRVla/1
aNaoEdX1QYTpzPPn9+nI63ucALNzH/OF40GGQ91pxdaFuZw21DcSPvAX4Oh56ApT
4miiWHDKM1o/cbHfBtjXjrHZUokDvSAAq43RhcdwUDLIwFO7nuyA7wkIXHbI6Eel
krTw7vIIV2Gh8DACHyvhvyVJ+nhvmrP4IwSy1pSQ6clmwjjSBnKHZfFM3YPnRQAj
oLRknzrdksl8n0BbCuehGtTS0Y0iNSY9hDVWGcN0yJFt0JFpYVmFa3t3OTJ6E/kh
AaoiPrZN9C7zHPyGEslXlmD8kB22uOOTSfG1rhQUAfJIbFl/ows/R9nQwp0jM7oA
4uMMaXKkWWhDkDobI48U40r0fGBWK1ANb2VGYy3rHmdWPH0uXOM1U6ul5EYz5fAn
sG6Lj/DGxRCeFfenh6aJ9xraVv5a81pL50GkASncUVMRnG7ORpHIyzv7Viq+0rTl
pXLIhgJZYS5Ek7YY+q7yf+cuyRm3vZgx5BGIW6fODWdvBBaR3PBaRBkm6OSGuURX
BA+DgogMKzx1byBApuh4HmIByfgvW8PMqEiIQDXkzcLXb8pYLny/i+G5rbfg8TdD
bzlMTU+/pOzqsa48f/OCeXstBxEqgOOvX6nrjdzaOUPujRd/tShl4zj9h3W+6Hv8
BH2N391tZgTqkQ3YFTDRLnH77m2ppJvTVdL4YalOLQXdAAdfzo7L5KQMRS4AJfAE
3Ms8o4Kdr7jtBtIx1OLUPmLX6Myl5SuA8V1ktFQD3M2w/mbFaSdwDYKhjkhd/nZE
OXDqUwNxsGY41ipzFHipFKJujynI9qT3Ok/s3zWkIeEDcsjiaHP8VTmWDyyJEvo9
dnV7U2Wo22bDLwSQ6b384xug1HXsECf1UN+Cg3FL5OTcFlq2oh6gWIuGYSkwIgmD
SMtATcR+d2hOOonYbwc1WiPvFPwghmCEZSeO1e959v9Ne3NB1oKDoLnGtk3UIrYW
GQ5cjJhfUo9+PscjCTTjVyOQufyif0hVQxMYQzNT9nYwdfgsmbINsUeGJWlxq7Y5
e1Amo7lWSVb8PYpZqkzpp5StzX0gvs2h1WHafYXFc7EzhLHyhRJymvd2ZWTwNTeQ
IpMPxgxRyodsuGHyp5NFAyanm4YgKIiUt2uqhbdPBP2dNbVhVJvO0tFkwxXNVC1Y
5DtwH1D+b7YiZdwXe6UAkhHjmc1rPdxjMG92Oq5S3p2ksC3ghPOK+8E655G3OM1b
+4VO/qAHSix5MgRvtA0W8382W52UlOxcJk0WNaesvXxW3U3SO1TYSCGqcqlQrTsY
zyYZdqzn0hEEqiCr4bHrne10Nc+x2xSj+qc5yHQkcTsvtAQarNFR7XTG3CXfAR3b
me4CLjokYkTLeKIMr513ebmbYCyFIaMocVlABQtTbOWzeRpCnBGtUfUoVXRk0Ipo
x2AEIREQluRGBFNOJZAsPNwEVtsA8dBdv6rokKHDiVq/g1L0mT2VrLRi2P39MQep
q5UYbCJoJ/+x1LPPn7Q65lXCg37buDBzdoFjeHEOvgdXNJrAGAcvLRd4TPpcsGF6
BiMVyjcMu5rqTJpWsslNLZjNkgJXi643iipBt5a/JVuGpsuFdwcqSg1U3gvfShtU
s2tjJhG1c7pH8MvfQxkKSkDWeBRHafYq+5ogABovm92VZb5eaSeMcRix1NGgVA5Z
Z3ZHZB0fqJRTJKKssIy7ckjjWnnOOzKqy+UqoJahrljvOygmKbg/V5vmKhAeLbxd
6EiOdIF1GBVLu5xWnHVs1xE87TPOaKdWVqL5eUoJzkTxrdQWdjWTHcqPcK5jR+ww
cxRbQpId6/fZ436Y6RnVZMzZug6NwoQpUmY+HhYtrougnJ4di5xHqUSSUE+qPp7H
33O22uawRODzUkUA9u3cD3e9PrCcC4LBdDyx/LQpYxGUq1xIw34WPdRNhAUXW0Dk
BRdBaRLoliX3mMhzLOwGeIyEUyc0/3CONsFO+UtKeDhQk2avomdry3lVb31yC9R8
9oEEh6U81QIhsd0EHaKO+7w7MDBoq+lSmYvf2EU6i3VZBR4z4QYdg9ie+w3ET2PA
CMYnQbvMN6Bvy5G7V6sXIhv9apfC4Aiozmx2tydR6Gu2dv0+B0g/yW3LNrtYo3jJ
pzlgr1BkDam+85ODgrsrHlK6+3Ato9mhiOIKFMBQtSECYebGP1PI9qEK5b5S9i10
3MYC3qhi8Bkvuj/ICqp7NdERJioUUwVbVVLXBh1KviJPeSyDfyW6lzLdObq5aot3
szJKygGFLbg70gTGEE+JuvVjs/XmDGn13BhaJzUCWPAsv50FWkqVlN8+4rU2h89F
JbpXdy0Z1O+Fd+ESnYE4sFIQn4cfNvybib7aTbeigKx3Q4Kf6bZOszFpVQXH26FR
prG1CD2mOglsNsDcDObdlqiagAEjbauRoO9BF36IR1gGTQER4VXweIPVvitZZPTA
iHzVL2bS+lgV+JE4k/uUjem/S13urc4WH98uYfMMAoZr4W1KoICfUB/WptQNt+vg
ovdtFtcn111atGfHiT+RqknLvFOT2ZwAv/d7Kz9dJU1xZcP8n6LV5k8ftkoXvXUu
L3dEKBGjksIQNhqqOHT5PzdVs8E/rwLd4y+CRGwv5hX3GLe/jiGEyB/BFcpm7mgZ
P7IsJ46sOnYLEwVKNvV8fwDqhgvnjGlWmAeKsBNbGbjF54XcSkP/W4A0BFNwJoze
YuvuB0UXUycAVpweg2sPQeH2hyFSfPzvpS7Bkq5GFHlMlD3My0tpqY4Qo1u8xisn
AUdSvwXlpuPeJZ/w5ySC8jjvwebctVqYAthd5WRGXuRQy7iNi3qKoYW6qOzzSspZ
VC1wsZHnXEC4qk73bP218LQm9lEsI9qMc0kidYV33qBQx0n7zN/d/uuOMmFnSflu
EFZFR7ib6oXl5Xs7v5iY+PgomVa+h8Q5Yne9fFLZ8FFHVwAYfoY7c+WF6tTBoJOI
VWlLrmiW5dLSnE0ATOyvN5omWZuWGJDH0oSxtnFOiQty8zS6my4CFkGLJO051T1+
GXiSs3FmxM+XyG64Ku99tNUhnBLMjDHnASO8ot9yKeGdcSCV0Rc/B2996du22y7g
BK4p2G1MccSjcBig2nMuPxZsQ89IZBWU6xmzua8OKen1rNAZRdrqMPofioetBvC5
y/l+v6dzKwrC7yEJXWj2Q3Preug01U4zmYZaUCUzSeN3P3aFUM9QBvtLh2+/el0D
9rKP4WTIlkjQOgcxL/T+x22WNFcfuodearml0N1A89FCYAJDpW0kdyHN/eCAkSP8
MABc3k4XPEygi3HSq3KiT2aAgvOvI29LZiyffFBZukFzXLWhv7UR62HI8bt09R06
Jv9mzh+AhpbbnHSuaBwwIPKAVAC1fE9OcCesDw53KJ41Tx1hHISifP4FgbD8WzDA
natzFoOlGENJYJGs44Il+yU+/ajOXrKdziUnLLFzYcCYTpJaRVh4CXoEAbfpLdNQ
h/xq9RBDsCvP0raCSZKTrKhV2fBgkpamSn1zS5PiA4iu4qZDkf/OFuCJ416q558V
mdjCOFEO/yOCCBQFJIVjQfcaPSNuM9wDjBrI7hLBwVwjEmvlshtfavhkYxWKEPfC
cNjbKGdaID8N9URauY/+2axPVQTu385cDS8wva9OhS3obxgkzXYRYor3vTNvLVzd
TGw3+CJ4H8hwXTTDGxFZ9tRaUfUJaPQ5Ag+V1QQaoNM0NTWmNUK/2AJTBxaYxyEh
tBoF9cAHrxb6pn1QYg0hL2hEx6oSRso7D9D7Y7KE3W9xw08DcfeQ25mAIVjxrqu2
MYc6Bvmspc3WNO9r+0GYCCLiPz8WwkmGuBAJkBedaeTZi/m9JfeY+PcPHdNdt96Z
QmlNn5JCCDbwSYgLqjSd+qHgFOXEnwOcuFiSt20MvIezd7cF6kRhWB8Ze7ZShhYp
O16vHWO6Na8ljGtYD8l6dgcI+km/xi2lPHY+GP9n8rWkqg1CsGAV6PhinJYhl+4G
Xl4VW0vbUaRSEgwgcUyNuPcELITDrC8nqRpDEu0vqwt0hizKYWtQvhSxYnD5ymUo
eI0hNIQXhCL/go8cSDTZfwUnwWzIFNw9GLgYVGqe4EQgFY650bYlnVWfBxgnCTH4
lv09xzCXjYxfuTgNtrSuLZXhmLPwt7ImAaTzu4+PZvUcTwhtknt8kWl6/4/WxpyY
4uLlLvaVaeaVRH6Ye9iGiV4emE1juRdvK/ziP5iBrfiJe12tKfXFoS1TRbl2NtBs
aOPERqO+DnUkaDOuPDqI9+8Qg0j4Zuq5Aw+RghFwRUca9wJ0pCWfybvuo2SGSs+w
vFwTIcxs6EBVrbXk/X9Y+4y027n/5o3gV4Rya/NXWslr2xNyAa1SmMmd+0cqwR0a
tr+ppzT8y3dKmH3h4wkS+SpLimKEl/CmCLaaVKEcmZResKzHXDPDQcpvAToIWcka
NvRqzDhMpW3Srft5nXIDQBoOpL0X0XB6AuKAMdwDotFyK3aINbOUBdxEsdhGNdfI
k2ITUZeY2GqP1FYfVA+pvfRoX0nYFv7VyPGalviHHevz/6AhVaz1G+rut4Psf3xe
8Ak/XyMDT3di12lq3G4ZnyPFzw55CEu3IMEiBBgxTqiRFPwwMCEmy9h6qxrjpccF
F8RfYoIZvdM2/1BJTLKYoIQ7a+rGJbHeUsTM2v5ltx9Dt/bCmv8d2dvoLJrpPQiP
fS99JpKF8B+4aD9WXRQO9S9RTLk07T3a6XScf9ATJXdHFkbEKY2APoVFJyhWmWJH
9VThNItE+CDaxSN5dD0D+5l4DjVGrwOjYPY/Xufpdu8bgj0n3P3ssccgIQ5OMGJG
DYnZc6OBXIYrrNz4bRFfFlU8rbLddSlkVZ0OGGwCIXkbs/5dy+7FJW/WwuOhGSFe
ml+D88YLvGbSdVvFXgoB6zg0lf6AcUgq5xcX/NbW4DEH61VxDyuWG3Erx0/cjFTH
mqKUio4gusAEAkQMFl4i8c8GzJDJqgm0imk1++0pNYy7zcVq2e3sHQ33pgr3orZa
2aR4uHy7nRK5I2BovCFs7oPHjYK/YTJAW2dIWh0aFnADaWd/Wea839vF/SBO4Syf
QAXtrRxYDsStohvo+ryUyeDSOYBuv1moKyZUBf7jiWA8jBig8oDebOlenqlSMux0
0BTrRAjIC3bDEwzmeg0jxV9P/2xNKE//sekiuEircGPvDbaIj9mtymxUV9lBp4JV
ft6WA0hQC6WSd0xR73oTFdYpJoB90QIzBKN/yLkMGCSAn/6HF0bU+uk9/QNiTHvO
RxlbD82bCjJGtCmNoIZcYtoMaRLIuO74QiRXKxQu20HzUo7HF/dXpGodtTFOpz5o
8Z9Ifd65JdFI6+U2gnJiJdYUPLfF2Rzz1nsUgdHw6tfentKu6TToySF93TAMptPp
xmR3TQdynVbwqu6V4EuRhzw8hGi/ZBqTMg3l4x9f2Bd28lu1lg1A45JE83bl++4u
SM5YXhmtif5xvx38bHuamfyqoy5YBV27Rp/eipF2cbuC9Pv4O+g/SCaP8nKsaKpA
DbdjrmkCtiFDlOJV0NbvBiyGh2lOqhFkijCPfUsVp5PuLxHCPR0tD5UkyK9+mtJY
UfQ0MY+PlDeWrUC3MHtux6pbDT9LqCn84UPwug+4olX9LIpdbypjGMUjcROH3q1U
7ptwSNsdMHxZFaFxEI+EpnvWkwu8HHboefLRBLOe+O9M5ndc2XaIqDtLDXuJ+Cwe
cKx3godz2kJJV4H4BHC6Jzw4a7ClZtXd0qIUuuN90WBB6PhuC52ymg4Z4D5cYYQ0
kiozGoj0BMZqUfR1j0Mr8I+X+J/V9daR/venoUh3PSaTQuzyuc89QnavwBR9cO66
puM00P2WUAT8WLwtNZMetQev3K+mf7uTayrLhuoCoilSi48dD2HQ81Z7GBBeai6I
DzI5hu/ja9Wuyi90WD1pJhUsJebsVmZiKOHVJz42PBvyI0BNlagfgyYk4ouOyE14
VgLyNkMlqywfmMWrgL6oYmud5OOoZW+cu9Xnj2igg9BmGFlm3ynxrEWSPiX8Ityw
8u2gDT8uFEn3HoEeQChu3r/LvwaC6Ibz4Vv12NQSlHKpoMa+OzpPSLkxgUr4CvKo
jKzCn4ZDB16GsOqw+CFJmshnX3p1i2SgUwakU5AfCBHCBPVHGkz/FRRP4p8F3Nvy
ApfxBH6o5rtbfD8yuhXeYJ/vS4UQ1rQA74tj3/atrKlpd/t/BhsZytgPe+2FfRr0
9cQGHz1zQOP5be70uGdkRnVgG56lY8vueXrXLJC0QoZ+yiisGh/R6xAJQOFyQgs+
sMKBBiOWfuLVTd/czXsSoSjSDkJcefZXf02MBwwxjRXlDoGi07MDfE9qwsGG6u5n
knIPZNIPUD67RM7t+4uz8KqukF77ARthbsYgsii4lWfqf16xtGwgAM+BovvCnkoR
hdaJMv5GE9KVy58joXjwwCXhrLpLlaWSiwPR67J+zHDMc9ikcaQPcer5VroRhwz3
IyJWwuo2f4+KljYO+TwqdxjsMMVnv4dZwyJ+RfuLOsrF9cBCuPUCDwZMktG6nDcu
mlVS7lQQeAGCoSlXte1EWblsHbqeV3Fo/fOOOgEw07cIKC+6BGLDBWC7gT8cUfe/
APJmIjbZdZnQZNF3rEh0VQSWEUMWpyGbylQ/W4Fbp3xV9r2Q5qEKGbwSEK6eylpZ
INTeQZqIsaJpsGDVVCw5v2xCYz2LvHfpcbK7YK6NRw0j0mEsdQmxxiJrsQeg33wO
bVanZd2SN2dq3MoPblyY9f6w96p5jpmErIyD+qj58AgnGyWB5oRsqaTquApVQvX6
WkGjq5vji8kebohQfEEJuJLRxtyQ4Bltt6FVD8FYtrcv9KnfcLRxO2dpECQBaRRu
QHV8XqwgSTYFq2uye1Ww4a4nXFVQPgWC/y0E8P2x0dk2QmzfGIA68puCe4jh4A04
VPkO8frXTghQKy0WhO1HEN6YqdEdqFBVmdmERDGbW3mLfiMuWIbVV5NhntkKGL90
QgvKtMDG3ycXzEP8ow4JtFumKBBI1SkzlCCRCNnKD6QVfTV/n6+H3B8Ic8lQF3yO
xnkYGvPuoXfCWOaaT99iCta/PR5NrfuUnO/mYoAjZf7xNfwjeRoyisLoNipm373Q
Uhq8yB3iM6J/mo0MxQnsRx5BXGZ6eFBparY7csBhcc51oxX9VBl3W1cH2A2455St
H8DKsm79khRiblQZHqEvXbGnf8/6LwSQtjtcBEjdT5z8pLzs42usrrdSOipLzLgL
g1UmqfHaIuIOhefLG39vgUyzl+qWe3Yp8Z/cy/VwP7CX+sTWaIT1y52kXAN3cEJU
wvkbevjV1ekLLOtLqBk5SntjYA6wo+wr6SQQhLfZNed5MrbxwN76D2+8kyx2XmqU
2ja/u8z5VSeEtApMxwtzHwK4C1dGDRgxbXQtlkv4YqY0VIXCU4SeK5Q4n4y9QSqb
objdkdQN7ouqSzPztvqJTVHWrwnI3cbf/U7PrMT5t6gFurzbSbJMIUs5MirXZPrc
cnWN8xgBaefCLtvefJmQY3CQlk9QPWqSX/nSzk0XkXyLKedyte64bHSFP9SjRVTL
/G2tmgP9ftHvQ08y5igJI+fHQ+SqVbJ9vglXiI27gwHtptjYLrnFuopXeTP6eeh1
XzrFRVzeMRvdkOjrEmAJPGG2SyRw0rfg0u9wiIlxi+BfwJSqGyDtaIlDvd14jLfh
Zv+0RIhwXjNDV7hauFcqoXndniz3OkPJ7EpQ1mYgV9/Zjyj8N2t+8t4zmHWm1xD/
lXKrYlblg716KGZpjQbTeevzygpepaCa07R3DZqPVygxOtfoUKDWOj4fvTa3j0I9
B6By5aM6+1F3+BH8erg1aYuZFmVodVbV1iUlVqHWj/SzTNlABHAuxE8BPhMGSEuW
TRy4gfQwLddKoJseGB5y7WKwdcoVYfSEHkF3l8nbpKTL67MbSH312ZiOLWZ7iB5G
CItAv+B6RGQH2ll+TVqPXpEDLm1CuI6xxWb4vEdTnFhBOEcarym+hwNGfe/YMnnj
99eOhZX3LiOveYhZ6K2SmRbNh2+Btnh1RUhKtKd2G3o/gg+f0ABwUIkYcxIDQ5cj
bSo7GKCrEtHPu4sY4woXFTtRkAVqEkbQ7MPMt3kjWuWJBEGFXvowrkOCEm7gGiZO
oq0WElHftefAgqd7kGZCDCYWwMCWjrAIxFoo7XeFhLhz0Tp41JKNgKIDk/FOE5ow
vuFiBOB0UbpvPXgyLIUDGhMmktpDjWspqW48o5CGurq2g8Wheo3oypifUo5oWUAl
V7KREbCBf7S1LTKzam1kbVjFeHIZ+3E4z1Po04/lq4kory9dXafkgyDIMSXwawWG
J8olVwRVk1wqK9Hsait9vjaVrNKUmWUl5barzUqO/aIL2krzdvqYMqCQHlkToF1B
USDkCgRKAxvCJYqfbOK4wnnULdlnUHpr/ZeI139yS4RAXels9lYMiy2bgd4iX/N0
aa7xKKVD9/e88+eYbRlUBXmnk5CARYFh2AY7JdYfARkBb0+AqE68AQ4YEL54rqbE
0AtUOMq2pf722cQrws3H0O/GA/kbYrJNZJXnw2MYWGbIPwK2UD19xMHCV2T/3E1g
BlbwjBur2W96/mgXjYuW8py+P2zoVvnXmjhIWm1mZvMmJ/4EBEPQy6Dtq3PVkw9f
ta/9f3guo77vGqAtjPwEta/f+paRarnwpvNEHnwi41YtI7xcGQK1Mf1eCtkE8EnB
VEt4xmjN3DabKw/acB5nW1TwI9zS0Cq/CDgteN66Skx1QXLdNfHYFxz2bNn4o5hN
PkvOmXz2t8353KgBT392ZZ6kfQzeW78tR2pWWStWC4WqY/v8OzD4+FwLtjze2Jey
U6cx7Oto/CPArOD8tUmrnGxewXzU9RNQSZHtIJlS/OkizTGwv6QyZJfHf3tNLXRi
e7eEdJt39oGQUxYXyTI3ndvBfj/uGrcyglukmbcSZDsx7R1Qeon4AhrUrZUgWwcp
lrMw7d49zoWPWaQ9HrW01SwuK7NC7fKVJli18gennRaQZK/JRVnIne+Tn6Ntjw/s
WMISLJWABqmKd0/I3CpeqlO2hQHN5MogtM8ZxB93bcAUjq+2g7ke0HjaNLnPnpW1
GH6CnVcRSLMyznhBgkdSBdCqfPmzVhGFcW4ta310cQzP1aFtsYpisbh2VdW4YPt5
KGUXN9uNh3wwjBKT1M3HqWOlEv+ICQSZKwdG1sdb5ecS+WAGGZfrAIZJzCDd8vIL
eiAXhRxP58LAMQsD9vD31NEeMAfUo+3kMEsgezXJ4jSAhvvjSzLLA7VpS1beg74z
Jzsx810p0PTOP1rmy0zWS3G/PRBFU3UQhjqkDkWQj340Gp1OqIR2CSM/3craU8lI
eBAJGiMYESeFXjI9+pXZaMFhh2Cs58+sQqCsTgs342pAqYaxC/XTq7f8x8AGfol9
Z5Z9tHZsN2d/+X78iYUV6Qzg6QSoY2VZr6I3NghDRCaXFo/p4vvWbvHltwXG2nE8
CNRqQquNE5hi+btOp8Wh+50K5MIwj7hXIZ/9+JwJUjgB4F5WR4BwC0YBEzJVkdvF
/Drtpcd9vXxsqlVD6jkWrl4walDVlTOI5SG8S++hzdbSZolfmNZ0ONph1VNJsh0M
n77mFq4oLGZ4Q+5v4qtqRiFi+XwUhU6Kl1tMCR/D5yqB5Z0Bwxnf/z0rNOa9+QsT
LWEzHxHLISfDSgxcE0QJDPHo4zHjqaPgqEEgXn7KINW715mKqZ1e1MOXMXtiuykj
08tYQMowtDF4zhzaEa44BaKXJn1GHbQ+QqQf8RgyaXxv1jImlOfZ66eUlpaO/wzA
o5GY0bXZpdMl5+ceGbTUkBDxtUetT7pJHBdxp/e0y4pbDE/hHr5cuAEvR+aNeLpA
C4J3IT9+HiJnf7m+FLBbnBELxWhtzduL0je/JidMNCN0+Eu+XBhN/GnpuOI7+PmZ
iULmiUu2PXr985O51o4SB/KJ9+c1pEKD4hVIZ4d9jyWbhVTuaOsY20XwP8juHPeP
0B+KsWP9GPUo4R1N0wCaghxBnrOSLH070RA7EI/ofY2cZt4UrvI4FfpmHeMv7u49
a/3f3XfZRQIO4kb3QP/VefTh+qQz3A6PKuiVhkPMQWp0ty/UjWEBhSxf7Ey9Ym83
oJ0Wkkh/ikzqkQdfATYUcP+QCT6vUJWVJjqyVAsc/g36tGdMmcCsjYQsVpcWHqz5
3cltR1gdvHhFoTf4C0hGatU0vcVBnvqMucynukN2Y61uds/1vmSyNijKvdCNSpsk
Szzzxn0Npw9k6sLgYu+ya9jsTsF2p9U17YGgKLFT2cBIx5t7qJdx87atQoCzk4li
k4tSHnKYcziBgOxJYOtv3Z8vp6wAK2NvrmWl6nz4NCDVHRVUNua8pNc6EftYZfrE
T/8u5+0ZV7EugYAr1NDTl8zAVkI2ykiAdLD9oG9fl0CAD7lQMVsm3jm5EOFdiFLs
hT4CTzEZ6mbVjRSwBsbJJ5YAkhlJdg2KPvg9V/StHUT/ePjs6GQQe/lzYpAKlbwc
jxKLjviwYxddYl0Pjxc8HL4wa+etyVHYuues7C2+pRpPcuyg04ON99m8qEkU40ka
QPygtBxQm5Iou/0CAUPkvdbb5re5sJXyyi2OiQKc4SFrA4zq/On7i95HANro+95v
uvnubDtBfc4jTULkeNyy+7QMdECrS7M/vw7JApGjVgjkD/VZS5SU901ysTxnpMm5
rHp2/Q9U+DPceNOiSsUANGqiJvhrEi3mBRI/rHf6/n6aq9/+rwUWs7hDOHQwk2Xg
wTYzGqwaDo3DNyZR9mln0IU5/p8NHRgsIm/1PZe9WS/Lg+85ZLcpXjiuy/Sz6ogd
6hADa1CU9CF/c+gWQfXLJ89Nnr/cLBXDuVz7AOKfwcST7i7fYYWUCFcaDMEiAfc/
vnqX8jA3nnXx2yeVdzSC+8aF9Jq8dbzWrodNgMvcOkiMaTgMjWdfTGuRXF7Zynr8
Y7xhMODfN7ZKZKHfWCIxfvUUq1yqp0gIg67lxbfLQVL+HJa6QvLdFJ3+Wxa01FGV
CRxLsK4DfnNADoCwsJMrFATtniun1p2QAy8gb1fybx0WX80LzwQVQTlzN1yPdytm
jXAuPH3RhTukR7Jj5QsHkX11XTPTfrdNcNwA+nS0o0RrKnajBd+NXeVsfrDlbEBM
y7TAdIU22pMlyoxHXLo6jlJGSwSjehQ/eT7HuN9OFYLUJ4IQHLz6Juq3y60FxsDb
Ru47ImjzrIj0pj9achMdbiNvUv1I0DGm4TsaElya0tsEZEdcd8wY1nQTjTibWE4d
ZJEviYXwsq7g3LRjklu3smIOurtGrzmSxzjZA2kWbgr6qwlB5kcpz9mBdey5QDAd
v/hBiE5znaVe+ucSn3KXv1n0FGOlBD5HasBHCRIMaD44++jcsvWswRrjoox9mqRh
SC6143SNuIvxbCLZ+aUV/4uqRSMf+Wr5BTqZnvBt1S3e1P9VJOENJBUtZo7ySjmK
McnFTYOBdH6TwUdvRWmqnTiPOBPIJaFAHUxjIOERqaG7nCdVROQKV2V8Re/iCGKt
4dXX7d7Zg1SNcO/L4PdxbHU45sVSyMgsDLMH7L2U6iHaR/D+1RzcgCFxmPX1XLcq
XgSJcUYGQi1scEJJJf7fTRzNWo/JCLiZya2/qzfkpDY1R5fLdPBuvXVrFdSXA4OV
qsqt6+0RmzpyvGPw7DEsSLW+p9LsZIFIYjL5Hi2UajYNutWt8iSOHCNcZpqDtoy2
XOfO5MY9nKkjitLgT7WUd+FVpqW/NulDnxkeSCiQCjcJ3eOQP62m9NmHXfziwCvp
o3ljHmYIimV2IRn91ep47FYdE531g2YsafkhWxd63ww7BkfLNoCkW4uQ499NVQpb
D2SJkAQfxQ4eatHVgcmCt6spRJKQ8ekdCDR0DHbIWGRYXgVLe2F66AdX51YDuVik
qLp7Hp62p3vVO2xRidmhi3YopfDGC5n+U9rtZsEWLtIWfP+56IiJ60u8K3XLN7D5
ty4mp2SKWUWkLgdKpiuHYHT8BXQ5lV+d065yRgXaYCCzNb0eIjWLJlv1vmG2q3cH
0j6J9ACr/fOHYoaoJG1wF8OcJ25+YIEnzmvzGm6HN9aU6qoiN4antwMrzCEZxLig
FKG93GgJG3T3YHf+0zzYlHT6l+Vnt3/YcQLqkFTdQ/oFO3eavKtruVTRwTO5eHhr
I7Wl8WxqQqBp5RcnFxZR2mKO77AWrW5LSgtHetQNszu5V2VPFc1XTQU1uf54dVAs
FEtTigCVoOotRieoUtAGLTIXMJ/z4DRLemvg/rXM/fLveB09a6udT4g+YjINyz1M
xXLpEJJ/AHQd1eGM/sS4LTMC4Y8/zl/TE1US7oa3uniT+SM3jPvHjC5z4l0h/Yts
ZXjVCssb58LRXZ47Tdr04qjNMGXn8xYDCcvnHkBHqECP/okj241zooRtGD+A9aAG
oRjIC3uB5jD3xDqeIqYEM89QO5MH1FupczcLnbikKuyagwYqjib8NvJLsvLy75A6
4MYx80FYR0nbBbBvHdlcvszHrMLLYuv9nKD9PWJhOjfvr674AnU9zQvTmlC7v8kP
c8ebKLZrBymEeJE4p17HWJouUHrEvB+BuUjqTqMcJF6jJ66SxERJ/TOC3787040J
eMQweKNskJKY93hw/hnmPFrxQNlp5PqSZv67ynxHXbcp7Daqj36dmFhKxfjUi1Ld
YFKBde3hgQu9hIYLqs5fxT5hGgE7p8rxejcGVeNpgDPeVoiFpACCDevNwr8qZJ7w
PfET1iD2lclueNhgRsuTZNQE/+Z698rorO4sws5cGs2GhXdZ7DiiT7ErSLGIIMGV
sl34ASn2wyX3Tuyyvcl906GgsHWerkWkitej2Cf0zayj+egsWwODJfiyw8XzcNsz
7RzNoqNZK5GSjU9tWiHGbib9Bqo7PoM8K/Voy8OeEAbC8eU1Rp26SuEisbm/FieM
ubSFas5ZKMp0sTtU2g+XCt7F8uG8WDl1LMpnYA3C7jvLgMsKFdAWWbdeToo7eF2N
GhVk/GSJEqXDOrkC6k8yAIk0iZKtsoSAH07OX9MvN3sEiDV7q6flRT9xWZTscN2F
AmVvRn3X6fwJA3COnu2g0dabau/8L46j2L3X7RF4TEOd3nEmeqtUbBJRx8AzcWn7
yp/OYjOg4jtTXoSJolUG7bE0h30NEmi2HEcFpQseEL5dCeUzdNgwPzGqRPejPoni
UR1cwOs4l9WR7v5bbyXZBSIBgmsBUUIKQFiJqsq9SojeRdWKm7BN8kwj8+LMl9w1
Uw5FXkbs9uCdHvU2fYeD3xHKVGaZBn6Yyus4/K07F1fUo47fAeuugwaRTxqiUfnC
+U6LxbpyFM0Aw1xdsiDRTlmiAmIZAx+clmvddL/6pf7nQd7y+1Q1daDWd5FoWGVy
65aLKvMRjor3u69kMlEbltIe8aHtKzxwAj4PXwn565LSr8LomNF4Pc/n468RZTnb
BknfPw/RUS+PDGbEQ0zE7dLDsKeljNN0jHvjJXr7pgOfOlGd2pNnL5Wt7qzzmyap
DRczA5H/F2qFfoRHj64ctrYtoxRM6Pkr1TiHNhu7HkL/2UpUh/DzWV2twDKyOUL3
s+1813Zmo4FPV2Yr30tMn7LVOV3XqDJNw9kkVz/rmsWM5aN6zeJqKwNYezvyO7BF
WSpCjN9kotUEiObYs2lZ0jhiM0h2UFw+seJYiIH5H/a9FAWEDHf3Yv9FRuMSXwJT
FXN6cgeLSIBx8w+GX3m5Gel03njg8Yr0bswtPVmmO5rjvYSl+A9KRnNtOrKfaEsl
GLPnkM/rjyKgvbEmzyfLAWFgzSXVzahv2wCCKL26zLKvdsEyBiW2bY2NJ2v33S1i
o12oOhPpTN8bDZpE3PF3KoQZwtTxkAZ/FpeKmWyGUPxNBEWCZWuZmdbadb8T/4Gm
bZ+EWd4NAL7FrNpi8XIf/uQaRI7O/XNS+4yC7VzHpdYgHqlwWMBvlMXuWl9pNEKq
ezElpMzQNIzTNHzmStuJf+pRTVvKYSYEN7QH236+V9j6YWf7r0nfKPq8XcZoPmJe
X2UmVi54AbErG4kd1Qz4/KqYJrmYIACjqioZAMn2TKttAJwq35KJtC+ZmCl3Eq2z
PuUSDLL0b3IRvjJx1YEKPsU94FAjA3SfdiLjMKWbpGifdQtKa++rVLX958q5MLA5
PiGr6X1EgbDvs2Mtsmzx7eFDSaTm423He+g2g+5K3szePStu74d2QZOyQ3PH6do1
WYhR41YeBGVWRAQDt82hxNUh+zCvdYjsGPU9riYCcKWsE9O5I+Wts6GoLQJlR28x
+ibHBHSt+WrcVu1itcEWCABAnqj3GUVc2od3vh0uzmRIi03Bc4HWwqS+VbE2aSE/
h+JqlOQr4eshQ5zfZ9zcxQuWjeSjv1m+XqyLr+v4XSJExWUjNpBQ/JiZxLNMMHXR
M+RksTLhGEnm7JHDtYRR75Uvsaq9TlTyqluXCCnsqOJkjjQNp7TV9CkDcvTohvTf
+tSY22y6Uq8QspVQojjFq2l/EtgrqbpnzvMxPRgNYvbO0mSSnjUfYEkqhTgW7etf
DmYVLMwnDvSwTp4JynKY/bmyLbh/pZQbefRk7IPZyakyHvGcS2GlfBmIIPJpLV2U
yZU8O3PaUOUaZtPD36dqQTHvgEnjXxVI/7mafkLPAWmnnWXa0ffRTR33wewZ+2G6
iS1t5T/0Z7rHKJz6nLUmehWNhsMjWu1MD48fYeRLGNmYcXDW8ZLgsiWX0CR5cTrD
FxLXmlcVcxxEmCUsYr3Jrtms5TmZAKxGPSmeCcER/a+7zMOODhVbLLloJJDZegIR
0KejWnobxqvDlQTZK+FnlMM9L180wqHIFxNMvf8JmBNz0shn0t4i5NVBI2u6vPxF
cNXrXiwiMsaOOOVaAsSDn+YpofZT8WiFORgap7A79nSsUvhFvC74Yxn2hzlvS18j
X9yNHHxvwbuL91kDBqliny+J0mg4YM13gKj6km6NP4Y8FhF9y6/hS9jNcKYtaUWZ
hKNQ28b7woRSlKmDRlD/Ss16zdxdYfAxdcPR22bSx4EjY/TMM6U35rNPJQma6xr3
WSezcc2UegazJFlJ0qTqo316wRj5xuHfcuuUKvbSV7whvHUynurpk6OlLr/oByq1
2LIHasre553EdJZUJpj5WiestxcwHKZoB1pDoefLTPvPorU8f4qiqkioxmQqkoWl
22RGBqsBOQajFmkpzPJZm/PVgf6jn22M97lrrHtaefFFd4WVaWm99zesXHOU0WXP
KiXgYfG9Dc4yegpJpJaJ9hmrUBsA6vIK7aCSJFvlp9Tc2tvwNxLMF6uWJqZwi+j5
rjZVCbCua+MX8il8gnaiGSaCbzDrXt+zI6rBIGfW7EboSqhpc9fEGorWHeXmQNlT
Ltw/kjbwnU4/shNwjYpnoENgGlf5a9Ec7gEQohlHYX0g0tOKvhh8um63cj+ChM3q
IgbzTORWfEeyaBlx6JmeiKlhQkM+waMcSAMt1t3QuIZmWFCVGaLNBvw00sWPZcBO
1bovO3CpeEurh7F8Krkoubyi6V0tUBs2/wv56FqI7k5fhGad4dAQ8MN31wQMV2Wj
E239nY+G7wo6q3sJZE5qRlL80L/35ZQka746Caa2Vm2tGtApuyK60qgqAbv65Vc3
eWIV+sMLZS7e4D4qoUz2lMRN3dWaQE8FVL2Db+PV2VdX5/Gsudj53BjcSAcg9GB6
46RgujKVi4L4BRBWoY6f0TpMjZQrEFMGtyprz77MP2IOuJOBISa2eWMdxRNTcLM2
BCQxiGondIaH0k+UB2H4Cw41nr6LQtWE01WhgBBF8NgSnQrkNMGPAPRuWZkCE24h
KuyKnwM8zFppveGYokhuc5VKwtRS7e4eFTZVCKm3EJhPnDPSqird5HUkDylP7F7q
2iiwS7X99TMw2QDkcdcQIlhDXFbeH9g7bY+K+dsjjiYLkkrvtLc0efwXYJFXWII6
mLvmoiGfiuABh8FJS+nq9aS6xn1DFP5fHehP+J/W2moJyofwZHlkeNtHC7LsI4aU
vZiBViHZLm/VLoamUixF7xT2vWyBTtmoQJi5aRMIOwvl5ehQevs50QeCHY/zHcoy
l7DVzTHBwkJqWtDFqUqnxvDiSzcCJy00h79MyoobuaoPqxriBxIpZtOu3mVfYXB9
MI1zSdw6JEQZz15+c4gsZyhK/tYTIwdmoKNn+vsza+KkvXQ9gOfCUoDXCCO0wvXn
fLj+87lXeOWO+CchUDmPIfHPIPLrtvU7fCA2jRuw33KjcOwW3lc0fsj1QNDbMQoU
sn4dQjdCzeJuR1Exul13ZtCd6igQgbDlnmNPQZjo2juwT50dG9/VKT7+dv53YvQ5
Dkno7sne1VdrSmC5gijHbjlaIRgN8asjOVaBk0o+NhI1Jf5iFoH3ca1YVzcoJhP/
9UF24lDRlt0qGwp1hzS0zyAKtJMqD5Iu60SdJwXzveGeAI3ibrbkCk+5aP2rzsmn
Byw4dqG33qYyaQ7yD4bo8tRwCfriysxaReRytzLFhLrja+C8yNup1wkoE9aQumNW
Ne8nKRZ1fMT/PYlrxoiSnSy9WcQCabC1+COzZCdRfhGUyipGjUOFuYXb6fdXq/iW
RGyn4Uum46MmPY8JHORing9YL0PMyUQUxZ57S9yFrgAhcv6+HNGLeolGixqGvGiY
CydszCvfs//iwlnvFo9pZ6/kwquK5/KjERp7fUgRQTaslAhfsic26fNwGN316YbG
YYq9DZtL2rCdA8zejHY4ioehI+X1ZzpRqT9ikwuoJgYHhHs+mpNEFmosdjGfVlPD
2WtoOljJ1OpllebMyvwtAE2qarp6tQ9KffTeRA8wzh8f992J2JxCLVM/0aT/nAIj
7S/t4cfAhruBjOSddalITg9sZhKB2RTbs8KTTahSEYFMJmxMrWCdq7ejyGKJyRMr
mYPkFj3SMsWQMH2fC0gkMA4V4LatVuUAP3BnTmsuLIFX8tFwTPFTpYsIzu8qRqQs
0c3zfxwoSHJ7tfFvse6i/PQB/b4r4pc74uAHSoiWj10aKfPtoOurv7ay07u0QEa+
47x32FG9EiyxddC7OhezF/HKlUftjTxCK7GBWgYauKd+OaUXLW8oiGvsJRsViSa1
cFg6zNH8W5WYPJgAb3sncZ/EJZoNOhbyB4KGyVnXCIRa2nk3cdFyksjpvG5uNRXK
Cnq9nY7XSlVITkrhXrNBpfLYTaA78c1Mk6NW0V67HxH+7cg4oTl6CyX2+aY8UNPr
EfGnnP6b+gDgfe6z6L4fd1iVqTv5vEJJ8sMjPnxC2v+nud0yFexcDTXjUHPforJf
oxT/KTlaFLVjugR500nRv8N/5fEiOjv+WK1JdAczpj8vrEqtcYvQny6OgpXIUQ+L
mO4PdrQsWTB9hw64vKShxOFicLqkZ9bykRpzsRP8jPRZ+ZxXeLC+JABW4hhXhadd
15XSV9b2oaMtLET/Td3dLf1HrxRjJsWfjzeePFOBhCIkVGl+4a2ndEJq2RlAw27k
6dj5VUiVW6aaYW7r+3dlF8x7vlN56CsTE35znuLfeg2N1cAD8D/dm+tNSeJmvSVs
DXzY5F8p3AuDyI57nWONIheDsNyQSWy3s8TvLSAKeeoIsprE1EoOeaT5fvmeVw9C
vxryvRLdHdD9VtRnl6YEs7/g2VP4vSZPdS1yJNGsbNVr4vyWe4lzPXTDb/A11xSe
XMh5nJWdk3egbHw1oLwEgmere6ENXy9KAQFazhdA5g8sTs//jPx4ly+H2pLMlaSf
BX/PIk2Qc22hhE7pSPdnJfDYayQLuRmpTT3smONL4TJcukLwjVHsJFk089u/HXoE
1tcCEdI1vrrAOhlgjjT++d+akBLx9UoplyDNl83mnsSxBCr+CzrCTpKSe83IUpQu
rNDWx5TUoeJ26uSXL8ZGq07wRGvg5t/dfBrCwze3XBFYK8gUddzqOmz1uLA/S/Z6
QUhn603NQ6ZLVjtDGNojBQULMKAIj3FPmuo++h6wSyvH3tF4vRX8BE7thjt1ckU4
EG9N8mMeMAvaISMcymfEl3OMQxmZn9pjOLJ7q9NaHE4wMES/aC1ZBGpLw8EZu1E3
3CwJLxxU9J02fZBPpuxqj+qcwljF65qN0kuvqYmRugyJpdlecL4fmF6+Vp0jmDkK
Tn44Cu5rHP9o/X+weMjCOfoIFIpBnuGIFS1ekZ1yPPnNpOZKPDIZx6/7DKZiSYC0
IL2M9t1qwass3KWTfQIYZ7IjbZJ8vUooPmhGunH3Em/hCAcZslTP9PAZVxzvWauY
uoWlUkIv1Gus04Z6Qnvsfy6uXiFt42J94ZrCBPWbfPe3sfZLSs2Um3UD7e1YWBR4
9Zl6+VjzRMPVv0OmoNLxar7LUY0iql4EAj7Vox/B1qE3pOmSKTuchQL1mBrGIkWS
n0EAiaYZdJPUR4rjRLLwCAFFppHrHXF4rKa/BrPTRurGXYteDpXTROi66f98mqq5
OPvvvoFyjHkAFh/+SqPBvN3AXeOvqDBca5tWmlSXHS0DrjxX6BXCWy5KQmejif2g
N4dDcrGuvFILMv+WfveE2W5jOwFFrP/Cb/aSZVXOeFhA6P31NsY0CPck2UduTgyg
vOdUsz7/Do2wwSg+vvpRQf1cCy3iT/L1vhLYvUL/FnPju9hCdU5XDtz0VcPIfZ3e
no0PG4Iw/OX4fmmJ5IfvI0XhXk1RSdKsoWLKBwTfct5Zsi8EKBnviSZSWEkq879X
p7P0h4R/l5KmOuHdt/tDQYxnUVsrxJ6RCyy/+23d/rxncCS2HBekIQVO/mo6V3U/
VhYOwKJ5gvdbGJSQspTNlja6PtF5WgUiGHvVhiQF1OPE/dO/8Jr9oF0SwhI4whrM
1A50dv+xnOLKCdPKbjFiHqk1WAECfzWS2cydPm9lj7ZjJpCU/rY+5wStvGHQrwG0
JBRsyckg1yh3oh1jRbdSC3rlFrqlrI7+HrfI5OHEJsOS4Jl+Pm6A6jUdsNcxPV6f
Vr7tn0dIwm9SjmnH92sUvt1So1HUTAJboQXLQbTEmIHJ6NPsCJNm4jhJ7ijU9qVf
kmsn/+eft7NfIS8RdWrOk8iCjiC2Xs8d0k78NGwp9H2IaCzZgcmhiu/IZ8UYxIne
Qcymi2d4kI+SW99a25yaXx/Y++B3t7v77rtC3GgesAdmNTVvOfy27heHcXV8V8tD
pGWvSksY8q8YkI/Wwiv8xBEMn+1wlGPWwdjhrNbv8nkUC9qiDqBO6dcxb5/R8YqF
15dgIdrpLN9Y8Wf2AY2O04XIIXNGHAzGZ53J++/OS3eOqe9P5+RXy6KsJvbtZ3BP
qRGXCmOv83P0cwfrLuCFfAr1NDySxTPC3xMJ2W3hsZL+C6qb6NxR/Z14w66dEXfb
b7Y9tmY60OT/NsdOPFvdlISYJQkB5oLpbFbhC1seyTH+Iprfn8dLby80uNEy6AaD
QupMRkzC9G4WQ3lqxMvurdHdIQ5O4YSjy+kn9GXj00IJfwZX1izs9jz1BxIgaQbH
SyQo8rrfMun2a0w/nsWjTvZg6vPmNXnxAmRNd3gqAf1ojTJVTTS43sG/qWYxpeEE
KGveD6F6xZRnxoN7NrozsYY/ESP6fAW1UIViJ7lmExrv8ICCXKt6on5z6jDshiYr
BOu5EmebZ+c1qE/P7pN7IMKB8YfYDDxKcpL0TSvp6MMNBjFyglGO4iHJq+Y/3dof
ALHkqOVwFLxEsA6bA6zdKDQVf1mjheCoFEfy4hdjG2GweJbhBue0gSVPWzGOoST1
32kjbAOx4Y1o/TTmRtawBg94MtZr9T4A71dA8xRG8sZeyjXBl9TnXXGZswfnOQlR
Wtr/iOXzuSrf1K+yjr3NEo42Dk/H3q7QthGFx3sEKPD+csa30Phi7Hd/bbB7GJCY
50y8fKbllSNtdJIiiIQfqRhgzJXF+BXK+ysmI3pYfEeDvkohFxUKRBWfMPrVTfsR
IghPDZw1m71hK7EkX1tNlsoF3rm8lI9g6exdjGWjq0AxLGVo9dSa+JEJiyTZ523z
7jgsweQcbsL731SAFgpQax5xYcgvC4lD3p0zGvnSnG0YYUuIcCLjqXBfcIiCm9g4
fvvtbwUW7uu6inDHj/A4btnRuy/42ptjwkyVrGgKbjAARSldMVA1hHudqEfuo4H6
KZZLOWYs34xPAii2+DQWm+kp30BQ1v9aj5rTCsRhaoFBT2E70UegDDrCvEpZFunD
k2D1vmW6D9J/kDX0IjZK2WKuyoQcDpnpB3646agAxjs9IdxpeiWFDa15wQ8f4bBW
pjQIcedhWdmAqwgT+YVm24Q/Pz+ugklXCJZa7E8NbR1ehFkVwqOKXSLw551wH2Zm
fM/ooJGlrnBmQ8fOpoTm7iHg7VzzQgqek4jZgcQIEZ1T/bq5zjF8Q1UuOePnaCl/
CncD9Za132wrOnRBDNOKcbqz3+cRDza8QEyoN3Km2udixeyQtcFoNFgCtGsfarRT
nZ3kAm/hAm6ExIsJC4nbNOgktSxAoJzzStlqh8I6XC1+rZtZiyEmlpGh6cCtnzgw
LyIPMc0ihGEDO9mJkBAkXLzePBZRDVErH+HqHyOYvdayFiOZ+UZdcRUoWSx67ha6
yDZWC6OPjS5/RHfvN8ygxDKiw0DXZvf87C6yfB5/sH4DgBmSOrbiylou7TlO4io0
rVTz5Zscl2hUp7dWeVhfKBMKg99g1A+jiXAKG5zScUQWZJNL7Nj1rY3bsVO3OiDx
y80cOg2OP7YI6enXcjFIFP+FSYnewhn2qhQDn9POqpupu93wYGuxdjzqnfA34xqO
viTRMnJ9UGq9yrwqmuxeNBsGVYmS/YOxQytcAZ1JHubwmH2QHXO64YoIwVk4JcFC
b3gEzi8GOpR0daJ9jJs5SohoPlyxTPL9vMtfSVfITTIFq725yNaujiwXKQY0r5no
3svajjaFG4C8Vt5/GFn2jroh6HbF3jg7LpWJU7/RuDuaIBd1D0D+2j26TgqAo2u7
xpb+ccScEDWQmk7D0E5A2/zKz0F7z7FzovvQjxZZpkZW8h/KH4eMJ5+WF7He1r6U
EJoA8vDHlIYVXCBfPfFc4jFMqa3RgbtuqwJMHR9d+bjEMQfcnef+j9/Iuk+xmof5
mGlyQEdaez3jSpU58Jc1w9juNQtuZhomeUGO24kP+ad0HbbQmV7bJedR7Ku2eVAn
TjO2sIUJEAhJrp4qmG93LJJK09WqY0ZWIysufjLCwq6AeCsNZXdqSJTZvK/5I/7i
aaNcNeRkAUkuGraPxT9fNIoKDpuNwo2jm/8Suobv2lE7Ex7pog70+hy9A90uWSIU
vJXpyIcra5sN+rtjF/UPyPNFBiILjStHTltxgBprOiRaqvYfizINHdZ0vdgdw/Wl
6XiuJIR1stlimM5MzXowpZKgHzZsp+wy/H7BXgjYXlJaow0OglB6DQVSv7KPFM/A
U2Wz23cYT8jDZuIhg+ks9TRLIQ/8n0eZPMp/RC2DRiCQYzt8G6KJpMJmOJ0ERkYH
p51bfz7me96JSHjhvijXXTDleAGVX2loH1dPmRPz0IgETcenOA/r7ac4BPZG4Ir3
scKzegnQYDTgYYHjWjJ74n5aBUdL2+A8SyDeWXW2IQbD/XWkzeipuDn+Q01BGG+T
b8xGnAr1EdzUPJNe3lFLjCxrFLSWA0t2fPrzlTwQYrzPrCQj/w/mgMsrJPKEZIaH
vcNzYRAksEEtpr1VztUWAepW1bNsCJ48Eyib7TuDRVviLFVH4dZbNAfhvqgfn9oG
lEgmJXuQLGdsfjoLtFCJQFjWsX/ZfVXvouTrMT73q58VzPeekvAMD9PUb2BBIafP
SLu5cOrMOeMm7I2xwfpkkqXJQ/ih4sWQZbofFrFl6pBOO3kJS8uC7hD4fZl7qNPf
1hAwWGD+ZK5QlVzlRSVZQiJSmEemlAZsx3U9SZdY5ftA3g5fGWJT3Fv4KFiLaXjp
EcAZjZFTYeeJexB7xwVvLgDafTNUkuJ6xn7xyvzw3p7q+rEvS1qbF38JiGBNeQI7
VWyQhnul36Z8Re9nTmEbEahcFBZVuVemMG0o4qoL22NMA+StBVLAlbi1K+Sk6On9
gco0dyb2k/ZF548afwrldnzeWt5XRqzcPnguUdLNunJjV29Rds+Dv7VBMfC8ajii
kMwkrr62/f+lXg9kEHiZdZkAO7XS/X362E+Bdjprb5z5JUpOQLvZ23RBpc6iaLMu
QuD1uXMtd0LuvyUmXYJNXg+eitAlHmNEA9H0tfxWuZqit10y+k30RDzNbxpEzvzy
EUcffcOGxJNymxAIzCzzVsewQohKmQXmm16RAUXdCVR85Jni3KoExt1bJ6cnzEO/
7MBDd5JBn2Ja0brLsosISmFu7Yn1AlgVv3fY2yUPFubjU2WhmUTJItrwpZgfB/cM
P1NUz0OYn3aE0ndG8vi8iFWMgrtLB2PNWWYZ/FGmSE7SlDYIf692KKkHYvTplIpf
7oPDTzTvbrX8hEgjjmaL5v9qBzeGiImh5+HWLYVli5yyzjTAsAT42A7YKtgRCbk+
puVE1Q5/IPonPNIhMVVOmpQnEoU6PcoWgjDuAzUGPPvZMKThGUBaA0958o0X3S+8
BG8dpF/YLGCnujUWDIvaRN5Pxp3Wv72Kt2MwwsS+1xlDwx0pDAQPvAwgWKd8GtQr
QoOKVTMokxUECfOG6Twopy+eOTekYt/y82N+by+HvBTv5E9KGwY1okMepWB7Vy3Y
cECPA2/pWOTl+ccWhWWIM1sshgaQeBhPJ8u6ixk5eV7U0AEJACx+jgz/5xQbn9S9
8apZe0QF5inoALGN4exlBknChgPv1p7hftgoN6Kvkb0EvNn0k6pVYZuWornk44Wm
aVRisH/VxJ4lPSHtwiCtQRupwfdR4gxIDZTjYFfrKLe+VFxy1bjKkdJre6QN0XH1
lUrHpbkrnjBsD/O7oFwL9EqID+vmgpTJfd7hnvdqVf7xKX5NnUJd5DJ1Pt50Nxf7
qlhEcaWjPMnmpLzBnjpBgOliN95mpmshsxlB5gn0WCeNIlsq5aS1KtGfdIKRCfH0
aGbpTpDJ0xOv7WntjvsHa8E+HpUPkYrTXv3iKZ18kTEbCLepD/ERtfYxRr3WceDR
eu9GqkrtcLUGTQaHcz445KrgogAHygP0DZLlIejPBGmpZefqtrtHRrkT7/uuzc48
2nsQfNJfrKs0GM59N+0Z9nFEFqNtMCi3AujNEqWC51KUJDcn2MYLYOYcT4kH+j2D
WxvlrAYdFWoxJoQ4usuIFyZ7JEw++qFXuzrCS19As5YWMdCSNp1D5p5Eo9sfagIm
3c+6Glw9zA4T6PHZH+04I5md7bteAhR3mgNYArxATgtbVrmx09zG3OOe0HtLD6uD
SoQsxXFJ56BKtSzvkUOnaPQOSnEO0TW67wLHzlWcGGKV+Mskj1JtrdMs+d+q3Hv5
+Gpa+nmgu54wGm5r6Jjo3XiJaGlN6qGgOaUvnGjAIPaWG3Xoi2i7OjJ73IBK8ip1
xRZhsozeuTY0nKLWKeOJYnCSgwhhs8tVc7voFyRuA/RCxVdCuCuLSNQTQbnb0pAQ
DtLEn4Q3jG4cW/zVLdZhSPSifTHcEd6h30hb57+5VhLma2M2txs8aR8F7W1VfSXe
kBByqBSoHGlhWjKDpFl3KR2HSzhMD2FfzNJC8+MQFyNYUORYItwOOD2I3LJlQHiE
yasbhG9Lham33lYqIb0ZV7SdU9L7cN7yI8hirj9U0/srqyuJd5taFfA1pP0Ljm1A
WIFcgomI6ZYVbf7qaoY2QpBdV7GGrsIWQPCuhnO4M10jqIwiZMjAtQPV9mTrmFPK
KZC7werFBpWMtxdJBxqE+TmsD7hOziwOzOagmEMah9q1Vvm5peIbC/NgTjYPU1KA
ElD2H6HSGuURDl9AXuEjn0xv+TNeE8X4SzhluIqidbUHqhjvSa/VAEQY7/mVbjtC
ORgrX03LpMpurK+KeqBx1TJj34KB7skl3Kt9bvTqaZMfjNTWGg3qDwNAl3DE63FQ
+UDF4cwzeq1WS2BzvSEH//f1QyI6+XsdTXS13a6E7tXK4z3mWr3qrTxEq9DUYTbw
SewTnFrtmP78tVOg9O3eDj4ydAW3qKXVeTPnwPdsLgrUM/U9cJYI1P2GQyIxh+va
XJ/Vtp/oYL7YxmronINvlWHtj5C0biMpLpQ5W/CbDmzxqhRgIVQkATaIdvYQR85v
dGCERHy3TLo6p6BPvgBMkqZ+K/hBbPusQKouDFuit8GtblWXJbNRuNSdCxmCeBzg
4Ec0x78FKw+gDKjuoY1Fi3rQ2mHgiiCNBP3CMa/114keVnnyeRkwjOc8EWzUM8Ju
QQtp60o0TrCsB2gwCsf7zwQjJ8Dn9+K4ODlm8ZPoWfStq8827urW5mUAjAJcnHTM
73Q+62nikLPv4e3kakT6y4uBcwgQYYN+ZQvgW2d8v8iEIdfN/wppU+Cyao3UnClV
kJiA3+dxwVAw1LmrRQ06RDUgvkVyuwSVbZv189yzZmwmIF7K9/e5Ccu3CSK5UBHk
jpj1juhJhwGGKgkvbTJZzMaMa8yukxfwiEE3QhGVK9KApwWwVrGFIRul2xxXWMmG
jUDRQxpTfFTejQKbKnI7zC40nMfZSqvmdyrt+eCQqmIOP8lfVilzgqvtIQtM6pfa
2/d2091U9FJ3Ig6ql/d9eKyT4gBCf0QGM2pvDzSISZibsPPo5UoXVwQTJYhomIcv
GVECQemeBeRgcpTnv9uylc0OO15/uAfIwjpfy15ssXpJtQ09NFEs52iRwnQkcuqj
FrRhft53OM4vxTll1cIoGgapmlfsEj9KLjsDWgSOawD93bBR5i3OINxdath/H1bI
M1LcJa9ADc8bSKbOIUhxVuGpchLhBZo9xPhx3yX8lVsvmQ2LCrIbfBKVifKs3qQ4
JwAtVDlJpHJ0BxedVtHnksbpZtGmeaNlxKUXHMWinZ9nLv143R8Q6jNmmKxO2jaj
Wxp5cvA4jGJSjbbuL6LtfrZ5tN1M8liMynz8jLlLu2MUR3lx/YecJMCyw4QKyROo
Hi2QPTuS+TvvjnggB5BibEBfk8Sp2FuSOJnFdSLUomSbj3TdIOLvib4hZjse9tAq
+uj9Q526JEHn2aWpRMhwHOLcwU/lpxE2v0DHPhhhzXI9ZrARH5zTSTv29bcABIM0
CcZpdX2KE/nrIMpq2a8A/l4aM+aq0GAeLGVnZ+zjCzKgX4248xh54BXAXUG11PKm
dm7mTTA/qGqpA61liXq53oSJ+TlA+ZtLGi3yrLQrz2lqGX9tlf9qDRCi7XYhShdM
hrWzo9w+dBaderXQUX15hpAKUe+Ys9WJKA3SNSdzTjZlvWF4qhyb84sAD7Qk2si5
L5D1fYvANN/MkGDysiYMl0oZ1MXwx7t4sVS0Az1/MyqaeGgjSPJSVT8yFC9K9Ox9
YHRj2enEB8NySu3qBrskU0FHs76de0eb/+zI6qQX5gTqEtLzJ24MnMXI/iaGg7P1
9SU3kGSDjKI9wWbLB2H8c/VpKLBGcQBlCXrqRXiPbyyEYsPKbPcyRFmx5v+HQwB4
2Olsbt2aB/fspaDvu5wFcOXFpOnmpBMSEmEAKpVTriRNDEX8lk2lgmdb/un7iLRq
NWHllo3MtFdFBQ0WhElJpSV61X25C32VlFzTCsKRl8yiKdOr56hfUupyvUdoqvFy
uwAoZFybTOc5Is6ZRGaWH4s6NDCA8wSfwWtZfSv6MgCz8wN58ozb2jzmfG8RORB7
QARTKhaxUrevUGRucC4J87l7DfSyABtq13VdQ7bPP2RcBwFFFG5bID0aUkBIJCi9
lDVnQK31TqeaW6jahAacWaFjn9MovsrcnbzzPECzYhOJRcJ89+yYxdBowy2Wx4/X
krYvwrZFOP14m2T7LIUBUar6BFATpfcH6gAjmYEpgjU3wJmMANuUP9U3qg3kf4Ue
K9j22yvLtMpxbHDvV4abqiAflAcrbkFSMmrIQ+zHNVSXdfPjUbMmEkI2nXuZ9AYy
RNk+9LtESHdvCXY5DKD+1XLG0K1NTk/ZaAQ6tDR2tH8Gsn3IYNS2qva1mQ73Ql7Y
KJE0AQfvODsmj4yLAHXHgt6x64idGjz0vVnSkbjQefP+Jkifeq4AdBCuAo+u+HP6
KDacpwjbKSZLmhkkaFZcOI20SFL99QOJcZiVrjaFnFxm9QlTzduTF+wHav/xUIYI
2RL8qTZ7GZiqtEzN85IVX0Lk3FzZcVxrFiVvqKWxqpeEh35G/ZdAGsV+ZGQu85+1
8rD+sND6WQUfMDMVtxv+lhlBdocD1OwHzkCn/icHs2I0AKOgSTXCnI5VREU2EEKw
gm6rj/NKi95t0DA+kxvQ/BzrvTIzkEWHe+X+4dCSs92kO6EjW3hJddcCVjIF/7O3
v74AjU1FiwtLPOHI4nzDqU6zDbPhTO9CqDBFWHmbURbpgdcYWB4D2hJxfmgBsC2Q
YpxguGYzLLoa8YQGO8bywrniemVPsqfkBySKtHLeT015Jes7sFfXhxQTbG9LDY7k
1l/4wxWG3043XFGhkUwvHVtQu47ZfiTAjuzAtmw7pxzRFG1IfOtPdyjSG9Gi72Kk
9q8LQzMO325B71vvpImHchV9PdahbkRm4SCef56a5frXbS13VhOS76d90jxIPrQb
XNwReya2dPn+/9/ulN7SGuWE8J8klMtBtokT3OsFE+jn1j43hyeb7OWVcLDADwNl
SuxVzGIcjWIr0Ukoi9JJwV3Zi3K5cIYqw65Q6UH498WlX00IYW7JJtZR4X6PUeWD
cJ4s1dkZC2QA+r1q9eSGyfjyJYYG/A5Jh8ZNkawThvBXIjwJhGSXNnS3uYmYyNXG
OljLK2B2B54t9LRn80yjlYIz/vX93Z7bX14vuOsHx1XB0ooUbNnvUS01PA/dng2e
eiJm0q1L9JOjVhPfXBt0q83mMYCZ00EMV5TUyT2gTxMqaMalAgCcU8w90OkFPgL4
3EL7ztUWXJY72l56Hswi1ugj/U04XJB2KHgHBvdVZZGiqonj6JcvNC9KkeIv5QoZ
xCV8Vrw2r9B3HGPfbur2uWKwOEj79X+dVlnmbybVfo8UDsdRjjI7Noy9Vh13zFMH
VbFxBFpB/7tGkmfcsZZbe30+6qGFyOHwejhHmlZ9yfPN9bKOCCugOGnBAf20ijcE
ARY3aixpFaJNbt99qVhf2QHC+tm2jaBV2yRgcHeLRSiiZidXHMa6nfkjNxn8P5ve
8mdlTubx31K4Jext7DRoYwgN+CwPBAxi4iNuaYMYWJ5odPH0u9rZ8K/taV/u55ix
pCMF2lJkXkAyK/Imk+/d2UEeB/uhTemTujB6QWpJyj38i0lHBdIyxj7DT9h/gDHr
uwDAubheAVOrO5gyeVh5wYtO41rvNFq+nmurq3A8slcULVgDt37xH+0r1HwdfxVO
NRQGVAXj9GUEeKfmf7yXPW1whq8F0xBTA9PW2ZwU9Sp7R8aYkfa220qGdkp7yWpd
ktkVhxwhtl8BqbGqAUm9fsKNyvEdzCKfXVJyjR6nEHrPh50BsgKVAN3TnHRBfgH2
0a+6WSTN9OJQU+bXfJy/owQz0b9bkd9JY3SVhCBdTAOz5t+GcHLsbDwWzaGi+1qD
wEa1OFAAAZlgX/AGrCBHiSJ8VKN9SAv5Fleu3n40Z2xl1VMRjZUr+DZSBYsIMIJ3
t0iBJ6HnOh2XwlMTEDMO9B3NIKB+RZpysj2cv/pdVtoCDDGsCNiywg9p8u18uwQE
aXpuYC42ddfzyyB/nCMAQtoTZlXpZfkztTZUNKWdfRGb8wLF7NKxkHTax/uO6Wqq
Yu+xs/KDbd9m5phgEm/tMIpJSKRvTpw8QqJcvioRqRlw/Gcvc87rsfnK7BmFWeRG
/Gskfr0acaaJBHlagiwd/eUag5RSki7s278+6tikBCkmiGAlYj+k715PLRxtUQ2W
8kk5pkArs3omFfem6AJ1ooZziUZ4/xlQUI0qRWgRETY+Zehx6JNYeVqjFXzZrzLs
PDaKjbpx9ZPZUYZ70S4loKwy9B1mwFPIcLByewVr/HCUULG9p/RB9pgcRdlsjI7b
puapNi6bYxPyNd4fMD8SowO7v6sVyHthp8bI686kx+2xdz4uLvOK8fKLI30uqYxv
jZxuGNj3Olx00Y/JlVoueSKdvtmqI4s4Oe2yzGTxIC0Bu/Bz5qER5T+IJiJ+ETXr
Mlj6gBTlYVou2q4Z7VnQe8Bmh8K8Lx1KXC/1DVG0DgZEm3PQ3KatAvFzxP4wqT72
H2UXOIUxf60WFAMdTmoO45D+FP+kiLggd4uo1nnazDMBJZDKlVgQIwOs3beOH9PS
a6MYHir82NfRv11LEwOfRwKhmd63DRsPqgQlQ+6/3MNhRS5GppvOcFw7NSE0hTj4
FKBKEEukeVlzWkr4Z7+jjMsHJ31RDkD75ckKQAn1oorE6TyRlKGRtQoOyuwsN6Oe
ZjqYvb4iWDJyIkm+I+pcVdLv7JGyTXcELhJLXrc+SUxhnQR82weEoPh2QAVitScP
g2l+7CRcyNruvTRwARwnjuXJjRM2FeRGll5zkbA7LyhbQhudJntrObhcX2Cgx0Jc
Zd77Xc4A0Su5Bo5ItNbNKcaHiry8cQnyOffW/apLiYQu6ELXIT9He0rZD2AUTLSe
BXvlMQ1ojqSqGWcO07T+JBjH8kAobf4MqD3K1Nqb7bFA9geZEsOr587IKScV/JCB
rlBuJ3+38VE8Os+EhFN/RZ8OUWvxncv0zGx7nHlXY98BGZG2dS33kSvzSPh4B0ll
muLnoMFbm6Nz72YCbsEP6ERdcFwcBkggZtEmEm/DvPV5CntNlJE35gmXuclfuqqm
D6sDB+fHyYCXVTqTEDgRk4cEI47PjTyQ0H0ClUMDDZmJZacYL+LPGMDM/H2kcBtj
1dOvWJP/LipHqgaTnMeP3t8B8NWMWwdl1csZoPw0vwgE+LG4AZDMjIdiocCnMi7z
WlTZ0Jv7KuxJthbMhRAhwsGa8Q0xMqzHhuMYkcJcC+Y5C8sIhAnmr2EYhklmRyto
TXp6LZxlCjzBMk8WTPmaptPLEQ7ABkhW+tKj5n+K/7vZE0HTeTHm924fKL52upgN
tpuZFCJ754LsDqpr9ghTKRjPPrwDKXigVAW2oTS2b7t2JaqWgzy+Quw1CC5r0k5k
0E2Zfu2K4d2X/d3QchqPpxX2qhRx9/D6f4y/4183O6KLeAONhQBOQ0Qc8ONK37+G
kmkRpi6h93Isul+M/YCI5mur8XbN/gXV0/BRCT+PdfytPW6iw6hquMCi1WG8W5bs
HI116rkzOMhVB7y2pOPLmuclNRJP8ssIexeZPaxE5o4eEskBmu1Bu/i6RTV2RdEn
EbQVKwEk9IQr8axBGP7xisEqywnj7Veiiuzhv4tK8+lxr0OHrrNaKoGk86xuZrpJ
1s+mv11XX57ZEGnl/4pwP4wv3hM371GziUrVZX7re93T/gQWzTjgtL/5HA/aBAAD
pOj3IFe/KYXAyN6GE/+Jt+lHvF5BogVlJ/5eLPdQqi+0eI6sE69py9uLYaOhWmUB
oxSVL1W3EMzcGo8KORG6vWV1s26D3Z4UsnjrXJ6l+qu77AYOlCAbk2E1SXgt03nk
Je7ZzFI8Gawnx86LAOspjgh0Uw4OXqJSodcGExIcq1VfKyz5iIeMNDlHuCxoHPxf
S8a5VSY60m1ump6BdP7yvqNihjDid9kfAOa3Hwqr3KSPHlNxJLTPwicoDkk6xy59
3avIuh2Yfjt8CAjci3f5dow35+rRmqabLt08ZaLP4wcjN265WDIsS+zPlCxGhRdJ
UhV2r3mECrGQWULpKlpbBlK5rQfArDfjCdz0iWl4FwAvVEkOdUxdHeUBOuh7yW8M
3PFajnO03wvQ44c/zmYKB2lYKu7lf0pDQzgwy1rTPA1+l35h1uhfgX6rinLXkz2x
qjY2LvtYuZrj7TWySFob0O8haEDD2Cz+lTOlIeAwoZXMceBnIECiRhSfJXuE29wB
8w5oVOmYXs1cwEL2Q9zfngB+Y6IKhuH9HFq/I4P4EIW8HvzCr+1bN0CYuZrvkdLs
cWdokSsIBRujAjiv/BWrLwNVGOdSDqpqRXWVDbCAm3SZLgg9q/swlbDMj1/JIWIF
7uXS7St/AXMEvf7aBxCM+HY97w33rHReZUZMXs3jSjlkaggqlKqwzGZcGCNqZEC1
Zf+KQm8QjkI5XslQUoyuGUD0f3KLw+KM6fzB0QvHwGmqk84iWsvQ0PSVgLYF12mu
r2QgIqsfeJciw1h6PAOerAkKambpjSt9Eq/a37pAEWUq2hrCyj4B60tKCdnY5Lq3
ueATxnSdsP5x+5CV8tYy9QJ1sdO/MCSRfDpp4D3nCce8LQRHzTPVBWgWOyqyQlJ4
kBL+SHyOliY7o1XimLRv5rezWU+Nf4DeC5iHE4RlPGGIAcIQPuvT0rszfkF6XR6T
ZhyGg/KCIPInXqqUwU5tbUys7adeYsWoENelMxuq5TvcEh60M47gC8Ux7SkuQvgT
h5/2NGyw8zhiXQ/FJkVH5J5ShrDpYM1UOO99/eTMrSevk4sb7kF95aYlumBgNKEX
ws9VKX/egIfoTsmM/RKqnpZeBtUvsifyB98mAvAPURBnBR+zVw+anvfjqev77LR+
OHgDUKsO303TgwvTx5iorZhLKGkrsTEUGzGlxfKfb3dMsnycwMjj1W9bqNxKDdvg
sZvDx+vZjOXepc/Ryygs0f8d207rfpOmFJ7Fz6WB7ZunMOQkGQxO5ZpX64/mVKy6
nMH+daqnAN0t4C1/MySUEOFZLtQ7vTuLY5ypoUdiE9jW6VdYEhT+Mx6RXO94dD8T
qfaculJ7xnogl5GnhR0MqwPoC3bu6DM+dkCAQK3n8DlmZxXaOIP3u0/9IEnC9lve
7fKQuh7vrWYPJI5/kOhEpM8wgixNfMPO3YBIa/agZQJpfo23nJyX9X5B969Ot2Qb
wJUHW6AJFuUcQrNM9yiTRoL//EMXy8odNs7z2Mx8BhMDbHulPKEn2GpKJF45wGLh
M6uFZvLNNNo9EE99iCy7OlQjIJ/uwS/2jlDOdXBZ7CIi/YT+acjR7YYkll9MGshM
AwIPh88PUQDaQRMAtz04BEQn+AGEFj9K7YLdJbsGiyoqtWRUdFk+oSVckj1+MTKD
5Lz2Z3EwOeBjeNLvVXpC8nolheXalSvy0+u6IM786YMbaTVLHq8rjKUnYZj+cm0+
SdyHbsvZgo2nlBgnM2qxokn218jfDsh5wAS+RUk2PZBWT9gv8rW+Q+BUP76SEtVO
ye7T/6u7uEypEUy1lXforami+M9vIwLE3pYRnkWkfTndICE8vN38VDoRKEM0/FX8
zGQx6CP68BOJWR0MWrA0b4r0Mu6TvxWy33torq9IhweQ5e+8IV/KUWNDmzRDMTpV
3El1VgzMzmT3aTZGvjLnyTGxqZfVwQTyZTZ/B5lZK+wArDZAgQ/sXihFE6Mjmn5l
UnEtDCHORP16kfBnRPEU2+A1gg9p8ZSoETkMoHGNuqxP4vgjfs/TW59G5MCKKUcB
5unNVdUIbG6t4nJYS0L3d6rTO7fP/5qN+3bh15dOV+RG/4zUaASQnna3OwVYiRas
+BntTE5k89NxSXk+klZunueY/gGcVdAPM6JeSxUQX6yQ3EtHw455XJbVcfNw7Sg/
F35dEFyqChEYJ6glNmY5n7FffCEGhXI0qSgT479TmljH6iO68SPDm65yZguev6Pe
uAUtILqydn1AqKks5Bc8i4FiAKdq9ThYfril+sk+NAz6Mt58+eRUTthpT86iUYhL
5xmtGXDoDhbNCDqpZ0oivw9CPyu3SD+vrdVyEAN7sMSgdTGW0E56E3pUIs8z7vel
/1yxZk+oQFpQNgjOOunqaKTbSr0WnXVZtgR/3HrcNiPpyj4nAE5cpQU9leGSM3jp
zzy2QYl93MSZrirxMqZ/Mdyk4mHSkzB1YfDv7tGW6qMaVcSbmoVkRnahaxyVzz+Y
2VagqQKOzKSYzkcc1ugvHK/lfyLK5AD9nMJgzrboXVU+aH0FpIFj61WXOQPIm3z+
xjPg3ly4OOfOKQjdIwTUpivHKX3ixPXzHt5i8C6Pa5bCWqyrOILubKzezLvqMnyr
R7DaSm1cBRflFzy+YFj/Z6whyokWypASvGIuQtf5YIFcQIuKXsgc29j+6hgo0121
6gSuPFXwTGBcRTOFavv/OaYNmzqv68X4F8jhltPea58LLFVtNN5ZtamSrzQF/+bW
1Cz5krjYc6FWC5kE1OsiliPthTV6e52KJMrXU1e3cIVldl+R4BXWRBMb4LQwDZ1j
g+tBZqSYmnCBC2+GeLYKnMMp5OImSAWjIMH/lJdaOVZofKbZ+2c6KycTOZzlgsQy
b2Gj8MtDXxVjU7OaDhSQp/xuwlgU4m+wiMkTzGuPJ8aeveWN8YOPUWU2H6WcNolF
dQ8Lx+qcXMJaDoLTZBC1LaG6IxMzvG1k5EcHFUB/bPd9TvthrMpJhZWKAPP6GeY6
Am8XOGxNfcqLBdzmszBl2OGK3xkx9E2MuN+Spqx13DWAQkz1DjticFGXQjeN+PEF
OJVItXlUKFXXwAFHeHQmeSexYxNeEZnbWaN5w3Ml81krbTj/Dnx1mm2f7pj9DKQ2
OlaQ7ZqMqhX4JScWDqbu4XbrS6Fv3NBMslZ4sTu8MQuot29gSWcleQw5/yRH35i4
YFFFOIhd7KrZHAk7sRDD11aIG9pTlvTqVHAoOhXKiilRwu8k+hV+oQbz8LhXuwkH
vFWDHa9YQ3yMAPiLorg5L5IUhLTLBvdBv+tya9GzNk2hiuDMNHhoYO5tWQcCRkiY
7YVvT9KSjMpQ13SQLPHt6oZkKmoRC5o5I0JxTv8CYlpJ+wYeJkLSTbCQptf6ldtE
bVsxXpoi37aR9RilIhkXM5Ce9oFNJQm9LHIhYORMDYv4s6thh0+1jgeiudQ3zKcu
IGZ4wuv+68UkeuKxnuSWhyLkbZrVSDfCq7HrbF2rMJpGvxZYdvRW+miQhL4EPz76
VG5Evamswf/lxopTF8nWPLJ5fTfdVrObll0uu4PCT3PyDZ0CNqynG8TfBeizaJ9f
qh3hKBW3HT/XJdlBZl7iGh277d66CJm0mtq9X6DzTfF1mg7PeJ5a95yRXZCwjEtJ
rjAjQFAhFHsJMfhSwVKF5Ec/We34FSnO9HsNpqgkOsoBdFvcYmgr06iIEPyzBgtO
6PMrM86A2iiNr4xQyrr5EsNKr9kJJB0Cy7bC5hc3INr4SyT4XZlEWgcMlJTE+kjs
mIZbbYYcTLpdhKVxmRl5L5fmYyk5yVl+HPnWUqaRPCZ6nC8nVMDQeEp8de2v9/PH
+iO0it+rGie6qT15b5YXf1maZbFZJW+ElPusy12M4vgK5dat+Abm9S/pGMskoVFN
/CgN0+y0IxHIg7q76BhZ1AnF4UEg/S+5+cSguAFWr09y9yTRhylUL3dvVFRrKFnV
uG4uOApabZTetav4rgs9CLst7T1PcmhkLuEvcqEPeWz/+OSWrjk9mWV+Ut13DKUi
lF8L+dfD0u5aMDw4o9T4Ebc6zU1fF+mGhfEhgedyUp1qRCnzHz8jbF6miwFyxZnM
WimPfKj9pcEy84rfqAcN8j0uWAeOlKc959IHyaPcdXUO0XMZMdH7eu7041tV6MiQ
Ob44m4GIBAfQS5OkOn2l6YtzdUe0Snm+lJ2ZLPdUhQejvdl8jWsXba8ASm0937oj
NIiqgtMYfRmE5v6TnxlJIMQWXNJOlg5CxwcMdqkrbyrrheaZLouh8C/QIZG6N2NB
mSoT9PsZf+2BRvzqUYBID2o1jMm0MaqLLD7FH6fWkmExBW+ZGuL3iS+a7FDU54zF
U/DRoUq92SSjATYwEZUvGy6++e6niN0U5kYU6fC6pAYsLyuJjDwhGJPZTMnT8grT
HRhp6QNofpuu1CMmHOfpff2iNqQEBq8UYHMu+Kx50ZOQTAFSKfGzjiiVS8JvC6UA
0J9+iw7RzuJvaQuK1TChIeWC+PxNBacBt/v2z09ToRy1ZZFAPGFMbWE+hMcKBYfz
10IO4MahjIH0EbVPYVaxz1i4wlmcPJPR56jyLMlbaSUBuYXfpQp1JoG4x0hVwynt
13vaeLUSkgC4BOq5eVesd9Sfyt+TizLOHxAA+6E+PxrOjWgnKUvP9IuAGfZ12sJY
r4WZnXNinoVHnqZPFC5dnwS1H5XZ81UYNMRmiGT6Np0SMX7eAKkzabFk3biQYMuo
9PmOeT30ZVqGg31n4k0hAbCygc8UxjLzLRVBjPVs7KFlkSQEU1I8KZWuQmnPy0Iy
lGAm/kc9VMOzMRUB4CbaSLfcClhndWmMfSVtbfPhWs4ZA6c2F/nauNvBpCpQ78P8
oa1sQZCoxJCzsVGlsM7e7bx4bnF0dmx3a2FREClOZSvaMgVetXbnbveRh5kDgdG3
TQOARZC0JKhgqN8QurNTs3bWrwSkS5Fdvm6gf82CTZlrZBhBBf3oKwosrXwM8FRN
ihpQiwjVMdTSsUZFw+MQ/NXNPYEm1HdPvgxRSELXQ1WkUZjEDzrBdFi8+TShpJIZ
gEOlngk6517dCntXUTGkKUuhIvoOHITAAjZrSWyimBoWYc8IJE9g5/PXMg3CVsC7
bcDp1/chdbQHyG4HLg/eTj9i9mSVPnBz92zEqdBSB8aZ7p5mOKKDCCHaZI3nYwPZ
AOCIt0u3JOEwiRkvbV3XoMcoLHeq5ihurKTwojX0+W8F6PJnqydeqYVmGsPkm0jP
MS5UuE5aqx1yCYxdwSs1OPpHTjy4/OPcY6gKDiVE1Ip+zXLRDTcQGCgvDTXT9lNg
weHW2GxFYO23GQgh/kXIuTKNN0tXFLLGVS5tHrQCb6ColtwQrxGnS+o2QlpAzXDO
Xk95tZOCZm7QlpCDzFAD+Wt/qG46hS9VSQZDsqyZ3cczOe12x3Ylcx+AqIQiHHIq
KqsZfqK1qehNTVqhgVfD+Zp28FLxqsCDs1fHjS+o0fPUrYXNF0QkGct/Gx5/lvw0
MK5srFjHq8HgANtUXUH70srTcEDKr6ECuozZ82WG4wQAwGz874+CMdC4FwVWCz51
wApPYU0+mPhCQVe6fXBb5c50gnrjhGZSlHMxqQIoDKuwm8qA6dDbFsZpk5N2UoVz
y0rCpAluUNmYqsorgqyhmwUomolkdnt98+Rsg1oupHSRY0Ul+9f+/irUlhn3U7KM
NeWEgdGzBeLxhuP1MLhGBZHsLkQLnf+rpqKsh4eyB8ZVay8PXaxRZPtE3a1HgTox
YERAsuFkHuCvFpz8WLEVX+iE8DynVlXT5/RldSUK/iohssQQvdfsihE8RStPK+j0
hMB511C1+rUl2GC2zdwvgGCYjT/ulEcRkbrng3lLqRjI2Y6bDMWNGV9b7byHRQs5
Dpn4DvKexR86GjMar9Il1OBpUIUqnPFo2rq59kh/X8Otdz8TFl7XBk1DTIVDUJXr
XOlor1K0DqeDSlbXTCpsvilRFeFfThfcLa+1L9MS8LOaGCsDXuhWKM66QA8XSUnY
vCOVL6AjY5xoS7t7Fit+LIwPPCyomxkerNMO8GmVabVbzyCSdBzxBdApo0YXa/5R
Jl917oTTpA5fZZqQ42dIr72SJGnbTXc4Yzp71QZjbLAYT4TNP0VRC+Z76SFn6Htr
e+7bri3PRXRXIAOL81gW14urdP1AHA5vqq37XtHQ+J+SWWBzmLM1+lE3QlSVfxXJ
38YpzzZwIJYSu4V6waFGI2TDEG7fcskr9hZMxSKh0+qq3uCO25AFIpzuMhME4cw5
q+Qm3Sy15ZYXIok5qpyp9X1ZMcDh4ZoK9S9oAjz/dXp1PEG0H8PPiPLCPprEhjHE
WLgtXS9m8YswDyrmjJEbf2lhIrvnjzwah/Z+2d28GvTPIFPu9ZSmEjMQWYDVBYAm
plk1+dWEie4MQFQSgE7zfan0IDybgGMyYSYxmjyLRP2wZkUPseE52AFWL88O8heP
0MzIqk0yEtA81wxzwcnv8RWi1iQdjLOmEsr9a3u0HC5SzIfYYeCHFHhBYXIwmWPN
W7cSwiJ6W8kVD9GGgTzsCuwyYi5Pm0pdgcdiCd5ZNuxVv22TC559J7W6VLBYQXRU
8xgqTaiXKCYzyHgyIx6KNPAk9qAL0W26G0l0KTPW/pgclGtvIfJdzw9dyBDjP//n
vV3yzURrOab6sHhxWweTeOOeSf/L6WCSxYxYuGwmksFyEYsu8+qA+FCnZYBXCTy0
VPxa1Hw7udEvIOiLJllty48k1wBDRPC8RDvscBAGVZeqzPlJcFZeij7yQGS5bguf
26XP6KNZfE4RH/MPVQySbwIQ9Ulll+E7Uji33gnOhlqcFxWvInlVw2tm5y7Eymq2
JWO2Fz4EgFH+gWKk/StklYd+qvxQ5RCUoC6r+4KMH8Uc80VE3b7EtUQ9WgmdxOBx
0XUOr5Hs8ueiRXcbj8rDSMs+fYDOK/IJfK0zY9BkqSkBrRgXuAkik3odttPX3efo
LwldmL+nf/yDguw7npt0Yg1SJdZK7hsbN+NlPUjmalaW3xk1SlH+u5mCAAWf0+Bm
zn7t6SFYXTuE9K6VGdp91+RfjGy+O6bsHUCowjAf1ClqO78Lw22kRBSOy6N2H6ZV
tf6y7qBcY3MEO2Ft2P2M7DmvMKH8f0I63HSIOe93lLESB6Xcrw41Kq1/l9uPVLHK
7+9S8I6u4XoEV1mQW5my1zbLFmcRw90JiGuVoltNdYgZTAZnJejRZn3qY8z6P/vd
rY16NlNI3XxtVh+uzhTra4E6O8CRHgq6qCpZmz8AUbITJlbOTskHecMuPcq4euWv
Cjts2lGvsrV9S4uvrP/gqdNlE2qaLNoCOvNQseTrYhqgeAvIVORQI/4AQTmVB4N5
MkS83LonYNXyz82ILfXKue7FU9DjO5vMkAu18wDQqPDcB0hHMlup5IO7D1g9PSPO
ycajdYnT8ONFh3C4+4RPRn6AJcjy/p+mLCDtL/tRuwd8A06utSL2/58C0KGU8PsW
wRUh4SZ26bx29Odvsf5toILAeeiZeFrOMtUoFdCZj4Wtw09g4M69FclX5GQQanHQ
uF4VYs46pupRQuPmSm0PpPUxNz9v8wvTJYYXUDep4mErydHzGp9VAh0ig7aXzM/5
UFKTNm7ccLv686vqIyjcvjqiraW60HjRLj2A1YN6/OasxNcZfRr5KOpNtblLMiWt
1sUVpMCFm74k4KYVXr3Hi6YHJVKPTVZtPkIJ6MFvlDVMdJIzQtHXDPOS3bxp5dXO
fhRcqSfjO3iRShaooiKPEvNqzCCOyUSYGt37JXcu06TRFQOVXJobdAAO2IVn6sTT
TbPMcamIldHODV+BlScTT013zQrz7wzOhuOJt4FF+OLi1AoYI4LWn43Zr6HMnJDj
5MV20p0JM32tjuoUoVSfGgR64hjIzsFvHYYh/vTHwQTiwhVP+Icrv6CUJjT7DPjM
HOKYR32D3s4dLuTrsyEQvCUOvitOFaXwIeJMFs8JXWIrvxXzh+Od6hHaClXWhmp3
1Yvz9etw2SkbRdtoYWqenkfW9xLhZXCvXdK7ixZgZHlNqrk8FFnIxuuZpffZRcNa
FtROFlONoEgqdnQNOTlUI2SoJErJ9ByY7sQ10E/Wa7bdTIBjrmbaGTgCavEPKT7j
1742WOAVuOfUFPNqhHE08iCREAAKN1aTHQN2xmR4Hyhp+///0XC8HmKWTZNhR2z6
u1VqDUvKwMBfBQV4wCr62O+Q4ZyhoVeZYCB1Fzyt/90n723Y3eeUqTMimgL8vGlC
SVr7T1hNVbcPO+JVV3imr2LGKDwnTBnmavHIjrijsfItdY33Y1kgK8bYCtBJlW4b
/tfAJfbK5IKnVLyd6ZCLhW/XNxOItO3B3wEoJaHIl/PaKCx/DZMyarqZzzgVbPo1
eGa6vhdXjpFiZQEV4ZePZgeYHQ9ohFDbO6ojMpXZzPJCufoUSCq7RYZo6gPKIBie
7KYKgz6vUGq+J4pgLmeyxm/i5XUkpaAp4+FFezS0ajs0y7Lo0kRXfsbl+FGcc0MX
W7tL/eD2phF5hUd6IojLKHqqCSj00IicwbkQ7/wSy3OjWW22KDuILvcZR1+u25yr
CCmNl2sSWxDquHMwTl9MvO/2NQN0A28cLnP4a0Ou78shP8RHh3XAHp/YlU69V40e
OLBHU33X/jsQwuf8QF7Io0h0iWwoso/e0tD7cyrBmQK95eEOGMx2gppqpRDsaefZ
Xv402CBnju09cPMcFJK3DXOsNkzJzE9Pla/IXSDCvUnMI55gBLV9kZhf1AJIaPUh
xHkN3ocher95f5YdyWLD6TKrmB6CQ01YDVnD7LrvYqMkEgvCeOxSEGdEnmIksGOi
fwbE19WS0TPxZJQB6BT0sbHiRuA6Pi8JRGiAfTEsS+F1hznIbR0YA0ywoxHwN3P9
4ahUtbeyDcjn37pBl6f/JyNFMdjfmt1O3jFNWNzmlEmgmNR+MpwzJ08x5xyF7bxB
DAHHJCFoYj1CHsONxsoSkxVZ5ZW9TWBPnNZVbPqv/KRugCtAfclnkdJgsarEWHjM
wmJVVaFm50IxHV41uP5z5DU9+2jq+7Vk/Srh4F0kHGONj0jmUt6IqAY9dFpHwuFW
oC95tBOdgzTmbbtwd53QKxb83vgC8NXGqXLXuH8MYL07lWuF6UD1g8TCnP7T2qox
yegr3Zi98fqgdeLzQymHANH0YxrHNWVy+l8kw3CTijNfxvpZqpLMyH/RZfspko+i
UICi6wI0yxQZ9inAeEd9QzRuZlNCutiWjwagExyYOfdmOI7bL+z3byWJuZoa4ZpR
kbW1tqy76mcp4vVw2+y+vn6dfC1OhzVLQ9sbuthhC3phCfTZky3SAiy/Oa1XeAI2
4OVrhKlUP5Zh+biejZAPpTj7v+S67iZi2Q8iK0fjgrKL3vwq4gHSOcqlML0eORfo
XUoeSTeug6zgdqJsQfelXmDWxmkmAmuRJ4vZ2pGet2WxnwT8nFVWQloLQ51YaX2g
HuUqrG/aN6uJTyvc+5u1/Rblhy9NvreENDgEBBmruTdbUsyyPlenjZmp9Fhbc9xH
cJQJjZNZFAfp/YC5/M5KBqL1vVdBZm9eSEyLzIy5EXCdiGCbd+o/9D5s8vJWiZKH
JmYXgdnKq8NC605c8OrnjUBsFYvxsj/BoSVSHWzzdSZisIjXVPKVAOjBS8AOKMT/
5hYMjNqXe7oCS0DDWa6cSr+mfzeCB5VT28tqAAkj7X+SvBl3HoMRYA4riEX8+2Nq
7viR2CevW1KvVLR3UfKZeekxES9j+k27g3m5Tdlt359su+TaKXANohfirxDlpBoN
P4NrY425Eh9gtqswgdSQyExFTxTzZ2EjSIr6nnweeU0Mk616uI9LLhN279kxTr/z
KO9R1UPjaFJ6VVfHkcZjhazGnNCbEW+iWCTBtUiblhvEmet402A7CRW1BQvWj5ob
+EjzHapGI9X/H3XJ1gwK7D/6gSZ7kJHMEdxkVbHJ+NTSEjuZU7FRw2GfSvGTOm6Z
w2bKbvMYMdsOYFSLLOnGTlEzS2/YGA7HXGUHQ+9RsaETG9aeM78MSUGR6LSDSF5L
QYXFq/tXAexSCcPMAtPTyEOUjPYzhTSP0bxo/C42sN0FfUUX6t0ogMdfpHTZ7R/y
aoc59huqtj8Xjc50kOl+zNZKabi7RF6oWk6PTRPC2Xmu0J4aCcikSQ6hWrb89uao
FqZF30PzwsaCh5vr6mTsURTPjS0cEugXZbKvlN6iINU3OfIa3YRGc3fKJn6fC+Oc
vtVto9qySTW6/7eiE+5br4Zk57NBd1crVzlbeClBQt0q9MAd4h6QXJS75Rl+/E50
lq5qL85FbZvKPYdI28ylT1h1jRcmW/7j8a4s+p47hzS/gQV29NIWsD9uasEi4JBL
WVpP8Hova6S8407u0rBubKoYRkjcVqyCjVn/7kZ5NsMC2xxdM+YNCaX5vkliJHkd
nb8VQUC49kMe2nn7o+KoLFyL1eJWRlm6OpzpugwQaBdrMYIH5xZSrCX07mCljbha
5nMVDWFFZt6+3qBYBS9RioD0MIbfi2x6Gerc5utbbOXBTD6cpMp0vW+gOUOnIJmG
vDEc2GpkExws/F7801CfqmGaHuNI+a/tyG0yphuPq/TxKfCAfVwUKBWMV5Rn/n8j
P/jBgRXsxAs3lxXLCB7tKJzSdj2tRsL6ZzeUqIePQFj+WZvgp2CK+VqUYZllpdkd
yLDj2e8THmw8gg3for5WecBgIG1S8XTUJoRJujyZNpDajlFhQgxM2Idak3c/7I5f
H/X9+ju5JC/n3IkkeIG9iIgfrtg9iElE9Mq7md7GF1szsl+2MoRVNgCU5OsQ62Q5
zerUPLxN2TzMVl+tdkAUYTsqjjbIRKzG1P6oDaVC0obJZD5299FyK2IMmqr9Qupi
bvNrc+Fx5SkK+Z5ExjvRYqmCX/JyI6TLLsqwqz3T3Hl5lWcLCkr2/hOqBE01Vxby
hNW8knQq1DzjtVaI1c5WZBQKfki3cyZ8srJQ7uICV1MqKZ12NMvh0070rdUcuDE2
2JswtlSSst2Mb+hrop9snCYMzO2xK//m70+27j6OIH95PCyukOoHhSJmLiiCsSKn
4WNYr9ieVpBNemaw+/XaMExDHEqO1Y//wHp5ASr1yynR6M0mlxVhFGLlZoiczsUy
KOk/sBecGcQ3FWwaPT9Xm7TP/3MtSb7oHSPfT+hOdsQ6/hAJKx4daxmpcBPH8xnM
uZdBgySsOZZO9uqaQh3b402C9qt/PfkjR7/nEEz6gq1h3ZfSiTYc9hg6Y11eq0gG
QMdwC0/hqAEUfzAencpTy11/H4pMZ/M2gK2MRVjkykZxjgK2RJItfccZvPwZa1wq
r+OLD+/0Yr/EUR8FgVZSvPIUdknE5IbuwsyXju8PmtvsIXGS53gN9Xo8Wn2jINNW
XiLQ7qbUEV2flM4b73Q4LyfZ2HOLDyknWqnP1finB3gbh2QvV7fraY8YXSuo0nav
LYS7Hyv++MQviGzwWDzeX+voD50IcCnZEukvIewIsB0ec0gSh+oZ9ScCevahHnUV
Vr2IsOPybP1B3Fs+75NVgrGgucaKOrrnQuQ0ml40byZNINQaiqT5+vB1U8JV764/
uKiIcwLsp5v6Cw+gJioYwy98aEaHL8lOHBskR8DNM3JPjF9+j5ojXijN2WT09Tyz
6uD/q2vUtsdYZ3Gtx81MQLNSe6uwlaNnpAG4XXqVEjB3cXNwhwXtPNY3qFoXoO1q
QoqC+QMXyfdV3iDe6IpjeemzDIKfZLcef7HfOkytAQvNWprd8qL/dcP+kYEmgYED
pX6xMI3kIr5YI6XLpA/EzWMSvBsqs6p0MQtokYFFi4KQe4OnAlD0joDH+eeSXnsf
DRke3OZOOXwXvUJGHU0n+BV1LOG0ji79UH+HPXdNX5/sbNNgQR/ZkXJBDHe6zV2g
zbvr4arrgedJXjPAAU7/XB0BYg4Tuh4jIe9EgmVlHM01h1CfJFN5J8BLG/hdzdnh
DpZozDK+lgddYwVG3yPaIfdLJJXnDhUQloDjnLbWzlUZ4Tp/XEQOQqn7pgKGIn47
MUQwxKW8fQeDAymhAFNEXR+Z3XokEgXtqlAaFQ1vWJEEt/VV59ZaARRzejebOqJK
LigozNaU15bSMm8WiwrPpKnwEYvEJcGTePdFAle8Da2LMpACYYHVbNYHN8k5Y0HB
ezIsadfQLP5SrHy7Dit0Y/63fWY0VN5vXpG1COGP1cgYFZ/ieSOXKUM3JnK8HVKW
fAV/faExp4eTZ5rVYgkAzJZcpYX3PZ+H29XtCxiLQXv8eit9Km687Dtody0DTx3Y
DpbVWdlatF/K2NR3M2ZQ5jwvO1qvVj9Vr/S6CmrdAPmRyIJVjA2kO8hGVpquvH1O
5st6I2IcKBoTed5g4LbrlpAtAHjARK9x/vJ0emo8EANim66WUIklyb0IwvwYbZgf
ES7ZEgQHguOyxYk+5FpMLtkKMxDh7h9FN+XIO3o6NccuGqAmhACl/+quSGAa2ERV
VH1X/L6irznrS2b6+7283e8Ds0sAaI3/lhwcMl3y33evhxE3PR6BWmsQ+7C4/dn9
9h3+g+1tuCZV5j9px59+t0SZfkDP6nY/IB5X3aLLYiVYW4lKNj8WnYfHIDE035KW
zaJhHftZJb/fbNpp/dgfIQ5I10yFxy45ZbUkab0C4M+jvJUnuinwUBnv9La5fep4
K9RmlIK9n1WNr+mGD7jpks/L3eSrk8jrPBSZ2h0snvh/JDjPSfauUhclsiumuvon
JNsp+uBENCO9bIO09MPYmtcYsvZYc9CMWhCjOpJk1jXrVBI81N6OcyH8Txrd57Lp
AjoBDjrd4itTHRq2ja8WyEyGa0BM8BPhOVr7jvA/L3pJC3XYTYqX6uHODnVkKXaL
GRX73X8Tw28s25DR4aYQhZewCWGhy9+5OoIy53UevyBsRilFYkkMg9xn0e2JbdUH
lsTdowU3WHiwRP/XdzPd3b+/5lwMo7Tzyi5aFgOXLwd/3p0/jOH4g6FYgtXf/CCe
3YWwsiVZY3gP9diCQmhLlxocP7RN+bH5y9lf2+3Th0IsJKsL3BwXF4tKeeJL4eHR
2qkRSqDy/4SSpOZ/aPLMai/ejBFgKtnnt8dEG1qkDLzIFGgks5BkK0TqayOsu3UQ
q4DxqbJXnyqMa+x5U66nk2ei0pnmmk77bizQCv7S6oZoJniMYki4NH14Ch6Wx6B0
CLwZUhaAZ2R55dKUTOKGoE0rAOo19IuDZMBbXOXnL3S3EFVTGhFc7U+Ds1/zbwOK
z7j8R4X51PVaXuuyC59SqNpLB963+u5E6ECCZK5LZlo3HmPZ1hh3kqlBEr5CtkPl
0sdiEmyoc+HGJHtIok0RYaK+D4HmFIV152x7xmju2bukBXNG/zzSFN3k6yKtG7xU
kyGoeEdiJRBl1hpzp71VnyjKDm3pVguB9JZDpJ8HoZ6CQqblpBETg21qb5tQag71
pVPlDp4NdWLsYNAVBMKKDWKH6wqbcUMGv+bD1oGPZsGDoSYU8NMcnoVnzzXhxLVK
xVtQBYTBmjesd1p6pYHXLM3JSf5DXA/lS3Ie3bw7Q3OHllHHLePZh47DsPkc9tOY
b3vNV4KRFA9X98v4dvq/wiQqG3ERVlqNtGwB57AMs0sj8/UN2LFgHkNjXM+xCjd6
MQQNd6E0nuaRYUWW6X2I1YJ5Cqcx43W6M4LTjrO4+nNTVQjM3IawelFGH+9TBX0X
KuVlb0Xrtw1U0jg+yU1zpoHUUe6aAmzPPyXAyT6w5z2IkNClTx6cwdok2vl+8C2w
2BIOPoAwxy+9H3XKO9MGtOvr42iv0GmcRunD8EGEENGCXLUa4D78/vR26aWSP93y
ijOY4FotETXzieZfbUg+CMfwSdAOFg7jNIPf6XWnBiWtSaiD2J4JquRqbGq9OGhL
r81q8zzHCQWRLPkDGEbCAXWU1qcbQXf7QzfvhOpuodgZ+Y/8mXJBCymqzVUKkNLa
mN1OumW4XXkxoj5hwzFEE3YqOy49a1cYA8AcR3nBXtph1sXt3YXChrGBaEmHkXGb
8m2yKuTmAyos227UaHcSPXOiSdjFfU223jX1VCqt3JjxT3AkMZ7UMPhSic6ZHpPC
C5v8SNctR8kOntInmjyt2yQV1UFEettzzQOlNfEPcP00cmdt0wbmmrWAW8O3hv29
w+SSG0D7kzz2hKhtx255crqjzrVTH01/2Sl/6m1z/mFWY/6lrKpHd3kEqkN5Mhwn
1DVc+rV3ngc2UunFywkbAGbm1Nyn2Sr+CN73ADIeDmhTLTlFjLLdT6RcRBEUJ9ha
15Ep9A57a+Jv/HZVSDlUsrS6E6sopnNIpwGXTPXeVvDbLtKZn02o2832IHaN0sIY
gmXFQuqT4+5l1Ja3zK2ZIxEJUfeX3iu1xA0L9Lp+utRQPQYvVfvZpcgu7q2O0nff
55yNdJkINrKXXxxyg1NNG0jzMbpYHM4jQ5dX12oiXLeVejFJ1GNFRLQX+7RocwlQ
ApGAT9wJCN1Z3JI31A5Srab9qAMrO60BEBhO6/NYOGwy4EImKnfU+lu8IbKlcTWA
IVxHhuVCN7LV5sPdoQ6Bd7Cf+IcLRSW4puyKalWAzlwMiibhkTRk3VYy8Yg9e6vI
PNsEd+HahlHIgtfwST7h8e7USWugGbeFWUbJ8xvpqa6dJM3zHjQmDvkMnRlXFnQH
umd11mL7MHlmPOb6srjynx4AKapVzoLnwo7a/ge//dUlHWRr7fERxrU4k2QltEIM
P60phYM7YWWUPQsdvioVdSPFVSvyrZWwYCp5LOkYVQbJ7/TsTsZv3hNPhiMXDBIE
zg5kN5MAg78P+8nkicFdLm+ojmF28GLSdKziVvoWvtP7iFQON4qAGszh3Ew5jX05
7Mt6VtQZzYBY1yw1NsrlUyvXeT/tlpVdC9XnpAjwngcCnRcTas4ZQGPXeqJrUyp4
acFZdOxO2/0qSKu+/09YJpphdwIkWuDKwtgwc+M9XrcBEDCzE92aztrhJRE8dBYU
jNYYHIBH80Vt2yXerRObUT1Z4M3JUOc8HqQzwtjq3Ud5R1jkkHov0/c313ygoXPA
J3Mpa4QJ757RoOLYFejFxE9dLzQH7HdN26Hk0EL4zyW/NZJZIALAfCs9NkhsMdPE
/Y5qGinSTRTzrycpK1oNHCQd5aLFXQI3TR6HgQJJoeVTeIVOVaCwVkLXaiTDUoZR
DpF7AIMfLwkx7axrmIMdwT34xLWVwV/mOZOcpbGQ/hreSrYGWDwvcnIrsY5R+ZA4
YYjRZkTee83Tgw20NC0nQUGMgu2AIlVvY2yeKnWCpF1udTCiIA9QbpsVX4Ealtma
V51bvXqUA/jvOKfj0yE3qNcmZ4mZHRY2cj7DdheBZhgrafX3qidgb8GceGS2iTXn
em6XvaATZTluRrooG70riMfHb2jiQx9Y+JS1T1EnmZCG4va22raJW7TgA14BmFtD
fOSht1UV23efqx276t0JmcKIrYFwVsqm6GKoRiVrtf0RX7HQB/yyLXF/5m2GtUM8
sa/X4/tAJGZI7/df6FeKldQ5CIvapLuc7b3H4SZxxGVBh1nZ3gfbCuQTbEElQAZs
Cv8jB9MO609CC9nsP7ZvacHf+z6NTqhGJKhgOXKU44xcmqyExqIyW7LjVmGw1mvv
oSWUUeCyMMTL0cLanZNpTUGoIktct6VU6Hi7QGsyEm4K9LLxNM9/9Yzo58ugWnpb
HCAVw4EGE6ynlNsT5YO4gBm2Bp9wDohkAt5/GNbF2ocLN04Aqko9AGhu7qKVfb9s
LIfucPMdWVvbSnTxfkQi0QW8TK74YaJEw0ykSAKB7R8Cyc5stCME+li20ppR7VYx
3X+VYK5TWbEWEi3aCt/oiPVK2dwOjuzBUFAOQTxARkYBwe7+TTlk0Qj+22bsCN7y
22bOI851u/vzIJxXBAOR71V2zbc/cCw2h37dpzKwDFWZOHLWkwC7o8kwtACTzTfl
eYQYaPDpNcMRrV6F4yXojpQzMlLuIOBVy0zYV4AEjHmsI7SPsbiRNzKJhoKOwYaS
7KuqD543sYfbd15oI1JRb2zaG72ZOjRbWiA6X3veDnafNyrMIEWUGHo0ysuH4Cnx
RtmSSIZWqZitGlJQSPVtRev2dB+v7LFPqAY1n0Lc5DyjgR6SFj72w3v1pOs8sLvV
9vaC4hhvmyPWegZmvcYHw1ytEdGD6YXcAZFogq3UDjtWSyJIRsUFsxW4zEF7mxou
tVoPBmi4J0PqfISWIQgChj7nC4ofeS6lxVw3uCCxUxWVG/qInX/jFFZEu3UZW2VU
nHdbcvp7/2vS76hSqao9B1jkRyb88/RYBFi7VR+L1y7NgVmHsfS3g1UqoUYl4UHG
3iWStCmvS7vOxY9POk0q0sqjw3FdFX1K958GzR1UgSQ1enD6wi+CeDOw/0Rr1xUm
569MJ728FUzC0zfKjgV3zmehiuTnZiSyTTcS2+8xVOk11+37mzeTGwamqsWMPA4Y
/swCrPvH7zyhrWym6JSa5ufEIEbJ2I/UfDSuW5ywqNmTgoCDZdIGeSB6Bq9ZZ2rI
4QTokgxJ0dY1VLHdwCbPFJKZ8PEOwi2ZAhcXjOJQop7f2LFfzhEcQVTluBN/yMlx
gob6ehOhqjdBwZNPp8Estr87qUYBKO0WXe4hEe2wQDyTwutXzjU2zZjDdR4Xkd3B
UYiZIdi6O8It7d8HmDeWYfOeX7UUJAdmNBKJK29dIVaDfdFJLCI50itKOFbvBp0t
fKNrqRaQaqBnZen/OyUo49fxJvu8UoyWyYDndhJAwG/TbncWBtcz7Hm+qW106hCr
XUGAR9P8kbgSNuuUQQin7oG1dfSLPQZMKUN/XqcTVstQIRKThxtV8YwR2wJJGvZb
YY7ZtiWaPnWs2mmmC0pxdI48uMuaBV7Nrd/a2f6twI4ISbYrS0V7gbtwh221TyEZ
U7YGWGvYDWnLNIA+NB12UxGMfiju9r7h1rpk35/QB+bZ8vuGhat4oihhAuneeQHO
IkPFJ9hbXnBJXw/gNOgtPurFSn8mwcyYSxTQOFdvQPb6686Id+x4t7ZN4HjXY33C
2/yAzHqWv32NLY+dsu7E/idqX6cBoZ/XQnsGtH8Ot/F2X0SBK1SXWarn2uOPax2v
sYl8AqqoLQa7lbwfxePFYuUfwtA5sYCA68twIyzIcKRZYZJu4pT16yy8WZJyXa6p
v37vJnqysv/CTgNIFDDuv/RlzV3KCYjio7DA39I/VUnReKi2XDFquUw32H9I10Fv
n0gz4E1jWly5zLCPDWZANjyOcJs6LbupncRLLRGhrisRRNszoDsZl4JRtHot8tof
qpjiYjXzrxlBPcDhfkInvdwOtA+zwFFxhl1NEFjZC42RcoBknXfzWlbpZj+HpWvY
idWX+6RqAT1QPzyoFqt7GfNTwwTlPZt9tGY3BAxVapeEEz90mgWk9rJpVb4uyrG7
Tzxypth5wkuO8yhYPgeC5rynLEUtww5FvhjwDLCDSwKMmWN9QZhjtcv0F2iLRLhl
nzt8Tt62BtF43YH7AtjBdvXY+qcZtwHkge2PAIWF1phY4GIMAAJEEsjcp2ekQSb3
7FO2Bxo5XLInq+6BKFs3U70GhHYE+TlpNSlKTOgT5QRszuCef6gvaFt80RBVWJlh
GBCruozF+pPoI754FDQTl1Jhatu9ZX+5t2UPR5zOKIjNfa3XHNofH4MqW0oVHCZR
LxhlXZMue/UEr1F9Q2l5BYAAjEeeQRmDKsFpXXzsrKfNC6K0dsGtG8pRZO96zsKk
7I0f46KhcnOoO/cf2wpMwQPan29y+uEcMK+uY4qpcpLGqq/GqINU4DKZLzcuyJTa
hYyhqSO6jXxQC6YPnevfpd7oe0p93H2fVAgmk6UGXcgxXQOpU46DhJAVJsIEY9uP
u7fW0/Dhwjk/ny93o41EFg2acwjPCClht3Q0UFtTbnxbEC2jcV/q5u2ixUHvLfNK
ATRS69RRSBV+/njeN6iUcgzKiWcvHuyamFU+xM21Z+k8vrcAdUZwWMt9pn+NQaN6
q9Y7NkljkstRGJTFLINQrqXpIHfVTSWxN2M+hQhmtM4K8KBTrHi3qaqtKLDATx+1
B5JYqGLreizvt1cB8oCSSUKfTjXo11mENoG641EEL3KVfqlhjalyE2PTgSr6TBgc
P1Aa3JMTfPhQXZDyTLHhNdpwaCXlb87wd8mIoIQGPPCjkMtrjKhZLqgZnl+mEGxA
Q//SUtiNmnUf/UJ3Bs+CYtVGeSMLREeIPpE/psTOO0SQ6oblBCLeoxVxbaHr0XDd
rqyzTJouROlnVJuHDLU+gV28l3BwUwlReiqf62e5lRGW99KsoCRv6zvB/gA3sKQe
nnenIOYO0dASdPM/WOs78bthVN++fmvu01zGA2YOeCEovL4J2hFD/el7CUxrBD/O
p4OpmjKS5Zt3t83QZm7fSOYHI7rgc8mOC8LeQ/2Io8tgTDd6yu8N7xX27jsKFzG8
Re80qrhPpjinofq4GuQ+urG3pRsxPSQMLnAVo/AZRPYq8Pqx/rTfVp+lFNrbbI0j
CU7lAdtdvUC5nsXp8K6c46hHOo5psihquC6PaN7L6w4VPCmnGIHpLidTTLeTBzAG
hq0Pb/twHWNDx/WpOU6b7az/yVXdz6hKU7Tvc0skyiO/hXiGxq0SMkYQizCFYNZE
UT1zT27l+82JmZqFiF9QvruLA2RfKIEnGkJR3bvW1FGv5Ew5vFx8erRuKA5pbbqA
r7HnCpGkev0O8BXM/bIeOydOKomYTpBxrtYW4wAF4ghjtrAxOmgNIuNS2mRPupL2
odgZDVbub4ZaHQ+rFU7NZsX7s7jSCif8655c9JLerNxD0oE/Kp3PHS79SIhBEJjA
R9w5X+McRHuSq/PM8kTC3S81kdp7svm91QaWBPVTi5Ig40IlWUbICstXImxMdawA
J1/ZZm4G6oMEqkwE4eYFf9qTlQAToChtnankRWxV6/QxhvaynwemcpXZmwtxtukg
+zNnzzRokuUcpSaNJFtBwYzE5sT++ksTs7dsFci6m1VOErNXVfveKHfejPRdbxJ8
8N2oL03X5vmMaoyYjqgnMXiNi/UayWIH+XBPYx8W+ufks+QYmGBJiCWQk50xuEuF
2rgDIXI+KineGooYaB1BK8ZtsA/uEnhkBsdJVYNd5jLYHcMOPv7JEtoHxOxGzvQ9
i8Q9xF0X1rrghp4d9YrvgfY6sDOf9CHf+1gkBvMtf8Pl1VWLD97UnU72wFhWnr/i
pGzopFzWbVfQdaOONMHKHAj3xAwhyMI2Kqa+Uo5naeKWz1zF4UuvpSihVbAD5w56
elZgOZIqyeop3Ml3FcWhaiOfyJQQZznZ5Mv4BDvx8MsKtb3osBH0OUfOzoetq5UG
sKd9/95uRo607aALfPxxuviKaUK0nyVA76FRbouNClwcOEN2TRrKYcHGDb2kGbBC
I126m26V4yYD+uWnK4WSYq6kAhed6yltC6fJprWPTfw0BjAdfDhXanXyTlH6c+lT
RC2TjPQQDj9iCVIXM5OpmLTh/Csv4m3usMfQF8WMKDdZYHvBEVDgOL1fkTc5lZ+N
cX0xntOxyK5KdoHoktZ/SEMAzzpEzNlV8Hs7tTxUY2Ws29mCnP2286Zl7ho6Xmin
xL7RQtrJym29e0nGtWI3Jmtrva1zoWli1fiGUK5qZg4jMx87dvgKTMLbSHEvx+um
R0J26L7FVev9et6tRnnsHjqL0kvSx2qBtH6UmbQPTkTfXHJXXDEJ6DKQOTGQ4xHa
y39ut1m7TLBOBxx9Yb4uQZny6TPveDi013yScq4aBF9vtFjj7oYFVI0Nxwlle8IB
EjIaN4j9G/U07cs0nHCSTxXGlOqpSA0q066WxaWXr5z2iop9lhqs4XtvM8h9HqHi
NssIy/y9HD0uOKPw5V2aUOpkwpKCmuRiYpxyA/QxM/x0XO88EZBzvrqIb4ZwmOtm
YKGHvxhybK8Fig1berEGeAxm4y+tsqUOxsOdpAfoeZmg3DI14P0D2A19DNATFRdj
6mqF/DOGNh/A7zy0aG+vr2mgxvBLmpM+nGxlcmygFl08uK5OwY7aD23QRZPskoNN
VWGNKRE0rF4Tj9HZzhFVkGblOX9ohwvVu+V812U4/y+N8tXOd218/vYu63sRZIDQ
X0yuhWJXOK4w7shycMGnf/zkiONWcwns7weVDD+jLeikG4wNChvkfOcNn2DyzKwW
FefJPkJbO5pXbWJsPbU2CAhccWW8wFtDzS5YL9WfH9laCJXEVs0wY0G8T0OPOsD4
sTMZSWVsqAxJ4EVby0xnh/Ir2nba/O4oeCh83g7VmIHX87LH+NH9tHk6UbOM1ZjQ
NZ13XqLs4/9w/LKBJnK+5LirLDecB7AccXvv57j9+FizxvbkOwoKKnYhqMgSHBUr
YC2dvvDoFe6NyEHxWrEcC6Fi69ucLsGm33SQMB1liVWziSsKA6Gre/dCQTGhwejO
Uts1hZu1GWrC1/N5xMmY60glFtrWMvKt1+u/5P5aCosiJV7RERuMc5bOh1XWoEHz
Bindn1DGjJ83/Bu9JXJ+VXerw+fuHqYGbWEPNL7Qh3R7oD2Y71cCGbrmMnYEnxcz
eoCp5pS749axsDRHd9Kfts4hA5yC/rvuiHyK3reY5/I8g0bney+3O979IRLJzCd2
1zm9EjJbpPE+XgKYWD80DZ68PMkEpy0o/mO5vTa/IyBwKC3U3AT7P/L341dLtARB
y/f/U+cTrLm/Mr5TnXm5hMFJBwq+LzOf17qcb8ug98dLxJCnWpixVLqHJ++u0yYF
dDOAv5bBbauNx/D9g7dmKDIYk8JZEpj5GzlX6wsrMh++KAIvupbAcBwVRVqjVz8N
RoJL8GWovBCjPBbj+PlUlfzUzjwMQcU0GBck9XOrrTZ6zoMUn/g93gd9Hh1d06w5
xVzud8/FAomwMrsYG+VBHGhwvlxVeLVFZmgk3DPMBJi9q5yfYXiiwSQ1CRfsR4nl
Jp0CoYtYZLHARLGIdupq0SXd6Y+bSWuXAJKksRAUME32xjWNoJQ7jYBfTj2EskdJ
YOfkIZBKkMDmM52WiBWmli95JU5qp1sOxGzXbrSS5TeVOw8GF0mhTIPooMEwbvvi
1wvdwJJahrFdWzmnOQCcEG9xMzXDY5e6KJ5ZmhwkzyoPJLcng94epCMKbQnQPn0F
W3g2POm1TREHlIYNLAK+EA2TjEGxOmtmSJsapCB/f/nN4RyOXi8F31BNOPsLBnE6
9tmI+d+nMB+x/xWxeDK/GJhNhzt1cShY+YVfsekAHFlD0jrCLeOfMkdnikAx/TLO
iByuXMRP0jql4y2VgN+4h7JwWfGmELMr75wGhriTihPKCrsANn9MKovjnc6Vsyx0
0m8DQp8cGCiDZsqkdZ7jlXVxzXuuR5/L8v5gzjcozqVWgotRxXOVAZyh3UGgNTUI
sEzpTBCwoOanGVNyCL+QwmMczXu+5dAUEDj03292SjURDK57hgJ9KmlRO9S219iJ
MKDZ++4xRAln/NrKSEU7PIyFTIkYQN1QDl5UKDyby+GZaY7x9/fOBb0aGdXthZ2j
1cHHZ11GYKgb2AD1shaGrwnY48AilpJTpeQui7K9ZotOl6v1l3Qp3YEk7djItQm7
DW/swZP1jjoU3OxaY+4qWEwr+t3JRKHvFdxqVmJE/v3q8J50TOMaWx5Y/jg9SFhl
mETYg7ggXYPEpKh4ETtiTOIcRk2W1bu9H02HSxEkFUC++vad/oNXUPvzfDQ1XQFy
2ZaMCdtLaILvTSs73aPhOMsmgeK1aHHcedJGAo2zE0uga5pJxPJi+xjjSuIlSGvu
9WVCHU5GSqQ0SsU+Qzoph1uzRmcNb+rcV4rz8G+5Q9h5zY11CKW6P2K/+XtxbkGg
Pqi7dpXS6pToLskTvQNRcOhrHbDt4nHR1gtofX8o7FyKQgyipOcn62YfBZhbHXht
gcAxt94NnpWxhvx/Eb/lupBOrO5Tw2VubhEBSA0JplwYOHyYAP5Zc2zI6Nsj3i70
KpOXPHH5/D+KKdABOHzoFyZnXYC8xI3tCjkVwDf/hxj/RcY5CqkMhjuXXOZUzCYA
zYOa6dUMGFaj0SY4S5nboTsL0o/3tr5k6eG6Dii++Q35gfcSawLZuk7Kq/jhv2cP
hXpAN90Bi31OGMS9FNGUpPZwsvI36ljYMhfR1aTB9sGpZAaMDb1kJ1Xge2SRzejm
Ze0TJxVzc/NLEIDzURfnrgYfCB4e857NlukdmTaKuUKtyGz64p7bk9kfMH6j6+/i
Gq/cGSeIYNI6Qjx3dBLwXWBIsNogvsgBwlUni5WX6F67xfvxQoOr71is7Zx50Axz
XYFeHbg5D2K3B3RjKZ+JsPTBcIfL10CnKPFtSS23jKWfMydgS0IDHnN0g7sdX1qW
pDh3NtJMSSxd05qVdftP76hgMX33LHXxWvaxBdrG7Dg0ZvnFwtBS04jzNOt3AqwP
znvGn6xgHAboBl2I4PduGx/m6tHaemwnZYZwI95EsZbRvZH+0D4eCF+klqSurk4h
C43PywroztmB1i0m0kXG/K/bq6xiDD3q5G0JHKKHd2cEZ58xf2bG4AzGQZV8t08g
e+skKGaDotY9e7XZyvDG89LVkyr079BX3K05SziiPc4rXy6OiBrKbWLc+Ri+xCoH
oysoDPLQPC5voH03iyf5f5WDUmAyVU0n9LWW7ySHu970DVnPoo84JrBIvekX/4yd
Ab9FsRbbrV+MvOIA4vchFj2zCbBrtYR0ZHvggE0OGlx+a5Ilaky7/LNhTwWiSBo5
0lFiFFk5UxxrmXeR12uwhh+76vb+PM0R8F3blEPTS+oLeir9P+GyLAek8SU9QRkM
QUrF9mtscfb8BPzAn1FwdcKZpslbsXDYcwh6FRlSisTpXvIynJ9TrkYsU7PK9RfB
H37b9IV2fnUtRkAplV2y4OL/x5+o0/1jsyE8E5htRv/PIGx2tGlphPzAOI0cNaJf
xMpAT4OJoVD/ALfBmjE/vPOe6NqRJvnIsA4CbRY9OQJ1YFUEaG+p7L18FLESfoUk
7SnK1MQHVBLt/gGY50iB8uGDDWDqmCldhFOJ+AUZsEBeeCoVcoMJf3NyQc+CvfbU
F1q3fZ3npLah6niN3bEJWxCG/OwbOdLjtPlZ4GGVJPSXf6ngTtT+OkiJxmvckRCF
3rrHYYoGayfTha8+wGFjMrqhSx9ZtFAsW1R5vccFUH9pA0AimQptG/rzrzCQ05tm
vPyqKlIe4Kl2PNIWGz7E6sYhbjB0qj3G2me+ZEfwFQ6KsR1BxZzxH7yPaBY/oW11
hKWQBGPEcw30gABFR6WEeaVYHpa8QNxu/OIwJlyXY2G4gzIkOsw8QQHah7tGYh5Z
W1bhe0yM2oUKSlbX0WzS5RM3yLNRdWAF1F1cN2Cu6Qtc80GitbXVOW9nmIEn5cum
/FSMUFLG4FIZ+a+IwGsNYXV1PQBuF5tGPxYGJQDDVMXrLriNNjdP56cQ4LZ/HpTY
/WlD/6P6KghFIEEag8ODTfQJbHYQQBjIxAf04payRJJAzTvYrAN3a/ou9/wagewJ
OF+gX9VbYVEviZClYm0d9tUtELYiJAWqMv7Q/9lti8BkAwkLRb8Vx/1ViCXsKdC2
3o5Q7soqLOBQ7+UHwci72eQX225GM6fdn4TwV6gRg294Sn5twBgdSz/Imyn4Sb9N
QIXoqAFM6q4oKJKlAuY2KPAW2Q7c+OTiVO8JRf37YRBQ0bNS8UnkGspalrcRA70u
DzFbLmqlOGiTR8vn6n5ZoNUBpnzhrsx7nXQLMtAHI2Z8047Ed5gTUAQrS7Fo1Aeb
uvYe+NeCwHCp6sQSz6LuN2wEqiWmhh3FZL01U8MuCIxZUiqzlKYYNU3BoSjTMcjq
rjEodpppo2yfu+yjE0vWXQ1PAXm933wnx0Tk0wWgCKhnT7ZeFeOY8nriFZTVkiF9
g7WArxDiqcaIYrs/ET29BUkQhCUEqRp7ux9nu7O/k0GUZCnbix7++iWRLZNxZOkg
qW3Y25qR0gLpAxBXs+LejMerlZyrtSQzZWDfELwXya44OuJrWuuHtcvfeAl836Y4
h+MLi95YS03rWI0T+D0fwx0Y+0cTtZp7Hmq1hpA2392/CNG+OYCYEgZy9WzbYtqC
DfX5rMB3NuSPOyxUNxwYGoKbBeRzwANHIFyGsclsl1xu4jr7KNH3wdCCYvznX3Dc
umpcm2HD2ljjHzrSYL+XqVN3FK8Gd8TtbLec4kSrP30F5Er1BE6Sz6ReT4FS9Yq6
/Gx7hzyoNvgra8US+0OiRq1cComh0PjrmvVY4w1uBdWybEsIBEtmC+GQosbhyCBk
z9jJJqPWGZl4HwWVzm4k1s92wLNrh8Zl7l2pCUsBRu0FHHEBE9exbkYeuhTqvQ4s
kUzb8Hg+8QHjCpd61QL4nMRVzewAVCgDAa8E9iVe2LK1WazwMV5bDIjR0SCOrpna
ovSy4m2D/pXFoqyqJGKuKT25VmBEk3ZuPf2VL/QAzNPkYTRN26mzPkUxPS4DZtWo
AbVE5M82EXIlRfwN05L3uluWdY4kzxOY8DfEx5jyxdJk59tp/Bor+PeKd3CRMKcO
VjoneYyq4IMLNZSxxuqA4LcZU3VwMzbCv93ATGIupdqTU+i/dByD1UWJHjjazszG
GkDnrvprGMXpiD7tCz4aD3ly4r1isUc6RkeqE8d533AINQzHjSgdtpw3ZKdaqrmT
mBZA3OLgZblAcvNufARDFXoOxT6tucUVo7Jvre6WJ0vzRhI7WTocwuJsvAOQke12
xukfyO2K0YicuoL2IvVeecaQEixjhCfw/O3wDbtXebfeFiBPTKNAjEvMxa5f9Jmm
texwFYJuKvtXcLIPoQur9V27OU8CiutTvACv67ei/tfAHOBm4RJ9/0kqJYuMoJcj
SqDhwGRT9etOQ/yYkumXkracmVYrE+x/h3pXHNdINdsUSjXhg/XRPV/9WyN5jvqL
rd+nD1oM9eGXyPyUBacWR1O7qNb/eZIwlaLyeQlNHFI0vLdkByv0Cf+0tFnnIAEh
HjO+3mjZMx0KMfN6UslSBJsk6C5QQRF04CyPAaitYLepFikBOsheWdgBLL6vLqFz
YZZTVbr8viL0UoFUzKBNzc0nf5Ngr77hlTGy67A9Mm4sDyiJsXnTnLLpjMjfoolb
DqIJk4epoFXHp3HM9rsP6Sbiir8SK68+6qYCwPn+lwGCOt5aU6ITqmYE7b7YIcmY
qv2H2X+4jiLg2F+c9ZzfuyFoYxCpN45wMyM278dgaOkqtQGjRX5fEFzmzvkSwei+
RDuzlNNUpNez882EZEvTheSE8H2CQVPGOIQCu91lLMLVJM8KKi8hYr5kiAVdihxH
gUsfQ6mHZNTprm3uAb8erQWFylwUgDTAi/YybSPmfADkHrptStcGzy5a1Z/jk3y4
Qn3yhwD3kSkL2k/Wr9QAkqbwDWkcDza0eu6leUr2uFRcwY8FuYYDI0n521P1Qj50
8ZJXKetY0FyJbgDborsBzMGJqvDaezF1WsBl2F1wBcaYwOTqfhherTVEWpCsT2WT
Pdj3C5z7PuPwMv/jtuEqkezrqyToY5hmLM/u3HHyjQfJC+cVPHIiLE5B3rcB3czi
WmsISrQ14lKU42bdWUsGtcBORGawE8m/Dp7I9CR6uB5rbZUTqqM+mr/puKGN2I0i
vKbIrfVwpMKF9bik24kOvFdXCIue5YB8YRAqKWYgcD2jImuJTKuIDbkhVSYOuy/O
0gYaX68NrxFVBYleF+E5RF7pV4Q+SSzd1ZSYbkMY26MVM4VZ2Tv1s0OehLFA05DF
taeHE//XPSJtde/SLuAsTFVAVkvo9l51DozaIFJtapEofesGb+M1kez5E69xKgGI
nv48nOojOCE8d/injQw2Z5JgKsrU7liSZEewX1csZGLJdc5Xk7y3KX7g29W+11dl
OwPDEefcHF/fa0OOvsyGsAkxeURr0CcTh6Qc7fH9qt8mAQhZvQHiGuYtdphxpE6H
00K5d2+dcory9nnRfFd22kYRA3SUiPs3QpTmc9Rz34nBJQi0h2FLFYou6Kr+f6cV
LNiYXDTfhC82RzDPe3c/+MeKZAus8lRILm2eKdC4rQeO6qwL53xzu8BpMGo8P8at
ke51H2JVDNpCmxiD/QePi0Cp44Xnrys4yQ/H7EHQJHHtMajsEv98PEQewqhAGRRV
fvHrMXRAqqloxeGuEHj8BAHtolcC+fvsBbdqn1JjUA/9JaIMwB6CJ5V8xhSyJh5v
8adY38c2MHjdhhMvxvYulK+YHVURZzUMJgyzFDnXySVs8xMaVsIgZDLEUlbj7p0p
SqZGaTA+O1U2RUUPsvyWCb8Ndgy7ISfAW85RB67xqATXX5OXF4PmOMeoKPLbWUIE
DzDCQF3j2TjSwYlMh6qC4RhnGfCyXqYbEnxtgh9vjL6cHNQggRTNM8kUBIHumuKx
Ev0CVzfzOauP3ZiiWngWdm0pTXi/S3Vl2ucVyvBwQSMac9sxgTYyIbl3k7aowLJE
zsGSJGcsp4NRAdGXZ2T4EmSIso4nKPzIBh1M1ws/NRqD4ZxHHW9xMsidpdeObfvJ
0UmKf9xPmhaAKs4M5waBJFFyVDbWtD5oDbrVA8rwfkXw2iFJpO53i+4C1DG6fgqD
lT0mPbP7u88G19H40usxoI5zTCJNTU7wuASI6OzY24ZKc+NAjckr3w/mBlTkde6j
XOH2nu6HnCbR4iaMm8jZ1fwe7c0lyO+zIf6zjs4Dta95r3j/AlBJzSW+P9nQ5YX9
KShDXqVuNPqWaufAfQAviN84GsPdm0Q93JuUgCpzF3JmKvPr1bzuKajyljktEp1z
qDVCNL9qAyxVssMKw/phmhosdClEA1/tvuZAH8pG9KvvSpQ8B/cQ9LNjeqZry6/o
ApZpj0hW93IXKUcC2tXN7pb2+ynucNhAk9hif4OaO7jPEzIht7XGtcFIsQ6Jtq1Y
XjYbODIH8QO0FhESYwB+gBFqEsmmngcLZLgxmTrD4PGjPOhrOZXfkvPeE9aRhLKL
siT7+wvBwXbgFx+pP7Ugzm5WNp+Sv76VVBAm6pgDrH2xXCkEVvQfmI1vJv/AK0zS
IjDpDLkQWizLYqpCfAIEaCvQpsSsW1xpVn2qRznv0W4M+iI5pVD8bkcA2acjb3z6
XkdcCkvSbYXm4Y2JA4etqEakogFfHbQe83b9aJfVUD0oifwO1iJZV8/4rCCE+THm
rGR4538uhrZ8HuQDskBFjcIxdNu5Oz/ilU9BHBwe4W2Sx04w4xDnF3V7bp0I/XOv
OvAvgLNKBmofqRm+VjcSHJvuN94rRBpmncZv32fvmQS/rNM/et5m5lxaaPxLn0e5
B93U8FCxilkoBot3p2l6bviG2s1zX8rIPIxp+Rw6lxhihWllzJk9Rn/niDkHRX/Z
AkYWSu4llgUApbeMS5R8Vk80PFsG4CbqT28HIzFj0j7VRRkjifu9qbbvFUq2hCzn
gcf+38K/dAuuRz/tkvkShhEJBQLQGauhdksO0GFDsHjIQaJcU3/Onbp/JeCEXXSW
rMGdmzBx1dn0t2LgCnynwYh8RmMzGe/1JU/3XNEJQqDz9ByJ1TM6EBgnDsG/FH4c
99W/iTSpOBsrOIda/ss2qgIkJpcxdBtN3pYyJHLHMmBFt2+aGoxZO2xsKD074m6v
eSyr6oljjXOYdpRQD9qjCI459I3dq6CTYXmJQDdY6rB8pIwrdwIEOD+FTRdJ4j/e
J6e7Idj5ljADrBMBIoFEbUhuZA4uZn4sRz5ceIpf7yT6DPNr5W10WvIFctJ2xgzj
ed0yGrjXWpctJpKFahKPEXrTcqlJpkrDhGe3s40hoL1s7ZG9keWoN1unr7jFAb2K
UfACNlU34l4V9IjvSPTnxaVr6amRtNRcb6OavdqBL8z+hEw/4bTuqDf2PdGHVIOc
gWVRqlrLlbYiEK0R47x1CJoPIa2Y+m/dz6ABrAOGUOzzU6IHY2eUPkhxKxg4/lCP
kLfcVfkjUSwGyCNxVCtUjZJskMh5Z1OpqmjT9qUGDcKVwqBrXuaHpf2+Nd6M+GDf
VO/LSmDxuXrIUrn/KY+8rHFdZjtRrre3J3YzLJtoEMEk4tn2YxOpPzGJy+DFHO7a
PVzm5PYLBuiYDade4n+d8t2eKBvSjfyhhTxiKmj4V6I7CHRlehXjrQJgaXOROCWE
9flVFNZAWuI+nhm0N69RkenYx1X1vEm3zaA7/ge/bwFkREzVKRwJr+/ZGbofS13J
aI/5BXrLHT0dvPgi046KaCc6hThSkk3HDP7lkvzxNsmu70G8jLOauKkAXiMvDtFK
8vPU3wgSkweQ1JO3JHXwycMs/XwaaSjowYNmykQEebXbKaXKaQeUmtQBiIkEjKw8
MQj3KzInUaYDC0vH+Cxo7hp8mcqylHaS1k2FtN2Zngu8dtrfyqv/QE75V32ptEti
oos/bnhcI9FTHknSTC9st7U26EewSiq0z2sOyX23953VJ25sqSg7E3c28OZcVRu+
n0a3Y9ff4PQ9AzUyNmmCF+dqW3ZuKPD/G7C1QCxkdshfTpl/JGd5vkRxtGEbkxmv
0IRyQKgYNzzOp0BGHnk1u3x4kpuj22EOJ6SFqePDbuvWNYqTmR6Nci1ALBInB1kP
Qj0Uiw58P7Az2Lf2sD+LP44TwaU/sZVChiahFCVtlH0XS+wjZ8zETMJ6pcxXNjmD
IsMrDitMLXK3pDLmal5ZsgR0qnjSJZk8vnUM0ufvzHN1lwYNqO0ab5AFmwMA3/28
EzRBdf0oiYE9vrGQ2PHRpphm2nbOG2CKGGTIsD8i4kaGe9v/8dyUF+rtiz6u5wQm
qqV6tC8pD375kiygXrPjzAnzEpb7xHl8/Kszv69eYHoK7L2usjrfrOiIpR8V/VMm
43pmCqEGwRm8qTynxi/W9nDAfxPuEcEolBz8/iEDQrD7DsRKpyCMbIDtvHTi33Lq
iL0ggJG+jIT2OgJxbgo9rgD7j46/rG1b2xhst4SxYbn62MHq4y9Qani5Xd8mshD1
yyAQLHlnjuxHxFX7KggRT16AxnqwWjqZIZ0JPsSs6c3kZF+8Rbu3X+3vPtWDaodu
KG1c7iAG5EBLDT77SygLv0f6uWY0rAIGnCuHDC9jMorEr2n2S+izJBODBqRwNF6O
eC0s32giV7NMS/Qsy9YMw5FmN6bXst2+QG0GXdDrvIHHVMSvdwqeFLggbJEfDZLL
SAyn/5f6xDL6/DtQiJ9dTTS0PnFw6oTE03DFKKw8RzAUNTbWArpeQjJASrCzIzyc
/yPqG9GHPvVEru9DDae3JrPZ3/UDQjfiEN4+ALzb4FGZuxF4IJIIEgQv+BYSUo6A
pN9UcqGrFQFzHtq3hxSep4IBn5vn55pCCHt6dEWm8CD3Hv7ggPXECGd6TB+AStOu
gcuf89XoHpatV1TwttcFMYnHcgaNliMOsBsqVI1QSncEVkaxj81SgYYa19VK9Bqf
etDPomLf2BzaLnIPNBNhHdj+TQxF25C3FrJz1QRsJ8cw4Btv6bfZ7oq98Pd9TILs
HeXaf/6G6bT2Lo3q7Zm6CoGDonYT5nwpiNG3lOyLZq72YPxkW6Ixkzgqx7WVwIOZ
IUoDYicIJbtCvCLwHejJ65pSslsev69fu0ndHWsDI1L+40RQQmLsbXb7+lW9sHSj
/zu/S6YZQ5a4gAmui+9VuLsLB5oU6dHQTvlhC5AdzM8NtPrGTvf68L2LYq/K3GKi
Oos7nno40ntiy2/d6qgRYvIguOf4Xf96ySro9eISQpdL1GXlsP6D8CvM9lkYkoBC
znn/Ww9jDs40Ov6woS6WtRQRnAcVuvSMF7DneE9TdJFqW2AuAm2yW7jZVEsuUWad
lglPsz4XInzOWpq1xdnlw4Ssi0TdMkODwOEpr4iFhHJHhpL3XdDdOJEQQsFzr5dm
3H1letQpftivkkUr59R4AuHddJoXvscFOr+F+MRYDzByiZ8GrghgyPt2WPrJh/+0
1dPeI7i+O/OL7YNRXgOzcU3rCbo61eHcabb5pSmXkwxYcnU7VfNa5WZVkxcxZOej
whULXdqwA6g6v/j3OxHTwExi/ZJS7aioG9nkdVsd76icaRlRDP//xneEXKCMpEJP
H/ObkJRPtJPA2ZGt+GZ8RfvTF9DLzQX6m9J+xmYgwBUkeC3x2XDEE5u+jCVwKGfe
D9rQefQUtsptefiCAMt3zpbu+BY5+JS1HdNNjOT1bev6uAKxEt2z4bYTTUg38L9l
iclNF9wosBJpwM0zUGeu5QunHCr6RspRlivTgda+VgnqWfZLnYTQZAppJrDMVKX5
dpxNM0JM+qWmhbCYARcztyEzFfz87+8iSVFHVrVPIjfbzbcp+Unqzsc5+sim57Dj
8fKKeYye+025i42pUWSJJWm3e/4RJw/9dgCY4G2TOp9zk5oGCl8BVgK0xUdDSlwr
HQ6hdBjqRYjS8xSfZd/USbgg5hq8txI1hoQSTvoB6112NSTHUPtKrZ72JefCj84x
tDRK20D7N0i6QZfAWAGjb6EQ0nNR9of0SsC5X5tKObopwv9G1MY4EXtwoMWvPyfE
678/1UQnX2xhSzTDy+FW/xPEgPTlSkD6GDDyehVnTFyRCA3N+44fZ4hd9eQSvr4b
PHzi60woYl43MoUR6M980CoISPP00oZyl1UeT2s9SfTJKU8OBv45koMPiL4hGMG2
zEHo1NjV+CjLy70VYZrANEr6kAqPG5jO/VoNDLNh8ysDorEAI1sYPDjXMShKc/2k
nCWzWN/KJg0QCuUTpT9CWBeJIBSt5hr4xZnrSjL5A4fDzoOHnp9UGPdvB3+jHVFJ
bHHMun6pWSRACuZU7LRsbxdiBRFSS65DiU4VSAQttW7uWe6Rdw9B/QTsKtafyFtl
rnloSa8iyd6ZsWYL9Bmv1Y9KeAcA+R1j8T9xwUEuHfblHNxgBhRyXBVFsU+RorNS
npwZiDXyA36+SefhsihFmWysQkNkSOuwVf0kYRuXAcNEruCqFoMn6BnzPYf+NCGG
2QU1OZHGm915RRWLCY0poRXkCQogyYItH3Jf5/wmga/MviJDKzowc88mdrJFCK6/
X/cnKmPoM15zsVqv44hMdN0UZ4R0mkoeRBiwrFBa5yqxaoGmL3rl0AbwbtE2Jtpo
2LyUoBL7Jup5Fa9Ofhzq9yoJF633FR1ajHWi+TDfO+Qy6w7CjU9XVyk5reYunNLY
MsnAU/sGQH1jHzn/1kginzbC+VTko0cOTrn4YJtM5O1p9qZpFmWQzz8PuxWHqwmY
27Gmc6jbfagdq4zeKrq3uqwhmbRtjMMx2EwtQgtFJ+8+EAbfL+s0/Nfwv+iM+Yak
2QdAu36FJ5XhOwgyPHiM+NqXcPDz917EGKVD/qA1jq27e4gKUTt6IaXvkroeMoQ2
HcC0+sajOQUFVaLpUoJ8mr6uFlPiqUQ0ka69lyRn6vGZF7JzXCMrek//wMWipn15
6etNAma8W+ieHCfBI0w4BZGiS8CwYGVivkZVBjCDR5jLAFvXBwkt6Yr3C41SLS6k
fqnJGGABhjsSFWt4f4kf+6wqd1eUGe1yKCl0orpl10S8uAmYKTuFNDYeNP8hvXzb
Mq8suS/5MazsDDzjOouYM3sdEFtyTHHp9x573xLNsmAKxGbJOuK/jF78zf8sH8mL
elA+CxNZjf5N6UlSDwINK7AlmGYCkgk2LNe+SGRU1tOlVEgFN2kOvbN5jUAUHd3v
B3Fsifj4XBqtYUmu29dxThnc7vdx7qzN2msLMBNo91eABGWh22EWuMmwZn3HWkFX
z2zlCIiBQpBcQ5IHfFZBDITsDbT3myC9JDDD0NBMZETsHUNIRjQyHHYUrn58+yGR
UNclKb47n5G4rCm5puJ8q6fRbXxE/n3Nq+lpSAdXRD3MQohpWIatPNF1gl36B3Yd
SQN3iO0quI7pG4NPIMYpmxQIgEvxW+gGcBic58TwNXBH7oIR/UmCB/Q4keWABvXy
ITt2hiE3BlgepJg2vK3KH59ZEglpMXWH8XcRIQe2OTBpRJa1Pq+ppf0gYWBI/Dbc
3bTEvEon1RYAjTi9i89wNZ7STc9l4AqVQ6W50U3p2UnnYKG3JIXwl24a67XJL4kP
0WiLMDv9xLgQeXstp1JxkKsI8FT4mkOt5+A65j2KXUkFZL9A6qGCnrWr3lOEfaZY
R8XXCCQ3+WqMeOKhzjLV1fQ5ffwOwCSOnOjr/fFlHaEq19cvIUtbh5Ga4m2MbZyw
ybfwQnDY5dG/07mT70tNQ2Ef6KYpje2DAxN73J5v3fIdjLmRjDbn7Oc408lavW4Y
VpkIahaNakvrjzYEkVX13RT4AGCnJmfloMO0xUcI7YLWINZxMXlgiRlc4iBGij8L
0rnxNcRevjD5VWA03FXXt5hvYOrbuXC3quP59WY4HBE/8r5+uiFvesu1ujWTVM2m
kAluXyPkZREeALoXR8tbCIL72UikrKy1a9sMwGaL82CqiXHiM8kG/mXQkc8Qy7sE
YDzvFZQGkUdGsR/WHj0K1h4br6JF3D6f1doIubSEU1b47sWkIFmIyTxsUkpJQUJS
jaBtEVqMjOSy5S9mYpXK8SwgzxlXEDBPflzwyTaLoukQmHd/8Eet4sN4alYwWYy4
rvw43F7+wXXXymB+NQrdwPKQZu1G9iH7+wDbrFAu5Xwu1Zr5MZoPT11/Ko4BDDaL
g2P9ZSgj6cucRilsXUOwdKpM/7h/SJ24DVXgkzpiFlBkA8OeRAOKu2ZrhMnpVgFt
sQj9hqekyvjGqthMUyPMS+SPvofMHzTqwO8SwzWRSgiO1ZV3JLr9hl/SmTrW/IRg
B7B4fHV3gsVeICLSp8WNo77Fa5fRp9G+RCKuej4utiOWU+RYmf7kqfrdT9EUwvK5
N4uGk9liLf2j9lXfQXFalbpZCm1MmrHzT12wO3YKTdwZjh3EXMn4Zls8HdU7Vki1
TTQHyM9CQL1Z8NSJ3I8MZrqJFTqmU+cvhw02IcWlbid2Kg8P/Tc95XBXPyfzzJSJ
DusCLRdUzIxd3GyritYCmwrEhgN4zCMBqTObT/B7Rrl7Cp36Buv1aj1WhHOk7w9M
CGXYJOx1y0eCyPn6/edG9stO+BU7p/fPbR6W7zQtBZKwyVBBLddydVDDWjibReM7
wGhysFgUyOxH/9IVksfu48ecASN1u8AWZuFf07Q72N9t+/7Uv4olcg+Eb7A8juGM
4nzXTZuTcYg/i4xuAP3Li2pz9NSNMSL5WdRqsWell69nXJVAdL5rTqYuCpQVAXnq
B0ZhWeDlNA/6RU+eax6mA/VH85Pob1t/Cqo6mnD1lAnBTHcCZStx3HvyZoRzrZc8
X4DITJ4ULfZs7qJzSpbqAA8pmPJgjbc48DIrk2MaSZnVbdMEIgLQsJRd6Xz1Os6G
4MlcHgvrqnYj/RsEp4DeYZ48HHt6r0a/cqPLaU36okzWFmtibg+iu3Tj9bPtHRfP
mh7u9pK/kas1Lw1MBP7wz9SS85pFkMh3VU7m/hglWbEriT1+NRXGEEJeSusKJjP6
mj5RzVTWbEL/4eaA6yOv8t1A4trr1BJWnclztTcOWDyAo4ljF0cdHql9LwDXuClX
VSZO5oBdtMrMMel8TBOWLgRL3C2ngpLCKkY0zW6+EE+OXaYs3tulj6Gk7Ku1P7et
sg4tPbqDP0P107Cjhoa19q8AvteevatHsTkt/HPQfaMIkv5CR+ma6ptG/gNayclp
HOza+NwZSWLPT//xZ222DCCK5edc0T2CR1o9ydRh0iUro2OrWNiVljpHdveiWYOg
opOyqSQZFgte5iajIbYaGQoWyQcLp/Dm4Q74RLRXzkN9SHRu4pIKm+ONN92Yvq1m
OaBvbcthmVU+oJcjIhvipfGhagU1apCSVPnadcJglb/VlH9Ib/JnoErrXB/v9fly
Bl8/iT+hW+x3Gx4RQbhxQpsRDIUB5UmRhfGc2hJZfd2ZYdt1JUi+wvknDjSz1+SA
iiV1i/LNIlFSFakknLKqQX2qLyR6UsvBu35hTg8H1512+fzm19W1lld9tvCc53wb
tvQd4kh4kTeKzx0jq2S/nXdlXjDK5aSfBzYm0Xgfr4ylBhMqzln5b+NdG+CPkgH1
EgukW7Q2xp04XQ8Oq9/Qj8ZZozfx12HnHqrOYejuWq+YnVY4iIBQngQDsDh3hUhF
4W/tZxng4iu0i1vzkU3ayjWVP4goVJSt2CUYgWa5Hb5SqYn2bkkGA15ghgrYFRQj
PmJ/hJDqPC5dRo6AZjphymdTinuMnfx0ZINAflUnG0KAGOPkKnb60wiZSFeai9Ks
ZR6V66mjPVF1nsxV9s7v1X7dm68DXJLRq2nGqm47iSr5hHUKhz7p3715etja2vFq
j59VpfZ9BUyYCNL1qHEEV0YBRziS+jAVohYMg37Q1TapXjD4GfJBsnqBxHpFx2sp
mQerDNyx8fRGGpKZUDaKvTHH+ZF+hGAikyS68uuMo+hXxoDuVselJrECQsbvFdB/
ZrzA0oOWx8CF884WVPI6zvfFc5LyeL1GOhg/lVG/ty9WbQ9v+JqbWCJiBTzs48/E
xGN11G1CrSGDa5A4d/n2/KkEj6mU829a6TZ/fhGKoljpDU2+xMb7pculB3aQPQmD
bXl5euTaMHDcLNRmPAR8+uZPwmq5RulzGkBekvlLqevbD0luanrMOzca31qFzPm4
3Q/eDuRWYjOShg/cOOEdX7pw6WmzqhpWeghCOZprkortR59AHDucf66RfDdcjKIw
Zaz2gCzygOmFibYxtr5pDvcd9BYzzyuqPk62jU6EuCCmkpJ9wYawOKrb12x7Kd05
zYQO6GzdKC9mtZlSZq53vh9B/fhPQNmCvDYneKhmkqO3uHmiVc8OEvXyNYJJ+iCd
RUYnoFi5DW1ogITq8mvn5/7o5bBOpVbwO8sqJPcvckb6dObywTjv94GwXIJYawGS
dAz/CvBPvZyxttkMElx5pMfhmbFgGP/A0COAjxjf0QiNtMOYzd5ZsMrxnNfaJqIa
DgHD+LigdBx+H1FOhFhvunSSUtAIAhEHwoFIjb9wWJrq8mz9Zguxgwh+yUeUqwHJ
B/OZbxKKuLVJDiq3upSUpSExr0qP8K2JBSxgi/byw7TL4LhDC+6N9o/hqHvqrEFQ
FJ7/BBDjou0PThlCP4YR2+a0M0Vddi3kipekK0DY1A75PSoExRx5iaplZJESUV2m
PPklDE4QGbkH6vjA1C5OgP2pSiJjP3y8uN/G3Xw2NSbOve6Gi0CJAguYAIQuFm/Z
ju0b4hy/5jL1Bc4YRVzAJwagMMtKzgMmsfVoi9tiCZdlHegbIQI5bqESZsX0jEw5
Kx5P+fYxZ8Ue33YdqV3iW5hai6HgDGbcLOjqzHvq/wBT/8Efkc5rDCm7CrpWaPHx
YCG1WBIXq/dfg8o0kwdm6zztf3IgBtG+AWlE8etwg0jeNSLD4A1Zfx1gsBjZWed7
m5g3GPbTb9uHLMFc68bHDpIKaQJwFQaRpJuhoPwzX5gf/1pKlIx4RiqblJwTENX5
eBIZRhQpAueJOCJRgYYFmMcUDvVBR8Txy11kxNvfhvin9HqcDW02kVJkqD4Odx9x
DJNphFP9O3VZ86erurYALbTdDDldi3jSdH2HIOxUB6z4gWcaSJpOk5sdvLyoteOe
Ufw+TCg9arHqIydQ4ISUxdaGvRilxtGD4EQZUhEPspuVfNZ2hj12OCPrg0sXInnm
fd2q/8kb9hNWgxQoVBJBN56+4iWqhneUVesYLkAV4f/J3SkGmZ8Wu1TffqX0oszV
kF5It1ESTHfrMfJS7kEup6Q36oVTG8KhuX3ZZiC/tCVV/poir4R4g46q36pN8JhS
YzySgluJ87sJG4p/iKxS6BqA5CtGAOWN6RrNQ322vv2JkbGreedLLiW8MABlzjLf
1b+NgwansWDBC5H3w4A1aYENvvfQ9M0fZakxVVC5FOOFX7r+yhRwlsajZesHiFYF
ctnSIYv/OYWLckUf8GLvmyzb5iv+8bq7ylwBo6Ti+8b7EdaIZWgUCoEatuqGk3/d
Y9nkHJl4tOAX7O3QD9J/mJ6NwGsOJnWhfL76xEbCpwhZ7X+yJE0X0m2BbL88emVl
l0WVeBr0/nsBzTY2zsijSHFSWg8XSuuZm1fzlwlBqenSJBEoTEtQTL/AivLUXbHe
a9qtkr+y7wUT8Pi8ZkBwrmdfhoLGMKCuujYF52ap/uXo67V8BIJXoTF3+/Mm0ewp
b18cgHU1lzMUdf04poPLWcte+ftgU/UYjZ/oKYnaZLCUVOOENlLBAM4zjpFfvORj
OI6ndcvDwiNMastroJwCubC6bmcUs79I3Kqwiritofae+05YMqk2KwV4lC73QM+g
hIOEp72dRbmUbvmv0bA4Blaj4ID28K8QTwwiyCsUHWIZJgoM1nGBCfzk5AXLubIR
bogiwBtgYp9Onkqmkj0SVUWq3n3L0TBqcQ/AGRG7zpsW7hahG5uWt0fZZVLXeX5/
EQpGMtNhr0LzZ6bw025+sBWtHWcACEtXgMztCG1GNJYE3t1w6nzJgYf/9O6hYoNx
qDnUaAmCOyo31kisxHc31PV6S7d022VTUPksaKMk1aI8y+m2SvREDf2gqJPXR3rE
scucUXS0ESD8g3VZhLhtXStUltdibAtBZW6mc/XownsQJqnCLOYSiv1YaUkgT2K4
eb9K+aXLUE3MfushfQmIbf4otbhMPGAEQb9LyL7R986JkfXTEfqFjM1ISHjy9nRE
9xiTBangHimdTzOTyeGqZqQc1fRVFZU6jCZT5Y8RieniNH0TcPLINv9RxiPxPYIZ
gc86PZNXJYjoWn7xWlJiS9MxY/QWRwHyrkJG3ut2k2935oWRrs8JU5rifR5zFIxb
d9LJy0bM1Gp2zd1XSrtzONmqzHczCuH9I/lcK3RxkZ235Lp9X1YujNWXCFot8zdn
zyPfQxog9l7h6fnAIe+VgRwDCok4tnbN4WEREXSBBJx6wE8wGDAGlnfS5ny2Wael
a36pAlR4p6cwJ0LLN2Or1klZSE0KZiAyerKX6evS3WV94o8wBD/sEsILDk5RPm8Z
RGWZZu8KncAKFY1JPzdNNFTnBN85TL45kwPXkPCsDgzIn8vYqL3kGLDCnW15vhTM
u56OT/QOAf8mwBaeXGFYhv19pGWKkv+YCBSDaX0ZB+B7oIG+0L0Ei0LNyb5onu7D
zd10ZNSg4M0/y5VvAl0cOXKyKIP3D9E89odAOSAaUivr1TsUlQE3gITnnuJEEcxZ
idrgXYhgwGUljSrq1aF9Sj3A2rhUml1i8jL5lmnXde7LWNHH2KJP75hf794B9BYw
i9dKuBU94FY9JXPFpvEpwBu9I3RfOkavjtZRJEulkuS8/I0PR9RjplgZC8Bu7tf2
l1zcl+eDd2HjLkNSIEXryob91I2PNV0Uj83lUu9lsSX7adf9yUJOmig8gO/zs/Vs
udLBBhNRXfE1G+sfh25ZKvUzezwimZndxLQWd4PmNH4Shyn0ZkXrpwLvVNvbXPWv
KjvKw506GnsEjn08REqVwkefzE1u05UJdc/ko/WMFKnDEFEmbm7VhYDNcMIDlDtn
OyoksuZWWLegtD3LNJIpR6e1W96XoJgG4hiEOXL+eHocMrIWKH3DB9IztsYpvq25
2bsWjuQ1hz1ubXjaXIjTsCQn73rZpLzolQCgFoiihbM+Dqi1a80flyhfhKo+6DtX
tTQ15iISvbi0Oje1jNh2/N+EUeEfTDOBbPUOPGwxM1zm3qu2I0T4cEbaURSxLj7L
Q84AivlRFJqQQMDcV5VAlrD/0Zh5GJpqGMQrMuetvzU5+PV89PTBRzNqRSg9jbqE
MVmqAkSCnvjRLW/ybLP994mi8A9jZQHprEsDTKBLQh9TKiJqzSKvQO9dBicvgRdz
gawdDgkSNZeoRxKlUj0QVKrGNwzmvzHxNPc+ZAy7NUmVc8AIvUZGFCP+MA1UqsKS
jm9tDfNAtI7zANjg3YlssV/ppjoSh+PzEnluADzILNZDhGQWYrPa4D3lkfr8aHbR
Ks/em2ZejBz2+08LnDlUWs/n6TQllqPW9FzNfPd7dq3Fpq9BUhfAE66fakmQAo97
53FmtfE8Q0vsA8USUVKCGZYbiQ1GLBo4GDldn99w4dMRNCJ8tzz37cD7aBGOPfmK
cE3JM2u8qpHs9Poo6+VNtwm7F2H9gotgqmkUHrrGpGrryGl3EgJQaZr2ghaW3Hg4
d1nab/Dywa+N/xCoPGX0+BjHbQAO9r0C2YjOUEtIxzQCCRSNqsPXfk5lAHRx6pzf
zbgTNp/9OLWDkk3rbG0WfrbHj8Pl6VD1hBEpDKGUPe7l+2k1JyS42K6E2zyKca2k
s6oseVC9zCac88zru1QQ2xwmhxcylWma/s/Xqw+GCYeM+9o+uX4JEfUYwashcA8x
rMz+lRBhfYjo05x4F9Ai3sX4Q8rsCFnV3dS2FrfVK+Qytc/On3MYsJlXSioxqUgE
t/IlR/0LeCXOJ5de5QECOdltvs8mLaHSC2bMFpwK5LOSmZI/l17voZSxwPWHgQnS
XZrYRxMHQbsxbA6n9HPNqHjnNGiLB+mNTCdA3B+zo2H+H41TofTiaSAiWN/ZfmjV
+uVKbKEHt/+yzntt+r0G2dadmglexPjndxpmECZHA/A89b5Kvecnr3+oX6KQaEBr
q/4KZcvV0EZfZPG0xw+HJAYVe/0dtJ3RsYFWUfp1Dji9h9CqwUrXJJPVmTVCi9S0
TDbxNUYdcVWs/xcSOeXMuwzcGTIpdCJMhxD7PSonti/xH1ACFaRnzxLy1cD0U2Rz
uMr5MIGVeTEhlhwqEPSuP0T6t7a/Uf19Mwo2CdVKtJujKoolxr+C7MFGbRpKcmJL
Av3J5hzGSqF/Rvkn/XAjq7IQn2L5ekkQhWNY0inwDmTSPkjKFOmkG98HDEbd0c2J
EoMoh7bS00NrwHZikTnsR1HiNheWEP/hzhBmaF7zEc1tvUsay1iowMsPCF7czKv9
UlZPdFtBL4/UCQZOettz2VBEDWtWl9cb7pWg+SQo8bF9CTXCEciT/oGzt2tDp2YH
yw5WN/71SXQ1EqmyeHSEBZLlMks6FGQXEs9jeo/SgOmP4MnqdkTonFnRtx21138V
fwgp8rBI9cXF42xrerz/2Tvd/TaPJdEccXKo3scg/NaaVZzLgk7ZVYGcxMLq2tab
PII8tRzpBiLiRgM6kg0XaF1PK8Xx/SyPuu0cPxjnuju12X9xSUxgktCyfGpnVdbt
4QdId8EF8aSvyyw6bUT6OdVKX0jGQDDSv0brDYeYe5FNRTuIhQSPr5UuuP1LUYd2
8XqPIUvx7rVum5WexSS5lgFGR7DZYx82TpdtkhFUKoI7dyl9nl/RbCB72eDZu8VW
6E8d2uQFPAp6P9S8Ub3n/Lwg9KuYWakutFgVE9YNTp6f7cpcmrx3dWd8rkZdUkjq
ot3HYrq0lqDcemIErOA8Ych75KMCx8oNYfqtREJFlN+HqrxF+OzzU0DVmTJOPsmq
rBFN4XCMtzZjywE/fY5ONRwppj4X9tyVpLCiNDAT6lGRO0t8KVawR5iELD7Bhuwn
/mMlHarKypnGcIGJ9h86a0m70x5y2l3YEK6Sr9fR1RfsTNw0xhTqR0kSBFEcsBrK
tFIa5jqcVSXRCro12XjKQ+eL3SwTndobn8YIU2FzQB9Dz907loUeaSnVnszXHU8J
qkSSag/QHJRXPjArDS3fKjYSGhxFlBt1droSiU67DG+xpyVgBsam89al7tiodCsd
xoRESVc+Pvb7v2LfnBsFNVN4b3BnTVRFW0K5ywmSAMuxWunk8yJVIK+4LgYxxfTZ
aaeplAzJi4A7krsXfylIgAci5um4atawPFQ9chYL5lkW1wIdw1HSGZXWlEpOCgmd
xh6j4Am5PjSVYSFR14JtpDiEke/8X4D4trk5vZnAmZeuK9nc03WVf53R2/kTfRfK
zqAqQisHfn/rrnx+negAczc4WaCV7SpnyxU8GsP7reKOVrjksT999YOMqNklzh9U
vN74Cn3x/hwWkrZHha4cNMuNY0XjAG2zcGk2YJLe0fA642A/qNGN0WatfqYpg9TQ
A1W/GSheDgDR5PhqDHOD4K1/XdRqbi70RVO0YuHmLrbw9d0EMa173aUomlXAwc7Z
1MPYwpYK2/MmW1Fq8BKtMCapcHgNLU+4ohGsX1Owv8bbarBfgjaLxpkbqkIFtuyj
R6HV3I4ZqsPKcwuXnffYEDcuKs/6Zm9dSa3ZA+K/aVtgE0B+TAHRc/Bmz/W+pwTN
UaB99GXOJTnwHIQCVI6/5c7TPI/MaOomXc5/5dq9w+ihXzZ17x4c3/Iv7g8y83Rg
OPMWudGFvM5phbGSpKycIyRtnXP8edJe9EgiP3WdioNW+PwC0SNFGDRGV0muqimn
mPPkqG/CMov9kMslRelwq2EY/2VAukxZDahgwU7HvgPfCgiI9QFurxShllHpJ8RX
ulIXEeVhuzkd62luUZvWJJ2kl2uzi9YwecKCN+vnLxbQKt1q+zXGq5IoH6IfGplC
1BdiQ9l+qdhyQWab4ZDMUx1aN36+UPNRfJWfaziJVvsqZcRVle1BrNtBEnmP0kJT
a55lffjFNHjyu1msFKE1XngBwBtvsP8ShyDSXX5mOW8tnwx7cMQS9keInSl/1txV
+kyptmnF/DsV7cbGSRszSHjpl5PPT8BjhfYnUkK2p7XXLJiatC5Z5hFci71OycEB
ObEfOtL7TXxyFfvc3K26PeI0PwjoNp8ZVt3el9bGhZhwlQirOUmhIUDs181SmX4V
LOhqn+o4eTJQGw+HcNF04eEg6IGGCtlmZ5gn+BC9xqknDGDgMbd2ZzJsH7BllqtQ
Uf12qxDX79XgwFxsmCPY3+nmD/jWdC2Py4ulE8SJqnKZAKCzgHi3KI1lXTsF/r95
VSNEo1JumUYA760RDYnEfZx1ygSIfVuxIT5WRVIM/1MDQEj+EvTnPZ7yqF6u6lxm
CwlBol0bm4+674kdRLREohvbtADsnRizc4/fjFrk23ten9gyGcQXnYjw7uHwKTEY
3On+S0kex4S5yM0X0i6eeawW9apqD6iXB2hOQtYdkKxFdprrH9++RdlA4Nd7GO3v
iiB+v81fcpoT2ziNeU+jjHnVZmtjhpI5Jga0PLdoX61pYrUoGt9TBuU3+jirP6qy
X69ghHGHzNMsuRux5xO8Zi1l0jIZBOsLciMYQOMHC+LSGQyyDUzrGhFnyhbQqebg
EkDA8YtTJt+Rehjx8dHXuZ+PaAKTyW46KMAq2kgCkpdmt3CIQRVG8O5XRNI03d3h
xrLZG0II85zEuTErNdWCYekUi5R8yLQkh2zB8P6vvuXXIZfmIEmn+Z7cGl+Qok8p
ptiKlOtty2evVJs66aenvV8rUZuTL/jF/kyY8JsV02Ymu8zWxMhfb4ti1M2+o5R7
LxSQCOwW9HoM7JqWlviele3PWLZAOTakgeREJlsI5a6YzH1YkVhjCsw0Eb1sC3ad
itiTQwcFaq2Lk4tDKfhoYzdeyPXXeENOQLNvtBJ+iF4dehSfulXwR3gA7oNz50zX
AbIi+yf+R6CJucsY6MsbupxZAy89ei3ufSLtkkZLyh/k2rFT3Uy+nFgoIjvo9JUq
8KX3IjGbVcRy0Sim0UBWUCETkUqjMQz+FOGUoJKceyO4E3ZTIeJsvjcWawYeDaes
y4PG+zmLOcqjg/UDW3zzZc+WxvvI14xIkNMBQ29G+FZZ/CpZdSmYvzQqrIhrdx5D
WLkPNIC6QsnlKWbGKKmi2DqEik/d9O5ERl/OB9Ty1ZFLHeyxyYZyG4Md0zpE7uF9
3W3h62qTcAgkWJTNyb1hDV9MJbqWwA2/v6W0qwdG2vsFJQ+ne9z9+67aDYih68VD
DF8bZZl9jQCEBg2tI0HPOzQZ4+EWpSp3j3VJEM9IYyrUZrzaiN59zUlSWKOo9dix
O4RXUGtZ7BJacBOX82J9mdfoEVtpHBaxByh8ZXb18URsjLgNEY2hGIc3AdoWYsFJ
/vICF+8MttmfuNw9pZki6/ZKnPiVdcjXcHPPYr+ZDTcQ9SnAaHdQHvoDmLehs7qZ
vKQGh78AuYG6mEwg7ROIqQm94fbjAp5eaSm5IMlAiAcDDCyRmc1bMHQIGmtOTkIY
rc9a9QDHU1t2T7FwuhUS3fZfyFwh3tb6QM2gII7tQjeIOadhczVqJbUinaOFoy3r
zlMO4BZcTFo2MnN7ApuFYpGUskje3v5I7Ru6OPrZEexGRAj2VrgdtS/qeseqvvOR
c+lS8JlPt073vDT/G5VmzebgUiIEBjkJFNlRGBRuEdhT+AfG7ELDwJCvohUW5nlS
/+crnt7jD9gViuOMcVZJYzStwzGNhg7qub71HbMJqVLJJn8kVWGUrTsl1Aq0bUg/
Uaqw0KQB1P2OCuz4TGWRP8xEw16WEgL34Hgrmnj69ak5Mcnz3wDnhQV9kfRmwZ4R
AFdglTMVBOFIm6eflhsaIyvMbrRXTzwvRSBB8St85qU5EIEu1HY5oba7hUq9m9gm
4FzMxFfIcIbtme85hH7bwZnxwWELZ4XHp/fqYsPHVPDGRXcCPz9s51+9m7aCR890
eYQ+YeZ2ds2KjBlLWmW+y9813/bhvxnuQRBsABE+2deEB5DfCcDWkzY+lhayYM6b
KTgPzGeY+4tN/uVEN+Oy5H8Gq3rN9BaXoNElRVC1zmGpKFPbN4MeX9acdmgzb63k
fq95GOXTqd31SMphuMHAE4o2sSnrVpUVg+zEyxsoUf/vmfc8UzSDu1xH6cYbg8lW
5pYsl4gOHc7arwjrr5jHcvNPkGMvaNVhDaiJwDDZfkgLu4ohJxcNlcXYbOMwCJ/i
4Cw0oiX2+yphngvgL8IvOrIj6Ij2iUNLoxQu/YKHsUyw+a4lo1OCxKZgYddIgotF
dFmjjloKwEg2OpVibaO24ihlB9WQ5Onsvq3a5uG/SsMTMKN1ZVzuJr84xCYTKDgi
z3CCi+dkg1I+q3XRZLJTicmSGIP1JLW93XQSyOaogo2tugQocBmly+d8HnjQu+6B
AJ7b1ph5i4ZXqONAysV6Y8LP3V/X4AegzBD52EqS9iKyo6UIpt8lHz1+bmaNWXUF
iI/9PCd8epgAxUXGK9gtty5W5GsFo7G/JILuneOmGWWIaIAuld0ej2qAGSe+JFFV
wrWDIoRBQcpH1pJiNHdAT461FybDyKet8wxaY3fu7jUF2VLTQl4CEiTeWmmvGUSF
Hdge/U0ThSWpgWcGjtkgsFJ8Xz6uADXdOwm1wu3ir691wZryGC8cG5QV6TAweE6T
jonXu15ecJe8sdrASbKYL/9SFXiC0Kqa3GU8fNrVYmb2kXtXFYtGirfPonUXaDWZ
K4PhNxTukC4J5f/ZmcgEAgu1xMOYinstGW7vSk6WByXGmGUUl82cN1sNDyRx5sML
jQ7UDSQjq8tQcELdYuJqzVCwxiqduTatVn9zi9VS3TdSM5SFidEBKMASaTWp8+vw
k1UzyhQo3YbXidX+5NenEmCTha/jgMtrDUNKCIzD243NrI7op51tlEYNBYNyo/cZ
8dCqIwO5URJcxxv0pjWFYWceBXiyIfUFFCp4L1nwpdr9XgfzQNrucktaURRNOUQG
KM3FgnarJSHsDu4cwmV6o770cjfIryS+iSVTHGXxfpVFMmwu76+Qry1y8wIc1+54
+VqEsmPHg2Ee7PR0SmLhSTOXFmuQaBNiJ4W+r2/v0CyBDNtATvvRLjR/E7+Z9cdL
ulYNc2wiqDrisXSDQc4WKZb9Uq6Q9Am0GBF7mKXiSyLGTGbfCQMXKIzicht0UMX4
DgcK4AFXQ80XNdzf7W0x+JXDrPHJiNWjUw6+ewvKN9PZdWiQ22SRaf4KBPypj08g
9ltUPiJaOQNyHpru6X69FASgCUsFdySTiw+eKTyoUnLrLEkGeW8K4hW2VfpXhxGj
gmpzuFkmkPq7gJWXeqNZh8wNYn44sKidGAxaHRrIBEaLJZe9w6GCV4m8diFVA5/R
KJBkLtuVXleWTcq/o1Ar+m0Hf2Yjv+eHiwCKe0lWc1/0sQ5gQDMsBuv2bJdqNvJe
CJECcNRO+9PTDKCkJdA3VZUVoehJ7//cYLLVVFhrWIdO/fTdktp5snA4Jwj7vooi
u4WPoa3GptexITGNTc3AtnU9QgAYI2/VyIzN33Y2hBEdmWlpsuo69NIHQiWp1rSg
tBD8CgU+J3t7dgvEfBLlNBg6tQLrKOLtb4yslbZY3A29zfPUVnDClEmNnfUKpP2D
OIBBbRLMfC+ld5ztokefNTGqcXHUjiswnsSuBljJFGXvm4p8Xitjwdm0E+WkNGLk
PaULq9SsFNtPrXBlZSJrqBgUCCtQVCipVUFhmLAnwhrl5MWCRO0NYPZsJ4+hSnid
vFMKx9t1+quJnLKPJY7aRxDOq5n3rgjdVkko9Kner99AC9QPM+sWwOU2UuqkyEQ4
IMZJ8n6TYjmw/hsZ2PnoDR636Gi6WefUFdjFxmeGVy+g3zxJyaSZ9lSvZx8THNHC
yGrUHaYLpuxrQ7z2RkaC/bKfHUqtS+8XPTsHO2JxcnRRDvrtCn/AxcB0y171vkY7
QjNQIV9JY0zXYHQa85f7BfE2eD47YTduHSDy1ShE+NkBXuANPhH4pnhhkz8LLsiF
XqO5z02bvqWH1H0adT7b0Q2OA5Kms2J0ee+YyVweX+2XSqXCbvU72pPvszFXTZ+f
UO8sS5Ch9UAAKl3H6FQu2n9Ic7a0bUKJHbKCtWDk62Syxc1L61JoyIFtBgBe5CS8
CP38GUoXICy6MqGDu8ePsCRJYf6mZ5WEZwlCeNmW6YpL4P7ZvvXA91T1aPWZUj6I
5XtYfyEcdhOSrYNI66ZBg01GG6DQClxD+iceDHouCtIG4HIiyjV8SIgtnBD41MJq
tHf5snfScA8V/eHlmLPDdCAELvzMIU8H2XnphXzf1fsOgvkroeN9DgVzx/8CFXw+
VtSCZvLzFyxjryZ1Geb3Rq9vaNnLEPfH8DYeOCXV3J7mnS7pfJqsag3WyyfquoP9
ZPOYEMkePPQHpGncpHlC6KngJVMZD+SaY2duTgOXFlaSLMHENZULD5NM5LNCWV4e
5tFhOrRCrTvSa3v/3r4GiShD0HqsjObT/nSWTjPGCqWlQ5auzj4ZfR4eMDHRzuXm
+mX0Ozx0F+40HyUxGUDnkIB/lkX4c8O1bG5dT6XAJ2dU2Q3vKcw793jQ06EVlg6o
2Lbxp9/qRNkoxwCjcT+m2T6xAHyt3h0J0uMekSpVi5IArUe/DkxD4RX+12qALggH
GBrTG5Cn4w22GNsYUzVxx2o+7T9qz/G89Oik+B6WqhGc9vMNQNdRQHVUJLScivFX
34SY9+A4oXrm51GFxehyly3FaSJBdi5d+wT+4d6J7FnFzs9iuP7A5BIHUnmZR03p
PI3ErjDN/yoYPvcoIFnupwY8q31/3ylM+inf+54nYH3dQz8oY2f7IZdbeKjscTh2
wT7YK2tAkvcN2JltvJz/W9HPWUHCc9Uk6JabOC0eh8c95/hyIxuQcyT5cAHyIFtY
ntSUflau6T/azY+/zmFna9xSys8wfRG3Asd5klshUBiMJ6Pl3SOKBW9ya1wAzu1N
PQJqFbUsb7Ie8GL/s+PhotEYve+fQKsIHTWZ6YwGxPedIRrCriMdD2UUoLCJq6lH
rtZ1L50Nns/ApnWdmr8Q/0Cepw6bGh79XwuHgNOErHU3XyKzn53Dodr3nJUudOJP
3LKxuOPUNZfj19nDbNt5jvzYOoVOZmGYYVKnfg2VOIJADymavgLD+oTmSd8d5LcM
UJTyma1LADCkuWDcm5gstrZBUoTqLH0sEwre2SklFxgijdawLJddlTcoeeEsqZ7+
3BInQP83XDfynA9NPFMxBY29A6VVeeMM12V9QIewhrKEBAVfZENUMLwT4zBX6m/w
tVCGt7iP0sbEwekAqMeYxZw+uHsImwUkh/1mKRsrDXqGv04nD97mH8H71F37Ja75
i450Foq1ffbeyaS9LJ8T/NBnRNjiZXk7wklqPhA6MdRZchwM32gCsva3SL9FYIwi
XinWqG9caz0TzNnQGEaCtIsnaZph7f0xB5Tlq/i2w5k2Xi/ojre6OZdeFusPUfrb
iP6+kQmvLXJxT2+uFnYBULV0Cb0CcyV1C/2lP9sdS0P7gxM48dGuBcKurfrKBGpc
tgFXzqjP2NnRfKcSI7tFezuICFeatmvf7R0lvn603ZTk2MenkITsMVDZDAGcKcqJ
GLCzUwohzMlwYJf5JksMQMVvdC6/AN4OsUv1R5/ExixRLbhOaYvwK6D5cx6c5Rxq
9ZIAezvsSvncZgTvKhynk+YWSCjoBn13KP0/yMk9Cy98roPNAD7yiIOJgDkz04Lo
0R7dTHYhPOojlqzT5n3ysH1sYdFGzg6u1KCjNRxX7CFLEHR1pgOsle8V7gKAy7+P
+7QMl2lcWHIzhjKRbcZzuFKsGgwMwUS9h6EEoDZeNLpIvMDmY9Q8ZJhJE+53BMEN
O5VMf46njk0NOaAutszcOd7y/ZRzaCxm4Na6vNs1WoMx0h+FSfRBA5qwALp+dx3H
gN6mH1VNvMUSU84NYq95L0mEKjuRAanhvrbSRR4XSEZLAVqL3pBMBVw/QcLgilDO
GXgQniJ3RGad8bmaXE37Xirt3F+LqugzgwmaEPN3QcbtErwjOLJGu10TD8Wd3nFb
g+kxndC3w2ksW40UqnRQNLYfwatNKr0gaFc/ENtWhjh4GtKxHdQmqfo8Ik25/tvl
KIkAersY/tobQ34V6sq1zJfaeqZcBpgDyIamvENIKn8PI0SmVnljE/txPO9vSnaD
RfrWl8kQ3pI1TgHTPlX+ixFzvyOHKdbaAgm0a0x+NMsqCCA90ZXQ9uMl3ksLyXm4
pxLZhUDXzWZGjx4ruFc+cR9sMUBMZim0a3VmkLHs/We5oezxPBFWJQordaIbAmi+
kB/gJpx2wJKaej+vYHAsXigwvPR533oJlSEHepHcyaTghLMxzWu+oQEjmHFdmOga
N3meqnd+ubxtIAsBXRZfQ+bjeFiW8VfHGBtYSuyUIWaM8UMlHwygHpnR2FDdEZkP
FEKhghY9jCOObVgt8GZ7ypJIONmqbS94j6fWls6/wCT1OaeqLMwQH2D3W/h+6v37
zR3PFr4PIpiJSHgBoMOIFaiZv7aBz9I43uy7rz6TSiV/a+/NUGAphqjyvw1hM1ns
isoO8m5fgULP2Li00J4CrK347CQ5wDfyjXEJhGyM5N/1I9ovbLrF7x5g0Cer2JHi
okG6qxsD/9HFLC4YR3h+bbKWszONeVZxEPe6xiOITvMiim22NzkN3rQKae8Wu514
yyyXR4081vrjgZ5N9HIhhHOslWh2jzgTXrwSav0TqGWqOEVSUpQ5xI+IKpZ5ZITo
VGvml+YYa9W5jDlFfdhiZMZdPhAr9N8idfcsYoEFT/LhniB4b76aFlVYdtAFLYot
cdf5M8O6FkeswZg/r0eQtIEsWu/DpWFJLmW/7yBSDdth5l7tGwB5VGZMuNVlE+qt
zWjbDPY80OpQtJFpSYBNZmYW32pQcX15PqSlyUqGqNVNITeFT0zKkWWHtfMJjhs0
oahQp74pMneOyN9TTxb7GhY+ptVF8ZwDbtngDXXmu6w5NM4wdqrBbRg7B769TDhw
Ow0YE79xCx/nq2f3ukRtjnrhA5V/GMYuGz4eV1oF4u894wnn2dKSVsuAqTnLfZrG
Du1tAaK0uEMih9071sPCdHvAj/x3noaKRPrCR6GaCNNJ3VxvHclBHkq46o0D5SYr
oPvRIyjwsWe4MTo9uJ/6WrJnXfwwCt3ZpUIKrpBlToCBDWgnNMC+0LtEQSL9voS+
uoRn/mmYKsuHv3DhrgBiVc71FooexIPgLHHlc1pzS8+LuXUmDRIptty0Gm/3OsZF
gwMfbBXQ0OHsZdhINPrD18UjxRHsPwYz1qZIzQJu3OKjUdmslWSbQ9QHnw3ysP5G
KR96C7KfTjXAE7wXN0SY6/e/AfRslOFHROQx6DilneZC//mptrzcpbPg3PeKcf/M
sSd/r7t679pn4hDnIyjUCcmyChiYVoFvc3kemghYo60FUBUWsuGCHy7qEAUuTk62
GNTN+jjsyw/RsFfRTVrHwGcFqIECLBxTPal4KJIOWhVgBYNRN6x4v/GNoHpIhHpq
GP7JKZhZi71DynEmXxTbXstneQWkUsoZdo5mnx/LEUxBeZDeg9ruRFgY73NRTuQL
yrtD1bRxp3wmdcdi/jTdNqelwEa7g+b6inwwaJwsGWt1MrJmLbm6YryojJQ3mdl8
KQhN9DfpqeOsxWCBKU6VBq9Rvlh9sO7ouglsaHzrn9V7JDFHED2gcnfidcvDmDfp
fMyt8Da1VbYGiUghBcm7Rzecge59GM2EPfCvpUlJQDAavkZUq2eOw3q1OJCHjuRt
1sfxEHli2puwNqAeoqKtI+EPS2vqmHXwjxj2c3F6SNj17EmdtksgtsfDr2+mHeM/
wWjaXhq6zq/STg2PPNCumLS+dpNtbEnP2Hq/g97+bVQDZuX/cVDWrc9os1zmhF3H
RO3Z8ebQRglOMLUHDGG8CVQLo9Ott6wIrCEcS99Xyc6MwQYr7B/ma6MZxJ7WOBTu
rfwpXb0mfgfOMi2Bd4R+eW3g3Uxfjxx4BcW+ALdma5OuCGcG8IPi3jY1xd3EGgT/
PSM+tv7MElNeItfICVO/6Apfmm6RxlVX1gT9dP3f62qNV43YIdAmNhS7cviZjmNe
d+oLtQCVHDdLqejQSrWqQwneCYISB+eDWioqkxpwlpglnJlk9JXpg8g/cgVrw/qR
CoZJ8sEfZo/F1bRR72fsGMLxqPh8sprOnOteXGiVb0YzEFOHFczXpva6gNBHVGf6
nwjETZLR8foKd3vx7+9HbvMONBGpyYv330JhzBI623XrTe2CIhynQOdXd4Uzwa+q
xN32CMFYand5tAs0OwBCapS9V+Vr9TFdo5qLECcJLRtFz+hJERiBSK3TciLcaxKe
lP+3d5viaHLAHyurF6S2TNVWH5xUwN5+37X7q6wSd/831ft8USCzIFhONQYQl8EC
UKMKfS6EDPVDCLOOys6n+00PQjjQo0r3G3I0UP0Y0S5wJ4qo5Vw8FPb2SWjzfbRL
O8Ejl24+0UCcWtggLsgCRrQEg1Uxp8d/NfCXsz+VNlKsjQ6vIqe/GfrMS5BQgWZD
Hyx6KaEGo/WuST8lItRRM9TnRmu6AobrJD8LfztmaCgm90RM39Z5USvuNfZp9Loz
xK0CSP6kgkg9opcsiHfUS0qx4kCMCl+X+7ArRmANZBx7huvWVEb06/Lt4KSrcuNA
dhzk6lxNQeJYfh5SZgi1ujUcFPgwo3VXkb/QiP8z9Pyclou42DBVgm9Ad8m934hh
SQugRq7tQnSz4a4JmCNGyLzEAoQvEi6mi3RB7Pkbc4AmS9DtTGh7r21+HmdqWAG8
HmIpmW2gBe4aiYBMAHaAx8zaj5JbQ0/56RUk5mbGrmvzjWZFAB0+wYGKAVNeY6g9
N5TH6F9lespLG52L5WZHX/faa5HFICn3aytMH0wDCvmOcQoyI/fVsAwQiJnm2LEY
zNpUW+o3/Kh/QYlA588+PnbLNRo0ICnqtuC5FbeFO76XMz9RWFzyCMQxa9iudhNL
/98SRrgRSyI1f82x3z4VjtmNteI+a7p+/jWQqDjRPALH7vHnQ+VtqIzZOI4Opd3r
PjHLPrhTkSyfRfF7c9uz2omDHMOBS71H/kV63J8aqYIztaZOfqUJBwgCsvCUYCOh
bydkNQUNfbEApOaR4f1mlRiA+JJeHC7y0Sf5rCQuQhqeHdjx+EmA41vNpS+ivJ45
Z3dMm7yXi3V3dybAXbCJ96OWGk6fbQuyVp4/Y5gJ6mgIYdk3jI5Tu+zdgtM7742l
J2Sej76K6QfwVsE0YtQDxdmo/jYLtjVrMntzWhkYiX12ll4FB4DWYS3Jp66D5qDs
564GulKy0WOonEFKKTK8HU/f2gDTGdXrz9Qoxrjkx9dDX7ZXfcj3t8D0CessRTDq
+/vruXG16kCD3qsgtyAsLFiE1A2mr7X3xR12DnyW3aYT9QDb/D2Aac05xoiKPlaF
SwYxgKWaKKVfIXR11iBMnaoUYtJ8OE+Z76PBn6eVrsPwqPWEH9s76kQ6Z+fO7HsF
+cOnY6bPXg9g1TLIK0L9U5fsh/Stonu4vn/EJ4YWmRdXmNUKTorMESZ5TbAaw7Bt
hZsGAt0GCCd3nwxTxwl+UsFsZpW7pVPUtZpaaSCkYK2V685u9nkm2bzYc6ERp/+I
T46plxQ+Gna0Dc0hijMAm3/53HKgFauulkAS7yVf5decwyqNn1BA4L7EJ8QJACG1
dZUsyWL++GZrPck2KPKLUgXqiEEYdE4t7ljydfYCFT2M731D9gvP/KDRZqAW/+ru
2kKpYyOw0Qibb2gUZdKRfGequiZ5K7OEv4p4tON+U8EBvrpRSBfIJ+slVZhCcLIo
5a4P3sOQCDkKG1CXieU6xUr07eLBTWpH9A31aYfsxeTIdM8aiYsAePb8MML3IFoC
+JoGyClEjojMH9z8wQyTmwzaia7VVqo2M8Sl+1RRG6PpsaWd9Bt/Ns8GheYlPPYJ
ZdpB1DeIa0IpODAiz1wUPBHTy78OnAFj38vS+iGEvkX79HD1i3zZQ+F4uQcOhrvA
MhsqEpgdoNIF2+AchLZoeMSiA6iXt8i/19jKzW9kG+XWMBz5Zb7zBtnUxIMrcmgC
lQAz5XGcp/e5R/5/ppBb1sjVkGzrQjjRXCE5pOcQMUwWhKnQhLZ9FX9RnDrTtBS5
lWYVsIjkudB/Cu0n3SpnIwOANOXspdKSFH+CcQhcONUXXDvqmG8eJavtkpbjQpwK
yw784r/Ro9gHoT4dD7poZdEovcFFo8gt2HWOipmYBsm+ez4awACOJnGLrhmuh5Og
cn67xtxxUtnqBe5UafSbuB8n2ecHJrBjLXo9pJLrqihooyiDIOn0FgzJa6rjps78
PRFgefnxt4yHhKmBut2DUFy5dTTJFlmRCBb0Na2UeFXA9TVbrqXfrn4x0+V5y1vL
V88ETW08pmYZ99eEZnSeGtcEdb7TGz4w0KL0jMNDluI7m6haBmcAHjcfVABz8htk
dLzLzsiUtOS6DgXp2n8c4FEbZ6Z4u1VKYaxZOrLwwLxVtvxExuy9fQd00/zEC9sO
eWQ+eMH+c5eYwvJOnr65io6TFD0KvrGsKsGuJIGSdgiV2FlcP3tnSo7JlmVXzbbV
Z6cuZEwTtfQK8q5Avh+v8MDUJ2nxCII8tB6U/hkJslBYntTWaVXySZCu19Jt1CMA
HPe00z6kfDuDnC0gKAVcRm9Aao/1KF2KM2WbLLFTOo9CnE7ucxsw6W5iSF/HBFDe
LA+pQwZpD7gc9Yupb0lT3+jy2CHMwCO3ndLkk50GcZsleqCgos2Xd0yuYYhicWrX
pUeYVNSh1YigkgcB3MYFdPSOAYPiixsAunGfOOcznUfWQvy9YHvMZCJ8x3nExcTw
YhSThaRZCP/IdbFYAajcuLWsqJSdWHOEqvq7Wy8w6i4jrCMHnQdsfzOG2w5KbKOP
PWDQH7p8Lzg3St4wg8zmB8XDd5hkHrsxukeAk4FS/dx1H4BJCkYoWgeNKPurq5nr
34c8Ha/Yksl+L95jT6cQcNk4WEqIE9Nwk57xW5njP+JhaJxJPfP/yf04HdmD03wE
X/yL932Yb4RVlImK2nOvXhZBAEyS8OuI1NkEyqky8xJV0v4hG2P+H5L7BsXw2ndf
3QGMbPP7dSZPzHWYzr7QdHRqb8vZ3dhGuFsyE0RJXEE4m6adS8ioLQNKiebk6pez
Ve9ozSulIZnc57JIz2ARAYlX/PWXW6P1p8bZMRsB4WEkaBJim1dnEuci7b9hrxO7
4n+cYGIcnwVGqek3/sNcK9TqeYD5dZbTaXJxBoxEaep29fxf968xo8dreg0PQgnI
L5J9dakdNvGBMJj0ECoVFe3lYGa6eXvk/I95MD8sH/3dG+fKy3NewPJjcFlCKDDN
5PzwnEb/hpruyNenBA81NcrRJPaFoDG6EtVUhrrlOy0W7jzzjj6kuB+7X7Apdn9s
OdZtcRquE7Kx3FFqyBlO1Usqz2Bc6ZRAap+C9EE2xzXuvndOFaWlxi67p8gj3hf9
u3Hl7qKsQheG0fB2iCynl0sTLgwNzIxIya2/mkrSMUbGyi+eDp1jshT36skxu47E
iX/HrGYG/sqNj362ghoaUsfRWqj/TqesPpFc5o+VbkB3ZJ01wIv71fUpSzE8vphL
wxNjK2fPH/UNfZ8oAL8cFCYaeOdkOg9Pyc+ZKKvBoaNMwiybkZMataLw02BGoQqU
JfOgRomidxQpJjSursLhvyBOG4ACEYMUAbSAS/9YDNFaOFobjOcFNZ3Zk3HxztrQ
Cj2aU/UbsCRQ/jbdN7+A41YYN/hHFRUMrTcMAZSL/wJDjGahgXbHHM+2lpLx2TfT
coR1IWS1gdryJeoYQ84F6l5v9KIG2AteLaATqXqO14P6m2VkhXAPRHAuirjI2sA+
ShXzrqouCuP1x1Dc9Owq4vH8MELLTwFzd6yZs+pacajcSzyHiBZAAaFu4rTuNt5H
NTODJgRuppm9RzLdcx20eRjOKs8k2dZ/3Ldpk05P55WkCCbRtponQe0+vu7TgQa0
L9ao3s4xdXK6tSCNAluacwF2PWBYrugmHYVH5/p82Yq2r+5vOeU/IlKJuJUhv70/
Yz4af4JP95hCn2S394vOqBkPcwj+fSj2oj9rLDUo5zhmVCi2WL41iUhTHdzKApkX
oOnlE80qYDBbhgSshWmYadEDQOTij6Fo7X0xq3hUhqO7CQTbmw8pubTzMGsRyX25
SPBs3MhF43xvaq1nSdhc2WQxXjdpACIYKMtDbX1nEXuBOCPfUrxJX/zPXIZrjZiK
L9H6YlIJZqLs0zoGFxBO5RN3xquqKkkLRSnpvVIalraKTY0d+itxPDxD4RAhgvHU
rD7W5phYOLtf3E8WFH5fL+B1xVPKHwSOH15Z3xgVuM+6auu736KQ100kRjZrivzf
Hj7wJHRdcgeyJwDK+ySKLiB3ZYFPUXABUWWMxReDSH/zg6jJCWRoWIJ3jc4arnC9
JdnFo60Qj8t9rVsoX6U02eYcOZOxrpA/rhCwUTfihYjEIVPBp9zmcDWAamLJqRht
RevX3yil+7z8qxZPGI21/d8pA+m5JE9f59Vr6WQmIJJcXpN/58COCl27G5pFFqUi
mHHJszP1UT+mIacNgb8XN1pfKfbiR0HVIG/tHu5WRhSX6y0EcamfAoE0MzBr2yWW
E6awsLmXkWewBewol+ZjIG1X5W5tCm0uDDM1gIWiREj3KxToPP0vHVD+VPdnH5MF
Jx8C79ahDRPGAb4LfaqMGWwcsUGiuPQH2hnkg679aP6etXqp2X0bn4pJuJgn9HZw
3QjW8GLU02O4cZqMOzM3ADi3+gCBnaHyUkESuDn1gIg2UF9rAMyKRdXLtOxGNf4e
uX+IeeHO7FozxGiqlbFcw7mHPuStB4SgAxad01csouhI9V9J2nq1P+jyltFLgIqR
C8axXQxnt1bninR8tGkmTIrI8FgOjBUvyU1+4195IbI6rrOwLmrsDMfJ/Nz4rhfY
4rh8Stg7vNmtPPTkYQhR57pHAUSgTUaxGUk1bLkHaq58+48jwKVnQc3r3b1p3frf
tagrvpY1pmNy9uTGmg6Oy/2Bg1ca4x9MwAq3ZePR+WppCCNiebJGCw3pxJv81P7V
w09YMhWh4EXcw+fuO7qlms1Hp+CRKYJ1yYyGR7sFvXuFaljLJatmdO8XHQEnSmaj
Jp76xySgHqcIQxUHRLSK9BfIQk8Dd5Uu2owDSjBCcey06b1woNFNt8WfnVeqd8Oq
SaPA5NJOTiK9qQXifVoQ4K3TXxcOeuo/kevwkNJInUcKS1ZPuVJpwf79iAjY+5sI
D6ttN39fU0FblyMs08DMtHpbfBlqCyJawk007vMac/nNiCqkbJ7qHBsG8/Cpx6jl
OIUtzgpxrCwZMyzlgDkjnns0YVjCUmJc0yXiEssLeFlBj3al2sPgvsxedqsiRQcX
UNGrYlhAqvCUhjHa3ho19UxLKnP1Lzwlx6IvUKMJFIfZTPCTOT7sRf+fp95MUe38
GodmV6Cto+E9KnrlrzKoddYTuvPqas+iN08ZqgpH7gw/ezGBRE3l1nzJiFnwkDVO
xZmv6Wb97CZ5Wbv5nRPSd5nECtyWp/CVgEQRHdGjiAqJjUF4luHvcFtKj7dI61/T
ZCcWTngxIvSaKT/qkN8E4VsePPUpsuZBF6SPk/Io6/8bu0sxEqENPIK1UUaG4Xyt
rLuAJyjwz3rXwWQOR/f3fc+hzzX0u19eWlyVCflmP61a1hLcCFDEzRNTz3i7EQ76
bHQhQwWpqVzRHxAPgxjfzx/coDkP/dVxygDp0ABFS5IX8UjXcGUHUAfOfN5LWE/Z
AUPDhkJ9GKb2kblofwFrqW8L329e+L3s23xqVmHkdTyZb+sbo63nWgyalash5oVR
wKfYY9SjMkv42CQrfR52LnI4TBIqBz6E6ipK+Uvrjngy2Yazpc4Hbl2zSxMo4E75
/Of+rqpy1iayX/BhjGTB1ZAHNFslHehhAERS04RvQiYodBWwE7kcCVGsK+IhIRYW
Ga5Ei23DUhKB/5TkNNFiaNoAq5RlW/g1OdakgpvkCML3km7pNKcRYdLCAzeEd3VS
bKF1dyfuCMQ4PiUNYM/pPOJNL94NRmNp3ePruZlOfSklAjaWvZAXlp2kEPFT9ApC
EIEctIWqgO8ZA+XAaRoJfxCdn1XQH25Q5Yf9zkG/BA0jisOmG+mpuT2dqA8xoecB
6Jfpa2Tap6k/v+BS1n3i3lKoII1ufsC0RDUMiLckY/eDkiIP4QsbEGwy7lk/UE11
525efYE2wUQdn6gmyisPLkHhKisqBSPirIy76xajEkCm+z3prbRjoMXolzqIgVjr
LxFBUTurAvXblLA10yo2oh38S0/wxHw2Da5DSZf5VuHQ7z97CO6A6WRVjaksjj2Z
/q+fq9/pT+p1DJC1FJug54dHBAS8Rg3PgFp29570C72HQmEUQ3wxUKi8QnwxQFg1
REgPENsRZWszJj6hb+XryxRW4CfBhnNBeyVGCY9d3LJczmNpjIyha0xbTtCoEu6l
2S04oXH4ulCNwqeqJsIRK2fXZBFM2YBKn9RoHyhXJTu4VGh02pNAElGIle0H7fRw
t060sRTbNAQhheWBJH05xxj8T5SGYeMuWf6MXuGkVQSuAlb6g/VnU6atdss8BvjO
Df2ap3ZrHLEuKOCb184EieRdxm8rQ+eb2z2p+5NwcEM/YdEX9X2SjQC6r5mwiM2b
ff5wMwzyycGKmpqB49wQOHVKP9xzhjhg/hdxM6DWBKVeenUdTed8a5Gym1EvV8Ml
jRDCNMlKUmA3VQvld1uPB8G7IJ/MxVsfUe8jK6iOT+I7WHZ+NaP4WAZxA2BujOLc
EYcF3dqPJXP8fZgXoiApmwM3VB9x3Q/dEXGUReBLHY/zDerNxM63zZQvKLLFYV5n
Kx/dLjjyWXUiEytdjhHigEMwkyizxyfOLAkP1dPzKyHNpklT25KlyjPDQCssgY2J
jQA/Swxs3/G7BM/sJ6PNYMbTxXm2QfxMt78mtB6I6KIJJwzrF/H5mJcIAuYLOYIx
Phmu+ZMGVpwjwMJG/oHfk7+SjJYBvHUlO7x4JEZNXn/+7CFjyVMxet6CzYM+M1BJ
LhuOgkPoi5haeDMhNzSa9okp2ypEe+2XtRV4FaPNfZtfM3kZJSp9LRCa1Pru6N9l
JEl4IeweTFLsZBTCsiaz4NlRl1q7e8AxgR+6zq/MPwUKmZNf+SXdtJzJ+RHnVymZ
PsHF3qyeauHbk0CSiQpWSAmPIWO70OvC1tKTBIvAp03Y81Ct2/0epzvIBojFaUE6
ySEGP6mE97IyjEbhgaDrhX7dSnep2Ad5fmt5/7hKuX08gX8G4e+jvFps5icXylG0
FVewmwP6YnQ5ciVceX6DN4NU3C+hr6/ZM9+fY1VhVLHl3hPMQsAP01YLNwSq5AKW
kOowuP+f5bN/tP3Vr84wr+L//gasMDeV6D9m3xA+Yd45vAnlyyHh+GAdSqyQySvw
A/hxLKFpk1RarhYI+xHdzT1z4LNDtc1fupU/Iz2NHK+dnXYk3hNoW0aX05h4zWPQ
tkoCtU/xgXeimOFbeKweB8SMSQPlfw2Y3abLiOvs4NOLW1VXEAZj08SczQjOeja9
BDdhLNdv0VfldHJE9a05qfSaWslH152USEM2p4Kl/nM0nzkZ3zB79u5HXiQjGYF6
5knKX9xc8wlmN2wAPym+EE7KqLrQ3G0N0OdcHdhz+m8H3yNM9kSh9YNlbHSqfNvG
aEOIcEABGrCo6XoT8OJdpcAzOQxPCYaBDldBlNxqT7Gb88pOvVFI48wwmLeeKQqf
mLsakTWGKBWgLP3a8aSWIqRgX+p0EHNBTt17YvObrWCZSXnnJX/6ftV22QstJzng
Sm89l+pm+Uc2TUmUZDxymIEJrqbhH49IuLJfFrUPHiBw44SxILCoInlWzGrw6vnl
pG3NLiWK+iqsVXYKe+x3No6AsXUjn+o4TSWlM8hCezyB6lnDKC393dcVJMDq8asg
zoWgjDlC13eNP/TwgIWm+FMLSASu6/uR38xltUDS1cF18sV+gvIuat+mBvBg1P+v
mk6oXJmwxCIwgz/JoSrXNyRfuJrtHyAIx9ggXHfwPVNs8KlP3I7YZeaL9WM8i1U5
6vOJKy4F55pKo8xtFC8RWQl4Qsg/bzHAAUluYA2jZ03Cd48DIipiou+jmkPcLeNs
MRqshi2/8zl99zLQERiUc5VV2zyfYTXJB7QzVzzd0u1a+EOkdA/ISMrE6WZ6QIoI
M4YJrKoVJNZb+2HFJJTzRduhTncNOWCztVoF9bMs/pS+DpDIz6qLKFJiHi8iUJkp
jVDxaocI29QZ9XG0g0CDgwzg2TzOuVDJafUjGwBcSdHyqPKS+bCnVlwT9OYiWCfn
N1DzDHHqK5NVfv9Uzkb8bUXP8QT39cNGi53K7d/8bMoLgKZbLcUqYImROLvjo9ei
UVOtCzRzKg6/87HQcG+A4UGIkVxM16TIJ7pOBACiZGjWwKpq7wk0N0Z87QYJDFQi
rCJfz1vBYomunQ1eQ7DahyK6yiexXHIzOG3CGkIcsW++wEeigH3eU8otEccE7Q1H
FUKYCj+Op3ZhjvfLb4rCAsVB6eFTRKiOUlcgnsOCrODbGe3XOqXAP3KJ5x59b4I/
+UMjw2xPxXurFBh3pC+Q+6UgChV8A0RH0nJ6nv+JL2Xd02gHGsOhkb8sCo+Hf+wJ
g6lB0M2312SDddhrXTL/yRMOdoUQ5pd5txsCoz5jhCTk/BZDXiq+zL7qtF5KE5/m
u70ae+D2BgDhHYmHFlCXXM/99rrovifZE797cjaMYL6HQdTbDMg0NNOVguIwG7EV
NYSJ6Hh+K9diuheW9N1uKt3pIUXPUJS5jhCk281bo++1CNKUGKdwYjAgUxw1mHq1
1ZKeK1WgL2Rv6cEwxcSJiiu8/VxvuaHP6xXyLicR+vGY6guwQZwCIreuYImiKuPf
uObWgXO0NCh1AydnTUUuiHfS2kfOPhB65uwCobZZxsfOipBVgXSCnkNiYJ2zNvaO
eAkqyd460Xmqkm/y7q/ZAIsij+N4Nm1lzWzoPK3mzo/E+pSmc7vj2cF3dRWl9l1a
jY0dlQBqJhfZxxbNh1fZojNKNryCmeX2+xhbBVRYzyM16DBVBcE68LW2RDH4faC/
g5OuDa2JxItfD+pf5me2SbEGyaOeF0UAf8GSENugujcJXcST5Xql1wlLkheaBStJ
Mr6QsK0lIuM7qRkaqH8eNAMmxBLIfOq4Vp5sQMOZeTXWQSYQqQVdTeEnXeHr/r22
sYpHgyhXJVi0Hm6kc2My3qq789Gu24kWwW3bO2mgXIRnqna3dmv1oIcYuaUwnaF2
HDGSjlnfVbkc+HhM7EuvODR9eh8ODVdYHglOtK93GZJBVUkw2YQynhzmQwGv8d5P
o06cJucK9sCq18J0afPsz9B/I2PdvjYhDzLh21IOqPJosP7/lF4mvgqE8qXHFeDb
NmmYkkY3tfooNj7S+/3XK0sBT+seUiPmUg2vtY7QrDtiIgF7FCW3I6zPlbW8mVW3
KswzEStRv7rZC19OnQeHREYAy968wMk6F7p6uTCrHUixUbIA5yk/bSf1l9GD5fpY
oWJTnk/xqWlqSrCw7G9vkOQEeCyvLxivrTgNDLYTuNl0EVRgQwIGZslR/xP2tOo+
MckwklLFR6elr6+YSH5MQCKsvdLlsYkTKsL2em/Sv4NteLHTrWkCtnyjRAfBEYWp
MpoQ694ZiQH/VskYbjQZhwtSrVZ95f912azELionypgNanNKYG9o25LQS/4LnoZi
D04Opu6ZoN3SzhC4uHRBWV/6zHvK0NybDHIwAVjAH5qbJSeey+jIwJQEakZq5tnh
6H8Qdv2IcUHZSFj9Kop9lx2sh8R/IZOofYBv7tx/e2EtuX14ned5p4q4EctVEpI2
xHpn1BFm9jLfmKulJXAVfQ8kJXBbQCQ/mxp8YqcP3F8EkJVVb5/b70NLJu2llW2/
pTq+K+wTH1+Rn7BOQ/Ik9NuYLeDvQn22yg1uyBGijL3gmhZX3K+9BmPBM01K3C0d
YzaFEu4qaBFRusZpWBZu3DVHgtZzmJ8wtHobKPcPLn3EWtrB/Dl0uwEDQSzF6Xwo
2p43yiTtBkNFQDaZgECARu0oEpSZfNWTEL00HzVGQGQ7lmoGcI/3D7cmKP5IKLsB
3am9KiKNn9M9nxSSd6nXU1pnEoCIqS1vFS4hiynAYcZD5ndipJLSRsIKkdc/WYWd
0DweLEbkGDFVySHEaTMFYyz85FJZyJOCGkhsLF+ZemJbAZ2jUrxWoCdeQZ/3+Yo0
KERprAz+QmsZ40psxOWqAaopXd5uHf50TNVK1Q7XWdAVxQ7tUluZXR7pSzKMkRl7
/X9ZlZKp16hAIhqMQf2ZWYuamaYGfb3AF5wooFtaI/VWL7SURWCVlsJH9sYu8Uuj
1q1pwsDzSPx0zmsQr20BtVRX6af3Mqwu3nXpIxYCfBzdBi/jSkbnp3YsMDwl/4oa
/3zPYb1ePTOTIlLHUIQyuUkdKYvo1vCuQaU/71MGrUUNk5P17G6xWRsKKzBlj4no
RgGSgM73rhLom3cgoIQX0FVbNDys5YBoquAm5roVlG3IERpYj89MNx3DVXegmyqy
ImjcVSsdmy6HRjP63/9Zj9lWhscxX/y4QNERqxKyQdnv0jdJ7+UMLGwGnnVaejqm
QaV2ZoZ2376I+Z99SA8yutqVbQQCxNGzR0MpLW+7daRkiqbStcD+IrWPKqPOZS9w
sXw2CKQnmyp7mqDtoM4fpgirD5+yLYIf4jOkLadX9NifWZD47cF5AzNetVgODJcr
3vqVGKjqjGLQ5Z8ZhHXdJ2FDa9VMw/+MIfHiZegQ2rdc0EV4q3ro4sTY+gzJOrW/
+kabWLlcFeE9LVbyhlYsz0lBnaAYpsGYX09+YAmBBSSE4r5D7p3WmllYxmAKjKNn
2hvaPXDn6jpRzD+1ypwA3jJ05c+a3CJlKfiKiZsXj7TLopD/6sN3XsD0lw4AR8FD
bJ8TRCRh1J4XjFKJbxuo5D3YP9LQ9oSX3Vayx8b+4G0OoezXPZ1N8mb1CrMGj++q
9UIlWk+g+SbxHvQTHZiemnAdHE1cWJr4I+FmTVthwgnC+uM0RhXarNX1J3wDjdYZ
ypVkisuXLipgkg6Q//sxcxowWWV7h7o44kzkHNp0g65QmwsjM0EET6kbfDoH+k1q
hz+YteaNmDuficfthrXTwUHt6xvNnp3vOoAQTumoNHkcez7nIqrhvhoKR7h0CQgm
ZMAO1sjnMkpFe97Riy/+vAUvfN5OZGEDaHSSaLyfoKu1xXEddp/PkdXnea6LuUr/
KLljE3rQrGGJT44lbDbYD5X6OPgPA3Q6eqnUJQxGT8N0HhwOpTUkmicx0Rb1EJCq
oh3IpTOBH1uDqIjBcjyw6hfKeAxfeu4gdLse+xgKHyIDdgsjktgCRGTjyvybIJg2
80MN5QWRy8j4ckgXjs9zKTgGX5No3LR9f+Sx+hbA7A9CiWhHYHd7/nXaeaodtQgD
VY46N+ghTeg0ik01Ck43bYTdL6N5HAhJx8eFsbzrQax6oxty3pD1OC081rWiVwBD
MC0IAoX5uAMg8Aw9GJfW1RSPLQEJ4Y2zlYuJ64xd5pQ3QxmGoqpo3P7UJ+2FENeg
R68ALL0rRv5Wtv+uNRHVii0FNddwZ/8AT74xheDM3vI8sSPUwZmIp7o+kvyP45dp
rvVVVCTOF6rure0R3Z+fY18CjiicALs5p4rsQUJhoIoGeVgnmausJcH3C8zK9LZM
4oTKleWckDCh+GGwcwD5HCo2um3kJMr/mVwmMgwOzRdVW1GSQOaEtlEBmfAkbFqd
z/czYm30wwM18soqRPkNyIRZrN/rkuuegqry5g5DbwoY+cn3irrIUJVtv4rPqW9F
QUJsxSj7vESQ7rRHCy5xzxCdMKJL48RDDoa231sx4/HFGwVOs4OyGVISexaimLfe
9rqoe1MAjKky1z9PvnFwI+U7blrSrh2IWhgfoa1IiyN106wa4Xu74AFPmRtus9R6
nguBpChhJ+pFPtldk+nn+7ONhohov2ZG7tUxw2gg3xSkABfhC701PiUk9v8li2Ba
0cnQ8AXzgMhNMHPbUqa8FiTyKDug5S+ee7PfPKkrPOfZv9zgLZLSDgqhLKjytGVU
tUjXzRAVGxcGjFeAW80neLgTRLiPMlKnx6LKMcovDxfVE/ukqY8X8fQ+Sw+3+pTe
sUUQP5ZS8+qkPZvlB03/WzUDH4NqMzAMS4X/NraWf+74mFTreMH2S2qYXLC5/hOC
QPE0XB5svdrpjRU8qzt+MpfQ3Y9yUrW8bVLGYj5kWHN9OstokprApIBWua+wnHCL
mBN16kDEbhv2hp1ANuNkIxtcgnAzXujWTLXL+Q4rjygi+0p9HydkNdEQg5oDKe2t
UFywNhZ6M/w/BwajhOVws4kZr26Lfv5ylN4x+uAxNZDIoj+8AUe7EAsm24I1D0Az
Aol/xFHdPgKPtJnDValxvJNNliKVvG4tpf1OGnFAKruFQAQiBavjPDZ5NPySJFhj
j6whAAelo4P3SrSEY+LdziP6zX3kTxacH7BpSsa0+qo3tZTggn5WUNHiZgv4NLOV
G5YNzTyxY9QLNbHUMtILWfrZHb3r5a+koTWraeAw1/0r/fIwFHRbFnINekVN1m8+
EqVvCOiUu3SoIMEcZBUmk8XkKYlmPWSBmlZjElP/tiK8dv01VulkAMdpuiYvd3KZ
qKBcHvrV+E/7wbGL1XGBO9lDyGq0aKQYWD8lyJ+k9/TSr8OhIB6mxF+ZLfDa3fl7
18eYwDdssO61KIr8FwZfmc9zwNp708IBHxNZhF1XdGQCBi1aGgCct4cfqckXFka8
8csRiS+6qB2vcETWUI/MiokFRp5ClSj7fAlNflYVjYOEuozeqxENwZ5hUlsnHuYS
xPGTzJHL53Kj4wf+uuZhiDa9LT6OnDgjBr/GT5MHVYw5NhLIOYBt7rwe/H5iipai
F3tbgd8uc43SWOAAzGwsxwIIGb359PbndCWFRmNxmubJiunjUzFNRvHg82Wxx4EO
bSQv26u6n4KFOkKZkrYAB3rW2DxqvyxM5xTL6xMcMqAzV8p0eUaUhTop9n9yC4Z5
EGAZifbUUBxjHIPP9uGcLA874jolPFY4i7XsJ3wKpBAxn1hiyrqhR5n9hrD6aPof
0NUG8RKSCrN9iaK1UCWWM45wPbOpb2UJXuEj6/bNe7armt/kGqe+lHJ+KNYTwrwj
8oCcDNC3paxTdBa/8EGhq9pXyP+VMzROAdH9nFNfIbVJQuuEiiRsuuGKB+QbEUkm
yzNQfxDPyrR4L1vmuchf+2T1nu4CTsjRbknOSJopECFCNUfj9pxRn6QUNxrdNoS1
DN47VYO2xScCcm5B9e6EZyRhDMr3AXYFTfFSnREUy36NBWhK60dzWq5TbxmH8ULO
+HGMTL53AuSFQKmSG3mGiabBHok6zLb4F6lCJlm6QHlGeT9pkQGrUp7c//X+Nnhv
LPxVfUUGDkOr9R8pAiD6D4/qI7p0D7ml/YZbBZSTqohXCCeXLq+xP3BTy8zuy37Q
sEYg0+2TD8NDgun4bATKJ9BWWnWbh05uP2wXCNzz3o5FHhVd0ErxFjgjW9GftCw2
BrgDvrWEKplFTocXDyL2xGIZVWPCYiqXMry5LXbZh2S5NC2jeTVbMNg0L0UAL6J/
d0t9Ov9an6oCyUfecsusE+BIcGjboNMnWt+UoGCM0RmfJExSk6zOZCNVmuZTHmAE
WL5e7x0B2ZZUAISYJeU6k41cSOWOXCVsqMbea6CEmJHbRO+q6Nm33i4HtIZQloa2
dNyPA8dUUWqG8nqN7OXYwiQC56XYI+1d5k1+IQxMNeHhJZuobM3FkmvcR82Nd0IC
vGlJ9Xg3cmowK/5yc4upJC/MegyvXNRMV1S+2DCOCMlgHC/oG0NFPblxAQ909zPi
WCVnkYGwR80ylRmSPsu2YkAorOIqFdqRIHhT4OwAm6vjD0Idw8G3JDdLJ6sUiM88
tW9UMr/lZQfQqja7twtbRGHE0oNf+/dagfxI7zVE6GUOm/9AQLf+CuFTp5lkk5JZ
qggzVegDIey07ivuBFrPseTjOLFl/hvAfDZUq0nKDIypOcgGVWOzTZQ8zXqg1ze2
92vXruVim7OAnWPIvAMq/htAF0+csGh2re8J4vCDcJDlXixw0u8ruhKMje8iUdeR
+A5iXJSBrN9rTVmn6u1m2pFiV2yGNFi2cMEUy2HfkbQEeRKHj5su6jpHf+ezO8pw
R4GrxdHA0ahTdHmVlEBKlttc93UzJ+sDM1IxlDePqz5o/wjoy/mmIPicfYtNRW7N
twTM7y1MJ3kHBq+VEZl9k09wXIldcab7g3VSnpozcYR6fpWzvQnlUY9OdpYqQVAw
znUvO0AMfPgiGIf3FGo8qxKQn0bbuS+trE48Bj+5tBNZBp55mnY/coM5pnAHiUdp
LwLodXs5ji+optoPs76/5S+QCXmuC9ek9N+GDe6O61e8EFg2GeoYvEOiAiqYgTLM
fTIrXsxPTYil7Krol7jzEyFo/irS+saDmdL7mkF0Y2HuCNw2t4RhIFxGKQU26J+U
13idpKRKPPWdoGGqc4ckc1j4sPHIrijqXQVFE5LrXfkfkzGJO5NAmqOMXmXVCZMG
BucRlJlp/gfxDw2lHwf0ejSWEFhEC/lg1pPNT3r1zEt7c+akeZRX1rw8UxxSgUKi
RV84+LR+Pn78dGqg5clp8/OnpMNP/xnvkb1+xZuJQi0tecW1EdvvdS26pQfHQzx5
zE6TQ2RUWkP1VWn/6ufLyNiTLfTT7fTBAOxBAT2MWkIy6INZviPlM+kH+gTrVziy
aXAZX7IQQI3WwZkoMCbejdxgR3+N9B75DSzjs6A8LITKIpw1AHNfY/KPLuL/jQn/
cCgy4evIulypkXhFLDa19/duQdtHeCc919Vouj0GAz2qakQh8Q57UPP6iTQ7meJx
qarJJRsw7fAGNM/Ir3E/NUZ6/MNqdiZDjMXqiE5N0AExXC7nblmgMPLGmhoHVurB
f7qqEUugeyJ/ngMwY0PfJ/no1fDDUwA0r15jsXrORV39zZw0ckqxmFmNNqRT9ML3
K7Cnwr5FbUotO+AQT6+6OgTKtffQZ+K2ZOc3Q8UQDH7r5B++Wj7YkjBuegT/3LXs
LiCd/Wl1oP6n8iHGVJZKVmOGSWVLPD8kmVt54dLeyKCyhMJ9gCIN3zOSDE7cH/6G
ulS7m4mA4qEG8088cwLG9ldpNmo3KYAQwwKmveTH007jDhLnXfBIFjYpQf7ZevLP
wDMp9Gc9aZWNLkmvU7YSsajdFwIm26E57cr5Ow9j0qJI5esq6Kj8CHDJfy6CYvoS
rZU/dp4rZZzWZdD+HAdZOPQDB/O/iW+DKOCBxiuQkhD0fL/9YiTfnVp4yKQrWuuz
lSm/SSqOTXlPtdGvwhDbi67osSupnDw4w3Satwq/yJh19eVhsNyi8B6OvDp5eNIv
64IWh0RjOxLis+SI378ebxjWIWfSHbSIfnFFKlCuDox5gIcUkzOYhTJMFDc2FroO
VABCMbwUyJro6H4BW+GmAM7MZJ1GVkIsVJW3yW9+6WJfl4TTWt55W/+9GUhT0uYd
ftkgJ1libDslAf1DmHUPtrlkoPW3wBviMgus/4vJOM551o07hYpSP0biCuIfgFyR
YTeoIFW6KuKB+XCZiN3VMy22ovN5I090qQgHATnQMw3y1X84iH86x7PYG1bJfYm7
0glSelVgN5QN66p7ylchXY/NRPLtAtDzMVMbcmKYuUQYveZVEb6JYPLz5y0sczrD
Jd4BLXGpuzzwmzShkqdxsO4AyMlQLDYB7IsVWGV0nlv/s9lsElvrvBnJold1loqb
uekXJvY/Zn0I9/aFM66tGDurAP/oSuMT9jQhTSr5y7x6dAK8eV8qHmC6WMNEG6OV
09OcRBVaHQjk9mMg62iq6w2eegr/4SgngLbpnyzJEqY05WCQbieIysPJLWAJg0cs
GmZu+cJ3LOEZUs+ts1p4clyNI0vr+Wek64Ut0Frbl3IH8D1XA5KXcLaUppg7WYOG
fr4nmpXAcpw5IzvUEs+y1of3QZCYEAJFdOIMr3voHX4GfpW0CFyniRQ5VbrsecjD
hBn9ThPyuSdRentf5/s3FEocyfdqDVnx27f+ZXS2CLxpZpKe6r4VmDKGBC5CxJDu
uqy97S1T7Y3KT3ryERggx/5NVzKdWsYZ7+W0rIJQ8fMJZKbF/kyE90jeT8zyU44Y
uVwf5jedYBQop4YEEU50bC53NhjIE3RcVWtgjOaug0B3CH0Pu2r1YX6QP5AtNVn9
aSbuUeEP/yaAXW0NXm1S5WpUBR+OTbjk+Dfm2PrKhFgOEmJnvq5yGciX4gGXgUo5
ZvsV34izUYNX2kNLwkQjGqnhjzawSlUQKmL7QlW6iX3kxcGqOAdUlLV66SEDVFQJ
8DnbuOr51ytnVEvEjrbz2kl06X3I+sQQMAOL1t/DZla23qlAW7ee7s466QkVqM9w
eRJf5gvgvVp0wFvkgs/FbL9g12zpeS23CK4Zy22BdiL1aULZAIHvLd978uTLfkg9
SOOS7VdVGg4KEgJ0Gaaqu+VlDiR1ckB0JY7fBLjtLdLDAAlIesFY2E93RixqqsPi
Un3lzkyYYJXjwSCEFBYBoaebFbe+1Mlrr8qL2f4SS/JDILS2v2oRO7DQ1p26TKsZ
4lxVFtFnWFI34w8ddYsk9k1BPDvjGIDMdhGZzvwMxnN3qjayXd0ANps+fosPhme7
JBQ6Uqbs2tvCCQSxvB0JBHIttfXq0PhywAXyvZi8D9yezoYgw9aCMKFvuEAxhZqd
rP2hWVhXiLMFCAj7j47wscoCf1MoYSJcUuAsQtBZIC3S48YMyO9R5o47X+QvFtKb
UDa8qvGY0OukxMRkXMghA0dCn23AFWTm0EwCjftQsJG8dOeq4yU85Nti1ObGATBm
E8Um7eToj9Ahs4G0Trm8BlCtJx1tyVS2b6YD/wJi06NmikqSO9u71sKbgGnV9HZx
VXR0xqFStHVH7/dDcPqKs2flbq6+f/lpW9/Z2tqgZWj7wIE2IWKEGeRgwDqmbnjT
lyqVd/NCRpukNF7pY0MUne51zJJInXJo+tOstuU+Lv35205eCzEclt3y+oOIIUBj
X7mJdniyn5pFOowZ1WR7/ZSEqKV6JC7/gQVnI0pelQ2zzLBt2B61dt6ct3+RS8Ir
KtqXTUDs2ryvhyNHElgY0hvmX4GSnHpeGfwkkn4jEfVzJcoxc8EQXNlld4UDRejj
ppQXeYuj9hntkgnFL15l7xsOrL8Zq6gIDcANIU6VQVmHw0eiKsLXyQiCkJAbJSCn
Y+8BDBDDFiy5R6NHx3zeBhWtsgF9YKwk5b6NoHh2pV6gRxf6Ot7Mr4PIBCqiqZuC
h27RsZSQxPYLL4v7eZp/FxSAXmJnyN6ozth5/ajvSd1BYuesbv4vZi1JTzxGb7FD
RLXg8LA0tVrFGurPbbfmt4VgI7+bRMkiMRwdLN7j3Nr8hzzvkNXz004d6dBF3rD4
oVTWmvlqGX83nWE/AY0S76vwEjFCIZZOCxp7sAy2j0LS88rIcL2qnCLRZ4Hm/qid
winTw5jeeo8ceKRPKuR04AuIcZVirHxZTcet0nHxppPfRp0sk50AmOLGA0dvo6uH
MpxLjOe+vH3eCl+wOCbJKY6xDt+AbVWy6mYGLp8r431me67pjTZozD00VJqxM9+H
wsN4QqCw1VYTY99Uw5GFkgeboZR/TgD+wHdyYx7U3XzIKb7plD4uEBfBBSWtRr/S
ZYsuAfuB2f9q7gjAaB/Z1pRM0W34b8s49tWKxTiW5cOLF2U0gT9xk7d1eNV4elhW
hbIvAX41buKAq239pOmNvYZHZO2UNcsMTO/zUvJsy+cyI1ZV9or9FJu9uHsETgtu
0LzHd99WCWXgVlq4C5cKXFlctThkLJMW7Ke3Zj2je7l/MLL8uokq+30Ncvytpp0K
jQ5o0oxA+G/J2bnbwYDQLIPUtIN4qwL9nKL8rwFI641+vQ02I96QTojdvtTIKhhO
OLSVsohAjHYGehlCuI18myIxyuf1GVmFtFqwxV+OYYNipnOl8YV3PnAK/SXbvktM
FkLjWSb65B+LcW7X3RV2hgKZP7NMJ2OHNQclekHb1BZ7nMNnw21yVJ/k2SKOJYXA
Fi5wODPUULX2G/Ii1HKu8s8qpFh6ADVDgJ1fNNX7Uq9P2dQqCLFQCQbybTCsIyg9
Q8zzhsNhwWAKuwlPjK+9kAjt7gwo6p4veytfdvL/Myfj/yTSopQvxtGM2a9I7Piy
6Bk+HG7GBVOmNQmBkPqbKOXpgEZn0e8KWK1KOXds43PHrpIKR0MiVBwYvUJp9AMx
tKPEao8/rHaxKHN2mjyHxv5vJTPC+ONCnZTNl94LpgIaJgvmkbAp99BLoeUjtUtn
/u/CkImMPaDMY69iTWasUc1xd5G417Xd/d3LL/RzlsPUR23s64xWuqj+HGHo5m/s
XO4hYhwIQPbpju6tDTwPsvjHEJft6dnjM28EzwmKll8vTFWzUcLOTtO9XSYxM8UU
DNHy+QGbX+5YA7cDmgNXe1pZb5adhRYJlAJD+64e0iDEdzn4sWFebToNuTNgW3AC
PITTl+lrw6qbfk3T5Kf/LtWprby/vgTFaCBt3MEZEeu2dF1K2HNoMIjRVteyuQA2
nu7XAA5hmBJRBZtZJQzHDqVz037M3f6anFB3CuXnDSGDbVf/2Y9sC7pJHWCELxN+
naa/gSXVl9KxJXTtFaGa9R4ZpU8kvf/DqPneT52Mf+f9kbX98T7vZJsEeW6/V3ue
Cfmik8RDJYjeCkZEDMgc3Ip926Tz0MCAyFfVnnXUMjeHyKdiB++TLVyMByOIUuiF
aOcd+gMEdGoC2xCACvlBbpIW2Pe/rFSs3S/1XlMCQqNReytOySJ25OmJ9lyqLeKe
DOK7/DdoLyE4++L7eH9d+Bgippyl6V/YhusbTB9ITYN6t7SZR8S5qQx8Rf8rltY5
cUAdaIw2yLAFIEVo1tBuD/5TRWwvKBgZEee/x48ntptA+pwLqM2Kz4FDfiiXs6Jz
jnishib/0es1z5z/eUU48Yr698VfbUv20rcUJPtMI32fcytZDJ5yuENUiTjLvGTc
S8YJMNKbl+Qcwt2+KmLcZDS9hVE6GsV/fXLwmGpM8bJIVaEGldyoZODWLctp11nQ
gqvZltvWk6iBmQQ0P31o9hIEUvFsCg13ISdx06W643VcN96hGMou5aXKgILQMhSv
w48Hh21tYHNGqNm916LOLSwKS2exwur9c3kcla9IYaQgYXqHSmX6f/XMiygkyO+E
MvFHH3ipfU2UhzyLuPTvDDZnqNg9EapXb6MNnQ1x9LqGnbwLPguNI43VtY0Kv6NK
ds7vSX7Pty0YXdFhpxCLecLxcSb8v4bj4v8szM9UnJEuxEBx67JK4i3rOYHjG2AL
JcpFFmMbmI9X7wYsf9Ln4mNojNtPTVxmzi9ayCLfW+NqEqSH/jAhS5yrWG7qI8pr
WZdv4/hcUlxyR1szDQbt85z12d0KRbloq5VOa6wBv+ZF1jcnesztMLiHieD9DFPY
YplHyAUhuHsvd93mubFtvv/aupeivxuIKnR8/u0GjV9awDG+YZdaC0hzfdfWFoYk
/jWCWKeXlN4so6jEtuPaP+UMSgN9Co/zofeagBwv4mKUsJCe2VZBy3+EqewUraEA
1GoyNiCU+airCETrnE3kps5UH5+7h1/rpegI1NRzayRg+eTyMDDGAp+NQxYeMRSt
Y4cJQlFA7CA2lPj1UWKBuBOCK3gaiDG19rG8/IkmfUOqExTQoPUF+8QLTk4PDVX4
7v0yTRxnenM86lmm2/rLUYMKxolm5I2PlDA3pFP0o5u4tcm6SPaE9ZhMeAoXQLm7
q3NyupOGpDvhXx561czdURM64Ccb/G0GfKEhJEhLJaT41wHh3E1Vu4Dz979z0F8J
UVxr9k7UWmXTdaDmyYGScqzrRqQPivjvP8eYDq3yO02s9kGUqMy1IhtGxJJ8jf42
Web/cWUGUfEQOWx7jIcqGn1RFM+WVx3SuOtwmbm5w0IaojFVqjVDmhlrONOelH0l
MVUpNG4phx5HFqs5dhDYvMym05qQ6lRro3tZEw0xl11bYX55Apg06iq/6Kt5xMWA
ICZp+7sSAJYD/8e5RYtC5tOA8vxEdhEzutGLZC3FDVZZiWDWdRfuJ9eHU0z7V0WI
kI2kStHqCPb32bQcSwtG2shceo1KcitzseO6iIDkGk+N18mGjIgvd6tdr/Cbu2SS
2/+VZmw6Tzq59sULTHCAdK61/bWC598InqBPocWLW73P/VkLv+bUr7+A33QJcWdO
/Uae5W68nVNfBQe2oqxuHNXa1EBze6FSpzErOvuKwODbIv5T5jbCGAtWIxGeRDaX
rPOwgXhatYNWauPIRGnCBdZLBKZQ2cLUnRNooo45yGQN+gTmPZkeByRmBEWvOntP
cZGGpp+3R+PzfUSpMq2/p0qDMkb1Iojm5C0aeXi7Fzsg8C88Tp/DJ8nBTffx+VDs
xr3D14+y7FseXhJgpfc9b0jEpLmSsMGwhSMfHpgW0eFVrWHl9yB4curzaJQeX7OZ
zQedOmTdzMS4ZwpA8NEhIORqG4BOEGZg+DSWQvy1bSQqItNu0ryPgW1LwTRqH1ac
e5p3jige7SFAqU9x+tJmkxJQ1rwQaFAti5XYtP3p8fl9ZUiZLYlvRhdVmx68af93
99v6MSZvD4RWmuHhTf/hnw9uSRl2JwnnErlM0ajXqrG6JnnhtoVemOr/bE7EpZBG
EkJITDeRPXSdlxoe1UyHMQd2kxYNe+EX48DSQebogL9VVThogBTLrZZzEve4i7FL
5Qi1jHdslMLaWX7TUP6IR1AfACq3SOJz3dcyYADz4QE5qZEZtY20TaH+z1eHFRci
0KvOvm2a8GrX1u6HZz+H41f3B2mNPUtM4qGVlvvdKRu4XJuBAzN0zS3h6j9uKz68
qFlVRaRWFS2Q469DuKa8taSbvcG+i4I/PH37mAdJL/j8Se1YoGBofb205Eqc7Bw3
zrZg2CsjXBLOaQd9j1L5sv1tCf7wPsac/5b2th4pTMDzb7VJwwIYnikMlUvceMnT
R8uPsCT3Vvd2O+XQdRHXcF2fq5hCq+vaES5Qd+ddQSp6+NfLpcn/a1jU4/vIf4hA
JLShtGfzxccfo/cYOMNRa5K8YBdE/zodySh8l2VOx4p0r/Za1KSKrm0lHuzNJAfy
GaT9t6VGxLYDOdMibNGF9xdAcmy4/vptZ7sLL4LrKCXI+wCeoQkseGuWyj+dVaLN
qIbaNZmckUeQ34dfP4+dPjyi+2M0kjk52H2jYPx5wFPjzIy9rtX9cfMUGeQRZGG5
WWz+NO4GX1R9D5VK18+SpS+NhQhqa5bn74UAC3G2+4gcnnA+dwLXJZKw7VifemZU
GJ/T+XBM8x3PcNXRuJ1xVU+KtTCPd9gsniWc8us4Nw6je+/3+0997QSyODtdu3Bn
t5rN3lcrV4IItAbHsn6NNS+zyXGLK18B2QBm4xUHpZJmbVF7Zaun9WhY6/22WR/D
EiykiJF/aQQbsLlZtVKBxcd8hLSZPEsyN7hXeIelCWZwZ4Uom3udRy0CqkCkygMl
h05QRX318J23k4aM54UvCLWHaTJ9yXpPnFgOsXIXeLBqrDc3lAvIJkHMKvCFet2B
tZk31tUI/ovKStV2NTCuj3gZ/jRJmVM9QrpQteL3qxMZWtp5p9DeTVUH+qJ7k24/
jspkOd5pa+E4RYGqNp4YcBMdhDq2F1nPc2Bsd4bm5khu5CW0NwMmxJlLciOBeysS
eP2t/JbEViG6vv9Htlr92SQv0+uYczGMTEyD5MtiRvL0JLZKJIKxxELU1wRwTBJh
ypEqn0fdWElSoNlWLcu2ZN8PbVISP+iHOkv6jqsVZQVjbxW25WSLwU8fMzBbE9/W
GE7U8bZNW73/+CsKl4bnhnHQtvFIksFcYrOuMxGOXb1gkKNcA5OmD8ca5IWY+ga9
MsekxO05EqrMtcS7DhgXsi9c3ahVt5aCMw51xJhcEykcVtDufzNaVWo3y5eHWsMg
7F2vN82ZnXchPjTqJryhmZ8ohcWrMy6IkNgqgKFQ0DWznfzBgU62rVGKrm+8iB1B
VV3UvyQDhmT/Ku/iy5gsApDI++4Y+406MAws+ifuy0VMLon/jXjjl1fMtB80Hpb5
iWql1FytKr8LdnHT6XWusbWih/SRHxVp3TmYlvmkaUdn/YM3T6+O70xGrNxm1t0R
kfAA7+Wanp88kSSa3OoMML4r7FN8lk9OkoIzBVCR24QFJqmgUjT0yDTcNlC0zg39
PiBk4MyuhhrmcNRyB+X4/ak/pgh43dgSK21ztPW1PtywkaopSVufA+qtpHQM+l6B
DoJDljWJyKGUOTLOmePdEd+AYdZClWrOKhmfN+4eO2YTiIK7zkhITl0ucqdj0XBU
L/omXNUVt7rJJ70+uZsRGZ8ubTKgIeSC/rK6jD2gPqR69LFh35NkSil+I0w80+ss
MRWuC/JmvZUgvlElGc13/N12yZF9I8nBMkhQ/ak25o+09awPKvyODx9B4FdPQAci
XJAHHsQM24sso2B2Fx/ju80cRCYqJuTshLztjFKnRlP0gmBt5Xm9N0of0Qd45fkW
y7MUhkLCDjVO2cFih/vSqM96vE5AC7MtcBMG3KBCDAomNtiSRYFAmoTFs0L/uAo0
73nHiWgKy6jFdGK5cxP5rTLUv7C0/kgdXOddr/DOAD8TXOjZ4quSOmldqpijrJ7W
ZgsqFc6ogbf2jcHlys6ZCAYoL4/VCAOEr0/P96XJcJg2ffd45CCwSdVvfa7dnru4
blJgPPfrODGSGIu6P1SK8mBnNcTSiRMBLzsrvqsefncNgZlEDaLiDyDAYihEd8mZ
TsYoG8Il2dkXdxTvV+L6YZEIv8hBHhmKuzEMqsUYT6ykn9PU3bvpe1OCP46ZN6Bf
zdOVFB1k2E7PZ0Ta4AISXJCj+R4qwE9d1CBGDAPSnIK8WzDLRh76DWNAKAizETng
kttB6PtNysQEqVtqa+ALZuUyjFiwovwdT1xrgdO9MNW/3qUVVT/HVsG+RA8u/Uq+
HXDxPpQFnZEVMiidQ+O2BIfqLvkFyMXRPhzCFH+d67jftjUqtTxiI9j+GSOwQx4T
XHhn0UDCD5psuXfyilpqzVeLWMP1sIOX3ztzS+C3CETkD/pS0jTNSBesWAQrwgJG
PaGckqfMsGWAVHJ9FQsAC8vPgRfamkUM5hM6TLPsAE48JYCdcT3ZTji+79vaW1AS
HElKPCn36PxH94Avk3DObWsvEc4CxICY72G1T9TLkHs9l+XrtBpusVnnbinmcNQz
ZO18w7bWaCrVA56IkHU0KnbFrmIw+NyWsUJmwJriBF1XL4fmOsysRnDEjzqgLiLs
DLCtkFjudjNDis+jM2Wb1DTVmTbdBP3Qny7L1h3ZbxqYyFkmneMdw2rIca9+y2TN
jhiUOQbNPOGm0/97wbyrfiDTufcjMMP3Zl62d9OTlJHtTL7ZBlXKyR4UEgwK9lhi
Qepp9Vbtl6MpkclT+456aPQRYLsGCWt1wrAforYpju2vySAjEUTAMOa5lHQjTXqp
wSBvTmWi1/9rux6b6QIVNtmx57ulOeI6KFBUJfSFoUnrfKO0JOAT02Xv0FCoSyA+
xkA2pWMU7pWvaax4neN6l1XQaPe8cU67h9FizlncKDSLQc3J+rbhFf/mdIYcb1lM
uw9jpTZ6ceRGoWDRqiB0As7F20w+z5Cf5nqyAZEY/im03TsPTHjutUp2CFbsNKAw
zE/eqTGSyolrl1MPtQkGnbeaHH2KXn0iMx9xi5FbcJMLOyLPq2RrR1j6zEYGju3e
0KNUWHrNn9GXuFMezSWye4qodtNJDeT2+keRXJFef2ALGoS/KMrIVLHMz1CotCrx
kzwQ3V3DxR5x8AKa1SchO4fE3zywiRj/HWK+cmX4yTiR0pfkcWRd9oJkzARa8ocr
s1zU3zPX/aaXg0/bD0dP3LQgxzyCymhDev/teG5uPBElvpD043RYdd3OPV5jpjUc
pTavJsRnU2yKeP0GAAbKWsGB3ew+NaJFxDpQ0/TUSpTxJCLzBk2SPkezQxOJNPW2
giupujog5EYtGsDOp8qXMKuR8Lb7wtr/9ANE/Qyd6293SJGYuGXufFXt642mjgzV
SuZjSNYTvDCHz6IjvxAfM+y+gXMJbyKdLMaFL9M5ViKa84t1TX+ST0EJtjCzjTTG
gp49+zagiWZ85uZiGZEtGCbOJW1beRGNJu4CooB0Dxx/3SEdUPMwrBr2vUyL0fYg
R3/vNwkoSs691PPIyLHMtQqoLqTDX6e6GqC3lTIErItT0riEGXsIrGRf1gqu/WgA
DSqQcLUBckcIpGi4ZzFOubo4W1MKlCmJeySrefIfKA6ub4NcFGccUiqNC8ab6qrQ
B+aTOPCk99OeJTK0doDGQUKuFUWIpSl1CT8ckNB1qVdzyvHmdFjJpX4+N6JRRnW1
GrERIWMaxDyoamElP7NJlVMidZi7AsCcmAhJ5XH/ynjEHFUPLoCVMMOrN1WzkL9t
S52w7nX6aP4J19MjntUN5kUXyxvM7JVjTISi4xk6MUZt6r6kk5S0rbbu1FsW5l6h
9568MMC5n3p9KL9LWMVRAs34X4Xrukky6ZYGlfxSDVkrO11KM/YYm78lQfsA64uL
EuZFicvS7rON5Kftx0XE7S6Kj54W/XrqeXB8Qy8coGhM6dpNBF0g/cCRKvrvFnBR
OFMY4JkSbdiBkbJOcMTKAO0GuqNGFQUK/H1+KIOohYtFu8FqaaXi3ba5iS2W2N6O
dPPl5kM377IJpuXFrgO/BZ5tiOak3Ie9Q7FmdmI56hVl8mI//bzlThTF65AY9nBi
gFaaNcEAPy/lYQ1mEEdXldMEnvHZNRcho0UUJQhd64bCWZmBNetfNB8EgRYpAhyG
T0Jb0e5Q/Z6GbfDr1z/t1VvZIsU6X33zZFUNh0aiVmU/yT44nZmOtlHQQRJbX/Vh
6VtQzOMygV/YcdaP63c94Rgj5UMfVyDbnbSHkVc23vxsGEueLZY4c0+CM6RK6Omu
L/LV4g1O5tYChKm7KP7LCTUda1YW+BRAd8NzK/rzy/y0IM4gMZ+HQ985VEIlTorb
qu2z0uYjzkwMLnos2nFB09ICkOBaaB1LZ5zXVg6ihoMyiyoExI7jCc94LTB4bYGL
rOD1i/m97KxEhmy2MhsEV20qTyLm4nva0MdLbLizMGNcfi4pW8Uqn8DDXQkwZtBP
m67sRWbc0F6NM3UpfsRCy1IpGK85OVF2VVnP8gnMzHVGuLfmmr59Hn7+dZ7PGRjo
nOYKvK+tBJBjr5bXhkC4wzJ1nqeORZaA5JsmNAhbznEkDmctE9usjedKFIHDmX3Z
65JDtmiwsxO7d3+IPONrzG5uesYda92YmXumN7nNMO2GKHmM9MshdWphuejUdvlQ
FcK10XgVvzQFyswgtFPJn6m+lnyGckXHJ63h4j3r6gX3Mc/2QwSa1BHNcJl/4cf8
+gArZj4B3+K4Wo6tJf8UxaUbQ0IXRFlgFShOw6D+PzUgLuuIAILsZc00E0CMYxxL
FJciulY9vQNQlUdo5VzvNT9zmxaLigyNzUwxevImaa0JWYi8kPDp9yPcU4cmL0gb
lXLwlW1SE/aY5vyNRbjBhW5Kblptbc4lUFx+WQQ9UnT74z2bd30dFNZoKT2gUlfj
gACW6IlVdcoEhM9pif9InYXbOgxfvJXWzgFCYVAVkuSJtTmcgjqUNIIOuwY3OHoU
KtoHsmendZHTW2XtnpE9ixLgmTjFUDXIsX6AgnuoVQ5cy2sNJUYxlGf5DDSxJloB
sMNtQYB1ThBip5Su78wjg7xOgAEWZkvYZMNVyk2H072Aot3bLviSe1CDomvkz1aw
47b0KJRcGuMvzZ5Vtz3bqNjokPhwM2x/WOCIOchXnuxsMxv4zN6BAUB+gWyvJrk8
ztb55fgGosQnrvONaOon4jY42GIK4LNNLrzryuUWSGrgrbm3ImdFz4z+4XdOwKIG
nYIAPnRkxiN4eueltoVcA9CZczDjQxIoYHWiMn+wmEia7Ns90IGWbBjg2ve426Ly
N8oK7Y6GntuBInyWRS9Jif3amLIUqmFXtjCMEEBcqB/er/w2QQY6xKD2Rw3R/vDk
f8jMDQUJ7zXculBG8zo0prFWUaCHocuCXHey4CnkqyOkyE9Hvk4qJWnSLBVjhI20
qzSUd2epo8AtKoiGCotOPiqVvXnKkt/QFJd8vqaLmRORcwruIvBQP1IVGTvihtVZ
XkL0I8wJb5I7hsxx/gfkhuE/EPueDL3Tc0oB+Io+Oj02DDlh8w2Uk/qS44GbrL7s
Ctj0HGhUTifpv4EgSrrUQpuSDWrAdrk2jwtTi3a7hiC2QfbjbMJn9j3Soyca9cfB
O+Z0ZUmgoGU7ems4n/QloJHFk0cJxvkAveov+NoW0J504Py2kfb8U8lNPGRx5ucA
mETvziw2iokl8Ga5H0w78u32FD9qsXeg2IkgLL/FLNdslI1zCwD3ocZhbCMyoO+X
cn2LgISU+RF5vKA6aRaNpvD2RQjDr7cJALWETIwGHlsmu0k8m0E0a0Zqc3FvbET5
RrRkG0akerXkon4bTqpYgR5kz4MccbcZP4izkT+Z/rrrxGnlUVTFbgm7AmXgssGg
Z5x+va/YNrQTj7BLBVoLbtRy8/FMOb989NBnMpVvxjdYTXsNJNkyIa7+FcPOirXx
7vu9B8W3fucdK51Wpz21yP/CyeRx6fOOwUPC7kABM0iQTXnMTT+0fRtUHrDrCGVZ
Megb4xyB4n0SeMRTuIrh16pGsTLfbL5w9oohJshH35Z//ZA948r2AdsMD7+iL7Nn
le58QYwvDasZO4gwjYGTpOO6wovW55AZtqQXVVw/XuVBji8JV2JPCZ+LT+Znzdnu
cMXW63beREY1yvWlKyuycs88nBezPLaB3p1Z605n+G5su36tuWn9FXGkOta8q4Ca
GjSYxv53XdTN5tEriTXrNd6ut03N2YV+hPeFDexu1BCG8dQut0EJi5X8RBRaHTUS
1gf31krbGSZHB08YL32iwYLCHO/qlZSDcBkz/uZvC/J8szfR5x1QyAGJ6DhE2tHk
Lmi5VDHFKxzaUkvw7g2UTI7SiPYh+8hcvomsY7F/dmaZrJpdlZD6Op3LJ5bBYh/j
4sTiY1ofn/LM2TzE9IKVT105G5YnX2/KaKMenrMGcwtfZzfDSrHAdZUgqZPHwJj8
BEo4DvV0J3wy3EkJ5K08jDIBN9tzuiUEzU9GtVTGqGVTEvw9RLELvM1oGwGRswIY
AlowfvTwYdy9P7Uid231dUkZiaqVAFTLzBXx9XI6N5QZ6TFEWfUc02HCS+OfTg2x
8bDwjvmL2BXphhlhDWTqcLrlBvJth2wfNOnnuAaiqicStMuI6oiVmIP2ylPRxkEo
bUcmETju8xyoJP6J1/6BWydi/LwIBZS6yhVaExK0GTCQJmFEqN8v1VY+FQibbF0H
TRKXY7GyZ1yUDt1pdxlYDqSYgOPxZ4yGrRIJVYUW70Nsw70aXEf7aSJQ1Kd72vL7
ISzPcoOTEhLgbRSNaWiNCIHzij5KaOvXgRgTTIX2FMCxDI98xDLC8ovuQK5PEK0h
eD1STnW9aIqUKCTvemwF1kHUFtrsB7XSuPR4nKL+jJP7O0L0z0PrkH9iItc7dLGH
Y8ulTmqdOQUmQzLa2nebKDBinf9bfdBeXmMJzDn/K+zbq0xT0OIYY/9Z2h256ld5
lldL21IFtfcdxxMUzB5Nj/DQDP+vDbtaIVeyjSzHFL3w0jy3pRzzsHFa23TvUBQv
qcmy4V4mCk3NmZK+tObQIuKUawVQEUWnCxVDf3kPUF8nA8KilPr6gkhNzf31WoE4
PXRGuajlfB5pQBd5LJPedaYF9x0xezh0LVycMtMGRbATXtNOb24pLzlkg36MnKch
czjcHftdCL3JQGOxZAuj3KUZMgG5eXH6dXz7ckYVsKcwPzFUQutqb4M3uI/nxwI0
FGFJdEqbdgVbxWXfgve0kgoZlgvUrYzoj9geH7RbMUkC69/i/risCiiovr+/GTsZ
hmcI/AymEC4JBxBryNiNmLObJZU4tO4iVy4Hhrpcm2EXhA2PAXMU0NjV4l7N5U1b
LYbZuY0FfPUHIlUTRvLFYVrKxClVGHlQomQA9zXGCYBdqy9fBlyZZ4jQ4BMcxXox
a/AF12jhe9EumK1WnUHFtN256zP6meghR6GA7dR9fr0ayfRN/BrKW3mqIH5eOTsC
aIImZ6AYh6KbaxR2pPm1a3Fm6QSFm91Kr7Y3oj4o2I4OMUHKNoNRUzZOij1stqNe
C28wwZTc9bDDdiBzQ3AFCW6UKSiKKfqWJJ0GETtJyue1EZMWa022vQYOQxDFUQYG
LU86gH3nzMiCRj+2KZyPyjPurWkwkpT49pLBBGma2zwjVHzzTEc/8kNNKHbQGBbf
MtmdKdlVK3tr6NocPArjd9aqA3aCdfC3Y0rHxFYOBhNgeO/8yACBvmlD5lfkZUYf
XMb012hKZe+VCxkJtyQ8R+QOI+1qdBmd+/p0QMzW2AStVOARxj02YYJIQBa9ukTX
wC/pGUeID+dO2JP0zJJFYHxMbabX9NzYLw+0GXZU30puVrOXRKuEwVl4/mrc3ju8
D9lCqqGZeakXAa2e+XLvGYTCGCw0nldjq7mh1IdiCrFvr/u9//WREaIb+PsQpdj6
IpM66wMyHTKFXr/cNFh2gBR7iQQ79T9/1jCd0oN+O/Ohh4CafaUj+rM0s/zqqTrr
aek6x/Gjc+ssYl8YgXvLebI2PSzwce8h6tIRkjxdF4Cbg+KvPHbzKVZ9JlrcnpjN
FXM823rufdAlvMAYSxIZCa+cdj+cka8vn6XSKKkJSil8i3KklQJci9GNT/P7+Mif
gs6DKejNDf2N2rKOxmoUSZjtHCXVSu1K4dxYFoy+HFd7x6H7E5Kc5F6HdNuaqPH+
wmSfEj/IkluFgwVUIAGUjUwed/EwOUlDowUq8DZcSio/1QmmtSmWE6nBf4IKremn
v9/ub+xOzkJy7AuyH1JtKw==
`pragma protect end_protected
