// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J3vb6y9h1CtBlW8W+RfONsiJ5xuWzfMtim+lq9agk44B+5eefK7t4F/cJpLeINlG
/gMxCpjUeKnazOWjEg02crtYPkPA3YX10czuCW37iWUKKpnqujYL8AjWEkJn8/By
kVvDBotJDvhawKJMY2c0BBdwYxcZlzUiFl8cm+zVUqQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10224)
XsfxYr4ES9+8ocUrt2vPTU4uW70S4pwgnqGN+QfESzDH/kL9l1BtxqYhWF8MdxPm
tiH15HETzhhORXNzxr53gaza0eoLIekblDXmxg07sa5Al4Wo8DNgTtQtCNBuvmb5
6vD6jhQppQQr1YilXeBMZxPnf24FkL64hvCILMCX8rwGZ/7kAPC16q2R6uzT9K5l
1BtmFA+5EchqpOC0M52nvi1xEBre3m5+xOGiWxXO0KuVq3hOj8g5TY8GyII9tyac
Z2FnohKasXp1epqVBOIVOpbEU+TS4c4G/8TCRL/QJxxXPV73pfqs2Mh17cNuqB9b
uhbBm1MS2fgix4kdF+J3ns70hspjgCa/E7IG+o7BadNTkSmu+bwMKz+ImucyTLij
APBsFmM21uJWWgO9pnZ7U8tUzHhX2nNDAdfQVj8CLwhGFHyQuBnojU4Ekn+ueYDh
wDRypUJYu0jIAP+knmqeoDQtbLs2qvLxeSGq1nKnJ14DgTqU7I6LPefrmM64FEFo
p11Nfro+vglKPMOeZwzdV6e/QJ+kRLUN0XNbhbGkT7gJrrg7GBp+S0jt1h0ikJXF
VG1AL2z31vYF3lS3OPZa2HKRanMR9iRTTtmAEraAJfa/64+KcAGPepgeEg6bQ4aM
z8hESQCiZSc0uGjYzMpuEn72R+07SCW1epoHhVuxc2CdSP5FSgBg5PQ1l5E+2a8y
Zv5RDeFYH/dbYFXIJbn+MhAk4eCFOgIa0FSD3KX3b0VUW4W7LZR7c7spNYVuuxaT
P6icsVCHVYywo5R4wFq0o3Wih8RDeud15+qHHf6MwB+lM1FrlLKHsAQ57qWndgve
ztgZPLNDwaKgWqnlUe+iyG/Boo7+PYuUPyZmCk2iC7gmF6Lhn8AZ46DZZcjWQsR0
NBUIDO5IMLA0kfvPY+sM6tjfkQH/E9p3Tu4vFCxd6jdcCl0pWb8HS/9a1mB+HJ8E
YXB4uu8inuqTqhibie1G5E7Ce8JsQJjh51LZD3ki6+7/QomT55lDxfFJicoa0MiG
4XbHirRWao4ZP7jIHc/rBd1eB15pq9gItvOocRFm934OolNk/Or9aTynVjHY4dAh
wxevEGyjbJdMf+YwbXPgxhrmIKBk3DjuGeAQU9BWSzZ8wYo/apl9MryPh1eLqb6s
FjiUCKljzW4v1oKQZfrLqCksopze5kf1M3r7BWbsokULrV3K5fsaIPJ+8ipgelgp
W7UtsZj4i0AeCt09TTqYVNx4tFpgBrlqy4/spSy5fP2N5A5C4kdQhxIm63XdJofc
OX1MEOAyUFN0NsOhL4TzTJqnX2IzjK5ckUGNoiIKv3dkdQw8wvaxkE5Ud0dUJ4tF
0DH6CmRtunWy6UA+MQgtJzpESFTJrp1JqhoIznJ/V4DbW8jo1Iooeby+6F/6EW8T
XDzOunaDKOHhIL1X0rGWhWbqney760iqeknWrlN8MA8gLdpHyTOupzY5JOx2iciV
iWu7UP4dQMtnc8LesVVlP2yF5as7I9Byj3VSCqbmIk/zUThm/fRUFCqEwoKu48DA
1sTvSPPAHa3kWaptEMBsXgIMC2OHnlJD4YP0NlLqFmefFIpTiLZ046ho9WAjkCB0
xOu7btfJ6q9cBdrQBpJAb+ZbkvZxG1WY5iRdkVW55A5d2rVdhRnOFifaQHucziLo
kKh96tahwRg6k8py+/wuGV3jwDjqfJgq6SIFWxT5+E/VUcjacEkWl/MYU0BjPir7
WvwAJZLlY5fiPD1lSFR1lcgSQFDE0bb4z//t+QJ2JYE7QHoTJNFqS44/2vwSCd3u
/ETNweP00RRYLpAyk/TOYKmRstxQxXKt+bBVVyYnTyhnQEJLvZdto2t+vStmr1tZ
pcJCGKAKUyghVJqz+TaymQp/6BUg2dsB8/RsfAV9wOEjI3rTPiMIts7r1CK1Rwi4
tGrsQVAaHcf63RgQBbHiYu7ln7QXU7dMuzUwApV2DwNYWa65qseO13C/0eQlnvor
xnMZ1RiN8PLD0ulZ1d9iyXfzcXQ2TjzY37bQfgLvHy+EXaY1XyGX53igzo4+6LEG
4pDiHZk1kueyTOh01Rfp9A/GuKO9gwKBoS+fpEjpk/gKcSSKMeDz0hjAWccpPvy2
D/y8MNfMLhwElndGerrAaC0Tlzx50yCKh4FkMMkQRxKNkd/4Iwe5jjbSxKEk+Ni0
i5fk40LrE1R10xz4vwJd5d62bn7neeBjD4Pif1f9GQIJ4+dCzNd7Boi+IUaQSNHt
4hstUrh9c7rWo6z+BFuBWUv1MPs0U3gloXc5cSM/vgt6VK527J1HJCFsmK9O9sYQ
KWyire0mkft5MQKAq/x5tMBIWMjFDvheUuH+rnn/kF6WkBTwOfY2XtwW0V+vGSZi
xux3MRBbtztoJo4JW+4noVdqQ+x3cghLUGUgNxUxnNsPbD/tL3PWNDkp3jG9Wm4C
ctALZPisqgJMMMHtuhHMfMyP8yowfainACGMkxuPZMZdkhYRPpV57/2mPBQoMs5o
nadaZrIEBi4a+JI81NKwEOhWWi0U2nEjmeFNujSwKiLnjgka+kSG+Em/2OosuqTR
iEXXIRtYRJJ+kP5wJceYhVSIrnaCxj1VduJ9Ay9qqvL4m1n9sdrYFRuYOz+C4Ac2
IQAjrxn5OF0F8Vm0u4kRflyKK22NWvMPpA9rEwskXaDLLfJ5Di/wNIv2oOPTS5Vr
lazD3gwoojGnz7yJQnpTnuPft12Z/2jHeeUylfNPN4TlK0qYcNScJN6/xNFSt7ml
xpVzF/MhM7ta+M3abPphvlkbpiplvUJGtVuiY5IBvhVt4fKYebfgehFDATX0sOGJ
t6bG7szWllmffMUnsDtTO+rXd6nGhLA6Iru7PyhdzHmdnP6stSZX3glApA6G75zP
+p++3y7fL2FDGLt5PKAnDrdX0L2QqPFe5D1H2glcR+l/WvCvdFpN1XfwSTPCpjB0
N2vPyeLSPMiIcGxgR3eJTF9NA1rHcMxFn6WlPSVV1+8BIUx+mD/s+oGPl5LaOEB1
gzhXPP5UHCy2dJ/EvZaaUJIE+Fty6RdgyKsjmsZS/Bmss3F1F4UtrIZ44DrGiIRX
BBYtfGMJA5NM7Cvr7lQucqaN893Q8y3hwh7dCoFL6uuGKdOBQQrY3zITlGg1s1uL
JtBc9v4hY3Op3nrph4gcsHYC5jwb/gJc9PaULL/k/eSsnQ21j+q23CG5bA9x0KRE
lbcT1f3ABEDTCK/r3oU5Sw1lBI4PbmOa6yeDAepanZJwWH7ciSNS0i19XUajlY3l
gvS9RxNZPdWIgY5HFGL3KNgVO+tAUcgHp4eE03uDToNS8OdjqqgUUFXydEvvdUk6
CBpVUUZ083Twe/clQtRN980iWxpVyZU3ZY630ABmai29aOfq5KyP+fpVyldnlwG5
ksWEMpWtQ7xCQ9w57uXXdehOJFCmA1LxeD02KTsHcDWcuC3UT+BgW+pRFvcM3PWZ
lh2b2Df4alBgqHb8F1ckpujwqzciSXTrMPwLnajyRR7tTthW5JigCKdOR39yIPZv
wMBHS4gC03cRNCRsoUXbuACBW2FraRQO0r/7Yx5TUYNL5jFc3pbQ9EwmMbp3hK8a
TrIdGgIxgV3GgflQfNPOUGCR0qSzreOCIxVhRdrI1Rb8t9e3CM42YWGgRoaDTaru
gul5JfqtlGxEztMWn+TEGbMQ9bQT5XFfqVbsZJpAfCgMdQt4+IE8j3AjjTmmrUZp
/4wyMS1aLFitLiV0uXDegIyJXQUJGF/jogpdIjCH5LqIAC+Hs7rrW05dhz+QVHvs
zoeR+DTnpEao+5YZjrLNOGGQQZFYSRG9VInh+pc2/6npsP/+hTvEwkZCiHtr06bj
ielwpeXjerwA965euOWFXboZbUjMuQe61xlhaqximaa8GVeBsF0GpKd5MpUlbtOa
9XuobIvg1KzzWvWAn1LM5PhSVZEu+DPevysRkWngYxH3CAHC0N3Qn5EpxexvboxL
ekrDrGBakB2AWj7Z13ed/SUFcYEsDjKguXBv6nW/yT/bEBzq3TbX6nroQ/VocdPl
DWhlL8/PI1hGbiDWSfV6zw1iu/bAnmX1/sBcspVwgGKafLkXKZ2qUxyz5rRv08aq
fLbU/egkMp6/1H/VqTBsrSYcFliuwyVBIiT0yCPcuHuN25L27aMoU4bBOpVXM76r
gRykCLxQbUEhnbvO/4V/Scjo1N6g2ljJnin0rR/vlCUO/fkwX6zmvcHYUIi6e1Pv
uN2ARgVz7hkxJK059XHtR1a1LeTpVcXLO0OtFh+L2mywwebNqmkJKhRkIVV3Uqhm
Ljid83sRWvgnrr2cHDiJsgS7OzuBliASSO3xxoIGTGCAhMX8jEAPHxnRzIVQRXY4
QmfujTEb0LVulV2wicvJ/4TiF7QZpCvDaTySO5HYGi/mxsas075Q0pqm6Kd4mjD3
NznwWdQMYlFzoMvSs8IeH+o7Dv8bNUk/fwaoYgLFsrnQ22PcrywPKK+DOTomQ0sg
we91GIjpQsfk2xf/ncho2hBzmvFMW/N+Ky6LG8mGXsgcZtJUse6SuJzY0P8EJJdP
Bwlibtt5/iRCEjW7n0MLE0Mhlta7kO9+9wmbDUqSGhRUUsGDYzLgsmwucSbhelaK
c7J9Y9I2qyqHjrKcngHkDS1auTGPllwqllP2Q3WvvlQQ1Mj1XE5ERXgZmk7XZJOX
2TqW2LmbHXa5hiE1GY5+h8YqfU62isBUheLEqn38vzvrtXPZ/2v+iFdHcxoNUkRG
7C4n3bV9IqiTOXszEkXs9u0R7sn3KGK5d2RDNR5rq2qH0Ed3TDFSJZY+fpmc+in1
dT33FjB6XB2iBBVRbJuzYqUMwKBtLxnA37AkismaU5A49xSMjx/nGZn9gaCPYGct
BgwPdluPj6ohhC7tcyZ3WvXB4FtxRlN3ieYEioWI8TnGrxbNLTWKTVy8yEIoSeE6
6MpR6mU6TH8eowBpKKlt91YxjhN34i67yj2PveicYAFbUoIVf5bkELUU4wFlM+nG
u/9qeTav87sUhskbc8g2eISzzpFr1tjidubF2/cbAj1bN50UUPj9YCKUTLUtte83
RM7K0Haiz5CiN9AFCiRSBRK4a78F8PqS0+jDwtjdoKliO7CyiTYNB9POyGEzHhGU
O0PMfsK6ki0U9yG2s5L4R3fFaUFm8H8tu8bWM3URiRNApcTuIdCmhS6jOChBmBTy
OV7niaSCiQUVD3zF8rmfobYuDelM634XcDW8Xqazu5bTOqvHe314DQ9mzZOXhdLS
DCXTyoZbWKmoSitV59v8ILRnQvUMABXNh1O1TKz3+CtHtDGLjTx9a1wIrsF4Q8C7
BpH+Y+eHcNFKvCmk1FA27WuAkK43VFIMli4tf3fIGgqFwuXVihJawvdaVa9qf1uq
slA/b9SAbDL5Irq0WIsD1Q+fu69BerAUgpnTBl2FgXoieMxd6niRTwgkzIvJpeQG
8aI5LPE1Q64AZZW75SsKzGHRc/7ykA4TLQ73OZkqWpi7afkrw00YLaUZSE+nm9DY
p8eF3mGtMR2Vwyd6/6ZHRDkYvK4d1T+QqXAkHDouEToCrcWR0XdpeVsQLufgMjmw
V7+2ibZHwhFDNR+4ofsIEg67vdp3sJNQhpyVaOG+d30Mnk+f9erwSjKKg4SeKIbF
qm/KopMltpc4FF8LW1P6gS6GXpCctvKyjGySlzub52JTUYwxGc4kkRl40ixRriy2
EhTqrujMfcQyKFiGQKBrVlMqcc42llIXPpLYGVv75uMzwY0Pgah8mEdQUTDMF3md
Fj+UFElm+y5ZFcR+p06Sp4Cq2ensDStHR6aMeNCRPSlgjXBJC2jfohhafKlIIbud
XvNuGWzE72GN5dnMjEiGHGamU3wTkqsjXMQWfKK49wB4m7VjWnt48ygrQxcwbk5o
5BeTuJUsCHq+nY9vzWmXnZt7q9xVEThHPx6EN96Z2ew5MwTH8iZr9smV2afkBNTo
GNJ18BEzKPchdmOmtoI8jR/0schLTDnz7osai6Oj66NNwP6qhuSeBH8upMqFKSPT
+XxcFgnoo95KeWPFpLx4T1JAmZSHDigFpQp7T8cHKjGbsUS3PLsJlxx5WQn76aBq
xEY6EwEU4Qtu85k+o0kgEzkiPrEz6r6ck+jS+dtZH/KqrEQXVF14yj92anaAI1Al
TTKFOC8tkVPWc/rsONSG5GAkhhRPKfzY3tPBE9y6gFK6tB1+T8L6+Hhj6OsMlMbd
UWOv0o2PWoroQV2lEab4yJFusKJeXm0V/QcVxSoaXDeVoBje6Vcu2PB/4h69Q4Nu
Ti8qOMYP0brMqwAm3cSn7huTPIMtckovKUhnj2QEDoLcE7kDZHxNUrR2YrCI/nzB
kwEqfktCOYNTT6r+dMyDXUxn58axOAGz0YDuihxCUzcUmoAkyJgLww69cR1O5+8k
jAFA3+XCSzJQnqjFBuR1gXpGts8eIry6DaD3pfMgN76dd6IoxKCMuUwo82N/doc6
nNPUNtHid6z3ug6NiBWTcCvJHy1MobT6BZHRac+w9tw+eD5aGi2bsbh3TPy2Fk9V
gYj9o5ZJVAeHv3b4NOheYYJStbdOZvpMRyRm7mJBFMxO2si5ibB3pUkGc2cOgh4Q
whnrTeY4uos+9fnEV06gGB+AwW8nvYFp3AV67y+4KiTXTIpTVqg3mZKtDgp43ohb
DEn0UvpNLWljrPJJ3eFbYfTLufRfgUuO3bWs/zbdXVl12v/Uxf+IpQ79aL+kONJK
svIGrCRmz2HTLgKBJDgcaiXYuGtYyITsPNNRc4TlAwEXjvvdSN1W/Vj6fmDYIl/1
KUFVrwToUq/PDmDKYJo5qBPlhGestFk0Mwha4+TvcJvWk6XGtM0CTSRApsY20GX1
+Owyxa6QipSeUQPlOwfOlYN4qINr5fiiJLmx3v7zvNly+xnt/9BBrMbrNWSiTGXR
m1IBsZmqWV9SYuKSU2uz6t+jVVjpSN3zwY24pozpNr0vWX2t4TFrZ77ZPJwvhv6x
9rkeYWYU1f6ZjtWjoZMnMGlOzdtYa3grnhGts0E7gL4Hw0GGkLUua2rvHZagc2u0
08KVndSgwssyEMGqb3aLIF4D1Rca2KvWhGU7ZsJe7x64XyXdrAc4SXD3IqS0Kltn
NqOEMzYya7eW+09+sx/zIsPg8MVIKyO49ztpPKY7JYsDZHgFkhRADgvsTCSBYT9/
q8LAUNv8knkWQuEpukAavbc/gdA9IcFb2PujwRXKZqCFZ/A7L+SuFO+LN/PXJw1B
GG80rYt9mdVTfsQmxMCEZvBq9EhqAO8xdahCfYqcyBWVTjjpyGLDbTXF1SrHrgz0
oIQACM6n7Ket50MrDMYvqaHiqmIl87Y0sqloANsUe914dbMvI4T1tUmjl2X1kdIN
hu/ENCtp3e+9rYzHjKP0NP3z8MLET2OhtEAMpUnKU+NsfwCJe5HyG7SPDxDsROgT
wp2jCgGlN0i4C9IU2tyrND2w+XRZwZsmRIUUz1tGN0s1vURSbDbolnf8vzg+q8mc
9K7oy7bOBefxlN1KLFSMj0wj/46qmkUccfweW8jRX1UAXb2Br3RWvC6dWobigASK
dTbj1SYPh1zYZy+Rr0CTufWR1cGhdHncbJKokOT39OuOAarjmHNfreOP2ztMO49Z
/B+PRC/ut2OyQG1uucKrvOBXHMFOBlcDFbyESvXha8cqbhQePO6Qp+5CLaEp18h/
7+wv1Yp/rPZYKIzqZJTl4QQf6uxOna+6mhSRdFywqj5eVeSmVcVT7ZGQQhNScAP2
F8YBQ880uiggsBgorS6sNiiIZWauU+SbnRilS1E9bvg7JIO32ugGWKBKWbgNL3Xk
T/00y9KnOBkqegUzxLaRxyUbjCseCVcMGb9CiD8m/UsIXvOvvPcHO6kiZcynqcIq
I5rZ+z/zliRwYstiQ2TiyZnP96hnr4mC3GmWzuPa2cQi6mE0XEo09ioxwzTvhE+u
BPnAFL+eGAWNcePy4GFrSAAX7NGjiP0lXxg+6ZD4HxFx2ONhAlQiq9CYgRkegick
SyPNkE3Euf58ndq18G6I8Wxis6T7NR1VWBehmXuccNu1Pt2eaK13fchh/KqA2G3i
FigGKqhbID6mnGuaQn1A8dW68r53JlAtLsgLwsCWPHbCjHxkrt/fFupCPkiftFo2
WBRQGhhWURGmb1L0zT0d8cj22gsy+p2lrp7v9Mf9Hs65mnZdZEeUxqggWvqPm71T
5O2+sbJD+TqpI6sozrurnFe6gUNAv6QAuqW9vS8DZbzTD/dAaK20jsjWzIvCakJG
bk3XbcUrSJPTDt6Qp1JZV8txjs3LST4cP0BW/rpNFH236L6D5al3Oi/bh0M3uXdo
gf8U5a0y3CyIRkMU9mMtD1rVFQiQENyGgo/XkeBSbYNNpp1ejVcj+21fUdj1ya6D
/W8f7e1dk3YAxMXOAA7EibUVPSpOCF1lt4xwTJZw2pavJzuzXu690MoqSvyCxhDZ
fj6/JzXY5w1Xx+ar7WaLdNGd01PVJzmzlUOuq8J3aNvamhvJEce5VqneU9VPtkRP
1d7bOnatyPh6waRb/8fX2k/bNkSsq9CGTAVSkw9kdAf54NOag5hNqbjG1nsd/FOH
5nDm7HD6E4roMcQm6z2WJjq3GpjCDkYtz0vSIcLaoYPQ7PamQbxiGO+itVB4G9Jg
CFRTtcrPzq3bOUibZ1IHKWEXdKEiPl54iv3lMMfaNvj5cNo3P4nHxmT7UNZ8U9kg
4zKleZbJY8ReBN8agfQx8180m0DM+3DqNWSWe45O7zrmv+aDML6o/Q0h4VGgP2eL
v5vJg46f+cEi5GgaRLMNHInH/USsCa4DrSAGkOLsF+4vhVBYaPKS3TcD+RztPyXK
vHT8niPQ/LphXQK2ahJscSKRiX4+HBiDjyqiMV/7hAZ7pX/mj99R5hVWdhcfV1z+
dGGn7naOAo1wVXHkKIh4V5ym9CVpSMZvw9LTduwGXbPwAYyrvplsUXCk0FQSvErR
9AFXkAxJlsaFP4yzQekSgV6F8cQff5e8nIdYh2lJAJsITuvBtY4oiclb+jMLhUy4
uv7iHxwgN1aTvYtPdaPGWAl2wkV09socMrnqhbqRt9d4Icf6SUWxBDiU0VL62Lht
f8BEDZn7/VMEmKiad0bHiQwt2uSUPgIawk5DgP+FnIJ63jrf+VGhZeBgT6jJBIOl
ItKXV0uF9qSP+6aogOhWwEqSCyyIkG2y31vy70bKMWxm/TAn3mqEZ0fFdcgClWw8
+NSVRhLkC0zIItVn7n2rU60ofawMqBVFzusH5Tay+371PPVpVc0wWfoIEdLXb4HO
MX6Wu4ML5Qioo4HfVgYIkyUsPEYC3LLEHGkPZ4jckUByfwNwIG5lDPs/GX81iLdj
s9AeHQyEr2N+V25l7RMjK6AMgT1Pi/GYrI/Kby7iGjc+E1Sd+t8+YlrgtfVwg4XL
28HJW7FYEkncGp+mrCAO2RJE5QKPNVuH9puz6vHR5lqy13Ot7xsCj1dPAWgY4qGc
yPcfKC+AZRUcQ00EPE/GSOKliAwD8VcN5DC0ltvLGeHI06EcoGPdZy78FRlpTNql
t8EVjlVMZ+vek92vX884ZBJhI+TtJWVg3ivhAXkcaX+jYygcwlT0HeVejyuLNrzS
U0LW+yXKf8swCsDNPjI1YVsIXp1jIHhK19GalX6lqHH77Jo+mQ4hlqxbJ1EoTb5y
33aoMTZASdlq9Zy/XSyT+ekTWOUwOEnXY/0rdbwFf9146TidCA4zajHw+Wu5vxmU
B2TcgofddJELfnxzS4OnhZF0LbXb2C5BUgnyNw+oqoc0DeHyBbcXErsdTOmqsw2U
dy/+i7/H0uC7+cmjityXdSmmAMCcQoNgImkmjU3OxGULtzPXjXd6g4eYKVo1OmUm
YrN1seK3e4uwgKJ22t5fOAb+aaG+MFWBY3ycwkpgx/QO94LE5iYknd/3vGZl7vTL
iMgAmSNJeaD23DHrQkiLTVN5fQbkP0Jhjc1bIGO81UoAj+nszFsKad+61WJsG6SR
2jFDJMqHFSg7W6ZaOoJbvmO4jF5ajD6UOCv2pX+AiN6Zg2kyB2dkvOxrcfdTLbHs
YIo0JfrVkbRg0ykIWE8OczMy5Tf3FqX+PNPPgaokuM9DkpMfOOZ+P14sXRFMIKt5
rsifC1JdD/EfBhz0G1bxMKl14n+XzFmUi2UvjJvqbuOPJZHWKJd5ADSqU7JD5uCJ
2mLkb/xVvSlo1PV1MS6EGSVMSWsXnKaXqgRth3PsvtAU9aTskoj9UTiSKo+HF9zW
DbtqRvnyZPFDG2v+6CANjSjb8QHOWihmuOzk3m2yYAyZTBH0dPb25FRdlD9MDiue
lqTjB0OWdYTMEZ5LLY4Bw3aWf55MdUcc/dpfBkyLh1/12h6EI9uMUsONsXOGhu2D
ReC40SN/aJ9T1TpxsA0IIYTuiUjCfxMzbVoSe6DEhOGK+OYv7o/gwpNq+FBU81qq
bSJAkGK7z2+HjWRnmqFwQxmB5lW52s7608aE3geN3WXyAlhB+nRGeO9TiyRZwA05
M/mIHN0Buj/ZXlPosp0jJ3jI4/QYjfKB7qw+wl/JON7hEceZlcad2OPfUG5LTMdo
2VyGnsdFZXYyeqLuxNHuW3vi5O3gpWqQQ5FRn9YCDUsZAc8pgIPN1Iq9iY/uOFXP
a71h7D94ZBQSXJvSeb4Cj0wVlRsPfcEzwssGEusx8HnLjgDToBjnW+XElxB6tiiz
yDSrCllAgKpO0SzIVM8t7O9DIsItSUWTP6ObjMn7OugjjaGrf/8/r+FH5/ubfOVe
qEOBzVnX7qq83W/iZ6G/jBo/OzuAVPdsJKIULVqpA8hsis5ReTfIeL9rTkFeqWA9
1B2eiEq3ECLdSpnfH85lbmEYPjgTp137sFIY9aTJ24kWn+RlqIw3hFZ8H73J5xjX
XT22yCQYdp1Tl1vMAGC/ryFwu8MVQ/v07Dnosa1rgILJawrIiDbne4wWnXmF7429
3YzENBh8MozPzFEnZPL3Go+aoWXnNfhIwCuuX2GcKUMQWQi8kp9kEVxZG5/cIl7z
6AEwUPiZlWVInFJl5q7U626MHox9NKmM7ad2rg8/mgnoZhq49B22dE/DRfXw5w4i
rFyqtBjM0nbgLeEJP19Il0uQzRJJ/Tw82q4uobh/T7/7/F8c4fvP2ivyu6zCA6fF
AxU3oI7C2hF9gLOdImrH8cvHsZb6EVsAfEXMP1xhknfjc4IfMIa/pgRcX0oPBM9o
eP/dyjfRKed/JZE22kGngEn2UBUaRx1PCFZDmqLgR8vbZpa3CZi/fxJko+U+hPth
hGoltFetoEfUyO/CU0KBgzaDt51fvnNGHvsbpMvyeDtJeUprnxeiLNRfJaHQMGOt
ENG+ivXeHOZ35sfPusYUDG/CC8RdSz/SGoYCtvHyXDNKy77/jc70NICizLwZ5Zgj
csahevuDFYD95Hxd/RcN871Y652nQeXi8nXTpFUCfn44J4wp+vrpLalJyMb+xyi9
zSImSqw/MafueKxlfOOy2qpbIz4TISV7jLlGaOH5ixz0kDCtai3F0DkSHB9fyEP8
SSKERFp+IknfU9heDv3QP8eRzSaTshjxCK2qsOaObrOo8EFR8NXhsmRnffb4hidK
F6kTNI+DDE57I3qhW6atOqHGBnz6/7TisTik3oyKaGOrQWcaXAvd6xaGmjLWaqz3
zbyOTUsbjwVu+Mv9UuiH/VjSeTg6NL9oPD8P4d8mB3RPj0B+f5sBqfoP/dyrvhIY
c1I+QOcyXtwdSzI+doAJiT9+A5Il8PFUbMSuIqlZUylW61Xs54aW88g+/djKLszZ
FXO+y5d/hj2j91LP+T7yR2FE/NpaEnysJr/fkWGHxT3/xUPdUYlFVObC/8DFAZvy
LJ7lPg6tSJKOOpowccDlvHTewFyuPmslBtt4Rq2y96SnTTrXG0bsHVoAH7fjtaqD
Ju6qXR62wJrXQKgjHHE23sLpV9VXXyJXp9MP+sTNamh6bXGN6cIIOEPJU5/BnMRh
hGRsOnbGikLgKYGloaNj/kZrY5Btd/VDna2WI5x9LUetDnQSKUBu6uYAdU+NNwUs
iUYnVK3p6n4HuIfjB94TkR2tF61XtM9DbZ+W/MrZMYdHoievH4yRN5Zd5aDzGxEd
OPhqEK8Y5yhE/iezpbl0I25Gbo+OKcCX0aw6UytfnF/u2Lre+7oOLHpUjqRtomYQ
TiGo0NchzDMEg94buijcscdUeHjIie/Nd7LTAtSqzu8u53YQwYT6Md4DqS3sUcuG
KNkeblhbU3ghrfah36bv2kodj2vKD/wmwZNVqL+DZyikNttWEFbyajx2IWF18k/i
nQqH3OXMMAJd/TcttGgC0PaVLVNWb27EA/x7h+frj58h2cfTRfKUGhPWeRvHKcTP
Ei00IhZBqiQa/xTQKhGwfadKndacPTz4sSVyJBoR1bf0r5lhZg1uMvaGR81GsY8O
wNx6yIvG9iHgbR9cYiZS23BtHiIf7sek9KOGjNqSh0onag+G87LS1tH31ad1tDpc
gZNlknTZQTDnXtnRp+fuhcjWj9OaS79Gn9RxcC44eIT/GHdoD+uI/uTpQ8X5HYcc
NNfsFedGbzTflsp3psmiS6iBBkgXY5rYX/nfJCrFtAhAyB3IxzmGv0XnN62EAjwj
0LqPD5B09HUW1mDbE6bghMmn+wPR8aejUZ6L9AcQMntyif0VKROZCi71ELNCT6TV
GWS+m62x0XvIMtp/NJz3/1Zv1k/hbPmbY6QGZB8Iaubu+EPipsm25s7/1p8OZ09Z
As2OGlOIzOvi8J3EMwKHcU6toEt4M8FzIuGQE2PNGsv1SX3v9Mmq/+oJBpPkhuc5
iaPqDfM4zudddQlYvwhtWK8olJqRbtaG+bFYxLwbXDdFwDKAqPlqVxnACgOIXE/W
TnLQmdrAF0smMDSOqrF3fjpGAhPFUhb2Y04/+Myd1PioYtJG7gMP1DFV8Tokgy5/
6cVckhsFUfUtKiWF1iK+efEk93MgLDe+wcopfULluFxvrK2NKNHJWopaPNKI98RL
oqcXFJMeBCq4QUoFGHBYyWg/b6QSqgmIWUkuqwMtdZ73uBK1pKB0tOZwZJ402yA7
edQ/yI14gLOWfYMaTvaj+Tu25XrGmLKy7JmyJDGTi1fpi6IfsgT0QVtqGHr9UfJC
+rL87gL7k5qkOapEpp3sB7iw3KEwofu2SSxPEn8iOOZFSwDJriQAgXAJtwL9eWTw
X6f6ob8RoKlmYyvw5BDWKYRa8MAjIDFmADILf1QCBU+FiMzvRhEGuIdIFkuIMXRm
6UPZ3AvppSQ+dT+84Rtw46uUGptLpmsyEXSPPSbdZP42FM0PtE0/1M/yG9GsuUlR
CHiEBw1uPRYjqy22W58K+3qfSr3TFciqVuqZLLitBvVuPUnybBGSQTj8ZH0RnIO2
po/LIXfYATrMTKtwyBwD0M3azHRReWVn6WWgJsBte//NRG5185l0vJbIEwAW+5LF
xvQI7JG4weveNX/F1kr9e+CjfcB8J5aQFO5Zv74xEHLgSunBKkcji4gTVZdnIKi0
hVWyqIovbwmpcamNF0Mdqe9pB+XzKRj/lFUGQYng1StLjj4QT3RENMzhpLrPDbYy
lWjFowpBtbVnsW9hJIPog9kHsO9UbtzOy8ZPlJiRGtJ9nm+xd+lJMlcK6ddH0Zoq
`pragma protect end_protected
