// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PRVW2T4z3RMWajaIhWdj2p7j5qBVlM3E+SknGLvg+GxvFNJ82wzP21sZ5ezJUmIu
eDGDyayqLbc/G1GdHhhpvVhThtGkmESGuNcyW6yuLntEmmkn8SJwvLVkuJCLaBtb
iEa9oCQzFhJ3bzLPGocZafJhbLcRI8cny4Bi4oWcDh4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8240)
yBNVNZ7k2ABFQz4zpQsV+N9Qb4ysSdbeHMg/fxjHrmdQCCEyV/TPO3kd9s/+d/Pn
k1xNG16VX9P7gZxFI+kw6cGWhdavdAjiYm0eKjeAnx6uBkucLq36zm8ex0b/DdBc
4OSBOFW0u5bYOaStMucudNhLttzXZnyr1Vlq+4jBXaKdyX8uZs9yqS0zwNb45Vsj
ObWkauENRLO5/MSEGIHBO3d6hAW/sjfVQ6faZiB83ne/Mt/RD4eEfhK91MTB/ATM
qqXWlidqQ3oi4e/3Jlkl17JNRcSLH2T+6jP80BQ8gfYQ0WD/LOrqmIwv8FclU3u2
YoXAw0JpZ2IGTpARq/eOm+zN1IBHyL1jWHxMAZ/9Np9rets9jG72Gg64IsQQmaCi
TsGwYUeKNcuFHaNnu4hq9YGnkEczFosDuHP9ZOiYjELPihBXM6twB3zvME2453uj
lAFftGGAgjc0gnXQRHGNkJdZEchFrYHr0UE4gCqtyOOPsUK1TIWg+raitAPZm7pK
oCmKxydganO+NKVS92MJRxquWEgUob3v15ZQd3oA3GDRjrusw0RuIgFoKhGr/vx+
Z+OPd/zSw5QVBfqOcL7YptF3z+VZuOoj46Uis7BEy4BA3rwEJp3yOcn05aw7cPBl
z+0vxsFsjM8LmQW/NA669hLiOZOitfIV8fiHNRCKwZqRjqGWljIAmuSB0ReMwdb8
xTOF8GZjrjKwOSJzgJiqGNrarkGthmMEhQDZK8zAgS7wP0gzLEPI6nCe2BDiOJi6
+Vrqfg6og3qpIaSKUYMDIFIFHLCfRFeuJuIF3Mc6yppPuFfvS5j5TrSkSKV/ISjQ
G1/Tllc46dkM1IfUeMXdA7f02DiR9bKZIJy53kuGmzE0agPhwtNQxD74ehiAjZIU
VSiiD0Ef3H9vFti+WRir/xm2AMH7PHPghEvS1z5zURyNkbWs8kkU+gZ+FuOuk7qH
+HoKfoiH3xZoZtXHIqwOHTIYMc4AJOh1wpdjP8MyEK7b4FFaJDdEY05TCKEnAPLM
jiVr+b3VUPjW4ck5h+24Mf167/B2gt7CBNhZQeQIqKvN0wLLn1QZri+kxbEh3jYp
QM1qKyJa3A9w3rRus6+Tj/Sj5KTB7j9hhWLFq8wstI1Wo2VsJ3J2ITJ3iishGkRg
wy9di+vuaQgZWTsxn/kdv+k74Kq/o3l2eVTAxQTJsHuG8rNcFKuiNkPS/3Mp9q22
LHa81IClIZdXt85XGu8u98ymYJvNiWlwAzgpENT6aiPJhK7WUceRSL0NHN7/vNjM
teTAQTrNXgoCBNfYgLDWkV92sMouxANDbr9J530xPf+HvqTuX0jVixAXrdvZOOAi
aTm2MCKjkhdp636VKHLx1DIq0JRaeOxJsCfRCCWQTWo7MJP2v8ZpIAfxaWD//SZT
L5/sDk4W3HI0jgrqZ+EAM/gxr8t4GIC0ZD6wwQiaGIGvcdURrHxRlPlhObza4CpC
ghLs2gjIJNpqtgF88wLa0ZMLh6wW5KSDyYw+pvXZIRjs2zXPeuGNmgjZg0zO+gNC
CBs936RN1eyMWOLpiL0eIW883XmDgCWbp7kk2q/VkWzxPeftnKFf6SXiID3JUOac
q71Yy3dT5pikxiEbJO0FRIQcfiwO0jH79nJoBcpGt1dHbkpMUjzzwxQVKE4J7PAP
CNDhQB3YziGRSLTRbZnZb+N+JDOHxWB2LmPLsfiIbfEZbUOk+pghBwV6NxR17ME4
P+y6jNtHdVKTJOx51jkG4Iep68ToUt5LIXX9ubIe/tT+1jba/315IaV+B3mOXIf5
i97bIKwtTlrtJdRJDKezuc76Ny4s+ifdaEwvltbsf9n32ZOxXHlvrC23m6GTimgq
I14zgTsj01IAQqzU7FkMTA50oOS5iMzYjY4cfcLTNBDTrlOQT1cNVYDjZuq6Hlgd
UfJ9+Iah09/3Si9kc13IpNzpD0zwTYVzm1kZ/lcMPYdm3/+PSx79T80iRMwTi6aV
46xh5JCpyIBJ47GLtI18d23wR2B6PbvIMc0VE6Canoz7vgNfXay2Eia5bMoHZ0HH
cwt54ZeN08mP95rDFw8AhwR6SpnQuvYQSXif9ItGjEorhT2/cStDowLXQ1YWMayV
GEWsJcfss+jtHKh5p26UqrSbrrRoF8kaKFEWKVRT9B1C5zdeC7KhfxWosiEKxl7p
+yrv/xhv7t4yT4GJq0LGQjjeHxLGXE/je300CBFgqb/CgdYS+jG8bDAJrq3xkdgq
ywNc2ng5gnU59rACeYqViH6ynCRGQhYO1TVnoqIji0eVsGXbeBwQrebAzwEhmE+x
awrwOC9mw4P2KsyrP7kgMg2zQebYOs4nL4TpB1WdbfUqmWS6MT9rRJuWrspYrCfx
TQKMO9+WyCteEp2L0QOdHP8OlgCVQY210Jf9Sv+ixdP+R/hIDowT4i9f9a390tP2
XkBVyOPCyFtKkVIxOaUupjkCsCmVMzmMpJ6jnFrrjAL5oZ54akUCxyj0hWkOb7aa
M8Y7m02S92cw7qvkEQgUax4jHtO5tZgpZ0/uHmIr46gORcB0CypGr0M0315+hO+N
cUFmBfNypn8Snl6Yo1uH1DS005EVH/WdUYt7DP1+asqiCAOjPpfCwAxRXTWROzOp
deczWfK5OslXs4jV7aSFGATxcLiHDapjOsUwbHCO1o8838qG3HWABI0DK+vRcCGA
0/QSIWddWLhyDN1r49nOs9+cxKGlzst6PgBZOIime8r6YkQ+GIvWQzAYbgUUoctJ
wrULXaJbILlQIFNwpLBxLGQVaD5kF8auSOytfN1CMcxQmuudlLsHh7kO6Eyekdb3
Xsy9kNZ2U8OHC+wEdFkwI5r7gXXu3ObrgTmBHhFeZgBxSKH9uM8qM1hlGBlMpCGL
/i4jaD+bT8gdfYcwyRwbtBY0/Hptw1zz7fKJvn0LI5VXbQLWO4cCU1y20V4qKQ0n
QqXLUdbKtamzWOAYmR3xQ3OPM92SUBj02vcGNHq+JIWG3xFcBoM3zNhOPvuoAWTS
43xQPFb29k62OuUDFPIg/G3muuVTwd6Tl8l0G/WvCNtw1PIynA2qB8kUnIkytyu+
JkLzVtMLRDyH7V4MPhpBte1kvros6Tvg5+qc1RoQW6LkC1V9ROQWLTmTg8ZWvFQU
VEz3QhUmxNd6bv7RXea08i33ZXTCUcVBiBeerwNwo7njACRgv3FPGXROPTUx7FOy
3zwnvxWbNO3sreZZxwwdkbWNZ+zNunvaSSvqYVe7YmW2eYGrqXJteuWfFtdn9ALa
5LcQiK2RM9u3ZZwCfaUEq+f2QYtsI+xeUjuhucDQKdzBl2Pc3Jd5In9Sr0cDMt8t
+nObOTZ0BwLi1GU9Hw80IpwzT4qCym6Fopjz/VW6rl0tPG/dNEzlVAVjGfM2trs8
PG7JMuCCu53U3POvr1kiUsa9nrfCQRW3LsndIgWy08ofPgw9TPwEzGL07TCkhhRR
+mashKPUE/famYX+hZ1EAXrbzxO/iOtOuBtnoaupBuYodcKQvminFeNEt89ezECr
COUbUDVlrbLsc7QjuNumnoJ1+R7fj6PFpjYQ9V4hVnzoOLZ+ZnDQ/gRem0yzb4US
dV8yQGs+C5in1QRmH9Iqibcd0OvBI2VMaUcU2XDvRT/93zkOt/mr6Gs0sLCNBWKA
KJU+htV6+noUpu53Xs/VDt1I3D5sz0uhHqmQOna1J8OQCqQZeNKtNU49RBiTqtgZ
D3UPHTQTkeE/nzqu63/lXIvWtlTq3CQfu/fKQJxTqKoqE3NMCSfnD6C4CLs490s1
JXDjB4Y+uKW4lda2DncxSkf9VBhy5CCPH4O/2mcQyXQ61hpTsjSCdYujkGLYwCNE
0OMsSqO14OwoHFSs7W7PY7yYzUiuseeezIcmxX3ukaByisS9HDKWNh2QElQYOR60
GkFYcU/ztCOSX2CCsNTPXODmSNa2NHDm1jXLJp5V2e+U+fDqUn9in1VmZmqYJ1vo
QEEP+lU7C6KELs7GPPGZe5d5wlLf69XiE9VrLZkrEYb43NF8+uZaCLBm4QZX9CC6
37uo+olLROsV1HzVBe7/h8uSnh1EMIXXF5XJ2xArsARx0Z0gGl5mMUlXNNcfkxs3
u1irUSuzpak6aYASvgD2h7xzp6xRGH3XudFgPR3Atwxpr5TeUQnDhq7eJyAWSeFm
u6a3mfPxm2d4uFntRHvhn72JZcnCuw//fCWBhbAD1L0OAmCNcwWeyF77P0Y7Q8EK
FTXQjXJd3QR8S+nTw2/JoVigQhdi06TDIw/e0nfCmOTrJ+FbW/WKfYKRjATcON4J
Kfuq246fgYkgpvSKAS3c9IaPryV2nXqyhxlSO/EWbnQF/i3KvTaCWe7P14mX61tW
/tMsC8zBhIPNgfePLmYuINh36x8aYLYFGhwrePvBu6va/JgabfsdV+pIcdTAx3RR
Mrc8OGZLswsofGbaH5wN4d2NpJvME6i9SAOOKPZjg3C1H4R+EePjyfuEU8OR/HQM
jE8+cyGAtzmhYaB+GHzrtu8prYL6axD86RiQKZE0IbENcR16vuFEJTaqu/zsQ23S
nNLQCVjG7YFewclRtYcIRzmZLhWAxvGZtgq18oWne12hzrgkAb78cQNAbKU6hbbz
yas63tmKKV7TZ8nKMnJjwPa3z8QKT/dVcryXOXfaLU3vDoUp69JOudqOhYWVJgCt
km4Za34PcYABeuOvRygjLTQN+qjkWncXsEAYdt7fAfVECYELhcSNhvhxlyUqQ9Ud
o8VByVaAClp9xcq6gaIR8zofqWC7J9JuRkQ+gGhBjUocsFxpeo1rQiA6LbNcjKo8
S/gT473IA2z3CGNPagduVKIerQiIt3B4Lmcj+75y6qBjvrouBtLa80T04YRm+r1Y
bCfZLUtK+xioF7/43/gd+WeYRCKbebDWMesqFzz2NtHmMVrrzOUb6k9OI7ctUC+O
VXpcLHUlXwOB55OFG5kEywm72kM09D3e+peZvGJqRieduNo4+Z5ODkUXgq78h/jC
raT+O1OMrWm9f/ml5E2uNwjAaH+urzwHQ8fvNoNxc1UFNHwvn0sNdBGopNTHLs/M
xolCWWCt0UQe66o73RWNUPY/MDkZi5tpvuBBp/VydS97b6q5nXPjJ37rJJEfKizK
VlLe5TKwchEO0mprfmWg1EBVHVSX7piwcUS/NNVMb3fwhwq15NZwDlISX5HYbcZS
VjOqGUfOY4s1g0ghCsWGwI0SoXiVfcfq3XzXn9y2lRZM5VyR6jiPuy+7nez07Csu
4MYluqPdyxE5nrCPWzt+E9lqxTnfj01xELVK37yPOk2xxWm+6+5N6/+yXcTiRHdr
yOLV9zslUoG5Y2t2n0ShAjiOC5Dk/vAOeV4B6n5vRlbIBuNJwLhd9jY2YcCshgMV
QKr3CAb4df7NN+OVDw/mhtOPIcuufoOwayYDWpK0Q0YzKt3bnpeeIDkxF+HpJMNk
2gthm5O5gDQj8Jha5tX5uebBhGFNKv7/ixxpwbtqtOyttaGybH8dl3friJA/xDt7
PJw2cOn1UcWrA9ynCfUcNUyqasCf6otn10OurhRqUWY3noAqZYjTOhae1vazMFwr
O/a0OOSc7JGRmMzWdGORNzpzqNSQ1O6IMvp9wcDGwtYoS3rcVmbyXozyewEG9T4e
NEzTeN71EqH6vB+Ji1MM/NuIvntVtQGld+YmzG85pu7XQHbEvpNxPuPsTmowZcaZ
oejnG8WrhckKZdJ5rS+x8nuM8iSALbVqHmd60wkeYCcQ1xzf/76FoKkhvMUshnlE
3PA2N1Ho1mFMDbIWPYHjo8d+UzlmYjAqCrWhCE0S78WoqA0FnGK+5hLjfLZHOWcl
4WeoS0CZRDi7gqUSV6dd/mPsmNrrmAOppY3YAOxcGwoxKEjis2y5J7N5IcgkTWN2
RzIwJvc+I3OfGwUC0U7D6LTAtLFZTtVHIpayRVbKq1r05x3VdJ0pb0/lsFaiXvms
pSICMACCYdx63tkmjf6avFXs0jeHrjfDYJoBtyqfUIwWJ5cRHwEhXmm/oVHyf//4
tu+22/Q+zwSd0VauWiA16hO2Sjc4S32Pc+24qO+SX3YPsUoihMXy5nKRXghhijWa
6Pfjs64rJ1mJwmLurTJLehoQaIRelmK/W1pOPDosZUKyIWTH+ao6Nzy1jFCtQZYn
X2gKmZm85jcgVkaJBLNxBbs78UwZ2ridDaNfUyHZngrzlbGjdLpIQ24hzX+gll6B
E9IaLPRVBxOALiOjf0ynyzZqe+vUZj0qlvedq++8HMX1hVScsErgRR+ZQorMrWv8
OIz168ojHZpAsQtAoftoRq4o8alYxYQKcufGtp+4F/KhWe2SizhbmJ0LbYZpQIks
m8nnc+VRXf3pbyBHzBq/FtxVeXjbODdytoKEgkWK/36s1RSlzrY/A2XlIjohe/S6
kcbUuTNm2i1YLM/e+T27NoQwo6ftp4DthVlle9gLK5OKmRwHLgqNkbQXzQ3mpiex
NzKMG8exrJbeDkNaqVMB3qUoKMULyKSEkCj9sBMuTJ4AvayW7x4hGZkf8NTnNfv2
oz+iKjed6SGQs8zyyxK/Bqte6KDIdIfjnxLDva2YLZmp3jKcnWs4Ucr+DpcDRfcH
vKj8o/QlskUcec/j5FKLX2IVf5VfDn5kVibng7IR9dEYHvLBU1NBJ4gfJG1sXvI/
pUGYp8l6V/UdWsn5clZIfvYhHd9BjOyy+nF0YPNsBcqywJtxZeOEleFemf9Zs3kq
D0fQRVaxQv7MmyuEm67EyUPfZ2xEjlT0me1yl0hcmZ544oV31Ube6uP89JG36K/Y
NcmBFPJQUElcSCVDfMV6h8jjI/ynExm0Ayz4HB+2zrH2T3OhlGQf0S1hclQUK+My
XHfkCWf6gU0uL/VbvvAuYblboLO4FnceER4f17iTvrZnksihqKHhrq86BXS7JEBP
2wXDtwvBENoX1EEWotHzhpHcwuLK9fp60Z//lq40KXYqyPRRy5Ie4gVEuOygG5LT
Xwcm1dmbCZsXzXSJ+sdqkDhUwRgVYHZp4+bkf71CGYo6tdDNEGl+S7l+kb8fGPFQ
f6fWk3MIKggTe583MVlOGEJWTTq/yMAjcI5XAxx7SeoMGu1qpzTF6NJ99rjZYF4h
3T4keX/6zpPLE/2cG1Vr3KWXYF7+yJEFZLkexSaRKqwMNyCUIXtf1KbGGkrrSz6/
shBqr5vFUuFzgmU+1zhZJEdGy5qB3r+WsOxXTtNtV34vCtJJjkYxDcoFx4yxyIgK
wyi/cHNzW7Arig3nB/ZE06WUSHvQ+p69JLVDySsrZSflTYLTzXFuekDywgIM+Mdx
cBLyqy3CTGeIzY1vdrJGiCpr1wZrkEH7v89Exl7hcIQh0VqXPzBBGIHzdjzLW90U
NElHWfVKujgDUvNvOAjNWyiN76fsgGr/UZcRL4iSW60Nt0CJFiVofCBHOofDxSFI
/piiDrRGjGMFB7cajK+KZgnoP6pcA4RREcGIq6bgObnGy5JbTd8JGkEX/rvD1jSl
QbBJIHtQTP3YyD9HH/4a0TFfFnuhUDbDJ+K9gfh/YN0gL7Xz4rQPaSwc2RUzUiJd
VOH6sHpH1MbX8JByY3GQME5+LMIolpF2NBOn9m2SzbG6i5BzCkI9FJnCjd47QIJt
3iY2lb/aSFFZ2AEdl/McaC+Yx44fDwWfbJwtOPTu0yOMpQEALre0MGJlmd2wg4x1
5WghrdgtNTEESN5JlHWsOSAPI3j1hknTxy8deCL/Pvi0DaB/U3nAho8ZGxMQLigV
DfDKWb5WBjC6Ls3H6r410/LcCl0qb88dTV5Gl/2y/+MHB48FKTXgWbyGgVgurjE/
qi1gcHWbq7WvlPcA/0Lg35DiusoWTIAcGRouHmEmME2IfZzwZowLWyFhukzgaxwR
uuL6daiozQwjUl/XH9URQOgVDl48EpC53NbtYIwWWDo8nyFO3iszod9GYtFS077O
xer7gdKPlaoJ3uQJazxcOVkQub0M+3U3H7r7RrrFLT9hG5VSm2Po+Vy3MQwPsCu+
hf60CignU2iNM2TSvi0FRieZF4AyRTdyUDHfSqNOAMqRxM3QOLV0cWcbJgtheci/
H021lQs4rwiWBV4gT/BUdpUeB+Qv9Qkx1PvVztmQda39y2xPKbZ9hG0kwruwUjR/
xgaor7cVngzcmonpQZHcpm1mC2Rt3ykdDmtt6KFlKioMrUsXD8KV8UJCqh2v3xVI
GO2dMUgyTircAIY+smMjAE1TKCKXou1wLAg7Wv8khTd1eLGsjWdIRnxisAOIz7Vi
g4CC5T6DQG4lT01NqOtPOJfpJBDrwH9UFPIn297swfc5JkqaVeS2eHePNLz+m9XB
tVXDmP+OQ+vIPugJ9Z6nAkwejgqtJmn4MC9L8Ry9yky4bUrYkLjoUjC8HmpW5hU2
pC4mRnsfNBpcElIP32W/ITHx28gDQsOUNiCZQ9UBz23DHqkRx2HtdB+eQ/vBweRS
nH+92iMRrnYSkA+/i7Bca9VI9tm0xSq7Y0wa7PCK74yM9TDy/sPkCy+z36N6odjR
GCKvKCg1mQT1wM8l+v6hyzplg9tjdG2qKBNGVF3qvqVfAIkf2oTVfhgMhs9Ttkzn
nPouNTW6skQJqKNtHs/MRzDAPv6ljLtNmf2HgJfsevUTxcSjRwfeHNy2w/b1OLCW
CcTscWQ/k/AYLnK68dFtQgTrxPjOEfOLf4HE+tgMu5bQk8w7yokyjyy0BIizC3DM
iTLmTaQWaliOAkmqCkI6EQb7hGe8xXg6FEgc1rHoCILHkeQ0eLKA1MCVOOtHlVqi
+UcqjWInixI3uJbPkIl1J+NJXVmOdK/272b5APRfprD9nhpBzwWWot0dsXSskFhi
hmhfY1LoXe8QCAyYHDHJVDhXFgwKHfHmUXKECiUi9wPQGfsx850fHKfIjD2ckh3D
Z0GgiU+F/nEek7KbxZh531a6IEMq8enH0sfIVl/tareXtKDPomv37GjzCjjsK2ny
BGMdqVdOsqilIraEz/w9zC+TEG8w77wYYcRKsygd8U26C36jy2+CJUtBMp3qAjbU
gNN0dVYfvuH123t8LUkQAfyF6fXH5J0igZvjkOlunA4ox16vxqpOi/CmvPZaLWtd
EQAo3RnHqN0X9aZeYzGXOks0h/KxrUNm0lUiOVpD9S3Z6ZUXv8g6OYC3Gyxu6BQO
UHobSke+rI1WsKGFDXHalfGl5QRBw8pVW2AaCBi6u3nNxrFAOwndgiTLX6QXqTjS
Gr39UZWvRS4zuvXLDADmCQtf+R9jAeFRqMLgSd50CIwg4PDIGpM9OGQT7aw5PMbr
DdAFqOnKU6aBEtR/JmhO+ONje+Px8jnKX2FUEcCovMRVkCMXippQIvN73WKHmSwO
X4ZH6kpKLdfv//5IWBnn4KyWd8R2skvckH4o+eHRiBXuH+It+WXZLCTslqD/zQ/C
2j1rBfRtDqCbgZVvG1ZFvk9fKEctD5Tr6v9lnxTXE8n1ATq/TyDeIogb3AmoloPi
/mlRf+DljwuhRYfoxGmJzeG4a///ZYhvi4k/un5la/aAavoUrL83iLo+9wztDshu
E0lVvFP2BZdpcvO1+dkpRZ1+JLRo2zofMLFXIanRp5QmMQ2ITBha/ZZOMYY/Aej/
cU7zy7c/kr9gq9hy6i2fLbGcuTD8EGWByil6eBY1wqYUnjxN8ket1NK46L+Xm2Tx
AFQOknkWUzgfrXGFeyc3BmI4OoqVMwzIHUoGrkUyomxtuee7T53u0TQ03B7NnA2r
TDP32I5GbppNV9aJ2wG06ycnQiI5G1N9DHF83L6ndivWoNSK4F//+nkmTfD96wh+
A3riuyurNAx5yBKtWv8uU7ymlWJ4CfgpR+Va1LO/1b4nezVsads+LYbCFQ0DQsIP
DgvHO8WgRZ8d9xKqURx1CETSf5ogtp7+B4FTSdDWQLRQ9iff3J+ad2HVEFJsxDWJ
Mnnx4nyDphV8vzGdDTzz7d6M15lguwi6dsved76EYThkc5KxnNA/sHKBV2xSJL6s
6JtFca3/AQjGuHhBTbfXGqjMmKL8r6V8KbAxThzryI14sORvpcwpn3SMSJPthmBU
5KnHv3wltF2Q6CGF/8DsHpA6k32xFNyjzPNlklAeFRfcXMVBfESGfYjeYKiFNzaK
l7Zm2APxZw+v2LfFYFRoyYG7d9Dmk9XWVG1/TObQNuDaEpK2nlVLmG7Y1eGkkhwZ
2Ncox/7jNj7DB/h2w19nNCcyTMXQxxR7pMRqA218LtrX+BFUViv52xtFej3nwozp
gR/+fdJs3hmCjKsgvLEU8c5ZKAcgUnT8ybOT9lyXOqA07ca/DLWRioK4s/TNILFA
meSUi7tBZNt0+1hhElzAGZYmOdlwk3mqnz7zLanC30V4ZGtyi0qftqmpwwkLfgwy
y4bleZ+vXry2r7mZcGJMkL2VSyfHbRbmMfhxJ5Yn3gQk69XyW3dZEwzZ/TjihYrc
GKfLDdA4E3qw0jVI0omHsXHJJR4vW4l3k6xymvH2hp6HBJAIyEe+iz06b+aV0+ik
4X1PhLcddhr7jj7spyXvulxzHxnlvN7tGgfs61EE1EN9IJBlQ3auXPU+xhF3PzIV
NmShLOYp0pa/vYGWhbmcFrLkX9Qp4OmYmqWQ0W7mGfAcET4oJOmUmMwXUeyDzJfL
wvoWvYnaLM52aoU2LIqHpRxj4UliHwn5iKgnzEGtiC4+EPqZbaJW7tl+yMpSo83S
E53d1ga72z4Fwlqk8MUoRVMtht3L+LRyR7aePpAz0gClvUllW8eK4q1p30gN3o6o
yXNYgqzWNBdEEwZai8Jatf96+KGfP6VjEeqNORvn6Rd0Zsu6q7ohsmcjFaIOClv/
UfvrOvWRuU3cpnoAlenVpcYjML1W8lNmoVyJnLdBdjhwrw/gnuTFSeJ+o/0zbMs5
0/AOnNhIimSjv6gd1+jH98o96fWmdttzUYCl2M1FEBUn6Gb0VVjdsky0JvGqgys+
BU2eezmAI/mq1tPT0fteoMrQu3LgfiH76uyuWWbBqsU=
`pragma protect end_protected
