// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PAbrHXUd0jA7B3FjnPZjDh79O8wxQFRBslJL+muL3uOXH4wHtFn4Z8hGfaLLuFOz
p/muUh3wVL0wsUKYU7F/3+beVL4lUTYdsmJ3d8mGfMvYq+ty/kpMrx7h/AMEQT6+
2ybby3JWOh/Qe02Xc+5zvjbXRBRMlvKz8dIoUy4tnRI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6624)
WwDrimQbFftEk47tB4BIlZpqQic4Gud8egt2zLqq3BmF3r3I/WiG35F0famTc+Bm
dGdGT7pD8XQHbV+nsWudMkLbhRzvveBt+55mv/XXWVEwgxIyATBM8fImodJdcxeS
+o5vRZPtrIoRU90zAoNTQ17MsFoKR7g4XvpNNDjTTN0b3fpuTF/Gb+xopnoSOxoe
XYRgTA7mRlRQ2rvnvxuB5iO0HfNpUsK8LQCNT9kKQ//ikDL1LjKqn+UixoP+3a59
1PNl039YFUA7JkxCenuiQmABJ14gu/ZSx/qymM5ZIiDhvNgZ/Xq5RcQ4R11ygKm9
y7u4nm3g0uRoVUM2aSWLodNUzo97bUha2waLCRJB34WyiODL2FM2UJ+VJcrGEIMg
WsG0ByXGoVdpO6B5LYxpRwp8olpEUzA2c0duIrrXcW1BtqNgEgxpjRcyQsM6PbNw
a0bLbP09PIOqqwFoVw2E4b3zkplhPGZtX9Mix1RDkrVQlr/QT//NgB64h8UoQ3qs
LJfGDul2W+FXc41E7m6WdXjKL3TEpLNEMn0l9JPHxFm9FLFOFHZD/SWtxEVHJZ1p
pTqkFDoty17hHKJLFfQ6V3pfZ7iUgIab7Z0kjanh8siUHdr5kMO6H4aorv9bD4eV
INGVt2LJuJpsZijOidTzdAOH/MtRYUfRmAYdYUeznpx8qwM3FQEHtkO3wfU/brCB
QtyJ4sH4uc9fXvsSiiXXsOf4bvSAnHGSirFtcvZZDXiEXjs9Xxs8Lnv42Abr7OSc
V1s4Vp+ZjBs9t06vny+RVj6YUH6S2HiVkA/oqmkkZvfRoU5uCz0l7YvLfv30M/6M
ktmmyvlJMKy+tFj6AYCWbCTxvTc+H9lW0il7Iyadu3p1wYGa0GY/AppZer8Wm468
HG/wYkVtSorjTSbs0yBl23Cp3MBNAGLwIo51H+dbAIDheph79reH/XcU8WZvoFcb
O4c+CNU6vW6Lx/ZsJTcYzcW1MWus6Kk1h+BIi+UmjQvCgZdJp/O4j/rKsWRHsV9t
Wxde/O57Tvfn8lEt4lt8eUsRoQ16qVLO3lOlfN9MY+tC/oyIMb2RdkSMO4DL/nGg
bY+9gk/1kEqtqze5+n+mODACHr5Fl/FUORiknWBnBzjfTZecNEM29CRsS0Gu7hEy
NpO2L4kJxGmYjVFw1Ie1DwRtrAa2SjOcwLw77o+PjU6PJ21Yf7X3lncZlRI6Q1R5
vBfrYrgZRnsbbuxmO6/iyj4+5l57+l6yjdYYG7vlv5oxboJ/DMkWPSY3RI7eUCJ1
EIufIsfR+7/6ikPNDQEMlr0m7LCmK9B0WzLk5Qut+InAq8utMK/9neCg2BxI60md
Xt1H6cYzsLs45uW4LqL0QlUGnS7QpxbNbSjXlK6FMAh13ptN9bLHwtKFAyqERGTy
Fvg9W6dxNeGUIAVHXcM0vwtxZ2ILF71VpI6zWk1CE0mc4sqfjcMEj2q6q7CWo06a
Dc9fVSMOQ778Bu+SMU+6GiOxpN577lGXGXqJrrj+Px70wUV3xv657eEn00IEJvDR
YhbCRWi9/KYpEkR1AgTOnCl0HfH8/QGj/7xcRa2VLykI86rUgrBoBR7zE7VjGZOJ
kbqinTOuODbCHk0lNh57r+A7g/k/2uyr5bOb1xqOS8JpTfcctXhH7EZymq2nPB/Z
4Aeq1ClEed8wWc3ARQU5RTAzmPxoyEvBcuMc+8BSqAmDR/RagXPQo0gJeCZ2xWQv
k7qamKdKQhkz7GfdC/cmAHqNYkNkM4oRWFiI0TdIZu0tuaQGN+kG0C66WkdpBawf
26IA5L7IdE6I3ssnQGn6lj4Z/xZA5L9C0IijbiO7PgpdLqfYCKZKvcix87tThfQt
0DXiFgUVX3i0rb8m+o2a4sFc0AYOhVix4kDF/R1JxbCKd2X8kob2wmRdLsQHGH6y
6vnzGDZ6biGLlbzROH+5uX1WCEv793vpAB7Fy4GS2gTftEYFIAtYK/pauEDh6fMS
2VzZIzRW2y6ql1pgOaU+1ixSrzq//10ssMZEJ4eWg8Y1tQfI+cBsdyWzvLr5eiCk
NLyeo+ZDObJSkFfh64Yb3Tr6EkFDL9pwhsaUsDc9uFWCjbA3y95UxwNmpnD4Zehh
MFsftGItfL/XAuVZVlCMbSu9c+PrgPmb99+C7jWHA5ImEJTGgGO6q7+ev/26oTPA
Gm2NSX4lfLZBxdNMAHTPOwB39GudgXJeG2t+nmOjPKR4ziT6/yi/Srxf/WO6MTuS
P4vKWE8Osv+xNBvk2nac+h/vmnQOUfqX3rBtSGwc08SYy8eKy9RGCOjp1I9ubrnY
05HG0aN8pF9plkWG0CtF7GLQYqCCIp6FGZ++CsgQn3xNjYqU6d5GgB+1aXriyLGo
kF43y7GAuAed5TDzwnDJU1iV1d41RFzNQEL5paG7EYY/3+gVATgkk3MMDpkJ5UHa
t+50Wqd7ASU1azGMIOcVnRiJYqn51/tAAIfTLiTzRe79m/09mgz0eIt4zRt4sK5H
1jgaV11M8X/NPc9Lk9oAAT7fSQEFq9lKFluA/Ha7OqpQeYxUwgPZPaCSaTAbE2OJ
uNYUdU3OTiqUMaFo7ifYaICQRl8fWyA7l/PLjZQb02bXlXfd3KhRbgmViztK1dwf
KHQlrBoM65xzZBgGg5WntjJXnuZGthGE3Eq35OTPoP+pV9idQTDvJGlplL9wfiyq
XcKkUrXjnsFPpVM7JwGvHS/qYhWnNUleWCVe2HjadcFNu8hcpOqEoToVfi+rD2kV
sTI6UeSbSunMyK83nJQryT5lQfwnvtGp+xF24dJvu0SMXBRH3ebdMyIxnFmDa8UE
JT3A5gHXyLLVsOv8GwKHju+1yuar+LvNadzqt5Gte8qAVkCKeL4yPdk5pri5/Y8o
zf6XA3bRTXXzoEgDGpZIeAaKWXI6MlnOse4S0M3APbESjo2W8kEKJ1j5OsD9y8ty
QPg0PrVGvnYgoDuea4JQGjOzdea3Gxn75T2ieNaFOpt19NszLgVxwCBdyBISiNEY
y4JFea6zOe6gOnswmCJtltBrJSgx92dJ875WCzCYxTJBYp9AJ4XccHAfzUBtwg6T
ALorfVfCU/6jRfRZyRyXuVlhOYloI9nyJxBoMoA+A/C05tAqIt9SerUJZRf1Sb44
CfRcBh9mH0Js0y69hGHjPeT64ih56S9n0CisnigydWSgQAiaqlooMwCMGijjM7s7
ru+2Y4S45eSj4nj74DAzy+Gsvc2ml3msDkDRNwgIEuepuXIKrV6SujUj1FtKSkvU
shMdrbjhhSAqKcr+cxxiVd/Dm6XLa3jZR10v79+sDQwOXuBroyio5mZUpbkgRHLx
C8C/7quMZXpNkyJ8aGabC8wephHaaTy5q0AOvnhSjCFlwmRhdSUUfi81fjVvC66q
avfLrTnYElx0mbt9goICO6jVTqREtGkplD9OybooIG7/AS6JhSaLe61yjndF4NYs
B9hshinivi7KI58PGwwAhbbvOaqQQedEop3Vby9nFVKrUsmEGXCnTGq7yhFISC+R
hkNIzdLaneHIQKvwA/9DWQcFIKfLiWQuNspc+FhohKKfrkrfn2Lof1czy7gpseFP
cIDX33CDUVc0GWkavaTl9WD11WnRdU2c3c4BHMWUr3kR9R0qy6zqlkJh1wu1CtSv
3eSW4byd88/D1jaoRy4VAJzUaavap/CUm1s1P5uyYOy4gcAEmJNfGWOSnBNfD1Kr
HzFxtB61/VerqtIUeI/jZ/xrsCnF0+jyyLgS5s6aUwzbWAXy30gcb0k6Ag/ur42b
ct3parLtMhy/gJKum+cqHH/PHuibinsBUmBGECnEZ1YB4mbn9LTtCRh57S0al1AM
Mi7NxdOyMkx7zseMHvX1Ll+dIwdOstMG9cuA7xcCG5wPVYBssbB2pIxSToYUkZw/
SC7372KMUjawlLuG9lCTtUfqWoY5gK4eHCoYEEr9EYA16dkbG/gktGJrXyn5YXNp
Uy6gTfvqPoOURBa8Xuyw+EHXMSEOSwAmEwtFpgriOzZqRQmfECp8RXKh91QeIuKv
2d3aLGUIOgF5spbVbjGhU2592Y+rCPR0cHOryWaMRzQybsSxOlZ1OB/8vODbQJq1
CN/judCN30XGwc8VLPLFMhwo1sh3X/dL9e8u/tgq4c0jtJmzsaLlBeZJBh8xbn5k
JstesWsXnHKswqgMsxTEW1afWO0ULHepVIEoBoEQwmvEIXPQN4ZxmT7ayGXRNGqs
Ifn11enP10INbhhftoqEXzNUsD7SpiASWFrDtH3F09+0oJNsnL62XGB0KraXElY0
iPKCt0IyPzMgCUZ/wfTGg2uzqs0ZwChoO/vQ5Hq+F1eEnoIwiQXKlexZWAk8FtQf
VVO3YtPlLB2CZrYM1/ADRsGO3THWc9lt6BBLHhwZSVDu5su34J7w8XWoheKgvn/l
r4ISd8H/Xt77NlrPcsykIheUcXTIXQGhvKvOSDNBjYqcgFKpHJSJ7UB7jGUJieLQ
qKC3n9xUeRZHT/LVCVU77Be6NW6pKAl3UZFnkNQV1yr0BEJO6/l0S68FqFmd/RJt
h/RkJjY6Xog+JaAB2wzox+eNCOkQmWQWIan14u455MPIhWP9far8VJiNXbTkrm7X
CCAy/6VN0nAu+EEjIztplx97rr9/DGbCjE4vNgiEk4PppwjVJ6XmR3Z3aL2BAQsX
td9UffjQclDmdtLmqOXME2X95hvo9eTqT4p6VH5ZV7XzQ9Yp4i3ajhxiZxF0+Wp0
xAsVfRLhuJPHBk+kntK1Mf0ZVjTJcjpW1pe4IDkHCMwQGjeKq/8lO64Cqkjl3LKi
5YQRuqVN3lZtfmaheqKIrK8t5YQju/DcBABOgHc32ZujcXfl2+47TfO/CSYnUBn+
v5lAW6lB2T1RV0nv22IZkxRnE2LaAnov47qwufxKMh0U9U4ZKqjWglOIUOKsHUnf
NOkcMoQov/UBlsPNiZBCqRr6s/H4FCROmjlkC1MXAtMqg575JsQNHDjscEXZrChm
IZgQyD9Hg2uvVC/IfDDLC4ZYsQI4bwwwmW0J97jClSUYLWjcmNQo6TCISNtfwDdO
Umlz4Z9PG1ov3aSkUWesuSHZk8XO8T8TKvstY+7e73QaR6KEyK7CXFTdtjO3PFHo
3QyXJVe+s0SqLQxq1XC6bisfGL6vO5K6DMJqI6iQYkvKbjjLaBmQKECe0LMzKjvO
JkQmXEG5Lf6G66P+h9PhYdC+K7F9ekyXPyY3HOgMzd0EUL/J7RvO8CB2R0mDnTWe
HEgKgcDwsEpYfFSWY+PaWEEegr+G0IdtQadnsGyX3UW+pFP50VfD4sVLN8qefdFd
clzxeDg7uEQbgD596TvJ9TKR28MFD64KxcbUHFG2xqfFdzk/SnyBKcrYUMrCeTEX
TTPSx8xJpGg4cL3ihlpetsik/6qtP9Y8SM+zpozzDh2h2QJ45atVtZ9uRixhtvfD
slNVYOwc4+tmCx3xix0Enqn61W3O5AQWGZ3QEucacV5TTk6tobe2UF5GbCdWLZAS
kQ+yi5pa7vIt2ikKg5ORUGOgywt2DxFk1+UM0/F0JrbI0gsgFUDF3LCafEVS+LW5
zqhK21qGYRyAQhGjp27cF7sXQ4nOowQnrqw3KDSH02aut0+qzEGOHtUhJvV/eJNh
qOyxIkvNB6vVXxhx9HCkAbMhXQTtpqzMP+nUxEGfUqiSYpul8CS+CKheoUwNI4Bx
ZADMdaFmP4Eupv+mkTaPh3Krlyd6dN7G3Cotx0xFZ39IA5fRhZRDHJD383pjr9pc
6hbsQMjz2lfd4jnsdkAthGNNm+zqNwrRuKuFgSRvQnX+Hvy5KdPXUjPMY1lLPPc+
8Gx6OqvTaqwy7/xet0scAZCLF5ExGVFQqNp9fFZpVYCQ3Ojwlvfw/JU3cTxkFjkH
d5YR6TuCL9pD7ClnOGmPi91QduVEEwQHzCCk0gtsrgqfJeLTclM4BvxJIB7c4+Xb
rdui0WUcFgsjK1FgGWyYjz13ZwaIlnqWQxOMle8TZYIOFM71CDb1clNICP1aT9r/
5Br9SGgZRmZxJ2UqVnTTrPLZRmB5sGYHBv38wUkmP1QAu8Wc86iKpXnW4MhJofNk
G1V/rvuSAAzo3/MKNeQib9EIc+tqKorSAf76u1I64ewRPJefLgv8prnSAn1QS5ee
VbK7jaKPt9+oEox7cWJVotMr3vj7CHf+NEAIR7njwPq5aYFFNZqpt3bQqq3T+Vyu
qSiipK1OxcCUSaP7VoBPQwcZ4v+EnB9Q1ANjmutqMwXgWLzJvU4/Nha5VW6ptvag
VH2AcjYqxUKK94YUJL4M+igSuutp3oUzhnkZ/sYTksVA/nQNeZmicO9Wn8VK7/Wt
+VIUH5LCPeX4wRdwkDyZnzeD11wxDyoTXaMfwPhLadwkWOP79di5L9XHr2uUhbpF
N0KA9IOO131vmY0aiuAFILyBAD0p5RqwiNvoZDg3jjOeCl7jZa3bv98NFNwhjhc4
2QzaS1eISlaV7LRDR3Q7zvgdeiUX4UQWrSRBEH+065OXm4KSLnlzSowl/IK47z5M
OaXHKUqETCNslGiDGO6FZBd402L8Be5/bSQXUk4dniS3/lM3TJfp6CUjW/qobXt6
4BQL+eSw2bt76KbfnBTHzxfTR01YlVNynhp3LUXVfCLOL+LSL6Cmu+4L6ClJpFUD
Eedf/dyqYbrcc4nkDOzTl04p7MOYzVSw13K6LEMtaWoAdSQCSHAuoDXma6x5pQCb
kVJD5B69o1uUNwmpREpErwwrag4V4YnMe76fSYt6GX10H3aXBGaaEhJNYNFVmit7
9k9VAUOfO+QTcGGacvvVauw63jTSnbvQq6dRF7w9jl22fFsZhlr/PGjNubbEonlb
im++TjJnERbFqbiGKYkAjJBE0LuQE0yo6KPSA49h5IoO4ZPgA+/iDk1poME25y22
uj1xTPCw2JfgwD3Dd7d3h379SWYBIOLP+ioKX52rOwSgSK8okRwLJznSLO2rn+qQ
caAln3fxQMOJs1ij3z9E83yGv3sLIWtBCJxUcE1oocof1M/H0IxasYvTFV6oOLEU
dYmUuyHA2uklHMwk/Z9JDH+Zlc5hXf2NCBruxk1/XiH9Iy9VGMT+uXngtJiJ+wJE
euOeVtfWVBjGGQOwmY3AV0xre4+9gy+pAbHbzmNokQCxTavPxzLoWimi9sSJrec8
Zk+6HNKOo4zGyYyh9O4uOQNLW6DiI5l2LBtaFE4fwAYz/3LjGF8VNKSlp5UbKB6I
SkEUonGsYarhcRmB/3S6WnFbAwKsFG+wZuGHVCgcdcWB09LSG0EaNRLYzdy4OgUE
3rCV+hhw12YvR9fm/jZrTyv1C7EXBi/XPvAxuN4rTH6Mezjfewdt10GWK7eKO186
celTLyrXT5XWyVQzQF4xsL81D0yFP5i6riblTnSQQ7l5SwQ0TSB9AwrvoCknF87x
Tj+FkpMutrlhci8gnclrNrNFjzVmYFW/np9lrPdgsAw3dvGj7m2Nn47scVTCvQtH
u63+glz33CH+NdJEBnn/5R/s2rR3l+EMV/UaC6eZsFbqt6cf9mbvDZd7kyYEtHlV
fZ2I0gMa+fvyUb8tZ5ocQKWNMyQxyNpEcd8z2VaDOf9p/DlELSgHUsJU8SWMJF6Y
5y4DzUS/wFn3Xw8Gq55jC/bcxIrbHRLE64U4sgGlouYalR+0JWr0XlKSIAxkS38g
2t4GeLxyMykaYyk4krJ/KMDyzdiuRL3mcIfvSNvhAKfXEbazSYx8W4aWJ+l1IMkE
V+ee76uffJw32W5uy3sDe8AglC8AHCceJaVhJvkiOBd9TKtkS6oGANYNuc4fJj0x
VM4sPH4DbxTrZxMBpvKsjpgCuKEdAmqgJQ6n1hg5W12VwlkfQmH/hp0mneifLfkU
F7cD9QtOGqoBUkznqt4JbZpltbr70lELPkUr/DrTOAKwaKFw/V6JCPL2Th3O7ZvV
9RRaQukOBQxBcjIfzEq262PsQXl4Cq5mbLEtvycQ2d/4qOmkZMA8Zj//X7SifUhn
SaVXq5QLYyaP4LLc9xf0+VM1ealankqbmTM6pEIk3Q2bQHjjJ4EDQayiVxe9gX1u
kJmJc873Zhtzd3x7tVT4HlkUTwnqTNB9gHDpSP4gDdWJ7WEBRFOkYZdqqiTa3CEL
kUtGx6fcsE1LBMAbauux+mKxfMoORlHKDYfyJSRCQph8Nr8UEFhNUtB9SzOhFt68
vrOuCWuK9vahoP9lg847Xf4b5Y021r429mlL60EN4pjKllCvhUOLhqUYbsgaFgB7
U2NTxwTAERMWIp5w5PuC058ptKYaQCjDZirHGwXBUYxvUGqu87b6vAiM84lKzWVV
eJmgmY40f1DR8rqW0oR48KxxOHOf/X5sQXqHEygR4vllO7qZwN5QvokQfRwXEHYw
4hHNBLH8gzc3OaUvLNd2t+VmboK5lk9YP0OQEDqKnYyuWuUjdHkV6x7vq9W9xAcI
lvMslPFmC662uC6qP2k/DwsFALW31Wgu+fiEZ+OiurgOI35cVSW3rCjgzZB1PIdc
9oYUQQ4PR7nZcBXEJ3KK35IMq3uuhO0Ig9HU2XYEHgmaTQRZ/irIN5ca05pJd9mL
b+1eSNCgYiE+M50oOhNbpjdUFNbKF+nZsba5+yH3vj2yCu2iA8I/iyvU+Rf7qoDI
Km3H8cBXbOwyI4tN03VEdGsZwBv7ydUojC0phFtLJzV/rDtynYgPLlV/ms1DEgjP
4D62m0g+SUW2njkJ4VsKxVlcZc8UjKmCVp5D0kR7UE4AFBDosJbp6EQ6im2XHe5u
0OmqFZfyDsFC+bWp+DKbl2jvhcvSXoRNtDZ7RxLn3mG/j8YEHEFjW2nrS2nWLpqR
`pragma protect end_protected
