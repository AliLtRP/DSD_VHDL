// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IgIYm9czHS3Tc1Kmfnwv8B88A4KI5V3bBkuvPM3C8VN2MbxhsNxr/vnrQOdNLuQk
EaIZpu2Y2E6tUW6GGZNZergZyrrs4EsoJZDpXefxPfQRLbDrybohGcwyktEC9tQ3
LTWkrHdzxJ1ItMZN+59g6BAg8tlukW6Vbn8hJH8DLfg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48288)
bG/YjhbMSgH4pzN8pJk0IZkNvHqWIPf3r92j542udCteWzCzpg9Mjyx8u84HmMSe
7iNoFz2C8vQUp6i5A7QpT91lsDv6mppHvzzui3ydVAQfINHqGpAQeRvfQCE7frbV
jd1wwK6bFYfR20a5dF/AlblEhRlosya+wDxcssc+wHU95s9mugfVTpwbfC4z+mzA
Wfc/mgRNRsas9CTbXrxseCY8dKlpiGXwVDVgPEP8iZdDDy/CRBd7h1WVmlj+dM9m
e9mTi60Uvuhgi5eYq89Lppo2pfwsubyBl3oDRYaTpLn09msKcC3tr1ZG9rKSx5QD
fkH8SonMhY5h6w81p/u+O8F5+PxqUnl9swdfbIcWWGSQQKeOf6zb3BRZ+tfSzofA
dxtKNXuhIYmiqlvkTkldpW7XDdNy+VfOLxoMU2KNT2x6zmTSsjPpa1bSN+c3GhYO
y9TXH0tROkdHBy320scjTz51Yaim42Euy3wPVY8913KPiAdVedIJuyjuNbSNCf1g
abLDj5uFP7eZOz+fuGwRQoz3s68k+IiqlHdl5eSeifUbOX4XMtVFo2yns5ll0/J4
Cl//AuGACApPkc3AQSIkTONr8iOfJto7vI3sLDR4VItlQzPErerIPXDYxKC87XgI
NUAub+a2lojGrVfPmKpAAkr+EQH5APfX4LMYDYIh3XXB7ga31Qz7Fg8ntDY+Voo0
9Exq2OB2hopL1svkCRfL4t3WnV7THyeYwryWNr9F2MJw1fVhk6qBetwqDkYtD2gv
ZmWvaa5K6Kf31e/haXly+L5WVL7G21MoR5p2aayD+Vdj6G9SxZCqlh/LmN4r9ECB
JGUUYDDRkX5V10h56+vNs9vf5Xrq0Mkz0SPItdTnLH6AWVCfobyajks9vUIIDX9X
8C0jF96paGnU/2BlSOFqLJ9ufUNtNwSXaB178xnVup/a1vIXkcM/k4TXlYcw3a/K
QZ8G3yxvJP1wVMdhtdAHQw0vmOd04yt0xpCviQTv19B42neeUgEcivMXBCsDr706
Ccob9BrAKyaSSZxfAHWJXyV9S4PUFApO8T/pdgH1bZPIm5cB9wQqLc37g0lTEUgn
kZA3EH8H0laMhvjQc7u1/+4j16LKAdwkYjsedKZz01giV/aP9VxE08iIKlQcpy2O
vzIXrfSciedHoy9f5OP9lflTkhm1G1+Sf9bhOIw4Xwc95wkx44m/0XHR4uZJ5SdJ
ejWQkYtXC4i8M/1n+vASekVTTM8NWEtXLvx/7jpbhPHMDFK1rIGnSWmtktmnrqq/
gSxMhRVLB57nufmUxoNf44uAQT0ujn66JmeWeJ/J2JF+jt0+Ktyd6eXmt5nlzoJG
FT8fLNhe+IGoGYBbH6H7p9mHtqDkXwM+FxC1WfbZX4uLvhjgOV6YMHFN5xVUExRn
PecDYei1n5NjtZ3LciSfAwJYcq9Qy1Pvfc0kBWPYDqneT8VkhmrCFP2RZQcvsYkD
q15Nqs8kgn484hRkbh2DqJnp55Lt5BKFckggHVsV4TLgFHj7o0yeqyS0jBtmL7lb
9Fm1FPtJ6kxi1a3D8rSvDhu6azk2SFPsQc7gvDQ1bpVuTA2OUcA9mcdaf1yIoJxn
1HKoUEMpPsCnLn8/dPpKtJtPehpY7X7qIwnx/HudZLv9I0UTrpj4dMC0VWWMKy9F
i/XKJMtGZjSa6fFLWXpS1TuTEdmDs8l9TP4kyExVjj4ZQ023atdEBOZZwWbUkx8P
+0Chrn17GIUKi8OLidy8Cdau5vSQcj1lL38fwZBg9WGMRF0D9DUFx90dEeBQU9zF
fpmmYgxq2uoa+I7xdNWov/EF0MNZO8/NBIo6B3ZfsewyCVEdMIXaitpdrwYBte3+
S2mIN1YKj2GDVDYAPGC9cOe8aeL8LiLz/QzDQKKJs5hElqQUor6UKUbn+b/3ZYDI
9auGWr5g6tFqIm617xJDIXcAlkpYov9IvEiVWehVvIyeLYmv4uDLZN7/rYN4dYG6
TFAzeiPhD0qNdTQrE86qGHhSQ+awyMpFzcyIadr7KNaDVx/LbfdZm/59gvBUDqbq
Jg8we8B1yA+NfJzT7jgFFobNd+9bxVB+lWzHUuxeAmtouaC3lvB0mzGSw297dN06
OEzJvJkor95PRw0/PNpfpLgw/eKV0WtviM2A/B/uKvfSQLmyn5lUejKbICsrW8/f
euGy6zRBB3vTqm8+rZLVh6IkSzGEN/bZ3wQCvJ8fMugPoduItmG3GemilrD1KXqu
RqlajZK8IcLmV2TZKfIJCwMoGchZBKhxtIUlMGdBdbBGf5yR/qs1RnUI4WAKAGOz
oeeT5y3qMHwyPcOkvwGloPnEHyAp06dNdOkmLkjmx6MJoZILtklhgeqzyOoAKRSb
1fTr8tZZt220dm93Q910r2Bh+8rv5pAlvwfiawa5VFvv3QVDqKWQwrDP07EtPaeY
rP7yiuKRmnOv9M4nRqoQISswYRawgV23LS5O3XJ7lRjE7hKQ/vEa4tq65SX5NhXm
iZPx936ewaPq1qVGwsPrpc2tfXqkwXqJU+vdrK+rY+wtwYgxyLC6DcVHcdkZXi63
SJYp2FupoNVNLlh4qaK//EeYoVkDV2Csi9ZlAiLDnvSSSe0++PH4hDVSa6kJmIeU
ai+ebfNS+aUt77LmZqAlz6OiEC5A/4oqvroWg4bfNGCTBhgFWlkiD1RGd3QxMg7H
9d/MpEcag2UaL7s3u1Sw3uExZX+eIvei/rb44udVrMT2of002Ye9qSCDte93EpcR
xARJ7ouV9I0s1mtnT3fWKYCXivC0bD7XFpFuoy86W/jDbp1HzoEkVYE57qI4Up04
y77k8G5D8wIgm8c8beFEeuCEl5yM0ceka4b5jNELjoTKH0nx4WMmzdd0zCpEDJAh
CmCYpvfKF/Oz/J30s7UbavdsYG5bB4XPFZohWz1hnYQ3q/6G3IXSVy7Bb8HzhC5q
GPxEZN9Vou5pSPfZbIqKLwssLGwnnc7BhcC1GAP2mDC9tJBub4ThEY8PK/Db/aiR
poAM6kRCDN90nf6kDb3Fri7BfjK0BIozbBoLv24Mzrru0i8vTpXZrESRSPHhOsUD
GsVqc4mk8MCV/B7UiPwHwt5XMMoPWTGPWyouqAqk2WQb7v6p00ZaodbbuKX0bHp5
mhebf+0DTF/lnzYSbCB+ZNhNeVR1a3v4TEdaePG+oMNd3tAtY8OLGNAKWx6cuATh
MGKuwkBsHygQEgt3LrovT16u4qubrJuEZ67MvddiF8FpF8f5evH3k8MHt4pMSlou
SL2/gwFWMpWLHf2V2TG7KhtaOlWeFpl7Umzi71Bdf28zAw6RK2+JOyE9Ay2WBSa3
MRFtpN7wvWgEOhLj2d15p31Jy15Y9A4XlAnvE9WJqP/EixcqUBY3na1rL48GEL3b
UJ3GYdFt1RdPWkVYvipJYNV5zfPtr8wYSdH19v7etSsZDR7wBBtNy5uf4az3rIoo
cKJnJn5JFWYx4vs85YvoMuwvifRhoxJH49uemgILY01b06/FKL+sd30esOUN7uza
BJJD6u4Nfv/wiG0h3/uMbq4hZ4pa9H+eRciYuHvBElavCPmPl69nQ135a99m5QU7
xKlEZbc7lLWVhbbzIDCFWt7zVy0Cyj1GNHtv6lcan0J3AgIlrK2YH5tHxQbHxu/A
ySdw71UoeRmMtgfpnvSGKLrp8KN4sJXcLu/bPV1HF70KA9CbzHCOM5T9+gla8eFA
bfl9ChLmSjZ9iuMEpaARVoJOxCyS226p+9js+jAxx7E70sCJ93G8DCdke3nUnA3m
BFAbH34tqsqa8+1iI9CDoeVag041GX7O/0bXCJ8z6lH7Zl1ub0d+U5OHjTcR8ox+
FzPBJrXGxJ/EZHM3cxlCced9eTB+XdtwGOGLku0djR/9UPckpz03BoSTSubB4qrF
i8fINRngkXUh47RTkVPDmSzRdGbfIkhtbiYvg/UegU7Nn0CB+4NvN3mmUNAG4iqI
wmP5QCo0hy+EPFEGbHbIC1du5FRE8DvJNVbKXO162wI1+H+gXsXOPgjJZPbkjPDY
CKG5r3yhd47PqVkM4imh2PdHSoWH3F+bx8eEtfRwgdFX/KhTF1kucglaNQe0Qczx
AsQpib0l/4GuL0jteb5gw7lVcjYvruqq9fogwM6e2JMXiqPfE7opCTwATfd9oeBE
Foj3pip12oF9MoWvAOE9HhBZaxdYZ8bv6MMDt7S1QMgaP8NNbD8oGg2wf9tvgd83
6ZtwDxIaTEh0wfC7x0nFOhL1tYjkGI9HddFuaLIovTDSjb6oHIe6sMPwk7ScilKS
OYQOymm3oAoPGFiUJeeR59GV1Nzz05pYeJhEp4KhdF+0jrOps6CdfguGA0SsJY4n
BByg0Nl0WrVXYsfvdYHnBLoN/FhhsVnypsib6lQTbbQel/bI6h1L1o3zjibhg2Dr
0ZDwth2fbI2ioOpR9C3fUHgtpxz+IGSy4+VurX6qz8BH+9mqk+njTaNEKWls4C24
vdp+s/nUO8kdpfWPe1xOxoG91c63CXL3ztqnCGJDaPzi2XFkgQJearOW2hsbu0rO
+rFoqdDEgUTt+6S8Rr03eC3zx0NHl8SG+kXWf+GmbLwPeaS3EDRIGRtLADJeD0q5
9bU0I5GmgcrSMF5zUIXaWywzf7drqhZA3oljRFc9yu7R7A9kWPrGcOXlqd8zZX+M
m470shN2c+BTAdn7HYeTsnr+69+SogmrMA/bBgW8S8vgqg+oo/Cw6AeHOLmbMU9m
7lg+r/Y0lnW4b7wbVWpzj5yLI64M1OJKxxttMnX3Oa3azgjjfvm327bibWnfXbEW
/s+9vzGI6cQo9YiJUpIo12oio4IiE8DG4MAG3t0J9fzemczqYuRedhjJzvZYbxUS
OEhuT72OHHYMg0EK+s4iAF3xxfv0HdQMlxJ7KeoyfIJFdn1KZWtc6lOUi4T7xmev
BOWEO8jDGI01bAVQJzmEMlc26e/fwqclRXR98i8sd/Jb6gtP8SDK35z13+27FjO0
mtKpKNA9NPu+nEZj+ItXNh9PnKV+uCdk+rRprlG1cWQTGCXKi/B+AEWKSDkKeNLz
8Jp1Mm6qcURKvAlOymap5yaBnjxRWLbEuNc5GoEcXv2NgdZA85oEcqvhJ2e1pRsj
DqR6I6LStFluwV3VXKJoq22QHGb0F8cUR7Fj1lrOmMpAStYfrXxRQZ2dK+n7ps5A
mkavb0rOS651QGqewmw71KrcLLSRkX3FTSyvAJp5cJCeA9WyBXZRMlnpgjybB8nQ
kq1Qn7FvlcCJ7cWrvzEJ/oyppW2/o82i6lAUq6FeVcbLAFL3KesGvzMVj/9OjulQ
qBbxUwpsl4F+v9WmhVMqyVsm65irtDPmnzPqHb9mV0xCCpxYUjDbOqpt230UDbyk
t8u3qRXZUT+zha3v6cPgvBMreJV7j3pTmaXSJmn6wf+W7uk0jwJ1X4OL1jay1ohw
dkcw/z9NlaV3Tjh9EGmSgTK4GGnmqLy1N8l5vNi1YG/ox/ag7JXQVAkg4TH+6KCd
qC4wjD6E4hO80U7SHyqex4ow8bUEBEAL3BbRPQD7djvfiKPHgvSD/PVmQgy+pdCl
yw6NTLtjSorOo3K8h00TuSLZJQnvA8S4hJqanCcsQuMxYlIuWzorCAosgUSe8hu8
6IS9pgnCcSTj+d0WQX63CTbskVT2AZEtUt6LooCetpi0xvdKH3FjyCZJMjjnGYgt
NRf+JaKpj9A/20h7lm8pjG+Uz26w3WTYweit+hqQvaqHxFUM8OIrWgHEHp6gkS9r
P0xHdmRiOchlFoyVATPtTPGYNr9i9G1vz584Kf9c2Zplt6pEJYxmmZnPjHUZeaaa
6GOehB2DBCaOsj3mo44O59bMYr83Ox82HwInXQ+jeoaIBa2TeqHHyPcTZad8E8qN
YJINrDXv3SaXGP/Hnsm8U3EEhgXnTG4lS4MYBVkLly0ahPpBkzRwYDyA2RfwDBcj
i9Nh/kSN0qc+xICNGpNPtxyTak3NRn4e/kRPSOAhpk6ERBm22WOHZpZFCgt7qBw0
EvrUp7rY6mazJ7bBjl3KNL9ueMptmiJmDy2dn+wNAcmkxm3gW93IPS7N1oHZ4dDF
379hDGYclNbH63NSHCiFUu649OmuOYwtsFDPUuZXIZFQFARQ9AKrLdsx1ILhMFCA
O3+nw1WoFpOI6pICx4PduZkRUXSrMOdZ4GjJF2v3Wt3uUBluVAv7EnC3kK7ZriOg
Nw/t43JttgtStUM+JowX9e6XfQ+dtWnMTaEVzcgOmbEKczNEzpJ6JGWEjC6mZ/he
+ydZZs3ghqASl7huV+YKwUoLCQlb2Kq8PPHp+ZeAQMakC6vgAriyuyltUzIxlusB
sPyfvfe/KJ72tTkS8jPyxGuHvp3rxR+xs/2OblZegU9uL40yu8wOxyMpwKqy/ocx
9PEC5i19ZRNpGWgt+MZQMHX/tfUv0p4KzoPnDWvwSKJ5K1x4G6/UJ6Uamc4dPlYD
0WIWGHd0zNnz7rxZWR90h+wY/KZYS8jbV0JRWrYKPh3s8s9vODIPp2ohQgAldlOu
NfzPqcUEIVrpo/Qca/qwYoQ0MNM1rxZef3/EklkRJeF+SLyQNqvxDIGpXTzF8Tjb
/UhFhJdg+Pnt9+yzdUp/kJbO5xlB4Vo0nyuAXRQb2T1IMI0TdbKKj5fBvd1b9YeC
9ApUGRxAVNfgm0/WG6MZaJVY+ZyNwsyFtM//sXjc/hFwrvhsCMDO2+zPtAVBI9QF
Vbbb/7M95fN/3CM89mSZVjVN24AJBGSH1APGrqkrVS6T91OjNuJQ3ZEpTX4/cOD7
wHrMH9l0hwn8+DANdodW8hrmtoczxpRdCGGoGJLW3QRbS8sb1pDzWO/DTVcD+t7C
etRIxKm7FC9B0AmD4gQ7+SKg9cQLxGWcTXogXqUhjQCEDoqrbbrDjMFYWmW2H1tv
r5PCRQhmzUSHzxg4z5WSZ5kXFT0/rCBhDf0XaX0G09pPZ7yGv44SBrZA40HOI0X9
yrEsU0ZtY3d54JNjbkJYm5jUBAETFlZAWCCrisEND0yizzfSv5CtaTG68LNC0VU4
a2ydY7dfWPriBfRWMc30VQILsf4ADFNih+pJPWlez668hxjmQaZVGuy9GDVxYqoi
PskOWWLeNE+KUxCkJvGRtFGxaZXDc5oOshl2QMxx1wl0XgM6yJaWjp5dQY1D+2dt
OqKB+fQEZmqrl+YeaCTkJXuvqwaajyak2NDzOexL3kdHD6ISgh+LSHnX0pFroK04
lKgTF8F0Js/KSRdVWF+B1EyFqtZcqXYxmn3YNl2kyZG1DrXwykPzMVZZduxtCpy5
MAOKA7liTORuL165B7vJTZ7LRW9hnabPBd4kWza+/VoeNDHOmOtoz0AOgwqyDwiv
uEkNZEQnR0wpvavjGHTNPTG5Huldcw4aFi4T8OvMtVLTCWg8D35WpT9+MXrE072e
vR/l4zdJxNTApwJvR4OCN6sA7mdYaDT2ypKCWWf+4TiiA6P1r1hbUfnc1UWTPzV2
LpovxxsaCOGLKS+f6L9MK+/ikAIOnkeNQ8GCNsYRhxpobJiLOF3IgwgbrUhT7pjp
rTMBjXQ7x9IF/TRKTvcVmdFR530UDBGpT11wqcRVIQZ4Bg2sL72cImOj8pk0L7YZ
wFbdl8ojkJV/I2XWLu9DYurAJaXSaM6euZ6/6rG4/4a+IN4zbQXlElJK/SJfQmYa
ueuXg3Eto8JaS11qiOMw6G6KTYdAPe0OUBxeJB+zYc+/AXS7lloVhg/mfJgBzOP3
q9z+7Vdlj5J52V5qtCHP/A5Pjc6LD6bwxhwGnK4uM1d9r09KjsWzVdJp8M6cQfJn
TT1l57gcuGDtfMv1b7y9jX2BgwJ15/aMkG3GGnnV2cB9cRfYqHao8IcVFACDT/FE
oNDuWu4gpraRY0FuftS5KFRP1RMivr8L7Gv2G15nuaQ0r1RbeaewwvnpdM1p9pzT
RZFvUx+enU2frwgD/GeNRY5LXqXCwMMCudjlYCpvM5Wk056hL4U/ecHMmySs3mUJ
1xv7fN8qbBUtQsOyG7W+BuZ2uiJHR5Y/qycCcoVuG0sBzQvX15LVul+Ndc/Opuun
zOl0pUgX+dN/9rIs2vIxmgWZsLX/JPPif4s87dFXfE59xZ7lW/HP42YbkNNy9bET
ete9VLifDe+iCLZNAbx8o67Tnxgjivj7MZ/EKX9KJmkBaXN+RghwLuVpryM4Cwmn
EIJKqvqU3RgmOuGNnm3wimZB2UMRfpQE7Sgo7LWvFgkwD/UY7onbKWYAw85bK4Pz
srO9814plsCQPpzF2psz5cO7nzKXnyJkLu9qzPkDrHgyXrCKwqERP1C72qVVjOG5
oBCfTTAfKHXO4FwisaP1HfgKzZws+cXvedsOiLgdrjRUubmpiMv2VucVcJfnr1gt
f2eIAPEbMgIofcjz1BHJVXP9zIB799X+yGLISZ3Zl6c1qlEYJXWvmtMz2xpT1uvQ
p6MOoPEqEnBc40vdwxrGSaiqp3GXiq1uN4enYoqFavZhvFPoD6FKk0RZx4+fp02Q
/faqtfTKsAA2aL5XkX+v9WPsZ/LjQ1A/zOPXXUtMxxNjUNr6eAUUXSiTimXjtKkP
2SGLF1uvlCrrRiFKQXrg67xI0q4lSaHrVW2Jxf5ANXOjTvw3h6yq+EGQRcpbpOxG
FXNHl+IabKe1VM8OZ+Sf5sVb8euVNxlovx8LBdi4QcjJf5AI4hLF/NV/4p8Vn/+v
gbe3AY/r7wvlw7PTqwmuTgWkZj1p2ECqzAZtatfIRI2Sv7JU5K7pt2ovj4Ttd2fh
eEqU5BooriOejbFwGWaQ90LXhYaQ0Yxta3onpYXP7R8Z4a+WK72YBL/kPToDlNpC
hHYhCbMEX4i9Vlm9dyJurzS+kVvy06cyaCs5YGYcITfDCemT5lqnrbRkHd3236JA
sHdpjRiGnHTTYNMOLezEPBe27PK56pN25uZVj2Tcmy+NL4Rt/ibL4po+c+50Lmnb
muiDVtIRK04T5Z6Vb+oYToAGLaF0gkW1k5KECQ86LHnmpXaTY9jIInatDFlkl/G4
dpvO7MlhFCTY18sWJ3GLW1qO3p2o1BDWqS7/vgO8Gsswi6Sa67j2MoUXp00GAUG8
jkB4+RuhKLo8lzpIxbwqeYoLcYBwUDsjXe782hPB3H94WHZXFwlU+VqF8wjPXnlD
bhmbNSyRYzW6m43znk1s8OrTL85hEziFFib9kZks1lhjchR0hxgci/Wn8kedLQpP
bA4CRd/90ZpziX5qzfaDwD0s8K7ZouLEQsc96e5wQBzurFxx7wTzl63dT9u2RAWX
uLKs5awyIS5iy6Am/Gd2h+zAOiOeyrq3vRimRO5A7Rkj5LVkLEP3A/lubouApvgc
ugQsO1FGvCUexwzonaf9nMx+GNNWjnNtYPSZxgA7xQKSkeT51mPS3JSYBTYNqj4S
4S9De9KDjYhvI5M6mbN9hciubmFvTgWQpSIQS8jvFC8w7Q8Sg+zWIa9Fu55mkyNI
iTeSEjUOWoc66glxLA+OFa3/b5ccu8eZNRhVb26tm31u5H2S6GQPyPfgttr59TGH
juRPTC8Jh4IgMMjg292kqnTg+esQdspFiDks4/jHW0IRtq4zMGSGQycZ9QD3Mx6b
Hz3TzuptO/IqyTGKEPg2TtHgFunB78oaHe51UylBotb/yEeY9mD2HWkrtFIHFaCm
WTE7n5gTNPHQgkpMKpkFglLwzLlzESaSWHeihq/hi2SPtsSoYNIcQzV+HLktUT2J
5OxfXHodVedHlwO+yGhLzXF2b/6tzyLxJs4/6bX0RwgbRot2BsU+130rhu/KCHNj
NNjKVrZTMQvLhhQ6gnq0nL3WBEZ0k8sFR+wwVO76x5grI2grzLCiEJEI0fRmRMZk
rqjOt0BiDwhbcBA2wQ2cWSymECnlpd9b5u2fQ+IpE76uSAKuBHcXmKT+6iXbZx9G
SwGHSwFRKooNOA0PilTx0F2hQuZF92cN8bvFreUyzRu19qff5qZBYieQ3vJ6gi1f
W71U9mWt1nPTMseBR1tare1e9krrawR1Z1Od2PLFEh1sC2RfdCvLn3ZdGuo7JqUb
1+s155WmVjEsqKK0A2cwsrsVHKQhf0am8hziYWX9Ps8pj9IMtaQ71T7ITKNd4/iI
/uWCFszI4PHUe2bjbx2VWrd68dGzyjwBk6qUqFmWbvAHhMQC4n/OgZzKPV60AFXR
ViB2YjRmNKiiuoLoQ/DNR0NJQqI9c1h/zhDkFDgKJlKSSezrHd+TbmqwpQKgBmsW
VwCFcwJiHvk4wgTjSn1B31+zhDJDmuvhOEVUTjmhgSou+PKy4WYjElTQ3h87kxuH
dohannF7idvobFrLnhQOYZOgK/8Xf4oq6UwSAbFcX8p8XrtPCAxunPdaqpCOQsPJ
HlYaT+dc0UInWx//vVBE9VaUgDVjiiKti7W0kXxJk2I4XNzOB4sqENUeG/czr175
MhRutLcP8x5qt4WGGtgt87vIaQw2FDzfYo2QLZW70zTJcAbUz+mq3sJJECVJL6K1
XwFV08XFUAzrFALvFfHirk/wmH1wjK9vwFgIknzzI9FQRtfFH5esB4rLDGb2o8ST
+dgO34Kk1tUX/GrAjrGXr/dWWIHeB83D7Exz5bKVDJwSRA9yTJvaIj9z38m3flyf
D2m1QTZ0Bk3wXRynpL7ZwmYauHuCao+X9xrDQU+scSayUxV9g7DsI9kZxZeniG5+
9mzyBDSksc3Zl9j/dSwpPY6cOWCyNzxNJ2yyzVfq0I6/qSiJkWCQTydDtHUkVKtx
mvPsZdiN864KeauXRoUHTfEF7TtK2bIUtvFYnj5OQOaVsYGJqhu1IpcCGYOqx+HE
G5BwPCIqFM5dHMv0UrReVsrobjFXofGAui0QQ2Z6T/CoaxELB4JLO1COcZqYOMYJ
pyvDAs8asdRVjMU9J61yoxMUzM5JPtPezg0ay7WNCmV2javg5xFbM83uygdPCBeI
hRltQaFiEGqynt8Yvg35I+xJjN/5+Vij2SxJEiTLH8Bwi55XUyP5+VHrH5ypKyRk
ggV2gBAorgbSBkIpsVbVVJqkdLz6xbJx/P0UFQY6jQgaj5gWq1ikYjTARNmEM3gb
ZAuJ2ILLep7nvuqG4NifUlslwgseeva5l4xyzhEP7Zufh801SLq7rD7EFqprxOgk
TxZo+QgXCbYejuFP/HvEEj/EzGyhXEKnR7EFVkMjc4Prox6F9lwvE6fR8793LrG2
vwzRXenfOVYXlPaEw2e/oESM+UoRlQA8jNxvRqljhd0AVx2e7iHmAx5/QjbMCWMx
6FfE7og4XUeJtpe+dDri5DZo2dyjjse7hK2faQ3uzzjXg3MRz3ZkBjPDFLyJV88F
tmkNQ6xiDoR3kRJhH7NxgWPXRf4Q1SBb1Ri8nrMwfDsXyAZKMer6VmQwOMLUHpeR
KYs1oOSSBtvNENk57QkRCTCL86qpwaZG1JN847m/JY3D1KdJF48Yo92jd54BuV2+
ruSU4Vu040FZwIp7xCPzS4z/M6pYRlttDPw+RV8of2lo2Wnq4SbnmSrsGSl6w2ir
5aRqfxYglgTC0dxm04zDkW5UKH2P8gCY9x8TUeoYGeYIDGLlgXVyN+mEIVchFRaE
r/CZAFk0UY7dKxuQ3LqLqo1erkiZbYn3NnAgOaEP4qhtUUcmUJ8r6YvSPqhSu+54
mwf6ZU9G47TXskTJkcZ1NE3bh3uzJIGrAhAfwTB8e8wwaXR3UmO64rj7x2pXaB9m
KAkjdaAZWYPbERTbhlNhjFvHST55MVaa4cQgoIYJquwip66JdcoAcXkJPJLWS8Dw
cboJBjS1T5K6enXflBLQnX9LIAm7v1rCGO9bTOk1PCL9bBML+2aIClNAB39pE2Os
Xq+7s3i5j5yhylNhbCuJ51XSSPBxR1xTUYTZSFcnkqoLHri4Zj81kqyvmykxPO8T
iZvr53abrlr7e328jzjUocYz0kiAzSCyAfebVZmSrrAFHzx9OpiAfGia1KgwajNO
Nd221dC60TL7BwtN91ASOJhsZEToFXI/u/6rNFRS8bv3HFZChDiKL0u+29WAGBhb
Xu9xfnJlNx6CdERIPc7kb6zBi23m0hsXfZZyvU+pD4acqnHvfG92RfAqmf85j4Pl
slGOlOQw2d+2awM30VOmi2HUWkmHCQFXgZ0c6OOsoTbw0aIto+ALV24OZLNWl7m2
CFC/SajyqgCDM0E4k85iIqATGa8GKxnWHZgUCdQlfaVwdtc9xBcO/2917NQY6l29
Ymg39FtrFbpOwY/dBzwkmybk/lwS8a5gazedrpUPZx9sucuR3vwN0+bdKek4u7mx
PhiUzUyf9H19D99GMV9kJn1y/dGRchRKyY9txtzbtB7Q1drFtZ/oWTee2+LZ5o4o
L/e4euPfnS8xrrCf5B3V8CJ6vK1kpKsPH1UK652UFrHhLnFj68qyp9Yh+kcoUTcJ
9RAQATwWY5gFW/gSGrej6VMhlK7Q9mHKRlK3Mctt7GG8ZWIal/DZDEAHgHJo5ycO
tQz4U9+iJgp7P82vAGM2LntL2yJdIV7aqCK8XIyBOJ4eqI6yBtw/O2BvMGXqQt9D
ps0N0eajzgrUvckv82XO19p1ut9hMYVmylix+IfbddTLUN828uQfckVd5D1Lp2hV
EPatRPVKho4Sqc+5DAHWJ5/2QfL/Qa/4ZBB5E6e8vQertHpxbxnrgAdpck87NSEk
QIJOotExi+GPPv6VQii20JIiqrovif0YeXP3YCJlMC4l5c1M1viO3CVggV5e59h0
JRFQF04ShW+aAsLQBnBUA1aYHp/N+pZR2N3RjXPtSMIW2awsIlDFttB1EcV+xWaP
DYDidVi2543cWcRtSDyNWEQPqozZdNxRoaAVyU87I/G8AyLnBghVYBvWEuwW6PbJ
WQmWeoIltncFKUsJuQQ7pozMyP+hBaJS1g7PmOo4+kiCvYUUZM6jdtnfDt0XvTwF
XPUFIwn9DzEsHo0h2T9YwCm5HGl6KCJjtRz2MBNb4h27k7nasqEH4Tu2SEJ0mDMz
wMOlStXJ7SUOIBB6528PmumJXzzVOa6+DOWUbUvWdh5OnHqHJ53js6KKT8l9MBhs
/joVEaaXtRUyTcWrGuAciNMpA3W/gcPDc1VVIogzJU/B1dufKdnUOHYBbYOVzfCY
oStv/550J00ujdi6uYaITzuB58KXnvOS+NO46GaboMqL/KuuC0RF2JFHsp9RMEVl
qz3Xp6iwMCnnHUm5swypCPAVFMu7Su69kwW5lKRv6SIZ1lFxJGNzCSLyRzfLzgqD
ZMYYryB93L2loihn4MmM931tE9VZYN2IQGwV64/xlC5zA/P4Dil/QUD9X8zlO5HF
x4qYjiyofs8EKJ+mppZRfyiGXyimby7UNxuYecP4LPL69XoiM2BcPM3JU60vxUce
W6tf+/l8lqp/bDlfHKr5QbN1PytsE9NE7bMkpRPXxVUTo94HOoUkH3uRS5XGdYPX
QMrylAWOwFGlPXSdbqjl4BRe1uHWbVArhIo7hvhI400fc9uZfDLjuWYCrE11bslF
Md5mfkc+ib8urdp+yZ7O2GNoRe4OdPGobmVpmsjJ/uMPbwJOiMIRIEDj9odaBAHg
u25NzgmkXj4WgZKVkqHpUXPCljf1py7KXVSHgZOss7Nn++NEnYdzRYa614+81gHp
EjHK32Zz2a1eCrWxKRXxSA5MhHK8q2+qf3R35rIkfckDYRieB6FQ2PD+fpHb+Tuh
Vla10yBY10uyB9bb05d8JEuYmzqytzQjBaQwZE72y6w9ehH2eFwMICINaZ0NzCS+
GyoS/d4DfiONXUKUG2xcGkGNU/g9NQMYDvWC1PaKeUf9MOphM3t63lxIc6q/oACn
FCujWsJadqEr1MMivQAYnW2RlI1t1c869nowX4IXonFB9PL0v63aWUmnvrHEsRgK
DbKa+jS8V8tc69RZG0PQYue+q+Xnc72vh3oJD1xbeOnXuYOJ8jCdhb/ree2MT8SU
oUDVZS6YbexvMzAHBkss98B43WE5kkY8BVUXC9ZUk8Fv7ud2iKpZz0YGAaWe3+91
EKIYbtByWGmcMKsR+0RVVSfonfPWeZlA8JfyGjpxlmj10XEGeg4T/Gm3jm1uDARL
Q1KpLffc6u/v2UZLg1qSeufPTuWWKulG+CS55usYaQGGGUJimDiN5z6yvYERQaCg
8A3Q3Yvs+XzpEpm2tW7juFTf9K5CG7Jjz8/Cw8iMGG2e3KcisbouMLFECcdCEw6U
S5iGV+vZdPJC/f66ybMDcNNfLt69iUMnoeqheFO/t5cZ8qjI/4ir/oWDMoW2hpgS
OD/rCQtuiM6cnDoiVAf7vUvFhzzTK8FCurHdDSwg6lB1kydUn/VmXiQSlAikviJf
9I2DXogpSkIh2MnOvI+MKDo73PZIN02gE8PVW3mBQxa775l9RIBTERR8vQvEAwYv
d6zC6utK5E3RLoeaIOGpgIMpbEj1goJ71QohtNnXc7rJvSVQ3HG/cLS7dpnvwDlJ
CNqv+hzn8MEhD1hE99tQd/HGmMPuxpZvtsdfZ7OXUsn1sYtncTCwPf1AuIihuSi8
xck3IHkOpgTFbEouttjX/NvndMjDWIqebyCrCFXcRXwZMD/gRdrPGzte9jJGB8OD
VQ1a06Hs1d3mpiiaRac5pESEPIncjP4Cyq/Mnn80AldFf4ioCT2CnYyYiOkYyz91
D7gau+9PUmHMQIZwwe9y7Ib9i1hiVIwDrJaluAlicZYNAyARbTkEWSjzgsSVvXEO
tLeohXD5WwErOXlkXm6Eq9N2xWjfQj3PHB7zAaJQrpZWKKA+lgrGyRkQTmzMIJAK
cKy0kRGE5/i3LXJw7KX1iCiJvxVFnY2XtJ+YhkgBrhUixvjv/FBdLeQnbqMUJ4kk
GX6Wl+GE9ivhO6A5ZpWshl+hPrShr1gNDXS1v8zDh4wsx48krBJmB0oh913dpeV8
sGNkO1NY1WdtWV11ETWtHdBjNgw4TerDDTR+l5awz7EQMd8jWigSrLyAFvXi/7G5
zE3xCSlac/pGrXqfogRQLAD1duWZIoMq8enlMBcz5eeOVA83r3Nao/blGkWM0lhi
zFWXyZElvcNqhwD84bx7WJ8m+jERl9BvBYyZp/cqJ9008eYNdeuLpp3oK+1qL1xQ
DHmZowRzwC/MjVc9PlGxN5qdwzYDSzlAMqlK/uOz2FdzJ0xsRBYyF12pDKKBbU3P
1K357PzG0H5KCluZ45i/v4K3/usra91R632Qcwju/CPZYHVaYelil6/cI8k1VD3D
//t5HegiXlObWuXGEXJWyntS+SLB65ZtuR6Y+BuVNRAxuJA8spPcv0lQpimhfsuL
JiZHnGdsZIUO8KDBxSMxTLDiMFGhly8dJUpuqhvdUZpRIJKCn2InmFj/uAGDVmrv
Ai/0B/Y6rgXXSH5360N5bSOBThWR1YeORGHdiwah/5xtS6JX6z+1s5zU5liTqI1w
uuJxsr9fXJ9jEPdxn0aN1gRRDeUO9oXqPk1SzJW1OnLscLxfVyZ7aBQHJ+yLx3hv
Hb7WtAiiVYo0nqzpIS8XMgvk/AxLaUY1y47nXG9MyDVs06MzE+73hyb9iHzGLF1E
VvslXBPtMPkj6EWsL5GQ3tL/hU1ppUu4iVbn9KS+KuYTuX3jz9Hger5Dd2ds0vUJ
GEfFJn/og4+83vKngBmVqCKcfNZb0/EsnFY06MtqK/Ip7kdrKVfwRC1lJndoXiX+
1dYqte+IvJQ/fr9nbZfdV1/rcfR8SrC0KYc3t4ZhuTZIAvY6fyjk7SgBBYIgecZw
lbhN3TnyVHiKfDotQa1/3m+LUA5kUcHoxLoDck4OzfVNiWXqEHmF5BIpjcI7ADfZ
9eic4wax/oB8gakj1aCQsvypyvRA8S822CVM77YtuYCYk3Jyj6C/RPCnUigX/v9k
BAqn3xpdXpV1d4F97mjlcbgpml9tGeU90h35S2fR/mX1XRv+qNkOb85fJmnRd7U4
CMcsLHHll8tAvJqwqQqtpMq0eWmpcxw4eLnd5LqgPe21tEZ6/E4+a3/791Y3J4/A
lcVk6RBpf9NMS2wCet8sZ1qcSr6ha/DOjRvZhIobPGM9G61H1T9nqUhfOyyRjHPW
H29T7K+6FxIffCp0CgVrVUvHy75cVpePTH7ChO3pT5+wBYPB4hjnkJabQ/dMrFWC
LC2EgSKj3aWe0GZeKkfYJCMQVKbQLUqXOTVAmAlBBSm8r0UlFUgY50GtTeSqHjh9
tFpOuPvlFVrx7d/+UGPjnz/h8Yo++6LtRLnJL2Pgk60JXtMu5Q7Muo+6xuiafcqx
XsBlwhkKwc2F3w9AEI5BFNcAlmUdlKIDR5yrL61oBctXpzjBq0XdHUApMChtqz4B
PVelUHFBqjp51JvqD8DQ+omHoD1nLoemp9AFmiM28obX0/5BkbmhRHlkRl7gnn/F
OxPg0dKDhbLAloHL6hQ5GrL2B/Z43OQoscR/6pPy/ikgPukWjDxESmC1gnw73nyn
Q358wYxnTMSWEe4HXl8CZqKpzW+R3EOxBqpXCvitakQODUYDl/ntACzFx+bXFs31
ZcMB94CpgOJ062nowMYdsaivYE5k1FeWlVg0yMnsppLItQYIOu/Xx9WpNUSGFEPH
AjZTFsEQsVrDcWfjQbAtjTsESOfwov6gfgp57T9z0GTyOingOdSZ0p6CPDCyXGd3
ZeHasdI2+jsIxRetoE1c+U5oLmKXEbxtjv5N5gU762qBDZw1G05ipl1bYG1OCK6O
OZqKMcxciMDzth2cZK/zmUB7R39n3CYiOrUxwtfw2A4yTgXImY2RAozOXfwHruOO
RdGJkzfTs5eMfnqni4YlDMtB0m9mtxfbnX0dvFkkVM3t4qVAJ2AqVjEqHOV+/8UJ
qLotxQoN/X7R1880ieDuT3jBiYToAOVrKfrDvh2RNo7VXo48Ll9Fm7kCxatTqv0m
onxnWtjtYrkHyR591WDl9qwap7XwVhoJAxKE/DBjFzwfAriO806464GuEE5U4YTM
EgebDE1bNeXWmXiWLCuZNbtVAuCWxXit8/CD1qrOMzZAU5CLvSZc5+T1U3Dqzi6s
qs+qryAd7BHfk2cROLQmYLo2CC7XFMEKP3texSkub+zaQu23KYOe4+0qupXFW1/m
d/zewgePuJ3HpBven/LiCnh9dHcDEGcH1mu2V9DqIFOzddciBkT0qIxqOoAQGL3J
brYFwVQpYycNpQdzTNRA08Gg6QIE9yjvVurdSiZI7CHQqa9dhGUGL6us/ix8CLKm
zw1Ae3o6rteMDdItzVqaaqyUEvnO67iPxvCipwVqWk/Y8FI04EcIx2fwra8bEStT
junvK9C6f0ror7ow1h3mL5Yhp7lo6f5c6HNkN4I8XWAeN0PpIxOc1sgDP2+74RUf
ZuwVAgJ8SjTpPRabcI7VrxTe0/xnC8bMQx3z9EApGOi64sa9b0zSlH9uC3TC9Y7y
2EkBVWVvR2JS+1GiOz4fkRpTIEqXn3JafCvab6Wgi2E7dtAaBKrRyRxgkyYXY8LY
S7XFHtf4lpSnQ3q7laFtZRMwGx2zvKKhKrFSmk4DtT8Kubz65EFQbOgA49MuYRHV
NzKcHkG/zdcIfe735LNCu/5BodQLJr3/kDbZ/eMgeif/j2AZe4OFENH/RHhuBMDN
8mfSQVw6vF2bDCSSAxxp4ow/31RBCbKrflsJDS2Hb+4I82H6Y8oXPWDcfr1WEP2F
3kKATJbfWnT+qBztUgvTSfVQmEJ9DDVIW3scxcMfaEPWkV5CfTaqI9aXdShyiU5O
KS/coOPBxxYmw3HwjfYu/S36VFkP1vO837O3Wx4KBx9vu5NkPJl0ufINphfEUndx
YJxcBBy1cx5nwMlvlAgUWdZhL1H60fujwwIs2q7mBe1hwSBN/IZMJrDKn4nM164Z
ukHhv5NK88yHqXv2KylLAsvD5XDenAG4/cY1JJOGLb6JqSc0t/hcjYE+74tMx+o1
10hOgr4eooCgvngiN8Jsbn8dgd092bTm/tBameWGl/LwzVIaYby2rzYu9HhPSV0O
G7YzKJOkvR0HLh56s4kyU4/1serZk2e+Sfms0NkFN4jnhWISNqTYiF+oPQqxCqJv
qP4msgSzEP9UsNuWDM4WBU6fC0QFFvE8hTvk1t1deQMkivUOJcg/CMx1Vil/eSyI
roFtOH0QcRxdTDYx2cuBEpLfg6nUpozX+YkUVk/XVr5eN7pY+IzY/xPpejOIMoCz
iOUkKS+LYMOKxwtocQ+5VQy6WZNlkQ02+OnrfiEO27JKF6YGp0FTr5xp36s950P+
ypJEzzOe0MsZPbH0SC6sTqmb653X1mYrP1rveR6TuCv6YOHVO24xR+UPZoFseC04
/3JLStLV6vfKWTV7S5caMpxxdyJSDb4t8j+AqoLNEHlmHnwGoQBkxCGMKnzByUuP
iTK0jWvt8eMO581IYHqCkswAVaPj7wELK7IZbrIz0eWMo31RARPNkMF0NG6Yazm8
bKg2+FMmuq+jgy/caakatrQl5hWmihnHiIiVGaqQTlPQKnIYz8qioBk9cnq0KpEn
dlyx/kNtIlpGzs5yOmSe6SJEaqNTxIIUevK/cpyCbrp6wWSeMYEvfm6bnsIvCh7I
fTKJLmNHAqPG7wH2uvuuuq5Pc6kXkiw2LyGI5PEolXEC1gVXhLbsUGnQb0S85ZHi
zKMgznjEeoQX/8WmWo3kulBmr4L+fX4dQyKyDEJJl5ryY0xPpOFyibeSf7Qxd1gz
vZEaK1euLcNH56JuN5GSjVmcDWQOjgc+wvPNLtmVHpjEE/YqqKezyXFOzqpTYAW9
8GlL/3MnzCeOGrEbn74AEEbzj0lHaAqf755oiW5JJU+rHtCGqb/nVtRiQIbCfgUm
1WGpNUrCG7osia1Rrp1sfRlfOWgdA9eyaEjxtStAqAbNeMupelKfIWJkdtkD7kEx
WsRM0Yd5xwHybVBGgvlYS/T2hFJu+dObiEOvSRqT1QpVMzZgisXh7cS9gAbr91y4
by+43CIyg/E1Yd0VtpArr5NwVIFkMqKIQgIv3qkkMW1RTxYUGn14/ieTk4l87g+3
Atr5sDoQ6+MjBM9Wb1ZBUXqg4XHQXUeKvwG3RLcU5iOLWr6hiSDSez6YFaSeDT17
8FiGPvuyS0xABWaNVAW8y5UQxsPl8dPFvbzSejoiIZsBXF/E7VCQqo8017jsbtBT
pkWNQOHkpI0ehe7rpf0WwjvEdNYu1DSluEj4C0lr0X4uH/meGBNGOn8fHiLNM/uR
F+CRt4CdsGpm764fTQSQKLfPuHqwt7oc/GSm/yP9Hwuvjh1KhV8rx6zOQJYs632k
YiUt0wADAbtVnzXuEIkd1GcvYPoSQty1px4rk2Gj86hfo4sfaRrrt/IoEfn8GjXR
XKc4baLU8qSnShuilWOeZT7Gt+jf/hxObXl0qNspA8SEypqYxQn6fUk8qUWKEQLs
xjWeJzA8M2VLOjtvic2dJeoHG7gZj1LfcZSRwAOoVBJ0/viYcSntEMVnJg7FiIgB
DvlQTIEWBK3hXnE9WI1du5Ou2lmTIag+Cd5PYbFI9HH1X2GDbil2iYrT+LcxOGWE
CijR0HrL3p0Qvw2gMQFsAjB6MC1bmoS3iPcS3bcVpbI04uXcFXpSqkd1aHcFV9C0
Cu+2gL9+AMjMkyri6yGWCUHYjzhrCwDQfwIGinA8MLmSlJXqVZ20n7ydp5hDFI1k
GXegs9ivOF44a06N1Vb9W3jus1JJ+Bjm7KbOMTlwPnvtM7ucdpgL63X6zGJu+ThF
4X/C+K5P/GtgqalLnI2hSD7rqVfnlsqZDQhNwB1Vde0TwRvV8aybjd0nGwjdJqtV
+Bk9uCpVjJo5JpOyq/lxF+IpDEUTZC9vg77GyHC6vRvgUeiJHIra7b9ffoX2Ko+U
DwTg4BWy7VyOseijAkFIVIW5rU2QE9Sy1z+6ziT75ds7zbh1cl/tXzJFEGcsvoMv
UUJmDjWbGjEtf80UcLUcCxLAgwXiE9S6+YaDLnTxWTI9lHbCMH/vDZreVfZ6mM6y
93gxjVDLiFakU/YHNsWBUeigL4FKVoNj/Z6okJEvUm16qeROWuiP25Qt4WqpWXBr
OHq0637LRiZnumhvgievqf5twY8+ixJV5d2mz7gDxXhjaBPJEndPBMTtU/c/LsQq
S7Oh6JUHr0uuE4Y18IcsFIKn1raASPq4z65qrn6eagmIjWfHGdKpvepRXszfmoyb
I44EBPyCXLGrQVNCCXh2JsMBCXvfEJPtDGLBo5UISc8vJXLp9U5Xb6+W0FtlVo3P
5L0EQ7LvZPF4t6smN3eIIVaUCgu2DU/dst1OcENnGTpkIp28957OoZ9x5BzrDxaK
TdctQu+0mfgjOjArg+IX8IfehsqTBtbUbaf3KSlzO3cM8/GrnYa/NzCoG9TWpkF7
9O+JiQBgRPHxFwEMktG8RaeDuzypEhCBbUP1OzuqKMJbBeN/XsQ8C/iwa8BRB3uH
sPywzWI/3KhXbTlX1OGWyOks7TyZy5SdKxXYDgBKBxk4B+wCPcbIjZuK0INwZ1UV
nmkNE01hK8AqD0UxqAU0cApgAkwV/3FHxagPgsLRCkNrd/iMyrzBdRh1SYLUsTbz
/z7hjwx352BsAXDZfRDycJ6q2WRbMbh2ujs1Wt83CIQzVFX+8IkwcXt7x/SXOH4x
y0DIGBFP0mlNRBFECCNtGmgRiwwmwcdR6htk6/9NGe53Prd6dazjBnA7FfqPhoRm
2HQdbtYC+RJoucPOge9Imc9OxWaWugNkZwImHlFw1d/HN+eJFTXpCiqNrrHL4Lt0
cxJVaUpehy9Ov9b3A+1GdHfaVm81noutYlglTEAJtX5PhvpToRt/w+j3efJO1UPp
rd1XrC8IAO/aiJ4OqGDV+SGit9TK6toSLRLSWvOEf/m4nXTgndC1OzJmzPv2yPjK
MK9fWTZrWenlcfoptA4EM2M4NXV8ZD7Ubh1epaLpr8QSXTnmZN6R269VIjCPXxTa
aXxcvdb8Znyr2GesXIWIGiDZAq/umP4zlrGZYNNXbegk/jYQr+I5tAUbUkqipP+I
6KDxbrekm5J7Y9tPEl+vKJ50E4O0kezll1NM/3T3sSohjEX/Aubty/FGLTTJ/BWW
AoPR7ZB+JcMb5P06Qt8ybc/xpDt2h9iKZByOwQzCb1xTQCtfVPc2yazu51p8JsRU
wJqnAnzmGTTsx6i0haAYR/deDgjE0Zp/5Oa+hlLtxQ6OoJ4VEUcL9tX/l+aSjLjB
ybInTQK1owYNITLoh0cOf/YVfI9rxE3TWWGXIXUyur4Wnzuh3LpNVMCx9E636jEk
PNwWbawKUSxfEeEH+SjK+YAq/UPgw72WAUYV5LffpDH8MD7FznEfDIyAy7z4Oivp
KW8XyakMxUl+fGHJqXKujH1THn1JkXrl17eIAS5EUn0Sgr+90s2ss1gOP8yA4cSm
EO7gvHbDOofTGmVPXVW75XnoIskMWDlERNhEuFHBhmvU4so1XbPnhR6GtK3afcG9
c4AcEALwhKl3XXHt9QrHs1m+gXih3IOxjFpD9W3Rlsz2PS1fsyWdUagK/aVjm3z9
lSSrDJGBZt2QB+ChPo/0uKSNb8bO/I9aXfa4Iy4Lq5+j5yhkgDyAJpVD4Nl4HelM
g8ptl4QUj/3roDIB/j5QM0IfQlcvUx8O6pzbkRl0oY77qtAwIW2FCTsFynyteqs8
PzdxbQy/ymLZyfts3atcSkjugIgtO0qAKR5ScOXvzMun4XWJrU1u3Q/H+kREjk/6
PrFkw8aIiorVlb2WWsJ/OwA0c7B1DMxnJRFdoIe7LJK2U7vc4gWGiQP9EFz0a5nf
KTTBpOSctUOpkBgtEZaiMdM4h6mrHQ7PGX/iL6KHLLjmgdxh14Fiem/x4vEb/mKr
ZyDhDYGkj09i3AGbJjlcafRF+nJtsYRArxMM2Vf8gj4kjDZpWzEKbkLUFcu8sEVC
SpEk85DMeC+EYAAnkHbMeV4BCpWJR2mV+iQ3LdOG81WU0qWzzWWf9WlzYeSnO9lV
HY730fv6eGImOIVgr/qLDaX2Hk7KpoCvl/AICtij7hWm4sJRPNX9G1AUT6eE5Cih
OUMAnIGiZMcr7Q3T1SMBc1N182kGUt3y+gIClR4rIwn2kYHWZNI3xR1sfLFbLXm8
kmczicuiu5TXQ1t3wQLXzv2J3aYbg3yQ4JSxP6wyOB+ChBJGIKdyYHHyrdbmlPX/
kTrj58Vl7lfhJpda5vJ8RTn0QFBrI9kBCQiAl4wFiT3fl7f/U87uiIVPJDe0NJ7x
Fveojun9FgVTFmOOEBuX9YUcuVwc5fV6im7JYuoJvVxwWbDkKsNq6T/NrUhZbdFM
Fxoe9JV5UY+AL+0TR34jvI97byIZxIb4En4fHs6GMZBZz9U42VeQs71tUICwEdQI
X+JJFu3pyOqaRamTrVAHrOiRoqEAQ3YmUQ6QeYXHEdPigzGcRhrDL5AK8FTWuMMd
p6fJ1GjG66qywD5zcwjHStm74wZKkTaV/d+cGfF3YbhIW5O2Ftx4diXYSUMtLWV7
2spxesD87G//wK5RAyYzzk00O3Dqd3ayEwZ2yU7LCu6YLGRdWODJElSTBjSy6Bl5
voxB9GVS34AuRtV5Ocae+Ktmyk8wzeu8abved8r/CMcoCoU18EsKJgUX9/NW9OUF
9+C2UrJawULa4PhedR98PaPMLjrH58NSlGU0o0ULP38gxc3b2hzZzGU8k+Lz7Xbt
E119zkNNln683LDChd1Q1/IoPFMKFwdbZNGDh+/4KhX2Fbp4WE9JafDsIbTdZauh
6B86pbGr6rYxfWjCNYQiCHDO6V0tLEe+Gs/8b6sBAebXbact5IfJML81Syhl/WJu
H7nMgKfZyZVgitfac9qNhEE3HwOdoUOWRofOVjl5tABNG14VNkl5dPfTzjMnmh1d
AskraLoihrWYTAX/nLjqugkfXHX61cYWEprbR38G0varIEDMpJR2defk/fVrAmxR
QyaQJy4ritVANbkuZUerPFCRfHrIBc9JogQD3IKvmaOUZYc6zNH//gLel1KmeyNX
kcsQyu6F1QwFf+BxsUTEOrfzsyU6mWA5Cres8qOe432lcXOUTc7aN20xAmVXWtob
qaWKFAevUUxM7GqrBh9/tGYtdASwp0wJ3CA9uT+DMOr8qiioHzaWQ+PwG3Q2tcEw
reFkRazSsf5rKJXz0hqGYELz3TmvzqHlV5YRbl1npVlObrNNQOr0INQu2nnU9OSS
ezmuBw5TzmgKdtLNVQSZ2QzOrhCunOJfjEqHIHIBuXB9Dl71InYLnSP37UVm2vs6
Oc3Z22zRnWwnlRG7ggW/RSWKvM7OlmbQLMRsCOwaN/GM5P0utOLrs3fh/F75dk65
x0D/GzKv6+qLd7yZcFkMz2725MIy3y2cdoXdoOHbYJabDKso1UCDa1HO8dTP5Phe
jCVVc5gWmiQzL5twX4rhH5e54hKA3S2QizRVjnhmOvis/UO05nrIPC7kFxT85fwS
E9S0ZAnJdJ9rF5IQfrYp1ZbnecqWp/rVCK/nOIwuF8jtpZKqfbygeFREnSaPJ7L0
LLcNaJ1FjoQ4MWXmWsKl2b0tsn8PrXw9PBxZpTJCLRKE+xP1VNpM2ggSgoh73oRB
XE2GhflSoYh9EJkGY3/dPZu3VjtPPbqRCGFrcUVQDz9KI9DaSQlR0jCjoZDMvE+P
SdiyE1sTGEHvex55ZdJ//SQYd8II6UMiyZcISALvpki1itxJhZgneWu8uQe7Zeuv
JTWC1CeTMR38+vF7Vyxc7bX/0mm+TGkgHofmESpCd0fCHn7QnxyyfBPF99Wa87Iv
qryi5IhPe0ohnobggsScfc8luBd2H87dJ4NxzlaapAgL97FwQdC2nA4ZTQz6IdJZ
bgnwkkyA2jJu+oPKgdfH+nBARYMEsE+G26C5KDPWAqj9IUTawiTiru1eHK6q1WFe
ISSxlgAGIbGAqcJmOVRN22cvJcoN31Jf9z75/h371TwD/qMXJTip4ndJ2DepcNtY
LEp1ceEB1V+Nqu4HP6ZeJQuQ0D4nHvSzKD3/Co7XAa+WfGmvbTSbNOSvlfA5XST8
vF3jYe5ctZvY2LJEZ/Nf8tVW8LfpH1C/iPGoCTPi7rrPH/CdxBORC9tbafF9qehW
HDEdykEStBim6s3a3tn3k/plrw3IVH2kbhrQd2Kwa5CjKNcXMlgBCDKADU9Fs8OW
p6CXXaofN4NsaXqjZ7QygtwsqZqsMPVzCSzNtxWIEQFqKlZRrRSzYc2S96GBEVQx
4d1za/UE13an6VQwh52xJw2zHR3eOUfM8NRMG4lS0CrfYVaTFTcq0Ws9bQsrggTG
XMKUf7Eyvbw67r8Cd93Vc6SB2prMJj/16hycn1xn7MsoKWdcn/4wEWHh7HiI3nwp
fpnKJz0mat9PBTTvi2WcQ3Lhj7jWAYhSq4K/wG++hrUqlZibZ6hXdWhzXIh2hDuo
/mk68Kh8AKVltOyIPmBoNfacP4nbL5QA/9sgWB5FgMRcgjH3D9anf2g5Nvqm93RS
H76zyYgUIq5LlNvcyaf0eMjJqMsfSLKeiS7OgLcOY9bGx+A4r4SIf8gambx8Tx45
T8zk2XyjRhV4FnyoQdbR+/SVr8MFX754ShSKfJxwVW5galZVVU+ELQG09VTihZNc
TSG/trblAN81m/m5WMHJfdLnuT0CeZLyF8MRE9UFtlad6GydIiODsqFovmV9ayou
povq+R+6AdcP02fgKNYJFrMDh9JoxrP93OGa6hRsXoD7SkA6l64f0ieso2r4fqvN
dlKSRy3454mO246MubGschGCgSgLtog+HL3f1Q5UtQmLS2tXKkRt8XnW8By6+oE8
aoFhcpIJTDDvLmRsXTontRCJYN8fYYPMFXBAIEDf24Shz5QjcLpVlbpixkoLISWM
K2YAvZ9B/KEOGWWTmHVWR9GukoMN6in5tt8qYn/hHrHxImukhcBBjDPHWFrzeX4S
GNi3XKfloYMKni6TBXbfNINAr0d256NV6gzi85ORTWiEe0nn+e7QcXtPtEoe+4bC
JU5gy1/2O2WYCh5ks2jndJb/1zA194tEuIBhLd27DC3ylGtAY0iPhLpE9dneObwc
uUUjfyupy/3m44GqGw/qplEC5eoS1CbNevYna0IgAR3SgP1n4Lge7Xni1/zTslZY
uPMgFDpUqTQjQ+AZFSbvinZwI02AoevUFT5RwACRF2PnQZU9wxTi5TlRtFZ3kVf8
4p79kpdIWqXwu90wm8JGjbbUNpGcmPbA/UFIUJiYtCTEFsALyFCw4G1FfKxpCLXX
lK/nlj4OgVnkzBMun/xf9VjBwOeTG0z/dQK2BIrXatb83hjyXlKyTarmFc30tyTm
oJI+y8DECCp/rSHN9XRSiyF4937nlZo5d/tEM9RbvF2bwpXpB/IjrKQhtR6IeRZ9
5uMtgJNDLQAo91UouKDDfpvM85tqwrMzEI7LrtfHRDPLbNSQ7Z2DJcEASzqfoHc6
62UjtJYO53HA8erPhE7g8+LZjTLzpi74ph+krT6bJA+om17PYKIFm/ysynKroVmV
aBlyLlUC+1jjk5pJrkRga4CMHJ6Yf2DJOQ6wmFJAXQJodeheYHB+SxgnT6RT0gP3
LyAFQntlXntQkXxLJNzpIKNvNBzbyGT3Y7tiEAOCXMRspFWLdZrmIuWq/WnEyJ3G
ZayULSeZ9kUAx95BOYYkC968QvRqWkW0HE94X5XR5/n0P43wv6dbM3lKLkUyyMvD
orCdNV0Ttp7fjMlRVIvUvT98a+NWEgKSQ3zAM/5Y0qv0Nz+mfFcnjJnqjCb/asRw
hoyNft/OzSLkVIRvMEZQE3L0bXceiRhaDC90MBJs+lhvAt5/m2X8Tw4SLC0zgFW+
w94kNzY0wK34Z5fpcy6ZfA8nLJ/ae3muqHyQaj4OsMvBIii5K6XpRaE3gnbqiYNX
wuLdzivKgKX1rr+PdYw3f41Y0FIeXbX/2CIXCshBgEw72GNGofF/mOeSKiKd+hvK
EbDGMG6GHTw+HpwQlHfRibvI/sLMumtILwS+aboaX2QH8qi6Jz7QYQzOJXJd9Ri/
3noj5qfq4WGnIGlCFremvXEN8vV7L+V/5R36iGXnM2EIZAG3SLuFmk2yg7tgd83t
Ju1c4ZU7PUZr4JLz7TP+Kl6mQv2H80NYOx0a6mp7/z52TkKbF+mZ7uzs8WMVuDRk
npzB3tGf2LpxA/UzY/spno26HSQDQ94tIGwuhMvkW/5pUbWs6vOk0tO2t4VwRlt+
UEt5DaBlHWFXblIIKZNSwX0hr33EvUeO/uCX4L1Pp3MwFVZ6C1gsRfdIWVpVMaVZ
ZHfcBzAq+tvjnScTGBgDeYFutwdfR9nGXBQGaW3Eo6MSgCmdDiJURRwgXiac7uxo
1OJ6Ei+aLnncrpGYZhL9HLBiSZ2N/O2xT+zPQzlmddDNVmEcrb0DSP4aQ/JYLJsW
k6Yk1RtCPQwaSIZ0LHdz8GimWm8qf8PDpu7eBYbZH6q8EksMVjbccxZG6O8yVJTI
VeHyqWrbYg6fl06Ju/kyPT0n98NqYEwSbDuoe6XWPGmmHsoMQyNmJ2Id6021BoBf
sRmn0dpnWVlSEdByr4r4WyzFqypt/n52IGmpxAGeBKYf8l347ndawqlmB3UFMSYE
1kmYCNmgNFuf+on2D6S5N7qwfOtkvOY7dmMYr2LF1jyNGsuoYrFGtOYV58rAjFmH
GvCFFrjXvVt7kPA7NMXA213T8l2OESvqhQ9J1AuQtgQOucPJpuQI5pt1VqsSpOEC
6JL611KN9xf87ABGqW8Pw3s18C4zQoUvQR1/9vMCT8hlr3GaNljNyDUGbhQk81cx
UIL4pVNiaN0rZviSaMe98IY3B1GNWDJ1hFdmtgMvSRdv+TkULZS8fBugh33xry+g
S/sJeobv+yqG+KrM2xLjLmnafkZCdGbSwsRSPZRk7gR7+fPu054zMvtzoC/rj39r
wQSpAPSzVM3D4zPUCvh456/Zh7anAC30TQaWSp+WSgEnxB4ggYzQjarjNQrd1lcH
z2V5gD4PLwhgI/AsNS++qcdHHwpwUg9Vp7IpNzfq9RXnoqL+JIk0CMs+wkdrrIM3
xjejdZdL8qNKmNN2IB4WgTHudUvsYrHKucymO5jHVlo1R1rq1rdyLPCOUJ3/MlzN
Z/2hANOfvamVc5Tz0Bg+wR8P8sE5G63BOPbII57F0tJCDghkOby2DtlGAjZiGD4z
i/UHfcAXV53bZUs5PV//PUXoE3x3Kl97gF7OaKhnr8/5UhvhYMxnimiCxYx+34JV
b0zbEQaVoiMsx6w8LkH6ZIJ2CS8y275VdgiApSasd4pDVi0ByE3pLyoTxYxjITo+
ilbx/ZcRjbKfiA4rCFsH21QncKK1eMcgOSslUvbhwCKA3Lt/le3ZRgJqxDzFeMvr
iA5O1Kcp4SkA9cwUFgabfH9CeO+bgNdhNsuSeKxz9vIsb2Hw8+LxFHShl2T3debu
htLyPE0AqsbrcjiOpFBIM6Z7u7lhH6zyAzG3UirmYKYXaMbRpBM0F3cvsrZMX2uZ
CyCjkQg9cbQkUVVMhelLt6/zRbQ3oRGk+oTDHINwlqrBCs0DSF4PHJ/RCaKhCjD1
7aXcJInRFBzj3MNek+y9dB6OLxTcXao3GosbsqMCBxbA3y/RINIWP07f3/pirW8f
qAs0pE4dMt72Bl/dmFopcZMoIXnsNeMHXDpQDn1C5Wh+yw6LncKEbQnNcO7OvlHm
GEXPCiECuLiMHI39s4vFc8HC8V2BJGZpzyWnH0rxBC8UbwbwbgTYhWsRnDx0PsCZ
cZjx0qiLeXSsYbvphR4IquU2R7BI44+Py39noJVlIqBcVMbJJ3tnB0JpfSpX0rf1
sdTevORELn/WejBGrcnEX6RUSxJwmO3U0mhki4pNdY+Pi/qPpaDQCwDGzhnPDTvC
n0OPYA4qikM8Mllo1PxhYvdbMc5fIZSqDpmTLR9dD7meKoGuECF7lN87xW600Utg
BWM+mPVBgoHi0QLMl6yQ393B1qgz6IVFWfxABEuzWRemxAqlSmyqHG+X8CYMT0+p
CkLPRj7b6ZtVKKJiAHq2Nu7sfbzNnnAFRWC6kdrV/6rHCGqY2euuhs/OiHBFKoZN
0J25TApCrhRePF0HBZNmOexSCeIPOGAJlA/yWMHOy0lc0D4L5UxI22ofywJQZ2iC
82s+zwal+9h6Bdulllmu7kNKRsAzaEZC/iBJ3249Wm6ngdqDYwK1VDzrN6oPe+WG
ICFVfhDMtpoFuaDu8vpr6BtqNp1cI0k+/7/Y1Mkr6vxG/oMB4+vjCMkLhWLniisc
tz/LuX5vi4/eLGDnBcUlx6NMuvUziWOSuTq2DHOd6LncyXaRl6acIJ8YUA/LnhAR
Ia7YWeDkT4uAKpb60IzXy1mVUQuhlOXzfvAYn3gu7O/pHl+v4rn7QX2jz18nqgB4
Q5zT3kVgLlXe1FS20dGLVxS/QK1EXmZK6jGRzN0Y1/ULMgD1Ae4+FQhTBL+dRkrn
i6ooFVFGnU+a5tegQW/diAAUbz18iRpa0HuGV7r0t3XNEd1JqDODaAqcJG3P69vF
aWeTMVVz3m9TLjaXMssS9ZR4mpcWHSkI6C7nn5cYvhnDjzJUHY2/u/u85IDtTwxe
b6WP3Lt6KbD1Aq9uATzqDSHopbb+2i2o7BTG9kvpIbzPxYAZsjU+SIEWu7PB1Q6a
sJ0XZfOTatI2K7BmSncPULuVhnMsNeodfC+igwJHyle10kkZBnjbVvXsCpS5e0e7
vX+pZ7UBM7T30pDGFYB+YA4E+8Yx+ancPha5kGDvYJVxfLcMYzgk2H0oLKINOuvZ
47AzcrjGBxacZ1IoTkZ8oRBGzqTcqVLaHhbIwNC2H+qHpa71SRw7fONIpW4/lo61
f8iezH+xVR82uV7uXJmvjZGb6HonWG4a1DukWhUXWmokwI7xUv3PqCCtJWZhDP+4
8fyek5BBcnADXrUqjbeorvUEnV09x4e3vf1NanyNHi0Mb8JgXGFD/E6Y7YmFHWwC
66bTqRPoy26Jov3pEO4vz4Z0d/3opC/Y+3eRutk9XxxSe88NAHf/8R1saCnhXV9u
kOD4f4SFV8qjnjE5AYn5u70VMScSMOEH3yxi0sjFiP5yLSRCQOneEAScJvYzwkF3
F3KLBsKqv2kHKE29PXVanFyYpAfs0SIi0QhGLeRXAx/a46d4S8pW8eh2iv9L8n7d
LOo0NV2D9hi7GpAnFDkmuxIdsUsAI8Mq2buEb7o52OVuTNjGajlr7WYmRTLeo4eM
lANGbAxWyh5ORw5H9M+o5s7BFj+/KF5r6WASRDNIpcN5pfs4PfBfxdjYlSGtVjiU
vpvfCIOKQ9CkQYxF41AwDdgKXib7hXk7qK6oDG50KrlrFmo/xzgmos6pWvBFFCdk
HhYHnf93JET/M9O40XCnrN56ITmyG5tD3iYjIhpsgMjr1b9NVTYo6CHnf5D4r6j4
ld6+uCO0m2JWfS/LNuZSy0DzG0suY37FRZlmv6jP7WHXcMo6hiCZUA1ZWGsV1ylz
COYpC1UJc0jkpfINMxzDASueOizpiOHydn3o6mB6SkJQoA2lVY4GYO8/LFgOLo0Q
lzsCIb0mS9VUcsXA1pTvcdoQ5L3IfklO9PaRKGObv4gbAcZdvV+q2sxr+MCDFPCj
0btKAulUFnxBmBbKeepsBJy3KzumyKQQvCe9J6hqVA4KmczMQaiwOjc6lg2yoMYz
0iSdHjdrqKtXYxOd+KKfDF4qCnnguB9tybQHxXOsZfYl6xRp9o/2OXIZyiAeQxSd
ptVJKB/i8QPt2+X+YMsq5Hq8okdp7RcYeZ7EYHPDrGezQI9HPIawMufbJrvKgM+e
BxzfWk5cGbGflBFKGgeuu6sR4B2jKO6PQFYOd2sl5xIyLlZ49XNkcxokyCKYEZAD
+5nbHYhIoGLHstCyouweCEmsmec5VjhTTqoOK+gKqB3Kn4YSJ+iZpQsx1f9q88rm
rKkRfdJ3tV+04i7VGr0L9wRHL5ydbps5PuOaE3AKmdgLzRAi6lSKJyX7BQzBQkix
qjT+ZGIeCIaa4FdJSChYtQCOWmMOMtQ//pxLbhxoFZ4n3R6XhXqdO24M+Y7fxYnC
0Flmxws5AEUjbG8UVsqXHegY1U2r85aJ1T3uDIPyeRV0+uVTs7lJBNouxUggDpMW
Ya6foKWH8Ukb7p6nOltSDFi4IA8FaV37mECFN+ytbr2jB6PfA4WoH4q2joj90tg0
Gd5iDBP2415mMS/tqkb9y3GiWP5rdJ0uXR9icwayfN/Pp68o7l7Fl8I8tuPgNOxQ
yOnV9BAc79ehZEMx0h92lWxOOuNLxB59DStZXA2Mot9rnMm+8Xof94BOy702w5O4
cPamSjied3IM8c3JPJkPcP3Z1gS5a47s7z/zcndOdJZ31Il/aown3Gr+vRQ2OoYE
jA+Jpg4pRdOyIlTgMhCct3jeQ/2BdvKF1my/um8ePx4XZTYXjCRZJYLVFJjyKaDZ
ayWwXTzrlgqPH3L57/t8LGVC402ASkwmVk5LfyXwynasgXJfEQV74gQzyxsZ7uOO
Do3wgE87CNZDm2OOmERopj/bEFobRlGXEMDvAncoRVnDOB39uopxQCLWcs5jGLf4
2Nxnw1bE/e5XxFtI+0/TRUG/Cfxo02GqTBXqA1tzcZrQDbDs4UXoM5J13PArUdKq
R9/AiihUzkuhvB7j6VR8TljGgMLaJEI/qZtCGy9pMfaOmB4xB0/7ZqvgiJPFnVvj
1sJmdxy1E5P2KVhqGdVuj7eiCJd2vRqhQljko7brz7hsFCS4EU3yvc3y6S7leCjF
lBA2UYYvFGnYmfs9Ni2nZZuo+KhIHHE9qXuFiTr14T68eXYfb6+RjabDRWIoGYbj
OXNpIac/DmpQIgCNOjgOzkoBBDRkQK63LEZm3Uf2DZ0+5q4npRMqh+iHFToKLqn5
n2CNv5afaVRFW+/ILHgdhYnAcLiSBm3nYO6mYV8CbJRHzBsoHS4WjrCIZPRLN6t5
iBhHHAdQ062bFCtGlck7NNZjuL8kAiIoPvj8kkaTowBvEnrjzb0RX35tju2lRWP0
1Yd5yWo/6QdgLGz3p3+s7aoSBJ6Hs40yXeo2U3FwxqOas9T+zPzd/xBorF/DRyLe
y60GehoCJHAY2/0P0p4ej7+iRibtImj26euYGRakCrh2tf5gFWnyO+F4pWEO8rkF
Nv5J/ODci+ltuOYzwAR5PNUNGqZK92urWHZ9sTr2rEVpVxUU3zEGHDo4+kLetWcM
oR6hKkukyZy4ZeDOvK5uaRTWB8cWe0iSDGdsSS/ujwG4ebGctynVYH6gEeAFcvvj
tuM96eWMzVCAhhNCdKqwhm3+6oxMvuchwPjApU9swXY+Q6crbDmscg0Zpz8aVNRS
ZzPiSc9I339kQxsj5bA8e0TdhOD9G5CPLjbEuMmvNjfuDDVKkhw8IeDBYmGgaVcH
R3tHXSLqLDI0UtV/OPsLn4D0EB1ECMBDmXZqbbMfnMENwMej176J20Td5OxfF/Bg
jYFG2YpxN7rTBh02stmer7tYMHkxIczbFpoI13QEBtSw1JNFCH9GzoTg/4JBL1WU
Ea/1j5/JkpEdd2xm62aZXNDEEdOgwoG90ogn/DdsujPU8JNztEkLs7/FxT41zbvu
+xJFtxlt5rbmNxZWH99+AEMEUFA3E/AJRo6w5MVvZVI7iRUhZHDXXk6i/P6vX9gr
pz34hxYsRdoRzRbAlTXmbq36c/BbOow19j4elfISlM7i1NjXPLEn++z4f8delGyz
pFN8M9CJiH1ljaRDOgjqFcKz45q+Okhq2D8WYnzieiHz4tgfTLSllZT1jDGf9R3X
bJZ/AgyU9dRs6fJx6xFb41ppojGE9r3kTYSaHjjGRVMnJuVC9yvV/n7ELd6OqZ+q
e9y/BrIX0SCTgJoORmDeGceEr8TeoJFU30idkhsNI4Zr31JNWoFZ7ivu8fzjBsv+
J4FoCBSRo8cQxStLo55i/pHYb7TkhSqzwLMvGD+W5UDQbsfb97xBigO/G2VV+FoG
GXc/DpHhlHBaNCFbYq7usybsI7Ufr2i3mIit6pUMlDgaPB2ZO8r5bkOIJmFcqing
XKZXH5pYlgLlxee3pZqREjA9LbZotlARzSnWky3c/9x7bnZLX7uELJZk+quF/ALt
2xblCuxUwCEPitsU68M6M8scImjno+VxjFRg2PgPFttrbqcvJav364HLRKE9uMYn
+zxweUsLP47XMcPf6SSY08ZKaRInpSynYuF4fauVZRxVSCshO9VbKzpzr1WY+V9u
QuhF5jTie89TE+eTKhWO3MX2UKf2DLqJ1AydPvCN1KrH0kIvxotgLc2AJJII9cDJ
VfN0qWEw0zJx3chpNiDfotmFNdeg624N99rnJw74eafrd5NiS9hrrMv06/yNm7QL
it0IPL3tMZDgULy4Gq4+BuIFTT16+AnYLGACBd6O8O5FwxUFTldJGDfGwCZmm3td
5D5VBuXHAosMlwOMCMkhDbXgM8VLYj0zqlFmBdGF3A5ZQLWEbqSKcJF3xgd7V85k
wjOtMI8BjbEow6QT5NxPJtFRQ4q6dgjk/QRKVjRBicj+vwHu+dG//old8gFghqrw
pMqLNuf6k1zICsDZ+sM8SGUCLA5qCSxlMqE35fDD6madhVCPfWu/ycagWSw4jIKH
ShbC5CnFzxnXQnCEl4O+OakpedD7xOwwT4+t7yAInmiDmEzt7RaF2o+O+D5GfVns
Jiyn/LnRggg+PhtxFSWt0DCDOSvo9wez5rPMM5Ut9qxRmSSyY7K4p5IcW7g68Ozj
rOAdRBBourksho/tOo1gCE218L4A/u1vxsKrJ0HkVWoqneS0Zu0esJbgHmZ5aRWz
rgdhVwqkWmGELSvhKW6r6q0mIWrPehGhY+tEWuw0Y7IEooBvXMF/tWfwtLZ+4E/7
a7s9LlQWEp7M4tFyCWb4MF/pRskpQw0TjvByTlRah/SM3Z+/zMzoghA5wtFL+8ZS
dWobS55bV+fh0xzpDqltHsngcNrdBfeDgVERW2aKXab84dfBtzfjIJy1T8c6uPUy
RZhH9YS7eTeoj6v2GIbtI7B5BYuoLF9cB0Zw4dAJYH7mUXXiSVqu3G1599zgYsmF
Zhk77jaVacjMAmNLW3Zow5gb+eiyBi+JD/Vlo7fE1kKObdQmeqL+SExrDaSzqpUA
i3/uYovrvLEOBcvRTKhZUwe470dHL1IK3SCmLIuU/odiSq2qLWKX49abl4MBA5Q1
FwOq5CYooLVlqd8Y6hWxd33vgArnfj0cy5XSooKzsccq4FW4P6NUoeuj8yThPjNx
QWU/aOLhxtj8mNSXoYTs47RVeaAg7zRwwj7yLaHkwqtlN4jK1s2acBvJZvtEvkbI
f9fHhurr5AoBVXfaZnSdaWr50W5kGVh42v8jWJfFrNe4q3Joobkp5P9koJR0wMga
RoeERNR1Ozbelp4rdwviJ7F0MqX9P6Gxri7iCGJXrZhS7HspVOmCTa4sxPCXy7IB
AXQJnJlBrhL4SMc76jJdMghzYK9DzQjue/PXTTTfBLoJUHewKkkfVPgfeQ4j+Nfe
mQGhUq9yXuG/pd+HHs41dVOf/KYKwqcCQO8FN9e+pQZ5nlNeuD1Og2R26qiVKYU4
tNn4V2fb9R8kDokpB2noYvDS0sfgyQooaa04Z7OwlUgMvn8toImOQEDRrj/MlL5I
7lgukAMhF4y8F0dk+/PpRwED3TFFVE/GH897fg8IYrjx4BCrANEKYeuI7a/HQvFV
zKA5znXS05zwsgIzjVF9zux+QCQrotmrUAWWTlRZRjSN58W1d7fCYjGUMgL94S7t
BoVAXKDVjUqXSMSmhL/ltZNgYADP2W3iFgaW+HcZNf+K6x/nn9SQUUwAlbQ8y1X5
78Nco7nrRNmzGHUet9bMvtKSMT1aGY3zdASHHkTQnQk0JmLFvg3YPYg+AzXjna7B
EJRwJhXEUWkuKn/fJzQTLvZ4vGjUn1AowY2umSR2NzyXMMshTfbdJwFYNbfwrAtV
+Fo/T9niKdzARy1nZMmZfS0fERBAojUhf/UX1t37kH6RRQqQkPVLeWpElrmd8KXk
sxVUNZIXt6IhFJ51NW7/sG/a2S7GKFmon5bwDfFEx/oF+KRgh1AkGyOdrdcNbcaF
x3jaX+bjAUk3gDo/RtVY9MCsPqkG9+LUAuwKGXF0Q+fuF984Of4oFzxWcZpQ88WJ
Inrx13ktaNBSiV2i2U32vxNd+L0yROuC1MNkNBk3WngURCO/wfcMqiS/CfX9TOnK
QUSS44/7i5K+jNv07JW5KQ8R4iNBHqv9elOxjHYDTyYVcncpPowbYAcwrI4tJUEN
5lu1vVBXD45Kp46XZ2YwPQbNp2r7qFsqHHjXbSbDz5lOnswy8T80O8aoIo71jH5B
hqdo8UzRP3tLBg7+rIO6SfqlpdE89XXOswJd0uVTEq56I59tr5b2M0agLF+fuJAB
KQxivnjjuE0ve9M14VXb3vBxErMMnvEA5m7h3FnU5PdcwzOHBM5dZQWpRyWf7aIX
Mv+2Sv+rgEO1z7AnB+CzXb8sn/DVXq8XgDXQHgQMs+tAutOEjvqc/QPTxjqKPePa
o/U7oJBxX1ygD93r33mT5ltQLa83UNbDaOMPIxBQJZnJQGlyTWsMX1Gu69NxbjZR
lMulpkna8xXzL9VFuaiHFfIPPGgfiwMvaxp4VQXNAMTvI1TyaWsfVtmQ5S4i6guh
sK/ZKxHqNutPSEPGgX4nhCT7Mz9xBh+sTjFtlRuSkkPjaXhZclXZFoiexglsIokG
pPO5THngOijvOxqGROACdOM3DtmHBH/wpKaFr4yhC26axXwZHsdy5g84UqXUa3Vs
V1TpQA3cAYoO1RwoFeuDcISDM0BkN0Xjz1dIaFtXVLkJNeFGtiGP9BOffyJK0tIP
KfsMI82ZwVYNAMXPZTFq8YlLvP9chi/5whxLMjGJuXLTAwXtzix9fh6+mGdwPh+H
svOImFiM0a+6FQ4A2XWHrLxwk9zAIig1NU7aUmdbaOOZ6iYrzr6FWyyw5kjCsMbr
17uWJ1o+BKjDeOU0EHJ4E0f+PgaXqefjCZVzTyDpz/yd09bxYQ2sRyFMJrBINSHa
2rAt6dGN4s6bRjBkJMBYw+WHTp0hpJimiWcARKRNwqmxnW7uKrMETM/pIr7uGApD
cc6FnHoNzl9GW5fbPfiPCdqCg9jr8KhehNxl9Jz+YYhTb2OkEI73W+mu293LJKmo
QIyouKCEjwMdkyZglCk9VyhCXfQAZ5HdAm7BEbL3NFVZAoJgzvoeKgcdLoXK0yYQ
QqZcqzXzeqxyzq+G+4cr+YZWz5crorEf9uCgl13RvteWB9SMZyDRY77kfhK5n3u+
ASxd7DJcoUFxzplW+Fw8JhOgVhfK6lgwuvk0ku2+N7OXczd0e3ftf9lWNwnOVlsJ
yFn084FmFHF14FeBfx0uFQht0mgZqXpR0WV2BNjjwYXw7WAF6bFoKLqkNFGzWqCd
XenX/NZ1GSZFDA9LYt4abJdZVtB8+BFBBFLfpeAF9xoJuvNsYCaTvOnq5PldQ51c
EIVzAJbGnpev1sqZuV5qo/qIKtMzoFmdGXCnkQHI8ADZD5vN6Uhcb9caSNF/vAuF
MUtsI45LYjMmZTEOVjtpcFr2k7RGv32fU+R98CefzWgoZ+kX1djXTz7JdC8BAaHQ
iHV5fJG/Dk3NiwUKCB8eRphIsuPOhszdzP9H6+a7HGCNOGVUa6okNLBLiXfKDkCN
gPCpfgRnvoz50dOazAeQBrVAqOxCYHlms0F+kXsLZ63JtPRgiqo1SK6AGMrjZB9R
E4Utn0I29dUJ/0Noj7VD6m9skdotyDZu+ODMEZTlgDj58+lq6DsDIIu46ZqStNoB
LptToVEeYk1dIyHja04yMWoP0eTUyfH7vgTat/a9KWSzCkufEufx4Irv/G1I/1SK
gslrwfQMLPWlI8Qgk16eWMtcahDlH2478KFgRTcKjTGG73+dHY1FXjSrmIEhA93I
Lvw7L7Xx8SpaspORsxOukqdJrZBAgQhdUKiGDrzmNGQH3tHnH5rP1MvDkyu6IFZk
ODM6JsTwbGddo40coFNJA9IZC+K9dmaEzA2+oOhwpxEgNnbsc0r6KQKqRFiYXXNb
595Iepfc/RTiMeayZg8HxHys0KAitz0zwLLJH3St8Ycmf3bGqzYlQSmOHFqUDkiI
xJ5ko8pZUUtROQUDGF1Bjm8FPd6hWMsG+6ZeWJiedHE4oZjvlHx7+qMRC8B21I8r
UVX+YQmBTQ64XiG6IQJ8+7HLr2ZvZ7PICTfK1cKi+ZmZl7XWc6lBox4GtCV4B1lz
vZpaP52Hf+YFGZUsEv76IR3VcupeBRZyiKrpNmlVLj3sQW8kIyy/uxgvynG6wVAY
cuOlA0OInZl5Ih9D4BjI7X5NGT3RPDAc68yWMSQtCQ9vRh95PlouIMAOZX5hbgKj
ETVMYoL+gn0AkdydM62JmX6eNlfnydBWAJBxyB2Zt39hcoNtCJnZg169IdGYivTo
ymHq0hZNQKgvZswpbueV5L0c86mIH19in4JjHiShq/yVTQ4RrotGceSm2t8TfChd
XicPhMF9v+ONKhyVsXgeSma3tlR0+qasHZOEwfaKWO34hDJBiGt4zERPfpknX11B
HEHUanrfbC1hqMR/S82AyTd9aGxYq+wWQaefb5wPyI487jG1X8LtczTakOwQ3Mub
Uml1n/URUVjxdcK9OnzJ6HXn88P5k7OtKK1VkWINYwEDLj7KElfiyu56ONQCrZzk
zQ9R5vzT14Yp1rKMv9OyEPKduJ+IClBmTchqzRzIOO08nfrqqQUMxQy3e9j2SgV/
gNR8QNVHAzBry9sJVPZHrVl0sd7z6mlFupCZkFOIwUneI1bYay5n6k9ZvA+KxvaZ
0I9GsSO34jHmrCz9/l8P0ggZiTZSVdGn7ikgjRoFmCRsX02EcsVi4WOUCtb9J9p1
cuFY8gbEzwbldNq/CiXvIU3EkHvZt8O0fgORL7AsXUc++No/+tIWHdzOh5jUvSbh
xZg2Y7voyrhj5Iy5ax3zj01FcjVj7KqHshXmeNTS9Eb640niSvt7hx6jd1vyg8gF
xC0HlgHsYEC/v6/xyF0eHctFQJGTxtuhQYb3x7szlzGzFEzmfrWS++bUWsx5yv1/
dW7Nm9O09I6zs78hUHFX59wdHyffD0KjCnxzalGgrcI0NvFkgO2vlGtsebW33OuL
SvlWLxtGNadPg1gErnKShS5q/bewM27VkHp8ZsFORWaJispztqKaQVseUidZa5ps
jGjZX2u2VzhPddBPOq/qfTxtvzXXHQxqBebwfcDPE5sip2rpa7op/6IjlM5YG9AZ
w78Al9nfvA4C9rhvZA0PisaU9NfkBK6Nym4I9yFrJPfpT35C14VKRGfK98QmTHD8
SnG8bDUb2YlBEpaeruy0NYuF7JzxL6BWhxK086djkii5CkKJzbpQ/06m92KsIAGp
tWq+MWqiPBQ6r1lURAB23+f0mfDWKKS+f5k1D1pDO9zHUwADzzvtnPnmXpwxYq/8
cXhElaDcy3MS7VSTmKBmuqgjEHvJQDB6NQx6cLRhZ4kP43okFglbJHY4Xs9NbbG/
rPSxfep6zOkzPsV3r0rV0v1OCHlNii5K7T6WW6F3veJjERtCbMS5XCPvaCwqHLla
lEqcLEzaRROQfbnXkJ8f3tiOvM9vQgi+8gSUTeSj/PrLlJpXt/hchFdvy34VcvYl
Q2CKn8sUw2tKookzwrl/kWphRiYh78WPhez3Xk69w+fwhf6knx96jVVoumH0/q9E
eev6z3gVoajm4zM7CBOObb/sG+77Zf6VxvDGatyen1CM0X8j4djM/MgdIrO1M3+Q
Eg46WiqYCcukkhwS0dnXwomXZDyJvdkK5bnmwA/caxF04RyamCzMJ843Vl8bOGNd
jrLCgrM0JEgQP9PYEIL3LUNvsoPtXFkdpzuShkFeZiQsIIcE3vfWRyfSp0onjElM
2HYS/RZV0awz0vvO8tDzS9qjw6SlyICsKujZ67QNPVccd+5wDP9N2GT6hJUfNvXM
Sv6Gt/c2VFnDDGX9xxdp6/XLQrHO9xZIM4ci1bk3FFQNHHhr8u4ubvr4zqd2RVyY
8J4XeytGb5lWsaO5di84fA/dRGMSNZCYNJcrGD1VE3caB7BoK9UCmuqfbQr98twC
wB47Y1OMogg+7sC5fzU97l1kcqucILCp201tXQJFe5MAOhKBmhzcH/7giojTdt/w
FMXHcJQkmpjxQvUm2qXehINsN+7xT3bPe9rtHwTSE7wjfe1b+12VvHSpx1xEBzsd
gkLhm9jaKTOw2VzX8/jVp4rbCfBtk0P/fkl7sj0rZBNUyaGTbpI5pRSK2KAtmXr7
4ndu2B9X4t3zJbwlW4NsMGTC194yEkNRXttsesj8t6Ws6J/+1ExDFQGGLRWOqKVn
Y8deQITYQ0XJsEKs/HjxddY+RcThNm6SFJgw9nmzUTEJsobnLyVUoXf+G0DN1vDG
ltaV2fr2Z1F07WgIstLI/7veWIutUfaR6R140KkPNTf+qfZXwdFE6SKlI4qoAlsh
o6lkxuqcwHA7iRPFqkyLBw9TKpFeCIqLi2RFe7hySuaO4YJ88aWw6EdOiND5r1z+
AhGCA7o1KVUEBrIuiz0rhn0drr3Ux2mEjFUigPxng9KHOzw/8xMovkxyWAP8bhii
FICQ6V6JQUmIu9pc9yHqifSu4PoYabzOU4v4hWVgpsUcTJkk48XxY+9so055Idsp
sb8Z6CtctZHPtKVoQ9BeKXuo9qN7S8ytTwwIxrC/I1weBlM041PTIeh46w+a84os
CDHeGxGXW5uXt2hwZMbvwOviMfet1eF3pdRGkCm8wwP3hZTuREikJPWXlm+l898q
aFDMwW0WkpzfxnTGA+p/e50wTcqlCnfQYvuUZLS98Quv2plenP9FnSK7QxmXLrW3
17YlesrpGXN3IRDEQnFriRKRK+jhSJz1AJawd1BwvXWseL5dx6mGKO7s4DTnKYQw
lGJTnnyd+jSbgOBuofZ1OX8ecYjx4T2y1vqOJf8b0qUEohFyLb2HQ7x0+p+n1le1
m4bxXDIdhr+rhUlX/qlKBbf3smKoPiywH9lXhUr127oIl4gJdcfSMXkwWWA3D1LG
boL2kWUGmquhfDw8jwPi1EqrjSblREnQDmkO5bVhwtGCZ3EGAEymLvjxVvwNJdKI
ZGLCENVtkFHKT/dlRrWvsGpCBQqvzh8RqBCl0NWKhWEAeekGRwKDinqThWNCvuKN
ovBchFT9nvj6cObx04h74WwPvQSogrdjw0VOnF5wH8OL9YcgZWEPexgEpelq7A0h
ULnTO0A9x5Jlpv/Zvs4VMjAJlzOyt7QS9BKhRShMH1xwm6fU4Ym1Wq0LTwgzPFmg
e5Af6ejIdbol2GLhmIDOb8qUWbvPxzK/u1/HPVH6nJE1yDBw2zkUmaXwMe8aTBUU
99zDrTwg0tR4PkPcRqxdrRl4Pax5raAhrFswCsKGfwX6Eeg0O4IuT/eFulz00akm
62kedcnzOK4lZ9XIH0x5jryage/Ulfm4nhBFhi09zh8h0SjrKBFOyHDUjcbj9ZZ+
nNHe1nDdOIO62gDt/HVDLrysFUKNvsHEDxURiySebLaGVVhF52GrzTR5Xl32PTJR
85sj40UBmMZO6x8lxGx9e9iIuQ3JFJxsMVkmeOZPthltehC6dgploQ29D8qSy+0h
Sm/oQco2xw00LbGmVTByfIonwGFcpUR/a/v4iqgIPKN7rH24RPIy6XYEJdUtx3IY
KwrnTwzSYfO71or47yQNt73g4kBefMOT5rknnKGgq8Yk7dzu4dqkVAGMreTc6mpW
eM1UwbFSAHWkcs8y5vGRqA51uDYWjT+R8q8YyJWLSkvz/OsDaCfsdrvjxcIIkZ4W
8/CM3YLrSqKhnK9I+Ys2w50Ido5WSTbXAKhPPQMCgC8E6fla/5eg5/F4v0q7L6c8
rA7ttdnfKNQCMiXvG05x7GsDG1Pf5It9mnBGsP9QsWp/rioebwhMZPVzSZXJ9QVo
9DaZ08e3HQmvogj0qmr0rH8z59kPgwci1RDsB/3n68xV03bZ5/Flu9Uq/zAiT7+/
6wl3JytelNEvOZjpNnSvY1K4ub6sy4MBExBzA6a/fXov6cfBW/SvdWTh6LCuR9lm
nEB6Q5/+zov1VpBcSgUHZ9+7jgpCCabHHOjGnhI33ZGQuE6aiUzwZ4jzxh9ccj5t
EZOFOTbnxZYly3EoFy0yezU30MIyjmfRQk/Iz/tCyYcSnKKnQe9LupmRMgBJLpk9
Gj5xKSIPD+YuxAXpz0nBItmr5QseAn0IQv/k13opEZX/gOi7GBIItGImx/k5L6P+
X/W4rlUzRjNXfBwEaJIGA/epiKhJ8vKN1dGS3aMjvpzuZiNdab99QSvGls73VdHx
2nbMD5grwd9GFjvFPyNBhWgfTA8+vLnHr2jnOsNjVOd2QDAPa+wtZSJZpEQaCKWQ
tFsFc8k4gv9QGEp3lLZsPHNaej4AFWAHeHSSLBbC2EIt/QyFrR6lgUiSuqS/TT/o
SS1h3C0iehyabq0DK2OkHPXB/4Rm/0SSZAcVeQGDRk/EoCvyoKRfsvPO9GGOFDjg
glOWtrL7t9kK/bXpR3cazITaKWg3JN+EmMKOZw9suKKeVguO2qzeFOB8GYLLzTb7
80xBqmoiDwZZL5rJ2Mza2MLYhn0oGR/+X+eCVnV/6aBKc3q3YKGL5jeNz4pKdEbg
csXjDQddLVR+glVuYnAroKtC92cgfQw0b5qbQYIOlVNRXpxX1UXa2Cn92LAdo7sK
qFwjP0yX0Prq23YMqG4g+bfozAX2slt6VvqZOynZ8HfdPVxEd9Wp4uCqSt1RXOTU
7+qfM8t6X/gK0PBarhEtCp0Yt7OZWgIThCoxMTc7yptacwsBMYMnUAe5MAVt8ymN
zUQodsm+zzfzE7pXoNhh5CcYDlrbDALCW7oQT4+WpXsVrwx2xc8v/8Mc50NR9oIH
DfuJds5npouXLhikDOq50mAfyLsRKqcxgBwYOC5fYueuwKx0nZAWD7Oxauu1v+fg
hOJ7X4EPVDK1px4Xu6N2NaO7Gg0bwJop3IB/Phu33CQbDGyg99Ku2JVSUn9yKkby
tTbVRJLNd3Z4BATDl+JThBZ8ajjadodPPaEfPHtlEC6PExZV9rhot9LWvJNWkbKN
iNNxRk+v22r+zs2ydBssVIjEk1/xdu4NwtbhBhses2dfHzdHBI9nep71IA2t4b13
e2D5fbtwiL/6ibps+F6O+7p6Fe+ggKRiJ7h2CJUJMLkzfHnuflnLljKdAsN5bANU
2SsyIWbs7jRrT2GgaTUT4OIxeiTASt5sRqWfaxJoK0rPVR/UXsrqS+UUCO0o4pxx
KRPa1gbVNvH0ani09L3xP2kUSPJK6qjCeC8BWKLngbE7j1SIczuFk1mBsU6JyWUo
0JIEHqtzf53I07PWlzy56+EDhjSNTmJfhreSK7gTzSBjrqyKqsIysocgD+rtfM66
ftZDE9OXuo2enDnbA6kbbgybsJGBRm/SXIFUJWh3uYrW78bCH0qLgdRFXQC4l5zs
a7CbT+KSTHTt0oUe7aiihKM5dXYcQiKcqAf2JvIPpODcgfdGLCsQoSGu1uZRQFvW
C9hQctkPAEkX62qCEtGO778/pL7f4UdD4w6IR4iJ0/sEl2SkBl7yCnQhQTKvWkCs
l32N1z8iT1lzFE4fP/Kugo3a4wc2V+lXm1CbfEEODQ8x50EdKspSl2X9x8HLPmc5
/yLWj4TfZRr8FjrUdkvBm3lwqqp1yWMCRksMC5OiPrXmOAtrfLZXjSUmg2VsF71Y
vKtiajR8t2M/z2vMaH6GSL0og/FSklcrV55itFSROw9iytHsetCNo2Xc2D9tOtWO
e5skX65g8lQSR8lz2FU9vCdeGDhy7kFZr9RIa7o+lzpqumnWqKwRr6jaTroJwEtS
2sknILPIgQVH/s5FOkZQAhAhb4KUE1kUreErKYsUd9RkJqVbOhYSAv/qCm+ZnCst
V+diyGs/Mx7WgY6yDL5vYAdDgxo3jYtO1JNjO9rzxvRBYgFKTQOPxgPEwgTEXxZ6
ILhRyQlDakC3h2aQE/X4/HYBjl3ItRApWqjaSvUN1k8dUOBvtklXO6OhbDGBfR88
LYE6v/brt04BwyFjvtzhGEv7ufiaQEtciT7kXp/e94JE8tr0rp8zZefhXTwmU6Vd
0mjxKiDgK0Dj7vHXai/8xbl16XklNUoj+U5yVK4GFhjHtYRfZ5xBt1p8P5wS93JV
uDszi2HbdPSpLpjUxJq9wH6TmXcb2nmk19bG/BraPxQKFfW/0C86o/M95Do07KQZ
H3IoVxz8ZEGVYLZe16rb6n87tgFyBJgz4QfAQKy2/eFYeTljGSlLdoSL6RgVq+Yk
8U8iMmlJhkzP+aBsUYFAqA/bCKQKFQz7mJZ6M8sMTJ/S3EUWYdeV5znW/brKuMDq
uxdh9VKyVVmB/bDi5YAlMd4Cma5hAW12CeQAIpSc1gVt5Qz3MFMxB6S/Oon5qmtB
u9RRMwIinoONh3LA5wjCrer7qiXkCrSuEF1eOm1YIEhH2i0yak1ZgBv0tF4z1DAo
q1+n6DTKAfO7VCC0c21xDnOAKgKLjKiljt7yhrUtUhql7ZfyVcaqXs05yV6Xp+m/
pgQ0xqTVZLyj5pbCijeHDiRFEZigj+bkTgPJMZQvQti/PTRsb6TJau6Pl2NUcnbJ
ABWy+E2cLV8pfjnmpQo5hpn+HXcyJvp35AIMabGJRYVPcBaeodeJ1OUi2PONrdmy
53FThtNgMC+ppqMluTHtpqpsCBLlFg0xcg/nIP7CMPe/kcIpyZAvuR+FM8KORaBa
mzJDavlFYT0EOsk0Cs1164NQdE6/tHQMiDQeomvsSLqwbP2l9fW44iPllV52/B5e
s4Q5yufGKpzD8o4A3ZAsmk20gsOZFZKcE2LXpofrbEynVw3TVhkLWjsRzlOGYW8Z
fixhQ74GdbgmhduJ+AKHRUMYk7DD9zh7FOtpGkwD8zaR3+TUYmIpJbbxUTBIbkAd
oqs8J5g1Tb498oUm7XOEJ/eUVeigTEdlR2BoIK7po1S1HPojUE6suYcFYv8su4aC
tFo61DRwH6yhwAzG/BgPNqC2TQFn3GOz3qda/3rIBBw/FX85wQQwdcL2cqQAJE/s
PKDBnq1VpmMRRkLDY/tChC7DrXRwXwjUwsuw6JoxWtD9/RDsEwhCDveZXs6gBEh9
DwH3O3QP/v5HS13ZUqJ2khFLajUuuPBqgPwKXY8fh5gMNdAJ9PolXKwF1RE77W5X
C4/67HjON7ycR1I6WDnhsxwkWKU3mrUUWi1OFeUQwYVNMpBMd3mRaokTGwrR679X
jFy6nV6GUXpKgPYRJBR/T8a8VpJsqa8ATzviyHhJp6bQoV2OY0KTcwKIRitWagcb
HzMmxnPeWTJdhoK/2jNlEgn5WiA56dH5kfscSHCa7K3WsrUoCqRK71WozjOvFv6L
Whv5B5Bexm0+rmZ1D+apK2zyUka7ux3SRbXYMGlq2GuOklXvrj/kgUakyF0j94E4
0csehpP6c85LFW+xfVvy5SM8dZAwjNQabQnjgfIeNFsjfAwQGuLvGNs0BT2UWFNs
VOY9xCYBcPmy3rq/qFGuT2YB55qJtIMrVeh+SbHFaMmLWiGutZB/l1CGjR/kh+Ch
sM9RdLElxRxpDofDGnMyIB4DrCokLASm0eo5k1TEInFqMwQKoDBKg1Y/qX5AreLD
Uok6M7+iKPDbvPPYSJNWvm8XinQ3gutnUK064FqU1pAHvq5FoW2Y7mCVXPKJ7Ycu
4eXpnR5gDTucvAdsYOGwVI434FnlnJ4yafszpfrt8Szh0K0fcwxupo8o9fL8s6uo
BCcF46G46YTlUn2XQFCWEsdc/7CJxYDkuzyq2SugS5SrML9KV2Bgf6Ierj65taWE
+nqOSfsoXdubvfBu2hC1Qg+6+0MUrGPCQYBVJnHLRFTfH4Ep9VxmD9h5xXZ/1YS/
uxQmnQbr/wDLhFQU/w7EALqqloNA156lbLfmcm4rLMwD6W/7Zw9b1TWBob0Q/kbm
qJCwcSQmrhcZIutQ7bJ3RjttivqVdGcA91NFRxrWjUz1INwGXe3A8gwd7rg8+wJ/
NEze0QJycGM0k/dNJ0Y9XWOQFVsXJXBs4rv8hkqwWR9wrTNSc/zD1OPDGmdYIALt
GrZij9WE9A+QtJSAc28d659nx/JcANCQdRP+Khn+m4JdLz6clnkwvwJ1nFp2YIfl
Jgv6n0nwqff61c9JKj0Or3dAezRm2lbRB9JlLQJ4jbEvs85JRygSmrRyMAEuaAzU
OTwZMwLAwQ1/e0FODRbORtxn8F5oSSTs/mOsZIiAKxqc5IuMqo+U0RQ4mI8ASnEA
Lp3XSHEch4aQsOnot3MPdp/1gFEGOtBe7TXlz9w6pCYBoctDJEH5DZHAvF0iTfJ3
REfue86aZ6qLoq+A674NYG2Ha26WTd6youVHuR+AUPogG1XMGfVGhy3a0uGPQrMk
woHQOGlndlQgL0sAmPMBZt3PZwPYqacp3goUmWnkxMCFiJ3ADUoSGKvNPdQQzawe
tqRqzOUTSnvzGmRYxG9A4bBxkjoz99av9jhKHTeR8z5Fmr/pC9KO00s6nk2DNmJi
4JjL3CHgBjGIBMTckGrUX2c6mSRSV0OmuNPBMhkJ6D9RvPliq+3XSfN8oBGr4O8l
IAaYW3yyIqsibdASsOmK1LMTBO67Cn4zCS3MKyOnBPW8Jp6dL20W6NJtXdL+RyhV
VHkgnYRqmTIJs+ZFO4kfVn6t6TITTXFGWxZy+d5wrWbfpHwVP1Ct4HeEV8ZrU9qS
KZENEUh0sHGKthvjgINL5c4N7JMw/IKlKRxtt8XNzEBOIsnaukVDsf9MRfJ/njsy
+sfEvmRKwEjZmvrUIqEz4tlndJA2jBztKbq6TvWeecS7Mms1iUJLpqjxq75/muyc
5ob2mw0MyK/BG+/zTwQmdeqG/+S48hFGso7VYT/djR8ovytgsKjisSP+mDBYXe+J
9ogy18jQF8D8aSCAi+7IXDbcbSz9ksVjTQqOriP5a2Ztek/mZsua0LSbTut3qzq1
9oci1EaraeIlQCZMHdelGWVDceWcqkeQs+KP2fqILXAgD2pyI2c+TtSStPbXlqfM
ILruDNHvEXLzOEKwx6n6ue7jTZV19md4vCuxBw+NA0LgUIV+BS+EckQ5utXbS9Fp
YTBy18P6uWonuMKoe2mfVXPZ7cs6o3b5UDkpjRQTqSUE0XXyIjBThuC4VdE6dL0J
VA21G0AV6E1b2Z3nHXKre+bEKoAa3uwc8ENU5VsPIxy7+YlQ+fLleUK7U3+5Nxj9
rb6dZ9I4t3k6x/9BLcj8VTQ2crnVpHhPqkCsAIJX38BE/R1RRbrZRd2b3gXuliok
P1hPISZIz/NbVXcYeZMe6mKHTi/qXBhzZ0g7rOvsE/h3KLAQ4BRm3APfk8IkU2HL
S7PNRvz0X/Scw3LFXYQ99MgCo2/vZ1oJ4MHtwFD70WonQT+O0KagCZuH71F48rnR
e4LhOJYJHbE2dEbD7uzF02ZsUp0TgMYwChfGZHU7J6zR2YtUwjSxPW1y73LWlvbq
hXGbHaKj3ATjQO+64tvboao3N58tSmgPoDPlDoq/arr5FsdBsTNnfleRlXe68y1e
MbD9ksg42o/xqdVrCNoTu0WIRBiTnxDdAkF4RBvxa1s8YNvB4riIK0aBm0/ncIF+
RTfYX5Yb5Zh/q0E0eMGLVjDpkMLlYkAa2HtmQ7g8qSRjTrmYGUmDoHOfEmRWHbs4
819Q7LmY5Fg7MNVjDYLSBx5JHCgA9Z37h12TRoPpeGm/hctEJX/uKPE9eMwy1W47
Jqaz+g+t2ZWdnB75PkC5p/R3QIIvkm6aZU5XGKkhIpvq+Iyiq+Bt0aIN8Iv/JXzW
jNTfqSUPSVLxMl/arnA1S0DpeVSiK3oKyboj/Cf6rjr2BcSAhIafRGXKbp4yajN8
tb/XRuSSGgTqLVPWMWu7y3x1NdruZraMIwMLz5vLn0PAX6oiML9Ro7k3VZWljyx/
6/bmYK7YPc3Y+pJTsxpi9PRufBLyfI0Q/ZhZzewDDM4I4GdP98m+/oqrqLofHFR0
gSpPPVurku+6yO92L7LYcH+IGS/6vSd8jUzncPn33gyy0ciadohcxszlG0WRFoPF
p3BFoxnZk6VqXHkFRRVFhdRb8AXwzzsAiIcGqyMWI0cpqHyKSmbknoacr6au5Up5
NX+JC96KIvcaCj0f/IzZW/ONUL/SqwPDc8lkpbDqDvF/0WbwafzpjFcWjYdgyuUD
DVf8R/SqzumOeXJG2mHBvhwmyvaHAcdMYlWNsft3seTVQiWeuPN5JrTR0DDgpYxw
2tvDWI7vrE1QgIRpUqPaQiLMQYW5X5WVyQsyDgaJ3Ovk5AJDeSpYUWkRnpBgzbc+
qEhtglG+2UJMVwNxpxjA6qxo9rj5Wpp9ta3mLhK/2GUxZOyFYm8iiZXx34m55VMX
/ND0+VMH/z/tlArwCernR+h/EoWpNcZQQN7DYg4wgnVtrsAASf6KneTnu5YaGnqL
DElwa3QvVwszWqhEEP4q6IM0yiEqOvNXvSEJ6YqOczjLpn3CRjMfN/7mp6GFlelW
zaB7LJueqMNPFSYH5s4sS7xSes7dgxSGJPTMxk6ABr7zLrLNjtoDXNmF04ZxlqcM
dJvBjJN1O+u3X4qc2cdNLGWnoJAabnxdMp/I9L4JUOgzuLY5UQ1jGaZ/IoVHPuDj
962jPzaot5xA86HJLV2jNcrzLwOYCRNZ8DyKfj/KaP/wLkGu5tSgYsIS8fdHWr9f
AUOgi0swhZCgcYjMIWz9p5+nLadQFusZ5w9OGLjaX2XENphb51eVL7PQbCYqd0PT
U0r1NMD5t06ciLa9dP6IH7O/xkvi3P6xkVlZ/nj45DQNpQpCFrPw64j5VpW7GiTb
vjdqtYuyxc5jOAbHDbm1Uye7IRg2HHH2rpDPngS2xkh+KKNd942fL0tb/EqLMocm
fnz6z1A7I2jKrgDDA5ARqOxRa0DBL/NHA5FZpN2O62Ru98re/ZxtdZ6Ua6e4gCxs
W6XLZkWoXGOwPLivjmzCbdtawjcAyN0JWfwr1thfiwTd1YkK2ZcXw5xoufjQ1dJo
sV5O1afL2TbqNcxWNNc3+Ux1Vc6dqs9wU5XPkXLtHxTX0tD0nxTSdfv35xelIZyU
k+ztZCvOFWGaWyCk9+p/AixzDu8e4gtx1zaubhXYrest1Ym1aQkic9Ti5q5EeMym
B10IedG3nEn1/WsCtun7/JnZSmjKHNAn1qpG6vvo0SknVbWAI5mx0muS+isfbrwe
QzdvJtgnCg3bbdXzb9FhWhI++8zE4v6i9W3k/FGPoqQHrPy0RZmkSTw4kWVCYSn8
fSijjby4BvS37CWkOEWwMbcjsNs8lTC1iahRr4bPbdEAZQpXixYpk6BLwi/P8q6E
hqnYP+QeznSzieuClGujVcuImhHUkxtzVo5sDGME0nqLh5jeFJ2KhppeiZnGz6Tb
TFg7GM5MN0bhTiDv6H2vZwSxFynBRJiLgeHbkvXHrN90PxS7lVucXq88iG1zPlNJ
AWB0XNVYW1vscnLmqWHHp5z0EBDQJVwIA5xoidl4lSWRn7ITPjlctxsId/eT+WE/
kSXXuHcEzaxCvB6QDI34VLTej1h3IaZtKhR7KAM5ZaAOcAf/wz6NikmV9E0kp+qJ
cVNkFrBqTANxnMQnXA2nFNoDz7Y1cTZvtXnq0nkCak6ab+RvVeNIG/esv1X5iyBK
DCb+A1AkoHRfgEDt0o7sNtCVtpA2G7bLSpafVU82tf4OVgrji3TVtjoFi6hnVxu5
g2uBuFaW6QU3wfezHNHMKK1iaOrKRGEWUDvuU4jVIpP6RosDsJkWzSg6NABjVCQE
C17ix9E5x+fve7lVylW2gs5NDfmHYeC8qG10utW+mGc9ZbqGJVkdoXIhvFdGSnhN
CmWu9AoRioqrEyTKVOb3BkGYuJxMx7qSaFOoWhghtYhyHfPqvn7uzylQycCbytK7
7pT4Clvk5DJiWkGCZhs2+I5AIJZq1roU4GP30elJVZQehl94mNtK2kPEat7t7Xzl
Sk8hTuOgCb4sRruKQfIJl9fwX95SAY9iu3osjF+pkWTBSMPFXQMWT9A+j/JYrPnj
VpFtf+Xi/Qg2yAU6JP5LHgJTlg8iSsX/zxuLtFWJyjHU8Vhk8hILq2WUh0dSXYkf
XEB1JLHIqIXYsBSGghw2nAYJ0IXK2A+MaJHTgVszZWAqxz8ZqGb/+FxPh3cN4MlT
BNlmZ9tvCWKurAkrK/c8UWsesiG+6HAQ+MK8isJEIlkkcCEyotaoxYmBnAh0v9Lz
Uvd+I3qji8zpQO0gRbpNMhOV/K75uK1ECnZVBTnnKr6cKu0DhhJqD79Uv7/MnVpc
DKl5U9emzROBNEj4uCX3edYjxMoENKyX+uFggXa9GutgUjMeaEgmQFEvMNZ6OaYE
h55Rhz1gz1VY++UQoOnO0NH9w1JLCrIKZ/euSXrdVfBXv8T9d/AegQlrTwWbij/F
lp3hwVU9Ldbc/PQw0pV1C1IAViOb+TFoxc0qQJTc3DPK8YHAjk2tb/sxxbfwI5ff
YD9Xr+/1MK8CAmislXPOO6Hq++Xf00gujyFCCavmzQX0vbP3o8ysEqp8ZVo4tixt
WnDx7iEoD39/2IbnLGpMW7hLJrfx5T4TIYJLg/qtF0uqNPZHJFnzTM6e0zxYUU6X
qreR2pIIyf1VKkmCey0QH3uyN2Je2eAaW5Hgoy+WOHctwU20ft4uanm9U49iTRUq
MfBENTikeRv+MOmpL5h0mzhieHvo+FKyNNy77XbQmE7cbyaqONl67rnvI5+cIuGc
yQLu4sW4/77Eg3bbEHmyi72oZYV122V6STdsa7oC5MlJyzl4qGF2JjKXNVXUiqzt
dh35ddnoTXq4CCJwiaEQJ6OE7dmBTSWLYcUEJUqCBQu8V2DLA8aEEqAnIKcVusPf
DCC2T9PaVBjh+ZDYw8n2DHe+RTJBnIL6+B3j9oPMiMcCrFEQDAD0q0TFeMo5m9Cq
ppkRAUdydeynuou6FPbgpfP5gCCeZbrPv/431j82D1uEAwsyH325nlb3j10OKTto
Fyj2ddM8MUYCG+CThdsFODaR3fxOUITU3cnNT515Um5oBKpRUmJSrHl9X4TT4CfN
arRYn7GqZMhRHcZ+wvEJZSI/ytI+9NzfjJi7O+j+nTXUl/aF48Is7vlsRFmbsCLA
CDza2TnrS5Jnd0BG7pN1vZuwfuPzXOFJ1F5r5qUAMbxSB6GM1IhCkbgA1PKzqPsk
yizSXJB2/cK6VHiHDjkaTDk+DTyAbL7ID1SDGvw5Eeh90YzH/1lKt2CQkzZsnQC1
Lsgc1DUCbmz8EazPZ+HMgCKvL8mauUK5M5+MJI8d2Ma6XsYlstPGJofT5jgFrCLT
Dk6wvJrwRnai7aIGCROOJHc84XCrky7RdGFlQ647D1uqTE+DZKMOW+geDUOpoZ08
fSdhtYBzdzA0T+TcLyCu4W8/+K9R+jCcBbuysKEwlGfKw+/rfR9Sv9B+goGQvMP6
Nzyd08K8lYwsbIuOIZYNinpJb979Vv5+k0a4BwqM8A8TF1XRFiywzJdQoD+TwZrx
psYO6tkaPIco/gaU/XKzY1tdioz+jK/DE7EDD6kirUqOE/+lDCRQvjparqyecRnI
aFhpkcP20Ddo69HP+vHzNQVuif/W9pa6A/1SiSfhtaulsevIWpoGtagsdncBE+ql
NASoVlWNfR0F9iCjmqSgV33VOE2bEzcvx6QsjpxppoRrKHf2fHQejgqcflnXKS6o
O06LvbP15hhQ1iNp5MA4tmZc5q7Ljol193FDn4ginrKFC+TBTyHFx0Opu8dRv0lt
vVxt1fgBEtL0Gjsdd8h3MdqAAW2OYiq1l/My4QvVBGMDLhkYUhuS86dkD0usJ13c
nmv50mXr3s0VL67ndv7Gt8xn6USSZjKEQndeLq2lUnTDAOxU3Ilq4zzDC4EDp6TK
CN/Jtlp5jpaarCHlI4kw2VfaBXhJdgbHbhubL6oGOoBTBJsGBec+ISEgEBTkQmzU
kPfjRCMSbKqosdtiOSVPvCabs/vsMIlnr4DAiew+GrlDzV4lQ+r36cARjjEkizHT
z//i2JOG0SpeJHy7+O0a/Kh+6hOVA6y+3jRT+wFb5zztIfnJiWY17qtyOpYMFrpN
lFmNSWqLnBm8RntLdrWp7887DQUpsqgYVC1hz9yuJWRvhdm5yVppYgm80zOUrobw
ve97rOKA15ueBN1P2L4L9Fu3EQvYnKqqnghHQDr6UlqqbHV1RTq3b301vmjELkgR
VAxO9ndlywG1YaKq/jaYs3ClUnWdrY6HjPqh5D5+wnvaWSrTjrNKhEYc7hFriqLw
QXs6eZMwmGC858rxBPwrvIsJbwFOa1JhzvvTpowwaND0dXAcPvdO2azWqmZR3hBW
oSk3X+3NWFeYJFSChDA5bE68DXRbaMaWP73GFooxfY11J8/B62DHH26trOBALpjk
SAROctNnzQN7pTev1SO079lUBfXZlH8nDz3QNsNx+EmJPnvG55phVRPXZurmC5FP
x1yzr8ztwzwwYn7tM+Spe+SGQ9DwT2kXRj0zzGtZuaOOWziSVJFHg/o1HSiMZjep
fv1o/NOwzr1lDiTZEMzrUW5gl/ggy27E1IfqcxODd8SrIeVBIPyjx3Fn8CfSB/y2
54LyU6DlrsPv+UBz+cT9a6l+8ilQ113myB1OUYLVLT8d9cDuUOcBZ5BxohfqEwQ4
X/8ZS9neDvd955CLG8OtpzbSPpDUDTIgz7jD9FZXNfg3ihtleV7bkZilIosY77NJ
6q6pGw8V1VKHtO7mBU3CCht93wQcfBiZz36CsHzv7CEQ/5ucbo9FBQ9XP3ZC24P6
VIjiTFamh+c6RbOJ0VES99PLiUlSMOBaqLYNwGNdl9/f0bY8j2TFykNC2CMiVqnp
+DB37VtezjJaJ3oCFzj5jKFi3ozGVyH9ugsHN3oLvxSzwnciUUxqh1E0LDfecg/l
C2nEkJPibot5Xpy0K91xLh8z1ahJR+yce/+eKwV9W3ojVD2ZKrd/R4+QtNfxcn+i
Auz2rtUxRnH9qqOlOlQ68wGbeVn/gICEDogT12OnJJXC64/aRFzmd9SBFEUYslWW
/pu6kEHZ9LNTPi1KbohawKjNnfMwfG23+q+bhi+KpHwzbhsZSgneNcfuf7phY3Cm
jlcm4aDzY5xMqGcjdY4MPFRdWhv53EscdlFPuJETVWuWi+UVtUtq9JPh6vEprc+D
E3fu06v60GbEHXvFUedRQbvAjdc70LAHqDiOcXyrNZvZX0xe0Mf4UqKkpqWffCO+
dbKKvu9LY63ZzBoomSLEmU8ok2wp9sRQZ4ya5QUgmmvFsLolqdCW7DYE2M8wcVX4
GEHHTqJqYpdrJ+ce5PaxKp4kvj7eJmLg+XM+b7rUonZqV+tci0iBOQGrpQeBAcg5
XaHFOIP/1Uw+2WexepQ/xX6JhxSnYhnms6MdxypaL6KcUmhmQ0x4vr7y4e7VsSp/
yO0ion9+uRPu+RnBLiuP8NM4PV6jJ7+iTdzwbuIF/77Sz9osS4cSPcCEV90dB7ub
0Jfao3Cfa5o8M99wC9lDycmwYwcUgzb/OvX7nEKGAoSQojYJeWeYV3KCf6JtNL6x
k3Z/5dh/NPqs3Md05nfqptA43i9muUSgisk+gaoe5l7aFVeUbRs4tvT8P1Z5GwaL
H7Tynel4FvDIaE2lQkkLJuu/N3M3RbeoKxNbRKsTs6qpEoA/4Zx44APnwF/mg9sV
4/U3mq/CmB34i/iAGAZ2/rQnEN9oiRxjNjULrCBsuDPXryUu509E76UxpXDWBnvq
EbtPLQUBnB2t8GWWAWuS8rnzV6rjhG8HVVUOMugXAYh0R1zaIu58rkv71lWI1cei
M/x2I+GBxzf3wf/NGh87cxxfsLE/ciZj0yItRS0XJC9ASU73a6QPxHQgmWMrPg1h
gU9kVseMJyhrTjgG12qKnT3pWTOCcZRES5ZhIwCfWlHjmMza0QfmX6Hlyjgg1uwG
sAba746wtB+09kZEkNBjEHkfQvplzTxrJx6tXa+vXbdRLgt19XQNlfWxRvNMThCo
+qrZktjwCkDTNpmuzHYL4XzeeSkP0UmrJa/puPXAmXi97HXOAWAY+CULJP4r8yoz
5z3hRWm8M8cxcuE359k5cWxKDgGONawC30btKbPWKUFW7iyagXaMXgRsisdZVD+B
gemXpB9bwtFIPeQFqfhJWD3lVShwYLLJYPwXTsmKre39c/Vz/bXzQFGLntWm098W
AswPGEgFWXcO3bXHiHHmg21haUOznVPfiQi7aJmZuirZ9NxszMITdNy2DB4g/xrT
fOT6LkicdnLBv1359PxXV8gKhjgGjWJYJ8QdzJMb/N0m5DgW6aXnmFXDpXCnP7px
nmQoqnQrHVVr6N65342WEpzpSa5sEDGmSzBblyPsM4O8BsaD0pYMaFI8ASTtB2K3
hXmdx1EfrRIJ+9tQNgdNqirxIeSxxAwwQWFq+5gNEER1fSMnnf7O+epX+byO35NM
IwCsC8Qbsdhim3+pYCBdNQFyH9PaOaRLnHPf5Bhqplt8Q0/G8teqK/KbAgVd37Ln
bBTrZIHNfswNcGcPi/bL3HecTKGhTStatfRGJ8Hsi2RIHXV+7ID+J5jhIAWQpe86
qRKRUr5fWZZZlKVl9XIWJF+RwtI4G/JKLmZsCAkAQ/WYcpm/l5X84Pq7rs+wmyui
ZyF26F4UVnv3piZ7mtLYSLPP2ELc5CgOJd1cvS3Mv9T3v3Lt1u4W7UF7yfbGq44A
Ly1d2lt/JVo+d+dzvPFWAXYQZHCfEmlZyIRWvZLu1MwahnHci9Kr/NxMicC21hOK
ZaqVFKtIatN/iW2paAy3x4LeszwMyLmmbnFFn55aRmSrO0S2/0uvyfg9qigS2HHS
KZ5J5TD1EXZLxLH2wlRRJO8IQ2+mywd1GI66GIvskXCurw3HNpKN/dNTQ0E0eNBR
5BgakcTWYCDPajZH+/oHEWz/YAmmxhs1Th0W6s9xMGIfd3p47fr1YcRYXfvKpFQ9
t3uVrnmhyhRzJVyR2HvH3gaA1oNZvopxqkyIha5KUJXgRNvbeqc8h6vkai0UKTaC
3zjlFK6E7Ij2vTq1HY5QEuh11nRmX/FOaw60K+/kC//YKKlSnC6iY9nr3uz3jjsM
+NZyCZujzv21A+5HE2S9MNHJmz9WT9Rjqf8bEOZI3fQwHbCeS4c+Go0F4O2abg1z
QOTrm8HvpkuJr1ySej7byDzwLAZaxtAOTCk/2fSA4Ry5WqiQeQTgM3p7LDV+6n6b
Fkoqbsq9a1GVtHYN58+OPleBzVjB2ZKEttb1fVlDbXy+PtZSR/ucLoxh1QSFnfaZ
MhFfoqdz2+Bk95KTcdM3ukmV9Vrb8A8heuz+v+j1Okfzpv1cmV4WzKyUPFplulSl
0kM4eQRDDZAJNVYy39JH+n/h5kr2lCamIvKdG1VbsxpZvaybt0otizqlhPBH0IKQ
HsXJyLZB/OiSpIo/xMSQZLh3sR0TgmG9ThKNuGxDSaHHGMYjwGjvDKF/e+l/19qh
2m6ZKLyU53AADm7FKhHohCkon9zRLtjHTPKA1tftbLjCqdIJ/RJFNpy9VmmZfFrb
zHpeZekmJvOYjl78sShjDguttKgCl/KsBLXbEDZ9AMrgNPSIYtQi1KkBOdVyh3Jr
ExpWhrEYDQNQZ9gz+PctNbMsTrDJRdhc2dhC92CMeP/0c0W0jI0AwyKf0ldBNrgM
t90R7PO2hV6tz5+bmvULok/OEfncF+cxLAajLXB/17nRPeGTa+VyoweZknb3o6tr
IJ5M2LiLAUFRYi1LE7KRzp0YP4IrI7QfKFwRtfrWU89vy7MQhs98b+ixFd0sl156
UVZYUoAeCm9gMzMcka23E5pZUPH/LCRFAPX7ffHTA07SYYbfLP4O9sE71YXoK0pb
HFjgCybxTIya4ktC0rn6dXsrvxIOBZSXr8gzl1FZXqJ+gUtfjj3DQrcd8B996iH1
B5r9jsoFbpAhMKG0YECZWC32mQUsqlpev2618cReDCZkC+PiJjc0nLeQesH5XA3Y
cBpWH1zIvPNnyrOwwVL8RnVMWYZzhUg9b+1Vum1n8lWDFFoD2J5W/MJZ127ReofF
YNcZuCvFMorN0YByRegV5JAmI5kLQfXJyJUuttk3k6sr9RSK74mtasjUiFqyvrn3
6yuSuBaT9a8swdue56fs570GBx5IE0oucN3Odf1czBzk8cNd6rhmhnkrBeHQ0twt
ROrQ3IYDIFirNHHjYkYsQXGl0mlLOWUXqpMdwd+o3jNMca/fw4/WoWUDFJS/pCaC
yl9O9PwSWQr8OcZ/cIA7znNNXIB4c77G5ptgHsSg5lHt4BS/MdnkSrqLZn2c/uRE
wzofMy3RpbGUDKUNSRF+0FylEXvdoTX9Gj5V/U2IMAVWvwQd0ZEHIkcjiY9k8GRQ
PTUlq6RBp5hmKQufnWJelCI6JjlyDlHFEOgq0ozDuYS8pZ9VaGs3bTFH3f2jzCV7
nPZ5yO2Xw1cp0rJkxOYODrZqSEyaJsBC6Aq7bEA8WvMCEEUWEQFvyJveAh24jUci
9fMOzwToJG9GD+aMFUGNYR2KPQNVSXimsjwGRf0l7bRiSWEo7ATB8cW1necon5Rj
KrnWRuVw9YmfNp35PWbFUFm6liO+xLp7wWUK551mdIgfYngmJvde3UDaNXmp8lFZ
MPOpRl5DH/HQx+YRmcBoqJ5lYC+KjdgOqJXVbk+lBogx93Lg8BykByoCYK3FJ57j
KLcwxBW80x9V2KoU5wiVHjRffJqtc5or1ysMSlityXugVEiyZXZuHRGRBzXvBWLB
b5CV58/5aGQr0IZ05M3TmnW1e7y2X9iqNmmIE47BdzIfiSQmwb2ohl5+fFZ9baO+
Vh+7Av+Fbefy3eGd8TKMwRYHmI7NJAKQ+QhfbRJ5aHFnCXihst7CJXEvnkyLvNYz
JtqYNZJtvLkWfPu+7KCVJ2vtKIku4SAFM47/9cHZAjLCS7U9E9gEfKzgyOXraclc
pAQfnvO+zPI3dvLnggRHKIoEWiYT/vcqbAAEvoYY/S2L+6pqOcc63AIK9EXeHm0n
DhzVaLfrktXsSkL1m4h5MmmNrGp1bfdKOVXwnBtQWT1SH23K2oAGFn7QAfRHQAxB
F82aqzzQqbPq0F7IOa6eS7sNFG3RohzgnXi2SgmaUarXVzKsv8vR+/3tqOYQq5/U
OkK8pwhg50DEAkGimKOIWqUFpFdAtNQKJL4kDilXRbrVduKHjSnuJHYgK3roW2H4
w73NcoDwg/k8JbSL6Zp1JEOSEDcp6QzOmpbOBw90u7HKT+JK8BSTe2q8+GJ7rkUn
B0bX2dISLB4zG+L2acNbcC9+SFtz71RKUHMQi9Zs/76cDg1VN66ulVqRh+JjMZzc
ZnmGEi0vNCjOGOFUBzf85M9lnjr0PIwTikqE+afwn7ab05FHf//7rh7kEz9vCe7C
Ipe3WxJ7WJiJGmjqEQ5PqUXT+xRmoR3YxMmVKhlgt6e8YaA4l+1bAmXi/QPvARpi
DbZnx0RN2NzwdSRnQdG7LqEdrCJ7hkK7bCxYqJfxV6uw0MJ8weVnjYu7wZyBfpYi
wpIbXc2ZlYXEXPl2MHfVO6OZbSZspU7pRR3sA+VzXKKhGhGvmn4wTA5BeO7iwpAf
cKu1blXB3kNS6BDJRcgAMlLnm2MjAW8Focqc8oRNMhOi211zFNbrcTF3QxBDZ3nj
FFGWMqtK6smSJ0wPZAbtS8XsiNbvwPD3ym1osl68yU0Vy1rGlQGZtoqFelaeCJ8a
hnVU+yATNULNHw/yRANFLSNOB1pC+1vEenWKqt5rkxV/Y4qZR3JXATZc3lJOlgbI
XQ7oPMYSbCYfmwEWcm+hRGSg2z10rYtM7DUIAo5hynWYFxS7B9k/mdYJuRzHxMNf
Dh2qMw9rUP5f956R0cnyhjx1Lh3OF/rYf9JvKiCoCgV6o0qOt9kfeJ2DcrlD7vYJ
UXWbtlrsFUIHXmJfD3SajsSLH0O2n67ebgTnZpOhl+gl6Wr03HOqjERFKcvcUscM
5ZEtRMuH2jaAASxLu/TrD/YOsOCJzsev9ZszX48qEvKy6wbejN9A9kBV0ulG19XC
YigOFFJeCXbreIFdFl86TF2Z3HzCCpJCHN4DFrVHd/1zLSuY5O+u9zW3eIX8H5F/
LUiSyWZj5/58IGCr5H/0glaunQeDIM0cXRmmJENv+WBN5j0OMzW1E78hHseKql4y
T76U9WsVFfBiQ8Cf1Ka4PonV9se2/IfOf6AfP2fxhuwFf8KVf9UYVDeu/GuRdYfj
lNRFJFk8CijV2N+VkG1Bc9BfjWpq5QEi2GLptKI/GeMlvfXdK+qKOZ72n7vZSVpU
FNTxiCWR0k7iawOp8SpjmIbCZXJ73vc2bemwxJ9Qi8LlzCmZgtkH5MBYFV4ajo7C
ADzikWRG4C4YUEU9hnESZIeuGnP2C2brbppzXcKFWR2BjIbgn2YR6Y4i08iGN0uK
QY2cagZXyJUMSwLeuD1phPOPhg+bc0XEkGrclwilzt3d2yZOtyDech6xmCs8Xqz+
Eib/JuUIS/dtRD3zjl/nUlGaTCvZIY9mY5uTGljIuY7mbfq89m0R+5PUbysKBS3C
9YgCI4gU3nyQ3EHV7SRpK46DwhOK/1gKFtr/w4donfEfD3SPAfynd5kMirHRNo7E
1eY5dyvufHNQC3lAwqxA2ipXEF/Q2CtGbVIOcZ6K4fKhmaAcgtjDWBtIwWeyAxcb
4dDMThBqD47zE9Xi2lZMmBEJfxaAuNkemOb9ZSfoYG+kLc+MyEHIovyvYWwHsjky
F7sLjHEXUoyl6ocFFe96IsgP/bRziknlN1q6HlxjWgAJdjm+9YZj9zQ6pJllANc8
ficV7ROSGM90QGr2lbw7Mk36XVDRn1liWh2ehhuKVRjZ17h0jL3DpQ86vznJnStf
yegRQAcnLkS+rxDTCJxAs9wrCav6o2EDpYG6yrOd8EGcc2qRCIqIP14bioqBFzQU
zN1Trzpx1lOAX/euulyFwIWbfIZCYC0AOjp8t/NQqEGtDu097HBoCSU3l6uDiSXK
jR+oDwamX0Spv8vMzveh6bCB6wvcSj/xJpGBQNewbmINM7X7g+jxrUnfWZBLzpQn
6Wpah9nqjSie9lwtnahtYi/F8v8rh86hroz54Bp2ErKPG/YLKoVAJpSlvJ26pcni
0SZz17iGABvkhWJA49kfrieMZZdT7Wg2DKrPzDrStzp+x2JlvC6qFFm+g2YWxfRk
sEn23msa5/Dk7+9YCUvwQMpC5jMCYRDRMfoU1sXDdnPmX2p36qouPVv9IHFKydH9
IXAVyEOLnY3psO7cdva9nR4ZtLbXSXFpJ8zrhT0Q/i/nSyMO6xkWWkn5uK4FU4OG
gKActeADr37jyj0fpLNfQPoJkTqX87vkMNj07MSVYO97SB/8SqcxFhvyp/k9XfbG
g8KjmLtpoQzPVqdIrOqWd0gH8U71ohajpnrYDN11sz0EkwWQhDWUP/Uy01Ocoaqb
2Me8r2r8DwTcwtQmoAgGXWsomfpSMwbYvAa++QrPVMXtIyFTApxXjRozE6aWc6ac
WAqKJee/L3C7vB9TwZg3tXK0BVKpHHKsON0kBgs/KjY3Z+GVYecRib0cl5CBCQI6
28RaQQMHY+J45ryXPTKK9tteP18zKAVrEJGbY3fVgAm3S5Y/RZrluDtcotUCuS6/
Mou8uzoZMimriErJKxLkf4zxewsIzhMczwG7tFD3jI18Kc7szVsEUroy+5i03QqJ
V6a8mkRVgHy52PgFqQNufYdRn7AmiO6OxMwf8Hjnnz58BW93V5Em7USw8x44Okmj
omA26/smkG352HZWSTn5MfeGrYmSdNXzS+0d5tg2YkfqqFaXpDgVdXcm3x91z2bb
RUfRgr8XiSMIFSBvYNYO7whkUt85QA0/YQ+7WRTW1BW9PbyUnaT/63pPQ2PwMjuX
x9U+WrwFIJWmq46aF5MGaTkClBVc68kcSbCxQzkgsl8dyIsmeY/+FPWX0gzbiZWv
33A8zbpnkQO2CmtzyA94TQ4QZbiFqMGMFWp/Rk/m5xQsO+arXf/nYWjdeDTYBpIC
sy+MQU7Z3h8y0T2v/sGRtUJmwsNVDzvvDi+Uvppbabejm0yfJPg3Ke0lzF2HNaCt
SbsjJ3Q0wvLCiYzcVSNuAagaWc4VhM827UZgypKUkofFcOqr/o+IfZSbPGxyhSH4
ypg3vPpolTJkCW0JJApLVBkiH9wNB7qmm7TiV4xsAkiRDN/fJvFpApvNnO6PKxkf
XLgRaftIvJ/hcx8pOGY3coZZW4RRH5QfF++94UUrIxmAU2RB+J2ll9CPoeIR3ofp
wLKYaDJ8u+70xL8tzIGwcSgwkgK1vf0z8ll8J0+fdJ/1XAFmuk8aufEz2NnN/DSV
VA5kdbJWxmx+u+HqwdW6LoB30jxse5Xj1d0PLaSn3gWjUX2mh1qlaRP6LRFF5KMh
q+z8jGRhB89K3YREO7hMiPQ+RCEXie9qSgQQdQMc5DbhIk1ur7Ln7CovO+TH9s9n
V8jkINO9a9Tm3JExHGsDNucoyRpJSJpNcJxry+8q5Y+gv8GtSXW/Flbe78qwaDxL
fq4F7e8ETJpLtsKfoy8qkq6T4B9kTYaG/v9550sDu+Gy/8z+ywOZo0Zp/5t+KJpX
QfO4B2d06PS6Lll5R5ezcX9Q6fb9zSGqIy8u/znM9HvnACC7+4S+slwSe/1Syqy8
dzzVmepB7NVMS1eeLtVxeRiYnE1Y30iNKXgb3gcvum/4+pQaLoOr3P36p8cY/TpU
iRaalIHaAZ8VCCZjVApdKky4ZCarAbXBloGglhWy0YYuw3jDMnpCHQiebWp/YgUD
NECdvoG4kUgpE4gY2Ri9klXHLy5lO3Ll7HfUu5bM0gKaB24awSYEJwOSoHCG5MAg
gaEHX04jzF3fYh7LTstcHMVI9nBlJ3MuSAMuLJlfgDyOb1NEX3twR9aF3FAhxjl3
iiF9XhyCjODQeMPGsZFQWzSmS5azy9XFjq6fZEPjo6NHKRVKrcCJcrxHTsDMNgHs
68a9Iu1KxsDZnsyp1HKNCU/9oy2uAaGaWxskteEZVJrBRlA2natlCaho53xXPCTU
EhXNC+kwOag7awIYiJXUDD1jqPhHE5c1YZxE7A7+HDW5AkuCxd9PgwrgGg9ZQdbE
J9TbgMP1ldambfIPxnlu41ejEFfWWmeisbYT6FCoFFbu54Hdv8Chz3LsV3ybrn3i
zNhO3QHfzpX+sLw/vryliYtOobBn4CJZDLA6GkHQ7mZLS+1uMETQvyaiRSx0BHvP
vBL2XZqLvFWhDe3xfknPH1qPuow+PFZCww2/jeQJlksDTbDI7Qf5JTOaFHidu66q
oMMg3a7dTyC7bo31pDR/qJm829GCPGipGwVfjttqzjkPgDKqv5/oG0RMGRVKKtJh
dFDoy3kxAIPnzOuS9jiYeN5Ciog0pmFPKuCTh1gxNU0tgiV06CSU7i0d4nv5Fyo7
Qu7zOKzZUt716b1nlwyd5HK5RDe3A6Rt0FMQeoqo1TAQQaMABJ1JF9MsSsOaZH4I
OvEh9x0a0+Gn1TxE6UEfoScqcy5TLy2Dg5NZZHFk1kZ/6eeZooOVnfvQy7J0CwZs
wL5ptvx0YddB53izqvHJ2Zh8R+VBeEFjBGJQCrO4n7pTmCo3V9dMYsTU4BusWRdX
Ml+tghoJJ6dKcS8dda9H3f0jCofauuEbXvlwRXT+K2SqjHtg7gwzZDGjXTEEk8FG
h5GSjBBZLWcDtBOXKUEBcZh2zmUvAulK2Kul4pUHNIlXtOmwti8AdmFiYctpvVyM
3Qq+yXY6CM+/LEGYJCnrtJZowcLo/YMObyO5ksE4trX3lEL3RUjBMKOaZPKP4uIq
7yrVnmmDIh4EqmAjRZug/F1Xgz/6jX6zmPPCbQ4BR9c5cVcf698QDTouBl1SyZP7
2buLt50tjrI3Pfq55U2MVQSuHO7A1rlNl2tiF5VFgVSQ+583DtkuZJEAfUL7xdWK
w1N4HoWjJ2FWKlEtTS8yCrnznWWtjGKhXutd+Knp30LplNljAggODhv7pNfyLL24
ZdDqlxi2qlZhwRktlLkIPPSWZ4fy5VF9C/LVWUxghbyCaKOJgpHuM+9r+BgwSrD6
VRlHToWSpeGrcEvApPvDCWdVFJR/71RfUmqHVWdzjbqrCJtlOxOh3DmP69OQxNJE
lvtas9AsGb167mYIcl3bTG7PXjlZy58rupanQ6T3nFe3S/T64zseC94Mru92LCfs
svstyUM5BAi5M0iV6HZPXekhg9pJg7rH5dthXhsu14rN5T111Ra+A8lSbElv7F4w
wJuMCDHQbgCKV1o+yHMo4102Rcc6rniVM4xU6gckWAr0wqoE/gKd0Q/9mUYRSP0g
Rnb4wE7ugjTsrLwd3SkIkJDNifQrAKciL2R2013ODFs1IXSFGOj7VyNx9lsXTqOR
Jk2NgHDaFwDLRKaMosbt4nv1lstRxG49GvyPHC98JFQdJ7aXF/DjyMAd+xJS7Tpf
GHMlmoT+cIviWOSQhK4Ln8pUNnrD5AopchxBXTehlLRquyveLli04Yz1ETpaRm0i
eEvh6rKrO6QaTPLuZ7DQ7eEOveWjLdJeF/qDF4W2bWSW7c+6cBQUJPzQzMxuZmOU
AMMCX04xmh4Pzf1bdnAvMtv7uAfiMY0mSkqmRA7wKqc7a2K27A9RcfNiT++3sHcz
StdTkO9dVVLRrHDU1vGxYuYCTPN44RAEM1bRF0DlQhVE3SsfbMTlxE5wSLi82J0C
UcMkTRJhgYldJDh0gq1xYk0M3uigEMIJhOWDJiU7iqW2W/HTzfmZYkBSP2o66tcG
A2mcEXitzFuHKwb7fqEqn7Bp4akqqFSaP4DJ0Rej4zV6hkjuHODlYoL3qau3MElM
ga75ixrrzyFLDazgXYYysNWF3JdGnkrxB0JE1sSbut7vxopaV25oiYJ20J4VdBIy
quraCu2GAIahJRExdjuIbaXHeiqEPwTMud4zIWoezBfZyfWkyH3jT5wd6m2Deuc0
OTXoz/tmCSFelOslfgG1/MnqisdJZ7LL3MCCGHirfRZAURvmfssKFA6c1C1gzFAD
oIY5PT+gsuRcHJb3wMWh02DJwmVVZpyrZ5Tg5u0tiimfBYdQ4m4oB6B2mLQfFKSQ
ONq3WJ5oAcOE70hMXyutYFITc8nziPqrZXgKG4AQbL1NQWSr2Ze/QJ83aqHt9N+Y
A8Vv4EI8+PNKI2gReKK6xqsBd4SWsWbi+NniXaB+qjsVzEjksqN486dmScGFNDJp
zeRsC0vVwa1N2DMlhDh45R7haG01DLC85wElq6qtXh/fe+oH/by/ahKKmpQ3xt5x
J8zP10Z46JexhEIhmgI8Dtzu9OZZENwOmKMrM5yPHzpsneU3/8uf1etf4tzI+jrG
fgBFXsQcuEr/OLv1neRoMlp7TkE/WmJ3lRIMPzM9J9ZwTR2IT9cnhtzUzmoQIkHI
fcRobNtl5ye1z6PNTeKof+lxMiFkw9Hy6fS7GRrb06QjbID7Z5l9FvjvX/XrpxgR
GO5H0OTIxW6ew/fBKr6q8ggZjXArx53EhFGBeWdhOvFh82F53P71J/jk/Wki8yx4
eBmSDHfayVSFzGtoEDBTEBYWOLnzbBTiWy29JzvCuNnhxeRMHXj0nfr5UXYM/Ofl
875kLSgH+HlFBezQFLbzAar8Ab2RTvO1E4wGvvkdRuJeRStuiuwzki0NTY+aWqzL
/DrifZ+zzLZNgpKNFQ/Wnsbu77ZebrzCCyqCGnCOqqL9CjlAPdJ7SvrRVTgpeT9s
qG/2Ta/Kz8xNyDl+3n/DwrJVFVjoliKaJ03iTPJLMDY5+lGSlCSALhIYh12/aEVx
kqJf0gBwefGnyfAFVcLjOmnJPg1IDyxSLauJ0aoWc0sWXoEflslQr6C2Q7rMz/zf
yxvOHuxA01Sf/7f7WxArhDYWFDzPxgMSR17EjVwdLZV5DlYfcU0V1yp+KjPt57M5
egvMyJopjWuv4S2GLJ7zv+U0n0b4iW86OxdxeXjh6SStWuXTxg2dpaTfHHZLgCEK
SBIrEjSbgYpUEGlOERMi86X7WTPIQv3JcfG6u+ziA6s2r8gJI37qUrUYr/2kzsxo
yQGjeFcPSxg2Hi5hhaY2o5pW62VE8UyLxyn/dP+GHmhNzEZ+4kjVwIgo+SrvGCkz
u4AYQsyulnuMrATqW5FN0It9FjHlZtAVpsG1GB+wSzg+beU02X3X6ilw2K6r95yZ
WdXxeTh+c6AnCV+TJ0jIgIGMR/Pffmeu44NP4LjgTyC2gIFSSyVIegk/PAf5ym6T
FV1sslH0gxuxfFkc1t58gnV+hJpr4n+eIwkwwyNxvIjeShsrnl0EFwQ7EfvgkKl1
pBAbfTwUUzq8zKR5xKgK0pWyC+L+cHeaNw3gc3yH6bySAXErs9pXvXxY6tDLrAAu
hiMIeb8QeYNxCueOjQ2bhYsCy0XuktYEgmvzbXAZ5YMS6rQ5lnSiSDn1YezREvc2
yeAnCK+y1zDC1TG9vVpUlMZFoutZT/u7AA6t6MJQ0MYMx9jEsFUBnKApU/BCLFKh
X1j2myGWRgq9IbCaPTnlGBwHIIQtXxYfXnDkAMYvlk1+Hv/SoLfDWLJRrDAP1tJD
f2CPW7Gh5AgIVxII8ykFdwpGuvsPVaAn3kirqURW7Yf3OvLxmwPIEwoSnLqrDLJY
detqtorRrdg/tQJY73HBD1wGJykxV6vo+rqOGbE+vdcYEk8v3hdzcDykKUWKgih4
AmMnVhNglVhbjDpufsVpZb95ucl0ZXxUi2IREzP9lRPZkKKiEfKMFuzsUTheuqL5
G71n5rpEZCD9QSAlj8pG0YC5wgRZa3o+3AtK4uIWM1rhMArUe/sAEfFXwBbbvjrQ
eCnOh1TJcCBkGVXR7dy6ac+GDWI0fBuY6E6BxLiTS+T0MhDFGp89IitS3jjTPI4h
rpBVZvo2bw68Sa3IE/0BfvaWcaNWQl5B6uWtQ0S98v9oGs0O+rP3N2HiptRWjNp4
qk1BnWY4t1U+6dQc20dHudaC3urO/bpfzyzAD5aiyhwIhvpQf4y8SWNP8NGyhSWu
Z1ZiNrivfgOt2zpTlkuXl+/e3A0kx1osZH1+BbVfUcMCDtgbat/CCE4iQer+BZZ/
wheSmPQ0/tGsw3XP8/c1MMKRgavSh1/jkKx43G6fyk89RyZZkW1VnOTPuTnnc98V
xtszqNgwtbqaY0zFDzm38y37lnlEYXk1ygOorU+xH3aq421Y9RuUw0zqBfnOnu3T
6FDEW/hyfojhrWET48NhBwtfipS4SPRdxBvWfoXSOghgnj2KIFGkKMcOpn0Gml0+
PZyel0X+PboLbmh5+e8Vi+Aa5oGspHhjjp9zya+oIPGzbpFIbViU94nmR0BXlqLg
HdUqexR+i9D2zplEi0Opuk6fc3EA6n4+YRgnBeGjkQIcnED3VJtxfYQgMWMmbiAD
CWamMFW/RTQUq4A+d3iI23TJzycHOqB3JlPQJWCcyp1J4wWWTY7Ip+kcIIhbVDTJ
+vaplRTcHb9FaOVtfcYSA70JfTVcKSg3odw1td/PPJZ9av9ozSu0uS7zLuHm24PP
fT6Ob/lRmATMuWyTGia8XqwC61yooxaHn3E7Be4R/S71R+SmkPoak6UhUoeixEUj
NaY/f+9ddRkJlGiSjM16eo6n6MzyNpZ/tvjaN2Ca3ywlH2oDfG7rCYQRrlUMWfdp
xG/00T+tZUawOos4iW7TeR1VwAB/amm/NgnYsK+BFWZfS0Pgjl0YViItNG/c0DID
ZC3hg221op3y/e5dM5cTBFvQBnBKZN2OKhQCpisDV/QUG1Z+MqB203085UPH91gD
BzRAc+282h3M8xBmiZM59kt4f/NtAxiQneRux4sI/rQnsYcskFMVQoKLr581ZYqo
+jFKUhm4HqGt2mvRiaA0DPO3BQZzpLG6G9/rDdC/3+j6VkrUDjoIr1e5wQcTZA/4
YnL4NgMhqiQG3/J6DOercKvPINymf5Zl+g82g6sbs5pNc3mQVF+7Csq8Y/ovpIUE
yRfnY3+nDQNBKrv7M60IEoijkXSL/6+3ZmJ3X0tE3VWU0ZqFW60OuxaGGTC2QTV5
A/1gd0hp1RXE3uxrA/QzDDzF/Xn+ad/Mr16fLyoAKagimHWSr5mNHVJBar6nvafb
9no87uPT1gBH4g5s9Yhst/3aqOq/pEdentk7TZ/JmYrEjkrCqIAhM7iaQ2AOJm2W
71MBUvy3R5j8thhc+qtsu6Www2EGnAq0poM5iiHejLXiio+4vpR1fEd6liZJhCbG
LKjM+qROKuSZXur2LGTelcBfa4ippX3rrBikJr54PknlfjkW/6n/3GJfcDG/vXyX
Bt2vlVYkSH6MWUg9X4TkFrlISLVICyj/sRwzAcyEn6+Xj/duE+F0dKAGJoqWOsmg
`pragma protect end_protected
