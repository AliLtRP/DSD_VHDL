// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n71RdthUxxttTdoyAvWBhNW2oswpHYINKmnsBP6xioXI3B1WrCNkH0azHO818ohf
Lx3E/kAiz6BBGMlfV546FLnsnCfapXbHezWIhK1WbdV7dyPtJIS/YoE/Dr6VBY31
w+t0juLsvYBOjqt28EmlkFa2cp6lazdkbPq00yRu4Mg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16800)
J+3G9pUrJCo/cgkJYs4T2pNYBocDbn5Dn68QsUfDwhkvp8lO5GwCnlHrR5ZT4kRF
2beonpAYczKMHap8Xj94WvHQB+6CZ8ziPgihBNo0J9pNbV9N9pUSXRr4vrpeudoY
J5pg7lrsxQeWlGZwsg4hQK1pRhamcRsGXqygtcXRj/t9QpaKyzuGTZI2ueef2AWD
fUurNda1D58Yqqc0NPsNN4e8VKieTjYCj0XQ4AX797LPBG8UVqLehLCUMF7C+CuV
yEw9z8xvSjK4Y1wGGPjFTFlci2TK+JuV9VHWqDv+4dbki1w0wBS1D2npAXeAzz66
cUQ4fq4TEO5ifxavkb0KhwTDm+Zp72Iho1mqFrd79Hw3JM8o49LoaGZksJ2UNGaw
8ruh4facLJZHV7iBv+mN8Hem+mITQGV1knrIwayZwwqws3poyEH+vOncq+K6cfOT
nvtgg38nAb4j8IhShntNpswhgVrB4Ri3fuPti9O78P8m7V6IK2/Uc9E44MF5pVxr
cTf62guChcccEcwGrbAyjvCqB1wZ6+8N78XTIKsHBoVRYwGrChVSzB0ZOUvQoUVG
8LyQB3B5yHPGPzSzUcd30ERPodmCjurOgmzdkyGH+8FqfNJYXaGdG8fgMFhCoMe2
CKH1G99weG2KmhMcPua8tLr7MKancQmIP1SRhTl/VGffAEoqZb0/jKOmxF2D5lQc
YDCPWWAoILucoUfwOnsd5b2ZqUrzaRZO2LGqWA8mfbFw7gfihySFFXXFmyrmhSLV
8C6pqVuNhLyU+dP7alhRPEBa7SeXZ6PYLnzgEq8xGpAhQRgD9xHpTbPDQld3tCRh
8XcWWg1c4deitLM+vHKppmoPuyv5mCc/gTS3hup9McyYhAisXIIQgMnDLVbiGA07
GZSMCWcITbXwCfQtCda6hhEK9Oyk2HlZh4skbpE3t5Y6N5Q9SrZn7kWtLK3ZrK02
dCjp2nmuHq8WwSr/jz4DHIZrwLmhHgq4Gvg1MVdHB+KO5R/cwGvk5Tju3gXopNw+
cIh4CM66zsdSzM3M5VD4HeE5ENVSi1gi1TWYVEJWIb3tvmxOiwz3o5g6b/FB0bH0
cfynSLho2LreGzNYNp4B4ch1fNGgbB4pZVb20RoF0VdHHLhD8N0dcBY2VmqZJ9nT
IOL97jSxPWJiypEs6/SbCVXltKp+trQNj/I7GK9mgYP71GB6umYtgFuspULgip/z
W813gXtoJUNUDeeIUWpWaB0UPYF/ieESeXhEeMYutEz3aQPROeYUvEoTMs+B3cql
rzsAQq8njZmRakihT6QmTX0UkaT6cNqQv/YGHsBTrMiQv1UxkVjRpwhCFSlR5SoP
HBDVSkvdrCHYWOYxK8b6E1iKoviZBDMGHdcjDSIlYzTLr0Oy5FYAHW92WfOWQAD0
uIJtNmvH1gMBcg1jdHxHAJuxyeRLeXjj7STA1Uu0T3aan9+cVYQyWlLIK6BqtjeL
kOfTU/A0fGVMEgDaQhg9lEyh+REnOeOxxZUPdJn6dWQUQ9ympvkFaWNIULIw+vSZ
VeM8AdVsG/vuXNbOE4JbsEl2jS/tko6w8jCCg8oyRhcv0vKv9sc1tFOta8z26GfK
h5UVsv3EiCtjGlkLx/rFecjfa1IEKLHBKFO1ato8voKgMhcLeVXJO4aNML2IRzKb
GesYXtw4s2LjRZ6V6g32XoRZy4xFU9cimBt6jPYOugTwdCQLZ14y8S9uxyhtpwn5
VnJfh4Aec4/H5DehSqdDDiyCuAGXbZO6OrhmCQRmA7T5l6bBQPVN//eM8H12zwow
JOYf1AzJ0+UbU9NJOeU9d4xZL6N/nWa2LFiRWcRvoUyLcwEw1G2cg3Cz5r9zhLmP
+mU8nJIz54+L751s961CjFq2n1MkXDzBSOVt10cAGKwPozoA9RAQVOgTaf+3zjyP
ziztJwqajC7fXUfMJ5unLYSPSOaOjThdC/Or39Yw0JY86D+f9vNRJjVe2PGZkUw5
sOKsMlg2evjpzU2j2KVg9WhVC53y0B5voUatnzXFLBXlCKw+bPMTiC1zuM+nUs4b
F7ZVx+eHhfdQt5/5SWm6BPJhDIzN6RREwULH1Uvul2zqYeK8HC0qtpMvQpESKFmt
bjG/c/KZS4uT0Ub4ZKJIiSeBaY6Onm23hBN5ktejm/fwIPbT57mjAd+1G8x8gTJh
HoFh1Ce6MjTGyaLlwycj8M+npdHsKqPge3hbz2roGXoJlLXAf47EoS7Z9fhHfGRV
fKG3jBkhRnUDMbu3uZQv9OgxiWpw8IfJ0e+nJConBS8xFJQsXskniQX0scpmo9IN
U6mfjk7MpSaL9JDxUZ6gpxyrPWgaZpernv9JwZSa6Zq+Ogl8zLhyL+rXY6jxLLxz
5X/9XHTx5FqvMZazml81/is434nlF8tryR7lC9HbUSzYj8v5N6EkAkdtKPbOhU4O
5hNbUVsV4eGg3mRAFMpUEqeT6CXO44pSIpJrn+boO3MW8zNIupJPQA8QvtQBroWG
wZd2ZuGJch/hI+HwzVyvErzMv8dEdY1HtLUZKYmVmRHfMlHa/Ka2vvNdj53+uxa1
f+YI+XqRghGkYimDf/bZH0ZW36Js3eYBFuC+b5QKjJY1f6xVcKKf5uy2VSSUXUMn
MXl0gQ0zJmHNN8Tu94sgesPqU/KAUqGyF3YJb8r/dHH+07MTSDGp+z8Zj5suLql0
Dp0Vqm7xVz8JagN9qgygir6idtfUB7fH5fX+WoYaTPbSInY9emp5DS9ViiJi9F8i
TF2/i8S4k1refTFVjNz4BzbmhH0ysh+I0m6U/cKf/24w9Dq3/+fxqECOLGjso6no
O3f8xUIEDgd7kpBTri32ofjsPakHQG+QY9Xv5L4xrB1ZN7jIB3v3qSolHDd28c4l
edgF4O+lfaTaHQghsrIlBiJKZe4V9Py6Oy9wH56vJrkDDYkomou5oXJ4y2S0Eoj2
2sKT7yGm9rKrKSr3yUy3uGB8YENoRjDwyTouCotW/EF0fh+0P39F8Kh/XiKqYUua
cAZ0X/IuF5CJbisb3L2d2QwrEl5tOiL+H8//+9ZKSw/xtXppMIqumkYa7V6RPFmk
nP7sD9vPZTUAxHqE9wVo/UoFznOWXsKoJicp3jrx+76tWp0Wgy+83s9FJQCrRtoK
cx3T3W5+zYoLAgg51p6nHuEz5Oa4QlnZeaad+vigaLE7wVHQH/jB2GwL7o7BJByH
WRY6jeZ5JYGa6Q7vcLaGe7mloXnm4QkdJ+l4fJhlZBrFkO0sVjtGlzIUXkuWG3yw
4B73mATzJQyE2BSdVXVliHia6NCwbvK/R2t6RPWCuxX5COyQV1lukS9uNS1Abjid
BqGXC7hHyv1kxvJgsqBCBxuJ3Kgw+uHJuQNPxG28YygVi7m79lxr2AST2bNKCQKw
4jrf1JOnGjcoZCOyJTd/JTgfpkAaRmmKbLz1pqdNYMnB/1e9yhjDlqoHOChMKp2x
KqqTDqSc0ClUSgywuAHDXIZMGVk4UFIgGqqWMeMtCS9izyM11muqpyJzzKUj/4i3
X0/zxtX/WgpfRIHIRvh5pgxwwFvQFID1ign+lhKrfIqlaEZmAXttvdibvFwvzdFY
jHzuOy8wG/WUv+AmMCdMCN5VxYmEQqaG6WyQyhu1e2HUgpsY0b9c/6I0owauW1S/
8d4MCUlEfS/o2+ciCvUZ+HXAX/y8wCq6T3oJFGN50z/sGWuFKzqwjfPPxXVSiT1l
BvxjwPnpNPb0mtEUtJufKdHl9s95CGnJvuKkMe7cLPTBav3/b9lH3JA3HzP1jLr1
ScyXlrgwof5opUnbTiY1yHHXs802qBUyc6Y1jaYgrboZVxKbaGZ+v2ITYbnPeMgd
V12m2l0MCVN/T/MI2+jcLxnQV+PZweF5GlfNQweZiUCnCJfKfh8xkLNIiLS0YfYe
dvdKIiB+g8fF2S3kN2pSIX/kAXZkWioGEba8XQVepEOu+m3JhD7iKaheEnqUyxbJ
q2aEpMOs85RwfANeLDVWK9EyH/mWXY5r4JWINVKvs1dYwDnq8WvWoI3m7BdXuTJl
r6IbtZxGJ+6KobnnLcdLAfmkvGRYK/mNmP/G4rl2QI9KBkJl3KSxVLuESnM8QyvU
M4LThmNZUepBJ+ZzT/vQYLoU6B7f25+zjRUFnU3jA1qVte1y0ajf4sCMVavTWKeZ
3w+wrf+mbm3c4h9qUtY1RL1Cq6ATRYhU2sRFiMOyWzzqPWMo7y4xnh8/BQ+Rxevj
daa9wRKfubPthOESNUQMXcbfpcyaEs12HTJFIz7R0Eg9z/4d99BMfb91JYKT84Zy
zaRnJnWQWZg0tqUxlGNHnaC8dV81WdyJMjsjgCM2MhTHOwPhnLjT1wwcHQyYS05A
PTnXCswToLfmeh+GxQDjSmEM9bU8wzR0siDzlnsq49HoX6pcwgnXYfOlyK6FvRxI
/AoB4JxRVpeOAtzSqD/LMET2MolARd2gsZlygsqhfjp7gFEoe+nUkKkp+URDxGIx
zg8ZguWnrVE5/Wj9j3Qd+WCf0BveC4wwEqDZy/ChO72sy5alGmXn7p5vBQzVyDFD
sWMuCkKBZx/IU7ybrMi/Vsb72IWkP4i5ewvZkiydmZVz+YrIUKWtpSVppudxbDLL
Da0ZRzsJcMOAqrmAiFsopF7B6peBgwBR2qexs9LWOP3ZCx9W9MNrBjK1nwoA/Gwo
RUZdyYEnmnvDLeC8+VVf54fYTwrNE9u2UFLvU2L5aSoT8V+jo0Yk3PBs2ECL97Id
g5OUL1VAFLXxsdgxqTuTG3LKZscL3EvO9rbmxWDz/DK9Ta8/VF80g04RfQN3H5qX
X7Xbr7q+QQETwqyREZ9n56h9R8wEpLvDH9crMMFqmJIqjA+JHL4mL9JhSnGWaIZA
bOZqZnMssvfoBfz06LxB0tx8Spa+zmqBzHruQh4iKdM31Eygd4H0oQIkFYx7t0S9
z/lpMrLT9FXZTwEU9cnKniAIeIbvSgfJ2W8NI+WP4aECitYHy3V40sA9+S1vQYyu
wPRuq/zMC7/8aMGDvSSxmAI0YCa23w36zTp5PXOPzJZl0SZNzSkqkECApGwezs3K
1c6hhSEnz21hQN9OU5oCo4ck4llQevSadGtTuPxBoV/svlBBHPtrOkcSMExIUbov
RcU6KLmVR2IAzmlYOVb70qyVONNZWlXSZgStaOgMCRmy0jzZ3nZdb5yke66YljEs
FCdhjeibnv+W4IdZnFcmz35UOufw4Hb0RHd+OHmH30Blrum2+J/6q35j0r3jgjjG
qoz8yoO5HI+XI5jwfdoZN7vnxU8b52/c5yFuod5dUNPjtSMjX2uvYVdbGJh9kPXB
toOCTptBJj8pgJAnBnpmbiaCf8fAW3Jdfm85H6FEJAZAa+UaC9HFo+LWncp7DusF
nwJhygRMLBELDiiwEKqBITp8Ce6J4pxoT0UCF3kdWb/bj5VYfzSpZ2qktN+6mjpP
c4lE8IGj4KdqOMPhZCyITEsN/Z8Pu8meki2VDPe408kfNsXOrVtpPiBPQAulmga8
3BQns/5vApy6O1H6GbZicJbv/8JdYH+k8PmJ1rPtixZr2LdF272Vib1OqXzEXISW
PcEEsC6RsOrQd7qj1QL1Wcb6/nie2G4MSeFXddLgRzxqd9jvLtFXi+zGlNTlmvcN
iOKxqyMAt9noiDZgtM/ZrwUenQbc+4ftAx2TnuWDo5qzN6j5Xb/MrTAtvFxmHLyz
fDrsgJaw3nh2inKmms2mBCco4pWBhCxEjF1M4Yoyvby2KOexw9hR0j7Q15uYIaSA
DeeVwTPZTpQXcVdlK4np53+BNfy+oYzd2CbjPX0TRfbUWceHjyDvqhofWtoCBq6e
uaJm9EFq/tnRxmDAQzY0qf8rm9x9tWbN+cobAa629mu3eFGTbG57s3uh33r4TIYs
mFdNe43ZrWSSpcDnsROVQTOg9GabUjkggdEutJUfvInKJ3Er8vz+H65Jbw873ewX
4SGDmBd3pKIw2wItbz43IeYTuTRRXrLQz0JJLMlV8ryvO0T3yfRxN6Qt/BhMyVcv
OUAQq3tHJUxkBFzltcfKVSN2ziUsWjjjnII0qV1OlvRBnhzhhIyT46EoLmiashfk
S4P96Rpf2TUAmCgSMhCkKr3r5XuSURSG1U/eQBj8TYyjtusmaVIC9D3dVrnM0hIL
G2IsxOzmdXkbJevqlrnmkuipiaMbKHtfr8Kyx9S6sM1VZGqn5pbHLQepQrExCRPQ
9ahiAChMKLgJr3GYW33erBq2MuSwvummlt+ibSaN+XrZnnmosjNkr5wb+dzcNrXG
+CCrg2DsQgZl6PuFjQ1RBqP/29/BIZakH6KItfD6sKRp3k10ankHl6lpkeL771TA
CGeON/QoJk/B8Y4t0t1VL9qH4B4jO6hHh6c3wUBDZ64PK6dY04ik4yNENOacviTz
4ckumaz5mkE+lg2z8QwxNyK7elTxD/aF9Wy65ScxhG1SqFS66K8xRBCNWXrvxzQq
ViSlMsTei64t8QJy06zWb9hgKtWBKuKnwaEozJCelFpd+JN6QeuzLkqW+27riqPs
dbIbDJj6Tg5XFtCIUEXOP1KAcpDC3EesewLpQbT2WkFlhkbWbrD7dRShyMzdGmEm
HdNYQbKHopOmhsAi23wy3qCUSOsH5kA5si7UQkKOSm+lHISM9y4lcbq1y2imyLAo
+gaEsvzmhyCJfE3ThK0/4oaqWd13jUD8mhqLpVVY3kn3xvu5fE02EXe0QqN25iAi
fPhK4rAI+2B3CUsM2p7msbcb6WLsJ4cD3nIVVlF9P8ywwVwzwKqE8V4MnPtm+Fxn
65g13DNfJAzO+PtYLfpZcaTDzo3iZKvN0mmQY4AlxldX03hrv1QceobBB6lteggw
jTIgX01QERz313MGSebEe17xM4JF6x/9CBXdQRnPSoU6iq3K/h1uVZZ4nHX2V+28
aaIIWuqkEZh/Qbd3QbXJtnlHcP94iZsgVlAi91eMYcKKF6gS8GO1eH5rVrpm0HmC
jUYE2YiwzxC72ZQRFhrbaaKqnNl6hOTMto5uFkOLwEVlJdUWK4T14kquoIRDt11T
dqB2JG1XKyolGsaHpDDVFt5oQZ9HskYb/dA73kp4JTJja3eNoGgFlRIda94VAkBG
wYDRUzxPj4rrxDl86ojJ1OdLOb90IHC/5ES/gwF54ypV7ZQu6IGukzbBz6d6iPbx
t51AcAgHYTMmCiXuM1aRYjnIftfkcgXQBYrSv0Ko74HWBBvjoghpnb3eId8hGnXE
jnJtOGUm8K+I0nr73sB8TTkUWfvn3y10MLM5wuHENhDBkC1l4xcGS96b+no9+MpJ
vYwnlhipik/1f8TRz4s8IUJcaZFuqYnGnLHnjOQgn9U4ryTrsuVNwI3/b4UY2EdW
HUzisIswoHx42KmoK+N2NmsRT29NwfiUn6aoJAANaWLvLzwZz7KpuG9jtj1urM+A
D9kAmMJ+2nN8QGLr9B63L+SR2iGUMSPMwW92dnC8jSCI5tgrjqORxg3YI79Br9rL
8IN/BtDvizgBetUZnR/A1bUVm2zUM3uila0dpNZuuF5lfPcjLfEUn9QfRlhljinK
wuUFcye56lfyT9o+Jq2+Y6Upaf+vzoAjrzXy8rcc9H9V3yFIsP+wnn+taiK2K9BW
EjiI8Bd7ME/Z9NKu1MyVxJQoo6sxIAsAGUlo9XKrGBapx71wmQ58glQxTpQ9jTgD
EpSJkvd0fS+hv5XzRi/m3qdELcZT/S5KeFuesn0T68HP1bLQFwyJZ0E8FysNg3rp
mbXDVmcEwAqw+fIJlvixZdRg6LHT2xI6d3PQAfvZc6Hd5EyW/WCEOT1L9NXEQJhf
1svLc2IfgKsIMR/mBi0f+Zq4HHaCXrWrfjuesU/3sPGm47XAFY3TpXNaRoyT73DO
ilSjRgApmE8Iri6kq4JKQ4YxtknPnO7ymSxEtdvvRzInQP1eWKu1/iKozMgldyao
O/65IGb0ofOON/PvVGIYJcXPXgCf/puouc/A9iLH9CwuHfphlC6JQivHxMOAjZex
iVH/wr4FwPT1e2o4GOXOdTj9lu9lHlUuHypoHaKHrQAVXUAHWKQp3kbaYyml86Pp
v6QweSPSCMoBd8DZJEHU6o7Vi+xqvgDHdQ+I0jp3oEizq0l98NGPbtv97qykvlet
Hl/koaB4D0uk3mSaAeDgP7K8rAi6woy7WSQySHAkdZuzrSfILE/GN2JM53fyyR4e
IL+gkQa5usprYd9Dtp9ShfcoZegDlRPsG9XiCt2qG4y0c8R3fQXKvSaao14i/BmU
KT/lgeDMl2WYim+1/4p/WxCUXVKjVqiBJXYsbdr91+jlqb44dXToy+oxFVSTW3H2
iK3vI9P+UDFZWklh7YZrXfuHBax1BEgq6FzF9XZ9Ay086E0wH5xvu3tsIUAANGE/
8J2qAl68vDN1qd8Jdmnzy6MR584qQidGaacuZBpJsfUCUH9V9d56e7762+lHJwlP
ub+A0k4y/jBoKfwTc1DNek+OWHO+i4PvS6zMtjFc5lWVZvhQQqEsYzPRrYetQl1Z
taVvWVkSVykd6QCaXHLHlnO6xp9XPmEzy6UTzCw47Oh+sThIwGA852HBgJ9v3QWA
sdDSjLyz0vD3cQmAYugVlwGCMf51rCBqraO2oqS+iPqugg96DUo/iSO2ai6fy7dF
6tRiFX0Dmw97pg/WxWAb6pWh+NitbOxasQ1LK0MIBTYKBC8aDPHszm2mfjS0rCnW
eFe9OhB2K2KrPpmB1MiPXK3Enu2bXaGnVl0c8dQeMwv8xMgYgKNu9y5Uw6VufW7O
lf4iidskTsmBS+8BG19q16GdCselQPvRQw5reRXAkaS0hpRjajqdwX1sZQ2nutrF
uDA+DxA82D5JyKvXirCC+ESuNLOQo8x0RbqGxL3LgGoRInqi+iXkY8jCzryRrAf2
wmAsfHMELCS+Cs6IVskPWhceAabsdQ/d3AMiu/wbR2xfS42WAPdrbUUFfV8ClfnZ
BxsKymHnZAujDGDoa/Kw4phv0ov6WIfD9pWkGpbIHaDcteRr80Sleuc/j7Q2cV3H
f/ip+dgu1gtdvOoPLUQg6RP5buL0t7E0cmuCaE6+h4kT2VsAtvZ2f+xIcwLriiKc
sSbeI+LY35ijz/MATTk9xKbRZHgeWdaIlfeXj5G1IEuF1SFmGleV/4Zld1laDSYx
Q/3/a4HEO80IPjYQMsV+/tc6mpABYUTTq2AF945UYVPHnkYQCkz5q4XMe50BsCAq
aqn3N5tbbKPWymf+nwWEyxhngv1Epg64k3mv7UX/x5HaJoW2R8C4Rt4KUzlRxsSr
lv1fkWZZduZ7OL+8+1O6Jkow/FafcnNjoRm6wlU1nxkIBtt48lV6bKOS5jL6bqR6
7HdbU2bczGdLP8sUoIfUXvC7HkKUxoyyjt+ZRy+BySZt2oKDUe8mOsRF3p+1v2h3
MgLbHl6YLc+PszveozFO3i884E80CWpuGheWTOqQy4i3CbvyE5VDAE9HC0B0Uroc
XFZ1Fg4U79N0gwi23kUrcCQD+81TruwHW8CISd6wrSoE/ECz8Mdof4MqGY8at59e
SdmT7etfCaSN/GgeZyCogjxY9bwMXes3M/MAmH+a0dPDsVq5aCQQfS/SaE+D09s5
+RSjUqR1R8ritWzQz4i0WGi6FOuzdFDjo8dmzGKqD3xFfGOnY0ZKte4nbdppJbkc
5ZmZKJPLG4bijU6tYJpD5m6ejql8YgpDvmdqRNheIjFMI0HqcCSnmHoFqPc9i/7o
U3yYG52/FFXE/flwM0u8Urz2sHiecD9+wgSzLXCdHrInQe5MQ6RHPRI6ybwVhwZD
WR4E4Dg9m5/MZe9OUQvDVkkMew85rirOVP9z9UpZFvmTFnalIneNyqLEhYlkF3ph
IIkEae77UVbNPR1XnPLZpyMgQQ+Gpgf5dEcmybsCbjLzgD2qp4WYKPsJwJC2/GHv
yuachP5VDM6+O5gbQJexJktbpnHNd3gWwv7qRz3ChuJrIl8HougvQqwCkHan6m3l
itGS99OAMzNodK9LT2phPf6Xwe8s7W/ppC+VApK+n4CDqKB8ygLttvy6z8pyxKU9
tXsg+E16M34aeriLksegbIQdOxcUuXNpdVhBZSbE2u8KC00CSYoXWV38IiTgmP8c
iufiNWwdFR4zQcpNbQKRHOWVx4zmXYAfGfiZrqA6hbrJunlI9tI9E3tc0UPEn9jo
jkIR9o931n+JjDaWUlr0pUZSV3mX9qWU356EFG8RJwEx5GlQA/7u49G09SXuai1T
dS3qF3u0xlRR79qiBi+8yZrCUTVTYpYWbnGi578xq382/a+HUEau3KOtEsMYzw6u
4WmqhQZ0Xo2OQUtorBuX2O4XD9oMcCDbbvVNpt1WEYw3exEw1FfTOJmY+Jv6b9rh
yhwIZVXHetfwGoxj5wtMv+5ZhK1YUhzSNMbUXCXonHRgelBujOv04I1VWn0+s3Q9
6fUjuNhr98Csgn4Ey/70GMCSfxN1d3GvYoH+V0moJ50NLPMeutvWn5JuAeJ4ckjW
kFKjJM4FbM+S9atwbpuyRRo6gyePUDuzowpu5wxRo0P8rgj+LffIG6pt9TeSNWQQ
ZiOzW3ERrNIOut3vZb49UenZBZnPT23qdsmRzjvi1QP9dvjo1k/ETU5w5y7xg2hn
ubBpI1n2X0lC/68bBRSBJft5aFJTV8gBDXsIUx6AFfCH3xLn6XuaaTPnlTL0OX5w
61jnO8yk3rnk/CiAU+niC4ErRKJOOH6oiC1On7V3zOLHYiOUW4fEiUg7a2liPl7o
5FMEUtsLKTaWJ44Jlegpjs97PbDuuzFcHU/SJZC4pcM9hXN9EZEtbFVOWukvQ19M
C9bNwwP6cBKIPHsH9R3MFJ+/Jam2Glq0sRPe6yPLBKyq42DbSNQU5Yad1vO1xH2w
JERPgihoAdzqPYXqN6UyYuMDOhoEQ65+9jG+WoMdu2Y1AKUQz4mHGWjekm/FJaFx
uQAG7P1bEKEqCs25/nqJKwTM02IXpgDzO8rPW6Y6yOw4/Tb591mVJn3hMtPNDJNT
MOdVd/pvTI8pREKVl3/oz9ULeAcsLExw04+UK4yPZ3F3C29V7SFTrmAAU9hVMs9t
abYQmbOXT5htt2ZW02F7kpsjo8CQ4D73sjTYxpTZN8ui1sH4KiXUtCY/PjSoylQ2
RmkiYSAWf16CHQ/rYGj6Lsp/NyfVDsfD01qD2RM584mYkw4uA4U09bNMC5hsEvo1
IvPGpIYL39c+zzXcijh/15QbeDNRBOe2ZC28ameEr5LQt4WA8nG1vA1bUL9kwpwL
uNLGCQvJaQyOAQLIAse00weEqPkhAf5KG728lOFYRRHq/n2SEKvrwl43J1Fzklpl
0PsU06NZExjOWjq925ig0/6K3D/ZvHJghJkH5AKJeiA/ZFoXxJBhfSy0b+aN8w3o
xdYnGLSV7tVnR4MvfYU/yMQRlRvoyVO2yGbn3SeeOegj/28joWEkRBa2LgJz21tm
vRNDWNRvV+0ybgv2sL5Jixq8N3i9bFiUt1OrZk6uKOKWqlZfth5xNwBGaa46XC1M
apD/LvjXxtjTuB0D0cc0WRsTxN11P3hD3tlkVESH0sWz+ooZqvsJ/cKBYZdBzsVV
bist6KTyL/EcKhTTrmm3Lpqn3lZ9mATIuW0ZiTMseFParkq3VNgCFmc/hhHmi5Uq
1ymlm1AtfwaLPUyo/PUpduWfLHHn3sKHrMpHI1zlZrt4OeoiFBmo1/Sp66fIxcSF
UZ7lX+YyfQIa7VuJYIYx5BZJzNmADGTREVFF7urrmRTcr1yig6VcXO3ozwW5gFGv
FEU4mMEj3s6obLSx/91eHRP4cvyJU6rQFS5KF5OkFjl4zSYWkqGEXK2MLxuERJDt
LFMdATGR+wIvOkIc5Dy0vmQhje+/P5XknlZtt5ZRv7O/nDciuaDuCcFqxQpApTYA
e/deXBERaKcYqIPaqH1M/LT+5jtWBLbun4xpxr45ASdYIykChGPmYCeNtnl1InbF
TGpok+NTJIyZBC874mNlaFuHO2m4nSQQ/tZdcCxVaDgwCq82yhfLigJ9+WkwS+A7
E+lQsVhYKena+W/cntpSk0IH+WbUizv6wAApVLE8Pf/C7SCzTZuOgPuacrDx7VIv
htv3/RNR33Bzv7vYoeVl1hFmKLofRc7ms9sad8BbP3gyAHfEiKnm59za9gt54+7/
mpzG0lohYJR5rPHe6Yy68Rs4HUdEKc23nsFCEBrJnx/UYaFUtnDEaZLS82PNVWEJ
zakGz7luR6VWg9imTaOkdTlIfcj9k0pEA/RukkGZ1snZYEBCFY5SgBz5d1kOrdJI
MK0h/qQtVnSn1e/jmho1+ilvPtg3MSBKgLFc87YI85qpCcBzLY/dv39mDNH7fOdT
68tznF4NrDsLX3N/wp5wOxMwelod0fhmcWrhKey6B9+1e/PgjRmPkSbbWvwtMuBm
cqJH6nIyO5M5mlKUZxT57hRGpLXLNmOfH/GDtLhQSBAR+INGMogFZKOsZHFYhGQ/
cD8yKa5uN3RE4H6HRddCXgcP4kpU1UGqYF2Nw8vNAU0JeyglhMDiYkgy0by2d3II
JBCcHpJWkeBMDkCcCiSRMVNwI+yWEr5rgdz+0xjSJnbtpWAETDknqvjLj7YV4Ltr
4vJ5aPn+VawVH/UrE+z27VMjOSKe1VSK2sSBRGb/CalI0mStDlFEGwNAt0TLuRcD
YkrN+vBCNiLgeSNXNa1cQstkik2WRHXG1jQnlpsZSyglbt2fNzJVCD8Iea6qGTdI
wIBDTe6tLFyNX0lJJ93+g7ek8l/iFdUf0++XVdzg0446BmmCWyhsZMKwh2JnVk6L
FHwVfejcT5lLzaAJzP9eemE5XEC46cPCX0PYTLjeNcfbkw3z3qXe3h5OPqYoJnBl
3g6+P5bkp/ohZ2TsOV/yvebSjGyFZ8WtE2///YxtSrFt7eCOek5uLAXbJL7JCt60
9EVtVqQbW8ZUwEs99+akByDwiHmo0M6Z5FU/ZvXA6orXv5RuiCyxCBxruKorccBJ
tg6g/HlGi5A8a/i6Hq+SFo5DimBxJnIYqKPIRGWUEDCoVATLr3QoeC6ctrw9uN1M
bhhTMoY4wEPiP0VbFZ6JSYOUkyumtqN6kizM32wTe5qhBclYjAjshQRLzIdabuPL
5lAF7zOhptm5rHrQe2F6p9QzARe4rN6/GxKTue6N1/xXZ4HSmq58lUIjUdl2f94F
5X/8/6f9bd+j45mWCCD+7eCqLy57jLstln82OkCL1AdlwjwQTcwYiI98dKqvsIIk
hSjq18LKA77Xmy/iDGK9VyagAuK31BuBF6ZfUrAE3lgeWX5+bIAdbRgcNK0HzWio
Py7nryTimJbEUPkIKZIEBb2hdRbGQXm+4X5fcokQFe3HMQvJZg8RDi7IdiYjyO3L
zMIcOMq/s05T2uyPKr0daeWsWTfiZtNg2clVpeu8s9SOMPb0c/ZOfXscpsMzFpHc
HOUxNDMfbBdrhGrJCvMs6P/9YADoqy0ymKHZcyvzaevyJiX7o7W2uy10kh27r/tt
be/6mUNRdf7b7F8VbNlsk6DJbriDrgBamuoH3p/JolrquygW0wUX3RsVRuqg5Y8s
3yA3X4LcbTkwWZk+SZ2rfKzOVTfrP/9Fdt6A5bbKjijfc3oJNp3m8gBbbNQhbVDg
pcDLGWcKotZIh4+Q4pPIeiaigC9Fa/P27OUs0hSp2tU3uYsxj+n+pnWAy7siGUYD
94hR2JyFVP8J3aV4ubYLJaWPFVgHfUJl7mSe4Oqe6dutLKg4DbewUDQqMHwN5oBl
R/X6HIvJ8tclwoyV+JXruYpXQhg/wGK1OV0knVgAYeMUyoBcdb6Iof7DsiOFK+3a
6mkagKt5kI3blZ7e0HKBRkDs67ShF51QzJ7dMaAogVm6WNHRR/18RlihV6F6/1RB
20a8H38Vgf0+1N235YJVVToOZUiQitSTPT303upmZv0h7iin8/8dfBTpkROhu1UB
J0GZIJ3ETYUwAG56YIGc3+NShnIqxIO3cB2VhXVNAizUZSa8dsi2k+rQ/JP0b29J
rNh4VMJBfQGH1YYxjT4hotaetiR2upyEVbwhB7Z3hB2B90vaIN62uQvp+442pikG
GdzhWPU8wWvLafJyzoY9XTUd2Iozku7gLN2TaeaCeRoz9ojdosSfYygFD5qSVRAY
9XpM1zA65vDWIoeIupHdejfB0+pvoqYDaqCzjBfHV7lXTe2E6TujGkwJqxjAC1LT
uYjkkX/53ZvZJRpFcyCAiu0daZkJhKwRhbUIFGhdUYpMpoGwTFM+1/Jo4mkHGS2b
HGtU272Ep2EM22eJGecbsVmX0tJAwklxO3he84YlyS7Bs7MOGB+3A++jkw6b6nXE
hoAlK8e14F4sKv2QHFEZYM8jrn7jjtdOoekJFzrrUxzqahE6oMSDbC2Ex1Kuo17x
e8uQ8bAsF4TYUCebrm39K0/PZM9jvWfr47+o/Wj9KKRWoluhr7JjbmAAfPiXFcy5
NzGRb4OYoukAs+K9l+9gh6szdNn/yztj4kMPxWANmwdXk/yo2cTIyhEvAPb7/gYc
S2SD3tMUlB8oJTudq8Bsj2p+8L/aQ58Kk1C2nCBMsgNGPT47yVI2vchy7X8rIFjy
ojrnktu9dL4oU4SOcqw71KFSlbJb+8UlIg5hF3cFlcgyH1FsgrESMM2vLSdRdMsG
7WORrXQvaBJde19pvb5YCs6+S1BuJe0aybJthc7iK67ntNCfuTmQX2VjbQBZ5K2Y
394GIS019X2W/KNA6ieSsYIWdsszguqFSxjLXcQWcQIqwfmvb1WTeIlyjHn3giWT
31Dgm51bIMkpOki5kRq60FXQk7ALVFdiyIESvxKLA4uYYXXD4YFksmVSUZ+Kylot
4oE//D0oQhvckJI3ycj51YQGDVHXvXmO9tIJFptKrq3snEjGttxBXG/meP6WgmU3
ouZOAcWbJO2kQvnmeskcYxYzQHfFghHXfYE2nanGcfKWOvQwE5iVKOEWPXzgin2a
K97JoNq6ypT44BuwHHs+mA6k13flBuB7LcDIVYfE1d6wtaShTt+o0o74e3uyuUyc
KFDTZf0Ie4EOM+UaxptV123qxhAP97uP8cj5JK7pa9EfDUWc/JREJPVAYCiOIVP9
n7tN3bQcMPZ5s9vBt9gCrm/Jw5gXQwXgjlcibJq0RPcjYfN/UG8jAccRRcxI0+Es
x3xUdh0HKHYtVK6e8qNl+kiN0GDEoVdJO/1q/EtrxLdpST9EKA5zqji6e9ewtWpF
x74qZmqFVVbrABI8WEwWDduB662g2Z5S0CesRQnF39QxFdfbtg/jlF0iRwr3cuv4
ezNsZuB8iM535WZA3WSy+TtZRHYCoDDfFfF/V37RHzdThXM0PvE5LV/dcQbdaPfv
DjyiLmPEG1l0CSqTJ2kSUFKERZ37EP4yTO/qx3U6COJqbrBGsHZs0PNy558zMdDo
dmoORbPD69UFPYltqElfZWxplbXWkzpeCJwbNJzWS2zhrBu4vomCAdAzifLY0wzE
Ryd4QKl3pSQKsQs2s8bOeFgsWOZb3phQM0DyqI5PJSwVeBaV0He2QzgbgYI6LNvf
JTRqawQNau1ZmymMsPbc4N2TayQxg1UlWcl1WZajXu0zXr5BVbYZ1YKZwwH6Fg2D
Ot5SdQrcvlveSY5fd3LEKZanNbLqjqaAvOuUII0YEuCVGjFiO0MDB0DmA7w2GPa2
Azg1OtLlr1dwxhMHXuniWsf/VPsvVoD+VtrZVs0aSEAIq9wmwYnywOPRrFiKMWOp
w6X7XNDOZoCvmK1i/b/tnKOZmabzy3ApLpoZciaVORsOBePyNIGugWVCoyHPXhzG
ff3QfEXx23rybpoaX6U29oVXW7UqIDJmamaNlNzwPxurwG/JsGtz/pCQtJ0uvBpC
Ht90gjAHpjmk4lM/oAehu08w1mX+PQAuo3vYTeovKbuK5mQh4fSVEUVnrpEKboaR
s8F4Xqvg0EWzeRLuMjsF1CqlHq+LTh5sWcDIPX7q7IxSwITbnOUksJQi7BY9YN3s
JtuYA62BL8Y03U8vGKO4wLp73mZOARoZfSnSFZtSAc0ppWkY50B88ANKiW3X06q3
DCf2KbMHhw8J4Yv8tE78x30lN16H2TnUhuWzWmRSkipECz1zAnmGYi0t9xvv2vAT
fXO+nSvGCoHzhqvKUImpTv+rMZ/FM6U/N0Vv04rjduzd9WV3zGFdXNnyThO5eAuW
5AA5CbH3F2AJU1OVjhQbJLRJ7f9/Ue5Kv/GN5lVxnfCFiptqsdBmB4jLJPtmjEYx
isDrIKDoWpkqurwYQGakYy9Mkq5Zw7lqaYLItN0h4GWXECxHa/Bj5q45hyAJ/fTj
+Xq/E5z5BCNJIzvVatkKC6pzyjt9PU+zFKn0mlLrLEpiR3PAqoami3i5qI/gVmIl
QOifF9x9eUtM/0yAOjEYRbG3xCeaqo0aHFmqyC9HVhJJIms9lDZs5tXrOQpdkxNt
OB+jAQakqFnpLPcCwvluvoHw4p5aMAjkvcR/Sdbvusbq6iDtZuzQTZCvT9Xu0AgE
DL78i7Aoe/z4CMOsM3yv/j7ioY5VpXfcJm2EYD6RIuuwxK0dDRN25KOOjW7i9ukN
cisrr5g6rhosVMDhSLP4kl0JI3XLAFSlRsDbaZ9yS5Km7iAOh6TjK7lyPDLDeaMn
JRnZnBubbXyPYcuct+2XSLs4okeVtFDOVL6hpnE/0Rd06SIhHfrNGRklpJ5daA44
gocBrZjdS2BZYJKGZbZHtPqyIkR0xPap3byaZl58G/35hafz4gjJpRh4jN0Lgxzt
NSuw06jhZhiVmVg9pvFsjAtwbdgoLNb7faWlTMutpdyIrXQE2a+Ea84aijRgjRYD
Ne/84FyKQfDkCEzX8c0yo6b9U6ZqmDDIFK3AA8SC4mLLsmTBTZnI3nnqnToulR6A
pRvd+vEXrLtDYXo4KdcK3v1TvbSHKq9sKxkIHxu68le7k1oWxq5QWEYmyhlz79GK
W1m1GpseKrq6MhLdTCYpS8UL47nSV82JpnodjKynP1+AfQODAUj2ibJ8t5eXFsr2
82E+IsbftiCHoCTHJY1+KJJY0GvKLVMcdAoJ89XWSh770DwS59aDIosOXV+TZDLv
c5vvBJpW5dWqJaC/4jOZZeLXYol6BwpN2EdAqQ3ax4KIEImhlTSSX9J44vLihzL7
+f7NsqAq4ZmuQ2p5FaOmJZsbCh4WumYT5Wm0FXB3lK4R/hL9ggbn+OeQRA/N9RXK
DPIJ5l7SAUCl+ovbyYtqIF0juCaEUwU0n8Zv/CAxJNJ2Txmyt/zDQSo1pRSgKuiq
E9EgGcZHHAEE9yv8ST1Pfn3W7MSA4eZVdEO8Zo0VLlbAOMtDfvWqWCXxYTc1t5Wk
i0mrd3unZd8cD1RzWZajM/rEBoz4czo/saqTCmKidvzbYHRPwjG7iL3ByZYC12ou
5mTaeniZSQN1xRvY2F7HZNu0WbftvtBtXt6WcrwHX/Pgvvrgsg6fDPW6wF1kagz/
491hqw6dJVefLg8Bk7F0D2pZZ5mIkoTgzlReRp1mBr/vhRwYnbZLQnj4ZMN8NrQe
8Ivc5bh9nSVSr411tK929rxsBWyIxaAab0MMs+C9En7TesfalEZ91JhTmfXjsudL
QoXQPxQxwNoVq+gyqaZnbb7bcPQpLbyfSKC3lUuvflvBzOt+jG3pgpLdUBs3YhfR
ihygXGhGlXcP72AeqqzPgOAp6WemjEVqbft8YVi9kO/mzqgV6Q9nJ/WH4PlsqMwF
Xl/HngyXHLIbZz7eNS2sp6dal+M7t+eR19f7tfJQey5lpWKBKCEvRwYE33hQGrGj
ETs9vo+tVghnUuGSkDfBRqOdcwSeHytzoHPCikL4dNd7Kpq8ebNmfKcOlOYAgYW1
DcPLYZdttTIB+Fr7Y5bu/EtZ2+emf2zDA2CSUHUWhMl28xMe1acKCk2+7f1/H+g9
VKrpf1/OXzkTQSiJA9mMHnxc8h+cKytYhkPp7tblNzk2wPEt3/TNDVqcJNkL9tbk
ouE1wSqMafgTUW+x7YHzgMj9i0dpIRjZLOEzgxFVrRdFuNH/9k32I91IgbEDxiky
4iNhJ0Z7jR76xqISpjfntpVjRaSJVyq1v3gZjMzI3R5i4/jNoV2xVLrvDY9gg/Om
d5tNR+mFpym83B63EaTuw/zj/EiiWPvxOsAuEsYHxlKC1FTDqLfYz42owL8XiAEa
F+/u+LzS4K7P2YoXVgNo9YzdnB1gk1HMDn+5spLOvXMQ2P+rEasuA9mcNEKA/TWZ
DU3chZe91fOJC3cfxmvnQGHxZhiPV/yP7UWtWK9bpuzU7+iiHywqAbYNxdAp21K/
dlDGzXnfDXX/6gQIJTpRc0ZKaJ6otwAGoFC68kA2hhme0q+vXmNVQaODutQXTYy6
XVHvPfqvBgx74BvFMVRql53xrFmQ0rsOFbEJiDZDBS+SSQUHxbF1XGzB7NrhTSSY
F9tbf5yZLrZKSeGHYbdOLDxexf+H/D83DZjTgVc4LvmhvNlr/XSbdHvpi6Lwo1jZ
9yUe/mQFb/aMCgEgHy/2QIYdP/I9Cr8rbU8ZFkAN7H8jvOd0dsM+yYWTiGK/Kgzz
exWZs1wywtyy0R73CucDUpwiRh/4FJyN0IsZBUqXh8YF+U5WZ1nf8BVa1jl3Ztm/
vvFRrE21iqFY3eJRWEAesT9IQEPjw/EBn3fuEjbugzvOaxEL7cFnhUxTfmoYtviY
6wOXk1UMkkuIQPKzlKlaPA8w1u4cRrNjVVDmdcSGauxDvAlK9lyKD31qA1Uv0J9o
Ui8jDcN/8tqmCnhHhzUxYzX7ul6sPxEkjX/ogtBUts//kcrVHMbeoWoPmJAdoqHV
LSEBaDgJ3Sm8B0Zyx2d9D++Qa5Sgy1IBMlCE0eC6Z6t1OoAibxH1lqspwzfVzGYD
dRvi7iSyblGPCkgnUDK5hWGLYtKBWMV5u+wIogFifx//EdX5miqgDT337hHlzeHL
pKapwMcOwLLDSYbTUPH5+s8IOrEroh8oNrHYvnuV8/0b9m1z9r3RM1hoL2JP7HK2
RN+57SyRviZnJi6Wvqjyb6gNHCKjYMLXG5Abpf3FUiIoKsiIgw5Fyw9elRYX9myx
mqNNwZlRXrVz7ZqGeXoPuf1YuvsF63szD78//K1XV/S177NP2eGufzZmPDVG2WZv
/smb4/7iQLTfAnlHpRLaA28HDzWYc9i5KXCN+iQK3JNZ1nzpGkE1UpPB7MSlCeSC
VeaeQXXuPuiDY5Sk1fUpNZcNck1OG1KWvhGQnzu3S++CabBLNRcCovXzOwU2+xvH
MqIBWTy6VFWBUVtSRgPqnSFzFJQYC2qicFWdgXXtV5V5adY4EWHKg49xHI9zU/lB
0GRTUNcc2/eZdJaSjozjQ2Fpf0y9xR+Zao2N+KEmZS00qEUX9Nusyq8ZOTre+G1B
c0lLL9AukzyNxj/9BawvI/0DXZ8hm2hTn9hiUZWzWudYty/BY+qEpwfNv8yLeMiQ
1k3zXxTR18HUGOin0c75Dj8orjtq3306AxjriFa6WaiC+JeavSbCzJkdFRe/OHQw
+0gKMyTVQyUWpDQF7iwnxoEJ9HIU5R/RwQpu8rTD6yZGN/BS5PpOO/76fWpFdzQq
+kSFeu+IRkA/9O36s1lAmlNq5ncbG8bWczin5KZpLJep6YByKgnoyW3UsxOdc2MV
PqRioXDLgCUCzbffY9tmHbStjZk1aMD81sjJiMT12wqdg9/5MEoKHIBFhlFRFSM7
b2BTXUGvWryCLrLXmiqKsGesjtc3Yu1xSbQjE7yvfkFo8OkWlwGushnzMh36ubNB
8cXFBlPYKSYDkjXzo8X2pIEsb7kkpp0dUBMScCett+X5misQzelY1Z5c/k0ospke
5/a2csVfnyvJupzW4OoGd4yq8YTeS/gVAuphTZEKDcCiQFp8SD4CoV9R+bVZDavG
+Ft1DujAbK4/rbZArD6GUhS3tITnTegUfHswzamTb97zcuPF85vtAYKJCMfhfpw4
dHuXxW3VPTQ2S9eoaLPCKbnSHdB3p7fdWsqujJS2JH4/scf48nlb+SoXzVrUT/dG
+DlxJ/QMnZ1o6rCkxg5FHyybA12StjE+BCBzMaLQihPfb9swA8jGO3NZ1R+0gFoh
zrCTTxDIsXH0NC7He7PtoQTinYZMct0Jwn8/TInCtR9WFU4fXT+rMGtMj+bpnQA6
LFyr0VRIdgpqwV28oqYOHP+FURJ5kHfelMzbof42jK8BnIvuxAgd/0FqsNezqnKx
Vb4QV/u5vxRA0j4pe/MLkMQVVtcyldRksEqbBPDg2XnGgtW7GQT5eT/I41GqZ67+
mo+XSDPWlXXlkLdhw2PbgUY+IIBeyEfSWV//pKaPzJSlq8aj8uJIVFB2pHuyy1xx
S+tpCBdUTj5MSA6VKbkZFV/OuRYWKnLyh3QGfODePZ0xrHGkJgKZPm6F6rPSdGRx
5eYbJuPXtMxUSzrPd/yH73HQOUNLoeLfi0EG2OQpj0dj6HpW14017QzrWNLlzZs+
DE+udidI+PFv60Yz0SIi3u+YUK3Kw/x9mPqXf7ot+oU0Mrgl2RDgvO6X9WzqmW8S
UVx0E/z4EIG9yqENyUJ8igSo7q8wJ4S7YEABQgY67mpr1tT2K8ffXKe79mJHVIpP
IqS5T8uXD03kTNb813T1aHKgme5wEHrDOHAUaNFygn5WcWCsTTi2o9++4aUfb7I/
KEOE4UQjiiPxbTy1tncWmI+mTdQ43AG0ZR2UW/40hriJosJLTd9I6DHfFkFSfPHJ
kpFGM5eVEjHGlZHNAxzRl47N6iytRI5L0Uf9rCoYzk9ckGMiRZr/GllVxNZ/bzjN
Aq0XaiSTzBHdsOKZEcugxMysgVrcZR1w0PYcSG5oTfxPyx9Ns08LwqORVUaB02zW
ROX7E5iJvKZi63TXJJzIVlwEk+i9K0PP48Bi1RvsK6r4hOlfHPnbfjAQO1mzpSNR
v+6lQ63oQxoGz1WCrNNbMvU1lkTlZyXfdQSN5hTSts6E33qk3f31+eNXYHLHFqmn
RsVp+11Tok+UMnDF1NtUB7DCHB5cWeihuRnrONpniSf73UPBYnig7YOsLWrVhisc
aUC4gqpoUv1BvsoqMZIvz0Z7RVCRN68OFw1WPUWUcTqw7NbeoMo8ajr5x5ptBd8Z
EZgoW0MMRHd2aZQnAIaabOWDqPrQmDlAvFYVl7nFZy1/bPTGygG7W8Dg5Iuub2vM
ChcEhyoTNDlIRWoNpPYlXIZuDzE5dbF7TH8cQT2WBOvPesoVY7UOADZP5rI23Z90
5kJWkSWaqGM++BZAwLS1BU9epDHQhOYVq0pNG2oIsZyeNaW1GGY/yOzmLsNPjYHz
1FdXjy5PGFWOBmUtjMaC2VKEFMZR8+IqS9i4aBrYRcbei94iuxVIC0ypeloI4KfM
vN1NSFzNiPZW8w9TbAla0oYCb0MDWu1KrSiuWh7m2rzBlcJxrAK+COXXqBGJBi0t
QpR3w5jLFWESOBha1G4I4zc1bOOU7jqdWl6P4Cv5a4onYcC1PFLAsF+UolHXo9/Y
OqlXfoolRd2Zhg5xnmmRS94yNLl4st6JPplt6HEQByRZ/+sEovTtk3kY/rKTV822
n85sEFSeUCjJAuw+vURH447Knqj/svcFP54UdyuX5GBynuKF9oDrusd/zn+X/Z+F
P6tAqtpS8AYfkd0CjI42fFjgnUUETKBNP8ryNrR2Wq7hUp47mMYOkHld25ifdwrz
VC24akjxgfht9RZyZ9hqEaKuKvr/MfMtzugfPSOMoAUbielYQtXqoAIiuNZ8/qFA
2dEjM+sG7EIgJDXhenVr8qj4P1KQcXG7NP7Y8RpNqeBdtwpsYrdTbjtc8OO6+G1f
bD1GY4A5dX+rf3oa531ky0zsoYgOoa4iikGmBmQr1X35Ey6/Iy/TxtI8gP8nFfR8
MpOL9iArRz0p0vGybmccYSY7UzDDKQls8qU3BsNPnHlO0fZyB/2Qq1nE6R4wsFa7
G+Z1f/RGW0v3UxAChmNq9u1ScvEUMnCV/TybMuUcCB+A79dAPiLh7DF4hTX4R6gw
3hGtmfXY0arNjIaZy2JtiPKfpvg8hB1iDsRl98wL080ld+EeoI+5VJDwqTUMAHQm
GesF2THVHU6Pdo48lyXmdpH5EAqG/GnJ/1lEQdk5UC/H+failQWpBOLbbDjbgBbW
Kym/8jaylpJaGs5wXSnozqLRGt4zV0O4aTI20y+FtESjyi5SYvnrmtVIMUgxHP3n
eApt26Ian05j+QENIqTE+2wkksUxdxl3zjrpmkBrRFuQXKUapw8tPDE9LcOl7vum
Wt71XEVFqjR3LQ7ys1xOR5HBsGiQn/qIjmViYC3qNCEmAXyxI+XXSmn6rUYIlzfp
+j1vg09fhX3xV/hgBOv7DuDO8T/GYQmfoNbckitRyeuCxm6+t2PP8VrehhGIorV3
`pragma protect end_protected
