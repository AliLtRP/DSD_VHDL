// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Gbd4P0hCEtxnQ60QwAnPifTq1brYeFOTbmCdIeuflMj9jYCcjxp0WIXWOXwUxiML
Wuew6KJ6HCXcWebjf+Z6U8vGjtPSHujQTEfdTf+ynWnysASslf83FZ5xy+zuB0jW
Vr/c9U2j4++dxIJfuQfpR3ECMIn57PLKbQuTsvHNCAQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
Yc4AB7a1lJaI7k0GhaiDTb7FuZz5tz9kQzQsJ53Zk8D94cvasoMqodqjKTcJphJP
34mMlIzmZkzo2n+9KnFrmq7F5S4xanJxzJJ1nSSVmTVHCx/TwhbEU0Og3ON0TW4l
zQFdP74zDAGF+4cvGc77DprcL/QD81fsiMsDO0S+59mY0inAAkjsG+MzcOwdpsKL
B5C08060agJkzavcHkT905OMboPhEnFLGMHLfRwZuqdLlWFbCo7StLTB9hYbl+Iz
SIN44Qh6E2ev14mI7IjQ+HyTQ+70JKUE+3UUpRcMmS8QDsjONkpPs7xe1NlbXgoU
ww8po62jjQqIEArov8ibyupafxFwKTjdhEiieasrcuw+n/I296KDH6WRKnkRVXKD
cWG2aV+Gg0Xd/RMo8Qeq7K7LWQwfLD4DMK7tjtejqqFfEouLvhnT1Ok4UTAUpRnr
ut9OwXsJyig96xV3WgFbLj9yterEqrvyveALQMkBneOSVPbSUdysy7KidmFbjVzQ
KzUK7XnavSuXwgiM1uAdv6LOrG34aRSv5pLqyNEoqfaBn7w0dGhGXkTKpyfGZ2Yj
lMQ3IU2o36s5W7S3W6HvTl+LCsOgCrg4FfY5Wk4fgOdk7U7Hjlmac0qPyrEVWNbV
jYJ0q+95foUwsSnrEq02d64WLaTLTJFedkBOBtEcdfLgzp6NtDHzKg7F/Lof5eLb
2cW5ezddsKf9HRmIjTKOCqkEzfa2+PPlxLG0nlmCIJ7ULoa+9BAtrVGMCSVdK+ED
AlCT0lgG0/M4SW4CEQxvi6MKZOtBOJSDGEupWDklTNqOQkGZ81qxPXFsw6Zpqegn
PULkpjO7X4+WJ0hHF7QL1/3Zky5Z2TLcF8PHOAHAZpNSfb4Xz5RDWYiPltPMhM+D
X03xHx3FoJ8xK9/y/RM8OFJhfa7EzHcPI5PRi2pqk1LLy1zb6v3RhOa48u5xSf6a
mfYW40dGXkuSjfIkHwoh1ddp+3l7oSffA1E7MTPq6CCvEy97sxh4MqeNpPfFXi6H
EKMcyAXuG/1FnbVkmfXvQhmfToBOLODe2NGTqgVzL4FrNI+FwHMUYFHCBE2waUuV
R5OkVhBLKxry4dlc0GhYQNJrpCkAqnwQ1fKNx0gSecAiBHxrz8n4GB0aOwX09IK7
wzblw+GHRvanzncFX0FvHsEy5XaB8dYjWU2xXQGBOdxvE4eHS0ZaXWe31RT7rkHP
shF7rFktn4aaabp/pYJSG1U3v0NExNda/8R0ZK1gJJKTEm8m86h8t5XX/GH28wcy
RGiOJBinvyxpcdeBai6VACb0Grd9eIkIU0ojXdZI48lMoqRV+GzhMRGAdcOIksMT
YyYsTZ9tLrwpLLHF+4og4M3okDtRiuNF1gdtTsDGgjMFg3HSi0ZWWReOmJ1914ae
EHgFvYJzuNQJVuAlRlfdFImw5CXokC021z4tyDFNHLDENbhIlAZKw/YprQLCQsOe
qmY2zZPaw5XPpXKQ1M7DlBIiq7YwUAnzMv5sZaPTJYcXqDzT+0jM8uq0Sc3L2iTs
piACqThWjChYsZcvDB43sfMyIE7p84NuSiBfiIGW5NliVu9tNp5TIIcIneseQLT+
Y9X/njwm82784PXXw/xHK8+xjYV3BRHYAGBKbXJ19ZW0QxbMorBZJtdk7WMbuzIH
IuLqtoxr1nyjXxBTd/b3hIYJzajldyVEghBIPuojuMYTLU1P55a3WkJ//RLowAJm
580ukbOV+M11OFucxYMt066yN7Ikebd0bxsDCPPQ99bhtGuVuVbX3feajpg+2gPV
14RpzhU2lZGiXv/KO+sltomrPJcGRbutEG5taEZ6HhjTbaBhpWL+kpuud4Xn1JGb
EpwmR2w4B5GU0/ooyuqtUp5hIUSsqCJ2voPSYoS9iLL2y2SbUw2IcYzek/CBWN7Y
5i0P/5Sld8p9Jx8ubU3FQpW9F8EyNcrEWSLTiqvWe5MkZmh7jKptEwWsMDqe5yuR
WoDWD8/DPuEMc0zCWGucJRlNdfv8nAsx4aRchLzIfgJXvJfri2tK6GTD9ZCk/sDw
uFF1gdH/BEoXfSQDTDcmK9rXVDCOgz6uV9Lhyv3qzbMPQ+Th2bHplSuPkjYHzlt3
X3w/KDd7XgEV6G0ex8qnvI9e3iqP0VyvC4ZGQ3Y1YpBEuryy0mwCdEe4bwfqlTeo
CEanSAd17TUCsb48wxf3BIGvkoJOVruLGgZ5uPVvx17flUBuHOZe3wylMOTnWw7F
b6lOLpuHZMucbibHoXITfcQvl/txkekp86/x3cComTZc3qcUyTHiYjL9ANO+L5ha
50q+ov1wkiE9zAu8cAj1q0b/ZIWRSYSfXuYR0u05BpMy1GyzB1MSKaHn7SSSu2Fl
yt7KxzEQ06PQV3wCKz6cNt4wlgwPDlDirrTN26ZUL87p0eQEabyeYiyAlsnARSOG
Xbb+90dUNJSRRgYRHP2pr+pAdal4J+GqvUWkmIisAo096pCutJ73TDN5QG6i/uI0
rvEyGGMzGzrP7CFLzpk+HUk/mjw4P9ZFl+NXNKg/YRVTg7iXwEQDycbFRiLFozq8
zHMJ2CGQtEzVC5PSYNc4IfiB00Dx2fOUyGQShII/VjQQvV9xkcDFwA5q4LtXoHXW
kTRhaeJDhkhg08GX35j5JNPmVaFFeeQY3OXNi3ODJ0ZKvlCubZ0vmp2ax/vGRwtl
JM2qMxCECMnJZjt4bN3QD8YfMQNofyoPaq79wRMh+/ViXRxdy8LokmpJadfJ/s7x
N3+HrUC2ahAnPLL9fW61+fj5TKYj1PYzHEBAEXJzDCS0zsVsUuHEviQk6OHuw0Uk
W2Fcv12oQGveIzcMmHV7P27IFgWI62bUXykLSZQGTz5aPGjkolu9eiqhf6ZQJzYl
hBu5eIhYyb0LlwlS+Mz9slao8yYS/1HYxZec8eckOhWRkMxv56OIMp6GNYQPBmkb
heHoPoKETYN5aDZbYqBSvGnfLAlZVJs4VwtFJqk8ZOx/go4Y7KR6Tt3lzxfNDKMW
7MHhhW49jYwzqMD+lVjoFoSUp2yZiY6zSDoq2jF/opvP6XgeOpz1TIKvwa2rjGNF
f+aWic235ifsKjPckls2EY4xArX0gY2hdz6SoyfAKrsTz6EMjS+T8XUw3rHfAOOt
IpqNZ6a0fj8yTWWATNcYVJgRi467Q1DfnVO3nkqRiNvfhgqwkKasctKY7vD1xxcW
w5tK2NlSivwUWET4cKyMHG+97zoRN4NdfiwBBw4ht4VzmSkaDs8yzTdDLMuxBGuj
srUuMgpS64bQFmGoqgUKtHS6x+ckWabhrSo5h49tYvLWRcSHicXeXdkeYNVbWhdr
eaZx6/7bte5/0a1CQ+UyH9dm4plaaOearrvLZC14n72If5fNZEJEXOyI3M8e/D99
ol/w0iJIZ2ixxkRKJwB+UeDomGMt40WhuS4dtVUV/84vScuGRq7ah8G/B5vVr78L
eG3yCgh+2YnGRbT6UW6Go5iRSxz7oCOQ4DPhv7e5VHWCZ3/Of7z0YnkN3NYBXuPE
JNreblgpcXfFOsQUyR5SYpXb+XElHFoUn8o3fO8oF0CPORbMKcKDPdlOZsUyt0q3
xN/roFxlHuWIOZAkq2EGkhU0QlFKA70nSC2IF3o3TK+++mnbEZv5xp13pAI84mAv
eUDhV/qCJ0Bq66q/6PaK4kClU4ySix0+1TRX2hlNIJVCvR/20zFC/lRPV3efNtHE
YPyYnOmp0TUHeZ8GZRJ6VNel2JBprOv+JFp4YXFFtxPxa6uUEKGO9JdBIo3T8bca
f7BpP0XjycGrcghKegGqLpROySuQ9Azz/7P4yGHrqlkuRFhH+X6S0bDK5oeDw1kV
QjakpEzVqk7VaRc41PVXvNNkcMFb8kxLwJmMOrMCyJiYdDNL+GCFIL/xNeFMgqzx
mpEM68CObT+6dxFqq2i3iwRPl2EPlMR3cFlchvSup1igdZieyxVuq19lh9XWiOQ2
BYxP0mBQKQI3u8KJ1IKUtNGmh3ocVmA7dT7I0bdcSe+hRsM+SGbRgquCd7AfWoz7
JRZqpVwkqqrCqjcorFNHrRFuNudm8WvBALWLJ6xKSMJd6JLkdk/2lCALKk72PYUB
Te4Dw3zx/sat6ZWPmev6sTvDBmFmQQGcxvku7Z72RtkR01MoBrKbL36EwNAczij5
H9SVSxsZZN45LqTvgigJgMljnE9VbcTBheMJ7LrirGxLH8O19gDeTm+n/hp7LbHf
Wb8mzXGJFMSgGgUIifbBydalHeqmuQsccfZ+LpEBuaNI1eIkALAzzT1IVmgb4/Qc
wqddzMv0OhnY7HHM6C4jl5sgPdm0oLoIpuc5KIhHxSrnbnnyYNLdg7pp8qwqGokp
2BljEk7OqtOz6pkpBRG5YzuQoILxFyH2x+514+rOaO5VqX8Gu8BZVnOewjPJCy3b
MHwmQPDBb0bJ0bkUqME8iIJ7uCEbqB2W5aMlRn11T6yKiSeZW9Vu/bTS6dyT9306
/wy34bov24ot3y/sj6KXV/s6PMoOxqe8lYv7Vrc1K2ilc8OrNPMreZ1Z1BWQfg41
0e9xF33MqIV+mPPoxqYrZW6sp2w3HJMFAA6x9PAjJE/I08b0CvkWWBYo4uYOcz85
2oQBR/4/u49XkdP3eDtyxVTUGYsEadPd5Lw2BHPnwseJHVqHefc9EAbOvKiwjpGV
MbWdPZHl4N13TDIR6Mt0HFxaRuPqQ94cKFnrzYzVEo42VBPcl0ViwriZA86WV3IG
eciHSmCnJtv/TDe/dP7mlyuznNjV2nahR06zdXVWJ+LU12x8poTOOWzFqz9BM+e0
p6/E5rhFaPMNTG5EpHp1XOq3+wYS0x7UrRxeP5AKWPMoI2pL5uhSvRGYRBDAZOns
oCqW5x4kXncL9RmKzgMBkOSxYvEbmcmY3yBCEH646AKU4MQhVyqm9YQ9xIBO+ER1
StVO4pj9cTg91Uu6yDaJtXxQ2c5Y2IzSaK7jKhIHpt5XLUjp/lGtNqEzSbYaQS+l
poc68pRkR5J+tr282nbei7ENOLQQKrhVGFZGeUlSA60/JcAHk7A+6NSbI5PtxuqK
Z9rfgWN+XyhElTDLQMVjrIXmnTbutFSN72GNYyXm87fVuRhQHlouaZ+gpf7aacuX
0NBe5YA26HXIjiuZ9MNrXrhPkl4etQSmDtUU0FiMT69X8B4Upb5J+/yDUTGUaSnl
7mIB8ow7PPxSbtfHisZCn0fJYsVfyxwynS5tjgea39ijbueTMKDB88bEKK6WKYt9
TCn9fXZ/7AtmkkXILjS8Z4y6pGvHjXc3UidUjijY7FZhDHbgx6j0fgIs5nJxtNiG
xui1po54ZbnmQRAl9zpGZiFdyZ6bD0WtuJTM7+XaLk1pEERsdMAiXJ3/TG1fFAfm
Vw1Y1qov4QFAvJsZPPItSKvQepJOiYL2Pm/XCnmrEFFeH1JlA8ql1aAHg1XggOH7
qlerCBygvTefaTicnNgQm5gxKwHjq9Zcv+VS3Nvq3H2Nvd3cnRa8IBGwUGZkduJz
jfgPsUf67tDPOC9It3tyWoBlKiCFJpnm8WGWsXHizFiVZy0h2msGurewQ6bNiWF3
rFCZI/Nf2BQ80zgUpbSoZP7DT7hreWllxrUvU7NYc4mrVN1pZdj7S2MbaYERAn5X
fLEeVxww1rxNoT4JY4T1KQJxpkJd1RA/bBHarkkYUHKcpB3v3VZM0eWgiK4UpZ0W
dXFM6TjH0nH3rkczz4IEIcaMhMAL1KrEJh8q36IUX586z/qaBZDgfgT8kyGx8yZJ
7ho3UxuqMrTOcoXG4AQGCrqkC1ycBxNg691a5y2qJaa+Q7Q7ltP7x7k1G8dVcXV6
YqUmWqVslNrQUdLdRpILx+BtUl4rbGubAjgYRKgzI2QrCwYm988HMnynx17oNiPc
fDHwTids31UUG7r/kIH4RT1C+RP9Fl66jTkBAXPLUCRPaCrs3+QNFn6Y8GB90ii7
6PU6x20hv7YN19QP6AY5f2faRXUitguriDmHWy5gh9wJWrk7R/rk0Ug4YJ6Bd5vH
MOL6uUzVwMyLahGmPlZ8bLSS4eH9x120u1Y1C9k7lMPeBafd/gA+TRwuuczctWyO
4Q9Jae4wdcWlHZ083MjOe1sfr1F1/hh1rz8pNVIaRIhdR26yJqSrQCoOTLQ6L1d0
3TCvS+LG7JFdndm9ndQtsHGc8cwiu0nuDNsQuijfSFbPmg+2uWsW1TBfuo9Hr4pn
dS8Aq1OMuQxgHsasM0IXHNN6WZxzhjP8OI1jq5lu4ZyQsx6+/JBJb4qGPXc2oXEp
y2AaAHXQ1invdasSGBR1FJe+2ujt3S02cvBTHm741lu84Zvp2VYfUzPWzEeoNaSR
cGWH8C1BNxmWVQ4ZRZk9xizvZarIN6YgJ+1eHsJ4in3utCMC6+Y+IxPKszdccT84
jfWyxle+dUFxZX88Nvhp82BNZEy2FoqkhjBtQI7XI2ij02kzZsKrRdJ7yu8luhPB
+1GGrp2muzJsktjD4qm1gmea7rhUuITVVSyormTKywGWaBwhfgEx7a8U815HxNW1
c7lbqkODNI9ebNx4KkPoeNABv6Y35zLUoIhSkBQ/2ALZRYXCOa3bbNxhKTRvL5BN
H5V0Y7yiyFZ3VRefQ4GY5LbZV5bnf2yxVLGoA2d91PHwJqbhQAbOch3knJsm5qFc
6bfT8SYx63IqZwuayOwCZgY4Lirg65dvZcHBBOvsTVH0R3WfDKfRPzdxwmBDJZCf
BOSkHNut3JvxJKeOyuEgBjOlvPocPX6PPpyOIJUMLAN3z7rn2v0Aj/18ZskXKemd
u5pDprdpcCaguzd2gR9NALYjfiVPtYETc5T2Pid9lTB9P7MBlv5fFsP4QnwKLHse
PPvHz2zK1VbGfG0KJgUoXQBeIMfyMXmCBBAMBoOo1MQjMI9seJ6e6jtYfhyWAx1Y
Ilhqtl/2V4xXlK1L+zM6f0BeZJvvfathMpbIkiOLTqRBc/FWc4VRReKRtWKZF/f/
1U9q6ZVnRwSfEI6b79In6nRmuZqeSPRgQXA75wHffOS3SSs4N+cJTJHvu+lQhQxx
frI/en2wW1hE05uNokbVX0pVTsrslCjdpmjBK/0Sh3GX8QGJPXXYCkNgPswx5hL6
t55b1qwAwyzsn8t+qDJ8Ln0/BSegOz73OhRP4J0qX1covYRp8VsCbkYs/SqYAyqB
qWFeGeHobC5RqjCeY6qcTRdeD+TPywlrruWxxJIo9w/zsr71T3omBVl3RtHN1hhJ
0xz+UCtmV5Usrmal2kd1xrV4MH1bgbEJeYHBrENKLm8xKG9XGqucKox35X2yIB4T
dYVw72F64o8NHuIkKnAyPTSTd770G5xQcxeq2chiGb8UsMyQAn06HG8hQ+xB6la8
xsvGS4G8+WOMn4vvMlngkIvlk7TBp1AId6fSxbdzYh078ml2p+rzZ1IcsDA11sc2
7EOc54xiMuCU2IoOSQLoEwcrAWo2CIp62bZ6T0ACRrl9nEysXJQSX9mtKI7cttGC
L3QEuFePMh0CQo+sbXM9pvtbZubZWtBwjjIHpIlgMLtz+fk81M9q41eMftkR3UPn
FDNUmKr0wCiCkIImP1hNYDUXmx7QaeXx2L/ARSxNR2pq5icUICbzfYwz20VvfVvU
w7IUth5XegFwoK9cpk1XqiYUh2H7IPRvwYyFH+tFct+xDMETmGPKEz2+VySULsFK
pd3wfEYSAYB7PBXElmJnOtFkX65xAI/WmcV0OCvz1wjRO90C5mtrBVy5AUOuocrY
DfaGnp6rOzaMGJE+lT3/yC0auRWsjJkSmLQZGWSWWwTFsKb9XgXX2cXmYzmuz9UY
DzeBuUP5OHTFDa5u8+Z5pi5pzRoZxXZriKlDkHpPGLYLUXVljckRrKiiLHrPiLeJ
TSN5nlQoU4yKm5QWJiUkHHJHNqOqQ2dA/JN4fhYYQXNzhr7o1eCRJjI0LQkBvQtT
n9nbMiJli1oea4f8LcMNBgywPDtxvdM53T4O60J2X2Xu4DangSZ3f6ITLT8UdWL2
529TtS0Xd7EAqIzt/b9lev+/reb6+CrQjKvYJ+hMm+FwDTNHfFt1EczHAso3O9LQ
Ub9Vg0r/KN94pns1KueaF5xKf237ynoepdQqBnEpNoHc3B9qKZeQL21lrKBp8s68
EwiybSmPNlhepKF/xh16KR0O3v+rlXYJcE1qRbTVy+Hv+LDR17InWPOELGaU0SbB
FgxYIi4bKcYypTs/Q5hJbIE4ryCvZyBFM9ZSeSyo4fceRZW4QqQS5c7EPIv87kKS
9YKVZviuwB998oZprC6Ssn0keo9b9gRECSxLz+pFYwb6NSU9F8EjHZILZDsidH4G
NOUkNOkd1DueGW51hr2eMOnFwPef8iJZlIh5tmlCDFx2haMKOpczXeqZLP1Z6NDK
/OeR2cdurW0PHCep6TA+yVcb8rY8zvkWbYJCWBDFQsObevmoFCVzIAj5dmVVkbxp
yTkOPeHMn0KJYC4qS78CdPZXAzS41V9QbWL0JMdGu/bNsgVevA6MGThv3cFgZDyx
RLTJNqZwSGSss7qcJX37bRCdKnXcEw+HUoGsAcuoM+c7/4Gg5HlR5kSp4D2lis47
uYob0dZvdWdfxsIyUT1fg3R/Tqc3o98vQM9MTvPThbB6Cn6WMKR2NVEtjsEbdUXJ
wYA2jSfjAYVxJNmYPjBzTrB1upmFuHioG4pv2H8VJuKrY24NQKY3uCflM/z5xE+d
I4/ZIOTpE4z1HGHlY5Q+gpvy3bg65vXTeAYn7NF9Ma9lhk/PQmB4y2Pi5x5n2Mc+
KgCkR+h9RuFxlMxjX5qXbKXfwFCbxe6s5SJow9NMJGuZPF2rwgceojeWTbe8hVXJ
t3F0eEsdkln2Jcz5+MLQp9tuCmsy9DfZCim2lt7j+/g0bgmCU9CAx1EZLsgBHqwA
zSjExhxACPemqd/IGdqhZKmDtXzpTgUcQeNnRCixGNELxbe1oL5VYIRFMbmVOOHK
fDInevvEtb9oIZrPUUyTql+dT/iTM23MeowbEUdLOJrED7gFpQudRP4nyVB1zy8i
yjTjvt0nT3ry1/kh/yvD8O4DLt6/yocCMFeexk8uj51IzbH4HZhbfRArkWO/t0T8
A4hQ/yc/BE9dxaLr/hbyMhFNQCo7lPxQqq3Oeqepdv1BV1rp8YOPGi0Vy/gMBGLV
cHMtkga2fg3pJbDxEDoI00S/t3qMQTl4mMeE4+DhEmg+tu2nNAcB+57GyO4hDcnR
P+z+Ox1rNW+yMyr/fIQVKUr7f8ez66CvobZW015hvGyqCck7Ol1uj3eHmgz0org+
5lzqcuoIgfoBtwVp0V9tmsCuYVXdZ2dJLBgoWJyrmxwbcZjqxJyh3A0KXGP1CTzl
mQdhpf3jSNbhvZNRr2REKa5g+qxr+Y0Hw3Gl1x2wPnCfCG94ZRKK6xgnSnv0zug8
laxrUjEIYYEf+Y2fJNG0bOGzFOF0L/qLvs5LT/wIFtLp0CBBvcnQMR39EudUZp8J
Je2rIrVGpIlUhUO1yuY8Ouot9oYyb94d8wgWYRNlYcZDpHHO4LlRLZpKIdVZpuMe
VT1z5v3zEY3jZwzP3OBF6V4p0F17fn/pyYXKWShHAolbYFtSUL9OhogF6YevN962
bpF6eRAdLmzdcwPST3uYMkQGQgqr3PsPDZG/z27+KdQ8eWolXLQkhPOBdt03BHp5
mPNX1U4jIO8wECSZEXkKF0F4tgvSV/qRTJi6HB8gho5Vb85qk4xCkG8cX6JJvtON
utSR3bdwoksuDmQLAZBRhDDF6a5TsovrACd/tg+7BaAHg7vMgQyEFYz091Aa4IZ3
D5XPgD1FzSbsPz+6+BZvKjyfWVCtctjBLYRmYfyy3VgNJkZReAaBoYgtyQ4r+QeJ
FreeokUoHB6JvlypsM48A1uRz2kMxtvPAV452rHUs9DxzejF6/H5VjiZ2WZ1utKd
9NcfJp7JH+WOYz/yxD8oofCTOYbR6sLsq7r/S7+GF7xyurOofijclM1JatBU3LjB
TUbkuwL+2u+WFxm00Gb+Tcl2Q0H77Ozg51Ze907j3rndbjYGR9wUd4ZzoSQF0gMP
kLfkQhKomc0z/zJV1lJrQ/dHN1e9tBatYdVBMw5izlj1FdlYsw2cs7VRdX4fcnhe
HtbJkdO4r9BMu/FtlkAaW7Vfrly9H09hDaIcrUbaf47jhdQGQ8ATXJgLwKoZt9pG
od7W0+EU1s4GJUl/8uT9Tv5pVW1ninecBUR6N71nRrwlUSy0dRt+BXupWdSqeiO2
bhyHAinqT+1j+OzO5vPAjsJc5N9JeVQWB7s7Sp0S2f2Z1NAxTiKQpIjV8cGGypQD
n/yar91Al75y+Ytk5gwvHJI4bQWRdD7+xmVWyRnellgf5bZIIiIUZZKZfUBFW8ay
mNOZaDv6fGv+9HB+JT2cHmvp2npEwlbBbbRtSoOtK2H/Obv0IPpoxy6iiiSxznvu
XtjUxwjw9kABqX58XR2W8msC1GeXBZ6U1ND2F788Pfnd02HGBLVa/rAAewcaunz4
91iAFv61R+EBVg/zh1e4/AhwIThuZjg9PAK3GCoHQa23T3T9POdD/Gn+BngXXlhs
pFD1kFX603guAwGkFLLPsZ3YbFeblKK5vqhYo7QP1E9gRIdjUNyTKd9iwpxx6ToT
pOPmgiM63UyuqHwAhfaRyVpR9/Jmyqfn/MO/QUPU/5QB1RI7Lo/s0fKKf+S6Vwxl
3mial+Wkut+phlqARCIRnz76QKIvNfTIBopHtSJJJPllLwYV/bPjpgTy1+cNzYS/
S0MCAxtPUvWpfrI6ziCkYo+r9TGbEbMrhHlFbHqluWB2lroHvHVdcQTyDJC3gOqO
REVeRiwr9Fv4N+TR0Sdkp3KLHIT16J9NNIAKxX/Icw286Ver6e/ElHM/hgHNUEg7
Oby08xe2jaeI4lj6jPOROwv33mC3b3gNaoaM+YDz1wsRgiI1syp173vpfMHCEk4T
C3lS5uoMuZY61t1X09/w/RyZWUXSlaBibEPcRS/ZoOEJMbt+0tdIHLmH5NCchT1S
NlsvxxunK8iXUkyGHJ7pbJUazu74+OV7a7Gnunk042ZcOkwbFJgx/iUanrxM3dcz
B5kWeygrpp3vWkj6EK43xmTdvmpa+b+6Pk7NYti5Ah5j8U/BHPQqk8XApa+rY8Wc
DpN5ubZUtngkWrn7KfnZ00Ez4QHn06ERvzdhkBjA2KL0kgHpKP7e0V+MjBASlWG1
rrSXSR13WMjSTXVt5VPGcPYUakPt78+a4x0eBLIekW588WE5ufiV2I9LICJ8B54h
mRFRSBHT8bYpJ7UFm5hYaI8vMpF1Bdo4l/m4w4Mv7zN8i1bgjZ6WswNSVVoU7GMt
Udvu4HHN+v8QakFX1ovV+hTzoQTraqDq3YRtDYuPYTFTcxMagXn+Vzy6q7sOyWxk
y/Gl2Cr7pWEhgfo9Z98YqKzp8PnFIMblcyMeGMqXIzSdBwk4k3hfaudz4ykInBE5
kmeAaOmqdWpmFPdVeam/0Z7rrnQB2Fr0MYXyLPkOP5Z1e1kS8iKyG2ebmp0UqEzB
wD3aU5Rtx6drGRnh8SAvAZfb5LcVcFE42Xzl64vZ2aB14vdtLdzSBYr7PZwWf6T5
w5tSvWJmoUl5T7JL/bmTZG8UO6gywVdbyAqROn/BNRwFRAcNGDfXnDKN4sVelVhK
7DzZ0CV3Lqrx2kiiU19uKtcXZuPty0eDwToZKBGWYJWUyOKInDvvrFkxldQhEwlU
u88mbtlUqjirWCFMbokdfxwn1CqPhWBCdJO48A1z7RTT96duE8mBAItFFDF7Ck69
TgS06/MGs/P5ogEVuwEe63m/Sh+0GNVfajjbxsCz4rpKmcmxLmC9oOkDOeB0LLt6
yq/pydqP1/t+XUPXf0T2GDjboN8ZRyDkorqrXBOym3jjsY9VP8k5u94I0rbI1G9i
kfA3FPa4kfJfPf7RAlr9dVL10kfLM79Hy+bp0rdH28HG0e5W8Hn2xdO4RtbbUyL1
vLfRvIUpcB1tv7vG3zvYCuf0T6erKxWsQRIzQ6nNcyOROJ7Mtntj7Z84wMA8G1Be
Rd7WSTm6QyVccAEFeX4hHVcSn5tzY+VkaqmRuaGnXnurlARVordntU1ImCHelL58
eZNmUxVrHTh3oiqCjXszJjRHp7mEDYdfR939egpBFMmdgo3ZyMtr2LmbLUNoFFeu
6acGgG7AQ+40sx3sQOwbqu7eBhsdQ4FB5xSRglzhLRdy7rh9A9peBBvZ08eycjV2
kLtNu9TaLAcBdZbAf+Ovg9t7h73fTrZy6ELfoli6lyOrnrN3y1fxAwX7Y8cKbPCv
epnnUBBmR/hZXjaQUGleXuiQl5DcjkNVLwbg2LQzNG8ayZZxguHxXh3xTAZBoh5O
nRnb1E37RBjT7V0BDjzak3EwZ1f5I1tVzSKmM7juZXytNJttEMd5X2kB2s2KHkUB
7dXKgq3Jftr9KR4QHerQXFV0I/rYG2MmgFaQaYZMLt3f8s4coDgUfkjlJNeIjojr
sZKWHQO+GmM0B4eFN1dOwH2PtmpQ06efSnJ586mbd4Um8yJevHwE2YUAmHK4Cxp1
ajlJjsVOqoAOlTxAoM22YJiMY/CBvq+Tt1hlPLfeWvIF0yf+iztxsEI++YTX+7Zp
XoTaKiN9JghUJjUXUl+TZXO3aTxzSWXSPEQZ/JgPdeDDRl3cdLsKoGCqGWzTZGMk
WdcnayBGM5v62cPaKFfEmZbPRgPgugbFIdtkT/hhNyyaeG+QLKWuw/fG9Y4y2fON
XL3WbLynw8cNvarYsAQXp3ttCm94J+SgjpQc9mg0yCc0xIGayyp/tnPNwMpevKOz
QPX6hd82BdBzKnVkNOK6zGv10/kMHOZAkE3Al7bjATMt9jpWPwzGOShvixTf9zdI
l1pZwid9JSOrzEVkUZcOB9daeDnnCrBWTZCk8yAD4UctZfokTETiGSe8FAH44ziQ
qMHUP8sq1BdoFN3sHQ7MriXTf48uYEd9TEV25S4QjT3R84+4WC0dHf5X5TYxzFyY
5DP8J0h1ToyHtf5mp8CzJjMY2OQ/+eTOAlnNqLo9pLJYQeN5GNsoFbzLKzw2nBmv
N6fQyWa6Vb9tGrGgYGP1vRP1GGsyO51bGcbHRQjuf3EjhzbBl3Q3yetFFz6hzGFH
dvFem01iBFrNP6Zwo3LY3Ccn+2ZF83N9LnyHe7aNQMJL+TY3Hyw6azkZYGhhU24F
BRVKDI7m7nAsLRwHr5so8Kf8idaZfLtOz3ghsrUQdY0l62pRSR00coK9jg0KDRdS
ekgZOrR6dBbmWoEHSSwtL1tfo01kW6CjZ4+wCaduh8REd7JrY1hp8mwSOeyHCBid
8Dgu2nqXv9uqonlmFO4Xu9rnUH4YHTqDIBTzrqOXwCf9EvHUoDHFgxVUBTPfTZYh
2rPSR0htzECwKPV90ZZd0xBuOizFbb7ddE9rsHuAOe4W9ijBK6Iqpj6HIIgE3HPv
6b1qDGq1W52BlfqOO3SrqiHrMetCmIG2eAkHrzl/voKbPdcXRL9zc97fJDyW1ElR
RZOvN3R4OJwsh16uzEDjWPbhiiunmV20wBEOBgkfArjX6o1e4JMEYNgwcr5DAcOJ
XpKk0Mr7bBWszgQr7ICR7TLgynfLtkxZ8xHYoINuyyMJR3JW7TYqIXkmX0X3+ZV1
9BFjzuNqzgQibWJIS3N0N2YjxsnQJTV7+kwpEtm3GfPSMekGQVyD71HeSpq+48i4
rtL4FmDd5rIOnkVlFKczcP2S5hvVU4w7eW28GbzIzzt8/vow6cvYMKw+WKzUxlZs
NAadVl3lMD9DZZKyw3JxT5DlnNqK3ht9RgdAcnjXbyIwVMy4DH/uXtvfeec0Jrub
h3RZ4E3Hd/d2+n8sibnnB+XrsscyNLLM/sYI/1f3/Cy1BhV64OIe11bSoeej1n9j
JjOz+/9e5VJ2jRHqGeGTE1Y8in0KW+jeCk3l7h+GGbg4TNnrT2qkEx2U8ukpPvDQ
O/QnLoSsgsVcJEXQwzVi+jHu9z7rQc+rbsxvYuFJIoQ46Tcbt4qMZmRNzImwmiw/
UYRjXOfzFlQuwVaipJvLQ7KjH4aE/eKOumpV4PPW4FdDIXFQvRFmFvi+/D/kUuSq
fZMA5szHkxBgIfuExAUx6carIvWe0k+QObaABl65l52+zxZ23ioKzoJ5kqAdAGfV
5HODfpz8Ma7cdAUZ8mLyCy9vlXW2+W5E28gNlsqI01RAVjkHqSjhlbem8b0qt/U2
UVxyp1dmulHvoCZV0UcCwWRKBdlMkj04Gmf8dXNaGv+28COqTnPF290tT0KrMv9B
Nxt9UiZiBzmohftAF2AJKXDxxbYx1CfyFRWbdvqW5QLN2dCey21ZmpBXmT+GFOkt
xsAdVkeaavs+ohfZzX/1wmKWi0qQM4SGnaxM0oZ/0Ubkjx1vT8bO3JqR71AuSCSV
Tya51hZC/JhnoCSoHRWZadixwoNVwpJOxVnIvic+wQzjMnG844yvn98IwljBBJzs
NTmdvF0xh8smIpOnhMwDBL+/jrwho22WYWdi8uP7iFYgASKVgw+G8a7ZLAkallmt
2gARPeXXc82+PSUPlJyblnpv/lN/MVmEWd4GzTimTTi8BAcM3jd8rqh0KZ2FEFHR
h+MEPLn827EGfoWQpY5Rd+HRKV1PxIgwwUm/dmThmXFmHDiTzFXyaNiJPB3yN4tM
Slv6owwbUdcKXy8RCOaca05E9DzZVDWfC5QyqSdsaGEsJWTbKm1ah24ZhhlMge/V
9pzHWZK/zoR5nvDO+uKXu341epvZ5iyYaO0J5lfu7hX79hIJLNXoRSLoqk2AgWHi
gaUdgxqyMcFN+88GXnIUII/37tlS43QPHbzt8Fooj9VCzDRLHPzS3dvlGcdaQw/i
ZDlopCQeNW0+MrT64FiCIZoSdFmw3XXkXA27kea+lWMP7ocAavA/SZ7N/rcBaOA+
GuLlrfNSFFd5mDmEUwWCv3LuhMqj6Nmb6gmvcX/Qim77sMJXv3IOE5ZvO3NEBbqf
rDBQsWarQMxWzv/F4eh8GbGMHVncDM18kxH0Np6QmJL81cTxZ+iPUvn4T5kX0t+G
MAx5kdSgrxE1dUGR2o02zymulA1RHFu/KWtXCebNQ9a1dYWupZhX4IZYd3MIe/Ev
gZ69X0aTYndOzPEHpX/ND4gXAapjT9l4Bpiov6obriaDoa7Hm7/6i5bMsYBGdnp0
E3lMhihsw1EZjlPnujGReex8v9XDjUbwC/1eqvTX2Bj9vbUPUWQzz8j2wxHknReE
e6lw7Vy0417g9NL3SB5DzqQ2MIfkLe3MCSVrTkLm/ZHXAZD8f/8HqhSRnP01aKQh
omLqbGFBSrAsyBwJfq7p+zpp6zFes/ZFv1PFbf04WSwQguJ/1+ySaMGO2XvCpAhk
/x+pXvSLZ15qAuuqSwUswZjLIL72I/5y4+wzxCrmmO3sQflXe1ONZ2n9fgRZc6JF
Fkuyk79BgPaL2Mk2OSvT/FBrCfESWvdKYciPdGQOK9PiO/R8rD/+DawGvc9v7Hu3
Twz58XyVTvZA/YZkEX48BjctCR7pxPlYx+pTfdYlXGRXVJ6kuXmKkeFEQIfLd9vQ
KM1Z2CTOxUan+ACaFrGuR16/ZA8sZqmpuEgOPq9v2/D/S+l6sqeVGPKOgI+41m2e
5dSK0SiTqPwj0109WKVnDENqAmZoIfdkTL8LmU1H1YIWLbNgsZ1s2JUmVQBBSNcc
e09wDr2fZ0LQni01bwQpS/UpNb8xscpuCj2sY389x8npU7o9dJ6RtrnZgxxtfnYx
yDluQukRJjH79z1npsiUSPWHlkI8OiK5+dilAOlTA9vxVpAqCT65oueheurulHnU
9zGp5ve1YvCrmST836acPDWpN73gDXABwx31RPaTfkj9ThBwUHp78Jn9foEJu+LU
Tp54kCdG1Q8y3AGjnO+wD6II4h3vPFRgo5JvLhqOyswBi5RFFeFH5Uhw6PAPUcqe
hESychbzljJk1xvTriqutOPSG8E51a2vHP/+0n41ugPRjdHydSTXLbqqru4B/bck
Ytk3kUJy0Z1MkYOba13T76qiRzsMA3CvNyepgg/ElYWP7ld86q31CBXblcFVnpQr
GCIVxF3WBC7nLB0IrLWqAnmOZ5y/mJO4R043Ql/nJlCzwIJY7lP8lOdhbVJZPKjs
jmU1PJnOD6BpNPlmXIEihyqF0iaviQ2gWDY6v5KIAcbeHFJLralBdSLMxuCobnlp
E2q12z0iNQalyNa3cRNdabW4vjgcE0rSvhd4/iN91ZiccsRHW7qWY6DrHRSAZ0NY
y5pnUtLFyKChbttj4Ha6Bi+vB70vyaXBkKo5K1LUksNlLTS4MD4J5DbMGl8XjnWF
wRtBOaeqZi5aghvq10dE9SdTyv52MhnMEaTsTERxYT8RQUIC5SyKNFVpKswPgEMl
PwVzWby+qYLA+o/UxkE/DHiNFfApRiMWlSANe9KY9Dpjev5+euY0Ow8t4HpFejyd
NENnC7AwVHS/EunhAxXQM9lEa6PYPPLf9Yjc+7aHQI7Z6pEcAHm/l/ny1P3UkRlV
R/NMnV3ktasL4+ylzg2ZnIbuMpvJaSwJMyFx/zAZ2nlKcc16U1pHHOEYHx8eUx3M
6StZBjPLMlG2p+2ijKB8XP31hasBxGegOM8EpfZ6f5jUK3v7rL2pFwzHQvHYH8r8
1o5eyk72Agzz7NUaY/vU1iMdA69HoGJqwMtNXxbO1xZ9jO3p0jNVo7EpfOVefDI/
t6woBp2ezyp+xrULqfNjjEFVBRq3F+oCaJrmfhr/ZbHseRJgay7W1PpL3bo5QhR1
17c1IdthGihRZCk8l5OmFzvbtxkK9r5soQRtsXabLQb6ctcZmjArJqhNo0UInQNQ
cLEsdxRHpLVObcFATCLuNp0Mop3JCKlhPwcDcvgxtriGl0y1rWiWMBCoG+whQpV7
25fDnxBwSwig4/g0IDObKQrxwh/MSu5SmXRZMbOvrRZzSFDsILWC2CUtdErEir3i
a7ygNHWJBQS4FidpcUZtxdpmkmtFtd8daqBMnOc6M5wLgnNwMWyek4/wu9lGBArL
u9JXY9g3z/UQoZnNxLE7cf3YlwR6kPFH7x7UugBJeTPeGXOzeQZMyVCMWCTZOrQZ
A0+rIuDNIKPcHTjI7r9la+RESS+OA135C7uHyY3hDJ5S3kPMGeNhv9zyUj/JK06U
3LY/HWrfLcuiojXzSDspzScD3kPdYbEi6+e+upcjxCQZRghEOKoKV5lsvPBWYJnJ
lnZUDWIHFa08umcVRT8IfZW13jWmdCBsQdbedakQl8TFpg8CuXjImJHnXPBXyGvl
WS0C95iVfq0csqL3+SSDA6Av6ua7t1QV/RDhigRHFbFdxEDFhAPf7D8g25B7TpYH
Zp9eqPfE7lhkt/Rx8wSgI8GxklF19Kc9n4yPq9DM5rd9dENqyE3BwsGZUz52Vdx5
RFyVImDsZ5GkpaDRCPc2oSHmk5XW4bQNu2u3kwTiMoVZn3J88ITFZOrRIicTft0p
BknXDs0fz+0Ye7nbQsW13BDuvYqnvHaixipgBWGZBpimweNHDq94rYmCWlyOg/y4
g9V6nGRg7zumnH8B8st7UTovswVFhB1ZNvLQudoFvckQAMmeTQFyEcyGRasFuezD
mOms3k9reOKXVskfs5cAW3Rdhk11eX6oJFur35cE7kzNo2hvlX44hQyPmwlkUeGz
lfCW4CcAIjMHGWEmuKhH4NlSfKZtLbcVkLqqJTzUznc7KLj67M1KbftdZLRTObrA
Qvvn/t5vwlbfmEPovHLEn3ukeEZIVjaMn9nQ6Ha8rmda8M5q/zdluvhf+YhgvFut
MGOFv+ykQ1rUAOlcYvckrsaffyDyhn1gPskMlMSQpmn7IH2ch1WsWTTT/Yp7Z+3B
7PHYC8aIfCqydgzDnEp8FHyH2DkOEpdAmouFsE1rQ6zpM1Nu9zZgKWRbZN42g01A
WsRXGLneAuKK5uku8wskxzaMSKLf9XZKHoEjvt7CVIwD+6Boq5o6yabhQWISoYc8
WuGEVzJVoeyypT8hshfwx0dcwWU/wsIvQKg5Rwup6WR8FjaS309ERqpfjuIahYpX
8EEq6juBXRJke7TJxlGFR2T7wKUdzKMOkrPs609ojRUMakGKwFiB6h0I8JbCYMwz
DDwtS4cx6PYVOLAg/u7K6GtpJN1c+CmrNKHs8siwUSGTlIHzQwRWXZUph56tuTk9
WSSD1dhWBMoS0rOxh8hHv1meugFHgr2tw2HWjw760tkigxwYPOICMnRAqf1YN42+
DCjU+8m0O1jVK6/O92u6LV/tuoF+MZ+mjBX/M4zV3mBWL0SxpRyxTAkDgekeT7Io
VA1X0tJj7X1t0MEkJLgvkurRH6eQSJ4AzJhzTTInAEwUVR92WJ9faNH0kuM88Dk6
4rx1lFfl7I/UvoJ5QcZfkM1GWk/IlpdgMg6ATOKz8itUrV2TlON0IJmBmnlYCIuc
SmPK98s+3Ul9CjF7QqjreEZ0v6ygiJMkX+ZxxKNpjLabYR0OmDxDS2FX/AIoPpqs
yl8g74NDTdz+fSfa0GBbmHPWoJ1peLy/nQrudQtCcTBaD3fuy2zHoAM7YoYlHEUv
2js5G+9kRN8Zs7k/RdCMotRfShjoKYYYxg9tyovPaXxFD+A0NMJsDbxUkRODyMUG
JZ598AbHBJt7Hj5IAKsvX1bGSW9Ci/+K2+gB786jOLMPATrD6XCGU7YFf5WwHOQL
wW+WHxOmsHI2hShh49ufe4vkim4kQw3AjNc7kdoTal18THGLJNIztjAIULBlmLdK
1NMG0MqX7QiiKAhVUvHuYWjjJgVBgMQnQZZK5yZ0oLf+JqzDMS31z//lu0BWjUm8
czJ/Dpkxb0VcksXLAAiMuqB9xsJd8CzTlVxxLpF7Zxf88DKzJJrTBVIqfb5rF6pr
GnRY3TUvXXYy+CbXeRvfrPJ4umT1cGNKML7lBD4wFBXxIGQnArh+8hedwBod16S2
9kj8ldxICJrDNkMz+k15o3o44pZ+kfwnXEALxaVCM8VJy49MlvopRBeemGxbvtWs
Ep6P4I+MRP/KINK7/JxDmK7S+fCDgCgTfjnrUhQVF22YId98BxnxtOQ8CQAFuP3A
ErmHf8EOMrrE8JrSH+HvU96frtnx1k4poRNhERfAfQDAAvhum8ZVUY1anbZ5PdCF
LfReRz9g88YWe0q9k3v2h4jf7PkqHA+Iq9cJGeSvZpBuXa65hUfGzuUpXrhgOxqC
yv86236QTi2uK6zvj6DWvB1U7fzmaQFEdyobaWk9kcw2PLXyLAwVIwY/q6siEzBa
ymn4806suSNYDt5zKwLd1mIpRLTSiik1Dn0BNoi3EqlkXgqcypvejw1idMCuhMWv
8n0x4VoCImlDIHm1j0tyGyc5Q2CBdofSfMBjW88sYw+ZFr2mpTDmvOAzkCuOyuNb
0dN9O0ynxoFj+TlWzm3en0bHfnEw/0ftFJ6xqDg/GKpJ/+KGcQ0wwH/qsRYT+gnf
QSKpJGH/Xqf0C1N87xnnqzqonCkgolH25Q9r9+BdnNRAPBNxP4yzY9bJ52nIiWM+
7DEtwBgSS/qLdPShUXOowuPHGvC3D8Vtbdc0iehesPp1OkhBmcvOI6/6gXpkejwu
sawOkxLAhqALPuMG/ilnywove0D8/tnhMXMyaJcikyynSa4obelptvnhc5EWekpa
pYiv37H45UYrH/BUL7uD3F2twOs6lTt/og8Cxwf7aR8+QOm1CdI/qGTGhwjO+Acm
0/EyM+LNqMo5cdT1L9dvYEnadt/0jwJsZOeUtiuETk4wQveMGwUR59M7CI5gkYrV
9gS3q3scKXXnX3jXbxMPm/r3q8JjkRRvS4UkbyJnnWVCa+YM2xvm4iTIuUvlHWpc
cr0meoMS8l8HoJOAgaBt769AxWLG3AOgglNAlFy/GayIhOodm0tCz7smQE89sz7V
FX1lhL4TSaw6aWHMmfh/EhVlUvjb1N2/rHEpyjpxHRHPVRCXCFG4F4CMe0S34nm9
Ewv/A7uPHzxHC95skMgT7e2pJhkfW50cuMpOuSfsv5EA55LiZOmfbC0dxxb9y1cd
QfxkEQsXbknYRM927YhYkxDOMOUetOFdspWaEb2mW7DmXSccj6Wei2Z+q21aE/c+
zRtOQRiKzEiX/QK3aWjJzO2XNqSQ6HtVACrWEG4yoEyQnJQnSvjEoeM0MR/HgyDR
Zmgmvs1yL30tOrsPgVGwsDHGLqcsroVChTJixeu26EuZTPkGEUAP/J/BlUDUCy+F
WBEds0ost5Sso9Jwvsl7YicDPduQnHz1Q9Jhbc1vtqRNqt29MplJFKzpuM34KVt1
CW17A2SiipOyTX1zDNs2BH66SuBH1e2SUHHmRzWzRk4tT7ePYwJOSUD+TVi88ibI
ER4b4T51xl3Jz697ABsQiPjcIqiN+LLEDkKWGHC5Kze/2Zh46iw9Icr1O22AVv91
8wBZeaNgkLWqYSY5bKINVogTS+LVY+NPNnZU1m5l8aC5P9TUXjXkmwUaV+yRQUpR
6OJi6EilDfp+CssmuFPnkXPPIYmFuQ7L0meO5D7TJIdJ/wzsAXYA8U2o0cf/1eaq
cRtBgaxLUkw0JPt8AE9w30fz2m1gPBdw6HJHc90kJ78EN0gtGqWVIH+wyyAvd61e
tNXNZ/71IqhMPYgEu3/ovXmLNEuTgpknqf1btoZa89MwBqO6Uucj8h2CQo4mZJUC
7K5gtcEhxwgoJLydHqa9BvrfL57eY5niHsmD+PE3NVF6Dede0Izp12WQ19VwgfRS
m+mYW0xYh4oCbNkwGtrnp+J28mqrqI6bUW+1nlf+1ZzYdEDOZgh9tR9es4BMYc7g
eIKQvT41yMLoyvehRGPoSRuH7o/GGVHSXMrBBl2yNOki6PyX92CICnGbMvJcWtHN
7dwkTPDHMYL5RSkhDDvH+ozrcpU3m4A/S0kTf0ngW5fFWXxNyCD2nLsqNQzZbaB9
QILpyMUAhcmnwmxX8hWKiruNFhmnlyKnGcgFMEqS1eprdQXde1kEYYNaQXikwfLF
1kch84UFZlNoqBr5P5II8uKkynH/hLntrqFsLur7gAWaKpLyixIZMBWTypGp4KhA
SPl+vN2CQoX6L6oYKJaHk5rp21KA2XU74O1Lxy9hshDzxNBoypx5vqr9FwSpmky5
LuKtMKJcVjlTOCD4yMP+tqIspx5/JfEItNhAEEpzVkH/y0kL9YPiW1+9HWJQHaK3
hxlDM5dyLAm3Wc970f3+x2tdFNRwBt2E0vaypHJ34ks76v2dW47WtWRHkf2i8Xrv
6nTM+I/NqO5qk8IKb6eAaIJAgXry5zmo8IBtVZXXp+9tBcBKAFUJlnXYR2R+HmCf
ZoFz3UDXRXx922CP8HKbGvmxsHNl3SihoqkRDqCAw67IngWDLMFhyOs+tFEaCBoR
Hw6Oaf9ITYajqaOW88oZM9Gq2C/zxq5ObiJQOQeE78xfAnG9czU8dbhhd3Gz+oWR
o6VFtT6XnSxJ1OCGYuwcofDeMEMXf/kelmdEjCU7FNsX5I6HOsnweKXOISJfp080
4jE8rgATTL3t4I4/cdqTR++yuAS099LBJEydV59K6654U+YTBxWf8XZ8wyFuu3pr
aNChFlrudhN9EJNUpEEVceiApq12zMH19XyxPDZA6eMis+Can/4ZhjFWXTTLPhnG
S4aadrtnEig4BbiMn1W2UeT07uB8UN2t60T/mVGCb+XPMiWicNpGKxpgp5we7n9R
hk/1kZdM3XEk/mSofwYueziJcCbf1WheX/ZJsRHfeXC1NqwaPppHqWwuEDkU48hI
O5BVj4oFFuj1br8qcGKoRdDk5nV8h8nYxzWOjgRmS/H3SuajkATLCxaBjUb9/eaI
Rd1mw8JgPXMX4cbtXdyg8gyLJqVNljIdeY8vcJRFrOVcr2YSxDP1GwLvWuYaGShU
WfdRBF1lMw+VA40RsbN0k6s+y9RTzRoBJfqTkB25fKlvAG33s0uaIJh+GYhDnb0N
H/3Dadxzn5SO6gVDBUPsBh6a4Yt3EZdk0bUpEMClEsgJuxX8e4knVLYvtrzyrN9a
MqYVqMOdICLkfs1V3RzYjybnrcbsbF5b2pVtYDpM8lIUiMGX8CmXtCwHnmkxTLrq
t/mhH/JlEOsIaCeDKHKex5S1CM8idsmp27nV6uHM2aT7X8HEt2Skdh0l1w5km1Yh
jGvgYoqzQ7jCosbjA/NloD2WfCfq7D1RaFsKkFa+xq92zR24ge+H5Y8cXwN2zCG6
jyru4SOa9nTfZnnvrIxsA2hbaMEcFNhVfOPFsbi0M4zg8SjKOlmrBFNVCtvNLixX
XfQetUR/TirVyA8Ig851C0e2ZP32+2e5S35MXVe46qQEvx3y24B5WB41ekw7cpK9
sgIGY64yUqePHfGoPHxwoB9X5R5/RytErbiUxcoZr/6J1Frfj9u8ee/OyywibiSL
1w1wjOgNxLF//q0SNcSqp0qHdxUxjzikctQtz4QX5jm/spSAt3wEo+BBUYAj232+
PKJKVntjIHKmxARmFnxNeeYdWxQNdhRHyTrS3b0eF96dVqqvE8uKsCZjkZgJNoaj
1B6EQqwoeZkZc70LIXZHxyQAtlNlCqFy3HLX/X2PCVClPm2d8bfkWdB1OzoiWdpq
cSz9vYzG+qukh9ggOJIYkfphDsoz+QqnnqPCC7k+whltL1ew8nqJXcmv21KUzM+L
oh6cN7k/ezXBohhfPuQj1YMQxAfq9w5bDuEnRB5a58fAfAmAX3WYi6bKj563/9P6
cmr/9epjE8fOMlLTBIKOgZW0Kg5ftxUF+JI62o5Mcy7+H0xaACMySgxqV4a2Gjsi
3Kkon5xXP9YJrUGbnCLo7TzqrJgDE8eF+RgOn2gUWBYIk7Eptyfp/w5V2r+JmeI6
3WyLvOqHY53yTdKSBlG2pv2VRyf1pjzcOnFfJjFxNRjSw/NlghMql4CDDGRNEnmL
kU8wdMFmdstZWxznEFsPMBI2YXHRhWcn0L1nYYi0CXIVOBtcEHItfiEFM+6L2lNT
DZqUOMCpYS8PW1LsG0+t9Gf17WjJvmIK3GD0vHpnT4cCftJt7WS6HjUHZ8jveQCt
VsaABTUGmm9wGAWOb9Vfy98IubhVjRlm/N/b2Rc/cxhEK5a5H3Btp2cxTbyczyw4
2AUlv7Nu2pMIhPgt8Y/nnNx2PcUJojNespHtgBKxQ1+ux9hxEffFvDO40esNF9lH
cOJrKj7HpyAt9z8HwFLygR3MSpFt2ELqqt+B/Y9gc3cDM0Hu/oifvv05Xpl/c+r8
YmGYsa7oDCvRriqIyXpJ2nfk+R68Z4enEgPe5i1I9KWGctW6CMRfACY4G1KMjyMl
own2S68E+iD2+aRVCcrQSaIxq6Ixk7sW873Mqpy77XGwGqqtKBpCWEI4qFiSvEqB
7jRc6ntvGxyGFv8212VkRYDHzNM+RWJcG4a7wYpPFt5Xr1dDXSm1XQKAiQHJobCT
7XFisjhRuu5jdQ+kVkEvycV36iwAozP7wB3Vrm0+aOvx0YRcyIPHOGNDou9GgdI4
O5gatu47f+aLGU8zax8GtQ+iubWUqa8nTZP9H0ZHkb/zP4wFI5V3FFZtkjHFReVX
0fDVLBdjSNUQEv6Ow4oSEvHdFLxz4/XsPdG5kUQqaFEe7SSH93u/YHDqSG6UTA8R
8giDj2Cq/0dtyWnLCB5h/OHFrMEh6zZM+wYONhcuSDBVKKVeKdep4u8+H2Pmpa5O
3aehziA0WoL+rSgBb9zTF/etZbdt/sv9LkgtdKEqq9s6ZBzhAr35Xqs8uOIFqMJL
JeB26NNq+QWAGdWVAX2TyTiGVkfFzA1IPIEWOXuZbC2f7C2zFZLclH7aCcFS4X4d
mnx78GeWv6XLANj5lk6ve1zP1Phxl8qpnFyP5CXe8iF5Bm+3QOwt44R5NoI4g4ue
lRVpnKIrodXEyJ1e/By0wRLL8eq0zo1bMDS/fXE03v2HSEB4ZYkfMDXm2d6gciow
soydlG9012hnQpeokY0AR9CJM5HT/vXG8qUFPFMl04b2dqsHdYmVIXc9l/nn3rGK
9cQWu3lBGDgWnm0xerjufS6TjcZhEiq89FdNRo5jeRWpST3RozHJyWd7s5IYVtUO
p1Dpkn2NwTq5P2aamQjNl5qi66q3Ib8H76OUFmFz7LWFVWZo5fQSCWIPQnT2ql6e
ShcAd7n4fgryOgIezEdzzmSG2RMuQayHmTcBT1x23TV1V6RtJkxNHjlx+UEvKtAx
QgZQwDx3kfLigXCLG9GhDH0toDtKUd/Fjb1IWsRnRVNsp9amDAnDcB5SkbeDulJ2
QaozujqUhtRVQf/qXbfw5nDy/Mk2kNIFr5h27Q4goZgV42aUXG2F9PmhxcZp2FMM
ZUZIc1unOvPXMFgGP8ifJuqFah+4CXlvrb2OYmjcVIIDvZ7oDzfTyjT2JWPbBC/h
XvK5pouVRxdM3OjdKBrmukc/s+SJVbjpjTIBXGQ046jCWpwSEFiCBm3+vuDdfoBd
3PGinhxLKbNqWb3nQbnu2lqewLYt2YftOAdCEx7ApTvQky7PX8DtqRnlzLdfjGEQ
Zj93SJXQ0fKw4xeVniADsbIDfyt/T68L7I9Mj7eSgsmm/50+I5JYrJ/QlXpSt2Yq
UEn+2nr2HMH78WcA5hkBOhSwb24MlChEwewn8DJEw2/c5ZmMK617yHjw87q4IjlH
3nZFd+dI+ap58Mv8EXjCLPjeSeU1eIYC9E9hwMViCDM+clLPXVi/OHm/ajmNP4H1
DlB0jD8U8GpzzzjZzS/TcUD5C5y+hnuvHHBYncJ1zSLvPXTV6mpHxqfGYAVKZ7sX
Mnn0wzolIdQGbPQUf+gbix7pYQFIQWjU/wxsFgqisoq8VIpL0YE0M6qINz9IogUN
deVj0sqnMNisPVsZttiHXcQMXAZMboWY7eGb/YYvwSb2CXl2qiOChDpIlZOCyN3J
6FZ9CyK3XHnKsCjTUz5cOmUTKA+Df/JROrmztZxD55sW1Zpn8FmlBx3+bxS6HIhF
+17akXfoE328dbRRDqzfqfpO+fS8wcvuC3LQNFyOaOvsgFnO2J+VxKrl/yETEosJ
Nu1nRnx7LOlHiO/UyPLs+mevFiCEOrNMwG40CkE6Z8UsCPvnGKNPc7oKgcMb/yeI
MNKi/CE85w0Z1G9zmeA0qNwAIPlhHnQo2epLBj7/tgyfapT13JcTK0bnHEyF4AIK
tZKzA6m9Pw6exyXYbcpre0GIRLkshCdx3P/89V9RnEtlpwREnYFP7wVG/+us+CHw
42KOwwhPzuDt2SQLnU9L0VXamPnCBNun/uaZxLI6Xrp5TvF0IcG9Y2PCLF7ozpHU
nMRb/OhF9nFGLFnyKfbwVRXTJjUM+lAcJlvHPcg7pOvj4AGGbc9hMkvg+GrZowXQ
yRFxfZIx685wwTLUOx54E9oZ6OwV0uyLr4AK+FqtfWIOuKYI41howCEUtmEI/9Kz
x4mGhCFI9P+4u0612bjPCjQfJUKbSXLxr/QHi0PSj/Z6odtXUGFrO62jPPaLrV//
VLETQfe18mWgV1QHf0ysJP6JRJKLHhhk/IVr1iePpgoc49FlVfbsvaf/1Myg3abv
DzahcNx/FztAos7A5NgEsyxzxXE3c2rPyrjP5CY32FRN7C3wpF0cHI44M+BgajGp
J3urk72uYe9IWR3HChF0GP0AlsnDEjJKL4Mb7ee1DXgUR7ZY+TsvTo2dqWnITjNL
or55XJwdfOsAu51OeIP1rZm/ZKe1iRZ62eiFXtSC2NWSLZ1Qd4WnFpbiFvg+YU0G
hX2qaQctXQK2KjMEd+F2UMMIE3xtiIxt36K9NZ6r0FfiJu/JpiEX8b8gvS6166DB
YY7mdk+72XxenFlfnIbcsSS5KnytwIWuBrNDJRqU0oH5KWVYUZKH03h89bAjy4gP
1CzBQilpY0B9RTjRObQH0mOrErrkhq1zQv2IA3uKGhOltfggjNRMHVzTJi5OWJmD
zQzQdS3gNK9i0iNjbt3U8etwrg+lkDYiKwnk8eVa5fqleSKU132sTUwAf19dryZ3
nv88NK0rcG0o2Pjc6V3zafaMbkpsVj9gD2nwZfPMhEGWWEM38Cy8958ZhFxMoeCO
DIWXGMyR0a2S8V8FD5WnktND0NUtsZXvike3nl1iZej9Y3XwFVhirY+Ov+AkMFqm
5hqievBQ/vZPNTAEF+Y3dfSWv3/pxobrrP/ii7kPGrQ=
`pragma protect end_protected
