// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
T0l38jks7O9CKDY8wVsgh4a3AjIYdZ+DjV5N3AfjtKDake/N1OjRu5yTctqp/WloaUkY88wHL4rm
0JRqUGHactVzmVBkceLugPd67hAEkR5XzjXnW0wnHdt95DLqRBt+3swH/xx8N8Xztro2BvC9ujjv
b+e7f5zbAy+aTrYqlkX7KBqB6iDiRc8s+MDGxmnKEtKJXd6IQfUgUfmNge7jhc5Xh9dQY5Q1qyxm
nVEB4rQ+HaH7MVKbSuoF5oQpXo/oZcQJYSEOeuQrNiY+/r/a89y3Aa4ytdw0txP2xGjXrQwBKWGO
aQL2iB1pMaIbrvEfaz/bnUJCRO7MwcYZqS9BuA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
QuA8+Tw6ua98srcnKe2BSk1zuHeoLerp3qVIgVMSHAO2TX9SJDiD+Ae7sJLDnplYgVYjct6ZTvkL
W6bXl0GH65tZnuYjK+kYRiOpfFSWTd57EpAc/Ku88uX8wydob5dYW9p6NhADvcIGXa0P0LuADYvR
wH5yYV5Ns0nNjwPxSJfyZ99Vku4N8Mv5KpVE/jTxzHjyfagjEoaMO+BWQ13Vg+QdaTfJkonyr/ys
OWd3nfwEVTzhqglKU7sYfPdX4vB12us/5COJFzppPEDn/EZh3Drb3ZdNshjth1v136xqV6K1nfKs
GKGywEGulTg7v6zxNPv16iGk6XTS3ToTO76R9YWcx7ZrIcL1MF2oUGeoJeWQxDlYReW1NPB6cPJN
a6qPK9e5j4G4o0fCFWKWSB1ot6MSyfVO/ZOxwn5faqIddkDpiIRAmF5LYLqI3xtSJYqsEEqVVyjs
NovIUc02yauL6Fi1BYaS5HuZ77f+a14346DKryiWQrS7i+AmpkQqrI0/k2uP6/ONWdClM0WxlULi
PdvmWNx5Brkwe7OsR3yQEjp1pzSdWWxVVBUdyKfZZYcxEA7Zjxj/w4RT18OENKOWh1gjWQpVGY7G
d8Ve0OXEdtTQ1M788Qtd0eGZ+hcuyTzOsbBxl0nkUxNW6ytqPv0qxAIrwejypfG4sfaFL/rSRbA/
Biqyjue4rqwAAJs+qKB238uT9v3CCxj/uNDx56ClSBp69cEnbzjY3cKlcD6m6IbZXsRNCkd3wpIM
qDTWlE0ux+BpYVuYHizdtrJByGFD38QTcX0HxyrH58+MtocqjHa4dZmBRLdDiyaSIWJSuvjsTJsE
yrxdLUPXetdOjwBrmQr8w9S/Wn6v7cjPLPkVWoN8RqEHvWy341SECvjH/vfUCg3/aKoMfE6DClN2
jzzr16zhYreCQ5QHo3wD1/8JT8EIe2OhShmxfGtHwpVsu2UOJ29dLl/mtvG9sR9Lt6kf8f7rBNee
eVy2Z1IXCZ28dv51bF/yM6WpHKsuzrB9G89aX2LHEaNWHDIE9F4+KF2AuWBi7aCJixTqqdCpTOG6
xDoD54mIfmWUCH1UWwYT2Zk8x+FXQI+2QxNnjql8Qb6JI1clDjMW771C2jAsR0YOgiOqvzmdl6Nb
crONTGTcypFLviYRocSba7hw8Jz3blQzLGfrsIN7te1iB4N16N6vILD4gxqGcrX341c524H50pBj
q0gNxgkQP/yQcIQZmT8N4SIFvNN+G9YVXQvELf4KbPO4ARj7hbcql3PpKFyi8xhdAiUMv8TBCGkW
pG8JDwtfBAC8g61q9+FUADgr/+t0Hh/fZw7qp8QRjwuHw8LI2h9hSF5lItl6gcY5ttQP6w2E9Ylr
NlQDjLywbo2wR2uu/CNilarh/QZ8BfPBHijU5BBPaG4GJLpdJzBDIUYANggRThgVMSov29hMi1uW
St4iQcgR06OV2a2Qfre1QUYuVRYqcafuhlzu4SJDU2GCDOsb5hEMQbRWpH7YY0Rl0They8ANuFzR
p4ZqPHRt4vAlR7HRJ5BRoeE8aZ/5XleXoEK2fO+tXGuowq/GEYak0/mVHXTdxwDbq23K6b7nhVmS
y6X8cQXmiyHQbwOxexPiiYu+P3THgZ4Y5L9inkrshr3eMWUbAHOq4wGwudwU9e/BDOqZnY51GprC
2kJsFb0EPVuPvlNI5TZKPRh8jK2x8YXhAnO97+7iJxtBLwXjpE7XgRaLQ/9PJycme1QhtJ2alRBK
5sytn3TAMYvLZXtAyb/9pcdMWn2qXdLKTjJ2EWmGQ2QTSSZfGGZcdcmQyDcTG38doqZxUY50Bny0
7Opb1V9ROISR2Qxv6u3v8GaP3f6S3hR6bryoAOJGf84y8FrJIPZ35OwEz/1P9m4n+rVA6QafEAgZ
Q54kPCuHHJSav+zxzmPqcqpEHsN4hswP5iF0s+qE7zxn8dYHR3BqU4A8YgQEy7VlEqGp6kfY0UHs
zTzBSzHSynUq2/GEXgR8tEyFOzyv4ik15WiX17i/uv0CX1Fe9Eav6UHBk8f3+fhj6V14fODoiwZf
8BbnHIxhb9IHwqP4VrxrM4zhpr0qSZgay/llR1aI2kEhNadjZumitlq2sDY4yuUsAUDKBgeXlSs+
UBozsjnEr+i5eOoJk+xdI+BnES2m/7/HmP6m1uJ6Ze+jyWwIqP1fbnCFroUsfa2T6S9o/A8YkXtA
k4XE/d2VKRJxDBEdKR96urVDqnSMDN7z/raWGCXh+TG8vH3pSY1oViGk9IiJKFZeG1/hDHEIC5BQ
/DnoPb9lIj/nl6ehvcj/3mCSHCHpes8mcXByAf/ON95w6aOzzBzi+zCDW0Z+miVuOIX2oRMQ/wU6
eeANujDBYVggcvnsgpW8Lc46Ybcmc8cglYPVM+WF31aeC8n7qk0VioTOhgktKoGwC/3+7YTqE0ee
ukjZtVJKOXGJpmn0HVCuX9+f/NwxFqzDckYvBvStCYr/p2I//ItJMMH1dH2+XW/NFf/r9MoySEWw
7hi1Gc6aqrD1GybsVQKZDTlgB9YsbN5BOz+UN9Ns4ceArbf5IexqdOf5TRfdnszAbznC4n0cOJyb
9Arkvp+1odZDjmT4vDrTJv97l4ecITBqkzP6F6K6xJcelHrc6JgPdyDUbrnDznjQIK75CmdcL+mB
Xh40kZXbWHBK9vnFhjt9Y+V6KeZ71gamAli5oDuGU/ZWj6adr1zYmxi8XCdrdFTK8IsV8hl8TfHO
ocEKFb7mKfGg17XOW83IfeIHyxzR+39im1BxtcqIwccqkp4LfKfgFPL5XOCTUZyZs6Gkwj5y4gUZ
ylFxSaJJbUm0LfxlUN5FmtWEvXqM9cvJpZNzMJWVuTQhKMbDX178SiQyX+LsAyREDFgMTPPHC77/
sXmERUcQ4bY/7JfjBc/zzrFIbdYhqwPI/mvt3CBcxsvYwS6/oPEiLX/0H+1PuA3wiA8fleUHU3qI
FKqjZtCnB7kCP5yI8bujuFm4pictOmMeZUKa0UwYXZAn9OdJLbTiMUs4K1Uh503ocL7yDzXq+cyF
zgijCLYYMcarRJQLV4f2Wo38jP0E9koucKqEn+Uc0/RDHwHkFeogtSDmVbdDD3dEmW1WMzXWzwTL
kIyi6+TN02a12ScaMgrSRUM7Rt9ReDJ6XQ8bgD5cVR6rD4sh1ExgTclj1CG8ct5JlnGgb/JWQvAJ
GjUY0UQuYcVCmZ5cDB+/bEIVqAvQAEJukPbuhN2qMyytJKWnFtCEcBEdZGCTndLXzO7h66ErKwX+
hZXjJmkrDlJXy7NtHjtv2tbhLTmFxs/GGOklfqQE5bw0v7p+EEEM62Kkt9fh+DrD+bmkMfTb7tRZ
l+tCPmBeHdrB+HrNgCW+aanG3Mv4aujqDkjC8BXL3cizjpQ0Z/HYkcd0MoJmJ3w8lm0+WIAN43Tq
jIYEYoGptyvybvQqeX0dF4+JoMchp0iY575q7+Mxk/6yi+E/oCKq1wS/rcFncKKYJHN9oBEEpSH0
qmtEzVuNhzBN2odaHJTOA6PifIG/1gRKbgzmLk7HhYa+2swv0c+6X63Dm92a7DxJFWvcSd/kPO+U
/zPiEXA12KmhDF3YZ/R84hmJeOB9XYocPvCILAsu7gMRNDho3wiTQs2wZGu6XwJZyXAF6f21yPfX
9RZgR9yRfw2Etpub8Ez4eaE21vtlF6D+oYQnYr/CQgPDR0zY9BQigexdZC1ERTmksOpTJpXzSQ3A
Ay1v5A8d49jWTRvI7CLODUGYCjIh/jSlPUgQYowGTt6R0gqg4+W9d33YW4Gw6962sXowlY693jJ6
sANJDVD76GC4U8O/+gFa0zmzZNCz4P0c0SI5rIea4KOqJjbXQbED9ZObSouXlMX1r2BRs5K2a7K+
AcXrCc25C3l5KKWyuX01wKc9N/RLMAcEuipp4zHG0Kgm0Ja72+E4/f9MxL44S4CuhUGMbOQ4Wo1e
RBKP+WkOXJ0x4dXPFl8HA/2KkiNkfV+kpvitilVtnHSZcAVpM3xpUt1xYdrE95BILvSe+ss/2pP8
9D04mxjKa2BEey+BwPTbKwYkZwYQz1hWK04rFhyqxTypnVQJ7l4MZ0TWt+dMJTVreB+Nxor0gMrm
b50NhKK21KPdfugl9iM42xh9MgssN5IGiRaDM1Oj/jQQls66l7VrsdMAnpk2K+qQQuDYVctvT/Og
Tqfvhjpl2wclhu+VRh7Qgh2+vmeH9VpsqXwA/EleJ6ijweP9awi5k2Zhmm+B3d/VSzZ1q+pjqm/G
god+y+5NpegXQWJlt30WaloicGgynxdkQkqhbidfbJtaF3iUFde6GFf2yqh1Ax3L0MMq2EJ7RzXq
kMooqtZ7BuvXK/xI/EPoMpwgb0r6tMwSzRXhc1OFdzqsyamhF4u5X5BLOyNFg1EpsNg1/dm3JJ77
2YUb7ouwF8lPtqwa4ADXNkZRC5dCMXmPJL4U01bk7EMEhrgIXE8HZHmMAy8USF1DnbrlQoBNFMNS
llaUBc2NzwXw+QNB5jbLK9n8q2yueJ7+zIiJk+8Zjm1EHuXSKFCFuw9m7nThj61D/jCUyeAskLFK
4ybKzcHjmTqgxsWgZqOTYelypuJEIKYShpP8G1gMfwnNwiwL1GGILXPpa/ntC78OY3kB81IgNgHR
k0wyTfsKMnWSk4xU3tk9Cjmvjombn5QMCcAHIKs0yFADh5urTmTr9P7tQH8yKnZDjq3U3K4k3cRm
Uj5pd+EiI1IYedRcVraHykoHD1QFl5Z38nNvIKhJuhDUqylsdxNSNbboFUZ+f1Z1P2vRd3ndFIwn
HUAu9ewuD3C/Rr8/IcuCR6SvhlE8wegOwKDzHQyjaWTbq61GsMLSMT4dNeXWxGLJYH3hiOsiMlE9
17oirc426kEmBzs4nh4h1P3JLioTVnCtWeHryd+nBlfBycorwFroOkpaGbhW56JA496tlnt+bZny
QClCyXZADjup8DxiIMJxjWXqivGmf+AP6Id45QkzjCDuNpeXdIkfCeQdMFGAaCnvAoBOs49cId29
+dShCTke4/IABcwwYDAMKmwkr4GzG52OS5wAeq+RywZZ96S8qZvE94SZgi9mvZE7xUHPLA/1aBd3
Xkh1hkKBolyTOdEMVzmM5v/eJh4FTFbPwwQUoHZRBgHHmbZI7gF0WfV323iEws28D6izaseAvh6Y
ZBwv0Dfk0lPcdYnNtTBx0skHnAr2uaHlO5Frt0hjSYJqPNgz0dIuJMNhTZ9IQoovrfomkfFIwyzP
AOoCT3L9jZx5edACyeAveJvYnr5ZetERXH7inpj2L90KtJEyCwpABKVT5JFaYNGkhmOTc37Na9fQ
EjZlrt1wjxV0igiO/RuefSFu49F0AMUes6aTOzz1pit1qLee0w60TKoAZlNSGH1BQdepLMe9J9Aq
866Kjp+cSvIwutdQbf31C+8uf/eGMyeP6ccVWKsBJkxsyGqb7bF7AKUgwtsyxRRqNpQplP2AaTLm
kZKacpiAJJ4ctcqrGHAIp9iQEO5tH26kDNkRR/JWFFxP86Qc0dm4cJLe0v7Hb1zJIgyMoo1TInaG
UHZlMsdgySCWwV1y1t3lzKytTVGe/cKkV5Sr17RxrThYbRgLu5ajYf6FXA72nF7sGuIMFLhv81wQ
3ix1KBUBB7xNDFjePWXA26ugRAhtH9ENxyZmxdSdZuaBmd1mRtSC3z7/GwWp2IAJ+6aqedzVq9NG
ZBhN+ao6znqHf+VP6MljF4qgeSrG8SzgyBHyPaIbB2rkoKJ9wS9cXBcgXYp/fZCpVfyBn0NP0AZH
OaeOnZoNyLEuqT8E09lkww13epYdJvioImEVZrum+9vm5z1lVeIKzTNAVhPlMDMwdVXqszP0qWzj
/77ksSeMcJAsOShsxYbisESb5A+mWA3Uu9/xQjcVBDMw+UyJ9ADhboEHseKLjsnfld5SSJfbvaEm
llajOArsnaKrj8jDDWkE9pPel1v8NhIB+pZS8hHu945flHXPPkwB1KHm/fTs6rhMjiIV1PotbIzv
h3vaXnW97sphd2Z17NGQhFlq8h0gPqMn8nPPDl6Jj+EovpYLoxV45xQwHhW0D3LHMHmlTT9wUOXU
tXBZhTUGtQHXvAh50Z32npVBMEhNCS5buBSBWbmV/GbnZqh3wgP+9+Qs/t/y+lH1r2gAkYjRmCwa
0Sr23BeOeJ37m3NjHHpon1L3ZJ1BFDevXbm+ihC4hInANdq7HHE9qafF+wLUSI/Ncwu9aR1KB+Jj
hu/iHZXj/FI3g+FdfmwKALB+1cTkyMWaeon9KAQX8xQ0SnjY4oOAgKgcKTxyjZLdqjsVydrY6+C9
MS2dJXnRuVR2JktL5OeIXP9dM7Ua3hKjdS9eDgeBM9u9nDcwS7npVAcUZFkR7heAMIyKoCg2cqMG
ahg0Bz879OSqXrSuNd92JZ7ONjbIBoSxhTekbEBwTf0u47g13/1X4kNCJp+I3CFKvhrir/KiCAd6
lmNOpdMnneExi80VagvBDxFUNJxyphG2mIh/6K/SpzaY9kH0Vq+O8vv8pznQk89wba07V0mnefjy
BnAFK2PDOu/80hFhW87ftZrX4DwxMHO63HFEUoE3KlQHrJTedmNFo5elMcfyANE7+jlD0BM3v9ck
I+Nhr+WTCtgDe9ABs2mQNmE=
`pragma protect end_protected
