// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hEfSy395ci40rWIfTueBJNMZN3+CTnfEYOoTRQSQOQhik54fDkCQResckGymvH/2
KsknxQUY1FHU+aJIQMXUABJWFIwvzuNcnPrCGXtnB2picPOai5yO34BB7nQpPkKj
4iucQ14RxJsTQWl7IqRj3hBZkTSzuiMPIB+gM5wu3Ro=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 41280)
/YmPaMr/1N9f6ORTS8s8V68X3nqNAbBLC7Do1q96ksHH6d+nBYzAIXItHajiAJSJ
DMtzZgHG4OKEskKGuTT2XW2K6cHcoTHuVv8oeDluVLbrwcjSf0KYMo5PT0sYBd79
Sajmx5ijjxNrRPByp/E0j4NrrdATKwbcCOBEibZofMBDc+0Xukn8236CYkPrTQFN
eCphCUP+YCZ+a3cpZF49VXgpqwEO9RH8xsmyr1pj2Bd7ci89WoHfqMu64zbxB2Z8
6ztEBoKjGZDi2nPNfiLpoQBiDHdTcmVq1skPLnm4hTaffhFvaLGxXEhHTPLU6+lQ
fL2rIPgqQnWm+IztjGE+8C3mfDQH7SBkYfxvx8au6XQjPY6SXOd3Di3LOO/QU2Af
AdjSifEeplEgZi/V0M2ovaeG489O9M10cgqzj2yMEd08taPFGhWLvmzO3n0fX1IW
xmEhRp7BLtQcPCiJ1LMMZ25EGC3+opncmAvA4MP4L3Ub5+E9ckvMVKVJHjY35VvG
v4hNLXlsbiVJYYZUVBT1U6u0zDMlVtqrw+1WyWjVGjQKQJyb8e5nSohLYfrsJTht
VCasWX0zcUNWOo5zQMRd4xdAFsjHOs7FmBWyKT0rThfJSfPZHdlC+tr7esx1I3ML
6PEJyEtbo0m3yGpEkaX2dnlku6pGuuPHYm2xk4/ol8mF2erXV7gZWXH3jLahDVPB
Vp/e7MnNlMpp0cpULEVKuZPi8xUdx+tgbXQNIZEZIoUgfieq4FkO2oP9vCSWAVEy
jwPMERue6J5Eb4WeBZ8zKejtr5VYUm0vhkbYwoXRJoHifklBDF/iLPddh7Ux1/Ah
8Tpx9sc+ei1JlrZwZBf4t2zlM1CYmASywlA5UDk2deMlBwt21xpzy1ydDgVEUrhl
pMhuklPIGjgiMUFtY7ZOf0OM2B9xhhkpIkN1qyTf0IKvR9ajWtgKpqztVdiFQcS9
TZtm9VNjC76qR6fJbUFJ3B7UDVwIoXAfyZNoOESSQ3V80kD+aE1M/dvWrMZAsC3l
P+SzXXhBzlHS7qYZ789RrVs99q5Q6t/qqdcL6LpGOLJTdvLJy6EGh+8Uv1jT5sLi
7GR2FyKayJVqa1EhFXQMJ3NqjDZDQ7vxJUXISRH3OMDfiWmsn2lG2iRBD5RydAT3
JS1+4PHCkXnDufZXMrvTA+RWQd3+/0uXdF2WXgOYY2HZdGrSTHyB6W2KUvVDP2hE
PQonLrQw8fxSepnDG4diGzJpy3Kb2lXzZTBMHTBln6o2DmDs16tTPTCggk5ySU31
UprowLxN3gvat0D874kPvDmUdrxObYd7nsnKOWS3XHZOheYPeM7MErHvmn7wZwc0
/u4DUqPNb8pq7KuWU8Lj4eqxOyhzvq5i00/FkB79Js9d87N1MnFeHnzMrS3HqMZ4
ab+hQyBIik4dc9/RNRusP+mO8tj/8L3L/xVkn8sUO2ow3NHsaGLKaNI+Htv2cjjk
WyqK8VHLlLhTq1ICup6XucwB/Ru/vnPZXqIiBwMUDrhzlJMCcBrz/S01KtgCOjOf
wett9iULnhiwLjDDws+LvN5IEdjipIQMHKmnWrskClry1t2AkvwRTsUJ4/s9k+Zn
g0/VZlTGTphN3BdIyDXrKaGE0zXB0uUCJbPMGMvyqX+hBzk1vkBNa93R2ToUbODg
ghcFMlPsMEP5DANtX03jT00INNh1ZuabWh8ObLnqBdN6YSzxinBMaTG5/y4vFBo6
aPFz2O1b64b0kACYPva2FyPnuKhGpGTccbxZPfjP8pumhrXN5IsiDrD8sDrklQpN
57PoZf5jGypNxIadHa7S3Mym1tFkzOhCH7rEQg5FEUvBv4C9yyixQzK6FCvYXW2w
8U1q4oWzbVRGIKZTJ2okTCzvw4jKqnOFohZBZqYelnavQwUri6W3SI1K7e1uj7bh
HXIgXXcpZBcHCjYBmddQzCbupZYuZo4HAeW/LaPdxHdbcgEWOwY4pQN5d/zh5Dff
TX+IqDK1Blo7usOBR12KB7QMXcut6SjSYBqwaTVRToCMeIu1Iw+il24h3uAVmH8h
WSrqVJwjpNNBhgwYBXDlTuRB0NTkPa01CP1cAw7Z3Wk00BMIibVY0oZfB2QR7mDE
hBv3DOBbJB0x2UZlZ4RFYVWAimXXV6hyLT4NoLMYmU/OO0GHEyZtGWysOe2Sc3lj
AnztgzkUKlx8K1Ls9XNvqBYwe8n4dUcGNwx6tzYekUAtfCHg9hFE54jkIeFKmnit
O0rjjs50ftUGlQoWhUwU9T7kX0VJvmC5PF+b9JnurNmVhEFq/39bTBCKvk5fWH0T
cHkec6DqhuAWjCmMsRitUcWissiWb7sDwsfKQudrs9AST+KkZ+XhDJK9NvGNLLeV
uyqG0+W2dybSgrOSVuO9w8Ji8tG8FMv2gjQZjR5MuDqHtTDY/ynWs+2wbLBHM1QF
H8HCUvdvXAELy2MunDaVoTazxjoT97uQ5NMe5h9m727ejbbMcpaLKlM8Z8oEwxW2
wmp/XhHEPjWUOtoTWP/JBwiJb+O7ikpVasKb3ou6WyzRZlJVjyBFTC1tUg2rdua+
CvL2eMyo4Ra7e/Jk7BvX7BO6isBWnAI94n3iQQuNePV8++gjw/z2kuJrgi8f2LAg
qGtlfItTaKidcof1icplFCMKlr/4Eoli0CHtHdLRPfc+baCpTVqFZVO1uncZG4gi
DswT0zFhoxIjsVTE50QU41b0QvIa0KtTMwBF6MJucOGofvVUnGL+IXXX6ZfmwZyZ
iqxQ9Eormo6RjsRxzBfnMs+BFquuXjBAH75qG+fqWdsGmiB4MeDB4KFYQXt2eNtq
WCMnCWix+jWp3WE2YYyCxH5DBr9gpryWIrVZzSxkiLpPyfiRiKEK4JLr4rbN74/8
YmWF/ubJee68hwsav9iG+q1QpbBXc0ctwZ2W8o1NW0gVBKNiQYQYJjJM9y1uLKgN
XXNJ2bQV8fQOQ+6Z8fR+9XNsx7b5Pdl021kdGhOIG1YT48QcjGR1jGBz9vkBOAga
iUKzXm5H+OXaT9k25eo6U25gnDyRPEkzYeX96mZZmcUfRBfXe2Y8xbh1YH22m2al
TbvSNocEo69lnFAsRSPIKNH9B9oa0z/6pbElPji6X7fvXDfhqOjbRfNaynpWvETZ
bkYUEiOSroVGnlJRDmIwMCKbhotqKizQdF8FDlWF7rki9ByPg/e8rwfdL/oAD72z
JdiMJVcQc9iB+q/qB4I2TlL5d2SWfQU6UWRs0QoDj3lYAJ8muixeL0FveQ53Zrp9
1e8hKXULq9Tz003R6yu65qGLD9PK1NXoAZERsIpajjVTUv7PGma+J69g3FQVzokz
++Qf54SRY48m+iTFtpRISZ7Z2c3ssn8BcSfW5BLTZZlJhd9hNTnB24k+8mOxCypl
zTkiZvr95tPWTIpW6L+4fJxs3SfTMivAKp0M7E5vr81Tx5ezV0syJszir7tNEVPi
6RxdScCLrbq0jqp/MgfZYmNQUU+IcCkVAPcspQHeE8RSKaLfradkrmBQ8V2UbmGQ
3+Q1RZXz9w1ZfXt8nC7vVwDQsF69W3AA3X4extNoIW+zwhSjjYFmELQb0Lxc/8t1
8viikpB/or5pkONhFl3IPAJvY5YBMndeIbZAj2/gihDPCakKfaOV1o98o3X/zdyJ
os1VZNGez+wjsLtiygHiVBQX7u2icaDkKGCPcgDNnDH2VHRgwUgi5MBvHZU7vILo
SSt63KnfZc1UEVz5RvwFxvqpM/K5uy2dnNfWBcLYks0w0cR8+ni/eXc8bbRSnFDW
lsvNiZRlgiXtypTwOxAdCdLo/6aQWNc241n1XKM2/cw82oYDNfBtdB/sn/gY5oNH
y91h1lvME2M3ESa4snXg4F0Ml8eWcrzNjH+mdlBUXBQPAY5NlZl7B1bHseG6C786
mnY75TL0zUqCvZb9DDy/C+RHsI1FlCqMM57v97UZjDJ2yFxuYjvC+llJ61nqlHaH
/kXDBqcjhPoM0o8ULki5Bt8P2I3YQKpMrGszUbjEq2/aKCnqxg5sWFxF6J2xyg+J
Tj4oYzLq6J1DT2zi01vpyLr14VY+BEb8UO+4dXv4aJ0cYYTE/SOcLkWmH80H3K7J
6YPzUa3FvocvHf/AByXFc96BzzoLv7JcYfTm5K2UTpTj/ueiIx239eY3lXHAa7Mo
e6hE1CoQDOaAf2SrG2qCfMHaF7lGNli9k1SmWTWovMZvYlwmN2rAboVSoRWJGi75
vwpaSitTCZfnfjVQRKm+liMpoGcxjF+bYCsmeBEMVfSKLBqTaaOnxi2QhrDhfLN7
q6tkzus9OmdsTyYLbDdGUbvaMzxOb/IHgQq4Vpovu974SbKjH/AbyB+DbaOUerPs
qbc2tPjtDK5iAEqgvnn0Rvd/yZDH3K/2MlQJRvjkwty4Z4jnaeECMzQE8+qtQ1s2
nGvNuTKmC27vu2eRc4qSc9bIncOFh0bqt0yJj1JbBZLt9aunxTUcINQ0oNUx18cr
XpHHoF99yHKsR/uOQMunTsE7lVFezlnJ7LqjI0HfyWqyS3NfTxINuxh9aKtnPlsv
Wuvl0lB7smKpnBav7pizqMRYfBqFKrgBzmjU9w/L4IhZCQcAPT1l/HBTvqRv6OWJ
WS+KbMEJRXykrRv25CP8jE8+dMfP4mMC8mp0WqYQ9j/XCPa5zO4lhrwlltr9Lgza
/xmWkHzx4aw2VDdre4UT+11P5XUYDeaeET1rFOci+K1Z5tYGzCjOb+ChY3TzvbPl
osLIN6r5Dej333aMI/iRff5BCYjr16sTpgfT5laOdVhY4LYII+f3pKrXaXOgWLdI
wFjOXkPyISiRE5TpIvhYZRVj4fPSVROskRRjCT7+b480cnmzokgTHJfq40KSsCor
RGL0Y5QviI52VaKo7bXu+KOI9kyDafg85FI5FCD+agCHDHA/UYJNoWsEjAe20A0j
9/Vg0NE1eb//vj0aYmK2WwJj/OsDa5J1tXmC46lULbAWuEQhgabqI/n+c3mUSzDv
AyOgMp8oZi3zNntfH/m7O8U5RB5jTaoFqBYdYL4rBhP1HHjkLC3QxLhzorr283TG
EPjcQjIcUIPqQYyV/ssTfmGuNuZ08j9jnVHJs2JfaA2aeYqOI5TEJesEeLzV+wXw
yUdY1BcWg1Mh5+KaAVKVFDPgUsvFyNizhdzsIy8gLP7FyJDgPZjKmiZ5/JvKgfeV
pXVt9qmf97hpi7p7JbsSMRWe8Bdr8ij5wK+XYKj5O2zJ3S2YA50sxChFNrrFDFNU
FacmEiKcCLlf462gmSjLipjzsNHtQztR4o9a27G33BiuMFfuMS8jLPBj9S33jHC+
GjqO4YoMvKjAPM47xKtrpt6Fw6dcRGsuw1IevIgq/P+GWEZ6JTDOSsHgaioCWzjN
2OU1VhzDhoDQxmpYxY1pyPKq6W9WinT6wk3o9AK0AphrPk2wJVnw3VbQIziPDUks
7RdPFcnvlJqSUyadyibW13Wlya4/pZTWLIJLExXMBDNU1rYi9ylo1uMzsijzxYnQ
yUUhPgntEQ3lGuCdgeUG5t0fVihtHRNtpVlsYTjujEcrUzcacT9kHgiyYHMcUKMb
M+mzzMisqExqEkhT/NYtHlu91hoGOfVBXeuaqOV0AtxBMLACHAzI911reh69JRVc
JXvipN0MgeEUxxeDj2OQuyF7/GsRPQR/kKde8mp5RuGX8/J6Ay2ZZ9x+rXi09N7m
+Klr5FWO0xT6fqGgadYs91eXBFZZFXJXGiQHYwWLjMzP4yuio5qZ+czDRb4xnwXA
gYVy47sdY4NsyLBxEjlT/Gb11iixQ3pDImABoY72fQw2NOJWth0EbmobmTs5241p
iiyqtjJEi0kwaUMWq3/3WLQYRRSxunMt+haHqATJl5YezRYmvhKCfncF3JFeQoFd
GAFUmVd+LgLoyRR19jx6zjsNcC7jA3nEUeFauB4c1vxBPoMnHNa2M1vnLJFwXiM+
s6KzkmksTRlXVEzAoLhfmAWqYDGwh55U+g1ndFr0XrrKPm8/Lf12nE5VFBdpRGIM
oTzaEWVU8Tui8gxLnzBhFPbo7/MjhXe0yTYVth5LPj0+KG1VJeCeIbsR183VrQys
pGPUP8aRWQm8dOId1EFxUQFrgmb28Gqmpq83utGa7gDtKIAI8MSzaeBwHXue1a/x
ybosY9jrjTf5aO94YHoHVsfur56Dqx9ipX9WfmUFPnf0Maya6liGJRg2RCPDcPt3
hN2aD9q2NUJW4QEMN6lHwcOiw4OZJMtQDngfsUde3qR6VOveuIkJpEbcaoSWqxYP
qd36kEy4iZnjvqMgpbQxLZnlRoAiXOgyilNwy8v8KrE6zzFGJrtuuhT8dSvdKmzO
/HoEFJ8wdyfmA3bLkSQzSfem+Y9V4rrVWJJ6q+ttM0OUb+myUSmV1s5QMQGetI3M
YHQZxuPEirsYyXidcy+iNT3fvM+uC2kb1Lt4DQ6+MjvtlJL9z/tUHGGvVzRiD072
qQVdfVpl940Xs8I4g30a2pp3DcplzeqBx70vujQ1yf7pPxW7WA0wWuFTVbkyQ0DN
fyN/Ymtok79eFaDex7C4LPNBjrxLFfG1vQOpIDbEtX46Y4dRiVypfERSMhyCSwvC
P1wIuEZkoE0EhWwxr0OKN4ZY4PrjPvFgQu3VQGgmJx8mYlULFylFAKZ91VRDBeg7
mOrAsxlmsMTFjM8x4QqefcCEEbyoaOxeBtb5OqNzAZ9wjHSPTTgLcIzl1aa01MR+
DhaZAK8g6tWcXJD+Na5J6Vdm6VTo0BRZ2oHznSvnRzqAQ+Z7kdFSfo4A6hxgYx0N
7CT4jSisK8Dxz18nJayBqCewJRwbSI9upI8IVjktQniPz33qM5XD0IeCAIK0f4Gr
V3xY9dQZExnNqA6xpEVmeyhxB8/KhnW9kctwVgew83J16SoD4FhKgKLq7uYgM4Lc
8peoyycoVJlbVaJ+gtsGLkC8C49FIp3XrKTvB8uYDWhutdhNbYkk6GSQ+v6TtUBJ
M5gnEX6d15WmvLJVR+tqfHqMTSXRZjvL/Cj0EzNp/7JIUMTq5iwoafJCeFMuhvvr
rkaZwkCM0Aof6DjcZiRrW9brmE1iBnpGq3luK4kZjlCxjQYf7vMGUDIwYm4TRW3f
soYTqrYUz/DiLOw37CiTI2/db7/4Koe915dqHUILtNh9ugeFmo/Pag/c3julj9Ov
AnHl0JHjHYw51ebAtYtXlr8RKCC0vjhpqEJmt2QKgG/KOlOunBRieSMIbECL6A1M
DwXvE7fwjcPIsn2Q7oeOaFMufIRi8eGQs6ZGj6t9Uqjp69ClQ9Ltx//DM7lH5RdI
leNCWDZ5xLPiezOeUeMF6KjvAuByK3hpe1qn/sG1OqToLPpVKywVENgaSRyRq2jr
0aAurc4JpZeS4s9V0vhGbsKlvjFTIJHw5M+GmM9QDN7HpVBMd4t39RYTfqQYbHvX
ok7ozlEnGEWkvU98YmVi5GxaDM+sNS+3GMO8G9CYnNj/L9gEx0Lsx+F9bE45hPeA
KB4jUlmuzElg6lwZYZiaVFZSf3HAHp9HDgEh/lCD1OFklMQm9J0QuLVRjnC4n777
1eJpKSAg5iqs7Q2bZ29uZYg7dOu3B+HzZXePiMZn9tzBR3+X5jV+qESp4aJ74mJe
CA1nGFxWMpiV3AFSnidOSdLoG7bHyG+DL83euy4+0wXNE0pbGKLQjG7h8k5aSheg
tJ6gV8JGqRYWM8ZCNxeNvFqjOPcieHyaBH76opBg/krtuvr7Q74X5BxnGJP8UyPN
LNLMspLCSr6utcVC0IwU85e90MEQMkCWp7+I1kt0F1iRNPY0HjKI6yq5i/UZK17/
aEwN8dWbg0YZ6MVgAwxwPkcRTADeE8383gps8HZXdb2tOFWnU4LaLPTzj/e1fxLZ
tMmqQvFHRkNOuh1BCWSiR4F+aTom+SiyWg1dVbJWNL1fQgWhibJ9AHCjIchXaz2a
RbXFiR0W/h9/My0ecc+tbtLiwa3OcsRjtWF6HEgtGqFevGM5xaM8HEImyj+bAttc
iqXzGyBW9BmppG1wIEX4HsBK4UVuJUEDXWKDVpGIsvShBuMXSn3xilNcqt7C/eAh
o8p6MLZvUfN7X0lwEeLai7ust1T6jZyuYm+tGyAHKOqP/keEFjrFxAn4SciBHmgh
yW1recsjg3MqT0f5c9ZxA4EJBhnS43ee+1fB8nN5kS58gT2PxIG6f+gMOfYYoOTk
puS9EK1y0U7ErPO+HvLOR6SiT/RUppMHkoeBlho7aHMdek4KcylA5o4USkOHSo8W
tdV1KgK3vsxAWyG9MuOKGvYvVeDvx/TAtGXfv9ddHTcqbYnJac8+16fgqchB8s1H
nb/l7kj+WtiA30vsJqPRVce1WpbPIW9uiiWkm/3JlWOzeW0YEHXGyffbUhlG2+DL
mgASIDI3PqW8NbErG/u76Il9hFNdWWFhEJpxy0V/dHIz6p6EwokbxqjfezAm/e6K
Kx/0qlqWRn7+a63l7XBvbPCQMpoqDkTBhx3SsLWDnkOVcGsFLhxyB3G2lEvmCVlf
Wj61rgwqTk/9DDyS8A8McucwiG3t+TavDIt2r7AYO9d/DN9WmsOLnNN2VGsp9ZpN
msOWTAY5+wf3sd0ZgCu678YIjC8tGzBP+bFURreTxR9sYrDkzZvHK4aJMYnV99ek
RBijLAKvTsm7+Zy9od8KUc18ftd7rHQCQwXWPkJ1cqe5AVQkeAypnrnkivJsjRwM
tt19uSNyB4p+FUJ0caYrbiE1bz47+h8ZAjxSZTOW6AvjFyr/VujpeJH63ChaFSg8
GWgupu9cK+Tt/9ZH2xM8zsIzl7S2+zNzeNb33dfni6+mUe0ecwe9OXmb+divmzOm
4oCYzNCWjXvrl4tqf1sjc5b2xdEz0SdfUjtFzqEQXWMy/7vKkaC37SvqFZUQNJy7
IQzcNWp5efYLXBEAnMh5tyhn32INEWdNyQA+mru2L2017wD9Xm3EqGRyurjlatPa
eqfv8vbkJz8/0Xtekyz5IPDP1tYb4h3dXMiwmH3ximCqSPc/jsu42g4R5BcMENv6
hiqb5YJJ7IZrgNwlnS8sKD12kIfmjVEa2/h0ixaz4Ifk7lKb+yT2LGaOjRWeEy1A
P2kj++9ODpPHJiXJ4IYdsDgsHxhdo5QtctdRsMp8E0KqrgjVYABcVHhdm08Ikp9R
vlxe+DWE6tAf+C72CJ/NHDJEG7NYe9yYa0B1ucylMQq1VdM15er+jQZzjupMvOP1
M3+Sksyr4+S/aObZvhAcMZ/KU5B3CopZf42yw4YHFHZ8OIR80lgWxhlhass14qMw
qgKNVF8Gi/FXqAJ9lEfoYcoJb/yGL5qoi1473GsXoDiZFM8r7O2Y5jd9JGWOcbS/
PgzOCSzzg9035pA3uroM2RZ1JJOrqFl42O4m5V0A5k9eBH2AXC2O1Jzb/YwxzyFf
MEMnFgwSh2TTS8q8rylWOKswBCH+mxqin9oom/tcu8REoYhanRmfo6iDmjJF/z79
rSn8dAFFvnv9Xn4TW0jyaWvu4fJ5SGLZcOryZFccd08x1OniKUpRCY6az14h+UBa
+yS53TjRrURN7r0C/6HDbmYqLzb4E1RiWcNnb2fgLQBn7dNtaR0n4FzT5Qt64ttM
7oeqr0HPIIZ5jefSFyMc2VLZD+VY8FZGTwCFtEYrRDPvzwRc0R/mZCRI0pPXmrs3
L1KVXaHrGhnB4KM7sbz8v7k24dM4CMkB/71H13enrjQ8ZlYANH/WIfWH92+BRrsi
LnjdIT2TGqPDpJCKuT2ooZ6u4JN6k8Ug3A8ahM57T9l2VV52GnZnKZpaJeF3ejYG
nC35qFYp6bESjcoCKXATtsksuJHYqLEDFOj2+kGpY2q6mS9s+pftBQ0JE783T6M2
sMULd52gct9wDmxdH8i4u7GNoJX0wv5zFQyw3MzTqrO4D+xd1hTB9UGbosVdMOBZ
CM9iZ5iEij7NCmytsVVRQAobCSAgBPYFSYbxdaaAvqE4b1nKldR1LqGRHDl0tVAL
bR4KKyGaVvAOfQSBRBzTNwIoLLXt6qz8f41pjERwALubOCFR5I1n1FK6lO3TrllV
UQSCKB8VOoEgcp5XvbN1Ljs8lpPqD3StGbsWQfsH2rXWE0pO98iNhhxoVO2Iw9QB
yl2zWOeIcTpfLHsDccTmMUJsCzEiks3isKOX6KPGOTYBTm1dzaBAVrqICaqB/+3/
ViHGMSx/5or06vzYdvwGEpBqIgEwDLrJSQmXoULHhFA1hBNvGISBtyJeT4Vmj0p3
WCJlvDAT0JtNNynFlN45xjgYtMQmjNZEtBM6zXbqQrBR7FiRhFhAjUi9oaDcT6QX
59EOCazoNNtr2bp7zrfEyC0y62YIDfgLaJDv8SrXSld97aRUHtAQ7ok26pjaOwyn
7D4m0c9fRbqptROneujOl60MOqu+wWMFPMYooiGrSuGPriiDNs1ujB62ZXkjiUGU
T0/lcK84d6br4OPUmuxj/XFrwEU8dxKC9GQU6Gn3oRufUSOQfvaSVN+7MoNiFTuD
NT/u9CGbM5F3bm2oH/pvAwXsJ2E+d8YdR9nIUDxgIPSJ1Ml2eCkTvfJ/RJeO3Hn9
K5eukesRKFEiaeYCdBpakzviNtol/uxNpXTus3GdKQZqeSfCOpf8Pq3mPIEIgsxF
Qd2De6hYPVmkCdBFaodqUxfLy7aXlTmyNnG1pwKCaHhrYxvWcP95aPubRRuydOdU
FfrDvbJHaynh8hojc4HkBRMaOieq218AsT9gzk0jBxQN68mr48NHIoyiH9Yaazpr
dipzKdYFSOv39EmsCgN74N5UUcZTF1F9/+N8c9NnJ2y1D21lCEtN2RgOZpIvyQSR
u8ThdB+M36WFFcPde4XW5Lr5HWI2GukA7rhxHGPT/H2QKgFQRrwe/sX8qZw6F+X1
4J8DTCA6p+aL3RGtfu7b9dZp+0vAoBEYiu9i+qvKI5EnfaGdN3kcA6m6/H+/Yf4F
nZePqoV7qjb0Lc6HBXVZTS7NWKwQYiIcVO/4jjav5JqX/afD+DPKTz3sFdAQ7bat
FC9TJ4U/EwnMZNwYMW6Uhz4VRLLF6tCA5h4dQrPnlQgU530+Sj+dET00CpFnbDl/
ryiqeywZ2zZR1i6C89avDbQ+9F3/Fz3cTeMlc5TfUm9qAIMe5sphomDgQxOKTnqO
WG1WU9RICz60PHctNJoO8bovQKDUDlz06+vuOdTGhoAN8/HrZlSXurmp5aO7fjio
xowgUHXb+tuEaokxZFg0KNAjiMWXXf3d4KzPqZxOK0opMpzrPCNmi0EBZ6KpM1AD
63aR88rE/zNG5N07kiKPrbs8qfekkbJeHnFTbb1h//H+fWJ9B/ELa9H1RJkEJf9M
kUF9OIX6z/J+E9/Oi5Xjllq8CHFKWQk6a4/zscsz/GpW65m0MV0vGVwitSLrElFy
3DlPwvMI0yKgKNn02fT/tIS/a66C/XOCvXcH/UUBKFWLnxmWfzthiCsfsyix+QXf
0pdWTqj9ORht4xoib/+6Kn9O5F4MIwE8HeW3x4fKDmMA3Ad6xzTQII5RwaOM6QIy
Z14BrYGvsXNTh0OAIseLNwQp0IMrDYVVqc3+TxSNzv7cdKm+cHQ7nZtUtB/qo6RZ
TBG8kkrFakhS1/kWu79qgUlxlQa5dqst6l4mEOXdjKRxtct+gZ6tKQCXnq2B1645
O/l6zzztr7g5sYgXqsA87H6te0uuX+3qs2OrxD+Y+ePQ96Ysc5GZlus5VgRYvLaq
79kOU925J61iK6qtZG0tr6923I0lkCzy5OPScZ7CtgxaUSBez0VLNmScnimzcVlS
4OXXB+rqolryI0uaVZJPfIJjkOvtnJ/590//kTVJcBH2AKEkNeMWvDfsfobSPvfh
T0H0ldxnBBcsmv3VUUvQ6bzPl+A/kUSc8tL9G7kC0rkhKUHa9CMRVihFI7J91wgw
TtXpCvEJI/maBXBzKGO86GG8DeizqDNUlB0C/Skik8lKxzW6tUHuHJE2ib+bYGYY
QCKxhaZB20gIL3p9ejv3WZE21BZHY6VF3jMclQZlPHu57uEwdIbxa6D+SQ5PohLD
GiLmv5WawJGDXSzNVjfnmj6IacFp0GkEPGtBP7umnXU7vO7h3RpMszP0qcGn5kEk
AVmpmA024fBwoUgodDfe+/WyzAbpLx8bYpCrmlD8TC1N0e+fn7sGXESdV/M7ODmO
kPV4TgD6HD9tZjUndBQLFnXECzvT1C8RsRo7lkFlAdKA2RIf6Y4XFmCeYw3h0VRi
G41yOYI/tqWCMoT805pWCk+q00cJJjKQQpU4kj2XdjCsULehWS4pp4R1RUFOhhWg
EWr8Sf0wZuAieeuBjR4QLw3Ng5wuGK57uvMMKpyRIufgAASwEJAqAuhf15MZb94N
FymHrc99f+d0/YmHUygdPcMW/yRdV6nMU3xckDgEaOwQegeNaHpBGnVEORB4GoLh
5NclFUJluKK6vYwC5DhVzbyuSP2YoMtmh0DXOFlWbc/DXH7etN60vziS5ghqOk47
l6ppzlJj5O+F1zohGQG76/95wzM/IxqYt8rCuQTfWEjNMuMr5Cu+6AvgHKKfVnXv
S/qEsi2zfbgPZMVQqKS6yKfsXY81r9+UU0lKiXw+UkpX9R3DMONikkXI4U2+yQbz
h6+tUZSUl32c1jfyPMmBZ6yrw3QybT4e13QAteNPm7cCRe8R2fUNJxmZJ0Q1D1Nn
WcGWLVG0f1rk4BjgxpEK4t21OkUWIdeH9GkBLtTwiNIeCUymvlGGU3tOV5oAqMAK
AnuK9sF4Gt0JFbz1Mc1NSmfHpb3cHMmqQySsGcBkQUyc1ZzzMN580DsDweC7Cef4
AMEXpSqcI/OeBkIbvvWKRH4zOgmhHtCe5lrlLN2DjTXYmH+l5nW6pkEAkmQubWua
OpzWFCO0NB69mQXOgQGq5oIByp3bcWbJBM9IM5z6KtdpKs+8UM86V7Vst3uJaKpS
6K/+2NhXaFodLwfqF+eSe2VvweQzzf1BpqGtOBfHGB+g+USRCu8G/Ngg/+7lai+I
DVExd2f/fEbT5fmq3vk654wiMQfjGA1bnaSXfxXrA3QVxR101ZL2kgr4eD+O/iM6
LqZbUaojiyUTFMMvCBGtvNrevkkn2xILOfTgnUJGNshaBh3qFsfOjiAMPCvZ2fw3
c8eUh+AWu6ytoePen92rdQVdxXE0a73yVLPfF1qImbNr+WTBoaFZOHv9Ia9pBJWs
4XcczIQv4m3AklW4z7UDUbaONcbyFO0MqlpTFUEMELPdZgKq9KhfBQZDPqi8t2SG
SYSOKUX+iZ91SxUg2Yioxh0haosbbOTCTkeaUK00q6Mk4++73+BTJiOMImyH2HDg
pv7vDFFx9Zr/BbHgTjTt1sSFWJ3AOHyPaLseqYugBoCol1zxWqh4TclA7rfHfuWy
IcOVnCbjUwpMXH3f24taeG0ojAyZer5qZhBuy9V1pJsymKQnlA8rF+IjYIh68pK6
fehc1fUe41QFjOTuWYwcsZlXeX2MNVfM2VdOylX+NQAxS30xzbqXIfwLhx+llxvG
NTli4qqJA58masGPB4fchMMcq2cI59fIdfV7uCDYkntJmcgrdej8ABc5SvJiMj4m
zAOLBiVAYkkbE63J4Ti1sn2zqfow6PXMU06cjj8CiUCwZsJ2MINVe33Scc3nmkCt
6f7baFcmjlSWoRroL1GXdu+l6U8Swul6wqkufNr9ykh60RQ4GSlBKBlHrZroHDrm
Ey1GRRRVfX1/xs0udq0PnMsVVbhJQ/x8tG52u0GFCZnUu+bgJgQ7w5GHwjaOsBBo
yU4QXupJe7EQS0VzTBJ9QehRbW7tF5OjxQcpRQB1sOXGQQKPVNsmMrNs8ciI+Lk+
Bog3fRGj7E3ni3MaqjmB48s0ayBymRMQY2aIdgN7PD/x30FtHpXLxRdYLLUUZtl+
2p2nrfe0LuyWQIIqHtPNdtsSsXTvWedclWbRilbgD+Kcx7hg802B0mP2+vsI2PeF
A0WJDcI6tsaFu0KZfE6xPFfrCAp6iOWLRNskYkBWhrqgHiimaROyokaL+jK+WDHp
9DRq8VfQWAICqE7kFvH0OoRAp/0oxADL+CfYCthdHrUjW1HIYgeYeFYFC8tOMoOW
VqFBfB+yxOojFm1umMgx74VBm3tsmUkcjlNXwbTP5QB993kWWLw+hEKAJr610YSo
qFOECFrs5r01DrNOOWV2Xz1uRFRNSiUpnt3VwBMEiefQ2SWvi8uaJ8ba9KICvFIE
UATgt+y/MMkblTeTgiOjbJwA0zYIxTTMUnsFz8ccX/9jI3ZV7gu+ThYh8oW8FCMA
dfuyDoGVK2dMzxe8cys04kuQkIr2IzYXCp4bXd6Iy0f50ql22Xr4T0aoOTti61Zv
hk4+g2GecznsHTd35yzTkJBR9fCdSvOR+OQAJobuJIHT6HMxv8biqBoj2xUVt5Dl
mpKcXDrHnFnrrqhFE+0s8ZAjY6GW7Vp7t1eTPNWs5oZ1ycK/BFLoDpd0rlc/HuFT
YvxhbY+gQ3S10MZvT3IHH1pKVMEs3hlv6b38WE4dg5VWFbkYs1lEuAvVtGN6yaGK
Sv23t1yfTGqzpLVBUIXTUBDHPulVeJK2f0zBdP6vIdDMngiUNFZ0FTmQtEKevVN8
xFrfBCRNMZcJ73JXiFsbjoBlX7yG2p4jd5tgL7x1DMXRjgY1CzckY7LQjo03m7oH
UPq0PWmM2C7QwkHjDG9eXpSrPT53USHxO7j2V4Cd1UygHg2W86t0envKu3aRVuhf
EwYaSlXcBryzJHmR6VniK9BlKB7E3z6XZzQMSgBFWoLUxOHWEKekXW5RZr+NKZNI
SR4YjM/eC4JZBAugkZBuqU6xuZln1zg9NMjfLv7By51WN1creLL3VgE63ViLvBOJ
8nVnG1hE6RgWd2vAm1IlTDr3nBmtg11k//RqpHkBxC202UkMIN2gRLRkB4oK1SaM
WxnpoTqV97HrkiCZNXivys+4/1tOXxCTJ86CUxt+B+LERtE5l3j1KumtPOk8a0ec
q0dGccJW1vI5qra3s9WVx6wY0rvJGSe1rTVeWBzACWB6AfACzYoXyc8uy96wRF19
4uNAdi2tX2hnaHNvyDxGZdtM2Ln5m57F+oF88t3w24mo3T50pncytYJj3vmxbHr+
MBJLW4qlsS9mOEGxcglEaJrdnsCCHt5F3j6BfeImBGfTFADzK1YevdR0S5fCpc7q
1h6oamN5Jej4iGbEVCZY3g2azwXExz81Ro7auV3dAZ9E1E/futpjmKd2h7QSXOCo
QmZo/O5PxHNXQyuHP+UU/luuZ5hpjISZ4umxF9dd/6gYkWSrmUjH6B4rQbihREgT
SkBqNjYKj5sMXE6oAT8KzzvFY9KwZUEG/8Df+Nz031bWesL0hxNFNmj5xqFVDjcx
f1qjHk6chmL/tsExOfmjNgvEetPFcGAWsfBJFaMumpa12MtBadIKQZBt/ztmcgx4
J1ndXRysP1xTGnR/88blVdlkzX7iC/5RmawLWTZAcypfj1ioRgKzK+s5nZ64RQaw
PtkPt4/5yn1DJNRr8UKVViP0MPxX6iIjjDJghJ4jRnQ0tth/gAaocaUbGglhmmkd
GB0UF//H18NDoQpxbiZFMrl10/Ulc0qxi5p5+iDiAer6gNy8OBS/61bUBchhBpoI
AcejA95+8LtYidubL/LIm17zlOate4FYwKpC9BLohLFh84qz9Ci/xMhWFJpTjZnC
mgt2IoegmhXyZT1fEu7zVsKNMBlaar+6YmXkgpZ4VlourVv0XPIi5kEB22zJlZeo
tPgprGbcsyAfg0xQ7uj+gB/bjLP3xc6HSmlZRwWpIcvL8u7TNG0KzlnD6VaDbmOj
ep0uzjlFmum4Sp05/bf8PDD5xWb/H8YlW9U7NhLrIfsOLP+j2i/JiEzEBQufiibd
4Cwp9dHux2Uet1OfjuhcxbfbLwvcu89DWpi9LQvOTIfsc/f6ubCbvAJeohLvxTt+
4gg5Hkz7du78jaF/SLrolY/cQbBecXIWhOmyRVxzYBH6N6UWX8B1ZHXVm3sjRe+u
6rIkWY6mhGI6foYAt5gxWYEKhQj8GHqurorq7bhsJLMCoeH9hW+MBHRgfazAFflS
pR1LL6JxaIafRYUVwh5mz4p0HZ/3C4KW2lxTYlBBmhRl2URtB8BAOWPWCo43NjdO
e/hq2omLex20nsJAkGJADNPiPjbVfzSap93IxIPa+xBkYuW/RfVZAo+HfejNHbG7
ylhso4yRV1VsKXejU46ryppEdzfECGu0T/2p96iXeCX7XWqRRKjdWwcL2EdPFOkH
LwVkyUH3USOgqyAaOIghjWsIC7oW7XDjDACibwc62SyV3+AgxT8isN0oGvkdMfOK
zcqFpy/6S3VFMzV9zzskHX/WSfuYF2lRbD2YDnJ/JniqNYf9ZPp4BL/poQXxrXsw
eJ0OHsEUncQVnJ8v2vyLMM1HLupJtuE0L7fwJ/tNcnidBaMnfPjUvTESPPxPCLUk
lY4mgXBZpm9lJMGrZvHvfSV74j30oPXP737AXmNjtFz8+Ax4KH6oNHTc0/M/QdUv
aIU+2PYFNkb5IeaZlR2mzHK5EHo69WHjRqZXTqTQf9Te6Jm0/DrlhlT5ujPyj1bG
w2RZykA9tKJBNr4bSOjbWt9pvi0fL1Ueun5CACrwosL8rm4Ly/iQ20Ao3h+cZ8ra
Gmoio9Be5B5RkCCzRIu4Vq69p/c9uHSoiLP4OSxr0MsIgQH5/vqjHucjGJq/bk7q
BXJH+juO5dxOUpQlTPClKJGwdAmO3Qu3Cu4CfD5ZIAe8W/QPa4Jg8NWCVkNLyD8y
SkqLStMKxpxj3YB+UBoy5oymBqUpSLA5w2F7q3l7xYCH4hIU2KM2zgZEfHB4PZcq
8UM7rznBYnT7wjyHdd+sEh0lZKrrAxwhX75Jno4aCSWZVFY5xYRazQwJiOl1WduY
eW0AhyvmOpNp+N7CILZWozHrYArewkKzslL8MWBn2H3wd2gIocIP6ZF7sgnyO8Fj
FUEwew1spu42atXrax3wm/8yF0UbkAD05N2TXQIAmhTEcFXDxU1gPq2/Bvl4V/WH
urp+62fOD0dXsu7+/QehhBtdoAysnPZxzedLx5VrH6P2ceMn452DTnw75DHXMTjk
qIAd+PTi6Deap8TbaivZyT0+IQbtUhKcFnyT0OF/sahwixVwqX6EbZQspqim9KCV
vPhPF4uTcif5glqhvvKJV9HygaPT/Tu5rhTc2pCjQ1mt+rDDo9099xRZlfR2phqC
vIOCKQYcxHOyAU+ZkaExP5Qp3l3oO/6hmhQ7GjoF8Yhdqxe2iKPm8iqHiCE3nna7
tf++SByuJNBrMLdnF+yidCMJEco1FrfgcidVeztvYKGZGEyK97b3FKv42iGfkP6W
+9HkOII2Eae2m01Kifeep0J/0TFJ9p5NP9nPOPrWxILsRs6zXeNd0jI0V2MhVRN2
/OpU/T+DnBIUPwFJ0Q58zsViUx8GZrcLMOcP8CfsnvuIsgYEFNIaLPZR9pW5NIIr
QUbBYVSHJPmWiqXLDLNTnvnejMmwlF7TAbA60jt0WVFfWwqYzGARAj4dwmutR3Yd
f8lRqhKg1jg3eeIKVxZzpI6IR/UMSCv18R9yP78BHXbpuGHyw5MlUQ++DVz3u/W2
t3moqO7fYfXeAB3UzfAEBw8hmtr0w+qQ37/Vw86lFyFZG7O/7ryvSA+P33ZBDn9Z
mt18wngJb4/iiMGpf4BWq3CGYqC6WyZI+vF21XNfQfw3jOD+rlqhnIkewqpGj6QU
74wZSk6fPYIALBHS3jYRKxNZNgvoNlitsz7A42vTkESOZLO/sSVi1Zx7PrYiCXUc
/yl//bH1zxNggmo8B6Gs+Q+3I4010K/Oof4udNI2ZfgXE6pV0X3j/ItzMxKNIYyq
E6u1ENVA5+eR1MPRXgxIEg8b/v/4Co06wdm5fC3ZRpsbYgdHDf4WuRGBAmHq7sBK
8gvnyOj0kvmASetjHWCcxnZFCkTEoMnUZTPe/OmZ0/TereKNJbdZNOdO7uQvZuOZ
Pyg2l3AlYXahbuu46Fv2Qc6pix7uXUq8U21iABAi3tFz23f08CUdymgI1ESH4aG+
EvgzJbQqI2pejKsmxYGsBRoLYQI3ueecmbrEFJgXh01LtotgrPPgnTFUg2NUSGRN
qI5GcijUzC6eLIKlqTyL+jgoc0DLPv4A+15s1P8zfIHF34B4Q/5goLU59boJaZhH
Hg9nUoRg3vSqHvdwHT8nzaAZlg2ZRl49gt904dUw8EF4f4U8gi3VVr+q6+t5UF+R
fN80QinLL+Al78i6XYE2CuLZwFPPYz+cS4lOIYCyNMwpNIocYrElLqwu980bEtWG
Jh6bOOef4/OfKccaqY+gLxkNxUr4e9YCTG2LPtXPF4Hkm2d9hBQFBeDLHZog4KCt
O4TnMYXxN+SOFLCXFU8H+6jfJx1U9k/nJyNxUuW9hADsk/rN30lw9Onl1cFCDhk4
mPc3SN2+upQF/jrkGw7oHbVelM7ZkY0JATbVTn792mXFA5fcf2FM2PVCbb3oyHCw
qH4PbFP3t2wHqMUigcy0zGCMRu2Rxg9aKCo6Ca5M52YCrJQTj4Gfst/XW+RjvwWm
zngYi1ErweWcjQcDqlmy2htMv3mpqZxmnAyvtdsp2RkdvI9NiK/QgqkA0Yw02SWb
0jn65UxTggKj5a1Uy7J9RypmricRDX+l6RP4emNPE2UxOsxxlfvCkd3ZsNKov06L
d7dFqXB+6xtZVKFFtwCdJ4yqzMhJpA+7pMxb1HngeohK//8qKRs1244iTcHawdbm
rZhBSTZWUDi2EMm2oMHHEvctEMUDfHMP24Sk6X8EI6Y1li8YVqnAQMDiwWBh41w8
pZvnLKe/dp3E5Jmd4t4KLnsOc8SaoGN3azYHd1syE49XWWHdGOD+o4JXNpNShBU6
fVceE7pzcQ8A65jYkuxqLtQJguI4UlX+HzgWcRkzRPctOI512CP67eYazeh6iCrG
KaL0vqq7cTfsV8c8KAdHDMSu00Kd6tMQTIbY8Xnr5/Ng/UKFOPlo5+hsQjL20Eji
RtIOYkf3csaJd7+otOwXbydm4tQuP3Zvlx6AbtHofEww3va22CRTYHTl1ikUW9D+
XGBoFZzsRCGfzVLhfo8HFEXuFAZqdyWqlv3QDtXe5atwRwverytXrmhh0I6+nQtl
87eQukiYs+lw1AkfXAzyAA/OkvKJj+th7rkEmhZU7OOiAcL/FaPhyy2mQUr1lDWv
uSexGz7T5Z3BDEP0gFj50foGhF3riH3IwHuDAwLVupYfuqckc+9Lzb/WocrE6m4T
Ao66hwb/uFjI64vfo2Kqea8AqKdxEeal9YHo31t0LXiAoqT0L8xivx9TarMqccYK
3T295R2ckbU43WbJx+3dN0FZy0uu10d2lMrCyua71GYL4nJiYwudkDmSQ9Z58+86
uJuQerGXanqug0EECrcYAdiYPyiE7XaXJ/nFNzxJ3BnUtHMIN0d0GVDnFONJafjr
JdYTEAZx9Xl73dMN5b1vkh9bFpr5dEzx4zC0qkwglfAWyW2P4JmNIaD2x9iNJ8qb
hiLNftL1eEPpcmPD+654VePf5E2dUPvVEKGFyPhKjphJ5EU+UX1RVWn4jR1nHCtV
2aBEcCjQH+WMXWdHy5/eTY8UAx6wxtYAry1cQbEJ1Wpobg2bz+fb3trP3dEo9SQN
AquLLzlawkabB+I5re/FzgVaV/Rj/lGFXszZcS2vqs8ouXLk4xkchtu5vBjsRj4H
RyVD4EpkwJHZS61QwdXfbeCDjngzUZ261WrgeIJnW8PnKUcey2KE07XpWZKVLezT
/029D+1nk6yljuS/UkIUjiWsWzACAxj96VOtLGgHZdruxC2mwtFt1ochRTaG1ccx
PuDNqJSQj7Ij60Lg/9+LWnfvlveLyjXmGe3hJq3pz8JCpV+YcLJ0PUuhDjM2zS1g
iNXP/ATLRkQ9YGBX55VDoU8/todgI+SxuGBpuSFsxn/vavPoOZxe2V9myiH45U5A
0t8EVFPt+NBwBqULrR1FNs+9Zmw0GYmK1uT4qdnzVLzi/HZNiN+W/z0UHOG+3y8K
FptHCZdTNDQbA3ku8kteiGLksCOUoYvVydZWgSrSWj1BlglmDe+SLKdXBam5cg66
ATR275e+KHzB2wBFO578DYzy8iaGIPk48Q60gyoJwXfWDBUq2YijI4aXGUsgxGyx
htBA6XWRekVVTNJDQEII4Dsp1N9CX9gFSKsghtj06o5GELWtQegFM3e99wZvu+aD
LGpFZolu7Tl+R2H2gqgJbt2KCjewrvNMHumVTNG5gVgkJKs+CVFjwf//k12bjzVj
hBtOVigG2/JkPu2xdyQwTQfwTgjgFN7NwVCqwDKMdbgC6euElJRbsmKDiWSZ8pXa
0n3tad2wKDIpGvQjh+olhu/nTICPBpIShK9+efhbxFPd+thjn4cJOQ3ITCVKS5Dw
3GkdDSks0I/kX68KGfQ9vIsLR/ly/ZdJb9HY8fvDEe0D9MHTwM0CLJYRiJBDQ7G/
E1ZNIe6cD8AuU0AqISp/XchU9uoweXLX2zLiBbQksLbbzSf86EmIosl6xLTFFwP7
LAWsULlBT6jOVVqQTSYHZxYdzlmQqMWhqobxJKEB3uCNP/5FHny7GDzuFwADEExB
1RQ/JoU/Edg1zpIEChTPrBf6h9lq5DCPfTsi3ceuU0R58k899aSKSrqv9SXB3eUP
IMYK7FP1rqlBkU70QUSlGdgvZZc45YBPiE/7Mf2icvSBzE/2tdYWfkgRnkei2AVU
U+fVTtMynIjgpsc8vN7ix8L3ToDcESkWB+he+4PoZnd0yZWDzyh/MU784NZ+vkNe
AIkqaSadesU2VlWpEhHZtsBzrwoSBImeLPfc7ZiCl0vcT+SDR1yjPtUMpp0GswTK
QzzU77ZlMOqvgPmSbdDMjjQ9/SAfhl3L8aziAFlVSFuoxFMKehMzbcfsqu9ndYVA
SZHSvlJXfryLXYxvWDbYoqF5njFlMyLYMtTcaaX/GHnBjo5/fgYYWwKKbAVNQufH
SRh/hd5MOFpMjdoUBhf72HTVXoRzpBxA4r8XdFyhD3V68rTk1ixJX309m/r446no
uF1leZjhpsK7DbhR9Wyzt7mF9aKp9OJraYBO8S0JUgAEZTG2SrXuSL7/2Q/jOeYS
SbPT9xA0IKX/87ksw4hNqvfnqgNhCV/RpfO1/WOMPpVnmGk6pSLLMAnyybZI3bwf
ylRbldpNrm3x/DGrzhl6uj+hO5QQyDcImx8noDF+1fJuHcPSkubSmZFvlLsytue/
qh/93qXv42pyI65I56ShjHmcFUmlQ/FkQZgaPdLlkuqFbT8sni65xJ9t/rd/XZyT
ssjI0jAJGKp38pMOyA66lLPq3P82BO5lvX5yepxANNM2yAZeCXI/tLTnKe6VXfIH
U5p64iupZQBlydY8fJHLqdi+I97wiBGWv8nmd3NXthccNBjjKOoWRqOSTiOSMQsL
PXbM4V1R5GFzjFM1xt7ckMw28uWrY7e2IDzavBlDRg6Rpi0a8N11PE7QMHE07h8x
jAmI6x+9PFrSHYsqSBB2H6cwUdBwJT5cLS4PDhvNLz/dFDuYPfz99IP67o/agpi9
J8+bfKMDDStlKBblRF1bH5/PucxbikE7OWWJNsRHsj/3XA9GN6QBd8m6XqpniGcQ
9QL4BrOeD+Vq4E455miXwj2SOwV9tZnocd1GZe1MKzcGSTl64573OZWgARPPiEdE
kxA7dQe0TxdJGjykz8CefrGJWPjPqKogLrCfLrseCw7OQUtBUhZL0TaZAVBYX0t5
IkFp589Y3+HRIbJ6T3VCN/o6l+IiV45Na0a1KLYURLUZczVGAMxYFEw2chBeBogX
TsfXQZj9z3hVBqROFRMHiitHv9c+bNvvsUcSYNAyYH0Fhc+RqwBBYBjB63OMPg/n
zNdVA9DgwIfavCsuiary6MC9oI6sOYizc2qRmMB9aWc3CN63+9dRtH04m4AG7VOC
j5XOamcOCS7r8SSl/+ZH8qVpLBfkP95X25nN3E3pIvHXX+OrkJfEKtAW6UOwUZem
bwziCQ3RnYrFdC+iKiudUpLOwbIOtybQcGOuunIbKhpc+5azA029KN33dp6uM7Fn
jkYNk4+XNpl/2tcTyqBJ8HVl+ggb9gUEbzbi3Y5qVoV1n4ll2k8MstJHLn6g92L4
nG4kpBhGYaFV/4Vdd95bbzjK7+JGiZsX2cBV1Dc6CFK1tp0YiuO0HSJ96QJWKMuF
4uC1esAk3MP50tcU9Y9EGhrQ6utEq5HDC3GuzfGgtlV5YFlok6VfZ1LWLbxbNAQV
0iCRXyT4/DK+u+POlMm47AMt1rayQi0lapEJgpJ+DgXQbkw0aDfFYz78ITOepqvO
eAKzRX4gkGGGDw9jtPjb+0j1GIbrot26V+BeUTaRNARuSt5FVlDChdh3JoE7/qR/
X+m9Y4mev/mqzQzrjeqGU/CYAWmDlHIcmUppmX3oFgv/nVDFZ+mR2Pz9yHEiGByh
5uawygrSCn6j/Zlwl6heExhF6568ogNsSiw+Y4PHCSuzX3KI5wGhLZtN2dnGuKi8
DzIQDsEq7BeOH6dDNhRQ/M4bNDnTFRZwDTNgKH4VIgY/l+ccgPC0GQTc06Y5hZAQ
wKPrzaDv12hGcZWqjuhwKcbge4BzTewIgoCSxOipIv+ZFFtXIT0Px231FzjJgtVd
JXBumqIFV+9j45nWcDS7FnoXIDgcLvt+LLHfE3Mmbku8YC6kM/skU1WU9hkIzK1R
3uKGAiT3cHmiz+BvuJ8ZxJzAxxX2iI9yi81pksrw5nsY5Jz7oHTMRpUQuTo0s8SK
cAq/s786Q52Nc49OHVqA8HALrK02e1GNdkWx/SEZtlbOHiNqxTaApXrNar5I+4Si
4UDOW6KskVoX7T0tZS16qHzCgr7TGZbDteVIAL1Q1Pm2y56AlBFvNG2xpI/YWyQq
K3kWaZxoqXgPvBDf/gGNo5WeKBLA1hw5S+DwYChgNUX6XK4VX2P9jDQx9FiH3Xfg
R+iOrz9+MLGWvgR66msE03espigJE88V0bETqTQwN5xU4kaqblFCH9gV3dFnIyPF
ic1y2S3CUqydQ188OyVXNcOxpMuHu69zXIpY1M/nDaSX1SVYtxUKE64mCGPXd993
ui/7hxwV5LuFXe7nj2X8fvVQV1lMZXA9bIcfMoauMVbaUTcflq7k8Z+R/fMcDdpu
54f+aRh833o6WV00/Aue9UwYH9/WWebHcT6ARyx4ZZvxKh8YBGGT6O1GIvZdMmHi
FiVplzPCJTQoQvCHDaK1Qh+k2RFedBqSO9xm4uNT7Es+0Ie6nrdbHLIP7RxShDV3
fB4fR9/BmCe3EQHtYepiWE6n+0qcHTuBT6TPNzlAywO86V9v/XK6QFRWUX/V/veS
SZE6jNIbZLlKy4TOmpubSD0Q+6sYwbojj36k8R6l/gjWAmRWxLIncXx+KQUIMqNX
s5eBiZtdAJZQWB1jK39W5ov5DJr9tJYArRrTF+s8rpJF3rLbxX6siqIN7+uYeHhy
75lvCtqC1pXqYr9/Yu9jO75pmPorTg4qoWw0Io1Sb1nae66hvJOT9ArvvClRKfOm
ILtOcgPeV7eoyznuBCgn3cCpfibIkcAPplYXZZ+HOWKqcgVtvnMg5WLioZejHU1j
CpJLqaRjlA1mjBPCbRml2u6t6oP5ALBg/z8SaM5F9FVCusWe7Vz8D5zYUorU6+cJ
cDn3U5oq9dM0vjL8TDjxMjq3b9giOQ++ZC9oFFFyZvYJ/vHtBSUMLvM4hEDYWt9h
RNmU4Y3T7Htjn4IiV+0RzfHGST75wWFo9Df5r2GA47JoqEIGQoOdDwVGurVcTEHA
4jyyGy0rEbUxQt28XvJKgzkv9W9CvSQ8k6Bkv4mX7er3qKbtud7NR+B0G5qCv1ps
4v1tx8xVv69n6w0ayN0v9zrLmyWcUAkP4ZEKAGZp47xWzK8VmovbTTWulWK5tgJv
O9qWmZQ2zEBzqh++OVT+uPGEwiP6wXRZc/wvddY/Nwuc6ALDWLoTxEbaq74a+Qfk
xII0GaUCiAD45nT36t9/rse7R60b/GA6ueBTSPkGxOBbBXcqDWeLRGYWxiwruNn4
Z1LYnEAbWrUKCuksKvxN6hGv1eWYE2hpapBIbSd50eFc4uElwKFIQ12APafL8GhG
ssioFHnIC82KQ7nheIZH37VA0+uUorS3vY28UjjyZKwoTiMG6vQZAHc9KOA4vHhq
G21EqyQhTVfvDJhyfP08DQGP9zZ6Yl1KCfmxxHPm7GyDjjwnrrVVZPpiK48PBCsp
f1ne306j8MLu88sX9Tk3AOs5UFkFGp9/KV9bf9ZJ/bOIVYk7IMvSzxRm18GyW6bB
YXQalLp+2ScqMRq6rfGPOD+JqYJdrfu/qnKsCyaSe5kJndjbe7zVYEZPuOGQIbUW
MoF/oSMS5NVeIWOvmE7D+PT4PQzNK47vvvnXB39VknPA29x4Yxx8tfBFCLX03IrH
zFyEa0Qa1jqsGoMrygDyEgG8L+sMMk/IXdAzqCxfxXniFS/KtIvwkHl6CVBdW5Jc
v9FrTZ4+mjKU3S2/zWoStvugqxkbDoUrYpczNg5GcSarvg418cDqz3DvRqlbzRC2
CEJmufXUp40b5Gg9Vjbh+uaf5RgE36whEH/Wc7WxLBUJHtKeG4pjNeoF61G3d/ZL
oiLLFJ5Z95ZcFImcIG+94nyixcz7HgNnMZe8pnqXu4diZ6VxMy0OAuI7son0uMfB
/y9JN5hxo0CI9EQs+7tm+kkEMl5cTt4KAugIkrnzAoMWEsaRUyUutMCyhvXJeQe+
HQLE/YI6f2Q398l7p0NNAqDKe4PQY6tZxBXQKAHgoUSvVoVFN140nktLaFdjTCeo
Kal5TcU7hW7olfYhMpYzDG6yZFNcLHGK3FcVYXQJTkfHZ1szKQuUHkRwMO9W2UxD
ykGgDrVPDsfDn8ITVrjdsZ4UplUDEk/1SCMVSsCLh+3CJTmDSQ2j6F7wLMCDarUz
jROYgqYhh9mEml7FwhVa852jDck2NU6OsAY1mxZ7345BumCHN5RyYF/qWYePIMk0
mclP64XMhbW4FJ4xK+HTIsg40sGArBgcltmOoUat/m6mBpbVyZn3kqu7D5XhTreJ
LiUdcyAmcMAfmM/dA1qPgGMmqyhzooxqipXqLilZO2pwTYdf3OMiHYM5nNTaUVhB
zEihYLzeiDZ7uBnM9zBcbzXqEb06kCrvN+Ubw/LveaTsIM1ih7gAmxBALZE2sYz4
Soz8B5XqBttmIEog2B08Y5DSHTKQgunIQBoxg7TPMunaYPUy1roaXaAqUzhaGsfd
55o51lir5FIpuAj6V0pdZ4y0viQZGUmpDgNzY6A08VmkIv0IJX92AceEcYqmTFZM
pr5rW5PcmU8rFIS46r/MEYpllwj7FbjN38wDkL5s1Hftap0kCiEc1phmWismQmgE
mOR5MHu6I7wfiGU4i9isBjBehjKcx6CpiceTNDd1nzFV+XM2R9egAIn3dDJjIJpP
4OZLm6xqq2QNLZ0PpxnHB6VE2xA27KT1JHdXufFrDsytsg8ZYpqfyc3ZeQD2LyJ4
7ch32qx96juP85xme/WQ6C2E0uJrZIUuM1423NuYlRg8X45ZqooFBkZhjxZ300Uh
TA6sXFWdtObhfRyILSJqtyGxt20LNUO2ZOBP8LGYDBYe0tSrYbmlTgIuNd9LDS2a
drb+gWuUuXtohyXC/zsbSnKrJV5c/1U2PgkHbCFpfTj8MvNfIQL+iwJlH5buHdvI
JheHKPLI+ae51UCDGpj0LpPz3MF72bE/rZiaSm4x7VCfE41LNKbRRLm+ijDD/nJD
J2bbpGeuoAxronGv5mnZhaMUZxB4LEEUO9ubQQgKGEWhNJqrXqEmHED7thcHrWLj
gfdwFNSfhLA+ylCg/DnrZrwqgWMLnmzW0jVh1pWL7AjV/Tt3ArHSWQ0pS+xifrlK
qtvdO+eO2S5Gf8WyWFuTZxb++Qd+Saesgh6/DzjlVz3l/WCsFE0jZrFR/73AYG6n
j3EJ+BOXnXoDI/XQOx6BIkvZAP1NtuuUbSqjAWx/jtqUo0i1r4OlZ8YRWi6tnBXF
lZTAPKjHKY2r6UlrHAULzXiZqkwCOyTLwSCWwhHzL4/2EVyO9EVLBoKhsiMetqqW
pzGsq/3voBurfx6D6F3keXaBWF8U6ZCYwIJMRq9ri1auU52xtiPIOYyYv9FD7wzY
Nhw5WbPrQ5e+DdCrNqSRYUvnekCgt8u0mP7mWKgMfUWcMV7g+DxPa3JgXa8Ltr5B
YlIrowEEuO5A9b5ZUdSWzbwZKYAD3OIjQttFBG1nvOjkrwhBrZaVqw8ru+HlBFbg
62KahyhK79wtmZcC6E0ggDNE6axCDFh2DXlVndaSsv2NrKaf8f8XBBlz6oSLrujI
mrpAN5WoaDHrpdns9XznFoN2LXnQgTpFx+1Lz3PBM10V7O6CHB9lAPc7QPOCDRP6
LWNP/k1N4X3LCuqqoYyEUOPczarJb2pGTB4wtj4U17Z0lcyBw0MyiVf4WF+JgRSh
YolG8Dm0qJAHWa2joTpi+U5E1Mmm/tPiskqF5bE74OIiQ97Ak98HTNo0cj2VeWql
eZkImQFkqX2Tzm04qs8NAFPgl6/vycRa7NdViwiHnvlMB8CbAL7zC+mh25FOSNZg
/YF9Q07DeTXlXqZfoK0f6XKaWsdscv8JQGAsZgwHpPTCxBB3TBHgOnpq3f6C92uf
CKIc6iQC4sBHOLUwShUXgT7Zr5K4qml6eKD3bpfqhbu/qZMGL2dN9y/z1pJ/48wm
H8+JgA3UqvkgmzA/rxHaXeQ+ROBF5VdRjz/8axlYfvIoip4XL+srVzoSIe1tvDr9
DkV86FbrIiiC0XoeAYDdSH74R7704ISUccltP7XVRKraLqD9rdolX0BEw561oyko
cBP7ye629eRo4XeGaR0A5ZTsB5zTHFxfX9xkbUzPa3rl4JcrMYKrxsZckQ3ur1X0
6fYLZe/RAMExRmPlzyYm4QC7KiP2EsIrCz0oxp93Ojmb6fie3RbbUJjqG2VwCjXc
osc2BYLGg7+1cBogC4IXUKd7tJxwBYtqDLXbUYi9fwwwGJZHpeyIiuWbjR7nxJHz
msfl0b6YwxJgilaxQqvkM9VZl7uHWjnyaMwS/yXek59BgXGlX+WYghp2yATOCshD
DxR9D+79Kg1fpoTrVz/RCpkkdvvi+G+FI+3/kVvOseUuPRYiAabAW4V/Uun5ybF7
wfLDKJczi7g9QEb9fTFvURC7fIIhdEsEFHUPd2u5hCTm6fGuUiAGmcl9vlJtK9da
fGAnTCnCnk+IiLr+4Bde/GjNdooBO3vfLb5pipxzwdbPPDI7VSq7I9kV/D2bcrQt
5lCbbVxA+pudo9umTF7MzOVGPCF6trb9cNiiPeJMF+RilP5121qY8lyALCHVPWEQ
/IPIHNx7j7kd1oooRHZj92q4KbUhyajizQvHSYUHpQj4ZNwSC37qVEkGT6KDidDV
pxGRnVRaRtSDL6bTB1ggf5GOWsqcVIX63CfVP2uy3ryXdCNxyQOhCIrFu5Xs30E0
ebf6jTg1MIOtVzL0AJeMrBi4EyEe4LpobnB0ukSe1vlKMBZrlCQ0PZPVSEZ64MQD
faMe/QR+4sdKzMVgsQ8Vje2gyfxLT+V9pfqXB+BXuIZJlv2YUxCHPnPGL7FBo3kL
kp7FXWdfm4ukhLluR6eIFR2LTqmDpLm9jN8kji6LZOhPamgAvVRJeF/bbv3jfo/W
FWla7xSfw/anLixkQ3nPjdu+n5d61y/D+squpgW2qSArYijTJCCkal4Vkj/6g3iW
7L8equlaLbP3NHS7VGkt9dbFVby8m07/h9Lz9fm7cWDz5QchmyAsxiBEhp7sj8P3
RaEjMsrxTk60X7knZytsB2qyiQXZAiEoLH8yzD8SLjzuiLU8PpTbSMlx9Z3MGe2d
abhaQLx0Q46hAkSkqvkjybcCeRGf6gLqZxjKKbRooV7FCKn3rlkp5BNHy0E1XuMt
a5e7Smi6AtyekstgF5uuU8P6J+MN5CA5VL8xZUXEZQ5LZHRlm9w2xsmZ0V1qM2Vh
XujGvf/+8X55VuQmMPdFvK244A9YwqUKcyUULBzeJTwwpVGxr2L9gprn8gijSxBF
ZUv8H2lXeUZgh02lgzwTmra1l614IqT2tGH8GvktJEtkuLG9jV4tvSqnW46L8Qc+
lmofrvdFVw1wIO0lGyS4IiKlfP6JTfDl4FlkEEHH1DslNBQG4+OJbhcUo++IO4Te
VFtv7jhs+JqkVLrOAK7SY7mRdP3033kdeicc7fOrp52o3/Pb95T37vICX0ifkedt
GFa0V1VI8XLvdiUYwH9aVr589BEZs/SbEYCmXnUQaUn8rDtKKO62OAQMxQofui1b
KQzo2G7I0tmEwoUkepDdXwWJ3sT9Jfu54NgkoRHYs6Yj0nIi7EzuqZkJ6fO42X8D
DqvdUSTG0WgSa/CJ2KTCp9mf153si1LaKQWVPlAdiouaaKY6gw17k7ISg2UvSV9Z
s65rXB1Z9ZAKEHeqrvoTU86SnYwOB76NZ/lXmmURB9WFYzEDzUP1sxuWFuqufKZi
lg1pnDkpBDEzg0YKgIUHWY3xSJlM8hAnTWaQuwktUxfRiFfEehLDyl+INfTrilpp
GFPgeWPYESUhYqOmYs6pEgTgVahYs+CDZDxpivkoOJd5EOYvYZ+4uJChxvr/X7sK
WtDnYTfBs9gSbLZtDEHoujYJhxBEWq6CLjQL2jgAGjVumJBvwyz+6BEoTIVjw2do
j4yQhEnN5IlVH9s2uHyPkntvNWG+6amFo6QXD21T+Th8w8omI+zUuMe34mSABVTE
CA8QzGBeuEKSYStPo/idXBZTZn+vZv1BAiGAleJ/o4lkBLW6lcOX9U7VVxNcV7qJ
/bUPdJBaV7fxAGMs+PnMruxPAv13ORx5oof1f2ecz11oi9aXupoPgSZsXAyWDpdE
bTL2Gj5diZPqSdagz5XX8Lt+xHW4xlXQ7QnIyXsi6H1ETnaafYrTygTBA337Bola
4X7z7Wl2J/KKsfE3u5gBJu9QVJXHUPo3Ep+UT6UZUFBZzUqug4GmlW6dsn1DRN+4
mo4EQh7yK6ubFQPEmffC2OBPFIl2bNDNQgbsnDNstBuBGgTelYUdUpVpB02pM4wI
35XFhUST+hqtYEaytQxfvHaceMhzINCBmyxj2nOc7nqVwnltATrskH4zo9Vfx0MP
Zf0sW1vHTqFppYKikLwffldKf3NaiXIjvWkeQLSa/mO34a6cJ+LTzxsJsMu/eP/r
DZV0RbulcYxEDxilZe9biIKSbMtbtIEwRiLmG7jCgPDUY7OqSBMfQZgk5D6pNErB
dWnm284m8QTSwtgTtNzjn7SP+o03k49Kh0d0eMB+83X0xaz0Nbaq3TE7/0y9Ps2P
DJs751IbzQax+g8RrnjyKe3lWY1fMrtvbhiDHDbXBNmb+TVhhS8uEPvLSTgmC1KN
i1Wi0Z1bfqXz0qfVhMfJwVPB4QpxEsGhpR8b3TjzOqsQxy0sHLhkJ+ZfkVBLMvp1
tC8TQK6lYOLidlzHwShem9QrlEwFgH7kQTc4hBhKCGgosXvMG71HRaho2yGWYR1Z
wTR3QHGJD2dkJxm/VZkBzBBK6j6e0RMOZiW2AVlKaRs0uU2NEmmp4uGbeQu3VmY2
CoOv88zgK/eOx3lAr1Vefcb2hZr2t1/n/ic/z4O6mrHxvGcRqZgD90KiPcVqsjWK
Rt/dGKcb5n6xwenj22BZMp729ER+SmH5m8QMeiaiXJeCB6zmaBkEE6UfXRBk/CgG
tm2JuA22sAe+Nl2V/eH/bx38Fn+ZMLEbaBhEJj0s61RVEh6igFwcilMFhP8dyNOD
KeOnphBchpe8IQAMsUW2BrEK5OK7df+3+etiwqqHmSN0L5/Basw2FlOnoMUtxVBO
lLWlfC7MHmOMLuMMyAaPrrSiRq7z9RW7pHpH1Oxd/g7+r7ZJTUwkf0fymKBwhQxm
X71vMC4KMhKma7XKl/4979rdseDMwPi1T1eZioJhM1bJHD0NwCNJtjqERPmKG+L+
6pfeZPDuUHOdr9d7vq2QYH5qHRV4UdZEw75eaKjUZOGQHKl72MjI47p7AsiY16qn
AESWnpz+teOJw6a6USigYctbW7p9xrWC2NNa+pvj7aEJLv2CoIk3hoqUmA62Ke6m
rgaQUtWiGq5dm17Vjyl38yvjFzS29vQ7lg1J55ufEUD3Zk7Jpu7GzHoBMtLyHk+v
lwohLdZTP+4ocndM/n+Z7c09F4YG9TZi3WBjt/QDoKxv3SImhP8egEhTZhJijhOd
IgPchZe1cu28Dw7gntnZfTpQJ7wuC9tp4LAWbWqMXPK1EJM2yjGBAqX9+SVghAy8
WT4ycA/sb2ep0oIqEFfmINGcSYQYJR2k8SXzwlRTn3hRbJQ3FPToqkji+e5NCJkR
8tkBDN1PenTDkivHS45hYMbMKq5IHRKl38ihaaw0OVbre2FfCcUhXeICFi8n0KvN
5e7g1inEa4cps+vmzsKSlH6GVmXPjEWgemB5xXtpScg7UKzqTQ4g8Z5IhkGmviTQ
J1DkL9tIfeLLDoRmxMyaRCQbdgwvybL9YRblTY9iqz9zoKqoi+ZdfouiaOdxZkkQ
hLP3rtJ0lKCAbkv2xCBy/WdU91w9+RWaHRRAjZ8tW4hV1HxYT9gEbwbF75RBeGyi
hKxYleHKH4Th/jdT0Ahvv6giqBkA6LHniWXKigQN6VWcRudp+N2OVLvebz5xMMMs
2c7osQqH9Oz0zHIW0QqZ/5F5kI7HWmagZ5yJ64GyIGAIaL1eAtB2qNvoW6DpVXUi
3HDCsSJFapAqBw0KLNgzjztwSBDdxNdA370PNMUyGIY/Ek9g/qHlEa2IOLYkQvvR
Cx25eARiF9kITwJSPe0SoOxzNGIliiuLiABfFzKbtXSP8972nI1Kenlr/0UENfeR
mlhGHnmDWfJTMH5gUmtyGX8iSLba8pKPcHNPEm06JkyvObwRuPQYs5Kt3bYOtJh/
GVgZ26+rstD2JxlhQLlzDiNkdDYuopwQX5BEaFls1KUHPQwdZniPAgZWhJxKJInv
J1J9oMqeWIaqO6QwJCsSg+BZh9SnuKedOkJRt5+LD/hqH3YJBsyfnWSuuMDRJ3Jn
yO171vLqw1fNLNayaKrbEtTBTLacM3jw+khrJVC1ks5YucGJUaHRNJ/ybO4t7nlH
iUWXaLO40KZG3n4/fGsJ1cAk5AaqSj+fVtT4CauUockawhlyu5QQzlPbMoI88YQm
lpU4seTBPkezOg8OhhLtlEsC6sTyRZKHGxJ+L/ealZillovBLd6B0BB6XpGcKuMf
DDbPfcTue+H932j7iLzjQv6wgexYiVz5tbviovRm+MERV6zZO1oKmodK6xP8JeXP
gG2Hj1WljD6irxc5ODj9rjateiwDM1WOLlJ2b9tVzDOln/LJU0pBeOQzeHNsWbjc
8Gg1/xn3vI2dyCQh8f5ifA5tlumnkuIEFmYgN5wsjpdrxY5RAGJrkmnErATSmlSk
uN/MSIZBuEYJWmsyJ63MucJTyEW7ZTGBZ8H6NajTip4tws3oUnNvseKj0BUb7pG5
jdAxtsQ1iPZKtikuvfSBYaKI5F7F+gf0LTf/wg/MDO7DvytbOC3p88AagIpD2KYr
DMfXLPpNrh/0LMfbN+6xNldvBGUCqwEn4Sd1jGaowuWJuMGWJnSIIDMiqSkLZaIY
09Vh0LMeLKI4mn4wsLTiWHPIKV+kCJnxRfU8POUnrVrTyyCkpfrs8yIlBQYIfBGO
JrG/aCTaNPdEJdIekNnKZamnLUhjNVv3UFnD7sy8Co1+iBHLRWPlpX3hDvnKG8+n
67ayqctr0CMd/4MnuFEbeyowYBe1n4xL32YiwJrdu5oyMorDzQOjgYQ7Lj7KCkWo
wMrDl035LQqgtLuMLnEMEGyn+kpzcvMJS78k3B02Qrmb9X/qQguLs9CdKwsbYfpW
CIWRqZJw3wqnOH2950JRPDZEpjVBlARi2fu/BXLqsb4zR8X6JDJWG92pKwUrmCAP
cgWoX28IKQhzOpHRpptQwcCPV8NyRtYh0pGJl/uLVqYRyflJ8E2S28P53qN3g6xI
E8VkQ5gF2rUqkaug7kkMIkZ8jsUEduo7zonhNcZRd30Quvg45GIMlbQdmRLswMG+
ioBpr/biG+16O5SBHcea0smKwAJXewA8pq/YP6+AIM884iJKA/KNg76EUBn/DjP/
pWBU8WriYVgpAt+Eu3s32Fu0lCXCEM4D7nfvis4RSAKnh8RpSvEYAzTMIdIgBPTf
338MpHdwcxUM/iHgBEZ6GMFw6ki3WZv87wLob4lJryQkAL5p3S0lZkKqtFxBbAkO
n6/BrllciU7/rej1DKaA+/FF3ycu/BhGFKTeLkNyboUJSLBs0w3XGrF83D49hbbP
N65TJ77Pm/4AE32W1JHYYFuVqzeExMurNqU9nQblDf3Hz9yF1b0mKhGMQwA/G4A+
j4i3XaxKqkfyq5oHxUv1N1p+Cacz9IgccCTOK7yMhcts8eLIbbM3jr7TUtWZ7R7q
fiq+RHJsd+rWxYZT89wqixmAv4fe2KKWlgm6DfrmoFW14giYY2kyIz0FIfEFG+5W
qr4HX9fe4pS4TG6UnACsu9/dRLDapcosdRrksgmNh9vJjXkB4KJ/PzggFBnIJWse
ygRowsZNfIIDYN5HZfL2a0IKEXxHLw/4ENF0ezmBqBcLWhqRa042xTif8jn5qOqd
jCiRv4rS718u7vJF0ZdCDiQNU3WCYVkgDOWtV+cIUwGokPF25ncEpTnHRq6gR4w/
U3mMYMeOU0LF73zvTKq3YmLcq54mD7zuYlFK0z4MNHgWC7+Jmhim0R3njz/YEBCR
8fh8IFrlHjOD1wXOWwVUOp0fyfJzLqp1AOue/2g/zxmhA+RkB1Bx856xRk1/ePqb
WocFmAUOiAUpSIw9tXSDxkytkoeMnKWP2mpTZTecWKdnG8GIjs9MtUJXDX+Qha2V
ulUQfBpqsft8SYqyduhaD3npWWWYAWbkqsrWImNcU1HyI9jDl0VfeAh0tlpvS1TW
zwmxkiKqWXPD2rLjm5bEeiNcnFgnsDWHESHrdw0hPqG3nIZ64BdJNMjkmsR26akY
1BwPSA5Uq2WggTjLVqN5+0OiIt1rtqhvaTSYINBjOjpq/78FG6X/kMtaGFhdD0J3
by4iDt+Sb64qKUIPlvPqtReIFGxNhk+2nKzAFLpPZ4lQ3SeIsyEsPkQf3VtqaNiF
aEW5sIyzIijOcvVnwDsFQIEe8dVaSAv6Fy8nNl5GPyNzo8wYJLdwxKwCXuTtrf2L
SUrH18coP5muQUhlm5pkFCfb7IX79Gg2+nC7n1kpbc66A8V+KVXU1eVyTyGNJKve
MB0+ZK9uIwWLS6s8o/LOql4vp91jog2aSYRaB4arePN6AzYAxLU/4LonwSbhjT39
WckLVFO36X8d3c5cRNaHjwn1Hk7EnZ+yNYBx3bbDdWZwNr3Za/la2ccn5ATT3vJS
TVV8neKoq/CHrIKVZuy/BwiHYDaLp1X9TjLN1LJhRwudWJb/T5RD7RnaGZJ/po2R
nawO+6X3dsBsTN2Dk0NCcWROxxzZ5XhEBPz6BS8gCVJXCWb6Sr3EjrICSt+aLN2S
Wnpg7EG50rh9Fp2Kde1fpTD9uKuxFwHclihnIShM4Ej2/EnxDixbP4s3SPYU00Ng
lZK4a1Mo4cvNaixLf85FkHLu983buHkggfLcm9mQ0VLvnT675Q+tkRvlOv6Z42lu
P7EipnbUN92gjUJrmVWNaDxQ/ghYOmSx8m7it+vV0cW1u4rGCvzAZ9hLQhX5iUwL
CV7ABLUsVcJeTM5wQ+XEZptIPTuyXmNOEyaRt8u4EDIpF9i+q6RuFcoewHVd2jqs
LnVUXH1dy6YDEWc2jGUOw2plDyDaeuzX8VGLbbINfkkhmHXk8F9BecOVs1tjkMNz
/QqW1AXXuUBcZtGLwfzzXQeTfkZrLwZVwAWR4a8rLZ8QlN/4SFplw9te3jcjc69m
H7QoqTaVcOk+LDKiFQ1FShjFdBM958SXUMfTdjUmMOWbArARNfFUZb/pjL3DiTS+
dD8G16hMUtVqawFLkp+CMV5mMsiZImQmw4IRr/YeTzGfrG19Aud2NVgAHcsQmDd0
cZ9k01VG+o9lFlF68f8J0cY//CRsh5mauZtNnBgTjpuleKbgQkzq9DKpFN8Zo+2k
hFTxCFVNwC2UXXLkEyc+c/c31dCtN9aiU81ihgO7UTke/cFmEvfBNZTwGER9glNr
oesy5n1pmku20Wr9M+1rJcJlmpZVw8KA8FTBOG28QeAarpCQEA2pZzYo8T0KoGlH
YHi8YMM/caNRC+6MPzFOWFArx5RFtymHx71aU2xnWEGjCcmm9zdfdHOvVwPSs1EH
TcJNMx04korbw0kaPj919Ll+MzNPK4EUqK6S0IBLU8BL9ByI3ZPlkIBA44cSO+yE
nnadh+OsU8MbRaKpY1ZZmKdx7NR6pNF7OTfY/UoJCQIBgFkFIAaBGNcJfEQ6Jd/+
IOuoTka3to1V8br4RWwCzdWu5qcixpbNXqHp0UhtdH9WJ6u4FVw0gMsRTk03B9Z/
9+FOFus7N9JOda62HJwC6f0b2R78C5P9IawLdqoF+uPVeOuny9Q36OQxC9KVFQc6
DgxuLvL++sqxAuFZlKP2Esnwnjatr34w5vAhgfupjoNDB+VhTrF0zVnpFHKaefik
ja2Ln972dWZxWlXXLx7kPFb2GGgI9xTdv0fzFNxMvuaPpTs1T4FKbOdqcMSMzUxT
xd84T71iJD23ZuZW5jw7XMLCjxKtPrDE5QHRTpX3SZsCJaGCltd7V0/dXsDUwIyc
SOsWNVxu4PC9LzMM7gPH0xM3XPoR5akO2twh8QdDkP3XbT0Zet9Ap1rM6L5VbwI+
dGamHC8WDdYT8wZlliWanXvKQUowENc6/iN/5JMuuUxr5P9Tx+bsLX8y+4SYW4HW
2Qzn+ObnRjnkIwW9Qa3YgHyrdm3cD4ioCW456bK4z8Vdz8uvzyEigmvKKj5oeW9n
Bxgd8pTsGi1nA59aF8cJ+me/OFSwuUgdZIf3jcSVWAD60vnqynZ+xVKvfIejDWcI
OricjfoYgE6uBemRbDip2G05VC+/+dG1ZY8tZM8y55hCxoKwFFgqyviHzzosgJSz
pAAx8TsFMqWQBXdB8BcVRbQ3VPpZk+/ACq4ea/LiFefSe9g/5b4EHRKg/ymeOAge
pbkBzrkU8yNK0gkdPl627luxBl0SrTQdzGQQU3JtQhzSJPwUS5RKf0XjmKSGyl5R
6mmhjfM3dsZG8aBJdRG69K3OgjgvF8Z5pJx4tegUj+WwJXYA9pjySJrbgYpgMvX+
l8+96J1hc8YUS86pJFT+FoT5Kkpu39bnjIA+7QhS2u4FCdXwRwVexfFTW1Xw0JSu
MKrTiMfFQm7mWzOCtQT6oLySS6+CTBnP8yrcP8Pk7LRspBmj2BYV8KK8h+AadHd3
Ho0ctWKPTMAs5hAfKQbvX9pSUJjdCly/A2Zn5mQHFCbvy7d3GbMOCzFoCZoPaghf
uPaUfBKvefV2erjD0wakLEfGijKgkCDa8jl8ZQClRCjk4KWw/v4XK9fayw1+oHMd
V1d7eYJBX972a68VYgY65vFMH08cXwypYrxjFWBokoQ3BM4sHWnhCFWcRyM6Kcjn
Qu2nZg1vsIAmOPPWxnoK6GHwvOgzlKg6vOU2tbwmWTkK+SReq4KlzhbjGKKcRZbg
7HUUr+WPAtL5L0pb002KYLaCUzRc5R8Qkp/hWl+iTXuem/ytAAD6FuY1ne33bJYQ
fZzZRuH71L4k4HqQ7OwT29Ycdci27w2ng2Bk7u34Xh0HTYjHAzxXwgnr1LiD8+Ji
bnKPzFRuvAJn5qIVqDcwmZ0Da97C3Er3t1FqoKeyQgExKh52RRb6G8RN2aa2jmIk
zILqhaHOhy41jmDvRBcmL3qtI5AlNgxEC3rTQC3vnbfYabAEJxEmwEq0dGxqzAJl
RQb+4RU7/63th4tkvdnNNAHPYKMgYzW58VvuGH+86lN2CtIWgQ4PrtJn1by8CmEy
59hiT0TkD+rAFfcoAPlzWi8VC8W19cVs1Po71iH+aTWwM4YmB1Hpku7BcDbteJuI
i5pGGH2b/iv3wmD2Gw7zIy7VyztLmPWGs/XbC3u3goS1qawU144+CrVOWZCinqS4
T9dpfMVJqi+WoLNR4a1lU0TbfJK6ndOCVm+DSZALf82eLSVYh/Idu9OaACYbi877
/b8eXeIrNpHP8cEF+o5yHbyqX8CMzFLE7ClVch5Jzr1xLd1hJPSd0pMYwkUzsMj0
pQzu6GgbaPUSjUwQUzONhKXt2yhsw5r1Bzi1Sg0JIj53wcLNyxJEUjkylC1IHZU0
1Ii993SHRFwZIQeFraEOhPymmWu0eSj3jldHwrLJRo/qlS55PTlxkHzsRGJNfWGA
6/bgTf8wOm3Hn1MCMJN8H3CC6z1Yhvup3swMiyQBLYyL/k9xgT9CUrfb6/xx6tK1
wZ3L0TvPWejG3uR0okpl4WFF52cOzOWPRT1AVc6Bs/zSid5MkEjumXAJkVEg1Pbk
l6DiCLsTt2W1qSNIhwHNxdRnsduiQMeJrHkBaPrXH4ml12OWpu1iCqeo8+jZ03oD
zQd0yl3oAmzXEFdfc7TmYfTIPG9UXjv5+mtLgEpWB8PmfG187jqjUVGiYgRYvbCh
seHc2kpnoPqu97+GnUMz5foJCy4glyxxxH12t37FLYbrOjSsBe3kusUlXIqRMqff
08Sdf94QZxqBMrQWlROgd1uWX4lV0mxwHhd8qiYF5w5gx/9w7t4fC+MJ9B14M5Y0
nN+bDPQ5qjd/tV/pX0IhZvoxkrwV0ZqUIuJal6DRsep2Hn4EVCnI6VAL1CXrbSXk
JwzobZevAl2ty9Q374ftEcCu2m0jIEtO8x5D1LADZVOilf7QWLr0Y0cmKz6eZHoD
Vu+2yXoDjSwfQWYBHEAwyLMh/IRRlAYe3TR/RPAnj0doytydwgyHptFFyIDlNmbV
hf3VnOi03Nygz13KeqrlrLbBDRv/zcoFT0nPx322Recb+hq/FoCTEsy9sJQNYNQI
RR/p4VZzJNy4W+jUPbHl67F5nkWl8A5HCQu54Ig4SIHokmljdPh2OFPOpbcuVyaP
Ywo/qvd+VQnRzdHkRJSOc8K2r1CPTT74Jb6rOThj5XJsbmcqmUV5Sp+HseI9iLAz
Z9zxUCg91r1u0MT45b6yta1PYOAHi9egOwuoBl2sBfHrGEEdb37sPBF+JmhFK7mH
BGVnoRN0BLK5GlXIAkRPQnljkpCBmUULbyPxcDcDxooFP2Sjr7t+KrzP06IYFAYA
IPGA+IuF8tx0rBEuO5pThABjDoJ9Feu6XuB0qW/yBH8sSt71qKF1qkaacto/SSoR
Rv3arpiYgzU73iUh6BjfA38zZjuoeThPj+NcYEVBzS/pNTKsB8oUFyrc2pKcmOIF
fC0V75RzYkGHsD0lqzG8tk+Ddi5AInoB9SllGKv5kBumuQLRQ+V++c3n++3v6Tph
asl/kRb9AM10vK3RlfpwUK3cRwjl5zUBK0HBG1ELLB4b5wUYAiWFT8hv/FdeJnxd
8XmpofebOTq5Ou0qqN1eOHco89HvU6Sodhm3j0EZYqJFQ3HGcAkZgl1/3rx7Gw/6
G1DyhwJHcjo4Zuzd8henY2ruah3BOYYBtkZNrkH1GKzhOURhjBsz62osjPIUgUm6
usF/KyTQ5oEB0Csk+X4pMKIh57Z/2nfFD9zuvO7AnDr1oJorBcdvEKyeycHjh9h1
BuNSM9B7tOibMqzuuBLad9cCpn9clSL/2NoLOqzy8vTXGmnDugOCOcVUss114j+e
KPdx6DPBNzcfD0tjCjq7ZPdWTHvbBtvaDHPy2NUwyJtBVy5zBFTgL5QCHsUtxfxC
M1v+OyH0tg8Jlb5Ojn/c9q/ncGNXTyaJQKCc0lWzN6cOlmBDnufgBAF3WnbFcMrT
HL2QOCbJbANzHpWfvk6ZrXz5pTXksXI/fY3LL9dJPB0vUPQ8e6OP+1m3KveR9ZD/
JCxFMPFoMEqqPMVghs46kOMEuAVtsmlcIPG/QzurlpkoKc14VFOwTabF0cJKrltV
I+yvNspQDTyrN9ZgjOjYou1L02hOEHaqsnVS9OLlix6k42eB3DoDd0hPO/jScMn2
lHvIrHMQvoBWYRKz9HzO/PvCr9g97X1oCyn0qq4U4Sku6/Bb9Yy92KSmIC1AsEWM
7KmVqKdoZrTFpQDBPB8YQIufrRixwn3/0BA/jgqCXfmUEMH1Q15rcqj47TfihxrG
3by+6yC70TdMYybkikvdCOakIwy39hWrXlrAJZFxE1TGDNv34nNBodqqkIW37A9U
JNd7EpVwR1TSUkgymBAl2teMNacpZRbegmLZG+QqDAC5ulJyFUbzj/1jIolsue2p
g1THmVOddvdaxmg4xxYS3hkTvNlrZEmPFxhyoDJ7C5fqkzksjwLimOM9M47cGl8p
0qbcBk4Mvhw6u+Sra6zuufBShttIm8NHznb6iRbqJSpo1g5lBZpJCB83EZUGeG9c
7B1G7vwrZ4JS3E6rJJ5xStLblDFgtBr1tFAXqQ86Ay+oCaCEzHwE9hSDtFVSzcjW
auVUEOPL1uI/sTD2ZpKOsfN0R0FHcIkYNfp+pv5oy6X+Nqgk6B54ovjoqqWIEx4Z
a6SCkDBkbgsIBzf9tUAAKgY7a26endJJIgE7quHnzBUiGMg7qgkb3ELXSCkuRr57
4C8UbEmAuBssbSsKGox6TOK3fTOkCV5SAM9sLSfEvigUoqSkaHCOppfXNFa1Bp2P
R9FJokvqd8I4E+6dTRI9gYZSyXpb3dUPgZbu1cZUp5+Dsmrt3YC9pIa5HAKobFGB
wYkyfXI/WANg+8ZcSUBZCHyHD/Dn9eYyYGqmEnDN+W6cPk05n797oNIGvN76eWuf
YeSLqVGTQTEify55EDBmxlWPRSynqV5zRc9DELTsmFXmSEj1ADoiCRRdtr8yyLJu
iK98C/z4wSStdGUuVXK3AXvXJhNWeAZEaGhOPoBZZtcbyrESOw7tkr2IXY7vUbhk
R7kCC56XQWsTkPgXmdsn7VJNHRh8RUmsCHZMnBwHFz6Yv62NIc//HnIxFUUkJcDp
a4j2dX9JOA1DubqPB42K+5mXHPmRzrrLwkeTYvAZAYrVq1lAFb08MHUnj/Cd8Elc
y40Hjxh8Eb1OsCl6DLkwYLhCZi6LmWwlrb5A/CXDBbgQ/WwduN2FbPUKENfMtJ9j
BCDeKIWksoQP8kwolJS89vms0LLiSQWHY1UrYEFCy+YFFNv/J+hB9T/68Alp1Qy7
TMJRF152F6nza7tWayoEu+MJPY/ekfei6DqXhpFsVX9CRlZ9R1NcR3FsH+pKG+8s
G0csoNLnX8ECRktgB3LtD4/s3gYIwYOu61dapJPv1u9icXaQU5l/0VdUo7P47kaU
fxUmRahY7I+g6wSY/9i8C19Iwri7Ef+u/T+tPXiE+kBkpyBoBQwcw5XNS65AOzoQ
RKYqvTh10RvnOo70EKmcfk56varQ1o3h4b9UxJXVMiANG/VTaUlkrP1lhU6idqHG
WzPBqSNlkTQAhbKO0YGRs6j7hdPQVG+lJENYCBLHVxRt9w9MW1/b8QYIlQ/qrVQw
F1i6LBrhr7A8stJapmVUe70E8LEIQmef0bpdIbSqaAmMMSspb341UG6pTHqOtoKO
jEi4arLAEJwiDPgn3GC4tfvRlFW+T5L/oyLrxK5m4SfMnjvW78JTC0A+UZbhTs1x
I9anuzIn7t4NlY1l9FPHAbMqpCUZ1RPHZnLSUxwgA758mvCha46cBh9g7Ya/6L6Y
pmnOn3/1C/+x6fxvUwwvXT0i0QPeOTiJ3tWQPwd89Lt/7YQpW/F6xUQodU6d8qT8
jsE5Vwdu2Alf6HR2WhuBZYn+Te5BTpuPHZYRQIMiNLII+TwrUncBuyl12ZZEjMsW
TylBKE282B8jGLFxXfZkRVkijX9MWIZ151QsEbVy/rdT9eX0vzVmK9ogExIQk2K9
UsOb98+SVhTiVFBs2JgJb3kF3CMczaPVKuR12OCpluv4OUtaC1g7fNDzFI16Lx0/
nwk6V1EwhZ75C1ncUdrJoe1h5IsMFMZt2qV83A0BFLPdZiMzvbuDHgN0hg+rc5E/
b6iD7y/D0nyLwuJ2SFpCparTVW8Mh7dsS2kFME1UTTiikkOJOOB6HomKz2sU+fGh
DDjZkMJsNPkvKZPiWtiauUQoDAhuLdVD2TftQDFph2U1Bed7M3imBnni9L9ZcwtA
1oLFUDJfofi1c5+vyGjhuOFCWivsTTq8GJOT5YXRyI2xKLLfCEY04p2Q0vljmUNy
zq3ewNgM2+eqMKYTDtJnmzjqx9+C3vg0Jrbyyj86meAxZSvw8MUCPhRSifpVg+qR
dnMxBa2ZHzSfz24Gov/FmGZupisW0yTc/u1To1u84Stld5irkMHFVg9PE0t0PeTi
qAYTg32leTOcwGovCka8lV3RxsE+byGMDpg5lfACAZJezAqnqnPK05Peh5QA9adw
EPU9yOividgtKUUTSy2EA9SEfE3U9eqihnp/7MwEU5iVeAgw7WkMuHvsaneokp92
KA3y9q6BWE1p55+NmVWqgudQQlGJbBNCVXjYev6ANlFboIJz793i2S9VYmyQxLsY
33eSlFvq96fdxW8ctcbhWedK7AFENz/bvzRzBSjgllqds6gL+63r1eI5m9mvwh/y
ivJM+k87g8ndwlqN68uyUYqohqXZCoePnTmVNsYW7aGSoerJdjv9OweK9oH/FunC
rahfyQXMH6I3HwaMy9js4nvog84FS7Qchm6Yt5F2gl5MIqZEw2d6lYPuic78Mmyx
38BswBzJgzqbXFPVrhLH3+QShOHMkaMwdlhvsVwHziD9dDMYeFBvMCv72aFkncur
3+8rYObPE/6DHl2ohH3SwiZg3RnbxPMa+NwvWWOYpx+xxjDEOYXd2jBdfrO38YVk
RsXB2PgjxWE7hVAd8qgq8C2imj8MXj2fCZkOFN9cogpnJbpsHnoc5fwwHM2EIWGn
Il01MjlZJ0FrLGxoJmEfX26pEAs+wE5NNufskQv9h/d6+hQfdXVtp+kwFoSTgC7r
r/9QAGuKLoMsVi5koLm4VGJaDnkPgBf2gToZWAxYwVCoGPfaMKRQptehw+Rvq7yB
nmSmjRYtXWBMFYFSD9kftC7Ci4DC2k5R/3TFmnfqU0uMr0vRZr01L5NvZzVY5Mpp
TduyZj/Qdapw2u8Aikvw2WDNjQMAjA2/edyQ+b/A9w2jYFEOEhW4sNLrQZFGu+ok
iaGVwh/ZY0ckA+4rr+oSBG6jlEEBr9quocAFZwoFB2dVfflnjARj0dWouR0RxJIY
h6BCn26nAouS81Qvew0hISZYm1KiQsnG2NpPR1weutp+wJPSavYC496SVhF9DpQt
DcQEI8l298RGuukbWZqSFn/FuKd6CAhsgnw7aDuv5AabIWs4HWMZV17TcX7AMoRp
glmx99q0Udp0JwbIh+0W7+j9EeXuKVo5WGZrmMJyTRRVMGaOW2wQIzcqH/FFk9j+
v1A2yiNxS5DHxC0KlhKKmC5HY+J7tPffr0+RAt6keiG68ErJJyW77jS13Cx6+STJ
1m7o7Ok/PZADSse0H+LR7g568CNqpd2m8TZdzZ126isQ6nAjn1hCtu6yeKy+C8Ek
9ThJXkWRDT80/bJS6FKparY7l5N05+u3GnIOCW2+EX9O0kARmTQ3+9Z2kzOV9ZvI
oZzKlUEnXh/mB/kHUtDj6PNdIKQwyIBGp+ebQwosKS3kI22mGxuO3Xh8Lqf28si+
dqkYwB7Cv8uM0gIKA/xJf6DuJolW7q5dfeM8k/9oPT4tuUMfJ2VjhsMRBgZ5/bzS
O764kE5Dpcwb581sSwYGCbolF+G5DB0IZ4wH/t31uz4uNYtHr6EsDvOKePmqRAGo
pRQH7+7n7yTDdnI7zuwxWy7j46FmeC0G8j21o6Dx3nAFYr/BrMwT1+aQil2QzbkT
a/CtAKAT7ZxDFSL1NjTlnV9X6pd8eQZUB382VNtTMPbsv9OLZw26c0Rcc0oEgq7A
jYnRrhFRn4YFaSXX9eFG8j7v5RYjutV9sxOKQYni/eQ32QpMMFaj9BrP/c4WjMA5
3IkA7yvnAbZww9WRyAP+iDpS7kymSoydstCpfx39kQ9hNPhsVtBD42BfJ2BHJ+I+
6G2fIstXMIKxIBSk1vknDR2hj4bD+PghIO+N060DBhKlFAoTRdctxc5peAUqeObX
ZNGZIIaJ4yEVNIuHlj65XDsTvZtDAfjCfk0uTG3d7laYcx6DdEVXKv2GCOCkgeHC
9L1r2wg8UHZAXrnFuZR9iPYMKvQ9Z9IKCOkdFNGInMgGZeAvMjkNct5mGb482zPS
MfUcDYbumvxfrUJ8HOCvkNuS6pO38ON+95P69sJSO6I34hitOvXmfOLUiWy+6rGd
pr3xwquAL8XmgIPFthVGtOfPwqNAvHchPGhFSI5E50KbnudC2vUsJw1CAFYDymec
kSxmOllKlrDfo0OMgc45nSncIx5C5kZ3LzD6Qz3fYZz9ERvg0ET51CZrfjm6IMKz
08gIBd5UYMubrns+JjmQziKuvIhtlANIy4BtTaPYUuv1KzF3h8EOPHCxuty4X3aa
baZ2VaktcDYq4FoDoS/3a7VlxqCsnVudmbB++Zw4IFeP9jldYzdsd2iRYdJ1vwti
Uu8blZPho340x+JC75fL4dWZC6Weh8Zee+t++nLKVSZVD9xITFPDf88IMUgTvABN
wZFl4YFKYwwtmmWtGUpT2zM3tZcoVoCwg/2yQ7goPcgv1NpSSUUEqHj5Bup1q/SS
jA+9dFxj36t8O2Rf1E5yQhTMxw5MGPiuz25xf5FpN+NJ7Z8YancE4M/c+Uh/NUM2
1cxI574w9Jv8Tr/Z7nEcryl7iSDqyDimcSALEqsx6gJVEAR7/UkvTrdT0FPKBzov
FRZesnzdCuNYchEXNJLTbOq4zeLKky9DZZZs3hGCL53irZz//Y8JeVi0PDoQmkDW
04kTRg8d0oXjZmUV2lIm4PUq6QIWxBuNjP7lAG99urqdY5hxc9lB/R/fc5mSq7JV
iVYvAjy+DdUNjb5tY0bQ4ZWqp+uslu/PQu+MH37EWvBAKfoqjd57dM7jlJHPp0rx
qJgr1fKZk8XAMPjVCA/3T8kyXKIg3LDSOFLUgr0c/bYRvMTmhbNUpqCDFMVb/Q+w
lHp+L+eexci41oKXySlNqxQr/FESfE4Y3C1bvE8r8j7RCJKPTixjWVfGSA6BYVTD
UgMCEcgtnxwjkQi5Lss2yWDe+Ve3VHk13y4OgRsV0UaVK9rCylm0jL0wByWceiLQ
wxBV26DiOu0O377l0qIVD9hang5YU/R3RIj3aFffofkPfiyEKDBuax9NtRDA2/L5
46fwGIfNpW8Q1CH8rPsFHGLWYXmjjlOsyaUCgmpJCwya6+c1ww+F2ACYhVu4R21w
gfmcrYjvony+15ilAFB/W9GomLUa44nRde2L8y2A9yAwNTeGHuIzQyYI4Ax/BGtJ
Zob8OhO4rVq/6/Ipy4lORqlTtJAPnD1OsuJ7UwumYfoetY/f1tYGf4ia4UbAyzLk
0OSfJ5AtJlsJMU+Fp+iMJSNXrAuH88JQ2ndBxxZe18+7D88Hb4lMaFKaawEGMN8H
hiYvWmsHz26HQ21Mk+cnDRM/wrMWvZj+seRnBcu4yQCUsTdc0tZCS30+mYGSRp4/
6Iq1cOvD2/8CEl2Lqe8EyraYsJ7XEvlfcDc0V3T/40qeeEdNxU69YZoEA5pvi9sh
G0k0D+vSBncSXzHzew2i9cFg1lq+m4o/eXoL2w581FnffGrMr67xerVcAYvoBYyT
i3w7feClLwmDcQM5DLTuHiOBz8axvL3cQVmoDi3/Zgo5HVnhgV/MJlZtn6TYh3iD
vwr0rLW9Oez3MDPcsw8DXyleubC2vO3wYRW+9XeV6gVBq3YgcSiyUdS70rMbjKyf
l+WWgMlqszzuNf11SPbixUfih24Ak3tocy65DAoYuEzP2WMwKXTwu+2yu1Oh2Q4I
l+FPew1JaYa14yDWaYXehGFsNqbNwPbnysuVcYnwkmZ6kR2xsRmVBvtn3VcxPY6s
w/++HSfHNvNIrcrlQ+q4TU9QWPe8VlC/JPQg8T47GPd7ZXKZIM0AUKpFJFcR6tXb
hVNT0VvtFM7SlbC/h8AXblwa491V8M3BW1aLtbVBzIqFJ3yrrJwkA5PRDIfPkfIL
kWS49uinX9aF62u2UmNRo6Y7Dw/ZkK7c2458afYhkKC85GJi+X6TX0b4JHW8Ff0a
eEdb0qBO+2Sq3OTLR3lRC+5dGngMGzmZDusyQryqzBV+lieP4a1IsmpDlydPETe6
dLUI3XuSCuGl4sk2zlQpRKbHMcmCPC9NdHbnuaN0jN3EFE/WCTOVmk69goYDIv70
PI+PJPo1hR6+Rup4yBTjGFqEfAtvU0Auda++9PPfK0oB/7tqQKYdI2gf6Y1uVHGv
J8toVgPvJ5a/JSABW+mNv+35HjJUcyQz58S2as9C+iSFd+0DcFo7Iv6JAMc2K/q6
EnoJ6BeW04Owmh1LlMjJ+rl/YrkjD6KpzoC/+GGfQplVRK90gNT8l2jMy+1QWRDa
tuJ6Xdj1mTiGf8ytODN8VphMpQSydyq+L3Dn3dolvxswrJriAk1Vc4WtwG0zjrQE
0PfIpALGsjFtlnRjflpVzr1KIWfrVTPkTLjwuHCu0iIw/bWyoQDq6X6Pfk//6M+2
PuvuUhZaKIosKZvBiqjyO5578ZhY4u1zrsYS2AOxvBa9OVl2cvm1GNWJA2Fx3oTZ
fpmaJa7OiqpaUVDX7+NFbMgFsCjppRToRVkgmAvGKFWcfm8PVKfccr/0zJXnpGV+
LXnFUentWBFoDLrxmmCkev8nLSCS9mXKz4Wd7CH7ZnTQaVeSWkzR/0tX058G1KId
rAfBMxjFOAJ6Wbe/ckDKHvm43X2sE9xJlUF6tMPtRJDEly66gkzCZK25SvgViz0T
cx3H79qkq8UW2xHB0n+jNg8DRgKWjf+tJuHXfejV2nHPHGdjYOIcd+BTnoJK4Uv3
LCJ+1KB4H/u3l+BxGl2lk5C7e2dCwG0GDGdJmyPKgsAkC+birV37j7EQPllIxkHW
pYYbrk8jCdarfxfxdB8Ye0Qn3qXWSm0bWcqE+B6bD5Ws6KZ1OrdnpDubHqlbEWQe
A8vuim98TXrmYZ2IraLEoZNRDeU3gUD8wPhrtHnAKcfwtl6y8fUZlQHMCRUWg6+K
nFyiLJMz58lTb7uCUMEb29mgLVhEZqlJwdL0YAGbdnppTVPGfnDvzPV6cQU9DIL3
Vc/2Kra/pLKpyhoFhoF0X1s1g3TzAMSgJrUW2NNEkC3FbkRVfUKeaeDoZVShQ+NM
CzQfmVxoyNjWF9QvkUzJrPm/5Iaj32luxbF/AaM9DSCRPWGBNZb8pGCaOaev4M7Y
A5eJ9qIk9CyEaIqLMS0OUQ5dqRbi53D1uoXT7G/9anTdbOa3hHIqo6C3VXciHfzI
2YyDxEE/XhaLhjg2VA25nnb2y2Cs4bgVkDRZldxRkGy+1aqeBDRHK34E0vKz186W
pIQnqtigYhRCjFCFLsNozjW/MWFYdgpn1o4GjY0xmpg9SQ7dpDbU8opxg+Cvpi2/
gSRglEG1Jc2H9/d4nr78UVE/JoNREgEke8jTxmAd1q3tSqm2aPk4/lrl2fycUN7d
cVGyXj5HCI+UWmvGCJVTMHmsAJMB8GTLptX/2i4Ue0Jvl0sLO0eUcwvQCzJWESh4
FeisbSo2bTCxRia/7CBAhr8a2ogFj9ra0ocatyhjCtS0y2x2uhh/obZZGhpGj1XE
Hr4BE4Uh9A79qYRJJZ7sV8pB8JMUzBZkI/FR42bqBKpefPoxsdUcaK888Cfad/HE
s+4NBLuSwsdFxnsFabRIr/oe5WFXtosCLmlwmPPPVRR/NmEL3TjboBup5AQr5zh0
IXLO8Mq8aH2F3U20wjCd6tURI1nbnCqFjXHZzJUTDp06JrvTB58jES7VnjOmsTPP
ba3N1+qsbMCsHa9DY+jaEVjoUZ3MSj1paDawd/uw1At2nRlgj3LPlVvZhwME84K/
iLV9uvNk5Wx9xYq+QXLiXRoCe/MNghCUgU94arCZWeQjCPTeIbvQUzjbvUcIVgHy
P8ierTK8NO9VvVID0Yj4/0+Z0m2ytApET9gT00qKZnlj5to6mfzKwkH2NUK0z0eH
6AmaoHlyIVMTjSaf2v+wGO1DOqs6Zb/Qi70U/oTNG7JzdLH1DBF4IYCCGZu6r9r3
bQ9rHAissyjbwf+Atd2rHW22kFe+GlSNSJpWInAASRFaze+xIikYfnBgenJyvzXv
lmWhCpCfEqO/mbpYHFvQveuisjWP1RA8sZlbrzuRUkwekDsGBBtx9j9HSCQS17Bi
KaKa1yDb299gauq4PMCNjnnqeRYLXA8uZVpUI0R7igBMcFxzdNe+0jmn8ZR3td89
M4s+b+CB+/l0gHDycZpDEPkvCQfyPZywL3PQwjUNAZx2hSsLuW7PpGwUTShkzJ1w
h1Y+Ihv1d1Wh8+fZ9dKdQBtPprPBKBQ8p7p/uRBrw4iYtRlnT0+iG0TIWtT9tSjr
TtUJ5lQpPD/5PrIrxQbbf3lZ9AIc5vBRJUmH6XHhHB90thd3SfASF3aEoqmI/qKU
niHgc6+EgnaldjaIAov3WQNlYttwXbOUWjeyMFA/3zhjytov87KMOUlv+FSqjT8/
sPk/RANGkHuCD0CTz9We0S5r46arg7ivI5KddgP55OjrZtnO48HnSY85ZFc47XbR
8F01Q37iXXgkWviQlfIqQYP3OzIW+y+QuHh+TyjTMK07aztveqbwIag1MHM1ui/F
+ngXqTGRBCv0tkWIUmBZH8R1wCWB2Bsdop/yLlXF0RYMr4O3FYWA9dqzyIkYJ5id
v7ry001/27Uz8Ky2iqcfMsArB/MSyj0eSyq/flzZyt7Zy+0aLO6cCUEP6rS+te23
Gs1iOJ5BrdA4xwmlmRBIeWAGLNpYaXEuXQkAwswNBRChhRCuIY9qrfrG301uFNdw
6eX/AIrx8RN12FYx5HrEKf3U6YQkEgXMjdzbLOA/IQfLYcAg/Q4RBCoF26QSAl3L
7RXuHOm4xNx+0AeXyAbdaZu3BfNEuF3EUvCOognykZR7COPC1Wf0dDf12vNY/3m3
xKK9dh+Nl8KIrXIzkvGoiGQqBsQFYbxELemblEYw+WscSuKuXSO8olr8lJHII9/u
Ba0YZtyJfc+h/3w0DujVaqtaj9DFj6u1n69dHGYap0lOXVERHr+u2+JeczMKh81Z
xWzI9aEb/mcPkRA89UihCVdCWA2p77n2vM30XkTigcERmu2N02Do/yJgYkNJFu30
QRtbe+8XnWbjsh9F87czpEyZ53gq+IqoWam61Kz88yT3hk7Mf9SQ8INI1Yk9uZ8J
bu9lZDbXvB5/orvTo5SfF6kPFO60LaGy+BD9ZU9X98ujXIvjCDfF8qQjJjKSQQU0
3jPPtM4nej7eqX5zTxlQb9Xp1jLUHZOAxSq93sMHjOozs738x9X9gOBFgkHHhyw6
uRRrhYfC502aljc4EmJ6nbAu8SCFjhcuGzVieqaXu7kqjoyvUY53MERuxlNk2zVo
3LkMD6TZMFwzAyhvKbI37t5maxgvfeovN4m1Tsyt5SQEu4anoNMg4zJFV98PGGSx
Gm8fmU3GrgryedxWmoIM6XBMyx/gzAM8P4Hi4CPtJtGWytDCH/G10jJgRTv+8o7j
tUNsj/D2fI5+vGz/ZqNFUEVJoFmVSiynzzvHAMmLMRD11PL7w+Z0ny7ynNBWfh1g
r6Jruk3GNBj7c74+7zbgdeWDbZyva8AW9TuyTiqcNINchOuNvDETxY8/i00tGALh
LiCbMfKUi6ZN5ZTAoD3zqNrztiMbdsFSaKVsoKi7PrbcMx8bsB1mLTCaKXHcGctu
k0aqO0BJ00vtsIKU1QuxL6j7/MyS0iOSvUOF+VvmrjQ4iFASsbbl7r3+41qzGLm1
QSj04Gp8dnyaO3epePH73iLVrf2wNtw4CBvU332mbn7kv8VpG01up1ZQukZuLotE
JxeWWhjuV9NI6B3mwRN+DOkTzxuFjUBNYQ35M3eJviG6kuVmBusfiMhYPefyldl3
WzkAQsB1d0B/Q+GptyClCLcaP7VcDWRiICvKUdVz/9B6k5g9afJzBvl1YmOO7xPC
nJr7M7I7YkzH4WCmbvo+CmsUkIDwgDAUAyEUUFobkhaPl5XkulV1ehyLP7qSZeo6
t09UWeou8CkLcgRxCLIKuHbDdBU3vfVR4/1Wis2t84BdN2KlCfGX1QnCRlfzK/KE
0+XFNW4/SA5gLJJNKI420uNdUnoL/uZMCCGjRAouyAMQAE7ddsGFUivMAxt7H1bz
0DD5lu6oCIKcMzL3l57VmYXUKNcz7tS0kVBpus2Y5p3xkZV5bfzmXIFTbX0kb3vp
/YQYuwoiQWlO89OWB9SPSgeIuxOeEf7t+4Zc0+apP1BZ/4tikFQHH2CSEFqMn+5k
dvcmn4nxxTJjWx+U/NqQvIsVEVSopPhZ/8glMy4WR92vX5c26d6smhq1VUsg9DJG
s2nXIbaePyI2Pq1VGvIsBm3hHBC3fHLisxT/yH9TX6UkwlrDI/YgtLrVxm8i/8lN
ofJQ1xC2Xogbqp4gatnJtUxIYbFjRepgUyr9Gok9ISAGmeU+8Dj5pfo3I0UiE+45
T8H0CwEfDnPTrqSPkMGVpbzyBbI7UFXaCxf10gPhFsfXIkxnZIumWo3tz8FklHkn
wyFyOk65uR5vkF3kER9egl8Q36l5CL3AaNuYH8p8x3dxka18sKd+25kBjASDgEng
flp1C9clgSI9QpFvp5kOUW7XFJmyACvTlJVqdlqGB4CDB5fKh0KYYkpVQJweO2Cg
RQWxo3jpz6HIC6hztKBMCQw/xO0OSBg2OzAcTSrrAqJvqIdGcXt5lFehTnZHTBfU
a+NVgkE9PEHiCzxxWsgIhBOP6ELT7j5EoGOTCoWPhV9IOuhq7Z8+ARHtFhnXgXgi
hI14GtOTlXhWKGJkYQDfvNReC5cXEdWqEVo2uEVQ9VXolg1Z0OEkn93a1fSH5awh
FPRElol3caw3MTK0wm4qJ4C7R7XAnP0FYo+Las+5xvBwS0Tsf1UH3aLg7w2+BTbq
awevkCVWRFpEi0Er8Kx3uSzhm/18eMATB3ThX5v0izAQrZDqy9nji5eoAOHYWNwg
t3pN4t2CFxWU0pZWQqo9udG/AXjlhrIpFGVkoV+2d1/wpu5xEZzv8ASbNd3Au4Sh
LyF/TT9RiFew4SE98YKwwxjpCWZF0Y9Ay1BvqPI44+ZXFYj/07oyboPayr/M3BNQ
X4PNhy60jSV/rcl42P1mqNR8dvXf35DBf/g9vo83e7bY90Hamc+4+MWVuvH5M0Iw
iWzgZGLrMcuPN7Q/LAhDRX01iWU+8slzfzQh1DoSj2vBYGlWPdWUv3lYhi+RN5mW
VfCDCZsBTS0bK9BbUkPzgE0ueCihfRkFLflXhwed+wgVHSd2tVblKMeSpYdt4bIo
ipLIrSJQeNsz2lkGDyHyVZ6YLlDzzKSP+hJTOej+TxsePyXMt67Jaw9t0dD7y9cc
eOKPA4JvH6fQPcB8r/sPt6d0MnB5QFJIHYV0pIhXQrEgq5IOaqMy7a+pUb9xeLtv
qeRhm+19VWGrWkkmcaAPDcLjiUrdD90YPrBh2j+YU1ExGzBV4lIamBTnFd1AbbCW
ydsnAGVjkmm0ULBtGwBNq+aEPUMi8hSLW2q7sssx26Eur4RT1CWJI9AZvAIUiU7i
XxvOfEsow4fc9Xm/XU+6u1MXSbshRc0VLSsed5TWyOnIh4MkXJz12dC7+tmIgZzq
wtVgGSzMQ/PPrTcTdmJ9qSW2Dj9ZASOyz1cYgSnR7H6ZmyIsxsnL3pdYX75WjoL/
qTwR+HUSx0nIbhESOA+FP0qyPodj4QLNbE2jQ8iG68zuNKMI64FxRSVy9588MOOr
ENW50+AriarnsrahPJx3bCYY9goWP4uGE2p7xjQVR6Yl2trxAm4lWP6VFaLsf+Zi
aZjKHo8agMMWlPT0WNNyFUXtc38q98ZbEYjQrhrFsN9EGpnCUeVl8Iq6fc0heax2
K1dCheJO/8xJXp7D2dRerNDV4uConGJfgDaAtY4/ovpjOm6CxG2JApCaQ05mZh7C
39Ip1SqTTpzJ3tP88sG9GByoeNfALD6gM0uZGz8JLCe3CzvfTq20DP+XAoehrAUG
rmJiz5GLbX2wmBQjyvlfIjvDplYHakjKRA8z1xpciJcu2BjEJX2rJ6iHYfsarbBT
FJvWH8N3i8KcD28lfb8cxTdE7rwIu/JRHmmPyiP9/gbZkl6NbmV70g/7Lf7EZDzF
euDQYR6vtZ8HXST8wBJyQfQS+RDFuXdqex2ASVKGmAr2ZVkgCkxgi/pQ8askjnQq
VCJ3+/yumo/ha3V9neAkBpF9vEAzVD6zrpT4eoW1DViTkVGN5inE5EYIln7U2vtv
600lC3NOG8N+F+LHFZZ7ejtopVLcsddsbszhDWpAgxsEbphROInHaz9WMx4sQY5a
6BDbIVF9r3v8o34qQ50EHgjI4vawa+/AKVgya2udmJfbEk59UCT7BU+7ToWLW8GM
j0aScgADG2G8qJ2YDrxM3EwhA4C0SQ4RM5E5whC9wv0SWXeqMfnUoJXeEHx2/qr0
ZXay2TXP0kwZeUr/epEHv26MyACpQ5WgJ4GEAtNcCd7TPUVwOcmlJeOs9XkhsvXM
kMD2tXmSu9tVRjOqxVWGox97WWTbmYQm9QlfNBvaPEVIM9sd1tCgaqGKAvPJp38l
FHjUR5b/an5TWVNQiQj2dBQwTgOJvLmLw9QsNv4Omm6Cf1qRJ1153ac+ZZHuVHBH
3cv8b1kaYM1hkdoe4gCtGEATGrB60T4DxygsTxq7ULBlD4cS6Fe7GgXQPkfstRwg
aR8DEOa8kyyI0KryIAfvA3W8Og1Ns44l+StRNHwyyywVC3XhRh1yp07Kswk6kAPI
7zfffRenP6BpApTxdpJVN5M8GVhP2aulWOPEVbCOt61y2WxqJ0UjWsV/pfqP5a/a
N/8Y5NA6yYGy3OMi6Fb401aja7xGe4GKSSZTKvAbI2t/zhH4KwJo8Sey80PR+rex
ZjSB25aX9Nsu1wyQ9EIeJ52h1JnnhQfXw2TBi6/tu1If7gtRa2A5ArL3GMdi455v
y7p3Suyw/7jfxsyUfi+ZPZcQ4fnRI/XhmNpjnKCipFggXvJpIizOxabvKOyeJFnY
LvbQSrScN8CI4+YFCt2JxpcnmNtNDOumh4ZsG228d7QKU46n5QBVhH+2LTB2lRTh
gI1W53g12ArWX7R2hAl0x7UUrUCgxVsiwbfnq8KhGL+qDSGGsDovv9OxMhHUF4eT
F/CXF9gTFC3Q9fKyLnKCVu0Y0PPrjiApWHT/sE25POfjk6S0VbveEXS+S+GAmc5J
ug7AlQ2Fz30NQXCXAT17nuuzuHO50pA2dOut7D8QlPNctuKum0Mrpp7dRGwalHIp
Ov+eHsxATZns2wOnsXzfgRceKsGAa/ewMJpEh/3lgZiBE9qKbmxeLgtihhdGcOO4
ntBd4pNDxQoD/GVzyLd0aUsWUWoC9KxHTvOlzqsLDloLENbpPaSXBn1WY4SV85gg
ee0xg36kZ1KuyTyVOvyHI8Ys+D3Ydb0BTtKgiYGFAjRY5WKyFr/3zLyXaNwwLMfw
yVad0GorPxMvx1dDAzS/tucBD8FY3+sYKGgrAJKbgm5xjyIV69vlKh7DM89itrLz
/zQwC/aB+6bzBsEUZ+YxfxQD7BDjHWon5hREc5cIbaIcjtJKu1Fia7orDATjAsMN
FAvSdkH0hb8ZU4GyYVwFI665GKe0O8EaZstHzeJv/X718JG7O4DuEYyT0fvqdO9l
GfPhICcu+bW9baMYtqiLYhZ/GE+U9cKziZyRWVwS+uyVSctHYTPgWODh+ynRm3Vl
MzuncqgeQo8wGbCAw8ySi5qMzAE/PW77gXdYBApS9trI3sFFu8eyXGuMSuticisg
dRURQsKb/W831yETsKrSN5YG15ZkmLRqU6balFbPFG9A4HfH2Npxc9v0FidQ0SEj
wGtciVwSmscOlaq3MiTrYndikjQPaUNtR0ig7yqZ+4KCDY5VnP1xe460snDlRB60
7rtxJyTDSHxK+Cn2wRTVSy/r0C4XxoQA8V0MInwrSu15MMqK1xWEjD5GGJfG0Wo9
aF/wPQJ0HRHdo0FemLt4TaHnX4QjvLjMMGyxKx3jTGUjlef93wgtUYWSXFPAIUt5
JQt89MK3ZwFo4QOxQqwecA2VbFw0/8aRK2AkEKNKPYZPj6Vlde5hGToxyyLYrMjn
fWBixLz4j13YxoUJg99qgcFBB20FpYC5n73WL7lqAvwmjnfQMwCX6y5isPkCCRST
8Jmj0x9ajfiRlj+gjBZ3EhjlFWWCg8ALE405L14yfWUtL4/7ZEnMtBHMGJoev86n
5rLP0dUGjmuPcQ4Kfh545caQPZ77go/woRYMNnBLV+kbc8ahsDbR2cM4gtLi31yu
DZ0aZuG6Gnz3n28vrtufKaB0ZPbTEWP6n5X8BgYKZeRbx0JPLZb/27plMC7xdpzd
6G7F4/S3R1HOOwsd4zKh4s9f5STbB7qxe8Mvxx/eRU9zKn7SDZeSAOsXDmi7M+U3
yZQo9n34Bag8YYBua3nZZo112T/j5Dim/wHWGG0kpRcx8ZwhYbEV9iPYm0d8+D8g
1ts67u2ryrnrxFoA6ev/wGN1YCybqavCcr1umak0OePsXYLPWvov3SMAMT+JUzg5
JLg+hmjTkTHlUwBd02Wuq21Fquap2fEqW9BNmp70PW8SliAF01ujJeeJV24UdQKy
gUhHOAu5wDx85x+4sqHFqCukshDrjLBlwnLiYs2HDwT5KZuPsPBsYVE2SUc6YUzM
EEwvVEL8ALRkQaT+5EOVLctqhUrFKMtgMKfoi87Qr8svONC4tVG+b+0wNl1NSfIF
o6POQuSvX3xdfamRToaAE+FHUR3V5MndHNqCG6A6Zh9vHMqA/0PIaU7U8Wf3CCKr
MLKDQzQ+dsPODFzAZB+CWpRbYagCdyRrn/Lv2lRDRkKVgMnS0TnN4YEa2cc01F4K
fLqS2ck0liVeFj4dG206A0WdbWTzuIMULCLIzBVVRV1TesRD/k+42rAmOQC6YsXH
oaGsarhnVaeFwcHPD4VzgSthdaEZ8s4K/c/pqgUUAFlGzDZ36DLtPHH6QxMfCFhY
tT1CIUz1L0Y9+hKqNjsCxDro6Ect/Qvty2vdCiPb7KONvzH8sNGMwW/3lQgwblsT
JFWpgi9uYHcGVI1jwF4xomJYwElSz7hnQ8vmVz5ZIjRUMT5IbOeH8Gej7NhF/5j9
3bZV2uXUhXSC9RoCcw2N55s6cIx9rZDxhwbQl2H/VPI3HNeoupavO09IPbbEAPVM
gLc/acY4cjdwoA5Lg/iQrtzx6LYUgu84NHv5eTJO418cDGPYYRDdmAba/B9KcItN
VWqPsxqFaxdxd4cPfZIFpyvgK3MKVYfgZxWR95IXtbru8SUA0fw7eKmPga+fkyEd
vhBuvUspFhsooEJzoDYUJVB5Y8QFBjf7wjfXsVH4PCgV9sBTwthMNCfOkmfacOwR
bgKMs8vnW3ytL/PaCoYVaVsK+LQ9oBx/ENls/+NuiIggy8CPDkIoqHcChC6Mk3BL
Bx8/My2CPPuge1/I9LZjkXzCeTj9pZp0r/Jzr0zu/bzK6COeg4Jb17+oE7k4CiDz
CbXy/q6WfVsW9GmZYC5yVBQfmF5WiUMOF5ZSHEY4MTaGgmYa+cRaZPwipK91jiBS
bLfsP++dXE39yHXXK+dvpci3XzIsDYiQSzc49IzibY/xO4FsEM2W+fbwDv9Pd/S3
sapPRg3dqB9oI7yIVbpA/VnI/pK7n9B9e3Q6YAlBo230d6OEYO1yZ2yZ2u/13fjQ
1uDgCb09I3D3U8BZAKUW92RIcfFWoyYdE/72f6l/bMPELQ3JKi+KWU/XKmL5pGO0
P+QUHbl33Peex65mto7DZU+XCjM7JN7asZiIpJAEyMK56qyNEFktcf3m2l1jQO6s
T9WfGeGE4sALz4fI/klJt4HEqzJTcyDQpTSRGjfXvbbLryo5SXE29L5Hghx9ZkMu
yXWRbAVfqLjzOmV1GxOt3PaZRGG6Hs62yxr6YT3wxLftMYmu8vbOiqvMIf/rfd9Y
dwqKKywP592Ut82b5GyNpHl4deWZCNljClY/p396ke8d9a3lBGVh+uXTnXYX1REm
FmTnNjt7DNh9gNpVle/Eg0wJ4lmKe+ZMhonvde1pANDpP/mKLmW/kRHI3EXbUV4V
c1mvwaFQci4L5PwZ4aEFNBxv3fH+FPFB9MdlPwf2E/a8XG6hRVMn6DtdhJtqkdoL
dHvHTJJtWo9nCH12dJwlK++fg5Ra6bff1PynGsq0YhIWni6pt7zf2pEtwXgRL1gO
AdYe91WsMRaFSjLjZZXuVdai9mHRGoNkiAE8jPPIb+gOd8AQJJRKqSakIz3kPKeb
848wuIg500KKDhh2FbcTdFin6FSp3bKxEBA2z/y2j6JNenf4SxXj/WOqFcHnbeml
1gXexUPmBHvJxyLfh/n1wC6bkwFdSIilVUPG/bLL+SSy8lSJRt6emuh+D5IMvZxF
oD9ptyMwM55BLU0AEAFdnWcWBbx2vkW7yuXrQDIabATa4trH5Ox3B5a/6v/Ho5Xb
NtjP0A2+pdEP9MZLNnmG9wYNecv5c+T5kKr0W7vpn+dCQ0uR9GRvifquSmlBzVxN
vtM9qIgNe7dfg0JBJtAYiaURwImLHMTvXmA/6AcYaIVs4ALKOFfQ8P/IJWjfimuE
T+1mj8dbs66Tt+jWnDNmKypBC2cqG8R7JRZ9L7DEoLGZ5EvBs8FN46lxT+snw2b5
GMRzWxSxXDc0TRvzrE114yavuKFN5+UDLhJmwc1xWGqiXHKCFRibZUt0Yr9n19+T
ALuYWQRejw+/iQGsNA+VCEWffZCqPvrTnlVh4/AcVuBgVR5jlWBCOFKkW1sXg+ZP
`pragma protect end_protected
