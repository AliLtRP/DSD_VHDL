// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e8/yejL79RDbj+YJ7R0d5s4/ZbpUpubzb2pyL0rEtVYl+NNP7BiE1E9sD2XYtToc
OpzmN82hjx9AM1Ac1XJG+7OVkrB65rf4YrIrqlLqfU82SwmlJD1rC2e4IosXiH9B
YC5T+UdC+6gNjKela5h789wWklDC3c1edJflvu35SSo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14048)
ZZ2cf5pFm5wpAyEbBDEHbVzI5+nrMOtxlJcFkNrwjluY7b9l8qhfrzyvymsD7cZg
UkJiPc8vq5Nx3lDu2O1VQ8k8qcGHDj8a63acChuKvBVncRPdbvDzp7lSAufpgK2v
zXQ5WO6qtC/0SJx8+GPm+AG7cY5/qbwcl7EgS8RaMp/yBEr0y7y/PEisy9HbNPQ2
tz6HCvbZrWQ8n50JxqywPDz5qJQjLMYaMXGbJVtpIVMzq8YHcVmd20V0sJBKb+Bh
HWGySPAeLgWFsfOh0R0TKXfcDAcaiB/egex6yQyJEJ5IEZjEp/8YXElev0/bzplh
xFQiY59PJ5WIU5yHVj2Gn8BVtZl29L+ZuB8vBjkGeB/PBKhj5zltvSr1q4Rh2GbK
CKD83QPrAyWhERHFVqJzLkOHjGwNytkmE1WKzHyfqmS9YJ6BB+rt5bqpB/ZAH5/F
BLnFtH7Pa/hrxK9yz/3+rnImvZgmZqu/mokyHTTZVobrrhpfnub50UyxUW7UhjX/
y6csG6qMm4wZyVU9Bq3/96jo/KwFheK7kVio7D/jos82zDYElhArfRy6wX6GIQKd
obTVT0HV0x/V2fipipUrlWR9iSrUgYLVqNiKXg3R5JsLYd8CX8R7YVl81FxMtmTo
gMV/sT34aKuRN7fMwo9F1TGT5am3ikraxp8hwFXCpA8MKNrmT+SeyQohkRpTjoQk
OTP0pLkHENxxTbedqng55JMc9jqsYehQQM1JKBScDftmwulCYH4I23d3C3t1Yb+y
MSSH1dO/8ATzDy3YH9pz3tZCC5lFq2EQgCGon95WVu1sfkcAf+nwzksTp9K+OJCT
3ISZvIjo1QUBhDJSvD/82QMWFej03AJKaP3j/TMAqdyMwvwXbzDzO+uLPYC9Nj9X
Z+SfDuBKUmmvSTWLfJvBR/gW2l1+CNmjJfsjdjyrd53IeQfci2mFpS82F6AesTZn
r5Ji5X+vxFE1ZeVOExtJBo6jzWl/ze99bPLXES8Lreu+zWFlSYHZNUueZmn06RQU
et9C27HzRIjtpLLT2SkrcBb7tPO11UU/WCL5A/YZQJcuttC3nKFKrmIk2vM1Cbfp
lBl1O7Eh28SqX356awdCx1Bjf6NQS5Stn88FbxCZHV/+ncg5ujNCMmpWfof8ZKqz
9Mr2T4MLOqj1e1qHBw4VZ/IZldSfMjL9K+9f6J4nA4uAWwjhPDCqicjz8/uh0QhI
6rbrhXz1JHAAf5n57QxPbHleSJhdWBnWbvV30Ovv/+hCZns1GS/KB+mepVxWiXZ6
0yb3rORsKYDn6TJGgXbK6u5WOyRNIsuQDRtI+vugvtenrmCyy3Cv1jFKwX1dYnlD
sQb+1Xx7lwmiVfkC3IyPHr2ZEzTlY8jZVpWQfFcnsy8ra1mbrOHlZzdfWVavx/sZ
0S+3rWGDoTt4ID6I7Q+blAqq9RVeY3nyjiybaYJM9RTZK8S4R9egHqocxUAwCJcc
ubrwVG+NxA5iWoySC+VUTsHEjQaaTfZMVMFhOywjsOOaXe7kOh+VXVHH8atYAe16
avr0vF8ubjsm1LLDeqrGoYN7HW03OG22PXzv+2Z16NZaUSzvpmvCGaTdCJSfILle
bJzlXBn0x7TD5wXownFJtd3DwJA0gcHEd8e+iuaLAoNQh4ofd+zBEsaqgCVg1mHN
bPOdvpJWFMZ6QGZiFB0qOIh8l0gXGguFNheGjOu0FltNli+SRaJJQb17XbkO/oC2
U2AysOjAJ1fHry+3uWbKcK+/s1tIVtQfbH0KaUnKQL57JxIc0hCWTV3kk2GhQ6h4
nlUrjDqPozgmsXnX1VgDxnQYelGFAs4E8vKiZNEA++QIgC5rjoZBvczoLzlH01uQ
ehcxj0gfC48/NSMvRHK0Cgd3JjBhaw3t19SuNzYHeEs7qmodxkQAipM3hPPRc1O8
hr23mouJSjIDb6ko6ZtxqXbG9TWacdTeib0EvER7hBSaLhzRhBgkbgXiS9vTciBX
mY7W7xMkSpmEZgHBBW9keygzCTPFLrMB0Fd9I6Fa+l6YtRSRR3+e+PZY6ynWxd7h
xeJZFL214P31+uC1AtdqcBv3JzzdXKx+7tZICZ4rK9FHYtMyBil52ElCC1jHJPe7
kjoZ18tNddiaRhKrrtrTrOEEdXLazgnE5iR8U/pyjbKWDzEg07zOD+0BfrRybSAj
tVwRktXm6C/T6yz5T8SIcZ9lXADwBOlXPZTGDeWDBs3lYC9dBOwMsBvyD41AwsLK
T8Ot22D18vVgc20BATCIf3hqiUUmBoDbVnW92rXZfZhO4Nc6iteJptxAx667Tij6
L4Jj/yW3YpIXgzfICS8+qjHD2LPTez9dRYQ/suZaOeA7fLBeG3C0/58v3637Vxkx
i77Iw1NFSrGNIQwCQmKwe3c8YmHrTKvu/i9pSv+Et7cq/AGjDe/f8ONJFcMs/+VC
/7hORq1jKKjuSavbQuNWUfcS+TlngxjLy99Il1Vb/nlhhBXZ1q/VJzr1Rp8SlRVN
lMeoIJd5KHOsN1W1MSXuBuYXpgD59YbPzV1Zo3/6pUWFn0vivkX3l0IzT8JYtTRi
GF5qoImlkCRY4BazaLavMDSzwPVJoCcAjs9dXp6mG9VwYb2kFPzDc7jOWmKTb8/9
O/ReFe6UPtZbTHfNfLFba5LQh/6J/VPGIwa+gxfn4cWJGT8RD03wLUGbIjaZFG2a
ZhawXmWpye11uvk6a2xfA57H5ylMnzH/+0upu4KZyuXLeoexf09BcHnKuBP2GwVL
7jQtpguROXmw0mOqtNzWQMxMUwS0Y2qseyzF/MhVLJoBE4ClN8SXxxePPF1FIupx
g4w6PmtroV1XdFBk5u6YQnp73wtWuquiA3MPgkzy87KJyr3QPyiRvgKk2/XrGrlX
+nLotzi4XG8wF2qlZUJfrweyTV+MoGyKNjUa0o1uKe6JEorgKoPNA9oc43Qjl2XR
kRuQgMVc5mnX2spobXDZ0gD5JF4THFPAEQnmBff3zwtaZJ8dP73RuujQqjsmsv9c
umIsdgb/ymFvePJFHRcb3iNHfr9CeONdd/5cpSWj9O9lb52R8z4baxUKLAhqRSxw
2aZo4BIJf8kJYP7c8HOyHXinNQun84O7nBJUkrSM5o8VAaW79ok5CAQSSCAyWt0K
9GVcdA/9I6UapbH3gWewLNZjgUMcIr7asQDdFK8jI602UwtYH6BRY2z+3vKNRgvF
QKv90unNTl4lIics+23YWyDkIzZPbFXIYeRBlRUH39AxfocfNEzBjgVeygdkQjg4
L0dLyFNS118U7x+84b7WCxJ2beMVxtjlKtvjvfzOtQnKX1EMb1AQHk7+uSW6ZS7j
71BFaHCQEnjA2HnNztN2K/QZcUwAZHNCmYtrjnk8NJCIAXBuo17uNvhFq+rrBL09
MS/+Bi/SjKUqHnfr5FE95v/asloVPvRifdU/xSuvfMUD0tC6xQnbxjLcDcdMvgOZ
znacoT8UwtI4SCLtFss/v6Wg6fO0aKBiQmee1BzbdTqq7lOog3fu+dmAsfOzDBkh
YuYQH9TjYs54Vo/vmdL+Pt1tuRR3RFt9jZuMq/I4gBfsXMc1TotD6n7qV51X1sjB
nXGJPsiF32t1x6BBWQXoWvk2B0xslG163noUlolSk31TGWiA9GPIRoNcvL9Ir7C2
x2g0Vr4Hs2nS41ImsenhlHyo+CnFvhg0gJLewQ6e9nNCE9pA0bmhWKBYMmPL8O+e
kzoI0+td9mHbRlNAZzUas7W6wiUNcPORFFwsHRl3Neix1NqHbQRW2mygNhlh7zcr
zpI5WeW33RO41nMdMaNDeUoMMxerWALbwsri+IaaIB4Yp74y9kruCC7Dw6V3ZSv5
bddLs0iIS1+qujywRoVoHu0y9dPEn1wc1TvVFhcozGlxLS0SSJz7fWTMZLjOojWY
lYhaMWzg8fjL2R3NeTPWbvB8fRFMF1/aZzAMGx2+IvpWIBd50O6KWz1OTl2/sS1x
exuxFPfbkuEGXcEqAIQEG3SpBoh0EZHhDVxwgzviXCEREKWTS8bKzzcWG2ncXf9y
wrF/8HEc2lqmbbX4IaNc36kvuNm3eTfD1agPl8TJ2KhagGolNI8WIJujEbXiMioz
yOwPZs0v81wTV6ZnQQdjFq/tQQIm9gm9jknQ69xT+DshvpXJa9RaKbOhQe0u8iiy
Y1atSE2YHeHQg20H3bn/+Bjz4oiPNhFHKi133j33+WTBSok5OCB1x+HJsIgliLKQ
8LN6hG1sdh9sAJlV49O4D/LSXPSH1iyfcQ5UkPGekugrvC/tO1Y9I3ANWGRo6lYS
kEAlgqOJyv2ilLSkyqesc9IyqCulqtwUF7GcFtCXN7mVGpkJba1tpt0ipJGDod9T
ZjBQoOGLUuSk+I9U0DwITQDJwEPvo+AFa54BZK+gS9ecBGVVLd2uDjCY9d3ps2M1
yw69spLrjwAwNp2+rh4Mnl02hNvw2TEdvDHZ1rkYNRKQxHluvlGpcod2Y1A2E7Hr
ygk/XrxG7sEs6wPpa7FyK8xZn88qhpmFOl4C33P7gIyO4pmHz05uz4LROM7iyr1x
4RuYML3Uzb/JOYHDt5RwPxIS3AMtewqj9cmr5YS5CmfFDl1cvYtgO8VK+vXoAvgv
lXaaUMQnaLSj2QpgtXosXG/SFVjts2kYiCFSekiY6YoywFAPYbyywL59Z7rD1gyt
PWuyDfC+G5Lb5jQ5cSo8oAyWQbE/Spj3XRASsju5D+IFXogM/Ovox/sLW169J5WA
38irFr/oD89iaTxnxsdx9OCLKadnCd0oNjVo/lsfe9oMU9r8KDFyZJ6bdtJnCvE6
YihJ8YnqaeIwPxJGjvygT0UEJu41LMpETdCH/9MnJbpVgbSXt/S18ftmDdfJiAMO
a8wOHPkwAvqv625HFc4vO/VuZw0WtBV7+G0eRZxYCPI1Qesd9EY118pdE9u/nn13
p8K0EEqYtb3ulAzxcxGP8iewSNiMAc6x7GvgBzY4frgh5W7mH+RwpBkNX+CZ6hQQ
+IPk4LvUs7oiCYnJRYPdzt3D+WfWhAT9kK2aWTNjhjucpJQ60fvvBHgRJTCJi+GR
CiFKj6nnC+gAXCCM+hv4zEToAAfkFMQbaUGKEqnKMTziEShKO3U1LQ0wNpr/FHZZ
G1JyicYYncm6UfcP7TxsOjGLWt5C0PY7f2+pGYlNdf3Q6UXC/rPqJVLLiStV5rlx
R7Hc12bamokj/sVwsXP3O/mm1fTNE4KdWCeTD+xyMOHYUcs/uIOYXf6YWbvQfwn8
bey9hCOZ23Yc8ErPP3uH9lTPJanh5qwxSZ95dMmLFc3Kyt7QRnTkFFkykm9uJUIB
6rAF1vpDVUI2f4lZlI784xdbl9FNmTbn7Z+fxBuzwpae8+HG7l6t5cpJO6ntTt3w
VkyPKUMqqbAaXHejg8W+dUh33mR9AQRw/JuZXtzzSOlBOpej96OztrNYEx6XN4Q+
jTxTeVbHc66pZRltE+2j6kcz1bQcFb9wbcndecHOoaWiwBOmWIDdwThBgsR4sgjL
pdvaO3zXt0Fbu3Q3L6sGY/ZW2Dhp34CZb5vUILEFE6ppawJ9m08iapDoOZR9Sx/w
Wjj5C61HVsnfU3PaACxnncJHnUKZ272nlopeLuuxNzVXgFRuvXqbbPYIyksIHJvk
bGAK2J7XukE4c34FHeOsnEZ/vwR4kOoi5npUE6G0burGkEJUM9j7jJciolNJ6OBw
HDPgDH5IEYH7elw+svBZfVuFVvP9+ptwseXQ/zFGFLoZOyo/rnnYUwlKSumHqg59
fWkJNrGmVa5G3inCCZ8BmcMs23HwqZ9+AgosGYvy5HJWXCjYtYQTSM+obRDDqMyA
/TPMiIyon5hH7B/XCP944eozS3s78t2eTf1AhpfAXsXsaQ1kRaeTM9CR1yoc48VW
BNdb0Z0LylrHqHhGscWmnJfu7WNzf/C0PjLLRI3gA5rYghIGQgWlGm3y4QuImTKu
jVb/HPYuapdVbfs8++9FJXt5P7LO8fvvYy6ikl4j/nw0ZJFEuvRV4bX93EaXh65p
sn2/GBCkcJwOMUCcBxJPNl4HH1zr3g7uDRB7HmZz+k1i0aJpMOhJsNrx7V6+EBE7
CHVNiWnTYiMmi4ggTTHzZXZnZPj5qgaIvUaK0hfQfX8Dk3tTbmf0cm85CwfFpoPK
fiZHNhPIh4WcN8lnIhk2t9cIEcNTUYynFN8bBNFYWqQnR8cLbuaCe7t4+bYTTAFb
GOWTqdhnSGrwwYqou6RBgslcEVxLE8unWeep0RKAOWXxV9EULn4krLT6SepfOjuL
qfJYGIJOWcqF7XaDh6Pw+j7+qR00B0lEW4zlDQakouCB8/e3EPDwpyDi7Ho2KnEp
zwzArZr4AiSff/jPh5tqzWmZ+0OPOUJGYmwI5qiV4wDZv/UL4kPkBgMO+CMorr0u
/4P7ifjyKT4qf52C4W59iimcOf1n8rQyocT6p7c70UWG+dVxdT6i84gbfPU1oMQ6
yKNkBKZVaCsbvhfUwsUESAXeBJX0+PBk5ZK1MmepkxM49Hzub+Oihf73e7h32UXI
Peq/66gQKXf8dQ+YMJQscxClP3lGXSo1MdRBCW3pp90+saRBVbp82eoOfgv2pDyM
4mYfiNZcYFbYtY/AHoCJR6aHIE4F/N5B/wDZfDQDywl2Xjwdi9Wx0IKo49KwgetL
rN88lVcg+09qFzkUvuEciLviNC/bRKr68Ni6EfBzhxHtA+ajIediyYdhwQuOSaeQ
CtuvDLVR88Xfzr2oMNFig5Ndw2ZJJ/6I5kH+K4lpQzGD0JLChj1N6+l4f/c8XLBH
lyaVL61hQrf8C4vKlUaIlD8FwQgnvuO/zsAjxsplKprvtGzEAqD+Vj84XLA1+5KG
Zuil0LFjmaXtpNTnyKFtu3KRU9XcyzeZlihXiK8hHyhh9C0KGAT3d5oAyvs342Ho
k11m0zx6F/Ic+Dv/pKx2//Z8bzqwXrHKGwkHbxkxKT/O0jaHWRNKTi6lSCko50M1
bZbln49uD1Wfy6b12TCrbJJURTyEgRfcHS8ABb6gPwQZf1O/aPA0d0hWS1WgAgqH
4h9rZIiC9vnaG1VzX9R7jN7YH/2Qo6tIeFGxL8mux00eI77rj/KpNpgdV0ZPC0o+
XUVx4UeF9XI5ERBNpXg5K3w/h31HWqf8ui/W6i2OgTCw7oUsN2yB+4jaHUyZgYQ1
4XgSXtF2ggSDlTXEjYouGgMZiklhhJwQPypzJ3Mb3tL7uIRBmLN2HvK4rAs017vK
6Nr+hBKV+zKpHcdNz0TAL2Ko2FqiSi3gxo20A9ly0mvAvUFlgzqkgpudeCRDXZDv
Ze+0wrrX8WkGdx72Ncw15nE5nQKX1vdG1s31dbJ0g6kmmsvJvWIb5VuGdxJ3vYat
Sgpk13OohMeQMvxlnIactB5WyJNQY1cyon6HddgDNguE/jY9cnU3+jpyO7lTRUuK
/gWOKqmrgOjACWIgq2kHz+xUE2/wxUseMFTFlqEmcyUu0MJEYkHBTj3jf69oOo1d
wTbOlOisgsbaLLVMgZ4AWxCoiOIZck4hlkFaBuqW+vHUZC5y5bsyL+gd7fgaUdOa
yL5vavW6l9P/wdXHfyXgQgoodJqKJMMttLSFfJsLz++egPvcX+gs5JbLJc/LT9cP
ZW6n7y/E5+I86DQlxI8XRFjsB5uL3gRgurFDi5y3OfRwEzKZ2ko33Tk5+LauNqDH
jqS8Hbe/KKObXU3y6ZZ3UTnxlgD+rjPEIFmpVeREcRFlSusUx4Vn/EaOgM42XnJ0
fGWkKqwVS63iSxA9Lxy+nyNy5I81WvXz9nOdwwQmiorjrhM/NB2U3ccK4D4yNNvL
X1Xms1hzq79MQTqepRpgXk7P5eLBBXP1dhzc8jzM1dQQL5TeuaeAsiD/yVbHI+nI
L35aYjhpWusFyvs8KASqbzkA7ROgSXLrGLLTQ50HoXmmxNRN81DI8h+Tu1BXU1Nb
8x5LfvL7IDrv2GHDzPcLRhjG9P5/G5F7wRSrnnsTBoDmsyL4LIf2QVhGDYMDyPsG
Fokl8mZawFb5+iAVMrCLSbyQXW6uI4K80DwnCe2NBuqNsM4XlruWaJUAkB1uDydO
Dq1Q31m+yMpA+AFZoGfey2nmYl2Hr+DcllY0x5Alm5JR/+2cMdkafy851caYHAAp
wEwi3sUAOIj5Qwq16O1e0xikheKWaGfd00HGuNGrNWREPbDs7hFVUDgHmdCad1aw
XsXqPMeGbexxj4hTMHp+DDwVZPCbU9acHW0XbuQscmPua7Yc0rJ4CYtE2cEJNhVc
N/us5oiMU9MdOWeekbMK8rbGIpmpd61ab8Hd5sCHZTEve/8rqsEhjlD9CH1U1LKP
6NFyX3hN2W+YS91iLDOR4K8673sBkdsJ2gQNl8j4n6qNiIV4aGzIOAP8TQEMAO0j
4HXQ9UGgykreXmnklCRQjx48N0vTscpuPatAg9bOogAdvSGFn8Zo8tQsl4z/Ig4p
xoamHoKyLHAOUH848QWTtcWzO+0w795itljhiiZBqa7qHshIXsOjrBJziYJIQmWQ
1cz4xecIC67thWm9GNz746nViZCjW/KUfnjwux/1BNJbnImDRMEFcilzt4PxHdHB
Coe3iOGfzgQiw1Id56M7vmdGHq/6jlj678gJehpbEBY8ZEzJ+4eU6lLwWctJTEnK
Vq9gDWx7Ut8nRwvY2pl8DIadQWqqMUhiKig4j4/ZJ38gD2gnXS0lzf0Yyq6drFFU
JxNZFt73/JNYchEsQNnnDczNYSkstt8pOeWh1kntou2HJgo+N4eQkqkQWas1pRIr
2XWlcPXZKc+Mue9wPdm9qm/y58A+ytCMM9FPYO7Mdr5qgQWoQZ76tgz1hCtzLtbo
wRFh/U4RE99O2xDiE/baGxr/3y3rQt5aHFwG9pjLYGJ6JiktbXMS8G6dZBuMlizS
S8cf03Qu5Ax5YiGByj0H2/EEO+vtSzNoTo9zTwWDPEsbcPXL9n8NqeRlTvwjMI+p
O0cnidNqGuFO+KIvWwQVKHNiRQfei2z9T59KppEW9B+yi979OtYzSfcoLc2Bt7nJ
E5DY7nO1g2UavTlkUnYNU4zK1cVR45Nr4RTtb0QHax+dqmc8dIkMYrpR8kNwSWpq
uF7T185bgAKWMa9KKiVTxoMnQss08JsM18qufd5QQ7fafQnvpWwuE3Z51j48UiQn
es6+m7RjwcXxkwjLylhC1qD04luhg1kCHVvcSYJT4z1HY4Mz1JTYn/2y/B+YDU4W
392ykU7s/MLKr7zL1SdMxA3aU2+/wqG5POVUiLB1XBp4IM77Nwj6xy0H1aIItgC0
+xsjjXpoiK1LDFV3VNBMuVQ5r6e6lMvtFwqo/AYsyz2TDg0TekrOD4Yx8pQiBHis
cENBv2IrIzmbu8Ms4oxT9/3lIkhrTdqSnSNkGgzQpqdchxWKQiApSTCBRVDPuAuJ
vVSFwKjevbgkgD/M3Nyg0xEyAVBo4s4XE1Ap162P0wP+VVlFaC14IDtdi5heqA9L
jDfdcd9vrMw7X7qCRVBkn7n+MC5Mc1O7yQRU44EcuYHWO5RSenhK9SNZPuyuA3WS
7TTcHdIw6rp7NeY2H3bTknEakfnx3UAZan0uo5AY8aOK5yZoHfsGaUFJF8oWXGRg
DLAkgdl0z6K+H640VBeyIIiIwrEn0/fUoUveQE5wV9w14WKoeExwffx9FJQ0/uos
Q9K2QoHR/9cMYXsJkcKDA/pQX+z65TjZCpfJ0CxmpU4blv9lScuW/px5Q3JKyGme
BEPcQAb/7uFHF6nyPZupWScCrDPIIElW1gaEooVsbEJ/T598FtAY9K2SK1WgpY1R
BK5yf3gUzlSW4psTZRwD2F5H9AGx7cJLb9ts81zLwpV17zQG2tVO++ZGmXZEiUgo
1CYXvS0ez+uq6LmmsUyRKxsR3ccKcyvenEnwaMaQmoPcX5Z+xWyGWkmKX4dIDTUa
1WQOgxy7RE6Gko0huBf7R4rl7nYocmSsEzatb8952hTHYhY+6+P3kSwMtfQYtFcJ
GtxcsyZFp018cjpbKibw8YAJr8FgEdoOpL9EutTVKB8IUl/zzqaefwRcVFy5U9+x
8CB2dCg988iBP0Wbw+eEegUMFV6mCv6SNynKwadLUOzHE8Nb0kAwNRwde+mpTucy
pEbrtR8uz0MFMzljD/RDQ8hjPGXBPVWpk1aFwQD3UbDmpwmR2YRZmC/30Hk4RaQx
Wws27yy42i79zEeGHZNECqLcg0Us7HZx9V+JlHb108qnT5D3ysNdORydh7mMlDMS
Siwh6yk4Tlmsw5b7lq8K0jRTDQUlzXnnnNJv0O2VyzXMQ1zABtarxyoILcLnfwHZ
+R9N79aD8Ud4GtZ2CuRZ9D/xRgM+dWE1bejnHshCuACLpe0njv5sFb+tUfO96Bns
4lhR3PXB67EcgU06B7nK2LOo+Ds+kOLn7ipoaO90erB5ZW4j6jdHMUnWB5sfX2Do
PKvFOzMKxQVqYJuQopnjBp2/dT40AJOmkzWHnm/PUE17D57IaHUJAQUvUP1QXJq1
s4KYpyXni9iuyi0DCoV8REQYpwwHvx5cD6u/+kJ+GDaUa8A1/KAaQFXbanREblDK
mu5ikrYXkR+/WxINvFqUpuA+YaEcFCrSZ3+XMQjbGbmhGsjdiWis1jx3tcGMDv68
qieyhd9ocZ0+6cNmlcvLeQodKjBighRdSN5eQIrhM7jrU7+7b32FyM+iUgt//bB8
TQgI4s/1/XToaoVSY4dTA4LPYp/vrZnVIrIz1G7M+shOmiHL1yvlNCqrN5FZ5ltd
QMvWZdYmfgR9h0sLS76dJgYIXwGasEtghpXvc/f/OFxF32nEZb0flAaW18HuMjdT
/8gFy+zlUhmHMHBkua816hnr8C95vlbs2uRxDwq9ib6UBzMqgWXocFPOUm/Qwbai
5/HpjA/YkC9edfB9s1NNB6eYmFhqk4TH6iBecenYDjl9Nj7U4SfwMo8EtCzEzirc
uglHIHGbyAMiANehvlwgSFLdRxoywGm2ISSxkza1x1tByfvZaRnv1Tj9CbIcFLd5
00bvYDzXjZQrfov+WcWJs0dMaOqO2oBGV8G/AhJtfEcCqgdeT4b/xCcg9Tcp7yM3
vcV+qjJc24elzAIrf+BYRMp+eakAGiVzK2NkR2jx2PBodifrOCYTIlM+mirqG31p
itU5wOKTO/OKiGxe7bv9t8RCtxL5mc+MPIVSbzdD/9cAYu1SekVMz6k9GDmGnWjR
kiDnSgdPpradRXYS2BWpcuoPpCfDUQtxcTxeDKkKNCeindgo20WmlRE9SZyStZML
de5K2EFjhz92AZOCYatm28ky6EEbb2vaCLY/C+1rXgHDI1xExc9HqaZPVmhRKM5z
BfGqSSgHzPTGS5spWMwXMtgycpDY5BFlv1dybjSTck9XG7iNwKhBFfwXNW7YzGAk
+AJr/XC69NRm1eS18oFsMFTZpN+8q0/GM1Z1nhKyTeOrLw8yaGd06hEHN5fSEI8e
48iUgKWYRuNQah2EqIjMbmgr4Mdy4Gde8NEwtPplghMbwUoltRaCukuMkGIpkKE1
C3TzbJyqVjE7ABR3iSfILku5aBR6Mx9Y8aWB91nHCM0WPTHKfr1p+2ioOKcNy+C6
cBivyMZWP6BpQG/F4Yhtu76JMZVk+S2Xr1jcS4238zy3d23M+eGfB/4oM293P3Xz
jP1IjWYMjvBbq46qQ9ilk+xZvgB2SbHQ2DEglt+PwyWikO1r0CI3J9HYgLI0LjSm
Km3EPPceXHzIFLWn317V3YPziObUomaZpdrZqGPA7Pxh2q/Gl7OJB65Zwi19SAqO
pqUkDyybaZnmdhyuF/dryb4TOwhUIRH0oVo541ta3dN8zMjzIxnTEj2VLHN5REN0
TuCHDtYp61LJBoueakJEdM39ItkJiJfM4v4OUrXgtzgiEmYUWAt7N/cv4BnqQVw5
ufA9IVCQNeGo/RjEE7gDHZ4GpKTYAX0Y34zj0J7xBneTumVO7kqKa9sxgqNdVBEU
eZkmJPwlzn1wpXHK9ML9CsCY9eF2MCUO2up+5J5yjjBFRX9G/bpx+b4NKGV5b0Io
lmRUsHrXDeXx+BMcMiz8Ty3V1I5rIg+tZOWtHgBk2p3lDlJe2w8S+5KL9dCxrQem
TtuoI41gq2+HS5EPHB8nMFhUqcvb2UjGeasBUJNebY2aGcaTxKtp4RcI1vpnHHqh
yLHMkLb6SZpD8vd6vN3ptUeVPwXnNLKKA9K4sK+wcVccv3YdzIhBP3KDvNuA/YJO
UO/zfDT095KY7mFvhr5kF2hJe3wiS/q1Hl40OGnQu1uwRiPjoHJrHqOYqgWXy8LB
wclxy69AACrmDIuZ+TYgF6H8GMMI+POv5JRatXlTgwokWwS2wSWZCaK9CbM4EAMV
cwvJa2l0kfLwZ5VEb25+yB9zfWHLwkWliuerSaZCYIMkkxkImrI1Uumy5jaj1TJe
gi/JUO2XDISWDKtrTgEMZmhOXaQ0RVC52UjEh+rO9v8yjizOHmBp0/1FYdYmEz+4
al4nLkWEoThBClPGTjusRzRvKYCQx6enYy7HSnk/tif0A3dkhH8YVRU/HKepd6gn
4hwYvxOovRvAbR8ue/YozAeEKrsXLqkZ6Hhhcg5GHaMkOqIK+u8zDzqIk5jM8IjU
jOPSHdSuQ4/C0vQolqCL1bL/+RvI4V7VKIlF2CUQYWhdALRUL2MSyCxafBolES6o
b6XzpL6/N0AtVuY274x7RtqTNQODmfvIgx4wR6/Ri+7+fVDRO2DTMKETsDAlaTWe
fPRHBtaStqaW/lZ7/o7OfzHhJequWQhxd3uJzs+TH5nrXwdZMeG1MsQpKphywYpN
U/Y67HCSgR2gd1AJ8nHQuDIJn8NLdnd/H13gOy1N6wjlNW0Vh4IaD1ibbvzqTLXi
iRb8a9S0/dtgcGFDUe3MUTmhlL455eRLEFM683TPDKvwVaTrH0v+hmjMb7KS6OGq
jUqMUjr7f7YW+NIzAMY5BWX+dZG/XX2XVPr9cdgDkZGYz+6YyxSVBBpCew6YaFqc
drxPUBn5NIkcu76q6GIgy2YwOL/go5obnRr1QQlu+0MQFf8L7nmGqoIcp92BXrAr
RiXe4SydmZhjIEB7ayd0yb9m8QgrAymudjTJ2QjbIVv1A000mHiA0NgE4W8Pmr2j
qFVKdtzYwSUyYvfiZ2r8bCziRrZ0cRe61IdJ84sNZluNiml7iZkoM7QGdv6hQNqc
LKhoAGx2i7Wqk5wB7ONVWbc1Gb1+ffErQjuAGWNeXS8qRA3QrioQ3R7U21afRDx9
5nuaKaAMFcdM0N+pqgBPbKaYFq7Z06C9eUDfs1pzr2VVPW4PCaiwY0xm5mxKHZMz
jP9T3ybiJ/mz97wtxarpzM12SjJ+xGmM8J7etpZNYvfBhy1XPwqyiIy/ow7r+5dh
/HWxm0+UoIkUIsS9sEDEVVxnUAjfSXXC9Rbz4GYEllYlCve67v0G+SL6yVYvmrux
3WZBb8LZqApDog8RJxCKtJoWgqAImooSjYSg2K4Rm9fTPVXnDEXzaEmf34nN2JxW
5AJ4bbwlezwkiSKcZLgoLq39YxOQkfh/gG2gUSdW4MpGWQccR2vJoDY1aq9VPT3M
AglUYwasPvTB5QEUTuJ/OfgLDI37WYO0wD2ulaxsWyek1BUMyrK8QMoyDfzMzzGX
QTpL5hT0qpciD4qQrSPq2BUUeWGRwGiEt2WuqljP1UN8KKchqv5KCO1ekBsKWTSt
rbtsx1SpFX7OwtOtXYRclzkFWCiYg2xyBUbV2tlOImFuL/DrGYBEAWWIlmraBSjy
/6vdzeIwtuK7klhHDRNnUO4PYOVkeVFYBw1LuBQE17lsuDTK2NPw4s1Uov5Xqtn+
vhXuuPtz1jKjzMJ+YCgObAWou5UO9MojL2bNKj6DcLloUCAHc4+f5f0yEAcZKUq0
JnWXYhC5P7EwXLitaNUmXJAKHP/QHk/LOkOiQcA2ayVn7RAXFYo4+xifWAM5ann1
x+Sjg4QwIb1PTuuxFFR96y0uewNNeJFlr8+8b0Ax6fQRi4+ZmYEUfERwiaiJ59Nh
Z7e833tW8SV67psIFEaf7/KOPuHV4j+CGh35F7Ac7FqDC3bi0v76U2KQptb85vpy
MSUEB8XevGfYl5ylY/fYXVdeW80jX0LlAwpgHgdsAKSNxGDHMqjcbi0WDGyEj/xt
4kf+m5i0JVZIbCHQWCsvN/lb7xX4KP4HunHGAfw9Bnel6m45sAXvupokuUM+9sw8
Xxjn/N+yT5/YInx8/gNNcZHwlhruf/xzpcH+scKan4XK1Uz7Od6QlSVUpt8WLRPN
i8t2h9TEqBVSXaT6eTPufnMrCK1KOCVf9PBESKBT+ovrJRjDDmbPGLeNl3kjTPg1
l7wOxx1H5YWRSv31XsXU4M1syptAj/dtEP6ZgF1JXfnSYpUqtNvJybB0im6Nv3zy
EzRo29c+UD5WArUEezpxrBLlYAuv2f5wd5phFuE12cbFafeWAXLbATvKGQpoEraf
UX0NvIV/s5Nf8qaVVf40qGFwc1kCdm0DYyHUdTkrmzPx95jQwm0fuOJYde1pPLzv
Uort7U5j5eoHYP9PAa9eWieKre/ZuLeRCkm88YedXsld2wdH7R5XRKIjePOnPjPJ
Fdu53YauGIkRmHdzpgU4WVDw8kZZKLtzT3xB1mQvHnMigddgkXj5igsgttKU8wFR
BZTrouDT9bQUok8MABEDnAXUgXJLjl2KM+sk7jb8da04OseqC1onscC1DoP0QN9q
kxJci9AvgVfvA0Gc0hwW5riNhcGztWRpnQKfSvGi5LI002vx8OA3cnBotuf7Jai9
HKR9iZt7pROiOlOZg3U50wtC6m73HZTqiNctWB6U+c1ZgWXmc3xF2YGCABCWU4ix
weyG6/WUtzYMurBh9YLh1STTZ0S4f3KDmtMuphine8VeZTeTVP05C/cv67tnF1Os
RHnK3O+yTaoTm+3mBz7RxN/NWEak+95V6amASx4lkJesLDa4Er1PtgwnBNULeH5a
6eVrfiL+dgsooxmwMhZblVjcpEBns7bOYQrRxkssqMifRTumIkUptly9xlNsLvkP
0D25D28jAKMX3O4NwFkHZmXS60DjEuiX/Vlki3LM+j5GGKBbhXlu5ljxbvFJ2lNN
Vlww9sJ+MLMTqoICWZ5dtHGNiDclX+BVMwhhqnPWAcyLUsIesk/qA8nuMwcBzIYw
71QaVasTIuWZBm5871MQ/FdMiiVM0ZRwLQowLvdzPQObnfA2ucsHg7/DU8zzRQJf
ltIo03FqDV1XcBuVGZE9UAlSOeG7x43cYPmUSN7S7C2mnd5crhBD9usNGFTiug9x
t83WKCWS9jWDHn5gDlhcVHyGH8swvpQm9tg5Lu+zA6IRmnUcdtnsKu8jljXEMh5q
jffwyIReB7LeDYOWIo/qds8uPRuioeQDXlp7kdvlEKOgnZXXY08SKjSOg0JEifE+
gNAFOk5T+8Zu5CdcV+buRXIFevTCCaJevDR6uuLgtecr6vvgMD2+lFjxP2sxyMvi
n0FdX4wzMOrtoG5tYXv8dhVtlU46oactGjzQwkh2XJ0llwzb2KQpXq7DaZGvfrE7
NK6lNg28U5RUPTRMghiKEg0Fuusw6eBZXPjuT1kQe3geuglAgymW2V0vX4xg1nT2
cVKlzRR0bIxSIzobHw5U6YP4pV07AVtXwoFnWREUJKU03PaufvmeRG6+yKEtUqib
W7lGKaZa62YSiS7kjxyIDsuGj2QSjlYPfOH8F/PJ5TpgWOYsX9tkwYLeIzHZk8CC
Fo9RMKoWrLG4vWVctjybsWj89rEcusKzM9fAi2oWfYeWTQ6FuBs0ALJncRJUrh2G
jehDy5q4WyUzw5e1AvdmMQcDV9SnJkvara0CnYzmOYOFiU6pRutl02hqG3dYS3mN
Q2GMOdMfJDQ8gSulIPkpT/kaMTGT2e2horCNppgZP9duZu/ahpyvZ+DoVlgzDH0d
Jv+Msu5grrJ3Jz1FlVlTpBvWbj98Tr1vLiODl+K2Zon9WRA8KF9Ebry7TtCuUt1s
kvD8fI/gAimsNoA6WNCbtgbNRCbqfKQCYkI9S9XEH0F4XSam+a/ih0pc3YtHFSKy
O1MMcYviW/xrLByxZZZRjn0IXI5Xkj7QQMiSayFeUUC5Hlzo5DUmrkJUArEL+tD+
IQrPi1lcmtowf1HtyJeCM1loel3KmNDslvamrD6YdU/VJYCloGUCmhZKkvoAuWUk
kcl5UG2fXXU5EduK8bHHhwuWSHFCbUn2o3khSnEcl6VMn2SN7q+MdF0nQQrlJOd7
0c8ov79HUiK4xhQdB7bIpOI+I+SGh1BGmKWE7REc6KO7zrA5FGI7ums7gEcyVKdk
Cca2WvAYhpifEPhM79ETmM/hJQVN8OrTEB6StvirV0Y7JiRU3gy3ngh3u3Rn/f0N
1fq3jss509esUqqLHdA6IH2mbB3JVASYIEWiSuNqxI/hekYNMyGuddZPdWs04wXy
H3sfvdlkphykODN54x6nLivtW1SM7EfFD9MJAsIDz3/lhhqCDYCOHmUqqo5Z069n
WShRei8ujVHZbPk3WyUUAYGmDTrixYLS6G0xtlBrJSF7rRZnVGJokmGmO5Phha02
vM8oALt6ApUzl5LXrkuIOrFomNfYhkoFO3XIx3qbcnb6X0nPk/871zztkWErAcAq
gtXJUHfAFjME8lk/YGSJdRjmoxCafys71iXB3VT9W+jsP2NeNyKR+K159IPr7MmB
76fbZIzF1VH6bwyIVX+DuTFTUj+ptzNWw3vZKqKHVbmUIgPkl1JFZJvXaE+OZG1S
ONiKOXbTHJepV9/pRKMV/+KV4H36g0rmZ8R0xWPZQ6ab57vyHupkUYcxWhXZ6vta
W4RBNVAYjYjujaxZiaQn2or8vjKaXsOQ6+WpgJTwcM0th5jeoMvf8LKI7aUCdKt0
Y894CjtFLgUPElPKV8fJU54ufJeGV8XlBrqp2I6ue2Tp8dOSWMQFiiLjuE27spBb
/df8jOkGxlwevIlX2Cx39a77i5XmZ4iVm+TcKSGjnnukWk6aM1P8tGX7pfZYzD6O
wU7+3HcRFpOZCkVhGe/7s5lNbK9p8A3T7WYKlAfzM/uINMfsABsN+QTkVXQr8d1k
LD3TnCPjsxCO1bV9/hZL/rO31BIFgPdK7/Erc5Ec36bYWa9on7HUYDV1e54Ld9bJ
1sb9mDXczD4rtsWxMfa6heJzZPSgJ7MjQCY+ZSt4fq/df5LSZL0JQOKjkhoE0VnP
cR+ifglHoSIg+XsLqVLisuGOf2T+Tf7aeUZI7xGzHvHrA4DfoWtNm4hYzYVNHZl/
HclT0CLEDgajwOZ9XFoxbhBrnxx2jxF7J2fyoFQ8w9WZEF+ZyYfKyOd+JMtOL0uy
ALBLyhde/sH0hiiaYdQxPePhsX9wHPHLnlIlRUdsphu1hB/M4cT2Me5FQanGKjF8
ZRYhBkdyRQg9WMMGJwuzJTIQUQJQPs1lkmQ4Cjc0B42A5M6ttuqQp0ndOeTbnJr7
OZhhrhj6e4SjkVsLAd/1zI4OGSJG3CokThUBnxUzD7XNqHT57BXgautQ6iW7CkIX
o9ZPi4R9CC69TDY1JgW0ixXlxw5AdNVF+LBIP3OE+dUyorOEhq42piodE2jCwa5D
Luw1+CXuHznJHLwiyL3dNX7Wq+vnWxYjkQrKjB9RFaLVFAh3RmELIsOZ4s5Z4lF5
gNNh/eJiTawCBilf22v+yWhbVITfFtEz+QO/OcNl/McVNDWQin8KdNROY9o6BaK9
td9INyV9nX4Ed8tbw407iar2TgREWEmoCIILQB3MzVI+ld8mX/gGcf8l2gECsnZF
aaytKr15tzlV6kbxMUbLk5nhqB99AiJ2IEBAGaggU/CANqQMoTl1zBmfu5xuQ3ZP
8e0qOOiXDsFcQeLnKRqqKBCTTIj1GhMWvaHi96wu+CVaPl35sBQvdeAb/sYE35/d
NTGyO94H3sdN+xvmcb2XlWnp5U1Z8jbLyvdjscVS2AECk/bL9x9J9tF4F5qS886j
6NHI+U7wxBvcPZ48nNE4GRRtBd6+AhFWQH6y40iz95CuJ8eLzlQLA4Vuy/KSn4pz
Nq/ML4y08tsqtQC1LXMijCAnRCoQFdnRnDVkylV2HOxbHA1vWQYLH5GitIge+Ikv
sN5n8pNKPN51tgo20C7DjBO0QGvWjqI7jQg5B9ZWNaWCnKmWCa+Ixs/TQTvO9zKb
z3OP3MoGGGNtwPmVS/Zbgx6Lx51xCT00StJgJKRQTYpHd9uMBEj0I84Q/axaW+Eo
1iH789hFcP6HM3bkyXxwcFtrMvHGVZQWQw13zL3jR83UaxvLrxfS/ePsdLJQo4Jp
l458PGqdXbvDidqOSXCcv9ZiaXpLarHFjeQPxWXiuK6HTKapIkYjmsBh9ArhOd+6
RWNc7Ne5wL7tl+yh7MK7osCU4NNZo4+vELeKgCwq0/Rp2VH+hlr17Hi2xHSGFfZY
WdSOdmUr6K3KRPTXgaqDsmMonBr0U1PRGa7aiN2dN3/K+x+7unYuIY8NyoA/6pAv
jFMRqo0McgendDJ6aiCgegIv94cJU8WGpC5dTsCl97BrpYzTe3xE51EOu/QNWL6Q
lruzPVgQv9xEZHK2oR7d3IX8xSxMMQbBW2lkxZ+H4VdxcuZrdgPJmJeOje/t4EmS
MVZ4CwSuhnWGgdarUmsVbnWJiMEdDnjOzhxxfwExUDNf6BQQgAJ86mKa58ONXKP2
A5oyHZFjd1yrLNBZpHUzVR4GoeSLjqMwmjucrqaTulk=
`pragma protect end_protected
