// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ii8xJ+TDr0X8tUK+QIYkBiO6bmstkSPm7quoPi6D91rT2DJnXDLJ7dVqvxSlDsu7
DndD6Q3YHxijgkZEBPyWgp8dT81ekoOCf8rdjRHcsrWZjjChTeqbPQsY6xgvsl5T
hfCOeoGNdp1CfFp2tK8nmif55eKLerqHp7bWKBh0HPY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48784)
adLDBI7ET9aYhUFr1UFTkmiMMkFacEmUU/+nCrjYRVWdQC7IZJGDa3yXBKEElfDt
2+r0PoCFx+PzEXKUhi38ml48VtBkDl822IukzkORfAWOStbhJEgFSN2n4qb6P2wk
UpJwwFlfrdliFh3TfQN3m4buIPH4ovsmKPkL2rWHPqCN7wWwy1swowRChImBQEyi
57w09HPkg2Sz8dQaU6hUja46qVxfUE1S7tdlki7TAT5WK2Hi6SAR+bAphgk9MBND
ybXbYb12Wk6R9Lag6DPNnOZpbqy13XfI+UrVNgpxz0nb7LKvs2PDxWflufOjPR+R
wWhO7C/OXmtshwwM63o+1qN0JME2dIq5+KoFq9rfc8Ag3PNT1Z95jqlO4EcDeEkT
fPNnw5sXwEs+/BI8C4eQXPkgcJ1MHPqWwBg3z0XMSmyJFo9jkz74eT8eVhioyMoJ
rIN6Yx4RqwGyQaoOJx13opNbJEDWUe8ouZr3RdevnWLoUUB609jU7DSZpw6gCf27
7Cr0zzf6FW+YpirzdNLEswiJdcQE/w0qkkqlP7pzXEGxElQtbmHyS+e5nlvaoY31
fBoWJCSdhXEhhlAF3jswGUdCu1vzIMoxv5c7pmqhS1CTPB3iDZq8yXxQw519qf9T
x7wkQkcDPTF5qvu7Z3EqRnZbcPC/aL1UQRxG0Vo4+HlfuHhgYnmJzg33fTPEwQlE
lKPs7aq4n1QuK5mBUcSs5Mg3DZZBj1g0iVfcf88gUTCRlxyOtmXuy+46Wq0u3neZ
Z9EEYI9PBSfqd840e78XeZhI7Q8ftixvU5OIkuIBUVybJPHz0eEzNyhfOHpa82qy
iyC06k6fhx8JjaQ8ERqkx3DterFB9wjUjYe6lKaCaloE5NbKkVW0UjjKHjLMuwYp
84DPjmKNe4pSwVf4pN/X8EA1gnvmDuxeBDelRHPr51kNsnEBwjA+oRqsrQA3OkYM
ZVdQlB/0/ZMznAnodG30Nrck0RVWYfCVqKSg5yOhN3DJw/h/XzGp6ZzAN1Uf8Sor
28YzVAbPZun85m88CZNjTrH4vTeUyNtyVcscV559OucznGx5in+7Ul1EOv93PWTx
DQj5alSNqNJ+ORfKl+t4U81n7EdhKbu7/L+f+/AuKS5EBI8oe5X8GSNkbS+wYPNt
+kmD1FEaFpNBbn2xvnrSAVACyoa20pTaNqA0BPvBZpM/aXX5Dv7jbgsT9hqZxhHm
dR3ujS89beAnUIsVNmMixXrcL1CdToyfqrnA/JgVs/DnJ+NoF99bvzTEBEnnPWd0
Lpicw8D/JkmIwxUsJxvOOHNYrI4WEcs9dtLZFv/fFALUwkHKuiNlGdMlFVtmR+nF
vM08iMK+KNlyM2AaLsqSot1FgP+z0ewr8ybWKicuN5vN1VRiQThVklMlQ3Sa/LUq
djkN4KbVfUOAT81fUVPJGBXmL9d40nTXS1AZCqwuKk1fvQNAiIVen+mTn1t9fPbA
133rHUAY0XZ4Nlu6L4goazZyy6JT7/UThvvEhopVCTHeNKKzmA7RIHmwdNyEIY71
xbJbtR2619HrG/1225gvT4W7ksxeHUv8cyZJKi5D3P+obERwhGpTQpPQ65+xjxTQ
6WQ+0jEbinsWyfBbt/CCRRFWbPbqdNbNhPM4xUPowbkXjReqC9nARAbaswgzZ1n9
CNNFAnkMNUMQ5RsehjXI8Xn3/R7Kk5D0n+jJVpci239as/Q7x9JyYrtfB04kySa6
E11YAY92T5k6dJ7YDBpC9WI+bcVWZYwLzCrRGAaTN2b/MPNQwUH/qytiVbxb/Bl6
EBb7Zm9+gEpBucR/ZUcyzmA2TyRz9hxyHl2zl9XraMHLrm6BTNDGbVPQYBsQn0DL
R/eEJ1DMrDMfwiWZtf8eh1xZAyzwTmVsmyigmrujv/zl7ydttGDFr6duxcnd6VjH
qLAzxrdP6pCmyhrSRuLjJFT57L/6GE+/P9yeQaggnb5gDjaLeeTfPJENTa0sRZ3b
OksSHAgHjbJYtGQSs15fXRjIZIthqieksV1xyxfWhBTDEmsgukJnq+XMnEiN7FBZ
5bWzczP6GqCVENil1NnABLT63ytmJDaOhAi2Y6V6nAUo9Nr/SOvcEzj92Jo8ZTfq
cg5bMvFq0qms+getCYTZJbGUIWFqBkzDpqHv4m+vTCQukdPSfOZq5WosCosvd/OJ
Z7WcKVEjQ2rms64SxzpjNKjYqwH1VaGFeKTzl90+bVbGEdNrBqCuFdRvdUwOKqmX
oNpINlzM12AwuznTYNk2SeancuUElb/HeTRHAJVHZ9Rq9SPenPUSna44jd3xZQ2s
AvHjiH49TOHyuSkUq42m2iP0ckU+TuJ5vn60sIqLQSsQRl+E2wFsgjModSD7u+O1
nGbACAwQhq02Jnxl56QNpZIAs6HVLlEAvYnWwhIGumzhAYtP6BLAONcXQHVqGJ2w
W/TmV2RB/THZtUuZy5L/7XNwfC8rTzdzvwp7+c9BZ7+yA/RaKFuNIlMByI7b/9Dp
Lj6EEGsFUCVRw/l7Z2NyPTU6HtSWbxbjcsMXlug1otabQ0bPrjTBnWWKJyu7f2Ti
r5MkTzRVUFN/Nq8rttd5XM1cEuD2tyG9vxWpcOi1P+KQG1zUjyb/xkgaMoTtirYw
VGXHeYsKlr/n2fotoDg4oRHeVdH3ck8ew18YHULgpcRdKggbwjtDswSoyUv2PBny
h9D00VEboTrQOEPhDLc+9PrjvgsfUgcqclpK3Cjq47K00+yfcbt5FQGiu8NCsI/O
z2ydYAwC7GOWk8rVxAeF9SkV1JPNnlg601QZO4FXSvaewXQwmWhaScT+Yns3XdyR
9JumD59ey7aCUnPVr842+iK/7MAt9AeaYWK+LtFAXZjH+umbKLEoeqa7M5FQgGWO
LxlTDIJrOURyQEKtjScaQGMkLJo+o64vPOq5YUd3AS6D3YbLoV7kfNwRKs0uvdwt
zbdviU1xeX6jeqBuc2OJV4FsKlJX+U93V3tJHCVWTbO0AmGVNCBHjgj7aLB30IDh
roSS7rMaPACy212cRh6bxQd5GtqZ8OLzBvRYT72bhKl5SgWBAjIrkHh9UQY3CLRw
Tm15Kt95YuFdXPLg/HHvCRYNbgBwsqCu+Rqb3BuDQlzFvBPfwFDPVviGLv7gtbNb
V9J95NHC+lOORrMQDXVBBzzWe/n6POlpGRUxnX2V3+tyej+PlFW3GY2Bex+LWAJb
LaxYYUpyox3aVos4JDHiKY/733oNd0G4pmxybUKPCBFNEWmwyVYDZwrL3LBztO/u
uucwni6i1h0Z3UvY33hVhZ7jkI0I9OxHCuZpH501YtY0CfPXrhvgACi4leto1ucP
JVSy03WBHCK0UXGTCFMX7qBjqPumBAoEgMwVJQxwvnO5izCN97PBjfhZS2/Rdp6A
92Ik+pAifWsIp6uHKssTLRFqwiCHgLIdp7MMP/znXt0VMbsjMtDHdwRw/DU8nop8
7MIbpXQ05W6lNn5NV2z9w1DTpA8Kke/7ivWY2xn56H3YHdGm7K4qPwsGsvKWHdRb
e8GLYfC+/bgBkDE2YB9T58lqyuSmY7AdtUQPYxD4FDQTdJvSfo7fbjWzDr+IcsXl
U7Eu4gJqLuY9EVR9hggCmfe7Az7vx7BHUseUdWWYAlJLh1D/fW0+tWtUWn6r5xCD
g9UipNY+G1ssyfLLhhKLcNL9btfXzE7j9J2SVYNFfRmUqmQTzixiIhBgohfuRO9y
fhieRGCW3ZFNS7+eYlrRV9Y/Akd0P7btnHeQ7JOwzEFg2tWmfxf3gS6EHQ8Wwzo1
Q1heUkWXj/bPhhOC80iY+9JzAydpfzPDIUn0kl0A4kWi3Iu8oOI79/MYQ66lHYDS
bvyzly+KMx/zl5hBQBmYOlMnnPUjmJRM6Cx9/eV3P9rT0eByESW/PrYFJRfeRnN0
uKQAKm4XLrCbRMCPKP7hkasYXCdC6Lo5zN9dgvlNWL1q9d5OZw0sx5zFDFmf/NT4
5wPj72rnv9yywmtj5zKCjwalH27205A/qXBQY2GpNVhu+ONX3UBPkr21vuinPcEV
65VGN5KMcbmprofjV1NVu14oGTZUYtvNEZXEqTJu1VSSDCcrMP5dW2gH7n6CIHV1
AKn10H2be+Jz/vmq6l/qzg49MUrRMAlvq+IKzJW74Tcyx3qcm3fwe3cnoWFpieIh
J1xEBWDVHnTBjsP0dTtyCH67fYFbXsqPt+LwSCxoWAJm+jG1OJUPv4/JGfHvYmnu
/FMNlkOUnU6bCGviOHdw/IdQyq7q9g6hfK9L5YqIHx6oBvZIdVvlAops0c7g88Sw
RWu21vGbHIJ4hlytCXFMr9ok8MuIxnvQSgqrWTTx65kDDfz54f6cmNWJZenpnVt4
RwMRmH76m6e+m3rYuaT2wTnvyqkWKpHpBHJlX8uUBB2ZQnRG56a8acexR50kyL7i
Mi0p1t7phPfVgdI8hTBWhk3CftY69bIQIKvYH6coB0uk2RbVx7KjqgdsJ7DVWYuL
lzsuX5hQiO/UKz1F7xbUX+VYZpErvkd07JgyPrfqCYeo+LAQ81KvW0EaCbW3cUhk
MJfSqEgmpqm+LSMx/myirwlG/TH1k35EtpBfFRzrwF+wKKTvNBHmepylUQbWanUu
Iai7sdkcM8n/cyJ/BEi65zGs4pYicVQ+dWlinHr451m+wyQNSLtzR+NMIArMzr3H
M/5o3USMe5L40CeRWwFqATKmE3koRV8zaqkPePYG6f0eertFeRggwIexcdVs+h/I
oDrElyEbUREwfcKyLRJkRouYZZnwUq3L4VtVdgoEKGqOzaQmjimDTsDPEJ0TKPfp
uEV27WNpglfnC5Z1TD8bdzZ3mNmV72UjsGBwNa89ibbRsavoTIg+DsWysZpPlLzZ
GYYJYn2MMQPweBC5Dbl6CVqWOf6PNgyeJ3d7Qe6dp6tvhrKV6+nRTZ89i3tXr+Fy
m4f5L3/TC4HDd1jb6iuR854Le3NJZ7qNMuNANMcicHTDUfETIfzAcjhbKCRAUfkd
Q/MTy+JWkPelKpfkyFEDB+n6UlWusIhnfhXontU0R9ciK3FiHVUgskxRfLOK8CL+
VoKsWEERw8WsDZJS/6MzyQRB6bTNS1CMPIxgQVZwhMq2c55FBdabuPzk++z9P8uR
KG9lQELJlaSSBaa5RGX10RHdJd/n+nAbh2R0xsazxJcKvgmcC2+BRWUHTqCKfo2y
FtMYeeWZLUt6AQpB8LWPXZSqj+PZlF1aNqcKVcXySMc+4Pi1qdSfTahMupcNrWa/
IkioIJEkFD2Jgfvl0sAzvgGpsjOgn63ochxeThOBAf5QCJmijqwSNI8eJu9Vvavy
GH7hJbuQ7X4D934Sf0SwhytMnsX7xuqlroTpViV4PEXombycMFhm663jGPeywkDY
W7gYDtAlUq8YtVXAvhTSVzhv+FEs+AhE5sZwxzhcPQ6NvhKagJTTmR8LcujgYJY8
je9mVvuYqm5ZaEh6zVZLRcx0hfScMXGKHjpZ49ok9N5J5dHXzhrmozRVuVo3OvSC
disGi9dQBZZkfysMolGgwgYtuNADQctKoRLHQWyVnlyMh+FZNJShWtr1rZuBB9bA
yq7wfP3EIOY167UBP4lxtzfiuY20s9P2rtuczH8XeukWLhwKXilNUkWjSq6aOqzU
omQX98uRI77IphwG1J51LrB/sWPg6o55ROcuohlV7paDDdYc+YkuodgAouSEoUG/
irOf/MskDvvSXNQcMHDBMVWYnj9YlOMcXylXWBSNiD6sxbTICJ4J21Hg16f+RQCK
44gkAlwPr1F72yf9NQWXsrVwpMeV2A8Fn3uHxfdw3a7+rhGp+05L+Umj08hIFUvO
hQCpHA0nEzrRayt6/AFJQhmMazmNhBl0gfXX5ucr7q0MqW7OjOREzmJCeXuW/wLb
wotruCzcd3WgYDOv4aeFwuJZNE+y8inXgxGI46bCoGdUYyVUlyKhiTZyF44Sh/mP
Xb6OYtkLc3dw72cODgAtbzArmnzot2KLb6Ztbq3p72iOpDtIPGbTLxXte+k1FCMT
wdqYhxvJ0Zt5XrN5tZRjKaSEL/2u8zkTr01x2+ueUhgJgdyzlxT0yzqymVI4v6Fv
LiRFtUQepRi9G8XayrINBmLMryBgO1aF6TlEXxIIs7aJ0I3NcWNFAoOrZuKu8hP+
MVAWvrX7Y2W/gVX9xQIYHjtjD3PalsiKViEu2n2TjVo9JxFVfurErTgx0MRT/eyH
FJWAby3dR/K2YXBTVCS0d8R++96nOvTQ5nthmdTJeeRjxjvIyxPHY2joGecWSyaj
ZgljE7FUw08+3WlUhFU3FQQbRXIgJQ6vdAheTEUQj/DxdN4vD6N3a2JOVVIiEUIt
Xs91lomsJOYJiAduazzXZ2ZD2ZUJ4ln4+csO5+7cnurInL5is1xjraBdtRuwJh04
Je2QsmDH8cZrbR9EkCLHMCUMYQ5L6NB4V99O29GajU264OXdv1NzFXfBxP8Kd+MS
b3ypCKGDcnjhVSiJ8ha8FuIFA+c+Rt9K1LUyFglDxeML6UdK99Tq9UzMYjEayXfv
qs1BzmNgb4ozMgVS/xTWwViMiX0yYxWMK8IwbWZcyAnvtf06FaBoxy9GZn88pYSk
Bj0rkcpVJhfSS2yq+BKiOLdDEb5XfwUNbfiuwbzxAiEDbGZpVK+rm3E+MHgfJrg0
BiZ7eW0bohFVxbXVUK9YD9g48gTQx8Kec2kXZww16J6y6yxgwv6oc3zIdltG/6uV
Rmlo3WvSq2JLqJ/4QoeZQdyCZ6iiVU/0ipqgu2f5wUB0S/0ELc0dKOBG/AE7VlUi
1rfH/5U/3/G8VE1MB+IAHrB92brQQdHxoX14ljtxAeL2d2ebRNdP5+tCRSpKxFTc
JvbSyvr3PsMNDn/f9ewIk/IEe28BzwXzhayHhLGxeWVkvuYYAF5NFxPV5XtFcwi3
0TPgBUiLTfGLDTdqPF6pp09rBgbvCMlfAvACiBvSmxgLlQa+w6vNLNCHlz4Qexlg
MxQwRGO2OLV4tha7UC/LHC1cs/v2X42o8D9mSX5c7ozCtz5E6Uckk0UQ/bVaqlAa
ndRbnNnlRN5Hwp5VfWzV4ToKiCAPln7NpeZb9B5jXlN6hnlxSgV0pEVRr8VQUGeH
tf8b7R+v92fwEJDawQs4B6dHdWTH46MznsLjLRBAPNRmJDPYDEHd9MwzF1BopqEY
UY63jwvQAtkSIrbIJi6qdNAjUF1ck0ebcU+KwjJ5jeGRu09FsIBVkkeTAhHba3ZR
3Enf/eLVzRz/YEvvCrd3IucPYzdgyvhYxfbYzEAD3uB096YfSzPTuSkklNMFM2we
+ZFvzk/qqjcb3llw35a5/DGKuoNJbPdSn/Uga9ALqjQFA7Gp6q7AVBM2zxozf4XF
uBjp59FbObGhGwgEhAq0E7JqZznhW1UCHWvyLLSA1kAkHhdBiBd9qvnOVC8Xs+sN
Ex+VxSp/SC9OENwpsbtby/NfaM4s25lX9Ai0mMtaOdHqe+qkx7jhQO6mBjXKyrD/
tWxYOajqAQ0M+zKldOm+12tSZK5zWNt2QQ1AdNHL2kjkJv+svytl7OYMpyBQWXiq
GQVZnqxM5z8B7GXESCbij+0XjGbyJCz9frHl7LqHMCxHa6MwFMTLTiSEA/iKfWxz
SV+t0LoK8zPK+F1FUgTIpIYn86XQoccItiu5ix8/ZwuPCTD+CY/RdUXLEhANT2P5
F0TumoIJjhJ68j0FdJMHjBwrTc3FKy0imyefH2r9dHpaHSlvfzedaV71/emAXamm
XRUdGak+v6+ZY++gA3lsrbkh71OZ5ziXVPD3m1GQT1MgFX95U81++TM8yK2iQ5aU
XycwVZC+GRcE5NAwEdQXXDQ9+vLZtyzGzRiFdWrJZyKqRwD4bIjCs76Q95l+G7G4
UlocS0Y4c5MNYOk2/CCtH3qt2HVxGM8KQ/ifgJgSkDxykVpJSKQ2GHMV9S2TSPwQ
fC5m3kgOM06fY2mcskYvd4e8cGT1tCc1UcEf+KecZ8S232X3Ilw5EBYTOxc8qpBi
/vwrCw8RtMEBYjBD6z6NXtEpyDgQZ2Yr/YTD4FJNExBOe7EGoKRZUOk8Apv8+9Sf
znu8sYRAo1lHSORsE+Sds7uw0qK74/UidqyN/khAvCsRfvLwUI8WkDwjBmE4nbd3
jWxHX8x8ypEloq/uH5NrH9CNsHAGLFAn0I5AIDUYBUO16Zd6VPXYN/V3pJmOfGJ+
cdS1bODMx3r73HJLly/sCSJSuSdABxwLWl/bM568Vc7tpDYEiEG21//xkasU9htH
PJYifzL2hF2hpxckUkTS39TAOP1FgjEA73j6q2HjLmY3/zFQVITrZIvfSkYsYHqG
fbZ0YJq5kmfb9pW9CvrJBam0JihnMyecXuy4LEfhHw6opait+Rk3meMndMpSbWV1
33NHJUljuVzTd+PCBdhPDKGfAZ0sVEtFkuvmFZ8tJpZ0ThUMhn5T+Kx4aYICMWOT
0PAqUol5zZztHUQsxY360vtrKX0qIWrb67aq4LCtlv5LdzsOz1gKdnrDHnzJOBHG
1Gsa9IwnS9zw57TlT33fcJ7RlYIhuP+squQWkkph9fUihPtx9BJeqpyIpJMC70po
8B46wqxpqOPVpaYYJ80IFlY5cnZX2+9uw1o4XCln+357LiOmyPRqxYxWdsjRvwSL
3Uc+/XGDb02w9bICY9iHKdBwP6L9DjDx7ENa7LUlEpeZDmvnV0iRUFjYTPvuSnO+
AoSdwJq2sWqfjt+372lMZr/9CsIp9V7BXxokmG15y6WI54LNEgUdk2/d2GWW5HPx
E2AmBU53Zuczf6qybcDYrT1KBEqeFlQ+Gl54NSJLMfyPWwZmD+FxmhIMNfawyNgj
clrDAfBMNAFDSYQFIVcPsHImrQ8yzgKDmHihI/T5yNrJNwizi0vaBY6BKI8pkHdd
M/KsIoB4A2RQhEoX5DiofffloShuw8rXUWAKf2hSNCPHMJkDOHysBKWWkq6WYy+W
csTqNXNThMrwTDMg1ZKZinqqLl85LF9/1EcgfL2Zrh8AuB+evGAQF5vtOzoTXIYg
xuJgK0dv1yNflV75lkFoCMJ+JRuH8NFrff+EzBRypYtc5MVKoGVAt8DyEGPfria4
y2zegRDtSYpCP8vuTTyOpF/sJngKE5ihjtGEBEFFFAVmnCEQ9fqsbNITc3O3Jmpy
qfSg4JzjRB/JQASErL3MMknYKaR/aXr07Y+Qsc6pN55334rVmfeIpCwUXhGSz5xi
TGl/BeW8PHHgN66vzb6cLA8OG2j8h81Aj4zG93HxW7khMwMyeuPGLKPH2r0btqKq
n2Cqh9GROl5oar3005RsiFY/kvAPBVSQCkR9MyJnpRch2fpESdwBwpwqF9tz3gMk
Qm5jsdH21gdFi5459/ZMD0pLOuLT+lUk4u1TrxN+XhyLA9jUdrfNOZoMOYxxsQi1
/lbsckNMu1HrmqNl0pP1knw4aVvuZNGZ3t2vVY9Hh5Ir+/kUfCTgkLJOAD6jsLbz
mD+wiPFGMLaPS+nhArL1DBBUscxQmVtXRC1ZTEhhEDuxQCuOCdJEIifeghW21oRs
bUctyWYDCCBEz9ZYL/mUOvf8rl59c/FsopcgGOJ/VoNvmLBRw3WMzf1qHlE11jNp
aot32BWbM3UlnYqZ5XqF2aKzmJGJypFSfuD+EteC5satuAE+osUHRMMAndIOWLvA
N5LN2XfjUrt7jw84Q3IKn8abIGBLl9V8+u2daynIfTSqo8gwq6eUcloeT9rxE3oI
WYpXxIJh1Bz6RAhyYfucr2m41B2vUOK7q7Q5y7nseZlYXKUpzWMShrr2jnkHGVsf
LbjA326HzDOQnJNFpwl/BPMqsoqhz91lxhUNzOwd8TbEDYS2GwYXp/QLjGVmenX2
WLfBOHmx3e03wdhCFGytev/bPWQipFWKhAS9ndJ/6gncziWO4Wytzht2AVCOLBiH
aPykRL4LJI1xazkvyVNhyme96fHKJwLXQIAVaodOEMOf8u01dlha49ARsvYEDeJP
9vhrkAhXaOufTdNajwb2KNsjG8mAnWbmLNX7+fzExQJfPGFS0oe4PSDkiewzSOa4
2wG8ExZF9medILMPE+jWNwsTXqPXHKUKd9OJd0WXJf3W/ibWuTZY71xXA98C679I
pPn0yvRMRT3UxUqM5ziEMz5wcficoG5cx2PnhEZC3Yndw/nTdo3Yi4s2Ze51knJL
TQ7OzoPiI1c5Fg06bxQmR7yMZLWTgj+DJHx5kw5zOeKkYFSHONMJpeZhO2OTj4wW
P4DKkhok7J5oON6int0gXMK8m9bccdrFvUTnsWqIGFGwj2yYUGP7qahlNeaRlGYR
zUVStEnBQcT9MKxoacpOkH8roPviTVhEN7eIYBUgmLvu9RYmnlOgzfdqUkozW8eI
0E7yeel/0LWx0ujayo7fU2g41sQv8xz+bG4ApSyL0mDeYsnTzrpaBFSgSjIpxv9y
1d/4mBU7AlPbRTY4oJ8aGS2Z+p3VjkgSUoGjbKwDIhuYfudVijCbJisYu5PAhGix
PBrlGMkKl82+10RWdqY9II+01soGghu+K4WaNLawgXuNJPpQSStazQk0keq1vAjX
gQTUf2mGTN3/k+p9GI5vvvu8mEItmJ39L38jhuCfYwP/K6LDAILIqPzgfTyBSjRc
E4A0niCsCJeHzUesaAmQTHQZVyJkH+uMgkOST2Gzou8g5FK1olBEM3Odk0RwpNdG
icp8/zYNtMVLJ3dQJH3GZh9zlyGo4iXOgQFwhjU1/xccMPT6FzN0Qe+XubZJXj4l
C/7CXemhK0Otzi67EMTLJeUwHGR+Z05MEAT3nKOWeNBRUCyJlETUeDblpk8BJPqi
N1Kf0X8OhJY2D/wKtDqlciDz4jmvfGgUTCnA5lw6R9nPuUYGQsBM/x3f+ApuC0mS
4tqUcZG5sj+dRKZwLrYyrVphlXsyeSYI08uigfTtfJUzq4Xwf86Fh0A353UBae+R
Jd5Fx5+ze+GweBGrkI6y4huvOegzznzwm5mYwUGFi9QarQYvJBbn/MmBf2X9SMeq
d8wTfGsnE3hnKAp4/feTYYVGcU2G/lFXNNwxnEz6/iVmcN7Pjo2vMO1qWNnTnMKr
/CDHDXIGOmnYb7DsTmAkes1HgpvUQSgR+bcbB0ia/mLO1xmEm4+F2V6ONFpBlhXO
MWIXlxrHYeJx3yOxzL9TX8hDRP8TBKxzR0CIkzjXDxILmLH3eaTXzlYhzRI7z4vl
G6zOQgjbzZifLMSCmtu70sa7y8A2pXYzzi8VU4FEBnCnvK9g6vTtANOf94fa2r9b
SwdyMaccD7HYAZJYi12jJuBA2y8Fhc3+VCYeEyzGkpN3PkpXKWm7dMjzuldX/Omc
FY3E5MbFmjNmgtFSOZbQxT1iYNkeAAINZaZM4zAnTJ3CjTToyas1mpoxhX4CZx3S
P295iK7w3WLoEELztY6SNtDbh/mI5sdKHSrm4lLyiDa/xNNErNlEg/n9117/57ua
U3WbD+75V7XM2rN3VBYJJim25L5f2e7AddKM+uF1M+WSnePUsxa+LT/3imMVwIwU
7VhgGIF+esqmBOoBMFqe1vNqV7/rtmyNc0xBuyWRfkDWf/EqUsulftdRF7qrpGFC
RZVHLoZeWydlhu/E8QsHGISbNUbe+Oaol6kAQZ4yiVAgb/vn0xwlhvWs/2GGsT+h
noDggckq8WPyhRRev1y6FWkfuzuTDVl9/hQ93S5eP4yYy42bqlINybntKYILAa7n
FftXsWf9bHF7TMTd+80De605IIStc/LAHEyRgZDV80e5Xs7/OzJX/8KsFiaHdmI2
WfNjPKA2LHNR2uZ+vtBE0KgyzK7JO2jqv7TscaVC9rMW4aNgP9xi4cOxH8DxlYUV
vCALHx+iYZLuVdGg3eMLyduEmYHiAuIQFQIFa5oeoE+ry3MwPx70fOXoSh7/513Q
YhtAC2iim3uoPR8EBPmmfK9gydsV2QVey+5rtm+EN450cNtn1sx10jIEGXlewPdI
l08VKv2ak+RqvMbt+MHT5GfQaT5FHo8sI0jHr5+8EVtFdoBUQ9bT5RKbbyiCKEpI
WsI6uel7bZl63vuDdA68VPjc4jZiY+z1Qn1js6/3XN6Yl4weAxlJE9Pr1KbBdpeA
1+J99QZPwEzfORfF4jQkKXDRXCtj73KgxWjYZplyGO0xn5GDeTn5tz/fBpjTMlBw
iYNR6uZ2HMZZdqXW6nm+3KWLG+PqlprUPPmlSgyPxxD2XiGIALJgCwZOxx6A6As2
0tIXn8oY02RIwHckHZrFElNWoXvMK/YUh1TNZx8+5x7dYk/WSjvkUimO40txUY3X
cR+SJspmcfbjZRXLyVMBurdXZ75F8+Oh/ISVxZH7V7uLvh+7yuBXwjpgdCBseR1p
jykoxOBt8dhZS13wf96QZd0YhEuCy7PXJdS4UwHa70wma5eHRIhIeSUnRGTdaePh
IvDllAthlyp9mEI0CRsNnQVpnMKXXYoSJ3oGlCpAu2JiGsg3Z+qBzlm2j9f0MDvq
Rwe/oQ50GXOffbz0+Qwqpz4hq9+SxI2AiyoNOZ0u3NbRwIq0rSIByMuNBpQDg71g
rB7J5K+JLhwP+nC4Bt6iHV3mDmhyIzRJFpbHKGXGLTL8fz5idk+1MWsl9/9RH3rZ
HGteBqndtyz479uTuDLYVhl8oKcNV1y92nM1OrUiixgPXwZYZgdFogx1ZFr9cNC6
8PHMopdRteK/keneA8p/Zw12EgonprTTP6ee0JThiwVU580MNmv+DMBt+m59WBCi
W5l+SMNyeUF+sLJAUqVvYOpOJ4HEPI+bd8hYrnsOlaRAzRtCbndURndhut5izot4
de4/TrfEXHpZGxjZ/J4IL/w7oGnesn0GNKX8vOcXYMSW4FwHkb3YfKpfDnRaVOEN
XUJOaZhep5cAAsPso5XzSW66pgv3zS9x81LowJtoGJG18K/rvcQ96DWiPQ5zlpdu
lANQnBXSDp251G1p2aASTstBq8Y8Mwdh5i9aCowheOPjw7eqB9qB1gJ8bEOMJmxH
4j6bM7EDb9+1H/dP5XuxOp9V3lU57n33qg2f90m9vZ9CtxX8PVzYU6ykYDKOmC1y
L/fErzaoWTqag5yi3ltCedltcya0fS0f7ReHJd3etJ8kf1gLkxvdKaLVbMv/UQE7
0QiDw2/vlcNU4TwtiWqKLtAKOFUBvBbvGmYThaiHpVIJCDk0SLS3qEbye8c8X/0d
xTbnZzcL0mzF8aPnO4fi3WLsyzP3KgxwLrcVEFjA+KGTBeAVg8m0HdEzU68j/5QP
lg8kuuXKfGGrk/ciJp9JxRPFfLn6buCyUjNdhZ1qgtzH7B47mHZ6soxEof8Doi6t
oWM6c6jlRmqiuZutproYAlZ8wyoFtTx43WLuOC6A6pir1b19OnJ+GO6cLg01tK1G
MtkVc8t+GOEVohfdp5YF1sZEfK0mUTRNcjL3hw2nIaGsTxFHVrM7ZJZjMQqBF+Wi
CBRJNWn5A7XomcuOOfJRHW7kC4Hr2XwNV8/g7qd6EcPDCusZh5xawbTItPDFk10D
Q7AjGkY6MH5juCb9qBrVk+eems2AYHyKoCap4DRja+KwT4xEZYCq4hnRtJHampDn
URP4CLa+nhUQg3KBvCq5fuZK2zZoAAdxwnTNcl2jWEN1pMp9UlxRjWXiuQGmSVua
yFgbhj4wBDSRxC4yW21M4dRqyUPxAJ59sGfxgIf8n/72c0tKZH5LF7JSG6tEa75c
ZZ600xCSjXfJzFAMVhxfasz6RlBT+XnvPumue3E/Hjzz6GpSoTPXM+/ib9nLtUVl
e8onB8EWiq98VMD9hNjsrJ9T/9/7Hvby0yuf/LJaBdVIkBiEYwNmIQGTBWXNUS/h
zUppAco0oDAl2U8y8CvIwOqBWbA8pxT36NwEqUgUT9vH2A/8NoD8mOVbpJitnR6g
qJkCmmCwZNSIxQ+Pzx8sLv3b46mzZOnBGUVbYI9U1bBDCvdrs1q5+41pSViO07GW
vqK+ZX1ozW0PSTnpfoUZy8/BRZQ8bWkYGzKnpuKaxWNSeMnhdmxiAx1pX+REq3Ci
ib7ykfLB5BtLfMWIWcLvdlE+3r/gg0nwb6TQ2zgnXj1gXQzDpswYdsYp7LU9uMsh
lMWDYPNpVL1WkJ+xrM4mhnS8zmt67x01jruWnDSXIV555O10MRGE1q2wosozrlfy
c+u9yD0kLfyTPsS42CqYqLNzWspIa9KQX1LNviRMS5lPrC8tPqiijSHZM+dxBui1
5AUbyIGs91D44CeyZCOwDdW9PAVMPBUlkw3G960NIdVwQBDIc2cUgkFT0+IlY16W
OCuuCqlIiuRdSEsEwg1QUBH3AEYJuhdChCszu7tqDKtZZT8pQx16ZBAYw59fNHSn
6sqVH1kTKk8zJ8DYFx/b5bpcpboUm5rjziIbvtDChMTD18dEh9u2bjHeBboFo0Kw
tdKsyAx/KK20V1fojUSp90PiYZ2aXNOQ25y7kNP+JR3m7+/bsvg6gxhCYlSm3/fd
5BdW7AURp2MuGDjWya5FUgGFBwskzT5MHNigPNQDUSJXZc17AZbPBgkYeBvaGLKR
BuFotXD/ywufk2Ru1RUS+rYmc27MPpwbiYwatnGGphoKCe4L+dtOYkIBMpYkqxQB
SXCXhYbdaPtk/7fmqOVXvkTgrkQ1y7sunwnEsKjKq235KKD1ChmBTfJEytv4U1Je
vRKrnWQmhCCco95VFLkfptPP7xopsQKpVrikT5qgY7V/8zvD9pMqkbXtAdecUl4O
73nyRJAVZbdtLMWgF6hQefdjpBrtCirRV29QcJr4zeXEBlAdFd9ldSi9Vs9YbhhJ
Xp6Obg+bLL26O6cx53VaDlDQSzruyrKsD+0e/ZWVHCRzzd6SU7Px1xPggG1ThrM4
78W0K9j52LiRGcbBSR/DTdyIFqvGB60mICW3LYHUUcR1PtoVrmkSlWWA6k081tuS
oKevHwccPassH7k2X9aJBzlqvJUahMejGrcugqxoa8b1GC427Cj8H21Kbl+6ATZF
bTULmYTfwT/BMniC6AoanS7hPJuRqCUp6pn1eZvWhMUZ7tiMQ8vQ8ek0AjrT06wx
ddKHzQMB98IMSLWHs1FPu8RU5VF0LBXlJZ7hf4qAhzJGC7CZpGmzyzef2LklQ/ia
/h+wI6BhEq7FhlVleixU+3lqMRS93V6cdWoTEKb3+BmYs0RGcKY1+tWaoQS0cv7O
0t86r7NEiKaFZGPos9FTY6m5oV1oBcmgcJL547FCRxOaj9Jhitk/SLi5v0AZEGnQ
2u6VTZ0l5QhfI31FRcdcD293NzSAgtkwWR+q3h0j8Tbj55Lxl4qYRqWem+dbCWw3
KnnOiIDzJ8vs+34sQijKrvL3HfPophdbqLv6quLOM/k9200xP0QI3z0NokeA8H0U
Kh3rVIjUsMCdxrM4U76QdxTBDIcVjmv0y/LPUq8dXP6q1BBPAunp+lMADe8hWnv9
mbzTkrBMte0h/+MHk5N9BD3el9JTa8Hrib1KdZ8Rb2O4f900vLPIKItF9KxDvDFA
I5cxMjcm7OrRPrp9twv7qN9GmXkckj0osQtxB5lAA1nmJzX3ibD7t1sD/p0SqDma
b2toPZHEAlf7Bn90WfGwdVnW0AHzdQjnNyfvmBwUpk3xDT0I2qx+ZCowdfTAQMJv
vjrbaoaV5NNn+OuHssmkU00nysXmKMi59eW23LF74bMX9p8F8Bjrv9i9A/o0u7IN
4bZpLN4CS5+vwwOTCbXQqv57HfMFHmDN+SAZSY6olGftazydtanvGgIg0gCUcKvK
nxciBPL2EB40Iyq5WGJg+HOxYG4n/3qEm30MeRn0wjePSr4CYnMopN9GlC6N++O9
rNrbHpBP3uuZs+9xybSujlTPMSM4C7teaHragvcyvd30/RdjRSh+cieiVOCBc3JB
kDAWI+jh+FETkFDx8DpIjX8ZmkmuyDgA9yG7uMobYWmnZkMiATsrVsVDLOhr+Wwt
7IJGUl00UTfuOp8KWfDb2kANeQKS6+oCel100woXnkFcEFF39k8UFT0QXTFmnlKl
DFDEfHwx2S1qJ6/ytF4A77nXBF2nE/LiUJ4zxaMysJKnVO6sCIjTR6ZjO/MNgUIZ
IHNiRyxKEmtKpi6SVIKtrSdh+dPmtnPRiZJMk0YIt+M6PFAOHuIRGElvOTGKGeIX
VXBhK0T/IQVGPD9/JonR5GH/vgKFmb4E6L1shXFQV56wHvz3+DaLSac4QVmbse7A
xhyloYj11++UpuxckbwfBtJoNGw+vITfBZLxycQXYJBLm6UjjZ92fV9BdXKKtdF3
15Ke0MiNP3A33URynqumVIJ7eCnAQbOM+14hJUxaMBI82cV7zyjhlPoV/GAv1cm3
5cQeGADkSCox/ackRxrneDGo4Z2HNASBuZa6vgWjAdJQrkJq4Xgk6gGbV5k4z7qH
/vVo9ZsPRY4FmUj2QCv0ctNcHPwaiWDO7dBVa7tRuMV8TBTrGPxmHR+rr06uBbbV
em78gYQhe6MnxDkfQYBTgXJMPhRvGrXz0ZddNYtJjfceR7Ho0RaHqExAruXsWo2L
62rbX+nrKKzE9OTbEoFs8kxB7mur0F+gCo328nHRbvdgIo/m2Mtu0dVvF0/joKRc
PTWPu6d9hO6Lt4AjtuV2dBj7NuhKjxcjdvfK4YyrClQlamXevxgKX9ouyhM41BXf
0cYAWgJSq+FutFKURM6XZP0ubTYHt3QeYwPbWhdx4qmDAigtI/RBoENxUE3kDBZ3
e5vTe2GKPkDNlZjnrHWGWB3OJyeIsNdaL3m5Ciq3us5gVJgn/bv175Ojxyxu3AjG
RIKGWPiz0el7lXtGMlh8+K4qllijqR35zTo+z/V98VsdGoCanFutswVWp7QdqA2H
MHMybiS1lQrKMsQ9YB9q9q+DQztsgPeeJ8DZuX/9xgI9OnHzYKhj2j61nYyaqidt
nW7WiMlf2yjOjSm2/kKtXmXPuyrtixsU0ZvFbMx2piER4Pm6dmiHGGrjEdcrfR/s
mILmfS2uYAKN93cl/7d86b7YhWUB6T37k7mwjZTKMzqZjY+d8MT1muDcEL0EEVOz
0kUN3NvvdsK/j7sPMx7xheSp85aon2JGjiLb/ybmnrsMMH9nT9ReAAhG+1+FS2xf
n62/o1XNeq1sI0VUElrakBHmsfhASDiiyWXmzjC3DdLb6vH+Wm9P7jwjpaOt71T8
yqgeyruInE7sWNwXSvegG5zHHLq57c6CN7v+Xing9fngfbOewqVqi11hiBTElWZ8
+YC8wM2ipN5Zt/OxMXSguRDTqf7PmbJePF3zQmYVs82Sgcwk6ljhjj08sHhBMktM
/OhVTPplBlFL/1cSYb0HDLpKtMyhiJ4CAe7FleJ9qsbfLmS6XXOW3mMHJloJ3qsh
cN/makhR85vWH2tX3OfZEoEH08Z2fwBNK6Hmx3l4vybzeY+tIVy6TBi/watyPltU
kaguGu8eSI9PeV8oqNJTsPS5bz43naEHpUvLmEbvvJ2GGwBydJUHntVcHwZcROI/
jlyofTL6b9G1cr0pC+U/Uo06m8M/2hoRhJQ/PPwOYrNBxHj7tU3lLdOZLiqP+paU
MXMt32tB0s7fJltggZBsTev5imYlhEsi/udl+BBNjK7KIo6fjY6K6gobTs07w47e
KQWTRTrO46SdNTOYw5mDsobLooGJc53XUSt1GIqVdchkakfBb2MQsR7SUP+Qb3Sv
0VXYOypRLJg4YCOxRibFs6FFBgMdg+SskbJWL8jztF0K8cZUt2wqlYFwCgz8qtMN
iYDUbOUivpqodDocgEHBmUKEcEjccJx/15cc2kFa/hh79FFpohyAUV/+Y9OByR3n
XrfYz0YNAOeCV3P0jPj58F1+RWchcKwMqy9nGhAxfqSuvINUU8px/Q68RD8FRkvM
V+s9wWGRoU+TcYeHAp8SI3316qr8ZniFyiSlGElv3YRP6C7OHlRznVvInmg13Vxy
cTMWIskFghsMWazMoEvnZwaiyItq7UAoRfL49Nqbjy4hac7NXoV4SLvPq8LqJc4X
KmSG+stowJCotowT4/UqIskddO4dsLqP3iOoeQdvaRyRXuABI/7m5/mltmZQcwvr
hiJjM9VUyk/h/U0y1WjM0wvHAGbMX9Rdw1uYRsJQUwu3we14TcEop+PoT/chMyae
9kT//mSXpnbhTwRMjwJYZpMX9s1qavSDzswCMxhEvhLzs2MjbHRKP72xBehiCZbC
pJ+Bn2B8N0/D89ZQF6+LUxDl5M1gvzSnnBFGp+x7uITpeyy7WCSGJEqlWRw50o2P
pA2OwKmO2LJPIvobiDIzUe6TA4azxZjuIFBk2bBCHU2c61gjWUj6pTch+nqxjk6T
csOeFIJO5sHrgXhH/NgU9kRajT+ZFuLp1b8C7uY2Gc2h+ZttwmgLcv1M+M9o807y
uB78UIOEnEpQhuoLthhKhMC6WZXNvsiJOUvD6JYgc2jA1DTFdH1yzKH8WvcjqBj/
HN0wujw2vh2WUM5hxPRpwzyVtV/RMiM6dS/OowaccExQfzczbazNjDLdOCqSIa2/
R0UNFxIJhJmrk2Vxsh0e/s9u0d+/Nj418eh9CFH+5ifTwvv14EHGuf1vt0Q23GtV
VMpU4LGZK5CWqoyidvFcBy8E9+Pg0bpqZYWwqa2OPln4Qll2R1fE5t6USu5IzGjO
ARqF16JgVpfxmO+ZQpyhg0tohS6qkoCMh0I4use5fWObzzhzhn8siDQyXrY3hqOq
OxcbN9N7Ih/7/H5jpcb8NHDAKx/uImnFjjNDiEN7U2u7ZQLZS6x37FtT17L5XcDv
wuelMJLcJwWJ9i/xLYGUoT8q02EoaefPXDsZe4FDdoSrZg95vj0FdS/BcJpV7iI/
vIKapu8zXnN0Xm37d/laWOiBleTXmM/k6jUm/ky1RUyC16mzJqkHYUPv/DySDVGJ
p5+vGeul6NhVqdcoF47Loq2vOUlwNG5Dnlst0Hqlg/ffMx6QrOGksTb3s1ZX6y6O
yRki3llFH01rb5CmanpqbPM9TevlQcxvxcGihJlu+r6sLj6XbLaRY34kVxOliIPB
H0M+YIndiO4JZqkfKPG6L0DBqxSD1QvUca+afuNB2ZSkG/zmbzTOlqcEdHj2v7zk
4NDskKWAjZN3E34nDvvo5VW6razWpYIV7HQtqC/zrxe5ARe/xb902ltw7BKKxTU4
LE9956hjY3PJhE73rT+crlBMfSrNf3O4h3k31m1pPIkzG0/pZqhHjb/Q3w1IUmFj
IO8YH86+7LupIosCTkiFJn7TFttehHz5RmSf/B311ZhhH5u74g0GpEKrzUk8Si96
UOQ/1BRGEug6VlsihPkx7JGPOne+fh6zv3HPqSqiTfDrRSVhKDyO/3JKmpq6xxq2
Km/zSfor4FeVA0eTSIq9hujA5ftQwf5uHo3qgiF61+vsIPnkSmj2yKe+r1keWIyx
83btS7OD3AlXBa0c/TGlh9C3Pa4paN8ciqEU6VaJZrJt+pxd6mEvdeEgx7D0zPLF
7pb/brnAykhna1A8T24zLIWvWPv6onnw1JJUo89wWoroKyJhXhQBJRsL2uGXw+tZ
/LIenX4XDxveL7A5D7Y5aQZ2zLPHuL1DNBEVevblF77dD5Y6BxqeIQRxFasHt9oj
TtYWATVaxFvElgN+DUpVjLLe3IKXG03FcxV8CmiLkeL/ql/dlyVm4y+/7gNY/6gg
U77r9W6GlEfoyMFAFXMv+NZ8rX9ClU+DTyL06/RH1qNSjwvxdbSMBU66lSjqggzG
FKXLCmIBl2bCm7koZahlJ2ls97rj+sGWkNdW5yPUCJJCcAI5xXa+Qt1VcaPZtpdB
go2FqTZlBaaOhTVCj0+nBpCJIlB+JN8nV7LwMe1IpRs6xe50IVHzMO4BfGFQhFFA
8aiu22Hn1UvnPcWXTB+79uQr0ENLEibAMjZc5sKDpRwuX0WzA1MW0sX1xnMSaDBb
rXLPSwB3fs7LwjJ4K76IhoAP+rsH4mkNVR4L+24p4bx9EdA4yKoTcYakSxUyiVmv
8tNgPuWVukU1Jw9n4H5apiZwg4gFVcS/nFua4Skpc3xN7PGyNfbb3uWcKAPOyW6U
JBEaKmxxZY3Jq+ZsRQ1uMikNIGSiPyR5NdKbRdOYvNg1luNiMEPhhiooQtqGvlxn
BvD/pQDJBHfAfpU5/H8lYBl+xFLYYr2d9FfbJhJu+m/0wLvDilCJZxDyUvRICyjZ
s/i9b3CQWRvzZ9L3o1BUfexfnIo1EpLpjDUmvbxr+QChqx66fMy3JgYVdBEtsI39
ozOL8H0iV4F1FJkEjrnKUIgleaCS2n/PrRm4D4Qp+Rj5gqOEsVQ/DmNKBDjheqQZ
e8wL54uhydSVqDP+XMI5U+5guhWUntGpdJ8pF1PLigcMs+eHEnrOYXAL8hmpizxW
AfXBhipz5/G1C9AZERz8Anb0P2v+wj9XGP1RYKr+yFrnTKvIvjhJsGn5Q530xOnt
gA8gVooCW2l7qmLXFsRn3IkYy65VXc29EieyV2A0/3w4fCX/GOFGTGfp/V75e8mB
Jxsq2ji/qH1cgQLkJG+sdjEFtPf74urjKHASMYj8AfW07vKf5BYn2QHVlGFRGCMT
2B1XCW+ZbRQ7D+tz4TOeSGoDOFCFsKKmMFqDUdlm4WUTZi6x5HF4jOQmSwtRaMHQ
qqFSYcvuZfZCG3kOHwdeFgCypsGk8afFkHFqJBAy7irtw5vpj3tStyD2+yNv37T4
LG7/FY8SKxgUVjnBvCMFXmsK6tPYzOJmfaKn0F/iNECB1wYuKTICAyEd2oyC4sk0
jMFIXst6QtrIRj+00MMPzySYuU5N0jOe3ou9uI3s8E4299BAPdQwW/jcwsk/FzFE
kSXaSBFXUyyy7OWBU5cmfsvICeYJPl2uD81uiJCSr//NiS7BoOW5XJttMbrOsNzn
v5WuTaB/vEHZSWcEzKAQysyluZ277sr4o0kWYdSqnBpjVV8rl2WDVInnPb8Hu53F
TiDtj+lQBpmSsEQIuTUaiqCbdCbj+Zfar7jBeRj149Enaa3JfBcvDGQ6zW6vxqIv
t5+uYusV0fE8Xbt7Yge8aK2ieWhOYyKn7TOIqM3FRDw8fcOqCrKe1wOEfEweQUgP
uWI3mVNxXt5bvnCgpepm014ahR+Nm2Ta2agiziZkB/Dtt84EbzsWJh/hvYayoRTn
5xHMm7rCgEGXd5bL1TGMNMLPVTVCHtXLXCmB5NBE1rHG8bU4NiZaQQwfD5sMIn1q
okZWwdIn4nXt9IeTQRvLKi6X+guucFDhjmYk16jdAtNanKTTXUxmZaxaxBoUi5at
0wjSgobfPedLV3mNzJ+ent5/LObf/C4jrOJ9yP9vJQ/AzAD2kND22JkMf/KhVqTc
ahch2MB75MwxKdMoInQdn20N7EIkDF8aA6jg2PNuRK7KJTBZcvSKKjUUhXbh0knA
lOMMF5lqwdnwldQ1Zup4uuPw2VNRrLrcwG3jJFRRIFWm9F9EDGSSiPCTLwhPiRZY
ZHqWqhlInrxCl7xye1ZaJfcCpo+RKQn//Y0LNrUZg5aHH4Et0TRjjqkpitlXTDtQ
gUkeC3Dw6oJq07xnJPk4MEHKavA63SthF21p666Ln2WDwnNtRj2sO5cHoLT92udq
sCrVb1qWxmcxuj/Tq+3bQwNRDGZ7kYlHiYJxPImpN9S8uC7YRhSLzrVms2PjH7mo
4eL4UqcNw4BQmh4hWIlRRs1uwaCPRmBUnl//9W7MqWTQgvhXpCJZE+O/uH+iyATd
EZS6iQZLNK3p1fhQVNeIRxQEVVyGAJUcSF58+g4vC/SYoAuzGSL+pjGguLFKwI0a
+5D/R3pfBk001kSMdF0pEhLFS6WYmAA+TdZUlR0swqkrPY9BuqwV/q9iZqlQlPLK
g1kZfoz/TqSeXjCXdQoxplId9FfKIXqjgPJfzLTvldJR1gpixXydP/quWCDocxIB
tzeow6CriW5INNzsM6B8Q2s6OxldxwRKxvtDcuVt+MgwMuj4JavuOl7wgrMjxMMw
Nj18Bk8uCMcfG1dfP+5x7cPS0xl6fzj3ALTdrSfVsK/iWtH5cJNw2toUEzuwDa5T
2lzcAqF1hhP+lqz/9eIP351z6CkgsFr3ENFMShuOePU+OHXyaaW7UjtS/KEk1Xgf
M7J8afnxMbuOxMqJnKD1FUnrInC/J0UdriyE+WuQiOa10i1dt3LsaA+1Z6s/1289
Ru2bp0Kt4zJ2jeHDC1cpt1UCi7UnMGiFGDKLJtWRCiH3b8Jj2toCBhUBTzlwvmzV
9PR5CwXGP7uuhUYZSAdyDKjIgs+1xoXYnJKrLjed+gCZKMaDpZBaOvvau3jdQgNj
DBC4c2KlKkH06cVBskfi2RsWb4gpA2LeM2peO9GMaDxd4f9mYYsZw1JecaHdw28s
AWNw/+o8kNcBPtLJOYAxVnEhNrKvjPJRMpiqKPF3ZHPvc+7aiu6WYjJiA6DzVdOo
w22005wHteYqC09H0yltMQeTWYyY9wbXyCd7xEBG1qvaaEL8XhT9wtVt56s2UY5m
REwSkZHqYEFBp+EoamwEBHkDmf5FZvwcjrbWN3mEKsqXMWQageNVF0O+1jUG6hq5
yGGN5ZoRuK7AgU/vCDskagQ30B5MyjTC1RXUlhJeO6BQxhZzIgNbgSis47Vc7nt4
wKsLeQePz+CWA/3XKUfCyopGMGD5VoXjjUNPFEVInVyb6YMN7srHGwNhgneGaqtl
HaOSuCXGcmm3tGKOwTh8uvTvaLzRDOc1kxDMep6ZICiMPjWmz/Y3lVTt8zG6+W7R
BMX338Ucmcf0ySwtlE1sxYlJQNFUIt4LMnyDrf5q5JYkf71ENF8eOsti8Vb3qDWI
hi2XiKkkMyDqZbVtnnQ9BJurytHDpsz06MlNEliUvscJMLfOWTVU2wtzNJ6/kfoF
ey301USA1x5twsotXNLiLef9FEoCcLj8moRt1zQL2+bIfHkTTowGiA5KGa1jNJZv
2tgDZp52mvVuUOHzLJSVbn3+307VulLP1uWN8uv01RmJ+/EqmX83QRza20gnwqO5
XbZk6wNELecrDDWOCRtFYUBfd43skiacqTg1uKpyHC1+PTFLYHD2hyRIEqLGHSbl
+2HXnY+w9Jh6prWuRSgnyu1CCU891Ohe6Mj4HaZHJTqKjdixWHx4BYc6hkdqKjCz
KwR1T8/7pUYQK1fGVynWJ0buaC6iVsi0+P3Hd/vl/b5TvyhEDcd8jiXa4Dl8jC89
VlY38UwV9ycIyC21IHhJeyclDpyxDJw3GJhR3x868RIwGmjD2lT/2dX1OBLmrSo9
DtGcRQdk5kVGfyXDRjNo0hjjYx2IDKDDA1VrOgMt1VN3KpDGLDJ7sEKQBIxBa6CD
Jq3a5hrcrjIBNU6ofYR4AfIHFdzoznxoCzr6IzKFNo5KGf09nUQIM8OUL2F8crKp
P9NYBSNaFgi6ZGHw8cl6NRHKwBCTznHfTBcuzCXxaa85dZHqkQi69aHHSbdN30d8
nqOr+hjGrl4Oh8KHGpHyzo9sa5OqGiaIxLmhK2sPCvOgijMR5Jo/Iw/vPeTJMZnz
XhYM9rtzqox5NfiWh7xYJw2C3S3bxh1tI6ormWY4CDGuuGcGjpYSyfY/k5XmCLsQ
tyRx9mGZ+4FXwQ3TkD1vx6w0Y38TqZA/8GPBVHak0/N6xCjWWqUIiMntbaQ4mDor
yexGNfaGGY3daX5uVstHIcCrbCotd9fTkKsKFn4azWCQO/OS6GphXEm6oKP3fPkV
U6LnVxqXDzWiU+ONrmRP6fP521Qe1c3R9dqx/pmCOeEfysnpMZO8o0fmFNiKaRVc
n0yuKsJCoBfAcWPTeLxsvAu5/srRbR66kdsaVU0wbXX6zclUDcBSZ/FQzQMTHgjw
KhJEnYXX3w18CYaigIp1i3jVsgP8LAF333WyS1fsXEhdGBEw9WqVyMT5TtFEu4MZ
W6QvUd3NuTv+w2vBLhjxilz+I2sGZQZOD7Yr1yZ/MBikA9Bz1ag9AqbbC36/Sjrx
CPRkqnDLDHdjqoqi71CkTDFXn3ggq/dnNEkIzXw5G39RGeYdmcbG6CkWnljyr6UM
BF2TwhId8j69bzC38Fx/TpdmzWDOtOkfKpfu9YwVkV0msHUSM6F+GWWWIVZsQGce
uDlqX8uprdPEvgHN16e4/1QqE/zxgPc+tX9j5FGOkOOOO/FNAkDSYBniv2VNZs26
mQPFR90hcCndVhQLMwRgCLW2lILPORDeIuzqF8oucBGWGkD3qXp0wKUWeZeVRphR
iwVpFEypW4G9XbJ+WKulcksR8R+A3rNjd6JDtS3iq6OrSYtWQESLw9zqll4sXG+Y
2qZgCYoLoOzyUPG+bVUTR+X7xAPNDZ3mMhaqn8+EXhOqZKSZ9n3Q5dLhO3UtXLvW
rgTRpwdZi6u9x1wc70bZZuVhC899j+H3CmZVMVfYfQH0XReiQjbYDhCzorfMlDZf
xBxN2dlBnyXHY4bQhpmYT78BEZcrFe/tNPTYR4qLuQkY/i4bHeQxBzWbqa1ygabb
17Il4fWN8F9+LqfhlrIppnEEhyJol/hURRDr48NN38QEgP1XnnUIWoT7dTfBVnOw
RalrVJVyzPLjHTSEsBlUbELJ7dNZFN+nEBa/8z26sQc7bMn4KowwAswjlglMXuMq
ne4JzccyDw7HYY5tToytMDPeXCcOxwlJhqFMV7KJxgQaYbI5/8uWFMqONKmfqkzV
Cm15SATgdCyd9KO/gHb/eoYkdrEHcc/T2RAers3KJ5EOM4ohYF5KQ3cWBncPGm3m
/vCFrMx4MKnwRgD/6BuV1xSwupKOAC4fGVeVSYB0InAfcoi7IT98PHUYfWNxL9h/
yI5/jIppt+mpuetpm9AmBpHgAAnqZFy8C8O/3FDSnc4rl9Vm52Y9qcN3X8rDxF2W
Ju+gr3Kti8Vg27iCZvuLBpy7rfoUFUDQjluAkv1J7mqB8oVVCJXWMuX4fvwuKdsJ
y98yxOVvFwhOHCKj2beP7eicLrXBkx8AaRdRCw5VVD5mhDaI69ZPB5MBf4jP3vjS
z8a8VMzOeXLvYLyDthMITHlvOW5VirKvw004RHQ0rw04zQL7oUi/mvCtUJNkDx4c
dsJyQrijEcbATtmBwATQ7m5DwGffy4qQoyxJvrGevJ6qZ9yLWnk6uDhCDnriDyIg
jUF+xw1QfEdJ1i4U6mDXLVbGuCcO7io0E/Jl+LnM42o6qbvu3gdj/sIAO/G0GjvS
mNDQqiK0GOu8EpMXKfcY67hnkt8i6UDiseVs1e9AyISDLaoLAyr10zEZWeXQGtBo
VooM0HbqnyPBweWIhu7CUILebPDzjHT7S8zKfOplptzbh/K881PT8goETPqXYCQD
upesofQU/ScYqJBgwQDCZuj0USQyaO4ABIAQOL2IKlE2rPaE3M35om91w0ORH4bG
OMfirCHbNQJqfHQDUq1ozDK5NCX7FgHe0sib2KqmD2Rx/QLgRD4dzT2wYd1Op9w2
P90aRmznMwMew+aGpolMIYpZNzzYN2CGKGsVc2NbkDnHkDFK0+pcZCd4aF9OVlA6
jIgGCgl/qF2tAkAMVbdvyYvNuTIpaQSpI1KuL8P8r5MhOQYpMGKNnhwCyKuZcVgm
VVTm3Wv1zUhRQSRU60Y4VvtAiBVqGaV9smBVMahL31hP3mRJJYavIzYr/LD7BQup
W3259ERQQEEg+i/KfZ22JCabTmwx2qeG85BuIMtprCOKvz8WNeS4w3MdwEL9+xus
O7SwnINwi4y8Sg8YyqA0YSJDg/gj63nQAISJLElMPoeqmDJGFxvdx+p+KryeR0iy
RhstKxI30XZiBcmLSNrk43L1fqGXfag3WMon9iAqaUQ2vX2frjdgyreQvSz4ULhb
WZ39OpnJJZInbGJRqUVti5JudJvm7lR2xMdwEakUb3BhLGSgDOYfAKRARp84kmWo
SUVmRQPmgd67/7Rqsz61gY6v7efL7uIIhuDMq6g53mj93fmUPhzxtd/kcmehznW9
zMfJe9lV2P91cKGKOvQYIijU/sYJbqAMJvjZktJCltzB3wlXUx9g7Dwff3hx+8p1
5N7/uGqCYYJ4lCGeVRnLPosRQaJOOMLoCshx/Blmj3bKR23bZuXBD82rzGEzO5YJ
+A6ToFIZcrrQ0jrew8sUMUIl167W6GWnNpTKjdAdw7WjabGdeZayXDblTCgx2KJu
bq3nx110hCiCqf80zkxQVqk7aL7e3RrogbFhtVqwMOsF7auW5KWyZjtZ8OpQh/1q
+YoWJBa/gRCa+KD1pWR9PxydcwWz5MVovUb1+P4MRLaQQMvavZemzqALdVy+9oyY
9rBb5y8HWs7r6Y89PI1333BTaF7kuQNGY4vTB3cO7f3vlrBQoe5/Kek2nnzfc3oz
6IVZAFPF+nr3n9noGRulEBzH1vgw4Tvb241hYaYxG58BcGgA72hGbOun284VvIa+
k99PP9tKHTTxB5mQlSMf17stb9lmTT6qsWpjj3/ZadkEtyWkBoHr9HtlGG2bEXb1
p2BBv7NlCVCXtOZOlk3eW3TFxQwdZOoZKl3MLSzUQrTOgGHkGIexoU20IWiUuF2X
Gqtj+xuVhETMVGWstDxC3Ys4dP0iZaUc+OySlB5+FRDk9Nc2BTWrURFolxmZUPUW
t2EDQt1H6ysMh+DhCElCqbL7/yHTOiDy+IxCuUnj5npESb9ug/HR+rbYDlNkX7a+
pODX5uqLJQx+6I2GWzl5QLoKp+iodHeID23iy8ZpxwG+yP14lT3S6OkEHmIS+W9Q
Q0FxsUbKwuID+MlZzvLMNz/K42IERr100eaMHaNMKPbGpsTzDvaKYyy+hQ0QM1Wo
aQHKDla8mV5rd20ghPntaf/fQBLvM8amK1gvQbcOq0s6zqqoco0EcgLWcwr0fsZx
aeu6QHqWiHjiXCgTg8sM9tiIcKG65pfLV1QoamgIPXb8CIgI5J92cJ+iJvwnv7UQ
bGe9BozMBDLAJAVqC+Jn7XRZCcjyHOdu2JK1ZUuwTUhyDqGwPDLVZYA5dqklHib8
td5TxWllec4SDuoOwJDIDLuZsYEbhS2y3gd5FYoSySGnpJorGO4K3RCWgaU9t5VA
vY4keAsB/0SYAi3LkwnyNat1NAguGkCTfkCjXu2fa0n6WtFysznHNOKS7RC7zVzb
JKWYnSyDkCpG2zCLz64JTkcWj7na+JRbWLIzeEqlykBME2iZHmX9Up714Y4TLoEX
Eflxen8eA/eri4T/fFRXsv++fb2ZOij1pvNYgZVi/lUVPCFges2r7HNFhLIaUOeU
wSpINwGZsd4J401hm0SNvrbcCyzMXVgY6GaFnkpp6zLit+Ru7MK50GCCa1tmvgVg
hxNYv9rdtjOVNXu9LTS5oO6cCpTMX3bUeESaWOISwhgMaVJpCKyct8qPzpYIbS9S
znLeMCHnkfgsG/qxle4i7hrkGozdLYKN+U8Ang+RgA/79Juh9trYEHmeJSQsKGUA
XGOPMgFkWXDbNLvrNzgwXTZIYnTo9QPX3pQOoZiPy9/+fJ5pOQm8J3TB4GzjwpNw
BVDwyjTHIOC1Y/4XY7+CZc3T7ruzARdf9UnMFEyU2ZIyajfPFlEGUFL5e63jmyWE
GcNwdXXSYp6+l0bHXsv8MBT65Rc0mbiDQ2S/Aa0oqJGLf+juN5BHAdWXKvaKCYsZ
EdbnWMVcmoT+s/MuKYFzI4OHXLZhGyqG5J0Sm/NyzWoWevNyyHlHk/Sdcuvfchkq
FmRywjYZaHk7R5NplWB4GMX3ZklmGy+5ytLCb+Eq24fOwv23l3bgAacqsc28C09/
FvWgqHV3s6PXsUBPxRzyxd9qNdZskgg1UvyLs/u2FAWI5lJvkDKz7/GVvWtMXJFh
KNpl9FU9/fswBDvdaU/y9J71smckKQJ7qg4dtsXuDwYRaWpS7aytDp4Zs4Tnxif7
yS3xF8uCTtgVzm1RL1ivLiUXNrCuAirlkBk/L9cBdsUBpNiO0IGZS7vbhWZYjy75
AowrEBshqUGZ6+N9IhbqltfTkxx3QD90dxYHUXN9LHcCiONjj+/iOvn3T+kwJ/Df
hyWgA19VgGJ5kDU8WydbeIzFZs5tAdD/xDKVXuPlVb7YtiiUx+hhxaaO0VM1Fbsn
O4hklpr5e44QHwVK/hTyJ33LI5WpckMm4XmuDEoQHAx7+/VXCrboTJy42sxthXTD
RrNBS0t7vnKtFBO2PJN4Kwb2k/jEq5vvzGkuY2UOqeLrNpxPNG4nlQ9z62K8aBZO
duhDf4pDqCaU3N2O37sdYbSOUsc1htgB3L/Sqk1irbsJ9tQDZs0Fu00kfxcFoMGc
mFZJoh9EOnE2qCkKYzN0L7kYQC66dyjr8+3h00xMi/5rAVd4WEPIlGL1MHtH+vDk
2csqeFzdmLRRZ5t//78Qi68XSbYl/rwEd5Keqj4N3AhAmLJI2g94asto9WRPD1zR
943vG0wUvMPWITK1jsLYmaAwBw0T833q0sNX5QZ9X9r1kM1dQxiLarheHrrZd8XW
71BaXTAh20qXveP54h5U/sdDXg696dGvZjHNtqfVRnWbGnXjiQO+xud4OD1e8Q6y
wKSRqN/I6yioiEt2ZAffwFQa4SN4yJUWLHFAonhTuGuc52Wbqm5eqiHIiU0535Dy
hphEiVP0kEGAMeNeOuVusRgFLm0EupSehtEWsZX1okgFGCOzZL/nymv2ML7ihebj
V/rhjXkVhmpoAIdzON0ulP7gvwCNvyrTVMHIwA5P8q11Bx5FSK+usDh8l3w2KZYL
aUzTVe9U7/9xXN9DumYMxZXIyzWTRxXYmYVkfV0hPMVDeObr6tYGuyJN+55v04lc
qkWKUvO4po7L87CnfTpstX7vES36S8dyTsO8YysS+YgNWkZS9lyM52Ceqc/BK1Hr
OaeRtooU7LwWGdS2V8E3rM25L8Cs3IbCDs/GKrH8ZqDvFhVkydRW1VrOH61lOpf7
mP0KfSjVhf4RBky9W2Xhjka6cJXC52OwGLaVncHejI7733XSDZVyOw8JCQEGnHZr
2ejZITA+LSqKimB9Q/cEGZwrUZ4KQbB8v3WwwvPKxT54z02gTl+2nUd7qZPCWumD
6Mw1y6/Yvk7WRlkeU/80fZeDAYmFvS3QN+XEmdodVfdvFdQr3BYxFGGeUfIOKViv
44AI3JIHoMuY/BuhvEbmBWVl+KdsHypDuAc/Zf2isg0iFOOsazHW6eqAGUjoSbZG
74fNNFSBmfrTDKiyIciSdx3f+IF3ARK+u29J5K/yveP4KDCK2fUcaA/LhLGJoLUy
zSb7VAwm5T/RGCxtu6S5OX2QOKM8IjZccS4IsknmhiOwvoNF7Qdd/UJ8Ap2bb5DE
oeBCm+eYZLuQF411IJkAmCuL7C3ZdtL+xv7X2P2NCiysFyAYDAuuLk9yglaEzAwE
O92KZMrKiQzSkLAllyr1mjlkRwiTWfliKbRTjM2UofpSFaM+9JBLbeCkBQYVDAwJ
mrrUse3l1eepU+XLd1QlxVeeD3VQf+OWbOI0ujbFrV5/WwbLueMVh5hca6hguhnJ
FTjhUdI7q26ZmsHRCHM2Ud/Ek/weQe0jYgMaVICuSVz/dPyUfumgCFkgmG+3v8uV
AO77d0Jtm0D6xJnEEX9Jh/ZYv3SV4M9irmLCr4PKzmj0NfGg+xNSf6XIB3Ri7I17
SxlaFaR0rtnNdRpzzwmcGitfq9SAFsM1VKE1cj0GXBmbqmnHmTpMDi7VsDIWeG05
xyF7XNATxcUrr26vt6sYRuqEQZeHxmEdlWTsbl5/f7Sut0Ns2xQAddTd7WzWcFMq
oOXj3BLF4D3D2fgpf2JUk2xYfFv09rGZh/blRCp58FZA74T9QM9LVTK7oHxIFfyj
utAwXHJpur/zttVLvwP4T+y4k946DaayKfljZJbYIthp2oYPpwoKUSSXNJacV0P1
Rl4uSu37NPCCmqVgaojjI7nlt/zGVYFHrygeoX+mDLBN0MowRWvn5IzJdBXbmrK8
hTX0Kv8fMnAkujev1LxlJxI5zdE1mKq6EAlLvKbaTtn5SrDUhS2lyNyyRYqRCTT7
eF7fOOcHZjv0J9nP2RCJxmdVR6go26jeh2OOP3JEG9FBmEIlmVWk9EwVOe2dgCYi
hQvJ0BdbJNjWaBpLet05lccv4HlqrndCCGIybgtHdKmcl954/CuY3ItmH1UAMDwZ
ZB//gCtV1zPVeTrKIlHbuUPp1eF6M8keN0NeDn6GRfMbO1rZYES4Qm2MTy2gA3v6
qxcKW7blqh4J4nEyFW63pV2V33nGhvGrh4Q5zQJAfe/BAris1H4LUJssKrkSod0V
zl9cDgvJPfb/JDdngJ2L7XTKElBC/gwmgs7zIo2SbfS4zNVBGEXq6iuOdyEajiBu
qQp78VtSHZKF1qs7pRdws1BgQnYRWR+6Yrh/gfYyjFjleliiz7rjAnzL1TORR3Zz
I9sLcdijA2jVOW/6Tt/9rfn6pFDViMqz/RW+1ZUMsBJFAyFRM7dNKDhDUp7DYJwI
YDZgdsobqtXo5/uRkiiHJKtF6kZEMrHD17ob9+E3lkp7LnyY43xcj9zrfFX7l4Kk
CJlRFPVU4yE3zLkM5OrHe6zdKbwQWQyIrh7STGhM8qjHXt6AVdiiM1zU2mQlqxc2
maU88wZ0kyneENPkS7vJisxdPos6jT2TJDPn893UPVnFnq9Wfg6w2ffabBD+Z75H
vvKoFFcafH8Wniq1Y6nhFT/AkEJj+N1TPKgopSNjkts3s239Z6BGBS/CDmRCPfoW
7Spzj8NOrtm/sKi0oxXi6gedqLm8O5RVE1k12YXbCOR5qn/zTb5Wz4xaBw+/sMQ9
2yBlpyMRi83RJYA+7NLkFzLP0GnaHcP309jrOc7n//0qNiFdnPT/uVzJjAVhzsnr
r64Oao7IdW1ytF8bQK8YlIAU5MKJn4i+/c6v2m3OBCNt0xweUJiCdUOhhfj/w61c
+fotE0quC7zQWscR176D/S4oXQs3rXziFzwV0zMDKFHL3nrvj9ovNfkPCU/2FnN2
Gf/7MXAF9kQqw7CZ7xkZQAS3NV+YQDOVkj1zgvBjUywaS1j/+QiG3o8AaqYWN1f1
GgfJrUhPcon6x9+T+c1SnYzfMlqQV0rKkyopvIYFPOnW3kkM8SLqATQKG041lZYq
MUuUDe3ntlo5LPtMW7vnAIsr7xPogkSNOTdshoCibGkWtiaVyQbzT829pNqJKn5U
PSLfjpTmAvrjLshM7ObFM4akb2CFDSj33o9pi33QgVA0i+Jk7IvX9pCK6LdinCil
V3pcUyNsvTNqWLIR5M3/hKzPatDD62iBkrOKakcWOnxYpA3HBs7X+j2Nbq1Jc3Mj
S8CoNq1zxvYNvXOjHq530Ucztq7PwUnBzA1n520xVodOW/b02PqB9BmtHHqG/31R
dK5IQ6GF/ppjc95nd7IY+p1LKW7y/Mkaaaddj09UAVjiw4NlTqO/2CK1DvVML2K+
Ch/EB1vNvPKgf66S3UNUsFUqMs8KAcHwgLAbj+MH2oU9rHVez4fjlFs+30Kn5fkI
1xT4ieBf64IRg+s7XCGJALeF53I16kxQWVKoqVDLevDS2SYjtofGeWIMFt9Tx3t1
LNCRax/0CUs+bkISIsMkQnTGhyApnNri6FP31oY7Qm0KfzVzVIO11Kj3Rz4u0KDT
VmH3vQ/biP+CMujMs8GZmpKy0vkr7zU5zUmsCbTG0eqIud7SAYrVTiBc/5gN1no0
tty1kfOd2sRnt17lyN03ieep+7Kv+FG4MdMgso5/YbO5jEaCnyXWSCWLowUtDMcn
t1slSPLfQ3AGEvTpOjosHjkZ7vYH6x5XogGVc9w0Gv1+ACMt0yUOLDyqCR3smf6z
q0hitKmwf/92s14p8VglHbm99i477YeoVN/uPv4UE+SNY0xP5ellM2GjZ4kJGQNp
dJ0PKW87U7wHBHxWEEKXRzvfpXKGIrriM4/wg7nCJFTSGp7+wy1KVFfBAyVLlwLk
udofqQaEwy66r3r+9JLix2U4hrmm2oT9uwGDFCGO0TiXdm/eK1iyHrC8oHj9XkdC
6xW90EsMdgF3Ozu+bVLv1xnWXRYy3XX65Zh2KmL1M+AQ7kPCTVrLQzePl8Lqvrfr
mpbytHNcWgs6r2R5UImLnG4y+CrE0pGwplxMhuplRNRhzT4U/beD5EUIgtSF40/Z
qetSzKSP5fLuwnOev99nHJZcHV94GHGahJSdveYUYCDI4HYAYTqfMBp5Qf2sOW0F
EofkFSX3M11OIXWrkmkBydKIcM/CxJ4CS0rMUC+DzzTOfATDiWV/gOuip31VvIQi
tYu64bnuCPMwc+3BpIRvhP4yoX/0Rjh3eZowadvQVHAz5wx6LvKL0gt48u6lwh3n
PFIfLUBAxnuw0fzboqwvU7k8wsFzmZmx3BVXxazQlOeatgFCjK/9uAtqtng5ReMa
uryw3E1cw/mXxQReYIwZG7gN1P/rTXabqmrsUD279uab5zWvukJUGER1GOaUxxQR
PhEi/U8s5diOY1RLYuTOvNPtlq4BsKSl9fZEIDz9OZqimpy+WzgvyEl4pcUXXC0V
hBQvvNaPG2Rdnzr/7ZbWkL1owu/c1GwSqB7bM01XkAIaD9emeuX2NwMtZ+qquPFl
RJ+AdGE4yfJ0e1RwXsZUcuAmj68IiORj4jJoaiClDDPVFhQT4Ax98X6qDvNsnV1p
Dau0lJPqHoL3n+mWSEWPNCQBTgh5BwddrTpRAc7Gj2d8gqjvUF25NYssZw9LJ4na
UIHeSy7IvOmYSwfH9nQ1E0blBEE0Z2iMZLUwsL1I4/7e00SpYDlBzCyK0Z42QvpK
CL4BLDpuTTWbdfwmYJclDvmlNzbioTi8ZAelgoxHqO0WWaFiGJ9EK2NKIBzzzG9D
4FjnDZdL1/Z5TIskw2ZxnE5UV0Vz7hi4EjWyrKo8PXbGIZdGSiiF4w7EWVkbvYrj
5Bd5O9oExV6yHwkpIPAWE/z8CsO3itbv8GDdBXRU7/cieSXQ/vXTEppbZCMn+oj2
uF0iPVJh65ugWk68aZLdqTK4yLrLuIEeAjfPOjGpn1B1sCtCNw+XsMtIc2QGCwvH
CivEqn/XeL2PftsmGPHPY35MbnP5kVJgRUmnnf/YUmYRs+35siUJQWhKih4mPyOm
gahTRAc+LMjvNaA1KYigMi/nDJ68t6FIp7IAN6f2Wvisd3RFBJ2Pi9DRusFEbWX0
15HyBXVa17bNLDDREL6RoSFoSYPhkgB/qzQcdlAlO+xpidpA+GlXXoMk21tGXhm+
43OS234r8wLX6iksgVtUWK8fJMdbqOBF8yQcjP5gewDOKsu43Tz32S0ppiczPEI6
tQHTIa4IaZ/xBRBiV8RWzGN2RECkBVuPTMJcNEqK9p3IuypZYok+gWg+RscpmjCF
mv9JwsSJ0VlAwMCCOcBy593HzT4MxY76bW3LONFepmsU4lnE9E0TVJ/tstztnylq
XD25I33fddP6e3P0+KZDRVXcZ/Zb2HbiTXmSQpHix7Mn+ZOSd1tDuhpSk823vfQo
TA1XXht8RYaKxi8otMkYHxNS0FYGTu8dT8pz1mxnkJRI6jTJZExv66pS0yccrwDa
spwcE/qAvtldF+Mga1ndY0te79qzGzpvgRT9+5XYx3CzPv81P9edGU2yMQFEsRXx
+yk+pEsZWiKqlsPXagb/dBP2+70+V8DuT6m5ScKwz2BOCLiH2pE7TBUtzkUKJOGR
gsbpGeCUuZhNySen29LRyS/22Ryjb0fkCrkGfkJg5jZ/RCIDBxA6Qu0XOiD4dDTw
/bkWSxjNidVg8SlmUsfhVWm2gu27TZedOnWtB2w4ML5nkYoYUu4/M9weoYEGBsF5
WBuPLwI7IVOSTmtIH/V6/ytN7GDaJNVoXHPkrtB6L6EJzdsTDDGOrJldyS2ERrVm
wEtZl/eq2t8vGLYtH04j58z3Giv2rHbOU2L9bDCMMdGH/M1MXb+ydh828Ncle02X
Vh1vrKjh21wqnLZVhCFQ7D02++lzzsSdeI0aLmL1/EtCDXGGV5CPSpystnzyaaEv
dlGKW9IPWN58h5sHFiVII6QNmdyfM5bp7yXTQdNyGL+iFdwUkgSBa0XO3AfoB/oX
Rbde6wERFDH6kiPuD0gDdrVLKyiS9NXUzBGnv89z0masOg55VrHAfcQ/4axhpsIj
CKSd1LURXr/e3X2xEBTpDIA3JyguAA9C+Ma4EgBN8u+YtX2rmpI2twNXiUSm7FjB
H31KMmATaPlahko6BgumsYoNB+IGCp0jhSypYlDiIeQjdkQX7hUkZvU2wdlc6ydp
w7hQvOhDDfbH00W7ETzrIp/9Sy0w7NfoZsSsrXOKqo5gXpCrTp2CTYE+Px8l57RP
HaPI+s5J8joVCSZS+2/k0Z2KRJ3oE1jf5gQn5a0a87dhAHj7UryXmaAOn+Wt9hjX
uo9URaJ6K3jW/BG6P9XSCGP+DLwcBvpK59eQkiuZyudJIqFaCSTKRifpFhHlpZjT
OQ7S0AuYV0Le6ghmJ9hHyCDVEKkHw7KZ+YYl1E3DSSVfKGmuedHlKVNchP1PVZ4B
YQ8BWo6bTK5Dw6gCSdJmrMqbg5kCD3DFIh7h3Om9Yzq7AYmUPolS/PLRPm6r7WjN
15qvroomQSKeHMgpn/9bVZF6TzbPrGYXo+Cv7CtEOKEOEwtvRGNkRns9EBnNWqvm
uwA8fqy9e9yVTYxwyPKV4YrswsjpFH72ft8wtz8Ve9VRPR3vo+39KSng/z3EjOnP
DGlFppHQFTJ3XU+2uuwB+yg5Tq2hsDIvngKdUkBbmRej32hEG8YelkkGdfzCqdCP
dMqIl0HrGtMs4I0F4Hy54zrU5uMuOUKoQ+lvrT4eXdlU3Jphg+r6HxwESIfu6zXX
eq1PtTfxPOL4dYYFStkGAdThX8gDgjSKLJ4neLIsKmaGgqwR7R3N3gakZStsWqxi
CCaAu1RhmPwPeBZ0eqhHCoMtUwAKNuWlDpPwTklJmRncYnFouvpVdNicZnk8+Ffb
appHGOiUI05xjO2/LBQbm+L1qwjgEEDI5pZy5BAY09t51/w6lzVbWxoMzBJk9mHA
jvUYdGtZm2ryW07vkqp1odRVK+44pVjG7ohmRTPIMqzoxbhcJ1OvspsMy9mlOhdg
fr2cdjpULzUQBh4FGrYN2qXGYAH3ZydH8BxDihjjTW2Tz92J6nBl2dpTEA+KV6IJ
Pkn5dByXTiqLaT8GXZU9vb3I7CyQbW2YwVrnA7FkwT/IsSifpVjyP4/T3TviovGT
wiz7/vQeGH/rMKVwRF6EWXmngD3FCzGXkeTpby0WAU7k5NgN6HvqnMwICSs25KwE
qMTucbz236tOil7rrNSUtXC2W8v25MPmzIAP3JFDC8ArL0NIbmZPzT0IQGflR5ct
6wSPGlFbnMQqM61VlsZOco66SI73+A0MPZKE0VtL1xMkV2KFqHIj9Su6wKxWsmmh
stA5lbQrXpVkS4O/vwVINNner4lWVEf/yf31b0udLvOfI7zbg/nbhFXyvHPXMyHX
A1hVNWfV1jbbsEChMbSWvPMDA2PGheuapnj2oOmbV3IYeKu1aeqTCqFimDyDy1vL
dvSrQmC03k0EWwlJvhxyQ3cO6wRL5XFk6D6qKD4VqHmyLnaXmQbDXSJGOLKbCef6
wsBkpVtXK52/4UepwXAKl7T7YanBBuafMPBgoRrW+Dy3ncWgmU0A/2isFKuzFxUZ
+NsbYANk678JQkVwCzSymdXij5dh8gV67144U4gB8FDNEgbOmYMtxv/b61q7iP7K
QdI7Qkb+AMH8vuMOmVC+cn/4UQoa71mBEL6K+TyvVhKPiC/BAEXntYjwQpJB4noF
/ajGvgP0iIGaZwXOZXnXbVbwJeigQ8p4voyt46+ABi4agkUSkH+dqWY6QyhxkibS
ACes0Bn4z4h0SLuQDneIgMFLd21+mqqMmXRIzmGvP3CQBMkFuDd3Cp8Eh4nNCbUW
r0BxFwIjnlIuQ3Chph7N8QJcSwg5PzCMrX4mc+yo7BQodppzvGo1hiBrsLjHdnzA
O5cMsqUoDl6bL7RZ36kfcqpO1XhWfOAO3OCirBqbFaC/1Q/Ir4ZmBjQ700WYO0l8
utJ/31I9lk3vPLwRU4/oINH2GoXpuD+0BMrq4Br5zwo72BU7GoKlrjFmBnkealPf
d944vqDTuXBINJNazPUvG58Htysv2azj3REHBGCjay/e/KALhtkBv0MkEYS8CGi4
utjGXi3DsqRb0jJK0hwHSgmEXoF1BItF4+11Vd8ZUzsgqLpPEeMx1Z9KomTvlUbx
36v+yYg0XZN7EBr1q74VJMB6PciFqLl3Hv6fNdWsKJdztgSnop2GbLH8J20XIxaV
9wkQ7sO9yzzuWy74360020c55SvYdLdxcPgu2HxLkCLXGapYsMmoyDgyH4s0bZo3
gjmdjLD6Pt4JwaaCa+Bh0XHfzMDh/5MOpULMZprcPq6avyV6KuiqpabRh+2mtvl9
efanc8j28LvpEeyPjQcKuEInO7hzHpO9qA6zQt78XZelCT07kI5663cabA4P/qjb
vQ6TU20VUK9yXJ++Vgm+kaOBUAAF6Dm60l+URtEUKNu4zG4WhTKmePqFq4U6BqtE
auAD+H7mZ2rqLBTfgopSqd9iBubL//zqXTuKl9hKCDAEoFFO4DCUPthdsC4FCXTs
upZGO8SmLCYOx3T8DvaiZr+s5g+QEhmDb4T7Nh0dUMfjMpWgZHxe+MFXxawJpFM5
s3NcT17Is2N5khk+HmgPHvZPZFm95jTNGtvATDIg3w23l04+Yoi4mgfkKK1GzqO2
Vq83MojzqVYVMdZNl0T1dzRoSr67R5sMa1SExGIV5lEkWP47CVrm4bsCVtFo4Xy+
KHl13/6JJCBh5xu6g5pgGvQzvqENM1qky5bq3UeBp3ZQPRMWUGA9ePrTjI6ev1VR
jFeAL1U7VeaXXhvqqYu5nlQzdQ7In3rW0kpPEfpkSnWKWB4alqWDa3imDy7BQVSl
+Ds5GTNRENS565UwO+Mbi8NmNLI9gml1ZxIN2C2J2dded+cqBXfshbi4yc2D9yXy
48dTSZnRx1eZPTHUeBoh5Vc7XQFB6nODXKWFC20356+v85sN0MV5Z/UOZl8d0s1a
je0fAlLw/rmcGKO0pM3MFdHoiZSSu/G31lFfBS3j9R60ExriaM+hVS3HZX3KkFtg
vAJyNO6GGoxqOiNSfNM90G5gazUM+ZfJSRoVf316+G31xZP7m2GdjTUg5ElW15Ff
s0ekEwn7k6HJgCbPvdFnkwqGgdyvl9yjdQjBad5JdCH3kMKeEqQKIXc9U8nVVsPb
4319Ndg1EvYuhD5mC/Fdd9vvUa4of52t/fejZFPw1EO23DEQa05pXCgl+k8p1vR9
mFWasNrcTViMmTLb0YhzYAsvsmNwAWkk3h0CbErGFe9/uQ3z4NMhACd/CvwuLfJf
sepcPyzqxtGuCI7u3etLY3XKtmaBO203nSi9SQ1hPqpWEVknjye3CaBR0+KdM4T3
Og6khl37FwCKs2pvXZjLeaqhADt4FJiMstgXhX/b4HHW3U6xUeHrp/yMqYYc8kq3
NhODsUhsCfYFYgd2xNO09NpKQXMq7KX+pY4yFPgyeZ5TFRdUclVg70d8Nn/2Pjdn
ehK9dHmroitkVnb+mepwbdfR/JE/BxCT+Fa8BJA51cXvjSxM550biJPxc1UmeZ0X
wlQ3gZSslxlxMlNnVFzJjuXRCpjw+37IGQge3Nr+UTDoOVGquYJnDsPa55xC2L5f
grlX4HRRAd2wYRr5ZjtZHFLnNB5jw1Mrro9S/fcS+3Y2nnBVrzF5/F+fqeT2dsn9
BOo8f7FqgmJIlPrrJrT4mzW3BcKGkTrIaXQxOzGlhljRW5UXXhNg7HQtG38WzRtW
iWB1SjG4Hf7P3cM7tqIFsRV+RX5eyEm+229+lKdgAVd+/AQf8YwZbiSLdL6YXtl2
wZ1Q6qJnIvif0e75h1ie310/rDst5Nk+9TxxoD4S9SU9ntAzm5J6UnobjJ1rtUPm
348AXRUda2T/X+mxz8PU4YkuH0oD09BegBT8P7J1JF9jQK4PpihIjV2v3h4LBRW4
uz8db9U6VoNWb4Y2vuAUsj9Z0gb+nexyAV7cxvUxCevJB2NCt1lwgr5jy8NxvhZ0
xVj+QsKiZIxRJsv4CRoYKm66prG4O/1fgoV9LY2/HSzQzMxCBOwhkeOOyHNYJZhx
Cgck+Sq9jUSn/EIID0Wnhzr4QTBBWdbicwNBBSCCLhJPLdT/KvqabYWf/ob/Hgax
3lvVBbDN3d53QuRNpFNPp2IbsZn/oswuHR1btOYGr7yO/mxtI9NJIsBzV5qDxqq7
FQxx+XzGp6gRcSjjvjGNCZyaZwY3kV2CIIVPAH6SfQ8ZuZlxT7lrJzvCufEmNzij
kSzBa0XPR+j5zBX/KRJ5awxEVNdX0qk0F5ZZlzxGSjIPkDy1yFqgiUpplW7cewIe
TjSvV0+QebvujlqvYLKHKsPwDbXNZVPkxQv2ndhoO7nyFEV8MDI/it/xj+jdBsGH
UfGAkUKwueWqRBah88uFj23hrFB9wmqNTw7HrjojJE1gilj5HzPdZN3gru9rJ/vO
qYUgFLju6OhE68FbATy7DLx7BY04f+rg41+F23e96hPcD9EomZT66KUtvV2tREyv
E0az6cbh3WEAtk9b18vVgYNMzY5wEAFlT5ecOkx43JkgwiZoguIXXZWFdrQtEW+b
0swCX5+sGmGv5Oa2+Q86yL1FHCNlwREE2t+4ImjQeAVqiZi5xHnt6llaKDowBhSf
Gckgqd5e/tL0VQ/AJmA5YdYw9fCRiwa9VC73hNWKEZWZfvikqYM0GckLYeKs908y
Jr4+x/OyMXxlp3lL4PQE46wDUopymkRzmmyjp5e2Aco2JpGdlGW4yR7iCaP5P438
nyGxMT3VFOVejtR2UqgX9nK13q1o1PHb/CrXFW/wkW/i/ISKSVgJgWHA8ZsTiaAz
FUlkvezDwX5vPBvzC4FYHQw7Isb3v+6ERW43y2f8LJF8n7DOyjNm9nvXd84nMf+J
yzK1B/wsvFHV6JKxU9ILhzwzAigGYIp/Y4TnWiyrS2rN+GM4Tbc65M5n56XOZ+Mp
q9u/UUmO05nWzcLB5u/L+74Y97dS+kHflFGGDlxeXJkHfAQJ4Nc50RGaDaWGkQ/B
AGc4507CGMC4RGmnpj1SOmABebhG4YI1Z5FTXytUrTuEyoepv//eRwx9KNoG1ngj
PCm+dQ5JdDV+jyPPkCsPLszCwsZbTzxtMM12cHCTojwpAdN/GaU99PC8nQRvakYY
+/T8xhfo33TfXYvh2nDXskLojlZjHmcEcjxoUwz8k3T8jr6lvIQY1/aDK97c7jf2
yWHT5I9Zf+ZFQuqMrGTpSlTBaduji+kT2DsyV7QaLJs9yMLkGihGSknhWM3dMLEL
fzi/zYUn10wYKUOq+wqbCCUUyttoD5mF8AvoWQvJU8wwSWhdV+Iofq7UZ9XnflCG
myAWR/vjM2MNPduaYDp0KuLhTjNLRaXRQR9Fzu5e7qSoGAYfxkyhupaur9vY26tO
sayGHzpOf8VMgYXFGi2xMV9Vv+YexIGJf74dq9JSB24DFLCe+Qimgio+XYEzPcmV
IIZyWYeGOqOHSFB0SCObncz++cVR7yq/x8BeYxUW6xIM90jf1zKEVPHFbOTJpegF
L3U7DPq+wT7t9D48oOxMKc/FSUs3G91R5rZm6kK+ARZFjhVIYCewAHVqR2bvx8Fs
0wcK2CfdNAQ0tPmGEv6R0VsBKLZfiXECvM5IXDQikeqo071fgjvAaCWa0nH7Uhg7
xuyUNUd1JnR1jxnSNC5lyER/PrWehVdStECM4cchSqK8D2dixm9dKZekVd6kSVZP
8BXz9SzCmPJPsdWe/KbbT3AYLtEzXPckIN+84uTCwphDGcqszNu5RmhdLbp3RPZF
5wdzuZlOOsW3tnpSMfEgi+fCQCh5XwD3s5owMUGvBfi1dqJy9aFZM5f/HIwWeg4y
DOq0OnKJNOdcrs0GbZFnU9ZGFV9EsJvj6Nkl6b9LdtXsmal0VyEp0MlucKtw+k38
gipiSh5yH8k0vqR7vTRzeBiSHCgHA34YCuCxNIbdFObbhi7EDRXif44x+dEJcJ0i
tAmMMFo0/+yMy7yL+wDCCT8NjEPlqHg1kTt+einZ0qnaRzF8sS76PcK+yTOCWp1S
JupNFznMhmBn8nwTiF9YoovnotysTlYJENfjcL6Ok7XdWJajeKQHtA3UZRdy2iJN
crUAG61VKZhh83bJGeGHhK8/d/mBIMThltSWw9p8xw0pc02ZqDn5bY6Ga5A2tNsK
2kq2JkQVUsbObBBGggtmpI8cYF6KqJEOOJaitCCjUwycYRIqSDB3h5v58fBiopST
17dHDy7xDxAYFU10kWJsgEnppYlT0a6P7uJSNQzq2VWSdKpUv6ebh0yonf1pOzIk
yzIizzvS8wOKJC5F4qiPfcKR/w7B1ClYX36zpQ/9xK/o9eQJNk+xmpsJbvVwn7DF
8vDycns1GNGWxGsISFWfTlCca2bvzxRNnBvDULIV/vb9L9qKxLMldGz0p+P7e/+K
zbxLtKYD+6d1+lcimgG9yMX95HWhmvsBdqAHZNm5tHGxsmw9CUqP4oWe2AAayn8W
083KsjHmpBBCtVpITfCB53bcCertTXWeliCZArzW8wZoECplBQeTxX5HEeAnr+Vn
DnYPcq+KjMeHWowNe9DUaFdXiCJ6UbH0+ouFCu+WGBs05E7LhYIVTlYPnhafjLHe
YKNC44Qky8VR2/ufUREVje85qrw3qJ5h9zgMYhnobU0Rrf5yg5UIjB+XMIaaIXVj
u5/QhaSAFiljp1XCxH6RzGeNzvUnO3IEUgY8GvXAMEy4fRNijAWM0M/1MVUl0vrg
TmhZN+sACO08xCGMDmHU5wZ/OT15H91GHV4BLn3qJJXyk+c7evudzhqFVx2WvZ3e
6PvLpXYsMnoJdIaTB5JM4WM0FaCe3wgat1VN8MRoU834zdPg7LQAr4+i3WRpOi8h
gzEUJYUWN07kATF7rlP24tNbgN7bd1uVgpRvv1xXxXz1BAnE+m03iM50/jGJlJnx
ornqHlkS9wsvpYZDqBgwWskeQQG/bE8uun170oCQlooEmNoNW+mESKlyLF7sFJ/S
LrTGq435GcaBSgJlSLPwWsLEsLVSmI5nqBukDLOpdnDl0KH5NtTOsU4O/CcyHM/M
jSj6DGJuDB+lB+EtaJI8aukFH8V5k98rJt4znVg5TrCmluuQm834N1qlYd4EdPlh
DUu6s7Tp78lcWJfKix3Eo1VnddHAGpjTY9bpkjKbB6EcuuxXn3EUYwOU2WLiZZwP
TUuV5Y3fSq1yWj9ax9C1+ZNYf4ddQwxF7p1QHMK6R/Wb/ZVXdHKc6DL+mOjcNItF
nXq/2BI/Ai//2zob/OhtTIEk9UD83LpXRtK3rW5kEaBgqVPKa7veHeIka7F40zip
EmnWcTgYkjFrqiFjQbjkkX/1sCDaC2OlfC54VijVy9CD2xo7xYxHWSOa8Z1Pgh67
dVHmcBZtUXyrJXpOzbw6E56mOuXlCGOtH3B4Uy+Ehl3973/r572ORsZXSaMla2rY
wcduytrmMBK2jbhYHtHoqClNjcC1hdvXgruaKR4K/49Og62/THOo5bbmbIb/NkB+
soHNB2vwUyTlAuiaH6kBlwu0PceWMRDBAuEVO7f44eTm8VD+U63jGJ+Fzt0qMI/1
PYRPH+KAuZTxqAEr48IBkJ05Ty58791hpQ9EbXBfJt+8Y51iILO8Figj2PbzO4pI
3CSJxBGXZ3Wgiln3QlY5kahu4DFzT1CFt+PtEjxCRCLF6hURCc+aeyLmMo68U6Qu
h1/omAop/zbixPHXkSZO3VylAHbnZTbi2ely2szsGlHCMKVqzXagAU3xxLiPaXYC
x2MyDhal7fKdywhKYZFUhmpAvwqLv2RJL37IlMM0VP2OJdUEvjJqqgSDl3wWVXO+
yJxjWWX2jIwLgp3o07gwUWvkxBHPElv7g2UEJGYDK04jVnWYmJ+hYEm55ZBJUkJC
LeZPxmhYhlvm+aBAzUa8bblAjEjpYfRYZK7XZqGTu2Nv5RSKLbFW9sBiq/MVfc6m
70lfs5zCYPysifiaO4a3MsSacca2/xu9RnWR2NY+l6Xrm5uTA+CohaxfQGs4Xg2x
6LAovRK2VbpcT/RA9semOCN/s7QEYqvl04duLQTtH1KTpIaReHRZkeprkvLVkQyL
GmKgY8aBqmR5ZxcfaCK4uqZ1VEEi+BUIEuOz2ugeehKgJdptfwe0tBUT2+jLNFUu
ANGVeBxWNITq8k/i1QZeijX3ic7RoO0eCbkFfwW/ZvQRaaR3cg0n3NSKN5o72SPj
0x8mUBJeMiS8vRhZIJ2RTQHE8SKyAmZjjopKYu0erDQBaaLfrL4x74Xwb9c/1mxF
s6wo7kE250wTdqsmMpU2NG/+7HpEpVf1W0Umj2jy2QfvJlh9NN1jhPMjT6yl9Etz
LoEX30aB2cTH+15isKbqrMNgd+YDy1YSFi1vB8/+AjS7i9ZmipDK8elOpFXg9Wbx
OurMIaQ0zlDVBxJbdue8OjrZOs76dgbC7sPGIthC66oe3l9xL86GmxvcEQ7o2S4T
TbnuXUfX2TKiu8ZI4lkIF6KLHAMil8B05vENXbgxx2DQe8LGiQ34V+H7Huw+AJaS
c/DvkKbJQgP4h6zezZMHvqJXscgCj4ONudoNhxnTP8Q0sbhtc3Cz+cuUGoCg3WGw
T7ZTnBrC6efKN+9QncY5qRVTdpFTfhzDmvCfYBSqn5yCLBtPJmmF0Q+e6dMRMruR
kNyWGoN+Ms505Vrsl9Qnn1bO8qW0QRk9F+k44UjWhth4NcoAdIItwzQntL05ASTn
5pZy/whGHykG94SMgAlO1lYAre30daN2sBX4aGDxXZJH3OAWSKrNzl9TA+FGR3H/
BPgr5bK+F2OMpTZg0JQ+fwPuCViGjE9WrT1g9sr1vodnAXuxXvpO4XIqF9KVtfJU
+1FA1Bwo5SMFBlhIspDq4IUmDt5EckLYYRR72NDx7lp6rmR9c2yU3EUwr06eESfM
jpjc1vKmk2+m/G+FTPJaYL5RfCkIgqJqSoSsv33YsPOlhycZ5e0dZu2k97WTueZx
ulUyEWLgAMWa7051hsjDDwgukEHPz9WRlcabH9JTjVV6XQ8lCFXHgx81ZdLnqpSJ
daGXMP488HpnXpmTq95YW5rw6It1NKLItU3qW7egNXpk8uTUHttdmJMPTpMkjqB4
QMXmQcqfZjam8WbeWrBlwUW9pF+4Kmu/h9H9lohrVget6trFThZb1bJ3x2OPtD7I
/Yl4UxWoCBlpN9cNPGjWdKcSRJeqqaUYAdgUZoc7WTYoei1sx+iiUBvSS4EKy6zl
QqbHT45DUR3esskfsj0YdPci4YIZCRc/4ZEvtMlAic4pSJQ7RXrieOMmOCKuy8iD
OOWjsHMXvjH15LaH1ffmQe2b5/qukBgv4N0TLFBadQCG5h/uffux2JH04vupQOoJ
dof1Fie4/XNrlGXwcD8b8bXxQMqSRijQ2FX8ICmb1+TBu2ipuxlxdsQFDUjK75SJ
mn/nAPM3jNvojwVxQqaKRigvuFVXr4SWtucVnygl5fdSEvh0iedAEyiLaz3LQxRc
/hD1xTCovRxN3naIr0xpkJyVR5WU+JeUQLXbdf4eQ8+yNvrUAtXTRLkPn8ORAsbW
BaztCDdxXXLYgqoNqVDu2pJ1xeWop2qCH7MMqgVWXLkS5+1Ev6OHNf4xya4fB70S
ECnJ+hZRFtn3ocQX3pCACexcNPGOKRS8yJPMsU91sFKKkeFurKaMJfOcGO4gd8NL
NZYT0BrnzuAX6LXXgUwAYiAAp6mtUSzP4iClIDXKDXVBAlUrrjvUnWZq+lZf6eVg
1Nt1jD+5kGBbQ8SuQkopzTX/URECYm+BiE+7URPgOgLoYlKIblNA/1/fqVGe/5Sw
UIkeQ+SZyhzDczgon8oTFKY2M3lQbtRmwckoOipgrpzAQEYuG7Ty+SVOOgKXAc3u
zkrQ19ADYktFCjgU2kbmpeOGN39JBnaYbkE99PQEpxdezNkg8mW3ELDW9Rs682QG
RQaVbuE1BE0VZaQn9mYdbck+62Z8BeS/oIEcN3Edlxj7lwKwZ2qBl7JejMHlAwYp
0M0xRDcXl3ynw8Tpo8bAzMYFrYZOH/AiLVNifuoTrTowp+2m1911bahoEYHTspaM
xR33GYUaR/MQiZhQJU//feB/2/dl054QZjDNfqpe7iro3TfDc5bN1OtJBkEK5Wwb
AlOXERt5vthxpY45jhZlBWdyae2eso0XVAu2+H0YUcs1jiHiCLEfPZfuTOlx51N6
ZA+1YH48sJh0lJgN3kex9ty/m9vS/PsmSIl0Nifsmk2zO8is0uXBE5lJXJ/4aHc5
QAlUzcphR5u/woKirrBFaGLhNxhACHFLpee49/yDHUZQ3zHahxZcfipHuKsaO42M
XzHSfD23mXgV78zu/RLvpvyuZCmIpOsATLv3brK1g1FWQzqpMxPocF0Uvxzo+/Cq
Z/V/H326RZ9r6xkdLxBh1Kf2JGKKk6omrddR4KEFWEGRXdt+ubxnR7onW7D1t+CZ
YAF2FKjLgA5IVZe5J+q7hbPIP0GWNPWvbGKVPtuqbjE+DDBHthlo2s2elid6sKPo
1zF9xip/deEbXyQ7qKrgdLjaXkJE+eCsGznrN2U9FOzl8FSGQT27UmbckQJYd3Zm
rjfoXyoFxc5NEJ2iP+ab+82F3rr3jj69w2jsyBHyzt7VeQkhwZWYw+N89O1ieOju
gar3r8qn51U2oO3db0lgL8n4CKKeon6GruLS+E09T7lJv2rxUxSQd5n1r+stNS1O
h3iqwREBuKc8fPWoUdOnlXEn16GNz1K6/3f6i5TAzpQy1JULfT3NpPjrZywkpyth
lFmSO2Dp8UNDwDmBJ09PJUsdRHyyxUuPE8Pkn9ARViL9EMAWB3fjjSxffA1uHJto
VjbGar5Xz84dg8/wZZmmAg98O0doYzwrcZxIDO9v31rLZFiJKwlTzPwUFTew2es6
KW0geFY1mSq4V5CQLcYyJHeOq7ocDwj7o066XJJy207aX0qEiAS0/czHn2jbNztq
a8zW+Dkw3gd21ZOZayjiRjHLt8B4knGPsZ+EQbd5Y/aaALdxCvChi0dd0+93Vu2Z
Gp1tRFTy08kizCA4k3GkukG9GBX4mxCWT9Oydd15EfUlCBG6gI9vf7uVnlIrGtr8
H21lys4l0jXRpqhfnNhvKyqJzJzo7eriShiZM5Xl6nNKO+qTTtCadXmnzBp2ym91
j7qh8I0m4FCcKwgt9KCt/uD2HlqrQ3SCJLwFng0usZNHxiggJEs5FAusGfkz3kDB
GeoNdGqtxCdtYf0/n2eqpRZ/pm1fxf1sv+Qc/FT0fixnvArDTyT7hAG96v7gNrDP
O7gbVniavO2SHTfcOoPrpscw8SyDeC6I8wGEVgBIbHyN1iGkmX+G31CKbleU5fR7
bloYQljoHI5r8bVaNMpsxOYRy7qnoSDr0CpmRiAJHjwZM1aey4kjB3bQ5Ik7/msI
16TZ3S+zB2Pa791DtzXuaYo5wDCZif+Hy0weUGArxfqvEDngVcHJsWheGEkfPqne
coYW/jt2m5oIOWu1oNFvMTi/vOw41OsgLdAUh0nL43ibW8QUhAsehdTdAengxbs+
tSiUmLxdpQEcFOz0BkiTBkrYPGKNitTBuLdiStuQqVd3ZTr0UA9rneL00s+x70XK
fSMsC1MhbFkY3LHTxLHmayGx7zaBftWD3lAlQCnOC2VQtntF5EWJqzoHvUxgAwOK
ZpLPfVIP1TiOktnj+J/VaEdIw/V6QleEEaoVx17jjJEg759Q5syv+XnFJjQhlT1W
NXxfxYWFt3VRk/PI8i30io2l8x+vbGREtXNodFDCAigq0DWkHXolpcTMTWNgCdwt
NXpb09f67p+Psv63fN/glJqtF9w4JUHclvmOO4VoWF5XMVDuZfIX9UIR//GxqukZ
1ixHMGS0P+fFAHVLNWRZLIYhIWVmmQRDLF/+NdtgLeo1bZS5FYeE/Y8xdPx5KONW
vWHbMW1PJ5yEYEiIxZLAQexM8APZ2S928pqqiG9Pt9rolwPx6mMZTdFBXl7i3dBq
NtEccQD2qPTFLigRf97vd66IE/qezxjQtkw8U8X+jlHRvG8Pmdiykq52v0/zGzWB
VUUgxa81dTJK7RyJ7flQbXFuAh2VINQweZPkrzOg42uC8YeWNZSi2irr37pnXquz
3mFqYQX2UUpXKMymgAKunHVmWXtUfkRetFvOnEKFYXBKhsapO57MTT+LW/HzYpcI
v/szBRjpmULPBBnbbZmgv8YmefBAc6dIhh+VPMiHMOQauEWLDp6gc52tIPzRfPET
2l7FnhPDOu/ejNCi3ncwkYzlnV5faexI2IZUD/9f7CcXT7p2ENaGiy5sfYW89iQx
baTmAcCk3HnctUXI1fux5CO/Yc584fZDPcNZzXl8cPFF8EAq6sp3ekwMzRcIZd6G
rKQBIi2V5bu+sn7XFiiBOCDZ8SIPtdz/vZUZffuCOlCaf6Za1tIfCVUPj5NFMwRg
q6fI7Pa90Lb0eUofcCSVIcwYffVmu3aLgo1cjgE431oYAbDhijmlONMf0fqZ4PYY
lPPkOWebT7IjK60cIxuTVP4sjTlwzMsCX+U/Ng9hGKdFA3OP1EwVdzJ/a16usuW4
y7UDvo5gztp+vKJobruwXAMn0Lqkj2mRsnSsJmVr3KrJssF/iyFI99I0X1kwN7An
mLzLSntc3DMsDyeler5y45pScyBusTywlM2vhV0KYA5m8q0hIk955XsFWu77Hl32
UCYUwkCtVz5jpVhbromrCA8V7Rnu5eUzZ1Dv3n9kVfXlcprJVR7FPujF53HKJvrF
I0Hm7jR44XaT7USx4NnBAHbUd9XoHruQQbGOdTdL0LtTt37j2WPQjq40yiqPbmFz
DspdX19XJxHt0h03LsYPx+lNLuINiWlt2UNjkE8LEDbFYbg1XJyWP2rWvUvXiwun
w8hKtNXwE91DUMefkOWEPHJl/NZCdqHPZ3CwyLmNSfCFpAn6cUnk9OMxOZUe2MID
+nrdNzAuJTY4jM3ydVjyAB7Wp8fFOxRZ6ZSCmE/HdvjgO8ftURGnlEn7C7+ayqRe
rwyEXrTvFJyTft83AkrsaOC9Apxqq7UDvfYt6hu4osRxHtfEh/R3JftHVLTwZXMV
+I2T4FDiTrKmcSw//t4w7z9tPrwLExWUBwag6kYieRWGE4XtHwq+V9lGze/0s3Wo
DteEGGx76ndpEZEx+R7ugFBCrk4mri8jSzXTOBXQ06DYYGLqF6siyjnUv0yrsl2X
Y+Oc5bXweY50iOirPluUdCrXLc5EaK47Xmzss+Dc9UU2Cp36BINySyPX72VWKpno
vfs+fw2hu4EZO7dEwIysRNhI7OAC+klXx0Mp8FRRcKjgTh7R8RV7ThKRxI2Zjlpk
wftMmpYSf6DMZPtEFkWZZnNO5PRpA+9T/wX+grQxxez8ZXZZl3BWw8HsS0+jWL8q
NZQOXar7PSN6daizn6imwPGc8eJOT8/ofmjIL0/UAQ5kSfe7TFCGm3CoVmVBJRaC
AKlnpc2+cJhXqRUGJOkWnpokY+iBvyZ3LFFkn/FR/UHAuRkDQygiHmiGK7Tj5pov
pdf/swFNzGRXreeJQD1ITUcNFNPIKL4Pp7oNAvoeI7brJwhtFzlpjrAb3COLABrw
G16noIBExcpXIsz2Gw2r6z4biM8QbXxX54M7TIRO0cD2UqtFWfAjjVwGpuGQ7Vx6
rznXPpm6ovOVCB/wlmZKYbtOzAgisQnnpn4aG5Jv+g8g6erpm3BUoqVbDAH+g5LX
fiCJQybWD7lF64c2KFzJpQoyedKZa3LjkNP2PcAPS9T0F3IthB2Jk3w3T1cbHK6O
gMwDUJCQdd3eQ0utObD8ucmE7tMZgvDZTodMdp50vwZWTCKn67gjVI2IGI0v49Ug
a/6Tz0whZWtZkDRUmYbn+VfmA9lbN1bTsadylWk/L4X8ooUdiQ3GkAPWoC7lN5Z3
D38pOS/7oZGaNhtIfhdxo5XvJan8BElACS/berLnZ9zRz9l/eKk2/Bdb3cU2GMrO
KUxLF5dU77cgDQHrsE4wARlBlpA2xGNezz0WF/R4SC/WAunoIf1WQFAdlVHOJIoU
vnBn/swUD5oWuc0x2Gpc08mjwwF1Q1E1/tTn5oIaIjDIx44N10MQbUyA1cV7tJh8
+iddDvBbb68iuk3SJrFeOAqR+Dkm+oQtMqlpoGCzuli3AShL9GWnKbbBQbtFV4J0
LO+DQb9QenuPcvZ3nsa5iMvmSr0+bUK9PQjie3nlkEr6RhVBEexpZV8pVfPf7N9s
O2vAGFcA8VTUPXc0VmITev2QjcViVkVUhTyRaoaeIYe8Pqeqysy4YxkpTIhF2vP8
Byh0kI9LWdhWCWxKTZJjl/RgBo1U+c5kjc4NAjTAyC+INZaK/gjXBQkyF+EQNUbX
N1m9uKJtRt7DhyAlBBT5wiSXKT4riJXh+UfGv8AQnQV+btiO7UvuvkhdMdTm5f9i
K/uGfHcayJBINh/KbpS45e5c/KJvEAZCNMtzC030WS2Qi736qSkpMTbAaW8HTSs/
h+EXYyFupUChqunDkEkSGrD5HpAgCHbqeFezK8uemWdyQIrbZzrPwk0NWIU5iImT
MaJLaxSTuCWeFtLFtLcAa59+JvYFVUXVVCn9uQqAlRvfV0ko6DtQeCyjF/bTGNXb
Yxmdc1PZJ2QHkXrItGFkPS/fQPNARy9M3UjYgT4zGy/V+JrY5LBkUhwzuLRbRtMF
P8EoWQlGnWsasfOseQO2EAFo4ESOpdfvS2Lba4EYziHzbjNXfIhhXk5d99glnbYg
k5uTzN584aN/DxnWmEBrdgpG8RmzwXjZPezHRqzyZai8Ahkz3nYXeJSe3S3fsaH6
W3+41FxERty6i6gx94vVwk8j+1ExOJKgIozOjLWHMoRYclB8oDhI+8cVE95W2h+C
qKVY/g+Eftxij4PulYr09T5/p6hqzeLOUfxjGhjzov93E8ps0vQ39e/ZeQHEH3sP
37SgvF10jOOzotkZH3SDsOYExbqhyPSWqBrBIVqQw16sNVx19UTHOF5Em0BYYbBZ
cIfrckcNKzatSRk2KWR+aGOhug+ki6UBO5lEAyvKntT1We6IYx98VJ1jVCRM2oBq
Z0zF9poF2TPqN53SBHLK9cevQYvSdPli2WQ40xzPlwphi8Mz3EdXfYX6RLtJNZYU
HSDvr46mtkZ1V/RkzYw00BNSE8aUlihp/3N+ShJH3vWdWiaziYWgKSktY1+ES2FZ
e8nGUvSwG1wo2U9eVc0ja1xd78OlWxzjsNS32/7WM3juhU56WwVemQrvZI/OO5YC
Bc+8QdwPs0jfD+g/nGoN3gCF1S82gJma/yWYxy7eaY0c2R3SkiqELuPavVNthWD9
vX+e6uzHbYbDXI/36/F/SP7xeXR6oKMRVoLzb1fSK43QIMyHVPKkBHSb0c//pogz
xYkjVVrgihqMV2eguHHxX7qnYLVaat/+lUvL2MJbxoZa51W4Aen3lRtrHQgJunj7
OQDn28ilpZFUSkCkn2n559n6OcNu54JtYa9vueFcez/2q5Yxku4EY0r+wJ91bzaz
1w5Gl1gfitBxKls/483kVZX1QupNNCyZl1kaDI8OBH1SO8PcgrO4o2UVBXedVsJw
lroB7ynsWbYuplOLdo3TF0fy2d/rl8f7lqEpvYY/HP6DhqyH6Zfq+nyfR2LOrAe4
iuudUIeN/tXksnMsZzzaDm6d1/pV0uVWQFT0+qoyVcp1r6OKlJUZlBehQx+Yu+xI
K/+ocrmufl8dZFtbCIFr6OkAllhChlSU8xliJDsW9IKd7vXsDr3yP47vQmXLIB7b
0a2qQzb4/IJe7H1jjlrhrDEEnVUBuVInuZasD76Epdb5rWQAbx70kGEuT4C0o4Dz
DJyIU19xA2cr8vorwEK/gqaR9pMShRX/fAVVPTuEXZ+5T6nJkv+LbKUW9pm7pyZz
6fbKklAwsXO6lAq5pOKF+uT80AcnrjbwpmE9vCu1Bl1FQqgyMsEBDCWUXxNpqS9W
Jyhu14MWH6QfWprYCRbiqV8S8Y6F2XFIK4bHPrU98KoxPAGkj6lll3acp/dPHqKF
SwmFP0XurEiDobkHSpVtElSaccZlUmS4ZB09IftpKlfLmgmqxsHsR99k7ofR0Fp6
cwB6mV8Yc+U/VjvaVkkRKxAzpncsERlk7wpggxSSuek3rXmzKt25z81lDiSMhxps
3VWZCvyI+RYkdGQS/nRB2QsbhoODwDLPoDUOl7vAhcOlsUYmdSkcj27dJJkWlt6R
yKIbnG/kkL4pXQgGBAqNqKHXPzaOb1vPno9zQ1dQn276ZLHeKIYByCJ98ZbZv5qF
58HdCalTqXjWIz0ACekDedRjH9uQviC0z3l4a3hfMO7D2/4axyrp/IHfP8oNWd/o
mjfLdtJpmvVEvrd2L0bP3qldrdMARnFL6zn5ZGJCbviDU29JGHDaHlh2gYE5I2Jo
ME+hGyznWR/wf+pn5esjfJx+kFggWSSripx30qLA9EXnAxrQP4cyiYCL8F9HNj6o
D91QWhqbb8fsjpqBRt1/vlGluGtLJDZvc1ZQpGayRAWD8nPI3L8ed9j1lqYbHP7n
KnsUENJ+kInyIqrrcfTHjzmstHXyzPdzlnthy1ZLTrqpuzTUKJ357osI4ZP4ptPO
jwnX6+FWgVGLqL3gdLo9TzNTvBoypCG05j+1NF68NZ+z0kna17L6PvEpPJ0oYYVZ
8TE+bFjeR5hEfWlV1rYghVCmadhBBEx7gp3366rTJfzmEHh3GX6hzoTNMF4ATSv0
KCbBL+WK/Z24cd3603KAFDmQnTWe6oFuLlg9urdrkO4hlTlyONZaWOvjG4KU8vcR
Wjhpn2vBuX+ygoBxpKmPBUqb7FZQM4zHgJYL1U+TtDRYw2gYG0Bbc7FQB7kwFCZ8
A+pmSO4JNn3/JR6x0JJ5AZ2wzf446QO8bpto2W3EAw2VEQ2E/z6xDxuSTA6LoYwa
RoH1SY1jI4/JEnpmd0tc+2Fb8BfBxiR9o7p4IyPm0Ojjrp18lfcYO7i3/T0yn1KB
b1fc0eeL6DV1SCBMED47seTnrhJYO9KTTb9eO1VkhuN8NMOQoovNHXVEbtvWfOYw
vJLWfYP0ET5sb4M6kqbjhprjvzlq10l67bwRMODQae89hYu+7LwTB3JbnAqDcfLG
wLtpmGOH1Ud43bt9sHnveQWHCKXusW60bNkB9j87cmuBnvbMFNiNE4zJOoTDMvjP
EWzVVWkWZnKWHE896q9hUeHPgo1++cnOCB2FY+vt7cnj1s5cH/5UGWEr4bGLKn/P
dAd3UI+V23iPIh1kyg5C1F4hC+EhW3RiZZrFwAvGdabEhZm57Sn5M9sU5lM87U3O
p5MJjRcBedq5b8vvUUSnETkFQEH62wOYEI/Dcf8zESizshjlkqMWEO2x0bVKUHpD
UhxXC9IBbs6HMfsjEqLFw7WgWWwuxLvWoZqUfcwabhMDoeKHy/zo0qQRun+lueJ4
AnUywDpFLSxfyKCsc/ZKDs8qm29X10wQotfAeVs1ZcBV5koMAgv21U9RonrAEm8U
sWZWmbhQ+DDAbv5KQRj4HW/frTxkzB5UeU3k3NCRe+oIe5B/NncQvZVk5J9rFWBF
+wLcbN6Y2qm+M7w+lvtq0fCRXNhmz5B/1RyJPuNOpssjOx67NsK2mGPGPr8SmCDy
BRuGrSJx3N0VytvBcDVH0qP3yk9cOme9QJ3s1OAu/AmkpveADKXh7opBPhVyQi2O
AlchfFCOjA+pcPmkI1K0Gp1Fnx/ssPNYRKJggRHEMamfdUrIBaAp6wn7vDEVbTi6
QvI4BjWOgJrscANBZilRx9HCDSd/TWQdgEjumoyL+j5BuecddmqcrHYV/+tCxID8
xcp4N8tpDqw7qj1aloEZ8ZpR12X6KfFfyARZscm7hQyJhgGbDuOWNmR/nsQZ66fC
UbbIpobkjFFA9E72e7CdNRM7OXJrUj9qODKOMYRQ2RNXl3xJJui2kUhiLNgIK9Xf
rbbv/nW2rIEjMzOBK6CaQ9Et9qIuZMZeLOOCEWxFJFjfEmzpfTnKMnPQvXiMZxsZ
cnl3Fg3CPZmTqW/BjnndbW655qqSb9OrYcaO00wslulsR8EoFT9DldpcIOi7OZZ5
0FaBUCy9ArLibC70SNjFsmKAVq2/nSUzbFe+4mctzEaJylvYqr6zJDvH7a9Z2nOq
DsPwcroLZj7JsJUMrRhXJ47UbJn0HV7VQX6yiJPEhVv77+cOGkoqo5+BxVy3mElZ
f4b4FvvMcRbTAAmWPFmQqUkEyqah+KLdCNyRAYN1Vkrv0AzEjtaw6GVGjZL/Jfse
erNjbGaEV9LNHU4pJQaD2EWLdReWbN/T+gIg9cwmfExUIZx4ohrEF+WuszbSUItk
VrZ7yXsL8bInVZzv1G/cXpR5IH1S0Sr+NjkZhXKKGcMj/nwUCDw+Tn1FNyEwdPcg
kTFU2sWf/LqfTU3wv7D9HZmN4KJvQaAHOfWG515cFt7zMQ17rfrnz6DFDzcP53UL
D4ShFFduMAzSlyJgi2cUpq85/h/qDGvpWpFdLHMZ/er++dcwlkjpW4b+tF1CytUs
9/4vpyMa2pUzgj8tlOR5Yi0qjkuG0YgAHFJIl1RW7++myJ99YmutVL7UeCEpXrDI
54h0zY1O9stW+6LtqSRhiipSjwI9YbKpHoSO9nltyZ6TXtHnZvVViXRECpn+vmEc
wtwjHEbpDI2FdU9+ixidE/Bg1VlmcdsFBinDNqI6wJRP7xhY9TEb69q49fdJ6PMK
2e+oVTs6SyzXwwN+KT0kEG2tD/XPqFDqzTlG0ejPxmHn85uA/v3H2fCzt1omzWeL
gnWx5DpugEhxJUsjj05wH5+Jqspb+jW8nVUwc5J6rerYcDng6BxYUeIKlEBo4Qes
DnHqkYgPoYYTdSZVKhpcEWyqzWIkEWiQ388T2qWzYUEKdCglYLVwvYzIO9DtUorI
sGFFzQKHr9k0IVanKOH1kUJ/6mmoCiGNaumX5p4O82TX6Nz83+NI6G6YUXDfd3Ad
BMtICdyVUZyeNBN6f9UAUfz47/0jXheGNt13Lg6IltUdUnKUBmwHXhZQMrTy8zZn
mrJTwYVFE5ilyJ/gG/JE0zd+j7ZHP5UzI2NBFyAnED1NMp4P2qryxF5FIaSVOla9
QTXk9HWWVs+DxvmGsIMNIZV8kcj/PpXCU1PWPUDjbViAC8o1fcKSQ18n8LJjQzjt
hp85A+2rwZhmm8EhPO3KgC2F7z8E4P0eAcY2nNYzXwFde6m3zcnRMQUWX/FpHyDQ
GbpjichN7f02WjLA12zxpfwxFSN7OCJ51JoOCB8zu3UnNw0NEH1mjYhHCxDsbZ+O
nyo1MRdtR3o0eYVLiwgbf3eIm7OSx3uULRH+3lb9W9X6rC6VrB1B+dxLZMrnb0lj
ZC5uNbwBPxZgejEye1o+Q92JU4SYYe4wYOaBF4dcaGidyY3a058wA1StsXU/P02l
MWytjRghTRTT56SWFO5HvLTDQz8PhmppU3gxiowwuWFYsQx6ENxJVTPZ955s5bD1
mXoMuUuiBs4FbZ9HSUxZfydlsPV0D4I1y6WFFAEO5hljZiwzA7tELUJHvhPe6S7q
Qd5pNOZ0YGoWSdZM0tVQWQ1uV9dKBp34+7f+sqdWix8Tcum3SCjoBMyTkLIuYHwS
bJ4RBR1I6u41VbZWL0IEWA7BadWTBNseG85YbQX/5gGq0sRcGlp/WdDATApanUfP
TacurfpMRY/IUzexof7eJUCoQOY9MUNbBdLjG9ZD7lRRV+eVdU4lyZmONLJUkSy1
Hn2fGB/C0XjgkAHUOLz70E/nbsQ7O6T4HjhBinzMEibhYcuXKazVHxf0VEzewAWj
JOrA1uVEuXob7SyQ3SaHpKlNeCiToo+DPevNJhqcfNZ8WZsmBXmVUbvQRGgjECyb
qWxObDYjKCc8bUd90vKLXEnXSZ7VDqzOIXptiUz8RlrF7vHgPL142TdVCVu3rqet
fLTTl8oQ9JJ+7aWJ85GZbtZhH+uDs2de6aiWRDr28+W36Id3fhvg1ebEAefATkIC
DqZ+7iwqiV9g7SIvw43j9J/IoEdgWCXiP6Gj53JtTwPgSgBhgHMuLNvl4sKNSQLF
LpFv3E7Sm5FkW1wPrGMgT3HG1Eh6WZxkPLWqC1UcApyVXX1DK0eVqhS0+nedfjVw
qo7CPUFxfx5MrPTZkl4ju3pm48F6zfh21seR800ssRgZ9X2XE8WBFMhc4MHRfm/A
MhRIcX8BqqMO13ppB+ZH5Zy6gzCwbMeB3P+6TfIGGEeMHWVlCIA/w4PXBbQC60+l
6WBD/+w2NmaFOedCyGkT4rjgxOieWBmlD4RpCIS/BqZpIuAqCavNpBTZiMwEpnVl
sxPD5uxvijyeYs2ZLkZwjgomsaq2r9M2/FWIs+LxQDmdAABS2X5RrX1Oe6uxOpbA
x6Mb4X8ZHymt7SjH+inEYHsYY4pCW6s47NYbhy6jXuoKLI/grLcVfXh4KJS51DDW
iP7XWR98cTO6ayfD0hv9G7OqDbcTfmBD9l1ejfcAwiAMqWxzvQJgg8MWKELcWyBu
xy+LFLLYeJOSCMJO+yCQMlvRQI6h4IPnoEh1wp0Et5OBzRJ/GRexfh+cYQ6898Dh
nrOeBJ7FzsJNpP/2JsvYxXOvd5dGxTXHcJ2PKjPSGP0mSCzmIfX81z2FN5vu7lCY
WkixJ4TtXFQi9sz4dUr3WfePw03/LshfC54oJKUGUFG2uHH9K3cpQfjwlH+d++n4
Y0vyXfZn9NX4MJEnJnYGNoF5PncjYhAVGBiJxz803N3HJ0knqS/kIqL4UM9bQSXi
9AAiBJlibl8LnZzbSmy5rTTYhnKWhIfSoEgFNTSVApafPWwIZyDA/afM4dZkOTfX
VIXUBCx6fr3HXhgPHjxm8vBkBbM/LlNOCpBHzhQjAdsdELPXmqSD6dSoUhH3sRwt
zw5ybf7eE8+Bnb3NbvKSxq/+Lbj0hYP88z2gRVl+B0b6yBvYcUN0WO6YBSpS0vS4
+OjhdMoXaKG/ntaXTPbZ/IQPSblAVdfZkfpxl7zgZEl64aaKRrYevm5nkth25Go1
om/s/j3bN9obEowsGS1tdFUUhzncA5FZvO8EyeKSVBm5X2wR2kMZDPVvV31Cwlu8
hz+StjgnSR6FJb9NqZ8EkITP7GEhDvUudqilTWmBJhMzsVMrzNwf/P94woxFswJz
FCj8C+qM/krL77xFeuEFPu40KBy91nQnJdXtEQrRptPpUHTEjiy1NBEayU/XrxZt
6T205rSLk7e6suK01ksYp9fZLDWUzQysPQr9uHUlwFyNBjBCtKlnLQHVc2eqGtiC
m5X+xUouL+DQSvwN49IDoxb/rOpZ0VDchjn1Zd2cmW4sPpHXXHLn4HvBwwIT2XzV
Hw4xlcpv87LswAMPgv/rb1ToShJKkTfBD93hV0ng3KI1AWJ7ENO8kbkqXUOO55Mw
zfYSPaYkmAM1NvM5LFl8dBOh6DpbtpYf7rnbH/MBT44TwZP6+kxI6BT6zzUlbRYy
2Btm8k8t+m4zQyM7ZrSyeyJySN0zlDCh3XAA6/RPURzJa7i70EJkWwgCRjX9DM7s
vv54qGH2sJolkHKZpsgFwG47qZ30rlP7MYXuCJuziTRgynI/zlCdHm5QSyi0NPsl
V1nNYUcRSg92jd//CU1RQcHl4xKl6BiOm2Z1Sk3iBpQDhMU1IeBpKPrKlvhE5Su+
ZUELq1/VWDMSKSIGd8k8D/jfw4CSmcdRE/1MB9AWz18r88yPyFdjVUedPU8VwLCZ
fLk5oQu1CLqKSNHkHE55dEJDUYsKOgaEkDaTA9YMTxzCumdxe3HOmtmk7qDejARd
W4v1O5W2CxlvXT4WyaV9S9l10TX+sSK7KSYlaytNJyvWrQMQR0AKr2H/8TdAF8gl
ZlSaZIdQwCR9EIkG8/dfJgM4mbK/MmO1EW7cfN1dqDOGvGvAce/ATGyqNmFV+t5I
Y1NlHApP8X7aAG6HJu2hmDC3H8RiDjOfXBXW+OHlQMJ37h5t4NCZFbGfEm5YuLRI
9EqJ5PcsFcjKsF0bj1jAkMeSAvCJoIMF9w/rTolzvf+7NkaLRyc+bhSWICacrAwE
aPSdWYG8ESDreO3k1LLWwQXHRQNxbO7tVjhWwU5+hEaLQiQn26poltQtsPfVOoMh
YFE02MAVnr27x+i4x9ArUd8BWOMDj9pBVhE18o+MRzTg195/3w8iGE83XetaOjjI
l6zH0A8sh33wufF9K/xoZzKZMtKXfH3qgFqjjM2weNVp8CD86O7ueQl9VZhm30s/
WUXCLjJ6y2ak0ytOnQoa+0eMj+4qKS0TwxEjVYuthGUM3c0Jo7BDqYXGLQTvLXvs
iDXY9R1Qzv8t8p/NX22q2ciOROj1+MUgLBNyqWTj3DmNN9qccIFOCvpCesDWAym8
aqLeMIXbSN6s0y1ZaZ2XKn39hi20vYl2Y3y0RzbbKAtNm/33V4uq/VmJJmyNNCNs
C5S+LSWjV0lyBknVloIk70kHd/raLn4WCFPmCia1AQUuQCXCDyRtf8MPuDWVTr0p
+HBQScMC+0KgS5r4K8fmwi+B41HOwZN2ilIelmWfLULLSIWksOCLsENywWns/3S5
r1+o3q+qSKxJg9bhfkcTknLoUQ9it8DFwOfXJ3dvO7vt0LR8Olzu0D1vgujdnZss
/YZVlUhLLuN45X0GSZBrke5JXZBZIl8Ast8Co9B6u5426G4wh19JbyXpQgB2jiNY
IhGikFbcyeE7UNNzOb26O/Sg12Jx0iB70cM6xfx1x2w/KiV48Vzc59WRed9k7SAp
W2tjWas/7vCkpttcDEoQ2gYFmvOXoZWu7mCxnsWgALNuVXOtnEm5w+n7NH5+Q2qx
gzT9D0oYmqXW99o83K7Ye+WQDJUUiKlq7SEpOKHptZdV+x1GF9t0y0F2EBvsyUzx
T3hcPrUrch3utS0ceX5pW0M9tM79q0l2Q4DhQp63pWT3no5+xCMZHdBOvQWZ6jzL
ydFxghCgiaTzmgmmZdeP4p3sqjSGovYFrSg2l8Dq6kiEr09QUywEjCyBNlO5GCJB
LxKICIY8ikBwzT5UEmW3wYfOz4/00yTOO3kKX0F/kIA5avMP/Sm/xMoh0RM63Fjh
OYD9VfkIY699ZBYDKvrLoHnI0KIbwB5FLL+tA5Zlqgoi2ROnrOQ+IRvzrD0ruMtB
Zi0YaAzgoGtAK+k4kLLq79YOd+Ci6ST1tCpynN5/xNj8olh7behgz4l3UAJOJ4wI
T440U7p+0MaL2xdfuo2Ldt/4voL/dER2Hb+qCyXqg4Pm3PvU7OE0GrPtB6mq9q+S
3+8LDQ7eKxsTfd79qVQcmvP0IEUYWOWbnjytHen7bZ2rEZW/dOkv+9P/UNoNgJdl
0Oq/J1YdxoVl50bdiQfMIfQ39zn0UPydFsk4KjFmVcBCaDELsPMBZsbD7UgfM4Pk
nY5KCYVGuCuQuWSAI+JZLuuTl7cV65/qjz2dXRMThlcgV/sdcDd5/obzKZf05qYj
0sKZ7ySpED2k4CKe5XKOAMuCN4MY5MbAlIWhiW2pBmctT9Ju0Vm6xvKiwp+mozyn
qLaaQdeFhXaAxsxW2ZymVu/tCdlq+g1Ag4erJbcmuqratt7LluQZvu2+9vitNagA
uMaWmYbcTOcz46/Vst28BpiyQHZwYkLbFMZgNynaYqktxphtBlT5NJE0VppFR9IP
SPZGJoFvYM6l7pv+O8D8ibNu0HZRCk49bNk4TH+pND28ZBiewHVSJ/yCumIzwbGO
gJRQb0McogYGZOKH2reJr6LZFZxK8o/gZa1DjmpBodxX438gqUB4UULa6x/pnzIR
y1p4cnwPv+lja4u+xbKSCh19vFxgfu8TY9YT2RlfKkXXWQlp6mif6Ll2i1ExJ3xI
tQwf3K2JbyA2YFUhse3Zny2hd0AZh/MvGH1YRe0NuQfvcqoxgtL6gflKyzvc1xU3
5qyVLEBmjlK9eMh1GqDMFf8TiNmQNSBYZJbvoQeFVtNx5ZdmPBgHiM+OpvlQ1zMQ
/rtJ5O/JZ+0fJD+x/q7Z7K6hdn9safuqv9iki3sAYEKO1rdnq81BE+wToxuj828k
si/XGVe/77h6KQdMcu+ellvuqYae8JyiCX98LoOuNlL9UyupwTQjWtettsgxc/9X
ckbRqozh8G2BplZtxWCioIBfztciG4xa1Vvkrp4968SyLp44FPsCyAfBCbbxOujB
cAM3z29ZL3Zf15mcrFc3xE7xtpH9NPsJzUnB2yK8h7fGw0N6lF8D2b3Faz+B5kM/
pCXuwusw2/U4KIb5szJd1Z10gwE3l1/C0o71KsVxOtWGIGyNny/5acpnLmLQC3Od
e6db6tYdVQ/p1+nqjFqGkG4aYupHamT3b8QjraEJHCDJF/BLRwgSr2DO2ldgx2ID
8hdqAV2n64Hix2n9zPZlclO63tETcgcvgZbXY0GKq1j01wMfYvsKYVd5DmqUnupa
8qO/E8WGawSofvH4ibpAD9lSoI6QNrmKjH8fnKinoD7Y6pzMuygFKbjLa8/26aOG
R7rgVqu4ET/6EcvSfPLxbAl7dYjmczugDVw8ZdtIAeKPp5rtiONVEW05yL0nwTby
l6hUPt2zh9cKF9Fjcn2g1SA7wQg5pYhp3mw37pImEUZ19qSeyZmMW6OjqT8Xhj8d
243gbQXMhjfFVOLXj4aw3YzrTrkN/phxeRtSNMsaj4fkQBRROoeAGAdIPKnvlhlA
9z6XfhoIl0y1umwi76ip4Id5eRs9yp823scUowqhcyRCvzB1woLNAK7RVY8R3UFp
aG1ok3uFAW4bS/EnzquSsT5WzXNkP1KlHOcF+jguj5aML5vX1KNJ3j6FOKVnSPRv
zthijJeAZTCE9heLJPMi090Mgn6pl+FEGR25mP99NvkaI24FXmfAEi+6oIMAIBF7
FnKg7buDxkWE5vEpe3iHP/ZMnpofqvCzeuorss81W93Qe6xV/8MJ5gCzlnsyZFjc
PPfDqMoURoED3lhDizPBdiJNz7YY3/wwMpYTmPaIAPEq7FSMorWonrOoUkOxkTWN
GX4b+Esb9/dZpEKBIAw+o+gWspHWYS4pi/Ygs+wq/5tRxGhGfpr7MbbNKgovFiy5
JXBLbM5IeMquH1ju9Hs+ki0WJTltYaX8kfmRsWGPF8Uu845bVTJpriYyOzMN45rr
lJgFwlAH83CWvAGrijVtKCogX6F+utC+xK1mW45Z92NwN5/DxuhJJsWb9QFfCiW5
8VuIhayNmvBkv9LdT8dwkb2sCa0LdOEz1RvgYonLMvAugIpWTMN/saerZZNy+QOA
0PXiCBq/cCQQhH1bsjLpZB6ouGwgufvBk4nSxeEkp2cSs1FR/tYiPUwyZURQ1jyF
mJV4VRzXZRjRgPhEU6bFFX6mlAcZka0KYNSpR1MxnFb+ZBSOM7lFeQBUAcynz271
uNnMsU10MB4q40DoKCNysqJQNeXaRaSTGWKSHr/y2GQSn4j+FWYk2I/zmHwKpCh2
hV8vOaT8iQldH8vlHNnydlZovlNlWVHDJwhSvrI291EV/2u1Ooo1STaMKGWrZUh1
2RJX2OPVOWdoK9dZg6Ane243oJ285I5L2L8abjrQxqOydQG6B20oJU2oPJug4sMX
4lia0ZChWG56T5h2/I0iknAMGQycZ3hpZ/Hcm5hOpZIwihdQyYRw7BGTm3CF20oN
qfkwDlf9og3sIyTZ9CTSzMbsngSji5a8NVuwxIzeJoSfhETmbrXPEWRuqo9GFsnj
bdrkFitdI5DUcaWX0Qut9lKQ1aBydcWsCgu3YTzn5HqvazZlApFPNCMzUeuPyHg7
RSjJ6Yxk4KAf1Vll1gpuDBlzfminBbP8n+G9U/z68utomwz5MOQ202Z6pX9gMjAx
fCQPIIoY1SfuTn3jQATcu6qkYgiZVTVB3L+YCirmTB6Yi58lf/vQUlJnTMAoJhyo
ZSUolTBKw+ZZH+6bH/X/+tU6/e65EP7+oOx4MjFe05LVeeWBVBJMLeuk7VJop3SQ
8pTQxjLWBh4zEcAaW4erU0wBj72Mrg9YS24J76Ugg6YR7K6JoNukM1tBiwmVe7iH
kRWHCW79iN6eF+5wyw1szy6li+g2xn3tcybQzT+c4G+O0HPt02BbkZXmim5I01Ag
Q3Sd3VpCG6rxN864c5cPHlgw9rdVevv9K3mau/uYYjqbU86UtQ4d0/UVNHNI7Qhv
NvKQSmStSHwGpHoyTbU249M4PAhpaQnukXdSL7Kql04vn8TIRa4uGup7hO2MuB20
LKZENm5UDBRCtUOx+JjsVegx5FtTpvGJJjwjZvB5SAglr2M31ozXiIAZVttIjree
IrebiU7jYfmnpR2+jH+ZmBfdKCP0PdnXKHTVx9vVtn5JZqO1GsUV+LB83+GY1LSH
BY7W7bTKAwNnnsvT7SR+eUrqzHyUY1T96X2Nk1VoP0WldG4GaaGyxhzfaCQtF/pi
XaMC+/H5HaFRcsaV1AAMWMLVoY13RKcMERyR8jvyt9DfS1WH1E3zOuTXpCK0QKfA
bXE7GGqJviJ5Y2OUc2KbE2HJKvhjL3B1TlkANu9w8l3xt6pGYQWPDdA2gqtrYotx
p8AI+sEkHwQywMTyoPX5TQRtvia8A2TD9/XkPJy/0FkDzK8NK11keGczNlVpRZd8
R40mWuL/q7E8Q566jphTrGtO/aF+SGFIC/DOPU9UVV6jguE8JI8nBcdIE7i7d5J2
3lrhucU0H5Vif5tCp5AccMcmPiw02ePVXCNPcCe9VOi7hfTcc6M5FUuD29H7iuDm
DqtcH7Euhx6dF7mjFmM5lEXwe5SX64uKtazGKBj7I1n2N4NsG0NffT660s+hia9P
Akz1pzivWuQS6Y4o8PxRPWtT4GxVKfWpJUfHIgcsIPtW1ke3OMJu3OToi1sj/mxh
hvPmC8pW+2Zmo8auWJFfgm9wz3zGdhTPDvk+uFmgCxAeqd5WFCig13jJiT/b4P1c
vV4694EoIBGZnC+aTiu0NAQLYxiKnroebul52eyn1vs0fe+ApJ2jy3+P3EwUd3qJ
aYVSe2S/ulSYY7mvq4NADcqLQ27qynyT6Fg3dcBADaoMfnwl84gIRxn621W6bkvg
2ZUAFQoe1uFW8JkWWzfcBJX8+SiwaAWDIQv13EOSbH5MnIPfRDPqvrLhxHu9B4Qi
/9AOozFNr3KxLGyCukA3x/0Pa+7sZW+unpwS+Kvlw5L0KnDmKAgkIBpph03sedeC
CX48aF1ZWoGXTjuC16aJNnjlxQOzPydVuMbIEQ7tw2pcSC+IYDUy3Q/IZcYQTKrO
muFbeUSm9zjTuE2NHPhVNGTsKTsA1QSgOv/+LSUBEuKPLgsene9Ofa8MX6bBiFyG
VSL7ZgU6uBqmDrIFwZX+Xf3hUqGKyDL7hUvzEiUG3Sg1DCIvzzWX8/vZcgeZjDlu
I9Yy52W2XL17l21yLKJ2Z4Oh399iOKJihE2YLt0cfYxeYR3RQSl5JwZc33lm3r3L
mc6PVyHGti9Zq7CFcy++drTkB4qGig8F+Uso4NLBlZQlcS/sFKvMP+EeykINPQAa
XtJhUO03XZLZu0cZ/pwNV4uOoWyjHII6rQJHjcXhIR8sQCT7VGfYBwl/nYpYz9MN
I2UhPRi22ITDNFqa0niu/gCER11/1kRxgoTGZUTUdGjir4OKdSSI79sh3uo3afoc
bnDhmEgX/nwjKDb9MP46oiHWrRBO8qn0wCNKXxSF2kKYDDm+FdUOvJEWYIAB9827
rq1EjcSKJQ9CFe0dxMceHAjxj5nGsXQKmFTQj0gA1xYodudNHfrH6UeU9SsQRsa/
QQDaB4+JF+Ls7+4NpHwCgjTbSpGZlUE9dUKW+nI9nsilQIhdvE67NH7gRDf2629J
StOBjJ3yHM9cbAZeUydmUNue8wq8nkflOeOo7FSTcJLrpd6P+SildHucX5dWHAdq
5U5DuPiKiOADOQCoACYRl+tcJ2VD4GDFFS0RQjWz24l4kCRDddQtH/J6Awo6o/yS
i2p9gPPATPEEaJiz7/n6Vpw2SXUfkJ3ZQ9D/io4SpFnXQrqVH6/f/PN1NEYeWM9M
NeaB/ZqdqPreXVTclDl2WKJmae/WvdGSxXmBcqpUXyMtIt31avm24JlKvyVsMrB9
GANb4rjv/3vr+RYjuds7h1jjS72dVjqecEmRzlGshvrGisDXri9u8YRnEPeTnXmh
sdfziQ4Jrn/LefV3PLGQgEETrKDVeiG5j46O2uSmrX6ClwU134laj/OdcmeLEqRt
XkuzBiRBAAJzocdRFU6heOpOHfYR1eWlgHiZg6YzDr7Dzo2FadiHAgzFYH7Xb5QN
ptiDDRQW4MoGaH/P0XPAtYnNH6YNi/mNdP2CclNx1iWkjGBUMA7KQolBj+xSKCfz
h2sX/hs3VuKBCBUukyUo8a0vUtbDU3G9o/M5XlSGtBchYUubodarMHnEGsqeRLod
8t2Bx6WKzZGjWuHXQalRmK91v6SDOgxCMo1TVfvCoxUBZEQVXrjT4bK+JWACOUub
4YcO7SHbKk3BFBsX3YdQ7H+Bvx3K4lFYbSrCaKpU6vp8OBLftWExu1bVetC5z7bb
2nCEyiBIXdECegd7s9sV8v9S43pCMqfnl7pY3+vpq6Re6EGg3+NtchM89PwTTsav
6n25jd2rMKvvcZc7OLN4oi/tqW/aywoerIMlrOh/AeoHHHcAzADzi8wfjsFlEROe
1/SinqbxSyB8geHrS3O4PQXl1fYU+VIHXoHY5DoP2soI9oOJllnu5dqfROdWh0Mh
YWq0dUvAStqAwhwNO3NXpeL1DiCMEbDaGtJ0JBieGJfzKFmvyhqN67BIfTkkIeyH
JszSbZZV3F3n/6N/+YVfFHOLlsrC6/oH/qBzHPgDtiQ7uCntowfi/aIMl4xMRoxL
5twsI8PLD1vhjfQW80BzLFlXA9zlcCO76H2jTJ0XXqxGyqHJdK5DTjJ47AftKOAH
k/xw4JU9+sMhK3tIa9YErw1PvrZqJH0bcJCqvECCHp3yIqoSlKOaqmmDDHek+urB
UPxobXioUjjAwfAxx4tydNc/+TxDwXTN64jg45Hd8dtEseCSzp1IogivwBijlQn4
5uxdcdDLdActyWis6Bgl1e4YV0PvPQVAKOOZHlBezz9L04CRUCYoYRrkGhYsotHF
T1QWj6tL7VLn5yXQJ9Ovu6I6tWMvivNctB8UgLzbHhcmgrXMxX1cV92ehmFPBi4X
VAeUoVRVY/JgCz/0Vv5omuVu4lhMBnMY0gAX/MWt3Y8dpTqhLxM+51Dy7vXt831Q
5CB0/8d2IZ/+khnWLslsB6WMm1H8geTV/+nQ8OXxku6c65cA1blfiKzoO5R7bLea
/dlqtrCL4zlb4yuu5qB4xCukcoHlc1mLisPZJoaim1WtjZUVch+K4VdvivVdMmcD
A7EFg9edYAQjriLJJxjT/Gp6cfkgiwALt/XbJI6gN6bPjIo2kF2HsLKQ20MZoYZ3
vtUhY6bitDnyTXrkDLBAuo7qf3Ra/LblEdWsr2Ejuo0eQyrVEG4+jZGzKPWQq2jS
X8FxHInRz7gsri7NFk0Ny8QgGDyUUOkvwI9wVnDE8Z/mW+d5rlZTLT5PVTPPQTLM
C6S+S0YN63YSgoDSW39Cb3X4GDOEPnRr7MdTG8bfzxszgreJlqpWp742s3QVzuL2
vueTmdxdYl3vs3ytUX+Uk+RZ9gVvSS0kD39WBwPARkdkwuXWRJnAmkRdiunw2kI8
5xsgXAvvLBnZq3kDEvcFv0FVD8ZeSTmAsvUWYLBM+r/H2dhe91QOFMCjDstWXtg9
0DtpIcug/t7mJjmutCovnJ8QrXaZKJvpAmqpOe3VVisEMATPrAmCAdBPUezRJ44T
0lZDe53UHwYqJpTVop8KY0zzI47amHKIm0WawJ4OQC38DveBKVpznjhIfHQi34nI
czqA84MBZbz51EEGWoewwMjYJQ3JcUOI2lacAM4/1MPHLj9zVRTkfrXdb/74IUgP
Q03atlRZLMr3kYpLFFA6aM7wLnXIUkQ+2hqYsmgPBIqn0syESKbdiXoYQ8re/OLB
PJRXLyn/PgTWHP1vptLKGfKp3KDS/YZDlLs5DHOGIWzF+W4mUaHftw7Xr5Qes5aC
cagGTnIIFhXlSSVi4plKd0RKpDU8DkHY9xqqQrbw857IRD+h9hju4lmZci8XT+OI
fU2z6ggiGwJdHiPCeIxcvXa0WH3htmXh54A/SBgj2s82q/hnog+WNWa9oyK9EIki
JwrA9o5Jve9Aoz9n0NZ0Yhc+KJmAJZvbeTMfmrLwCbGugAAympDXHYP+5ZyPll1H
Sgvz5BwolGoJsyWpbgm8+B8/dcql4yyI09D5wzauBlY2injPymDinyfU5brxucDA
UDqRvXR4tP7Oc4VmRKUVUAB4VBkVt6tAlmouEIBoJEeotNsYsblZrV4QfYTsmFtk
H3xw6MSGJx0NhlTJwCS38WpDxjNOvATC0T3MStocgd5eDjmHvNytslwRFPJ6TnYs
WhiSYvtXSgV6kmeMHvE2VUc5WiYkE014jLHkBGE+rOwMWF7NLWeBCN3WEGSFy5Nc
dE16Ag22Wgc3LDvCXbLejoZtRUAF+JQQ4COsNy/B5zNksdOzTOUQ06DbOnvf5mgU
04D4R23sfS95eRkyhr/UAKBv4IpTBm2IupHnoSLwyivXUllCNihL6thIVHrP18kf
j0NCROMBGSmEDUe0c1yOjDEp5lYbBLVjrf7T48Svj5TfILw39Q7QWNkLV2NpM7JN
F69h4QT/J9xwrC+Y0p0vTctfKtTKou00yVkTVuy8ySrsM6pdCKCKnwo6KRljQpK2
O+XN0qYWLzt6Z+GD3sDfGk/SYwjfQ/aAyweS/tC80/D7pHnnwS+KoTDxbyq+aFfG
MFglxDEAWmHOJuMGlEtG9akrYPWTK4Uzhgy2GVBfG/ACBydGIZe/lvHdpcOOXqGl
hQHfJOs9+LyWPAsrv8/3Kxzu1JyJFhL3uYDn8qrW5pypzAhksXws8HZN+Pz40qFr
fu3BWpVxPJuVwQ6H3XVVNGdFdnSwScGulRtgD8FY1SRil0pQB+s9LLFyhOWmLNGB
x5VIKIshIkFHcrFtcfxgkQ==
`pragma protect end_protected
