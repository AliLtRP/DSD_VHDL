// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b0ZUVNwoa/6Eq7Tu2XfU3VDlhb+97+V0jwdYAWOqDFWw/OaH/An+Mpxxbjf5UT7p
PXK7kMVkWQIv+hYk6tIEiMRNT6BOdjWCaOOwvU8KZWQq8OAlslN09cvFraw51FSy
nwcbVZcnHOjMYrk/GpH8mS5QRkZVN65IEhzDi5dAEzI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
FgX+jaoy0Kc3YIAXtV1C1kgtSOu+sDBba1NSwdyRt9NwcDgM7sf70GC/sCxuMhlP
KcgBSjSgW1bT6JqDTh7ygSIo44kgCIs8fnQfPDezGDCp3fmtFB+luP9RCHo5qzoJ
lCzThihLFS4r11wBfpX9WDzuC8Quz3XW+D6Hq+lghPT5Lb0GIqKrbhhg4tNtHi47
T/nk+GE6FWjCEgGtx23r1JSVBTDVek8mv5eOJRIb3e6CqCcb/F3Xlvgax5ljtWap
FWlZUKmrkM3sy8uAMZONWpaAVTmS5tlZtiGbAWQUNEJwI5EvIRbi3jEzIyJlyfSI
u/qWcwlSYBlu9rt7q4bpbo//l563LV6yt2zEJppRN9D4+fkEfge+3ycuXDA+9y88
9SXoafBNMxkNU7JR0ORlHGbUcqypaaaii9QY7yZRO3dTsp+aRHn23+Kd8VLWOFDT
OFXsQkbgTZZumwpG3+F59J/7jbz3zLWDYY8thoqPoG5pvh9NBeowd+wQctXedr8c
lpwkjgVthIn8mjS/4Qo5lwPfSmq1xjL9N0ZvgJGjWeuJvnapu6RH1e0duN5t7pEF
N73XGYSbMSkpLulSynoHmwX4Hkdwg7LDGqhoKikH0FAFKEfaZU7FWejPmE7K3c3/
HpOa+TD58iY1U3TRzoql7pw6er35vEzzo0COQEXYEQhUe2UjLg5MfWCiCtO8lIop
B8EcRAmkqoRyu6RQAG0koAWr6vEQKy4ptEhkFUfEf9H1SGyzLIFln5CfnA2/Dz2s
kn3/OVjA8RZvzG4GoQJf5fDGGTBd20a7sVBWmUvo/fu8MNRqvr19zSh4nybJOdPN
j304HUJZejJBTcGIi7Mlet78arSNw2V/Jlpm5VwBj50NeqjsklnDedw37K2rvw49
rc/dbQj3toGtBh4JXvv4bB3la58nlambofGyL7HBvQIcovci/Gg8tKdOw4wYVZN/
pXjhSztFMQHpKjdSBmtfxMUzD7YpWlyI5SnYHRTlle6na/RNCw5ExkhAjX8N60sV
3mmLcjoImYAtqpcaBAGE6Q6YHD0+pl3RfEb+xO/0j9h2Z9J6ZxhQGlHH3tKhSJMn
uL9pIkPDcF3J5zTdUh2HYa8rZQZP8dkAudhtvThfoff7mqO495X2+MndvkgzwUuC
PA2LSrzfoefwTbej6T0pW6mlHBYPaV3m2i459n/+ETql76JrUrWsMV8l7IjSR8+k
CMcNhGmfGddHUGuqbtCG6rvwb8ReD2iMMSnIVvCDP/+w2BtHbkByPMhJr8O0hVa3
KSDdGq6+o0sG1uNbyi7B4gsnm4Fo2LjvtijC+xzQOPDwd2DEl3jwMHeoLxmI+1My
p/cFyblucv/O/sD52K+U6WR9tx/2s2e+N5Phw9UfqvyRpJfBRC0IT0iXuszadbJP
eqy67PKqY++cwj5Wb1psa/jKJuqNLL2v2OwG8k8pIVB1kg2h9yKJbnnklKIqK9dp
p6ofvcxfHL74bGPjOU6uay7wxMUbidGsT+ss/omu50pBnoDGRX9mxVCs0ABOI8JY
xPrKf8fFFw7W3POXyDKp/chdIvKuTFCHbqTJFIH/hMGHMrdWlP/YmXXZfv18Il8R
u/L2NjVYPxkC72iKa0W8NxWQl0+lrhkgtNQsZVMnwU84MXijqcHmwr9yQiFsHXhz
AqRSaeO8BLHt30czvIr/DlJxrDSO/Sv0OuF1uDP6dfm8loywa2B8vSCK4QrjdYaO
I8FVjsByagMcCQuW/46J8jK1ZDrqF0Z7RKnJm6CW1r6zaAINvgUraMGUrYCEKA8a
UGn5+Cn/YMcwQ/r08oUwn0e+7gBKQEbtXn+vJHdN3NEWNavX5jYJofx+QKUb73KD
CB60WCblRGp2KtmDUiU/QELOCNVZRjl+mwqIxRQ0MN06le7cEh2UMgfoqScaM2WC
8uuPAg5fWr5zmWWDwVDrOciuFctc839yOJwxtGVbPIXymrtiIYFSNCHnusQfgiHt
RdqdXeglTdFpihsQ7prO8fhHiKa4j3n46NsyqPFi+D8jay1GrzWHIndJRxwKYjsM
lM/UKTib1ohAz13b8lMdEcvnTWx027Ki5qiXEteicVzvV4UbAkYsQdIa/mxyliMz
YZmRbw2MqiRtUWrGLur5OUbBPmrSDrQpjznKVANe0He5O01svtPWONJmynezSc9U
pT4NfCMLbGvkpOWQkOi9Y8pvTzMk2FJz1KXEyobSo8+m0AGDiOt5wulc7DDSt8H3
mvYpt3/xGru6nfGH6V2e5U30wDKBIWb+6FtRlPdGb23qsZvrGpU8xYa1rVVyvV5Z
qWHPTCvRP7WmopcXwpkfTK/i5FOofVt9DNejfYZeYHFDZgYR5Ta36NfxMFjNUH5J
J2JxObukbx7oDfaCoyFLWkZVcCUEMaGUfEw9bheIvtwQy3lxDZpNzeeCUtFOlUrI
6T0TvFb8aj1o8Ej/GsOnrCxnzilAB9zXletAJRFHIpaSLe7bs1RzQC6iHdx11NhR
ZV4o1kn+25wWtTM3ToFODzVowp9cYRBOnZIlUd52OL7YR/JhIo+AvFXXcmfoxWeO
EBger/KBQoQZYHWN75gFgXiybR/jh7FP/mLnUM+f+FvQ64RQdDcn5UbIBbr0yl1+
56rSbuSJn29utlskyGQwKPDJQTprJ30KSAGoiaTz1Tf7SZaEDG3LoUM2rhOnBUXI
ioqqPenKamcHg9MXfjC/rsiq3l+rDT1VcX639/mxNci9USih77XfmXiuJwp0GkP3
BdqHXDdYiYslVbzUZWfhRWxl+zbS+G1BdwuIcd9s/Hh7VuUArBkf9Ge6IpPWSzid
8JwaUIa0XXURfiTd8pruY6+Oa0KkRQa6tvIIj+RBNmRFTpD1t0yTXouEHG/pjBur
h8TRqHsojyvqxr4XtrS/MLxFyWf3owov54r14fN6Jyovnwqs8jNejw/ot3dtKBnv
/bVwZP/oWEymC10s6Eh3Clp3vWNHRDDETSZyNjj+7aGVdYvEA5SWZFfHhFNjCc3i
DQaPBWDH5BhU+FeonjI9cYyZ4Qk8P/tCe4mqfcaEm9JaLrghWB/nGi4xGXPHs4NI
Unnrb+85OyF71IRzUp5Zyhn9jG0YgTfhzE+CUohesHFWdN+o2XiGAhHhmlJo8asi
5KabNkNNkXSgxy+Op9vEwyNDMBpVywMvh6xFBwX5HwMnDDVrqAD1ekRCtaqk/Ed9
AixiK0A+y3xRcCQMMFSjIrvtcR/4Gn9Qkfpa/Kc0b12iLkC7yFqdtMrdi4FguapT
`pragma protect end_protected
