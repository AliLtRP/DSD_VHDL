// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kx8ycYbBrx2U7gERMnmdw2AiOqiKyjGr7K6nPVMj9pLQJ/neJJRM5M6nmvs0RPu7
89mMXcmtgYw5OLZM6q4B0aYMxw6IbwlAVB7l7s5ERgir4+2e1GTF0D2kdHufzX+2
Nwx0+UoWaxh+HUWgAF7SpuIrkjEZ5U+tBMK8XylF9go=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48880)
yHApA3v/lg5uOc76KLlV/hqHCxvbXH747U3Jgn545IjlpcG0ppgoI2qRRc9pRcnz
zTJy2S9RnJhqWtMjkaxn4PUWeEdpxKKo2O4mYzKDSFTffgrvVzx89jzGFBnz+cAV
ddKd2dAorIXL/bTaT1kqCREY9HMYB+bIucemBWu83wmPr01rWvuRqzJtRwj/drLc
ZGwWOmoCFbcuoCNTbi+I7apyEN5Icoz92VXOSsS1/tL8ZwzUL2ijhNmLyDy3M2iv
Y8TxdReiYo1X2YThf43eC7wbwVoH2ng37dn4cm2t8H9nX1R4Oj/D5UNKbYiSHdtg
1VwbGO55Ozs3Ed3cvx49GhkyHCc39KAFCPhuRiTGBTcOafK2m/kRfx9ekINVnYSW
WyqzzVd0oNa4BRmgZaATU7tkEKgCYghGT4ImGxNHoWKE9q2U6av3J5k618BupKhY
txk/tv6Zbwl6wuxJU7fyksvz6R+4o+61T7rzsA3E1ocoiTvH7YYq6W6cLjkS9WQg
ZAhMSkjslv7XVL+NIqmF3HUpEPbTFyizxh/MQX5dxpRcIhZuvKckvUbKrpx4TQFP
djsux8cP8eH0m/W19IvKI2ZMtyW3Ytr6a7JEwGRMRaMRq56oucWx3+omYnJy49nX
EhxCfCuJNeDeQwyCQMSGbL8Jez0wONJ2/ujpLcxfZSS3M45MruSKtk6j4mpDvunh
V2A8kzooNxSp2hhWjHdJdwuTJz7kszyIMKZNSwCad7p/aKIPTyunLP4s7STtUsjI
470h0dgS/TTPld1irUhaZB0lH0vx+K3aAnijqxFNn/QK2jqG5cJvP2qTEV2WpIoe
di7rvCppTVLRVZB/oujZmxmNCsqUE9ZkYk9coZw7jGwQ5QVxFJZxK7BRPzXYOrKH
tWXbRiSoXokhbiCF+tXBunzxupAWubYndD90AZAkNrnO+FH4OzZzFDZvwXVXgiiP
kk2iCuaWb35LOa/1osqORVpnLQwgk+4aY3xzgYNMSIWMYeBcuDPm4/mJe2t9EW+o
2+mfzyVif24nY4locDmK/LfCjrV2dnuAE5sRADVzh293rIH34jOJDfMDSu6cOQdO
6VL3RwC5QQ57+bP/IO7TZqudzg9GeQxgzkrm02EUl6O4OfBFtfd3tN7ER3OekRHC
O/qEBVwKAz74kLlNq22d7zFgRGA+DhADwxPtMw1oy7/jRQLXK/+P5wToX4QuxJLp
IeEgDvl81ofzK1qdWO4BcoKbL4KYbFMOxR7QolDQQe7NMWJjK4HL+EwQTv2g1e9y
afOXN9qycFYM6nCGIyvCWMF0kCuNBFaOVFL6gy9wrEnHEXpe8bhwTc4P+YO2ZrRG
TIAR3aiuyQF5AriYpA8zVowc87ZWzAZ7aYoRe376Ypde+5sb96LO50WzB6Bu81rm
kXrNa6n1wPojBsJjML649K4/fcqA3rKiB4AbN6BF/02UcbvXmGd5M8FnWXMlXljy
OiywXMN4gHqze/ee8qnseD4tQNN5Yu/2srQQO/w40CigWfI2Rg9jdfLpAJ2QByx2
gRQlgxi1XvgSWklrnFOR8ZYyWid8H/5d0BpFd0dr0FSXfUJPGl1GJeOllh2pysB9
WXS7czgRBDvCoL2pLNCr5PS9TAq+FiyBVA3ylgElO6fnRxZYyf2cPcJjLyYYX+Iu
43nKE0cCW/XItDbvVUdvJPJSyK/xO35ooeRHnrB0ixcoXK3cci1Kz1NkPVje9IF2
NYCFb/h6X2guhK8/P5wOkIe9qNFpzFp6Tenm4nTmHSuy6b6iOnHZYCcaBen6PmA8
S3ctXkSiJ4h65SclhOYkUNC5DW2JPsQSaOTUcI+T5noT0zoZBczAsFDIewr7Zr8B
+JGpV87iMassDWKyDgBm0bzxvxHCqpQlcBw3+5i1/ofDApjcqQ81RaHIW7lFKcAH
9GRhZ/M3FutxhGe9M+QweG9mr2H3vcpq6V+9ZmlzaZfQBtQu1zXYZu4+H7YOoFVN
Nwruh6O0hXU7/6IlTrMnAQgoWpqeelGNA03zW7djpTrSoHpWCnxGnjZgIn2SAT0H
+tNwC4bVyBRpuhzkT1GeB31pvudvogcyocQMtqHPLoZJcqS+Z07+RNThLy8VCAh9
yaXbgHInfo9z/jx+N0uTuxHG6HjH6gdNtitzgEQvtyvKTt1gxrJ5bRKfvydvEOf+
FSSphajF2YXs+UK+6unqY/k5OAVFl0TsEd+mteJg/16mtqJEGfM4c7SsksZrbkC6
Fk9IQqzzFaUvSC2mqcn9vckdNZ79d0f342VSssp35IXbJcdnFftM/KNVxxj3FRJf
R8IiaTBocpr60JiOnFqI/NrXMLUC+JqebmBcGSFn/ZewCtQH8Vy4CjtZ3Mlpi3I5
7Ksqv5wD+jW7m3po8X+h2tzv2N8azTplKQIYpmgxIKe8EF0Zo6pp0V4QXB6OFMHf
TFMY3SHs7HBC6ZuGrIhPd0H2Wjx/++vLlaOFPbXK6NZ8WnUWleqTRoA5Unt2Q3kt
nCNREcUlczHO0cHWrs3eeol68zCuPf5rcWytXn5fbkQVxUd0ICbACmC91F2IRFai
qcCEv7CyriGbVt9T7UH1pGtTuIlGGhT6lcEC9/+ZI6uSH9AeUs7eMN92bN/cbxty
W/q/iJ6VFohFOQ8o00ejQKCXHR9xpc3pLyueIv7wzbr2iNQC5dLhNUKw5zuVg7Fm
NBfJ+KHbqQigDsa9tssQ6VZdRnQIRYpacJiWY4Qu3pzgPKiDIUJP/ORzgtRhsTjd
Gf3+YFT1GBOaLvPuMHC5aL6tlPbL4qMqsJqvP/IjEsU3nnIV6csyKr4IzkvWow5e
S8j39bnSzmPhvVbkBuDPhbwjcttvgLEEbkKpHYBVrEST4iIUCM/p3Toc1bg9tL5j
wsHR0bd+/+EQ7aUnhRPESfXJ57Ncrm+nnAUj2Go9Emi3Tt0LH0z+dHLCuLhhrBhF
IwqM2iWqpXuTBT2dzz3X1kvyQn5ib3auO0ylsDPt6dAsXFkdjB605/5+FnFxlNAI
kEj2buJMC9dah/XLIGa78D+j919QeTyCfblXNe+ez2DSnJFuBu2pnCYBghCrOMK1
cDKS9dHUKCQD+CP3K7b/Ul0UYPePeFZggCQbkQeJfVhttCn2iUvNxwTDZa3mkH4I
guywxRqYPPIvANfrZ1qlOCtsaLqFKFhoM4d/TJsK6aSvzjYT40G9D8Hp4Z5Ebnq6
PP3SHLaXAyKXxWREXfvFxsSs1YKMalO8icJ5NH3kxx3Mfdt5HbyaI0nEzpbWVLdH
d4Nh5drEGfuyfX1yYDnqS7iAwRm3rd+lj5UkCBZD1SDa9wp3iLFzsEfE1f9r/p+P
uWmKiroulGWrEMO4YCGN/bTFCGlw2vuiro1cjMoEdOanzT+B5SWMoumGPYOtGDOS
4d5GPZNmA4nU9yJCvombXN4fX8zBn7K6eNRKR+M5Lar+Um8vLUnycOLbkWKhk/Ri
DCckMjZn9jm7CeKKB16FFK/SIFQRf+plTg8n66N8Ed7+x6rNCvGCJHlYXFRHc3In
1qZIHv8+sdkWeyrOMnk0oJfWlITWG7g8LIomONER2ccAk6kqnXAIpV7mCSFK+pFG
vaS8wDNk0eJnpGu76YgSJyJeREkN8mwknLkqEmZEs1Ki8Y5eDOd+haYs/3KNAA9R
uWWnlyApjteFKSIUXHZfdox7tcgzu72/3sqYWl9rd0zGigzE/ZOn6rHRY551dHAg
QiMbeUN87s40heDCh4tI3PKo79iAWtspmwrpff2f28URspShkc/D7EHgPKSg9zZl
XeHYq6u2b8n/ui9Z6aQ1AK039SS/NcqHc6AM+UFyUnpSq2MD5z8YTGZ3ttOT78nJ
cFGaUNLyNujXQzeJXj+c9LmZeL1/iLCk59r20J8wQ10VFHJ4cb6Ba2BSqdoZD1DM
ETXq4KIO82oBwTk6rUS+Ppv7QROvUwiIUAixeRBUblIX7FVYRfkkPog6y0SJ1lwW
jPT3NmwpslaAJhPI4PkYCWogNeFQOv+SOcZ3zrhsoTROoRKcWp1MAqu35v8NY988
QYVeiqwpwqccN2VMh1VBy2S/jH2xdZhp5EvlZxXclHg78DcuuoF9YR/wOatfsK55
Z47H3LzGluLgPc6PmivHpV78EpERbYOh4VKjnSXlsyU5V1X/NBTxK1Es6HoUL1bA
X4fbdOSq3pS34wxs0vroWkg8SQJnquNj/f7obWhjOamrt8Lnj50sxqEUT+SobRnX
ZOfMcFFsNR29Ud1QMHUQloSxSCrJa4ZNjC3UftDyCNOQ8Cr3bgV47CwZb+8PDQum
AHMIbhstiw0pelFhr7decNAuoZXo0OQlD0zZJwZFBRbYuYoz+Kl3pWh13hzyokT2
IsGrAqykExcFN2KHDb8lLaSoY1u+yal7MqyUpMG+d2lOaoSdiHedO6bMfv6iLKJT
0ksCWeUt9AdgTUpnLu9XEQPdQED8/p4wpiIXrIpNAliCKb9e/8zF9h5YWEEvaoyF
vwH85cQXy3tR5Fd9AhVz2+uiw5tPoHXC+6Woy1ccVO7ng+80RSrLdOY1a/QylDkR
cPW6rcA3D7AT5Tht2maFA7lFczjM/I0gRlZv5c5vyXTzPqnMivoYJEGtEXK5xCsv
/tlb9pIxMooYsLamrznPgR7wjnXSo5+emKVKe1KUHVgl6MzQcCUPNQmmvw8O2nLH
UXFrJYDo8gLrhd3xCUQextvIbtARfOrU1nvEsRa4RfhuX0h9MT0hIx3eNpr+9DOl
BAM3/8zlJdzubQDDefWdL9Rt0xrca3xZnF+fVSurOfDMTPjk1epgFfvtmuOPVaG5
/cLeZrg02k+74HLrCwGr37IaorGiUiwonrHypwpKm35pSSDXa7VclMoo5+9kE3Bu
hjve4eXokfR9MPdI4uDvGS2wpMOBfmbiS53UxHTahHfS0il2QmA2FtLIUl6xRJ2m
tPTS1rhWwwQNzkopjSgSzrkXvxrv+UBbY3/UInob3EbN75hfqA9ft3OIyaVtjn2h
fpE7GSeETo+3eSx+cwxQzFTSXENJ57k81mBUrVqY8iTkG5DRqkSmvLviggfGtMr8
+9LtGOIOayE7uTZ9eEAlqf9ASeiG2D6BrCZJe6X7i77koIdr7DrRb/1mWnszh7tE
euyX3Ske00vQjWwx4+2kfJsx8+xY4yu1FB0oE2E8Otae6wh2t6UsodRgxX610FiV
CyqDiKdOJiHlqbjs9XNgtFvsyC5dI4jFMsVXjyUsH+mZlKoM1Hw3spOW1cYAYGCj
+faf/oryxP7LAiiOEtAQ4pUfaCN2KxjaEDMacTlJX6Fa0qgIb4Iw7lbGtzNjp/yQ
KsshHkxnH6TQuyBIZRcPlaCwsmwf3RSajuBfAFEwkVL695V8vDtJzveY+EtOYqki
nnr3Rbuh+d80mLJx4c5x6s9a8Lg6/j3XeMQODJXvHPGvMGFUsTnzbhgdi517UiDI
vS4wZ82wbFPvYH+6k+f99IBSPKX5xokRXRzK6v+0pTmnFQdTcmfhSZ68AJEbQ8A9
5S9nCEEh7Kzq0EcgFDOI2p9LcBL8kXiJNchdpo0lByMT7srKej0HA88Kg5PWjm2s
jpL7wucU2fZA2dZrk+v1+u99smIiPU9XOD/gF6HNsRMpCI/wogiOsKOe6zrbFXVM
h/WuXu5KlknSHP0F4XDD5pdcKhYT/EdraAkjXzv3/W/KGAVv67rcIBBJLvejIOjw
n7y8reAb7WPlpbwpDafTp6ZWbDRzMrpE/rVDzWq1K58D3Mx7oaqpJpvZ3rayXut0
JaOhmL8+rh3E85kXZcWkInK21Nmw7yQFuhVGNg06+1AnApudcgBUN+VLYafLroby
DGO/pmiJC7765pkOc372jdEFwQXiYoH2tT6bOyxumbDBGrSpME+TVQGSnzQuwsWx
g6iRDhOziTYjpT0Tr/23wGWT1JL3ppztRg3ve2eMzuo03M34sK6BkJ/Vy6gMO91C
J3QVtx+BbwoKcDjnS48JAfd2haG5XhczYtUJvvWWg7RHdhbddzI3DcTsxjMrNDPo
o1DbTW8J83G/qDWMRoZ3id29vry6hxeawFgeSQVYMFHCqMC1AfJaUoXSDq0g65O1
joJpF24q0UuXgVlsHzhU6vhdrrYw1xGw10fSZNsHJSp7i1OAyylF0PZyxFjkHy7c
xdFqL/1iTnmHPmw163+399u6S/AZIhidkm8M4ljWPbtM8aKjn9jIoMh9UIWZXafV
MScdgH1SHdeYHZiotQxXPlZvHYwOwg67molzso8ZO02VFdo1J/FltwJ5zFZd9DZi
DZIkd//wty0J2cwU4L/2G0t7bwge3kXCnQLIoUeTO5vNnYPwi6WaHqf+t5yVE1qr
i6wL9+Zns7uZBbHYb86ZTSb4MXmD4fCjV//6gLej/irqkSkD9BIoZvVxj1rTM+D9
oR/e96rU5/JOs22ok8/lK17gULVOnYeYQEgoKx9v4s0Cp0hLlyJrFzz3B5/fDuDB
jXXJsJmA7VZ4quBCso/sr0EfRj1nEHGQWRoUTAnB/h6JJiZTMOXZQxYJPpOZxDfm
SOXdQ0Bs6yVGbKPjhhMpOZ1HVZJ2PjbESp5ol5F2eLuDJDp6XT7h/9oQg5he3l+l
7QiVKizhw5Ammy4RKWS0KtIK2Lh99fHU8sqmWzfOsHNlxEiUakdDjpoGrJ0xWc4f
B0abQQUZMtck41wXEaB2IXtFuhochpMnJD1cO2MpVxLVaIUsGojlg8Oy2pb0Rf9/
Ev6ajwHnJIP3iiI88FDsUxJchRllaTVwkuBDokLHFr60HT+eICcXXYrAvTqADIb4
2yGk2NxlelkKL1NybMPrF7erc3ieyeB7TdbMZp5ltp7ALDVzjvV6CozSVDJOYBDM
3Fqfq9qOf0XUaBjqdQ0KAu6zAOnElcknXCJMlWTZghipKzLzhwidChk9mqmUcxwV
EC7RPCHXP6hrTe+CyCXB6dpxsaaFw4bAHBAxRnAlCSNCN1qSBuCQklJNafMWntgK
xoxA9cvFapeGIADdrZEc7OsYkb2s9Dx3IKh0ScMWcV5jI78n2CRBlCgb9cbR2e5r
YceG40jZVoAWYJa2qq3juTlnFg0/3vUdfHoA6mLG17A9ZUql0AOXk22+QSbR7oPX
ZWZxRuF9vyg3HZUAQO+MGVWqfNjQ0F1iz8jog11Dqxc2VXh5KdAEvWjqcn3Vmq+o
cXkWyaXcMaYry3/9cw90uMFyZW7MOObXf0CQ/KFQ6mD+Z7R4VuDe2fgOUSNuTa7K
AKOlZuZx531+LcxEd1nU0dOCs6HYXGVWRxpUl6fKbkgq26Rf0nbp5/eRhcHOa+H5
oQJsjnozSHtMcWa+E+T6qTXPTzv1rrkWMkCb3r1MWt0X2r88eRZs/9OUbxA55Xck
YUw0emh57QLfn7RoZuTYViqrIbZwRGO+1wQawDt0tflHI5+/qgxtpGmWsuiP8z0y
7wTY5Rko6BZ498id5lZ8GMkurirYIVgAEaeyYtJ5ZFkgvQFeDLPyPx5DgVVf0bqw
Wnd1q4gafkE/whnJvzaFV485Bd8mjKXrweS4f0DGr7AvAggpK2aTXFaf1fWTEkmW
7DBzhmnS3sXqtjrWTqjYha58QREbXl0jBSQk1sGLEYAsOacrffUTUMHp74Ozf21E
p4U4moJviyyXe4E9SMVAcIKg+P8rCLq4fDz2x40O0tmPq+zdw+FlA6dKCaL+or0U
DcB+J+zAZCAf0sLkCuKq3t8XCQyKJiJWrvzUiIs+T6ZISL4n+e2am3aUrjdWpLEN
ltMM87L8+a8FE/QmejfVvFV3PtldKti3qIhKNKQBtl7QzJeiJlz0CMwE8dLruPRJ
aA0rMufZAKE3iEcY+AqCCC9mN6Ola7PpY1MytzrnNO1/bOKQcSiu5iIhfxG6rr8k
uZgULo1tFfs4kepyUrihreo9kwu4nfN8wiNy7Q99dBbHzLZdS6uqPEeislm5XbEj
n7ApnBH4VrGWcGsEwcrhG6x0+XKO/kCyg6GBSdqn/EPtVSGDfV0hT5j8aq0o5htP
U2wi2vER+nhGTMwEoZ18cIwZGnZAYBgoEog+BmH0NZLeVAfevDscamoEokFlJC8E
nvClBYs2a1Qvk7mnETAe/cil9ddUl0oT2ApfTbxKMwvsio4dkdh4NwBF8Cl3Y7+m
bJXIoOdmGCTS3TnPp2LCiRMnq/Wy5R9gY55Qt37mv2cUcgjEPGImskS0pr39mjPQ
KuaJb9T2ght0GMHJH2jw637JfQMt0QYIFAykB7F2XdkSQhGXA+waKCV+tNbPoc/o
no1I0l2NmDJ1fDmS+oAfe29qJ2cZohV35XLrNNNWfLL++CacuVBj7xdxuI821MYW
oPItmNx06Hu6RuVaOhXSM7otli8cSDREQL9BMRuPGC6GiOkF7tTjlyAxtvcG9l+5
nkhx2WjkRUFbVhJRsVuRsfIyXebbXqTF+aayjRieRd8wsNXKiItkVzWWBwJuJybs
5LhMGUJaPvmpYrjZ44NMlkYM6OKngJbM3P2E8PZl44pRvija8yIZzLi0LcBr92+0
3EWmksYE/sGoIp9BNtUXzAWkhI+ZAfq5hz9b8FEZn4PbYeG3SpTYYXPLgrmkAsrj
sScEhQRRIoWueIYtbt3D9BGMNuXppIXkbjP2f+QqYpVKVD9sEpF3pVhjzxe5m2aq
PdOwcC6+ECL857rcIecDElAtD962FTSj+50PqgKrRhyuIde1O2ZqSwjm5VLmnR4M
KiWdO381hTMpgd9P4joRd7xSFSVwTFYoKX0/1EohkQLG646kxJjpRbWkMdcGc9nl
so6eO3l8pXPbwqMcnyzz73RF4JhKB0ll8bptTGWe5y6TUiLV6lVfw76PrbMMRac5
yua1Zxmh7JRQPb49bnyh/bL4fHdTY26pcBSjK+d6ULnhbhxkKpI7ZT/Ww0QYsdIy
DAT5OEjWfzYz+F3JPeq5B5VkMjtrxgAY+AbZ3p0QDmQNbY3wqDSSaXSHFWpiHz2P
kxdOmyuxod7cpALodKXxW54OoE1GLxmkUVW8CPXAsTNlvH3a1ZbpKZ47r8Y3noAM
Qvjm5Nci3cHXzI+PkRwHW4eQxt4l6OZD5Xdsx3/T0fEbtrZCf8CxoH29sSr6UhUS
6i4SatDb5pTWDc4fmObLTG9OxpkoJOCpPrWHJBEE4ptLRWxseYLLL5Dne+ZZU98r
DwJbhsdzRNbBl2Egdp6wHGoVzbfsFvcWdPPVYSQGA607owP8T0/uij8TcVnmW4ZW
MIMp9tsal+UZNigNVRH8vpOH9j+Orb+iDMyGQS9J52DmINLWQ0o+7kT4iIVdoXDF
GHpkc11QIdLgHKKKNnVZjRjZ2Wn3QS3VRWNzM7bSb6/qE45T8poSMhIu3Ztn1EV8
MGqZPaMULKQIyunaNcTukGtIa306t3AnGpcEMPrThhMCshIUEAtq9tyx4/SOaBtC
w6+vjsxIFXl1H6n6gvNquKT7HHFGpFlKtP+8AOx/mx2hBVndYQRxVCDKm7z3mbiX
aYe962m+PeauG7VFXJ86Er+Meg/fumriI7bO7xY49+U9bh3O3RVN+morhuFXRut6
M+w2PoiaNoEoCJ9AmhlUxuHiKTQ/c9qm1KkZU8FO2ysIgF6wcrS2XqtOkDF8buD2
/cE6iD13S3CbntRuhS8TKWX6mbfY+4UqWJ9KMKLA95nktnaGSjE3WWTSSCV+OPuz
xZg3WBlcQSW159kTTzc+aByXaed8r6e7HNUAPPgOTF3BvBpr4skjQR4e9JiJF6pe
33NhR4mhqgaUEbpLJjUMK9+MdrClaE0t+Foo9i6q7M2Q+Es1S7GpGxGTEampBFRY
IfonJ6ZO0sz5Hz0OMKqfvcA8vM1JcJ6xVUggXO2NBivhBEOHxwP9LFUg/YH9WtnB
JJ+lB5mSIne+8Gttw2TznMZd83dCFqsqMWY6KRrkztsOCsnzoXMrDERMDEFHSh0i
f5yU1yHljOcgnaO0GXkesodklGL4QsQ3DYrxIeRLVzV+p+le7c/omBc9YdfE8GK6
z3Ut33wlno9Uyju6+URAIDGzeEtZv7492KxSnKXo5RoGywokqpGm9AyXNJCKPE1y
E2lCHd3MKNBkMRCEqPkoc3m8p++wIolAtkUm9mAKLObpEDqOW1BuFy55s6Xz7UK/
3X/ExrneHNr6a7JE38zm30Ph2HB9NkahPxoI4gmFt4zRZQyradF79Mj+0LOEEOwj
cgmCol2hlHTZ0dQkyU2LpS5ZAdvPuVfsNcj8+ZIsNoo2Koj/9vKhJBS9MpfXhM9F
OakNel8wGfjKhP09SNTcEf3vqwgkzT0MMcwmQAY+yzsLIiiKrDMGSH0qTYCtqO+0
HpyahkRji+IU4noV87mskOLsHDbTJKet4tnvXMTM+V8NYrclPbPn4dyXEA+BEfYU
884igVD1U3w3FMXkEhlIKs0xv50fescii1xuIgmIBTzT0dbx0gx2A2FXRXfOAaw3
0f4AZX9u5ITgyiuy4HOB53pmvdZNFX17vZjO7xs0DpG/hItYrms0mOWbxXE0PpZr
sjvOtLqE144v98Bn0t7YeUAqnopdJ+NXTdTUHS4bAyEK4FhHB2W5j5Y/BdPWNw1B
DmkiBLutmraZgrhFHcVJ39C1bxIVAXoJ1DVplebabIeU7Mf9+jZ6YX7rzSuPDcMo
4AH3oR2lkI5bazkquhDU5WbcQ2+8eTPNXhIstQut6KLffxBhIVsV8LRqsKAkou+U
h3TcUMc4FXF8lWoEGGZ8WueqHA+px4zgLYqwj59oN3GIo5aH8RIPhoNcmONbFGcT
QbRRZTLGvtFeLtUiZ4AZTE8ff3kfJQ1o+Tt+fhqoo0Oqof+sjVbpQkAnEEHwtJag
3B3aoWGRweexU/yMGI3ertU9Hvfnobr0xfhHStxRywKvFlh75SMZ8UTA9lPBCwdn
MyJvYWJHccN+OKM7yrOAF8SYOJiE4gO7hY2uOViIjnFfNA41sEsQ+z9GPWaNHVas
QdkkZHSoqaIO95yliwl2Di5mMnEnvHeq9RSgbu08Fbr/NePV60G5oHaAMnFNf6h9
6HEaCtlTlEUdtwcYwtQodYFHa2r/j7UTi8A5ZzYPV7vSiYVe9Ttj21T6m/Nb9ytx
nb+lPugbrC994MwAaN5lX0pGC6w6LEQAULlhyOMnBTs4yYXrVagrLwUr+MJo8wWE
/OVr8wf/12iSfNzTX7c6IpCjTMDu46n6t5XDpbcvIFfLXFcFGYbEdNMIHtExtYsW
uKnxQZ+Eolhji2e0MnjxiJ4TN2Jo840es5ndHGR2yHdXxIwbHoiZMwnMiV+cNgfo
9A1OMClhIH8zKmjTreKP8D5BOHScZ9/CNrwSnVbdXN3PwWc7vQvfuCfKvMssinwL
K86nAMQYLInQ0c2PvCVsalN2W2rpc7PwXzK2DznGTgyZB5w20HKZ7vCI/LSJiJT3
ZwTdVzIEa5j3zQal/Zm7oms8JhWHFOHe3wODTeaI7JtX3vLG7cyuo30QzwcMX+LO
R9miT+XK9s+cFVxLWd8NTrhBWaQBWYxqp4iKRNPFZS9p7qtwB5zQGlrvvl/AUqRx
hc7eYtQQ4CRaU+6bE57AGnnre3xsi51psSf5NR7pIFVxy0dKVRkkk8LwEGdmla1R
V3KExOzs8v4GXLGXRn4LT4YuMsSsJxAUV+ldlIYxPjrb8hW/N5lFg/Uytsw+IU3j
djLSwV/pVnHs33WhKcbyd9t8xJj4N6fk2aps/R17ekB8AXfyK1g/PM84d5+/ZX9m
RkSKAa8VFoq+rhOKDgJ4SXzvohK+jpcwAKG0XcVcZkZxjFtPJo1cazzBwgtKw8xl
hnY5yIfaJW+b6FJKeeY+N8IdOO0uUcSn+GuINfbXHpT4kYoceg3CcApUgA/crE64
SAVu+kbkb41WDRTlodJUdNt1kd8WHxja/hI1tbiC3sX9PQotRHRqH0jO8pHjPzuZ
ZtRFViRZFY9ez+KtDaKDzD31tqql0T6ELgrtVdIQLAj3n+nJ1uXCqg7qbXkY+eCH
c+ONgkke9h+tcaZxQQvefnv8t1jfTRNAyJoG7gQEii2MgAkL/m64KqdNoFS4FuS1
++smpCZr6QkpdehT5F2kVmPeETszAb4L6Urxch/1I4qmGNyxlfmx5JHQt6Awhi+e
YRQ71jie6VTePLwk6AdoGfgUIkAfZYspKP9dw3XuuNmzpMkDRyL2CxXSVDtISUs6
yE5Ki02tGpKCFwncKb2KdzwJt2hrOSKIvXARrgQGLcRQA0Y08J8IZ5qwFzSASf8O
+ATdi9bTbnPr1CJLSWcEFH9GHMHEx98ZucUAUe0MBY2U8GUDno4/XHQtqQfbNLaV
ELITLK2JwB0Si4hQjU/IEa3hsV99igqIgUWV3DoQD+dBPYHuAE6+rEeU28dLqjmx
gF4ejrywbT+JyRfW7Mcfvt7DH99+zf7feVfIlXIutSuddxjafIGXqBHckpRZCnDm
Tri9sO+ns/YQWm+sw/mo/bi4IGQGD88eAX8YOLa8xb3d1ldu7vkEeST+gpaWP5Ne
inhzwPnEmumICbhwl+qJ0YxuxFDLAostG2wiiFF+U9cC3HFCJUJRNtSsEDb1dffH
pHmHKQG70QqJDXm/zZf7zmsUqkoVZSIyvXXRoK0yrlJ2w01wNvwY5fx3nNsPkxlt
rir7uHf18pVaYhQzhvODa/5BRDdPwzQ8X97arL02S4pcsdABK6qJlN81ea4/0UFx
hG1zeB0QeDKXbMTayi2/jrLcIQH7IyvCKh1G38TjkM9RaCaWTSxPQl/LmcR5lUid
vk14xQYVBhjzrLSoIlCaN16h0YSm5Fhh3EnDosWynv1/Fzk6az5HBOgayuIa2lPs
8q9sXg9U3LNzUm3c6DTGAjFcda+6+B2ffR7dgKWUfSNwA945fEhG7EXxJ5JhjJqA
nhXZ9d280TPXD0h5EQbgQW56feJmEIon/dCESiV+DL4xQ2Uv3IeHeuOwSzB9mUdt
Lkpu008RsjwevNp07Hgyr3OixU8ooLOsyAwLkUVywpW7EgBwapueCeLDDYhD6Ad7
NnWnLpXy4GtMiKNrQPyaZ7G1m9SSwzzigB36v1e9kb/36pn4afNMrVTRxN774x3J
b2dLL5o4lBTparAeYVvEm4NJIvVnaHUscaLZa5tHXfaufqnxc5nCRqipekS94U56
JgFroeOUx5F33Yeu6Gp1WgzCYnyfJMvuLMo2COmZ3GxqR+mwQVcWEMoG8hnxSvQD
rxObRtW1NzC0aZvrKNE0wQ0c8iENOQReVZTbfx83yB829pMp2isleSl6EgFEnhd3
j9UkhSyvPGp16fN0ftqzfvDQK1FyTdeQvpEHG1LJZCxHQfWf5RlAB4BO4zs9DqRv
JzQgPiBfXrpb+Qvwj6+/HVAVcoM/CYfOI93pEy5llcHD9iJjNG/f2Jp8/jXKf4/+
4vaXsyNptDX7CvoXMwAnexlI71Xo0/ZaCZakOBS5ECK3RQMbyCdUXQPBb3Eeb9CG
kvRmnwsRq73Ke7/TPcNCoNSLtwzBKMabEiIjLRMWblQxNgk9bdwCZjWxC0OxMWzS
NJGPRhDTrvn10A6uYkrQynh11R/mi4s4bBM0xn0hnu62ppbs8PmEz7fnaGRifim8
T+VV9gF2VZyyqjHM+v+lYz+6T/uIjgEEI1+xE+/N5SbUUmweO2siWUCZb4AkukJI
TzcuJnENnwRQJx/mUATkcPBjAJ+yvAa6MJ2Fr0fzfUZKZ+XYtpqfvr4T/Z9NP41e
xUBqOVgIwEuRaS8a0roeBi2wHWoxgcgiER9m8eIaXQBY7WTqwWQhhm4Z9yl/2IFV
Z8ZQ4WxrM9yZTojelPXode6/6596V2xPdcVRLyREqIDudjVtwCL5+RkAjajLUDEE
EyAGn4f5JOC1Oa66SrI5403HfCWvLajWT3WQae7IH4Mp5t9O6Z9GT6MPcKFAvvP7
9w2eJOwToN1ukmssJiAmlAY8mKl6Gubo2dHnOodAkLm9nceUO3a8+7c98DhrCaRa
qw/6qhKEW+heoljY/kRka5P5suROUHgVr1B724H+Jr3CmltKY2gvPsORCtxoGkSe
OMV6Ba7neBjGFO4/VRMEA9LShanJdK6kPcQYP57hdhl4ZtF9TIYWsyk6xZX1JCXV
+kZ4SMsdTWTHPxyUBbSUMVu751P45d+HnZULzITIKS5jZF6wekYRcQknRJHNeWwq
50HSj/KXuuMZvq8JIM412iZ99MaId4UhUoORCZiR+YMO7pHPRwA4wO0/H+zV7gtG
39PHVgFOXIBFJNGnUt6oZ85rjsdyDXAfm+vaFk9Uw+XGt4uaCYYNn6XCkbDsvTPR
6WoDY4zQo0rvwC4gruti0ITrMak6NWx/osJXIi+rBJXypS7JfQwJCGg9S8ny1Dcz
AREBXjGYfCCv4AKsWB7V5rVvu/oX+yblY47xNOrTFs1ccIjpALxYn21CLKze7tOD
OsQXUCZfFaXZ1Ib1JxHPuagpzuGbpr7Qp8PMmx7oN09l+tv9Dv8AFszd20bzEcTY
4Sse5OMQ/vyTcarHMpuU0ryiY2COAH3cwmvfwTGyuH+Y82SgNF5nP8vFFQ4bPJZD
LbMtPYUT8h3uE3yg01kVLiLhhyMWe9amBrtZ3gf1rS7kJ7/Ag53svuiW998hovZV
0Lwaq3QAgPKIoBZSUFKvkn4cPSPQQm9xmhOxxM94yjam7+SCPR6I4J6DAP2I3bZ9
IS0AAjCDpdKt+Crww9W55p8faiU/xdv5rvUPd/oE/pGC+8sW+74PTIrhUUWFk9rQ
7oahvUsHtgTrI4dt1LhWrmteoSunaQ4Uqs7Dm0RaDkn9Ip+Mtyp+zBE/lcVDi1kW
3VJkTBoYeSTvIiaJ8JHFwXZuCIv0pwrpURxaqw1f1GsmBye3nmQTLO8+B2hvqZbX
foAdb/DSkcbpVGweI4Dir94raJww7zDz5wzICecTDtnMlJIYx4/VoJbUas8Onl+U
yk383rp2OfOgWCVUz8OMiUaLPxsKIYnLQJ6ScPn95eZ9zVWly2LgM8qKZWl29ePm
Xr9Wj3zCHAXuNMfcRtkUypdYgD2zR00JqDzPo47WoGmUxjOr8Rkke7LlAk6ONplv
CsgD8iTZFBjAn75+vBZrfOXaM87eOWIoDoE1Yu3HV3l1go3CeI6DQaCgun/P8Eus
47qcTl0Xj5HFLbGw5g9uzVRP+u2w2dGwjuFPgq2NwI9vUFjmdV1EziOVIey0tllb
OndGxNvJp3DoqA2/aj3uYHsdPGyumaoVVPR7Le7esCqpr8swJyt1QOj7XDy+5Wh3
wgTJgUhzXGL/HFY4/M6FKK5pZQecOUUyMtFNMDCYTuWWfBfUcwVuvF9j4mnMgSEe
QoDZx5gs/co14HQYZf/wdfXDLL4j7d+Hp4bn5t/S5TOYXeCNNfw9mFI8eP06SLug
Xbj9iZcJ1AfhCOOQBrEgnUZjx0MKfk2cCWYrwx9SByEBd1qFT813qKm92zTgroiy
KTtoUjRNeT4LVpvF3T0LGB9PDstnH2LRbNOt3YxNTYCjWP554mA4/kEuvOrtNSLn
Tza4F4GJ7ELBX11lBYIWCXPpV9gldrcSBjkqR7sOKqkIRsMueWrVTqk/kLt24E+x
5ceFwLKJ+o1UcsKtTNFAvdhEFNE1DyoyeV7a3wY3gaCHjN5CQcZTjdsLjnMoEo6Z
3dFLtejch9pA27LudyWHjifMPe7UvKdJvqFfzRXmIIAurIto8ajeZPkvwRrmizp5
WeZziDUsedNOj0NOoVWNLGTpFGWVT5/nd+NK2RGY5EFnx861xp912YlyjcsANpTQ
Rhv68H0HF0K8xtUoaKALp9YA4hOADCLlMUmbiYwLK10tzpcK3RF8YIdlBDibMh1g
b8FqdEIi1LNnAQh2RGW4kZGzljmlUKSXF+Cgggcxdal3yLR2ik0TLkt3u/jLV6Ed
nuURNEtnqtHmgI+79FNv6HetU0tsN1LibGghgwLXtJchMrX046vKIm3yKhqo7c8f
v+l+zdtVS0fJU3K/i9W3bqvNrUx8xYNOlbvw6jTITpG9ymnuASzQriJJuf9L/GPR
+iNJjqmSaaWe+kffMnoIY0mRhgN1/QQazcqSMGnXKKn8X+nZyjvOFkKK82ZAGc79
teIClQStnT4eCuQA56Oo3BrDZuyf/y1CoaGaDEgQOV+hI4xpJGEn3Ob6AzEl7ccu
VyFOXu4v63z7x6RyKrnxShy43Dor75dp6FaM3y1u6kw7P4596vNkaccV+2dJobVz
2i2DX35ZRsTMjr0KU/fkqTT3wSQaO45rwkn0e/n/Enka0yKdQKnXLNqNNUFXK6oI
q4xmAuJqyaG7r/S3UuyEF2f04zL+IIR3VNhSW40r4uEQgXocmq+e28A5wclSZGxl
HygWwWXKvZ6+8G/mpRceEjCfei/KOjZJNwttkODWYrMQ7dpBoHeE6kDrNmbQf/Cq
3iiWTQGiAHcZ2I1BePNQN7sIkPDERcPmHwRI0vn85lqfBlKUuI9d8drF+1oqxEGD
2u/+I7NEif4IDS+4otyfJnCO708JRPtU//wQEN0YdNr1ClIsUhfGcaq1esou7sTq
1n/bnSVPLYHEtBtDQ5mCb/d6DcXZuoRrQAXiqJ8Q90vs+qgcZsFTfEoqhNOJJwWa
uf6D1zKYbqM6paoNnh0MpUWrcx4CTrbOIoiT85lSZxlNqATYwpjRIvNapf7SESWW
d0a38W032r5366nhwraLaCEC9dysYGSf+pYz4lQLYvluWt11Q8P+KTYFEw37SUQ7
ka48YIqQ/z5syKU1EmvdSW+iF+GmLW2lpVLe0O5WvGzFVMZKru5dzfiVBMA7ubr9
NB6JJbz2SuDDrNmrG4IapVHXLCHcNAszSc2qhrTfDmITs6QRHO+zcQoWp1jm43hJ
kNqIrornSKYFwRwrXUuqT6/+x9VUdkTTOkhZLPSxdq/9SnpM6dyR7dTFvf4nqk4j
d1+yw4VZMUw5RwW7uF3VyQtgYlLm8r4RrihTkbzdw2Z6yQBezIIJgXnbcwHKi7qO
FsYIo7XDW1e72LfaMJ/3n/XsyUgsTvPgGPTI2iK7mgUOjegfNHuin7qzT3esQu/k
v+eQJ+60FnhU0CuVO269HID8wc9rq4hSdhyKbdejbB1KAvTk8ukNiizbHWMZ+ExU
W1QRjzXyHcdFZiqHxdrTObjdI2+hGVGMxWwKjRnZ4v9aLKpnNeePxzTHwLy8Hqf7
ADJCGsI9JxM+LlUAozZ1DU4VxyRv2WOKFvHWuGtfVQeZAjhIEUwayDUUqxfEQBjB
kOcoV838r6yYYCBKrexb6siHpolge022QaIEQ8ME9BAzTQt/e1RhhWqZ3WKpWJTv
r2VpDOTX8nb8ROXBXHDTSZV12w9sDEM3wvdOTqyCBJq1hCpz4JJipVCaMvntLQAB
7eBX+XvovB39oOtPe7wPeDF4VbxE1vS3h1GrJViN++opC6qN+EFr/FwFMsv4g85p
/DsBiyT5OxAOjcLkFMcGoW+Yjy9KbkEGunuiXUJz0D37vA4WZ3Ff2XKKusVrOnfL
m9G4/rUBFxxLRT6m676GD/sBet77N+aqR+w3uYY1u0o+3YAA0FacDRxyBC+mIjWJ
cuR9CHDwuF6RFBgwHZ/d0/xNlX8B9RpsDVsjdGFyhJVKIhh87XriGgV1Vzjwuv/f
rZa9BjHyZ4KlN5kgxTMzyvL9rDgSUoXVx4z19Zegd2ntkZQMKNsBBRXEZCEk/C6w
MiDNDXuQAg7Y0vJhX3HqHCNoCdRj9N7mi9Do6nIdyIJThv3YTDUrIi9zy2SwFjYp
bEVOb55jC4VOz5N5BzoxAIv3DyjxuB7npVLeid8PnbQfuXsIFgBSqUVuV+dnEemp
VhabKQW8MeoK0ztgX4RtmXXCRcU2UtYMAJtG03qLY6LXOtuOd8MH/uShc/tatQqY
qLi1h8oYxdCQY5vEUIdQ24K5wcSaEGxywZA5nnkrKw0+h3VOsKSUgCJqOP5sdXpD
NEe9gJcc6nviZTqU98uhRzadEwdDhW4WkLtc6cPJs6Xk4qX0wUejM/TAhniXZyVS
LpP7FC2z9TmTV8fVVRdKSK+ReOYuoFOfLrBxHFmthLRvztw5eMZZi3dTIJL0bRUe
Uhl6FrDnrV6zHrjwjelhhQJJWwkpVXVCKTuA/3ZajMbWJ7T89LK1souYgSSzcJf9
em+u0Y1RkF7SJrLP8t6cjCXmetoVepVdtWH0x8ZaDmFEmKkmI0TmhT9QKqklczAi
88/nqcwwHW8L0OGtZyDn9TvIccfGEcNPqYGJdvn2HNb9qZA8tQ5RuAm65MbMNbj1
dnURPAbIdrNw8z283gfsjX0UrkhBznvC56l6U8n5w4GGUMX0GmiTxyQD+s07RIt9
seT2BF3aloIC+K7+m/JLMif1ZV99zd+xDNLXUsSjIPcxgnq84cYvgGncrn/eRAL2
BJmyeyM9T4E910WW6ySoC+FfA6MUCKJK+slxdDY078QvtwGNDyUcT4c6gblGUTzi
MqaDXAhm5P146rDKKDWDPzrFISdD1T5ijf61LKVJYa2GUsPpzTz+J7Gt7qyZhS62
WEEdAdDOHbqBHFS8GkD1iK7qxxRd6MBQrJzuG2hPv+0Fr5OZ93IDTTjwBDE/dOfo
IGM2sPannRd+pgqcql4h6Iefod7ceS/uA45PXN0LsFejODuAXC+FgOPFFurPiPR6
0IvaFezWvBEkkc1RiAmvlqFBMiKpq6Grhk2fNELbgKRdb2oEiAVwEH+XoB0FVOtq
FacZOdqnSTnLnZeiKEjdf9nuN4tQbTnEKQQeDdszoAdvQvNlMuCJtYgF16QJ7ZbA
CDEeIXpWrv21qXuKsco51NnD6QeGpnkkHL/ygXKBVs/4YE1XlZ4Ao6tabppb1Wfi
xNQZr6jvEgJqSQaETG6c8L+sYGisXfIWbPkBL1MGDTFPn7TvxPxmqtGkhSrgmsVk
eaNRC1EB5Lxg3aEJwHbzn4PeodE/OHLWmApW2dKmp2wDiK+jBsjaCuWv/LF7NPzQ
ReRfRxomE0G9f+NdPMmsjshpa6AeA7+THWl3LKBD9RIpQYk3RD2sXIsF9CLbYJMH
qR5MtL3c+mCfEAIYeeKTYy1DdjhhRKLvBn24A3xm9CGnvcAyMbilcc59qOyyjmkC
eKHr8p3teE9dopflqdufC5VVoOZlDn1ZStdlLlezdm89YY5NIukA88JUVvwWQBUu
1/rYjnPRrTxgCEb2gunoz/oUgjObaCfmvRLb5cMGQeX8pAH7wByQx72YfWG9Y5wO
FeadkNfwlJd9gUKuW428qR3p2l9Wl2s86eRdfuiYn4yDdkCHm2TeDJ+C2Iz3bV2d
5NvQ2YOseo+56s5Uhl/zUPKhOHAl8t58v7uh1FtdUeCSBGEsesV9yGYJYva0m8+a
tB9xk0/ZDXXtDFAuMTJfrBZLVkP58vVoPPURIw3x9bY1gJC7qKlgxtqCLF6o8ngV
l+mJqIbTWysSbXRbchuMxrws4c6n+OgkV6MYnmQ/Z5jPQdX7TqXl6Tq5DuRvdxlB
1wYK1ifVT4or284RNb2jjIyVNrTA7sl9OGFdYiSBwPC84AgR7xY8y5kgSVR2Bseo
u7k9O3qObGBi5DJw66gtN0+z745HROMJhi7s4KIX2NRXUmCHMJ2EovhjMIey79IU
8K4ShtW4lF4Q8KwwhvvUalE9QdqlLFZMq+DGDLIS1pJLrTUazz6FIZyIbjK/hVNJ
HRfnf7N/AaYUvPtcLHbeN9eZ28al9LGfzauLUKOCzm6fU4RXYOsV9PLzpm3k4rmZ
b5ljwg+2j/89o2ZeUgvP2Hg4yD3dzqzhsnbccVvYymxbNq2GplCaEs3BBhl1jv6G
Yn3NuVOEHnqAHY+BK3gVqzdEAikqBAxqkADjrDSMIwxo1qaCfH5semDpkynLJTd+
8/e14HfL11WPDZ47uurlFmAbQCj1ddKbvq9uO6Q6mvWN5n+7tTWLvwHFbCVOvNbX
IK/9srfDGv/9F30nzprsrn6lWCjvzBFvXc+76DPTV5g5d7NReOcbuKJBX9KCVWwL
X2ZgY6Ugntsl1mi+ERXW0q6vnvqdlP6HnO8JDLR5YE1ztbrB8Bq78o8rS5grxCXc
r/6Q/PeWxdkapIs71pVFjBtVke7/pqgIcDZoHEOEAiIBERQxp3nrwFvVvDi9N8P4
/pX20UQojb0mcomDySdQKqDN4jAPHrdW7xWqtCldQixMYDj+R2HffxqdI+lYXPOP
Bf1XIRRW7ZgAqPxCEVdH/4eiOJNEvaRxRHrQp4u6dwhIqPyALjN6hsMbrmZ02PuJ
3OOnfP2xoECa8+0r2ue8t/cGYW4EnB+UiB8m3GUeyYlTNOvIt6VX//8XM7mIcCI4
PqhraY7wmGfJXjnjD95YocARbMTtyzr/rNrgL+IItpX4Qa71Ei+3BL62yFqZ98q6
RJp1s1Z1/WDh4xho2xJIFLm35Bg4EMOOJSkeNWxlnYgkAo6OLW4EMZa9FxZcbeZu
utkymZ53/LecT4unWnqnaac/bkbXilBcpbkTCD7OlC1vBmZfnAQ5O4lPqgcA5Von
zMiXwcm4GpT9db7EosEOUjHzSqArG37cTOtu6uy5YUK4jM7QeGBO9PPkefuooBt5
FCopAfFzYLvN0oFsXdic6DMuEyjwZNlo7FlNWdMfjr2tJiqf+HLxS0/pvkkrMCT4
w0esgq63IE/lr+umLZfk1avj06zALhmW3nWCqDuF36BmXwBLM2U7iqsIJQVu0C17
wSxveHNr3K4JmlexQXS8pSAOul2YMujS3e0t8o/mVe7ul3Z4EUpSZP+yCA8vaFx9
NZvwLhp8aveyr2a2ueV/fmbVEFz21RcL43uyNOTF7JBk5JJdVrkpkKKLhB97eF1W
PPnZzCsunZLiCl5j2h8ZMETuyEh238tbyB4/GEjaKByB/IxAlB76I+yb7opNOsMU
CVdo7CfGerqxHwk7V/aek9wuF+APB0wbOpbjF1M7N0n9UIJjsppvMFAijetqiuzX
9EHlT7ob8C7ihLuM/0gMHn2sMWN8w4AeDDnHpuvH8XvQ6GJICF8lsQjWZFypHj3q
ZeWFNBABlrxSJ2XDYB/dkmf4ix88cKmDSDXBtNBTOPLSOqDYtCJ+nfTOK9FjsLvz
bPul/e3AtBDhFf2XlWYdrN2hcXxfkwEdzTGZ87GXp6DqzIeUEjXvV+P1465fr3x6
cn9RUZ+4fCd8cA+G2iqqxRnv8iwSBtYPQTHog9cWfPPt7JJteh/bE6TXyT6dxjL5
mOkCjdA6FIfUZ1idcCYzQ1NBXoHhn4nT/JktoEp7Pe/2egX7lmmVAJ4CmoDU+x9F
0xtFp31tBp8gplGgjfx+GO1C5P4CwuiHpGt7FZ7mPiDQ3vTdb5Nagq8T+Jh3iFXU
61JwBH65zYzTj3q3qxcybyk6tI9EKsA1vToA947EBdL5iD3XwXyr/5Z81wt5iGWh
/jPTfE9ucHR2va8ZgtnbHKq+nnk9EPVkaCkwx/3Q1oeaF27U19kNDwZE0IfnI0ar
pyE12UcIkeF4nNSfiQe5QWlfOJ0wcd75gTmyiK/5LlZp4wakUUzgD6iOksgeg8q+
CcvTcQh1tiUIWTcOm7ikkCl2X2h+CX2+o2H3Ap4v8l9UqwvM9P1ZwWMzN+KbzUnq
bHgs9HFKdmZWVV/hEDPJp/gf9i8y1ism5G30XXGdUDcAJI7M3EnYgMlthM95sFh2
AE/gar5MwmItu7yx5gsWo6yFwFYhGD60YxqamJS3OIl5Hbf5yAHIj0QoS7/G17kT
1/CiBk8eg7AZvWJIWtuw6WVKl7DwouFL1fAQocKXprVzy/rSEPFT7edzt6g8+ost
T02eeoV4PwUXsa+Hg5YZq/OR2XS9eVl4nSR/Tb2lAzS3S+U/Z2n/yHp8PiFBKt/w
03vy4OKzR4/cytFc5HNsNrAQ4agb0mYyzsOSe3Xv0W+bTzBqvywBGUyEYeK154pq
SeGXO5obcUhW44QY0w2oSSLK3WaRFz3lD9ZVtcvBvj3eJwMWHDnMLDHJ89pJ/cv+
FVOCPKN/9USsse44DTfQs1ihzfweDy/eW1fIEdCQan6c/KJUc+97mfP8pP9v4pRA
xEt1Zt+Vt+lFitK757M+jv8vw20SPq/q5P0w8QqHra0FbwdhF3Tp8rU6VHW/Ribj
jYYhaHeyX9Z6rhTn05N/Zx1kZj2HNImDlftOM8PgbhpJIzWtdYEFAcDw9g8FMQ9L
MGojpVOs4CUioks6YYCCG7ZYAi3XhaeWEyd1Hkhh1zzvMA9VD+cLgYm00I4UbiJE
5dBbUEyDrrIvVvTHKrwHtncm7CNBck6OWxOObkG/T7bYwQ5synVwa/hUBGgclDne
hMN0ngSm/3/VM1V+uGl/EdtV2pVSkHoUZmF71XnLYK6DfTgEGJh8fuXfwy9mZdFJ
7ds0HY2HUpgYjerEIccHjUN5iVXr0nTaZOyqBk2nLAEQZ2/rHDCKla733kAPlDpL
bB4OldvrBcY3J6OEg1aWeD19qhYGhizlWi49sk8Usl3RqXtKetv8PvXQ5yLdgBUM
FtiRzd6/xu3p2NrNYVeMUh/S4H/h118n5DXv87Qi5thEueai+izbHuPHrGdseyKr
pqOQCt8+weIFPD3wIcOqbs5bnr9tejT8IUeByxOVcjuVrCb4hNhE1qt5Ep5yPWRJ
U4JbtNmOsTYHV8hKTja7X++foywFBasiZgm8Q5sjLiyBJ9JCt8hjj2pO64KRF7i3
yOnbf6tqX+txnX6vTWhkBW96R3f7aXzHSfSPxX7APlFOslCdislK8FrVhGm8c6tn
czJkaUfQwe35oubl1ormMJB50Bfr6K+iCISzYdE+NDoSYAUwtN8Wx5Zz4xBrFTBw
Eqah6Dy5/KaQ44dT0FPn+9y/FSsFJQM2l0MudqIO2o3HFSU1N85aE6SRr+4ZtW81
M2NdNSPw0hp996G4XmLVnhtwsaLBvvsvGr8+wGGC1QZFUVsoxbU5YxM5NEtLLE+w
sNHjNwBgL7BKRj5yFWu7U2LR1dlSh+gRI1g4cgufpScBJfUKlZnCiuZQ1/OsTipx
8kSFD6vuIfpqM3Luv8d/R8fcAj+dAWa08eXh055IvoK1p1685KGTN/Rxa8xcysQk
gx1vR16DA7Q+nVRLbUstO0knb3n5qh9aEPs32qh+CRWTa6MtIpSg4QkHA13i2Et/
LKrZLl0fp9M8Hvr7Oyw1SOB3yA9sqv4mIXdmr3tQDxBDX+XohcgDfFxS7qb0Czgd
Oxbp/xeMMjHXU3Si/Qujs0p3m//yjP2EJMaKeLZ7ZTqM1P1wVe48CCAyrMBmCEKa
sUmtpxV9c7jV13chuRcD++ayxl5l7engISihBnO/r079adAInqd99xTYckBZWsWh
p5ospsm/0oDyszZglNsm1eDXvnsWRvXYNeYftezj/GhOX6PuPFWnuEiF5lhPgQ06
eZdUX8WRpCYmaYfxa5MtmEGmdJS11laAzYPjR8EzRTNyqm14jArAwSRRWd/H9A3H
2U4rq5+L+7CMAScOmJmIgjVdOfkLz9cCX3ZRqBE4wVwUxpGf1IMjkN1ubzLytCe0
9cLKNZKFofOytjM2QG6WQtqa3xIOF7iUI/PYv4C6TuGbbexuNuYLVzZE5T+g1Xdl
oy8FR0KAJCji1sZJgWvb9zjGB449e45xgAJG5X9tMMj7wF0ovyaxSSwiBw+IMRvv
5up+YtiI/nBgR7N8kYGXaXSZ2jc9Prqc4zC8NhOraC44MSvRuTlTfvjAGuSVNcoI
Eky/6pDqo4ELVT/j6Y+EcopzkzrRVD6hrY0ZBqpIkuKJuyr5qQ06/W/Ud5EUUWf2
HarzWAjeCjhRHuCTrB2b2WHPZoUUjtaUekDsJhs6KvwblJWxoloM5i3LUdu31c0U
JdOm4m4fxceLQmOcg1aWZ1HxT6e3HfndM4j/62NTcBqmTI9E+PYrr9O/BIfN5vA1
/5gQUQRpRO5lRpkX5YOmiupR2OAA5nF+momcAgbnWfjaAFFWnlAz03wTJ+7VJPpJ
3la/QOF3Mh+o5G4zPW91AdtW7NvsBEjDhh03TK9JX2kv3HkoKMMQI36PbpQ8dT/j
Y+ICfcmyCruHBkMxstQKtEMws7oEqEf6pz6a8jBGMSrDdov8PAz7SFS1/sbArI7/
lTl/QE6R3NlApGgW2WQMPM15Oq1VOEW2ume8w2IAtUXAiqOb501Uw7mZQ8AIV8cj
yMp8hrp5b7N4SF96/iyLEMVh3viGMo5xOsHegkulShokDbRlqFDxL8BJeqVgmJoi
Hf1hy1exQXARrQcdEHOe1EIc8zwp+K5TdJFhgOFd6pDUM2ElykkCFNE09/w6W90O
kej1Mmi7GF5Y3rCKBo8G27Xgtn02tSvMCVwpbhnDzini6yHUqR4uXAck+qbPnshc
iw75l1dJvoKU6iBQioMl1s5++KANoxV42cVekQdbztWyzguK9R+Tm+FYJlYDblsh
m6VweWQ+gbLJcOGiS1z9tKJwUXaLL5CgsNdy4sPtGVoZnwBRt46mxpGUAiC//UjX
/dRsywOCv84MZ45D9gRjy3Fc38vK0mWnOhKq6diJL92s3k5W0t7fTrAKmWwkkkgS
35bP8/Y3wQ+fpnobBQgAWMZEDmhJqLBCONDkVKQo3rCAZuw5QM4uYGaVbd+sUF8K
kGZpYykCpNeiFbZK0vcGf4Sf5sCiUiCs3h6kcamZCvu+fM60sqtXcIRXbxXkjPNq
b+uitGp5FyKX4gC9N6O2Q/tKKSdsMlwSxcx3nZ/GfPgBB2Uz7levUTa+P1oveuil
HoG3b1+btpuNLol+FEuegg5Zzeag5OkMhk3MjjuP0skvmJyA1HxIX8GJQFuunWTW
NG3XQeyNA9FQcbAi9ZpZ8+LnRsAV3DTtbeU7mu1INmoiNzJhqnHcxJYLZeSpUu8F
KcT4ORDBksIi5JSVIN10Dc2EAmvBzjM9ltEK+tkpyVlSL7eeKABnKYHpQdYbRfXL
pQ+SUnISUgcY+6s6s5b0m1kzGNIcKT+LFbR4ZFCfc9vZmf9QideuV9Wa3d4weyua
cP/RwZVh2MCsHBeWURsMeVSHrjjuM1tzFQ2GBZhIDo6hTrWrSQNTHqnXba8ocK/w
3o4txTks9Brt9sl/89DIyVNC2At1YiBt2Y01WU3Ok6rIDpzZlr4G4WYNnjWt0fFl
8rwqR5S5LdUSQH3tkVjC0loH4Ln1isOxsV/6MFLf0fcu2ULZMKcpKwIXPTGfgJRr
Ea4YGb7Bjxfr9rBnp4DQNWVIoISMe7YmqSIDDHd71kZ61fZ2/ojaIbAVlQCbWDo8
hI4GUACP19ul85C3rnRxb9uBEb76I8Dwk3aZk2OYeWzwo17cHQzevVKiGQ885zgt
+bAxQkT4tZNrPcQCP2caGZWfhWdfXsPaAmkpiYnzqkbv+4Ot6Jf0tZeoLeCRu37i
FNDM6NGkVtdPkSbbYm5BWkpgtGuzyaU3sEjBuymsnzNcIOpjtj76zRQACTyhxFEG
vtbK9fdEhuLjtx8IvdJqbXHIlM1YukyLx1b4psNzwFtDS98TUKC0A0BdwW+trZKS
AeriyxKUCSuH18WD+IJIPqVvq/AlPNgow4bpiTxYENIUxePHsrGopbxQxVfxOSFF
DQhRONhl65e0CgznJgMpqRHBy3nNaOETXYOI5gHEOWLbfuv1SFF/m9mHpGjwOa8w
8hpuvW1YZ/9Hvyg9PeTV4S43pg3QiFERUG42s1UefOw4S1zMAicJ70jvkYIdgpZu
fPbL5ZuqJUCkNTtbA6nYDDxffv+TsbC+b3xK2MpHWOV98EA/UJ+1ZMdtvT9WOgmZ
7zLtzvDtu3dM4U40SClfy3ppEp0W2tMCtUox4/WyBzt0EvgvPvqWPoJy8nYcoGgV
z1SLMnRLF4zGS+HEMQZvmJewLX6ZGHDeelUGQrBXPiJv5qz4VXYTi/hfBbLReAv2
5cqM0azXjwNvZyYzall7SIHQ6BRAwp5SRq2UXjG40xSP6wsT/me5yHqP3/lvCbEL
GHiZ8wN+2Hfo0OXAGjnuIu9JbIRljH9joumez7EHhbe7sjQ5XhF+UFoq4VaEd9Ls
NA2qXdaOetj3LtudUMpB3mlfBnyNLGfO77Q13SkoYYMs7JB7TVESQlSQKqv6wxxn
nFlZ5yccs5vDRx3Up+UeCb/03BaES12f/Cai0g83YTJBckFEKFTCZ12yh871HpMu
kJfbcP9vka1PZG0C3lVAu3437zEvMZKt5hFxIhBeuE6Ipj8fOTEStmk4SXTU7Jwe
zPF+2XBeWY7mCJbXpmIwmKSVATUC73UZYhAistZhOovvtQZE5z+OPipaEK+YCV0q
ay043KeB8USv9k0+5YqpqG6mMGkBzIcLHBuVIjaZFyT4MQNdZUhZBx7lI7J59W0n
aEQH6taUEK+TQPFSzROYsbSvlAgUUnZrnlbkCA9h9MJxKevHm/u9MyLPrB85oz1t
Omt6bpqXNEoMBjx3+TtMdrgcb4ZX4AWvmWL0vDpEd5HvL02kLRSafTzvE9QsrsBv
P1IPxl11HxXTjhyOJ2ZA2kOqrN+4tvpp41fw97Ngb2820UtJbKpCQM1waRyCrTd2
+NOWIP0fFVuf6iUkwb0nXBjjibah3NxqzhOepM+6GQU7gRTseYxjXNFTOgqW3X96
h/iWYmRMP8JL6B6OEQAe6R3ZzTRLyIEPZqXjYcxwT7rIwqIIt1SZFJuU8VyK69Qx
OArAr8+4ob7tJT1UNmEGpV0cpYPn8O8IH54km4K1TBVJ9NlBAvgQSFVHDtl5UWFS
BuCRo5LNlorGdOx88UqYso4jBzNO+i8EfyfLX5Pf0tkvMbmy/GfHsJYzF8iTQ2wZ
xohuQCeiG/8mL/GyyshoVLfpLgrLEbZsCVf+c48IQXpdwDBWQNFJ6QcDSa6ugONv
6AJuH/CSE5aPjh55X/3Zq9KiggWMeRlUJc01lVPu6aOll5NPrQg/rEZtgtyhcdal
wTiSnkJOIZ8wglQX9eU9pdAF7ZRZ6rWDqEYjQy7nWTxkz9MQmaAxmwl2JWdgqHT1
1rsc9WZn2R3z+RDIeqohVB5hR0YlPTZ2hwtsSfd5Mhs3HtwEbf9YYb/muN6eQQhd
QrDl1MZ+IsjUgAL6aNBuNtENsSI/gb9ihMEOL8p6JCWE6bHoFgGsJgrE4TT9MJSt
aHB6+YRJ1mrZjVNTRGM+vbxN6WsB0q1U/4NfCR3vdpKCPOWiXbfO76JeV8f5s+lQ
28X7JmJOgj2IKEsS3mvRendgb5FA+T5xun7ulibMOBmPTAsps/tpXxckMBXRpknp
DI1fRoEv38FTo7HMqDNCEwNxRmuG/J6XVIQVvC21QVYD5hFY6tuz6T54bkqQ1+iV
0fcrCj6xvhUnewQH6V+ZKbsnLngAFeUS4X9mlQvzeV1YuInevl2YAXCJiqVTplV1
E42g6fYYFNMVpvdaGnuAuUpcu3ajlNaYTJEjPxAiZQ69cr/TGzWiPyGPQv2nbUf7
uwY2z8pBEzePmE6Mltf+qaLX6VnHu+Aw6nZxeBFPzEqL35X261rtm4yAzSthf0gG
35jJJ+KArUIreNRbOC+SmBp5u+7gAFqhMwhpLFs6OZra4DzHFVHlJFjDqpg5YvkX
38V+Me4LAkGgcYFT4N0wskJWIQ/sA0ZJuXGhFksR2vTceWR+SVtBIdL548zTcz0D
n4ooq6cWbkgMohR2KUj6EIP4Kn5y3Z38DRx+8M9YdRYObjVPA/KdwkGvbtdYrWrG
cV0iJEncbrxFw78nJYPW2R3Kb7bE3l1Npk7EAwTVT8MKNEq6gKUIkg0qFrpLRdg0
mjz46Jmuq5w0JMWlRDk9KfZO3UYZuSZPGS8vU50+3SfIzdLMgE74V5+eTVgJeMP/
5XlPJO6Q6Ht2/a5KUepPX70V7Ne3wYhpsrBqBVSDgfZups0nkVf3CzEDdeiN3A/o
T7R/kHWZKuWbAM5aBSbfuBI5d3+2qEHVaWM9DZuTEbsxaZpEaeyYX7fPq35BQ02G
vl1zB08u61WQTv08S4x9Is1hj6+nP1/G0BaBtkOamU2EyrRPISyMXHQ0asXoF0s3
QW+FOTEYu9LaZoVEHqP3UH6HzrhuK5z4vmNxPv497yeb0Urnk0KbgmTAxroSbPWH
RPHVbuYxFcqfyOf9QLovJt7ljcBJ6FYOVlwfe2joB+9En/SjAPzLXBDW5j2Huy5W
9WfLT568uyxp9UzImNy3SrIn3ztIWQFIq+qDbHffO95usZAIU/oCzSRR3G+g/JVV
F9pie3KZzxMEaLMeQ4C7VyA33gHS74jHoxfi22i0qlc51OnzT8kNdBeUSGkcXabN
iSjXxWMm/2sqHhns25ZqCcdxtVBQh3Bc3hRQCcshF0kroeEpXguvefKV8fIX5Q71
Z8vEoHUWbD+4ylO/+lICM5QYCrHPBzM5gaUAy0yWVrSvMifD7hQYxEc3ErK8jBB9
uauGg7MaGImkKJJseXxQP3kXeiFD8p88lMveS4Kz2DL8tp4sFu9SrCfsJN1zp4qQ
51HoaIRC7fD7IrPYSQbM+utWkFSUvgcLUbzWPYajOrP7BdfxQl+pIrH6j5Jae5wK
hZznK7D/tcucHx4nW7c4sC+E+1pZ1fpt+xLMWsN6vOPotmbEtAdjgwNGApQm5ZvT
iqUfSNR2KLkwKIlx6lrOPh8M50feFGziATTb9J5XwsNuifj/icNAtUoQJvJHGPJD
2fpHOa1xxGFs3UqSzy84CBlOscTj4vq9l6SIadkUBLCgAyIDpAVITH9JvdTU2QTg
TMtO8Odj3bzPZSguc1wN1HZNOxFSMlAzkvbfqn1FsTkhDSJRJQ4e8K2hijhqXIkC
+BioaSFFjrfF7NeKWNUPSXouzc9mjHoE/HaFQOIx0GAZy11L/QzuHJr3R9A0z51p
srM4s74Tcfy/vY4D5rOCl4xNuKuJAzz7+gQcbSdxqd2cKHivilQyrR/1D4wL3ATG
AkVyXIl3pEMHVQpTynZhA5q7J/1r1PyBzoZ7cNJbZt1/yyzWVOt9IB1lrnUFyS3G
W7Bp0Vo63makmMbnPRhXsmoVcm/KtXYJkNFMc4fQjI34TRBuSuyBuT9By92rGlQU
UDjRigkyupAx+V1JxFwqKytlQf+aExuNTZldecDvA9U6e722Qon+OipwMSRq0kPk
ZC/FT5OZOcqhqXXepwSN2TGdM2lbo6LCmogAXhak86WEe5r5bvRzh9ykhYbNys1e
/giheGFMOvutXFwIz+FBE1bwWML1ZR/+CBZUh5cu8GhZtmbPJIDFYaXmGO+Qq9Iz
zbrrtb57EyLQ5MYYN1chXVAQgkhyStRlSvGdIw45Pm5DvIc/MYnEkQPQjlSrNcOK
fQDwYUbZIsHfscZ/E4+RwqchZUfm3LW1Nvtec2TfOzDkfFVO2D6WuNYHJC/10PWX
2ORUmZeX757hVLvQAqdB5gCnfU+lc0WJ95hbZkfIyjqvONyrQwMdWqbn8rJMSVvr
1cWm02qbLGGQ6VnCsHodoplCRGr5I9nnUzr0ErTYUKNStViVHHDUFSrCERUSP0FB
3bszEmqLdd3y9Z+AQ/rs+biVNTvULVAscjEakfLF1rixc9XJPXibsHKjA4JBjm4B
F9/eP/vXD3aZrOuy79tfTmjLyFFLJJqNaBJZq8zlIpKHBOU14xWfElsNxqWcWlZp
t3EGBznYxf6cQqMPjFrRxrZjkWoXiF3W5hfYEYQj+yP2YD3NuR+ErSJsmfzHI3MR
2XODuQyVqGSz7Lb6Cd7Y1z6m3tKpi1RHQlLhI/3In5flaCUuCYwQcptKaJK+tfa6
RjtVFheg5jlakaoYZ1Xb8XaXGHKYkn9M64KTuhc16fiXnPR3Z+WqxhlTSusoWP+h
7DMhsvuLSIBNfO0ZLujxbzMz15yqJPtMzOW+hxsQY8n8taOqaITgHTyRDyNVH+hv
7LXNrBfeta6qA/gUzRYKKdcvqR/3OyagBf2e7tu22+mOpHDfmOmV2jXAL/wd9JXR
E3Rzl9pWjP/wg/wJQJXKQxSGiYhnIKEm1oLdf5A/+RJQW4H1egFpxymzWMrL8gUz
ckxHK6rHGfBBAbQa/TqukOJR15mTNEXwCM/HMknNszMHb2isew27N5EVvYsFWcf6
Yu2/igUOmXDJFt9FktNI8x7EGjn5ktHVUuRIzsSDLcsLK2SFcdKX/+Vxqe+KvLzF
PD3J4k+xEkzUZhoXuLmrbLyoG4HtiQpfOcpeoS/lkam+DxiUuvNKIEIsiZ1kR/Kz
uD1qBkLDfPfgpEP9eCkoOnHRHdHtOfi6nwCa7IjN4uHRImy8RmjNGetvlFYZwq2H
8J6RFw2oTLDgGoyNoOqUQ+75X8jzkoqxspemDhGABM2C93chUSCSQWKuzLLC4AuG
f/1LHKuyFHaDLOsNd0177eVr9JC6M4l9O5RyNjr/0v6NY7sOPIpIN5NGLg1996bG
eE63zJKGfFM+s3MguxS2/Z+xfJWvnTMjTWQq2uUhuTGpB2YMVEyfJLB79Fg7BG2e
5EuGLo0PzhS8dKItslMQHR7Uvzf1zJOPV5t7OQVRs7b5mVZKE+YQEjXdgLG/AsGY
roIzgZP9yydIjp9oTJopfs6X+SbEbgLdEW7I2ahG1Ob1/t5VNio+30X7EtZ/OkMq
d3RjC907StmHmmngYzu1l49xFYGFuSSWgZQM3zeND7H7eWsBdycW6+5QxrRIR3ko
2b0iQYhsqz9Kv4pQJdyyTxVIFXpYpVqByLCzRx+I4jit1dw7zowAYsSoWs/B4tGi
hdybrkpjCtr6sgOx5HECn96qrNGwR4jAhoGBO2OHpyD4R8AkrK1tyFTK8A3q4Z2Z
FWKkPNKo6gwUr2KyotsGW1/NPDpWQDyB3BSxARs4aASdFUJ8heGuM2AYCZm2hiPe
OHadnSYI3S033VRxikBkflv+FxO+IvgZZuvf0XAozsjRDoomTzHPLbpZRtuml+cR
Eodr/K7vXYHOpiKMlKc1ReOj5Iyg0VXWMSVZklQPf5sefTpWsEK8Q0L7hM7hnGIT
iz7unnxi4PR2tFxL92OrhPhnwJsF7KWo+CuB7u/QhxqDfv3s1fVzXYGyiSy8i4fw
uiH3ZI4mtlIHLzo4XA6R7AWNdcYcDT0d4k/DXp3aiO8tQ5bzgWDS8znyeCOgWr9F
LH6Bz1JUDHHbIhyJZd0xnaIr63/Uoe93D/25+LugjpmmCHQZdYqW6n9opjPmkV2F
8BH/vwzDDsZjYLbbJBG2T8RiCbra9INvzBmp+GjnMOum8mPkT0vxigEaluwCZFPZ
JZJpA7Bt6bqa66WCjq2YutGwN9mCPc2m/EOtdP2izInbaWhqCofiipcLEgQDlOxm
vpSxexGGE7L2YQeH/3FSgIsybNxE8JvRPimUhHZOwiGFopoqKfl4AdDAwWSUjTpG
RPR0JpdpusRqvxLuiQh7Kf54uf2CTcv1nMhUeNcg5ecV3KFXZkSS18VZU2mmtTZv
tDfbYZXexbaMlshcHgL8cd7iYgOx2vVlnoXnEVqE9+UzcIRZY3D0/lCO9fhBTuvC
GfqBMNDnsVYVepM9fDr57Mgpd4lfAHqJM9uhNkUhwPvcEeI3yNxKkvIp2cIjOYAT
jsbnthdw+QYBrBb9cEGqidyjjUZFX/kL6uUk2x3Hn48RUXJh7rPDunUKxsnbLdYB
mNEcic9edJRnnjpIQcoA2LK//mGs2D6cw4rmWL8XgE9Ut7VXWygTdcSm1z7fqmvK
JT/R7InwayEP+SspimrxlHhXc0Hhuyy59a34IhTMn7d7+T0bmEKC8nlV5VLRsJyp
e5wKt+nXH/JNlxdJgtumKO2OR+uU+MQpm1el31PhBKOngbLnb5rXRpOOXkdWh1Ms
/Q1L/XyYHaQcNqEwXc3gErsuh1yUBtOzU+u6gXjJwyWdnICIisCxlT2KFHvSS7fy
RlGviyFjnYdRpyVWr5P0h9VttnB4FYMhHdoHDuDX56Zs5EPhitFIJqckXiCC0/AB
MugpPDoM4LnI45dQFwys+nE6TgHqchVtlzbD2165gT34IZEzF3B7/NJtjD1B1G6k
YQgMAGl42jAl1BcjExpgB5cRBe6spwrOpAWe0ZGn6rXvo28DdHQ1GpC4kG8dUID+
DUZCyipYLP1EGDalsG65CWAqYqxxU6PoA5ddTcxKqfAOJu42JssIMoAG22QzsfeU
PgBLJMeIzVlr5M88xxdr0hxfZj1bOYMSKAawsdvAkGtsLIf1CVPMfRAc5adUJcRP
FqU0R4zvvvcO1JshF+na+/Rk5ipkE8d6LUcqT9ah+NBS7oirFbXS02VHFB9oMFcN
46p9UWiS/MUtEq5rEewcG2f/OoZwftLFZ/ttoo2XlVvNv0NxZ6F06NS1Dl8uFAXb
hbxaznqp4HmcAZLrhhYc73tXkSj3o5Q+P3TpRbAQtjp1ADxY5Kf9Csoaf6Ol5V++
ZiERbdJJEZKqV2dXRwLgSf7IQWwgKg+tl3cwcjOQf7AzMTHYaLaPh9RXtaUp022a
UJ30+OpFF/6ZqQ/knt9lzLqitDEJ6ElYlPi3TuaKKa0mWO7hPD6CUkQGYjF8OZSA
kh7jomI+kD0Jytux9zFWoqoPGNjFlOwVgBpyCNBIjnN4I4wG76uY+NyfVjuigjQY
tj1ncj1R+/GfFXaDC+QB4By4vFsdPziMGObFhn3SM/R+meOvfkSndmX0ptM/9dOH
74BG+EUBQXMYoTGaZja/689WyobwC6Fzu/6inR+tBin135gBfEqYLZIuJZC02nlb
e+QxHnfEvfkePWlRZwEegk9G+Rx/QXe7yXSUSH9++XNlBjRPO+bNiyIRPa3iBop0
nYLC88yblqrV0oQSMEXrsZuqO6y2ARqEulTHQcczc4YBDQsl/h+WTVYIyi78lXqF
J5J8YH9d0FBSP2fq3JvuXuTDvMOdKHeIC5Bqft/r0ykIWMDb/cz1lLyMdW6DWfhZ
1PF8DgFYIS4JH22KKm+BVrzxjAtZMH5BU5ieRESUh8jIeWNNRH3wxagtKYcQywdC
+qQ9H9372SMe5WtdK1YQyTxJ7Z6EdjwaKmXXNVJrAY8IrDWO+6wFWC1Yhrtt21o7
5p1C/Zs3KTcjrcVhv2QAgmKM/4v+GNAUXsaF9M19cj1qXSlfOZ0rlZlUHQpBqGsi
mCZ7NtAGvV4FjwtfCWgvr2xXCLmlm1XCcNdc4wtGz/Fdcs1N+A30faPqxVMA5phG
FXZzY16E0tIm+8ymN8wDHN+gGPWTzOiLAzGiqDtwiO9SbgmyKD7ZwEygqjUTojL9
Yei3QXVLWIvUbXSD6EnyM1esYbHJ13aiDACnINGGa1HtXs5PjRYKDAzWpyYB2wUl
L6n8lpA96JPvn1L+1OYpLLQHU1nl7w29OVVHZBVriyfDwJRYlymRpaIslo/NtoCm
ub/fB3qgSVQjDO8x851AHr019DihZHQLGFcOeB5MRMNVlVLPLfqQ8YHZBsnM09Kj
+OYsz/BESz0uGyYBDKol0RupXG0dFkFPkwHgv4roC1TJH2NKw9IkiEC56tHaAgFS
1e9WiG2dreOXwghU9TviTk5Qugy60a/YQiv43ovJv8eczXC18k5wz7O4oIUqIjac
8pxI84hOP67iECLAcogjIM1AZGxFnR+p5mwjE2w0/RIrsSxI+iI8x34NMb2EgCJT
GtvHkIRbmmTUBblQxq8NOQDdaqIQ1rqSk2zfbes/Eb+y2538FFdnQe6jkI+LIN2F
gQTmUPO13/tk1IkkthFydighnP0wsUXqgTQQLyjyQaC4rZL17X+g0d/9B/diLCe+
kTFD1EZK28mE4Xz2ulSi+aI+8M/DLJy1Y/9nZ/j7/VIuQCBJTmrXRWi69DNJX2K5
AWITZvwpwNP5RSLQLlmH8WxYQhIg8O0bGv1k5NwX9Psb1EeGoaQR7ymiNOsBL/f4
BZe57LAtOn+Dq1Vk55HyntGYaz3KXsaDrfbo3gzVs9O1cn6I47PDLj4KKXEWqmq5
MgmVy39xZlIbZtkbqSrAhy2AUSPENR69ppW73MohhhFDHiT07FuBWySLhLtluiCf
3JLDVNHF6VadR+rREFA65rgVcKJjzwI5Be2F2K6WRtfB02WM73FYJuP2bY8R13bB
ndm6st8pnZmS9kJ6j+By5CNOr9EicKsKhxFJVT2UmaS5EjN68qMFDTnDmlHSqZaI
0s1UpDmKot+1OxSHg9GJbVGqFKUnAJ7RztE0N0JykkMBxkt6Ky9VT/ttvI6p+xOV
nLP7qZHb7yQ7QoYmhyUZ85VB76K27cJ+UrXXbvMGryo7AUsAYFwr84b294ppbIku
tawltgApJW+iylMSgq1xPIClH+1KySKyIl5DXDeSEuKuUrVjuTcNRCeHTB95gVZr
a3GH2iTW0mCuyfCOlX6VKgBJhQ2aPzsvn3mKLZIgbZ9a6Lc4XZjvpvAUwmbQFxC2
ncmhD4uxvPDivDsgxyWuuS8+LyQghM/FojdHcl4a5uJSKp+ddyFLogSMpVvSKi4U
OfDyJtU641NGXltuOcjxGnxEAvInVeW6wFAhgVMwW7bmp1CACNzxTJixmz9HJ455
vk8Ifnn4V7oLuMgQlSk/ViegBqVZbT9pA8F2GR3+anq8D1/YzbUx91NDWXhftSZU
deuZ+RudGQLQEJFyNHo3jZnd912kiCf20D8MRi84ZquRCeMX5sTcs04bOYaomVVv
IqDYNDwao69skc77/o6p8E3RNyFlx8Ui1Cu2XPd80Qj/Om0jfxyOWyhKJK+a1kRv
kXqqH/IDnjZxzoErGwd6LvKcA4kZBzU8hqEJBqrbmMMO1XRLSRkMn3hVoTKKMvKy
zh2XWopLER6VPvGS+cXJCB01EKa1sqQ3gFMRYQlWKlEpHXF+tsbOsQPbsw6WkTKB
6Tf3b4jAO+tEG5NqO1YCOqtcsoeFMxrQkNxdG1HIELTSfWJqBeP1PqLod4RICaI3
SEY6FssbXmbGi9zBX68DZp4CwD2haFQw6fSzPvR1e1yQtaUG88GTPDWmZT0qJwVp
BvYvgJ65FFAnWr4DZG4PXb9IRYkCVBWORADqoOtXuSMCkr5V11vVXzS82Z5NZDS/
3l8mMfLTNJIi1Li2y/bCxwmbp+F08J0KBbG0fnKNCC+wPT6JQcLbaXdNRny9bdqu
gLmBYUOJ4VCiWw6eZV4vzcaH50KmRjZ6lMtz1IDcfwn+hpaQKOdq5sapUjtq+vWP
SKjigatwrPKqvqACQM/ZpzvUxRzJ1TPZhUBYN3GxGp+weyQ9wnH+EvuDtXcrfaVi
ZPrYXcDgyAvEjknr2/lPJb09E4yJYm95y2YK9Lu3BPpyJzJIkz6lGzBjYOl41TF8
1FUf/TrncgnA1H0ZLqwB9ryA7WJQtuDkPi4/sjvBDSAAqtSczWVvgifv2mOUqLai
Y6sajunOJjVKiuWUtr3XgFQ9BFdV6b8NeGxzkOPMANfp1mT/bO2Ts8r2NJwT3MJs
dSOHIcSdEIW3dRZjTWQpPhnehgcDOdcPrL2KhcoeGqCTt2dgZGNQlh07J0OvaOGR
b9mxvv5ejak8Kki3BJjAVKP26JfzQhze3W4eghrXhakHzn1li28iBuiTkPoJ+3/V
kGX+wpnN1mY5nICECc2fUrLdP8AWsSnreJbYJFDbFxOA/QXAqcRGIA+a7DZvzTEJ
NUFcfuMwOrm7Uo56qZF44qkcfuN8vN7zifyW4vf/6Iu2tMear1zeG+U9S5D5lx4e
pVzQIXIKIRaT06D33d7m/A3uUwFznHllYauPwfi1o1lKy4t4xhY1VOlz35wa9NfC
tLMqoyxgbope8/xEA8T7SK796fOBUdqlssn+ZSbTkKqkmxCTXSA+6GLmV7KRrhmk
d4Y1ztVwhIIE/BwWUSv/7v6bA1x1YDPTbWDukkY3DqDXzb2MX+8N2rMlSROUnXUp
ZzqSgywGMwqJ9tZr6+zNCLF0n9Twg6cElH4IoknCFBURVEi99SX0RNKHYzJLhGfL
PhmAMt+5e11dObhlq12zXuoEHj8PLAUhe4g23MUk0vzTkVoBofhWkVY9XXyralcH
+wI3I911IMtYnwDMlt0wWiY2l4W3IHGcLd0VcasoqWwdz5Tn4pZcPPZw8m1xtfns
5T3l5tdcz+JaMaxYVg/AG63mRX5u3wPxs7v8zveG+qMxU7fD7mTAcCA6hi6CeT5C
uAqzrgZ8dlWxhTBT/6HXw1n5H4leSbdBFmfRmbuaBwd/4EzNxKOS8lNV3EsmBL3T
H35XDa86PFlkPoest7Su/V1ZBOP6dBxMqmZHBdk43PbQVZgSmhwGbz1E0jusQ75Y
CJATN//lL4+pDdQNixbOuh7XbWfo1TIUcnjd27rDCRHg0SIvoXI++9h1r2bj68hp
zOKxlfxyiIQJpwdIgCoXvHUDFTHVQjepqr1A+jz2yMQh/BigH3nI9TIHQbtGR8BZ
I63Q9VxUOzqCCjRvxDhws8t0mxZm0ntYO9JNRCoL5D9Mb5r6z1uppYodBTHDz0tz
ukuGnhzxtdc5tqJXmXf02fSsMT02qmQpt4+SaqoDJnvw5KkGJJ9A1W2NQrw0lVpX
vCJ8UUqr/6o5umYCo+ypVByd+g4D+eCu++bV+FmYHi3zvSr+pVMQkXvXS+Iqiqwq
HSOQktWwqUfV+IvvkvuML57oWPY6ig/l9dVn4d4yXAI0SD8irdXzA2LfL6VtbDsQ
ggyPHsWI2R0PVKNbUDtkzJpqmCvp79i2wXUrZV965Q5wjGVoAYLRKQkNVQ0aUo5n
8vHrsgf0oPlYcJpuNAGgPJfNDVjbUogD5zb0yo/hGVdoMS4SVvZSHVxx6zDaLT9Y
/qeL0SV+4/kV3XBSKMOrw2hRYxPaz7bx6KHetdoKe5lAmV/KcKi+fZlA5MWzxbmi
2uNZb7+PxVzVZ9HtLpeApfIc+aq0MG6uHF3IIaxlURKmAU3t955S851naD8ohOdA
sDMlLV5uc+hEhTdQzjXp+ooTVc7N0h/G9lo/ajCSqP5e+xp4ZdkLs6UKcWHF6NuY
JtgtXT8zqsv9DoDLM60Lro6mVoABMXOw+M2rC8U6kYUNjnvfY055KzPMEYlH0b+z
aF5gXfmMYnghCGUcumSgRCQOhBDdkLxIopY1O9O0JGPGedbwR8hX5ysA24EL8KO8
Nyi12jH+V0OhWbEvsyht/QDXOHbkSkuhfh6TbxYkLjBG277vNldtZNFQ747iPRx1
jWMLZqqM0yKal+EiYSItaI6cx+O7yF8O8zgdUh77NvZECXbihJMsruUE64c993TM
qiZcS4DS8M5OWO5djEQ3/wM3sSvs9E7YS8FYW9AYb9hTgkkbtMk5Mwv0yIYT0nGb
wduwA5DjlSfW5uax7qWDOzGIYyKTJcwe48otUt6vNCeS0I4tScJrvqPr1MHR+PyR
rgd1yYNO/KqjlIiQFAU7cjfAAwsS8VpKbon5Uz6XUbboXUssoHbun9YnGXOBKeN5
dV3qezVZvEJzpeS1QriY3/Q5aBY45Ah97Q/eaWY/sE3o6leeM0c01/kaFRD/VJbP
R3jYUJzTiZ+15Pi7pWLHQEL7I9xP6m2FmHy6sQuHlYKiQLe6VNII2SxKa0YCC1Ag
i10aVeWyEyUjPk0DYv4G2CiVjGaF+fEwj79emThe0x1KuWK8yOVWcbGM+hZoi7K3
HIIOHtg9sS2/Ew+ZkOAWrI7Bg+2uHf0nE3eGu3VNRTyfoaBed9L+HOtmbs18f8Y7
AdAM3iIaitWfhu+FVlLnf+TWKXNH/MVxz1+tCuhoH5hRLOGmd/5yc/R9sMfX+gC/
TFtf4kMD3lzzXc/0GwyvBrm/X9FBGBMzbuQ3GD7xmkOKthXdrnCUm/jK3MlKyzCD
+uGxezLTYQMUSmI9+UUHHVQtAlDUp/aHtl7KmNPLAM59FhGphI2QPegHdi26C5pB
Esw5NnedUtxC1/xQaDavsCiDhu3JEYPaGYT/uJVt3mHZr5rEQvc/+K0kaOtLQGb/
iIfPrDYqepI39544+LAFiHaUJ2MSldxVFaoe+/a2UlNMGkYGCWL0HHsDvdTh5u+o
oyVo1QQtizFRIa2cfYFoFLMPR+BRdELtj/QIzIe9u6eZjqGyxNfBPWR9EyH4yMk8
KljMUaKiRDgPp3YkAKyrzBIQEeC/JY22zBjsX9X4FaIubQLvCAlwrRW639EqIaGY
b/wbD0G/wphR4ieKf8V3Ug0PQgImj4t8stfhM9zEhDaHQWlXGJCiTU8gZmUFi414
v77G6KJJARcxRDRxAf3/Ri+VH+kiU49VXDg9RCW0Km5rOtDhbOSic3NJTdJFfgSQ
8d1I60NXLnX6dC3q3iJxuKGl0cPvIayYtXRkMd75RoXMRYqR13EyJq98IedNCJIV
ywkQqI2zh4p34dqrOrujb5os20hECHSq5LQX7EEvdMyw9LpijQdswwACyrHfE27F
BSiCrvc+SduFUcWfFTqrcuWFnCwo8OMykdMKWcNIF+YdMNzqtnCMdrwS9TEaNRRJ
zqoBBeSDpQUwBashEg4fSMjoY+qsCuVyZVgljyjJXWczMOEkzJPDAz8APETGrnR7
ngPYWALESCHxBj74QhENNHrZPs8rMUCwQv3VlYJqDXXoPqfOZjSVfJVFMIbEt+ZA
tg/Y3f8z5o3iRQSPzasat6zlYBzYQTpzRv63elpAR4f4ErWQeidfMbvNMdp3HSYI
5ykky8Il48G5rcevO8V9VJrTQf7FixuxtP4kjh9I3h0zeRQ/qpzj+G4udgnxgoG/
BeevDLiDvdWF8883Js6BMqc9hdzPQBLlzmaaNBZWvSrtwSZWn9Ju5ldcr2hLLIw1
DKrrg/yZ0lqUNj82+kY2oyUaI/9RR4fJQ0FYZs/7T9Ww0g7c2TPcIakzYjMNhiEY
/TbBMF5VpHuu1EM4BdDJYjao/N+0xIINjd3NXplo1fP4xigSJI5r7uqha6PlVT8W
Uhz/wKcWnqDpbLQ8MVINjTV9m22MUMg2sXs02hGF7rWoGtCeQg10+sZGywe75yLD
ivk0V+ergUQNF0p1Uw3WgWmzG23hkmxEUPqkeWtnCFU9Frkk6WZzyfmruuNutG8S
elLrJh+BJEUC7/sBlQvHXNLrJDbWUJtqiagtPgBA7nRAWO1qT5pUq4US81LSzWon
fkg2fjDScXvxKG7UDQDbh9cSCK46aYFRJ9RauQs4p1q0CTSa6yv4HgGMTMR3HOvs
FAlM95VBg09LzX+p4O68yclbSzNzvn5eZ4MkvoN+1fF4HoCBphMtANFiuAGRBAEl
3iyiu0FdUt8bePgXbu1h10iqLDRQVDULOnqXbCV6SagQ08z5a7AonUTDDbUbKPgc
O8GHYTV6q6Qv3T0OyGyzYRHwH967Z3pXZRRsIFJ5O0b+goO+7Fn8Y+NSGuPFvBnV
zAFeVw60wqfiSXt/Y64DPYUY6M85ZgQBJfVe6Yw0qHEQVAYjaC8AnJCOblXj0a9O
0p52yiW2pKisoAr1BlfzimZRidierin3f5zWV6/VT/s2t8lxbCefdTsr5aza/Qg5
fpOzwKC6+SIM/IQ3Ls3YPOlXo8SovrfVdOq6d6O9UXSlC0H5lznDIbhfalVVK3qZ
xaZrD5K+ByRirxyONBHLTCI0ZCSjZF0kLuqcLgtpKHcwZY64UrA3cRte3Z/3rdFa
2Ou8CnTVxvWtEWO26AI06W0mmDQTJqKyynA+BNF1fTM9gpSIgz+armrdn4Rlk2UP
zTj0Twz8yOUbVnKd7g0bfR+mX4NMiRYXAXstZ5+pqD4RZwPMLqLCgDCnWA0wYZKn
NlJYcRuEqj43Iwm/NphxzO7V8PGRxgzbDIrpAys8OTWP73NcouVZ1MTUXoFE2wfW
6rghdBvB6hk9hgIW7/czHvoY2SSqqDWjOQ+xtDc1MCPrR5DfJr1oWfhqDCS66HRb
07zkA3zffe2E/94gU9ScRSLZWh/RyZ4nEJbsad6+KHMVJ+T97gdTrjN6Wd7KpdxF
V9v1VgFphQCSQcwp+cyk6WFORBNsKB9Cf0gIjvqJml+NfY2dE7A8KScp8ua+6uYd
lzOqlw4izzBL7P3Sdpb5zHykLzgX4avzesfOfZ3dNt/rMRcpds9WFRDgw4D4apST
GHCE6a9D0aQspNuUr70tjVkfYdTVAdEAes4PlgfwL5XCIKQS6p4I9n35BkN8ipoy
sgARR9VlUtsCMpW34JzuhTFqJWktehX6+Sg7U4nB2HlVGy8pYdrIZ6HTDfR1o8wV
WgITaMR6svIzS6o8HFrB1rAb/qnIPD5GjgRSWoryoD3CFb9D+w3oegkBojrqhXUn
msBiVblDGlqAfBDxkz7f4Ma5noMnFubNQoIvnP7PLl7Ss0JjS9j9G5ibr5Rd51MP
cp/yQrBI3bur1pa+MhVSxBkXYSl8iKFfQCfqc468h2WkAheECc9ZvnZrY/sXQcQK
pqsopHWLqcHcjSxgiJD1zcih+ff6rxMrGzqrlqsWr3JrODcgS263TdFxpwUp5acw
y1zogwWSw3Dtq1jV9tQ/gUCMF3AfSahcmql3WNHSHAIxIvHUal9RqoG0SLZT1xMz
25edxpRodkjuRGzt3bcL/k6w7P3d8IOm+WN0DaRpP+452E5TTvxoULOi0hw+4GaO
OnlzMboFzve4eMo6aAmuriNOGIcXikbAsuD1T+WsF/c5jE8yPrb1RDn53NCs2Eq2
MDNCcuzQ6eRJXe0XCAxbcHi5A27gCgUWxHK6rEXQu+lXZgNLc9PYbW0LSJzfem3Y
pRkpY0eTpdC8uFw3Utb7MLSUmcFUZIrm2hQc557oIOP6c9P8ZOHZ3WKDsvarg2Rb
tATi+Hru1xHMpiB322kHlpl67yr3KCasLBns1i2ex52KgGSAWhMtftXjbZvZyONQ
jWWyatmJs0BzlIQ8tsOOeGwJmh6WLE9/Bdhe5TLn8h6vU635gk385U90yHeNqdaO
+ZQbm+dN1k8X+9Cz5G9BdmyQSFxAndqXE7hvakP4kFIYZ+R6RgFBuHh1fCo73sDW
awI/WIUku0ne7150IeJ7ETZTgyITAKnev7KQIa4mrt9IUJ6R4/zpHXzvWUCePAgr
SN4qo2jcHf8fLaFNHwHolxgxjGl2mumyIi3CFswoM49ywkn1q54zNZYBzt4i//W6
hjwfC2yn3r55KvFw+u7J/vihmYDpcNaciQ5LV2u53Wmf4hjgi+XgW0NqkHKjXEch
mxCIfRoTA6zTr9JmIn9A+l+3tRRM7SpvByEg7KS4L5dldf7aGInZE2sdkxggs0rl
iE59UtOMcWwp2tih5fI8UGoZ5Mur9lZoDiCkzXM0MtiMNe6D25Tu1V7282vjpGtf
C2s1u+528Rv38FSvHPcm9VBeaSGVFQVfV+S8Zm/R5WfUqnEjSu/BxZ8/3iTN9kUb
fqD8TV17lY8R+5KqrF02OcAfNKMOiqR03vkvaugRp7SnMNfw4mIzm6B8cFmFvdRm
+FtblBtQJA6ECIIQcKesdg4SRwO/Su5aGz8svavf/z7nBFLhVz5GwEPZJ+iQIwk+
3PHDZXlaL2nu5UH2xog+jaxTixx0dto9XsTsIbbq9yL/aZ5q5yHc6Gmr7BacwVPo
dtgZ4X4fymaRhjdOf3WAjL/G4XblbEPFLG1TaZ+n9rfcH+eutmp3fsMDmoDsFJvX
xIYJWXCCHuuJfT8uo1Wbeszr84gMu6Zitru1TDuspifqA2ALZcntzwqqWZjZlRib
fahlFVML7TFJ/fesyLJdRwiS1imk5uw8MuC8TFU1fCuoFEicIMdjxFdBm/d4DGQ9
5Frk6LVahk1j45Guwlljk6ZR3w/qOZvRcHBZ51uwqzYIq5Kn3Zkdepx/SCLSM01A
zDqKUf5gVi3YqSLWKu16ZFzw0DKxRztxjXWQoLfwXfGDCy5GvGAYgEcXVoz4Xusn
qGBDCGEd8W99xRtcE1LIT3R+hGUEW1SjUN92M9NrcOWYljDgA5U7IXaSQE9mbPgr
2JeejAm2NX+QYcVvSQf8tFFYg280RL5riMADeJOHrrSjdDtqhnmbicg4l8wYi0CI
ZtRh+wh+0/dzBJ6xmWdDPNHFXao+yer662S+xPuFxN4JNQckRsK70VwpC04lY02g
Fw/Ipen5qJoCYi8BGQMy6r7Mtrx+0+n5NwB5Juru5Kc/fdPRM+lI4riG5oGG5XMq
XBXCJ32zRbcrSSP/QGumyV/WiXOJ5Jj6ws5P4TR5NI03lWXVRJYpyLVpmOHGWG/z
IfZcL580qm46+ptB72+GTkp4S8NvkAaoMNWeseDh2qXI3TEQ8locaL9wr33qbJqB
H3xykhNi6xGmVA2FkgGWBn+gX+EsgiVUavV12c8rxMRKsycbqKUukw2pm066sNYx
r9b5pZ7En/6tBjUcmDF+t2LNeBccbQkV0WQQrPFsrWtMbNBx8NoboKYKN53hVu5H
iJj6UyPOZjPpjCaiRILPMxWn+21mc/+86deuxqgzkYzwMIFvDuSIoCwYG10nthJ0
pQ3OQoZI00NSkZomTf3xS+8VtXHaapBIoLMUX6hiHO4PLVay0uWePiE1KxEyGksj
XuZIIc94pGF1QMpYa84YYLuxzpde8da4IVDOnpaMgB364UZVi4+MUStwJ2dnBqrC
mf5YIPXlGoaI9QFceRn8BXFEMBbWYy+WEUx61RZW0D8TubnFBYooJMOVEK1mfWx/
iaZ56fXUSfR1X9FYN2Kd/z0R6TlLzMZXYWdJoIpqI+M2Y+BVw+CdRfuDwg2h3GPR
8Yvb04+xXw8oe54PbROl5gxvM8rTn9GSGSp9t88+f+A28f15aqeIK++aMMErnMem
5MoABoh1q0vRceCWC9f2OZGuG1gN5J32KpXucy8IOB3nw9cGkJHsdKA1hOPeXLPL
BqtVT1qgZehr/a8nGyaNSEav5ovB20WGGnRvtjSoJIH2IScD0teljUe6WHNlGvE9
FBvupd6x81Ou31fLxCyXR1bR7U2vXW4hE0rlgoUJLejqJtd7NAaRqOA7zQ90Yd1b
LJf/hyvffmk0sncrh99YmDMwQ2LR52b2AWG2V++jKtofi+u+kzI3kCSkJD1yUj+Z
xfwXCwtcvDkr2yqsSV+MnszAXW0Sb/mnj/c9cAcpQUWz78SrVM0iu1Of/9PmjCxP
vKSXET7cq8q682XnrtdS0BR/t/XbQKyp08ATbN+2gDxOQLZLFW7ZcM5mmodu8nBg
Nar3SsDFK4YsSyglZIhs5318gWdmulrXpuM6D6j5TbSRjQiE4KiyG8+4howODolH
hNxLPUVkTCPMCUlrJSgHS2hKG7g4/Yn+sMQoJuWV/TlnFX/91td2t0uio7/Y8nC+
gLuMxy6klKcrbSC7F69s6TefOPA0f76pUQHx/UQ9yCbRCNguQw/CHdK0RHU0T2Hz
/FSsR0NAInPOJbVqvPrBw+sJjWADFCnFUD33fhNx1mQ/kOQEXWRCo/+W1Vee9GhL
ilhyQlUEUBX7WV9W0NrWEC2B2RfejrFkXtFbhBlNqGLteFh6ekQKsEWbqyqBzWQu
eRE+he4B2aDB6J7LWCtHmALQgcx6AI7EkSF4to5LTk+4VT4gMXMHM+Do0lFD9eF6
YPBmuc/Fsbw15qLrFnANkHITFg3jocSIEdKUBjT7xAidKNTQjQh8V7CmL8yFR5Qw
PmKEG995bSzUFCUJ1viliSQD9Bp1wfUBgsdY038kx4mYA3L646x81KZjJEH7kqCi
GhLpUM6ekyGyTIpW9fde5m6zZGfCOqYpgTO3J5GOpDObrMvzMg/cfOv1o/MP72VV
XYBC2vaTvY7PdwwYLVXi2286iK9uEVVzspsPLnz6K/I1jKhaIh1yrYTi+GXjqZ1t
0mXDKdYm/Qb9tHug/qQguxTIUjjrp2v9vd2KQ6wqO6sow/zEdqraShUQ2cqJvAtU
3irYgRb9sWVhMbSQIy4dikSHa94g93BAvkXzh1yy09fndGo45XP5rWAaXhLsJi3Z
uiRA4EeOLuUfbEMy8/6Q7UjQVA3JzrD166xs1eIVOhs/vAToqDu9IJfTNzFoVnu5
gmfE59cpdysqA0b+1MjDgGTAEGWri1/dhgHOI9qlK6Vm1lz81UerArWKn+PRMehN
g1KGktJvK4gSaGywr0er+2Iyb0D/93w/rThQfaS73d1Cm5FlO+uRf9SxdwcVOpLE
SelCq66tyjxPGbZMRLHcB0OR8z3/GITL+bpk6GLusw3quHEivxvBrtsXLp1CJmi/
yXABegovnk9OnC4IpN6sr5PKEOVKr13hotKKCGzJ5WLuZHCDhH0trzAat9CEc5OZ
CFk/OTDy1SebBApVk3cfCy6d7ID3cR27dvnb/dUVNpW7VGJoqlLnJLWxudZnZNVy
ROudx5iGO0XV9J5ibgxbAJh0xhSDj83FwRvrIFfIYHUjxT15E8WuKAQRycUEa1gk
9nEJamBceSHggHa2+/Qd8wv6NA1zaKlK/poE93RYz/IZwxMwDUi5djTTAvyg/sHz
pPlyG0s65LSCPvBdHhBpID1M7rYMQATgPlyuHCSskWc+bSz5zwo36wYVt/i3M0Kn
8aM3jwSQ6HR6odIljhxMuP17R6fv3dtObFHJbgkmHE7iQQxyJVWuUd247GHi4zBh
qWoLV2qx2dKXjglfhkyxC/oOTDN0CDIhfNlWTgC6pe/jQK3KIg/W1hn000gRD0Nx
22VLwxx9056gG7s7Gx8TaTfP9WkctWJUyzNtGT5br15oLJrDAsi9YvgMSP1f0nOg
TGDrQz5o5FgUH97iYl9OKrh5Uqvz5cXQPZyixegSGxoq+86+D4rA8kmNBvlLPwS5
1+FGtxWQh6eIzOa6OyUe4uQRNJ4fZEOGKAIQKH9tA0vbbu6p0kiVjFT250sjKiBj
sT2rGtWtnTckGsQR5IlivSCSfxi/I21m26u5nNEIkxvIPlSDIAM0HZGvsPYHWpF1
+nXZ0rWpinhpGnblXqfNoWxOfgYkrherafSfqK0YJMrwAoZUOPPbo+lIoGO4V3q5
7KCkkGmN2OL+hNHp/Fz/13NkPd8KNJBGUtm4OXQQm8W0OmdLszXjucitHlmaDONq
ZLKVRAEFWYh0QXCb0hgvWVnPcwuNwYLVJuH5qv3srk6KQLgDOLY/kqWxehgMvpQ4
e3Ci0NwvVcA/Ee8JwoeNLHm+/gOeXytcNo/mbHTJGd9ch28wjuVhiP2yFtHi1UqJ
eNbiJL7jXUSJr/GSDEiOrj6NtAa1ryhD0M6vNEgji50N7dMD7jTXRBGuQpU6QLez
UCyhsyUApu68kr40CI6/p5celxMhTelBYGx7XEswNTff2GSMo77ONhCqpLIrip6r
Y0YuGx/BlEh8+COynllBv7moUX0N3YAErOmHS/+6tb31Pw2r4PV+SToXFiAlBXTe
gL6Lc/3oQMEVn9RdNbp4KUNw3+rHEdRZSaZkvjSLCmVrmKW6ZDQQf6zx0VkGpput
pQEq2dikBbNYC3xm1HsEyp9Pc1sbWytEkyE5U+6HgjusCFwGY7Vu3WCGewo3b+jR
+2D9a9EbX2X+P59wBGJdSgvLgeMxz+OddTScsamDB+p+Yzn4dP2nBDAc970BMGiI
6ARaaDBdq21zaojfSYHyXkicqVxo18sbZVR2vI8+G+/K/BIculK8qoUZan+T/aRd
BW4blVzZyyTv7aSLzgH48+QBpDaCwwwsURBnSbZPJMnwDItm4JDzpZlrcHcvrdga
7VxI1KOWW4gHUNHvgs6QqydvAgptUWE7ee75Z1RtwYH9k16mlvsD+A9XqH44zfXG
3/MoxmXrXhMra+Pk0m2pFNkMz1hW00JMWMlwjWm/XbkISJzU9++nHMnhhBhH1LvW
HPynGeYe/frqGvkG6IE8kWlsxYmNUh6mh+K8N/2pDV7h1IpYSXtfjFpgilMTQT15
6xRZiZyd87PFEIpncHNR+IITJTAWzY8ijXcHkLWJySNFVnOXAnT3A088mKUzGBEc
k51Vg1qgCFxLhth1HzPU/silWbELaKgx5x8St0PHJMTMz+P21eq6JWl0dI2IvUw9
C82BaqsLJvWstVyYreC75TsOwB+1VmMy6u9LDEVIYDAgxl8ORPeGKP0G/9KTNa7w
g+/mLrkEI3IrnAuWNIJDM8bMDu1s8NZ6jpqPqPwcVd+UWuPlzFVmdoBVk37k2zOM
zIpBX1spRBWPJmwROSntHg6HcgeGMldAWdr4JN2LJaqXSD/UdLT3Hc3HqErMicBh
0E1KvKl07ab1o6928ALAucfinTfgqG35M+GP71+M020yyJoCE1w1VgmQUCnZVi4C
sHqOFx73CpBR63KZAjTmSVGwCXu2FpFVF49yXVJJjv/+FSOLDB5CJ79H4Fud6uk1
26BFQoEPT85HfAbD1kfxh8Yp7iQohvhis+f//UhqvLyT5U8woMtUqDjDSy3pe5zP
3hMNL0QT83cdCjtKOZ7T8IltsAy2zgk9tD8N9T8pLHuFvjeWoW4n0PbgIaBuU1pP
7wSXc5DRgCzTiPHOwQ7DjUhJrymIRu51NUJNa8z/ayuCFtc65Cb/CEQBMdrfINcq
uWNlt2E5OuNZbKg/Z/TYk+zl4YWIkssIZ8fv8jnpTNypHu5CYCLysSnQfkjqnyor
XHetFQTyZIpYVPqIPhDEQGa10RlsKpFfKZuZt8Kl7ABuGsDS4TcQEb+NqZJRhq8+
4axNAR2rd+0mGj7Gq3R3pZ7Ac4YgZ3qsVNil2MVfRLKTy3da5BkKlT7spL7sfkxd
Iv2KwdrjIn099IjHJy9wqbs3aYF8KbQ4ntwqLSTeTWy25q3iRmYKD+A0FjuPG9Bx
yxo+E52hJgyWqiB0KFEqljUOaL03c21dkOLeUrdTU+aj2Mjlhevt/LY1BQ0NNa8r
MTLktC8EWOIkiVaFfjRz4aAps7afuZD+jE5zcxkRuP+BgyYGjjeBa1OwyRn2l3gR
rr1duAFMvrto7szQSnI4OHyAQFc+E+Qz84dSuqiwRz87CLlYk7pMQUqGgt3A8Kim
WGepLe/UTtbqzCVI8oNvZKFTkA/KNEt9IyeMjVceltuOuaf4urZ8nLhZcZFROk+i
qn6ZZv8sajdrc0YoflXAwQ1EuMF5csuQT0FctSQRcCP+PQiu09suZAMnaGc2rx0c
qWBa017Xkb9nDkgBVY3Nxnfogi127sDPC27cUUw1QzH1VI7mzgwOpUSUD/jfnTvZ
KutH5QeS3i5NCyt1dhZ25tdM77CYIbWEZx6rqRMG6HznrOZOm4e/XP7HMfTQNlkP
ywUJUMCjeAWEoTP4QK/YQnwKuLY0zPK6+C/CXzmQ5nyrLu6UsPe4EUmCT5SbtSsb
FiFOkOoD7Gdbc1kTutRC+Z1lxX/zQhtu4GIXQAiB3AIsfuzKXW+SRi/bA9sZG5e2
dNq7n7USup6PeaFjpl82yS1hy8n8jKGNhsLRXaoF+PjI5jx3Tpln8KD9K9SWWtZv
500onU7iMbrcCenKUsV/TRWFPdJtHfp5TxjRnISjwtD85BRka5+rFV3UjuPveOkY
+/neqZDc/DxTrLJKxiT22A87o4ayqXN9yAK1PwGr/xBoPn8PLq8TYNOZ5UazwmDy
28AYggr0RAFkFbzj7D7Mee2F/kPeA5ZMfnhNXKnAA4k2s/F31B2rq5CaIK5vw0ek
B4CH31JakfwX9LFw+FEpDo6HViHkyBWLq6HJG1g0j2IH/AZFQcbrhZFq3wRde3cq
J+d74vo7i1JBjqzy0GchoGnSWpJq4f7xAQRa98wDZBJuC7HyyGTJWrbBJDxk67oR
tmqtDJzmVB1y792sLy0ofFmVq+0Cpooy8Q2xV8AfFpMhF42rgdDm8cTS74QyujAX
FMhKM02nFs5E2U6hiMYLJ+MnKtov7yLdkyXFey0GBKKeCRfh2Uq2SeedIGvqSw1E
6ROs+9RtBOEWi+SwFQhk4cf+6t2UqYLHLaAEKHPbt8vN9z3kftCDG4/ojqb2dodN
jTeBH4J0OJjATWW0fRmiK/+VqafzqQDDavE+vLN4upj8eWgdj7TQrlOFIa0K4HUT
EE5ksy/fF4KKPvPGEsZWMYI218eopswnsH4syIj41PIZHd8BKpTJjTnmvNS5EPnR
JRZEMa1uKrvvjvZH3HgBw2YUgvZZv28L4+JtMx5Ephyks025622YFLFO1SutnvrF
9BYVnwiW7kB1NAroJGAFfvjI2jGNJFRq0FtYTMZVKL2yNTRVHejyNF57o4hDrXnD
Ky55ySyvtV+kPQVsmExaEjXZLR1RUikvn+/qrOH9u1pn/5zFunTgdNthzyvWXiGp
Dt8ctfP3TFeSXbLTLGKtxuTah54gsOMnRwMNZjt3PjAgprZNFqOBRC8bWysR4vaL
1bDNb2lT7MaVuUo2KR4X3EOOQvJQYfplPqxGSAoXnETvGS4ENihJ49KqKh5jV+w6
2DVN722g7q4lioehkaJ4CErM2c4wlipNkxHFl736YpposURGtFx76wTyLw41FGYF
9v+p8WR81YKCGN4yKilmkczafNaARQclFdkGnOc/m0MOy6lVJJGI86V8lzWH2wOq
tzE+bHzje0ng4iArrELwv+NxQTF/4DWYx3isoP8jJQgA99e9lZtxC2v9vwa8Ze1f
MxMg3UbxIVX4ALVwVIWjBiXp893lAHGJIu3prC67kW2oTRGl86s6T9rpqp3GxJFW
Ay2p4TkDVciY1HrO8YocsFGQmDej3ly4YR9a4OyQUrpSiv6zTn+11ETbDS6FZ2H3
+rv3tXgUsfJw6NdNMsqiNwPFScULgE3xQt6/3e75D22vAqBJ6cc6e5U2A6wstp5Y
upe+t/Tq0508MJa+LfRr6UaVPtWfkw2iUV7lWI+pV7/nd1/wJ0uDK+ZHIrlSdhMa
TjeJRRdfKAFnsFZBKY4zoZrdM0jHAtorWA/oeghxnFZkxFBm+mJ1G7TFwraidcKZ
nmCDs7VVWnwHCEBEKzO0ihOwUU0DQQBBofNf6Ajt4VTN/RZrE18sx3l5rYP7j/3/
DWP2HGb210sNzePo9I0nvMP4d31IiygamTPLFSE1IynxJz/EHTvR04soEklqUHob
B84CJrsNlVHEbtB4xbpT17ubS1ClVA3GQzsELq+w0FXchVgGC1pxfuxWeNLTKaEQ
pAYmCvHMWjA5sH0s+JwrY/V2/vsb/7vmMIRSAWFgMiVrViFTr43iC8ESSL/XIUER
Lc06cMcKp7143kluR5L+6Jj5lD9L8I7aWSREofAfEwV2InLvxV1IyWABW6qYra9N
ZgMJSpbJfM0K/i8Ii9FoaXlVI8iGNq25D8RwhoSQ+9ao/gM2MBHRnU0RK1CUzmEF
jTwA7HDViCQZbs3g7ALWFZbv2CwdzWzLLZ5lYSoKepYH9Rd+AciJTJ45cD92f2+4
9vgU0ZjNQJhzBmYCCZshN3b0UJiRoVc8pG7txKuM7NhKxe89PTEzyt+HZDUB7VVE
8DQIJf45nWh6TdxFrVfAZNmyp7cmox511hnfbuFhZE0iQ3RxhVOpXb8fwKaeCjcN
v9Mxxw3iFvt1ks8AvxDiFS8yVPpgpOjO7GJcKeXKKz46tM+YCFA1/xQO/orQcpqT
9y3NfZbYf1UXOlyYg5wBHGwzICaGPlTzXCvvt+Mvs8JlpVwRp3i2t8yNrWbwuxz/
pSzV7YTpf6vhn5rpOy5fvL56Ij17bZcel1H7p3CBUXjjYLT3MRvGQIGJXYLlUmXy
iBy+aNmnoSotsH2eBEOt3rRxBLjatIqwnOqYyZHdc+uZFSrRB2ZLorpaUNMy99A8
2HOg4v0HY9xnHzXO/XrKu29jUqoVM7UnCijyOuziRrXRwlzfO7AQKh46vBw4cGhW
gIEenPQtdGockGnyierQrrPaRZ0RWCS6DrNF/3ZSpYY6sX5PyWcOVmYBO8b0Uod7
7tNgXw+krwvqcaKggPcY2MSKVNiQ2X2Jxps62tAiLFQxcLWx9NkL6rIcg0viPCdh
KmButSNRiVqQY4a/wMFYSWA8piHmoU4yL93fOE2xB6jmf67Q82JkOS4gB6+msacE
/mMWvh0ITLxS3OoZ6VGiPtjYoYHkr0jhnVyR3070akI8JmQ5pyVTm9lptJKty6cE
91NDblIPCFRPR1R03qU78eXXNdGETHTMxwWeUprtYm2583sTGkWjN4SpNnaowXa2
gbPfqEFuEX2VhsfjkONprEI/JEu1SjbbwWBPo7p/y+4Ckw1vuGkDUAF4/05fNZ4q
RprF1DakUH1eFiQKQH0Pb/uGXrcICCuIvJY40ZC80fCIXKeVLPLLdom47/Pswt+g
95lT+wmDElKsGsEt/7WE+CAdWjvrnxwly51tPI0PP94+C4JBFGnGTTToGJkzwFIn
NNfZc1lGM+N/Ww16AZqOWhJMbSs+P37d2optf+1YUc5rWElVbFpfTmfNbv2UsUQD
q0mG7SuglboWyeoUmbxP8ue4TbiBCSN3sDGYCLT2uiXABJdgf4AgAKpScxGJ/qON
eegLH1HgpC9yHScIBWzmL/BLQRLKBNzjNybpaOkhhYvIULV2sPNcdU1JG3+n0EXM
TakghYWcaxc99HNg9LBpge8HpJFlnjn+PaDYCsn5gWnTgbZtqqeNHYIDX4br5Y7C
8HGx52QJgvQ1hwoiO1WhLbCiJdrTg8wAM66R6FB3ZICFyao0aO6SeyUiHLrRCS01
ZMJP9DxaVinbDryLo9pPncNATaNef7HCOkLjhnErMMHvW2v4vX6F3uStl98K/LvT
4sBbRYseAmftnhnzdeiyvDpPvwSLXfTVdo9el8qJTJ8tdgOVnch3QxESBK7twZU7
qgWUk0ewd+ZxBizGGGsGC0+FoeleWSrIkKgf8eSKHF8oJXHbcW6T0lAfcbp9ts5d
79W1FiE9L+I2lNFMRe0mu927tO0h0bsXnbjxZf7VxforkXrnyqjXOtS4nRDptW+C
rqsBocffyC+2Ka6FLTgblmczBKNraM9YR1WAonsqFKz/u5I6ur3ETHQNLHehXHrS
UO6x6ZQR1kCjkwMEH4zQfPbdRx57A+wpsokmzEurp217rXFzN4I/Zg96OBy4EwtW
3MLEm3cKX0qrzIVSXcf/q5+LAZwkd8OJajXW0kThYlZvMYrjxDEAjFajo+kumzbv
AWLB9dEDjcj/yK2uGApDEw5Yaz+n4vbkGbu0XdRX9rrITYeD0ffzHQLlHEEPG3K3
zCEg9bxDNuyVzGVQZ+kmUUNEXkiVP/jzD1mxPYUI5sNp9vnjdp5LMj9dkpMTf5nC
Hdq7xkC67qArpQa4Z+D61719ehZ25fUESht8ECpjBlkWSZ1lm3AkAu68vCMmVekU
lp1eIOrsMfFTIABRnsinlpYW/uq/b99Kc6GJcoJmsgHMKoEttS5BqNwEp5+H2XU7
p1xnJDn0jYSwqts1VXtLjebixgMljGKxFlvI1/b2XgckKayAq5dEzbmSd5zcSd7R
jX37po+wrvp16ZD6E4Ci7e5XJVVt4Z7ydptdczvb7Hqj9nx4fw1wlXUaWEqpqfJx
ZSyGLDySsJt52GJhhUdPxavr/EgBoSQvd/I6B81nxyDcoczqU0JgTqP68ZU79aPy
umvqfrdwv7B3m3IYCbef/CXFNTv2Z97sKRMHnkB/MZZuvAMCnOpXBthcBjmrH8Ad
Nx3oKq+sij10fpjH9A4exYaCfuQxBs8XU/taQNVqEaZHnmr42HSbvF4HkrjTMer6
nOpwH1sFs7eDTAAGEyfMlVpZjekYJ1+qUYgG8YjeiCTpww5jPoNuBk1aVrKBY72K
XcCxVy4IhwBHl+ZPBrv5VZ9G7NuK7E9QAh4iYG6AHMI5gH82g1oeggkmX19jIjmF
Kaq7x8oIYtofGhLO+I6H7FIfbpUCY0yyF/lwD1PdifqxB0UUDommMAYjl+LW5h83
aVuASfvx7d6c+Oi8KNlYYNSHdOMgGIkhK/Fh99tNzC3XSnXU2859AR2P0DnLGAGu
R8mfldIyXyfVyCxiTWwU30EI5IrLZ3Sdp6576pAH8RR2Da7jN7X6z6fZZpuip2Pw
/Nw39805RmcaElgW3seDxRM8ixN2SDCZ4k16ccY7QEHe9CoxVB0aMeBzCF7m0ohb
x/1aTHb+dFfu9ecLa7D/xekEKy4j5mnYDYCmA7w48uiiam6pkyH3bjr6BelAftOD
HnAEfBBRy176st0+80FREjjvtxcFUzvnqjvbZe638KA3WLDByxJFg7vtxUuupihl
MDPin0QxR+zR9RWthQ0VGz5NX2aDd4viCrojE5kGlzlmyeblP1uIgjm013mhU27q
j38XXaEgKmDCSn7K3jAmXZvn9yGa0Uu6rC9sgvJK6jqjH6De1gECXzRdSJ0xgWqz
s28hQdUWQWRsWwHS6ddJO5SZ51kyRtHjx7TZvGOjGnTrRTdFoCFCPJ+OcbU9um87
L0/Rg62i7CIfbqIZep5hRM6THB6Jna8oBlz+962986lTmw+S7SOlxXd0O7YrDvbA
Y3hYyaYb2UJkKX8fLTpQPi4wpsqb2ExVKTjztDY14lBQMa1kv/ak0nFbKgApGu9i
5ChVrZEYUPkZDT0KDtP3TivOlb9FzumLGYec82P0sVE1zJX/E6bxf+8CzmRlpMX+
GkVUv1ZpRzmShFsOX/hjHXo1qDejwCfgHIlGXwdmuZLgmzRtJ4H85/kRghqKWz58
gYXNfnjzqZU2jaTd9yqdIXhdvAUVFuqIBPsvmASkLgCJd8m/ngGaB7Xv5v2CZ8hi
Fm+sss5hEgDopxxzUvGaTUrF1NB0R2e4qLvIlqhWZQsgWq7f5NkX5ffUKQ/QsanO
XQreZfCD1Sf+AoBgGP15RE7j+lBN5w70Uc9ly7eDBdwfPSWXwIq2FHMzeHzPWRKA
bUrtGsEY+/xdq0tQO761PLTKUG+cbwP1iN0zWuLQA0DMMAMPDxFuHaQ+uW7beF9H
2fbxKtAIM/ox1yVvHUhpM8uBRh/zNyPc9L7EsyiMNM0lZ6QYrJW137wDHnFEGhAE
w6WYf2ntix/XUh6NSdct/j4qMHyeXxMQ+tBRWDLlaVW+aEAGV8YENbIHdftYg0qA
EKEDg6ZbxFo7cj3N3u/bNJ0Lhv387OpFkVoSNaxK47li/7Px5dgtKExoENgMAnak
IM5Dsxwawo89e6Vd4ydN+pNZJonQXQX8D2LJGQypUMT0JZPF4pMLDa2lxt1bXmZR
XAouqjOefemzzmczmZG5c7vbpC5+c6WUZjM/HggcsRonAq5sVJKKikRxPcPNe2H6
f2sImQIxlWWKR4DfvLJWJlrsqPH7Zso0UOjhy2fXpFspCKD5SnaJMi78NVaZxQJW
46oZ8aF1x+qfoXOQ4hEsIgzgarew2JyYZ49xeFs6u7bnvmLWHFnnBFDAJeXuS6Qv
Al+cgBmvcOAyfl2XEOmMCaDQoWcmRzfb9jrGs0K+ca+DC6YGjz/AnEqWDLMDpxuH
mcaiE1wK0/jw5V8Okhe1mpelW6LsKXuXq5tLzv8kr68yHh7aYa52Sy35qgqr2m7N
NxuZOTg6PLUcF4Z+DODF+pkwaEGCCmBWZRTPKGG2q0GYUnpdV9nEuZNEua7ewDIX
zENW+8SC14L1uzRqX7tq7XGMSe0RMDm+v4885zdoS3yJ+pJUCtAREkOmZeBwz6NX
lVMXCWaRWpe0WttbwI7sq07kPoHg0fbzZQnKkcR2OOLGyxLgyBZWUVBbJjfehlsX
NRMJMBZHYFZIGygkJyxP3K/cjfwrXdAhW0ckDnW+4tPyDG6Ksb+UJQuZyRJUnZ6k
Rd1e70e41LxJ58M3WeKZKwfXEYuk0W6ZExa4wp7y/QcZHJWzMWfhP4VeW807gTyj
JSO7q+Tmi/j02Rkv/G3JKo+NYZlp4gqSSOQ/vbECPNw3ZhrNwQrSA0IjDjxgIplG
Al9Hfa2ERSlFoqyjiS9uL+WWL5FVNlHslmc/t1woSVH1m/HFZrSqqP+2Fpcm88QT
RhzU0ksO1t9/cfDb+kwN2QBQwRkLwo3VI1DaSnS8EpGJ5Ss8dpEjWdPMAO4bELdF
O4wSnvuuiNNhQ7iJHCRkTWIT3UDn+01hq92LugSQBg2LPHdOhy/2jo53nUIkml4u
zn9ejMaVvrN9oIYhoJxEJLTyqo/jvMjdOe8NzdE5sIIQYjdvvj74A2JR07n+EMsY
X+D729uzYELfMu8ocBV5vbCuD2gmroflDp6g/YsJW7QKMo8MF8yL1vGYJRQLcIWI
mz+Az0ZCJF9kpCtn07sZ5eigmwThfIelmzSPUG5EIeJqk7AQSq8GQDprZZ4iwEq0
fY1IK5J3TbgO0R546oVQ2klpqFYTOGHZds/6JuU6gnc7Z6K3P2SLNrlIC/vf1RCi
/EzynuXiGpTEHvMLmB3PO2GoLmsCjlof5djse2BuMa2Lu2Mm3eMgZ82RgIiDK50J
yXSfZ2KJcZtDI4rOXI5hl0O4tBaiTEz7TAJscm6mGrpu2yoyJHnYkWcyHSvfq8BQ
KgbPSdZujRKCfQXxOj96mm2z1qTvxgGB0iI0whpfEhISy1TmKKe7SLsFYWDXTy0Z
JqB8Xn9zL29auAita0pWfbjRwE0biBuSPnj3ZVCPlVLIZdqippigKBdiA0E7b7se
gSBSOVtfwUZXSslOzeQwtsNBvUhRuB/QyVS6s6Gyt6qXHkfZwqSj2ys1a+Lol685
5vjZHYKU9ZnB4bBfhUSylD4cIqRKsnAA2sVH7Iycy1K1tDzRr8uu0Klnh8AuksAS
RaMEtY/wg6oCJzrUXCJz/1+MHoxcktoQUdHTj3FOIw5NtyjbBNGAI6BSnVV7yU8C
51dWbppriPFEcnPizY35JFJZ45c9MmI32kRV9WrzV9GxAkcduNFmCxUKvS4QPMua
thJMVK7QOMhBZOSRMUV2m6kg5BAvsIyoibWsrMSqOXgWhEAzjtarrVZt9QWnh2U/
BoU97rT+xqxj2cZD4x/b4QXPLMSWAAHo6ocbA83g7gBD9ATLohNFN3qvIAHJrRMi
HAxyQOUrAAuJxcWBjFTGtunIn5aJp+n2yBMr0Lptb+9l56DMPL0sc9xDLMgqOV4b
pqdzegiq3bDn7JeRqI64ndv7x3sZuldarMhA/MqbV131vI7wrc8h2TkMv1srY3n+
S0zpFbnUYjmBKHhU+1qMvTXBTGo9MPkB07Yy4D7t9H0H84AndbPfJGgmlyQb6Cz5
a7Skny/w23riX08a1z5Dgsu1FJDmdb7I3EqO5jKqEZeOx/+2i+SlEeBGwbrMAyzw
xHPsfHsGRM1aKaEezTuO2pBKESd4jHAoFhV7t6NIyExuAx19nHARSHc8PLapiyeC
EQV+D9G+etcraegoko7I+/cTZPpFejqWuLzHU3U3HQSEaacWSybP4eXzGk1qSvRB
GHAqLFHncsUKkFNSUBrrFtHExXE/mkZMCxoE8YG1FScHbw7XZQIUyepoJnlslqnH
saJ+xrt9QMoQZGXMaUihxoBrNGUGzdTlsSa8SnIOr8aCfn54BjBOUQuMC2RY//Lw
LC3btH5P1Ly0v+GERKY0mPHUQUwUAITmf9qhzueThzFo4XQxNyMb1jFWVy0OpTRU
oC2yllkRmrEM1q/Cr03UYJ55HjphX1FmM0VzXi+7zlWUPGsxuU4mAq/Es29J25tb
U05zdIJd3GmE4o91Dg0X2zxbwnf9fwCbbwfDOfqKAcJhZyJ1A3iu7v4fA2XbHGaJ
nq5DnDcK7Qo4KZKzn7mPMhJIr0KB6at0SfSUfJ904O+P9mTwNt82u5L+hQhvUZPR
0D6GWYa3rXWnu3Jg/P+zb+OPFVTUxz6CweZ+aiotUbh5Thq6OyTeSEgW+dKrjODE
4anjNq4Yv7XQJz2pQNsm0Z6AAVm2R8ut9LZstpEWF5scAwCxS824HbFENl7Ibzn8
KpBkbCDOukFga7K5OJ4k5Dado2WLSNB66a4Y62+0gl/ufoW70U0Gq1Gv4TmhF0SO
NZYLPrYKKtl1/VmtxSiZv/t5w+rswxz3rT5wTxZGnmks7evrA5/odxhqSj7rn6rd
zDbFCqjPJ9boq1D09t38wr3zqcZdwlG+pnr1lbEs7nfDiYuTNLdBwtGNW1ja3E90
wQbZO4QJJADR4Htusl82FjiJ4YsPCYpb7VXXW369WJWbwvE5suAKPiBkOK9qrK/H
FLIX+J7zBYFpY+ZmXM4+42MQxh8CCHMNmi6qxbNLh3dxs4vT1CtxUsEjqKeYql3H
J/VBOIYS0wpLyRhpjMq1z9rD0vmqeQ3YTPjFh8/ODUAJBrDx3G+DMvrdUVGem8Y9
QArRTRFEpBlNg3W31r5MLTtUUjei3yIRkfrQVhjXgdOc05e1jhi2zL07tB65j5C9
WGr9EFX9WRWO1W5IJ6d5XET+NxVVV4l0q8b4BNJ0DrrQYeSki0DXUeE++HL7QILl
TA+0Qcq5iIxcc62aRLkNTGYRaHWcI9LB8eZQWAkbDLWaM52kvLp21E6m6/fbdjq8
w3gkIELTmj1sq87NQAI8laErEP1C0sAa3eMHTiWGI4YaUbgczcnXSl9o6h3lsUXp
Vm3/E+5rfydEtRn3gOda8RwU9U345yTcUe3JwIwUq7MW4RrgwoPwpRuFvwvGjSe9
32B24i2vIWdofNGNnp5INyrhoZUzvLPTkvuGFiMSrzylSeokhHWxhdTgNMvfCB1z
rUbXswQcWs6DHabuO6e3jI6zjchT3Guv4/GG5x3PlEnbv5cObMq+L0gUfsvRmOec
9ByuPc2xvqP9GK3SIJNL9004I3AVDC7v0uuUNuP88V073YXYbuOBAPSjffKmzqO3
YCZrjMibypAR2Fq0cl+lXIaEG2Xe320OkBYW30cZhPNzYPQKpjNcSC3gdw7WEwGo
9HE1uGgPbcKLJ5YgnCSyp+3BMO3GwTpOg/28gomaIMp8rfrePzUZTX4AcAqDfAmw
A5+8qDdjuIY5Imyf9mDN3ASHb4aJclHRVXunWGAKQZ45XyHV/4hsMEUiYjhBo1h+
FcO9otXo90v6LAsIIfr2gQExbJF2NCQkyIcn3JbtLdzK+YzP/Al4mDcB3mvemODs
B3A4UpBDoKZ1ff4ZJviTZdJNyOWDLWyWsTEeO7U9G9t6CAcg5itryFdqdYYSin1q
r0ds3vwJnTZ8AcXHGgx1FkamZeHE+QMrbjk3T6QgQ5S0hFUiG0RDiFpXyKUvKJ7t
iR1tZEzuIPjL6Umqdjmx1MmCVjhKm+ycAUuHsZtxHa+qehhRkhLj1aUJ0ITTwCb4
gPQTVLqk3vBLrsV2EyyaGeM9cYravhW/PU083rsKjE9yX10fJrywiDYvVXh7NWOb
jS47qy83OpseYwpfGSEokNeo7cFcWEvef21aaEFKLMMqNv7i8Zvo4nDPC3T2UIFk
QdCMPidzmvyuZL53WThUZKpaPEJRq+DzfMfehCxHZ25tZUYo7t0nkCj45f/sy3oa
UBp9rsLIBrbsPsphTKq1FCPeszGbegaKPVgwP4a4u+eGJr0Lp3momUhaKRSLD6yo
rnjormDIVJjno1ioUH6P4OlrvsDSxML2985Shznra3/ZKX4pOqNhx3ZL+2PS334q
eskjbXvBxDC5L7dyBU0Eoo5ThdNcwR/6xWqA4pyaZtnDk2N33PTzL7CswAv2wick
JkbE8FI57q7Yn+0Ra7JdG3FxMGHj4ocCn+qz297ESVZHFTR667McrvdFcco39CTQ
AUZLz317e4JtyIFfRdwMmMwms7O2dz+jLhp+Js4zxI/G4ybpVjwK7BdShqh3oE4E
RRGkrGXCx1mnYKfNaIOALH1IB8B0WbV//b8jOvJaEXkrAeOk1MjmazTuf4gVN9Wg
SB32DXLhaQlrqSxjO9Bah3utNa+vpvnmuH7/pJHBPqy/z4gZQSEpwbrx/rloSK0P
NrgMyowByVUR99cydDMVuQDVKqfVjQC+JUN967v3TpdM9MkAMgmc/8MRifd9tAWv
0O3snECn89CrumROh5fs4glZU52T0oZp+tVRid9vN/g/e6seF/NBCOLLaFZvDaq0
AXLiyY7/+uTN9CPjscDUwpUHWwWtyTkEP1n3U/iMf4sfl+b4Fh86llYGWiJKOk0b
nnWhlG0G/fRSlCxbQ+dtIsa4lvYRXzbZgSwNRo4dfRqrQ0I4LrrBYiVzEZdoXGGk
SuMTR2Ele+3l+KSOEGWGsYPI8BTSjgzCw1U/e5mbHlEQE1vUaLwJzpRVbEPH6LGa
B1SnGkBBneELMNrO85NEzrPjGjzRdTFPG1ctqCmU9q331N5uyaQqZ7Pu1k+630br
v6TaXtqGHs9ZTRC0WHtTwHEtCAcZE7qSXf33Ww2tYr0rILmJ8ABDrLv7B5/if5y+
Sod9fD4lQ9Zbo5DV0bD/j1R1vEEXXOYfdSQm3IMIXdo0weKt0nnxgP5/qiWiSuc+
TZO4zOCejm9zQG38L9qSMwM/x/aJMWhk1Ltj+bbg2uGHCspTYCBvHb4zYcNqB/g8
ksdkpLqyx4KMUqU8gYe2jGBb0E3dD2q719zHLQqGt3q2M74WYl2Y2Dz/5rNrm77w
plsazMLIhw/Z/TnjoDNQX4ItVoGsY5j0b8+4DCYe6/E1Xd7FRNw4UMSYwFz9bgYT
zdFtQ1G7ngm2owQmeUMD1S8YBUlGL79CKMF4uAZiYBwHQHkAU1gRFdaY8ALaNC8v
aps5byuzXLSAVJQ0gE/Zk4Jv4wBELZHHR0AH3NoiEglgKWtPResyRaDLHqduMkVE
pIIQoZDpkEynz0Z6lxaU2QOBx5z+uf2uSLDXWdPV5Wj/5nki9+P62Pb8nkgW/Wrq
8kdA39Preexyl6G3kuAniwcfTSvQx0o4QUiHmBAN8xgoQfEOQsEJEIhWOUQU4QT4
ako95F0oWB6nfSQW6U6VPaqvGGHeqAY9L0uQOqbFnd6zdF8YJwZ8ncHWZ9Wv5LRj
rLVvO9amPN1LTR/Kz3Y+ElML2ghtCVRuWY7vIlpxhNjalG9eocn5SM4MIF5zBbNo
QpMG+t0RR3gzybnJGKfeoswTMJa1xswOc5PC5a5PFfmpaYFXE0smfmgLhY9ftalv
MBNAiV09MooYmC9Jy9VKZ8J60LpccUasjBdEWLlnn8r/ECJTx/06QT20t9O1GxsO
swYx3tADuUwax6IsKcXw76VKZ3rUa+klN5I3cxIPgH0b+MnBASgBUVY095/MfJrB
E45E8T+qE+S2sAZTkzreCQSyrOnsy0r1IriQmnep+Q5AswDKMgYGDFtf4VkDGISO
8VI+Lf5yOrnCkaLKCYb1wFfNpT17NbNnWbXsDcANJ/wd+dwHU64EjdyG+/PTiTkK
fjuN6e6mFyhQcj+TXAJ3IIyO0MKgFPvR8GnZxpv1dzbvhQBbJ7kIGT8TFCQYWsa/
aJj4BONWg7NwfDXLc2RSYhfgWXyOEUeyk+OxSoooT1p6GWfe1+Ar8kMKWM8sO5MO
yZ73DpH48484pro7KBR7UMK3Wb6H3xGW/W4WPuqfADlNcJYb98eZ1y7Rqa9aBI3J
CUOKYOgQMVblmUz7d1OTh/kuF2Ee8cUORq8MKWhKA75sjju9ze1g1Fj+mGwaQsFi
kmiMe+dbr4X8JRCVT2vXJaaFQhBKunjggoeZ7NFlabmJKHP4S3+KN2+SqwxezTeo
ihXZ/RWQ3juPDlUP3LVe2InBnp4bhzsB34nRvqD7V9++iF7SKKrDEmqBhWVagx7N
qnd958kVeTXVXPTj5cNE6LLMmfVWf5w4CKKkBWDjoxgHzBfrPapSIAziAdUc+D2z
BaBbuGhTTDdyW9Q6pWu0ufsITnkq9VeDK5kNHaBycWSUiyO2FqIjnq3J9GnoCofI
JZLV1ZrkxFUAKML9NbFKh7B09Q5cUXAag/vONFo8I/EGk1IgUUBl3uslZRRb3c29
ayZiKOgDe/6y3DZD7CYVf2vLPeaLf7lhiQAP0Ngp3EwZD/HNi7058VRtHjFSYrtx
pX8Ju7iGz0GtiHcUxuiSFpD5BlqiSAkKzmYsZlRpTd+glo7F/q8vt0QdfU16C+fL
Rq+VxhzbhEHf9NqzyXEw+lRGLEeTS31g18HpPzjawyIHNFwNgqJ5SPvZURNAR40g
vo6EsVDmHj0g2qhfYzNn3HcPzcwLDVY6kl2iHXvKpUXV6Jgo/sATRVsPtkKV9Crv
qRGcrFaxheUOVsvvRf+PH5VQhPRBTAu6fiys/Q2h7JQqXraYPG46CZD7P/KgZd24
05XMmzWEi+xVHignHP2R7iWTOiu5rLXPfGGMIdt+UGBiuS3yPhRKYXHXllyVv6yZ
P0GjF0jYrvJZOEUjTFkVASE5I0TBWRHcAewurHZR8GMM3zmbLTJnIdBtUuxSSQp0
Y2VtdJ3LhS472e5iEpiB2+dQLc0CLmH3MuAIUzDSYaCkBmVsPSt8fqa0cztFKzdf
5cPU1n1gZGPj7IeIhfI/L2J3DoUCBVnkzExpIGKYibn4DvbuOzOWuBnO+9H+veND
MpCvOxvJZJ2hIB4WYfysY7LhA+lUztgO2OxBgsmtNYV9eiaQRMmefMBhr/rehcd7
S/o319m4kvaDOWDoJpMMyGuuisAy/uF029BrMB64404XwNW+Kb7QwZoZvikjJixR
k5OzhdfJD+68+zMZiOun/VZzQ7WLjewa1jo6tCyhVxdsGC5XKNpkHgS8AdB5XBsQ
zdVT43zcv863IOFYG5r27hgP1W+2egYGloFJppcNmfkl17mmI6BLihnD5VFFvjKj
kxDzNIIpDpFE2FWam/GkZuFy0oCEvRDV+YTDdNRyOdPXqykD7SharcTDjIEnaRAj
cFeVEBJNaFDz+qZjS3KtZrSwSKt1EXVQZ8TqkFOcICxIQKX8pLcJxLKRErixhnPy
onMhgjRuJJa8uvSQ/DXV0lasfhY+J9+EzXACF/BvSmYLgfneWFedkL09az7wHOVr
nhffpdIpFSVMZb7F6AAty79v2fdjuTy0jr8vc0VIH2zHlU8wf/AWLz6ndXarPFBD
8NfW4Oj2zeQftQmX9f6qpcQDMcR5H2nYpFnmIhuN9pLuF6nfotaaKVFtQG42N1PG
e3ohSuP9ohADmRD9qYC0oFwKam8SDx0eodrFVw4QEeQlUhaIcoIpTZ3My6hxp2Hv
9XyR2tOjphwijRWnPHfbk05I+UwZdosfTnqF25MnhButaVJbPM0dlGnh0znwNjDQ
sr/urH/6Y455mNP4ZBJNsHoukfbm9MjRC0DefyaPxR1wPl4E9ugM8eb4OJdUIV2b
xRTJUy+hhgmT6HOLEROFjjXIZf/QxIDZkqUmDhRkqMvtiUuZbn6aSc+xL5Uy+Rj6
8NHEcKHV6vgy/iJIwYvazyJyjHV+bRzSUz97OJAJrJ/lpzNzAcxSN34xPsvoo7BX
vokmkVrXuDDkYPIImyk0/QSspMThLQgo8Qhpod4WXJP7a2gljgvCymUdTC9xXnE9
zb+unVyXU9Rv+po7K3gZeuNr5qw03YByY6/5Vqj0q/mtIYZzFdDGHsoxyy6PUDOA
iKJV34EmlW+yKwnemHLTWIj/YteyVudWyzwRsMmvcMqn4t+sgRK2UHNxpCg+VQed
bG7U6KiT1lZ22GmOVIu5nfDZg426Hp4v9Bv4cx0L3MRK42Ohz6h5CrqTEGhEU18T
2fLNpeHJhJTaNxIhUGJC9ZnW6UQlZlbQrfqBfI0QHmgdh7SY/39XHWPnQdi8PGu6
dj40qaPwhmhhBEKwu2BRMGR64q7jAQkgCn8NU68GGrkILOEVTfpxwE+8adEc8kG0
KNgiKp+5Rj2if5kOPdgoIoc7d+Dv9CKS7giW9A9HXC4G5vFgRd4dvfua4ZkdV9Hr
THJBIgxcNtj3QYqLKv4vXioloeVlw7DUs21b5ENMZhzl1oz2ey2bl1n/NliB6cbh
eujH4FJe66q66iQ93zrzsoqew7kjAGXagrVG978StzrTyWbEEfq3ujUJ52WRS4mC
4of5v0imTa4pdnNq9h5j1EOONsmwQw+u5N9YSDirvmrpsx+DYngj9QpMWgIw9y3+
P60yzolXdeMqzlcZAmSh1VeRMB0/JFjNEXoH9tCRavfMdhMUbsQyHyNo4qp0/CW/
EANNRg+yU4OrmtcCEVGpe/VcU+e6rVbLdsNuuT6bk7zoo2KX9PjhGY7VxHIdHa6Z
bUwnY45KAfJfERUyasg8wJBC/WU8copuHoEBgHXptQhj8NS+LzwWYZ8fznQWtUj4
VI5L0D0jFKisWxy1ZkXWrg+48FWRlP2SPWUNiu/eFw31D3TWTkXwS5OPPEjK83ZX
H696g5AsbJN7GqbEo/3hnu3YQcD2eKanTb9g2DtFnDVmFHqppRN3BZJ/So0WYOht
IUThLVJsHPlq7bDcgmGw1YHOlRiqyZpOgZDtFDLrNovt4jaqD2AEArozPhDP7b3Y
tSD6DVUpGvx7KigyUYtoZSJ3nMuBrwJpwiRuKtZdWBvAbJASR/RYC1LL6Q3oYYS9
5pSX6tZpRuMdVwxmr7bI70tHFMVibwT4Do8+vAFGk0BykqmvlPsz13tcbKqUa8y9
PNWHT5C2H+vfGm7qCAjq9NnY4TU4Njbq9GRZe7WJ9pURMeBCaxudAgxCDqoGtDea
KtHI3WfsmXXmIvFsQ4DYG2Znvrp6QcFkP/5DdkgHaKpM9+xZzwCt4plgI3XaT3qv
SxcACmKhunwpeQ3B3NMg7h1kmdHXaop6wVh6AzwC8K8wD6IzY9aBr2BUQxekL35O
vBPoUq30ZCMNlrUKiOA47Tp4uNtoPsFpAmwiohd/sx3G5zcV0KXeb8RuNfAkyyg8
pBsFPSizrmTx/230c7wiD8ubWFjiMWrf+XHHblNe3H/yftQXSn64S9bZ30Y9Ucuz
HRd0FKUfXMpQyl+TDit0sipWljIekxsNvUtNxnqPcdwxQ+iHB13EottJ93XLkQfq
mFAVmaJ0biyMy6ALQgjDqtDaOWu0mcaKKvI1jreQyQiwcsDyYjyAxxnBA9ZJiVYk
V29ewn8kP8GRoh5rs+SjgkimuPQTDLP84VHTElbvLVflV4TvkssGG6lqVMXWSa79
K1znm+CN5QcOBj8lBR8Aqbxe5Q3MpAar5a0ggAhaElOfpshSVzUNlcwx9WDAAMJn
OUk6gX7qiqHtQyKhwEGiIkPqEhQoh8h+cIsd1GebmYHi+KciGhqEl4E1/F/TQ0Us
3XqlNWPnCCYpsu907QyBrukbUmNFp4RjFscEwt/sTcxuMlhD41oJr6ZAZpU0ct9v
GsxqllYdbiQFc2KbrQ/jCt5Faieh1ktCujlUWBvm68ndHW6HT5X1qCi9Bh1E4Phl
zOjphwa55dj33+Ir0e78KecpFyTUWHqQ+ftG4BWTiB19G4hQV2U9ZvwI8Ze356i/
5xgmCTu7gaQ3bCFSVP2OKGlseI0+ZdP+rzSMcxeKENxVFCZKnoceTa19bT4mMoKu
HCEPuvk+IcbN/T78EhQRGzDYAY4GDuBBZflaLRxIZGEAiB+lUcezokODjf6wuW4q
uzOX/6pIYqL6SN6J7TTmQE/GJV+uj8UBaVfhFrRyQto01Hre5WbJQbhcEsZOrdzE
/NNtzJXwaSUqS4SZ3pT7Qrt+4YLxgsoWcansM5ukRwJuEsApuLy52SfRAlv5kw+0
yj1SyOlQR3IG4vNBSJhz9eaijrWYjjhNlqEVzHJuzswAqPBriSk6D156AHOUargh
7QI1u46DUGEsim/9rDoy8pfKqludK5hInyYetXH2DJbqhaBvwhJilStKHEIjQHZ6
G7Qqaxf2MOJTqu1ROARN7d+ZJaoqwAoG2Yc9PFiSBIMUkzSrjkkrCH4DoE4hMZTS
Yuug6g+JZiPRYd1EzW2IiZXiFSAglQGDY3QCzK0oPjZN8U9rpXSL7G1NjiXmiAIN
3qC6D5NWVDNsw/827B+1udhuONQBAUvPM+Xat+MYchqMbcpVUx5Ll4Yy/GKdx+eH
G8Y4vONivy2Bw4gdWZTFR02ae8amxb3IGFCWgm2eUP/IaOR12k0VdkiiT7pwSN+5
oXLKMMPcJzDZXSJHLh5tDLW85ptrNnwWVZ+65QFa59QW19ks8ZU8jJZqYlXOc392
Mnt+npAoBuGZe4KnhF7/asVv7NhWEumwQaBjcOSNcPbRcg7Sb4bve9qPDq3SSc3R
eQTGKQFcWsgRuKwNtL9bkwPzCRKzjpLi+cypANQlGZSY1sQ51Z8TL7n/nBEAMmPi
DrHjTIJtr3AUM6xU5svEC9iVq5+Q1Mhlk9gkuo89av0uIFwXas1sBTJPURHgydbB
MMnDyNj/mlSoN5lr2u+NBJR5Oqd1DvSjxCVEtnwrZCXg/4/GSrQNx9sUcrXDUdRL
vtgtpcMuWbZTPTjXsOZGGYDLJM3OCxOnhbI0reu6EBzmfMMtCg8RDZK5IED4kIc4
OnUOkgXrAz3zrDQGkzld8ZY2PUdvlDzrahLs1S8x+nsD1SYrSIFz9PXk4mxOz7N/
vM6aMrGtOQ2B7UJlb1JbUm46iVPE0e/4TrqIjCwyOHpELBK++6K2KYJZp9ErL4qG
bWxmVSD1qWMqytQHedQLeR2IvovUKLNPLUofElFKkChXA7x7wdbLA0cdYniJDjKe
BIwkbUh45mHhWLKbLCtahE1goeBpLNkrqztrLCUinYI4Jv2AX4N+2OSXC57g45k7
tUYHQs9bu9vFb4ftc5IuYkYTw1VRJ1yrTfZDoPK7TDzQ/MYnjYzAyK08hwD17a6T
wlIwB21CLeP4szNMcnv8q3k2MyPkX6mkV1XIaKm+BsKBg784AP+dW5OxVOOLiNZx
MUz2KVdIZ38GiinrRaAvW952MpNtZ3nH1o8Ng6iQ1UqyX0XfFs3Yn78e4Hs/UFrr
0pML67w9q0cIQpYOFVNfcodukpjnOHfQPR2HByaUvNixqj5MxUIL7hv5K2Szs3pP
AxACxeCjrYTroO91Au26L+nB1UwOl6NXVe6G7qk/xgDMdBAbJsgrOwZfSPhTrqLI
WbE0igImBMfvPPCALGUhQ+JGcHn/CwMM4pj428lG6tP41YZuArJ3EDpUqXhn+mw5
boQmMY9E81RIDzDEajqM6JS/lIKJmZTWRTCdGiQDnLiluFh5/4BcUg3Ug7wat9yl
EmFgnm0Qf/SJcECwRSjDAXG6YsyLya2u4WK66N7Zy6O/NUWi71eW8+0BalIQL2KU
ZCeGoPr50HnS9c29X+ZjRQavJ+aQp3mnxlb5VZRdaOD6kIJZZ0m0xTDCqqxxblxz
UHqrFBtIPOMZT/FLqZZLDlr2LPRiK+PJF7jxWIt1t6M4HhBmo1XP11xXt7fCX52s
6dnhWxKW39ez5h0ZTjckC7O52ZxcUttTe6v1k2tjut1HD/wsYyMh2GfeuoRrUx8M
aidAY5DrUrV9rF3H5/osUHl7EYju8PTmOsWeaTTesNzuAG30ybHgxW6YuUeIX5qe
SDA5tc1zuj+uphdufzG2kBI5HtIChYJiqxjuXUCnBLoePfOGi1o3zuB+Gkt2BnSF
N60MoCMWgq4zAwdCMVcqjQ==
`pragma protect end_protected
