// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UjDcuo+vPcQFxdXL1TvOUx8ZgYlWzMLrDwxOSWdrKW81MPMXJr2J7uGsxgDU5pAp
XXmd8SVU9LOx6U3rEMw172KEUUl/vDsn6h3uRRwuddbQyCdGX3uac4lPuu0cIObE
hix3dokBKLxk31u/Gve8awJA6jEfjs65wULaSlWbDjw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8720)
Cyq6yxQm3JNy/+rKJWiJjGfpxp4azy5KioueQoVEEj3WX0VWMrhGsd+HYe7THgn3
quHiw/sjXEqHdbI/4MssQ/y7zt7Q/90QUTVVk6/zm5pg5F3DOEmkxI71B58ZfOVz
BouL6G2bYk3hDPHUcACLRMaLg4+2tXx/iAKH5HdujiGFwLKv59RBQdaFJUlaXN6+
NeihQg9Rc7V27huEFP6I0R3BW11t8ap3Qdx7/5EoXT3KVboX4TvB8FcWui+JKOj4
H1V5M2l+2Ceb43acsexwqNqp126JNE9YJJEZsl7orSuN8YS7TuroblJ9sqnxsqpQ
ptsqQ/lXdlo1BRJQIrSdgHDexpIUBL6L1pt/xsYXYiblX3yQvMlObJVLEGoTwLmX
GRMcvqcmRssnRDJeZgk2bfYO+owvdw6I3WuWys/5H0vp5IDPUHaahFHzjFIuk02p
lEjbKtJ4UBAc6HmG3ChTjihyjImVNKT5fVkFo1X3ozj10VhvOu38g3Cljq5VGDxh
ICNvPipE55DZ4xHAXU8Bun2kTTeFdIRZ5sgVB+g54XAHR4GrOu1OeICStFs1qjyQ
aUglmPW/lii1b0CnC97KHUNpyAKhAOkAmWxP/JwrdaBE/jsS1Ah8XxPiUEpYG7aQ
9SNfC2pEe9KMcoZeQZQxMsW4DVfznSZmmfWf8SYSuTDch9CV49seD1lnajwv97BX
kiDF+sJHZE/5QQdz88C0FrPFQNOyflGAaqeJ+FQ4hiKeeIYAPaGsPEwcxmq524gE
32Dtm8NIhvDOs5J4yLKAv7HvsMc+P/oSvh4VZPLtl8InzeCdYjfhO+2Weaa9zhgi
eE6T98fgT/E5lRxyfdCNpa2ynolwXftWAiQAF1smwmPX6vzYgeuykUntrm0yVOKo
cXbJ9ljxgMPrzCJ1T91tqHREQpuQe6lkz7+aEXxTodAK+eeqSz1Swi7Fcye8vvrg
huxqbsjFYjVPdkJ63jCoB5zeJVLA23qTllddlM2i8PE5eKPTn+1Sxd2UtOQf3+GG
yQcTN0XaTTP4NLHuMSB6bOgS6+u4zZLyXraUvSSYPNVB7r1cnITYnavVj3Lo8StW
bck47HbSAq9mOITzF5wXEAyTQrgOKY3+FK366CCgbIh9W3kH2JUARQGMYPIgjF7U
hTKyvBpa3MmPJAG3bfb+bGCbmENQwzJbTaEFZxX6ah1nxeT56gM9nmnHwUIcuUlo
oNUT3IZqnd75SAV67u5ULg+96uHynFM3dAO6hdko0TWsWZh2bT8+/Q5Bjx46m7Qq
oV0gKtmOQaLReitVjZc2YTxxbNEjqYBm534G5knxwJcqTCzqa/kdC3w7Gmmf1lRE
B50EI8hwoJrTw1tY7xwEzDP0iAwa6w5AJ2FepX3wVvRVajUBzRWrTrBRPVV1NI0k
xJAGrsmIcchDpnP/A3FAGMivBRDLGHR5xbeJq7OZ7TUI/EV0W3vrBTfA2Hd94FGj
+cMeflT4dgL0yZYyEWS9mYeDg1qTEKifJxXWp8ZsQf8TCzIGj1scbdWFkayx/IjT
ylUJgZ5gU2BSGEKaGJmvuhC+xNCHjzGNMGMK778titgaE9TowWoOmCyk2avySCVL
wzG2Yj/jOJnAz8m9aars/MdB86p3CwnkZmuCQzQA8XQC4+yHSTCXaSoAWtrLd8Td
3fK63mI+0VG7i01YZBF8VrSccnNwzHRLr8EzWlUFcJJ53VS6URU+au310I0dNmT4
1KM/zU2CsVfBqrIDoSHH7tEY2tvsvHqYY3wrAk2YXEUTbSQqo8QW7XUvd8ypQ5O8
whiLCYwik+d0rRlBFHZa4PDb5dxPcpmoOq7sbkXhk2MF9E8XJiwfj0TXJupW7l01
0dh8GbhZJU/REi0z9gq30wqMIzvu1IDQ6UFUzywGR82TjnScNqCuwSMY8+VB2VXu
KXFvH/w2wwIOUE6ZlaHh7cevQO+cYtlN/UOmUJaNw35xhOaZzu2qG+TbWRw/qffw
fRiO0O2uFyco6I1pCVSv0i78Mbt5PgaHlJysK9gPAFhH1I27/hkKTpO9JaKPUgP4
gb08ze+ruM16HaMHwjG1xkLQ9JOosuAIHTKTwCM43OqNik+ddmVem/qTuARd4fyo
7p3Y/Rd3bS8VxwFnHbroSu+ZQf4UxZgSy2tvvaBEraZKdWCIdGNwdzJ0hjc1o0FN
POD0uznxt8nzMr4ZYpoLRsQQzQ2e2Qfraq+1T24sGyhdWU60nayvVFQjZnvMnsYV
D117IDfGZvxjIah0UV+rFBEAgHnonjKqJaN6h3Z3usNDJhlySK4lvwL+SH5nxvHZ
FLlVLKPMwTfLpNdDRHJ6mareIVQVyVdRUieOW1mvCAG+sCU00icRXRgz1SpSVZ6l
kVq9WI0/hUkXA1mNi2YShgQsk6OQmDaMuAU6SvuAGNSk68CeoROKbmRvA7lboDZM
OG47EqJA8eyaUGRQqUfq1E1NJwMPB9PhgcwYwiQjYAWJ0rvIT5UASiC96kCgb8i4
S42hJRdE4AcTcg9I68iKBvMQLZjiSKSQUxJs6ku0MF5LZia3OgFcSY9olbjaJhpZ
Y1Z+zzNWKuShJmkMXgH3En8C3rfE1s4GM9bYLgXfThTKuvCgA3yNdrtRQei2hy2e
TdK+TE6jZo+aYtb6ogrmjInMyfFlwizX+bi8sh3jLs3aqOXFLuK6hmR8Yb8P7G4R
0hZ7xX7geAn4pK4K7gfYurjO0CfB4DwMleoOvLAS0gZAqIhOXCtGPf7bUOa0pzfb
5B4zxlH3u0i8JOEg6edDElVC1UGzx+GzjFZSb5ER75Bm3TQLTOjvLHxR/myYJwH+
sdcKJ05JNb76Tl41JLk0TuMgnHeEuHtmDU4X+817O/xykdQYXSy7xrdVX7cGuC6M
PAKVVKBkrtmXFR5M3ZpkBmLwluzPlF7rzqOnlX1WbQD6njtpiqVikmg+LfPNdHY7
tG1xbtgqYMBLIw26z4dJPca1y6GoENoZsAmRy/5jfwu89nEk8vd55d29Yw/hJQ/7
wl3HaZ2SgtnJ3iL3IG+SpQsLLlBbgX2DmNapZjZkzGIW5oBW2YNmK+oUeFBozp1L
QAQxVpNOEMKgw+XXkCkG7ztRYCKjRnHwkAM1D1L/UIrC2p5ZSY4q8OWxgIYUS9qO
fDEhy7RXoGuyIM0VQESo+GLfhxF3xjDdgF+MIduWqEAU7Oua7MEn2sb5LJy4MO36
ZiZQX6teY2fv5nbaJCszjVghDHTif3jUB5TfdV5EK7n20juZsVOFNJt6Y2gmKbbK
yPrQQQ2li4EFh8GkAu59Ku/WeHLYeL7h9ocqw07bPdD4ylqqw6tyidAJkfLJgkcX
qcJJgyuh1YXB62v2/z3sQWCRs8SoIa4joshd5QVspkivqi9AORcc85fyRoc0wjb7
FfPplvSdLBv2sanONpV/B1/B7TSLxAHS3S5o08hiJyxQYgUrgulrYhFZoabqDETw
2jJSQcccAmQya1qXyK/Pi84OoXkmDqR0WUQ1V39Tpnbi0w+yVvaSSnMIY/v2p0zc
kk5PFeIjmZnkdBYLsR6n3C+BO7kVa1S5ed5ApCdlKsZVPKBCJwtVGGkS3Fzr/mzn
UlLZRf8tfEoeWrM5bigas6MRyoeEPwNh39hsFq7W7ZfQgMT4lZyo89LMoWd0EIM0
XO3N8jCps+mnI5Xydtaz54anyPRhQ9H0otwD5vEqNXoWIyX9SVs89SdL0tLlgR2l
oiHf1Ci93qqzfAnfFB6hwwZzTNBYKSwwMY7cL7SIZH0Tk+JOfdjFfivRO3AAFi43
SDoK7Et7peJw0IkVJvMaupdQsqGXoTFvmgtVOLYzu6HinMrQcLzUq1zGmYzCSF4Y
CVfqso+GlYIVJH67VoNo/U2yTP1tbaPTrG5JZmTPEeED9OBKrbuCqxUPZj6SUsiS
KGkfQBDCDKO+JJuhDyjL5A5yO2SLJ0vgnm9uOVQPG40XpqH2Tcxwu69bmr2UhDe4
dfb50fb66ywUnega5e24NhZvsyAPQvbj1vCmPp62AVoXbe15uQN/BCCyT7b1jiP3
DOu/jiY7bbcUpdEMBBot1rX2ZJ9eKEy9GnEVhgt8sgdkYODrYxn7p1zjKuF38nug
kqddi5AmuTw0NP/bggHFTiWKoXi6IgENZO+bx1tddRshW5bXlCeqj7a9x3yExBQx
4TnOGRX06GtOCTTIe9yveN30MDCO8jeBpyr28ZSYlFZ916ASR5e1rdhVDrkcFaaO
WWyNvzGzRnCUIA7kpxB+rTkj2CgcF2VZ6Hknxh3Mc6s6k8up8umFr7B+/AcNofQV
tJwUR+DqyVfSSV72jTTacKqwqEV7argPIGtz7dmp/JMiJWkQiL866eWrd3ExS6X1
4B7zonjvQbykJYOUWS0pS+BoVEHqh5mFv9SFiR5t5Neslo9xK4gkbzFpH7g/ts1z
7opECH5hiYzd8eGmJhSAmf5JFOtFg3M3HLGNPECo5azIfBhGjebL+j7DZ3/9spyt
LEe40EvcLvutslRhPt9ZBtfq6u5hvXGoGp8Ml+V1B83QfXp0GI42e17DNLvogHaA
fXCDR6cp8abZItB+21dP4TU2yEpv3SbX+3qLOLOe6JweaMMT3QzYrU88XmY3Dc2o
50EIo0GVu/l0fI6cFc2QEoL9OlnnDzaV1n8oF+Iwee+u/HSmfvGknKwKiGBqsGgz
xGPz1med79s5gMRyDeO+aYz2u4e7t3MxVoJ3f0zVY1Q0GXROB2YcaxjS99PaSeZv
kuVj2yWk/kNsnD3cSsMkft+beEZPRoLR+yY7F4Z7cds5XoOKvozZfHYpIYjeJcuw
pm+JjKEHCgsnZf24n0StDf6oO3e/uAAwGuhMXiw0ZO3drInQJ8fz6Pc+tvYce+S+
CYqX2iAbWeTgENNWe6qdESqLQDXDaxhfYbpzXgfsz9jCIxkgXEuMQIacTEjizVvq
m8KBhuO5cZPEqH7Ae2p27iBd0l2X16So0srz1pBHnszP320YmhRaJ66+Fm+OgzDD
G5Ahqe2Z0VJ20TEAXioKPqDJIPqMzIuyAyhw3JOBjyh44axI+FHKkn/U2/p6i5Eu
SCh9L1P1b3Yn0au5zqDUNyzwHOtdnY9cSyvjpNq3dM7n1Wx9/VI/429iXhlrzMpE
MO584KuCHjNHcLqczH98bAm6gUXsGfq0tXoSqx0+2TKEmnAxA1NXnZSLDP6xUYJa
71XcXxQQ8eN7sI3ceXsJDgHmyKdk9LM6a/fvtTxJqDrJnR/8Be5LrxaGJhBxKtUp
nHyvD69XKtGEYA+oxPaESdJfSBh5KLkfMvMAoWWTfbQPB3o1rIDF60bNwhEuSmKQ
3nZrjy3RWlp9pOXisROt24YznlISUX+WXJa9Ry9I6ueZ+M5a/XE+uJwvYhUWhtM0
9SfDvt9aXwJHsbUwfJbhHpynzaACzRYW/avTZc05hpop5OZtgktUNoxlAROHhOsw
AES76qr2QEcafAD+2wgixPttHBbraBs0Z1vJ0s6gv3mObZUZp00OZ9THt1Xn5QIn
u5R5Y0xUtitsbhSE32BkDrg2eBUi/tnD0Ob7crTcRKa9t/cTipyP2ruDQXVljHo3
1BfBneipyEpYMZfW9l8KqYn+YEPz2zggNtxfXTIDoo8OiqcmD5D7udWM5QS00GHo
ZWHG9oEwszT11+vY6ZrUDzYwPmkuHnmmBHTQAraA04kkpWZ1JYgZPhF8UySCHHu4
b5o0UYHNJzYoMzVUxHzrTW0Q9BCrT7THCm5WLHFfwWBWs6VJcDfQkrVdnq8Y8yVA
FFwSev5zyJiVrnxhnNN8441g3BruQFL5azE6feNbjf6oSkcAOBb6Q9Y1Jn67gNIL
QxXhJvCKrON8ctL82bYaUtZOKupLCeghHyUjTRCt7HNME4D5CS9RXd1j9mlI9kh4
3tMF7KF6bnBi/VCmKK2ozqqSSDedt4x4cHePjAmSLeagWG7/9nxCYt/l3LXFtFOC
u9UlP/9M5MeQBZj4B+TiCyK7bBD4G4eFuZab6DzzbbqxIWMZ2vJ03XAakBU8aJhl
3Z5ir9iPcm8zHrPAok2DNINAJAGzIwosj0EPAJ2l1pyK3yvOtlH+EHfKbSepbPME
dhTYe5DCKEzcsS/b01srAQU/CIPbTFbQXfZiq20qkVVUwvvVAoJUJjt5R2vY6wPF
zZjXpRIlwG1UZVrqw7yOW5ZW4xfsltshCwkfaqe0Fc7U2QN07LlNTAdh0neY0/JV
fEyr0t9IV6WzUkqBs3godO3fERt5xDbelo7l9LlmAnMA6OJ50JIBH/ZcuKivMq8Z
YQJdNIMXGFEy/PvnPC52B8cwndeNnu8sqSxrtwb+1wLviImKxTms9/qWIG9R6clC
C7uO7fdLZY8erboKdKx+htUEZ/uEOU5Al9caYXWGSQApyxNQCbDILYDtuUUamI9P
BxrsJq1ZiqTRHddZSrThwpl6vMiveuR0WQ3oO11URH/MhFt7siYkJowP3AB8/Ds+
EuLiyraNrtA5Yc7ve0e1OFnKnVk4pOHyIhlf7aqd4HOt36iC4I1smuwCFND6hVBK
yJTW0MurMrT5EMyjxJjRczFrFu7ku7RZMlSG8+y6CLM3mftPet+3BYaSHtJDOd3j
VNTUIBMu9Hh8cIXQvmUpPHoR+UZlW9Ek86yaunb8NBK573tgXcvUN4sYtvooEA7z
01HEaJCi2ooMMOiWegDMEsdsN6vVAiz7o9qBK/XXEuIWdoX1ig+bkwI1n22Sdurz
lHZZPm0WBC7QFX86P5M5IbuNJJoFFYVP1qu+H3dVbgqI0T7kYD7dlQ/4in7S/7AU
/fDStuNBtAsfIfIci91e8bvTr4VE61kl/ybAsvkOjM538+QyaRax95DZWfSL3sE1
Eb8Xb9Ym4Wyjc2knLmtTaJQYmnbFhSv6UKyaUe4HMcb+zVOIQJrKUbQynFVN80GO
4LiiHtxBaz2EVm2MZLfgIBwxyv0iOdfHcNtt7BXm6jYCyJIXwM3lmZ1xhXheWYTA
JrXDou8PiqikiGE/jjwairboOwElcz6eRY3NnhIHF7zq4YeF11FYdaKuja3WrvcF
h84yCMNDZXMItcaJ75qhDTrxJnnlIaV9aBHk/rkhDXCywB/qECSieiJ3i5ytgaft
vKgyLA6t4hdVdgp5m/U2YKTh2Axn3iFhlvC64ErYwlWpRmwUQUTpBrU4A1RLizfe
NmAEaeBwMTKjK51/Eq7Ny0ig7D0l01b9TmQjgewhNp3Qroh3WsnDI1CtbVIM8tKW
B6xRcT1Sb+Ncp/xHjL2Ke8+SBe77zCXXj5qTdffWBNTZOIWTnujmsDzkFw5RJKnH
Yh6cunwaAeYc/bdHWXvxwtMvF5QWxnXasHbhNLa0xGESMCg6gZa99QY7VPA5c7Ib
Hcu26Cycj0OLzitTdkMWn9oFGlwh98cY1lx5dyCOKhgnc6XdB4QDjeD9SHUhCfw2
NkzzCS9AkMueSdi+PFflW4x41TN/3ETsQyh0My+j6aax98vMRJ4+QmKCgV18aEak
iqev4+/tI5arFgixgHYHRsk9tJXYmFJGNglSV94tIDQJ20cg0NijX8cN4uTgjELT
Y7Oymk4AAd+Z5m4y99tqUNFFJlw11L9ZWjpd0+eWECG11KxJ2gSdv5F7sw1m+kOG
U1e2rvyggYVVFBKqWlBE9iiNieLbjPOS5Kat7KDIUhDo3O+SkfV1uojoy2u6gwWC
mjcXOScp9+QY/HFNeluDynrg3IaBBu4wi8uoPm8p3Hl3CP+H+o5HpRHbusWW9ENn
GkFkqGgljVOhNUuTEl9blf9SOO25/ZnbWxAkWLHkhaP4atpAAp5yJAXrqUpCP67W
syZbDLARMQu6jISpyybBSd7m5xsR7RJlYvePugZ7Z+gvz3jSolLRxNov+ANE+mE1
O/zx1vHBcpbq5bYni3azBvfhxuP4aD1LMCPf0z/NlaOtK34Cfrg6jpvfFvEAy0xi
5yxdK9thz6TOJLC2rzahcB6gYGmGB7+r4wjI+j9BRFU3tbbIJuQad3mC0vhaemDq
A5pM/0Dr3mlldpZIdaZf5C3vaf8nkJdpe/j76Vpl3pXWKlGABy0CuqG55so/ucaF
QzCY4LP32gi7nVCYR0n+Y1SDqNWOaIHZ2emaBu/jufByFXSB+S3/yx7fS8znLOFg
wJNbR3Q7PvahBo/tmyzyaJ1shB2cZ2jyxF8rQlCTAz87uJQWY3B3U75qsH1wfHtG
/JnaX0fjS7bm/GnDQJ77sJNDjHNoto150UzHnQ2NYgMcWHzf1C76piTr9W/sKOap
XSVDT57Hf4ecvNi8+iWFIhpjWH+kxMou2/Eqre/E9G/RrHPHYAq6uA/JqYReFXE2
YB9jlq1x6kjH+OKQqkrc8yDgNWwoC1uLTat4FTZ4f1hJ70Yjsvm+Fu/xKmSU3bf5
XfGtfMmEWamCQ9zuPFESBb1wOrALhi1+mqIkp3P36YRldx0GhFfkai+E64dzkYD6
yYGq40OBHUULolgwUPndpJepIMm0RWAKGaRo7LWZFWXyRXjsQ7vX1utko4YnZi0c
iq7/svdc4kWLwob68EWQFqHQOFZsPie7CfVejwt3jJHOkSh6c/Hd2QVku1j8aZ5L
0EDlI0KIqPFwdONvt9FwBAghvoUZT7PnZ8PIPkGqfnRmlVyvuidNK31q1Jfceeb6
c5YQSHnlRxYE20VfTj+NlLT4cTd+DIPCzmD9IR1FB3eM+is3r02ijHCSFmF+FSdX
lRlL4KK4W8he2sm8eOEfkO6A2SQf3PsdML8mjN9+hiY+K+ZqRhEyWrxK2rDF2rS+
QfZct7lD0eecoX1D6Bdwn5Cf1jz5d2I8NzM9+DyNCw+Q/BUIeTtV96DVF6GVK/J7
iaSc2mntuKB2PDcxRU1dpR38Fp58ll5Ka2eQneZ3qj5NWjM8vrpsCuWQ/c04hUHO
YW1v7qQzF19cY7QwPfhfy0ek5DFfTe47J8VAyrtteHjvbkYf1ABqcqsh0VB5Ocv6
Dr+19m22tZGWhHYQv/41EVjq23dTkax/9hQyJ8AAcrlQsxRd/dQYfoH/5HQSiH36
6nVvgrA4D8GP2MNqxwIuQah/ef5+jNrqWCyk/IZsSxFihK/Z8Ouk17WKm8MogFUg
Og6VRuLyJJ4Wtkm6SkBj4x0Jsqjh5WkXNPeuk/hjWM/rHIQgyP+9ZedRv2dC+sIK
fF3the6SlwGG0Ob/3qKHDFz8UyOBQ8BclddKWMIFHlQ1VJefvpDXbPRHI6AWxhQw
4ZXv6CgLRSyeMmJSGdATGnZFjHTGsmY+NJVoguNpTJH0na3NLibWg3VhOra0fgCP
TuP7muu4i/L9OYUsxG3O3FW+qiJqlLHtOe/gxfidp4lu2T6T1e5NKXqQ9UIMKnGf
plLVfn+54By/7tR36QZNvEc2O/oIFPp+akmZc0+GR4XlbamTQVx6VV4xOrGbQy39
wHAiJXcgq2KDXwb0Orqv3i8L/1Qt3emPVUk2AaKYuixQuSEoCHMkmU+/SzfIY8uy
Zyx8aNptK7TpMhehkQSP5EEcSRNQk24+l7MLELsnrN2pJ7qANtS0yC/R8lyqcaxU
ee0iCOxhj1ZzvxwSkjxs2Z4LAkm4YoreMVTDvvdZIUThAmLFq9U4pUyfHFqFpOdn
TaAE/8EhQW2M3fxiAnA8TjPcfTINShBEiWP+pmWqRbrwXS/ImxGgLChdZvBO5X6F
vkFaIJKEMzAP2fOGIHT8HgfGUmcLMGlPJ1Yz90MaBxmUN8uMcbYHdTSS4T6NKZDW
OjVDU/cvCpuHsDdMSd425dWqlulSLMmL4J98YoFGDTssTrjdTj6CMuT9P9Z340CB
VnF0Yh1UELgYnhyOjfe6m5BPtq9xJ+9nLLPBvBO+bNt8uhrSVsDO9Y8fjSKm1ZI/
2SxlduaApjfmPCSYXHU5vmXJJjv177fcie4byhPIdaA/+nL1b2Hx6zatFH9CyDSy
E5+otd4K+GoS4DHHA4zF3YRgJTT6RZSpHdz/eyYMSBLOkU8JlTW/X4Nv/4y6wSF4
M4VGZ4Dts8qImuDEpDW7ReFtihz3qkPMDgCagYBMkKHf26mJBY8Ai9GzK06s9FYe
AcTRDF4PtZf7hvSXZj/+mOuDzvWmKGp8Tyv+nKGl55OD8AHlUDu9rcc2MSWMJk20
fRugKVhgGW3MmP3uy+TnbtwIBZIM+kO/KkgcqlfKteH4wGS1OEHQm/DnqXmPel8g
P1hYTOo9Xylw1FwvdiYKImr//0RKJFzZ/bJAbUezeOh5l6i2tLEHPQVIW69HWVSU
1S3Hf3yyOmjjjFw+qjws2eKtyyDl3hrdK9kqjibdhxY3V2+YPTwqRku4KYxIaImZ
GcC0WbcNQFnwb02uzEPifqTB+bkLIL2QjYpBCaKbJZZCRNBas/2+v3DoQa7hZCKM
WoUJlIDRssrsuyFr77rdOeavlieopUHCZ7IRaHI0vPK3EOTMIJ1Um62imiqwSPj8
tFjoEx28Mjm7TFeVXdz+3UTMPT5j7eKgShDDdjRzvIb4Bh5+A6lNO78pGCVZ5jCb
5V0OPix4pyuXArQ4EMJk9sgW5+jdEcxiSCKJPhG1c1e3s0U2GjsYUPvqXfESpofy
184ymdJjqYmvFejvfxueFJWQb5aZC7cr6LzljuxLQMKRkqw+Knv1NvemWrhBC8cs
KO9Lo/Rsj27pwwCi63s5BLll+hh+nP/gceb3hxTM74EOo5xQTe6Qiir4LIwMO0hZ
WOYh7eiADegmojk8Qx55+IovMcJAHqpAey0EJ2hAmsW1shE9FiIH+UcPcpW57dCi
6vpEEEQoPRlaTIEbLl2DkBfIC4LcObR1xoBflOMFr1gdTgCZpe3srGET4jWKGxiq
/t9n9fvMbtVhhbCEB35ei4CnR8czgtdZcpgoTC2anGc54Om+cEorOtM5RUoyNtKj
ilhDLnW7N5Dm1M2TngKtNKXFTGkaUiemTelM1c1nM0B2X72FvmJyTk0gXVtXzqo9
qOTp16PNj8EDBGa1ysl/RUHt+4muooOBIjpi1ztHtCT9SUcU/RY3BNy1pmCniF/T
90jWjjWJG/6Vg5pX0z04KosKjrNZnOmJZsd631pUMe+CA0+V8Gaii6E2hN6s1afN
FepQxouakf9p3BucYBcCzt/gaOfRDoh/EHqivD4vsynnvhZE7RIVgxvc7D1GykJz
YzbZg77tyX/rvtunVnYfAi5PkQGQqszFtqcQoICb2Gg2jgQ7RcN2ItryGhCtaHtD
qXyFxFhwiNv3TWPJxCf0yEBMKBI/Z26T1tNL5CMgKA97CmEquEDI0rIWYum1DzYe
fBZprQq8+8HzGFvvlX6wXojoMXBhDSmPnmB0Ekg/W87MxjA5cPRWSlElMhU0eIii
U1sx2SPL9Xkd7ASUxbPu5bS28rQHLfUmPBXDtHU29s99WZ0mh7yLkrq/YJGCW1BN
i/uJVXut/+LWVc1KM39/jz43KNJx1hkXU6eA8AVrKBAhrUJcj0HoiAsV6RA5E2iR
emWoRRzLR082s0yMesfP3rXZuMfLkn91AOyFWsn5RDhkjRAF4dNjmZROB4CGb+ar
oC+H/qRRzZLzEpVowE3b6VswARME68TPB1jEA9XXuQ1yzFs2rOhR+lfBU2fWljkv
fYswf32UYxZ/5OevtBR3K5oiofpsK4Y2ug1SeIBmy+s=
`pragma protect end_protected
