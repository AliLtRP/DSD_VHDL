// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
twnk8KUstTWpAuMbzrzFijGp+JRbC4YHzRRvAfYLs4rfAROHiiyZdupAqcd45ei6nxZfYzOcD5pY
nXOldBElogzHCx2PbkcGjTBa7AeRXrKyDxkDsvX6wvAEwEQWHOce0IO4pU8UYpEemYX+k/STwB/4
fraJ9UHjoefQtx08/qpmkeJmlFUlRntBbkkKwUG5CFJ7640HWRvN3qXcVsKtJagU66lEB8OlQLIs
nIzIY5+ZKXaNRO6VF7WnOhzv65XN3cBj8td6PUcT62wdQZqBLVVHigyj0hz79IH+3LG0RviXpebS
Dkgp/REWpKGro41NcHRr6Dfvf8woRhYwVVP4wA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
km/y4wfATR4rKFgCxxxSHUV+ovPFHdg4kt/ReF47QeNR1yT4TAJ3sNlet07FNVwd5NG362hckO/B
7GvLlJPZOdJY/kgyl8f9mz+bhqnbaLPqOzca5BU2wgCyFPsTc2vQ3neqe3DNxS/eLhGXWIpcy5JP
NEBedIFbrG5qFsUO3F8PM6Uje8rJFFDNcd0gk9nwMPQVKGS7y/rNU1m8Z0TkiAOvdkxXOHds+Bh/
lB36fPzL5IzHUG15/6pVQ7/3EgXkOCsaOyztaZM5GPhVrrzgdNM7ag8YddNIRJSVDsGFJbNrEPHc
+xj3dJAOggvLzn8VNybe2Y2KVZWBRTD14MU+4qCopFa+ATgGCbV+1BPDrowob4sXKaGLcwXIOB+8
Xf2maDqaNPkqBR60MvYijD+IekK//4PTaFmJSBG6wr2ghnkOUgd0wFPVw8Ly1LyPeYtYXpGASf+O
35QmG6JCVmoInKre6K94U2hCjLc39BzI48wvybm9zo7txjNxqNLAYH37p4nEWcwUohxiupRYAheD
XB0TPSvhHe93ZOqffpnhnh71k82Y+JyxifYutQzOkcr4I1RmWXELwcpY1Lvw8eeNXkIgVqTx7f+s
N5SSo63SDm1qOqkmiaLFtFCf80ny4gSzT79NteM4vBIMtrIyt5e7Eou8o35xTp53e8k6Of4hFVKy
GV3lsW8amf/wVdu369iUFS5kjTslvNe9RsdxfpmThk3ElcbBkV/wHVlCWsk/821YF2FzQkNmgNVw
QylTQ4+IxYLfwiaxRRMAm7r5YoDaCSg4qUIwEPNxY+18oEAE6/MBct83HxJRLZ87FKXZn9SW3/I7
lYc1pmRg8hE3sKhDsVmDHhuxnJlqssDukb02SbIKSB+2htdsQkGpCidD54rszB2Zc4qdL5uq7Xbr
Jd4I8MwYdxU9Za1nSAAVE3aGEoRMsqRoZtVQKIGiH+0xOAVx96CFmwJjoJprsj+NPoFowHVjlKQ2
YYSP8pkvETcFwqYzU3hRg1xHJhDW05OY08IVqjLa76wab/lpwbcFs2R4SW76sKu/dTwBGfQ28nsN
w7n1LjpruByOJfXiYI5HLV9IiEwUUDwmyhmjpTSfYMRPGxMyYUaOZD8hAg3/ITS0VmnoscmP6dqk
iCQae+eggDaUiSXnt1ns3IerIU6iDJXjjwbbda5sx2hP+yckKFnnDzwAsIcZ0sycExtjqhypHB92
vk+xgVytpPBkBrCjUm3wNGnX9p8akiZSYgpwnp6O0xVFgXpV3rSu+Zai6GoY/nyEOAJoCLVkXiOv
nGJmOGLa5xrfq00l9gFlcqjQ+E3h30Tq8J9g2w0j8ndgbe2s6V6BaBbhb/oAO4IZ4leHDm2zhSNw
e6TE4ulkvPVaYkOPAz1o45N9QKYNnPmSgTK4xbzPacCxfEYg63oa/0JFLUX2FfFfh5/ZMSIjEsMj
KSLAQ2e/yqKN0+jI1tm2HGcEjkBUsbcpXvDUUaURoGoq8KWvhNsGaZI5POloGvW2eFkGdCxRBGDt
A31FXq2iwzRfUsBCidyrZgDbCVV5vd1T8HTVITpIxx3iRxrRyKLSe8YcZGoqWVfA8N6hsd+3KwQJ
HmChho4vrZmu8Rl2L9BuzHMCvrfeKTCrP8nksb2DG/6Hdqae756aZPluJH7IuauJ7INRkYHGlv6r
uNK7qj3njQrzRp2tjNx0EasTOxVLyOZDqdSIy7XYDzYVueWz0n4K2/Vkm8ylJM7ECyKq+fa6QOMI
W6ND3j9kjhFnBdVetj0UQpdvbNe+vxLkBeei5uCIqTzYtJa8OkZwSDQNVqI7vv11dHTwnmIzuehh
kD8VTDJPl7hyszSDucDBp6hezbU7cRE/yc4xmyJJxS/nV2HgKXfDk17LFrprpxgJj5NbV08byzvI
1xpc6wf1YzROyyqMIu+y6lF372bDum2cyVj+MfWDSqQKFvbo5kS8UHka1BetBZAeekHNha+8qlcE
8dD3e687/jLw2IYIp3FV0tc7tSc36iQN5IXqGg8ndtmVNLUR/doastwcC9r3pT6DIPs2yDkIjWeG
ESNweTHkOFqbimd9sida9tzCR52ZbPQtyIWEJBUkUOMHddVqhqUnPGDQCYOhALBx0XuZEq9322WE
OxL4l9djkAT6/jCn9wSNL2Sw06RErcsHcvOU9VRBXdAEGTlgRQ+ziL7Oos/IA2l04o+s/cPatOc5
0vWWY68o0lgRdegVFgfjaj68C7LpJWQuaw9+mAml4q3CD9KRlh+MkJmsdMxfYNNk1+wjnP+BxnPG
sD750eLjqifBD3dUTmECgLZQJCzdtDovD330dwJ0k12uNlMoEX/oYTjeUESWUvDtJ9+yMHpZv3Ks
3c2NLs6IiIZa0YSdLLL2aCXv7JMHboeyAGsW4PZVyt3yKIRDFf2ZLE4DIhsOOemLuZIKm74nBR5Q
AIDA7xuYEt1aVGyi6cuMugd58aM6uCh9wQc5n3WZUcqg83QIUWZKj6Tx2L2AqOWHQZ8Q/BJjVIU3
TYksw2GIKxFK4KzlI7Hb9OzzyhY6Dh00PZlRrlihlg1aRgpZs0AWrRIKEVOr5uIhCMu88kWjl7dd
VktOgYIK95x1cNpnCi5+0RS+9P+pPuWqSnOfQeu3nHbnfswXKHSAaKYHy7j2oRsrH7ppEUy1sSNi
Dg6MOEG3qPzqr/YJ1+IDWwaaBNjdhSC8vzCJj7t+v4Z+JXaTL4s2aUc2YUg3g3ZrWrDAqIonOEyM
qTJqW471MTtr/D0t7AFkc0JFNM79yA5qYTecQ0sbj4UFqzXj0uOJXS0vhEcRHzaALPj3NZZZ8ELu
WYtuQeCTNGF3tU38A6cm87xFw23269gBNtR8LaSXc9+eoXDVeSErCJxzN1fr7VopEuY4aR0cd1pn
kmspOMxg/hy9eJoXvo3XR4Q/JFUgophlzmEJVC0hKumjkMW1ZWBuDB+LhtA6zkwio8mnO+5HSIKy
uNvnzqT0Ib07RJfFOBIOwQG8EevpSWI3p/xzThw71GF0uexdMEi+NKO52DUJ98M3vYmZQiLgwOCh
kYc1WL7qYcZ3bSaR1SRtoiP/6NwyRPEKQg+Mtdp7IBPgGvcbOpVppDxcSUc82+SNKaDDNRAPz9Ox
X5mkbx2grOQCUErUSSHliUFZ41I5IL8WpBrT3tGedDB+uERq12Qc3qEzD/EH+HaGuDFBQf4fH2TA
Fd/ffWFVQl97eOpU7gppo57IJP3f5jO4H1CI6EE5cRE41aVLcB2OKvRWodHmvQIl/mciHd9MI0ey
okSZUkRi3Frw2YS8eoSLt4OV4iIPKeL796/Q9xXaB44g0Qk5fBmaxdGNO/WVVz1ESETwcmGxutNT
AwYoQrWg9NegYXQBscLwjSPVgRES64duNqwq6rNzfhMgk9tUvTRBcSO1PpMhYZ/+PIbl+ST8s48r
HiOzXsSyBxG63BuLIpqYvjFHLOtSTJglwA24SSpn/hWtRBIW4QfypgjXPNFShcsmfkSXgdYcN5e3
160MrA7kqlDRjNzdxGLwIeIx21pAYZX6hsZHlj7qiOAwnCKnSYPo05XfgWDYYH4BQEsFZjOxlV6L
zpvsOOK9CMg/lloUjNAhGU9QTmGdKENO6SfZRIbAYx/gU22W7wrEUR7VF63eUnRH6RNJSbYbU5l4
5v2V+Qlm6H5eAf8IsJ8+hAh1bpg7nHh4V3bShn7c09jQhSU3CG4fQSt2date84TODCJFneDO5y56
eha6U7AQF0vHJaGtOXSzmw9Z7HuTEOrr59CbWKb1NeVLjN6yTv+kMIqdZij37Ga6En5ylKWP8UAs
OV8l3ay+oXN+YxQP8+ECPkVruefU0DzPAiggxoZfGMaaujqxNtCAyorAgeR0NhTpGC1DFhM8sGss
IWB9+Sk6ACwFD9a2ZlQR3iYWGHhPu3sK85DfNk83h86AqsmX2nmHesV7RoNtfKe1vj4HGzuLIN6S
MZwknrcFL9KAQ67GM25+U83U723mMuspcqPjjMebGq22m7EkS4ItGRRGm0yUGAii387TTVnQnKDU
vV/HokuVuCe8pHLChIiQq4KWzrt2SDdqEzvKk4A7K1mRZoED42g+d0kvrKiHbTgTS9gBe7CE0EPp
N2Ips+4lU3tHPAd6NcKaTlhw6kAiKhFS9A8A5GW81LV51ech53mOorKMW9kjAI3Jtt/6Vudqj/n0
vSzw45pAHZ2ddHJOjtKKBCAttO2f57H2rWDIdZL5rkVHhWYQbETNuNPp6ghs/qVpggKTj7ER9Rim
rTy8CVu3gNJjCb8sVZ2iDoOMaGoeSXr8D/awIqysP0SNWPa18Hc0bavg7X/COzcr6saotAZhbj5t
oGy1SYKkl9kB93UQUmnANuWTXqf//KicglXmDXF6LXBeGTU5aqhA6WFzd+MceAj848WfC+8S8+Hk
+s0ru5FkiJ/8x1NalK6HD+wX9Jw5b4AZNPRR6peZgcugBxCJrKMC8fuUhnDqnbNnWtcfq07dETqS
kPmRYHB/kYZkF/8yglzpacLtwiqpXKZ8KTcUmYBM8jhW4LzXk6lIEMOONdHv/n0alL8tTBGMN8Fn
SruLObaakDZAAcGmL5yctQ9GK9Rsb3l7gkYIweC3romzPSzWUpxo8gWrbXzyCYXjGugKw2+JwQEF
PMJQZ38F0hJJ4pU1JBjTfLimB2kzAUORzy8lMNsy+Hd4eyJp/v588zCtsitjzRx/t3EPwfg9V2CY
k5rs8GJczJOPTL8rslF1AYOd18Kn7IaBrFjWAEboz5DKWFAO0obXlQ8j0KLnUMMjvFtQX6mJYhFo
91WNB4bx1hZ8cHQ+ofr3X3L87/NDXhgqQR+x9g4MNnaXrUolne1j76j0TbAckmOvawK+JFe4yPKx
aoQq4n3qpIRiYiLAnI+8kEzYemGAvzd1XNdKAKYQkNbWM12KTF6WyhsU643Y4bxKG2i1ygx2mCDJ
szaFUbVjMZyzYXWBrwndar/eZftyns3lTzC+MXCGBNqE3UZHTn9p0UaCHDjqJogoGHuwVEK7ZhF3
XS5K6ydOjPCKE8Z7BOYAL2CN5Dx7K3nuAAZhe5zYe8cgECqIgXPMF613LFzi9XivinC3fEz6A0WD
QpBU6MD5FUIzgOiaMEhIuTKG/j8Vw+NaLFxaXREJpHhvXC0lK4+suVTrBzi0WaEyU1cF/sqsTNqo
pd79REzt3RFW2qsGHS8lczszSpZ7r/dugSNEU5M6lfvzWKtNy9jlq4jzTrgkMynq7qQFP9KY0cFh
N/PZdWSFOCzqPbwzbUsbgdnO0+j17jF0gICXdqeTHvImhjsCMwvQiHc/TcZNWGm4bEwqp6NizOmB
LJDjHNrG2dEPxz+dDnpZYlynLgmgrlHr3dmSGjz/qFA3KUVP7bI9MF4U4goeh7v9L7Cg6noOESqd
P7AdJdiHxKFfonfiE/usFo1sc15dHe0nObpLKvZzZwKAC45yGqJuxIl5181f1NsVfNj88p6eSrt9
JAWflK35h4OpJ2NqDVXjnQOI4LJYfhWwdxI6+z8HSky6aCcz2kM6JJdalexF8CEHMqZFoxHCQGWl
Ktd/j9Tv2Y8+KEe4uXoWft7oSk7aDsYLq4V6WF8IrWDjL/vNTGtN4J6aBAwcDMqAz80jcpU45K1S
nbGae2q2aWa+Sny/dtnVbIWR8zWRu2Up9bouq/ZhMYmMC9P+4Z7BmfB8tBfJravykr6KbuBfJNDV
jHBfuL5ti/PNdifV3cbNEN302B7EDi3TXvz6HamQCuXk/JjQfUZ2Qf6u5d/AxkFwkdE/MK4mJphc
wvDJjIns+BM+O48F4gCef2hhX6qi13YKvluCSxdF7dAvpp7/Lbr39gieh92ycn/aWm95tV2lYT4x
X7QSnCK8B2vAp7/oD/Xxr2ADBJa2/JNUwifvkpSehutKVsXNCcNobDbTxXx/D2QdIbsyFtSfDnFF
TFGzgBfMa1K12vMMM6v5RbG9NMBkKnj7Ry8sqcS2DfvaVnBGS4evM/dcz28WkzAOd8pekhIsEPV2
2t0xjyT64KqprE2rTfhjMUWhGIlBSm+RvJF3Xjoj2UVcbxB59zqbPhCK4b+ksfYTeHgs8o1ozt5j
PcFbZyM0fFoH+rz/TniuH/8uP4ZNr+gEs5jW7YoXpFKch6yEi6D30D9SkeIOJT7LZkeWFsvsGUxi
s/fUrzkitvUT00iAApIhf0fOeulplK+/95Md83yE0H3UHgMyt9jRAL59lz3ixeGy62mxkZBfgijb
XVzYMhtL3PtHRp2f/ejpw7ZwDjIIltfPsjldVRXcEmvyA+96MnMgnsMR1OhZJQcAAnjQzSV7ZjWu
C39BWqiZ/vF2Wq9c9o1Fe4VK46fQEqTq47GcHKbNoYy7jfoCARok5ISjSKD4Tny0gx0oNrBzoR6f
DhbFmjCwiDNpXfNgl92HlCcv+iwSSbc66H0jN3lKbI0Qfm8Ef0lGhxnuTdqc+URObRcXvFnC1svm
8ySplGcZ66VdQ443xUxagVot/j2DRzacvm2AXhgzosvcX9805N180eittVXjGg9TiyC2cbz7Hi/a
zzLaATRiODzpgZcL2OskA9P165JxJtA/6C8/2MNUAHeV62zr3aEPgoGDpeWdyBB8NVLSo+nIuCyx
TAloEH6zQxzmChMV7OWOjBYPtA0K/n1MR8xWppyfI1I2HV52O+o/Ra4CdFN03PtM5eQsp8nPDHIS
IJOLPx3aFJG7VVWAI6xLfhLnqYbGJNKxKPNnMm9TRk32/R7Ig8PDyF8Vr8gW8tTDBqN+judrHnHU
hHzqHFPUNImn5wZ+CZfdxnaS4p8l7gTi34vYBgHalmauVFXGDr1aHWZNBc8TOBWdG0M3eCve1DXI
7k0mlBWy8sslOvLVL5ALt8zSNDmliQc0Tizl8BHQFG+cvRFUFsrOTqx4s6FbQLoepvTxu+PuV+QO
Jce/qP0/oDXobR07LZcB2f+GVwfxYLfMCjry5zK9bSZLXmClUo08BLQwM6K3cstzMnSzer60rTtd
WnRJ5dCyjriKaxAEVwjqJSlFM/2t4iCw8e/DWE6HuALXcqp6hViU385EyR7oIMTG4OrT/xYY61sH
/roPcBFvQJhCgtfBJflIbF6cSBx2AjRhRDMjhmSzbFuV3JcNzgGJmIaURtvgDRpvaeLOkfpqBWeJ
cxRqDtc95uJsA4wd1bfcnsQXHdkS3izuQs0mePklS220PqLdPqLVN8g9zeqDMaJWUbTd1mJs4pG1
TQEgj8Q8DzAekksnjhoGeDBP5aUGJ6zNvCb6feDTkpFWpTSD2eIqb4VDbv5hQlI7iJpPVZph8HQS
IHIJxf8mvf231kiOCMtzCLLo2avB5xY95T6Y+ehyqbsMVagW21brw/lVCSW0pWjjKbPRaQHf7xLD
qwD97F2ZS0cla8U8QKUFtrFy+GE6xk4vd59EnPSJ0HfZfuga1x8u59Ly7O+2RsQsYBrJ6kRKeL2U
GBN2nJz65s27s76qPhE7WS6iGwXLSrRBR6lJGbaSsuDe//CmtOyieHyCouGoEbLJ1Xt2rKXeMVAk
lb1b1dpHOFHGRdIaFz290sJ4Cyw6EGRHVugjvZK/U4gHPsNGYbgS14WfGf8/cEWaRZySyZQWOeiA
Eg3MemYt2EaDqpXji6J/0CTe14zrBz1v5SDry1Knz5xMAh17gIO1NA6pmvdpk8x/ieLs83hVI3JK
u+1c9BRsMeaNL4zgJQA8BVELwvHGdy7TXaPiVqN23sJwGmDoFM/BCOl5qjzcOQ/YwSfKrvj3pS49
JaQdEEzhrRL6DqQ/j5KnlcVO83zJEoRqVzdqeaPss6gNGBqmQ3X5MQ2tUsxJx6/RieXHeuHK7dM2
R0pAJzwhku0yGUZ1ylmL8ZD5npZNqoBoSjwaz7ImQe1EZ1o5cRKYrdq9yGUccV9FnD02Qvv5gGB1
PkxeIxdOfx34n7UAWIIHdOsCwW+AXEgZeFrm9XECsTgyySH4SSey4D//WerhNR54i3Hn6trqGcr9
yyouL1LVZXbuiXQCK0qm6HtsJy5Sk/zczzNv8KnOuESr5kGkYDgEFafgBYWtUqsFvvPkA4UxrGxd
aaEO4JTvWsgJ32odlxfeta+MvMkQAoKVn/HTs+j4/NcPZs3klF2/iyTN9aYet7mgFGU4dH5sJoc9
qrlADBUU4knaF7xhVCGph7b/X4nV3HRS3G6iK7JiVdCWqHjjY0XbCqcRFECYhV6n6fiOoIVv85ZM
ytwxIPxSGKoqPbb5+/ba/4J3bTMwoNk6QoQWMGb7YpHxXMw7rKqjELcD234gnW6Gt+CcJmn80qhr
v5rU8DsPm/n6lzug1fE9TFQIzBDXywRglNKJc7YWPfELkXjMUe/U9mSpNLHz7at352Cg6WpDXEqv
mjZhC9ptayAVhZA5oLq9FknGUf+HtFZsoij8W5vXHotL+2f7nWK1Ys3YWsXoJ3Z7TJM5fmLzYjh7
o5uvMesT3R89IqgYOVxbMrV9VKUaBayW6SFm158pnqlg3POUUJSkyNGTEXjqAbA1Yo90lvQGNU4A
9gnVnjeXaaWwKEtM88bmPLWU79rxPzmlIabzUNuZuI9pnMJAH2J/YpAbeVdpCSHLkYEND39ia8Ow
VVgXN+3wLiKPj8bMz5sAQe7xFRWJaPQ+LDUJf0zvCgtyGepZeU4I+hSzbF9eXpCkJUFpx/91v7Tk
4SUw35xyDfl886WeLiiMG36Ay0pzYk5OD7whKDZrk2ywJYnJ2JvNVTwkhicJjv/+QwTlEIoDmdKa
WNB9J73Q1KOswED2v/H9A9N7jn4i1ixNifCZu+mLbrzdHyMDDjcWkWmjIDwH0B8IEGxgfzMloxoH
rc/e83Doj+TdR0aUzixijJJH/9mN60V5Nqm34A98KkYV/rnU9JcJF41OLWofgXeg6ogb++/7wjfp
fZ4/o4GMgrp1+WxcDdOyuxsNiWotixiqRBMlM2I8DWQNLqP9l1hkzcWF+jRCDNqK0gfklZNgDRKk
mmS3fL/ZfFPiuP/neEsOCq/HigYzhfyhuPjg3QSEXrmtWRPxEegGN5/zcFKgPaRPINhU8SdtnkgK
Z0M9ABWAHg62KclCUbQ0vTIqvCWl0DTK5ifvQHUZ81dppxtu5sD6EJvU3Q+7k32JdQPtYrvHso8X
tFLleLzu9CfsWvGWHk2rfsi17+b4PhVEIxa1fF6nEysZM9LNRCFYA7bXzIfH/MKaNB9pP3TbawDN
HPhoXAErzk6PMzqQLHA0FfHiDr++esiETUVfvVetejLYxZxnTOBxtxfFpdHHfdHU4nZlQ3wd5c1q
0xXwKtb68bMfoV0LnSRd9C3FB9rNTDMc8kxOcuxkQ54e28N7o/IJ12v76SW6+I3FRZxS+OQTzEYu
96AUgf1jtp2LWvpg+haJnjGj+R3gCj5G5kplR+uB9GfKCApI3MQzOQfmpCJQPgs7kK3YlWZ/FeB5
wFPFsaFAQQwRFAEoJRHfmBNOGDs2blMtanQP65wTupgctEIg+4GB9ob+D70BWzPN1jXdhCdvNinI
l3LfPsMxWk+MRCi6ZBAChcrCDfmblmq+dAv7VTh6jatpfgMqRLyRF6BmAg5+alOjgcUMj3O64z9R
FP1ojm53rPybxImHs0Nfzp9/bDzS+3INBGUaJxCEZn9tMFfZUJry2dJq6VaWQs6OBDmmntKQeI5Z
zpoRKmlzFmcer/bwy8lIebloUkHvzzmwTlQFCprnDW3AMg8yW4cs6ktnkS3EkMl5Gco7fccdYdrf
pHuei2EZ6bi71YWuiTw5jtf4TyahDNvj5uXTaimJGGImyCTLsvCDet8R0QHyBuF/eQDQDVbOyMcW
sAKDjW1de1RrU8JLnSng8IvAqkSHPkT9wPv5hptVHBQqfMnghwqJF6XqFdHZe5sbhRYxx53WhJ0j
pj/bQdzh6HFaJ2Fc0ysZMz7faaDe5x4Lwr31RAlfZA46UngzpHFR8wamRvG93lHILQiZiANR0l+W
VElqepgOjPbktxa7qxYMUy/OTudzt4GMNITE1MZp43WVKVm3+flalkQqI6V/mPm1rgx4IvtmYwhW
ud4Gr9B/TtgFHsBpsmCrL/tck8oXISP5SPnF14rzXpm7PM3hNDAvccA3vJP8PEgpk1Ofna43ni7r
EmjnRJGQ03n99zQpl8JStXGcfAUp9YGKRa9Mr7bZeBZ2kqsslDn2l3zSLY3Cgr82P+VPs2s7M2eB
zXJDCHbrAAbmzUurdYj1XEBP+S8strhfpXePSIx4pIT3LMXG0a4a32HmK7o57TYFHUZQ8pcKEarB
BZinQB4p+5BWJIU2R0SzJUKI9JJPEpCFdv2nd/Pg2xX4QhjNy8BF/R/vvBS82MSDR0TtWjQrgMeM
fINiFcj0iTrjI5PJbkOAHqa8l6dQcHT+Xroyt9rTSbadZnqDj+nMkedWudl99nXCaVAjmeakisal
V2T/KpiEZYTudKmqgDX1KC6djjNv7x3Xv4Dy0zwtedWT77hAks1luXmDd3hIH/zjIwtyzG/xVNue
w5cOyEacC66rzlVg7d61vLwjhsQXRVyopfPfIP7KhwNV8CJEM8yPGksLCD3Lco9qhqgqKcOUhjkk
Bxsd0EvmZXSM2sFODIL068d4I8CGU4NcWCo53HaqONJxyiaQJyqkSuQ7vNQX8oSE4VUHP9RUe0nr
VLVYi5FbVJGQp8/7KotfaNt7NJSO2OCCFGnTzXmwYzILrweSmoSeIxQhRNt7cG4TKKvpITPSTIh3
G7uMYyE+GDTDz7jtXwCPO6C2Lq8fPKZYmcBvnw2aRFUgHfPusQ7f0TPOQLF17bW9MWNk9JMdG5nJ
D1YKSSk2TUtvY+eq1PFLEih4d/RR36FufTnTIY8P2jnnr+SbHVgT9hQ+KotGu8xtoioMM/OIDAqq
6AoiqlOMui5EceiGo6ljX1yStU4lVNg1M3Ic9wgAHxO8/DXF3qJS9oPYiXFqv7HmatMQqAvW6y0S
TF+JU6Kzf6Ied840OXauGyXtq/JGtU01k5BK0R2bCvkiqMOiOEJkTxkVwfwcN3zqhYUlM89mDjg9
exwy91iao+DBwuTiYgiOnHqmtFYEa35T2GaxHjkPl5qet1/m/wVcnRYp3Vz2NnrAsMOyTu4/4OI0
dYcLTOh8rd3IrTXmp4RJgh+P4Zg1cz8hLIAfDNTPQLnzLbC5qeytBatecgnPDn9TJHpl+l8QRLYl
jZRLB6jHL+SCMQXd50GF4wkjszVt5Y43uizPoXyOQ/WYuB0L10ROJ91TE2Pv4NAyCbrSGc5sqfGQ
yfk2p6AZxiVdKvYax2frnWJrgSSaq9TOraI4Zsqjn+3DXAZIYfb4sEgOHiOMZPpJV8+GUEHz7r9N
qSh9H2hqD2EH2TBvsi5jjhHP9rw/BVnILIdZlCU5UlFfQrGaHoi5bGc5aH90Pl6DnfOTE0G/+EL8
GkI/NBIfgdE9XD/cGqa3hvLXkZYpcuzD8STbH12RKBDfTbTcUS/PYL0/1XWi6TLnauPZdYaSha08
5idZ98K6u94LYQofpmZM2eVxBhZCvqg1/7GEIrmGNU+qczmNm1gF9/MQgwlYavhYFwGuwBsqr0Ty
6R7ROHPAFCg+IemVRlJboVvOzcE0TCjX73J1EYYERGI5zKkQa5TnaUkiqwK+0g9vi+B1XIbsCuY3
hpqdtY8qTionoYBccw1cJPl+mKZPZjdFlBNqYboZWCWU2LVQoppAKhNmH1Q53/rBVZ9Zvg6b4vcS
wP0h3yLVWs7LmJjkxGQF7/lQnmbXF6ER4VmfcKyNZvtltcPHbhExplMLUQOeRtY/aLrUi/agcnuS
Lf1mBgsiL77bXrjk8zBUxSuLT6ITjvqfLfWZI+n1mw9KIjboEAyGLS9AxzZUSHsauMO8rxHslFf4
04nvcWy2+MSo9U6dClEdo6vYVKwHIzz/7m27MQ5ZZWj3rv3e3H6Y+Jdbg78MUFGcg1ed32biqJeK
4Rzj2GsU4N/+U/KsLfTqDFAgFgCbh0R0F9j0XERzSBQpqV42NnyY3yjYWL4d0/cxpHOqWtZL6ANN
YAepWQV039fgIn35DYNzGOq+zyMFv7uzbHvs0YQe9ADEhCIIMIxfxZNQsXHMvCOTcdzNFL0WRzVD
aisI2NfXUvWNGUcRZtjRgk6CHvVlqOIXfME4z1Tj087TL44HXd2c1bfS/cBlzhdTMVMhKqUBDF31
caLBxq3QvoiJ5m6mjzL1C7Hb+eFTJm3GR1RJFK3cERJzJWOW9ztTMFD3nBdL+NtEBwAwqkciLSFF
CFUdQD0aLxq/FNianI0u3DLavL6+CDvPTeVxqdYV4u4yOHumLKFx1mb2w04L2PEZr2dYyzZAXlqk
sPMiCaqqB9V7llGRHzzlaXG0oKWT0Kj2/pKYTqNgVtNz/8F6ZgO0Zg/eQK4WeTf+s2f30DVL2Bab
0KbeXvcIKVhoBM3PTNOvRMkFeOR/ziaJnLyQdQirUmxzuqc3OjYksddc2oDy9ygaOuLAqfCRoFc+
FhlY/5i9alrtCHbQMuhvJyZchYV72bxOg0VLGWpxZnmOcsZ0bTAX3C1E5J5cvTMYf0VslJFyvXze
P5zN6cVMWxU/Kzptrf2a/78O7wqaRNo5b/LD0GjRLfDdHbH7NswT+e/o7Lwulh+RmGypPcK81/34
AW7o+tAXFemH8AhKZ0KQrS03+36PkQNAgWCUroTnG+isHybS3DslYTWcd5WQWrGtNdv1BemdNudm
yFfKu8LMLBt/8hY4opjG9hAT7WmBB1PITaTTDjUrVSkHB20RKxcYqwuyp1CyrWNN2f0k2y73KJex
mXe+5QlDSmLL9TAjvGpTVuW4/BSoL7M5BWcKJlACT5BiPOdP3PmB6FjnkDfDg0QpjOYKcfSMLoM8
CFbMekMilhFEDwMtrt8o60PHpbs7pUajpe6RiAnYcXeKKGST6g7WaYvV8nVNzHDn+AEVWToZaZFP
ON+Jrd145ypcgxjEL2JydJqD9mO3sg22mZrzDgCH67tcQGcjjhJ18t5dp0fr/0qYWRZG2Pzv2Gm/
vdRujs+9uaNjuVKzyU6YHHh2xdVOuFpXVispk1kec28jhmR8vWmoUhizUlCocNxf+V6TpE4vwhgW
Ib7a7lxRyD1djDXQXVe4HF7sU/OiMJeJcOhDUEGXAIpOMffWj0ORGcQRmja/cIX3ufZ+qEa0gMe7
NTK8XAUqHzjQuHqhfCSmm2leCVbv/UmttIYpTq8fq2j+2dBDuzOlqrOIS5q4yw+EvmtNNtjvgVdl
BfFz6e8AmQ+rozJiuFtf6ieZ7yDUbzIIOvlz4X/E3xEO07EVR6QQ7jmr+w90tTlNiHJF8i5dkbRq
LGvPVNhonbh9gJWY1zLGZ8s0WzVByb7d+Ns2oGMo35h8e5dH3QPZpu9ya/Q2qKYwEr3HURFzPuEb
EUJRk3hZC8FRD5gbMdxYbrQhtCDrJ3sYaDXpPzrV788XHR8UCYnY5N8eFWVmfVL2Wbu4Lou++MDc
wbm+0nWUuPvCzxUWDPUUR0G73MKX+BWspgjuO+2uezgMg+lHzPOLlhbouygk8jm7jZs8yT24mH01
APie/EZvxfwrc8jSNziy7PYnNd9B6zNft1xGZrAers4fwwJeVdnmTJ6VJ+BRgqOCNLSwee0FsjSC
wIwVCCnHnwqPPHp7MQWw/lIb9Q/t67tWmA0a1hYzRYAW6IUWnLs42tlmSObqNA8F27D74/pQT6X1
9qEECO40PIYhSXyfOUjX3oBoAk+FDFT1OPl+Vnvc+s556gxcQ4djrjCXnAz9rpjJWNJM4sXeqK9+
vhnOv4gNB0RHXh/2j4d1oLrdsJ+89iPICQz2Ldd2VSDZUQYUe/ezyWKC5amy1rB5qOVPhcB5Mxw4
QfnjntH1XWlPU9Wrovi8y4E9YZCc2CW/arBDVd1qtmpRA4DatGp7itcGBIcDRjVp0Tua/TVdLvOP
d7mBfOnoRz0m5xNHm7Yj6mDqt9mI+flWuUVXaXN3iA4ckSNJIL3nEb13K+1eD9vDfJKP0S2m0NbT
urEHfw5HTz51WxNNmLemWy2JUB4Hu3H3tusXTGKUUXktBSTFZCr5EvuBeGOA2K9LnsDqIDQD1+Fp
41yQ77o/xwggGESqTIfdpJSz3/OTSgzbYtYJ2xxgMfl5ygvbUvFzyCxTI0z0Iu9VFcbqW+knPrs+
29ukRU3x7O0EfeOlaKcIt9sW8BQQgojMlPr9z+jMnxpxJ+E91urlqGJBArlzxyhAzY7TYcz0qqWp
W66JFmuKlPR6oMSWmB8kenKT0rvAht6NZH5oz/+uDmSHdBEn6hJnzzPnObKOXMQtyP6rdqc91hZE
YkRObls09JqeYbTiJkZwkYTfWECMzJ8Ymb5CXYcVh1qSOy2PR2dnvX+TiGECYkdtMcNSIFpMkedH
4Jczm4rni4QzqnDcZOwZ4V8YRMyKhRLJ/qRvAChrf/Jpcb34Z9yprRiudZ57qWhsIc7k5oAmRxdB
+s7Xn+9QTlILk0jvyDqJXyQFDetr8RoBwui0OOSEBlbVPUZwLurz4j1GegI3b5tafZkCOdZxNf4U
J/9BS7p2TTsmz9L0x3/rggZcOQQVMVgYntwl0evYJ03404rF39164z7K7CWfrh3qP8ZWC+41FJM6
o+Y7XSUIZJgHhhZZIzBRoHktqwGxnSUkQmcrYcPVeqmg957H1uFXl3HrZEfkRVDQF7PVdEHyAjua
DcidM0XUnrmaX2iWkkVtZUYejJeLSAy7YUskhwqdTjCLwOkDgzPyHXVJmuVv4TIOAXwYKblCuABT
49QPQYlQp243p6UtWqjaRLCVO23ZTMUYdZkBT0OxdSk67G3xg09cnkEE6WJQgbmwLG/iFfi852nK
BepwSK4FX6wOY9tbgGxjHtI6qnAX+FTwWeMLNrNsKAijgbe0S/9TCCv/nbb3jZ+y5GeJs1hUhdkU
4Purac9Wja9VL4fzPu4u+jOLlSAwlNxUEVQDyaMqfeY9R7jDTlS8706psIj0oTD4KCFHBTD/Uie3
TUFVxvZTvnubD7Cdnhn4uqN5V6H7qeles7LPj28TzpAllJwfe32RKT+ZgEDXuUb3Btdt87WCirAK
R9wpLoXWge4i8kbyzbdEVi49XTDmqxd/5GBy5wM4DMe7E+hezJnQRpv502vR0vVi9TzLqorDDn8Q
7HQtsFTnlyQq7EvZ5EdbEnYX1RaYxubmFHwVrUXJ698DTk2B8C++Rwxge6sDFbWnUDXIBBTA/vrd
cWReC6ELqYHBOtnbU2DBlcqICjIC+tvKvDMIdv53bkAYFWIaG1KlVH3F3Qw+AbtQM+beaIBHZLeg
cOyNQgSELTNDrN/vabwDiY0uAVY60RQeGR+wSd2ExFZXDekWqen1HxmE1oWhqaUdpm7DrwNQygtx
Sgnaq6CssTn26F0ahft7lTx0yphu4Ry11XSw15d6Th7kOfoROkyGGTYkHA1SOfjP4oGi+IpZk07H
EXjF7Z29MYgPgqReZsgz54jxU2l+QqmQwF+xOH/EEsC/qiEXUz3xTW9y20g8H8Nv0vtFvbcuzubK
LUWuUTiZXHwMsvdixt0P9Sc2c8PpET+ff5XiIgaAEkIROo7Dc244C2rE2T6SueC5xM/J/2scAFsl
BejeC2cPhX8WYvpABc/MFWsxBqBgdmztQm5edCa1ifuXtxlMFyTrehehsI3blCNWTrV2F+SJ1e6C
h7EpYtzxk2AgmqDc9OuiyIua4uDQ2XCdmYNE/Oq3we67zMuR2kAreLqBjjlXVnhA7/xjHM2Wi/hp
1uSAMLQ13TLOKti1YsK7ZPa98FNks2nIJl2NtUaQa3VE/Wt6t+Sr/4v68N97oIH4f3V5onakOfrl
LvR4I3udAHeUzO2i4nUke9CRlPP4nhrMESDYLNhQHKQsCw72d7l3Xc9Xfapd5DMdbl6Q4vvy3dCM
heX6WCveJBJ4krM6GZR1IPQcHwUtBxw3cEJi10Ei/Ky5y3/dhwv4HHKir02DnnMR5pydGu9ovvZ5
HP6DZMhnCIJBO+TYxLfgVZ+wzm2tPsQReXM87FM+7B2/z7DyurwfUvYhPQLz8Jz6rVodlJaPKfX+
WglRXckThD99cGRbEV1vLewItIlZo3/LgwpcnVEJOg2KHHImXcLbzPw5kJV6HljKC+qwImcXgxB1
suqDk7Hb8DHIrASdQHOVzM6dHBRWvdJidg3sszcu+3BiXWepUOc1U0NlVssICoB2h28ew6DTMSwH
Vxidbmr0zO4NG3ahYdPL8Kx9hV7kGqm0Y+CgUirYxSlO2ch0+QMZ6nDGsV9neLb9eUJW30M1t6CP
+b6zpolRuUYOkae0i9jdMDDdiQWd9sgKT8JqxtvNo0I/DmltskZdDmDR27ESG+JjAZpVSYIgE7A8
WIm2xiXZKSlMFHojPNVWL8Ea0XkWsHb2JJNgzXJ06iSQUUamNoYkKx8Pp/FkoqIlrj1yz8HrQ9EQ
zERPeqP+3WpAMA4srCLCpR/xUJNksrhsZKvdkEnDSmYNyFkSMRdYd/RuJHjwnfrUzsO2xtqrvEx2
ndiWd6de7954GwSLgRnJm13OJL2gS/aGvx7udgvWwht38Vbyvz78xnNk7Nfg0HLwGw0gcJLsUYEA
mzsDTpLjPjvnTb1DyE7KbhC85Z+EiqkCcIFZXEBeu2VX9fOgYmC0JqmuK5hL9Z3ZIRufrkOdUtcV
67P5x+J5OcQaXP3f8ASpc0qzUK95b4x7bpd7m+qu55R0tQsDCsVKPAsAJzNGaHceXbMoiEwcLUcf
6nUh3e0vxoPO0LPsh4fqFxRYkxpXDdayI+e7OODG+fsdMz9FRvTZRoZdKFpkv6G+KuAfkZUG7UvY
TYf/weE70iva6KHFFS/kZvP8qLLXt9kmzn39EPnUgCOZXVuCYzHCWN/7GfdaHUxAXJ0K8Jbzw/vI
SU/Sg1Kb5z0iX+67fTTr/h2ntiWQaDAF0sUoXaZUOwICQb751y7c3BPtWPaaGwIMUzzSpo/yxRlG
thdIHWHJa8BQ3tqoRBLWL2wGdl62G5N8OW+MhCuOi6DM87dT33RSdhoCEBXYLZ0wXKW36L3J2SEU
vrpNG0qPefKeKTNjt7JOqEA9soPqDwE3wmH9VNxBz2V2TLx6SEu75Czh2AmjMntnmAxrBLeaIRri
z+j7tM/NELXEnfC6gr4vuWfeevqrclCO58UCSDhAWRYNN3Fo70dErPs3dFNBxwYMnHOpoyCk99kX
OYoLpziT2Bc169u9w0GkaRDhrd2LxaWuNHkgHnu2SBGOfmCWNKs9exhIqw6nMfTXlaMygbxt9wYt
ZC10YtrdSCYcPYO4ORamSVqy3gJ+dGs1LlVmYtEGZAIq5y8eGNaYyM4WUlpoAHojZWtKL7XkcRSd
F46LwRmkzYFJ7ulwK6Q5sQa5m0NM0jo86I7fXAnleNVt+eS22hJKUO92IEZk4cTiC1sW2uLzvXWt
3xY1EWiGV62sGHnhjY9qYxj50PWE8GYcGBaYfx03WdoXR9bizIEzJFcStOU0OH2C2iO5Td3zqeAA
wo+WQBW1RtnW52E7YuDFfuDBw4hBGOPV7Pc1l7TH89BLZh+UQOTGYzSp+njr+kFwr9B9V2sxfPDu
BgDsvsCcruSfP/qcGL4NFgoZ+LC+jR+PjPGHZF/nwsIV5j9SM+et5AagoAA6M+IMlHawhLC9EK71
WrKHfyCCP4xIBt8+P4fgJAkKQpw1YGWGvBgChfGD8UhNSJLzP14kWW99qYhIcXEC0uBExHDebvmC
/IIYYjzKLXCp+Prkb3DypPIRq2KsU5havmxBBDLbryApy+mzt1AC6xLDS/TSZVzNnK+TScqV6gQy
OIEiFAsIIfMDSkg35JwBOfYDUUoyCbHkxT/E4diwRImfe6vYrJv05BQ2Pa3JIzZTos4n1P28bDzO
kVlA3WhV/MULD5apWu9gUi0vMge9PIUgw2LPhIB1+CCsn9rHYFgVsb0z+HXXkDCM1POX5R0dzHhJ
uzTnJ60u3EI9dWu06eI1zDEDJa188wTXp3CeTyQKMJEFPQKXM3BcxJ+/jKT8nM2rGE7gihBB809Y
2P43SAT8uZB2/1gfSVc/bIGEgLfFKaUVy9yRsweXY5SxGsWooydVHoBC38yamkNckpX/wxeoDeqt
QzIuAsttjyC2Xh7TPN0oksOELN2PbYV3ff9rTDsMj3vgbnXwdA1zbPSaNIxXU6zuPxtTsKPdnSmx
XvMFP6wtLAeS2NRbfJSUUYxZFsXeT5hPIFDvwtYYVTIWZFc7wmWUnEKL1u5mkT5llsSoZs+4V1/O
V94rD2db9OfpE8A7yNiITxRRGc56VclzwBBp7h2Plf5CaK9WK8Vuq8fd/C5OK7ZU0b7nMPrTq1TJ
uLOYXgqpc408nlnzeq0BdXpeMEirSl6bltKowc/mzAYHeK8phRaovQEiFSTKhCV8bVlLr2ZqioQz
nnUwH2ANCaydBIVUEfx+hh+QRESUxznHk43Q7j4q5K50DfV+aE7622+T9n+B5or91PzLSGCHU7r7
sLoa6VIBi4ocOmu6+Oo9OYb83QCPL0hZjZGeacWXtLFemIc+nPJ0840YNUYq/jUJHWbB82sNUFdm
HAIysfBbV7KJMpuR48qxh1lT7yV6fRvgOcf+HBfGBLXJPPjCKfs/ESR/jVgyYveOmhOEiUru2dMb
5REdFch5cWp0tPjv0du/Ot+KZRBWpCqKV1l3UORBKXC4kVJCl46nu8OhTdxCIPmr2ru/XPrEwSmy
mQFcOsY2Wt1/3qdUNw86Z8YoPyTrPoffdFZou/ZZNZCERgRTL+zTzD/YB/qQO9J1ZqoPDuigs1Es
DvfKcAHdVQZ/TKIYeeQj7i4lTIU9dU2LORR+OrDCKtTl9M8ohVoG1wnsyzo2+2raxdSUiGH6rPL2
Ah6u3mk+BSa8DmtUT7qPNuNv2lXYLNcDrdCV8nHKnuTs+YZYBwCeFlg1m86sfR19bfHtB2myAC9G
tPteFFnhM1kiMJJJimAaJbMvAOHUvT5oCtIDStWxCc0l4aJzaT4zWC3fgVsVT28lPcfkuJB8cT+3
AOiYXwL3cFdPbgxBTTuiqJ0R1r4rvLvPZRd0yLtLQF+ueERcs0/GtErRoIu1IULF4soFCWoEouhf
WXILKzKjZsa7gYeBZeWv3baDPfcZW+2lCFmwV4t8s0+sLeZA8d4WVJcaGxG+xvtAKRTgzjpK6jNb
t/u2ALLxLz8w60GOX8mdbfE+EUxr3G112gIq6v4lgy9mjlxMP3sJBz158Z5T4ugMCUY4n6hV0joo
5c+Vb2fR8ltTKuZ8N9sUZ6dshxbXWi6VkiLcY1rZv7iUS8JJU29YWp5ZLwWfKcf85t7IQccfQ4yy
sOrKQxnx/ODMQpBx29vi3/FGmoGJGVQlzktXtwDO7LEFVYZvhxv+sCOZCE/oZT5TwTd2g9z7RN/8
TJOhqAy4oBnia478zAvWLijfuOu2YjuHmXGaYAlF+Q3v2q134LL0OepxZLtWnleFUR8D73w+zVrx
+Ir3bHIGwSHsJKcRf1bZlRF5OgEUflJpsVWtMhsocEsRpm29aerhFxhegwNYayB3Rj4IRZ1IDirI
UR8LQY5Oc6eQnaQGi4MhSYJSqH6cbtt0pm1yBwXXGC+2xyqNY3U72JlY8mE0HfFQ1NKC3QslhH5+
pbDTTDDwpLmCBIqEKRMi3ejbGKQIuj7Gdts7tRzAdwiccvLL2Y4rZwuKHpbrJFOcbyiQwT1utf1f
QgqZq7RfixQ8ZVOnPnC6eJtNLQyxk03Xe43F8LWprxqIAei1kRfEKCg0CUPgGJ+4Ph3sFM2Z9FUP
OKPVz0RE4bus8UmVnayiKh4PZ70taX7Gkn2bhL3BOM0hAKEZeEyXV4cFli6iiep6YNmSt2eb/JRK
6f24lO7BGHom0N0dtrPGYf/qj/noDGtVh5x7Nbe8WC7/i2xkIE/PlSb7AEHfYAvLfvScqQWOuHDZ
7WpWy6NQ/VAYUBaFL/+Glr7xOYr85JhZEpBntAViUgPnHXoty5maML5b7s3kN4aTuoi+DPVq2qS7
dCKfb35jOX5osGcgDNRgDO7Puf0gUNU+icYMbugkB1IUOGdLaqyN3T1mrjDLq9s1HrO/lXvBduwt
yAkm4k6pzhvYzwq686TQv5VoFsxbJt3Kke+24fXJ//gJ3ZQ6JnkCMX7D74M9dO1V2kSJXHOM/g4+
gqPTKXNdvAmJ8zsYcn2MKEVaJw4abruqbhg9WjM+7kP2q74JFA2JtizVuzobbqvWKmCJcAYBiSlC
00CDmWmHMhgSs/Ma1Y7u6B7XCWpmEeEn0Hyw+MO/MZezmZGOBGRxIDosiF+w+D7W+LoPrMUe5Cff
uxQkHMUHuQ8nTDlIG7AC9cCPw9UI0UuJ1jO0VeoZ3E8iWeNKieoBFpB1eDW654OhompzsvQqEyE6
xERBXQaBOG4L8vSnphSuohVEriBTlfJO55xGMUuWfMvRYVnspeGMRpOW09L5RV08dXIC2647c9FL
71BgK/5wByEljpr5vfc3IkEVxqjJg6E4QsWx+cZrkY64wHSxY0yvS9SVsb4eQwZt/jaiETXCeea7
WJzoYj/y89KZvq3Rk0+qy+urmiYioCGN3EgSAujWxQxvKPIh+2fthaTfJhDznTLMSCZ5Lk5p4+tB
bGzDN5vWi93GQOojCy7fZaBKlWx4C8/tGNZ2JcSrmBO2NZEhW00y8yU6vbZ8JLwgpYvkH1JHuzpU
iefyd8w9Qe5xWrGJpGhaJOL1ujdFJSmsZl09Db2ks2zeTgSG8ZFnjyAmXkhATyFB0FLeK5GIvccm
jk7aQxz5iYGbgKRQgoEDa5RH/woEEaLCRV5uQZ6oOdgifV/VkyeptqGb6s150ndfdTwRTVV4Rxq5
XWu52CnFNH1HTH1ZXd1Ltiz7RRIW7es6klSzWc0qp/D5Z0cIrLm3RsE7joMXvJT3867xkMvTrEqS
k07EKT/ssfrG7IO4SPacDnXsK56VorjX5IgXw9QQ51UlpxEnvsG+FPap+x4dDo1RxOr9UeiAvAQC
49U24nhzN2ES8vfh9PyM4UTbbjkHESaXQXCyHOhHFEkZCJZJby/6H9YHw8mJYlkUq8T1Dyv5DyFH
FtWs/UCaojm7R6aJlehgs261NdsZhZ75xloQnCVg1WsF9bKdlINp7xMntlN3vg0PNXt3BjgDncBD
EeEcMdsoW4nBNLrxkX5FDZHAuWZlDJlXqjYNpB4LCvNShuqZb5CyS3w28iLbBw8xe6nYkoDG7Pgl
dns62v4H1NxvB8n6buDQyK/qwbiEy6dMixPmDfDXUrBghI7fcHchfWfwdX/dDERhDNsRzh9/sN8Y
PrClEaFEkeu0yiwP2hnQD26iXWp3deb2P29PHWg9uIpg3dMR7sbS+qjox5NFUJ3QlQUPUFVjhXrv
jerJDqEZb9NKaJoglcTUA5eF9F1Xywj0XxFUfrj1i5ohJvH4KYIrOKKIUWPXhCIXqHu8OF348yb+
U6OB3lxe66hcRn/hD4hEXQyfkZ00mvoRe/J6Kp9CT8g6Q/SgQU5APCj2ng+l5ELT9abuw+Ueq7iC
ulqE7GXhSrApPgAw/FrCjBsvS2CHuwpvPygkvAmKj+ord7t/HiqXY5V2SUs0ZEf3WPZdx63WYyKA
z4rxi5MFilHkdH8dEGmu2KciFDwEQMsQNKJ11gfmUXo1G/tktnbkkdz7KuQDrqzD53CQU6nD/ynQ
P9aquFrRL+hbo9LPAOzo+RS4GSn6DwSue0jLdtK9Qh+ME931bK2VKe5kNJrrY5OEQzJU/IdeiDYG
TO7dRZhIjb0pWFw/qcad2tiVUJTdA7MaA/xR3Zvys/Sh6+eGjw+6mubTLsnG39pIVQuXh7SNzJ8z
WKO4aWMSq5Ob/rOWBVpSP11LGmOanVHec0AEoUuzdDSBeyZ8eSiomrtFmOb6DElkLYsWsp8Z78BA
z/2/RMjxsfawYa1ZidlTYaCqyt7+YYaU76DBAUudOFFEkF3S8DXevABzfI1fhm91Op4rQplqc4hj
gAGgdyamgVfGNYLIoTd0Pn6dHQMBZa0u/eS7IIgMBCRNIldIs4hXvXlBeWMVz6kz268hVmYTEOpF
MbYOtpndijETHE4JKxYCiLtWIPjtfjgAxFRG1bHkgnVcJB4LusYSUlueVLRO92okXWwZ38l7tSOT
trQTbOmhYvX1TRcuC7Ee8BrKYwgRhZrGmNkA5CIS5/Rm0X6reNpqAfmkETs3B1jW228iMCXkSQhn
uhPWSmbFjTYeW1Gr2k9ZeiihTSqznN9PtEvnZGczJa/sT0Xf8rQpgU3S50LAg0QlSoaXhQZfiCo9
4y8PpWqjI5QBzLRTO87Z7xh8lY8V0uT87bhL8Dp5bNftCOJzz9trfFZxtOUx1MkL1VutcuyyX6jS
aT2YtBPdRXMbR4Nkef9H74+Uh3UwlaeuKh5z281QxtQPT5u3E6MoYwgqmj9UDQDKJvSRBOTEcZFh
mmA2W7sRB+4oxG/WSr9LZJwtOa1OBrG/yoC5XyWQDvyWGPHzIEE3RXyfUggy8+qvSxqGGRlTNrIt
gpTifhZRUQMN2r1FikVRdRru4nWMGq2mgoTds1DgYmN0DuL9E9XI0Xjjg7dJx9XzMRoLNv2JGvoa
cVp9GcvJcAAOo9WWS8+Y5OZ2FZEwUzuHBC+paQoFfn2paz2WYgf/mr7tv0IbYGkMAjJvxzR7p6AS
Bef48cJbvytBV/CRvy7IVhSZCIa2GyUF/gBWrzEkeDgxajAyzqzNKVMy2QMkBigDsZV+eHoCuKc4
aKlDphjJSUuvDB1EM8uUNn5eIxfYwIic+9wBTGaC9uwVgtrs65yBBVvCIMNQx71k3koupNQIe+59
HCnW+vidJvqTcaGfKb3dqILhnHQkqzAdLvQ71N5RzzHlIEURcI+7WUpkeUbtoJt5w6s+7FwkJjm3
o3Sxbimtx55/s07t66WljZJFFFHN7rBy19GNvzjc7xmnyrNtfYv+8ItnUDpMgwnsUXGQgaVrBXgM
yAecKaCrGsp+hTgc7TJhCvcux8/s0w0cRtGrYZqPVYy8dnE6ycjTjONDvvYJXx3urmcMRHtbrwwg
fPd7ycLPF2HZeZMcHVSJyg2FxD/QJCjT6P9rDKLc6EbLt5YyqdR7iLQu8Ih90s4QoTbWufJgK+Fs
aIL1KgEGcM3xO8+Llmdv6t4sI5hALgCIVRyBtA7Xny8p7PgYmhuLpXUR5W6OMdL83JpKK0fHpwk9
Fsv3tcci+h/R3DpH/vVloV9m6X6bL9pVHBhZrDaMg88dQ+7JvgikRkwDfwN/fzG/RRNdr22q4q36
6b4ayd0hmRMEsYJLlC2V+WKLp+PHWfpxTbRJiOue/mLOVmoyhCzsNszCw3MoMEqJT17KJYEAabYv
4QR9TrTJL4EKNrKb7ajPVEpMuGTDpRVNq2Hy1oHJaHYB36pQC94paq+79m3V4/dyTte+Im/hEANR
Nk1TRTJ4pRC3ikRRO/DvQpL3LRrLORqFq2S3a2LaeKfI5mbR2HKTBJcOcGm95B26PUfsr1q645kF
bKHCs9hF0sWaRz87e1x8Jcs4H4f66Pw8bf0AXbSVh7pd5ITcUbXSS6RGXBJRq5CgRs6zzNZ3ESCi
Xh1z9rNaSFkwA0XkUf00ULCaEqysppKyTX8nBoH0O2XCPqDBAOd/KSRJoXfQxydn0sfIb3jVCbAh
BErrA3mbgbceylrL9174UanOnTRAe3h0DPagYorDSHJKCwsMyyU125cY4Cke0x+edcejK3NA5fb8
iQfRIHRaNySxqc6m31aUMIq6RJg/Fjn18xc2YZcEOHZqtPUDleAdSiPALhoQEz/syrum07tioD1A
xizmUM7PdgFSTaxgxpIp3w8tyozTk/mR2xpcCxhErs0y+UeehqXCgezR6VUD1nYQOLNjypLkAbL7
kMeYiQsj+fXDAZz3ymHXbV5JGUJCO2BZMtqqs+GAjwZbr0NzLnyY+Q+TrWYuIroZ86I0km9heEXK
XjhIm1WnfyV5xLY2NfB6BV0lhWSItnIRDR7ZQNIB/uoXl6yUAZtBK4JD1prOuLHZ6ugbEmQOSuNC
XHgIhLZxqD38YKN1iZc48PTJgpU2lhSDwrHvjdUP7YHRE1YaUMimI6v5vMXVkPuNfqTZrV/74Wqe
egEcPJH6bmDW7QB9hTe0LoE0c4edb1HfF6LfMecKwlvfQHi9C99N7NDiZSFfRmnXSdDGCOn5HjB9
Dm4TWg6QrPD5VyqlxnkjajpfGDZWMYaicMPe0tAlwIjFCKTKtIjK3bI1yErI13jJSYYq0f/99OZt
A0vq1Uo5eH7ZJaqpuBk/Awrtz6fA3YDmvYqNXI+Gp6Gnan+3r8amvwP1ICr2gSlyQ+FL1X7J58K1
IzAKUnFCXyb2IiELEd5/4ukk6kavcGh0/TAkpw05Sre57T2yuyD0eA2WPiXugN/AxTSSVKYUXrz9
kCo8tZpCd6TzP1NmDYqCJKkcr4516qHTVyK58M6p4Sn//BzWHU+tmFAOllpKqG7uAB5z9R3aMkFU
TwndJJNNPcfb7ggaG2LNK+dnEXBif0KWlAQ14O6z6H6pM7Ttp9ktxcRJ6M9VJFruRcm/B4f/zG6J
/GHpV/7q5tZD82FKAzvf/shQYFewNAaIGYoMPGVMD89Vr8xUf3XDvBi93BQgCoH00Un0nUet6tfD
iqljufGD92zWfbOu6sbKKyEETRPR8VbeZt1LJIZDIOGBHHILOgdIzPJXwhjnvONL9OqNsJrNnP34
efWLolF67BWFwTVnECCCXHKpDjswMs12d71vMrINqKZ4InFEEvhDAqSiGrWu/pHC7nkBmXTsZOxs
0cOU0EZbXcnqCxZUYTajgrctXd7mU8E3TfQf9VR33Dz8lxFq0xdh+deazz7p+AW8qws2B2vAaY7B
gflgZFIxTA9IBB2rpesXZ0ImcojDoFMFHT8MLcWowwovoQ25vsh+tK7JqPbxsqAGQmGnykUMxOrl
/TZRz9NplTedqFKBMKn/EMMo7yMtaRDx+ZNDsRsIQ0sqffgjfgDzkbzSJs9TMTqoHkKAy3HP+N5k
e6mXaQrG+BoQv1BSxn508Xnm0jYO/tyJMZDIoSJ8get5s7dKX4GQHTVlPvul7fCmMjJrM2F0fpTa
IOl+6AC/fjesM7DoYtYN53R199Sy92IpkVlalT9ySFLbiif1CLlgdGJ1vNeS9y8MSuroq+/5CUzs
gp+XG44jMSUxJjdsMH4OUqfA8uwxm5YWGmPwyVOqoGMbxVryYg6zQrIshi7wEUXNLny4GJNFezqa
PvmOP2bH+iokio7K9IWZ9Nh86vX1vB2YsQ0LX6r7M1Dy6GS0KmfQgj2wtBzvOTtQbA0IVIOmr1LG
f0AImoczcnXQyNWvpKV0k8JM3z0wsvY/2HRbsu/jlKPgXGJlmWb8g4G2v4qD8GZA0q/9/tIv10g9
MIUFrEUxGnIVl560+Gc1BNsQiAD9t4gjUnjMKXEokSQpmwmD7v3LmPL5yZ9MECvZePVqtVlXLiic
40ddmgn46QPp/qA7hyC8i/uxvVQ1zHgBMMfL+tpvjvPYCGbCowqZnv26k+ug5JKD8wgqqXwth8XW
rfIn/JZaiWbJnB+5JsgMJnQlyu0IxFZbrobttEGntgGs8FQwenyFHD7+08Ol8qcNWRVvBxYbAXC4
PF6XWuc8wzMaIftn78++P6qAfg6sXW0EcmgoFd+CuROK1Igph2+o3hgi/zh2zwEHh67+lGf4Y8cY
ihdbsDWdUVUt8emg2ZGwXDxQenkPsUd2Hy/dGQCmIUjIOhSQHMBtEEeacdLPpeev2RC1MVlPbHLH
2YYv/p/7tnct3vsYS2p0rQgjSZ8rAtrCmVwxgxFdUWVUw6oYcb+XWyfDy0bkRjCs9oCC9vRa60nN
psTPGIVwIC/7UinhKBtsejlMiVX438X9zzbQ91fbmexbDPvddkzqDNsvSvHM/lHu+tmqMtNesYG9
IsyLIydcu7OScVXzkKhNRAav2sqrY/qlduZF6iNzDWuRkojRJF6OOyeAU/uIwsB6lMSM2KoOf0UH
Jrj9rEr4yhZ1HKOwDdvhkThxadU2bjsZC40MS3PoAPM3XC9YrNGZnFn4bLkx83D2EF5fJeeEpz+e
W67+TegEQwQZfdFHNcjbvMysN3IZ02trxOlH84fG3YrWO3CslTRZKOkGslcanwauzp+sSDszIsPM
OkmeIRbLAa0uGRP397KyOMT8W/LWwBj9XRhHp6A9dQVzfWDKdFjtwDMYqqRCHfSfEQSrSNIiMLbQ
IVPVCBF4EqwmV/DDMt051dhd2oEpmWIS+X0xFh5vqr3AQl8u4Trs68FbbAkXhcAqzZgd1sWo0759
vsrbo7fNX9/xhz9cSDrA33UhCBMVbFO2Bfavbz2dRSIqiblfUERmmZS2ngWv6DGlzMBaZloEE//Z
YSK3B1DDxWEOWUk/BBE3G+4mazxETGvLm37ybtmjPOSdpTUjKLlqlC4uBudAXL/9UvjMpnZIO86y
mxH10X4HI+MI36iwq7MPX8EliTIx9ohGnQWMPZQcRh92uEZZls9ttEsUUvj+tkhUQaHwsbjEL1Dd
gblphaKRfIYD7ul3PKzPwqqAjdKQ0MSg2bGPkHnBv/xC4zjdA1nDxWLPvtsEkfFaLnYrL3PMiJGM
oE44lgrbVRMCryri+q+oTGk+NGJVfJoSC7jmINwEvu1UGhLHUGpBgrCSKY+PcgCJkfpIPn4BsB/6
CU5O0AebA5t5eF98YSuIjuKjLIo0YV99HZmJEtZ4chJ1UkgMCuHXMwHxJLl+xy3GnyLbYdK8G3pv
DgTnkkJy2k492yQx+PSBkOJXi1CLt2/8c22zulY8ijsnDOWRZ4Oi9+a5Lq69BsPebP0eN5rxOjiR
K8Mo89mcoCCnI8OJp8VpmTwhO0HOeherE7EW7+r78RJvIk0nTJRa57pC+316PFwMdRgGeFHWZxE6
Rfz8E9vlZBXn8TsXew+f3PCu+4JJtj853iMq0l0QznZKA1HPTSVDDPyXhdEBRIGkrvtWhWQCi/ek
PvT1KOeJB9B7jhMsZpylT2NZzd96XHQWncY9KZlBb8svuKHWJYpizHoy1OGCOc9P4l0ljWKIYe5I
rGuJJ1C4DeKPJFdZhG7Jl7XNRz5fdiolFK26gNteQdIeWe+36Kgwog069j4FDbNR7M/IwjU0pyjb
gqGO2K9Qky2HmrdbqtP5TubUib6wpGQLm65ay61s2zhOqghCoSa9o6dipgTsiXgH+d7+9+nAAHhU
V+dNNLXNYUXVZ4qqaLLuI/rJ+Uys9byznLy2qLQdfinZTtGVE9BOvL9ZjS2Mb4HzLteuyk3nqe0O
mwCU//eaq96RAjuHfW7VniI9tN3s2cts/wN3n58KGxr/tuyRC7Okiy4NsBZFzNaFMJBHkUDKz/FM
YkBES/kSWVUEqZpKc+XbKS2vWv3W9eKAjmX4nTPo2eqrU2JLOLDNPdi0nlbWq8/Ay8rSXIQ+i8gN
qextw7x6OYi/kZbwxu3iGy9ZsrQ7eyoFBZ8D+QvTfRcXbhs+A32SfgfX+25jA5Jw5SsPvhHkMrgP
NIuQ+pTHeNDU7SdSpjk+oJQmUYbv7Y8nzNDD4styQNognFIOvaPBxkvjkQvegGCpBhYPOuAAW8Wx
vrvJynEqLk3pUJ2gktsbRbfpStLwVGL17/iJJBDu8yoH1eMfCBmsjUUC9+K/N5RkFu5AsZLtSn8V
X/KlLJSpvl1AHZzF5Df0nIrd8m0Xnce8XkIrujTlGbLsIghjQuBXndzSU/bvEI9SNfrGcT63MX59
2XeNMAlCSmyHwMhNCpzbrqUfItAZk6MNxszBHiFiXQ1Iui4Hev6v+i/W3DTrkCMMnHfZWHugDgi9
/Zkq2YZVdZZAcE8x9gBuEAJgGjPsqPXd/e2e462fIPYs+Q6INA7n9RDo4b/Fc5h0I8A2ruu6cWBb
u8nh2k5e+lKpKQ5d+87HVB3xibm5dfXv6/lrD/YHtsr8UBQGMVnrF4NkX1KcbApgny32BzSTSWCZ
RyprGg7b5Wlvs+50xe8J6VSJkZzDDEHJeUgOn4C7xKvVIgR2n4blqyzMZSsWYuENy/J1KzcTWIC3
HMFFdnYREK1YdWZhJfSx1Wn7HvyGez0ckzkpq0KX3SVDz5Hs91S3+E9CrqesdHmiU5npmkuMULW9
lYgrPLpY2fxrqFmH7ktZYyCO2b7oiIHmVEn5VG/sD2XKh3a7UJi7ydIZ16ZbIoJLXq6O4TjU3mbK
lzCdm78OzFDuB3QQ9PDjQQOtQkxaUu5CX4cfGterJ+QViiyQ4YkKn4cUCGxXtqw9LgoIaFffW25k
bNVu5weVYLNGkYN7TwfiC1ohJLDJ83ZC8edlQizSOJcDSIPfsETjJZigw7MLE0xuIjPd5la5l54E
bMBVmhh3vCrEI6CEaGRL7asY9esin36Q4uu/lWsWRP0qtBo8UiMFpb++euZc2A6/Ovjx0nBgPQuj
i68XgUCKLUVBJrYNh3KKJFXz3jWQslhEvpEDgdc/kPCidsWpTB6xhKichCTKZ3JgM99BGl5gq76/
bfgDREYmtPM14MW6jeNe41hGe5Akk+SSWohAbU7npSJnte5vvZOf/C4eZw/zGfiBKlRm/nD9TlG/
c2GTAFP/C/7Fb1fprrH4f0EfEh0Lk5KepyiiBs3+Q9jDdjuqaSF1Od3dDPUbJlAoI0UWoPJ27Bb+
5UD9T7zsYoyjOy3XwzYwhkw7v9fCIc3L70y1n15QLLlZlIGftEwEk/Dtv7eylOqo7R4BRdMXjriZ
ydCa81wTTrXSEuP/qSEX9lUH04JSFF2laQC99N25HvoYctkqFfX7QKwzg0qf5OzpPleqLVC8EaYc
tHawDz9RsfapR8vIPTErvEtL6TVKbgea0s0KSjhuwxRkx+OrRjZsUT7uUeN1
`pragma protect end_protected
