// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
B/7f3eeHDbzoGmxID3myRcTAvxowvjnkU3J97/K99kXf8zTMMaTpj8qOxJRg6bLhkiPcCthKoGzq
wbTY1fZrO8xwl409EPpE/iehDjgOBm9uKTQZJ2SsJEQDhVd1gTiBxNumxaSjRswvwKYARyl2oBry
GSY/wwYJ2kmZ0RF96WcK0nPAAPym6T3aVMxTzQrrHSQ8yM3Fl/sN7iGm35jeXRyiwsWqRwh+SPd/
h6eU9ODo2eFKZbSI3JVudhUjKFlGlaMeAkDMi7qP88rJPgaT+WMA09J4uYolmt/Q1+PYzTNuDn2d
jZ3Fz1BBQxovpI1JONOVcTICySeqgZimTwyD5g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
d3Xhpx3qcvinYr16UeLpu4atnY97LwaaXwiJWipbG24kggDzPsVF9wjWhlDNwyyRn5akhjyBWVAE
WcheRGLZwBmOFxVMyNkF1yKJ7KL6EqmYw0uXcmC+GVmn9HGxTTT1vkcLgHe7VULvUBtIrhmgMoPo
Jk6sdOQSKNSqyFYKJVAxglLA/373cZfoJrbug0QfnEvF3vdOtmiajNfFSGabiUsnakJSUOUP4/Uk
QJQLsPjFRB1d4zrZNTZEhDLiWdRHSckrjsXcBEneQ2jMM5OBZyFDMs9j1VV1Nnhw7Em49X0gtTC7
wf8jjmcx5XGay/xCpbQ3ZF+QZLjLaTfgdl5eNfK+JJvjS1dy89xaJ6RqSzLh/Db1/KfyzkQB1QHT
47YyNRNegT4oUkwNMKmAX35OSZmDRyCCiignTvRSOJDfcBkdwUwcUzJowMiYVGMw0hBLqzb17arc
QUXJGCCMC4BlIeOKqdfDt/wpfXTk5L6ck0d8cvujfjTzKFFEWE07AYd1p49WqlcHhxd/wGhfumxn
sghIwfucSJ0JJtjJJiXcnNm/Acb0ynyEda1bv9lP0QGOJpoaVz29Sc6HC507CUqwUKh+6XFEOLwg
xT9ADp/dY89pLCPdlloKA/VHgT2Zekcwpmcpc8C/lMtUqXUTvBF6BMP/uaoob3D1BBDvV2gEXlC/
SlPRI5pRP9bZuytCXERH5Uaoe4lUB6mqaA0SmkU+fNPycfPbD+J/v2DQPGvEsYLxPbr9TvvljHFC
zg/xj31MNw+H0BKY6cHHW5ckvse7H5Fgc18QSKFq6Wqi6YO6yM0u1C4Pt4EY4Vwgoa6ebSaGVqhi
3V72AU2QJaGSPzQzxgItXHyJJqauCD0pPkmVcIi0iJq3oHiq13eYdOys353pMc5OaQcG8wIOZ84J
2qcUbgDxgtnRsT3tp+SjQs6enVvVFAJGpCUk5c7j/lQ2mjnS7k066Bx8bY0QDzHF1LAXKOJb3Xb+
/7/tJJrdJBXWVl9MfXi3l25cb/v2hDd4Hnv/BSc2dZHLpF7uvp9FYE2HzLxPaGRSCb5VCFZDtEx/
x+zMpJE3uQR6SmBYCcclAKkxgUtKSoscd7ow7CZZn72jyumoSUBbwZhgYcffOR1pe9w4cEHha1cy
6ept1N6UjYlrZYI9w6yye+7n1tlG+vmUfptcj7eDJALg7uNlLFrs9+bWwNB81emQoFAWu44g0JMy
WaLBEmfuNddGE/j0OutqWO+aGTAYYPaXSeiCRfUDo8htGmjSl8PatTyTEEQ4cpndolbG0JlJ8Td8
jcqsGasKPdfyXQ5D+zvPHq70QPDeX85/oKkpvnvmX0HjoeUmVFUALxBs0c2vc9RjJGTNhQAHvHvC
ria5T3DEf9toyNtB77S3NVyZ3XR2CCZnlElfjA7MF0d06u0YHaCSpgd5Q9zc74QoF0bLcTf9eX0R
DBfFspG441RvAYZUudfjQjON7M71jQBd4aq2RjsNmWSrjt3g7KwOwB+53FcZPAnSItk2ULPNpgCp
RBCs0VqSpeyZKHmu/e2D0qxpUcpmHCu1UuBQmxzDp5jWGal596tRaekl2Qg3KxN/zkVxcxZkhMsO
DneEBJeixuAS0nTQvcB+ABHEjBOR4/Gc50nPeGuTzwHG5S6xUWniQH7USJGBTGs94VP81/17+rCA
cpdy5xmN/TzTSLl2qYJ8M87z4g3y5q9O2ff3y5wYQTG4Uw2dAA3jg0XkwjmEDXVZMPOCa790HIPN
oyyOf+r+MC1ZQsDZWhlF+3RPwP6TuSMH1F4unwCppZa2+4B9Rwlx9po3/+WvBUXO2Zj7k2lswPl7
ry2XS1603ZAg7RYSgjxOiUsmr/SOdY4V8lB8WZGXqxoD9UOqP5noTau9QVsaQyjKFXUZxJiClu4X
XI+BbJinTg7XUnD//7D1Q7W3ib+TzBSfS5eY5RNEKz90WA5xLQ4ZSk8Y5VUKhMghiqZc5/0Fg5nw
5PCdx2uKanlzynSozbq9hw7vE86OpPKIUpr+I1IceXaOrWfM1NauWYiAiSn9U88aGINCkj+3CjHA
iufrorw/SuyBUx0QS+mKWIJHnUJhkK6mqQ1rpkjqUTHT4JXadppCUtSTsQatwwIAoVOWhlEDoqD9
giRowMDBlZVQFLob96SeFAOQlVNMO0PhGsmhqtAU/NONb5i9Mwda5SFPUq8XFGUE/DpKJHE1oQk7
Bow9grVedT3kX5dQYw2k9+Qd7bzB6b9ZQ3ToTrRxt6itepH/KFNX++QQ7aw6vnWhe4T0BJ625GQW
CRoK++xeP+Mq7Tgv+JzqU8wt1hIkh3dVU5UyThvuRGv4C5lUzMkY7PMA8bc24to0KYlhvfGLHxpU
+bFHrEIrRsutf49r67QlvPdDggdFj72db2X5KxbEzlDtRPdzRe7GRGvDY5FGz9JpaQaCrqHIVULZ
K4Ou7koaTRaVSNBuxjHfsmp/MC7n3l5FgTXo8PyzCTaJjf361XgsNvczHi7b/de6nHXV/1rbE0+8
dNlV1NmUo142BrjfTq+PIey6ThS550YFvaZJRDWu65qJCKDEDQipkZh+KUuFqoVj2FFhMHQ5a460
vZYvEIRLSBx+i7lARv6BrEBfnUNppQg2nZ09XyrHF1MTcAFguY8FIV8zjfP/cSFg3MYDzEkZTD50
Bgo1qnkeUBNGtwTX7UHNJk1xHPsa4pnC/V9QsVvHABeyzp8BLFn6aJ3xaRJ8Oy/R67MqxBcefCdK
T721t5C1iSRRbCkoGEGqMJ/kZgSUCLX+c3Q8G0NauNcplDrDUA/8P3GK1XLHHBFVcT5Se+DCC1iz
iXxg9OAMnEb6n8q0QBSdJPaZ958o5CJTiJ1eeJy04cY0jKLH1JXBf0lAN10Wz/P77pnQFvWEhucw
z4zbScWqh68ogfVrgpDr84xt1Kwm+xZeLZ1v9LDZVCCCiDbBRPoM9oUEctWkcQ+ROaM4ciMA0h92
Q0epFEgae7UUz2U8AWxvShSFkOLouXsN8dxeU8Ho9CZTtBfSYpkxqqd+YqBjue/lubYEzDdkM8f9
NEngQdlZ6KNfAwCAvtPqWeOX/Jnqb680cHTfVxQSoGCFIqfjbsHZDAYIr/ou+OzUj4h0YPkeJBOa
rSGtSpvBlbrIyAPvzi8xdVWnKtN6QALmOidvkYziaBFoeQcp3HoveuSRyeOSk7E1W6MIx8sK/nqL
0OQtThMFRXgxvRVmE1DdeJdxC2UxBGJAeXj27Ta/5FAvDklLTg8OdHVVDbIDo8/Qk6QK9uyX19Gi
X1GcBQYiacsGR7BJL3de2LhwYsCgPMpTeLSxgtZuW3n3tX5gXVT+HzKwCvYbly04NjvVt3AZ2G5m
Mycyp0vNMEBEA6yLpMweeAwReteu+LmM/5cnacM8ca5AbZg/xSq/YkmZF3hkt0XEgiikpBaM2Hqs
Ko+KrUD2s62bex0zN2FzggcmtHhrcxr4x8GCWL01pdTeguuDbC/aow5nCVoG9O7DwxjCQi+XEnuO
/vOMTtIiY08tmPNBBjQRWhd0iHpnvqmAbTRc11hrSmEGoluItPj1bFKDHTmq+1+umwLH+yiCwSyT
ZDE0ABpTp5IsqQ8pbV0HdMHl5hWOkHZ0TpK/E11PQdCXPwVNLeG4NA9t6M6DEuGFeKDsN+2ho+zj
++Zgv3SxMjmyggeObX+91vRANqo0zDgXhYYOhr/9tUpYACfAdniNKpLQOYjMtKNAei+xxOjaIIUa
6A/+frS3GK4v/Qp58aRjDMO7fuF/wmH7yi9DJ+lKaXykWdNDXw/VeLBXeoGyLDx/HK1JO+MWC6an
L6T0cTa2N1k4nUnR81HU/ZJfgRq0relrWwBSPaoxKEt0XV7BZELmurQNb9gEnDOYY8RihT9m1Nzw
ClCuLtnYdABxo3VtsatKCi2G6mbLfD8hvn1kqQ0oEku3XDyBUgttrmnDI1zsUHZHBJ+3vVcVEEaK
Hfn1oCx4x1/5kM6FWyTPwcnOJbxJ4n/QxdudBgrfej/4FRIwsCCyOhL+eExKY9DwbtDfQRBkG/B0
F+ZVSIHtjbnhWoR9ckr0kIXsbcem9XCIaaPGcI730H029MQZoQqAfHr/JJOWmVG4Et2/xhM2zgrg
PDEsXIdQR4Ldo8V88713rOUZvNsCntep3tr4VzVApROXKr+K/vWvpMdEjLx4UoDi/asL8BBbNGRI
exYe/mxl1eOcl1fhGw2GyaOFBD8h1/TRwhz4RIPoaveQ6kXjUq1Q3rhFVTKBKoqTxgTSCYuPgLRT
YN3bCb+wkEAa9oCxQWJMSry/LyQPRN0fRQZNxzmVxbjDcIl3OZksZsk2rjmSXhvX1Orw+Yr223eR
ztx2tfUpthBVJ7NoliSqzBx0dc/i9Z23MdefAD0RYr5Z9f1I0aB1x25PXRRUlU85rGRCdmPQTVKu
m1B6bF3sJ/8MrMttyK6ur/M5fr8Utuz2PvXPp8AOCJzUTPAVujQUJD8JUeG5TuKvG1lttbkA/KHZ
uKrdj+W3o6jZtBDZ/N7PYarIRXHXYrwMe8Y2OZe5+P10m7NJ6v21ZOckJKUo0vcDQofGPl6SDm/l
So1f1Q2hFQ8DcMuZoEgky9o2XTym1yKCKG9owmsBWba61m73QThrZhqRlvLKbSJLHj40cf06RwT6
VlaSmKpLPnE4dF0bMlkR2eHpxzUIJm6EdbEtJv8/5GWEqNrHgVo/LwR6D5CIDUi1YaNCSl59a8cN
LoyIpfPoMTT4rg0o3DJQzY/pBTfbBHbapAk7Xgep17uIv5m8KiArHLo4earQOvxonjP+F6Q/buJu
8T0FoCEt06Ila15z2rcKym/yry+0G6uSeayNfcJHcg74IXiGuRP90aGmdf3SKxXHwwgU/qTDjJgm
LOVzfgYAAfZD3BA2NCiQTkishdzvPe1aKWrVKywMG4ZMoXkRTpows9oxr7eeysKmSKsLK2Q/umDj
uwcQECBhh7TvwGK0cN4jsq+oQN1WLjRoWA3WfFRfdc3PsmGpKUpLgNe4ZoDvNVS0i4RY4v3FV1gU
PUhAv94WXqF1cIKCoN3Ebxmq+v8iXCqkznj28SnHJdNPivtMyVLJS5Gf6CNApxluUqLBwofEzuMa
4VjUh4LRcl/WbhxlEJAkOPdEXapRywVR2mhAbis9ke+OnirdLZh8S9xoQ7mk6BL06V4j8lygbivK
MaWvbvtOy8XM+wAuSwiq3nxaAZPtnVpZitqEda6qtS/H81NpKhBXYwGjbrA7LLfwD6FNRTMPMhoP
s7CmN/a9HTg68wfmo7WQcQwtYbvxF5ITx+fk5mL9pR1lzzI1xzsbryhX/Ksmgj6bUDf1HcyLmPdl
/NUWa0/5S1ITcbmJaXruc9v8aWxQweNvO/ZWi2IjmJVq9po+EwxqOybtW39YsOB+dSJAFdTwQVnY
lCwjVrL0ZVvS4PALERLBogaEfDfuUcCP7i2PXEC2AxeDPi/8p+EVnsfi39W0WQ6+tVC8Vi9dDibe
w+uyZ3RKpz5L/v6/fAtwgLYA4cNw3JQ0DvMGsXgWgJPX1Og2arsKG02HW005r51o5RI5gimD8MO9
TFnQJIrNb008pzbqjK1oKZ89qMCdXwmFFhqGM81YKXSbJxxOZHoCw06HXt6GtC3Zm42dHFIrqjwa
qw4tRNXMmSN9uBJZ8x7qZlaoDH19xttjjhBFxdsApWTqK7XmX6pk6dRxcWoNPf4AupJRgpnKLdUd
IrMfiuVRV4y+YojNLsqtTu0EJzQFXDY/bH3SX6jEDoe3cKuIYcFU/JWjNVNqvBF9ZyhZ3CeEujLl
SdZyg00U4/xQrEhOV2jxM8DYpWQYL2pqMhPlyXb/GagMxKYGT11ozVMzoSM9aSpLRFAWEMQ0PPHj
KyqW5AEvvIx8aD8cXaoHgWb1fN5LQQJnv4nyarYwuZa7Ty5nh/vVZYZ2EIpDpPWMOl0Re5/h9VdO
K3vTsXtt0qPa6QLHrt2NNTMnhPhhwtiwdk3PVRjLSvOStsCxuEeOXCSwIfuCatonsxNnt+ldD6/r
GkE7hMSN7dCl4QrwP6i4BVnd7L6a/KBjjq53/PiIrQ47uJJvscS5uQPidoYwszSNtZ3sMw+jNHBe
cjDQm0A+llJwjLqQS3rYuqOL8aF+jQsAsYsWurQMGm6SY2A4Ko7ete3J/PD5PGDS7koOmfpJiquw
pgzBTOyLIeCgDsIX7AFs8lmwgPiO2TChReLvNAkJMs4wobe812kX0YYjkJDfIt7rnaJM9lAoMQWS
A3bItS9qanRHrxjKkcQmwom95BW3JaeiY6Q1ADWeUWnxGFJDU1L+I94qmrUuj1eY71uMFGXIjSgP
gK+3rjBs+MbNmTwSo/kE741UANQOgwoy8Vqw0HCl0NOCWJtmHXmlGEFsD8LHGoHXylK0K2XOJkd1
GQSYpK46KiFFGPaY9yNNR+ON2ErQ9lBlRfFu8d1xfvkvmq4LtvzYLlD+cxHjmWqfgB3qv9BOBr9W
+pnAjqDSoIL+47KSrlrnWp0TuPHS4y3zs+CbJpq5Iy6V0L72voR0unuNvjgKXZ4DkPo25IpmAHO1
7FkhojX/zcVJ3WW6tyrw2WXi0yyVfpjptYr0D+d10capCq+o55WmfBLU1eOCuU2iCJbrDqNi61tJ
QlCRhEKEhFRaBam43qLp1sDawn4r362xvGbUMHMd1xkwj97evrkJvR6I92Ws+Hl/AZUqX6H9BN/Q
yqvu9O9Iyl1fN0X6yJdWp4dKXvOdb28G9efdbqC7HwfFAVq7xL8e5r7D9XcU4CdMrgARlyxnvHLt
UA5IZj3tiCt96zwtREkTxKsPZZVppYwPNy3amdsezCdJcM3ix+/ebKeR/+3TURQBQoC4itdlvE0q
zscqkjvGhKcwFucIDXMc7/pK7fla+RMGxGR40dOmNpqg22uWiW+RzgPquOxcZg4Y7o/PxiYKCzdr
VaH0fTG9g6d5QSXn/T9v/cF7j69hRw3wMea0INkNZh136NFZSq9i5rRKp8kmtlwkC032g+w3uuNJ
ne0m/TSHLwAsCr0DzUXFzUX/WZT/q0TKEbho4LUFU0M3zz3kMclX7rT5jWSG3rEOSLPm/x0IG9E6
4f3GjY0S2CQPvZKXMNG7zWIKwrU7a/L3CIEMG7B/ugK096Idby7FB1v5hkAQLya3KCo+Q3PncHgg
dvjiUORbGPjqa0Ulzr5ycVVopQ4W/ZQ5VzYx5dDC9+vLzuQicj2enChrHNmlWp9xOurTAfHuiYrI
pYhMnFFuH9I/TGUXVobEk0TWOccx7rQUZ+FVacHvReU4T2kg5H4A/raZbGrFNLeK/ERuGWM+Mr7a
JiLgdzoEMoomc+0yC2Xs4VUoJNKljCjhoNZfISPcXYxaOVK3KWbNDx9lbDAaFHzMPddw8QQRjDfX
mE0oJAhCDHzJE1D+FMkQhRgAVVL+O5kU7LcYnV+DdTDAeUpJme3ht8lVBDLZHNjf71K3/VyWS2mf
6FjrM4W+brbSqLK58PKxugRf74sPnzOpbkDOizHxxOGzGGXFQ/OgpFVsQqiDKB1EtrZh/C6V0FII
C/7MntoGIFENJBueBT4a2w+kz9ijYm3JJiUL6AgILSx5v5fGOUtW9VT7QoV99MLMi1B95kXOJXSM
dj7fRJ6ejWmFnLeI94YgNQx+rePOkC5CJEoehe7YZKGDS1HqJn+OzEV1U+AN2jlDtCfVn5nwPXrq
JdeEUeOnIy1SPXOLSeACehfLUdvruZTQEjd0BYYjq0nUH154BtxmZ7CdBubiDCj6bu2Gl23cIOo5
MyC1jaE6yi6eLjRa48rpnJl2RqHfc6AQ/zQteHQ/kjm0v8wVlvpICApI1fChhLszel4vhNeRBNPZ
KkSbDSCJZ2GSRun3RVFGn7yaxXLRJbGiUupkAG2kFbAqy4dq3jHC25qiYZNxsdtPL7/PlmKrgQlT
duVtc7k/ppbHJEzd4S7/D2mBoBTpLIusItaOPUSvmk6ZbEi0NaQ7OOOTiym+s/rcaU5peJlGdVVt
3VUebKD8rP8R8XbXPxsxXWq2eo+V1L1WJUVTIN1bRBXQzZ8Dc35iYGM+0srkvif1qvf4dXpdVKPp
1+ix5sVjMB3w3AJb5nqyGxJ5glU/ixW7FJ+XexNWxtDGmftJFhpcC14CtCnmjm06GhAsPqjDgdGH
Yv6NNrvZv+ZNmikQL7d4khkzj/ZibvuXLH5c8MsUrPE1iPRlKUVtLdFK53vyJcBiqcCRpytOMaFE
+n2IoqgrejvFi6yLVbAbbdzDTk0mCNOlDad0vbfEF3APJInYuQtzzr09oTmV+ILuLA0V0LOdCrx6
8ziBXp2Za7kA00utzOP5KCbqmsLd8vrplXCifH6oJTL9f/jXFbZedRdpty4loex8fWwYOxfewMEl
ai4RH9eu/2iA00/tfw3B7l+4pLv0nk40lgkqLtOocxBnKmWSQ/twu0kCsj6/L6QK7hngMq3csYwa
J/zQkrJSkCZqFBLUZDj3k+fyRJbEI6vXJz6p91iIjWAw4co3PymPQ1bb3+qBeA4OFcNbw1t3abvp
v/hDU9zChlOFAHTWI1WXl1H9ZVapxgqkECrVlrH9TE01s8yo177o9NvYdnp0+y2Q5r5wnaykPsTr
ZgjMjmoYB4TAQ26GJ33onkFVZeVzeQriy5w9esZc7EmAH7wPgYYT3GRWgBcHDJBj4/ouq6WL6ft1
Qo3S8IMcxUCDdUcakryQalTWL2zkJS0kTBIaDOpx8mtdsOcytjtpPN1dNbJO978NG5yxY6CZj2eu
/vzLs9M8ZhLV8ABhwQ9uLGaPX0a1Uj8YVZ9LFcu8UZdjtKcVrN5z/qjS1588TNuH/4fi3tujexRR
E81eyF3r0EanmXXRMT8ZQhn/tUtWedamalXuavhre6eS1QuUAAwUqJ14PvVWPjqUC+SWJPWbJm+Z
2Sxlm0yqXpBKEb9vYLbHJzMHYw5WCHfq/smsqSZhw5dECypwpIKKKDDU7PYjMrqiXuF+QIclxg7b
g2HYI1QTQGKm+oqjLG0KhkCQSwrjIIap/YkL+lTLyHca5l5cspT6oPCWvsgenmhQv6mQer4yovXH
Mlp+b63g3uqkTa3SG0QjvZ+OwIBdsgAXsF0CM8tn1ihTi4Q8wrcca3wE2vohYuXWg92b0Wzv3It/
zx0AAj5QUC0Tjuh6CTk14+TH3Wh1KGAcrwie0n5RrqB33Dpilz4RTb1CCBbC+NXsSsPCOR0dY5RG
t40wh3aH5QntcDvdIxdq6NpecbS+Cwg0yfz5Tt5ZO5WGPAXRkJ7J2Z0isa44H739BZqXD5B7Zviz
VrQmtmiU7L7ta7RGuVuA/1b+GmXlemXUy4futCZoZmyQXdhM7IdPKnut4MQqbGlYmgg2QtA1UJRv
ZGuKwX396hN0lXUeHo+++2/fG93CvbFwqMwAwtQDXDGjGUF55GQH9Ju2qXWdEsvVDVzJUZ32uQg3
ig/ihashTTwp/6umjfEKOq4V0CdR3GmrwOQGuhHAWlK5ZbFabPfEd5R96iXTv7QFCYQu5yTQyTQM
yTBtLXPWruInR6TAjWMPZJ2lon7S7s2UKDal0nsTfbEV4Ad08OKYz9rpB5P2HJ3BsWkXSv2EfaYf
6POiF1OiIArw8E/GlGVxtpCLKJuzZ08IW3v5cWegiAuvUK1HY0mJ88HQ+Fmr9ylBiTXaDCa+z2cY
QR4FrroKSV8kV59iF3RN79g8zUn64KajXtYak+W5qrG4QhDfuSYd4YJfJChOByT4G+6vTvl9Q0d4
ktvMogCFNLxcAeGED+w/eMQaCZIzUwLoi6deD2IjZU4UiCG6BIiSUQKjPbwWAgiepOo/CBypgL1b
l2nYFokGGLzIyS29ev+O1QVxBX+kVtdDPrLXAg2DVxgEF2/atMejToMuXzPBoestjjVdOuOk1Akm
Jbdk/m72bPufjmBRvPyK9MEvBnPnEFZTdCaqrsT4+FiyrqOGyXewU9lG+luPZEv2At9QIxN+hnyW
Q7NL8CJPSXEMOtxCGnZ0r34wSy1PaJM1an+uf8S175aHs7oqRyjkGxsxOGcVlqsX65vMhcDq0urz
gRvF9zacKGmrcx3rDojj5nZ0oY7LFlIfYRXtpla0n3fIRugAHKRLdd6wvsGJLvjX3oe+Smgh0RXT
PtqAAHGCs4ud8lLVjhy5REZYURadm2T9CwgbE/svZ+PzMJ5psEiIN/5L5kqeFQKyipW+mkwr5pR1
3Y/CurfM2hVmdHOyWOaD3g+AJKiq+8Apms2lhqFVJzXtH5CDRyoXcjGoQ+AaWMQNwHbB2cNaS2CI
ButP3gtJWcK2hDxhMj6hRYnNL/qgFv4tkL749PW2lFSdPuYXfkoamacC6Ibvk6Vqc9vx2/HklsM6
hySnKRcPai6RtXi5Oy/rLfWTVivDHRR7/YFCpjqRydfycyBVBhQ9sn9NyyKQPOrJ+AviPud53asc
IlZjoi/6onQc1GIhAdVzCtpAjgqqClZoA09qjZ+FF+KWYRpVMo0VOM1tV303tpUPdqS+XfA0cYEO
E2ICnguvYA8k9JxOEchXxYbMEgmaE1dREejo69QuALkVWisGT8mD2Zo8LIcVoWeJPonx5ZaOmzfa
+j6QzglCbb4u/fRXFIeleQoWZ7cBl9xZfrJMwNo4FkA/J5cMg5Bqfknu0ivwZqLRsG9fHjiVfFyB
Z5yedvfDzK3lTcReo/sPCW8QztEEoYEDbFTCyIKIRAt6Vjd0fvakILDqQhnoglNmJqQ6XaquG4A0
BOXXHkO+4SUAtmqXn8PQtL6IFfU54l36wDZ+c3Xu2RBfyQedmYeUbjrSD5v1DENzPxMpP/FV8JLz
cWja/QGIhmhGEwjV3CTlv1PSFBjSGzxzA8zJT4cekCt5mWIZLxltDfB0VBZBzTbmCH4OXg6fBMb/
HJJHpEITWUogL7SfZ2YlVBiSvzNYxzJjtLhniVXJKA+adj6OnzBVflfnqCEuk5vtMeMvxoZ3GEdA
91PfzhStNBvlAhRFEqbg5NyE8N2U6fR3pvz2cl0kvL8nnRtil5t2Aukrp7gI/h66rHEVdkLf/Bmg
x3pdFDI2Y+o0Phno3iP74v6Qa++Rw+ArAvaGGf9zUDvC/kErTHxZ+VqXKFmusH9NiOjXOxacol6V
345u1bViHC0aPFyi2uyCaGgtfXvDsQZeiznP2d3vJqpB7gBZnrdL5c5O4BPOpGRBRReclx3CoBSh
CNZcq7a8gvtdzfHRBd+syZWqOQKL++eb1eKZPkc3HN/E3/T+DMyEBZdQsXXUkSqcGF7wwxU+F5Jp
OsREfBIJocygyqVo2CdIeb9l3mqaGhL1vUdBf5jclC3XDCZK280YU6fHQpI/REMVyIinRIhPlBhZ
9LFWf/lkYNT0dTIPX5Ekwyfc+GATFGx47bacEIrvhBtFJn01ESyNoh6qh3Mjs25zM/tfU/ctWLwT
eMqZstYaH+RaDETQi0zHtwA8KacOWLNi2N4YHz8QfTr8hROVQ1zM1tDF2dzoVwWwz/RxTEKAfHQS
wCCRfih+52FMNR4g74QXOngI2S2z4LMXnnnoBJQj0+N1DiCPBdOO0i0R6r/BLFpm+tmI92j4LZV/
J6LhNt3iS3QEk/5SSGbYe/NRTu/wFbSyQtGUXyDQGKPAPJBiBMl6rzkFTf79Ii/QUuT2MqTE28In
J8NSSrQqk7r6xdp3D9Id9aRqOr0BXomUEEbV+TB5jugu5jH3bbRFY9jnelDpb+Sr0fxTs2uJVWCJ
ZkqL4KDwlT6pFiW8V/Zn0O9+2zxIsWlbJo89RT5JZYTfPBS3MHqBrEd+o0ZJENF4DjaQuvdPQzD1
4w+3dfKelmX58LeVWPesq3lmT0vFbS3K91rT+CjZ5eb9KdcEnyyS2MMTROxaH4A/JbFiDgn8r2Av
q4fnmOz5puYDeNGa06BNSrp6munxaVKWBvnTUo2CTXM+c5Qi4UD7xZlIiDi/FT4nu4RaEDLTHV+y
ene2H4gr6RCY6f9wC7pVebNhfrEBorvC84Srxfivn8luYWJRVQ+YH/RmKbXuXLMFxM4bTpiKvSN5
O6b8Bcq0RfEFcxIdSO9u45KwPHSnmAfJ9LdDTUe/IDtbsLFGzoS0MiGoZaI3UNtd8Yl8H0A8Gd0A
RnifAPL/UKonWzzeVByaTqHCh+y8tLhYKyNENpLKsRU7cum1gbPwwkAcalJ9RZMAcyW71JVbDOuN
gWg5DDHJCV+F/1fKiy6Y9+v/0UyxQwrUz+sSfF4dWmalaSq92qBK4sH2p7iBAvSlNTGGUuJJtUaK
9Uutjmt2TR8ocxQO6vNkHYExUYeIecGChIBPm349jWQIgCh4tHuTnKI/3tq482af6bOw5w4MksET
9B08O0VjRkjNG8TiRZmeaYC9tmONdrMDGVDKp9eGm60mJtwscqXGJ46AqS5za/pahPgJXiJR6BaM
lXIYvny5qu5lqAOafhpKfPuAYtrlGokAsUn5xjZEq3euWk5FjHkpslByVHsstHf5ge87w1nJgw6v
/iNck6zq2cuQFnnSW7vUx4ryXFHyd80NzDahAv9yd+IaX5/UFjzizU1HsvIsQ4pbROkWCCzvbG88
aGteQ8gWIbM1kXkcgJntMcNFiYX8NPbdYVYf9wSx0RZhkXFPM77/tReMnLuJgBMjkKjyHkHI6idl
n0rQlqeZlowzTpDnAeUAM9bKWWb9IGUyarvfuhf80UGEzAlTY92XmtYj7lGFR1+hcg0pNRNkvNMS
8c0ad1IjaxCxz0bI1NNcn/hRik5O/U7FPKHLCwTpFr1DFCcj7CO8x362Ny2Sd3iaKNMacZrtYH4L
NQ22lcTzYoDmA9OPrdgFBuxbkXTKG7I6z08AixnmBn9JOqSuIj6gtcEfSwpFlp12KyNAI6r5rmG7
LdYatVSVtVQN0sWDPU6akE8abvsGaxFnIap/PfnHMh3AxwAG7TUEp8X+Ie8o1K6WDKhU/p8kA9Qc
aAyUDEyoxSGkQm1U4CdO+ig2ybmnt8oW7LXzFO1bcSQ1aZyazC9nl91pYsB60WjMol/PANKWI//a
gP0CUkKME6VxqWfk6mI2rFjS0IbaqS7XhisVBiN4NHENsBHoWojNfRptEhl+059O+7hsSLOuCJM4
01pk18QJY3fFNMibPvCVa5ipDds/1VZExd3ERvl31m4K30Pjmj/YYWK8PYm640TLKcI4qbSd88I/
t/IKbqg9W9IuSMwbRlrOlGLT6XQsGaEbculrYV0TxXE1JhRnoy+cX+829ro7GXCAoho4gFIIzIBX
dWSgo8LTzTnDdr0S5QlMfAIW3qtKZ2PArAaGX51ASptbjaKKA8XGkmyVlbrEm72XKyH04UyFavOf
KSJ0nhmn8WKQlySYS/7Do5cV+/TXXCT00Kxott9f64zVHPVAk2cmxr4bK+UcHqk7akj+Uelf4IOP
Wwg3xhrctFosQlzE6/DASbtTroyKZjoukzZZtiVqhBQyRQpp2pl62aXHXM3LtkmY9lCC3qHuU9Lg
2oP3NgevF3SwYIskBmxCJo+CWEYpQLDCfgBCc+cWiJ/iSvcyKwLUIfYQveelcwt9ZkyzDTIcG1Sz
q37gOmEGI3KandKaR5QpEHbcqWYuiQLN9Lw8vhB/lfAEsF20IjeNU8MTsU/EJN42wnYdmJqTzBqk
aQXZEqmAnc10YAMrHvNY25PY9VQf9yhK0TOD76yDTA37qfPK4aeJe8pAEGntId3+7QvEnG+9rPVJ
nGOdLaRzRguCcvaJgvdDtfpNq4TO8wZI2igccKB8r0EAuElONh34JoWyj3FZS6QKDPXLrLZr/yT0
Oe/5Zzjh2biA6jOdNKGRMy3exz0O8uSFkGdX4sGTg7gl0TgdcGWbClc++pee2JV08C1/k3Ddw8X2
EfDYPNPmQeNktLE247ProScGgQOALmG0+oNu4XjTluSdMHezyrCqvKwuiWwQQyftW+Gq4gowe8aF
vNYQYH/0C/Iu/mpAi+IBp4ZUg7cVlkdkWGQ2KrGDrJQK0ssQrV+h8Y3mlznzvmh03Wuu4Jz6ohZL
vFxE1L5te3uh/RAR8UtcRrDrS7zMb/lQ1qiOV/Vd2QrcyO0Qod3xoTPkP4t84KanqxiGfGxadqiL
30NEBZISaxKP3Ndo6SLVDMXXHdQkQNWktnTvqJk8X5uEG2ibpWmseg8gXu4/4gJk+IUvPBrFNhJT
JFqxSxKp950UohA/Cn6658DG4p8NqRut2WFRJLXIT4EO219iPxKXDfwccUj7WeNCnU5tEka1ubLo
3ltLUCCXcczJt804WaGma4HqhecB574pv1cf9Bt/+gmHRJB2SDI9WAZWkO07Og2KE692dNTjIviQ
fqa2B+j/vsHey58nk0f+N5t2A10vZZTn/IdR1YEtbveHMoISeZT7xylYp8qP9d36Jgk1Y36nv2R3
eHKRFlUwL2wuiJbAaYkUZzT6h1p1xcX6Y2iw7J14N1PKA5gF8dSJATTsvZCPk7dVgqlo/0O7chyN
tiIr6qSb45V5SBomSxnFoqQCOANEekVcRjeUpz31fLcP2m+sbHA9aw0w0BG2OQDmMMpGE1hv1vnc
YIWjOmBCa1GgU0UIZ36D5aY2ofYo0mrHG7NbpTQvCy0DPIqsHStkFuAQFGLGNl1V3i2I9iPX22+z
Dhm3pcaLryRGWCKbKGGhb8+QY+qapCrkZB/24WZXCQzj37RUgI2etocvGDlO+lzbqDuGo2aqYw3G
rxX8Q6qjJB7wP2ORwC23k5CWj7bXgpePBFqD9SwwcnZl4/ZeHxXNIO54ZKQYPArzGRvESC6rWcrg
m1TAEhjLWmDtRVsfF83fRMUEczcO4NmzEsURF+9iilvH4pHtY6ZgyY+gBepDlRmyAmfWeYX1HOdY
uqo002oK6tGF7X8phVByobVaEnLCrLsB+QhxAYIqti9mV39At/kd0thaH7Nc8rOwsM/GH3FHM6oS
X2e1+T/gsadQeltw2t8bfgwr+nmxp1LBBDjEg6ztCT/B2rG3gEeun0JaFh3BnREgELUg9yhZc7bi
EBm2mnlWguLkXD/LKDpZKlFeSoGWj80TebXbQuPAeFXWiflEbr+KsaQocaFWPVwx2s5XLe7mSfg6
lBlgiGoeACDvdnAFLzJk4VB5bCLhWnu9DsUoKZy6mMOjQCdncnnUlVsPMHaH6+hUa1yVqX+9RbCU
NzRKW9v7vmPznxld2ndlFGdwlGu0ELqesVfA0s4Cc85W2Rd4w6m9qcmjVSu6WV8NKQPiBXK/8tpo
lCsubMfea8DcepC3RiZzeBoYmrEhLruTZOtR8schbEQXUhDjd8A8nIGdySN/8qOFeMwU5nkB9GCV
0YxSdOGTQfr8afxiM3EMSMtUTl9D8pC48oBQno2GrCL4q44iNQEKVYwRpDiBE8CTUCOpwzSYttzj
gtGTLMSz990hk997Afkne7RYCYeSZz1J9gBTO+fxz7xtmVcdeaLOtUBnf7o/drsd1lKfqUnWKi0m
/cORZOSSs2/76Qtm4EjaDJeWB5p3qLX/P0Jg1Lw64wkWtpArQFv/ct8eGm0jiTQYssOPr6CLrVEa
OsJ9Aspy7/mlFfyRZCVSI2oLZH/ByoQpDVDke81TxEuRlE0HLnGuBmVOMLLI84osi9iuXwQ2Svta
rsEKcil6TTzyHkEP9rxYL3SyB7iN7dYuLZHfNVQJMrNrxulhtwHfPT4YWIfyvoOxdhbcKGSvMCBp
xygKTqyZcdPtVPc+o3bvKSLeTa2IhdwG3oppWK2URlynfg7153/nskobAKFQxojpJgEBj9lPiSvi
HJlgHsbVBJi1XGiMGcFDx5lYJ0VPJM7tygeNxHran6CvysqBrY+PYxbw6Md/Omrtki/dvaq2pHsD
MKjOmOC2q+v/skvlo26o36QmPP40IfPzL3ALvDzKVsQn+pSyppFLVlKCDSouYvqf/iiP5prDaUCV
zZpmAjdZXREg6amdIqTzY5CKuDkmY92bRJT82W9gtwNk8HZgxN+fRRu2gxxzZPxrgMSCZyMXy5dM
9p2GHea3RT+auID0yiQIwBaTqWOsL7p++/k8G55vPh7m+19CZjX+H7oLyRM0++Bt39KDHZdRW9tE
JDd0mdf/JiD0qFDR5rvS58SMEXLKSsKtt70lYGpwkE636Y1L+v5ONDU6tkny5Vt6kicV2d2Rdd2l
0RRoccL0F7WCtpL2+UvQEq0z8m4MlxAM+yBmk77V5TIns++uOCd76wHwUozedBqME7DeP7QwL7oP
JXMyRvoV8UBDdVdpbr3Si1vOVCSXnnjbXepyuPYWXsHVaEJIqpC2nHkFF0CYQJj67svTlEsNK2aI
KBfoU8uBU/wfkhjwsW/BxqAQbcmG6HwHAki4UMVCZKKYyZYwu8HZ5BUaHFzqqbErjOOR2hiheg/g
gULph+TiGK2Pcbbz2ci9BZ1X74nH4AfHfBtvoZryxP4v4JmTFWrPOTGfaDhvcUklU5ldhvtXqyyO
XbSO+Q4YkOzdQffsEaRAqWMfoZ4Q2cBppL7bU6LGz4HrBo15zuLxaoyXCu5/Kwdz9CVrOs6B9Ciw
3bHxjjTul2R1XPts8JmcIxoFLByMHOAyaLkb0D8nCBoOVxi6M3Ht+Ug+DmyrBCdCgGMsA4sGHXgr
wRjFRbOtBevmgCk7qgFG1ie8Go/RKBd6L5Z6Jn7n3etQURyloOV5ShUSmsLAAIsahmMEPJmQSCX2
i0Li3docfBqd5TwaBidsvykdGU+oQW1lHjJjUAj0viucK+gUnr+/sLm2aCGLPNoV5mqISTuvs3Xo
LbD+3FJx8r1QgK72sfsuMb2P6BRW1IOdX64UHfe9LyXCuMQ19NuEPKOEob2Czhq6KftJxuJ6iL6Q
tof7yy40DvPoQVInTmji8qqFK5QZ5sK8gsXTLkC+q9AEqaaFTb9nhLZYg2+ikIdY96VzI3sht934
tb047gjYlUzqWuEnRs49gf2t3DRkl69m/Gi2/aUIAZPIKdnRNQAVuaghyEaQA6ZlAvhhjyjjOY5W
4gd0lpvwHbNm35O5c0HxGhuW30MphHy38i+f9tMpNnuvWq2OOn23lLNlQNKlXSdZBuMXWEiXY42X
1zKd4wjadEgvrEmgrzCJTmib1JnGD1B4/KOT12lv1TNHSVBXx/curXZuiMM44WxqiMSXzG0hHAwI
YrdfRQDQE+brgg8T+j7sax2PNLjrRYHyrcQQdLsj5I7Bx+ixpR5zXC+BoZ8159ud3dADocN39ZVg
Fp8udq6MqxjCgoAtKHbNvrmvM2Nih8KncmzaBnfzzq5Y6mtKh2q+H6bCINEfetKRMhzHaI5XnCTS
9/E8dxazgGjsF1bFfeE2KA6AZCGj8q72wvfjAdBiBRKmUiG1XMiSnLbtS2goRMxV0SWuOgRcvGU4
9hVebXDOg+aq0c23uklYtT1pdkgsuRagJf0i2G3RKUn2ly/a3IRUuFuXmpX/wNDB537kfHlHvjwa
CZ2fCdlcfVwzAAOqZ5Zv8OmsikBgEsDS/eHDJ9aM+hZUIIZLaSqiQOauijSyKPJbGDQCSDi5AiOd
tbwI+RGqny6hxmNnsaYurshgKz+JjyskT43yxYZFwQl3+YmTmJ5Lm8dwtvR5EA0Tm11hwpNnAt8X
VvHLPnphqNTA+yOUZenEHZMNkHIaRHELqJVA+Y73GoNpJm+kwYPxMdcBbApMMx9chrI/oyvrxsiT
ZhzSsYS265mwk02vVgnqQlrXPvAK+KbYtAHwjUFi7kQan1+EzGL3lBvZMG0ZnMEJ0QIK6LByWtSH
YuZqhtVxkHZ362v2JQdNWj0lwO/GN6zBFsbkiul7cvGnxIB05mVHpMCpBlcN7m4/0F+SJ5Z0579g
IfU267rS/IMX2hplEIT7efxe5AAkL43c2er2eR5VxcKzUzOZy3cgc1VYF+mBP6UEu+V4Hiy0JJdF
Bqny2gerjyUM6WV4k/TkF5swLe3RCE3MJp3in+yAGNvKTDTS1GBHROf1BXl1gY0TLVe2RnfsGek3
rPaiTCSNLWuGU9J1EHGbnfAzr+dgqqlSy1uzET4uMqtOlMofvqtiI1e3khbPyAZCWNAChJK2grOC
e5Ih43h5IX8qnANI+cwvDRMXDfPDBMiH52v6iAVcw8yZgXp8dX+0cb8zP4GZMFESW+8XoMr39Ky6
J4oe/kItvl2Oipjhw72sou45OS2hxcDl2M2PymnOU8uR2YsKYtHg3vB0N+mJJFPuxpbXH5KgwSwD
4ptlWZAf9Qnh3rWimR1TMvMaqUla5czEAN37xLyppo/9VXoSBpwreXHdnk6iC+3aAtsKj0g0p8aJ
yfq6E57Ikod/ibRMc0fEeJXB53c3B4xAgv84ZDe0Qtx5v2SNYZINrCO7XbdYveiC/tZsRotrGQij
DTuBhwGVoY8BjSbGBjm76T3MdiTXekph//rOWHy9Iwph0yuYS9lWjRErrkP7P2afqimr67M+7rEb
Eq9eGwRRkHB/enZla3J+/B7yZ0m2FC63sIeTKnYLRW7ZWVgUG50W9amibLnaxfpgcrYZSpkyEMbq
xnRVtOxllOI5LJnLVlOMAatBC/7TP0bK6L8HRqPaGVPRjb6Uuyd2WQ61uxnUSXZkMqh4z+4w+yjD
5hJ0w6iJx5OcHsgfNAxrlPZir1+Vzj4ISlNSGc9prN39EH8tw9HPN3nvnw1jnTQ7qqTpI63FtsgV
jc7fMIbUbHj0sGkrCzJOP5w+UXmupraXTSMr3DEOcpH6EaL20gLMG8C+FlQBKQJMF1kuCjUNjt8r
SuSJGt8MlpM6n1n/+SKMgdg/ihtw/OAOEIEgfFwSKpAsXySekiDWuc798o95KfndspnjgSBg/nzG
5m+W3j0Hku+KOwX6XuG1UbkPVaEuWuF9PJ8YpXblnXtqYwM3/aTKBdQqus9pEXZwtVPpCI1W/JXL
iV/XfbqrcGmN9bkdSzlEO6VOeexXEq822q76IdBfQiivmh6qgKLbFRT8KJ4kVeX5D+wqjLvioE3k
2V2D5nIeNZpwIdMji4aOcteqrn8QP2qW2sCuuoPfZ65MlOivU7MOxlhTrByDerr5M+35HrpCkmQ6
+7k83J+o1EbHgd4cODq3PAthaand9Cnc7KC6bOkjSvcb/LLIdYVsGKzeMvHjvqjbOl5C1ewFZiZ1
7irEvDaFWJ56rvslDcmFN7USocpscxxbIYkghMF/2f6KMf6//LedyD0rl0KAMItYUeXkpAtvbkCN
B93C4OZEQQhB8S/4nWE7rUaB0iD0P5Aq4NruH06u80FmzdZ2CXwG5j2fhc+ZCrcBg7XFsaWhh2I6
Y1QBR+gz2i6NmzwBh7wEcsEbi+q8N6e3sd7D/1PyW2HfRA2F8cZoSUgN9ACBnFpclxSw0aH3C4DG
yZgsGmgOx2NQbz/hrWhAFmugrFVX+wi7elDj3AQz9I0pFk+SeS+svmlknwUN92PwQq9UqZ7aTGr6
hCIOUsDhDvcKjal2Pzed6+VooAe7aGFPzT9dRo/IPCQk13Sbd0SbATOynkMEe1sPN6GSUDAvJzlr
EUn7Sgals9tj/BZNfUP1nKEgGQLWaLwJSEAG6RZuCoXgrK4jlyUGOA87hEpNR7GO7DwXLyWZBDua
u4O7ghZZb4TJDmEexWfzZIsnPXGOBEVj2icSswE7kqBp+ie8rxF+FPQM0+Od4YY+1k0ktZYOHEX+
Fqw/TH7KVQwarDpvp+zqQd7/v+Qplw0RrGYYQxjY7Iofu0ocK3BEN5yRgYArpcG6eH2dfrtyX4I9
icK41Kt2H74dHcuaEtenrkWFMvcq586Zu8iItpU62VhhzqnHsBxgzSUqyEzp/z4c0tOW2ALvqPLR
zd7bIQr95TV3Qwh7N0xR4cgTl2oZ3ZccdAforXvxRwowEiTfBJvHDGnXP4IkoEddcf4gZOhICUaN
ZjboabVlT6vRphVYzNHEKj4vqqIYL0jcr2Eqwt2Fg/D0qFy9a2B5zuFdasl9daNtzzVh5pPXxGxa
14Zq+Y2vS/iep5knvyQpto6/RySX4LFq3F8w24vl8BXi6ok3WEexSbYc9Zp6sX5bJeRl+8FbMe2J
sGkcC6WTWA5K9PQj9fY+Io5GyVvPW944CcABM0obV0QubhmXnI+g0tfXTWhtqQrwsE1g2MZcr68+
UQcbDMgYuLpyqgKQQ/10cybMsqaJkka5Puxsoqj+dokAm+2dfOVRlhJM7KproUjY4jaw7uoWfBrC
Dc+PrKs4p1RhF8BYMKfljlmARBuoVBrT9emNpLnAeLe6EiR+jFhWVlu7GTY75IS80C94c/zP+ku6
kUUdvKz0zCq+nVGeQjh/qGaB9YdbHSk1S8r7keM7c2uXH+bOqf0GcjJ5FtjYDjKcny2rtRp+/dMB
VMMgQqSnFUtsSSMqfR7wzjyWaHWvPBsWxPKA6W1YNK0jcDK6wkbr4Uv2J8eKUww+0awM5vsTTH4C
h4/dHKJP67cKZ6gN9m5whEJXtMy2M30CVWwDW4AEk4t9qWvmWSXAKCrg9gLyze2M7PcMBTEG9QUc
gSs6ezAoBr0Yx2FUuROOBvyEuvigQk/RsL9Ky7RO/v0AyCfKxg4BJo3TKIxD0l4W+/1XN1e7VQUD
65NVqyYuBcV0e0g1ssg4wRQDtOR99es/V7sy55F7CYkcW1A5bWtfViw13PRpRxcawRIWRAPMqyVy
Q1q3Ru31/rxE4ECv6CcXRQu8Q3WafWka1HK0Ym7XoNZFC98Ibf9fb54ixYAALhGj10p/Hs7ewFk8
MVcvGlr72XK1+BF2vbPYM1YE8vg2kNzPGUqMImb5JrwiNz8YSOIvcGV+CI/NKejViYw821eh6RpP
+nahl5uLROaL6O4/KbG6bqUfTEEXDG88gmfhUz/Io3HpR5HHamFmG6DF7dt8EycWbSjbf1Bu4OCg
U7UCl9xRk2lRgRrR4ykOIi9j7s1IgZK07hok5N/sMBRhplEaMy0wQJHhGX6wS8aLaUoKYP8BRWvi
orVhdDJd+8Tg8TcaOD4YL1VjhJPEkn2eQZAIgaZIm1ITe9LKulrW3SQjeZ5VjAtD524XZaIsLOW1
K+E0PWi2RQqQUjn2fE+fhM6hVoXpRBCtV7TisMejX+1FSHscBOAcTy6GJ5OznCTCiq0EuEf1yj2d
cXHQuklmzk5ytx70aQyv0IlpWqFx/z+puq+32s/ZCTCtoMmkr/3O8b3CStka9A9cZCkkVUfvTh0s
pQsvPFKjJuN2Ow3IBkPrTuBMYIsjEkv2o2p0alt5dmt+U/72Fr+kgBfPVD3ygCAmn2nS8ecMcYHw
5r9TBxuE7GV6kCZ26BpYco0+i2Rw99BNzSNKgQmTsF/Bt2TfqZBz3EhLyPppC0yNmj3cL/vd7QIB
r+eBbEXZLhuPhqTXrXX3DuWAVqxcmHCrPeL2SO7oMDULXEJ3wGermmemgVVVXSIh0+XjmI/J5HUr
GzevNnvFUGmPWMB/fEkCeN5FtO1sWvJtzKh7zHyU/D7Mk2D43kIQOk65kNN1+hV/JbGa1sxQq7jP
CBDAZpMbtt4nItvNcqgONZjADYfRyMe/GpWH6LkFoFIOUDHLYFMsBtJnT8Ks3J2xKu4RqLaKiXsF
qwbY0aGccxyx4/TI2qzMwme20TXSFoE37fYJEG82qzdggJmdtgyFmc1xydz0MaEjFJImyQ3m/53J
9j00SWYENvPpl5QhY+KeFjFKmIX08vKjdKkicYlihrmH9Sp5zePU2NwgBdbQWwh6CZUVjvPQbvo5
sdWnA4+WftZIDE22p13UNll2aCRaRbKLq1Dl9PZWIg8hyVeX8tZmSAvMzjtJasGg8P2trwPQkIbU
ktcNXjdXwcqpYQBCFWZhOPCSGciKNy4D/sVvK+dZoYsA5nL8I5wCp4Kt4bFG2ahthgumRafbZtzQ
8fc6DZIGiz/dLvXF3JEbJJtzpAyvSQkOY7bA6Cvgo37buRdeXz28ZAHtibKY1xfOyTI93L4PVLab
yjeiIb+1mTzTUP6BNF2gyz/BPhUjRWRNvruuqkZABPsWEZ8Bz2T2e4qGQDNoWAiPAKk04K4vkCQV
u+OM3Zu9rrL+UwJTsNkoh5D8dqegZyedVrtWMIJkQD8c7RiPQGLj2dHZ7ByY1SMUuIYVBBQ0KNtS
zMhFUf/bSKtcP35ltaXI6WOqYwOklgrmcEjNceKfHXwE/z/jmd6H5G+qN1Kxsyhvl7XgW+Mj4HDN
9mFkkxASseKKfmgfl5xjtDIQsGlN78KTpv28DwwB2oDiWZeZ6obU2abtYB29nsLrliaPgsxbBajj
nDvJil3oZqVvA/tuwUcE0Ufn5IMzv21p2PSExtFKXUQGOJtLcIdNUuH7YE2hJeRCAdKozjcEjAYs
vkGwrrtQFA2FSXXlz3I4KBQ3UXNTK4hu6tCSqapaONG3zWSRS8Y3XpVuorUTqMuxI/LAXY9mVLLE
vzc352v71kU1fE+oPcj5DKdykseInczcJanhPvoeyzrdsn2BDN3PKjAwA7ZD7GAWQ72HMcMOMrzj
Y63tZP8bnbkajbUXvEzmdGhnv8p4aN0w2pnExmSY8sT5OoJnNh6kwxGDMTClnkOoLt8Ttuec3H22
V9tbud7JCNyL/Wywlbwyq7bTBrWLAhvALZE2UQNrFsLaeJzsnVnZ6Hn+/dcJS9gbqcq/6BJUi57T
l/ma/4RZtT73RxhCUjaXKgseTF+4d0BqqSrR2LdPIT/7DwkxlZCYHDUwozTIM9LnmTruyn4fNYGS
S8UCg16QaID8/0tk+t5omI0EX+FAzeDJmeJcMWc/2A5pvIlAGKZJoq1Loc549BXaUFLrjy3A+7aJ
u5ViBuxgeg4VsdI7hjscOKClCNQo3aM6lQGq1m/ztVJ9Lx9Rm7qJxk2O8LV9SykSjpMj1EyJvqSD
6FM6/ufpToyfo3Ag4+In8shOvsAa4THs0yTfc4/mX8kp4Xfb9LqiSWukWVMBF6TC8THTHhBPAHk2
BBygF244huBjRFrMD/1Bk21H+zhTX44B9hnXPMabkTIpJemMN9clHeNmrYGB29Pho9CRrfZ0Hylp
F3R8oZxJRpuvylKmfNvp0RY27YfzXrc0uDbMVTJmOFCIocs2jaexWAlwC8zW9/YopSqK9x1H+HKi
WDBA+n+itgHrLdBNkX3RuX8itb9/A0IRNyAvIegK/03DuQ59CKpwtYsX9Lru6VM4Olb/41ohd9l6
pQTVfpAI84zC0cBeISvTqlz7RkO4sZVHDd1Cf7xqjfocJVfuOXMtZscEJreLiHm3rpRHFRzSRIWL
3nlSj8uiJq1hd/o8QLkmBlFMcGrB/8hp4y2Jra3DEKDdGo0vJscoxVPPabf+oYLTSvWqGdnBwFQf
hp3TsqLAsKifKS5DrjMEByeWRx1xRo02rN3lehicM/N+0UHF2N72BAENyIT2ANLRDZhSp5xbZMXz
sxubsRw0jj6AxhSzl5XsDQZkUomjkJP/LgIKv/05cNaqZo1M6BAU6LWEat8ZozG7ik6RATBx0oHZ
/zjpyqkr/Cr7tU48bj43gq40JVMEWRB4VDEt0cn1fg2/9V10e6dzKBgDaHFbBuSZcSJDq5R9C/Gl
LwlpotWr9VaSeCWYLQFFWz5GXCFQPPwcBwA7gpn4pJltIZ0qDiaYaesHgyi6iqsc63JzGixNf+m0
aFf9Gn3THyips1ZvmndwxCqFHLoVy5ZzRENa7zZkwBEoaVU9vwecBhwbV3/UZTqLXmyznqHH2J9A
Hz0Lkiq/9OGo29jMR6VG6RayucqapUHBUniTKUHkTGos3a0ACRLPusKd9+RXHxauaIfg14iKW4Sm
zgNjtMAv94s4cnVreIhIGKANxedOzuc8TfsxACau3mroNBsPXBwJHoJmW9n5sYK1uhvRD7g5trK0
1yHyzuWOaMa5/DfRIag6z1slieeH3xC/WtBdnbQGTZAkpk+ZKuCVqqCoWDbDDv2ZBp8qWhLJbmV/
ozM+sci/APLHh3bANhUG+F/dYTj3X4AsDX76YqhjEL5aLzAupYRdDI1zKr/wljqJOQk3MKRJ0Suf
5qjUjHZJdii4A6CJMEqfCCvx3DtZv4EUw15H6jOLTflyUGj6sCpX8VtqRgHFqvYveWw80HjvHVUg
FqElIfFcTyeW7a2TwqwGkC2w9qQU0izcA8zEuFIGqVKaULpjOJUgOS6I5gvebDZomEShVRuzguy8
zuXvMh5oJPWmxyTuIbU72BdAYL+XDxl2SQc+EHpTp88bxmTZyhuBgh1lfeasI08Igqa6o2UmWqkq
CU5htqNY5jPmnynluNrM9X+yGdPlgg+NYowqIayTWm8iuorCX+wLfj/Tf4F9kdbZlThNoh8iAwVN
eZiCGwVJyMnMk/rkUwoPB5ZukJhXoh/na7CUP6SGM4+1kBEmN5myi5Z0IHiCg55A0oEA3vxRxvI5
PJ8qiUDcRCRDvmcxDd3jAJ/zCaj0YZ0A6tSOGEoM6WP2LrkGhB6exi45mBvMM/g5SA75hbql9Kub
jEUNSKf1gkFnabeO1M8QSuhS69h2c115P5zvZP0uvYx0yqZCZlwxWwhUpwm/n2WgP9VhrnK0Fy4H
BkWp020XyU+GY7lRlB+hdanCKDGZ9K9ZIu/Fxg8f89Hb0Ao5P0/XADqzAbgjJd1Evbp8HafpdFil
vaPQ5/onHhuHZLLmoR0K/n9O2OF/1vLjpClZ8uMUQFlo5VabTrA5y98OingTF3UQcZqs4Wl7QkAj
GkObwRIl8FENkhgmAy/K5wVqzraLJLhW2oVu1YeyRwCXqTAkd3sRAtPnlbdHLACLD+SW5rQLG5JL
GIUydySUGZkS4KzEVVawdooX9kJLE2JxMlKig6KFCyGCUZf81w4/0OQLOPNAE80vamWNw1bk9XtX
vJWn0Qt0qd0ldaNbHr/Uj1NdOXZPZdIHiMfVM6j64c1B2y0ii06h8pG0S91O3HYkVc8LoJGEwJJF
AJXyKBPzFrGD3lEGzfTsOwsBnrfycNdH81Oe5ADNYzdbpthcIMf9xT3/1C/04LQMkojREck5Peym
aEbYvg+eReVNGZXU/1ebisCOl4ITUJj39LYhdVD7GVDIA/Vc/RGAE4sxZZD/RvTQvqe+SuhODrBj
Ct4Kd0gHyJfWAoGwgu/owg1kxGVouYmLxP+/2Qt+Mjd1pdXVgliRpT0cJCXpat9aMYZUE2oHgC/J
wkGCq+6Mm3pxjGj/ZTmzRe6gQVgGAk7yLwlBWQgHdZqhm6H7YPVsPAxbjqPbQNchc4BnD5oysfrS
kH0FkQnztqfJXhIJ0sZfQ/GsVFUHyd0V6rxqHNo836TuGr+VOfdprB0Dsds7rs4BXzHOCTAzmk2H
sWQGkD1hyRWxUaVia8SKJFXmLBuTrqgX/zdimZ+bIaC76T3I42vtoiuK+sm4gu+GKlg/2LONM/GV
xIF0DwyMn17PijK2XBlzObnDXsrsj1N8XeCwWHPCsmifbFuK382nZ4bFx064Ft6lu1Je4g3erqTV
NqQ+8ui+oa/hT2bwCyA27LgAywXoPQ7bnawCPsrv6CKVWLS8Q65jFe+KWDWVMOPdDkD+WQfZol89
IUNMsGjzVvPMyAvv92p6z8pvM7E6gK4BpI/WkyjqKGyC0AFTj2KmUMmB8GAuRgkfDBKCyVICepJF
TDpeXdiWdA2dt6shA87xIbkqmsD9PrgJrr7Noc76hG3qQzU7mavPlCRCcVw+74SXQiHwJjHQwtpz
X2GnexE/T6PjBBfS+y4tsvjjXedgQ0KjPFQ1RO4HmwI6pIbhQoThNcjne1sIVYNtOk/tztJUdeEY
upZkbCLXWis33qXM8a02uyg2dszubHXHGfGpoTBmhG4renDl4f/SSBQ5Zf6BNIlSVdYcmCpSZq3p
kbpkvcFUMkYv9utxvIrZC1uNC8SZxKVvW18w4YfoCL96QiVtiFNFLYqEyvxW8TBrG8pIpJ0/Cphb
XeKtNf7fjpfNwCzdSQFFNhAAGGN6SgPxt5TXpAIjQkMxGa0x/1VC6/rq46dc9oNxPXa4jICtdU45
AE+R8jcaTzRyGuCLZb10on6GNxvOpecp4s/UFo99n+uFh9gVRWbXcjt96+DNcN52LElydfZqWKlz
rj1rE0NIZBF0cUD1ih/7c1v6O5++7XNBoZKQEnEYKNGWbnvstiZsvppr95SUl+8RamRTxicdjjUd
KUtiNac97AmbrT9xdwfIEqBfa1/euF+A67eqwziB5wbLyj1Vtb0GhvWqK1cIVumc+v6BWRJKX5Uz
DgK48zu/VwvnQ/1MqzzmboWEMaOhRiN+OZFm8S0Wgeb/dS3yYSclN5DatzorXiFAa+0ChIPtHoru
EeMrbbDiH5bcibw6f4MelJhEHA+sBc1sPXrXiQiTdIjnN2HaG+NTPbQ9I8QTWb7PnQztFoSYqlmi
EcGgDjPNjO99MlHTMLZeRO6EwDgV/SvwmxR3DK4ssk9x7nZ6iMoIJQEIy544c1Ohuoe4S5Myd77m
yTQUP+FY8Ghg4f3AXtYFHK06gYxO3sUVXx2WRDEnb2w4fuZq/ybXm/Piqj2Zl0VPGYOHuxPj7391
1rsB+mLPd0/NMP2XbLsHR2Thmtbu/Xcibmz+XxDreEB6yv8UKp+yn1nHp/znbYSkqqngPkoiMywK
f4Hj/sZL/RfyhWZpMnoA/9ZhFslxS6v35YcdzZDgZ0t5ZFShl0hcscs+Ad2alG8hTZa5SKCqhXww
8xmsXryZMWUQ967nvKp1Rp/zoe+yoPPw6N0TRe/LxDS6ZQl+etJxYh5buYHPklHGnZzc+ea/oSSL
Bg3y+JNCW54di1t7+CS+YLsAzgURCdMux37Klk6uH/XAYkRTxvLPWz7xwKUS56NmPzRwgtZzdNqc
QPkiHEY9oSpoC0HdBTnKFkZYsS6b0crecGMjyRYCcjtCCRp/+oyo8/S+sR4slzswxhUYd/5wvOWb
jovSw7QzxpezLSxHCKKWo6sAnIPco8IgSu/CIn2tzkg/i+xVV5Y2xGmj1PbxFA09+z+9CHO03I4K
oWsJ/javiEiZ5KGSP/M/gQMsuUypdbYE23NESWk2sodATjcqBHBFJTWn4AXj14fMKnLaHWfnV2cR
2mWE2YQA6YSMxpGWGA3rlmQPiHeNOIFXrV+QaCSE0CV2eeOBHt3oMSZyO9tTHFpcux/fcdJUXPG6
YFiZKa5RsVIWGGc1o+k0KpTdxpTdQ6SNC6EUQUd1ahHsKL5MAf5+mU6Oeo4vXMf7kg5zXPwicQ1v
97YW7oZ5+yfzLS6llzVFbYgFoJ2oD9+UrWSHYTKvcnnbi7sC/8W2VYD8R1eZZMOlpT/NqAe0Ogwf
wc1WVqvO83h1hFBjXo/Sk1Pzmgfm/IXobkBRJNe2BbPrdX+3P8oEERBaNNTybGxuN35fVRbb8tvP
6pUUQQe/JlQhNRz2WJXA6ixAf9X0YZ5LgBk2oOFZjGGOn2atAR1wOLnX3dmkkVOt23yY8gmfHOJt
joQD8/9qYuN9TByP194mV6idLyE6TetR6J7wh5oZuIK9Enpb9lXF3JLkZNqwzMpFBwaTQqrYcZrO
xh/K0a7/ghoXm1QX9R1KsaWPk1MKK3BhNh+P5Liv3a4FiN7/Px42kcalJaOvmVdQXbWsei0YQ+KW
QA9/fdlRyQvHE1mXKi3U89vOjHcap+8SfItSbZ1iYsz0S3LeHHFTngTs7PweiAanRk+CdmpxhWS5
KMaltxoD8iLAvjDB7cLCKU2xpeIaC5VpLxxTx2KmIOGAWfjNYJbg7qNFK66b66PGIo7qmMNnBPZm
DPnEnWgaHRQLYf9v1ZXjl8sHVIOq33V9j+2Xh177dBlj0E9l9V4g6VVqLuNhW4EQ+1S1r2ubryEK
wvBMOZptLCis1TMYJr9OOI9FN+HDr3LgKFQ2Msa/6ovIVnn/0b2K/cD7cssGsOsbL9/lycs1P7Ls
DqKRH+K3n+OR0rAH2xq4QMwz5oZdTMKyWoVvPIfq9qkjHX33k277j0xJB4QeTIOg5NpKV6+BGpMM
NogkzeaLAugaYfformKSr7Jfwh5iKv2MwyHWEgUoHEZV516xezPk99OtSjqob+CTtrr1HF8o1uIp
fmtkVzzIbazCpaLiEjxBE06RMOgCypnGUYMcpT5KL8PfCSGlrQ6RbJA49Ry/VwcC0fvMRwSyHP7E
bYZLCFYuKLTHkjRgAB3i8OaQybxMRWOEztvjQZfaFO+gDaBozymyPxOH0cfBqUYlgzssThUDVkVh
NYzp4K3x/T6a4VUJfx8cFzAf60NWK/Ldi34kyaK/nv8mG6JLtZXZv/z8fz8fLuDmGImnRo5bQowc
FL6hOVsZzQDbo9Cp5Pfo1BLxf9Jej/40sdW4o6b64eo3Z+2Cu+641ifoaZxp1Y3Ce94PaXoyoRsV
ty8Cspk2SmoVrxP6FKdYAhl2pIldk9Bof8G9AI7V6mN7B3IjA6ly8dSrTDY3y4jP0vF0vDF30WQa
Ftl88yQHQD3UruB2Pb5JmCZ37jKwMM+ZROed38uE8pm+oEwFrhz9RgQSHUQ7FdUlhXNjscblo/+7
zzPwb0dU1mr2sZ+Wpj7RbRYNk5qk/0KDlZcXC5qC5mzTNuJF5O8+7Xr+3PBztWFGuBFPofxGc+ih
v/qi2EB8sn/aIpj8K+kAea1PTvsbH4CRTRRDkxNMKxPjGfYIPbQHDM5KN0yTwc9J/CwAG5g3W5kP
7fa030MvEyJG59NfpUWn3hlo4IiXtsrsj1o3cTb5rfZy2hAA6NAAI1U4JMRUVB/qlCh6hCIXivbq
0FX+yb9NeRfblDeNJzfjp/4bEeIgC5pr4hZA+Ca6APhRgwnCQ6Qhz/SVLifw7q49Re4SIN3ye6Bn
o47g8pYlm8W5EPEgnSbyDmYNLlIPAXtfO4PQdkd7Xnw43xoYxMR5s3jko5gTDCCLoiNKU+dC6X5s
+LXp+ETUxSNYY0/1d2s/6pFCXc9KBMXhm6kGZxHa/QMe6YgNmgydmi6DsGlEVnfS7ShjgO2IL1X9
FsdS44OGIIpRAFUYO143XLb3J26IUDFOfX+tCQIJp8KnUX7zJv7g3O9C5yxf/Wx9zIPLbfcykuYe
PvqaemUi2wIFtzKNDlic2ITtkMnuOAgdyeSdneaIAfj6wjlhIY1ysslmowvNVnnlfAOtKq2UHZDW
ngTKPJstyujdOsssJnNekeocNLkyi+SCPlB11a7FZEVZRe0LX58UWu1i2xm8b4vnmwI1U7lTxUZ0
6BHczkKApDURCfoc7s7nEVMpKbKFzACv4luG3UrcstJduKANh6Z9ss39vEsw37wSmrw6EyaBQAiP
bC03PNzjHSf7vC74dIuvmItCFwo0fTPq63UqwuTlfz9HsG64Wh4nzr4H9QZNJffb4F1tOLeiK9SV
DWUgJNHrTCAz9NmH74Qo/GEMGjwBgYOZPyaGKxh5iiA1d9vt2wEZsnWfoy0CgLO+N8qtskojx4SS
ZvGJj9/G58mylK4kVKWrJsK0jBeSuingY/PE/B96K5Lxd84CFJrjlfidPlu1y0oZWsD8N63fU1gG
qnlAsIC5eoQmRRwkpfQR+VOh75i9zhDcW9spabkoWZ237V7D1jUydcBHCR7LhyfjZriImHHodd8B
jr1WLDvkKir+qX+hlirtfxOvyw2Zy+bhhmtrVEXltxdWs7YVxAye+45LuX8nA5DGMmeWrsU1TUta
W5ExcOaaL30eVxFPzsOQSy6XyxhE3gnLCqL083Iu9h0GgKAA6a4nGpIF9waqL/IzlpXEf2r2AGNZ
TsfZ2yYJ1+JgNML+pEKCgjCCrekGsTr/DC/9GLvL3lstQSJ4v7T973RTAJr2OM5TA4Okh2r89s5b
rxVLUwKfrpNqmG4MM7Cf7q3yKltOCGxVPml9qMOJuchb2/Xih4i+82rGpHciS5/TjYsP+BHYtqG4
n6YXbYhFWJ0td+6txR+dlcUoI/x2ArEmXjpilPHYgkeR77H5FOUe23uIorcpWL6Hld62nMkTPXLb
4vAeSiPYqfeJGs+8bbPe1Gwskj+tUNniLsznLMy9d3EtmuiG26jSKajeNSa28c5ooF479qoNhIs7
f2A2m2T0FGsXl8Y7MQSHzLrEsyvssrfrpLx6keMmbcMyjI0DeiuNbaa4HkAOG32kSxyGVMzoq9tq
0PsogF5+UqlWFW3wDkWD9PNZ771SsWflywHpiyoUtj6RkseYP130e3YQsHB3sgMZoqofLq+gIFTJ
vvdLXLC4e48v7vm7qiQawUeyq4nr9QaUzx6KFNA6JJ37+9FJKnTSrHnwQU3LkZ29bCi+LUSbrjGY
Dr71Duc6NlEnqDsQ2dDvEd4meYux2lcMUba6z6k+ICBfEvuh1u/fAfeow4lpwXRvbxtvKcywlsA/
m2Opm/Ww0/vYW1yVbT9GBumadvQ9VUgPhrkynwrlXGLnIv2n0rHXmZKNh4kFoGenep0KFFDCbW/Q
0rTvcil/8wo4W3+c3aBY4Xb3+pabZoN+HK3VBxLRhngYOV7yl5P3G9KRF0Sx2YAwUVP5qG6N3gTC
12dLyjt8KZGwDJW2SbyhfBVxneMZR6hUWwZ/yJVUNoK0ko0UkavC6kMLeTBtKzgfRQJEfezMdPHA
RF58geN8Lker4/S0tJKFZ2J/VVhZuF9h4BPWFgvDYntkJ2kYvINk7OIOTJ72ni8C6a44/en67lYN
YZNAUIYa58+E8QGcGkJLYUsyNCoHkQ3PVUt3rUQo9mwDK0FalYLUpIeGEZfjmVBLPPXbtQdXKiQE
c+0gfFzpk+QrRqHvpQCFxNyluyhH/rd+c9NdZMsNo9oYzG33Hsqte5JHmMDnrL6FRE8LM7BGliSg
MHzBDujZGfScabTJVKhBJJxNhnGgULtX33nuwqBjn+zRHXgV+SyAjcWa5fBWcc68tJsyrOd4P76x
HKSIOKs4jt9q1qp1ucqsLMorFzX5ih7SFGISa0FONtSoEH49GQpLhlqy6wNiXXju8esSKVQEcmkI
qPxwx+s6oOvVPT5lWrRhA4yjJEcMF45TebhxEtqvX1Q2feJHse4wpAkTy+hqoBV/t5WpcWMyEf9N
0LRI05BHICzTqTmInk0H7bAbNyQ3Qn07FJdSVQUumYJhNm1Wh8knYObakUVGGlzFdwIRgg3O8IqI
aIOrQujzE3ohenpU+QUmGS3a5PNDnEuOdavWgkAXnaymhE69TOgDMKdfAJrPpBaeCDPiW18z4Q7j
9xKz0r1F4wOADJj3REykVMuxcUnDaLXj9xtujtjsL61YWk8AOcrhOjZxt3/Ty82zusXaBdG4u0qe
dJJKrRwcgYMSQP+1oSHIUQuxxutx85Ord8bDH32SIo5FNsJZajnL7TNRdaOhXwx1nNbfZf3txAh1
5Mo0bupdqzsSaGsESQI2lBDMlre21jHwZdVOs3/Qq4T/LsabAx0c7fer73EjeOvAY/Cz4/fkkW8H
dUOuaYPDToQVULAE9VJ3OytCxYQx0b7TLOcO0Vz8vxBDI0usniJfe8hQFIyZyMGX+s/aYbr4x5WV
KHL8dsnbWF/VJr2QODWUE4AiIgzArllVK2ynCGz6d9kSAk/MNGLym/jfk+03dseEOxLR+0FahYUm
+3W9I2ybsDtU1XeAnV5nTAaDyzWNlXK+Q4poPNDNBD2V6gZ1MWfVZOA0LPhWAkIq6UvmsCj2FlQL
E08ivbiY7ocy3aMSuJMzyfm3TXy9EXBMuQGtYiM4Tsp9Fg0l5zYC1Ups7xSVxyQK3oRym2jxwvlL
uqvMGaXRVUCVC/cpRlpWItQCAeLLmgO64szVWctG8fHcQ3kOLTALK7Kj/zpVPKz7bch6UxWvX6tn
YJ4L4Kyd8YvVQL2nm4m+T4h85ZaNi3UHOzvWTlZI+raUPXXENeWbMYEvv0Gx/o0d7/z/qOpHroR2
S+oSPxYISjObeDkc/npNr3c0skmKGwqEm/ArrQ6D9jfWDXAEZbCjwMdQQ4d6TJBJu8VLlyfcTaaC
KM9loA0IIDM54PSgVcWl1rsNbByMjLYQCH4ClkUQRWenxwfACTkKbYebl5Y/pFFSxDgmec+Ky9Zh
lQTRr1+BpYJg1NsJWUc3PWD/6wjsGrPp+hDqk3CPWjj8qYWZ6NgtYh/BsausUW/sgFcfHaQk6Ql9
PcBF7pmHKZBvv4CwYZWWYby0JYzU9cTfxrQSl7KEH4TYaJ1uSoMgOQsf8y0LkJdm1X1B11F+2K9y
HTAU3vyit7RY0eyihCocy3nWXmX3H6mFMC9pQeG18u70ldFLxRCiwEzzlb3Pg4/WE9pkJjPLtSa6
P2NhJKcH7HqzSlPGlvTcKLstrBOQnM3mdPEM2czuYQt5szMPD/qKItyETg0XWJMIVfbwY5UXoUQw
tgB50n6JtdhezjSpF4qWmPuPlI8KbI6WoxV0MJedo4WeUhhk8I3BWYGBiJeLkFb82tbE+SOQVsJo
ZAzKd7hdT0bgAHGM02S2iNJ4jzOcgtmVL7A+//9IJkbjpRIkSGb4314p7hclmU+KR9Z96hXHrxCi
pVT9sOUIMwVaFR5rGARBx43QnRq42D8n6qK5q/3MkMAVnuge1kkCbHi+V2yH98NcVCt7r5GvndYm
Gt+4fonRpeTheIEkuOn9SP4SXmBYEJmurt/qxfcMinkyy+NQfsMXhW4i+0QeOXy0t7f461xfGIN6
EpKkj20RQYUcoRIlb09S7uyRp2u/JHZ/cXSNS1XhAV7xFiAeXPPXOjrq+p7LmOSsDVsD/SEVT5We
GfoiMjXEk2ERIbapWF9S0EP0WoIq+ym7wJtWSeKJIKBRag9jiATI1tmyKOtmr7aoFiNA10Po3Dwq
7lvVD0vi9yP3V8WsV/C2i35qGTGbYoe2CP4HwNDTNpcJUz8bmrBhg8+afxmVGAIwp+auvIVyXaSE
KLLyvE/nq9a4VC+ecWbtky9yqNy8/cu/Zaya9OC0v98tCs7k4voevy2hy0W1rORgZ2A8b0pLLpTa
PSrgWO5PeYI/LnI83a305IcGHpZMUgf497NZ+AsNCvSe7DLuifR6rOvzrtBZ77uqdve9287D6h1F
KraB7Y6Jo/zNmA69053a5emoxQMw/gUD/MQR5BijlFFSsh6OZnvhAsXppwcIJzcsMw8pnTWBIKpD
YyiQ4WzApY0XpsresbHOU7BAsW6cjPiFdtR0pqw4l6xGpDpx/4viD9ZVFJKFgqGYJ52Yc6yEz5Oa
A0+FCPmxIrwY+s1duqvyrpU5e4aznYdNNf0+Q2Ggl8N/dDOEPHuWkzAlpwd3POIm2heiluyRdQTt
8yExxynCXqnaArUnTnb+oYFX2V9cgSyy+FUgCoXTLC6ETZHBpDcdo+d+2NF+4bN+fB9ht0d6L970
/BvOUAUwDzeuezKnuJEtR4Rf9fuJyw9LxtJI8ZxYeBKa0ObDlupS9nPhHOfMRaNONo/8guwDaduC
IMGhNudbKGF9ehGVdE4XLKjZ4+vYe03ajKYJ+jvqmchn9MF2fAChhLQFOWJIMu1Ini5RII0eK3Rt
lWDqi2qzi7bHSzYmUflg53a7rhY1rJgpZkc37RQE/eiO9oTCPL81VcmPD0SHa6RGStAeBYwTD/UT
A8tnAy03VrCT9sQzmnqbcZQwmOQ3Vgoxvytp+U4Vyq66N/gwsgB6cxOYgmxjl84E5zbPBw2WDglZ
DNpuQdNAemqBMfwUljE3wnFvP3bG7gviU/kR44IT6A==
`pragma protect end_protected
