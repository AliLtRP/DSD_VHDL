// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Rcgeba9YIsn6JSkx8blDxZasByj+ensHURGbsHpHwkY8O0qdnD2ftRlg/U38C3Go+yAY0+XhAHHE
Bd2bnqQImuBC0ah6bHYHjeMuq+X+VUHwpq7Je7bn+kvARcwznV2sNHIRKFI6dYCcPlO/324Gafrh
b267kg1jO6y3BamQZhzxw7inosZ+uro/1b351daZrAhV9ByY1nAql1J2gzQ4vnQqlCfXhoaqrgjC
Gv4DniFFm4lrZWpoFxfVjb11JQEdtkoqm6ptlYo62NapjURcibkoWBbSXb0y2cxXhwba2e1ml7kE
w4i6T2+VY9aUe4CRcydej/kHTe0DHaM+Z13/Vg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
s+lzo/7azM7qPeqUJHSF/JXuAX+7q8ag4WxX6KwFb1uwfdCLkPgamqoWqNdMWNUsOudqmZ7Ga61B
YiIdEOwlJ9CklPUW187ioqpDWr7PtmdFMAZs0ZYA3X3kyMx+/gzJxTYG8dxb+m4xybZJZwKq+zQH
p9yAL/C/wUHHzCCXvtpQ4ECj98NunI3kxKhyG0YocOi4GCkfgOaQCTR188RsSGHpe3MM59DzTP37
sQbcj903vDUJulY8YsD7kjfvpb0IUk1sVY05F/Bzk+UtGJ6pVpkK6gm4VZZS35M0Srz7YjQHbkMp
GDg/avExnSh8iQ9qxfWA/fbiObKcV3X1sf980+BrSh6zNK40WT+YTgQma3OiwzMLe7NU0aWXLzzJ
yPK9yvWjVMk8Q55A3W8CkbCQsuVpHwYcSS4xcJ21oF8bOCwty8Xmkn3YqaWh3d2fYFCKlL06ixYo
hTiqHDpgU2p674kpFt7jmxVHneVZxNdKa7AUsUlZP/q6lVVPp2OZsYRYQLRmSxdZL3il/A9P0340
PXOeW7d+MlH+oqT1X6DUvxGQ3Fw78N9cJoFSAM2frEGTuWlLrjFJBen5GKBW/NXsj3tPBSXdDHsI
V4M0lOaPkBivCGfd7eOqnFtAVJdgN/v1IRauY+kcf8fMyQq6ygLFIbr4jDtpaX2WYYZTYxnIwX3t
jIeUE15z+XSL3JYmKnrpb66kNpjlOlR1HM+CcvFDg7CE6ui+sTgxwsFzTLh5BdVjqdsTAG4hetWO
9ccSFIHV2iS+54gwjwyiVHgE1Ur36KxtwpjbCmTJgA4S/tNsLt50hCvSMeMFwqh2L/xl8h3k2CsD
0NUavBVUyS2UajP00tbbMsHy6j5NkMwRnM2Y48L1gEbm56DLfRyIvE6DoVwLIJYdgznYDent4ecp
UTbRCNYa/ay5AqhdwhTnJdziNlq3vlxiyiHgheJBRkq1rhqCtlnUYZFa2gmnQuKYE1GiIbZN5VeQ
GEBJUfB8fMg4paf2e7Y71ChafMyJHpFel+TRKSgc0UzFH52Y6mO0L+jq6RCzqQfJZ7XAv5mz05iv
0T18tbI897kP0HU0+ULHMZ4WICa1t0g3wpXAvzrPdhwsMPqpHwZQol7e+YV4udI6ijam9kaiKL3B
3z08zcBAng5ehwUwCQOVVP56CeUpA89mPIg1EnvvD41RqDxpLgugO0w9k/XVCk8Jpj8LtlK4VXa/
pZ1lc9KWS8eyut6Wb5EgFPexxOWggdNmcgcn4ThKDUdW5h9g0fVEykjU+bBg4Ut7Fb+do5kIVb8Q
nR8DZLgTDmHPDPh1RGnkppS5W5Ln7mUXtWh5YMNUN9vJJWHx10nTKgbzWtfHya+FCzVRNFRQA0/R
PlrPZH9Qg+Pauuar3EEFDOEQGrqkIj9hTOeC9lIC/7ZRFB+x+l6aiBtR1tl6sud7fIh+61OXJUwf
0J+GJTjWk3RFJ4zYPQUTXPAWCSztveL8ufiQ4jOTqmtvufVB4Ysik60cCRIsR9/L1pEH0wuypFb/
tF0jKvNUn/4/6jCexd+nF/N1O08ucSn6+cp47rMDgQBeX72gsFJud+apVFDJpbIig11bFgqHyRDi
yVwdzZGe0xPrtHFIuEDwRygH3cckeKCuVUczMxvB0L0QGZCNblFVTG73xLpC/7t7YbuW25Up78PG
wV5ReJ7kLJYSbuYv4w+Cjz0Gku/dF+HVMql+M2iAr2h3A3kQaHGOO2sDWHk4j5hsw90JY6pktTf9
sUCqDDgzWcYdPzngbEgwTL4LCoMJr+6XNnDzGYzJwxltxkXaHNQ5x7pfurH1y7wH/U3Uz6FK+Nhw
ZjO/e80sYK+R8KBwiyLaezOavvMNl1GTVPD6y+gkx2l/fo2icorBV/yjP/aBlRhJ1pVgvF3RTSLi
GYVk9IuCyYFCE5cffJ7cJVD3r4b1SspYRovDRTbsv6FWfaDjDzrIrzLgaqyHptulemSpgtGyFSs4
DiT50+YfMlY7zFPLy6EVA3wZKagqZFlrDCAWzeAFceIgdCvMorow0SfmcRkJK/514TObVTVG6aC8
G5iDNTEcBbLLFajaHmVJFNapaV/QO2deWEfQblUWBuIq9UM6yRgPp6eenTzbBrCTc7TyjhoslJMM
bZrqB70VSPE0une6r2SoJMga3bsMfREU7HzjhjVu6HdACNNJz2fluiefZdeMEhpiJr3qBErkKyoS
YAD2cf8rWbBb0v+FtzzbqD3HsrKoRfk4OyWB2yR2JQ8dgZAGd1rT4UUi3im0Q0QOiABo7JeZeJ+p
7HQaX55Obyps0eFUVeJtt862HS9+aG2VyDicWR6O5Egi7q/XIEIRounCwSJFWLH9Oayocwsa/fiN
iLSgpROol/jhm/aTsxx6yj6J4n77hkJ2FtNoqTLXaCGpcFhQ2XI79AYDCviFtMSbBMIAaBEWYj4w
3Bytqjy9FhpRpVeSVrq4WeLTZkysfeNG/Dp20t2Floqgk45JEH+6Xvhwbf9bpTLR6WiK0S7vukFS
kpa+MIOxW95Qov69yNdJpurdbOTtAoOCeMYSP43ltUCAr92ja31fvFpcC2IRTx+Euhe0o7RvGKys
UhXg8MMophRVmjCzO/1NxXUBxNtFxRLYdtlXKUrvPXQxt5l/XkrL+srnopp9PY43TSg/V+HOYK5z
bZXo3dy2k3dwCFQSSNnZ834GqDNAMLNEttergJsfeh16+NEVAoSBF5eKJNJ9fgQ4h1XRAakN3to9
kDclJdVIMCm+Zg/93RauynbueX/b7+Aec7/1kpNtN15PEb/0gJ3ncgr8Wj5tlrJkhLn3UPgPyNbF
FWge06vMeHxyOMJ5tcsis2/zb0DMGCx64H6X4vo+hqlH3OOlMXPPbZgmyqccqCWuOMXU5ACKDtkC
CboPrASE8ye+XXuV7mQRjcfcHDzECOYnclZV9j++C8ab5U9ZrlNpv8BMMDFWN8zqvWERwkfFlo2v
dxLqqgrEuc35zFmVcXMfhemizUqtQ1jd+WPErPfxzdgTWh4ilEMMsZoZ+ObnG5q3dKI8NEWeNARH
ZdUS0foPz//OmuNvp3TnvpI3NV9kR50o3S+96F/dqMVrk9hS6qgSTLjtSFxK+yTyG/Y0FHGBgPqO
Cv1GLI1f82H6DgXliQv6Y8B318rDgZirRTeNSejKN1W8GhHB2lLBvsR1FEkxnY5y5KCk04T8JgCY
BvelPlh1PQJI9LdLqfQ+jyDWBnV8WQE5uhIpt/gHfwDktqlIvcX8KmWoUNJsxzDh0u4eg6Iaao4o
K3w4u2d+MXNXOHojgDObfM1aXmdQb9G9Q0B/p9hkFVKF9btnT21OG2INJEzoP+Qbf1CFArHFMjFT
sye6eeeHuzmfrnOaHIHiq0bqhBg4LRnLahuHpfNOWA/AlkbQheNmEyiuW9P/A4l2Fi+4AzRaWsJ3
UFOhuTIxzR5hHMoRJxlInKHCPeRzY1p8w8DCcecWjBdlByf95AOPKAeAdE3Y4nPZD9Rs82BIWIce
iHTbuc1NuC4sq09zSwl/WvqlwtnKHN5xVtut2bkzAU/344J9amcIIrRcOStrG0KtDQBFxVpVK9zK
GlbWYe9DejSxGS11P1hGkfvKaU+BDiR7NYQ+UHTeGrcL/YwsGwxq8/mQ8jGNUlZ3bxTFCiz1LYai
L6w+8s94LC7XwFSCr9kPe+9pWuszT3oPLzWm/0ncLHf0wXB4Cet8dWw0GwVe5zQjjl0T0XaqWT9C
lI9nfhzmXkAAA+ffZth+US+eSvrHNAA9m9zW3JYsEUQ/29v/QcmldOTMmo2La9PmxTv0iVyNG1RD
bVgnqTTmjnUcyXSfdz5Sy1yYG0nHKHHBFh6d5cNywgL4xVMlBLyv+/zLvrOlgEWwf5fHV/jqzdSS
VAupeqwDTN9+jEY2i+2q5oSzXTC+5TkgJ7+CuclIucyt6AunpBFc+oJMWVWTwoP5UhQQuLFZIVgI
lApC7XJX3S7G79C1GHy3t7vEXeJLhr3yStksHHWk2L64e/TMnCdx7xIxbzVK6Zse9vQCu1vyrFgQ
iWYB8xVlpxKrIHtKMvfm/6h2L+CzTQfQtr8FGoXbrlAE1Lpsseq8zOFbNkPfWMfqHSRDrxNRg+N4
MbH6Ntm+txZ3chbUp+8hXUbYNpXLL+vUsR/YnX+wrMfQ3yQtS5OF56su3RzNQdjyp+3IY/3qMDaD
zgE6UUegg1CI0MJH0fwlNhPd71D7E0TjWU25W9V7IDR4ES+KU6hQdQt7IpEBa+Xq0xZqU0ZzAMAC
W0ZV1YQg1ofCsBzw61qFubtlQXepijwt6sXx0vZEdS9P6iLzI1iKgmYFKMAHayUXEK00dZxzEDxJ
KTo2h6mV1jl+Isy50bu19BsEdiUGWNNM/xoGrftTmgNgjEDvlEQZ18UUs37bkMWKCrBL/d9jNF1G
IYXzFwK6I7exZyNeMUR3mHmLgsGz9u8HG+IGY6WLsCVumYM6K9r/5lKYFlcnvXQ9+p2NFV9nIec4
cYJmyPvR7r/5OP34NaF05C1KkdomLySnkNyyNGvJkl4rmwG43Pl0qYZq1W/nLvfkyugZ05vEoUSw
9s+XapLG1WACb3cqP1MsYuFrsLHPgs39eOAHyMD9PIXx8aasAOSWJMjVawM9YYL7+5f9kEyPFKw3
UspqV4V6f7XuL0k4eBBsow/38pPNf89ULlcG00RNZuvIq8Q/cVP8dlfN/P3xp+GmcRK1+zkYirtm
Va01vja+NI4AS6yHdba1NV+/UsE52OywEpe4Tvf6v1sEexV/qVB8vRErvg/dEpPRoyuFeY+YDLP/
+KXY6LQ5SVmIpojxrCbabO99hW4vNHsighPEq5eqqxj+5hhRp8hcnJUwmXkGvXhfTZNxK21OjQ9x
jPvg1OQ5LyI2+btAuJSzGnU2ds/kWQV7gc2JWsuWsF4R26MBLsILH6othBsySnpUOopUWokz0pON
pn9UWbB5vi7zv6TfnO/ZcdrRwoT6J1LE4TuVcrv8gdKUitUR621chAYC8RPuuABzVd1tutaEqDzB
Evb+VQDKBrAm0wqocSGNXMQkBmb/I7XubXrl1uuOihYWfxOhYSk9v7Mm/Mx7pJEpQbZgNBQJK/Ue
gzpI34AeYZitUl2SLK7WAtQkXmcLw3kcaD2ZyLJWjlvO+WWSQx9dvWaTU7NMc3hgl+OCt6EKS05U
BZ2aPr8zcbbFRNuYLUYeFNYLMg0W73Zg/HnEwaSD8GyF492HacjqGR0rjpKjonsHl87sj2ASCzfK
7rWFp++FVmeVsedHaBVLXwPaYmZhBt08FanMzjPJfsjjTqnl0MbTy5P588fB/oX9KlQWHAGlxybv
J5oyV7GwaUnlDuIPEhRb6K1U7+DHwIQsegHJFy8N2I4gieIisEFU7rXQcyW5+oelWhzt5kTzl7+j
tsIm5UhhBbaPOSA+8GOzUPdc7VDPS4ErLI29qbAYy+kmbDO2TwVjigmet8bjPxvXr/R7Vu5shtmw
8MbsJv44vi7YTAp3FsgU26mAHg+k0PutXs+fZWR+NU7PcHzTOqFoUAMLmJLpI65AHfHXrqFnVHzZ
pRT7FXIFyh3Ud/bh7BcrVi+IbFE7TGVHqdD0YQCd8ah2G2KWSkyV++AX/ju5kaHA8fHgNQwJJgIv
s/U8w9LsGaLUjYs53gZ/VaGf62XAo036n2MdSRfNOAyoe6/+REtjKY0I1DU8C4Erp3lUexOrQmE7
ouhUsJpAAysf5/cKWiGYjB/6IWuQLH6H+KV6aQs8NyFeIqVFqGoUx9ugnwXik31ypQPMNXoK+UYl
B+HCLainrdf2KFq77ImPf8vZyf+D3RXLnMvWUOyQEXf2g2CAdgAferxnobSZ5pvosndXfupELs3g
CY8QcJRXcgb+IddupbJCG5ZYxpvVDpXogGpDUVfj+hEhBm0O9w/sOsLMREbnvKIeB/zi4pQFcIYe
oYH8WitW5h7xiWYKR/hqMa/hj+HJwMNCRHp2ILz4M1dDPjMpVlYs7r6NQZK8+n/Rur7L5SzFHi+A
7jhxxGqGdGmkT8RbKObcqGQ3CGZqotUG22O59A4wvkyklq9HEW9/kIe6Ww40xq1S1VQgoaiN71qv
seMlOh3dgZ/FgSod0vxudsGDpbNAH3MRSYBowwlE+lyDjqzZ2YEqSBQHJEimkb3sWnZLF0nxmRfw
L+EVNIGkMg0vx6Gg69doWCRkC1PBAQwUXEYvwT4Q3hVpiBJBJCpfVm5V3eAUVnmZKb37dvRrco3D
5qPGZSoP8OBZAAP6Fuln/8YCwFh6DgRtnMDHWiO2YTJDZ+okNl9QfPe0oYAWHlI44D5LCcASWM5a
S4JkIa2s4dlc2+bqDtShrPe7IQ2LXp6AKUgOfjmmKCTb0Gz05wfvni/yO/jhCqDXRruj1oLmee4Q
Iei+7WzsMudsvi1t7HbwsBQQqj7hptUc5zpHkzs9TADr1PLmU1FwpVZX1wRHCR8Lm6uuRc73q7Mt
ahkDO9F3M1TvwFHVKkLQ2klChWR8Nj08j/UhQa0UViomjnV+LZPU/5rJQ2ww4dXiSxnwB82ZHgue
8Tgf7D6mq+BsvmixOmR7AT5WjMsEER14zc1Ap+iiAeK/aZN5TLMvQxchtumzv+e3/nIlV/VcsfrQ
oGF/BWBUlkRLQdI4GZXGj2z7/WK/dIToMrM9QCBuvtbYfDf//9xueS5kiaYxn2Z77bnmfW339NpI
g0xPVP1SH20ki1BLfuD6M9f09e8BJUIWvZ5fih2oi2QT1ZsRzYZhQKelQNAwxSUlDwgjgN1RCmuT
qk19lKWFOTK2flCwY6GfOArXb9NtnjHDUsjfBgj9TAC2VukFEfUY64dxmk4/UxAwkRpmI7ninCxe
i8iXxpHFAWWcs4H6bMmdLGCDA+aDPoWOjsNN41L6v4V1pmXQ0ya+EA5llo6VMxErWwn26gJyq7BA
/wKR7lP1meM0Tn/7LOEwqb0fSnHWqPLWLMvvBMCltHK3EsXwInIadSlyeu04j6zB1RqSA74FRcRc
5VhI+b2BtrY7mLjvDhCIOrAgAz1gvur1kReFA4johGVgwoFxpT0IsmVsMsRT1jKtnJ9dpYTIrvYD
WxBG2oFhMgbkHG2oBdngpKQK5pmhmz8YQMHI+AdOacRbIrH3FJ9VsiyWxM3rQabSovv+GguTjIrE
9drprxO9cZaItHYeReJRFKiaAieETjd5mfsPPHJmk1fFwzgKGsGlJl207d1coBxeQtFSnzU3nidL
Z2UdxXcFQauclXDBL5fBvgAVE6BrazDIKi/VvK9jFA+cIRiX56Mao7Wuk3X3QA5I7qtLx0gYXI44
HwAMJPIwH3HgDcjFVWcw0VyOJgHoC9kZLxI0F1eaImhWbkaj4uP9yoQYKOkCVlvv7hi+s5hGuZ7s
Rs4OX2XLEkOTlc3LQbkwJKShdLoENvI0aX0zN4zUKhbEMFCSOe0zGXPxhd2rauprF8lc5U6h415b
ei4C2IB8RqihzQSB217JzvttTVDfFhraGEXzE02ACzizFYlPaCFBDGI5uvUnErWChmmUzV1xC4b9
T4UP0xh0fGaxTDbzZFhZ+ovwVM+GxXYgnzu1TJ1cClsjTPo7BxSyuzRW/fxPvkZ7KN+zLEvYbK4d
uNGmk4ZKL3T3KcrmkneNqDUOUlxcy/kjCb6/mWuAZ+/KEtNpWRNks9WBX8W5Olvg3LeFcnQcl5F6
mgclQtBa4a4cY34fEaJtHihY449siXRoVdUkv/G2JOPBCHRBvn+rfeS/A9hmlPUHqD+QmLgdw/zy
JBGxRTB1jdk65eulhelVj+rshzOdjO4YGm7Zb6qDAe4JCqUMCMPIppvp1oCPO4ebq4/FwCSnf2yY
0MC50cF0YgXTQDBPhYsFxoVKAdutkKtvf+F1nhQTZk0UtYQyBCo+Bnp8I9twbUoQbP8uP8CO62S0
QML82dQTZrCv9Kl37s/Uw319c3DKbiyKkelHIYCvMIXgqbC3u5EJcakOM0eO7VQtiqjMfNuczNTq
3dw6p8zQ53is/OwxOzMszzCuPgL3KywWWTcu5fNaqICgQs7my1YkNV8fdyoY0igPkRXVHGCVV3xv
5WXkGYWu8Z3YIHaB4fUwGXc4S5gZt+vpKoUc5SyS/HOO1QsojUTrh6IPknsuhIzNixX5llLT8P4J
yFy2/Bxm8dEeFwkOp1MUDMDRkaCjfCGyMNcSzcA521/5jhjGcbtf8qM1GrPZ7K1lxwkB/MpXXC+a
S6XrfyYoHfzkp2spVftZsDBbIRpLHV0lSj3yq0UNFPOn/bKR0imGzShpAx2Ix1T0vJ/PHnfaO+oq
mGMokqg6KZwNkSrMuIWWj7UFAOfQAqsg+mL8ATuO5ddp4M9zU0hj51+Z+D4NONkQw5gxdN5rXv8h
HPFNWAaO+1RA75xNZ/jQ1kAl7cpXvDI4y9GNxaY8u9BuFv2dwuBYcJ56MVzxONROuzoX0mMYUDa2
J8UcO+pUaclgKWIKyzHonMO3tW8CdWzNPg+RP1DFbJiTc1Csv9H0u6xYl1Op6THg0IxtcCbSpgur
/ET+6/fyldXGoBkC1K9X5uXUzMXu7hZa4ILpqOcK0/MmIPLElxoTX5vEVY5Xyd87vmYSC8qFa+xQ
bpIvUWBL78UA8GaYrF3VG27XKeeI8uHubqDvOkYcyGUlhHM+QQvBCd9yOHq8FTSpehsyJdHTke6o
ljfrMtbXPDFC0+EXBGz6yAotmppEulDd0X7sbqJLZwS2T6MmN/QtT6Zi2oaFXVfoY09TvjQe7TqM
wKJkzScJs3HQC5XNdbE2wPsLontxH4Tf8LBlndYjJh/wUiNEzOePl1fsiNbekfOEm1uaK8KMwztI
IArm0ZKo1KW6Q9cb+3tPbzVV3w9TssPK3z9rNpwIg3H9k4EM9HKtvbtsaglUQKpZ0Vwq8k8BjLcw
mRxEz29qg5a1gv8z6KQbnYbe2+860jRI9QLQviVtYFObAVM+9zh8h4H68eQV69EqtdxRwH4JFyEK
Wme2Qp3jwQDfZ88zflAUniEg4LE6jpDnaSs9rAF/saKu4CrbBSCBfF6wUrLFWcFoMU2RgqQwqstc
3C8ux485uYczLmJXFMNDeNp8cJSPABrWDzg6Hswf+VoFHKaasJU41hKxYGTN0CDH/3w/SR7C9YgH
SblO3XMYifb8gOygiX6peEWvEwWvEstXr2kynekK2R3Tx94R9G3xcZD6qFu2ux/5X1Nry+6z5BI8
JNo+2YXVd0x9siCyOg7bs1O/5XBx6aE+coQQKK5YclXvG9YL7JybVuylPBhsG54fBefWaqMSBVXi
gWeZh+KnTEmhMmmx2FKDdS16gB8fIuGoBOC6UoSRlIiRDVaN2OL0S/bwAxmzX9rJEvcm53yUi7Dy
hq1K9CphrtpOp7fOS2FXzaTVsRrO0fm/2Fycb7MJyuq1Xp72EDHfwZfjwrzZ6mFrh8qSpcop7XO9
C/CBWwxztps4sjUyIazF9V7Q4R9y6Sjw0U3oNvFLbVYrvx7SrKdyWusYw5be1/PIt8xVbY7/DDN+
AHw/nQolj1oSQWOucmM2T34/D2qIpaZ9Xs35N6Zp0oHvGf7UW0oG7V4MusnmdNRQiNpqmoyLVyRI
UxGiXM+apNxAW160DT5USJ6GwMroLa8bFNW7MOQrYy6d0XpkLzIe3SKEPivAChcpIQpdfRLpK+Vf
baL6NPQtWu4XfuB6kKFVYkQbVoEvhED5Yh9nN4Q5JQX6ojiCCeotWcAlfFq9d+8H/nCpO2QKKFLB
hkl/M3BIso1rOeD+tha9Er4DxZ5IRMtauafFFt16jNwtPFTF4jMq/OdRXTgnyylMI2E3MX5ETRFu
Xux8zBzDvSzqfNOsGQt8uacQM7yL4YJcxdzmv0ktsNfIYBUrfmk3vMXOA+7A7QkPtpMKKD4oowHg
gxyQ0XzQ45jeNaHsyBnSgfc2D4w98XPqBJPwXvJXgm7DuROd2/yRRlY0zRFAT3gCR4jwBakY4I3F
+legyIHKhd15V/s1ErZu6PmNptlSZsoIwtXNs1xNm+mo9XvDfpz6Dvj11VntN/I/PTFka6qso2Mv
UDeuwaWxZkZFrOyFUWeTjfkLUxLr8zbR0KTWtwpMhuaA1dswAecuV1bhFyazfLRzS9F8Rw/Z2fAd
gEycMjjsUSbrUJnu4jGS7+PyXl9G+q2WTk4ZFmJ2Js/wnpqeUVBB0FmJMqWZYgd3nwcj/rTfUCzI
GlldisM/jN3kF1HwBMsvHmk4bSrVl27/26P/8LEYXDFnMGH/CtAHj0ynZmdCFWbe8pt2HflaPHB3
ybmM+i8lMKZvFwNwWgiQfIj9swFTJIx9oq/rTB8Y3oHrVHi2iJRuOMpAdPhiOstwbyRNnS911LBV
uVmfnLmH3Q5+kofW8KXyGM5EHl8FXbQ38p6flKjApZfNfY3kuORM13THVmHiOlHaq2XpQgjnlegC
eZcCavIGA+DG2JziROwKJjL14tg9crICegfxR+NNWDZw44oyDuJVdqFJwJtoleIEge4dkUoR+zpr
pPDVxMaM7d8KO2pVfZroCw290flnV+uOVJ/cQusENMgOhjPqv0CQwCZw63w3sO46AhSEIfbWXKz1
ZSNlF2v5mwoTSRRHxOPx4lNbarYEhUPIRPvpcEIpBWosnTo5UD87gN2YEuwyt/EnGiOyu0oCpJa6
z+oQKWXtw4uSnrJ8FQErykoPhv4FJLJb3vtosoSKSla5qt4sfofZ+JPHjb7QBmEvPKsgLH2Pvb28
FomJ14KbOGsXDfFfhzKIMKe3d2HSuH8+hp4js7D5ky6qi29Fx5Nv8yG5DkdZY0NLFSK1khjxWxCO
DFzuwENm2ZA+TSziuVfsVX0/QHgKMPkMjuC4yWLNRxeXgLj1Dp1wJs8OgRfkdy9BkBWNAGa1KG01
+pxeEpD15jyZr1AKC5fJ8RFTN9N5+EQLdEO2kVhKS/nnSc7QYMCWUdPcGkULTjHYzXPzsTFQJTsc
BsMNDWdGCmtt8Yx1PnoZs29c4SuHzSKqbP4ls2vKs95zZPSh34FMsh4ycNkIfDVW37wRVJNkTKsC
InMatSI0WiizrhhNXW9gBd89b6DGlWzPEyNvlpsOrzWRC60ue9cj1usjc4vS/59jSim/jre/qsYY
Uxh04E7+/skpnXlo4FkFJPa97rmYen3DO1/L2epIcXngLJ0wUjX7Aa8j35uJIf73Y/SOqdFqoMqK
+C2l/J8i9cl9VWrUJ8yPvqGDwnPjFJFDUkQs+anJPS1UlLliWrJYqOc9xY1L4jy2PmcRu5yVIbJP
H8RqtD/qaYVoQZbvde5zlBy7U3V5cfJvU/T1Xh7t70pFKHLzpUN+aC+QFhAtVZ/IJiRKLL4PpXQJ
r1NQFoiEcRJP6DBDmfJJGw1VQVEAFjrKif/OGV7bZzTjvpDE7bsB7xoopqH/PFFLG8RlElrdnjP8
u6Qp4Tvxaa44mN978r+riKeVauX+W3qLyqcgDL0isrqpoupWtnX/prQm3QjAUag7UFZ1Tm75p2Ur
Arx4f9pkzn+Y259PCj1EvsAcbO5cGpd9NLN9hkcDUeGYfy2BVCSgg1DCfjQgF6S/WCVVXrzcftGN
21pKM+3hao40aZxXVbcq3kQ9k5XH6/Tbl7FwOM/KpyX+QcCFojlbURi+M4az5SBpgQYhEFmojpf4
YwoT+80wWP8N83W5X38YLRiO7xVhnhRNluC95sHynxSarS+kTW3gFKdRrG4v5BQe3iyDUmvZyjjo
LNWK3GXwk7OljP6VV4xSt0l9Ir2T/FNTZTIxU813dtgQPX2U+cdNg5P2CnL5L2XH+KbK0wu7kLoW
A+daXGIB6F3+u0qXJQOiya5iapVPzLI3qHlUJXmjXP+u9xHiryInLD94XpOGkh6KLyf5zjViH4/7
pw9AiGCcFIkeMA68/YTyJkS4iS4sDN7CcLyuhblBu9KdX8ihkIK3gLNVg6/iQxebtyaKnwm3h5l3
nbOm4OQrZ0T1rN/MNXDfNkIhKK67ZY+nBVgti7xhso7ofWgcoLj/4R6afhSOcXf34WfBk0OsdE44
GGtVmKgyqyyflzZrp6fFMIhoB/QVeoJbxncpLD56rdD9WI7siLaDXUcvN3XXUbR1oGupo7SNdG7l
JRkTK/etdn3sryRTpzmaaP8Nm1Nmqrl6OiXkklNjGQfEfES+P4oUcK3TmlGxqwKE0rLYOO27Eip+
G85zzI7QSk0lliUKqz73yZc5rv6NSwb5oYwxhO968VoRofbetQ3OVwgVNUrbUzQ/P4B2pWn3I39a
FTcsIeQhxn3ePxHBP+RB1h7aZdOMOTHaxNGKjX5hNxueV02lq4yTUSWl/hVBEKzlqzzdJtbY/GQH
gDYKqWvBPIXkbat47+dMw6Pp/vHvrMfPxNXPxYogiH2VMydLh0ymWbGZvIgUdpGS/O/+SWMDLk3i
l5+6aZAJ46usnpa3zh5GqXYcKqmSJmPyg9tLCs+YT+ykxSQcoZNA9EfQzDDu6omom5ZhuqJDmLdW
BdZYI73h2hO8+94I/OxWf4DIg41ZAFiHc0N1q/qdQjzdi3FOE8FeuN/5oo/sIZNZhm1UQCKgBTRu
7gztBFp24S6T1kwEuVmXZS/Z0upq1Kfzu/3Ye631FX6v+dcJEHrXeVIGNTxeWC2vLKLwPaaYZMzf
GFB9N7Nhj23+1KEzDKO5zQS5Xcfb5wzQUAI32qaay7EMjKZtNv3w4FXsC50iYbW9wp+rYd4ddli9
bpTlD2Ej1DwwV3CldRyDefhw/n/3XlGfOxuU47s6dIlk8ZjRDHor/omIGPrnmIyPlbmPd1L4//3z
sn0QIGcpph+5NouYY/diVUED1qDX55WMe4dVhpecEtHhFHyz71ga1cJVdHBpYJ/i0JCv7hNwdwWi
aKCH1qjMTPMi6NyDv+Scb7hkAWNlR/+80cf8pQi15D51KwtCwup2Cd6Wv5uca2FrYPk1vIcnJRDJ
nLmfhuJnUTwqezPYrDy4NhaSQ9FS4UjheE6jeu6jqLTFC06pBaP7p30rnulJsvatMw8m4/1cfrej
1hM3rUKjJFDbA+RUXKcvfUnSk5j9O19QB8IGgLHfo3uuWN9VeGGRZrBJKFbGVdMUWO4XHM8jlcbS
zSbuXV2aYvlEf9F036VUtA9nCO7tMIQt1v6TLEbRYWJZWNS2J/M7SAth+3LmXBuYOGk5/7+943Xc
Z/EfQjWi0JVqboKr46dtJlp5pgw3fBIIYXcz2ijm0o0t11hM6Gl4EyM5JZld2Nt3ldgCGvdPfSGV
49QUaugg+9YpSR+r03QTnfH+KWDBFEswVI1tddvZe8QlpVXG+QcyB8FyqT6L75HIoceo5NFtnAZj
Mc4fifvdvsXjVjzzOBtZ6Ce+W/lgDxtCe9xk+G7VL+IECkO+QupVpDepwMi3KklP4zEY2he2Wtw1
ARL2UkcWwyA4+LAt8b4u6GpaOMUWQr9OrAo1GSSLUId/gXSkmHXTq0sY1E387czcBOdE7PrC7YH9
dbeFjxFPwb2yUhhpm+rG9yZWer3eSojk9ygxu9SgU4bialWYHYLclBC0HPx6+GrBrElon53tjXN8
+/zXPzp0kk+OtPKMEXg8AbuDdwAekqaYGKaejtrQmSjKSQW38PS/frAFKybQlx/+Y9hTIcezRyCX
S3eTNL9EN/2DhlpOh1/x1PV4enCwo9kc3pDrqV35NmeBLaKCTl74WVusIu3QybbvLcflkALrv5Vn
lUIaN0GbwSsuVKh0oaFj7rtPhWHcv+CJr+EnmX1YOG/fwAojfticZfSxjqYkmQ5Oa+6mwtyMnsZW
2gQZVTVTpnDE+PBYw897rBxPEqAuISBjsnEon0atB+hh7VmRjXZ0oia+g8GQLHHYniyC91IC2wE4
NnZFqETidIsuM/y7bLiVQ9PDeh98KF8lai2sKVhDjWZRGuiueYayaTOFyw6zAmc0V13mVgjSlBJP
dstkE8Fb1pHqn2ujf9LZrJX24yLLhGcXQQseVYc3zRYobSrUu3hXGAUV7Cz6OiiWLG8dYevQV1lS
iVVzdbYsSI4dUlyG+DWzn442ugizVsUPcZzxuYQTW8JvMXlvszUBJj8+97XNU7JqtNEz5aXvZgn1
ht95UbmUO28Ldw5VRxFd7dgk/1AX14H8WSSfkwpSNS7v5P5YX28h3rz41wVrkh9PoJ6KXW0iaDjm
xtUA+R50xLba5W51YDb7WOEyl1KcchJxMro5vyYhJILIe/C87QC/HxhX9TINFdbOdF90TkWzPxSD
u8XrdVA3nBeFM7HkVR1qIZjuO/f1QGH9kc1n9+1km+0U1VsPNTi+H4vwj4ioxw6IyXQUrzO2NaBP
ncskcDDds2UbxBrQyU0RkIyCsn6jhuL9dXUL4uPc3Du+lBc7IO/32IejdFKiqlM0bT9DDhzjcsvV
XMpu0XRRQ/4vCgnJ0TNzUOx4Rapb15FXNZA5uGsGa1JRkVIBMNBhiir62SF/FeTOEi5N6+4MTrst
GX+cC5KaQD+JJ1bTWk1Lp945nmYyl+v4vtVtDbqYy5RTopwEs5YLJpXUYyGA513vmaMJvVjovG/X
+NcC3+9uhi3MOSNuigW2n8v4rJt8TMx2glc3dqMCmGXhD3p74YX/0uY87myS3SY8+JXgohZKN0fW
hzoyTNXeKfnYALbxKVjgtscnhmCdy5hbmMOgOmUcRKwgU3yu62Yy9AZ0OsueUgJJgSETezzgfjaX
9EhUJduMfbpDXQkprcS0ZXAQIiTM/0n6iH748os9PFTYekRTXozco800xyMDfRyBaZcdDHTMWJln
61IK46j94JXK3sGblDHx821dJVKzzEIlcBUBBWBORv4Ocy5mSXUIn6ndz/QObAt638n3K6KQmY9J
DF0hZq7Q331m2Zwb24Zc4axE52b210RnAxdUBNOwzoHshRG50GS3wNdU+xWZNhxO8gIxirwpadtF
R2RlPQ7ErtgsAVkZqqf7qSYIuOIx4elcATMCFhXwhU89YwZ6y07vFuz2nV2OXYkyBIrC5/1TwBqN
6/c4z7cwM9S6AQPoqlYeMF+qxJ+X2c33cKGqa6+DFIUYLbQqAwGwyeXxfKURVxqgTQFZTOF0DIpC
jUysf0ngvLZ4QHs+FV5DRywDouT6RUX6/s1RrEhbqYFryPpyuUUoX86BLHKCgI3VKjQWwphdfGgw
GKH7EMkgE1lSJZQ8/Ec0stC1EjDd9YT6XxywxCD/kccsvrdQppsh3Vf5v+x+vfpGpHSP79gZBDxs
GrbMgq/u8ZZ/ZDDHx0o+un+nzz8NDMEFHGD5OHfI6w3IDqoKkMO0Mfd7plUl/JbcAQwCIjx+xE/a
1WkaejK6eldtZTgqfvABEad3wX28ZrpQASQfTKVk2KfWSVQQNyWa4KBCCVVWxJX9k2S+gomRRe3H
CINnJ/QqVHsUFvWJVzG+B4yJIE0qk6qtskQp5PkX+0LV5Adx1f5Y7MdW4yoiaI3Y/mKjgYh4xFQg
GcvS0SE4EqapxAh5TJfve+skXq4AAT2BLMkr+eRlDY3Tu/TIkToDoPIfRuZxmrwBOk0npGf6HOe2
KeLfSrxd3ZHO5EGPNxYIzd1gb6YQnQBaB731US+VjYAWfgAiEVjweFEwRBcRURFYSTl6nL4A6IJa
AQxuDXw5d7MEPwRpeJHdebG/o2opU+oXzni9kW42YfbuVcakrL25UtV6sTghloAkEebSClxW99ZL
szfUq4Dy3VXGvJjjC99dbJ/k1n+iDGjafLQgShx0AWoiP3TsNB+fI2E5lKovAma7OSl9ZylpRv5e
J0HRwiIc1C4w7bIpUwRd+UDtv6sDpqEwkaKu8BS5YxFtIMmLagmfrFheEA/9tJh4VTW1IUTe6OrT
1vpJLPL1rRY6V0w9vc0Kj6hiKXZBjXKeM7xlfVSVnH1M0PHMtsqhqdf6h39AI6GKjpq8lRMibzPa
4X5mua1L1lwbbhJ/TLcvtnzFKQG2CCmQyDRw+XiN3A9WG9yXjm2WkXkXprravXE9qbllJv9n+JA2
Y1nraXXWB+yJXTuJ/QN6rbhRF5b0Qs3jLh1bkriTGEX7X4Ol7rIp2Ewz0XpREtaPZDwCSXopYQKh
zY5U5cM/Tyty/SDPEON0pVOgILNdiHQ8pE4EJJZR2m9cTxNfvJMC28uCHDXeAoxIPZZRFBxxitPa
ApT0cNWp36VcMLRYJtuez7OR5nOHADqeeOcOZr195RcQc2m6O2GqtvciDHkXrgXrVGp9GCuvhyyH
twisjOlNB2PuGJiOe7ZOCX3bY1qXARM0u92aVTjthkJnCBPhpXN4zuY/8Pl7l0m/uz3PSsGJAgQU
1ztCcZlwwxmzlS3A3+vWHGcbZPYNIflUJw3CQRxjA6vt55CfBQjJASciIO9O5G1xzPGKOSh7uYAJ
hIZuuII9qsYI4lvDWcU8WS4866uDKZckUjPUBzk3Ts34+pCB7VsnLPtVDl0kW9OMBh/QdN/M1Iyk
eNewgNi+506AaQ2XICoIn58R1HVKF/ifYLgvubZQ7h+EVzKykL4GZP0wRAD6kuiAg03XunCKzguE
28h7NJ28NDbvErLr1UVFxT68UZ9H3jAIqevFdw+xBH1JJYm93OqGE8mfGxx9pTX4T26hR9UxuDEa
JihjL9Ua8l97UBZifvBbO7lCPylBckyULRPV3C1ohcmNd6Mg5KDCrDptmiUhulRIqoVYY990ShYq
EBdrmMdlLIw6TpkWXngv2mpildadVGV6m7EVZS/9TBZd8rrHNU0JRN0Sxn4MhVIuc1UgWTwEeoVK
tswY37oJbCYB7oNAR6UPVyGJPuJyCE0x8K687CAn8RtCYD4tcnbol5ru6YGx5Kb7ssV2sB2gWY3A
PGfS2NwpCaYFuZ8E+RP1BpBYXL4BelCIBJB4jaR2+PP+Mfg1TzNR99uvfY0+oVEpBzF/1t8HGdGz
bj/ttVWV85oy9a7k8C45QsLWfB5GeXVOn/1laL7LnHP9pCY+Dy58qUHpVahtSeTPuBCfwAsXhnrm
Arre7YE3X445pxAG3qCQVamVzqKXZoiJNGXVXVL+DcExoeLJxWiqf3dfXjXTegztpQJs9+wc1LL3
wEzZc8M4BpMCitNZxwtB7jXSbJp3S5RqF8vU08AZZKQ3gNQfYAgendQQ1udkJPKPk8ztHkrmL0ZO
6OcEPXlW9FrcoM9M1RIVqnOtDWp4tMroeSk2THmSTzZ7sbQDLpJPZhMMixPvM6jp4hpXOvt9elSX
bgs4c2DbUo0xkG7WJkzhCLLji4pqgBRrcuc9auevHOp5ivlGWJwNPMWNFeRtKxnZLgcgETSnvCG8
fwoTF62GwO+h1GskiJNIHNaTD8OmmZZbQMmyQ2j7wYIn6p/jlZ6Q3WCiSoMQRarvf7dyhwz1P75f
zV/BwsrqW46UOZWRFJ56XPsG8+UvCdzyWr36mosS7PpjqVAAJyu9Cf06OBRphvZuUzbTUAyZxEcR
4xqHw2Itf+n2225MIr7hOdJiyZkfVOM8f6uHWkZuRUSWrH/t9FtnZxPqgnp+KkAI9ej8Ev/Wjk3s
u3UBxX5iyadRCvq366Ehxdg1a7Sncq+xq59B4kJDV8yFGuWBfTLw04Ru8NAsCZfS60T9/EXIWihc
3jnowv1bdIZ5Ivx62T1xhk9o0kcDBYJm/PAF4vCiIs0va7fkuth5+x3YfjyFSNrrVuVrhL9QhoUL
FdfkMjebPqWPi4XnJgzgzXwzypXiw9qlfRuogvEuz4N09vXWuX58gmbC9N+tbxb2Bpgc9oy/FB4I
pL/8N95QdASL2/8ocEYuoU2vQ10/VSeYtbYqEmUkvzlm3mzDuPZZ5wIQMd9O9K4Xzho/PGMeJH/E
wJDSRbY12jWNOT9YUyHUIqDlwqvq4Wz80LUeSefN30rtdBkgUyufhUKBs+F5QjsA7Pf37wYdhuuJ
A8k0UktyU/nIooOu0q50iLOHunrCJ7s6W9su6CtpwBOXl2FPtapB9/s7WgekFW/GBxlzZ0PRxE5P
ujWPIAk2VW+ZRW6OQ+2IgHdJdmGr0eVODZLefmUf7RLfBZi7ONDHwT5lAA47JgtKyCjqvtwJ7mO6
ccLA18DI8+zP7pDL2hlJI78B8ASL21Oir4rgYrqHJe55pYX+NGFMeUbH9dGm9Q1edQ0gJwT9EX7O
CjNelrJ16FZ+me0DSxAa0kmHrhPXiSdIM4lA5Bh6jLDDwL6kw6KYDnwg8HXX2y5Z2AKrBgk9SQYs
LhSdLt6EMc1jcjHkTK3pPAZYr5cUCdOCbl06Uf3vM45mc4jKTwFoc2XauVUzxeMKyjPG19TpCuFx
L5XkFvOR06J15FkKn9cW2b5u3q7EXHoaY1vnGncyJ9hpa1hygJQJc/vOzo5keLbPfZE6npxxLPpU
lIu/qCVOgqciJqh+7TPkxONe1rXPAFwWipUbnsKNKtQGmrWc9Emr2RH/OFiauyMkamV/g5LzXSYD
1JyzcBdG5NAJ4dyZB0KvTvYzrPpnvnU6Om/5bp3NG03nXOKHZUAw4tKRbyLJ+ZlTpHI+TTFCRCyQ
6XbmBoO4wyKIchNHULDgjVIBRrDLdHDNoEe8cmraaz4iGMOVhW7YXhtPC0bKzl0RmntWznN28Kcu
eBSoWxzOWoKgQKYnF2gdZPEMB++WrUvWCu6/F+k4uAMUSjBp5e5ddeZPKkr7ovrRZrLyW3vNpwqN
tjXnhoIjIlFy0G+LqJfuk+ka3YpQU00MAuKDHzHgVzp1I7Iond64v/tQHKShtdkPBeaMuYlrWX8t
i1soZLDjSziCgfhggUMbJfGApVW9MBGKpJWdpo51jOBbCV01gK/RYRP1OImtT55T5yR1cFn50HQl
M/Z3T9iu9B/2+7rSruSztjA5qoaBsqCFHlp4wtWTQeJDRlWSHmsIlMA7SeXY75UqL5XCQwNtnJN+
RPXBuyQa7ham80KWbEGeMfsO5OCgDGhQhc0ruubXpBc+KMfHeAhsmamknssKOoki55gaFfKxDBBP
Jb8O5Et0Z84tWh50Mi23G1UNZ631yrcroWmOQ9qrH3hHqdAwl/2oduMh/JMWy7Bi1Iu35l9HVDgD
Qqy4Gb9beJZeXGXhhp9iPABwvrEwYw+CxHTPRy9pzGfGrAhazfZejG1MVDaNAPlcFZ6PmCJzJQ0l
1Difjsa3SBSXcBb4QPvYlPyNISh6bRuXtoc4CS8NVyek970OtUJSBqPBT4gjxnAs3e4WrV6wFyIj
1NyLoA8fFUx+8uNcG5/BRh31F6ra9QTUavPAwrKcq/pCyfHTgw03LWMfS8/ipB5uSQNiZsFwI9T3
hLAml7+YIOPHlyVRWfKDoMYxqlpgEfPsMDqa2ZK7I0+rV05uxJsy1MDGPQkOx3U+7dfIXM/iwwXp
nhmtN2GJMxppq4gN5guCjo2R7AL4Wnx/9q5uyVmCKFqiDeEqD6jEIjx3uOc7hdvhHZAdZgCODKEt
n4Lt4tjJK4gn+x6BVwCRGUW1pY+rHKNOYKLwGUQ6g14c7Rd8jPHpYlN4BtwuObbjwI0UbxMUMfja
giV5rKof3zDnbr9IYiICKmPlHB8ZB77R189IejICME81YcGgYTc6XjdpV1LhiZaxzVe+cfa7pqa6
SMLOqECcpUb3zm+zCx30xEc1FS/aeEq9USBo2bKJyDAvM7yi1iuO8pASClReA8AtS6eidTLMP7+5
uf15gl1txAOQVWm7ShH5InOh4DaMdLu/K6Cvo1hpmGc4ZJ9lJI7xew0TEip96K787Yipz2FInYii
jQL4zTae9EioLGssnW+c/E+yvdppxQzGV1EQLeO4Pow9wcV4PvJewKk/Eg6G7qOvtoxA2g/IrkJ6
2fRj0yfuNksx8pOfv9f/ey8KH7wTJ2lQRRcMncLg1NFZVuXUU+K/JN1jNpkDkGirIPFKmaVAdxs3
7mAL8JNIcqId117+6+s3zu60MnKZUNPwYi2v/JrTCQ852pJngS2XkDk2UjZwXBEbPMM+ZQq6D9l0
U07+lH3moSSWvEYNMu/bGmCw+Cy8xcp9X594jmyPXvCIYhmF1QOPcuQrvno4yqnCkd8SybJIH6gp
CvtXL7nakbkkVME0wi7vEUA+cfK67c3rJ3SU6VZ8usNmf96OIc1V+UL1QxBkUyIMr1COff/6LSp5
rElLrkTEj5uMI2NvTqq7DpYii0ckuZTs3ug6xkXhakUbWIIL7xdhloZWcLji4V2kOxbY3ZdAT+jv
0WxlozmK6KESOIkQICMqrLJwlGVRw8O/VyXLb5o6etGThV0twRRSBUlOOg9eM37VtOzQqEgkL/9s
eu8rJ2mJoS/PdotT7blsSocXnjGW+ESiwb+i1FMwJnRpE6Re0Hh5nKw6a9iAUjyo68Oe70mSv5PY
mEpAFotDObSIBDymyCNBww5phY5cSNZmdRS0kZwL4o5Y640nKDiKpuELfqLFaRJZNUwY6ZUODZtL
9t3ALo+xKfen3HGqhEhrzIAOAr8my0xPDe5O7GaOMCkEkjhbi4GoHSnT7vXLLik5LrCqSFOgLyaD
HK3opVVGEJf0RrfP7F65yzO8JliGun9m0ymzI2IMd1A6PCfDP5MH++egrtddhuPgqIukzr2EqcK4
OOP+u08zcuq5F09NOXhSCA3F6wQYinp8ojOFD6sVIl909SmbLQAoy8XBqY8FE8WXTpsR70mLy8e5
Pmpcl1mhv6jjRtqfC86Me//sr0zorDyyVKzztXMKHHhmt3Hm8O3nZ4DvpTYGDqI7p23FfVtiu2Yb
tsOtlsVlI50Aw5kRTLuULV6yJQsMwFzwLRfHB9DrpuuULOCChbd2aeCkQ1I3MWr62nBSJQ1uY1nG
y/uXjopDEA8hMupGnbtJZQBOET9vmAv20jXkzZX9chdfQhz/25GoPBpZ9rYRQFjoTRELgkxZK9sv
Bn612nhYk6i6R7RyBZuafYkb8ewm98T3a3rKkWZXKFqqNircB2fMyv3tvI70ArerVi3lKLZFkD21
LIlS4bKp6rXCM4u5a/nQh3mx/GZWwXFgWn3bgrmVbyDZSIvtz6SLB6BIupF3ByFOZEmvWENZgucD
Vll/Ac96l02jWnzcFbHqI+Ykj+DLPLKbebtw7WDAijMKeBim2uDs6J6yXlH/lY+CUXTfC2ZrksPd
K5Xx4XwRPRAUTto9VEAF3oMgc9kHE9yYvTR+0n83+9UXVkwoDiopMvDRAUrvD8T6hYlmcRiebetD
I88GgUReSOW4ncTC2MS1rhqr6fLRZXVrbNGC2VtrgK1TwUsBkJ+w5eW3FBC+2nCPsdgtk6cR9oVW
97BuQDCJM68wiKge5oaghn+iiU23TUupzFk9elulw/qcGro9iI7mS+fBbqcTLsrPjjNY3zE7dQH2
mZdXGxUPxaTI9X1Cq9CB2HTiAmjn3rWrXoC5l+8rATYEcizi3OSPrRKJW5UoUIy2CPRAGmap09sU
Q18pghgk0E/RWBw13v/DNPrLbkfiCiMZgyZXaHUrN2+a6U3ToCDpBEEYcooeXwHICK7doRuIrt2i
aan3jZ9UMvmcqz+H1rFsj5lclHRNfLWj7XonMNSPw3mp/v6egRtuu0oGKP6mbKSDLnXyvbj+ZwUa
VzwbBjK8KWeGzClruRy7MNrEAY9KVXx1VlU5oxB2EFKfoiOK3v0za/ya+MeBc4ZEqdtIlPh+7hsM
8y6rosmXIw0z3BArNLeO5N1859ZkgIe/Y7txJe2NU4sWD+KRHvHutbmk/gXC4bdLsNyKPpNDrj0r
Rk978kz9MDwszOUqfbtPAacOCRfm1WpQ+Ss9PV1iU8QnYNSL5gmzTwwHKfCv9Xa1YJ+CuFQuKZTc
Q8uIyUUdg0fwUD+cQTm0vBLIiw2/Cpj66uvqjPhU/T0wcFxPKBiA5wHOxjMdoymJ9F/TOORsDhi5
jhAgTdoY1IoZ9rjldeuibPYzrj5YbPhyLKTEbsv2hrA06IpcIV8aq3xKYZvJLa8y8o9wdjknyFhD
CAOX6MIWa5kQ2FzpJqwGVGxQNHsiLYFbX0SuB0fz0QxlKWSlLo5DeMytUwL6rq/XPTBooAO59//y
bUR8HHRoMCaX5TbzIc3TPyF72nd0SPw217JSY6eSY3NzbGH+M23BKOnEAcho080ay6O7TEayPUBc
pmqWrwM/0a7wkm66cRDcCq/y/nGvnEORvP5ztzThGdsDXdxbw1+kN8IVspZLqezpOjp6FGa3KCEe
AbgMC9E88tCAZXH+DxnkJq+yztWTSX+qmT7z8LJXxjxmbJvWdk9qvt6wb3hqh0DUsqnf0Uif/Vvh
5UXy6/tnzuKPNAY+pJhopkEdrU/qWTp9+c/6T7DyIFjRqnHUnpmZDki6e8MI3N7Xe4jVWwAgFD7n
1szK0dbmPRX8lhBL1uMuUpSyhE8gd/ArxSmCQyZnmy9Kc6fOO17vaTQjxG6J02Gl10lm4NXB0Ovj
sPxfdJVslwJzOBcykZeT2TUvoyBNTD1NtLpA+A5lVhDMJFjOuJzXjZLgZiQuDmPd5tg8yGiBFDr1
sKjtR4BnyjQVBTXpUtLim6ktVFxU2A7Ot+8Pz/jAhm+E0aU6UkH/6QBcKWT75EooN1s9OKnfwW87
sm96Pkq9k3iDZYBgKu3AqqTdi/8/AlEsiCu/KjiBcZxMS0G7taoX8uGBIluIwJzD2C/jgoxaxCB4
c3lr+HhptFTjZtFzo8vee+MOvbsFD2a6LVvBARzN1387eGli2e0AWubu1S1/3C6dJp4cgk4G2npj
83HVTrFJvGrb2iMWaK4bTXqqPMJGXjIG9BFRio2JGzPnfYBTAkE2QtDf7WfhCEQIuIiCx7O9PPX0
Qulpowkg1y32CrMWm+XDn/NevGB2NNini7AhBRy0YbxDcM7KPsTFcERU/NIzOhFCm8LWg06Q6kuh
sLJ5AhNHDTbQldLC+Vq3lcwvjHth/uzN6QK+mKjqZ3p+W3nzvb1/+7wpGtIoYUOtNJeW7sywpky4
qt1X4DgeMUW/vi11kLLrAtrULRFXvpmk0bO16uc1FoQzd07/HahSvGi9c6iew+PlG/Dd8Vgwgms4
D/wt22lMgufCpMIgZ1iWWIUybLEH/PW/Z0uDPpLThLhF7IaJqKBTvIU1b/ZTsRMoYpNkQDF5SM+Q
3osnEqYWgizIj2DmZWda0zEIRCy4h97X3PkHItXm+HkpOweC8qDDGoQMc9GoThAmQQPW/EJu7LcD
aBR5KWFJdNi8iqA4gE4pGvls4vq6F/OCoGVbaOhgiUk1hPsMjpV0EU7SaFhhx358LJd+ELMqNLhb
xEmPX2HOGSsAJp12yd8YzNZBQM2gvgm2mGrfQyU0oqqEqDTjowwC/hCGFZVuFfS329dfLi6n1uUp
WVEPrXUHbAtWil68UPEtpL7iXbOl9jXyBfdzNJ6T5rELZAbHnlTgZ21oNg8rDDn3+6KBp8X/YrTz
VWjKz2Yg1orUKBJGoqTW7vBFIBYKlOZ9gxeZDHGFqJo+VSLzvhLeWF1Qe5mMztII1EOMXOvioDPB
E0RLaybI+KH4yDKFQiKPfMrVvn+92i0TjeJ5vzPXbpXPWRQHSwTOtwWq2vOOLU9Vr3G1N1qK8BME
PBSmKuCAtOEfMhnDo0HkEREuExWpIanRjcmv6nJHgHQr/wF9Jtkoof+CAZPUsg1NYcWRP4ygfOi3
i6fR0AeuppWCSAZWtIgQLmdmyoxtklSdY4SHYsP3gHDfG0b34ooLD8T8tVMNp9bUa4VLsFzvD+z+
lg8rXoiIzFCHiw2U/PxkpEG9/8UNdD1HjvOrsx9NTzGRAMG33SE/mo4/84hmz0s9yHlvpQdPApb5
dLdwwqJ8tE/H4I0VjE6tnCVtb/OxLtCbC1Ao77uc9L3E56/Bv4mTnA==
`pragma protect end_protected
