// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YlsDDTgaPDfQSrLEKorv5lCC0kGrIIbwX3egRncU3ochzdPTeKuz43p2KFySi3heKmNnGJvlvK0/
Did/QnB2s0SYa8uJv+FBNFD/t2XMA+rpZUK6jzJLQPrfe/Wr2xEkWdCVnpTRVCZwIJFMU44AF5En
UEpw/LEf6z2xQ6JmiKQcfWPSKcgLgo28fyy0MtaPqyjXIUHmqplHKQYGBFMIZ37x6VfS1tOORuHQ
D3MlYiwZqqKUNU4wqnPaxxqjKWgrP7yQTXoA8jVVjMJP15/XVDaaofODN5N1ZJakvqA0f9wZmK2z
uOQaOT422CYOSp0dMaUyLHwfJtbeDi7Z4zroNw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
JU47139peXd7y3TGeeOb45MkzMXL2y7yTbgDQ8JSJ2YKJTOE9h7QgPgf7ATh/DEts/H3eawgnaOQ
LbyqrENNPRmdLd5z5Nkc1GR1WzAoI6dinXiUapaii5nd6aK2gbIcg1+nR8ISCzKHHMb+BmK/r2rG
MG4CKT/t5fo09lafHnqBYB+rrMH7GiFKUTiflb5AjbRGVui6WROE/xt2XMg4kE7QuUlOgW+ydvV5
DheuXUVE2icJVgOmtHRPNNZvr/aSZY4Gckr6BLFkYw6WdZzLSEXNSoEyaQcuhmwEL4NYRtxnfX4R
unonCe034fNAWKx/z7hqMOosSAwWYaVdxDRQQge3+fJyFY6VfuOBP8PB4cRHRnqOa4Uoej9qtLu0
a8h9j1AWbrx7MR945qvMP0xgEPs6goGjx6NdMiT4a5OQp+Oh5EWUToIo4MGuKQe0MDkO8HDeO/8x
9adgT0Z6A7qT+UCLD6SuB4pXSS0PwFt24m6rBvcLpvv238ijgJqYAQ/Zv+ScTLdpG6sWSa7QPHGA
vw2Duye+JroNLgomeryMqKWvJN0NFfRIsjA07tppYaMUsQVTVbTVHT+//d1VMsa4vpqwgHg26KJJ
Vb4T8zX7THLnPFon7doPo6PvVgC9hAjyVjByvoxvleprAEV/0N+GYMx8Savb5SbrXKzxHdxLwFRW
lLeTIYQKWbeykfcInrkIECpGrCsdTDZXcok9ijLIR41HVPN8hb7SpvRZZDARvmSlpY3INqo7VXgh
wgyrQA6h5nexrFr4kGG3Fc+LDgQtq1trLlhYb1CXyyEho8DQQ4OCVPvntXJhotOQOQRfGqFA3D9S
7Z1YvRhetSojfobhuvWj5bw1zT05fQ31h9B1NgCnCIEnVnxzuzR3+TEw43x0k4jUePGwU7kHaJng
TOmEGi7EjN+3Y2VBtNqVKWna1Sur5y5cp1etlxGckm6zgrlnqECHH5egmrL9v+/kv0XFWkoalERf
eLQUqAWRIHPJH3uxRayNsAvWBTGt8JmkmWtNGVCpuBhn9tHhmoRFbVi8Cx9TcFD/hQF0r2h/8eAP
pie0wnJ/w4UX47DCqgRmT+RshH6ngZpolCpQhSf+FV3G/GPPFYQ/HLJ6PakNVnGRcUHz2SOcX82b
8gI4IQb6wW3OuPywY0fyKI3g6fB1PlXra3k4/JVojA9tDF+AKLz5VMuFBSjkZDwaQbdi+xXRuEkP
Jz1VwkxrpBahdhGTKw7lC1bR8LnOz3zqWZoYUXboZlNlKXjNX1JoUbLijegMof9x5oF66lVljnbk
jVjwHHwJwQe511WytXS5a06CB4pNbZobyfCzO6bVafWdRUQvbExCVkBJkdHxe1yNzBJl3ncDl8qn
DvmD6lnTA+alkpPLyNG3lShoWfPoAxDEyUbNPGPTtHvSNfrwXu42W/gW89h/cOG5T0jxTYdV8oAB
cRrYY/0b3dLq0V1Qeq13q4BCRhJQRBYY+O+HXuW9nC7rCSkm7dPasEeNxc1SnGwwIQuvhjCHfJ0J
NByDqQpxty4UKc1nhW5xjVB9kEj8loGrqDuQIJFAok2+pMPkA77Fu1qukN0YPZ0wMHxhTxiNqCLN
V/KefXnU/re0OObZE+xbqrViUufdv/kQDvo5CjH8PPBgHODWVtjq1KJ2RTh/99lWtIBR/rkEHAxx
X17qMbpUVYnRIG5t9505wZrA3UZ9fRAgwP770taH+gy2MSsGH7YrfX0gyYopIVllDZ0/+etkYEaX
aEVQ+6VF3uR546ryGNywwlvbD3sBxANWVjGL92bi/+8e1PW+PfTI6HBXchpk0thofoAnM7ew0t8y
0HCBLZQzSEtD6CPbsG0eGmS/Do9cbbId/Xx4KcqQmC40s1a0jRjDQfJX7MXGzv4KD3aIXf89dAAx
cpH3iySbr6Q4ycO8/BEmb/yfQmKLFRdi7+uSUdwW+Lf0eEbEnRALlsLW9taR49XTkU3ZtvZq8hJ6
ACE8YkwL2MkqcsYNcOdXE6vb4vMcuxYvMvNFSI8jqoE/uOzDUzCp7KDzrVvTJy9vyOW8mp8Bbs8Y
6GnwYRsS9V+7LDV+2vHkJU3hDiOBpJJJpCWGIrN/IWyWlpxPMjawtHV/nLdTiSQYP6pvanrTvWyw
zr+aC2CgsGTBSMZWpZg0nGLXPw/jJc0I/oBegrNBqcAsTLsnVhcUxCwOgBJBuQSZeRDTNo1qya7A
LBHnGSuA2cJ2fnKgFdVIod/AZ3EyTjtfwgKz+/2BPraCF7R7xjyMWGGVxnjaIkC4rA2VFc4V8fMk
XDO3Hzg+8kqHHnY9TxmCdQ0zlZNKRViHhpH7bvhrNreyRN2/TIpD0k1E/3qQivOHbb4Ww/wHfrsu
eSVdB/aZHMbQQLmmxeQbkRKoj+TZO0EMLr4vzrJI63tUHy6h9OIRk0elGcW94ACh5iWPYDELcgrz
ormo4eRI0jx+Ac2lmMIJv7XSvtn1BMr4yjURiJ93bSfIHPYgmXfLhSba0AO83XcjwzUV8imEec0f
mVBk337pL+vRKBSfE54MkLNKpzLFN/q8O1fLzXtlAFUECobVV9qL5mp3VsSOeEYuOaG6f8xgPAYK
peCJWyr1iMR483eOitGldTp2QHWPV3/EZ9yjRquCqvu7CfGjXVO4pUQ2Hr54Cfnlq+OOXBqv5vG2
AxyxW9bY4mXuQF4Uj85RGNIYhzBI5wFRg+6dqC8vJ/rKCHMjJeDfPlAeTDqxj3l3+qVdLPq4pHNR
amIdqtoLAraLqZDNAxd5vWaufD31vtekumO8orSrVorbROmmwxhuVD8TzAkP8gGOfdLDEc8U2iuj
vY4pyITL+ZC8DeFKmINe0awVcE47dwZ3x8hNbGJu8GxBKDVjHmfffIAVC3AF37m08N0GZqvZ38vP
I7h6OZLIKOkU0RLtAUMz+0heF3vQcUxdz8BYrbypU4i33XNT5F56UPbB1tULKDJuWLcAUY85cX8v
PRhwYncz9B135HJmyRH6SFksCHfKOahJTEBIdyScFo0pCFl9MhIBXejjmJ8iK/3m58EkI7+8+iyp
UhMh+bVyWGJPXtUMd8Vz0m70GvPWoP1h0UtrP4Rg3hAC9z8DSRwaFd8v+BlNscj93sK+w/N3ntZ8
5vuqhWz+H1KGbNWXQy2QG2WXNm3qaH5/oeMFgFk+JqDpjG+Up4C1udRu28HdIxtnbGolLteGufNH
tMrgxC3E1clQy8umaV5+wWjMu6hjkowMp7omlZrryj+zJcltq/2E/+c57DU+sOTtkO1pDbN9iuvj
xsE/IptKM2SuGzhLiN6eatFbZqF4Zg7vwHohFa2KvO/mxn/dOv1CS5v7MNXAR/RhmaNqg240SEeG
GtDeplaokViMIF+1G8IUtWPBwx6eCjVV/au6JC76PBJnk5+zJ1a3hW+u8wgLJyoELhA5lTshiyZL
tcl11lnHoEa9TCmzFwIOG1CuFcqB16Nx7X0x/t6ulQGxRwat3Xgj7aGp5dcitjfi+NT6ZSh7Tj5l
kfOaNj66nO+inRn5mdkOE1/JIbpsCciG0oAFcJNIjsUL2WjMJ5SrXk7PW0+fyaCKsN8evMm9L1cC
qtO1vUFOQEdQHRBjYkhIQ+B4Pt7T+SgGUsdR1IbLC4t06sMulAXa3Z3fbp9W2tbNi1lpI3HcXmAd
PqgFB/QDD2V/h9FR0l893s9OQQxyK+opbd1UwoQ2xxGK7pSlVT1lw9HiP8X/dc1BVnqSV4L5nWW4
016siu3zATL4Qjr0OvfBa0i/VpAQTDEaMS/eUCxYi8o0q9Fi5R9qAInprlBlJeKj6ogVKT5SWjJO
NOrQBaDnnLYeNGWRixlL8mMkBL9rABcCjm/6DXeOSgWanIJj+jmV/4YygCJuGZfPKK7vkNggGEFE
kVijxI5V3cU30yBTcWuP6nCgqFGqsgT6tLLF1MQDnHvsN5cWv+FkXbO+nhSHOHJE9pLO9m6HkKEe
xYaAtZLjvQx4bJerFGatTFPash87qxMgOL8I0SBoamgplqSMBTsRiWEUYaVfnHl4I/DsoxCJFVnM
zFfM5wdTZDJM/O2jx9YInkkUgL9zr8FAiI0tES6NIRHWnzKk1FhL503lxfhpzFHrzv1695QDab1J
5w1afgXbbDSy2rJt1uVrBZ/vH97mVMIjhQvCDv54Y7/WrTBoktC4tvf7kxZWPaX0BoyXSSZMgdoI
DRg9PGVMrPeOa1/61ZL3M0gy63Ng8nG/qqdsDTxlf+RuJiDR5KmLHFRdyPBO+h2TmafL4+NYRwUs
4gbTvvRmgVq2gm+0xm4EA8MDdhXmr3zUSLXoS17X1Xzw411goSEorUgSajUwVilVmoRBofrTV22b
ynXUY/bnbKW34m4fvmdIlvXozjI4q+BA+VvAwlQ3qeSqa5al/k8er+JspotJvxbP41BK2OM1Zv5d
kRzQbSSjUEeuZ/+CefrEWUm5E1I7Qxp52qkz0NkXy9Yzf3lrW+kHfJCt79uCKxTOWAoJwoFkDYEz
NC9zrcGZrtTa6eUa1+MIYLicXKZPH+QgjPHV9n3+JdfKez0Gfd9tJk6xqaNb5Ph/d/uT3GhBhZEy
HYfw+VIxtgor4ibPDKO8gc5kBSoUSsYNn++dY+w9ND37SEx7BZlMKsx/U3cmNe59PQr5a+7qT9lZ
/mdDjf0tYB+85dcUdEU/8FGeQB/5nTvDiq2FNxy+By76Ju1Q44+amuGyrrvcWS3BUgrk+AeY3FG+
Zpbl+747X9HoRVGuyUJDMcWflKVodeNhgmhn0UAei3UOz1fjYmy3MZDp2AvDkGO4hiH8kG1CHBKs
8FSNCtVfUvYAVxmeQfqNm4E5pkkjEgMqcFyy6Lb1bJvCA5BgaruIHrO40S7oz1atAhjGqh1Yhyw8
QHHXxgXat0ZWyacM9IYnD9J+9VFTjM+B127xyKRjH7oFxLqNXqJOwDX+3iFYoWivP6s2H+nYqgT8
UBU6FRbfQSbAt4KV5pJkHcKpzEAZDH3eCQQ8bobYwMUA+EpsTJGfuFklpdNl2cJAE6BZDuw3SaX7
Li0kUXmnQ5gvB4qRkRJ2zRgXqJtlIrzbQ6au/1HDnDZDYsOK+sTPpHVsg5ChPiJKSMOQSjvrvqqX
bAJVO+iibB/bDgnUY9tzHEzzRlZXiu98tpjvaq+1+S15db6OGK8KEMY8rT9IcC9A4xY2hafNq45y
1yeK5hwWSDBUWmhWj0ch5RUAsaMgpdxod6ifE8wrdD0f7izIBakug8ZrSB00YpbsKZq7QzdaUDci
PU4uGgutWGECUjGT++wHHsTLwiOCieFVgUOY2RO/Wp3lhY0Ufvm0vlwvggh/Mm3Zp+5vGEGWgLBS
ouT5wCV8UkT8ZIw6KNA8LTByxvW7/FzyhWmgEnCLgeE8y+SJ7GHwB0iYbRckcrvW94Otdn4uTmbN
kqHr/s0lHDGnZAp9Mva7cLYQyLRHF+5CTp2lkQdsnu7XqM7IB0/9WPg0iKWb6Dg6IYlScjo/dAt+
OdS1iebbWzbwlyecmS1KYdnUu44DzK5BhICDaTGgaHY+I25TZs7jKqZ9S2X5ODhN9B02LlmFTkkf
UUWLmV717q2PhtI/dA3PmW7mJcWw35OhZSwvCl8Ius++Tp0saWMYT4g+GYGjyuIiLCVBKL+RxlW3
+LMyLo30ZMSIptFnajGM5FTmfkKAZZ01nNvi5I7kdHaHmyRuQIcbhYWZdADdkDE6pr8GclbuF075
L5LQucOCc885LTp2S7QapCiaoLaOQ5CpMF7EunPsqAS1iNk96h4OWkhtlcLLXnkfuQnii4D+yoOI
jsGVoIHd9Hgwy2joXKgc55WNWMSeNMvt1Vz+vGeQBJJdOm+7jyWi7ew+44klHUIpXhKs2a5liSjh
aWWcqGPnZGbG8r1l39BM85vQJWDcKfyDCggupmG8iU2oQQ9afYkHYreLl3oubER55OvN0RA4fFRH
vFEIOkLaP3u0MKhjlb9sJcZf2goz7DR7l6mELvz7M5C6PtcxXyfS11sTVt9yP9/go4jjDS6dfW0u
B3oELYAmxZSTvk+lgz6jxXTyEmNDeVE4/TmQEcfxpmMPHpCkxX3bUBqF3JohHNSk+sc9X9NQwaV+
uRMWd91GwE786+mk++ek/BvYhkRQbZDLQku8xxKxxZcbcGGEYAkOaZXv1hyRhuXpUx/rOQWG2kGo
GCB8G6Ev4Inewgo4LMpwb0YSGqgNSUjdDPmN9vsZ/oqzGMkNh010YlYC8SwgToQy+P80PgMWgIlq
bAFdewy4jFTbgpjiIc19TvFjorT3IxDL8F1IR8FgdBGAQELK+QMbSGl0EKeDXDDMZBvn7Y2wW4hQ
ZkL3wv0Uvvb7+/cqsJpBHXj8qeTeoRQ+/7u5zdHngkXvZLlxctZq2uinSExQ86TaZtlK0208J1oA
tFrdEQduyDicn0cNXamZ1DqWLBiHZEG1OWYqFhoVuLdBgpaW3aMNfzCqfDv2GFBPmffofCPFEfTA
h1Tzb95ZUNPROdQkyB7EXoqvescb8DE0xfCNRGScKkyBdNEjnmLzHYFY+wOGbSnUFXFBmfgJYYKZ
Mr+U/LLfG7tbcMcI5OW+Icv19AbZF7m8+jQIznCvRyAfuUUBTPKfrPWjUNQRtZe/AwI/sOp8HseX
9uZzDII42h/BpDyvFVROVVMmX3x71DVxJ730gN2D73WifWyrNFHLzcCRf4rPyI7fZJMWGRmCcEy2
1glZKmqP76QE2G+US7X/iIM4FQHKYUvS9HYJdSg5eftvKWwI01mbRX1Tu5X64nRU10FJSVll1jbl
bSxtPJgUCyMd+G2oSO0pPM1exBHDM907tRqzGU18CZcVoqv+iVavUwmrO7sb3kX10OUb0DKnH2k5
nargy2a3gzct99mZN9O/eSdt4uSO0VlDkdRZETRv6oX7YT0xGQOBFqlHpfaLehL9E/xUBAt/0sOE
kjHwfJ/By17yfoY/AWmSk4ycyukJJQNNNxct0ry4Z3kO/bBqloOVfJIgqK7syN4faHSDnN5sf7Wn
71tSZ+edX+jcUVPy9tqvL8IBm1jSMXwARX1pvMZpFa9IaVKD9yZy9fNacG0iarqS3Ki72kH63cBH
uMpfgEqJ+pxljRZZFcmx76Uv7QrSI0oAolfpktXGcFdIViL8uHt0F21hcPKJAPv4cpBjAsY+aXBs
HXe60vpb0auBSOWjve+p6bNAfUFiAOK9VzwNYicc02GXGOaqWyE+E55gyGWemsI6ciMM/O9yZJHx
d2Qyd+87viObJ/ZCbTk9nMaMplmnKgK9k1S51c7+YiV0Yvf9L4/r2Df1vJIsw/zYcsTN1HVQOxYs
/XJq+l2FTldldldAN1nGlxvBcSGNUrJvtLrfpxcZHymvlrf8EVgz246VYCwAd+0R533Zi6rULVWe
lqjWbfQI5t7lXJ3fIoRqzEBPseewriISnXiGBbrk84qFXuo4PjGfrdreCju/NJ341c7m4LAoHQ1f
JH6mnoN3xHyQuRLU53pW201F8BtP6JvSAnE7CZZEAYQyb949hNnnGNTwNijR6bwogLLs+THolgB9
9pfTUHq0FoY3TpNnuJAAmbe031LDGyvKDFFwOYIGKfbW1qVp0iJyMS8vh3NdzNq3A8PFsBBKrImC
lC0r5h71vnqTweYvEH+Q8TMSIfz1r6v6jnewq2uX1jCvDuOjX+VdMTvpKQ+1Kw1OhkGaue55zitF
NOKDmd81ea5V8CqYMVW3ZSv/8JWZCwO6wpYUOrXKqeR9p9BDfspqtOH5rA7NKwy81Zn4o2rD3Tp2
VaOPDQwXrkkmgF2vbIW/wZy0cKdH98zRphT//St+H+3f4BVHLJutVSvYExZGf/6SsU98bHpvuhNQ
s1nH3YLZbnLEp5k4yJjYamVj9p4ygDh956e8PuWUDR9tIfPcnIyec1mHlge8FwPYE/d8RvSgDEeI
9+jMpxKV+saTVC3D4UKFB9XM8taINQLEZAnC0/hPrE3nclGi2CF5MUL1WT4rCGj27X3iMk+dLJ8f
ip71sYf/vcq0T2ygDVYYQOZIYNaYi/kMdcOq3ImMv52yHOxGpa76KlH3BfvmVjzgy4/DikqyYzrB
8w3BMVacqXaang/x/WWX9tjotU8D/NSckHCesmD4/chskB8REANe837APMZ8SbqKoAsPPF7zvB82
HT6EMaMit4sBnZ07Gs+CNj9/M4pqktAi1DBj683lsv2GPNt6vVgPHmTAZIRugbGv2b2snfLVMUzD
zUmRi9IRcSFfBtZBKGvWMwC7nfevHhvJF5AillQl4tOYK1VSy9KkIOLuCtGUsLyFw5N0hpDh1FLi
uEyAxogD/hUAaPbZUg2yohLrwMHsKITZAJu+Ft4B8UL5V6n+URGjB6pAnI+lzitIIgy92SJDeDgT
RJyTbzDTyw3ozGnJSu327n2jnTPQybWGAQBDs/vUKJwbUP02PLt4soSW8bZTEoMCeSckEremIHBD
WL1ktd0iv2A3hqL3xIWcqWIzSwOGgYC3j9FAbnd3LZccJ4gJKoYgFDRCiDmr3P89RKv+6e/e0OuM
vQg0W0hW2SclDKTzFMhFYWBBbneQqXyWb2o53Qh4wyrXQDfA1zEPzcxV3uQTtfeNwHZG7hnpEhqv
WH/eXgEGfbbL3aDm3rcrM8yhUyQJPwA49MStU4JbFTcP2VieYo2YnqaM/aqOzDHENLAFbqfhxxos
AhaK+WLo6zj43HHakO3HvWfzFDC8JSE0TKklA9nm0nP+/LkoB3Qa/PKEIgByd6dc9QvgvYuqFXXd
l67nnxBdF1dssl55rN5S9Gj4jSNafigTtwSHL4m7xW2RmImvL4UEzOqX0oKRg1Kjpy2RLxco956H
IQ6MgI55DOtJuXdZsbLTFsUQ6m6suRHJ07uJ0f/kiJ8jgauoFFArETOLkanDTu9xe8JEjEaIsLzS
GuwDsHEuHbY3+oABmmDKVg1U5QPjlCRNJm8szIb39wu+VBwV7XwsEe/po1EpoW2dbJ02xTZqWgpv
nLcGSjhsaaHAQrFJ2EnAL75/FBk1Nl0V/Ps1bQHPj3M3WmbcLtS4IK2BN90drXhBlDNTY5D4gTmA
aLxyPkgRPCHKV7aJfgLh27FhBrA/shsJsxBjhGIHS0eHwgmoQr2lwrcD9ddCz76cZax+uKsRHNx7
JvPpLTZ3O7lUDS8WYiMQsFEAXOY+ABCCiBRMDFhYsgXOT7a6egonEri9SvF1O5e5zWdR85oL2qce
pZHJBETV1Ek+OwTUJfWpmSVnCNc5Ua8WglA5zCix01d+zy4z1MDbU1XN5g4bpYV2NPFDQ96aPsf+
PPpCvpJKMdVDMUVdm1JDHxVLeUuXtPqmMWMaEqc5j+R82vD8F72J5aPhCcy0RGnSUzaO4TT2YgmU
bm53z23TN21Xpq3llvrP2E4xOoBavZWWRbz0UUxCjY60HGIoVEH9DhlVDa4H3bCn1b6KlR8SR7gw
Ot6+yy1hOzOpiPlkfxln/4RDh7uScdAi1CvyTsUr+xgUipWZvaaUgcwo1ItZCgKwdY1bN5apGqqQ
nYx8WJk9Yw+aHHJ+1c/CngtP9ZY1Q24PmDaF6GJqTv/CFa/sCLuBIqRMbIHHi8oIPo+rqcstXlwj
oaAxTkK/siH0Kpmx4MD4zA0lnaL3hjs8QpNNKCSkzv2zNuhC4OkCYdiafLDK3MuoCAvX2Uj+Qfrr
X4VYPi1IXV11NmoZ6g2kVexfnH7DF8CVzQ4t8VFNKjJI/W4O12yE67YSD4A1YiwD2x7ReOgMBA2n
gqpUF7O2VmTWET5sc8JV1ejKC2aGjMw0ibGTSR9J1UeK7QfM0s/Qk+bIbIWr/NoXjM2RaIXg+9A0
e775SiTQhCl/Ah8kyoHMvZI3+c8PnzHwJorZflVmf4/N8rUOsmjeOYUYVJRUOeP+wsPDZOUU2jki
tazhBsljYNsZ0AZooK/IuTV7gmpOAOndR00nW90SUUxsa6z8KctwashaVh67hAfLhCiwDRpIIKCG
aeqHf+74C3E+YptAcIpSRpfw9JloFHJ33DD4HyofZwT0IBlNBq2HpusQWDNGMio1SBI7BX3ZPTMj
xr0yG/Ixpb2tOefaPd9IKjaXDkdXHnxUO/ksjUaEbUsx0KDEH0r3E2jDqsYL4WSArvw2J3WzCMgJ
PkcmuitgBhfwe2+zqRiJ5KeByiAMFAJVpSwhjON3YSoGoWzh70cKxmOaEL522s+sFP/pXq17+lVg
PawLHT5ZJHlLNGwmqb8xpiALcXF+78Bx+y/DuJKWcygOcvvDlWYWG6rYdCvVyYFXdRd82ex0u7GD
fLXmvk/QUFYefg2+65MNwV13zJrRMu+oEKIUdskItvolzZBkDI6VeIyhEF3XLQiti96YR5zkJl9M
WsvHLqyclT6LtPZBiWy2Zw6oIpIbCTPxqz0AGw3jlCw3Ca1di3e+HVsEPyghTz9a2EevXDcVN3aD
oBbs9DHaI089U83TT2FTg2Gr4z6gPbHAgwDpxZzlFm2E0isyGUqBe6J5dHaC/zT7ikvWgeyqEH6Y
+XcjWAMSlR/wSEmwghO7qYDnsRElklbDsbMHxUJqA2sf7StYzqTN2LPwe7hJCC96XosA3/rZu3xE
LqcxWGDNL3TUYaRoDObMDq0OS7MrOdfDt70iB1yYGrPBFEETqdGIjzCgbAMxjj8JATapBWu9NBw7
ZxvBM7SFK4Y8yYqn4iNPIQvkgkbI6UtQy9tNoKG2M1RzDOGrobKchhdopdkO9IrOd6J9Dv0pWSCw
krdbw5ZUTt81tzLfDnFO3BoHTiAJdkaAVppqlcuy7oYmaCTt7SDeAXZ/4zNSAxqpFJbTdedwyAIk
JdOG89s5eMy5bHj1eNDuidOa3qaC6hQnMiiUctXrQ2hsuZWowaJXpsCC/JYhAM4gHy7PRFkR1pUu
26LgiOfAchL7dUNyO3IeArOnXy5piZmy7h4kyc7qtKP78SwGwq+KIkOejOd+mEJvEiCcbN7F6q5M
qy21qZR0LH87nMoMXcv9vTWopMTqx03aLADMh+/rlsRxpfIfZedVs1kPizJ0p6+moOWjReWY10kk
Rj1gZ/WCc2FGptHiNNmO8O9g/Her/n+qGKKVktbN06Pk0nFSw223kYFmUnWzettSikWPOTx+G2pZ
SGHnI7OjXehYapvd82EROFW+I/MnbtaFww/Luife159JMj5Xoh+uM99bHogJnq1nvcoNEuOkBjFb
OtCjEhS9N5pbSk+BlZpMpyuW7xjSZ9vamFL7vDwokfuiP5CZMRj9u/3/ynU0jMHug8we8V/saZTN
FL7Xi9cBAyEJSt5GGVOheK5WK3lzIqBJeYiweuVM1MFDq3I+4rY6ePL71yUepqtVf+ve8DlZWCp4
Lbc40mC9L4Uh56PztdJp5TcjXhnEa0nHp58ld63Ts0csKhMSjp4ysZ9fPt4zekhnHgqCpfSGf3N4
McFc8SSSCB34mbPd93VrjznlIGDcBTx9kApbtJdWxJ7ju4k4JMjZgMUTgXt2Av6CD0RQMThHxBIz
R6fSdlE4Om+tSOEWmq3DRZ5/EBIiWPsQ1YPArSfS7o6v
`pragma protect end_protected
