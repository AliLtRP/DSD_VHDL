// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oVj79CrBbjY8vUWRKLIzZic9wp4eqB82hEl7Alxt3IavdDMUcz3y/EOXso6VDcOr
3lsWriIEGH/+fEJbxMxSOSA2Bqu6GSYQp0mJ1iYI12sZoLwIU8h7teRNsBJYxDnD
3/4MRQCwRrxkI+S2aJNCL7UDsYxV41bnL2OngMpVeBQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19520)
w+I+2tE1LczPImIdAVxNBTfLnYIWDTz5I/GZUooxtDBKMGVAFCfJFRQyv5Fng+pO
61t3CQQqBEnzLSpkPvx17NxM56sH9pC9ofgTcFX5NQOGm0GXb67v4OJ2pLjkspWS
Fgk+Y3z0elBTPZaSVikceS/RpmssNL8vBzEHQCwd22Z1f6HOsnOxL80Ah8KMBqDD
KM9FiEYZNyzBEFNi4QlPwGhZx1KyhMd3YhYvScb1iKDJXYF62v+nLw79Jr+q1aq+
S+pHTaworYMpIfMnd0BunVFuKPfRmA4bnRBAyBK2mL6fgpfW80cTa1x7zFzQRwWj
8Sxfh3UcsA0IiCRCiBwl3JVG4+soq64BZfhKCZJe+nh2HgiU3RZAp+6zAzWhO3R6
he4lCB4V2YFJjVdxC+ZNUU9iGqyBAC09KcWIL1ItBNCvpvpBRAZEMSMjQLQc4hYO
8Ys9fVjEGHuJkT7teSn68niCIe9I6fWHqZFwUXEiQQgT0CzwGuVu4pLs5iT5Gchr
J31bJycXOMiDxIjChIeGMUVIxb1KbkUpRmDfGNUAGz74RDrjIWJshKdp0D2DEoob
I97wrk0PyG9nGujPb+ZJwOQyFcOf9Dy5nOjTNbzbLjX0Nx4oRZ1kUl6v9v1MUPer
PaSf4ePvOMHglBZeG55wUkW7CW0wRLg7j2YZ2okNHyRyyB3M3mHfkJ6bGrxmrdUK
W4Hkd300qtc7BOEg+D5TCIjUU9vI1f6qxHHg1WEWhefMMV009PlgA/kJqgW0j84P
PIe6YRP1Cb1mlMz2+gB8vMNVbyi9FpqooD+2isQkUApJC9UridQTcZFIA7T1TEKS
undxmPnlg8gcWFIYRuDDpBiXHnPHH5HX8/QXOv2sGjbttuixmnU3B8jqiFkfsDcT
B80qRxRx0PkWPP5q6OuiIE0/Fzbf8Ycv8gfxmvM02SyqvZ+oCvvm91QzziKyCSMH
Br/X7njgQQ4hy2/RJuErevztwixNk3i9GSelEyY1RyqDeJRNF2LLRAAzQh8rlHlv
ezPHlu/j+Dy7QYzwQ1qJUFSqi4VyxinPKNuxQP71/AcGfUeti0ZH+ApvqbYO0JX1
+WhEM98YCIHDDhZVeyByPPtw1Due+p900bH7e4tv8Ts6VDeTAW5Ij4ViN9zgsX1k
Vydhmw5dzZyim2AoqlEpcmfh2+ChQpMJE1EsonVx1UNNOAvikVj77tfz8niXrmdQ
1rNf2aJvhKLMJoo7T8Y92e8OC1Izq3GDowJkPUcRqXSS5ss49FyqIUgg9w22huKH
jurp2yRc36KTQ4q3gpRSBUU76oG7LSDtf9YaZer8hTDYf1OFjrI9TKEaQNPOv1w8
BVHTMOnpf9uwEsolaRoAQ+skqldb1UvS1yTN6G743MHYTm30tIvhGEM2ySZRlLlD
A8RlSfS7oEW/2jqvZ8O3ZmvH+kPbGMhvQxQ6Mf43Fkg57g4egssUbhHcLQ0rq/Yk
9fMm0cFJL0pAt+JymWwKOKaxt7YC6b5Dqjk3RelKVsWbN+ZZ1XtviQsF3mDcvvn6
XkDteAkLH4uQNn41mp02UCptZvWsyl6RtPZ3moMnQm1bVodMF01tZ3Mss/5ujioM
1C3BwJo/EJiHHz1NsLKoVS411Vm6YGtgYhf1XBZwGnV4xPq1vu8XerxIuRkhPgsV
qumjK5qmQjAY/olETbFAgrc4OT+0VstL0WZWK5Ds5pfb0HWiewL1V4NkUKSvud6k
4QXx8TDVE7lo94uYTkXqtmYDQytyE+xWtS/mzJ3aJrJtOYI0uDyu82eegoKL6K5j
euyzRefHgK0G8mt9OpJVn0yIFKQgjNyTeq/auvufHzZsxHfQwZYe4c262mDhdwsh
OVTVH6AOFcSPT4lr0zI9AgEVUZI65H1nFlbRu/isnTciSS+GkzP1A09L9vL4139R
iVdStiBxdmYyJsnG2rveU8jBl9D0AuURuFucXQDKDRj+qCG/2x3yGGI8EDzOlgB9
0brx04DH+o05hmfEj+/D7DpBFKoZWqUouRLY7nqR3+h2LXdTDe5ZEgmtF37K+HM/
54f2u8AxJx+Wmbz3aa7k30A1uXyfCBpUqotdh7YDF+q3AFCJ1XKu/gHIXvx1FRl7
FW4j/benEeW3NkEd/7ksbVEZFKZSvcFrtpPW2nYjcLujQ+D23UF9dh5moYaFIWs0
TKZapVDqaYXSPB5/CGFZLgikea67TVrEyRMi/jY5vihEC84DoslsjvmOVWdd0va2
+jw1It7UPJJd0piCSLEc3MLIQInxRDdwZG4jjmBspT8XQ4JNpq9e0vwTxzOOikJj
GwPeQWCqSsvqk/Mf8NfZRTMMLuTo0+npJ1cYnZ3INcdoY5g1jv5xl5nE2kdpV9kZ
foKatwjeb961poE4Eqg19At2Ajy/opD4GnZ2ZT3wmnoiA8vplVGZIkW0uoKaYcf8
moQj9YrgLDWKuJHTZZSJ9OXhUtX7FZcqBdU066N950bxe+ngMDB54c+I4LdWURp6
Yusj0CnxQpN+AcGoUU56h6griy5sbYqKAispIa4whmsyTUBD6OdPMEHguZFSiBNK
M9m88USss4n5JiJRxm4SyygqfCPlU8MV0UxHYU56mG6JRDwAcu0e0qNPj9vPcViA
SR9rN1ttz/mUoYTtWjNokXc64jp4u56rivsIlV2LXHn9RsjrBPuzed93NvqE4SiF
0e3IfQv+l8eTu7TxOk3f8QPWSbobdw8PfgWEab8D9XZJiEw+XDOnhr06lk6ncHi4
g2Ix5tojUQSdlKGWKABYUeGMhm5xplGiyDsQNpBoApp3euFGT77fA7p6800NqM5T
xKyhNKgxkihfn1dd1a5v8krCqsJZonyzbwLH9B9mxJtqvWwn/F/zj4ygJERes/Xe
ZkHt8P2ZPs73B8Eee2z05SxXjbN9fwRIKBOWuH/AorrrQBNlVLvkyxLNshThC+4j
yBEU4VeTpBiN0Gt0bK1T/ddqxE0VutwzLpaWzwtGse8BjVwKqnHkkBKUjVjBBFHK
TcjfFncItlJZFXAWLReJ1eOMcsjgML1Wjoq8xPF+sPxSE/fLqOjUYVVxfVxpRMHb
UxSLfo7F5e8bF0tk0YSkFDpFWx0sYQdBdCJCuzPLQ23aXJY8pSCzpAUs1OQwynBU
X9cVBWmTJXrdJSinW6Piyp8iG9f8nUBPtYJjpn5RPC7O1ryKbsmYqoLOeVG5kEn/
Wmexght32S/VtiiyU7WvDhUzOaNIsFTsiteBK0xyV5bPPM3IorOyCOQM2Ypizi19
PllBBDcoDsqzlCDnQ7WEL9YdhIAQKaQLb/NBp5NAB2amaOANY7kRiComqx4oXxf4
iOYkRFpS9C0fA2L7bmJSGOlvisgkegf52j3LJ4dRVlXP0cFsRiErupRIaQhfnb1O
qBUPTVbGN2mqPJArvCbXmy5Z58akZ6P5rLylG4ZB2VSY9YE5U/a/55wiMhiEslVO
0DcUwjEzWu+xR9wiXePVrYniQY0/I7M3xy2abGBBiYMmJrZ5kjr7ikr1EzD/shvM
CSEJRoQXd3Dq4UWMdoYqhY9bFEqLGJsf1c50rVLppQapnxiJcr60TVX/a0+C99Yb
k6tc/a4yccyfxqZYeROMbuS8kDn1RgR6r0RkaYaePoGRW6NvabnBdwObYyJK7a+q
hY4AzTFe8PaqskAVu5SKklHR76OfoyRe1wSh7H8LygYOPDO2eTHDNwt21EErIUSF
RDTJSFkxjG/dHU08kggS6eiKOQA6W/RnBwk47SWbQnoCe8xy43uji64AXvvvG/8f
RP6evNKtEV+amfSnO7o5dr6gtWW56joblbmvliLlyxyR/W2iP5JpHUDxFCKSESEy
Zw9sL04tsQLJiD7St5WGMHVC8ARJcIz+s6PbBmuGxF5OFxCXMMlcTVt9bBR5RlYK
YACmIFnpPxbZc98GUttBc9NFe4a4YDDXjH7zFTVwiHcfBnfEFSKo3QfUE3sVXGsw
UHZsXH2QzRK5LsURWzUR1FHl3DQ+Mu/Wx4uYvKcvk8CRfue2VS5+McgSuXLTn10P
j05tEpDfLv2dTq37H6ZdcUUpdc/I31lEQAPI0xgzAtsJZgXfU4g1ZPb5v4eM2DjH
1vCOL8jA+jR9cdvP/B7hOux5rLBjwyJ3fU7seycJVdfao+2bnaJURL7/UKPZ2XUo
dTKH457+IiQKOsLAdEy3LVVGGR4yQzbfFB6LCbRrbIUeLsqk8SXvh3C9fuDLTO6U
iwv2G5qS8NJo6Ge9wdaYRPZcI4qAn5HigPpzsuoTEwtje3yR1EdfDz03s7VY21Sl
dI8cPR0ezPUB04cH7yD46JqND5L8BOatQYStujvH169AoKrvgfbYKgcoRVm0yGne
kLZrBC6FrMi30QsIZAuHr3jboSaZaRHm1ZBLsXJGaKjg7qoZGTCJ/g45io8ePbEw
SpjZBRb1PQOpeTLte7jN2pDbtsn33DpZDIpX7f7sL8oWTBf0SOzU/JXMw+q7QFqd
2HZUOWhGhN50T+ucQbf+k/T+GIpdioLMQ5zfFkgAE4p7Rz2qbmGh11J1wO4kL12B
D/qQww//iywCekgE1cNcjNNJnuY+1WKSsPbGDD4l2NjmV5u2oC8SE69q6Ts//vJv
6eh7tYJAg8kJmga9DcyaNqITGYCK53aS6QjNcc965nbreI++QeAjWyCb+VpP+blD
M6xSJj6MNCf9cvrpIqYrIDJGECi4ZR71Rq9xW0fTBUjKAEcf0wCflf91UjIxX052
Ck16zuGLGRs+OBt6RCK511RNxW6egrzlBc4xSBWvLcJb0MELo7tIlO/5n4DK78WM
lYXDdZw9s6Hpn+E12+CeD/Y/kjwYioOMNnK2Ty3ZrVjN71onmy6vqCHhle69fe9r
4gWazDaJ0DntHIikVBM4upAZByxSCUmJ+MrS0XO7IH4XzoomAeNDwhbCFzpKRgaX
EUseWGhhnYfmqUPbD7QQKAcTk/2/iu6s7Z3CH0wqiEhcPaI0nDk67u+OW04QD+O1
P4rUGdgfGVafaepQjJq5WuG8X2Pg77fDB3HKv+v5SexMzexVrIK2dDO4HfRIG0LL
kad2llES5UCEBEJ3n2CJYR0NxnK/8jHMYda/I4lHPYlmEwAvzuPeeuAjU6536muC
ikRZ62/tNCIQ4xfM1WC9s26s8qEOXOE0VYzDYdnOO+p/BdxacBpjSUT/wmojH53z
2Z7WsK0u9jPx5IecVYa6HTTxMu5fbVa3kM96chhcfgl9MgNO4ZZrf029n1ksA1zC
sbtE9anXbjnkxWRStFC4MoM0wgEp4fbeuWeOXMHgZlGTWr2NoG5SQCO7KPUFEhLc
vRAkYQvtjOPmG/W9IZ2IzDnrFXUmBbwk7THQ1ZV73DU9bRGjfP880Ev2OIa2VBYP
Md4YJLO1QAr7EUMRrWo+nc6Z5r0QtSeb7wCD46KElHFoc3rV9VxNcU5UZJ0GYKy8
mRE9DoqYwO6bA76mMtw9xqx3thNnRqbLjzeMVK8wSgbu2eVyrCfeEQpywebOQ3Oz
TbvzuWhOHlCWjEjNVJpGGfobJ13x5buoCdqwvvuBKBIq7CQJqjYiKa7+Wtu76/GL
2QfE9AyVXHg+2weHhAuovcJPgaKCv6zo4ILRY3pjbDG7KeDWLx/xpR29JiONXcI6
mWYJ7OuE7erBONx3Anf3xTod4DolPqEFAZ6mZHUF9zUW8lIJScJCKiCp5K4cKFnq
OoNMs+jCege9nprqDInMqFJBqSuls5k9T7SNOYQnhPh15gWWXmkZeUjHjytQkpp0
rhtSz4Eh2zshM7XA1uKZO3gB4/sPVqN8t5L6nq0Bu4BzLX6ZnKDiwpcobb/Rp23W
dbjebBUlVUJVN7Vtwl1EArW33R6Zl7co6AS/nMyc7A9pBllN7riYskzqg38cZ+E/
RRhVWwEnOpUi4Ye8pslbDAvzj9PdKV0WmpQ3YiZFRpX2o6ZU3CUMX64kkUNZDjTl
123IPSuzuBqtdIEvdq9LQ4OVhX86IXgsiMz0gTRNadk3QWizPpLrf/M2AH6J1Q11
gYHCmBGtP3xyWg1bsHLBHiHedRkIrvOdDkRMIUwt75+hGMw6rEA1N1PqJw8Fjm/5
8hYKzjwrsjwd9aUqVoURKJg6+pEAd75rifnXhKxbtguRSN0n8gXYdCrqqNgqcRvs
VEUm5Y357Q3Fewt2t3xmriapEmO5WiYmFqiUr3cOzKKL+/+AW/tdub4SqGidrq6q
enGqev3F1fUw0P2/C9i7/X8aqgzAQdnEVOv1zn1ljhPMxFmxqgDEvcJiOh4Eo9wb
hZG+qiKr8zlp9iLsH9Ua4U86+ffi9GXKYBDa5ntACsBUlppB1PBLrz8Ejwb3eylx
DwIKt4xC0MyvvFinA1d7wZV05qumM4bZgebhesXYfhpYWleFe0Pz7S+M5JHCyp6O
9mFAw49yGe3EvKtRxg+RGJL6th5UN2avR7VkKIBGvBwOQV7NH0R48/ScoKhmQVqh
e99mfHccBrNl3iG9J6j7Sz0HeL9L7pzUprCpJh6FBhIW/DSwgIbQ0LRrVvZtm0ez
MTAcl4XvrrhY4imAEoBu+n5f4c3Xzw3cm8FgPJiKYxwN0q7wGeA3ySOxNyCOjhWZ
+9HS8tIrg0u9FWYRSUPg7HSsUk5kvLGVkbyHo+sjdBLwgHEtxQsJoXbgSKyC5Zv0
42UwfbYyLi1DNo1KCIYZTY+h29hmUjvzed7PJAZI9+dpVlHlJpWcGmEQ+Qo8pE5W
pM64M6/axBUCUwRdZ7/3cgfU73rivPPm1qqJcCUBx4vaJe27IAmIXwinkt6i+0r1
hkyIPYWh2ULHffHSqIZXPKKt0bON/F1S/eFky0qLjooEA54I4s70Sp6KSSrMffpi
Sy6gQwe+hIW+5eweFQ9W0fjBAaFjb6kDNIGQtkjU+041vYqCOQbBLcb/cOG4CdEH
NnS+7XZJm//b0DS30d5xc4LD4krERlu7581ONhSqbgDiZbG9DVPrD5cgzKPLTVyx
mxm4/04uZ7r4E/J96xvclBZ5jVYlkZZh1M9MezstVhjEa1WXIWUOKmum+Lhb/wKt
znzNnBNQGvDRNfjf8YrpmPOhWXU8Cgr7G2sQ+lbWnOFihKrTe6rONGwKaVitehRX
jZHXMXUdzKwCmsj1Qefug9m/3oS5Q1c592j93S/BqfEoigqfBsWogVE2vgrGNrTx
54j1qUV2k8FBxgI0iwEqv2EvDzW1sklhvQXHaCJ0iwqArGPueeC9GscN+/ADfSHn
9hLohxQhx4PM0SEGn0jytqa497bdKCkTMI/6E5hk5mmYM0Mrb0p18HEOjSSpck/C
m+WfBw1VF3ReFYQCJPk2QQiSQ8dxZf4g2aA0RcJ11rmgq0Cgq+ns5Uew9DoUbEZ2
iyIhIC6X/uGK1O1MtMdToFu/kwTKCkmqZYUEhDvI8hih9Xb6g0+n6MiZrCYRO03M
M9/vaDEKGqvax0xyXse3CCrPZSDvRp54UeKvxDA0DJv/Tax7BNGTYZrmuggQgRqk
jzBj5/URMEQF5IP/sYX8ygZMtyGXkux2cTB4OVOH6bUnbHpnxaLRu2TxQYiFqgUa
2YAMeh/IUVyOYXdGZRGdS/E+16+bHVam8IqEzbMqBmHj+OcI4eN1lF3HmgWv3AuH
CrkDL8PEGtXSEyRpm93DAsxQg8E7jZ6Ut6tGhmSChQ1pWvh9iySUyyHT/0SogNft
TwUM0oDzqGKLnLvelkn+8TXfxgN+8Iy+O6NnFzOAvuot3J53P8ZNfsKABQYApBbB
tcE6DtvK7zsSI30WNr83ga1xN2abtIlIjHQ+euUhSPM0FpkjFcfrhmNy38jpKkTr
2CbVHwgEmHa8xGwVA62srVAYSMUeBIfBgQTXcA2ypk3Ims2WERF6mjQfVlsagX5s
RI5ctPaglozE8r0dwmEb16EE+NuZD5XvgXwbzjmLPAQ/9t5Z+gV5Qu40ZkBfiF4t
nrlvN89lNb4GK8QhaV3dlc5CYe8p9Up+ZhdbwodwgsKQUTz01UZJyJQkpcEKTfgw
iAi6f1CgJ+9j3iBQwLW1zFoiL2nAFUBueSdK29F5Lx3EH+3qatypNWxCPKXaE2JA
AXU3Y8o4Hh6I8MkszzVCsyqu45SEBe/qBzYvqXcikOxtEVM4HuDMR4SrXsAdP7iX
LJ5DdcvviHIAJozD3ZzAHjaQebf8eklqqS7KW8/xv+OZrzGq+0+2xkJwtHsbB+8w
V1w5tnAEKA9EElW+VIDogTrE1gZXgYSFE2h5bPNZLvrvpfBPHM0cewVO943GkWy/
h/rI0Py8a5S+Tcf3t1i2d4DUPY2S+/btktFNhHnYJWdb4RhreYeHDA0AT+bOg1ec
HMe+xd69DNDcSkWZTKgJ4A1SzX3VLHnOCN8ra3HW+5zBYkgi5oeDOXCrmJp3djJM
iu4qj5fK+vSnkUM9PWjqhtMq4ySacwE8dr/0FKcREVSasCTJMp4GiQ/1Q84qsJdI
GaEPpthPLEEzKpVKzmL/paz++RZMbxm+rlL9SbanDL2fQ2PnXmKMlxIDGNBplniv
XatfMzW1FktiNRVDpDKLDIe/oZoTRxFV/KomTwNa0puANQ9r7S2PPP4frd+4DIRz
vM5agfdY/16ogeIOEAtifKBhX883DMbP+lNRRB2muaMpaJ8o8o3zLFUaBoLkrAR3
dbj5MnXx9tqCiZqF627txq113mrhDd7QOlM4nsUzL7UxfvpqwmvG3xSw/i11+eWZ
0WN8HW+NV3U2GyDrutL2oTdLa2Z0VrhPIWhvgK//42rEwRH8P0ktiwCpLLkWMpje
NCgHVn+CjbqY38kVwOojn+GzYg0lGu4p5iMEfGt2Pnc82n7M2gBjbKYDzUZKhTRt
uTaLLiDM02EPPmB48lonWzJxoqVZGWvvuxI1NEpf1+O/PUMs8YRvQZBwzUJctEjC
Q9C2Khy7YmIMX6CV4I0WRDS/F9sRKsBNdTRsN72PGs5O6DAHE4s8OyvUOOTp/kXo
KwwfQyPluh6JehbHz7Ci5iPB378FMMrAw323c4bONTp6zDJny546clitAOw9WzJd
dqqSHfsohzt1FT73a9ycFRkKw0Gi91t+xH6BU3siOdVHgVGNiKjuwHeUo9SMh/3R
WE20frQYHmzeQwifS4WsLJ80wK9oUp8B9Rvt+Tk6KfHEoyW7Y/bOEsRXJNEeDw/H
rMo72LoqkFA6JFqgwHh94amDwL8q2ae23iKUNes+jd/5YlYb2GdBeBctIXbxO8/c
rFl9OlDyiVgasyTCSqYoV+Ov2HJ0/BfxV9QnsAtX51IKLQVRl0YVBLb3BPwyySqV
dYEoaLvtoDI4dQ3FkKjMXQKwDVN7GDHGIjyEV3FFBh1qrpPkSbw6pyYXClWksn3z
66l5y5Fgu0iFP+Sc1k3d5G8/Utk5onERqaO5uzzhDSX+mJT/o/ctfW7x5c4+j1UL
rxmwdPzmpLbTpZXpmYZuSwFafbLbY02MUXO3oalChsSStDhefr5DTc6ROoF88QtR
yqaX6KRLK14Ktizfg/c64Qn/bNIkOK2YtMBxEOgwwt7+un6edkWPZqOHUGnGY3PQ
I7zMxd5OBx4awYsTKVBqH5NjEYCpCh2DzlSE3x+zO+L0Snq3BT5fMwg+hJa9ODWp
7muM21n1oE1QW2rO94LcaGRFh7xX4jC1razKhiJBPLpHf2ky4bh8WjTrr3RYXe66
BamI1kt4D+z/wlv66oxOpuObd1eIxV9qqqkFzjxMlY2utWPUAhNwE6ZM20N1Bskl
D6pDqwr91FkwZTMOxQZZTIdn6KMewoxZuDH8dIsqK5VDaFru7llC1JpC08cr+Ipa
AMCD321A7UsfUSX4NGGUPrYc8ZITNgdL70Wx0KuCguOGYVsM65+vUrXeDwq6hXn/
C0AOMrjXt0tzWJxUTHEHaRDTFJZunc/zxNTGprpCC1gnlKrvMg8Cx+EmWUbxzBPl
cR6Rki0U/z7Unbe89NnIn/tsQ1wJJXvPRHNOBl95NtVyU6jwItixDb6c4b2jpELB
5cLfWkhfJnMLmkBo81/f8hlsHsKc4TC0INvaoNgdySqDlXwqz43yqy/tt1AjpTtb
hllZO84drkPKINw/qUQugUeSvDD1yoVBYTB3d0l+WXGSyASrPsnZSritebDKZ0IC
Uj6UsvmUoR90PAyra7w7JaotMxtB5+JA9vHr43vkUwTut5b5mV/nBlpDzePq4CLz
iUazzfZsvmcA6Sltt8WOaWrF5cxE0CSpaP8wxU8BZPXmUOcEOdN3C/Xv+QagtfMU
moNOFE4kVOKBeMMwIw8BTHUr5CLNhWCgyrJxMVpgKAs8EgjYUdd0Kfg5/1H0x/KF
75gkF9tN0XRlIjaTpkEwoygbS8DH5YZMIyGeIOAu8OZFVxOLJoouoDTyLYOmW4HT
VKfl5DWZL1TfGNxtW94z+xZn3/5/Gcv7ZQV+ScQDG97Pjhc8MIeKW8zSjpEqKH0p
SDvrMNlEZ19hW5DzUTASKGSi/clhJpQSUipvktj6Z7s8of8B3LEEvAeOpUD81VcQ
P8hYxjCz45TaqtMOIAuL51Eo9jCH/v4zCKFFGS43RJGkqSRdfqJV433MVR3Fcr3p
dk2cbdLH1usOqGnNGKZcuhAy2OaSWBf4Zqbgu41C2Tk+y8DVPKFZykwkaoHYTWbi
dcsN7frC3rxhaEgNaSk2HT2ZKFhOaQcrfV8OdMyRTp+JYiZXkSJ8PIHhjv24+peO
u38PpZ9+0xlb2LHJLdC8tBatL5wijIpx9QNCnUTlEMoIdX+0Na+1di95U+by0yWx
c3F82T1eCmP7Wcf2rBHl1EgdMJIAx2GrRSgaup/U5DjDGLrAFn+QZ9WnRDx0RXDT
bkCIT2M+PT91ofZkCmpuAFkFz8gB9qpLk4p7wAvoQITanGuOQTr7E046Jy46VB9F
nW08zHJlhWEa3YBCUdg9BJN2ILyG+QfJn3Zm0BcQiR8N65vbP7J5JyKzgVIHRyzI
T7WL9eGmU+xt6LcVAC2IHDmPjDXHeIWGMpkcAZ4qiI6jNQAYJQY+JflbR9C4axzx
eRiyB7sV0GD3k24dr17fNjw+X153R9h3curwjisJPLkdVYb/PPxk4r/a0CyfTHIo
dU4DlLYuCeNpVW8lqQp1Y+n/z5p8Q28wnt6yrC2Oh2Q0crzclbfEW0Shw1Sj2yPJ
ZItG98Y+mN4rnmXHhy/qjFh34QVqKy3IG/QAybv/1+V3q1lldj3yV5LEIjuCX91v
HjitniTRGVOMlL5hvtgaM4FUq7b7qDn0WoeATSuv2X5m5/22vdeXvGamQOGAsKHj
4TEav2N2sjHzph0JuKtmhFC0epTLaOMKkQJY7133ap6mK7p1+yWaYBlebBo77IEW
DBPLTo3JteotQ2q5cdMphcCa66XpfsiM2FTurk5mXy7kgilsV2fQydDs+61K7Qt5
A/o4v10D0OTVNi89081vkPT82ORQ5A/RZjwzXuLrdDSeGhnnhGN069ynVNxCVomZ
pTpC/rCWCNvTav21hILDkdkATUMbEg0uYPTkqXve0ymTQXPm5X5nLXzMzqnH2yzW
XehzVVFwtsjDTETflZNn9nNUHZqZulQ1GWtX6o4lAdyKk2achTxKIiwTqRFgemI6
lCIQ6qeiwc9idveVOkksP6y6sRRC0jGLZ0Cer7h0fhjM222ZpzarJuKr8ggwMJEQ
8tw/MTPrREAvK/gpJStnsVDaob93mOpGdxhtLT53+cXebkUVjEdpACyjVYFcadOI
8zApB3+9/NsuDwBSEqE5qCdzmnJ0+M/+LXPtR9J+eDe0wvlvJyXJegBUb5bp8OWm
7TZSQHr/K/7ao84Qowm+YVTjKQLUBMhRMBZLSbIC4BrDEenE3uunNeH0CLkq8cn5
OhTyhNQvCRC+Lip1whhooMD78VhNIbnSVVWPTeZmPW9N1/H69cLDIdXMxs6Qeaa4
6TwX1GgLaGhL45txovmM1THfwraHrv4RwKc1ABUoE9MRmAwnuqIoq7b4Wl4zC0Tj
Qcl2w8rV7hWxO8H6YEALxTD5LCYieAJoUizCz+qtFisAjGrCTqNYomIcfwvGxZis
+RJWVJ4Aw53N9idESe7hstRFV6b6M5WGYnn4zaPsHo4S6hO4UEQH/+VsCSARewDB
oIRjS45ZqRLtNV7R4igSyGAdKZbFXU8+L0vpkIgWBqRYpuILDncXLeSzi0F8mB7O
Ur8z0h68B8T9byPRRRQCzD59LtslDaHoihUzYyamb3GCi84cH98IAyrN4pzmcmvZ
ItoXitRFuGUDMbVr1mvrYImBDWjiLXX2kAnarA/F/CB6/Yo19bXA62BY2RfESuOR
W6PMhPci4LcJRPdCZeGncoTJKGbIxzl19cxcO6g+ylrsDYJjhnc5KaYRl4Lgu9xp
SkYB3c7bgjlzjqmhSNs4jDMjUlo5SqMoKphXs2PcuX4EiLHx07P6xJdc2fy9Lemf
Zf+RW87NIclOK2tSSPfOfuvelL/sp0Qou63tpC1LvwI+f0Ig6+Qbcrlh4cG2ybZD
NLVR/ovjdRRgKmkCcEh3zm1ZyLYe/ZeO91RIMuBCEenLVwsX2FTCk9p5p4qHIEmL
XwWqhoN9L5TwZ2rKMR8coMRLa7u30wRYiEqApkmVGYuV2oo608hfMkh0qj97k3V5
p5EyWuwsLgnhS7OBtgv5WVJ3/Cs2nefqaBo3bthrHiErAa5Qczp+Ke0RDpSeWtaB
J7CgsveH0uN+Xu/5GYALdyDo5JifQFBb3q4tgSyPM/1PCw7iZqVXhPN9CfQcVxgT
xCcEaNdwdTrVNVP/z/SflrZ9p5vV1sfrFs8EQeO//G+CqwuAOylVGWGJP+HL+rPO
esuKcAfksHxROP8OghBj6yXc8O56zsPmNIIpaO1vBhvS/rvG39sApqXF83YAIeAK
10roDofbuJd6FwHxvrUqmsxxMVVkQCHwycBpwXxAK7WznUZQI7g4AcgLy8vBIcx2
6gSnaI6+lQM9w8maEmICzc4HckOiE+xqWF9HJhwsmUYp5lCyhDj+150b8vwOcrtk
klKWooBScFY2/M0rfnzQ/7Bvnlg2Za2JVRhHg0D1s720OAYeVHaDdfUhtF7bx4W5
6HzyJmbSWDPtqvSoLngqNVIL9LPwiggyFiQyQ/lFKm3i78T7u4lYXkSxNhv8VGAD
itg53QEsXxBJLtXPlrLMGbOekULN5l1dUkxsQKerRpyxBHJdGXBhbl2v2ltF/KYr
vMkSMbmIVaUQf7KqIH2v2o3C3MBaNmv1MCPUzYcMPKWbcl2Rq3EHt1HgM9MB7kvx
jvYKVfJfU7wRRvjiNeQxZ7Kz0q+7QoBwKr7Fe+KzSXimmfks5+GAapkA6Wr9Q9H1
qZUFw8HMDKlrkoaF/RrCQYOe5o9uGORXiqJH6XMDqfj+ou3l39Q63WDe/KqyoDeA
Ahbc+VO/y0xeeS0buBeQ+yPo0TibppDcddWaSK6EFbxpA9scgb619Ipf/HTRXlgZ
y1DYRBckb16w5Ekh+MKTlF4HijgdM/UP3lr+/bwsGTijYp0C3mZELKGoer6ri5sI
EZnesVjRin+F88ekTWuiTuIpItSKOj6AkURPhBoRdLEiuM7Xz23nEo8QxDIKvYUC
rQltlt0sIMRiqQl1cNt9aqcF/OM0uaTdXbxeE08X5l5xDMFOTO7KkpLV098AWS3Q
FvlN5C4XNipGDOoa8779uxWOaoijVxr64nWw55i7DFOOLDjBAWwuNBffbvX+6Jpx
ehTxzYNjXEQB2onQGm2hP+1K/9CsG2VG5zfhJbKkzey2QIxsdcQi1nMiifjdnC7/
yeC+W35Yw4xJO+Ab620ZEdF9TjETgBEgGakDTTas8JDdjOn6ZA7yDnQMSkyFpwpS
LIKhs5+05tEjGR7PyKkQBT4hqMqtBuuGu0WB7dt3FM+URaXJ8TAfNFjwYJlvok1I
50lP+E8kWBg2cCsBhmG7F5SoZkoTL05laUyNi8hWua9a/PwBRQq5U/rt1a23BGBL
Gba+K2CPCmit3ZbQdTXuBv7Z1Hgzruk4bKI74iKEqABZItdULXKw7u21rredzjOo
TSEkVq+iPXKTg2lGZfwyq0ImKCmi99qurKrWDBPaI04228sDx1hgDOTpiaiRMxFa
mKCdsD0203HfQPzbWk4dWlnc2MTsNIOfk6TxlI1TpFw8OL+OoqLBGBmHyQLECfK4
ahcUhod0fjecJAA3p2kXAim7AHu5CtpI+E66G+NMqP6VkwIG/tMb9K3RXs10Wp9C
+YsB3hUd+qr19jddLJ/Ua1oxfVwtxl9bh2SrF7la6ZuvZKB3KV77lOopbtgDbLKj
uXY20aZ/5RP2577aaeobz3r/2gDuFz7LKhh9W3NU3g/8CuVo+Fo3tQzbkv0aFjeP
kAusNJjPsx4PpJTkXn2GSMuni/riK30Mjj7ApKjD154o3Lf93kHv06jPz6sPf7fm
xFPuZL5QkGh4DDhHO6+DbWDavh48Gg8eUs/jaWcGwtjjnY+4J0Cd7OzdWk7QZD+g
Ucds6DOeVisA2g6JlDcRZmLynUHwEs0ofUdMGGBcCyrc3qre+aKIcKv6g2kBRCgr
n9i9DojbnnFZyR1CwocjYkdRrEBlM5tZAtAazpbX3HCBjP4jpr8bUfCp+rtsR1tM
BSEsUhXcNTf7qHkXtw3gAKQralSRobyMuiiIWiZD3xpKDFq3Hy1m/wxONqJRyf/F
GNmPuE8zl7Hrx00QVFpAksZBe3JzT5RxMse49QsAQHFRbgC8VRtSIsHs1LTN0Lbx
iZ0ioM+/zsAVZBVIcXl0A85hFmO5SM6uYalNXuRYc5V9PwSnENSO168unOVGOmQh
gfyuNBbbmkkN0XpjLtXBvRBqWZ4vR+96w6YbYuETnfHMhlyBpiSBBLa3c9rPrBpT
duas28DEsS96vuuF8V2CWb3wLqiHn7oR27iHnYgyCVYV0KY7Cr8E1h+ZpCSoDSeQ
8kZ9WL54pnlp4pz4t7xUBFloqJxk5gLKGZ0K843uVTT1sdtfBe6kEbTG8EQifn/k
RfHFNR+MvjofK2hBZz+0Bs9itRPxGWQ5n9ir4bqxs0UvQkDcPnDsS4/UT6sJphnZ
4VlmdDHvpEJqtH/B95GGgKz7eguZ1ZG9IWymipC8phoByCuWNm57rCBxevkRMFcN
EpcaOevfTSrra5KcHFIy0o124M2pZhNIrVzpHtSTNbgUwYLNv4mgtomKSeE+O6Zn
wCGtuOqscq2FVwhyNPPcql4d/nV5v6T+4KtEgvS/w7l142ilLqfQ1hF2YniuyZOE
jttq6oopFrVxbjPkh56h1nGm8LJ1XQuGHTxZ+uo2CHrIUbmXCWQsjO+ctpNZ+eAo
SJubi6FiHJkAZ4dZ2zKobqnBTMVpuptHC9S+Vx9GotI2mlrOjn3Fw+O8lLe6XQja
jSyKLBcbJ/VdOqnbQ7ED15vAMlXfYJFkB0eOT4N92WwbET/WN/jbNnGzoZ+b9ib7
ysTkFQRS6ML+O+JUFsIZ8acTSQVJppwDV4gQFZj8N9hGQ0S7D6t4JasMiEceSHs7
jKnRNRqj3TZt9QS+Uh95goWdLiTv0E3iwVA0EiD6u9RG0brYjhOI1WlcyErbF23E
hYXBZ3g+RX1PVM9Qef/PaDL/7Qi/8tM9PW2mf8gBe3W6AM47DXG05hzFnTDEyeNH
rFOBCcj1YEhSiY8M7MBuzkp1C7zOGfcDINPUFgjPdcFLPnzXTBQN0hI8R2rzEM5w
+qXto6d33RSy06G7k+jCWo1NE2Wntsko4/8QBwfcqbxck7JKVfaqeYoP1ES3VQQP
+yt+ZaM91ZDk4ZEe4GKgtLc5ICRptsbf7khO+Lp70dpaI9QL/eFkmw7FQE9s+rOs
bNBLPv/TKaB0PDVMQTwRoqcHBx2L80UnJvltGKMa1LQQchBNmQLmAx7LOfx76g/2
726p449cvqbQ27aGf5C7Ch8OwiUyCKDtSRgXdqLTpOdQ/Fvex9iAwsuMzaUQJKqj
JD8uRHa9Wpxn/TTMytdLMQE9cphvVp9TZUKnNoR/acsB86S3uP300nUsXFBf1TCW
WTfknMqf+U7/5crjriUERDqk5xIOos92HTJ9jlvqRDUEgtLLVU17GhcmBCH8B4Wb
oWY31QNwfytH99Zi4/NpCWkpHftXDo2Pm09n3kJR/ZqBEzZInRaO/R2jHkM7j5wa
6JwKTik+xftwuTmqG2jzDnVd+nsu1nxwje2Itok8M1MoO4nmRv2hX4hnU+z1E4mK
Vq9+lBBuQrlQIGnNoAENWP+VjdoHqPNOJRxZ2bPEQCCwsyDnv73UNomh4skKyZBF
gfUC8OoutwsE19op22ywtDJFk4Y6FVQThdhhJjtvY6LdXmgamr57MfFv2qXKp5GU
PM9Bb+fpoh9sptb9gZVNiBAeHePBr3+4KbfhHT1EtKNR5VTzSBm66plqs7o9j3TL
WIw/XKlphCElS7E1dwzZ8or5INDdJK2izWuvwOdQkWUG9qQpHxGbix4IiUPFrdwR
F2CELHQIuTlJO6Y3DDd7m7ZQ9IdW3PwmrNogX/0ZMsBpH9O0HKnh27x3Tlg4SSR7
qwDaFTpRayuYQ3Edo/Iif0NKKxG3LPIKxR+I8lmzCq/ztHueuZ24pWJkvWGHgq8k
VydFKiXOrYlR4ZqrPUgcWUWosG1lQH/ELddvkNh912LA6eZUZMzHZqDb4KuKBDI9
cdcZOBDLHxeaVYZVX4DhxDdipCN/2U33FAIwf2VeKu0z6bDClkoBvpAPNS+16ppw
dlq2UKzULbg2Xm5TObk4FfFw2tuiUFf3h+oxQR2ErnusG9pZQnZl+8yAmRsZkp2L
1LfrMmSWVTtt4nwP9dMqQaZliFNNbTA/sb5XKyhwynHDrMzsOq1Jz1zLoBOqu30H
1l7EA9JC2lKpwqucDHJZc9IKPoPKDJF7FqOyvYiHNdhrnlmDNItCubjEdHMfaK8+
ne8BK0kNgabcaTEBKfG4SlhOA/uwrnKsvqBK8fFXQIlXRj7zRKFNRQScw57plguc
TnQzqm7+2h4qbNP+pJnFRjhMhgMTyKAxVNOl8Et8PEOj72Znbk8/mwK9D8vzjFXQ
U9p8cCp6oqe+DZ8tjAtXZCtgv4oonLwDeRoE/uVEKs+axC8VeCiUV/WWbJGVO75W
kYLScDQX48zJJhdsnAl5xxRmYsc6ioCJG1yI83qCU9VjKl9cIjWTELPdooWXQCuR
cdgVTE910r0A1fRO8yag0xF4OTSLkiOUCp2e+u9bTGlqyRRLORr5Qzb6yvNP89Ba
8Rct0J7Id4j6VGplYdbaqApe3fxzk3gRADowfpoq76oEjsnbvh58NeCoQxNR77nn
6bS0tHoz6VXiXTLiZ+p8uJIrOYvKqUYJRWfO9DAkN49ErsBYRvV4NmI5JM+eRduk
VwHEXDnzuvLwif7z5HcQ7dlsqz39tG9d5GO/Mqyrl1bAqIo5f603DBCmUmBIrT2z
FooctVsMv2LVgJVQA2WOug+eCb1vXoJSP3FDMHQliCIcc0FcMQ/C6B178Ndh528s
kKg184UpzaaGa+MFrRLkS9tWF1STVKc7K1rskqn64LCZuBCsiQUtG04DFspLgcrj
JQp5p0RR9WwK5myCgAvdAull548nIF5fP/+lY3by6wPZj1Iea/yYsDxdyTYSw/DM
g1XXpNO5cFj5595l9NA1X07JvXwvAPNmkZitQCrgClKy5c3J1x4p0c29QAZ4v/Rp
q7NJOy+/5R9tPlYL9bdHyCGTCgKHj5fUuaXhdRVMYN38Xs45+X0fLVMxPYBoK9Yb
sI22h2fyfCeVT+klZLvd1WvkcYDc2MaKQgfZBUCzfmUNmcrLIZwG5+1n2bCztw+l
pj/8nCnM+9oGFs4CC3hG5Xi2veDcwrI6n7rWbZqVj+cANLFz/dg37nEdx4Fgoug6
c5kCMADiGwkvVW3K2GqanmTLjc6OBI2HXlBLKVRXQIbpRy8ZPw5uGHy4k0rL4f5Q
vVeWVQDf0u3v9JAp/Vc2QF4cwcKDlQXzqgCDSRUITwkJup+Obr7pwNdiMVqGMTY5
AXpll3bbtNbSDizOR1XEzgKdtHhc933NssLYBA49wx6lvblu2UF6iLHmTBFEXr/y
Lw2pfOTzyE+4o0nWCX1UECiH8aLqA2MY3nF2EH78fUXsoB1KaQNHu1QKhTHCP6/Q
FGmdYspyc7Q8lXJz6sNq4kWlbK1WMCBw4nmdSHfar7cJZXW+wM/IXzCUZVHvrkzd
S92X977GBJK/BY759be+rMOXrlSrzBf4ujiULLShIKLo3tDXW8OVv+u2bsrkjPum
2lNit/zew2i3zEnDwiPow7aZLLtMziuNnk4tP+3vGjU/EwjfukY1fs27jf+jzZ9d
Jm9XwBEYx9xQ8jh4vKmcmYFnVjGqq5nthnx+xqGmPu6Ft/Xo/6Zo4ZlY7d3ec+Pq
x/IYVjqZ7dLytjw5Gz+UkmWybVYo6av3WnPkIrSVVnAY38Y0epNxS9Rgti3xlFOf
C78AdSJBtexiJC0SsZKHjhVEhNJZ/HixnUXYIHv/9dXezaUYTajwp0qHXmva6vZL
t7WmTrAhd4L1g/zcSv/KYaxmz7WZwDB2t+dpzfpZje7juckNgc5vv7X5NT2oh2yQ
8ruToAWMlYmMPzB9LWk6shs/HObROGI8NsAbDYZnH+2yVUMzgGdb9mHJ1zL/Tnii
M31pa0lf5zX3IFL5wQIV0MxaLKqqRde88HDcHFPbRWccSoI1KhNmugLvC1OWmWtn
tAcsXs9NsYx47GJQidgQHRNBCvsVqyhdX7IHNHi4j35hIj+Z1sIreCS8ueKe/CoV
/m9pgzTOPQeyHlEHK+GiUqGzNZTHqwh4B8dA4iqiOOnoKf5yGTQfyLycOHFbK6RW
SibidmkjhJy2CYAuqb89qy0imAf6ijfcW7y1PhasR9D87Ehn3rXFIMxrKrUj4IPz
u+p2Ar5KvFoaAwGizIcGryRgOvsCMZoEB1UNM0BMkYcL3i5teIUbUDBHPVp2vySV
aUafYWItw9qMI7aWjGX8AUUCdfnmCQHeomZw0r39ih0SZprFufNbu/wxwU9MqyH/
T0xaXSzMaq7oU2+/uDxA9hrKVHASeMN4daTUyC2OEXOp8g1/v7xCjZvAdFn3xnxP
A7dS75amkBA2Wwo6Zsoap+egXFmbzmy/wHZk7OZzx4M8sgHrTlg3vyqQBCXFgk6A
iZUGeWmGWILz7ei4ixdpjO79qC0fyMrTNfe784/PGLdHELOZcx/BbY4H6PKuuM81
gyh3ZoSrHmgrNkvXDlh8XZ5fQDs4c6JiDoJHkPbvdIJ47k+nMTvwLegRaagragf7
aEl2N8Apgv4J7YfIUNZ7bOp4fRpU2z7XOocfy+wv8P+4ZL8YZCSHCgujrxmWCg/L
QwH5dZiYe0bu7PwAgnYCIM3bA3cY5QYPbVhMP2jLmEpJ26FbLllyy4Af0vnFnWLe
mFU/0zPEsh2uKR9t7dlcZp2vrZy0e5rr0h4FKIv/TxPfY3tO9o40Tii9muWx2g6u
MxJkxiEKu+DCXOUGFX4UalFS21Rn6+ChPRG5zfdOC7RpjUK3hrbooF3XIhbDxzO7
Uig8XWoy9J9IeBuceqjGrUTUrXwWEOA+sDwAZwc0lA5dYBbb13Y+JT5IyS+sDPni
xs+k27GzkgJCVbqyFHOwRfzpL5QSEZo5GdPNblS8Sr/cFhgbSsiQVHdN5U4bX1UP
fCzSvkeIwU720OSPaUdWWJD380dv/F4aJkSF9b3aCVKWYhnSQE+C6V7ynylW9/Tm
SeimRZOjMbl8iI6QIMOyBvBM6hhuZJ0CR+3TnoXq205FB0hNPY2kfqj3r2cH70ys
2SZT29mVrgnP7SoSjp+VLpXlNgY2GlOZOLEmmoZct9e/Fq7gBBK3AC4j1izCtt/Z
8SETrXVzR2BZ3kpkAjx7D0T/UFX/5ht3tQi8ziy6Fojv6U1WScOnEvKuIvWClXvi
c5catPWSjORtmSutQzmtTrI3moXNAO7mI2kADMANCDZUV4G05zHEQ5jhF2noqEPR
mgdDMzVqkd4ICIn30BRiGSBFoCRZQam75D9620IulovjYkYobckK8Lp4Y295nLEm
zM3SZSBtX+kCfb8ZTbzuTQpPxY5BP91R0nrNhzHd3ELMbaRYcx01/ieQa1f01q0L
HXxFXKKV8zV8wvs9shYmT1C8alXgTMauO5t4FOv5gCm2rYG1a4QmUPp425Dxc0I8
Mwsosr6QBjXabH2+BfrPsAp1qjsM1AwEWf/DXPhR7izNrxGQM0o7u/dmy0JQOjiV
rgDCvGXYCJjf/Yj08UISGEqOAjHqgbaWGd4Iwyag7ztjyZMxc9YYjoCkDqgsR5RB
F66jr06P7Kc5gcaQ6m06L1jjK+aeEOqrXvsEan1u5x+8lxrOJhz/EOpcXezEkN+i
rVSCTrqx3+59Plsqbb8+zJRT/VnyuS1aJTK/n35sO5MZdQJIIasoOhGTq07JFR2q
vfPhdFbNoXoBrwFK+4hagZj06bLGqVxc2wEqYGpHttPBBRXCL14FuBTFzcCUIxDD
QBJPt18ebScBxAZpgeF70roelS5kiOWGhQuzgfL5B3lJF9LJFQnpuKP1vNbFY9GM
+kbJPOjxGBOsyjDHlbU3hChD6KpGnvkt9ABCjEEezhNQAu070zsS2bn+UkKRv4//
2Y3HNPmnMFIb8uyC8SCrSgDiN7kHwhGKtaW6d0CZcrcliTa5hNsYEiA+wTEqWmqi
AfjbHYPs0d4QJJ4WfC7SySz2/kOHyWjJPlwHhHktwe5Akim5fnK3H5p6hDJj2A8D
R7HwtDmFakP1SIbGFUBS0vThCJPoPH3stGxcpSuxOwRn8ZxuWDeJcP1qG2j4IBX1
OkPQEyRlBo0GxaiOiLHneE1oqGtY6ZIkocYfB0gq+ALPxuPTC8MtP6qHVNeniv0W
y+h5J9SEjZRgRn8przHsy/7WgvES/IvKtCXtOAfhKmqlQArZTu2OWShOWZycrrTD
2op5gpUWXZtgzZCtjtdrbGGSMZHYRcBPD39g8rXuB9vpDswaqar9lSH46OiMq9mH
rOWE7d8okno5PVPZTHqgcEoYV+VjcLUFWCa8Dvbi2zBSiHdcg7TPRhQaJoWGxvTs
L6+7MyzW+cZ6QYJWV1AxU7RM1LDmlTpKchsstd4impNeYuwH4fTz8MtKsiRY848q
cjVGwhNrvERDPwGwMmW1AgwOKlStB5mBESDe5HeQ2N5JC/NghNTOOaRf8j5O4BkN
sccDK+amx+7W2xn51XJUtkrVrk/Lm/sttgPZueWj5M1ybn4eGh/+HQ8kDBkChS4Y
hWqBvhFsGQLpC86w4x5OlcYKDzuocfIFkb7QIuXWcFTi2WY8KB0uttxnICvi/hoq
vOviFCz7C+n5axqtA5hRh0dMUlQLiFNxqcejaOqYq7etXaqYhUtvkmFUEKWet1gV
O53+qrrxDdyfX4QIsp/bOa5hvBIvVFPoWMKO3SQ9DeviaYERgoxS0Jki95CKUuri
KsQj60lOM8f9Tvn7RIv7+GFfxY4ZDx6wLGwLoaXFAv+oHsXjLC+c/Fi68vTfdfnG
MLww/lv3oTOJlIA+ofY7NNzTskAN4vh6TtIODwZXEL1Wn/smHUy0RxSZP1Y/nZmJ
p6ujCIOrAw55XjU0yyNmyvWEvorwkBnPtuTwBMF34suqfjPw8IDltbBITxf1m+y1
/mNp92hiBVnZ0Eo4ec5psIwRdMtyICSBq/STczULxzJLA02iiqHwD9k7lOujay03
bLcHpDK9Nn/ZXcmIsvnJo4NEARZ/SMOeti89Y1P/Hfep9WEnnsuDZlb9EYExxwMY
8zJqIOqFfVkhGfhfij0NxkUfCSG9kn8Z1pVUswXygR+rJk1g/sPjrWNJjMZVberE
7H9p/TzuXIRXhIUtvplTzaTMsKKF4eb5dOyODSIx4+zTMou6+RrX0sdPmSEj/SgD
26LONymosk5Q9CxmE26s607gUE5ixUPcN+DfXdgN0JpZ0Lr7COZZH/4mfdGhgMou
3gPObjMxvmmkwINhcDx/E7GVckvEuMcmsNFiQkRbJnlDCFuJLtbeROQlvd8rGy5M
QeJWCh4hBd8tVgsPKiHlpgNHna3VoqHS1uB4U9TVyAGcxle36SXzATDBmPXq5NFK
OXzGDnwqfNbC77h88au1wp3s4sCyZIxZAcV/G0H881yCfdESVKq+/t16gGU36x/S
/127fzE+7fejC5XuDpACQYACF9cbB0M2yp5Gq6oXkL//m1bSshAkO0mseF/sknkW
VFNWXZSczOiiXIxtHiZM1ATwm5NW6qLNbFZZLhMBeUUSNv48xlAyefPwbXDTdSId
zvvuFHObhBgg4YMu4Up8W4kw2Vg+0bjjZpVE6KP6/pcGw9hHjDF8XECz53fKiT92
xdOYN9K0qgsbC/4W9lS6WdreRT6jlSltbHfvMe8ZkJiQsikA27+a4juncyrF3nqL
5daq1fZa1cbt2uBmHGIpLmFLhEwXn3b8ar1Vs3fbJttHIU43m5zuDE7SOFCMeUXd
Uh8UPqHOjMTyF0hYMGCZ7eJqQ+BxQ0mG93FNTWrhLFyM7531cmbAHtQu4REwBBaW
J9XEFGSNykSvpB3FmMIDoII+tChoSMX4QOboXDJj4QVdkrRyBOiQCvipEvn9cfYk
QR2NZMMLJxVSkso+oAi9F6A4UpxwH3JVnfXANCPoG5yh+8jKlkg8lGIiytDnMKeg
q2UtNUl6QdlhucKacV70m9dbwqcl+zv0I6hytv4T3FrLHT0l5DdmaJtLwALgVhRW
YY6s/mRNaUChNUF0TOnSXc/qW5Cn1JY0djpzDG+Ya8tA2Ejp5GpU2k+C+8U6o+hv
WocR5LkQZKeWIujcpGoYP62LPFl91J49wipGncaHTEQhL3fyBy+Wwb8ituHhu0k8
zmB7a26C+yMjVZh7abp4vxjLeCB56HchPP0id5XPktwdmnjv9xXtH9M4GHA5/mdW
Iei3yvxOIEvFa9ZBH1l/wEj6dADX2K6iboWA9FTDutv/xT3qFHPbeWFGBj2IPtJD
1kaVuWQlnSy+v7ATLDqY9ZTVNDhQZU8AVVh1qWDzK9BJjWoh7EOoHuVnn42ifZ4x
53Wr3zLo3PEjv4jfCdie122bZvnzy5IKdWw4Q96zyzbu4x36JO1KfGkTGlT+CBla
y+IkEcE7fjAn6EMdlYzwSguKYEB9czXiI9YMlc95IaN1FnJQmBG+2Om9Os3QslQV
L2YDYdkl1HpoITWRqffY5jhypndtEl/37DA1kOrFL2HK1oe4Ng93VSdFODsRRfOh
Hzx+J/BstA6EVGSmXQrIhcYOsYzbA4TWt5bMLi9j9YF0NsV6Ew0gy5iU2UCInJvw
QDfv+EuPOYfrKR32cQyIwjPDC/Md7A3x3Sl8hiwcbowkffOHBd69k/AvZ2UmREAc
h/QXR4dd5knzmnCTtK67u8CTEgSBiqsp4pqLj7j3WZxtdDeXmI2mtFr7BNEWId6Y
lCbAOZ8g1XZGf2ZN1lesaMV6dcocxQWI2qseebrzYgsmQuVZxWvAVgqrZ5alMbXa
Pf+NEBbYAWZRRe0nEz7BCNkSxPInWjjo3K05fbTjwdyQYIMB+kF3NHYipFoteUq6
WtEFbKPER1W6gEZv+rWdh9sf5HzQp+X9FaLs0Ey9bVgknyQNwYmGnpHfJwW+3DBJ
ROUUkKMVDTnV+qa060cSU2uyVW0htbpGJjBREJieonMB+pt0+RFw1LR15esNFTFL
rI0n/nAVnKfBJfz8Dr+VcbJGOGs+drT92rCKjmyk/td95aP82kXnB9pfV/FSp3e1
PA+jdU/2tGlvvDD/XQh9hl+LPBaOo7dXJoY33/Oy3er7Nc7m3FZVY8Fq8yjyzxj3
d3aR332Pc9Sgc9zk6N7Pd46yIuBlbi/Oy/IUTBus83824SVFiM8XP9IpnqLsPe/A
i7UsmNnwIgYgixo1KKTaclw8VCrg+X5GtLBDDbzzofo8opwbAAPoEqDnssMQ0ZTa
Ndz7N0khSJd1kb9OgPARUpB+2TFu4MiRHbDNNoHYfWaJ0bWmSWL65M4VJyypcIdW
SnK5aZuwXyMIzNQHI9VZ6Pl29Wv6RlDE+syQ06tzFZUfYmrrlebthWiUxoIcFp0G
KN7viLwAD2J6TLgF1BgGq1XmG+AkISsJEgIhJce4F/2wr0exXfazvFusL8X5P7FS
6o8hWjoB1rHDsnIhn9QlDuZlfFfxWGw1LbeeYiOXN9bzk/DBJvxI5D6qKwnZwZTe
sqFUJR2IBTdgfhu6rFvOC+xKkvROL+UibAofs4GLga81npaGvIUOFNDvjqCzF5fi
LyLj3fK+pA7FpV0Tzcej7n6Kn1NSOvpkDLUun56plbiw5Up72cIQ/YX2OxjYyT0J
k1J0wBWYRqu/pp0rwAVNbsVZDHktTx0iKTn9jKpc7u3n+Sey2dxmt1qvgxnlHgJx
WGMEzc4fmIyCTa6/XepiC+sz3Lqqzx4nuFH3CZ1Hfz1t9Gbjsn4ao1IuH1CXvRpH
xt4PToohiZ+LVpPmZE8ugZ6xStm5vVPbgLGZMRNM1ZXD4115EorcM5/7ymx+Z2pc
PKqrlFtF3D4NRy7N49UA9zidhjvDin3NxEJahb37OP30bVSD/+Mqfr5K13fGQ1ko
nLMa9RSGd7Zguv1NyghmIbpkc+pofv2ZCd2w3bjnu6gAZRHJfCM4RsWLK/F8xHwo
oWb0kImWFLQkXzQEVG4yPbwO9uMpsRfue/BFcRvVLB0QDkPLuYlhDvIrTysXNKik
XTnIhxNp9g197aYaVU24TCbbAJ1CnLSQJ//jXn90hVlvtePwiw4mnBHg3d087vqi
TdZmxSSHdqeRBI0ofHMUN811qwzDayQm7vGZwdiuK9CuA600/invxrjyDMCEChRI
SiuoiFMzi0xD5GAGNr8rikSeY44YLYLFCzxikHM7A9obMTRbYJnZao3b+gYBRCec
gMpMbc20sucXXRQwJC+39sVRV9ypgNBSVwBxZ1BXaBAdsuuilQsn/H88jeSaZkye
hT7h3LPXPocPxiUCpk3SefFJex91HbD2WK+As2JWpug6AstQb1bOmH+1tLciPvMe
bp8avGXphleXCpN4/GsTCsDUxzKl1Y5W95HCTE8iaH5rvM8EY9Wa7jKQ9K0jxunk
p+4RQTYKe3qcDYZeqBVbaMvCp5uGbwMNqSCamvuuP1A6bRvEs3951v/0v7Kc71lp
dEdHf28T32hpUjJzrgwqj/aqu2sq1IxHybqyB3WCeYA+yw1nLd2eG7D1ZsuqIqva
DxNxiUqUjU9hBUzuuMP4HyFT/s9p34oWjEjnUERqQJw0BFaEjUY4JFAfdkq4SgmZ
pLCRXyExOzDybRA1bbCkz02lHQ0UsjaESQdnqJY9myNHFOJgp5JTXNFZzYgCvj+M
r6Bv+8nPpBt4jHTf+fYCjMLmH2hKZ/FBAZXoXIB4MGvpcTqIj8kI16y+Z8E8KjW7
npgysA+1jsMwFY9/XVaBwzW5zF/yVVLLFOIWFrafH5vt2rXAreBFIFwq8UoKxbcx
cJjFSVRAfJI1mGsuLwvQAbqn0vy9RATYqxZk1tXaiGjzEThKT+2kQCpQKKf1e8IE
gE3KaZ+9dQCCC87MtdcJtGTY8Vz5bOSERCBx4XBI+/ttmptImx5/UwRZZIIa3P5e
TDsyTK91qa5Ofu/0qie9/2g/mMC4yI9ByOpNUGBUy8dLCTsRCpdXk+O1ONwVrS67
K+qYmBFy4aUIZ4eBolx/v8xs0OYobNMpC/2IIGRsSYqw7IINnBkbYp4huUsR6r3/
ZeC+uGGy4EoABnPETYLWapL9XzNxMv2OnaPbI9ZKoqg2vCSBNN5yuDu526mgXRZV
ii0JLGv7ZQvbmoGe6NlOyqB638oE14URR00b0p9I+IbqxXuA9GpG9r8Z0IzA3GJq
gHK029HoKNhEA4jFJRx7vIbVa5gM4FhrJalzICEFapvWxBv5Z34mKMV8oTWea0TP
VDFrtLiCBzZCUUviK1fQToGQGQPU4C7/d3xAyGkaCF63HHg9p68OC8BJHKLRWxsi
+7dkldfOdqn6JnxI4H35IHJULA651IqGspeR5xnxSYE=
`pragma protect end_protected
