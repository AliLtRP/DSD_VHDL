// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Lttoto2+LGcItodfs3c5ViK36UIiuoXaVoOZ2fjlAgYiKywl0eKnhGSjc9C6yFRu
LDJrDQiQxG/XSFq9yGBlp/4k3x2cFEAWgJibfumXuyDAVrZxRXrTn7lTcvODVJCz
Od7lot8Bxo9BvZC7TqHTkPX4VRZ+qv4+pwGnaTLUAi8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7600)
+gMHMaZHyDUCJLptkoSw3mHtJKjU678uOYh94xKeSJaimAWTpo5DD4KaFDhQ1pE8
Bh/V1YOrww9sfkoa78gM4OFAnr7HBLBxJr8DArzcVa6t0pqeh7R1AV4ZCwyjoMmc
8tEgwqu817A27DDwb4cdatIHDAo1dohU9LTd+Eu4nPSxGffTKRrC2fe2yjyyL16/
jZQ4VHxM0EFHIONJOkqYoYBHzYwhMEkJvUCFyQR6S+jsunLwHmKf2cZwS6eIfMAE
8Su9zYtyx/6t8WMBUGGXdPUNdFVUsKML7y4YMf4XZGXyA+2L3Jwn/sizgyfBUfLK
yF9ngOhWZBstfALqZV8w5+LFildxbRP1wOF4aEmXINPRmOJ4sPVjDXMy095y2JWO
TpVhMoML30O5Lpg5/F2cVhb/ydvepckMN6fdKfByQt3It+QWEMQkki3M4kIODcRr
ij3Aj527hweVG0LnKOZX0Jxn7aR9p+i7tkH7LgTcnyFM2Msz0b9dZlypcflIQYDy
Ml70r2ewx1xNhNlQpeCVwbtbTJz1f2COF+TWKHiVFOhFDCckHDso4F+iK1NTGMwc
xauQtjqndWGaE6kw8JufozL6tIQ592wwo+ZMk7P/MOkHG7T62p1ULzEyeoYfOYDQ
n3tdLitD8C+KBlN7rr/8qvRdGnYeEG6kXSJVaZumbO4KodBoLOFnddeI6+EgeO9R
XWqf6fV/qPVvt8pVLt4FyKZc1JZOxtEYJrvZNVSmmkTxAv88QqSWOjL+vpa9dAs8
pP7Un62LXUvg0yTgpZgJgxd9Fg1hUWHunjsVs28tw16eCoSQhFN9gGFuGlh5S355
/zYfAZswTFLsCZojbFWWJvrpan9zgdOvyqzQc98TiSQVd1rk1t/kAZ8PDYL2piuW
ZzMGO0WnHnx9gEQm7PqgL6Rc7uPjeO4mKCjlZaO0idNzJkzR/fX/6c56LWhCmCm0
GWn3qypGRPD9fq90cJMejn/AHB5wS2qEDZGcsMi0fznmEa81SagwecUeG8UvTyAd
QwKgACFwVj9x1EHR7TDzASca4IQR3fhPWASyLyLn6kKRFekVy6ZO/TnAa4A5mk4r
otrCs/5fGQorToSace23OBmOZREvnmv63pVHtJyPc9f+Wnkc41oy0O2lEvLzhidE
BbHQ/DBTZnolNTbH9b9oXTU1SE5M5sv6XOIALD26matJjDPaa4p6A9RrUCDEQP5y
N5QJY4nnPWjrTOxqyFdgKDSOQDIzBHeKZdarLgRVEoNG4gEJ0jmpkB2PZDbWOPht
ehL13OZuI6fx2M5Ojys9LqGIO7oyHIiQpiQTvoc+7Rr5U9WcnCJZuih4mKnaVEax
8dRD4e6FYnYVx7xH7WcRl5uyubX68LH0A0Kqy6pTDY8eOsBLRtm13En/iCPa1gEK
Ldmo38VVToOtvGefqTaLjO/1KzoWCJF2tQ/kI+xuJowYeU2RAI8YYjKNTgTk+fqs
LnEOLI5USeF0bh8m5i5EDom14610d4eLqtyjLMvndQJ7w8bQMyDx1mCX9Zr+hp4+
C5KZYElnLlxGHfOTjCEpNqlKkm5x40selLzqO3aG2i0XDZEztR4aStOyGq8SZ18j
pXZOI4kLARhDLpWEEEMDHOi7pA8SfMK/SSlOw8OyMcWb7dzE2si+LoHTZ3OTAH0I
XqD5Av24e81oKXhlpvm3+P1tIXjgnGcFYUvto2AmZ8cled1SUohUNyxi7Zzukmm/
uMJa3Nw9vHCCJLuXTdKot06uthaDrNE3Y1fn+qXgXI1l2ltKELdEF+coJP4p82FL
TgY4NlRrWZSJX7HhP3zB2KRXylPuFujGzF3CVs/J8oFGPCYnCJ1usujlnudBdF+W
3y4K+j/YZ67rqnkBbec3eauIQG7Yy3BpUGzSgGswSINtsvl+HokO/JLI7F/pyv5e
bY8hAJrWN3J0QlckrXNp0nF2bMF0ZMWW6wHxA+y4Gy226EN+KYteRKBFTaT87SNm
qUiDofvg6VxCJThz1RBEKTgjvnEcuS586MLIDy+JCQ/bQwdFSqLFWhq2AQEGqb0W
lOePiRZu/N+S6XbmRgcOjFtBRZpTQHjkql7d8pbHs8c22xA3vcgGq63i8Zm/qLae
prGIPep+o5F4QOahkYZeQhbpBvLiQQ0HZZb3iUbR42r5AQ/CeGJ6Sv3yCAz0UcVE
c5G18R8ujamM+q4/8W6gIQxB4TUOFsWtNGJK5SAdif57MF+SrqLEKmSewcFYCFx+
7EksLVJPBkVTbmvp5Z70+2WX/J449ddfR2aW+8X8QjWuiX2ulN/sln+3ZuEOhVQf
nZ20p9d8luNasy5d09tRa3wxKDEUY4bSL6r4gphBPiOmrtpT0QOWTgdnJ3TbF5J8
z4ksFbRocdUOOd83+WJhJPw5y2okg97e8Pbb47xjh8TJdxpHX1mfNTl7StN7ikYa
CiveasSrmcbnOimJwbspH7MXFguQ1nUh5EQUg0QpH3dWzVvjhwgh+MVmVt6ElvsY
c/LHUxwbL1nI3uD7xprGQKu+vGs+zUW3992m3t05SUG8BzLlxr3kte4ByfHbWRCl
YZk+44aE6JiPu4/R3qesubWaclgqYMWNGsRMIwRbu/H+a1FUzbKFBskGhRrHkEew
HWtUG4vB1cnDov4H9hupFSIqmm9gNHvhWYXiwVXUziYSSSZjXCK4kaZ5ku/ZL5sg
qMAwQcIk/a3jLmYZhQMQB17si3LgHhnY18m5gfEOKRJTPTmqOi5w/6Gg5/e8s0xp
ZObDohBRZPM/pzWpUKEkdKTjBhhzw8y0FhuJ74MLd8c2eiUO5Rf/alFHGyzH8kNJ
9Bx3sVsNScIr9jF9Wedd7d/njcb28WHXLoHmKrxPuiL2oR5dBOY7hH0wUMNK4AYN
uV6vh3QhMZFoxBIPbKaH6a4bnt0lUNAAveRqpjkp5WfqmkXXWpbTSYnLmVHqvFd7
3Jop/8PYDHleQSbUaAM/zjGUd8KG8xhtkJxhLhGXXGKMy5cGBD9/VoaMeG0lTjsq
AOLygzz61zaCCv1Jm6UbjVFUiavfv3bvDYW9kBmitagJJ6tlL9onJrN534xFAtV5
fctAPkWR8WrPMqW6LL5mOhOFybIjb1CyL6RcRPoJ9aPwn0QT/ER076mDFNhVNYph
/PXlTgByOOIBRvgk4ihH3ed41w+YfSDeyI7c/rYHZBv0I5OmwHyTGYxX/RAvkl7O
ayhOLKdvrxMcD2fRhIAlxZhBl2X4NRAuEVWpkjy4VCENupUm9QTQZk2yaGgiiuyB
57kBCynGGOQmpHN5pldrSBVSARITAz9t2Vue/lOygTMkMG0sf+q/xl7WDivY9hV6
9i3vRBbJS3ahy/3jlmOwj+uTJdFQH9v/AuCCBxCay5OqFB48KqOqGTnIEdIT7PlO
PNtqmY5Ucr32tTtzB95yS4E0rM4Z+zjcVYFGlNdZrJJTPm5c26CnHbsFjTalDqMr
MKoDD94kEGOOP5F/FLoJUdQpk4z6CoCCG8/w0iq0RLVBurdMCN1pOW8GHVTQg3yb
7YPkjH1ijB+bm6tpPs9fGS3LKMWLeWWgIoNd0VrC5COsnQHwExNc9vlFTaJHfB3J
5xDFEoRqsgwixbx2Vk6KLu6yudS38Z9W/FD5uS5ZbFaX63yKpg9yWW3f0hGcoFFu
B4kb1qldM8M8KZVeXQKboPkn+lT1JtZJOTxW54sYptTge6Cmr3u9XbbMfwibFBeJ
hOkDbmPt2OOnJKGyBQCBcMM30GaMRb8F/BA1ERR89v1hN7ZEzJOiseVkKd3oesH0
lmautGIargAXImbGWnSqMI5kmeSw4bl6ZKiI9D6zd4M30RePtiRFy4WOTrHYWjpd
wleSFkIgU3KwLMuy7nsyWUTksF3uE3clwf5nCJDoKsQVCuQlTJUTB8X3nmAMdCHI
6Q71T4x0cd0/cUdCQ/FwVSQ0sTOocLbEGFqt9ev2euYWzHquPoBq4E1EPZfJYEH8
HF2MtYOTreaZBIPzJbi8B0DBMljfm/H6JHHwV9F7zGSzMJdkgrSj9j2yjYa5ugvQ
tK4bymbHguhLRwDqQBndG1FHjCTTA2imM8vmFS78irRCnb5lVsd55cxs3h5kJB1t
B2BE4eJoLtw0J/9BxoYtU67jRIywsFu1eL/JOfGKTXOoxOtDeNxy4Y5wswP2YP52
3UnK7h5aJS316r3coi5HG+8kI0IFCw4pOdARbtmXhsMel3cIeGDLD+9+IfUlKL4P
LpxAW3MN1D88QKMwr2BRhUXbadGt2gQfTzgdErIJGfYZBcH072RJYu3yn3kIAL1F
XTeN7g+buYSeltJZs8XDBSeSsg4NgqBXwBhrRj6dkD/AEQuJCY/L2TmP/5XVqW5m
YPhwe9Xvq+9Jk6H+Gz1P6IE3wl5Za02B3vmn/r82jkKQZ0nZDQ8qnzCsgypPuA6S
VpT3muEuRYxZOabBK4J3VZ+dENor00WO71khATXOXLlUYBEHx98fVKnCt8Hx7Daw
bzUQ22sUFX7X5Q0DCEEjh7xLwUAXfiVYDafBJSer1mnNWd1wEVRFxzZXund09wc0
bKgEjvwKh4aQ0HDDz8Th6LCTV0tIdlu7dG9Vq/5MXrjZi1RTLkj3BYM84kJNJcx0
GOqiU6QSyOxuUmS3sp5oevDJuYV63MlAMIKWwGxVm174C6g0R+cYr5cKkTRYb3qN
xqL0EjKycV6BvKQNwwfjKtY9mDJu6Tm7zGQRLAKq5PfRWTU9CkpLRZDezn2thb3d
H7zJ1swcsDjTjQDIc49nnRTbBEiL/hm40uwOP1lEH4nNVLL31rhw6IW95UOmqUk6
DEIkOCdYKYUPg+v5yIViwJ2EBt6iNcibass+w78lcNyhfSZYhpLJSdZc9BuoD0G+
yDX2/kA4VKwrq9N6/QLdl+QUMRXoyfYEl1AP1vlvJsCd/xgbMdF5tDfMbN0RCs42
P4Vo/arXwDDWNG373ApiIbs9f1eHC7NwDICSWv13DL+n2zYIzuP6h2UHVBC372dK
oe6Vc7pbekxoQpVkjn8sF6Z3NJPAUzSYf79BgKTR6KwnAfKQy9dRBrHZ34W2iUHP
ByM+n8DfUWCwV2TKVezaA+JBhgfv9LUK9Qpqbl9LZx1V7lm69TEzvI4cMuFxA4Ym
W1M/A5F40EKk7TctKZj+gc7jQr7LfULoPXStq+yyFLiBXuJv0C3yke5lso8m0A+H
mlS1lEeZbrGnMld6kr9Aqyy8Sqzat/Q7KAJfldbu4p4Ed1YBRZttii8kpVJkAtCY
3RKC3S62GE7Y1mHLVY+BED7eQqtyhr/PKB6ng224tEmOch7qazPwMJyCU+4vSyOV
5x66LJZ24lQsUzr381esxmurGzgIJ09CHHtOqM3NBBhYF5gBbvYjdXP8IG36/ZKZ
7hGzDMPzhgD+LSJuTK3dOov8MSRSn3pPQzM0tynPqaSVLqh4/oC/Lf9dagNtMkCO
Lw9M31Q1SfLwbJgCooMoDJyrHfnXqxIRYJraFfzB16rHcTxEATw91+7ASN8+Ru2x
62xirWMx29hhbIUgrRj/rWYiukNHbqTS3p7TEfOCeIUuv/S9LlhNxP0CEsJ1Wkhr
fc4RsE132UeBBNapPt4wB8YQzJSKltH+zAtzphgMDbb2/2NtD3nW+lL+IzeJKlok
MEoL+QXufUtHp6xvs9nXOFsMqW1SRuw1gDP3TqSmZLzJr6vxZsiG363zIikuZWbD
vcCphKVdDw/800sBepVZen42HEojjLGgoEjUyNBG8o8EsncN07jeA+VuBu3rO7QD
hneRju1SpEtj1YOSYPJgOyVvXyTbnhunAsKpf46mU71onKAR96aE9ixxvXTenkIR
yvSaAaR5kbJ9xZcAhJ/JUQfLLMxM4rSCNsVKvk8wWaX7yD4qJSomwkC2PLBoIXu1
iPFVklLPwsjbtKn9Vs2YIhGimX9ysyBfo/97izC1/Mxi560uwYPn9wDijvwyMMTT
NYQTnfs1POJuvhc7N/6ieAeFBTZHuuqiUkKyh7JuPa9RNLQvh2DQEgN79lGnrgUS
oU+ciQ7sa+bWhm8hcGQ8nFd3Mju9c/Ezt1RoiwmgY7wwW3NoLeDvKygFdh7oylbd
H1ncfbo22Mu3nYFxkSkhEq36ZYSmwSanvjDr12k+PAHsrGheZq+U0s9PKZ1UP+w2
bzZUeKih5R16P/yF7nxLEJqF9a+4ZcHj7a6B1c+F1PuEE5NcQobgqsWv7YMUTbcU
G8AAZBcRgcLof7sDxyZYW5VF3l3C8hcJUuVe39fxbtE4bP9ygfGwH4Hsp4tw/jes
B1WmUMM8ay/AcDIhcJSFfi4y50Fw47/sQT/BYsktGZsV39Ym93C9UIfAwy7lh8jX
pqQXfrKaHGwNlOcmAhdW1Mv3RsBE4kFjirIaPCfiDzN/jEIBVIcFLQfVJUISPZeX
2UVOKUrSqdFtzDFs4VQN16lidzgVXpJ+GGYkm4uCA/UkL7DrfBTmVmqeka2RE9kL
ZilQ6dGuE4hekOZ+y0ON/8cH6CwmKhQm8WEE/EBP+UHF4hlJ/MQy+4DwiFrALBYE
RJ4eKECqErpthvdL28Z3G1r16w1Mz63+4KUwxZWB+KMbY91kRsMX0EYuKnBRkiP/
aSGvLXgKpswRw6/S1/sxwYy5BuBBHTdwNXCMt1hAsf9UAz+2WhJjr8yJnfTcB1J+
CEDj9p0HATbC9GtQLmANECA4dj907x4g5eyePI0keQ0V6YqAJ1WE7LtUIxl7wdC2
Qg9f7j8cQ3tBR3IpoWoOup5PAy+1WhcTdHdPtn5YFCRwnEC4cwtrHCETWa290BhG
DRfMLrsRmkHSIzBNYLp4wsXHraM8AgeJHx/1IwUzABH63BGLloPWYO4CRlkzXkR3
yckmO323fpNfWfBUe35Zbusv2UkPdM3aZ4JVarBSTvcLiVrSUgDO841ETm8xsz7h
qDR4/xR9XoNAAzAKSfj34MANjCqJOpPREJYLamB0wPVTks4emAdIwehMCQ5vcfF4
BkwNLgPHSJXHPO/mS18phHuMplQzP4avza4CGGR0/gWtVnspoNyXF7WrJM+Uywlq
mjNO3cbvnDdX93nctJOyF9808PDuD4wqFZbu0T+NFLb3eqipKHF8SxJe2Ity5BfQ
7Oa8Vr3JP7sJ5gOHyMdrOrsPP364DuwXI5Bx4vyAbvA0thQ5Ivjoa57eAXzMmzs9
HragxvRGCA8UdIiEXGP1GAFR4n0yMNiyNHxfmXg9hbFwdMTxGH9IXzAL4nPTt++5
ymy7VRVCqNWSKETcIbDnTYPt8Ibvleb8UNrM3+RZ5HrDo+Jvk7PaFFwMx6Xyr0uy
ctBIZGseDkVqWc3k41YvYzoOrLbR6T1k6mcOA1BWqvQjnu5ctoUGwa5X2UtrgDAC
CZlqOLYz+hz2NSxXO82JiaaFMK7t6aZhlSxy9yt8oYAluuki9VgL3SH0AsWd1JdB
w52r1LLf3wC4PlNKbW3fhLCQTqugMPMmYqMvfaFTe0uvSOUTBoyzzc7FU5vjs+wp
1QOjY3PBYg3pq9GpSPwzkY7QOv35I1Zhf5ycNhMU4KpeTFB+GAT5VsFVIQ1l6C+c
AnZ0kQGOfkRwVzLKrhTDPY+uQZhvIGpYZOMmNVDfv8qsqosjuvQt2PtKro3pIMYm
iiYlIvcDdUniYtzhjvIRlbXwNPIfRKTa+AaNYvMcdqR/i4QviSCAFgX10pW/ln6t
yOomTfZ6PxEVxBnXGQhlgOn2OGHknAopynQ5VjHQWttv9eLVhelcYn4xkd3jgT9m
sZbv9HrvsPvDHfxcxTtm/JKet5c59HHc7KGpTyufBmDEfwwTQqL0o0DJGtij7+dF
tZa68vH3IY5dsaxeVfUpY6/XYypX00e02ePZt7wPwP0yvs5+Q5vpr4ljZVWXTxgH
4Ln368jpfM/lKr4Re/B3s+qVPDkLBXutqhUiuNTgsah7I//mg5Fl7jS3Ozb/lzDR
rpGiFcvQumGlmes67B78lTOIr7mc9NR+7O1z3+R/i/JuvUjZInBOJe7be27zc1A0
f3fJo/sEjkYANRe4RP3/XaSnmQt0YAKaIgxZ2RqyktRYmp3ho2+qYo6ZrGNwTE+0
FHTv0tl4cdV9Ydb4zLfTIvBtB9g7hbAy49N5CQm3/Fx7gMZjaXbbQrMmr3lL6mA/
xPTtBBCdIa4PtmJ9m6jrihDbXrBVk7zZjdbupPGV1UdnxtE3uy8EtJeDecqHiVNd
D6LhjORW99lQe1e8VSs1Ho2iyLCGiXsc0HpKJr6GHv1FBiCIg3LEOItJfoD0O746
IsDrIP2KWE3yc7fIZeoKHsRxLIzwMHD2FNy61WFIOJK7Nlb0yQnabcxSU3kX5c7c
zZs1wymQESA2idPOD97AyGleo7IoLxHTRI/yTKWDfI33laDmmQ22m4foWIykVrt4
XsDbltAs5htr3Yik3L++SZxU1v+tcoAmAmZ4iBUE2YzpAqqVzz2hXbkpAZlsVmTP
Cr72Si0FS2/sIAVqzicCnslsqw5bHFRpNwLe3kAPn4dUx2TZhTSZf3FoMpLJLdbC
xlk7hJwduRaash8jMbVD97bcbsvq7NK6NKLxOTvc0nktOlLApvW6bWNLNmDtWBtQ
8mALyeI0LiBeewTjuH72PUJXwx5VLUa6MeucjZ92wp7UEWVWOUkwcTQABvnXcVmC
RnowbA4UDxdgDJVpxADV3fAgD69Pygd7z7x7puMZOkiacalytUYidTGtXz3YCHH+
HdOUrRjEFzoCW4KsFXhtfnqxEEBPWKQlwrKgeleZfiDRbyHJ4Dr30NOtQWg4+gEd
xVP2otllWbbrQurQVFjV4RZRMZstGeSC9dF6dKWmNR+X3xiUlX9UONYxRkcyJ4Vk
riGYaRDsMyB//00RDmtq5TVhhPG43cRZJ1CmQ6zZq5ftWaB0GCsmyaXn7O+c9lgg
SKqPhn1DCSPgfd144FN/krk7bT7iA1qhRLHkWQHzblEtUiv36HIYCGkclXcr0Ii6
KP1g9S1xvEqk9FhucmFfArAaqFe7uNySkYxm5tDfMStu5qjBkso52jWGQzVQN6dB
gSiP1Q0lpS05XERx8FI8hH+JILBt6Y7ZCf/uk6RK3lVVRPo3BrOcmWE84YdXs8bu
KknPfE78QqJ4VN/2urj93gGCKvCF9RoQ1FJRGvZYLmo4C/2e6NL0N4o4afdtktzS
ddFQvQPEkqAlrHWiC1r3H1F1jOVAldDLHGE+eM1GR6rlHNsphgsCmmhO5c6CkS0G
EpWzzrVXWrlXP8JznqA2DX24r958kBzOc+TREuUloB10g78jckkJvA+aF4qmJ5z9
ob6+CLMpXT5d4BHsIPRUDRLcuOkU9c7i67tQSszPPtlXI7H2YhEEwhTcBCk5zufL
wyFHJNyQ8o1f1DuYwMks9W16ih2BFbohnGG1CJZIQe5+z0HOIZE4IurIggQupc7v
hOzfTxmrPl0PK5kPh9dC4xIK9DkrCiLo3hvZKBBucOpkRs4YktczvqeSAtKwpLEW
ZeFPiKijz+6wuvd/VpeMtFN9LcqYNPZiZx4cN00aF34wUiKhB8MN+ziPAVXUSIdi
1jLYcPloQSYMoiUdY9DW4ahlnMFU/YG/eqBvNFXz1B2BObKV6YIE9eTrG6O0sbMv
YsjpcWRxx5kOanuCakzPzfGeu9U1eTAMXEYvKNT63pWeEC3reONaHwhVy+mYkfWW
gzjFkF/SlthUr9LmdCQG7GROQhd1tw34KBAEkTAhsMFWZgokENWKQlr7+7AnGb15
6ca8LAMPcUPvysh9GGNaSvMcSyLXOS0eKZ/Go7Ew2/aFiz4hUFR9iWpadMrPnv7h
K+YvbbbBwE5xOP6wrq4KBupt3/eXiiVJeYv7vl/wodjGJfgVgkVl066F4GFlI7g4
NfHns7bN48mzVkP8ZfMH+65PGVn4Ymd8N3WQoiFcNFx7q0mvRji8tfXrTF+2WW3K
+v+Q3Du9dJp5LrFn96d+XepKdxiYwe45/ICvxt2FKGffkv2JPvs/UzHBFS2sZNJV
cFLfivxqaTBEgh9t4Vp/jWrB8b09hNJRxt+XGKiDUFwrRhvTDO1yaXjzquvHKHkU
3xWbghH6t+qc0M65yoE9/7nEnTgLkpGCiZehhOmidQ0WW/3k3zwuuiIgdUI4FDlx
qMw5yt3rrGYpYLCwvzrGRA==
`pragma protect end_protected
