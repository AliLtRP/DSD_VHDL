// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Hv+Xf9wW8JBxwdIGbkMnaMxbz1b2gI5fSwYUw7/4JdiP5moOeNx6jQpEbVaLXDZKUamfpp7Wdral
2uaMHgZBNpuzyYowf/OuaIo+NH9OgUbDv1C1bzuInTmy7A5jSPRijX5lZngZ1KgDzwK8UwQBgI9A
eX5SL8sc9OODVWrXhtz89D3688yv7Nc/JSIJBPG2fMj9kGFoafvtX4B2e70u2I1PH8JAokhhtDRG
SNGUSmfl3IpUtYZGtvy/RzpAjeQmgF2HAX4pO0SK4bKhcS+h+WmIiVZQsxHvJXDTHQAcJNi6SMFS
g/kHEldKzwQjSE76ZHIP1mT/NaScrV/dwcRa6g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
udITNF7mxPbPTmvtfx0alz6liwstdobWYT1aqs231fUu18TD4JxrsfCOj/c3GzNRq+kJWnvysDPG
B49JgjElKq0Tztv6AiuoN8AcYFhDQoqfUX/WudnilUKpGe1kh/7tDJgx0TZK9ljt7Fy/ynFG4r61
4fNTvdFXXz1/nTPjpVLAgLxUvbXRqYx3rNlFf2JEzdYARssiekVtQfqX6YmNOHXusnozVD2Ehano
RKg8vSMk4ExhUf9oUivzAxcmfN0LCLrR6ecD88gt/z8MjGckkDwRVFIEoeCblIg0vwlMIlGvv4GS
kOYApEMC+Rmqfkkc/C56a6e//B/+GhP2Pr48IZr982VuAPYuBcbW0uSTwUDqkrQSk4IcvEe29OTQ
HJs23inADq29zWEpGRWUKixvW7IgHgnSTvzZBhNpEb9zWloH6JPpz1qfO4Vdk5LMYDmX7hfo+yMA
UjUvmER+QBD9UNvQGW0FpAf0c0RjUxJRX/K1HkIH9KgV+5Tjlqp6jFIf8K08eeurSHYurXih8Q6/
gAaKWpqZjM0dhKQerip/k7tbgDVkms1+KQb7R1p4fp2DBdSnsxSblOUczAIJNCnKNePsx9gtE6RD
izx3ekg312DQhBhZgB7ROwpzZ/pS2hcZWStqHih528dKY7CCnFm13uRXP50icB1bPlnXqPA0OWm3
wu5tWkyLGhvvovFx3SnPQLOBj+HA/VF6NTYoVWhOXuQgMVqhN7Drlkzm3F3IecMUDf02SGtEl8dB
NzlG3yCbT4G31SREizGE4hE2QG1LCpY8x0TryejoMALR1JnlX/IozmR+PaM1Wz3k9fNltRVoZxVk
16VHj/VmYWnF0ov5BbNZNkC4CQggM5l7Gt+qQH1sinbbzG03f1Rsf7AR8Dezed76Vu6kQPjMNUMZ
fmOwYbsGN1tZes0ub4/KCm+kR88mbe2sWvvkMf0bHGDZ68EjGSKAzcrzDs3vVgY5PzzPdvXkDXJu
HOODqUP3Du4DvCAQP8+pfA+JJN6ONjLTqIQW0p3YsmcuvDW9Ov/LPiJULk8/HkmNfVkDWnTLxlxC
S2nlR1Rz8mO6HSe3uyBrVzuFR/t3Oh0ilFBvc+3Lb4hhzP72lu6jVu6w0NQLzZfWzoRV7yvi03f9
E65DLqkwE0qIzaNR92MM//bFbkEzvDDNZGweoSQdWQc00mTsi9/tDIxBLVBLfPb0O2zDZKfyA0ny
HEYjCtC0FoOUhDwrzRTUBFaFfGh5uGuKiRqIbBIA2oDFaboePh99aZL3S8Gn8REdwIFxzbU4hz7x
+JucA/ekOEHUrKZcE2xzOsXCtifoNMWqbhYhWVnMwnGfeIxFWQWLJe8EQcKBTAvNFE5rwRZyt/C8
aJ53PH4j4xwQTB/1fz9mOpqGl2l8CrTD6Fwjdsr8FjbghkHqUicH52r5oKj1TzAEoX2+4Aph9Zoc
esi1aEZBM1a0j3RG7HPcO/rvo79lfHQmCu5Ha+8H6nwY/3Q3ZKjKXbGia/hN9WAxvTrZLOTqSlqW
f0ghl7hti1pbQnF7SoW6Mmohp581cyKajQAlmmaL0iBOWM4zfzmAaXrTwjXiIFFaMw3/03mWne+H
MlqSy4N5Vxg5ftVcJnyZfYYGLDnWScuc27TtatKnMW2xmnV2sNtttrszp57yxkfaooTlitOlyN7y
uQ/Vl8GFfwQcbXU+T4GypOwsVlCgSFkQbrX/Natf9Pph4nw6f9TgPTcvxXO1/P/7Pa2rX9XqoWoY
9fdl3ZhKInXPnZ8Q7f3BVfBH8SnTAitnjA/wzYau0u3tJ0j6TfHEYwkMrKLYG6pMbyjlaJHesctM
LUhcHcsSVVhYMhc6Kgcy3lJ8m9yiVZfm+A+8Uu4eo/N1OaCaxku/QL1Ia4PbMlUyhxxBZ6ZGYWTP
Re38PaGUV87l6jmMv34mIshv17hYim+0y/MxrGzjToLE7tPx+AB9y5uHnXtlVE83xEp9JRanIlID
ptuXJ3UUx/thhomRktg6oPy3/v7rUJ+LLwgIc66aSr6S8si1XXhb91BEuP6DaV5YOPzGFF1/3uXW
SinFqDL6ZHHI17NA2RR/K2+YX5jM1k3HovT9Z7Y0Ipl8KzNjaYV/wAziot3oeVDaIXJCcwVpXrgK
KZ8/GYICHE074tbw3cvvUvZVI7e8pDRN4FV2tfwBQ3QSwkaMT9JtJRlVVhu8XkujMF05KjJJ5xoF
owZhWHwEEiF+H48aW2ZYGW0Fhi5khk4ZVE17hwxIilkrHj/60/gZHqkEw7dSUhaKHR2HG6MIleyb
xNJFiGrpx3jFyJ487O8+gL+uvExUBHeUnhAMWVZSq00AD/jge/ceMb2RQTkhboOr9ty/GR6gSphT
KLWDJBCjjlJWbkN8h0asqY0KLgLO/7xR/n0MoHw3xrd2i6yGYTUJLWtd08dK0wuKUbul8Y1yeGVy
oizOLw+cSvmXbZkutv/DzbyieWnN5W7hx+8vsdKx1WxVFHTN3GdWyKgBOLJMCjogJc8nzesONOTr
Z9pswdJL7LgcfBo1XTh/r2EDwCUgbaDj//rf/sH43zcoDo3cu7ri6QEbGpwoDH3PTzb+z8I0oRjA
H5WGxaTGAPh19gtT2qogB7ieqEpSlnG/88Gc69slxEXlglBUgpUPkd7kIX5OVYFd24z8WXrHI0CE
vjagXVBXIwyKXZwDxHkS+6+6uSNovpMOfAWOwUqmnhtp6b92n6vwg1ptBuFxRJVf8wdZG4T01lOH
P9tdnCWb0E06wGeiJ2dLSHBFhj18Ac5SRp1AfPkmQHXWy5VSyf8xlwcWZqTIyCihD6jNY8+IzV3m
C+dIPnRy9/qRl0Rr7EEkRLHqgudgki73ZEMfXArVNuWagJZr8iY+0e3qGiAV685pKNp1FBvUjb/o
1n0sPHWGT/8WmqGam+BvsUGLrtzlDNyB31AEMbzmVRf/odwbadQHBV2KHEwPwBvpAL7u9d4Myj1J
BjFcujQJZry57FLWzKt4b9jIaJH1WWOFp5xS0ZKZ8faAY3M/hL5e+xiue7qmxzbNiRfuWVdb4jqd
NydXeyBweX3KULoLyAZU7mnfqIKQrjs61uuKif77FYHQUJP9+LKhmWsg6DY5Twu+9ux0eMpt2m5W
9EOhZSjJF3YvZeBT/67RC7x06JkQ57g4U3Kmg574i/QEg69HPpKxi9WBEWE/8luy/w+fFVeIAtPh
uXCSmgQo+RSJWawDE4kmQrtZyv6xCu+hdOndd1EKlKhN+8YP/Bk2xY2KQNJZz+V4J5TS/IFwjwpa
R3Aa8M9otdyWxjc3vueyy4n8ulktSuxd9OKnfNFFMONmsXcOm5uaUmwYnF0W5SwyVBOeUmpZI1Dz
bb05id3quACFQp9RFDawyj1Lx8RAbBuzpNCBDNfhV6sgGSDYmv7DIxSNnfzJ2l2eYzQFQNP0+O/e
9e5287GAqIVuxzhO1WIM+YrG7afQVtU9eolOgu7sULFVmucHIdr1NFVVymYh8dRv/ggiyWa2tSQt
bfNNl+jL+P8WZjgJhN4wp/FYepT5TiREM+I/UCNM5Z8jLkT8uVIOVTbedYKCOOJ6Poe5UmkwqJZT
qyhivc05db8JLdVygyFYFP3U897E+RWkvadrA/ObCcRpl5qdOY+B8A1SKJWMdXWvms/7tyrz8hMo
KdEiIcWsWngmwz4JeS7eOBU0lK+OgK0o3k3bGkwgO9hfG6XRngXmpxH9vGFdzwo28JKBoZNFMkRZ
yNQNDHOuCowcJ5D2EAfTxpoZ4p2cJCkHZWRVOCn8DF9PMRofG4V73cCZc1sg1ic3/jCT50mqn1ku
Bm0Q2+qyTXbJA8vUdX5j1OvaHMNRCLGLIixB1oQWAfpT7QKw0+gzyTuBSxWjx4IfcC+oAJFhubtL
qgPVC5kWWPAr2FXnXZBrN38OJDIvfjXjkliP6V7U1tjm5goVIAaiCia3jGLfZQPc/SkbJbPJVplX
NKgujcnZPeBNP1KoBWj7zhuWKCRyGglAVLkurxe1H8TQkrNoNRZcPqF2uYZfG8hIe/TlNuirt/gA
vXjD0SP18niC5dspdi5bliU5oBPqwPJF9w9rwF+4wB+r7u15gd0tt+ot5dei4IP/s0S9CPYaRTft
NvyK+LgiHzHhd0+AxMqrclovg45Fn64eeZKUCJkH4CFbktxuOgFnER6dzmw2Z/q0h/9Euw15Zyy7
Ke+ebFeWOvx5AmmsByEcsq8cL9KQnG6yVvIRAakfEQazn0GvG2VVRCEdvRYOlrplT1JuEpzRQjCD
9b++kbhsqaDgtEeLuKU+ZWrcFj35BwhOtUAGQqzwzyXGhoyNbH6qfFgNj88K7QJG0F5wc65HmEjJ
FvRUcWXTPsXP4JJDDAdkOq4n7BLLefe0WyrslzfKUcyi/I2/9e+yb+jssL4rnhyJyw67C8os5JuL
Y2PKv915/qO1ztGNjRzqOmofKVsITA9znEaJ8hvDLtKEwxk//CT6uD1oGGLQixNSe5Q2P8S31r89
mLbAQtm49xzKrN5CG3ecgmkhZgzOt+8OdfrMN4+6832QWeFBeKry317Bxw6dEal87cX7t4DNAn2J
KFgVj+klTSYz2WjxDvDqCpjxni6vJrJUtwAxloK6Y4cEXOCBEub9W9VPuujPLCKeiPUAjmG9LR6T
MZWbZ4TV/2vpXYZEWzQQAiw+DVXNdr4FaXwNcQ7O1IlZeX7dCSo9w1oWSQfutuvb5rjFGiQYAYSs
XwKgIddLgW6euypt5E1IWWiRZG3BgYD7IDfnPlKjf6geTG2iJrkWW1MDNc3xleVY6JlID60Mm+9w
zbFmqsdeNE36u5VLMuO3mfACO4Enbe6WIOHvv3JEXenf+4Avbum0WdmHOc04tOSF8XPdoc2IzAVW
1reSLkh4/cpDqZu1rR9M9uGCnU3pM5MqV3p4UKzwhgBItUOcz/wEGZ5QVBK4bcwq3/O0Kt4yxoyz
sf+wSzZsYWrClXN2TARvGeRHLCCXOrxei4uA85LzyolAYftekBNaWKr/Cbd+nxSEWc1QX1tqzyoF
/ecPyHcTwuJ0WX0tarmXwK2Y4742DfWuz4Itmnw6LtJQiYJYzKlmXd+QsdA+7bSX1pOxtrFhzwUM
zYaj3ILXWGoUxA1iKYPlkGoogo22BTlcb/NWS4hyRr/gzBL6SuUN6ZxzSiAxQun4hCP5y1W+znXV
yqkVxyvW70QGSHQ5JfdYeRLhgNxSqr/yxzcJfQLymQycf8eOO8z3j2CTGIj3/cxaeTBIBmSIpu2K
ELR9A7LwN8wHlRRtvQSYvqqsooVRvNybTgIXHChnzqGipf1MBVSQYHmVB+mhxxL2Vk7YjwGIT+VV
AUHe6sTBLFgCAAyf6Zp8cXuBf/BBPkS+rqFyJVFngfcLzrWwc+bcJ0CI2P48/yKnC34nhTz9sxY8
N6rwWaAO/kDqalP+T5teT4VAUUIyV/4tnodovQsLLVLqoXgyaCGL1IXWglo75lzG5+3VAeg6nZzH
mMsq1hM9y62bXHeWrEhU2C1Y1aE0K2frZiFiuzOc8X9+FvWYw1MR/rlRihBOazXOYPXvMC7S2QzX
l0e0vfjBnZwLDO6oUTovWJHdRULWm6WnL78fTGQzwbdge71ZA2r9JRbg0kvcV2CM+LpibhxPIfX8
M26jUwDYCdI1XBU7+ByD4/Pw6L9tZ5Js5o/JZj5QfrAmhqqbepbbOVUHfVki7HyKAUaOGS+Ox4rs
MMWodTSwA60jaG894ebDlum0+gIFNXTGBAxVfg6+WkN32qmdD9NiRJprWCSs7mVTUhY1ekUuhWNl
elLVySQ0W8fd1fqT6vCi/xqH1NrEsaPRXS9VzgLBlRBCcAS67I191IzPTkgM0DuZCI1kThMklfSA
1zWxfzs+pSUIJc30stiUaRD6OoClP8PRlUNZxKRrmDFmPx+rrNYIPLHSmSuLmOp4W4HpPEBEXPar
EZNPhqjoHBNdgwgX0GTSG+NxNkFrfnFd0qUovi4ZzS6teBbnzcF7hpeXfLH/kDsmTqKz2pW59PpJ
FdtZMuHO7HOYvIpTe0jrD7Tv6F3Q2buwooN3dYdcGXa9/KzCEcUWpkHkZswILZzQIyntfW0+AvPx
EaGksxronccbhQyiurpj/UnP9uL0jz8QV5N2plwU7bAVe03IOPtShUHFC+MfOJ8r8u02F+1vTUGr
18Xuw0gaFtKy8dmgswAfey6UJt/kv3XHW/023IeNgp90NERWt2zjcQwqt5yJOa/gdpq8TSx/8NLX
EI7cnCIlaAZWKOKE9oRWA5CxtjeHN1ELc3AkPwYzNugrD3j6AmLrxC3GHdljJAJ2dDgLBdEc9TZO
JyFBvh0B5i7Pw2oKFr3DXOWtyKSrigIx6nuRqqhRLJoNJx/y9wLLfaxGQbElAZgNTHiPZzEPjlEq
J33oAp6ANAwMI//SLsN1KqTtVH+mAHfUN14bpT3IiKdzoiV3SBdiHDCNDN0q71Ynbrm/NDR+vv1W
q9UBnACLVHXmw/TfW8tSGnZNT12BRabpeUyw7j012M4iTVBB9pvbnxXSBt5NvbNEjiaIiqAP426q
LeF0HeGtwDmQDTbd2pI3pFgwKZ2FQ9ng40Pjs8OoAmYAz5UX2GzxGcI1mYvNWG4yqBGcNmZLEpM1
DZ1NBJE40xEhmdddUoDyOeKGfS3axoAEHrxt5v3H2+0q4dG7t7ttRMYZz+T0vlinSriUapg6fzGQ
KbBLAx9TRbdWoYjm6YmCouToZ6OcU4yMjySPR6ayi85SlfnLa1NjfYHXcHEP/778JcBOivEuraGx
VlNAG91hYwxCvJLYBxBOjDg1WOcfsah70I17Y+3HY0UKRXOuOpIT9qtxSb3IYXepTmYUgBEpz722
FqRSacGXS81v8LMExOcopAV4jzSBbtNX+HcBBNWbF842XTl+gnbPyjngalrPCB4SKkq0OVbweCtc
ps4zAUQzDM8ncfZNfRlP9jGCTdr9KcYhAnYnamWLsStX+LAYD4wWQG7flFPzW+Vu3jCPw6ythysE
1NvBWg/omvIJwy2OnXY9fZzBaB5k34gjD/jGcHW4pBpjey1O2MsOj+PCUtPniP5aqoPVVOCRrY9R
681YHoZTS5qhGfGHPmmk21VYlDAvWFNc86YpL66lsgdN4wd9h7xTD4F7m9ZkuzoA4Vs72nDzX9Lo
5dx1/05/whoFLeHoxM0j82wX3gxK1sEkfUiW24Cb8WvtCuzoOT+Zm7rbjF+1FtAX2Br0WoujccO9
wPaWXsbLwCkp2tEz4UQqS+TCuTXBG3iDfvptxH55C4eVQpQ4l1Qmd8CYAZDJg7oxfIzD1BLfOPAR
JDWzbhNZdR6FX31gzBpk/cYnDN2KolKkQFlgwI3kAv09n4fJbrJ67WXUvDCQ4j7v/wZ9+H98dSj2
sLJr0+255jss7gpIqrPzuByZX57ulAX3q28lzR2hrZRD3cDW9x5Yq2nkegonoslB2aqWQTcaQog/
1JWuQF74OjD+hhQz71WlfOIbWmJ4q4H7TgiZxGjvRYeaQuu8RPCmGRRqM4UcNWZWNet/WKZjdWj9
+woQ2rlenj0DPVfMu8dPf+o5BixOUTXaucLT+rQppEg7g4Jy3tnLmPII1YkjP4DgUCs9jAieyozh
GOrLRwnn2/9nDhc/4I1IWTt1cehDguNnkwn4FQxosflNmgXAS/Ht7gEi8p0R/en3e1FkqItH+QKS
LsKa4q3wUZMMt60DwiSJyrvKD5yR/xy065x/i7cv7y+7tUzsI/XrUtt8hCP6xBG3VrZ4ibCFcpwy
FS0Re478+rArtfeztkHFvncJYoNyqW1iUTPSlFryuzoASIrFzHg9S+I3P+5BJdFQ1BD3FiLrBjEO
qJkXRCqiTm3+zXPkfR5peiRuhqQKJvnVmq+FqVgodyoeqMpKQ4wZVxdaQdokgFR2rWxBXXiHaif3
Xh7aMl7ZktFJqJbQTjWp9uyVC4uX57rdJG/Vb9Lf6pOmCu/MA1mXSdLLOWOZlnC2wCk+Ayg8NZpg
SLeEv0aOGFr/dBBHezTS25DKii1bxDUCR7huzthJzix66ZPzR6ST+8dXZxZG1CQFENrdneJD4z5J
RyVtsj8o+zQpVQTfbA5ocEpoLeVlX2JvylTz+VVSSRsDADDvSEKTILS+YALmdjuKxGiN9xAfsicp
2AAtC9SedgwdmLeFj13bL3fTYU7FTHSUFQyQLEw4b1CBzRfFDFXKzTLxcsu0e9x/pQHFePJWA/Ig
Il04/JO1nRu5eycRg6DDJ2ajc/UTxfuGBuSEqz9ioI8eNMDPB/r0ppoj/7/Kr3y0l3dl+1VhSB0m
MGMFdzAPW+bCwdIk1FeFhZEkUyD9IN12IkL7MrzA0O03x6NOQQ2dW5yPZuk3FH6Hl/Rzj9JQ4JNR
YwiXUGbq2GWqqD4K4KvTimCyQAXpFDExQiDxcHJ6DY7aIXob94PczSgybB0oGckdNjT8k8ImOZus
Tcljzq3n6z56qU9DLPeyIfkXy0qYxDz32RK+b+H78Xe4bBE/ULzaSfu4nafAkxqtdWjuafPzhvNR
n4HN3tJh/IvcKUGVJRPWe+tvweSSzHKELM6AMB6D25OMtzTnIF+rn5rakkMCfCvFsaylYZPeYE+u
YyJUpn4J89vlKc09alLdomV79B6cZDtJZvNocrR5J9WKIvCk58N2yAKlsle2D9ZJEs6UxrbR4p/5
4C0d/9QNqrBD1k/pXXvEbIaTVesT0x1XNxMVEbnOsU65/H+95S0InQH44CoJ8hVqDRpr7WerFWI5
J0Y66Gs47P++O+tNmWYiGXQT0e3HHHYCbpv4PvfQITdMlJs8Ka0z7y+EosqjkBZ371blqNtcINjQ
eNVL5/sctUCo9VhqYoQw4ejJdv2HbU9cDMTTPe7QDqwSP03hiMMziOqsBOWbjw+3/NGz7vT/bGNW
47texNNSyXRJTu9DWb4ygKR9vsG1lyZ3AoUunUdw1zyV8aLNAaC2HGnu5APr1QrQ3imwm5qY7mIt
tQWEJJiEmVMnZixDvUF6Obnqg2VPNDjaOPDjUAuMdUtTqo+xAeNtMdAK9nfTBSQCHp53ETmy+CFa
l+HsTYu6E1sGY2GS0BKsgPagW8FPmOgLQSuyjRHKu1bwZUZy41o7au0H75hnkq2mqLX7kkeJYse3
RLpS4qSfu3lqEwPCeRuLoFtyBDJUGhWcNGEaUImq9vkBHuJ+dwnGvJpTOIJvDu91m0tUO+IHoeoi
EJguMFpr07IJKJkrEXyBwd4jK7iHw/qQc3BEtefzWPtsVIZivqGIFQriB4swU+ioYA5Gf/MGs777
sHxIBWAv4FU/Q38BysG6xa3y65VBoWDO1J0Lg/hHXr20gxkbkYY/J7HdFLktnK6+2TJCUAt60u5e
j5mnshabf7mmIk3HjG6kEG3eFrDvZIwLMTkAD8Qk/rScBipnEyEga51baSc29jzXgzsye7vE08Ly
kJAdrC52uaajTTFbwgxlhosls2n92UHYXxHo7XQpKVCQfgzZVf+Y8ODzcUxaMUrnHGJ7yrGeug1u
HO9/5V80GXzl8XA8Av712imsXcVWeqDucTop+JAtflpffqtIOGSLZ80GO5NP4rDjbG7kKm7mm6df
kUgZ7BfAxrCjjroA7AbTe0/4RlI0v07a6btmZ1tLV1P57DJDVjb+HVr9W+jthNsyx/n6IPgrPK26
b862HH7aAvb4BgE4S8fQhyPwb1dJeGl/dlbt2gq20VqfJhAwHqiBiTsJaSsy4C+gZIEuaOo/2kFh
sxcvrF61Jf4vcjSUj2rGJ8Hm6Kdbp6YIxkDGUbHPVcxbCzwZvdufkALsfXkXvJGrFFTLt3S2865v
11VamNDtxcYPQ1BXtRM45FPgCP4xIs4sxzyNB8BrIKJIjKWq+XCzvmIlrh+8Vb9rTQc5hXWMCgrT
Gb2MxpMezHxO2T7HVrAKumYTA0WavXPZkUyiI/qEqbjhj4Y4e4+/SX+/lD9b8p5bmnIy2L6avjKb
ygt2H34ELQG35mH0FO3FNEXTFSCSUD1rhkWNQU22uJ3jPE00qS0XCdPvak8M3bUisU6LINHSuZUP
3O9A90aUC+9wqDD+fb4CyOVJe4KYUvzoDIg/OWBBW67/v/YuojeHH6aqmWfDMIs6XuVaEtspYhi/
pSu/0dx+amG0rl72SNojOnspaekOAGakwmHZj568CHgIAiwT5DpBr7KVJd0yOUNFaJ3mrgXPBz1R
mqqDVMoh5PPgeazbghA8xVOD9ACcV1clORtT69IC+6TNg7nHid/WAQlrMRRWjQacIYgZ2q909zjP
B35YtCH1oZ6WUt8jWWMVg7Wft3FxaUuc8nafdeXKT6Z+7iL9CFk1BXZEYHbhL+KmPL7nlUKYYoSf
wPcvyZCx158eAdUvdbKM0qLYvhmrhPXjwVW73Dq0QQpT5mmEHMYNpiDjKNkl/oZXtCJzbGIpeB77
TI6/Qecl0GJjTKWDj/vslepi6UXmGZZfU8Vv6ORsfiW0ec2awQ+1JNtXYKcPL85IBulkChwN89MY
h3vKRmlbLkwW9wIxR01mxHf5g1Oul9q7H1ihxcD83L6YyvsLl1WjHkbNrCSHqDalTQ611JAlCy4X
HLqApC2G7qEnV0+sh7EomnvDA5oUKaYmtzdovUDV/ZP8gbCEW77kMM4r2LzVc9zWfDLbu/94CJ0d
EcnLIldpc8j9kKsUtmx/DcHOiKD/a+biBeyRXtQfLcbix1V0ixglaKnR9H6egm+RQitNkNjySl5n
oub8oYqxg4Zp/rvPHLCFN3rIr0qs0bEmlKDxaTnOd5D+8DgCXUQYDgwO6952cD7FfWsjdrovyCNZ
wrBk+ClR8GUgJ9eWLxW7DkTUZCuF1FA0KbXmsSIomAc6X4tNAdcbC/erts5jM7CmvWArIIVv4zwD
NzJIlq/x3cvODeQM2IDtx8S/qm6RxHaNhTfY4UQyeC9fFiXPlAa2we8JLxlSv7mJTvoE29zeChtk
N8Tlo8WOFYwntPnbHAzY/SwlAR9DMr2cMrE1OSWFMSvrfxKi4eZXULKWnGw0EqbpGs4+ediArLy5
VUaoVGKeNwg1RI06vmh0L4QhJ6GyWfaSIDgD4WwGLsMbPo9B6HA0sk8Uo2Mbl16hPiBqNt8/2RLj
hszy6JC8KPVDAKx1pNw5kKyy3tXHKVt2q5N8h1tGCiGd5CR0DVbRgmCZ2h62sE1epl+L3vSnFf0b
LEQXRygVWwdDfyvO93MA92E74E/Qm6DVz7NcGOqXzJ5Gghv3GGF+M8Ge/OVurUG2wX7jGmj3wSFK
w4GsxuI6BaK9ZqjEgVq9kxr1Gn4o9/Mi/tQkl8DdBBRwduNGbftH2s17Jgh+8f4QUCbkbMSadx/f
w5xredL6X8qcjjnRtiwa37/ndhNhOtzapQH4Lk49FRZEddG2hAY9t99YjLEj8ZFr10U3bc52Ypl/
TnKjsHBqjQYt9iX7//JBE4cAQQ+S9AK52IUheHPka78v7gwByouuDTJ05w5wooeJGqqOBu/z2Ohg
+sI9O+tSd7yfNGy0bxNbWXTG4rTPCVoaHCwEfR6mMOts2Qk62cy+qnHfXuMW7FeJcnef/39yLrix
VfqWjIez32CjKgN0fomeZG2Uy7XAL2I/YlXhXHXDNBgnWsu6o8QsOxnh+DNzMu57RyF2c3qgFuIA
4O2cTB/cYcra2MrzhLNoYZlHxR0x6UpSd9PlLCK32oY1fgSSHgXjrxiBREJS++Ka3Zr1IrCA6IOr
oUztQwfS7DpltTrwGLjTZjMScmPv1rNVyYP2DH/hrVJ/ge6Ui9ZSQ0xn6a4C0rARZqs4qlV27pMp
L+R93G7j2i7VVc44mdB0342pqqbkK3WMYpxIGFzKR03B7GfvUQtf3Bl22Lqk2f/CyAE1SzEccKBs
FbDC0DyAtRRCEJTn3gN1kgsoJvIRaus7aq2isPbltXWUobAMZayigUg69DchkNIqzfTs+x7Ypuiw
d+//IvC9sQyc8omoJ8vxsXxd6MmcePm9hMaq+LyODF55eoNh8Et2AP4xwhc3Lo0ZRik1ZhzNN0ov
5ZOyTg4GiZAWuwr2bpI/YrrHgxU6jkTUCeZApH8WW9v3HT6CTc9jjfyaLpDaoHxKZGoo5ATS6V4c
cF1Hl61HcJEYWjo6mcQmjjowmiQ8YqKMeY62OWk69EgFsuJZ3JaibDtDMAcTVQlgmFvRAXswXFkp
+vmtPh/waY0sVqEJZp5k1fcFAEyC5HPtu7eaGwUl6Hzh0Jfy7RRfc7+WJ7n79fWxgcAHRf07rY1n
nOdFlGtTzFAz2RB2ZQklY394hS0FgsvmjVMf9nxi0YIi/qvseJ8iiU9CwqfDVhHbBa84pJDNcEhY
9RGVQ8RUf+ovK4umHLZtTvWD/BO49MeZMyxvk3Vbs/vJSLkfx/h48abg8SD4mZ/yG4ujDZjjlOLY
XLPNIQt5xu4NkxAnmEVBVrY+rWOHO3OiGvIetYpsowLiutdDv5ZGUGGCtnVnkJqJ1M0UXrEOicnQ
XfDn3j6ZtzJbOUw9/X4biYGX3cKHZ6jDFVjIjsYoWXh9pz5Z1JgAVsNT0i3LzIOGHpfd0Hc0qTmM
X/0GYlccJgFGHmnIVp4MuQT7/01CBdbmThmFeELNskgTlV222+4+d8Um0+/JB+GT/8lGcya/RElh
JNfvgwAXc1DJGmKJ0yU/hQju+/As6oK7GGrX06HSq8SbAqd9UAznpqJq++xWo8NA2ZUxXqmjPVAY
k90/G6zWSF5cGsga1+xvZwiYedhbgr/qlulDklNxs1WkghqvIC0KxWZ8JvQ6KByZFy7e/8nBLS2N
IZ+L4a50LbWKCe0d8S8CdjmgwDGaDFXvGmoonLfiKv1axvznCW58hRFfPV15nKfAmw7/fGRqXvI9
quK0Bqekf51KJhDQxlwtsZ/hbbQABdg8YHU450XBz7LtB3ShBpSaRRTaXW/5VYzuLziDzYrAfkvN
MGBV9GgLDJUKsY0anEi6Qd9uy2Z8DwiA6AnmK87y2SCohY8Ad8RCCQ8NOVoKth7NFLQVsB2agOQ/
q3r9Ioaq6lIGsC7xncgChDKI2leJkq90hH5ocGHqzbfGwlR9i+uxBufyGbRxlXzmg9MDcjLoO4jl
Z4jTEubXLhorsTQXJtFzKmAuYkPdPJNb6oPxc0+CpPOvcSJwiEN7JeCpz4JkNxzrO9JJHr3TOOwA
a1t7/NqzFiIWetiqs9HIBKhYMmzDcV79s9my6dCkP62dlCNAtIhcjVGZ3hqQAjo+3yFG6z1KhIOR
8wvsKl+5MnEdL9NVaTTzXyyhsL2fvMb6fwah8YkRgu1NIHFyl0+GDjHD3HBwLvHoEk+8+K2PgZhW
RBqnSf/Ze6LzHi6hpwxet8w+QJ6R3Lvnf4sJz2qQrR1zxlLLUvtSyK12aBBYhEWFJCL7Sicl+d2Z
4ZpMRKn4sdEequONrpJyVofN8mb39+4Nq3HMF/R/Yoh8WmbbZ3B4Dj67aCkxiMImwTgBQ0PTf1kN
kJqsRobSXV7cYQg33o7230I+URd4U+X20qO/nQpyyA0UQseZUAII7nnOhGuXcHkTC2rvuTydcs6Y
tN60glxgzBnmtngLGjYBGj7s5hJP5zqNR3YYuN+OV8YsPoHGAK0GEKr8gt+AtGghhfz0WdJdJ6NI
7x1vfFCMuROw9FWHPXHmDGgjXZIo2/+7euu8R8Ubt9hrI2yIEhl6uah9ViJaezusCJLsHTqrQgo6
l2AslR+QxkapYCAbqYEVSzIPrfTKb2nsh3Z+KMAnIjzLIfh4gjBT3Tx0ctEtthc83A+Sj+ZI2RVr
4HRGhCrkceohJLVWuF946nQvkQt9II/WWFWxjawqUNYRiyJQ9pY1vaTyCCfV5o5zzwIe0vaUJJ7F
7R76dhQCtMfQStWXn75qOq6BgAVZM31vcARc8XW7oIgtbx0/fkA4ftuPbVuUEwj70mMW5rHwjQo2
cRMlEVhSxYe9UCGA8VsTZg2ZcIquFphBF22Kja+pR4He3Lyz5+g1BxwxlKwGzts/1d1nuGLqOk/U
tG+mh1aX0q26aWuWnz+5pee3ZLCMn305GvjrhYwA7vNoOC7BCLzkbgtqnNQRGNMZlHampQ3oKN6T
ND7ItR/S7ltESjfNK5YgEm+FNtEOkiEqkDzsopUwb3fye6hd0DLHsJq7efc+hDLQbnGVJns5nPLj
txmlyZxij4Ixe87OGO9eFRscwYJa1nevLxjEqbE43Cr3rBLXJOxU/iK9namUosZPQe6PaaaaTXh1
PC43P5Px9ouk/tKog9VE6N12p8/xDq3ZrcIksGOG/Rjqti2eMNxnpYRtnHvBDO2xeNmi67gZk74X
Gn/ZqEoCmMJfuJitrlfCANaNhdMXb0ULU70tjPCImBVCWS0YKInoRGwF6FAT7MGgSjEO/fdq6qZl
t4GMONvG1KDdkNOjmIBEY3Gzfvsn7j/3Ix/WOG8n4/CoQPmrL1NV5xDKT3i5I31/EyN/x4TiPCik
qrOygxPr/doCXccNAhv0hT00oKlmvdgLuASoGPipEE21CwtXewjJ9FERKb7Eoa103m6PiHtV0cu2
wtRdOGYYZtLViyeyKTp7uyHP5C3gDbrxPz1icI1Dw7UEtBSls3srZh0A5AAOM95/nI6LWWMv9aIs
nWNEZcoi3SgEpRpDNIM8TO/dSxZZtD/MI+H3jg0HcwxPEibuOnu9hiWPt3Aqryp3njpxSy5j0zbM
NB/H46dsRrDyPx/SpLlxTsYj/Yy6uTqddw7W1Ug3SUph9QGEJ7LQBvnGvnjJs1spbRCCnZ3sgiSK
x045JvZtiG46cjhIu18R7PDEyNRT5BPA2DrLwEOYWu9bMjiQ773PubQDcfVTLcAYjzBOd3wO6N8B
57bw6RifYa687ZnfA5hWLzNLFqaO5LTyeiEFaFzwSNSvB/bq2A1FrODVS8ilhsh6jW9m9Rq+UD4u
ELpmkzu8tGrV/Np7ogUzQ8cyBm830nqrQXR/sQVoFQ9PtG+pm94xvFP/d7pQv3xTIl4oYX86mxDQ
7+BoLMzUtZVMCmTc0XLCDIgz4Ot9RjY/n6sSJQx4JVoDf6UE0094v1lar6RRx9MB53HwGLTGrXIV
sGC24/S/P8dPJ7uAW1oY99ZsAURVH8XuNoQBVUpuTSRBlnXRYm0VCrcjR+9iyDRhV10iJ8sGXVLI
9ppjRDB4Ce3mPEfa5sp+diAj7c1Qlz9BorU9wFfhXNtQBGWYPZFMixgphit03M1sb4umR01NZn5V
ZpwEO/i6l0dqPlW1wxgMs5gwRY4E2Ip67R0vzwIqufC1jKPXXyuoynZNZKpezr5E/seMwWw2G5G4
FsHPiVrWlK1sG+Md9KQiULIUZAKclXVEcP2ulBkAGOLLdyIgOElzATak4gdBelN1c7UZJj//J4cp
MqyyTg0pqJyFwzySr3fQT4mw6EJ2kOvRJbTbdI5drk2uNkXlkGokGwYM/uwWzxIuxBY58NReWFZ3
UCE59oJUWraNTT1vgTQAcnJCn60AtF1eyEUv+g+KdEbj8rhE1YSw+ZSgpwkbqpo9MQDgcQIEUFLy
gMMst9j9ssvHRXqzqEhxpOHjwQm2WpzJ4RSqqxI8XULlIPcTby0c4IUUaAjE9IqspKafySG03h5q
p2TwklIgnORa5ZG3rIBXsQn9zsQ46LQnPo7qoYzOBYs8vS2p2SgGR1hLmCR3BrFeBxuLpYzFzu1r
Kra5m2rDUmjS4quNr0DK5WMtyXkLBAEW0mFyKMFDluBg+Pn8ihsV58iAK9D9+m0bJe91z9Vy2V37
sqYlfDKsUcGYG+IThy91tLrbHBnAHYtXOWyMrxStb2X43y20cFHDhcGQaG0K7rtKVUtqyEuzq/q3
mE5VLUH0ize2lg078GovGgTZhq9uhVPKzlOhKY7rLNEYkiS+zb+q9O/w+MTiYXoghSBQfopZ1FJB
7GQuOSpd/GFpiN+96RN0QH/S0RQkXD5E9GW01uSMDXoYvi2pv5YtgHyYh7a2o2ZNTmMKTnwbACTp
7Xw3fWYGQSwfevqZE6IpwHiQELeyRAxZOfhiKICdXEafMXd/iBK7vHkiM2X320Sb3WOExniY1q89
wn6XHnaSHMavtjNhbNJP/xO0bZHldpexeCij66byGD17D8cGVkCrQZMey1i7HOqRNYaIxvVq5GNf
NtNqj4oX/6w/ukXXYlBItr5wmO/4+/k6piBnp5qO49SmzUNw4CMKHT01XGtCl2a2ic6S6ywzVchT
SSXv4j8n9f0wEn5X8P1q+q79uD/SlawyOMCqX38nyMyG7aRIEQYhuPMZ7iFz/KxJKn1l4xohqH/W
KRKGNLtw6neBVVlBviNKKcf4BmIZIAesO/a0bsXqmI7wJCHF3rsZLR0AU8UX1Rg9x7UYnfUmBOlA
3zFmDQPF8vEFNl86vsdIvnND0YOiXZLlBRdj1FS2NY/LYW/LyjbugW4cpDhOCyBiEAsqwPVp1L+s
yENNol2OeyNTWsNQuU93TvU6W5t+FsE4aDUqaPMa4DiO+otdwGSlxEj6jUVbsfpjRHhBnSMrWjlg
+McJDZ0rlkkyqb9UZ7B1xZWivogk0c+g5nV3q8zkGRSgp0Wv6eYpZjb5b3bVBGcRoMtheYpYkLfD
jsDpz3ZfyheRnQfk6e/D5phg2610+VyIqjrxo0sgYc/as1i9yVAKL7bKH0zgONevZsT5vrZ/6tnE
MZtoli6MaIhKC5xJ+fEhqRVUTuT8KhkmZGPNOvXFRmp+dmQ/kmRq8XXhNzNV4pqLBEapAJd4WD9o
i14uzMTAZFFKAhjHfBS7mHh7yUlqAM59vEpMwH0CPsCWzDfe4hcrYCm40531RN0Kvs5VDbIUvhEn
w54byMgQdiNG5jQXZEzQ3rHvu0AmE94e5DpMww2/SnUEwr8GaOjG/F6oovk5BoDUWa5jTnxxvfAk
iYHLqQ9kQDmLoNbNqB6oQDeIO/+8hHDVZggk5k/C/ddfKCSZbQP4qlvXPvEWV3S3qDb0Sm1fQdWB
UnlpAO9d7GRFH5F+crA1W1Ts2JPyR69omE4Ud9vULlY6nCRHoUNK2+NAYS9aRT0qYIzj5idPwBR+
GzQWzqARWQLcpbdPnB2PReMSl7EWtJSR/SkGJA1iZyDexvWLqzAsPcd/pK7rudBWp9LPDmgtQ27C
JjXw0L0vDo6aAdNuPRUoBvdLBRPvjCoJ2HP1tdekg34gIpRC9O23n+96A8tj+rKDy7gphObsvX1A
54V6C4knm/ohC40t6mHIsZScn4VziogSmXn5PlFYEMRZfYLXMQCj6Id8VmArDBQgxVmBe+fYvZLJ
Hb5sHch/qznDe47g1muYc9Ayuyg+tCxkJki6FvRrV7SSGW4ulYRhR4KctI1TCq4OVkVpivNddTMR
WfGWgCzsAXubp/4vtLQ3SAsrSv4UVYVNk16v5r7JWK48dArK3P2q/RmpIHIoqBYBbXAC9pqh4g1H
hr5tH3V2LaHAXS4VZmJRHff+PERrx1Y9yheLjw87o5EjpdeETsYnJW1IlAJQKgGOT7Ea1ZhrsDnq
bQxZTrv3Pomp8D2q3JbmSct4D6NnSmHErRl3eHdPbMuFu0Jiz6JW1XkKKDhvkizDGZtjb072V9qC
scamK1gAdbmMniEYFz1DJa4PjJFGdbtjrZ0nv37kG9FrE8tBMaKcGinQXjDOELznpwFhO6LXCOvx
jAAtHAYvjA8OHL4yopN/85i18GNrfOFIESmIfSrclh8wJ1937k65NEY4uYPD1WnAxUBCj97931MX
is/ZlRYwc6Vz25eBslL5wO2abjTvaHkDxLf0l/F86uzdg4wp7NXgsYkmj5tnQgZ6GXaFx9Z/sRON
RRj4NJ+0LJyqQ5vqXLtNPcLMl4uaEO54bWKH0O/RiZl7MQjFXDzXlHcJRYCFYGqhlLTN4RiMN7ti
mgGQZ9HzTIv9bTwdPz3+gSnLY/InrC+BuLO3cevNbrAIRWT2ZlzTBR3a1XOD2QfXJrMCCmuja9ye
q768wucGIEditerBa1k2AVKv73PAnSkhl5AXTbYn+gyDg+7K8DhuUoyGEkJCd+WLMu8nXmxOP6ph
w5yeg8XbhR2Rusl6cKw0GOvbdaZuZb+Tu8E48j+WVEiiIxXJJZgr7qXC5xNHEZCDWLeeWHu2owP2
W2SZAl/uv5Hf/707O3jkOhfXIzn+rnYseV6J4GgA5rU5Fh2Hr163uxzxQNp+NNfURLrgBYU1GzMr
dl+/pHhcEYA30U+hwRnj1QJAcm0Ur9ee2SJwKzLr75LZ/qeUPp+j30rqMBlgO+apxnpQCn3I9kti
dISyEnaPig/R7Aazszr8k/Qsv63Nw9VUljFO+kzXCfospFtgVbZns5UsGP/f7vHdR07n+wTwTtKN
llrQ2As9KUaOcFVj/zAWVxo3v9GOwKUQvhJx54A7vApfbZ+os6tUKNuP2fbtAUOy+gYiFttoJHtG
nmFDyr1rKmgs22n2fPkHNhHFohud75E20Nh1CH8QTjTKzsoruyJyk3j6gMgxMRV4U2us8jgU9Rha
4DIEk/wEykyED0ou4uOobOUrA8X0HaW7Fyy2TJnAkrWQIIEKpomZhqkStiI088mwB9DpxvIrRNJX
5ypImpP1Aed3vVjKdFoIjFNbaTVZrdplyDb/st8EcWlCOr/LjZkQtAYTyYrZp7Lmajw06S8VG72m
n4rUxNQW+sPbNHNnxfSAj2kFvPiQVb1JqLqtrBc1Cm58lTlZQg4ISP9iqfctP3wtb0b+N0zPtPJd
ccM5NiAdwbr58b4o2cMRhnIcU52WRf5Rxxw2oc/73rqsCVhOC9T9qgEQdKK+C2b9paHqnOZo4lFl
58srRVawtFlKfYWqSlmjQK8fyuN5xC/m1BhVE+NpfaH83OQ4WWqpKl8gs9+KmAD8U+LFvfzGQVxe
1eq16AyRXIyiIf1yQnjsN6Vdcm9lV+c/paoNr/ejhreyRVBI4MD+nuE0aKRv+oe7a53QlU1Kfp8D
o9E89JX7lWcq3sSIikmN0QrgrK5oI1ylSUHacgLcYRKJMxQL/DNDruu4ZexBVw1UGXF+w8xA0nkJ
PI1t0145Lszpz5TrCfnRFRMqMxo/q5QqPTv004NK/dZMWo/5fCu8/8X+zOG3HiMOky/yHYSP8xzJ
cjBr8TibUv04uwwY+lGKAFmECwZSQti7AgsZJeQR0UPzpd8Kbreyp3s9/XdXiMGCdWxPh5PdYSW6
p8wQaA2oJ4Fyyw7CAso0grb7DNyrXKaSR55oOw3lTbhJ6k/Y6NL0Q443n7wK4zwQvLmTrvphM8VI
ownMIJZrems+PWtv2O2TX0Ta5CMP7H0khmIWIdNYq2gg0OqXa9suzdZFwFu6sbZb6i4Lo9Empl2i
uCq/9H/37VVrPQw7dkHzIxnhSyVbLe73syspfbkHipH+H+OZd2sSoP7wW0aMOr3BZiMVHzLBuTNS
/3OS+aG1MSN9qcHHgNn1SJ44pVf40dSO1yn9sOXezYrD0BbrMyHfzf4geHDz5rCrfjKqZ6RtOqBZ
sFg5H+P1AOWyAV26DBw+ddMu6is11LSZ0YI1sBvFJM80tK0t2J4NEOxSGLypmgvbq/EKswYkMN4p
Px0G6dQmIX6ONcGVDtF/JqxJP5ZUAz3X5tV9PFquU0TteY58csJyUFNKE3qYe7n9e5m1St605l+7
qa9m8F9HYxUFgRAH4Y1YGYxBh6Z6waLGpjsWyE9AEI8imeS6MN+eN5WPypQqKXr9rNtARu+xZ53B
HTJ2pfPwvR67ZaHZtSLOGLg3bjZABzsYJM1b6Y3Oecwdm3exy0c3nHAJ33zfYV9tHgreUru42D5x
duwqV8QC+xgeDL7j7Glgt0wj5WqgCqkVCuKYVwJw41iwqGjHh3H3X1Rek39tTdWhCMjMGXrsu55R
PaBdkwYQVF9bW/7mvfqZyJVWQ9a3Up4JrlhImG6n5M+vMfXjiJzSY+XH3ps2zJnPWxcJh1Y0F39C
Z4z8bORMMHg0hlyf+DnL3VdylmHjBOswtTnWl6i3n+4jsanASXyUbdRIj89Iq6xb0RleLsZHBfPT
aa8Mu0AI+AW/WFg9ZKq7LrfhgcFOZgHl56SZLu2SHusCTpwvC1AOo0NJFe+D96llFSS3ccAiJKU6
+TLIzA74i9AQtgX1k+j4KhOFAf/AapisrQfuUme+dJdIFi0Jewy5Wipc/H+KBGTNrxkxG7Z+eMnY
HCPGGHdg5+cJTmNThmSIuKX7x/6VCjfAtvN8F6YvECnbYG1z0DlVRr8QI4jG0J7cK9JpXVuNza7s
vc76LypDO3jUQGQ3vXhB2/gNsnpOq8cmR27Ak6o6Oxdi3RIMbLKaNAs4CQmZ1pyc3rh8U2DVHd8d
AuTDBHNGVFmZCfZSPavwdDOj9mYwPCQi9mIporCY1a7fDR3b9HH51Cf7DFOUbM7PFoR6zWJFG9vg
0IcWwnefgvfeRnhg1VxSzv6Jh3ZHQCs7+Oa6cEYGJV2jhGqHOb17zmtaEyN7lSCUVeajVo8daY3H
E24jRAiLIXhS7heriez9EMJ81iU5za4GV1yo47nV0b6Il8OTzAjaZnrWGxA7fgA78wSF73r1OYYo
X1xeKGZKipQ1TWuwbt945JH5U4rYQ89QpqaP16knXJgi7gCu17L9tTosUAkaKwxt4pfcO30Kb1el
QBC3XF79U0on0xCbibf4ZE0g0U2ObW5EJqA9sUZbTYyA9nScZqf8qD5S+6D4VAojhiDBqEBrb1aU
By5OiK/2uIAhw9kUbSeBCAvUcOA3qacQ4O9VN0etTe64khhmYzQ9t3C5WalvwI86tufTfmDCc5WC
vYM9xwhHCg9F+G8USkOt6NxAdpy6wisFK6xC3LPekG4tmfHUA3UvsKE+DYY60iNLWgTn4PTDupSr
WpP/SewJID7s+JQGnd42HViT/FwnmjCfHdyAEmaOOzX7HfowXcYhCvi7zOsO631rDpFPQdf+Xr9V
wBDihg+jocBFrkWTfdesnow+vroSMX8FK6Ba5YCwsl6OL5R14E8oO/AOoeE1eF2JVzvTvlBXfl0W
WqDCO5IysCYmqBNi43/WAnWUfJ4jAKDlTVuSpCvntMdPkUKft7fItMBoNlvYBQ9maUpOUImqjWbt
78DryUXMthEZ2vXHlr6L+0/0GxQdnUHE9vwJF9uvukVv/1ik9+VFvqX74eXP6kYzvFEQXE5wugon
nSJts2lErAfGObbTSKAzqYi+MHNOEf5JF1K51W9DZOhJvxmDiJZT88TjKZG05cvwaqrxFVO98gGn
IEYNOoXYW6jpS9y7R+/elPBJLA1Zme6BjqdlZQ5S+jpXZQXfrOiAJBm07k49TkJGeB7n02d3pzeC
psU9y+2kFj1Kq/BWwKsZ95IEv6DX5o/kR0CbVpqbLnPdqMRGgQsSVVr6etG5w8CAO4jt06j2O019
S2aIfopd3k+nZOSQei4EgmKHHrc95ILZ2ngt2OMc5bldCRJdrx2pc/HxgnSquPSa4BBPGzqGBsAs
ro6DcEWW4M9Q2m3WvUT2l1S5/aO9IaqpaXMXZQapXtZY3A6Zb2ay8aJ4gKWk8kdgcfS0ZShZhna+
hxTtualTCDMXJv/h9qXrqVsNKH6Ey35OsfVXM3N7vHOblqSR82jVr++5XPFOTEl+4ORK6lw6gXGy
dUdBVhpotjYSVKsuqY6YnjoawAe6E7gaCAipGPYxtNtgvKQB44qUjGNMMvM8anWF5AI7MY+8n+cE
Vk7JD3/Mr4RJLbRUvFK0zCKuhUkXtmRpKirRwgtdNVhrpQ1AiswAFYrgL13/JRWdZKsf/qZY6xKz
YB9v3KHCVouuBVeqn+vnAvv5lzWtD/HCw7OYTNrd2OUkQYbRNXAgtN6YmqgW/XtiWkKmPi9Jq39u
dpD+VpOXrcu0eBpu6cmnwPLSEBhahINV6ntoXKdneYfeZv2Hb1SPGIS2P3f7mKxAIzeuZ0/lbI+j
WKEQNbjQQju03yGJppQ+b+8M9COZ7lHoygyIB2Bl2Q04HgopluRMGyw849EHYzYpGfVDmIcPbzol
2dlQVwXoXHWdpny6Fm2GTJMj1O2yuNzRQHNroPDC85D5QiXcQVHeuFeprj5DImQIaoPFLWwC4Nyf
UqZsvJfsregXJjN9GOcZhAbERhuwTnphWLEF36vJyVoQa9FaaX17MdESL50dktVgujvW14ArQ7E5
P5HdRerOgCAudUtcz2vEY/j5rm11wJIdY4yWqAf1lYoaH3rxHe8ezdUwxQ1x+gpVDBDqIjn8E8jw
o+ek0YgCEnj5sqqH7gD+EDLDkc2A4W638gKhoPjN3qMcKg8uctC3sF+ukJ8HQx7xOyG76VrPUPIK
U/Ld5iP1g9ObVsPlRT5FCaW4i5ol91tCGOTCXVzO2/3tMK/0As75dHBK1Kcdq8276p9dpqzz+EUX
U0zInShGq1tyEp2fK0vhWhRZYRZf5B/TVR+a+aiMbXAS6P+d6HYFNPhZWxuy31Ck8YdTchVkCuAc
pk/LLDpu248+VO5ddKG/ptX55evcbYR0v5+3ULhy4lQURw5k+gsrag+T+OwRvH6LEdj77UtlsqAN
FiTDJWbgVLQW1OagTwVskTODKCUhbn/PhXlJuib3uHKI8/ogAG/pVo5slRj+ynjLkvNYhCLNAdt5
gx+B+EpTK3fg0fgufbmMlkQmo2FsLqcyEeKoONExYZK067cVibeDhQQgw8k1BsgORNDDPtH7rrMQ
B1H7omn4tLFVDPiTXLdcC80tSuGXEqCq18bzbepSTNC3Mo8b4fFXqkN3KWHJzH84/IetJCEb66DJ
Nd3yfMQvaMqporp8imTRsksAUlwa3HfAJdobD35q2T+MtbF8Eo8Z/ftkU40e4AjEZUTgImZJhVSt
XfkxymhkNqRZnqGq/CKg4oyw4QNKHh+09VM6F8fymKnub5G3RaOyHUch2/3DrxT1Uy70ZnuejZNK
T5uq4WXkhY8/ABHTeZHJcwI2afvJzg168RvSHLZb8wAm6weBMx1hwKpNl7P3okQ+k2YHmtmWuDov
ytIRxt7mkBDjo3JXKZlZKi2NnUABx98GyXxKCKl91Fl/S3vytzo0dU0y9RX1OAi/jeMyoUYZ/HO7
c6PMVXpFIIbOx9CAFcRkNsz4gm/+B7lSPCG0EuzNHv3EUH2764vKQbDJ/8sWNKthtODeqVpYSKJH
Cx+WDyH6jAIVmZ6ykjfOUqFR2/PdqcFObj2A3BgvCsTAP2zQ7pGghBClftWZKQOhlksc8tsvitJJ
60G4G8WNoy7LmO80zs9QxkYANieWaMiFj17wtqb66eeU9y1wS27nFUcgVSlKljhdKRjoIbSFtZo1
r48/kzmDWICb1Jq53/1ae5xFErTAMBQxPspdJDuAJii7EKGMni0WgHLW9KNYy6MdGQeGpBy7E2Qz
72IIahTQ2v6i3CeISLDSXbE0/6TT8pV4q6RcLQM/2wlKdf7SWfDFybjKrn49VlWeFEjzFm9x/1sJ
k9CcXVVAYoS+XN9FkiT7bHAhBkkDy7xekgEYi53hcLJoRDcGfuh7wnI4nrZ4AVlKNKNrpRpCkL+D
OKXGnYoYF1/zVpIMIAtadfGppmvjcBbBVzEE0Hqa04+1WfKuZwSF9qOxcLLLTk85L/g6e3sPieNT
Ty4pZngW6jnWPuMWSKwOLHL6HqJp6fLlFEq++qs6dlLFB3W2EPdt3OysT/04/ZpwrqIWPrDOVGDC
zoJDj8kH9mgFDthngrmk809nwIpjJ8QZHTLWGbtUH+TPfnz5TRNIcPa18cJPKfFym4A4ExQ53D+v
eIAR+xdzvufpmO9JwySlxi+hBayuC1R7c1+OQ0GCV/L/xBcvL/J9rHDZ2oH61mq4GnV0MxaBipLJ
8pdszTTfZFYVwcJKZXeRlxXmO8nSQDrTiBzUJD+z9Fc0uBilFlXmOWxXKQTywTS6AaE9HCqaUcFA
S8lid90hWGBd4gFjyKvMk9NbZ6KZ/PXm/1xiOBHba6MVAVcp3POY7JS9/DODhk7qC8oqaCY9xbVd
9SB/XyuVxlMdJ0xmlosLQLgmyJNYjlLQIZ50hbc8+TQ5vNINiPCW5WBXGnhUo5D8g07EYEDOHDQi
xnYboWh8gyQuGBVk15nNTjKuejIcrJFNb0tjU2YvliEEjFCc4rkVeS3dyKNOqIu88YXSo7x89XQ8
6Ymua3jdUmUJCSVErM/UdNueYB+BWL+asxtDHmS5AciuJMwacvLGKtFam94oedS94VNYJBQ7K+5j
GoIkoOkGMqt09NaFCBlNqRcqWC6oHAgqPn3EVXlcQHmTes86E41BiILv7X9BQ1yJXzuBOY5DnEkh
m8lIvB+OVVwV0t2fbh7qXZ5u6gtjTT5rpTO16EohVXXcyAURnVJpedH3ihyjwIkWiwMpc7134JOm
rjaGYM6aQNGzTQ4dj+3GKvASU19B05JSTcFIJT69ak9zC0aBCT3lFn2o/HGhQHT7J0cVfJy4nt0h
5FMZmDdEckF4fTK09Uy2+hMqETvAYGrUyM+bkAHryahbpWf5dhELQxlM/Hf/KyW/SQXRa4k24cIe
FWqQaxJ1R1NVYL+PLVWkGieV15um+kn8ygaItstMJHVEJbneWmhmHG4rZbRaiY9rFC5DvpnQjGe2
9/Q4wZtHecfOSjCDlQgjfnHPb0rwFuwCD1l664/p1FdsPw6i2EICaH/Lw7xLW0nZCuVEFT3lhZyZ
MAn5uFrN9+Rv5n5FOlZ4PgqCXp45NB+bY0K7xcR3PIPtpTHejYYlF6V0tPw5faI60TjfkuN1DPe5
LQ61VsV2UUSEsWSUEETllLsriCFJUEbHmnvV5JG3Ciun5qNprsMZt0Vjrch5OmqXM82/f8hHvELT
RP7gCSdgq0J61olZYF+U2mHZ192pw/5porlyKQOjmZZCdk+IQt1Hv7b0EjkK1gzAc8lEorHK+duA
1VUfEaB5mu6CrYbCn0hWncc+2diy+bP9n9Ldvlh18KKZOaXCo+JdKf8AJXivtFmdqgj/TFHM+nAs
7RS0ji/eBqtwCNrVkSOiG5c40eBngHmDjJa+T05ebvQABzOwZeXQwLt5iIJMPNlEW/aW0LFrx1fK
LBUXb02kHvwfG8Nf6lcDdhdxjQIij5p8xH1F2omjv4Gmv9e4vnATKsJiRMc0JRp7bM1xw2YbvZS9
WUCKVZsF3Mmgg97L+VCYYghF/ExCDPpVdea7Xqsljg/IEEFTPSmH8AgDYV/9SrYYFN2Z0WqimmSn
7tMUdXX4uhRjzLt76UNPEvI1vjkJ3MSVwj7mawg5UzOZ0bfOZKKR8qi/0KMUqXvVaWxaju0/GfU6
dt7kZuQWW8zdpP49RvNawU6QbElnVNRtf1htVgL1zHH4aYAIXb+zHtrE2r9ohpvR68F+c1VQZt/R
XeKgHxB1wuAMYCdTJv2MJ0hhBC70MmSrqWiFu+tp5udLbk4tmxsBHxc+1xIOBKDgxWjG+bBxfXU6
lEOW+jMtreJj+q03QY92KXmYag3dnN0O+8LsCKrEAAqVpmLAJ9JUn0zJANbFX+mu9n8zArOaqApa
C34PFjQZXworm8xwsz/o7kJ3KB8otDO8KAjUTEIKm0G7lZwHmyCDdcrWU1xkI8XBfjGNoGugptJm
DqprNXp4w6VxXkgLsM1bkXwUAgiFI5l8NHsH4YAchvLPAOLWEgQSA54Va8Zc6EhPNwIXEcDkHYNS
+DILvP2F73WsCi5MPrD+oXkK9tyx1dDlEWBSzw5waz4B8ut5hgzsTcEwIsY8ZLn4rwyKHHYueT1k
aJw5mPfGRQ6BBOwlgdScp5qqsUT+EEF2hn9D6lWegRt26VEM197LBwaysTtolO2Y2ls8ZKp77VwW
qhjuZUCqN0Z+FKqKt4RE1GDCLOECA/PV8ICWRYcw2DaV7rukG37lF/hAwVzcDIjGV1tjwAZYI3TM
+DslH7SFQGRdV+S0Y1dYWK7X6g1dSD6Gnahp2B4cZrSinXFh7+BkGpFekEJIf/JUsAibyomp9oPr
rWwUCBn/CTd4LbOOZ0jNuwpiVEg2+RkjgBo2/vkXi1GmZ6p4Kusu+PEdLVAWWKhBVI5y8SKJEajF
51p1WuClnlrLQxRIw04sPR3GYf11LyYdHFzUM6mSGl1/BQXYUO7u3TKSgMAWFjalYxQGmYe7wPVY
5vzoZyqLjMEj810TK+JzWHm+M3cBEE14BDG7PnhSBGI+rwN71HVAwEcgCIqJEPV0vSOapAEnUC5L
i1I2sniN9dXS8UybZp37NDpoPSsfuPb3j/mblf9+JN8HdP8vkbqM1ACxmXDzTK4p8sRBOgEQ/vBE
kBw4og0+C6GVAQfIzOKTCgBpK2ncpf2lB/Lb68eEZz4YcbvgM96XyjwX/LEMIh5+kZffba3xDg3/
JyeTmAjclrVKQmthIJNdJqxZPsa6k+T82GsfvPXsUh7zG8enFwG8TS8zrGlt4jMi864RsOGHYwy4
1tF7Zwta8wwVCts2UHEjIbMQ9AvA/qlg049tTTnSkuvAizpZjY0Y5NK9Vy6UE89WnAam434AzWgJ
zjsgcSCDuZAeEwmcPFdQDc4sw9herpSF+p4rliHmRhYvztktypKO9/L3qQG7UcxHpbDQ+cFpnYQD
ZqMWVo+lMj7Xq4R5W2s+sdzSTBVxfdGePHGuXUkM3inlSlWmcg6JFtIZGKxAfOCRu8h1mwNGfZyk
HyidJB2IKLDzCbt5UL2CGX8nH276gSXYC2VIhRHs2kXCcMKwA8RBsdOUZcFgzeBrQk/FvdESG1qU
xh0bDxviiFIF5iLk8FDQOOCgcXcx0Yc3j8jR7elxfzvXkRDFen/1J+llVtExvRs3BsduqMSBfyhg
/t+KXqT6KhWhL5mF23uELtodfKisLZ6VRO9cJnOsyqbtETd8D2qN3ajiTj9l1GgWs2aCJhFFyEsM
bdisaahD+irCaLT/3lJEQNFAABvvLMZImBe1+aLQ+eIttjdmw5HHBOFYXfwnVowPJgza8vgwy96b
n7sCirxCQmnCOdsGE3rz8XzyUL1IVdPHTwpIosbVyqLJL7wnESyt5rFg04nqWn0EFswdDoWIn+IO
QEY+3zwTwpWt1UpBhyIMF/XlgtH5SwTuq4Aw2NxTistNyEJ/Nv9E9o1GqAdbaDHfQ3fVYhL2L86S
5XCNRK3yaXp2OOg9jIFVZusTUDjDXKv4at0QuEMoP8Ghsm6hJwPsfCvV82tkHYfzJXPrb4ZAxkWO
eGSuvJPLlm5FBA81lacZ4xzYgslSq19PICt56/UQPzzrtvZa+zU4ppMnlRK65/Z23KliQGL3CHsz
4llD1i1OJlBhx+ZRc9sBCHl926VSdqqE159JTL4DnD+ajxRxzeNT4GxsArTk7bmfEKVAMJ87ecGy
LzGZfxqZ5p1cbjJ6QhcMLIcXouHAq9rc/O1YPHdiOy4wEWictCmBzNo7SaRCMsf7LkyNwLyvPYu0
SuYv+w9nd7kh+Hq1DvPJGIlIm0EgWt3EZO83yulhnXXtcb4XWcXBD7F1v2Xy+IiWd/cALkkiNkdU
5w0+pnadw0ImGwND4F6dZQlUbjJ4kMh3/29EvhoHZaxOnkIOS+5GDer8QYuTNh8OoIYqlHTjsn2h
bbYYOlY9s4+08MZJeIcylv6fsBAJKWScwv/X/9s8hUZurBHULAUmjvuTBTMsFAs0hbthqr9UksIk
Iv9YoA+yKy7L3B/9ymAZrbPhRLPXNQzVqKVGkJ8RvmeJoF4QmN4HLL4yWxDj3Hb9QpBAlkG+355a
GwZ7iXJgnRhPUivo9kHy38hmIOcOozzkBgtiuT6PogVnyDHJ7GOYBxsJpjivYkMXIpvvmASQIlM5
fz1a/wfDQOIjxHlzC2YupNFyXrxWnD7z2ecsWKGqEym+erNKS8tBumt/wd9oKbpuApDJXnOGvIeX
S5cLcZsoIFIeou56uMnvqUCJeIAyacm0FmFs4LfoMcW+wfi4LVrz+8FePg/4a4sLxabQmHxLhhfX
8385tBebzlA6OL/gBfY3tHjga9dld0dg6icNfsfQbZC9nZ9fZu9vwaz2SRirFt2w4fCIke2RYn+X
q07R0amT5P4mey5N5mM+Zzp37LdfC89vxSUYhcShSYuvmqPawG1vq+0xFJ07UY+RKS2Go/r0XLpJ
F7fJ7sAJTVEshMWv26TlygK+sZ8nwTGO5IrHcjLvJ+Rd80+sSggnhiYjD7/636lVwNLA7TixKAgK
Lojg8v6sO3Czkm17uii6xXpwtqZyVfacX3jzfNtaaffP+Jq2g7DFkA7R9eXrfknJMJYFA+XJwvme
gjTwnB7CZTH1mMdB39O+Ipt5j+8oUK4+dq6n5WjbMVRwocFlJdKMnSQ3N1Wir6W6J7enoQ7RY6Ng
eua/Chb0SLeB8gtqjSaCohu0AqP+JhOfBN+BvsWHtcWXN9C3cYx9L/RpQI/E67OxK7XOaukmZzTy
A3G5lNhv5NPE9CElLwdf47uJhrS4COkit7t8wSJZCF85OFncmVmClztTOjcn0d/9j14qpyGNWBXx
XiV7sfrjSc2J2wKn1v0jCW798KFfektvebV754DZDvZayUFmjGGGZyjpUuLszwpP7v6ij7hhDfbX
sn5tGVQOAmY8yvIdFu+LQgof/G4oApUDf0hrEWJkub+62eZ7jLtrNau4JGmXgColqcqm9/fhHU0H
8CI42b9eye5/UQBD230arJACXt/C6NoOWnS2ZsxLj22WCkdXYD0W8hekQoCiket+h/rWbMTZJ5ie
c4IFzcdOospSFckhWor34HntnXavNT4uKcBCfUt+S7j9VV7cvVSnq6Rlz0NHX6vdqQcwiOf7kqfU
2RBxh72aUIEvztyfw3In44lyItQzFv9a4CqQUIDrQpiCkAJAqcdPGxgqgYgiKArVVJYkXpu/MJID
yuH6CQoh01ckmx1Ok94o2WDkaAlLfmrJV1il56dizvOuR3T8zpNsxSAc9/K2QPNq6/J/UOEUg675
jqJq00v/xdiNfJ/btpBualHn1/tnHlqEu/Uaf/vSw3iA/nPxBjWyaYzjwqvtrSg7GIO1yzFzD5QS
ku85wpIfGuSRRISau4bY0jSBm1IoEixTAVEuc/S3PdGlu4+h3oh4Az9dBny8XUF+nf9A9fwX39I1
+Z/nkD4jzyL4keAG+7q+Zr3vSEaHA6uyZtFmQTjdTgcaiplCpGednf5w1Gu/Fh3bFL5tVvAFBvBC
L9/UygMvGem+F3K8XVghBPEeSCvF2Uekw9QbRmqupxKlzEoM9JSTQgIISdPvqSrfHKWMqtPOy1ka
7+BA28iY2geEh8m8QTaObQtlgNVXpl+FAK8gCFmd8p5KXg6Kub4Pr6UpOgr5B2MFaBAumuQ1VHN1
qQTZhn4WC67qIbnIJ+juP2RSuESFSPsi3JZyf1FreR+sRNWdXzIyp+Hg2AblCdZH9sqryNUv0uuK
YkLsdu8e//bgl1xB79o8pF59NYZ8Zv/joCP9GeuOYsDvRFTKVVYxLpN4h7C1IdL3akv5X5PuKohf
pSwxZvZ2YFpeIRnyAyEvKD7Qp+gv46j/IcAwAReIpdvImBP+Rj9h0CDhGRMZTgwNvVShP6OfMb5T
Va7uwMe0xu+O9jgRMnZPbSg2qiYjLicsG0VNd/75ywKihO8TaP2fVfcOOIQ9d5/i3vCV+9qu3hAw
QBYeWmC0SmI0eVQDFDF/BEwBwRtIQYakgP5S/RIdBsM2Ks4uFeIenYaCLEVIllQ47C1vUlgDGxNY
N7Vg4Eciax7QVwalNRgzsz++kNIh9bkd7jVf0hhFrxBs4sIMpNFg58wwh2cdD2sC+N9Q1WNqBqst
OXyD2g1D5VE7kVtHDv60Qc5cQ7iZPXnZSleEKNpHQo9nRfHPh89OMGqRZEra4L4jbnt6fJQE6iy3
QUWgL/whYZhuHEeHXAQJBmviOlp8DT/x0/tTXkcSVIFceNG7S7ySVhtDf8in+EI/KkN4hhFaA6V8
ThbwDnrJyRsg2Fpu+H704maLLXkMAH4iamAuaM07vGGp8R0+2AHtjGYDqcjOPOrG57OYbakNbmQq
ZTY8lvpZgU1znVKoXMjuxX2XSxzkkDrCOTV866/a0WILMsEbExDHRk8Ku/++weKxq56ORoyj+V2S
q+8ydmwg+gNNRUAnfawu2/5HEGjeCI7cKUZtIoy+rnI9vgOFfpdNR3/jq1PTiZF2RrXPfP4MNXQ0
PEAfrsn1K1pxRm8MDwmmIwlk/77h8jSJkxI1lVLeHaj53vJbGxHLO4nc0CpJbTDNYlPMPSSHqX0Y
qED7lxAt/p4kOw4ZBGrxIsOGcltbi0+vaFkXp5PS356mhGGXBgYdvp6gtwvVT/h7KWIDqFXdFqZ8
nl9WZ9OcBTNMSl8jQIqe+1nhMXYw7lVN2mTFbEBPRuRlOR8gXC7aTOAeOJDygfCoJvhXuYS5gdkj
dQfwSXcAx124VKlJpaPWjE/T/rcMeLScVnrB32CA2MsesR9N3WMP3E38gKJFy5axZbb1wlQLJLvx
4UH7BT5esA4UcT/lfZOtQ0MYzQP+/h96unvENhfaN67l9NOzYBMATlDrnYSWyuFyxpULVroldGPe
S2Lxq22rB78drgjezL+uOeWEUF9gWtSrooK2Xed2WqTw1bomRZ+uDzjnkOkUBCH+LszTMRHNpGGP
dX1rdQO7oGAoFypRESYYv8FfN5jWX/8Uv7nB/mq0XF7FZedk8CYgz2AUFB1pJgH4CuB8Ce/zHwSz
ib4yNa2IMj4rGpJlUAhdBSAP3uZCUAxrHuqJFmmWjMJYGlHY6yrTDAKBgK2Wo+UCmQXvDBoKj1lZ
DR5WpE/fj9ezK4D7bS92hrcrfnkf9sydsJPiKs29cUyEKKbWKTyKHNdgtawBHMS5iXO1mcvVqaLZ
Kv3XBEOP0AAbfMdx2xG/9kEpwr2c50YGCNmGaet6jtsN76ns97ajWzqZCZ4HGeuUwpbPX/iKNE1Z
I9tj9xUCJb3l5rDMxLSBfNH30+igkgbS4RZ6G7NGEJ1JISNJTB1wpC51beu5rULOqga/1U7Yi2QY
IJlp5YzGOV3cKTl1Ecdrxjh+MpjCI9AlzLaZgmhZfFJbRSHWye+AsJlkSEJOVpYkVghlBwunpnI7
YFkkdBLngE4pjut4EUMzvnCWzCFMv+KrHlzoZDHYg7mjpYOGlzXf9VkazL+J1u3WpS57RLmvMotl
yvBHnK5e3gJK1UASa/+0sB4zb+8sSSv1vTxWptSpaQjHQpn48m+EH+4lbDFWddpKLErhIYics99a
L9qq94bz2LpQqtjvuRykQkgnTbZFF9vooB3BIog8pyX9lrTWLw7zNVha0nAZXtqxDt/lWoInpfo8
u4p5adNIU99eGbdRng8sLYzZ8wyYqBd3rW0xnkDvU6u9qUqeKFYm7jAFcS/93OFF5ceJy0WI072c
c5tWCQt2PS7UL+eT3DljMYMT4lZpNlNe08z4PAIN8VVExwy1eNQfi53XrzUvnPhPPl8l27j1ou1b
sviE0qtGkFwicfGS+OSTgjoBCjdYOeH+0DknXBi61aMCrzpucfBc7QCDkslr/OZZr/Gb54sfTDrA
Y1bHPDiExXY7EgX4qjZEQ0+LhkEwnSX3aYC4DFrwpm5MR352QLBz5Vp8C32ExnEio+/WWQyICd9J
rPBIDWwPXm0J7WHcvVROO059inlq8xZngD3kRxvCOtiBHaMmJgYCSq3rrSI29Y4OuWL5mTcNjTDL
Fx42CJZA1/r7Bxt9hFol4yxFiYj7orz/hPRJtF/es/mYXQ3Nrkl7Uc3lTLEekZOKnVHVd2JVTArn
gPBepwC/PiQEuIAZ63vidgORP/45s/1ehFYapfceNxOiaHBXDoCYkKR6FS2tJRzT6YxH6HNlGcuU
zntaEffD64q9mZl1qd0r5+8U7kwgc/VgibHPYkScqj8IIdTQHZshsOu3AhRWvMsfhueFOek9ChUp
vM+oMsT5MD1FTNRg0Ye5w9LoWgXttShBG2GZ1pVE3OWU4rBz7vvcsSIRPkWKajd0JnTSlxN6OXzQ
BhwWew2qZpb+t6CNEY1oBJKKv5vLw/7FLXw5jMtk+fZla7fLiHEoT14/sBc7BKvXYAEj4w/6t1uJ
nb1H3xni0rPAL33BGXG+/cVkCKAL+Xr2ZDT1piqVKIZJOmUgL/lc2DyKyX98UGukthlkcq5Yge2k
NE6Xuayk0I8rSRoJOKebsgp/cVk4K4CmhEn9uX9kpVYfljvu5iDck3QX9Jo8nUFhqW40JEF9TgKU
yxvXO1Yl8kRcaeERVlg8LTyzCg3rz7M+b68OWDkyhPe6gm47yPEOJpgAY8r5gEq3WlqicfmqMJV7
QL8g2RoT+DCzb6lYOBTJMEWX/3+g9Xw18J56S6TgmzGG4JoG+dK1VzQlkyGlmSVRXU9CYATbBq2d
7t8jlWnLIpSMSuXF5JGnBLY+KYrXr056PzbJQjAkS3/pVl4FAJyPChT5MwpClhR+kMxoHX168GA9
/AU4bWyyik4rdBBp0LPl8RJZxToDScCEugPM/TcGN1M2v+ST5YHmWIGX85yZvvK+af+jSeppr3lk
lhW/grh7wHm1BpV8X5diItasPS+dr2C/moPf7MqdvgyRFpmoyIFKJR86OE3olnQQPXUlQ0nS7rbC
lEk6wszL8aLBpMLPtyO8MsC3Ckpxk3gooIGK+KPleaIdmQ3d3Pf2NHQ0awV7cxyNw9znigy65XdA
jF0G4YZi2tM9+TZvf4n/A1wq49p/65qlLpgJHOiwg5UUvFqL85Hcn7uKVWxxQerzzbmurNHtnM+N
LXEcB/4CNJ3pdHkwOTf11CazrkJdaIkAybm77MBjZrJQLtQ2z67+Td5h263+WcxdYiZJMttgd9Mm
9UcZVRWai1xqyMo6u90RPnclSnkz/rrqQm57vKD5/3R79GWAv8J+AoJcMlTca4nTItDDuW+PAaZB
X4B1EzHufDy2csBqHDPR2QSdKO3Sxi/xnG0R/kxjwtKElMrvWVLdgEAODrC6X8gEnAmEww1y0jZW
7XwNdFXxp4WWzng5UB4vJXpynNM+hMibNBqNdOmngDW12u4dPgvGwCDax1qC+ZXQko+QXbdVowqm
GaPyNxPLdWxeWaIapf0B2Zii3FWMUUfug5XcezhvknJYPbX7bt/iR91m39p3KoyjOHwuowXOxFc8
xNN1GP67YUlPbEXcDCV/l8L3w74nILLwYRlQbu+inyVwPexZNRIS40bhGY6fU27NBfQU0GJPHa0t
dTIdFduLHgA3RrAwnn6rFgSl/qY4gRwm+04ZSs0RjnXqy9Py7mhks2oHGEV/H22a9i9iY4JLbVkS
jJkjXD0zjsnwU2HAqHNcZuGJWEXpNXwqGZFLIOg1wL6XnzqXeCGfeWN2ls/9eht65AS4rI4y5l8d
pDuW6tCsJEPVRHSt7sJHz3CWUn3a/8eKmggVYOhX6ZYUkjNQfuVJW69JlO7sA9BAJtfgHs+cFD9P
m6284UPRmZGkm2jWT/4K0b59JOD8OEi8x4U5CjShavGds46JGhwo4F+uSsoTgIpibafve1/LA7Gq
LmHSTADYVtRI67yQXaTBLt1kh4EP2rMx15NBumTbkTaKRlhFYFMZ8PShPBh5Cr2Yfu2NtGvI9zKZ
w2fJeuS3+746ZN6pj09GogdjoA5BlHQCFGioqI1K0hhGFIfn/kQiMcr+2e7+kMDp5aOM9qMp/hDb
Jl7aUGerpwLgqVXXPzX9Iza8Vx/BKs7nYrMCKHnp5npHRX7TpNjNgHkaipR8/ut5Yg2aZiTHSNNl
/S51BQ8fGrTGdedRuhCXCWUhGNxCesQDHiz6BFgF3NakeHNA4nJErRUdhUNR31fPNjWEh2XlE4bJ
PEex3rAc7nTIDvqzVJkU+7MG7zq+6+O/Dcj3UrgAEHhHAmNYT7hgnjaJknn/Fuh5R00JG9A0oKdU
pBUtPYF9SOteYaw9Idy1v5fFGVcRx2c0ZAVmB/HMbmC3bDFc9BM3DER7h1DG2xH9kvvG4ULPrJnz
4KBjiakCgJEs4+xoB/RN2fmgNE/8EoOOUXjo2IACR/iMs3bjOwGqFCd9ihl7Qf6QsdFXbg6xOI0g
+zNTpRDjaRhq8aA7/iOAonXx0/F3dDGlAS5G99ALfGqTyI5340V1ZKVYSOCs0Fp8Isj3sDfjZ8Ux
nhfjGx7GDMXfbrsFEuQAj2BWFjAMJD9lTBUPwvCkN33dM9lP67pY8WHVHwXAhKfKLl0B6J9QT3ai
Zcf+NUaUhTwR8cLdUHEAYZt9PYXfdtBjzGXwle4JH7dldLD7SYL2YAyLcpgPJQ7by0clyxYpQ7um
xZ9hiNjd2P+/aDdI0B/UGMUGJlY2ObyS+AfEy8Qp31wlpmIFTQWh7vQZEqg2Bd5ssYqRaGFpkVp4
0p0AIQ2zvtDgq9U0Vol9HAsB8y1GxndWpOoaX1U2g91L+bpS0I6NTMS7x5HIcMtfgkVzoG5ndt4b
c5DZQz3NCA6lehFBylnvPZL3VgIUqcsXXVCFIacROiMjCfzB11qPg+LRFaIWZps60saYJhlFuSOv
hQp9PmsKagoKRquJckGpckbMVCY3llKSUbkv6v3DsCLrrAesG1RVM6vl/L7sOQsqUoUmgBFNpgIx
Dqm2gwwjFghAqzZnSjznS6l/Hd6ICjcHxyV2Q7okqVW5CLnd9UJX8pYb50eYdjeTxQrmIHZShfgg
AlQWdBUIODu6bLSYmjbOO1Km6BAGvIADp3LEh9fj93uwvyNtx+cFncK1YG3OOQWTWnk+NC1LBlfF
yhTP3A6osR5Q+ETSkXHThB6I+7z821q2DIzt39mTYpPHt4zZF0052oU1k2MYMrcB1eAsvmD48wq5
yaeTgfS0UzfoZ/5uh7IyKeEJxDjpC4PVzaYAPHOf76t14s515oB8vgws9iCCpcbTT811TB42RNq7
Y7hLS7TR2DcWP5PT1AZPsmUNNd5JMNl42ouBW+Ecwmu3FX+kQbJ/zTyXXu25fTmKtstzVk2mkiRq
ps70Z7v2OyJCOkZjAsxzmAzuzRUXXU0fLq6lUY1uii4FfbBXzyHGkogMDS5L8fl2buEIfUAdbYAW
u1SvD4ctzs06oG7YgzQJnVVCUwm2csc73J9xoz9w1SVn6XGjPhcl4QvQjNTttOmvKVIqwp5g6xdj
sU3tkNOds2zGB8RfmRDsVirJAwwJ3jZRcZV1LwJLal5x7bsiCfS/fYN2SA7lrIrO3jcLBeTT0f8Y
z3pT3tHHpSQ8yqTXDh4bRjvRtgeGDwCy7AXXJzbi52B6NkM66Dey0ZwzupmbVRiVwhUDMgC6ENED
r5rvza/TBOcQdL8vy9tDIUIe0zVFSvFWbvgqt1iKLxdqJORd1Z1MK6Lo/xN+ACpuPvdv+FRfDIdq
CltKU3Wi0PKRhSrZwjJ/wvNJzl+gEmNb3MY5fAodCA4mluHCDiQTYagm+UyrREcGSxrmf/u8MXaR
RCn842GDdDnkMwFHHesGC71kTJCAgOJ3jK3Ibz5hm8JtZRmOfZX6xhr45gxx8TgW9bqEdO8lyRUx
IM2ci2++jzezVYzHnc8hQwSFckkuFJm4R/J5bmS9jCyNbuAp5VgDl5WAx//BNAHA/6kSjZhj2K1O
axRCqPQbmz/gTkHwgWuEiWzVBgHDOJK8jZ7rlKLJxX84eK4r6GAVzEKgQ1GVqW5woVpVw3HQEoAk
Utz3eMCYFaA8b68gC2nb/72nl1I6pmR2Y7fvF0Nupwao66zm5cO3ATOGng8CSY8QbN67S0QbMb8t
b3Vrr5XO8u8LpjsLLpfkR8g/4zzhZEKvb2AwndJJVpolakMOvhNIDrdcjPBVJm8/IJie8UrLuKif
2MqK9LZ2g5DfHWqbATeq9snps0CTYs85VvfxzB3I0F54zujMZLCOcCijVYYrrhVMbCoN2OAVtoof
NqGZ51TghFM3s/AsPBIYEebtAGrmV01AIbhdUtKF0Y0ae4jzq0Sn1VfDxq+XIjNkrpKf2jsP3Dbq
QH5N6rixSTIDr+5EPDOxBNqSC8WuEcfJ8cNnMnHBTV0VWidbBgn8J93NMex5BMcS3XordQ2/XC+1
vz6bpYzMEklnHfwHRBmXmjiDyyRzIBCdjZDWfBF+8jQkwbfx5V1AGq57Fj3uNxEUTwHnZqiHzdqW
zS1D99LPlfbNPluruzCucJsha0kN5zYPSgx7DaWSdQi+7RZRanpUNe/kIG43CFPhcvwy4QJaX8yz
Ic0NttZeTLnOeOsB9pDKM01gmBD8wb8O0IGyl/+RG4jRis/hHU2lWW0AtaVoGkkQ+EkWc+cQVvwc
4gLOjZPVA+kDW9Ryh4BkzWM4La2PmKI4c5z+1qHe2VWCpu5jdRB6zjpD2nWdZCkw8GRN2ys3AS4o
C0OpmKTzVdZXGdGh5qM16K7qGVfvNa2rj6bXTFGASRs2ChAHl4+4r4OV3J5PPG3JP6ObxLdjWvUK
vzQHrVO3YAsg+yFfPc4GNCVB4tIT6SGc5bUHheeD7Y0KBG4kz5nUtdkS6nIgRfTt/av2LwVrWzqp
09bq8/2BevYejBbR7Mi5t4BV4/pQGTAAFG+2eEiuT1J6GYYK8/SWeRR/V4hZobP1yAhgVnVX3Hkl
7OPBnJRCoi2E9DvAtmeTekgsvelc4ZARw6vEHNfkWrJlMfNbeKtdimPkPV52huIB1kImj5H9wrs2
0MQr13zyoA66OyTvwQ4A75ihHzebAi0Ny3aZBIo6MgufRrQQ3azuftsyGJj2yGem46f61RZMFnoD
GzL0GAC1KN+aqzY4TqrIXJqkuycD8S8EyaleYV0W4iwKAu+Dbjcxa0U+t2oFzwWJzoMrfb2pUGKv
BdUqusZhYRA3aHZoqmNvR6t0eIH2kOhkGh4hwJ/4UKk2HjZiSYKhiyN9nR0v/bq09lbOx79AoXtw
fiuTUXpvURfQ8GY6HDBDHXbmMVvUKlGb3w04h3JBQc4REMHkfHmcZUnWbaxsiNekZzxvIPPtpous
/w7JajSqpVoXpXi+PWSNXPt3tVyAg3jPqrTDrMvv5NNhnIzxLbMGEAOL6nQF48RqJp/VoOH/rMn9
kHF4haU8kSsrRMGfdFt61fR0iKzUJIOqbsQQn9YAGBXl3ADf0fglZyQFuoAyJft+1mVOa6g/TD3T
Aa3PWMTJY/x+bllblxyU9ZQP5d6Sen5hi0DVz3fTTn0krNPpgRz+mOOefU7JGqkD0moGN2N7+b3M
v6k0cbouO0o907O6dwlQiMKvkfePA0Zl/bJefKAWBMOudcr8BzdMxwZsKOoZYalscuiYp9Ztgvuj
aZZCKQKqCiCrBkydp7NvdpblNOTeHsYkzk4aFu3Tp5fgLoYrYYG0hB4cYAhhJPRz4X/cOdddictm
W1HZ73o30tLQVDRqnVXWByeeXpw+Qx5ijiSDtEmmPyRv1/vYb6GpyP/lHRU3V2ALR9bOBP1DRdTU
tqn2qEBewdgC6J05VDXpPpNmVEqp1SrzQOtRzWPhjIZ2GnR3Eu5flYTXkt7OlrSaXPbEzMUAkJGL
abqmsV8+ChEhiaBUe8dK9dh+dWLeAOGa5sPQNoLPctNBPT0oWHdslBw1bDINfiEz9Yv4UiSU+ILx
bEYizR1rJJ0H3kmFL9cqxnSiUXJeZgAXf5dAiot/jA1pf7t0gOFSp0ZZl6oh+BGd5R4PCvh+dz4T
thwxEQi93ijDdx44yLT3+LOi4Z74VmBp/pzi1MDTKzaJdxi8QENUmBV95jGWTU7luIQqudsEcQ72
Q4q6ztlRW8c881530UJEqSDDpjJOkHZtETIyVyyBsrHzGwjHqkwYBM5TN7G+/SGMT4YTPwKpo3VU
X37TO6gzce2HEI138HABPxDAEMwdI2ji22GaHr58kG4c4lKKGzQ9R+Qxf8VEKJ6lzsTP0zvOvoGA
VR06aYFPDlXcX5NrQYIuoUiwUTu5ySt2UnsThLpX819ZKWlM46ZQ+4KTjBg3AKloOn7ueedbvAVz
+iYJlD5vEChuyZCbgvzc1tVDBl6w/IrCT4vu7QzdvLFJSZeMUZIGdC6k2j46lhzk/NokvFYJyz2H
BBFvqgIYfMJ0EXQtOfjU/q2j1Jxw9WNxbDW3f0nGcdwMmlLTQNjj/emlhbe74/xqoOgwFag=
`pragma protect end_protected
