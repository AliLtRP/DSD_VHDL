// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HAgqF1FUKn9K6gqSIGcm7BltROttaMCrvTkFBMJ1prS8hO5GozKCszRc68J8iddR
lXTcTy2MgVKH2WDBXXN/lX6e7xeEXTW0i0NOJHR75UQxjW1fpZtH/Wh/YDFhyJUX
SQobkr5IUL4bi/EBEQCT+HFJsNq+q4uHQJLGAURQPRk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5424)
RzH/sCXZFkB1t7JQPEMWJMSvlBWd/n36I9tu3LzmjzjUKHfUXPGr0lxQgmGe41mx
FstEAF+xAsNxC55Tb+1KuHuR5LDubUv/m7vqGxK3hVwMlWWe7LD9un+8ZmIRbE/4
3bjNvAs19l88G/LGYxMwkmakWsQ8YP4pD/u9Gq5ELOIFaLs6dymHDjLASoHvGdqd
DqUKHWB6ozu4CBncqMKnzWMKMhnupZeN9aZt7NVpedttmJ4pgHj9HLjt8tmNIsQM
Uii2yerJwTo9aWud3Is0h7r/qzv+1MdXs7x4wy3MW32vdFYuqy2qqXrMe7VfQ3y4
N5Fo51zMZAizU+1oJkzVFc9XWi0ul13amk8HhxGEQRCjJi7WDnwxHZzzde1VtQuT
WNCdaP06jTCQpiZ2kEYaNLiMjHerzEb6oMs3a3u1ETlakp5D7Fj3h/0YhqEHHrbW
LQS4viFBH+4hwD5AlRq4XYv7lkzzSzn2vF3nxYajvUuimjCaEhwUcM+C3hoH5CeR
ZPMdPmql+yZSjgB/PJwhBWb6BJoWFWzjZgXcs1HPp1QPV/3gG2P3T+kD4YW+Rfj3
ElZuvNEYPZbOY6rfxLkpzIQxUu0GJLeGT2aRtXy608g9int66oBWVBzejBT3spUp
ynqqvoAZ9LEmfMCF5+t4tNLL4wQ8URlvXyA909TgakyHvcnEvR833m1YGxedPPvc
7iQR+L5pp3P4OsTJxFIxp9lb3nuRY/PAFfBru0sjWDXZh3nVRKvUDCn5nBgIJ0X8
JG9EBMcb0dd6ePRZMyG93iU4CayxlsS1Q8LZX3KZk39a6nQczW2uCKWLlPQLLm01
FSK+YhKPGei7ZOsmcqAJFhEWzTFBPpUoVeFp8iE2W1ilMJ+3Pmdje5Hs+0acr7hi
HcARoGwaDeP4/aVFH/HOhMVDnqso7WK0+w6W2jnStr5zufyQ/1bo6RHzo7qnoL+A
/14y7LOmWK6FM6RGVs6KM4iH6g8ZmXrE2ltRAd85D3WfhsE1MAi2qawdIMkUs77W
S+HGQXXLHRY8JmyrJ5+kA/w4Pi0WUfgAnvJ7AAJXjy+8VrFSnSfex0Mo+dfAa1pA
28zi6hwjXK8qf+sM2ISzdGOJh9erEc/BNvGS4cmGsvtj60RZ4oXgHGffFnkSb2/e
yPe0P5Wb8VQfMYcSkTyQXpD9W8gzSbwUiIDKam+YiMbmd9/U/tn/K11m0QkVe6Z6
PKcGRiEYcLZi6NVOIYxaqr5Y5OkTAk7BxZ7g0kJeWjq6PBzDke5D5mlpguq+MrGS
WN+Hi80Wr/elpibnIx/vtqp+ZMndHAEP8Dng4r2Th4FBUXgopMI487D1TYT0o6+s
tCJI3f2GkaQuXVPqw+mDEYooKnNoDqiXkHAcCfvh6lXO471dQf4RVMWdsvqgNhSY
C2Nji2PqfsrF3LcYFFp3MaREG8I2p5AH6utqATGpjoFGQkEIDFODd9AqW55CeVFQ
ES2OiAcUkQJJfJpYhGtn4My9q7q7f9nUdpSn6zVPlvuF18FQKhZulmehv4XYHwXA
dvFZeHGwMGm7p3+y46Fu0sTP350asYpixJ2ThH7kLrFttnpxFb6hMHGi12QSi98m
E1ZTsL4vI/ZXMQAviD4ZvkRwSechiM7g5c8A4FlwXpwL8cktZB5qtlBIhkCaeVvQ
oGIvxAt5I9cIFytzdjgUuQQret+SE42leMFu2BBGJgpSSIl4lhbc7jGIwaPSBfB8
evgSGrf7TeEZBSxawlxJ2DEssYMT3SKFb5yeUMxpE+S6KeMLctk0JXFl++71PcIm
6uPBBTLZRonXpYv1S9LeQS0+ToBLaWSRcgAyUjhfgEMkpkmPZol4Wuk+o078uFES
UBgDOeo9tYTx/LfE6Yf0URDkZj6Wfoq/RjrKFCam7suUjU8ixqhP+wgZdvKBFfw/
A+QtLWMM2H6hsA5qsm6Ygj2ATZoM2jpYI1/W81x6+mR2umzqt5H5dMbBOqPaiaRX
aH5lpGz6mm/87uBWNAvN8BrOcNiye3q5PzJdtyyvkuiOrX0eFPUL9dgX/BpS56nO
AhG4dIBunPsZV9vM/sUWtak0Wj6/pC6VLOeQWNI/GG5z0vpvC8cvD59fSD5fGyH/
j9aojVrCCmeSCClNrEt433gmhv/YvmjXRezwwcX0t5gpgRzxdlU7gIWXKOcVlkAM
ZRFMDkehCqLNOnNed3EtIzHCClDdyZoj2vVJQeOPjnohks8Ouxo4GlWpCDQJsNV9
9HI0n4bAb9ruvXOu9jfqEJ+upgvDgOzayfT0RbObQU1b6IEZoLQhr6DSFhABE9cI
MFvcKrgUn+YxgoNWy3t1Xwa2ZmpJlHJNCqON0TxkPXYqjaHTIXc0G112uK5MeSSd
tKTHGBAaIIb2An6evKJq2WYrudnq+k2aYJUZwOuQ9oBEioPLm7d4tyKyjECj/8OU
VYDhoEWXTvWHgU+tAASKvcYydl+8EQWyI6nkYNAvh0M8JQq8+1yhoGJjW/2UvOfV
PDq9TBty09lE+dmJgTwG0bHIKk5OB384kuF90lZK3hy3e6dfr399YvCoqNDQwW/0
JsBVF9sED+1tF+WOxEaSSKmRIAmKuEnUlOvPLfpLUvhnBPboq+l6jZBrbc4SIAlj
Afd9n8/IQQn2aB1OUwTGiyA8+NQYIxtx/gV/2ZuZwsCRYdee4WUEjz26JyMwiwRD
TAryk4eOs4Lcb6brGIEnvqAcOlBur+wpbfmzxza5b5YIiCAHlAdUroEsryvwcB2W
1uDv41QZXBDrLs9cTOAf70tHOV3dGn4zU4entp8g7Iq2/SBN6ChWGgQSFV7xNOfq
Wy/PQlTpj1hHOedi6UOs4CjFLwJhhTsalikV9rXd/FQZ8q3vu7QzNT2mNCgg3+CF
EpQVnGtrntoSksPhqPgHI2x4U1GLv9nkFrNMwkYkoRmHNRThNsQspCzJ8EoAEsi5
ieC91dK1y16zHvF6puwzB+Ep0Tox8BRkSw5gitbdatgYymbsjSRss/YokYqRgj03
0v4vljBZ5mK2Jorl0Hcb+nvd4uRpXO7pBjfXKojlHqXYiPMbxDF5LKWLy6u6qUHr
LEdxqmmMUXC0Cqj/qig8vTi2u11+dq/lDgq/lyPwpvTfXeZgJ1shJhYDr9mVPls4
wepzvKBvTd3CXOoKSwpzSzDPphb8125/K4dKq6/V9eNdBinsSfu7cO19ciXyTaLZ
K3KjvfzryAOlfSu1fQiB8p9xy1wnrSo52DR1lncCrlZWVBJ8N7l7usmhoNX5Jj3g
a6E6IVHqQpsCj/v4BI/FWBP9+aPajLZfuDM04PHJAG12uMRyJ/SLqOXC0Jshdyu2
lvQMYGm+ZFIFjfzIjvCtkF71XweIcFMSF/cYn0vobykWP7tv82FEa+A4CYnFvpNK
B+bUG4KGndNpwZM3R8/V9GFZakRe0vBeQjNmEADHl4yV4p9IJE/Z9IK5GaXK4Sk5
DbgbkPozB4Ta7qkAjMq3UtxQdqi70QgYzR4DLbjub+At3aYGE9VNrUQTWQqP37B5
IXSOowqDwO08sCZyE88YTflb2/YYJKA9HgGt9djlj+zRNgAK4cmeVohVAoKC5XV8
qghWODl4BlnDg+yfaiqYPUpE8Y9kLnghKvxRD754IQCsebHRxnl5UKcWWcdAi+lF
zLY/1XclrEPmMplPcX7yUvmThnffmzE6F8ifS/YDv8Q7UgE2ZzMUBGMyfq76Pumz
PfevauvNmvJQunPP6bLMc/Za0Lo/iWKApASPl4Se+jGTdGnxdtwS9cnq4aNtFna6
tYkTJUf/AsJsVqYzLy1WUjcLnEfd1KZnIv491Pe2yGaloUkqg99PjXsuQ/JiRF0c
jCA4p9lpxniwef/7DEiwMH/XRH/rUyQ4jdip8a9XYiDTkvVlSd1sMYG33k2dRW76
7NQApNOmpbT1D0SL2tZY8T+FcqQtDW6sY18/oGTQ7odu878xqSq0u6wqPsyWtt0i
puNzD0iKR6+e00MR5WfKnSr2ehhmKsfsc5PUNtiNDYi8qfL6LAvgRnXYKga3RQ8Y
iS/WP1x240R5bgvcpQPSUpFY7MLYp4ECiHaQtzS/xkfjW6sn2Vx48CNr9V5x/sGP
bKD/M6KoofAZljbPDIvAaZMS6RAR4GqkNSdgZRhG7IFkeYg98tx5J++b1/nboqae
6u2Dej/2jc7DeEPeULokP4bzsbxcW+7iKem6Lk/gbCCwkIW65WuFdFdDDeQbO/5q
tAr+4HFOD0vIT/pJyJR/U3vLhIH4W6TMC7bdfYGbPMfi6YBoElcyPXayzvwkRP09
2u5PjaL69Vp3O31PbVzjjePcPcVKilQ3+QpJvrsFDoEB04IaaoVdNqqOKpzhQgD5
0zY6ORL+xaWRaWMWIX0+beT7D65fJI9UR0f3hAj81VaXB1ir/FaI1X4C+Z9vMyWe
Ss6tRnv+s3JtzUDJteSuA1Ewwbjp4AOR4YnPtdw4++txlnAWjdObgHqJlFYCFmKa
4f36YVX19cCg2GDGSoqGe7xH1tr1T7MesRmgUH+BMHok3iz5AdjdPZmo/4b9YYs1
KuVnT4apW6PcDCvD841Ieuahw3eYpXtNMNvGTHe9IrbxX+DIn+Rr+2+KRCENRAQa
DD03NoN/TDZoT3WMuJosqVKCr45szlanSZ9kfsyhmpIjoRNuj6aEFDpFMfbaNIBA
DAICiIFe7A6t9ZpGaheBXg2OGnT6YxA8GVPH+m8Q6lHjZWTFCMQPETgknRwiEW9p
aNTcBTFwWtPunM04kjN7s1wphoCmemCsUfvwM5f29f4aLyi84wh1wgDFHu2rGOPj
AjAu/95dtyZeFdl/PF3BpsUowuU1zuuXqMXwl/QhJnfeJOVTUGugxyYo0WvzRPFS
f2dczg4JZSfQ4R8jixf9TI80gMtAG2yywYJd6diaOXyLpc5g97tMEdzxZlwFCddx
GGPzgp71iutRytcZMsadaSUrZVgFcoD+e+WLIUpu3uSSYXflhMARWl55iKFMMrr/
bgC+CFbskeJL3LpWDeJfCJJ2XsaMh9QxTFtZncqhXS/AIb/EZzl+IvRJD6Uklf/I
EGDa2JADb9tySgtEtkvxub+Jsgi0g/+JdsvJaEvQNVxx8YVqoz8evS8Ko1WnJj6k
ZM7Atss07QqRhBx4R7UU+KUZLgKIHVF+9jNU0mQGTLLoEf55eQUm+E+mBPqgjLl7
AGzyCEWDcMEPJgIuxNvHz+4oGQwvnwn9dfEzuubuWx9W5B7h5opuDJQBTfHCEOUt
RP3aYuchvLMsnd4O6SFTTC//Cd3GFT5DweunQWfmB6lC266qLLOavbDDJGLQLMyv
NWkbZdwZAeuKf8+50PQ4AFKDs73aLFXedmSJ/u0CiEtj7x2Rrt1y/jS/mrBadvIi
l/bP9ydVNyeyVlct0r0c6/mR8EjDu8RlmDxVvw73o2iDoQeONZSBLoxcT9VBiZYU
rwjPRgENzJ4bFiTLHrGD9LRWRP/pQ9XFUkVpBQphkbyVCYVv1QPAG179GROTFnPn
8I1OOEN+llGyVUt7L0emJ0GrJv3z1HBpSsGo9Qx+Ai/3zGhPsLOpyOJ8fzbbWR2o
JEmFt2nHaHGYOWzDjJ/omsvgJlGKXzAsvoXOYAw5MIt86ts/L86x9bSGIz+nmEhu
XqhEP+6ucykNURMxDJwCw5Kib2+qXq9CLMAa48bivN5zeMgYcqMEZ83s86haJZJq
ZCFfXvG+5J8VrO9CSnPFIk3FsS5vQL3Dw4WRSSZwk2i6wU0CaIM0cwAYQDawd0Aq
n4cLmy0uWJPxNJmAURNEK1jenliv5wjHyBiv7iz2TvQJua/YzcxsAb1zarpOsgTP
nD7t8zY9TFY2/wFJFOOuqBZ5bSUYpQKqB4IujV1JUnK2D3zIWxOthb/UDPaaJtBW
ILyTC/HQsg3EtmJO+az1o5qPwuElMDVWqLgYsNpfUOO64aeqiZX0I3MkZFIvjp/3
oSjnfIS4GK0Jvku8Pa9B43ty8td9dUt09i9r58QulJWFoOeUHGCW5PEaddtgb3Qk
N6vakiDyhhM2MrYyLXfK8LdH7S3rjrPO0Ng7GocrCR0FA3bnPaEJe2kIj9nmfkEj
TS4nF4gmBVGGt5gAnW26MqY3wAxb6Pa05+zWFE6Vt/mz48nQiSj4IsMRqewnChx0
Dal5V9iZxk5DU9qP8K42/xJx7YOrhTBjTnjBQoXh0ghgi4c74UjVv3LpCyWOIQiM
gf1TItrrK91UxnMzb39abCU4J8wHVo/RNgyBBTLh/u22wiWuzWyOOphRKu6vjRoe
oCQoWP9VSvIFEJhRF/dCisNZUeeoW6aBTesBnFkkXn97P5Ewk9xuXbpVK8srJiuw
d3F7pVeD7LUP0c1Bj/K6JaGe6YnUknLpL9tCICSjAoFigJi+M4hA34mF/pO01ggJ
HMrCIEE/SvzF4V+VCCI3YmLOd93NAf21vdSvvDaqMJmT8CokjvpeMcJWQYJZqLlZ
k6sF4xWI5kJn95ZBIzjhBeF+hAbOCy7KpNuEk2va4GS0WGjszmyhChBde75V9WL5
/e0QDOK0dF2bwn2nWaNvGCM5S9K++6yxg+wTPivbUe/3KBY9LR30i5iUbZQvSE8Y
1nMFLaIANTQ0P3yyjDUQ9HPTk/dlDh9fRFlIMsMBrUg3kt5p4LWP08O8Gz+6iV+c
qVZhcuRErOl2V8/wOP9TYmbeQ5JYSHbbiriWoLdKIpyVFK5UtA/Fn3k+lULDj0fk
/lSM2OPDvzbd0zOIWJ9ZJPLns8uIFl6KtzpL9D2zh8kTwZkxrXo+v3LP7CttLYdA
PtWi8y9iRX/H+DWxd+mhQLnHCKEixntgaMvpBL57lhzIpxwZklgr95oS/LF4DM18
uNKFzBjyE9nb9AK8oXUA6054yzW9+qpJLxr6aO7GdSjXcOzQbTg4/pWSSehDslRu
E4NfV+zsd12wLGwmNzhB103CDfhVg5+2vyAvWE3m5dbks1T7F4C2x5G1FLKGCBG7
yTHRYWQPkS91FcSxjiOmUnYBp5czLk2+htpdDQ7x+is7bndCQQMtcpF6/EYgDuDf
uGGq8Xg10urcCAXX9yE/DcAMAB6EYg3GUkFmxPH+ZkDp/LRMJXNAAtlXN+tKHL2l
P8lXjBMjrcGt5+j1Bfe36StfyIP4xj1qPM7N11Kvo6xV48g8GjsfiCVGo0JZAt6a
g3U7nR0UBGD+1XNJx7jGdzsXTgcdLQxkhXCTxa8ikh+Mpn2GCftQjhMPTwgGjLQf
`pragma protect end_protected
