// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V5lm6MwawEJ0YdCD915EY26CHqXkh3tfQgOBxX6YVXlhGlad5uBmLo24DUgLxzqD
cEG9w7Vc33vcc5FDK/kx/jx0uCz3ejNz3bvV9AHZA2Q5PHddtje8ykPwV7qrU1fq
j+iHjn7suI/ITxlzgr23T1UaO6JknAqLCux+yffh3Tk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62144)
WZnSCIHQ7cOfXNZVQYGwvjHN5HEOZ/cg9LsdKrLIXvZs0Ug2oXr2+9VUzWtdCkZu
rhcO59u4zprOx9zyIcYisweqmho4a/7a8+xBmwG3ownTePlgLKgwwqoAFXFYXc3m
t6L9AyXJsm6pmDh76dog5LMjLes7ks+b/YT6c8kCvp7FL5rY+IVsvpXo3Min8Sdp
iI2n46iMCKn0PCgr+8o7OF9o0zOMnqsTvrvUcby+sUmI/m4v7Wwqav605E4o4BKl
JW9Yl22tqq/eRwxyoOOQ0qkaK6sssUVkuBHCa8GAM8ic0LrmBACQnU6yGb8LL4gz
CW5W9dWJH6eNtYUwQLL9C+RVLGgPyMKtwuhVvD3bGwo9ptKUqVx+OPTk3m16poIF
O84b6zSZBfYjPjuNEnEosRkrALk0WmeyQQWVyNP2OiK9P3uus+eIeV0GnaP7zyj8
4ttYEpFK6zRHA4FQIqu/GD5WEk0n6cZSKn5EWpsuxfHpKZEd2771T9JY79MzHEHw
6yctfaAyHq5q6XRDl0yZkvkD/y7MibaEaUjRHt1ka1TwQ+kIMnOtlTD8vNgsEvIC
WIvxoYQxiNatFn2WqRRQ/hw9gZPBihgW6KQcmA6JrdOa6zZt/kSyKHDhnyH4t1gX
69yHV+G1PMfYEqL76eiF/zgByWvWhM5AYlK/GLv4txSMAoKLA/0EptNnVIoXZp3z
Wscw6Da7wVSe54v6yji62AHuDPcEwyD4xF8aYC9w51lZgzBZv3vRVbNlMVlAZ6J+
sOXfY9GB0kN4jE+WzEiPzISYGop77IITCvkOdK61xrfQs2ISjlZik2WKYEHgMmtx
AMaEEo5RCF3Gmtlz6WwtE4HC3P/3Xpk8gg3EwwUPOCE1YaOT+IBANd+x85DxbLzG
FHrk9BS7zYbjP7j3J6W9nLOFzHcr0VmGELfAZzFeIcXQomAHeQSJQKuTqnBl46RG
bmqyAUSJWVE6n9+SqbFNMZBVcCxkO9DsDICOrD7Gt7b2yX5bwWhn8bV0w6Gubavu
PCHSsqCBBRZGCFO76aVDnufPoKTGs9hrXUqztuc8zX/3BtLdNCd3oo1bry89T2Hk
Wx5cfIUDuHpAo1Ser8adN9Z8yv9GTaNRntndz1tIFZjBz66btV/PFs+adYDhPnlN
0SI3erMkSKKkizcDtvGn5J5HomBbQlVjTxYl7yJAQk9XWOqD2gbdHxMPTUsGk1y1
2LVKMggGBE2p8zeceCYMMch7UuSZppCqIOCOwkzd8JPnx/d/ZhpoSw2VeCEwqDob
09gO6k1zWj+s6CZWDthB60GOL3k6qE7HxkvimVNdeMjTXFnKrQrfL7CBbfWeFLQW
ZyYwzYHbS99YPW7vk9+f7IKfXc7ZwLOM+wmQrigl2ABNsIbl1Zugun5/Pe6U0lut
+vVdSKIITzWGjIaLGP/dwf00WqXPbQCHQHM0UNXMYMGT91KbJbwcXAwD56SfETpW
qJFlyxW2FszyT8+n1NWdqxD5MI0AStfsUNNq9anM8oXqmKVkGLDnrD/dKqvhFHMd
8Hc7X7roOPqxjbOZ0Kw4dfR/uNJVDbT3EDKIDWe7SroGajaKrqADmkY+S2exdczH
ixcxOVrlHWj6a1vF/5RaabkJoxVxUZft1lihrb5SYFs9edibKm4kxP1f2PFTJ5mx
DGSLCmf+l/j/EHwP2F8CE8VV4ZdkBxhWNA0R7MIMUPDZe7NUBQhiGIC5auERoDqd
3Dk/KDiQH72rNv1mO1ek6/2MTQ0i41FAfb/UH2Ywe1xWIIfrvnOt9dy3Q/fur5aT
b5VpBc6nm9aJllWs3gE2l5+vX9Baq1I8nUIhJWGQDI/iAVsHk+sfLgnoHamRxsxG
V9iIVkhOZtCvblhKXMtDwpwbUI2sY+rjBVh/B58K41oMwzdguwv14lofA4+zDKUq
cfg5tR4QPygP0SMoyBvyxGWURPHWgYbqc2gXKbpmd+/9lC4MHFS4sLe0kjvtIKWi
pQcztr6psOem9apW4XkkGeZYy3ofCEQgvYfUKXeZUJbnBQ6BA5NJQhi0jiAxbHwt
iwlMTqNnBLnwfbls0JrID0sqrdkm+wZAo1y9+fOBmweEwi7fWiGjucLhwEmP9oZY
TaghYCZJOglMjAZGwNNopeI+3wDVuUG6vh0jDaJL7UvfHPU2wtdVLQoRZpcFR42L
CryY9uZ9+wR1adXBmg7XYn8OWQ0gaKMKEuQ1P/+NB7xexv8x8j19VhPr9PB4nr1n
004c+IDMN1vhEB+g54EFZphsaAFYGMIZyA7/CFmBShSNvdgHICJ0w44fzGafxYoy
xPZoktzm2MtZh59ro2jPxHiqTV898NWWI6AyX26toRqfu/+q7J2IHBT3NUC1/sRM
gH4+ZDmEd4kqirxcdNg6+1Q/JFooOEZpZ8tIAMSWx3ZXLhMDpidgdDwMIf6FNXmj
w8gRtS8vRjSxIPK3SZkDdbk3cLxbSPFATAOq7fJTtcWjWoAJF28vqv7G1hSqloVm
2/5Fg1QHCyrsmbpAcFwhiZBY9xVhqBdx3mHyPToze5gswdgSnMPeJHKJbP8ghk2t
URs7TJZBNKb/ISQWOocBj139gJkC3pd6eNo1DLMrFyuhvQqDHjurihj9X4QN5xDH
h88SufUStd8UbfDkUo429StBZBam46IMoHkCPqu6XIR4OOiock7ngxVNp0Z1NNT9
vnke/pEUjjqGXyL+5NOCNworGgfkKHbjWNL3lBSenvGXrnxx/iSkV+JlZEgKUB/I
ZQtDIlndNfK3UDkohxP7coBZQEexzqZRrn9hD80/lAxgdntf3ApHssQ43cjQYp4S
b4Iiqcx5HSDEC5uRiKJG1uBSxZ9fnx53VsWiz5WjAOgwPVOQBJm72X/tsZd4FQmg
veDZrBEvntOb6heMIDDiYMOMP/3BYqqnRYuboEl/bB9Xti96BWSb2018ypzR9ADl
YZYJaDmF2JEn5KcyrNUkN7l0aJmeYKGVgbKMBYEDL7F6LCEb0J99MNk9O5wkLHWm
WZWNFd08YkELj/fwVqWLcPKHtbHN/FuhS0AyN4tklKnPcU/OKuN11qwQtSRuRLJU
tMAXRBE+YqwkwfotgNRml55fyEFM0jjfA2kSwXu70EU1AgDv7h8CdLMe/KhDcWjo
I3N7x4RPS0gW6LLe055nApo7Ld49J/32QjVKngOsRMQhid3ChxV7zGqponnDxX40
9f6LmxBJv69NWwlMAWFSnrMq+ZULEA7+HExqA/UAojivEtd+F4DRTlK141KS7tcF
RoJjP2j8lrfkciEG9c8P30wvYYw3C3MDCyfe7ZLMMGotCgscWG1z+GIc7RLHvNXW
BUFNdurcTaCobEAfCTCHMvnqwf8BvMlh8hpT8mI/fVbH5Jky66h2gS4lUIUtoUUC
tXNKZR+YZ4JXOXc+yUnKV+l+jstcwU+HaC9GbuG2FyrHVGefG+CMIaYMhbNFpWk8
FfYprz1N4XlSpMMARCpxang7mWab5OYjNTc+IeJBf3uzpX1nXcMmiTqSc3tarQh0
DkqocSF4pEfzzUvCT0px0k11iZRweEvftBhQt2WZFaotaImg1GyRoloB+dE/9ea4
ojzozjawbtoPBT9EqBVv3FhBtv1DOt3ru3sDIcjfFK60kkcVQFp84lEbvB3/SMuC
GXsE9lEe9dPYIdVKCl2khCZDAVM3f7iwd+L4gSk7/BrBSo/SyNeLyGdMAZHjyEDn
S2SO18y/7BjafqLrdgu0InhPMyXa72cp3Y3FD72ngTiOa7MOnw2rFmldMLgNIx+A
tXK4AuUzeMCsJ0rIAmA1LdqCM7RvFDyjaZgKnviI333QRvqGAZaOf7Payx17OSy7
FDBNRnxJgrc7HWd15KX99aj28Fc2ZQ6YNY+2pE+EUlNR8Yti7vXCQyAvy8rV3KM3
+MsZd1Wo650KYZM1FI4PeDc2xpKPj4yPfC5VqzcIiAjQ3etZVwJvG1Qs/wF1gRvX
qKjMfVMps3in0Wq+3NLs3LV8UcSNTQRk2sAEWqLXglxOmtihkZIWQwgyJFHw9hoe
2UvrciOvXiAftigsoPastOFs8Q/QyCiOcpcRhI/ZEyFbvc1gxiZCTCJybMrp5w1H
xhYbmyFxrkhpSXaSi2lZD/0RuO2/ZUc3HuDO4erxBpQ9Z66ke239/lLFG3B5E+Uc
z0ON0EjepHy7gIAJH/hhyY7IPoMgIpTqsxLFfjJcMUUuzI85BGNwj5S+FS0vfj7U
EQ9jpPZJJP+KLbzUuayJBcK/5CXVWNT53SlHl4s3h/ZqfywjAspwq/NkAo8RICr6
n290445t0BesYSGU8ToWiOVkJnEOb9oI2AwEK8FOOF1JfDClFYIKkaFDh04AqskU
4HBCUj5PZB0fzOYIwh8uEUuchz7VEWWS4aKyZBk2lPuqEM7WrE24g+GBvT2XY6sr
SyzhOKFwgTdfaGqQP5pwnx2XWY/DuXwgme0bj55DXnWnd+lt+orL+WYqfKb8giIc
oK4dwHYC5pIaQPkrK8nWJpaFNB0m1DVnW0SXO2qTKey1d6gAxV3W0mOBgFploV8F
nuIpOSrM4FGaxY0SRlQDN1ezC0sMdyDgGehCDAhhv5kGYIDY1Qe5Z39KjzfKo7Kv
5ISMVteIBUTVsR8micdw7+DzU2qAEitfsAYLrz8jOBRaXUyjg8iMza5asGSq1XDb
uSfA+ptD77VxE9t5Ag7cr4NoTICcsURaTQJ4CTfTVnYm3oMp71ff/L9Lfu/RUgXq
R6D4lkPPFamZBMi/CxpqYutyaNByO9sVdafdykwjfmGkGH2y8xUwRIAU1oehtqq6
1V2JPX5FKB7C9LUl0QxsTplWojtF6uEEUKwNNYBXj3B0wR3S5Xnb00BnqbOes9EB
DOIWu4czFwYsBDPqGawuaz3o5MUKAKWs1mAaHh2J/UdjROvjhVAVLk2mz0dSYny2
Bfrox7BBaymGQUtptfUGXUf3ZCP6Q1lUjGo5Z9eUDV4j0V9GzbLkarUue81IoVxA
hOelwld6uVRQrRIj2h4YHox7glm49ueWm78j1aurQ5mLffEaXVpA/R4xEHVCGcOZ
P/kXNR1LxirsBrAIi6f6Cg0eU12evbEoJglZovT1wkqSgMcdh2cA8JRnxak/cPdj
Px8i8aFe9TNOylSZ5tWkj1KEtRQSTeEE4SyRDtfsWkZJdMaCINVRP12xuZc/NQR4
T4EQiXe/J58EEbUF/49Lt2ZnP0CHuel1kum+5nhgk9iN4C788pYslxMRARgMwZFt
NVXoxcucFJbrj4tMJ/8Q4iTt8RJxI5mBf7aE4rjv+8kRkDb7KVdw+Mf8uozpWDIT
xvRS5COHEf0t2fsOc6tYqzGcDeVqRuO5c2BnH0XAhlfS3sGdFweNhqVWLIQ86/DF
1uEWLvPcza9+TuJEWMiL9igJkw3BJ3ug1nUBK7PtADKUfQxTTDoxwBLDjr/h30Y2
ANYiIb/N2972sh0xiBFMdRZHo+yH1LvT8pEw9PqPiIKU6L19U8XMcUnbCNCrLE15
5eZD04so5tKjrVlsqP37tEBhR5jeXVNzbkFruEr9L4dGhtGY2cGfMW3hV5yJrcuj
I8B7LHXn2unLLd3PvnetHgNlBmD8MLQTESWrJz9VsQkDXXtQK6UTJ36QpLU3H6in
WuG6jeH/Ee1htsn8lFiiRe5fU+A6W8uzj+BLLADN6UcQcksOMlft9q2FQjwv2e2h
c64V0r/9+eyq+d8l7tDkpunmaPfbjY/QV23YJGNiSBIRYZQLUSFb54m28q3l3VnD
6Lw8DF7ZqgqcFkvUvWnRwc0BDHHv8o2tRa7/c27i8k9EdVsatDVGnM+46YTRPyuu
ULhKFydGAxU+x81P/ch14VodMjIjdgZ83VyZedlC4kHy+1H7MOuhnEr+dqDlFaAI
lwmxF4YZemFTK1mYvgeYWPgbjMLkJ4lkozjlGG4j9FRBoxX7B50J5FQHtGriNezX
HShQE+AvUJysV7OCpLf2S9B55BXNKOciC+JEl91DbpVVea3V3YWQd63liTKOKC2T
gOZ603RluBpdt3+x3zHraIg3M27rY+PAl5Sg5WFfs2x3c/DnN9tKpNuoRWZaNoMM
N4xlVx0PXsP3xthSCHgSG1acR3WRpgnbE0mxqVkiMnhCiNDyNHQl/n6Mhr6XUTan
TycE6Nyqojz95cEyydA1eRU5p4VBQ+00a8Rv5OJUkEzswWHJ/Q4PnAweUEm6HZX8
sO2l7ZyCp0kORNoIysTGygaeygvppbJLQaH8u9Qzjqc4miZKUnPv6AX6UPeSRGPC
RAroMuYLercFHVpHsIWld9rUYichE4YRpC1hApknNkMUWO+Fihw1fklVkDh5EmVt
2RLjIcTTwiWql52GtxYqgNYrkdC/ln3Za3T0VrC2nPckTcYXLCRZLt1AabhvXoXg
h/RxBusC0BRqyrM+OjuNBaULKijQhJy7/BeAsX4FEOumLw1qWsAkd0lK9iZQvIS4
Ees7jy7PZQxceibliBLkg9ofoAr6RU9eobygt0ltZHMfUHkLCHrGiaahCCgpHSaT
BZiaRx4LS8Wr+qzhaksaG2U7qhLFztI7wNGjLV1DYmbq3069hUJ5AKiQbckJdHJH
H5L9+OlY3AMjE3O0oOPddiLtl2tQZWZiA+wWiXlcwZpi4IueuSuJxlZaak+sBh9h
LnFkiNapUP6viSTSPYyYed9zp8oRxLHGXqhYm0TkA+YrZUnZ2UJyGMsmi0OM/2to
7aZ0BXTT+hkCsDbONmzT2WcK/AEzFjs6wGAjO0ceninyBi7OLfXnJZ7Mwi8rnmC7
kqBWGRPtXff/kwfM1KEIxV9gP8hNFUTxTX57ArHr7EAbnAzpItrSpkLAKTRc8r61
QpzQzR06aJ7LVkh0id4Syrt43o2VxRDcV7ItzTWwwy5Go80OgAd3FFBqHlZCkoxT
1LSQdTo8qF7lENsglm0XoTPIlLU0VCFSWeeKNQLNJ2OGxcmaZrMaVqoNmNkvOKJv
rlEWioOBkI3OYhSWCRSjmhI2JBIbW3JMdCYJJcpHzDys7B6cIi9VktcfASQdCvu9
yTxC5bUoRkkhYaPZ670sDDNRbkm+O+nRrq4v6e20lkDIBeEgFCQuEZA2ZjskQpQn
jfJPi+Z1JirjP3K4y6T5f/PpL7KOTTqDbHgzdrOQasnZrIkWKetXAFnyeU3UsL9Q
uRs2uJcPFcKxErrCyTpQBDL5xOUUa/v/9EEroYMU+pAN+dDA/vocFWhEA9lVE/Eo
YC4sd0NCtpg9FEGCHKWAZUlglnA3SaCf2pKe24N/gWnJhzHqMOqM8F5S8Ol+ex9X
Er/Sc96SCSpKfZBmY69yuf0Pgu//sbXsXu18qQICHiwCM19FWQUJe8cEktEEIAVQ
YlgjFrEBN81Shhp+x3S9peqyDwHgkODBmtj/PLGqPqsaaKNXHRP8vBEEqY7b6zoa
EhSEgdeb+fKyVNz7BEWkotW7R+Km+xgtTsRUKku3eLm0EDyOVJ5pI9hTg/GFEWbx
ksfp5FFvkUVtrLb8EUOJ6fSk1VrUBXxhdJcwSEp3CFa0QEtci4gPqrBxidkk9YVL
GJsBk2otMAR8M4kOgFRIIzrJJC0yM9XMPlKZ503saFywgodqGjRRpZLz+4gTfA9M
PJwz8LLoh8C88HNI8wlpaMG2dOBn0G5w/yp/Q9j9DA+EWlhx3LjeZP6UfNTPhBhi
ZBKBb3xIH8dFUaKnhsu1HZAACKxcMW8Ka6suW3iq0Sh3qzTjYNkEvFp0WW8LsZ+t
YcKoRmxJD4Eo45dPfgYUsXqGQMylmuIhTqQEYvWGjyHq8rnNF8Y6Zg9ksoOX3E8M
XZOpaWsma+0u47Y4eYpzVfjhhMbRYxMLjUgfoOeL2fgA8/xyITn2f4cTvxRrfRPl
RKwe1zlPdcFzJc6pcLN8ohLPbQe25iggOFmoOXHCIKRGtu4I+e2iS+6pEZRmoy0m
Ou8BmsGojQHYQ2yUW0+bye8x0g6204e0FMRAbZU12RmmV/dbkR27PoPaoefbk4KN
68ZYl3VCCuhxoqV8C6gb0uO+F1Gen+Nbsx3HTGclOQmfVEVhkSCY7gItJYk/o5C3
xUO41IUwC4bEQL5jOgY9EcVZo9CUGgcGl4s7ClDOH8JNARktbe+mrj7Kq85HO4nN
aLLcAPDqeCL6UvYp9pdQXEN1/WIC+RfyW/pT/W9WMUmb7ull0mT1KBbH/2afaxLH
0QQLgB0UrlMOZjmLNZZB+hxHCw1l2tHa7auOMNfO8EhW9TH7zfPjpv8D5MGHGHMw
kNSeQaDDcjQo6W1Ai9mqdD+9dGYji7MAj/iqoLIvaTQLUWA72PMCdqck24Ix1XRV
5MSV4Dy2LbdzYqtPwMENk0miR0lZQA2fwRvahgPKAOl/FmTQnBjod1kgEvgoAUC9
dxl3y9ebXUq8Rw++MJuTJ/holB4mYXdqi1TYAABu4sQtffXzGGQjQQBrF8v2Fr5i
Krmm2rHNlITepHmM5Fj0RtGHAqC+QHYU14K+Ug7HRXr+z/cKsKENtK30tAbQUZ23
w+fziWG23K4iTx0TcisIFOkxW6S7IFxyZRsM8dceEgLJ9yupiD+P7Cfmw3plgoC5
rOXTnB7xZr2z03tN7wVj++6B46yuHgWQa4heD5nUWJgAZmQKHxPJ2uvNdYsYsLdA
kdn6YsQvaRxl4PaD8dS9fz6j7CSo7ET7SsQVIJDpH56U4wyC7rANSrN+ErQwUvCi
2ZtieJsr0t19fPrG4rZ7uVf0IKc4UDSz/tAe/I1YxqUnW1U7nAN/HDDP1lq0H0zk
gDVlfaNlAuWx1sizxr9D297CfuV7NCdIwg3OxSNmYpmOOkf4SsWcBdPFSQAEywQ8
01RnNwOlMzm55Fh0havVK7viQV92kofKYGGhRh8/Sdu/rR5N/Bgwpv3Qelt7q2PC
QLtBmVp854A8PBOscC2Nv1sEExFz9lRqNfZA/GMVDNcYY1/7K2a6oqYSwm6N/XKx
SEUiG2IkI1jFl/1rpHT1O7jEYD5tCdY3HCg3ZhjLRm6uZX37KDFkE/R8+8GwkoVj
9utb/L/v5YyTSXEXsEE318ukB01SMR3ApcavD5Lo8wzlpg5T6NpvNfp/BdT4KpJQ
v4QRLPaJU+1aiwPHBQdg+nag18ErEONDXJoyxi1sXXa2mjbtn5iR+Iwy+USATkgt
VcXdI+A9AarQn27tbH33C+zCWnOLp4BETKIdyoOr5pgLMdZCNNPM4aAPFnF6cR2g
PCQYy5k70tSM21EdaDOGlIRiOgRrvtEvuK/qICPiZ/AiWSQQJIiTYdGwxezBEJiK
IYKJx5M0tO2fMpmTfuoJwrhb7DqTy+NTZG7Pcta4RhyVIIdiMHV83n6AMHI06HNy
eTrqS4fqbF90VqTGli+FfuKfWScVa/rOo2CM9korG8llH/cws5iayyF0WMFhIX2y
PaPkGqmRlLocP8lBuKoQRJQZd/u+7P+sXBXbI2Hh5sJt4OoT0kmN3ErKmHnogO7r
ngbNEujAO2XFOTLulAcTCLVi/aYV9uIPLyl6H3KwqsWhm2PuYk88+7EICv1WY2cb
RowjbyuKe60CyKyk+Fk3rV4zdtkxBYvBaSSb5cfp2oWfz9E7gAl9y/CNB1Sll6ZF
Q24sT2tgHNjd4kul5KNGkEfM3Z/IKZC/zJivFylr2jZFZg4Qa1/AcFRzk4llSKfK
U97a2nC2zOnRA8M+v9pLpWbXBywi2J/cQLx1zKr03VzMeAdk5JDa4vNq/TdFu4Cv
+4TjFdn2o3r1Ij3aDH2IsG8mZpKsymC5VGHvqG1AX55iPXJ60n4ZQWTcJgzuOnyS
RRQnHBGTdG30yw3GyIVxNYU9Co0VBCeXT1KRSCG6LHRsJbutj1Y53XTSfE2qKZN5
0N1clQy1VaHrigckMrSuHHgALqE6SS4Mf2mT+KHaFlIHz7zL+ADWKLcB1V3U0B6T
PnKELqWdmx9vITefSqGCdIcr3iR/6WLqzh6HiPYl4C0DQPb9T1KnTJNP6ReyMXt5
5yKsT1m/zxoUkaSsbvmm+kIHa2rq7QIUK3BK7t91wYlxf88z/EvoLCMWNc0pgX7E
08s1mg6s9Q6w2VLoVz7TmRvW0DdnVvkZiESf3Tc1UPCobdjIFM64Sl3oSDGMYz2Y
Dc5aG2wh/COwYHe8oh3NaOq58VOiXTpEdmFREsktFPuBVfKd4kdRVoCZWeXerB+X
T+SEs+dLCR1BJipJYeSfNLBrTGypMT1cwuEjxSh7R0cHYIElOchc2gHp0OVrHtMQ
wAYIyfuvtNzitW084eR6dmpj1MpWyXOj3/dKsQiWm6JF3HwXtVG+TlGuRJKbUrbF
xa5PnnFSOgPCt/vXBTtBL3uah69k/HtSzW8wApNwxekMIJawqttGUCgdDnAWs6Tg
h251Y/6U+StoeSE9UvO4p/vNRdMAhPp6GeHOEOddUmb2HT/P+MO2ToxF4dfqw3Fv
XcdbP0jAYBuFDSbzAlviy/0/MVqTAdZGEEIxBTOjZoBkmAdnr7K5kz85fFqrDgMH
cMXynhmy3dfMR040f24NKhHFDzlweEVPDDsLgLfOOcnybl24HUUj4HwPLWTD4Pv7
6bP0EsJdDW+F/wHXeb9D7T/q0E0Qpi+duJIe3D4ovNzB+ktSsVYexNiWxZyBo4/Z
5nsVEq/HijwHwNfDtczKYA/7XVtf4+SVETx1trVTQ7txNXmFeW78PeoqZCxT8kcW
mA3FOdAw4ByB3adKchTsK4siFQwj18xRVGLIm6Y6YdTaVpOIcXpoGpUgPmj1zrzI
SEMX6NXdlmf7HsgGueKTDoGXiGvR0DX2ovzC1UMGv9WlvFxtnAH5xSs4qt+H1iRP
+32MEshb+aw59Zmo6ckrzJenyO/qfk6RDsqLjN83n3RNinW+ImpIz7is6g0png8T
lVozls7zPvhufDGmJESojJqEKAjnoTGMfZ4MxkEXiq7gfSrlWSvM0s9ij0CMDCD6
SGoShrnP9rVqd8+1PaB+CPzgHYw6swE/KCrZl5vC8qZge5IsPQ9pCg7756QYOr4W
ztfKGcRERj0cM025hMRvKU4VKW9gqxFYClukjB21zRLOMWFfAMUleDKt5YvcbCE8
AcUQj/o9fo7Emmoyo6fY8bYJTH6RvqtuM6XYmNZWEUt0iYOZHENhD841JuESTDpF
hBlq50+hqvFQLXS/3KDG3PyTYz7QAljtnSjMZFnA/smvr2amPNXYJcFrx/FUekFJ
XUPWTD0h/gVucm5zFm5TGLZBBcTwErYOjy94PNJbFwPdiF5/aVnHmQhBWErWp56D
J/CGqnsl5bFZ4dWz4PipvndV7OkGIKDTDQkt7c2vPeLTVn4si64yKB+2D8qQhDvL
Co0XVUuH68hO76qMygo0c8igx7Mpnf9TU9X7We/CDSV4N3C1ukap2QT0eTdtgGsf
USeOgxB7DL7GCBORad6aqrfGC+DjCzqf+yIUBbPvTf9sd7/85mDi2N2yDv0cmEig
1nQRVsKaZVOAg8+PYCip0ylqw1S5ImJ6J0f2XUea3QDORJ9n4XfPL+0CvKplKRKM
m15HdBrWwVy2E0IrVGFQdngezwFs5Qz0wA++Dp+M1pTcNJLSJsjCew6TMctHgEky
ZsNa+tr9/+hcowHmeCtOutlg8hUUAFZOEBTKN2qqlfzru2BinEC2zk2eBvPB99Jv
dhM4+kaFJfhzoD+dtFurYuOWDgp1xipip5llAw0ppL6d9loBuyhyTkP2zqgHTi3s
R9R1xplN0RZhnR09+DIUfIvMbSDPxE1tjSwfXoN+6cBYOxFFQ7PQoxDgbe5LQM+r
9sd5EN7tVBKS5WQwoeHdnC8FjaE54W2qF6nK4JDngwLXC6J5x5oBG99gdGbcFGcX
rsEvrg2Mthds+XR5fugTzKIPKkvv65Nl1d11IqpZNyfx/JMt2HmpCHBD32F0U3lU
xkGWG3hgy9Y3O/bvk2n0UbkUBeQIDM3Y4pWPL9hX8VdVSZZlbmrTo4vfLVel+4EV
7ysye164x10BkTUH/163/Zh8chkyUo7r3wuuYfN1JIqcO/kOB8cLElJbf04l+QpC
UU+AVpq5n3Qd+rP3huccozeK/uRA42AeDv6CXwlnoNLiJ5zdmiTb0nQP2UjrvJ+o
xt9Cyq9zXEvoxMUjzRY1d2TVl0pjf8jnl4QnyB0IYPneIYDw5GDi2wsmBzQcJxlg
yd+6+in35NNoWttbPBAHDbRU03OoSD/dZmj71yYf1AALRpIC9rXnGFARuH25OKKd
SBvG3Jx+rlsjUtX9I5F/eZminRESmOFIWyDjOVp3JHPGS4w9Ojfg7e8+8z2MvwGz
9Xh1xS/GmomvA5AnSeKVLq/MO+6F2FGDemkgtP3YzxVNLVs1f4OQG8U4AvBw15T2
qJC2MXEIdid9yglbGP7hjzc+OrmxngHJLggSgYBIsHEB2O6pCNYGWrPG7jJsQfpv
hzfEOsCbIEeMAeTTDUT8Q90bqg1ZQsVoPzJZPggMCvNrtMDXz6540bhX6xqDrqh+
tY2FB5SQF1+kwzyi749VIuR4sA/ioOEHVunFWM0yUq/dz26vPRHALZweRcFDgbGN
DLOUM0b5deNxtge1vcrocqvU5x/RpEZ+SWjhjymTS7HhOfKQPBd6eawPeaLDV7sO
qgJYO89ciJU7sriH0sQMc8GoqTAqMrLEpppwhX3T+HDV7IXGMbggxIZnuOUnHtR+
GTSnD5b4qQZ5I9k781VTU03aXAZEsUY+CVYATi/zRlw78sc6gp0IZKWI5s3WcerR
1LKjBU04nnmHDtfeCljo8VQ9kZpKjOjum8cOx3gDCcaUpTt7h2ctcRtg/1MIwTJg
2gM97ffWrBDhmm0QIMnbv100Jqf6hAmtRslfX5Ud8GBKehxx81vqdAqdEsbJJcPb
eF4iIlbvS/6H9k+2133AeGykt0+l3X3+4tW4iBtqGVjlTt+KnrRWy0hJ2Md0baUl
VwtDiqP+Q29bu9N9aKGliiaZDVywMUV1RG7CcC1AGQX4efolzO7GTSKzU+zqNXve
QytkLkvFqHIW+ruOiNELLs3RA0ZDiPbSs7GMSpS4ImQd4/oREZllM1qXASHlE/4y
hgzrfEUwISpKUQ2s7p1i0EAKcN47y+Uwfzmj8F0tsaWK5Pg9t9/Z3UGMewiD13ve
8mO3QFMqdmZ3CXv6p1cdArOW2Sgzuk8/dDhXs0yGItJjzwp4JP4AR0Yyco5ckqCJ
TuIGwp90zWavFmWNRdOtyOMZqemRxvbBo7aHpPb7ZhklvYyD21axk9dkv9+ZdbtD
qfFGF3cvyy1XQNhhIfJVhDgXeiKeLDsa+PYVJysDw4qWmOLG760DOjPn2GiAZVx1
Jd0xcChGhApIrLflcC8xMkXigPKjXTi4UJkiVItECdCUapbKvCwtiU4aY1GUbdzB
LJfo8r1zrSuHEXF9nhfqxIuUF6L7TkmQLz+4uN9sAegry3iLs8yy9+R3aOnyWXb5
mNK5NpJWrPX14jR+MktKyfyykEHIkUQAY++X8Znag0SuQV5GOybDpeLSfv2GnOKc
vo97/9XkEfw+Ileq6tsEvCzyHJyzLkF6ueuWhH/RvTr8iBggHYD2ug/FbG8wD+f3
Jw5McH8VWsodJatBNBn0aYPS6UOr7zWGg0iKqjhtqtHR3fGtqdNpgoZ0h7VvPV39
dZrPEuPJho0CXAg0+uwyxnsTpyO4faeVnlKf3XjTb3mTNrxRGhYnfOPECrRoBBp0
G9OFnNRkin71roUtYDQU8uMR7aOvXR4shhBMUBbRh+RP/tScV2f5Fgmx3PEmwrty
k3KrLVe0v1UagPgx7Tl8R3XvL20O3CBjzBB0Swe2WjRnTgb/DKEbWnrfo0zBk4Xr
yVIm5XQGzrljP1M+FyYiZsYPEW0CzpLR8oA7YmsTec6X8gGBAvoN0fASa2WmYb0y
f5FY4tfh1G4IEcST0wlg69d5i3i1ab1aZcYT7AVrxIXDOqb5tfqaha5rN/eSu11V
jXuMbSx0k/tamjH01L6T+dQZAVg75eMCitX1zSA0DanMe36J+w/gmkMLsB3N+NLs
QhOy+ijMHWVYXq2fuGEFbEdCgfOh9o5he0G9RDRO+JIb2BRicO5yzwDUgNFV8Mhn
Sv8lf1+9kmximoNcaNZgvDwbg51RkQMmkrKU24huQoYhTYx73H7UjQumcJNHT4sd
l4RvpBfxu+7poB+SDGu3h5+Y/gEhx2ZVKFyrZ07+x5ACscEztmjc/ibdrMaJCSaZ
MGJubGMk8p3EnmNdFccd/hSAxBsLUBV6nrSmWSfqEIU624Oz62sSPsHV0JxvRss7
dTC9jq5VA9hgn+qvweIP8DMDav+0KfjfdY+5uTwch+BSB9g+U7RW2P7nbAejOn32
A53fKc+UP/2HB8KOsGeRZtFOrGq/U9M+Vh9yhWtoOrXzl43N1q2qssFxLcvQaSWZ
F/aHCn5I4ax3DeLZ0ZdxUQLdz+yRq2/bt6cPoZ+OsTwJA5uQXBmVL/RD2ZLeXpwR
OYPiIw/uS74qKnpTeZ9+QI+Y+Om+k7D5n7RzzYDW+I0R1ErtK3CNxKqw662LS7gg
A+RpXcKeq4ayBydBzGlVMR9SNMmQ9AHPgWl2+gzT1JIwOz59NRM3Zqz98lypGUTk
y4ob+1alj0hCQ5qg2UspCmB9xEM8GhBKaLwe28K9Nf2JEmc8e+R3r2d/zth2xkIa
8KDzZczUoAxdMcb/xwb33OImGRtPHE7ZTcS/TnyltCpSHq3fWIA60mTYTv1tXDCa
GTa9yn+E2XMs54eCJ0qNq4Q73cy3BXobkSeaGXHoH1kSmJm04M/DH9QkqWUGtaLA
KRtZ/ZwYSKNeMWcc5WDRHK+wLOo5GncDY0lueFg0qFaX99Rw1UQrEgTN89RDxlmZ
MPxPdK8ZHX+CYkw/xe8h7uY34ENvNsW4KdhQ/T1sroXJOhvqB6hidZ2rfhXKVUrE
hc/o/q930RxBCOqpyuZBPjTkjYeFMxPBTrrJHqby+cvSdPmTvUKw6zf7fO44SQHK
oAwW8pxz8v0tyHXHBNmtjlZBc9Saq29uYC4flfYtXCHRx4EagNILJ4ssir21bKkt
4TmkT4jc/TZuCzGL8WmfnRbxYpoVF+HQds7j7I6FUI4AXrF9E4ckyVEvIIyuOQV9
Zr6CHk1yh9en6mMWl04+kj++z3pfwUxqXIRWC1ZJ0ZhZQLe7DmByJctDLJTi9xpK
R5ar09fM2EBefmfg3JjvcOODAHb6JLC8lQ5oBUhvME8QI+RivDZXPwsWXepzHe/r
aNflyt+vs2v+D3NjlYX5OnIhfXdQsvf6UX+2bR6nx/1ESp5EzaK8Rv+zue2uHtce
C3cLGuFAGdrJLy8BmOU+R3q8XxmUAPNoAZi+/7JSxDWYcC2Iyk6BVpSSzpclC2N+
DlMmQggDfbKyReIWPyFeWYvnfX8nterhB3KMYM5jUxUBvtP9HfJD3oWhLVPM7cAY
5bxmbLpmUxaYsLPfICox7MakIDBFiKqgJK2+OuQy41xW3K2S9NoaGluZaYJI1Erd
EHjIHjzUbkL5ekIHxjH6U2YvWGgB5ruY8V531rZAj4f8ebUJpkId6L9x123OGC41
ETqCulmqa3mfy12nVUlrEbAqgFE4uAlZpAfs5dSkFp65r2JtMQRIlT/GSIn20vzI
9CMFkct348L+EDpSoFGudXwwUuRXdpKPs9fPoUY+KNdsqdaNloEFVV1qhhiG0l+N
r6S6Kj51plx+PlBf0nW1BD5i0qBIMQdgh1YYIaBn3MR+YIYgRR3PacoKCLpS6J5h
5+MwuvXylEVgDgpBjNVYjchs6Z59aNZ+YUePXm6dQ9JGPYo8IUezUmI9U9GDKd+B
zTBoM7jxBX/ZVp7d0xar5OsLTPbgQtnlr2+3RQ1fbRBVag63iBsLJuy0lbHyaNyT
X6mnjLDCJ1xaJh4pBzWg4IkNdVI9vd5Ro6nGYe2+nCny31TFkS6ste6moqdwWzNA
8/QAElvmBWgHgFrwNmmrPpMkOruZPruVMjpcnAeXHE+eTdJEhHQdEyy4R1jsdX7e
c75FrILAlBbPxOwiSOTaFxkuS9OXBaeMKPYwH1DEBJAZXCDbVEiWYr9lH7MSMZUv
uO2cr3DN5DPdrOdK/vYrsfC7Lr9DOZWi1XNMxGxJwwpwCkN6IRvCcSTUByaE1eqV
YYOy4Nmo/oFn3Yd5/60W4AlmmTeqk3sAXdF9wXagcQDc8KA5ajwapQV14gEQPx7a
D3dF4DOXhjKt7/wHy+Y76qPTYurBW5zkhNcwmoHgDiNbf9hB3QkHT0fzuXzldNqx
i+I0le2vsc+OJmf4yHvt9HQnSur+fF82Z6UfdI5Q4QNBPUWac2+FNnXbnT43ebdv
uEqDH8shtjSdnP1h98H1k2+3Rwaunek/dPrITWHGdSBx8qk6JKZ6mJvc2IKYf+tA
3OnKx+tBaiAifzqX8Z1mRrDLlXx6HFx8qnkFdori/8gRLmguDEFqw5T9esvjjP43
VfA5ibseVtLCF2hL9Rg9KnRzpWxcu8oFaLlqX//O91hnNt4lRoqpih3QLicGuPkF
pnu9cJOtFlmEdxHPm2tLDQxymfzajce95AwPysB39Hwn7RDQXnCBCuYKErZcV9Qy
zo5yFCwH95kv54bMvdvW6JmVlC+3hqPxiDAMi9eZWTCZr2c283DvZilruXu1bR69
O8psOSZXgd3wY5XwY5+M+G00whyZOXuWvj7WwlIw9y1dhrsuMyYxm4q+g8u/CN/6
Qc6HOhHpqhWI9kJOm/0ff1XAy6/sSaQTsLgbDzirsV/qumDI9hIC273K9VnjmWSv
PRlz9yKG1bDOK05nych+CURNbgPyFfimXgGKiNA99qQk9ZVRvgp47x4VDDaS4DOn
flyUCiw6i2VJu5+urCY+0Bq9DvZIuNPVIkTJIZl5mNIXR9HwIMj3egtMc3sWHvb8
ApTtnWFklJNflSLtHr/PgUV852WU6/SU31132Q5sY8L9s3ga1m/tMSUNbqpFrP0u
2RJS9FeB6tbFIMkI9FhQjm+annCA04SiPmFove90prfrsAU0/vGtBUqlLEcYqVuS
IrnG00V831QzW7WOfh7Uv5ScvI/4Jpe3jSeHtzrTp/spAt1NFpb49152f1OQgbN3
uZrByyx2lGGeLT9aNbqZzPY8E+GN+/YpuZunJlrUDvWvTOxyGDEJIZYCfwgNZ5Yo
srz5IdiPYiZaCUaqIGAUdOu76MYpMEyNuv8S1yAB4wB2ml6gThK9PPJqfIpQv31i
y3t0UYzoOoT2MW5Np2pIriSVZc264LgUH/QqSKU3Q1Cx98MVPTwQ/qOoOiwXlg54
odw0J0fvs3Tqx7KpI5TDXpTmBdB8OjU7h1mAJuFODO4BqCw9wSLfBnqAbEl946LT
ylfq0TaXOSL1H35vLUL/f/zTS1hHzWkrFrftcGSyl6cP0/JmdqlX6sD4YG8Rhry+
+lGc7xKnJgOka9IBxxlN5yh3batntMcxDK9A+gkVkz0e4XkLew5OeH7DX5kLS+Ke
Zs50p3xqsmbzkLkYQWXhm8hSHGnkGqnj9Fw7aiw+TYfAQtKU49cXw1cXwHlWlNk2
VqFRGF858yuEvto46tJa/U0BxuXJFn8gE3128UAK2Phrqba/a+0PmU21hQ0QbclB
QVihsCb+jz+mwoTa7bqhc0lJW6WyCRdtttH/HxDrgtFnj70TCrtNSJncq6PEU9e+
xmEkja4GUbspbG2lMMppJ6wlbiX2R7N6gN8YmhAjEgjgWm6S48KBWVMoSCECef8i
F/wADydVyVJz5pwd272f7TXbrPkA6liXrD4CnWGtxu5rzGVo9is5BG/zoaDc68GP
vhWq6bPfAJiW4TSMP0bVbEqLhku+q13HScbd7z41ndsTB6ggqd+HhQdV73RqefIc
nq47f+g8VhD+Gk42NNjOf0YzSRqHB1EubJFHG7wC+/t7RiF373SREhhoq/z+pEF/
7+l/zYFIiLxUl1h80W6O+8iIB3VIsim3hJrepOjiLCkUF4jyBxiNJp7hotoxqfTy
FiJVXB0eeKEMJo2Dyg8wH4klVMHsLO5L5B2wF4gW9MRbwwDTy/9UrwUKh7UDCUoW
GoDkITqp5hzsEPH+wH2nWcMxCRjj9hNI7QI1AJCJ3+Y+QY9YGKDF4z5wKQhEim3X
ShuC7Yq7u6UemLa0OV52ldYlrmVSivP+zcLBEcBRtQbLMPRhbW22+z7qJPn9hm1/
KEj+75QbK/G4jWBL0t41LG5FlyljTYfwOvEVk9ZGCd8hpjXsRlRBiap4gVIWArDa
To298GuFOblrB5w9SsneXE48IhH/GiT5aaqLzwGwEd+mn/JvaB9gNdMz7/Rx2i3I
ZXbH1fa/Af8+nnzrMWn65E9uMVmZOslZFTPWcWAPK4ITh6zyvvvcTJ1ai/4iYJ+B
lj4uK/Z7vGCWFk9v585aE9N5l1LLjw2VupKG9u3UMFJrsQG336t5Law3+BIeByXt
853ljm0P3eLtyGxzuIDr8YrTsQ26+M7S6uCIWhrgJ2kJLOlRd5hnFLi9UVW2OOM/
mcuPz1ZeR6jJn9uJknJkkNgAjhpst3xKGLLakgdkihVoHkiyZ6y3pP8WUWsbtCRn
lGTXISutrQQPXjJT7EzK7bivIp2UNXMsIqiTTcRikvU7hOhVx3D9IEZUqI2+hdpH
m93dQe0WJE2r6ag8KE1ArRuPAmOk6A63D24ozm+aCQI65duFNQUJFXkI5dqZEpjQ
PNG9nSdLc9gmH5ozs+YHVv7ELFPL3w7OIXiwM733oDu9AklO4cLbjpj420HCGDf8
gSJdZD8HX5H2GLZgQoKJiEpf020nAN51vQnuS6eEWleWqnOy3CM2nssaU1t2k/7C
Cc08TV7h7VK/YT7LqoplIpGXpH9VaaoJ/IjZJHlsAXLNQfsfKT4kWBRHxE9WYC/h
adDXLrGyZgkJ1bYrndYNN2vuUMhYjw6/RxXNezKmOVEWumTAJmIOasvA/n17INby
LHmOeW39x7o5Un33s5bQsiY3sYSe0oUaBASscesOJ+aSVk6UToGRvpG7v6siP3R2
tj5M11UH5bvtzftcYxDPyGkm+bDH7MD79aIJmflN2A5AjwXaV8li5MWr7Wj1NKSY
MfedSPWWHMMd0G6w/ycjJFfR2ahsQHt5h8LFHZeR+PV2cv+pndFUGgeDK7ycFGHQ
zIl37UfwqghWeI1ztMmHhAoV90xGXeWwyQHXmYnmA35UzELXJcr6vxKHGxfS+UUJ
TO+kmd6JBkUg/+Z5X0KUjcKmO3t8ud6h+H4mW0kSrGwuoWMjh100qimC2QixcN0g
fkffBAAATFsyYdpILyG2c2V785isbvayeQGZU/sGfMuPm3qOrj40eA+/mgHtTTzM
vJXCSGkTKFZ0xn2XSX3TvctzxA1Gl7UhUI2wVjtZtVjvyGcrstg7ccg7P45+tRgf
FQTG6Va+s+RyV1qcnGSX9F1N8kNLnYPKtLMqwCT/CFTwdTD2dMOSXHGopAgc1x61
IYXclxKmdTtZDEoTFP1PSJBaZVJtJgyRQSyO7oE8FkIGqLVyukHMXfdEJjWeH1aY
DiIrAyu9rFs+d2wq/sgCuouFbWt4ClhmowFadTv2r7BMlUpNxxX0iHp+cNpIFSZY
WsJUDHzIryEYr4VdEK48l1wDIIgu5iZBteN5ZnM69HoAstfaZkSBCbFZdvAmJFEL
Ychg1mmC9oTZIM/DNiR38pndSCDaY8zXi/c/RUQonNP+2hMNJyyyyx58oBvIJeS4
NtW4aPgHaDQLFKkxw0/g6ramSe3rDPAk/Hnn/mzybeXo+SwExuJ5YMPiNHn/eyW3
fVydIeWvFSzq4JqwiwiFX1qo6D0uvHWZ/lcmj1vHrjypXioMrDqW5RArduwyWFkr
vxd+nAvW/Vw/QNlGHWYLYNs5JBpAxItBh8ArCaCfmy3oUe3yH6tFAnrpSpPH40Kt
CoeAfLFbIcqTFhnCEHPVcJoL2hvrxuIABbYWF+rcMkCqEbbYjJKVUSKTvKzva5uv
uNBTiKEaOd2NlCfRcNjSyyAb2uXggZh7xTgTBellF0TLYDirBwF9DRruHNo3EyRc
l1NtuQELSNR3E3bXF/ivThRSDmv8vo1/gKB3NY7s9nqbBcHyVhdZ6UXBpRxOfCUb
AzjJDmugM8d5lhnun0nHiOeP9cFA0Jz1suLSbYTwMng78HHQkLnW+4TGd7mZMc6q
PPxPrYrcDRig+7XQ7m76HkflEN1ZJE7TpVx35Qg9wBzH1QsClN1W90l4qo/sYcBX
zhd7LiUfxCD0DHATp/M5iYdcIa6W1mKSNdIOqzKKxCc+quUxytAGeycWBNxMFzlW
oCQK0AmPryjTDugf/tMvcIwIK5Excs2dIUDzXGulg8uX4dvoom1bB6PcUgV5MKwZ
GIY10tSq6Oti3b266QAZSILimnYDqfDRApmGhBfVv6OAiGFQ1RUb+KnFhm5FkdmN
hl71cfVEq64jSWQLDo1jOaZoHnPMlCg4G57Sll/wx24DgGEbTKRS/Yddmlcr8Ari
1uXmxyJTGTZOh17K3a6k94lMSnOHQm9MrY2F3cp7ZmPQBW2UksyPuzs1osO5nwJz
AHl7Ouxx/tLcJyAGZ9Ne1MK+ycguFFy6ZpeKt6tBMJtVCHUkJlwW+i1Gx6+83aze
vpn+S7UFgB8puQ6DQMZaHhjR3XBLxOZ/QPzKLwwFb/JQgEYRUhGYhIYgo95wH7p0
cN3mRua0wxY6uvifpL0ZRBcUQm9HomEE5CpInujpWVSuWmbz3p0HWF2QAysv4C81
Usfz8IddX194eOVQ9mDHlEMVbQBiMfu7LYmVgepgpLyp9YKFFC94qGCHo9lkOz3p
dAQUKT674qi01W5Mr6Yk1f5QZRQJx7u2DQKB25mzuqdJvwSFS3kNOegjc0DB6Ms3
o8+LQDjAtiu/vg1zeGB4+SOrBdaDR2VnJVcqc99i+2cZKhWX5R0Iq8VlgdwTHKj5
7UWzk0Rac/uEA1m99uelXKZh/FwF3BDNNmE49xuhA+0Qd5rI1v9kORrP8nxa/VWh
oLZhh+7ta/G50HRr2TBPgmiKmTweerSvkS2dlallScj+JlugSTjoMMBxVeAAG6uX
SqQhpTysxfBnOOsfJBFF55n++GH6De+izCJukduZfwxBmtsoEw3SuvAgrL9mwlrh
0d5qKgHOWfk8nB/TYZCBLB2XqvEK4jw5UzO+QnNIvbYOvohFI0utYNOgdGvPhubs
IuW21unWainOSR88Zj1hA14ZHJQMViAsDB/qVwBfDoQW8jo1gXExPFFaBYgNKBk6
y3fxcoUjbMTIWPWQjGAdqtkT5OqtUVfBWlwIk98AiIbAQRWB7UVnCuXVWTeA309U
+mmMQkYidXofKBE8D/5PZvSutHOxluCsryMWyXl407JFex823QjEufGMzjA1Wj3G
C0l+d9GcHfMbDtpOZT7LPmJhH99PZqGO/vSWFOuKNWbGIaTruE7RUcXGZeEEGppD
iAWdoak5f1HXxEYIUCaBNDvPpGdgOKAv3dl9vV8zv0IiXGwHcKJbB3H/8tH63+dU
Cs+H21aIYX8CGMN0AS5Q+bciJDiP/xSat28on/tm/ffbo9u8E55pEQjlDWn26eJT
NatYLJ1xBT7NBmln9e283ih7LP8r52xv3hBBe+5sZFEiNvUj1pgi3xTKh4fKPNoV
u5anqKzWBDE57ELDFSMjtdkxZsRMDocpIlFkzW64PFLXkFpys9XR5HyjeNRAW2Rm
NFgoMWmgXgROy9Kevu/ueWii/eV6Q22LpI7sY1LC5PLw9mrMLLLKzNQK4GUv4MDi
yT5gTy1uONdfNsRp6UJGiiNGlmxQJNNjarFSNLBzocU7xnpyIB/IfqHL1sKp4aYG
TMZDRnSlyzTEUqIFftk/pgxrOgTZZ6uk6O7DMY1Ur2H4w7BBw9fn/UDBNpD5a71J
CuYueBzpOayWfXJxssEQW1oRK3970hmRLukBlqpxyKgQbKS8b2UeM3xiBU2OGZLt
kHUYRmOxEizxjGyVXZg3GV0BjPQT1+A23V4IdLBXYcZ3slb97mOVsIZOoefMNJDA
RTQ0UAHaz1RhsGwtDYkZgXrIH79vQ9Nx0UBJdvU/84h+/d6tLCxoOrrPFcBdkxc+
uM8gKp4gOumDQdXdKmcPKD1kieYxnVq1SzUu1Dg+bgRbCKfGdjcTy9PtBSELnrPC
iNItXJLkk2wadYVsDBBb+n8p11PKoFXEl72CFjGLDEEqGnEprEEEYBjZCuDYK0QL
3f3WHbaRv0cydr9+XDDoBrsO5Q2nHGD+48E33L3v6qNjJZ8L1Y+uvZLtaMN9lf/L
EyO41JVbWp44Mn/oVsXG+SCm1x+naWcDeZXIA+kSony/soVZ2nTy/Tnc9t+KIQu9
BSIASFxu14B8aNOzj2NYsr+xIb8Eqdgh6wfIHyzmeA4UUggOKVi6p7mBkPmWMBLE
1sAohElZwRgO7V2JuGg1K9uzSKe6unCq7ZM2B4n9OPEJcFzLLfoddm9iQXC0LmDg
TZGrf/0Ahh2QFDw/d7/5nAvxm9Nqn3GOHkWE+hxnpRgWJgQ72aQe+1U23o1tAmih
7nQXIIYTS5lbvTzngdvlBOdHlUzVvBG3MdZbw+qHMbTuNHg172H+pd/VfXa+RpAF
DHN4tPeM7MbkdDEGTabUbCSon1paTPxncO+lQOufFnExW+qr11Jb3or59bxjlsOd
4ufU3EE2i2ym2Fu6j1I1sU7tDGhtpv0/24/vCfAiwSsFQT5Zzenn7lxQ7b2uz11W
11MS5IMtlYOCWuTTUb1VHhjKl3ii8BvmP+/wRY5Cyu2zOgYfEkZWLezDikh9ssML
6S+t4M8Av2sCPAqGwmNAzmQYWg27z/HKTNLXjSzCAdIOsGVOSnsL16eW+HlJffyg
OBpo/4GgPTWZBIMLoreB+nphvQqq/HERg+IF8uNmRq+HgWLKbwub0Xu2r+MeFKCH
IlHnvTQLa6NpksauopuKgLkIwzh5n5GLjg0WgZtprHKw9yKbGp9fek0nf3dQ5ej9
Zbvi0yp61ROsyMiMA+YB7ut/1I0gGjGCMeATTePs7F090g02C1Lf5jDtydA+cayV
ZR3ciqmdP/lNbrrXAHzXe3cJ16voMrCcWsSkUSnD6i+51g+WIA2mQ5Vyjr96nrqj
2kh9eXyYoEhBqsH5SGN7akC7chIRTajDzmDw1i0e151VfwRVA+oPgf58OGak28oS
3qkUp8Dm4SFivjcVnmMO9CWdMkhlArl/222FviW/z9oc83Xl8/iDlCC4s8Y1EpkH
1Ja/4XH+x/Ye2SfmYexk34UiIQ/Tux3txOsaOmujLKmaT+vQPgSRDIpyUZ2ouuyy
9slnzRniicdgPUTRAKZ1PQ+wlahQ7t35858GG328TGzNoN5e2rf9xL82c0DTZCNt
IzpwpGvC/TC0NGcZC20V+BdqssvThTYAatg8m1vWQvblNgnETY3NZZ/f3DuuHX3F
qG+Lm8UJWJ9RWcZE01ubzWclqskigqnzPhjr3O46ufzMtR8I7klgLVoRtsb2jNL6
zTryOG0CtW6Lop+R4odUfDPLaCqYdGcmzEzH282DtKEjdrFZxo8tDNI2qB93Fm/k
+VqJeNoav/UMlXmR4QsRyLBXVeF36kNlKv4rBOpkGZznULL8t0VWI1CHaayxwEsI
8DJN9u7/ZiQYLyHuM7MSATl71U3QCC1j2PKBcgHkdVjWx2nMt6CBhJWDHAux2aOY
Fy+UfZj0LX4TD/YA8xtAMFw27LfoVvV4PjmOgzZODDVNQPmTY3ph+HD82cirzkj4
UN9mjCA4QjEecH9pEOE6DhmR4YXj0Sw81/K6axGtoaPXXDsjWSMCCKAth+Jg7gha
QnscxIXQV+Mo1xXBCADUXO6JXQ+L/lyB+cpepSCFtaOmeiKd3ZzTKyfFQlbFH7UR
IwnPBkTjO/NiN6VoGcqpUS4Vb5JxpuJy8KimaK57+DAVd1IPf+o/LtaqxBGZ6spd
A9BLqs0IW438l4g0OJN27ldoDsW9GEs8iQX6Lw28FcuJpaQEJYbLxopEYVSTl6dq
lMup5UUKBIHJ0q46JJgvXfKJkP1sUYvsY8XDLfRId4J+SgiqC/PrDY7VMETBx9SM
+6iAJSYqH0s6BLKnFRPboWiIMmiSHWv6t8gl5dydI9gcbogwQi7bBDqO9l/WFQQT
TtLWR+jsihztlep0v/fTgILWgN4ovVdRMjcEWpwUQsk2wFL0mcY00BPP8JcRVOeS
PGqxIPaT7vLr0/hNxiCtgdWRSEnWV/DqevUN9P9DapunaXcfSKXT0r49BplUSGzg
9fdKq5C7P88TWOPnogBi1thaEUJl29C34000rMIboes7bjk6m/mHcZS2UdlMvbUD
RXyFY1GsoKlRViKUPgnZhfu9qb+M7Gt97W7/+ZiLLTwvgpKop5JG8agn+nLSR3vv
dMN1Jug/LiGMtRFxXAM8Ph11RD0kbTBgwaK6foi5kVsOJZyNULsNJtWpS3c3BDI2
VVVREir5fM4vm61ruXHUOq6uAFpXQoBRM3VxbQCIoET2zA4ogDpT7ndcsdG44n4v
z7l6GuPhO2qG0GXvJQWW8hjOYwJnA1v0KPRhQNIYXNccUt/JVpncYTYq8A+GVM/d
nT9aPiby1XH0UZxCGvbE/wLLC35+DOHs8uDNvBgH/YvAJT2OE5QmhPs2j/dMDFZ/
LmC2K8NFNhHJZXewnII/SH/nQV/BJYBKQ+t3EYft5JnaCxSvcy8kpdE5dxjwk0GH
YFgez4s81/GLYJ9q8r7Zzq17IsygbhOes4vgLRxqG9I8l40ZtEDXutieV95IKYP9
44NnEQApp4OeWsBR0Q408sdllxSLq9eoQ23zrcB8P7f6KVh+lYC0LIxCEvlh5xgv
KGnzR9bEa+CYQSoDqEfY2YhPke3CjcfWfepnRZO/UmCFAnYSsExEKGSXxlzFVRRd
RWGL3+p1xWFvHrV+bnZHY7NOcLNBUCvk8H+Z1AA2E1bzJY+QHi322OkI3uBV+IJT
VT8UJQ+K1vy16VsGz9HYcDMxdYdMhsVm1x/eArktjn1o5tely6vbi2SvKyo6JWpD
o60hmiPu1Xw9oLw8sDKo06h+Gz7Z7KwXZrAgv95Q8r8xD1MmiHSFzKv0SUkU1pWS
H5lHCpBd6JfDVHsqniMmOwy97uuu608ODMmW1z4vGt8jreShzjFc35pA1+TZ0VCn
EYniySBeogt/YuY/8JKXlpAe72ZTLpI/1KrkNThzc73ZBhNWTm2yOK2/SPFjIiDt
Af2jCJr8KXJVOlxgNse4W+vZ6IfJ50EMtQF9O7Z7iyS68uNyIYKJrZccipApwsuS
abv9W2Cbpv9Y1nNf1PSI4eh2a6Dp1qPF+AX4kbujc/xXAUFBhW2J3Hw7DvTRtwat
TaHxXI+/WmPspD1gzcP+pjl+g+o9F/sk+9rQnJns9mqLKpSd/m3cuhuFLKrJEK5q
ubzDwFECy4YJCFtmh618S9nKrAy8ib1hr/CYfj6A4JNC9LjR0yWMBFAoXJRb8lDN
IYRBwbK+rnEjmxBtDZTodeQzLU0ipoBFdvTbIDj+JNoefBS+aSbfPvb6sH0OzyhN
EPRViRzv12j2TCCM6rbomKvRVuqevjI8HIpGbuz4C1obSsSaqAkalWin2SP19f49
8dtPS4DMXeWbHB0JOZEGs9XQLFMHZ+VYtOJRF63mLI2kMAW4LhF3OUly5DGdQj7V
rLSaXJQqZTWoNPlwD9AaUSmgwximg8n2zJyk+G6z45ltDoq/tmgwZqbv3expwgKM
fOE33dUzPaDI3K6OBt8QhXBGSMc8GL9P/AyuXxVNb3QH97qBjCJUmrrW5FyPjOKz
zbzGI66bO/6yPyUsDyCCOcIneoQ1V8uYwBYdVEbh5DsTm2wAt5mAXsseLih4SnCf
TtlNCWqThH+j4Aaxt5CbQkDYgtucMupo8SW+GS34xWEkDNL4uqGoNP4vACHuMLua
5c725/y5NZppyb+/wRejV4U3Ts2FqX/1Tm+i6JsPvSLiRtGkJrIgmuirVMihdruL
Zi+yxWA+ROi+DusMrX6g4PV5fFW2L+l62aq4UrrG4i7aJk9g7FRTtkC8y65mF/l8
WntCSaXxzSF9O1HiTnu6vWB1NPXmOJpb7qDDPi2wm9L5Rm4vW/EkdHAT14nqE0II
8CjWXAg9IGI8rPlO11FSPgGhvikflxudN6ADjWs5mdc5+KBkrUESY/3B81X7sYPw
yEIBv9IaW+MEnEHxAs2pwDlZkWnlNlVtWjNr1s2F8oyRc9Huy4Qb03veXNuQF8n6
T3PqCKdcACgRzPvqlfFHkWco0eX3841J+km0nB2PUI0mXH87Zbp8qILCimNHUxBz
SfVv+bPyTY5Xtj2/1Lem5Xv6Myd63LVMSGdloVflsXtTytJItXg6O0EiY2nrYsNs
dl8qdhcV2SjswsyctJiMjO4pwjUcy+e3tz5xibiF9pJGx1mNvcAcfzHItRo3Ww1g
Qvv++A/JtrpioAYMMvCtyoQia4KGL/qmHcpyvb/thJH6XlOSPJt4wwolmwhVbOQV
7IhWHFUW06bJWxemvSCOlJ7V006qIRautuBpAIEftxG+ZWK5B5fP06Z/SA5+Dx5P
FV5kWtTWQBMIK/oDqbieBFlSYgtCSsjJC+Aw3CNTv5aiPmQWLEZIap6zNQmbn686
t8WDvglhqUVkDuyiMYgdqeKv7QEXgDY47aH9dz2kucJxeaRv/QSMWCqOR5ovWaF7
uGJPrOzRrVGyURTZXfZWOL9+01WE5cr+keTSKk23l0dBIDllZ9HENUMfAgQoHBhV
TkRUPeu00W2C0XE1UOSvBFzDV6+m7uKB/5lHalZSuCPeZ+kDOrbxXJX3QE5+ghZ1
BZNl/evFER7fNgr1qKH0LpxF2uDnmeIBi9EsENn+F3f+g2EBzYhocqiKfr49CPJX
oFx7qLNEo3Zrh4n6OO4sim/pMKZ/TG5CKzc/hR6AxpkEj8rtyqIHJZJk5+vC2eqb
Sf2bWtuto5i39QjSbHI9dxotf6H3+yrAy+xN/sHpBW7Sm7w8ev2xC+WhwBpPIhta
KLu69YLHiuMvvI4U1hZ8s2JaNgpR/DEyLZYwhf2XK2mgT0nOQs3aJaZMafFJhJMa
n7UAB//9i3OIO4eYNNjEIZPMgRfXSu7gHwj7z6j2GVRvS1/dtREPJLSUNz9wW64w
xo8y9VPiVse6c7NDVUxAOqo3fyt1zm+cQbf6LK/Yy3PXg6xUFkjs2h2xIcGjmDgx
gRcz22MiOv6Jx/yiJUeUAxgTeuZWh4q/okGJDvR9HKn8YxutQFDouvU0hhWdvBPu
e0PtHQWKmxTDnFYuYZib8hfcV53Hlp18ZSk+jLr6rKuWNksIGxPt//qEXYV1ErOj
1xnB/Z2cpk73D6JF3IvlRwy/pAXEqYJE9x1pltLOU+8wMN+m1FVfp9wgr8Q2sIlI
8s0lQlTbTLfcyrLhXbvg/PA0zXkmdl+o6Bp7NU7Eac8sgsNyTLMimEIePFxlPtm9
rzQ3soZgbzWNpYEPGtU7Yx9Yc+l6l2jZ7sGw/WkC0vAMM6xZzXBSsuJi7PXu6BgX
ZKBEN61Rm9EHs+lIvxhxPVK2Yq+/YDVLtpskEE5neicNFFRK4orxARGn0WvczOl1
5Q+ssoJHjhjQlSZjEYM9s1sCIbvaxBtPIUxuE4Wnfn97mWcuEkkIagn3btwxSB09
ZNef4QOHTjkvJmQH1qt3ScIMBzOKZmal7ehuDxZVX7CFc6fX3/1pf1xi9/pDL6Ti
flVVvPpWkxKDAGLMcrNSSHcO9EjRfZy/SxuwpOvsIcZYE5Lx0000Yw8u+2LOLNeO
+YrN5W6FLH12QH28+QX/dBh7ZSqg8Zzfl+nuoo/5LSScaCWF/NDiV+r6V+zVyjhb
xQC0C9HsJFadPF6BSha8Wr6jTqma+pgxm965u0CTAp1Mj6j/UUbXx5ReuaS9eonB
4KN85vZGxtRORZAqpX+zVl3otWDPcgm5ErO/EZNj8LTU0aEx6IV/O/NTEtoiwjnT
ZK2xMstXUOSNeiROCqPCp5PVSTghb9zexl/9G/YU/tZ2eIOKbYYXefjjLjHyl4JE
B51k4jpKc0r9GnT583JwL0M/RIevmoQHgvhyHv2vhdQ+ScoxBdVRobrGWrisgn68
q1l6vwqZDGD6NtBrWsSSgKnVT7PhD+vMHXiWBRSZLyOIFQQUf45cS1QUZ1WgdLXQ
MbeP7TrshWXWuq0VL9Q0latSCzid1ab3weEreEClLH71AtqSTOEw5NDPClNXLjRX
Z5ndQ04JBRZRAT83ftlS4s9+g3Be0e0CBuzfbzQ+U3lidz9gJM/E2Vo33MYlduQL
x12nZ8XJnCJEBInyjcEXd92ArU/vCnJLuyZBCFkueB6QgFVZOHEzAHuH+FsegGUA
KIZ71Z3DTilz/2j2CmejLbBqYgpSVRs4c8SOsyU1AW+5Bsi/3/hjpiIe5bKrRoPf
yFX+u+XsH0bGqXHttbkjrE0O+Gj6qfIuiv2SKA3qYt7S1iEcIi6s4a8T22RiVUGZ
cyMALNQ5OMQkkxccJtLTFiNBuyaTFZ8wFgew+/obeaQKqTskcF/VKDhBEpVvhWej
8eRhUy9wMPrcyWQCQExJGNzTvADGQuP7fXzGcgpKtuMnImPefi+sBZ+rr01PlDiW
fVrTZB5KEB60TSIpfaAQUlqQ8WAENPMoebTwEpmXEMidVAx9S+XwFNyF4PyTZzBh
6hN/eWUinUTHcL7F59YI3m+8DePNPHoCMmH6qVWZWLWkJW/2F1fT2MYpRk16xA53
zLz3/zVS+Jh9Ae3anFZpN5EI5r9MuP61E/iZSgYat+8/yIbSMmO0x4UgCaC/wL2K
4LNWLUjgUxO69udKL7J9nCqsfYm1EKK8DpaOq8Jf/DhjJNn8DM9n0DtqIqGaN8MM
6n+hYaN8mOiqPxqC/jV9f8nDSmKKEQOl05Pzppl0MKWM78FQmb31aZPIPkanTrqF
zHZyBcBuu5CBiBjkaG5hbdE6fBYnikeaeXekK8ro9wx5qmLlwIx1FRfJ/OssSVKB
BWIpngE/kwp1C6WhdXeNVF3TdVsKoAa9/bXyUWxx35ygYk9rm9/Vx+ym75btUWsT
taFIbUpx+owP/mnn2nMVhahumbPs7TZykopS2hc4YiCCzbHGCcKa7sKRyfhPwVvQ
T9G9Tih3pvK0hYw2ADXZtXRZUjou4AYpDIzb6wGQ6pGyVnM0AASRJ0TAyxdG+xKR
9CL20BVirQBQQLqwG8krOocG/JA8SWecthbIQr8Q6mMlxt5zMk9FDyc/7VIJRXes
Z41dJA2/AdyRhSdPbe8XXTH+4D3cFQNcNxOerUtC0lqCXEvtLDjg3iY1cr/KFOQs
QB6mIJyLIqiJqIUZwnE+LliUIoTyI53BRml+p+wRW4VCmsNal4aj6H3KGZw7xTYo
Rvj2Hrw1Pu+5C/lk5PFHAqmp790QV1aldLpIbHgpBGGCh13ijq2UPsi/ZDS4vFsA
35lVMjCEUsB9sKLOwsx/efdr29Rs5JR2mA236mNbQznY6nWnq+ppt0K3JGMaHNxE
xoWAnxgfgLnqi7koyOUu762f5Hve4FLGMLvMqK0e+uTzA7+HF5e/W0gRgo6A/qFm
eCm0cDNfn7o+ySzNQ/gsMt2hFDSFE3Kq62x+UCUD39XxZWgfxIL/r57Ko/rJhCTB
t4Hd5hDp2aDuOb0JqeIGagR6j8zh7g+8Q0GzmTR+YCQNRUYczqOFmBZxhp9xFbXM
HXh/yCEJfUoz7C6FLsCPj6EHAryLnWfAe4gp3gfpT+BATfNqN5KNn9lmkmx+cm0D
h92gOG4PRQE6Sv5/oADpW6h/B+tCpfF/gjUOJ3yyJFhHCRUVtFP0Zc4NAkTkxkK+
FSBS31iblGsQ6acKR7rG1DRKEgA+cvDDjqNiIhpPG9eKIzHUic3dNC9ZolGbI9l1
Vt25rnaIELB6vcxBBYkSd7eDr0Up9k9WjRpJ6gtyi6nMxCnxkjmVM0hjiTeKf4bH
iatunBL9SoQZeTRh89ExKzsaUsZgnxMshpLJc90H5wHn9O9y6s5ca8cULh8j2IEa
omIGvMXDyiCJxxq1o6bBZqG8NXkOW+J7dyRC9+6KcmCEUbMufgoRJOd1WVWXvFFy
9NvclOaAjMtAzACflaV0q3Xikl6/qy2k89utIDAJNOVuDP0wkDxzmeuHYy1RTibb
/X7wPRKCURvRn6yUJvUk6HH+oIwWdwy+AAH0lqaj9/Y31gz0EcKJC8Ha+BRf57ew
j0+oSGa+Cg5J948RW4+5IP+6SThowQBVUHEnCTMfbKXTmd3kNRHpCNU6J294RQm3
8ymYmtXmiNT+C9ziRqebyqT50Ylfib2P/rtFXEf8Yd/8x2pC15C4kk61EHfCgDBc
VSBnFjrl6/w5vIi9iSVMGZZGFDJou+Hzt+Cfr1osJkIG5ymmLyTxcvYt+9scOx+y
g25oSipYYhelkZ7ojPU0xv/8VaCbAzYrDbWjO53mke9xLUabqw6WxbbSHYYPKjzq
W0dEbAN80U0lpcaTaKmRmxWyeCWJgpp+dc+fU+C8LwFJGbLaT3bXQChCCTFLWeoi
PVGOr2V7xyty2AfFryx+BBDi7c0FU129ebn5KH90MOnJrxVWnyCuJBVe+vB5gDEW
xy2v1SgDSjKhzZZYBSBXsSn3VFW4FAYjVS7n4/7/dZgitF5iapWIIR7jiXskjJMr
2BTWrHUZtMPlUCN1dqbENS3Q9cKOK6Zf2PLv/0bHq1shlvwbMbkfI3SZqoT1Psh3
YWo4AV7wBbJwDhPmd2bVqDi6XF/IkVhF//DtV6j7QcgggOHsA9d9rdx+DT1lRXwI
mFsBcZNiEKU2UEHN+tb34U6ksx2PNQvaQiMBFeqsMcK48ISmGoGoQIMG5PZeLtRO
BvUMTBmmYmSvkizxLVI5QVnmCztLMiJYmYsTbboJ9SZRe36Xvx8Im/vmTrDxpZXa
hmE/8zWS8UpDgbakQe2OgJBsXiQOX6HfZ7kH/jB1nuVcRK9g0puVCCf2NZ0tsesn
If3aTUkgyYLWOtwnCvTBzLL4E9SO4QCQ3YiuI9v57yyi2IIKbaI3XhbO+9VxSJhh
OdWCcigJCwy6uLj9MsxiQ50+n/RAdbroXCqwkNZEdMRpW62cwma2e68/kyuGnDXy
uqqYCxO/Qztyqv32wHBRxwP+TGNu0jaMiBvS/cCbURXFV63wJCPo7nlsnI9blXCm
0zAL6PvASfCM8/fkXFdS0+ilnoWlNM+Mf+M94WEyndDlDtOcB1jfF8uGOhjtPaV1
/FFca5XliaUl54FkXtgm/2yQ3oeUhw//RoCj1eGXwj0zO/mmc5x8jP6PnD+q4L+U
JdDrAcPYBAlrYO2UTLWsQb5a+UEVpOz09az2JqPKHlFt4yLtm5HpD5cO2G4sqp8/
z+BocdlplZzX6dKfVASkHlXbh3i7vLnzjKz2mhopCT4qRpPlhy0z0vOwWgADgb88
o1iOYkeLqOB+hk49RxRaLv+yJly98aZJxuPObV3tf/QwXtsVlhe8Gp2FEs5XSfqf
YJuJSDDR/lkSOM+zBqFggKoGxbP4mAwlPQlAkm87aNEGNkPOsTnYD63bQFLeNc7b
44OKU4kuAQAFQevpF1jB+xefi2ljsN0sbql9O+jGlTFGi1tAJ/z3Q6eOVPZI0pFT
Gt0KXvjtfS8LsAr9oowyREq/vm1slfofMeVv2a2HqCKiOJP6FqAQ+PiME0lEBkGa
DnEsvi1gz6e7Ytc2CJp3jjU8pmhnA5DMzGBp/NJ8dXKWcuKj+nGMJwltxv30eXNe
b0ibfveBlztw7QqEgaPxBpykqBMtoqzjo3TXnQ9u/RWe3SRCQIfyyRKLQ+Ne7MW2
aTzPd7Jd9LjvCPYpjuQn21kZdyp3FVUu0DFGQaL4FVK/fz2k1QY9HK8U7HElGZi6
IaqhcS4p6B09dR+s/lVwpQkBa0cNd5duIvtUOf4W18KL5mm1aCWwGuTDUB+WWjsY
Xv/7CCjUcvgSEB1mY4pGdMy/vPXxzC1v2Cp4AYATXKKNJ6w05o0NdcrIBUjBR4We
wgXIQOHqlGY5GO8644wQeHIDmoJm4KB3H13rZ42IncUELGZjA2z7cVx0hqnTcmZ9
F2F7U9pQdbESuU/afg7808O/1I2/fCDeOdZwQCB+ydayHReeAyiz6Czdu7xyAVkN
xB95B+YA3aFtzEDP5rakazzGLn/zPJRfesZGjT/iFpymDoiK7Po2tBSHB7dtfuwD
loGKLf1xPaYpLM8BCs0MH3IAaN65Kw03BHSkuv5ff6Rc+rgA4KUkxUd2ab6z9f4d
Deawzuqfv+GPPlV6gKVR06meMeMt1nHQ3l9vaGcrvkK5BELi7W46sGKAlG1tfi85
ZEjBjk1MLFTcQ8qYdP1ALFNwwj5FfTAvJaqTtbrf5GQMeORbNqkDGssg3getV5X2
nip+hi2qqciID3zZRf5Z2qmvSTh17+5/E4qfzGxhjSFEp7n1TgDhUPizIzCud1KM
mcStajGSybNJUjRVoVReFH7ipOYLfFdjJNUuej5L43mRdjnA4dn92BRuADs3K7C6
3Y9tJjQfZafhwpJA6j6Mn7GvydTsyX1PnaRDFEqH5uBHIZejhr957Vo8Bb2yYRtj
1HFDOegY0zF/g99BuV/+nPbPfwR8KxL0aYvNC+AYHDMeRoeNLL5/bGYXKqUwOraR
Yb8LvI/JhfLj5YFTRGAs34YgI9KNdAD6X5quYYw8fQf77F8gAnQ/T5DgsQrj3zJx
TaRk3tor551xjTB9U0XknDwzksoGQ2wPJZQLmCFSPfwRqZFXSLZZACnlWG+0k8Xg
0EHkibutw7Oql9//5aLfqlRtCBIYBzIN+exgOA3YO2OPddpJfzufwOMgBnd59GST
FK7FoBwQ5J5AOY8MchlLUNRXdbKKSG35KvX2i1hLP/FAcvJMsCGWeTOgfKdEpXJ/
9Xv4EMamJVmISXtPmGZs8YW49Vu2NDXifudr/6q0qOiye2J1tQzvqXAcArqDkcvd
a1mLuvbuBLe5Iwjv9C4doXfyZF8ycm3yi+tbSZVcCAw9cU68pE2dWpH9pXJya5GJ
JK26tn5MnACV6U86Pz+WQK+4vZI5PLz4hm++a+CazpHmpY39HWHNuGmfPdQE6J3E
AsGkE9DzAF5uoCAZ6VnWAr1Pp73NBGnQ7C1xDUfyRtoe4ahl8ksf8ILU0rHX1o5p
noXKGSM0wIzgRmerQELJS2sEOaGgQHVZ6PDXe+5q5ExH61J2OJIWUkeFIeHGb9kI
HthrTvBQAZ8FUKEdWr+oSN6O1y3a5NA3/F9n/lBUYfo/HNBbhBMlMc7xfciad74N
tsngKcIfDKgBqQhsMzVadLzVy+OM9qxA2rl8lQv/87EL5CeF0697z0h+Up+QbsIV
QXFY8xCIdRQlS5ReIxZtd7EWnPGT7cgwB7RyNUyO/7tDe0CKaP6OHeYgdGOA7Qm3
R//4pqhTXXePHJKkviN3DQeU+YXvpv4Pzs0t1gdrrbfrSQbs1cOZDhY4+VzMjBOY
AdgCiuJn/6//CusI+ct6DIIhjNHa+V2CadJwRoO3VaYA8CARJuBlTmZyjkq6U3Qr
ZYykqMpFQ8grsSF942UadUx212UfQ2P7YtsWu91p2W5htwPjwsfkkcFZFUpmIVym
m5KcR3hfkGnORrv7HXBkON/AEb5KZzA/1NEI8If0R21g7q8tVeBp3/JUq4TGhGe1
BDwF09LueVDi8zazQQN1pWV8FbGtFGO70O9ARJeW4GhnJb+g7pVjX6tut/li3WjJ
05FNiknypVlZmq3KJnlzpVtMmDRQqTMdYg/n1m9d3WLAnfsktyQ5rn1NKiApN4DV
QMI3c8bb4BL57DeHwLXfue0LDLXYl10bDY6QY1Px4WZ87V0tJJgqmdXD0foNErml
QA+K60yqa23tdeWLH6l+/HRgweO2Q+E76N5mb8LGXEQ8AEEHPH4uz9b+qqplzsfe
+QYzZ0o6goFXNbWDKxtBnlG6QcAcIE6/nHdl9SXYp5p8uczE9rL0WxoFmlje4a/Y
ITgS3bXpvD54q+hZxzJO+IEdhTBzI59aXTeWQ+mp/NOsjjdnTj68qFrxTFVizVam
4fMuZYm19PAk687I9+AD6rJ8Z8hMTjQDBc1kSEounK1RU+wZyihO5O4Wwbj0k6Dg
Xoz8fR9oh4v6Lth8AHGaBbIMPIkWCnbErwQE5FRTpJ/VtLBLsea2VZJiCqQlS+sK
25MpV+s72eUvvaidy2HHBAc/sqaIvIpfchtpZBb2R15XSexnTknRGE1wYuMCGh3v
VczS3x2Z2Kri/0uJuXdG3DyRn1tEro+kO315c78mnDuYcAvuBrWtJIpYOoKwn03t
YMl9526ox7T9SdUtEEV1N756tv5GGitQAis+hq+oxiLfx9GcyH/cT/CAJ/NxiJD5
+iwqLFKXBl9O5/f1ixKoQjOAomEmkyqx1i0TgOciOwwwuYiL4FrVt8vk+6VQvktI
XFTlFvqQnwCsupbLUi7N1gM42ykE1zlkqYpXWspYzNGEONvVLCoZvpaj8BNQFejm
b6Av+8FgwjEnY/ZS76wsJeI1Hx8mynqpJp//evbK8z/vbQTd71cqCwM5yMfh2+IQ
1TmhOFSVMKs2za4HR60qq1+gmyuj5wdLtPAvGjOOanSDtiAL/MpqSAL7tVt5NGFq
xHXpo3ZDyofdZq60eGd4wSm15GCFfzspYIht1INawdsmN+DslZGtCjZndCLdREi4
ozTjUtVn9P+tsYl6fetVP8b7l9QM08O3H8X40Av1aC8AczG9kOOLEr8hSJCVFQlz
c3bpasvMw9AXQ6D77rNhQVVJWM6Hr1U2zPCCeCMbr8I2oazwGB0zdccyFtcNys8R
bOVE/EuMtCOJeNFlZijdnFl9L36DLq7eP2Ykvg7wWkU8Wgs4oecZZTSmOSuESXHt
iMDh7EDokkmb97Iz1VXq9O8zOtFnJFRwcthIMJ+Lf9hYZ0UXm5b19uj9c7oO5fPx
5YsLoYdURpjxFNN6Y5+lakUP/dPpsWVrvKRW1Dii93/XbDcGqlpFSSC2xa14Gxmd
ajcFW/2kHQ3Ca+xXwWEeaHVx5rpixbdLN5QJOQsq5sBS4+pPFeQ51H9F78BwHdlh
jDtYjo/AxbUZjKr0oam132wjUuPZWJnTh3IlhnthRgwRjMxaOkHaoFYwK3IQwWdU
AFjMV9EmiAQKVyW1DeLAYprQLQ4+StAp1AwbU91UI5yT/d8Kb/KMU3DBUuySigxg
MGlswLY6tXpVCDbC9WgdiBLCh+KoIw7M0Tdny1x8e18cKFhoM4tIl/a5SWnOyj3p
ouzA4dBWH6C1cyr9ngYcyP8sIDlnSreGzZ9oy5v92QZ/pvgY7DsCRTfecLvt5MVs
VfHvz0HyZpzbUNeeOc/YLWPxwfUP3OXcB/62hh6pX55aY4W0s76iauKnp8sdENY1
muL7+UKI19DNmkWa7ZfsT7VLCqZlYg3vC1DYMP3kEK1rbrsCORYCwMhVJFXgZ6lV
FyqYAFCTGHwwTc1+dpwi1Q/5yrRJ5ihqGzCRFafFF54/Lum5HmJrsFWG+3G3k3SH
8Jf+cvSa4Depv5igrcxZkCvgTG5lrcEXNOUY4I0/VsbWFUuS37h14koi5I/IBuxu
oLbXESOWtKVCKWHIHsuwRJ4U6sphUKSxBA6KVRGgWrcPCHp9RzhRr+1YgWcIdFZf
YkaoqjzufbgpSRWaiJtfEHF1g351z6Jlo0XWZnKQqjXZgsUYA6LKO41L37nb/J1L
VG11y6ZYgtJG1GTuvbiqk8m7zNf9OvFCDCB/9UXDhtQPOgF8N5vgq7nYSFl+f6wg
4rYb4XC5JnqLG0hWz76FuC4wn/wY6zpodtxBkrVeJnpQy1d3YOdnFksbPHmJ9L4i
kZE+P6q0wza52qqJpEyHvsTdUBzqOc/uCnETbRuP3lpeRJrOhj+DkWMxhdi30wa1
jOzIUm1HfI5sDkiyaG032WsPr5Pc+CENZyeSeIa3GixY2uWh7cDJ8ZuvnpJPEUEG
4CjDJTMRD+OiRW24rs5TL3oxEShSk1LJFqx54VwdXxcrOAXbsLwR/vtx11qlfoLG
f/NInYm3liWTQS0I4CEqAJzxV2UxGGXs8QNldBPoxqCb1+bLQRMjdOcunS92HGxm
DvbCZ6vPdpGnU9Ve+CKffoVjrzEVYMpbtGW+0Gqk8OmQlK+PtsWPW+ma0dfoD9Je
OMdQqrJombebaHWNNxiz0HLrlWiO0JRSRv9jWRfxEcGvSNeYoHd/ZkXT9FAoHFwT
xlSFAzwziqKKgvQNbs29pc4OJqlFuVBVfDPd/lC70/QhiV9bDjjGJ+DBIhU3mLXG
3zlSRE2caEUJJI7htd82lS3AObPvNWNN0jCh1Pb7G1dzA8a01aZXskbFZ0z+ecFV
IKs/3jyvpK5LePmirx3W6EorwTSSv5ygmovR0IUDF19AjR14z2Ugfhdh6mR4QA1a
i/dOy+tgSJTyDGRWsSUteF64cPA1106fT6s/Eyiepdocl5lKUFLnxOsY47XGWgv9
KdZRqhzv8T/TcveXwpe1rZPOnQo9JgtsofEfjlI23VZw/C23MKxJRIYW4lFK6yck
w+npchWLsL7k4sZ1+TW1WMEYYW4aV7r5ISo15pPJBoViwDOLh3/MAg5f5+KNjq3h
AFOTmh35D90qX4mkSSpgiId6ticbhoeSeTNaeUXu80FnzLtTIYH30OYlIii9XBBb
A2NT1ApQra+LrTlSy8T+zbI3h1K1oY5qXRgy5MXF03FXhacDHr4wdI5fzcpljOZS
hcYQIODIOOPSFraDslk/GL1IAC8rIM3vSoOT1IEtJYZDWmwIJE/bcJfeKu6pxA3M
8zT2FxxNc1AKju2En515hn4ql3vnRDLYFUQvbGgl7UzTqop6f1Wo9zl1Ol3/nP9P
hKcwqL9nzSxZp+wjpJWTXwRfb/PJra3wvcs+lF3srAedQ19tF0trDVtktRj0FpV0
vlpebFZZC72zrj3fXnEro1EZ0ErkCQZpSn+tXOXxTxw4tFuJj4bshE7/tbkY4Y93
O08T+vnezvPdZqRIPspS0eLIxTCIXoF6BSuAOWTU2O7k63172jJLmhL4RulcYxm7
YtxuJaVLy5FRBcDKUxpT0Y0u+JxzszYDJkdhfTUZMsgeeCjBI71NF1pcnU2ANw3+
LCp8dtm22vGpszCnI2DXLDjO6alyXQEwyjqobc2JDnlvVo0FOobHjwaWMxWHlfMc
xXxGEIYaHUCHaamJ5gwgYEuSIfzX7DEMcys25Ra5jRUt/t6DrpXvkh0LdRjLfg6e
CzFTVpuPV7eQ/3vJS2MbPc2J+T8pheVAaZX+5dRQiLnhgA0VAVDgYB3gmlCtNGYD
mMMkZEQ1C11c/mgtzPIgN1PG07XMx9TJeDDyD7hkq8GivV4slfFH+JI79/dBeAfr
7H85rOxDMnJEmK2mz5erojdSffPB3SU6+yKBGwP1BlUQopHWDM1byFOMsXLz8IRO
gFtFuNxU0VJ/UQLuXikyyrTktCbujwAElyrVfg8zBvtBKbnLEFB8MQAFdGA6dZlW
1eaKjbkht7gKOgayU0WL3Ec3ARQmHtb1XEORnNNEoFp+sMnVV7QL86Gg9dAjbTfK
HsdzSOdAoI8XKp1Al4pr13ZVfxS2KH9TwezKdWGdkCE7eoCubnngLfz1bNvNEGDN
Q9Hwe1PsqdUdOslN/xfU/wSFjNfU817HJrUOSqSlt5NFDmT9umoOo1CvitpIEcms
E2uZgQ1Q3NVGDsnpboj2iISRe0w7biOHiW+XA5Fp04Q3b1OEr2mZ1Cq52jrM2fAD
29opcqMnNEpp+rYNTp82UpWQaRxjb+3m2xa1RnrfXJuDomxWEgfZfmMqJDF38TR9
R49/SRVhQ1TaUNdOhmqdL1TbKNd+NM+pcuU/jZNO0Hy+H/HBoI3g3MDieP80sbyf
9F2WaFFDNgUDM+vZ2UOtzKdatoJ4tz2nklDPNYZV2d28mlge1tj39o4TFAdA9n7h
rWyed4cSOTJSQr5RKX/lI9xVYCzlZhYyDfOsO22kNVC6HZ8Lmzc2JfxgggE887kU
EhVzliTHk03ikb0xZ/meIQGNrpiXAC68a2HCr4D5VeTjBm2USC7GyvLnX4FaSOKa
+GnwCvOnkVVPDsErO3N0fwBufU4sfBF8WlfgLOYfqyVaOhPm122uDovd2stBIXU0
k8aDdWVECpg2TBbf6xhAfzo0Om7mLxpr6jZChAhPbJAQL2FFlhJ2YRIX/GQS0Va3
HU/uB0B83/4S25H8/ImnACEVkeECIJ3JwU1eyBU3SqQX2+kf1tn9k72/SM6Xyq6x
7ICgocULZR8aYNGpmrB7ol3eAluPaPoni2I8Pca7LJ/OcY2Eo8oPjxHeDd1D4KWt
xmjtAgk++Kz61AXFiPHGcnrY25xr+VCX6q1WLjNTWc4fw1m5lZ+DHkP/snojB5LF
I/9g3HjaAL42NIttBufT4Uxkv1YrnoTndpsAZ15GUPOGEy07rdesUKUBReo+drjd
5jWJXyZ1suH53Pviyk+jHk8XCc4errr1xN2w903UbD6k23Gpx5FFRnIa5Qcka9n7
g/B1VmTGcwZOK6pUCyK8AAK8obCFaY5xXcJMw/60qr828Bxc9Vd/ydWFuDgGuvdm
H3Q9BMzgItqTw7Nfo7b70BEstIQzSz90FHbJTOBovfXhm+qfnHCjQWXFdr8TddT+
vdjb4kHMOyuTcpmKbW2pPKu6yq4spnb4HLkjtP2SbkyT3QsmvcM0C3RpCeMJYum5
nGuH1G4/vDjo2usbwzdCtlH3P7LGukpJ9aRIizKwvvHL8MLJThcX6JUXlTp7EVjK
Grexx3X6VGLlrlEizieuI7QW7nkwFQxFFEQo6sSE2lgo9TIe/mgmyxUQ7R2OHvbH
7S6iGoM3GX/KsFqTxWieq48dyq0/SUq9aFxqFSmL9aAtF9BJcE0X8+8o2HHyDiTl
c6hJuv5tZNrHFqj8GC8JwcH55dfmiZQvQWbAdx84r2sUvDUZ+m+K9Qs7MnxnyHZk
wpba85ku6s3dTOxEHw2adwA5zqn2wF7H5ZpFRZkdxyKG27r7DLUNlHtEn1fT81l7
AD7p+4Esb4B/LMTm+Ly8xMaoVBaeDPk/S/2O7zFC5XFM/0JQONR+iHqPTunHYdbD
WTqc/NKuRtEtggZJUWGTeofttmX57d0njOBTe3tbhmX+1/zlojlWH32qrXUiGy3T
AzVdvxs4d7y9Z/1bv9sga2g6IA6HMXci3i1wo+o/GrKNtJvjpmUK+F5oOLxq+bLE
0Lzd8LUwSd6pfSSK+KSXBI+tStQyln768S8uygi6EvPzANyDdcXmQg7VKpKd0/Cg
BrAxP3ChA5RERb9cv0HpAUQKIxJKLNSVCu7v6e5pBoFJoZbcTgHXZ0L0m7SA7hNy
evaOmZasLb/bg53/3jOBQs3giL8zLXoZ9QDhpxji7i69Y1RW4BOEJ9yOTVrit2Ve
JlM2nsvfUUbp4SAu5veqhpIsIfyuowFqGhDyT7D37Ym7dIyUpAYpEBt0X61hK6IN
aE1Dt0/C22woCQysjt830l15hPJV/58f2nXtopCE9Gbcc+aIuRp+ZrQ6hpXGxjmI
3j924QWAR+a9BOlF2pHppQyjiwES0zgoWOXAowOKmna3Hu6q2nrVtygQrcPUF8V7
rtySkI2/jD7Mt+X+j4GKQMCc7wzeCI09JtO6HfG43pcebymQEqMm4LiQNb6IIEFV
DEspsTpioYESTFHkYLabKBdTTM8jL/3ye3GYorJN86RezeF2Et/SiIkEiAW3qdSF
L+lRxr5ih6FO98ikDh1NYs4+w5H3ei6avukofO3UbvpO8taGSIs1hsRzEzhJjVnn
C7TldrJUgJZkT2huON820nSPJ2ilxVGgMXqoYQf5Qv0BGWKbtyJXo7xamhbOEQVL
KUgMkzZBZoTv3ziPqGednTSJxJijGHiExxOeTmx8yS+hgBnl2HgocHbdWdSo0eec
IYo+Cs1gLnd+I1S5muT7oaOxMXvoi7cZp7CLM6RsRPUpt9Rixw78cr2tQ37JRvsB
Pxac6jDtCjlAHZkdeBztO6s9krbXoX/5hD5qPj0X9KxiQID4/tLQ78lnLkkSu4vZ
50UYX6fXqkA1eh0ygU2j02EwLWpGB2tqugtKubbEaxLuR13D10PssptFimUina83
Z6kDYe64usXbOesIfbXlU/SnSPIKmNbSFjHcERW1YhTulaOff7wRl0TTIAJC0PSj
K57IWB+OfiAEpPMnUVC0a5OjUoxOTaW/Lj35f9HblBi5BYoqHF/TOeVqOwaOAJqI
1ZblWz21bRdfHWQy8JDcIUvhZWt3obo37JcDSDi1V5xuZprxppCmAHwvNm+QZ4z/
f7r1PRZE+fG/zn/yNlbVNok/u9n/x8YBncuQZuN7QL3kdIsFdASWLBvbfcFZoVTF
tVCd2w9PoaSbL/XmnhjmuUvys2w+pQyBatYBIGr1Z9HPNmeuqzkahopA6nFTK+2A
Y0XrCysCTwiWnL1+qtublEKmRgfLBXE7M7I29RXu6X/bGlSBhSZbHS4MoksFZDRt
BgVJu5Vhx3nWw8Qql59T1UeRAwEJ35lqqC8jdsGlrN2wRAfRxdrhVYpmp311Viad
2Nes5DZ+HzTnxWelek39+04LuNFgUFcrAEbx5Ei7XOnQxs275J+Sh9AUlYk4toLg
L8qznyX8cVnvFQQAaIGEmBTNW1hsVxNcia8NYFPL1XoscYEfo2oRtQW3KBKnrY1W
gCkHchhf/tnwICdxNMta8j6L0TEsNimiKlwyEwIhVxmD9powqqTX0neVJgOhDpmg
5vxxzTdplo04u9pj3F76LsQ7aMh1JAvurPsL4u5etqcSrkq1bAR3QkGPH8TXtYL5
TdqC9/uXKHX5Hvp62WefOj5S8ot+B5wGDuYYcuxd7+XxjCegO/l4N38RiFue/yux
spxNasw2xj4a6m7aP9juZm+1GyIawY2jP3TC0MlBd2tg24Crh8fNGQfF3hU40U12
zk38hSe+hNfA0UzTnyrnHn0iDFXzXsEjbCZR4wwc+QUaoKpmg5gbttRAJN7gp03c
WD1NxyJCKfGDh6/gZOyyVM2t3vzAu7qhSZuiTc5bEuuhUtM06uV2rARaUHtg5L2K
8VitbG9tF8Dsws10kgwKad3un6JehmGJqFShQT1waz004krh5kswj4k7qXrj2XzJ
RuEuG6iiT6/+J+maI4pcsZge78pGwfv31vWBSSVh2BsUDzouOrPDHqDe/UR9Sazd
7gd6MipvJWg5SRds0s/doFPh7Sob91/slxr+QNK9i1Np/kewcvI+GTK2D1lWcdg8
yJbT5CgELhivl7+6TXlNSM+XQwIzIMmoacan88/49n2VFK45JIAGhfbRMCxnGoFU
wz57PUvem6X0yScn02S7/+txlR/QtWB8MAn8Ja5nJ/iy3NdF2Z83VlO4BYw1YaN+
+hTR7smQOFGDB+fmrcmy7IHeYHP1xcFqOaVcYNUXAyhLJ7Z1athhk9hhrEwHldqG
n8Cu9RR62wdhQ3B+rmU56gcAFW7Wf4Qdx7YHBg15mXS9sY66wq1Z/OgZQjYZWezs
HbUIQE46B448q+c87L9AfONktdoMZbz4hvl/qETDQxFzY66AtTGrsNn9ZOTz1FFY
ONO4d28sqodpAmoQe0N1PoedKcqwbbc/nTsRZaoKZvDIhPO6at//XbMJi/RU6WD7
nkxs8WO7v2s9rr5ckyWoyXyKmytzGnGm+fbruRGn2xZg7WVvB36sPP0WaojBCWC/
E1BSyYqjR9wLutfoCYnEpdiV3GwZYjYKpWjoNoyqTpYXETeSikQKhws7bfYsOlnA
Sgfn6DATHrOfbiWP+LkAg2l7u28pL1eSSVJ2poiBhEe0vdyoElJsvbCaaD/syiWO
wdaQUjP9GQl9VXncabI/mwB1DXOEboau6LBPZg54X6ndumhnCEj+wXK1zxQsyTaX
RAb7tNJ9s9a0iHcEs9xwhphPwMLlLBlDBHVWPdF5zrfC/230KEOdUzBwYnuWrG4O
W12eICLjFoK3ADtl2Jbv/SjBXl9FPK8kkdVisXehQBIAm0/hv+hA/tVyumx8KYE9
yo6boX3A6OB/4GJZHsFAhLvGnrtcybXUtIuOX6K5yddvLyqquZDWv7Hj0U+KzzK8
dpv+B/nZkn1SmHpjdHnOmRDuqaWlzg27N+jFSbfm18yayvyM5+vIwe+nKf0tiApy
8Cf4oDSv1SHYUAJvDoa0GJyu/yIhe/NUlj+qyEkFd3sMNeF7ZKO5NeGWZ6vq6O6/
S3CQv+XHcLUEilPHQ8C+H0XiQ0pHQoUWKxfScL8IdISU2LLtdfzcjZfSl1udVvu/
qCM5ijIuXoduPUFwfjglY5casoirehHL81aGRCD8TUHdl23pMahWuzKUnOzcdu4w
gTleMCU0UKoBu/e9pR7jEk51baCDkjNxFglIvRcOg7eDb3VeFG1ebrehSGk6c4S6
7cJVPAQrWx9M59/uAp5DmbZzliJPH2SlsC1JqkbMnjuMIZ5NgppIYSl20gHfNMJH
FXLPLOwMnvxixHgMqaeTH/W0Ak3IsSoxGmlK/E7knOoX39cycCGe6Tww1PwrUrzc
mDw95Gjots9HcDGsLtpo9tFvdJL3AJMO+v/oMTkeuEdsJeo7hN2XnLVV0gbv6tOH
GYbfOdM+O7kuboJ5W5eMjC/u9lkg5Vprixl/0054365tX+yNi/ciSQh+vaxdneGk
gRVbus3q0G4SorJgGq5R15E4/BmgVqJJzrRfDdR1QH1ynei6wLFzethes4oJxBHV
m5KRofZewC9rco3vvu5oDpPf4EZhiG0R8+P1grZZzU60D8eBZ2WRQYusJY2NOS4m
mSGtnw7BzMV/pJ6s+ISIBwz6ndBPwJRsC/dYp2hp+4JDhHomSCLUvYzuzHrB+zKa
p7UJ8kkxEd/tvnd0R2gFr9pBQoOnUO7XVmkiqccvIUq6O037Ex783SZi0FikfoIy
8cxDGNH0PU1gBfjEDKT3l6aC3o8lVedtE8Ov80flC4TSWxJTWrp3hfn2KrcjJNqq
B+80M/2OrkhS3WzHtmcdTuqM8US7iOX1KMp7fTafXSchY2u//EMphzC8ytWlu4GB
S6gABrsZVDaOa+jpdR649yG5rVs3RwP570sciV5e976v8QwACPVZTrKSYhms0SLZ
JhnMFFMTUAGYuSvnZyWZSah5xhu0Mfl7eV/UFUiQRljMCWX2YMclU9r5S1tmjHrL
sNUigR/nmPrsfTutPe4DYX8SrS98xw62hpZ+6WvD2W5mqkM+vT98+ABPRG2Lw04D
srjHlRk160ItKU7hwnbJ34AvWussikNZDcV6OZdFTN7bgrB+TWFbYvr46+eJ453o
n+HeWOe7mkKxRIESI29EWveVO2n9p97s6LnV2FHnWoz7BqjlR+LsCvg8auTL85mI
GOKBP50Bls3nnmKsg5D3gok4hSv0xwTnIBCNoRQi3ZDaxZluzRVVpW+b9LOKxRO/
sjcPYU2oo5CzCOYgEF7R70nthrs6I/pBRDBmQ7LQd0RsSddXF4YSwYTFY2Sxnnvp
ngmYDGgmJA8c8NDJu7ApfbAj/hqNMC7358nFk29WDGOzjuJ98zMNPk8YE9s3NCQr
Shzu9PNexXydqkGOzLi09Swr4jvroA5ILg8WOi4Z2fsjPWWHRvk3o/jlIjSO9UkG
RHW0qXh8NIRfF7LXNYQ4i83hPLnlPjNB2Q23X4jSCxPSMY6f8gHPv0JCwDLIFZMX
RxDLJMsmT3xNAGOumJ+YL7t9yQdNdj3mZed6m0h/dIo/sXrkRub37cSjJxgEwB3y
QuDll0HNk0Qbv5zhd/OwlEf4A64hFf/wS+b9/rKd8GAhpenOskQc4KQd6PLAelWN
wLj+yoDagPIs6lH2L/IDPp6ZrZAvikR/ycSEvn7uy9808mZe5rb4WtcVEsuUO9QV
st39CQrScOPzGrWHFieiz+D+YkP7nKOTAeJZYMGfiHHCbWE3d1ogqvj4i11ioywS
NNsFnkg/0uxerZYClRZ+QDXGwbjwYpCyrAXaVGtKT2xkQLcLAjF31d+B+DHImnOE
D4hEyoEnKbPPdfFE13FKoAWenjNz6iLdsueLvuphmkLDGuUcOpBzWrvO/nx0u0MT
UrADVRuKSBMK6MzfayR1NMDeN2aXgY1d+F3sZ5qCKSpI1L9u7v6vSXAcL6VHNONd
X+2m73Q3rXb2lgiUSvfa5i2qarElVWXuSTrsBe1uobSFv4iloV1NlvDVmS5BetpA
F3MpXqgRLAm0VgOxOAHBgx+OG+WaJ02lZJ0A3/bDQb7QHgSvlGSS98cmy9Kx1kHX
lLNaKz7wkm40n7pBHtlImSXmt7M/ImnNBmNURTSJuYPkuP2Nl0+D0gaCPFCwl0Px
4QRv6woZaWneNHpaGRgGikBrZjbh2iXStpz3Yvl0WbcO1dGMBj9QVeVj+Ymn8E/x
P6MKeX4qXAuNV0QCoUUfTRmJCaouxIgQ/vAKL0egUsiy/hQK0FF8P/qWWoXar3x4
qea2FKXrb28R6FgwPIeNlX19Os8P9UmaUqAqm/BxD9dgOYjrFQDfPeHyqlc6K70I
GJDAgbdDTgH5rQ8Y+Kmm9mY4TJK3OtnlHdH6tsSLpFPbiod413dF5MmNOQ51RzDv
CHnOdgC3dWThmwBnyPlvgQTUO/UX/VJxlzw5kTFId/6BvBfRwdjiYpU5F86dQok1
BrWPH3JghEwFUNAwK5WaXacgPSiTWnMCb/GHFzEF9W1l1qF8m6EavLBi/kzU00+S
+1uW0odbhkI+Q1fJpsMUZ9KuQJY4pr/7SXFk2mQhVtUX/z1sbNCdionR7QISy/gY
rc6EczqT7ZsHJzeH7nLMJbw24k8K2lH3D6CbyDb5ySch6IQzFOCveZokZi2FOu8Z
Y77qOHcr/unfKjrfd7Uj1ejhlHSaI6pI7ySe3m2eSfgxM29xe3Hykdv6rKC+aakJ
Xfwudx3l7v6ci5XgWcu2HXeM6kOSoAj6kxlPZoh//gGoaZ+uXbi5k68Hq8qsymN+
dYpdWEAMXnaA3TA71lqWDPd1vLn7d2NlrZYSZ9iukH7tThlO18TifBjDg0XhZ+Kn
+c7JJTZPvfy9wytv4uiUyKDqGU5bGs8IpvoBXEfx7PB1wlIgt/qHvljxgZP0Gd8+
2VI5xpyiP4LUMuwTB2uBp0zLHw2FEJj6yC4Ey7S/4gzp9vNlpp5GsgfpyIvIZWgh
KqY1wQO8n911I9cXP2MFxNUG1TY4ztKKtJMMNlap/z5mHvK3mu7JV1l97QUvD4f5
o1MI4Q14mqfhnpF3BemRvVR431F7LiLRgQEU/KuOY4O16X8CZUYzb5lHeEQCjbkv
fEDKAATs4bbFHgA/Syo7NVnVk2JXE9FjJ4C6u7KYpeqN8iEYDJO4PAQxeF9Ln3DS
YdrtosEI9u8E1dE7NDKLGUSM3tbIrg7K/EukxkLE8eQL3azjcSfJvoqw8akyfKWp
cP7X1bkPa0mUbIuuAuBpUQrR6JrdNchCEO1qVW+QmTLbUtMM+IxkTVcPRH91v7nk
p9au5mH2stw7wzhnXFpsAjzT8dg98Go1nIz49V/GlvQ6+ztRvkTauws4GMtPks9S
RmtbR0hZHYbmCLHmKu0a9ZmhbtElbq7pE+tUEbKbsVhrg7MpiPJEXVRYs4msFGET
kbGhc1fxhnxAYljVpCqiDWzxrJ7Avgo6j+Wwlhy4c2PML+X0BhOlpyMWQi+mE8yj
SbHPl+k1xkC+QPHzpGPvBKTt272oKaqUVoD0gnanJ7kAuVzCeM2uFy0c/Xa9L746
MDYR4gWjvKojxCyaZgCjy+ixGvROqCVporJEGdSZ60tc2z0RzTm27/S89Vbuu5Y+
Fomtc4qq+BB+bgr46zPSr0e5tZfHe/FfHmJUu9xgePxomKBFKA9k9eGG522MNhKP
UvSpbyStXjSku1k05R0QXovX2zb/WCFP5aJKsXmDUyRW1/tX3kAsvmWpuQRxjz0O
zQT3gEBIwrRxMDi8tDiUHDZutaa55G8WHkMPNe2hXvJtJT6FNcKWlODBcekR5DaN
5D6ZeVzxXCbmyaSwX7WNlF9DNIhFTNmnCXGcFOX27pNFv6cIAfRxtMicNfxDJjAy
VymGxj/oPtmWaH9776vXjXJyjlp9Enz84e6wC0ZeCMPbYWiz2nX9bXuLrv5DA7/z
3gbMBEbzEXlqxuWkwv7egDgJM8OHL/Gnpi5tnfPsD02LRVoU5flQKHEMzwZqGa/D
E2zKCpNoUmPgUjM2TViRUCchh9pM+07tYnay0xCULez7Fzq+BYuvIoUevAmOH9IB
q0qAg9dOSblxe9FHHvsieHHUOX5zQiljeZYrqtCQWasKusP0uECPavAFsKouMKPl
7AnVjAT0+NNtnAMQi0BbqNxH+N7JkjAAUknGBQ48pTcOII++wY8Str0tNBrs5/S4
H3UEqmqHdolFFgT+w/msxk6X/aY/BDi1N/t5sHmC/MCpT+pu8tCIZV+pObFxXWlU
s6NC7kG5JZ4aVLS0oK8N1CW3bWVLYsQlDY6c5eEHenSu8R1rJqFPEgmKWci7N6BR
ksqh37ZKjC/ppHQwtCZ+SArWRmEaLWnTuHZqzijbN0Ax3QLXJQxKZM5Du3Qp62JY
nngn+ekF2KXFs3PC4q40g90ZRpQoliTSkrLX4+WfIOLSj6QDSFTIWaQzad4Vaqk0
jHbVKlPYEBtRSlYAIxPEGImmOWOZpBz2qNhTwIBTm0GYuu4Ix8eYpoyXKDyV86Q0
S2S2FgbNHc3JXG6CA7HBMwmvZz0ZWm2mBU4qrQNuILE6RvVkxRzw4qtOt0/4fCj8
fKniyHJDBRvI+DYXIIf0/NdrqElGkE08FGxu+W4uS4++8VuHyURb4/gLCuDL8hWL
e4EkIbU5m+m57M5PolcmoyA+GXvjnanVTq4bV/t9XMQEv8ukdq2YN7kfDfuKD7/J
jdYL/JyMhnZfXKUnVXxhrzpOm/EeG9cXu4MTnth1cK1kB9f60hrtvIXXrfuMQau/
rY2XSgcDU+9JMbEDh5rP/BcmUZU0cYhxKSEihGh06wntqdNQo2I8aBrptM9SQzf6
MVjeY9lWuhBqnQOrR7hqI+FZXjTva1sjc/ufXHhGJGyCbN92XUYC9JZJdWDBiwy0
KcobVxY2ZharXS/ysFo+HB0UM6EgpFONyKdxPbLUPeRGKukDCQtJJFNPB4LfMzLq
rv438T3a55r/Xw9xCyHSdbNG8k68dnHHG+iI7NHAdAVdQWYoN1JIhQZPmE1WjRzN
1b0jTiCBiT29RxXsOHBPig6bokGhNmGuhDQehlf14yuBIg0os4X4X5wTacYcySS7
AiBiZ/nDlNhtxgl+VJcJoT2LGZKePKD42hlw0877ok/JWvY101U9FYsfl6kJfyHC
P6JgGedNQDFko310PLhbMmPaVdIjvt6UYJONXW2RvuDA8/bgLIJ7CFc0qsGIHu6Q
q4t2oXjYMTiTG1n0M5EHCUXZ44gbotDTqVQ2ryvjyMCrIYZB5o+pX+8OB1IWopgb
RIc49/ZvUoyH7i+O6waJNj/cc+E5BX0r1xjvZ0jhURdOh9eILXE10DmfKQivPSJj
ul5apsTurZuNHd4kZ4T99I+N9UYku17z2cYXBujjrMOoSLelaKdwyM7nicHiVmru
G70575M3r8arM9uYpd0upR7tyEDbDjKVQBpQETEvIo9nn1f3vefIXois7VAauO7Y
e3nx/z69bRy68HmykwaZFPRqKDas/hIrNZxxVz322NOg9zwzqku1M+G5roUv6Q0b
Q9nyrnejnQqPYOgh60Rn1PINug9wTZCuHd+1FYCpP50m320Ckc1xt6qZozqNATHw
oBzTHF4qSh/mJP7uUmToi8pFDFfmnOaN5qr4huqMkViKfvVlQvRHo4uPtNXIHtkb
SFcfJPUENopAiir+xtClFKJInueZeU77mexsPWipDbac1wfl5f31MNkDjtkNGqrh
KBSwi5ykJ8aMyETCodr+9yeSv1tvBLg0cPCtuxGU5g5RrCVAtCLfSqchf6j38/YV
s05SrF0HheeIQeZt/uwqZnaZCySXJ1JLah7eJbeDnNj0mh0dpkW6+5RH9qilfOqt
hqGVk2EtW6dLG/Rn1UU0+IyMxPNzSvbio37gIxyv3M3qiZ4fyMY7CoeGm7miA+qk
pJuhELYKUgbTvKtPTisNcX2G+TLrq2D3HKtpVID2VctbIm7Z5ya14adQf2SoYL/z
tJYP6980JP4T9bDcITAtachhsphdYTPn84pa9fCYsex5E+3dM0QxJqrHMwyr51Mu
uCuSSsVFQB/MXxUyb5P4W5omrwv73U1iXTD9viHF3y7dewSMhGaYI931YcY+J8Aw
4MdK2V6l54dUjpdvYd1mbcrih81ixr3DE196/zDHeieiyy8tVcMM+NhHuB+WSZH+
kDQNdGH5ehTKyG4vmewHxOTi+TU9pnf6CrrktGEUkz3EJZNXtlWW49YHy5Ba0+lP
kJV5TftginldXk8JvnO5nnrc9/A23KHPTbbcqXoBOtUrcum0/QS1KlX4vW6Pq2cK
fh1HwfaZKdzfOKfgz0Q8ZupluMH4BDEZ1cIjxrz+4Qeo0vqzlQgacHZeAFQUMy2T
QHbZs4Zq1GelxIJYS6oa8p0ffHtJRIizZwE9vFGTCLEN0y6+k6Xy+I144gEjNIPb
/hJnqXSZhleAdZocb897G7WeJXhT3cX45k6oqymn1iP21ZL3hn/iTrjBe8VtOiPj
Q2wAnmH5YCOjpEBz0Vsh9CC5FTP2NNBcPqU2AH9B5+9Ol9cjlu2xGS2ZRIH1aZK5
1v473K5Fks8ajMZzT2rmuFg5F8SDoMTAdIBXkpgRn72DmA5iQKJPGAJiGD6sWpwj
yKd52ujZv+pilWB5cbARtjXMjJDnMgbEk8fNpMtCOuBtPC9mBZoCgOmoJ4nmV6r+
O3YNRGCNwkbceivuYwW3LFL7myMc7H0yEZlJvgBd2ARGzjnO3D1CjIcJucBTNZQq
PHgfZmGoJRbX2P5O5O1jsGaoWFQz3Mkfdd59yJR7tyDIi+aoExdqqyE84aaPtr5l
L2nZJth4vvagUpdQK4uhTWPIOYN7ACHRVK2IYMkVT0ZnaaoevafDbjOhq4HywRD8
vSj3uQXkt8Sp2msvyeWhjE6m8Q98utkungnJnORHebRDQ3r3VXLcpI0ifzuXqlsJ
VShaYcWmD3WxJZJ2DwJblyVlIou/cWvM/gKEr71dwm1MgbpznorG71mExMggdg7y
ebzDHKvWILIKlF2AWKGkJIai4hbiDzTSFlFBJp6HbNBjB9+LcLClWaKnKuR845QV
5mKwUtNox7PGDHUktmTj3+ngTV135pMkgDboGVBJbyMMapPFq7uXMVMexhRTHO/B
PpfwuidLYVLt+mFmBUUKETnP6obhqiblek6i3+FQ6wrxUrRbHMmrzgxNKEqwNhpI
hVePHPw1uasCZEOWGqqGRJB6r1E3p0qdph4ul78VTCRVwXH5pQJlUJJxVDnC4Ye3
6OyFVAmrfJtuZNnpJXV6H3PZKJ+9hSnjDqz7qnNyzCeXtS0Xk3hMuF6QirvHkRzR
Epw54a23UTEHcGJQbe0zZYB1YN4rPXRH11BLsXsvGQEvdpbeJT7hOjMrHjLtd4gt
an1S2JfSNxBc4lPRazUEHRzWnZTTHZ9QSnuLAVMevyO8C1HnJ3LOB2BAJyZzT0iw
JIWuaJrYp0cNJoDV8vuL8zZVt/3+a+ySdCC5XwOuv+47aiDsQLle4WprVr+uHKi1
sVzxle1Sb2nXxx3KuMTgL/70kHiwzqaxiMlNSaeoUW3NINqIMczZscfRgGzNpalL
Ptr8npFBO91aSzkLj4yomo4dryGGI3p1YJtG/i2rFXdMN8kgTch3kQC42A89n9zN
W/PudVYXSXytYt7hvdWidFy3T6SJ0OgGKx/hvujqwJn4kIM7DEyyrMzDxUTb8TUc
DcFWlg7DZrzJvQoL45FCzzcfGsmA+L9HX55Gbe3pso3Pm9KV5mvCCSYz5L3yl0lx
S06hnQ44J/zekk15NY4I06Q7PPEWiHrt+kAmKg4jY/F3EWNpHhqnc5/RRcS/bkcs
i+uKrokFErAUWqZVKzcNiZy2lKUx3JCp/oWQ1WS3sUoACQXoswJGgyMQpmO1EW+Z
SZ/0MInYr2iwLy4BrcipuKk3wqu9/fW0gXq7b95UkD7AiYzos2jPx/NojLAZ+rE+
ys6iJoekm+BEQrnK7ou3mJPfVPuQSqcioRLtL4RgtCrdcfqi4UMAclwuoO32TE+1
zPB2VtG1iKK6yyoXf1Oq1UvhTh80G9lQpNEyt/G08w2ZaSQmMK/muE6AnyIX6QA6
6/Diifsz0C4XaKRfLZZH0RyTGEy0t0zzbCdogBRIHEWaUbk9JGaKx80z3h/SxWHk
HdsKeweOLhlCDs/zswi6Ahb5rJJcMbADJeM1PUcgVsT8Ex1ohsUU7P8bcGVCrwy1
hfkTE/XmyT+h0IPxfbQfrv/Pbk3gIq9rPKOtRE1rgO7tPLrBlbY2JfVEvzV0GM/d
2X3XbC6sL/hwMLM4F0U04JzbdbBTFJaHNmPbYVIiGotV34gA1Sw5ZMcxF1AuNOb1
IQoRsKiipYt819u2k3wUlHxGUGt+3PY1mf5CUyGSP+QiTFmCn5pZ/k9bE/Qzk/hh
SLjr7aW0gGSzqxwTRyNs8toQTTnY+RHnLxQJcGgkrCMGcTTRfalQKyepiFqMvm/9
Xvw8u8Q54lc7LX4iY39pbiM6rDIMEaA7DkrWIejInfgbFAtzpS1HOOO7PEat8ICY
9UN85QpN0GqLexsihKm3jwFMKPqxu7MITawxyspkv9U9ZWZgRrJWtlWNikOFnwz1
TYx24yx8bJag5vYm9kS2wixz5J+Uv5veIBYfzqlaDyXLoIeN3Mt6yZJuqIaXVTXx
I4KjTpF/feZWpuxJIrESwoSC2z00eKFgwwn0GYaohmfz6MlQ2PEw0xmGbkns9NTp
xDqDg1qVCTe+3oeuHXtZQVjS4ESmIAKnanUl06N9GDq8uKpg2+f66mqCA4J4DZJ5
MHCwVusYm5lc0tQLeCvm0XzXQ9ygWyaMnlsKdV56gADddVlSEWk5WwvqTbvafJIZ
Ino/eXfyT+Q22uE77Y+6zjbb34gUxlHsKTNcT7yT9EGKIR5Gy87aKFtX1j+HJxXc
r11R4ZjqdWc3+sso/qiQjPmUC3JgpELct+vMKbRD6cbsEyRz4vaGVaaQal/LjKJz
LUF8vocwPSt0JEZhYMd8AqYshwTQ0m8TFIai7mICsxQQ87zBVJzmQl8Iocy8VWH1
tLYcxpYPt68BuBj+pe4owc684ZC1+/4wIEMoOaWQPyyePOj3dBBFGZOE5hEdVpcg
XAxX9Ne9sJmOKYfswK+K0iAVHhPfhjsY4K4M/cbh3+yPt8kYW/MbYS0AXdQRZZdt
fMZ3/imzt1jSGaeX9TfQAWHDIZKX2zJbALAMla9UseCA31VFiwFFjpm4k4ZqUg7a
XiLa6O0tjLREE7x0LNTwfjCOs9p2ZcbsRqZ5mf5ULgY5KAhl9HTElz4kRh4KYagt
lK4wqe7x9GirJIpEDsRGV5IoolQ5XTEJt98bBC6aargMgYjT1iHsJaoBKkhj2db6
n2+tEFyqWUbRQ02ivehgDggzfNtFMjmhyBVZJi9kyQ7xZEv1V2sF09GsCZofLTCg
6iBUb1tjUDD/qTeiYZgvlzcpOd+Ste2Z8pZiHlui3b3wQqsyBssxXlgBudNQJEYe
2iLzUrIGZWivBmbaMqbPQUbMbzpfGfr/pE0TF6j+6p+1GdIlPjeIkh+Jv2DIzeDn
KEIup5tRxJCuErQFIXvmaPFhrMg7g/3ZmV7v/95/K8bCrU6rRdIgbXNEs6ME97Jt
pvpA3iD22mI+XHFH/hLXCgNs+SBrE2A7sOGonULAod6owGxpaxcXJNM94hE5t6im
wO/MDQg6u7ZqdI9Q191fP2DN6XE7oSzW7V/Xw3mpwpELzSZkRlhHAhzbk2/O3xNA
GcMVQz8VT13jqDt6c3mW23+04IMv1fBeuNkw+7szGIYj/3U6N+jmukhkEedNIub7
squPi2a/UoKLLh4SYT7qpD3KaeKH97TTMdQ4sonM0gqWSL7eZ7Dc0sovvK5W1HPA
hLbF58YON3oS+jnBY/DgZLkVAyKBordkR7jKlP3pjL/SoWyQVOyR7ba72EBOrg3t
fS29sj7jCSajRXH8DNoIzpj/T0j7jAMqJYS3KOa126XWOmY8win0vgrznob0ri/8
k4tAsaE4cfaHFWQNK47FgzBDoPTbUqOlcRlEvsKd5rrh3NpTZccrbU85P6E8+tzU
eE44FwvZpif/h+bG/TRLz8rN/A2vhUZNXS+bMlizC+zrHVI0VzhO7yb8a/J44cs+
0kDlJ9fgm2ILMC8y1UdZYvzE1VNtYsjEoUbc3RN2zk/TnD7fUmNzfdbrvYKcu1dH
eh3mK9BEeZuFdKnkkAQg0iyYoYuB9ebeUZdhhDAUtanfHvDNclK75O6d+D7xl1td
Esyhyv5AhEZ9ZMTRfsGT8DfikHKltb83b3Rc0983R1d85ahXWvCY/VqMtSkpNkhX
dy7jRpQaBPqGu+Oj1k9ycc187v77rRI+ad2kxk5MM7Wp7N8hNd770fsRmTRk0Mxv
qZ3gKkt5ZUnphkUlzhLLzByyAc2GAkN4jxoTe4dYrgcd4J/G2UOTThq7xH+b4+S7
0vSsewZOzIWK2EyNd58A5dGMLeJWtDagNu6YkjWU9491ofqlDqU2NmmFOCdLyis7
ftxKmFB4J9Cr/HzMIuXHHxYzVjYnF2vMDRZUL7gSQUc+jPzQPx1cRlCseSpmThr6
aqbw/FASBwI39FMgI8dE1z8aia/S5CD7hflCTCoKeVTXUH5mHVk/nZBty/dbdeLf
xhfsMsL7dJ+9EPhW2KSAqNyuWPNmTZTKEvAzL3/dO0U+fngX1PeTpjHJf46lhE7W
f2xSt7boKQ7YjsDKV91DNUM22o9QSBmuyy7dHFpbjcrVNJmUhqh/ThbCTSYOPxGB
spvs/Fx+w2xBnJvzoeXaVqYPVt3vL1pHT0gPUv43erA7ikkhAD8P0i9+bGVJl6L2
AXIKwHzgWLQKT+Hw7xVo0qxE3kmSAUONyXPbucvPPchjL4K9VLD0DGhQEGJnAGkK
+CyqG5FY1drcuCcGXEq32GEjSCfV4irUvVxeQ7ZLiUSL23h5PI0ILIcrZeG4bPoO
Hdyio37PqTEuJRJvEgpjCHoJN8tzI5Xc4lDQsL9bQQS/RcMGKt6f3pkSVJK8526h
GwpNtGQfOUQy8gOXftn/nzH7vYKV+ZKvKayDCcniQUu7WiOvq+9ggsWPUvqJsfRW
AO0bpQcRp9UX6PPpPBHuO+UpZUQ4Fv63y6RBP5fVEIwjMGiv9TF8gLChC2r/3Kg2
4Wk6YLfT34MgSL6uL8P9BeF1/9SPKq11jfjzAhj3f8/w9s5I2wy969qoDdVqOM8A
0379IrIq1O7rFKtuL/kMVrl5SNcxsXv38osKrogOhMEwswZVZBZtrub+VZfY9QXz
zZPDxLUkHicgGqYflwzpPXwYUofiwthNvyXAQdo4BTwcVNEdHWUHheSk1lDP/06i
XdaRfjccbLov5eLeY0XhfqJFEXaOTtcSd2qUPYiOnGjPuNolhie86yIus7gJS+L4
KNJmWJ7+3Ld72nw3tBAwb6ouz3b864PTOINrGD3Zn9iAvMwNZZRLuw4TWFVu3Fgl
W3oh3ugW3zc+qxnNSOaILJAFBtP7o2/hVTE9BqT3YPK/U4EDCSUogn/om8o9VL6P
pXT//cXhO0UTon3BTeWX8uMTSX3VTeD1LctOORDtJEhZGillEKbIzauX1wJIRKaN
VgpTo1/qFJ15EhINwNu1pWSd30ty6z5oE24sNLsKozfCwIN5wmyP+3yODpT/WVgA
e58nH66OUPW7SUt7aQimUJfcsL59niyMPqO+vmZ38oIM7MJ9fiQsIJeL90F/ag/c
ISyIjqAVKhGTnEmn6yECP30lhDnbJpVQod49nkP4bVk3cFM8HwXQyGOm8d0oDbIg
tqnz/BA4ipE8El5/DK9SNcmcA6bHCOjDa080rNR/VD3EBixMlUacxN0Js3W30X5V
RcYlP5VB1uhH7EtKCbZDp6jV0bzkC+1rnQxeJrnVO/31z1teq/Drk7HXe5X6CBif
oszu/ZiVnYYGzoNMbPCXYs6u+SzRw+tjWcU2UJKPifK+0ccbviyqXsQmLu99eMuA
QubXxEF2pR9/MOUAG+tR0DwtX8axrsrrK4sHbjt64raRFF5FcrnkJTj2polu0EhC
s+1x+NgCwzuZNgqJ8DZGIdvgpVGLj1E4iXlhugrlufafeFbL27IMFopXA9//gAmJ
ji1XC8ab9AR+839h+Vr47IFksjwyxkvFDBWrXdyNShmZPTf0L0PIWUKCY+pKoAsl
1BrjPU6NKJEmfux3JmFrWRUGZdNACjgjcWkMwmU3VlPy2BhqckXo1fDMJLoU3bUc
mMFXuAIUXuDbkqQnbfiMnDL1WBjUKz3pNnKTXbeJe55UbhdkyrcAPJD/gc1/zkUh
z8QzLjTjEApO5EkIMDsXEvGpKdZxLwJehBcrVN0h4xi5ozsQlZ5DcEqF6I1qiBaq
8SNlbhLOKMjO4cF9/Wob+9OeV7iIyVjQ/yiKg3B9lKMoKFsi883dzBRadj4x907q
0AGJzdcdh6/maPzUVn2pzcmyvU7dgYCliagORiQ6dn0FUHvAnwsvGAgcfrhBz2CW
ea5aTE/grFxTX9GPOtDS+T7fPoaGoQoser0I5DUXNIAU9pfwncjSeMKaE5aG/MG2
QZw4Q7Vl74Uom7/N6UStGK5/bet30rMnXi/VIJP9QMEWztQFTbCu0UndAlNnTCrm
AetNEbBhnzGnfTB1YtwKfzIz7vozJpxhGbEBCpJykovOC4lkpUbByYxI7VaNQ3n+
ouuix9JkiLDmTuS+VpsN4DGWA543dgyEPG7a+gdlQ/slvS0IRKOA6wKwF2HOYisv
Jx7ECZXH6IwRkLq4FUxXQ4tTPV8PbXOGMsxoXY8vCeow6gImh9HYhVt1VZDNoggs
mo0YWzP8qw9IPYHS6UlfX/Ptvn4uL1cjMlN7jxS3hrbDG8f5hJXRhDGAeTq1+RMJ
jKGqBwJdT1PhZ+205fqI7Yg6rXSFOBxbG9zki3s8NVg2FnEeHDZ8ZbQ7T1vw/LGR
RX8zJde2Y/1zsUy/wNMeMmATWNSHVL60ZPkZfvzvz76bm3vzuWMS4XzR9xvBvpxF
3z5tkPNhE40fRT20jnqi/FVsd8vUbesxhR2jfNs7twA60yyddeQuEI41SLlXZ926
j2Qrl1lw6jMtj0NrAOv5+P61s5R8cthFbzsq1NzAbQ5g2Nfdk2diVl6NPWD7/3zx
EJB35ArHUOD6xNYnShJ1DUOxiiI88nkoyadlWg31FPewZIsZDXaPW7b9WbtP3WzO
aicdLa78lqf82xRjV6k6x0XYqO/lJFqlJV/SmZ5pAK3BulSBLxv/NjyKSnppOxCq
XMwRCS+6B6fRF82lwHUFXNOYyJ0ZVCUqpF+AzESM18C7pCkhNavMv5P8AhexwnQS
8trH+zvXtbMOC1EsSc+fNDfYScDQnSUEN9aig+n0VAO1C5P8WNlZTf/no0pwatrW
Jm3wrI7hDgAdR53twFRSOD4ZzflxUXXq0fELJnOUWIUp+Gh/JPKW+j5aleWkU+9Q
l9kOtt2GHXZIDGtjB6na9UlQdCq0GYr5JM+whryS13cnG7j17vaMnLFEUJFWwgMk
2zR6XqFK9RqCYSZi5hq4IBBM0LaSpFCoPZkiJe66pO5Hn5RdoaGWpQtxt0aEG9k8
ZI2LY412Czhh9juXh4m6qzgdgsEBGiBVNlgVio8tIlVI7AgP/o3MdAaeWma0oAuz
U4tP4RosoXg/Pe2WGXc3d/tKFK5dY9Ep34g4f08eRt45ICsSUt8YFf/3fyzg3AZ/
lzFbTDjCAcGmGzVLFHDwCzHhbiOkd5+STmR8RuAjxU4Zi/LOgefAVOqIAbJ7pxBK
/0WRxDuyWJb8Xr47J+yRs0Gf1nrlFzV/YQmH2fXaAMk90U/pOfoOisqAFa+ACgJ0
NKJIc8Smz97+r15upOmbTcdnker3CdGkDe0NYyk2jy66Jy8YWSKPML69yfy2TZ2i
O9f97LywZ/oM3Ym5oRJs0bColiQchTpvgczyjqLt/2eeOGq9WIdT3UauLgWG9tbN
sR7MNgX/JuDBfPD1cyjsz/Y2JizIhk8mxUpuqWxsRP4xlqcSK1Yw6C74qjS1NvT2
sSLlU3UWzF37zVQmT+a7C/n7hwMdg3WkP5V4JrVurfWOpqPbBEyHYX/tR8yJQNhg
t84KuHOtM6eA8sGULddHKSnD0QweJtFyq8dTakmSoxHPrGOmJKtzKYUoOhkfMRuM
wY2XK4w80zlfcYcgu9b8Avn/sMWbCXAy3iqOL07PjGtRzYOY86OZlgqPHpMR9NwL
Q7oSChOwrUApChQd4XuEEz2bgb33T6kPbN1UYxCIzzWBLPfV4Re4YTaeOoVmLxKB
j7DN8PnMRb/yaPrVCkGotKsKVy6CMt0ZMvtr+hXRq1cwuW5uAq39fbBExnGvhs21
ZJuCFhG/b9rdnYhBinW08hEWiYe+6DUBPSsMNXl2/XCb2aZdnRfsq3m1HSJa82dW
/z3c0eLT6zG1az3RX2AFz56yNvPadzx8QiHIczPmOf7QoUbuGplFe7OexVBbXa/b
ioY7h9MLXVq/c2TLgyCpnK3irpXl1MKkIRj1e9rMOCqAbBusmLUk0fSUSt7xoXnB
6kB+WttEd9Jm84xY21ZVNgGmcBRmwVfb12i6uDumZRj2LvLU09v/lbf5GSGwQ/6n
pj2Rv2XL/XlZlvLc+grFbqdFcclUbgUa3CQzCRNfMDgoc69Oah4jKnLQhk8o5TOn
kiwGPPPZhjdRPA62sXckUA4GgNKH2JEt4+AXiO93CCDpZJz/8gOzKWAVyevo6a1F
pTTZauwVbLA1V+Slsz6C+otzS44HnYluS3uqfE15FOVLPCLr+40ujMh4zXPma8DB
gxhN4owEcAFc7aa0Vev/1nfjxyu2EoAVHvHxUczSAftBaB4oUUkb6xeV7/q5CV9u
EiCvqO4I8xUVkBStroq4Zxbxab8A+j6rj6q7stKyedkACsuILhps3rD6YSZV10tQ
Jc8J3G71MPU/rWMMWKqopTRc5zUSFCrfIKPbEF/R2B/U0VvVk8y4AiWWGbcJUAYZ
wrmVMiTARZnmTMBthX9oaffCVwevD8j0ytxnWYuWzA4ExKC80YOX0tnQf+4Y4bHe
fUagtvg7nrGCvmBFxz4xaRf6UdPgCBDzRqWLhKY4Ls9ZY9EMkMatv54RdSocwYLk
Ii+vleDdyN1XlvAMXCgJ8cpyem0UJjXSnvZc5ixPefvzDK5yo1p/7uNLd+gtFLXh
qs9Ta37n0IHLZqUJY2c95viGKi5vRYF9pjZ1HH3kyINi/g9H3LgTRRgReKgCG/j9
baWQAqNUwXYUT+OJGwRpB1P1OvEyN6tspE34cZUWOrMncdtJwIaKGsBcpxz6BIVX
X4HMwm8yzQdBGUumAsnc9pMrv1V45TmkrQMS2qxR3RGWljcnhqzSxrphZuKS3UH0
vrCY+3BHGMkR5KmbF2L7dOEWERofZUd3VC1wLrti+a7zINVvUl07Y3p5XqARZsOl
91yc6dKop695cdsgZEzcreg2u3NZImb8XP1+5Qpcp5zeTqACH1yQ+mdNsWoq1ucF
PBf78+2WKMWL17GwNZ2CiIQEXmXVMic3k1Ko2tPzW8+Yr6dg91jdV8A8I93EgabQ
izxLcRYcgjzOC47PMtOssyBKlXjzK55xRpClBv/Yj2drBC61IIXaKx/i9Z4uLUDS
1U9W6mAh00EJW6hesOjsuoh/FA4z0xLzZpoOpvsxebFC8D9X6NPIre8Pd7Pq1mef
+av2sEPEVFBgB7zxNQ2lPG8rjhkp7YycchlOiOxttqYuaNJksGV8Eef66bBfg+D7
B6NZCCFlnkCrs9yTpwQabdH9H96qgtO1iQs6H6aW46Oz93rg9dEI7Wvaf5uF4jyL
SnIcBczTkHFcICx8fiaFeOHXjsHEJo3vu+SmbiVYu9LAxS6Nncf5Xd+TCqDT2aY9
nWQfdLE/SbEXAfZkkXoN+jgS6DCXemcfLuAmhGTvgIhlcD7YbvdDrdupGvQURi7a
+P7K+maixS+ViZklGLuM0OlozZxfR8zs4+cAm/H71jKo60nIiAZ6IU5vVCdAEf+2
WIl6r/gUyKrdbSRezgDGERjjzCJYAyJN5sr0Os9aSYOz708guEV7QW3cxpCMl/DR
mULPEPiNYLrOX+20ShfzmmBTrh1OboiLpd+kb9HNkE6mQHbE+KKvGOM8Ze1wbKug
6mp+wT/5lkI/x+CdHkJ4NTJ+C10xaDPOgIPuCfF4SZVU/tOPBPYPGTMv9/8OgWet
UOi1OamsBgPsa6t+jFEWGhAokckBWtd3TKYNclfkzNhAdB5HQZgdmrd8y7aAfltr
5LzixFULr/u2LYzfwEJEr22MhRNJu9QtZIyfgLEyd4qH7yJBTOFDD0B3JzeN91Lz
GnfZIvE3Xj/NP2ySYM1yS/ySQfATyBTkqTBcL8i+4zb6R69EXh/7pzzuySgqc4rG
iW5bNcukPGLkG3s1LouWF6Fu61OWcAfmInL0UoyhDsWLNfYUsYOBCzYApyt5tBPd
aOE6mR4o3dx73er0BxlODU1XYTkndupfuW9lVmRiUpKQ+AqVS5glSQ8LKUAsShGb
aXokB/oyScUm958M9J8I9xWqe3GOO5B5pDqXfLFN+7iv9f7i3iYUwxY0P/SZSYbL
PsltCQvCq4jDliLtK3OdY3Sv2uC/ormqrvseTm9x7LK44uMXB9hHboZurf4MOi/k
jmzDlgvH4uujS1fhUJ6zD8x4wAOrAFZxrTNiHjJT1dWT2e/LgXIYq4eMOiTzApeB
fXoecyN8iSuRe5FDSeyCFl7JNKV+nL9KvnS+gtXhOzUX99NmoXhgadidspPmSoyP
z9HB2yyS6+anSOvxXBByfgpsT8HjVeWEBpdHOelFn5R7ZtFNcCy30Ycum1Utvma3
fDm0QS7mls5EyPxPQuhApMjd7Sz6WJ7EwCZ7PaPym5XjrxrLA+uMGqCD+WP5jT+D
50f86aovfX7NNeEBW2FtBJdYD7yMoz8n3LPj6EJ6u7PqyOAauQjywlzMdZCd8tMe
pjqpY8v9P5IIoHUCQl1FbQHn59OGEzyy1UhRjYu9jenCrTpeJ8E5fUq0aDjFmjcT
GNzeGFlYGo/pooLwSwNRHU29bg0kHx4BQv7paCT4TX7aUXZoV41Jltt5ruNKFAcC
OG6lkPwYGdVwNTSHuTC+ZHy+mbjg0jVlgr0V5125l+6xnJucRY3DLsMV2SOfWswI
gV7dbagRDGOi4XlszmuNliT+SLTcBIAsRR7aGvexa2/kvo+WZwZzuI0Joe4w6btm
IzZ3Y/twwEtEwZtIYBZZzZbo8m7ubH5pGGqUbF2bG1VgEcrXYF6WRxtNOR7a3ZEi
Go24mW0A7LK/KR5BI2EIiXeYt580CfPsWe2AxQ9+O5R30audpxQSaaeF0Uez28RE
JMsOTwXmflHRlW2FJ1fqYqaMfPWFVsQ2JCfzl/hr41aZiyXfKNza+7pS4KObyvku
wbvVz36LYONJ4KLFDkNPI0Ev5FYPCbZxwnBHRccdUsrSv7LDhY1MlOJvM7nGhrQ3
dP28rdb4WBRa08U9DZgjUPNgcdPBabYDGSX4tdlqcIUkhBXgB62F1VCPavewUl1U
g5d6K9On+HqvzGVSNDb44KcmArt05VJCqYNhTTGDZ+Sy5VMoA86FWqcJWumNJ3On
vlxbYd57FEmNYqXl/u2ZYecgHOTWV0dfm+O4sPgTFCxT533u7WkWNTODeylhCWxw
HHsOJdQCGVKifyESSrflmBpC4oidJYJFnFLyl7HbrhknW/51At97tTWuOy0S14KC
gFwqSMkPTCeAgyShIqbVG5dw32z6OblaLPMx1Lv6qvv47aX4nPZbnjD4zPXrFT96
YK3puy/v9QOIPTJar1EFyScZ1eEDHrqCxrPScugA5AJSZWgSWrzyG+LVpDZSzz1D
rl2mgTsJNBlBciYEJOoXTY2y9xkHxALLlMcbZZIjvtXM4urEuOYWH3FJd/vmAPg1
9JxGrqWiUUB8ir31Zu6IK+FgAkr0hMSnZ3jU8LHNaF6u+vqRQ+kwKpkVfrOKAS8B
g5Bgkz6WrBJMBYooMmcw4hjpQnmXemnRPpY3vOTlJftpFJdZTHwTffU7jE3FcukI
s7c8GzyIdgGK1xD92d0VW0Ne0+jh+QptE/5LOBCvMRWTSCXiacU5Z2v6j16LZB6o
7+axbM6qmSZDGS8XUha7BiQOmAD/2pYndKimJWexH7dR7Lcuy2WxndYxR+QX5xzg
RRtek+nxBchJ78cGfZp1eC7twBGj1lJ/gOj0THxpeKG3zK09ddDfLNb8F+iiPFu4
PhePwyrd4SRzlbpMxioBRRebEZshz0J/vWt4aa3ynIHAig08AgRGB4TFgr8p1uJv
xTJld+0KrA20UzuabLedyVauaFiQ9haN1C4TPQgzvnX8m0ea9doX650rcoeuzvox
+sgfXrhMDB93wIUQl6cgruwNBoA4OGwHjmgbVjxS0zagwSrw/uu3gyzp5c6+1ro/
cnoGYo/M0M2K59V9Z4l5wQ6cK935PQtXGqVAgzNyPb1qU9p0d0rJLcxIZkcEKs7h
sCzWw2JHYuZooC8UsukKUr6ZczWexxqtwOmgpcNZ34+t4rdjvEoWjwQKTieXPPRV
b7d0fdPQegNtJXpmBBcGmuLD4gmNAF9ADHDyDbrkLF2coXh8gqswbYf+z5ybTBjp
770R+BTz/qB4y9VFA963i69RFbowHJV3wGOI/jeTxcfboqbWePd07KI2wWHe4OWl
HG56uVMMj6yO0fMvZk7kayjLEwRObwT7qQxxxY9zxYGFVx9EqiZ2RvS+YzXRGmAP
oZQ11sb82JWI8mEBRMSSGPCJhslyLhLzDCWOrM4EA7ed91JmcO77mACvNBmf2TBt
lPASsLzPISRD2+59wctgsxRojHWdaU/ryBj4WJW8djnWTMl9jwjHop9iXdbp5PmJ
2vTiqqoSko2G0SO57cQMdFC0rzEwsOAqOSdkrV4AqsdsWJAFc7CcJDj4Ql1X248F
kPiOwYhlkDCGKs0/ZhRQ4XlGPEjPktvNllpJl8F+R6W0kpD2X+NQ0W2H575wuWge
Z4MWzzOMALAURxq37rZgb419JdGGYSJFMx9eVH3hvTleCYIETPqyTFnEZDbongli
Pz2bQ+9Lmj7X5oZ75PZxbyZbA9RzyyucaO5AtsDdTsduRVFXLYFzT2KNSm8Q6snk
74JFS6Cy2EBFpkY9KVqMs/9RWh9A4k7G8BHZ9JYfXQIigNRtbAA+GCDiy0bkBeZl
+Q8m/11jyV3dFQ3apYYbIDxtKZZDFj7iUdzTihWNIsYk8xh/ju4es3hb9/YIrcGj
auqrioZ42Jpk34qDTIqI7xDmH7I49NVE+9bB2YwYaiGxHxEY3JN0n0OEHRdWy8af
1QEuseFmO+xn7PZvpGm1jRabk8QLBXlxRNRGmXxNtWd7s0JpXzejPLtfOrSIDfNi
kSaTF0xrtHYd8y1eMXwKuxPj+7Sbrg8qdiRrF2a/0zXthvnutAbiybdGQ5nWWy2i
A9W93+ZCvWwyw1Ejwy9UINq44EvIX7RTzb853UoFeJ3ClHA7S9ryJH9nW/10rcsf
hOkoiUxddV5BkBXs87I39HTCtZ0wYMYa/qX7N1P4kFyvJVGMM7nl0DhIf1+A3dtT
zbZN4EY9aJgaD4bLU0TZKkXouAUjyKI78Kbfej8mKJ8hc2jm0fBwWgmN/3iIzv5U
nfbM2HUKVQJ7qxMnrwBG3CEXAPNkb2QYkACPYSI0JqiXu/qq+Zp/CMaskdrqbOQ1
yBo8GuefnxhvWfbmeclSegsKoIh8HPQqvS/hY8jt8ClelmGFncoJEEyXGCDndEWX
E3KcDbfeiIv1m7Tg1dfeAfHv9DtAYP4HnkzYcBTGHP1eMS1X7FTy/OAllyJuSPN/
8X7XxvXSi0hHsmr0BBGMN+nvNkcRllBKd1ncHK1c3M51aK3edWGLVgknNx26I9Ot
72wpcy+Ge9ZYIJAXtIIpZ0X4Ihs8OH9geQoNdRrhzuW0VCW8hvW1UKfDFcHQMReb
xEqB8t9D40yFp0jKV6dGSqY3kv+dAraYPP2tpXu6pxGkgBDD0OZ6Io38Xax9DDQC
G6YhUxbaw2i6UbSfd5GIdVkjet7LtVrXX6vo2IH3pE2xwfAk65hhekCd31wTwPV2
KxIKFFBlvYw61aTBgg0LEBxqwYX6qBvm+4S/epgxGy1HtKqhuFRo2FB2Wko54jH1
jhIBFud+Pb2JRMc/EBQbDc68JxJ1yWnmULBNOR63Sj6KgplLc4JUh4c/HdewHjSC
i/lo38i3aekZY2s6Q+QzkUZR4a7HuwHV3W4AXktOWhJfZ6Uf0tWy7YfizjjysBZp
IP57g9UZZpl1n4795hBMyTiuFSzepN1sC8V5QNWAJnfhYp/ndNjJ6IEeDTsrRytl
8pUJuDSuVCB4KPgsryDtFDEXNy9REfQIUp6BjxD8f8NJdC09/08XVM5HBze/8eEK
NoNa/k9SaPd24hCCpI7UBXiCCjXa4N/xW+kBPQrckluOE/0vIABEdf4HILmzG9nK
0dVxV10PkN53mRxdHBqZfVNaCAdy3myDtElGJK0YNSoxUS6t3QAuUmcQ1u0TZd1n
XHyfd7o8ifij5A4m9Jiognl7VEv/LNo2+9ACRpDLEIa5BLmHtHEgCJQsBLFpO/yq
/Czsy89rltsbHMFMAx2OGlBe8yKzIoteScneycgSNUp4syN4UD0LAk9CU+Sh+Q6+
N7uGayJwWcBxLOVhApSLGAXMF8qLi5gaXM89hcbQGNDnW2EQGqg9kq5bH8bWBEsZ
A3+tVJvE0jmDm2A4ElzAHsE/16lYqM03HjqC6rDz5VxJxoMMPEk3mVmkxs/34yS+
P82O5D8awLEKo4a0oxMt1D8SKo1aZidhQy5X7bMPFlbdYEKlXA6YO7qDJWw93j3c
Qa6f6a0d+OJPhThkZFvjdVPtYkrCOpvy/V5/9YsyGEF02B4t2QuUYXdFytxX7x7T
NhhxYrobu7c+VSKID1sdJC9MRT+vhsw8bU6yQUyHXmqZ/0QlLYC6gELkIMAOAi4+
KBN3cIJrU/uG0+zqLqZTOMT+J/NoFaD0DN0eThjjv7VQrP07lkyd/hvpyz4/SbpU
V5NYXbnQawo8K52T9KO8rANoJZ+axLPOivZzQ4l/l9nR3ElV6ygo7gzfW52T6jT6
+Oqjvn6+vpLpVPm4gnkDLH4sE/pGw6VbcCbIr3DSAUJ0V3i9wbxeFADoFO8wRl4k
zFznemAV+K+PfyuZ0pMLgmHOpPrO93NOTD1Pdu2dsceSZNmotSO1vRTtoFbXBl2w
T0xVzC94Ksj9f7LsETrJcM1tpIrkk8rxBfNNpgYavlny3vqqBzKAHwhWFSI7MJF2
LiKicEdXesZH9MDV827jAQrJGptAUJTwminTy8y2a5CyidmDv62xROgdzhqdfLca
gE2gRwPEZ9XA2JmAeG/PDNc4BEiwfPa1Y+6vSFabfiHlz5vkOnp/T7e4LlfTC6rT
NcYkpkyKu7fAgNDDxbkZYGqocBhxWZs0etoLwc+SgDh90eXPz5C665FXKpYZmo4O
vujI6laOyArvk7qmBOv/yqzTed560zCjrUl++gTm6bSiQhyP2U2lfL/QI0132M0K
XU2rHnvDMBDeGfF6QUCM966d+koOAl1Z7ffNzgX951oNs+Mh4fRQ84J1R5EV9/9p
hlk1iwgAe+Zz0W6O0ueDKzjqoGM5WY/sA2x98oplcZmbcITZD80Exm6MYXPtAzUF
t8Jdk7L2uUnnTWj549dVkSVsOcYd3x5D1Vf60lsQP0QdrIQ8lRYQMjq3lfkEeXtr
Aaoxj1pc8bOHgrjpN0Qg/HXcEDJIMTKLcaMtV9LmWQsFLRXQfAA1sRGVPGrrHZnt
vtHhbdU+3yZ8xXyLQIA1N/DLLIpurR5TywfdQ8o7RVuT0TvyyO6mShDjD/Tdb/01
fhhsxCnYg4qQe9fhNI/tSysx70iuTZv0tQ3UBcIfyfN0FwVTFI8lBFhuEh4YcLu4
02KZ+4Wjnhr/mF+HrhviszgbCpsUAHA95jsWlCJEaiExqVcPTreTkZ3h4hdA6/Gs
d2Qbat27HyZhyi3SK7BCyYNS+/5B6TjShcKhizaiL32PdLiDkSnrUNF7+Cwd5k/2
VB1/5N6DD6u+fCsJD9fsk5t/jlNRmpXJx1Js3U0tK7Peu+9AFCjB28oXjEt6K0yq
rI/dhCPN7vQ9zThVRZwQR377BiG5I/6Bu4k5H2may31iVQdRlzO+3gGQacfVWgHj
+wQk6xKZA0G7iEIdesdxPwnKAHNvA/ZFKLz4TO4iCQd7ZrZ96ZJ/Td2VEHvu6GsE
RiWYKeoZ8wq/kOwqWzmlj7G1ADPSA71HAbZVVx22retn/f1B2FCyHAwgWsf7GQ4A
0n3aD2dg+apel0xIRhFeXKHABX2aTo9y/xUYHBmEtKUjCnRfAdnLIZIyQvhPEcSo
FstnrB7zhJtLhmVjYEXTeEAn0zbI8hrQIMQu3i54MrWK9om3KBaQ5DG3K3tG64wt
8aZNMIMuVCIGsxmHma3LdUTQ7swx8kZ53o+ipQxE2gnFDaoFYRFwcVyv/czx002b
dcJMxiEY7rS+L0khSQkAQAzfB3KPfbllgJoXY9s1ob1Aus3eUePU81mydH5utlql
3NpONnccp2YAeU8h42piwwDdYotQhhwkxWfHO2YvuGiUzHiAJ2ltPC/3VQVFuJCm
az3SoZHGHExKZyENkdG74f4NxumQ5sn7jBXAPmWJJsO20ed035QbTFHzeX2e0RgL
4hyKKnF9sNOCnf2EMwMSasWf9r5gjnp58tTL6U7R+C3pseYBleJ0lFPNfSbuIeXm
pAa5U4ZLz+Veomloiqxv1pQ2qvJ2wvZZfiuZ4iY9ItTD4JXPx2ROtyfDNm6AtoHs
HLye5hyu58n/SmWZquSNV6JQqoETiVapIWnRmwN5YHD7UVT3ptWG4fwzwJdbsWXW
LPeLxIlU0FtYnQknEmxWoGqD4er8uTnmUydMYMLDKhdWE6cZULfRQCnmAftXp1Mw
81JgFukU/MXmWT68MxRLvaqu/TYzu5+e1vhcNvSCeUk8Fhask+OJHllLTq4wPAWV
G19GW8iSJLOC1f65Z6zIYBHMqWEzbvuFKH4vLmPP8GkAsFvB0mf6R6mwfpHN/mAb
vdLq9CTgjgRYbu6UjPU7xOebZjNdYyrQfq6uhpVqCn7HDOIu4kO/VYRJbMMWPJKb
stCQD87IkxlEucOdMeagPfmaPiiDBuD682Y9RiLWpSR6vg4hEskFnki0ltEITmQH
Kg3dWp8X1ZQzXvrXij+cO6srOhTiZPJW0DaDprdPaQIVFmwRIu9s2SUB8bO5JXAd
YrU8rdLRTbty+W3T87oIOFBDvPPqdafSKOfgNXrgUCWoQ336bAgAr3kbzptfI/kc
8RSK5sfoMt7KgCgkDrOZVc1ZhqoAdbLYcMRe9LT+yPbwAvQ+jy3TfOyi/oLtPPiV
5x2vFlPix/qhvzBsv2atKu8t1NyEUO2YXpFWkMDfU5g+tBV+PXZR9EB3Kzlf2mtk
fb4xVmzRrkLrGqGgUBHHFoT+RfVfpWUzLPPeyLHc0wkRcv9VigC8kw0aIanpF92Q
U7XyiB2k0PbMVdg1pmIjxtKNcZlTaMs6hS9fch/m4jeB+RvVgVv5zPa6Xd1REnPo
3/YZBWbfVLpBtxzo/pWmkCNOZM6KQuTcEtUh/FQ3pzsYaL6ryVhXhgPLMCS1xNWL
K9KsEkVwteJumOGx/7lD6WP5RAb5qE8PxqGQAXCne2xgd5gmyCHTma5i5YnrRUZO
2INDdGtDQoqZuoAlOd3g7uQ0kXgKzk7oNzBXIa2hhN9V0nrxlNGN70J5E/vhwQtt
y0vdYN96ESSi0IOkodTsYkneddXnQxrWjPDtkM6uljp1kQft3yCQH5b1SW4oXLQK
Vqge9X4g10mYF0zOhRuwfBQuZVOvYBwNnJ1HzlxVHbaKxPM3+nj4EPV6kUEiDYWE
6IMiAKrWXwIeIZ6o6CcW9tPzhFWj3nprzmj8CBpZjzjeXmvc4BVeucHQ/hrx9XAc
s/xNfrnkC6Du+roXigPrG7GTXgy80ctblguMkTPtFs0ttH0VdT3VnvlDLiSwq8o1
SQKG4vzEESEK94i+JvC2gKFEn8VvX4vg1alzTyXs5w8EFRc5xLvCtqbTITH06lFX
ZCRFAVtua6Ae8xhiWepKS5QYScGZdtVThdbO3fGlbNtbj7RJ/MbZFwZtNdx9EmMM
bTUT3MWz/ejqHznk9YlY0Sm/qmTUZqlwl3Q/ZRk05E3bUXSD2rUfSAExkUsRAIv3
G7kLGU8A00yutTspDOhg/XtxTpdrrTi7887hN2pYz5Py6zsy21Id2iCiS2HoGn8R
yZj/GylvV/5iTrhpvenuXcQx1hLajGsom+juTX1xA0yIMy40nP4K4N3lyBuc7emB
Cnre/+4AmIbAOSolsnU0UUrkSW0ZTbcjW7hbuaFP9waSXeuCPP5HPErsWSrroTat
DGfwMwIRQ3UBY6j/uA3iJ+p7M4EGqfbXWe3VyYhdM2baxYixzqkPaTuHSaJxetS5
0ddKscVsqh4RfIHuDN09LqRj7PHqvPy1hM5hlIDkuUl3r19uW87vkJHOzsvKTjpI
YKLZVvaFJeM7LTbCvH4TPwHwEg5OdcxxLnz6KxGiDkm/Nja2u8bqkFE5Z7M8XX4U
RbKA8PEckt3TV+oMO1ADOxcwPR5BXg5+T8680etuxeW7PuwUtnBt3J9RMb7PobJp
8hUyBF1zrvoYBNvYEJGeIA9zSUFhX+HKi/+lisCxBiSDzJpQHNW4z0Ged1ducP5o
LqepqVILebEa+VTFkDTaaLavHpwPPWpPb6KT9jk2CJ+ikoz5AqKtS8QHTbrbzJb2
tYnjBF9CLKMRecSL1vhWaRAVYc8Ewev31k2wQTA2bPov1uOg79fg5502IwQiixPM
tYYAVUBhqDWzvZ0+lcTsjl7OHxa1M7yz9pGULvAW7hlHaW1BBbvq9D1bke7QPGvG
ZDnNvhtbGHw5XrPQ3ZrU6C80HcUBQY75rBnEAKcxi4UbMpR43Hi7CmqxlkPyL/d3
zqic81bmOoqSLU4Xai6FVOKHT2GEqh8d4zaJ3DbyCeQN95dtQcr5zL5A4c+8/Znh
W/YGU2G0s4cr0hqeLke5+OSpWf6Y79uWolnaSx6D1hVNKDRLcgtV0o+LC0NWET0O
0XdZYYluFsBqBvlxIcR63hENw4rdBECq23GDa9XsIbsMV5aCd7NNOnhKBh7otxwb
NzyyxKQpg27rsRqy/2zcjx/H/XY46IX2EGE++j4qvpFNKmOyuETpB5VXSu+sHzOr
Uu2eaoz/1b1PqE9mAz0SoO9FYOw5E2oz7Nv/x6EHUn2NoGqtJSNYmt1pHPMhA3ZI
3g0rNkb0BIPgAQg2nG6ICwYcTJXCfVItS+1Vet4UdAn+NF40WGNQN2ff5JoIoy7M
KF9fGgfC9sw84iiWCXH9X48ObmzOY2cf/vGeElO+sLyN07yI+nQKOuVtGC/8QkUf
AqhsFZw6vhAjY+uNQDqm8uKY4k7XRhmdwEzQQ7KgCggq0Jwqm7WOVpX6GfsLRnbk
Qx2+EqeAWmATNOh2JKqAkBVldR1YpJ7/UxI0U2FouYSetJy11T9FIgGG+Dsa1DhH
kwAh+gAFnNww31qtzYBK3wFBA4OZwOna5Gvoh/sTfsg+yKOEa2xkYDBUlgDL4Wut
40HB8LryyRl4xpGc56me2lTUoTUd2bhEYZwdPNd9orA+piM8lxqGHloHD+d9/cTb
gS4vIVraSxnBBDO257vtf5yd6NrUitlQRM69HevRoTW6RizhzwOrLqDdUTOYh9g0
kLSGPnSDVPwIP9lrTR4ljondzXEfUuzodtTXhHUUvxE40i1+y1VYUwRtm8wwIzYN
cNataXKZSlIKIEfO5QWaDJpTKuGvVMR2H+gaR5XZUpf2oe0ufZeVeJeZ9incUMyQ
gX6GHgLkSXRRyun7RwCJyP5mzDl+gGReypTrKN+Yh++qR0KLIS/QZBUn46RsLz+Q
32awC6IO1lepICaLezX3UZauB1oyAcAzCZCoi8olxj/qADdjYtrrWrmjvExGNvpj
Yy8nbc0RQSTaHcyVUCZm5Jgk4QKYiWeHzbPnRxr9k5jZot1NlymTStM2LEZ4DEwc
clWA+FWPErnosbEuNrb+oJ/TNYk1ILfo+dJ28RZq9klGxMcCjF6/gvnLY+S2SWB7
RbwKMx6ez6qjNgIiK0F8Q6lNKGKJxNLb1i3jugI5wnTsvMCdHbwveoW09TNwc/DW
GtPe3dROnycI5jLX8+tsoIduQlBQ89Fr47kYup1Ad+w8oFNuvSKV0f2Zc++SjpH0
GjMf59xej1XsnwpAKwRJcSbwqB0M8mE9lkXsoegdtPOt+y9gPI8tjExUCMW9vqtk
PdjAdWoZSGHf79dajDyTD/u0of4ydVz0yAzRH+TzpF3Q8883OH58Jq5H6mBZ+cQu
wBwd6mvmiGSEJCcUFvRGZv5F+PIEjdu4AhTQCTBtxhR7t01taos2J0kBH/pAalz8
xCcUceB20tORznIfNGGA+11OiS2lSHruz2PiDdAsfVYtTDLnMJ8zbVKbfqEKWCbo
8p5TO2RMpiPZVVCFQ9B0W23TiZhFUe5ll9WknxMomTtNE290mcWTNvWnqRiXGKHV
jaPHOmWEdNO6zLLiicSVz3je2dcfdj4hev/6/sFKyln5hJkhJzJZEE1Q0U2Zh0sk
FFU7z1H9ADjdXO/xKAoiBDh59ei3ED4vXsubLSFys2ACosBGhPDFrOWuJmCtIST8
6ekyBniOdYD2/PJcCRV+atpnOOioODW6jYm0p6SNR5mxeUFvck8gegHL3JgIGLgx
g4oUQX467OlqlGcXejlLXShBlb/gv/5a8Om6G2daiA9aAy1cfGTX9rBMxvvswZ63
MGMUdcDegl3GrTOOfMyDKAGmDZy5khqGnI5fU/hLEvogKueJBiHQrDCDjZ8SEHI0
hrzUH1C3jIK56d6NbWLePapXRQNsC5PLLoikeaZNHtcaU6gKOjD+RW6NTlAlknmo
/Nio3ofwrBhoSNlmhQ0rCLrM4qA0zRzeBCsRuMBoRCDO1i9MuGxMVD1Nt1RpIH5Z
CWCPrG9AdMmb+a7sY6ZmFka8jkIOfN68xphmziuyQzNuyrOcWIXNVOmjn50uB8U5
7VTHQloF8ewS4TtLK5InBQn0KvlgHJtXdsKKwP6YpzNCtAsZDWHYjodPVcnEtXyO
utlgJFIxtfFT73ru6Unpwzwl6SvEtlyMZ0+sRUu9/k45Yh9qSscFunbW0B2LVTUb
Mj+4e1ezaYZPOZVMXsHt3oWBABQ6FHC4I6VQtHS3Z6P/sMoDAtxaAf0PJI+nyud4
RbCqarar93iXJfoMDSy8/JYOAIklp8O1apKMEmXpmqvgaRBtTSPjGljxKdF3wbAo
ffrq0m9hXBAAfZRH2L+Kz7oZ1g7loq9r7rA6Tn0UiO9xx0mdlslPPpfYu0kap5AT
fYiDxTkgCXZvevqhgW5Orvn801St/uBZJcLKiQK+0wFseCVW8fWag98EecbQ0blj
mCHOIny5Iz9k+t0V5fZb9T4gG4XO+kgw+n8yZP3a2MhBBCxgrGIv7vkvJrJ5DY13
s8CDBMEojiCnSDUFC6R0e7vRe2J8DkWA8VEgw1YIz1bQWVgkaJbj4tWEg6wWwvYO
U5rHY4RBn222YfU/HFCfvvJVuDI28b9suwClS519fjU0Xbo8WSH1wNHyqP4QNn5C
UTQtH28LKlxWEa3fDqzeLgjuBn4sckS6Jx8MZlx1qFf4yI7de4fPHP+iDn1tKE3c
kStMO0oxPLhV0R/caaLoNX+RsF3YfcmQ+kKjnGvdAWtyZvv7TXijxw811ACg8+k2
fG0XbxDYzHPl+U7qrUvobaj1V2Lj9mdXEqkKv/bX5gBT8BGVw7ptzyw255ad00LA
+ZKCQ58vcsC1M1qD3tW7c6xco0LhWglwLpUdpF6r7hxnUMjcmZKP0mZPWTczLImV
LtavFtat68wLlCqB/ICr/xGlbksXBIS97zUD6Zu7ywo+1yULdeR+HWvsaAPtyEF1
V92juo1mUwkWdkgtJXmRPHYYE4f6Eq9xxpMnywNkrWA7erRxn8SzFF/d52wrQI7d
FBUFWUin2S9FtotFOhvNFA7C8D3ZdGUwh6ytigF9xZ5U/+ovrV7XOMMVoOnWmaY3
p+usvg/W/C+3BerihLBy4sHlCqfbIlIFP3nstuRsiqLcJzhpXqrn4y6SRIAc8yhh
dZOKN2sFutkkH3V3Oe//Cl4gxm+w0bf9vr+/hz4vuJzv5zucJObioy9M3NY3TH+9
ZYaRvomLK5Yoc8DrfjPMoiaFQCsXnWKgNJfNYW2kGzit82MehwpsFMZJszvIBPEh
3YmJx1umzs/1vPRCq+nur2Heats6dZnqtrgtk5wvtwlvJTR2dQTNJWfj805V1+ay
u+mihdahc7bVitj44oPRyH8euOdq5BWxd3J1NUhVQBF/aseF47kGFFidBU7IvFIv
dPgzWwn0veFB+unMnoeXZrnrbrRkM91HgTQ8ShbumyNhuA4U/O1eOeeG6mVuwxd+
quckLoc6yY64p0LrvMakO6+5U95dnGTTXVmOn8awc2COWiT6huq2g/YxzqnKAf2e
NhCkUC9+Qfy36J5N4t6VwHV+pDLuKfIDYKOii0lZTnGyj/dg8b+SQmkK6g9+pk8z
dYQniASMilAgVzJnDDG2db716HH4VYkFs3iHuygu2xUF9oLH+6S0ASbfSgIuEkz0
s3ntRvpHpFfZJ7G5diYGjk91xyq0R3q1M78k47FkPRh/enUMxkt6w7APwmb+CcGj
NSG1romQ/flzKqkt8r+65xAgexFlgCU1p7ngycfA7a7Np51d+z4Xas6va5tTpZHj
rMlTH6fg+1Hj7qTAfcshEJNT2e6zoMUOnHqdF/FWAh3yTL//jN4ExpJAFxJqbK5n
bXHidzM741C7dlapuYONHTL3wEBHmuLxcVZnaHCVuSRSvLndLKklPnehxb5Bt6yE
vOVMic0D49FPcXG2LPEBQprEvnU8qyFaDsV15m3jR7VdfdiuscfYczpycPAf449G
rsv2/p5m0hKRvbtHiiErXm98yXyOqjH7CMG+t6KYLXv74uQQqMEEMiwmoeuk8uFi
Ke/uHd+lnjo292DI0XT/We6MNlV5FO+9gvs/fV35W8xD3jZeP8Augghp/ekiXfBo
vh4widbxuStOAaTbfX5ESIaE8I9qBuTl3J1UO69bqS1PHRpgu71Zp8JGvkydhJKH
hwNlYPyrhZdwYcPNDahKc6dSFK0p05B/tLzHVbuAqO76Los4Ev+xF2zgb+czwrCy
yH7m1kPtzwkmC/Z+nh+gKvisjt85jAW/jemRoud2ykXRCdvv65lmcRSxZAI7ZSyf
Fql3lqG0o8w0XvrHFiQQd5jdMA8MLwiiRdvpl25PJ4IMOqEMMwp0i1kIelMzzJf7
Se1gQpYCSuQzOODzg7wdRkR4u1590v2JIgIbEhoQwXfmt+7lN4bcWf0mASuCqb0y
Eyl3DM3H+KGNihLYnw/UqbqRKl4kvB75yvdeJfhn9x+fCDKceoztGNkZ73r9MiFk
plbOjBKChj8Wg4jho5Ibda8Y8pMoYtAJxfzIq3Gtx3GAxY2awG6oAsHbVK7g0Sz5
xpoZH5/UrfFcr/H40NE9Md/LbICUjHoGd/vuKrLVx4JzoAmg4mhVyMzO73uK/4DX
GDPKgFbhFvTRrq1G7BYcMFaJsNeCFzbaFVowLkIzmGKl8PulYJh/2LZavOIYx3Om
Ny3wo01nz13DBo/ZUKq8KwgYRbwLJMIMwL7OW6GC1Tc/tredUX9E/MkO6AU7sQ6h
N9F/bgvN1LzBdoZUddqyXF/R8Mt2W8Atog13mSETRoPgmToD3bfc9t/O2LhYNtSC
obfQO7nESeB7pWiF7cTmBQWHX9wPPn5ZDJfmWozacoCXSSFQD2L95TTBYEXCGQPA
vxx3EF7PPHdCbnqchGH3K25ziC57w0vjdEFjWnkJCb2BwwgyPMudY/LR0veUPZJx
uzJ1+DdFDa41fVKyAfcPUrjx0SwUdbiK2Fo+/U6fxq3amZHBjkZVCzy2j6gkQ+58
Y9d7aG+FYm/jgh1HIw/hKMGHg/mmeSwGPSnk902lAJR4nI2APg6zUSabuOzEIMA5
MgF3AGKjpqWtrbhn+qsNSUJJiZ6CMAJ4JUGDAb4hyOWUl85lQBSibaOKZ0dz/3Hn
uIMhbyqYbDxMAEZMZXeLmrFPZ+5JygqRMQckM3QUvXYOfiCy4pE7a7azek/K/Xbv
wVnVZdbjN9VNZ+xr6yhimpzaPpmz0Yj4ffsXt/UWQC3MefxndebDQP21aJEbF7oK
BY33Dp0bsx17DbVUvDNo5gUxlNt4OfgFGaIw7X5uQO1k8Noj1OImzXn3Si7rLqfe
kqtfLwLWNn6+exeZUuvS5/9ROdk6ZxMEo+RiotnCX1uMJ14iZSMh1S2pms+J3UYV
LWHtHscoF4IH8ZBL5zuhBD46g7NCAEcxn0KOWBQ5Z0fW/wnOkab6gbaReTi600vJ
kxRgy+K4JIBfM+Ps+0eYHBcGhESD857NI7W0bK3uTvcKIcWnanN/K7ay8woFZb5S
YrnCyXNxSDaHl6IMn3l6WeCKccY4U/2ZAPSpdFpPxcOH3rbEFua9JcOwUeRPm4gc
n9T4IxXbi1fMgFXnr4rzedfh4QNzPD7ExRaBFwiUJcjYeqBHb7HK7Hg7jnRYFVnp
BYvJhVQ/8xuw9yrR+b2IyE1X3x5ULFLSVHT4pG1uI/LhV81A0E5am+c51p8AsNJn
024dRgOqDy0pYqsURLf7ZeovF/+mzxM5egPWaSVMl0XZdPqcD0owQw+R3GKPRN7J
CbkV4X6RVfWd2Al06mCQeVSeSVjHcfI2NMFUTWELwPKtkZEg7yMX1tYh3LuD4UIW
3+M6lZqLo42N3ga7II9diw65B8vF12g/2ivoWTCMUk0iHcQiWGEdY2y+sh62uDG8
5gxJbPQ1gfcAE1ZoedmoUdgQEaQJsbZBLpNXOk8nEq1pVQPMFF/yMaX/7Y6Dhhqq
6Alw9KkG5you/IMFV9X88bOFRF6K0F6f0XThuy81AbT0pleb2vi16/Mbpt/4Y876
t96K4j7wemvXl99rY7Be+QIi6Jd9LAGmJXYk3iw+bMYbPuCnOvuRaXXwk9/p4NlF
+9Lo6ET9cosU51N+BYuwgW//X3mmfJi3gF/X7AH+CjpbJfTwJAFJv/0hqgNLMEJQ
4bZtu/tpPMTXmJgXAarYL/oBFHtQZuAxqILQW1W5QUyWhk6xQSCqJTkTJbxrrST5
afCe5lJgdfD9y6IdV0vTevSXwgyRVZN0YeWcLYC8tASFtcyt5DdCL7WvC/UnWdH8
yz6lyylPHmg5PSc3rl6b+m1MsJdctkhTR9awMJBUwPLDEJwISd4OAc8ytvkFsfcq
wnDiKS2idXydpKfBTtfC0SxHjJXpMrNV25plrmYY+NR204a2Em2wl4Vjh0mjbA3I
6+ZPbtS8Mhrh+6ZglfzybPQziDUvaEtFb6HWxZKscS0gyV0RI0UTpR/thWqFGOtg
Oyl1pVAX293qMPOk73+jn4cgOzBC5LE1lFic4wcuIiIMHx9ZSb2ND6+sssYCJuA4
VNnnzB4yhw1BooZIYR4ujExfxRLO0PbOXOFxJQVF+TYUP1SDK851Tou97Z1cfp54
xwkSsza4O78bEYQIWCyU3Vwk0Z8lO3jPfXsl5lRAo80yJtoOTbH5u8rkGTt0slpz
5Uj3cp2MALUU/DILj2RXAgI5s8MhdwbWQg/hJ8swU3Lr3vqylX0QdQA6gYJQyDjc
/l2aJxV0tateZs0paQorLV9t9APprzLPLXEnX5PUVOc+/ahMh6it1zkajDrB4mTy
Dl5+rmI18kuRlb/9Gw839uKr2XBuM/8Y451cXOJtjACcSF1e2bNXUDn6CYp3XlKN
A+KAuiy9XyMrnR2glEAIXNYAwEYVwiQTaAAi58AjYnyP2CZ+ixDwvA73MWNJZvyf
KySJ2w86c2r165kyFszl1q5pF/pMeol7c/+y8e0sII1dPGCGWVmGQgG0QiOtatUX
g0g8H5CWdG7qeDb7BPrTAkQbO9uUsk66W3aLlffvMdrh11fyPikjjG0tfmpFjGPp
HzqCDnw7Bapx9Dw70nHRLfjM1BT9/25N+P08qugeQNBvIPawToKtHM+FR/zzH6WE
1Ij0iTNb8ACwf5GByTdWbWOK5ztBMVGLw5EsbF5Cjn7ZjqHrdRGzYrzjXvYMPSCY
UBp8hCl1jirhEY5GcGQ0NfDYY5gGDfMVdrXKedYgFmmgt22UOM9e0Z13L6D9Klpo
oEwj8lxcwOgUFWOlCWCgg1gjmSjA7Z0X6BqssDnpOO0ZGabdfoszr0BOidJsgxcg
z9ZO1hT4l5DJYTwuWFx+H7s8XQlnHNAvBMajVy2E2uTz7chbWGdqxbDalBySsGy+
50vCjRv1+1VBg49gPrKsX7RNcnsdqDy26iF94VRTE42ImliBvfx/BbhGzzva5DUQ
572yLRViCk7KKruZy/47238CGTlU+9NOMvOPTT5GFvAdr/YWGdBNNJAIzFpM3d9/
/SrzgMU1XDqFy8KcCiipaPw6dTV5148OkaknPrMgohXzMIZUhnRpzglqHFQ4nuPq
htj0IPK7u116hXjlIRtAt/3xdAloVnkz7XsTpDGBShA+w3MXMLggb1aVfdIlfceW
RYF1lXvO+f/Qaumbov9AQ2QDcrSUxO6oNCVjToT9JbqJFLqAjAKUAage+z5gZnAl
tqMFCOAYcbDdgyJxJOAELefKe8MYwNEPgDXkiIulzq9T7umHAmi0wnHyFL46Nt6/
9Var36huXynUOFYLW6tQD/iBAVLw2xvm7tXl4TVi6f2/IMj8giO9g7paSiaupuwo
edVFkwKsddvBn09xR1Y31Zg6CH+Ihytr/Ek7gC7RU8DHtRfUxWeGQmedKx6XLTqK
Tfsq2fdAwFZMVZSByjh3CaEsqDCaj36h5ok9Vip6kNnY+9/bzv960FrYwkP+OnNH
YvdvBKzt1eBsU1X/Px8OI/PV2aayuIzlmXhQgbfN0IekRvqPXtRz+xKrJpko6ptK
00pUmKWhhI+9K/fMzCzlLlZ/y7ZaxrQTL7Gid6104w3+xTWJyHN3B4ScB5Aund/a
hWleugvHFzYBQ+PqB5gdjBmkXwI9A3WKSEXPd7DnoeqZ2Sk8XQJ36YzBx5MuOKFF
WlraFgGfRRxWcNLHAt6z4mkx96kRBninPRnOIFBhIBIrU2Pp1KSdV/OinacY6tDr
ZIfD8TOqHeOWvWyQ00qwbrbnBWpswy5RfAZXExaFnyzmVmSwDd/1wHKZDLMa0kgI
K0Ry9zBwKT0kyWqx9M5Sg37MeEBUMH2GJwAnQTNO1CFskBNiHP2SGxZsSYRzPuKv
qKKO+FGfI4NVw0ElimoI7DAbiaA3ae6xwMRueKoKy61VQd7pwTDJJFZnUDKjBDkb
+99d7Y9ajvhCg4gedOrkk9aNq/vgq650k/3brxGS/GnFWtqDtMwEq74kXncgX5BA
teEy3ftSt58JwsacZVLp3AGsormtKip4Df+d6+iptL5DCQSKs4z1EaynsMbKL/sD
78nylPtpsbmhY0Zoe/xpy31LLmJ+sQr/r7N/im5ITjKwkzWvMtlwhrkNfaMoeaJs
RUZmtAReshliJlUu0EjzBEva/nR6KJGL6Wfl58+YIGTWeCx9kHiCnAxb0OUnX3xb
vDNjCFquidFDnJ4RaaCEshb4FBGb/pr6dzH+csV4xZAH60uiol55Ve/VkcDxt6y6
iV7feiGxtkc0d1DtVdKJSf6iPeSckHNz0U/vQvAnX+GhLoCotmesof17iryeA4WQ
wipum6p/Tg8UktKqfeFiGpAbxSQhevs2SJiQddVa2qo7jj3LKJdy2FlT6G5t+jwW
E6CrO9CKF/1Y7gPbHvlRtnzgz9Q4v95SBJuJOkZcTwPNFnU+2BMs+u5vsuvsk8ev
PHL6UDKSDW/ro0/2y5B25nMBG/5lmtqhwpFLllwg/kbaFiLshARNOodPzK5RAC0K
r0Oje+xXSz6vUb8SS22WCv18s+LgJXMDmJ8X3CWkkovZBttd9aHqHCU+jJV9LC1/
RJ7jTrj0QwOFxa07VirqW5uVND7hTdvQLAhZLOHAT0CcX+cFWRd7wEOBR36fjQ7F
mX86kgx/hBmBqVkZNaRGCbO4uM6vffqfD5u8ktXhO8NvhosCcVkqXZMWyHD9hnWy
QDn692Hxyo1dP9nsqwZRrit0kypkMlELZKD9eRZhRCWyLXYOuRnkAnwm0iVVu9jR
T2ZowA9jFsDYSV5MJMxSPuyVMd1dDy1Aj/uzLxvnd2i8HQRxWx+kzYUbtv+qPaAf
JJi0QiAjvZSg3pem7rZ2ELc3k8rwPX9VcwgmACf+CBE17LVViEapww+BpWrpqywt
l0l+gFtDzo87t5UDfq9pVC2eT7gRnKiNJbM8WaNDyBmtSDWnwpC6tu4ltVQs2JVT
ehGNTF/oZwQhV94BGySQVbw3mKlf+CF3lulEHQ4mnItMNGYVBYFmSVRAM90fvt/a
kncqNllaFGUa+tWOTkDkRnfdDZ8aBpASZwIlt9rd18Re2okY7uDwznqiBoUUn/OB
+GEdk1yV5lTwcR46guqUsFmmJkvf0PkQrRVQf1mqwMLLiQ0x9AFd1sFEvSRK911j
90NCUesWXVAnJrXfQ/u0A9qGY+Sr67JQsYN2wzGVAWCLruv/fmN5S4+U7KHM28YL
mBxPd6hZjd+CmzsAtzA8S8Z9VHmPv5fJFCanSbKoT1fYvMWpajvZ1lBR1jvn6TaS
V4zzojr4QeOQK3F8St5UOPA0X8yTsuBUmM1w73uk8oaCfmwdZzlr3s0pm3GkZ5UD
G3Ws9Nz6YZShM0UY6a1S137ipoj2JeoeBJBn7fAK0GCtbHm1gXfGxdVkCUf8UqLf
YcV9ozrqcEEG0U4PENQiUlpgLrGTfi1Zg6eFxohwAS9Lr5Xp2mK8ueUmQ+yxP3Oz
6M0JuvZyEXqs2tBkvP4C/LE3STP0IEjoHoHggrNOrsP4gmBJwdc1Ry2AmhAGD/+s
AFicTupQ9g7pabXV3Smtodol7RQM43mzrWWTVLHCjdQXCFKn3rn4SMXPj12LN62Q
PM0gGoPmuQK44O8j6uuM1tlqTL8VA8FoGclOkF40EmOKGNimWjq2pwzsSujxRQOK
/7hLHCgUFUvJc562x7kmuYYG9/WHNsyLWbVN7nH83UwASz9Z4o7e2m/nGzbXAk4/
Q6Eyro2T6j7cffKsEY9KbPWz+noNkeHF4p96t9laSJ+1WuQI0KsyjZxc2/SQBBKT
dEfRuuDCaX/HDAGoNyFywzuolX7Itq5f0Csr5bCPzMDINome51c+fyQUGf6pTZr3
zSEvomVcMwm3RFoSxj9N0tIMzC1j/EqXal7GECga2GsTjE6vNHo/E02q/I+V8fex
mQyWkzd+cXMAujvypdgE6vKIeb4eRyAl0dlAho9KcMh7rb7cAHiz+M5NOh77zVkE
GN0FlJOAWJREOfUXGXuJExx9Z+aKrjFCuGQ3Gt17kdNeTyaPZ8RBIhqrWW9Hi+Oz
fdBwr0xV7XMNbZ+IIT4r/tipV+SUSSwQYjxnORFHgWsoActF820oDt5/2OePUQ5u
h/BOUn/Cjf6XzXbHeiTDX1wNEJQx74HDJeyRbW0Om0xzWK2JmvqAPQ2zY1EyNnAv
XbahFc9BuvZKiysTZbI5BPmX5ue11OKMqSRQ/4ae6zJwC270IWebO5dDSpcQVmBd
E94g0h/GbFzVO6YkDONA6nX59E1dMLDwXz52GwLR/41TGfHoAZou5kIl2taRPHZB
kfCsCASKRlNmfbvJFe42YClPblkCUGknhPUVOb0mKqOJ90/USzofU5J4/f62yCDH
VmVpQIJsJa+mJM1XYirAN2ka/gYkio94TsRrkWGOb1dWStNlNH3QwJX9L65jaKAV
9C/YAHhXSpJlf1Uy9rSnwJ4kDJyiyK/hoL0Vz3R21MEodx7aEoZMLBy05imp8RyW
/x5F0KvlchEw/R7G/sKWbP1EJps1Q5Dp1S5lbMjUCCTljyZrWkBJBqTrDojoJxTA
mhfJcb/mrvaLmCxYN8JYYB52nD+k0HuHP+O18wMk91j57UIfhot5cSFQYn3fzP0F
VkTrxGKgFpmghQ3X6O9CBqyujGNldg3ey++MJiCaazWFJNGfGOFVLKrdhGhZ+JHY
GiER8MXfv2OYU/9dm3Mqw6irQ4TBEmOfo/v9YPG0RlFxYysy/6G8uSfQVOnReJQz
uwCczriQ1oUXHf+i8psiGpKx1lBL/v5x2ebbTGa8qeGeIyAD/WSZhiJQaJtAaSMp
Y2DiCHIcLQjG1OnPSgQS759voNDpMetoyDE99Bj3BV72RvHal1+l6vCjAFJUEOzD
M2OTwhe3LDYnk3pVvmlgcJ4onYH6JC4iH68YCi3koBpPT3PgobRalaF/LzLswr3l
VMV4IIlm8ZooJ2ZZ0WbA1WNL9WugCL0PHlB+pQ9eYB2w2tIFaUBOGk/hgCo/7rcn
iVH1aQwf8bHtzQfYzhsGsoUDUyNZ7KAX6Q4XdMQdcvyfBoJdj/nrBvR8oC8hkVcy
AFHy0X6QKXiW+qePo9hLrHmjWgNGO27tu5CL/1vVS9PkHLFTaqb8pGvEtZZUhcwz
A6btcQ0tKnIfvqGRO5KjS4WPPyWRyhnD4pQyuKrJrJKOKw7g0MHvcwgmZwk5XFhR
VEFVasBqzjUDUv+VZPVeVaPZZVL0tcCckAN+qqg78lXnXUQwrS72hLQ4MsCXA9yj
73uul/NizYZv/SHqW87e4jo4fYxZ73/cCgQOmVkgKtu1kNf5VW75QR7Pq4nk8bpt
m11I/wF6zbs7AX5ZhMwKOPyu5QvL1LmWiQ4sA0y3IF2xlGhB9FhdEY16zpPDdmEM
5980jLaIWjW5wh6RxLKBwCub/2cqS/QzmKQ6qaYXGjUP7kvbhdm6FHZ8qy0YfLAK
hXbKNzjduqTr4W/hGz663TbpsifsfFi83gZd7jeit/vfC3pFeLRlvAr4nYcSt//N
xUhybU2IYNDNzYZEUqnGB3FGBTHtgBIT9CslR+VrQYC51WADVQy0TnE2R5H13zkh
T1z8BjzsT6OaJqpC4IuyWZ+arVXdZpUH4j7dvUq4rgUlT9oX+LuStPbDbJ7rZpZm
dOgZhghjSopodRxaQzuJmOHLdb1J6QJv903Gswyt9DZTxyREcWLE6Rilg9UiElvw
3ApdP3Ja1HXeI54m8zzwKXEiaNLnrigmhqpUs4zGUJEQ8mBvIpMCP/NcU2BtjY9V
GGL9M+LDSEcoc/n/KldTNuJJwPVJojkzuqecILZqGJR8zoMWoP+Zzhcf9w9/fZhc
36+JqpfDfm5oBx6cyLcKN8EsnYlc9/wXID/rBTjy++YrcHEK1kLXPWS0ssFctiFx
DT+FLZLZ65JD9RZBb/k1k8c9j6tNPxiz1RCvMtAuKo1m6Sr9uJmxclGHTU5vrcap
Z78j6Hn4k7Fz7L7lEzUbWzrBSzuoXkzAAXUYALWk5iOZbpNNpNwCsnUxytl+gUh/
eQenXbYBWo193EU8PVVRs7IOJRHvUcdFkeZqgg/5tR3GTu++DJPPMHDqvh1K2ny4
sD9BhmOvePqjdWSx4MOQE/ruiZp33KwAL+1r7vq7h9Hne+nW2zUQaJxjLWLdSgs+
shCX4kl3EcRLJpRIRmgxi4WwQ6ixezBlCEFcQVQf9/rGtIBkkDYaJX7DlVdhMVjM
d4AzdLuC2dx5Q4w3DA1DUQcBRVaFCkYBik4+h+YuEg0UQsh6yoNwhwIlyD/X87IF
KyhmXpXOy/ll6fcq1xzQcEQz3QZXT+zeWy+Tyd4vFvqPhYCWtgTr+R1c0hzAR3Mv
LSjsA57dDtQU7WR5aOCIz3dDI1AcSjh9dK00PCh8NHyp6OtPSYB+9TeG/JhxvkqZ
A6k2O34vIl0lIRzoU9lDFrVKp/UOkrjs3OjXP1McjjahaHoHBFG4zK0lx2GquyNO
KUgWTlgjmkJG39erlBr/71rewmE0GFkDDZUEcRHc1WDK/wLkD1BxiF5YSutlsiA7
5kFj9bJaZ+UcZN9ePcyf6TkMFGJFAhgfxq0JKO/PC3lVFuRHOqOFF2SRrb7hZZpf
Y/gS1IiL78/ZYqVy4w/Vgvl/9eLq9n+WmL9VBDdotPRc0IcqV/8oROfYeFxPRgwM
qDDETmSWIXYEm7mOKkd1Q05gaOfbH+jPjBD4Zg3Y4Ihs5a//aaXndHRdB2mnaIwt
tXoa+VK1lbTq3EZPwhKVsYd5g3BRIy0ipweIG2pCGcXsVtfuQpuX/I7wE99kbE1G
rWoOh0vFc9ve1m/PvKC6/2gtp/oQMGzhqDCH/Hx3ukHrYBToXIapt9QzQCl9L49b
cu8kbQ+4rVwxBPPWZB2rZkLBPysqqg5Duart9i81o9qu631RWeVyWFxwpRLKsWm9
s+60LdC+KCn78IkDGf4ghXaQQsyyOIApBPIDiXe5qBCAG/pIG9+dGq3HuBrYMbW/
DcWH9jbGGq1/0NF+pjeMs1l6EQuHqiJ2XqjRZUuLxTpwDfgpPRwgyHaxLlty5oJC
bQnry/ZrQk3lZzJi7yXMf/K9ISCDUGEemiauxGzQyJEWc57PAflAHxxbI9yv6nlL
SgbRnmEjQBJTLviOovAm3M5sFucbaF7W2/Nb4JZfbHY7vluowvFiCgZR3u+l0hGl
9cua2kSakWYIXcd04mrHggUmYtL71XMuiGCUgGq/1QB8JrmXynXxJzUTpOZKepse
knkQsfTKGRsgdYxCGCc8teX6tiInE9+kFwE+GWGx4JndcyZ5QEZmyCPjVVg18C9R
rpN/fVZfPL6dCoFKtDhEv601pDLU+J+phKiOZT2TwiZ9lgR+Muvd94mIcwA8Xq+e
cGT9XqWCoLbn+oSF2HC7tQWhAh+2YIlUrPt08DhpMhxaU7kaBnNuTeaMvTgESQHS
yBI5iosRugN7CHdt9f/5wB+MmOx/FsZ31sd22Kko29JRFsPtrHY7XTDUMLMBX1RA
sr3b3cBWJz/+i/bRn4Bxlcm9R7nrGIr58MG9ndLPs7sJNr/KC8Pco7UKXYZr7At7
EArsybnPJOmawH6bGjS42rWQKOAADJjMkpzt1gVZsGoNXZjXjrpHIVsbPXT/ZuOS
zc5dUVcUEOQB5q6d2gfHsnI42pQ8nNJq/dnFckd5nEv5OUgX1LbFQNJ+tJGt2fQ8
9p7C7yR+aXE647H8Dm8ZXmmmzrQPi1PK8LOVes3aaMOHrRF8jEobgzt5A4VxrUxs
UvFMKWq8ePz0NKm4Tbp6iuUYbj2riSJOUJDEkI90zVYwjFlAws37bwEq5aSs+k6b
LDyqfIbBXg8Lq+B2huJ6/JJPyJMd6wZPc5C54fwTrj5BpQYNjGSqhZ/jSsg4kR0U
2DwfvUzWqJh+kXQbGH/i8G86ixvqw3XYnEabkri+94Nr/r5CsDyFzymIj67dEMLe
0g7vYHHezqxNswFYFsjgtn5WF9PPGyOYt58Aj1zVt64QJJqjvCrk08KQY5ZK7qRv
IDO4JMvHOJ4ps3qEXX0mWbcgVvh9QN4uh8jPbi0ZKQ87ufkzfLD00OnFhfjeRqFS
fqO5QSD8PEOuGPnPVaDqZ56RGigAI4TAOh8VeknlYbjAVXV5GLe4zgf98FJ6L2Ky
j31E+JFUE314wnE8UU7R2eOA1gWqB8NQTj0QXRsVI88+JBMmx192sFptOoQNTTvi
q0kOd26iYGz+HNFaZtIowON9g95AWgBPGVu317+OHnDwH9S+17aLHgITEugDkc6B
DTvx32wToAEjHIjKPxXAxCNTB5fLSDnb39t+Hwg+l1ovY2eA0P4Tcr/hh/DwG+WZ
hd4ijEntuAOWGs2YwPpLnMBUlpfngqTGrdONgdfycZtNnH/bQp4mYZUWhQuTyc+o
2nwXtMGCzsWG6ygY+oEUg+cB1L6U2liZMi5fRvvN3C7iwKQ/WkY5bEgmwz0ZYGZF
WiZrjao37Je8CnsaN6tpleW6aYEDBXgwDhzFS4EKiHj2jE7VYXtV/mqgYl8kAtre
XWQfl7uvdE0eEsOtDBXTxzJiH/nvZ1us7vbzouTEE/KvH64BEDxDfp8wULF3WzGi
Ea9BHXMdWII5i0sqtsJLUzvhBQoySjSjbU7ZwtQp7rXO7N6sQZgidVUmmReazdXz
YlYIBs5e05jEwx6Mbmhhuef7TFrXi3N0VjAdMcviT2zq4GSvh1ZlGf3XVXmZnN+/
Ep+w4Qy+atjn5/TjQo/LZH8yPTiiXpsMufK/877FAiUX+nJMRoo0yv+AUueQswWq
wYPvd5GkkGTJKpXH1Sho0QT6pvmybGVVs72qJ+CQ6ylk2jucgjpUJiukuw+GjE+v
GoBtzRMrBssp/2szzr9k90XSt4saQAvMi50ztzxFDpJ2kWoGif04h71nC/L0NY2z
iBN8buzb6FzCii2g62swk5RsTndIAksOL5mn2pEbs7VR4Qp9OBG7xmFKfxEmkBse
EJKr07cpNZQgoxGJE7raDqTmsI8GB90uzAeLiFi4JGFqA0kiivbrNLjmDNMhzUOE
/+Jr3bGNtaD9ELBHMgShaAEP4qxk1kY7EIsBw7JFe+g=
`pragma protect end_protected
