// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jQV8lQ3/jRUGWA/x2u2DhL/zMKWg7y3Zp5itt572EHfAXfTcLh+wT49IDqLyMdXp
DqPvR37jxRqRNfNOMmt7VvqRJXW3UZQrxeRt+yOMp/7OLdT2ichTP+M6tKe9LjsV
X6yIfKd14LJR7I15ADJZBoai5qIlrJDp9eJtX/LaNkk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4000)
6TjfcGOVhLbmy8/Zt7TrR7ur0Pfv/4Vx3ZmyKnQHoGx2JFXPNq1GBQT1Q7VNWxIb
fUhzvraUHCsY3Afr2up0k95ktMytkJfBI+XjS3vaL48JfoO721R7FfZjHZT2Q2tZ
8WSZR+z+BKCoEJsm13yCgsrpQaquSmC2tDY4+EiQytQsMyAw/zMbqQxa8HCdZf0R
bB1cBkQb49oWEzhQaO8hQPp59irG1F4YUkT49f5C0L8CRqY7uVunpHSG/ay7M9Ax
p+Y2gIOUHOG3hrNjDgKCRY32uVDi15L3a/Eop+ukfX2FRMq98rGPoZknnhLhJMn+
sXlrs8TpgR5zqIqfWNilfZp9D1N+U8XzTZLkHXXXx2LgS9dyMTBhDb3JAdnCzVil
/V7wu5mXDMPB/rQvyEwR2WvY1z2lYzJbSkZbOx+dQ5pmn2jm1pajVRDFCOYOxoja
1BrhWOuQyUI7uXWF4q5kvjR09QTXKXlzTqFbnl2N3eQ+l3VoJJvn10695KdiOLPw
HCRgJg7lJte7BmwqSjqYlZaes4nD6qgY87k5uMHfvAjUAA92xHiPxoFMKRRZwNbs
C3AK6qemkFO0RvdeyEc0ROa5ECyrKP7Hg7vcNwnC2RNi97xcmLsNHasa9iXDzREW
MwR0PaSiJ9CN/yH0G17SJJyGLu4esirgLIqIe3Vv2KaBIVcqXQlWIBKJUnocbOAd
pVT04o+UGS/vE4BGj9sJ5hv+McMv3T96zu3dhqbdxifdcpX7F7GMOibgo84nIscR
D65gewEd3simEnJW/3n2x89xDpD26/SN2DUVpbxNabCpVyB2k6JW89KYmHb5U+oG
QmtciOj7GGwkJugwjFxvaHXhDT4iUsRoFMkbHUvs0O/X1jTLW7008AE0FwIGMyKB
DgWPLyHeNujdoxkT/e47aBnO8izz84vJDLgZEtELrwABQw560+cUQ0wD3rpnw1KE
W4JnZ60FO1mHmQ0FSdLZFP3z8M6UxfZqiI9TPxCuOb0q3jt8e1O1yE0B1E4ITCwn
UHdNwDKoVV18ynjJM46k5XAymTXDqquZYf//6V57oS5KOWKLMrqG92EuNmUx37ir
ZREq/94nbz4FrPmAX7CAYTyoPksfN/w9NlS4tGh4ZPuX0xsffYpjSnEIIpYF3vV9
1Tzhyfk67+5sCABqdVBJ0Pp+W/jApbKIEfTf8KL8n5XnF8vcYxrYA3buPLmMVXOX
XB9MpX6p64rBUcyFmoF7Jo7s3qhVP2WOZW63g9lPMEhmoYScwg5vOXO9BxzACC3L
/CX7dkCluOE1sw5ZLTvjMGwhGkqi1SfZmsfKjrKlWyfmxTGjRUoaUjXgBnotlIZc
bO/ZC75HM2FODoeyfbdxZrxnJjr6H5iyeDrpYtYe8H4dA2GfUL4q2Bg8CMdAuqz3
04pS1KkKbTj7KNKnNRTmVMlSAEyKLsyngNUfVg9pzBW+bppaJax8qeObA/MdTkUE
lXdqt/d3A7WgFYlT+v5Gfp5+3bw/GisTAIkLM8fTke/5B+5A+8q/XQPYonDI9UeN
F0P6imRVIYG7y2ZhXpBHz51ogL4Jwe1IeXCOV8e2w/rvmLiFnnPP6y+q/+Mpvi+5
hmpVHF0XdXRgwAQAeeumXNA0BYlALlX2qtIqpcjC463536tqUqtjpfnhqe/ZFa9Q
ZegKu9JddHOX2hjasjZBhaa/GzHm78NZni3lrupd1ZrO9rlis/9RaQAGaWnhfqvc
ELxkMgmAxL895gJqFk2+jh6z06aOZPsfVTBNzwkud2gsV1vDPXPJ+0GWY/6BKEWw
GcmrzhSsskFkZatA4cLll0R43bqmZZVxSXYFLcmptAnIpWizIdqZ6Gak1Z7hRJtG
u1RB0vXDaxCXV73/RCXkts1hEtXqPZT1b2zo69up6K5uapb1MJkxMn4z/lQV1jwF
tcUy4nm286yOgTF/BrBEZ8zVamc5KNRUWNFwSQcnIp+u6fOIerHmtQXeJYHWPY5j
5v1YofGj1/YJso7lDqLF9VehdDuGInWB8q/XM3T6LMT6Carf+fMPgy3hJdjA9RER
Qs0GzoQZ6eSH7TteAKQuk/xoOWGyzdfoH5ZIvhirKknZGLiniCg4Y+xglPLhVSQk
QZs1iAkr00ZBIY4hwZ3yFJ4dhtLOnP/+qZllQto9Ib7+PdfXo+kcC5zaN3c59LXS
9sFrxzydcmdnHQCq6VAloconrAOXUGEsVuvzv+Opbo8Pc23eh8LrgszXeU8HaQrI
HnHvilF87kq7HnltLsIfgoYbfQTKCkeVKYnizIV04/uP2sajZ3RFd0xZq4ZJVNNK
sTHoc4dJRSHoaMaWoGHtvZzRajpQwppkjl1fDxlGPncli4cWsYO2mLMIRfCOrx2Q
CMcazHNdGlF3fs8KRCwO7dl+9CAw9//O/vggGzuUpmKWkWahBxt2vsbS2eglBkrY
RrnpzP4a5n5rVNc97CqJefYpqXmHcc47CnPd78m1N/6I90DuLJLpwirjGO6KpcdY
qWKn82aMFwBWx4wh1iOnX7UZfuirLHy39wwXeRy+zGWWwSaHB+kBFcQ0TbAmCv6T
tGj20w69Sb8XUSpfkdEPMzZrce/8seFScjKw76X/yiS3AMj0eQbY93bS+IRFzB+f
7Z8VJ2LfHGq/d6F+bZNLk7F/4cdhBUyEONDQPdEz2AbeUEOLuan3NhpGnDzUgJ6B
FU4GB3BCzEjbs5dWTcgcDoOzVA2hKfIzcw4/Xwi4Vs+8K0ZkgNJNCd2VhFfJxsJC
X4hHbuRyF6ElHEy50iircWw4AISDuu8gAW1xOqoBC0Nwu01T7H/XaAG7UeR+Dv/o
xMFgigi8WC3zf8ZkaRHAvoxseGXCI9VkFxXTbYDKqqOxGmHZjYPEOPq/vWcXS+kZ
RM9NXjWVZ0ZIKZQuVDyq2d+7bWj1kbDeFuV3olFJi/8M3BvPg618icnc9DFf0U0x
UAksBfoASKecdPPc5nTHypTjfPO2hEcs6GIe1+4EZbaTytQ0SliOYYzEZNxSx5ff
ioPDAe9ePDf5ihU/gzJz5wL3sTeZBcXVR3+hIVIYI4IBVele2rt0tcdXtJ0F7vL+
3LiqvjrERvth07saclO4f63sJWU7ukwYfVnUhNVYXddfraTkUj0eB4WM3ZEqN1z9
pJ+EUeLQ1n46b5bx0BMMiobSNG2y3bzJPrKhafEOsaIw+rpmWA00x7G8uqQOiUXW
+1FLe+z28IVa3VnlIOTErXwnAlCH6fxiJDXJqRAQ5a4BaNTqPngf/K41KCwRAXwZ
GABioSd/qGMj+FHI9fRJcl5PxYjBQufLlLMFxmpsqco4EpFjZ9Qkaf6NE3X3dOqb
n9NoIWJKP49YNYbO+elNpGKW1uwujzp+xrjme8M++CkfdPYdPfjVrDP0DM0zsZ3O
Cbn5mkqk+Y2PsvXHQRdO8YxTnmJYhtOmfkz3ahxG2h6qdjsBA5PG8tk2UI3fooS/
G0A3LzC0bsMzfHSIdYqC4Z7wHIOswMfecPk452hcK9ND34J3vj01Aks4bSIov+3S
Dol53/x7CzSfuUUGgpa8z/l41D1+t/6niiEabiAfRVnEpuwCHJNPk1+aGSNAbjib
JmLXKOPLo+gfdG32wZ96yNQujb8pKN+n1xCmgouc9eIe5FM1PKESfHUJJ0h3emU0
My/YduTn1YD1jRJOuwRSDkIk4L4/02rp19Rd3jTOttR7mcqCwXw551DTyBFlbNek
myaOcwREhyqge6/rdqTcCRugTCYnO0rvOeLTIXqsBTfAmLm7SCFtka/7cRosTHOU
556zPYtZ0FweIR83dKMhLiWWBGAVMXWN7rzDXWdVABo8ukC8n/IVskoEqzOhQAs3
8uvClUEoSCRzeZjcnu6U1Zb8q0N2Y9zkVVEUTJXniDTeLnN8VRCpr3aXqdoznvF2
nQ/vS60bv7/1tml5TFzRhrNXLus4MlT2/5JXMLBESsRyr6Sjs+MmUoI20z7YQsPq
6CUdB3ZB1VcSjgzRXVDSMSPiAvjDc6mGQWYcDWG8YsUauqxhlVPDcaX2JLcfQxCz
DRKjoXPqhmYoVwAgZWkOqyP8dgWLuzHj2skqlvFkVY63JjlCv/Ushw8TV264UJ6H
aXtfOI1uc9HjYWKR0KdnKeJi+RWpvcJs2gzHays3DCmHoE7JZ9mOrcwplSTgF3g/
8T8oa/O6EY+TyWP23I3kEnyrjLlYN5FgFeSixrPjAJ/7mhPgGfpFLiTCvTAWv/sO
0rFYVTCxPNqrV1y4JMipbolE6taFMzbgJPn5O+SsdE8iR8z1wkxR997yesaXAXyn
Xlyqh9KtbCvB03rCoVUHMlJOl+os+C47N2UJHyQQoJ3ujhE1V1859Z+apZMxMu10
OuGT2VtDqX6FowY8Mz7v6Utauj0jhLqIDDZJqp2HHt1lpKVf4dXTqUSf1FyBGL5h
Eq6C3VX8XBqdydNRRITjmOvpsr/N5J617sJ/COn9YYxgY+p+laVqbWNBPa2+ZqgM
+YMQrDFrKjxhD/Sn/RICiv9CvwlT3D7dytUW51/DqMN0LPTJTZWOGpq5aVp0yJXL
fWpSf3zckVsBfZTR0AahDOetOlOuL9Iuv+6rdLwesbGabhYksMqB0eUJYoV3Vith
LiEifzD32iiM1scmm/GKhsfiCHjiOWrGUgRXiYoqsvlA501OMRMXsj9YlqDNTsR1
h6SwGDUZmBnvSGQVyi6f1H0vjuCBaTm+Sb5jIx9WI4tLNSqfqOvnmBDSiW13SzbG
tQQV2TlLJliYwTC6oGf4BKASUGlTLEyjk1sIQJ+TcSE6KVC/HnGH/PJTIVKCryq1
eiF9sAtNuQnG4Mkzu29pyUphbWZqx2eGsFOWMoOxxlgNeJr5CLPrgxO6jZ8UU7AG
UzPe4EWU2w7kyu7Hch1Q61AVDDrSddW/gzd5LEWFKgeBbPjAyH5hpuOCWlebG1yq
lWdL5rE97IImcrF0HlXrSUAhV8BrS6iM91ZSrzanUfBUymi2sdd8wdWwjGg6ff7F
65wlZy17vImu+zRJ4bZQoT0SD10u86lYvHsTn409//owHsvrpP/sLtdALuPe9VRT
/hv7sFUti/m802R13BL9bndc25/yXWjjwbmLwo7mLdDOobN7dgPy4fZPUpNrIEQE
FUMgfWOAXWUcXTmmFfyLIbV8xbHt64jJLy30vzMTk5STjpitKFdYRAFvbl4DmxJE
n8mvn4fDWVapyVFUd5U2qVxfRd5HrZ3K1HzWsc211DCB45SE192JDMSdiKUg2l1g
1X7MQv+jBcRFNWYdq3bTC6izX9jwm8HcKtAe9tP882B0WuNigO5+EaxmoLuRGYY+
baX+slZt/ZNgTPsEFbbv4g==
`pragma protect end_protected
