// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AabeTgVPwXAr4qjWlrSiq44574Oxtrp1NKr6STgyw6tRB8voFwbWClyFOBOw+p4E
+c/lVbM9kzEC8IA0MM1/eRmYwsLu8ji6kPt6HDQhcM8bwaFyXy01IHpHO40IQpAN
NmnNQ52cK0x2Jkci9r264V6b/hr8JS2t4BBM6eSjpIs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26688)
UUZLa+2fyTcmWYs5OKjn4/V23FQU1gznImFpVrqn9aAkDDoIdHDuNWHU4HUZN6KW
JYXYAI3avxgW05wWBYA+WDem9uDFEWT0K31eveCRX/U4QWkbrW60Ba7gh1Zye+NX
XH9thqvapzziiZ6K2549+Hf5mfOg0cBnAtvUpm7ERBw9+CLXyL2ND5C3e+kIFc8b
Bo5LZG4QcyY1yjXSEJSWxzeWx+E+TM/J+DihM7kRsfqLYetG3eEtmH5IUJv+Qqps
gZ44HJoyg03wKv6TEa6Ou/XBZ+znI9NuQ3Qh9z7z/CCJ/w17WvCyjYorp8WrDLgR
4uHDst3Ok+lnjQjCyEjBTIxyCLz21298m5KGK0c4/zdR8/Tf4VFya5ss9ytcDiPa
sitBubdRMHJhwnfV7VE+GFDmCrTjxOIROzokQRMiUsTyFAJXmORh8O27/k0bpxMj
HY3SQ1tXTZ82k0KvnAzpTmeZFzA5ifW67mk0e8awix3+HdVu21acRdAzpE5GzdfK
4xj6N3oXpJfPt0YJsNInGy2WNo/0WLv7YMm4YtTmyinZVjIDywutmaGcRWAkxZqR
qKPDg1N0KyKFgyh1jmxya2FpNODGejSmvySP2xwgcQawNoj4lExZ8Sdgpk7HziEI
saj0YhmIIoF1H1aSPP39aiuqb+xpwG+Xd7TNNSdk8ueW/draj4QpnqNt9ath6OmE
cRcvDWPyPcWymbpGrJmcMKNy5gDT94uiBN/SadF+2LRy0u/N9IzJgLhWHwU6/Lj+
S5Y1IpWgR/VBDA1irdZ7IMpdiYqa94RXw8uhfvFU20589h7fgQCyFpsAKGpy/J1j
xZ4tDXeRh6TgucbnQxQJKcCwy+u7t/w0tm5/9Jum0GQUiMUrSPOufSFMC3KnbQ5n
Ft9ycPeyUzNKw19sktuns4E0xM7s5zezMlGQQt3m+WsVUdKTJsMYzSIUn2sP9J7+
Rf/+ZcC8jC/vOURyZmB7te9EvrvOKNLKiPppGgKg6P6no0kjTJhQYJv9lpXpuX3V
NeFh7Q820XS8ltWxRqY+Sz5FLXKEq4BFrurwVbVx9Vbg2XWZL0Nouv4T5tFpyVVx
xu1KCoHhi6b+KmETUip9qCdqIOY4adOd0FjSdjGfK64OiEjo7UOU5FnI51LcAItx
uhCwBWLn0s11uHQdpHIRRDb19pPcydz+DR++/n5ZDyhCcJK0jX9QD8Tx1Yi+bcxv
VI8xLNciYHb4pQtoCyg1FQ6oUVsIZU1LOzj270AC/+fKvtCw35F1AkKYVL6S9dcW
JUgO87y1Fl1nym6TwEgkUrLYIKkxlHqjoBr6hCBRuo/DL7m5WE+XyBSIYAANTErS
JJSfqD1gNc6C95Zeq5LlCM/x6yBluTEZl9+jJ0lZQUVEbVN90JUXqX6/egh7iAaR
SfJlftcNBLk7KC3N3U+tWJG1vTfRJ18dmgDOpiiJexEXRn6cBoQ7a14fBWMK2KTL
DNHXaDPkoXXXbYmNJthnq5ZmZ3ZB68lRELaaUwS43G9J+b1a5i0LJJLBwUb6twwr
EAmWVUThIo2vHgv7tg1BtWMltkfEReX2fZNU/QDHgMCFw4XnQ7PrrPy0f38s8tZ1
/0bUe0kQ/YwtHU0zXCs6POUXm90C8modm0PSUYZRQzha7f861bmGkrLUDgWo7CEP
FzrmMBywF5rIgxn6erO8wyfAqpe3aib3ZZ7j4lEPaoJikNxd0fv83wu/TI5nOSnv
TgUL2SO+g6gCamzr8jVNjBo1r5vgnNbnQ78uH9CQO107JGkJgOotOH8SBg2RfSFn
8+co+vgTXXeWezffyRaq6zD4HmAFAU4dycICVULVQ6xN+PeIEHh7EYi8jOhiB6d8
7/oTndmMvQKgFZd2pbbunlISECEmx/jKFLjjtdb+LA7mTO5IshJKoBXwgz33qRSB
whQd6lyYv63sgS2coyc++VV1ebb2frg5TJpLxGldvT5fp55zkcz4qGz39D0iRa9g
LhjpWnmZ8ojBlaL01/iu/KCC49i13d6awzFXLYk6ICn8vb2XWeU9/iqy99Xy/vg9
qRmEM2AsqBGONbn3JcmumaQWSDqbXQMMfcsM3ALa1HvUoTtVZviUDVMYaj7iIfcK
0RpvfQKXfzEpDeGWpJYLbv6vfyucenuW91MIFpisHhPt7JNTLTZiymS60d11HJj8
R4dBvwXYZ0QcdfQqdCqQkYvQycWwaReuFOT5vjD3Pu6D+j7dUqEFTMLf/XMABpba
FOkZGOXFKs5AbNGMLmJI3M7xH8JbHdHA1EA7dS4Szx5gx+SBONXgHjccQbADQ4jR
Zjdy0f/W9NJ6r0nH512Mv2VPyci1AgN8DxE0KXWGjET6ZlRGGYmb5hPiX+wSscG4
dVzJC/pZdkt6ElO4eu1C3OqL9fsp5ow7waFedqza9bKFwdWNg1ELAak77bbkWaIO
gES/tQ1HvCKt699TmPGDiQfD/zqjOX4pqBXIKgbkW7GBHW05hNNg7IlBF/D1Ktoa
xKvJWssDsFX5XxyQ/w55JNqLa1M0ADq2e6EUqQCmnwehlXK6GdzEQnyz9fTPH9Ru
ysEn95diEajQiGAHciUN8yuRxyI8Uov3Y2rPW7UsYraLJ2X+tsFUoIlsY4g9RcYT
uelqqIPH+vtwq4bc4zjJTq7mlaA5CAIiysOgkVChraLfF85/8QnwN73IYWUSp2CS
VOTUoX9+GzjHC1acGZ9jHOVOWkUQ3h00aCn2EepTdtyc9t92S7E8afRAQU0UVcpO
lrOj/3ieMqaGI1UgJNMdcHq/O0VOBY8TGhSnQ35r7qjmGGL6fW4D9Mqxj1sw2adu
J3p1zhvSIq17rov2w1TNRggJ1gv3/qfuXvWxcGr5BTVIzFKVKObMIfM+bqItf8EN
KeFsSwFAtxTh5+3auK0EBUmuwMgo67/FSlHGzx98zxY2s/JJA6F8fjEXHEZ7GAOo
Ee8kve0P2yywwU5wlQRLHJUd3v8W1sBtJSjFT/RiNqg6fN4QjI6bBUAxdqJ4HGP1
zpFT75OhT2eYC3oB/ebfut57vKCr+kOiU0TzGRumB0o/APPw3AzxV2N9hzVSXEQF
W5XrlAVxw2rNm0oNR793a0fYBh4mkhonlZFW5oQru6X4nhApYWLGXz08bFz2wgbJ
I6x+ne5jmrQ8a98/c6z1DT2XYaNOMwtshCDC6qjSlhK5ONCSQTTX8x/66XJNHfGr
6KioXWhAHOUGQC2DKmIzC7fi1gLUvfQeETlBhahmoNd/K6cWODl9Rn0qJ6SMz6Hv
Nf9iaiTE+S0+TampFAQbmq6TvT+cZzh0YlE4aeNECB5Qqy4sobc/mgUogtDjDoWH
0wJEdn7t00Bqr19jv0bo58TkqLijV2PuySFShnUKatMqUN1Jgr2WICQ6jYRPfis3
3KmuBgEQC//L9ice7QfhwAQ3YiYlqiB5vhXeHlrFw9DSb48meBZ38zduzFNgoDXw
cjPhpbxaqCRsFZxqyl2WZFMVfopOOFgf4xQeXoFjS6QGnAtmkQto3fN4KiJAtRGO
UTwGcJ6wQBDhCsVkK4zoCOcVd3hxUOuWK5+EXOT46CSNMJUqGrbJ33xPnyxvZMAZ
j1ZIs+SOhnzEV8XRC+9D6dypPEX/RxXPCa2wyIN1ziXuW/Qg08CTq17JglDBIlNt
8bblGNJd99QsIshIJaGfvxozJXDU8REIaYkZQJn1+kU4hM69wHHiOcLEoHXuGpfw
eSl1GkCnLBmA5cKaD8fOlcD7NVfOVMAoFXyQFgRy9ti2nTDseS7a+Bevaeh4mxoO
VhPnsZ7/yjf1nvK09a3hotWHTIJWg4NH0HkdO6RPOGjuEwaGVI/RrgMCNNECnSn+
4HV29KxV4uAIZtpPw+9MM5+P5drF7190SeGjfiiKIyu90JDc8z234w05St3M3NmO
oEFZaaJ207Rb7VccghxM0WUwAh5MJ7H/R7qsORk4na7DqUNobl1t0oS4sh9izgK0
hx0FSKFz9yGOGjABbesLUgUfA9Z3PhLHzsf/LEzEajhOsUengRDopMVSm1Fh8xne
HGUlt7SaCyYJEm7xCcYXyBojXaTqGa7+cg1nFVLsB7xbdiBa2MBiMiT+BCjxgXCO
Cum/BJL0YUOALHJfAanusr771Q3POcWIqdO17wFYLLWcXNxUMsMz1zaYKSKOKl0b
UROdrWufPjABlNBtj0HuxjWaqjGWillyPuFXqnQRp5ysV4iBSkvsHe7VAYJbY77f
5rHUIE25as4NNGeF/XrmSjLSf4tY344je5ftYsAODPf+lpBDPETJ+vD+sWvRYX6n
Hb3SjGeTnOD9LWW+YyQW+BLz6K19Z+aPITzrTx2rYywsusiF6TQT3OFP1eAnBVAR
Y+UNImEZbmQoYK/L6rvnXWGa51r/xw5k0JzYOYUEYD3HmXS9BAsdQwOm09RDDake
ERWkBZ+kytyhucOHijswDCOc2oXQdHro9tnhWpFd6InXrzfB3nS+qN+KIJ/yl7hW
Wp2sXhJNlX4a9oH1QW62As9B6X4YTbk4++wqJu4fDeVfup3z/3/vbbNW1olnlYdV
lp2onJLVaGucabjLx/Xbe02us3gZ+hn/aDnk2xp/RprHDszlQpsZa3oyOhadWKvI
Z4NU7Aq1LYfAuuM4UK+qKQAJ2q23Iwwllm1nG9lxj5pW5PzRH0nMMTmBR+Csm8fW
mCQ3zVrcSOU5f6lQAEkialCP7/NHP/t0JHC/WSN5o9RKocwNQ8Q+84aF6EtMFLSl
FZrK/xfCWl8Wwo1KRqqaSyNAZSmhdW5vWEXVybN1xc4KSFnWN/JbgDhCa1cj5AGj
lxDmEMWVFrJtxyb3DWUie47iYT0VyasueMYQXpSoM/X/vi6w2NIZiXB7IInYwGZM
tHc3xuU3Cu7bXMSBpBApL/+4pQRRLfjVmnvvPFcxdjLK/oevaRGn+9BiJoNHIHw8
0V1swbZahom3Cuj3AaNaxLY3GlovuPbyYZ03dHbqQdltzBgK/T76p7ov6mRIja4z
HUPnuwkjaGRRraiL9MVugAUYFHqQoH2gBDa9cxRUR2TdKlx+Az2rGhUJBUK4uYzi
GU8fYleum9Qu5FUWhh2jDrJPkVfCQOsieIDe1PvaByNeQlvMC4OwgXgCy934OijY
Z/vOklthHdRnfQSSVGasvJnVX0RvF7IV+MTBS3zEwTdsNh9G77y/XhqEyuZ7zBHg
/DmWIuoV7xPcKUYVlNDKARGvjx7Gclkm8PDvEp2g0ZaP9107pXQG3dnMu2tftUVL
km1zjDJYZrIJfsz0ZseieCpUEdDLNFZIlgZE9C/yZuM7FMQuAJMPYpRlEojeYnhh
deuqKeyFQYMOk2paTxBHo1qeVTotxmjCV+JBWyAp9pRJlEehUrl2SSzazDWrN/AY
QS8dRcIuMQYspu/y3tOcI4l3Bn1+KhTkMKaHjxsnhKObMQLpZOK1jmo/T/BVXy2K
DDd75dKD53/wDSMXdpdMFcFX6BPk2QKTbVuXZTThSqV/vy44C8fvVlANiKY1MDOS
CIUEJnqxdu8iR6D3J0k243bzsZZXe506DM0yjt116T+nZXTkYNTEd13/EuZ0Yj8e
ZIysn/A62EVphW6deEQxP30hvBUsDVjnWAwU3Yu5emfLYcJLGMM75NGpZ/DByQpC
Su7svbFlPa1RooSneuJNwJ1LUoCUoZtdt1DS5KmIN5nlw4nWH7BCnKRo1mOsnyDL
Etdgz4HNUZDmihsPFyI6T5c7NvUQc+7AJJVbJ/SoXE2/eGRWBaTjf0ra7b/m+4Io
wN5z4Wgs612sFmB5/DwLk1RCYwKkwLQAd8/+ch5r5im0GlrCg47NmQ5CAaeczIo8
wDLUHuGBbkmfCnXTDc2LuKp4GusVC5WcPP4DLk4Eq50HfH81ySt7FdhaR6XFm7Tb
UwhpaBJ5DqzyOylu0pGcISXcGsRxDbmMMB4TZ97K98IqqKGxC9yVmaybkFG659Dg
9x84tmPwyDo+ymyf0ID47MPijcIu8UfdOnFkL2+Wl+4uVWYWAqIIH26akmPb2Ms4
YpuioyhypFxTNli0nO/TsB1kEBATBmVMzPKHbjvMEe+fdD6v3q+c5oQw+4ztcE1x
tzJVfH0RftXFCxT4iwBZf3gBgNdJk6vamjfNQTnQRSNyi+42KuARwy1BYcmPA80A
gE5xhBiyveeCO74NL1uen81dKuEiPznm//DIOpSNgvBa/+MHqcQV6B0eo1rPCiQA
mMinkrQm+YDJxWbbz8FzXksvh5oirViOhuI1fphlO5eQMhTf+GNOX908zEwoBm7a
0wM3KRD1lL3JmcsVauOfmDhvo2cAorqeQIjg62dyCoYFhUVR+4+/dOkQX2Us0Lx8
QjbEtdVIY4wAsccPmpfuYTm4VseXI7oFgF6J9PITcfpP4jEQ8ot38HHPIiFsI0A6
FAO0Ji5I81DNUwvPAkUUfKnOsR3yu5WJ83g4yJwzVV0AXkg7CpASyKGEXHlG0peX
CPnUmUCj33kaqoWEw8xqImXsO99qLxesaHET40d2tvEaax21fKGhME6BYwo35KNh
lf4Se+pAyY4hg7mm2zas4HtzMrGVLzKMrAAVUI0CbIjQmxAKKAAigjgfh0T1R9GT
hv7uG6UZhAmBRKPrts7C2T5V5xlRwXiVzXZfAHG+Q5z3DgN7Sn09e7ZaDXcL7LBh
tWIvCu8rpMgShMjjY6zwg5D6VGxn02nfvz8l2nov9nlyaEU4MPoBUyN2Gua+Hr/H
TTHc6fNjyLyg3hkeiWglkLxl0lkxDAKNNO0XwmdkgSHD8lPCU5D7fcnAUiayhFBn
D7o1YeJogZARbhYeyONPBpuO+GvNTAK+OdgJiFJvjr/ENlY3nhGB3jvjJBl/JFz+
qCmsTP5PRg5eNZP9GOfDsKpyzzcxkStI/pLWmNb5mXWoQxg0E+0TAoLO4F1rIgiq
1t3JM/TUN85XgFvu7sKd9lJlLKmEP8/KsdsELuRky4GcMyQkoVuF7G05/yQt8cn/
/e0eQS5QNYLjFXt7kY2xvB1wNqk08QEw+Swnn0MHNvQKnNpPdz+gMu4e8/KpM9is
IFEYiLR+SzJh7jG46EaeflS5FQBtijQoiGSGHDWJUgH7b3fwGXk+CRiUGw2st0Eg
H8AWVenRbPyHuHAZ9nAL27v7BH55pBCiPL1dxAk6eM/WWH/IMUoKJD2exp/Y/OcQ
PgZ5bTkvvnHgmnfcRvvdPoqW5LJ8QN0JPmEFOdnLhPPWIYzwB3bhDFpFr1YEgtfK
IkYjORyvjZR/SwmmxkTjeiOV4pJ/MUd4nh6cOxu0KrPzintzJAE9d+jSXFtWnc5v
+u1i6W9rPbaNSUihVZ5ioUtWtCTzI8XRtmPyaMgq89Q0j5WrK8zx+9h4XulIjq6S
19eP2jMNn7yyuRnYOk0CRv0dvtkHEqRnjKIQtKxvMWiSNT1YEDHB+4mTiLlxJIK4
hQu3UsAx/8y9gLOf0EY8kOjaCWYfcs8rDwlzv1qpzmqiB6l/hlO9vPH+C4TRhh6L
n2+SeootcSRIJknoxOhsKPmUQdxQISNyMowH+36ICsJi/lfUSI+IBUFdXXbC9/0V
OzxkjjZ4515pp19zX+0NM8MY5OXwHpLFhEVzF+uDx8MBXifKb1qm2BUYPb5iGuja
/p9BsqC4O+azElttCfx4WbuOnKNZX+Fz/d0wVXfK9+VeKp2q1+GEZ/jhe1Ji2imv
WmY/40d54JRNjqo+EbBquFzoHHjPO2M/Ik3t/TFp05X14m/PVSdutNtMubMjDJoS
6CAsQzLCw1imxBDDxDQIfor1WxRgG6nn9vjCZ+S2W5U39cgB8azkVuCAWn7lemJK
0dYKe4j2HyBlk76pQMVp6PrTdKmtIyy3uTqj1vgr77FM2HKjcfoK3oUMC1C97KU6
caESjGoC7b1SEICMgH5LZ6WinXt8lQOlYV6KvR9F+9dRjZH9GN4eqIijEjM3AEjM
iIQarmm3nxnlrTpxeKUvvOK+cCARrEk822j/sma6f5RpW8WRq4sPUrPgT0MYrzTB
ZhKaOvZC1ax6ifcwtA8kjv2guv+mFOMEAFDr+ocs2/KQCgAlocm0KhAL59Xxeuwr
AL52OIa/+b6X4r8M9OoPatJR52UcwmC51g+jBHx1jux0Kt6TdEJN8JyOse3UCKXV
FVROCDl3Fxh2/wLuCw6LV250f0k7+0yOI0sVCtl0iyw06S0K4Qe+4uDv9xU+svoa
CgFzZ2SHLdeZ3JME9soXVBTkiTm/DSDqbfQb/79HwXa2WlJsH/hPgyJAy0ja/JZD
iu9PwtjBWJuGRybe5QC8z9Oi/6KeVQTAPDyryDJC421VDsiY855GVS8R/+3+P3y6
RmL+QPNtnmoX5EXJaLGt4RgzKnaQ8tt94pGLwtOFxamkFxORUJ6K4qUFXMtDyOEm
TiT7WAeub+YDRVJ8zG/fvj7cStMJ0fBvcbKajJVp7CXcvd+RprQNUZTEeFfd+89G
X6N9XMqdauurc4plP3JZk4/smznIzbV3rEjot2FMuT1LFcLjkDRyOpCojvlHzoMd
5MnA7eCdcQfB8GPZsQWJlRbTGyebbPOVA6vHJjtBNcwcoEbIBSl9Xg4ADK87YFPf
Omd9GTBueoZKLlSNGB01e2NfyObp8XJf+UAjMpYG9KKEL5OL1jQTmIY9ljBAhu9N
VFqtSXHwbaxAME/EcffGldTVgske7anjJoV/vmb5XQDrR8qH6u6UFnD2HnRX8vJR
QI4jVbaAFO0RDBgncgx2m7IQ5K5eIqEdVx4ud1NpCNNTDbJNQgVsMjwzLlaEzPa7
tB+APNwRsDm1drqVvyWO4tdUtK77fOidFqpO5Sgq6L2LcQjc3QDKpnHTiS2s5Zs1
ylEuqh0btGGKym4czbaHKA0JhkybOui6jGXoiXc3PaJNRQG16JUEqz+t+O0qV+Ov
kxLKB0l/DP+bZXTadKrXgFqHX3KLZgR+RGe1cYYsifzYlsXBrqd86VELYAkv6F+i
t0T05ZzqxSfA+BoEg1PEwQUAfxvqpXNHmKUtA6zIeycULAWqRqIeHjsbl5cEzxdn
XLk5VdOrYDIz7tWi8B51BjY93y2Wq5Rmpv9SrNYiASFT8Csj+0uR2Xdw4uvJ9AYN
AzgubwPLmB9jdwd2DNyk/zekEvgDH6a2NWV5vxtPk57DSlTM2+NDTl5+2WdPF56M
KluLIE9pj+XR4ONEIL31RsotZBJvoyxfxm4IBdIPWduAwkScpADWyRAgfXZUD65M
A+g0W5uwKL2xrbePeTDzLUi2Jk3XxwYpfuMRo6B470m+EF9pGE8dwk/HY3p2sIGm
X4twFmxc/iC7mLGj1/kY3RPnCXs4wrBgYZm27vmy5Gvo9NmHghosQtOEgkkT2EgX
wsUaOeBb9NHBR4vpuL8EOCtriV82zCv++jJnsrfk8pqww+4x3h2cN5p8JNJqzJ4S
wKrCPkDmzO1Q8g2MxapSrP+DRrK4hE47T1zQkMMvA/ONUwp90qVK2LBHO1y3qTV4
cLed9BbjphxLv6NPLNYqSaALJtQPJYY+aE7KMSlf9Z93HMKZ9LHQ6hGk9Cp7kZ1h
7XM/gfM9/guCtdz0MYjZ5DUpaKBcBRHxT0Y6nphlxJrJ4qh7iKo13Ywr/98++l3f
n+YmPqHyZt/dxi9Egt2YBdnOW8aaxYFZSzQvMGVQHqku/w1NTuA2gijI+v6pGejS
Wf3snqyvZ4r8DpNSI3ouwNYe1I7RpCtGb7GfF6WbabeyJ9h3qCOmKTLwmeG9bmBg
YjkMh6PxkAzquVS1FS98zJNtEar48WVLnXhZh1zFR+iPz2yyeiB9zbbPkbVZn42Y
GVzmxswfnMI8DzyL6a6waFwU/uL/1jFB1Ml1lmNl2IpjhaLKEze9FDaCK58wLK6C
83nOkgC1INBK15hSSOrTAjEElX/8hQgbgdMUWK5EiVZ4QXUUFFcZxIO7jIEw5RPw
XBjy43NwYISEsisM6cL921/6qVBkIZVjDUBBT6uw8glwzBHfGYOOCuwzUcCKROPz
+PLJtu69sJbw/Y+OPnp93B1q9MaokJZm9Tk1PDXcDcpRRV1gdwmJdzELl0BgLYRg
PafcaQL0Ar4n65QV3Ygh6eziVovEh1SW8V/s+9kWb+gMPs4XMbCRHfM0FHBGAM+w
TnZeDlazNpJVwimfeFNOP7exKYwISejO+3RHZ/3pd7uUOBt45PhlyKStbaKcmvTd
UouBH5Gb5CYg59c4I/eOpcbLgD7XpJv6uCthwWTcWu01BaQiKSMFcaoAeqC/R7a2
9xThinsKU5Y5SKaN/5Ei5bGJvWIO1ct4+AtD8pJUEQyHQbcQnz/hHuqKXHerrmuz
k5oNGGnnmRwxsieB9rntC00YmRQVm3xs2bfeojt2ovi3opwLS8/LJ5Pn8JhL/3OA
x3VCGgN4JBNCVYpH2XuMNWw5GZAPdq3i0HOZMivkmXJveSdMGngAJtBnH9c6Vu/b
nfKnUg/aF5uqadXKL3to9l1R0GKmGN6wLDevGSO9ptfVFBFsnoZnbOFNuBhuxwv6
q3rnkymMe1fguaC6TMDyz1XNctYzyYxc3QsiwmXsmBzts2kOG9gtupVVq5cuuQl6
TaBvthyAdl26lRVDf2aaNMwz48wLChQWCCyWEdGHOSeelvLED/xh4knbtItTeSKF
OICyG1HS5KTTGBMLSt3NfNMB17VKgCd4QjDhBXfYLcBc1XrA4jbilb6LKejEQtpf
Qwk4hQtwW7BDrp0ijQTL8pfeeC4nCHpkCFDw0mjJUe899IieKdDCF9kXpvpYjMQO
YCLI1xl3Qc0zAO8NUWjBkjOL2FLLddNrysF5F40udN+OgIxDobymeMOqH21W9Dgn
gSCV0M7AW0BaQ57aPXbjq3Y5FCdNliF4LqneD8ka5EnxWbUpycM0ojRZt8RDbD0E
oJeNFedo2s+AsH+HGzvWmfyNQizKlCOTgC/VNtV32v+ZZN8uGSzfAnby0osMQotr
s3TR41/36JXCw5STWJe3USBgRuxKYiEiEcG7D0Ops1SPMpnDKdSpX6cPfPQZwFZU
J51akY70zTWbIM3qZZ1Wb3pYWgsHDWIbhv09nQScIS8EWUYwnDHUzZxJzh9bGCOv
Mmc4rNPoZBohF0R9YszuM5BRthUMTBfn3v7xj3cCQ8bOj5KdqBTA/+WnOXA4MZnT
H+FGe/+eDXBsUHOs9V7VerDlrHxv3xfFHJ6Glmsl2iMjcw+0293dUq0tbKwhQhJj
GH8MFjWpZSyNQleMq5RvSift7re8Q54CfX3DsomI55oe5L/eVO6auI90TMM21RYm
hLg9m+tV+L5SFV+QlKMjUoMe+P2NOavt9cu8yKM4RW7jJxTYtlYhP+meF0s7A1UI
Fb/P0cVXgYcDDpFRctbsQs+5JeA4zaxMYWz2GXTjBcKwSyp+kVNvaKtaH6053uka
kFvRFPIasFohpj5iBvGRrFXeB3a/kJnbXk/+msCLcV3tBP/KtFzjzBt8V8vX/Oh+
xZf+LYbdbikEQpEvCJ2+wF13vx7BDH8ealexFMh9NWKh1oNJqbTHFSfT0T+3eOaB
zH1/kLk3XkWwHDdE4Aih3NWAUhyoVe6B9i0DQW9iRFn3ZEegs3ev1Jw1ynDzUK7N
KTQLtCQtzSYnPKegPn2DBSXHdWNwxN5Sicwtyba8rUIzMjgdrJqco7HURJ94PPmI
duRtSJAi50BW4s8VrEbkrw9TM6do7fTKiDqHHL4LkYKgdcDWD4I39l/TA2ziLuUJ
QEps3R+950g+oh61eAEYG7OnQdVPJvcmEzMhUpdGupp/ovdBtM/8LsWurH52cxPq
/dmlxzgIgV07/ImHmzDU7Hxpzvax5LZf3bi8zRD2aj3oZIkf2PoFuNEIwwFRA/LU
gx5kgZBqK8XXXkGxHvpCEry5nejibNWzz0J276KBQULStcA82oyPfZJLaoLMfvFa
69xjl3C51XRhsgDvLSL/po++gFDb0KKFAQ4iWn3UKa4W69NjtdmYz3+T3sqXWJuQ
JEa4+Vcx+SD8r1IqiycJQmMJ6bdIZxoweZofjSj9v0RDP7L6I6Xe/HZYWNM2B2CT
3BP3HTtUluiUlkSjtRUqxrntE6GGsUYsdI6MzC/KXJmBIynm5PMULtPBofk9JNGX
GUVZb4CvOSHJK98oFnZzEN+qtBb5O3Rj105plmxJ67aWpHXMYnP9D/JaNOcM4ki8
Y6ygzBwu636nIPEoYML49vG21FeqIx6arORuvPPZO5JbjsLD7+dBEuLCrYoegPOi
YCN0CDjQHGy0vREr9i4DmvpV6X6oyQBH37LEdNURGSrQJGt5CE4Pv4TtpDBIsAus
fG8m1bYybXl+OYTJv4YPfFChSwt1QDDc7ivaK27KEK1vugKWT5VrtKrRLa81v3uS
XWc61VlzsThNyqTdf7hBnlu2UJ6hjmoNo5CEWxfXdtrAuBf4AgYImeTQyibR234v
fgSPnI8iYQF4a4aeVRjiDIZULidl83lRFxW1A745CtwHtnP4FL9HkgjUIvjnKQTf
dXxlAguhxzp92rz5g/st5sj1xrJCpEO1haTxKCh1IAEIUxzy21NQ6W1UMJ87/tuB
sChhyiopHpyxOLUauXaDOdqxqpB9U+5/snqxgXANW48GazyW9BYdNdt266CMOp72
9hVSc0GfOJPLuNOkScvxKkGxZbQBG5Ga5qUWefw+yAbik96LveGX4rJ9CRVF88yT
gI7emgFYO+GsmjtJfFj0HP+U3/NIJu15nbnc4sUjP15DgyIyuDAjFDFAWKJYeofl
YOL96KoSIPuUWZ8cGl6QqvSLYUHW2jmbo2RYMvk7S34La+3kEpmhVpKvn1JKpHzZ
qzkWwTJT6JfU67vHWkRGhFaqsGTYWHu9wDdLE6HFPVl/0iy30WFR1fwLL12dryGw
30wOewjNiXFnSFUZWYSssBnnxFgWk6W9bGuxk63i6d7XjOwG1XVJbE/tTDQV+Cpi
8gN72gRVv/ChN/Xl7VldJB+yIWqxqOVO32SxYG5OyP14ER9uF0cQLjjpbFsHYB0v
e2OSnaAtJx/Uj63Y4kvkkad5LV7pYgg2sOqsCjhuNmSP2EpXO9VMkmhnv2cF3na5
O9mI0nxNEWHAJnZ0bTgKHhBxWeuMb4DyWAGqT6uMIRTE7rdj8PXME0i0nDJISbmR
DoTN2MN/SYiwa7ujfmRR+VGCb6tZPpFnaekibSljx9v+pkvP3fzquVXr++zqcUhB
lZyq9YAJuYnDnZ56iyv+p1DRHCmKIhtYM6vj6PvJA7q7dgT80J3lzTnMc3px4nTY
xh4IYGk1IkDYvIkWPsiwFimK8dPKnt1f9DmXHmAjOQ6ODABAeFHfuYLwQG6ViBn+
S5VProfSgoc0J0EpIDgnNnJGZKYl276VJSAWoIWBEToYVMl5Ti/u8KIBxLyz7FaH
D3ErPKqxu5O+lxWPXJIlIyoryVbAC+TyGXpV3MqgTDRLYqSGWF2P10U93ZXv2/l7
ThYei8FjbP4mydZ4ckzlLhtWGf1hvA83u7Wn8a+2+o12IRCTI7vcvmUowt16xtO1
llccY6s/yLfsOiWeaRwVquLdtovDhMr9p2JXUhM+9iFz4ltLeuLNWn2WxyOcSPKe
VZPa8kgma3xSiQJLIUY2ODeYv8/RY9LuBmqO4FnGmlz3QAY03ZfuGxMxvuWW6Qjx
VaZm4NTa/A6MnMWsj5h4sZMLBoRlIiitVa7m1SGxoHLDEoHeRq+I7ZoJnyNJl5TI
mGM47+MKEqFrU44HbidGe+nQ0V+YsLDfO9YGmJIBWwKWV0/V9IggV06WunvdI5Dh
Z+Pfqjjacme3O/X0TN2lybwu+3DGA+Fjb8cuwYtrXOe/PbpNa3ePNJGeDxEy7fkU
GiiQGn82dC1OCRSrqEo49qR40bFPwIQPRak2zHv3TI92kWF5pgXtBBzrKvuwArjg
7ufM1nfDbjli3wU/0wEgUCm4gJFnQ6T3awHrvvFho0pLDIjvb2CFtUg83GscTUox
+HyjcpS//HcWH7rzHzCJBzfdrOKENATrXxrKttNOc23EvGincUarEIylY94+7rxM
Q1gRn+B3k0fFX8I8Ebw1a5rw/YFnivb1clIT7g/OALAICdaABDotqQZgFlAZtLX8
HgVl/PvdtpVSM2m9geqpvm0bC6YGcpO2NDHM2NKm1tx7gR+wXpkvGF50O8q2G6m3
QAm7SwDZSHvKnkAbBNqouaQFhiswGfzRm0mcGC74beBLoV/4WN6G5kxKTLaUOanU
hUu4DiNywBHwPGiflMGu/jNSyBy8bgzvY7QfQmScNrDEhE5c7tskmyo7GhYMrQAI
PiF6hzbLEN/DRfM2TJn0frrV00FFKHr9et631jThZHzoDdj3LgR03vDU850dyLUf
hg9+7nT1Uy8tkI2vWapYLOMJQbVF0zgdfTJwdByS1TvRop1fvfYYzB8k3htGcs73
vY7r2eOik0NKv5XrRT7y9LwxB9JhMrTXbbvY8G1oZqAa111Ny3k7m0WiyW8y7aea
wrJ38Za7BnA2VcWn8ok/elsd6ttU2l1ll/y3CkyzhoUlDSRXduuYAJ3/d3K94IDn
BDPSF1tuD3qBDdvftV2dhBnEq5d1tfpC1B3ALi9G3tJ/eBFieICltL/LuWJQkqyl
FA4l9XfCuBGFO4a6ejVbby1K2OsXALkmhbM9KRgJuO2932NRAESULXdokWvKns4B
Ni/J8UtSfgw4F3/NwPiCF1CAla39PuGjuqA1lGRCqlwkcqVB4TM97xPlVJS0Jxjj
p0dLRmh9GodUfXGVd2NlcS2YokstJ/yVU1M9tMh1zcLovTpEySRn/hFfaiq8mgHI
FWHsyZnY209laP2npo/vcpaqLTtC+HWfIAITnqH1tggbwjFj/1QuEN80kITJUTBL
0HfkByGrTPl59bQ1xGg39mx7NWyD381dEIVTSCMda0NuUZWXGUVYpBHnEHQaQbeg
TqojPaDIX+Vm+ZmZJRqG99jElm9kkaa0noFGjLuQ12xQxELqiJyMmYLTvSlfiAEP
bUwbVM1pBmCleqIa8dtXtwQ7ZlkG+MnJ59GFAEyEMGcpSESafLqt2BSuyXFFGlsk
jaiasooDHfQ9vOxRm6ZOl8MTzE75C9/O8sBBCm83SE2yOEs88k8IDeiBW4qA2XSk
aK2m7yupCy/1yKSJ6TnIIz1QtIxh01fg/EiD5LcgYUEXEhIu4lGfUoR38hy4vEHk
49pThMOxodvL+dLQwtOKvZjx4Sup1E69keZQs8Wo9LrWwYzOUxGw52PGb+/DwS1K
ez6oPq7g42pGU3u7+wnFcWGXBVuNE7rfgpMB1Y//yDU9E2dBsL+xSDRDprvB0Nmz
qySdP385YVx34AUMRs3/PoV8AQIHA/1CcJUMOapqaftGJCNvu10xmn3J1qiTk6fp
uHMOqdQBw4rjl9yoCR518taGu5YsZlcZkFq2qPcT7g2Vp5pPzaspgl3px7ipLrh8
26CpM0tdqLn1uZZAnn3MJiQxaBXWOsb9cSAfE0ZEw5IUEUYYxoBz50NSj7x37a6B
2PuKCsyhiazQCYLaSiaVZ8iv3HlU8kGDzJMp+QNRUMxTQA7iaklX8Oi6DXeKpdVK
LlStVSu4bW05psKSBqfWxhuprR2RHFlYXDONt0/nIuAD/FBJ03QTHwLdRojwn1pX
MmKrgEJoiZv43O5zAyJXEa1obrFlOhOxh6qBCCXWVAlydsDe8KaM6xe1Y/NrcLNg
JsmoxeeCViQQD0ZdcH4Z3d2UfvfSIxTHm/TRT+bTjMQ0qo3Wr7g+7hJXlXct/JsG
DswwTL7Z7hD8ZV3EdOQwnxxnHmsFPOc08ULv1JcjazMflgk8IlCp8inDCjdcS26K
VdmLyROYVjMB9jTF4szXJL1j0YXpC7E7i2Bjy1d05QlYmFN2PKXS8+Gxh4l+Kd/a
z3Skmdn/I0/bnQKtPNwzjj2B/bZSVkHU+HOK3LYUDqxuPH3Zx7Ni1G8CtG3CD8dy
yw9X78dsDNNGYplmLVWGo/qC5s7wNjOmI5UPFeHpaNe0CTNAI/mC42wiQq1PlGRL
QjQt4xv/cyg3Q20n4CV4duqo0i3jfjPajwedkwGfXZfbMeK3LTfWTaOPgjoFILpW
SWuHHB+KXhr4zak4qCIh1ZvGyXyP6n5TFDjncfjSHrEXVhmwOt1sr9YgqZco4KyG
81uwZYL8d08tUcTrc/34rV6vtHvmf9Sy/TwjLzb7HHJWstBs7XBEa0zC4/r7udvV
/m4D8otEDn4ueqeEIhCbnoUoRsn0+EqYE1hbYBLXVQfpmqosku37jfSKLmqskXSq
A7StQJmnEWrCDRQZcg618bK0qWRNuJSiyGtia8kG30OKULqFa+8AZ8FbtAZvVKVw
E9I4EP7CNY7PwxbO02B+nNEM86jPKoVJDgBZuOXb03UBW1SWjR6bdEUObhnwKp89
NUxPXGQoEbnsahN00B2KcvXhDHd41YPN2qfT20eM1YqM3OFeruFiZsxPQZ8rSqrz
0fZsyYkkg4vd4fN6SULV8YguOZFyy8htaH/M1GtP7kIuQIGUXPsZiiY/uYEFNSmx
NFSr+Tt9Ud/fTqsnQHPwMtIw4WMIMHBu4CUDyDzjGoXEMg0E/WAHlhqm8wF+WzWY
4aLlVCMzBELE4838oe61dIB3rFqHNBgPQgNr/TfFEe070ko6o4Gr9FIg9ogORF0B
VLYKHjJNDmjBTQsa1V06ZvGZZIxTRDe1/qaj2+8zg+PMNDEbWcxA8S38/ZW4i4IW
6MggZFh953DD1m6JYVCTRLdMpb4hS5GRrcZYye3ql+l4rzOFnOeGO97Ac/xc738I
Qtp7uKTIe31TVSLHVFfcVEdzkCLy+QVjL60FjPdHpZDY2bxMwe15zf2A1hvCtl4G
6BlGLdBEoikbwtShzyJ2ZXKDfqSpEqczcwfUXguVDCh5bG/HJAb2KLdaeXIpj5j2
GpEnxjBAFMut6fedXwtlqNDDQNq7/rgon/UpMN0l5jqWDB+g11syMd/+k0DV2Hp/
Zc3s5XfFT8lmBeUBJ32q/DsgbZp/xRlsMjHYbgyf3t97DfiloU5JJ9Zfj2h6YxfM
eRaJuy0kKeT6Xc1ryUmBR4Q5p1bSGj1bkuXzq7m01vb4y+HXsWMCAKlzufdbhMIs
WI66USv4aHGPFyCA5cGEqecPc1ElpxtwYIy8wvymB9+yILlRdB/LHuYKs+UrVTeY
Yzsvdq+bVjq1d+STm6A3ZYDbaLpp94EPo7Uyziu3UFguOba09I/N2bQQ18Tbyb3K
Y5SdFcW0jx/f2ydmouLGnSyiT4esC1xPlnA5lUpnP4yYuF6RqtP7qUFVuY2WJENS
cR5igw4yZC8Nkgnsya3Daj1ZKwcw5/Fp+LVjByNcCw39k5pExMhEgG9dRLYq1jhG
8PA8yEoaHLosbS2nAUWarJry5q4jLPTSHqc96k4Z5qndlDJWp2jwK5T//HQgqVKW
Gg1sXFWg1gAebKl42R+7BwyWLobxmmiwC//MNeaXqsMtPyjJusUsmSQLtU+zE+yn
fgrqFeluiLWsmsJvHFTzTyqQY8XUYVm1FMTFhrsa4LPb6vLD4QFWHVH6XoqRh6ok
cMqvYJCJD/w4dfeWdwbhlsIDq/cPZGlXPNEViO3yZottr+7FFCXUYqznr6vgBJFE
6m9jqjrUdoj7qVJfcHOcsobf4ooctGwytpJa5w0RjEBQSe0l0ICXmx0CINwtj8pw
cF0yu+71tdbXZrscfq5b69nT2aLCiHjKtwT6ZwjnFBNp5C/tgf8O5ffKRsu9uX5G
j+IaOMCd5LVsSaM8hVFp3Hvi6lbljb/DvaiQz/3yaQP4+W95EsLGIpUfD/+tpaFK
ZKdEnRKssyGY5JZ6wZlV4VoPmUXIX7BWpvfy5NfFt+UmtW/PSSlHw3tqMCqNntQz
mYtK1MfBLeJ7TyHFBVR7N3wKFCa3+63DRcoTRW6jFDTsQdaVvObjTvVDfD7kr0D0
j71zB4OKQjrbr/cyLOGwXYLLvkpLXssBGPFmsWdgAiRyxfxCwVFkNZ78AxQ0CG/x
dOatyDgoiMvFIIEy4r6cbCEOWwGugKZgl9ZmzybVdXb+F/BKO7uGeiDigiThsL1q
SNKpnEWCZBmOCZoEbwJn2R25zg7Mq5TZAnrZfBAoP5/++rIw55DNPic+MED1idk6
EVr9aksCuLYMPgtXGS9S3+XlHOooulcMcrAY4TlM4rgVTEbqtk3kO3QmahfA5/YE
TmrJm/eN1WZSUdROUTVxkVTOSr4r67kvCdHYNTmb4AV2uKaFudQAMxr4/Ft+OtvN
Orfq0ytf/icamTxnIREzPtsQLxinmsOcTucwZ6/3kqJ2tUvfYt9aOWZ/bQ+Wfo/r
B14/dVRRhOqmMf40gQIVS9VEoLRRK5waig50EMNJ7D+WgLG1jfgQJLwkQ8bH4oc9
mP4Jc11cEZawA5Ctvb1CojcmgJCzNqL2lE6L7b2fcN/eH7RgJJFkO2vOKuAQ55eK
pd3rTNLaybAS47s/IKDTgKgxNOFVPGhF4DROHb8hXv5cWJWVhMUSfAspgyKe/qXc
m7+ALjKF+cqjKWJjPdNSWac3BQ03xcripdKMYlmvK0IMjKZpVnH0k2FPswCCN+V/
Kbe7+iS0oGlmwxQhv0uWDqHHAZLhyPXewO/YmuzVn/YVbc66pfcWpiw/6YSp79Jp
JI4/ZHftn5GEQAGjoX4QHMq9vSl1JfohAadESyu2pw5nbDFr0laUy4zHW3ivlI+9
j28qOFo4TEd5t8Mk5P11DDtp0/M9/om6HhfZf0ZzVdCVBtQXG9F38yplVbJwNcmp
pbqh9Y4QB3X2SmADqC6W677C/5jtmNtUhPRF/nwQg11bLeKj/80ZCN1+X7UO/myt
y4AmqtGErGCqBn0qKVxLFlQu1aXEQoFUgzrYUuk8V6aGe6jvVvlh2izLXlSPo4/y
OXjis3KDLzU5i7SoCyOAqZtKkt1BLOh+qVOurx9evCT7VHuojzZQ3Kq4pJ77Zcs+
yXEjqdATd0+JRMY0jWfX8Hpw5KL9gU256Ql1RMu3XzHqWh0T3Uhtkz4LrUcvB3Gq
odFX//VSK2v+wASUuEsI702fYomN5htJxW88xwbUcQaJTg4evcf6UX4BKN1wnygb
yFEpOFVijInmiGDjEbTZje5vi2z9FqYtSThT/qcjt/yBXsfrzQP2iXrXQj0TG4pl
lOmk6mJhanVGbkcAEXSUPb5Y/OwebRPwndDl8v3+HNDDUMhY5fruMvr4ms/3Hkpw
4inbtcuoRG6v6gP+q7VN0JVAzxFEmF+Iz7H8cqYJaJAW84FUZFvNCMFizMyTfQ89
vynd5m02g9rWRI57UmUpj4VRsiBTKnYbKkB+fFt2yyi48/oK9fkbEY2OEaqbSp8L
29WY7dDO2iFb0S7YhoL2zXK8LIADzfuzbrbSJziMWsZLWYOGUotHWv4/qEas5yfC
tOY1GWPT6GkR/CEfgUSchU1/ZTtM0N4l5aYOOwuWAIgVrm8wCeNa/pIA/lM+BhR8
Guz0CIxQwrln9tAXTHbzL7/Q5vKUO0JdeW6lQGqvawCIosxSuiUIv8dAsdLPs51a
UESv9dmYdJLpJDzDAGrQFCybYlLQ2cUPKJi9xNrZ+OOzvzqR4feZYiMpbdQWfY1j
NE9mqdKrFkLn377Ej40E5Na7kZQi3MRQBHqL0p0v29XLl2flPYo4v811LolYHg8G
ef6j7LwKRlcASJ8PpD2RQNifLk+mWZXiqrRV9z5UuAx87frfwZNQAeb3dw7M8nhE
xnd/1v99l1R5p9BFkWOwccTdh0jFKlN88itsitBiffoLAGjVvZlPdMOuduiNupQN
Uw9EbfGJj4mWA3imr+m3Tpx8oHg91LebaGHAJ5VtTcSt6FE9WBuc2iTW/HV/ODef
W1Nha0ruJdgyISYwDKu/Z1YM/uqCLNH5DggzQmZ1SEeV7PBOtmwo0MghdCqYsKdk
5CRJSrPAewHpqSO83qmSN1WramBhyaK1g5wbb41tZDqmgaIGVwyN7BGr3xJ5KgzY
Bm4QNzJXwyHL3wi4Ld4fMrzXF3bz4Y2zMv/7X7+CCojDtBKfrO66GZ+29gOGaXiE
qq5trX75/JfVnnBZGloEa+Ng/uvP7BluF9L380MrHAAawYtuOfVRRsHmwj7vq4TA
Zq/TEU7fwPouuYQ0abjzAqKsy3ioYonhrAhuQWKfAUCXOQRFAVYQyK0spo+6FVAv
1S1RrCwFdhTLx5grUeXuY8dJhLj+QvrJAOtz+NlsYmgal/dz+xZcT2IXWdJAD7fR
ujDKD9esbIPbupVku8Elq3zyk7L1KvusxczE+qBgMM1e8H/3QTpqaZA0CZ5w4fZf
Atnon5CXJEHZ/gQOLoNZq2UG0CK4hUKwNG1sh0uyion7YNzDQseeUon1dw+RXKoI
usBOnJ1o6NptlC5iii/GK+a4mthiPg1mI4QLMBGs1nIqEOA0JjZJbYr8L8+Zq8D6
y4zjrM6QrmPDK0KAjXE+EsqhA6TSHYn9EVag3zalR6yB+5QXCBc72UVD/WL0rLaV
pmVAgaRzitWDpjlF0166tkTF0FqyuesdoJ2Cso7xCmR+yi4RK7uAVO2m1F54ykrL
HuPcrF//AoQq0kJWI42iN60QxxWhCb+FM6Qy87hL3Xy3N7Lt4yJMk7DEHSnBJbh7
8bYj54G7l08xn+lvfk2pA6Sbk5EOxXVOHBSErDEIuqCrEZnfuiH6CIpr7OESUqoK
lGzGMjwKRwhSylsQNLJnn9n2yPiJwq5aSKgp45cMRBylcmkNm5vWx8yWz37SWOaO
rs0DwFBH04kuspkKN+GMwV+9YTuCQn1ajFnLzMoEuySGoL2+F0TIkbaCeS8Y8X4X
IrzUu7Tp9ETIScim9ME2SIWtGKTNvRoZ1/Y1ZLo37mFelodSN75UVnQ2L4HO4U/3
Ea1mawR55NxFE+jihVCQdKjcsIVyEuYe53T5Vsw7Q8GA//cuC1JcOY7O4RNYk42l
7eedCWvYzbiaXf7qeJfk0MCOK1ADuIN9g9YuorrXKcKJ8bgE+Xh3LyZzni+uTC4o
+8on+f1358AXbj7qJVFtQLllbdqNinWHVenWU/0sCvJMw/7/IbTE5uVOA4Ygpf2u
xnvk8r0sfcMI1tWC1VQGFCZG+HXKPcEQm7fcxPq/Lq5BhYfKi95+Gl1MxRE6+DR7
BTl5o4Q0KzQV2SLeaBuOB+l9FBeP6CWKa9R5Gb1pW4BBxiLCBvbZT+5U21VVsoEt
VG+RJzs+L4tgiQdo0ravYpftQyVortFDDXMBIoa7e92cyu1B70W/kKdsiK3GibNj
GfeyUyp+INWd8mf8PDgx/My1+OGZ5nH7vgYw167DbwvgvXOk5KKilmZed1Z5/5n/
knxw21SB8InxKEHHif0oDoqOEEIFpPx0v2lZJ0tzyT11n2VSg5Ye3kDLt92tpL5J
8HRHD/1S+6mxbe9tKvJ4zf3Ls/eIcf5amFmcbO4PctCs4FbjkqZVjlucMJW85Yhp
718CvN7MdrM0Up7rsyX61ruLJRobk5mUH6cbTuLmiQieXrOmnAfDT0t/pxxDtIXw
YtqG9Y9CQNfNhGiyr5qUGTmiiq9eWrkI93E3VE5MOqfCEJH4SQv2NaMxD4vCcEwS
yCLdm0z7ik/3QYdQLATU0rOi9qHQjtqYMZSAcwMdH/kMUcNBkm0MnLEkf/HPY5D0
GO1StrJAayxvftTppKKha8ZTfF+Vl9edNlXVIRhIRE4aW7XPSfUcau9vR/GK+vvm
vRVw6N3r5+UEOMrc73LnBUVSC2zF9BKfoleXyv98MXybnyXc8kqh2fCS+Dkde+b+
/37rCTO2N35d60R1rzw+6JX/bauendc+9r+dZbNnQptPBsn9p3osVDbRd/vjYhrZ
uGufbDpx7a98kNlG69DFyrz/uDVxshIriKmlzxONCo747w4ZiK34F33vjxG99f+t
4M9fMfMqjPM1pqDseYSst7U2kzqnWNvBx7NX1gAAiC9MttFCHWOwNB/WAfE8dOp1
phse62DOIM0KLMTpEzpeMzUKSKm10KR9a7gCFXW6d/NOaYmAuWXa2EQJqvvUaWnJ
9Ly4DYi+NOSUHMN9CRvy9/bXKjZ2vC7dRuU3MWt04O6E2E+VoA2nRCjPrltqa7db
9JhUfI/4golvhzd4+ZWnRG6fEwe2BVpyjBknauFxEQr26Z3kDxWrzMs1UI7lc0Lv
sxE4/nRE+h0/sJYWTrHibOH+up+o9XGpyS0uiULfvC000/40jnx4pBtBcb763WDs
Y+62QwJDJcJGIIZbPLijdSk3SSFnx5S1K2fD1e787hJoc5dbtWCBcLN388ikMZ+N
rVUdLsFuYLyRWPkVt//vLWu2T8SVpCsfsRVfaRjWnEip6tlR8GfSTx/4k+dkBD+3
jAt5QGVBwSUMBghozWbG9DpD9Hj6C2mvBNt4YHA0kCENRaio4aMRWHHQRuEeQcDA
5VxMnn7/C1PkpcDSJBrMORUvmeYOEVvg6fn4mPjXoNMo5VGDPNz1FRmcNB9+XyMB
z5d6h03cXyZLosjrneVswp9UBz+8z1I9xr2bDAkuQVr9Ndv5YcMM5z2+qpFnHQim
Qw5YxKni2nvTHRobBMGdkXV5rIaRcQT3Y9JXRYPCxi/kM0Kn3kV60cvswEqtSPLs
3ubV7Bor4ObnIQmAQ1KfbZraIRZ5WFNseQE+cJTad9u9dOuxffOJZJFR+ytgUEHr
dWSm8aS8+sBI2h89ZEpfK288PDSe1zaNJxLKE6OywpooF5jjnnfuG8NTg/Ns1Mph
pyWqDaduL7ltSD4RmstmN3liGw0gWxdUxH4Gr8oKeGUVUcBps4pYkuRaTmbdklBV
MRlJ2MOYpCAPSZzM2iR7zsjmntZv3BoeTk0fF7nsIdz+qtXX8B+zjQjBZVaXgFVK
BmhEF2Ue6HGS4GicZeFIxWh9Q2iyzs4yQG0cSFWBE/rz2Q4PbUAAlGkwuneUDTiv
H+7KcVxAEMAaYGDGzcmXm1Q6GbDAAnvVpXAvHDhe4+R40EcFxRr8SPeTg4rZayqx
YX/rlAG2OmIyfkA8HLz8OUYKBegnxQJdHPMM9a5rTtpkZzZlRZo22totwzYUmplb
AG8qa7zk4OOgUK1exA3MaWsOvaNLwZ285ORGhabMwaYb99BGSh61u7mki8czkhku
JzXaVqMKq8HlmkRs7BZLYVkdQYhQPHKCC/MqVgNrARL65GpfUSr7/lIwQrYDUh8a
fgMrI3UOqyEBTgv61BkIX/wQqcqutIO8UE+oC0TIW2qn3ZBB9RtIRaW1iBJ4BSwX
/dXNbD32mU/pGK/yxLBMmDcwfinkq/BiIW+n8Osn2UXVhZ3NSfASHc2iEVzQMZQz
96opYtI0QoDfrMxKCdt3Ja8xvJV+vNepDoiAdCIjq9oxkPTIp5ps465vUsLJ5+4j
jsCg64P3/ex4nyu4p0RzsNlx/pZklkYvebNLnm95Pi4sXoYto/jbFaoOJWGQPt0F
FsM/gqS1iz9d2jb4LEjEFNOPIWhNvmp0aKE16j3W3FC3cyWDvTxJsDor9Pd/mveT
nrVybGg1ko1O9TBqOTyIez4zmikKbKd94N6wz8WXKKaagM24vFCe0mBtm7jrBAjq
5cy38dDR5QDcws7uUZdGhYn4ZLFmDo67xKRVBTN4Xt5rzhKpZKSRRT1QfEXmmvJu
6D+q7Lvy5vsdyyHxsYI5OELWFWkNnkGhjOXM3X11ZJUmGvm5A7Xl8TsnM3OAiE/Z
/jLx91FXAtSZSpWeLRWDMFkWNi33J+eiCkvz4B41znx9lDLYWK3RSrOrbfootIrl
ddyuVtt4vtDB4Qy4kbUC2Fg6Zzjoe/IwJa7/naDlrk3vhJCXMwyXyXMP9+HvUDHe
VHaNuZa8N8rzq3hF7mpY0kHzQn5H4CFa10c4UAQjexkvnshJRyxZEGu9B5YaJKpb
pSimXm2kd26V6rDZs+9q78DR2C9Eu/+EO0Z4KURScsGpcAe0fG/apcUnXjdsVG47
BEztuFwjA0s/x5B1Tj1PqGmD+ED+bObJtn20GFGopCp+mo8C3jrl44gT9wI2Bk9o
AE/aXvAQ4scDl4KNj5wsHSm6zUpPhrk2PUClk/sOzZRtNsafEBltjoZoDpcF/QCd
0FIUY7ytFN4oHfQNDsrRp3hkdkPtNLkEn8oWzZka4oMVVzglmwrEPXTjXUsZpPj9
meuSVYL+9NGqrNzn9URkO6gr0F/Jb5ZQ93ekPkg0jfPr6L+UqgMKqXWfCy/1jM2y
JsyFQhONHPFMphnKYZBnQCtAtTEz39AAdDoQ9tHn4uoPRI8mRip39WaKbqD9vMi1
NU1gn5zUd9IDqmjhhANhkjtygO+uduPcQ7pFt7MGQW26XvPnCMuRx/OFXdmkkZsq
Bb57mFbQI6o5BC9VsjbajT+gDc6IHyio1dBzGZpGoEszU7DDpHM2TYczv47Gg1J0
+MZpF0/o4okl38ET2FzKFrA7MX4uZqQSoE8dxoYJaI9QwrYrJXxlm2EiKoCh9hao
6rfwry1fq/9Ya+1dWHjFSHmonTX6Z0TfApEx/GSqjr6aCSIhi3Tg7JSdMTfT6Ia3
Eyt/rRZzQ9cDvuNo+GQE6bAatIdDRyk25oFWfLJ9YXS5Mbmbk3yQbT3zbAUHRUax
jTFsfGEstFqjOfYfteYApFjvwZPtVPLRl3Ayrp0VJxn2MMityWU+J7xUBy326qxz
qgZeaSedKKddAiI1oPJAq9mKjpQlEJuJuMGaphAVx72FZ6QKAXt7oFEIr1bPZDr2
xoHbyLN5MpuyqUfPlCQVYJ6C5fpejp1lvyE7Lm8tE5bHxbxjKLWmeH3cAMHAptwL
zQE/P0xs2c0r/Uk8wtnyFxX+OL6GxjQCSyRsunXcDYKJvhe0nDGZgHX6KQSRHbvN
BYxD+sYMDPP4awhQbfCOW/unBWViHlvf6/1OA2dsleBFl1cMi+GF4GYXqUa1EVoZ
QsINPM0mABBd+Lir1dJOZJoPvPS6HylExgvqCZeqzPICRIVYrkskze+xN9GOVK0y
2+u34KH8DozL9n5GNyKk6ZZlE7A55tF9R9kdjgndldjMcbjjAT5q3D15PLkMMZ7y
3GYKcLI3Pwo5a0ibkI7k/ZAvv3n9UpH7gPReMd3XgeczUBXmpuFagayC0JDXJ1kO
7fIBdIZ601MsqbJsNc67Jj7b36FwPpZU/n+O+NT1Ftpy1dc362Mzr5OljdA8mGv0
I+SIvpz9MIRfgmAAR03LQRxmaiZS1WYm5i9AGeS6jUA8mWRsULGHnJHw6qS3RNCp
wxM/1hyqrCHtJY+Bm/wjJzeuw5I5RN3qaGmhZWDrhj+xoapmDp6N0q7dcDJNgCXd
zWT7Mkip1mcKUwFBFjFsIJ8iJMi2mQDov8uRxc35uUr7MaI2Qv0wJ/wJA3EqDGij
lExOYssm4XsBHuQBihvb1l77VQsNmWx4Hu6n8Tz+r9GtfrGLP8UhlN51/wU3rX5Q
Hh+A9Qpb3PjJRbgTxHcpD5LolKBe7oG901W7sRpBqVa9z4TR9Lh+anONjt0N0MMe
c7NUn7rlSVk7GDWHknu9P48a1v01OFUVmCizpJvwzH1WE3t5L3mbDQILdcwzTCrC
NnKzPBVQ6jRgzoGPP5WLFiH+yp8tg2pRoTlqgQYTOxed0d2eAmEsH4nWkZ+aPlSL
Fm1zVdiDlBqpqNLbBKXUK/Q3jhy/0OmoU9zOqht/6plUjBgjPEhXYaiw2E+ODAWi
xHRkAtYFfKhklIGn7U5DqLPdLkT8EzBh/zotaDy8A2Fcg+zaxZYGRAmI8X5wGuKB
FUPJVLCu60D8P56QReQgi4gRjmTMsCOrshrgTCFIPS5GWRUbPQy1RuFR1KIBZXQx
NZf93xyNMbl9D8822CijmL7l7ej3vuVj+Wvjc6R+3ZnP5Rbu3SV0xQ5EpLW45YWS
Shlwj9mTM6Wzps4Z3Z3fyZYZjhwKQG5WUjk1Hk/rA/1ZfKhZhuEG9jYVjJU4QQ1K
4ynAwVmYYoiZcgpfEOSV88UkQ+IbR7KP1fU+esLVrOVs/pln35omv+72iF+JjZre
g0fIyndPsYJVcFomDkEFi+tzDVbW0tLJIyGuzSJqemv++xKhEAbljf9Q4tFo05Jc
3EqJepBj2QU0XeNito8HsMk2tyPKpnDxp6Ssh4Qo0qiYHNTFcTAAZrZZDI51c5OM
Kxndbu7IXm/5fYqJMIhpQZZUvrkbJipOaNi78FyI5Mt8X+uwJ/tJogNFbVDLSpxt
2zGQF25R2TZhJ60t3Q3MSBdrEbg+ii2KYVpZ4KHwTNcOH7wAo2M2XYWfg7jCCc7q
kNRiNdq/TYOP5VuznM2ubKQzm1+nMEMqz0tBVNhEvPKHJk7RKpXWJWAZtMfvIHHC
rAfPgq8Kfj2r2tv3vLXvg1YXdaWmq40znxVWEwPYBWPmmh3HEizNoOfNhyfrLH39
eXiEUVPZyVg7sY7rFdgE/KsoDfzh/hW9GtUGkFsFeYONxwsaiLDzr+H5iQCOmIjw
PjhCuSm2TwImS37zvcF1C+QV18QlRtDtG0p/Ia13Sa1aT292E1Iz1PPasITzyLX2
m+YKrieHw81Ot7NtDUJlMDa9DPgnyjreGOVEh31a6UmAJfsnpYdN6dBa9AZ8bdxq
D2CdO63aIdgTi/zuItI3bTXXBou5S2o5Sj5oCXYsSIXm/YshSd8P10DNg8veLBMY
npcfvcmgXOX7XYGRUXR/c8Eklll2F2Llvj6I+CEpbkwBHCcu49hL+6lTAl0f0945
a7nK0KwQaLgR+sQuDSV8qoJSoxJQN+TQmB1PTiBE8cqQG+yVhX2EM+Wvvl4mIfYu
Lu4yOsDz0ztMzpXV0KXzzkVNg0jh5Hu4CTOvVFl/CidG0//6yLcvitNIRlDbYGgW
62Gk0N33EgO3Cu8c0roJZu2ToFWroWuyxD/IxFY8fWckfiSAfcQIWeYlV5W6DC+Q
gQ9jbJUvWEwGAgkS4TpzfYBIno17lbMYmB4icLORtWqW9LeuKDrN3Bwm1UBPYt/f
pfmW/gU2V6CMP3li/yiUTJeksXVHBuar+1PAMzSZNvqRKZlw7VHH4PwzvHNDoopc
+9m/xaJtQxYq2MsUeWxuiU3ClAa3x17j6ZGlmpYm7i3KToRxNQiGn0CNBVwmqoGd
D2OpaQlubiJ3scpCRqlnjLvPI4FMSjhAP6aqda+FcD9lSwJ2fpatw96Rj5XwF8Af
S6GOmk1v75maABTLkQzWApO5sfzdJObsiV1Gy0xUvLQr9oW239WnVFA6fqZvdkXK
z4ke4qCNSS/hRStC3Rx2PX0yxI95e5SGwCEpWeCd3fVIHk5OayP5Pwy9Lw7OQ6q4
4H95+w85Sp6G1kpR7h/xYYYzJzVnCu80bgRC86BdJq8aE1iXAyJ567fXjCpCCWqf
5meybnRHz2DCRnCLYINoSkNe3gYInjsyjWcu68EqXxrKMJM5BPtucF3PImPEmJNN
h7a4FlsH4KacPp8HadOCSJxBvOK7iOsEus6/70CWHfUNwCm+mgWf2XH+7iI+5VNg
gucY57ZhV0pzXRMWA0qkB2W+tVKN6H+0ZFPFDKXqPkIMBz90kJaS9jpHg+XaI3f9
fYNSMf+YqrDLJNiRAm2YktwqFKfQXnM/kfRSaMcplhLRxxSwcmD48osoyFpfcgrA
Chbq7PxzQH0mciBFU/ku9Jm8B5cavmR2k7Ajh4/W1UAzoWCOwm2KfsEqyq1GUQ61
TC2B9qrD+1KRGRhBK/womDn03O0zS65ox1ngdms1DkjVLDnBc+oPevAGLSrX2Kh3
7uCz+P+Ob056Un3SocT9OqLeh0GF0/PFUCzG0bg7yVMaqf3Dgce2S4ZPKaIRUDQT
OB3LI+dpNCXnwgCrJCSZcylfsKMkB3dfavz/wU4m091AsEJtPt5O3ukaH7X211sb
q1EBLAQDu8IDuWxLUFcZd9AXcs5mv0wfl4xjzwv+PRL9rK6hNWRCV6LG+w96FNqG
VXBXWaVQvCuvWQV6GpvBHD+np+Se8Ggrk2WD9vD4llQHJuqVN8FaBRoglYJ/jnoT
MrfILz7nikorFs6hr61Afjcttky1wi6uXuHnKmZQcJY9DQbmoUxWxNvy31Xpr45s
b2AiLJewEKVJmZMVdyfnZ3vLhNo1WRpzlG47cr+GomyusbOjd/PiB0nz4JuWH4Fc
t14WFPDceYX+4lGic4wbKvoOsU9827ePv1Uwv1kiSTYNSFQncfm6Bha4dUWPOkPU
PyxoCg4OLX8kONRNmuFeNQPFfULfZtFJ6QVJJH0BesVsuq95C5SHNBaCDWv8aeWc
mcF3FXKXWnRDSEF16Dzeq1DP2VkgIfyqfvz/9rReAp6pJm9rS8Pm9K0bq7wr6C2g
r2x2ycxuLkNaMLaWilK6j4NPBZaazt7pMN1cc2ocTkawHhPNidImxJYs5v4YfXWR
zpq8Eze92C9P2v0F2lFof96Ojs4DbHcidRkdBaihmxQiIUrArb7BMdstayOaOKU9
vUwf2BjVTw5rnEqEtpUlTogRdzETK2zUf1F+s163dZXToIXRP716xYB1tT+KaQI+
Qg4PdQDezwwqUXD2fyS9tMN49hR6QyDz+5iDOgYmXEppxLAplg06l5T33Yn39sEx
JXsMfDqtyihzhbAzeLVt9tnqQU0sZCYFKkljLU996zKu8G22VjGhNxBr2LBdAFpy
OPDcTKgJIxEYoTgxEwSUfbmIySbgIseXJAKV8oq7dq3xVlk69OB0a8BNAf6NFFDk
81ZcOuMkxArYyS1O2ENNo5+ae9VJMd+fK0A2Pob/aBAk7+bImH88GC3uKtGVqTHJ
Xb+Wr8veZvqQPJ700Pg3g7Ud4FCE4WpEvQHzdM6i7334pNyD0XlV/X6w9SwL50HK
gSmFy3XmYpVs+vEg8SFkEnunEt5tYfSmBGVwq5p+RQKmJDh/mVn4iUtiqqM6Whwh
sL4DnxwLhkFynSa1gDLbdHgTuN4WcEvnzuAFfEN4yFCB7XYe+RXdP8Gacv5A9DYE
LVmJL+kjp7Y1NfOoPWv+OHZNVRPzR9AoyDrPfpbOYkA6C3jYPW8LiZxz3lBWwR4k
VfNGeUEQFf8TR3snkGUBhnIPVXKZ0ppsXxCmkom1dq9BwPtzKRN1ZIsmgB9gdbQo
6Tzm2LlzRBymgtm9XElv8ad5CQcSPwpY71OwtiI/Fg0ZDKjRw+R5aSdIKK4auxVy
eMLdk+q7QU2XcLk6EqBN4V+2m8NDDHy2dLuZD4uhtyn9ijwMcxJJeYhxCuZRvgUt
YTrmxFpjw59AMsdTFALhmKdzTWPaWJXsZ09tubWWu36aLSwVudy+Vzt6Q2J3ZVOB
TOc4Zi0QULqAAyVEnF8QgIcarz2700x1FJd2xfemsdvyoFDUWLbMfq9GIDhVJwC0
bcT8oIdDR8HzQTxGSLfEeZv4MUpTG5qh1WiHnrRBssleHpeFRMgDK7SKxEiT8m//
k3yFSq8HgAkf4rxq6BeIu5AHvEumBkbYNJpbDBT2hVRYIn7iRYn5PrTGzKN5j32I
s0LOIWydPhQzkBlwSBGMTma2Ej/pvA5mFVrxX0U2T0tUB0KRyKbmx6PngCVELQ3Z
scCyhhlUQidxl2t7jurmUHQmtgUSw08WzJpBcZO8AYvPkHoZX8ypUE1CRX+YT8hy
eDfxQmHYEDB102PaIghC+A6j6ukD0n3R6PCJgrmGC0ngRWrXj77gaEvcsuuB+4Oe
gzkHXu7AbAj0/XBuuA2EzHVkPe0ilPNZryvOYh5u0nMWs/Tv+gM+zoAX4CDXnXiX
sKHUntdxTmklrtYWAG/PLd33ERVNiPE4OkXYjQklzmBfk98uNsQgvcmQdzsA5m/I
mITZl9FV+QgZ/Zj6sZhCiMkYricRZ18USO5XzWpLW8qdKz+E2flBCWs6idiGGMaT
/1Z7kycKYrmUgKFOP7ZBkYGfUdSv8wJR2uYErTnui1F511UWw0shcY7tTA+/eywk
0/aPVHuNAHRv332wZOh1ufV5AmB/S2sKV7Xq/Vdp4ogeYhfLW5ns1XwvCzJNkdH9
3web+UkUQYr0MbeoqSqips57ul5UXbivIbNCIz8mj0bVRi9xus4Tz9ftERYIDZ7l
YaaKvTIc0Oqn8MR/f1Xaa7JzYuZZSI8EXZEbd8HqDC1FniJDrpAP5i7dZcsasfWk
so1WA+GCtzm+2qx/+pnQkziVo+Yl9f1EayTsWoMvr8Z/TLPgnsYRZeYVlRD8GYye
PR6mGnseIJeiwy0VGuB5qy3MgxoJKp9MZXXhdJ0I85aC4k70GQIFNtPJo2NSbGzm
w8/CI9OQMlTfo4xrAQJ8Q6BVw4pn9VgPGhKEkDORFQzccUW+hsaFOc308cpwf4It
dwCZdmaEjY6uVzUrnmLt7SFRuszKLmVn6KYAEIny9reeT99YkaBtnSp74Rp9qI8A
6Iry78N83GNYXN+/X3wiD+Ecifh7RvNlqeN5MfgdFtB/VVnI4XFuRzi81917tv8L
96zck4uXryQCou4CPNdvhsoGgcrs0B2w5sIokkn9VTfRcBFsoX9KVwYjlunYq149
rv+LIKZe9csoD/7fXD5dKpjSUwmcDAGXHPB6hoBgV1bLwL/FcNO4lXB1U2MYd3rM
JOksTnpwL7HDpdJjqlrmxIunHaNrc9sOURA/0jjVzT/iouGJogxpDaOtB3q2wJBw
mC7SpmcFIJmpJN7hhcGU0dxOn5w5l7ttCbav/O/TFG5HT+prwtUFfuYVesYqcJWc
2P7W61GkBix/7nmXsuytzphS4fE6SqzKi/jBan6zMRwKQ03v8tf/V9aPsoIL66vg
HtGOyErTNl1v68TQ0or5pW94kedkLj6SMPxOprumIK03tiRqIqXzM/z9EAYJOReP
2/zKuJtIu90i9FQX+fwGUv1xJYLSSfaTJdZQdEI3G8qv9hGw31btRev4+qTMZ25i
ZAdbhJgJhp/Cs7uj9DfWgteZxPdWWZS2V8m5L1cgOydtbqJyuEdUVDIhtT9cekso
KOUOitXdEohLxCnaKWqCdhXicA7QI1j4ubWplrv/nDw/GXnDu8svEQtpdGl48yBq
B0nx13Yg8vldBNJ6XPWoAarWlik/dmpG+6QfRL9R5FVhEQz3b4QVo6uX6ZFCclm0
VKRSblccTJaigZKaY9yx7fi+nNtvJ5LhAfTOZGOx1z9WDc/YM1/CuImEeY4Llj1a
4AdZMN57XZDyL7DSdVWZvldNMPiqn+wy99cpA7iarr4Tz/qYKxV0pEthLdlQllEw
Pa6aA/h+211BArgeGPS3Xvo32bc5TXSVnbK7AIONsDEjb3ryLe0MxQGFL5mrTRSh
Z+seIy+E4XvN2TvOquXSemOnrJkEvJYKAroWgD7hWQiCdZyztUtUmkTiO6rajn8V
pjqABo3hQZnwhDWQYZElNNBFLExDWoMHo5sq/tLWVVDEmbAInp9cMF/mLs8G4Kii
eS0LvQiqcVGx1TL//rftiDyNzht+P2pOY//prRoNuCMbNoZ42sq+4A72JHtjguos
iDiqpNavN9QzvMZILZS6iXTwJuAXe8FRlxJtyYGG3truxBHt1uA3AaT/TUdGq78k
9i9q4pm0mHmCjETPPW3g7ItMm5MxbSdIBqlnSbh5dJc77ok/zMNU9Oq+Brxu4csd
q9xPQ5dP/fnKAoPvWvUoDGbGDTlNxmBhm6nQFvnNIt3L9zPjCbRPzPbvNvQBKaas
PGjSK1QYap70ZCmZiD7fLc34ObEqygELgZ9q4DKSfxr8ISIxlqIwOXW9eFhOeA+Q
fXNjDIYLUWHnwk9UWo0Vi7mPFZ7iCBu8UNkCmoF4G3poC3/+yNANs25TyF2i1sU6
Od0p70Q6FFP98iCg2bm0wzR3zVNXYZZ14D0UyBMFY+pbBOCvP1NpnzIdxybtzW7C
bVYgirNqXOSAXYhKCO7UwkKwwoy+o2ItqugR3jj1/imlZ9NfBZEhugBVkxFNmemn
v5YDgrRZCqCwPqF2GU42f7zaaeEN9N2/xMRhDTZX4kJcAK2DlXQukP3chRH2oSgl
tLLPG23vyXdrSJzhbzRu64QGkE4IiyJo85mWkL8djNGPNpQ9erSEBG10rIRgizWV
/bybNzBS02mbcyBABJDnZN6ZEUOTnV+yGYr0N6ttQcyrKuDzYoWSPERQtZ3CZWpZ
P98rZM5R0TVuTs7vPUBOD59NEXQHo28k1jNM8P8lOu07U+JdOow01zmhN5W2jOHu
cJbUEgtUwZXg/nrrVaRjcenizUqHskV4bMYnzdVrjTG+rDDcl8vaolteLDvNQeVZ
4dXyORWOlRVTzkHunjvnLsG1/eCWk3ed/ppiEnd+YiS65aUfqCWJI44rdP5Ob8rm
2WtEfVweU3gddEoJY7Al20c7HQJ28JRpdrumX7LehpgNb7PN92gjXjHhEQz4V5CE
Sd3phTK9m2SyBIRwMojHBWFIDyXGwu/oqUtx3c6Vmw0EJuIWflBPgxYjjtAEUIYZ
kR7sWpWYPpMiAo0LTi9xIU8FqGR2Yb75h2y2gePhaT16z73ArsNGLdPrZCZ9GKSy
z4PsivWLCw8AxMSE6f2ii2HmzT5TeFFBQ+JAU0XSyTgC2LaTpUfDn+bpYXVsEAT3
oWVo2+Pq7HUKNK8T9FTz4Cj9HKNdx5Y2tzdU1q71NxkIQzTp7UwBpb7ISd7Ap7Iv
ILTuEcjMPi7NWvISqoarmubm0XbrjUPxFTAToOsN3wbszfPIFrH1S2IMbOz5JXny
lAA8VwuY1kyDxAIoNVY8asJ7qIsHgV0JxAg6X9uUK/EqKOcdTYWl2JNIQ3vti7XU
5TqFkJ2yViAV36+zRrOmsoC9lXGHCIOfsidmpf3f9ezb5rQw82FNw0wzGI9rx0cq
Ny21Z3nfvYYaIm2OcuKnxX5oG6iDEknDOmV/oPcIVlOLGEmVCPuGERhYIUS1Mb92
aWn7P8/KHBt+v0+WpKt4rqGTeWIeNw/NqABX6Pdo1frZqXAxk3Oa2TWLOcTljpBm
CfU4k9E31PitaKZPdpJWgvnX+/fjXMC/nBNr3flNXz+Wec+6Lo0TohdfmHcjJoCT
Q0O5N0W1tRKKtFqBJUfM/C8rtNmrhMvFdgQLUzx+fTwrKPkLv0vJ4yun1n8Kg9fW
QZ0XM4U21/qkGbF2eATAltDH7yGP3yDJ/FSczm7XlQ3VMH4+MWN4AxaLVBfXJWrs
9BJN8n1yABmZPEOTpzlq/Y79bb5PrC/St2gZlqDJ8SEtqaGatbwKCuBGMdRebi6B
fq5nCLvqo79k0WgxNMf0++foSw4ier9PTw7NX+4trQQWrf/09clo4e8S9amkdYoE
AHRuM8NPIIGUNsAvONxCUsOERdAUycHr5tVQxtzsIdfTlrQ/+jY7Y4EQKpEQ4vze
iCtW40XfHl8UVYRs0jdlNeDAUQ8WRYud+jBeVvyMZv/5jj1Q1BUxslNtX341Z1XQ
18yyi3IpR64KaZhiNhzQNFk5YHMGQngkibwl8nKw0BjlmSnmer01QZp6s0vF3g6I
Rx4rwiab6q1m71EnMJmi+fcyi4jzvcKabIbHzgcyglR+HJCfFWLllLhYgVvsiKzE
wxRWbJFzod9e9W1wZLXjLD/iRFPX9cQB0w9tHMgFVzobkOpCcv4+CZ3MOY38vWlD
nAVyQL2T4qSy5DcDpPjowHmJVrDa39+v0uyN4KS0dvZMfWDEuyBae97Lr5TgQgYD
w7KGJJHCWfQmcxpwZMa/MhjpKqnd9coTJ0XtvV3qPgZffsqyx8SnLLrxbg+aRcfY
NXF3zwQADvXB+Z+JPUiEcXt2Dh3QgGNUkN6LtDLJrsPHGUqBoKVN1ui9U+SjpSqc
7LYB+u6JyivvAx5vXtjRsoH+a4qaZYudqYhM2GvZoT1s0oOXBAscHcMbjVH8keD7
069HDx3ucYGkOqkRKic/rCS3ls9hwI+QrkqcO+RQrYJor6Cx73lo0PkmcMgxqtqp
xuIynsasXjgxg5emaimlNQqDok199d/xdx+7KFb99WkveYH1RVi4U/+ycjq+5RKp
WohtW/9BbKm1eKzBSv4eIe49b5KqwW3AWOC1ki6T4V+dd8wIVFQUkvWKaz6+Gzx2
Q0CRIV4O+GsRyHhaEkIJCaqEnBcPmSeh9uCyarMh0iJt9pHcrNHt8P8MNphCLvEw
Zkx7ySnnQWI8Wo9bvyMj8KflsqPu9OOKfTE1+CvISdZGm+nwxkAHls9rgjfPEsQY
SNl5RX7W2CID9HRH7YS5OnWZKXKMLxsxlAlwIkceT0YdPGjJ7OTEpcGm522q+fkT
MphwvE2CP42HjRsB76UyIUb2h3JGouRWSd7dnJBUUc1PzuzZBuGyqasQTJfnBHx5
l7mi4fFK6it4V4uNKUbTmShkCipuqyitchaCYYs8xWazFysY7/HKEnaPrGQr5ZOi
3xd7YRDKWbUPthF+NMbde6az0/O005PEjA/PLuMRbHibaXSxO0v4fzz8P4t8sgPL
nWuJjl3YMvWZgaZezDuzgvarTDKWTSavXqH1ZShtQEj0X6++KlQcEvg6NpjMAlcw
5ksnChdThxH5rxWjEq/aaRwIZqAnpc3Z3tWl1QQRIa/fGnF5SmtS0yQ9OZyS5Mnx
21iM5yT9ASD8UeLidtfkEu7lfNVhqa5ul+YYjj1ffr+c7XdF1g71jiw3lL4QUKZK
JDeA1Yl/XnD96Sb1qSQB+lVKOJFwYJgTEX6zIGCLnb+LP9NaACEgWfjTfM/6j2bP
MxG6WHJp6I20WSXmzOJNOZapXgj1m/KXrOCi8emjxWkB75OrahKiDfID6d7hxUrT
3DdIxFZi815b3PHrvnfDnP0jif5rWG+yhk4KRq5XATRbfnD3GHPQRpMTewUI18BN
/Sh1Ytn+K9kZEDqWJvy4kD5SmSoPxoHESsyZ7zGLna7Q6DtUap9o3viPzt4vzKm+
7FKBfBmqXHXjeeUWGK84TMICcjATdrGViyM8+UPkuMXWiMzBNusT9LpTBnZQZeVU
WAO4bFfTwybeXR4BOsF2PbADtanQKh0++zBqRwPPMRprBwifd8IunnPT6oshnhRM
ON79xW+rPZOinJnIdt48T8Z8ZqtRn+fH9dunJgch/ZY1xKw9JajZECJhx6B7jMOv
sT0ZWVu8TS33tWHsj5AbUkpYqmIPOepRs+q2UybL2iOyKU+MLEKyWsKov+/uY48x
UHoH/KnnyOYGH8Tf1SQBNMzRXWiVW5k2aZe1qYtZ79V6O9gB0LcqYyedthHryF34
4xkxskY3TGxGT0V0mjXs+TPc1LjayhdTz3RT9rOubjovq8ECjAs3O/VhTuBfBGK0
cE1Hzj346Orh+zszdH2iwrLG21HXjRoS1B1xlIw+e7PZErwhfkA+d+k3A9Jg4x6y
RfrjMckNaKKKV0jQZ2A47IAhihLzdAh6yMXoK3La7WBV5ucLoSMSE918ghJzt2DZ
pHKYxhP9bIfzzTnjnbLoPDEW4byZicdoB97ssEaBFf9n4GQc3Kh54YSD62zVfOys
FxiwLN0TSyBjuIC9lm663rJfnAwtv4j/NME4JSrNTBcTfDLZm889r7IVMOvqVn5i
Zr3TD8JcP2QPIHw4RY2U1sTB2wDCvItBimYuytRhr2XcuhYXbNfxV5t2e6GlF2EN
MUMieXlplkjySdPjt6fwiEe3sz9QHJSsHvw77zVKv9TqES/nD2yyVxP6Q+jtUYz2
`pragma protect end_protected
