// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
kCOBywyAE4q3sAZE/bhCSL+pMUegF4hPLuQD1bRLbc8JMYtYt+7UZfUsSlWwIe/4/Q4udGxYbuTt
7eyFZ3eXBRX/w6cCUHF8s8AYHMN90p4OMep+z46xIKVRs5PCTuHP5S0vRSfLBV9Sc8HFP8kDc0G3
1lLnPkoB8unfuggCstm7233ccn9yVXToYfFpwEoHZ7/GhJewXa3hZL4u10wXpVlPmA1zsopZ5oEl
VZKivpHB0QpixENtifDvYnb5x22ZfZgV8tA6DWuzMUNyu3LVWzNDxDYj8wwuf0kSU7yEnkk7EKYd
BRsJUTF9Zlmt7pRZqb2RTxPX2gHzaX1ry4FHXw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
AsnjZ60avhmjN4CE0vRqyidYEeNazGfXja9xpf9wEivqJv5T4+Po0UFIgI2Xwi4RCjTEKIeMlIHd
zg0t0Zgcg+/N+eN3lJRAu7adC2QNOTaOxlR4yeaO0qRPbCBpVUiTEuSfQsaOvF0q5FZwpAipsWkY
k/uAuVOrwobT22zz6oxHiWdchngT5yTiva/ofHKB6A/43zk+ecoDrJEyQ0O7MtZKWyXNRkTVw1Nf
qLIlsKiFhBOGOk7o+8326Wr0ol9xz5yCyBq8FY3Dh89z38m/Ka7j1lG9qjDY6eBRL0y9W5SyUwnR
dd+rr/+Y4HNUUwrCjqpUGNuGbTkt2fHYbj8CisG27j+cF/4U8IDYdxYHeQmWgf+ULcif3ffZZMBT
Lp0PREw9xYSxXopvNpaHM4uZC/a6SjO6rGLw7YinIKtHoJNu7TwmSpHcQKbFI49PR8YJNklEEFnF
V8t9vpCT076nBxmKK474DKYJ/SZnQGKbsN9ROKuXJwnqcFX3yTp8aFW/nbeDZ1epsDW4BncmVeKF
NEo6VSGYfH1XYhNdDmhqsiYXqNVpSlgUiaRVH+PF/5/BnOZWRGL09VzBUZLc14tam5qd0K8Tr1Oy
grfE9NAq8k/k3QmAJBLOz1r+YY85SbCYEcAXQynBPjvs0CQtuWQnUeywXdIdGmWS2vw6dpb0TZkp
eQ2c0ZEJhvC1+qO9Xs5Bn2EycRo8LE8ipYLa8jO6FlUpABLP0HdtaUgU2mv2pP3IvtCckbzvyo/J
AXPG9T4WaA9DovzyYcwzeXwreIaN6OIig2lVLWm6B2uh+64RDWWDegwzD+Mr4o/dadIoDJto8xC4
C8W/XfWxBV9OMjGHSZSeRqJMvocehhPwiyjqN8pII98EkKL5ejB3O/IbM7srVvco+hjvC6vEf9iZ
MTsX9RDn50ThKjsuD2GFj2ehMVH5PIk3x0cLPfBf1GWobrVIpCVHoW0d9g2uL01F3SljeeRHpF8J
mnITy7vt63p12HqnJb5Vcfdjudz18vV3V94/FJO/TF/DAlDStAwrFkIdljeRgyTBd49+9zxrQWkX
Kd0XKSS+j0HzLUyRSCtnP+I4yQ+0PEgL2mYEg3+a6/3txC/7ypwd/+cGNXJlZDH/z6zie8JkLn2p
216q+vr/6C17chZk6z/IV+5Q0FTWPmfCPA8nKp+2jk0KkodXe50FgwdDIt1YJD6zjDPfY6i2Qwpg
AdPxXDIDbBqt3XolYyxTk7NAj9XXIgnG8hmrVWpVHbkznincIJCZNsO4ATdBsMIJjXvLQKFtm8yY
8QdGMgu1WlY1I2uoNxCPrKX7bHXqMbFarHBeV9mpe4cWSR0iRUHAwtiZqm9Ji4/1ubIbnd/sDFvh
AvX0dvxd/B43446qodGrPn0J8DB5Il7U/0SnSCZYYGo9fI1ZeXZA9ZU7NMHo74aKOAuA9/XtpTsw
PT/a9bYsrHgH52oQ+aMLt9Z2dFusUSsVf5mYALHQoGXVbKbfrPYzfjsm4ccuaXPIiIqGPMyafeU1
o8X4wWxWMTZFePp3VytcsjvIhotoHVDWVkZZAZmqQX+A8uA7sLPtXJUs2d2ZD6U8vZHE0U5j5ias
+sIlZdQj7juzF4Nn40PTik3sWqqjRUJQ01tI1GKtE86ceK7q/iWJeqd0rEzo0Exlr/upA03yiuo9
ObekaOpumhpANjUYPEK7jvA9YEwBN7X12WrW/8VeU0o/YsZtpy7McoBV22Ve3dLNclv4SVJFUBQV
g/V7W9AvY99i0Hyw8lIwYIYQ4Y41AG8GI49nL/CRwcPTsfezQNr1QE3l6mWSuxqW4hH5HKGLsrYf
m4luOJdH4tYcu6vZ54X7F2Qq6k2Ag4RRJYJ4CYMKzc/IUlckRz2r0Lks7PkIHXCUe3IA6n3SY1jm
849izUoZKSzOj7ABinYkVK6KbcttyivPzbA9EsC+NeKQ3GX7RFnmFLSMRaOdCijXsUMiHGCrgpzp
ELX3/hnjvPS8ea1UYN2CwwivKfL0NWVeJ4RqHenDmtxVpMDTrPtnleQmyxVyOkagzzyaDOyqB99y
jcQnQzng0G/PfAXuYqg+yosvr/N4mvp/jxls4/0YNL66ZJrC3+uF0BKGViUrf8sAqA+VEHFWh0YI
wSKD0iiEGV1auSkzsRyy67+RUwmH9ewRIMWZEwwTmJzMt79lpeHvIvXqXpy9duiSiVVM2vd7ALXl
mqAiPk1Aumtn6GfEmQ3haMsmNRG6XEVkmCCYbDS2j5BKKn8AIo/Y6uzrpBrVP27E46oOQt4ZIIuN
tqvoiuLCMPD488+S5I1yYk2TQzxy6FCUsfXTe+ligNxFHUdHyHt0Rdykbi5JuBxmBduJXBMGmTSy
d7riIzpVSr9OFKgACZKrtYi5Pkue7zqa3REk4cMuxB7fFB1wh+MlDmtNU3AUSzAncZ49y6FaeArv
8x490SRstOkgFBbzANahlFxdpaQoPRGjHQ1ps5jYiu3gl/HANbuovIxRDeicyh6iGb/LPn4HBkQL
gsOUcHPDUu+2uKxRWD4k+OPdntunhGFNUoF0iIkNx4aa0cCfBnP8L4n4SXhElIV03pwUZRuHUeU1
y0wdRk/8FI9bzWeS0GocJmTA8aQktsovppRtOUZVCfn88066rSVfhJYq9z0eTPR8m43QRXHzOXA6
3Q7Bfa8yPlOM3nFcO94rSKT9lx7hA62LroyaeeBNcNC4TDQ95ssHjMY+Is4Muv7XPQ33cwEdVfpa
zc7M1Iye8Adq7QFcxZxt4MygnWtvOUTIFcvFHRzEPRTnaexQ6pHULvPxR8g6s60fA4st1NAf5do4
UzrBVxSqib5Mq7I2iMSrWfxDDyi588RHdkvA2FRLqa6fjcdepuwtt/KUEYTvnFujd3O8DFsiO6L+
++DLEbmlchb/hpxHoD5VyuMlh9Dr6PTPe4UhFcd4o5PYyAI6yWhxzFUwbiYqdUDdvHBkekAtW6L/
A4hb1p92xPunjAjC7I0eBcCDKiHq7pimUN4zBXFcjSMPk8b9AEItyVu4oq+eFwYU9H6YaDM/zYRf
wof169rA4Wvpq9DxD5ifL01E+k5ntExH207UUoNHJS2YT5jZ/orOakbNivOrdfmKGkaiqi5M8ey0
BkB/5DBFrboOba9SLzizDhYTSd55LkneTnzSvIYMfSEa9Mi1WEDcKcBp5+vN2N7pAi8EUBeRmJQn
C4/df8D1/UI74PV0XMB7wpPxAijMxdVH9GF+bS29PQnAgrnwxkp8mLeB/pCpfSDfsHoaUPA+txLe
hxzwW2e1mMgotG1B0BMJcaJnmK2rDX0MiqyHCw5rtB2CUCO1PX/mMtRRfUYMxNLLfh7Gny5f/0uw
ruzdt2N53gLS6uJyLx+uFZnrWP0Vy3RnAltaHpX2GgX2V7ZpNC32PaZ/IDamIvEiDfHAvbD6wW7C
kJzRYesE1IT29cXkVD4HeKgCBPJcbjoG0kRr7q/aArjkWhUq/RI+iTUVA9xZS3A/qxE/smJmEko1
j9iwmode8fwcuhQXbFS6SHkLjop0Domuob3wCZ4DBSJveiTa+6yExNlFU9KTaME9KVI4kefRRpGN
zXtCnxqBa2qERe9jTXxu1PGYj39tlDMpP8TNSY3usQe91H8u9DppJprJsccX13Qg+ZfEzTCQnxUv
fp+IADeUXQGQN/TiDH6kvlgD1UWYr1Mpzt4EFXWNrA2GWFnIUl1LWI3D+b159EGIks2l3UZAdN29
N8AQyXG+bRavf1SdzKFZXpjNLpIz0AWagMbyWdLWO+8s7GUmenIvsIGxh7ZiGcX+CPwllcjEJ5P3
RGVc17e0dH+lV/yI/RBxarSLNWHt6Q7n7fwULbxyKNajZrZjz1x8U0U5X2NCVZciVcnDL4viv9t/
xOMQKTfil+b5LirotGWAwYR1wUf+Vs4Z2HMbOQlBUcmc49qj/Guz9OroJTyLyacQi7JxWBLesMi1
+sA8CEnYE+EgAAEIhqAdMj+OgtD3slTTi7bV4V0JXQ3vjiQwcqAPowuDzYGUrHENuq1wW5GzLDEW
7Ne1rWtmxd5gT0+pIqALcQFDd9fStXs9vqq25elyv8T+ozCC8O0kwkiAmKH1QQsLwQQPNhV8Knnw
E98zqMbPS4BFSXR2P13wfuDhBe0FiO+Yf/JhqgXV9LUOi0UPgPk9YmA+rJZhJ0fgWlwPpgtFYk11
p5hJZBcVBsMdQUDYNJdONHQJqTPmE5q5Gi1TWeMDJb0JT3VZVSb/0dhISQL7dX3s42d50CPti769
2kKU54WDJjsc8ku4w47e305B1siWIaRTmT8NGKgtxXMoZGHI9TC+/I2fesK3jryPzk42b4PDAxH9
KRe+MDHnvd86rGBsU8tifw4sa9EuRMAftnVVwpeCJe9NtetcSxy0roEtsct3rx6kFTOWVHNPy/mU
wTQY5nX7thg/bIACudj6ONQVOaxc4PgYD+1JJg3axgdVzAC5QkowsK4IYae77I8CfraOEEIsns6V
ZAXsnpx0JF0OeoXqBjkl/NZqNR6BFJndAg0Aay0FijSGC1qyAwaY1M6zplcGncQRjb5S6ZWlDIM8
cEt0lTqfCUg7Sx+P57JTepaJM1TcIrxJBwoMRuuSDSdr4zZMn8qTIDtawQ9IxJXZNGmiSR7CqoNM
v6/HRzhvoVmCZ+BANj7Vlk5SIcnno9m/Fucm52DrPtCfCJwxmFFfbUbQ0qnaGjXNvwprqj57yQ29
bNXtIhORCq8tdyNrMtUpw20GY3XhrTfw+NJ+00x8AuKsokCAUPnv0HldzuCygk+E4l02mZAeJ0sM
nayfO2QgpRaN5adbqsOyuQkDwEiJfIK3SCqkPt3FRv+8ar4x0sulzchFhFkjvTJECXFrczowmulD
o26lUr7bK0/VXO5MjN1e8berryG2NPVRBuK20O9mSMLcgtivOHYw5asYrIZFOMGG3nc+4spGvzF2
F/AW9ezgr8XWlmFfDrPLhCrtUnLvwjvBcVbiFrLTYm3L0Y9JImJ6de8eOfJ608UZmRPWiJ88blXO
1JGYaXLItZiJjlG+iOtP2Dw1LNTyWC102ZesPTIMRgAzY3due5kW8AEwraT7C3soh4ha5Bwq4dHS
NAW4UyR7wPe34bR8ziiJa72k0GhSgpAxZcBq0PPfO3V/aMUq2JJTJEqCg6JBtpvh3d3ugO6+xx2A
RE7mTxbk6vZA3S7ffLpBD4rk3VPHEt39L6mXA9RPM362Cav47QA8E36KL533j6WaUgqszcC+GD/H
adaDENRE/V8sa6tkOA84ammoEJtLcQINmx+hELKRszECNQIYVS5GvjFBs9l/iEZQMfw6Z64IlpOv
O3kSME+2SfqTri7b/LYAOsdnHy6MtkTC+qi6YFgncO7+B5qfNLMZ0HzXZ7tCkmwzVGiB2u0FTvF9
cJfVOyJBMqeHniuKbhOCAv/S3zJcwQz0i4clRFs3V0hQljCrXC3EZR1o6Ii0dsJPbiQMhW4I+0nn
5IU1IUkfRcyblK33rXIdm+AbCY5nauaw5ywU299cjb3jro2tgbf1l6DpXkz44sJoSG9LLjtIygkN
jSqDofdwvFQNJXK2Cfmin1LLuW5j1UWv7Rw88sUHUP23FYDdjmb6Qm5alEPpgq9rshF3v/e5Z5XC
REn6MzRkDTEKY4G7RSjLXZTBfDqwlWxGFgKVCL8HvXDC/wCHTIinbp34OrSOk+XkC6EYHOQXW6tP
vkA1AeNy5ijpEyvblZh8wpiWRtUXNiY0+8NOVoR7eYYL+J9w88PPZN8oqMAI9BhcNlQRcKvyYmBa
jS8FvM94xrolpZn2AGaSRLx/OyqKJCzJPcJOZDAMrRjYRFQhc8CjU0Mf7mb1AZ5g+9vgvSO+N/TT
GzW35Kf0SAEBFQdFmyfZuRxnmeRZUF4Wdq/ZqjVS7on3321nFgHDlmyI4jjPsz5cdxrkiOZypJvn
6MM8yRbQjrjb0PkSib4iNIBto6H6npm57Iddlvq1zfThyQmgcOG90wpRBVYyeLok4bkU9yZyihYn
J0gdX0dJSXwot8miEXjxCyWNORJF9jCiS4SItblm1vSIe8kuH21z6pHICdmGOzQVlnkTDRLY16fW
1QVaREgRAZgrqUcB8WenOOp3kzxfuA9OU68c6PrUQrsowmqyF7iY+cTpVk3uHUG96K4L+JIRuJB+
FDeSHhIHpJR1j3dBiS9rESM2dWkkmDJHoVUvYEK+FO+v29fI6aSZoVuxrnSyTTrDGPLisNHEBBHb
3kjWJZEw42+qLIX6ckBLPoCR+oEp4w4CBqKpmomX8piTKe2FUgvfN+HdJ+JhiQY2syzimFiEnp+3
8c+EH6wwA7p46VWzuos7soWbuPuqIfscHsB++fAv2zJq3YbbnXmlAvuwvKSot7ZC21A0xzTeA5vO
D8DIgagzlhSiPwvLzHCbuCl1lUDyibmuQ3p9qfhgB9mSSZZOi4Qb9yIJPaSKjgWykpstpjsGZe0E
auXMwIg7qNGdiP9Ds2TWTqEIcnhgEaEw7VCMhE+S3GSv5h9vg1dLAcaTH2ti+HuVgMSkSuiFgMe2
OGyWpSysbxr70HSUaPvLWd6IEGmvqg1s+OZn+sd+VZ1d+bVXk4ptZ1eOsilgIQEbfSEjJx2iddtW
JRuZx7A8TM3hM4Qf68Y0EtmlLymdru1jQIdNTAdlmK8lM2FLBQWLqYVmHGG3GUsH9rzfa9206RsP
srRHYg2D2wyZAxLj0DZITuP+xGLL6VoklDpj6Bi59w1v6ikBXXUqIVoIqaGxcMgoW+VjqYkg/wy7
fVQudQTrQDQm97PkYrKOzWBn8R1bb8sIxRKnldgZjjGpOcUE4t6xMt9KVvLSmWX3MJ4jI2HN+KXh
fpnaTZMcm2fOruzBVuhXGonq8elyUEeC8fWZqoF7s6tZQVAnFsbjblhwcjpx6SnURj/cv/GvqlQ+
M+joULTu9942ZO/vtxTzj9E0T0h2/4Ev08VTOXTh8xS2p+fEU6OMLwPtIkVIT+7zEgD5NSAQUCFO
hjrM+dvTTX9nBRP/ieHjsEaEdsjFCd9J6uwXsI3aw65iOKxkVeVtU54hojOEII2YIuai5JZWyvqi
hd/4u3xG6E3wHogizZb+w2yU6ieYBygr+ncJZR8Frs+p2CvnWTE2WcIQ4VdB8HDWk0O6O31LoetT
BmL5XkzAfKs/7OMvii9Wxjmsj9q449lyvwOkxTHQsaISP0OU5UMI+CcMuiZgi2ttP0Q2+vTQ3JNq
KyWZj6BFSjfmf7iTK2+kIHBu+092dt7smyHWpWDyAvY6yHdOSmgku4Hoz8KtrMXJbI7LmzDhoFid
mndwJVcYo87QWbpOTLWxeTF7h8XgqM1FpAvvseGaSs1x9LjBOfBVZBGhc1c7usmk65j+aKJbk9V5
4CTb/k19j199tnOftjNr7xxa0m42NhPuuavRPUolcoCW5803DVLb65uQ+nRUXIWdvMQXJCMfvwPM
j3NeAGRHKCm3URpHJvTQp+fOTKGnVSz32WBR3CMz+exmcr7gydf2mBjSQfQAOJBGJVdZwrWcbqbC
7LOu5NhRVW9EuhgCANSG+jGlL8aU7CYkxg3M9P7xcfUiPce2RvztqynsR8Hj4O0ZMUhu54oncLR7
iNQw4nahBmjJRLO4nKndmTexmRX+A13bSIOzcdSkFRSHoZeMaPXW2x6eSrnpCNuuANGNGVg7vqNU
Jcz6i/NvmhV8/gPhoUc6LbZIsuWYkKFwrrgZjG9hoKL9AkRkCACfZwGmMEqsidoCaVbPb47FaQEc
0v2XyaepRrtpAM4+j602PRqsRJcmOuvJx1HgIIZa29TF8n8dPpErlpJauOhTNElLLs4eRP8ioWeA
1YwUL9cnqpTkh6XphC/rSEPfAohUYrmhsfDQP4UWoD72tUWLxt3bQRCPiPA3C6mXcI/1vuMh8G+z
3FJdGhvuOP1KadYN1/AxZgWy0YHFRLTDUn1cZroBwX8Fd1QaLNU16Ooh+TD2n+Rgd9hGInmSDmiY
GdZpdJs4oEfI++RUFgY3jaYiSXFQ0eTHaYfMsQSrYHPkR0uP4DBkBf3OdSUQUurXVjVdE6S0z1UB
Q2xhjkkFwqMEIw+4TpDaB2kaVO98g3mtN1WbXpgu7Z2dN5CA0JTnb6nyQIknBzV3f4FPQseE919S
4ZlFBYZB65GJoQnwCgOHXMVp7iO0PPoISRePukbwtBj53SK/fSVEnbG1PndJBmNWHAavRFgI273t
6xTwKZh/lQLoujJ70hGhzNQyytQlu9wGvld2cmkr8YD2G39FulvaWqZHGphZ50h5FOn30wZ7KEYO
5mTTxcxyO2xz3Id+WCgDWPfbf4ah6JrjdZNH+5d39hFqPHoHvHRHVod4ed19AcZK1TFjL7F1AmEn
KhgUfwSkJ9IjpEBaF1nbEcN4+nmU8XsNZtpOMDTQMnEByjisNU+qi+wDRyKGZysqUwXM9JQdZwZM
QhaPOeZ13FezyBQVnLdDHVoZmkXj/955cy45h6H3p+Sk4lDn1Rk5NSy/N9KVJJieB1qJMmMYPxaH
W+8DOUvUljNXTsr+89bUnDWTxsFTL86uPaby+MxJFUoiexqXikZskhLqRE7VW4jeR9rEyx7/9Dly
hryJKYjwfMW3xXVMd2jMmm02n3jhJgdAQk9wQR1hPkG/Edz1+HkvIqeGwMQWUQr4uR3/fjgfZCMy
l5pmi+IwskkO3pNXM+vCfrMvxRqU4YskiiWqPrDUCYkOk9YevmBazJ66pC7APZ5rzq6h747/9ZlX
UPwtq0+A7Io4WGCd57/f7oJ9ylliiV5iU+wJm4FM8SOh1JrEIgNaroSwILQhHKLNh1vt3Ks+13Cc
1cu+a/iPeRw0vqbOfbXkYaR5gpHHiGDDuLg+n0Y//r1pq3+v9gqaIw5McI4fYWe4gO8nCbCS2tAO
CQJEWJlWxlirI94FeSYNPo5ZCxCSJDoxy2huboofJa+qF5jn9R8fnHpdiRWvWkePGgXS1OPa0KZt
8krVFsUhxj8oyTtyd6Zbtrn4+azA6978spLKGeqKZt/tioP8slAa7HTToZ4IepJE6ZJYAJGVRm/W
XtvRhAWLW3TaKFVhPiHP4wluR2yE8qLanNHSv+fD5ZAUyYvgN3w4srbmQDM6L3dy5I/hgcd1Lsze
8ZWF6CD9Ypep7xLSZTOvokt17Kg3BewSuuBl8scH8ssqHsB5CcbuJam2pXh0NbSRK+9w6YTRDqT6
K9w/sbqeQpI+Vk/CYGucw6xV5dsdsK6Qbcs0Dn2weDGfdcwLQrgk4Q7n1z4JcEA0GIbAST6/RZ/i
OvMnycMtws8d1aMPC9ez0jJ68P3tTCdRnoo+c6wa0v68H+3/xKFVUAxmE7ND5aFkI0ZTv5mT8ivx
s3elgVL7nwnkUGnFnNYQ/gFZ2TzhqPdnjDytO2asqLuvno/qpZZokIrzi4MJDoGp6LAEX1z5gGUF
Y80hpCV+m1GTqAOcBhfhhJbHchyXZDvLCSeAq1ic33ggeaIPpS1aNbnmRPBNg5N9kYI1OTyaviqh
KDEvxlyyLsQo5xXpIE98sQTt6RfUzO4ixlxhhAikJ4oLicGgFhC0T882rI+6nkdmZuipOkY0yTan
qcqbLqNCrbjb+Srlsz3FxAw2M+9FctQb+IEXavJyhy6hFQqi+KE4Bz23fhUKv06USF4v8HuGfO2Q
AiDTKB1tIGmvCOwnzN8yU61+rgkjcORpYDop05Eb/gtSYIZMb4JeKU4lxq5toElhkcBDOF4abqXL
BBdKAG7leGzTR/aBXkXaVEyD8AAQHmU4Wn6oH8s6p6BAYWfGl6thxD5fN0DdQHufPPAE5JSO04Y0
vw6goXrr0s+8e+3SsnjJHf6otTgD9vAVlLAdfvX79Ief+tv89+9Cv+CQu1XUh9U6skgK63s7ODvv
qYJYWahdBUva0I/H5AF5V8rRAVxgC8h9AATsJNWabfOaFLTTp9rv9oSJ/QYVmjwKxpXQQ6I1yzgu
sTnWT9Zuo/ozimdvZyClHa8oXsncY6C8lsz7b63Tf4RSCiviDfIwDd3RXNPdU2K3G/r4tDtDFv2G
Ku2Xbgcr8RAT06RZoMRxAiluWYbb7IHhuf6JYCZkYcvy5x8kKtqXgV5NGgr0HiVdVkBfXe56lEcM
CS9ZVgUctxoLbcUuvS086ZlfVw/9QLKPmKHCz6kYWwhRzXF/xWiFuaXjQ/hDnA7JwUgOxHrr9F+4
x/BpRXqEZB/wU4Ve9HIHtNbhtRVdUlkNwXpA7KP9/xCtujBvHbjvpISroL0THdmRf+aUaNR8F36v
VfX1KS56hmZCzw2BIBdhtvS+32AFfQGpM8XWpfXc/7FeLbCCkBdXVzLp7eWcPfhS118xqEpchhuW
ib7mFZFJCe9h0tZDtpXC0ppFv+8UItztQ+v0tj4wyP2Zipu2dv291oL9aEYLcKBFUK1ZHW8w5Rn3
r3bZZAk8GYsZgCrvf5KUZn+9vtnd2dhj+I/yRBB6H0g3NDUArw0pYUJYHfgaKOY=
`pragma protect end_protected
