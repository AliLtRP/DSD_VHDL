// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IAFLseb+mNs0ZB5zUNnM3xQpqpu2Mjd9aIsADPR0YdNGIXUQ7l1X4BYCn6unZr7Z
NVXJItMv13w7/4Me/QGGezlO1igEGi/CUHl41YWaP7KE8yVkTk52BBMnCGjzHhIP
Q3F1QhC7t7UP+qz4z8b4afd232hFjdeJDQRIOS9L52s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27792)
fs3M6taFh7cgh3IbrtzRPVbpJ6s3NLlZ5n/8S4ncBrqOjzsrXtkBU62TOKE5grWX
R8eAGMfNVUThTNcLWC/D50sMMfv+4xgwruwN/+MLB4sZFEesnZHRrw4WJja1rMh1
N6U/JR86vPCOJrQB8JpFuqFTQ9ffKZTnhiTGDiT02kJJq96SwKQ6SBxPxT6JG+9u
7Es7RJiK82u2qBxWY/zaP2KOrYEbkbe72xA2re2eMl4TQ35W1oFBxDqrXTqnPZH4
tZO+p+3/so+SoDVprn0N/1NBYzTw+c7bfbuq4CNR+rqvcM0PjQY76IW9n2/j4KmZ
n7AHtgkgaGDqs9ZIHQvowIooYyej6KinZ/1V5Uw33PToL6Ny1lNUJ3f7ZnuU1gZI
LDe3tprGbdBtPTItB2+xNkzPgmSrM3KbS4rTp3rDsaH73izOGCfgb6qszufass9C
P1FLvH2gAo30GYgGxMZQXUvWdHgZfyMQ3hVmJLlZw8zEYGLYyWfA4Yu6Be8iEmxs
jcKKhJYxj05ddCrmTcQ8bHOlfRdlWEspKYzUVSjmT94ZiT4cIDOvIRpQimxqFfaC
e86h3AZYvh3ffXpNoQdjLfGvmUaV0r2X64kqg3Xlxi5XQW282qX7OH7Yr3xC62lA
6hs7KieyHELa9CMnj9WFle2dq+sJuEiV5QOCGOgk+ovUpyJ3JuZHgF3Xyg8qdoKN
eDK3xWdkJ9dNAdcgwEORHyTgi7QsirXKfjdgw9i4xETDEv+3f05zBCUbElZKhjZz
po8uR2BbOJAqrgDitTsTJL8do2vITe2A72db4e4VqDtwNHEg9I/dxOA7usR3Azhx
pLtcciIJ8I2YTtErRp6uvv6zI9fTG8ri99EX6LxdU2tmW3Ub39VZYceHVfx1aQCb
mEDSrwkSa5caWGQNjYQS7xFZMdlvVFu+VDI7d5NNw57EM5XWH9awwO78uDpaGUbe
HMkfPK2vx6Izvs3cwt4LDGgIYkoozqBbL5FBTk9fDfze5lQ2ukj6cJA9tMP+nNkq
G/ny6u57peRdeUBYwUSx2M/JphCT+4wIb4AVXpeJ9AkGZf2Gsm2uo2QLDCW5QfXJ
pyXTWdPALAPCukvgGZBy4LJrant7Evi+Pd4Uol+iAqorhg0San0/nhUqC5SlOxQw
jqMahCuLBYR3Xm2ggCy15R7lgwoAMNxs7RVFq1+tBkovc+Wgpb4yrPk3Xrb5qhkv
KhBsFNCbaXvWi/FvZ/iXyjzHiLW2nA1ZZ/PdnSDlK7WY/lUeucsrt/abMBOvNxXU
IHUmu5CCe4JIdU3pqc5/NXHG5UjhMMAC0f0oVz6Phk1OBkeqnODa2EPdk/1FEbbT
NI0wP1flzAbVMa/77QrISzeYD/MYW5udcL8QRiojIlogPWLKMpLtVAwIC4G47tGl
k98rjM6OhCZ2+U4ZJQXC9nQvHnLqBfx3DtbBAviGFfhj86NRcHQl3OChc9yIyR0C
VH0HKxynqYbxX7heuZ8iMF1YAUBTxlfjnisWW7V20fu1TSA4m0GazefDYvaK13zf
Qe5in7TK/SqE0sUsxiH7Ss7cF91J6SpsIZ6RM3xNNhTqV58SFiTttyWIvmRIyjz6
y6TznHYHIpLIin/erp3232INVBFIrWXcJ2M/qo+ATc6JufNkMk369pEBM3tiiiZC
G9sYzzdwiLxei32BixwzV+hm6m6HC/rp8l6MhgWp0bKBIAZaSzGpldR+4NY4Ir+0
3oKv9Vq7yJYSJI9sTgAVmVO9nf8+fQP59cbAZCsk6F0hCDj7bvaGOjArzyDY8w3Y
59E0tYAvMcQMEzb1smKg1KJXBJ8qQCouapFdNXBV75hp4+O7twIITbxfEJHXpjIH
A6Mwg5zox3OcjFIF+8RkHNb4b5fMUhWeFmjnApMaM0CqDolQ95VOBmVr/rN/3gXM
AFIcnWoOa4mZ8vPB9EJqlzKflsUfTnHLC29bYGJDLfvFOp4bu1j3Bz0SJTuZ3BU4
qBtsAAOiIiotRtu39sJTGRGFsQO/z9N2Iit1SxcEoFs7oCq02dEEhvhMhRiLy1Ej
R86YxgsBNejZVI+8yabi6PwMVha7ckWLe25wc749Cx3fvM42Wv2rzb3sgcGzzwTe
HLhGZ5/15OYm3s65Fa6QqDs/LkvC8M1WZUQ3MbjVRkHiWV2qVJq2pcK4OPA0VS+J
GKpsNZhaVYDz3WTTqan40U6xvesUGFJnP9JBvf3pd+yTtRks1mRDt8ilAD6HtINq
FAMUNOu4KuYX+lFE0sfn3sU+yZsh1ajj1EDuDMWnwT9cv9/TYuouzS1kFZ0clTtn
JI1Vo/4Zr5kWaAzBuRM5WNXrSHH+4cWUW3jkpzwkpeM+dYm+kR/iC2y2CfTHtT/X
2O6tShnsbhfa7JNqwXXd8TjxTAAmH+HOU8JZFOSYNzVcRtfTYgE6h+ruU8mmx0F6
HeNP7hRDX0zFXB4W2gLCnQEoj5XT8KOLJHrKafwTAiRseK7sv6JQdrIE4NeIuj7a
UHVaNF+Dik2qnKNCCaPoEDSnoLo6Ot/WMFuKJiko+L1shofnuEykgm3Qv7rLcaA/
n6aYw4ssgzwrRZir2vGhunmoOrSSVmYz/NePLVgQImgvnZIFAmjS7Vbd6ZCxAM3C
XgdrTBFZo4NBglvNA94g9GKgIDi4oIDtsZzrhhVk9Js5NnlkgEGL1z1TekHvSkGj
CZiSAxyX3UBTnFU33KdI2KNQGkymrtZqvFfSPZcKiCyK6aKAi8gVgC/Wt1qzzLdH
Kd3GbGBBBWgdtgq3O3vo2uyRJHger1aA/6VLuwbUYuU/kPXrbeq152vFMvsanh0s
6cGMXVM+HEG9jEA5IE3wNpGoXKpyvyyd7IK4tuATVU7sqrG8DbJOFVY3JGiN+GhU
6nGhXuqo7lo5Tvp1EJcEpb2IuHS5ykO9xMJy8guv0FIZhKw2J2yj2QMoXJPV0c5n
/tqEZ1QeGhZTBRHJqQP1ci1/Nvnsr8T0qA5DKGhNMP7FwHFI6uWCiCIh0ofOy+vs
KsEc8bRWfx9cqNrCbb+JCHHd/7hHK/RcJNfPPeQU7NkPCCt8TWX3lHnYyLRdfna3
IO6FFGH+yg5n6GnkbNCyVn8Mo0z2HFqn9O883hYveYVymeRAxAbJ8P7+nslYCLaa
X0WD5lJB6zNlU5V5iNP7n1Wv2RDjYOaaorzP0isI7nb6rt+mvlW0V57Q1FCkKNae
uyHL+8wIgjXk6e8ww5xGhP0MCBGmsjNV5DTHfkVig2FPzJg8vr3QhoOEkiBuyclf
iB6yAVAvWnIx6S8X2cOQOshzfq27c+SVMZcgiBF/JO0n3K6ujxCVDvfJoECq/QdO
nfWLycI0SPRXh9fKCWMft/YB0Ax4ON3XEB4Zp/enpjvC+e5ZyRFDkEBPiP9O8GAX
tSAEsZeMOZke0Z+4/fbUAH94P+gf5bKNQZyzZUGHT31RQm16acwBTitFCbuMq+t8
aaWttnq17hGgu3zVQCyNi6ExHOy2g9MvsnD5rzslMLqEUDx6lkX6X2ejM7+P2ZCg
Y23n3F2ldP7+xrgcy+S4DNmEhs0eSboYL5ZIWpno90YwLLdPRVDBAt1/lu1ydAUs
9O4wxijs3G25RERG83Yv6RulUaaDU8UQ9wXgXxai91vhdMr+5M70+WKT3xd9w8a1
l3w6uw7fQ6vDTuGvUQbfrqs0WbrPqlza7Q9eSs1Ka0oYHk2P59NZI9ZUwnlIwLRn
Zbwphvvir4h5PavII8xmzA0Cdea/nmLv1w3UwG6WKWWQ9LHHqrl7AcZnBWkGMDmE
O/8o20CWT5eO4C/nutwXO/QVL5P7aFIWGMiAicgOrN13gcbqzo/fuC2gOYRvc122
hmvoiRGwN422lLeeFSU2+0HRxX0NHNck/WCE22rlMxrFFNnqSNLVb7TIBCXFWO7b
3Hx2yQDKDhofTpDCDKXtiL/YEKgFyEUTQDDZ53hkaaN27OIcoN8CtAc6IiJd3szu
rfmS3p51/jLJxWbJvy00LfwkWB62yW/AKDT+lsSLoxtUbyMVO6IoC0r7DfF1IGPC
ccSavBoTDSEwxnKzj4cyma64a2pDdwBWmflcdePbLgjWP30venA6K2+8rzfu0aSs
FQ5yKA0cjzvM0apxT+/OACC221CVDAMBZfKWrgOsdQ8V0EXf1Ep5D5x0JIGdtvXO
8bJJIXYzOgGLJZf8MxsM2msf8L0ayqGLf5dDhoOoQTlRBNgQ2Y4t//qraZ9q6yWD
bN7iFOdBeyYKkfwjffgIzSgH6TXOXngPOIRXy+CHljli+KYltmklZcFq9xwF5VWC
kTeo3NzKvmrst/Ky4ZcKgdjlxZJQxI0lD9yyaeeOo2oBWNEp7Xac3vkfP7hf3QNM
GqUJPkV5lHezU+fziDoKMtdqJvQU/eEt02Rev11V5gc9vWUtfINE5CZQwt0DmFTR
4P+LM13Uc2ViqsF7wZVDF8HZdm8kL26mczclfHgQmZtwOMpuyfhFeOrzZRg1EItk
mwkb7cBGb2/vrAfAFtu+pfKckYtqfIFdICZ1N1HpYidq4stigKSbL9T2LFoKHK2+
t5NxDvT3pcCGPgI5Rl0szvXQMEAwJfy0uiot4PlRxm5TDRSeMHdV5MX1S4vs/00W
REqzTDpqRvy1DGMzJDDoTu/aI7Ej9+2Ppyht5NCkOr3SofnAWcIazjRqIN1PQfHl
wqwQ0D81FqMsQxW1+z9monXS6FjOzvZegCCXWFgFSg+V9lAK0tIzqP5rDdxOaUru
mzaIqZHMf2rv0GubQbbTmX3Pdv+sAAuWxMF790cE2tMzQxEpT3dLpXvulLnD/ucb
8hIw+p/1+QNEeAX/f599jqtdk02YHjCt+6bIoTfyCz1Yem4gAmXPNpBU4wY1enr6
OSGIOwryo+k5tmQYKObEIFWQGNSwz4EKmm+r1BZQcEskmDsaf0cJz9cm5WwfIjbe
EAbo/A7zwEAxJQoz4CAoToEbTS42y2Im1WUVibJNCEc7teBJfqQw4B+UUvwHUoY0
jF5vlKUwed4ecgfnfcuFMMUF6yUni4PFWfNlzZYt77zvNyOELUIa/twlijqRtk1u
7EHC/bn9Eb4B3lm35JLNL9zQ60+vJuJ+9FSF1mX/ChMFozjuh9Q5IfnjpkuYUTFg
+xfzk5vytxCUcF2nkJr8P+LbHowyEJ0XHK4om0gNQk3cP5wQUpzmfJ8i7SilWN+q
nGNajV8FMf4FH24eKZIDhRB8iSVuPiUBwa/KIp5ahHILuNnxCsNe0l2m9It1LFY1
UbsqtPNZ7PpqcrqvaSobZk/Xgr47/3nj+NALFDvivYk+yu1k87+f/ZKbt+qQHtdW
HiwSUPGi8XsywD4Gf5i3RDpsb+QXQbX1LVe/NuWfAfnWhZ4TyBTtCiVQoQDf6sRY
0sVn09ATuOg6ooAsA0T/s6y7pNtr9W3ooJSQr1wHthxvp/po5jA/kGGG38Ermrk7
6nIvcBwtssXB0hD19+oGHrWlqTMIHk8pWh4CgCvgZmqtl93TR1z21QwGV0U7/u4X
wQXXtMa/QyIwSOBhMaZ+uwFFdUlSAnYYHDc94antrVdiMxGbl5AJ5PKlC50OGWrh
/F5IcABIP+AFqLLisUVW36HINEMyXVR9sFcAyESuGIaR6WCsi8eVYnt+3qqs9+ua
mgTWS+D0CNEjF8GDwdV05uCXrAqHhUtA07DTGYOJLdrE/ziu85aaEvyzcvqBhIaT
zU/jb858oaLfjCZvTJqGT0Lu3P6tIxBv3iaBkHcvwRoumNb1AysmepUIwTFbYwFE
VTC+jH+NnRcAhXRliwYca0sqJ5F3TfLL4bfy+3R4OEoqYYEbtxMGbndc1GmVlxai
emwK+knQPl3ukhbEDj8i9fFjQhiJTz4E0gGrYA6/C9yiA7fx+RO/hHrfePaogUsi
dukdPrEj70aPHnDo4cMI21k5jSznU2a2pOL3j93MXz7Ko+Umpvbxn4npj5wDVjIJ
9B9k6wy6u17snE0MjVCVUQ8gMiPc5bH7j89yZp9B0OnoFHmOkC/di77FoMMximb6
lhqaLVkNmPi9uEqU1fjYLZxR94PcWv/U4QfTZpFODsN/6s+kXCCOfwpsQ8cGcgH6
n0Vb5nuATxMJFFclegu5TZISnOp06dJKtOvXq0bv47wHrDymqXsKDJ75Cjm2JU0x
oKiZokwG4FiTMu/in3ojz78udvJsIzxgXLVIoDlvM5YTfEVyIE+JptZn1hJfqgAx
8GWd2qswaxD7lvbym9mZ+z1KdH4sOF/RbbpCJ6vU85ccO/slH5nHOFYS0btl26KE
B7VH2qm9BNI5owRAuXHqr4+TIAW8lBS/Lm3n1qjltnTAnHb1L1ec/AyJkmP4Z5YA
V6TbCpT56g851TqxE03FqU81gul8q848xbDu1YrPuLciXlF/sUhIcvN/RxMeZxYP
IW1JnYynTcWM0nS/ZZ22dVfzBdnrOd1ZUMK40hPKwtuRYqvQ+qvFlyYLAJuACjWP
TIO0w8uhVNnDpsEDVk9P3AJFrOOCqkp0QNAFgjMwMmjq0pA9nsI856PUyq5mwtE4
35GAukHTXHlQO/6GQdqbRYIGTecbzWmOWTLzf0ZN2isxjYxo9Z+N+JvI9kny47wG
5ujoMnnourcQEhOkFqK7pdBnCtpNNJZBJxCunr7fFwnrvVgzWpPXVSkpFge2Bh3W
RNDrWMAPLIbyQVqDOwGFriPEPQAMRSrc5ZFShgCRWYC2o2xktCVW8L26fg25Ro9+
KkiNM/1peeivm5c+Mn8BJS9Kvyo2/HyhGX+BzOzui3i0uFx3xCNwKT7Siy3w4LTZ
/69/mcOBT9GGJMKCqxPiB+4evSaZsZ3pTtg+EJskr1YjpTqWtbJ7g1ewMYdJKuNA
AIt2vWqcr1Q/luVYBQ9RqJhQuVvfx0FI5nTaEOPrfZzmzNFOzhBKNWATejokc7Mi
JwUp+0Nq0SmLg3yzcaLiJkK1WgbKy5LMSU1oYx039qrN/aHnU2L3HY3Sj8SfIbSP
XyamxUPQw0/jO/y9QkM9imLTU5bwAvgqR8u9o0WSKmon573lQbZ/wJ579ha4WGSV
GUgEVN985aMBKB96+IIOK98Bm5GaLBIxB4+xobkvreBsptt44zKLhGdmDsbk2cDc
0fZGY0ci6925VLhnx+kedsZbwwi+2n0XO1UpSl8XT/isbvRtZNVasn6Meq8UEVJ6
u5LsMJL+W6KLmi4aQdz5R9tTgG8Jgrx+M+y3H6ecNacfXJyQdyzoO6iJ41amgYbm
6rK+9cV3yshO06iy5sfUU4s4XSRxlw56xVYZQTdlJKMiTklqHh0vKHoUBFNMZE8v
feBKXQwhzAFFD0QaHIuJjkyRFCKch2P9fUgdmSHD9ZQT1OA65Kne3mWcNTVw99gd
x5LAXF1yzDqBmmNdccRiy/ze/5JwOPxNZuh59QWVBTlh5Cc86OkSWgp2Q0dtvP1C
F236TEZbk3f4hO+x8UWjAIZ4W/iBYiUdALMmgJgnSyf4bKqmULHjdS8MSKTdx6SZ
Kt55yB8tepGgS3U0Cmy1U28JdF8FRfY7FqTCA0433CxsPi3QDEz4uEW6fSeQ0sfA
1u3dbiy5E46ZOJdzh+SpdjnaqkXsKwkRFXfb9b2oN/aRIjWjUDNv+XAgaq7MR25f
F0tmPN4DfWM2SSVlIWXe9LudU5nXvgpUx4Cc454ztZfngiDN334l20UzmlJnoJfi
mopLwnVEYqyfdD/AuVnZtnNsGlD8z4/grFVqiazG45BUiqrbMhQzVr67OJfhBZyN
O0ZbbWMqt+jns36cdcM/OG6LAGMXz82cntkZwKS9YcsD45wTclLgAP1jZGe79LLC
L9iZSgSAWkTywIM+MhWM4Svwz4bFN/k+WQpBOdkl2UEDvb8gTujmDvCEH7xkaOhL
IckURoQsDb8ruxMb1av1QEfrQ7pH2997FPNpDnIkNzBeQvMJ9oAbNz4aRRl/HR3s
/Zj4TC5NxkVq5FXS8t+L3ON6AYYt6RnlVRaqn/0TvLmc0E+eV0Jf7DGXHrmzadP6
DBevcpt1MAbK6w2loBVBn0E02sdmebZLAQnOdxpw1O8cJnz4qjFqDflY9Zv7Lgzj
nAN5NhfHc2Wrp1G4FLur3XCbgcTcRSNvf/mV7FODhtg0zXROOIXaBLBY5ULk0vlQ
7TOIefQjR5ujOIuEKiyfyJqm1hgKsEpq8gf9l8sjWCs9wzgi+nA0eCFuUhQ1bTEx
fG04gDEIX+mJejaRU1IoT0sdQUsEkFHapYMz004HPWsB1GnLQ01QeWBwSqZv7tDp
rV8+nQQDbnK3BamAVDrmRCJ4J7YzwVHoAGI7HTCQtPHRpX872dCT4kdSw66HKYuX
+ZONv0J0FvLv0x42+J7Y1HDZTeEhbzmQ5AlXfXzuOOgHXzrbFejEBevVUyd6ZTpF
7B6iG+GKccwuKNQgdbUZJU2aTc90t5KCmnviM1MR8wwGZdtwKX/7wMhysEpZvxiP
vwW1B6WQhSLiTlesnWQJ/oKaP0mtS+k6sISo5UIZrhua93OQeDPG+Nibj2A/863k
pv2FKOo2AuL8LnwTcK31EAdHrGlaZZSdzkGfTRfzi4hc65bSypsb9QZPDXwQG6Ie
HQLlf5qYZxmVgYVo1fJfymjBD5fBnSVvYFxT7HnaSIfkHoLhEqcMtnxdBGMNZgd9
U/8Snm4eDd2yirqRpxL/Oynb9Yyac6whPdOn+ROPFZX7b0GQaWN6fH+runSK8fPH
loHLyASymRgey0cEtH0ck7HCvlTZ4r5IlJ8N7OaGswPlbGmVZJbli7dybwkSKVj9
L+7UM5Ca8nkyO+Fsfi4n/0TiIovzue8bzj7t/3M/qZcuiwvvpsznm4Nb/XGhBRwX
ZeyG3HZ10igAMrLj0Q9t/JqIJI74qBY97xZjTS9naOELjG1H8deVlbpomn3ohJ6s
SFtwaFI1/a2mhekOuISrauxKZoZylMiTSDoByXnLmclgFvVnXKMS5SPRBg/CWaOl
UrizTC8WpOW0frDI+fozhb4IXDm2pOMQl8zNfiPoYcytGGBjL9vuZAJaQgl68T4k
W3CUB2ppSrsZprRWRnrmARNfosyazsZM7D+9eVTCWLMOpRApvSziyFwksFExk9jd
1ORfnKUlPotIZhLmYeRXBgVU6SuSSzuEmI1dtFGP27ZJxOeJ4Jb1/p+75LUsnyCa
wOk4RAkBZ5LFp2esd+0qsajgjQ9AO38qRtKosMLqiFDcnPQQ8O4QHBfh3OhV0U5o
fGl/1keDqcS61qjMpRnudIe8Unfcs7OoqNNhXn1IXyxk3NIqms+GGtcAQlkW/w+/
v3225Lau+wfeAHH1LXgKvK6pxUMbSeeMEC1cWz0q0UTaMmmHNM41783cdetuYF0t
WWOrBAioyDFmkCM6mQJrLrck85DHoXp04NppiDE4YbsYEJIW1SULrbkWySFlRrJg
Kun3zMvlNA7p2+Udr/QTzp4S2sXWu2jq9OvcR5IekGjzYTTzmBnOATFII5gcSrSH
+Tp8VglBUL4xr4riDgm+H908i96AizB/iwbaObKHmYtDAVJUyaAp/rb9HE60vVSm
JGoNYpjhzutmsw4E/N4x1kYttez9NvPn8WFDJGVGZ2LMIpGpFULpIpKFD785xG73
dP4kFUsOkvsZ93RLABO8IEkdFQA/pUNch4qcM0xtcEkSv6LAWrw2KQAa9QJfqfIP
dxIccU4AlCs42fwOlj64aebd1fthBh9gAxF6w+jioBSl4e5r8iswFt8xaRIRvgo0
1bpCawtd2HAq7l1alhnOQpezd3G3kbXWwMdISP0dZAgTrQseMCq9JL1TGOIyf56b
vSK/WsBU8OMPSopnBBg8NXZg5o4XBaM1K1/YYmaR2d+zPUM+lYm92iyV0eleZaQ8
+g/lt9+Nb5xDK6AJsb/LQrqImzzyQUu1+umtWYh7+cdAtFZ3VNByWa3wFAExI9ny
f+T6SFevIppwWEauMduDiGMiv0VXQqIzgMZ7J3IifOVA61xN4jISgqJSacxyVh6j
u9PSz98rjnl7IXDT2kwDMfLx152foSFYYsmZx0Zvf6SKhOZuEw1lasyG9FuA5HAE
rUMxZfg/M/++SRvLM2NVAF97m0K2KI7vy4P0+PoE1YXT4pagEgZafNiuiGiNu+Dd
46+JA/wuyCbU7q0jDTGCYuT/7EbOTWXoe2qI70CcXuP/uJA/VA0uCcmB5AAA1yrd
VspqzI8tPEbmqVBhHI20RSAS/kyo46PXy7ye1PxjY3+VZJkRe3jHILYJUev6htoH
y8j9+qBmLzBKJ4ZoUh7+6dScZhKQbyBsfVn6eWECcOKrhyT3NoTj6gN3Ybsd9/Mu
9/zBwErUom3zGVVbF8qQ0FJdfZ6M/I4PFBBnogB3V/Nhr1SIijjzXjYPYSxkvOMB
9Mwp5719zvyrdGDo2WUrm8OYOpr/x7InN7WRmMntAv3SOqRjoASgqSLpYyOyx3ZZ
xlWCLfMY7KS8/12uHVa3e6TDbJHEQab8fIVsGTxXuiizquBt52rYNgRBZMZuLpZD
TTqyxmMgDgQIkfxRo4XJT/Ay3TI7G/KviQwqj11L2/P8+0ZFPQlxef+oATs3XfWf
Y0gkEnQRqAGIRlw+i6GAwhPtgscVZphCoiR6vnUEw4DbkaFcYIzEpzpGNzUdTXuS
8gAn9t8yCxHwgPIQc2oboJF3DhBd+Nr/KsFlop5IFz2gwXW03g5ld4ZP1YFr5YRU
4C/MIVGd3269zpgHyo1obhpg7YPeVDgFX80YOz2K/SjH2P3y/DC8YXpOivI8shRA
FJyd7j8Um8Ha1U0FTQiAO/k5REfAkXKNnI4L5KeDohJjddBjTfpoMsqtWakxP1QG
wSOv6JWIDLYhr+7E8J+16N4MfkdKD0OAiWwyDcYmnqQczDgRwwX1vZHzL+EqstlY
6Pa3N7qertKOmRpFitez+mTfbukcXVe5xjvCK0cb6DiBRN3ePrA8UEkqKqpaPWG9
oNSJF9Sz+TASUuIlgwbEG7wTUW1OuDMjwgOOFF5nlQw5Kj6plrvv6xju4Kur5s3h
E6AzJ+4QeCEniR++NLsnJjn6yYFxdjtxoUwar9Clail/kXb0N5+/NeKe/AgL7kde
b5IV5ndahCumP89C374boaRw6yKGD09nwtjs2Jfte0DnXTW0fyM4Q7E/qVmEO39U
kqacMukZ8sFdbVLJTVL6k4EJDaChYQXR/TF8Rgj2+W82FJd/nVLX9dFy9WcAg7oh
7Q9feOz9kfsf6dFfW8LgfZ188MNCcHY93aLYKfjbzYqvbCmdJf48xnGSF3czd8mR
C8HMDRoCsR4xWMcN6Gg/MwxTdkUBRqPnFdShLEzVzI68Yrsr/aOXSHM+7Rd87sgu
NLxQqpnR6aM2mi5N7k/sAs1cxOxO0Dy5aFopueCQIfpjo+lmqhTFdZZ4EGktufwG
dIsUx7aZD4KRsoNjCDiXdLfNGKH11NqYgFjaTUzdj88gnjpte/fsLJApwEzFgiSE
SYvVXI+/AGGQrODoFpHkULbojd4n5IxwoTNoT1nID4pbxZ+iBtRTdktlt3O1fqX/
UsoLzaLG1IjhUCmF0kaK5ijsYdivwErmoettpRb/Vp150AxekkS1mSo2oNyyZsLw
OXNAtYxaXis8qGpbzAgKrBRqUDU5Uhx7/x1RFEe1KZJeeOG9jZc/UAIbJhDH2cn1
lmQi9dQxFBGVorDkRK+HTi+F6Tli/iU1MNpx1b0/G9Z6MqUNRe5S2TNUfOYlDJ7K
AZ9ft4kDLK83VZ9hbeeY7gaovGwjvK6VqIbFgakdZHbdKbXHjkDWBI3pIZkm2Het
/1g50VHNe22xtNBd7Gr5D4DzMGdsCYNNVLQFSsozC0B3VfkQWViisR7f7e4FUxvM
Kt0g0amTq6Nbvm5FUARWsops0chjKaIr0a4kt4s8w/WYmqip4zyCzqQKaqXPSnoA
mJQG6j/ArNx7AK3Ow3j41E5tTavLATQx8DLnDnbQ7ZC0sh433jGAMJ9qlOJcXCl/
cU1VjFkSNidKshHML5pAKjQ/HOiaSTdSCWtnqpzkOJIUJy3qTfo8u+20d52L6479
y1M+2bc71qbECha3n03EP0So4mvsj/OlYNvkxCzTK+NZB1jImxCySkFFmpikmLMO
o8Kaa457r54bwwtOmYixC50wwqZXzl2uB/i7HsVDHtlcxPHCiTcTP5uUsEMv6rb4
XfQ4vpKXlAxoAnFyyTE5Bgu1M2Fj7B78KpBXX8CoUI1wPowaDmQqt84fd+kklrk5
gF5vJPXwG8iU1rSusuJLbPSjARwPDoAePcgUSHrekaGn6CKZI1tSA2jI1A8hxe2D
LJrMsEJbAaCMy7gUvbcevLhMo9W1aoO7G7PGAfMiGEh2M0uEXb58+cctPgOoB5g/
WEUkvmO9gbz21CjSG5WRODXAHqE4nFLBIOL3NhF01y2ppw26dsput3wWt5Vhks4p
k7FeqiXXvRDFR6IJYZpJMg0/lSXu+/OEpjJZ/36sxTRVatYzireQriVGqZLES1tE
8Ssf48mcwrvJHP/oQdrrMwrguAF+e0ALilF4HOF2uxulO1lWNEIi9V84eqhWnh47
YH3LJh1BNbOlnf5P8VH3ugidqEXXuvFSV1EcUBfAGVm0bDe1lkW3w+pDx20drlmD
6RAEYmwdXww8xAD5GE6Qv2QA/u3Kfqtt1MF2sYqxexRoaDZN5H2yECOw/+yJhnWr
Al4SHg9hYaBNTLH6Bhrfp7qpiISez+1LRDKjLE5uXLZhRwfY6tZeGSR2We9nRyKT
twf2wg+E+PxIrIWS1sunV7KwrXvAnBpzmS+R5t78sY72b1Y27nwGnEiMCcdem5di
cX+mwUlV426tdBAeMziDxkmRdCv49aoX2riGBG950Kb4TVHUKZgIWnOGqYXOZ6sq
RVZ6zy9eewyjb9VP2zOAsqBm/7Z+iRpABy1Sef+B/SQ/odYSKO539rA4FVv8HuxZ
Osz9Z+8i+o1o7eja2gKvYZuViNbvaDef8bH2esYFhOeLoM1dM1l9UGB8DyqqyUcZ
VHU9cCq5MvDJVKE7PNb5NO/VmHlT0YtbHvpvWWhY9gQitKq7TMqeZZiI5g1MAi3S
Z2JMNdg2FITT9w31OIzYXzlZut3dP1ETwzYEbY89Yp18OiTEHMZwXwlUqW6XG+ok
RkdUJ0b8483deXrBOe2cJX1b9sWnmg/eVKjhtpJwZJtVaHloQMTnwzsNxiQ89sus
KirqwXtUtCnwxn7KI28vexJQOjRUYm5E8xsOA43Fuy4jjdElTMehxRZknQDe9cQo
iM3EhtU6JFXkpczppWrHxzpxK0waJQ03neQf3czj/Hov2VC/KiWPebEHVO+AI57g
iHR+3SAw1q7Ng8wi1W6NENFNHhMWW6x9VVxdtPqkBUYrnwmdRAyJp3piIi/aLEiN
sdtC5Ej3INjHMbp+tpUY1wSXNf4D/mP9Q2Z+n6vTYcqVjW1nOGH63DvRV/OQoSnL
NWz0ruYtf99cQW+wlIc9FL5ndckBt2VCG1AU2KxwfS64fdgjPCdk4sOVvNn0g2PR
w6HE5L8BpOEZdbeEFiUbC98mZlaJLStH8w13v84xkiNO/WnvCTuO/6rzgqLYdRoR
ytQWkKOMy/bVFweYhnLNhdOh80do+nrKkZFGMYSRtPsm1ge/4GRc1oP4LDSUA1Ud
TsxeDL2LrDQM9WsDW29+Ip19uBMSRNnDKBnbRa8JNoxkjx4nBmy388SaBY/IySpQ
icmkX4beWfooNSqcgvG4oL++fxIPeww8Zb+NLDucSDA7efSqBW/Et5sEtt1PJBKv
/pLruQ1qkx3hYZgz6VsdCQHPHrBleEkjMKr/FhyEX7IMWc+pnDMXNNK/3tCBEoRA
2T0E1rPTM9PXOYLBXSnQGY+SSCOvimEEvAXPYSJBeKa1jhhMIzVZZMvDpkz/Tqut
BXDq7v2iAkk8JA2kAb3oif9rxxgVpcxJkv9sViW+3h/H7Wq+A2g/hb7iGtt5H4M/
Mvg48ZcJk37no85TT6fq+NcVyfzCtFpvmIdDM15NgduxXwD6XxwcCIf7qv9ecY7W
LmKCB5zSbHE4PsCJHiuILo4OPSuWf+J0gp5oIqubKZtXh6cRqa+eFvzQF4TXx6+3
z4JQCU6LvFx79vfXnwnS0E99msrriSBrUPDIHDLjU3juyBq50DkG1o+5LxfgA7ce
9zw+42GzW3D1RxAzyaxAyR9KzgsNiuu9oU3gYuGich0emn8YemHKuxWav7YbyRKV
mJlSsK+EwrRJbaveWTk7/9Ky1fkgBrhj2wTmg9Zeva92YXaN7YM6WK5TYCXJofzv
VzyFgAX1Mkr9+9kWgENLWSU4+4bUxVDsZhOQAumYrrTPiagEp7d1K8OJkQYOkNmm
BIumpvXpzZlFdzxrrtpAhXO/M2KGkzQfD0jR2TVLVQUx/fRlnXYask2hxoZ0nIgW
S8hbHIuAWBM5ncaJb1RprVzkF5yNpqTsBnPj8qPaLwKiqQ2BWmO81M/bt5dt+qKU
fUuep+rje3SO5kLtYpazFJnp7ihFnnGDI7nd6dpfv+lBpmEvsPofa7yosz+/+fxO
GR7m4v9dVa6nK8LI8QsltsDi5Vi0sI2dyZDUJjDOLEgpk02aQBXOjfD2oedNMSRE
G99A1PJrJvaRM7FAamYrGvvEigE+ROAy8K8CgkmcZgLYhScm7FvRZP46eDlQoqpP
3ZkLoINPY8gBdN6J2VmAGTtCB+HUde62cNW3XM2IyOF7thpm8a80rEhv5HBGU/OF
ArRsiDxF/CrZ5Ut2J5ToI3MO3H0sjn/jLPpXac+4BAmE+8NMJJtBC5RSFoey4gpO
3E2+1orBy0lUPmdYqjFDgCcjtaXJ2pn2NVpvuVkAfwYLjxNPlNOoFWmvnUFAgEYv
Gg15xP3LiS7ZXoN/NOcQTl3rj2dHwPrQ7VqyeLHtyMIcMpLYLe8uShHQI5UePnUK
GC0pm3bIaDIi8vrLnWySqA1WkCWs9jbuN7LK2HH7tJii+uCMgnNqZfUCz+UxV7of
t1c1HNcVLWB5wkQEmznjXNNFiM4ZMj3dYZteRqqjQykt0tcUwkyuGHy3RijFOOkw
1Kr5iLJ3c7NbsqhU6XuV3LsCqfzQhymO5a9tApMyZYG/aMj9lya+mx5cHjRM2MKn
JZzt9aVg1PHwtzc5N8LqRCmL7UnYtgzZQ3kJTmuaKXyDBWKSpPp1KnQ+/Ese1F9s
pJzPEbQu2OLpvcCN943pqr5c/leOoCfA+1S7JPrxA8S7CoiK2JOk+JcDI71j7kJ2
CbTsk0qmHNg7ZQQJGAYe2sY9Evvep2aEVSJoh6RyhlJUsZax+t9PpriJdGYIXTZS
1kfFpJHN0pW/iIRoMCePviMqU1dL6b4klzFZjhbqdNwebv/jsN3DRB8VXaw1d/Hx
5yvjWObDnGzzSDcuPd2r4LVS8lEZpauKdM2unq4eSLJu5ToaahadQEsY/w+8SRWe
k9fhnfRaRrpNwAzeW+iwswRBbtntGvCh0QWIIFOxSj669l+/09TW/+ipAi+Vq4MH
+Cna/mpKfeOHZKtREzLLYNLhocdDLW3e0K+gho0djBdQNyNin+MzybCyLkuqN7bY
KMCcLMGg5TMNB0e4TGpeomoagVRvPEPqHoaR+8FJ/gnaOxPGKHjwQwg/6wmmPetb
ldaYybnlKx8g718Rbx/Ke9hqDTqr2WbTxPU6UFb+Xi7Hi+CXAcLPMwZmrYlWdC0a
80Wd/+EJsMYoTH5eo5CBf+icx+sfAEcWq50tnQCY4vLJbhAlchtOFO/lsFgoYXlt
ayZQ3it4qehqoz6A5DZ0u74Jooe6yrxr6lxHyS367RUP6nPgLCeuExAS2VulmMKd
CkuRKT47Lb8l1Ajm3UaiVh5CS5vlysCp/qzVccXWu5uncwEugbivuZlAraZm+MGO
qP1rSRk835KxicLF+W75G35NvEQoSzLXkhc14D2lJrVUKgc/HavNCoihJ5gp0oNy
qFd25HxHH7ggH3enwcZKWZiLPo+200Na60rfd3TtHRbjP+LDg0+Olv8Pht9yRb63
I+XipUxW7kjR8ti8HrScO/70b+AOdI161YVxNYg0VU3DbwXc/oxhPT1SK+ceNF5h
2Tfxo6fYuLZaEWV5/nZ5IN/Hz4tnhJer8EV9OZi+dKOv/BCpAH479kfSUd922yxn
Zhr7MVxFJI9qwrL6IYKMqi4sXJcdQYCKTJPkHPe7obQPK3VQlk72F/YzMob+shj3
1bEzTKcL+ww3Oc4j9q6+MEMfLHjeLE9uRCRPIfQNocqaJ7TyzBPacp62gZz4aZLt
dDsbctedGDiEjwVx3KcBQgPhLwJmmYq1x5o4r8S77OgVcDnCj0TDIq7PzX9z6M+v
dCsEdfKc7l6jOhp9GdQnrvq9tUyHXmvE0oHpcu4CCoC7uqKk3Svvf304+oluJZVA
1MBn81CmfyqT2UrUOyGFcrTdhmJPjHHRT6whJTaSwi18ApjHJFnm3FflPRVS5gsr
DrA8tc7MkbFK762S+x8qnqDsDnAPxwcEIwkYAE25K9rj/gBX6j/8vS9cMp9Jx9+g
2C9fg8p2Ym7K4loYvGW3CbiojoJhIlQK9trDosbe3qkRuNoE6c230eBdIueV3D7e
6A/fzL+UH2fs4+9CPp+613jR3ZVywfuFO4Mkpx2pkjBNjtr3BfCmQfO3HY9pCKG8
Iwa44e0azGNZhO/CEhL3t95vkjuXs3odMpdY1hZkln8S/Bd223TSaYMsRVhVJpPI
xVCRqJ7Flen57qiDAdRwmDxbqnJVTaUDsB175W1bg9ObT1WybQ3Hg6j+1VXSUqIw
NnvOoR9KDEysR9FzFsBxCGhr1308K4WMxIDsipio75Y5eqM30djWFxLnYhk8OL4H
sLq50vW6WsFWGrBr9D2hSkJi/k4ZoA8aoJaGcoAD+0FHjZQqXZK/uGPYL1rSWJM4
2Tnwej1xptT74D/12WMEmxbTOEW59npFqvtR1GdPyffAgWFIGRW39IFfs7MYcyQO
JMFKS7lR0dieWbBXFoHzrMn5vZRpCi6kiihX6Cs0cxJPsmmaStT2kuAH6WfWakjl
fErzDjWlcMwMXGR7McPprzeEkwSIGsJnzbnTk1Lt4MOoi9qVaVLvaoBRCB3THHcn
5ohfmd3oH3ti35KQlj7Cdqr7aGrQ4PLN9XGZBl7/axapSbRDWKOB5I72QLcaMATs
1+3k88iAkD5AYpwJIw+LCMgDpPlQdXF/Bj3lUkKWU/I9384ul0X3TfgxkLrHnZRN
oN66YWjQMqWbAcZ8BHOjSuuO4c6uZlctKaycdQfwqSDAaHbi6SAoGXnL+FTiWEiz
P1HT8SoEFAvvuSNmuTO61QtAQ8cqMwvkPflVx3Ks7M5AIFBY3gRjWMVXlD/2nrFV
Wjxj98OodD+cbW1jekOhWzXyiuSNGCdTLWC9knOuyw1MjT4iAaA+oU95MrZb5r2F
aRUGhPKwmRkypOlyKLuRM7pWG2ZZGrF0vobFGjtWBNu/yN9IA1+3eL4ViOqCvg5l
b8RUYj7u6uJZfj1qIPpJ30a9U08MBnniN1kgCfktS8+2+JBbRhZydq0eI268AYxC
uA0yT5GQyxY2xNkKV/R1iI2F/A1ogG8oH/NZtgdp+hAOo+dqqoMNEKx6e+GgsvVx
4jn7tWV9qDINAQ3qBGiKzG7T9IUiAAWwBEgcACI0rZW6/fUjE+o8by/o/U594rLZ
RI/0n3qrIN1AkhwmkPwzSjzziPX83/e2IaB1hJ4qR+7qdQXp3YGOi92AUF17C8Yo
sv3SjTPqRmKzDFGPM0MQ/bdU16th7lacm+WvDkMoH2jXLAdMWifEhG7gNr1S6pG/
CXEOQvndjLkaWYNEDWjZIWwQnAgHtd9EwFyHhgauPM0ojq5VC8W9PQGJ6nUndGJ1
q5d3FAUtNPWZOPDxxPNrzeoUY5ECZc34FmsIM0l7ZFXWomjopODre/hG9kDsoFtL
3dpQxvire1KpblYsj1qXCsAx8RmqxfsUIV+zQZy5gMZHZ51nvQ3zETje40PCWPAk
sWQICACcju7dBv/uz21xn2+0ssUdyWBp3GLGwpvRTXZHHbn7AcIpI9TaMUEJenOk
d4CZs14hZyKq+67bwML72UfW51rmfN7d3lGbX+F2jWXP8GAUKqx5YnsSIwO4YGrE
cecZGYx9PNnIKEGOp4g6lPa/jg+eYNAZ9jJpLNVh7pgcIs5YBt1rl51F0/HFW3Ap
F1jPI++BXnemaFkbKZSnXQdiyHlryH3oEXptbwkbhKJfO10BEOrYVvWBS9oZ+7Yy
STjqWM5sMfAvA0XCGXWAx/q3bb2EhcRm39K/+DUCTLqMg41iY6090to+BNls7bDn
N6h/NOaMnBQPL///YeUt/J0lUQKPqcfA0NVwNahnHvDLLk+8xtsU6K7M6U0IxdOK
rd6VPecP+YOrYmdN/dtmChwISl8atiDyyeUCh2Yobm90xKArZfJGPSQbci+6GbGp
NVhuaxtkCRjKkQAwHWF2NYNi4CQBdFzIVqTfwKT2vNLjOoz8AHvIgQCkwLCr/X7E
Xe/0k6Iismgm3NnexyQFuq0U4LEmNCvHNzR0vuMBQFU9hZyrodfhj9B0fGfKYum9
Cg67z/GC2hJnNFL0ooY9zPXBIwYUKIDzNxpk0y/FfcRX52ouQ1AmSPlzVQ82bSU+
gTLI0NX6NOFnH1v7kxBJW43esH9mN6l+tPo/+5R0upaQ4lFR2Yh9EGFZHMReeHKi
ewVM7EbjCxLqaHa0SBVzg3IBRUCQkqoQNIVtD1tST+cvhJxMZ4empMQAbg+1J3Do
JZ2GFl4idn7W2waJNsnkiXcmWUccQmVln6iqKLAeLqfTrDaiH0Tw0NyKKtu63TuV
j/ISULl9iIpM3xk6FIYsb7GJD1websXPJwwFZxj14e4G7vfVCoRgt5ACwkLdDc+5
O6Hn8PP/ya/9r26Q8q1SYdR/2eOQpa0Qn/Gu1Rl7cbPkOvhXZQDhis5F0j2cpvix
tP93REGAesL6fP0Dk1uLY9rPA6HE7S4bLbuMPlgYPtzdq9V/oH6AfBE6yrWIjdSU
mEGlgPDf0vPtuzCRAxJx6sLL1xlsRlEQbzG4bS8xtA45nIuBR3c5vILN0UhLE6OD
MBxhIDxP3hwH1+wXcIFU4elgS2tVqgbOCfABLBP9ZDtR1YkkrNWV3M+vTzbiqxS2
kYNH3G2fwQ83nkJfQOC3xrwHynpsmE0EI3g1nHx+DR5lKllte1I0ZYQxzoiWZHvU
SzqLLqY3j8H0JKIo0o05Exmk0It8q9SAqR9ZknF4AEZA5xxNgGpQuPKE+iKk1taL
3tnYOm3XwBytEjjGtUhkFeGlY3l0AUzjxgSJaXeD2bulC1VHr00SGdqTl/Gf1Vug
/GDKU/TuTpiU52MX6x7zEbI3aa+0s+0+2Edu+1wJ1zQ3Qm8hPUdJjPjf3eAh1+ll
58X/CaCSKgZc4U5LEPU4s/IdRWlNCABOopHxZ8350sUEi3WNiWVWvQFXj+HrkueW
tYadEpheWkgrg3ERIkC04PAdQu/LzZzUl+Bi4LI+UNCzJXYp1bHx2DEjaHOEQYpb
oEkHov2/oM2eVFCAyeByEkZIOwquvmUlZH017aF4NtDHx8sz4rkXaNiQe4fmpOzV
Z4k5wi2LSbdKkm5CcJhI8HsPdoFrFNeTISCG5kC1f2BIGq9SByOraWWKZF6npovE
fxdQ4xc/lu7i/3ZlP28WS99ci1aN3qfGqG+TwLuGXsuDBwl0GBIaufJoqHUqRoZO
8cveUzPkz4wHk5CqXwGwky3J9dOZvGEFteoYV7/E2KharRPnzCmCEV6V+F8koM6I
ffxjvrUtQvwepRm12yAOXijS9chVGUXS+rR6xREpDFqjQEkNambrs/tLFf3Q2LEI
oNOcj2w1A1N4RGHPmJ4M3Jd3wmheF6vac2VBGZqEDoW1/bn3NfBRazIAtE28R0Z9
kgU3TRy2zo/PpCxtzOVUuTaJxmncq/y1TwQsjT0fGk/77WJLeXrstcDBakkYKZxJ
9WIcDag8xDmETxE7mrYK06EsLy7w4SsgOZ0Zn79umAekUU3LvqozBRJZHcI+ICzs
a7gEonSML0OYHsDGo8sVFtnr/UWi2pJwAFmZy6yD1hlZxKTNl/pURVuArLF5APX0
0XJVwkD4p+ViT/FLXD3Yah44IUrJtp9VrpL7JD054oLHXx9eHuX3FoqZi3O8NWV/
T+v2fQDkNFKwBH09KCl3GvFQ4PMnEaJIZeSkXN7WljF2luyfknnTxuk+adsTHEdX
aoiNAEaiyG/FWaSdIftbPR+YfnLyaTOjeXB/uZ+X1uCgu3Ttx8wr9rsIJL/lHnG4
S7K2/7Uj8p9BidhCs/56WCzl5G7UOyMO6Aotls78Yd2+/zMA/t3voxUF9l9JiNLu
+fugdV56irg2tZY7dxot3kHkEY4hIc16M2ry1m8EImgN9QOpJv7fhJIq9MD7ZmWc
UjKuod3ahq03dWFkoyNDrZjEc1Iaqh0T11I6oSOAIN/nA/0jiJZ78bCms7pTJtI2
cP4XK6rDJI0oHt0oSxdQA2hTr5T6T83ZL/pKGy5oYzFLPyO6NjYZk2EZ4fK3KM4w
mO4tcdSBOuSmDWC2LCDKmnQIyY+V2UCPiVN7q0tmWj8gHjyeCrD+mHnvOQvSdRKh
HHDTw5pjKNM1c6daIksYNAahQdv54hke/c0OotjnDlXPD7BfV6lS3Y5Bcf5h/kWM
ZuL5pixG/tMwhtL58cOEyX0lKoebCPyfzm9riZ4+ZyCLspaT8OyFAlWKjycFYATi
f0fXOWrU6EI9XhLCIhuOhYQfvsUkKscvnsQWHBzLUoN9UZlkTDvps35Za2Y88ACR
mowGukN6ZZMOYHYbcaMPV8PofVpUVnJ1PxH60y+89jm/m/eswizQSacu7iKBu363
IrF3I24RSHlWoMftiKY7m9lesiGejWAZgTGuBvdjSqXQ901RRmq0VQ/RRrCZM9Ny
F1e63F7yV5AnXQ8n4h4hdlg6LxCuGk+oZTLc6EsjjIx/3pPuUziIvuhbcIBn08lj
tBSyBysg9M1ls6vdTFu1BWgv9HtG/t3YXjGaVUyPe9hnRPJINjNpvm5lRC/6NgZc
JiXso6xYUEp9KBzhLQAud5ff6JlMJRrdCZ/BrzkNWF0bZoW2DX12D57vb/1Gw+aN
CFNy5LB73STWCtgc5HKcSGj3q5ms1gF4NPYlmr4HamjHEgayIAixOaJypfIpImYO
It+uSMb5AHnyeEFKzVsQQRgAumgX8XgwpDhyUn/XiJZE3twZx8rczfSaqfLaC561
SNfxJz+R36RMEvY+aiV4dKQ+wqRfdF++/un3JtlRLEWOtSEOMpMVUaswZGg2WQfm
wlKUbCDygVovcK9fKliQyfujEkEnTQBOb4dvr/lc5E6CoDXzfbGii2E32abm1whi
Ovx2mEV56RRgB9tEAJUvLvfxOywWJKJ4m2kCFrqp00sHXQvOUqmUzwVzrQe1tnMY
d71K0KPZ/G0eeti+pgmdUp8ePo2eX0Qeh3WM6ZfNfq8jIrYrI9ghFOUFlgklw6hA
YAhkGX2/Addzj3rBIhhhUI80oX9HAyhc1QVVGkdROBVLh9D0E+Zf1wwsBOYyZWH/
7y/QnBwWom71Ob3D2q1MS1trOvgnhwdDly/QdIPvGoq2Pq3RHwZvs18wskd7rMjO
SEto2TkPApK09eY9RW1lycKF89qtFOGRBzO7St8LP85PP4v8aFXAdnE6Uavxvqj+
L0F2bG/dkLdQilxJ5czakOKlaEk87R6Zp/N5SRk6FwSA8ZOk5NkXPnWicrPxQ5IE
BIjfRw1za1DVZ2MpazJw25vF74MqUpK9qOIP1hT1vt5uJaSXPeWw+1c19Vl9HeLI
SDXteJuVhWYygT07Oz5VkhJC1LJD9RQJWxam8jVBztIbZ3XWotGItTe4Jl2w8uTz
j0uEu7j7fL5HLYBSHtQIUhGxBQNei6ZJTXNYME8qhwtFYh/R8hNve6bB2M3mwLQW
rdcH+DKb26hEYGNu7awsO+7lLw0AKVsFPJAvY6f038M4tDNwrf1tTF2lBcTQApz2
s/SDfXynb5L3N62C6UzMjhHIFvzoJep1pXeUZzOdzbYmA3niyco+aP4KumNb9wmX
e8qikDA6BJdEC4evoJomhAjIfO3PKR7huFkQDnxKVIkL3HQjMKkj96JCNFy9sEcU
Y8j5wjanePzuQGWkmBN2rbdwMQ9mZ4xQG6vzTmJ3LQh4TJKLbLkmRCISN1NgSkKK
vNtYDlF5lHMdnw1EefX5Zizh0squ77i1rcZd2e+8TzF7wK9CYCyh4nhkUsXaP+eD
qXZ6Bq10+e+/12yZLEUbMY4QJT+yI6evTeg16JfLbDVPazji4XjIOse4DO5PwwSd
eKa9eYpGxpAjUEekYdd1Y86SggTZJXo4nbEqrrdrV6P6qGi+Hpg9D01PGaGmTSGQ
E5FqDIBMYoNp+N0z59KqEOoPEVMpX1GSkVGY5SQZxPD/eNO3iHksJGXwA25Suu4L
taDeBteuYiGAct60CQH9RtSApxJ9OTH7sgLUv32EURUoRpbbKWZKLBM4b68N/HA/
SoMNqFO+qxbTRTh1NM2ohepz4Hg1UKj0U64a55EYOkFJswPSX0sU7D9RTz4fJD39
zZLuuMb3B+mnZbBRwCJaW6XsMKwOGLPMI+VJzciWBnAJebkuM6P9oZZLTxGUm/Cg
0oCBesRTN6KbVPgX7Jz16G5944nFa1jU8IJ7qpwAdnXXHZaJ33ARIzwEWsDf0PwZ
+FzUuWpbHS1VGcSIEoDgcFOrRmh0rNkF664jqxbIRIlK6Fwg5VXiMFfUzmKbX6W+
ilR+8NxN6ScHdFHFAg/s7DxIcrtSP8dYgUY51GaVwsx2a5gWT9z/WlMVQqUflM4Z
oztjaxLIpDNAQ5x1JucIh0fnoy3zIEHwuPRn9c5nA+SCg8dCZKyhd6HgkJ2ykrwz
XGXWmJJPUNO2KB9qhjucP9DeU0qqNyGit4u3EvHYvpKiT17Z1/MmsA1AIItdkcxv
WVGBVGchAuwMy0OvD+KdV8VJmBM9LvLDZoPhtDeqLJkTsY2LHhTPP6nZKpub6obo
/eRCbKrlLnF1Wd5kotORwV4StQxPH5nKcrlg9GJcCvt33IseYSypmIm2M0kKGxxw
FJJmLJJlt6hjFC8W5K0Ji/kh3B/Rtmp+GKbpqtSj830BxY07EEPXBoAVUoMH/8an
60MArqj+2xK1hPfxIgemzJ2YPZDYv1n5up6QikPepLPKuQT9NZkR95it05IcZ4R7
W9eMKXlJ2Clxg7D73jtCMNufbXrm4oH+HM2QKcg4tybWjLywz7dXN6rcog1MWwbC
LF3vtwiIXY64OYomICMaZUkxXc02bLLfOYBRgugEi527F7UKVd54cYA4pWLNwg1M
yPfd2Q3rReUtLrTAog4kaVPyFMOALIyeqU7RpsE0Mb+2qb0rcUQK+pVxDb0to3bP
HuaGW9XQrZhqz3k45x/CSjBn7MMOpG2z2W5BkR9jWvsD0kImgD3yL737oxNyFXQl
CPtqBzdNv+60gcY9SAHhHokdN/i2fixdKaLOC/Ph4RqPbg4Vdsvmui2kW5p7yjr2
qsamxy51yBTxtLZzphsdI0kp3QVpcY/rcs009/Qe/D9G6TTVSPXEo3rZFDHSrqpw
g5CoyCAqXVreQffPJS53JPl2r+jCLGL5ApOgN+2QSGWmn7xYBmlgWzvo+y365hFU
0aUXjOvppGAjMIPZt/gVqGMALRGYAOUGADFxcvEO3N+QiELkj7ZFELjU+MfRZFLU
+FDhIOVNqZEAdGIr0aDa+KGg5sbxCO2GtF8ag5tPkXRWORiWdmgsiK058lMeI7Mj
OZ/bqvtqCbrDfveP8l6xHkxOdnEK9C1UHbUgfMNHJvJwqpF963gVyF6A1UeXsu18
UolFcA9qwP02piwyTvbZzA9rCgxFB3I9B/SBOJDjQrwZF6PV89pBAVGfktxxQzJv
Pf40QAGlX6LmjyZsf5GtyBu+5cCNyeRbbqkQ9z9WrkDRTdUKWQnoJT1qzwQ9jdqa
a1oIGB8Oj8bfZasU/R6qlh+wOR4Aqzk9jc0vlI16WVbpOQq+k1clN9vy/xClqZ7o
IL53VApMOlbayO/CiqqwQpgpuz0k1rxPe7uh0ibdjHYM1ipAlYsDjOe3csHTLLHm
46XDMJJlk3w4zlA+4m8+/1c7z93R3th5ZLh7j1JHrl8ZTBGtHohP/gCjRT5hakH2
CHVv9kjP+uWEopdVMoAAXpElStuciT3LQurqeo6F+9qs6MIHXfvT013uQxMtxdrb
jjte5ypYUkIS21Y99hwoGPPiYemdzqq0UC4n3M+sdpNNafL/cpGdA3BgPPDOpwGl
+mwJPFSh5kNpQCuD2YUVN9MKPx5Ws5kS2dnnzgUJIK/Th1Da1PPWb+LP8veKqqJs
mOfE+n1l2Pb9Ew926B/0BACIk4lT97E79/e66wgw55EuklAYxd6RNQCpMPkOm+ct
+6xGJlgXlaHnktulOjBF8HzNI437ddsDjfMoWUjBbsdmJpuisAbq1uAfPd4KNeSl
wPPutLwwPLGGzHhBwn4sdHd2v70urIp9JIaRL+m4pfXzc8yj1VJgejlNdhQR3Zz+
SOym7hnprSrVFwU62N2PI6yaUC/edl0mAlHVJIg02l620kL7m4Lg8a6YC8L+OEtT
OCCpDjOGW5t5UcMFL/OL/ft92shEMKrBW4UHDbYtXU6LL6PbFM13evLDgqKBiYK4
4q9Q4oaRYwHxO6YUfD43z+G19BRAuUaxUGjk9zIL9h6nQVV1fjJdmNrHNq6kdUvy
fTkgvu+nw4OfD9MAA0lSXe6tX98c/FE02BsaGeEKXZJsDKRoqkMa32cKKSAQ3ULr
ILladmqcCEcuIDEGNLfjX2qKzHCsN/vV5NTRAz9Brh64w+mT0TTqbXvGvkkHVPUl
VawrY8Ok+lxiZnVAcnaf1ZWumOOzDzQ+ZbTryDWD0jLAuPekq9cu7n2xPyPUWzv3
BB7lIC5DbyfFVDRkPiYhAAQVH/B5LYkUGheoaFNsTvLGGimwCaHspzaMao0K2PMy
VvPoCd7l9OVkPFCZGAiLciEx4rU1LfrKZTwr91sheOZdiTnQGdupnR14JY5wSh5+
7UcCgyIb1jTYZBSKRtUVCTxO2SI6bA0vU6HCKiMmAVpWe/XGZtu70qH2aJhwTk1m
CBSxG2cu6SrbeV1pqbgqKpCzdmeCVU+qG1katyicl3ZGYMpti7IL8skqqQx5eRVr
ix6nbnmEzsZz4yKviVdartLCn+wSlP44syYcr6VWkwIdtutKbcvAZbsnTbOTkdL9
FfEBAnJfqKM43zVa4yHzTAKVoKsb8WjkGT4oEcz5IPeoZ4RAAe3UHheK1NoAIApH
LWWiH60Tc+0VI7Llxa30gfZYkpb79sPKiUq6VKAKrJHWbdIzpjiIxhO+DWsf7hSV
nqKAI+4lFELaUsbM+WcqBbkubhEgsp3tQDHodM6Kf4K+q7nvhq5jLc0g8a3TolnQ
6vUtcfni9izhj4qot5QDv2Z9d7lp4mQwzpgwWySkpBbrrftbGpHbCgwm9M242ojx
ZhlrEZMKHi2lC01JuoUWbIuZIf5+vvLnGCTR12peQqSYoT/x85ZwPOzy/weIZ4O0
1/E1cBWKRIzK1v5rj7MIfC43n+/RqLhXqHdz53ystP6kv17d2cUOvz4vU9TTvMLt
utv+OPoYnfYb/7TsntDjNu47Svc85DlR5cr+Vvq4XdMUDiAwTIvcKQbneXPgAg5u
P+5aVUcRsISYlR1jWFbF7N1xbNAUG8p1VCB/oXQt1SzpJW9u5ywRN3rr3gpA0Lu8
2k8JSbbw0ar+gppPGkpoLls0m+vWFiPZmS59A/BA1srQqPTj0dh0kS2aa1SqGwIm
n7en81NlCbSxlcGGqhGFsQH+3xiwj2GcugYhthLCJncnn1mwVVE7YsO34SsMwZtR
eZafk3WHdnZipAWL9rh3nV8iYcNEvTG7pLyUtuzuviOzts2bxX2d9iYWRy9GvKx+
QDtMBRlapxAoKBpdO8UmvdqyvPdBcC6ln+VRvL0z1jqHcJ+1ONHqso4traLgQs6l
Zd5zRiWy6Ty6vC4Lqa12+sxp9N/2Qg0BC1++wRyhMks4XH6O0qChM1mQWMzq2Pw2
SP0c9rlEuGC9smqc8EbuZOSweVQNCIrRvRBfOQmZyTu8v+Wv+/aHqviWVFtnmqGs
f1et2vUIKbAHg6RjPa0dajOIbH1GOfEf/rljXzdE9cccCchhEvPf24wTYs5l6xaK
N6ElCbrYSl9EstGfBInzYYHkzvW60tRcnZMK5cgNMCXXAYDEoMy4NKfumbsryc0l
hhC3a6HYmTXRx9vAWaYb+tqvCw2T5d9EM3t+MuRwOF58lZhrWZugnMTG9us8+evn
NDW+h7DvPhkMKFhplAmZyDTuHewqPjhmPLJLQGoElytuGu1hEz5zwsVR+TQVcyed
L1hi+1Y3V2YjoeS+haEOMWNLTYLPlBtLPyjb+Y6DbUgtjIVYcp7kz3Es1n72Z8Nk
9UFm7yoOvVrPeCNbrcMG1uP2eB4+la92/WU7X6tRarRas1+uJcZf5dW8djatjBXf
Adp+RKYPYZDAI05iD0JzClsIRScfJ8FOY00gmiVV+SujPqrA8fHBOAAIZNmGKeH3
oc39Ew2SaQyDn8UkoeyM5ThEqZxeA1RGL4wsYRPgU17GK+d+t+ro47hrpZNAUw1t
1SnC/fRUYoqpybhkSPo2lsrRG+X9dTNwMidEUO0/d6J+oBLeIXFjbYhLzxS/XFXm
HWXI6IGz4xcZlo1+XNdC06lU5SnU3GuNqU+7/NiZBpzLQtpwQhNXzrKbmneaO9qm
twRdfiIfLrnfI3VrUhYUAv4pXsVY+ZEG/CNMAC4LwSDKR6wsakUqYI1TH7SBc12R
pfmlk7FfuuUTi6cKcpVoKavxJNcO8JOPZ1sxhI6oy29Bi3aRxbJ2VTd3N0WzbDt5
dZOZZMXskcl0Uk31W1roMN/GQzp4Rx9Qnij6rAZsi6B13RoJiSqhG0kbljF0wPN1
NuyhNsGtl+LvCFdU5/VIFlbk3UHhFuRfl2HiSO3GK8+Lsaqw6GmXRjgz4Avt+rrj
f9sov9Y+1n+fdd0HFcHTWFpMzJsTFfxw058b2/hdRmNjZ/fkPkyr97HyBSPJliYf
I8O95RM9P9BHUjEMZ2MarDK+fZWp1nbgGtKC1PkpbBQDNSGZSa7v+wGGEG1kWS6M
bdbhfMtXuxQC0eg+BSoq+C2wY1o5I7xfSSgPxrSrh4JR4mFMxM7oiePjEMMM1PkU
odyR9jsssMGOn6+g8RJ7Zd5nom/BhGg+aXalM1Ytj9X5Uu4jmMZPpZOSNW0WqhiA
66RJRPZXBXjZCC+NCzW1PDaTA1rdh0VxbH/ULQv2BWTjlp42sL5apwwyEs9TNSWB
s2g7dzMxWrk7XrwKzBiha5ZcubGdah34Gu/mvfUjC7ipDDOVYeRxol9sPu4TavsL
mNlEtppGQaVj59KFyvheVQQwcFgv9VVTyij0YeySXZjXaR2dWdHlZbZc+q+uWfaH
5JoqPnDwBqqvIvHbvc+CwJ+eqZVqVEB2oOpSGZLu4d9xIqSvTewydqUDozCN8oz6
9ySOTxV3dYbuxx89icmpyko8SePL2SyhyWswnDikyZdABUOI5RrJbVZPbbtSUK54
o4iUmPyRNSDcLGjCWYH2kzyxJV4rNXJ5ctBQcH/Zo158tQwJ6XfE6ffgF+r86OIq
sC/KDSmJygl0vNywn7JrZOgEycjsK7ggA7F7i/yuTLSDs4jWiIi4fzY3ywmv78HV
JbgJrZ/TEomBxT4IhTnPcGQln0TPq34g5ohPZM8Eyh1bsWl4IGUF3j/5C94N824r
5bDB7YsKmmSt328UoWkgg6SxDS1si4a+Wyn5L5o0RGXn+QRjn70P5sOn/QyNwzPU
xpRdLSE8eSxZTUkoM0+F0/zJUZeDPdcfNwsEOFJLV3XK0AzMUR1b1l4wxzrFztfe
NFT/p6h4xvUI9GTPozWwMFqv6ko/CXtfED2x1bLv/krlUi9PZLGErqi5TKwLc1O+
k1vXgeI36+xaZdHyM4Ml94OdJz/nxkTCamJBstyfY3IPNe0N38iGOSkNlRreqsO1
P0KMgi6iIwrceMdy2at2z7sf3rcxhhb9pspxcAtSDbNnHwEdLdn5pP9/SJ+0aClr
kPgceKAIlqnxba8oNhBOLMZJVOPFi9XCculPfKEH86WBTT71rVBWEQG2iApXgeE+
tdEfnOeAB8McZNUlAI8zYiX8ZRyqJMfSRSj2Z9pVbPMH2Equpc7z0ueSq2PN9ecS
1F+jvv/NGLL9/1PKAQXyenT/dQAbmlpkfBkpvJmTPAz6M13Th73/OXeeIHgACokH
M+w465vb1DAju+6m4hAIgcwK9AHRD2wTB2dRH4jVlwsNsXexMInowS93+mezI4s7
CLSWeLSIl9jrxlDpj/TGmQSTamIn90vnMBg+GHyMkcEAPd431umqKJ5PuWo6lODG
v3OcYRrFcSN5K+54/fGZzPblfeL7wcI7Jmb+W6WrY1uFyJok5fQcGqvKO8F0L0Ea
A2gnkGNPcsyuRKaZJk0vlJlEvQD/DqJ/X5XLA9vlMkICC6V7H9EYof2tUJF/lvxD
lZqrygdTyH8ZLQ7Wk5lIzWPuW+4zDNOj4a3HAJvBPL+jGIuLG8dYbzVXAJxykGNA
b6H9BI4/Sr6REYBF01XdL5N4TbzT7GWIx9/je83CkaUIi+Iz7IAwhUIjr6ISeJYf
CO2veo157nGTdWrsLjE1SuvmDyhgNj491l7STsVzUKl4Q+yFwQuWdDAzTIpD70Q1
hWdprlhDwFzjqgi76N9oXcCo3kMZdZa3oZng1je83GQtbDldi/t6n3JJgRM0Hmo7
a+ThgvF+qVjaSnEgXO67n6Up/m/KXeOCuxRD0sdaLaXRcYGZjrnc3nz38tMNjx25
F14OSM5fFvkWwU3qUlqVaMw9N3SOGge9H7AqHV+fV8U6Fo7Z+RGIdb44Z58uwZKK
eICOooiAQgUKq5vEgVhnapz4yacWJ+CDRtS9heZ7HrOZl4ji4aehwBUMpYDjR2Vo
sTcPHv7nZOYzfZgEblSyzZko3i49zsGVYA5ZG8RHWeOMbwUVImbw7/K9NkFH3RE3
QU9iob2S4FWWgd08JAhAm9f30W26lVBMua7P4pk3OlzZDViPqC59NJvldxraobsw
T1IOeYNUdpwBaDYYJeqjwZlnoxnLGq9iraqQXv67Cb0tY2Tme83iiOJLncqPkn7l
9Ch5nEo5Z1IUFXW+4HCm0Ez4VURntK91mRLnDUKCSPOc6xb03qltdmH4XvOqeVmx
gWNhENXrFUGMrHTkgUxMZVOjptVU+QayyJ+Et8UdxpmPnE9rzcRnn9oHqXY+rNjL
XcSieUXkznBfVBRNTY5liko1axRqhT/OiTkLBs9CTwUphsxTzTEaEDNMyGPucRyU
3qO7NJ4NS87R+vGpc0jCRDA2zuwAkQ+ZEJAso8Ot2J8FnEqHZbuYdGyU002+RDc8
MWYhR3CBfwmOBef3e6vtPCwbSEHJCEXynqgROuAs+dDaIbGJZbf6pjZSFS7OUd4H
s1RrhWaCr6sLusCL5ROgjl+i2XLw1H7AYsZTTlFjwBIP4N7zzbTEEzi1wmIxqmSE
10yo+pWriWHJH+AKnW+QJ1q5iDLMlaWsWQxD8jHxXng6EXn5//ll2G5HwLABJpHB
7hmY8NLJd4GqLeBFEfcYI2E+yqLoDUJjCcfaejR9M8SLxjJfDtnSXFG72TvacWdp
wYnN1Ca8Aj6bElEStz7VhLsDZ10AtzoI/zfLJMc/l3Djqp7A1mw0KZ+sOgG1bjZf
LR8lyOW2Oq4FClYnmGNh3WZPvqScunGXR8jEB9AttICSmDRq0LNWtuiHYOWn1ctr
iXxFKuoCmGRuP1LrBIMscbUu/kEWxl/QcS6BocyVb8lGoeNXA9zisI4GrNoh9t2B
LlQQWBUtrFWdPaTc8CHEdWGEMMKtEzYprSJzH5JZojfuL3m7ZqCIl0FWdgzIzdns
M/7BemHtgiZuuG2ceOmr4btT4KhGYRNvdLfax1DPuEsIKN50uITRAwDOrmcX0f3g
vgmntL231J5x2muYyiwqQ5Gdo1s9X/U/RDFFN8NdcoiJRbXFzeDjB6igWhLjoCIe
8eraMLa7bKGKT17pnPIdtvI23zbAbTVvnwX4gpTZAd1sZEqYcM5ReqM1Omy7idss
hvkfIwrgl0gnqGrZLrTIbMLHwGzGFNlBL6a2BRoK/i+EPkBmssR4bf7LWuIc6Dxy
Ie1dRSiHx31uGy6AVhX/4JnK3RCt12y9SzuzhboyD70ZGimZ+prFQ03+TcF4088t
61zjdrszLP/W1KIUnwdxl8dXvCddWsT4A6WXB9jJ0uGcnShpJQ6eo6WROJ1IizCW
MLUkWNBm+Ym5zxLRQJ4j8XXncArWrGBe3ML4aJ88UUhhN84DTVOhZgFiT3X34cNH
kM0zsMYQkYrf6gHHUDJe6lrOVyPpyoMVKqLKnzf6GajvfLh8XNjAXY4rShB6wdBu
FPeXPfQ68n2fOdCqgp66D1jGdmI38eYQEMPdv+XPtzVYk7KwbHoHycNvxST3TrCD
+FKfKRnNFrbYNLkMGyYR8710Po9wAcC0Zv4YN3a1q84MYy3p8pudEFgpuhGlfns1
uSbhfUR/n8Pfna5VVk0L2qjTOqnZ3U6eR5oHY+g54KDpVy5Ji+r9y+nttSNQr1W3
/SnvEL26dvwvkvvkEo/jjCPjm7wIYiXRQLVxgSapp0z/6aI9l+Vgo8K2w4J9yXiK
v3zfbrBoECmolnlt+idb3wxvDwe5Y3cShjJ92nGFklJHZQNHVN9RbmS7yfV8iIHS
Jau30OdmOWshbPiBlYVzeCH5AubQuOgVuBsA3izPXLQVniN0PoE5SbsXmF718dGn
+/Ltbsw51MwMF88CI8+8pXAianKkarRvRdRcLODe7Rr06KPZ4TnfIvrA6MNGIl+4
KklNsCSpZZAwKNJwQRLyE7XVbUtWdEUWzdhn8t1yyTJCINHduzGF756GEOH4c6r5
3LBa+K8rPof1GlJpVqxAkmnBu5xWBJHS2hTFQQnJBQDosKdOA8ho7HT/Lnva3+wb
GIOuMaHf3TgC/DzWxL5it54TNgrUNwRNXrib9owlyVlibEglC7oD3VDoMlrApSzJ
xE3LguINJ03WxxblyyewqXkDIRc930S4P2SJUID2jc1LjXryLoQTjwLGWddw4WJe
8eg6GBNCJ8KqmUzlAuYpjxWB9usfZ3BkTmzRKF7ReVPTl6Yz8pzRQZGFDXRYvcu9
y/3Z0KqHDITbLERXNvbaUFIkm4dO4yjoFeq0QocRgn+Hf+UnA3gLOmRvpYmEPA6H
oM3ncslz3lWpQnOHJszAwciXDP8BBENz1IeaDqNXtoNp8osUWUo1Itgu2OHXvGYq
i8IG1M8RcLN00x9EhrCyiEdBHnhP1KQ597YE6uX4KywOc9Y6j59YS5UGB/lHFhfL
LW/BvxyN6pvpG4VF3XnyiOYqvuKvjoLMeEAVvPbucgsOdTnSXkvKcxRMJOPz/G9V
t0KNpsba9XiJcyKPTR6CdmTdaeXv/OIrwjWhPoXGg0sLxQFM9BOI2E6czKORRC4L
2SEBnsyOlpvQXrIsY/CQUyMINaEqWivJx4ShzjEIfqPqfGYian2v53ILKytK4qk0
u8wvWu+y9EWxmFI04RjQ4TgrIKnJbDiJtqmpdQ9Wjq6Nt6SZIjilEXmMBup98J2M
7mWYPe+y0vzH1DJBcyApFfp0zLPd4O4W9IHR3457xFL3Xj0mi/kW1p7ACL/enPLY
4cZ+cOpfFjPc0iJPbZtrUZY7SdiuBnYo6XjIB4hya0lGuAnhDadSSuO8hKgSg0H9
BG3njlK123ioaVHEUk0tTM0ydaR6jy7mOJRVUV75fLgh0ziYnK3vd0DAhIWxP8rZ
FP4bOr9plFlg5dNHrAPIM7Hr6Sdh0RQqkNUswVBpAHXSNTowYFzy1zwHuc7i1KAQ
Smtw1SJsKMqn9O5A2CIsePOvN1slg8JZq/P+YhNNOBDl/nUzJnmx/zkP8Oj6/x5M
0ZNntl+kdRAbibTpL6UdbiNY7psw/xEljYWoNuhSwV06Ql8lNg4/AsdPry+0zgui
w6a0xSGblo5uZU/Oma0PV42Tv5oG5pjmFnGiyPF8ar9sWF4Xmsb7vdnnLBswtGGu
+sVLALLFcaKelbeoUYYCH/lF4deLBY/CxNFHtyivVAhGM27cKH6V8myvLBYxmXnX
8pwMUbX2wlALPO/9NnsNbP2Q+l8spP1vVPUZt+efqlgruco+Wg/WUjvTcgSawHqd
kZGcIt6Qks0fjVBRUX3BjZDI9qW7nCMTcrXFRtate2gYwTM4i/+pEuR2CpIkkcw0
YR0YBYj9pM5/veSy1+j21sb/8myg1EzSNaSgEwonn6QE3bkaX5CdAd1gV/urjxt6
JL7JOJZkWc50oF5G20Ubvhz8A9V+uamPEkryzEPM+6S90a/0x+dalgeHg4RVnTWf
QfPHONHJ0Kjx0FK2/hpMluawAHkWkAsm4DujU6nSNBjw0KLXtvu4ad5CqSv/705j
c1FpMehhTwuv/En+ap2Kse16lqE9N8JGTO1cxIJR8JUVOnfjGge32wIWJlZDXKTw
2MJlVzH/YvNxaY6gDwSgoolVaO1gHPsoobvQx5O3yF7hZnjFyRRO2+N3El3iCX/Q
v1C4Mr/MtJ2hEZ7jPI0O3gT9Zdeb78qz7R55EZS6ci41zuiKDXeD9ItG3Sw7rKaz
T9X7gM9CbXq2WrUs6YeM81SDPOrKEEFgfgxb8aXtrEXq13msIcEh+kXs8xxv5+Hh
tmY5ILV03UE/gE7h663Zzo32HW+CHXCs5sRiEkKgqD3S0unU7/HBJxMDIB2KuX6g
IQw1ZsBD97jLWMwZw3R+XH27D1kwFc4b5Yf/askvBaHAy/6kRh8Kjp2GayHCay6G
+3yXqkAXChntnand+/NqpUF66OkjIfKrsuee2qjsikxpiqHDw83HDTb9SDD+zdEJ
aSY4WjACiH243e8XIHnNGtP4r3qgviAllP05ZXFBD3jw2mKN+YuN+mMo2bOE3duv
5oKZHtMOrw3ucMYvkEntQG12dZW7zFw4EXDNCfEgr7KYyUH5IjZiAGw7MTjvztPB
ekgX+bxPLL22djRehPbEW0EmA2Of0755FUojboy2H1qEheG/nJrvljMFggiVRKkN
L6RiblZ/ynebU8ZaPoj294NHKScoK7lMWQmrs3KmHLjyzzcE0EFLduzVKOze/dBN
mprIKYG3t4smyKOojH318cxjIUFR+c2GVRq6GFmTll6t9aU9zEJbL1M2lU7qLzMX
Jbvlc9ZDesdktkquohijhCCYr56+jjMV9pcKvHHOKv8C4Do+13+u2ru9jd7p2t9d
Js/6nB2MFaWpYrSk19Mg2ebzQg1cSG9oywLyGpmMucdgn9dDnY05lnpxxNI6jEgF
eeearRp6JK+fKc4Qo+jMicr6UPtte8R/QcWSHBU1FnEAnHffemoWTeSfo5HIhBOY
fZTRKOZAvvKA1Mab0Fqgk7/kB05pU65ZPIBYC0hrSnqcWLNyotLr6PccYA1+a//A
+Bp3EoyCtO16zGr6HVxPWQW5m4HTu7pplrC80NteQVEwQrQMhVP8mu6yflijwMdP
qRDsVcsgifpvX5bG3+r9buMH/hczGk2XkEXPLtNYdFt2uNwMj2S3AT2dQHu/3lgT
FGMhyzyUTuXwPgLGi+RvxzK7b/QEcK0N0XNymssgpmONUoNC0jBoVJdCCIvCH8EQ
TTMhXic6/2lsXjNWr6gNNlDi3EvpV6Rviae89zE/Wf3236BnlpLvpp8Ey68dJM8s
EPmVJ67f8aLGbmgTqx6s2kCJtB12RjkFxcUbsshTj1UsRk5I5Jjio85cCmjCU9dw
eJR/YJ/ekYWix5aeUdGRfHL2QGLRqbid7wGoQf4tL1NeVx6c8Fmy+yexoQjow72t
eITmqD+ZynBqEFbwma19FRFj1DgsElPeFMSh1Suak/UKa5/VJVD9fN3gdgNBphta
ZlIl3ggTY6Sto7cIWNm+ODgDOoaCPeBWF2vRuTo9Kxv4XpmtuF8I9/mT6+6/9v53
xzcwFFbGVcfF9M7zwaIhvoySXN8X8o8v5ol2JLbib4MxumU6jir2e9q5cE107sIO
XtzikEJXmRZij1denRqI0fJtoGflgzc3WtgExZCNr1LojjAV8q4TUo78yw8vzdo/
IW3LIiGGiguGYyvVwPBV1r7Udwqwo/cT5EoLYmkyd0jsIJ87r2JeVM444/FabiqP
+I20AKhpPPOmaA+IU/O4A7FwDc2ed05kAWRMQqiIdXrOEorDSQQu3Z7HUH6M00DA
9BP+vQgPKvWqhfGr9LvB/IkVdrYIL2/MznN/VU1MSFtLxJfPXCP2jCVKqB++8CZ8
qJNl0IBak59IDqE93RiGSAlQJT8Jt9v4zVwvwT7DF/6mJNRKMwAPDP8iSuYJxeYC
xk91gRHbwNekxjTTD9Fqz4yfyPk/sr60z3jV5TNumvnhu81rv8j2Qbyz3BSz3bX3
93FTMn2B1GV3W3c5oxv2dJ5fKoPwb8iPE2jpLMtxee+2GJWhtadAfJ8ox5PV11js
78nIjq4e3g9J24DPPnRxu/V2tdDyI3LVeOX07mnUydsxCl8bo73yuvWu4GZTetZB
rWX1LyP2khW0YaFNw4i7DOaWy2GYOVZZSNdn/zivEYkcjClLa1T5Jm2DQ2aX28Bz
m12d3LDDCLMe7ZI0yUqbAwVJQHLrgV16DdeBN9xEsz6SUUSPkcZ9hFYRmMoZ/Trf
YR9ENL8noyyPZzpvLI+Ra+JD773fwuk5jg/z07HAFz5p0ig6x7NGI4Yu7oLCYBXh
H5sneSEAORGqlke+n57IM0y1lYtKwVhoPf1gS4lqltezm5PZb87zaiIRW1vrDpkz
COGkJ36JiPfZY+D5YLKYD2yd3P6MHOT2aX7FPFPips2+QxWKLVmtyf9ZrQaPIIia
uIHcik2UseoDb2yu+CAFiQbd/+bMWgykgqSoJZ37Ec4tpnTaqAbwOVnBwGFKAq2A
RQcHXQXMvtwIjSZdgFEn2q0Iq+59kW3LoHXKjz6q8W7qz8/cYJY/4NYa+iDj7649
o2nUGhWLdzoMLmB2oqPZIKRxEEy6DY3gwrTvR+x+tuZ/ybOoBnTiwaP0f9dKlIeX
1oZmop7GxI8PjkMeA8nJoMikaCBzq9ZZjhtSPqBaxcMRS6MMogH/IbhCPbw99jpu
0ozsD48CanLb8pk8OTfwrkpb2guRThkf3e77EicWQFzYgFFkUV72bGNSVgwbNxiE
XE2EEv1KL9rebyXHfSFYMALW0a3zveUvxngb7rDURs7zWVSkNCOSqRexx+LxK+jt
bEFvz7wkLZgreKbbZoZRJ3LaMIixQk0/ZzwWybx29H3awOaCNjm6FnB5QQAgEEfk
Dr0JEppa4/hRenMGtYxt1Sf0gVzvPPoGUNCGbtEdhVwccUKeY7PQIxMkfEwQ1Uf7
MKItcZx5VAagEf+zkF53P2iQZ66gdmZH7I2x8Tr0VRfC/GkC/d0FJbp7DLqpo9eb
dujr2Nea04B6j+DclrBswtSTLNrdCQ7ojlZ9DAesNDDt0qupmqaSUieQNMhmHobj
BVLMwV+Ql5dC0sC6Jf2CGdYEaR7cBXNvHZXC/B5oQGkPCWZrVqirmY7YOXhQUTT3
T62CXesmRqiUTOpn8Fv1b2U6jLLRZtNEFeoo5qvDpsBViWleLU1Zxa2hdWVv4htt
8rIdEnVg0//XzLNkMv2KJFgzi4E8DqrVMJcRC2/O6JMrqEK6n4t8JNHgL1egImnq
o8wjwwek5D6sP8BJygL4ShrX6QRPN12ZPtwZC0VMfJii5Y365xGu6twukjQHlHFd
hRJkJQ3Y6W4rKwNrawoURDVDljiN9QjTI0LLW2rTQc21h8e5mRJ8s/CDIDbghK2m
0znDp6haO+iJkMDXAk3u2rTV6OvTA87gRyP6HLPzoF+PFBO0vLERBW+dHmv4ddbb
hJQcnv2rwcYTa8IsKa4Zd3/ctqTnED8Azw5JroKiZFibC71a1mCT6k2SizCRWhnq
2r1mP55yGj4rKFgQSq1cqm598k8TllCM4As4mU6N5IcCDL+k1dAIzb6gy+D/EWfv
lC0WV/en0pXsZQCtc/4vYuPKaChEx0P8azWF7I0FC/2YTd5z3dNXKaW687DUO+BE
9pUb3goTZX/bhaShmphT4P5kr9WloBcJFZvYYe/vK4S3ttwCmzokSN4olILWqNVI
gGnfM/uH6AG+q5opoqsOqcRMZnvBE9eJWv2K01JZ+RWWLMPgir1qG6vXph5VFgqw
b9T/ku1DIu34J/Yj3MEuK2uVNEPtkLa6aGzMQSmSWX+Wi1TP8YVwJvet2eyNQ8TV
SqqXcHBmqQv1CLvjtQy6nDCk2RAnRtyijpufAQlXIivMZIWJqFaoPMAMGH3Pwgz7
dLIM2qqMgDM5Wyb33SOJbO+fYB5UQgc9zBEWCA7+hKCrhHz7iKjglQfvUV2ag56C
Q8qDQxQsfpdmR5KXSuHL9N1dzSAljiv5wcMB8xfYYhMALxnwgAPXffPRcpoYdFNj
uMAWOiE8jwJqZswtn3cirDjsolVg54FlS60nk6lv12TRsTJ+ilu+WDPc6ICX03pm
dMflpKAcZmkVT0S8XV2XDXKUh1YHr2tnl31lYbH/v+6gAQyNYEwO4jQVS0wyzACS
ehrakn4GrNDNlJOOYtV1FMhoFv65+2wbd5in6HgS5iw1vjFFw4y9spWuYXGO+zmg
pcKWkRW0S7LToD/WtSsN3zMmvd2LIr+/FC4tlGBEQhXkXAZzAfV27qR7cxrce7xl
cUg/PutCynrm+xZSM9TuKp8WDU0Nhk9hYI5rz4Bv+sQJon1HZrAsNB0B4t5EqkS4
siGX8yuAJIuU0pSD5B1ro5uqnEBHcSEsajwUb+jtRGPleX8MqFoNuyhdVxavH4n+
rAqlzC1Llpn2ws17c0QCdiMWKjW+JMPoFycEVfvJ8YfM7dWjvKZzhXOyux5gBrhI
`pragma protect end_protected
