// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XQthlZNWbS4UklHWQ/EoioTrvMRn88/FFM9rmCupTix4apsH0WDbLinEl7yJMuNR
apZoGfwSRueZ697kyueRq54x/qT4uKtT33/wMkVHfevFAYw28mvZfNpynqn3RylG
UgHkL0PBm/7d7JO3qCLmjS1LCjzwkDTedcwYa2hVTOE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29056)
82hPmQ3f/ice6u7x70TZ1ziL8jUP/Eo2JP5RJmXHz8lyMT3ztuzLQibru5hmwwyX
IEMiNxPw4PIZ66rKxnWYrUFPd6z+25i2OA0QYifumDexfSVXDKtlwyWyVXH1VpCV
JzooMeguCr6thfPSvohV9N6j7d2gumRC9AKqHvSLjZzA9pE9JQ8/7uwstg8K5qmB
5DNrfRdlNyhBDDOq4/26cY3rCpHhfztJQi1/z/foRGaHZmDvKjSttSE2LgOgWm62
dM5mLgt6Lssbf7m7g18R+GIfVG0VhOQTygbe9nyPnmMo0o+DF00bbygCOzEePKbW
jAvYE/FVVRK0K2RacKZo1uLOWUedhPxFDF6Du97o05uE6dHvfDzEemVAe5J0iPLa
kGwgRSsa930jXci6UDxLPEVcke5878FJQ/+lXkUhxKDX1uS9ptx0MvExD6qTZleg
ZEIP7YdsNd+kVz5vqlobQkGENf5qUZTg1j9WYg526lYCI4hCtKMor5v2VQ9ge6G4
m5vJLanz+yHVVbqM/SIY/E2X1mrpFgYnYgHgz+CU673II/JbFOSjxOHEgMs+HboD
VkDjgLW16xiy/M4lgkdyEHtTv4MSOk/RXHTACxQusk/6pgUN8UqGDgYC+3+6YBIy
YlS7j2y7XFx8m9jij9Mzizz/kWEBPyOks0xHSAdj7m62Nw5YyrI3UOj8lFTPzhP1
U+uqCMSUxNvakx05kgjPgiB0i0TG67gBoHsTu/qzYTsBJ+Zg/gE4R6361xZd2lLn
g21rTq2Lnk3mBx808kRhQcc+vMJy/nriPJ7edgfVMV1abvYMN+FFBCNb2+krBBT5
k400gDxnHbzRvQh1D/O9rgkW97PYe821W7DODRvs31M1WMWfFp1OVcWoUWpMrAOG
ZVAV24uHuX6uS+s/YS1nXqaE/XFvOp9wdcJqvSxvtKWWVA1ySqWfbdWaIqgOLbpI
9OhXfaJ4f78UmtomCuL5cpAt9Zkq2F1iBq8KcJtxI+X37TC03tMbX+BGVvxZgco3
Q/WaM4lZJRIRhksHiEwi4zBIsmoUWLgqddC0UeUPfvoBRUQWoECLrlV+BfDFw5Vw
LH4AgvF42q5GZ2FHHaZxC27ZLp83NKopdpvK0p5LofQnkJmrRaKysuNAZONZdOGC
68NrPfQKc8c2dl8XZyWxKR1DJN9ozm5WWUJqAsIMCKxaAG2+bBmvT/hPZzVGV9RT
uQcsOzDaFhBDOo0PwtqxgI/81IOA1xOvp0By1Xx5/trkepEfApi21l/TtNALTFZC
DSNsWaacyDx8RmsBAqSonYqt1BQViTufnBMT/RNEglLkZfy3Dwn1xJr5Vx+LcU+M
yt7IiIGAgvRHp4XhleXywcqMqFA+l6U9DVh9GF9yoPNV5QzRF2jP67L205YLEqDi
zXgqE4c/aCuMVi4cN6O0dFGsf+qszJZZrjOySB7m8GlhBtLjq+oicdIjM4F/gPRg
biSX1wWWpGjvvYxWCNhDHxDYw+2ZLj4q71L569AS199oxdjeSInZ1WjzYdp4LI1I
QgGqaxlegOM3WXXed/sJVfIpUya/28VZcFAqME5fvM3p9JcMNFMx6TsceNSiPl99
Ksvf89X0xJKMz0PEI3dZiChTC5WkETIh1jLCYbo0cOcq8HMtpu1KnMung3Ctk8R6
XTPCphNTjtgNf/L6l2ib2qhHdVDvmzmGX7rO0TBlwEAqacpxnRTjMmuxaM0sUgw9
kTS4IkCGQL3uDsY1W0j9SQDBquHppL/2ZhcjUuHI98tSrscyQthLJwZqTfNhGOZo
u70S4s8EYD4cHuIr9IsnjYidbwMvV5SZ5xqWJNOZ3RR6AxF9FBIZvzC3FDukRmfl
FoQOxIFLCz01BYJD88IVZ6zOMpyLC6gI6Gj45f1G2F0NVwPU3Pld+zMy9X+Hwjws
DfedtJsFv1hdyeBhdkP6lJYWc5QcXGATZ/53bJ2r5k54QTyiA3Pof9GBbQw6MFeH
v0WRKTWZ9wDymzXUpMHPIBN5BfpM3ek5ehyQ3cXkrMxGPnJGnDsmeDOl1ZQyKjyC
UCHmdkk9CWzXU5qu6J5mI6EBE6o7lAYlJGqi5f5c1z/mx7VqPydJpU/m6cNY4T4x
SjniwIGlVs5MecAhICmNk1GIhbmEqeQ9DJq3s14/XaXzL5zdrYxAcVNWes/voZ7Z
hHWLy7gnVnuH15mOo+tsSn4kGRQG85Urph7xDeXe0BPJGFafFmK9JrMVR8U+TE7D
N6R7+l7RbDGVVM8HM8ZVqnoG5iwGX6GN/XAmWsCzhllxou/yjnEr9AAS4wBJwuWt
VGr8Gg9497Qt7YiDbxOAzQDhtW1p5oRb4Wh6hI/Efjpr81RWvk6powgDSGDC7m+g
5q6BibVLobCohF83suguXJTyg91Hpi+v1aXyJlHHBVANCqU2BQJ4fXWxxC31/iAs
xhTgYgS+gIg9JpPQMYEIdEG/xDT8C11DPChlVF6o3B4VWbMM+NPbRYepeM5D+/jx
Uy/xqi9esiDV8sVojbmWKvg6NF1g1HbymGZO/5Z53nsa9wNVK/knhEpgb7/wLuSe
yRMl+1WB9pxSY7deesNPwPo1F5vjHZIJ47ILDo8bmgFQbeEg12HcVMl0rywYWqkr
nrrkCfy7ps+cqmFvkaautPUTqFMLqOMyjLKA04NsIHaCM1Es4REYcOoY2KUSbc/U
84IHZvUgGlX9ejabtgW4MFXKQh0g7Ultk6E4IHSca5vr+KPv22AgY4xA/6zAip9Z
tjzZQcl2KrgiBd13v8qj9ChG/W0P8Pv1QgZGPotuKTQx3lqOkzy3tHIA+egFQo8g
Wx+Ki0ufO7hOLZ8k2pklf4ME5txRl+SWQm6rjb0pFNcv3eGtVh59oMVcwqrLZBoB
bJMJ7iljgA39HXGmBgN3WkRh0w8YaTv58w3VnTwxe6nNNvJL8HmeMzmwsW6uWujv
NJA5YWhHcuAhGz8PgkVx7hoLSZzXkyK76sBKPIs1ZRaVKnWUS7yLgJy43kIRmm3j
JaAE/TRZ4oW77lbkskS0zDYzul9Qj+wXXA6yYUR21wbDC+9fOOeeQ5aUY5ehZE8O
RsCF+kQgdaN1RoHmS2DjpnM46ofTdKYBaDwjKx/yw6ECFy2i7DaCulEpJIwJWsiH
p3AJvJZXqXJXLupB/IzWBOQqxHh0jiibTKKVH4swFZNHvxhDdIPTrjiuA4WB8Yag
/YU/1LWwRC0zR9S77615rmeyZu9QoOuMweExn9QsQG2h3mzxHDC8X6AgkNo/jmp6
ufxvsWFprxJdrGHKRaXp+J4bZ2xUGTWgS7+yfMcjR4XW5vRNfHx9h+1FfnRRbqT5
kYyHftxAKab3icuKiN6IBu8PZLjmD/imeH483ot41XNtkttDTdZfh09jTj6HkwC+
MT5ICfeHrsYXze9W8PHTj5nhWub/SP4K4VDsAxsvN+FH3lbHCF5tlPw4yayAJIlF
xSxNP7GKHWBmnBMfKkdaoeZHLVoP/jhXgADOKM2o++DXUapriVzJ9Zdr3W7zQdpd
pRj6iHlLCNzAL9TdCumKsR5/2nh1q9x+1boTjT+b+BmP86OtVOEejeRSOPLeE7pF
tdSvfcmd8Yyj1T+fqpKLbaoWBt6gv4E9WVTjOOuMtXjcOqiDfC8ql1FfbK1EoTze
aMhi17qnW2pxJeA/lboGr4Bgr/TAnHKFpKd0D0PGleMlGqiWaqVf+6txChAgVhGu
qj4MpX7jQQc3vo77jidNk8iux7ZTASfqFITqh4KUJgM/1sNqp0cXSGsHyQyxc9oU
yCtBzNFnzhpNVboJzNioGnQGnwMYkIHTpElGZMctFiJ8iAdWcCgUo0mXS4ixVs7p
ou3i4/u+Pwntg4OjC6bnKXUHMye+EL7z6H5xC6tK3Nb1wi0hYe9mKZOBgYGpDZuM
2IoX1sRPpJAaoXMOqNoWFNdDEJOPG0G8RChuPZBJU4DHBczjR0PDrIS7/LKjdBwk
isfu7uIxa5ypbcnnIx7a3l6gnWUTUPy1kgHGl9mQGbq2LO23wxcwXpgG6oY5EwUf
0OJhbFnrMxPlAiL78k2jkYvIq3ABRL9CW5bG3NMdvJCrf8PTXV1oqlCSoRIetZgD
/4SC9mN42j7RjNkM4Ibtos7SxJ/bPmxME74sJj4SA/J/EquFZxieQ766bRZIH617
Gk2RBSS2aRe9HUh68XpUFR1uusoJWha+GSWtUQZfpPdwIAcs5+ofCAY9xfTfHgvz
QS/wnguIvooJ2AJWyfC9n03SGn0G6EOsdA20DWHlgbPx9ln//YTl62itu5JzPSpP
v3V0uSMqNSBpnuKX9pxs/sb3dWWDtiW11/2ykd5Kh9+SY9SxOS16O9OJw6KUf9rY
SQOZXq/R1WTXkGFeo2pcTJyKis8kE6S/piGNPicFP2nOkAUoz5BhKts5/4zrN43S
v5EWfLstc+fvvtO4g7LgzdgygxAjcuoRMcuXRVM5wcZD5MxvAlX2fSZChf+MSjJc
J7Nb7CoMOQvfCfI4cXiX9v+UEWHFOF5tYZ+FcPW5egqP2tC4+7514riJwCQqBEzq
yravVfcy4qt+pV9pfbqFSk0FFfrJzUTXe1nVj0Uva8v9BbwC/Gu//dPdjgppJpTO
zPCL/MHOyHKChDOdylyGqC3Nk085t6NtS4I4wGptL/n3LKMBatvNWniYroiMEg5L
x7vrC38sP6m4lY3Ti9uJSgLodXaLunC4xtALhNWn8TVEPs8GxgpL3LTDbiiHD7sx
dMNn4jsnJk9lrBoyD38NKhtohmaBBHa3lQEcfNP1ZytMW283WX8rxGfKBCb4BMJf
uLPBP3ESZnPZU6O8yU1M4rvezYDQqT4BtIlvRycca0AAhmwouQLms3lTqCGzgmrL
bwFn2Fx3/+/PwxZIPyI1+d+0DHN8PHMlxN5RQXelb0uDaOZRB6AJ7aszNlLqOd8L
q33n9ryHyoEJ+IuLhyAHVnZ9j1/vTc6hLzyDLR7ijEUCq2v7BTsSvqyzqENbhSAa
siCcO48CRYaK7Z5iRmcoD3ijM5ocEfWedCTfcTw4w/CYuMWaGYEy0DXH9CitK7In
e5ADzowXAV1verdLXe3K60eFM9fb/htJWlddo7+wK5t52LF/qFyV/HlReAiCDKrG
5Vb6Z05bJ954hFN/uQ8qM0tE4fPcLJjr+bi4NWMGr4wAUUjvaaXNNQQ7eK+IBBPt
L6UsZdNdKZlvZhvNyjJB99sA4Ef2M5545UHDQSm2t3evYi0aFqgAr4WpUrbp10Fs
TKKROOZU7UOBm/KhyL8Qkv1J6UiYpEkNVkn2mpiMVDY8ExuMJ4wqCZtPFCOqX+Ov
vAX9oFgHLVjz+iPuKTBvO+jLXguLyJzJ4rtp1mV0PEZQMstJnc1mNeYbiEVG5DyC
4zfgz4z6Xu4Ouv/wdmjTb4cG4oHeqqrmCYuze2dtbpJ2ngLT9FExdraD6McZDy3f
h8I9wjnE/kqCeg1sw4nHrQ4K1usqPfha4RLXsbbu9afiC/O4GKA3S/jKO6OSqHN0
NmqgfQ0uBqJ9r/lvelqSl5P6q9Q8FuDV1/utX88kayYWBGn9eFghFZrrKbYz1653
0Qa7wPRmkNgA9vcpJuTFvDAUeyFXbCv9f+ZDA+QFwUYsH34ab+gvHKgGOIdQp5VY
lGN72yckMcONjdFrYedKnOHHex6eiptBQdTSur7wOTebPXgG5fQys275hVjXZqNE
QiJNeg39ux5tC8iBKG21DwoHNoaahs6l2Ll0zjgE/s7o9da6/lvMuxGKv3DBIvb0
yTnvmfsKolJm8MmxPUC08NeJCmJDtBLEyVAlX3lEla6DzbeDfT5oDtC3Ijm/tVFU
GrXC0xF9svuT8cGL1LJB+LRWLhS19EaXi7wmSAVQUx76ciBbZiodL2OFXsuwxh+A
PDIjb10nYgqZHOPlqlI+GGs/YkD6Dm+fhzdg8Aa6Ho7TIT2SiilbvXnOTSJX3QHm
xXfy0A9AfHL1B1K6WRfBerITlnJXqZlVjOwsDHThzY5DOV7D10q5vxbcx2Xm6pKk
+mRLI2KlyVgq9kmlPwrUGmSNaZH4GoZ+nEZ+UIo37kpt1GSFp+vwI4kNW9FHNZ3x
3TmSpggsDbsmGaTR40+15Dk8uH9mQfO6WsAI4GHoguz0cZl64tjlNQS9PqngCWR5
Hwk/RSza4qY4rK7JZL+k+tMittVhDASBco3n5vhYBH60Cnpn6TyHahUsHyebWig6
Ll/w8Y8db49mCePmbrJVO7zPBqu0VtBx9WVBfxA8igNgkZ8LyEFbBPa99FZ5dwV6
yqRld9AvJz1jm/jR1S7vOnXO28ia5/Ku4NGSmy+TNgxlGrq+h8T90qzOtjMxPCiQ
goR5OssH6g/D7UPeG8ciWcz57itKvohL1dtzsqi4PzPXAQHyH7x3pp7fm13x2IIc
xQJfDPoQO+zCF4myQ44lq6+GA9qH22q6wvDQUw/Xci9qkIy/FTe1tIagSkpvgtfN
QmJYGtVliQIvVp0FomD9puTjtUSr+NOPEaSKx3U895JK+8JW2n7/GPBRNJK5u77V
6U6FTKrnchnDMMszr/nXc7JLv2WgeO2LDRpQhSRVrIBJH7UpQPx0NjTrqresSfFn
HUUbv2m9v44uik4MpEMPOpP4xF8XT0ENNK19/zTY0AQFI5NJEAQLQwreSYlhSVKL
3B+mLlha4IpWAQkcAWKHkIL8fJ8jOUD3TQ6tZsBvbQQOdswZTTOBctXeAhqAzstM
sDxHmzwTMfm6VRl+QatUQlGksnpM2OWRlOLGqk+Z9nUJeAVH029L2bTA5aiNx5Ze
Xp0DvMRS8OAc6LJbwuxW4IEkW+IGkbkPQreW5X4DvpZYHMyHuL0LXtgG23SLXDWW
Nk4Ty6hFSy33BqVRK+jXoPNfW75H11F68qxIBFTEXe/WxTPW47lldRGj0MgY1M28
aZIy7Ibkilp30FZW9MvvUxjA3ulbUb4jKqnr+f0XGkvVH+Ci8rPYbCR4ciqJoily
2N3HkiQ7aEguERcE7RonrYr+95TspbigWGpjh2QD4E11sTFAgvHbSOCAL/Ryag6T
aZsHo5CWEmxSY44g2eAvfXQBndHW0RGEdyUbW9bxf4BBDShhCt00wDzxrJYt4ero
IR1AlfOVokEiIXSLTkcK5lwnRnNUuFBI+GqtXGrsIVh57ljLvItvUAmAm25XGHP7
mH4VaEbKIyXaacbJL6ZMLIvn2h+AhewTCOMxSxbrXe4JoSLGAzms5+ym0EPyjonG
NVEXLjynJv7Lzn8XToI1loCZFC7TU1CbnCIfIx6cLQAJGMUFPsRnpExe4jPkmUxy
p54PfkTkW/xSXJ4ro4Lctg4qxjy25YqpZnfDOfWCWjyH8959Fxf3YoujpfpfN25h
91X7Q82NEHgFMlvCaINQ7sw3h06RI3RFdktD712Js0q8t+v0vTW8ZhKJ+ikDU/h2
xolW318WbooROnl7+5EIUl7eXDJwn2d31HlyX3K1WrBVKKpRo8iiFaEXzrNA+XKC
fX7/B/jOjuBJ0vvZfRDPwreRJ8kYIIL5pEqLolK9RgtUC0A3ne2mLdMnIDGBEoiD
Y83yKpT6j6TsgYFH5tpdiLslbzZ31ni+FRKflnb61yeAVIcn000qg1U5rxqwAq7u
SGzDAJ+9znghidjq+OQfkqAiDQPERkNYk97Q3cyjOO/6FV6RYuwieMZdkqzrGV7T
IdXG4rJqx9DrATkIbtOhq4JP4f6TH6J99Fh7WE1wpfQr4VQDCAeiUBmt/7OWdc6m
W8Wud3xWJu3EpDwqBKN6R5er2cd/ifUjP9Irydtwu6nhO08NLJPhIr/nlcs029K2
s8MtgmKqbhDi+KtDXTkdL+3cFwTPYgdeNwQTtVtp+7YsPhEJI7el4Sp1UK7ELVE9
pFN+YiuekhM0Gf0F+Guadn3KxpfXO5ZLjTogzF1LiE6R23vPKxkOXIDTkJktx95Q
ygXLtpL+21aIES+uvMHyJVUKW4r2T+vzAllA8XHYWW8iPmmaF0mBizYQNNKDFviv
ElnBfsO6Fm2QVHb2kOWTTGwD7ZpRwNgXQ+0LecvBTWJMjLodVF2mWiaNir9wcNUd
GxW6X5hCfSUBdffnFaxj02YEKRlRIF0ZyIQuqEEkrOaTUXzZOBzjaVAXcEN84vcW
ffh8S9jMLBX0dNHMluV1opInVOZsorYUI47A4dVPzUY7RAJ//zB5A+GUEXB2/uB/
YwA1SkYGrkRZ29wsjwRLTczuQcKZBDyR5DtSXntmtBa8IJ9daVgbuCuapup85tmB
yRnQAAYpUWMJo6FTqbRr7ZMU86yKO+siu2X9hZjknDBCfhkMnEyJW/xdqcTt4HHj
kgvP00YJNv66PUUvk+dGt6zq2r2BSidW0vFknR93A1ZTzB2HeCU14CPE/8Mnq8gG
uGog2oMPM8cL7K6X1r4JZJdqEsMFMNkfp0Q8e+IS4mQ4BTlEzdLhr422c6qNtF2R
4KRJ+QVRgQqCKh0N4TsDzWFcXcNJteLwGQqqUmwK2nWxmLVNd3uNOk+Xd4s+Kjjc
1fs6EiDIDG0nWA8Y4UCpmYDA6x9WX/7wRbwYCAA/bx35EdeeMKsSVo+Ou2y4Wqsg
zj6KyAFky9zYhSysDipCMia+OzKfnbJcSqE46RiXjfZP/L8ptw1GygYm7a2KLjCZ
EAphpGtp4M1Dsd6ll7WBQ+s9gJ507BmirZHeLd6fhADis5diyCLbSkPY4xj6KTX7
YfQ5A1VCSWibdwri+XggPF6xsw8yKcfyZ9gJG1eMidPguhMl3q+p7q20FDoVG/a7
9bqVMSgIu8QduAgO0ZYvF0hhxSS/KZIHv7CKkcMVNKOidhxNMzxGk7TAB/KZntuI
YyB2Coa2M8wZwJLT7jet1QY2JS69fEtwjD45vam2e3iw6WQEEBD4GodHvPrt+mJb
KCcYFH0AjZ6hbm9yfBcu/8Q/wtjDqEcL/JjgP4pWJxFUMPERs+K/9+GFzeIQnD7Z
59IlIUAoDM/CQRW4szGQKIXxQIB2k78lxdF/W0fVQs9VU6FIyuSe0iia8CLG4boD
4zQRPf1PeI5OP1eq3PfcVCvMl3nZyqtyDihYeXGvNg+MPj4tfFqGL7Om2UhVwhyo
Lp8/86z6vGV/jG1L5qpJOpkp0IRB4WYgtnvdEfKLEe7vqe+0NG5ue9hZrfQc8Z6R
bFkED6o+MhIdzC306HlbhvdlqvXqEttmP34l9cBCTU/mhsKRqpBqYhayyssX5rh/
zJ1HQ4mMljkX3AGuAGcHM6yn2vtUOf7FRvL7piDA5B8O1oGUmbNhYadVjRU3kgrv
k0k14Fu5KVZCCtzHdOO90DAbjRYXb23Q+9qRmN1lpG50irPItStlknG0eoo2dExn
fmIXQKP9XplXvXMMw5Ep4pHVWafaDtkf0vMRyOuMqVeZarJCmA3jJ2JorgxebtlQ
P6/W8g6ZxMUZuhBk1clqFdjTfbkUdmMgTfEIQ8Ti/U44NB+n11/JCXfQA6R83/XK
MwDCyQwcbHqcUDObbynxJrtYmJwjZ0FCWRmzKCE1fz032qzj8+YQTzVOjGZpP6lZ
/o8Lbubzt3jNXlGct3xxnqqiOtfWhvJgjhMeQ2p9BRJ0MNZkSceF4bzi01dxrmz/
uFIcK7hmnr64NjLcEqg73jllG1+pXpVu104a8kcRPwTv4Uac2MfMunXjYDRoRm6y
akN68a+Ql1s3tUy0wx2/lcYxr8IG1v5+qnsSxWhQN5EJk4fNjKnA5PdTblUKoAtM
aKHZemki/WfvpJj5DhPi5KcATTlUnND1mwBI8u2UX8UxJAM7vGBv0KEm8diawoF8
HBMbTe1plP0bOmZS90/AX22AJulGz49WmDby/1nKKLaXxwlGrmZYEzCUuAsbMSBN
ikAkWBrDf9XIRgAGGuyi9uEJinv9aEdNheluXkL7LQgvbazOPrtQkoEcRHrZBEqe
red10DFR4Sy7w2pJ2UnaBlHXXaCDFH+ZbryfSLAqxW/GzIXAKILGq2uZ7QsEo4LM
+BUmV0eBiK53WxINzmAQBMohcwdJ3DWWrEZgikLdf6koH/4spu+BUwmN8ML2CJKX
zymRQHQLOGHw8qv3XCX7NxXynwujrhiZFfyqswfX+L+n9RmRQCuns4ea4ZXFoEQn
z1GTcu3MGwRrtRr+UB1mrha4pGMdQXjIWm+ESqkq7XXoi7wUNHlvrmLFx7swPJ7a
aShMYfbmMeq+MAyCaIGQ5kDzuhQVpjvLW7YS5vgaJMqNTqQrk9jEZMZ/4qOd+nEt
/1m37jcVEvJI8g/Y1eXODUa7eEjeyw2R2lCZ1wELyBdITIRehzZA3RTFIjrqr2XY
jtjfeSkE9MbBXsMgzLlX71Nmk5iy39LEsJMIoRTT5xo6IWKJafRv+AiGEsa38gNh
LlwIatc5XLQMPLjcckl91y+9ze9B44/oLF/f0EOXxUXCoLWt5w4dNzMHh2uy/VCo
yiPWeUf4w8Ei84PhRXp0ANC4dM0npE5KDce3rb/SRel2FVLcIjQVXmQblLAU5PZb
a6UqFzjgqlrjulk7aXDXrYIewymATvw6j2qqoME1EKaeYuLYdFXP0nDeINtJRvvh
LO4C3n5cKuUuphZObnHdVhmDrAWnGXVRNUEsAIWgr2FTMfHgAquKCrcIJzAYlY0g
Ub+omdsCXIsCtNFdtpHTssdsoJJBZGYHELzbmeJAHNJkzemnS+Qsw+cb6+1cglAU
jXR0Trhqc7JSPyTQevn79PTh5hFUN8Ayqiq65EGNZQUokhIpwnAYv6Bc61S0xKLN
qlLtUKrb60FyCY9UBgXamAQNBmBOm5n4Mb41OqUFGcVOYNRckTmk9T9X7s0T0yvl
9Z2IXZSPx5Tp6ZOTve52BrScKyD9HAwTohCOVmCUAqlGxJY4mL/RVVEP8bTV/mgx
fCLOyK88LkIlCAQC1fBqB4QF5z6qt1K6p8jESbEGMjiiRaEgSltP/w/M5kldXLXJ
Sx0dmd+ZKJJULRVFAudJDOzg2yt9esRX7Z/0hnJCcjS55YqJuOKQfdfKrCt5JnxX
Y4w4ki2XfFCo3wx8SmA2znMJIlXqnY7Ry1rT08HWNbBaGIgUf6QqkaE6waTGsHKG
ZszmQ5nytUpQa+drSgeMeZmLUvXXqFwfvasm+Ncd2L3QrqfPkEWQ0fXGbcQ6HwNP
+2LEJswKeBNd5DqOiL62/9eXgucN4x/HaqIYaTyK4YxUTaZ77N1P7NErDNWKg4Nq
LFnnbmnjdU1z217H0Zwjcfg7m4eWPP4p4M1lX5oKOH/yIhFIK2ZV3uOaHbxK8LeQ
Tg5d0VUR5qjV6WnLuduPWJcKHxIY4Pe83wTcJRwbnHmFQ2jVdREFZ1cETRbv/61d
s9nUCZ4N1LDdglT8xOyFCaEwyoqTT8wBPqttyBwmigtR0gqYU7WNEhj2A5AGwY2v
/fkd31RMefNo/28++1gw3yzhlX/33mRuyLDnba/bfo2qieTQ03xo2PEHFh19FL1i
141jAYed2fu2uRypbBB1k0OYMozqmQfY9YSpuVegXgr6nj3icleVMek3DaDITpBo
WubMt0fu0ij+0ZoRjqU2fS5dEV1Ob1kgEGm/UWJ5kbQGTAlK2tPagrJx3531M4oV
XY7M0KcVYBAIYjkMj0w5CqoxzWKWki599gZZgTNFrRpm0/j1bCM6BABmViO1JC22
HSO9y6pre2j0hTO53/ii7gGKDDPNZTkU8boy6DbHEC1VmZxhbdIAtyOlfXKnqWXA
Zeo/yVxs9OWCmhve+/SHlAqVF9pPpZ57b6Yi3Du2Ro4hgXnThcJK1OQ3IMV0R9f1
Gm6O6LfH+ZtZe3nWy4/plqBVFXLsQ/MRBDA3htDfl4Oqng86r7PTqp+mvHUVY3Kz
6axQ5TXgyywJ53/9rpbESyjLQfAZOlQwXlmey2D9hw96pl881qGAH0WvJaG5VvYk
PBt4/PSTQboll/AL2y+o6gbdohg7emtFkRc4VKKOsrX8AY9KjTZhIIA40NxwIj+C
Lx9xYOEFcOZFM4O3dahaib2KsfWP/b1SVmZqiDsqrG+iNZGpaEVKscX8XAwykLQf
t/b+sZKLnVkOG39M5Vu9BvFDA4LJZuhEfauDY0SZhhOoRV5EyDGRmTBjkPrBt38y
g57/DY0ewVm6mFoLuU2kyWYIbacZwyC+9L1WuO8eyMDMZWGcAlQIwwnTVPQcVxLq
SJOXl502sfZZj8wOEW7RIM3qh7FWXBgRLXaMvi3Vvx0iwqkHqwehqnKM3mTTO+Z5
xHjUlTNcIZpVnK/crDJ4yv1teJAmmcdr373NS0ygPtOF/iChCZ0NNknMiCV1TcXz
/gCREWa2wF5K1afs9TRdGz/ggP9KRKPu3ffHLdtgHp1PW6DnEoisBDvLeaqY/pWS
9XZraH1HmNgNfaaM1OGlidXY8XOFXzdWHaYU1bxsD36j1BHI29BkoyiLUdWqv6gG
LXjJttdWfCfMv5/blLB5s7MuKVm3xrPItm0NgcDxlTnC/ogCN17TiAD/bdkhjpqp
A+UE5QOG8Z8B8/uUk/99Y4xmJMTwxL7fJ0RLEjN+jzqgOPqYl0/tw2M2UZCdM9Xv
mXaQ5CP8vCP3BY8XyfD7WzylkFHU7UBKwcdWNwBDa4Ejp2BnUEqTmO6kpDdPBPzH
14NIsugVkAND7hKUnJkotLvLn5QxqXBjqqYnjiRWnj4Sln0az9wm4YyUxCp27ONg
cP4YtUVx0LHQ8OFtKbHMDxHFvPhYGkxBVQ+TEHr7A9xsCnl1icnX3iQQB7hx4g23
PEJ+hU45JlYNJppgmOX6kJTxQ3piTktZevzF0GY6tj0Kt0ynu4YaOn0AjNTtrBNL
hFw4tDKTCXR5FYU28IVLim0uSbAbxgzYNk4oNKcLvKRkiqdWAryMxbjz58btph1B
RxZOu2I6JJxhHBOftqRQQfXO4aBP8vDVLWxXTQ/uHVxxU1smYqnl8RIg0ybSt673
NImRDkeKqVOZzw6l9sSiljNgTNxEY1y6VJJmaAyimA+Be/4svjyq0q3NG+T2sIRe
oihjXzSJUfkT9G7pLMlY9UZ3hZ6w6hkg0w4PD9EbUBX2jEj2zXf+0lke5pNO4E4F
z+noy3TuWznXBBPEJzStiey0ErIDm3NqSH0sCdUUKpsFUnL2kQeTO+y1drbJ/WUj
Qa4zMWliOqT1OuWZZ/AFz7aIdfhAdmnScfGNDitSbWp0JfHKEhbDU2SwT0ybZWEB
NWCSDHM0McD/vNwA9ucYxRm1OoRpqJXueP0YqoJDHRDAUC8noRAJ7rpfF105mlWv
aeLBXoF9z+71Wdj5I7UbUvsxxq5a+aO1mNTn+m6OvpddXMx0kXye3JpSVYkR/S+3
MWNvtfwqDssVy0rEx4lCZgMSQanrHmvAP8CmKyNmG3SJn5Sb6SmWS6N+63EZBDsz
V2v9+Jq2po6YoTnqTdIzrEgvQwTc6rnpkR8f8hdd5mYSTC9tRYTct0WcSbWXTlof
nv7GcJZHHvyQApEeo38SIrdRAxcK1Kf7GCfXi9rW5rSZUcg7m0XgOtm2lNn0yyp4
HTWa7jjxGKuKYA0CF42Sc4JgMUFgQuTrxDIjflhdWaSW0MKSyvhJsTQnz0uxlxXQ
6k3mw3cybBR1qxwWBxEEOVtD4jcGa2MsOcs0yuVYZKq696XLmauBv2yLktIeVHRM
bbB62JZ9PqUI4YFbvDdsU2f0swMgrn59+eM5AYLfPBh0XTYj8v6cbKKO49Yf4CWV
TNd7lMRnqzTQj1mPZ5Iw0jQGZJw7gj1Ww7r+Fhwq+81QQQIHJWhfCKmJTeKouzhZ
s9NkaTYxdONpSNjzxNKWjSRsLF/3xCMYI8S7orIKRXbhPi1ShGx3SLotxMRBuli6
yicUkB5LjoP70hKw/PsrW4DZ1zgYXlLJR+2z2QN0UMBuUZV3U8tEnV3CdeNXHevi
wIviOvMu7IP/V40euC6Mf28S69uTCSx8dAl4KML26WvbRfTW/zBwHpsuhvViiogH
F6hHOaoEmQ+8wl82WuipTDUDyD8m4rSbrbRaJwY8OfpWGhBUCJQw1ngu7AesWgVz
XneqR+NTm+sI75R+dleQuhHp3W2LMf0IWfhB6fOFoaRPmHv5tUA5VrJVmvtO6yIG
dwKojkPGj+2a/sOHAyAzDko6ejUkXHkElUS/g1J6ugNysKg3j+lc6kNRgOS1nQ1U
krTZozi2wrQa4EdBnJPFWyFbQhWHTJl5dYfPeuitthO7IeRso85I6swndgGltwIf
8CsIVm0aRZynAbT1w4mcm5SoAH3mV/eY/9WGg7m9zXWIQTuRWK2AxV/pdqGUPjSb
GDzkLkLLEVrePyJ0/86Xet73Z86g41g5+Jy3YM0ni584Lr6iS/58TAgPY+aHM3uk
fgEvm3BBPgRxJ/lS8K82aKDf5NCYvaHk3BmUfpUpBw7FJ6dQdmet5BVpU8t817eV
E2YLrfguxLztI0Zn+LrE+MZDmqjX0yo1DgFJEcBrtKMAmKIuFCmIDZXXQuWOfSW5
HaRVz7MWHGk/Z681gyuuQks4bqQfdBIsrL7H26Y8wFUPXon1IcpgKuH0UYG2j0pU
TTbKgpVdN1/OUyeBJ3/fgFMrWTroGbEqqF9KrEQbr6vZ9PWpFl1Y1GklHNQH82uy
WK996OIQtQEE7pjHS3WMk4Gmnl31+kRoFdLXJ/qepKhUkAbwPasNFMjXsX7FKe2g
WVLatFiE1kwSuJwY7zFXaK2bE6Y+eYv4rDoZJW3PmyolQA3y062YHpsgXcDqvJXG
oOFw1QJeuiEvr9GYPR2vA5w0drf7HbdUJycT5IBAo8oBKEnJ2lKA7bvRk/bd8pXS
lqA2SQlhX7BNzDfGjMsopOnA1AXaVzgEKZU/ya3bhGaxg4B0nMcGJXbl2s1M9Fzv
8f5Fp2GmdKLIg28AawmHlOtl4+yHaBqhUEtI59pr5gD9VNvPFEl8iDTDoCbptJ6f
UK6EhJYMGDC1rjdc95OkHPGQqbJg7KttC3ZqpwnQu5BSu+q1C6+tdIp+lVWm0yDL
KIN+23rPxTUQj5IhSUKZyGM2X4j9q/pQQI+dl9nLQsjRk1j2T2vWxELiFqGJBPrT
2ISLLIvLecLVQgkavpyN9lRRaMdOnP9Ui5QbxUjVl/ur6sQ586Ugs+UOiMdbB6f6
N7rEexq8P6/F37Gt6CbOguDALpIQPrGdehlffFPA1AzXvsIEatneehoaG/bco3lJ
rmPRIYqDxwi1VXSlaj7IlSFHAP0EMRLc21xKR2xY0OpHeOMKWeWOGR6/LjfEcS08
Y0werkRBDBOf0DoB+wgIlXBVsySUSxRAdMaShPK7GoonZRCRR+9SXpoocW8Kkj8E
WLR/SV28AQ18iXFDx2nhIh+z2Wg6AZKoUPmSTc3CqnEtwd9Ve01+2ABS5HBZSqFR
dHrOWsXF+90VFklRk+h6RyB+ELA29EKH6Kgg+2/qN63v4NTxNNmGRAS/R9I68Q1h
wgpYS7/w22eTUbVGGYBsMeascu97ryzhiRjCw6iol25lgewSV4a1MpIXQPnbDq+D
OmDUj1d9tKWYuUMHu0BLWTZmAa9mC6F093bvuzU1+CXtS846xQsLywfljDzisAyM
IgJfaTdrtbUISvjoHUTaLxY5wLxNeXQC/x9mxTORXNGfPJMYA695n+hL17pKy/wD
2UBySGWtCxYGnL322EfZS/m6r+yoBxe/8Qua1UoVpya5ptI9YKBi7500raAybmux
WBpvZhUPwcw/0DsEwHX3E4Hx8tDEtKbzEz9G7JK8XkfMu3JsMqraw1CFGfa/6sSy
zNlMagcZEfZs2n2CP/hDRr1fk1dLnrV0rtH8edfw/bDBZtg7m0r19KzqOxg7k8/K
Y2JLsUoKgJIxRW05nu1U2UaYHJpdOkX7dNxcQLNNH+lKl9OrcARvbWqaYPpoiz/+
a3CNW0K9JhonxAY6VWYO9ZiOPk1RRQiuXJhn6jkh/QhbwTmXABYpPzhe2/UMjCV4
R++VlpiT2sQdqpsAEXe7zBsbNAQ0YtWIASuMAi5Sdvoo1dIa6hX3EJIixcohOeSA
S0qKuGn6ci+r+9ikpV2lzS6Fxjgi9u5nfBRxgey2uf9Wkg7THfRzJUXRXDr8JZBz
q4hpfCpKn01mQWB3lw7maVUQfFGRj25En9gnX73zNA26ZdHnup+vzxeuamjl7RxI
GVbiEGWNgkLD3O+TTPon6aiRBW2sBd5B7VL1TiRAMYx+WLsIMzLOkfHXg0SBv9O9
1fln7+CR5quf/9sGT9MHl1dcpSR+ev99533WSpYfBJ6QayJSg4+jF7ghTfdfqTqM
sGuRt/oXeP9GcnyJyNZCYfXM6u7vdFN9DdazJeNNf53ezkrTb+7hBiarwQs2pr0+
LrD3N3fLY/qkadji/4mcsB3lHZiTZhf1ggOPRnsPIX/QV/rgkLoGvuJQu+qLfAHv
DUnJJ9hGUV+siUIkYIJjIVURjgEXvqnNlVebj9S7eBaM0EtAFp1OSIfXXso01jjo
30dqpTk+cAwcrCxaALruknqvMhEvxBvTSJtGBDsRnpw1R1T1FlNVsLV+j/wQB/je
E4TcJ4JblTDtWkVk97iSv9Fdk6BmivDxcjOEAWX79OAjIVdMRKv0eMqNC/uGIG1b
xryxEW0bHvtyUB4D5QGt1dcKTesoNQHseOT1flyq9T94HaYn9mLEjoSrCVeaMjdf
rxeVAcaCD9H4od6ztk7tpH0c+WUUXx7HJRp4ZhgHOR/F9Bm64borc14GUlJ/8fgj
G/K0uetOgQtK758dQyozgz0VZOH8vO7qxjeiyThkxI/1o+i+JzzW4TnO1NW/8XSy
Be72A5a2HzxGVqeSWmaGBFdHuSR6j3rSEuusERKim+t5Tyf0zFJdU4Gj9+HbZ5aU
2SLF0//RlBjjikIN0bgaT7WrSB3m4BjwbZzaWEqwLDcrrPqSrDVmwbDG6ygVZZiH
gVn9Pgz24wAuvCOP0pKW0OCeziDBkkuHG5UamRJQHks+/5xWKGZolR2REDGO6f7x
jKRcwMoGd8zmKQIA39cakfOZUSUllLrZsTRO04BTBp3Pon+PZhTCAHCWfOijnbm8
yCT+dMWFF0+PGUhXP/SBbMHfanyJTFcZPi1al2VUkHvVjQ8hIpeOu2jNXiClLY6f
NFM56HAmAbS18RCaX93AJIvlIB3M5JszKZeI0rM2J2Or24zfQWzIhfB/FJCC81yO
OP75PqtuhlNxoSqWQ3CLf3b/JiVF1hjR9au8fmetxfNparp9PUlA/sCyZ8eo3dax
Ts0H2WY2aab634R4A3ckPtLQ0jCNlP9dUaMq92KGFGxkgyc/AYNxfDIcPVv1lAaq
xdaF63UBYSOUw33mC8vNbwUYWzU/Yrjz4zKpiNGm1M+ImepVReApAS5Q+AHwfSLv
mtj7D6nOigfES46o1zC5EoEayrkSNXXy8jzn9Q4NUi4Nrr4iMxA+KEVuclo05Ryh
tALwlihgylWhnenE1B9R+bU0NwtYjARNbnTwIJWgEIWpXgk+C14GdeVq/qyUnR5q
Uax2YRWRMiK7ReD3xbiQaVkZxfwXr6nxJJmuVIqM39gLJDzuvszZtAe4yLL7AaWW
UQG/4m6wog7lmWoRLmJBcnxXiNSWfMGBYLZn5lyP4seGPDlB0zSVWhyiuvcAjtGF
gboHTIVsc/+pwO8mSNiJQE2re0DGFHjVHvZoBi3GRUBisYMga2nOxrclGiCp144n
vVwHxUWu0Bz63Q8HQ2A758ktkVvAJ5Uh/w+KzOYfPwHHYivKNa1q/FI6n3RMJ+yt
4x9oooE+/GRVvDPbn22DXOs0rv7GMJzk4UcGbhqFNUICYmwU6kTXJHgG2yuEjSLo
Ai2vPoAj2kAfV41WBgxv4JUyWi+1ukp694tqIeBrkzzzGMlL2ZR/dzJDiI7i8kT2
cbDrVMLzux+uJsFKOrzvhzgUN5xVXwi4t1M9bAlYZGMFupIescG1q5TMiD572C2H
/konZ7KfVF3VJZqDhEOgo2HZEY1ZKUVKdUT8m4gFq0naLFFUzGdaoqFaBQD0mSun
Lqp84RX7jHOQIYxwVIb/DoNx2CZJ9TCzmuOe3xLjawFO09SD/FDKVnRf/T6gWWqc
JkKbR+1EkBQpnAQ1kV4i5ovJb0ierK0TMTcSG4MTxu78K61dDsfhr+qZlugRqw0B
OQg2Vw7ke6/fMzl4/GqBNzuNir9UAJVoYtl9Sbw9rZ/oHO9h9v45e1qluxIKDd3e
npKlTeq7M1Y/gYb+MDJmdXnC19RqX8GhwVkmW0+PNIq59Ztzg791hyJG7eUy34QN
cvduAvQu9Gm6DthLHIvAjkRjcfVEMrfzNgo+Ly7q6e22L31bqHd7xpHciD4bydxy
FDn5kTKRwoLUDB49nhND1JsBUCfXoqneKvuiMlioSRpBNTRGAeccnBoK/D0gUhUc
ZVhAojzOPiLfN4Vn42ZPQndL/lkNol9iTxFnwjGhTNqbvva5Bx8bdQIIfh89cKHk
fKlWDKazZYH/ErO7aKBlCTIx+z0ztTYZ4CB8V1DYwdTHgKhsVEYXZM+bY5/6YXbY
nJWLS+0zWutRwUs0QiCcEJikPQxnAwCBre7U5Ab2NPaQyh98L4pUQBLp1NfPmc1a
ysB7mxdbLQiYG0cgYBJSdHJrV3hlS/tfYoZfLW2cbmU/yd9dRMZGkw3tk2p5YPDf
X6J0+kz/kaawThxmXwoqvxtQiuss72sVrD/NRxC01gY1T8t1Ne1ARJgwZmzuihQG
MuN6XPfZTh3iqx8sjCMQzlM8q4mkuY+/bPDEks/4mK5z+0UMmrRFXPpG2s+Wtx67
hwuM5EghM5GlDTNBGd1IweX09G7nLLd+gI3mzhYQTbjgGbnZ4uZirnNo9lXPxU4S
VIRe/KuZXgGbEuljoJTk0R6UcVXqVLv8tJMUboVbtRcfd1l/PyP+Tli6Xqz6u4TQ
diPsuT05yLEs405YDS5RCyO9TtjtSs//yoBa1rTGmYB3kyQtUt7h3tNewAn4URQs
HDyMgrc1HkAw2RhJfWt/jF7x6hOlqnr7Sg11M4GG+eLTPw+hra7PWUymyqgd9fkR
lLrTj2zoW46FjY2RSvcOxKYJl+0iIymdzQAFaQd+OrE0LMKel4Eq8wPDhZKpCjTB
5E5LwDw7cH3hJZhluLSKQSij5DiwIYRXDSZ+OsuUehaXTDmHcyr8vcH7eU4BeIby
+EkLKNNQUUADDTK7G9m+2tCtnHMuXdqRelHfagHApzb5osroPXMC4KNIei6U6Btl
ZpMQtNjbR7fMDgwaDlAw3u18frTc9XmH8NZ6y7RKozgVMg/TInufhNQrEXLVIoV7
QT7zBB9fjQ7Xc+Hxfn7YeJgH/IbydVURBVPOr/Xissq4cQ/FizHGDiURw0LDFvXi
h8kQjdNXc1BRhV1htGfp/yCVBM6SH8WBK20TZG78H+F+hTvDymug0PP3FQ/vOoP6
/+FEv+tcC1X73/T1qy8WMyxaJRKKx+tajbayE20BDeATbIT5CZAfzUu/lXEWYiyd
SatuNm0n0rdT2jqMi2lP4Jg5IUhHBNb2ndFgt92mHRV6DRAnbALRFRSSdtwLitYF
CeuH/ZuQ+4mA8VSySffsnWuHvGcG3fG3njSC6I+eSsJh3mrVVzUBpjjQSA5HaJn3
9YCfaARQwlcb8IcKHx1j8iH9+KPblNwhZVaw1Qs085i2SRMWuzpVkIx47zBFzOZa
rlUGtop5AMbTTyHTJuPT7anSlVG5bp3pXofE0M3jMoxCa3f8ROo/2621aeJytaBP
jWg4C1QTbYbmuu9FGCeB55VVA+Xc1fMyKbU38aSonYzAtb8W3Q3FiTVtOK5Mprpy
D4KiMzwmlkddDXsu39oE/zdIE981ajVqn2wep1TwTjxO91l3LPtT+kxHs4OwjxcH
j3AAXeTwYE4TVgtyRjNe8W2ScpZ+5h4y69lWHtJdwsHsf2pSRS1pdcqtrBz/wvg9
wR4bUdnnydJelr30c4SJZ3EGX6g76zoTRwD7aRsbXy9nebuIULBzZU5uE6dFh5fx
0Qq6J/I8KTYJdOsmb+MrZVaH25/ROINDIN6K9O/yRtlxnP960RAWB09kGAAMyLvc
xcuEsntoVu9ttmAZX1YWDY5vkx1/pPJm5GBZwh+xgxrde73x0wmhHiSKOSTe9KYQ
q3aalvxaWSq+n6xr215zwVZEe/hiAZ9vR7OOnqKQ4+/wQIc2zuQ6agh3uLxtcU3J
hTRd0xphii5Wubj+o3xhuTejibtNNRgAUdmvfVoVO9Li/A1zVGXrB1wqQNJfloW5
Y+5P3q2Lat0A5UNOeflGQnRfcZd5L1z+/+/gfCQu42bX5yfTHCDnvexB1qlzXHhZ
sjh8KCY+ErDyxG0LDd0fhRqgysYrd0xdahIy5KET1GULpEg9uIa7PTUu6j3n2krq
0no3vOSL23vuY2tVpDMs4ByTAnJNbB3q0gFdlZ1/xVAlDgYnya8pQaXapmC98e2I
c0g+c7KObKKXMWc0YjqEp7PeSY6tfmjK60xJOyhsO3n+dYD6gMBHwh1OvVCCQTML
UAr/YDzEl1HamjEbTzQi3nUcEags4Q9tJRs/8t7k3PQsHST3mR3EEh2LfqRe3fsP
lc67PNDr/L0WfGy6U6+e5qOQ0ytFvRapYsKZR9S0xQ8d4itPH021zWIzEcc4fEk3
7F2ynVhKXmdNpz2ssH2PQ/CW/vfQt7bo1cgfLn89Q5RggTKJ5XsbTV8pSXy2quST
JHPM2ZV4is0/Uv2BErcKCvax7+pOd/urfBDi1ANZE3jbDo4jGWdCnry+SeUDGLcn
C9sQvKbncGMDxMdaPx4u7oTIeK4hDLXmN1AgXOIAUe4NsEu6sYVuIMzl5f8XWm+4
cWHgZAFdPOggfQT36zHkY2GZ5urtpTslpheFtZPlU0tDt1WgZM43oHvns7NWr+Km
eyULRdKKKy/9Gpxqr4QYFd1DnFWx3oa6XRiRRfabjov4HO1Un52vGT4FBmj0XbU0
P5tH1ItzVrN+p+CCDVRWSLc0j+FTMeo8S2Rav+nBrsnpabmaHi0W/jS9Ssup19yz
xy7ehz1Y2Yk3p55FUgEpruaN8HrUMEM3Fr6AdSemZZ6/qidjpzTO2ge3s05ap8q0
d83wDw2Nyr/LtMPsBt4ceoExCyXOE9sucB+2pGLiB9adRDseOyw0e1uLmbtmqXHT
iHLLy/4Y+rKCs6iv1gPOf+7GTFOdQUt6+yxD/+LKcnzvG2YwTuhi9TvsIWkupkD0
bdW4HpkTFruuaDN3hgOCufJK9azbVB7dX0RPgLG4bw76KAsz+uVlz0Q6VlT8+d55
zJLltDfEE6iBbJ1rrcllq+/QqqX37iHHLAj4MckBx6HtmBYBlyJQqPcO8lqSsZze
wCJjhO29+Z2s1YHFFHBuXFwuKhcevsGocgsm42D4TbvSU9EX4+dob2BgB0A/G4YU
fzvg8lQd+ytCsp+/1wUmxU6E5r/sOCVjnVhfqGZHPYMNBfXL9ae44zOfFUQn+lOx
TeflFBkIVFI0PgzpRRxH390Zdb75mNvb1przu838g8FrrWBVNQQ5mLgwAkY7lZw/
Epk9kfi8gKwvJv+OVSsI0T3sri+G1JS5hMj5u/I85erIEotp3QfvVi7KlE2to8UV
RPGFlYJ7VZc50ek+nAgbjiaQYDXQo+CfptGkoS79diaVHsGzVhETRN8bxp4CeGsb
aG2BvU84WBZkChppVFuoWwLIGZw/WPww3qXGQMRPgd3VBNoIHcf6QuG09d6MmeK3
aJg+USs+dKoUdsFq0GveHOejAEQv/v/zfg/u9WazWTl3NFHcZu4wWw86LJK3SS8U
Ihyem+auk9yULdKLdmU6P+I2+VT9N136HxTI8tYv1KOqUpUvb3XtrGBjQ8Pk4BxE
rru6xG3ohbQgcxgfiytz4L/2MkIC5UliE9niurM9Sj4nOFDLFnRqkFHmV+MZZJ48
PiPke+kdHeVilKh2qnQo9/KsVPzb+cm7s/jytoGPdjWvgly3pwhjIcI+jTaPbFiE
P+ZuoOKCq9cbel9lCvfw4KU8xXLoORrhdwQjJtg7F1/Boe8a06ej7wUhzLuwHLR/
tPk01utL7HNGrhunFYNr7uO1c40+7REwKLLwUB0cPxOPSzO//5ATOkTe1dEF3Qm3
Ocq6otxYmb+8i/+a7nRpgIL5/rVBlqNmh4/CBG91OAFe7ThbFwtHDzIxDoguCyMd
ELbtPvgN780yauW49QJjTVXxef4IVYajfvzLikQuxhtE7H0HGhqUvz6LQAvLkIU9
yAh+sy1nQloQZe5RjEdvFxzSjtJ0eo6p775z8ZDy2FZ5ZgSAn4mZBHMowWIrEQsi
R6GVSmwqeuLkC1XM5xOdxL3Hb9IT1CAJtHIPbt+Pxh+TAR+kPVXQRVKNWtawsFNT
IJUNw1PnZiecNdEynzMdgT0mDn8vlDjNifvdhdbkEBsIIqFGVxtX4pNQf0K8xiVt
StuxGkApcb8Fto7ZAiVuuCCSPAuzQpcbOF8wsWWgATCMVVUgnUCVYZAlzCBkoh9m
aUCtu95wvrdm+csQZHDGwOie0Cl+WWHP940piPWwYDDtBBLM0k9z4ZD0o4i/HWDk
fzgd6B+9w2EB1V6VpDRNwNPF3fnm6abWk8Ah2B+8xZvQni1pdKNiBhn/avLyDs6L
F3woKmSrIaPs1FdHJ9Qs8GAP9sjuYd+olcadmUyr4aGfUsMbqJA103xC2HHYMbCJ
pQVz0s0O+laQtu6rb7dL6d/nKarp1ukaL3mIZ3ymEXCJcCVg/LwhGoy7yWA8eXks
npwrJMEdHtFh9Pargu2GmECkmpQWtatiPYvRjweVwAY9PnGhI0P01iKPkoITJeFR
SGL566lsDME4+ZGvw2J+NWDEii39HcSZVNQvfC0KNzdrIZcTkC4C6/y2Z3MNWPae
AYvTd2/7aPAwqKzcqmKCCmodrUj/L505hC4bg/60d992RioWk3RJnLil+nd0rPfl
dhBb29txxi0nkjTOUqqGcx+xl3wZaBk4fjsQ+u4ysUHT/QtEa8Bzja6+NT0mHrO3
XGrQp0fa2ZKrHhz9bx1fjkuByootbKarya3evFkabaq/IuidfwBlLKPswSyhzmXO
RsQCf/+PeSNzjatSSGYdiNhvjP4fsIk51D9iUunbgWsW1ItBHtETp/9aeEhyhSrk
JGtG1eClUCOFOIz4a/px+mELPjPL0vKBO8XsQbQgZGdmDay9S8fMx/B70A6rv6FJ
7wCZKRDzmKwWFkZ+Xx5AD51HJ3RaLzB+2YzKKW+E5NDpaoxgxe1ZN5N54UDOcsTv
uR9ox6yRH+ar9NVfYTkYG19CSrlj3FQPLAyEEfIT2tflZazn4vFDmFjVWHyK8/Y7
KQs0U7inTSnbFjbF1B71/Zw6kh1aERtLDOTP885zCKut6bIU497r3ewzTwbdE9L9
lTPKXl/jqe/3WLDzA1PKrTAYCrK839l9ca4jcNoU7sb4hy8F+ZvYGbAQ3w4MZz4s
nmc/bYm2oF8O5LdfomBC6XiTVKpE1uMvogsja1s4+pHDAgy+quOS3xYYkSgWBR6y
K2gTSq6N450l5KIZpZNozmncaqXEoADJ4/pyXotN6W8q8AKmChV7TqiqWMe6j0lv
IqggporuGchs5dTl3B0TayldjmFqSQQjjNt6xUfQuzLvlBzHe0uzVCacSTDNrema
4hTDzTnq9PVoFVc3EViEBQF+G7NVqCrJzLJsO56TvyggBYD2x6I0f0Y0yEp0hf+4
J2kXX383GaPKornZMWnoJKhNhgekOCm6iv0dGmbAnCX/zIy13+CxUP4yLHGHDi/x
FREwd1yxyZeqkmZZ1J6j5JopwiP4L+nr019PRz6v0vsz8Rsv+xygLSK6OSsEqxXl
bmwjbc2oCQq9TxS3g+kgdc471XCPn7AHUrGXRMaYND3tilfCAN5LRtEUVF14FvIN
SUASIWl+SHqDeTFmlntZYsshf4nYxks1OvAbsDF8JPHcBZBUOhShft/f+naw2HA6
rEmYvVFSMaDuj/irn7EvpWI5vihNRxADKEjiYlzWnjq7XK7RXzLF0XhxdcX9RpWx
rENsgJHW/JAOrl/z3/DuiwTbnWflmn1aVb/gxgI6Gpfs8GwN+I5bBGzKOwZp75Mq
loZ3svExIPhX94JvEWiRD3ghPdoKBQlyyMYovIE09fqKnk46myX4iSWitnJA6Uci
7DMwWXqDVqjMj+n3wFRzjzqcvm2M6Jxe3RLlab1UYToTseFEOvU1egIEjPuepYjE
OlYPDKgv4BJVOzlzOoiOJDA2JaxtKSMaRdkwJyEUV+RvFd0ws7zvdhmgeLiEA/Fm
ZF2tixAcRlbVCj3xvZrKKDc164B4MFEAtHYXEKkn0a8oDuf7olNRAiQ53KiivPVd
6j+E5GgBnlmy0YyRPtuj3NUw/SaU7oNI0s8p9+bpoLxY34fzEE5b5MzKxY1nYYS+
2tB+5gIH+nMMsnh+YXjVmmHQNqMjS7FvnlM9kslmrI07yIlQ6vmx/r+qfmFIQcdh
d6cyJewGP7P3Hl1HpHe0jip6ZOS62JRZrZ252RWlLLUo6HbsvRm1b50VaR953axp
wkGT1ewfOSUeBwoBhH86qKPiI/lBLEWi1/pEKGjvQrqzcVjJoAF/f+bCZJ3nHh99
kEb7zn0PoBhc5FOG9YAE4IhTFMblLUvhINfu2Pr+0LxN5lGeWkJeZHS6SqxHnzsq
so71iWWtIbsmQftym6iiUngCcBYQypK0iSyCbSpvLPjGuGESqta8wDk9NB0lUr7V
xQ4/bpcPh3w3SmWQlYLvlTHvzbsooiAq6SsgM0SEDDr0ss0gA0A1RHIVCrgTPAd3
wMJjpPNe7nmMGYqh7+tkpaeO59jDDexg44qVSazzSo5LJewd9sAcYgogpl9guUGi
TZVsq7w1pf3wbkADSJiNMBfAkFQcpCNvrSAixxaENI24TxE6SSAYqV7N0FfdyC+T
Ov6VYYA8TEWTUAMIEK3pkEa3Tv1VT01R45A2WUUmNlYudkURjDg7j1vdPee/3txe
Vty5vXmwM6PmUc24odt4veo1981/607Zm7awlPeojO0z8F/CUGN9LWsM1RW651lw
oOktTsqg7gbfY17oxjEGXHsEdAiJi7AhY0WzMrzgxAM69XNeSPzKOFVCdRxuIc7B
7CS1hQLNzAL5G+0WdnVsEXTfId8od4vUiJdZs9bDQnq6tHxbnKskwEwINY/Orxdd
g50yBeRXDzVv/Ver+mntdxV3llLlWlOHDuFpz/lWyISVwZW4GR2qJxV7rha++BX8
8Y5yTrKIT5lSEN3POlBPfIX4X8Y/tZCODSW4WeEcd6tIodRGF6T11TejM5MJQh0/
gb80yg3z4t2U9JVxLedWpoY4pai1t3NX/D9FMJT8S/xIXhZj8yFPQ27N9ZHRYSnq
tW8rpGc2Ec+hanAshwOPjZXKjFS1P7rOkHNCjP1Paf9wVQU922bk0KtmiiElGery
A5/tvB60cWycZdWbzgwGthsHzLyR9Wu/WjuLVut0bkgNVRwjVasSiQid21LR8xLC
mXcrOg5gu3IemEkZ+4kB1yRGhkLVdo+RKDtuNEN781NuouO1DJI3ZtRMMYb9jB5C
pTuzWzhNBV4nliV6xzWqcHgpMMrLqzQrEc1UBgS3fXhI55/PcrN/JE7tlIoDEqG+
CgDSAj3lK1TwglyIzNMW3flqlIbsjyJt+jWmtjrm0RquHcOFR1d1fCDOWEglstII
BGJve874rEvzEesqhEvwtNeJxHP+pGRkPURMNCN29xcfK+LYsHc4i2m/JFT3Wi2b
dmSv31jZZ+iAU8VplM7cOK3HYqqRQ4G8nhgTfuL5f8zxxgPGMsJMMxwPHNafzP5R
e13PCvksdrnpVhLtNznjx70lp16KXZHejI8QtGETPt3r/NfcDd96jL2JxiMUxXNI
MRRyY6bYpd1LoPp/SUCMC14xJjqgajf8CGDXjo9tv7lidAIhFzr93jU+qIRmhvi/
+Oky7b3am//7bdKtMLxJuxEN2B5nxUsg4gpLIzEfUP6uvXXfJO0E0WaXUOaTapMH
4CkbVBifNMoLkLT88bCcec306l65nrpvWCNWhh7WzrzgJJBA+2YtKB0/TLwpQZrV
cgCDSb6EHeLasS9YcCl1gukcpoA6AcjOf6eAGfgHCSVNq1T4IC/SA2Vn93Rnu/yc
peZ15LTbIvZ0TsvI+u5ATbFLHncAOdK3wX1ijVz0oNH6zHax0LCGvbm898VRQrJz
kXpVL57D2fcU3GcvkcoeaIIte+3o2LxwjIsf1WySua/PXwS1UZvl8g+A42HKZ/Ax
0VcJ/0MtkVMvEpSy0IId6z0ib9/A9RrW/3lTJFd+sXGm5E6Xh3sIxjSvD0ByOFQ1
OOdTXlTA8sVebqMZN/9L1Glf0dktlqRWbK9FUHFAznWYIv/+Y1ddWRGSorQDHhX/
BAypE2AOLP1xsKgpvW3wumG+wI986o66ykyOwlqCcfe0QSevgd15lqUmuHuiTfyS
5BLohRgTvXHT3wj9lf71b2hdaw4XZH+aa46y016UnmjjnFeC94jpXdB0bBV3pLax
NHFKd+n3IeEz63NHQgtIOcisBUwQtwuppAqvanviFkDbYfYnN9VyQfYYJ0lyUrZE
Kqwn65aw8wyOsZA2LLBR2YAotoOzsRSXeTW9WW1mhmDnnjxo28CCtpu1glzuEqDx
kgsEGMD3W0BcOvFAGVW59t48x3yuHEH51s2SavKdizk9rcLOcWkrbB8iJ2qYUa1S
GCUkgDspzifSpSAKTymAbPZUa0o9ePZ8mXWS7g8EFGoEL+IufEhLbXCJD4OtlOxc
Fqqqjw4pEF8D+X/Nm6lK7Lq8dBMwCpBG1YqXHRLTMYvCms9ESo7FQB9D55NR/uuy
T29pwbTdq1ErGorL7IQLEdHoYZvM5jeYZfSHDPg4DqhAZUQYxzZL4K91VQPsd1Vj
K6VqR3hkuT+1qSAFiXTCFuotk7AKZmFATX71M/E4/oKqAoy7BAjjXu7eox05vTur
MwYJglq5kI2r/bagojYaaxHe09UVaefgzayGrmex1f2gn6HoL8QODNAuPyxe7fnh
0Z4HgJxd5nThMSsrvcMboNM0BHzuwh9PCOkiVIn0se0XvJFwDwI8OCyK87Q4ErVU
9rzy7kMVtXNoH8/l6+MC65pbPxDzxGw+O4PYjc4477xQAkVl1fZceyAGMuGnnbEV
tKmc400IT/mw7doalmpuyMlCtABU7rXPCoua1mJnhM4H60ellAMY0ihMtpeZJPQ4
XGlK3tlFqnDkuIV5HI7p+TfKBbpMS4JOzx4oDyMTHxLI07FaT6iGjA6lz2AeJy0M
0RjxD86zijXJrMoC+u9peX/LjIM0HFjmInnYroj1NFi/gxhs/3BwjpJTNGVmhiQz
eAHfFMY6LaU7Jci0ld1VWQqMNiLQvsu7Ng2aE4g5wvAwcu1o6wr5xxq3Bylr1vzt
urNuh/aFDKTgk+akOO8/D6/+MYK229Y2HpJJRiQThdpODIfNFD0TD9KzyD/tKk/q
H84ZPeP4uA522zpUSGovTrY5LPVP0kXVlR1boYba3c8Pddkobkz9/ioyVD9EYQNO
Z5kEeFuU0HQy06grV46f1rQzhuk2tu+pE7Kel7F5NjmBi8HutWxp6vZodqCt0Zxn
4xwxl+NvaygMvhTi3Zx8Obnj497qR6XsvgCLXj+iqDQ+B7+w6n4uSxKFzV0fzZbp
BP+SC66aR6lQ+rx2xeoCzFnfoZ+z1aeibW49jv+heuVfOxg4cCUJ1qG4CKFQghaz
fVhyyg+WmxFsKOJhUSCS2xEGhwDBTbVtnEYQeIPMtkB96fUQHZxdExltOsUI/o6F
83o3Pg4wy+gYDqCzmzKy+KpAeTubWrg0VlewauW/sZk4v4pFKh5nmNW5wqfpL9lu
ftpr/DFvz7+i9BOzbt1xwnGrGNN1hkWIaX9+/ESAxT13066DcFWFEoEyNN25r3J2
8Kw1EXGbrStdm/mlM7dK+pvUDSQaHHpZldX9avADx/5Q3yz7tH1xTuEyvvvLsTcc
zS9sTcHs3TrdNXbQxH07x/Rc+A1CsuHLBrq5bxxaxMx3ISErYX6JStrzvacL6fQF
yRhif7DUwm4Rh3wywr/8z9Fk0t4be0dWbmyxFo2ehJTDo4WB2dcyo4K3HQ4ipqtp
C5u2qeducbivnaYSv+Ox/DIK53npa3LrIOsQaq65lioUk9LWjkOUZqQu2bqeM9lK
EWU5ps7ihqRfX5VXCYmPEGEQkeudKkGSxbKTlTMYY9BtsFd0unIUpoL6vcL//uWu
8swVgWmr9LdSMcuFYMg9mKygG0F/yLNgSvVmlXwXlHnMLo5uv8YGCsaoIYsanfdY
WwGRZzLDmu+RABhhF7s6QfoumDquoKJbyKsNJsFAt/MeF+BmYlRglz5GpWHjjdml
LDISl0YfZGUmHu2+DagzA/sg08/Rvh0r6NZLA5WAi3wc/qWcLYRzmJrmzKw6V6pd
28cMcbfTBJrlfbe6kDpMIbBmMB8Mdkx1CYJBQOorWHbvt6u3+SGI8bqhGAtLW1qQ
Kt5uf6Q+VBTag6cDvVkoymB21GKs3V89BmSgNFwmHyKYotEWtDQiisaUkc/8rFDU
7UfnxRxVfIK+zkXw4y1O8oE19qcWscK2+ogd0imZZAL9560sSKF9XpR0K6CbUyax
y0eDcA+7B1qmuolOZ9uM0NHsaOyLJTWbWPXNWStaNqNGFFMf50DhpDomg4WQssPI
Y21ShbtEVtgOuyASHOclfaO5i/EfPDAzRcr02pahKKwEalWnVX5bBXEdQEtFiMdB
5JEdeJrJFRKG5tM+3khm/1xlRlFGmjDYfp+wQo3GrKp3fSdag9NglSgJujEgV/26
56rhifjjxivAAHJSUPP/6iKjIydiVgKlK3vJ9mLKzo6F3C9WbhcJMiwplDXD6LOK
XJqz0dn5IFaLxH424T1M0nN6jJH1HCbpwQAPgxhKfHh4FuOM6/3iuON2Z8udSdyF
o6tmCfZEXxvFKn4ZzXrU+7kgTsf+ky8SpEoEa6NqHQotsvXxX3+taLNf0JY25k+s
bzFsA6heZUcxgyyJoKfNgtJjzNrGyi+D0YaCN8sLDPOC2w5IlWMgn2SjWBEHvyaq
Tpb9GFj0v43PwWnf33PG+THG+voxQQnvbi+x87ZEzf299RXXeQFTaY8tziCHhClX
euvF07WIM4hoAAc8VRxSqLuEEgPce+3G+SuQNMYsxXcnypPFVHRbcZe43HCtTT6u
xl2q8zPZuRhe31KSZUcujb1Nyp6dJLiZr9Zi/DT816T5RAjOxs1rmaVw2KpjQMS2
158JPztOOPN9XmriW9bP3CxCOAb21eGXSSDu/Wy55AOPSbwO8JFgnvwkxFoMRF5s
tEnYF1ddf6+Qnfbw2GLzdExilVEwQJUoXLETtJ4UsfHfEYE5BUDVD9sAkot4vn4H
11Y+YZwEUx/rL6YkHxJ/aSEMrfTo50Exl/VOYc7hyWJo6TqlpR3Z77blDfYIZ+UZ
JCJqpCPAiPzxTtL5NBoSJveOwHAy6Bjc7hkmAvQOe9clWaD0ValPGbt9NZwYK70Q
DX8u25uDNBJrxPGyFFTNmulyPD7/t9hj0gOIkY4CuTxMbBaJP4LEqe1ts7U4Vezo
LhQRFcCUBGN9QpWIoLsgCw9gnuLeTRsgOZTCXnu5sZm0bCfJjwzJt0LTjb25KJ51
S0CGTNGCkj/XE95ETeFGByt3Ir/7jITo736ZePED/HmoKzHuv9dDEohmxUks1aor
K1nZaMY5SbkboRVtQrwJzjBJC8Yi3As7ypw4wezWj5AoMbkgDWq6QhHzabVQqEXI
rOaL9E4ZdibpcOGPJ0g8Ah70TKTNBrEE/Nyfidkg631ZRZogCCDAZtmV974v+pah
uEaOsBqmWoUoMt915IrtLMGHNTrmetL8EygiLvrbD/UmRsVh4KWH9w/5ds52xPmN
ng/IQ+EQsOwSMV4rsgZyG3DB+0yqFt44L0sL1fAZGMz2WnmvZnbNafT/IhK8LPaw
HOkq/aWaw00VrgeoP2PUcf8rLCqgxp+qauSCyj4v2Le2omYpWo3PO6Z6jhXkw6Vu
95Qa2oH7S5U3PHU96+RN9WWg4F0eopUqNJIlQrN0g9hvYNRDjQpBfV9YXHZxHPXJ
WflNkB8wZkTAGMWNZFBaCP8p+G3UqSO7f9s0KO3YF/2wFu/tK1zDnGXyZTmZjovP
3BzM7YptfVHh+u1K334uSIdzpVpz4zcWOcPYIFFnGY3jAPQiUvAKqaTR0qEJf7k5
+pxEk7VVrdjkWv5WaX+1OqGKrzAF66jcFEPg8wk1dfA+VaDawh4BZpxGl5yd4Wer
Vf07jGKxv6/24rkhQ5dckqZNUCWukwK1wx7WOxEYcUoFUoLRJ2Q0sX6894Wd9Arz
lHlRlEJX/9vZWSNdpCatYVwKF+GrJiS7bm5FwvSAh6D43W4vaAAaRywEM5Gt9S9E
0rjIH7gBFOPLi9+/F1Oeg9sPRbLo65x0y1H8ZDDgaqk35799RG8wtk2dsSAbfHIm
FMmaw76VKJ5S58B2BqWt2pwn0WosSop2iZTv8MTxidm8uqcfBCTcOdVsgmWsvJNS
fnr4R7GGAkR/s5DUch2WGsj4RxbfdeJJ7n/BIeLeLqCFttAlw1uRnvgQbHiaVPBq
NEQ2OGDyniYRRkWjE+Mh6gWqBmTF8rDDLTCbOEz9PmSf2bNyCPmomO5Fu+2VuuAl
GSFVBvLs1aDvEvBkbBh7WZPb1bwaJqN/WAtCDsDKjwtfRxiH9nsZYZx+oukX3owW
JZ/60q2RxikHb/71TUTb++J/vemmQSDM1St9CboBz7zmyxRI+BujmWBquA1YsdS6
ReFM7y43V0L7GuEdLvRT64Es889NWOhUHdJkb5DKaalP4ybFupLwYqrekijngsz2
3wB7L68GDYrn1lKF2NpTWuAPpgF/kXfHtJjmeHpe5nuao0xxPBFnIq3iC11Nyc4p
fCmXQmESfYAJ/S9/eszgBfprfoZwJTLagfVrFVVhLj25v+RMbCoxVkr7gbF8FOAG
xSTSz+lO3z348o+AYE+ihZWknz4rocIhLyIV7Zed/f0Ke8FlNrrhvOXMYdJPAwNc
TPw8DJx0g1xIOJpeR0iuuYgDAYRmjWpaKk3YPhZXrfQFBZxxG/xwY4FIAQeOKOJA
k41NWzOiKzTkYm1Yj1sptYwuv4pfXL+arVk5NP2/kre7GuWIf/qavmconDRgyBMb
dJV/avb1+tWQ2QYlt1V4CawLZvoLlrvMmFU5qyb8t8qcKTkDgtc6P7jkw5RlTGGX
2fl+AzOOuhBMjl/7CzSG+cI18kqbmyzRGORgl+voUJ1nqPA6HdNPY/ZoABi1qYVN
U0ZobUT/xwBr4e4I+fg4c9Pxh67N59lb85i42wX1EmaQ9zXh9pp8kF4CzFQmRDNx
KynlqXrcwSxG+c5rVj34XDNPW7BKZ1qtTF12lz5q9hEML+hprCf25mAt2Mz6bLoq
maDLpqlYhk84mXn1FggkXGWVxNhC9k08p0hAr6P26VJT1/lBgb2kzgQmaM11SYhk
tv41hwygtCzx0T0bHgfrl/3k98BmB6UrNthhcCKfb2/lc2vPXxuVNagb+eTb0IKt
lqcen8Pad2/wPPQylv5DyZJkBDb2KPO+KlecCmLGTNvyqYB3pSSHeaOlA4KRCxR2
cYBH918jdFtPCHzdKjkzriT/h2I3Pb4h47K8WkhM0m14V0x3SdFXUSVoJniDfDT0
Q0wZ2+SnYKSZLtInF2XrwhiO2BQCZ1mAje0W8eyoDL4zBeFKHmQkKvXzcEtYwD7u
Du1sv0dVFKKyIBL0NATvHzN6ETe+rwWQIDQ37f8gNMKY3LCMycRbmPapzAHiqQyS
LPasQGe1y+tmEDNsI0QCxjLU4Zf6mFE9S9eYP1fhTchyJISkaM+Na3t6ZDlbgHGC
OirAdGh9MZ/14zeWDYUJai0UXnQxjV1GDL1uXe4MM/nCVNyD8YJAAygDa01iSAIq
TnB+Ezu1+8CsvJfkJKuEQzgfSmzRw4v4cm1YgiBQQMU3zAmj0Xc6fbcYHFaZaJFr
SIhJPuGo38kMtdNivzuWt1xqSBxaaZPsiR7WGadFTIRUaWdJ5AxdwhPgr1uDdMOq
TR7lf3rAV19E/QSL3wZXegb7EvYnUFpC/42J7dCkQjGRj7AIOxxCFMf5r/XLJuz+
8wMNmgabpvMjGQBmSr3PaxfPiaDPh3PGL/WIq4AzvLK5yxl2Jg9V9vMo0CtIayVw
ohvsD6sV6/VYMywQPqv5h9bBvlXsVXIP5wPeYOcA07n9/Cg2ieCxRyQylo6ha392
hZOR47jrPyyPydi/rYWq/h0FVWxFujJfDoVKU0X2zW8u0+XCBlS3HsmiGJkYW/ay
Hz4q+54nL8EdAZAy49i4lWa9D7BBVMuVM0P+Yimri77V+B6cBJpM3XkR3TIE0r2/
/M4M2SacFGpgGoGlig62x87pnxCc0mRlOwgG7U702a9Nj8SwepMu3onjUpoMr6IU
4rLW8ODa61h2PVxRiPLQX0sO5XHtUd0Q5grQaYNSO6oNfJXRuZESug+8ykAlY6+q
LhtGhuwWdV6sUEvSUJ/XaGdozhG5Rs2+bfsage2OlzfbgFRKOC1adDcpvBQjDeUb
rncICPrsvI2PZep/bwAD96BT5qFVsfY9UVrlbl+9ovqUAdqtQ2i5/qr89f5TSSrD
OpdmFuVwrt/GkX9T6xta4octPMFxZuQK37S8AcaX9wXZVw4v1JsA1PE7ArgCUzIn
yMVvhaXYBIXY+4h/JFpLeyIpKb2tJCT8QVrT4iIZ5QVXWMH3qPz2AA6lxAH0mkJx
y7q8P8hmVf859QYxsTduRE3z9AOS1fLJPnSOu03Si2qN9sR/v7Jeddyd3M4OHjNj
F9Ad1P+hrMOqpA6kChgtvR3uDxqvvW+NaO96p0hIE5P5UeeuDDMZvm9yygcORZVz
T1ER2qGH3INglOrN9RQMfsrd6L8EsqjFBQO/whLVNOauwVX6kXVgVvZ+TXEsYMuO
ZCCOAUBinujGx3ne6KoPSZFRlQbf9QmcHU3HrE/SZiOTOPrybjfBrnZ941zw6uUO
6vWJ+3R6V3fRz9g81gZbb5jyy/O/4vyxO3fI2eaW9Gunhk3PGH7cVxPlcOkJkL71
c5VbiJLsqOHUdPXjtklTea7ng2zO2cL7ENOooqBCdrRJ1f96Twu8eHIQla+gKA4Y
8LGKDuPyYuGI6zWFjXbPr8RCCW5ju8/HDCkibwUvvA7W3t4F+eNbHEjusp6f5H63
/qlYWQe5rh705Hwe9hlUFtLy1H74b5jXjWB9ZTOaczkZe29ftr+uOZrCpTJKUUJe
3sQ5oASkK1p56stNtKRzo4onF6vPnd1B3V2euI8JiGJA+8B8MiUkoOOw9fNV745B
jNPrSHrZ40TEBiw7ZYRpxbIkJqX8k3HEVm+wXBay6KoJZmNXZw4NPzUYlX5V4dKp
7Yy2AiEmIwVT2T0sSCbVhhU25STPf7gj+9KeRKsKNawSODttl8+UFBiCSCYQijay
X5eczPtNkGKOCqHlY7xm6zfPlY+TQxGZSxIXBvatz9Fj0COyPCFV/uqeL314izNx
1x77igCIlQE4BtEi7E+KQLi5LVPjbOj95O+agomcTYHw/63kbPKht0UW7AvUZfbd
nnLBYzQNZN6IKK28F4YT+ZPx8Zgp7tKXsqRBqvpKUDDQ3lULmhyWZyuN9ftqRj+4
w/koF01yMKsGWRkW8k7cnzHu8NAAx+zaD4/iRkSyi4xYEMeYuI/PuQVN+r+eQXZi
pgBXMdVGklTN5ssZ3C0dlqhwrPG8MGdwLUeH6c7vEepWTe/IrYaqozKq0asC6v7c
2J9tfJ+QNSCkbtSUuiiRvm8YtavVlecJ2X+tgzhOPEbyukmq1/n/KgBmZuE7Ei2d
L4OzsmyytC7arqUp7BQOIA1BAUtwpHHwGjlejOWln9s+ZQx4nffKwsD8fzAxm8T0
BOpZZp09msAX0Ay+NRVOumF3wtE1AYKpqE5hmxs1rFYI5q0wR/rmoLNi2O11VdOk
u5xB2zyt0joZ12g+loNZRyrN1ksnIdlB71ExVu8b8RnfJBuAZTgn7s5C7UIrgnJH
uqajI/zBVQ18zLVsXDsZpTsfXA6uurI9j0yjIHAyRZaR4+Ccmv7+Cy1DfRVcksal
0c5gJTC6+6MkOpujNqBEzXDPgalsLr7vSBRykIsOO7dRpVTiAewhLhXjSblMC8QW
n3mca8TtwRObOfJ93giH7ty33uJL4frFe7Qt/Ahe+5zv1p/VvWS4oDYZSmBUkaIb
KUKg3zAjCNaW9PAWANWxKdyaqZy1C2sqn6skMvYsh2uaK1PB0Bx3jw5b65MywaV5
V0VNVDqNvTQVTQhX5z5M5MbzRmi0H8f3G4hTmqYUQfFuBSEHgkeAjY/XLM0f5n1M
5JTd4NP9VRPvaNVJRR12/KeqDZA39CJs2QxT6oZxHFsjOwQ6QDKDATQhHG1nRC+x
9PmaxA7khSeS6AAzURyq8Dzw5+49fvNxDhIw1/PxtoT0RC0hyQYJ8xmzaqa/PqzO
JPaMor5CaCk4srG3/dOer8iQXc8uNtOnH7QfJiCmTxHwZxjlQ3mCdDDKnla/rlos
TrHZJ4KEGEgoQVqJ3ckazBkuqWIW51sVpS75hHR3w5hjPfJ/SO136OhLiHaOORGV
fxhYWS+ib6MiEjXf1q0JGyb1y+cEfVCz7QtkDmKKL2lNLUBLwRQEYmuK4nAcoF2R
77ReLc430HFrLz2EF/l3gNSGZ4tgOshgbdTuuH9AE0vhMFjj4nDpx+YVqE7OJ3oL
xiJMFMgaM9F4PDuw71M9LpNYvwEW9aK9kUa9YP5GXJ4DAihu2H2kN1bSZHDxGrJ1
vrPqHpbnme1fR/SuCD75j+wCaDqS0JshVKc6mhIRvQQfMB9UE6tLt2YijoQuZ/QH
6YG5BAAmZoLXchAeNeZOrKn/Gkqk6gzvAolbfDXl+5oZ3+I0XLYG4IOBA6yvPH0S
2EfBwhVwvIMPRr+Zg8MNeGoO66daP81Y+SpE6IF2ur7wgJqMMITFrPyXbm1tLnxF
I+bUZm6nPPa5U8F5KR0s/UOnC/pPUDE+4kJEzxjiT5fG2zT6wE8z8IsnpltBcLR2
mZCM6zdowqlawmKPL3LK3MFrRabsfTIOyyEmluJzWPqfMQp1r+n5RnYpmb0B4Eb1
gRLEpoDPxf2fpqRFrKsYTEEiwlWpsZG3eMPv8sSKOAVaskSPvLMDsWOQgW5+PmE2
zJMm+rVYVP6ey0rX+FOpKFYdx683A60LVzgAAfqBHIB0IOHJNsRTLKsFwDumWxq0
BzdAs3BVoJwrUgPmLR02xXC/RAcFkGtNiuyYwSm5SQlf8pzPA+eiMSHSWv630nlt
tYyUuaShRVom56w5ZqSESugz1+TM6SPMxWzNwBqyGL+dGQd8uAynfL/IqhUJneoV
zgKsMZ4RZZgRmXkm0hwWKtsyl+1Hpw9KAQ1JsdM1QofcTMf3U8PmU6Ow3vgWbc2i
2xucxVrzQw9TnYJbQQshjTEHCGH134rPQf8LxN4m76zEkmVo9CGY1EigHKkKpu+I
9GXvYKu6koUN7F/zKWyINSJNQryX2xa4wBcOGhriP+LoJ4ewoCabAPj3q3NsIDO1
Z6pFeYcbrh3CSxTIWcppusUe8LjFQQwBvfbme2W0MINkiiKwUIBG2rIR5VmM5pEr
VXCOOYe4N7n/PnGHkTiW9ZDsqgkkY9Dzc5SImJJ3civ9IWPsRVFaZtOj4wD+34lD
cHFfkk+dv96trzRnICGUDDzldZ2dAnwldkiPU/cHr+g1y31qqjMYb7NhHlWRLexR
jzabjIsOzL+IMZo9xVZ+xKMMFAQP9PK2DZZ8KqKqjTTVK6r+DSkspOnxNAeHl791
oL7hbfaRHASh1M3kMO3J6Gxwr1jAqUVl/Att50aBOPMFEbUAF1+onFT5ZyDawMQw
3Wm4KpKRjTOSDktK9BYY1sEThv/BYRxq29xXtSMkARLBUhXcA6TkiyeXrHJguJEp
Y8YpHw6n7LlrkF92hmvoGMryAoAh+6uG9SSVRTUteiIrGvXz3+Xz6Vb/wOqIHQS+
V8QDTOPhM5I/VVWMbw9bUvXGT2z/UKbS+UcOL7onEChBm/JMGO0/YC4dciVT3kfI
ojXwQWq2BkVxzCSPcuEX8vuGKVZ+0mlKWDhqjUusq6G1xZeL8r/35WxJXlfQsTaj
RB5nfPKq2BPBS93bwCjxbJUAVF16gYcgWM/aEo8cQ3z9le6dWI3MdzVChij6pHC6
MsN6je0zS7xnzJv5nByzjYueHWYkpBU8YOPZYdVC3s4xGJ1JU/sEUD+1BKMrps1v
tS2IwB1cJonW29VTmlX2IpGG8o6JHeU3qtAG33V1hCdNP/UTbd35BHTk/gqAjK1q
W3y904p376yhuhV9AKKJl5Qr4t20HTFR1j+ny06UhK71OvBp1U9rFtgPrxEbYXPZ
+5I7rI35n1YGngYPIjuZV+Nu5NA0UXLkw0T/IzvY2rA0Ikh4y00hh1C6GcrslILU
od0tgduNRjyaQu1KjUOktqY2fFlPKsICXV0253k0CQC0TFErQB9FHAMKWWEAniKU
Vw2tqj7AbYQirYSthpsOhAk4Xe/J29cdt71An9XexEsOZkhlyOTHEhURKlXWSGY6
R6lWu/Nhrk/vvngYNfI/x0NlFedoZGHx8tNvIBskw+c2bRKZNgbUR7+iS+apXcYc
3YWkU4ceVQH0TyB060WfRtClwswibVUL4CG0NAAmEflrRLKOBu3VYwLeG8ovE5Lq
zJDMvQVWYhVKB9f2gsCQhNX4sXgUERyg4aL0g0pW13JvhJ0AGhPkJhwNhubqbrir
awB0RV8VH1NLeGMDcD6t2NprAbSYAR9kQpskOnx5SaUboioPqrcmjME6blxIXq3D
zCkc9vvpLgN89lvwNizmj0BAq5VGPsSBArrxheADVKmgj/EAXQeQwcUwW+z2K+Qc
Tzg5xyAmfy36DziND2p2OB1ptQDzFgOZrejgmffBhCTOr8K3GVdeERsoYFcBvc2S
bkoRjIzBqCZs0Y2vKOKSKbVLjEO97OkD9MnkJ9g0/FJSRid5JbhAJCiiodXchjO9
PppHYSphlwbBDPdEUC5ns6Jx+xsYFXxSip0lvXPhTzm40M9sDk1aghYftgUvsna3
HSBuSLy9udK6x2UPJf4jZaeO+BUzycO5upwb4QoVfmmj1ek7W6KudTDR7cuIBDAA
1cVexrR/M9uvd46AJlkwobjwR14q+iWonRN4xQUjuLh3+o6i49c6PnkeGOAUaFwB
ZC04FIqfkh+FVJfP+fTGrEId9V9EWsxQnilu/+SxDSq4ZQ98KW/1hk/qo0yledZ0
TWucegaBkm/ZpTXT7rhKC1jsooFBtmj2dP/JsxZ7Px6Cg4552pgCb9UeC8CRWlsV
lS1Ys/ql0pUVCKSAYiqNQ1BNsVGx8Y674r/VVUOSUdw8nECBiVij4S+VIt9NSZAw
vtUZwkiSOUOuCk2J8hSgFGOFfaz/2fsABWKoaLydlJ68+SFAvI3wIDvav+8ntML1
4jpJXigQD+OxAloDzeoC9fgOcXyKKYquDh9Ll29NVYxOiyYVU4IoBmbTUBeBzV7X
2jT4Jj5RTeCPxHbPCvp7HR2FwGM/P7MSlsU6jL7CEotzfzrXjslHMx/CHwpO/FmR
X9erdllJl/ZlEU/AhiMonBNiIOx/s+4njR2S/y7HnmUCxxEr2z/wY6Vy5z9CS6/D
SxL1PGWeSp03VqMo3nwKt+gVRs290GGhzN6375zhNwlmuo40o0g3AK74nn+1Ly7J
k/PxSj8aiQsR+401c0CzJKSRNHEIasPl950DQwwN9OBA0gWxY1fBHhmbpDYyYlZa
4LUAR2pybIwEuEovy/aKPMBwksJAgq9NvIQpOsnaZiucEchbTzziACkpsvmzGxdw
jsKBCNYxTHwarvQwDQEWfvx0hwj6vv/3/x4WbQbWT5GGzIKdL5j+FP1AQY2PMEEu
mt0xtgj2wQH4VsQRG7sITvfTR6KJ/dl9f98hgEhgReZt2P/MKXGEYVbw65QvofLV
ssOe7pF2LbQsfDy9/o83doWewh2F6yRc//0QdrF+6G3456YrFTPN4BcqA8hDxuJp
0n2cDQzQR81hlaWbFAE84kW3av3qYTqcyBU+HXrAwQy9kwbUO02uK0zkYD+ghHYl
9srt/7kiMf09lITHl9fsLyF83BcrsfUqV05L7PQ+KiJJ7VMTxcdOoMjn1o6gUxU7
sPn+mK/GQqI2PmKcGrPgU3kah83FtHBk4OWBPsh/8Y3Spfo0QaRAH9UsPxWzSEz6
UE07o7LA/MMJJD22XkX2JaWQaPheWqAt5O4T/tgR04uB/fGmO6EZ0uvv7uP4jxUX
uO/1Nma3T0AyzCgZPAP8QouGngC6cpICklwK+larxrJdyQSAk/odAqiYoxdaxSiC
KK94bVhAefxR3wWARVk+bnUjQc0UqE24NMMsGUmpvczHewJa5vxhBbxiS19AhCuD
I9wlgNzGVEj8Xq7qT1h1XBnYlv0Gt6I2RxVs2EwbQvxBMBi8Nn5GIk4grI8TolJB
evK2LAOPMvKzaNfPfbbk7bmfBl29ZDVmQD8XACXQBBZdZOXowEBmiWCdIOl8IBoy
elQbimN+Rmn+KbmlI1r3PaJq+xpRxpWHafkDVNkS3BHQ1LuAXwdr+avOIw4/8M/z
6As9gVqfUUDJ/VyXl3vaR2eqTpQ5DqTfQiFrD9sC5vqwq8PUHV0Vc5MDzrYWXSvr
EuaxXHtGQHAUpS0SMrc4JQ==
`pragma protect end_protected
