// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j9MO/AI5w823suYLMiVCx1XH6rvyDsF0AahTiwV4ZBGQwBes3I7w38K7Lj9k/DAm
BCaskJVSJEYZSwdMVmF4ymHmW1VMkrCt+n+kjlPP85fjZgj+oTulwf7n60zoobbe
etfiKNXbH7Bxe4iXYwPj4DNsMtb9Zc1Ady+jIJDbrXw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10416)
lh7NcPoj68kyfI7Xvn9848fhbE2eaDSeKYI3NKMuBMLlB6fgw5XzZ4BH8B7b6lLN
w9x7b3ESdwsCUKK6fZiqD0HmnEmFW742zOtkcVy9lgMJH6vJ4d+kXD7/XSaLFJXe
mmiOX8LhcdLUWCTHB0eRqrr6aL125+EKZm04PQan1Rmry0u905v/1mCdxymQ5Sby
lS3ktp81V2Rnz4biKk6jOBN5sB+XQ7D2TQrRH/ZXmKnXgdVca2ge+zrm3OxBxhm1
mYmZMAFL7ytNpCLFunmkF6r3UBe+HLe/U0oeck+IlYZ95oVEAjvwikr9NSuo9wT/
ig9VhGW4YdqFtHbRN3qA8AXB/l1soh9nzwTmP3QxJcNj1bQNaMjPfgAVJyAlGhwY
gEUlMiWNTyhmNHCCxV14VwzExvjBj82TVg7uwTuqCtGJfZmuVrpmH7cLxU4OYAvH
NNjFLoJ3JuHFKJXa0bKk6szRzeSWv7BFSyjJQmRivhL36SJ0nU1zpvokwTh825H5
G7nQ+ynrPlM16btFcXYou5sKVu84YdI4g3QSDfq1ngSa1buF1iYJvCF/hVkm6xsV
hbFrEd/UePfq1m7vGi+DZD3bXIUudD9baW/Fh0x+/x9kNNW93NXLaAp1989cTdBx
4twKyGokMfUHk+5kkjHxQMqHgVMbYPCyAidGo97UzrvkVN/GFpJLRcT8PgW7IwH5
jwuR4b6zd1obZBDzFlVPGFUFD62t5NJafPTb/cETtAUzMZxVk8d2MAV0TEj9ISps
JI4aXO7JEG38yTsSK2PHrLorLL0skHsT3nSjZupGMaLQA9+2igDBQPbKCds7FlH3
s/pKbnXR9CkucdAAEUfZi3xMm2WOngtIcghsM9YstCq24e7CzlNIwRulGGatEHFh
Di4UgVz4IpykZEEkP2803gAI6IVz731KVrVi8k/K843zHseazryQoR05LvlkMuS8
NY6PShubiWoaqh5j49xNJ+Y57jo4Y8HQkiACIRL8JZypYWjNuDiDEUa+BHUJwi2n
8vP2iQp+AD6JwE2I5qOv7TxOVmcyE1xSEqTXxjgdvSpYkPXTBGF43ykUPvw4BOs5
zUJRbvOEOB4t+FdWNj6m0EX22Wv25CBlQbWhOjC9za6anKD2ZUtqOx21pYj+iVP/
2g9o7QysL82lZ+gtnW0viQoZ0jmhNVASzth8DppGHxx9nolzR83RET9vY4lClQzs
Y1wTKSkJo3z7dBjJpyzR5asr2STh8AYFOYOynq/QO8sJbu0or8ryweSsuITIPaPL
4/Ub24s9IJ9i/r9tOdeGYQ9VTglxPtvUOQsHvSPLBrYnadAraWd+dOyammC2y8nl
3OHsj5webeSm1BUZILLfW4aa1MLOqZ6asj1YNul9bXr8dGZl2fDuCQ8zae97JHsS
O2qsfnV0VncmD39CaWTX0UmXi6581bR6hnmxyoL6m/V2BLgu4pmuvgrcugXJgrcW
TV94daSXUFJ4ZBHPceo3fXcL79jvH+tuUeCzdVcrrxLOx9ZUSy5rH+Oi6kRODwX7
WxFDN0KdRSyKatWz5cMrKjh9UVM2QejPVngcOtk0WrsTPAcj9hyGYadcAXWAiKCQ
fc34lgxi8yC0t5EJTKuZFCnWwnWbPuPAEv7X+3txuFgpON70QEUHAluRJqFwb7sY
cMFrjkPIZd5ARzopBP2qNMD0Ke2JZQiIBxQiFjlf9pcvxaTWuF5cwcO60cosmuoX
dLvZxepIX8KCU7i2xsaTfBQ4Sqsf8FmV9akdetTXXdXb9QycUoAQpkuIGwljOIO9
1zyuDrVZLCx+fJ7z++GxmOQSGChuji8JCv+GtQxflF1vD4FNQJCMCuvFfxQcNQTs
C/lA8503ZFVfwphJefrZpv96iAuhIP+GaPe052oSdTKEYZhPtUQAG6fc2MzhK/w/
TsH8NaaP/Hfh4WpmsVz3JfPzZSl2c5+45+TpgTizjcj290QR/EOyDyHfjenxUaNr
Frg75uSanNbQfWe8ElmT62q/e5BnrpeILIkv6NTEHN0ko/rQrw7cYt2VS3kQXnXU
qg0J4ctFhrdwSl8fFXd9ZhfRYvn964+0em4/3Mo9psMjXOsjuavd4yiwkDRzq+IY
zP7YOQh/04VKc6dLxx7yDoCn6Q93LjbQ4oWiMu4qe+qB3FVG/x3hE9ulp8iq0TuX
h1wF5n7OGIyMDxRJxXzJDXL/zcxWr71JQEiKSQtVzVJhxmYhBVGY0jYek5pc3S+/
BQdtD4wEpvSlIuVT0IYVUauKPc814OZnwBZIrNOsyx+6MZ9hCISebEgbaGasS6uu
FjKagwu92Nucwit7x06B+qcrH55q6XbFmXOXMyGPT4BXRSOviOmb7RAxpG89C+cq
dF/M4WheZM7/1VxA1K+f/8+3XvdHdT84ex1H9okDIOhzBE96q1UEbkzbdHpWZjKK
W9FbL79a+lJ/FR3HzAYe3gmZcpJv4JRS/ZywEryKxxh/JpZ6ttHArAWy2EZZEFYU
7Q6lqrk7BBdEjxFpNjOkqKHj5+0E7odZz0m7ErrDyG1d2qLeiRBP+8Qf+fF5FIGg
Uxdrd6GSeCVBabeiv15xh1kipYB/UsCVJcBo18OHEtlKcPjXl1oGemUgbaL0zPZv
uMJ2WRJxoqvgVwBkIKg50C27ff/WbbgRKtMi6TqZ+FjMjWUMOeMzuw18Ezwt/1Vk
O3DIgxAFbVNkoKcAiuiytVRat1O8tkiT3zCwBB3Qb3JqSwCfPU+73kiEul6+RY4c
72S1iwCBKfCQA69Ql3cyvReCqvEreUJzIxJaNMJ8o0JuLKmJXClmXCSEmn5nLSOR
/kGGircEsvna1NGjFBf8O1htMhSz+MD0/nPWIl1YCfhBfsb/c1lBQM5erh1nVFRW
khME1x1Bf5yWJRSNiyRfXW08EokhevzcvqrrdocWt/dSqqV0wEE6PjIBLpOWHorO
KzONFidoi4iZPayRdRUaexlIhfOBWaoAnHrBN0wbsLW/jm7xUMFfts/3gSVzLhs3
pltChLR8fKwYEVTKgD1pWVuZbKntA5Yz7fA3CxteaEX2ZcZpQRteIJur4X161u6W
Tki6+nvl05431B5D+sSc07XtOj1sFafQ10UM8PH8poyaI0A4ZR2SeVtvMZ5JP/hG
jGDO2lGAbnGgPvxK9OtHUWnqikCU8WTPXhTaj6rGlC3fhXaAeam6moBysLhdsKPF
9bSdjAGyEXdO++namaRltH7y0EZGb6iuZzCjrO9gsnmhiH+RmiKUDTpLuQpv7cG0
pxGU0kt+3zKtPuQuFuo0oFQilX4NuX7veiI8Ac/3J2o1PXImQ4XOkZDWnSGnnjKJ
6Fp5Oin+Pg0qCFILj40kD1oHJq0DdpcW0xJvGclGXt0Xf9ny2YJLltWTynxpyFos
W0YQ0t6QisAZBYOXUUVcOtXwMw0w7gue0IaFuD/O9Gv0jWsm8S1tXFoNZU+Xf0Sw
hL7UbPUlDPWAdZnHudNIpYk6GsX4lPg7na9GoCvDzEFaXafGC4WxZD31cnF0kiUH
dxXcBlVaB0F1d4lxDQtfaAW3a48fxYykbCDpH0xUY1PhGI9CgObt8SQKa4/Yv3t1
X4DquktNx5zAbw/kgo6UgqKKly+aXGq5Maua7+rgOeiH7NvZXM3RpNHvMqQdsQ41
F+ok5G/QvgDmAZ3JK0ODlYwjEuihvFADIGTVDRkrwU7M5WduqeOvG/Y/OWJ08LT1
MZ8BAdmN9JtDo6oSyF/EPhmVMpz9M7JZTuxGKDKEIx0Ec3SeejQ1FqWhTV5G2F+q
46muNRQwMMR0Wx2A6JZ6jEPCLzoVIiliY59BCR81/Kbj6lruKkfluDBRpky+SMcA
jsFoA+6H5IjVKvxSkfpe2FzVBNyV4IFWm2yCcsDyT5/f5CZfW9bv9LYqyEhZ33B0
iAxqO1NuRTCt/Db36QK97YY4YUpK/OfGJEL3QtxSIgvGLK5XN6UXE0igcqPt3mVa
FFJTYOALykpqv4Th95g1xjm6fUfH8ipvly1mVHOL1o1j2S3Sw4sSkgJTSd6pbY/y
/JT8aNazoV8d8dKFT1z2zN7nJrn8DuWqk9QiGrb01mNNgo2d9IhpvG+yjDJQa4G+
6Vz4042HDzpFQAJ0mvnPDvugh8OUfYhuqe7ZWcj49TCLA+ftOWP31glkRsRIUXh1
CaBW82GsDBd9MnrpuE+Fwf0lsHxYbcZLUzM18vW4C7LYnsfCX9gfPBB/qC64RHbo
KZzbKKhjDInm7ZOWLEez7uRFAqggOwXKkqPB8Ssbzd+CZ7ybNViuOYUfsC9xGVmr
Anzj7TMpckXgH/X2nf2D5IxB9P/V27detne2HCo4ExLxfeidTrUosXg0A7ydaP91
w4muwMe94QdBsOBYDJIg40Zq0Q91bZ7gfHwfxi3Wo+bysIFO3J3gsJqVCHqQoyDm
rphOSzN8i8S/kCLtBG0iTVfcgt1IQhD5TEXT3gRco2qCj1BmvEYl/UlUENvhK9rE
FI8tlDnP9/O28sEVkRhgQo/AVdL3kjxOCKISEGdnWLjq5r6MrKjrE1fBgpZ0IlWL
z8AyRH/m9huCfmpM8dRAXGXpswIiOg5KM4gBlvhfEAIL4SEHH8aLqgzgH3KeyCuN
JpZOhNF7Db0ShdbQVyzePM5EyNToZWvgdYVajZrQ9X4fe5ezBFlRgRY+1Ip1eRlK
m3/RnvJIhWZYuki9R8/JuQkdwwXBAc7ou59bjQRexNrsAnYZHqyp7xSP0B+gwvoi
G59HoxwbL+PTKZpj/PpEM759O2jn3+uq6Pt5Kb+wCOfnewvY0JNkoUoWU3V37BsD
oYv91WrbHXO/4svYsNyZKm1PebbVvFnSFjNBJyyPuXnRfa6BQm+CaQq3KU4nPH62
avReOnkHxORq4hKAFj5dhsYys5jaAIZN/Jt4GimeQQFBTmg84rgevjepQ65Pj2A4
ZG3uQm+vdhDmANkadxRlLL/qb8FBSHuUoD9cFSB9hYZ8riF0o5wzx6hbFwepDnze
iea+VBEsKL+lefrMzyU00dF0dCUc2GZtqliHnYmjBaXCXHf+eSCQ6xFOgHDkKSt7
YsIl+7JX1xykUeGtz8dfplpcdsBMtYQ7I1RPJG+DYOOCgHOh0zKs8zBSrQQaCfFk
BLt6qYXjpSWM6puKVvEcYLGnoGa4lex64n5387x5dYejFoquAh9E4SuVyPpyVZGT
tSWGyFiorbHkc23C+8Dz/pPiElJvxy5uyO/AlPT9tf00N+/pUfGlDS6Ktb6AI523
CZtkit3VEsWobcwUXtbhR7OvVq2FHpc4adONzwOMDHCwGxN0qxT1948gNbDdHXXs
SPLi/lQwqr//MBij2rlHokvaxv/kcEzB6ITSBnGapfVJIlFdErpiZFkm8DyRlypU
iLwoIRGoKMxTg67530/ALQ8jOz6ix9JQakH1asQR8wTl85CFiZv+fuKCJHOGM2Fx
MIVd4/0Qi0XcOsXPCXBI4cfZzs6YlMDUbnoHXz95J56yBDmTyBu4ZfLC1M5a2HA3
04sGRf62jG3USB5dGVljlOHcFesHWh76ARmBPOoA/0td13dFdfwlpnKklH3TW2Wg
+4CWoJvBMKd+peAgnnY7TwfbBW2/1RxMnNAqKrWMrD+ye6H2YAmmBig74V5JhfLg
gQd1sElJRveiXRBAToedNlze4BWpBCk8jvpo5eJvGYOPFlAJ0PbHyQ73P3tyo6dc
3G81+9lDS9sY/RMOoArXFBnphkg3y3w4amf6EEaYNYKGr5bcXFfBLR0haiHISMlI
EGTIR7fA9aPdf7pcKYrwGokU4hhl+DLLhAu/KNVvTut/KhWxQx12r1GuhC42J++l
6hxN4+J+3Y7xERjP2NZp1ak1HqHlxq+6h59b7UFM0UEolpf6OKIJSTmr/hveOQ4S
IY1kW03Z3WuDSbo88TfEczS8AGiEKX43n9pjyKuCK9pKF6+gzHCd1qdZwKpt5I+E
9rrbfPseoI2AIbzKu2xJlJeRE1G7Dnzgk8Kl7h546M+GzB+VXPDmWoO2pp81TFI8
sz6ie26IpiKP4xA9f0V1Ji1tRSsYypWEm6XgSzZZFgEI6XmIw34iSpb3ngvFh5Qb
+Bn0dvEfMw1vVU5J2tIfy2DE/fc/RnT6AU907fXLmeVWzbRbwacvIuasWsbJBbjw
pwV+fJfcymSiAH0H5RQ0BEK7eyY5rXehL36gW9W2peexRS4rz1Nt6bUxB/T0IH1n
nMm1FAERL9wdCg8Ri4kiuOkK7Tc1/AG6PGIJ0xyRY99l1/mNILOwe8c6j8TuCKUD
JXfiHKVMbKHd2I3IET3diPrTYNu1zoTOfJ7+ZUigPziB/fioAEt68BcAn3Bvu8Dr
pQ36EPaoVhYon4P8FBYfXr+mO2YxLSX2c76hPaml4AX37nbIZTbmXP4QDYvNEajw
/AeschaAItQHSJMmNrCB1knBfo7Tgox5Qc/HBMXPYtgSVQ8byhTTmkn9i9Y8g1vv
7idDPfctqK85hsoMO7uasqnkAwAOFlZiaHxXSbzUETP3zILrZ+go1lB54m8gbAfk
3Uz9oh4uEQau8oL2cOZiS7XHJ8iIpIUQ1qVPI/ZaVa8VdtdPFPTUvL4CASRL51PO
WIiIuvLPYYWaQDzNL5z4ggCJpN0QuRJmClA2RMQNWqIM+rK7sT+bttMMAkbvg2b2
GOvdzc8jLKWwsOGoYH+5IJHYQ5RuNQ6CmXGK6ElNBDhbyFJXxF1v53IUlbFQ+Kfg
nRBrT/9K5dD2Y+TRsc6m6xdaRsZE+FYjdFLFNbbZ5Ic1oRSUIPh1N2+Bm/O5PH1W
G7nX9Ue+jkLv+E5+MjHPDWHnREyt9hQ911QAwGz81Cu/o3d2E7I8hprY7CNyKlnQ
kAbpkuD3FOzOGKz/x6ZrxYfafumM2GsLhNTr0LssKAJaKCB7qYtgpaYDZcjBo65d
YrSfm7JjKEPfsOt7zy9F6MoPuQLx4vAnXoGC5RlnpqJkmIIz6ye8TZgGmXcGI9yH
tBlhF1kQ9v//0aPO7sKt0fz7WAN7zOaXeDQHaftBtxDXzgD979+cwysa6KBB0JgY
mdSvUqjqQTsAYmbFng78t4injbZtXeZJsSjfU0b0tQXqCnU0hwwfB73m1glbxS/6
1jnhf3bYB7T908Q2kg5vudg1zWtCLFfM5qllUDuXvHYrwbVtEm4nhtcZGMzhZrmp
80YrQSLGWFKovdWiXcVKZZl9q5zIUY1dsKS39E362AktdTA2+qs8Sx8Ad8BJ8Px+
F20gkWaSPS523+IuXs1UBr/ThSKFxFRclll/vKi6NuCssl+DwxoPL+dsQ1JBUUE3
5n3aN8R/zaX3hyf7qxitfqS++gDhnv8kjGb4N24GAMyity4ME3RQXQD6dAUJcbdV
xWuyBS4sTC98jFNdRZuIr9FCjtx2emjD7pfE/P8GIZLIRTvMdpjtMkAs/L6TywZm
W001XwOkYKvpYSCHQhQt49v+AvcfZAj+BllwIer3ube/PCnbc4eSlhSnRMRhI2e/
NEUpiQv3VUZdP7Bzt448EnHDZNQwf0ekjXS3f1mi5MzFPckxSMPZ0uhZ3K70vVtL
3t6a8CPnx+6YBlAoTYZA9V9SQ0NWAstdrRg7P1wrp5y6hRQB3gMVvgIZbA/ZSduP
NYJ6lictyKTBO7F9VHLKTyKcHnLNzlkyjyaADvKwHCBbxBqoBw5aUwlxQ66K85Lv
Of2sAmYc7QmmPJi5XCHLeV7F3ouRDMhkmu7YQIR8DWzlmV1GDSnIP2Cuc14gbdpS
BaeH6Ln3spZ/noeJ+OQL87f9UBywSOvpcw7T1G3lRvZkXxso1/ggBIyrUwB7SUvu
vB5Jho49ogfOpGujf5aX07iXIv/YkHL07GqjRumZJv9QI8E9Z/ifwG84Eec5TLvP
n8HncEu8r4mnVVh0C8t1Mq7KGMyZsiHPdbzzVxWQKGrUXGDT3334a0sFJUUBi380
FFGQJXTrnIbksEPbuZDz8jRgO5qxgOcvu39byzw6tFldLE1uhII4UJPuN1vhgBuh
+XK6wh5dl6EnCkowq/m7Q4sj9L/KRW2qiMwjL3NRxY8oA5OcV3kSFGdVQ2Zgl5d4
rALu6QGcytSg0yALZDE1qo8ocQ6Ksoi0IxrQfwbZE8JPuoG1DzFK8neb2Pd/Hes6
2hNvVGvNaL9CS679oP0+CXVX8tWUdx3NEYC6AraGk6J79azdwTMvKFKRpH+sWHH0
n1L4+QZKnSulKD/zc5eCMZSkYSbXokSUZILnZxkE64RkHz54JGWOkmxAg4E9MFQt
vpRS1u1af0Hd7pgBFAjswbgJMbIs0Laez3aHX3L8Jihyz1VQ7Yhov7yFLZOUeof+
0J48JNZG2bYu54PqhMaz21rwWSthqvxdQViT5+iU1g9P30AHi6KXIyUfOjr9UeLy
1dThIP9qk+9p/AhlC3DFteUqHUD9Hk4MiEdvukeaKFpifpvTMUBw1F4nv7BajE9l
TqRKWXl5A+/2MYI9vLURCKXV47J3YybRtkUZUZVR7giXaGbh/eWT4b8ZOO0VgYDO
gQJHnjrfqKlU0pRALX+RIo1MUD7XvEPj8Uk8olZ/LHuLuYnL522ksEmXDfCnhvFO
raMWNdw+snyMpxEdBGv32hmIcgL80fzbfw4QtQNMXGkP+aqR4HiNSzI1a39/HvXm
346vmcJHs60InphULEpCZ/MqlC1ooWnUpqoypcdZxZ7KUPv+nOMlcn+VdxW8MkJz
XCJ1G4Mx43j6OqOj0/+HEU9eSOjYlnvtLo6W4tpmCJm/vUYWsLNv6wjI03dPJ4us
LdwsVzVHPxOozNgzWmREh1HaXNTG8+KfQCpj547BKCXnMrEcjyRBj2TsdTxLIVwE
WX5BEQ6Pvckh1nmPUPym6g3YqrXIf4dLGsqrW6lECet5loJkr4NQdCeaqGemU8Dp
LT1vFhxhHEO7KK94LBZFvDUCrWRqAI6K5cvYPyauVh/a40/WFpDCyA25UiO1AuM6
AiQsnb3FsEcKW+zeO05UAd4U33KfK3N+kEDahpkQMowzU4VDmekgoDq6Pfi8kvLD
+FUQpNPoIwukACRVoNaUbQ7xwgkEk7/wDNul1VKrKD6CpN9eu2D6Ha9FNQtfHN0V
/z8RGPTC5e1MrCqZyOPEX1zsZOCkU+RYQxl+ClzI1c6rmucfi/QMrOo52umH9XEf
sVVHUcvSeaanx2lLRaAzBZHZrhQnG5qcgwGLKqXiBukPeWi/AoDgd51XiBiOolbP
iYYsReoC2v8KMZ7XEITSDDG2Pxx9fwZFBdC1Oy4CKNoVJAsNOmOmXnr9z0yBlQYb
7Ng+YGUqy5MOcI+UOY/RJMJXVH76+viWgYNpNCImAqaed9XfwUV/7iM/uRrNGUu+
Sy6giW79FyOqY/n6TTrVVrgPxeYXlK+P3XRvuN9JQ5I1j5WJB4vTv0qF5q084qR7
5hsncCCJmyKHzI4QtDW5Nba8G89rm9CuC9nhn97z25zG3FK5lT/noqg6LIno64Zk
tct0OjzjVXvetI9qeLByEPZstff8UXph7qJa8NGUAwfpJbe3D+E3oKxnUtLSF7Ao
eGMM0RgQBFLWoL1tvu62zUSYqi4FVLf5klYkDD+E9/P9haqrVd2bOGVCEEA8n67R
3ZVd3bcjR8fUAdrs4yNCRvNVXtzqIrBuYavJZt91vujT8SkELubpLN3UvbBSdKOF
UZbdpCrXMB9UVthERkrgcv1y6Phl1w6RLVPVZTuVm2HmdoE/y8xUm+0q2/FN45d0
Az2TNf783Bd42A3SwtENpeL9XL7DjU+AU84DZ7KmdA0T/UYOGreaoeccnD3yE7Qn
heBVr4JmlJ6XVBD86UW86FMtj8qCd8J8HP0Nr1zIVaV7ErhRnkvFBKVJqzwoQMQX
e0Lg/6vEEQGWM084kfAR0o/ciNswHH7REOWw73vKAP+tktmohRks74FbmC51SzVG
FaC/keIn1djrcI10hiQDhrcM3KXXoODSNuA4fBYtoU2ciojjTxe9rn3Lb0Vla1ob
sIBxBVedqV5YgkSrnBH1DS9xDIIwy53E9TTbDpuiy41Qq4PffTOSPE281Un+SYIa
yE/2qX2+M4JmJyoAKNOWZKa7eQL9IO0wTf+ffYDYmGpDlTuW1q7uoDyehEm37uAp
n12vK3Ky8EvjqWuxPrmdo1UQZTXErNdR+60vRcsvqNza740OGxBAG1Joj7g44pBR
jYoa9Gryx7LxP7gLc/ERvB4c87D4lDXHhjnI9L1vbtJ9OlME673s7MIn796J12Kd
CcuoDGrbdVtR/TJHjnrcKRD6xT9U5dmIjZUws5s5VPAEwBSjHI4TlyY87HUVagZX
BOLleIKyOalRKOI4r+qVmKliif/BbblRr7YewnTOmZ9j0UzF/J94gzwzqF6M6/mX
ta+9e4Cfm9vwnaBDI1cF2VZL5BYk/78e+GBOB2fcRDbNT3foCp1ibsPTJJyWKNHa
8mgYJms/1madyHy34hkknyrHEhYDO3fmf0TXsJ9wVY5RXs9oaFI7lhte4oSDqnEA
6twv5dsVcciVsJ2NCmtHaMHLNfQQ54CBo8cSYzAobU0GPQYCvHxzTKf2DNg8qG2n
476H7D8Dn3v9ClfpVHVqEWNmGjrctJfVYp+zITriKB1nNZF9k6uUaJVc8xrYu7Iy
7ZMlIRpyAMhPzcfK7Eb104OomFrXja6mM15qTelWI+FHt5YkO0lu9qtJo/SnkKDH
Niy5FpLtJyizy/+rIFrMLEgyZNjc79siWR8seyZWi/Hc6GWwcg71JVqQQj8zTcdU
X6EUnI7DmP0DBSkdTJya5YO+r0dZGdAEgmJ6TRwE/O/a0BWsQx18j2RqMxah2ICq
yDhgJBGS9M6F7ZTnm7S2Ud9TJyj3vBv1TbKbt+F9fQ+9zz/zxEpuUADGsphRQg9G
SqIVd+f6y6KW5cqAgBClq82zQJH+iHgU7Y3SnfQAVo0LZcwyzmWcu9UMjy1JzRtl
/rqISCB4KXhaYuJl/WFPaFPD+AxNl6s4cs2iv36Tuen7nXCyE3vdPXrHA26iwpPH
gmHb0d2kBWoOnd9do43kcGjJI+ggelndmKDpQjyD0X20ecZG1/k4z1yUC7BPQVe9
oRSykTwZojWfCDFYTaBMBWWNkmmkjtW6gCKGc62Vr9sblzJKTAgdzP68C9GSvdsK
4HdIRfw1B/CDTvOTEgcv6mOIUwlB6emdQVnABKBbd1olYOWCTaxm6lBiTY5CZScG
CgplbMgVIFx7WlXo6zE7zz+cSOniZ3LLpheY3VEEENs+zXfdrMaGjKPKi8nfBybO
N/uk+zLsqbyWzYxDDjmJg6uRJ52vXnZPLQK1m14atWWGOYgAHue8yxgOYOU7NAxm
c74nH1G0GeP/9pDDfVB8Bwn+RDQWyEcN/tOy5jiVCx/N3iV9Y612mM27NEM52GfR
Yw3lF0fjbPqOwSg9SVOAIXu0JuQO+XP2cXPCtRLE9ecfEsRE8Ab0aSHeQVVQCRe4
d3rpTZQTc0gq0xbJtvavjn5C4anS75izFcklTVEHKHwzEG1bIGvqXvEkn8dmjEJ3
I3btVAG2r+YVhH02Oceo9LK4a39lq+LjJlwH4b4rCUzeOcM+JqFri7fJ9ETp30tA
GD8QvzQv82761xDmOjg6ZDiXVREuxxG5pFLwL/aQ7jV2iy3zdZrb4VNSeLqfkMNZ
x00APbtcmUzXiZ8jINOO3H5Zf0dzE4m6HJvGaOJ48KFcXcgEG645XQVPYONK12J7
hzrtnNfpIREKid4IjJLb5mswOM+tClZnenrXucuPdD5XYfamRwj3Bv/1tyuUxEI8
KMIr6GJsFWFJpw5j9eXNIZWEym2c/Dt+wLk7/ZufeWgsS+7/YaN4K69peuM/iO+D
QDQz9jQvXLWeimlXpwXdoNqF3rq+xnl3WECOsH1TeHeda50b7GylnbB6PKDrh/i2
5p0r0wZSbvdk3MhecTkDgTAZp9XIzIKXJUNpK32gmr9XRFV58y4614fEhdrZ3D7L
fJub7+8356sVIoq0CjNJrJui5Nho0zK/UCFtalVia1x/syDb4jgdoacdbToYVKrw
ZU+Xsa6SspJ1Igx+kkVi0EvckS7HtSGZuKg1ICnsruxzNYvkHuPnNQf14CTJPlzx
gq/hqyz7wXnZ4rfxAddUMuIj0KfWZ3ZhnN9JE8nMBYCREW5qF+38ZpWaW265DTnZ
yrr1RIcO302M2tikeY9PoThQKdqFxY4ihL3/v5WqozSY/z1sFP2DsdwRRTAtQGRv
Lt4ZZlaZAQN9rOVlBxFKLKsHIIFrMICQC0S9JajLevY0kQTwy8n7vKGfEePbYoyc
N2AGSDug5gK8rI7myqlMq0ObO5pqq7vv1J4HKlZh1JymfaMWFGclfWfRSug0czWs
vRTso2ew/QbF9ECf+XayQ2z8Z3UI3JxnJeOq+cljEE5eWO1pgcaT5trZpgvaZwz2
5yPz4CshWno52yABIJWWe5um1TPJmUOodvT3zlPd+67ypAwy3qHGLXe4kNitvY9Y
tFQjvsuZJd/6fiffFIKRKWq813NmKTHoe8n9jvFLbV6adAK6Rts9TPvn2MEZ+vwk
Mz6qeTPYrbcBlysVSVbNdOJ5zmTSrrxbC2nhhsvvlClj7R1Llai51dKbpUfFJNkS
ECZ4fIe//sBoHzAQZZwdKGbnO5Za7P4tJDbO33ZNyIFukoc6sGKviBCxl1XaolDV
9fJ6Okq68D63Ee10PpfNKDE86J11eX0CUIF1mrB5Y2k7/O01qIR8nYp0yaRRqrZq
rwmFL6wTgcPH6YK37OLTZmRUIgb/MAu34FYcieUA1EyWji2qmP8vOLOHivOHU6TU
H5JLnNhY/c7R3V+zxtjbHGrMu7V0wkv2yTZQXsC2m5V3C3w7eTCOjF2XCArWMZFQ
9djv2WJSKEabP7lQ0DD+TK3hJgg3M0Vqu+3YG6H1Cb//PPhb+JNM7b78zN1RAUXg
E2un0nGSslT1jBUorhUak47rE5T1Jp6mdefNAI0y/JiymNAmz4IovY5RdjzUHvP6
oCqwN+H+VlLu38UIvmmPvyBE1XiKSlV5QFLLmLcU0cP0mHt4Hj2uKPbya9ZL8E8F
tb4i4mtkdiWmLKoFm8RPyiz6sd9yCFUhejihvlOKHLLXj56RNtJcldApnUs2ttQB
R2jBcyIhlz5K0DmNdfmdibX0cPHJQfecsMY/hM3CNpe6eTp33bhgOapS5q6+1Ksk
WsnBhHb1F1pAmpBagpIyvEVLrMrcpZ2/0rbA5lS6RbU6zkAV+x8u9Wjy0rwZKXGK
2q9/DVkv9haK6sErBOM0rtYNciDnVZPYj2bBgw0IHUR82/hL5sRH24bY7vJONCwx
sqSDpgqMqNB5DAQs1pkkpmFPiG8WqYouvydMdS+FyrfLLF9SCuiiWM2459CTopP8
63RqXLWO+QgZtOyZbPVZ5ZEqcIT0U6MaGbjISeGMihKbJioldCSJdxVyaW/HLjks
deaww/LXIl8PIlb4HYqNCzQ3J3mXP0ggeZJLLTWGdls1sGaHb3d7xJB6WskJdIFZ
eEwONhdwJTN+xqjawaOWyfbQ9Z+mFFCTAY+ker8aFtSUBWL3d4bJczIdHgfzzKeU
1uXwxES4y7vd0q5tNaIIxpJfX04wDG+kGcweK7IYI0wBeB5Rogh0GtZJrJjLh9Or
LUIpsepimXqOUtAzphN7cDZ9uu8T4hKYAaHSfTwmuzFfGMaMyABhh2TbWd+nSwFr
jpOe6+r7U6++LJAkfW9KlCemknyctJkwafnY4OAw73IPMRMVcoYdHS/u/LZJroRE
Dc0qFJKGVwI2kovuKNha/I3fOCWlkkYF9vAqJIJbuxs4JJm3cq7gnTpsQ64f7Xg4
yt0Zm9x8DSd8bjV4D/k/0M/WvhxOEe7ZF56lyvxKX4YDZezkM61iiVcXjH34goMZ
`pragma protect end_protected
