// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Eq087OWicXFNQaR+4xFgsuq254QApQgDvsatNJko8NECjK0KP0lrNxRQhzqXsRSe
IHUOTzxrdyE/2gIhgiBxQbveJa6yIWSjXHuc0UDfXCP92QogTzOiG3g4k3LbKMnm
qpjSB4ewOoIpJzjuIjcT4zQDOuBk5sub1kJ1ENzZsus=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8624)
inkUtHojOT97eiwQcdZ2pJnCwJUWTBxQ9nZNIg+e5B+WvSuomNVkcQUTL5+oPv4/
D54RcC1iB/Dxo2vTPo+vXBvjfpLyZ1d+K1/TdVp6jjZet8LnegqJ576vdjJzNrrb
WACp9agEaI1H2DbmgNDUMLoKgutTuiAfXFKRHvfjzewAUY5V+PDCMpw1yYLd/xGO
m3Ei09zOOmsrbx3Jy0RUUqXm6x7/FlH060TcEb8+JVc9qEtQ1xUp+azcC0ID6dnE
kjkZoOjgimresozWdPfT8SWoxsGntY/H46UhFPIZTWRdSqKnRIGWfKBv6Uzh+rOZ
l1k29r7GtfJETct174qYUZ6lguEkolBPY17DnezBxdqMfn9juWo407pL/5Nt6hGC
c9SK+IquMAs/t/Uo/0zqvQnJyMZLEJp59IeoYzCCGE5VK7H1oPSJyRTDVhtAwl0c
wgjCpzs0K/NtRV+0d4E5Zi3gkueSeiaZvVASoOB+ZTvtJf7ioogzPxBpnsuFAG7m
GnY5ALu/tColGdyonRZf6v2jJn4GKn6CtAMosiKOMpQd0L5RgNwyVkFhp/OFoLWF
B4B0L4MKweaboOaNi7haEOv0n2YpWTh/CuhowYe2nX4mUvGQa/yiOUemskBxirn3
OJfXFcyUI8Y8nK+lEPxxKJJM20z/j01BxlhC9o0F9PRL9bDcDygkFiJM5AxC3zFW
DJLDc8iX/6YEam2W0yayasllUAIUeDqbCycSEyR2U8Z9utdn9kjOmC35u3PDPHMm
sQ+QelfASKD1vhLyGH1CuZeRRmsFyOKexTLAxX4Wki0pakXjbcv1W7rhikXEJ+Su
ic7kjJbRBUFkPMpM1VDxFeHI0SdosKH/FSMIN5bhEit5rtTy6/my7wtA/YyUydKg
vDJppFXwbM+5fx4N92YmcD4OznZjo9YaN2W/nGydFSU0HQR7ICTCB3QSs4dG+ZQQ
oCrzX0wmJFm/kBzI1LqujfA9mNqu7WAl9xKIyaxStfbbVna4SSEAv9n6C3Tnwj4i
L2Bpdyk+5W5vaWQkGMzDgC6BTUPQxG9kMUj1k1ZYyeb30SoK+5Hp2QIV1cmV21Wr
fYvknIcP40PnGbNVbXoFIw+/kMD6w839CAd9f46FDDB5DxJDXld1sX7Au6Yx2U3s
+MQqcRN4M1eiTSXQ87TGFtrQk3rNR6FJ4JQ4FQXijVnoSKZ+sNKz9RXzZrv3vXtM
W0W9wydTVTPWEMTxqFrlGQMhfTXkidudWeh9kocXZGhJko8M1wKpdT8q8QzRh3CB
luKI1/TFbOAGlStqdXz09FFXy33PqF+VxRChjua8lh5cqVLkiDmxWJMPFnhhsYSI
J+//MwUDSyHZvxOHAYtrBvlZSRYsJbYQRxK6jAyowjslsK347Y8Z9YFiSNRAvloo
rOaUingxgG0yVGpmyHBitTTzkIffVdIeaPpcn9dIaoPXD1iaaoL7+sjbX8I3023T
Z96D6vJn3qo7xW+le/b6fN6vBi+2SdamzSDGigxVzNBzv1iwz64XtiwCUt4E6EE9
WQx88zJGO2PacuFAfV3MnZdaacjMEl6HxSI0r1/hSuKlqe8GJz2boamxUzpdoC5c
URMcIdAcHttixSS4spevdBZkZeIxavJpnAK5+Pf8TY18s70rdILZxRSfAu0ICYcO
V6ZaTkpV3AKjaJ/kz6AMX/0i4l5ajqnSzY1ukDMBqoKmujMO6HVoA7yO/Uqkq8Ez
3jfBZb0n5LSgLZO0M5L4+tEMo1ax9NfMaNNmqNTy4qPVrnLbEI9PRam0xnt6N2jV
dbeJfPb3R3D4+XpQUzIrH7NJcuIlw9eWsBVlYFPDhEALhSJ3fNoaVViMibtEzxMC
Q/FlcvQzIOgehwB/7GjaEf0QAD5O2c8z4yXkjwZa3ANqu3yU4vtIo72PaiVQMvj1
VHE72AVDPbvyYp8FmlC83MNjCf/Q+CDIRFtJn46BZyUxRqZrK0vb/Tii/jrUocUD
ZLt/hpiKNVyNY/IHulFdChdWsChzaQiSF0Ueex7BgPloxFCXOR4ISrd+S7P19UcT
/A6xMJRnu2VwnHm/8Ca2zjd67h+bHmnqg38J1PCAREHcHGB2H9zxS8Kaj5fTskTh
vAD7INtCg4UypRVouNl9g1mHViWVa7Mc9eE++ynsQ6kBH3SzdeWyPN9MJFT+6eUt
59a13399Oa8UXyrcIBPiWdH+r/LJCjllvgiLlfRLL7zgzZ8TQPSvMTX3HLo16xoY
BwcdKz1ZM7LZBq+Y6gJw55qxqxpKxH/CyLLMWQVtrOpbg+TfSZdOMOBaSEXJRel/
xw6U10mubGS+aA0oV39+Y7G1VMhb6csgGWyqmXmxt2bQAHCQcPR/RKJvI+EHVzYV
qHWj9Y9IucFD2egipRiXzvRUT09NnqOljAOZUjR0N7vLobLn2n7mhavJNv58SKD7
hLpGAumNXs9N5hYdcVnaG05s2SUflaOgBxC1Kz2v91ZwS3Oo/6DDs37Yt7tErrEi
rN+fmg8UV1OEY1k7H+yiFlmBm+7lfJMJrEtd3SzXYUjptC6IP4syHJmrPYOZtvtS
p8DU5/VQGg1ilIc/Hw3RQYhJ00dtySWSlpFEoeoeShNoy152GPp+uyVMN99eTAv1
M5xeAPdnbalfGZIqW4X2U4OjPaBT50MD2FHf17BkpGrF/u9pMSJHOi3sB7Ogbyq+
EwIfopLsk4nl3fJmlw96jG6/i9IHqIRW8CYjcTuh+U/fPqQPixgGz556suFCHKUl
Wx8p2rdlqzKD9JZz94DPapPhucB+DcngspIJDSVty4ZQCxFYcoz2iY1JlMXRKIfK
GvyqgTb2Pz8ga3BQmR68OLiMx3Sm4uIvjbuXJkh6DtbheXeMJx4gOCOlgwn7o/wT
CsxHmy/YV5eRvJuTf1G3JsrVB3Ks4T5F84188Qn3xdlI53haecYd20I5WnXkuZBM
cxufydHo8sTKg34N+T3yyilQFzCCmPGOqc/YAIL1XYC35vw2kmmR+oWfQ9DuCcRM
qp5w/bkjpj6mdo6SsTlia+VWk6W2w/RW2TR1GA8rtMgk/+cPQYazuqcZrHUvbArV
9fibe7YtsNZtGHe5g+A1eAsXsDhZsJlnihFE6/SW/tVnAdRISc6kaCIV+b7M99ZE
VMdW9TjMLZ9ApU+2jfcUcbBjLkbvI5/d9P7Bgy63h9mkiMdWphALYScdcj2ks/Zh
ud2iPa0XFSBfHKSmQur+uOLRKeJcgkyMazf0p0chujVeCpXrOU4Ej5THOajGC3i6
Ra5ZxnksxZWSqXhGKnPxrelzOV3Z8oZJXuLpkYxxFfr5MX3du/lz+ZDEADpQ747X
lleu+eJHeUeNcTP94aSl9kZ1ejd7o3wpb1yq6qwsexENm3f8JWKWyc/LpaHZ044C
Q86/shrPqBtLcUAtd0ppYStKhNAIF8YbmXaQ5XFzCMe27Lz2QqNXyJLNsUmpfaqE
OQy0memZ6HOtqsJjP8WNw2RSwfyX/kelpS5xXCqSwPq7fdwNV8d4egsIUzVFrsw8
WYEcdT5p+Ms/tQx3bSmcsYg3LsDZpBmQnycVjvh4QLapFa74M0BqVP7lm0AusO3B
ke8Up/2VWOybcXtbjcB0H8DUY+mxYRQ/+sFzO3Xa7HFMKs2m/1nLZKXGpaYmXLXa
CLyyOPVDYYDaTZHgV1SQqNoslsvIe3dQ5SdXRYNBtDNxkoWyKWdXWMcDeb3wxZyC
jHLyByerNyENehNxbi9pW/THgTs9OBUF1XjPuiVdCZH//ItEANbuMAJvA8EpJbph
hm8YhxBJpc/Z1N/tnTGeI3modJicjYVfjFzhnHBJ4zwqdsBFmcU8SEaoBORlJVsS
rs4QrLzOHfFjdiL6U0R6D52z1If87+xNZat8/YdTRkPPIjef42iHU6KUt95utUwj
2bIBRbNsHi8HE90QeuuPFFevsEVGbntlT4kd/kpNbFOkckXrQ+3UMMG926WYTwJJ
bChwZXYc5V+tFxdMc6gVJnZSrP5YqoP4pDkUn6LtzKK79eTeufnsKKDvfK14M2IZ
UUr3lM47/AeXcCQJxQXtQL/TZdKxFWyfPBRsJfbDW3MHhrwLXsZgHCpdO5d8COxB
INdor+D0GH6nLrGZa7MFIM0r/FuWncCnDF1FFLaUriJ1ONBy68bZEyf5nAmvkQn2
7DpyBfMIFc7MvSeYFW3EZHb1SCAXJRitM1AqjN+TN+cmGCtC6MG+3CcJ7EYjxGsq
JXQu3jC/OOOUlzZ6yIxM7CjLcz0zX6xnNMgI9iviWmzOPfYejVYFd2WYHAMNZekm
IfRV/Jr76HuwBriR8PtNEGu8qxR5hPGHli4z7XO4NscGa9wFZ0OSR9ITLfZbfV/1
Xa162dy4jKKQakKE1Ub9pUwygaVjiUPO8baxXON8MHGY2D+qyT5+Wa7qR5cG21Im
OhrqsKxuZnRDv5bMvh5TwQYQVY3Ss/Z6sVzeoSWjQK5iwETuWcRzfjf6I+CFfhm8
rYcbL06nTkX8n3N/snObj/zpL/BrHdp3IZKgj51DE9CYtRu/Um+oiiWaeYqE26pt
KMCS9M5t3vh9XobDk0CgzcQzF3usgmuAYgjXtlvMy7Pd3F2ywSSt0oMtqzdJ1agu
SIMtvSv/RsiX+XXe6rkx2Ma5gGX4fBfdRqTIoZA8r0/3W2NObWYF7RgMhUUaOyf6
CC1Wx8QlpYwuSkW4S2uH6Mk84Dnzn4KWIx/C23eCLycEZSkVDBwkj+DCxTp/78Kt
FgrGMge4HKSzCg60VVXJ2pi77cAu0iDVqW6dF9sFWgZyqUwi4dqLTVguysMKXHTN
BKPdW0DD+5bnSajpnjZ/27AwTUdq9iwYoe2j1QIamZt/lViSn9fo+87yJaMSftqx
6oqgDvWqzEL1HPJ7SbDsNHzm7e7+07WGR1XDa1QdgJjTZi8ytBN6s8cqLTSWaSkR
fO+MWo4WeCZqu9t5HUY9UNG80VcOKcesnTHkQ9Iya1aZ8T1jMqtnZ8lsJCeUmuIi
AsvG3BeMog1b4l5dlpKOi1e250ptJi0cDof6vMl/N7Ryb7JaeaJN2MEi3DGjfvqB
Aiqxx7Lbv7eR8lNKHMegvC/lOXDl1bMwOBFDw8CtxFr6pYTd407u7V3xPPtnxWg4
oAfBvwfmBN88yTDgBNvfq1btXdE85FdCw3vz7eRf8FGv2g7jj2k0MJwkyOz1EtHK
5RmiOPDJMe3zft0NbLXrDb7Lkrs3rTyZP+bsEwRRW8A8IiEuIO38T/q0ypVP+vOl
aPr8d/bMn21mdzqpYvAkdNvqZ7CfFeFril5RGVlI/2oLLGGLJYjjFdh53Njf+PE+
8i11VKu/w16O+kLgUWJKswxKVBHwoeKURZN6oQThP/6Q5qZaUofU8nKFtL2jNEmP
8GJbJXGfJCQJMusxCbRN2LUvR8ruJGz3bxxyQVNpll+zmhFfrfchKDfO7ERVZvfR
KQcIiDzHGs36gy1DK4m42ZSMAG8wVtKVTUNrt1Ej8HrhrBOsQ1OHgI19Gw8waKJy
raiCYTUz941PqLNmxzfB4Rd+dn17GrTSgO3+9hy414bNzeSFpqwprM0n4pYK+QpP
YenUBHoqaRP2GWzDVaP2skRxli7xwWeQhf824uU0njW6RQiNLazeyA+490eTW+b8
sJZ2R5n7nIkynk74X5cRVxvihz1cPLZC2hkgiIs5QOwJAYJ7dALBTB4KqLK7N5ZJ
sJmAt3or7kRn8C9fB8EmONOC0rDV3sL1v3iWTRgAi4xiLEABT4E8RfrTb19+A4jX
XkfNEV/zDdvAg9rt5enNqV3xKubY8BXQ/0dbGwJMx4p4WdyRG8so7PTXW9G6Mrg1
WYt0UC3Ltd4OTEy4055cQaiiL74RqAdlCShFF+T5qCViJWwwaRWLDINwSLCkq05y
K6MGlAdzbLSRyaoAnLrq53uJkpJuzk0vrXSxUkiDeOoH9M//8A7iuHPqFmkrYX+V
XCejw1B+qE/QCoYVSip2TrIJ/zTr/2WnrzInTmcdBMrXCjZU/woSVaZNrn1fxOfw
1EDZ7uav0yKA1thD289t2X3BKoygyrkdM31msTSvuhPo2rmEs3Nw0WVWquuBsN0t
wbI6ZIhio/8zKGfeyVGQOO6OJgAX+0VgAmsiRG182I62PVOVwvNZgCUQplopv6OS
pPFTh+lurSmVSams3FlQeFLFjTb5jBfnojfy3Dv9t3tPCIh2eVYvWT1yDDBy6M+P
DFhD12WDpBzvBSv7X+RegvCYsGQivXf3bMyQeUo80hOZmP57qb6lTCplQa7obYLn
xOLJUwvjiohwpHO40DcTmjMkynatn442t2o1bXSTaxMBnXTDn7IkxcNSQtr13gu7
HSo3C33fzydjQF/+NFMVrjVHhiGRZa7C2i8rs+FGpYSEhr9s7OL1e/w7TP8wZR7o
Fzx8XtMGIJPmOqP56Z6qMi9tScEuVH1W4C+65Y4g3h8pXLMnU2kcS7kr5sB9VSVB
vB4Cu7ZlLosgggVnGbo63dyMMB2xwI6SlUqYEMxXe824AiIfRdU4uubHhbNRQchz
GV9xDDx+QWHnqArBKwEU2/ZaqKJzb3dOy1q+a/rQKPuSGsboSHQ4i9x2EL7gMLXZ
+7bFGDCb52sSntB1WTuLtVTAidX3fErjK/geFZipNB7npFHbmES4FGUEYm4Xdd21
rfodUPHVmC8EpmqBFlnPmQgDNTZ/4ElWs/UFMKteALM4HlG6cT5Z6CzH4sdnUUS0
61RHGJv2vUBiNwh4t1aqnQ5iET2ecQKZ3IfuYAeehqZKoGAuvt+OUKFqOa2gA0wI
i+dshnTowY2HiNdlwaICDWodSOAgDhKtTPwN2Gz0EcdY5KqKC8nvoIbazyPWzcHv
bAgqHzrNEblER4fsn9WXlgraNFsZ/dvnfN/40DtsMAUL3cDuwdb+InanFrdqc6Oq
UdgogM1Atsw1BcFksfgYi0k5SCROuuoUNleriRTEWnusowrk+I3mbWLY+27m/xtZ
+nn0Lysx1asKjNjBV0nAPVEj+tuPkeCbuneMkmgrqsYey3+XnsC6rwyHueUEsqe9
c0MHN9m+ZsU7t6TqBUYeZOr1YhyZC9BMwiKkDdLUxcBU8tRogJHqrnZFyjbWTJ/W
P9Acc/oI5m486n2D9Wq2EcBDnqGuizg9UhozsMlpdT/Xir+5WSDyYv1PhCjyCr9V
AQOxfCI6i37CelKD8y+UcunaYq+1u0Zznz8TKiAB2X7Eq38iJUDaJ3KUAaPyVD2R
9TkJt/Wjh0fkUcS8cXeKo60req8zo1aOAOMyinKxD74uUirEZq8Ejnhv4Tqe9fSJ
NRn/h+pDyEObIPmDABJ7uscgN3BmmZ99JNLi3pzBkj8hdm1iM2GGEu1L0z1u+Yfq
OeqSLJP2CDzUeJk7g9Fgbaic10eOuYbMlHtoVkBZwYqG68hAnspwMoU38QPmwcwn
F+RgUnseptwLBcWC9GmZNcODNWxY/UmrCmQCYD0PytO27tnsU1oVUrSKLeBl05y6
1fFbKQvayQh6cd0PaPZkjzMcLM+JyvGnYYKVQVbvGl54lwMWXTQ5sDMOXDZ1U9Dv
+wjnYiSW3IN8t5cm21FsQiJqmDwh4hDowxZR7Dxl8ii0+P9y5DTf4A1m1GXGqywi
tKNVwVdKZY5JKbIp7H20bRygwr9FUwhhFQpkMF96wiKdQB1foJM3r91zgOJNG2vb
8c2BCQQC0wpjZfIYhL4vAin19iy9CbYqkLKnssPSzkZpgRi7G5XI36muW+saGH35
beAIQhAFHdQjqLq1kjkLL/9yvVRr8nEorNTGY5tnIP2I2pnxmUaHcxm4S6qtE5VZ
pe6N0om0GITck0shSdBgsk+NagSv6FLv5OJ6wG/tp6eDCBgT7pUZH3blKEuEnxcO
5A/ozg+EJkRZ/H4r3OZHCWg8l3LGy9AKXmb22XXfz93hq1eqANPbQDwe+n1Gr9u6
NiLgK3touOAkuBy/djyvCIhOBiMDTq0H1wy3Tgk+AVjUcnSDvo7lPmf2HOUjwE5r
Gtdz3ZX7KGPcqIY9PtnkDFPrXgMoGFHGOUGVKLmLyKVzNTAkYxb+VKI6SAI3vKv1
IiPSyYg8GBPySFiDI4zix+RDAEZdsW4A4JNjVYcUtzP+IhNfo1FR0aGxwZ0ok+KF
0cu3xJG8bEc+c4K9jMIJv0OWygf2pUYhzuCIalFZgmvvZZKhdTL6i+mHFO7myrw8
XdCMQi4q6XBrG9l1XfwK4paczrsEvP6aLc/qLAIcPNKC6OWVvRpp8mZn4t354ltQ
RWyW660lhpxkJ37bcD2o1D3LqMDdmDP9oUPOrv6pCY8SiH8GX+aCxHT41vh2cGJ0
/5feSWJ5hTSgUXaWCkI9hDVUia3RDBrmdJ6ZusTFB+Ho6GPTXQlM4xkOciy0xmKD
E6TRvv62bIxcbLQnV0THmxp7/H84cg7Y2hzhRHxd2fZbYvMLq76uhQPgpQiueql7
m6A4c0DF14MqskpnwRk1YcykA+7TBRdcYr+bjra+dG4jdRbdCdvJrSH6WY2SMRK8
opTiK0ko3Xn88F+fpWOWK30c50X8WQwON4RSvOMVQpx/vA7NX227nSwP9jwb7rJq
VAIMN0pPF4wyQvRuT4yTIPsxuEhT7tLUO2AOYG8+hIllEiXLbV3mPBrt13t8GPFV
yu3xWz21potKby3Vov6KfzjEXqQKmnaSKZgzcSRkFchO9qt/kv/KsYPY1zHUB8ID
7qjMk0KvhO5ijCXKOGQ0obmoktOuvInNk50sjA/de77DHiARuP+2v85a1U4hZ5Bj
quFG/5GsXMFZcrsmbnKGEC50UIybvGqAefWlXexhbEhAWOrTJKHjnarh7qhGtvLy
nF1e3UTdwTZbM3javiVQxlRQ+stQ5h4/x5OpAaxpWI6QIG5DmEpsQdTvqk7+THDM
G00FTb2ewJhAO5csrGurU0HlMo0XngKQTOmTkGcaJzB+FkSq0KkBl7FhDiJ4wknJ
JLdgdj/6Ia6/+WTs2Jyr5gA/u8C1JGQvEcZDH8lgYnUExucV08jkVqtAqItpfZEw
ZyZfDDIKr5J4QocHv5sBNz9maq8D71b5HJebMd2iYfjmNc5qHO/guzOakjLyWJ/H
kRoTHVMMCzUg7YGp2YfZjF9Jbaa9NFClPFZDHaWH2IZImOARjwRWK3DAnex4Cpsh
rYe5+3bIzGutR6yrGqT+61YOaXXrmDydlkRoqJ02UiBMZ1fpJnVRdtlaMs7FNh7m
Qp6r4ALKn/K1XLkxVN+LfPYFVWKlL6ILMDISaObKE3fKpvIdMMdhYFOsRRXBerjU
GUmC1J+s0vI+iZ4AOlJMskcKbeo9kgUnBRNs7og0Zm4Ma9Rkv00axES4Kp7M1uIF
EnSotHIjS2i0sYyFiVvHB8A9tjxDBGsAFYpjEDG7aLpce0yN8u2H0rtL4SbYHjz0
0+tY4ffNz/aw1YBoTWs7yw7kU5cGQSPnComWUO0SO9A1W1yKiriluVLC+6tlSNMY
ZSTp88sOTOD8C51LMx/6MBn6emTF1ElwAlp5TPsEst7YpgdpQd1uTUd/ZtT40MHS
9HDMbTGSVqzm3/eu3P0CGI0zxSdKgHojbrrRgtuWrBnaQWIorNBj79SDYWWC9VlZ
iC1YAkfNGsQwToIsIMIrz9RJxTf6FNctA6qkpE+plYzsptN/QZwWk0ZXmYZmSPVb
yWVotM0hb2sSpaKVsFiOPIAp82C4CY3H0BX0YuPrMmHo9ie3gioEw3EwlOe7HfRq
v/SwSynl/wY7/RkqCWO89Rim99+GT7pNw4R9e+154nH7wq3jAhrHJMsmJtQ+8gFy
U4Sl1NGAbUKH2Noz1iDVILt3G8S1gGJwnNEyw4uGpyAAb8nle/DREJkKoNR4DI5U
qGP7opazzNiOju0k7VIM3/K1Fm9o6nSyTDLjnCsMT38J0LZBnPyI1Wpu7vbCTlRC
8mAI7BlypZHgzF6rHPIeMkWjFcGQShi64yhSC4zq95A/zNKUVWpnztTVp4BAWbmx
SuNMCIAlXRHur3Ob+cBE/PlxV7rjmJa9TcioYDpQD1Vki0wrhzhtByU22+SCojAx
cN9fD/6XLNFmEKn+djvkANqDAC5LftlcLb5qqYlPofuTLoEzSmE+zU6iw0/JKj06
h+5UST9eYCvugOzmjulDtHcSpIc4nn17KmxWovLnPxBRhURIt03iQeiAR7bdEy3m
YJlA80n/eiPEs6bBKASp/8bDzAn5a57gI29/9ctvCtOyse88XVyZUG9JqV86Cs8s
gRXM9lt2eGuX+2xkEP8otf6fPlaqY0PbjwrIL3IiiSh5S4+x7eXpqdJGqGh18GQ6
dqt4InCeTSrpecHfdunQZd6Fqc2Jp1dU1lkSsM4FowYfJ7AB7dD3KIgErLdFyfx1
XifZClRYkXG6ywfFQLCRAsD7a5K7NUWH7dzTK6sa5hj+Maw6brf+pzGL63fWYIlW
tHpqI3+hSL2J3B6RuXG+AEmbGv9DdsVQ7353M/fDL9Sgxyk4F1mGqd4CaYhRz/OM
UoB8RYLyXboMaFMlmDF4PxTbex3Jt6+gi9l6DB1POvMzker9PiLAgv0kKg9d2wDm
09sy9n2VM5ypNyyYKWx4KMf7x7G0lPV5U6r8IJXdzlM+Fe06D+QDH4s6LnquYGzS
1uw+8Pr5fqjwuzidloGr3ZKvXvzzylqeszCb003SOCeYn1kQKgbr31+lS0MevQvn
TVXyIYgFsCGisz+P3oHbcreSkoVFRNgiC0QqoVrawRDa24i42dAx5V4UBNfzMS4F
AZ6CeO85/7FtWwjHShpFvz0EXyycnXIE1KU/9lhwRImlPWhc1+47MrGGX3TMMFFo
mNcyw78UHBwsoJAQTNW+biKUfZYkBQDWpfsSrB4+2tTMrwWgqMpigZ7/vrGXMXDl
EqfMeg5GEU0dcvtURDAxIygJsXUsAxRYQakAkEjUoZJbWdWCMWam2gK1xFEiaM4a
VcSIJNyfVzFEr0VgtHe9qxlea0c0TGM4Jz9jdU0iCxPFHbMJJ+cwV6P362QsI5fQ
syaVkX7KBbGXKOdCen3fA61Di21GmLZ+X1tRv2vM3469AWeYa9zbCBabJnFNMQ0j
kjAFfYmHBiGplROeJR0MDJ161+opWTZpJP8qDvU+Z6As5lbtCU3cj1z56ZKS6DDk
efXNwiLzWLqeBiJ+h2sR/jx9fPSwUkIWZMzrpeyoIRCqstZMvZlAcjHze4zXBr3n
yU1OqGhAm1lRANsB0XLdzuU/ECmlrZBhax3MZ1DmDrZZ3VWWzIx2VhpH9ixXjCsn
WB6Hf3a+ndRjSsv36w9xnfP7fshgKhBXvwkPsQkuxaF7RX2aw0KL7NbVBA1xZWLW
cPuTTmPY3EDcXV4sUqANTJXnsfVIOy7rxCsec67w2JPTUYGpQLZV3Ti52L93j3zU
zWmyq2Lojw6MpJgvuaG+ZLCmd3c0da4YZFL3mdTrfQMdZnz+xFU9lGOcWTo37Ztd
ZD4KSJqU7Fe23RfhS5ggYwNj5xMKd5p9kq2DLjS5S0c=
`pragma protect end_protected
