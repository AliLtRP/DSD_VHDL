// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YxJ2SObTEL9Osj0zsjBpNaZ8OcZ2kcj29WOLi52BkezUrFdqdLGrWr7aDF9YsxfJ
hTXKiPvYB6WmbI9eTydGLThDdAOcW8iLocskHblSFTS7GdGyJ0yroonYgQRK+hlY
mZfZd82vb87wpKC/VaQNVjB6UazJGoZOsNW4HVbs6oE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29296)
KZeqQrsEvhzATXomVOe9k++L7elZJ3NrsAU4Z3fBhCwJ2yefAx+cV/In5MDx/ql2
bChKKYUf7ZyCK6p3gxkFDrUt9MgPku7jPVqQIU7t1ajmAZWf4/K2xvYd7elLJbSv
BjDVtdXAJt6XomJhQFCGVpoidS1084L9/4LmYOX2Bj8SxuRyAQqKne5gOc2EbpQz
u5oMl/S83+okoAQEdeEn0q0R0fTIT+KTVQb7K9vZcHunf4b6OnjrPLzEkxAINrhy
eele0zkMXJ7NfPol+1rfSsk1OxV/htxhnKQKL8vW4kY4tH/v3trDsnAfumJLu6/w
wm8UQlnZUGmTuEnJAK8LzrAVYYrvKOLkWDplY9Cc/AZmpRX/c9WuIh/ShgRxhGdG
9fuCZ3HMja5S6hV7mWER+FGSmMR073EeWZn9ilkNSsAnAogYsKzoV9e9aPYf8u+x
AYn2jSv9fenweAO2nqJakiqGCxfWEvD7Udn3MtfB7Xlw0l6U6QwQYTRnLUHrP/wV
9WSIXxeyccJxCwwN/zKZ9ds+E0N60o7WKhCD8m7VfvA/ALzVDQykIwrXiOal9RON
Qz5FJ65DYCyiR+jfH+zZQpbEzoTN/KToVHA1mQVXKmPQnCYAQ13KW4Jr6NF+1Kwv
w5iKeYjG/8u0ryyondh4ni9Z8YT+C2g84gWN5sxow5jY67cqCzE8B9ivQO1dSwwr
zfI/E06F0e5dL/aKcjRGJMVbwAZoD/iQVhw8g8ZjzHHAbu80+D9BQMfv0xBryxxr
ziLQmpAYVUuI+yTHioP2rt1WN4ZzJoj+dfA5oYrZrsx5l0Tg1QHLJhpOsdntdgFG
jNKn7rVHtbUYYf7/jsBHqx9PZnnutB7i7E3aIRx/NjY+ZiyGWLkazgSmwlVL1wL/
ZHkgouCmadtrQvGxF9lc6iaAC2DARi0TYZ/kVbGzeBwRBHcpVkyRYeFYnzU+vvck
/PELEuJ7UY1JZenKoPZXhS0Kk1uFZXk07f//gkXqMl8od5jAlLa7RjT5sm0a9dlq
s6utz9uyg/UYBDZqCD/jGk39vNoqrTPTXsIuWT1UPZ6OlGM5kTUsnBL1oDzPLyz1
oPeO8IFaCgQem9UxOLW6sVGZOodnnA1ZqWsptO473inZ7a3vLIkMNCWhTCuS1BCT
MNMDe22NaNHcDZoc599qI3ojoD9Nb1jCqFKp80NMxfRhoJSGBObXTtqLSzLrdkn1
g/c4+NfZdxM7h0MomljlUHUsrIiIc0ETpMVBUotvE/MhGRmAiLav5Gu6pWDLqR+3
+uoK5u1GIsNO9jY6t//TCrb50+Ae6+TOrOtkiQ/OosH+MIuCnSxfPyAeQHUIu3tY
mqmXmq6bIUbqmnVyMPpN2DBHu2eopIvO5MAfeV/2/ZpaOolblCF9OA4QiZ+blUHP
jzZypskvhsSPxR2PAg/i/fpWgbX1HPBYAUOYqW4V2RagstPwSxOeTpyD3xn2U37F
cuvhGQIuLbb5gMHhm2zqUQEg+4+X9Lm9Zr/uPcYdnRhrH1xsih8XDYwjVNIEMzcJ
qmdukiR6H1i82dqX4foTPcM7DoeyuwgnePIQATQtVyrIIXUVlBIj0nnqwDmc19DD
J6L4iTLnhhmh9vGIKc88B2d3pjhskPVTNwO6YzTi2g9SdLjrbqoPKuqJf6LqxwgA
CU32KsDdAQ+FfiHNWArr2jgnqMKFtXD1cCK/azNvqRhJjviuHfznJr4Js54A8JFm
0qSPtBvgTHoyKX4B+C4jL0R278mIqAM4M9as9n91BAPDkl80bxMvLC0ribVTMnVx
NfeMd/omyGXfGoe1ZaFglRDjna/ImT30Q5qUbpKd6M7ASKTXcm+yBMklNLI4bbtT
LvYtS9vKTvA+4lNyx1OvJ8TOYlLuFJcG/VquqS3ebOEvLK0roac0i1dMtomZ18kK
eOSb35ZnwOUw+QrbvDfgwI78jbtt89NLsOg41T+tidj+aZai4Of/hec5C16UbLjQ
ZdaHDOnu8atOuBmafkpzTGMUXZOods4eclcp7p9dFUdHlocC2WzbSD9XuybuXiug
LesGMICuVQ6ML/ack6H2YvIAiJnwtix1fPYkA5RYpTnR5Bo6p5TQZLcqDGDlJfTr
J+U3CrW5JKB5QglNgD02YjLyMwT10MnuuPhUsQTzq3cS8mfHQNIChd5Nzetj/KQD
dVoue/aq/a71aPOhHrfH7LJSrI7hYi1DAr15Usl86GMy7FMVm2doKICMI/Cezxp5
QWwhCUZ4iYGyChE3b/MYPNk4jS2ohBR9NPXhMf1hodPsWocwRGen8pk/JXttSg/G
Fhqc90LF9tg72bqw4ctEbMc8UrSku+NATMWWu/k9kmvqSFeGT9+cvucGDx3Ix6jf
I8RRQ2rFOXc1C+uAbqC96cQbFsWYHNMwq7xM9G1h6cs/VfiXEaU3zEe7cANxiwF6
lU3TMaMF4ysjFLQAOH2nSZLuGqNDfnLUg+cwDjzgqAg5sMGeZBOeIJnaVBgyzEeh
I2DYtDIPoSY7MJL5g3rhvVA1kkt26IEyKrI5HoHE6Ldzh5myxyp1EEOPYHIOg6+N
B7MUXNMbZ3W1qKmR94O8MgWfbNMdUZo8gkslI+znTWfNMwSK8Qs9bcPbJWncdrkH
snjXnq1qi5aZW+YZqfjzMPp+Yx3Rto8Dh6EzT1RIpbvwiuo8Gzjwr8GFFzYFfRJh
QyZ+dRp0I0WO46vuCDWPNeZDt3AHHzDyGg/UDkxICeTtoundgOv+LOLhs2tFvuTq
0XvqiaKAmyBO66JDdVlZYuZyDAnz2/haBuvbVmjGuKA0wsgZOV1mXpMDQYiqnA3M
Y+KdnFZJjkjKFdB8MzFXOn/eDpx5O33G4w0zKSphQ3JE+0UMBaA7csXhqD6t5Juu
Cl21sbeZIMQvMxxGVDmUFrRSa8ip9z4Zzn+qqKn10JLhCYZuZ2Oo2vbC0EVakU0w
TtIHkbLCZb4pwyyhmLbmXfYMhBn2QvEIYz1c+yrdnsBMCHxKNfDJv8y2eDEl2+l5
LDCqZixl4Vtsf9iUb2nP8nkkPGhKFWZNE3aFNckTQLp+FBECF11olbhjVPfz43Un
6KREiKdBLRBvjj7GTZUfEOQytVRu1q/ug8y5z4o+9BW94IQ7oINLEoMNnsk6VDqb
sn7BKQNdVBFPYZJUjErRVSJ389K89Tq0k/WB+Quc8wCyeGc7O7YDKUDjw4L2x2sa
BOeYIDfF2Mq+BSm+ZGG2GmQ8VF3/RV1+teGZCGm3T9RAUoQ6fxCr73i2v05Lp4ZT
bs9jwLmtufTMY1FMPQBF+kgDjevOd2KXOk3PQLtuNi4HFmvOCMmzytc91piReLhC
Vd4T18m9SuiuRIoRbFFAQ/xP6nHbbOrdcTM4egP1Wi1oRsHHG/LJ31KjuyK6X+gk
HPt0ogyOyrzOh1V1M7/WjfNRoSxr9jrXMNbILmB+qy+dQbUA+Du7JbQkOzSYM+BN
YnqcWtYsDpL5/H7R8aEQLP3cjV+ePVTwFAz6pfJsrm4LiDmWtS5H/ZntZIN4uQO7
mdutPcZV9jo4Bk1EB/NVmEUIz433qof8+x1RQH6ts/CWniHEaDLyYfj068c61yUP
ZOOKZKyp2xUurd9zYbRe+QgAFLdjsOew7IvjwwVXK2mLa/W3PiLX0MSFHTRPax3C
IvzPTGMcPGA3fzSeL9cqfWVpbsIS7CnGa5u58df8MNgLTZq//Pgb+q8m5oz74QP6
EQ61tRRrAd6axTSIg0GkYN9BVExfE8Vquk4XrKvrUsE+yXlr9rHDcxMDKOkrJk/l
iEu8A1/w6P7wm35GaR569oGCCV7eb+KaLT522zqmOLLY9eusKxbGadSSuVHVeWqt
JF71Ozp9Nl5GUlRDFvSayPVuxT7W6M5nAcSwIqZP+X36nK4yS66KXVZqbHQ4aqPp
VGzVvsqg8kQN6cWTNxMlGB1cqoQJc901dVD6I7/Zy1lQ48E5jxJn/Astx/BH+75w
LofIWx6iLBppIQjwhNo8lH2eDU/P1doUgfA5fw3PM+4wXIUUM2bs167g2wpAzU4s
SoF9njJI7MKWxMG7A+fuVKtv2yJed/UbIurGexPrirLB4i370Hf+3s2lmKDDS7Ov
5lPvFdIhF2m5WJMCchkOy9idEEvPD+Owv4ndJROr1qD4Hw2zf/b+Y7O9sFEKDrne
cNlcZbtoovNUUYbPpMkLV5K7S5ZkpYqBJA88dKp56vG1Ijvg9ZEB2N0IYbjq1u8r
JvndVA/tEzvrhnehBkv8E/cM8aizzH6Q1psHCrvyW/dn7aDZ5ZngENsQ8Ktr+a6N
uwGXZksDbga2/2mBhFAw14iDR7p5LpekLPUJkY+cMaetSSoDgVgrErvHvAOgDWqH
eUulOokvteAJxzprU6u0Ep4ej91LfiaM/KLRDGXs8cGBf+P4prA0/3NlnEMIBfAo
7SsI5UAsK+GgHfI/I6ZhY+m+FaCcWp9qdgywqBHut/b9cpeDlxMH2h6eiu5ZKAmR
AYr+buETjfEdXwnZUAn/OX0cR4jyWN2Zws2FLw97AjTqhG3Fcsd+yfXvohicsNzB
DR918o7u7+eF1NBlo/MdsGxSpnQ4marcYHQIGoTfS0qk8ZDkSSyBphIjEuW7wG7F
IG4NnaNxk1lflnwFJ/tCoSVMRjkb4EzOg+r4mWB3ijoYy5rJo0c4edQf0ywF0iIO
FK43HBbsuqBTwkElE/Eh4Z+IO0k+PFW+Alh8svZg8kmW9BzWX0+RkdaSuH25uqO5
xyObZ6tgLU+0esZd00LXhOEyAhERv0HYNKkbTvdTodaAAGfrK4CEfbIf0u50NE3r
oCC2havWJfTWPvu/J9avWcE9FnVR7Syy/YTroFbZ/p68BkmWNLtlwSG9SEreq88g
IwFjmFFar99BNc3i8PcmBf6d/XZL6k7q/HX97tCFKWb3O2Rl8Ul2VvlPxm5o40on
uC1WSi3T283xQ9JAq4cYIB0OHbfeUkKsbGRVYmcYNKbq5dc3oUOqmmxwD8d/C0Mn
f4chJcaAz7mKuE5NXZ+Jo3CBaVoxZMWA7JkaG5+CMMXXLVEhEBr0NHwtBT+g3J4f
YEOzW7ZQbbGX4g7wHxPlNYC20i41NznS+hLrJNXnxHxPCLV/IPa656NUpp98TOn5
vyHMECZsZrYRvgzf9osp2JYMzsaLe16XkdxRyoWbzomshM/YJslEWURFZ1TiGwPk
iLcwu6+FFnOHxUX+KXgQnIkXfWrfiPIxnHjf5jGrZIuJ2mDe9zciyCGfgAmYWCtp
fLrilRS8Gw8HXCjpjtwufD7GF9kKeVhUTM6B0PR+7vpdblSAt6kBsUqAfeu60How
siU+uPSv6hhzp+shBt3xesx1mTMqgB3blVlTVyCKI23mJmgZJGH7th6/2trJOjZM
3M4HXGg6htZd0CDQTDaj9r14MOQHatN1W17U60UdilOF5VKhZIk3M6qOutxV2/0O
CJiDoMI0B1FwSS9ClG6QxbCw//3avDX/KifLvuLI4qpOhyL4lHlAIiM98cDPjRft
md5HRoRcKvzO/67FL+STP1x4X1SCySNK3j/KLkGwAjAOlrVxvZwWFCrdKdUAcey3
4UEO8nQ1OL4YFn/iRTPfIOKZlgkaZZmJ/ouxrjMud0WLMT7BIDojSI0pvYzFHlYR
KZfyFAB7axpGU09rRtHv8zDj0hYhabsEAkH6e2I28CNRRX/a//FA4go8YNYCMNsn
5FSHgMDnCT0Qcc1523dPdAnQxnGc1p3DthutIKjsyLF8QMO7QBha1JfooDnhDpgi
eTlS93LzdquXwwROwRZTZZHlKVfAZts7TiCBVeqvJLsIurXonnlmDM/yvaKqDH4T
ttl6S6eCu6lD6ewkesUIq64Dm1Kq7FgBDFU6R1MDnELUGS/qkKBNlp7cbHQ14MYx
Gs+ZLRMeJrfccfGff72zTV4EzsFAPn1o/Qkw42wG9euQUOp1DUV5ioEKF7hX7bKi
fpk/jQljlp6hvcoU2oHA3uiWnDUHhMsRcr0zv956kGykAY0XSLeieJdDiUZuCPef
boutgYx9LLudQcGPdSGp7D0DQ4j0a5sycJPfU270ByWrbWuk3jUeBuE9b46pMq0f
NsAFy20Q/yTo6g6SiHW/EMSbIwqxlM5exTEsL1hv68ohYvoz4zBT/6bRgVN++W+t
B+xSz8ZBzzrgg/9Pv3Pam17ssUk53EB5lUyF9OnbRP4d3wqvPAYiLDzxUZy4WEjW
4ozCs3dKICcQBrwe4afioXkU+ZNsYSyvysE9oEqfyqMjtdaptnY6hXcaSHjL4pi7
G2qdk0fpgWvCF3Mz5lwryXiHsKog394XkbmDqmHaVrt/WNpu5QPt1a2g59L/v+i1
rmiDJQHCXUQPHqFayT9kXBGAJPGJIB3ic5OuCnYE/bE04PIL+c6UMRxHqX/Pgm4k
hBNNXNOO0YmT5A43JaelIE9gNfqs/WR76wlh0BGK+9eWzzeBb3qSFt4t6Dyi4rsT
ConwtIskW26L5XeH6fsNlcLe52t7hz89j/YyfNu6r7+sU5klJZMb+i5KLhTWE5yJ
5GpLo5ILlQPdGQ8/K8nWhj4DSjaIZicvlXMyhiaIOpQrl2Gdk17Gbqd1ODCBsTNn
WZg4ZxUK3bQp+fMRJkJSAE2LAB10/IbL/2HrHjmFDcTs9O1qNql3kuRlKh6jsjyV
V9ObaXtUYAETRVwCmJoGJCv+OH2ZCfaS4SJIJedVAVjDfLlDduMiC085sPSdfkBa
VM4BnROr3kNU37+Y/gZm+TyvVdNlJjBl79HiVscJ0j2bLUmhNZ0Bv1YD3VJduIXn
PkzxccWIQH18+EhvgLAjifJDkEM2OVTgrDG0OfYyp0h1o22LeZERdpbJfDW8nKWz
OxsHJ8aAapcsk8FxM44BbtqYVUw+qDq9Z3uSVDGZTq7gWcUb+7bLe5OqtR0VffSK
mOqn3UhnhFamIBahbClF87+oOAToRGejAFjGBzMx1rVf7d+HlzhFCw0mb1RWPQNM
B7zm6VcCxE7ZDLG23flafh3w9KdITLl/9VWuoG3ORstOsszCZ9aooYDlHURP4iV3
1KcX73CizXUDtG9pR1b54TzdOotQlWRIWG+fa7zzy9l6UgQdl900K7lzpqgem4pc
a6jYZuxLpMIo6CEvJm9ivA+blLR6MnFyCDVFRzC5AMvsUcug3/nbJSIgApYpH2OT
XqFEVw7rO6bWe2cV7YokUMmGskU5JkLALV8m47yccroY1QjrE0WBY2Nic74jZdAi
BVM7pCA8j96jC1xe7xxEIr3+FHhxhf60l9hckl9RHSr9Pw1n8yj8m1PN6e1OdPH5
Ju0glEVGK+UjH+6uTgkd35B7OgBzs/pTp9RoTKkXG2uM7HPFPanbwDJ0c/E3G2qi
ESKqWjQrenokvSaxpFThwY3UsgWZCVaMK+zPmXwdmij8BGhmu83fom0kWO7c/38j
YwiJwcIW658/9cj/inkAjrhla9qKfMuKefVmoGR/YS+m4A8+qvvoASnJ5cGj60+t
Q4ycyMgrrFarIhfG1aVgU4SO0IQBw9NBXrRCLz2OHp5SRirdHNBrzAswKIENdWFM
VCbnojQ8kV9jyYNYDoa0Jf4v7e+cFS8jbQQjO5Aexg2oSzLefRhs4DXW4V63lL5V
TeDowo7QqNflwhlrKHQWBj01Dxhu5yjS6hSEDPpEL+N55B9sdf45gRJjviL0wAoa
hnIOR5QIygMIHiZMYog2+4JPEAwXv+nJKnrILCgmf9EdHtMGKmmJGTRjxIWSsycH
j4jT8QHXzSo/6TT03zvprYkh+Cd8xWE3xuQxwuUgtLNgozEQC/TdWaM3smMTSLcZ
ZmQ5OO6FwtH51JCywB7enw8C/isFg188efyzoNnDo7bEjazt9cnOUmTLUXRGNLWR
bD/4PFkxcDZkBaJssNAf3EY3EA52ddPdMsiQJ3VCCPUKzMiv4kG5YhxNqsO5lVKo
Tuma+vnisuaH4A2KsfdrpuWcRrWHkYfhPwVRRo8tnoDOtpFQOWadvd9P/kWshr5p
F5Ng4yCCk7qf2L4NIvyg1h1eK51/yOLfCP2H5YpFvjEppLPMJUP7rFcSnVYKJlsW
8pBYOev5AIefYfQaMAfy80ymwST78vtp/30Z/apv9DnSTo3PdYJiN2UkwT3uEbYU
C6RlCuHnQ1q6STMfhTrY34yssL1yqSXC2WRCjOKWJo+x1AazXcB5j5n7Zy6M/RRn
oqezcxyuWQZrljx7NxHlRH/C5jg+BBgE8+uP0OUgwWLwwGBQyK/MVc3fQ75KXp5b
9yXCJXRdXsurWvlPk8CgI4HkgcYtKvmStRkb55Ch6m8BdjrozAalKt7+pmIa80Wn
8HyKMs1Xj4nY1/WEiTOuQDbDa56bnzSfZe0dUZsasm/xyEh6p2W4sCJKUfq4FKN+
wGY7FIXfboNoUQoCCrIX9+lhnTWfO85glymA/7fM7ep+2vCWots/wZ2ttGxEWdjn
yPLWkI2ew5h1OMPCRsWyWC1sWFLeJI1fg7BwE23ZaOiSDgOk+XdLkFz137/VN5AP
9TZ/bHWcYO1Ww2AEnWwFrDy8N/YLX7qysB7V8l9TV2rfgr87qMn9Qvfqm8RanfXr
LmcKMqd8P2SFhnWhigceo3OIUjyACOOekg/SYOCu2iRGgVppdtj+OJ496hiQBHTB
TD2dErpCSYNye0SBlKonx9Iu5D93eAi7zGBcRcN04g4BZox16jKGvZOf6YMDuHST
qBeFzRCE9+06cgeamDzJoYiyo4CS5ZVT1g33b56ufswZepA82HZLrU/8VrwNWhaP
Dp6s5mgV3ChbkncflHkrWTpx6/sMq/pFNmcSDvGWiobzC2UBgdo6Czxt5PrK1jHw
yMF0Mpqlqn5TesMw6b78uxUxD4Vq6m7wCQPU/u4MdZKa545jtWWmyUFO9Hel1aM+
MSiQFSiwrhiNyYGGsMFowsgjRP2dDRXQfMNngn+eCjw60XZjQXXPQUcfPje6f9ng
i/CQjBlK4CZ/2vWVZXTo1++BE5ZH2F1r1aN3wBro2YyhNIKCp/aTdRaNiDD7b1OB
7hZInCP+dXmZ5VQt/oZgaRL8ev9lTRRA9tv7bUv6lndZZgNmixI3yaDW62dvcBqw
irxHFh95QVSKA8ywbQXxBJQXMTQ5JmlGbek+xfodrJ0neLmtM4qTPkLW/jD7Ff/q
bcKC/7WP+ntsnn2o8znaY9aM9y+tvBNOcDvQfv3jk4fou9MPm0dHVfad/xe6cBd3
5nqgqKeRUrfqZLT8J/sK1KJDjKYs99e9zJEuPg5oWy/cUseKicKKh7xL8G7ZWJWl
vCgLgcMIp83Qqt2PYPmQh+Bty/dAoQGQ/Fzp8pChzsi8NqFhIJalOWue33BWRfMf
OLnIQcDrzDcqFK+QGP9/pkxZEwo9a6MtjL4fMUuWMqc7kw6G7TZ39vEyfGwuewF+
vVhhXLlJugi2Yg25qVYF8sCqvs9ejuy6krseV9U9HiYxrXRcTD9HvMYA8vuz24+n
46vn5QV8R1H3h8AOyfDPmv5OaV2hMZQlZynVjEOE+ZbQ9O1h4d6fazHXw28TyxXU
Yldea35XxCQpbi4Edja56gbqsuVW/LKlMV+Eb0iQPXG1wXmD9W5tTHz2UQXQRM9J
iweGlO7cn8WsUv2/eCXt3SrdLy8/Jc1KFEsbMq1KRB2JBZeCzKulpC/nxLPBsU4N
K+h3WwqWm+w3zesbq1+e6c54jcNYd2VyYKX4QDI2/8uSwNtC7uIi747y2CaU/EJq
FYDuEtWrgkt4ITwNGJqDm1JJuqdILlXO3y1tZk/Lor7ZUee8xkOGufO5AGqseMrL
DRKoy7aqGy5rzJQ77umbwMdlribbm1KHb1+eF6ekWg7E0G+/FgTlIR7yAsSEkMS5
mFJDEXkGyp8F00bXPcIgrq15QBCYZtP0BGI/EctRF3BHtvrnPQCI0efkhgGHasAC
40wXrGHZejOboFAAmkYzVsTtn5tqoKo3MB+WV1VBTKmXgkWBR5820U4i+XmfR5q+
51NVETBgpk2iq+gmtZ8UIVderFolgxeag8hNP/QOXocLErz1ebk0ihR9obDAuqln
51TB/8iNIS2P4AlJRocgxsK+JUcpPpIJywpmhC+XGr7H0nArbmHhSdn0bCVfkxyf
mlpN0T2NaTPvwuJmIGquenXCtsN5dkoSk9HWHNCYqhoqwDGsAScQ81i2Xn/mrQls
PEl87f/PiUs4jCTIL2iJ77NZTYDjB3vZAQydss3JTDRmCVrUWrOvZssNGlX09i+H
JurbAcga9A7P/IbWp/9QwSU5clhgrbo2j1rlRQE8/oKmqrQn+fwhcNbWH85sPxU/
QVnCKzTUMWuA7ZXY83PfW4uQYfrze+j87lW+xqQDfKJ/GIEHNlWHkhcYeYUIrDhg
PscTDweS8FJXb2yfGXCC0diLZGUOxcYV4/ixZCh7XxA3bYeEyolQx8GkHJ/H0oYY
Nm/B1n6hV1Qer+So9JmBVc/VFHcisRDMcMKmrkkLv4Zaw8+dbp7B9qthH24V7++B
si3hHFbAVYIYwqBAX8bAjw8PmSHqX+5QTpG68t+AbLSgImWtv3XjUufxkfimBvoI
8Qz5mPCUI38MzO27u7jwZmL/MEwgnFMe+xi/uAKIFh5bcnp8ndTXDPV5taou2n6V
Mv+DadERFqfw0FrR2MnTcXAdvIHSAxCHtlMyB0mIgALljT6VGyQSyQ1RN0HWFBrr
m5NYd2LsF4mdYyZoeyW9Cd+XzIPyxZEgG2IUmFzp205bNYJ7Dw3s9tB7HoGmCSTY
ZlS57ay4phrrqhfEb5h0vDjcrolOHfNsPCBzn664pmSx1NJuuMudRmhEsuK+U+W7
kjj3ARj/xPM5OTqloq9IdEWKTCN4dtahkk4LVM9QqOTXMKF4NhQAfI8SlnBPqG9b
TMNnfS0m3GaHoLJa5AWqmzgNk26N2t4ECEbFz5aY5dBaFbRegHQEjle2cobAFc5i
XniiKCT6y1W7PHxjUGaoYhTitBG/FI1A9JDgseUyC7mKmC3WPEZKNyCOxRMjtmLz
eMlzlipyoYwCigUrM6Tp1uyxfcEu0BnircK7zc0YnjLNV7rvHc/82FIQAdn6MpHP
Wls58Mhi5ymhlPzgcvzbKWwYsFzUEeR0of4iRjdWdCr0ieG235RWy9ouwpzSBKZy
BVYfjt+eNluAxaVVJfupD5pVHYtuh2cqHrnhMeD9htqY1pswNvCasvUeJUfr/3aU
uPlon5quRSjez+3vTSJW5WEo5Hzrq3P5o+13rtYwJ6pCi2PwL1x3WG19eT3/or8s
Gs9jK3Wz0+0SCqNB9wbPUo91ZEDtvrwlOSF1OXT+WNF+hI+ceLBjRVqKgF6Kwii4
pmeTO64aH4thDfiCSBtW+rNggv/f/CtLGz5DJcOxWj560tWI31HLa9fxxlrpnq/w
Mx75zFp1pAm+DyUY4yTNNbYKcuNBS8tNFDM6YTlTO6oDBvSoJVhpri16Mdtfa425
w5l1E0YDLGSkmEM6NwFDBJVYXdr91ogS6ovPxKdDFB0j1/yrRzN9qOoJZxqNkKJI
q/SRnCJAVB4g4T4TPeTt27WmZh6PusEnj2oyKhbjuVv4HiSdszuD8hRM4Hpysnt4
rjZe6EHcY21nD7UrzQiUqIWHYOa5Kv0pl2x8ZbXiyZs0HaaFiTQf2z47OoMRtO9l
KPJoClHA+E61XhrgYbp+f/WXLLhqm4xWoHnM3GrG1iK+RDRUYkZ/J+22rG4tjAWI
jUkKxhJyN9jml4qb4GHconohGx6a+rQtgcVZSow0EBUnzy+XWq/LAzEXvQ8wsBmJ
220+YkFSMWwj0PbqhGPICqkKus0On+cfhsBG/fVoAe9Ku57Fi5cowbxIyLB8GZpP
pxZQwhT4yXJCTduumT9Dh8pw59Sgtn2NUacDvToFwHiKkJ7vQgCwV0OCFjKf258T
qdZEKauxQYvM49Lz845wWRe1pfONhz4Or9KlLJMeF+GocWTUmWbDKa3CLygzQm+y
kn+fc+zhLM+54TJwteMIOLotMTaM3GhsEHK9tHBJJmgmPlEyA7JzFMAKxcLvkku0
GiFMXWfI1eHq3735ODs6uMnzzF1u4qJ/cfKM5IzUv+FGRUkV50cPHxEtmnLCElFd
U9XdL4v4HUxF2HREI4nD7MS5Ftwt6I0OLNq4KJUf1/L6xrHzBGYds7nc16ZJirNQ
jp8ND+Siq0d6V0kC30nfLislqjF30bxFhKldpVRyFHswQ7nxP+XRhebbdB9xQ2kD
GzhdWalL2faQ7Q22NdJE/PJ+WfvUAA8xIaKGtuMoqXHoX1on44FkaH3TYTwEOE1Q
fIDPN8tBh+i83uXyV2MAHkQtD42vZNw+bzd9aDNoY01jnJZoCzY/HGliGKQyUXq1
le4bojWVw1/E5N0xkgtqFe8SYp0I9ibzna+CzKM+QxxfpXJlt0T66gRDO4Dj2xZz
wlG2Jk4tEHBltUsM0eLXkPxYsiP0xO+oGq+eHSi/x3k30NkgFgIQAGLnF7dO7duq
ntE/K3Vb+5ebf1pU5kid2ZTFklVh7ZSwWcpHx/F2qs4W0fT/UmJYlianvejMMH/f
viMBuLV7xPeodR7I2CjYaDuJwiea+LD3/QxuXWvHlif2e8oRNnibBmC6lNDJZM/v
Pd4bWTQ+7Xzj6gcutjk5Du9KrmAqF1SD8p/+owccoPE36wHY1xFTiSRjD/Q6dFo8
2/NQwpNY1CWkaYyCaHWAwK67/MxV9BbRpC3GaHTzFSZ9xTVbiTWYVJCXjQ1JpcZJ
xqIpB5AGGoHBao2aYNSsHEXxmdPeq18JPywuktLQQzWsSFqY6lupoT07WdhBMXkp
6GNZ4m8xTN3sPWeDBOevXpJlSnAbzA5gxvaPcE0GskE8bEx9tuHUamPCoY8+4TOg
o5GEDIL4ise7TPb9FurzdTm19P3rBPiTk9KGdm+p7e5Co4f33QzW+xFXHp2zXdUY
KOE25WaPrW1aC10SWkMW8TICDK+e5BJot3hfWCA2qWEtdCWtx/n3OWGz44ybPZAs
q1+k7sX35PTF3xaeHtvF1BfaiOOAGtkRFYaigBvrix1Lch/K7CpC7rRXCXg0zZUD
Vj5tHWqp6iUlAGen+mP5EebaIHIPmWg8e2Kb4UDy/Rd4x1cGgircsau2Jk7snMlF
YtCJZRLJd2B9lopv12dLqh0HqBe4GVhtYe5U021XqfX4QWWX8tzmvjCxMmIkuZuD
VZznBjJY1Wt53Eo0qVtGgCS9EgD5ZW46TWsxcsDU8bqp9L0CP/upSH/dVOf1K2f2
5zyaymBl3yfB9zkrZ/fSSdMhSODpogQIcDNN+bvgRHvt8POIkai/1UjjcR6+uOot
+cyuAiP/VWyVmMXV/rmpkVbzHTCHtRuOgsxAhFa/I8AMImMK7gRMXIyCRwAna7bs
3yV4H1zvYo3QwCitRIue/wdBZ67DfwEroDbA15+YskScA+nItE3d0Q6SM1t8r7jB
mqbtgMIBx15rBuvE/5/2E/8MwFnUgJoXNTxHDVsLePrGKum/mH1aMzmZZjv9d1kE
vZs31NrLTAAwlxeXgUWX5sJAX7SliyjIkP1cmR+YIdacSqk1UO4nG/cMCGlKzlYx
YL1qEYWW1T6zScpdHIBZbstngzA6qE37SJcvZH4a+pTvAAmRTaitJGcxfUM23hrK
SlatAY+VAWfIih3FNTFCaA/84F33cUT6r3C2AnoGbto5TXYFltGtO9ZUcyimPO+h
Xb1HN4trswE6lYXAzc6PwFk+kE3V44YZ+zfl+1WbuI6wkOB8Ht7b33HAqZQBThx8
aTt9Hd7dxvSyB9hyFStGbpv5uuYSKm0lLdXuDx6awvhj1IO4UJcv+Zmt+rA2hUgL
WxKX81bVsrZo41Vz6BTiNZAaeHYFwj9LAYUHZokKr+ykUZGv/ru5dC8Sae9mGUmI
hsXGacfS4yeInrJSl/Th/3uxLIe6cO9f9uuff+4V5tyK/caiTVGTjEQs4NRH12tR
0h8rHjXyNHcfvEku89Ztor37F3Bjo2E+9Q75KIPQczg5sFACIMBDNlKz3ib3NoGH
wk+Vvgyg/bLHQpwd6eg8l5ezE6KZM3uoq2hsAMz6TMd5DpES7dbkUSuga/Os20i0
5QlixPobKWuYanDATxPN3cRcgso2Ad3uVwdrruf+FzCzVhoIYwfdF8fL0Rbd7Cem
9bXHGDsogwjsRuuLKA2UEQaOS9DQ+I+xEuIFE+Fo2fBo2L4uuzCBzrXCztYIk7Ci
H4cM9h9LW2m0Z9r1KPIFvTHcMLhRHNGsWuhCMSLgivRi3NON9YuWj3WWyU6Wc4xY
hC3tgkz7D+uvqvisa126lqf0gHfExMsfOah+l3FtQOHzJid0qHqth5YcDGkRJnq4
gSUVBm4vNoHMbYT557au3eJXYWmjnVxYwXRmAS3TGTRqWkQo3jsV6eRyGf6dyRlw
al1zAxcN+6qTXfe9hGzLxoxeBFYWb0fYURx86hGE56T+DYcxD9nO97SyqVG8Nvuc
DmOmK3xPBClg5GMBmfzc6EYqQjBwwipOfXslO9CBpPIOVhOhVYu2KxUJBLlewytu
SOWgq8UHOrgvpHe0R80ENun5TVmSCzgaE62XL+T7jokHDuvV7TcZdlYLW0W8FhBj
RLmUJmrA/yf3EIeJzNToVfCx8NuKi9cTjIoKU6fO9iAZ/47I3qoLwPQ2xbRFlaIQ
yWsP8UqMxJ7peq3d2IMqTMnAoIG+yJkXOWjtN8fsAb/nQfVeOjJ7FgzWEy4SNXxV
Ftt9U1IA34xF6oRk0z41e6LGSEVrfYN4T5b+l4Oak+Z8CMrna3KU/aDO0Xl5E1S8
wI0Sm3/arV3AFNfe23cK1l1zj+2HecSc/bA8FzuAd7i19j8jxGAjLrwER9EyNQDu
WKa9yygEMuV0pE6wlxmi7IZsWzO0p5gIIGFoRijf5hoHDd+ia75BHqnFk/SLJlNn
guGmfGXjfHK9tSkHQdNgvSse5dmzu9OUfISZ5BaFNexvBhTFmRTB7uJTyuS3Iobt
q0a5eQ/RWa7D+ubwiDcOqhTu74D5J3PATelJMB0fI4gwDYN9pkA8t6m7JTcVtlOG
dpAsZR8Ol07Dtsf5wHIc6rR5oek3vA3nVKRyRQduQ/ZLkrZgQjmev8e/elbH1VvC
PTFvwZS/OD11IJUnwZjai37FXbm5XFWR4+GDd6YkMHOyRlYOqj5t5MYYyTDrDeFH
pJYuAdv5QC3J8Id7D/elGCshY8UGXFm/oTug/DbWa4cIydFTlD3u9YbGtjF566If
3X+iE2o3QXUnyF0OhwMgXGLt9OQfooW+lTZ7LjMLT/rJxdIm/0DDFNxD3OlQeeK3
k7swc7K3DEcYnzPQ/q4RVfQ6U3Lrat/a39R7P/VBK31JNV0Y5m7zsGyqtMrV73Fk
jpeG3Y706TMjOW3UnBtAK6q0MuH5A10oOHGucLjXH23geNhErxg194K1nP0+T28/
A9J6+pd+aRa7pQjf+uSf/2TG6cNXff5aoh2f26nlGn1srHqQDim4BERpCp0eRjLV
Jv/Y/F0qTChAuWixjYzP5Wwn4PWF+shL0Xqw8NoUjeaLzgxzMw9NccbAUJ3NIB+2
mVtnWcvHJPZgXe0+FgvJcuucUsbrkX+rd3IJ7+pzlhXs1xn9pomJ9vjuCL6EZP29
dm2kwMNjOF8nqel7irivpENU4zsqui4NSaIMX6eKtcCC4fPgeVAFKjVvcM1nw70s
6kOKzm0SUqKMfaG0iWZH8RMiGgg3jTBHRFYjEI0LUHCcdnMQUucxgU6XtzF+UhIe
LegUlHaVgumYJBC68x1b3Mo2OV2Vzm7p3upao7UwUF662VgclCUVnoWUYYDwCAJS
JTLEFLKDR1y8QYdJ5vGpcK1jYGnivOpx9yufLEV/L7hXXJ+TxmSD8pjMazYAislK
8De2AUH3KwmBNLKyURRNW2AsXIUXkT37jfpAI5L4swCJ81kBc+ZcBFPb7vsoUgA9
bn6pK/l8CGswvRuiSHjt+oncwbkrrNO5CbyFNK0u/0+8Q9XSSmDhPixhRSG5HZrg
tgmXJsO6Y4heNjlCVXPtMVEif8iQmX0mL+b+NUipZ8WHXVTOEY+HJuDCt9Cjt6tf
634wbL+kLfMf5DW3KXb1iU4RMhkGW2lA49LymDZ7AAkCFAOfWk2FN/MKoTqkLTtn
8VlLkkCMtKFwrITqTfo3MfJF0uJ+nyIeApiimUoU0iV7Lr+CSiDUtyYBdzhV4RO5
mMM6BqYqxHA4oMU0eItsIauGrWxTrQsel27FGMJd6VGdtecB21CxEJVJC5BIxx0R
h2ig6rh/N4MZJDdjYYFk1PXdH4iLZqZWAsBGVfXP1fG8Aj3RAPiqmnq8zglPzKkj
thhZQ8qSrYhoNM7qU9SuVkB/26ZHp8kMknbaJQ1sHErfmaSveryKe5vkxAwXgeBz
51UMviEI56BvJktuV3My5El6ebuKysA+5Q/sEuaq/dGQv2ps2+j1C8Kp4hlhXd4/
IIrrUQ9Z/idj0UQsDrZvHgXJgXspFy2m5aBHaiAWGeKmRv8rsXi12AFnxJzl9Tuu
VslFuU0nvXM8XuynPwBcV6kf2y1dtrwuak1ZqfCyfIvC7Ropmgo02QFf4lWWgdUg
QZyYpbYstBiESLXxJOpag1TQb9/cXIuewQ6xM7YwJNwz8jgKVuXnuKDlxkNuWEct
hthK+TxWrljXzZs+36Z3o2T1vXmKRuQsbU7cdB00OBUAj6aJONQnDUqGlg94fwEO
IubjnbryQFrIybrHs1TYynFbNmtUuHfDC4U2NarTSxOY3Jxp2gwO4PPfzWFU/Z/O
+Eu0VaY7NxLvIAzb2C0XM0/UkVOe5L6ZE09pDIpDg7iuYtChKVg+Xbpw+2ERhKEk
QA+Eu60QOgSsLtC2tITgS9LN/eSlX/Tfc6hwlO8ixFGfqSLLhPG6CVExDf92WuBQ
8+NDsMJGkjBARHVWi19T0CEEuxIhajNt40oLLptCrVO6KRfqazmxw6DO02uDOlpf
odW2hmKOCq7sM+AvsIL1shK/nL5ZEfaJARQANyrjNCQoBlcBf3/ZNCXmlmJrlxxV
XSmA3XSj59Y+6U8IBy8WmuSfBlvGi6j7F792T/3h1r2mw5lrh1Axlvnq+2Carur6
c4WTjXs4lHN1KcZ0TqEgC3dCt7D6QXxSzkp1kNc8NaMV1elu8eia20kv6vOs7XKY
TahgzNTu5w3w8S9vvQ6x/thE16y3pPaO3mZ/V6HeHuX/cirpUrZCIVfiMigRaWnq
98uC99scueER/Rg8iJg6tRIarynkG0SRW2VdK1ylkYUgu9di6Ce51/0WeP/rILpR
YwhWqLzcqNqTwHokVkxhUTLpcIVFXGSRftWkalqZFKsNKeQFACfKYLC+Y52mANxF
AkXmCMLYEZv0dAhXbAN0McIY1UCw7sBuKXhWTQpCr1e4MhS5vOWV1zVVsDSc9jfC
vN0kPTht3mb0rhuuCLkIFZc92gID12vaOpXTkO+VG8HWsE/UbrjXc5mVVLIRsS01
FHWQBQeZTC9435sOYialXEORHT8eqAMTNTtfkg2xF8p9/6Kyh9Da1Jgmb02N/Z1v
Oi3UVBMKxRm4oY3IsiWEGeCW3TZY6hGEwva9dAk4LY9iM7VnhfqqR6LUSAlZM1/L
GTXyFZgSbNKA/r8KHzSR35XN8zLBNmOHuVsU6VoBO1S0SGj12gVMWmdMcmCZUp5N
wYQ3nTI8epk2VqOyFy63m2MLywfvLn6uP+L7qCpvgDujTWnb/iLNpJN1lncdx1Zg
lLA8q7lFSnihFiB+jAZaaHiaWBu6gNdnDdIycXmncgKWOGN14/8TPvUCoReKevbw
PxkZYt6Jej5ca1Ony8tBDGiZa+80yxAS+DtEM6IACoaNuDnHy2qagRTim3RbbHJd
HwHC+3zdOJOhPMe+jQROlUZitHzw1cB/slSOf9DhDy6xM4FBk3ytpBM3vRlweTna
hW6Mj5yIanrFt46YsWACUwLFEHf7Vaa1QgQ80w7EvIyWPEcJYxP11jryfw0eAwzu
HL1+jJECQBD/KkAY3N8IU/06c/C3bkypErWzPF3s1J7FsjEoguCkj9jrcVi9QZwX
7eRpfd9IN4hKjn4bTkoeSQbDK/9b2/S3FnkYUTV3aTPWK70t2neQXdFVTEW6jBNd
0WZj2v/cuOKjfpA3+PtczJdfm+loPJty7Dy/FRkyxfGaVzThTF1WJ5nyjoKC2ecb
HsMEgUeQL4R8J1Em/Si07OEbKU28ZBMCkSgUMMT+wKMQvhOuulOLQpXEDfM/sfLT
xN1x5FUt/FEsi1zB1jwB8PLty75ZLn3NQZZJUAaJyK8cGLLfI+ZxQP+9oBbLzq1p
Rh7RNz824yApOYNWGvHIM1yFxAvUQ44BXS/10MSC0eycAguVMheH0+jM3NKq3+Cc
hB03WXlMc2Y7sKir9Lt2lKGKTHI+USm29fKTPdU+CyktFUktTZoCPGu2AGzVWTPu
Kmd7wixQoPufGxZ3tKEcv2qT+WzvH+s9KFA9BWMKtxHeMdVAduG3UXSZZ49fw1NR
W5Z9QaYTcEeVaJDmCtDsI+HE2XChY3AtzfXimxOemIeK4Nf3Zlml/vz+QYF8hJeu
W1R6BJhJxXw7+b/K9r+ybs4/dXFqlh4rNzFAS17Vg2rx1jXDg6T+NKVjk8SoqT02
I2B7nBsOBxhj46sujxSwtJLpa5DMDPkKrcYnV0QXPgyunN7wh68d9yvU2c2b8OH0
pc90wY/QnUVcULWzwfkiBJXZqmuCi0EIbP2855LFqvu93WzlOTLunbwwetJ3vJst
atuWZw2aQ60zb3o7FJCFmiIlBM6Y3Ia2Z+2W/2c+tWn7Mfk4C8utIGqaH87/7P0u
IRfTmm22k4iy3XAAy2z1Dp/gGP8v28oArpr8DSYCT/nLqznOwjaR6pGcw7c6RSxi
5dlPN/x4nh3tuxiXz2pEbzEp0TdSkKwyWs+D1Fbi0RHTR4/KJBc/UGsMLijEzPG8
pfob8IYYcRbNYqTb1zF62zWgMx4avDUfejvVIDietufir+ehCVDuKjXHJGjXpBS+
ehqukEro/v3kJ+qXuWi/0xE6Gv48rnmEg+j+rS98PB++bMUpgNNJIT7sW/aIbPef
VDy68OeBi3UIob1FEp6ckLgAp6eDdxsEFTsVQJ8a12G3MdVI2xiIe5kWDWOWPxHG
0L7mlz6bU2vIRQvh3uffcd+eClfogsr/vQm0tsu4N8X/2lRNnyISiT1588tz0RcK
ofzPL56rXf2U5SX1cQLCqjrhfjWMios1w5YZyUwP43KzKxYS55HhibEIj65DIjcK
1yaTPnMSHXSmxwbc2f8XU3FTbaXWL+/j3MiZgPi4w10GFaKJ+PlCteIb7mJRTfW9
JEs705P9PKGmbC+mU4WEvs7KhgfKCEGo4ihuX2RcwByQG4mJfYP1QgOoaMKOjqnH
/P3aFgaHb6+WYY8uGPuD/MdmDsZ+oO1w/Ksih4OxBf7pdoYQ5/JdsEfYt3V+teJF
hZVSTGdGpWlbKGOmdslqA2n6gN4k3+x9ul/QgY+TADoYcu1mDabmJXX0ZIkzFFR+
VOBcB7Nnzn4QNX3fiWlGryJKJ8/+rPvDMQ4A+1NzgCYxIxtsejbCh3LsWZvK8Uku
uhiBbilBEbW8nCv9lfgzmpM9nSU44XYrZLyBuQza4tnKexJst4R0IxQu1D/wbKPi
KGPDDkLz553b//jfzOlgjswXuqG+0km6zLubqat67W9jZPuuybYfHCiuHkNZ9zff
cXvcSz7sm0V5nVLMHTxWJQAx75PZck0GPehvchmx3L5cC/+3i19VXTHFYALwVgqu
19gSElPaVjZaMhsXwT1nscZROlzQOSAsf/RU4427pd5DOeFbhSNzCCpc+kzKHOnJ
iWF/BKsrCnO7ulpJwNhaCLjAcoCs3EfKwJzSjkZMAYhWd4bPKbNGPSXlFp49MEe4
wPdSjZr06Iwcl7/RqXRqxEfIxCkcf4FjUdvvpPEVoHXLeyI3uS7Wcb21vkGeC8cO
wkQc3Mq+B1+C6mHMlaSy2FDuLLkDX0hT9oENV+Ltb+waSZc86pRMK4lW6Ou1Oht1
AGvCh4LRoTEOvCIPLt3nIHiqvsf06ZgDm0b+Z6eH/zlt/PlD17dSR/vcwMgEyKw6
8aMQi6Ix96w+2PReTpo3coAFsFEXXlfpfjzsjp5hiE2mlME/WzVU6K9J9/WakqOo
xBNlgvloEQnzDBpip64cC99yeeS3Jg0ZsqlBjLUjJQe7Akx/c4VBKGZvMpKJj5Yk
p6dtCsgnBvIyBP5XcMJvAmiae1YtcdvUxaVjJcQTjdSoUDUcgS7CRRK/5+zKkMhk
zL5AS2VE0DOC55etW8cjI1oMobtY22G1WGsRSooVehqGth9XzLd/hB0PyY5UuAFb
u5c17drc7WM8DAJC/lMlE8P/rhVhVlyjnSg1WAPhOa56NzsSCEoyDOgWam3+2JLf
HyksEOtsxStb5ZJw+O1X7of6uECveWFbPZH6rb3/pBWS1mTKiynrBJvc/FUsku9f
jCFfNRRDxa1QxXhIEu2GgHIwivZAYYMSORA7GW2JNoW9fsdQpmfBqt/z68Tyyc+K
wSjlTSn6ZqgqzfpIhjlYx1ToPRGBinIK60Q+m4b/eHiifu11wliWC1cicvyqmORm
MwTK0kVeiENRBIf95Dz3ynuPE2f99EWsCwYMiOxbgDackOyR4y3ZkuRQEhpsgRsJ
jMjAqclVR05EME2+BV7JYlE/ZZ5NmSwPr+i3+5ZUejjeSiykVseW6chO+6720D6A
mk/qKyZNgbNoCr2xJ4qfhcveL9ZeZvPWl+LCp6rDCWLM+eg9KE3lGjUx1qt+okor
mCSWYT2gTD09CJJbRSlhSeEZxsUebRKEdSuc+jhPzXTmHus1tivBygIZACO9MHbt
3BFmMW5yjYchpJgJNheehSnWE+qQ6B2+eJDAvLxfzRAE9FuD0M3JQxzqoZlLnI9+
yQkhfExXUGSihr8bbXgqPTPtNSsRlscezbdTidpT7MOdVnVHxe7T/KZRFhtPCFW9
9FOlPdE7PXp6r1YBMNTpNACIZKDJJAnDLrNN9oKxW6QOtVu3Uu7E26FunS5/FXUM
d14dSgs5y3on70Nl/31PlNTX7hJ/S97dgbToEINIWR5N+wBkJ/rNLZ4KREM1dEHC
R+MJRwDjAE8SWopSyv9yKHSg5FzdLX2D4+t3/JcfNsnjsuNzfV7R/xN+AiP7/Q6r
BDZ25ZDZsG3b96yGTQ0FaTp+VSqldEtHbj+wCtsgkN7J+uu3xcS7m4S9DaVQLTNQ
L4Z/0llEaliiHZZfLGMbnhem2XEszE5ssHz10yzJ6ibPERWhNfrrqYQTytCE1+z+
A/ktmyXSRxrFbP0+f8FEZT9thiJ+jotZIwvwNzSZiDI7EKBdTa+w04Mu/djZLCB9
Wc/uMMmRR8ToqC/SwxD3JAiwM/qU8CZBetkq7xKSfcW7A8SncFTUGBv3Yce/srqv
QU/6M+bou8XmNs+Cub+7AW9lw9EeOiPF8K5e9EoTkQh8lGvWgzzCwbjaW5iD1N1T
RLJelLkNLlApVB69jxy3H5Y0sgCd5GkhGOSTGgmHNLC2U5ThRhzZm0kxtkBdr5UJ
kLozugkGCWRkQLQ3ShwsA4wTcdWsxyHc+xLdIYIvaB0agbOk97jyOk92x37RQ05T
yda/IZuFpc+zE4pDuJTYeFwTfAOP1EDy+G5hbN8amMwo01nERiAftzPjJG3XQWj0
XnXyiHP4Acwk455HrYpZXY+lprqjJAzLM2aMYq5zM+TTb5q4tfUXACtc/t/reKGd
CHk/hF+Jbo8x73yZ+rDAMUpGs4NtOPXdZwNEl8cKxCPXX9mqpAND04PS2E28/WXI
1yZNhDMtN1/U9oD65LeTtbWvrg4ic/wg7aZ3P+drF+KELdk8n5SWE7hZBUR+VHzD
ExMYfZyBAGVJiW12et4kMR6TIhS9bYAEQKZY87ndRMcspWOOfcXA0bxrpbOhrNx+
/pCOj+0FRh/pSx+pzOw/bDxMX1SKDKxamAxEIrkShW3n9aQJgMJ7Fy71ylyHAJB3
Xidgwuer/yEeit+1WbzqH3MWrmuN9oUxF4lssSNV/4RhXXdzzqW2vfXZRWkSg+Ra
JAB25aRGWY3otOAu5QhvEP06PDMDrCTBebDoEXLM28eDeS51wukCIAdr45aXSqi+
I3oysrFpoW4E+yw/tLSAH1fxXab7dibs7b9cRPfUE8lvDDgdgdJNRSrG5JSORXgk
5Siy9/U58lqNH35/Bx+iyqTizLVV4JktorxmuLiBBoeaHPPu9tbpPghqGB88gjrW
bL4cZ7MxVxR5ti/nDvNLghXa7Ffpfyeo6x71jGaYJrUG2IJZHODeDBD46XYdHmO0
zPUPLar/9IxorI4egdxJ2B3jFkMX82YDvJ+X38Jh7aifiz4hbss6HxQyq6OtD1o9
Gyd4n6nIZR6pY3iFGVmXOnFjHnZXeec+134nFc5gZZv5206fNwBnA1BSpFZGfVdb
8FBHGmUGRNv93rwblr8G7ZaeJXIjt2T1E31Q4v7ToYOLmFPDVlu2lWzrFQlrzkcC
07dlblyqHNXBiuPdc8fQOtUgVR9aMlWy8e1VYhslazE1qJEgQ3hRSDqf8MBp1jBw
+foORhV69l2/9eLXUGpHCgTl/xPMERbqPAilc75LXjrPiRKgAxjHiVtToCywXFNo
KUwh2UUFdq50tfapnVIs4eipYCogqM8XfhLcefAXixJKQj5OYohe/doZQvpGJg0C
LRDFpmLBcD/1UGV3tIa2EMfTYJ4RZ5WGXH9iFHoEb9Pz3UbhIO0Ib8jbCKzj+dUO
muvmT8Eo1ax0p4kUua/fEeREYiiN3L1+R/9r60mkvtRvW25CQMMdBXjipnxZETlO
dRZHZBSroBCSPe6UojdrRyBCFNJ9jt8agClaPqAVOrb4xQXBGeQepG75xTILFZD2
EkF1OLHGye9WZj7Ku5SpOD3btVAPQ9b9cNqF6PWk5k36ZGsznZquI86qP00U1fWl
glHdiNUbHkVtjJgrNMy1VYgScCYPL6fqaPmv6IDUYExut7V7iyIVe112mERU0PzP
m6tah4qWTrH6WzzioNlUg1S9Fl7BkY6INmhiOySnfN+cqmevTEqyJ4SrcKK9u7ng
1a+rQSxdznSHCvjBhxbN3yvTtAcA+jgqk23OF7y+EEWaykYuX7UuidhD6MVrWzyT
CUCl/61eKGKBJ+1w5j2yHLg+JV+Gdk6zsgO1SzxnFZpINx2lyMHR5L0qgjQrHq6s
bByLMN3+v7Rw623M1vcdXepEYi9kBBio0f02TmxmVLVsFX/W6A9U78mKiei6BnH8
SeC5RzZQA88hfJUPLgL9mxdCwTtyRm1qkymxoyk6rY84rwxwurhTqX9Uv6vj6X+9
6AiL9773bvdqC9cE2Aw6Am+oPX3kJhcpuu8nsmk3ZA7DzrIYQfF5ZE4i/7mZcvwU
2YVEbQS0ZUqOCl/ku14dSLdEg2E4ec3hlCg8znWkB6vkVVDu7rBk2yO/EWJNQF/c
81ttsDGmVxSXtvmdFG/9slIY2y+b7TECMmtwnc5BpZCasDKwHwSVCDzBrZskwfcH
gaY6jRir2Zt2IkQYW9H4lCpI2Eo8xDrGXXsOrh2GAHBYQWLTgKC0C962YiN07Bbf
5N+kRYmZUg32pOAkJaWtklX5MQrdckK2fLoRtGem+J6DL8L8FAovzWZw7iL8kkSQ
rV5ihnEjTjf0IRrKIATyQwDtsCkRKY6Zb9TwuDPBVKcL+TYN5W6gl1PWpE39hzE7
c0RwD4i2Tz3CgC5Wvcei1QgoCdsqF51RLhOChNYzwhdcPDNbt0+NvowmkY+pmHe2
7FdaVK9CzdATX8sCkRwFm9hyybPXYvzyiMa5ddf45CjXdTC+W3qlBrVA/d7CdUCk
a6QACVji30/iMd86Hcb09kv5iAQ72V1rkyWiUd2r6T18GVTbTsvsNL8yieFawq6n
3zGYNFGiRlIbFieLaYPN+I4OdCqMkmeRcMzCkz5Hi6DIXKdL5y4ewjNf4Ry6H7lM
/GPZcdGiteoYWB4e5Fy/su/DBBqHkJ1YwSj5ePR71zs9DOsVdf2VjmUk+o6y8q49
MHlnwW3ZL4OQMV0FG0kzYvTNHtc3oR/schsoMQMdfmQryRJFwC1Uggq3xhvMXgLs
pBnfM59yCmVRD1ZruuIgerP1R53cSrnByY4sMp+VW4koKavZiu6yJ2UXUpuCZEeF
RZlU5XBfJDwKt/7oI7RI3u6F/TuPCQ8YSO0JHr5skysvbrtS+UzYvWf96QsiPnRr
/fn8T12rYhfC66Fw5zZpoQshNO1E+z7opnIyaERUdZYd+DJznACyPeBsCDJJs0Q8
hwP4QVf9SehlznjhDIXpzZEAF1df1FHv3y7Brazja5vZ1SySxZca726u9wtD0CQx
NDzjzW8K7LNtdctWxRMVN+F/yzhshsSErSjkfxaCv4Kxh48oSdolRug0MB2fmzWB
tw1UXTsiUj83m+HQKjtIe9Kr/9udRF24MqU9H3scbOZeyZhbIrIgxzEliOPlLQZ7
LIJKtWw5BIA3j4QvPyF144ZFkqwQLlGL9Vqdcc6LglfHipjGDLSt+/wOwFtsTnq2
iRMsEnG9rAf8BA7A5LIRxRGnV5jMUSoTWY5zI/71kCVrltv3lIIC9XZCspQ8RpJ8
/WZo1ab0l0teZE0kIY1P2DEFUjukxPpZ/4C44qEdbFnc565Sw0sjUzrRyBhrV1r0
zdSrgS5NNpf+7WTcmYTJjtsQ7xDr8ZnPk5YpCSu4NdojqMsget1a1B9HdO4ad7mz
gIrHMQIVTm4ZLAeswZN/Z0kKy35XgOV7Shx9efI7D9ycrE+Ozlk9AL8ZURhq1Txw
xdeqZSIRMhL3osBb4/nAjqZNljXORxecK++QVEsCw7pgCP/x9J92mfMfMOYSStf7
4roRhMgmKGhpf32B5U8gxVxz9so0uJFKnXn0vG9D5/460PhFXtCqqrAlb97+Fyq8
jVrSQDLw2PEsjlB507tCg2R/o/gzBGCl2/+wzkgMKVvIu4zGxCGvPtNkWa5G80/j
bInFdX4lDOdG/iksJAgYrSyqgITc6m71R4D+u45fSIDY0/0Uve8Be6umN02zcoEg
9tNeAQ2wS/MPEu3gkOTObFDaypb1QETdtlPnjSMok46GfI3wsCDOjN+5XVV8x0Ll
17kfOv7wKuAzQPYSwGi8ZFfT6GniC0f3NnH3hAbwciAZJKmyc4iVijdfkiJb1woN
I+TUPL8RB495ZoG+4+B3hze84xZKtoVVcu2Fx7h9oW8frdRl+2GMfPR+IGXgJkSj
IMOQ+B1m1oJR56aOzwI4A3y5gkKNRqhyPEoT+VK9CcYnaacZVA9cA2iamzQFTJs7
BG0ww2+SsDrT4f0As+0FF0FeV+ADzfQFPbwiblFG/JmBlI4j4H7SWdrWYDH2XtyZ
3G24EnvOXpIQETJiOLmOHLS5Xn+E/9SmZfVr3IusQOiamEE/H324IFK/QLl1Ur1g
frB/CbtCNhvvYjWYhG6xPt8vGkh/OUvyw3wSkZihPjW1EGNf3XsSr2pwk/QpQEVB
K+O3apY6qlUWVnfOKa54Ul9bO9F64tt5/hjKqemXnmjmS/1643G0FyzEA7VrfRmJ
qqtLrhXhgdHFM1hDtNhNO2wUDmz4BjODTkqf3glO13stNiudXjTC15G/RppIRMx9
NUrxsGpfzXws5mz+R9oRgywcFKdwDgDum2sJSgjk7b6+L3nhZDX1GQIQ5s7SDlgW
4S1ijEol7KCg6YyvJIisIB0R7lM28Mnf7IzVjNIhIGw858hecsJz1wwLGA+fpXEY
DxQ2A3WvWMI9d/ahE1gP+WOI/HEGGS2upEJTLwxAyH+YZWD54WzILdYOegV7gNRe
W4DLFqCBYt37oAjtErIR7EgWe3Ix9u6BhhioJ2nK5nRM2MvrtVmPsByXaQM5pOre
k+GTfTlQDY7wAk1t4td69jmstcZT/7tYGHYfEv+yrhEJxOyKl+EUFkyiR6zmBSVf
ppWmAa+c4QrYDRy42V90R0zt6ZChsIkfUhcdR81eQMTyjECmUrlb3/5+2cqw/aXz
6+4vij4zFOkJSYWAEPR6eXHhI6zcG3ulgahIbROcOT66wAJiZ9ErXNihZrRz4jca
eGZpSNT2o/kGurBO0WBWhH68CsW0mbG18+80/MtoYJmwXR5+6Z/XanQTgDHYFBmc
bP2Sib2iiekVJfp027Pzl+e1oP/rxc5UJiOJJ6fwW2DjMg1J/vhkPZ2Uyw06LZdE
KGwqIqKeNB1P+VLUgfCwGGJkfo5vkzRRpetRf8zZ2HO3wh8T3oOpbB5NtJdFqviF
j3iD6E5E/IwqDAi0etVksY6MkvgNk2largHjvvOUAnmdpNtQ77Fl7wBvKO1yTkwC
3lyTIFR8R6eWeiRwbQtxabr2FS0cd4Cq8vdBEVRZTf/vNcug5dzUTfD5aLrE8li2
S7cFnVWrd3wxABrPyRMOzHw5uIrPiyRLfDnOSRhyBokKHd7YRAFzwXsqQhgpTE6n
wl1gBFK4iMvLzT8FQcbXqSNaWGuktLdo3QToPUcMwC570X90WrPInK/BQcrrq1Hg
MoNZaM/8PlO1hND4xiwhOz9SWnubcIZDfc7FDC0tRHYELp+4T8m/dqXkoC8Azj8r
a2ipbtLD2WqYIckRvbeJ5J9Tmp+qML3Ju1qi8RtVWmqI43+yz2h1hgXBe7WyxiI3
z9hJCoaDl4iqrfEDCFITbqoSMdoZDiEgmJKFSRo6Ls96j9xbSb8L8c8APLn052Z+
XpZrdfw/6TRuMY5qtQ77M6IBSUfjA11nQH6TZotZeWVtOBGkAJ8jYueWyVZOwcO+
bjbzzz/vivEiC64JGOSehN7YSZyIyCWmOuvDxLrA3FkKRebzlny5qJB/3WF9KeXe
3GXAVg+/LTmb4Bp7Q9QrReaY6UkaoBn/2ENb/G8964PyEAloALvtFQK9gUq7qNna
dsYjEJTKIJViE6h3ZyQ2VJfH0TR0uzG9RuoIgt/utjkdg0qkTor1sg2mIqxKJTcK
2SLo/KJpDGmVyjEOrNftI2z4PYGWag3qKQ4shk5CDr1gpxg2hZ8HBtZhbrJRrgy3
EJH1sA2CQyFRPwvItEMwG6ZaoZAQiLMGKOP2XpGcWHkKcF3HQx376WJllFBkz0/F
zCQZbW986SZ4IO5g3Qn4FLQoQZt/imfrW69aZX2Fd7a3JDN3ytg5BH2PYS8ckt1n
7yM4+Dfz/0B8pJUZxHYH+DwBwX0O/0Iv6HyeU88VuNhUvPZPeCABQCKf6Ap9Oc42
7Q/fymK5Mg/yxZOjB0w+NIccJL3FxocpXAANwinRMPpi4EgXcH2XGe/7dnZIs9TM
xBTcZtvoWXXHuHUyouKMF8SKXRvOu3GNzlTGWuwnN4R9aVYaE3iVED9r/UUtTlvO
K5vbNI/5NmxYKH35ZX/2VlqrdmYw6RkYZ6PAtg+McjKYSR5XIrhbE2zRjbDgT1Jl
LY6nCp+OmP99dlpArJsA7Rf5F4jEkXrPGUexmQdS+N6yoFJe69FhWyHw1i7SDZGw
Zqvl7KdcElGblcZgn5ObmpHwlP5YSDvyEx8nRJppRpCWer4Eoj9PqNK9DImGkIZx
PprnYJQi/dAVkGisYk2tta1VaAvJBHtsKnhnlzF0uw5UXNO3HQFptj1jsHYzDW4m
EKpnhKheoOY9DNC2XwjGEljzAl4NVnMfG+fx+w85toaXQKeCRmNC+F8OoloLcUwV
DbU91sEiYRV1iLDUOlXRovZy/L2b3yjpOCWbjguxrRPqY+KsL3lYz7NlNUpBePRj
HJTCKeI2Yw52hgM9WtBtvNqmoAVaNx5Efz06Byuc0icMhmeTaeO/R2JBWkIv3j3s
w6Rc3iw7ZRH8abFbJX0AEvZ9z3aH7Ny95RyPm3IG6RN7j/++HbAr9UhQrSyzoi04
foHUlW1HCgZi7Amuv9JLk6ur2RZcdxfMegkoz6aCZ0zM9wtnx/outovJSoUwDBsA
n9WK9ysAPj6tafFNI097FwIoEfjfCMFgS8Eh7btRbqe6DeEPnB+b0ZQGFWEyDGtQ
qzNU3Z5YYixEAdGKHx0RALRGooWDuyzWWuwaw0uRyNF9OWMkRgXtlCBCj8A1MHBO
CUMh4c6acTyikKaT0KwDAvh8KSL+MaQfdWw5EE+fEG4GGPTjpIHJT1RDkZZJXeGg
QsJe9e3eJpHKE+k32anjuhJvARiTX3M/zgU3gHeHOFpwVlt+DPRMD8QZWfGyguJq
RDnGEwN8IcLAmZUn8/PcU7NV7OCy6OXuZe9PyUAVae/qwlgy301p0DSpFlUuSPgR
wEO2dyfNB/lBu9jOXp+XU/7I5X4zDy+ZFUNoryNi4EOlKjcSThhR3U23A2Ei0AYw
eQD5RPF/rYULldGCVAupNM8vCmGWkCYmFV0lqT2AmH34iG5DMPXKi6YI48OCsJeA
bueOxNHYUoHj0qqQDiNCjnJjTv+BqBPOi2t2zMmask2PnM4BBX8RAIMU7Msb0QtF
VgHC1TQTZxO0A3Y/g/Oi1OdLgvBiCIAfCnhEaiTxxj7qCKYY3BJ+RUVC0OA4YJYk
wByQtzZKRvrKbeHfInOJaBleVYoMp29oBbsh45lj+39KcIanZlXj0okj9Xmcwr3v
aXPV+RkeRqViuYG13G6hvnIRHd2g0d/TII8cgBB50Tcp62b669OwUEahXTgGdFng
6S0G1G/qB01MA625VQiki/ELg+FGOEjLjAi7+KraxlP97GhV94UxpTMZIgcLo5Vd
PUIMMsHhsZP+s5B9XADO/t6TmzBZrnVljLmGFPCw342GdtzDgYc2R3roFzt3NtXl
yPwFeVvxao094j25VfQ1fs+mgJP4vq929uGhR/OoF2HE7upGmXRtUdjR4YRZoqxY
bAu+4rjAU8bfe5GS7mZKFG+xRabpQYcez1NOb8qXSJFxFREC2fONeGxCrurH2QJG
Q9Tjs8zvr8AnFMWPrzB/rc+qp7xxlKeZ6CJcFW1GBtSAoyZBaycy9EcqLddRf/yZ
VwAnrJMGdd0vxmBqEmFIWRkjsJniD0ZeDxNjABz5p7p40jWfXdnS8SceBjciTkA9
jLMW8kspDmzyXsPO0x2hZ/U0Wdm1s3UNmebtB+ZN2fHLIj5gVLxa0x7hWvKydDPq
YZw+7P5sNSGXJDzwgfidBTqoy9cPmcib/Nce1UaqDJ78wP0zPz/+3Fh1CCCCLK1/
Oue1Negna+Q73HLxDc4pE8nNYGmZ8pBMRuKUcD5sAUBfXQHJ/h66EJ9/Ipst9EWy
gpH3AQ1wsnp78E06BMy05Pk+9kMXZXda2fOW+oTnlSKB1Oh2PONCsRzIZbhAuOIw
RpugLaUr7455Crmf3zJRIks5UAFjDLG50I+2oEnuCb7qkbvOcmAv4XyJj0Cgbs4C
5KnCBulDuWhfAeHK45hIte/a5EP+Dp7ZkFE8t0D4xc5E9f5jMIqcwIcWidoXygNJ
dkNMnemLD7taqZ0vY9UkJ/Y/UfQcP49H9sS/OgDCg0rCfS65wcuB+NANYZrtpRtB
+oTASryRIS01egK64308HLcBcv62rANGQv4LYfNUH0v2FnKWBwq/D1Dmea7o+jxb
dAlV42EfTeSzCKiZpiFXFnUATizj1TrjZYmhJpnJvPykWYKQRN1rKpdoVucq353H
uwV0leUkpwTWCa5AghUNmsVbPkQOz8QqPdYF83iPp8EA6xLCyyoomI8QmwexiKDA
VA0ci9HGMXsbVz1HIcKTPFdKYnaqeC+JE03ryhJlU/5yCcIAu/Cdvn/u+mGKVoy7
Kjquc/+/vORYqaWhPR7t7c81znMy0Iuby9vfnReRlT5vL0Q6ALLjPjazwD/WV2HU
hAdk4ntEhOki41ynqxzjun+/RuQ+RPa9ESxj1ioyQ/Sd3Z6vgA0H8aOFuCpO1WtE
6Enw9uYTjuEDBedTt3lSs59u20ZWdDI0pNiIBsxF2C35n+QHvJLCnX15z3HoqOVS
H3w9tohcQCu2yGBYyKAZahxG0CcUo2vlkWKrpys8A/pS9N5tujxbJH0V1RT+Ozyz
YX/VfHrpHRFS8GzBHvhGGvNAViq2ac+VIAa+AxyOmljLLaNZvB/S3a85ukZH7DEw
DSFkZ+hdIgCtqWwY9TXaQ0P6/4+Rs5KDTD4d54cC17y8v7lnIjed8yYbOFVPXL8W
Bmb6YMaLpA4F9vyGC2Eu6Pz8Af5a1q/UX5dooCs/OrO/JDp0LXWXjcesULUmFOXa
UZPFd3MOblxTRCdscP8jbBEANz95KQjZmv4XzWNvypRlvIjUBrirGHH/+aI5nLDB
Mg7y0/EzunSWOOUPKMxsqoTN1XSjylA0A3CWPE2LAzBE6I4iQffoaLf8wQ9Gx2HF
KyM/53aOdKzVLTfBwdDZ5q3dvEX71JGGB9u9m6N2juJxdu7jJXE+OpMsDxXVL2WJ
wfK4SoEPmcHACLYiRN+Y+twTzLcurtEdHnOthgSfeAZnm8naprZpH8HOgjEoQ5wM
v0N0fCnWxU4pX0tEs6byw14XhKEf7OcfR3yvbTxulKUH+GnQAijvLR3ucSLfGasR
AsPfEI6pOsLk0VhlXO9zWROkfSp3kX6o+dtMjwASbGSHYBdSVVzQw7dsv+PAT7Lf
mZ6nGhOFLczuewUkh4fsyCLihjxDzhIQgmLQRi3iL+aZm8ML2m2oCDPrjm5Sc5/v
+hnteLKl80ZLn+7V+gkBqBiB4xf6nYAvKRMG5R2f5D5bxEF9Zx9L3ufDUlhH96ck
vh0k8PVUkEFNpKLq+szec3yQNBqiEZrDNeQpuAWpnGcbTaDl8mcH1+fPGJiVa+Ik
tYaPMc7g53FOJJWErtE+7zxMtTO9xN4SMmHfxM4t1zU0sGIiNDxSCw5WqsJWy/k4
lBHEUU1eVprmDS+SYQ/vn+BMM5/qNJqMbifgIWYMZTpnVMYWs5q1OV8TkGfSUrbu
HV6/nx1WquMdqwM6T24LlXfDqxLU8x6h2Tv7eh5iij29OIG9UPH8+af5VNmMmXHx
zrH3GVNHZ7HJs/fKBf5GKbwUlmFEcaACGKeVXQf0C//rNQAAcQ9lAenhPN+ZOJGJ
L+3a+DWDVtamMMeLGr7Supd1iIX2LdeOe+U9j7H7pb3fWD83/un87VfnOxq5cLSx
0gfK5V/aX2FCi36nbns4so0CIcF4wriojQIiyyVI4Xcf+utTEIm9S05obD9D5+Y6
f0U+WEgsuvKrJr4V9kbcBsLk8kE+1sUlFLS86SVGNuzlLBEpJyk0qL0XGVFf4RbI
UkO+mbuGs+t2zOSBGm0Pp2WqHoDLQmZM+UwdTP+/eHsoTN/9o8YL39stCuEAiJGv
AcCQEeUNaZh36P7lDu/D1RIyV+LDjolYeuR7RRl0VxcpNLU6FzYvhj5sR9/QFF8a
DtXL7vowrE1IdlBkR/xoc6AFbpNPcyiOI9IMIoYwbSBiF9lzHOUxs3V//u6SuQ72
2li4lA2P2CpI2dcLCnsjcznzVcYk2nPuo3i/wTEZgtGzPwcfccYCkWVpF7JSwSYw
6pDAIBpo+1xaMbk+BBf2q/LOC/IDHqNDwtyK51B7uU/59lqj4gLh82SR5eHhqAYD
4/3mKDKuBYKgsmGiNY1qa3qXLygayGVeAWJUTtvZmjRnA3t5bmbCFoqjzBdJIrYt
Nyc81QodFucAH3mufHZREXBq7zrJeM0RPy1I8GgJqUD4XaFTRYIOj0HCWp8kG53+
qickTTIS3oIjk9+XSvdUkoGJWqF6QBA6d+FXbFkTJ01ai6ZaZ6t76nQnINh26ZHS
OLTxMMjyCv9oPh7GT408FQWuzzj7u+5dNf7ICRu5lHWjVd0jwn4/+vykZCo4s+dN
Spi30HEETMsk4s9JKvAhUGeug1WKd6Hw3Z78cmnDyXcGbfY7MgR+cRns/K5dcc8d
NGEcH8QpNa+C2nhzfJujEVGBHmUZIWbyQYPt+bXyaTAFqwL9zo/AqRTxjvSgSnlB
i7N7lrXCmcRtG4szCq0tn75+GyiQnLe7z2XQ1+SBBrQbAvI4J7frb3zcKPuQbX76
IU9PH9q7r6h5AMcaQhUYQY/EjjJWi2wfXcKsN1LCetHXCx0dbXPOtpJHghRJCWrB
hdyPfg3lgJEZU/OFyOkLv+fsI7nbInJBXlPbKQfCWQmCH57/vb9wC4CVT6ozQgUt
zLeueyHI6KNQgoUUgS2Mm2aZw/Af6IrwlR5r5MFSw9lEbtPbHLACg/dX0zFZf7oy
r0CXZRqn1Nuy7Fx6sGnKAgAAYU4jmEzp3J8mw7QZAu6ieMnafpTGDQVQ4th/06lf
KgO8IbuJQztZk6YvRRIn0VovKoWHdLuxoReqHFTQTZv3og1yrayYJiykZoJ0zEB1
4hJ9WbEOMhpmtH27cVumfZgZ0t16+fEA/FJ7Mo6xs5VmnKDmloZ+nZo1kmHyPgbD
Tn0cB/+wkp7QYXzxtjLes11t9XEnLVzzWs+rD8DYchBKKqePOQvcBaG537vaUc4h
9zOy+ACWtGMxlyIYIVGLYBAd4LvABiAtVF6J2b77mvl4OPlsw4Mlj991hWWYO81Q
0gm75FJjknKwNlPvzIUqsLvDS75P6s1Fkp+EA6qMXvHv4USuJlPMirDmtBSzCWXQ
1NVyNQsX0QsxwcVmfrA6sxkXeZSlS5gQmZH4MQvB8aa0jw8mtnlBfvnzSH2Faeer
eU094qf262JC6z+moKWfWas5V1YfhM2gI9facVNzt+vI3xdeXrZW8ITaLge4H8vs
rlxOS6kLJG6XNhrsMo/tmBIYj+3fxmX2oxja7fQUQIIXU1DO8mdW+NdEjmcDFLU5
GxT8PqCfkaXXD9SwUavq2ubXHAR+Vv4sG7Cul2Q46YNkDZ44DCwwWQ72cid5ksUU
yD6dsyMTtlmDiMQJhDmjXX5veJyXYVw5zLqLPdV+EYTAelEEpoOynX2jx4DochEn
X1B3UKT3LXG50dQIXT4bRLy01NjXYeWwUBhFXFJlvbBCfNhC9x1rGycai1lgjwtn
yppAp29w39HFFTd5PhwIuecBYVEU8crDpw/pTItieUeO+R5s0NLmmcXmkBz4dD7W
0GGXGjwkSkAb0XnDA3zn/e1HaJJ+jTj9LwWtF1Bbl9TtvHo2mYx3eLZE5SUCS5zq
x1jEUTEmcBlUTLzLUCDx3y3XmX1dVyp0P/jDg/nD1rzqt0wsxtqaGtGuD1+4sUYR
Qlmb86eNRACAhcKc65p2SlzdEuRVAwgu41VrCBqIo55dRgFsXTdEZf1rH5z/xvTD
ighnnWzkpVv92SeOOnoFoG5EqOUf7uj814Magsn8nTW9oKOMTyjtxQ8GDdvE+mrT
Hj/wZ3Hga0DO+/vxXhVGZznGa8isgAQW/W8Iww5jxm6brqqoOUQ5/SiCcOicHMRl
xBnS9M16p5ItiaN67GdOG2Sg9XSJE/2J3OtpqSQ9K6TW7LbvBaBV9whNjDz9Z5c/
DDFWu2/URbgahQNP0G+FkLEHwlCvzArjEXHhio/3CjU0HcrIeWu7jl7eqXkcDFIG
m0FZO+C67zt6YD0Ln+tGNqcDgHWapBbWzOgogS3CR1TQvgZqefHNC4NRIfDhsn/C
vHy2q+OAuQF75V/wpdlARFi0IRXDVI8sxwhu1VulnYkB4Z3mxthDHpJvrBr/3p7q
6xK/+lZYIh7+SnahHg8jHRjjmGt/KUwVP6NuRbHX5dNdlcyCQlhSFr+chg1N2iKU
1VYflIshZEPVvTZUs73HWB34AppElQfIVvQolAzZed9DcysM7ejPv23V+Xh7uJWq
nBRMhTXYxDTXZZBgDa5RHr2mRXXrOp8Jb4019VYr3+RhylfruzpBLl2cVRsKPKwd
Oog78In5FCgnBZCt2HC+Nn/hgMTFhexwjLoseb+1RnVBmkR1faFMj0tIg+M/52IC
ZYR9miP0CXqLFnM2SsS+/hUgcN6lhJgAc4oQqTE2XS6OhcfZGSCVkYDB/30hwLUZ
304wpVxBeTjxc2A29Fnn4Wifzwec+q9yWPQb6CTINuEC53cmQKYwjb3gcWIO8XPg
8PqkzjsDmBbUTCLja9R+y1ynnMZM7vzG/alYHSONTV1ykKkC4kqfwdvPsMLpZdHC
xToE9l/6hSd48N/kOWNJqERj8M9uv6ntQmewjFQ4RNuA90PIY4PTQ6aitcs/flyk
U/Q8fOX8oFwGJBh86FucqknbyUchcPI2HBx52bEqpXHbBBSzxgY1n/633PCrV93r
6MWAiT88gEQ42JRPurNs2Rd7ZR/iHDoyypf6KJ5OcnBg+4/h5w+W9F2labxINn7B
D8P3087w4HBnxSYg8/RNtjuUmcm5FxGGSGe5YFUdXVT8WOIOwY6qrU2rWL79RlCj
cAUWN2O+Pfcy9WZfkAYziJMxNJqOm9z6y1ncMx+Q9pTK1H/l567ZUra/iRyBtDMP
+ls6mGwJmsDR4aAkpLmA3oTmNKEeIEXuORfn/PWeTvha9w47SHQhkIXZXq2hqQGp
NuWwCXg5VBELiiJ0abUKQs4DCH7Bv1rtD86phUT4wMm+AkdpwHX7S1yZyXLZI0k/
GRc5ZlsyCuImvsMVAdvgKlrQSQi/w72I3rdrWYEDdQTjmcIlKftfGrCrfR0QQL7R
X6Xn5h2HTRS8Vc1+0CzGhzJykh/HnzM8A3iAL4OndWkJakqBIfT6rpeCjwmvD841
AbhlEU92zC+k2eJwwCjeCAjwSLFAX4ywxTfUvCWgvpPcvvqcTXIU+mGhLrRecuN0
YDBUtxLzQAkGz2doy9biD7B0hxK/pNZFFzWBOzAP0+EK+VRNrriZ7wLZo9hAgoGG
bPjlGzRIH3olV39oMaZsgWsI6LHYJd+0wkwxhJbukLZtFHFDETXFZI+FIciZrjqr
dQm9/boAXRX5WLwgbv9ZgQrbS3amklN0D76rQleVG2CVlF0qaSDMy7tHwaIXrBZz
N4r8HgpJuoHfq8adKHm4ewdfSNQ2XI385xc+YBA0p6O+TQBM0sMr5iNTDweVQ8LF
9n9Rnm6cC5O8lkcdeuWYunEY84pQaZ6hLrQ8aJKXX2eNJ12ylNVUXgNm2XoZRghm
j2ARESSU0V0l/h6UwzvcYS8JZ1c1t1gqiav/UWsTL3Of/25Z78z5uKi+Xi5CzzU9
owkd9gKLaEH1FAq7ZutZJfw17YXkxmuvZWVk3BKGp+yAvCqYbr1zrCScM5OapDhO
W4EtDN54nYDEfu/PxPSCikfqyHgUOF/yEuloCDoNN++TuFMD8lChSBHawsefqAKD
n/4EED1tZHoCNBvd0FBZb9JvlswfNbo6a9SmNaLc9332X1lomP77PiuLPjFGxrG0
FPPQUkmow62yez/0gt4TFCwj+1xJcblyFXQfOoYZfSGkW3TUADywgRWRXRWzILs6
DCZdwPfo0mPXVSKztVJ5t9bBBRErmZjvc7fcEtpQA8C9pgrXaeTppy7DjsbOOtZQ
6Q4PvOnftTGntjIy1Bu5P7X5MnMde/CFyQKTi7YoRXDA55/fFBe0ECr4pBvbDwvH
j8RGavD9fAWWkcarQrdiui0EmZBcjjMkD/etVo2dAhYP9S5GfFaOzg1uOCiDB6kR
/heezNrOX3yCLKwwb08aCFoyc2iL1iDiPZk6kVcJdO7Szae+Rx6tvheCsJNpqx0L
cRKPWiDEBV9rPf5Y7c8D8pFxI6FnMVOla0EH8RgvJfTqnElv7nLSC1Wgap3wHIr/
eMK+3pEAPRusk6gWxk6ZdcvxH/59YdzYcK7pgsDJT4ko8jgy/u4KVovaGuRdSprI
qdTEeB1IgyUEHPtm4mQ968ZM/sB5h1qfjE0EyBg0Uw2Nc2/X2vmw8leJFLC/GPde
4gPJD0bzUhECUttWeNdDwG85jDwY3GnGQhW+03XkW3WQovqRf1ymYWDMZ5TzZxr8
PpedxS1sdtPURaKUndjG513BasyuNX1ENcgU5f85FJGvf48I5+8h/aM3shj58Uf8
NPWRsJKjfgw2peWVO1FoVSCOfnHIMY+xKtUnjv7xav+MCfIwoid3FQ3BygirCsqt
bKR72eAqr8HkzqP58gZ1MWOqcMbbUfabkdBYClwwDJvwTfa53dAl9t929ECejqUo
DQGNChgNAL8Xo8/7qjCVXfLGHtHjp2UqQ92CLwF7DnAR3B3hjMR2C1PxInYLHD6q
SO+LvZ33+eHjd+Awx0Wqy+zWPJr8UL/pctrKOOhs380xEZ+PNRu864aBXCbK1Lui
/jTQR1hfpm3R2Gyngpw1RRiqbSFsxPDS8rZ108lG2wEiTZGWLFk0LLwnkl6jdMr2
3FRtRl+j0V3gHaorg2XQ/I3jFp2qozAhCHWabF1/PFMP/JZDWqbtjxRIJBXUx30g
roHPj2rghMaP+AWBdX6PVmBkpW1LLFC6HmTXiSnsBTLNdKDmylMzb0ToeK2hRX2w
hjT4wfVF7qDT1mVHaV+6FrizPevNro9P2h6qZtqapf6dOCe36StKHguE43ruDv8m
HCxcvtvMQ8/RjKki5TeXU2SdLqK6JnencBM2WRhGIRhOCYirVycwZ/VIqSH7T51Q
yZ12Yb3I+bfC8soAitqo3gp0XJkTwhgHp/Pam/mv+T5wEg5nCLpnKmJUZU8uoR+n
kGEE7NLbCdzEO8XzZ8GLmTpHrpXpjJdgMoerLXeq+6y4TQMiGQcD+OG98NM+zICh
C+K7F6Ql/cHsxFh+2y0ojMAjHxZNiIqIZ2JqzNC+DrTvVYo2IVPVA0hBRcIbVKKL
PPKB9A/2DO4irRR5qm4Mp2femiHuucBMzrufSPUulo0CbfLx22fbg7d15MUHm+Tt
Lcjrdyb+XaS5j5XqpYT35QQPRkTJtzJjttzZXFYJtIcqZJ6tuuyesbh1z7/ShgYD
bEOfGchLQSmgBdkJxXyp4KHud4rBaawRVr3HVFKi7EP2XPJppOAq8OcVsxXgcwGi
34kXdc/TpvjTqqaKkGx7ztgxpc6lOcWu0DDasdDkoZNE7wsbyNsj1GcffmYTZgrZ
RjOMyMRD+DzAW4aYstOoCn1JvFWSmWPQjv8BQOVdndl3NDz7wuyiLVir1xSrIuEh
B6ZV9cLpR9+/0Urt+nuM3wEResGkaMzxk0hcXr7yE5KF9I7KctLTnrZxQhoZpkQX
PPjm0nz1ZEmr4Z+wQzW2OwRUDbJGOrmJ0ofrfxfdSONWQ6P71NYOQLw6rvNLqj7T
+CINmcEaidTWu0Jf7TvOw/gjbAEvlYpPSMxQVQvzinf55ZSESq1WiBtNSAY7M2xq
nHtxVScXHCWE1Rsp12UOcwNszaV3tuf51gZUAI03fcyPA7QhSn4uKu7XvhXwLR+C
e2Mz1Z8Qgb4jLByBlCUwT+49UQoXqsYtx8+CMY1ju79qYrwqEPIWP8me+dphKPby
vKTbr0un9hUtrbaxP37Mi78sJtIk7ZMfUBtRrUUGfroiO6fxCFlIvxj3Zc0sHyzd
kxMWjk+PEkG3teeJjyhxL9Zy6EoB3sMepiYHKDfFzKGovnDruVQlOItaYvSzgMp9
VYytwC1qr5DvkoZOf8nv5uaDL36LnSXr8OrZpxuxiwTdg1aNjhDaTjcyEIkZmjoO
VOIF/S4g322ktjKOMluaytxeuCZo7vCirGAriyLY3LZCO9WdMvRK7IyCVz/TotCA
Xt2zK1v6YiHZT1WJsbphNEppG1x38uFgLNWA0hLGi9g7/ryY0KD7baJ5Y9up5cGM
cmGm6brXRQ71XkzBxLsFbbZijHWQqbyIERkvw50HfKIcvsFT/bUz7IlO0ZPiOn0h
UwlXX0qznRaCBo281cmG0w0nesZBskJHxOzKQrpZi0ic3V2UlSXU3+JhxHzHtblB
16orYW+lmOq5KPUdM+MYSB1Im4LOTHcRMeUKLY2xgReRmR7FjJeknlTUvIA85lxR
8zfCvZUvWIK+g4CU9VqOtUIIh4LwjpTU8YvltTR37BpMIKqLuXSLu+l72sJt85qU
qwc+J67QsVkE0BE7mXG8MAOsdEoMy0QWaPj0ZMkblpAfG/fyqmfd7QjeAYUdT+6v
u+h1+kKdwVNi8pGexjktjurRaAsF0VzqgSwYtP/kjdES0AIRpAUKPdJ5ALVfa2MP
4/dbVSufmec7bkzwHd30akR1NL89qfD8x6ia7YOWkTZzVsTDZmVXtD7DbADkjFsR
tG/g24xfN7Id3xKjFCHv6vT1hTGuOIQmmAnLzlfZVpEsEh7yFs/jTcW/xxVy5cup
Cc2rWDDZmWAMkJzsr00RtYxZscjmx33p36cMp1BZ99VDwYrgsAzF7d8I/lcj4QTN
TqQDsGTN+mBu6EcgsgSBdo+ntGEXvq1Eb52mXwLQnHDzM01iPJPXsqhywydUM6wc
YrkZ9wfBnM1vEEO49j3fUfeY2D0okG5vKxD1JHYkAGgbLY8V3I1uN47aUpA9CxWH
oUPICQd1ocXs3zKANOCM/glaH5o1VQ8TQcLwvBls55qTvQ97fMUoP/BdBRw9MSVi
nMhLfATXpeVnzZLUKTu9amQzkU3+HMUzuwp8JXkDJH+G3ugaDQJKEV/S5mtLeSC+
GzP/vKIRYt5V4cEJq5Xx1+SUfreTBOCULn/d8ZXZEbubPKBscpIZhLqYhDLFO5cA
0FbxmnKqj0iGwHhPM0V0slp1qAmm9BY/D7XmeGI4i0kTN1izEFRbiivhtl+GmhfR
XHCPEF1Ee5lzwb2Vf3OFcbdkPFB5JRIuEAVwXH6V+T4rWiWqlKCeIx+akaxtCRak
ooc8MTBrYXpLmzl1FfcvcnjcjA/PRNm/JhIq/grloKkMJerhNjTgGLvxc2+m6xjR
/lim+c/9zUqQX6wGhar3PoNv9dvPDT3CNffDvm5xtaSiVi6X0nn8sKUpcpUth4NK
faAmlDllKBxiwd5T3XdH9a+ynNx7SVi9L1FCRybSbdrC7bLFcp9vjEjF3Gb0xcYl
4J7C/KZ42oZxsy7pwQCKnXgLSkWnxj4x2JO8QYjjam7GdLftxPWHzVr09D1vCwUu
lDCqPBzqDJtpAC23KBoRuRj/fm6TUcDe3DTOx9OcrhthpEqT0QPMCjpmgGkgsQn3
P+qmVaszpYNYyNonjvwJqsFgJ1RrCDdd4uVvjirFgqOA8K+h94X8YJ0kKNBB03pt
Yw1Ja9ET43H6us1vQQ7vTg==
`pragma protect end_protected
