// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RlGROK3i4sKZZfnd1xNuKcijjDEFVzqV08W0YHAnshGqW3AhThkyz8ob7Vqd5W9+
avpkbzncVRcn1RPwznGJ7+FPbzyGTtAMbeoHrZkRthUO7MCem5PQjWPbDZCt8Gyr
ar58J4icszWSVpYyqbJbaItEFdVSAzwivD2e+qeJ544=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4960)
Fxpj/Lonu504cvTqYU59EpwQW4fNSz/4Rmc5CiRhGryg0rR1+7vBBnzDohtMqdNx
gQOECyUuc3uZeOC+eikGInlagEXJPfJpeD1pfZAg/K1NKcFFGDwZXea4RXyeU9cn
45k66cuaI66ScCk1TzGPr7lvIfxnLNj1Gh1owgXZ18ZCBAmpQ+nbKx1Vf9plXtIm
tmd+RRTOGlZVBqPoUfCUsjKnkV+DnhDQOk1Y4IwJYWrHFhDtILMTvFXF2/U1J2Zv
SywOfHba9KMXPxLi0SOx5+Tud/e2AfS73x7L4iTuJOH5MRCb41hwAeFxsvXiKfON
Y7qdXQ8h6jRW/nRZlAs3A5Xyp14y+Hm0tW5wHJUA6gQ88F45dxMgWqSEF4RSAkrf
aVMDnZlTavxoHmQKRD6/6DoIQpT1MVyOWMhoXRn0loUWUeWvKx1AtuIIuL4mG7Mg
A8lPstTVGmPBuVfyhQDiFhQcBA2MbES2I6vC4eqx+L0vt9sVlZRjUhNBboF5AxLR
rca0M+ZeubfPzEkvYrpRdRlBrAzdaALJ3KqY5junCgjmaCHvpt5ktLcMjTTExx4z
tYBp/xlzWIsejSTZO3/GqIZ3dkecvcV4U3B4X/s+ZBReI9uNoUjl47qLuE8FwSM1
QxcuxbYGzmoZIkvASm5dwt0+TQmArtvrRexWoEmHKikrIRZ90pVqJmonWV79pi2i
nvyZ3+12/AHZbbjqNd8f5MN/qbwzfSj+Q8oz2S6Sik8Cq7GLnIAbHcbPxeKE6TZM
aldm4aGofvoExy0sy7+a1OEX0t0wJiHBUgIUifoVO7Vod++OPUmFB95dkWuXYrkM
Lfof/Ml0CUhXWrmeV/D1MnhDE/icAzpHuJVdL8hr1llosAjMv8zHuQj3v2erZrCN
1E1dPFui21MTSktuGvgQw4K6aMHzB6wRmG/l1QqHo5StgrB5LLeBi1d2o9U+THC2
Ud8SfQEZVg+tTkPzK+sszdDB36kBn9zHArYX9r9NNuG4cF3HXeXXheH0R/jzA7Hc
xh1W+F20krnvk7VLVkF7KOGA9NnNqEkuK5byGSiNeKpECS81VrimsmBZBTcqU4BI
LsLrDcScREn6G63+A95g/8iaXv1SUnzTCLvpBIvrcXhQYiGV0Mt4MnhXufKdh0Ry
0FTyE1ZGXkSHL3ASUmlXO+LoUQ2fvT49444aw7p6iswVdcVbCC+O++4+Vqc1o3qv
hVWQN/5GTu1/jTuh+d1nFmg9Aop0xheyJAAxxCzCUid8Uw9q8IP23M/7iZvztLdg
pgfoV8neVWxqjFvPAVu+ZkDglyE7wgOOS/2jb4PuYKifekUdCX4W+nnnPNAgDQGH
o/LHc6QozEmU6R1KmolG7+yuz0InaXzLcvVOQrg1WJhwJwAjyiHQ+wHkgTsP1i1U
Ns3WqAwof8qL09bnqcrEFniYsORUx2e8IusAxQDmub36wnufotjocr4/QxI8jVHc
3sWzDegFLnCRxyHAu5dP1baDdlaIs7r6ARFhzMmd5yK+OMvvCzpu5xKY/uFg5KIq
ygqX+r5tg+gVpoIilnBzEI4uzEgrkI/LkwerPCQ9aGigjzIQyTPTWnhpFv4mkJs+
tdP8Ocg4/PAm/m1tg3+Qd1fV3bbwUVbng5gEhr9gVIUbP11AGaeo/XcoVgBeg+gB
ZFDoaFiSa6iXEuW/Hj1awm39V9jbkf5ktDK69WsOuSFxJYk1Ei76ruV+vWXrXb0H
rO/iobX2Xah+fq6exNI9Tz/I6H4IWQtd4iBFLoCE7MnRIhxl0X1O2Ftu1Ay6E+9N
MGoAEIywlR6qfBabyhsa4pR+n1mw26EycI9dz/IH458O8J4rjcl6mhiOJMZPBCwW
DzzjmZztCYADBYD1KFfUpW03ucXGD9FQqSa09BaX2ZHdNAu7jvFDDBj8S0pNVIY0
DXCWY21ke7EHMNgIv4SQySd0iJNE6lAuRgSm+3cIeI5ncHiX9dBNzIhvK5+d/d2A
AAdZDBPnI1Js162mtLGdtviq9WXKJwXVDW45Fsr/UdavqTpkDohBAvT4vQjKKVWi
gdWKk3OhsATGskrBgSu3sGr0nlPgrIjTu4iPJbQJVKH2PKjwllyEefwGNcSAqwg6
BA+JOqg+/a4f0heawA87k7JbtVJLLuq0+aDchN3vL6uuZVj9bXOHidOqqKqtJU5d
5puTo0hHl7YVXXYQY7Y9fvY8I+y4Ju8zVtVfITe4as11+r3YFu65cOUX9yjuhswP
h/ybVt4jpOam+RVQCreSX1bIUUlnLvlOEmLq7oKpADbRiIO0S0JHBmecoQZCo+Oy
gR99ZEFMTeHTIBSRwYK82KY4Un2G5GKkdOlsKLgAU6L/5VHL2ABDGHA31KqJAC91
TVX/EJPzAW0mPy2wGfcrkx1f5mfzcrv9wpCU3Id5D1UiMmBIe9arrcdzI8Epl+GO
EReQJifYIXM376WqvoitMJp9scvKU5ktDO1yUXMH+POsE8SE8OhK7eiK+B8gF6jv
tMOVv9uZHRkxW7wYeBugKN33kNBZ3E6WD+/xf4KEqJ+7ZYiDT743UYFuRxpi9HWn
45dlCwO05VMJNZEJNoASmyyF3z61uXMbgJZbfl+B6tb2oCgubVz7j83HhPmMENCl
UjW0oXI68BaZylsHk70dW8hAWKtJ14BT2j90UzwUJA9li/q+3J9UI4xH4H9/3MLG
ip0i9LcUvztjMIFtwn2ls1muWX38G2qEL1tpjktryt+1iZLVoQnf+z5D9zb2i2Sn
yZLOrkNBEu9pj38pLFInTdDlXQqpjJ9PIGiCBXWrcYTbdmr0VkylF4NnP7G9QMvk
05xp+TwlyjtUq2V4zJoOJDcGqru9Uohxqat5p+Hk6fV0b44aOYjF+MBqowPQwHg8
k0IXvEdI//fDzc2M1bhPHlW6D/7qGipR2/8bkI4H5yRtjztC0bdzjJM4+EAkSOfe
1EaO2Hd7L5HvjPRJRvE9DEDuwC82en6uRGmT28aMKPK2zeGhGnzBKWjWpZlHZUEZ
wce+lQzYSySegmoWzO5vSM4OUAbuP0bgIeJRhUlfoB31B82qDUUsntHFFSJ7zO1e
Nw3ciJL/+eKV0XfbCMg7oaia5pwLkZbRT6cqjpPxUyu5v2RUsZzkcR/h0vMyJr/f
fCADMttJBVUjUsU0Au+qg5O9+FBKfvkY1s3IGumN5LH9HzwGBv8nrTATYS2VjiyA
szItx3LgKpXpSEVSb3WfNP68Xfm3g7OETmn82yzpu8FLlqWirRQhOWo3xo+i32OJ
exePzF2sQD1t+Zx6ngKnuGTbHqqQLJHT+l2NsDLxMTWEAtyaFwL6zYOLBs4ZMQJB
jR2FrpRXZaO0ev9056sVCCOQ5QEsyNZS3qCt3wA7sebj7PFHl8FJzOmb6U+kx8s6
Ghnv/CTEEi5SxwQpUxSN1vv1JWmqJGeW3NdUZJJLGvMbT9xmT4PrCvW1VQhtXrB5
gF6QZWHy8oywa/ACBL0Mt4PyAxhWPxpSsrzi1GzSiwQ3Iv4/+NV69WwHlC07/jew
EH5bKyzmfkbub2QtHMhfjVQXT1LPRpFeAmaYYcEwHzsUqpcOperY1hlzVsm2HWVK
aRYPbxJTW4AKo7gTerRCm/QzIhamcFdh8S5Gn+dBOXJmCVvIVO3ITpAFT6+Jl/BR
NQXjHwgfcGeDPhFFOiTRC1WuURQH36Ajq5N8GQu+RHpyWH4ZCm5eA64xqOJqU7PV
wQDTcJHJJ0jqritae/QVOCMziTpeVg8KbkOKkE4c48eOFJVKHCMlXUF5QVTwu2V1
2ASfiEtC4YYgYA700iShtcoePw+c4DtLrIUsY5cqufQ/nQLCSlE5DCSc/l+537Yg
SuDMSYw0eerdpEN0Dnks4P/JP0rwj1z0O3L17fGHVcQ62rrhVbC3N4m3Qw6CXCku
SxseO+54OC54BX+CEc8GTBQTXdJyMqIg1KK5XmcTEyFQC5ihQ6RhRWpw7DrKJQYE
V6DcvPhbd+i4HKnNFPorp07rhKEvKjH8DFm8fmYxFxACtXDfbJORpJAsQL/5PtTE
st1pOfe6kF5naeNIdU3dheqqjs4IXkS6f+DsJYNBJI/mDcHTVcqv1lRRgbg4/Xsz
EPO12jZDPOJYebE5ofNv5GGWPA4o3FGJEAB7YAa0M7YvbG7YX4BK9GZxUcHUwGvj
jXgqpKrOMKezdBBm90flb6a9gCySn5QeTNjniV0zznvTo7XteaVVPwx4RSOHKJwC
GULrL1ZC9/k94G3hkMgqPZOZ3Zd+/qGZzwDPOqCv0quuLMDfSqUCJxZ3BrIkGinJ
2mqIlCelJVYr/kmIvRfDvaRLDmTAFOp3JfShBN9T6IXZTYIT/UEtn2NyNYQuNhvP
TM3dydqODnTaHn8yByAaWtX8Cyx/9eTmP+Fk7nGaVAzAnpyOrF9VOrAIFvcukMG9
+0KE/O4t+/tNEZOAJNX+ZLIJV/IXwFLBPcCtx6yxgXDDmAJKFTtJ9jUFBgCAsz9p
sYy0jPvmHZNNdqQNIeQzMVetgE/uPzeQq0bg7Teu/rhcz8I8qlbe5V/y6mHIJoTm
9pJy4DdJQmtdCipj1mD+DFVWjl5a7PLDhEQA2D5OyjrPaoaaRxmYvcJd5YOqFJ/9
L4XhSJ729xtBmaCYWBOcaOzbSRJ15biAdjh11w1mO4zT0oKRQrt9q37W9UTEboVm
Mz1f8iMcj0U2sKNeMOv+WhshCeS2ZPZh61LrLI6iJM7KCjlMD2RbyAX1TehToWqU
jihVQa0B1lQgWVfcq7WoB047NTytAzA91WZzuMPHduRQQzyW83UvMy/R8n4XOVgG
nH52zRk8BZ4U6G8yRX4t1PzmJPQ1FJFIuNZrMsy8NvmzdsZcGy6ccxfZkhaesuyr
+kkYo/LB6kIVwwd4/E5lDAynmurBosQZhC0Kkd9UU/sUGPqlAZLvAYCoH2XyOKbe
miv9clqr/j5KzoExtTkhnYdIiuVeWtmJvAsDdkYbSwvskxgSpHVbC4//25nsUPl6
Ic/98/w0JC0c1cPvKFa9ZAyhmN6JKcptaQCe1czrLo9PgS9Iep8jpzW7HTO/rWer
eiv/zAmaeiJRQwFt4xlqMGUrXptxTu5enRFAEI3e0ILWydLgtBw5aFjF3RPoCvuK
0up9QZbkN1FnEKMLhier7xJPJQf9NHvNm0QxeMO86arjjT8THvReEOCMmDTKecPr
166LZjBlhEWmfvpRX6xVo2iZS2ze+mSb/NMqftVnctqTEY6p+Z+B2QS+PSWopHbk
cnnrW8NFnx2oxZq69o1EEvj9dAgrZ0WESy6PkFmIE+T2Ptss5wCZIGkUtslO74Xn
PhtlI8IZh/AataOnRIqW8c4/rTVyaig6pio+3CiNBjT3YCssQdNR1tDAbJJBg34h
PdUUV6V6pyNTF52QMfMNJ9kVaPQ3uEy5t+O/hgd/nEYxDcJlAgecic4D5t2F72X2
9pRzy0DKbqFAi3So3JY8F8+dHI54h44c0KtcgC7Y4PzBV1a4tGnqWSNm1wVPYExj
hItCI8n2ns8BbFveKEkccEdvxCR33MzTGnRi9APmKsnyjMDYkzfEW2mrAwjrUcAr
Vcz+52sQSpyuw3BIrLd8pEL/gs3DFKHYdrjDWyUjb+7p2ux+slLUvZfKZJ8t5Kt6
bUnbFET/hRpYo76ElxThHs0SJlDurBl28DokzPwxUcnhUCRsiEZZ3a9UPw8Km9yx
6OZvZWEFs7P29at9Eln4J/XXTn6TvU9yAJX37Da6/pZWZd446GwhDN6Gf9w7UucE
mWOgAWa2gpmtWgzPN/CWPW4h/rEDtj/HtU8cKC5CSLQI1Nyi8kGIjsWgN+av6ecE
2OiQnIzCYWQBQ+zVV3zfnYU/yBkoQG4I883es980lMlHjk/3ToVjKdw/M/qEMm6c
PfeN5IVCaC73YwjxYh5bhTa3GrG3QCwlUR9e/lMFoCqcTx0a8UaG04iIEmveH/7R
Ino1t2rPBK7RjTRhgeK/taHeDhgYZ2K8bC2rPh0aL/5fKOLcqZYkM0vhIp/HP8+D
PG2b3v9u/E+KPd+qbzKoGCjwaogKysMW2al1XGrq02sN+8KJtt/gGty3gX7B1wbe
qNRzVDaXSsSDdZa2A9zvsmczMDW664xgz4t+rjlhcn7ZbXsLvFNFEYytcEUtzrs5
taqIn++Gh/z2HFBwPEn10CIyDV5OUiWPsX/Qm/T5qx5l+RkV2EsvfrCy+n3LparY
zAHXqFGJE+ZuLS5cPqiBxiXAXwTcfEoJ/tCLfKc1gNmB6W8sZyKf0KYe/Rs4ySvU
wq6KPuC9mRG4dN92kBup/ZUxU22xd8p8nxAHEh6uylkmbTrGcHwobEXElpKnlq3I
voTW0fvg5yhU5HhFENS4uXcpAqf1P4eUUuQJptxM26hckVZVMzsoFqWZEq5zoXle
6W52N3LszS+5AuHUuujlBDO3q9k6W7bU+DSc6vagmdUa0wsgivOqMNYCnLQPi4Pz
PlATM1pbX0tPYypMTzlFMRaIfgRVFJk/YextOYvrr5T6R3eG0YIi4unfEqaz1dqT
mWjpdqCHR5QFZsn8CdHCFrF46xDKkUulOevJ9lPhclJeKR+aEqVbu6SmhhqqQKTb
Ibu1tCr299JbGpwREY3dww==
`pragma protect end_protected
