// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
kFgDz1/pOOG68hED1iV/aJqUSLKGiz0LBGKDqGQZYMpl7qDZUgP7bm8t8Nwl6aj6G+BZZjOK3zIV
rTgJrwIZoexwy1vuvKHcJDimgSi0fazPy9Rd0A6iRtjvkHUp4iu6KTE+ewhKlgpks+YSr5bPa/9s
t0puBcPXRS+abcZlazWapx3voBJw7cSQY7ZlKWBUFh207YCqAgjpqZPsR1yOcMrRzYeiduJVEbxO
IaBEbubOzlsekAe5lkn5e1ThSZKiXnT0UpAmoX/Tfo8jMTj0nKRCYKBX5n5NxHyjZRwHA0DgpEjP
bKbYrvU+m6sLolylyhaNcb7CSjc1HYu2GzlXbw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
MiN7LM3kSBr1X+hyYKTC1i/4+Jvcc+TircjG/bDzDS287ijiYCUmwloizISfHYrQCyQCvYb0uiUp
3iIOH3AoK7id+0IZMLNG3gCAHUiEqPMNzSx+pTppYiwIrmL2RfDC3vcuiWcyQLYSu+jv/rk/81QQ
siGry7hKj2nRifTOtePVygqjq5ZHsz1v0VO88WEq5NpEXWrREiTffiMa2IGCA7Gh4FeIpZWz2lzB
0hrvKas6tK64Djf77sd/ZhSQqntmo5WWIIFUMYKj7RJiFXRosXRDV3uyUkvDsKMKbfA84R24h6TE
6+gGhTbeUK+eYV0lVCWqxXArHf79pdMBgK+btvwW6MrUCV+SKB5mKq7jjqDu2d0amZXzYbCr7ULB
7kPh9qnN+S9VT8xyAUXTNwwVrOkAUK61wl+Ev3TLJOGXxDK/Z9eNrwYnXfUpqOHr1N1wVrQ3qbAu
O4d7A+EjoHrwzGmQVNlrPAbMjf0MKVYa6Uq6zoixhMqMW2hb7oPYsxyqbWVhXZUmgNrIrAYG7f8r
8HE9szCLE51H/bXSwnlTap0VatDFpDcOd52XrJYJYSWDrY/37ZhbU3fw55eWxCeWzBAESBtjaQGK
t4jtqYojYszp6/gXfMXPfJMwfvesbTnMSBJ21XNG2AgUHpg5c0fyir+Wi3MPA1YAgOp/E1TfEwhB
C/PJC5mfLn3FSe5faa+u8BY28GatktzbRD+eRY/o30Zra1Tta7wcowYSg/V84GDCAWPlYj4Dz+IO
h/SwwO+TqcOMDc15cpbiwIy+VYlwDr5hzBAch+vdnLk/4Js0ohZYaNCkWG3KAl60lvkcL/e306hN
SksJU4ELc51w0chdvmDHl+dhKzpXbxNXIUtGp04H8k1jpsym0CZYTPNdTX8xnCUv5KTRNH8aqjNv
kbzOy1pggX6HdnLoe7GPaxxLybFlnNnHjEc1n0S8cWaemJ31BVNaf/dxZTmMG/ZTUQuHsc0zqz7f
mPzTr1GRrhU1XEve2ub9P9uAZ65fDVmIvz+NfljkXzJFyuswoBrvrR4Bwc+zpMb7HrF4z68KclXQ
8kD0UFD43m/OqwLfY1arL6CaV+XGVvO0xmcJOgc0MDHTAIRry8rEgPaJOSLhKlymyXsXroH6R5y3
0p+cQrKn0UGcmP3XjU+hC7+OPC10FYbPMCHRXAGBJQwEiyZjizgi99qdc+fl2kJjIkCFcVuuz1tp
jX50UmAsHyjqdBNVFMIzYbSsFBYwptecw6wtLpWfbTEdu2hXwAQX4abYFtB+o/rs/27DjLTJpofz
bKaW384w1LkrWUgr1e2kA9OBe0I8tkQh5NLRnx0fPcyrfyoELz4rFvbg7NTqTv2Ff2pbDLbjmARy
+mHnW5SA9Q/ZT4FadC4UPNn5tRXVb9vUxA0/QMY04M9Ynux/EAuD607uBUHN2VKKQvoYuOmB2c3V
4YKjVcIiqzl0Lss6981zaT25n/1s9jhWgT6HcVQ1WkWza5HTN6gS6BGbfHi9J8qsbnzKn8fcYYwK
LvuBcK7VYRm9B1czMnqo9c0nRysRAfJbajHIWY+ZgGi9i2FDb8H7TJlJAD+EyM//M7XZhzYSAUF4
vZH22HY+1FJJVpGSkkFD9nOcGZywvtHeK3kIUVOsx2wnBiN9srnrmERRHZSK88zE1pWKVW9MvN/M
6qyD64MXuhxH7BvaZ2HDEOsQW3ZNCxlkHJGGDfk9CzmVJAsmWzkvYCtT9nAS/yelViHcdyzEJNk0
pftLXldivjNzY+aMmsd5DjX2vVCiU8lD4FWPLSG7XJjxdqSAGNqzuvIGobQUov0pPmnKqc/B4/rl
ZDhH3AwyG1jXTvQl3UxQ1PjTeT3fTeiZGnKEOso7+9ENyvak2vyeSJssXpm5Y/BNHcEQfpaemg2H
GrqsLkXsGtYPY+P+LFCTTUTDNzMP8AXsn2mEwKlGa5W304aCOrZ2dN1fr0ru9ez8geMkO2L+nhiZ
UfS4zFOk/Cf0fkuIwPiq3krt4BwrdWbPNb/8JT7LTJvEMweOQJt2DZb2Rbx9kZVN8QMrfvuhfuqL
UOEtwWQHU4LdhQp0BNCbrCGuOyBc6hfXaEV5CGOWLJMSc7/plnjN3XZlC3qtRQlVfZLohupuDK6K
ptPp+IaCpqCl8Q24xC6V+F+A7+YyCo+czpwGqg0YuWtNApyYE6fqZzMTwHISdMflL4SW30P7QVej
tXrEVuqhL7oVgC0ay+i0uteqDMVusqp+jjIjPUFMc2QA42NdmpV8JRmb+fAivuWkJrd4jISBv+zS
U2If4lrBbpDpubcZJ1qAnA8m9669qWdjwE9/79/0OUO54mWLv295YCtQ14PQTo1K+5i6rj12Vm/7
upDMp099kgQNA3xuMO7x33wzYwXhi3W9Om1JBrG755u6uTADvEc4zRHtahcwpUgqrj4/bXELNpKZ
/ZfTuFrXdwmdAnlzwAt/DnZErYRKbNZxSWTLelQck9GBFnpkStpKuiZVN7Uxebh+0GXIFX+Fitbo
u2RUpO2fDdHDQqKGvwn/DFe/ypOVEoGw0opouNNa4mDRp34TBZBrE4WYebGOw23xgPHeQq4lO5cG
MiCq3JJubNJovDnqRtHyxXUO+4+eLGXhedZfNtbIxIkdVG2o+IdKLA3ttuw9DL6DEzM17G2SViHI
ki4oGRgUn/WUqAfrvUKuu2Bny2Uhg44T7hViq2iw3lIgWW8ypnsKeCk1pygmGx/TbABWscmraMbq
ez4FDMu8IAwSe9rRjAHSmoCj2FnLDxzOvULwDZLVlEBTNxCSNMw25XGNPdKHIEv4dXVJsqhILtPq
tThNCpGg4Ht8EQlp/mSlRzvi10BePR6sL5NbEy39xbyFwnmSbP3IQpiildvVjN3AEmMnNGimeyox
0OCNRW7N+AFNCAD+fAC2lhuysa5TevPqRhN2yvGVUOCCjV5w7AIqZPpWYaguhmgx82S/vBEOzWpU
npvSCllBB67uuoKDKLjbv8Utr+jbaU8JAffnZJGieDOIm/QSwTEGk5XniLhtQDpV2Fh0xjTFcca0
oKoYkJSjPrxN9fEGhz8RpjDOTt4+KlezTQhESq/1nmkIzDs06u1BM8uAbwEH+hGepi+sRYDV+xf4
b+A6XQCdkCt8hXK0S8/rOc4Jtzp1vGUJW1F5YJ/wWkNvZHlt2UhKjllPwmL3sjJgbTC7eVH9E/aJ
lkYAfpxktktsldI7WZ9KI2cOhBJFiuQ3MQVj6mvzmAj3RYBmnoMK5rcrTwMzP6FN/LrIkS73JPPV
oUExF673JJtQ1Y8vJlCVmIkxEKVF+K1LgEAVM05vEnUqk6PZnCvwsug80WmchytLffKS7eBZNj/8
S607dtPPZcMYpQ4K+iNTbzzeWalGAttNh7Fr1SV6m0r9e1eOdrLy6b265Ub2bvCXEq/E1KjOeGhb
XkLKjdCh5vBFZ/jZt6sx38Kd/crlnoeeepeO8uBJ+UWpAzLjfyGZ1zoIiqxf84crhgtOaDR64Ky+
N8nkFbZQQAPQ7mgg54jQVgKzbuPXxBv4C1Wmvs5wbdah+dhDWqU64wxSSHHeVcVJX2RWZHHM0vnK
OxeFGcv7ZPjAcIAZpd3Ei7JGDVAa1CA/DYPejudtgJ5W0JRBJm+Oc+ohCb+SupZQpZHLksh8xJmy
RoE941FGsQ6imDOOEyGmQLoyxmJyZWv/Nl6innOJIn0UgkdIZXaDTIFpyRHBfd7zF93VEmSMZ04n
ZxPJFvj/T+bUJvcu//d8cgtogBDLWRSre8hUoowB5cRWcaGvkoRXKMPXymaX9XZnS7567Rk1rUkg
HB2KwXQ5GqewAM/lr/SZDrth4ZY25U9bun6cV4yAFbl6eXyyq4zFqbkyxe6jBIeZwBV1ddg1Wigh
nl9RSOYB1Pk3OI7HU2vZf8irgV/CXwleZqbqiUb8RXRjsSuzZu4shNHVjlpeGeod3Ig8nAkAP9F+
WwtUZROkmjK8lA/BTpVuqdjQnpaFze1lKSkPIynxA/iidBYffeT3I8X875UAd8An2RLvv+mAo49U
JFaBlgftY83wL1+/r4tYVGWNY7IOJmZp0TcoQdjt36Q/sKKxveAAOpmBPDBjXtZoDarsRafzrl1u
yPR8Gerltvfr90C8QR8EjMzb9LrCK/yvgHDx8D8q/so2WWEXhlkB/jftbc9WsdIUQ8DadM/zpwVQ
GQamJEGGxKjwwWuv5ar1oPLHHctq3tmGAiKfDv8LjHccg48sfh7U5lANXNICFetLMVV52OZMhNK9
ntFTpKxXLzNBc+Ce+ujL4/dfVBA7cWxspJ564/QAKgmf8fGOvKxW36Y5eOadu6ippZheZWNAijGI
6WoFs+ykxkFd0CWuSGwHtPAx5Gi1YGgevMGQi3tU9UPdrie4/K/7Ad/DS2Osxh27fAKKTnXco9mc
GjpsVPW/ihd+jQSouC7C/dt7kz3Jhd/lWu5QkArrwPXsBmwW83F1hKIcA8VbNMPqC3pwx6umjn/V
/266iaCfBKN+6lfTfvf17tkIvcS4jq5JRtTKSAFZ59CDEm//naWALZbE7SYP05zWDndNVg2gqUwY
pqpeUx3p3OK4x+a2WjMavWM31u4604cp77M/U8oPru3MJfkpKUBiDynW5ZjkYPjTryVhi8uMjIYR
Mp2jfj9VIdcb3vBiR60rpAJf/4eWkEKhimwcJliOcLgMfXbi2L/dkDYQI1Y0fvhPv4M3CdDcHZru
vw5SGYkhZ1qXdFldlRs4idkPPpf5Xx+ZUyJ4SMjK4wV0JrpctW6c+ez5c/LAU6vL8JTDTIo84+Ux
hVXD8k1LJQW3hnB8JZWbK95I35+ZhHsdDKTZgf7yEr6b4yLk+0ZHJFMtjPCWb/Wlc95gkImyNlgO
8sybBxDJCRyARRz6qnHfmLJc2ZAYQFskZB4/+bus563hfDx/rgj2DmjR0Mr2nN8CAw7MzQStTVNn
ryFdi2dnmtdDugSYoTAcu3EkvJj7X2blC/vMVbhsCt03pmDDj/CfsaRejsdRSAytnMgolQncK2O+
RKOcDijtp/9Q6JB5784FQFnwnhIwji+iv58SGAJQ0RS2OAEAFWmhDnNrwubs7rLPZkTq1RMcs1hG
/1qzktjNIhl6UBCiTzoXHTR0GY4jrqpBLGjiOqp3l/EFrUjJBpcT+PYodKlayPySCwqj0MfzJSnd
tnnqX3Nm6k69ncQQZP5KYzgnl42kjPCgFtTNCtaCpMU8byxuNfdgxmNTo+ZKMGoRU1/RaQpvv6wu
31u0sd4ZXZdirZI+D9WfyU1KgbG2KrzMKJBnjofi86+FdVb0BpcU+qhGJSjALXZZcTkUECxro9bL
VCzh6y8zTGo9DQcMQN9VFndZ1qcsyltj4Xoc5yDQ0zYqgB2vA8jihrcjl0OU4Qm/mFWsM69vZkhZ
InLX3VdeILmDgKTqfgxhtOKfDPfkqgKN76U/hIwskysI1dq43sGGOChUTssXieVdbZjwFLTGMPXF
AhGd2ftp755A2wtI7Pubdn8V4L8qNx91rg7JwafdGam22TpRFRfNoq2iWUDeZ/t7YVu0/Q0UvvUI
Wv2lXhFEreox8WfvMQNlIwNOQVX9Gdll1TsFwC0xyv6iLgugurypND3pLF15v5CzinVabRPem/fn
vvU49Il81KblS+1zhRODW4iNhPwQqbCFNJNR1H/10rXrt8/wOYh9IpaVb9ItwepaDqKDcvcPc4sV
M4tJPiunhdX0WvCXn17v7cd/X6LDLQ6LN55n1O08Kd8pyNz3Oc1G3tz71RZbnsMKCiDgjj3uau/d
YAXbJjvyXESZKTyt2hKTxOXQwRMLRjGAb+g3zmnBGCVD7eqBWx5dySdAu4xPFcjazXnzGcWsV5J4
SAWbaBtuJgwpMMUA1sBg+IRR9Izz4Mxg1yTP7/zl6NIMdAJXiPjsrB5JhgRsAl0cgaoC61+n5VW6
ek022uBzcDW59S6uoemeZc2EcyFV/dWAWvbfHJr1QiIBTnfIrO5j7ozqc4gwMqm/xlMzSOfx3HyK
o+UkUhHSWGFsq0Rd21bmVWbhKf5T5IjOtXVoVyZN1Hhvr0sExsxHe5IB7o3qtU7uO8R6cjc+mPDw
wflJlAJTkeOzWIsEWXhVgcq5aNurHkgBwwfjBzopFYzWlL0qsrOxz//92neM+JJAb99Gdyorpp+Y
NVFJTTUI6moRV+QfhG4UhIZx+ooWC2yfHdKOpYw7xPLI8pvfnKluMVO6hCUjyy2WjJ2OJjxJMomz
tnfX8YNtDvP022wMocxnkRUklcIdPLRlk7OX2Kwk8AdbNK6yilIOw0Hy01kV8gqIftnodifknhyE
jnMg2NIBnkDWias7/xznf23nH+H0+T+TspZiqp6e18uSBPYpHtrlx+y21sDHy+51QkH0HP/uFYI1
WcwwsXNFMk4Y5eW8JX3pF2OKHMJmuD79kS+DgXEHLfIx/Hz0qHF+BZjfkwfpwjLucLM1Z1CdMvaF
vfw2BnVggHyDlaBsHRMGcX3h9did8ce+Ru3TqXfsa3TJj2r561iiBH7itbR9NPvFzJLKRgl+lCtF
TRCkMnv6WGmuH/ZEFeCYpS03JL6IXcu3rZeY0oEdWdmFjoWAmP++scvWonjC169L2QCQfI4i3ZkE
Wb6Rvtky9o5eyrb1gyfgWSQBBSJ0dyuhuqe+SrEqL7CgKU2t4tWS2gzjPgKpNsphjcoiVdURQ18+
eBgqK4P0CM8hIvPrEn+zti4k84rTjC32pzSbGeZwTLS9HcAScAVMF7oZF957T79MCLPvxWf3ZB7k
BGXLwNrONRL6lwIRUZfq8sSbbUixW92tOhJiJpo3ldGD+LeFrjfUKRtOCuRGniApj+rEkqBCIrW+
Dcaeq/v4TSfPomzd6GjVm+EGNthPD7xx+rnY8LjvT/9hDUZmrOhzw1SzO83sxwDfxfC47gEOm8jJ
zPWw78h67lsh4t4p4JJRmkNksbVwv5tIbqUopOIWjUHFZ0uZIZb1fUyjw25klKPOazYcOKmWpLk+
M+AtAs+FZv/1hi2x+R2DnfkdnCSd7BHCflXEU4JG84QHx7Ao2NozbrBsl3MaYoag9LpAcfe/2QXs
//ricTc6QKimA9fIoO18z3LT8U43Bz9Ltfc1jjXin61c3ADo7Ct+Lf8yyPF+fN2yMUIG5AHUAgfJ
T+js8dDQd5oH2OJ6l/PTRZwl9LUWyviftacF0K62ZwTSdao8rVKIDbYFN9Bf67bS085BYsHQReNx
9lv7gbVTNJdcfkoCY9rdYfiSTi/3fCXfjo7zFydMr47kG3sFGqGMcgUmzGy1F8par7oMyXU/HxKF
VytOCrZlsRoBcK5XToErrs5XtY5rOTPXE8tcSGxD8AoE2jZOrn5aHVOInvs7B4AZDyYUApTsz09V
6exspOCTe201w0S9mvQsRvENa1ntgvoUTlgPi7bGAiOejF9S4iFMFyYi+h31zulc96vFRconwM9E
QKvaih9//QoQRLVBU40KlRBrsrW9rtdJvgyrcTqboyIIVw+U/LjXeA6Sm9FPNM/Z0JEu7On09GTw
bAfKR07dsFp/oYUVWob8+WV5mKT/5VVv8spF4Q8+LSO4A9WOeO7wEA69GyS9lVd1iZo9Rn3XFojg
JO5Gp5l91ld5cjVaAeQTN6qSJgpGRJXDM6aXS5AbK/faxR3t/QLZHdvqDzDio7krJMbwH0B5hzXW
9khu/h5+nhT8RCmLjw8tOxhI1F1ifUUlnInKaglEv4zXhJ95TBjTYOmWRnuUcjsJldlhywx2nNYD
R9goZtHqeQqC0brzMGmq55aYXE3Wux/1CI1F7Jow4I29b6BVbm+GmTy6+YM+qf4U1I7/JWly+4NI
e1c+COSXD+Evb8sIe6mTzQEjhvszLUadylNPfHcJp4ggc/xPNWWanFT5gzNf8inMe4LOh6eqsMZ7
c3K7BgsvzrPWLPpEB33QpmzH2I5JyS3yLbZh4fyiXDvXCblQ8MF/0vxydHzYhFItAMGHdlgwl6TA
BM55g74+mHW85ONhFZ/1VFYVDOpsBkfg7guDhttkltXAa44m5yjgAZMGiUvdkEhbtEI13tkiXLj+
U030wgXZafAY/5fS5nVgnl6y/QqAlc/TihN/eY1k5P0oiG85WbgawLlHIwz3CuNqEH0uiXmPf7XS
nuKCqmGi16qrfMVfD6OyYfmtXwdUbLIWw5Kw6spPjdqTaQxhXB4FCFSkPLMd5tapcUCATr0l+TBP
YCb1042GVrRv8zvd4u7OUF6DldzLgm5+kCHeLTnBpBgw5oNs5zqkfU1wX/tFAWrVA98VPzrJhQhf
Gc/mRDYBFT2oMbVdLX44tLICjOPX+ZrXp6c4ojI+RajOFEU7nfy0x+GlaxlQPiwytwz7PEC6IK24
7F2HEm84VYQifLO5rEvqQybZLVF6FZKUjihqcdtxg80kxIJDnNMgGMsmy0B+q/UB2Q7ws7bpOtO9
FZnzZKZ5JbHPt+hulQyw96uymySd7ZpqFDRejGvzBUKuz8/yYt7Ahdb52LVNVc2wt8vJVGuoWqBB
tyg8E7D/hHdNCHMtjZ93C77GgjZuwk/OPrqb/uDQ1qdvvhXi3/R0Bzk+MhNartSZfLIZh2OKa1ZF
jfXAnx2a/WW5x0rLOROGjXcPSeZnPL/4MJeYyII40IhjVo4R+/bzZFpXRXS903/KV1tMowzYhQAG
Vn4NU36oqf0xCnohBbEfiZYVf7OZ4xH5aDNLQqLQYQuBNUdw7kd5D0C8EDI/MP+K/EHqaIE7yTVJ
9D4Pq4+KB2jMns0ie1Y3qShCO9TfBjjQE2jf9mEZOKGKjpkqt5HRmj9X0rVxVjbfKomUPwK92p1Z
LLw5Q9PvQpyH8pYQ1oD0mzr8lmcwQK5K8XTMdmrhQbs0RVADX+43+MEFyn8w2kDzPF/OdTfW1tBd
Vq4wNQlfJVgteRxzVwspNmQUqMjnntOWzsN9hn/u+WFgLk7R4pRoLEKxTqLnqHy6o5lGv5Sr0CxO
e6nlROS0sfAWKCavjjLqxXiPBt2tXuPFU9Ry47tBoeex5sj/Qmd4NOAuUkCWOC/q2W1GO8hqJ1VZ
c7V1UtzP/a2jEFOSTy4DLrrG5tL3Iv347EwF36KJA362iaISi9S4Dr/IsSat9L/otir3JX+GDORt
n9wtN9kPqoiQvDf7bYFd+NbFND85SPtSWMzhnTF+wxBwVNimNcKAYxL0AxFISI8mXg2KN8GaVKmX
eu7BSyIBcFVu4YutpHMWoo4YljnUi+uhL8ntAwUCBcLTTt+m3mlKZ+QiaCg/A8rZaoyp/ke47GfK
KpSrFZQXOlmsl14jLy99O/jytxCDdbzwFBfV5yuzFqTvVleksROhmnEvTtFDgaVu4jYmNvpRBJYe
an5Y5HGg/ddyYd24ZEbrjWrh9e/H3HJp8dcs2vc3u68lDJ3ukY6RmLuCpZphGRkurwu/8bCoIaVX
nXGTMkdnhkgu2tycJ9rL9Ou5SyCIYs1t4iwI+ympqEgBtbj1YtL1iYNrCJKLi6kUlRB7tmfaX8Rm
CDyWfaKYh+HTuSY4qZXm5E7XugDwjmGn3B9zBeSlPJqmQZBRax449kljo4voOKvqmrEMgPyX+Tfc
BC5AOSXheFGFKFXdH/xLHTxu+QWUgjVJ8xSqiImrTimjbb+jHrQQYpah/M083gXEh7AF/mfVQwMf
+KuA9OpWVZHI+93QGB/OeMoxGp6sZaN66d1M0AcSiZF30jB75K7SMQtkfDr5pyiJfrk8HgJ5DFFX
gjQXTF8I4X0btBNdvcHsnn9CSj+FoJFnZTooo1B/PSg/oQfi0M2/kJ8Bc0CXn1FAa8AkZkDRiIoE
EosTNryTH02yx1UKJ4UIkUBjrKV24pmE8oQ29uZ/MhrX3xUpmfpO+IMLnaAfStyEJs46qfranzwC
Opgndt5ZWc4yh44AbyZzXI+ueytbQYyoK97y4jylerRDG5WPNlRwPWSztWvBxkjx3gJiW9rMU45s
WSO6tU2zYZKvMmz+mX4R8Txz9jS77d2wnvWQTAA5nWJcBRosfSOJiG6kPSvz7fpSbHaFwhDtHOyu
0R4YYXV6+JpXdsBIXMVS3qSsGoOLy5ohYTE9k+FCmiHOWSw71y+eQ0YLplkiqiAQLtCSAiiBF2+E
QOKETq0oroQB0+4ijsJLGiGrgxNtAHJugioYGd2ChvdDbb306nKRXkOWe7laPv332ShciAPmTBCm
AetzQJ+syax2nJgTnTeLW3AX4xFcoAS1jNF6opg/BQcdAdcyO/Jo/bt8XNu+/1offRoYVkAX/ycH
0vG9iaIgsW2qiRrnYUvpdN2H8eJ+WRKjr8d/9fy51zxofDj/C+NGpPE3bWDkTJvqAhAEL39mCmOW
vkcQL85NjpOUeiAZWiDObnaGduL7eX+fKVegDSAaxb+6ZVD9kfT0I2WryYzbg18gf/phx4SIVJwx
sKZ7uaF2NSg8UOaDYPK5Pz+buq6Z6e5mqgxCJVeaDI5qZ3dhlS2832VHmFCPZVniuR3kr+SsrQLQ
LLrTbX/zkP/N1fdQ3zUGa7ZKVaokCiDvje7Nh2GRwhZG8Z3VwEp0V4Zbc+rqLUBMsfFikSBwz29C
tX+oJOmlc+xkmlAKE+SxJRUyM8TqhXXUD6MMMfygWspZXuoEbwTiKDzj3ig6cyxjNQS+Vd80Z5Kh
6ZDEh9aLE+tZSfMLWFWD265pwRfabkBRp0eXSr7OWbKPfuq/iB8fh9hlsCWAvTl7dsT8QEFxUz53
ybaDgWEzXSUB3sSbggqobqEhGerSHzKn3KbcDPWqC6e65NqdzGfsC3qPtv+ji1D27TAP1imzguNx
GVI8J83N3B9s4uWJlexQpsicMRGzl3hMsNHdKf3bFZoBUe20+Sz5vFTbxrvxFXEVtAFxS8L/jICQ
eTgvONHdp3xyd3YwZyrzQ3YBwFkC8Np00bPsi+cj4LgjVa0AnIToBU/rHAecx0azeXiv8aWQI+GR
qysR6SM+WYfBsPNW2WjYgmXofmg2O/RYzuGqL11nHvUxnzHxZK7IdWGQQfBUcxyh8WlLcRmgsvT/
76YtmWDVJMAzlem0mwG/7gQMZc6vVmBsVrbQ41e0lNvJSHec8KmFe+8g00KJ1rMHonqQF2vk9ls/
C3kgQs7njhiqAMuxr+lw+3KegJUiGk8Ak+K9mN71W5Y+JHHSw8IWqiBQenoofpe1ScaH2/Bz7NCp
ajQ6HBxCtdFhtzui7gOJVAK1SGhEu4oAhwja964rzNs5zPZLsvl6xFLfaM5GfvU3b8/rHYtCjrg2
drGhpeh7OMjZdn0ksXtLPIQDskqwrQCES08vfbWdwgNyFIvd763MdS8LMtR+kLxlAaPClDQ2/1KY
KatgRzU2VtEPGDj84b3zVry4LUAakzYeIlwAz7GAzsGlNVzms9bqaDe/C73ILrcT0EeDnhWHHBau
YkDBH64BV0iKY5u+yHhZXTtxBDtkYpAKCNx83xsg7UEC4QzZeFzDFog1AhKdU2ESxtLSRk6smJmH
SGX/A0oDsUots7cwEnAhmVGG2FjuOu4u+AzLVegrH2Eix8FSm1JE/+yLEg6zF2FOBouEA2rOeKHk
ahnXpMb7A3vLGWwMg+9gOQm9gP3K2qbr6SS0aHAlC0fe64G14xvkXtGqEjQC2oYw1qWCYQp8AQiZ
nH4Kjk/DZ5iQTdmR0hYHgdG+Ds1d1jCP4SdvbX0ljkOEj76bHUAekX66tbaFylXUBkrD36al6+rV
SxQakYQMF8EJQqy5dZ5pMq13EXvMKr2rjgJMi3vc+8lFeGz0xrTydNkiLi0uLrvKWw0kR8PIOZo3
RvDh2tVRhKc+HGldfY0H8E4heo2M7KyfYL2a63/194Nr1y2PpIx3y24QMdWdgDqNxWDAjsF7OduZ
1FepFVb/9m3OGEaOfywEQ/90EZl8iYuTtOx4TazccnwseLaN4tRsB4H7ElJb9Hoh5XC4u6whKrTw
L8kwr+mGNU2nU37Ty3K+xKEU9RsmMEQEP+noheG4zhWULeEgdWGcqwW7HvnIfdGcne5UnDz6F7sB
da14LDNpDsnTaRCT4USHrmomL0TwqWTSD13PWZ1TSYkzcD+vhfuLMzeS9pzqVclpyjaXoluYmHfB
NFulj6ESM5RabEZqk/4a/hRIcAtYzb0GNev7Awzz6Pr3SV1YzgwN5I7Vp8XJ0u25LWxjz8216Sk7
umxEVqvs/zQPU4BT+4pQ/TH7kB6jDMmREcu+V3+wvShWf3AbDAa16pQMufR1Q+FQ1FJfEgYCvAH/
A0j/WUa/3e6T786Qjs9upG7tb0Uu2RjXshln1ZyupLev2d4MV166EIn6DUZXY7fQwPr6/XuYtUJl
6+DChLIqhi/Mb52OMhzSL5ndIJ5d2YgUstsJTNbxU0A75vx/E1jB/DKex9G1WhQQFGPHhyFzzLNr
Is3JHJ0goxfmOc7nC/9RTmyLI+Bnav09U89kNt/gjK6R1A9yQdQ7j9rOQld3wbPCw4PTiBk=
`pragma protect end_protected
