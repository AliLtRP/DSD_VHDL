// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
cEBGxX/0O6JZ5UZ6FRyKWby/hE9StRDKTu0LT2sYALDgPHDd24bOTw8XxEc+9FzOTkMerNYMsemD
sSCg+8A4vqQcX2Ruk9BvKJWMWUFeoIAGl1JgXWFfcgg1XfylgddZyGz6rpuHZ3ma6F/iaQSawRQa
jVphLAeZi/cEOdQX2gMPIUD3BYrlMkpCSb3sPnc0Y7J6fqvb36ZB4pwBooZST44YyeF1wOs1tvng
+kTZy27reh0TY4YwCy0T3NPYFhG8M5s+c7BduFB8IWVq1eWvWGOFS3dGDVt0qaTQX0vdomVa+Uf9
XUKWTsduVCq0UVU2un5TpW9HhKRd4gCBILXM9A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
/Otq4ATIazCpFqgShmqh2TQPDS3Zl2U/bLtlOvCZuOWx91YTj+qhmfI+yCSKCbUk1KTiamGbEqLZ
sT01CVvRrD1yO2fLxjSicUry0GLtUfZKdfS5P29j1e5G33aVa3y4wafU/s4CsOhdgPyfrASZ5kL1
zxz0kV4V2SgK8J6XS3kXI80/LdqvDNoiBGQfFDdVYvteM+ad6xjombATlwnei+WMIYDfWY9WS3SS
cpKc5ZFH9KDR0FKKE4imTR034rOu5h+WXWXPVK2VaLIN3PZkjRnM+b8a5WhKcWMeGiy4Z+FofyZp
FeNOcGnSvXgUwGnK9tELYlIghgX0NBPzhv0oRYtI0cBE5WFhnaCciTl8FpajufuCIzCFTMu7Amkz
qO1lAidYJipFlAhHz/AhLrWy2kYvOPCBeX7pi/amp5FvsoeVM8pmzQpjJFn/YkAcNbc196JisWIK
4zu/sHIqeJSg7dSmrnZOTcVBsk/PtlaJzO053aZEFfl/8dDWpf48ituG3OsRa2gMB57hZOCZ7LTc
0Py0Nlhf4Qncsiw3S5fUOneHEp0kz+RElJTPt7UoUSa1yduStynF3PUZ4qwdueNbmxGZAFJCKdq2
b+YiCfxyMoi36uZ5JogKjyCk1NbvqETARHPeqsHVtPSeLvcjOo6eoi+9eZNGby5a+kA6MIN0lnk9
At1oGk+dPguHwBhXDYaetdJu6l5Ckrrg2tReKIlgkCcaVu3GtteI4Ku+ehs1R4h8aMh8EGmR+o3k
aX6Mk6IohXTagBXUrbdBq9dkugLnea0WU3UR2DQH4dDK2F3f54LQ06S1aiL3pyc10Q3zVtzHjzgg
Z1iwlk38wf0O30sVs+PmamvJ1jyVwFc7tR+HsdKQ0Cmjk9QSZUjqgtyp0GG0bbbJiYmH/6UkHFQi
tzlDCBu0/wVipMHVfqX2Mc9tb7tDt3LhOKSZdypWxPwvaLl5xv6DmCnGd9bUWbuvfFo8c0zlnusq
XzRTiQIRY26LuZUMrmLcmciI5HDnwcPNQC4Ojyopx24CFnyFn93p27X6EB+9OtXdrt3hZ53WjA8e
5stUSbJtKigxCZsqxTUnvfiv3UbVuNpXRw0ObFU3NKdK70NI9SGEiKYtq21JwKIfBcpi4DB+bqFl
gRbhUWuZN+cSEUmwESvI06+YfMDB06mIu5GBzMiO1SOrMZrB/y2w3TL4NZLeBCDeZGFgl8x86I2M
8oHeJZ7M5WJWwk9ZO6xwgE4Ik341AAtV2at5I8SYVN+6qphr1EkiIBUkASd3/dA+Z5Nsr/+tB8g1
g5Xdv+69xXvAaITu4Y2zq7G4uiO3KH6ICuUGay1tKSThIDzLodc3KrpjXo7xChBTgcOGyFtk82s8
zuIOy6aXi2DqT+bFPkLNwgmfBu06CyZ5QIGSmpg3JJYTkF+8J9zo/8BRIfi+UaET9nP/s9oKfd7s
xoNtfmE8BLUaiUSZy145+57k305o9Ye1elqGyNQjCKeXibQ4s6v5o+NwkQE5zvFXQBWApvCRwywB
uQ2Duw5yIbOKutQEf1gfJQE9d3+7G08dEh/XPA8TFPhQGo6nMu3oa9F6KIbqFFVN3oLVHVBxZnxP
19O35hNEAtZjorP2tVnlhMMUnLvc1UvEGA9uy2hizJe1MI/eonT8xoQykQ4NOFi4GZF51usKAerl
YnVbUnwj1ea3hurnr183R6hEgSOY/ZmDVkSBPujmnOOzAVglQHJKnevqZmAtU/LgShyqRbzMiN2v
0HELbvpWuvWCi/89OwT5ezL7k2S9ozp8Cp0mefmEqoJeF6Y/NfTvR7cWkTFYu2+UrcqAocbbR8Vo
q1UHUPc+O4em1C2xzoUwwvbvkG5loYsIleLlvk+CeZT0Q6xJCkZmTZmDrC8IDryLR1DQyqsDbOtS
o2yPfDJtR1FWlS3qsB1X2Jo4/2NTlvTs8FMEeelX/t/Wkl05hdlD9hAYn3JEFs1PDh8MFT+LIVfk
v6Q9Fvs2fGmxICgVswLSZEgTSrNHsnx98Ig6ZwZnruhC+LmKHEK33DfkNxzKXfmbazCSbfJxKtPx
uEYFm7EoemTdPfGuDSjz+uRPYMGK/1BhqEf/vSd2UNeVyRAF0SJW7pWS3POYffYarDDm+3zkNmcl
DbJXM468BKrY+r+aRAKw5fnfitILSdEZDwSslFhuknEcjyo02QsLHeYmy2ZHI2HuxIafWMY9AyV8
i+X73xR2c529+rGwc/xHpSy2PdYVBKZrJBskl8xnLiiixF/IA0MYnI8ZFFF5qivQcnP+MAMVoG3G
xs5razgkIhic+RhKaLv8LfDk4ghrb8RVGM/SwUFKmk4DBKSv7ulob2ys7hq5k23o2NtCh5Uuywfj
YIPZ+dWUtg0N3zpts/nM04Vvw2u7FuJgo8zeM4HAICVyMQWkcqnlzR628fT7ZybiI+6AD5yc7jrD
yYbQrbwTuw/kb4jP85hI1h1l0IxEMveh+2Hf6cn7Ae1yBC4wJnTOF8N1A0HWmWc/WCW8j0Ip01iv
LPOikJ8xjL55cq9qbp8Ru7djMZ233GVtv/UzVQXOK12wuffQDJ7PkzsQNKWHOuHJwdL0TjhvFaOG
tnOS4ix/AXNUXKPOQ5utrgSJ+iTkjq7GLKf7tO9L3j/G0Q6j8u/CgeL0IgoTOPjSs9mw0LQiZI6R
uNM9ZdO7sT9if760mYg/FmxwUoqLqe+YsxPLyIq11SsX38hPrPw5peFabBg/tOYT4SXIQdGtvkDW
PGLZToQ9in3q+XrJIH+Y21o8anjsmU3aFKRHi72yNvNNb16RVd6KlCAdvVJCEw+oAYyP5YddsBXr
ToY3NatM+/nbb1w5F7qxnRHPvWd/9ljHOF+kTaET/gQFJssNSOWJYal9Sytvbuw7MQqb0iCy/6Ya
ejeQ5sFIxvfO9iGXmYrrcq24eOAlVUWNsG+CqS05Pbk8rSufbjn+tPWqLk0SjjhR5ouk4nRBxVau
GnZwUSu+tnJmNvCLRklFd2UB5OJOUp51HMiIU4/trWQJQdBhHlpUZbRhiMsZZ1iQvGW2WNblomTv
v6vEs+xiY2g5F6pNN7/W6iYuI6OaeE+9hdcasvc9L4uH2ncHeQcd3MnktacmGR9fMquyBGpbXYdW
QPd9vKokQlMTnFI4LYBAfTxHZMaQfgkhuFXksXbukqYWvydVA8bFvBAAHG0858fZCV4zh32uVYVC
8Uab/8Uu3EIaiO2W2o2csjAXUO4FcgEMsjJet69jil0XdnblcNSQJLBzLLGfPW8MqU9A2+Z6cwJ+
YskyHRbYoCzP2Xkrv7NM+xoDlRdPwG2UuA4Pxl2pqxCQVYT4XqmkmVtKmwh6HO0qNVxQj3KIOQDI
KCRwUJcqiSKS+KyYvuFzuhQ+g+K++1HFdkdtPeHBOvboZOi16yC+VLLXrUWP4s7FiEPow5YEy6YJ
Ot/LSVXYUYgNv4ydlTFd+IFdH6GJIwtbGxswLOAvzub2SEa+6NxSMLTYyXMldPfTq8ScaN2xvXYq
IeOtCaSPevtY/laPty2afmIXAfo4Yd0lUAHTeCrj9lxI57fO9bb3rnpj3Sid9CHWKM8mYRn8SAlQ
jWJ5P+mzAUwrQtipSNihriAuFahoR+4EjbtDBFEu/fSpkgeQtYFMhqinPZ8+wB7jAD4/NgT0qsvD
c47c0eKTonvuCEMZ0UzaobPRlGKE/rg0lKLFfIAg6k2KPaNWzK9DyxXm9mq0LhGGlam/L+KmiC8m
oUiv4ytx+BqtzO/38nZ87SE9BZZPg5Te+wWkkbOZXQk/ZsILLrjAe+pH0tLp03BPH/zn5oRt3HtT
ilhrVv1c9Zy3rGGDUt3CVyElsCMDEzpx5J2ArdX69ZdjpYFz1KsG+YQWKXz0NB4F2Ksb5uRhgZjA
XVGuDnp2V3EV9deEc3yH4jSfrULcX70yCzGmq6cm/ih1SUFcSF1a4GORZB/8VMiBcjBxTNvLgtg4
/K/kPdeOHyJ0VlV5n2Zz8RpEaKjs2XRrQ9vOJt/1WOaBOuRPbBmrcj5GPj7+pPpVohcq5RenBfS9
gW8fwSc/0UUks4ioqPZZpkoI76nVc+XuZLkx4xGh6WWrJMWABHxDHnortqFVnGMrVJ56yetKpmu/
zYCvAhgDmjKvnefMae0+NZ3JY1fPtYbOJUkJycjSRd4FaTsTkS9bOY36KuFSK3DR+yWfR9/WVL0J
P5Q8sswkgL6bxmuRhueJhJRIQpFQ35c92wgkoGOynGVaXHKouqivkoWli845ep7fHqAKconHHrAA
bnn+sqaauq/c82F5xCpfigZMN0ur4GiRrlHvbjpPf9rwWjnJ4x2qWsGpoGKASNvJec4msAfupos9
SUP+AZQ+/rnLhbhhGecQqk3e6e6VeVIo33o+1TWQPUryDHmrrYxIzBTGims5V4O29fygBT7N9hul
LMufJySbj9AneHh8UVtP3j+TDaGxMHDcW0hT+aCKXrAaVtBn/z27TZglRsvqFfovS5PPCdYS4vXP
Q6OXvJ5BU+S3MU1ktOHXfFM7PzwHOYJ6Bo4zAimdBsYQhfCgK3EthpKmBhPwjK9vpi+nsJbEzWht
/bZ2xL8B1VVQNU+aKSPP6rbQonxQE5KrBcH4Lgoz7qfeAcwR+5caz1ztGyy36fEbNLNX0aR9WKB1
3cxik7pM2zw7HkfrzgsvFX8/c9eMRuynPrP4IxjJdQBQhLt7g2Bkn1/ZExsyJVy6QG9ee1nnZJYf
kW5wnHcMTbtDrkI5fDfi4Oz6zm2LqLV8SJSl3jJlOBEcOB9xRAU15CtL2fST8Dx/afEG6KozNHj6
TbZZ9YH711nLELdlNityvC2yllaQzeUYz3WlgfBgMHkE9Eaban36VwE/oyQG1qhwpHlMUTzWiPLo
Pw2gQyrdw34mlZHx0aIqvqcgAX1p49F6Ve1yohI9ByEkPLY94E29Np2ivQftPkCUJdExx3ALU/cC
f27tV5xzseryQ5qvJlmTSOCNBdsPdW7LmCTmJbqNXINFnHRjmqADECmfYqOechYeQS5+bb1LFUes
M1t+NgqN0LCHR0h7FqvmRtKkYM2QpBAWppIgnzHiPmDHGK7CMLimxU5Yyb91mS1SLBMesuRPf1JM
Ocje1gYL8+1CLnV7sDJSG6ixwtv/WDp6xxosvnUFjxUrDfGmbwYQT18fMIzC395Xcc0bUHS9S4r4
C3m4ZttMaQ+o1iMXVgwkldN70yOqQN7ARtbA+i67jkwweIYt1aPNmvl2sk3N/4hn0MCgwUMXRd4z
v00vjrwi56OZTY4jkcC/i01kz8EDEvI3xf46qslm8807kfdD3Fg4Q618qJW71djsu65aSdi6GKVy
JgAw4UC6ONFg0mnTG+Q2tounWmMapUJu6hTu2yZyp57O6CV6P+skDRyKTLjYfeNtuub6lXZbaaQn
Q2BtR+yjy/aV//wCTXi3flGP58v29XenPOKHFe1LcJNLDbsUIfhh4WCBnRAOvN8s8rlIYGXV2dVl
W75tTAtxACFUSCfE4lQqJWtDvIJOZ2fNLSjlWG7DEN/mIJ6Twv7w9oArQ43JAjX2GbDCf+i2zWjX
WZjTcynhdoGpNzkEXq9I60tkoHajvmxjWmCIx7hQIQxnyUZwokrbH0MgeXIjA/qmZ2Ofrpg40KtD
z8+khRBveCcK+ikO9O+KXlKMw6thmTLkAjbBbHZlBdyK76Dxb67DqjCE7RbXzw01iSCSZOxM55+r
WntLZwYuVQjQdPX2BDoJPCQr87cjyUchQw+Cbp6R9DedR8QumA6bGwunh4VLYkpVKU6eyBjiN/gz
WFd9l8a3Q9VU/8FdTwHjLJirlqoCR+0AcedwXCAEIco1aCj8ACHvNxvBc466brXsG0VVSDyE+Iyl
ZdGE1o7pEjs012Ma6l6X3fsKGfVyitx47owcEIEzDdSl0QK+eShLVjGJjq2hbpFaE4ynUGhHcT2x
6fNohWiGo7vCsMbgnsxyz9ZwJFzar3CAt7MAQ+7uh23wyNzf7gcEACvB2rW7kuE4mAGxWOd6BNut
oe+1w9xKveBJOsBhqJVMiHkQ47ZbBUH5ZyzXh/95LWKcYt6Vxz4oq5S9ABYFR+kaOYetcN1HbxFI
n8Y0BBoKhwHGcqkpUurmBlUZ2twygC2MkHlI2zw2HPodZNKCgkLgxRHTwB5f1L3SX46oBRHuVBrW
hrclUkLnq/ruVlRGzvieGWrTyQmM/u7+3gudLT+1GHaBv0PD+l+bxClNR84yEDWX/bjbJWeFy35E
2d8tf2Hol4GQudtvcQ5Ld4GJaygW4a6gLEOigez3EhXWltHcgf2WbtOTRFaR2wtDbjwZHHQivkeX
qHtX3JkDleWqhYRe6vB9c8fODqw0gLvZJHRy1UCQhQYLp/sl4LzNDOwcWy0TLxpZPRU0diVMfvFX
jwsPuS3uMMkani2ikW7nsvbET5iwMMyPJpghM3UP3px7nvTcY0zEfjZaMnyNzSy4T5EFCbq6Jt5L
M1kNr9luCJOvGx2k+sUwKaAKPYtLDLtMfNmdx+hHfm7JPsnyJuGGLpOb2bj9H9AB78NaUhosMN/W
xjJT1yNTJy44Rjf6r47uxdeyBREFplI6H5JKS1I/Ulw3jWW+YVIFgZ7p5EgTbUieYSzX0pJRsiY5
JSP5L7ty6cS1tqiWqBvcXK/+KqBEcxiM3Y5wU9SR3BxeEyGEtVuJxsdadFXdj3ObUoaRFvvzFR+w
aEXC4xGhjjiFsGnBQ4aXNCg70APFp+bKlGtEVWn1fL+E0ZMe65xOUZUgRkmUbLyc5r6FI/xlWRHy
PYkG4sPb1FSyo2i3nXyyp/8ANESfst8QdMm9ymcEvR+BzYbuGwBgKuaPItl/jYUQRuPKeH7uCgnu
9frFpGKXfezfI+DNqG2zt25UN+z4EEMLQ1gm8tHdctGlmhFyCs6zBQDKbz6r1WXkB90vkySZ/JAO
gk/gHyJrNFXwtxM0+LZIz5r0TZ7PEQFjnug3wTTjPDdXwfdPBx/4ed3TFG25S4qgNQhIOouRJLmF
ppey1LAT+74FMzzvtCiwx7FUW5kggGKkaJB22C3Q9BGWDWuZ87zAdcF3lRFJI7rM8FtVfUkkcd8l
dwMHV2m2UrOeTLawIJ7h+Ie7pjoFb8Awx1hEsTHltVG9BM1JDZ8NSNe9784Oxs94vW9hCOEXyW3Z
b1bQX0NjqNpz/g437J0OINTsFK67hZ4Z8Fw5clNuuXBhm5BowgotOVSQA0AGuMqsbmgAeNigygYZ
DrUSbSkED+C6OqLBIJBEGFOcwkRukv1y7cP3bnrAFyVekC9I8uL2ymZh4N5MMJdxC1FfxSuUUcHA
TnW+zR2Cjn/qjFzZg9KELmKSeUihRoqinriGRgOD7ybYXSJiOtyQM19tELaQyus54jHshL/UJw9f
UNjJqBkA8Ygw/8Wg4v0CZXiLiR7UnhTQ+XKo+2YI+gcIsLUfVuEk5uXLf0Mv1ZQttF+Z7XKnfFir
aZ+IjTOdoKWgkIOeW2AJx/n1im1C/R45X99GgQNnwHhfJKB85+TWKySjYhDsHJs0ZGyHrbb99Cpp
2QK9CL3QO6nv9wVnr4XDctFhVnftK8jvPjSpVt0g3pGOvAFdiHv/U6cuVSAFI9tRL621oA4pz1Iv
D1efLuqD1TjNUb9GwZiEz0Mc+pmXHU0uyWwdAhn/bil8j4VOS9a6PrS0Ry+kVmtDYOjyuQl/HpEd
FUfY4jCpCicETC3dHvFx95/w9SZfuXd9Jtqpx/vqKFrulyeHUWWwvn47uy+ta4e7uNiSXZDjtqUU
Jsdhb68J6+o283K3zz+Ejy0GlNzJm6CSVD5vSFQI9PCnK2CN9+lWe5Vssq8hVMh/r8DLbbUuumOA
Zug4L11yz1Qu4QbTtPaFgrp4hqAHNnx1zY0iEbf889gcp/tWUmduLnKjBSJ6cCMEtLD5uCzufFUz
AL4iL/2dQoRrIsM6H3DAQdp3R2H3blAyqfpOOLMU3gHqQjaWf920UzREfHbow6+nCwQbfU5bewSZ
vAj0UTZWtEf89mPp+UN2TH+dKkHlAkp01qyZb7ZToILRyIRFzeu/tu+/rM8wtmWl47fCP7Zub81/
1P9IpwQrBfarHWzBZwBe8K5b0GxsNOTAvQ4YwcOYxBkzE13f5qEThfnzs8K0x4bqskl1to7aCkn1
4/Cta6rGm3IePoS37w==
`pragma protect end_protected
