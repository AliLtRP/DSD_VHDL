// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nXz0uvaSOB7azszzCjxK3mnnbXoeMIZ1yyMePl8XsJ0manLADdJ67LkMSpFEMJ4w
xU+mhg1aFwMcuzs12kv8ZKRNGHtP83JgQJjwHCrTr3sQ6nbP0AvohLvn7XYsFEoU
QoaroiW6pNfUEZ8Q/t+P6v+gy0BmpcGsjvKqAln8QF4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19584)
04qPGExE+6VRv4XTgQLZdyzkV7jn492vGtbiQGitQI7gP7cS5jgiIiqz6L9R2xqK
oaNIvITrLQjA1hHjhTwnhNUL4TkwK5Q9epcX5k/O2DCnB5T7vU0fEOTsDmrWWavQ
GYlBFBHPd8e2Xeuqlw2MOUvTRuB+9gHlaPznRcRaUpCc+FpWtMkjkTkH/y6pbsxF
7J2qBT+xw4h4cIGQ16GluAEzWWSxlBLJb7AccRjj0t0XmZoeaXo6H82ksT10NSmC
cmcMAU3c+vkmkEZEtTe4+tBaHFJu/Yby4FLQG+wnlnbtAwC0TBJvp7jrA1+1sz8p
IaP7BQ+jaUwDreI3kLpGTFF8I8UVgs8S6mENhkqs9vYy3DvW9Il9GwGR4rupgopb
rbU3EACSBWOpggfdnrIIruSfU4AYszKz3a29k5mEig3DV9Oy7NwF73ibIHKP7JVw
9iuZcR2ytb+AbA6ycPXsniXJb7aNMJambOIIAwfSeBA96QTNifgikfWSnpkKXwnj
qDoCIFMmQvgZMSRKppcdBkneGT8jojTISH+sIMoDA74eJB2Sb4nR6U1ihIt1mKJR
kxRPBnZEiuX8Q/96qGKvWCX7KpB0E0iGXVp/jrFFLPoyEaquL1S00j/RqYpENspx
HjyQ7uRPsx/B1xnmPxHlHqARr1oa7Ns0LvPePca9FdocbHkngob687TpgDHkGi13
dgsUhGrBDf8zcIo0Y113hXUwCcW6ig5+KjKG/cc0G/pxiB72Oj1XzalsV0eXSqfM
6TAmqmckg133De5UpjrgbbCvbJpDbruetzyTKXoLN6/Pt3hjpd1opz/vhrzdb2Y7
E9cxwpAoN6wC1KM5F5VJvEJhti5UUc7/+WN77FNeRyhc9/W5DopbHj9GiI4UNgOv
cVZwnEkNI5jEyELfmCFPNU3OlMX2tWCMVmL0Vm11geOYLwefJ9EEG+btSzuQqqeH
z+e9gskyWco0K3fEunVLX7qYMEMdEeFyhNWOUOQvvTYw86lXmpJ48e7J110trHhf
1AtCN0R/9tYQPs1Ox7amCceLBugcA3cLF6aQw6+2h2WaZ57KHRhYTj5xOfpRbgr1
7pNhL1RhL3VNHiuFEsZcvhWhvdGRQlc6nkyKsOMbKc6GWSaHMUUNusH+DweaTJ+v
mmpHizu98luHiKmN1QPDEltc+IhVu5jpAVqiceu/LtgJvwotcwv6NjUi9Fk/sBoQ
ICgOu1dej7Ae+Vs0nfbj1F9Lr3hjRb+g+O1fm3qDTdWuh07BglGh9B7wHzfIbR6b
F2/ufT/hUWRTUHXpkdWFEZpdKmOuDMEN3b3IJj2ifCON2j5JsIgkZZXeiC5wDO+k
C79mIelI/YdnsgCVf8cI8eFQPJZ+MupLnay0R4av/PgNDQU1nDsvbnBHTuVxlLh1
hVIt88cFZunvpqN+j3J+gyEbj58FYkJctFxbpABr/lccN2wcQak1R4+P4ImkTqk3
CPULlGN1ChjSuGMp6eWLDSlcsR9OcRLU+T3DdxG2U0NYv55KY+6LbJZ3YbPGSEqz
5w8/o/Q+t4CXu3Vx1jmPzmwXRbO/CxCdQS05zugCopdXMIiJ6GouUd06MUFSpXWu
4NvVOns4wgr4P3h8/eMKRi0Sfr5FdhLVuzwPovwMM5d8O38H9ksTeXVIHPAUB0hc
vkpvgmOfrol0tXyfJX/gU0JoWZoddFJuysuGFt4Z9mf6skooeDU0BY6ZEHqk6EDe
cCetG/4shOMIFLN0f1ofk9MWEmkULlZpjtrS9DfrW4DqyBK4DakWVBJzEMxZxgpZ
KIIv20/Q0+pueBn2XU6P0U4XN6jbfO085GDaTp+Vdq7OUvWlglQuwDRiKgXgUi2f
B7/+t1qHVLmH3alIltneSi4rHQwUTCwxelE1Tvbr5qvEOB1a5Ho/55JFRX4FEk/g
7uwjAK+0uKx/WCuYIdkdmkZQjLRX77oAdW8xP1icqe5rKcSpltK+bjjDehP6G0jQ
aLznOVpMdzPTXyZvgG86h9tEzPTaCYVxG2rwftJwKsMt+w3QyTvXH3zYHPhJ7qxj
UHQUo83qjQbuWipFGosNrctYt1q/2C4NDsfjuGFyEZeTEh3sxxCDsAWveq2+cItq
32vJNmcR8JSf/pgrfTQV6gF/Bc7R+hJNxSp/oP3Fl/AFI4JgO+P6q9voFYowgfnw
pNq8ofOuxKWJFEps8T3TwI6g6M7txqCcwZHJWNvPbFLLtyp8GNgBPCS1A/Qrepoj
E5+zEYPBci67pHkUgKNR6pqWtXQH4X1lfr1ztaUpmVfErOtFe76YjYKK/eG9uiD9
KFJbB2faeqo+zacXt/ckFPHsV9Q+oTnXcvHNFRYxDD/JtavKXcoQsjjTErAl+J9P
lSSjkgYPj0nSMgiTubBkUtpLp40TlqoSbCyaGgXXPS+ST8NB1tqu14SHCGTD+ihe
MzeOPIexDEGV2rY+r6qDZpVFB2BsKRwNeGVvdXupNb+cVYm/FDgqpWyIb9XvqSVz
/0sy1z0sZD9MVrwKjiJZ7IPLAJSXN6zPUeRY903k24bQ5+uwCm1jgH/QemK6SzBT
6EjJkp8H5HAvnVEeaLjQr86k16vcn9HsThHaIQR38xqSelHQUMsZfVAXSATxqVVV
i1ibDYi+76Exea/Qojy5TeBiq+R37diErTFI1iTbP+Bp2tnl350sIx6p3rcdvzsX
0ALsg5Vix7+KUO+eg46ZDRLFFIKPa0npoc8ed1hBxPliDreICuihG2MGoezmCITP
2YZD+JodoRh4YRDZmSLvW+GZBdxWFWsDEzDS4eVDrqpYYG5nwW77j4TIu1VAT7bv
sv3T59oyKzdiqCdIW3GN8eE0WeP0fkbD8YUSJTO98Qf7hfLtNugf+gsAnTuLUpKk
LqtZPNHkPJVDcgS+pfLHDgL6Ir5fZ4nkilgbBH4vMrKko4ESm/U3qX1HvE8fBk5t
Pb6+3XZmKLStwhDrZa/9L+nqN4qruH2e4vhYdBfOPWKLPDtmcT0rbtHS81S0YTk7
aPCAAUeCtzsK+pTAos3G+hDRjgjFZpzOt4VAUn56NMXIakU4+3zNIk03rYt4+lSE
4WWS1NnP2vfnScLUBGn8QJj5NpGBeoflM2Q6pRE5UQMufmO1OPc16Llb+IYODSHT
oNlqk37XIG9eB+tXHqjlk7VTwghcXQOEQCjBdK56swDju5iO5Yk8ZOAYPRljksTx
q7EV4qgEMHwB0RFZEvb6U4nJQcwTOZMk2tNxCJUxO9CUxKumGoOp3gpZ3BpVmV+B
thTSGKPYZDhjv+P2w7067A4f03IsOpZIRuVGHFjxi8k1PPWGHehb6zbDV8D/VXN0
ALBQllvw3l4YtcvKD2M16oh5aInbpmZ0BLw9FfQCJRYxiy4F1E1NjLEnAjOUtBar
CXl+09Rl0Ybx5+jHhIGQZ2XVelCxK8d5nzbKz1WUTLrYDHWULtl2Zi/v6ioxpr9p
Lvb/sddS8e1Wyke7CbLNmEHF3FgXydoUUUsXbm7/nq2Nb//EDUpDTRMs/dzV8o1S
flghkr0VZil5AMwIlQgnWzHX1KRyr9DnOkIpc2z+0/9xu7eOwfTr90u4uoEjtIjc
C7cgh0YvkP5ECz7e4xtoTEGnNaZNpHPh/+Q85+4/zvryEeWHQa6GmmlH/rXS/WOm
TVPdqfZcQLZgWpbOU5AsU9S+R0d9mL8ssS07w1CWIEFXgH0MR2ohpb2oR8YxqI0W
rvU+Yt3AEIdBooN6ZoRK5NxuJ0Pse+CVjAJKN2JzH+ukb6sHBdCUXbwRH/UGY4n+
ZIEIAgeT9GpGrFOgOsD2LslSJs6Uns7gE77s/Bb38yxosMDUtbQ+ClXcR99eGRt7
zV33ulcLcCQBznoif7AxeRS1Fy/HIOCoJdW3LY5dundreXKNiLli4JYNlrQ79S83
3SRPFThEdAOyCWY+w6TtP+buAJ5GSqzPoMieetD5LGReJs8qcTaGb44KbIsRoQKZ
TXvTIlu6I3BNSV76b3JRwF3wNouC9y4R57HZZJsc5mJtDai2zbIgTP9WZPIO/QH/
K6xXvQbxmB3zw+htXK9lKgm/DMFqkye4ZkHtSSZx35YWz1VM3LwEcNOpQaCi/wEY
BolMaoi8u8N3ZPjDKvMPfEZCeSkLIPDTIj513+7+BfIeAkuvdbWczrji6UHEOCnu
H1/XKDEetJBW5hx0OJ/t5kISVt7FeMRDKonId6r725BcMYPoZ9ZLXAYuSj76rBHU
KblxdSlFpFo/GDh3CxN2fmFd7R7TWxzgNAoK+Wb+0Rk18b4wFGDCjzP2x2RoX72h
JRkYDPrdBEpn5FCBCAEVA59SMqndl8gsQFx/oiUNCditj8WInIb8+xmzE3uDfUlB
MDWdjoqkrJ58qG127Mmt+EgQxe1eo0MYu2XLsGW7TxY3pKiBagi/t0wjRNbf/Yxz
Sk3TJAN+BlCI3yJtCSUNvv4HNrBkS3yMo/o+Xw0sryfKMhxv85X6DnW6mG0TJ9zE
pT0iYNAmOR9rLpY7i2oY9GeIsUZ9QI4EAsfDEMzZWX/0MCoIJ2c63VCVqv4OBPbG
DZfPE5pneNgv/ud7p92u+zHgjY7I5rzDhZzElFWrvA5MsoUkbQc+e5lvnQkTN4gX
quCsD02T6CLJo/oEiugPEP0ipqYPM+fnKj3VFYh2AI2Ab06LR4m/X3i34nOmEk3U
ObGpKv/viKf/JfYnUrqPhnFYnYJ0x7GV2XIazs07IaSVv9BZ9Sv+gXgssa8wVJUA
cJ2wkIPPcdQwsyAP+IjGBmFN9J42FJzP0JRFj98kwC1l6v0TvCBD2pBJG1+fVoqC
gcmfBK+zLhXE+4JBT7cWqQQYb09/i5gDhRMW0cGmo/Nm1upF6VzsSPF//cOCX6XO
D38W0rHKtPna//sBzfuDgEOPzg3+kpxIOhedSvpEY1fqw1kjmptG/La5OcOXaiIv
Jk5YkQIFHIomWacxbjbu4Ce45H0+0U8uMTsY48qBohCE2lDFgDTjq7P8n9DnCPCo
8V1Fz+YuvrDEtqM7UPr/EURoJJ5zBI/7Hd3xnncQuGcM3C/jdAef/yKnJC0gRJL5
ncKoPvcniAgiK2BmuN8pV3y88AtidarQo1zyvyE9bmV8y7KGhhWy8uEtE6FP0TyX
umB9NgHo2UhYOgKU4PKBFGCVa/OeL0jPA2BlUatB2FWQEv2aJhzu+OK2PVO6WG3d
Yt+TGQz1m7SgS81tCl1JBpMjq4icYXN77DNDq6CiskenS7U0UR8s/CQ9FZW+td3I
hXCnacW4VUSxoHxfxPA2OWAUgV5psFpFYtjYRfyQPVeYx8/29U5Upb00h+0E2Vc2
ZeYxEWWi53woDfvkEPOOwiKbPDG7wycDdLA+0HKHlWhhf54FYSZMrfNfjjVzZf1n
nAgftweJfFYs1UHv2bmXCY8ZRTHUUwWagPU3WN2gwV/3dd9ISzAX5weGE9EUc3Sc
K6griHdPFfX26z4KQlKWhVhFHwVOTudUdfERiaaf7NT8px+kNVSmiJ94KO/XtqYE
CRh2bT0ZnhpDkUJZIuWc0cWsZ9Ze47r01fM1+U9hWNXMjPa3xf/ye4pnCDPaJd3A
RWmXJ4urIUanYm4ne4OqFJU/bPvsM2uRpw57KVYqQ7FMjnvjdeD6pp4XzQTYDfxq
/1ttjcXueuCvKAAuRqdTrdj4/Xsf0Fh+hPptzpjJO8rYrQ0aTMEmBz07bYUkCghs
Rgb5zlDEOOXQWQYWCWBVj5nb/abBft9sFb2gBK3wv1ateSwniSS/TTeCax5nTNAZ
QxD0rARXpxLJAWV9KyWAhGEY8z0k0Obf/8H24sdhtK8REUNUcj5huzZTHtkQ4dtf
gDPgslJFTedWp5/DIldvDGRTSkJ6g6RG+LfJwOli9LcOl6258m7maOpgqTs4BGKu
mAkcvN59boq/GOOZAfqFPfWKyWFgucQV1ovy0oAWQ2AzbD4lMOLwecCdZSflYk/5
GwJTLsqiYd7gFG7t7TBUxNAbvrZg4F2zdD33sqiVT7Ff1xxYaPEFItLyMojXtWuX
E+w97K8m1EZyS36JDYZ39/INJx6IvJeZi/OBHPcU5fWsg3RSHxkufCF93Sud35mh
Q+Y2L/nZZdHpC3FQZvIDo8GcNOHn8/k0+YfypQEErDYjXRKCGdKtS2JQjBcS0+LZ
lULbMHYpqLO21Gd+HVYVbdfkmNYBfb1L5ItnEXrUlhXhgxkDJ6m4P6BJJngwIGDO
6iwIe7rAsXb0wAul2GKMzbHWLA48fDJYFo9tfyvlkoPcDp6/XjBv6yA5qHNuzAYY
8gFq0wydSEDZUsBeOrpY5SzhSMBHMhcQ30Bzo5edgMY0Yvphd4Yz5SLJrw3zeUCI
pkO4h2JhEmY8F67jsJOsv76luVmE0uW2ws1iw+0vVdCIsPUnoz4d0sAGuCDwCMQS
6XPyiJ5QeAxa2zP7SoqvX8GTHhsbJhWI1PafKZvceMsVkUr6HYIW/erP0FakU8Hr
eca/uyWtCC4J3gKOR0sO9ENXTw9eLqzQHOokd8cUyO65m6emPQ8MQ9FGncnNDRIG
T2fDy/JbiJ1LS7JS+Iv7jzPf1rRCMpLJjYquNiE2c1SBO5Sk+EHbkDK5AiqqI9Ps
Fuw4hc14HB7EphXYzYkr5dO3H/3pEU/+mUQxEHIdWlXPeJGaJjT5psFKz1va8y5i
jILE4zNFS5Wr/6YXyNoJ6HKvz+VNM1doMpjfZnf/RDbKGDn8dt2xEvNxeRRt/Wkt
rGNchkK/FDdKaQOIcbWWbE+fFF+Umrd1ZnL37mVWcjuijr2tK0D8Am7cktFhdp5H
8Igw4It3pR6cPqFGbhqYKo5eB8S5Al2oK3bEJJ1BgCR7MEEcyutH2EK42MeTcQ2u
UYxbFgID4Zjk3tBAOYCvo89H1ugOpvEz51fi3GIwhpWyQlv48yn68UQZ/glpUK5u
07STwKOSbiu85m3+K8Zj0/+n12b0pyBV4cfXB/hciFcpBAZ6gchQ8jwOzxNFhYna
2HLmSkqTYsFIsr/XVLpRXPWIyBkBU+eoMJKOXKOVb3D3xgjG7HHYHUZp+nhgW136
EvnuJckLQb4Cjjvoig2ab5N7QkgHIi/D/BC/iwIPE2W8fUYoMKM7zCrgIXxcCD0Y
FrpfiqtPcMMDNGHdnqISmmMJnEDC8sWX7qvelLsc1Pgi9D+KDjxCpB04HygO125Y
TdCXdp213jEfLv5a31Jw3qPdd4vl44dwN4Txf80Bb90++rUM0hniUza7SEcfyVtK
vUy1mvW5XJz+G5Y3uXhc6Z1vrsSBjadsM0492ZR65lkdF4sJxlxd+rq76YL6DCuI
xj0tXzTRw2xOTaELR86vuzC22IgoJ6JV7jI5iu05Np2HaY5i3wLfKtQq8Lgh8Psw
xC8mgsaYeB9wkswyxsk3tWHHvpCch1Qp1g9WFp4+vEOOi6Czw8Zi7rjkHhU+AjaO
OfrFCVyCVxZtx3psnpaEVZaUJWr+61YY4txx+yrAXxfy9yzhavtFWM9SywTLMC8A
ju9S+9nTLmN7koS1Z4j57lwiTdTKt/r8QQASqN2Z00IZ4HusDrpWuT/2w4YENArD
j43YiXI5GWzTrJO/RkhoAJtKAWMnY9Hs4bnqQfd2OGwn/rlAPQJ8WuYwakv3ysfy
irchHFjWk4/dQkL1cYWZYVx9MN2OifqtK8EfyaJlAka2BtkJCsZ/1NGz9xtfWND/
930MJJpF9cuqKXF4DMM7flpxre5CeglMU54D0veDfOGZrCCg2lAi3Gt2z9B55yKg
x+rRKYtVRXrAskF1eEuVZ6XF+v9xhIqnzgRLISOZ/GkvNpigbhtbTedurWqZ2UBI
b4fmYrulzxChCQwPHSGaEHxA0xInpUIwBKL/b8d3E+iCgIijX2QTCCpfIvUwycnW
V4tkMMprFxdQm0QxHXwhOxg6kxVZ7wQEKPyDUNPx+Gm5C/n6NxoOn78mJEElmTKZ
HO473lZmy66Ypw5Pa+KW8Ecm5gx3xz3m42+9Kz3sz8bSrejxdGjryblibnrU/sao
2ZdblMnLnPsBMWVIbOP1teuAHxRBANXvq5YiP+cSCp1FcWSH+DyJ6yW7KZL7jkQy
ELFL93l2uNA31Tp371BnSkzP5lnOlM1L5XNnlfAQPrEVpHMCH+ko+4vC3RDdhch7
zpAdKNwrZlt7PwCeSSkD5Dbot14FKShIn6HHKz+Najvw12jH9gk0iiGm3xSXqUNJ
cEsk34Vcii7rOg8BKii4ubSFosWpi+4kH9G9WGpMZghMzBrJnOutDDCqxbvWxc9m
rO0BhVe4vXBgFcTDdY69/9GJyXJTcLRsFUMyGtIXrpVDE3iWgN4ny+iaAKbwu6m4
GfCdVCEfAdWMsY7qvo+9opX4roXMZvPKErK5t6zzQ1Wiy0r2ZkrYHotGciuEpwyw
A9yXOJuAU06rXfqIkNxnSm5DtlgzFEKDp8SIK2+b+qOk1123noLSl3Y3LkmgKOcX
TeR6GQKzqEnWyezzhnmNA6OZ16d4oQc5h/IDTuNuarCKRVC5X0TLW8v1FIkEl5o2
C0+gudV2V3xNm41Jg3KeavGPcCxEDW5vPcDB4YySfIAQDuDKvrcKe+MFo78CU+IW
uBLgaVRXWRuvbe7LUgbACv8Npfi+L7H1XfyYHj0Jfm+/e9xbV2g3eoAXisxwfI6c
1EFVaVMjPX6Ya79jDUzPf0hpHw4n/9BF4HQddFF0fMuyuxJfh+eknZUMDJobQtmM
b0q6jO7bdAik588gMe61d/q/K8PK5TJvJcw7hOZuyoLu1AVx11RtWS6TQaBkmAg2
S4Rmt0AvrXa4djL2Dt5AjLg1wWrNq173spPhT5y/UJiFxVk+VxV6QaIVBeVEBmCT
l1dV8AeBlUkp6bFVaPof5D9aeWJOeNdd2/rWjfj411aQatCT4atzRxXmZPrdHrmz
3PUm9tj31sIoC2CWsLt/AefIVE0jB2boKiW0/V1QEBYZtxHr4wVcTX84S362UxR1
k8/V8XDjft+JLKoM/msOcEM1Ckk9bbjsYwhN/ABk3dDxMKi+UnC/6UmC7+Ii32m0
e10p2lfwrMWKRrHXOSPQ5yL9fBenQmNCu2wp3XiT3Ttgkp+3Ixln7ZoVMeAjU0kI
ZIZ8qDAgvaFHdHwZ5fc5Kli+TJFcI+OKbg4XQfRC+JzI57NTsXOf+UDwRsLeitTk
snczioJfNbRnfg1iN5IsTYt90+xDSwS4HU5prpL40ItApHeLtZ6o+gTYxXwoqdsl
0xWLuXGC1eXz7xZWfsBHImUMAOU4IvPxBNgo31zPuCnYzUizyPJP+qIjmEteY6C/
KTkw8RchoMW+9kPe7AHv6Auei0ZNmkHk8FYjwfH04q2JZ63SyCWTf8CISbTrAC2N
ui5hHdUu3MSuFSzDc4tme0g91Nkvv2ZDN0e9afJUd4mF1GRBLPFdpxsaU+mr4OWs
8LONP7822Ml2ET20/nKxErQcSi8qO4srBJDOWCL9rmmq3CezyYSRfve0nhutIHd5
u8x4ueVTg06m148ngrK8h4rpMf/jmNb9hRe5ZXB7yRfTbgMcq0VtbyR6HqWED5zy
yvg/q9U4LFahFt737Io8lfAUurYscGgrhBHbBS4gEj/eMOp3ov60Oy6W/31kTwSH
u3g/C29WeSrqYyzy1ksL89kSfeBrUz+910UnMJNXoPxcNpk+leQBrByIUoQJmUD/
wObKIIpo+XQSxnlkX5MOo3GNCe11O5oD6AJIkLAOfwtkRTiSct3xbCHiXyH12G/W
Fi3468GRg2ryl5rKzMQPgWyqfbmhP6RTrM4iiT6pZwCaVeQH4D3iNFkPZEpCqhC+
HWHN4sul8GMKE0TVI7mkEEmFL5RaatUnLA7JMUPiJeM+QUZkaeAdfCEc/BKxIaIA
JgrgWJYV6ytcbJ/x43kuIjCRCcx7s0u1WQHjU4BjpazmMR40ir4v3oWHJrxgOoWz
RulCq1/OrKYPbYfzAG63ryr6ZH/c8wY1Hsz3GyGX/auUmH8EOX2rnUTVELSfqNsQ
YOOLAvl9oFP6CE8Ez3jLcNS3NkHP3Qbv+DJlcYWNlkP9iUY8ENtq11BSr7Ovq6fE
eLmjhV9cv6Cd5V56u0rCMpXC4l16qTen5jRAKPWHB2aPXADnywyeyFHDrstYt7dK
oHQ5OVG9Q5iGJ1uaZMhIZj5WlNfY6YShefERmoBRtZQsY98AXYv2YnMhOBe+yMyq
ZbXawwAaaM44p79Kxs+4SGsBPT/sFyXTIVpBoQJAUPDUDUFSzMAI6YGa2zV6drXv
YmVM5i0UOg5QbPK4cavRGLN4XvBfXtoUnynGgr5AkgaBMt7jHpzhtq1HmAMBd6nJ
NDC/J8JwxKTsUG/BcK6ljeF2+EHItSysaj1/oWxIpiiKp6nckJGklF9UZIHZ4Ss+
kRn14m18FpN5s3avzxS8BcQJuGGy8q2LaaAtU1w4RS+t54P0aulX2n2RVbgvcxsx
DsoAIEZ8y3FOrLiSbOCFOftF0wJzFuZp72LO9TByooIorQB6TsdVp4KXZJNOS+eK
elk5Nw2C9i13cTcSZ33SvFCUjqIp3d7AHYC11xPnjNTvQEDH4TUrwHR8oVYPiv6N
M0V3WoorHlcmM02oFoh/h9mV+L851/KzEhMVJu00rp/kqtqoz5bBHCQwvJ9uNYru
2rGHiFr7ImvuKVaOaqm4XUzYstLVsmcOA4963dGyc6VajxSn07SRsRwEu21bDAjU
c5Cpnfr9lzfuIxyiD9MckAaKO+lzO2P11dwGp96Jc39Zw8eqXOvV591gaFM3Ax9f
fy0cV05vP2o6hlMTSw0hje0ZVkzC2EXRFoH4QSp2KN/BRBoJ3KCFqQ/E5cP636II
HZoduRChIKQ5HLi7KKXyb425ADa1oLFlI1QJ+B8HuyZM67TO2znLX03NQH0vJvjz
5pYJV8UYGs8lraSxqwOtHOEmSF2ubT6Kxiudv/LbvyhRlnUK/paGnpFFafj/0DbN
vxZnWCQBIDYRKl+OgeclLbDyPzf4BVgG5PL2mbwpSXjdTZzdMhFyeGkmu1uP+UEG
mFJ9GCsR78QaLyW9HG/k3dLpuhnV+REYEphIKd2kIroZpQcQ7/gYpUGb6Pw0PRTI
dN55nzB0U5PMnlCehXBTh/hlprqjp0f4QEAODRKPz34WS3ku7j+2CHDeXXUHsKvt
iZm79aAiP49DgWbvce+9v7eKLP4ew9hWvO6qfYWkrUbTfSYDG/nb/vpNQYgrO49R
YZYWcQC2VIoPD1yEMAqNs7b3YONtw4NZllAe0/69Xu4ZY0u/pxbSANDyEG1o43u2
b0I+6wzJnMtfL3wmFNBlhQA59s6FYJDuq4rMDypPmn5lUtPjs1DR7LL3uX6VPbgM
eVEeaOkukngbfU9kE7aDfcL5ssFjF45iii6J3r7U+Ir3K9P/4vo+j80qcGViuAru
c6a5FYtQxO5bl11wUHRucol55HDwLCTSW4pXikhdCDdtLSMdSSkQBkb6VNyJ+KXE
7gt0Zz+WoIzRmPm9zHpXho3uQl2E1kbQbuHoE1UMelSDeXlRuIBV78h9XHMtnfeS
DY+UlGyf5A8zgnxeGkZWKEBiaDuKkS3W/g8eTG2EGsX4/fwAA+hLKq5Jk5nokDgu
IFAp0euJj4xHJ5QX8U05ff3NFginwfM/c+0zwmFb9JGjcIxTpNrCjApmSy7B8wLI
Hj9XM4Xhx6wIeR2Lhk41cRDJv/Z4ognTo9fYi4T8fETQgMCYkFdCwM/GoiWl+yao
hIWV18XiKFTUxLSTB4YdpTHJxkyPp2AE0GXyWZwwPCa0B5Z4QSoeMha5Cj5+kWI0
up94CHw/JrTvvUAogbFf/lMtseUd3g4U7fzWyQxdG6/6U0qZ9eOIkQjsoPRl6apr
JZau3thwI03Vn6vBLzImHzXVEQrHjqxh8WMNYFARtYH6aumQUX4heeqsI3WZvekl
Lr3xKsxCMMX2K0yE2GkwKPONoHLd1XGPoSJPZC84yq+7Bk82kW8FNRotqqepdHCF
XIVBMGHFd/CnmX1sRdOGTdZ88J7B9KuS1qpBCTeNO1EORIEdmYF0TVjIUkA76NnI
GSmP40ivhiu8E9YL9jluODdKtI0YkNIliqWZOr+Y8ndpMZ9jvemgvY5qm/AbSpXF
m32iq44hLqjUA6NACJE7ZBVAXJV+pvbkpZklcFYga8a6QbkemvXa/PniAITxDqYQ
bZfoHDX/puepu8qVFjjTnKD3o33SYZ+uvl3gdett7C4Y8+Ktt1VexdTKjPJRQ5FU
8vec+kWnRNxO+4t1bxnNX+o/Ei64RJvxjiJWsoF/ad5A7ezXDq6xZCZB7XH5FvF3
Q0f8mj8yO5tTggnwg9nI7O5GvJoBAT8pNOhHls4Y0Lm0zcLyVyhpgCl6wxdHYUkC
nzuX2i0To3ppkfRcCKv0/SLMu2SQyWwikzS6WZiNwHoR98ESV7Yd8uCPjCF/sHJi
hVa1SyP30NB9bPguVO4V9dfeyasrD4hK0CrzWLcvqIiyYn2quBKz+qKqNDRC8bwt
omp/w4c02UcqK5koasJUyF1oY6UYLvTYB2+eg3v70N1kGnD4ZRo6rxvPZjliBePz
1DDVRMrDbd6NGY3KQ0xGe+W63Zm0kbbDrbVz/oV97X9mIpmNrOOSBrOOCR/hcWYz
U6E6rto4FNxYaF0BS1pby5vnNO8owGtG2s0ds/s6cjTnwfLiSJHVmXy1oMpKzRfE
ckX4qdtGKs+QgrHF2WBAq180jLvmLqTzc581r9VElr8P6fDVdyZIE5JZ4WfxQaEu
zWdFl63z6YajvyRw8vGzSKB5mRo7h3WDoxcQSqNTaNSKn0utQlVhGmajLpAvgE2H
lQcRouYXabQH4fdWYlh9DQB4ugatUZmpjoVEdQbpoaWz44fmhyWg/CZDJGVLwrdv
fqDapLLe92D4LyP1FHCvCFIfDp7F2ckVlf78sfx2A3/hyw4chwCb/UyiuRImUECp
C8P4WQyj1MBvwNzysxbJ0HtytyJsIvgU46e/uGPQEcONor78u/yoC9xCAQSQzkUa
0e1z0A+N5rjHPb1CBNMZ8iX2FB20WsS/Q71DtZMddAXvhQah3/uIBGCTbqfz+xfU
UCQ9tDGKLv5gChNp9fgRJziXqcfLENJKRw4N0xfjkbNdMKJ+HUrkY4DfKPNMtyEk
dOQj3H/STAGy5PSY1ePwAeDy8cUSxDkxfftvIGyZtxcr+Kl7NY1qzdInAbU3BUDd
fTVE8p+34nW2KrSvf1LcrVN9FUz/entP57J/GHHxJxJd5UHOdZTKTYUjlL8czI5y
uOpFBclKgEjJHFVudKjD1+t2sF4xpHoIcCB6s6gbQvLsi4fXL6oRx/DKPIUtWcgE
2oKc0ZP+qKfz+gQEMUWhMTE51mDYrvRR6asq6uvqSN8pMLY+3PX75RHneWWHqdNf
dCCdPFIbntNCTkfhTAsauH4fSpzTxvJSqWvxs0NwRLVLqgInSSR7/K6IDcqxmsf9
s/9MNEqcWhuomnrWGuqQvTQEKdDK+zAExRSGC1qzI0MaFPNnMxN6r+z56Ipb6YfI
NrCGDH9XXolZcf7uByIoXgy2IkgXbNVyEtgSzwkfuu76eGJDlFc4MKuExK5plOw3
9DEWxu9/U+HAmB2TcwhShTP1U7PX6aHKHtuALpnPsTtJljtpwXQKhXBPt86zfEMX
+ebzCCpO1l8Tna/gFAXsOfIqGIfU2kpoLEiqkGKrol9AJLg+WIfPhsXzUZScWPwT
aY0j23/SFqVghVkzO9RDa93lWzS2RPWnb7AGTPre8bo5yp2ncKpANBIUOHAbhpVJ
EvTHU8qd8qeMg1Uc2Oqxj3IsmtgtvixVvV4GZM13KBXpb7TvPMoLWs6n2rlYbn/3
dSBbihW2k9vjT/HusxV3U4BIt3bh7Ob68+Z6NK3zQuo5sjMtkMK5zjcdjswAVTJp
+zJRBvmuVB2ztzK3IG1PTXYYCwcySKSTxuo9ojP5mt+8OgzxTM6s3+K+af3li3xP
V+0K/qHRkhN1RP2dyvMt+ctQnZ3SMtF4sWigp9DVT16iQ1uA47PPDZ06glRbnoXf
/ChJ99s3MMHEl2hLfwF/eF69X+LUCoernsOiNaZ2ETzCIpx+16bhJMbXR8S448K0
RPCiShqWRpK2M3ZH7g69kK4uwEk1LH0ZyRJd8rvE/SP264Jzd+zsm7HVBHIWcts5
o7XtKV6tgq2uUJnToD0HKo3qEZZJEVDz45gvnXTsj0LtP17/JMhYpk0DOysI558I
1T4bjuYqtdt/U1+8X1MBAi7/ywduvd4a0c1Oe8ISU2wgvLQLAj17SxxWj9ZcwsGS
gH/CVjwW64N2x54RNbH2Y+ijjC6TBNRl4rfuYjxyDU0uyB/kdYvLK3l49uI7Mp34
JRCLZ0OCOK23LcGIBiq2pjEt7JT1TMVKUJMttS8IH5Y6jOi8SM02z5MNsitOefb3
w4Xo51DwIp3fIZZso9YDgGT1O/32uMTy1f3Ci1cZ1Czrhqyddppth3xAAx0ERGD5
oqLyyMsyeK+1qV1Mm43EM0cu2FJM51X5gzlxg0uVjq8vTRlwGvAtfPLVm5+hpsH8
1kLk0laK4dUlm3vtoLil+8FQ4XU4ft4DtyKMcgVikHtd8KhXWuMJgodVIft6WjBx
EKS6DGR+jidbcg8IHXjuX0p8c6Ntj2C9x+zeUE13gvJu8YS6VPGfTgGBjixsAEBA
Tok2Gqn6XudZ9oWxiZtxMcY1OYxGcGm8aHgVNtCq6hEFyyXbUO3AnnBEGapdnwM2
V9s0CY1GaebRhZZxg6CDQ9WCsibqJZqlqLbD6yRCfGeCLYp8tDq8JxXCK5o2miSL
banMUyPu0jaxRL5gCsWZUcm9IkZU17Fy7LlAA7+2Ne7fxt2rEXOXRBZKmqxQS4L+
vJj8hg8w9A1I32HJ3XFq88UF87JHZzhUcb+wASTwfCR70G1U2OYknf7TWmXqeZAo
kY3qZRiHnB8aJl4amHRj8kIEySsCO4qtyzW+Q6RST5KbXRc6qvz6XUCg0kcM4QeF
f0EO7jEKbRQuGZB1+36EjBrg6jR3XoVMLcFOrB9YEwO99zQrzIlzxesm52nHsGSH
N2Rg13vNzA+zifmulAKpJNLbyfqZWsUorChkiyXVPptlW4vgNrPGQVr3Kaz8QfoK
3W4Y4PED9wwgGTmt7pJDUjR4asB880r6w3oo3Dron2bXE/2Ha8W7bgF6m9pfWIar
UzvxC4FpPv805MsFJ/+9aISHJe7x7iwrkmM6tlXQuLQ8qsBMYu2t7NR87c9sy5AV
Je1gIkVEu9JSh8qXTJF+sMLQDbeezPwzKx8BrngnYur01PPDEiBf/CPgDoBc5Buv
HvTCKoV1hphJUYO7UD1/yMuslBBCaHySRdEMbiLFaM5CLEEKhTDjNAHAsk6s3bH2
2B9a8Jk2LrCdSn9fRBB2a+7KYVk9JwmnwWIbbwdPcW2u+5cIpZTkDATOFHZxdcw1
JS6oCYiBXmhcs8Rbp3l6vhD5cX2NxLKoWJfbC6gHvb5xRE7dkfba9spzgMnCmkcD
UEgTt+r5KYEnf9i8q73Cx2az0OabRfc46TFAROyuBSDLJUXACNbnbJjJCBw2/Oit
KZo3seVEXNYk4n9Ziz2cu7PY90hI1rYoEdwEuzt5gPxzo0HoAm4VcBB0jpQkkSR8
KHr/fFIv16r3lNagBl2qPQw6LqUrNMA5Z5AaIkT/iH+0cpDc5ucGWf7o61FsPsLC
ePCRJZmwXjjzRvMC/58EsXPDERaQwPQiQw3XNDpRWf7Lc5x5bIJg37b0+AUGHaF/
1l5Ol3CdU+5uG2NOrN3K61Ib8oUZmG8F8JH2gr8hMPzpeVp+u86B8cKt0MDPQgfA
jY6xvjE0JaucYhH4Up/aCVCu1aERnmW2cCLuV8Pf3PjnngNZF7HhUxNbDgY0eO9I
A2cBEvpOOKRBXtgEDzNQEoPQAaxjuV9KDaXPduMAXggJrCyCpizFqCHEt7/D/nUD
K67dv0pdmumfCh1DGFYa0tLJ35wdTGyLDMH7VgnwAjZZYUVbbpObSLf5votxDoYj
3rp0Y7kr1PKleLcWc3V2uR67q014NBmmLv5L7jU322F+SNy4huanOVXKNBh8mr9W
rakY6QpXljxuRUpqzDCEc5LtAgo0djHQ8PdxQChHaLjm2hsFBnOQTmRTcz190XZz
YZwQY0Zg5k1+ndHEzA2qGQ2eSMRVd049zk66Zyus3d7bdALVupUKwfFP6MKP9QOQ
bIwV3SYrckSF9XL/RBQV+c0gw7Fr89jI0glQfNspWQXALKy0DXhZtcJsqScr8XIy
dlKsT532xqtW1ZxNHm98fsyFJxz7I+FS6ymBTXWmwni0+9uSqmhK2Pjb+0mgBfsN
w86wiUC39/bC18PqD6mf5tnYNJGT/eCf8dCnHq6ms1MxOEpo7yTVASEC3X6lW9T4
AgDoKBIiOVXkyin29LIj0wb9Tfm5QKyJqBsgjNkBAEF4nQvqAfZ3WbhdyH+UjuNk
SfOpZ+QsEbDySW6PiEp4VrsoBR4aYprgXfY8NCLTNPgDXs73xNZMeejnoPb7ku84
LICu9BR7coTm5AhbW3N9dJRlxEfrTu7baXo5O7dbnExZc0ttqnHTyCXn7e/VS2VY
Rl/n5mwsYF/iFNcNwcs/b5cbTAQy3/9MV3aubT+BNjcLl/PYUlOzwqDD6an8Vqdr
yWUdbhsMErkrtQwgwy8KyVSS69pfxiubnN9Y5DUn6h6P9vzLMQJ56jQF2yOBaUCu
HnOgKx6/Wxq3UqVcO/84CjDsUWbt1mFT9+hFdI3JGK7fVwlTliNv1XHxFZ4aSWvi
3R98suPVYZ841UyR/XUP94iDf88deEW56MkOSw/0NHVN1XHMOhmJ+HTr0O3jX6nP
qStj2oe3YTDO/79FsgnfP7c5nWzP7ZnJb/GqC+AoOO3pql0BARbsy7L/32/wlw5H
AOCqc60Z/ZbP4SsFGRQtfzvvuGz1QpB80V74Fzng4xsbpBbuPa/QtT8fBNtrq7x2
oIhmTFgy4Hh6wcx6rY7xCp1v8VfQ9CCAfhJ/Dd3px1qTEBHT5Qt8pJGOfYk44hEO
Lj9DmvDT4l5qRkhiryMKRnX9h7ZICBBVGmaGQoVY4WUgZIxi/k+GMRF/wStKMpfW
gnB/dBNZov2i62gpLAfET7k3ZDYNimITvaRVqGtcAkqJvWmlkbf5u4rPCpEIbOwS
A5larZgnrGQeBM+gwo/mUgzJgPfv9syJXlicxyRW9tY+Fc6231WIcyewS7d0srnd
a397r2S5Nk+8HuxKzPoj1qX0dGQ3CvxWncTyfm52mCY62fl93dZ7z09a4RFqJZ58
Yjmi9emXl7XxgAaL/IT2hZOC9QLw7swX8zJEC9NmRL6ohBPCqTsUH2IHDDzbZ2wZ
+izvkoxhYOMDVco9c42OtNcFMM2XiStfoMEazrlOS6wtXacOV9UfodmBBPI2YZH1
w73vsyj1ybeL09M+327MV6aVuy7V2BpUxHZjAj+JinQllhxbqtXXEF6enDZh2nFA
07X0K2pSOFRn48l5Df8SMc7DRvQWZWOKA0J+H1ZQTRI51375pGYbBViS0A6Cznzg
KYtnlVPGC7iozGGVJV7a2kkctfHoFu+2sn/NPVDERBPE1RkYXFcljVRZ3u0KWWpb
tsD689VqUlr7eMDs9dQb7lYb03qqqVlrQlksAfaKZLUi/t8sDIpfRXaNYrvP7SLZ
fq1+nuTwDALNWsS/e0N5U2bBZfeeu+HBs82RMr5voEz9NUIcBU23pQ50nD/OmONP
o7erE4ik9qU5U0G2vn77jGc4Klc1wngl3dAkxnsd3bvZ/xpEHA45D5usMbsOoZ10
ffjRXU5W+j4uPI3J75Z9CdiN3pbIerA3MlaVqHNvOX6NAuX7wYFPshgmuHcVwP/2
ZhFdZ0UIBK1qQAePy7LwXH26h4L8bV4B2zZSUVUyIVnsZqXT/Unh5iL9BIckL4tg
+iHZEkZjZURIJttgEPog/q8bvsqt/AOB9F/5ZJvond27xmrpLrW28/DbnKN7+FmR
e25MmuBX0ixjavJQMFHveN1nyhw33omOLyLcXxNvpAU3r1PQaDc2G1NkC2Aee7Ic
/Dxz7JzcuLEe/ZljsWpHNozs0SzVLpuyYz9OLitclC2D4RUcFr0w24KT9tYm6s65
ZuAxhbWxynAsoh8NyE+rYq6GRDYOwDNSjzoi2A9ZzigPeHKBUdn3LevitcySRou5
2Vdj+ebUTNW50xW+RyBn1p52CWsRpJg0rIVIAh3wsPWJTJf+8UePNnSpC1yrhtNl
0clUZO9Y6dQ7Y4WFURR59nkMeRzGNQRcM47adATCuxLkGVYwHLONJogRmhA7DkbO
39pbABK0vHByOk4cp8qed9n77PRPzyJtva+W2HnGGCB7UI2Np8rBJtsolkLsOzoe
OaOrHvg/Pbz7bc1a0Z03xiZzfiGTRAyy5BaODcGoN3RFzwzt0adYBzkr7tkGJJHn
pLkscq8ANqhd4MiUUQa3ztPjxYKz8+b+kqMY++2eSDefYoiheE3GvC0D7aSEpCgn
B9sW+Fh4itasPu0NcGo502Nl2+i+qFrB3tfkW798Ymkvh+KV1EjLj9CojO/CRIvV
5qc9hK7YGF8g4J1YwexNy0Ne+q0F5qxiT1JSzeapKOvNhbMWEjUC/83dQAmoXxbv
RXjAwUTsEI1IHd9+ZnOxPPNAEStTn4nEQu8EqAJReYQyrWQgQIyKEUqxNYSmMgDz
fT3L0tt8hH1lIzx4riWlzN6igBLgnq2/sALkJFJf361olCObbz3PRFhPsBeMb9FK
eQ3cLElmFwyIkwj5nz3Yxz491MnMQJRAdrjjPmu/nfnqdyzQMnbVIvK88gMiGY1I
WcnNX70fEseBQZ57kqG1flGJDWxj/jhyVE0nb96WZZ4HIMAvGHI6gfGAvbGsMs0X
UHfuOzV/jAZpCroE/UCwWuO3w4X9y8TZVkHKNaXam/K0c+tTSQ5v8Ye5SrNs3UMK
5pYkN9NhGVsCqvx9PwRR5hSEYjki1vanPVlsKp9ly1silM1XLK/B4HD7Lgz+5lIY
STd8X9T8GtVN08SHMDa6GBxvHM7T1vNgyT953kEX9+lLLbQnQvbJKbglCyu367kv
cOjlFV21pS28ZOb72xM3Ege4e8CfwhtZL6kRXS3Ffgy66wK64MMM7mrvNwhDKamu
p29gUpoFzECrYr7xP/HkDt8NqCfU93tGa2f3kRJLXVw+A2J5Nd5riJ2kl9aA8+s3
gLoLXjEjcMpwiAbNaSr0XeSF+yHTKFGy8xtPE8rNOpEH5GZiz5nJxbWIdF+DijRE
OciSFlwlCU6KG2uUrIAVjRd0xCCeZl08p3to9cLJ4m3uUAk2WKdR858gdzUO9SWR
oT09K9E4FdLb1DQLsHQ/N3/t24VMvz7lnUT0Yyz/K5zfs5/QJ+6OXDGJbjtyf0x4
bcZjgVwZz2J2SsStWScgYh/Q067jU87E2ISy4LISSznObWPPfa/W9o6OPm9P1t04
AWRhYXVV/p5Do2W1IZ52CD4kvWLDLx03GdlJSTbEHnhGqewyODBGZehnpbtb+IO9
ek2Cupg5nwdDwxU/2q3CtxFwCqqTI9T1oIDwKA5IjVLzTccYSaXBoklPcMSiIP62
hYFLRF7gyfbo/t+ytSAfmil1sZUsgPxvy3cJFz3pMgq/X/I3YYt3ndV6p3hVtOZN
kDaZPplmWfXMUwfAx/oOXWAeUZQHrpfj2T2BhxQOFpAfozP5RR7OeFfO9v5HTbVV
uZc9Qpc9tR4HaXzrQBCU8iDnkKzb9wC4nK9kMnVaDNio3yobMH41FfRd6ggW79fX
M/tx8X7HguX8awswxx310F8secaf2cw6OKFlIOAJ1ebo7DB1bXcVh+jdh6iFzAbQ
e2+x7sIDxlEvdzKM5Tn+Z3IxkH3oSMRFHqaf3mSJUItFcLCNTsbqLRqOfz2Js6V+
HzZtIx2GtYhBCoGjpE3+ANfub7ID5SAGi//bv/Gn+kZ4xmeCYEOWRSOBIpoL5qQu
r6bF/6pGI889c/2+mQwBgaU1CAR85u0ICwASm8slmJcwziLc1FkbBnT3Rfvo424n
mKL8NCJNCrIbuldb/2uGr4A4RBssautiWZkRm5CgUIBn1zcS5bkxcfRfo5i6siuj
GGGjb0xAKAnEwH46LB5y1/L/EnOaS+XLu/2MTy67Asa9NO2hMNkf/h1L2Z6IheQJ
6ZnkWRG+IgAr0K03hEjmRxw14XSPVdNkXV2yiJNTQDo6MWLIGflsLJnutVVAfXbw
hA5/f6+Ba4utQD1LFJIy+OZoZKTd9shQ2rn7PblkQ1WU8dvWEpnTuLMj2r2sYJCm
cSRlThXmkwXsuRGgp7UrpDGoZEMy3Is4jP6v/KHdhGJyhzgxrXTp6uVJOEcj9T5J
qgsgtVYkIxQjlLfqBGI1FF2U1wAKxZJsAzKdIFr5eFlfNS09qnQQml+V0A3YbKGO
D+x2o5IVXez3VWUnn7cgOkB564VIh2sejnYOpHIibScw7henAPyEXmQYS/+HCFJL
PvZ9PAj7hjlpsGFZgjOni9RQNYKpMZ56ChqWUNIsR46rV/+QbXzJxtsDb6hO5xJt
VM1SGpzQ98TVHX5sHbI/wTK3DQeaJGjGFc3ax1YXLSmkhVEprSODH0iUqldPx/t3
E6Ei3NCEY4vI1MybYwDtQbQtyu/oKBMyu67tbq1PSpZ0nKFujM0hfzw2bmIfEuSF
78BvrmSJ210erMJF5hePQOpODnAU+uGaetu6IvVjJn1elM2TD5VYZXBlyUHu5ECg
B82p7BDhb8KcO/EHRkNBssq6H19XsIUfJDVvMBZSyHUFDfxoTHViGt1rOniMjvcH
pi7VG7H/VYiH2P6LmAI5fHrcpstPoJ2pwIuZIvu642nczs7trBDjUbSzuncPcq/M
uib8iPfCbDJGUc+MnUAuDevfHqS3nlUQkqj1WRlRb9+ZwnSfnPmdBYfFdiQbi10t
i9jojzSG0aqDScp2GRgdV0zGy/6xZPIndSM+s+XTnGVu4TLh4n4BLTEDNQ0QG/Tb
qk/HKRxayPzzhpAy4W6MCjk7ZLXuDyxKPIy1wtTyFodNe7sweA1VCC7mzixm9E1+
g/OpGgFUbEEowUpJWLeQ+8nQrNlsniaq1vvifH6qRQdJ0I+sL+aFixX7y3WC5/Be
AXBtMuFVwTNVEG/I/bC3efPhBDqCVoKBPTC+3Lx1A978ga/knlnAGWGRCNTdDq1a
beBaw8N06uA8UWgVKyVbCBoyozdtzz26Sud8PcIC/b6lAuFqw9wn4uHuAN9MW4MP
t8ZbJtbOWe53rRQY3XWdzKZKvpjBNLgsSV3qlX1pbUQ9eSIZq0TB/BHEsCbo0o5K
BAPHsWuPpkQAGsfNEV33FtZUABRyOpi0vNi+q9QZTz8Yjd8b0P4OKEWop9TKVcZb
HHePSaK0mSqyrwwDhMwope7/hH+jSUIo84MQ6EUwGMpPMNugLXhUI64H0LpGQ1fO
fn9jiRNlX4FZq/UcIO/0/sQ6jaC8uV0nUj16fZZ4JUvafSj/RDB7CGgsKLvGKyTW
ERVA7TkOXMqhDR7vcR5qhsVGtK+t6Rfa95MTaCj1lmcDRcit7165QjhmVSKGz5YN
IevWTD/93rJLi0MGvGgy8kPEqc1Pi2FufeTiYcG9aadAN4gp6t3btgn8qULA9gqw
gEOZslzJcEowTKHO0BWtfLreChyywWHU8Xt6B1GfIJl9Ay9FbxtlJn0KJHCz+WUF
aFxLlWEJ+66ZZ0sV61/MqW5vs71oWivge1hA7OBLA0YGFOuUh3c19Y0TmYXuEBSF
JDCxLaSq2reOKgPOe0X4NyfPkJpij5DD0UMG6JDVGuAYgh+g8uZwFSXj3DKofQr0
ou6EVE12M/DXEZe1Pd33conr3iH2hZDj76YAmsyIhBQQmB1QJyJ0IBIpL23YHxVe
BCFVz1xk2IfUa41aOnuWz3pRR3XOxbnMQMgSkrIG55IG0ESeQSqlHJwVTfC0rHt1
RjM2uBWDKOQHRDW/yGMMAiNcAoKxbyitkq64xUK1gBolYS7MZ2r8P3b/H/vnYAg5
Lx4IKYpeyH9gthY7vYjZPeTBwE51FMtYgXyCFhAj3thk4g1/6YEGz4rDTU1Oy426
MZ++1PKqw03Sles+M2soDemrnkuL1UM8VEvKspyrDbkO9DoPcQlB8qinGFZt7VFK
acxMIw2YMMw9twQisqnlQPwuLmz6Uj3KZpnHme9Jiz0uUanqVEbB40MsknMJJVQ1
pZqHAly0YTnhOyG8OPU2MUj1LkVlFhDQZAScLSo/blNDxxh8yBNCIJlxcM0TlLXw
Sejc3INJQMsbnH3QNxrNJad7NPoBM5GMyUgzHdzXJuVNVRGwfwocafTjSgFUmdSc
ISEZ8eP4xWaSGHtesm13zvuYK3968OcVqMdJCK7u9jW1UPDpVcIReyeoXgvUtam3
dnn5WFkns5jOmiuNcAbkl5h0n6Eoz8v5wRb/5+Aem1UCqHK17Dh6+E5Mrx7GPjMR
9mrtH3oGaRc0HxAI0+RLXiaxqYDm2AY0rrCWaN+MIq0SxhqWfH6WOln7CMyu6mUi
666ocJv9YR32Wv/bHdBkXkvZV4CDVr1tXXZP/l7tSINu3kV7VTj1DOqaXB/KVNSK
hUjse/lUXrUCIWf6pQvDLopXwp7dvlJcRfa+g4qXbdGvpnGuEufVaNbkCsggRcAr
Bq4KtJ6s3JeJJr0mqD3rG7fdIm0yhZPP/rAlY9e9mVFIEkqZ4E4dabxyRh4+Pco/
7jsydaxlC48Ek8Q4rMSMkMpwLF5pIBuSNBo8R0thEM4/2dcfHJvYZOG/uBYXHqXR
qvXQ4n7RppPVY1TA1CtaNdAgasskmEMmNJ7faQwTJyAtOegJuGQqwbASS2D4q8xU
ISmMnrfWibyvldwA5E1Po541utDQHLeNiATOcHYl1+b1NRLydk7GDR4hFChZsHhG
IyfkKko3o4X8pmkVs8k2tUoWsHlBW2JT1F6XLMND/MP1SGA5R5/MDlT16jTliJhX
QKzxSl1GxEYYyjsPpmAdhvrzTMT6nysx1jdXfH6GlGhuO/FUYoQjmUM6LrydqJeN
thtBnGpvMfKsI+YhG9nmZFZBauMeziZMFG1bHRSLNX7ndmR1o81v272+cdvCDEsw
NFz9ZWWtQRd0tPloOe7/IuKI8Q7FrVcAIF2K8gZFzYMbP4at5aMK53kM+3b0L1h5
XVfBNXUfLjKIFTyrhA27RxovssO7D0gFTPLG3XYotOu86Ncvvrk/br+1UL0Sx9wH
ZflWs4K4NTZ/d/3mez8s6DBumrMbt+eMOvE1I4lXtNQrlPsKRqVbGctohyp4/dqP
HfLk2A7p8D4FyxY6DeCF2WVchQCpHMAWLKfdQMfmFcYIZr9x2r94M0UUy+F1+1KQ
xuK6b+S5u2hkNkpJY7b8kP+ZdBlGzRo7tcQ+cYITGxP3BW0R3eH+9gx4ReYYWUDP
22hqUDCwLa6zm6EVYrUaE00VZW9AARmXtVYrAITGPRdYgmjVguCcqCprOUbp96xk
d3ugnzaX6idw+FORd3HH8H5Ta+ZfIOIFh/c8kQPwF/uhHTmkWdrljOeFgo86xF5R
JMGGLQKZent5E2YkwtJeLkGsNNT912rNMJ9zuY26LahURRXV0c+GE0J4ojp2LtXf
i70rfJGK48HbtCM2u+JlyNbx+wD0YlGzwRedj+mc4GVYnwguH8JxaPQESNyOZW83
dW0AZtvyXtowMXQkJA299/kG7ELszWraoMW+qqGJ+abEHiEvj2jkhZZYqCWRrSYF
F6pMYZKV3nibn7T+m9PYRr5cvERvkCQFM+0q5upsdJERyYXNbtroESI5plTT99Oe
XI2uk1ZAG+FE+p32UoElZ7o0XQ5Om14WuFwkamwSUpALTOLoJ4xKPEE+EOiBvi1r
nu+Hp3CAbTnAr3WmmSd1djSynK015cvLWkUkAfdzrWhAh86UN1BUk0i4GNhTVIxz
HImuAGeW9IwB+QjrDEOGrkAXGpsHsldu43L1k07ms7+1bmjHoTVgdpaJJ5hUr/54
ESHdDhA9AZMOuWYLVVuY1y/kYiRp8k0aM/o8YtSXVFzGdsXElK2czHHn9Mbvw9a5
tRxvETMsylvlRexNNrIWpdSfXK7eF9SH6bvNodPcBWJ+14dCFcF+5k9kDSJYRA6O
2DHExUeKG8esRrgkL4u/eRCurQcYjH9d9gq3NX/u6RkCZoHFU3HCZSNiZ4RD1+9s
Hv8oPJ9ok9Tc1BPJF4p03yP2wFhonEEvc3wmj+htRGqT1XlL7fsV2pRdyfJvAG58
PxK1bvowbA3skdft2XKcGv20bZ/gRcVPxvmrlsSHI2PNsiA0g/X7H79FXaumVtOp
BATyqDpTSjr7qYP1ehvue3+0Xq3a9rJ8OJKfSFoiEAexoxdJ9cfP++pJJ08ShAQc
5Bt/6Zfa3vCvsjDLyD5BwWeqU/9PjtgdDP5YDlnpUeMyoMjkBlEEZStsJ2cgfQ0V
gTsq8UY8VMXZrfKG4quaChTQxsZzUswK6Cnk3dMOog5UugE0OvLx0NWtJcZWcXy7
KYbpb0uemmHRJrfuvmQ5PEk4agqfd91ornLaacny93EoFqB9+EHs6PUpxqQ/tesD
h1YoJAu5lKZ2q3Py7KymyECCkqlI/eD+DZvnXTzeP7qDeBKmLeavnbPy2ViRU+NP
/BjN6lQXuna0rZP1REYJdeP0m5W88wxSe3cNllik0U6QHmQsvMU7PTLtzzjc2TmY
89j04TihFnQ4MhwAhum8FAXUgrleJHgQEFadKEczVe0PC+eJefAbxDDImn6Hj3CV
EVSqt25E0k/qEoMhsxLLQPl+j/V+ic7R48hZBYEMN216usCwMd8RfGIR1QNe9AYi
8pM4g472ynsmE8aTI37h92XeQJMjHTB7muW5UqlIJeRl0kFNqgfA7UW9J+b/w+P3
WXoVpMQ/Ufsnr47gnW4Ubr4YF19oJUOuKxFWe7SBjdW5It52mRZDGI7Z77EvD6Gu
uWn1uRsFIJ9XQ5uyfRWeQVY5cvQXaB1Q13cZhTAr3HzvEsvXZLfc2tBj9vCJ59AF
utDQsMKw7JDCYC6FIPi71HgcI/GwxN2F46VTlsV/tb6nvfBqdw/lBHv9o5W6mnEU
fONFy6B5YB8/DXyqaR9+i/We/Um7hyO3K+fkJ53HC14I3l+V+2oEBospkkGTLltI
W7njQI9hpmInMjjKSfZBS8I6/NA/Qufh4BqNwLY90SL9A2og3jLAIRZwblWq9wIB
JWSuUfs1fsNjepO7UnD0O1a3QgP0SpIiolrdHdQt11DH2DI+BFTiXn/29+pnd6M+
6U+wKfpD0zBPtBGj/ggLTsXF4AVrvOG4A7/dsdAsE981aJXfO6WEqUXmkb6DnzAU
/ffr4A5HKX+7JY83Axog3PUxrzu3gu5Xs3BlU9T/h3kVSkmz4L399OB3QfS3TWJF
/9ODyefzXHGw5sMXHNJEGpMVcXz6DDjNXxLKnF3m9Q1CENqMVoeALmgIHXOT89wb
lYyabB2V8ztEo7gq+S0M5tpmcdNstupod7CTBliluMIlf1Nk45slw+w59dT1AOan
CWQJvw7dROrQu4MkIhrGMypzvu7tsjFuOmWL7dMuuSG8CzVZW+EL+RsunsmInpo8
N52rh4jhWWrzAiaJ9Xbs+RJNBfjicRc2uuUfsEQ/I/ZOGLxgr21AWTOj6zqfDTvj
2iG6ATs13aM8sSxbfrFYpjd3DxSQvdb6cZ9GTsbLx7xhw5sGM/X7JDqT/ecxgvhC
M6dUuti+ikOa3YddLCMsn/snJj5/ehgvTwPcrcntGw7l4r0bUz+FccYF156F/1YQ
rmFrHSVRwsS6t21IPoEIRql1NAWzgm8xSwNe1PmAjyoyYZzV3QhEkQG5HnB8W8P+
SZp+HAcIW50kZacT44OW40puM+kVwdzpkddUpbzhCSILoVEsMnzHGTv7KRdGVIsR
rROSZ5Giz/CR0acuxQeQzc74DVz6iFSj8RBBx28Blk9RRFbyGTDXytjuHcGF5DDG
/Rit6+nCWVboc4sWe+zzYgR1KlwMuMN5mTd8bKMI/+Bnk7yFpFYt74NityqUvu6g
8vpxwsrkixz3/LvblFL3QW5bsGpy9niyeTMjRimBSc1scsUXP0Npzgngpawfsqz/
`pragma protect end_protected
