// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SfCsW0ZMw/ok/6bcuktFLn+jrjA7MRbPtVlWem6OlStztyfYPWtotcLw76yTUuNG
S2WFdM5PmSK9BbWMJQ7PhogZiZYAcrt+2zQJbTliPsh9rBjnN0ixi0RjzECzPhJw
4cAGAlVUIS8POtkroTREeaNICiLeBl2DQI3U6JoP+p4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
j/BFO3mvXaMnaZ4BhuhmPUOBfDMoUVj5vqENWQiiHXnot5xVR5rp91ujY66OUcDb
7dIGPccxhKz2yE8rLKDg5HXgxU6mIKDVRyEQTjYJpIBttMpfXqVuvsy5ZQox/In9
072GR9vwBUYIP7Tz4905ZrKrvZT8GgCeZ7Vq0/wU2ZPzusKJK6uP1wlr3DVIz8C1
2MdmO6q3iNczSO7oN/dXBJrTKy1xpuqornHrAoEgQvmW69LpYfUFbQf+XL2rxIs3
im7yA5BeD+VevMTpAZDFIBQ9ZznGgYJ88AqXmAE2IDr1D/HCeu33/IMYpNFpnMbD
HSO627DUUJiFz5no7XHlDxyxTFcxwrSZg6j2tFvI9aplYQN7lkp9j8aDYmjigZk2
yOs00KdVSEu0dDZ0tpSRzgWRSbX3fGkMm7X+SqRCEffI3OfNEEzNdtWqQ+XC7Meo
Fkxvjfhga1Hv4U+CVXrGZpHS5EA8G7aJwsINTA9OXeRwuNx1cbNUBRKKhm1g9M1U
KDkmqn/eyrDDW9QX/sUq38kDaxV+9tbaH7G3YF3zYfbzfH0maXkAa9rTR7r+95HL
wLGb814jXFdkKN7sPzY15rlxlNSKMFRz9KpjcCYRz2F/9Cl+YUmetgz8Y8TxaF2i
TM89Q/7z7M0d84203+vAVtocgrJAJPHqBsfHFR7jKiFo1gUKIPOpY7VVDQtXCh3z
apWwsYp4LG2nS6nn8xbL7yscffUcuFqJXUqujwSsJaVf+dWRHRcNT1HkuGxlB2p6
5X54fFcU8aP0QzlNc8YvTjRJlDSigPuwA5BF3gMpSvjVWWojIT8OrOirkU4S7NRq
eMBFlXf86cAvTsFebm1tKucu0KkRoFIhES8FOvyHen1fDFdJB8pl7thvEbvcg7Od
EhbZB/xlrc2mRRigySPWok4afnPBELAreZ4gp6KCs1OE9jJFNDdc3wZXC/Nsh1k0
BXkf4QqFcuQY/ax2ig525JAL5UXt3FXM+B23M9su94FrstEVmtzS9XOH37PYE2mK
ANK/ocqAngq9lB/XobFAgkABnswnuMjHAeGDFURLQXxPcxkz5T3T2/22A4/TCP6O
+wpbGAdgvdE0MFm+ySzUZ+++nIXFiHnQT5jB47MrK190lCfHFbZmKjlS8e0O7Ptl
d83QmMVUoniaUEbR/74nBOfl3R7MtOU4YjUBmzVnUqXQgvhzmQU/bj93Nal/e3yA
SpSKqxwcbqcnQ0HkVeX9l+fjbCvgW/IICz5kOcoLjfo2iJ7dNte72d/SLsQUq7RQ
RHTU5r9kpm5l1rGjhiK3NVJ338qQgJJ0CaYHh64VqfrilGuuzy6lKA8W76cckLju
seGZdtG5E4A0rynyB30nGUab/E4US6tee3HbqLkB0YVhTlE+jJ/MV/MurEtdPq52
wBoWqWRuMUqMzPA1vs1a5mHMGGHnSdryKHbCMyu0ygmPx3p/iqoI1sAMzFryBkf1
25umWNyltatAA3zE1T+hvKgHo5mNe9XlSQjS8hZplljLyf9P3ySDYv+2covRzj8a
4Gn96ZMmL7yxOY7e30b0dJdSl2fyN49Y6+yB5778HFPhPICMboABg+XmpxKA+NHX
V798hko+TI1fzWQydhi2NDLQmF8Asjzu/et5h2HxXFt6j9s0Mu7VIxJR8Ld7M57Q
DjEXeAiSd9c8ZkkZ3lXvlDBpvaDZinoyFKhMcAhYsauuIw1If+3d4wkPChQcQDxj
gr+tcSHh/HSeoD9luZt16zvBIoy8wD5Ezm0o3r1xYTfTIlWt9xlFq8CY4Dzj1YH8
XEVCcWh3+TBRKvFjP6zop/+ienqhgzpdvuebaVwwz8Vb92xGF1ebx8SjzCW3Lz3B
JTQIEW78ysPpNr1/DFGoBGUKzMQ3nUGaxFq9HzF1H2KJF3tN2t9jHbvT0YSjPRy0
N+yvd6D3ckJO1x2m5KnaMuAUi+XaS6/p+pEfejeliWhPI2QPpjKSIQ5xI6mjsAhV
M+wWsQcfFIOxohLYTVsEiBZQm26i2PtDcSq9RePRqI4+TLs4J5enjqSfqSa+KIUF
MZGHzK6q2Oqc/IHLGuyfcoBSKE3mFJ7qncSjbmdNWxZI7iInEzptsCFi959tec8T
B+xAanZnfTdPcolOLnPYIqI3/uyGc3oZeCacDTzfRn94MqE58tU7fl5uvfhuNECF
3D5sZWwTdrKEQ/eLsHGu56QAI9FSZkWtLH8V6C3LtoJEwDodu/ZwzBLNJi4s7Gkf
dlYYoYnaVGbBEGiw4UEG3zkL4N86kvf7LLUjGYhTowRmHkef6QqYsSD5tuyz40C1
hmi8mtiNaFukrrnnDFIQCQ/rxhRxNofBwzK3UK++sbKzAZhYfAx2EuR32jECnPzX
lFZiKe/CLOdRbQnYLvwcB4VSv329Qlx1e1rponHWc8CNCDZKJ+Jbx/DHeVSSwsV0
/aWXccFtK+YzmhK4uQdDNT0idXy7+q01QvxCiRQVw/ldIa09LXgekbEWuhCL80DH
ig8kfA4MYwqKXrauyDlk17JOPsR2BSZuzPl+MuVJ1Fw9CgvBJYZLZrYG6o75NVnj
zI7UuVEOlAgELmQUXCRYq+w+W6Kxyfr1u7Pby1YYRkzncMCLkZ3XFy0fLs/orNwK
d/6msc1MX3ZNm2WJqzDvmTZAs/P4mdWkgfJsLkxpdjuoJgzwkjkFnEyOYuEpmIZ7
5l20/aljCIz1LyMfVF9tmh5I/5Ciia0kMVwvYVAj3nm2oYV5dF46f61T6hWMtCpT
9yC5WkigVXRZ7exRP3IW/d05lbEhPqee5dlAlAgHEVZVOZC916PoRbdvcr8FlFuv
BcZVKPHsLVsXSpwGhTwaISxD658dre2PPGj8tJhss3wFV9CUTmvHld/+ULcoXJUR
pQzVHrb+UcG9RJ7fw8lj1GO9tFHkvkbyjhQwUhSSDIN5tvLOV3lXCFyEVbwEBoJv
qID8VNPsETwL5as2DBt5Ow==
`pragma protect end_protected
