// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
R3T/yq8Rhq+3QsmK0tN9d30BTunsEYxpiHKYOey46KmSoXoThQPNqfpI1aaz13tlKvI4WLlK1Zv6
76MCOy9bnX80/ya5QHiewN4A6iiLaYZwdV2NdJrex+DykiT4Zb2VwCYFULeONMpRxauR5Y8DoB7J
zcoZvJvYo63vthndfQo4vMvJr9+zGxGnMjsUmElhDayFPl9JKXzuIzWYaXSLrzUXPDRYWeLGHqGS
v0JqXhzvshmytohzWu/ZvlVWxpNMXE4Fm+jFK5BmhghPi/oESJvJIA+EcwKbdl8qmAC93ovVXVm4
IJObI2UUPCF3TEj15YYxLon+2IYzqNhW6IPYKA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
jMQQoCLNgiqFBKcnOxDI7EPyQjWWjAcjtAohMQL6F1ACFPX4CfNj5oQTcR3n2/J0UpkwK5t4fUWE
55j6kAeME4d4w5UC2RF5HtmQFY8lOwkNrwcbVDS+1k9ujHV7GD7DOKi9g/ptRE1u8VPcRudZMqtE
Gfu7rcMKnHrurBSaH2uvvR0mZQwJsggf1lNF7bkocGhkAAUFbsi+YxeCqsm7e1rSH9TM1afZe7Z7
xYKAY0Kh+8/5ykVl/lilJyTrSyjmVs+RxeAKf/8sfn0soKgaRK3C6kP8ZbH7yGUsGEdJy6MtN0BM
bUVvV+HUVEJy2o0th8N80TUwpGLP9rV/5KcnWDVOK7pqzwRAKDtNNd9q51KTQkobX8n2fpzo7HVt
aweZzSaSzYAfpVZmOPADWTaLc/VbyjRSD7L1skblxsrgwSVmxmAvUtTg4KALhztlBNqQkEKtB/dX
pDyeP/yxE/kY8a1C4AUcaG0XPFq0kS3SmAYw/E6qQp772pLwPFrc7tLwskNdy/6zSDneq93oWriR
rZIs3forkTyAYmACglO58jS830shkMzZeIehJr2Iz0FVRCuFpAI+Iz6QcKHHUshaOlY3VuiQobHs
155yd4lp/QEQvFxq4zuQG6B7EkYxYH3ADz4oyDpWq9CbWlZB1JEhnykUUwjmiSqN2Kqp0OeFCePI
9hxcRRMDcKmOlotEi6o6SzhY3UgvW1kHchjljo/uW1fzjFQIl1XbYkEEgSLeE2Jt8beez933WiI6
tWGi8vQ5rSXw2G+J0gt7RrXXTYpAjY3oQ8J1oHIpWmUJzFMpAoeZA27qEQLbOTUQDhhWKK/65shS
YyIsbdmbJZUikZyKcpueJMlrGyCmc5x3XtTk3DQqnQkSN0DcjP7C9BKVDUXjuibVcRrJHbIjTn4f
gSBa4oHtEc01iVkOj9hy/KrORfCww/UDb3gVw8Z01Zzoa/5Yv1gwBX5wQmogMJabCNvMz/iLq0o5
LD/p1Ejl8K5cfQEPl9twuK0fXBM5d9W63BZC/d6IWL3LpSzYvL0CS2DYSBDYkOJWas55rM+HoBtI
UdHU26DlhVf5D+zsK/wh8zimz39M8d62VjfKfLKcwIZXL+LqY7+uoDOpMI0fJPE4L7ex+vXHryue
b+UUhAM4l72TdbnM3UKNhsfOxQrfrBnCXaij1r296d+B5xvfx1yurs0a6hP+D/8VZ74QDMdtGiyE
rFZ20XyK9fzz27HoDXiJ+g19HJHnfRR2+uRj4C8KWPmVIQt9SmCk8d3IFX2ELMSJserTVaCuF5nF
DyhUkz9s5r+e192g1b/EF8IHTpryXWadVvLkb9oJq7X3Z2ZBWAWfdQRDczXyhA75tOhWpajofzs8
JmkbUxcZO7OLxsUDCFbJc3heQWiSSNtpbziyFSPkw90UWLU1lrq/9Bf7sKHGa9q16/8v5I01FA3p
GJluPlEQoVkC1xA5q9d2wF3XP5IlxEjgn4iSCxiM8lmakTLpPGkKIZneQnRjkBUlXJ3uHfEY48Yr
j5pmVQnxpFcvkhwoGAIhqsQHpa01hZuAD+p3bel+mUL+UndyW2m9wENMlmCqfWNz1zD4v1ETe3jl
NOnDCd82vWMpRgnEaxFlRBl2iATeYvlgbrMrXC692db+ib6t025uoNooLP/fkPPCvS3qoUYJE8Kq
aZsC0UqCq39+Lq2EC+sY5AEbZojPzyckSYFpxRqJrALHlPlFQXXmPjIP4T0KEUVeRHFuusmEPLa3
oHnQBRoNEqw3F1VKIdeEcUOV4r5WutAccysZ6r/kw9ew6U9SOmD7yG6wmg151EMzA704LPGMrIpf
Irdjb8ooTEQfmNlUKbPkkYyWHcAW+ZU2/baNOdFIN+2To0pnZTCA7Yp352xWev8KChgSGfx4T10h
J6YQ/YIHDzgs+jAXTWfIeT2WKOGVYB2ml9sqP+q9plzUMumXkMT+pBEwuVBbmKzsXfSNsgibHuCb
PEu4qMB8YGk3+gMWXEXlVDBoSARWZEDYXtaUbL4cIsjAe0Lo3lIHmB0METgC+qePyxNt7N35XqpO
6t6S8HuCd4ueZt48bq97dhRPvHDUS9zH0Fpp8fLKGvq/moP8vKfgCZd9Ue5f42wNTkSzwoVhNYQy
t7stItKdOjX/ZNrud6A+DUlPU42TKK9NylBl0JDlL+NXFzVIj/20fq8F3ldPvLYN6ZqudbENhHPK
qaGUgoCmawo+zKuuNTivul53B6VOS/heJ05ZLgCBtEt6tDhY6JjWT5OOssqusfQXAdYIEWagq/sX
xgzsp47I0weEFzlaNPpIld0UiZHk+7dlvG9f5cGFA7DJfhabN3ztB6E6Izo4dMF3jobomhJTPOcB
95e85817G3BeiVcfC0oq5bkEC50sVLcFzeKDVmP3C7gPLWgWVuohX2jEyvgre1SLZHTI769PJ/Qh
WcVJIzmRS3Di0uS4o2m7jYnwz1YAvO0wOkYiuxmNBZy56XX7+Tee/3z2yOfAgQvIb1ixId/irAtR
3rweVNthYLs3gew1YwzybTANoPxPY7O8OGrL+nYYEZ9Ev1movk+cxDjHkmEV0mEb3g1fF1qZ3uZK
GDwfD1SdlUIHSsezRI5NsFizCLOx5tHXaa6MoIBMecf7RDGSmx6MN7zmYAtVgfclhHp9jpC2cYLL
/7Md7m1pfQ303CWpfEv5fCvuSTw3Tl6cIeCoGMU05omFpuT+WBZxjSv3wSMdttWqISfTXUa3lGCW
CHuOD6bzQK3OLJ+w5bRoGOFnMEldiyZS2jtedrSm6ugD9mCgSEKJYRP8d4mPV2lvNzgN6tImP6Km
uOdT7XFLK/gwoLQl7RhiaE55RAKlOZTWVI8jnQMhdNgRPbsUu3RdLloREte1Bwl+EIQ1MAasHUBs
A5cbTXqQ73A7GLIWCKmQNdah43df+MFNzAeqEjEiG43j9bV87kuFn8Vv4+SGmC0O4NsQkT74WfPg
W/jEe5DBDjqhP11N40XPGAnbc2kwGggXrW/InMINTaq0ppMWn+p7PSUWtB3ofBLtz3mQR6Q1NXLe
/bRrryDy3fpWwKWuiCYMLksDjhCSjgXXlHZr0h/rdEqN29miSA504BIwc8uIrG5XjOjexPtCrL8x
d20CwI9zvI2aDyl3dS++4V4EinMMwY4JDBp2JH63tKx0LfwGCxcVNzHuH0r0f8yQ+M6Xq/mmngid
/OSTpjKogGbkBUDRgmIQtu4Ortpppbl46k9nFvd8i+VoUrPDLJkNNel2cg/dySX6dA1gIY74N8QK
6iXHNpvX2dRK29Bs13h9BiCMpr/XWeHocZdejnHP439mTov0f4ehQ/B95H3Cx+CMHPu0t9+2lu6/
e+d6QhHfSYOGN4TAYxl5fS24980lulJ9wpYryH/jpZs1Uim/eSduyjrAaJ4gdjtK++BfOZzsk4RL
OecAkzURySLIvoOR5alq8C4eIyciKnRVkrhiAnS4vlXqRHRg+E/N0+VJ7o/WFjUzMzHkWvKlJhv4
7gxwdww0cBtZVc7ais9E++XGkrEoAGfMVHYn8f2OF1/Uu41R3DGhgaz6FKAjKaiQmYFNiJi82kyQ
oZi2sSQagJz0uLQFF+Cw2bka3ZlseDTZCsiyR6Ldx4WfJ5wMrMpBGsPg+we3Cifpa7RN4MFm/QmB
0BeNzAXpYW/H3UsJf4EsUhJhP1R5UXvDdGp1iqW35zdYfajlrpkCE95tqb78RJVhhvIndDZHurHs
GiMxPzOOZib/4sC5TGOLe3CFTi4ZbPdSR10dNhxflKpb0ELjI8Uj19np8y2R/L6qX7lChgIjt3HU
T0P11NycVtTvUprTaBHkYIkdcI/mugo8osQns9LQrJAYcwAKrfZnWKzm90gQEeQZJ2Enhrfw5It4
dUGLWLPF0h1dyPHcfTW/TI3amdHxihKQa+O9VMlHzYV2MWUe0sAwB15ORWdPqi3U0XqknPDevM8f
71D+h0PcIpNj1pN9Pv6ACSurz3Ze0gTpdOzCWWgg87HQwlrd5uU5TzgX//LlPMKTRAFyu1a4s52k
cMTwl9jG6e0D35cYboaLY+btYSzVfeG/T3X3lO+B8TAWRwQ/YKshUhMQRpNvOuGWW2MVp5toOzbB
pA3DAwwJmf9gKevcgDygqZ7WZZl1+1H9jE9OhlqcPpVXxUIywT6yb/2ahMuIui+p+RpVID0gLGSb
EAQFQt4cAxLNktSN8IpoSL4ZDc8VsYlLdXzP0/YcVk3a8yyt81bAgKZJU08Oo6Rx0+gHqFrzaPTV
fQoE8q6sbHMXKs5Cyah8VasqiCqsVSbHDDxyTnLGg1IwDax3PqY5CgSOg6rhoDCiMfFOspXtHJOx
YQJol2h9gSrnC12/ujWBOadktUrWvxtbLYXC0rzYxgaxyI2pCoJzFuFk1xhERwhupN6C1ITQsrUb
65Xu0/n3GIMuzgiJq61kuIyoiGPkf4d0vwrDvbZhTXKOCccwoyqrDthWwA/bmuye3X5bYfIUOp0+
DumICkssAk8e7j2vuLmweKl3zliCIidyPjC6BC2W2LBVBOP2rdNPPEN+cTF4gXf9/jpv05HtAjU7
WTiANc745XTIWOy3JIaJJqC33Mpq26UySyJEoaKl03YZda3fqfLjKxPy6yv8fQwOIF8jd2FL94Vg
0P3MmqfiCBIGj8vKXrM636OyKtHR+QzKzQIlAse5yWmrj5im5Q0QaE1BBERzGqnr6w61L8T4tttq
ytB/X+LkaadKeuXhh6muXAd3p3ti3PjTedIjTHLToM6yWUfHJMNExq9dP5chjS6YOKgscC9FcjbF
5Jyc/F83pUKtNAlF7I3g0faTD6OZt1HRAgHZ1+qfU/xvkC2Hl8oiz0uidgX8Vvp3noMKb1oQfqdT
v8QFDTqUktz0QAlwvUYDzaJBXE32RzI7pneZbRATqJ0SPh6m9nDcZMC/1eRCtj9J4bAtM0w2RBwF
3cRXqpmTLbepXN1jpcO/ZUaYUW/RmzvrrJ7JLz5e+mTnYIvLS9rMfJRylSV77EC9QFi5zJ1QsVo2
VYwZKIoL6/gTxXbycKTBtzE2MzAsdEPQtQmQt7cl9xT2Jk1MAcNzYkzO311CknX478ejA6/NaNAk
BWhrxT8lntR9VHS99mLtJphPKd1lTTiaLVkdATGiXgF+dTXKcNH9LeKRnjuC39P3iHsYveeyWga/
98YrrM/wUMpOdekyD+qz6xn4vVTWacRGS4bKW+gBWujn+XO4mcdmQHanRMhP91JZK90C007qiKDf
AL7zsObwYt8VvUTcvXh2VHSka/xT6pKpnFgpt0JS6LRjvswNEPO7xLU/mquNt1HA7PhifjomjXKl
V1D2bkROdoWyjnU4nQqaa2kGb2oU4Hn6qK8iePDyeaWuq0LQKvWTxogk3DBCjxkjfg8p0Y9do3JZ
R/crHpPvqlUY2V8rZVM5ZRqiGExgoH6IROtfR7zMpIc2kNvzlCXBnYQtkoc038ugMUX/7vcrTHUr
fDEF65MddP1ghmfeGCwOxNWeBBL/f0IrUDK6Kq7CQuxOuRu6KSqTALyV8MPZG+u+MQStKiiXVwAZ
id6OsylWfkHY+MZ9zUh/pYc8sQgFog8rB+/4QDE6WhrEE+fI2bdZlDvzBlu+qga3f4kMzyyVoQ3l
Vs9zPJdQJoaBEwud+l7s6YdnAqvq27SPSTPPk3QLcBwJq/KTNcT04OCEN8ZA962CGWLhUbkgkhaP
VIE9W/YQQrKiPDVJVQUbk1uqAjv+N4wskgl+yi1mULjIx1tDwf50/ukqan6ny7bN0BBfvM8HZu6Y
2njuNfwa2/ov5TBrQfVA8K+2oXIV5uEHhOolcO1ioc2+qYKA5ubm5rUbUGjQjE/qB65yFkVBT/2E
o8Ob66X8A+2IVyfLxzzUA4TwZ0gMpcl2ptYcO/bzY0wwDl0WtSDlC37xXNu54ikJ8WamOFW/78s3
nqpxg7eOs3viZynl1ToDqNN2LjdfzhSTdcniFDKnNcuAk+dAW5Rw/QmOhEUpisyDDA8Dc4PY+BZZ
CzTigRxasTaKjBTN21moHpthNlNEvDgN6Lug/wxLKPY3Y+F2YwDV/quXCVd3MnzvTA2VMOiukbAA
nl63Z9v6ldU/gXE9oaKVgUoIPGPQ6Bs10z4LAWTdKcUiARFexiyoz8yrOdBvdBxAt6qh8VGAQbk3
InfXparEjmdpmFMFFXiFUECQZ01JcG8mdwZBo+2vAka5YxKbm2WHhHoKMa/zzEK5Yrl2Y71zsAHf
RyzjtCrBq2JSIk+oeDt3n5+nNJqXlJ5q4U6BHsCFNHv7/Oe8hYh7yi/tJuDPVJJv4zmUzDIhFNFI
agTF6KiMuiHLn7qXNQJeX0f9iDN+JvJ6QV9NZ/rEYye2jBbgdjErcES6qBsnO4LX+ENUNBlSKYle
oUEmraL15NXSqiJf38Q3hLyPRfRUJU9/TLx8t6Vnr+8Zzx1RStn/CSVKyyXRIxbBx7/rcOIGxG6A
qNdK7X1mAtPHh5+TrSog/DWMFN4SicqJSdhmRqnMbAY8opo2vHe/NlBfuxM0csHqT+4FTO6pUJzO
Tx+dh+7/Rque2dUhDp+tueiKkOcUqXl30mGqzNpqj3THsxnusAkRliwUJKMXL5VZB1kNZrvV6bRv
Dz/zcI/ODggIXFKAl/vdwHFPSZr2X/rO3nNZFJmXFtHXms1eSJgyH3H8etELkS5DruLL30q/6isA
WJvqF0saPOU5hhT99Lzj1bZwdGzULWjq5AwwTMGDhVyCwxqRuc7v2cJ3ZEI5JEulT/dsiRdmeJd3
3iug+ucgNgzU+6gDW0DUkca1iPsHU+mTsXkKNfI6NZ7iuucNLVuR0A0R4niG2uv0JJQWqA1+yNOq
CVJ2NqZHHOoJleopqOqvVbt4Kqs82hjlGo4qKBdfly84TFAQzbZ49jtdarTb0f8GnlKm2qdFsq9n
/FC9V6f+KMRn8XieEFEqiGIprz2fYWwwns7kEnbTufTZGqLm3K+cfbsktAWh0ECtdvzajvt0eeNk
aZTHca8phcMG96h6JFe7AcvxAqIgNi2vq86EZhaZeXskzTPP6IwlIwVp2daKkeLneKNldF027Z03
uO9XurMwXXrWEZ36kQg01E2gonhN3uXVWNNIpwWvpTBI3ATSpgEEqGk8eyoodeNK9H0XYMMCYUpi
lCR5c/kouB0QYSzFRWwSZ35pTnjeEtajMQ0YCIrcJCYkkgBdWWMkXy0DN82XMw/asnIrR09FLSiE
rfMmD/MH1PWLcAmjeaNv05xkExJlTs6H/z18TkusuCYICnGBA4iLJmKFvtkOyn9r6YdCau38YLms
BejuiFTvHliUiiN2pFlwFo2o6q+FStaBoUKw/XDy1jZI+rzf2UA+Rz9LN/Ih+8vnD6VjnorKMBXK
oqtGIRKAPlEHABmg1dCtxWu7fG6EfGO/C6UM1cIB1+mUFPeqaOh8KYbqYLCmWjNPTgOGh73p8JJ4
g4/HGch8c7YoKE/Shk06bP+ISCNMWs6aR+KHA5idj/vCbqsM+0Axh8RpPjGQPEQ5mgQkNpj9Lj+Z
Hpbzb7V00GvDWBi+Oj/9HxDyAAmdCD6XBddZjyv8lR9pN7dZtghuls/6AAKlpM3qINeQcWd13Bcg
az8oENV4dopcQrJ2pXFJ7PWZqb2u+tCgrODewoPKjk4FTv/0Wx6hnqM3FgtxicTABxMxQBSUJPhj
OXzZ2Px6QlCvd/hqOM3nuwp3KcH9C6DibHcd75rrKVsgtK88ZPNyzVvARDyjJ2xzxMPlBvkNC0fi
H0g+z3z2i/0D24+yUPSktDztbYY0FD5tTaJA6Yw7+UNG8gMU0aAVIFu0RCWlGoMvkRKzoW62H0qH
UFf3NPGdKS+Dtrqetu8N1R0L/sObK9EW3rTG5lMINh5KtmpheUB3W60dTq6cT36etKwiM+oJp6+l
lvasw1i5i8vzhZGgo9S43EbYPWuANDeX8EhyCD/bGNHlBrtS7627HZct/QOZmOSD9o9JU0VyDpK0
zjqJQ/tm8PUjujgTUHjvYPEeZ+Xio8iIuvsR+74dM7v+N3fYLgkPTSvHPMXk6VKNnEeI7c2OPsNi
iQ3i7LFWXDqm64FBrIYFmTu64vduRvTat2owzQN+Kk+jhApRdS6ZJ5LArxKMCiSs6bUyqp3cWIkT
E3oE2hnwLdL0GlO0LDjZbvyB2HpuRZVY7KGd83jaTgciznRDT0AXOPL5awH2xnJqts6Ow+jLbShO
vxbFmR9NJp4bc4QqP54V1nPZL3EuUyBUcrvZT5uiX+x3FKBS3+47Nk3zkI1O79lBlxcZNLduWxar
lPRQDGnGn4TR+eGzA0438oDJAyIwuHINYK1THh/iCGtCF3qe03ZLqJcggLSq9Bp1pyvtH5hmiqfi
6gYxzSGLBM5OK6NSldv6EdywDte8HgV5YiSAmSJPm9MBQ1tSySFsbqSZaJ+phQE4aRMMKQqxqndc
SQbbMhh3DmZD07W+STml1wcg9/SKBJZa5wdD08LBvFdLX3BVQRW+Pa0GMaVPCwB+9HItB6c3HaBW
ry2BhcAUl1q1SVDdQ38Rm/5au+wSa7W6aoKJPDLG0FmNrVKri+XPWJGm0qmPmtnNFzQ1h2unJ9nd
dwPjMPw12ToBc/9D62yeFmhJWmN0oggY8RQL+Cw8kCl/P+Ovh5VBGT8KuiHCCaV1Y0OWvOYEy9TC
hrvLRySbcDmaA3zpZBtVKKptmqzExhWrv/8qBsXjs6KCxK4WaPPE5c8xCs/P563/WfGNJUo3s5FY
UDc9J/HVLjfZpTE74mz2N6XffJN8QzP8x+I3RVBVg2GpojbuoTcHyqHu6YKt+vVZSVkKGX2F1sqk
mW6CBBdm+p7TEA4/Lz9qQACFBOxGtxlK+TcKOYCFHC2cK88hHTzHE6sAuwiwldWwJmAYaeDj4M+m
22/SLzY2sn4b+1n9SX1o08KRi0FzyqNpseOr1ONuR4ACqb/uTIVkTR4bUqVveAI3WBMs6E/WJ9sW
bBPtfgv3z5UcOHb2BHdHDKcPq5ly5l0FFCNtv3t1XFUE0Bdw5nGAAiMnuKJieyWoiZWNbNPoXHSD
9QKwYp31gtzjAfcTdE6N6+BcGcQHqvAEo4/AdOazs47SD3UgIKR7opgPFJb0EFU6faaaDOUOpkQm
g8TzEFdCZfP46R8+5LMSnyzqISY8pkNfiC1Ies3KjwFfU4NcG1NcrfxHmS+HvqguGI8cCxBruoxg
exVq6S25TLYUSEHj8ZucpIpvo6lr3FAPAeL2ptLtISHplEZSBZ3KRD9vnEkFasREc/9AzIgZxPFV
YORl8DQkoflqUsSBUlURtcLSxwMPIa+GopB6A3gmUyiFF7CLYutxjxPrtmz4CkRjTNu7rUGQZo63
CMDCE2XJf0ECFYoF8ybT2OUEriviblLxhol2ownOZpS5R/F5CP8LxWUo/WDdYj0qo32PD2k+/dQh
cx5BDSodwu8FQFD0P9vSRDB3HfFIIa5BZUihtQJpl0OvY2RVooejVJfb0A6GsyMvwoVtI2icW7TM
1QT8QFR9uD6vrrWyY19xm6hHkIyktEdvooavyAF3Gijm9KzhSacQ3maEAIwhM5dVrNGLNM9oASS7
cBW77R2HL3UXCBVGQOJfK7QIRJDQ88sbZ2OVpHxikjNHxrwFQPxOmKuHmlK/GZlJdSCvjEa+9FtB
8CEMg6JBy046Y2pBiHZxrFEqDCx+P3V0Cvc5KjwSXWh077igB9BRzmRXsPwOWVw6zjWL488xngLq
08dwNrbJbUl9a/tzkrUJxeZaHm1Zs/+pc6Eb7gBk9XYN6BMXMg1chF48rrNIRhQQB36+tBAoo0z/
RPV/fntJyNAPFj+FnDdUovqIrALlVu1/uPm9vgy/b2YydQ8F6H8oQlYtVGyky4dt2b927xB2OGsN
yXnOUvqeOequwbNnkji23G6/awpAf5uE9BjrAgYz/sFu5vwfFoqF6VgK8oOdmj7RLgiVD8qHvdb6
iciqRcR3msTYigtkalxUIroV7O1rHvjFUDQEY+FpH/4CQjdfbqFhz9YbwBhX+2dLQHlyEgzs8vuH
9gCDdTqwBzj2dOSx5GJO/p8sUm+8NEOWE3pR5/uO5NnKghw0yFN2KHj7zeg+4LzUcv8GaydpZNyV
V6wxYc8bByqR5gHPJfsuL57Pffl7nVzq0KLEjyZ3FsW8Eq4jH52tJBHrJnlZh9mwOUGJRTWegiVm
Bw9dvEyB+9p2H4cVNYPe913MvJX2biGG2LzosZyXRk8pyHXk44DLlhgT26UbzGmvKKswykNJrwzr
EZWjSYv2FKpQkEOtYawOcsTKtqdtnQYXuwi62bKr+ofPJuqMe9vSKorFnK71CQr7CXa0hw95iiIZ
koh/LOBA6m6jH2ds0gh3Qb9quQPd4yCuHPwWo0RF6a8bO+da+uSCvhwMbyA4pdAgaUz8ovBv7Wfs
Tkuji5xWk1HEv7LjYoAd+7/wK9OwhbDisIcKB7wR1Hu9yCK68rnMMwRhFCtcYkTqNvz7UB5Ax1je
ZtdIv4k4duKBjEYOb3d3nNzlC6FlQ7fwtCaQ7x4CK4GDN632uWmNp7ZF70y/fnLXLW2Dfz7jqLKG
B+gfmTGp7p0nwaAOB6SdR+Kh1FoZzQCxUkzZTNfVtbA3F6ymF/ppX15+n1lf66TnMgPbnY/eV8tR
yuTMJJPvC8hdbz398G4Yd6ybuJPjIpjY51DriWb2D7bz0idbecJ/8ZzffdVzGJCuOA+hMEEatrgF
JZHC/wdkdLvW2RIAO1ZKLWdoexpsavlvRavwEln7Kzm0Pwwo7nhesKJc71pgsXQr0kTg1rG0bWdn
T/MitywuW+S2hUfZAgn1z6fjuK+ijMuHzXtChAPLQ7lH2yACWDDlqa1zehUGgCvop1DNkJLr0oHD
nWHQadZ8GnjOThiE83bfx0gmOY4AG1BxRDNmPTKjtg/BVCEzmcJW9c8mRjrqhZm70Kw3SQVAkx6R
rgCBnikeFlfI+VvjKEmAFXDMNCj+f3cXlQ5v8PaIr6Ez5VA/bVUs3Y0pjCB60NibBy0IRZnjp2P0
UOsABi7LeN1ss+xtrek2QxjlS+ZPcO50dHn8sSOK9qoLE/FLW+4cwPnwY7XAf/s7VQgw+z8o/qAy
Edu/Z73tDDlPaPNhte7JVbw2K/fWOyANI2L79N/NaxK/2nWcq4eCRKd3why3FzvcOkCnpOgdojB1
fw7TggnzpzOEZEa9vMs9FcnEBt8jo38uEsFs++yAAzGlZ3Yo1VX/5FqYXXtcw2PLvauPSk/A4uwf
IHE3OfGKpD0b4FRvOS1bYsaVeXUc8tA7RrKZitFBYdrYAy/HjGrodCnlVHAuee0xuBxTSUZObpK0
46+xMQAphNEzFfPd/wddOp1a40PRnjyl8BKh27BpuaWbUWXIaLlC67cgLTlJRgQAQWVT5WZBLhJ1
ZPY+Li90O1sPPO0KaYGcpjVXc1bd6dEl91ZIXBiQRH/ZXRYzfIhT/rthBtMniqYvUNbbG+YScnSr
2hrLHg5FYU3+r+8vGzElOpZB/CppVZZSqwLG9zZQlHZ+x7acR0PVAMEbbEUFybV6zTFmRo/TEf9m
/UwbWOzPELTPM4oJWxJLNvnLop4n2i9LA4K12dr93UsiVkWBqlypOSkr7BJd3cDVkLqKl36ly5P6
MF0c9cRRClpdB2YyWVppkueny+2BFtbhrWxYmeNB6H5g446unuj1Iiu5y88LfxAL2/weHQwuL0Fn
BiF3BEAU732hy9hqhAag3cyNctwzvgoSxZBpX675eSWwfjjWDJdyKatGKj5vhZ/BWhDZCYCxF7L6
iOAT80MAogzjVIcvay1MRgmYML+J7y+Jih5+tsr9UV83jH3/VfJeUelGSh9w3sK1c7SobWjLe6yP
lQ+QYhE1+J6qmcEg+ZNfUfFJFOw55FUq/138yDQaFtf/eBJ2mPJiL6Sw2W0bbD1jq23y63/+afu/
bDsZ2GRYc0extDm/zaH3QdirBF0J8W5rib0p+V82yyk5KlzvYCYq9lqt47sCRug9zHOyxD3tzNKm
7Auaz0VpvpuPoBGUmwBPJRkm1gH5/RqpvxMMjt/86jbhUvYuxeKpRVXEg6fTutndcqHke3wDVAzL
7HaJh+Z2pdtVkPUDQUIXTFnAZ3zWIFr/J3pSo6DMgvHkXeScmlpwps6B2vKkNPbeO0mJahJmucjf
VWM5NJtEL5wiV+4yrJI5ZbaBLhs44wWk/lqK9DfCvyBZAWh7A4yoRzQv7RzsI3+Rb5fd2PPpuNcz
oyRAc2fneNfKehhJNpVkrzwVjYUg8Ej05ZgFpAHJHy1HUzue6JZBFWPZjU/cgfS9tiSTFvqLubFH
ADf/MypoM0YUwJyuBekp9foDyMFDe5xtrkcqKNFMXaV4zDr2OABvaJa/fkmb3gqFCGjUGIZy9H+j
14T3KnLVS4lxLej5E8dFM1q4yZJq8rlb0OCv8JXEw+Jn09b9MvQg4Yi7Sl2tL6/I73YX1kxOt4Re
K6n+UET9UUEesR45lmTEBG6/8pek5kqoi3cPgV24sNFEvRpIFvddX4r0ZyK/gnR2GQRwNVciQ4W2
cKcDkUtPL+ocvmF9w4zKjJypcFKoRpsut2De1PcSMwMR7HsBdgIOj4MGQcBwj9j1hCXEDOjrP16r
yRzST0n/y4dhZ0bKeIruDPFhZzximOvZ4PakJBMAnhTqBPWoZdBKQZaigOnJKKekiGsGkYsmXjdB
Qd+YeGwGKmv9yVYE1Sxd10Vrp/uV2S3T1cJJYg4B4A/p1zu4i2kKlj8HIvkZKbhxvRqs8+i9+4Cv
NdYzrbJMZ6DvrOZ0MRW9d/7N6BGtwucVJTAqvemRwPQwhLlCTHie4CnwQlR2MIkTie98j6VVUZfF
n7RTGEWLOTo/nVXl826zfVOPl/Y8K4xDdms5alfISXI4wJk+90NV0FobLPZCwRbFXGWpR7RccBWk
/IuU3XQSsIDp6k649YWpF2xEdJob6HrywevzLLbfR3J51UqQjd/wSn22Jr7dW0W2lhroTfKyarl5
7jbDFB/yrfLmck4ikD3AnRrYf+F+5xQ7VhWLOF809TIsse2NvRiOghlrDhBEf0kjfeB8Ds6EBQBJ
XuJL1g==
`pragma protect end_protected
