// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DSJOSvSQKL3LYhVypZv6JIxHtqQsvq6TUelBsPlD5xn+sqzIWYWUKsv0ui+xBXyT
p5vR2hEoD/+rgdEApUDCgQC76HLAh7QtJV+SJYWzKRI2nZpxt3ooKm6M9z5mCk1I
ox7tcvTmgOFtE48qbfRNI3vuitnWs5onX8QeICiH/Ns=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9168)
nfjP9/SnMFghM1Zbi1daM2ZQpOU34AvH0YIaGWuVe/VG/IQMSz7Oy76QFT7JQzLC
DdmSZHkx77H24YA8yjCMiC0LemuDYUlu6/5ZZeoPDzyLmewXNmd07ow6v/NcYKk8
w0jUY/1EVc7cn4YPZCY71EUsM62dLeMyF42HkMB9qqdTYjla5o6yHhybmUvfJo6W
l0D6jsrzFlIdsuM29JqTU8y4bFfhg6jxsho6krvVlOgO+74hIn8XgIwaO81Jifhg
1HJ0vXcIYi5qOI26shEQNWpm1mjhl+LDjLgpopkt762hBZXpp5Qyz+Jpg9Lpcpgt
JOhHB8o2cgaIVymaSbFlCcyN/E9sCTwFdDQb1GSfNhRbA5NZIKlUZ0UnF0gvyec1
ZSy5kxyg3Dp0IVzTzYszYIglDPZLPHwvL61sI6qAn3bfsQGsnQufDABaENtb9ydO
rnTejVLLSscRokNnpkBpl5s9h+HoxTFWQB0o2mEGiQPNRXzSBl2QATzf1+Wt2EwM
SiYnAR7bZblZLBErk1BpaHyaMKnJCg7sz9iNTZlvghu5o1+PmOm+8culNhxVwX0i
CwslxzQdwsy9iqDo1fRFhJO+z7Hc4RkGaTwpGpfmm8Z35QsiaLyn/E1ep6oTazvW
p6jQTqmG6BpnzMCnOZu+O8dtiNrJ5gJRsh1RUsyue+CIgZRuJqXfkXuBP9Btlh18
GcGV4Pt1RpH+C5/r+TlDPnW3GRg/AcmKK740MiJmpeyrOztOwuS6LG3otE4AAHh8
0tf54Qa27InDiKyC4ao8XL4UtFwvjkIK5w45IXq0hwbWz5crrNdiTsi8LhY1+24a
N+9ykpVKQJjyJWURTB/9QKbw2wnN8DhfEcZ4qsOlHU9CsUsNQJZGGmUUP9ikXb4C
6GYO17Vp7K8JpSdI+p0i4uOYdHY1dki8887bmLlS0nEDpRvGYI5cB+kvDHpny32A
1N+pZTLzhHcS6Uk1Nik444leMOPb3SJEHQTz3Dv80bBvKHDSzI8hukM6N4zse+AK
y1+YkQ/pd9W8aJH0ZycsJpodQPH+SRPQURJgPL1Q4bATe4v/saQ9F8K9h0pnlt9J
BjLt7R16ltCUcN75aydBCaoFtFo/OhHtu6YM/zGUTo473gPRl5a4BEOu1OhA/sR3
jKtU04vJzWfpm3qBUTcNRQmSLmzkuTfIYN8q8TQET2ghIQEglaK9XqZ2UXogdKXN
cxmcy365P4R5y4wdNKyP7oF2Y20dXQRPIZh2srQiliAqd3IfBg+QnXL8qIOSmHXw
oI9q/3+2TnuuRfhljwBi6KurnbClZmtksWA2DfoCTlLQgKd5NIBcXx+LBjB6pP2Z
UN/vUED7ER2gRjMo9fnjtaC+5St1pnZx/5e0re1Zo/92fleGazszXqDTfWHAe+ob
sboio9ZKEGJW4WJ9EXDZRfA6/d613/qHmjeYWHVItwReuktbDWelocf7hROOy78B
q2bksyxP9L8DQiU89OqqqFa5lsicOfHxJX+0gfWInwyv+nLXbO889+C5Ky15oEQu
Q79+5EvJxual+06bmfN1QuXneoVUdshzN854aN3Y33KxAiCnYjPoIfJuOTktZ3rh
zcn4W2SNPgIpygL2fNV+rlKCpJ2oadUtN4MzxeCz60cDbQmFuODKliHDG9GN3NDY
22tUUNeWLLoeezl0ZV7P72aBmtmUoXyD+WmfjG+zM2P3dNTz556JYIddQsdwu/h+
jiVT/vA0oWQVVxoqf9rPG3eYl8HfLgikBQ/HBHTrUvNtVVNyd9XdyTm9xFSrIN/t
ORCM4PZ2e6LnV9Gi8grPZVMPdSweX5GJMwUw/wunNMfGdf11JZhjybfEeXFZII7g
f30FWb/VDWZx7qLBrJXwquXEq4iTxt1kqtD2vCyhlPcuntckgGkxBA9CGwlNXjYo
kQbLbnmHLD5xFHi/VAi5WLum800gamyt58hQiJ9lHHtpBxNwub5c3cEujdOpB2Bk
cXMKf0hanVjpnPNkA52Z301hYPERhUsTlh3oX8/t8LQjLwWmmOCN2E3xKVeXEEUz
TI5auTNNAR9+XWm4lkQ1CiaEXT07CKjMAh1KSzHEmqolPTNWB1XTyK0Np6CWqiRD
ikj0waDYQn0Fz8hC8iPuHqUHFK0s0M9cw65sD6XbK37LibmvfbHJ1uwbWunapRPO
BVYPdvxyJO/740HBT3CQtQSJpf8DdnxcQCldkcEaYfPXSd3fhMdnCI/dXJBZt7c/
HJ+H/Nkn96bDmzTHmUEP9sTzehv+Bgzs4pfjQYMv9YNzqCz5I/wvzEeKDe7UVGn3
H6les9D09KNcJtgnhoTni+Kk+WEC6zob8R5bvM4pUHPG07wjzCwVeKqNtRZVmxYp
bVVOyL6WYAy3AkVDq0MI4JVLPk3bafol7iE+jpg1tPyPvAT7xzl0bZvNpgaxV9Lt
daQWUXWa1O/eskudlmOI2jHYtmEa5ir6vQG2EDCUpy+iWYoqO3Ji3JpD9xFIUoEM
dJg11cy+POXp3QIpQ5XY5GiZPsOh7ODN+voA07PDmm72ZxZ/Go0MeO5vWA5SiJNz
SIwuvcTi/iPmz9C8gHnpr2++DYg1g5v3VdblnQDyUUE5e3Eo429q9TkSKmsqqmoY
GLaZZ8COB3LngnR0ypCC3RqwImzodUm0sdfBI/OARic0QxRpnXKKx5yQKkawRk5h
tpK2VksNBJRBrndJATQBGm07fmODMN3ri1I6McyrO4ybl0hH0kLuRD4f2G50ktxr
9IwxhPJOb6nW+s8o+vwkK6+UuDuHJRhPdin/+nwLGFBSZZnV3AQdT4wFzDzLOFFe
ss3p+ZvnY1uB4v2veGc+YY1piF3WUt0XzgByLDigX5XWJpTBc+EaYznbdD8iKZVB
FiQFAILo2sZLiPnj8NmbyXcLK93OjGNLxbrsMOWYZ7r0RQsfEwyYktCePfwgYWyK
CTYlQTLWAi+1Y1S2C3WD5p2+YYqx3Q4xSVSYDQ9jjkQelxR8vBSm2KVeERHzJzun
24AcqCzUu+w+x27gr+n7/e7sXBKZ3HA//MlpXvQ1N+32HkZhmAupx5/nqVIws/UE
6mzQUynRZMx3nlBA3BDgeeA1T73hklD5dHZp/5lRcBA/FV9FhMJ+P26IvF2XVHT3
iz7WwcQfI0xjCSZmV8zmsM2FhaDGoXEk0YcnjggWtZv0DFl266/zwXap6PEhpF90
d0P8GsO7EGgayflaNr4Q+KiMRwrQJ8wWVrVjikXSGKjyOOb74WQ2WMlSQbXzSjq9
rOOvc+at/eJqUMF0gMRFhvHHJ18kwRxURLPI5REt/8/7RJXOMelx1+Cd6jkyCRqX
iaZ6JWppYPdAuZBzTvab6A2oUA/VuQ0i5Ra01eAmM39jwnFNzwdmL/YzA8TqXZYb
m+8JYkgufXYDcoELUC1/NxfDxnbMeuxyxa2iYhlKaCnxXHiqWIbAF29YvDQMet1s
knyJswdJzQzzJ9pbDTO4QqDKnTzP0pN49Q6zrMMznUouy+RDay9xWhTJH8xk161C
xzWnfoIQJkL6djgUU8J1G8hkwPPOIa1NV98rm2KjVXitcRddRIO2iXfGXk4DexQA
bpK30SSjhvfa8UTUT03+uu0qY7Ke83O8jr0FWRmTbP2UC12mGkeiYnNHrfIc1046
/bl47KyYMPd4bibllAx4fcfSw1Fsli0J2iNbsx6jSf2kBm6dLC0z7BVJSLu8rPmC
MnwtbmHBSZ2QGgxVVz2IOvfya2fObl+KIcgRcSBRRZHPplXr8o3B5VPerM1UFPJG
c5WORgVz/Dusgvv/7Y2KpwQU59gJGdZbMVZ0IsWl7H5B8CWNF7e1aYKhs+f3+bH/
gRMoa5vl/U3xH1cOG0SGIw3dBc7dEkP2R2euS/j4sg8ZbWbySm81byhY2LZCq9B4
Ff5ITcso89YsOqLIK1ombiaBHMJ9QD9V7T4EDY3p5uvtZG8jhoABlK7W/eOTuuvt
WZ7TQUhyVY1HfrrsC04GxM4hQ+re7oH1ut51RWD+dOkfsGg6/cfcqXUsVH925/fD
TRRVONxj9I0+6xDySTy99w1+5+bEsq96ToJa9ml+QLTWOP4eZXFybVl2Aq7xdvJh
kOyJARDF+xNGnOAyPCpfBfIQr2izYvcvinxaLvVouXXWB8QEN3PXBoahPTFMGtAL
2pnO0XrGJT5aJxA3cwfpvyV24cWSI+K19BXjyDowgZqsiDlAcrJvRXzZdcncMD1c
o1gRAxkdJyjrYJm2gQKUw8sOibF0EzMWDlaJqT+OnIeYpJDc92kYcTlMK3heocp4
80fqtbOGZ6ALRbDPczZwX34hmE0XnuAtKd4adY4mQCFIEuuBjPhW5BEZCAz/aHDc
IeodyNFFufPN+h/nNsCGo1Gr8f7jgPjTJhgsnqAE1YLG92GqodM1deu/U/9FtUhv
FZlOt3IWpyUvAKtW7IS1c8wVl7OO7/Q9STfHiPQ8Ez0bCK/BLD2ZEC3nGKHL8N5D
EC42vmAdtSghBt4eiWhW3bDDJZmk3AtvTvo7e2Zog8X6wQEIx7EFjScJlh3gqeU+
T4ZthhZQ7ZOvuTvXS3tvQuDTnsB+i4HdOZfCQEa4sxwZ/xueqxOPSHOeCnLHMtxP
4eC89z6VLLJEdahzoYt1Ga/H7Jr2m+O/9LZW1y0yO2yUs9re3aVtoooQM+MsEauk
/Bssker3FYNxjBC5zkMGVHLc9+E62BnAbhXKgcezGRaxiErtK31Rt5BZDbFSdx63
3j8oCJbDRUKBV8t5kI1Sdv/cfNUW5/KTV1EhQlWk6GWPsKHPqU5PpYe3W6bPF55p
wK3zowLheNvhUxyARRWNZ6RhQe3lLaF6nXdEB4zNAG/4yKez4dbqqgtT+JO7m7i/
gUYcLA01MGRx9s5cIeaIt9zvZVdfhNMDxl+urvhTlKs0m3N8vNCF2XoAX7ij4PxG
62Y87cRz3bE/f4RnlDLSoSCqFhFHmKrbylcSaWytcO3bv3WbXKIcToZRahtvD14J
twe+tGueuPoyuZAwt9ALm1md4Yw9r5r+/K/ihFrndQ2g2EjSNP2+w5SsjI2vj7MV
C1ARTkdEWIpHCciuw38H08mwhUremifMxxOr8IJRQLrwb696BGX5fbVxyUCQhPwx
pr8azS2XBJPsGvApqakgAijCvUAzvXtnRsljy/zWoAHW95I8/NpBIGU9i9pZFaed
VXAhHMZ8FIAJJBr63mSqVemAHfrDvjh3car+IpVNY5Fq+2Udxv3NzQL/BMUTyHBy
OTEM7h1bjpqAj5kMrN58Pl8eoWgX2QM8q7TKvBnAOA8c7CId972/uFgbxBc6HVhv
QkjlYhqlEAb8auwnVnhSdt+tZ4H9q/E3M1DnYuNPlb2gdHi85UT/juC/M4XqmjZu
AwbrtnsAfI0F8g47kXSu9j4K1+c3eHv1Svs5kgpy5j1Iiaj9UrgrQlNd1HXjLmbO
O0umlvy+XyVtPLxyaIZ9t3jTPur7moVmfX3IuKxr7xutWQS0REo57f+xDxZgw+SH
ss2b0Cl2rYHz9Fw3bixksAL86TIp3Zf4dVN0t+0WCNDrCfvQxXgo9593AsAmw2ac
z8TTHRAEOo1bZDyeq3L9l72pmg+Kxq1vZy4/LsZCXyKJ5k0Ls0FIfstNb3X56hy1
FNc+r04xRFUxM/hTwH2bV22escbI35D3j0a3lKnm1QnP5umydi3zj1H/+j5LD+rr
jD5jku14YWRTOEWdcJXyEUxy3rcdvBRqMY0D2EcbgqibQJUI1ErlVz12ogLD7Vjb
j6uY1l5RgeOxX9HyL0rgrfwvm6t1eJmuW9+7ExsgvixSHVVrTepmcxl1qX0xUtVy
7Wiab+2+vvwHUUPVUNLMnX1emPG5F4ds3Us3OikTjRClaU+1Cc8wxQgUMRNFSE5v
mVfKC4iZnPfcmp8yGuKbdeUfWkLf4oPxIJloYDx2tvVZWzjdWp2Jkk+6NeykwmtO
vfllvr4h5on1y5Y9wjOEzUsUjYOmAtFYP3QDXcZGZk1eheDv9/w5oR4rXVch3ENp
FONcR/qOUvBVSgA+F1vYvAN9yUQ+kYNknTzQv0Qkg6VbLTfTUM/T/1nu1ykQXnAQ
w+CUvYDT2DoO9C9equ5nQo3UVI0yN4UOSH+6RMcW/hG7I33+gB3H+QafOsZ/oosv
6j6PdPQsCZ7zHWf+Pq5jpJhMmqfO6a9IgLcu3O7djJ3urf9oTau0kYmS9itkgVt5
j0Z5Vl9cRJBFwZRqJvaN/cufUAnQQboX+xSWRBmk3RiaEVCQixgCtyyA7Yg10ekw
zuMR65P7q5QAZI5+zK0PNYHEVdaTIBh3zuz7Ai1m7Apuho4QFNEOlSciWVuPnY5s
bHBoNr2z7j8xDw82sxfyyFEtc8zASae487WzhPoL/x29BbdRjZv1psErNzj9hOhf
7UEIiCynuAPRDvPtOGG3YyXPZ2DxgwscD85xe5USnK2qtKdx7QGveCTJo5CCBNKs
KGzPMN0VWo4z8sfyR0G05C8roxtn8Rdk1nA42qtvS6iTn+NhFVgVMDFl9a6Uvvw+
pCoqvEzKhZpTqtCEI1dV6oy3mirfEU4csrp+NOaRNWIeFRu+s/ATnmtiirj9yEjo
scZNOOU/0c7qM4QjPIK0MIdtQEHnTFVfTcBrlM/xfVlmPEE3WdLHQMK1CH+5JByp
kLxIZMNduUQwiaSGjQwiuVVwcBLJu3cqOa3bkJX8uY23kCRUixzXhOIOoG1BFHWY
On4S/0R4t3hmuqD/LWH0xqWiWwg9BXwNOo6LJYwuYpor2fPV9CbxNLeeBqbTVQ45
j2I5yIyAqTVSNDhhRvTDIN101wovLk+qOGuUSdC0+3BUXKKaL56299SJuL7CqXgG
F3WUCtkLxJCZL2vgzSBsDFk/Gp+KPWa/t0uwirycMl24cL7NGRdgC2pNSjLlq5u+
b8g7/ov86FSI6OtAIrHX+7PqjXuHQQZ705AYCw5a7Q/CNpnWixTkc8AbvCoIw4ue
JhLeum5gPapZwE+x2hiK2RcXnQKePHoNTSX40sh34XyuVLFtxUg5yNSAiFL6q/2F
lX6i/pydrbacJ0VTwBlvLFA/EBhXIQqvg+l1kZ09iQq06OXlJXWtKE5rl5wIgpge
SioPC4tUCZ7GC1DiX/uKcwNRhuDGsnaLjUEil7rOaAsgpD9lqg0PSt1i3+yc1g+/
9j2T7sCZi5SC4xgJeGnGovJ8HBjoZeqvi+Ugu1IU2WvSfvXu5eOpCoz3miXLs3dG
woHbU5D0tyleDkOYQIkXPnNvJSWWCwsjgRUhtclzG9y0Bsg4uFNHcks6f8iJVnHA
n3Tt3MJUFpzc6rS3Z8vEkFAjETMJo1wBAYV8pPWsmlt2gUWKPisTzRbzVucVaoL5
+mTj/FLzpe75yZXRS8SuvRzUFpdaV4ZY7o5A7gMzkek9oyDpLWpAvd4DF6TxgcHy
I8b3zSqObHmgIE6aRPcHHsFjJQHE1ib6YOhbSKo7y7ayWWAn+M57pFVeP47E2eJ/
x/Zpzk37+FI6E6+iACcfWVSXHTyV9V+33s4FuLB8k+qA3+9dNLKmkiiur9EexOd2
gbHQCBawilYXLaTLg1hEfRJuiD7VYtS66ZEEcdpFhIy3ah62YHaH3uva5qAR3oC2
C8IEVhAiKOr9vKz3AXG7m4VDKGgbKruaB5xpU0S2SqpWiMVYJVxal59t3lmeKjkQ
qd0eEnBXMZTFKBBPAh9RncsBMY7vPAGelhJotJGLwL2HGBX+QaouwRtReCT7gpRD
sx4+di1Z6WFBUyb+M3qqn93WESUMdhNfrbE24iA6/yktCR3tybzMU65wpf7C1v6q
q6yqlDQXKfoJz4vSbWTuLPEwexHxv86l3JKAIc6DYixq8eatB8ercVHfLbxmEPyE
sZHPfi7my0ZuzMnJqcytZNlBcqlnwvAUF6D8T+hUeji9rQuP4umeqDKxGQpfpPpJ
YSVPseaOAlT8Dp0FrQYDVjISIVAH8hZcHehZkRD5kefkF3R6ZJRmdqrijpc+W8tQ
x+PV6xNkpllvc5pCFWJnyyjm144hB0Tl07xfuWc++DSKf+wblzAKixLg1VT1z5q3
oyi/q01vx+2yzKthlC2d/E4552OwmY+tj+tVdavILJc6PjuNjAggjhu2Zbyhhuvg
9J3HqpTPlq4vZmgDElFBAaCAl7zL1+9yGrkfeyyBMY+kgAfXJSTS8maUzpwkRX2t
lihe0uUUIv8KxnqnIQi9Q7dVUbcrwv5cxU28qBk6cylBpeNZbvrB9jPogUPO/eFj
P/N90mqLfgT49XIJpohpmtoaBQ+XP8plJJQUzbNI7iF/bE4HAjWI6cqJj+pzPikL
kc6Gs/pmy4/k3GSqVEk6GEC2UNHkhW9vNy6iwpRJOxSt0GUoAdA5wMReEMxiBIyj
itkO0X3ykr/3JU9UxRWlFjt7nlW0WsI6Qea9ZV5vAI0IZ2QV2Rh4NnPXrvE4vK3F
+eP6DfhGnHopt1DbWcoY0pjhdzhIwY7MRQa7RtL7GaTrPfaOrC4Y3sTm2wjsB8kp
MBq93O6teW7UrXns+QD47VqKdiusUcJWZILQP+BSihvabEU3dI5tgAmO/NyAdmfV
5KCj+FPmKKKCy8uiyvrDXFX1RBcN49p/QzjZh87LaePRAgWVihdEMPI0vb0SePms
DwdeFLN44ODcTux9bVL0enU7Ky1MV4i94ge1xZhiXc+m3S9ga0kg5h3I/PYGiSh8
aqKyTws06EL1YxRMAih+deFm8mKCVO+WzRYAbYlsFn3ogLt/9zgFQp08mejfaPbw
j0v/wcL97GxA9sFnjor6oQInHpYEE3xhq1bVeWOrcFmmZCbAA1XrvS0AfQ9sNS6E
QKAIKXd7CN6UHRV4zck6AfbaM99x3H5kW5cuB2q/uwayASPuIS0W87jY5gUykkS4
6z8l/vE4MPtM8b2Yg/sPIDksaTR/kGvRrgN+RTL7Bcvc5ryrxzYBZxKZrFR4eTQx
Ga31a+B4ZHtdgjQsz8ETxOVaY4WL+ZZ/wuv5c6RE/vu4nIlpaqaA0lSX/FzgZRXU
3LgFyeku8H0Np2huANpjzagensqP0p/nJBQ+easFt0gQ1cly5R5LlL/99lpaHwa+
Vhm1dkCQN99fMVvwBUcHbgKbsxwZ/wYLoxixjihpqcCrrx6zaABEsQztL1dBZpdx
hvOK46wqz9BuwTESFdOcNxQGsns6XPG/5XgH9W4jnenMoxSNZZwH724nbjaqs6U/
gtXNVYVFS76foYwv9+kexYhIjyEkbj7KNmPtE/L4F//8ZfAMpsRG9rjkBm2vUvZL
BhPNn1DrH3J71lIGcgXujo80NyzJAD2UbY6yCXGzim8BUNbB12p5lVHPQfSF27sM
zaZcb6TgVtZDVIDqjKT98nOal/67yO66bx7k5YZW3o/FSNyPzUasbHU/a0PElBNN
q8AkdxotnJ/Df7gi+Tsd0/8jDfNxyPr2HSdZPdN83hi0lw6VxwnQ8nzf1rChhHce
tzNHT6gcV2SoyMFH2sUDQbrC1oIj2KtDDyVbqW8SfjYNOt8TmbLku5L3wdpO5BeI
vd+3NwAL+Ul5B9ZSU0eS+eHjGNKfQfX4TRVXosjHTfNQLDoVGSkM4uBiZpw+UXA2
9hMEi0HJCc1wA5POIYJcHwXNxNN8mtXrM2tv2HgUrhBPBQuivBDc1Ti7MEvGXZ5M
aWfUX2tNKfDgq2SNiMsXDF9V2q2uO1im3XPJshFYwY9eBa0f969/WEsaCoXGh7W8
Yu9SOO3/a1OsYEiHtOX/1YwLbQCMWkvkptCsUO6vOmSFuP2KrDEcfUnw7+ybQkZd
v730kaOY0dp92YKhxVNlup8U2GEhZvM97+UrzUnkr7bHAoY5mKh9k790gSJTtGms
5Siu31nPrIExtYkcThLwPk3SZRK0jbFnhq3PT1yOeHK7AR0QFWo/gNZ2+rycqnQL
klaJwdXsJMztOkzW2/9tuZB+hihsVgPm1pIpM4l1REBmTjQ97rrlFTt7X4foF4xJ
y6wqro3IURXTfZFqHDVqbb4WFESiKZP2hD/yQ3KhFvo3fpJrIHcHJrF2f4aV74BU
R9g+/z+/wTRKeBzzYSO6JjX+sWhl2f7y0fFi64IghY4c4Tnnt25Cg+S6Ua/7JC7w
ZZ7FGKBz0XCCnALw0XR8pK1HlublBShZtYj4APFUOKs3YepHExSEp9qF6C37lRNA
Y38I0mXIRVo3jnQSal+0zUt6QyTlY3uGFrY5kFf6uXiQxzGqaLb8vJxyewxtj7el
sYiCnyI2dTooGHs9/3E92CIaoqxtFkUbn9lZh8pqxHuZRgkS3p+8YUfDVPgYgiUb
Wy6dknzzdmobdzJx/vN5Kr3lA91QYZ4QOtrjpBKiPC7zrWgGbzG9t7nzRYeF4rjQ
46OZu4lWv4dwJj06TypeHj/URLOEL+yWdw8ZkvuRljXgZxfHbkgtX9cHM++I2ndB
z0NTvSo0mNmUaf400/9ZV7+nYAsKABE7kWlWPwjOOca2Y3xKKtwj17BXyWt1ovYo
hIw3Ud7XPpo4CdIVDtGpnZ2cs79HIxmY0mVyYCeMcQ5rtXBMRy1+ScGqNRH59CBi
z/l44/vyYGB9hWVIVrPlLi/dgvtdShrRpVKiJGsIF8+wy46LRRav7y4sw4ZagFbC
E0raVzEavVFwQ4FeXaBjavlF/AYGEjzBpkLLgpOOOKuGUwJpkHvmLpZ43aiGE7un
e7giG3CRNRL3Xdkh4GY/UlshbYLI1lchWlK9yOfZFjJG71DQSE16Az0TOugDI/9K
HpF9Q65K+1uIL51IInNN1zAiy1DkzaXI7n8Ix/9Z/Qmj5G0YwM043K7p02Y+fUkS
IiCkzac182C3gu3970AAVUq4zTQayKhrGottzJIySPtzjvZRPsh8oldEo3a6pzpx
+DEiCJjgUF4xg7K/U8XmDJamyUh8j3s4qLMWK9BkJvdg6zdTB7XhVlSrlIx7HlaX
BNxrozWH2QDIMzPyEW+NSUtuxUo7Vd/IIjee7iaYfRAMkRIlNYozE3Q6XNvpufh1
iwXkX074muFfIDSk67PqPKuYDW6EE/ks8eOaHsy6/qfkWBf1tljLDBzKV2Q7YBnc
QA/hfSl5m4/Zf3LmxRzoosEj5cRzF2eCyj8+164s8fX4MMW5221NIcLnnkLDpQce
AuSdvvrC0SfXOm+knZUGN36s08Oc3lkfXkOCMHTecMxgslT9XTAS/ZvNFX+kDZ0U
sQXeLEPHsKd0xSoIQy3VELLHzl5GSwQyxPmmSDcgNsjqbAIF1Es4t3FYtuu8cb7k
X0vJWj7mLRoDe2mpS0hFvF1+yo+m/5ZcCcd1CizDgGY0yTwg7TRZSj36KbPdzhgp
wM6E4cgjWuqJRBGxqnOiK2/7gGZpLsrOsNUFOd4qrPt3/DICUonLa4nFhh9OQY4/
TabkbdyNqozpjoJ5sOrCW89UefNSD39QKqWEWcRmot8meFP9BVQlegHJKsvzAw+g
s0Zum1lBuaKJnHGVLnSdrVBAXcBcDWMfWoxRkt0SrqfOBrJaG+aQR+Dole0HJMRM
Qgw8N96DNfhPdDNVgkohPuAE+Ub0crJFoWcVMBjo7dG1wHEr0mpvJlQgwN5ORSez
CoNaixFEF3hC4PfLlCemeHrq/tkPDnZ3jnacoT1nnquR9hBVIFrTX19muWe/ZMKN
xNfoofOf6FxqF3CxYioNIYejRaoBuiwd90ZxTweWjVeLqVK2pdUt6SuUwh7p08qC
5CxB9vcpJcZPeUf/bhic7B3E9qajzj6sRqKdSRftZOv5bFAZJnwG19IHbT3scrqj
Y+XS9dqHymQnhhMfU4PaooNapRSCW7SQeGYKMLDkTxl1FBK1ZA8QUOkAVt2NH3YC
MdI+cf3j2GzIV91Ti0qC8dM15LP82M18PR3mU1wThbE1vegitnXIxzbfyFxrvV18
jGCKffj8Jo9hfMLqT5j9dfNLEgrUKHJmDjPfs/VXKCMSobh090xTlEepoj9Pnsa6
XAGpO0TlyfJxocSiuSCL9PgHtWX52QuR9oMA2DGAn2oT0ASw06anbPrcrZ4xJ/if
a5T1Amp/vG8sQ7OJQtlIMWigI6fOQNaV5XRK/xHP1+w0V6ND450R44Tuc6XCo59P
7J8tYFjNyXXq9ibLmC5YGIgd5b0XZ2VoOa7efDtu1i9Q5kVkkalo/4DntUHmrww3
otz76bXQJDY8e8Eh92oPLonc2PIoETUqhC22KY8ZXqQy91vkfeu0YXlYtIlK5P2R
`pragma protect end_protected
