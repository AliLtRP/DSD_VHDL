// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
StrMDxMTgUo5N8mDG13qabkRbIX6eIOZP3OWOxmTZbXvyVWKNkOm08ljgj0SqTQHWkUF4IFjycmB
KAZ5aaYHbBLb2JOAl7Jq5xNnPXHSERR41zIfGrV1AeDXgc8O2Ei0TbZXH9FfclVXSLWNjM0G4TB/
VRSx8DI7aXy5rkx8bTch7gAarTAWeNP9vI4k4H8VSKsthQTjciVFnJcjWo2lSN8qvcUOJ/E2EMiI
TTG3I+GsIMOpu6FukZjzzAT1RoYv1KIcRK1dRWCxuA6pa8PGte9lHbNSM2rdqHyaymeqsHpRY2+E
uvIAZR5T/pz4MqI2SORmdlpkwatJFxSkVrc9TQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
1EgJaAM5cLO8z0drIYpjjaCKc3Y3VPmAipJ4m4X+G4eajl8bPxzpRUlrbTP1okQYvnVFGscRLhE+
RGmV2T8uPWFBSGIfxXq0c6d7U9nFcmeXFUtNTWMuEerWrwDQcy5c2yaSSY0V1LP9INx2I0DMlbEo
mdM3m7ntquKlnQc1VyZSbL36weCfWFOSEX1Spqj9eV9oVM+iBdUobMDuy6bcy41OnKgmj9+P8GkR
BMDAirqu+a3GgaYd79vpAPgIxJ43XDNs9B09lTGvBzs1hHwSXtXH7/9lj5Uvd+xKxAMvzTZVj0zj
60GDPvFIhAkyGt0gDsZ8sLUaM+nFzegtZatZOsKBWsgzTvqc6EcOOhnkB4sR0PJNycDi9yvlwQ1d
FPkJxkG4lWmlJBZhvF+4er3UIV+U85fZ1olvoSVs9QkiILEiOrmfTWdfGYQIzDI84XLtJon5fY6U
4uNFrMXiUE0cZdqCEBkPsZyau9UYfCsqZcTkOON23HKFZ+V0L6uZIqUd9UcuX/mnrX6m2H6/JTQg
zIkyFBumy15FzP8M4n6Ur9c3rZn/k/lvZjhjtxv2p6+vVPFV3F3nElaw1rohMc2G9lImAqrFsNky
1L58JZBXmcQBZnI7YwaNOFS6fAdQh3wk78IwsHz72MRa7YBU5JGnOcbOgbARu56FNVtS3Rh8RTMK
5wni34Tx+CsdAmanUVd2QWr9xto4FWNuNYIq3rNYz8dpoqvxZ2zFtXEEEJLSwSx30otm5VChqFPZ
rHiK8kEGfL9pgZ2VO6woK4SpPvoLvlsd7tGL6w0OoaMEj0SykzV0/76SfR76zCMXp1rqX3zgKqan
wTLvJ+nPUWn7yhGQiU++HRajOzlsG6NVwtMwfzMtz4f+krAgmUf/CRWdiyeof1YL+qPMaQxN+OFn
6psvjTDQiekRYUoTyjWyfctE0tBR2eEMIBsWgjKj0DSiuwMeY/VlRsIHZ4CM/ebH/tymApmK1as5
Jz2Z1JCtI+Ka1gUZRC0rR1BhioMuC3IGD3QWih+TTpx1JM5q5GAcm8vqn9ed+14XomArPw3/U2fm
pLJguNOxxoFpWjC1B/ICwe5mxpwXf92hM/P3S1WlnOt99M7xnzUdfjLccA1U1h69aCuQVwMiVlfp
k4NtDbUId3KmcIjl3ElcWz5C3Bd5lTkjUKKClGXxYWIb4I4rnxcqMF9z5gJiwj45F91w/J7dqvWm
jaGgIWU5fddQKZZCJ/B1hR5hGXc6PQoitPgl4ewi+IAQ6R8HKBkSgUQDgbccbjlagrFCj8UXtn+F
v9WxbekS7mrExleiS16L55mov8XWzkMF8HMOep9iE4fPUjivm+/MDjFxkUUrJTuvlm1AQMvOwss+
9HKhuIAV2mIa+MDmR2l6rjGPY+9O0aK9I9hbiq5E0+eIIC9+toC9tnY0PGeMmCywIfpt+2MdgbAx
zr3r+HFAE72QdtwN5FeL4gVO5xFXm4GFRK3GqqMRQ666xipn+V+AZO904GB7TlI6Fk80DjIj1Iug
/pDDLctMPt3PbNTNbwxB24lPT4dAk7ruKxe9lrGiDEyf6RAmf4DWx21rljEKGnD5brlcp5u7cd0Z
KbI3RpxjWWWYlMt5MZpmne4pEMVuMZ/59uiyHX2c3JVRwqL2JQ+dQ2CvCS7lzrYO9oYvse7nEfMU
D8uJt4cBl/v8WlZO4tOmJDiverE9ClXpdCw0EVkaLA3MqyXjBdU9xibJ3OnPYrBA8AHrtH6Cj4IV
/wDfUWMHnTQygsFK2yS4cpr1JVZGwOSNDw1NiBHhYflf1mjZWfyOULbaEQ11t1nue70ktCMkYYye
zjn3ixnSAijFBEtpBMYq5ryQlsKVUNEZky0nSboM0vYcY2y7LSyyFzc3SZBADzvc8sqRo11pB1kA
z7BDdiJk3y4l8u7qEJRB0HZAlVKUWAJQ9MsdTJZ9sw5sAqfjtiRvtsAsl66nAV+6fX3t+7mkHUxL
xs3bfYKF7qGP7nJuV0tuANZ6h/KfK22FGK7DVMj7xflg5ppq3h2LO/VC4rRUOsk3RX6iBuxnH9LV
r+4P2KM7ysZCdyeZMZj8PaTSRwXpKBJb4EGKryCj8VqQe/0+ZcZ8nS2zat/ie2ZMNoIa/jUnsLyp
GUjcUZofGuxVxTq35goFE8UVDicmQZP4YziCh4E8Y0Nb1zZP66n/Cv0Mx9/U/UgUMaWsCNSVPErd
rs1Ulfm4sxy0prI2YhnuEU5j9jlieP4ldV27om70RGvV25/W2sur0yXzrAWC1Poh0/xg+2Gz/TzN
seJHc8ZWUljsL2vn3W5JMHKe4aJ5qDFDJdWDMbafAJHQEz1gcBqsSm74EIWP2Qj1zDXL9Hhn9CBG
0IALraTkvKXKgTJI+9cfqDb4YVhgHJuYnlqis1FajuxxmWA7eZw4dkOF+FwdjzlK9UKp8E6Zh7Vp
R69ZAE+gpeOcZ0Hkc0XVjhJDRH5mhkjVAKaCvlk3EJ6VJjoNhLbWGjlI31Yw6mpw2IgoeTZrDsec
jAj2jQg1CbIID+tmUOZoccYa5HEZYZa/8ma9JCuTdZGup2NIBv+kWCB61pI0kzRgquRqrGQ4WsYG
puoRBUtyo/5urdIzY/cqGPqpd6EgVrz7P2N0cTy+jSJ0NaagRFW1CDX2q7D+a0DgQLS1fJpQl07h
w/ypVQgGat3OIomKp6ygqMKBYxlPdv3ba6Bx4/n4VYW7HSHmZ9dZLNP2OZTiOVj/813Q+ZHM405Q
0VbbQswpCOIDFAI48ULafR5QZ0mhZq4jH+yf5+keAsSHMgZIiK9pLSb5xKQJbqVBekdGDk0T0BG4
r6oT8nXguJXVIm6aQ8G/auS9AqPc8LpfEuYMjwj6Jzj4hLaVZ/PYaNTlyD82FMCEQnM46YP9F4rS
RY7cvhY8u6n0U+dWGWXCo/WG+3c35sLobAXCPCjPUARIi/+Aa9tq+Qv8un0Q2irqaqgyc3LbS8/+
b5wghpEGUrGHVyhJ3XReRZHdh/SR+nuPpoIfrJmr7TnBw1z+5JG0CW76MAOBjdqijeA64UcLtAyh
mO2zFibVJmVaFDTgq/4hK0moGT5JI/YCAFjLpQ3YbZ/kH+KZEfRqDSE7leeuM+ptX+7NqaEDVMJU
JCDr08BgdATDtMPR7OxY5vnKSD45SMtwTiZCvOHNsP3ry1PLqmtnBGFDzEExFKDMtuGPwYMCWNeJ
/dV1OZdr1c8IHczNnkfPKEW92nyTUUTlJubsgBcF/b10N2cFgHByAuGSxJbrWUOrintHZbYhuOp3
Qut+HaZ82uUCTOXmjyOTwJF+ccOb4DyZLOCqGlbsWh+cc+R9xWJpGIAFrDr+1yg5SbQ1fkR2Gm7o
5nyQqQuq+R7DZ6QE1LT6UsG1tfJLIgoUg3MGD6Gx+uqD3Wtuea8V2q9KgHxzMJop5hv14+6j8WvF
u18bd5jLJI1SLf65D5DkwTqV6UxTGywjAlPiS4iB1BSuyWPfWx8iaGVvke33e0G/K+Nfuvg8inqt
AR56VMf9B0P5lInZUEz8Y7idThOC9GP7AGJCTMoKt/JWjVMjA5IP9AUYTtYBuIwdR0MPxYbhfk/c
5qztY3nL9QqhHPzxjAfG1EeAHAiFBWTFy7FKbhPfKqKukgk9vG/cAMAfj5KiRFkYvk26/A3YF8oq
ifDsIk25eqsqKGeYLPpV0PSeooK0ObpA7wrT9Dp/L6sQ8SgoHsk6wgCf1nd/FFRFeenz3DG1+zuP
P6YWoJp0Y54Cf8Pz+7o3x2p+PaCYPyavnXV9ikoh570mO/akX+REzQj+OpNGul7P9Q7AbswQlB5i
CiibHxqmdVDKCjp5uogi7bt1LtmUcvTzdvXHXlVaY4Pw/RMDbZHG5jN895pdeZ8zrdLBJg/DEgMy
41RzyQoqAVGdty07JQFN09hl65zcyfPjmOgko0NML2257P0i4efHZzHtMDIf/55sp71qBo4iiJDz
5nIyDNcZ1cFyVE1A1SSDV8FJsx5qHANbltgIkGi+YtEAj63pzWlwlwDkJvOc8JypNr9ZjzkuboEF
YV6RMTHYGbgmZ7nJecp0K83d7gFgLEfKNGmd7b5GqbZWxAsiRPAk4oZJeih+RZTB9zjNvWXrZmzK
dBW7MQCbJ+NFI8gSWG5sGioU36ra77VhBXa9IYuiZa9mktg4rT5XkcJz+HTqfxLcjRKs8/uRfjCO
WMQEJEYJsxEVxKANCJ6LEuX0LHP0pQbCajyhSA9e6bCsRxbJPXQnpwraLaTMQm0yU23y6XIRWVyB
xgEhByuNZb0wJnfN8Bkx5DXZs2YtIq7RYQdUfGvqIMt7Oxy0bX934qqoRdKwIWu85rjLw1TS77fP
j/c8H42ANWgAopLg/eax47kj8/yfscOJOzCfonkXuBHIg5zxpU4oD/3jEqg80oqN6dPKrgJ8oUbt
NihMRyFdoB9pySbdFLgEMNcz642D3IB/oKN0YRJwoRjwz9QFwdr6grf+k1AejJCMtrW4hVZFnvgK
b9T0JkbCmCWJjtoGW18fGqJVy2TFCIM0CRBr1R3yE3uP4cVq6VyrV5pcTEWmHwITAhrYWmnNH2Ld
awmgtu+9g9lWYkmC0T3u+wtsYVJdkvTCZhJY+CAi4Tg2RuUjp98EwjgbfhZ++vemQp/PUyEuWaEq
gs0AS+lsqW5rEih5fsyGfIukkNMrOThA1Hc2vU7VxyUvir1AAIWsKAisoO7rNRiS9uEZsFo5e3fE
OB77QM1wSaT9MUL0h/iMd69EZLgAZEXudCuaGce06i+SEgaMmC1xV4NVjqhrsz0nP3Y+Pe21bu2t
NVUwIp56UwhlBTAK79wXE9cG7EPY5KhF6Rfs/+AQMGOhOMwq+pc6mJ3oiINcMEuCtFFWl08OMg5q
KWF+Q0c9IoZNqv7yr1ZgQlKEg9JBNQJq9Mh0bHSbLZlB2U2BlO9rpw7qdeHY8gA3Wjnse1TcFHbM
08lgBe4dBHke1BkRmi3iMbKKws2dtkfROjQAvM4E3AP6i5aBbqnCMh5Jk//44ho4mY3SVjIwWsH1
vRgsyRZCmNVBiDEtlQL3zaFpvoDDUkemFdb/M9KvboNsNrUVtWkCpxhY0Fz0BzTShVmKFPzW7Zgp
bvvdbaAbt9uyFYd85RMorECMgG7nAh/Ul6jXPV872dFQnrypiMwKxB20iw3w7GSzlujXyOLYDYF4
/e7xh5erh3q6dnYrxBO+cHvkmuMA8DiLKkSD2P7PmiGek8QOQTWUJP0+kTnlQGoupob4Vbq5H/tW
ew9m22A43wAOqobW6EuNfIjDr5N87eU1QEDYaIyp69txSVbqJyJVMM8Za5v3n/dKV9gjHYwQxYlo
+JF6pdWKy5fVXeLvFcQbYsBTpoNYxXkK+KwdUq/YyKxcILWq551Z/4Hu+k+T/6f8reJWjBK0FKtg
c0vhaPn9WV6DQk2limIK7LiGNFdnfNwfVTQUMVXxd7syW7hSukIFS3zO0oqMiI5rjLrGjpwU4xWj
iV0hRw5U14f+T+lY2WOkYfcFNXRE6eazhgJnX1GllE+NYxzQOEMA7JfJHw5El7NipV9ks6nTY+vv
8BguEaMNej8KFb4oszKhu8VBdwLtG/d6M6s/yud+WDes5etxkzwXw+xtAbIhbCXnM60+YYBHbbO/
LFvKpuSnYY/Zd2UtCw/Vqyy1Bf4PlD8DtZ+HgLfGRiN1eCIOTn6UdRmEzLvLjGU14w0LMeTt7nBS
18n/4sVfAjHSD/y2hlimIfdVgDRRWZ+T/jixRU8hmZZMTUR8zZtpdOcusvPZHDX5kaT9NgB9a4R6
mElw7TDqa51+EkgntPMf3jiF1k/7u9Qg7Q8hc5vBJqBTyU0UUeICOKtP4CnLW9r43MZXEqnZqfnb
9nR1XoLMECgDADy7gHlDAS+76+xtOjYIjsDfKrYlvNhw7NwkIVmvdCz62xKafOSoBLSgWEF6/ibu
e4NbZgNklkaDpNNYJtyBQoG/Tg3K5sCNvU2zrtoF/S/MIsxTfkgRkhrDNPXcGeyhiiKlZajax4SW
k0Pg3l9OlGb8jQN8MiE+/tOR5cTFCDvIpRC8VyabgdZ18b6vBI+f1Y6blDTL5pFib9P1Sv7+u6NQ
jxRXWqYxqepYsC2gpSm7bNaaljwY0Ga1xy32bsht5Yg+QaGyAxuaoxa/9mq+MXOy8Ci/8Y0tpQn1
qUVtvzK+w1w/PSKKbuf+6S2SxIK2ei1VyNWtIISrboVkjo1T43L60N9Au5+c+i2I7iMUy1egyv6l
kR8Ted+Dz0Oz8yO9+ZGEiHtjFDvI6ScspXxSfjQo0E/V4KA4DanMXyxNKxKusxUy7mCQkDFcVFtm
umxaNFgNaWMmijgfchOLSTsrqTaSb16G9Vpa5TGXCUi5AvDbSXEtOzMfStGNfrf87yhVVjSaHUhu
ZEuTdoa5Y4gptEk9xQVIqPWSIe+c9EDy0hMNbV7WbvaD++3HmVQHPkFoUK6SvymVloJZ2dx698SJ
+/mJClN4+A7I/BWOu+LN8MIedAMgpRr6P3BgWTaVN3ONJx9JhGlWAkRulXwj6osHga5FJ/CS6tVT
Q+XS3CqBnDGNmV0G7iWJafRA2GSpvSJ0I9xiwYgHJ6F5rHdJpJBLd4e/00Kd2n6lz53jk3tc6nF0
fWPI5T7Ho04KYo4hDgYzYBMfOCCRqSF6eat0u9dTg7wag3QLabM5TRM/KS2YuwVIROpanDjOA4lt
vFW2qKgnRcB+yk5B5rlRP+M/XS5Ia6PqWLMkJvqx/VoV/1FaU2kQNJUwYlQL1jlHXqY/4gYXykvc
E55qNOyRJKsL69IEAK73kXui8J4hmbA17PaWZKkpmN20JE9YLeK3ARwimeg+/DOTdfymVAJrm5OC
C99kechU46aak9pCZOgWaJagqtpeRfJJ/+6oqXif6Ko6u1bWHLfE0fu1Apnhdu33/1s0g1X3Q14L
oN9/lchf6Mf782fYFszIHC87z245SfF0vaJZHA/1J8ow/Dc6Z1xKfqu9/yDHb2EE5GYRNvCh3jyx
JckuFpbPk43ORzeX6AlexQBiDVtSNxKk/T3zb9E1WvLHH/aG1BxQdo7oGNyoDcT4FqWTPJkkBzZ/
M69JEazBNB6VJujR/uBA5oX2Mdk0KCBVCMNOeJyyRzXfLIKweKQDLVCcT3F3vGsnwkSCuYOlnqdR
vzBoQ2lUZb+SoTxbDEYfgAVbrJfRKYrLkOo4fUeyakX3cVd3QEOf32ryLfvEAhI0wjkE6h22ZeIn
kXj/Dk76HoXUupICyl6vTUCe4Fsai4ERss189rtxCWPx96TBQ78NPg4JEQ3LBcZRgiBJ26ihjaR6
XgnHH8pGZkF2jpGlDc4yPXpRj5AyQ1/UkcNZIAqsppDM3jmILNvEiKSOo7pUrpKdrBPqi5IWnUt4
LlDUOItdg63qJxN4G0pQw+f2odWpXtlAUI3QV2ul694QC+74gvnrmAl9I6dGvQrI8w3lhnooJAho
Z7JqfMJ14QRC/wOMQRZcHTMJpdXGUZpBg5nZyny/MeQceLjm7NgPQG2P+m60eSDyljxQsqyn+7xg
hroPswQqLK/5RpbLzK+gMw/m11Rv7mD5Nr4Gs8GA8js+jJhZyzILQkF+3nMc0E3etzoZCmd0V4e5
Ht1jdhGPnIp5xeu++4XNsRVl0L/DTNNDm39VmaHc4GUjwK1yqqyMWphgGGXDO9GbJEwWkte3GaeB
H6PcBqLY3zpQGA+yxd2zLGiby7Jd1b+M9C7MOTZeLD3qx8bAZlDTn5KE+ETCETBrxKYlcr8ln9Ne
3RXk8cI4Zaa3FFQeLsbkCe4KaMcQzWeC4nQV2X2fymyfKCdWjnATr6P6xM6qzyUm4MUhcsX6+LAm
LEsHZG5YFWKbog86DXp9hclYP2za3d4TP2R4V/ZSgyBBcZrhhaHL4RgH/yB30JCLkgRxURDShxkJ
EE3L6Y4YNIeQgPVo9FyS+Y9PTtkkfl+jV15ds1vd5biDdcy5x0OEq5IX+PXeFXQ5Jc2uGZFL0I1F
qNjrs4QuuSUO+chLc0oF5l145QYDKWyIbYq0lqMyUZIzPg+N/iw8gBLctORznxz0h/8ClmiBs2EY
8Vqp487VVlNHvpBa4gzGkyCHTUKGHQo9NYg5NdOO37+Ub7OjC6OOi01MsAOhn4eggyLUcx6QyL5b
4gUL7PluVeecX4WkW7h9PmI6OLGpfcUif/wphl4EFw0FywehUIPc4mI0kDFEDUEEUpwkC/5TZhC1
NnbUEuFyYZt7IbffPIP/zdCNojaYCkRgRJ0R6s4/AQ6VANSBWaNse9KE3DFL5/v1O1CPFrOE/k3q
CGtC7DFdgsZ6Lk2yvLAHap444pQCO4uUP/UKsL3IwbnlsQtFTTPpqIciPOAysMSUjgKFtK3yXl8U
BzAlVNI5en2cEC0zpHIP0by1C5rzG/sZ8n/o9Yz2umtXaCld2dBraarQ/iwHrYjqmOo+R/+bNjnE
JtK/BlrSofnddbdjytWAKujwNyoO+/8H8wfiZrdpS1R+E73A4K/4Vne2PnBBzY9Jy35iJxsO2uhV
hSGrXqWXDxV8I9pNAkHRPqbNNEcO0HlXuxRcJmFukI7tFFe+7VBL0NLUMaQrtXNVhVb72k2jhVYA
OfowCz4S65Do3nQCwFu1sl6YI99HcATRjJ1wNpJHSoIfhuCd+JyBTqaN5TDN0f3L07sX2r9I5uT8
xMoidaEWEeXPkfMu6hipTnw5KPC8MvVKKevVDJYT+4sfp1Uo1/8FfB5gnifCZRKUon6cD7TMd2am
CYKasATmOyjPoC8PD1XuBo/8kxx3U6liscXajiyeTee/mlSEVOjamvFMopdZWNEnspwZfqSi+bKr
YXskNuU22ptvrAsEVvWEFBIxzTGSpJuELWGrefD8jaD2sHJH6jlPaZ9BueeQbsD4RBYm9m3XYZAv
nZRjatUNpB1Fnqa3VMg3pno6YYzUu82PMeagmygdbf/tuUBrXCV6nTb37lCd/3M/jK8L9eLUibVY
8F27ACuqFVN244s+YAuO3uu3jN+S/3OFJik72QrKXAB0GoFpZUqGe16L0Q3GVCwjgosEtXYpnu9k
1Rrv2hU3c0Cm04BmyD75+eNXl0m59b0JoM4+DWxUanmphaZaD8O751J2jfEOod5JCIHb4oG7T0wx
oxSjUGzlxOVQ0dkORzyErojapoT3/johpjnNLz1esDBwbXCeYHZSEoOPJYXLD2O5CvNx4qTmMHBy
rfdpPimc9pxqCPmGArdkcC4Ux5tDldjKrhwMkoDo2UDuKLXf+LqxPOcX0/AAz7GyTqqPsC/GIWOZ
h7cA0hsjFHeEkEOPSNq7+BiQE2fSGEuIGQN8+2UKwlek3wVIjIdmkXEb1Vt7Py8QjHJCEKGR7Vpd
kYO5x6adMQpG5MlwJu9vRJF58wuWmcc7pepik0R3u+IBptOzpMn15H86ndo/RQsDSOj4v4oFbMOS
aXjxsZ07DUWPYHM6Gkb1djyZP9aqEvwA25pi0yoR78v7t60FJMeQhruYRuTaOaodT1gxBKUCZKYc
yNDn5Nf38ObLMYtJFqU/PxokvMux1crJ5CLtmp76WbD6nQShCdDdO5wWFF/jxx9xdpq1TohLQ7Jx
y9tBa3VDX9u0XgfKz2QvRSmMvekMJ1zs/i3fUZq4iFZHaLLhoEVgtXZD8KwEMKIJeGLHqFSczooe
FZ4Db2ZLq3/KbSIBP24aXA7hNikuKK086bSB3k4NV7HgHR9L+sr7FVa1hTCQqtr4PX3rg4e2SOix
L6BrNAv6JOgIaY/lIJn2m+YpS3iQOswmPfhm6VSop0UmJ1nuEQ+D0XUmgI32xBAYuObRHoiEFQYV
fU1Z56EmjBurkzIw53wkhi7zikATHZDgXuXT9/alSwBWQD0xVBP8LGjo01e5wJd6h/6/Kesyc+p3
goVqLsNtsZhRyJt6j5MQVtKnTkHY6zV8jyGJ0A8wN1Ver79qFX7FRyAATwwLG2HTTlBmChpvk+Vx
WuzbxopLrBzEqidRqLW9U+VvHMqTkgozGv/HwLFq61HXAYzrLX0s5aX0yB9WC2uiie86ja3Sk91u
iKwOrr+kggBGcxKiBgfxSQJcvLwV5Y9LYlsqOzMLx/x2o8WqM/DoZI7lxXE3hV7W4Lpx8NLRTJbg
GzyEXVP1lHjmDSno+QmvtV9QXaP2NdO+FnlOdN2FH5yq+RryIbtVLq2SV76XwpmaU2wk2ABCFMdm
fVaXMLFtwdE7uy7yvaoPAhwtDlgLXwJboL5NZIvsRMXjRw8fKfzn+x+Vs5hy5tnZHGv/XRJaLqy1
J5XWdGC5OdJzo27h6r5cjUQkd5Yh3s7CY/xREneOq0ONPRs+FkIzPvDzDwncMjzGYXLOL2N6MdDs
pHy+Lm48MbLpCcoZdEX7c8htKQiF5DJzjhUGJo+jhUjcyIt2ArBSICcnWlWc7NsCW0kTOYgMq6l3
tfuKgz6PoliHFJLgQCTnV247Cb/3iR8y460F2qLcViUpO54GfesDrWsKT8TvMrrUQoQDGw+w8wsX
POgDCnU6eaEOc3tTZt9RIhyGeBRtskJa1H2OVhhs5G6fgdCICAPtFJwt5P5I0OvIoEH/ijxZ2Swa
9pu5Av6MIt+iYiEsnYjc0xGlO81TqPYXZDHyxEHp3UB8FMvJCDKWkZNlqwAD+lpV6IqhAu6XsjpE
CAVh2dJ0neKU4GiqE3Ai53zoBwvcUYfTopBuMag9UieKALu3EXPYkttctOxmi/ezvzBMD7mOHFMY
iwYMuIwVNXluy7kZKFs9Jg7f/bSE6Fe/kf6P2gXKAUO09ZKuxmyF1KBlrp4aZ23BKwxFuuV2wV0B
dVXD1DP0Fx0kagqTN/nQZI6APK9wzMH2vuLZ3ccYj/Ix61arwIfSWlbO6EUdsQuaSQZMEKdRzpFo
HSyxyrEN2RBveN6YaTvhF0243W6kLwaW64vi6dQHeF626YpZRq6Ze52lV96MMgsX5msc9hZgzLGm
rxfFf6T6v55oVBdaoTMffBxokMpz57vHgslo6kimJUOPi4jeZ5Tjm4RBeUxZoQc9DjPSLu/PVfwF
7P4XBewCC3IoiQA2k9sTnL4AAUdTfEMzmJQf5THiPsgb6gxElTwtKpi1rMu70mLunVnSNmHdAprn
ahNjkxOahoiC8iRTH11f1fj3sRG69++MumNut/Gr2dxC/9kwvsyOv5GQbhrrXnBRtYkEZG18CCdL
u7vIhfP7x1j9hCdLNIysSG0ITbEa5C0GH7roIlySopdNnho0FzNHWwUcqUleEfQ2c+63drlA1L0x
yKw6Eeyuj1MRDEh6I9gOlw+Mvnvd4uEcG6NS3HSzncoproQoxBU6delf0810dU6YPWqc6JyAkkDW
IOZGWy+09z2B9vkf9O6cP5K9WtxPhiFTg2sX4DVN93XETQzWocjALVny+JvN6bjUbz0Lc4RGXP+A
r+0eP9b/RbpBUVWMoBhhu7gUZIMWyiLI7MT3j0alingF60rEu5nA4HmAxhknfM8zhG2n3qJ/BxRj
mqSioYTYBkueQ7TRnB5xsXa+8Y+JwDwWIie0hZwZBzZTAjv8JacORsoIAOrcWwe2BS38C2k25FTD
ZP99I8WMIXvN2dnMMalyTkZjoRk//y+zDtueQ+QVtinQ1ha+B4uhTp5tJjYjkORJ18pwjjp0BDbb
76OsRlt6TrhEz1/Go6LRYSjOHQKtlfoR/MN0Ho+MvucYdai6ZgtmVVIX+liWzUPaiScLoeITlI+A
3eXy5VMPWYtn6QczwDQBKP7n6gSPmPux0va3MkkaE4fD7anngSv5zSqo9pPf98Uf3yUZEnD9DyXo
xd4pADZbG5YAaIE9SPyJPr2ZIle6L7xbBkw0gN9yCG8JAo8eiUyIT87l6ClCLeXk+IJph4JvBjs2
B8tK4JlBbas66rBXcfMtVNmnIl3bz9/wzq1ieggiaVMR6pFK1t9Wc/Sq9kTf7PefO3lprAowMvXA
wvab+lSfcPOfpQl8Md1SQjZW0sEfIR+UrcnTcB3QVy5Dg/rUuqVxzkay/sRjj6f//t4qwhbglX0n
swjrktwPmKB/pzZjwo9B8vMWM3cXpF4vVDcF1gvWi/MKmxura/JtpDRfwDx8uyxA6uPlGA9/vMSW
e7UFP47qKxjICSYN6X0CUKcZX+V9KcvIHOhXbVHPJ2GeRmAQrcw9xXMn553IgHA3jE5lkR0pLYmJ
sVGD+1gTtTQkh9YG77qcIhwCasl/1fmCxwYjGCfHSlKCiBfScxI4spWWbDrehvjRZg38f9ofre4K
z3lGficx4U68AdXhG2V7zaEkG8m0LbYjrS/K3+AeTIErPHk2M06xVZuw7BaEzW0oDe4M+uaJBxNA
Ws2eH6vpwTatOemxGwy/Uog79Nm5lkjG4yBIV8Gm8nfoTrCqYCrv+M55Bh3oygwO1oLxTg8xVtq+
WtAf5Zx9b7ooNF/C7GfZrXOChHhr4mr5S5hlJ4Huuiyc+jLdN9wzrVo6qwA5TaVwWFqnwzrBpln/
FG7R9U1PINtUKnxD+O0nfk5Af+IsrntZinqDgfWPx2WZYSywiuuc3DHZvXLeUllqJ4eTi/PdsQIM
lgT3ggnb1d1TcrwzXg5zIHJxgDGY5eaoSWGvshC+Irpzl0aT2AhSMii1fgJqwb5NWYHJhdt0Nqjd
zwIMhI7Aj+QZE+qQOPR4f7/yrdNoIykNYBWS3FCeoz976g79iEjacW8JoSoJomODZT3DEsWxBxCy
VUJnTiEQG36IcGHbSGfG6sj9IrZs2qZOoWqc9YubXsXaSdxCk1GhOSOx05Eg7b4rXpNBmLMbMdM4
RK6xqxUFqV2YRep7ktc26TgXyl3811KmuWxBbkKK/puru0lS3QKZ5MpaZxi/XxjJxLpI99+T5Vaw
mhpvL2bqP7FUwHgNmul3B9bsD93iNzNpFO9ym+a/KUcZTaGF0SfEdFlmglmbI1E+PZrqG7mJkvQS
JcnB6djJsIJiN5IDYIARbklh2sejXlU5+W4iHbAIZRdImBS8qoQcrrdRVRCwrmpseEyHGLaK0LvL
jiwyyA+L0EXvEX9syQdz0mC3LJRw75QD6mlTXez5KhCTwwTEi7P2STx0u6L//Am3RNv2krLH3v+W
WnFC6BYJCyLYosaxH8mLWAU2QKLy/E38dnemv2pqjFmxiB8KVmT/RTay8d3tYbt1cYn7jTGgjTy+
zXReNPBZGFdaQfSOwevFeTGBoY23271NumhDK+LRTxtPl8LbFDTmXc2v2t6gjvt2joq4ld8T5yfZ
7jSndriC+6ZUCWKKfhrxnlwH++J9GRX7vYfhLbXzl9dlYtHGvRD/waXJrr97eranSZPzOsLURWbU
MhttqZSgiKjKDQRC6PHAZcX8XkBc3UMxvml/Wn4mpbeSvGGdHmQi72VnhgAYb7nugHQvfj7/7Rxd
Y+/9jw8E7FBsjBoYlWtTfd7a0d9IxDRag9wBVG7TCYdyXZn8csSUX9KGxJTBefjTrOrLytcn0Gk2
i5heOX7h+Gjzko1RcwsQ2MJOUXyMAYUHrBzzmxEgYxsp6Wkq+FrsUbu5Aq2x9NoPC8gS9PjbuqU+
s7Agqk+wJCS7lxh+Eo/NiXeY9nGUQNcs4XJCGpJw/lril7KSAc67FfV36VhfRYcETlzBhANCXdkh
IR9dkC9keGk8hWvT2p7jrJbSwihJQY7nUrYVNN8VRBfQVvGDQLwpitqQe4sB1RhLEglLvYgbNr27
fMBGQuoHKVKz1ghz7QKiiJZBO/MoEDwfybG8lG1yWQmk0niNOtN4QDbRQnjDxGaddTlDqbGwYg6u
r+4D90AT88EJcScmfOgQ6zwTKbxSz3XN1opNHghRCz70MAzqhuEVL4OT3q2ECSyHRfCu24UrrzPg
ac+dj7Igie138kaKCArMmW3Y+QCPjDO/WzvgGoZgp7E1Ea1shq6fdMnTS/286xFt1hdS2EM4SBw1
gBzrEG3sEq7+zPj8MeVTUWi6L1zD15vZPqRVts1dIlgPvuaV/7X44GvezXq6W+yO9wV+XGf+AZdE
jJBNmi8XIBU3Us/aWPBG3fZJu2JEb8KJjkC0daNH+4u2hYvvQ8Kw6QgfWu6NXh1XtqF7c/Y37qEO
PYBL0NbRahRLfOdnyblV16312IGzikx9RPfErxJI4MGwxC3HBvT3m9IlEL/aGuxJuC+jDqLb0BfH
xy8CW+xmMjV3cdYiBC69/QOT55+yQkkJGyF4qqRibu6rqXF8IHzQUu0dAH4xsHXrSM/iQi2MLc6L
LjfJB9htSZKiRqDfN3xGtOpcGd1glXFpWD6ItjFH13lj/ucsd02TuUhdT6JPqLxkdlc9yxztN3B9
c1DuKTUZFy77cpbaI8qLienbW0uhfBqQ87cQq1AgDN+0TLO5fcGM6EuDJ4kIptw9rYNarRplCcDO
3n2fUlZjGbnd8q514dQlZbb7y/KmrCPZB3t2skDTGxRdwv75ehTVquqglPugnu7GiHYwV31SdLA2
Cgz6GsW1arK9Yxkb/WNJdo4FfhBj7kT771im2SQo1M8554as3SMXURg/qOltKn9tQClZ3L06hO+G
FsgMHzEe0DanimxEeP1X+YT5dWaFhxxKiJlj+8OMVOGhVz5H5K3MpTTBzkVlqtY7ZA6OEsOlu6Z4
eUYxub0pkGftFnvmgQmDA/a28YPcFiBA9zIImtKnhUs3x4srfirEHjeucGvPcACPAAuHFke5/5Fr
yoXJyna4bfrIwRZwHkk7r+JW+W1ILzAIqKJ0GQCF85vufeIbwTBWDZOujaFrOmfrHKrexlqHehCs
h5hCfll9SyHjjHFJYlDiuvSJsRByj+/dPJPTd3VVJkQJy0sviq0xzpkUxhR4u8hmu1RAUB1DjdxX
7HF5aQaoPqkccXkFSNxGFNJDrVqb0MRCxAQTE3qe+juBM5jBMEbGDwpOLRyoTh+Pp/6q5eUxSYUe
ZFIM/APw40Wlohop1Z8O9gbcCurDhF31ity6PCB1yY28LBrpImPq7actVHv0FdGiaKSzz16icqGX
wqimUornYLBRUBHsnqXn8/e5OFCHEQUL3dQf2aJI14OlJ00NwbXwt2hBPDU5ndsIvl7RZhjHl8Md
G7JNz04Bi1r45k3IhvMeLxdI2lMzDmWP6xzZd3VNUH9B5pSaaGvEvqVV86m8apuZIhOola8FEn9a
xi1WoG0DO+eqPxB2Ev99dn30MVDIEkJGSW9u7JmsxyckA83+1vAvyqlDQwG8u4Qf6njzjC0GFUGH
/LUDZq//m4LVx3Tyi852iOyyuj9gFsC4vg5fKjorRqykdV3ahyRnc8z6yJPmr+/vW+YW8do1VQrU
FIdq5ntsJgQYiWnCX6YUmyKb0kwjCDhmDteW8dlfY3h9+mP+trzjo2un7eRfhqy9HQdg7lCtRAXy
Y6KbvRp0ZIrbH2ODl5RM7lzxi7w9xvyVdG4ZEAYqq7A+NQ2ZZAAiqjqRNgNYRlhQS1D6OSPZCEHF
yAuym5gIJt13+idw/A8Q5kuDBmJMK92dJq8llgWEuN2pivB8q8OyAcdteDUUHX9+REvM/k820eET
52N1Lh4vB0TpuuMF/At3QVT4/nHNrPjczHG60dFttkFtg5NkLcY+YNK9goY7pB/PSr7+r1SZJuce
FQN5Bx+Z+LSFjp5lHnuFCXVfsPUk/czgqZyzLrmSEkGGwc+QJm1P7JalZh/idiq4rAQkX3bwScr0
rX8XbAcHC+0PywMupx6oNMIxDmS7YVi0sCh7sC4Z+PessGgGsuCmkSUB3ON5lVsz/8CtM235ccNX
LX+aaTBHWxQvSJ45PULbHYf09ygbEGjys6ry1x4ogrxhLR09zIYaoi6BXZ+2k8lSQdXOx2Tr790x
GOTVNYE85QMhYux2LMHkroXY9iaTTHJYqN1rCE9ep5eMMRuGiq1M9hh7BNwLEYy2FWo2rxR9juI8
iMZWs28NSIe+VvR5ydxYZWXt6lYimqtLdIGRtjDLyvIVv3RR0bjWpq55PLJN5covQ7ryJ2wWaD5N
btGW+N2iqQqmgTQz/llzN8X8SnKxysLPgU85yqbwhUX6eN5mrMyIHplpxY39KCAEG4ADnCzBBPhV
bYotOHE042mIQ4Rwgfjk2lviWtQ5FR+vzTnpe0dnYj1Do/7U3z1PgXIaDjFJn0JQmA636XSpTTSw
xTbbxL4Ro1uNmeA1xFKdaF9HH/0EbnK5QyMnwF0LaxkMT4kUnZ/0Kj/O6jJ+Uw9c9GYNAsA9U0dB
XC5RcSId27udwGTD644HVz/11VbTFUY6IqRFejZ8s7hwBwLfEdWgXPBa2576DEREv8kZMgxVAcfL
SVg3ppbzoPhAKGfRmq7U6Bz1naMO49JopSdz68jtEylwtGd7Igx0B/Oo/eu48c4Cq1wnaoOwNCJq
5JdBrv3v5fQytg7x8b3viSdAFFXa14/ujma3FltYdJBh9u5obtMajf+MFks7n36ttQpoqwKDs2ux
ZMOTekbUJ5oXPfr3HPxpIxlCzfn9DirPq4XmyBa6d7WDHLwT9bp1xikJobZMh2ZJD6PsbwL+0W8r
1TPyoZdSEiFa+BUeR+Oyk82KsXkAYZM2hrhYypOPdIUwjhNVw9NeyQbtvQvL+wVZ4OHY6Px7BA6m
n7l1fZCisRHz13Cg2AGED8txJcL3cj7Qy0niZ5+QQV5ee9u6XjKC9qZ0RGUTkGzNUPfjp2d5DlJo
ElA1GUKY/HlhGDpw1elBpePBwbI0pnq4aHGvkRiM8DD72Ll83jaVhrqnHMI6auq95QL7DGUsHRLZ
iCz62AL2UVxDT8/0ofU9aXADnBjeydEGVaj7ws08OxjFP4zOJ6zJBGbk7eEV4poNryJ64gObicBP
QWj00L0gYGEfKoHCkqyITsX0JYQLA1tnElAPOoJpEqdb2ifgFGATK6t3eTGhJuoPMBodVJlqrONM
UG9vM09popOxvs8Pr4jP+2MtWJaJ5hkMUfHCtVD6KNITogaaiNcFp45QgOntZy5Y52eVtStea/i5
ihHSyUG7Rf0ySd68PVhP4yEXZKCv/zQyYrGz7M5r7f5ZgQ5j7CBKxqpOj/NyCetykghIZdErkEtw
dxDb/bcwXLi/EAKSQku+CVMBmLOMx7AU/Jso4flhJZu0Jfy0C97JIepDpZuSgGPomC5on0tQk0vc
lgQvKvFlUyRpuOhWYMFbS+nTuL1btlAjsajn8fUVehhZPAhwwwMKkMwjCEpEcjHLhBU8zMBkYoWU
yFvIzPGy5nG1MRGVxe9k6AmAs1G6Nmo+ip3K0vxo8wz+pFXf6nEumroEw+Us9p5uJbtxDCUNpJqg
3NHlGDcjmdrsf2a3OfxopgSqYl2uTNeVAZymi1n9g5Tw0de4EmGXl2xyjLmJn44IwBbE7O5aIPbT
61tIwo004C0LWF4sVN9Q0baJ6TSLLLexPelHSjTkm0RNq7l1Yg0scaRVMPNsA7zBN9nMqKG1Nfvc
5t/K0yENSTGxjVmDlMENmGsroPvpOoMiKmgF6/AlyacaqePPv3BAKsKcarAAyNk7ZIOybcETl2PK
O8PrXIDjMnjSVCD0btz1zBU3knV0WzjUjfqiD0TdwZIcLc21Q5K30OR6XFjHR04zp1z23ZeyTnM7
zXOQnSn3hBqLZUw7G9KpmDkwN28k7KPfQ0Q/2pr8U19kyaEDUJk/HjSCMraXCtapTAoyErO+TrYn
yW2SgUEEgauy80Wk9QFuFzGXp+STdHtGU4NrV5bGvxI6BeoYlDglFq9FJ5gW29rDOd9nK3xDkdQw
gCXIXXaMYEFdSh6qcML5yat3h6ZmogQuJUQM6K02jJ4m20Q5TisV90iad28+AxC/OL1zB4CoSkH4
P+3GKSOmcMDiFIqZKo0H5U0h51TaOlYe/5caKeV12bW8GckgSgG4iTzcu7VFoLMQ1zOxL1rO41+S
6Qu3RsNl3kEf5YhFvLiTNyVer3CnRPEXyhaVS47grt8NVist6EkkCflwEkpNoMusZYQzf1OSqzGa
5vlhrQ3AcWODfHyyyptNN0bHSa8f76ZCl1xsStZU4TR0OG5x/F9UjeSNSnorXn2G5ds5lyEWyltY
vV1rqVG6yLzyR5yy5PsWijIngife32Ee42Qoirj800o0jmT8InQfHfUAsS2WUEIcTv65sy0qLa5d
f08cLDruymnFYgf9J8MVz26VeJk2UulJAJY2CRsGlHpQJtqfHvo3We/0eG1yRyP+s9zMaRi0iZkk
S6YACBv13pXIrkfXN8PUAACNuHZHlkbD8XAHb9S0S3sgm/mvBz4eYmdqlfCarF+mXgZCZsLemNgD
baLv9HMMst1pGCr3vVsQuEspMeIXYP6W0nCyuH7oGg29wNQ96NMl0eXF0c8Zs9yIfsyK7IJ6TLm2
HW+qodRg+Jc2FUIIuUZwXMsK1W//1aYwAnR0eIuqJl9sGVaANPjthREkRGJ6Jf1MzNdcV/UvhTO+
ikRQQyr3joO2HsbGZUnjD8tFL0ICIbhRyDLjFkxyeWed8XlntCAX3mRDNfv1nIbOsLCU0UGMzH+3
ebM9m2+Rue6zWNQFvqoj1pn8XcAr45Gm69nD9VEI4YnNO6MImfj33h/dhOtaW/1SAYK8C/aklbsV
mypp87lZTx8WJjrBPJ/WeTiGJQ2hN+1dQS0yfK4c++JM+RdmS2YBcdgr3RyiWeGlMDFfQwv6jIKY
fYim+HP0Fh07xeIfVPa0hsdDSB03Hq0+42BwjAEfLoHWSBpPqZa0AV4CR612MgVtyHef7QcMFO/B
C949KJ7uuEWsSEubCoiPvezduIikHCjp4g3nPLbeEL/CJEFIdP9SrGKmp4huzws2jNZVfXqvyW9l
Y9+BDdLtmEWH5G1h/vHgyNhi0sBPJTL9gMN5i+MOJH3HBHSwBvIGinAy+JJiBWBwhlurvLokz3MA
U6fuJml/e/uXFVnOZvO/UyJQytElIfNrW28ADD+bhI0duvrEnmSWD30cPE+SXW5Clnrg546d5yQL
R4179B/CrBV9jv1OoWQSTT/i7CC9ipS26a7nuNXUVO1W/xcDEHYObrKuNxC1OaqNoFbWdodlcs2n
AMZj8ZDErZ9Ei1TZRnTjVk1ESo1Q0W5/kF1n0PVOQx+wkWssMheXSxUfBOYfYxfXInA6Ml8pSXy8
vi7LG9u2zJWut0hYIesn05qzQE6mguEhpCvCMs1d5lSEgvcbZRkLq/EsCzV6qPFVKTjjHWsmYCGm
ICWaLoFlKvEnf/68/VxdZMHq8mcD52jZhjwo4hIYTxsQW32YOL9Fxry1GllE/7vSvbJtT3ppRPY3
CiOYCSwx01U4TjyrfYEnesJhCoZXFZMEjs/vqR71kxIt1VyeYC7kp+Zy4W0CoGNzgBJckXZY1m7s
oU9toWWOAtBQHVwvZ1HT9grmr/iRIvHANM95Nme+p8FtYSKZAQYnnSLrWw2V0O7/xwmGR7nSVnPA
yFYqltf+yiS5gcUgw0/TyyR4pmQBEdraUM4HAZ1khAp+jDCv9toGt0JxQ1Z1KuQsGUTaaW5e7Nhq
CxYVnZgpQFlxZa/5daeuhSwzEqQtDFHnNwl23b8X7oFGHyqkZscuNRFRK5G5ffn+sBjibRcor5p9
RsZR/egWEUE4EoLGCLja13NMP6h5hvmMj2k7s0lzhvruj+j5T5zYzvWPWbaMWbZQZXAxMM4MT0ad
1Zcoa1EpiU3kbHfTqBKNDsbcLyafpdmH1v+nKjnxEH7OCeoZ9YiWn09GCBpNXYhQfc4tnC2y/VmD
CbYxmrwmlBi7XWHH/YBjjIkCgRiHqvcuNWsAwtgGg+hjfyNJMIKz++NQ97eZYIle/ckSwMvm2Gbf
7XByFYRRazCrwbI2AuBUGZ95plUbCmmjtRYOO8YR60MbJdY3gHUB87F9VviKcxNj8zP9L9xfLyUi
rGjZcWGmTzudS9r2TtnA36xaoTMz0wADbzZ/4V+W5odEAqoVH5tb2TSzQzdMignajQN671+Ya8iZ
BoyW/YJNrNHd7I5s0pm0koQd9WAGYCyBYUJMrd7vdCW6VcFmSLHllpF+qUIfl8aAu14pD5OHyv3i
a9s2J2jujR3l3DhJx5SgHlTkka9tWBN1LAzxXghOGdQkneqAOaEumuHePRQz6r+omEZL0eY59ACC
5K/p6C7S8O5yiwAPNE8NbvpIPAhZb0nv5af2Q0lddqCX8bFuV1PKTgcyqen5jwB6fyMW7+hzHOVQ
rYJnRnnR3Dpaq23hyF5tJk5JB9IPYda72omt8q7rFf9xgClosMza5nDIbXIaZnRpI+/PTzOJpCE7
vy6I0VahPV2rWHipaNuyDlZR3qV+DjcZDDdgz57BwKroI3aUIK4CLFRDaaRu9YI1+zEDdJMSz3WM
9ABhiAWIjAR8cFUzuf8sujmRhA94u+GvEbvdRVqIWTBCSDEymDRbmdxjOynggYhQxZQ97LfMHY+V
5vrPiOSTa6SSdSWEKW2L2lPhO8DZ/Yu6oD+dadONAcn0p5mgw5/lKe8bR83Zk8DTE0gm0UvqYAN4
aPmz9pdF95NNaEKdeSxWoHrdS2uUOWJBRNy9AhT24SL/FMfCFDDravO0W2w0AD1KHws2yGV1px3H
igzr8GXM0+JRva5PeO4h95ehqi32ZOFI9aCpZm3DjW7282VFh+QGUeGO6d4qA5O9TBtZUAZQtex5
7JqoPt5eRW1pSh+NynvrVkJZTX3lCVa/vDnYnt/dwRVtzxZayJhZSUn0j/rmcT+mR3YBnYBMSC1u
yel5itmdaohzIcB/1gxkzw8q6vzwua8eIMKwg5xv579NEEV5OszrZFtUBd8VxRT96jSvoUMDpngo
FMNMJ/ochUzyENaVDKVjCvqWztIUkcJI69kByQs+pb5Ecv7Y0MrT/Os630gtYm3e0fZq/qUfPeuZ
ezGgu0ipbXSySSPh951YsJr+KNyWMlTUl7DCycZch4Be9EStM+DStpY/xKJYeFKcAtXwckT02mWD
1gOTc0a5tNDqcBoMykwRm05dqS4Gdc70aj2oFiaaAV93A7raDflbN0UulXf8ziM2FK+7761xjZQZ
JYXKnVNsLAVgLLDS06+49u8ocnTs9KyPu07iOBDAs2MBSD7f36FOPWzn8ahS/oNOkZqlvdoCPOAU
eWK/hiolOVBdbSpLCeRxbowfZ9vLQiniVNFF+v1Mf1JsSFsXQPKbYNupe/jw6m0EjJYSsgHxx6be
c0JpAoa4nImqVlUhkMcy9v1ynai0AI860IicgoIsrpWQO/e3Dv/GmLSMACTmasgMcvCtaUiDnvpF
BebgK0CtmS0b+3XFOd2onWUeIyy/HbHwRwCsRWfswLVRxzW6kK2FG60Kh1CcF2Wl9fJgosZPZ8f7
R1e8vnEouiUKyK0RJ8fS1DvPNW3Ka21AHDCFp3u7/PqHvBnOs48SR/rJ1LDM23l+zNDxCr595fsV
FFbTLts437UpxSHvzk4pg0Qgcl0TN+SI0OqDE8h9VcJrHbAjmX1xEDq8GScMDXcxsogl7Sg8xMbB
ONauo0B5rJkHZ9kxI98pSdpwZqrWKspjD6qg0fZPKP3DJb4xSemwWj+cs9tuMOIa8dKUBRiiFuX5
8OB5Fs17ZGxtWKR4rMFa2JCvE/EvQifuBopFDVfZeDTxl97zvQFXj8ethUofkDFt1k6It6PIq+Ot
F8bZXCEgHi0kCFK5Ih9RJdON859OcGokdxO8VRF9385KTiTXtgGs5LgttzV7uE6Kqn+k4XOKSfbW
fm7rGghTl8PphmIy4mqst0/L4g/OZCI/y+RQ2BlQCk27eNRKvDsHJorozX9Lnno5cguD1/1hmhRA
kQmbZPsUWLsK8lrQpXuMI4JcrCjnyhloJTzIXEdqmcx0weHbsEQnpLBhmYsr3apPY+zmBKCTISQL
g6AZYKYsnWNNvle+u/TRizRAwXfvWSbccXiINa21RHadk5pDGjyZNeWVPBXUNJoHprfmBf0lWz2A
aYmIkxrS2/vULPf7qjA2ztLWbq8fn+et9lU2iVlri607GHN7RU1fsmlFJeONzhE0a9qGH08uWTlr
COabYvFBGriE2uV/JI2XYO+9JQxm4L2r3GyGcmktW8PebDTIUjwuF8rHaXDGxyRkqdAXBn1yIkgL
VVkskm9lhtVkxwNPOD71V0367qpSXclIoQo5cQv3FeZcHRWfVz92UVuatyy7OxYI/mb/w/LebSIz
Luab6+RS9/fq7LIY7694oMo52sIcSaXbML4HsXTSnvZKcJk5pjhChq/sOS6pS83wqQNvbxy4n/ih
EyYF16tVcxR3uwM/s4QrSyBLs7mg/DlqKX1aHVVG9QtJxoWC59iPmOPAggjwLLKgQW7ezZUnQQCr
j0+AhvHyg9+ubwaMJViExTaiIl2Amox2Y8eZ0jYWam9OvCIur7Ak5vmCzm469s3qgAsjTclefw2w
7MCMcsYRrlfqCeBhDTFD36kPBGOtRmiMzhnhMTmWzyAVnWW1krbFeDw1A75mEA5so9lSY58lXlnK
ON54bzDfH14z4KfTkcW5EdIrAWRaFEd9zhilDAwD+W26GyiHhpNq/gmDphMdOHI7ZjjtWeS2v378
Nn+CA3r6y4BQqbomSde5SmwViK4TYv0ZEUaMW4ToOgsKQSfwEnn228JWoGqwgYISBQkbD14Jz7tW
lx0D9SOOQNccqMgwT4Dv6ZN5Y8PlW/rP3Vzp4S1agU1C4vHkWNvPafg2nNUgLP1bUCHXtmU2eg4a
OUlHYiMIB7N//PyfJk1+R9vueUcghbKr7ALDGD/kj4Nfd/6iGGAoqpPoNFNzp7woYmNW7oRPU8Tc
q/BM3XbEIKdTbjYRITs3yPPDNe/rOdg0eVAz8E3MNGUeojLWpzxHB5vKS8/VYYDJd8DWP+Dwx7YC
RaPCT/HQg6gvecHJ+rRT9XTF9m/UMfZncYo/5z6Tk1bNSBjI12Um4YWVwybYVgSZP8wFoCm18BLB
6kzX1qkIW/yuSiEhWsn2SfXx6wfDYXEjjnpKr+tEI/xE9Ij6gOnfq5L4SF7eqU9r0WzzkJcR7f6F
6n7z+eWUlkAOvGgvozFHpXAs+jZ659GPziZxHikIE2uerw8AKJYqAYUyrJtwN8PIoZ4m5wjMzSoW
bocMdu2DBpTO6QJdYC16KOn1MA0fiWc7o+LUyUjgwJBRM3f5u3PeDbnH/NCqJFX6MRVsbsE+7r1z
qqRyYgEpDRlLieTPiud7Eq1XKGDomg5jVBitDGPQbI42BvwMuGjDB8Qk7B03m29SbYvXrNAa3XVI
kFDF0unArBvaUR6JwPIKKWR0AW3PbkYGcBIvzQz4Z1nti+HRmtNW3Ge9wjFJEHfwIIuZSEflg63T
IK9aBQVh4nd3nFWvggbEVMo3j7gMZqZ5YUEHFlVhOYVNlWRa51XZZ/WbXlTna5Im/qGtBp68ZdjP
pw746fkXcOIo9z8PymuHrpz48HyIrFB+vkwo0kSGRnAhZgea64BQviOh1hn/8Welqy3Cg8zgOypa
iVsK9Tz/ojxvE3ae2z/FsUsTg7YMbd/lNuvX9WtORlrEPXCJ5xEha778Om8QrABzS/CpJGwCPnDi
nn08Ak8W/HgGhnHyVnTrtavefTIxrGEY4hNA7QGszcQIBHOdySC2PI0a66Z2qP62lKss5xWW2Fn7
z7sI7sg+yVuriiJVKMqT4P+fLuoqE2WB/z6ogN6XoIe4Dpmp4KP4aHlGipSEK99cV/kXY9lLclOd
UT2YRlVmpB+RkEZ1hhsFLajtuqPUqUtpuPAy1Yzg3DVbIPsUY8EawKOspXo8GZZ0ys8cVSBVI40X
x+tA2SoKZHD+0Mmh8t8LXNzVG4sT57Jkb+YW3mZt5k17E3ynCvPuMoFHrd+UkbGxkQYdsHzWx36J
JbDYEnMAmLZhavDgQma+s8il4g3WUmhtnH5p9NRuSu1mQiChEsILboW2YWcY/6iBUe07udv8PCEe
hAXK3TMnEtJ7qLTV8GdvTzZ2ZB1MUUpymwVhygW32MoikZtbYBijqEgMvMAP1XOnPSS6lcGAmnJV
6vxrrldDZxJUAUK+5q+spieXI1w8b7AWybDjjqhxZ/Trb3KYnfCaKHlHoXbZP1fZ0qlWKYEAoSQe
Wejfb1ysokl8CJwuLSj5UaWlHQp9ks+P48Qrrj4/NHDTKqPVGP4+RgNnKEWoauSZFWi9NjN3x2b/
4gItaXLWEmd6BQsRFUKJNse89VGpJnUUp1l7yDtBLN0uiwPpFRO3Q1EQbynSeLEP5EIRrQWYUhAc
CU5fdec4G6+uhgbi7GAasbradmc6oNwGVqA7DRi2XGMPJT3UD2k/ghB2BzK6CYyTplmFp9HF9bXZ
4aaUvNnEM+xa2AMZboao5GZATduKLeK5YLqzEoJhiiLMLyiUYOAL6NS8OhjLUrstmWmIf/IGXGUS
u2wv1tH/17e9YSF7UhGYe7gUPExxX2mBPG7KjRaB6mY915WcQQOzz9z0ZBtpbY+TfaCEWMqRZFUE
Iw9TCWOoOwMp9rszfiRWWI9qOMjOXT0qF+8jlyqSVKJG6kIcqxYAffZz0MXFYl87TDmdF4xb9kVQ
H5v77fORM+POEYk4IrAWz9vt+JqVavFzirVa9Me0d7LhBbuOc2zme822rX3sGbDEF4Mawq2CP6g9
vJ1U9NbawaYdyMYQ4nFebA67y4c4EbDY4KzIR8glBpwgRXCKF5RDlB5oAWvl3P1/KHNUU5KOtEdj
ND/JQSNwso1uj+rukD8a5LIx2KXKc9UbXfSt4JcEOlrdi9Bsc7+uK4MxcWh9vRURCQGhr8O2qHGC
jgkgH/xZh6wfQGsHZWRTm+tDOBWPghy2uk7uZgpMH6daylPw4xlxxvuWKG3K5r10Pkm0LM4aJy9k
3+VCopPTabXfObn9LxgvbR4tkkIQKprFUNj8CJF5G2I1HOhiCUslrzG9C0Z+a4QlJ43Vs16wkq4z
x5spCRY2TMbeDDpsL4oO0Vq3eV7qhblhe+0x+xZnhEyLLvHeyOTNsp9xIz5TYfnP2jGFedwCIWI4
85jvcW63hZe+YYYjLbYz4xPa0LgSe8D1I3jtmjUarh30kaIT1vLZIMBYZV4HSfyXYjKaX2E90LTH
ZljjFmk1/Ixtcl7sTW3VYZ4hevNcZVlq0tYQ5ckCTqmGgezjTPU08Nc7YxYoNnWaitbRmzJmPge3
AkQXMLltcqowmOsQGauqBzk15yM+j8OGukGuGvcfbY2yHlnAhxXrZMsNP/Rcblh8wNiBehxgFp/2
jCtSxnykNFRc62P38L8FGb63qv4YYwLqAa71I/F7XQW3hOTx1VjISzJ62ZFQo41OcG5JmbzwFQ+e
CkK2J2V+s/E06NCt2zToCKvPJrKX/QQ1Vl6GOxw5Eod5YFEc3GTW9p929OQRS5vq4aYn7bhmpIxX
K7PULTmVKMlKNOz7gcrt2n4eR1cvsEa3ln7RSWRTLCzzwVV0sLCzjT9FuJrNlq9y6jNTJWvkLgT3
cvjo2KV/KVE0Aua8Az/ranNtHouTtb9GTSBsn00djP6/27xaVU2yg19erMTtU1ypsvDubkYAJy8J
cF6coNftM+n4ZworZx/jtClREDMRP4QOd8DupzXfuX+ZX91NeATYkyqn0ZbG+9OEs9HhgEHgZKvB
BOdCmkPxa1AHAeZonN4phaK+Mm+A19UU02awigAA3UVZo17YqMxOu7ZR97Pi2rqJnjLrp/XOyv/c
SeYcPXpdtj+baidch8IK4ebHmpO3+oX2lwyKaiF0mPX5H4cKnM6JYy4kTlxQdaePfHOAuvZrVG4M
+NBjXW1fhM/+sSP2uueXRqTa0BCzSnEVWkVnlX0oieRv5AC4NGnd59xu48eqpU7r3Pf/19zA1vYm
mZbgxvzGHC51euaauCVCP27Np9xFWmutunHSXBvuHRumwF7CIkCFFzQbTKMKmk53QQGQbbWCMTks
abiwclw6jsorF1HY31uXSHYEsNndfKEFJuUvhW4LTO/SMyD+XBv/l8dJc1W7Jpxgzn0WprpR9axy
lKNQ+hseDmm4sSjv/EuQFCXsWcDZzv6rAKMXyvuzYAzq2HjztB9VAwvKsWkB/k0UIXBPYstmYC6h
+Uj1aRW85nF71085Nr0UB+Rq2pN6O4Q0KTvhNGyV/lsdkOKXTzDVpjqjXl0uhocCJEtBH9fmapTo
vh8gu5UQRHQQcIwpy+mV+7w0i6Qlv2hx5uMNmcJ9msJZUC28i5yRsXAV0MM8CFxa6+A9ulDGavac
NV6gGP3iGfb+WxRyT4QQ+5WUqtskTovWPITzP8VFAwLAbO+V71pIb8G6YkNorKbf1gq5iY86JToa
PALDZJdAVCG+kCQcFT+aNfntgzZnpWjYnrMsvDZqUiIhg01N59f2LxxZlZfaSfrF5UAzybV+8wDu
DlROTSATYy+FTwnusNoNvmN0dVUMWohqVrynz045C2tBlMeegKbLFKDWMrfZsdbZeDquUGHbcjAI
pkz1DNZin9RqZFTMbBD9Vo/HpWCtCYhYiW+4Ra9fHOKunI7X5onVTgpHtaHmtehWPeC9xrogcpkb
JbKb352m76fVaHRX9qxo4+J3mZwRUJbSWGz45vU6FJdboVfx5dBsTGaxMCZknhtgKr0daUWMJ+jA
ow6Yf6BnNgpK3oLEMrImjYsL32L1o0IPrR361gogjDvbc0RBgkOZ95b331psPPdBcdNpBSvC9HkT
zLCxIiqznYrZUODXFR2HeSG0DWEVAe0fu4VnFr2CQqi7jHVhTtwsoVyHCL/h4Hnu6O4KbrwmH0Av
YhSnn2LmV5YDZS52ezZ5Q+lmeGtkUu5G9btU2jdEhF2b9lynLlwk3b+nsXOJ6HxOOt1bib8+JbV8
Mfh2zVakhtgKEzINorpvN35nXfmIT550TaXUnfg/S+lupZqvEo3EDINDfSRHcG8gJlkBBr8yci8S
sIXFRY7pbrKs9Qi+aT0xHOmgKyvszfNgF9iYpqhhXZPRnE77bztmJ1N5IPrtKfq36u/XEQSA/4qT
ovWmUwHFS+CGqeVjbSmnuvLTAEwS2ENEw520uqoXKmqnR49iT79lPj8CygvQE6FNIYHUEyimXTaG
RriP+w8+JM5k9QcdXb/kMfZF92Iw3SUHStV34cac9AHvyd27UEq5+LfyugEpkacZeyTOYvos8vti
eObKzesFVgrATursOUxAxh1NFwLOIc+NVWqwAWgBFctoepwtvwDvXESMrwpQKkkMcv+Op8OoXbMk
PWK2xzQaj61VyykVWfnwqgXCTF8ieAr/HmS4mpaI/tnuHwf5j9FKhURq12XDM+F2kKcQPzRS6o+8
b5G87qnaRW5qafkz0mGJxG1+GaQaji7ItoeCi1hu16fIFwUfc9qYDn5MOOLyJDrR5xzIQApFj89h
dru7QWPj0G7WWbugp1T5ENmWSu8buc9oFw9Vm5/pe8LT43bke8OHBskT6Bc+cdXmZun9PmC8fP1W
5KD1tzp797u/mgczjmLQR66erg8LwUDe0RTdNDJSn7h0FyKX/WiI2BfXKuG3ZUn0fyzL8sgJQOVW
Vaxx+WZlBSoEbNB6EY4gz34RBav6kz6S5DBzBAreIyjYxLEGB3H2KTpL7ux9aUQvVCyEWKKSMKLt
i+VtPSWLpaaI/5iBuvzMB4WQiMOFAWVMY5cA4bv1X4k7JJJjSoLV/vIFba8U61tKD+aMo+KjfDgT
i6SIDEDB/FdDVCfsKQw2SzOfqRwkAKrFuriYsNjv1Eufz727OdGY9JFHATUDsnlURd/YcXMCOiSM
oWG0bobK+h8rPZlipV1NVIGFf3bH/b+Ef8jO3WTXHgGSK7f0vOGRqgJ6lEc+5aPcbRbXv+6PSq4k
mCgrodN/8BjYsMfLIosIJEzAQANNZlr6Q+XTR3D+U17uDF2x/YRUHObjp2Tn2rJhuQpL2En09z4u
JzirioVk3QEbss5J5VQ9sub5SMzt5mFko4DdeHUjsjqLCdSp25HvVuC3woYn+iT7uiljlnwtKgsS
0aloWRH+XS0JcQycsbeeI9Okac5xJqWuu0EOnRE8gIL0CvOG+abNfUdThwmiBbVOZJLybUVFFfYV
x42DXAps7NqKUM4skCkdYoXFF9+cOGgcT8mZevEz7tMoDUG7Jtg9K5PR8rPdYjxDGVTgdkqhadxf
u90dHjJn2aGR2P1q2+ZcDvkehGPHWIZTMkkkfWutX7rJKci1bg6NQlDaY5/mA3yaV+BFTO5z28Te
lzXx6r1yoJzMptlxBapztfNqUQ5okp13y34xK9IFTKheOpLxgS3DespdWxNYTXFgj9J2+GAKHTNo
1js4xcpizCDsTq9ja77Iu8mEtkkYuxAMGmE0jElduLmvU8JXVrMwDCKEAT8CLs7HOZAd3s+QqWwI
KljyPB6MDToYZLslh0NEK7/Zj/ZbW/xEr30TpSo5SY+u5wRLWp1QR7paV3QiuL57W6ol355DaV6A
+uuObFFDlsZ19ficcOUtK9vm4o/EKZqI9GSMFwXpbTn/jsA0MwQf9pgaAuR3HojnT+sPcji+umPg
4KsoEgtP94qVbPme8F71KaNwuR1EHNRXH3Pu9Ol84vThDDQw/21DNkOicCvrYeJDqPNBOcsHEnPH
tobkGpPlSv+V4gJoJbfMzTKoX3CdgEZ1fbgtB6bStRbzhSi1cYfBlsR63JZO9le4lH9Lj0Qamc3c
Q1dcrcPNq+jll41SxPDxA4Le+MPJN1Izca7NtqzON7El6bM4EUenFK70CVYESC7lqN97lS/iJeHF
qnnr73JrUVZdYYpRKa2ic1tWDuKIDDag3y6ScS0Gk/YfQ8krMmLYmKkFqZ2pa4EmyUJYu2pMLMEB
jnbV6pBw7+STAlGN2rNSNUj5Vt1z7CQyGLLzo1FGFZ01fdv/lVkuoViJF5x4ZWLyb1rbXmFVgLW2
bYnTaDvX4xUvxpe6hOCeXkpvu7JOgfOSczm1w/77vtizCwHoWDCkVxe2o9FJYqgq9UtVvdiYUxQC
JMgUMIDEymWf11RL+Ry6t+8eSWwB9omjUlNZka/hPoQn4PVc4v+q6ZMhjkrqyeA6nm/fj50qensS
L+xkGnz1ZSwYi3ZraQ9a+D0E/xTYUU7v6lBuX3q6U0etWjDQYLEYcro0EM53HlxMGJ8nhUvmxzWb
7qeCelGXl1ab2eXLO1yDVBzPukPH0h24PXUN+uFmXe2kQ2gMjqfGJS7cMeuKsv1Kwv6Kqquvx2Ld
likcBJ/yMULFIFY/KM1yrytualVsJK6rPic7m0tfsoE4NtKiAeH9+vZa7T8h8swUoIsN8wsp2aIf
Kc/GEKIRr7NE0WI2ZV1V4XP17S4QTEPlqiDkbH5f4X9FB8vQMDqM7UtSYuqk0oiUxjO5gcMjS0X2
nbaYSiMR/ei7C+WICUgP7tCdbdrof6P+sK2pQmfLODzjXViO/0N1kOYvLl6ywdp/gDKkcHi5v4xw
+iBhD7XkvzDAbZSBoCpyZeTSiGgWzNfA/F6bpViYkCCcOXy3YKR51EI7rHTpwHQUieJ9zn30/s9E
453dc+t7uZ9lrT9eSL1F7XjREA1ZFqmOzjMdmgvnxTtIUi12y20pCOxh6T87s4nxmIq994jCuf19
gxYydst1xbcFH8MBMJHMstYSkBbrYpPpyfsKjc30FrwxNW+6/RmSLlDyI3CAZA+CBqXJnp/yyqHx
DUE4PAKJwfYlITXfTq7ezt7oDD7irLybb16kPCBZEsaaKXgLQpJGkNHUIIT8WC/BCnSIENroJUYR
tSHiEFa5Xkki8oey9SAa3QSYXFMS1WelLb0CQMNunaHG/oVszoyblf3oR4Qaginnmxz+3IGcNTNv
QClWUI4ITj+YG6NrDjjAJ/fRBKAMEK8atAn14vkAkRL4se2z79VT9cT0J2RO4I6qZUsUPFS9vX9w
JE0HiQRY+9yCvfnIJVEe+bo+s5VWk4zFx1kuQdXHqDdw02RcfzSF6baSEeFOx9ifqpt7T8UpLtS4
Tcs3WiNlEoH31wUAOlulrdQ976CcCDV924AVW/3qJBPhOFzAHo+tXLz+2HCEBx4UPvQKGlSprCuP
eavOxgzuWIcOG2g1d1d0kzBnLtlXC/Mx9iItEuZ2Z7+i84d1C6wUG/Bw7xnsux2hhYzvu0PVgKA5
81nOpX0mvfvQzvSZxwXZAPijQ/INAZNzvK9aam4qkB9JmG0GFOUfX83+gm55PHCxrUthFrI1GIlL
n8Cgn4L/jiV4nriYtMfGQ2K97mqbz/Q2LqPwBeJ3dvPc3NsTnouFENwHOVxnz7wdl+Lg5ZhRgmp+
OAwcOiiPV+fvgkZoJz0NZHv1uxhz0l+O1a4qzOG6zAaOwrz/eqfRHtRwd8UzYC9vg/QXt69wbkM9
FNpPZ15jBNW0Y1ygfoEp6/0/78XUfvkw2WoF12qohTopBO8vy9w6q0/voWA87ixN67ang7Af1BOV
AZMv5BWsdksZWVovCuBHvpW3PoTb9Un/2XSELrglHUkYTBHOIgMzCIQn+1InqeI96fQYWiGs8/37
n9GIkONoCwDBTnGsey74/o24JbzufrTAtN6gWO48l4XkxFxyJ3vOL+qu/nRvw9gPTZzOR64/evzq
GIGb26GBGW+8IS44w3DzBFShfgGlQWsJJdfwRbMviSg2VaBCnuPAacs7hHaZf9gVvLGHqeRoqG0n
Ynfd/KTLvqDqBEsLWlmGaSIeJt/9uiOh2ZoF168zoZhZua8AoEE+rT6PJ/hvdcUOkX9hAjvEv+d7
priir7lY+4+MKflT7z72HaNpT7Na3+d0LUi7vkrWuJwjxHwLi8bfhVK+oFBkFNVX8zxd789wr/8A
jP8ujmJv6Z/Z4GFH32HayhesPfJKiBuzQDcarednZmA358cyI1m94OB+8vm2KbfsHTUe0xayNHez
Ucq/d1prtoWrfkEU6IMSDMGH7GpHiCH7+4o1Fq5aj6mIwdD8+haO2caj7KiwrUWynvZ78uxOa697
GE/Dp9ua73Whmi7NihClDHLwDaAxEgT9tgo2QnH595POWEexz7IFMuZWYKhrTXPetPGVzpk84A5a
HcM0uqJXcnCGzJe62v2cK1AiwUGe/S2Drucg555Wy/pHkd/jozj7RC6jXYWEztzBas3FeWuzWDlE
QFMcz0PHBQy7dZ51wOSXmlNfjCO1xJchgwEZeedhn3Qkii9depUzJ+ONR9s/wRDjYyIWD4LourB+
lpL1SoxEkzYR2bGynEhJm8XBmGSeuWhrtwx7nY4EityxNGUlwg171zHfnDhF0uXvtXvW/QP84871
P1SAnlpLvwwY+2N0zlYR8ziHS9f6BhZmITqpN5oxlGXhkwvjKbvcjONMhgTV0RA/AfzOxUhdOtRi
8FFmBcOHBR82iKmN2hG3f8r4xgk+dp0FIbwMcG/ZgcgSc75BbVze0rYC9zL1/KCd/NnUUKjY0jwz
fxGDkWO8Mktae0EhJeenwRszUBkHh/WZsWvMyuLc7yxH9WcjZgclDb54rVn+mRpmftVKMos3viZu
L1tAib0ChP0wQ6zPNGvmi0hsLikkt8Cc4wfJdLY0YK4TeitwDq/+ghtUerzYnIZaDpxrK8bGswvj
bvwMa8hNolt6Rn71F7/Dsregj5PYmiej8wKEw7CAMvJ496Vuo0gFPOkuy3iUO/YQiYBLOSziz2d4
c5Ppvk7KxPkcUq8qM2qHCm5505/ytpGXWL2Vn0Htua9zeGlU9eFPHlPB+Ihv8bGdcQHkiE7rwZ8/
gH+ClMeT4xVSbpSGt0fXw17wauPWP5zBZpg1ks6gVba9IF+tw2E0xt79QR3reuVIML8GIRlRU/Fa
ix+eUwDj8f+KyAfY146vCg3FUge2B0o4QmWwitADwIkd7GeSh2vikSPdzhSDMLGwBIsDg6TbXE2s
EBe0YVhyq3rLlBK87YGvbm84hjrWJvDCTsjribqQo/NEq6Oc7uZj5RDjEmaFzqc7wr5DmeMHESSG
SNY1QrA9WQ/jpWXrgdUVopUeQxu0XB5XWhK6tef4O9/RYJKmE/VawyCGuaYFHqxhL1fdOoGi0zLI
PZMQST7cw6pWf8XYtTdmXRRvK9C0QUUj9OuZjLWw/0cCWUX7MP09DedQesGf7bdrF5/3NBIOHSSO
4hT6EzajMNFXxtseKIr6mQhksCr78FR7ybfo/JDarko5C2a0gVQPbhl/sgIafCxue7uJUXRUrd5P
x4Y5iDGXCxtR9Mrozn/Yio2gwevqCgAnHxXiz4oX6TL+2tpyQ+p/NH5w/rc/v9cdPLdCluWuj1aE
ATSlWpPNMMiZDFhK9AGI62pt1SEZkgPv/2WhxLlAGz/j3o8ngG6FOQZZ4bw7rviTDnxKjrLkx98S
2KEJQ3AlWNRz9bdSXCn+ZfBTVexk4SFjJncV5cOLhJaXgYGbz7v8cmOlkUK0Dk0bgyhkXZwD2rZv
uGMW+4zON4jHDuTnPKsMC3OXCjoGBKkbffvLKy8g9D3kSIYFoYMWIYunKp1LX9hS0tXcC9NrXsnz
dznlL1HCCV8I0Om76oWp1jyvXnxReftBJXD5bPwIDrYv6yBJxZTfzwPggrVON1bPxHXT/Fu9qMMH
rKkqb/212TS6XEUDr1m+n8LBxtEPjd9Jo517qjEA4X2FDJjwQidyiXPI//T0FeG9+W9QyT58UCGC
uj8McW+/DKScM1h2CsXBXyd+xZL4tS5GLc4eKVpe0+fPFKtiCEzL8r27GG1crBTgHUqvvdLdiZap
m0gpHIZL137czEmvHIwSwAyXvt5/VJGUQMLOmk0o63jmhd8ML7yqkA7hsjtUPPBRYw1+f1ub27Hs
pXO7a3M4nsHqvW5CKw1+vE6/Fd6VS+3w4BI66K5i9OSiHPdwbcSxhLrErMK+B/jQKNAC9DS5ZQrr
JHeciCkiEUP2EU7CdzjNCFj+z6ymYiRx9QN2edTnmnTdE+JhM4huyhJaHqsaXbxgreKdGLONry24
tO/2/60vzNkllrncTZNaIDVQ3juFkeHOgSIJ9Z8LCnk08H/9eCtzLWv6UIDHXGqfm2uzcPdJTmNE
DkcitVMNz7zxF7wdLCGrzqvkKFC7sn5nbcp3J1VeaKdp7UbMNYX0+0UZ+3IR46hcEos6xaVVWYGV
xNinTY+r2rW/6OvkkEaVwXIYth6jbM1wFkzMS7TYPWyPul/X+rPcaUhvFdk/CmAYputdBQgFDNvM
ETN5SigLV/X4z7hslz+4MOxkHQFwFzZoWCc9qYMQjUugfI8p5Csf5ABRQjiM+DST3Y6xyS5MVDiY
lmE+0IJfn8RP23d9orz/RHV2oWNIi2RBO6Bx7LA2vQCpVU9+xSXbTDTwFNhFdEjzp63neIju62Hn
MMp0HKH3WdQt9YPklvWtE6hBR89MPDNrYtWIHH9rMRxEga0uLSFdLlnGjCIx4c0gaXFQi1TE3/1T
+b06MNgUwOhnHNDlhmnijpQmGOo/10e3A3pELG8gcgxk6RJQ5pYs1rID5lKtCToSu30wfIV5zLJH
X5btyhV6wVzY4prdz8lMuoOEFkJ7QI24eVtxRK9uijVhn/Neg4lfwgQGe/b0e0JH0MtpwP8pGvzQ
xS+fNAA+ysDrHG9p7qUn7SQ/pKMVLfXDoDMG31IxwAfU4JXb4UmzHOylDwsJ4MUHL5MevUPtE7ZP
3ZODRmB/60I4cJ9p9KQk8/368xB3Wr2rMzIZTMI9AhjZsVsY452gbS3eMv3QIa4Yke8QNq9xBoIf
QqdtL8IcQyX/EaFeXMB7MfDWsIzttaxQBFniT7sVdLz6mGSgRIljKmrCrUxkmxiTK73C0Da+WLAy
dhszK9HgTrbCn4GhPXYSdsEYbEUAa5mYXNwOZpq/ffoXyeI86T1A9G4RN37ikmElH4blT9gdffQi
kEPdgQ8+jPPqGyGeSoEifOBY+W4a0ChEvbMmFGNLDfvy8vSkRU9+/sfDShbsSEdzyfhXe8MupToZ
cigKo4HGFajUaxokTWYmdeB2sFIxh+kGesisXBSQjrpT/25f7nT4INs8IamMPfYIdBdvHfmwCcPu
n5YoFgrrrhiquu6q2+me1FGbEMwHodE4M4f+AuPFz9wx4w3TlSCQGscxuMxC68RM2fKC8IpeljYM
J9vizuUcf7VDE+jx+0yj/jctQs+UJmEUR89J80zeE0n2su3tuusHJiJS2t1ApNjZsDVWYT2+bRKx
pq/xeqgm80n38Olc65pID/X74NgTPMXiOYYAiaJQnjzBWeXYLxyD9oSdjNJSYBiNA7bHK0m0a+O5
7zwdjgMqN5C4aymLSsGa9aYZYuYb1tGNRRa+qi/6M2Al/aSm6JLvb6+XOZv32Ztg0ZlyC5T2dTq/
MLesgI9kcAuGLWZKAf22GtxR62LdAn5xWCL2Pyig4+oPX8YTBLvr1/zp0hPds3qXQN9rikzRLJEY
TeZKNL6Y0fLLcBBgZTLTovnQqgOSKKFeO67N6AshtsEffK97BJ2/4fSZd8nhsf3YmFOBVjq8IyAt
FxU4DCnp/SY1/YMY0z5gmnf+N4w4KJHDgbeY9o/KM3o01tc4bwD6aPSUv0cKspV5pGh4UMIGSASx
vNvdGXHfGvSRBfIoPkzTQtc85PKMLddW0Ke7pR2lWqgZQ6Xgjy6xWH3kHCzS/exWTWSh/JLfq54H
v4I44WdEkobOW7EmtzHV6PmXPWBEp32CLrAupu2RHD1N4gmRiCBfAnxqsfg03BNhhjJVI1Mj/Dkv
OQgIJtQ7jxdFrp45Hs1ejhtApN9D7OHYc0Pd3NI4mvGLFv597bvdDshNfcwOitUKwoKMKJ6pL2np
P3xsIsD6qt0Vz3gw6dbg8qXoWmCl3wYXE4OjvF4CO/f8e10f2I1lz+lO8cWomTcRTwbahteszi2J
/QKjaCcKDWrXTLNQ0leOERPnQbOr3y68Ub5mDLAcCJQaOISwHEy3X+wrElS7Ca8MhglnbPDn3LXX
ullL8PdmEATHoUAnm4cVI3eC1B3r/78PPZ5JyGWGEEp/eerh+m5N5bGxfgC0+v6+B/QujdUUZZpa
t8s/wnxHD47av4LjEYNegtjaRU/UX8tBtqZgSZ8IPFyGQbswYAt8iPLjWLVawxiuDsgzXKIj2omE
zdBc6Wl+bIQz70jaSFTbmuAOvvO4xq4jXksK6ZkApZYgZrwB6ohF+yVyOPLblu1hwCF6XBDRdzdk
jyJZk1+zz8qcycTZWZ6vs8OV6tA68P91PABZmiN58xMOXDn8PGUKK9q+JdHbrcWksNvducJ1+CgP
Q4q2k3HqCtavq1Ish/GDjRyXKZ1/AEDdNSr4qlDIh+KpnWNJpm51fdPiGia9K8P7sB7qUVrk6vdS
JmM0cN4GE+KnzGlQFthjAOKo0735a3MhoIm+f9Ig0SjSE/RgsTAPyaOkznxsN4PUPGFDkDTOXShy
1GdMqrD0NupmEZs+Y+qTYprbL38zn6LjNs0uWfQJcAn/iGJddaLLYYjWRiEYdz6nbmmZsIH9TS70
6TFR8tHq5Zo3P2sH8wSK+/BEKFOKsmHKqnGvXr5c/UfJ1LjCAiFzeoiX/n3mGZ1hvHn7jrq4alEP
9XvlrS8X2SToTs8THcI4PG9Dp9b4tkVwhXqM+n65DJXhoLfFbYjoRhLAGp7TXu64fbLC26zW6Ikp
HBP8WbaNZLZ7QPtkpB7BPZUaTHcnM0NG0BeYDhxiQGQS2mnijf0ZHOz5Btdy5HNGceHPvb/qNjnP
82AAVUe+oSUOEQuCwiGe2RN4IDJsRxbv9v3LAdXhV1SrIawSGXUlGY7l8rV9IRpjwfF5wZ2uudHi
ghwuSGvEFmYkal90X4pBZv0kOGR0Godzmo6w29Ud2PBSm+USQQqFybGnc25tZ7BDUbhAwPoBs9aT
2fmVNFXnpZMfwjH9yxR3/ek9vJYpeI4CyBa+56YhMeHK/pFcK+4NuIvEFWdOo6Vhw7gOMjrPp5m6
PObJQamktZYc5VVKE3S7/wPO+cklCc0yYNXB8OeSfiPZh+w5tMhO13fQQBjqiroWxGjj+ID1C0hE
NNt+mokNDlRrAzzUY/gEE79cK/RVx8gJ6P7fi65q5mkz7SkKFY07NkPDi7oXVDsIyGltCLWjh4jG
a0dQEgX3dN+Y2aVU8uvFoYQOfKg9QHgoERDoxAetsVIrgWSqMwKGWA6B7us9KlwlqjYnz/PqkjUr
ebyKFJ5F+Y6DB8xmxA30lcduhuldK4uGbng6/uXyTTuaFq0GuCqqBdhymZx1kbV1OAF5ZTOXdeNe
yC4Wd2/S0cwOSQi3M9cy1awLcBrMHm2QQYA5GzCyRMt1FgE5y6XvNbDdoUoqOKBplCHkbOHMxvha
k9N7cyXsA/953WcCi7tNJG7UvTNTrMfNPCfFpzLPC2OWSxUaBWG1hlwMMkjWSM8czjMzxwfjUv4V
aWokfPAdXh1T+fXzGYFUNbFugKBITok1ZIqX61HBRhKhwcp6WVniXtBAezPFsN1EK4QhUbmREMPW
lMKUzlwQTlV+EzdDQNfYoMlqONwmNZMxC4qXb99Dxc/MiRNQi2CSQalGeENFJiZni6PtxRIte4Yg
bBleb27ijkHxHZhm87qt1uZTK+bbUEm0MKxwPVSc6MTeyQYOZHJeC0QQXREOCtm0/DVvBwLiPnv2
nKiEaS0QCuTioEOg0t753hYyBlLwfN0Kv9NG+gtOkrFvSGUkQYpzMxbbB0Q9mxiyjaMHmdvdfpkb
+OXU2Q2h9QaF/4kPPW4IQBMrbRCWDEQIFNUl8IkwUkwF9IOL8ErqrK5DS0mZHgNpZhJN+xmCnrsu
Jv7dsU/joy6+frfzy05jjJLxWBR3LHyg89ddY19BwRfNH+ZjXDYoYUimN/G1BdtGfyGObQT5eN1t
kupd7mlI7VOnQY0In4gm4v9olPUuJjAi+0fWjcjOBPKzntywAa9QwFLdeGyql8Cajq+84Rftj7vI
5WtcnQw/Fk44zB1u2dDCOYYGdUNCI1iz4GBwo48/OknHA7d9znkqwp1w4CAbThfP7hQByUC8/A6Z
AjnOwe/QSV6QKlht6E0P2N+c91D1ZXC7YOVxb0zrBkYALAgBUm3brntYzfk50DqHcqYXWDk8D8xW
BFXwxJ8rEueUvkcmKOO1Rc/Yd1mIEJzaexqqwltLJ0NgNcnYKtil2t5n/9zzxdGbReY+kKaC/g5r
qDctF+rbYMzItU5c6qnochFKy29Lsrz7zQKxvZraUAcFF1YBwNFTOkVzdSQtsBJvPkXBPgUXASF0
mdZ0uSZIvQ6bCcVze7gn71QcuMZQ9nj6nIOyBmziNJRugXYiYJaPb49/OYgrV4GcmuW3GTJRhow7
MTd+xzQJWjkUBY6IBVC7CJ36QKekTMpNsIT2MvN4n44Dz9aKryUjjuXjPbmZuJvtprrc74cAU8gn
mPo2ZWyaXPTHJ/PgRvFm7PW2O+/CakDQNXsylGjE490VsSWOvj0pqHiFPC/QtHAq9ZsGxTQJGftd
/NhSTju8UoN4Sf0mARdp9ReLHyIrnFOUNjMFGAXVsg+WJQqOV9EwTqofPD9/tSKl90yfJd/GU1kg
KgBxqAJc0V+kw7sbf7YwPcQ0Vjj4hfaQNFcEj0njX2YLG/QnDBe0W9mUCbRQvXKU/nZG8RJ6y7GK
RQvb3Kc4PZ4YywIV1NAv5NXUhqU6+nnNAqfEy+EcqYg9KGHJTTHdZ2G9ISjU8i53F5Oo/Po1MRjT
Jusy/TjkfkXaM4KjdLUCLi1XTS3bah4V6vbQyqCePTEUslInQHHHId7VaaZ9+og7ZP6diKWld6sb
99fnBfZJWjCTo7kjNRT6//qx18PbEYkuEBkWXhhSfePpnpgTIWf/xRtpNknYtHuT4VqK+uTYrMPf
3qiW+pQBLSe9fp3SI9D/lqqdathFLV98jHz/5vpcQUQQArBAmB2dsyyjCygpVJlhhzlXJKJo9Hxe
HQeKmO5lkw/Gbr2a/fUDhqST+scP1059tH30R/ojiS6UE/cD6Hv/gDPBmrODlPmEaB0iT+6ERFmU
NJLCOoR+YMVV4PjxzN9RJN932/jRRBy/MOCHrLryoNOezjApzlkw3cVVhycfZB2uRnrMi0oIvCuw
NSpdZqcm09+bXUMto5zpm1gvkq4ZosJoZfMuJfQam2X/J0zsFzKlRMfDK0FAtLE+w+bo9IpDPH61
g2qpAh5Ja3j9EeJXqWVXJ8/3ctRhlC56iZGz8tTJe72Fx1lRoGmCzQE2HmJb2NfX7S2qwshd0nzk
NCqAJZJbn2MCBQ+zFzRqKlR/5Qr4MX1Ke2icv1Z65Bg9xOqguG6kQSffM214Y1sCFsVCIc/V/AgE
0dfyur6jd+ZzttJCdJIilCnDj5R6SMU4DmC3CwVpt23SUEd0IEKFrF4DyftL6NtXW3VrfFgu1bZ+
drT+lOCmj5LAH/0iZ8YOeZmK9JMjvKztYQZIV+7jo7PrRsrebJhY03ds7z0UVb3ek8H9KlAL8YsV
jc9uG4R611YwR5u9DFd1Yp8AoboHM2Gl0aqmCkhiO3Ku16ivr8mQJ67vfyKC3u9FPDyOrlI35E3X
HzLQ3kIxc5FBGjdIUCZvIYLPb+qTvMKKfUy5e5ihC8jdfBlUPG77aCoG1jGjKovwKDTM8biYwQTl
4FKHyw9x8CvgvhSwSYKwQNOy9ndvypUj4L8CcFGbM1fi+0N+r6vXnnzcivZeJszMfji52Xaqa0ly
ar+NUJZeG2qWhmYVR/cy9c0fat1FimQikFK4eFDmqrMwVKy9LRvhSu7fqDrtBQlBBxTd4+KdaChc
CsCCwBDQ12Dchyc0uxvEfkukswWmkVJxRtIeD04xMYpnSdD05t5QkRtdiTo85HQur4syTxopdaBP
eq/ek4JeLvcViEWsyxxbwmyusyg9HO7RMk5iYdQmvrQuzQz+I0APHPs+YWNnR5X0plOUskwnl0uh
+n0kA2i78lg+vAkmgbfhU7giSBDR1TqQZPG5EwJFuLOTo5fO/uab5va8XJ4TEgxca07njOTk1bjl
3oftN2UWEo8t9cGs6QGUEMcJyVlmf1EzXn4Rn6l0nY8mCfpjm+xZLsiINWF031W0So5JBLqVBHmR
ct1fjPJdhe52e7kz84vh5HttVuFWJv9mBO6i41Qabk3TMpWYmGu0u4BXaF8jYS++Pez5d16FIk8P
miTOi5B6BGM32l94TADzesWNcbQpzSSqYNIMUxd5nd3g45beQhsLsc6QuoA6yRG22J89rABHVtBH
lmMh97blplll8XKF9hiUcyxtY5mGD/xWuJd48l7G3JlsKD3cLSz7FZHRPbVHolzRaYBA4G1/9/sx
/3u2gVTqkpAS83Qq+ojlT4296NbUQFUgKGqEcCjdSoYKp3RNTw720t2WDLV+lBhUSkFMwhq2VMKz
wC4nr7gjHu5iYlkNJ6UYVYXHZPBOzI4exSUJD6Y+x35C5KOnaoMHGmUtMiy2VTCJe4c1uDYfe6FP
8npieGZYNv9qd8ni7QVglUSLQqX2xe7kCgXvO34lJanXEYTD2FfV5mS/TpYQchMbfjB1fleEzrTz
roQcYnN6UHCdNnWOtiH1ARb4pay+/tKOsLhcnE8vgjDi5FJUs0ZhfzYDa0LlDiqNYnWXsWxuNrgd
wxi7oaqbFN/SY6aAnTcUfyGZhvimSuKqrIasMT4y+T5QLowdx7dtB0AQz87lNPOvQJsuW6zfR8Jv
CpeDNvQa0PZC7fKBGWcBTNe6R1qObZyaODZxLWVtlY7x8xjWRa3m44WGJ25XbtJhAPebgblf1nFL
wNx525hSusKiSbPL8vGyOU8FHeuKVVWMs8C707ZCpVEANkLEYaA2mhPIYjP4RISlnLn375txtKoV
CECh+qdsGy4sXuXWEcaVYDwvff+cTyeUF1YicH5fKAdQFgFxe9nqcrLTfBJGxk1NHp3DeSOQbQoe
shoclpCm96fBLP8KrSOq1z/KQ7uMjR8wNRuZayD8m+3aig7jOtx6rDZE1X4Jt3nBQvoDuzeS6FeK
MyOX0AZ491lY6ke4w+Ia1Fazac/ubow4kh3cf/CjJDlQDHU3107SMl548950g/0BQsaXL7cmRdEI
0hcWi3dP3Y6GVqpwarKUGmnExN5e3x9Sn48XwF2GHkjtIq4VdbQN9C9oivbFxhOz4JlPd0GKLmel
JPxYMppxStUNYWKMP0raJ7qC6+AzE5UF4Xr41JOop90L+s+nnF8dtYNBe+1n/jich7ZTRKQPnNmi
pMQDF4BfCoyNpKLnoEWDKysx9vw5xTyuv0j2EKjrz7uTitHp4CITQ6KutApDiy5pqzquM1TJ4f9W
cv4zSI6ZAdlOoqGU473ih1Y7fcBhLaBB4opkj6Qf4c/Bu4LYODljWuvz8/Lr0TPVCNcEEiYPut5x
bW2E8QrIVj6i2hmq/pIqoe7PE3QxHJaazCHWQ3hhvjkLDrnWL5KuXAYS/YU6gO1prWKJ+rAiDGdK
DY0ZJPUDRwYsMuBWLwt95zBGXLBeUTzHrq6RSfvZiO1JSpCg68S9aBrQ+PouotMyvt8ZDqjYR7bV
1WGZxT/ygD+2F8Z21//gm5R2fEL6/jHHRs1P8Am1scaWS08Y1qnw+tn58zGZtH772hpIqZzJHbTW
/0EiZ3o0DKlqS6IOGgcSp48OYebgHUtMQWFLLzSOUWCzEAyIHekyfcB9jQH+yDSyC4MlFxdwJVsj
qHECnqxW88sbyfpZnIA6vaBt/KnbRbNhp8T43LPV6kn1K248KHa9EyL8I5X6mC7W/PtpgZxPMwOQ
xF4r3wAIvr3OD5ysB01Rx/Em+xq1ay15F6lI6cQG5vYDZaKIBt2YnD3oqxXkI6BJzVyo2oxZyBy9
gfeBJikWeeHvKNkBLnSx2hqeaeIwVVzwQDJfbGoAskx4RV2s1/UmYNsjPd9frI158AKRmuIrwnsk
wIxSovMFyEcnioXet3rvy6DgHsPLNGU9WEbzl+LijrFh0InYtAo4H8xX7ZimmWlyh5S1EdV6dXYr
aNOUmj8krieCUTXB+UC8gOb6xTFwZEKcJNtBOs5NKt/lnT6+rUmklmcLjtLKMfvwu96cs1APNji8
bESN/a1LXG0bRos0EmEw600h3CgwGk0xaULgSXEn2qputGXE29YFmxVQ0FMYMA4Q+SpsofJBrH3g
my+ntm50JAI5ejd2Jz2t/3AXQw1CMQFHT4zQtPwg3kqZRd798Bp6qJ9Qu+XZmKXaR6lYXvGn1caO
WabyMsohy2LM2a/oMGEQZX6qsRZKCjNX9cV72M4eZZ5kPNqnImBu1iATrgHF69XjQHgDlxVdj46L
Z2g/qi0SCQPjwNHGM3dFM98XBVsViYJX84Il+31GA6N/KWsVrY9sJ4Vdt7UqObYDO85BqOiVrc/X
PlViiUz2M6v6a0c5w9kr7TXKgoWnd15D7EyDUGaLwIVPfPBu3q8rxUF4Y10NLIpWeOt8Qma9Sk63
Gua/Np0xAvXF15nRcwaIYyjleyX78E2qUsmT/FLUkDBjbJohoKTIKIw+KQTc8vVi7RpX9sLmesrr
uLz7E17kr3dGvIIyxzI4fdx/3iaRfuBiICNVMiBpajfrPyoHuGsabWG3/0oVIdQbVaJg7MMxoI/n
BCjlD1Ic1EjLTak2FPWp4uzzTiUMNha+O4gKxBY5O2oovk5S3td64uFVZ+FqG1yoMa2vB43bo+ek
CDA2bu1FXMchHhsZOvqix5Z4Gc/PsJqMJKrRhyQBHFoL7EYsZzCdqc1D1UF8JlSxCPg/K9OA7xW6
BHZY3omYkYjCxgSaMHJb6MhSE/CPZfc0fLuVhFDD7JJLEqI+4HgmVaHf3RYqsZbOisw2U1gzLvFi
r8iyZSxr0RsDfcu/ddpL6x/n6/eXASuzNsrgr6s6oVyroBno6OCysTGKY7lTbSbmWl1PvA731zwN
UZKcp1TuRqflna9hA6f5PxyDFW3Xt6f2KEXFXMVLwcp8saKtseWB4dLpRPX0fJOoRuwxfcJWXpso
6dbp4bu/Y4H4ODdsdfJ0wdzFSaYvaefaJaALAPM8sJUnkAXzUy1Dp3l/XJHQZO4knZ5KsWb8MKg0
/YfdKKMGIExrCaFX7nG1FET0Lk5QByF3W4posmYA7BV6KQZg5ooP+ZZMI7QMwpHyVhxoPJJAq6js
62MnfJsHrEmmAWSS1O06WyfrnWS+namVvuaSNbmdZ8IrlaPlLPqA8hV1qLciEP6StuEu5q+DOkLh
v6QxX0vq+0k10ZSWkoyys3mkoJ0rdc74trcnVd8wwD88wzJQumeZT3ZQhtEU0x1k+8CbTRy5wdMG
5RG747rX+1r2jaLVNQy902yObkeWJalV/rc4xabppwSM76N8v+Jl+x/XNWvygVUjfoCx5Hc8T2nJ
1n9kbgJDVtS9yRCWt/uqTbdm4wQN1xKP2BDsGmJOytgd896Ri+wz6+hCOLCl19iz/ivjS1rGwwhF
UEC8CUdItsIq6257Fc05/epbHznwPaI+2wm7uEE5n/rbPlpQE0e6An7oIr8VjquewQ0+W+Kjym8y
YkQ8KTlOTlJ4h/yBqY0N1NNoFFzSNxEwsNE2K3XjDqMAU4wuQTPWfirO2B+VV+2EOztC9eZbg8pZ
r8IK9k/1l6sWb4QSwJZOo4YsCy0kos87sH27yddrn8ASF5zjTDmah+GRm0uWjeXI+nTLb23byxQg
82fNbaT+YCctfZl8aJEmeU30urnpelGzERCuxyS3G5k1O0mbugv8u9wWE3AF1TmSxJVb++FjxIG0
1iGyregMfNi118sfXEMquHctgk/7cRW0ZzZlwE2ZF0aKfwtV9WpJ6vtMCkHCu5qedp5owKxTC5dD
y9lUlH1mc+ibTIUDCSN76Zlg1UO2KlBXQjmVYhsk8xlr0MyKibU8tu9P8kDVgfr2RGd+ZQ0Y6fZA
W0xzYJM69axlhmivsEIXIgTg4d+2llC4j+Y2OUFHI6L4L66S5cLrAo/msmsgeDcd2Vqcvwq6CeBO
LDcO8Tw3ky5VDKjatKSFGEwrABpC91tJUP9HaPsYLri/U3tcIIsBah2hOJfn1MsoDPpbq/hrluFt
cNefBbgJMMeSlnKGmZC6/8TDIW2kmGle8/dzb1/fayHhJru1+2NsgUD2m8gFvq+scltX2t6lOdkW
PCIsUnfDJefOTJXdKicRG286CqUUVHQVRctUy+OziJePbcre8eEGhWssqxI68+4298uD7R2sKgTX
L2dokI2YqHpvsyv6u7OtnGy74kSCAH3l7iDOK//SCM0A7Gbg/w3LBA+fJcOZNoaIEJ9TyDTgPh/B
eysdV5LNPNdArLYfY7yqdfxlzuHnkVBXh+Q4IS2Syr9RpnC7kNJn0vritH6ANWDJ9vDXowJwL3J5
BPN82LIZH/1JcCzGfxRXVdIZl3OA0INL7RO8og+bVHID/squ6fC6ODDmAJEXvH6ocerrGAEFwqSK
bmOukfaJlyzZaLNDOiMxo17+Mth6i3e7Fy7X0mBdSsW7M6PXbSPmYZ9NO28FaPiSbI4rcsn4b818
f9LGSnO/SoyRiXrSxChsHsnkdwiDnvPHBffCpiTo3+FQfMeo5ZMbwhy1hmFqs9CVxpbViioovrqn
RZjkUG+Kn9JVMY5XxuVV+BT4HpmytvAW1iD3CCnC+18PCcODeMyvn6Qjs7Y9Nj6IRbfbxFo33RMn
L8xEJjGi1nxNcBBF9aTc7qhBUohaZiGZFYtZjNrcuowoYEFnNBVUYmotdzyittkqWDT+GzgwOMRK
LIKqsleq6n7yYH+BCGzYuWs+nTEtj5VWhxHRY/x8MeF0ahUWn5tyhzQuwMEK4PqSb5CahjNklYxr
TsZ0oqy+G4QDqApdE3UnSESzedlk2HlgL0g+mIHzV0WItQ3QWpte0bE20x0lzBkYo4p2BnZCtIy2
+9eRRfhdPa1shjX8PKkVADAY04cjrrFLEQxDvhQOBio2EL321TQjgluZ4QawSEYS97bmXDmPY5jF
gnGn2uvvwpWcP1DFSyKXsDrVySPnwq4rxhDoMaM1op7KRCG/8Joe/qYB9CXFEq2ndgJKKVduYAvK
RVv2BOPXcuv07gU66pmaXZuoKwaM3rCk/IPbh4Kqm6llVoqN6SXQVTY3OUR1gJF5bqwGkOF6bbgO
XHPbQBtQW/Wfc5Qt0ech9QRlNAjnkt2KPUGAugUCH/7keqbJ6b+oY94wtkxYQ1MR6e7kvrqdvlIk
D5Hv5DyxmZ+s44Yj6nqU8c8DVJ7juiouzS5QVM/vTT74Cqgl5ghxWMk/hXUK+SRglygCYv6UJquz
HSGASkafEwo5f3SySYrmY2Ay1QuXOm+md0e7EOrYh68hvnc14uqvSp4ScEt9fp4SFOZXKWcCh1cT
WCFkginc2UNDZyer1+jR/MmaHMkaF/JdBZnJaM/bg50AwfZu8DEFha1N8G+X+cfHCkgo7h3eDmUJ
fAlPtO+n2d3yjDfJFKu8eOo07BdNThBYu4va0GBBNvL0Ix7/1LQUp82UVLoOKkq268sIYvtL4bbQ
8NbcgqqHfMRiESrms5B9PPZOpPDFfhBsGWJ4PvskjPQPkPeGRFadUq8J6itcsCwRNNu8HYjpfYH1
2dMJxePw98RmmtDFLFq/hYe1aVUsne64WYww5yn+WJdzXLuD7RY1BmYCi8aXWAzNgr/vs+SX0jR5
XG7FUIBhv+ioKwg3SJaH1oZh6+9IzXGuU0M+qWrxnPy3tk8mLuQcuhdiDDcSdRrqxdUO3GvdMa35
WvM51xScsF3zeNAzIQlvCe3H2Lw+qK2TL1KqZqkON3ZbN/UR7wTl1zqCEuBsYx4LtM0yuNpZFkFe
/b+9ELGP4YPIvHO2TMGNlHPCOVVrFQq4jZql9etfC/sbjMhxc7PzQ5qijTEPl5Hr1eABICBsFhI/
OK8SQsoBNc931Dt+Pf3BLpOR2gmpawspiJy8mQhKIIA2BmchO8Ag69d4KhnMKhhK+2VdZRtR/qyZ
N7JInPcoqedhCLqBkg8LoLueQzYBaGzVsKMDUPuWS++2yiQTiSnwykuh5vV7sd7NW6zDu8fFLt3T
vs+L3s52/cI7qdJjDFuCf0fRdSnyeOVz5v+hEwTYbCMfHUZ2P1RQXvMuk5hEj6fjPWjQoD2lCGdj
7OupcAbMHnQlsDx+CITe5YRiHlii2T2n5f7iGeXEjvEoid1Ax5LHq83lWVrm7qXNsOMM5UpI7eT1
+cncudt6HZ2PqdXIEBqjrGSwmpxI2bMJB6L9WYlnINoJGL3mgqpn1Au2oQ4AK4LHEW8VPRip5vLO
Okt6V9ow47g2l1Q5Cnq1WwlF6fV+J4lAf9jIs4agO3jtTAdN+6OpjdRI04ZqcVQ6LkiWwjp55OfB
LRSZT7/pVUIbSob4n8EI+yaw+32pG8KNcYtjkarZuBraxnmK5BUpxAw0gbpzJfQ2/FJnkKYimKlK
8We2Nck4uMtlA/95bYMU57YCuQiU05+nF0ahYp0xYDbFvuzNQM4kQeB49MjnPGnIjmglwbuz8frV
K22WAbYW43wMaFIxjRPuCzYUY/OudjTYFrmlMoi0Jv7C4XqGAK7caijRBkfUSefrKL1sldB+x/jt
oqcRWQelDMmUlTjlylXU6KG8ueDVCYDRgd4fLtGquEkCOLt5mf0P1wjrKeTPhwkGL+v4yRQj1VLX
UFqPTKcYGVQzyp23kHC24Alp4JYsvTqIN5g4h1rbZm7hZvTv8ucIHjzfZ2Awk3aVDDxIp0J0HKuu
lAmt2cG3xAGaoa4bRE9rqwzxvCcnJo8SnRIpQoG5WOWqniuMaTQIK9qnBNs8WBbVgx4Yes6Pui/b
u4MmK1Xff3YWIwOP126smXchQLSAVv1yOI2yStXCe7MGyD8wQ46WUMRYV6/nnoulCVFRCWPUQdmf
MDzpmLNANllXwZSCSR+RkxS1lEYNXgyRh2JN9OltJCR7xo8uP88e/Mi7L0RpKkpJLEjZrR/fIdp4
vFCS5rywVUjQ7LdtOcAowUgNa/41H9xamcqN9vvN3r0ugjs+xcC78/oWDUAIyhd0TmNzWkQey0I/
Ri2lc2b8twxP1Q5Pnr5/f7NY1z2GaauLkELEc57lftEmie4xEgBdZymaxU3QpHm0r+yAtcCW5oPv
m30ufv8h7OfQWgskOOONMN2TuvZtezbm/GUYnPghDlr/rW3A/vT+NN5QQ4BUATFSgGYYrJxg3+64
wX3VhmskwglQtp1Ed9R1ahNi6R5LLEVRvYpn+G/FIi4G5OBEZXVWIH5L7NKxl0bmzC+Jhq9EI5t6
tBfZpGC3CTyS5h/2F1DCKQZN0BX3NUKMY5+ofKrkjwkLPl2hua87TVU9DW0UB2K2nnmD+So1SBH2
vESoLLNBhjaDwZyih3kv2DI8sb0/T09e2HdfNJ8flxvHfsPZKgP3/rMquMNQJlI2nUL2qlLIqvUR
fN4+GsgofrOzjW8W8XU8365o6wbwXtKzojbT6S0rkQaBzb0XzxKKsIlzdOGIWSmMl3fdnrziwsx+
qK/KnCzN/2WDesgHNlT3K5ZWp3fmzUjwNRy/iy+bnlwTnn3XoGQffiSG4O1JoJ/1Vaf5GjDshUTA
R2w47NKcoWSwUycT2FQgB3tyGLCDb3hq1na6C1RXJ7nPzZ1DfxUwHtYkgaGmul/2m5XRlhZ3rQ8d
um9w3Yd0RvNkQD8nevcWMjk43pdbOL+TqWtryWNJ051Vu8wbZ5mmibpa34lbl+nGfCl7qjspbpLg
ft7Qz5OxtoSjPUYn4wLtaCGhe+lsDTH9XWYAMJ07orhTA5k7XXT3fCg9/ndsjjrv9BjjkTGQHiMe
Df8CoodyCgLmbAhT1FG1l4SUvPUuvq2CM7JZqdbB6yGZlNvkt9bAhRCIOudPQTZFleTkjSFVao/Z
Z5jRyVelG+UQh10neyhpSptR91b3t28s7TBMVvNAah1M+Pu+NhMCtBo969Iwinqcau5rVzeGyBVo
fYIREgQ772VfaBvLz+maTII+5T7ul/NqM89gRkAKOfhToML/SUJVRqHntc0IhiEE74u7As9scNlP
pGchD/6x3YQqdvzZV+/KCpHQq1I9WovN+s6gLwY+8DhWKStDDUAo5tGZBWazJynDVmO+VNOF13sQ
hDucFqilraiO7w9RYeMwYdnNGEDDX1Zp3lXqyj2wExHg+oG7cVhdXEXFcf5Hb8/TudUSnpmgE1Wk
dCan/bN/m6UkMXvaIkX/CnQiGcKmkLsnv74XmWQ+/wc16z/J9zl+KcVyZercgkFvjBDIcPAnrcY0
wooLz3iYkZxanhnBjjH4fiRlmOtdHr5RZ+F8dEr1IKSsluySH5SZojBhPCwzjp8i8CLjp6IbAN/G
nCQcnSTlFnlZ93PJbJe+n/pFK79s2hUVPhXZiA3h49W6NHD8AR3P5QlEp9TKD+8pBHi93Mi/C/Gz
gN3yB3nb90fb+GRp0oCLH5Gg942Z5xo2KEqcnFt7A6Hifs1lbNzsHsg7AsLsqYsCNpCuxx8hRoEs
aNFwX1AeHsWTsF+ywA7IwdIUPyiGhgDcgRu2TGTPePo1zyF2j2QxY28rVjYcfKBnJxdLNuOxxxUL
ATLny+++b6xyR2o4sCrg4TM1o+fAZ/dn1Lp7WqUVKk6+oUtq8Z8+PeiopM+TXniVNtML2G6tr/z0
cUPPkswiPdUG35QDL7/R/1rT8Sstepxm/cFW7btJwlAJ6BNFxI4KE4k0/pKO8tcIOq/tdYc7Zmct
LJSPhSQzocWA9FtQHBgIVnIH1ZSFKQdYTycbw0gatc8q5w7EE57I62aYhRDgaWIFB199PqGHSNMX
b0hi3zXWETxKbhFTMSSxUIijxGdgBVXqibdfF+VyJGybgg/e5SP4vVSEfslLge4uJt3b+RcUcO0g
lofUXQ4gWISOpi51PV0f28e2wdgpWd1gP/+XHYOHbZ5S0jSDftlwCCKMfTSb9jzz8wjQ1jduOjLC
AQuknYHT/fAQJrRDcZl0RY9sjkwLhkdaQWqaloqo2CDgR5bv9pEO1FbfGwIGgCwQ1O94e6oC36fX
xseI5Gjq51GVJ+3y5ztpDgNZT/R1X/Olbegh2noxyObTdYPKau4yulKYAMEws6oxEV6Z1KplTLhP
lj0dyajoaBd2dXY4P4w9ROssNj2nGCJzYv7WK91F7LxZiWi/aYbGM9llHoZynq13jvphBZgSgj84
nhY159cnJ+9+MMvTFPoxTDmrhS8pkeA2xZLv6fX4LmoT3Aqg1vhWEL5lYbXjDA2yiLAoCytpWIg3
JpVtRymmrvUiThYTAZY3u/rhLH6QhYPelrGU+T6Ehb8/gPKUd6kMo6xqtKWHPMnpRrGPxsSWVAIH
MgcQtPTWVW2LKPpKuijqYsS9pbU7jNZhDMMdlgvXzhbtBaPXznf3OQJGel8VzfAwPjl0HjbItHKr
ZkWqtv8+JBavG4Nr+fXvoTKMsIcYSPehnhnmwP8fjApBGKC5aFh51y9qFp+lrq8uoc71FzdbiT0M
7Qpvskq4kO/Tjb1nMakxiJZKmjU4i+Yjes3zajfs0b/V5LFgZfvRr/yWdGorWahaAggLReBmtWDW
4V5KCR5hJILZdi5sK/418W5i4goxoiqlO3Xl9ug4kui+6KN4iL2ZF8m4onC32Z2++8LyDrF9aCqd
vCCSvI83TxFj2gcVcwDIcy8Ak4x5xnl/4tLSJmSNldGs2InDgiFFc3jKYMRrwje/g9tJwNrYiZuD
Y0tNnFGNiXzi6bbQprpX7qu6LwWXNGw/2rQNiITKfm1xX+DRgkW8TRtqwlbzpWT4840l+Tu4iZYI
8GTVdcPYLls1SzveZFXBZ2rvlLRdtwpaY74bxXMDPsvpJ6LDR51l1jvWbXRE8JvkX683PVd/PeR/
n1AvAJdXArjLM8sQYI2W/ir95sSG9zHFp+czHMYzwj0m2HErNcEfhU2D3uNkhc7QzCzErJogS0Vl
tL0/Nj6F1GYy9rXaedhhXq39HXa8XH23ieZAwH0eMF4T8hV41eRkxJq9RZMMKdpXMSTddH/Me+Bh
S0lhSSpoCagDpOX4jM21hNqGiG0H4vefUfSJI9AIE+MxHd+UnFhtu/x7+4woFO5dV4ufA8bgO7Zf
n2jSQIj++gimb41hpWSys1jzJuOZEJsDJKl5JYkTYNNCzd3ozkvFZTa207bE6sAaYM7+8Wlxgbfw
Fmup+64uXH9SLYB5HeQ7hMwaU20gvCU0XlOnElpnFZLeQyb9o5xAhmnQ3vtJJVOMBJPee15J8fo1
j1T5ocrzcqQaULLnQ3uxva1hmgGXy1FsFOKEOAGtfsRO7404e22A8rcqSG8uPRyNGlVsONBS3XZo
jdsB7o8dO1nJXKuspOyJpYV1KhJdyU7ELomsPh2R5zWYDwvFe/agIear+a8CV1tsGjzH6pN6jbnH
cOy7ykdgRYHxJrqe56+C5bl+26vExA3rqO3qaZgtxqShLLtSAZZDm4NX2ASnlIHgkOxCTzDENj/B
+SCcuGdqbbh2Awt42cIPTbwlueK0PuQV4QuU5JkaHfTO5Mb3aLWetovELOIXDk9nl8x/pl6Eg5et
bwlYLnFMCeu39HaWAcGfUX2v+2sTK48cpU0xJ0gWxNLiTS0fXARDhSRUdWTTXrkuD50vPcsETeb1
USO4ocTvyn3g11eTtDUUp8rThXvvAnBnaSOfOXPgm0NgLIvOCr9s9AIGYNIbTGfoOTFcvyMV+0gF
+dhVFQzzw8rpl7n8yDYB+yHygrxc6xovi3Lpspbmx52C19Zf//WrjW2GHv6+Evpr1GvtN1RK+6wW
NvnzCpW3Z9dq52u5zZ+AJHsocAdVr3rB+g6ZLFGoNUliDiVUR1nWuN2adjxSzGLHXozkkosJnoHb
AYLZGnSSpVr3Zt4Vt798ktgE2VPGsiV+V6Yk5+76rT5mescS+YYliqu+pF0YgzbkwxJJHJ01N3FT
38fIbNMdD5v9njDNQxk92dQUzXzIMetY7v6H/wdIW2TrmD5IHQVNaTWE09lEKrSMqR+AFIwNbWks
p9QAhPhMkuQu8eTfyRvG2dQnSJ6hSLeVmUXlmYS5PZ23KRaMoqBzY1TO8sdOWMJWhXh0lYWuyZxp
X+JepedOKJrDvM0QJUfbxDKhBo9pXHsh8tN1nKcW55QPRlGYMKNl2/TTwKLARUCjj0r9Bppmj7ZN
qarzu4VyGybVJExpVKWaQ6vmlbfkwrBUQnhsrFXo04tOXN5hBeJzaSLhhEiv+bjtQN4QFZHHhkog
RVsx3CSj6zmaNjwfCaHzwWlIeokFqmPW8yNLlPQeWIiBU79Yt80hAiOwqv0sIhayeTp4X9lXmDKQ
3bQENmJhVpiMUPv059CryJkbXkPkJqm3FF7/d1ewABbRSFGskZ/BHX+KH3Hjcn2+M6jqDqz4kXD9
6tS4t5+HG1MTK2E3Ow/rHtzTZACO1kGIBKQc2xY9DGHQq1w9z6IygxDD2Mc0Bd/tu8DVmchU/8aI
iUKLuUomKpDjkvzJ8IZtAs4iVRB4N42CKtU8RlKc46k9yAtx8R2SMc520iXd1e/L49lHpiQmHVfL
I0jfAqiPPbNNzOgj5pXzEDypxir4XTSm/3gPbKgayXRV0/kYNWPRhDZIA6S4ssJYAIRw80CDWABQ
ZMFBl62p6iQ9+hwFkXo/TOTefMI8Fj4xNEyviRGhiy6nO6qVTaQ1C+OBiBTlOS1esNHOnXTjc1Ao
9HAN2eRuWjS5Y6pNnPQOsSOvkIk+Knmh9IEE2CbXw3GRSiISVSItPWbRo0rQi0aHrzGK0Bm2ceQn
1J/9TNzz0Ta2DbmYpevZFFr/ykXz3jpJM8PtVBHPX/nSxiuO2kn6FHuu2L07RFMzi8ZbrACg8naY
TEnUgLmj6ppnOMa66hHTRWlsImi9YgyDjlEPLUPDP8X6sz3DaHuaj05AC3Zbs6x+sXcNUX52xJY0
HcI/N6pL9Yp5WTwl+6cWmEDvhsTLCnkjjUwD5QBuuUQU00NhsimYGYZZhmNHkcCh3mhkP2AzbHQi
vmbLLzOjqF7f6Mt6d+r2iiRB0F9MaaUo9/jhfsNmI89Glz/CiTv8t3raP6xnSMgSxeG43v5/bxPp
1lFquVM9R2ZABWqE3hETllhCCRFdao6PF3tJrZwTfjp5Sgpdu0Et+XtUg8PBzAAFl7sHAWmii8X+
XvGLV8PUsStfmRqVPdSvkGHvvCc221M3CYUIXCrFNjhlqhhV3lwLz0ls/OmcD2fkbtxAIf5hS88t
/uThJ63qpbcqDGKQCwFgnWfOEQwH7UX7BRjB734FEC1bwqcEh87VJ/K6Qg/kF03xpS1LY5FVIMIl
cNLe8A6QJsD2Ym+uDTjdc1L0BCwdB6wYZ+EAf4rt49I3VFvql4M62PFKXpcZ4MnQLfzHiGEC82+O
6O3TlE1GMh1BwHLVTv/BSBvUye45QgGGqVBI+20I1MEb5YWH8sW0OQcy8fYEJqIXKqVwp7tRbIMP
cBcHz64HND4QUtXcQ7jsUffDmgUKu/txtGAyYgZftG8qexOAx9Xdv+XtfdvahJzkxx2mgAUybuOf
ssG/Rkgl1AwCB3Jua61Uql2NV/XDC+ZhYUwCV3rkmtql83e2gf45bx2bcE8IDcFpdguWk70mXyYf
3pROdBkY20ZFZVjgPgNkKEGfahBzsGORXCyEmA0Cc7Ut7yiS7FUDZKyyQQVZcz51oT9Mk5QZSilG
CS8W0Zni7pUqjCwwH2Z1DsnIad5BpBJgxMR9m1At5v+r1o1Tgg40BxJM/dgCP/N1EAzLqs3yoVGo
A6B344qRNDoiw6qVEWrBmrN0E7tmV4IKypZnNsA1/m6ys3WJGbIAQhPWK17WdwU4a2cB43w9PCal
wGxNR1eOjtwD6i0RnUHXJEhANipdFTq4DKSaNub7CartJ34O/ZtX3D+GJLsq34W7t/zNTpdEC+Wx
H6hjFIST8eQTRWmBGuviEeDS+29cmrxs+PxPhu5lFgOziPMsBmhcPPzD1LSxzQ2cOtTjJ95j2omB
oOHrTHl8U5aAecz2Tpua3+JxiYuCyE6v79ZV/NVdALL5fuiF7uaUNQR0kPyItIeBIo9rguNkkmv8
Qs7WA2bxzbxMLeb0A3qsMpb+41XEk2g0ugN0YXURjnO5nPfORgE1u9IinGHg/rxl/AOs/30HDGvz
FO2rD/qZFNo7vkag1b0rZsVxAKNkzoSooad6ZUnqzQrg7U/XDKKpuqtNT7s5ggNobSNZGnDW8MrP
TpQcDNKuFpOldS5mGuklDnK4RqL69GgbBr83WC5SCsAEI8FZIibrj5+Ms/1iXLdZoYjoBL70ljHB
xUnVN2zndzxXWMrXtu7tVlS55yHWFUxG1qwM2D9234WOtrjmJPIY3vhXUqq/drandTct3yC+JCuI
Vllklu2ZQn+SFCxIQkp2yKZJphoIcnluasZs9js2bKKch1fmJLNufTbZGxUQjSGVx9bu1axMD7gg
uvn44IrGXNJ66atmyPUZFg1c4VJtXeww5afBUD2+dfT40plbZ4Jw6rLHgyqMdJ+bSbyJXqhouPlr
SkIycigd2jK5DeYnXGPymENql4Fzp7A1NUu3syIqN3BszOqdQIr16RZpstn4oJpgCN8sCLnLFVKc
+6Qf4amcfpZ+Wu+gEf/9ZOFUZknHBjJGW8XnBrIKR7407LBHCLzCZdEhPNOjTNbv6kpxphRuaH9l
I0HrvxMKdmfquGdRTPcO2CZCRYjWMe8hPx0Kasw1oZjZzYQbA0SO8iTmPOd9UjwOeLQiGfVNHfzO
HhcSNKaAlgguSujcAD858DGe+8VGq3lpVH3WUELm0rsT8MSSVOrjEGtJWjpdY2Kkib3T1F9w2PmW
GbRcP4C7ARUocBfWhQT7yWuv9rY+e9JrbuR555Q5WdmeQ0+WfL717nbaAnI0LzmVrzIJxZ52mPpE
6/QZgqDxND34CvFbM7v36YiqWQrE2jp/vYrTsBu3pR/OTUrWj7NhD1CtRaVjRFOUpRJhFd//45ln
q4FnlrsUQx//CtkftSstgxhu2UBMYUgaMKsUtSjzV5oqurV+vWfzL9EoGEVxb7GKIAYDgaOkGvAp
6nt0WbEbShE3Klhn55hhoXsWB7LMS5EV/lkB3HnUZ9SN5NWIrpA+tQBGHM/UzaCOf1TqhNtsca5R
sg4pSYvdDvHL7A1Iz37llAfUVxCQoxv20rEij/lHmVkmZm1tSgF1F1BCgMBfRAQMg0ANIYk/Hsp/
Yh4KCBm1UFpO4qvYAZgKq1oWc1c3DEViazTzLVz4SGByCRbRSZn8lEbKWxL2Eo0SY68BH8Uwhz6d
ljtAt8qeeS6CLwntZnx711AOxgRgvrzJ03A+57nDGJxJ67O1JB4zPmQqKu95McPtLLW28nxxuOTx
CQdjL6rr7BbKWVPx9mIdF2xvJJrqTWQ54aY/VMocfzMrBevf6zDCaXa1HXXj230k6zlhqnXwHhcX
bITlzGhhfrnZkJoUlQj9hpdTQnPxpDsLoGb1emMZGafXdZlLd2sI+6mOYWcSKS6AasVCTpd9I0mf
2wFZYRhbbEHhcT3w3xxFWll5HPvNdzhCEAw0x9mKNgwxnTq/MmYPXb3uEUY1EKPztESmoZRKf5L6
hYgYSmcApmk5Y74TxtFGnDY5htPkA8meU8Qh6MKjoI1+lVnU5ex0D0HKqhHbH1TM/BDPSUUCPBsf
mmozDB1XTGWMIEOBROnKjF5TGhhixd0rHsGDam8OmlGvjB9GY45Ou2VCYFFeLrmEmEYPusf9v/NA
O4hDSHLDovqT0XQFnPyblyHPORjkYWph/Dhi9J/B6oPq3n9mFt7o0ZgfSk8csRVxF4A8DcmIp1N7
ijOSob84km0D9ohD1KdHJ0ZE+3t9p//D3AbxY60E5O1QFbI7gr13HUDrieyQaQfbUuFnupwwJSYC
Nj8RMxeeV8nQ97780i5boEApenu7Ev758ajEFN1lJ7ioj4HfCNxtZDsSe4gx0jYORQNWdI4e28a7
34CuggXghnPMQAg/3XGc9V7+q9nRZa98S2rmV5cwlsMBsq+cTqIIkCxvx5CkEgZA+2f9ShFRHqQx
5V9Phzt95ku9qZvXBkSyrq86gLrk7AYqaC3sRKOr+qf2ADpR4IHjLSHV0KJbEVNfyo6M5VVB/aib
WTHNxwe8dBTNfMSi/yoBUsQpM15w+sTmRVL/3sB0p9Owx5gGtQuqUnAEsXZd0gpjHx8ZCqGNV61+
EgHRj3SNU9kb4F1LAcsus4kd2iIwGnYEuGBs0Z8QZipiiUtd3/tXN071AweBUZ+19qnAq0iDdaEV
tX/nej8nrLNfLA/ZSLNCDtqx28ghvxPAtE0k+iKQHs9PEaaOki3FURXSMfZe+gMQwuVdUP4dAVv2
LhT2pIoyOirkbMOpgP5rKjkAZ7kSjOhqs3EUvPA8xY3zVPw/ZYt15T8ZdJwdFTPeio3mVlMN/tec
yIIzvjrgergomWydjY4NBcIQP3ui5HEZ4audDbd3+XrjuosthJ+g5DUaN7Ihj8sjvRTP5b0hq3vB
GCPJLhH8tjF85fZDKMOamGtD5dT2zYf1J0+JvkK23CyemaxubGEnGaqHGq3loHCrH6J+oPPtvA5C
g06vua8Mgv1U35L2HGAO37I3aTwaPzD1A7Vx0uqef6FIM0STm5L8mxJXmV/19XLHp53SQxaLgrG9
ouPAfDLiFn0JJq/U4RkQyDqeot0+MdnlnvSq/vqQDLg90fJAoBdpT5s4gGeJziSWneiJlDqD/rNj
rNFlhYxaYpcFKIeC58TCQ1+qubIY53nfQGYSz31/B1IBu+lCJmRl9ieNRSCy4eY0qSvpa3f+H//H
o/AO5Dymy4xFHCkPyzwxn4ptC8x4KH9oU/GK/hgIEHEQ+uXyoXfYoWO8RzmhH8rtXFw8IgwQV/zx
PKFryduHlVLoYFIjcYkyFJet35Mz6g8Oivy6qU8hUpb3qOSSnhBW13T+11Cfdor0E+kSmKUDi1Gn
yuKonux2cvrKEiFfUEXLRqzWjEzVlFE6ubSfxYLbZJSo0b7M5ORlDCD8PbOGOq8pfbefkP2ZOmDh
GfWY0/PCtnyGWescmdxcTj9my03rmrefCQAgGVz9CrTblfYjP1BUFICha38l1fK+9/Xp6epZ/4L1
vBzY0OR2uQAq7x2bIfK9BQzLDvXTZDx8KChOpy57AQZQGeQwBhADyqSBH+mW2GDcro73kr2cWL5Z
Cr8WYgFvd7GlGY7EhMur7iEdpiWchKPO6uEMxXsx1gwXUPChehxLd/ipQ3/zFw0gjHpbWaVMoGlj
uEe3hQLH9Rp8HIEskuoG49LXVdWcca75Crf0zEVFmy8rWpHEw5G6NmavJvrSfHttA6X370G+ydie
XKwtvlqUeRYSWiK1VeL8bKp2jrx08YIgW249dv88jcJAtFNI8re4xOoLJboiXKsjv0p9PebCvAoe
EpcEMk3XfwVUE5ZdaYul6DpBX7qsaJvlshOAHsuRpRtFIGKC06NQV/Hsyps4rvMloj3JFiSBbXYS
n5w+bbUN/RAkdNmvrqS9aDaHcLBUjrEGwb+kKjZ9DBUDOVihPUDYVFQCncpCf8QHwJPi1WUj0Bd/
Ybeb7el0RkcGeIYETxn8DtT1An7pqMYL7feiI7OqCzr39GCHDRDh0i0mhkYqI8dYDavgcpIW/hG5
f2ErWF65HutOW/PrPMRz5xcXgeirme1BdsR5fgaVA6Gw+Arn0/GKMTSbKmOzyb8jyv2Jk7FKEHpb
/pKdM0DlYctotNaEfv5Vnvuv4nd6bvxDl37zHnaxRfLGEaVTshGmKqvmzwakiCuSFuKcNDAzF9Sj
quypog5tUHsdYksfFcp7leG+Hz26JqeAs3aNuQGtgs3KDO+K/NUvWIjSpl5Pvq0hKb1YR61IkJCE
VCxIS/BR7UcbXoU2Y2bYAFMETE7zx7Oz7YL6b4mw5KmL6JDKsVzLfdYlXiRleiVZfPoo+DH0ZnCN
rHLkfzo4p3S4adm2+LGhfhSq5l5lajiLhOWmEdk3CsG1EjVjL3w0h03I88iyTz3r7m2bBsaLWehj
ymsIi7HEW8LtNN+HEfW6sfFzBHN+zGqcV+5foO6M3aBsWhcP8oDKXANsP/zFaLsyVs+8wdvpDduN
m2AvZSNmx8m9RCsfQjDJKQQEeGuI9SJPmLfMOOaiSDvN3dYzswttgiu2jgDpeUNem28aWF4QApph
pot4cJfE2hYHJ7v8i6580TK1aREDTaJ3UPfyCmuEzPhS/f27cJillALF4CnEIlCBHFBNE+OF9t8l
X+7fLywOAfxbuFgo3Z46j/n/rhERdPw96s4gBs1IPx3UC7M+r/z3J+tJEvvfzxi+arfDSM8DWxiJ
ZPg+dyV/AA+sHhqfG2RihnqPaTGUSIvC0EKqiWhf42wlyhzSnRjxxYzgvpId8/RYmvgFN2coQK09
G3tabW67SxA/VBsMZxebMr/WafednxtJ6ahzkOoel7Lqj8G6DgATh2/agM617kZUkN9X3HkuLFjH
AJil0XkMT1TzUvdWgnqYr9XkfAt3r8pxmB/wPgHsFz3H7nN9fl+/t8tHJ4JdlUWFlFWvyOIUkip1
0DwvWsRUhFXffDdJ+KIqd09YkhmeVTDFvwwMGYKIBJgeWNpPQkOhIDHYuOtW26DHubLJ3OosB8Gl
Tg4uhj8qRzytby/haIkUBcTE1TD9sjNqCBKu6Ql5WbAa8CK0DqaFa6bWvZnINcmnmw9vyxBMpr4w
nO/bWzLydjyOxLzGgDP/FL0fN/4nWhuF0Rf9VMLbkb/zywu9xbpmb3oOrV+9l+EEGJio/JtsqAHB
jbYpWT4BCMofqerttdHRSQ5H6ywRYdqLy1DywlKGss3TUF2+LE7sCsIMefF54H/29jq+vMoQOgDv
xLA/T0NSHwQHRwylefeAXLfqeXn18alrqcS6jUI+4twakf2HK90MzCnD3uFTCOy6jZ1U00UAvv1E
0JS7U+UvvGyz5Sgy40JMyPJwgQn2vH/dI+hXFa4ANhWW58yITTe2HGV7qP9u31jfDAAyEk/SC0HF
aZZ+67sOVnVmz/RkFR8YAqUDxbY2UclY4jOfeslS8rkXxxHXCNU1cq+2DJvaT0kFtiD/UlGtyvo4
CfM3A6Ta03ghfbmdWrfWOMDE87RvUZ04fY1YMeueqOyHTTX7aGRUz1gUa85bwu3kHnWa2eqzLUca
/I9q9Tq2O34HBX6kEAUMbVa15HJ5gE1op4pC5FD8MUmdmc8rIMHOzdurom2JvALDC1QtVe6FIlQv
FOcc7ZOTyegyDtaF9iJkWy/5HJ49NFoOlqwbPMr2fd6lG+NnhcvFwb6Q4pXbIe5X6+bq9BGFEsez
Abi9DgWBEqMARFJW+w1QDMccx5XPjiLV+hkUnAYBEAS0jOCXQuZjBNtqU/dD5S4C3hzILY2aCXtr
oqGkuBiUSk/JYXFa8s/4imOOdRNFTMS0ApZ0ospNd4tEGwmkE/TqlbvpI54u+/+woqPMznJeVRvW
0G/eK7Zf1FF2cEm3T8uQ5MsvNLtBPjmQv3OSQ+gyxuBnKitw156CsSgGrzgb7fQivmj4k2PhHQx+
j4B9Cnqt0eZRU+F+nGq9OADmTnGddNf7hFZThHwYU91DUUD5vpO+N9a4EwFB/Z3PoLmOks4Itat2
5DOK1In+CIbLsZZxVj6cEl2JQGn3h13rNTa20GXcfaC/XtRqWWSaHehmoAt1OLoCvlf2TVATfdMl
KRFLHNfZplnMpbsYWIXXGOROhHJLvrXLb5V1pjPuik1/hf3keu1/8udhUNl5+MB6hDgSVNtgKzSX
ShblFd1I0Hs4FSzQnO3FDl7buZpkN+P+pY0m2x4WtsiPg10FBac+0ygtyjGajBNOwCGnvpqLi9Hg
fkY8ecYyJjBEcZFo7Hdy4wFaVF5rdCyJlRbSTDk3JcX6k9Q23+KApo6wJ3bkcqd3yKlNK2Q5tLbx
56UqTsXGNRBd3WOjwf/i/yW/H9sMWPxFrEafmZ0Y7n29vlFllvicOzMehaFoQvCqxXvWlLHMOiip
GBhGMnVf8m1bw5kBG2Hvb7fJzber12//mE1CHhmQPdp16h6lDFmzVpsUHpWVwzFF7+alXGHeHVb4
ben5BtJT0a8REOR/0AgM0DzkElQmgkxzLndA9RxXCGBBgLKoDPzAn30k0N+doNtJRUVkkWg++jrL
Q46MRerRmFh1lcu6qCNW8PeyLCUIGNLNZ5Q5jL5j0Sex+/7cS+/bxf7d3EXrZhmW5LF/aznckXT6
zr0fB2xI48N+WoXHrRjAzui8ptDZKMAWXKHf0UfyJDqxGULaNwnXZ4sexiPCE63iLpxo6C8nO3iy
2KFOxQh9scOYGLAuqCICk2jM54237HJ734J9kPVLNm61mGX+FH32FVNagvMzMusxqGF2YEFxFc3Q
gX+yZA98cZYJPr3R93KaFHgmUGqwBNVMKJQluwaCTLw9Az/zIS0LAhVclY4bvPwNHGLtL0LImmrn
iKJtLHut7rigKbMpHBCeYljV0VGHdfv+T6xmF9svCyv+nHPfk2CDyQVcbP4X0uSZeEpTKswgZMpu
l7OCyPmvC8DOwAqfFpZrd1UW8CTBGio/3tAigP46VPvcTppWxECfrr9rCV2ng4glkPJGdZG2jDTA
8/Iqb0AK9okcBqLpShXKPC5ixNfdavq7Km1ZEEaXeDF5RKoFX3ts/ZCRgoyaDk9hK8QffzXeDXWG
1JN6hhzNTOBpS6LiM9w5U2AvUGmWsC4NZVcw2Xsve5zp/0UvRTSHzKnuM11H6lENxhSn1Ac6Q9QR
dkOkKLS1j0X/Xlp8JAhr/5pP1YFeUOGxSUr46PxBTPaDN8gjgSh7rY1yzwJMoGB/+8WyD91SnnUq
r7/VoqjzMQVDOrq2+ZSJDoUX66RtuyGfTGcBVB/q4fSjxu/xhJEqx1/HnR480iyihx5Wen83jNN2
8XvwWhvWceZYO/5LMN2c+Fc0hlif/r+AnuCYaFeDJ5G02g5I7c7fiPiGO2xv2g6n5mDaRN/SFnlz
i8mKAxffMQ+vC42Ova2NgIUj2JEC6ZN2AXr5i2SKliBiy6FQ3KvE5ZzI5ceJ97szVWP8TKRUvYay
tMO7PXdGmpvnKoRRMdyTV7iYgEHxRZdMWwhwfB/yVnVoj7U8vWFarJOGZXDtS+a90LJuvEJ4pBdU
0r6fdaahXlZNBUL4G9JAJ4VHJ2bLZk1mwug9IyEuXeFVXFa6yKKm3z2BM5xkngsLPQ/564m4Ys43
fwYbZahFRqKfIkI2nSE+1dHMUgXdCBcxtO6dUFMGrVJvIDbM+Bdibo1s3gf/H2bvrNjFFJeXWyVN
kpzBxNsr7e1zigJBcEwAqQYJDsMh1TH4vL1qgzFKy7vreXAHP8pEYb8QFDsiUkPal/RkbANWBUKM
eH2RXKZTVA3FZ173yNnlWxKaU0xpRKS6369BwPgU8sgHWzhP4rR2m78H/B6GKYhDuRrsAFohnDqw
tPUoRHC1cZCje7zW7HKhiS0ib6JPCiIVRgTgipYVweZudbuaIeITBSxtDZ9UltAomsfcFGPpFeDF
csHNMz3N702g4H3p2Tt6OkXBNBzDI213KkojXsfYVJ+dJhSWOeeC767Yh05dT707zraLdlcRyReg
BR1QrSz5kBoLKbxaaiWw51uYvD8ZPvfBkYTH6z95rLhH7yojToYXLt/Rjy3zdk4O0Vt7KNHXxnVz
rAypaua+WGAHsKnKyXhixHrcpuHU8fLbU15R6eTqdqZ+rzjxXbYFiTnlavQGUSYaTtI6rWWfMJRI
jLAxuQ41rNsr04dtcUPtr6RauGlnfXTf2UDLrATq7De6qHEJO94qsY1r/Z5pygguNyFv/o5nBwbr
xUQ1S8Oy8k5ZBcAwb847FSr8nU/B2mBmmYV0iFrlP7URW2LZefC3EU8x3IQ3C6QZ0GdwzADnXiIp
ibV8c6/LAFWgZBlfVOnyEiO7eFHRBz3h8oUm+EAxCTIwUgWu7l65YF9r3NVBCENUgL0BbcqXXKtV
eDOUm/+5doNSYN0pU3jUVlTGN9euvpWgIaHaAj8x0riTFZepOfz6Dtj45PycAfejWscJ2Ew30Ea2
jxQRB4OToHVQ54ZFi/vXvmxwHf+Rxp1YgfXi3GAegNv3wl/PSbtrWVUyIEGdnaKhKMryOb7v0Lo3
7pmA92MGBbZOVLA/9b629kPDvaP9wkIa4Wq7aFMv3ey8U/D6TNpRhk8u51n035ilHI932ESFEOP2
8K9gblyxl+xq70ZrgOeYKSCLHULycHA63SUYlYZFetEgWN7JotpKKHHpmDIHUK6xKYBD6PKD0jWq
E++leI+rmIdz9eEF309AE/Z5RMZ/bmlLFHIPrat+HLtBwGM8HY8p5SokqRl71dhpBSXJC+hQg1o7
WrxDqxSEHCWQdojD9e3T4Mg8McMBuVYFfGE6yxEC3dWEgHrwA6EZSAzBPhs+3nASf0zJucGjNDtg
R/XJzAFTh61xmwhplMQ364r/wZCr8huUJjzlJ6FgLvEpFnWbAsjT5qocESc1SBpo85z1oKIHkY09
n6q2+kUU4Uo9g9FlECo07ZWRJjlVnuSsnRc9PogS6O1aZFwtZZxwrAXbuHnaZBnAzKaPPPHwBv5m
Pr8z+HER/2K/AFFjK9dbT+KA4H6gFcFobWyN5gof48yPWA3wxBHQlGY5rkmVY2nrPlSuI0XRzuN8
LrCkvpDfEsHIkxhsgsTUHuPek2FAN6lG7iBtP2krIodeboVAAmxK5wHclIybHYRlMFLPF7tFrTgC
59KhOTRB7DRbI3cvabzou1Z+kulxWcGN+/Z16oLGbKBbTNwae4pT8bMYH1gzmsXLpFhRT3B8A6On
c/ZdtPKCde7Xt+TMthRFw+hYvOLnQ0ZUk9Ox266aTsF7jYqXpbYz+t92CYuG+ZReSRckYKQvlo6o
saiofWmeHOnY2A2wiGgooxdwjZ2LDKoB7HCNlIJNOgwXa+5J747b5hIWFwjZL9IJ2sOL15e9863B
pdMJ3sDwHYdJ5zd50So9L+Pcu6HROLtCw5M+Ofikm9wmbetAWf4oV0y/T2xyTggBnHfsNWZwfB1t
4rWfRuMCVeqPGgL7cZDHwV0cxjpbU4QdWFIKYBBfHRmP/2AktmqCdSFqSCV/4nD1Ykc4T9dZVUje
AuFX+jSDxvUKXL1S9hbtncHsYgmdbeopqwMGgVCm8FQxqgmhOCVAeLLC5SH3LP8oE4sVXY6JkTiK
ZXpMAwE954Sf+5ccmhYVnlMj63uXfIHWjoRgml6jr9FIdWW5VeK3BQchC60Ka7uUdQE3SnClCUE4
D5PlSZOVYt07Y864hnx79ovUvjxzrFrPgkEYSOzEvt+hAH+2XUC3NTMSSVBPSJmJN7BQvkNIQSsB
+t9l7IqPDdgrQFZ98NELH/UA3pNhjBd4CETv4UBJha5YD6oqJvljCYJG58K6bgqMmPoctVF2awYU
lsa7AgQkgdNjjK6PT/Lgdx69CHKwE8ab52j9LAR84BC0MUjxLVscAlEraJwsWu0nkfzezdy49OzR
SepeJG6YNHZRJ1KZ1wZ8yCseo6XtWAe9LIEMYoayF+u/n9LgMpuEcQIgHAHF/NcEXFxAwdbcrXMO
cUi9IoDulncZz+T3oEULBr7LBC/GNy7N2dKosngvwnQh0CkxNy0H8HDwYVDfgOQLbanYMvbdx1Eh
POZwQItEMceJwv6S2c1R6IN/rD8CTUy9B8D3Vzk0dJ5INXT0Wk9tqSmedYbjjG8wTcZFzp67lpy0
eHkhu9I8Y4fxWtYar5ybE+G8lvMHGNa18ayi75eAhQsgjNy31vpyFoQaw/EHe075+cpJZxuSXAnz
jqqm/AZ2fzqNehm7xYl7ouuYOXp5AUcvuSyD0wDoDptP96VwfypPR+6Ji3uuCmLbprICG6Et6W80
7qCd8ow3v0lEYe8fxRXzKAWw9ddCciEs0oE6YLi75PNdF+9rKaS/oCHaeg5Fhna09QXDf5303CLV
7ywbuJ4KX0mxle6mHmDpm3Gv43YN5kL0QslIuKnWK67hWGjrb/N/mFWhDdlSCwtT7O/XkKxslA13
gGW2QEELd0PdmX1NobeVU7f+m8IZQylnNYTv4pCbyjpBkJ0VEPcUjiXNeQhQZL3Spc6T+puOykMb
lojGQUr1vX96irjS23sMeKJj2ByIev0FlL14mNW0Pxt1ppzl/JW+vghrjQIgrkvZyB9KglQspo+7
pZtbkbsSZJNxzeXnYqD2wJaPeX5OxhH7c20uUBao/cravBUTmXL29Ntzbq0HdkTFiu+Y0KdPxygW
MGG+ELyrKp4H4PDHdtSAX2LIqFkmGlupRXOW2CehcBUZYE70UNNKpX+hT8u+4Z4eWT44iIL7829i
Uv88zweT5K7MwJNV16Wg4VaYxODqfw86/L+nhJv4xiB7skN+uo0TiEGitkH98lSRDd4CgCJ4uH0M
GpYTwiNPT3F6q4p32YYYvIHws/LytOOZhREqtTpzPj1vqiDqGAUtVQT7hRamO865J+5JVN2J+9ii
m4N9lFDQp5Gvl+I+hyhitoCO7M0qPNat1d/uzSZs7nbsRyV4Fkr+c6/F5e7z8oUdnEpmkKQZjEsr
rMkosu2dwpoG9z3g+XfZPdSzO8RL2gNMPYN10OvqVzyVNIsuSOPf7kf3VqlIOOqlTEzHGqPqEd23
uliou93rDBfTYknKmovOkyn3goreyCvIfcWOeuonM99bkb31S5ap10/hQaM9ccklZsGeTwY0vHT3
K49aeNfUwfbV4HtCb9edokxnNxgIlR2OijQ33OzwjfLzZGKVdWqwgVcVxWvKvKfrbcVPCjrNP+2u
mRMC0OIeSk3S1opJLkfVeEO4RXu2VhUw+fYLiyUHu3gLnYEKzYRn1ZQi1M5J9vi9B+7euI+UMTQb
KRsvY5P9IYq6muqRNQn/sVeyAkZc+2634s3xkdRUjlUw1x2ihidCCYov01fPqYgHnY/5ux8xkCnl
+GhSL7ZVtfkr9JDSH3amq0trtLYv9yxxze28GbUYYr1MXizUo8h154LI1wAWx6KUNQ9+kuDjK7O+
Cx5+RsTNAtbJ+FontJ3bZRmT1+eTAO9INp5IA1i0+8fOxmL3OKEWY3YmyNmQ+/q3owHCUKDrVs5Y
7cOF9mfV59dTeV4SngWebXHF+J35lAkFHgrrPZ5R93sa+znfAKSvoEj7ui2C0J5UH2lldhSUFl6d
RZeY934nzYlEUZDz6Y4ZiieqtjWDc7epGAsDMoHMvoi9Bd50tsMgMw2BMEtdZyqHy3b2IZgGvlHG
MbCORafNnR4RHTqgUlynMOkDTn6fK4YWStjvgWDZ1MATbYvljPwQOReNODfcJP365isY8Z+vuwGi
K2CoquLthZE37yPU881oSr5w0qZfvWwzmAs9BE2QHpzNqBcanPIL9uFnuDdNtLc4gzDUlwpThLZe
NfEfHG8D8m0JSssLMvYjXAHG7GN5tIXNUZ6BjdyTM6Ni8sx/0EtcPW7JmQYoBoX8+OQj2ejLqb1c
Vv6OGUPHIqufUDTw44tttlNGvnNV+tB4z2x/3Zf5kHw3bBp8IstRwrQ3veTdlbBvrEs2L5xZf62N
Bg1K4Zq+v62pBHjTAcbpZq9cFG3OREsgaj/5C0BMBQ0g2IXndTeF2FvvBaHg8iwnvudCcwlPLkeK
45YVQIZyQ2vx3nNmAaObqfXIC43aUoPdkYO+Y6UAN8scv6ZKqd4KZBUJC10H7idOidprwuQyPeFP
CxlI0yEZxmNUa42zXBHga6DV/APGnnTL/LAKFfNdDT1D6galODLlbqDTbsGI6fSFB8RG8mcfJqb4
GOCPaDzzODvrvyIKEN/wcnLpl6VBeyLRq/20qliWHIeGEOvxo0lwxTvM7WtXuon2k1SPWJrAqEgB
juzRn+nFKQynLEul85ldwGckLeQ4sX8BE2vrFPPCSbmzsJJ6TXDEyR6PX5K+RhwL3h508iDeaDpe
Sto2S4qSjbjAR6I7qAZaI4jc5in2Gt25yFrbx6g4ZOaxP0PT5ZydqCGYa9Bywp5HqADB4sZNyXix
WyugOIrw4jFtb6cioZoKDmfFnts4pRMxPwVipgBrrKNMZwf2F/EIS2WZ8Eu6whNMDe9jeQi2c31T
2mt2zI5SpVW61V/a6ATDca/REVmX1uILvpZytqFNMUSFwJ6HGsJ5+ovP9dNpPbofeJXeqqxkL4qU
Gu4/JHj0Au925AsURpmz7UXhWCMOsOqSyUByPoPRUXwvwClEebGyUS1DOBa0o+FGtF4m5WHeCYEz
EZ70snbXdbYlP5azHN7LNmRPipWxu4MWSd9I/Lv1K7KCthb/jZwSB1CyBzV66/aS/7gidzgTVRTU
xxBS2wi8OONunr430RtA/OdgDPEfnaneHnq6IqfSmZ5BgQw8LF5wW4BPFAGHVL/7sv2yKFmenoSI
np9zhg42WukhwgYqf8B1nrZ53bHnvrT5UhgmWFJVC6bbvzbMkMmN9EFQ+8Oznsj30LVLFhk/PLR6
hr/C9blFtOCfV6Oip9g3woxfkgE3/4onhYSdsYGTSgAxHLcAbd9U54wVhq+jWGsIN/Foh1Rftlmp
M3d5ZhCnc35sLo11kBgsUNyQRrRmqCB+HSDl1ZSufdt5cPsTaguWIZqi7Z6kmT2iUfIme5OzC15s
zWPKApumh6A137t7frSP+y3Qvg/+aEadvBBDG0ma5hwwmKgQnHW8PcRhyj5qxGQ5gDmtCH4/O4v7
mtxqGh40G9+rec6gIduJng0cnOWpxf9pVoUe2GNjf55FoQhWjAv+e8lFTrn54sP+QooW6vQR+weL
JVJqWvkaRziJW1u8AEU9/FpH8OljIiMnET9ZoFhEmhYTzDLD41FsqKApF16rGAwusP4vUppZFjcL
4Rsfc8LohlH87FPELENQmG8fEhVaJ7Qa7nPMHG4Owk2bsWAGhy4byUC9yMPOu/K6EUPQcJGCccW8
EWo5LOJ+SYk9qKGM7Wt7hrIKA12AMPuB5kV+vNpbjVPhUcmut9yzJtZWeSrZI5dlGwdcoU/UzaCZ
+sOv/GhJsNBM3eHG0UmOfGYibBYKr6+LdJbqFhX6S5cBtzuL5NhsTNDVwMUswmpzXPFVetV/WSJA
kssJUPIlrq6RPnSF8JkJ70zUhTK+OcZc9UiR2ZvoAQ+U4Phnj/zWd8v/PpP6eFcSHNBFJg8a9nPc
UPjftD2VmX+pr6EsF9dF1no2PHxgTqNGnd6ZSyg3jsZJWxV7Z1Hoc1+N8U3hfS+gBkEeEmS6E+2M
oXt7B3D7qvWde5QryzfHM/v5npsFfdo7+7hz6/z/TSK4QKDwM5CH31ecJfHMEMvoERnHrzxdSDZM
FMlZw+YGjwrzCWf+4QHefFpPq/UJo0eX2RyuW2Vmx7jqcG3bBLriAThIUPQ/hGzQVSfFgknDoyC4
G2rTPy41iXR1O11FVacB5qpXlilh3Iqtxwj1Tc1hC13vL5IvvvCRERiGE1d/TG/Eh1rJOvIqpL3p
nQVAgJNEk5BHylXwzzsjjej0/UqsJbxvY4R9a/NdLtvYzSMAadetDFNt+8ILSnE7b5ZIuUWvMpIz
wc6iBnFF8CyFhvF7lzLEwmrlAXxNEq4VRFFf9DXflhYRPHwd18C/7ARaNhrvJlTu0g/nuc0A8fwc
FzsQV63vCMvKN3Ny7ORhcMsYmDcSodZTm56COYpvS43cBYxnlWdNFiEqmuH4Xp+Et7rEi2oF48Jl
VqGctIjmaUB1yfHvQy7GKhCsL/ImAjAKA3HJc1x9RoavBcuy4N5QGeU+yt5gcJy/Q2H15+lzUUIj
XwqyBI9NqRGfZhKb7YWhPnwIYjU3UGif95+Xy2ys4+XYb73hgNjm4hSdK6dlfB9Tluk/dgX6TTe1
Skp3V31VGcjzHs6Iz64bqfaWDSx2g4tqnfPMFFHHIqqrYx1eM786zmI3Qe3rxXcDi1hFSepaFhpH
5Si06S6VmQRur8bo9IkLYvY8GI5uA+0zTc0VnUwwArGBL72VjglT31BkHU7IPQyFjmxeVarDm8V0
tn1/ca+kvP8UlPQXeUmprzu2SfzMqqSt0x1K9tdGN24iUxoiEqM2wG0Vy4/NQdDUN4xA+XRMhC8W
u8Qkk5d5tmx3q+CaNEsZ0YFd7UyS77k99RuLmNz3dFTRItraHgg0Zxr5Z8wL45JbpM10k0YCmLXj
hk0b0H9ST/7viEVAhMIigPMrRS8XGpb6Wsjc8PJY9INnHu3ZMyfj7mKG+UjI/YYf7C7l9gMYA6K+
2K/0ZK1j3dD6cuCwMvOzTfsrEd/C+F1uq/OVmHhHrzWMaaT92BqGrmhjFj0qjGKpyH2CwGLQy7fe
M0UmtISfwFX1isgXrS8Vi5IeFLDAGCvUUVVx9tc13DbgtW89+o8uO+isGmLFe/QrCjD6FHZ9E8Vb
mknSNmmyTD89M3EmBwGjbOsNFjJb5++HDPtFqvxrf6PlQtIRvOcYYIth70P/1oyZjcSICgw4OCN2
MZmncH5sv76Eg3kMceH8zkjfW2DxOUdBtDnuP5znHzpZOehdsFEiBM/QWyrurDVlhUJigcAbjpUX
334Afyo2C6iD7d7R/DZcVUJxi91IesRBvaIQEdQqx0UNPy/+oH3Jwrj8R2gBhRh9LMb/0JFUnmEV
k8j+gVqPus022GOBeddcGXWhtDlPjD3r+ay0KQ2lRPT6khmXu+2MhNADdaGJ/F9Y4VBIqH/kVKu7
BmDaRjQx89MHJO4e6l6a5p3mukfPAal4qtsmwjIAmkibaF/VAjDPq2xXzcBZnQKsCegiH8ovmoNT
g+i+t7fmE3OS/8jw1GKveYBrMtm5QkZMITQB4EmwfaKNiETthVCJy9jmE+Eb5Hfxts9TRdEhCI7k
s4+W8WW93eNUK8CHGJi16ClTxLOoOdilWbdHC4t0TrRd7ytUKpRR6Ed0hlM8lFMJ8qNfFZl3vXIO
Sj5KvZ8vM3DlXzfmKOcgn468vddXvwHkf/OebdvuK+o5xZlu964P0P9le8AeaQx+GvoiNAoIZK8y
Knq2t8SQD6MLoQj/I0kAX0trpY9vK1zd8G7kXQINfARlRr7CGHagroPmQhv3kDWL8PmVPhZMW1+H
YD9grKt8jdl8QIz+yUDXVbWz9nUsTARzHagvKcJuoAELZlHrMa/uIAGQ3Xpc3aCgm7/4L+xQOypq
BVsUqjFHCj4z6jc4GCv/GTz3mCUrLOz2vuryC6zCyS1SG/ZcfnSOnnLxk0IxrkpHCfJkZbTxX8K3
/Zvu6I5DWJEm9hFDEHQHk1x+R4QFf5/Vl0IuhXs6m45aZ7m2NpvIUViqjbHowNPD5no838V/tgKE
l3Lqv7y2e0SksWReXMVYsC8oc0niTxZgXJAvqJB7ghRjimA1nL+kmZjS+rezCTxhO0xrJw9rnixO
mLuBf+150P75bF2vTiZocNHl/EhtAE7fWFsHt2npUdhgNzc2NvN6a0jPx3gF1TobJzfVaPRSP4EM
YAc56TIaYA9pqkf9gJ8dgiZb+kXVlREoeXp9AQgiel/nHalJTcrbVyEowFP02UX8B9M8VWpfbLZQ
A3lIdWO9blEhqLqfDVGsZUlwYEaZX20PT4AamGXsVD1+t+MQ9q5Lak8X5Cbr7ecZlioabzeaTIaC
OScYvOX/ctOPaqXX7w/XOZseGT7297PfrMT/GX8QEIpwGi54lHfPCWp3EgQ7rydl2x5XrjQLEyC9
1gG0YHwdERv4n3SQM4UYDA3g/doojWf2xy2v7J5L9OENo6MxQDTIlKVgYararcLFdohQeR+z1DG1
WtZ/CJkJBHwJoZR3JKrAAvIAlYi7RJSWE5NK5fsjbUPSHvApN0//7iRo54il0UjJrMXjbvVOzjgq
d8aen14N5jpi+1boQ76qDzI5d6RAlTdgP4SUuTiO7REIrdLQ9W3XPP+zOgYLy6e+SkAzf0Efa+z0
Ee+fqWyN4YeQrGq93BX1v0NZ1DWKq10cBUUxP+lhoqkBsbxesZNR6cIli0N3qeGWyTe512UeRd4x
zAyzeQlfvfxmko5sAm8P4Ca4MzwoGm4YfxtNMuRpgC0qIrZ9/+8LZ16KKrQmup0CSiw3u0X5XeBN
OvMOv7192xylBC3M7S9YbpnXLm6TLd8DkVfpX/Q1jiO8m4B+iXB9ofd9ix31cFy8CI215fyrKOM+
eS/GMBCZ7zLw2Fm45IjbNCAaNoOxByNPuCOLq5Oa5MYZdB3P2kqRfAWQ2ZXgiBB1CQgiV2sP6lRo
Pi1ZSDHzhCngfAvWSxHczbHAAOM5CZPCYq5KUW40fN5AvxPG3/vw1JHWN8hrYPyOWAfHVKQVKKPY
ScJbPae952bMIcY0EOwGgqMuR8+4TQD5UVCeGbEEg509npUw6SB8CUcxVceLviI3eEfj+FnId5G4
V3qyC17DmojmJffNwbzXS0ukZf99BAqo2BkMx4oRto/mDJpFkl0mkzZ1q5058nbGUDBosuHNjNll
x2h9JkRF6mjpIiIFr7Wm4MRHC46L3OZt5vgwAto4gXrZ0JFlS2qO2JBqyQvolrAVfBrBwVQHFeDQ
rO6Tqgim2lmgtIdDsn/0BVuXXjwExc/3/2bfbq78IWKY0PRUhhG0aACIApHtaJm5jggM3cNXO9J5
dwNuu1RieVDqMMEP70dooe5Cop9S5gGXseqn6FsI51Mp4Aun+NLxjtWJ7DD5srIPeg2B1MIfkQ0I
q3xdfVup9Jq2CTyt/Gt3wyWjjOhiItUGlstmmrsu3Kmcus/D5foqAdZpVtbVLXvrXNuTkLmtkted
w2lxxKbb5UyN5hT0DSXIR4mAn7SV8u1hHXp1UIvWTrV8+/yZmXxj426BCnQrLzQDsnGEUdqL29vN
MyVVg/vIkDmYSXQrTtA90R30YGHNcIvPTmerRcvmQbetwmimsS2nsD7RjSHwbxfvEie0RCVGGvy3
mv0ALwQXUeONEheR7U0iA+tvSj+a2uw1bQYq9Og1KMGtWqn041ZQPcmpBsQpnRN4VH1XiO1EKGII
yWvNpnf1bkCOJeg8Ve6USvVDairtesT57Yef/CE8rF6wKy/zalwqDih4FK4UCZwmtkB0bW50mYin
32j2rGoCl1gmSu8MPbOg1PRbn4Vmx2ITYeC1K4QGem6xDoJ1IgO03VJJOPvXaVfGN8cvLgDigUcK
/0ayx/DR7lNUTddLy/dz20S5GXfWpJQ4DYovMZI+iuUWinn6Ui8QPZ1ogEWDLlQh2rIU0tiOkO12
AGu5OyTGgI0z/hMqulLUsIZQ8BWg6FHD+XPcgrP2Z7P9/umVwyTqnsDoCLpevKWEjoh6InbLKG0I
MkVEeuh/OR8w6mtVuUdEf6XnVqvxgUvylvPv5WUu/JLs2MMx8sIodXl66dUUAKJlpAAvgdHZlrr1
vlMlr4PFgyupLlqjL5AbXjyjDGgrQJG1/vWuJGXK5NuKEAD/ZLlAVEZ1d6ZhoVMiX7wIwlbRcnIz
0PevxvmHJrXoHHy0ox3xqBVccEt4XFakxP9lAThtyCShPT0/pqxzGj/aMSjYMqCnH+TjpznON/Vn
Q2EMGvwJ2PJItrnFDHbxSzq48IZNTXNhir8lRTCPMF+KBQ3tsSQQpouWtu6rminXa7jxgf8bph7w
2mgiSD0iFzXag8Gy90JNuyhsIWoBhwSkp9tiyzQajkJUJHi3anNnVEsnJT6apnVZazMI9hJkKlud
8bmDfCcObmXVLBcgXHxa21aGWDEY34jI1DHbHuRXy9KOZCzStH3Ox1KabNDGMruwZIhtEZEvhlOu
s0CYYb4S8EeHd+vWjuJpd8MN7Ay4r5QNQX9ytkWVrkey5j7fAkh6rFWEw6KBz7dazWzqzqU+Fzj4
nkoMfU7E3W+64SV4rCrVr2I+is4uByEfeH23HY986TVSxyIngb5FGCy7FC+o1+wZM1D1JT8XtlhQ
y7/roE0//zhlMSCuAm7z7OT9+cUgJdb0yHYgGTD1ARG1CKKniEkkFEL+Zs8IeZkNeWVP2BbvupB1
030Q/qjf8/iY/UvhknuvSj8vqoNGFxlXZ+NQ1CgfjCtmCbNbcJ5DvDwndTcCwrxCA/k+BZk4/8Lu
btxzQNP7Kutv8xWo6TzBjQKFKUT/ebLfIbqx8MVCAiUzusuMJ/52KqRIZhhG0X2zaxcCP0vyjzbd
0PgAYMxqgdRFZBa3mkS5h+I4zCAX4AV5dCylKYDDZ7USuguIiLv4nsprKxOtXXdFGko8ltU/T2c7
rGazjnmno+Kb+dXJ+jn1/I69Y8hj8Hm6ILQVjpAiJJVmuGsGPM/tsdy079H1/IoClvAcyLczR/fn
+kjt3S9qZ7fUyJwLGFaZYi0GHEz9CL8UXHTK/5m+xHaZx2mKkMX3WOzBprC1y0V1L6zZBYmsk5rl
4UG7b/zqJkXAG8pdV+yzU1Mmw/1lz30X/kjkaoxEA23v0qxWZbiOY53MTYJKg8Vd82Z7NlC7MAbA
b9XqwVy1b4cLmHmYM8nFCmCo5U/d4FEDo6B5z/MSZa4gjoh27r4QRMz42buoxdOzaVSAkLzPM88A
/takleA1bZVjllDZorkYs15RT20hysSTSyTUf+iZf4h9hdrMCNg0cbwBF/RO/rewDqPG6lISP4YP
h3N2IqAwNP1rSAU/3rM/RoenB48L6/qmpPYSRyTLujmNHvqSI6Bk7QSzClI//o2Uklw1TQBl/jM3
mVbsURHvqzPkveGeShx19SYTM8kt+ZX9csn6aHQaatxSAqkW5Nr5ZZJ+E1f2tuSbZAcu+aZsKh+e
nS5F2xdcLjO3x4v2iKMiIe7014LmnPhIUWX/7/AlJaQs+5IMcmrolgFc8u2rtYP4gERb61nRSgr6
8J/1Grx+9ZBY4ctl2jnIAN/yjN8rZQqcx76rr+aLLSItg7KI9B/fcJiGf8zmstipLO5jGDZFVo55
mRiR0xoTeDCorZWxNxPCvsQrAai1Q6nKqeZevgBZCxrQ+lQEuwoNKmgxgwmFNwA5lb5zYCwVg+yw
EmqopjCjy9Aiyzh+JiWcZECVqNLHYqI0tVRU813cDx0HEStyKfmbIkd3tvBgm/9GWp8cEjZjkVPk
OzvNy803lw1ddKyVymJjZ8zYyk6TZSQX7x1x2jcD4KQfUl4ZhMin5oHwQM3FbLnyh5GMuYVu1GRA
M27v3qGZs07OeX1Da+u3nFOkVx/2IWVJrcY8nYSlS9U6IA+KhAPAk6DYxiJNHYrHECXZztompL9P
3TMNYVYV+fL8PMxKuG2tg+Neh+em1LBQY3P5Byj/54WP5Lot7NaNJn/joLhTWLKVq8LV/EDEPteK
GAhkkSUnYDG8vosPmVR9KVcI2Wb7NBr2+JcqwDQODWLNT6HQpk0uKYFImdYslwXyyOV8KtFOhR5I
C3/MFXuhm20nzAysY6I1G+87Z25UHlbdV+sfeaUXpRQwojdy8Cfw/wIdbaxCI4sCoG/b/VaTr4mj
xHqUjFTcSxt1TTKv5ynnYTgJnD3m3YWM7hgAng0YYJB4m72eEEkjzMhwsIuPOhxaSctYrFBCYFl+
yzWOuOp5mxyluO6dt/MBa1Np+3hqsfc2Zmsg3pELDMBm1L3spve6WaXg/n2VPJija7y/1vLvWGQ6
tFF6csKGPofitDreS+0CxlIu/t0akq7Zd2/Y7RNBDxOgJK1qiFNUixOxSy3KikPxlBfi+CmupGXV
7Ri4cS2HxPGm77hFAXZqrdMmHXjkqT1hqHCBZ9X76dtF47cA7fXygBehoCBTRgZ4FbDvGhKMP7E2
l/BP3iSXdKMSI2KLj/Z1Ifg/0fNeejxmCUqraGl91/LBqTcL+6Gx2QhX/KoMRpbPqbbmQmKhCWkS
Z6atjnW8E2B1ZlzRcNyyog+zdlh8oy8lz6qUToVhrH+W+tJOF07d2m75R3pnV7CjbAbXtEn8w/+W
zC9hiU1g27MgwyuTa7nlSTJqlKmdI4p+2xmtWubImzKYeW2tf/sDOArSSIWKEXKbE7be/UPZMevq
eRUQZ+TBfrhcxGtFCmjggzQOazorkibtxwxAM3ZddxN46PtSU7MjlReIsL3KWn3fIWELMqnGRLuO
d1i7gyweTkmF9HNQV5PMICZQEd+hfqdVKjS/PUPLWWlhdQuKXfpT+E0X71CoSh42f09di8EY0P2g
BmI00xd/MjK3TUCjUvOcrtEO5uZWzpaPUnIGC5zZAv8KC0xhaKLDHWGVBVX9jdH+g0Mv/TTHRLoN
HU7IvWall9L/r8OzuOPu3J1/U4UvffsmIZP0rncEITKAtcSapzEp8ToL5NBLk3VGzq8maYVT+LWp
QZVQKcsl+9BJ+th2Ff8oeyW9lbrooGauHC6o8dujrFNVsE9upQ08S5XwkrcVbw/KEI6oDR7hN1yi
02KhQS4Zyr/oHge1NETGfjkZwHJ64aH1GBTBpLcUuMIJm9dBPaDRLZPIfNzGgOei3kvAbh0jOHkn
IzoUhIJzuakJuRXV/YDYjLRyiqWHT4Wmm07x9cAB4bpOvDTjDFDjc3u7ksHHM2UxXXXkbj6l8hTA
uder/uCacqtxY+ZEcyKEWmPKG7KrasRIdKCT8Qps5rbVusSGm2FY18kXx3DIRiT5MVZncav+GOgl
ZXl6FaULfjvW+7VTJKsqXErZmEOGFg43aOnpmIZbO+NukltFnC44Qi5MhoA34AGkmONMdH31eGvG
fh4qLqyYi8eLrwzq/Hux9EC3rWhW51JWhfhAOH/vvcTqz1Si5hMV6sDWRFmRYHZnNgz+k588nZpk
gxehIOwbA7baku9ZHITPs56M/GVLYQfbCmryIQCfZQkxK3uiTHDenhFRdrEFbRpkuWn6+vdRO8Ru
d34WMw2sFnusCgMoKMpdfv0FzwfpzNvU42Dwi1z2iWkm34bqqF3C2iCPDCJo2mqzyvqTQtP0g6Cm
WbjY1f5OWRoy2h6ONK5LRH0P+svehLPXQNGjVVUpT8ti4xIvbdY9uOIf/9XRyiUf9JwTSo+ebhl0
XWB/t8jhTu1WN1ChCnPHo+FlVrLMtYYcxE6QkBOvKOgCEQDKOAr6AUh9Nw98g9gKC1ZEBeOJcZZX
fWO5Go5qX2OePn8PFjJUGkUJi3CDe0NlscdI9G68FK1RYC5hO6EkcE2D8TvBTtUn/TeYrHY8SrhK
ldxfj6JYw8VepRO+2SNQ3aV4ktSCa61iBqXUrkUV2H/8qSWVyBnt8tX7B3nOYekV+rs0O8/Tf+uK
eocD4kbq83cUbpWsNu0nlDDQKJh0y+ehQS5JVPjO0bYP21CkXiy8TpNeb8nz1gwKA3TcAimZhIu3
RaIvnCwGKwmPIpu3OvVidF9ipVkalhijLybYeYBIpQAQ6LVFpSFixJwmEVxaiLNWSSL2dQ+ROK7P
/BpffoRKaHPMbN5/qLchCM6Au3GU8f8jK1PFxmQ6Z2SDjiv5Rv9sjt/Q8IvRLtXzZHW9WCFW6Nah
VJJH9mGXQ2sqFJcQAyEWg3oog0WjK4k/R7YRj1j7fR7qB6g/4UVJ12lDO0LZB3W+rzoQ7G1KIZKo
5XoDa1g1s3jMdHy7c62xU44udRxk5zeDJ1m+1pR/e1wzYqQDfR7fXKBDUM7wLEWcruIt3f8p/7bQ
sZeIIB1UzTLVCWDpUJwTQO7XJRyBiX2isBS947wHR+0CGMzQ3lOd8AtMi46zxqY1T0EvW5rLike1
rywReBfHiu0ozENZUry3eEeDIk1hE/QFJEvu8ESHJ2AhiBEv331AXUWaNliUx2G+ARt7+9l3Q/pb
L0786kuq6GqLgd3aEEHxzRvV1wqwkLlDMTG/oYds9wzj/E4pLOjU2Yo8bPyt2ewxngGTqTrw6mM6
eZ44V5CPz/ufLPDsqBPQka3in34zixyUxQA52cr32YduU6GSP7n65yP8adKTYcSS/6W9DbVwuGBh
VUKmJidUj0DEum+7HeX22G+xbOk4LWBFzIfUTexEaOF3Ifp2Px6tnJlCFdIZl0qqqpPWkwZy+8g4
GH0wwRj3jaasQuEuddyi/Lxso+7fHBCPCDlTXRBkvbQyIS1leHv56cQAV393LwnQc1GX+2D+Bzny
Ixz7TR6zjowe2VOgIjFT42/1l6YdB5MkTli7FI1KL0+ywDgop7kPV+juAg94YH4FFkaA+/CjprtC
+T8izmrTlaH9vrYHRyDFoMO8yDjrJx5b+DuSfuKAHDJvOjJSlead8mk+6T+p+blQfhwmM1jfY4u6
XU0ZRRondHDd5YJAAGq34MzISdj08VSpVwFv4TdUlwdcMT75xo40lkmt+45ILHHkhs/OR99FqQqP
FnW66mX2zJbe2etKppgmEC6aH/oKBu0mjugyzL8pkh9klVce4qy/AAPPkiZPFtYY7Me/Jb/zeHoO
syeKz15LsFqEh0syH0sROXQwd6qSUVHDT+TMwpDzk+o27EaFW5153pQI4xa4c+rB7geQo0EYUhmd
BJ+Wsj/UvQTPGAOmBjiO3n38YBjqW8YOb/l8Wigv+U30jWSEaYSIR0knYmRBoUV/zG1N8i2l/prO
Ucw8Ll2GxA73vdzXzr2XmihrP+SN56m9yx4goPzVQfXW1s8xha0BH+fVCuUAxpYh0bMOih5yF/cC
70cIeXx2Nd00Yf8WAzxyquzX7ygF7Wno51UmOlfRlD/t5xy17I6Qq8EywnntWi1U3tCCMUyYYolY
B8wUfv0TPwxdTGKK6fD/NAw0qg3CwmcaS7d9pOz29UYP6Nn5pwuH2iAvU1eXRpP3/lD1tmkDS/i9
51UNwQzXI4AJvY/lHtlJmBx6Gw1kV34l2GRKYpx8SciPLZdB2R2T0v1EMIFe9uOhYnW2QZt1n08R
fBJIQTkxU9+y9+SrxFtW7IxRRbYcDlofQrq2inv3spWRlynIDz3VwAac2hIRYUsvCHwOB0WPzlLT
XWB6S5UU28CQQA3HwB4qbkQA9UwMg/BQZlCB2SEH26bmBUuERFL6+aC10LpflXbg3pz6shms1c53
MgEQaNJJkR9w1qK94mdQdQSEe+sEtOizvGoVgG1qdpzJdGx7IFQ5CnGV7ddWfcsNQvNwgqLBZpb3
q6XxEoyKkaXxnPD0HPAOoJtKUUrDZBU2lp3MIQrDojNyVFRyz20iZpKN0TNsHFEHLBGLNHxonXWx
IbXXLy3sS0LTp1+ROzlEeGSpxogIq9ovVy2ZLitIhHp3Dp0bWeAwQbDN3vU40Q8t5vSENyNj8cOF
DWkvia0JuIc18t+35BV2oJTAYuhmgJphcFTZyQEYAxpN0dEDNjeY8OjMEvRcRm+ZDLXLL6Ghz4TU
/7AQ+BRpS2sK4unJGLq5EU1CGRmTTokfBRdT9XVuXCh3BgRobAfR4VExKlc4cn7ZJAIrUd2Zv2m/
qcQPAqtKiBqHvMIK2QEZEopckPfSe/FHG5Z32DlwdQFipF+RFC8ZvkYi/vp9z7l0YHaxizwryLYG
WSXXodVXYwYYuGo8x7fNxHi8fSOGyJ53zTbxijdHT5VY4y3wDKBgkWkU5DtO+zt/0UrTk9HBN7/O
hvSqfBcRRt8Zx60V30jGk8bJgXV1LtYQ3RVcbrzZo5or+6UkIKfKzbRa5j5+xlrJq8M11IzWvma3
B8Lar/XYfVhgs0ZpkUQ8YeRRp48yez+FWw86oujkWz/fhQViiKzAVZliJtiJ8ilz/mAAIsJdsDUT
mXHs5JjwhrB/QnfY8NzA22DEAKSZAmtuOMvNr2X05bmdq6j38YnErDBAQ03SdQ0K90VcBIpL0Ss0
6xuC38k03LxlgiJeLycySbtBUjk0vw9WWniXp4zEUeMm6GH6wnhSaRSpkM0z27nVCECMpyrUWlX+
Qh1JYkLrd969WOlkT6RaqjR8bo2NJe1s2mYdVHdTA3ti5d3/T3szu6A7hiN2+j3mXkbCzhyTuOkJ
viOhrRGXBF7QbOxAfW/F3V3iguuxZgSBPyWv7zf7+Y4BnPFaeldIsfQG/2qJ45QouYVFjlatIP4e
d96aGxf/Ez1/pIJaw1Qg/zTo7qltobjfChYqzL0IFMqHjbXIKckRgrYfokZ/eSbXtJq2G3CFqNLI
rqS5ABo3QENJIB36y4y2TPp69LRjMo4FTwekQq3P5WKi70/c7H2pDmoY+kLzHz7n34nLBeZkqyiY
GEeebv1eEA99ICgzI8jgM2DtGnw6BmyBTijL/W12v9O7vEknVbqYFukXzTaV7SQJeL471cajfNo7
x9V6+KZ9E0KC8TYLlMU9/iBkZvvg/hL/b+j3PNygXHnnbT0lJN0cxLcAjpXaBK83b4hD8F37XSn1
KYIGQvl4Id5HT4mUoxYbCzCSpgBhgMULZDW9N7nPACMklRW6jWR/0q3HyiHRWLhoclQqJW54D1g4
Tvlh07cG+ob1cx+8ODsO7f2zoo5v86x4kPNxGz6emAOTXW0i2DZsrEXlEJblsLHWhTjH/F/2gPOk
QWP7SOAc1//i+CGZjOA14IjWYv58OGBEeKZPcMpAVGeGkq49kc1kGFrbdlHSyUQTO3Rg9TBc2kEZ
HAaE5ZawAgh7r0zza4EsjQhCh8OYEumTmcHyQmUnmG+FdFegXfNhA6qDWrqjITSuIqnbe85JLBar
hidcZcfVUrIrmh007rmPTRiq/S+xPwJP/7dk39qMD/XwHco2C8eqVS/KAQnk3yu4UD6xP+eUi8RG
vrx+W+wXqaHsZeW90da/ioTQR2WO3RXa7s83NCal9+YHFDptO2TnEtLYxQifshHacn5IEf0YviWQ
cMAI1FsTEqwiunajSFo1Lbz59Orkxl+GP1cKq0iAsOh4CbPXbcx3DrtajgwWyJonFAszA4coMpMp
5P7lw8CnqWQdViWweEcc9EMyMOx4BOxnKJ8nJO3Y4sNjKoizsWsxoT6xSUYdhAuYS+uTrDWoW8Ba
2GeEeKnYOQsfgIZpQmwOzM8DhrILrrAb6iRT7yycpzGsJwAbZqGJ2oBeZIt32G/2FuAjLVXIAmgQ
Ra46nweS//SmzcsqY6LZ90VsK8+5g0b9pohQTXZ3fKKoON7dtbs0uFxJzUgNld2AvlBypfr1wH7h
uZDwXRVYKew/RKGRdMxn8j2kINrQ1+pivbjGYj/PJ2mjy02Ie1ECnXYuYuiQYKKiO9Gt2gInaLkZ
LJt/AjU4J6fQTrxL+2/AHYSr8ytcio4PnzhoNmnY6hgcn5cJ4dJoD2NamwKpi+C4/04nF8muOeXw
P7Ds1cfeo8PJI5UQhEa0biF5JgGqldO8cg8LS3gv1Gkm/Mb3Sqa7+pdi9zKKFnifnJkl1uLlVlq1
70qUuaxaC9XZoifMbBYeqKO092MW9/Je5Ogaawo75vnupJ2nyVYgoMUNL7e+DM8jMda1dMvkXsaA
vAheX3LQhg/wsoVzijHp11CKgIZ++Q1jqnf5zknYrlx06CHWtQenyrDQQdkK/WDn3qqoxtyeJcss
LhsPIWFaQCogIZUxEjgSiHLUEp2rMcMta6zSuHEMe78Ow+uz+IGm9lfOunsMo27y7l3V97Vs4qRf
ErSvqyZEuKvpC7AeTCmThC5GJejVWFxRVkJqDSDs6D0zLYs4LZ1NIweDOfK5B5LY8ShZomP1PctS
8aPVe9zlOfEMMlGyL/AiMRbo6FZeClDx2xlHnBxTX4NNRarA7iBozaHFQDP8FooMgccCSdONDFmC
nG1RxUv5XOyszo8dKf1ah2G15DrozvC9rM5RLngIG1nd40UMCLyu6G5SmNU0GSA3guFFjoxf3J9D
yYOG1rHoy32JDOWI8wjJkba41bddHa5DVcGk+kYCLxFQvOkktfDtsv0LM07qQpYWm7fQvKIoaOic
mlUN+rU4L9jUwX4FWpyx6ejYLn1/2+nwY/YZKwyTpVvtVbWgjpHDQKucHtlu2LmfZrbETa8E/SH/
lSAuAvkvoC/u8FpVZ5+Ieb7tdFalxdlyVaaomg4ATkDF8AgA0rNko3NKaPpEpnBCZ1eugziST/SJ
GyO9skSUO/BWtq16LBByaiMzrDNoVoFErtn3u10u72hOCtdU0wr1yQvfZRrWucp4cttkBpH6NuVZ
X6EmLCbEg8M3NHwa+UlMWSzIm/Q8kpRSpmaHmKxUMsTFguQQx2xjhfV5AXJjsLeQs/hEJ9MMbJe+
XGLmrr7WlZi6rmquPR1Dh9Y+zkK2pRg8dYxf6HIdFBeE8MhFokK/uYQ7Nay0PDl4lY/NbkcTDLDZ
O7VUF5VH9N+eRScRNy1Ig/CQ/x7xjeHqZ3KP8ZNN+oQSeFgmZluRXaIVoYvUbN+XN1LYRq6dovJ9
zP9zVBsnE0o62awf1GCiRFFZmMkB0Zk4eHmkZxjElEKWosSze59+aO6SeEgLgIdsXqVvvNU7/6l2
XgsXQUeywwwvhDOn4sU8CLBiqdkD3SeZoCnhCRkFKHrefrbwODBQVIveoZOBMe23DKRYFhkdW8KE
tgubNDYIfHTPgP6dIHXGCS56SruLWsDglrdRsZGtr7rtdr4l5hYRyOe5xxgGCc6kggaIpRfpHswS
AodhblhFavy4izu8chDWREWU3IULQkONO+DOU3Znzls19WXcvcbr5dGzSRIbl3KuJeDTR2sBRYwH
cvnNe+O9wiHsWBjqeRaSQ/BohzPyNDgrqv+yfQRYOp186hpdxpCbC0Vb+JBa1qmL8QeHsJMe97i8
JaGzKxOIdx0uFY5pRtvYYIGd6CTaL+1AOqybUZgwHS+7V8q4S5ORjXHwCmGc3KVVv3qGd2wCunXW
xrY3zUn9vyIx0Sp9q5rL4+l+RIi0N3vfErV65KxrqF7InBjQAq54fP0ZhS6m/Q5u6WHYYziVLsyi
dwJ+bdapcxnhjZowW/V6iobXmuj9O8oXDzdj8ui0U2CZ21CWTre/3G4nGqfVpRsP2UIpIGP6C4zy
y+aoHfUPqL5+xOJ0bRFsWkyLRGaBtt+psUtUS7/ThlAsNlr2JQ0zXAiRowBsARYruGP/QXTG/H/G
rY2O9x++xJjqCSfoLiFSdsHeirFiSX/U55/nHG0OF1X2iaaMYeTi12vjsp4yNyVuIeTs0gtXinuD
PvrLWLSuWG5yLg195GU8L/4+r6iUwUWUiCk2LgD45P35FEr8NlFaHiy5AjLTrko9PJSkRx+dCPQu
MOOgdtdr6FWtHLeQXZ8paOsD8UaKLEGdF3MO0LXLvKFHi0B9WjAyaCipInrgTmzFmr/sKYgxj5WA
eH/lubhmmbzS+6WVeWAAaao6W6UOE3+wl3Ym/WPlcXHpgnQ2AevsPYIJI/xDtfAeV4Od02f8YMV2
6FsttWuc2QdCl0bVk1oSqvndAotRnZEa2yu13LT4c/1yJceL7240VjEFAv7kow+irCqSIzbAavTE
gbfxaJSDb4sJrgRyVXcdLWCBBAergO8jJ0y3eBVh+4HaTK28vT0erv7a93pNhxRSNhCQp8tMKHPc
W2zODk1qWohKHjujbvmzgG2dSNl2D+LlYP2GlnraO96Ku3pha0yYN38CgA0RSctJuBW1lzNd7FAX
BF+MBeD6+2MLYmN0AVLBR48Zde/WW23pT9F2ejLf2Q1p60j8B+Hm9hlja8/I0Oum5vq5M3BotyOx
MOIl9A+u1J+Sh9G3lH5CM315LaKvd7ViI7ttbDQWgEKgpqTxTpG+yyoE3sUUkIALiJHbnNFcF8RY
ozDNp7yipmYjHHBorEIZOS2le7phOjARCgXcBahNvL2k1DjO0yjiSvwWhixlvRX51naY87QTE3Av
4NGW4GXW2xMgAEihc6ejcltIEI7LkpBq+mxQ9lVBQtrS2qj0BW7eUHPUIl4iv1viBSmD5K3kG8P5
fux+w3SEaiflSLi4O1WDh5j5bXIuBYo91b3MMmZfmA5Bs7/SpE/faRAWH+UOEoIByPNp7q+fKMtK
Zd0bs1FVTnEvFGbjzRp6eGfZ+zEXp76tKZwZi6k1NTCBtBDqyFX3X1Tj3GY7VHpBey9Y9uLmHZyC
DzYjROhOxLw+Oi/t36swF80kxs2Sm4+hgOGTC0zgoKbI+HhWatEX79h4XmfPfebPi6uhyTadfUkZ
3Nl8/hRAnr4Udiini8bhg7L+zoiAxnOJtZYqDDvmoAAkDB++ZxJF85XOCy1BuVxpMQsvGae7eT9i
Pyd1vwdS6VGFxJHbqnM/7Vhgts88WvewlBXd0NttNcYCUSiEFVqXy7Oe/PUflHwQHueHKKRvgRjV
9hTAmlPd3JeE4VT/iqQxVC01d23c40HQVrG02mzwyf2VGw+dIbzQVjqVZi6czEy90sE9RejNdmyP
9pmPqMjDc/zvlnUjmnnt4VTDai5J7bEkmVFPis3txk032LhlZmKn7VX06HooE8cWb5Eg7lFm1zpb
80AS1TFrBoITFkiSj2qOcsGmHAzlF3y5I0JIxIhhj05TGVjjhCK1/t1q/zRaADFSxYM61UBU8RXD
9CrVNUFbIUZinTLIZ3yFBKyyNK8ynXPE2vCkktJgr92fvduomc68vRuOZW3PfaM+QflWjhwKYHOT
MFek7Nb5wR+0+OdAblG0BoR/+OGw8HVMTLp9W+WMt3CbjQdg8w7VxdKfDMZNQGU4OZeqeeTQiINA
0VsIrKij4ITdcGX60DflG/P5W8J7qlO4zTSTAeJnnWswMbVf6ai/kxlqAHuwxDoliXPxY4FlMte0
FXYGRka2SlKSwsdWFG1v5yIkYfhDTyn3R0sUScZt67OHo2wD7Y4eGFP2t4D4oxUn99ACxgEPNCHA
Jo90r+119EUtWxiuD0aJJj6ZQNwbT81aVUgSTyM3F6SaPLSg1rVl8T6EZ5okgnY3YtezSMH71W9M
yBvTRR86j0lgVTCAg/47v1Qnl3nc+hkhhEzUrHgilO5n9LbApPjJLXmtxskdQ3GlzqDkTxS8q3OC
y41Gfaj+6KXXW9W60HZyiUMF+fDymLlGVe8xhJ2Il9BEQKW9VrjIdOtEI5/uWvLwXMSqlimSBo7h
I/kDZgkkArvYvCUGs/xm4iRPWa6NLLk5uY7sUtujqZ+OyXsbDQseeVJVI+9KJ5HocABMlYI8fMDL
AV6oNwSL5ke2c3Of3xM4tpQA/OrSuPkZcUXSQ+pQlr9VRnEjulC5UxHER14lZxPLlti1BUzwMXNY
du+zaX1/8rF71zZqrJ1T7Qc+gt81lbwnlzmo1Er5HpBsapDPtags6elP6lZZFTv/E0Bx9ywHULD6
zo3SmMLuWEXnfo+bNrxwCE27TdMfjjEq6t393wFAzYaj+/uOZcLtWtxUUI9TtFM4VIhWyPDjj8F3
locpj8gyDDqGsu8CVBHB+wesCpUmCg+cjOhbK3yNuehd1zPFByiVTKLLLoGvnSxktpI7uScLbCs0
rywmdCIKxJpwaMlVOB4ESrcGmBWiEmLsx337UsY41cp+Hs+jqKbbFy91ohBpaLWsgn68RwopmWWz
xP6TWPjXAwP4C1RsoMD1RggWE+qzR0A0y0PvyRXx3yRS98Nka3rgl7hUh/4qmeKV5QcdDlkbWq/4
xk5BcKOxd/P1SNt0CYojwKrQCO9Wa/XB9fCTyN8ci+T/vD3HVOEIue68S9QWa/0DfC38BnUW9Xnb
XWLPWTAHf0YUX+uVNquf5lWTzTr9AF53tM63DUDvJu9oVm/JuAObQDTyESaVwv0fPeS1aukDtoy+
3kn1uL1+A5ax6J3lifs7vz62MEalRqDBDr2CPVUDf5z6HAtaNiZd75210Bj7TbfR94Z03S9BDyYF
qs/4HXtusf94sRX6f6FVZM1z5zRibAZT0CJjAJ1FbHrUnwejec9cCtzrpYasndxLXnssfxyM/4yj
RmotGfscCh94pjccc5OdPRtYm1cfss2xmuFII9pQJY9DPimnqFUHufQq2Xlk/s3VKBLHZ2UqZ4ok
gJIYYJ7zB9e9jzAqh9ydXFvuW2/cTJw9u3dylIP6ibiFw0KPtHowLq0oxxIZlTRzP9bCI5LSdT+T
3qADPBHrzcN+Y54awaM7C8kTaDPKnWzMLiJs3VxuQCIkpCi9sxhikdY7efVpn43anGOw2L7VoeQJ
puoCLaUYelpsBw/16MMN5X8FTF9qntRxwQ/ZBTJ5suiefuXQI1kB3UeGxCXi1XFNZ6HRGM3AdSHY
GksEHz9NU0yl4+7Vvg9A3PMsCAbODXen1xUlgdtQZD6L5UIVLcv8u1Ef3PS5ZmBOwxi6ig5xfbD5
dCcM9doxmgKaPDVmsb04xfvp+oBcQrxt3OjLnAwqJHrAtSroZlPVnIb5g4KyAKT5k4X8+BSXmcYD
BdzWrut0zimU2Neb7P8ZoeSMt2QEfJCNMALh20gYXHpf/ja+I+NUbDFletFuALN0jm6p/dWrjKrY
xE/N77J4swiJypiyH3rC/bLp2D0JjteYEClCod0mHJ4alZ3flmS0A7gUdD5gDlcMyIxiH6/uVkCG
bm9XA8HYEHmkws7f/FLfP14dfCDgaVOjleV1Dh6Oyw2CYbMbmsnrkPPFfeqX8IlsMQHVmryX/5SY
1e9wgAPwkChnpBR2NScnQflvOfj+QWYMTrYMcxRX/CQYNtPSNqmT3HDCKHEsAqH8vsnIcuiYHX8y
u1jRR8DNYE0lxGSKiAQnYvWeFgKI7oQD748SnivFEid61/UWKvYe6jwTLMXk5xLMlecx2hQBdM/Y
m+IQI46md10L7dxuUdj/GZnH6k7cuXNLkvCA8CzNkZEi9SyhyraAbf5SSCZVRFuHAYdDbwaHK11z
1rFCBTy6z/MbA1bwBLQkxIq/+pZRUIA8+KHIooYJMuffQGCIMh0ysfqhdelamsF3jWCGblK47cVP
xEKLh3CsofIF4K4auB7f3pEyW4T5rsecRSskQyeQF4EQRqJKVOtmZjgWCO30MeYSs/PFRJDvHM7N
J4r6hZhUZqs2TPb+8mD7datL5dqyCJO1thsS0eBDg17gdq3WB7mbfCxTej0AEkMWwNb0kWme3pBC
vrlp17pijrdJCef9PuPQIqalNePsWDdap21ZYN/nNT1DW1Q6KSuz41ltshRsUn+arumtPG1WJEIH
4HcimSi/l7mTcqGnCVTyY9Z8egbk02NBuqswa3i+sb60ZUPdnr2BZlCm4zHSsJB6vapSc8uO3Zkm
2985bVQkPGMyQ+0o4Rw/Ejoib1zFrVulBFO+cOnNh7AjRFTTLMv3T9jF7z2BN0ZleDrPYXBVkwh3
4Z7lUwVVteuEnV5YSXoOF9iwMRy5itBHpoQ+zRBhqHRdzRPxpycx8rhM6tqvFXVUnzEU1hN9NTax
/K16mXmO4lnHoTHBinpRKpgw7k814ASHeeoiIoMs8Paw3BGwy/v4RoJgzuLw+Gmjr/DffA/TqcO1
gslRYl7dCXdNvnuGIRX5oZyBysV3X7CjvAxHFesf6C+P6P/lNNsUwk1p82uIilqorJ2HbZuwEo9M
bVf5P4bQpzcyh0JWeQqLE/F9sgtHm2jv5PToxrKICdLjc+B9bW/X1d6SB0EZpuSkE/r4rrCK21lO
F9DsIG50OOnoj3ayf+EAkLbJBp//B/oiFN+dHz9vSHPh+5zGjc5M7mvEnpHUuzw2QAlp5/nkELdz
FnnZ7uVnFOXI4KbfGMU1fWkmjiuIFtB3yR+qzJURecjBAIii1eNY9eNoy0bKfFl+BV2e7yYR3x6Y
g06xPB8ak243v/kiPtToO+xNFM59UDF0nqzNTf8ml/PRQkVHos7C9tn136nMzk7gRXcEvC18gv0S
hlw2pbmgA77/wL5axl4Uvm9QhrKVPZPp5Vp+DjVeOWWZ5hjX/yO+5lQLR+eSxAY1AkydD+Ccblc4
745/f5kRo35laaROgYvlpYNGade09waRJtjxxckXVKN0/Zc9TjEcZ3js90MDOA6euSS2rvauH6d8
wjzYlpZOqccQvOMeCXuArrQnonrK2pA4qxUi1HI5d2WHhFonGPiD+GgpSHFZzStJuMm6J4/KzC6O
zTeXVIdye2pTeH5OBNhZYE5rmX1AyjXYE6NbKvbbeSt9o97lAdfLlT9J3GWKAvYg+n8xhoGe5Nij
NzM6CF9ST3j3X8CI80m38oc72EftU+RvifW6D2sRg0yCzqPmSO99BlCUPtYK9vRHiCDQtnxQoTsQ
EVevkUlMAQuE9TIkuLx6JjWm65kOgrft/Q01M8XUrttZ3S1WshMMrvsbVBVKqiXiaDoWwDwFZN4e
UEQENRqDmnTjtoOjFpFVrmSMsrIKTZbtTEYngALpN+c53Zu4w9k5DLPgUAJ0HR6YtYbb8Q87cNFt
TbaDCeS73Knjlc8RxE3p/VBCTzcAYrxc/NKdbUeC5+dHvX2vrIpEhJPTK7Vkbk5SE1qXLgSQuh/N
w7OjDXADnFUtlSfoJzjgPzfj1FtM69a3C75QEkMkGkHAosIX5SvwUOQKX5dhy9w4UCxWGceyXAth
dYT3/ReC8+Wjaz4YtXMCZpIx4B0xBJXgZ7WqszBCteL7hPolbz4XOSlZLUt/4HvFlaCPEyqOm4Ko
fdDojKXsWvdseES1qi6oPm+X7U9bxK3KUW914cpQkwy+gSU8Hob2oXh+buxGE5Ee+4JR4R3XZQhb
LRYfATCF/1otfZ3YYdzzAzn+2BDY97qlsv7urvpjS5LyPSCRP9DerdjDC+8tlJiFaL2k1PGiMicd
xtBySHcN9Ca/tmf+K/IZBITxHsz4CBFx86VdOoEN4oLhfOJDjSNA5kP0mgsr4HawPW1oI/Rb++7d
L10aRGjSwT6eE2Q+4anPqxtI7P6wOaAKHsn3OCb3lozrlK8Gg9bNYlN8okKotMvkyuIrTtxuh2j8
8WGbjSqZF5UShSqvShzQnMz1iQ7SxKx8iO9g1hm7fcPSqMIjPXspshhN
`pragma protect end_protected
