// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ViiXdNVOSHdQ40gHOqf3s5kvNmBzXZjAmWbm0sSWPOc0Wf/toTUIOYRkYHQHlKPKTKNyAXBoJ0Zm
dD5S5d3GKothg6/sSYF64LSkVeUaOgF35KPGXUUjTIDxTvJClSL5i5/YvnMu5iT5X4QWBbN6QS/C
mCAUri9KwJYLzTE6sd3NWP0euQ0bOTyzb62yDNK9SmFgKFagY7tjyTEP+qU0lD1wyGjE0NIBFtpK
baHs+H9ZirAAut7qX8e2GKMZuS/br/Jfb5gYiaXdVM+ia6qwS9VlPLrZfJ4A5OsjfrXfu56ij1g0
TeUouPK200KYUj1u9L9g/RjHswuZ+V5RhmkQVQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
vS6FWQkEoN2ko4dD00pWCxrfutvqGrPmt/vScNI3UWSV/488mqmOF45YS8oktBgLvZ5aEdBgAXmX
gFbRuvb+VGpYVjrSvEq9VgexvGLOclEH5ECVd16mWSYjJFhrUncPYTANnWi9WOphcXEEU53v3oTV
Z/NBHK4TonFZfactvHKDorQAfIFcRNTOlHvLMm1LvwYkSACopoZAk5Ox4wfAac4w1zoKC8GDRtzg
vqWMMoWNAobYCvrNGiqAXEciDw7M5ft12RfGdRWOVMPRiz8aOH5FmCaDegTR6DlaYEPhnFx1VK09
YjkXT5OPsrv1WxJvs/Ye8sQ+fVLEt2l2id4LOT1D3dvw+bGZqgjSYRnwri2ER88w7cAwX6sC0AOK
8O8whqCxtdLIUEeNJFe34Id1S94ew8Fuq/x4m6Ul+IRig/TT4Uoa/ma/eh0QeQX3alvB+LXBle2J
1tJ5CWcKLVbNujUWaKs4OmL9Ixp5ecMPi8HOc4QgfOQDgY8JEGJzmk+6MLnn7yuypBRvDnIoLTdH
SLjn4XUloRTDkQ4yCxlhmrupfhCKio2kEPN4PakeWVTOtFXv3vum2Mfrb5aYHHdlr4YSWdHluGuL
02VFnCDB3Cusx6ANoNAEZ9wIvBnaVkhkmA2x/pfInqYyM7gHFUO0TdC5kHvYNr+Apt12MmSBp9sW
cwtUhM7Op1G/+yv0uCNDVPrEmmmMI+nBGQmI9EcTs0sRR7wNDxxjlaPRxxIoaGFrYexjMGSZdXV4
HCqn/eWlDyCGzcgpmdBCgjuf9bShH0heFSIbwvgwDdGYduXIWxzmiK61z48lZw8d/6Brw2VROQM9
wLvJGkUVQ6Gsa3St+fICzaW9uh0EFbb2s7T/E+dhoRP6gv81j3hGC8ceGlUzGr6boiQiXr0ElXbz
KFnrQGUTgPf/d+ieGOx9r30xGUklUmzQRBHpfL8R9C/48zvLgPbpAQ4U2jCtK7aqkQ+zfk4gQzlf
9VNAz1ZM76GawFxyNd+JlD3DrutTIHpx6lEl3DrHrEwugQ06RQO8MxDGqRShVdgC0hwaVIa7XtQd
32ekZev87dfFF+junPGYTTVnemd9YaqUuazsqrXQsARR1cTbj3sbk21+FWjiHMnJYqEc2D/hc/ze
t1ubStJxH7iWaG2R4tN/piwHmWcCZG01GDJ9+/EHHbE01yCsolx37eHBKBQ2MN1UxssHKd2A+xBg
BGURrRMqBooRQlVJ8MKuz3sPHweVayEOLh44rDJJsiTzCocBmENbT6jXjyWRVyaCSAjl6v44rYjt
7rflf33WNUrITInpNM9bjE8fkZxzgiIKIvq5Oiu+9c0IkBW70uKDecfINyW3/9s4AG9jEzxdt0xy
TveTgiABBEGHGm94XJ5vwl3mE7U6Yztz03TQqcOtuNyoUDddv801iWEp2eakWXzyTwVlSlrvjNe1
ZVUmvOBuXirkli3eYSAdqOa8v6oS6njJVBiVmJlYmi74+CyAmNyVIqqtp4Z7CjFnqgsiLStN0PWc
H+10N1yRpOSQIK5B0yw8vKg1CoB9qI5/Xg4btUlWmYZs307W62+BFaxO2W4Wod/XR2uPlmQe9dk3
1/pDozGX3+DfDvg8HibfXMuzqP/9Q+N2Ie6Ic2EDes4kU1H95f6VvVNOSCcQuQRZPIafIytmj8xK
XjPY1HZi+eFOSTscZnIX7z3BWVWhAR0v5APIq4Hji5NFFqDJ92YZLV3idqwfnwpD+0CkPhPEcFxU
e1J5SQHo4KEWfOXCb2y3+gxOWpdurR93rSkY9ytZJQISeZ8ZKGhizawxkdBbV6GL/vSamJv3Efsq
wu4O9zDPSwNgvrms4y+HCo/qBy70tNBgIQ5MFdpxtI712hSNGRXZkV2XRD1Mn1BmUgiSn9e6p3gy
dGWWnIjuzPf6vaWMY7GaRrsKvJcz6xEaIfHGyOw3UBEueCA1463Uch40aYGAXhpG0Crg/pTaTr9M
QZAb0QeRVvhFYrYZR5avrEaZTI0X9ClpXzOMRkAOqm3bLrdiG2/uAN/TMsiDsw/FAWzXn4WLskqk
SBzPKxOOh9OqFMzJf+fBk4djRJdE8wqcVFE+j61YWhUU7mRELPVqlprvhJ21E1Mra4DohEeDbMT2
OwBb4dasxcni7rPTKCWGzI6s3CH8Czrh1qQ4YR3qxDy9IanGa46pJUi10dUg1Cc0rBPaEdJFme1M
S7vuiuDuEziqKjZeKneAc0f6XFLKTrGVK1xnV1+sX8uIaG1j1zHLs9ZlkCGbTyzMaks9iYN43Hru
ybsMq7cMGOTKVrqJoQAhxXsiIaid8jaeLFs2sKKonqGyRAAFYQWJtuZnc6fT9Jc4Za+HxMI5r0Mr
F9rvycJLod6IqKbeF1aS8wI0m/D6wfDrCkPIqIXu/toGLfXDJXkX4PYrEXySjIliBRVJQHQbsCXN
ap88A8VhZHFhAnNLXVEbwwrBeG+dK/mCjVPTeeh0PitfRHB7O5nYnFk8EaPZefxe5wL+RJPEmzzY
Qk4BQkeY6a7+JSn8ghZQj/7cMD08KVN14SwmdH2sPVkw59IFL9ydRj6Lcxuu2qQ1qIeTr/tvOnO4
hfvJT3/8fUa5IwBF35QMkeTzPQBBvRRe1N+zCg6eJ+0kXkRYSeckoHYoGmDdWJoUzAyz3lzlpczm
moIzoWGX04woxNsyMG6JkfZUw4esD9ekJvcdP00DaJN9eMR2vIc9UfV16680rCT3tby2DLS1mW8o
i2XJoOBI0dBC2LyvylLmh3OqTEgkK4HDPPNG+oAE3vJK+WIkY0ioxudosJjcLvnXtfERz70/wQ3m
rz6YCr4KCjTARmNcsp4cjHCNlhk/HrFZ4AT990MU0fxW3fvdo7sYKSnon5PrNs8TfhFbzjK8Dc8O
W7QYvULPYcZe4rbm6im4WWHjZTyrTvX0ief8dR9irRVV/GY8ywFAMkqf0C+FGmgigoV5H8HG7W74
DZDyFp43y7AJQcfZlSHcFqocPxPqBS6eguVRuyP5jlqS627vDFipKzHzGimD9uSxrrZHZsigcOKZ
hubFj/5lyuyU0OorlsfYtylR2HB+cmKkal16S9NohXdBkWEp9sXNPaW4uxSGB1zQ0gnrWmcIu3mH
WF84UHcrKqawoTRuLR7/jJYAxLm3HeV5GwfYcA8f9p/P3bWx5UpLKKsmB6quJwxHwbUcTicU6VsE
fNaadBlC6Hm2+7cxeDIEtToptv5WR3vJTNgv5wYrpa+//xkDIOaFqqWEdFqrOpW1pMkpJnwGiNRa
QLig/t5W94Oet6L6xqeqRuwZEIqbPUz624bjA+Dt+fsy4z7lE6KwGdb8WMkT+AMHik1GzWzWW++Z
WJ4EDLSCJN0U+XCEbE1ILbC06/3LDiangWh7ivhIey35eQdY923RLc87lSI1LvuNKU4x7u/puTJS
yK204668x1zloHNRqh81eocfL80nnyoOOaxWPZW/gjpyaxf6Jw9VTru0C1h/S2hQtvdaq93edsBk
2mqeuYZ0VOoxCPpaVWMdCdxMeiH+hLMkJSvPT1+pMvgtwFJB3aqQO9/sPfKDZjdGxF6lAm52zorm
6yxERzSo5rKy62CNqQwEc349bwJ5rZZ6ZPLSt43tojeAlK21JvPmK6dwZjuuRdSfdRmrFKaogGbW
0Js+ALZIUYOx2T75IzIb9Qj1yt4fuxezYHB9gedwrtPzDkDHLHpDLFlmgJ90IHf1ihu/0LE5ROBf
6OxobW/lPA/oXqrqJIkpfOctszEVCjec3xGMTT81onrUhhfriExcnrW8o7zirZAH1bLDDFQwCsi+
59oFuIs0+2JHhEQny+XO08aOMruPNeApkUwgqOM6h6B2u+fh9vODJ/TNm6mhGZy3NuQz9bqQVDnS
p1xe2OOsM41JOJlBcgzHSl1kWwCwootonsuJBeTcF2iOI7/FBO9CHNC9JGZyG/En2dNwUgAAzzPQ
PDhRMtLMBi2fTb+2GIVo2cnMLla9fORcftmr5h75009eZ5kG+DwjnEk1NeyKW8ed8G5RJT27ypzG
FengoAGJiUTZ717jUW66RalE4XEK6pBbKGS6z11NrCBYbkUIriG52MfOVbbQo1cOBPvDRV4VRD/M
nMLaj9b6EFpyCSkmxH3eiuZA2JufFKmHYk+b8aU2tO+c/YlXC1Mtom0GsyDZx8wxxDGRUYm+QEKU
Rg1pBujHrPwLPDiHwXVwNy8h/+g8R1Vjvc3hyjYTaVSkDSv7DpdhA3MW424Qy5Ga0h7J2cK5mXWP
KrUhnzGovw6Ajilwi/7bLWlI3hvaINEJdfMDvAjID1/bEAEtY/xWtO1nMLTmHNLilCdzrdYriz/e
JVp5S/qX9rvCctB10QW5kwcCZ5Ok9UnVpYMwaa5LbWdqk0b7cAjgTgjsDkJdVaMbGzDE1L53bDWg
3+nwr3f/Oa2vdEE/YGgwrvvsDwTscw4bt1vB6gkSaZUabsMxSZpeQjba2MKL01La7Suq20yeEZ21
Q0MGUpGJUnEzO/fUCV4OMjxHuOiStWWMneAEeFylBIc7BYWhOQ6paCyr4YjP1uACJHGBZJHio+RO
00JpFRGaSiss+t5aq9sJKT0pj3+GqAy7jSseuV4IUZsXjq+GDa7oX2rXCxbfInxqsgl9/DpzB/fs
UzEvUmb7gC7f0WABMf2KiPXu9lJo/TJ6JMKXhzdJZJVOX3HmDeF5Z2Krky9AEMLc369zgJelhEDb
UKDhe3ThOUYzsrmvgRJHywY8OIBpt2w6SZ3fdLtmoDx318jax4/iP+SUulJgMo96dh5ggosTrv8A
4RStS7rlIyOpaHEhsUCMNpEztURof0rTczCMSqcUP13/RUhTIBtyrMJY70s/5+5M/AAE4JwdACNc
5GIPXD9IhvtZGI5CSDY2Kj77SArfVhGKiY1ygD0DvjQ1ujcbzuQ5grQxFqwxvscVEPoEPh+RcjDV
yFmv3EnznV0J2j3bMfp3T67zI2nM6nED4lZvvUAicCO36+dpPUWPObFs7XShuUOypAfKtBMaXfAp
kzD2gr0NHlYfWphK22embE/fTvrYZp9He87S0zbzmfgxk5d0qet4AYydTz6lexAjGwmOIShfeppT
/Zawlqax5TgefGlzB6UjgqN8B/8ZQSUcGwjJWYdmLvuUNdzoADHc0Gq26ljjNpil59VxpMy2EM5M
F4PlZA97A+gBJsFK21KJvjIg3rvvhO1xSXRkzn7N6pktuAE/nrqHUvJNwhO1fbaOykRV9GEEOjnQ
Wmuk1g+8Q/4TPvpzulZhOaObFgq0ZY740HKJwmQTjjt61jsw/tQ5MgHkrW5wOPEFtIxuSrH1s3Rc
MFT1VW6UV2xTMzjJyLCJw+cxYWL11ABNlJW4Qh1rS8cMYr0UuKjh+XkS474HEPUUk6gOAuJj0zdB
l0UP5lXUJNPocah769eAxtTb3Wnbh2ar2gh53t9Lo9114WPF/vY2KVF9D5nbLZvs16ENdcMzGf4X
IoipEVxn5Wcinr55ZJ0rbxqE4ssoc6+peO8GE1Bv94mni+HIp8pN2t5V/W1FBRSv15ZqtrbaCWuE
BhNhN4zGYNaMDVDZPM1Xoyag8PKTQzxPYYYpTquiK9G6rPycAvGi/K7avjfDB+SrAyvsda3uMPyI
+Ynx3cuP879f/IIiN9f2Sj6Ad11JNbiS4/dHIA2FDVngbpeKvLmC24GDBkKyoy+X6KyP+mE2Jafq
N+1w0tSIjPbX3XALm6xH8FtzEB+ZyFuGUob4nY8m/NmgNWDa5hOz5ncPpRR2AQBL7CfECoq3L9GX
/dB79cC9EJ4U1et0dBKHdVh+JkaR/l+OeGd1oYED8IVzCWk0vb3qRTTD7mnP/smtM8buIQP18uXf
73gn/3j2Xl5J21rUYI3au7a6wn2eibNFOHyHlhOPDlE7rp53cQA15mZ81Pbnh9VMq759LV7aB+9G
9luWaIOEKNCvgn02Y4Y5fVo3g4hSI4H29GHsT372/MD/r6RGWD8KZQbHYdpZn/8nYs8aeau7R+7m
DaRFM4GWrrKAxo/vsxxgzLwrwm4ItTZqEA3SjNziRx2Css40YmJLRoOE/f0mYp71fbyQtYORJQio
HUjVqiHGir5vXbVrHoWHo5sNNub6slN307B6HReRNV0iAawbHIUJ+O2WYgiGoETqpcUmEhYJRgmx
ECMTri/zA7Clpgcm0CQvTA5Pgl9O42hNnbFBd0Hq6LOlPdnMc2ZbfuRjt4sy2p5y5Oi7K/Qv3HIg
/7YjximUn+4+77I/wlbYBojwdkOtoCCq0UhGjEsIXMPgqe3gTgdJ84VX9XH+RwMQnz/uMAYUfniv
sbJoNXW5GLq+Drg9XB5Lv5R2W+OiHN7Nzq92YNcRx0FA/s0wIJOWkfvfTCoZRnVeEJgGUNGlmAKG
sdxJ9E7rytPxalvFQBswLAqr92hOic3YQDbZcCqmaO0Q7X2VQWroIKRy0QcHoXyC1Vr4P1WUtizT
o1obqn9KVUa7QMPYpZ2HNXtavyDvMEOPFXGlH+povdfLkWrtD1lizaGdqk2vX1eQFMn1r991KDcA
TUEVQSekeAx+/G/YGC+xTdSvUYkjuWL3ryF/m/3O4JcMJ7RQ+4MJEHhhI/Ew9PB4PEiOyvEOM6eL
kq6LAM57xWMy2lQFhWOaY0GYLp26t7ZiZABnljS/Z84voNaSALLV0oOwX9YnAdvAgYooMbW9hJhr
xALLfBhBiiJ9CgTyR04svRbrQcYmjEVVTNbWCS0wz3rMbyFyqBD1zZ82Mk8U9Hx4okxZixqpoQRP
MWCxAd91Tr67bmamgdd5atXlI5ZcNZogXu9xsfNqLdRxc6CrARWBPIVEifjt0ScN898twQuprqs/
X95Vj445JP/eaxEEBLjCYrmFUEL1RazxfduxPdZZ6A0oR0HdiYcSiovZ/w6+Yw1sPJ/8b8UwFTz+
3DMser4gRSiT6UcO4ITErLq+DfblLfSSUMRCiRgSZ5PrCe1isbM7ar1sXHCIZOqUTQY6CiavbHLX
1uHOciuNIJpzQwHGkJJzC7Ya+1dFyTrMzmR4nsQpvJIyS7msgWBfve1lYbsRBk9mkPRQtRZDMvrE
tfCIAjVYBlB1vy0N3NPdG73AUuIHuuvQglZb2OIzSvB7d2mLfQw0/mzNTUNLGRjV8mM5icAQsUTh
scLPVjZf+aJD+Ag2NetTJdXz8f4NcJWrsUV5uKWYhAhMRy+DAiWv25WJb9G2KqoBUDhFqV3AUYFI
2L+leUCtrzQJit7ekq/tq/c9updl9yvRvV2ZPz6jWc9997lanXjsSRzeryKnvd5K9wsES0YF1lFY
uJPBqXjSoJNjdzsEkzb3eaDWfUins+2/3sgy7ZWWOz9WZKlJpHNN8jpJgGEKtcwzyQ2Fp2Al01Ej
/18RlVnqthwDqPVyLMU+69fLzL7SIlSXO0yrBZFty94fO14IiFrpqlwH97lT1NxEs630n4FV11fY
zMjr0shconG7A2eiVkKiG5h4Or1jzi3bL83y/s6yefvtMX4CT+bTKU6xCbvsYhU3/+r6TB3enmGy
yNJN3y9S0G4PW66AheFCy269wOSiknXzUUDMVZoAGgxVfoE6Rowp5TuVNNKAAMRbx1xEJPZ9OhH4
xaOOZWizd748INmNBpUDIMT339WCqW8zF55bP3HJtOqmjhAylDBadcYKHTPWagHdmVntaVRuhHby
0C1LpfELwQHvTfQO28BK7O2ysCb65qrK1m7qzf2pDsXYDf+1VpvypLhQGTDOFbeIdWyDuDrI5noa
f3xy7Eiy8S8N0o2Db8lUV1oIvVeSn/JGfYrmVe7Ln4K2+5Cq4jIDTJYW86SjM3sBP/HWvwpPSgjP
W3jkgBz8oc4VmqEhtdt9Rnfmwd5+8ixA4qDTogLHOONzOrfvr7PDKu2G0n7gro+vK5ZqfumpzKOL
w6/Y1hrLzzdWdPfa43lyc81+wXat8MwMAjzAQKphaA1LMt44JRw13gpL4VfvDeEo05vKPa977uh6
kQHcjw/k+CglD1GyaXt4fH66YLsZvU98tkYyoDzmW0i6vgpWghOeLTWbCVTS+9xAAQFPvU76YePX
MUFXczEtVTQCDnO54GIPp5zQq0r286Q1f7232S9B6ZDxKIWAqs2Hs+Bf29iIqJcA+wvfio8v+zSi
3I2G6a6xcqFYLV9u6wYBXJDXJN9EdOR43twVa53PQ9o01hF+eEOe6x5JAydeUfkntNIwWPbNOFp3
celRr5/CtWjEhwSCvmYoJ3kqbmj8/LpACGoNHUchsTuhEl+UzBgXca4CnVfq6Dyy6Zcwbt5k6FCF
2aOswK0m/99aW1KKwt/CgmEM224ZOIcNTIz45w5QhYpbsiNH28Yn9KkC4J7zwXnXUV5HOORib7Zy
D4KP3aWk1KuuaiCqB5iTyCv0RICiBnMymLbQhf2qvfZxW5pc5HxLFwUlkSb0NIRTjxILev3ZB+iK
D8Ok6zhr4q673tuaE3/hJdwyYs8bLOM7km6y8hgnw1+sdayRjIrDlpjof693K813w01P8WaoXdeb
t5Z/IKliQPO120XSS6OAG2hLcJzpwW4BIkl8zff66dbVlE74NW4tEKUDBY4EiLF5dqvdcoZEpXyJ
GiEkewAPs2t+AaZ55PeQpF1Tn2uBJkbsw6yt20VTkZiVus8IGOQnPNbd3sikallHVScMhB0F7i98
XH2rDZic427X7CQzfpQc2RBUZX8dLUH/0m2QNPOd2NXy3tLWLHxTUj3rPZFe9nbEFwKDBhTdly2I
YwNHuuzwq7TSsUqV+83wzj7Y2vi+HYIxA2hNBCEstr72oWhNVvpjuNfV2FRmWJzjv8DE0CyfosT+
pREQE5ywC9Rngv3lPCN31y7j8s4CKWLDAEPVjp5Jk0UyWtLm3fSWuWlElqjJtGTVZzrhiRnj0jU4
Nrvq/2E0FmowK/Hb3OMuMFNXW1W9eI3RCvvj9IO+QMLdXRHx/hS4RkQDpS8QEgZ0W76WaiSsRMuA
0WsiSveQTU4eTOhG3xGCtl6O4RD45V1xr7wu4CHFflEwA75oY0qg2T0gYYIu61U/PRFfhip8011x
ohIa7AMMoldk/1sYtOO6TY0Fe444CoqM3ONNK3OF4B8dM0DJiDegd5ojjXTpaYjPqfaX/UolNTd0
E13CfMR2sCDtDdm5oVequmFAW00jZskar2DlIYuTjftGvvZ1bzZkqAn8pzSJQhXkgD7i51dKUKQ6
upNeq7YyDZYJscbYQfTNmdQIhmK1qfWct0VLEVyx96DYuVVRJ4siQY+LhnWkA2pRXSWKR+h3SS5t
Ap7t324BsPkhz4ciZbROEiOngiFSk2yjn9uoLTa6bsUWm301KJDEWP4cAscSYf9RNx9jUYssea0G
WbaBdBFVCsFiADUfhydhklkvS0jG7oo5SlrzSJobkF9SJ3DbaMUOothhR18XokxHWb7CkwrVsKan
OF78cA70B7vXkY8XR2uFy3Jq0WZbfCCONraz8Y1W6LRx9iQ7KLWTwX9rNFfir8RMcUBwgl+Kjv/u
/JoWmd9kM5al24jf+lvLQyDB4kCmoETxxIJKVsGZDgHShn4L31rV+CAid2tDm1AKpzXs3LW+8MP1
K4AokQd0n2BDytXu89US+uF19wDj4pjB5NOximPgSqNGTWxqSS0PACaEVbYe4ogujriqvtvdKpdL
uEUfV0M7k0ORcBxOI84RrhOb8/D7DDtBozACsItj5WwQkjFgUIeav/aUx9DjD+crq0qfcdPEfttc
uJikZS7MQvmBzXIoeIQorjO1A/VMohprpsio8g41p7mdQWTWmGsNKyaezoxMWDJYnbIBCoJGevVI
i0tuWI9/4pNG6f83uo/MtQX3GvpyHN1mAGF2LwakodHiEVTymZpoltTKCBu57ozp+0AIY44OB5v6
ZHypiiE1Pbr2o/k7RkUIj0f63ZsnGoE0RmxafdOFxfmAiOah5LB6XahLvrFIChFDk3Dq3BRicxDd
60GVY0w1jHX2WU9K527gECkpZ7cXZ77nEDcPb3CqwjSKQsfxXKQZaJQ0LhwoE3oZFG14zTJrVp7d
HzMK96XuG8Skkv5OG2JXPrHKAef4huFPopwkgJMDFldrzDRYyTU98lA7X10vIxIkc3rGLSORvXl7
AiAJ08gB4gXxUgtsjtx8ZoGKgR+R/geQM85v0gGIs1XxYNLbPr9VG1EBtMRz0I5z5i9bHpMCW8Mo
6AyqEBvZiBYMGwcCCxtEQwVCDiWSw4m1bMZ6nRVnTZdht8ynfU2EYwXviyPygIDqI3UnGscAB6/c
aRcyDF/kKJhnCLwucDIKhhMz+rKunZ+v97Dmx91zMbOMPREo7esEbbz97DkrlEYSX0GmOkDFDA7o
hJqH/Bx3HjGnzS633phyYalLokQWZ87lbvFBxS8vAdDAJJsKe8Ehudkw9viJGhe+Ri1ag90tlnVn
Fb4TMs+8RhNTCc6iSzX8yWaGLFDeJ7FHqbALpVpe/cdnMKZoDOThRi++3rcn+tG7ILu5Ocv7DceW
bZYrgMLa+i5jNAwPsMkmlAuvUqAX84QTDCVHJq/PoyZU6yF/aYnVmjL0CUo86RIMH92TpR/450h5
XYyJ6jIti/YLeXOawCtpRVgka0ET6zZW4Y0wbNYhidGBRKLIiNacbsQj9pG8P/rc4QZr3EIrk3Ci
j32O1BaMePB/38RIjFzxlhOiUo933agFXZwewhLNMpxDl6DtHUbsQb3/prX90G3naq6+OE5SadpI
MNBhHKVvhF9DkgLCtB5AXSHs8ZY1VTXl6gGUpRzYSlCiifBHzGc5mgc5h2Nz44H48/Dk1ly5y6QH
AkP1pWMCemcZrSlAK8GSm1C5Ft+VSbGOTTcX/lxXhkDfPEeRY1/KmkKbWvEYkTYW/nO2zrU8cTdU
iovXEffwx4kGE8wSylfx3thTNZDYiMEOjS6ysXXN1EeQHPmNlEfepWGaYTao8JPBr2WlB3G0SRgr
IECqwJtxGvjC2p5yTSG1rcoeMY8H13YT2ad22v/8gyJbIdrM8QWoXTUud4lP5qUNfnZ22Rq9Cql4
tj3xJXgtZ1Shh4IgEaO/63xJCu5rz8alTwWXMw614sxBk/oWjxvw2gMBdFSRvqlEsZcPPaaZo/x4
h/jwK30cIL+li8dAyH/ffiQ1pvIBUgU5k2rqPydM5hZHqKnTmhffq0hyzaRfBlxfh/hG+a56aEUQ
1d7OStv673aWwrloZq+AdIsIOfqgPtCwegl93iod/Ymmxh5W2XC1qpSH10Hbs06zEU0AC3Au0HWx
8BQ3rrwoIsDMJzRrD79oeWVe7/5PO61ajhDzd2IZ3yS/0QwxzhUI9E3kU16xlXRDTMVeDv8l9Cc+
24vBxILFRtZn9VLTlzsH/ImayiBZKavo4ZcdrHEHl846BsV0/YnIsp1kdMjlVElVbHytnEByWaG5
KaNZRxPWfD+DKAM7MEzrrWgKxu7CK9Gq4pBW3NuxeZPB7FePSk4noTu2/bRM+PbpitL9VU7ZjET5
Tc8MUD+ie4AZC3ObiuQcgnD63ImcYO595KUx+BPQROzI4XPi6REMtKBnTxf4bxvdOuRb1wc8lCKb
0+Ku+Twcmop/8hurkxlmjORmiSjMLi7yGMPiNsdN74NoXSvxmBM886XsQwfy5tkCu/6IERuY42k8
oMx8dGTyO6eDA3k9uAVJ3tXYyf9kYWTeKYeMG5gDaKVNjthVIamE9LWnfv1aRUrfffbnvcY4aPNc
IoBNgOHnvWm3/vbA96XV3jjCmHXDTST2f3YFheVSvAsq0m4UFugWqcYU+TKOtaA2oQ6aISNjBgz0
n4qsxMYwo1DXb4oLizpAumLPS/FD581JuWTjhxCt28+tRE+3O2JiR5WHZhDpehJZsk42X+B+3x4D
KvzFHEuvTfJwNqM8rH3SVdGrjEzgkVxcwQGcH0gfB5UVKs7NHCZVWsASO8z4Al4pByxG8dEh2D3W
d6lt07I1rPTjkHbMQ74zb8OZQn7d6gx4qQ6KEsxHBjKrs/E32jjx755tfOlEb6Sl9q5RpS7duhAj
wDUS/ZoZBHoJL/a3JSIWdQfUfTA0Kr96bkGPJfsZ91GKc9XwPEJ/vQSYp1f5l1AaVmmyilBwVXql
iChr1H2Kd6HBYXqfzM/clzVzAZAR93JPiC+mcCOlcdJon4ttSJlPvZIgOPSHhPky8RBvwHwAWBjW
/JfLmvPcFaAKg+STm1wdy9VJUlmu9cBWvA9fCGK4Bqcf7Un0MFxdeiacvnMjOoMxjO68gG4aq03Q
A/TViQN41bXmZWF8rbgrhcqdMvDaVkVqySEusS6yrYvcv7J87EKnSjIwXVJr3RvzUeH/tFE8/GG6
LCkhIUEigwbqAjkiw7uR/v7zgW3/WOGSMdT8NYYescC906a1d4he8jKHoymGIg9WKBKt24HSANJg
2Q4+rCOTmYs3Nx3A83AYKusX7wUXvJ7YnKuhRjVH1GkarPbjn7pECSf+8odczqnNFKFIKLYL2UCr
9x4BvuaEOdJASXWAP9Dw11wNMqA6SphQWH3vzG960AHBPnCDxatuiVbZWs2inUfQ/dW6OGJHM9HI
hHVBTLG1nwZRQ4rtvvTGg4wguvTJXSqvMrpiiZZftQYbI84jiJP7/X4GCmFxfVW0s1U8wg4FWPPR
5oKHWlMCRMsnnzr3ncChFJND89KT4TkibJVb9psSESonQBsebZ0e8oIyA5A+NSx4ShAYXF5zxPMh
sE13WNtVBmomil+chtQXbvVG+Y6eQn89sDQdtfwXZ+SVKXqYD8nVepKvYOoAs4MF07jARikweT7h
NR07IwvdEMMR+udIZ0N4YK43QAun1loYxOD6O/YVOmhHhb6sMXJS4brFMyMKHzS9h9yBpYqMc/z0
q5CcBd2O51WgMVAXikc2vyvYco7SaH5pUhFtu6uCnKEmBwHNF4CulT2dkUDqlc4orqtdn5FX8+5k
2MhWAdJ/A1nPKLl9h4U6drRxD0N9GA9HxFzmwBFkO4SKvOhd3kGXchtTv8/unWj1fbE2Xg6s5wkk
O4I5b4CD9pCmFElQ0t469HsfgGiqe+d9/sUCrnNG/jB10hXSxP9uB+qeB9flt14ihp19I2OP/Q2X
aA7jS4tFwAmcjxCeZ8V97/iTbLlmwiy53wzJntUsmd8SPtgSnx0pVk7E6xmFtFupXQiQgh7NEHr5
joQaI2meplZ1FaTDW83WxODs9kTeNVBbhBGHo1Uj5ZuFk3lqECNDGLudvnmzZv9sNXNv4jdHSQd1
HVVw2zwaAKs5f+UYXHtoZxhOHzhqKd0eUenR22PqWY1jdKm0/0xL73vcoKkbibVFCMEIIfqbCAZ3
Nh3qramvawPKs7CpdlVRLsjYqNIvtr04zQnrDEGO411apT6pKaWlWt44/tOJYVjk9PNjoIiwf3SR
hlffnDtvL+jh5/MWw46IF8cc/4/tLUAYYFzqHWXXodemkE4lp49gailxMfaltuhMo8B92SQ6QlFQ
pqrfuk2sNv8YCNiuygky572uffIdVECzu5kBVHze6rxlWm0VRhm1wl9YyiwDwP7FNwICbfL8FpNi
mCls/3jRF3olzYh7MfS8eLL56Tr8oAWWpEXscLQlJbPEWGn/eYPR/1wyIeBfOdC5vJSDtwrFI03c
HKtKicDGou2aMXzxHsKZJErFYdst+lQOoyz4uTjOzjUM/1tHhsJPEC9x/XSQZt22y0ewrf7+FqJn
LFr9akzXOdAgJX6gOn/bqC9xDrMhmPcD5uU8rvkHshMTNqdUH1QO3O+bLVb492MoJ6AuFLWkl9GD
kHDnRRc0H5QuzrdHuuglFWQP5DIyT2eU518YetKxlxx8gyywO0hMqzljFfx+sfjCqwjb4JsAZjAz
aMqAInHXjWg6hwAcYRYVvhTILD1Z3pOMYNRylWJZQcj1yyDrZWCz24m1tUPIY9uh+Q0aWRJiw8+R
zSH9ysVRfCLYzM48I9BR0WNkYKAhCPzfXpUEFit3QprLxduPfbXTJ6f7jKUDlCWkaf8B5z5Ys+Yt
gGfn0MT1Z35Wjroc6Ul+xvFymY1WyrIuNqA7dRBkvYnIok6AkYQjX8qYM5sC1Y7IEKu909Xtvucp
XqElVaGeDYVG1ccpSENclUjzwJiLp0d++XSb7Su+al573lm0Gj9aUfSIFwcpsoF9YPJFZ31SODoh
bkWa3Y8WdABN+1J6ifHAoqNBTB3gaoOhEg5WX/13rU74/mUzlDME86HRnIt89qBlowfHKcGHuvfH
BGrb9zfe0II6PSzds7n1fEJWxtbJewJRyx6FVX4yjPrMpG3IMyeAwZUoku/D4Lz6G62H2WnXIV1M
TouRU8dxm76BdxQ9nb0BALCuEY1fs4/1W5CknXuxwtvKM+lDElTFpeWYBh2z65MaI3IDjlXiURol
NMvV4iTDyL5gqzAwKBVTosIHj72BZyr/rdjydbal1HSAZRO8IwVoWhbVvykcJk9oY0sh/2CYtMbF
qOqaENChv4/vFx1lbFNUANHyFqieKqjtWO9TE/0vcnhZ/F6ST7QZyMN62Y1h7hr+2XBurIWZj4Nt
p1jR+FpbSoEiXsoYhBt5vrdIj3pclgY88LiOntGD+2VQhZprunmdiLv5GzS/6ard9JMkh9ftASAV
0z3R/DpPEXbjyAYlXBX9onzkJtfAR9hiqBQLbUKbMkyIQAloTWDS2zBUW4FDwSdwvf4egNduA1QZ
RT4wKfIPv6EgYgCHZMiMU2Gt4cdlHYy7QQxDUz6Q1vrSb8zrB+Fw09FTy4r0eIXrwSSfMt9Yr1YH
tki4eu/q8g4TzWV3UHkFHY+t7/D6QdvWjdDM5cV2XtppuUjnIkTkGyQtmw/E/YiUMhBB8sRxpWrv
tV9SDynofWA14mfpBfJncUBJvIa5LHOSFPYUQI5ZX3lj1EJLxrtnWHAOru3+RwoeBlbufrXRDVHt
u/UZQnMJZuV2kwTXMAIKcETuDM+HhAG7vgkpLwc+e5o7uOEXDmdPr6Ss4NgKEpp0V3Feod/a2Mll
RTfpPuYgvIzawIJqjWtfvwlYWHVzbBr+v2d9BwHgSWtbg6REJxrj8dpukhCdTpczF8kmL/7B5Bjo
PBRsY7mwu09oqotnlcsUtZTpIrfR7O47aYIRua2DuDCc4GxmSnE8liYn3fH80FHsXGZ++5M5y2+t
Dr40m6UJEZFXCsc1ivZKQaoE9EjyXeTdB1g3zsnki0JFzXFKtkDDVvPyFZC4A+/C6bcLAv+mnZVQ
10i9tChycXGLSCUtq37D0qii411B97olsLxDA34O0Aw3RxmFzKSsRvuUhGY9hBonpCLFLEd71Hp7
bS65DmlfDvHwomIgWW+5jzJzBpgj0MpZ3ykKGGZUiRq2kA4sc6RJz71nfUXqL70uWHRduCdrO9Yu
Dw1uiK6k/SnXsVH1MVvT8aTzH3vFpidLT20ye9UQOyaiM/P47CGlEw/3UaNqN/LodLL8Spu1IpJl
pP3Py+ktyFwNwPt3oRigwS7E7d+UY0DQZ0jBWbrYbX9lu1XNNwhx6IwuK5E6FvDbK64cLvmNMkbA
+XKNv9rWJX1Fk4/RP1zu++bOx6Ns+KOvH+Rz7F9TWaPta9YJyw3T4uvZjB5Z5jaDRyGcKB1Bop4K
WyjWiPnC88UfzWLPQTYQitC/sABkE0AIa/IrKQ0PMkVmb4MF2po4I1sKxvj3/F+YnAzxfTEHqJnz
96OvuNXhfVuYxiBuTCf/Bu+KKG/1fQFRomeZbv0UPTJcMRLBIRkVc8FyH8y3OwlRlNtmf6uKC5XG
qlNLqTl2kkeVSP9LwDbZ4sEbV2A3pfUF8k8UGDZS+lu0K24Ft4wegdJUrboCGxbdqLdcmYFXwcxo
ywBBs5ucxigYp/1V/ooQaaiymnJOUtYMXUqQx3k+apUcERe0JHRuAO1PQ5AToN97rcrzGeMhETgB
R6y6sWMKze0i7tBrBgZmzNRFNKTlM0cQSZ7/Sj6uXPm0+vYIOS3Kh3psjcQpapuWBv4318bX8udg
5weFkHQXwGg7W6zjtTlvALKsJ4BiyCfpN942e2jFMOITQoJDE7HTasqYXjKn+SSbmuI+w2Fg8WFR
S35qxCADk/nnzWwdOkA5gremna6TObkSzaIxTyN2CW1ufMvtVjqh5c/B9vViRud0z7i9B0iEg27Q
HdJP6scBMlyXl4Dm3II0zlm7dBgZyQ1iDGmy9eL5ZrwaWX9vwtJBPIWkhrB2vGeqpHwKBjcKZ4Cw
RY3tlemJwZZSWWMNsBONg7xCDQVIaWY8+Z77qXlNwXdtGX8ND3n3kBPEGZv7an62bfMDcRDxuKzJ
+I7pBhTmaOe6lw0SvzzjyrgO2a1+tAXsz4CMuMPWzeBaOGvMRhpltzQpgtKL2LXaS56W16ShKak5
Tye2waOgXZh7z0tyDWEL2areEU/W6t1GFLStjOde31r2eqAw4cUVjCbkcj4oky44g8ntH/1FwyH5
Bpqxr4oMcao4Sf4hF6/87kjeZZPEki+POZD6QGKNqiNEEaOcxOelAXKktwdQ102ewiEvuGHny1At
t7CPmXgigS2xFYFVFC1gQkbZ3/NYJKAGH2firv6MhNvNVjD3K3U6TgNeSxcwh60wMPymDxwunXns
lUV25SGqLbDsWIxNexidcofYCrxOwYwopAtfHbGdKP8rx+hj0VABlr0CaPo7DZOaG7b9fRzZ0pH9
2jJPie//izOdDIiEjMFVhezrFJAxefc89xQkuHwGY2NhZKqZT6hgnKKHiIo9hIq3JG29ADIzRy1+
n9U7tcBqt43hLjMTIwIEUrt+jPw7jOhdzH/2vHbsxX+ZjPvgPOEQwsjzA0NoR4Bmp9Tk/NrU/oGK
x+TlFviEsmIYbNOXZ+5uyXbmneLzS8CC17cjvYt8sxj5hchcYybsb+qubfKla9/WiGzNgbVsMMPQ
xprXr5DGUicoafHW6eor9x5eZU989JD/9b2ut08DSJu4id2Zhdam/Yn8RYLx4WxLUbacHNpYtvhu
LMhjqSFmf5UetbE7MZYuhL6z5szMJ0r2fllFDDgRiOwe4tI24HftQp5w5wDZQsF+KUx1WEe/Dic6
w1mlg/DV6HzA3vjcDowjJh3xuoPOvrsJ+sVMGBudLKOX/6Kg49qaAzqArzaIUWiQAXD02UORlMOw
Yfwr7tdNUn0W7jLuUfwdFuZrMhsld3MvL2VXAGko2AtXtRRlngsAxkOmC+ZLJ6PZoJ2IL2XjDOjk
P063Mia1wtZqA/n97GTNUWxAIzlNBYQ17OayrRqpgYusyvq5KFbYGXEXRuSUJhjsNCA4mZNcEesB
NwAFyXcphVN1q9Zl69FZY3io+tprrYgQFS8yBPSeze9ED6Fy+qNXS/LaLi8XSaHWWVhwy1ANQ50l
fXVl2eOFbf2VNQxxXOg0W7301P7PvPGn0QEKcvMcBy7Db648jRJzGh8bKUL9YScakMlH96B0Mhnj
FS9xxjMduKTDa5XRTOjyumNk/sYD06+mAL6cXAP2KpiopVvYKzjiUXTqMyD4uvBzFRPZVnuUpM6h
aq2L/39NU80VFn4yKHa4xSUV3V+8bz9AQ/Di7/wm+nGQHJA82vSmiIB7xOHqJra7jD7rWQnfa6LF
6Q+VcaLQb5A7CZpDzNy8pOuxgfCsv0Paf0omyaKpucqbB0zyppZlVJ0vJpdXVuwP4FAt8/rlS4yV
WFbEdg1Gczv4RXMpQO0472MXKjMu0kw99a4zTYOm+sK6zlunB9Mk4ogvVhU2RiWHZKHZQEM3pLRO
ojKtC2yo8ivYymcitMB9EMtaVIvTCdy0OdXwEbY7E5GVPd1meOu1Hk4Xeg9NVymo+yxdavDEmkxt
jkeRJNzFZCJfQv7TaYHrlSCmBKTYnieYF3zarH9t6ls2GS53JhlXymLi/byjZL5XntulKwcKF5n+
CLW3nQeOB/4ARWhuVtXQUx0j8YoJyglXyObrZietCrvKWxtXbjL/3J9aynJFUKDoX+/FMP+A5AEs
kEs/0ClUKI8RpR1ti253POW3FPzZua/klNkGqVzcpIEIkhjoF0f+mvral9sci43DdwU3Xpuz4C2S
gqdq7pyhZdVhzxC0ebiDign2EG0MJy8toqSXWpWFPRq2YXxiP3R0QxF2im/+qni5vAqN6tC95sVc
KLoGtz4Cj5U35NzWMgwTl2U2Mxz64meuoJlObiTxLc9g/ZvuseUrcesozya7ZLH81EOMULSaG23k
kyEPzjVXcDQdtfOJvRbOFvA88OjyuJHt81CQSfkLrGbVbhfendwqDmcSHJKP7LO50FZMBxyybP53
eboZHR4GtgXOG1FBHKrQqIiDZjYAq2CY6eNsKPF3e5SNDknRzR4SQwPPq3NjBTzLIdG49ew2zrEB
mCK5U8jYrbTQGCgzOtxa3LSIQgXU2NGENwCDh5sKF/TCKxsbj0bETrCzY/e1hBIL35DocnWI5LZQ
xCnQc04etUOm7saGP59M+9Ps6pBBVWhfBjmhWDVaeWva9auZYHE6aXyfC5XhEwJsBBnXnAdY4+zv
0WNJ4CS7c5MiR/cK6ZSTH+0kz+9qG3rLWqQvDjahD5f7rQGxK3RVPfMt9FPcP3HY79CHyNAtdCre
jGWLVd1Uv7CC7JLeSy58IrZyh+ZyUp7I/hJDtLmZ3o1tRK37VQ4Dwexvd1nTsr3BuGeNfUis+qHX
x071Cyw4VUHjsHSO4LxM3fxf4c0zX/Ey7xWiaQ98SgEcQm/3GYBAQ7ju0GNVS9p8Nn3AD48o72b6
Ue9NjdOLqTEkCunua2LkoIV34uJ4AVVeEW6aNqsuHYt4PVHYRE2MmtyIj3IVyXBZpoZQFeQ+yl8L
Xc9CCD+qACSFXNTdDUSD3x1se8LQxxNtLhzNyeAuo2dmxVlr2+3EawSV0Q1m2nZ9KYKPZrO44Ivy
MAyQ8WUzh8yLbpQvxlbzBLFoZb3MesSLS8ToxJYMFY5GkyKxNUlI5W5zxGBLQniDj0smoxyxiQRw
4KlBlFFwlzLxCtZeeP8eWoqk/526v7qPsc/GlEVgWMp2ZCzLCYcqzt2F325aAIhyJzyMS0/l489z
V8Avh6BDKpWRLmgOC8fVJMZE/4IUJI0wzNXONwwoALSNKWKL1M66eqFFbWT6cPgwYQk5vP8PehWB
0EIHVUQGNusQYGZuSEKpe157oqAPWqOAuyL+ET/XCTqEfAPt5vG6tjXpFDbCCMMOh+bMsEgELZuF
c9Pe6riubzO88hkPbOB3AmFF0pvW6eV/WzObSdhiapw3t6vxR1MFu96TW/QHXJjI0tTa7KB6VLg2
vDOvPW/hMcgYBOvCN3h3LW3ma5vqEBC+Q/wvl4gGRgSFPQ3c119A5vxtU2i+YDjGyv9leN6ozRdH
1oy9W/3oAa2oDJigqdDRdsxdj4r0j25rx2o6MGNBJgcujw+3/a5xv73kOODV3+FBP/ac5DCuGWjh
RGN6hEDHVyvpRqWzQoMH1ABa9UDcFdvlxC6FMJtKkHdn8pE6HFEMhTbEgBC5S32ECkLD6aTUDXTz
/G3+08mFtrh9yfzsEjA3ymFaXLQ1wVwxDJm7dfGP1l62MsGA7Vf0t7flro+hVL7DeIv+/hyINDR+
oe49NrAjOuUB13CjooITZIaQMCXgzQivN0cvBNpCdAgbKSwZdtdztX7FKqqcaGkAWXR6DhR8WhF0
VZ+8WjI6xX/czY52odNxTkZQ8LOuj/hnV6owIocwojp976kQpmzXVQM9Y3SSetao3+3KzBQWsdZa
6OzYYX12DkTPPbLRzsmy2ZOEzGh5IpO8soteItb5Yk+3rKKaBW375rEelIhSrwByuw8NAwjn3IbO
ICGE7/itFle9f29QPQUztMjuf2wYMCz07xDrMBdQs/9Wcl6k2D0as6Ob9K5RGJfIt0cbf1tx970/
+1ywwWZNZyvgA637ArgQ3u4gmbJeoGCXlQ6xDih+o+Bb9Qj2WYoG6MFSiB0QbzehNIhKIhRrqUPK
1DzwFY9C9QtWkIeFKRPdU6MBOtHJO5vhGGi9LPk0rGjHIbZ5nis3VcMjcWw/nXx13NpBntWMbV5m
JHUKmPxc17dKmdPCvSS72smfm1G8OnVv3brs9J8vL79PAprFvZQN2y1QeiEuvTRVcyC6niZTOqOG
wpytR2R1R63M5m1NsGn8X9UV+bL+F6TGIQlB7UZ36T+SVzKcQUAFLeSG/eA7t3+OABkhcvLA5bzN
/EjvWdAAZSFRvKX+NxVu61Wea6KMXNzQERFk79XMqKPIfYzwKFpddJs2WgxNNey60F8A3WCNKdVj
UXMGgfXcr511d21n8We2H0QBolmlj+7OZi/NavKmnpGfvJMFtz7tPD7V6SKnx8YhhamHDZAYWMjE
lZDoTNeRrJCFPLrrQUUKRAwU4+AShpmmM54zH9iwRg54JNpG4E6HJsMUMIS/yw7BaYcjBjduORjw
a1SuYWlDMfAN/nPWD0PtKZNWiXScdky8ufCGZwQOL2ol1kTw1c0zILESk3ag+dzHSB216o6ATeSK
kEO17wGoXn/6+7ptuOBudi+a8gaX6yetvYYQ82CJg5e62ukJANIoZvGroPf4KPX7iFu3CmrBYrYI
XY6JZlUzHfT06BVreIHEG3TA9wCeaheIThZ/z57hRGF5/jKNJLSDqXoUJbb4MAAW2nPzEvZcqUNh
y8WsbUVTNcA25eHhqMIvmn+sUvOH2Ob8bjmZtd6JBmBgQrfU8K4ddL5iGIOgo+82uca63OyOy7w4
qY744OPHcT/18PWpW2dRqUbr6q/W9f70qzX1r6XpYODxT9mgp+gU3Wa1PT7h3mJl0G9FsmOmv4Ts
7Nfz4HjVh74grQO0/kFaZn/iuZDPwm7pUJ4vYXepYEowteqnGVSAJ52RKSNKVU3Ordg1Qx0mMWA2
PlaDY+v0C05jydDeW+f69iMkEV2wYg89lBrsVkAip82jOmYHpGFeie3An/JLmhgJSzf/8kfNhSTi
Ir8VwQFy8ngxEvPgjNpjAOrltQgqg+GNiWxTjxjK7RB9CiRFtEmu92a2fb/9jRwcXpjg5YxEPwgc
JuhwXGpmxBMDxk0sFdhgm5NEHSO0mZ11q//32jzna5RlD0XpHBKPjW+WCBX/9jHM5olJ6fPctczx
C1jBb6MJlzQE2fyZg4pQQ1rbO8/1vHGS2a8gyXY6otL893wWt2Y2otftJtTNWcCHHywuDD1Rp5/k
v0wfP4acjXzgU2qjsb2xFBD/R7DRWMRBLQsm8Af9qoyDGAWqbEpGZg7LeqytkV9ez25nALRvXbeM
bTcNGOayvvCCWyxUdU5f85ejeGjXxsK86c1Dm/P6Rvg9WkIwpTexZtNr5F80717kU074eLkpd4PC
v9sfigyhIA9XcRKkRA+xte+RVnmaDMM6inEYH3V7NL45ronEFm0IA1NwX+pE/d3FO6WfAO4kxH/o
kDT4RRFR8rmhD1lS8vOd5PbzYRoXL5eOEDpgkJIeYIHiCuSkuaJkpfygGGpc9zMFShG6WdeFV3j0
CuZRpecxGFX+2EJYwsQ3GV4En/E+6v3Q0Yo1tziJp9D5XbJMW9gF+TNJfOAy0pRMCkqLUgdEAs4f
hBQvCQOEeldnBSl3KxeeG7sTx57n0oNMv5T/gpqFQotmVmNxhDvZb+pXlvH/pE/ucBPWTrhWGgy5
wZSqLJulRi3S+znMPbFXJGIaJc+NDpc9Cs3uR+bnmqHb18jazUimC6tk54W194iMU6cIaDfohL2a
xrF2RqIv7nvwoN7+rjpv2og4dHU87meD7rfrr/H0w6ohj9AJmZK8JHrRwjSTyzChzUjRefEtTGBy
PD30+9HIt9lcqzLNZjrDMqG2bAaebZ+v2tNnJxP1fRaaL2tMtEaY6Kyiqye3WqBlJ3pHihJM8fYG
J9B2LT5kPCv0/fHfhVmxb+pPMkMWjgQce9tCLszFkYFqN2iXVdqu87NI3EMiAufuHicctpJbJchI
90zd+ZlQq3QPFunFQJryYPYyFexSJ2NbDtv63psjerkGETXzWZfqB0EmKX2MePK738CnqlGWhOLQ
xs36OKOhLZogredvE3K9e4EtA4+ldQl+hHBYtutIauqSURGp/qU/PjRIemZMszazreuW9vZZKN4X
YqGlFhaGbvMHWhLslcllYpJBzlVRznfkJkq1r3D0VUj5RNvR6M6KDfs53p1vRHlvk6PL6lXCJydP
JOyORvzXh937iiEcNE0W8QrF/pCULJ+CXtSXLzoYxnHf1gYcEe/fMXaXeexbZZOlNtPN8eaC/+Ls
VQUMwNYFl9jIAiMXoMuSDzey495WYPbXqCBDgpFO2jlxZm2wlaMiP4GrNY21A9UJKjvkGU15sJtd
1tO5QJB/X6YHG3ta7uWYgiFMIvc+pzjCf1x1OccLSrZK36NYMeoZbTNOGOnzi1tFoFwreKHSco06
2UfK77PayoJ2IRV7eGIlo2W14uzp6H34LNr6eIU0wrJWx1SHY+gZpHQkyU7HXXecQPocUM1Jrk8P
Ack1cuknqXvY11KZDPwux08h7PGWTqWC9nvdHHwDLCCqrPyyGaIp2ZsfhwamRv4CgfGWj7rZ9ra1
ll+jyeDLNYSdciGbGcltlaZPMZkeYH5gqjUotGs0j2Fuhrnx6SzBsEIrniV6UjF3bTCuR9yDQqyP
NsmBtT1RyLHsyjTiPPkcCHjYhkfaUhY8q3NJQKFqGzoPXSaf2Ud/7S8QS9ip5YO2laXqgwuiNUNh
Y/exUytDxEDggz6lkPJpnz78LBE7ge++RBv4akqgXJI7zs+T35THbxXNG1V+HhBEkKRJKMrbgCzF
LrFIU+mpStYVy/9hgUUFd8tZZ0vACnAzenzmGq/8BxEBIgdSLIa3X/XszsDSMjHxg6JWCCS6a8AT
V8yAhl1o4yWFNwDJyHgjN4z1Q7DU6LyLcK0V60MoA8iIwzkvYEipSUj0pQyg5itVSqLIeyLV1DNy
ATG8V9+7fNUJ7XbpUyW0LaqAPsL8uKuT1j7BLDp7cdAxwb0/ZOHrPZ9R5fH0m0CZcyyz35AZcf1B
LWgQdZDaLxwpG6qnwhIYdwBEMXQJqq8R3MfkN4fzQO3PsZLngJxABBpYKHDozqdNwdhwEV2hQqJo
RQL4UxkcaoDcFslmK8S4rFZqPX1G9KlvSDlTVG4StmJ43vPs+B7BpZ0dcPeqMxmVIyC+LWMieW26
d0VgnS6Zmk+xcWcwgcTsW+F+Esy/YOE+S2nJkTIFENRJMDz5E6TiVee5///IT/v4IIKPufwN/nqr
i8ZUF4okqBUbpAiG1PXXSIdSR6xYIF3fC8K/3kXZIUUVevf6rDMIHSt46f8B0OHCDojYgHNHX2Vk
QhMZiCH4N5ArIl9ZN7y/RRy3Sohze+zNhIV137NrrP90T8Dq76LWq2d5IBwWCCYV+3jWo6V/TnNI
9M/lCD76eBi6/g7wd6Fn4oAO3v98JRy6+DQkcsGJ9cLvsTbXsTba1uvV1cw4uqHMm+DFcoZXnsW+
SwE0vq5CPKp/9528zmrHmS/pSWPycmU0P2wGBKAuC+6SvHqYONNFN4KNQZu5+iTB85e79sYbrkDy
1SV7Q9xmx4Vj14p8JWQNxHIKuNbWBMFNOShQ9FbQtbZNw7FTW0ugDGpjaOYfnUCQa8QrOEcX2mCI
/mJ4pVvRdi0yCVAPEnijKqrQ5+FPAkqappc310btT+J+LqSnN11bj7MtnFkn4gz/tHNjYFJOdsld
dgX6tTnISn/ffXyCf7WW0XKOvRrjZBrfoNwDIear514rbP0WhOWNU+4lhYZrFmgcaAO61eSgmjar
T4kQa3VYgfSb/EgprqY3VERTHkwagQ+a4zk2/SfODKFx2UthM9yYazcQqAnc9RUXnCgv9RuSQlAf
1eunElb0ux9ZfidakM+NgGvqV1D3VgzDmGxNmqMxq5jYXO9AQU2S8PglM1Rulnq02Oh5fQWx40NY
7+w9r7jWyXFuj7a7YwIH/QAcm11C1onLl6VxWzR4cIeyj71jSu+r9D7aTP8nHF0DRgnhUYvZBPtz
HAOKaPDEMaFCpGv++PD7V0wxiAI2hKa5fM/JFXZwgyPdGV0tHQwOBxISs21ZS6f7EaNevGbK2/s2
/yDOSRcKgezy1MTM9LvmJpy4MIOCJaUz6LuYjims/ZgmVKl53WyQXXVjjVU/dweAIorUJi7zb5iw
NfhLnmiapr5DWHvzceW5ueDygn/f9zWrNZFAqxBSpOASoUJw4mg/7bIyHw==
`pragma protect end_protected
