// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tYLp25a1jvt1+F0CNC2QJdsfDYrZ06qzP9T6Ga2Wb6IqJp1FhUEQ3iJaZB6zN7y8
a8aqA4fmO2xSn7z3Qzo/BChSdyq4JIGbW9chxBGgigQzbcfW15TCQcyMM83t/OcV
K9f6JOu3jDTciDOsDn/laCHofmFBEz2XrbAoFLvlOgQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9696)
YfjJKnmj9LeOYNj2+q9arvvKlmkRTXKotOFOz8nMhGX9Bh5mBQKl8xJZwKgcozA4
ky60cvO3kVW200c3IZURlvFHbaLKMACL83sVxd2ejdGBLwsjevjyIVhHKRGrPGTm
K0O9OJAVvilIZSzKLZsSeSOQCyevcpoXr3LFeTQaM+XTwlAZqJKgSc0ZVC8NJGk0
6WN/3xlzCnrEh7DLzk9J8IBKNuyln99VWxUYkSUL1B8Gqj8+fCDjwivM9P6Ed1Q+
KFdyd1xCnB+4ugDiWZPZkg4Qz8Gc8Nkcg4+UsYT9OUC0RG8NFf7ESOGkNpFa38oN
Y8CI6Pi9vHYEBUm18rST3SCTtwav7gOSD1ftoy64DcbVitdO7WB8jNicr6x5mHBM
vqYyML90IN3nwFQ0SnERp7CANeCn4VPRW7gmNco92horUgR9S2hTuZofgr/rtEgY
BFXuswa7dZfG4cHPVsEocXeEjEJVzFEHz+LrXe0S7ZZuLcu+mY0C28NhlQEKfYcf
dairHyxLvmd2qendxAy+fRKXAaT1hkplVUK0NF9oICvbX0Y8uhEH6qQ2HXlSHCAO
T/jNlRIU2qVCMk8LQ0oL+rGJfyvIJvX8MyyIadgyCjV+sVv1cshTu3Yw38rL2uH6
h9k3URs9vkXo6n++i+7o3Rk0GfkAs5JXn0z6Z/sJolYgy20WC+2SICRRvrXZH33V
BnXrLnDOwsf2m6+Qj2/l/oQ7w84X0V3sXtmoEiSo7auVgJp/Fmchp+yZNzqc0IGo
/IuhWmR7qM0T3MDiWFLcUXIbcUxsqLkMdK6daAnhu+yxgvU5ak1LOQreF4mEvzXO
dnff7vNtYhFbKNROk87L/JqKbnjczTeS7p0DJ9IwV0hiONfyKXBkfpsnVGTMgK48
41OISatiYZb8tHc1BtSv0n/iDj4fSgpLBpesk4eMjoJAxSyWiNfUilrbctjJlJKa
pB6dKjsX3gRqHDkyPlHFCPtf9IOE5NdVTqZMa2Ix/XBK7I22t1Z0RAqoCBkMDH+L
oYxcguuvkX2iv21e2kTQoebFV7sBpfaT9ej969gLKOKjWZpVCsDNUE/NdZ4DDT2j
Bnd2IWUIXDNHlqqs+qImToXQhQI93iRQ+cpIF1SGl2axT3f2KAMj014jYYU7Hy9L
kDT9OiGBrKIlLtX2qCiJ9zvfxcZo68S8ak7PmRn1UsrS0PQw6WvEdFhAbCcD3NdY
jQWYst0mDYiZO026kEgjMF/TOuW6S1cJWTErdwD27v+0zHjKx8Go019lisHGHOrT
dbIN36WMc5gGG39nA3yBzAEiGvo2Ibov1NO6gAZWJI/6Qcg7iD9CbqsuYKoh4Ipn
OHPFUQ0HFTUeA1JM9oOdPn5GqQorzwvDOtkcPkwveZ9+eqCLIczx8uG+/0CxPw3/
hINT5vuzT7sqH8Fp2Fn+K/GCTHXGPiyOU6GVJkV1BNHnBC22jmeZUJzW4huJoFkN
XLKcb2z5AdKHFujySUVocLNfNf64hpy72SV3S34ukcJfwnHomTYTQPrx9i9Y8NsE
5OPRNFgzTNbezI926IUdAO1hMT28qbqPtOQ8w0l1C4UWa7fVO1pAfn+BCzlWkJMj
mpO9UjYWAVrm6AdQYP/oei1xjC5ngYfDNyzVY3TaxNceUiDrFVJJ8+lhZkS5JWFN
+DieI2M5JV36QaibPCgwKgB6rriD95Vz4bY0/u2RZGzvs/DpIxmx3MAcfjAHOMpr
USV+ltfgjqhVA9zCNCWx4VEgfgnxMrPEbQaEzjsa/RCJf7GBrLiJ25XSqsKFtCIi
aOivb3h56DU1RQISOpMR6vni7UqcXpRimddtI6AHllFdz1xg53ttDwgcadoFstHk
/if959DEkVsDNTH4f5fzflFXWEI0X7RWO3doiJ8S630oCIMO6rynVpbWUZV6/vew
dZKnPS7VFEqftAvV+7WAtV7amSYRCgai7MalswokJVK/mov8124tpXKeesx6kx2H
BfO9jwEW1QR9KmW2cUgCLiQ0zjQdul8uoqqVyjNyimLbLAZCEoogSOBgf3MI0jEA
AetlwN9PTw2RO7nNrqIzBHrU0tw9BmMnqJUT4w/qHoTxGC7W2/2IuEYAG70BUgLf
S+Vsh24sAopHPGBEJClJRq6JpfQNBHV9UppeW1mBAgXJzWvELj/N6pmpmCbsmIer
9GOeQvect3WYdgmUH7SIFsq1g3xQdDIPumz0A7gC4hFNeEebRNwiSjeGSTqIqI1M
byL+JMAzsYf1XX3+EaJo1zNSELJX7mmc9JTXQx63d4mzTpKe5LKN6/5buIQdV9vE
vYO13HBi8xRsFE9qcav6m0+b5QOveTiM6SvZmgnmxR4VQ6ZrwXDU4XVYPu8AKmK4
+pcPq6B8N7LqZ+4K3TMPBKMfptNo+gN9k4ZDkGSWdT5/G82Ja022MfOPP8VFjN4T
KITqONZin8Wiro2wjuSR2YeXl6aV1ctcQpAk864bgycSxfqlnHJ2U0kcJ/eiCao7
mH34wJ3IjazNx5vf9cjlw2/nl2Zwjq9JTMgLQFKqAWOmUoeHZi1MTkbUXXoHLQdN
ihxsmRIVP54YfCX8wld93mZByDDNq8b5hC7REXTRLc/JbLQFEhT2EkIlAAKjmUGz
6nY42A9Y29jAsygFzTvSEfi2JYcC3CK0YjL7+C3AtOaLZxMIGdQzaoBLDq4Ek1y3
iDRf0T97CSLA2X0PveYQlqnTr03eFwShEVgrJ8QCEc61kayHnGFnup7Aq+fswyUZ
frR4fneoK2ilWSgAn7VtYMTV1cpV0quy8kpC2IRFSv2+Y2ocwGFnZAymdn3NGu0G
tj0WP4w9QTRpGTdhTmngAumY/dzbvfKZShZhkUJWlCCAHVgzImlRNi81UBDuO0yv
yFwP7ren+E5jJJgPmS+9ZNK2Za0Wgnv5Z/6LmiUpGW5WCvljp4BCukIbakFrVcnb
zonx9uvrArq+mPTmqY+x6+gXxSPYevqq8h3iQVsc6s4G71qi2YOXNtmF4Uuv/3ZW
m+g23Dkein3MxqKv8XlyUhx+6skFHCWM+1ruD5+HyEW1xwJDf/PBP26ZQIgNgeoR
8XqRa34HIdkZCfGUPiGigxxroSGmXUEarxbthchiA5RGhP9ZMcKgZyE7mz+WrL8h
Jo2TKDSAgKoCIRUPmqrEBpXfxzwxnZzC0E5hC+cB0YjKq+AJ1RpPMWdhhml1tV+7
vhKzPf8w+jvvw/XRcW2nbFDwJ6WE497oMDJ14215RFmExI8YoQ0qOKjicRtBo2tX
fKJHg3hGVIh+f+L5+HTKDibPaOk3uuEta47U4ErmfzTlKNL72NL0nW66J/ks4lUf
W4BsCru8SRYBsHGQHv9/BGGjAO6LjnEmp/OZNNkU7a1EuEfl5bK4e8J6xXuMV2DD
KZq8nbQphGDMdFf3O9mS+n7OnjddYJEoddq2b9zwAvzIrKCzxQ5FAU/pFINTmpXG
5X+OEjy6WzekTQ8gEt8wxUYX045ksMwmIeKREr6bsF7kQP9Kn7E2nR9RC/p7nYhY
hrU2Kwn58zn52CqF1vyfLKv1nMNzl1T9ZaWmRg+zxXlm6QS3JIMZ6HTlvL+g1wCo
gEbdddgbZu5R3M/amsqQYPZOOzKk212zjaqc4kaUurionyAu8gHiVAibtCM7fXej
zlsDxSW6vFfyoeha2LBNzqXFe09TWOvZ1625Ykhqd3gZrJ6XyrqYCYSTngmWXxmV
t8cDsfsOfkwQ2dosvtPwlfmDWdaAwelZ0/QVJK3/ORrMzEXdp0yVx58k9YM+/IQl
asXyLMXo7vlol6yArpZbMOWRsJmfjsJ4YepLgsQqjXlbeFdPUcfiTV7rT3uFFPgp
CEcKeLGjpuNMD0rF7kegw5MOW2bI327qvXxOAZ4V6LnQgXCr+YtnoUQVeXaBMQq5
7KTtbkpQgIMSg5sga5T7ynsV8SZyskFZaGjdsSZSIWgT+gQBkkfOQo8RIAcQszaH
VI/E9RFmWMQIrlODNY54XPuiSMDrClwye/qIDF3VTs85iVjCa8SZ3Mt3q9+sf5X2
6axs1s7YJei7ZZr6BkiGFXM69C5Qlvyhdgp5lx/MUpMAJyuUEVulLTCDkk2BQBzu
1iOyX85cFFPqAvRVWaDux4mtOKVb7aZlMG5s4X3Aeumak/IdFKA5SXhgPb91E2CX
ZjFNUlMr0VP9XSKs2lho+1xKQs2K9Vh52gBaI791Wly6u630tdl/JN17suLEadZX
/K4jy8YjjwRM+yuUW2yuj+yoNbpt5t1nRvPot0FAkhAzbM0No/1JC97pDlajTaLe
6Pv3KhAN4BHlVqeRkHcqbLry3xKXt/24D9BigxzAD3PvChUy5yuqn8DPiyY5Ecg1
24tXkesAo5zlu2QJXZx0k41Sm2eyEHCd3NWcMqJ7OcdF8LoxTdQ84FwREgD+idcJ
kKGu5hDoH6PZZsxPS8AE16hL37vA/LOiUWa4dpGg31EtdefXb5fY7hj0gJHRlX7U
Ze75o83hrZ/WA92oPB/KYglWsiu/Z+BTHwwDgWruH77zGRhoMcU7MVTQp72/pkxn
PlbxJBq4j1tQESdmseBtVH8ejjlluxEy3m7xCbKEAlCYLJtvH8HdVCrCFclzeZbX
ANtm/UxGfZXh5YBqDBHzhMLofqhFhMqhZGRP+rGYlSmUL+2zVwva2SpTpn3+yWqV
Z6e89jkZn4UloC6mEiTYndaKvgj/RJPaiesx8gsiILuFawOXsHCKrw11FWcDMdrS
vnbYPn+RDu75XzHo6j9MgogFnbQvehwCHcBbW+W2BmXjMIgTcTqrv4angMYOM48F
nQwsDaub1NwOLEQBO1EiH1B/bLjd6hA55od1WWAlOdi4NpbRe5S6tfA6f4nKugK/
ND7wqs/SQeSOCsler2UiIJIWE9T+ZUx3WtfVZZXHKd/jUfWkQVvVddKMVpuboLQd
d9xs5wTNFbC5n0o7s0YJsPJJHf1M0Jta3HOsYjnGOZHs//aQIhmVzsXlLhDNPfeH
77kIUhUo3wwXldzNFfhHGLTY5Y/sAFRrurHZ5fxgAn+JW5F0lj3rPe0vlI66nx0W
5BFtRoJumS4O5EJ0xWUNE2DGksj+MNd2Sy4n2AjiwcR7Lhz5FmaxCPY1HPzD9Rfi
d8EZNx4F4IJ9jpWZ4eNgrk2bFNjXjBgactvD8BHSrwKlBIXbVD67BNaWW4BhFb+Q
lbrGOR1aBX3bd6qMn8x3XoSJ0/qsH9Z7VyYpr22JatRjzLVVTFuD4K8YhcMqhDkX
nE+1WLp3mR0IsJU34Q/dTKKwOtzEf5AATxEtxV1o98GQ07CzDWWeVuBVj+AjgXNK
GuC2WoHUbi1JA1o7MoIhUDQvDKWhNjeoep91RntTU1AMaa2q0WSJ1rI45fCt7i4G
Lqa4aBRd0Vu8yXvHFRtjtteU6zDkmYE9jm42+msuSzMwGKKzOlyBS8S07Z1zJUve
pUpDLWJP2VP+pmlWcbtRJICeHxmzHUHw2Osu7821AkmLptMsagSiyemSYAOSddTI
xifwKRVF/SuTyfimzFcM2e/wL+rHQ+a0fNo76gaqR/QbJtuYVrH1mVxkvi5UecLK
VVl8+++4Oq5HD3+PvUCFwKWjDrGuLJgzivWGuiNH3+eiBbbqzpwlAliFDWRtcVrm
PwJLFR6R3Dy+dKW3fsBkm34Nx0pMBrRATMnVPEKeqGRMrDui+ehrvoSxDYealDqZ
NW7rJnnpondJV7mvdhNbRqmNPOrz0Fw+cpAGD7sAH8RvW/xEd+dQxxV0luhlNCQf
6YR0asARS5UQn/NYawVcHofCDKARFwaTm8orF8CuWp+aODmWtz2pKLuAInN1qAp6
XdtB9h5dNxxVfOfgnvZSVvoPd45M98zTD1hYJQPPl8lf8S4TwNZv/UnxrYY3JcgV
eA/uu6z+1q05ydqSG80ihQIS7P43NXSBzbJ2oImoPxW/FZ8sbs53w0JVoOqrShML
fP6FakT9mE3qVGem2Ii17aw04z67cXZBXCs7D+xUSlL2ObqI1gO6lYwlnzQ9xgdf
0t5D2WDYVRUlc0yCGTL9hQpHZkg77aWlEoHvS8zigDARh0NUjxgsK0Lqtrww4Ymh
KNcScuYfGC29kO+zmPXqYgdyVzPflubCKoauaC5PHkPi+hs+PppHRXIqY6bg5QUe
t959jau9C7byu5C9hg0J3YY4uBPEBc7Z+EkCWcejvfp7IWoHcEKSXdfSdqz/v6SY
wk446Pzn2Hl5LSdh4IJ96fL4mm7j1jQMyHJzgqsTpoWaA0uu4NRIc6jx4pAJivxg
02+yo5ptTUOGE4UAUe8+GA4b59oSyDsWKV7loRbU0z4x5Rj79awnWmWi0eStK2jv
bXYxDMx0hN7eJjMADQirVMnUkALsURM3aeb/gxMpIzoO4n/sbKwr5FBpUtFVrI2O
ocoYOsb6iJ21WVS2YGdMVTEFmB882qcDpL4D7BZjduarlGNir/jexZOQxqNCyGzj
XySZrbt+3txzjYCx/+9n8YI9fkkz0U129gL9vPCaxoVeIjAgmE1cc6+rrvwE896z
OybFHz8TTue4i3l01MhMS+UuXGOUWIF/vbe6RfEEMevGs+4K8tG/A4xuoi4X5EEm
hwXzxx2qDpeAcVIjYQDzdcbkMPtpd3dBrPxJz2WzL5FFLNgYZPQESBNMjRYndLSW
+XkOuy8JBNTjqpI69RrWWMbTS4bkpJ18VmTCXepodtrJ3X2GRbGu3S7nS6mPBZx4
f7BE4kHRPR3vIj/Y2twIKT1KGXLiYAEXCMrmO0eWUAKhku1+9meQVHye4U6Ru1kk
Zfq4RqFNybfV2y/9Rqg1yhQvIKuNou8xOaANtv0CWayJIMvI/6JCYd+PAx+JyEHl
zi6onqIcX1fx7leoWyX/Zsg9UB75ENxcSkSoPgM0jH9UeO7bgGXNkyIJ9zqJt1uk
cVPoKrSSX6ZpcCnVghVz5wss4cc1Zv470hE2lCevms8Ni6ecUwgFdz0QzBhRNOFl
ZaZM9EO18u7iUtD/K2Y84FeKAgI+2V8fYdNO5T2qpbELqxiU6sbkXb5MAxcPq/9h
yf7f+CvVmYbWQqbuL1raYCZDMkoi4dAKgqnZ67MqTWo/oaOf+BHNRV+A8KCBxDzo
7gmZ6p/hCG8xWd2m6HmfCM/qfmzbA1YykPlokuc0Rb5/2Jje+WH6s5ahJkL8Qj+h
Tvl88Y1f0p/B/7kTJOzbUQwlyB3vZGtFF3ZGgzlAaMEyZZq/NtX/zksFzCxb0qW5
h0wigV3Br76en9VZvfC0k2xy0qSytHjK60UGgjGqLig/7n+bbWhEK0V0vKdJyrVU
RNk1rZiSQic8L0Nw/SKEPTcX8mPCpRSzAI9BW1jGEwBeYQDlXmByu+wGrwKgzNyz
LTfZN0GBMviRgcVS4oFmF2w2KB4WxyhWqaKRRIJKT8pQA1wrfDWUNS5N1aNmLCvG
loPD+UgtVsKxezepWl/Jg/cW90aIcVxkMrQNWwbWopkTJHZh6uIBj/J8MYOqe6vN
CavqXwGKG2k6TFx5fN77ba6y3MWHCQ1q2MQpZL8vTC0hArv0CO0sWu1imrsqoLez
o4GlwVLCPVFDybs9V3ZNFof3v20Ya26k0qNPiCr1Lms54VDrgOnW5kbPUFzf7ViL
mQOUjpr+zZkm5DsCFz59nwJP9ZZZW2MCoXTDKASkXJjOeb2qPB3jUKLvoIU3gnRJ
u6RmyI6yOvgFaPS/wUAwxCuuxyk05S6ryDU1sGpVeXDMNeg7IqcD+bJO7/LofKHT
FKCgZHwU204NLrDpbN6yorbWRNn07+Lvnbti9QiQqs6D9z8jmPIjvmxl3WgsVdxX
h7Z4ZNGQen+MenjHzM02F25NATDQY8BEGxNivr+b4+6BHa7R18nnMsKdCxqiJqmE
a709LOCS/k91n2bnxEr+z3H/QIDND7705JzTO366aoqxbxz45wgE3eNjzPW6YHiH
Hr8lUrr0o1b9VWkQhQKmX2EdCUVm336wpfN692U//S7BNOZATJITxUKyVxogqULe
b6mZA9q1OfTqbyYzQ93wt30jm40IijSQ7YiCXo0N5U6xnjn0onpwojjGzBcQzd2+
us97UBT2mk6GS99xPjuOg+MtJIz6dRwp1ifTRAMrlv5PQDZSYvTJWbvllwcdDsE4
C4HOtKCq2EFL6gM6oM3cwQGbbxIuWuVdmIHRaLwOGpcX9+Z8mmgMOrW/pzfImSUr
4LwzWHZhsI0aR1XlFlpk6zCw3QhuAoBvdOOnbSZqWJydZ2tHbb6nt7cDtnB15GWC
pfwojJTws6JSoqaUJAvAfisQqLHVfK9e+3eWIkdsFKXImkrremssgOXuqaYJPN7k
DPoNmpeP7b20gRo2TiF3Pn6aailHKf1mQWkoW7iM2xtKV42wvJ5VxPgJpb683092
pATzbVnS2nCCo9xbENQT78EedTih8Y97x2digBprC3kngnbXlFPz7s2qsdMLFY3o
wzJkOr//ef68w/w7hI7ddJmZR1CH36ec9PUbGmqgzV6RpSQcHC4t5Rgw7EwhBt5A
Kdml9fxGfJMhAasV+mZPgDS9X72RTe1AZnbwQCkiQEv/CF0JoiXx2uxCw3BTLbRK
ByldjvKJnBCS4PDR040OnQb8ueTGcdml4mDsVxAf0Nvrmx9qVfT1cfAQQTm3XDkf
Soh2dYJUyAvmRJ3lcUs2LG6lqWc//K0a6JQ/PQ4n/eRJwpENi5oIHgDpKJRcmuw0
0aboZOutKb9xs9K5yA6Ryu1GjnQN2gJJsm8JyTwnlvYV0QA/x1I5XqODGxp8xpy1
ILvOJW1EU5LXfPMFIcHAnvwGXdGqOVjOHj6ESf2CMCW8e0O2RzuxgSt3ic+snjf5
kQvs/B98a0VyMVhbLZm665W26gPNEp/wniJ2hyaCgvIKHppUvgVacFBWI0LcG7Pz
gxnOuYqwU0zUp32W/tYHCiZdbWApXv0JUFrImBcSeqVNGjivl/jDVRerWxHjNuIV
n48jOd80YvzvM94o2Q6/dJ4JcP3ozV2q5+9iM5/OyB+RyIT54VzkL3y7iiD2NLz4
rd5biLNokydeQrvYDpuAgG7uDnflJ4y2Ejy8N8exnjNfqpTTqS6hx8BLONVHB7NG
sK4/6C7G00Cu5W4T+EDOhXQsoKgYlTs0/WofLr0W3tXnAXrzeaB4d5vrw1w+fzVi
5j9asgDn3wv2fBDlFWnweRxFAIaPO+EWbHRCICyTtd6YXm+r7lgPHiWRDwH71R77
cvcqnypwUDyuU07eqMjvce735Dv1BzMxPlhssT+ENQnXVKuF6Nib7Ti8Cwh0/84x
S3DjrjBD5MHcCfPef2666bVcUfhRPBuvVECRvUGcJT4B8IzAnnSjoc9VlNopbetA
7tGTUXBXITsSucBrz02wkgpClfwQ2EU9bpZFkOSEOTsiCaxmTTsZSc0OxVJnNLa8
k6ZNVbbAGLpCP1sILLfOJta0YI3kFbxJzp0YBiFUN2/iQ8k3sYmnYZnypRiSI9gJ
SiAfinJXwKjcqkWkdMt8FgF9PY2luvdB4woHC1e15NWZxUQKpPfIjS0Q/O8Myka/
OvrrpfLSxr1Fg9HdnQErMvB/gCw2FXfcoSYjm3zLus43elMPdIgC5rvcH5Y5SJ8c
H9ekbj1EgpdZfT5vPXMAkcEWPbRA8+CkFqmflIX91RUm6iOPPiV6V+wblb0H7nO9
cOWq6odZq7ZN8Z02+RZd/9Rh+mi/g0YoGvp3QVt80XGxj1wErY+Eq+bBc125hGKM
x0ePyO0yUf3Usx8ZZ8Tll8wr/ipQwjgBY58SGOezC6mqJAWl2ke/wx9BkHeVDLS3
Po1PljvRa/sgtlhpnub/V+G7yukBXAU5vYaHVIBPL1Hx0w9dVLK5ZBciTDgmzKIj
G3HNwXTi5Xe/asb6GvH6B07XU6PflWMJSQIZ1sG+g4UFn65LtGz/T3dijFe2WvGY
UghtXhWVaqf0yEW+ncxih26d1RjdZURxtDt1xbUHsLIg2ozGoO1N/GeLGS2VVoSV
gEFt1IxhksW6Ouj+yIWzQ5IUdLqg5Fzwmr54ltoVwHzdhWqeuwzpjdAuY7wOy5s1
l6jdCAmSzNyNkO58Gqp94RBrRfuFNm2GmAmRkPesLBzFNd+si5UxnvIJGogiOvpB
JgIGE8J60LB9T73mvmHdSJ1w7U3qnVsGxDodNmqc+uQSVmmjBU+OokVP8fe144zd
6vwWilpcETwoneLzfTw9XGU6srT8kNwE0RuXScOYH3yOYCTlaqlxM2kEFQQPPkIq
LdQiYGio8cznl7shuDiX5Rv+11qCk+znBfT9DoZ/eSIcnAYKRioNkd84+/1F44Un
DZQ4IjApUchFfmPkpnBst9vYsTPK241SA3QgEhWJQ7p0zcQreCtGwaPhWoxCgVo0
xE6A+ARqJpwkGzVZcTfkdgRD7Jw6gvpJbxq9OtTQ+mGQ4vmpRp1NwbafbDsCyjKf
12PMSoANTE2vqoJ7I1dqsMCgPmjODiq5u6cPQtK8id2Jl7ZuLPWWVk+ZpeQI6VTp
RWfh0jpCacaAP6sZNABFJekAuotP39+chMOOgJuLLbvgnLQM0ejb/bDa9PLE3pc0
os/O1pvDGjay9nyoiOQwMPCZXAA4Sm3Pas0csNaSAWx/QG/dEBljztIi3wBc8KNC
wFLwcwlql5B8kEYvu/369sPPQoNGu9sovJ1zblKFm+x2M+yuUer5GLCkYNJtiQje
iS+q1WlhpL7oAzcVkD50SpCieQtQZmJHqjeXFGXONQnNqyv4sNuip7pC/UbxoJBY
0QGBPQ1SLSxoocrFJpbbj+8lx4Gi4Kz+yKPX77G5kACl2bHncwPa78Gfhya8zKT+
/I+v3LVJACeKm3hgSzTVYlP35m2YV5Yk48GuS79sPZLdbq20O7KYAugIjjhgOEgL
JFr79P9YRXOuvMjkD4QsMgksjqf0GK2i50PPRssx5C11is5aLaePLz7wnd5s8MGY
HcORI1t/VhZDg3ujK0EuG7vOt5h/NNDL91+BRcTNh25xRyiEgxDSHv6C6Edh6VD4
90Mj2C0rUNYSVQ29TTS9vDFgbHaL55ifqLjgouEcUjwCF+7yYprvaBl3B9xiccvR
jV46nRrsqPlSrX24/erDJnW2ColgBge32h+lz3ZD1SjUYnytnlsuXS3lN0ZqbmgR
qItzOgcm1l8tx4xPW3WWBGD2RmIRucZ5YbQ+ODWp3f9wixGv8KpWEmM0t8lAcYMa
0VhyL8TNIsNrm5iQBCtzDE28jXh8DGZ3l4IRkxGH0hgE/6ffH8oLxXIggxaU/3Xs
O8yZaiJ9fuTUDYvU7OX9XnXTIcplCgy07Xq3LLW6pXQU5dXZPZgPgi97bu94UVLP
KGX4YFv5osbVJJCU8R0M8liLj8Q8MHz2aAxCxoJClnrO2yUja+TQ1ONLA1h9ij4B
kInPPIx+jTVoFyxAEBmqQvsrs2BIyHFF/MRZ8oJu1PX91YVOeadlA5aQkvrYc0L6
C8dvvNuhoKmZw8ZnLFAnrLmQUA1PZ2JhOvDlXgGIqfoZYsfEJe1s/U+1uv8Z8gSS
VAjvVk4q3L3sw1dKBRSl4EGyS7dCng5NBFLuUXkis8Z13tLTwhiXxr2paiJuVL6J
8X+jK/vTgYyIj0D4gcqeW4uY+ImDpys2gOCvi4Y5mAFuCuhrEw1jJ+2X6v3E+I6P
NlNkmfJdhVuzFgrTP4G5ho4F+GiLGxLZ7sY5aS66vqdAVh3qYBoZQDxj+/GOv0+X
T28hdM4I0bAc8ibpJx80qy+f98V4F0xBH+yOUQmNX5hI+mRNV+uaIPUGbxn5eoT4
+Yn/kxKy4Wcxt+x8wydu7hhXVDLchyOJDZZJ4wp5SKdMLMmTFl3d+SfKfaiKbnSL
YnYor0B0r2dorg8x5GrkUbzAbq1WbukfUlpgccF3LtlEYz9fJ66MhO4TiapQWiui
3v4CodhQXcvoGYA5WwdHl50+M7Xw8vBvwJfWfrFdsB+avnEEwyIobM4JgFrXGca8
1haN/K4ZrNt4vW6FwBGmsGMxh+Xzx/723HdPAHlTQh8rwS5FHjJbUIi2BxUV/zkl
uh6j3nCgqcpOk2ifkugy0VfihwY3wkmPg0LKenFlI4F9/hhZjCivENDqCLKTkRoN
OMI29glW45FZ7EWEPoJ/AybNIfwdhppI44u6XoG+6WwXSXoyhmtAqq2/B1hS3qJt
3vH0E+1+6a6WDdzXEnYCWDLqDUW+ndYJaPQJYSghH0i77YzhOmw5Dx302wxLNohW
BWmPnF+rzmJNlI9JyFbJsnSbhJFYWq3SKn8Q533wFBKEiNxFaR6AjnDsPZQkvOwY
ja1EoRDanel/ArgdKrGt+CmqUOl/QegolOHYCBLLiYcKXfmm/44jF0vgCEe451Ga
UXhb4NexqQ8K9D/jpG2cNUxUIloh4VEMUPbRJ4QeJrgDHf47DxrFBJpfY/qXDqfp
sQBeQIQbJ2SBNMk5+x2v++XhDyWmpTgU0PAshAv99Ze20tvlLhg2rROxIVMAoI3h
S1T7c7AF6LLS5NB/gHdADy+7m9WXzJ6rBz4LI8batzm3wv+ZxdEOZjv55O4Z12Aa
Cykp/nzKPKNFYtL8j/UvwBeEVGgqyrQXGHXC4XzB1LUInmJD6tBk+8P1yCBpKk4t
33MLXiqO+9flGC8Cr4xeB/OT15dh0pYlek++gueA9f+7rP3XNhH918sApvvgMeMi
qomEGYxNduGM9tfFp157zva2PytuoctcLwt3HCcb/b4USdbptd2EpkEmhSNYuCaZ
YOJQowZJ+Fk9/FHrNIOrf1rDUXXK/qqjPr9d0FhaCd3ZrwSj5LwbBtfu/d7Orj/O
vmlzImeQIdyZnR4oTaH8TBCnzAiDoHGvBppRDXGhqMTXG/GSak+L3gTV8ut/ZhDN
Whbd7T7Xu4PTD6XFCcbXRbuM/xR9tHPBB5aDSomU9ZrWpz2cgoJE3DaFY6wdVKTa
`pragma protect end_protected
