// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ERIwjqwHIaPHTKdL9wdeXAR//OcWFbx8xVQ+mKgyqN7pySOXjOZb+kn2pgxwonHL
jio8QhC5Gpk0bGvwmTaifWolXzPErZIlXNHZHRCf2gSQB57oKLrHh7YyCFIf5ug/
JNi/WPvBTWx7jZxzDuEsfQw5JBxZSGnNIkvVqEqKOcw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19568)
r3ksMU/Fag6yIPtM8tsYKQuCdUTYtvH8F5Q+WE9DjoJKh0KjEfubAzMrjYGFKkuJ
6ixHi2OucUDGe3xwoPc81brMjrzkQZ/Nb1ESrG4G66FfL+3ByiedxfQ3FVfQqmei
ze+NuGIA54skXBq53//Nnstte9wGST1sukwQQOQ712XkrwZ1IcOWbpiOoavVhv7Z
OEh0Ts1eZIk5iKR6+I7vqH13R8an02AZOvPjocSVqb3cMCufi6UNah4bhfeUYYVY
n+h0DycZLfj/oOBRCb6GE03lwCbXCQ+RJbjyRDlMQsDhQOv8V0NSEDirJGJdRRuh
dEOv86P4+0UEtMd8bEYXPO2StRcWD053uJFR/SykRgbHbw/KiMDPlJqdPnvO8k5k
S/1164agnr2dfFU7P1Sc0hBxcqVhT5qgM7eSQoVEvWNWhTsxFfdRqumluaMTzZlV
RfKhe0GqIXqEku9oQW/CbjJDqv2TI0LfsfHKLsYp3G9vsNYvPYmYI2Ibis3QJpqz
H/2nlHklpRpSjlShmqcbNoJgxIGbv1bkxAc5ujSZh6PA0IJivZmQs4iPzszubvXJ
avuXLRVkkzoMi/Hs6bumYJyrg1lcyEEp+6Tf+rdPvG1Zqdkr/D38uMClYlLjNk6C
GzQNErkKwtoIYlS1ISMAJxbrgnKyAWE8iNpQ+rboAOnn9g0piDqVAZN9qVjLPllx
uVYdFQEUaDwxJfAoytt4Nnc/CsGr+gH8aaekqKNTFeRk3MljzkdxhNQ/0cMI/O8G
KARl/V7jog6RP7aG1IW0st8NYJ/uRnZ6LvD/epa9Z4KzXklZnOfpGsJvWo+zbyY9
KtuJAcPD723KBueSCiVq97CYq84W+s7w43RIvNZVyAwa1IoZSB/49veNv40A2DJc
N18uwv/2L+Ulj8tY6otZGTKedSFXGZfODfzO+0huaOfv4NxPFMVom0Ml9Krd/fAv
gW+UavHNVix3o7fU2aSfBfZ1x1wdeHgFzb+vMO+C0jsnvHtn5a7yJLoabrb7rv+8
hwKS8ktx8NdkU+OOjLUfuoGpUxTzGmX6yRBy1EJUzIrARdt83dKGSdcIFAJxQOow
0FDjQpMo9gxPTOZ8w/hHgZXd5mkpdERialNDbzyyTUqHhZ7kKZM8gl7mt/zcNHKZ
/fZPgjWE9J4ZIvg5HAHaEOXGzzxTSu46ztkYJgSLO+t+0YXxF/9qrMig+n2zIPSO
44Eosct7lWIGxAcl1bZ52+FaZ6070Q6wanvFP+suL++eqUbbsYD1xAaD8jP+VgBR
wTzd+bvbUcej0rdS2DeEcF1LsVJATHajXpP0JWeX8upBexivAoX4WTNAz42Xeabp
2p4DYA79MTqVapSH6SCfK5kvxaGNHyisyCGMEt4wfIYWKpl9vb/UCiFaynPBh5N7
iBma1WJCyGagxDj6bYdiAChq0aU6AUL7aoI6TyzJ8a1oVDW27NTU63rNvd40cLj5
1C+3J4TbIlGbWHLy0mI97/UIcMNndh87Din8gb0eUYtmwQdDMAnRfkck4Niwic59
cl+mwhKsi7l0QaJNqYd4IKyFks5SgePW6UYlAqTBsKbmnE/c6GRH8/QUOmy5nAAO
PEFoPd7Du+zck6WFKNCf/MEmXNEcrTeHtzKo6YohRcA1TXwfpIF02hV1YufeXMJe
krBts3Nea3x+dLJK//cJ6coxlMp68K2lty7ioVaVXS+ixoEjEWiZoxRASKx8uyOF
hkyoJ1O5ahRPDNaHJJrWK9f8GC1NyBjILuTJQsAdgn9SbTv6XYd14U8X+VKTmJos
mJIM8Byc7emzoYtt4+1TvJWRGUK4GUiAhRg0rzDxluEulekP3i2nBXh5VyLTxQ1Z
tLoZ1djEtK5H1TV7sjcY2/flYr2EZnh8O2KRPN4NupcVLZ1vXOOW1FCw1K4Pm8nV
rqkMpJM6ozDyX35WlTszBulJbuxSKpNeOe702St1L8BxVeBrwZzru0i/y5t8L1vH
D8SWr1FjduKvwQRd9+dx72igUuA10cJZ3GY+RP/kdoAqCHu98wBjvE1Ycu+nnrDN
Bo9ABVcApba9Bvr2lLmuWjjoi9r0AyIaGgZTAC1cc7BCFOV46vIFQFih/rt98oDM
xngU/wehbH6QFfpwLfSm05ebOS8kc5E+CvhI/TPsbCUSiZO1C0PPmP7gMnfuzbav
htaAsVULflbGOnvCJ2h005v/NmhI4HpV17RyuIapHzUlfkdBIokD2NDBBwwQS7Al
C5fiRQqOkaSAArFzFJp1JB/EbEqQjfImOHUO8ycQ+c9u8hZOwzQMzIfMoMX4Chys
TYkto5YE2q7ASy9YkGCgcyM3+Yn4eAebyDncwujjm8dF8aASbmXgqPzCFASggdHu
HgsLMIHYE3D+KTJZxdwUz2i+9VF77FDdFZLXp66343gpr9VOzFVZ+pdqnLdRN3b6
CncQVn9hnpW8WsKTDAmM6b9+B3X+nwc4MpP3AVpDStwTTk6ABYh+rhRG5T4JzZMk
oNMOgy0o0NEruGBmILuBq4Ki4W7fcH3DnzbRlC53vFmZ14qZBoW+ZqCjaaLe0wZ/
qu+ixuUYIPT+sKR2SaLiH+yO/kweitYbPhoKGernBB0GGYikfrP9JA/4cVIBPVFY
sAr90ZPirAmDHwx/Q3+aZNoef5ZhH16YFEOSeBqgjcwFyxCAzFy0epNJb8BR6Hwh
WXvd8ZCQnAeHRcY9hClMe6EiQ8aNVNCT5MzK03LhV3BypTEeePA3UWT2vJWs4FbG
/nmXpeScR4GchzvObnw1WjOBRKyzbHgzKuEWyaGaD8B/fAKKp8TYOu9fHyCwz+zk
OGHFL81V128m+XvNqDkOwzBQSwPWDiSp4o6rLeVc026fR2/paZXzpnSrc+7olYNV
4Pi/lpqrt5w8TC3h0Jox6nXmNAgFzJCYfUyzxay7P20OLc/OgNLr/vTl+5Yjqj3y
v4A20dg+D5rApqS4LMq0fwDKFlKIuTk3k34r0kLw8hkuzhl0mDRdza+9V5vYIKR2
W59H2TbMoK78I5TrsHfy6UTC3aZyCnQtT0YFJBoZQh2p8OkFZ0iAAvofu95t7+0S
Mxvl1q4oyLoEiwWS0mGUgQVuaDCQYNgyvqznG3hMoSdNPOEv4zfgns4D6Zpoc9J6
HxhaC2ayfT/LotPe+TQM10K8MWnIh6poI2ZCI1whfKsyM3FU69Se203bL7njxA8B
SDJ/ODEVQs1emTNWZfO/eGhD4+c8VWu3Y6VEfpPO2OJcN+Epy2lC2dUpSK/AH98A
uXuvI7A7LZAIzPgrE76m8eGhWsGoU7c2k65duXz6XyH0TBYwUOl5PhoKygow28wL
b/lVCgR5xNKBSXko/6wJx0CGU6+Qraq0AWo6wgpOPPpcR51Nqh3/CqUDSV7org9+
yfWYRfskAXUxOz7maxC1vA3mAW6mQX9fqjyJR5g8AxJphp05TZ9Mlf5XTPPzgvtm
pNZZZ0vIxkBcDW5c3/8xYT5WJX+FqcbL5WbObf5MZABdMrXkTawBYg6qV+lCiKxU
EtNXfXDtC9ZpSnv5g5SuKaQVkIdtq5pML0rIBPYHFSclbTad+96qcD5jGyqozuCO
jtK2ElaqwEP/4T0tarSoko+Tm+Fk6tms/SsVK6VZBMzTjMgawibeoTqPoAaITD92
R8cAAe8tKB8JxqRDYK2NVFZxluVIPpv2EAJOCfqHTS9dOyo0wb5qZcFUDJWAJjd9
6Ld4heHka+VfAFX3NriRz61yLzoVQA/ux76Yf2a7QjqXKwWX9P95bpzenKym9hwm
3NGWkPrCKC6qVZXZY2XdXk2+orSj+bt+fq2VLlM60uSZEz9/N9+l22czX6xcboB8
mLMJpwHfrjzbK78bf43X9nnNMJDAVa16/oSTVhcT0SUr6XmFBNOw1iPySOqbiu5X
eV8OpZOWoFPRPzCM8ZQI/HSfAghpPTZ9bBfeY2jFjgvyd2gq1mx2KrSeRC9/XSvT
ID0FLS14WycOF9oo03EGJX8AE7+wwPGE0B/YiWgKDORhrl+tBZxiVo7kXs4CTN0z
ZxzcwcEUJ2MxRpyObBSPpkvC+BB/6bewq6l7LmIcCnOL1YtsM+2JrXfMzz5d8ksQ
4Tsh79GygvqgufNkdTDVcbqI8TUO0l6C0ekpIQh6YFYblPIn/OZksKQafXEnmIwI
A0SdZReNqhxaBWX4ZHjYpU1Fy9IZPo25anq+zG2PhfZGw7uxTmE7+GF1+DwrpaDx
DtUYgE6NWcGAu1CGxQOEqUPIQk8Z6Y8uCuArs/H25Ur5JpbK3FwB0vJU0qZzW5Dk
jRsNTASKcA+XWGgd2R8npIdFnKNjOannhJCcAJW5N4mC7QjTXNUO7niq80YPpqEb
FdfvyfAd8YWalFNp4TjV/Dz9Ti3HOTO5ZMAsMcNzO5NdiUJ73tmvwMqQqOj93Fau
J5f1o4VoxBLH0HpxUADYQNf+lZQbOrz7dVSdNRXVEvzPk06yO1jc7skFPyS3F5DA
dp6xkzbI4ixEtO5a0/15fCIl7s3Cr+03sisDG74zpaJmkK/8V53dq6K2yxm6Nlzl
wZuM5QkcZJARv2mjy+5nWmOrtDzuL7kXOQq7degUfzq73Z4OJBjidqQgb79+7Awe
TdOkmNAKD9ZdQgohhYveBrxjnOKkmP4+g/pn+R3P85SEnLftog2ozTFy4rCKpA+y
1yEVx4KaQbfE4ZhDNoZQEAaW/Ht1XCKQ3HMzJl4iYBBn/3fAGxNwQ0fJrJRjM4/P
gauYRxjbi1MYOAa3pSLVKUrWM6uc9u+GBUdT5Y7IKCxp3nFjyMQbogmWnnIt2L8p
xqBin5NMTzjijPQV4I4C5B61WIspSzZVjdI/0f1Z54kAOcF0stXau3UWpfY6IbyV
VKu+1ay23p7EooDbjVDMVu/LdDndjlU1oULAsCYT4SgvV2UxUHJFDUdkwIhngnVQ
efjYFhlL/ppONIZYYFIxWwTjlYy66/58Fkn6domY2fgiGw1tfcxDUDcIkWHFNuqN
zaW6w5LDBuqUPf45UGRgaQ/9fCEMpLo5AwK/f1q87Qgn7wFSnALz+obYR5pTAo87
SDlJOZzWjj+H7G+SyISNDNdkxzNE8/sYNaQiC+sL15/kO0QHJ9nsPtob/vJYNjZq
mihFD43ZIm+U2ZCaujZzsRUchF8z9d4bDypdQA2tzRUYItBhjJaf0B6GlKSxW4/3
fl4/3dlvvoQBCBqviciILobWG8rxXYTdFCMs4JSx6A8gFvPlKCQQD7KZyYwYBaEe
In7wciVs4INNclc+LqDaeyfR/09tfGSToCbs3Fv7SoqlNPrr3/6dU9xsNlgoTAme
sFBHfF74EExRBAJ9NgGkLfKBOMaL1RPrIOvE0Gf7U60PruChC8M0NgJExhzw3Bg5
1hHHrIgrPQJFjKSVgnxxmtx0zOwJZuoiiAtezT3ASGwvL8mnQEU2wGIytxRSyOeW
ASgG3dYxlqXHH6CxHGZ0OcnavSFHx1lSXLoiurTwzyoIg7eVP8rIM9UCpjVkz97O
Jdbyg1IOZQxUS/vWzBMSTpmQuwJEA/r6pTW+QT9nOkAcY+QAUxzbB18vCbNfkddY
jRCGB1wPtfe7+eh/KdNDASBeeqRMcGSnrGKht08pSN6ef301Bi7JM0naOChh4aW7
IjFeHz1TbKuToTdAwDDhE6iuI8Ue/StZA467Ur/UjN2NmzdX3TIJ1MYXRk1+ZJUU
k0o8ahpn1q4iwt8m5zVfa6ldaDLkiYxA3R8lk//RUK9BVbKoYtGJnnH8l1E6UcFI
m4BqjAGpQix3qWF/I6L4BMr187aleRh32kH7/j2gfEkgmQLmo6kFm1BRuBYNHMgS
ME+3N9T/rxOFxykK5Sox5ig9E/r5s0QyDZs4wjLQtvGUuLVOZ4S9ozWCJF6zTH20
aByDKowe9r7b1VHuxV0W2NOI+eYtNR5KoKJvWzfTH6MZlt8+1ZmwozWtIU02gR/c
MNYlg4GxdkQM7rHNHmb0PxjN/lwyYIxJhEuIzehS5/aCBKUjBwwmHzvZF66yVfbg
zVC50wElIBthWwqS+EufwTqVvWVgmmQ6+B39SlvEUiGwrv6LzGayqeqTPjnGOnTO
GU50oEyC2u8W/uJA8LqwfB1ZZISKxVqJj22vAlRSUHiYn9QkpaFn1P8Jx9jilN5C
54Hjr/frrfwadGrSjrcUmtcYTk+aY1Evo1b2ukGj7pbTxoJHTxmyzpLMFeupdaiu
/e/V9dzw1v32LwB/GrpHN7nXwFOkPZZ6tSrkZgmlnD2tFm/AMAvPsS3oanrixnw+
IF7PWtUeUjsOjOqYNBMjZNkyLX32rzTMSDloM9PIfsTdZeneu4VTYC2jvZOmpu89
kH3L3ikBW9hTDmCILvXNHudrcKxec7FJYfj0crYWmKBzZG8/ijXgLCSFHKRoqMZp
AcVpUER+uKQRWThnkizH6uEgBT8drzYjHl+gkkdvYQ5jncrcI4aWmVaRuA8E69EU
2vqmopgrnYWVWa4k5zY6U5T4icYyi+tzSz2mEfUz/uNjuFHWInWQ1JlhSBEhgOjk
kQUuVInQl378UK6hXnbZ2UtpJfMTlZnn1qgA0s6qJUEKIoJO/BTrXUm4o7cbmTpB
+ye666aZLInimcdxYz3PiVbNhVM7ZjAkq7xAPn8sGYfbs82IrzYDUYIvzONw4SEK
cM/VfEx+TzWS4K7/zIXRaLrpXcZjZSDRy1O7kPTaascKAvbLSxCTv6p4rMHTY+BH
tSepGqiHmKmRzfy3b1h4kJHn3LCOmb4uWcrcatgy03EG3ZPd3dPcpMsIsgLfcgDm
oxm0ydQpclZA5Pm0ldzni0/9wd/12P4+7PnRhjvYszg+E+d7y/0YM/Z1cX07rVBe
BgQfJXmdtPKG11pcEcJJjb2c1rLTC2SOjsaX+9LfoE7nYdfaMr+eMxO2IpToZS49
X3IBFVVzGLSBRhYSJCErfbZYq0s5kn3rih1h7hFEc6XEP7Nb5bv2fCd5mLi2KNJN
H1+roGWjoERGQfn5nG3mstJ50B7M+1tsGcl8MTiclZTU0IEeDffxBfY+nc6Tv03A
cWdnSMQvhqlersrylWyrVhgiBads6usUR1Ymj+IWXufZ8X10U32XeAGGljVhUJAN
PwwxW9ab+KgUf9I3Y13sOD0YvqllwdEDlPdVCo7bgZsbTXG8aXYrx2oG21lxUqDK
FtRzUM8qJ2dDmhEu38xrPhbJ6KFU8w6uTs3WCt0JZeexTIDRHwg80GqF6Vusphul
U7m3RGybDO5pRKLaGOhoxULN5/6c+r381I2uR4IeEq1wjF2gb/bbnqQilgmYQUYu
2J2pRsWcHyG7jISlgDV3hFD9lCnEVi/n6bYVvM0Q07WWFo1PpGPKcE0JTiB6Zar4
YC4ux1IIc2i5MgE5+bmF0+Om1eYaOmY43vuGsfMHyuK5fcOaEZSEQeWSsaoJ7D4b
7FaPAzTTx2kaZ1AyaQ/vQFozEF8jZ8tpEK8lxS2kwTPNp24+zL57i89FNQAUwgqy
A584e8025rsAHt83BTzfqaSlDG0Jy5Suvva9muPhYGp1RZjJSDH2iaxQiWEJcbe2
6AgLOyxeRPVxLjjzO60e6Mzw2rmoL5wEIlafQmfrP3LLuACLiWtlBsTPAHU856Bn
fEYbTLv7JhoS8Y6WQYRHS0BL+WFFudJP8pfBFcBI/DRbUR9xmcypmmWCtOoSXJhJ
wtVRfC5WZVt0cZVI7UMTa//wRdnLE0XsI8eHVYvuNBGS7wudifH1uHxx5QO2i8Ma
0K9AWSlltfoM5XGbyIqhkK0DgIF812+/33Y2wsS/ssgsjX3v8yA/y+D0LC2btSpu
v4FeIyVGWcoKKDQdzZAtjpzKFM0L1jnKKYJgY+8gE4DkCPXl3Cl2HPtYe+8vscBr
SQVZWeJh+AsMslp1WeKuF3xzsyWLMUBjFRZ8hg3pYA4GI9WALFf6i5ZYGqTUmNWu
AiYPht74IB0oPLTWCN2j/em1G+aNHDLDHZ3GaZEjxQNv+ziykE52wZ+xGvqIDIQZ
hpLK4z/oFKVafSRfnn49p5zYf9IoE1VW8yXwtUSWHYa0uaIhTsh8fZXBQuRWMGNf
uBw49y4EuqefUkYgO1XoGx7gIb+/SCGpEZgNeBpjK1p35AnrakqtH3iz4OgCxsk8
3lg3FW6SPTyQpGvES2z8AOUqZABPmo/ttRiFBGH0qxBQCGc2Ov3ESUkx0YnKUnlP
uQsiiOVT/SeugbgX9PB2RyK5uEFHlRgsxT45z1QJcwO77Vf6ShVv42wMq0DpnmNM
SwHKjyMn29rr1ZhQEdYRgXJ0VprCPW/X25iEgC66AoFAqYwXiWQy7TI+mcOurF7e
z5cjjARSlg6imj0ClMe2sdFrFWmfj34lWTWohbDsLYg0VgOWI272/Nwnhupj+cIH
cjHTOViW4lKKp/AeDeM0yS0B5r9nh67sXH+OmP3cg8uzu8EQfkXjXivcRgbfL+Tr
2S5RVjGH7OIC5qY95TPv2YSaNYTYYV8lP1hUp2Ps0FgEG2cu6+xAub05jymysBtz
UdemursQooKRfnYQdCAwbTBAk+C4Lanb9HddvDXSMzztsg17He7WOryxGCd1pVhp
vByWGcrKHm59IqyyTzIrZdrWx6WfP0VO4wgEZ4iDcrQWJlS7I2z2hP60CpZYL0iu
0ZFEEr7ddPjehS54UbNw7RYuuxwzG8tgC74dQOmlnue7+ey3f1xgO1KAEfKlXlJ0
qKoWxdOXbe0kPg4KGt91lDU80d7hJkllnnJjesp3m6A643N+x9t/tBS8IDx3Xg7W
z/gCdxB+DQMeuQ4p4G6p9/11EY/1lf9XcoL9E+QTb7cqDEFN3+SmK04u5MlsAPMv
Iu8mLtVWzbPgidRx7/1ZenJQNs2w3QXvDtLlrl8DzBlAM6Y6o1vF94yCAuSKgZl8
0EesK6P0MENj79UpUh7+LQgs8OfZN2Fy2Z28zk+GJzKfS+O87eDvRe4N2P3jEIZN
2CrcWXTg3MG4dgE5giCA6h40WP7hPELOOyt/D7MtYr2P77I7awblBtgxBIx5j36+
7uZ9BMkMJBz3K5fTR4/zFyCU/r3WvBbplQv3pYOBDNEK6BDPMuC3SBAaldzpAbUF
K2tJUiZAVPceDbAwvKUEBVVIz6b4PnV/q5imGoXNhzxACE+otoh2dJSROzkYXPU2
5fpjIVPmEUy0iYJSLpoj83/85x+B8eW0cUc4yPEAEuoUz8vMUl82BkrycUEWrxjP
rdHkgtKHJVfmaHYuMUUQcFcWNLiWnsI9Rag1EBG4MwyMNx+BsWFDCxmNSvZDRED/
UWg/s+QHsAD7vvlocZJNTBdvLdAXdvDbw2/tM+T+RE4joPF5AX38dkzq6QfmYJn2
9+e9DQ0OZ0wQRw5cPK/laJox2LHRZCrG+j+njTRSc7eYQ2eNOxlNdP+qeCr6Pytw
fxRsRBZZWlaxh99rxMy7rOrObgWZ5b+o3zbKJgn1zHZ1AirLDKcbm3gbUb/S528V
1XBgI4iE7WCSyI4r3j7UKkYdA2gIx4hdumSj0IynzZzK/JNjKOlWrCZRSIz/YsPM
we4YYw1KOc0li6FfoZMGMVw7C1eRCStzqcUkt+spDx0ODrDSHw1SfxOrdVxy3MQw
n/HbIrKk+6hgR1HU0jVl4Z4vUde7ha4meTkwYdNCaxyKV2IsHyTKMlS6El/Us6XC
vuSjcDVJ9MBlM7vEaIHJbBOvLIoBy8jjstw9lEcT/iwjT57xUyccyBOCXPXAZidb
nT1R3k4VKz0vY7GwbOxlOpbauhaJ83H1gxLssKXTm29XZsUhWOKyr6eihpHhzZNd
M5wRSaQofCAF0PPQ3CDuQgLTGo6cLnCg71HSJlsRaDm/eujRd1+CGF4+vU/eDA07
jV3jTWjBnQOeymjMksaX3kIbylksI85wrLi6LzvErxdgW2X/kI2ieBWFhXBkmLF2
yuz/HJAvC0f6P5tcIWQIZEo/r6Tb3ploxfWHWWmkol38tjO5hw8ejWrfYN7eAUD6
Yk4mRU1lv3q2uRihS9T6kTE5kLZ+8YBWZT0KRh8yInTK8NvoRP/nPBLKRQA2w+QC
ZZm712ydO7K/p7UGAP0j9vcJzxB1A2rzGjVALBFSGM/AInO+ggtamU4OZY+vJMnb
w3RTgXOGllnk8PpsWDuIQhZaDHj7GC5tQNnz+In5pY04k+Angno8ts431CzdcRkT
evgR8lltXWzL2yOK1CwwtgYB8rtEw5MTrOH5c6Qr84TWalp1TO8H7/Gq5eU31Szs
AX80qUPvGEeWMkBRWzqiFeMI2jOrc95NRdypC/luSVdKs6Iz7h/SNA4YtiBv6Go/
A+aSD8rtVnGqgsnoUDA+AutwsE6oYIwkhP+P7MYAY/m37oN01AJhD++Xp20XRtR8
XNYyhot6zFP1dgfLHsjydrE7jTxf8BleddnKB5QTNwFKzdP5JBg/hH4MmOaj1QvQ
1vdCQk8TLWaLDHBVZSerVG/WM5051Gv8r8R5VvtILJlsDZcm+a2JRboKbNY77l2f
zXlXvqTMRJEgZZGs2hoTJy58NWBfJxSoh3Lrz8maW/4wuL/BlYxEhxgrUzGNiOcy
2N0A0aXAw3PQITJ1EaORuyInYi8X5AwFtXpFpLuqMIq5lVDecikOFDtsvJ2yTDN9
YSrpZPvmmpBiO9XJwH2qXbir4tzoHDaMxOpNXrYT8m5x+CczisGhUpyMy9dDpgjn
2M5yRiG2ul/MlW+zWYNrNKJ6sVa8rc5XnxLdHtZaGOhDqYsZyYVQRQND/NOe2DhN
dKaaZUiACEQyIIk2TvnDWBf6fe6H/ItJFzs8XlbreDgPrvuO2oThwx3RAA3itHcr
VT2qOILx7dUymPzzTt+Pcy414P9Eq0N4g8h3ReX9bhrnWn0zCcR2pv4ORjujUl7P
xZ47toVs3Q4XBIOK77By9aZm51kdMt8I6Wq+Pq34MqKP6g0QUUzYT3GCVgwsNII+
hTi4n/1FfnmbQ66xwutJxN4Jzhopo5+09aJKPD1YuDxkA6FAYkSV8ccYGiiPpiiv
BQC2xYG3RZPudpKkZgSblayrbzISMn4T4RiFBlbgLsD15jO0a442+A3Wdech5ED3
sjpVZb950KMnwJmiI3SF2b4nZEABESoo4pm5/dZDp7ien1jkblEVwyizkio551dO
iGDa+h7we8IniP79iEI6H1hvFGwki1gbDSJYTF5h4VbGNYHS/KoX/vD6H4cJMq1w
iWKcpijmfg6BjDdITWgZaAHHPdISX2umLE5i2rF7zha4OBJeAPojyedNDJ+iVB2x
zpcz1QD6TQbgNEzg5yno9sklGv0ajqcs07MGaH4+hf0+tFm9/syzB7NI6g55Db72
IjVpgTqNYvZ4PUWCt+4uAWlTTRT9UORDsZg2wrRxkrgjsbdpqftzbK1InvZf9qO1
134lrdasHcSBgZbJbO+KIBOS8Blyj8afYEw4aOGophbcp/D8ecugNgCrF7fIJW5n
HVLuHv8QtWe9nQR1SjcoEbDaQ7CJo7AbNu6kDcx9UJS9UFZkzuT9Tj9R2wkLeNPK
HNjW3t2zSo1w6E4JSrT9evRN1+edtOq2DDWjEPoFX/iMh67WI/B1qjVdkXGxJIQ/
pGKAJwNLiH5rc7pg1TSal40voQBwQLFZBZNyP9S7Hw1f/ShASpKG8f1TB8sUX40z
WDOfGxjm5hx8nSTjtY+7VQtRT5zcsXz73VpOdUmY16gDxTcyvr0oySTRBcXT68DO
LAIIfWpoNHO2FrGUkjWlKwE3kKpqUZTavHXpXT3h9r2N/NXWNyVFXEI9TmDwvU87
w3firSQGsJHyZ7hFV6rmbWclHdcm2Ug7v82YlYAKDopGprtfoUoJRmhqRaZv+YEN
5daEc2pCYmOYtdmhWrq762H9Lysuf8NAfhlyc3QRpMo7zQNZ3t6S00OA4Iv4iaxo
LnZD6tsG5l9HxB6/ifCkUUHZt1iz9xaqamDHEP6R0vwIINaviSVG/vvuujh06S/O
vpe3GfgsVRSPqODm0lYV482pWj/Sf1gi3XfYcsY7zDxjf5EtJnxi9R552CrhbFPd
4ZQmDRs723mm41kOaSOiR217qIgYbYKl2bs0pvQtKV0tyLZzlSCbblexZiBwpP1X
E+plJ43OJRndPRLkw3FBDC7dm3HNYpWnKy/tR7POZCgLT6SrJ/ZV6vHhSaBeQ/Pa
ED4xhiPrO/w8YAJwCCDvdCAok3mfeSW88tsQMxe+rDOnj5AHJULepUXaAKMrt8oP
wqEQY9BklhLTQkPYkA+Ou7IUM6BAVXvYwc+gdZ1lFZ6EHzqBsi0ZZ3GUE/2jt8LY
QBU7ip/xI7QCBBXJKtHKvlES4cbii02HcWlKBzwVMsHDfpDCgH6t9R98FyetEtCn
XAROFbgNqCtVkMK3pYF8x+m9AK7zEuN2Nd2WG5Pggdw72hYq6Wy7e0qInbkw7Ye5
8vHwM/0DK1E0opa7qreQU1jEpUwUbMnM/wT/loUNRfNEmIk9vgjnK9puupy+5WT3
zxzCsIX+8a7D1pXsNqrg/mEB7wnIKWfjkM3RZ+b3xJAhxu+DIluPt6pTH+ddq9uH
ueWqBiJ/Z3HV5C6ZDI8vq5BeeFipjBPO/dPWPLggkeWw5FiH8QESEaICYMoZXdBU
iNUQ71E33DpZxg3ZZYHlk8xUaLbefYVxNbZ7DUOVFVO9f8Yk0PPzxZzfENi/A31D
ga+MU1vsL8f3x8/4aJA72psk4yQc7WdavX8IpXmh7/irDTNcSedLwF2lXP1yYKf7
xDZ3Li09Y+4qTIJcH3bEz6TtX5G4aOCtaQs1wA2TIZZ/Whb+MLwQOmZylrLqmkrE
UZ25uP63GE8t5CmKk5LcEffAwdujD7VOc3+x/YUaFoMV4IHajeE6l9LoJgm8X7c8
wc7FyEhFr7xZpQNBttJd93aUg91k/gn/39a4k79dSka9OrKAPeYOGb5fO6zOzycP
x86I3gFbG2cw3/nbffwrpmauDXUOHxAn3uhx5MI5aVrcjb3QShsOeF9R4WIuWgQU
NviPwSTShHbe7Xer9b47E2KxKrLyVvkf9SqkWGjIx15+lPwvoR8XDTIwghkWisL4
/jXA6jyJixZ0K/DcKBzH9d9z1Uh/ccGnx1MDoZiOPcIDd/9g/nK+Y43GADn8GHho
fAhkC+m61cCBLgRlY+2ItJdfUf/+loI29Qgen+vtAZnAA+CTeBlbYSIu27O2N1z4
+g08gYk8+mi8s7ys5i1wX1Gsc4n2BggmF1fuZExvKbmcUaBK7Fq5wwiA9g+0vpVg
O5mfj/u6QvFEWDuKov9tYGxWX1k1e0DD24tmLlZ61ykcnjPxhyl9TiU2zL8F1fKa
66iDC61vUpn4qgMCaKt/NH/gk2ubm3gzPJ6QZ5wclE1lIk07Z/1prPA8+k2t8siI
r/NMbckzT6dsBxPNSAINvIwAGQSMLY1H4VWZpmR/wohvbfwulfgOS9caO3IC/zIs
fQNQylzxp6yXdrVxfRZ9hLYIsY/QLfstcAKdR40WXLK9Je+F1jpMXXeirG8EATDf
+ohSBP4BuQJ1zL5OVn7Fe0tmaOZF6CY/dvjKJPqbqSSoE6Dr1pRLBBQ5rKohcC28
Ode/YyrMV46BN61nnzxgfNk9Uqlgs8mK4sk7yT4v1zvSmVL3WwLVqNHW/bG55u5c
22cCpxsfm34pGPG6GPIUcUAizTScJ/B67LkQzgx8uCjqoA2ZXwt41Q2OHPqk/bYI
Le2+FXcE6pEYewf/zXhH68q76hFLYRDuks+zKhZiCWOwMErwf1SzCA103KPxr2AV
vXn8SCy+oe0IPRE364vFTYLrDe0KLiRF4yAWkrdlJAZ2iP5ROvX/NxMqic/ZgYRO
7Rp7jcOFLyq4YfNxAmgnaHOlBOa5C2UYICKZlg6WtoVLs1vjQc6UNS9BGsfCUnAq
O2sNpHAqwIhEcpY51eBS8Rn6CPZtrr2JnYOKciKp4kvCQPUtpJzybq5USaAIQc2O
wDlg+zl9WoI8o4aVNo/eUG8CW6E1jxt/4QkfIgHqykZ5VN+tc7FkHDgFLWyeF5fU
5vbkylb6CG2KB5rAC8WLWEugAAr10A6Sm6nFhpPZkYGh8wbEqYif5J7CUynEsu+R
NrujCPsbqSN6RGGi+WxZ6VeWetlC3CLQ78wnP7WKYxT82SwNUpLR0w4ao2I0Hbme
B/Zc7QUFSeTjD7vH3OQ6qRWDIfgkXLnNlnmjK1btuhE1Rpi8To/7hzke0r/WIZSh
FmvWei0MPi5t3BRI1chDZfybZps1C/dV7iHZJJtG8Xwb7MHxgz+ksUjpWvq79XfB
YabHgIQazzIpXIw87xjBS+jZ+S1zS+GTke48sK25MsDwwY0EQaIxDAxFuP8q9NxR
oZ6Gpd7SjwU5KaNUBWgqKXp+up4T7ikcTsyiSXds6EXLvop2e5TZSkBNYtDm9YCI
koCJD7/CrKgOwM+ycy4k015QXbBC8XqL/Qu8HcWM+6MJcwvKDpbtfLzqZOv1W+4f
NXSvPYuiRH1Hu4MVlVY5di+XhYkuE/JvKhr+CiI4CgmfRmNMRuFQyRpF4REX+y0S
qAZmbZ3UwEWLOmhiOz/muiIS3zdN0aUW1b+PkBQG9hRPnxh3C4wcv7KujWfqJjqo
jVnsXTQ0cwWAgtN8e+onbYz/Gb32aZVP3Axtnumk3iTJGrngg9gx2GgEgJ/lDd0d
ZK3Bb7nxxqz5YVKZhbB4xmUFCHYeqnrmZSvKfEYL2dGNv20PKlgkLdTbCweJp5iR
8569b1Ws8UlBA1oeMzcdmj1cM/LsQ8mV6mRlFMVe7bnzppC2VjR7uQOJ0jZnUvoo
b6lrFCPHTJ0dWa6n7LdT70LtChNvKN0raYkofJCfGPuvwLSrWOYgjyEhn5Tqw7n3
fcItv/ohBIRZB5Rub00eUZ3t+tJ0s3zbEDPd7P22CmZZBdHFekIAeN+WpYbCLIKx
zD2oLb9a86CwrJE4FhQjBhPVe7+ykOaEx7k2LAL22f8JYDsthaz15SJk+T1LCHHI
Jmdu0BIj7EAVedKCJphOStPeLFfzu9ETkliaYyHCZSCKf1mlXW7NLV/T+LhTJfW4
lDHLxQLx08SlpYFUy+PMjGWx5TaIwaaF7McsytBPsO0JgZGdhHzXkgMGlTJaSP6u
PzAe7CfHUZ4gJXi9IzJLjfQ4FJ2AI1WcljqNIbZfDODE4EHb2rJemIFqd06I4m65
JeGESC5Ib8nB5lB5df1mjbiN9ocBPKxqFtL5POj7UO/PB3naDiLnLEjS0OykIZk6
fESAAe8I3xG5+cO89e5sUFK6b66K6/3Dl66FwVvDzIRvb1dKuKjjiIzklhn52hja
DQ7NDPrm9vM4IJS00O+LgQg36fmorYAl8GxeA5jrtNWr6vERwMngaDP6HUUsq0e6
fLaIllcB1ljCrZi4fhuGcVS/ek1STz4/l1eZguPEgfWW1tasjDHVrw1YIz5SyZ8d
L+jb6QmTZ3zcrcfU1qluAR47JJ16xhB7j5PqG7c7/QTR4vvgaP3yGGK6DkDmpAjs
mZ21S5JeoKiwAONbhHWrs36RS1ZomC4wDsrKeq9GYcEaLCRibgd8c55WcrngyjNc
hI40ra5QAgV6N/9Bp6zb3kZl9ToXHnezWhIDJMMcFQz4hOZnkDiA2PZgfWpH0dm2
nuAPz/M7Mk1BmYYn/vdc6SokCdg9Mdz/xd/bvlMy7yjt+ZQ+05jHeXNF1ZCQVOvM
Z9a4PKxz4F5TgLLSBhhi2A/KtvmvJWBXoX3Gk0H7q0SwXGQ1b1fw5xeeR6qqd5fV
vpo4zn5DBYn9I2CtxU2UHfiguVH4MGIQyyRRGzu+BgAqxJJxPjndY0DD7IiTPHdE
M7l8jXqyzqFl+VIEJnmQklzAzkMLaD0ajN/rnWMB/WQzDWrrgQ70wK3g5gBQb212
Hjclosqk/yHn9v8+hukx6P/lMRWnUy1OmjZw3K4D0bxgPwitxRhnXgcskD+laDjW
xMybTuKgxeNvWLbsvI1yUQ1PKcNUfBy8ovXH3EuJEEvo4xosFIX9F2e7wTiJnKyz
2rUbDTAgWSTODwnzhbGi67bVX1cp7yf4hsG9n1RDR3S4g2QecJV19gn9tbl7PX3p
gQ9TlKFgbPaFFmr4YqhHnEAMSBbteRMeahf6pCudVM4SPsDdTZceBP1IyklCWbRW
e6nqxGit2UoL9RngvaLi0uHhymOSZSGlUX8Lr3ZUyiah9w33pvzrSAg1pC7IyfhF
ivHcr59dxy+JpWCTk3fi00vYquPgMPk3TNM/eey2LjJ7mAQiuWX1xwNj3rpP3SAH
QXIjxI+LRjk9M5iPaKb3jQ6+56iCXJ7Bikl0oDNBHz2pCXReyJG1tFsnkLq/akys
HxvmNnDiEBpFBJAq3ovadIKxU+4h241BQ74Km8rUhCUX/0VJdILwvsyn48wJV6aZ
us/3cEgwnvOA8rnJMxeKVan2Tu7W2W6z8adoPiFHvygt3TFvecp5fwHTfhPhlfBk
GhluLLKQeZrM6sHyQbzFh+lpqjIXqUYB06mEt6sFciaxmfjFnoT08f/CqcAnIWl2
2tfgOPGinE0uaF3uM4L+7eWHEynLG6VqbT3HLmMCMYgqs+vyN7rKt76RSmGQYTq7
MGf8+QeWKz5DoJJOLEVEb/0YWnhTmE/5j0GMFfoP8NpUIspe4N4hnSbKhvYvrcwu
vvKLfizZc4RyP+7I10BN85qudclKnFbgBQ6ArpVaReBG1k0aR5ZRoypk8JT9QTVv
TZmiL6L3DwKjlHUgUXYkqu6RBxs9O/e3MChISz/e6BPDhBpkGoEx24oZVH5avXuB
kiWx/+K8lDoykXO7N5wdOrkx+UIiVjKOaitt7cv77hqinxO/8ZRx5aygqEqhtS5Z
LVyvL82sSIraKctiNUVElrMAkaar3Lhr0W80dqFy/oIPP6Ak9NeN/m8afxCmQ/wV
f983+UxbQDIHDI9p7mdWYfVKS2Ex3tUJZEVrIrCZ9qQdb5ENb4STuSxst/0EWWnr
sMgsrG37RWX8drr+Sgbl25W9TKVasFsRTyT5AwbLhSPD/Db0+WJox8jQiqU1axGI
7ZvPLYlTJ5fyaezdL4Y0ICSz6+9jL5yI8VauDiUEQe+RZYEmCdaJhEjw45DfdkZ7
buMygyNLKfBZC2iymyOZlwQ/+U2tRJR6Tv7/QHdLiQpif1exPct3PCGzFLrfzw1V
bdcworHyNlrgdIOzSCmatHA+vpgrcinAJlrWFQKQx3vJEZ3ja8xlF4oYL2b8+nS0
CTR23I0Gr9UHQ3DF1AvFL9VzR/CPT8H+vMBzej2d5DTnon0o8lxGMdN7+xjz678V
yQ0tGw/FFxvR5fCMu8EBCSXM8BmdIlSMnmalCXmdeDBmAZUF144RrXOQKNKWe7wo
FHnkxQtxvGqpPS2+WrGjK6Ns3PkVfhKBpabWgWb08wrr+scXO2m9SioP6AmtnTcK
AYCWv5cNuiBA9T5WeSb+14AjQPfs6OWrUiej2DNB5MW5IkrZRj0fde+ZKGHqxWjS
ZttXLbzUW8N0LT/KxErw/zEsj5IogM70iWwVm91+C/mXiWUKR9KEDx+pJGoV8dwO
iLn2TSauENuthi5FhQUr7mjv/pukAQhhuo28IdaZUoBHIDX0wzwGMcZJSR4x2Yym
xJskEKap1Outa6Br2gQ+9H4dGk4+owTrc8S/YOHqkRAPXV5704lMtM57jIxoCLtP
9zaFwBZrKpsMyYzpUohEYZsIp0HzCK5uFAc+x5YOD+6RWBEHTssYRzaTnbpL/6Ui
FZ78YhtkJuEZ8VbOjJ523AbQTJGZWX0c5/6QcZGiM1PUEaKq9pY+nFXqCs9Ix3+Z
bykGoYxkGHHLYJjsdZqqCmITrd8A1IemFkwCZTQvwlxl+drJ/4g57+w5HmOSE5iO
s/u72VixJbhs8d2SpalE0KlRG96peQb5zUpdTTpZtjBI25wnbdtE8F16+3CmxNlb
SemGHa5jjy8KvL0WbNKgv/FAWSSA6TMcWSfpGxet8d3l4G0/vxHCGQnp/HlA/qpy
ko3a4OCmSu01TOSPbr6ZJuPZawrarVSFaK+FY2bvbKpPmst9wxYVrp1oUF2aK6uC
hIOBMJa9DCFesHSVYY2xReLir1+i3qrvyCralNSMeMDTmCJzH7ne5DTCMppIBTBp
Fq6elVXU573tvHo82fjnB47+mh1BFemWuwDzsNTFMUe8d+t2hxZzaq9WhSUt+vij
Jq/DwAUFXzYOCTRvWZejW+zGS/OxgwjFuPy4aa9XY51pMpKliuqNRO1oCKFFOMDF
drDPZkW9qZjnwZR/wApFwhfzv0MdK+r8Pkp5y9zT2VVE/SxctdijqdDGHrD/V6dP
QKSTTeaxwP1b+3Hnn3UPNyvPt9oQeUxMowWjktI3Czh5YXw1o3qWnTjzRpCBxvgg
M+CStrnLuGIV0Hqm374DeieQQxSdSQsKtYtjCfYcRG6ifjw+dOZNtjv3t1Pk3saN
1wDfe6tDMXTNwQXC5IbiMhAVmGM6SU0YaGxrMSf0Jzd+L+ZWx5Xr7YyqWe0acVyb
ce15LSqFa+3cDu/5dAZrb7Ol8Vuvt2PB25XGVSV+2CTMTaPyZ7cp1Z6vghXsEngl
BV7X92ntmUAZYBkpihi0Kq40cktnKK7fsm6+YWvJV4E7Q8S0PqZc/ID4Ut2RUmcS
Kd7OBU0QwcG20U39sntWnX1MRvgG49jftWjUu6QuwftVTZC3nkILtYezFaz73LeI
zMxKb3+RZTHRujyorwXp4Q4YLnJ6dQTTERQ5NQtlnsjulfqGmTv2QN3HCHh7E9Lg
g93m+j5qanmLySkcomqJz3FnGvRXCf1pjYHXSvGshyTwzpHyhwpj6Fao0hUMtByv
pL5EqpBp4Gxvl6r2JGqN8MDVa4mAW+BKQKgSqDIBfVswrdXrHOG302+MrsJda/90
x4TKB4TBA3g+++RnaeSRFELaCZzCb7OkjnPOnBQCQC+Xt8d5EJSTNaJMZWNxntja
XTamTvTO+RM+tjtJDz9QhUNHo4r8EJLWkl7kRFIoaUKlDbULZSZ4pD6/CVV7Kwsi
bafK1TGoMTU9pWu/SRXEkpjuc0NBYoYQ4iyKQKMvQ37lzZDWoo+VYs0Bblbv4CLg
N6IMjEq5zmvARL6P0rbXujs5pLaje+C6j39pzkWnon4SZvY+SN2JUb0SnUB9y/86
Q/eYr3Y9OD8Ora5gqXUbxm6KAi2bp28+sWUrfr9L59Ced4oxjTxqmt5ewUBODlaF
B+bJVI95wI7uxTP+iqMRrkY1LQiJDCssVmHWbY4TGBarTKhVxXFlZWBbNn0et2GW
LdDvtgEd2LVf5pnxJWPLU7B+aHQkb83qcS+9s4dWEUhae/+Ct6Y45MoGGlQGly0n
xMTZSpqJ8uUi5bIa0qWBbrTXYsLUt6t5NgP0mgpPpojLIWRBK9KcawXFrLd4oe4+
0u0r/Cw2N4+ndw/P4rZz9DaFng8ywI2/JtIFIQn1G7/6o3g67S0Mma4+S6Z5gvOE
DSwkcf6Gh/oyTwnu6yXaOKu9XL8+rArJ4tcSuCSUxVLs2CdStbA8l+zGnW9+rGX5
O3yv1jcZyVoWaFd5ng+JziQEUPEvoqnIG0rb+BQ6p+E8ju0jPlJ0wtVhE1oczF4x
8aQRuEkx1xwJsm4Oh72IpZavqI8ITFWsnIAMCD7LXNzw+vVYGD6RuHa856LJQ8KJ
yvtWj0+Mo2J4b+oO50LtJxJwIOx/EbMVRr3A6uWnX1iNdyOP+cbcb6BmWnYqP8YP
YoIQIG/vj9q9qyCrf2Eg6bgfFdbisUsuCnr/rcmXj4vlZX+g20Dk8zmq+22Q1URi
WhRJrBzvMysu91+KJhJdES4WM6ftu0EbIMChT5EVUzXbw0fVNADDteAj18T7H83u
XyhbFti1GqQpM9DG0qmmFooGxZYYWSbVTkESvlzdS2ktAJF4h7HShfiu6MNmgMBI
MlYAgYSU+u7zbL4xInrCKMfp4Hz2hpxYgyLbDRly2zdMjy3x1dSCyFDPH8+O3TFR
L4LOmTenoTjuTgd/+Hsy7Zin4ywaQyY62LkADq/cqYks0y/1f0PWtvg7f+1KwXfG
Jo/n/10qmoMpdCCeg9WOQRV2pNRaTor/Oiw22r5pYui3Kt/IPbohRsIQCue6i2vt
nVKoWik8NsuL6bn1tFvRHwyxGSznefxRCz0bLDsGlb5Qu59RAi6XcVhcLFS3xBmW
DWZtoIRi5PhPOwJySy1SvtlwcVJDK0DjeENgBHBWgyZtja4h+mb8kaRv5pJEiX1G
k3l5HqsYqN9b5AJyONILKV5YSXRrPh2VL2M6roy34jL4Cx4ftjLTTS04zVvw54QH
JhXv2AaxkgyznWdQtMZBAZzdqSZXlFGzoM9bbYszdQ0Z01++crU4Kk/IS7JyCsez
9q6saf+RM9TXiaoQVuFuAM5bDjJB0dI0wUcq5v1Hoo0J+J9yQsF4Qghj67sAXuS3
E895lbdgw9jFYzdU6hrvFxJiOp6rNW+qaQ2lYkCHVG5jkP/ACH3uW6IEqbVNn1B1
YYB5Abnb6owmX0RhKUrzMCWK8lL3RQg5W4+lqX7edk/DrdMDgMVJEYnQpcow/3kp
xI/tO47OGvwRbdftlPxgsBExhyXcLL/F6zqNjZCiILWqlADjRtV4BzVy0JqF42bP
LVkje7AGz6YCJMU6Efz7HAVipoXLQ0xbNcjfFct238Eb96pwCsMr8YIYmqPtJdtE
lW+e/OaB9V9ODdPQC/KI6DOBFDGwRRwco6jQkIGnqc8/G4Z59ADHq17zBz/TQRux
+1nDwODjWblIbQhzM8BO7zLQPRsjGzxl/r0UK61ceCE7EvcHE2GMYB8X6xgeoEtg
poHpP/3xBEOmrh8xXNRdXI4Xss1edao/kpYZE6ol20kcPr+ioWvag0Rmv29vqkXF
lMteKsUojyYhAlUS1jDlbIY0T/DAj3cSaRv9mh6pQq8adXEHbpTlv0fnqEw0JO6Z
Yj9cA9khJmaiYtVmgDqJ9MOjDPh9Qyo6KRZm3cZ21nw6zqb5lIOBWr95/QCNVVow
nB2x5oey17/y2uHRkwCKn76RD8jPEPQ61VYnf8tHd19EH4vpJZJBZ2oDxn//kuJM
FRyRiDVo8RyHSDfgXkjf4meAFgEPzG4VGMru5LAOgW9jzfwGXWT1HXpbVENfmE8L
tGaLrls2ra1yUixDWd6Q1LrGLe9c51wrGaUOMHudmZmKWMd9FBWcU5MZh8gzKB8q
mBaNJIUF5xn5nbd10CkKuwxBsBxzBX0VdFYnUCc1o85EkybU1x/Emqhj3RjO8H9x
UpLcZ1iaBMkU8r53zsqd3YjzgExK70396LjeZsVmmnKjmScntVT/MlrHK4PRyZpH
5MRKXs7AN53y6tKNy5Gqj9qe39OVYhlksatN5bdkiqUF6AjzW/aJIuFEtSjug2oy
2no7slu8uns6saXAfs6TFvAi/4Fa4VZS3aLYfDbWxmXgH2slvO8mI84QBE9IMNwj
shqlAQeAKw80aBYoxCVRhk/yN5EPGYn9VGEVVLiyzF7gZb2Dpr+3seQ2oqkpiEjB
tMW+vEfV3MlbrXkBte1/hDTp2QQr1V9Js6fVuKvWK2oDxooqg1e23XAf1IEcacDk
SESzxaR61s0+sgAHgqXbsG5b03Crl+ZNNiz5/s8dm/mKscoOZGlqKM5MQkzGWY8u
9gaAs0hDjRBNG3CuiirhIbpPh4uwSJNPRra08eATLnaZWvHw2b+2KoWhAGEGjbWR
Xg31gWBm31LxzXwPqLr8jYptI+ujfIvdati+OJErmqM2wiU4hEnF7x1eniHIGaX6
epWKt1Z9s47p63WyQenTelFuDVioLF15/c0vLqFnOCElikaJRvN+Ixjaim92DuSZ
kQtNMDL25ArAShpU2k8MSqA9ipErOCh+kjqeObJS8HKqp+oepCxhS2LCKBmmxeXI
C0JS3cjJ9VdL24vaRA6/Rf5SGkoomPxS8k4h5PT00zbkWDX71lqTnhDn9TgWjZTa
x6jQ1wSpPanlCFaL+H0Lo/tSG2uQ3L4SkJdKccZffOu07qOnVddFFvRtD79qZal9
xVJL4Ltm/9bk3IjjgFu4BI4Gyv2XJKpl+PkDFB+2tbmnsvAZZl6+iPjDRJ6fNKFt
fbwK/XnLyJXFyeQyuVrLfeEUURglSs441eeusgJbONBorUBOHCvrHD9xlHie0/tt
kbkus+U4heptw/Edvw1TYYXGDULEEGkHywvBvqS/6615Qc9QSPID+FJ1zL0x1d8y
sL5Ob1EZi+rZLCUSSoEcUgMX5WNidOaFt8teSw9UaU0YaDWHY4kfq5CZtqBeGjjV
DPW9hCWMMAT5yaqZjMKRt+1n3puekNHqo0/rlM/GSWQucUf4dGYIj4JRkLWOKAv7
a7Ir7wjRUrXEQxbai+mjrgvG4HNzOJmJ3IDti7J6tvvUU9ltFy/JhTkdO+HkHhGn
uat0axkP9u1QQYjv/YY3+x9ZYJ9dRTIwwdgiB05AfvYNzA6UlDGfdU8j2E7fMe5t
h5WtJ3z5VThv6yQkMEAG/Dwh67N7jZWB1QqJ5D77MD7L+LUnTTiI0Sb+Y3dW/21E
TmCiwaCzahUokuSXDJrgn/K95WSaFO50xvzeS1SL14Z4ligNakz3LqZo8UJwtjf2
W0JzOcDwrZOkHi4Zem8XxZX45zMX21lELAUHHWOlBXeQydZYLtUUUTIzYYk84Y3X
U/bpmU6az41/oAvopjE0KE4fv+GioanfO169esVCAgewcU5bRRFuuExbQV3lalFl
juWEEBd/przKz3oYla/NQPx+j1q/HnBPnM5pS2+hnl3vUUaqA1gSPnqgqt6QLwRE
jfWk9BSlMRtOPST2whi/7WMBijWuBojwwUtw3MSxP/HTHzdIpppQp507Es5eiYwb
uUIjdeDknqsiSKFibyQ/ysP2LRogua/2XpbvnDlfFPHhpp08Kz9SwA+gci74FM7g
tv/JDFcnUb9WPpcOS4XRe+lRJHnMHCaYk50IpmEUS7m9ly9j72tkgURSNX1guEWM
OisDDHbuc4pCNvxIh+EMWCCvkIaOcKjSRw0K/C8G61/KRzVHeUs6jMat7shfYXnn
4/L5CciWMnV5wHgacipGetTrZKx+gz3JDfexkQ3TbE5uxmkn2FqPI/M9WX+BdbNn
fppfyqPP/1Ks5NEmoIaNA+IYKUOAI73Ou2M1qw0M7APWPgYKNbdokwRKrlF9vQUw
nf94BhrljESSHv4LgrXfzx6e1g21Ao+MoqPkN8/xMgyYxSVFb8ngHqAJnFvKBIxz
Js2YemvZhZ0W/TmWif9/xjGQ4c4gHgOmYAXfqo+XlGGz71E9qTeTYmj74ndLLW1C
Oz21PpYtOS+HrHfiVMA0itev8+PeDgtl0PCUpMkF3CqNeRyGNHLMSg1HuOubMlwJ
l42gV1VC2/+BbjwoYZBuMBiThqRcluzO6mHa8DtGR4nXQBEHvBxXwxZ/HALUkuru
r6zSl+ighnRp6+SlHf/LuhuoPOalcbNP77CKR1kTCFAmJPd2hoTI7IIyk25DHhCh
wtW/nYwplDzpeGrr7ri7foxy6L/qbynCCMoP6I5tltu+1FbeWIrXwd3CgBhRlx5W
Af1G1o8y7mdO3OV6HLT1IedPI9sUhIo5EgxUqLS3NL2LHyL73MTzF6NrO6WzSUMh
8h3PAiowxsR8vpLb9vHCbiWdMFIwJyG52N9EBXI7t3wZZTgyomI3b0Kz2VDYnT0j
3rIH+iOAVFYikrDuK9zKbqVT9jfq3FdJ58ATiaFdXLQ6jFC02mgRwPN1iE+eCT6g
OHmOSgFJ4I9wn8dix0YNIQU1Hx2DMYXfC5+3R88j3Psy8aeAfrmuXB90+kL5KCwO
oDrbW5QtjDuFOXMCVQm32pAulE+Pe8gwYHkiSbp20mOJHAIJc+7Rt82Jnt1uf2Gb
pNoNvrC55alaKPd9OVX/YlYCPN0d/SjLHg+5WCxIsWIWsD5qIdADXAxiU2gVcs5W
I69VBCCSBhdenqaRRHpPNTzAcC8mjDt+JhNYiqj+zJZmHAGAWBvGZmmRou2mfch2
V2/1fmYL97tA9+A++6hygAexc65lMXfPa907QYnmOxn306Mr/PfQJWKvvMXIisow
1spkdPgnRO6IRe8taXuI8chEfBydX9Ty9ywRTulJ2u+RoQQK3qvLQYHVc911UlA0
MvGR/4S9iorhLu3WRDIXjUWpYBVMaLLQUxtO4WYHg1YbmWrkooeWP0oZyRU0NSZm
QRUduZF5raXq0J2QfachCMwERzQ7qb00H4ivb1YpPLzh7BnnKM05EzSxtrkmTeRZ
+K8/W9kCfKyAcrQ8cmFkuKSAQJQy0yaGXB7oUhvpXwzW5qNF8hNRKj+5JVVezVyX
YGJdSYNiLv78Hadcg0ulng1P+zdaTPtwP5bgb54vg7ydr6U/urtmq5GjAK51owVc
aqHI2Tj4myP+6959NVA6SCOVgrk+ytunJKmkoZNKvl/efsUn3HIkGeeipCIrXv+m
PsMKJnMgQ86mtbW8zrydphragXtslWL51p+q1QPt2jmuyoWP47GgWYWaD/Iwi8AJ
+9HrMwKGrbPbFXIkTTA5N3tMl7VyN9lYirZj/3sEYEQq6lnWr1gk9ZTFmOhhElr/
bHTHfeJ4ttHZC5nqaeItdyEwBqYJcm0nBLmbP5Py0jQiY2Dqc4tfVOnLM+dJ/deO
S0jQ9PAuVZxO+1Lgfnc1UXdcpRJufzE0JS23gdUfHfrzzwZEmVFyQvr8ZG92883m
GQkwhfP4Bgg4QYdEUlInByb7uqatVa8DUhdckFVpwpj31Zr7cuUsEvuOL2CkXLpg
kuzB2IRERHiwRKH4l1D3SgVV2vdocmiwywvmxvpUZyhE/5tJOgCB7IroJuXepT7I
jYFeyWlWQwIvysVFMKmNKXK92y9Vke6FIHqxrJ+UgUbi4PpMihbhz5l3b+TcSDNY
HS0Fkk0kMwVrfd0GHLjm1tjOI/2GScg2UDFWxPdnYF2y0H8Rb6e9GAODoxI259oX
LRhagpzU4jrkwnHBAo+Sw7I3A5RzbyvQDJtZ4Dw2PrjIGNON8EH5l1xzKEtg6jdo
aummZs3R1tDLhU6Lw5kBlXBfZfPoV3obkH6ghxxO2McIdZZp3LcdaI2LGzwRuLa8
jUR1XTROvrhCMfjafDsK48j/2uEi1aLZgxPNo6TdR949uPVNi5oeMTaAIfNiv4uQ
JmIpolFeqPPFM0NKAt9Mk7UcRZkOwtUqP9ZCnYcxmKfYyBQL1RMZhuOnOijIzUuG
X9MX57qa3sHfjsMHUSQyxGdiY8TU2Lz4sSaYgLMBbPR5RJVl62VglBXjZDFZiCS/
R6XjJYLMXUBVdIuNmbfdXAJ0gAgwf0Us11Ggv4/rjfBOq5sdLp19di93S3PuAbBG
xozSVQChaqk/2/lzmD3koavZcMbxOv7NdsG1aW6pZLjkbKGIS6FdObz06AF5Wcjt
5q0VtYKtwbwsePGetXfoZw8OQ0wx79Ljfs853b6CC05zge5J0zUsHCI/g3dj7QWy
NRMexlawJ0nUnG5LmkRZgn6NpxKTXRtRNAUnDKVSJZ3EONudCG/JACRZPpRzJQNh
7/ojYQ9MHhZm66G7Gp1uIsxfHRVAt23Fw2jYsMidX/uc2xCv+nN2ngjbR+xM8REk
tEC95lOTiAB6vhccIVy6V1vhpFtn3wyMfvrnSjgAK+UR3xL7RP8sKG1AuCQR9683
Vk/uQqYduT1NKWAuIth5O7aTdsBB++Rnz8Mo+azpheG5jAm3tj+pbG7Ynasw2UXi
Zwz1IRDh8mZY0Ne9ga14Mn1Iwry60CxXTeJcNCNilUZX/g7dfsGw3ABi0Nat0lFR
aLOqswdtWiZAwewH1K/BgRl//PA6kHQE+9zhCVy9qKJoUOycB+5EAVKz6kpbAGgY
yPyIoNBPq3vS944cZn5c0sl/NB0SU5OAHPkAx0mc5vwll3QRphcXRndIUZg26Qdu
nXftOwFouXtNfmMbemIEIr+jjKN53LW2vCkQKdgWSaH+wFbb3T/DuMnUFgxdv21d
5JYGZ9PelLDb0Uaz4Ugr8T2L6nwIbqCYhFStwOcG7v9BcoQ5wA/Irp5o3yJq+n0Y
9GLh+kWpCiLXTCjVHVtVk0J7UMtwm0mxKQhk94z4QoQ=
`pragma protect end_protected
