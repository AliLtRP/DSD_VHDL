// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VDkUviuklo+VqDmL+eT+D3RfEubWBUrtw3nC9NWO5g5npon1X5K8LxdO5Op9Rjj1
yLt4F/FzO2l3NweRf6qRGqwGPD2LL9jYEc1N4c4f3QAXk6VUIDA+cyvxDj+nD09Q
KgKwSs5HzxivRjuosvuSqr5hnd0QJWG82EB0ofGCkd0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42960)
n1+hVGP32pUPAMI6w5Ey5siGIW7Ecc1H0+HsHDljOIxXaoM2iW7bPklsMkokHEgZ
YMxG5ABLcI0AycwkKInSkP1aZxUiKZB8dwMBlyUeFoIkG+b8WL4F7mOSyH6ELVLg
QVTpVjt+aW8Z7krWktVf4qRk4r3cnh42I5y4EEwOWVStN0XWWjqNDDokwVkLEvZ4
lUKFOjJub2nsKWDZ/Wfzh1SDnQBJKRBz0nLieE2oysrcL+Oqu70SSNmcLJfeo5ap
m/SmsO14ptcM2aJuVZ5qaV4/PaPE5jwOBlctr3XsIYREeOhLbRBYIU2Y8s3yxfHd
+DztwGMm+dI2Bs/hgEmYgiqNdHnKyf/IVPZYkicYmeEK1skT4pWWX8XxmFNQA6PS
AK751sZvh/xjDcTZV1VgWMedOvFQAUt6RJ+zxrtqyya14zeDxj5ahCh36t3nhARG
ytQRJ3VnKeBE4qVuzGEgfRF3yXneuZiIFpdlrjMFcq+bzwrzKQKClrrCTcFlmf9K
9sUnvvOdMyRD0LPnoyN3FaXUeV1fffG25fYZ4IgzI1/9qllYupZPyaSdv7WDEhT5
kr9Tbj7Ca81x4vjP4czcHT9f56vH2hOt7FkxeiR3YCyqZDyC7JsOKaxZ9MWzTSfP
88Y5uujheM5koUn2w4Efhl1BzNafsrfacqiHras4Q8uhnxECPxePP5Uj9Ba14Ult
9evYTjzB3/G2F/iWpebnfSWmRfilLKUBgH8CMKWzIFtKQxVbMKdS9SqGpHOQeKu1
pkQCqf94hTXTeqZuyK5ZXix6FI5z6ysYjhW2aPhC4WnOApxFpIgHmPr2Cu3IbNS2
XPkWmpmUwPI3wzqksVZTVcmSKUbLrX3oEXDluC4ye5MER00R/YJy6WP/tZ/fOQDl
TPP8jG41sOHnpa3yUO6nYWeQjKRx1bpM84RAePGx2fsUs+176u2yACP7Woew8OT6
fRSTskdmy7BnM1nHDbFri/JgTraYBV+Jyk8Bm48mUQzTcE1HfsBn7iuXO8vMLF6i
ORJM5yWw/7fxbZM7B+GZSobDtfPHfiG8yixTPA4nBXY3b711o+cTCZ3+HnANAisl
Dq4/RXqIkvks9Z+tgYjke72Tvogh/u3rXWzkR7lBewhpprGHcGaIwlCZEvHM7TvK
RIznxczzkynCPMeFts/l65IXa02G8WqI7HiT5UwOoaS3edKlK/d+e3Q/fa8y8Xjx
Q3t4oXGZRyGGpjvz8/usskg/DXOIvvFP/hZZb6SlOKzB1Kajy1tKaFlC8ek9FZzH
4euBy/aPTEX0a0Z0XFZKMPQSPy9fif+J7NvUrYxTUKncdkKn2ytL+v95BoIjPkC2
nXkY8WAhpB2W9Y1uC+pPxIumSnElhzX3ODVsnUJaHFiaalC9lYnYLltyIu2Ayb5x
cAAuya6RfuBAPZqpoqnBzLqisQQRbwY4+kasS9r7bv0dUYr+KSuFTQ4E49fZfREa
IVvDkd/OQoWSgsI9JlL1sU18dfb/Lp7yX5pgZSAreu7G28BkO01P4/4c/2eZvJ5t
22y/EQUB9rUFgpiHk3XgYpBUVbDptbFQSJr4wGOyCEIV1Wc8tpfy8tLMDZiyNT0y
2CltUTYDmNGz5EABd+aEbOcG8Miq3Y62qTuAgl1j/mQ6PigBimYdIdUevz0NJVmH
3V1AY31So+Z60ziDv5L9AYNxzt7DPDKmxxiuLJ/plFQMcKksQ2jYkvWfEyc9OoME
yjcAQAki0nn+RACaZpVNWa4HRy30BR+In2g2AXVHgZ53/8d5x36QryVlkM5iE0uy
uHZyL18zDQMCRqEjdc+PblT4Csnt9zbTiUmTqrBn6hU5DYJIgm4pOr4kMtb9eg1K
CLWbH+bowwuu/Djte0dYN7ex98DjUf3ggLD9WCGzveAWl1S+twcFJ0Pm0Z3God/z
/sc8sTZeold0/htQk056YJkKf2EBcvimc/gGTvY12m4kRO+NClMNCaptX8Z/1jmb
ghq0rbH/wci0OwyqIZfbOxlr8QggOGMrKQBrCr7qZFAGpFkeLLGHZtJkjoUJWMg8
ypceQFcpG8uaj4K+arfu3m1prU0JyL+tU+WlDlf0LONwDLV0XvfCMbNmV6cmqGA7
JfsiJlrui3NPOGvUwmPfNWLFsP8LsE9N0Rib0e77M5I6oLTQGOcjNLmr5cR/ByEt
rVPx0OB2tHzLtVANKO+R4gTOia5KM1CujdFvGdtml3DdszGECmJOnmz3AphCMhf1
cTWRMKJiGvP4oumHgnb5U/+kGSag6+EY0vTHbW06/LYpNKP86mXqz5DAFZLxoDnK
JDfRiXjt7re2wW7btC9ZhNuYg5tcFhtw7tDnQQkbd4YpKTvUIewvVE/4OAwC5qxe
bhl33XKZot+8wROV8fNlFXR6GrcTZGcAN9ncVwjUhr9jTF1k3Guk2GNCXPt9fprY
9MriMSZfs94GC13HROuu/HjM/1HeYI6c3yf1MGWKF3iMABATm7dCn0/G8ML6e8gl
Vyg9U26oYNWHXdgl4lY+AR/g27r6kntS8E2Iga6rod2OCrUwdUJQKDETzdn5twyT
8RRv39RNogaVPut33PUAp76nToWk1HDGebEEqG6G3TEYVRjeLFy5CCUt0UIc1zdu
rOSFpfiftsP+86ZYe/nZFqxeQd+6tZfLEx792BJd1Dn1v+9CwkT9Xox9s4LJvUXM
Rs9ffKI0WWuFiXUjFnVlEiYCf4YHgEv5prJSbAyiOJ1WT1974u9Z563/pL2SbZ4I
qo+7E51EB7GVoiUqdM4AwrD1x7qxB1Qv+6d8KmUfk/nX/rWoLuhDiSsJh7AuYSbW
gWnqzWSaCnvUMKh0bqKFSTxGVYrjaMIhyA/NmPQ3UnOJmbwvWFOSWpAbZ8LYxjId
29fKe57DMP20XBQtYqN7goaGu562GJf1697W27UXYoKrCOiBNkDUwmexV6tp8JDe
kyVfFQhGjTRrvcLoksE4vR9CQqKgDcUhoX0jALRYS3I1wcqbbAkimlEZuieVUNGN
HVSCkbZEcZF2/6j/N3m0pHoey4hnrm1GtPpYuhxGc73HSd28GdJd9pliAeUbl3ke
+YMTg35+xK6+czD/8tDa08gRonOzUfv/06I0e4YNQLAFUndxLG7Amg/I7VcgoGnq
EiuFq65x18bOzA+XlS5OK0Fd2GKixlN8meuj4BTu4Oep8BEHsySU/2e1sJRoYkBq
/xgai3xbhCMG3gV1auLzfSy1HJbjk1iTrNS7o+n44l96QUOuPcVsyrz0oTwDI0Ns
56wX2MnXkh99SSt8HT4RNDbBUk9SmLms2X8EO46VOHBuE0WO+jlvOZkjBOMheztB
o5Su5ORbLzDZdwUX9li6fO21q/hRQ6kTf0KW30HZMyXMoOnKY0kWreyXDgsbi/Cb
nV7DV1otOefdb2xMCcHE9Pp6/SpdCCRjtw8l/G0NiSUe7/fyN6CHB9Cng3kC396A
PjD84GaMSjj7JxzGRMOSNyQfTEVCY73iFjmWX3nkRp2QVsRzvnUbmLe0aW2a4WUW
fWhs6NqmIyt1IhlsbeHUHxMofVRNNyF90QrCvQSd5KO8TyX8eBjELjC6p0nuP4XZ
6PqhKTGBFpu6Xf9Ec+027v23GJPcMSY/+0xYOa8a8JssaKGBNmSJ30a6UfZpBCT4
NcY10AKstKOU1SPCR3dX++/IVCwW5pTqKJ3itVQgJ3SuwNnBeel3u2i6UtEFNgTQ
HHTYEn04o9i2yTQH+Q3KmHKVqN8x+kmIcrQ7Dle8mfyj+HqAsbxszphh4cuhfjfP
2MXjZ69HFn2D7HJcaGp4CYrfTeNEM3jfryQuGFrPn+FJDEmzg6XabVXIQOoNmeSY
DDL6Ic4QgYJnQa3n04bUuJ3AZcJUPJvfNKduAmMJu0Yhmu8r7a0ahdzlrwIC09es
y4Pb3vBjDlpoi7hxZSACNuJpFnfQ/yYMdYBq9vGYK9RD1qkHLUH66HhKCpgeO24o
o+mNWaNRBSso3mUx/fkL/E1kk13agxwzuVbqFbig+NH2H2CbiBZr7oyKLjPsfyWU
O30B9bf7FoqQOV3MPvC4KkJ0o6kK1ucjHts1yq2ympFSLINxuXyTga3UMe47GGhw
+m8tSSCBiNtKaJouipqtD8nyFgS96wUvJjdu+JmYPA/MD6gX3KLcTPfowi7HAYb5
5jPn5apjB9tw1SenKXhy+bq9EKGGatWB4rJiI24g0FUBk8vZcq7Jp574oi9ddiL0
SPgakoyl7rYwta2ryfnrW1BxZSUrze7ZDJCgKXTlLxvVVFNTp+1upDozsyEYghMx
xy8N48IzTfK8ibIhVO4kq3xeONo2IV2xygz0rtf996hC8iT5BqBXMO9ktXzqoWxk
8riBhtSw0aT8RbD4LXUFTMdU1JmR8JAqCtfdKchqGAZ6qCG/Q2zngc+4UohnOUt+
6DAhRT6N7HYfVBRIl6ahe1CAhootRlvYzmk3uInIycoddIhHeUJXGjNvSoH1bS6p
oZVpuKz4xcO38SA3a3PvL6l1JFaYhpFs5ffywhdvvfbdjXNVTOMK0LAmYtJVyzLA
UKADQ5CMHydscPonV4hO1NL8a6yA4LioK8Q7aabzFWYpm9eHrMMpVMmdfHaITphj
6SJsUaDPhdWAAtDSkj+WutMeHcX+zSJoqXt/7/0Pqf+KT+Yy6rsyfAXOQip/YLsn
4ywuFo1AkvudDYf2i4UT4p97Wy3owD5IIEi5arQGkGLFv0pFdZ2xEWH1HD1VbhJY
L4Q5cQkJ2mvePKOoWQiVIn9BiT9gngag+H2qnWQThLSVDgmPobEa5VUDw68dcH1p
h9cJpCn18iUupSK3FUlcr8T+kg3FCASV5BW6JMXcnvk7ZBb+riA52o90GkGVrjtS
JGOQGEkAqr0toV3aZZxix/cRWH4Y3nrJ95WeaQPoBCiZPL/N6NVjixUODOSdlUBA
sQ35WnbUTf1X+s5VsJ+nDfA9WusdCnW4OB3HTJZDkZYxDXkgfTBPUiX9anCdBgQd
wd0GEYjapad34O3WNbMqhxzCE2yJ4wTrmLbCNxQ7AlV56YEBjjxOaV4yTcdORgjR
PIIuDoWfwq/CWmk426LLOo6xR37y7VKv5hwpiXTyuD8xdadSfj6PlkTkgCr3DPiM
AhSg7s9K7RaXsbd/1na5bhMA4eQ/tkT3sPSOGeofVvEolvIxMsV/O5ejzy60lKCq
pmOjy/97bW0nyyRIqm14iAaI5GVeRHo5wtmTuRHdto7mmBzgB/brfsXUFTQb7xjA
TS0Fe6MbPTHcbxUBw4svFN5KMITbhPqJMY8FKKMwUP5z39h8nR+3+oUTh/d/NGCv
tsRWJEyd2pUhv93nb+zwpp8rtQ5jggRQQrQW6c0uikdWxq778OVjXqW3YGJF3XU0
YE5npFWRmL4nG54vzoCcA+M9w+l51E5zqwG3/ZUFgX6H6FJaE/kyVsmc4+LEFN/V
9TFRKYnusEHHM+VQKTDG8mkuU4IeoscQInCkmtLwesiQqKh11fO7UA7Xct+PN/gN
kkCoOMgIwvDxwmzSynB18Ww+omv6e1jmMAoq/+TQBcDTKCIg0vfB8ZHVv6qZ/gU8
v2d5tF94nsqz1dqNoD6aFGgcE+AwCzQD6+pfqVqrHt6a2IsxpPxtrOn4IuJP8Xng
jhdDyb/hvLpmeQkuwOLN0PCBooGDMtAM4Vt6wZm9FmwSIXm3A85YG2JvESExrMMI
WlxpVB59t7U714u6cP/TMWRMryf/rnUymT8Tw0cWdh3ixwfKb8snaS6wg8au4EwT
sFjCKWuemXAlSbT5CkTYOwzffvwq3wpbfBIhybhsF8mPY8Z6url3lcOOEqvROnEy
T8KPNd6k1CLKIVZQk9ZMnFA+C6EwbkfYy9Fs/8w+iCZkua3lOcPbWB+51RB76Qhk
esXWw9MsPMU8614XexEkqOGuwKH9nz6+qYZ70l5t1Njl0nlc75LDqtNeuznMddEe
frBmaD+dMZuRuBA1MepLnNptb7Sg4oM/aBbncHHoFqFbYAnb6+2d36w2Q79nFT8V
bPxJ15N+VM9E49aTsPXUUOFDv/iXednxKkK8Qt3MuQas4O4h04r2udpor3hfm84q
VUHHIBVpXCmUPHB9GfK4CxCDo/pJ6HeF28SqsUxqKVOaKsg92d3YKyNwtvhvx1ZD
avf3Ano4nGFtIWLwbpOYYD65vBaL20XhHkJTgF7VwWphiwyyQDCT30u5mVLrVLRv
beBKuoRq99+czZvP7ugKU5md5KV7KjzwV7rormmUCJBI9WWPhh0+41W4dKwf7daN
2iZBMV/cnoyTLncIOUfVseS+rm4TBtN8y2VDjsyVmibimgu0XUfusBzd97Guve88
IEfXf+Gy8OeUps6HBO9bGnxwL+pRE6fJ6mVlrXnyowsQEnuTCyPNVNhGPE6Dx5Ba
BCJq36PJyx0m8vFNQnWQ+DiJ2cvlzrhTwB1lu45c16llvFSKRnbZG8B4tQjDWWtm
BnF+anGmNRKx5pOxl+HyQSi+e2yq2qxf6IL6UwldcqyNtE8frly4fqTxvhk0QlhL
f7pmOEwnq4Zu7iWt+sJXOWSg9R0+SzkYRWMVx8jfY1RCTxqttG8UZVrLidfv/yu5
F+2WcH13CHyoCtQBC3k0jIDryPquOfnLkqVDV4PS2RXS15Qqp1sHFW5MVgkSlCz5
OoLXsO62HaiK4MtZROg2LrmXRQHdtfzsAMOOhLP47TbAsySPls+yaCsVlWrYWFVB
RaFLmnOu/GVOh954uv+DUdtMXv6HSuFevWbK+LPolsPYH8pRWTn8gFedKwR+A7Gz
frZNhig9sVonVAeqXElhZSgpEzW1Gg6oLgruCN7Ry9Ea+KDjoot+5lIzd83G+ja+
hYrWX1NSNZPgSqKzf/BfTATnxuU1DOQMUVFb3LQTHh9DVWht6e3kZJHa6CeSIwbJ
iamnNapxgekK7n3UzKeU0FgGkKgO+boDapsgR+6aHUE7o30KcmCtKm7yHC8kS4Yj
1SXD2DNMgsBvqBtt170PX3WOD8iOvAInpRjd9CkkfFMUtftRj27mhbOt7nuLM59m
nrFvi1AkfGp9BiPAnn1cFtjShhdbYZ3yO+DDWbxglz0cMVgsrGVwd73GAncC/5uZ
IgUtpku8JFew7gwctnt0zKGOkqq9bFSPLvav+2dSqSdhey0/1XVwj5Siik9DwbK9
6XtPzg/c5HXURau1sf1+9w3243QjXUU3Hot3cN4oyWs4GXhHI+IF4PXXGfCToXdE
h8x8n8Ees7iYrAftL+ffBEBheZ4vWodqSSEqzpaKq9kWLQnpc8xySQqnnjrzqz9y
H3zdPJJXRaSnkEUSoGn7eaMl4xdnhRz4TxCAHwJNYGKpXV9HqxbfQeL2DNpQhU6E
55c915LvaHTXB1Z4DWICwo6j3XUfYYoKSkBmTanZrUnVhimkMj4dosUOTAfKSNwh
2otNVNQzsh/ui6ODopNCTzojToUE+skPRdlvSQLFohST5F+MDfFc2IflunW0I6Wy
p0anE3lSMvz4Sz4Sb3AWWbByIeu+3LGBn6FSH0+SUaUDvkfphMOgzV/2JtGkmSx4
+OM0ciZeUrHzKqZX2pZRXc9InqczicIfgCCbOfi2bk4zRExGD6PncqDA3B9FoVkD
jGk2GLQycA3tjjVnqiqyuveDqUl7N3Fu8xCemqmpM7j6b9Mjf3rJ1PzQBTTuIcsN
QCAnKFAT+ZZ1KbFwlsuTPMUBLHVzMNoaJict3n0UE7sFaFX4HDvYOzJ5mv5qyOLb
iKTl5sDklW2RBiFJSp/+9kxlSSNv0IZg9or+zai50lZtLybn1SYn5CpTcNcrN2hF
oDRub+5rTgTqjlkVVMJX1yjuik4USm2NHdiQfiOav4WvLsQoXyG+iCl5PkH2PziJ
jv3F8daqMJjIQqhkU1peZemtk1vAdLs5+KUHrfIx5jgqM3mi5wqQWiWAH62A7g3f
rH70E94MvSBTPYumOtJbull/8O1//+M8FMyiibRID0DiKVpviZ2vr3I06t87CGwz
JCgkhg+rNYbdF7cVkY+S2l+9L0Ofj7+0fJ9xTC/JQmR7cOHXCuy3HrN/L1sxVcTF
oWmuIBbdElbdy4mEJ81+rw+RsgzIdH3GQjKlSozQ1+XkGO5x0XZqyxHLxeR6yP82
yIMJgSylNwQyDi2u0lvKT0F+zne1O3iwLed3gls2s8Sdr+nBg5iiuD7R+98kPgWA
pi15jXff4xi3XLM0hX29Q7z8WqMNXbGryoHwzfF8avgcK1NbT2QeU5weysBjmSm9
R86YL1NW8cM0NyN8HDwZ1XupZKuwExL5DyElqW6gR5Asdi3lDf8ZA4wh9XLlj8Q5
VR3MxAx4cb0skypO7buEboslF/qh6tsE87NiZvA8xGNPXKFJ0VAwnkFF3Uq6SUo6
Mfi72/++WMLatcYsFcwZr9wyjKpP7Q0KxBbZ2pQZN7gPUCHLOvsIF3UjEpzdIERD
cT2rFXTk8jWexTlmJsxZfKfPMqW/hwEeo7S1yFVGcAaB7U23BV4ECCzf2e3omWDT
yt9/ffXV/7SETWaVO9yefeXxyzScyLySmE25UV6OF75NjtphCYPGk2fdP+yoyJjc
ONJJK0GpKLDstgM0QNWn1uWTkL+Z8CLBK/Gld08ikAPsk16SMN/NKAQBS7AlLyK0
bERwQ5Nx5TMn25tWT/bBrZiuzbGnjCUiCXa+kfX0gLWV9mlcRWguPgCyvkaY2cI+
oyL6hy8/ZRgmgblsxQVRX3aam9A1swoULrrDiVyBBG4T2IR4t1jLMbum3rkBthvd
M3hODoVO/AYaUstGy5mSuWiUTJ6aynD3TlvZU0k5APO0HBxQUU5zoGR+tYR72zfZ
H5HgROJk3EcqXneOnrne9k2q69oGl+srI601e/pacwEKpAPk1jDWYzdzKNKU9aA8
XOgcg9SaEP7S5s8/TDpS47rQVq1N1u1GRxmHXGpbo9+fZsM3pMGEpcxZAjWormON
98nx0gnrSj5rXV1Hsy/fOU4HhdfbwHOO0oM8prnx0jxA4JYaD0D4kqw/MLwuWnAa
4op5HvcvKuqZdq3048NkIRBesPuWTCzur8jgfAcTEhH6umnI8mfhj6oV/SLrzsUe
jK4HtC/2uvPltzIw4agA1qrsfHrJdUpp3XCiK83S7CxwNwQRo2w5YUA7YX4/FEjz
S5EFTA+cJOKiTsYq024475V7HWZbRy9Loxwv3iRMOMux+fAGCu9krkXU8hbGbADW
e/DzFrJ/YPTL7im0ipXOds04M4JUyGzs0ABXKWGY8xehhoRL3x/lchR2fT9Qgw2x
MR7R5JzbLu/GAt2ZbgtQHuXPS3v83jfmACzL2KNIbw2H/3sMXMxW+sWEWoPEjJA1
H/IZEOyfKWCN3JeoBjUH/jNDvxd1Pvo3AoLpMIFvfyvRBKhL3wg8M15PgQYEslDW
IQmz8ANXazb4dmA0ozA34UG3wwr4F9BhGsyATF7r9vqL1CA5gz87iJ9BESWbJsRy
Hm5TmylLC56yXrJjhOOOJuSMwXBOsPQqRsd2Slh5iWwQ6qQllwUUFlZikhTp7byK
GxWEXdr1gF4cceLlWCgs5vmD9pX5wsAvBp4MOOQyYW3d4et3cNs7CjivQ+EKb567
HujnkJSlf4zvCn69DzBjKEqErNSIHU6F+nEhknh6jj4A1mZgJvQvtyPRAGfiyEFN
9IEc1hxHM871PEWpeCnn83BVSmmDcvAq8KnCFZVJpwzGwe4iS+IRIfzOOi0ZCCgu
/NT9WRWr/XoqmsuhgFOk8kkMk4PAdMxvFs91pjd+H5/GrPwwvhEDcj9oQRSCNV4f
pLaQlzjo7dcCUBKgUk0cneqJ16FrpdLSf2RhqncscLYbN5HahYXDRB6vGdk5m6KA
WHNm5e+x/TYWotCcKEfCejZ69Q3ugg6hjvAosDaMv9tfDLxYdhiEC3zk+Q7C0e59
8l9Toi41av3OJ2aqbcvjoCJHCHNItZ46QBiDyKzMtr015VmRsIowjfqUBIjvKKED
wL3yOqHghpYZkjB6Pd1iPvzcDqkN0rQyaVPlHrjlndED0T/C0eTC8Az6P/yVGpan
TrHfN2DfVNlY7LplOw2bq2C0GOIUSak8SY1I4IMr0EzgnuY2MxQtjbgmXasUp0td
lzE+JDLO5qRsYeY7BEokp+h0LQQeRCYPo9QBmzL+o3HqPKtY4IqTR85rk8hLmRYF
NHpKOjDRJ+u3Mt4vkTvZLmQIldEM5YKxj45g44seDaSLWriiefCVXwKAKcz4cmRy
ZaGMWN7rVAQ6UnR0Ox5T+jMdAzthpLEPbw9EH+DZ3s4LvBKZdeqh6uBwacu4g5/k
YKQckwBkTXDVrd2d8gWOPHmnUDI0YQX3BiymQVtnw7axYmPXuicR/td8t+8CC7fF
JIBuSi2HmKUFpfe3yVyRnmy0zqLNTn6kBuX0fNJRdlqoBMRC20o4fa013qU6SdJz
XmYEeyIdwS1pu5KT9N7XOdvZMIOBe+al3786Ve6jbnRAt6eoiMn0qo85ismK5ajU
TUmXNZ9RR8ZgtmoR3x0EPUf/icXy7XIRxKjWCnbm0zUODVIfzkyVGTRJVk9hbhOt
cBx30wKmfvaL5/k0i16PYqps7dY3FtKhf6XU49Px6J823P0M4BphgCPyLoI57GNX
THAmp1g8Gb2pMzd4WF20aGtfu1aLLkYLjECBxEsvQg97a/642l9Q7lmi6JAkONqf
4DsFkxG7iH5meYmvHTPKdPjDcm11qLPSzck0MVg2Exwtb6OJ36gS5nAgvg89j2hb
v815v2VinURKV6YF0pgLlm2A0webfAuXt4AimUI2wnPWJRMvg3NIxEkCr6LmLeOm
4EAaGFfe2m7iqsAtVEjjiSADlJmXVpRvMfDTXHVrYCHLRsPwtEE7igK3et9QAE7U
ey323RVV1ecUpTSHJl7tme7Bl+A6q621T9ahAanwmM24POXDAuALBY16HPQzkV1v
UAp2o4W/GCmd8AQ1kgqHJcJ7YdkW3PDJyj0qdn5Tb/r9J56XlgCwVC+C/7Uxy3Ui
Vjwa/pCGXX5i1RB90JjvYHvlN68+5SSy2TUVQUwbqvN0qA4OucZV826O71tBGvTF
3IVWyh9LiLf1NFiCvs1z8ndwSG51idV7pA5+TGDf9SFBlBKY+IPwD4F/c2rNvo09
wh5Ds/rFr0bsbpRU2Hs4obuRldgRENbcT/YfnQGAwMaYpmQ3bMEv0ooh+SbTmq3F
qYJX2c5fKCYCJU3w+QDoamDeH1utaJvqF2JCELC/ZA/8uuXhlDONjudcGBP1QFD5
qyldA2L53OCbcx2FJAMxbAtiw+Vw0CLcTK3MRgcp43kOKdGzF0RkIkBtokgl/SmV
kGMThA/8YKOcqN3SmCXKzekm65JxGBTwY09iPiRCHm60M+hkfiqdTWe2sWPgHeTw
Dzg0Cl47//8Jfc0j1JB2+434u08AgMAQBSwVu5iY+bLVRQSDp4Yn731/wLkSMuvn
FCMpQ/YyxdShekWBsi9XfmSpH4aLkHlDzgxqk0MXMCpXqsU4lKGMj5pG32ffZUNP
HP8MfgO3eJq97aGoM29DM/MZZvbG4Ec2CAp03tT9lYDOgaqGly4+bw9EJhGEB0Ch
ytIK+v6+XuZSnRRenqV6A3iJBzgQrbDB2PQ/WG3s1RMaWsF7IeEnPihvK47tE9IS
bF7C0WlcjbGaqWPTFVHOVsRifIq65iXGDXfhZKFtoNf2H3vvVwlq6iWsnIOKBT2s
sWxZA9J40xrRMIOyu2eHNy6rrfz20WCzvXreDVw6uxXEjeQGnJye6FfknNsuh4EP
Drz2NK/6Zj89KzVKRoU+j+rumLI94ruSn4fIFiubPl8+rSrMv2ZQIjmupEbKX656
5pi3YgiJ0veKH7pRp9A4skb+is+Q+pOO8nefSbddMxNm0oZw/uyJFgylQIQBUjMh
DSWg7vmSEOAzRAhrscaMlYdIrrv7W8aFxuFwAJFTBtJrl99DCWinxxwAhx5BsU9B
QYEOYv32RMTS7YmfYiQV4wB6TqB3fUEPenYyO7xv7hlGun5sr03N7T/F3wAuE5vn
9GGeUns5xzSiZ5y4r7Ly8aOocaffoF5qkg9DBdoAwpLAUmcVXgz2FGoEnuHa/IyE
BK8EBMvMiZEYKwODL+iwUDQUgvjS3UNWGJH91YvTV3Os4qccQb09tTStepAFElnd
VIUT0UZDWfx3qzMyDR3Q1yVWWRw2XVYfVYU6lNVGFrEkv5uju/pvrDCupyA6we0X
yJ7DZMpk67Q69FRANEykASDYhn6/B6bEL0K9KS+WbGPhY7Ytq15OInENnrE/7VsD
50EAa+SyYRfGC0oX5S+uy57LDext1egwRX6vN3wFqQyRmJ73keZEL6QR3s/Kc6bP
UxQ13wa8HxDWo/Z+bgVRkmvrmrZgTIy7JcwwEg8L44FNRgCm0Q0+DUWq3w+UukEp
ilNSH4Y4j0SGkrZ7qjHebP0aDiI6uSFPbKEVDrcZ5VTr9e9i297Ve12ZHLmrCiKc
ED/Ksk89dT1KkGJlfjAlgA5ua7SS3rpkLApU8UNiIOnYAqljg2SiXuGd5RUNV8gO
11TYFLtwBW7ncyzAPNzxiOYhG+1FqYkGKh9UjzpqgO0O5W5IV5HQb2Zy8Zaw8x/z
DBYqc3FrA9Wf/0gSXIGbHpbV7qNVwGNtJDy9VKWQSqDNnNJIE3QBQJCdTjlu8LmZ
P3zWHIOqSuOitQjbDTeSX2e/nJ7m1SWJHZfAfo+oTVeoNgA9seEaQCnL0DMRpJ0v
4WYI9+VupBJPlpoed3dmrRmVQYYEFZspEB3FSKjEBmQUv1Oz0ZAnVQk1m0IsZ5VW
BpcYSPgtf3xA8RisHhPRgKUxFDbg8hKomhEb7qIlbcNgeM1vuQTeR5fpk9yY+aIu
0jxhUiQVIvAsH8JGSMBwwKuvvyv+6o3eaCZwl1r2SVhXEQKYhgd3f69ZgObmKsd5
nplBNqQYcsD9BzLBNd/dpsK+pq0N/n3MnK+IaMaBeiOaFXMl1x13OEds/masSrZb
wTMfbGqJJPnzoHKfEGw5ZjtgUjOXny115LptpkSwQaYG/4sn+dYVB+2HWusSKMAx
N0YnvzxeJRrmnIIdxoc7Vn7EzAwbnGG07wWxYK5Mevu88KLzXhFQe+3Ue7Au7Jc2
OxnVTAZpVqVWO2WdSVZi/NDWH6AL+bpxIae441iZUkrJH3bdqL2ZLHf0CUnv6MQ/
qJOLn9c/ha8r+2WDkPsq17UTHzfYWtyOBJ+Ua3QOzum2BBASyl8CHLM4UIovXVsZ
h0StmEE5Kr8S6dQfZJ7yJCDqJCF2kZmgTjoAlH1/+v4dDlfzXH0Xjh80rUh/UCKa
Rm8oJ1UGdcjsqDICKp6cTW3+SNxEGj39tVlBZmMJ11IkvknpoZaXNfNuvtnG5xMZ
GaZPaYVoEwt21TlFo21UZTuFsB+KJmTLo8YzCWV4uFukzZbz0zAIm2/x3TBLBVyr
HAgFjxK2GHNqwR4PTpnYTxruu4w++V2ahf/QWsNcZMy0ueAoAGV2zxzf5ovrBJ12
/0jRKYSIXx9IzTmuMKyTJuKp4tFe9Z/K7C54lXb7EUvHznvdoNXOpVvXW4gRtxsQ
lRwk4H9iOsZBnE014hLNp/IuTCDQYyxLVbBVSD8in5uLIwl8tGuZY16LrV7rEgi7
fdnEIv2IEVljZ2zKTrb2xE6xnvabRV5jRhW2npUYpme1uKR4pnjfC8fONhjcW1gj
+Ke7YkBNlJKCLKI5w2wvpYSA985VbNt5IwBjBSbNAPWYNx+d3K3KVzZEnqnac9vm
P/8wIBFId9Gcx/BwX4AfN7g/WVsc/Jwn440NfbeyLhOVB7iCNxGbKdHTn/anI1+W
FvDxd6lo6v+8SPXhdX2DMQbxxdI3kGGzDwqcGM2zn4h+Dr3v/H5WTmUxw781CgeN
Z5cPHlg+odHMOS+nN/22aMaD75VSgffCcVulBvWA0DlXCYnldz8tN3+bLdENAWEF
R5ocBebPHDVLe6GQ/Vg8ZvT7vvS6VHBMrQzFBWJDz6nwu1HHy9kLrAbGRWD65u8d
z120i3PaGRgGsGZt5XFNvt0jBBK5lfRxyjrSUei0QbhefnXDxRGBXForzgJPs2eY
ho3KGmfDmgxlfVCZu2BOfA1v2zCxOPkpql2EnapxM2lw5M7kFO3VFSFXU7ODhPCr
qyjpa1GVdoU5h5umfRYry4PF+ekIaxAVXFz2WdeU17jZuaq40AiDRzBtWsDW4AcI
NWtEciGYmGDvwo3xzXJmVna4isbCeuJsMFvtfLtl1Cyuvx1dxALNSEAu4TPrul6R
ep4xl81oD1I6/rZDovGGYeGzFpo9hTtC+NQnpMOMSsUvYb7RMV4DFbiUO7a2riki
UvnP8rkpxeoJ1SNPfnsvNH5iZhltcg1PcKkfhJyvH/gCcVczqVP6YV4XUMIgF1Ku
GUnuEshF9hkBlZUT2NkSu3/Oy+7RybMywlowdSrgK35j5Sp5AN00HYIa4bFxqPvb
/yQU45+8RktmCIhxEsodnEhMx+aClgjc3Qc0AIt8urCMCtheKR2f+2ckVDeRzhaI
KlAs8rpDsLL7ftBLR0lLSDMSpr8S3+EnUBW02jm+ng8Z5nkGKIUJxUpnq/AF7z+S
im9YlfaX+EghIh3/yeisdkn+BRGPoE8gdf2mrrMd3Iul1r97Mv2lMUir77LNTHR9
V2VPi65UGQu5+YZKSBbZo1c924PR8Fco0ig/8gz3c2y4yi1PCGU+98023XM5szhK
VmVcoFDjZL0v2ljdwCRlwvG5iVskddrjirLclESuG83O1xDCLhITgrbV1pyTE+Ab
yHPztY6wE/wOzXl+hFAspCTjjN7GpY6/2FR4D5nvpm5UDlGIVItgPTFq5pFWCU/I
1we3B25xyFuxMXV3xTWre3x/MRAEewGc92d4OT0FiLYQvQ2SpCzRHIQmwnTk2Xl5
2Q4lVoL0eB3hWIHXV0kgFassQzmQoKPWZ5hOpQwwk6lNB5DIMtgM31ersqBAOgnZ
mIXtcrXruFlSy0miHU1iK99wwQzSIq2UeOSU/k9NVnUEnxTT/6LNns9RJfD+V99Z
WWez9yUmb/D54KhGbUDSrt8sJM+Mu8gFmPvVnBgK0FL63XIw0dcZtaF7XyYOnVm/
mhNtGhr2z0mi7zthOp85U/b0fXDl9g7H687ERkVUVcsTWE/0PGkR5HFemNlNtFH1
QU9w/S6a6fKCQrBucJm2ysK6UI1Kg81PMsFNQdH2CO2VvMrWH96Cmgz27QzDIq90
cFg7zdwGMC8dyxuW8hSC9Us8jSrhoJkE5wzMbNpJTQ+mO6s8lE3PETaAp6NR8x3B
xvUM2ephU0h9szcLoR6GVa98P0MWsaazsV5qp/S/sX/hzG7YdEgnlM1mJBfZzkqj
q4TTabKzqmv+RwOyMl0pMd88vlCzQIVcpnFt+/qgNzJYdcdbfxu3MJrGMcCFOhmG
Iz2za+yjHy6Vh/C5IMaLT2Dtua91dtHObkUmAEQQLSOkhy8vqf1rgg32TPQERGHc
DNojcYMkXSzNWCbS1P94k0Zg9hNyfagQrWdl5Vl9JM73+dDecxwFKjDCBhdZNKe6
zP4EBOdyGlzjLZCYzUvsUajv1Z6F+mOt2P3FzHUoz5qZSuC/AP/EFzrfvRXDlBAU
I+67FTg3JC+P1TrnuTtFe4ow7rwuc4bzSsC+wugWWOYvXMD67EFP2YAY1GPi4wfG
tNId536oi/G3Pap7sATl44T2dxuD98Lv7Wtm3fNiH3e4QzXqFBNk2Qy+n/7QNfSb
fgfKNQzJBsdQ2pNKLayer0mwYK9v7CTZ40Q+YwrMGCFH/M7BCyhcNzBaYEnozvJt
oRFQRGzsbVzJJviuSU4FmIaw79CXqa1hlde4tNwed5SIWfFvgM+uMu86RybfOnto
lF9Wh633Vm4QkSqNFuP+oiSobVD9dIRCKVYqxCUpdh+9mbhjGm625rXPVnp8ebMF
aKOQ/KMDSOi2a+5KtbY+jJPI+f6Lvi5yFXkrZo8I6/Dt0T0A1suODsbN/shMPoua
aVY9cF+g0pT47qyVodtjrS7oO/86JLUCFYdCgZgO5JDOsML6+faapJk8IuQUNuGj
VTu9va0RsFf3+QFC6dbiWyuyafNVFQ6H33lKJAsheG4Shx9P6mAJPf3M01Qn3g6g
ArAabntLJ2hs1nRRkVBrBV7gytVOWaOZX/kMuQLLC3/DTmKesnhWBI2jsBE2e5a+
G9g5hbjJM4NcKtzZ9zMDvwrJ3lYzMF/G6zax/iwR6De31InuGbiRoMUOfl0SAali
t2OhFKNoLHBdHl3umC2G7uPdFewHEI/t5gAjNhk/9qun+3anrQ5e8Ajmg7jGgiGQ
NI9sn8UVLitGHUlpY/0k+iCVDzuXTKzlwk/pAh/FQ+V/86wnZwqp66KG+FEIsgdJ
V9UzRk38rrd9watic28ZexDzmSjZVI+OrQoccQM9gZM7KcFBS0Cjoceng65otc+w
FzY1YpGU8/sissLqmoYYDviVP1kPzXTbPG8QrrZQrTaRDRAUR3bNth78vooL3xkq
JNZKc06/No38PL69QVc8sQ9LdBeNV+dSkrtnwfj3dUmCiOvoi6syXW4yq2L9/oKP
5wSyTzubd1+NlDwDusOSSUY5ykxVNJfn8efnR98IU97W71gdctmhmznDoaRzAqEO
Y8yZAPwdoGga/DOsnP4Ju8QvGjhB/YHzIhrENuJDt2KB/GsIzm/w42IRA3aXJBMH
bJorDaa8eLh02LbAH3EVQNWJJBy9XAhaIPNf0Mmy0U8eZJ8cye5iJyXAsjgMKjV7
LOH6crKzgV3iKnGgQq4L/IjJwbHUQqwWe8UEupIFdbyw5go+wuQEuUUk42ZrsMdE
ah7sJ1LQwhpX1cUXhEGB1540Q7Ax22/aqiU0V8xSsZdep7XxUig/92inzGOfSEEL
iollzKzEoNHGk9FmpFKLNbRy3puX2gMIQVs9vC22PrzDMDZ05+BG5tnc4RbAl24m
UvmFc0pZPcWGnqZ64Awi7pSrnxExvCTFSIZGgRzQq0ijh+U0Pu6yN9PqhpP27CQH
Svsbj/XwTUsxIL+VoV+8Kem8Jn/i24qyYK2BgrZWn2F/hPthDv1N8EB1E8b+hVDF
mflj5OP2PBxK9JdvzFjNTJyCFjwcMpeSGAvHLuGDzB4ftsZhuQICb2lNoajP/Xl3
vrp/lZjbcombNUrIql6gbuwMvU2alxFSHLQRYuqutC5G1CWg+qhbCYTZjc3srlUa
tGf8gNlL+SWhMgV0sZkk5jeh5NxNVyJ3ND5SKCTLjsdTvwZKrguTf2ngI7xuyTKQ
8SSWpN0YvGLjcqdY5UVy4JxshslzcmbR+R3zKjoe6oeA7BPoU825JBEpzgCtdu4X
b3QgwsQ3taicyZthwIM/Vl/xImdNM3GKFORsOVoRKQxAgwLzobUdJAAroD9GAHjd
AA6RXhAGsfL7HIuJF6XAWAzuM2DPch649VgFNMtP8kyfrm9fd6LAkPMrwNR6uR5c
4OcYuYIOPPC74J9yIrOjerci/ZkwHKYE1UPcANlVVWeJx2pD85XOyHKkkrVgrY4W
JYcpAzMDL7D3sY5LgmPI+q9PW+H8tkpmSKJ8/4M9j2UdVQQzOgjRv0VxMsdeLQly
WdteXvYUIs7fvRoULg0c/jmME3YU4ZJ0sgarXmABNlDoA8lZFW23zzNC5EWZcqWe
YM4oDMRdRg/D/56sN4MZSH0TiZnvBg3DIgRT2cTmee8WQ4e4JQ1TFOdvXE4EgrRC
nwgKR8G3rdRhtgqJWDVLKjYwxCdNgbnlhqrr9qqm9OiwnOR71NWFCD9YqtODZV9E
2gsuG7G5KYvtikfPnMPgzK3adSh5Bb+8IXE0uBeanuxHjvVnkAHpEOUuo3gjp65P
Epyj8NtODHeSw87zw+VEj+Ke0Ckdxm7rtUJdse2OZYAVnzxW97Q3dZek+am/Eq1S
Z4SNyF6HYTNX9v3NaQBfzweA5altRU2HC51UVc2l7RM970MVwDI03R7FID0NfjMG
Pyl70YKaZAjZg/d9SEz/zN9Hl9pBU48t2u3YpV5PeYvTXK+TNQgfd5udSkS1WWgA
NAEPDeb/r9sSEAZCqicgeU2uMTXlQ4afLZ/1CncbaBWg0ocvbP6I8SLasi+HemRs
oxsC7uixnCMGAmdr+iW/xLtJVplGtEF44pbucqD0h0mTKOS2c3/0D2Nv/7pRJeVK
8z1WGFc2s0Cyml1oDysZloJFWCoVTTr65tkVvUxnE0wd9G/qQiTY6YP9DCUJOGnG
FF3iPp12OBn1z1D5VJ9mDbD4AKJ3lH/16elCYuzxup+3TAyiRkBCyfQzJvKNBs3b
3wQhE7NaiMm44kZIoUdilmu459nc+GhhFRNg2c7nD9baBu8VePrpq7gDQLnaWEXB
sRpMBAEXoNHpYB1K7UUBvF5PhQDasYTqOgKtQZYgleL8kVkQR2tk/Hx/k+1e/xAh
J2UJuWsxAGCbe6r7fB6ZlXvxt1/0rHTn8DKSpwJIhRRaUY68GOv2afM161TLpDBK
ym0tyxIAv4g3kv7QfXE/ZLDfv5Pt0VM5/60PY91LZSwdDktZ5lH6VQeu8Dp6gjur
06EtEPkDJe0G5687C1aw5wq5l1eaH7FXuSD/qTkdcAnSFJB6/ox6g4O5KNIDYkr2
1ZuScGVo30Cvwqxv3aOkzCzOW/dzIiEV18mrCfrPabM65UUl2TExM9xkDV4xC0i2
KbiGgqb4vtg2oCIapujAV5moiwKdlhKCpV8qI+4WgJdh7Dz+KxIVZvAQxiMCsmIx
5+i3IR7GyDXqE8fsIK22WbuCbnTPqcQdCrqo8H/G2/c+1/JMa0T4dnsHO91zTfbE
xxCx0N0C4MQSE3wYhNENnAbot+rCb3BD9Cg11EdcBXaDYou1soPje5iiPIJ/xu7D
RnhICPYhbqgSeRiM4VKrYYUyEzj0s/Vt3M+JF8qAiuLo2gXAKi0fydr0IYK4LXxt
eEn5mQC54OO8NwG7s2sMbycQc/ov5F9oR85TgGaVG1Reep1GrnLSIjZIJZQTZWMj
9vWPkM29Fzp5A+hibyprAwQdWNmhNiqEzK5YPB66r8b5H/Bukl32aeguqs8haTNs
ETM173JYsj0Y2F2/PDpH6oOL1Nfsf35TbA1eWP5yNb0+5fCve5BZIomfuW5vI69f
cKxbQWtCSW+iWySCvdEtfnX39NZs/ImXvYVh2roHrR+Zz9732OsMV/Sz6tMDCXpz
Bmt+H/17M0rB1L2mDeSnhp8BW4AcRJL77Wl28CjntI1NdJQbRHcIt+EXTIIcKXCO
Wk9M7t582+IhxnEfNQEMk4dVC5k8fFvmYKTrklBD18xCk111AqLqclJ1HjLOHMmZ
fkPho2c+Nb6o2GkDTFPGRXsLKIh50vkNKhURte6O9LOtBYW4YcNffn5SFKvY/CDh
nvxOfobIbl31T8HrkGUHp5LG3MnRPfWhzv+x62DptM4Y5Vjmt/I6J4baUjtzoPZE
DULSkxTWoH1EMyuxdQmCQc7H6hZs14h5OJOZJ/EGlv3av3FiSnObNhALjI2ruj8X
O2qW7Pv4BwDXPgKBmuiSpHxwl65R05gFUE4SWia5k1NsW14+LjeOpFvYNGbrTzDv
QJ8TuJ0c0OUf47MiEDVW2tf6hguIk9cbLTaJk1hVW8cHf5wKkeoOSVbSI4FAW4BA
JBr/4Ou1+AMGOxdRA+sA9LIH6LOiyWKG3AoHug29W5o7YxzZ514dNOKr0epmfmm1
zhX+BUvS4oOVJfnZzgfJAfSK9KrMhc5X9UELJZ67x+rASoY7v3vRe5CYd37w3caK
7XItB/VYsKpwccneWl1bcDvO9uiePV8jVwFnk2FyCe8aX90MrndB78gqE839aPJV
FZZ+a1fP5mRv71K7xVpzwgPf9QVstk7lGloJ52+rHopqfMRIWBG28gNTy+QJ6Ma1
nURO1TiVVtIit4HGO8JBRqLbPCHrz6ALKQwnqgq2YQUoU0UpTtXpz1PkJQyP8grK
K09399lGmoTtBxsEUR5hEK8mbcouWqFUVfJHQnFIOeTWaT0u0OPXWIxsQuWwlArv
sNdqUuJ7V8sHs1MgOLqnxt7tuMPN7pr6hoU57Oa2Pa7bPi7To3ZjeO608uh8cgM2
Mm2MnGe5DEijRAfcWm7IRFnvdclBucVYigX2CUs7/a++L1+SfeXf3MTKPf8SOgqA
KKO0w7qAXpdng/IgT7hGK2nUjoThVKesj6LTDc97yecEVOXFledapVOIVUyKn1ms
bTRp+v5eA6bAtfgE+urmvm1VHne9fDX9qKAOKKiFadueBeHFUFITYoXgHvKmmdMR
5VK3CZTqJU/zaO+fpThh7QGYJAS8eYQadxtHnwnnmmJ4zgspf3eAyPR8K65PPDLY
Iz/KJPd4VYPKxCIlCp5weamdBsRXyNq8vvZOXg9kqIgQaK2Zab3GUcaZORyPIETJ
YcN/ydRz074bSZ3UUhN+8ssVIaYCIl94haCY0GdquhwHAYHPuklAULG5E6xFOCzn
JxB2hw1iBU9At/hGeTa3O9Nqa/VfraZYe7Zw2iZo6xDdStdlIBhy9f0NgsYM4tIv
Vhb9XmHHlUbnegtnPJFVqrrZncUhvspFsp3HCqU3icaO3xecr0vBnJg2r1ED7Tum
zM8J33J37uAORWhDVmCoYveiW3iVqCxkbtXcMTrBfcIGSt1B3rWkSZelBRlRHreD
HqckkxkHLIvL1DAJO4hDAimojukNJfQFVDiR9rXdznBAZ1YJuXjJW3UT3OdVXjnB
gKY5sHc6QB5RV6jkAfQY+3/4uLMp6ep9SklQqw0yILqxQvKfqE4hUSB0hS6TsZSi
3JONGCEx/L5OELWrGLlqo+M3RO//1LRbAKhabDbIT91L+1nySwYv5E68RLzpyzjP
9vIKcu3+ToTedSa+vDa3MXNZfOEOXK2jMu9ZwK5OKuC6pgaVrgA44TclBh97HwBp
gDY2uCzBohecZ1jdl0aB2dBqHwT/Ij8kMftoc0ELKhloSG+EQ2Y56TC+uvSZjqXO
KK61mVGUw6nKxyB7jxQejf5hWAPpz1Gi2aZmlpeDyfa9M08h8WfjTOB31WrDB8KX
4GjarO5b9aXiPumCvF8EZn5XBeOKB+rp7qQUS1YvJrFGUIoUBjxUsp+Jdv1Ty/5Y
5rxIXcVLKBtdA9O5X9bA/JT446JIIAp7EXvM957L6k4X9nGZOXJBQtoDYHAsE8Vi
PAVRUVCGeC2Z6lZoKVrUmaNIB4WZCvhKJ3zLg+Ro1D6/n3QgFbrNp46s2YAYF1cR
AcHKdgyYOO4hJZwKMMuGT0p675Gm2xDdmJTXqM6nDqi1KKY2A84BAAkw57mNzyxj
ZhePLML8VAy1New7zXHxTI1OxR5rvyebEX0tfKLB3J2hxyVUrwCmE7GtF1kqEiFo
HJc7NCtiE6lk8E0v8z+dm01SOgcQ/+mKP4rnD8DiEVLkSU58EZZSsa3sPKsr2YV9
c404GDrsutuR7OW76vjEDqUrLyCCv0Nv6UCDjTHzw7eOYsZ9tpRrlk0A3Zmn+DZT
g7O45HLKuI95HKfj5jJJINv5lAYrdtXME7ZpspmgBd7c5aUE/nyA/y7blSubz8FD
asq1oG2C0osAFpp1SzPe0APs5jvwvGj2H3c6aVp9n/iZ+RT0/gttE/H9GtD76BeM
rECXwwWTag4OEgaL57eWrzPkmuwg8aJ3Ni/ooYKZ0OYD5+sy6t8/zXOKPqlxXy0F
zl4AlaLbnUDSJ+Ff1PYQv/i/6c8QKiSLyeXVJPZuSKvHVsrWa/cGtBpvY5ykgaXj
isghbH54wlzRr7Pf6tLb0nEmrbSsVngLeyUCUcr8cS43KNcehKGQ+zbHRhUFf/GX
u+gr3LQhig/XkH/CSJvqGcbVOjzEe90zObiytANixizJ7uFRDuKcW8aCa0kfe4Nk
d0KyfAVLRSpVNzvtR0/QMXA5hvo/RWzMKdckSCV+ZwGA6oWPPSB5/04zq6mASwOy
L1xvbIOs9Il4fBuXaOtvd8Qidn1Ffd0PAYDxZ3aKnGFCk6sRH69htc3QCSS99lEw
rDFp6oJeFwkwxCG7vZxNRgOUsTUusua/su3dJUkvtIjbjq1RW8h9qqKl/vV+yNGR
2bgreI7ykF4apx8m+4/1jmdmfFhqMx5DgZbkj0+N5J4xVgtAY6tzr3C7TgwdJv8a
CPZ3L6HlhF0JMwSsXi7yH7xr5AUaM61pdoN5jkQyQMkCsGUUP/qwAzWKNnlRBjFg
FLz1DmQkvngF6IxOnBt+2RgrUYSL7U4whG2nKOTyhxzOq6p8Te92rsiYPV2Ief/H
AsRVa5KXCOgR+IpGK7T6HLVL/nmOFWDo4HITOWS+iFzJiDvlyYBWIos3H0RgU+P6
yyKUjNlVeB3miNLnFf7WTwyHvkErqiZbPDw6vf52B035FggEVjdkTdxNg62nICAc
dsSinH1mciBE3vaiy/nEsEW8aJA7bLTbexzx7lH58AzoIMQrBklUoWucdxUfye53
n4+G3LjDMmkmZOGTPMCNjGW6CCFYuCfqdBiUJxhTz/DcTAWDFRNWuXXaaSEA8r0S
ehhP8FEfJ/CzWVRu4vg3OV4g7javHkebR+Qa3YPDpYnmYy5p9ckm30+UgHIZmQH7
+SdHk9//jI/Dwg7ipcp71gP4AmsoYraxusC+DUjbmc0o9qhMcx7cD2m2As6u6t6F
wm58TCwg1ZHhCXM6WAxATzvzktIYda7eEUCUWQ+NDHyJUx4L0teoL73ntnn3ARGr
VcYXCzfhrwE2334neuZrwLc0Y9jo0Gh3SqkxV28pDQ+J1cKYN4yQMFbB5AYfEhK7
S0UcATHOxTUJUZqAEb2ROhjALSr51GUU3lZmi9F0JV5KQoTqJce+Jn3sfc+OP+xD
8A2uHrRcxyfyIH84eo3uFpGJhEXe2O/RZz3qG7hPRnpRdrCJDQqzKBPKBMhqBtJV
P8KKZ1xq1l8FfvJoVy1G4ImW8QvXWEdfwaRUh6jikZ0Dl8BXZX05G89OAAEcAdW7
ALnniap/8/vu5usbTxJOM6NenIzjXMuHks+MKvvPoa6UIdw8lq7J3pKxstRAz5aL
oXLN8Ax+I8NrT1SZokzTxkYIByKr2WAQUtSpb2khvTQavu8A64l+5OF0Fh5svbLq
+Zlx2mw7TUSj3jMRDSoJ3LqTjqrDnppPiSk4h02alG3HXyumK91xVIn8okYa79t0
8VW4OK3AO6ey3HQqyiTnQE8a+Bf1JoIp5rhlTq0VCRxxX60ZUkg/UpDWJOdu1Bs4
DH4PMQlyQiYN1ixKC1jUAF28rSOrneVf2M2BU9vTSJxr89YbW0doOFWUx0cVNhsD
PRjAPK8MBJNy975iMALj2+IE+ShREVh+2HCr4dddBhLIigEpp9BpBU2Wi27qaafQ
807lD+fRCJ/H1vdQ/sPDYtxly0GZjTpnv2vJcofqNyh2YhdH2PaJv4rOhvnf10Lt
YACt9VLyy7qF2HlgQGOL/hV/LyHia98fZhNeEOro+9ItjkLV/9W+qdCySYY3Ph0h
d6ReXU0iRflusx80caIDOT6m+bh8H+jMlde3wS0FTza4j1cOU5JyEH97F1O3AP+q
RiA3IGCIQgR84x8LmTZgJ+j0+oPYuXE8oytCtaZcRy8+XRE3aEMjU2EhD7vBaxn5
h7k6a1XnEFIu1YKIk+m5iEkPOvw45yTcVx2IgyjzXH02ZhXOlmimTCAQkb3ccafB
dhoXafMAVNQAzUpLbKJHtW3LFRlUBHGMKrQqCVO1zavOnGdapgGdEk/gehj/XZiI
ZnMJrXMUaFke741pkV7x9bYstd0iqB/TGHu+SZhF3Q/RnZvdjcd6cknJ+VOeBbAV
b9LN3J8kVWjh0diJhx0oNTOYFahaDYgyNVj+6kcL3NWlwfyCLFOlOgzM6fRZZNSy
dAcuRv+U5cJxc/xmkiMomaNWPtKuU6Wj+NsV+19PdUAyv7ELtTecjCHlm0yB1cgf
QAn5JAxjz1YdNyB6Es5WObdEKiLDJILocGRnQwiLZ9bmsiVMEMcAL7Yw5nqNn1F5
QsRH8bBiVVcGUvWKInGurXQ9JakW8HEwK91tBTUXpdSFzVXVbaXYER3roW0kIuyt
ARid9xql6kAGwp8dpRy98SpCAIKrZKnr20qV5fRqoC7mohD+CFCmOAJtnxunkOOh
YZ8kiFzrKQmV2kDm0uDlcatgWWSdoohV5N2Rx7LvcceA4cvr1pRR2C0b8izelsPJ
v3TWW0mrNym7Xug3F8T3EpdpVuxFeC/x2pMa8HupYnvQx9U8jERlVlZDoNUMNuak
8uNNH7YK5ZGVzwk0pfc3bZx6nKjxLTNPT49sXgdUsNXiPjhv5X3zEUdIWgVkcfr+
iqwFGxnWtifUHHi9iq/edypCBvy2S7fowpJLHpmr3OgvEHFYRfEDqL3EJJbsdP7o
aRtU6PLkuJGN1Z7v5Lo7vvXrN1wqjCT7VKLgaIqN7eD9FCRbjevQ4ryS3ysUeUvt
2cC/FteiKIJbGeA0XjF8LOp46HEt55NpEhmKNU+nnE7WqxF48+q0m3hwLdniiYTM
Lcw3GOaIYl6YDwY6/Xbbg9w1BWyDdjS0oh+TyhZt/qRY051duWQ0mwUc4ldATU5C
rseLlLRZFKSK4Jsb8mj/a1O5qvsZIQuMTAHrybVXQQqYS2TBgNwWWYsA2HBB1cqz
3yegfzkY+lC92zEdZawNFCc7nPxS3wySpRmwko6goW1oHXQqAD5eAbJS/lXRYloX
EO5MdTtwlbYeww20VpMxRvS7BJubQwLUy2iMr+yx4HKFoY9Yu0Xa/4E72Pg2XzpI
zdZDr6VwncMSN5/x+Kq4DRpacpHr+5I6sBsufM3f+5zWabjKl+Ul9X1yl2qjtHNA
HiJn6z6ndwKa7eOzEsvy1/5FoclWFqlLAdwLUNVi4f5DdFPHWSXyseYVgoVAi0l9
CVqqcyR6tWSxMSOHc5s3TYiDnwaWYKqjDpp1gFl17InUe4kmiyuTkflArSiP+S/1
l/+Y0z9KMhoim+sNiupFcoqAmwu684mYnbNQpf95JzXo3b+jY9HMn6i3MstIA7vx
r4p44Fz58C2WXrXRZa4Giq4Cw0Wv9MANxj22ByT6S/NTwJUcisP2xCznYsdyLWIS
sslp8HhQm+0CxSVgzTV2YrX/I23IpjZdDCtfN8pCwUwFrzxWJ5atmbjSAgqRdbAW
S/u390F9WHPGVAXM6dNlP8rvv8p2/gDAf8Y5BIEwem41NjmaF9MW+NOiBXpsTFC7
6pHX+TbmK7S+wX9Xmrn4P6Z9dto+R0Kz7clXiCppu0YsG+x0thtud0SJsV+hjzvs
WSxsYZV2Q6ZdFdHtrusKg7wIFR2cZki3UTBJRGBm464V7chiW+B5mkPEfCf8AYnb
0eplrWM2+rnGs6iYv98hooFI/4iFuFkU/0LTPc778rJCevN3rHT2LTtoZqxd5xe/
aCY8BrWO+FJgUvWL3PlnKb3gfAA7HHnJ3vKlPdgMLxqK+q5/7/PxRKDUgtXR4UBh
9un8+O9evRYtPME+S54jGAfmcUEzAQ5HLtdRYWDVx9FBQITR7z//q+ejJ+CsjGtt
y7tE6yD2Za8Du5eh6Ohg4sm4rnIfGz/gGHMsb+v9KjodBk9sipncYSEPD54mwF4q
+cNbGR8jAjZpIBrfuFOXSJYGTG7vIDZ+e1uWQd+o0CttdF8hFuZgjdXiGBxAQthz
/6vf237zPRQFBP8SfiLKzChD3oxJgxIGZJGRNOepG7n8q8GH8XJzYoaMhLvtIo/u
cNMpiOLyQbCP5sYcAzCfHmALdczwF5EAQs1lCrsIq2Y6bW+68CAxnUqEFJgJQY3l
86VSKSdfsTn3IZXNeJ+C3qkq2H8DgTdXRrqQoMqZCdY78ob1cFw0lXaFcy2se7I0
GYTWAZQry4S1hs8zdNODTCjWLh0sk33OqSA33wdpRl5wCHSYEoJZlNADfwO4AQtp
2HKGRwqUGO9InITs5Aa/JDLjrDeeCAA6XU9EqUgx5KILLAo9m5iyrzIWfJE6AgSp
jzSD1yDbSMLMAYLKhYq5O21B5pFCRpUaoFe1ojKi3wPbQjbaTBof2iGW/SmpU0NJ
M9bzlhkDVKR3w1sYXrlMUKJiL02xCveVM8szbOrTTH+UOSn/i7o62QjxPRwwz7rv
OFsDn5uswMQ4t2MVzcdzYLtqZ39cNG6q3WbyEUmOZQGAE5jukce4M7ntXe52MlgZ
S3/hOvSo0IwzeEqxvl/zs+e8B4ZJ7EH7fkilBjYzGexEP5gSOL9WIXCxcFoqgGjz
6xjd62PwuicdAd7WjwyQX9T37E4InHzQVco4bK7Y2J2bnGjHKmxD/HLPQBGL1yOV
mlTA5wFsO1cWjmKRrA9VIvQ8unQE9yACPl0OOXqDycInb4U06itC3utQd67gpN5x
ZhUtnGfZf3vz8eUuaGTobH35BFmPV2SMUjRcwKFJ/5VXdahHPTDQPcjN6O/arCEl
LGkOvH+HA0m6vxuAbwHJ/DOx308LEg0+gTpl3vixxhi2+JD9bxCTSb6n4dBx/jjG
LjUTP/T2+QiVE/bz2vRwYiPioh7QZN0EsauLRnZyElrdua8aWGUQVgACCL3BY/+f
O6IBdb/dSxSPmU8SPmkfvdo5A8s+785hEqm/X3sNJ2lAINKLma14pJecRgM8+AY6
zNbONH9W9CBjuEMBwQbuZ7jPB14fWGyNRIeiPwEauGZOSNSXWVb2FChe50sH3haq
aIBEA1HbWevN+0cUzmle9g3z7B01NV7XVg6CT1A0XspNDm6cXDMnbw5kUBJDYqxO
ZjmqXYisNDldPWr8Npk0zO62Inr1eXm8AU4Bt/eoOUwzaLCHeSuPj6klCZZ3yb83
LLuNZPbxwXnmHmz1ZNxiUPdHbffRSYuxgf/mcEKH1zUCkGWz3skV+R5+9DT/DyOQ
7fB2pQAYWzYRkrm/CTPQkOAeyiL+2OfBXtq05wCkNYxUKsaTb7Vp8hJwWfzZBipN
tqTt2RD6zrEU8Y3M/7Jm2oRjMJBp354QdNX5YebtaYTbki0YVGI26zXUPi7f2XcD
JBYn5mPM0k5Y5yOUuHWpwuqCnK6c8Zkljv8YYUghna+rQP6bwWc4UE/JF6oFcRD0
L2wfKxNghtC4hmqhwdIvGOjK68rZjTUmyhFebYdEZnrCt8+QvQ4p+1iUGCDjK2sj
H0hj6FAOj7dDdVJyUW4Ru+VUzupgErioSMw3iPRxyYZsd7vG/vB4NEE21RGmTdPs
hLbaTpECmOaGVPAVJ9Hhk7TqpluIF2nY8OFBenQSe3/aWawogcFElit9XZaUGzzy
roFjrYLW6YlqTXV1l/DyRBmsdLrXYjjYXeqvVauQT95P8d0LbCIZgxXJ2BofogCo
GJCqKFtS4YywlaRrVQba9OrOsDOjQBWtcGwBUSXHmvvH6zF2yetzprdwsWzhfgl9
GFz8204PoplffaiMtFZQsNqqnnlatRU4IJ+zPFL7pSNAk19RNNJUPIt7XdE8wVyb
giageGYd8pnKy3r3rvoUqxWDEn9G38AmTrfszNN8Q3JFt2Z58NOmeVrEYthnSY/L
QTGGe4XFgeZ3qOO/i4ntasG3S0xNiZ4JaCbXJXL0w5BJfTV7wd7EaUFYSTXAUf5D
e06J3TJIrEOjULHPTCZYCsgenlkPBFt9sKvrP0hshWFMpllPsazg529i3AkIyyzj
3gBtCmgZ1XtmH/pBPguKCih3Rk3UsHy4wdU19Yk3vpWFbiBJXTM3pT9xdMxUSA9L
e0Qs6BqjMUvDnhoCAb0ocfgQXYfUPvvgzoGSXZTYKatgcxPWzsm3tim1AND0OLam
2fIizr4OSue1kB0VN/7JWxn7sFsVu8BHthXuGWreaElCEqtntHV9BRVw+FRxDc4D
KUz7/cDCK9uIWzfn8zvgV04GRRYonRPAAbFX0+tT40CdeZBT3sEGdBuYPZrUEsnl
+a4STPotyIU3X6DEXjGgL9CjuaitEdoXYzzQiA2frQMN4M0V4yBkA508pr0AKgbA
ozSEIygo2HN2h0X3u6ssFqACJ3rmyIjPmUPAttJppSMYEodyL/lgJs09hx9gaxd+
EE3NdilYR/tvGqKJFLNCBDcvmKoPxahTQymaWy4/K55HF4G+0yN+ks3hXckJR5Lu
LqXdjp76y3NQrJTDtXwpSrc0OXWy+LtGroBoufrPl6GyojouBK9yrn0HVCIwJsnv
BaALuoFG6ZjYYWYD3m9e1Ugw/cyUvBImNoLpZxee0PRIoHwbs9s1giYyAMHGWMaT
EUpzCOGWsKqea0qhOq2ZBRDdQl6VGnB5/5JmAVRYaAefngKRq6iMgVwntneTCXBx
6dUox9uP0azkbC2JEjTf8kE2ryCuhhdELRjuxDmN9JWO1TP5H3Fa2Cx5bsTu3h/W
hGxgLRoqm0JxbbMqBABMAiYbsxSB2Ck1/wnIm9agML3lcuXzOBIq9HCv8j3Hqf9N
vxHm0rUUMwrRpbkGsWw+z2UqwB28dx2BXs7g7BANrHRIEw+7yLtP9617xGSdsrg8
FUYBxkyceCSRf+ppAVc70Kv+OJnJxlmotJl4g6OLesOYslQP9dNy+hV+ji1Rt6FX
DGFZR90HV+YiRipICBtVpii6UObHNbRroyMDkHBq+/lgfXcuR1gOgz4Sch/6aZPk
J+em1bCJiyJ4mcw8r4k7FiyDdsFktB/9ezA/ORIa5BnEeRS6OZNtITF37C8hJjGL
wmRgnqP/ygsFo3R20mNb/vuUpjb+VAsABHZ5c0EngctGctfbyzeXFEPb6xFPvcII
2KiTZs1cUo9Rq5dl3pOZ9xKKqQK5IsL+yRKIIw9GhGk+k8yr7vPN8IKk4Yyi72z/
oHoI8puaMoAVFRdwQEVGHfv1Suk+cRZpe9AqWgR/7s/hHp4RwE+qbdxm9lXS52gH
qjgYcXrBLXAvfNMk1AZNNbbRXcqKfX/E7iXUS2tbaolZba0ToJpluIjzPEc0tof0
PpwQKStyrOKlPxDrqBhphBHT/Y12srWbajdVmrnz/EwD7hvHNZ2OJIopp+hUG+Uc
bvOysL5vHcLPsvaU0SOqejOSR85wm4EfyqroVn+EamBwZPy8eAxJpjTJRol2r9Zb
TGaOE3YCWuIgi/uBzSTKAkOFpTwRY4Xk6aNplWXMxftTpbFYKBslKfoi0GgbA2Nn
V02yBhQZ9gy8MpePKx1rlvstgM3PpzNCXdGKnCPoW1anhBwFJ9B47cUsEcnuTTMk
x6W8uMn3PG/frOc934WoASolCZYFjo7ULAAQGrQ+SXGjAKu/t7UybK/pMASx7IzM
6JfuqF5bhjKnAh9QrNBPOOgS/TbqoDcNOy+DXLkxqEpDSuOHXlwstP7hv/NkwMB6
YgqoEsSobLPOI/QbnIgXgfOoiQAQ1KKjJXz+9ZiFyNz5eij3gX5oZSAoJ9zK8MR6
JLFrmgqr477wT7Py3qLcUJJC3DzGEwmph6/bW0r4BAvSyd94vzfNQm6CzVdjqT3Q
uwK0VAo+v7M9lrICTCZo5QHraG88kVEDtcBO0nXl99Sp0dnUVcoaiaqW1E5O6J76
KrU7lhdtYSMf7fYFdTyevs7y9p6lSFT8wChdGArsuzLX0JdcwKONSAXL2qHgeA1u
2sKklCvp/FCuRyo3oGHvwPMQuRXkGsDfmhn26lQca13N2yIz9UU1ZsUGGXcOES6r
94D9MXzNihEC4YXUk0nhYi89EF9jCK6VAvl9HNWWPdzxgVGmgDGgEb5JNY04dzmV
piHpTO7wue89zyoMO0nLmPg4BsLkmBH666UdHIlajPkvwUS9RJ/WD07dF3s3MtbB
ru8Hh0OqzTgmCP8WrtsikqlgT6r2OrtZoEihvhSsfV9e+xDtqVZUzdnngmUdp+hi
PTqRtaN4mBl8+1cuYLwn+kY0An8r2NS3XrwpC9ouNvEsmjTbqBrAu8dL+d+PgqiS
AkRh0o4/UZr6dgptubkkSSxAMO75lzW3Ve1dpDcE08N57N2VQ2Qd8r+2fkv++E79
AonDIzW9hhf7RnevJOu1a6p0qXBhOR3HmHtJ/MtVPSoosoW/iU0Orl2bJNK4+Yyq
dzY5PInS1ZGjn1R5zZZZZMP9a5CF+2Obo6posfAoDj7xukbe5+vPu0e3C/7LrtsE
IvteDh7irbgsX3aWlMJhkceaD0KHiNLzPiOeuIFycgCFS82nVndr/r/WyB9IVhkc
A9ryi6zbkIQs5Dz5+C22lDYwqgDZ96TA0BhY5848MDqp5Q2DnrCRx8wWWgfLoLpn
i4JfA+KgzEvbUdmMR+b8nh3xYMeKg3R9qi1T8S3cV8I5Xpza/TM5ZhhfTUDdy46c
M8kQ2z7PZ3CVRcLttnAMaKk3+t8B5+0xEZ9C/FVcRqa1AsZ+7LQapWptxdASr7h+
zb1jyU6uTD9b7suLTWMxdPiWrAUyyI6+FBx8UelP6Bc2LiAZWgQFPVdHrrw3B4qZ
JO6Hm+hYvbwAbIVYso3iN39VAVYzb6D0dqpNb6BIQ2z73glrDynzcsM6pUnOgV0r
TQwGcTh5B1FIuZBMqfihlYWgabSYku/H1aGCDG9yu+PmXm/pmx1imns1irBkOni7
ag6S9yNrc2nkiKT88GeKygm3ShhuFWcwM42rGbJ/pqjRVAwVmNCSng/Og92c6ZAd
BqbnGOl7+8eiuVo8bjl4cvQC8ACnhliv5UqDLlMZLjmhbfqCKFAJJ2Pmv8hkiihV
cvTWfteIlLKYCybTNquM4eTUudoqHKueN3yJZWJdj+cbL+ModsPx7DMAUn1caekM
B3PqRqhRZ6f9D4JzWvjZFk9Hlz9ItQq9vzWHQEUGmS9eVMnfPByFWIs1v4rON6iT
VbYcB4wv2lszNkVUCvlKZ/Xw4A3mdijfis2OSiyDG0Rr5gtv35Qtf5+VSND9Y+yY
UYyORpLnE1e7r/wkCa3ZAchHKDNxQLfg38wqEudUecGAYLyHCe62oRD0p+A3ksHH
gWMDulnHU4RU6d/AQettw+9JN2L3Ajrrvm9Kfdemp419K2O1yniw2LIx2sjvtf7O
OGR6F5zSlrLGMreyMnevTESmXwqPMtUrlzZ8thUCJxrGgXPbkCWeo5l13ZVYe+VN
9aDo9DZsHiMJrls+GP38rJPHgBtTKotWmbqqlhqV3hlWPQWMAeBDCyJif0YBcNqf
kINFPVVPYe0RQ5JIqK3IlavJIiydinP4P9sLFfslPV/Buq160NYncHFQjU/AdiJ0
c0ZCZPKZrnUPrsBZEDyU44QV6R6MgC4Sz0znrAyZkL+kQV2FH4Ii3pPHwUU1o+Yg
RvZEuDizJTQVeFQvy11uOUk7+jwrXrNAIuJH3kN66m4n5X5nmYiPGIXN/gf6XyfT
iIDz+bV5Qbz3rpE3Q1+rc2YqngrxciTJIne30ekcz17Lsf98qR5vLn3tZgsrL24r
r2BHdggYdWkubUApDOgRwmGJ6UE1ZCbmQNuuMV2cy207zXE1r3hQn3d/rW1UgeCC
651pr76TjsNY6Mc70ianbVR5paiMTyncND2/eER6j30TcS7MFP97Fn6QMEYaZFgf
lBv5Q3kKT9OI15hWJTVWjEFPDEhLYlNhAYvDKh4IXGR8KJw/yyHnScZuKwkWIwXV
sO6Be1GBXArGiLLiXl8qpEpZti5ol61nnBe+WUEbuIZJVEpvbRyCK4QummVjUWV1
cp6NjrdE5vXxuESgIP3x2UppfOqedRACDqqBAHustiqLX/HMPeocXql5oiQwU0Zp
Sxr/42D40QVqcPGMTHOVl1IpURggVUXBg4m53BmnfjYmB0qHoMwzB7f3AgjRUx3k
T4ms7uc4jsWNMmk4dP823AfQC7/6OS86kTtLpvtT4ZRSmgM9ua5O/pQhuBb3witl
KzIZ0ebWsRVArAKnU+9Z70vBBiKYqk8mGGt6VhLFAzI8OkoMfHdV2Gtd/VAxxblx
rdBvwzOsfPzXh+V5KJOh+60lxTAB28KhDoeTM90YAHFEhkondtWYGQmsezvy4Msa
JsbB+FAiLoEJoREX8lOvrLXt2hczMAjCAthc8Th/IeE5wOoeg5VdjHwd6vnOtXlJ
ajxn+LVHm5mwfsN+jKmiA9piFCbHChUMoJNP+fG48D17Q/0PLlr5p/jryswnws3e
asf9e+YGBj7uWqLgZpxDjwYcFB/WFZ0i6Kz+HqSJneh070OOdtFuyXehw0Ingt1j
UAwevHTTkxkSRmICz0Gj3FKx/Xlp5mgTmNSfgLeq7sFSUTMmFuAC2aaeq79voPRY
dNLfM1qUCuDIjn8AIFx428GCGL2b7u4NCFpWgK28ktIPs5esVMko1UnsuzuUuJof
wE/qFb3fna48ceCVfCNoieXlkftn1/dsvzFjiO0xIK5vGzcWLGEjRw/CCIEiN/HI
82IELKTt1HggmVXBfE5p3EWl9o0II2AA2vBa6NiW3ipubkQ+PS+x9/C2w6eCxTwz
5ItCvM3r/2BIHOrekqjtywfCw+NoUuridedI9nGNszDtZO3yCaQ6hL5wuMxZxc33
aKfdPGWE9u+9kHPveIewyDybPDMe35+N67zKfia4VLiQ/WOGt+V+n3yb4u3v2lGE
45LwX4cSHejdUu4nxw52UyAWtCQOR4AUx7YISJy3uHUsUY6UcYJAZpoFWvKNZGu0
FYz9fDTTOfH3/6kt5MFv8zl9W8eVXcYQXo8IsXQDa4exUX2Cjm5LwLTri1kwK6eI
6sTm5sF9tbo8aaN3J0AH4l3lFdFzZefKpK3IEj7gMgvgDufsoz7MX5qKbgHiyO1s
zX8DxwAkdInoIZ4V2bpTurclQucdncZMUoLq55AvqfHfvx2BnA20cPU4GowHUXZn
ri/n0GnIOFkRISyGoP19yok5lu8v1KOsoNKrZARQAIQFXZbo+lSF7Eepr/6ftnBa
9IN+/yw0jf34c4tWXMJHdhTA/sgr5SFec3QifysUggx98Ti7MDwS5JxKyWcXJHUo
fHrASX8dPIFv8b/b+Mxq6rOWux3bcsZklFlQ7V8mvJ+gzp0k5GkZ3ILo2+DlbkP7
fJH0hSBkFNTw2BAlXhBAJdBzs+gRd+nax7JT1KnjsnhNb0PELRlshBe9kQEQNYi0
j2+rGuUdi9kF5CsrWEIPx877XL1W34Bd6ssLHEQXAloL5IwSNuybV5k18tT4A+mu
mNgltKAnPTLRMHwzvYNcKBOgSyq+WY5eNwqtPJZfeDc+7eT5QpknpPwYK2Plqin1
cyVHyzL8HguNEb+8LRRG5FxnoM4mZN//ixHI0s2lomdb8WSR5yGleJb2f7mC8Sjd
nTAyZynzDZEaV8iGq2cLYlQ9b+IFQgJBt0+XwOs2cckBluBR2LcqL6I/l1CF8tPH
1znXZvleQB2NZ8pNXbRQB1nvqkXXEkgIYd6B1bUva3ZjIWb1BnP6fMnih4E04AeF
hOZnR6wXvYXFoiFUPJOCi+pd2li1lNffGOu5oPgLbordzei/Z4EVAIftz71qhPNk
uArJ+jo7L3r2el4M7hxwUkvqngnJbG3DhlrWmehXPEq97WQKNlQ4vuFGpyjvVsJz
hJPXowu02foBKk/2DNS+67TUENTeOo7+PAACOKD0SwTi4IAGhFaxYZ+HIJsw40UQ
uPaOl/T27ArJ18uYUv2RF2hZOXVpnbThChz9UMcfyu3BwLR8Z3DhUZcs3A82MWH6
HJKvwBYcdKDNC/hCslOv9Tpg5RKFE9+q5bZAFVbfsVeM5/a1cwydRTdkfVDZvjTG
m2jOaLstpFr0yHQH9uCL4HA27mTf4KFqc6zJ5uudqz1TtVZ2X27+z7YTtGAnO7kV
7s8LcqGJwF3PYJE7hcLr18ixBz0Oma+7w4N2+VMmXiIJ04O8dnxJrW9QeoLokTfL
ap5nCISiKsaqylKimIzA75kYjDWmPWQLgx9YrHeY6a786oc9ghyylaEQ3OY57u9G
aNSFjCmBS3H43TuZEukjDfJHY5HR/gzKRiGSudkAmZDnS705/BjrnZfo5T22KANA
oHmxDO4czAMt24lgQYXh86uPLjo1pKhhi4S2SItM1KVEEnssFNMhOdnkpd/MmPzB
qpPMUM7Ow7cgLgy1uitGpVbbxQv+Po2qeZmNvsLIT23o7s3qVZ1ZiHNuFJfsdvkE
/LW8uQ+FCg2NCOM/cRduvoLM/+S2JT6aj6r0BJ/rOXUhm0pahIoIjcoqTOX/8955
6dtxKKgWzLQZ7wul2TzaRXCziftINFzsuBjH6GArbhR8rgFWI2BRSQKxMdnifYCf
92jec5Pe4Z+HdE/iMSbnmtZvxZx44O6Al0x41wkCfW3E0vRE7PxNlWhyxpOOyF3a
BOTbp9VCXVFQA4mFAYnnmDLbA28adohUsGTshoVaIeDFa02ketOwDRlXA7IqcpLC
ZwbTsKKSBxqEgb8CgqmZ9SjQKDhgKBq2wkEB/1nUg1eVJgdrt6kNiErMwB5PANAi
T38L/D8D9krIQJVERekPT/Z8INxLc8hQxTpPf2cWDbuWzYk5Te2G3Gfo5gb5xypR
gnlOs00p6p55NJtStmQI10XC5JUzm4jmRhwiDRgr1BEJlUsc8IKRe08sSpbuUxhB
seoSsA3YZ1MPWFXWME42/913z36Tv8iKO9YIurSk1v3fap6b4xBqS1E4ryjWbvOT
C6rrYGPhq6qBIDunSC7Nt0hpFYCqbnqGKBHjn9IVQXL7Ywmb/TB9qQG4U4M56sQt
E3L7tFofjPUlaRxd8YPUQF3D6n0jnFHn/wIJ5/G4lylvX8BpAL984i8VGLR3bB/T
aoRwsxsP4XSzIMQBTzNo7GN+CkQ6pMiAaY0CfsoXXpMuXuvdjz3RDHi9VRxgzj+P
Jedqj8v/TYKCNgbg+YCY7xvHKc5w8bClziglwiZM8eWj+bFECztGXoIIzOqw0Dte
leF7vQCAz8RcGTuazdzQdbMnKgLFM4MlFvZEZVizf1Tgqo5CNuIEYiRxOnK07gBA
aIMHL/CKC7KOlkCPZX+zC31ptiQwnTMCceaHWMy1pWQa/pR2FBA2aQukLVL5mt9s
56GDKwuIGVEOJgb+fMEKRgCuVuDLE193T+4L7aAbS0G9CpyEL7lXy5eep6yQHP17
/4n3B+w9rRQKsWRHHH+/RmqTLVr/W50pgwau/Y0fZY2TTBUA8c8auKhYzOXcaXkz
MYUKubqk9EaBHH5JEItgHibjvglFKWwzjrZNajgtEc0LSWq2taUshZuMPc+eQ0bt
J13TTXHcALC4EyanU6KQ4bd3EqxaAuduZLUlnQ7OnPMazyrAmq4JdudbkCmiskW0
wEco7T8LXMnIeTCFhEJ0MTDVogrDH9ubNUkeaZtHdWBElR9vel5ypWJ+11bUg3d3
HwwF6nNKwRPQzK8YKxvU32TAJrVnZNsgPwLFl6bh+loi5Lx6OjpEOh27Rur/CJa5
83PwzevD1DhAyKIdt2ggf6YCo79xmeAjVPfaQlygIsmqSaKr23AUuSw16e2Rrj46
anop4uVkXD/vgQcP6NaL5hD0Gm5gPCrhP6DiTfDgOFH2Ep+0YtXe32B6e3+zRbQi
v8bf9mL7bxlmQk5TeV7HbTsDBd2uJ3d9PNXYvDlciNtu0+4jQl8NmiQx04soN4S3
/cPpu0WLFxd5OtpJIaU+sFWO4qK0mQNxVe+6XgzJyA+TK9Dp+i/ajmGPUUHMKDIs
EKhBmhxCRTqLYLtkSUgeta36wiUgXzcP4z4thrvOiiLZt/PPGq1wLVdb2QaAE5NG
PkSoCJFR6Ll+U/adwDxzzaCdax7Y8ny/ez+Jvq1cqHW151USvqM0Zlasd8YIodZ6
C1wwrn30tYYo9KgdbL/2seQTQiof/eg8NS1G4Ln7E8Q6K/CozqIblnBR9cOa+GQQ
15Fv1YPug/QTDSKrR+1EqFgfgMDNQ0i60U15GzVJT14ADN6rRYLtVNzBGDLH3aP+
BETUTvHXXkMqozRqYTq0ScxJG4WMTpJ8gU8r3GPghLe3LI9yXzEEQ9i6zGGravMm
PcMNx97h2hRLNaj8DZujm2rHNXs2WDrZo4AljVeBtR0M5dUplfRiYZwV0vUM0zD9
vGGcW3n6TMrrQEtkX+tL9dyMbv7KJ6qSMMk7z08+q54KsvXTsC9PyeQMQTEBQ1X5
kjttApJIdDjGMIv7KZYCXDytwsg9OeRRHWhfM5k0IMQRp/y2/51vEy+9At2X+ZLp
BcK4TCm/f0JmSyZGTlAWex3WM/HsiL/Qgv/iDctyjOREFMRry9g6H8Iiq90MPPl9
bfZmU7IV+At2uX9a/CcqZ6ClACG6WZvo7VTCEbozKWKaSq+kfvKNScoIbP0auYpy
F3p+LNzQ1Jr3XorUbunJB/ybKa4KwZ5cvf1TTtakimsuaWnlth1NQiP8D/+o6TYi
YL3Jhr+ekUbYk+HW9H0TpsKb6FKH12t5Y1wJiNUUfA38buNk8yr2fMLJQQ0epOKn
H8OAHJdkJtUydinXZWp/i466Qz/B6yHRJs3ezr7u098p5HgC+5tEjkmO2VixKZhh
nCHleZ+1EZsu1SiyF/FddQOIuW15820Eq/tE0rjW9Y88aXumjQSxGek70s3MDtY8
iZfwg4rEN0R4Wm+7y9ta5XLv8xv9mvr0nGUZFcP0WGWepZjSP3Yyvj3xg+djVYIv
tQeLtXx3tAE+BMw7cy+OWuCjoD2esy6y1RU++3wltxbFcqNbBZ0+LjS2jGdTmFw6
+p1HSBf/AkYOQDGEuahLHKkZksjWVph9fgTKTpGlXqpHqi9TIPTSjW3818lUyr+2
Gxf4QfjSwaa8tlWUiLhnf37yo8q9a7OhuePD8LsExWJ7J+Ul9BXy9qorYbI05kbU
yU8IfPSP1XDsZwe7pzQg0uXVDkz5x0sxbd6MREfe5hFJGaqvPdQ8jWfhBwwrqJnK
diorp+ZSIXU2DkDksgwSiiqXHs3ENnGFdLYzTNAhyYuVrw4aPZYMAfaA6ieYtywa
vXYwNz2ChR2nkbjCTZAPsr6MOs5zw9R5q/9Pjcy/Bnb2lZKpooxzV0iqU3ylNEbo
XvALLZ4GWxJfEqq3iyiWwyVIHGvknNjZhl5Zwno7zUheqYbLKcA55SEmOwNTFujV
tZ9MdkBk0hBrmI15LCCSCRjIijxQIytdxGD+LIzFStm0nTIEjrasz/IuX9IQZhBj
yviPoU/nDE521SMpR6vLq/JSi5TxyPSsCZ5USzHa53Vh/asYYjNz8BoVhg2jJH5V
xw5nT9NXNUZnfnjFbkWTtsrda38OBvg7O9GBVnCiSP+zI2B5OBBHcAjX7CrbpbyN
pml9mey/IHPtk4RmAhCpFZQTnttEwSBI4Jjknpu4kAWw4WX0rGJponfMYT9uSv08
53eXAH8P+OMgGZr1G3s6c5ExRTtjmWeXuQbKGEvms+vZ1snsJW1gy/J9MlOAs6k+
ye2saBjuugcfsG16HSry9MlQFIu+9udRnqpPApqVLB2K2W+o2QSretoNBQp2vBSJ
ySUbLM0DJTyQjFkAz98xTM7+RCZsTsJ/wTUwroQqXGGUZu359BMe+dONjoDRDjff
KkB497C3HrRgr2DNLu9/++T4di/cXkLVTKgu6ejl3jkGxmB68izelyi+JmUdI4in
gOmp1FBKS8CtbsFKoEUtXt7/5m8CLOjS0iduqlHbE/d5JDEbIuwrb10qankOnqLl
7yAYTfuiznTL9Z1BoUhwdM5JcWLcyU+qK2xBclEqL1BkBb+SzGggLmQiQ2bw0Cn3
ofgWdi8G2eoH6T2+iiTnYijFwkolVEjs+xJRy8978PzZ+asXlTfMqlafFhLYZwHx
6K6siHEQvgei4oBTpOXutrXhiTtiYPzNeWXKyyZFbZN3cb46FAje9JeFi2YCklwd
pFZBeH0solC9PAYbpb1r0Jsz2N+HDjL2ByP21zJDforJdMsclD9QsXiQ5QSn+LvQ
JAb9q3jrr25tFx6Ojmt4a2ushO26AS4qdMLFSoIrTUs90dvBEJKM50XeJkWYsj9v
wcuNVO1j1ma2D3XxUFSBC6Ce+ZhZZBvAM4Uh0RbhOdUqhIcRX8CnSXe0n6FqyhVY
cY7LoUCk4WxB8+8vtWOap53fyGMxvhDlmOX/12hD6RQFkgPcPet6iEDamy+HjHIT
Ak2e1XXeJHsidmd3BxpLgccr9GC9j/UbdojCCUbTzW8QGVwx97xvLVYOM2p4bSXt
JwCu/9+HkgesUt1TlTgvIZI3b5mEKJK66Vvfd9wHXmtNyTLiIBFL2XUGKTMaxMus
Mq0LZz0sGu/bsCw0AJd9fDHDR7G6WVNuinziFha6u+jrby+Ucxeilju67qGLQCzX
3BJLEyEuqY6RYIaOo1Tj18YNwA/QOW86u4HBZT+XGodYaTLxHTQbP9ONsC3ECvu/
KWeOkWsCUSUcOG3sd/2ETOGS3m8K2ejUo7SECcP2Dj5uBm1aBwHD+0/zIjkatIZE
D8UUK3J53H7UaLN4r3uaJfUwUjmdd2IApE+miFZraCD2q8Nm3MCIilLFFOKNCmdr
mbj7OlbvdEMspBlH6PEqkjFAhDrqV+qN+9C3vuOzrqqn1wvmcgANq74WDjCs80Gf
nnQD07fbjuxhWzbMseXtk6hbeoIFR33hCNTrEMu7s79eGUQJStWHjBxCgZS6pPty
1PAUaWIkTmi0OmyUknSzVNQqQbsmzW19TUgk8BCKDRw6gO4pfN7kUfuc3Pn6Ubzk
kRnJBkbXyirIT8aBr7oIkA+5z8rjWk6lHXbd5Y/sWwszQYT+7IW1PRGgwqjvh1Zs
sNvGJhcxjO1zekMLBfCs12nAIKRXnaqq/f3XXFBcM18dXKQquddjInw/WZkNuQE2
P/KYjOersjAp2aDiDl51h/6mXvId+PvGXZH9ylPXzl2b5Iv06hwsRuGH/dh+ojW1
+ahHxR/KuDd8ROfeSF3uGpCVd5HrvIOykjpaD2FlNRFjzKZiEO60L692+Jkwm/vn
rGesD5VzfXOY3Mom0RiYtVYcl64JxUH8ktIDVUk7zEH2G29p6SenGc1T2idY3WTY
6x5ZWDku1KWg/2c75CzKx/OPBi7hKgzQ+UbYapc5+iRPpZB5WTkK7WC7g/GxH5xi
phTW+7NJEGEsPekp+m+aPXwCBZ9Hl3dGou0aQtUzTxtrfNPgbyAdUNTFCJBdUONi
nkF/NfHXDS0YlI1gwk8vergp+JVYACj+tmJlI7DvQnhZEttkygWvf46Yzd9Q80lb
u25Kw+MVRuJoQs4CV7aXiOx5mC65NtiIXY/8fIMGwos3XksePre/9YuqNXOwFz+Z
oYmrfIlyRbXOxyEcxpmZZEpE+nuW5VdWXNp+jTyXf/1I0XW0QvPQDdZzI9jdI8+S
lUI9hmjlETJRGhduNOuhSINUUdUE9BSpxGrFhCfa29cC5+1r/Vom3D454+dpkcdu
WBrWGp7jPjn07lSvfySRYcPHK7D8kJaHqlRRUCOK3u3lBPt7XHrXn2EG6rDzYhR+
jCzCfHPGCk8jeWQ7FdF13M1D8dTtRyHwTyecf2G90QB08bCBzirHyZQoFovfTQ1k
Wa96L03G265Yye322xxzjwRLsAaWz0OcV92k18QXiijpQ7WShysp8cfY4gkLZur7
D0dNNR1cC/Q1DPDF04Nrr3xly27SUmIICJxHTk1r7pYFuv3eiebUodaHT9p/9PFG
JCSf2bYndP+y7Sv+GkC9csK8GIqNjzsmsj4Ytah1huKOwzEhbyNCZLwI/JT9vif1
ao0hZr9+WstONcTUwuPVyxOVqaxho98NSo8t4nrv1xuD18FXETanNZ9+R+hyY5tO
bX5x9hg5g2tEu5tInA5sTRqiWXVfx7jpC8viSWOzVzawV7yzALQGOXiJfLBJBJEt
5vtaA7ctpSB2uzw11nsFqJqXddptoVJTAg7CQkTsTqvLLSX33Eeouh/PKZVmLWj8
1gmk5FZXGNSvizHMbqusLckpjBAnWBKrgpkRGurp20p2VFK2tpGRd8LEApR3T/Nu
ymq0BtNkwBWDNxLUF0van4k7+vkSZICJaCgKLb7y/F7uQxTR8eOZLuOQL9CmFyIu
lPS/nCu9hAvR3CWQgrK9Lsv6EuKPYPPtkBx6aiZdvo55euDNvtwZEs0vO8886vG1
BxwAcZgmz7X4tvdpxjJ1Vbshqll9xY68k6ExhUZoldXWctVEwT3JXtQhK2h/E97d
o0rVYPkdsFUitcrEuH2yew9E2AzdUeCnKtTgwt9RJXR4ugEK1lX1CctfGCWGWMHD
SVYVEtDQoYZP+b+sz9EazH6eiIDkn1X10XWFC4abKOjOfU0k8QpeMQqg43nJAEiL
7hJgAou22B+3vmWT92JZJpniYf4kW0DRFFfm2aqy2030V0m6dI+OJcenmpVvw2Ry
7zKKKm1GKa3LCYOAcEm490Z3ApFrDNipRGikINio+0EtA5qeMQyXr4f9KjmBueBV
yhr/PdtUVJSel2+LbV36ojkT0Wuo6vt+8X/vvXoy3Bj6KKd5ClJvICyeS5t1qzHG
Hd/tNcZyzZoo2bQ5oh1S0OBg2d7zRKuQh8J/fvPWGYueA8QKr7B2Z9dsHk5sBm1g
0oWbIr7eWIeYux8PwgSqCVHm8rLkqsTQ42hkGmSFD+YptC+3uMh24u9MoDxrx8+v
m31e31ELxIGLSnhb8hw1UL/mtBy/XnZ7CCiy8iBvXpgHHGIGWNK/ViXt0OgJrUrS
GrRGdX2fo4l0X7esBS0d8ZDoglKLXdZbASpNPnzRdArUgOVJ6XYiqMDRexivohon
OC8NNohMJ9p1cEjoDNFmS+pNWle+eq4rvpZFpwredu9+c9KFZ/MzVksti9UN2Vqt
DvVbdKUguURW6RA/OoRURNh4YkxMx0kpfuRsX6xKcb9Ontb/ILn1AMxymGCQu8WS
PWeGCuvGtjbssVRrcgmfu+pwNX9TLKSX6ob1+j0hmx2nhfRBNjb4uyxYzWkn1ETz
T+S+ZU/mTrXyS3XsWMK+1+Ex0L3pG3BvWtr7gAyTrVCucTCzT32Xn3jLjFZaaiMB
nMz4jLj06Jpz50pIUUIOx3Ux8/qRAYLegIxaQGjWGRe3dYKNkqYSTqkgpJr1CfzD
bc8dKjy4oxlPXt/9ndvx+EafE7fBnf5flX4VZm9YJuqNGvm4MT9g1r25VbWbfxKr
1dasGJPJWHgdXD5L7D1mLkkaA2Et7vwzv5uPvAf6fapstaV0tUMHCNtiErJ/hQ3f
G2QuhHFrXzNLL0yyKtquARu6EbFQwWmQ8M/UO5ZBK3jHe07VbEAe4S0r6x7C7AbS
Mcn99qI6936zowVEKXmmaWURvR9s1nf/2h79b2LrSODHDT7No4SxMEohVgUCs2dt
duQtTzWmhr40n6RuhYdDmB+famU4lcdgIo8btuaKmLwlr3AK167/gEF6grqujCeZ
RfMzMoMhpiVY6EBzY+XNTJi1oMHseuvlr6UG2Ud/AZrZg7i8z3Saho5ZtBV4+5oY
/UXACk/YWQ/oQgN0axsT6P1Iktbqo5TA0RymnVlLhpDOOF1s/T5Y5wSYcg0vIj/r
3z63W743GO3izlS/LM0XEYK3eKQgJp+LNPqNR9a/yjVXFKWcOk/YnTCA33hgn+wQ
6kVVcKkH5iEUCzRqWIo7GB8LiWofNYNwguMDVwVUTfidhPvB4LbiVx6PDOPmFh6Q
MHpOks878tq3kKD2/Poqy03OWbPu8aT8b//iviTKxYrXXKhZ50DvLpzgB9PT8bkd
PfBhRwjEB8sOpAUW9lFcyIzm7HbUFpnCi8uDHPD3je+jpPaZnHR40ImomuMt4Bgy
JyhfTJ9oxNqE0Z5/EgAjQKiXbRYGqRsUpvRPbww9ORqNT4LIFehIc6SWolSBZxWw
ZCmJdfLfxD+fqX3c4IJ++GKjiG0gLUFLeGoPgFnr8VeY61hE3vwu9WuYZP6wOsSN
hiTbkzlqFt2bThG5Ian29u0XFG3E3TR13vWDEi6ur6ZAZwQhI9qtf/p60ZUQTi8r
zseSJQ7CN8X+J18DnG2YRdxsPB1sdALE7HOxFtTjk5UJt/8dQ5gQqL21KEzH7p3R
XR42JkR4+00uFSwfJtQgkPPp0TSQwcPwpPTtEUN4EfWnNZUeI895yHJBwx58U4+b
xMuyXV+sELYnV8thV9GcETa2uONcTT51rql76kDttrqhdCeFzteimFzYdil/rSGe
9M2OCp9kNOxNjaIbjxlpC/J4BpfTNXusShDsD9rPGZP96rlFXuuTizpJc5MO20nT
VYBwoJPx6eKaGByzTiCrXjuUOe3p63sG1cO6uMhSbE1N4fsUoYRQmt+tXLCh7af3
Ms+o7hZElKV/mSazsxCaDwipq0aCTkSiuL7IjSL21bn/YGXCk7jldbWv+F0vyTlq
zip6jTKyYd/eVkJRBOe/vtihbuAVVBFM5FV6mi51ZGZTfpTNz6ZkejLIaIckccBd
Y6NudhyNM2zb0Ze0o3aYlLXh9dFKSC3XdqL8CQIRNLiJmiR7hc/de8wqKvHsGs2l
pQgCLywWrPIKq8Me03ck3d75dbKyCksAOwkz2O2irKa8HuzkRqfMkwyTzUSttRRJ
gHTdtXPCXrHgEjpdzlYVuieleGWEZ5RjSUYikhU6FvAv1mZq8kJPahOrnvTm08xu
74Cw5V0SU+tASYXpF4iDjCvDpCDYGcvZHRWlXCqQE+AkllrldlPd51qTEbQ6TG0K
q2xxvAh8Tyy/WTGxcfG7WVjpBakKlZ+RpZ6ucR1DVtWJUp458c1450g5XN1DWGQJ
h33yZfOsjmKORDL4SGQCNgUp7EuKjzVF3I9cDg+Jt9C0x4uK1StK4qgDYgaSxsiF
Y6V/aatLSf8tDcgumQQZ0IE04JCqxGddo41KimfQN2Yo8lAg6IYkqlOSXmDLRJKp
D2eMCncMq3/jA3EFUfpXq+CKl503PgoP3UvQ4oMiTJbWiDz3PzBq5UIHs8dK40Ru
hz96iAOqNp92M8eKIFaWSjaS5iYQtP/qzA6rnR5vyS1FeHndVMGFq+HHng9plu2+
TbwNBzOxjhQRQvDMoAY5WZXOWBFUgAuKrSXFRXyfEK2HVEyqoRfyYShnnTsTFERL
7WHr6BNmk3E3yrbN07Wt9iJRtV/I35GyEPLiOfzZqdC1+kdamCuDLpSjDO99+3CR
snvyAzWe1x9qEqMqdJ7OYX+x+XN9LE5oayjBu1ZvdbiS04BG8R75rU8MNmn7Nmks
a7P+CVTy/ftuDm2MySgorcNZrkg+MD9tdQ0XZJ7lITxmhFMPRJVz4O8OlWQ+m7n0
hHZKnomTc+fHPvK9M6NVVoxpuMx6vWHlI9Q8c7O/6WE1pkmENUEv9/c+eE+BxXCN
FMnXtnn9GXty/vsi+uS2rzq85fYklqrVMQBMM9pNr9HTr4bUNp2BszTXXHMCCt2F
6Fxt+nuyUHc+baXM1jPKWBNk2oWE+f+jMrllRo91OAD/6amQMOL2XXYp5Xow3OEi
UCaKYLaB+BPM4AsKtpyG8wPrGBSiecT2niP+IRjWyEI4V39y4T31JA5LnBb4LOVo
5UIyUES7jDbHMZAnYD+LBNqr/LWcIL+1ebNay3l96dM94NA8mC9DsAqKSrcn0rQi
wHKYY654fgZMDwXvt/+Ixr4AwoGKcoJb65xDBXf86wvqHjLC8aV8mdFrdPVKDGMU
AFT0KWD0uvX/xHnhe3uXDiIIedYBpajobJyFU742M2xI9W+SgtOsqSO5DCTfOwve
zrRQrZvPO3vR+YmhwbSzC9tsvBdzb/2QVp4WDVisYSxAh192c20LlslyS0htS3YB
n9n+ULGalN/20E9B+ZW+fzpfRjraPOBCC/aWg/1qf/be+QUtpayc/BxQCoh7exiM
b4XR9aLtwspNsNovz1nlcim0Ay0eTCmjzQxodhGw3VlWJX39sKuBZy/BWYXI5sm4
b355Axc2xVVM/FrrN/BBsoUeOlmNZSvyEs1Xt8QPb11X/nSwSE80ShKd63GHK9wg
/0Z6ajNG7Vz1RR0LvOwSHJLgAJXmOHm6jd2UHdRqVLN41bliPE1msVYDb4RwWXzk
GUGv4poJK3LsDiN4XX8LlXELGkCjQWpyMOjzF9ogPB5enesSDtex+0E/SF33NA5W
kGJ+3FV8tB7vS6KDGWEI0ukD7pXpqxczuq47rKwDZRbinvadEKW5Ddkzgk58WSgt
k27Pi3CRqcW4dQXOuHplfzzSHeOk+MATjNMJeq0bfV1zvI7yDyBmG/nCakf1xk4q
G5af4YpCWILtJFQ7r1n/nEI746AmdTnDvxYgni6GX0QFzr2TEWI38D5FHp9R4G7n
WYIhTAQdqvtR/tamG8Pw8JbFcGEyPEJZztpDzNWk3OVboStuFdsI5u9q3npiLUoW
BynG0yEe35Opl7H9v96daPe9GiFT2e3RoOYUdVd+8utubrXBgHFNbXR7DTCeNE+/
G2UL0ZzyrvinMjfYn5k4fbqMH576A5XtF3DK7uwYzaO1YNe5ojEUhB7KaijflvfQ
ze93SDGlcavYTy7Jvt+MjB7HsBJEhL7NXF6BBk2ASiDmh8loOdmGBBv6XocFvJLG
f63kjxh53JVTg045gjU38mAsBSFaJvUHpkrv1gs0EHDfYdY9jhzlqDbgwvg901mw
YhpV/ddolH7jWfWEiQxoHLFYm+XotxiFODvh3Kv2eHYg3KIx/gj7oXYQQ1WVBO54
Rzx578wIcC/Yy+vaTgJTYh3IdHPWPg6JB6vhMZoJW2U/40/FVVacQTowREnnE0ra
EbEnK8ggE+1XK7rZ09XLnsgCExcepsiaPFwuOTpjN9nhCYIDNn8EatKunoA1aJVT
KcVvap+KJiuIvnI6hf9jW+WXaP51wS6N06Ep9EPTeYUvwprhWXEBOH6UQV8dhSlQ
yeOay+R+mlvDTrO++zb5NbppS1fBsGskQrKlekRHncO39zrM9Sm+HPmiy7+uStur
LEp14ei4OZQK/Q7uxSGLcQLgDlG/vLdp4NVVLxNOnY3FryyKkgUd6rO4cAkamOy1
7U/9k7jSUeaQKmut97jUutmja5n55ljld5Dw6taC5D5Vj5oY8ZcUX5YLGe8ZJwQh
oIYx9X+m5YQnx6WhKkIdyJFAcKRVCdUeqLI1CtqUeVey7otYn2CTeCW15hrNzKpV
UWi+HyUSBKQ/sp82wWJv2ZEpTwChTA7vtYOffkyoEKohnfbrS7RAe9BLwm4Xt9x4
lD4+qY4couska77KyPjvOqCn+S7mdHKl2+VjnhdRhxa4EBMS7XLopMOQqGqBgtGN
6HGsVc82+dEG5Vd3peQc2lch6Lv3HqamYZ5GZVOiC1uo6+OqYn2EeVIgQmRai1zz
MCDdXXR724w0dTNC98n7aqCxxF03hC0HQLNWETGsJYlaoE7cldFe4gd3633wMC9b
Ns3GFsSVbiTX3NhdRaOVnnd5JlE9Y5hk9G2fD0I0Xo1R7jHME2wnFCAEFkiJhJ+f
H+/2DGyL2x0Y7Oz24rYMDwtPUk9ZkNBaD6GkghZldpmeq1ks4RioEDqunSiywAmI
+W1ALqKE8mjG5pM5QqUe8YAbCdiXuvuIBaMMvUnQxyud+KYzt4WK97o/X4ji0xsw
S5aLe8IJcSkV3Q6ac1Z+5uxeRe0QXUkpwt0UeDSJApsPsGuE/yTRKyJ5v9HMcX4L
eJFzw+95cDkRE8DQxcIMjm+0Ok3rM3pbq5ATnw0sMN0+we+fqT2tfsv/sOR2Kuxw
g/PgIfkJCo3sIBUF92Qz3MtqpNXyK3/UvQJOSxoIgf2+XuA0XpHF9kWnPtE+t2Xt
TkzpnWudiEEfQs9fBJl7rDc1v1OWhbNd7mtdO7CeUdpIIn6zdu9AlWRcYxuxIcLU
oxLWDBoxY7b8q9S5AGe1MDbTgw1hmQtUxMKwqA1OqrXZqnkqSpPxBE0eX/PzIrhd
ESJ1sKQOBswl2MVG9+AoyZqISwHixg5cL+xVPd9fe+AHRAXJjhbauZ+pEC68aJBB
eN4nDgnNQ3WUE1eBHuxiRM+7pic1PmPEZJpbh9hxwO10WxdASPrSzvjj577Po8+b
MwQRfFRSvvaboe89hpGtjcwNNxCURicG5gO9y8CvEVnF7fOfWLviASaZaZa7IU7w
YhPdpf3V8DnLAVFktKc7kh6ti7Xf0ddcecnTMV0qrN6TtQogqMETj3hpjCCcgd2W
82T8fFJgVxAIMWl/vupzzGKhfG5w4/RHmrRNv/GmVxEjByjQVC37rKosh4OtXXkK
4Q4c3UUW5bgUVjhijDisLx6cXQOM7mZPBQ4yJE61gkYhkGb+Pp9pQRW2VPfFR37X
E+WFTdrIuYuEZ8BhuoPw6hc83sa6G5pv84Zt0e67u/gkLHDBJDdRzj7VsBpuQKwX
L0ciCBMyEy99opmgrMArYmu/gTDOhsdjqeD5oOkC/ulCyzlC+c1HJRWfosax5upD
uE3LmAT4bBzHsRGhmUGzDCj2eVxbhQ/sL+ZDw45mK32+cIvo0KIp+gvZYL8udsHz
T3lgDXqTG0hCF3OqCfFN4hVPis7tCS+3hLFWgK+6d7iNhMw1GEPQViqqnQn4AQx1
C7du1uHx5CjqU/0QEXW+VDiIphHFwJsuLIov0e0UvFNugsP2q4IsEHDCRj0NaK6A
dWyFxn85gfIVeR5n7/zxVo2zuZSSjexEH0PRlJOpvCXpke7yt58hJORFBSdNSqiw
pLHK8+53PzOHxtGfdKdCA+bgkGG2jIe/aiVh/BDmipC8CLgTT+pUGsgeE9t/efz5
Jo0J2ySsJBd0opf1gHF/XtmDKY5zo0gM0WIjv+4MMu5U7zPTh4jWRs8WM5UG/JVS
4UXspVlyM1JgY5QIJJQggHKxAAS9IVC3ALHNQ5aLbtcpmiHiao87oh4Qo+5t0KLL
mvyAMXKiKrD8NpMomCrcshSGi4xjQLEszEHxzOyjWJFpKOeNl/HSXmw+hdDMKFxQ
Vf1XSl5ueyXsXT/BSMK9/Ho714ECm5qaEUXQZkaRhNXvRsFfBWvf7hh6HYeCqFyC
Qr7NPfGQba3yOUHpAFhyFQ98RDjTCG9d8gUyfeot3tJA00WRQAovi3wD2u0Qk33t
zjFyCUNaWi6hIGcyyBYtpiNx00tOvAE/jXwaC21BaJMP24bssx6rdWvFxrOvlOwU
+Ttgf5ElNduPbvGGldZPnSFEIPP6ZyjHwPIin8O4GmaPvJjSuiVR/jqT6En3gKB5
lXNqir9neHVlCUfFUXtHUcD21LiRlkUb1oXG8k8/xz5KGjkDtjZmaow2LTQWLbrF
gW680Tg4SDLETAVFx7yRk7RCT+p5Az5OqNP0b/wrFzPkmTfdV7Jwqygs8UPrvonH
9YHTXmc0CFR+K/0LqD1z/zmDjekSiJyZY+cb+JomlnyJ83eCYGjIAKOJGbq4/PBI
0HPZ1m22snkumJTQUDYwrSARbR+hV/CoR2MZfaJGmTaJWYrAC2tNSY+Swlw3Targ
/2d15l3ffzpvcKWBfy28HD6OyhgLLQtn5nd/14I/VBY26pTMrCOoWD0mreXvnA1m
wxRCksvZo3so9rHNCSMAxnVuE9JyzIdfvQdvwIq7OlYnmY6ZgYy9iSElBF8tKtG8
zWpb0WhomljZtAz/eU/Es7c4PP2e6u+XiL+7fAIGu1lsHTMjx3gwNMadZE9OyXNp
D2W2/z7fcGzr3DCr56R+AKeWs900cNsqb7E4qqDl0+OQWW5IZ61umdK7KiQqeSYi
teKS3NV39fTntihHg6tk2rvkp/5ZPwhosVMJSpSoZVQ66c3ncrcUvSzCK1vl1NOc
NflJ7yiic7xHqGxY1rzmyJJ8ovQXmyNReDkMD44cpT24R/Y05Fz9/wHcSZYON5zs
Tk7S1mDAAlOCThgYBUWUYnQyt77QuvGkxxbvTmripiMx1Nly6MUnBikAORP5BrUJ
I2a2jYUckYKfwAJxenqIbRFyqonF/OxPiMJCIDxEL3Hg6Ghg/45X53AHMAMYdsmY
QFOrQgMD3XM3lh7n0NaBwlPmETcaWkq80uTx5T19QnAL/8bZMsCwWN5R6ouNAhsh
SPDDhyBUPhQZ3zuGS3qpIYg3yu768OouzL8kpuk+V8TlZJFdFB+GGEF292TY3xC3
S9qy116wwAwth/zAkp7Mkvm5JmX136cMm94ZqnWMODoBdDPdfB7PCugq2Pdzk/bl
loGo6Yvs9/ri7iqr7PbrGygNnXWdDWTYfZxkc9DXDe9LeX7oTs3w86R6zqgweEjv
p/bLO+v1DY0UFuxB/msGwsoTnBlL0nWExHBa/Jnd+oKKAXUOk48JO81DUvKdQTYA
3xaeJPAaa8Dwt7dPiJvEw8emN8sCPqMsHQZjmRgIcbx6jvDAVG0hXfCNTkDH3hBa
IkxN+ljVCfgejObldHa0kBM6JU2paz9IizRSheixqzlji1zGZSUUSC9VQIOuKicp
ezHIDs0uJVtD0O7V+K5hJtNiNhKbDxff6HdyYNDYflPSTknkzKluIsnLfO1ffSKT
yMmf/kjuu8kFHhjemJWJDXhyK0fS55ttEi7Ue1zPSdd4f1Dpq4ev7Ab3356/EyPH
tFF/vXuSvv7LFqOIXB8YHzpLp0udp7l2gUbaCQ3AZQw1udO2YKPPfGnBV+R7fO9Q
Uui1bTLEE1WzTzjeeaGLEhx9sgaDsq4JrH5xmDjYhUC7ZHTz8dsb7IupC9ynyS6z
1cFAaKNmNoUHCENmvBb530QCZ+sLmJI27B6Xm+aCfUHqON+2zXfTFZIwR+JQFLjg
5o/O22c4H3t1fzqNlsxw8lDd+KzyHgmUJ099fola2zzaIOGuqiFI57cx61w0/g2h
w2r75+Xh6GbukYsIj7bepQsXV4IxlFqPTbOs9SzwaE9Ox90VJ2ZfseG/zM6WLkYD
5Whlgj3pi3HfFPy0+ArsFfC0NRAqX9ku+NIYA3hR9KNvaCx58DsXD+aHyjjhgYEJ
kCPxCErzE8X7i4PWvG6Q+NSGHfmIAX5D4m4y+vdmbb4YVwTcoLIzBwtZBqUeH6fR
ETQ68DhoDw2/IJ59o2kn0VGgT7+QDRxY49vOjcvt0/1OAIJkdzXYC4x8yDBuvx6W
XpW5hbOOGGgOIbF5ZXVTHbv82VD0FSrYWjtoNAjLXy5AQy1YeSlqL+JlsWCbi8Lw
izVV3aN5iYte/ZjDaEPFpz5qoknbQOgdPJmFPhem+ywNOhb67uf6Ae3gi3qKSzuH
T40fwPq2/ZJsDD2pGPJEcKKVmRn9mfwPCiDfejSxQQpwdA1owqOf/6/+TBQrBIAe
h0NMDtTcVcjpnL0kTczEJ0P0OGVfmehTQs2+0pWD8W+WJM2TmPQL3RM+npeWszz+
snLUYXNNPUv6J2yFnDOLm+bqqW9rEHdHGdkaGP0BON8V1H9XbBl5VPUWXE6dQnog
M7PTnTgSWNE2KmIX1qsMhlzALWfJ0vUtX3XbBX1CIcA43/9wQkCTrr4xbbowHoyl
y3GbbMAQhOQrW5JVEBr63G8JaFwte4ylW0uvA3Hc6DTWxUsLFFVORJassXYsyaKI
z8h79tr+PIozckracBRKnMu383PktnPu1wr/HKvOyUBUOfSzgfJ4pE7YKvZo0HJ+
m864ynjp2yTat5IOI/Yo/adlEnW/qQMBhzfSxdpb4kxmSCl4U83sprE5vYBU8jz4
vKb6Nz41Xjo+uteWQpQaHo+Zxo+ELMC4qyaDe0kcTEXLSYRE6LmRuT0pAqmsVEL7
r6d5SaVJILt5O5rqp4ePT3V8S1i8V7g9u8uH6nbvQF7Gc0N+5c/sPCULLKBO4KJi
Muz7JBsfMfMD8lK5FBv1b541/3MGbqiUDTOwF7ryVc9O3gmnFX6/LxW60o2tXtiq
oUnKu2SOZQ9YQbdV1qiSwFfhqOXUqG7IdOPQbpwFK1TVdvkyuTfeJJpdWIfKVenn
qgfxX+xEcI/0QbyFQxorFBatqvfRVxWXHeFcTypC33y3w2f8+fJ6FVEUPM+FBotW
VVr6jp10OD03xwgav1cOALzyrlEE7K3RRcZ7R0n/raWS1ZS/G7L63eYH5LOBl+UV
tUNWNevBRzALUfBoeSjCcDILRfn4Uyf10hhcDFNFQ9M7UstBQe71POxFjuDjW1ZH
2Uc7RgMIka1zDdLrdNlkGR6R/KvkNa8mp9yz68BgfV0vwJHEDZsSrhmUbHmZ0QHH
WcsEb2N8z+9PDonzIqb6572W/pYI73x2kydaL2ZyJUkS00gdEu4HRx0WK8OtHfHH
PQpdpPFNBbK+5BCACkPRPg4F4tt4FnSe0KdAx4EYXliCtmv2b0RbyRsquz4GdVP/
ljPrcJF0jXO6ZJUcCE4RQ4HlUA+IoJtXPoctaztHKQaepkyKbnhlblgvhRVUZk9N
R9NjVBh/caz8NuTwlNLZa0pLif5MBftWJm45ynKtvo1KzvJ47DLzUZl4HhRz8F16
1cedyNqRMLp6AHfZChC68TR//4gL5uT+i0ulx43RI/Jm65E2KIw9oEwwExGDfyEz
V44QmAKoYz8t/AfCKkxGdxJQyv2405zV0efXGmYZNLRY4Wiwl+clW50Xr995wyVt
MNzWcjyFZmUe8VLovSBXy+EMVYX6B/lpla28o6wT8pJ2zd8hoHYrZcrYGk7GGrwb
0hzxwowyEfWTshIrcTZ20eKK2v9RWJGhaZtSTv4SjCAKaZqxY95jBUl1hLwM8+AW
1diuImRDk1oB9ylT0UZOaUjxwiY7CgMNC275XYX1gLC+7FEMKvLA3vmvNqE/IblQ
WGxspODggLVaYt+n/CDXG+ygCGumAXaJ6CRMeSVgqpsTlSDwcPCniPnKHtPglaZo
v/8pqLRxQGYLzIqz7UbtWPO9PikTKhoE3IRRB76Q1YV4ut8N0mFySiSQ251wid3k
55z0Yl6CMgSpRyVBZGxUxWSPjDp21d9RP/ylFkA7Sv8VPFcs6UqSy2t+ePFGh9AB
XAXNuKTQso4OxwW0gTEsa0DAS+8Xcg6tD+5E29aEiJ0Cgh4OZEihOto2m6qN/KHt
z+PNhUu0krncVZfUHLZM373tYojmgaTT1p1T5lUlVDaqg1EaTq9JStqrOfXBeDX7
+7OAy/dk2DhWSZJfxEobfduPaBX7Hdo/1ybDVnmuCJJNIFrZguryL7YrtlKG0Qwz
yKJrqhZA12jjkuR/EftZRVFUG/Yx2L/iyjGbtTHGb5w3SqhuTme7LFDGWNVwz8IV
7tZ8ijDVnNBTSwD48iz76P9YBm/UWtjgniEQKER1lhZnL75/UfDN4lz64xk6GSIg
eYEA0t47lttRuYnwhyV0Lps0VqCzZ5v0C0yJ0lesuZQqOfv3uQGF/+0VFZsx9bfI
+w9gFPOFQdQI0xXkKPG6py+w0qNrp0WKsfFAS5iJFVafnOp7sHLEHR335fkWzGFa
cHBjN5NojA8R6OzUET4cqtn3BVpFwpaUOu3POv5ysd08asV/1DLMCWfIQJ5Pj4vb
f5NhlQAFUteCy6lQYL9qbjDZ6nFeqq05O/q9RZ+Cefg9kYDJzAHyr2ccTpcJpFCu
2bqMS1XSGufq+UJvVrNWypQFKxSX2Ztys8a50XHPlvpFBGvnSLKIlkpVvxO/zh9u
fGXBEKj8lndTuVF2dlJDvwYR2bINCXlV+6/vSLRLD4H6KXDm/yeFNNoSClSsqxxI
3tDZ9QOlCVoT8X0azZGex6lKQanRVodzs/+KI/KxbCzhEa7B2WY4gDmJfA7Dt6ZY
ctysbeUpgDwWjkV8JQxHKOvLCsiLbI1IXJYXhi+K/byoyu0bq/Xp7T7HceYEMUFv
Usyil9BsYHRMG24I8xjME9ztU23ofq6qEhE1UN36BSCDyupgGmEDEO2oNDnW4EVe
yWNiueuEc3uKx2B03KFn5NuXF51K1dIfGI3Ys4q7ianJ5tTq5YuXh0CCwxf4re6p
3Yk+BQSqvYMX4Ho35H4w89cLyMtl6tP6Q+UlPv3Q6Od7kE1kD8H2xbcA9dOxsxTS
XW7EaRmiY7UL65gAFdWcJreePhmwIQsWgQb98Lzg912QD/V4V8h2oPmuw0o03gg3
olXs4RSlvf4vo8JFXghHTekcW4On5A/Mg69p9JYJobhEPQfuyk6iodDcEWP631sH
gkkg9xPVdCMPFiA9XMx7laSGD+9wcOdDlW2jmSzRA1CbGVLf0kR4bqtZMUOUQcTp
P+T/nr2dnU3YdAtzEQ1RAzBwUls+U29WeT4/Mn9uKSGqfoLTTqfZSchaeVc1BiwY
qyW5XNbOZhTGkvBnk49E4iDRgNlkHbV1FT/ICWqzh080a2aqfr7PVGxo6RJvtuUy
Fj3rrPZk6nvduOlDwNWXo05+uVg1SH3WEoSaNtaIA3BDzz1d/ZyUUu3RQpfIoWNU
dqCNqbxIDv5QVgyp4+KvUFQHNBhl9h/slx3j7WsGtAkM4+DwqCJflDntWYNtnt2U
HGcMex+LUJw2yzw6F9o0ssmSr4M1yPLy2ibXlwscTUydCjzYIBJPEpJFPvcOJusU
fA+SnxPgqmdHJKRm5Sg8hD7PQOOg2V9XV/7UHkyedogj2V4LdpZRFIlfC5264RGN
Lyb8AMyH2uSz4HODFkY4Vfr2Eye59nFhZ5LTqEyHf7ekF29tvBFhORXLdFugK4kI
GMe0QdCFsdSJaZEH08NgqNJQLuCGxFDmvZuI50td0LQUqqmw6eV+3GGD5h9KVoUN
Ci19GjL5c4EnKNs/h/SuSyZzAEJUestLWuAK0J+NnAjyM4eNiuN1rK41ZFeU5iE0
/CoKs52TVWH0QiyM482Vk/m85heZyw/ilQ+slz0Qy3W+RgDj+25SV3GjlCseaC4D
Xn9lg4S7usvZUlT2CO28m1epJSfrAj14M7VxroxL5VdpUz9yZyqGWQJc0HYFVjOg
q2z3lcAMGTX8D71XJL3oq/dEv+anxd1lbNVjRt96jaOfLJWWi4EVEiqNpqilmr3X
PPopuaqqQxmwrCWYTX6iByO1HA0KfTkbNLVmClQJvrIpd4l16JVS9Fx+sIFX9DJS
ccjUodx372IQBsnII1rIaNvYn4C2UGDYHeUsQ4emnZIw0QqMj98WeYXG8oNTLScN
CgjDxY3xi18+SUqAI+xCDcs3Wqww7XPdlAp+wwn3O3Mlk2LsNfppakTc3h7HqKbZ
O+jQDpTEmaHGmJ06+AbTiC4kOQOYNlLdBfMcs+Y5s2rshUlTT+NJa9bPuWPqqs7G
4Hp7VkxvBlC7A5zecLwsxcNkfQhx6uvBMTZEZP46y1ATkPvVWHYyBYWd7Ny3CEGB
SIkomFVef2TLrAhLTFv7pKttUxxrO5DGtQpbaeuZSbq5PUmyrkaR0UcP6iq5ALXK
03eTZ/JU1FBLuELf6z85gu64bfUqJT9BDU3JY4w4MFQQmrXc7mhySsgUqVFemjmQ
5PcXCivybyvHvU4Ptjemd5VPAOUk6cOo1793BMjJ9E9ZJGhLLdpVi7LMHNb6dS2u
fN0i68o27TEqI7iWhXYGEVx6/hGvkHCsH8iMl6qhDdsZzHvY6cSSOC8Q74Q2pG+H
fWpJGuuFI+amYUrg9oD5vZHem6r7Gyhd/xidWxlluJyLmlBVir1hFsiAB5RYbQI4
ww+n9oXscCz0quBlGZWA34cP33GslRCgmF6lpIK569dK4C8dECSBVIrXHAeU5WLk
Xpdlw2j5shpW3xoNNj+0BHJlGPtQb7HaGgBbr9ghoHauS0zY2PY2DGmhtowbpMW7
kuzEwcGkNDxpa1x/J6/GM5fVlGdE3g6/R0jLmWVDJiGFlOirRQeR7HUBPFLC88aH
itQOACGMSAE9R0xBto25UPu5HYHjFA4e5mMG8cDJVLcLgoCYivsxWJ7i0t98cG8g
gDNRVRG9IlQFh0HkVcRbmEoy/2oWJ0P9hO3QDRsz5x9tUfbHbmf0qSk4W49NvRcd
k+UrBjLhGeAg0ryH7wx42K+3sqSCG6UMJLXl/KcrjmdgFeTOxOCsMViQMEqA7znl
kirp9PT6llfJhTLFKvWv6d+PMgqm4ef5enl9cOOIczdTc6ohCegPKoIzmvzJ9CK1
8TCSzpUlEGuJx4wJI2zbcM/UTqQVWrooaZ7PA3fknaH1jjunsOrKGdVEdlejIGaO
GJEz8c8+QfOt7S3LKbY3d0Qynw04bbrQsAhNIV5LtI4zUgmE95ijl564FCIbF7A4
a2L2YekVAUlXkdkYzs5MYVxiMqBUapYZFVhQD+fVdSPtiMlqSdBiKS4kEC+b43yG
QhB4d97A+K6D5boq++boDtv1fuUACX5YdtvcghLGtcVMFloRZzw/BFteb+HUOFIg
uysoaLY5IeEBim8JsJ2454vvZ4Lj8H0bgbTUFi9SK/o82c00P4lQaZm3WsjiEOlJ
jientoVtSbv5CwOhW9BYQBB+huNcPkB8G9gK1ujEiyCRSQlY3WJJL1SJYJ1BGzdg
8jphdsf6FjY/owYTRvpEiNsbR6OdAg7XCu9afOp+wpBccbgZCC9a44IYyViwXpz1
bsxc10GnoWZ5E02S4zD+g9OliUS0dTQ3v5LJAamSE+Vao/rVdOew50uD5i6PuhJT
Te1d2LUzGK7lkUnH+2m08MV2vaPbomtHg3lHcz+CU+aJuXGNTz1eT9Gt/4QhfQkY
EVK5fHNb2wHPLZkSyHx+/QJs9TJR28p72MjfSCZffCRAi+avOffhcARvp6tNE8mO
bJx2tkQRtGovYN7y4KMi7ye2g1+pYohCY+RC/oImYMZmtwwoaopaEq96+G3TjEaf
ML+1dPQMh/M12GpgG+UrX2R+yAmU0ccYwDYslM0Rc6LOg8d6JI/z++aXc/ginATe
/DjxyEorU8JX9vx4Pdfehp/cKUzAe0ioCemoroDLrTKje9946b5HcoMKbaMDeSu+
QIUau1IN5FfVAK4xK5kNqHekqG2m/hY+3C3vhMXSCa3Ws04b1Rp2LGrYTQs9RTF/
i71B9Mw217Fxk/PS6rYXp48MP8U4yAmoDDy981CHMWethz9yE+m7eheYv1Zr8Di0
JucvR60MzZxfjlB/TkB4xMboh8JN98P2Z5qjXITbWFDeGi8uuiXaf2J/IxLqCQFF
Lw9Ad+GY5Uw1Qc82yYfK3ItGAvgEEmghgU3VMgMVBsTQg7e/8yZmx1wyMLppggTA
NfbGQYrkJN0t0Crjos5WZi865hMS5ihoh3SSIrUqxPAFcJAIUgQNPiBL686sSumK
t2z3AEmZzs1xFgfYO5MffDv8QUCpbFTES+Pf5j6VtBXhqCghTZKJOJGQP1Q4fBgg
3sRIOdNkbThvoVMqhtxzhplzWPEhQyBc4gwJdeOrJjMbXoyQwB8lb1or0nWynDxy
7wzFcx/mZvwNYaEbUoiuQYeJ6pJAjZtPEBu0T3r0XiMbUPROcHV8N8bqjvyzfp/R
+8KdTF3vPF0PEhv1FPKudbNIBvxwJI4oHkgY7MHVH/9XqyRpWP8q9fn0aZ4X2Kmp
P55KYy0wdFaOVScNAxqCdMIkfzta5142YzMmJDy9AXxN0uYoYivKbLZEvmZcnXco
HXlxd1NKtCRVZWTjgh01MzJ/Nr8H6Kj0o8heLpi/1Vsq+RBRorf322A6Zjtglbwn
5qcX1Xzpzt4XmIPcu18njaxwmG3AuGheuuEHqaIlekNZqSu1xEAvPiATX0gZ38Ss
li4vksbAQohb2pa8Dk87PnT+dW9++/NpRWcf5E2mFD+LoTkxBNbP7sbtU2V/J+K2
iTev9cWahq6z0QTc2Ph8DPhCubif3bYYcf+12m+7Yxzd3KgEcaRabjyn+blyEqmE
9eSdA/JfV7sBEQijLWKyo3SHoXACVZ4D0jmjgi4GglnROhm91DWwCoQQtSQ1e7qR
NzDgUYim43lCVH1ilitCXJKl2vLwDC3DYBdFFQ9TskkT4CgPjXDG6ggJwuidyD4v
BMFSY6Fje46u34PVCsySPQ0MT6JfQ/plLwoaWyFQWr+0PcTvUaPyqjLDvP/R/vxd
vspLC6+9Plib92LqE7COHVXfmBgJDfAhuMraXLBt/pCGN4yKCp94g9iczO73XtVB
T7KV6YwL5yH9c6jJNOcKdBc+DeAQ7k23HtKfjzcUArgoCu+CBkluiMqVPDXTxOGy
B3gVjC0raN+uROH6zjO0K3vc/3004Ylg2hlCYpkzRouveOWGCXBRRv4dzhqk/9X6
59OpVgM+KJJYmVnrYBx451PVt2La9pT2DzgqZUdVKLuJe/yU0wEh0DduAc23xxsq
YgTmS0tSlz/uCokhOOmGkG5KQ6ybhP4aRvCK/3RjyVrJJ1gies0PCL+3RY6GFStN
EG6BAATPpnuNbpkSjX9frv4spfFZO3lOkGonT0v2kkt3laPvvEmiN2mJ8BIa675T
LdmPiRrNY3ITGeLpjRxYsis969Lzhz3GFc2+GW2rVVEtM2rXf4OnMoiUQIWGjOXC
hKunBsHk4sK5MAhJqEZOM/WEaNCvPFDx0q46fLARTRVe0pQUQ2O2f9F2ae/H+E0t
HiBWvzY/84n8D/vFPbaK16BBr0CNMVDOXV/EiYoKBT8kFwCOBQi0qQJ7somVpCra
/t1QIWArOgomki4WzoEj3A4eONV2ZRfpCPbP4xDPtbFJcdG+ouLTjn52hZOP9Scr
3lqXP8KufB+lLTyaD3Tx+bhQ2Sam6Jjpfve196n1org4ZiPLNs2TCG71V3L/L5CS
lMggsaxXZEFukpfZPf8bAAGIBwsij7SCcLh9EzKaV9SseSZ9q+Gz6BbbYRVCpJyy
O68ALibeG27PPEntGPdMaw1hqD9C7nnus9fAAFJTMsgSpXAQ4h9qgy1ZSMzNsOuA
BWKf4Zlr5oUZiNai7K7Krla/jmXDcdUYyXY0USR/AoJwu08LkD5HIxCPlB6xb826
5If6zXcHG4KjpM+/Cg8Vsu7Ixo3LStSFGrbiR531V/LJm3swyBe6H2eW0VOkGjFR
7Q2lblbPDbVcSVDjVf2fX6J80jE2U82J4nb9q5V7ZN8f/S+roDIlL/F3mu+6yBRU
vd8TlCfd3m7si3Xj48MMfC0tFuL4PiQoTHU2LWRkP9z6+8SpAg5NDWKzfWHRGa/5
sdKAms0LsoVih+yRG3B068dJzBzRkmIc5qTpbpvHyujxOk/DblqbVWC3poR8uUl+
XFC1oMEutmE5aCkoVPuoHcDWe9a2LTokyUu1b+hI6wgNUnJhqXz8JBnUU7+fVK84
QX1BCedIc0wlo9d3qMa0m4OXKGELUHakS7eW3pAu1t7yBCJL1mDvL6ed4v85htLt
BqPpBIH9BQjM4R7mcbGkY6JsaIstL23OPBeEUe2rkjHZvmpukuh1lHYBDdJK62Il
j08r1fGkiw08lxSCcWtQEI2zopJoFzJwb9AqYsRhM425udHEIybgIQlndudXJUJG
IuO1nFpSTID3lBLlkYkl+oLmdgobVvAXF4mnA3joPNZ0oxFAVUP49W2+cFxqSnup
W9+B4oJvrXk0bZAqIj5UrJm3PcqxPEOYVwyt79VyPL3v4eGGI1G/ZTwlKCeioPK/
`pragma protect end_protected
