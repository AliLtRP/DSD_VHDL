// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ND9lVEkPXieJwknPxGDZx9fe0J7Lj8X9qDmXhz1hR3Oh1y84KWJFmnNTWHDi5EwT
cETJaypuomIGJsj59NC2MGurJIRggS1UVNANURmexk0H3+Na7p8sRVTAjGR0EFKO
8L19RWIniZYiXMf5JiISMPFdi8Q4zquSavbFdGDiTY4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12288)
XLsGQdg9VOaR9QZrR638ciu/EHS0wMtn2dbhmQJsW5ID6FKOzmGvi8eUuqUvyS9Q
PWZsmWaGSL4Hxv1JB8aljJJve5IG9HKHqJfmwO3cV53sSzPzKlawGHq68w8g5cYZ
OYeKyXrLIOYqJlyY8s1dtHDnBuq8yGCWbTiOVGP5PKD2Rm7yM4JG3Se93s3iZqGH
SacQxEDNOZVKfu5MLT1YeOdgSYkO8rfy6QY7lrSWCDOnFKKcLoh1B6GEXXOnvBC+
FpBnlX6CpZwOmfdfyGDHA73HT5PHVALeX0WO/ssPrwyRJanN1NUYam15Pj9Cxuyf
ohaVf4bQ5yjGGM5+1+OBdvvaZXQzDwKLUYMdBgYaK4+nb9Hg4TVXCT9y+7JmRd+c
6Yo5ZVWqXJyKI4jUQkOL1ubC4hPvwI+mh6aehhcPuTzh/GagX5Ueht8wMTEgZw5s
r4pgdStfBivOmze9Ipg5YkIgEq0/Ol4aKO6/7Gr5jlPTen68+6LcPU3KPu9qFvP1
h9cdcyDmL1wKRakBE39iFUy/UZ+EPedqdttdSwjesn2wWMByOLKrC8wngqROr7BO
dQbY/WNNoHVSHSjBEoZunZVdvyg6UtZBTggtpEl6CGoTw9N3U8lbI6e6t73PPugG
sHKQZVkeGX+BgsTWoQkn4dneS0WT0XY+EcJWhsehC0uZxpbcXf6P+AhP+cMHXB14
xSr+iB40fAoTmRV+6ID5C45poOmecA/5Fsdc1JQIa3dGxxRWPsdZ/fXECk3BUPGM
8HTERKopm4VDntgyzCzvvfO+y9VxkX7tlSjGtHbv/wReWYwC5OYyPg44SAKb6viW
vPTBvCvQBxTwuRmVtS8XYo/Jfj9uyUAMMlh8TwvfYu9lqcUhzkqQ9MWsENL0SRkk
Ytz8HfDvLd2XgFjQg6kaScTo58jYOxbSFyvIUyyHcxdbBCybatO3Ir3g3jSxZOGG
6U0BuH/853602FOkPs3DNFvl3gL8W3Ub3lGCqJ8CSVqL/VEgKseesEQEIpXPKue2
pddHJrbcQ/kQgyro2MXJprDQ9DMvpjxmSqWjGQ5juFKFely2agdJXWzbINPbh9gN
89M35mai6je3apGD2FNjD+9knvDhQM9Qmlb5QMG766YGWO8FDDnrMHz6muDtEAWA
aFOjJpdc1WXDaa4QN4aIzcvQKWltQnfy8eLoBPp0Er3Q4P/aBmYbTKtoAIlVC8BE
ImzmN0FqW7erSHCRAQ9MJeK2JK2NRrF9twPrTH7rNJRn7HmExPGuD6kt7e9/OcnT
5owuj/3BiUXvf+Kmr6Q3syyPxE0JeI9vhfFScbW72QxxKWCewzYlHjww/ZH1egNu
U3ifhNxu+t7skeGFy4VDG9WundtZhZmE5/xlwmqEqzI5bRDaGM41WvLXEcM67QND
AJZL9odQyhgV14N1QWFMm72lbEQ8HNuw12iSiAnits+A95eHeVHWXviqfqqpYB6j
vfbQb4/PI5WQ+yX3UgFtSnnnBZpHGWDzfRJhwJTSqX5ALJxBCm8TjO+PGS6IEvUj
OLs5JofWNHwHF2wqHRtCq7ctomUW6ovl0J7b3FPtuCwnu1UfGJT7lklQkOnoAcn/
Oa9wmSV6/nQmX186+KNJpGkDKHKVpfGJeIa6XGqTvDvAzAxxU0nfDzB6BCqMq4dV
i3wsd+xbyt3I1Y1j3Zb+ga2rHT2mj3RIF5Ks2Et/oAGf5kKq5J0CyY4Yud809Fi4
0F8v2UAxQZfs2M+52utSXOjyfvrMagOKL62xua57T7XhxntJIrV9mDZ1FYpA5Vu2
GVD6OFwb8NR4PEH8AmJz1MHO1pl+63pcdrf2vzJ4U9QCtMI6wm8Fu0GYn32NdAvK
Uov4iXo9bRwVxVgyFWcyMeRMCJpnvRvuvxmTENrnA6ft0iqUYfmAAqYMJhHK47tL
r4xpuJ1z+WFZO+9WqBkGguWLfqqjyKfm/l3caxKYFkYystsCSfSNcjfPog+xJFZv
lUqlHBPB282jkFFForByPrZKNFOzz7K4yVR/Ms36SqZyF+bwOrY0Jx83llLtE8rK
c6Z0gF7RAHfdOYx9XkPDjGWdB9aa1DgKSLH/5NW/Usz55y4hIp5vxp/YXHeGxeyO
DSmtVwOaXF93PTtnbInVt3XYivXpyTd+PQO6K9xHN1j4QDlpoD1fD7SM2qxdHYdn
EsTGrFzjmJ4l0H0zJtPqsxr4N19Lwo63DJSDjHWOBLdJh6Z56VbgYf5wp07wM7X0
60lh54RvScb3+CCp979koWVdQstbaSTvbg6JY4TlOMd21YGsfBd1/2ihqbz+7lhe
+KKDTyf4N+4ddfJeGqq1QvSjGRb+gdNn/g7a01mBzCCk0dz5/84av0aeR/LAOhWp
iokVXvnmp7t83+kVtvzM4B8FJPHx076sYWgP4wjtbRohi2Rstb92JrYXUeUGvPXn
SERZbMOV6oE7ShkEhuO+m4/Ytb9i58H4uF36rvHVKVLkUlQGIt8n2IDkEs5Z8PPP
sCJq2+h+TAf0Nr8O3xoQOb3u9gl3t1dDpSOoIGNRZW1Mw8j6XUKzQUYrFqeBR/Sh
qG+TfYh1z0GPaGpxtW1ZGlohgcVw5BgtNJ2mNd+H/G+/PPA4acwDlXBbkn8uRYdl
vda/UOtshC8FroJh9QX0GtxZmkD54di9ivrLcndIsRpmcIYC9uNIOxcK2jlakHv5
g9povr5tK8Dn7a3RSnWyfu4wrRHv/FAu9VuAJ/krcYWOb7bMAOKiyHB/k8yuauvn
hw1chsYqb+4Y5N3XG2xD8ofrSOfi9CaksNM2AI0/vfHjLPxJ8AqOeyn/sgY7Qnca
xeQ0RdSDcEjpoZTLytPzzb/7Y70C9tgXgIBfR2hVspLTDi0sqX/JDswOIsOGbGUp
mWSPDDpdIuJ3PVWo1pxOHmb8mbRH9zNceSldm3n9h6dtDhuc1JIvALVIGK2kJa4g
YJGVKI8+/q0Uj2dihR+dculdJuDrOc0kA0h3/djQrvhipQNlodrDl9fgW5Kh+2DQ
zzAmmY4cOWEQBeewuF76J5mq+IY5DFnLvGgRll84mEW4tWwU7nu9Qt0a9iMOsn5R
+i4N6KsZO6OTEQRdj+NLDRBD6KKq/gxsRyQmtanISbQQr1Tp8ZcrPdv+ypjJiIoU
uuI5yteZSsCCo3UY1WhCXQidzhi4h4nz1TiKZP6vYrD57C9/JMK9AGebOGp17Okz
tdzM5nLGg+oTdWDPitx1VmZHV7pTqGTRwzSlGhz2CeHnhgkxvnSlE3pksbtGpJaT
SXQaWNBCymn9YlYSBBRwy5xvuigXqv+bZfegCEMVLR4zJO3Jk5Yb4KBBNX9CkdTP
u1mMQpdoKx748S0swtpW2n8KzgNASMkPvZnMAsnjROo3dlQb+RnckHdO9e1WXjsW
bN+4ov17bO/w4WKKj8Ow5eFuqwHbSUouW8t3EcdkqK8GoT4j2Yu2t8OrGcomJVjJ
haQ1dMFE3crerIGCn38X1qjrX/FyLG1Z7TZGR69KefdCeLMx9+wHG5VoXkZVdlxs
SM+gpn0xjrZV5jD8h+Y81neeTsnRNT2eBSQ45qoR4GNWyfYj5Qm1+cytjLZDY0QG
3ffTJUpuhgbGnRlogNMAh0x0p6oFH7zrMIpEe0XGyLbiN3iZ+oP/Wg7ywXpLmuH/
+2YQPoK2ICloKFigQxbXeQsyglOuBNw+hq+yApQpGJtjf/95geeL6X+Hx/SNh8WR
O3OfsFh7IQb2pI8pgzu7tIcAgLqM0iPbuGng/6X4hJjvF4j2Smf9ir8+lsEMrcFC
Bx7YyLnz5Ns+OmCtTlaWlyQWseSeyxkZqKinter9JUUNZxLh+2QGIwkg3XovVKsN
bAhUvHBfeaurjV9UMbb4YanDk9DDUThF8vwtdZmyNdyAGlr0kRZVveGuRAL3my5E
ZisO2+JS2Yi0B8N3UtaDsYHrTbBprcygkVZhIwg8crJAtz9q3ROnQBT7WyZWMeAs
MVfDvM1siouC+TOIXpxD8Z7+BMkvHbZEYjQ7sYiyeyczPwXiVuvhp4GTNv6f/Hns
ypAXDuI34KgT1Q1Fz3zpW3JOTobBnT/eNCuw927v68CpUJUduQv5qo5JBpJhlBuC
R5tNtQs8o3C9SJczaLDRUPglMRSCZsEO/RK4WYtlPOeCyz45KtWU/sZ7K1hNiJp6
zWLeQs+4jhZ2WfU872v5cco8lUexcyDo46zXRCAlcM6YQd0OYyebUUxZKenSojhu
LMPObAZhVky7VfZoTaVRGLcwfwXaB1GNqHOedO0AjLtFGFrG8ElGnZeSoTjM/QHq
1bWCORRdVOwmes3s7vc7ai64N+AOCXhIeqSiHoZnsyL9vu+FvJWF5Dhi2yVwqIEs
oZ54gCILpJ4kHJ8HVkxPmRVkM6jdvDrXAsNiplxgYTLwoIHcr44DgGFPzeEFu6uc
uT2Sch9kQknJUmpEo2yOcnDFYvckO+LyRbbTDWnWmYNhdXUeED4wrJ/7J3r0jbAN
5UZLe0WslB+1YZqaLrVs7qFYxiI979Yk2BV6YF3lwINyQ9JPk2/dBF7MRFLQRmV3
vJcOeR3+uuWqWiEmZdbDXceaJF5zLuPpK4CDxvASgi5vbssIF2l/zrxiO0AQ+bOK
78o5ut6BPsnXaCXQVeBn7tYhomUC/f5mqu0Jv1STxa265E+QUrP2iAyXha5c95+v
uExE6TH2YdX/IowXVUI1ge+/N9TgrNhDxuSR1wUe55v1iutLS1HXN+t/BFUorkuY
oB9NKdWPzfeS4UTXuWrJ6G1kinKV4Zv47zvvDT59KDvOI+IrFHqXQtmT5dNIT90O
vMvVT3Fh+qczisucBBo5u9/XuePqlEJc0KykQxGdDhFHtXqF2mC1nYwwjZD+tVd/
H+csk4AJLKME3AJ7d2leEicoj0hZoRWSgvWmdQh9i1zQjBwfUzbuB7nxyT0t9L7c
FLCgBBSINuq2x0LKg4o21Ljwt6QgdqBfh+HJCJ1Ohh0uNRmcnNBFI8Mj5kej4REA
34HXS9C6+fhaqoocAWtlMvUtc1kbvdvkLZDODVPVTCUHJUZx7X5jRZ03I6kDAJQ3
1M7zllG0UPaneLGWtQmUiN6PSbGnEGDCxvNfUXGuAhnmGqRGc6hiwipoCdgN2yKx
ulyhZvj810Pustp6iOXvaKYNdqF5zbl83pTiHDCSThpKLnWw8wzpqYS02e36PsYQ
YkZLZ2BaUDslv4GNZfbZNVIGTFyD3hb0xOB9TNtNYhNo+YQ1iSOgk7Cg7tK3BgYq
aEcNed8rlcCKFeocYaq+hKkE4L9MgEwiRCm0GCRkwRhbhVSG6gg76zsnC1m0U8te
wkMOl7pe4A1heULAvOaaVJE7gRNR/KS1ERc10rdVE+9scvvrKzzqL6kDYNHh5+7G
GTiFQg4OWwo0HYkoHmNY7jGqj6hJFR13W/pQrMx04nVPFcTpSTr2a/QocehB7HX/
KIkbTtjcwLQfW5jjhmHvH5f0KxYIoYgP709atreycHAdQz5EFXs8RvfF1pn/hoyP
+mVOFyDQofKtAWy1ejZljShdQQI1WWp6NqMLxQg0kZ4oSbZ5EKfzXDQXLJjvh369
z1hs9prgIA6Riq2zawiNEtYeQGaH4jBHRYez3ttd+UAuAzwIxlWxg6ippjBOtevG
lVd6psuqA4gDK3oi0s5/av9y+kh2gIzruvt5CFqAK02GWT0Ly6s2sDNJKl2YWD3g
b1ygN1v/eUfKMCykQ8+5313mbfrkk5y1OrJqZt8jJfa7leBqUiXMwvdoAnyI3JBS
Yyc74UIAvMYx+0kprfMdox/tON4gQsscxiEP4VYNzYBhtxmuIJ+GoksC2y3XhcfU
dw9xVPV1smXTiYaY5xwYaNDhl3yX9d9lcLsbFfDgdiOngN8ro8MNsARQ16NcJ84F
wTQ18BybWuA54WCDNmLqtseGk9h415EJJ1ycvpMwC89Z7cjQKTYEE9Np21Sw56n4
mF2VOEKdf6MBxT9b7JnzgPI6w/9Tz05DAoBbLSZ/xl9SUs0L73PWIgUMMuD0BNaj
Pk/UdXi8B+ZF9ETPU3lKcV/pR+0AfkfV9V487yEwbr2cCeJkhssTGYqO38fAh9i2
qjmWx6ku33rsPUmRv/y7OjopOnYGQJHMuh9mrkAK+GAzHa5LnV+Qq79XXTKz64Vv
uyhcfp0gv3hNDGhEKFkfKOHXN2vdiJ6xZedY6LCsNYTTccDJh/uS0Iym5svolN8X
uGWwv32L5+QT025p0WN190HMpkhhw+HM8xuIp7WpKmWj1wtZgUZ6aEZNamytxvcl
Dal9MYdNGQPNURxoH3uax+Q4RedALEpW3odtLhiCsxY0tFBnUSyb4NwDLLjEGC5P
Wfky7F1CZb4pvtwvi6TUcIbjJdPDYuOqxK4u8TNbGluANjeCechUHxmDz+GDGjc+
ClztgkIxfgaIvQehWn+wnkBijm6sBAOJtkFk7wSRGI5qUmfbCza1NxOr5C4GUx69
EQESDZ3+l+KM5tSC/Z0SZnFWPPVE7x3pkiwRdWTiRRB7Psl0cKDe8zI5qW9XOl63
xPpY966Zl4RfOflOHWNd7cUUA7/QeOFC7sM7lVxCXS/gMu5bCZfUroludhuSY8g7
CWra5lfZWps4RxgIF2EVD6pQdh6gBCArdtl/YFmDQvbWZdSa3PrjFagDwrAZ5HnB
OcMQVmw57NT4zFqH+zXJoQsF70K3q6jcJbcV+ia9Horn9FlwtipASZiJNIxhP8q9
ww/90P3pouM3A1qesQgXYgTEXuZJlZUKRpMXd5Qv+YOidfQ0pT0BUPxif+sXi9Zr
IMZNJXe7q2R+5OLYTDMtHckEzQwA07nrEYpu7lfRJKLwaT6kaUjoFdfOoi/KzR+M
mS6zGnC+2dlrx/guxoBcrSE7iw25TVMd2aEjcXojHcG4fg+97ciu7+AdWUxayjLR
oy26emF9m6WqiPFqItSJ1oJ51J5WOsQVm2LluI0Cs5B0AX5LcmVfmK4Re0yryhdn
o6GcAGPkevtIsi/t21H0aOmjzUVNBq07e/OBkUW0L8cOCC3qU2Gd1jCULGNVUC4p
T5o89QqrsULEtKAjsU7Uep69fHr3mm9FyowPkOvt0gL8xBFo2Lfhp7uYGoDenCmM
fqICYgy1Yt2i8C2eIV53tkNy6aX4p2ZMXfmH3YSLrch0vH7w/iUvf4omLY1/ucwl
L6vjUePLdXOGJG8+Mk8wWsDTzzhnv2fxSjSvj4aoE/lx1Lzt8RdPeLVLarXDr9kG
MQdNHRfxryY00hvGneU9xKNqlIc7qDb9s0Qbe6WGZNqXU3A9T7B7OYgs7aPzLHEu
OJEVSk2O/tMSC+46eVDVZ3L4A4lvMJIKv+xO2itXPici4YvPM5EEllDZkKhyFnpT
bU30yaz02z7/bnMXOTgjmp1NnFCo/EC6ragDixowqA+rMmoYPDSmeJOg1r6dkMxK
kkXrCIy+uzJTugM6Y0aikPf5APnm96KUy4TnKRDqVa7Ar2qSFiJ2eIEheXZIXno7
5iiGvezPxm2jXwIWPBx/M875kAN8R5b9QRaEi+52to96/tiTsqaAB4G2XCujw7aM
qZYiuiwpOPvJ7aPRgpvDK+E6ENkDwe+5q+u2GGpSEmHKti34QTuj18yx9tU6g7PU
Mc7pvbGl254Nl4STfTDpoFdRMvN6J7A5xclthp5ddCBprn1MEI9zScsxVt+yDIQY
Ztrdr+1+I3m8eMsTtJCwY/2HmJSMuur4z5SxzgQW8UHhcYCF2Xp+s2t2Zmba5v0S
LxBVL9P+Sx71qXx2dkFARLljc5RG2bcqHuB97IdvPS/PJmQ8SqvReBBdvYQHx7fi
Icop+VewJvh4heotZ8uisgJfKX90Zex6iBwrl1fjLWxNg+TfUPHrFSi8ibWoq5Lh
7+5R53CAwkfWtXO/lkpCm5gLYLMXZ03dMh9JYIYyAGLn9ZuRzN4Zxj5v/oj1OLz4
X3rMiZpJqXpMa1ml4RiCtB6iXsnuIOLgEXdCKeqKnBikXVQG2HKy7NlDGg+MIRuh
h8PX6g5LlBK7B8oJ1PbKZklympHJpudp51ywGE+PxyJr5Pi1/7C5ddwskM6q8lVo
x4KYQYVkPmAG7ejNz5kFqPxxGXD82SDtNUmp5jl8vpyOwBLCXjl2NKd5WXPCd2EE
Qa+O3e33JIoaVZzJRkoJleKWmoSAeAGzAf9+rhsEpgg8ItXO0Nkl1cudreyzUooo
iqoNuthRX6ve1BcgabgSOkA1p52Fsx85fEscmf+JzUwtk1gA2qt6khE4o8SBdbKu
A1fXCEphKsdxM9m+IyohYxNZp7LVNHw0KRblyq829qMyYW0VBmqY3xZZ4Zysg6kB
ZtqeBtOno1xUkww9RxBA98y5EoVFt1RddyLS+RAmY+oKMqU+BI3Fbu33yHUArkrn
GL2++GUkXB8WT5FH9vpAo9kALtFRVc/AvgTqVm/c1H2nEMTp1imo7LyNmKCOpQf3
fVjUhCsQxHjie5jqlm4ZEJpnaRYjOgrv7WtW5PevO0dMn35nFFiP+qKJLBAnKQyB
vbEsayndIakG0IOAeNjmY4jSc1zMX0v4oe0EQWJERQY3VB3focxUAjkUDaICvW7H
Tq8AXNM3BrAmAZoDEVujmK4hQ7idOzU3P8vb2SkkLRPKz/unFGDj0JU6KXn82Km9
7RIKL8Z3sKeV5MS3VOd+RnnXjJR9Ew9wweXx/denfWIISQp0d12tZZa7+IrTAL6+
11HDvVH1s/VJKV/NJYOl+r/7GIuldQWrHGabnY7f1N82gFf534+F+/X+vESNrq6+
OvFqIiD7fvJEe3grcNK6xH+1d1BTFZ8tG3dtuUAHcLdDMA95KjLchAJtJj+Cr33F
FyJUDHIRE2igeyMpLTuJOfapQnGPTR2IA8q35jKwSHQHXfeLhZmSWCdMgZGUrcsT
EsQ+1jpf5OWezm4MW6CoQBVNwP1rXBoYqlB68jcMyvLspt7DamzEtW8Gx4S1WV5a
NJ2ec6La+wIIR76m0WPn2DCs6yDHBfzAJMpbD72rKvMc32moXkFxIr1OdtSv+zlb
WLhlno+yZE/SL2LL+Qk+FRNuSVla24AaW4Hgx6J6L6YGf+utzjxabKN19iZnkO+P
Q5MlG1bhfGSeILxjEZwclYrrIwCpKNXQ2HdBjBo2VbPanZMLOZVjGPbi39Pdjsw6
R9xwZoheFRLQgHLqcXKp1B1QLwZDNDFv2+Cr/F8aanaqrSiHB5VHImymr0yF1qpX
ub9eUvjQoRv5b5vfCuhp1LlwxGejq1fMDr+20aoamY4mTpBfPhJJ5rYke8YLSex1
w7AVVv1JQJfBRI1h0Mex4MeQ2MfIxWUpDJHgAPNmd6K7CWvG3acGUhxyC9yG1yLP
UVu38cUIKE40+OpdM6govP89Q6WNky7fMhXA/e8Qc4OMDDb5UQstihIl4zcNZwzX
5sxf1WjFN8GRkuhhFWw3ESckn3xRCgRzL/FobOmNubtyRBhggVP71gXtryhtaNqx
XYEUdVP2oQIyHbyzHykitbSbqLZW1cAWijpz6IpIg4RRgbxzhOj8SnvoSNhAUhjy
WSQCEonhrL9uumleUMSPJj69H/Z1ZqhSq5tHh3ixcVwA7KOcI9OFhmbz15TSchWL
gKv/XI8e1yigFxQgfxqSdV8S7Ufm/eQXjpkPrwLWad0HFMfQWZ8YeO8KJ+TOcduv
4gtjKoa2C4K4Kbz2H1IfRSCFENkDHuI1fKBdDFT5qNnS4MEfiDeIz1MOoic65nWf
+O9vScU7Cl/TMaYAYLa/OfGD/WFis+bDLw3nsg44DxXhYEkiGHbkB2AlBvWXkn2C
Jkm7V1I69NM7kju9qOjvhj/a+iZJamrjg6J3rEUIPkXTZorpIvihBly3JupPmDXK
aRSfGtKwylSUsoFdf8EUyOUzkoj81eMerlHdGVInzvy9fc4/QWMkNus43TLg5uaR
v9CRhSqvzrvk3coy+VQ1KjuNTQivqvM6MlD2JLATCc2UTwP/oPZUjsZwFkj4hlW5
mRKz3NwCv1Xzs3wWydm2cgr8y35tCOu7h5onM11sMRAwMrluNvBXOn9H/OsQQ32Q
FQz0syavUXlB5XBY/8BP1eAD1z4/i67o3jGxvaSPiMo44ytjGcU5SNzP1Q9MTJkA
1PX7zutV+CupppP33Mgkkb7rokNWSo7Sl+6jsys6IO8WOpgq31JQZoGf19xPK7Rx
ZSu6E4qNs7g60dkSh91Q2NRMCovkXDNrG8LEE9H+cKheSyRzbIR5IkqPw/DjnHiS
ZWQT9RQaCCUhxfsRon2Sl9zY0CRvzuTrGMiJYzTL1R9nh5f6t0oZSVXxmxjcKBnN
ccn/Fjr7aLthGi8helbzxdczg/1+sFG+lK0ur2uRk2sPzB2uaEqynSuH2Dt8aq8L
lf6Oyv58MKHi9H83ShfJa87o+tLaYIwb6KrC8fPpU/Rp3Ipzvvwhzby/v9I/f5fC
T1eLGIVX10aqNse2yI7hfeTbrWs+WfYMSRT7OYQRWuQ4ChCWabTAU3jQkT+Qiqp1
EVnsQ0dj4dEhsts/QjXjFPtpPkdd7uSScmf1F+0B6/NB5oQH8GKqYSGEHnamX/pe
hPBUgcDa1Il5z/jhboCHPfEMeJxRZB0mkXc+P9/T5l862LXO72QruPF0lWuj72vB
SKktd09EfLQ5ffNO9UGrcPGvNk0r0bjUITwd/QNZ1n3Igh4gLsmbCUEJqifG4rAe
bq0Bw1L2lZz2AQLpZWvkW6ur8dYZkyQdDgPUiiS+GB6TJCygUA6xvFlA8/JElKyk
BKAJjEIceYuAK92RVQfN7qcJKM0sYKUc/6hYP+IKfuzDqXJER4HbIM1LtAAea49B
mAnKsGFryruedJSkg/oQ+Cfw5+66QN3oYBRZ2L8MY5qRInhcYzuwX3MHnA5RCAbS
yjAEx5RzazD1euVdkYfpYAHYzvzXg/hNJIjbmj2opiYuC/fO55NfB7eO/JLzVtR4
+7lLio9MsENkvZQnZYPhy+0GMXFQbwf50wuM97PsxKCV1u4sSaEGuFvxGobGErt2
JEaxzGLoMkQTSyOV13681/fGZ8YOg/3nkJLyko6ebmiKYDssYfbTcRkH95drbdCH
7mCWMfqLXfOWgxHHqdFF+iuaId77h8K+2Cegmsg3jr1wikHeovr2dDaLWeEEblWb
pcuD0rMnbQrtlhTdoAR1p8lSsu4KN1l0R/gMh6uAX7jWhVj6qDurmE91fDvtZJZW
u1gGboYGQMMcQbmJa9EfsvttT3CTbCEpI67CiuxQshz1jfdB44PTiGkmzAPEFFpk
4KJYegduIi6KzarmleXbRPjHSzWUYIuS4UC9olgbSHSEzswJyxPYSgQIpMD8j4/v
1CpPUZbuxYyZlN4NTKnW0C0UR2KTs33nqDU8eyKnyRX2Pc5CN3HU1gYJx5aTA6Cm
83R/i+QjMVrVfHD5UnrXCZYghsWJxSIMN9cDzgrPTX/Yac9x85Msk2VrZOkJ9O9V
WEbuYy4YGTmEPPrehfzRS89oPrnF8Ps2Xj6eNB7/XxL1qdb7+Wv5dZbfYxehkCAM
AZt//+AgoeB4QuMgDLrxVrgJzMZXVsnYyfvA1Q1XqxcN6xOy6IKu5DY5MEv4kxlN
rU1mTd7yFSXAcDe8EX+5OERr3qZAhnb6+ZnKSQ1Fh5mwvtlR+N2Yv4rCEYorkbzr
0BIracU/r3Prmo3CvHhwawnSo4dXCP0De9t76ezQpMSm1Dp6syEBEEE6P47ufRZP
HmsnT7z6suB9soQmhsRqG1YTDLgH6/pT700QRXjWchgNZfzo5s75RMF9unwB4780
1V9MNQzLY3mI/yR4SJfaUuG7VwwEEZvTWMxjDhWy6VONlK+qdDtpVk2aShxMvApe
N/32OFb0tgxjFMgwvrXX5L5UQGktYEnQuKq+GhXpxa7OWOZkTbrhzlzAM0ZwfR3q
KvYUiyj+SWhXwaw9/lu4DrTqIcj6GfeTtNLAVIsMsBmJrpFYuTzHFBdbkm3Hu0iq
m0yk7M7O/XIE+KD5YoA8tzqbVAODR5He0sWtrvrsayytOXUhSI4QhhWtqIxd++JP
/SZE9Pa9yzOa4URVqOP7N+z/bevYaVnAb6xqvftIpCrIkoi6tCUp8JDUknCDVmOA
WAvpH/QokncdZGIMLRIah7W5rpjKRDhQ0BT6wecAaIxBvuCvkwUX/uhoc+q67jlF
rdXBtoxVULsdkTsWAd6KgwOa2z8Sj9kgIXE3laZOzNuvKPdFCrxxXsOF/DMsuCT4
9SyvirOiCEk+/kZEHopAZKVwRqccRU2uo7C56sKeNMuh339rAT1jbGFX8rAJLu6F
UAJkA7M2W6eKkug9EQ4gBCNxSosJdkZ7z7OmNYUMPkq8r85FxeP2tOPi1GQkHXSz
fztl2cTgLoTxf5o5pnjRcjPHcqUPIJ44nLgzUcFL9lxtDQIhUXo1CBRa4lrzmMBO
sCmjKyTUnzNJYoOuloRmEH+HIwTTaFaJnyiuap/cJm1jik8mb2/kqTBxUuOirH1X
k+aXOR8SI+gakiezFVXfsorhrg3xm+YPu4/RB69MVuS1LL80nJji72DVsWVA4Gih
g3o1z4Za6Jxz41iQ43kxaNnOIU2d3v5W/saoklleTpUWAqEm7wZOHQzsiEx8r3pI
UNAcufDYYJf6fItZSfmO4wtsRjWPTINgO62S4g6qF3+senJgBHEM7e+Buvc0ETYS
TobBvW2RhzeG4RNDAyNTvaAKrY+ZQHhr46UXe0vW6SwzwH8Qt+dUujITFD1gUfmF
AHYtICZpy4kf2Y7F3H3SUOgaFFW0+5+vreLr/nVliAR0rsDmMY2ow4qJ8cvC/oJy
CxZJBEfjdXUAAtEYPBJlt3yO5s/VjlqdG9Fv7m/YcocnEb3FlXHCscaDU7A3EHdV
ImcZx97QQ+ovldxsPTwb6wiFCo//KLHXGACyWlf1/srEPSAerEr6Z8NNljpMUk1Z
Lx6gqyXVUwDatCSXC1nPneScAyzYdEyzSzcdw9DoMNlzBW53Q07Rs+joy/3gqBcI
S38I3CxKVG6J0oSBxuXbnECagY21ZqVEEXyeRZVbMG77WGnsrwJ7iBtIh2Vuo6yw
MopnZq4rms2BuGgiT4ObNfsVbnv5IKFGzDY+BhUDF/pKgLTvFS26xFxvhlqtSRjQ
L+Pfbm8teOrgsUg7ZW7x+9loaWauky2ldq1L0Ua6CA8hJg/IihM5NVHEhAKOTv2a
ROZGehJjJbIEdzuNqYyNKJ5yQarlnAG2fIkgQDEeC+Lm2H54IgF5zyABTMxUvJjT
9ZhrDI5LsZ2bh2HWpXCrpYJoSzPT7iHjMz5dmI5w8kBEgDmmeZunMdmzA7tkyGlO
wF8E4w/pJdOo2QuPR0ybbOZdvwSbs4JbNl6Y4qzwr/PfW+GYQg1cTlErfPLleObs
Xte+6cV5Ja/xTir/3CYKer3SzQoA+JogKfNj6jjheKCD/daGgYasBZ+1Qx28+1Uf
PrVbBMjZNZYIJ0N/XH5EFej0IoOkNJud7D49J8SIzLcXTnm/QKnCxoOIIMtoXyUg
kIJibs5fK7HuhQMN4bh22Z3UHb8waI/fI12fJ90XyoAAuTVtmGNyHgwFjYCA8LTD
Z9BuPiZt0mvomw3P0boVjY+8gz3AVNnyNR8/Gn2hNrqjsubzVvArVUlcyot/6SGU
Sl/H9/jRMhoPitDb0opoktvEp8rT4jgNZpypc6n4epjYWzYijoYM+0xqJ55dgvrL
pcfcwLzuAWqF/wagco9eY2m2PUaSywpWPjiVm1n35NRnnJqPf9y3PJpQag2IW9Bv
4oIy9kpYqgfD5vSm62oMp+XGX3BotYA6k3aiKwoNn5npWmDcxG95N4f4nYXnybGN
dAuT3ncGU111NyfH+uAEUiFpFRZB9Y85r1zTF/msQvR6l82juZCKF9pz+CQ6PEzq
MwJPm123TBs96jDZ5tn9yuz54pndwwuLV3R5xwwQEetuForkU7DVsc9xIVw3Ba+e
NLdApxLqQoduOo0SOh3uh8qQo8kebpITA9OC3LngHlsVcMmyVO/8bzXRe4eUOZju
02Ul+yVVeOVZHlzvhPbht0dSATkvollj4dETpWEeLvX5dLwEHreeqiZ7O2NBjVJs
gjHBwQoEiSvzbQKZC01N8VDA5fueJNKlvh2C8HCeCqo0GijPznAxVGBSSheNSJ9j
oOYCpRcvmHGL12UZOypidnHkPNW4iMm5n3jef2QW/cHRHrDh/IiN6xOr1qVDgjZT
iskNuBOodEKFDvuEysMMInRQcFbp/tXOdgWopXsrCQIwxMJevaqZ2vTGS2eVGlvV
0KRcYZKhkG6gzSxiUdKKUkH6TwP/V1UVD3jLQIPPoCn7klC/DRbB+b2/GUqZL+q4
nJYH/TnAq3iLiGFD+g/NLWT4C782q1/HAqJ5xINu7XOaHmo7wVsSknJ/dxi3Lhjd
2+E/xwQylUEUFZB1LJLWuflDslI3W+csf3we+iKuXYJ8apIU3AUd66A+9tw0QhJM
q3BajMB+NQqSRzbLtS3QTwaDfgzZHrD8RG8MLnRIP50d01hFgiNajEPI/R0Ao3bA
61ma9rf15fct36naI70id9bkxo3m9YRK0CkZqXFOVxokL4OXrbMF07hZVo4etvzc
RPWgcU175CIlrDqUneXRMXsU/2lLj8cyIVP9knI0cfQPpsCMMAM1HBHI5maeWx5v
22mPibn4Lc/8XTxZPZcqy4lNJQ2bUc0gZVaY2ZFwjoRDvaNgN+cCuawDt9jM2oKK
aUFxR+bJTPgm/UpE0d8IBHAkQF6ZuZNMx7G8GWQAaMEnxmpZLQhyfAG/MWb5cY3c
TbAFRnkMlIRM5EVokwgcmy8eYSYAHlk//uQRJE2y8yAD1NzOC+b3UuBQKiI3cMDD
zBuJzjkNAsTwcEb6b3gmbmicKR7ydnT3ucjT8xTMiUHoi/W6BR7/aRUZ+GgC/xOF
LfxTrvCRcBTUej+yOmgIeE3pNKbqFr91KDRoiYB4VF8gStCHSysyPMGQ9ZcE6Iyy
NFYtmMe54Rn26k0QG0FfPGlSxLyfq8/M1HQ9NIx8x88wU198VzcM2xDHL9reGAPW
2pyXd6UhsDqdMaTO01DG6K2Q1+dTRPqzM2k60L6BFXU8VjHCsRmfVGytHNS/Hd0s
cY1n0rzU4FkuUBu7rt9oUyqdsCRySPTmY2QRxMoTbSeYlPTjOmSwFJhSAJBzMsyE
74liXxMcmHSuNmBlJhT+5ok0QwINT4QZiLXnybNwtDEXz9e1nEsU07JbBuuoLfvL
d4u6JDlNDh/1Iw8fmCbELpqW5iXgXOHEABqzsdl8nc72PaXjTC5Pn8xfA90jzwz9
7XqkFmykA94n6KAWDSicl/In3Buh5hag9dFS9czfpiSJER4NnnZNuw2rw8fHvpKQ
LCbQz2fLOgLRjXrDFMo4SL+yForwqsF59cLqBf/+OyuIRtKAkB+q1YHX7QYW44B2
VL9sxeanUmu7MzFySZHq1LtrkvF+KgL0um+IguLeHALyWNN90ogKEAAJ/Sz+UswL
YmWOOvunz1xDi9RAkFf/BOtBJB0nUokxo9Sv/qh/BKf3NuAZTAZwd0DoGBE/iX6r
u/zGnf7xNlNtTgN+GQ+XDkcpYWEfoq4xvzXGqRHLUgPaDyZdh180wOiIhJ9ilCF4
CWK2Tr28JKVj92e8tsdtoVHeqS8TDIBt9p2tS8yaih40kMM9Qx7PET/W0VZtuH8M
mbkYLQ2/qWpk+sr72mGQTr+DsXD9nV4TgZMMP2kSeqJzd25a8nZ0bSa6Ngm9DoL5
MQfsnQ4tdOCAe/nRJ9n1GFNXloD3SQVAHrtNyUTZviLw6Be+m+J/q/or2Cyjshz/
v76vVu3b4GEGBKtJWcPyxu6cFrYGm0GPDXPMfoyFsFAcyrrjJhomHejv/jzGvD3e
Xjwhf5LF59Oo5ZAwPGlBrnlv5sl80Rgzi2cExQ/jYihW2M6UKw0nfv7vihB+EE6l
gPmmptxzxTk3BvF/XjdlnlVsthEskijkOU/2qaq67g3u6ePOFL1PMTfOsWkCV2gW
1ggfhEX//fMMv/mowJa6DP/QeYBB09TOGl2J5uvnQLoNzQm4SXukVEXh4bRfWOi/
HJ3RbvHH5ntHu2qHSkhWcdQYJbDz0fmkiMCy/HrXv3i9aofnL3rfklPta7+tDzmJ
lSqHAuwDE0Ga9BB6OABfHCbkDcNw6XMAtsOdKsz5ciXsYH7ORIijtvRHzuOUlS+Y
IZssDEZNphvHdfIMxgdqTCL+8evFkSFceg3fpFQ1YSyZlsnWrLVWw9hqhiKxQVh4
B2niu+yJUyGDE1FMoUa8mh0fUBrWzXo9C9nL0SOgWjYU9PVjS1nNgYTouyMei3cY
rNMdSV/RXHZESg+MUKXBh0+mziPWyiSfTBRHdKtZA/1RmzBoYpdSRxYncm2mXJ22
`pragma protect end_protected
