// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tyzHs9hJMid4bOTTskOr9ZKj/owPpUkeKSYZo2nADLhjNYUPs0eVrBUziush0mWv
d1rYcd09CTCGlZUT7uZrKlfDB81sF3NsseImo4j5HsaVk/PrqJwXlcpfN6Y6sZn/
6TIJH9rYbCU7k3g538SRNGkuP0iYBkIk8xj91upKU08=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6384)
CfE4JmkIgqorugVP+U2oTHYcU5Yxpop6E7VcFqn2T7a8dD3EDii/IsSlOQOzIESx
TFpRM7LauiwdaAzE1keMs1s/P+ssX8rAbhjxRppk3Z+fsyyodiB1jl2ljfkk3YA+
JhPVclLObWDKw3L0q9mUBD2AitBYPn8Yfwf2E/r+s11cTIkkE9hxG1Wtt7t8RjfN
MgAd02b3VNc4tiBY8S6kedc4lOUlMgoKJb7FjbkVh7AMLQGJzIhqq9/vT06u9nL2
THeSddK3OHr16XjrRahJ79ZEm2OOzHqwpV8eo1qIM8vBeBZbFpyM80ZubgVtoTi8
tbPg+lM7gYV4I6wK4o3cU0oZJqMzY+QJetHcQ96vs4YHzK4nyyodEhcZ7cAgqBiB
4cG6MsTm8Kbv7gvdaehFHo41t19M5W9NV5ZiQ7mvFNHTwZGZ2brVah/JgYP8nxTJ
6pbneLeLmyufRodTOERkGlNcDxgbuCs/nCssrLvuRP/dgvJ7VbL4kFxdpVq8fvHk
ZcA+fKviA7OPO6vaaBfIko+T1OvcY8Jg5f5gWuAkczL7coMoII3BjVGIne+krHG9
qWJZMAbyd3oV+hlDtcaPwXpSVhsAnva7tko+leCn93WniXyBDFmtY9n9uo4QIhaF
YuELCGxr0Mrw5vNrhcmUJNY23CCg9/gEd/ef536oq6vFmpgSP6YrKTDFjLQjTdOI
mOYxrHAq0eTIXM/pSgq+30XsdBtAQS615JrRJb6Mw7vGJnoNN6NMzeVol+q/f9p/
Am/Skle2JxYyFwT4W334FKNieNMkoidwfHDHvlavTfkVv04bSR6vLrHLGWq0bl28
29HJU5rFE4RmeIwIDr8yoppsDGchnsHLsFNAdvYp/CTl6MzoHLx2D7/HXik2dzvM
CEOZMHBlf8RSlOiqQGQtmnYiG+DtcakCOLeseyahXUlAsA1EtN7qh93ciO/77iEJ
4MNybLBQJgN+xBtYvRKot7DxKC7HQ+IE9Wws+I0JLrka+wQK2tnkSs7Ucn7OnFSo
dziM1Y2oWCKWtYfFWLiS4T3IBcuSfLMwPTiDQ+NQm/je+QM6Zo/hbHUWJfpLTnEJ
5bgGCufzY/rLNSGQJ0Qno1Ns9KG2yWSIolMOUL0hA379957ahAiCl2MSTudPI3CL
KsRUDeK8bNTTbO7KSR1o6BjI8lbfxX7HKjgLscGQvdOs6aeHZNexAfLjZyu0pDVa
fvE199vxpKCnQtF2+ZiMKfvw3EQojKlEvUFgae37Z3fgDh6B4ZGrFkBi2rDzUWBD
OW22N+uK8NGn5BcQwGcg51GP48EMXcUxyXbHpnaqfJ37ivIN79nQkm9z8cNSTrqx
90WWK7SVkjv4VjVwCmrHEwv0b3m2ha7d/k0v+JHX78v9L/TZ45pLEBIITZqZ+d3g
XJ3Y0ya+eo1e+HkoqtSyQBmlkpF925tTGrJLC4qsBedE2CdMlG+5HMv5+KE6P/68
HPt9IUWg4GdEm3zt3W0gmktLZuU6pMU5FHKhDae6/0Y8tYKWUYGo1U6Dyxu8YqVM
df9sQBdqGQlJXMgMchZh1JQSODSMiAXewVo9tAMTy8cxqr0cdS1XGxwWvdbbjq8x
1UzkCbZrxabzo7PiftV7j36TaD46V0/yoGAMQkXKhZAoUJY4IuZ88eLwn985tWCo
e0rClS2OYCHKs13NPoFLwa6w0x+u2/G0TZ7+lohwszTQ0QmQLCQ5XZmFJS592XNi
PglP4gyWXOaQfkL5Zx03x+k6nGPAXm5m/cY10YzEy8sQn5uoqelWL0QjBARzA9ET
pys7IjUB/qw/+ozz4iJrTSh3AG67CKBcLW1M5JgykIF0vsqN4Jynz1or1/Cyk9Y5
dmgAWynbVxg+hxrzd8h7bYcCAcVdE5HyikyAFrJimojnTaK6/K4u8TWK1f/tnNf1
HoJ+KDn+8lTN8596Lasm+lXuz7uo428kguxBFjdsM3x60JozV1yC4DGdPw3mt4M5
4Mk0BenkWbcb0pRL6SO0DtBBtavAiv/Sl7NUlvyoAlwidblQj1oogqo8WY0kBcIN
BlYTfARmbtYvsTy6qjqoFRlyRiw4h8+eIkaQsnFbaqFelXWCNmW0TvYNO38vXpso
7LZCUSnAKy04kqoGQ0MQrqSwSORJxBRxNcmKawpS7JUKCw7C3UIUyyOwF/xMNYIa
P1xtpA2Ntlb8vtcVQKiZpHxx2j8JQjV22MONPOYozTgELlnbYlcVBLdJvEOXO5rW
Fy8GrG5EkF+KE0afhLiqnHztoM9IMCxPIPIg+Iz7stx0EjYsNzBUuAE9hh5f2uY4
+Sj9ZWXtEkgmT2+0Y0HhVaLi0UrqL8EvqCWsHGeK/GENcsUI0+rkR9Csgn7HTs4A
FWFZuA5rxE57Qn7hy+ljCtCfI7Xz9IkHBU0mOPpSuR10VZ/ugpG79EykSIz+acRF
A56ml129CW2O97Jx7oTMDQT718rX/wXN3iG4ZlBjy75Mzn/Ybuvw9paKXM9F4UWi
KHc8cX3RgEZEVpvQgkFfUUPXB71FgZyXJlrz4DxcCNriT6tieVEZlBAmTkz/mr9M
CQJM3tbHHKaskSDBwLSvA8WNZ3KLgvGO2cbdhEr0aTxLWBozUB7cHCvIghAUkBTx
ys5k4D10MDM2DzNbJpvUHHiuKr3HU78VqtnpSlubaV8TnOy0N+nf1qNBOKdvu3EH
D3/bV01RzqsPYK6A7twvqCTxj1Ipz9uVlbQn6c8RbPCquvEn+z3qdGsfxr/m5JRv
EZvPUk15ZoPCzuCsQSlnUDXGoGL9gJb9v24HE/YQMisjDQAXcqgnxgp7P6q0Bq3A
O7iN0rg6hm3dFpw4t4bVu32UWJWZJ7Qi8DjdPiWPOoNxSeVtW1jwhw6j4EZJlfQu
U+KZcAe5jxAmB1vMuOvILFp0VjXS3yXg44L5KjcWBVzeoKQIfRhq/O4AszOMrjxq
YIX/ziLNJ2HMs4OtpN9PEGnrdgwzVIEaf6uUg7v7LHxkfoOL6FqTaP1wN7vCDVqD
TQgW8ScAaQf8IsZv8JDIBa7vLdyRgr6rrGPcahOsUS0PUwIFdOlKlQE1//VJO/W1
gft/U81blDK8nGZSlVn6YBu47OB/+Ku3wxLUp/odqPWqkWQYgdgAY7VwiLENRy9A
dlFTgI1Hv6svitUWHGsCU+Bi1h/eHx+q6r5xzA5GR7u46HVoazQ7hvZtTrRNqux1
uQcrIHjDu6cKYwvXdaNEIEMtCL+Eugdf72d/068EhsSr4j1bak6VS6Zu+f4VKTm+
7IDDTVpQa9ayCfF3Cy/AYCeED1rA1dbb9xVLAVfK5zwuH3hXNhkXQn9QnezPFE9c
krT5nE3FRma+3e4UakVuh054ieaGPuwpFyuYVMW1ae028HjvNxRxziCkKHl3aLXS
VPayHLxAFHod7GA5I5ZyXC08hqppfFC+5cBOL3AHJipnGovW3szsv6sqkPcNX7NL
/Nd5zJFj6kiOFY+ZSTjk1sxYkLTY6UYSo9YopNF2QPAeSThMPU1DBWtFAEbdQ75e
eebKwxYK3cz7+SVxlrRYeWUt4fOgRxd54klHgqyFJvF6OSlxwM4xP97Z75LpMQuM
rftX8JjwljkhmfEs4q5rXbjfHMI/9DzKJY1WCnOyDYOYr0u2ZCdsaH+YKRgSW8bz
hwecPTnOX6LxYT2W6h6k2NbLrYVZk6MuaW6d1lBapTEBPk/c19Rx4t+zKSZSRRIq
o14xJ2VjBIZK9umlakysx8yQSMnNIkwZytWIir/2fmd4q2MIsurX7HgNIyVOhn7d
lkfJMhUOVyy/Nz7PJDv40KZUJf4eKq0JRpFlsfDyEAMKSy2DlSFb+Cocc0mJYEN2
MObjUWbx8HPE4VrBt7xGbGfv21I0HaeyDtXdBmp7xjOccLTi6KNKJe+M4PV44rjM
H11z9skWxAgM9ah1oDTfJONOCV9H8n/P8oWs8uomBoIzIpKOFgD88xjf/GDllkRt
xkwNrX/xBIC2Ut00/VGolyKYZu3OfPAEl7vBMRDpViVCgz/CEDJsbwY/yq+uSeyq
dE8N2EwaYwLcoWbkwEUIT7REc1XFN9dhn9Vnwg8M6F1d/Ptc7gnp82F8B+oCdTAx
jpHcHxzMV8SkaGeh6cSknXIlVj2MfweVhUPW4Cuxm84owABbEiiASepeU3ochQjL
Gp1DuiaU3C49mEU7Uxq1T0ykZ5whg35EbAXEuUCiOsU7cKhjyt5KgsJgx64eKvPh
EES2qAzjSafn7otomvEkKW9Ab2b1c1wg1OII0kLiBWYEKA2cHJkdDENJp888A7pG
LdPna4jnsHSL+pJro272Y4Bz0wg1LhMo16WRxKTYRhCk7TDnDDwGWBem7jbeKxY3
dC8o0mV2dM+SDfbmV8l4osrMZfK76ZbcVZPH64zWP5BG57nMjXAlJUfgrVQGWF60
WiAIOxM5ZVaE6FlLAgzj3uUVcZGOHNL4uNqjxS+1aDctBDyEkBL0eD2oYW1e/0KQ
TSMi3HfQeNkOtDVvkPSDJS5hTm7t3ZHPFOP4kmjGv5t+G72Ilh5PoZJNW/iss+Og
Sza2H7skNw/yi2tmukbuzy6kM/cZmI+vFdx1AgPK9uaQJ1yk4iVvljBazzGqk3BU
K85bkXyPt2DiXrpbve56X6sli5XlGy3F8jpgdYX3BeHgo0aG/T33VGrII3SbKTZB
MoZuT3zXMQhVwOjo631A55iNLCE1GHk1sUQNCSDHvmB+T2i244UtKe3+cmjnamfN
h0S1+RvJMUkG+kpNgp6opKBj1zWunW+NhHSOxpUON7tvPoFfTyMK005dvVjoFL23
8gDaf0GoqMNavYQnHxDSKA6j9aE5j684ZmMQ9Ew/+V3KyMmlJ7KT8B6pZTIjZcsn
LckHfWBewTdqn2+U5tsqkveH4vF6sh3UWCsQgewYuAdDHCnkZ/AKVXPpKIeK4NxO
68x8GTNvM6KF+6pRa6eMK9a5BTUQ0lC82jk9Y12/VS0IdbAW/Pry5NPHOGlnGMWB
OW/xWHMa/LRtW1gkQaXTqCAeJMbHMfuF4lYt9Ny7rSLglaj1P1oX6g9Dbrcw11Gi
wtyL7F8Q7nqEREzdhUsg8G2BN0I6pR7Gu/Jg0QsINUx1xpvsz4a1D3Eci/KDdMVq
r4YoxyQXRSEbf8PpqcqD/y4znz3aqg1AKVzOjvoKfjGBwtCOV3L5T687+Os7r4NR
AfA6OZ0KtAzsU/zLdp246d29WW9u3ZGO+Og/qXzUmm1k8MiPl8oTNwQ2dvXKf3ZF
LW5GE+Y085Ijbi+hn6OvX/nsON4mlFKGXgGI0Y0lS1gVOXeh7rIZH+qjpnrPaQtU
cYQi1bkOIPi6aOYDtS58VLllOi+NKEJMm5LnklDle7tNkTDDcHf0tDelaaB4YKM4
5EmjqIX3nF9KaVDxr3BzeJScBtZn5KuUi6J+t8X5xZpOFAt9JRyq6+vAiypBF0v+
yJ6EXdvU0AxonuPG5KvpWCjsOnYMWhpRvHy5QCImCsSR8YmxHLCNPoPGPqER7uwe
xkB83qYujzehhRjmMe8Zba88UY+9f5AYZKK+71pjfJMXNqGiY/bAeJCceoZ0MznB
NKUAMI87HG6i7qO4W8VL8an6baU5T6fW7SeqbPBT/QhBlLHRfOQpERer65IQNw6X
lZcZu8+Ez3mSQeu8IQr5zCQdf9N3QGNrN0vj/agbTZBH/eqz8SvL8+hlTJ1zbXJX
DYvAWED64mcxWxf/5PRQ70pA2pA05mYA2H/9OFlKq/jiieO0ks9rvIwyQqb31Oif
HIz4pttjVelE6qGCh10msKAd4mCntGTg/xNpzelYIA/nmxWSGum+2U9VbqKqsdlv
n7WGjVUoQY4dJDU3kxRDLFwDjMpirz+lWY5uTgsufwwsSQ/ZPRVQ1+SbtX/ApkOe
PcQ0uu/Bi8+1ShCSmVBc0ZYOgkXGU31Os1GXGeyMYYcqYzn3Mzfr9gLxaumP99gb
bz7v1FptU8u7MirHPHCca7EMopeV2F3YvC7mh0+7MrLaeO1zyIUwioD118Dh0ge8
siLJvudmJ9GcQAe7L5iNNMDg/q4zUVmCfbrnqBYXr0CKbnZuSoE4Ii9U/Nm9pDWs
ZMIsbqFuH4pNEni2ou1AuaoOIhL9eohymsCqdb85kMYMACJqn4VuK8geYSIpWjXP
zNYv9O1p3i1NjpcxZ0cFb1Fl5j19m/8ildkEQE+bsq3WOiXQ7y8AHfVmamMbgzU+
DERLskrOublq0zek7x1iXyCsBTv2B+4Z6CcNt3xIkE9LaUcQV3Tm7jKANSH/B5IH
TWRzQLMIu8X9gnNr5253Da8Q/Nn5VlOdcOtRgGhEuX9Qiw/AjLF7VXGJ/+yg7IdD
vGyRC8iVrjFYMMLjbcq5SDnHcHeVh0XCDYd6ewbIn0iby9PxvtWehUoKrS0DPKM4
P1Ck0m6PepzTVExnznJl9TQ2493DG0Il8c3ePOGa0x0cOjbTxE7QI1xKN0zSeAOG
oFr65BaCFjQkHStxi39NAGXbZCUwD4HgxEn9aINlTmHhZB6eACib3TwItjs+iOgi
Phd8elJQUJrSI0Mdfk+SuGsvLMvfK0Gjjq/EtFwpk7g5OPnTLFHwb6ka93OrlcTz
gnkw5oKKOdt1vHG0vHA/en1NgkV+4ZoVEUBqrHVeGitpUPTPc96aFHOR6sDDpMeE
pip7jQ6RGH2Gw26qGSBkeheEI5FMeXUlXPGbcs/1Qjmu9wlRRO2yAwjf7SMaIu3o
k9b7a+HwKM31eTtgoY/cbeMXYoIdT+6jinn0OaHAFI1KGis2ASRvu3P/NFtZWUFz
blbU+kYg4z6K+WMyBl0YddEeVEAxQNOVmZb3c6s59kG8Ky8T/3v2DVvGFESKqKj/
gz3djd1f5i4ilPhVJ0FnO2Te1CfdVOFA6IVnFPpWq0KgLCGbkpVu2ZS8k1HhdUh/
KQFBS4ZVDjBTFCBEHoyAZyrObYdin7fsnWjuS0YekYTvVNB3XYGqkfZHKwLSSZIR
upx5UBgtvDMAKv3gm3nuJVbrTy4nORNwJLb9vEEhIcwypVYoTUCcC8qDTh7Gra7u
dlovLabtqSpU5/doGhcfI+NwEmbXyAnjprSTPJjwhYS1TOoNfSdEwNZwb02I/6i4
bmGQ3rDFfQ/R7Hq/GfIsUAgRgp/Kz6JBTzx8Zvvs9x4FcDcV6HrvhYJYP6nJ8kem
eP//4dy9+bdx0FTGR876kCy1FNMzY3LcjtzutZPtjnIjzr00qOtGe0AxMld20QOI
JkUQlsGPf4EmPRyXeyQ53UYBJ0Zmmvlp7oY0gVKmc6S2Yo3NB6+0HfR5VxibhRRR
OwXQnqikfsk/HDsCQLsVxiZclIcelZLN9L5KQqnvwSTqqY1kGSZDRUBin11T01xf
odV7nZupTGC/HEDLHqhfGdVUv6dN1At9tYIrwdZVTDAfnSEEwopnuT4XErYZdJzh
ax6v0gETOs+rv5rt71HXz9xEtKMrXGeqL/ApDcm8UUleL/m7TSdJE3YcUE2Kv3gH
5/y03f+c0qFezJvJy+L9NYV7p1kPro+lI5RzDASpCm88JpCNd40wuZZy8bycxUzB
/4TgFsMdkFvrh81wmuwW3WtHcBdAwLBYeVemPlxfP3v9VfVEfVT6sAQ1CkoWANrr
JLQ5t4+GevMg224VJ1XH2PctO/sGTR6fiPnfQb7lzwmAzfcBb+SMYyYL07j33Sfi
ptAlJmoq3YN9zwszl4OSC/0kRYicnm2EMqUDcnqx8tLDTHOs/hB/Pw8vUITU7WSc
7h4T5aIu0MtsbPqzzEzqY/8599sCPYFKk6uyUjAkPWZQTKlffrTPwO3IJ6LNxBHr
kPwjvN3bmB/IVRQs/RWnQPSwKg7T0jwZBbBoTw8W+Ngn36c/dPcwAjMnCs7iXqQu
u9juEXmZu7CqrIZOlDc+0P7ILwVW0ZpqKgTNZd2zQ6r6XYsQWdbdzJiPC44r9HSH
LtsNXzNKUAmroFLcOXXcwagC9YNADKqc2KndUN8/gV0I1TRhcdYd+u6bOFGP+dX0
eh8AygBm0Q8iq1xVUyzNO4EtPJ0km9UW4UCFXoW+cADtmzeDMghnM3EJayPSftjc
5bveY+sEIDbKSqLJuO3DOirJMRCIpjV0rKVOynTKTRp0yNcW6B/hzy36Bu15eJ9/
CSceRCPwX2jspoMSO6m1LTEYP8jj/K4ItywGa6x52BI1xwl7UTQew0B75VEaDHEx
8FL3AQfM5nIAlol3i0hARgBDLm9gGcrxNisLfv2flyWn2Z468agntfIOykg0u9AT
fr7Tog59DBsajj95YH6wTdLm/wsFBsHnzdY2HWRWXCOq0HSonhL37jobQj2U/IHU
tKSQnaIWSPlc4UuuHuKpq4ndRUaM6OVyflyfxe1gs+7+/Fyh9DTJXDUTuNMpc80r
GvPN1ZCvRyW/TOselYkMkdGVU3Nf+8IvlPhRHJAw56Q6NYKerlq6+504KGCj9RKL
9lGhs3bEckFp0QBRWfmtJjV8+5CxS6lSIgM7tmT+yOB9xjw67AgqQx8bGDTUto9a
`pragma protect end_protected
