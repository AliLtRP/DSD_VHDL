// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k0HKWJtPB/utNb7oqJBf53ywTlN688BwSN2yOgoDk7kckX3sF1snjbX+hNLLkp+y
rO2aGXuVeG0kzglqueod65jo+0FplGGdSSLITOYtB6GlfjN8ZhwRwV/4xaGVdyIl
1DMZJuOnaq/YZNK9jV8Lc99WOUPurfnC+KMpQaERJ/Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32704)
o+IpXfwjC18OPTkYbjR0V/S3gdahQOGqgRezV6WmHyFMGkehXoRWCBVkimRTDrbD
jnfH2MG0czT5p4oY8Sw9p3P+Dlaq06gtOok+SCmtTn/DiP+IJx4JgoiKBA+Tb/Wx
CQrtPDx+5nBU+loK45QtmJzdLfmtNeMc0MTbdfbbJconKjZkWqhyN8QjmveOxdEa
UaUSMv1UMCPnPgCidHzQHvdAAYKQXDMq+miSVss06+NFirZN7tEtMVSyFEOxlBQy
ORNbB1wc8MXBjb/QEYJWiiy2gkyArhuz4gEPMw+wKpLOvjCVbSHiLVyaWv72tMha
0S28+XGD054aOF5MsW0qWm7FcPweKbwAWuRZtSn/ZbYYPqD4xzlPBLOgN6GuEpC8
l8ffYCFQivzRq5O4BBuvM/Q19sbu41szNPSpTrLIUQmgdKeZTi8MO4S2EDVFoSQ7
CrIoMN3/5nbp6+n/VGTkA3FGjlxhYqmRjfoQOGbD72gcYgsQg+q6gYbBwrQm5brO
7EgS3ZVtSWYRv/pJQAZLwVPn/JAfGOUPeoEq6fxLRfCzSlkpafPGJ0MEt3o81+k7
Qc6E9ctHGhlO/BH+zRTdbEtqtEk1UuZMOnauBp92JaMTSxA+Qo9JjL6ltrZVBYwr
8xuDUd7t3jRfchyezAOCF/jY2XTvH9WtlPnw0v/pCfxbpOpRrj9uoR2GFoQQ3Lkf
/ihjLGofZR48yoUa/5FSkUPGoOFaMa5fOAU2Exm0umPpWgcLfh6j/lGlkrDPsNNk
Wj6I5it5IlNNM5hxYF/DVex5TBYGs+xyOrQZ2sQfrk07EDrQL5eNusqfBTnLM9o6
P2dGIDzCooDwVnfo0E+85fWqhpLO2NIc4THuZySyyOJFfItZu2LqtttVMIb0I4c4
l/PP72NjOEbqY8VSSdYVYZ1gbnz3PF4O+clEjFAGM8HOIybTq05J62XqziT1shoW
AqyVk6cFNxY/ttWJ9J95Ko2FuXcst7ZH2zgmEg1mK9GU7I5MXcHo8h+7YZlC//lg
8hDFHBrtIChrWXYjQlpANSIMRud8YffTqqZa+8Xy1D9IzX+eVGJqJdBhveT5A0rQ
28R4NdCfiSIiaaP/5glCiSIXIMQUt7Ppg6EmuANX0fL9IuGplWLBe0kz2MTRljvX
SnYOlf1St0LlQSfXpgvtTLOspCa8qRCWB5a3qNXt3aqOqc1Lm615f6Z9kS0nHG6r
NMtFWPJjweC9APkMEVK0of9OGgremeB8RC/IfqsadxlVePy5QQKQ9xT4HHkODnsu
IfzgNuJapL02XiE6ijYXLSVtiOO322OqKivNVXyF/N0nrIVHrh0+/36pJ3htjNFS
NQSzCQAc75fmUIDzH4ANIOD4Lg5XQNgP/Gk3JD9VG35k196lx1J5M6UXtglDAwC8
bBJWt9wKfdIP6seSqL1DMdyR8B5uSNVmWJtDSsO8+mC5QmdUDTNUBXAPb0USdr6u
xVlRUs6HvL4otWf16+5pXEyjeWf63lB18BCXiQt3P6KMk+mSVakL+bcK+isN6lDJ
nXloV7VuxUei3xK+Cp86i1/mNbTUCEOqZ1REKksVwBVFvHDxAWd1KM/710xqEvI9
Q+EitX6kVA49AFfshv3m/8qkp6OiBHiGx4amNxRI/r/Q6M+rGj5uG5SspDLZmBRC
V6CQqMu0MNSxIUXoZteA6nNToqQRl42bpJuvKWT2J5wT+kCL7slJzEySn9ckao3I
Vev5xlJ6eVSZm2Vj0sh7yIbuVOzPWh+cXsvn5EaV4VqPA2W8ltwlofIBvoEd3LoM
IXqhqcmEY0siaOUaIrSaWt+2k2/70QqccFsqnnBdBknU5+NRwzKMThlQsr1sgRMb
i8WZ/uvyiPyD3DSEUIRZW4g+MyUUbdMxu32yAW50nuFvjqHl9Up0cg5mcVnSfDTh
4fiahpzBWt1KEl6tNU1WBi4etcGoQM/73GTzOdpbE96CHA14G8LEVz7APnZoXGor
4Xj8Dao4981H9bSrg/RVmhR6bUjCVccZ3ZjnjI2v2ZAdVRmmwhQRge0T+iD6FyqB
hCRNG1l3ZvaHijxPjNXC+s66vUVI39ruJKJnfoZP1IhtKRGAIOx9Zxyysd6S06hr
wlVi8afneO9Vn61OYYCj1bAVIaWuhvKmKpYhI1Pnah0VWyxpKDWtVkHaMNc2Aiqz
7eD2xjO5zPz0IpVBD7tGE3einok6Bhn0xe9pTMK0AcVOHq/zcKequ+9avzLQNY0C
eROW4xQVJOlf05KmRhw0uM72uBhyWTcxoHpCVWE5l6apUMurkgLZRQN7HK7hZmMd
n6tKguri5XnDsYcOn9RwmB3UfxY06tQ7iu+JvjIgZT0DKSDui4liEwiPbYswsrQ9
UmAxQ1C/897CzZBVSsj/mEN4FJ30rYb0P+bEBNpGr0TFJ2pAvkMkyeIcMFYUaJld
GgqbF2jaGjXWYm9zgH754wJ8T6DSrMIq+3tOYRE6jm7wVAEHB+NoXNAYPDbBBTH8
BYDMaFJzeEsPwMTDYPvm6ufTqaJLMKWw+iFvZyNVXv2dlhXriwagsmeiooDgepQV
F5HTgttwrJIK0EV6YOnJC80qLWn+v7aMckpyzV5tZrKHhOglHogAndwjI8qq7o6i
Endy+pyvIexTScL5rn229A4ay0MTCplRLs6ICvCls91HtXXrTIcotVkc3LvEzcXw
k2Haiz5fuuyyI6EHkZbfdlnq4c4gfI7qf4TJUHqkeFh7Fb94wQxjxEEK0PJ+1aG1
56gp5M1o2Lf00gT8Lgr3BlfycQ5J4EThsB+mttI8gW7Nr4JvT4SK4rpRfjB6XjDH
z/qZ1he/kq5jPJuk0SXtERBzuBRfIvaGD1MSioOK6zxqLUuygxZiB+8/snH7oroe
aI7lFo5eM0sjo2hJUu1C4vth9jDMv/UBgpMQYJF5H43yd+EnPHY5C59rvd/pItkA
2CTrJ2hKmthfCuaoZwTCZ0+Wlklsm0XofK8LKWABu0/2x5gNZj0azCZaHQqSByyo
8OvOCJTjEYEpMu4ybi6VGDLxoooKRA9p2KlnQNIPlav8oc0ss0yiKSxhu9eXrJ5R
H9l4iXPCMx/PU+sZ7zASiwAzg8xChUrXyInMTR2hVZu8TeN9MW+jrdU0GaE1/PuS
X6RUiAjoAghpaZWdhKPMTi1y5Xt4gzGznQN0YCFe8fhV9D57zIqBxzk7NhcrGK0T
8mkE8G4gRcs1tmrXhwiEpQEIo3gO+3q3lPRg5YOOG28RVbth5igxo2ljIdgaZSQk
AZy9Yh7KzbiUFbWQvCNazYpPReDeKsN411Ml748bRInLywrZJCnRYj1ed0jlhUmj
oZpyq1k9FBzzqBZR7y9IAuPpofkmPDnHm3AdaWqFOrc1bVa60PHjQm+67rpKoJh9
TNMUbytxC7iOTmypThpT4AcRDpada0qdEysyBDk6Ew0L+CCXN1uqG7rzYKgZQhCp
WUoc0NBPa1s/QKOnxAZG8RLE6+ae/FwwggOq8iwzvo5/pWER1feBBpC1ixDzi9Ji
Z/e02lPTURrtp7FIRY2Ug/zagi4kxswGJbhs9Js2SlV9miAVkTVVcdlNXVxNezZm
MCHpU7fe9zs7DJYJ2+tmgSC2XhSI/T/RekLjP3/ZHPVThRecP4d2HlntugLsrHJh
7Xw0iUEgOvTICMsg4xnCMWONQua5T+gH55kl99XaZe7uJkfDawlOzNDlkvYuu+dA
awwThkSwLiPAkQrKQy60VTxubK2PpBZidAyZ9exJpIfca7ITQsCm8T5jikncm9Ts
qaoh/K8A+E6wMkoKzsaNweuMt27Z1tV/P6F/7Rt99AsKc5mLlW8JPCTR4vLfPgz3
sHXY62CjmLAuv3CZhSEymhqBVyCNCW23tsICepWKT3s020//qRk0GpBxiRBaAevq
YXBZ71/h5lPei0XIN0PS0IWLiyiBtheEifwvfASV0DNaIJ5c93oJjb+v9U5qydfn
rfhz9QNwG/7FQNa8mGu1sP27cj39AmEP755bdlhqlvETHihsenQYAhso8SOsbRev
yyTaWZuG6mw6Sigy9i2Gt/NIet89ZBDeY2vqZE3a+x74D2DcU/oFycKAIexV8Bmz
YkBF90t3HUp4bzzPiT/cmErqth+ywcPcj+OSR6ew/AiDriqeDXl4Ik9UFCAjz5HD
1xK2PuoJTfp2QtXpzVULSoe/doVL5Vkl3Qoglc4ZpbFQ4rch9z5BxZ5HuHjjshVd
xdnP8JHkQLLJYvNVYhx5AFazrvruO14S8Go4hNllD/75mNReoChvcMe+LcCIpAUz
KLKBPRAXErS76Pn9jARuT0fg0iD64DJWPNypkwlVwAe6mvodaX65ukMZmZBVVh+o
FvQefHYaFrgYS9rp29mjeO3KmwoC3kcX5N+dOxzcnLRQynfqzlAAhpPBdc4iUIEt
mpEaDQSRZruYnX3rTRvjBW3kdcKOTjTEzAZnjJk6fxlaEKVvkz0142onelqV+wJj
MZSCId1vC03xDroxh8euCa3wJy8Z6rmPjbAwtKNXuomIp20uDGAsiQ4z5Rm/9oTc
MrjhvXvFc95CTRLG9KZoyYpIGZjBkTTGt+JQjmOeAlCo1uY9pmrIiDdg5Vtb5/BA
PUysgylJYEOg65HsHLMRkBXYt5d9uoQIPICqVGdMTfdc6TSaCawW+H3Yv0304YBr
NBHhi9UAhC1Pjh7EM53ZpMF9QBIC1vm4cDybqrMNdc7HSVw+ClY8S0PxDZwUzrDj
2fUnb7WYcTZgAnGdyG4niYpLcYroc8iLP84vFL3Do3EuPcFyQsfYvCjAoKF04X/+
5CEbFn8xQPnKQlCMTb2JzrEieEVJUbgqLC9lheHuydpmN5dv7a3PNot19uSeHJH+
RjUCzTupZsQVKUU6aZFBBjf+CY0vSL3n0ObdPES0GjgN6OBfyxobWJHc9r/PS62b
504mfaOLH+8Uui6EdOKoizNo850LMm4R6MIaSp5DehS9x0cwyKMi8ULL5z8e+/fD
SyQYjF0ZXM+xCc4YqW1baejzqLFeXKrp9RQ07Oqwf2bItOapM5tZINWn8IDDDCBM
0nY7gFt7usRJi8ix2pwm0kF8PZmZ4iEell/wUEE7xRI0D1EgKS9OYpfFs9sNuzH2
z8i+tqXr/p6Q8EGXFHGZbEQGu+UeMzBciRkCV8AhcDmlENpZUGjx3JwHReOoW6Dp
e0lLgKvbg9WsXAD/CjclipQBU0xRTHoAvBCSoGcu2FygXwOPV6ZACc7EtcJzX0/o
fHXYi5QMYTZ8XgYR700JxvfAi51bUEgzVvLIp8yblNZL4VW2tjvA3DHBTxeOROlw
G5Hxb/Bv8JfCqrW88s0MvZsuRLx9RuDgJ7vop3SepXhxRbUqR2t9rXsXWhi0bjR9
9ZGRtsSlnZm+zhWTcAoHeT/DFJZOMnJdTHXuMOWtOGJKdXgMp3BuN4URSHSJ9Ctw
x1JCv9O9ehBzkjUEc/ZtXxuE5u64GGSo7KT7LiumEndLJ8P+2CwBvBJy74ClDBt4
uHyGWxfQWKa0VqRc36ahtUf84WqUg7hb+sx2bkCKH+jNio65U1GnTayhKsXtTqhN
hJtjeIumbSNRU0C8d0GFwlpLMxQo+I+YGhOK1fo9C+WIRQFViqWv0SdCRN12IlXW
gPGgSM9gv9CqReEpxID0EFngi1GcSUzVQ6+xW4cErJbB0hdA24W5GO5dGI2LwCXQ
ShVnSIjwa7+ogFUyPL30R84pMgN4iYpFjbJ6lsefnFT9K6sJkAbU6YoUEjOxMr8c
//+MnCYd27jWUzwPb710Jz9AVfV/zBlQsvmwN8yqB4E2121xB4vObYHESi1j/w39
P7IAEnWGmT/zhlBCLSsA/4bn4q4DS7wgY8eIcvoirO8SGDW817mz3HJzdxCflOHs
EQ/9WCzUtw3solccVq0NQDjzZVOdu00PylXQcVX2QDJiY4mRX8HZJfmJA2PoQGkv
oQs5lvNs/lBV55DSGX8qIWPKTm/6FbN2f5asEyNeKbrydcGZ6QuLSR/p3caUI64i
OyuKmsKkBq9dzvCh8rS9FNYgTc0mmQSEEUGQVfK5Ha+BsBe8Pr+gfHEU8/QzsEG4
8x0XSubSkDo87e9lWmgi4SOIL8653U018MpGN+tpRmoTjxz92Kj/sNFpvHka4lmm
SfYse602KZlfXdsTHaTpoG9MbReBWeaSC21VX+QApeTf6fbTHXwmXbixb4B7d0oZ
QioY0YgzxNx3+zCaSlPfbx+tg2rq9UydOPIqWgBr7pZfAqNWfbqsbdYeH5QN3Zi0
Biy1Dsu4WqkDwazKqiqkGLDLW5hxC2EvnDih+Uo4Yk6RG5fmbGB4PlfjYbUJ6nMM
I6NIq/KgK0K0w6+fo1n/kWjuL71BWjmOv2Vs7yFmaVyfWssKowluc7jDbw+pI4Uj
3dn3QeeLkp3O436Mgj4iHQyQ+/27YrUJH+lWfN2W/L5rBuhbxPbVs/dATI2i8wzW
Xc+d3q+aw/4eTqiiW8WyzAqespOMNV29atVuD0JKiDvOcMR90XGkcW9iW8sHqXkT
Mw31wErCGTNG+uhsemeBhHW7jkTDCsrqtdoWAnl4yernAtfKpQIylS3h33/4qT52
19+jo0+ThLEXW+L6y5JuVD91+cP7Pv5IRlU6NMdv4nh0drUUYQ6AI+45qKSetymu
jkGE1T3p9GZx/osJn2O9vvF9Us5gyyZ9NEmkmLcyHjlA38kB1DjfCH/7ybHloGkX
on+rdiWGdAJzVGjwC+zy88PzpGzvZQhpswBbvv9tI/WFY2KSgNkKh2b4BEd0010j
VhXEyvylyMMzeVOI7BebE08B9a57MN+XRQZlp8U+aNyUzWi0/9elXjMWJzccgPEJ
oFxN0JTt7YNb4fs66qPKs7iNzVa75KHurScGKqqT24JjIepITLFyCpeGocTKQDWF
0zpOUxnOd+aAB1FMu/YMd4qYGOBpm5lpLx8h7CZGvlKjY8TW09toQ2JQcRhZEKZ7
cpZV1ybV/mab7E0oQDxcV7JoxitC+B6ydE6o9CbHLXNVH/kN5t6ID8cP2NHW3v14
zPNI7hy9Y5Hmlt+ahsDIiWfP8OKuiJ7SMD4CojYww65VI2bkMfCwnyQoHzetUoow
JpU8jwBkEFC5yZT3jrmGl2XeHSu8iUg4IS7fXIJQASsLi5C7yTEWyPQLnjImC8ru
IkvDCWsCdx5LR+91ETJr0mRIWTM+3zisubkTmJCLFki7y8Ceer11C6sdVexgKxns
B/PK/0AKWa3MP5is15AN/G4OeLf7zEzd6mk4cNovIbaaUmMzacz5fp2dMA0G+6FU
4ZXchCOmNyebIlOrgB+/2m3Jfce6BBK/98gQKb82IiBZSEt78IAwpJJsvTdMbCYv
NFx3EUBsXev9J4C2cefiBAIxESgLxEfPrCVnYl4SFGd6uerVuWrdCEKXM1Uu9zGE
kyVTy9WKSbaD6+EoCI78t8tKBYOjLn34Kka76pQhLG+XaNBQt/adPMSlArAMNp6m
T8iCZIYb7joNe6bYnIodMskPScH2VRI4MwkuI9I7/zULhsj9Wdj8zGleuOGUFGZw
I936v5QHk2zGjpZHtH5tlH4HJ8QVCXctTWYbXAnV7Yw9eHE2mFCOdg5rcP/fJrk9
3p8Z4b0opLPlAQCV04LgtsF1SpTvwpevqQnOAhz1YABhTyfSrJ4QIGHVoaK4qvDh
pmOtap+GHt9xnPuV2FVanXeYnPBwbmLs5qvRjUUxQg7q2PlKtpceNIWI/BfSJ2kU
yaDiT7nBUEoYnY5jWGCrMR5uDQmO4WRD/QDy8hdDJF5nXx8b3JRpQnMVKmtFmcL5
BgZNwLjEbQ8yCYsrNeqyI2kGqnse8dd2HirusUaOvsNSsiz8cQKGAzQeQW6LXVrO
Zy4WUsLhB/k8x7UnlBOFwauV0P8fj5RRACXhiTImTkKK1sH1kbhr/RwWj9uifame
Tr29UqM5gQHnJ3gTrnzuliYQ4Vnge66wIo2LEITlVXoZew6ycF043LuLcnVNBLMp
tABm2FAPakONLkLhL5pzG2BTN+g+TN6b2ZDWhQkCLaoEmVtsKtx/D6UBTGdUiz9i
jHEK4qt1q8WwEbajx23/1WV/mojK8rplREdrXYJRChuX8IDkSgBQSBfSkPbd5JQ/
YthgaZsYolmuvtfgp8Y83qLAmv4D1bN2zrwpzcb3Akid5FfbkLEmk9IKL2Vra4xh
mFgHWp0oSKc8Z2P0299hLRfk4dSNAMA05ntb00Ss76Q9Nl4ZSnBog/VxLO3KdMYG
wgrT8QJMdqu/i2VQD+l4nNrNEwpP8+ZseIlN4NYOjpNThbtRZKTeICoLdBtLvmUL
p+J/0HF5Hm8uxFwFQQfzEH+HxSeK1xn5jGY0/GCDU5G9O5Eei+opOzvUpGCZk7qC
PIgESBJRh3CrAwvlV7cSwH3vN3mTJ3BWfqHzW+P5xsEP/VsJyPg/MWzZex6TnZdd
oJT9+A1quP7dRT90dmtlnwekwliMm0sS7r095Xq4Q7QBV2Tth/7iWfz5wXCdWyUI
sZ+icby9LgEIvPh1eCM1Z8ESmXeGo3eDd8MU3AOldPEjQE7TOVgnEfX+psu5vE9V
nBtXtdXil6iwUcloMo+nLvc/zoG3jOAK1fk2/7tHDrb7ePbmXIaZpzMRwiaIPBzN
/uoy2F9CDgjxvCNyu+0J+2j8QUvS0sFSNE2M81AiRmpdx4gU+f9JK1bM5F+jI77e
9TN7mlpMjiUHeDSm8iYUM8fXoGdjix3qhe5KhiJVa0+gFRGFHvG4DDduIveF8+Kr
fIAC7PV88qy2EpErEyjsSuyh2Q0WdhIrS0Ej/5rsBfUpjFVumUIDGyrADgQdOjY1
HwRua77QUlCgbX4+p/9dtNVN1Okjz6GSxBiF/guCIQGYiOQQ2d4LAgnmBbLaItk4
fwvLO0YNPyd7hW2N4MvWXtaKouNdZ79ueUBmuGXLrXqIDYsEPN9xCKHLultK2+uj
WPrCNUQVwiEv63NTlURymT6YHlCQuV+hWLB3HUxGXBw0+nkJUhQBi7LAXwX7Evw3
qSQKXVqjPnqZLYHOyM4acm4+2yiDMnjd8wIGdEG7ibz4WwGPKoGxbeV7AhEhO6jR
PNn+wMWH9D860RUftcyb7FPSEVzHbye4ddk8QoVhsPvT8ecpBEteThQRlAG3CzlB
1KW7sdHTlDQPJ3nesrMS8W644VrqlZ6RD72zT7i5CUIM3NxapclqCcECdZRFpI1C
Uwqam4FfiqYu85yMV1z35K2/ZpCBG2fSUgTm39Gw5bCl0CeAXTKXNrZNQzDvLEHo
TfS51rcv566VWFmJLwJ9q+x3PQDfuTJe8noAu1DUkLuhcxnivOe/44ugqlwxWAXy
WXVjPMDBwCoFZdSSqrvZPep6nIkqRLhdvqchZx8YI4J207pgXGIk2/1xrc/C4dI6
RQXhbSpNAVye4CvaOtiQQqiohZpeScEtlEeNhvo9mzpwjCFZit3hmjdaorgy6zuA
dE2k/B9xlk3HYvlYsdo+TRzriXWVjmbUyPTq4ZRXyyKo1Xlcc4pnVY8zaL+h2kqK
xS0X9d6yM3z+VOyIlJq+qvzEFDQLvjCO/yGksmA6qHM8vRhHVmfCvl1nE8RpxVXh
z/zHWA5Yzch5Wy7QSbNbFEsgtTW9Ewpjk9bHbr9+41v7F4gD8BSAYVZ1X9Jd3ziL
/695frqWORoyFfY6c9FAR+QHVKr13yr2atjoSRXA6VXhozHDoaBEbb6QwEjgkl/r
GhbEkmXROs/D1R3aKpTH55KW4nsf41ltcgINnr6/sBCcl24sY509oYw+8esZmzLj
RoQ7LDa0XCKI7ervBmQoLlYEuKi+aUujPD3Y+c5LuHoIG2twpe34s7KSpwCnYOYs
EuOIo2Pn9q5Mahu21qlhcTtBCVeYCLK+ql8ogWu66LY0rkqNXWVK5IBvaZtjVVbe
2sr8BM/H6j10NoWomQdH6EWWDNzeXlQf1tdRbeyb0bSMt9IQtC6u6J8VXI8Ut3hl
1kEnPd0JJ+iS8Q8UNyqeiaClU6yb0EkQp7Yhj2DOWpBJMMFq/uo1fyj+WrBpxoLj
3XA9rnfVBPHViQuuHIgoak7uRNURiE3+vgDA7fb7H9VzsPfnzjdAutejtTR0wW1x
i4/aBiDhPyJwCGt86h1ukwMuERzEnpJjdzEd5z9Kkvjk0rVuTe9+c7uqNQU+BsNT
SlpqKUjtOFuMiYUr2yrR1cUk7It3kSiFDuLfWrcZoe7k22ZxWHfq6d0bhdfocUWm
k6uByya2krOKYaviq9BvxPlfgmFZIipYr5ZpbG+lTZpQ+6HviH5W2Q0mx1F1tJ3r
RBQ+L+TAyMqWoP+dEny4L02WGtkX6RrrgN/u8Qqli3RZxUBlaVi/+pRQ8kln88KO
ncLJA8wlMyF6uH+NS9exIyQ5Ru76Qk1uCN8KAtEjO1RRzla3zU72VVeEiDEto9Bv
VuwbhPhVkquJRT4gAyBs0RgNuaAxfKi6dLJL43/mAn/HrViAp0+uRjJnBEyY8F0O
TsWCTfvxtVUQsNlOlCHTZFp2PECODoDBMpYLkBE2ILu8mlthZ+dSy9jdT0pjQLaT
YffQVhvHYdA9rJm9sCjEvbQoBEVPqIQxSjn0eBwD/G6RgpsBpG/zUYPGiqFeznxa
KtGNrp8RG28hdMDfV82QpJ9zqBpgG8GMTEsRI+tjmIhLkrJGs5ZwpEuxQbWaS+Zw
qtXaaIU5/3hjAadj0cRE5TC3PoMywXvgDiWryG6AyaK2/1WN3R8Qn+q8Q/6wQzxf
3+pu4lRjJXyNP9M8PLVi8kkOKrixAlznSSjMIUYK2vgsB1s3FobJqc+E/mXm48bW
xWB2ITO/wgAerSjx/f+ajqN/deCNX1QG85FRjz1ng3ne7GfMwfiNFvyLhaMuOp1L
u9Sxf3j0bz3UDlh1xPv9duFSlBUEqBfIYr3qmG58u+y484pa1eUySnFMYrnrm7Hz
pgD6j4PGgxcP16YCmr7pZPkH7e92nMgu/3SHqnn1GgjdYVocHs1rNGBF5zsTTxhB
Dl3wbsJtEdGtAPBxXYz55msYszoL/dFnXhOwQ6J85yNd6DjsKS3XTaT1Fl0Enyv9
pthGmlF/q72KQ3Pba1n0mYBvLOIpdASoSjQUfflgaGi9hwVOG5j+e9b4Vx0wzQRP
FMfJJS62BbyC5finMSX+Bg2BSz8FF6TOqaK/rule7nblVWjOnXAPXRBmMf+supWT
C2MsI6v2IKkfnw36RF9s5ucaB+XHBOjnwqvTzCaLIev70+cZs9vlR941NHo4xd8/
n2RErWcwoQYodfg7HIcBRWNS0MazxLJNdoocRxaHMnLgLQ+Mi1qvKYj/rp56suKl
hrmjcRKM3kjLisR8sEcF8B/9Az0X+0xrpCEbtGiyp+VZaY0gCwouO0zcjC+fm7MS
YWnCVSvogHPiHWlGmt1+1uWJcvGGOm81UYE3qdKJ9VhZ5LriCeJXvV5qoNvy8PI7
cwfxSx81ZOkDhc6rwUDA8BrnNCw2pEEbJvv5gGX/KqMd+rvgX3QH7Y0M+p73yX33
2SB7pfNt2+WveRex0EwHhIM6R9TgSchNl2UbBPPrT3bolkY9RqvXcFqi/Wg2EAbd
PQZBLrcx2wG2gfFCte4c0CQH6UtN6C0W/5dEL+314ALl+QZUu5cXMqxmDwP8uUim
fZ27si6eemJURGHGAFeRsK5gIguiSuavlrw/EQUD9ERxzb/z4v1aEE7UNADp5r2B
F8DAZcK8XgqcZskHBj0noCAGteI7YRMOTuTzIu3acQ5zxJnk9OSN2e85DZmQEP1P
fXYylJBFVtF4OCoo/7AhVLBZFTwcapctDhN/Ta+iCyV9+w4cybPdO9qWO4tNEglW
ouS+fVlbqp+3sD+eB+tD11BDpJEPi7dupdb6tThNnA3t0bQ7kUuidhqvPXPQbI2Y
ewSQHvUEFk4g8bBBha/UE7yOhM8PR3nUaf8NdwO80E3xHFF6W6hacLXcR/mKUodv
3ufapRolKGRoJKVZVWYpV0TfuW48RMPb/T2wvw6G9D7hVl2auFM8igahRN2x6KJL
wOdEt9GVCgychFFN7Zk1xgzb6lkGyiodHiwHsj5OnW6VowbPte6L3EEpFeLsJAvP
a7b18E46i9VvFyAD2cPAKxhCO9oXtwo4RoBvgWtoPoWeJ5daPoCmMDd3Ot3xh5ux
P3BB4fLAeXlXLm4U3dHKsVZfh16vrwh9tOig1DKAmYY7BQoEcQCihc0uo0es1mRH
vCbetdZZkmyhyazh6NsG7nlfZdp/hcl03sCN1iXiOGhBRI1wk1YEDzwderq6iRNO
B/u/4u5/VtVk2NN9fuG+wRaov95m1YOb3r4P9vFXb80K91F+UWeM+3w2JK+1/+VN
l0QRFZBwaDAq7pz2mFo38OCnzCUV9SzRFKZaDa2l+kBH/Umz0MSy7B9z2wBtGseV
l6H4qMsNLMUPvKKbOtkZdy0VN5f9H+Z1NhApFGBhjYVS+AkiemVivUwSg6vgk8R1
lyzwtq03KKInKm4vd8gOvemv7DUqgG09swcYHbues7zDdPih2pkjirDCz2mgnkDr
DvKiR+eQrQRGzWbb8CFpJhrbyJFEdVcKpWCY3WHDSpQBOjWu4gzUe1j0SLFpdiD7
dNDH8oEesNmmnY6uq0dhgPs96KuXbaLXwnTOBckKYPH3WQHF7NJFkOVWSKYwO9Sk
6zA4iCBvAbWn4ry8cc95XJncYWr5vaJt+vVROnb/ZzABYhUz/kmQX3+fga1mBCOe
uioTZCAjQJxS00qfoZSJ10gP7wkpofuBSfQ3Yrvcawz0WlMl8xFnT6KsbQGGapUa
SvdYYZeic0P6zRSP3B+6P1a+0nBr6AJmsyZJnQFBxRkXh4u2iBSTQsFw7lo9SLC3
VOOOaeIkt78Z0mBXk2MvObRw3qnXa5o3u3Oe/y6lsX6rSTRW4s4HKXrFL9VrP+Lj
qgDNkKMBnY9EmGR5I62zhm8lSJpp56LEl5NtB2tWCeFJFOzLcDa2iq7xT6aewGld
15DbwzF5GqvSRtEkkuSux0ybbjPl6n4vS5nSrABrDgCYJXIF796QVtcXtY3mVWt2
CIDfTskIxbb8GjJdqZhiqaQFDqchQuHVd65JaHCJdUVo1GHWG9+51CI3IjhjZ4Dk
RIi/ObWf5tur3OSFUrBwDREQvNq02oTJgLflYHbfU/bpGvp5NVOu4QUTGhuR/kh5
pYzYumn7SO78UZM+Q2iSVW56O8xm9Uq/BC/7KuGmaDY1LtB/26xkFwcCNTcySnyL
vwHnnK5xVrmqTQOkzVVpghf7IbWmG//lwWtmbUIHs+9klIcvxfiMd4LnV5kQAo/g
jrsrnqz2aKuEae1+0mp0gqdoD1pd67Eu+7vNPFQiepeANpk3fnojVFgHrnVYF8iJ
n2eVyQBZEbUalrosYVyfOazir71xwbp3AvulCAoFMGJJ09AMr+/UfX/eo5VsaS5S
+/zUzq5yA76EaDW/dwtNWZFOsHtLVJH/aD2XodigyBshps+8DqiDfytrHX0/Fdwz
7AKSsymj4NGOvT2QKdgXRV/hkFxmc/g6a3ruATtm3/sDGPsXXZauekgWTOP0BOPt
0AIqr9vGH7qxITSbWQhjqVZOwVmantSL+Z1OjRm2HW67xQHymVO1rSpyQUoyBLIC
4nLd/1CDV0ZRRz9D4LnuvZnx56SN0fmGQBDodOtsOKLd4ZWGyvKbOlUoqioVH63j
lD2XC9orWw1tHMrteXqQ+aIsPiGOsj6SuKGhsFc3hV+uvL/XoUtvHDs/q6a6CHra
UeKY0fa8r+Ya3dhx1cEudlbLb8VFTKB42UJF0YhGlaYrZxoT4dqFIsOASkieRq5f
IYCPdxZpdMez6pYJKm4l9tqcrSlbgVKnWnjeSiFUEiW+tZeMs2UQUfbcWaN5bGwL
yCPDUU5B8afW09C9Q6WvO8V5F6+a2msCzrciMSvujRyf5MEt2Kw/mSKpX7rmIin1
sqAbPsxXuhdL14BE2TVrljVWSfk0aiSD1pdI6K3BuN8coNVcsVNDNyHWzWtoHy/U
jEVJqc/47Kr34MZsrfPgUrN+sXSMqJ8WoJ4fKpa6GMlkLabDjvizOZoePFyULEfI
xMrkp4blhPRYcLp2qr/Nkl+gb+M1bZGUgQsj/jZNKc4pAlbJxyGwKwRknLAhFUxB
Q5tQGVKITG//cxAyeUIBnacfgfu+6hQZ57W+VkpFOggcxqzxH+yDjj5YmTeqEA1y
I0F9N/ov4P1ayQY+G2uDNvk4FB6ErxSvhu41fSxyiE6kLW1gB6hKgqlxdGHJn/6f
ivCXmHQSRGrgf1QyLqDhw8szb0xRe8jaOzGIjyWyAmk4aoN5XDn9rAfnDRRIhWRq
0nTpiG1uPW0CBrjF1kE3trjn5oepaQxx+YpMhubZmw4BV//0ux9+eHTbZU2FWFH/
ZeOvlXcWWTxSWsP17wHi9TUyS3yA0DdpgrqMHufUQv2E8YbT9E0rBSvNkdB10ijb
PkjMosLtzOmM84XAomBBBDe6zjFbZiSjsQ8hjSqyfa+D5rZd1lfug6i2gmK98gY0
1zKa6pyXpTLiU0dWqc8bT0bFer1VKqFtueHalpXPAWq6WK5bpSz17bidIBJExzkM
CeO7yFwAzon3YdALM5LEi/hqLzL3V6/ebZNw7tjwP/u78RA6Z3kNi/d+67Udl4co
v1/aa82zt5gfEnfr55NTRBVnJi9Ct1kzFJMn/Mq1EIH/OK99jy5u1BJXDjPNj+Ag
W1+t/v6yso3QoA1agg0tvf4AVPBHdofrt2LRlvFQtVFZDQD+ErBEGh16ZCiHP7HZ
6eyLD7nut2zkIXgPw0xPuVrRvVs0dGaP2PC0bcNyOcHB9MveoIi/HADHpIaEyGAk
NtXsqT8iBDbjak3AWOtZpUJN4y1mimb2omU80EjOyH9Xnce5xWCg83GIYj3MiowD
m2/2J4hikVDGiNa7z8dDcWOksf95ZgcYyy5ViSIbwmdRWCd7TCVrQH2xf7H5qRR6
KhpGncxP3dSgpIw7xXdCJETRocgLh4Lp3eQ8rWlsp/o1vVPA/O3bdqTP6eW9XG64
5c+6LyJlssO0GfGnIrCumEMtjE88gOZfhwIxtJBOn/jsEqrFhbK1OIfgYSi23nmY
TOkxX1GdMLA7Qz85OYbkJYCi4T41MLg2AC1xMTgm2t50aEPBfWyxmSDQIgTegsc3
SgMMiphIjZQ3QvoEgBRAFycHWNBnf48dx5UBp/n8S/qpSFcm/k86V/RORtZnPHUw
2j88x21ILu4APxmUHfUiy+FYk8rwZgoRSHhNq3HBmOo/fM+J+sOtdz0q4YfymFJr
WP9ym5P3c+IwxlDEhRnLOK4lqmXCVV9naCz3eZ3fZh9p+yyUoajZTCty+lecZdm+
D4v9ATORmNTh7pDgAF/qrrfYAGGG7MCb1pLDK7/ngjGSUia+jdASStRwoOyjqtys
xDttMU/f9rztbBzqFefbs5PLBdvZG6SbgG+gx+wqubNEOSQaO87aHCfcslb4toZ+
3eNvAvzbUvcU1OALMp9426mLpe4jLObGd+P3jjHYdOaXAukJ+XT+K+qTfCJxJtma
vjLUZGF+ITidl0tYfXeVLnnPAnwXRm2DEwaljY3r8o/iGxA15e2BHHBD3/NykV/g
k29RWZ2NyKc7OX1FnKEeJ6c7+I5+t90M+i69Wu5yMC4lXrP+SJDJgglexOwQmcQC
QVYCsRCsuTJ6gpKYeHy+7KMh9i7LFuxPtsTpIlW1U1hfIGe5Y7AJHmtd3yD67l8P
31OLRfJKBGbQTwFFMIQCho7oXTCAMZjdtEGR2MiJkA/zCOdyQ2X3n9CstZ+4ms5Q
kaDrCl3+WkNBJlxyiUSOl49iRSoZQUgwsp7J1negaToSGNQAl39s92OZQespdq6c
46nr0jfad+JD+wHVclsKBebikpleoKKAe7C3y3uDxOUBwIerjCjec2XV61sIZ1We
4jsphwsc0zE73059GKOWrj7SJnZpp+tVG8wqOMtxIBn/4ddBXGkNTyDHiI2HSYD6
MvblI7Ji/k/amSLHIYUNUssxY9ELpbiFaZCtfQa0/ZYy3gOOdvGz3ekT0akXFk2S
vInOCI1CMgC/bz3GF5Y0RNUbY03cPxMSzblREpXMoTEoQor5GH9EKr4c7Sc4dyvX
wt4tbbEUdrfxCo+Y2YzrUgTxDzDjnr8GIzXnAecVP9ZSBKL/wmVDASgfIzaNEVi3
ZtvTsTlUiC3SuLjpbsG88+GqXz+37iTiwA7wZ7W0S6Rw1mWl3yTysIlRaxI3fW/N
yHi0NwmCYf5vhYgSnSDhjzj+0c658ouNpvvRpcs+PFgbEKiz1M+1D9YpazYZZijK
NvjTo35Xd+aqI/+pSKgahMsEQqP2Mv1WVNWz6IMKYM3ns+p1pbK8IF5OjQqjzpGz
b02w2qeftUxhWiGXlTq+Oc1z3CyFyDb78B14/fjE3UEwmVvHe59XfsBDrX+YMWsS
JgTIPgdZGJ3QrmeVD3g1jHtqNGXiFOByfgGfi+2Z+/soGfonjchb080ddVPDeyd7
Elum+qKsr1/jYs5/BfZufJC/Be1hv1fga6jKQHSHLG1PyfFNVC6Tti3hbPO/Fr4p
4etHPK+YFQO+t1534NagUJxDE9RuWk0qRPdFx7DysuCZ5tJQ/x3GAFA/yPvmRfM5
1Go+o6wAFz4GKczs17jfDmwmhtW4bkTZXsNP/8+nEubLDsm+jj8H6fgHTarnqPA7
p7iIr5jgBrRwXylfslX0zXO4z1nVXBtZ9h8k8t8loGjHxcU3aMv1zVyr2gXjzgis
qRzSynQu+E8RCeYBrkZzc9OUtts7UE6gtJn61CkboZadGSrhAKIKOBN8i4B0Sqiw
ObEwT5CRhl9QSbr3wSNGm8a7Zpgn4BeSzcxX5yZHW0+v6INiV0vz8AeJydx5AE6R
Asg+muFZauuKLNTWbf4FiEnOAV5tdgoOG8KDpMf6htREQW8wpa4hde2sTEx6TIay
IedFv7eejYgiN4k9H6HoiVa3MVNIaW/EWa0sfSz++gBvRWAzyckeXwBwnNmsV7Ae
jh+Heve9ixi+rof6cQ8lmzj3+QHOE5xeyTy6VNt1lT7+6PQeF/NkKuGpRj0G2ST7
YplsMeR8879xXcoJIa0sRABa8DPMBOUI6UoUCWyYyCjeD3+dYIlQV1CDbLVt0QFx
YUZDj1TlfbWx6h0Zj/PUIEt0yRT0h+/Or3HRao09nUQXS96Y3gx97OeAI5rMUJtD
A3blcxKOGtnYi1+ZQse0yMvTBZ0hqTavXIQlZvDqUcrDjKAz6EL9rFQVMvV6zYFs
pHyBaFSY9FXa3l5m/urM/MpHEEWFcXyTxsiFrNLcvmz/QrrZ7KBCzIsF8c2G4W2y
edV2KLBBaE9vPKEPeaYFGm7gQ+Cs3A4j/IPEqzDxB1iJJRXTo37M8VOAyKSpF3Wx
BMIwQDDPZJSlogdBaKH3NJtiq450cBtMeeEi0AA7DuKAV2RkzqZHFPHLPSVz30IZ
ij6dwoAc5dtmZ8Em9761kSOqBJVSe0OWTviKCAWAIengml+VgNZ3fAD1h9MUhhrr
+REwSasw4KpXeK+Vpjd2YA8xOQm3obEmJH8Q7gWK0ZZedaJ0N6f6JCN7cWdmomQJ
VQ0CWkVFM4SaWL7Q0qCMCKkxlSlgKHJBAri2xAQMXH17DFJHYJG7+3IXLITcJc51
66T+aNruAILfKT51HFgeAR6fcDkSiQKVYae0Pha92x2ymyUUswY8rGhtmtzxzKGB
04XRa2rJJRQXZucFBzXjfsEuMH1zwYcgQw0de1/3+ggWn3lvVnbU0WgB6wPQAdi0
vrQY/59lDYw9ffr4T9h/XHnGUlIgcoAhhpqZWnTJlWvt0xZgI+wVq+o3dyICG6Td
mA9MyHW9m3HLaoQyfzubITWK9LOyoGkORAlFumF/lCd4hwLPy5EMdqaONRqBQYe6
MVq5kEN3E85dnYXiXKVDUj7wU3tDL3lIMuhMYegWw95W/4FQ+G3VXeRIJcBvlwxG
xGizJF6RwWTPrczGQBrf7iBswRTQ02Vt+xUAFjW+BKiXdAUqYZyxxFAFz37Afzc8
augbDFbGrcW7uWOZ9IJ368Trij7okk7GCibfLLrCTBEioOEFmF8Ltr8DZlqF5Yi1
kuxqaNXQwXKEya8NWKdkzI3pZtqY/9EIodiBdeQQqpdyaaVpBeRlwtStXD2WHsIh
p5luwTk3YWIs9SXR+FrrrK873j5sACg1Gk64/D4RMyOXXy3rVKj/QcCk5i+JAjkH
V5fG4v54iH7lwUIA0cowLOYCXZDNdgixPWR+Pv1H2nG7yhS4Vqlq8digY07hcXak
wgsxCsw54IjW/07hmGrSAvXa0Gj3e4RjRxgG3wNWVmJS7QElMGNPOj4aQE5En51b
bVxup7bIMaqf+V8m8rsoQteQmr2AhlkbskfFCbs6f9ZSXscFaJgIajnrKBzM+83G
zXQ8agEHj8dJwsVGT7oQMrgEsllcNiVynXq3XthW3c8TppV+XaWvxUKV5Pv52yAS
sM1KUzJeit2nGvIhLNLm4UnsQGZXveoT1GCtAsvrUoPuXUkSoG9sae0Jm9TPBGDZ
nqq9tEgdLl4CqKaEeCTPfhMhQLUzfi21YObVNuSL31b5gpGlfypC1hZcLkbePYRN
+MCpXkwuUq0hgsF/3y9aPavPtbYxZMmzxMiPJvaOSuVWjEK1q+RFriDkVelhVCHg
yQOvapWHStxl73YMWzBvpJlCQIKkiJtWSoI4YcGds8vu8KyT0fYl3flHvcOVC1MN
z/KzRq+RSxldz6fOWs4gtnGVpSNB0dnDvC1VosnD/cGGrOVNbopOekQy/RugYSdF
Za2Ni3NrUs2+ECiRd9yamY0sxSeJTp0kz/6CmiyBRFndW+5LXgRmVt8DMk5fqVM6
u7/rsaZtcj9Gm0D+u3vaL4+QjTyLhcLp6qbcGKAwxbk4zlEoAsWtDpKhWhyQChKQ
8lF38KXE+Pc+us1pmjsybSxB2joadlWQPlUrML3jKdXrBHQxSzGsiAjXQ8Oy28b3
nM7sc8oyb3EmhBIgsTLMqUYHgWzmsdQCWhYUvMe5GpMLoYY0ywytY9oYaRtkbPA4
HJ66QkWb9a6vOa0l2zUQEAKZcYF+GBhJQxP4jaYS0xWDvZeQQLeh7M/WlmBak8a4
F/wSzbp3dOsBoQFfv3lj3V47XniVCmIEsY8TAbVQlnbfZyiRwNtXQyJBwii40YP/
1OJJhJwm/pdzVr5G9URf2h+SnC2NN8pAUveWzy0ALBfh1NmYA4ElVsNiqhAU2OXi
7QHKmoU27hoN4Be+yhJfuL81pC1A7lwK3AaJa8MWKcaypIBtfp++fvqrazILdGp2
bktZGQ8zigi56qpeWwD066uXeFGKo3AB/lV1H2rWqnnmrCRai6vt3By3CVb0dQAW
D5QHOHrR63ytXWvDKmccng9kGvc1JjJAeOq60phjXmm2pwv4DVGeB390QzbXjc5Z
MqU1rvIkyPiwHOmO72zGx20GN+r7yiIfQw9glNEsxI2APFbybNCkUMmxJ3yZxfT3
Ry2Sbub/e6muGbTSlfkYlD+5zq2lU/1XHlOZutiKavXEyx7fBP7yLpuSUvjys1Mr
QaT2lEWpJ5I0ylutslFNg5IIkUqNUCGVLVBPWQeT3L6EPCt8bxTIBSprZT4myGvZ
OoACDgQYD0IPJAfMlLNE9jHbkrLugDsbfNV9uwRYH/jP7bMY0PHdI3Cpsx2HGyUt
OOI4lMKq5rooV3kzuLY5io2PwOAqCTHMtOJnxRmFEZJczVnt4xJrxeHEwI5X3RLl
YLBJyaqBzsH8gYC5vARNUB2kGH1ziTfDwzEIhve3BYhevmzOiwnOF9Vzbdylioik
MU9lVZ+3lWv3lO4sCblzquJAf/lky8OZFK0Q/8ph8uEuTGryr9uzk/TJ5+vjZTtw
KgrHx6gXlWGy1aQ6k+gJBAKsBHir5uSpq/Uen8R0roHzy2AGMWwhTthmFoK0b+I4
M5Pt1GQBdgS185LamomHmAZ+ezyJeXn8NWKtW65QNPkhQT7HacNr1Q5qb/8EDYL8
CPdGFLVgcZvypTAwqbK0L4uGrqHM5JzPfttiDGvHiUi8TaVE8ik+rbtXUOify3wC
hzx9OiYK4MZpWmPh3a5VRaEvVrHgQU/QzNwmTiPykCwb/0CSC5z/1r7eel4jv1tP
QCc77JTf6hHeflh4WwbIhbz9jqjki5cKRXktJUmjoPCWPg11O0W1QDmZsNykn3v/
eHizsQsnn+bCZKLan1lJBnwG3OqH/LDR1r8Mg4ayzkHtQnitbcNtbcHbRltorTqr
guqOezQhgB7QVAZkzNINd5bTfjfqGaqRr1wGQvPeKcqgSNzxL3sVf9IQNbnrfQq4
OxE+gENrO928Jvil7EIM4CX/c95MpLALTDC12ElPs/6c30hV1aUTyQJOga93IZME
Nrtqf712oZQsszJGL7VkWwFZoblvftdEMkShT89REocDW4GSXB9eXvzyFCiBzm+2
v8n7cMWQQam3ybV1/vYRSURQOFZ4/zdRqfx+rIk/fZl/sSr+Gyd1OvDuWozdPkK8
m6eGyPWbq2g5MF1B66EaX0Honk1iEs40WVEijoqdQ+2YE81LctvyGFMiso06tYAA
g5FQL+QdwelQXYDwYYQ7qN0FK+KaNzWWEj53+eex1wKJqgxAmPPOoCdo1O5bYpM+
9g7TejI+xBScTqaJqAcyvLWNkYOFwOuzYj3SsgP467+8y14F501GNya3TxWeIrcg
TgLyOdu+95w5trM8GfOy5tgfMDZNtuh1JaXsy+eDTtaroxIgbHHqgN1wehLAZGO0
H94K6BgGesp/rKrtjBNtW1Gs8XaJH4zwP+FJeQ/eoh3XNaGacIKGsmoiZMnJiZ3Z
KjKoRkj9ThRWI5cA9p8nRivMdK+mdo2EpPE1x0LQQiNR7VrjtXm5rYPcXsPYYk6c
nEZITFhQdaclPky31R2kPot5IwFdeUx5aymp4kbmSUcSx1VJKX0bYWQfX2zOqMfG
C4JxIbLFnfF2ui8JJFTmW7QcYdcWQZde3vIRug857cFiWj9Ktzncd2PswA8hKRUo
3kFqmAMMDuYI3HZpO0ldWQEZ++BcMXFXnD1NPlwmWstALU2WVEdyh3Iw+3QeSg/5
ew+lee4iV74VeuFtNs72Glk23bSqFFgwneOQJLuDA8SeivsiTXtWg5DPFdY0ntG2
+wQ5u4AMCdh3qmFDqZ3tbd3VZ8pq6ypUrsnVwd6Aw6bBFf3KvEkyIRcinGDi0w9r
O1kV58XXKeROvkbOPkzlZJwwjOrCZNnZdyVuL9Okj/XW2inEtbj8dfY+mABwjO36
aXQL+8IOTF7EHaWKrvnyF5Tt+dXSgIrzmreBBjRI9HVVPiGy9tM8QIYpFCk6YZki
Y2bfNDdh09XvzkVTgoXYXgCHaAR06UcJiRviJ4SLVbOAn3kKcmiTfMHJj0NYmqzo
ftY0dW61wRAgeDEb5zxfDV2rYtxp9lqAQgI8/zs1PwXjOQPG/BY0YU2auDk99gsd
8HMIYnv299rHUR9LaSgntFVyhcgEYNgqYeqvelDkkwNYCUPW+N/3ASKI6+CY5T5A
ntGQBVlyvNho3akAqaRTActxPQudT4pX4Yc59j7xfmWuM254UdP/fQiD5UG8/DYX
2vozJgw0jDQlZaRl9h2CxTijksdi82uGmQNXrfJDafNTmoZuGbfzeRBetXN9RPa4
ydAt9FMZccF8gwIGuyq/pG6AekDK1I1EtdPATr1SgQYE6jh8Vq6QHqelBi7B9xCx
nf2m5O7wJsxC1s10j7YR9jPmfDR131ShlyeCkWYzGQvaQi/g9xQo22YElBrEhMv6
1WiaYv7FgCg0VcPWHPSs1XdJ/cwUAcjtTbgD15VKcNsw174yFSbO48sn6XEe0ZvO
3LJPT91o/OFjqdr38jUVFOf/P22hLvR8hIfuKnX/6AFmG3o/V1oQvLU9l7LHNWwU
bPdnUIoBCwOt52u507eCwIsV26gewxshuZmJoALwl5mZoNCN2dXUBEmtSkS9B0Op
RH9cleh9Ry1izWWp15raUCpKlysX9t1GGKmoPcN2ARbvbOvObXxvA6OrLBOak3ke
Aq+K2CGL5fyM3hm7NkEqlPCAPLUzEvL/Z5Nk7wBLG/BrXCOjqE4H2ZnK3U7FtGcH
77pf2KyukQxvvMH395QLjh9oyKpA6K3fyDjdyc2QSXgpUkg9RlCfXVs5VGPGjine
FVd3AQy6eGYnb6C4UxmQC/WHcdhwraWI06r17x8unvC4MqSdnqcdY5x2WcatFfYT
JojPyjQ4W8Os8vdwPov+pPVJNdLEzyHh8h0Ar07KcArOlJVG0Fgp5eWTBFUvoF/j
mR64A5xG41B/GsTEAPCzQ3RmIGYbMw7no+9Nt0Z21+iPyToCyrJ1pYD7czTa+EtW
j08Co2blwgyBEpPtlDVW5rCMaPBTStLh2fchru5Azc9IxEfvgxtcgE2sYIlhkDih
LPUVgzOg98gk/FDz7Xn3HAN1MvKnJu5K8phfvybBZ4tPW9EtTjHBpldUwXKJEdnm
NLUdJMpWTx35AEuxnzQLc3M+mdnGhu3ybHzecG+CZNTx6TmkpXd6JFo99HboJIj/
c4NgSLHIPZQ3PTG1CEkbXiWDVp6iQVyVhvFRCgYkKfOcjlN6a4Pvug+moy4C+5Mz
NIZWR8g8rrdiBREIXqHVM5NUUfAf+gKODbRPMLHdugB1tElYSdaw9fkN/gBmFDFX
fBcMlsRUYdxAq1VJ7CJtpNDlr5N+KO8Z5ANwi/QecOuBCGSDpJxoBdpMI+rOgQxd
ya4MUdR9F2T2s+W2DF1iJg9Q/14YrMkkkQwyMfecMIa+gKyMRmoqvAyjWBxaPNqL
hHKTHo9a+UQ3NruK9fRZxWqnpdQ4a4c0TwkwTh5fZR3e/+VJAnh533SqxXa3m99z
3NNabQPGqaxD34LHwN82jTzhIuwwxAzJ1ZEaJs+1c//2uBdgUiXLIlgI5gsm/WLH
0/xHAcvNjlXP0V062yPLrbzYWAFblBuFOJrNhgCco5LKbHLfep7MLbRErpEjdxbH
I8lO4byiWaRRdfThYypajNi7GpzVjmREXch5yxG+IrhZoQO+Ae/3X0Q6FJUW2VPg
hXl7ttrFeeKjgDpj80qihRVlrjbULQ7Bk2h8F0pV/PS+RFy1m4GswR4eekDu7wE9
KFwSCYFvBwpyC/O7SWTWnHCSV8UR4Y6EdZTSGCVztglV6cGM6h0PonUkoVK/tHBg
YK0JDgftWnEpwZf1K0D+4ZJIuYmSS3YxmrpbwVOzCBwhiEx3IUlEG1tdOLM1xSGy
XlrfMaIvxxM4LX1SDU7tgmT3ju16juck3W9/iG0RqPPmvGFE9VLp5TmZ1p6Li3Gi
tDnqNeDYpB84qsQNMnGkbhcnKqNiyQh4poIr+Zstzj4luH1kTwmHkT1Y/dNUolMD
GwHKCb5CFgjmgWIMEpP7xHJE5JKotpokQ+N3q9gu7rWoXKXr4CUat120oCcFa5TY
MZO4aLl74x3O4ND3M9vpWomd7Xs3ADM9JNrrukaX5CDrKM+U1LDsTg/DyQnA3jcp
bDSkTpwOT1EI61Y0VtcXsXGc4dOZgGvnZaNGOr9LxKqe1FIyDe1uqEH5+pgQWqmh
h0CjtTejwuQdKxktoUkhlYgGXYnGHEP64OtaJcHit9Bc4YA9fY24vZPUfUUgmbSp
g8lJelfAXsq/IZWY8n9/iEJcBrDjEmjlNbvC6EWWLd+8+DKPcjow0Y9KmdDMgW07
NVVo6ppWf+zfkrsqfMsWxqq97ku/3enaag76YAF3Nyw18ygLrgEfhA4k5M2AcjIN
LLgXJvEV9iznQ/c5TlsWb1zzFIeooQeeToCkrgot7X+JUtQyl4qAjbQLGUOZAes0
XT+yY4hPYfsuyj2swdF9KKbdRYZHAAs0ZJBraxSjGDmTaj6ggeUv1PeFEEMmnlX0
pDDclUUiVMXQ41962vyrf16+ZS/ueuOF6tG94DdmU0JU2gVla6xlEi7pZDyrFfVI
RMs6RoP1F4LWO+vk6/thk2HQTyL93ikcW81dMOfoHyB9CpB1yD2QJcpCAWGS5xd6
rKWFqwkqX4o89lNJYo27PsNZ/PkA1rgRihAyW0C8d7b8nJdNl1akxc+5YKjis+7s
ykrMORuY4X0PQqWXUZdH6vGONJJa2ohAm/T0ZTFHn1R7rxsgIh1gFz+8GFuXOTJt
y8r4vfSD9t/Df2V5M0JnHBe/HJFbP1sG2+0Y9tZuTor2slkqZ0URmu5EPbAWQfLp
yEJXi1OqSqHHKUyt3AGiefLa1h1bwJ4QkOjPpxvoJ13APUxJ/y9GNvalfoGMNHgm
NPI6PlJ4VPGkCuWckFU1fADDMUshYMgWL9U4HNg0BASJA0WqKXyBxm8jL5Jh8ozR
jGS096LTJgAu6aD/4Zx+kv8X2eiPHB7rwMpbf66Gd42rLW6qeg9cKq2QOhC2b94C
Bo7ltVY8laovdh6kCEJn5BCxGQXWRZ4SPjQD+9Y9+/d5+moCnufNFxZVIX6gG45L
jlKy5UPBr4v01+RZVXh6YCVmoYLv4sXyRckZ0P6Mo9U/0PkSD215k/qdwA1/u3O7
cPErHPypVqp6+zxROrFy8yy1lFZLTaXOpFMYWQE2oHd7CWYbhwc1nwMwQS4R6kFr
2Ukeg27dPDSd/6eeW/5mv7iwp2iy69hFtHw0yVHg+0ab78GjI/IPskKqxc4Tp4qg
bOCyiTMo4LJRc0honNwk0UV8puTR41k2hEvJLMQePZKStUWD1tfxY1QYQJburMUj
lrTXtP6dGQWtRK54wYixbYfRcZcy+/rFa9RCmm0E9MSarf4WwCfzxfCXdTIyAgAk
ihK/tSG36LzgHv3hfQ4plq4f9caiobZ1nqOxLHsFsGeppCIdu0Bpp6mBe6iHyXTO
oDy3i9Awps3oVAf6gOmeBdqNJr4/M3CBng1sp9ChHo1nBu5H2vHecHXFjKUPFHd2
V/7Y4A3ld0nQ8CTfS7twTStmI6AsHmImRbhM1j0UbO7cWkaUVeTe3HFwXQOOlC8g
4df/1R+Rl54OrlZzCbT3uzzJZpU9qhuQtHyU39u6iuggoVu7mEZYXf3Zj0uNdkpO
KbcmnCVwNim7RdVOEL9RH2m3HT7iNWPxIUKY9mc5gBs82ibv5N2i9KL4arr34xL9
AqeYP7u8xQEeKZooHsM8c9EI5XXM5emgQCfu0xxYNse+/aQX6XZ5Tv1QHY/eVYoH
MFmxPIE2VLj8k7+ZsLSHtNaA6GVLevupTLK0a6Vp0hxFqHy2AxKk6iTOPLBirivI
xdF8C12Di1E3FIXmO5Kg7ZFia44WMrrs9I1urmPyzvJ50lNB1O7JEN3L/8W67ZNL
w7O+rr1ksxxnVzKA4kEEK5tvL507xCylWVnQMan5xptjAHmvuZ9Sk3FilGsB63Zt
JDwsapoFrgD5FYUft45MK67HFYyqegbPorjTrF2CKNE6IUO6+l31a2VUmNmSjsiz
SnyK4EU/fHswwFMgRRXkchvuj+PCCgCNDjxoXt9x6imp23ZGlIiwK/nkhCTNopa9
Cz8t4E0/Sx0LVIx0wt5cmEmguvXvWLisMvhPgkBlIwcSDkDdB4Nb1O3LvR4zH7VB
Te+w7JB3aRnxS918APO3P3u+Djsa320wZa/QuJ9q7kCYXpxeU+NqonqGbDfV65n4
EMwc2lZzUY1Ve1MawW97U+9WfZ3qzksBoeVj8F4ejqRjreEBJMUn10lsNGEvyhIZ
RSS1pgn4tw2AncyB3ciNUK0w6cC9iqt5nlI9Y3pS5KmuTcdHr7WgFtbAKB3nkCOM
sixBcWctgjc1QqSxrN8U0GE+R3nzCnqVDH8NuHfL2F+7/pKQfGxCBEX2dMBsBORu
4XTCZsONB9XXNs+PQCQVrNh0isdUMEuFg7dQYY/NxOauwXJFEhXRVCyJqVol9zvv
B4y3uwCyOxKdL++4LZOopQE0S/a51bBldiHtytmXIWV8fWKFjjCjZUnkirjNVaRd
ktcEXtAeFes/N1WBblzuooNdxtV0+kN1YRtQ9dpsB+1QtXKNkDNQTgg4DHcXe3mP
9Ib/lkiJrmEJtVKUFidKDcpWUlK+lm83VCBTY32iDeyY6utzBPcYQM3TXyqco4vx
k59j45EdSZcck1byE5hK/tOVC9cDLOo1qlJ34p135wgUROb8sjc6xjIbildBmwfi
ghZd9StJxHxMt2PkWBcyodUlQQivNzeW9gjhjuLygXIFAHLr/3swmBR+cgsIqqGN
pjQ6hmBMCF2SiSa/DJyKgweVqcBvl8/8IG2HCjflt7W7hYuPcO3mR9QS2Zh8otuV
Dyr/GuExrhLRLpK2BtuTRkrhiDhpPKrhM/WnkJFoB5dMaoA6gerriCq/7t9k6+gH
0X0D7U9yd60bDkxPquhEHy1NX7hGDU+8+EXMqbIv+ZH4QVx7+sZnPbwzOIEotsnU
9nXbBBJsjfRhwiNH0lQdrnO6No+mDGh3NrJLxk1Q8tce91Sls8+G/ICpNd4X2tcB
a0OM4ahGvJ7mktQ7FdrVNOlW+lpmH5ZvVMdSe7YIXvM0m3wqwOxF9JrVcdTLkqR9
bxgNq3J/lW2dTW4woxISdPjMPh71wzFd9zk7n39dLdv6YLsPP1ktNTGtjLOlTWB0
81+DG2Yi1jnVjtuGOoPJkhJAvyDCGk1MFzv9V8CpKio90npzhhKWmwtWtsCyMU3C
chpoLSm0oDMWDnY8f/pXGzJTaK1c79WUFmr8nsRc8vzGhREfPBA51pcAL2WRUO60
RdAaRvr0EoRZEOLhQ+4dlvVoEgiERrnPgnhOiWDzvBI57qGBQeY1mtCiAWdhh9hk
1EID175vmXFhLndHDU+HMOay4zXHsfcQQCCtVKimr2YGD0msr02GTMVhp8bnuTD0
A7Is1GzrMjq0yymbLnrYzE9hzqM41P3GL4Mk3sZg1SmbgQ3qo5BJd7nqeAhh3vKP
KBat7J/BzOCe21WMh5FAP90+ELIt/VSz12HYtm93v/kd0NSKWvAUje/JU+hGXmYO
6H+uv2SCXD+Y2FXCzcCeAg/zIFSfD/0Ipi936ps79MR6OnSkKu99mx01fo29jPiA
Z+zid2vDz2TNwyk5DGt3hqUErX2LP86B26FVa0BUCHQUFoFpNSKnTeDqyBcR3hE5
QK1BZgyyt8EW9bBT5G9sXWbhlTyACcVg7oKJxo9zBEzf3dmIIIu3IE0Aqu2xhkCH
JDYjzth8ZZCjw9iBmJPL+Lmmw88hI6ScymP0zq9GrLDouR1xUHU0v4RvRRP+uwBK
qHWbV33tlPVptLMd8FmRDYcuv0zrK4pZxLK0kLxpEI4SOEXc1F68pBP5nW2PpwLE
MFTt8fZsPyRuiFujC7nzeoa+a5OROnKaFkO0skEq9lZ8fz39wrMjYFTrNMtBFi8F
kj43kry6dYU9hO3PBI6/OpG5TwIeDdRnINbaE/cnBY0d8kbi23IBya/+6/yHQDat
M616zAuqsOLLT+FPPjHkx4ufIYm26md63obtPJ49Mik1BBWL49L1FtHzGcs32kib
6tDz23+rxsV5X1AVjvIgGZ0gVgNyttVKSkgnIS/9OZdHeMAdGmQAN1URjFE59LT2
XnWfCjxkRSg0nJ9a6DCQxKEKcsPSnLtEHtZ4Iobr6aSCViwDHo0VO67qG7VTsrN2
Z3mK0PQag1tJ8sEsrafZfCHa+MNkGRBEZ/DEMfVKM7huY7/47xxP3g6YwwI8bKub
SBRVi5LsQkZtKFCJYlG4ZrYFnZWFU+XnpZftKrYO2BpovlxWmGhP6i9f+fTV2yhn
br/I7xEMiGyRr3cYn45DZDoNKFhx6/dvTv5GXAiENuAzUnPOEmpJ9Lp7zU9S4HIX
bF7UP73gYAjtbWJAKkfcRnJpC9NIxLt5BQC6WgPSoU73+iQNwvEQ/M0YAva/bUil
T9gwc1o/TcY8bRM0YuoN3kpOcRti9se2KywG6/vnHKbuoWIUwOUTVcpST1JriY9A
OEb3xaW5dsD9T0ikUqKGj5SuO3WMc8hSzleYA/75GJoa2kRPpuZMNL7KHmGED9HE
c+5Dk0abfonlZ6BZXP4S7V7VRUe1iebHrxquUA11/8UKHM6uSLP5Z+kCxatWIRax
lIxLqzsHPVl5uKRrEbf4dAMvXvcCdKvpWdKJwiRQb0B9Gi5AxXSFaqhU3yzyRgb2
o1O7MH0+itPcDCbdQOiRsGsGb+wJVp+AjZnqY6RlRjxXVnS9F8AJkCFLNU71QfIa
YYlnfWiWLCs/sks8ATZqqQ505/MaXsareOhBdUyprj2/4EPAQQebbMi14HNwI2dZ
1W4542eJ0OcLh8dzXmn7qg4b7T56xRFyCMj+fuooxGiOhvXeff+fbcfvaWM3Wzb1
UvEGrQDnhOk8Ft7it/TIcHl1257cmyXYkGlEjeSzmYlvozOIP6i9AJScr99z2RY+
6Z2h5/+byQBKxFay1zuNj/waITubLbjjt/OOwGm5cmn7kqFoddiZ3lTiltaTlYAf
Aa39l+uV10PArwEiHVgGUgntvE5qimLOsxylQHdw3I8/Tvo0p+NX9gAGo3DN3t1D
BB01IummSeIeoD15tkvlwCFJfb3afgSW+tgrF80ZFsfS9cbOnpD0V7wglO559mcr
1UJE0r8BAyNB340AIjg6gJNSyUx0rIpoAoD8Vel6GNwTBRmdqeiRLU/B/FNqHedF
7iov/9oP/6Gu8nGA6uf1viEr3u88KzmcODtXSKdMOP9PM4yaYIYe//iNXkXH2+zY
B24b+MDYluoc9rOvuDrV8UjcSAxwzGrm/LNUdLdwAYbT6IalMwsLqsLQRY0jPBzM
1aoAhcSxFoKgApRamggFjXeh63x7VZ3UG3SPYSSwB1CfiF67rJ1VoBQF9Sr0J2F/
nZqjSqhFBXMNTKoSeqxm5/mBBHKIJGOEBugn4fwwm/Wn6Uhx3RUbG+1UPuAnc99G
yk36QFFBEHLwzbH1b4PZrwOR9PYyW8XAmyuVdEKF9RHyRfbynHFz+MchkUUWbVqv
QACWA55ENsRDaA5hkget4OIXRT8O588UMvQ619y4PPRK8FU7TyAIZXPOXJnz4rKz
NRGLnMw4+6ivjuxaoLCFUHQbAhzxal8ryNFUYpDXrA40FMCTueYxL7q168qh+8m1
UEm5OE5elCFJVBGRp1tmBQvRUGXLVlOjKoNnOxVtd8dWIYHhw1YA9qLDT7/yqnnQ
wGYo/iOrdQJsletWdst4bFKHc6OMOpAgGW7tp65aKBWs7SYGp5blsmJXweMv9gKg
CS/urCIBJ6i+NiwOrBCmWlN4TwyHzvF6hs0OonUItmZ8/pndXxQC7B2+gl9w2XSS
Fs+ojd8JsKLpa/4oQKfF10LI79IBvPiUf/3X50nXPCFFBIF7U9fg7fnt5aWoc5cU
rLvrQ8SVsEPj4K9RX8fv0tJUFMR+9Ms10H8oP/ANtLxIx6EkuGblRqX+zFnYqRav
ERcRx+OAQggrqQPqUItWw0JCG0R2PrruOV1H5owLNorLB0iF1qmFt5v/dSUUTVoW
JRZKJnAG4AuIAJXJvHDANpn9KSr0HbGr16beMrIaLAn+2peeHnqeuMeRWhNu6Tr8
vnyCsjzfIxAy1nqAceZ2TAgjE/rMHr3QrxE0LAuVTun9gAPB1UNMFkfCc+H/h9Wp
meU6xWCjzhAP0zAgB1T7cyetc8Es2Gv1oMCHP15kztSmUJsjo/gANlaVRxpaMuur
WFq743Sw/KCxstatjC2/Cb72Uxjjn75r/zMxEdUJJNLQgVUmkMArmnxPYJna519q
yag9YmEjsqogj80PFWoaJlYz57IcIXoNzNTSOHlGFQKe7esbiWk7uz3PP2ShpxLx
8xTD5N52r18937vd/jjr4c1onD4rzDX2PwWUhZ1uDmPqEey3hEvYQ+BLpNnm0aSp
IZ+IvyuBLSH6qGWcg6DEbTDP0/Lb6382kzy2kjIRRVzIEOkAIx2EwokoQwcxoWCf
91S4rICgWZ/7K1R1Or5IYmraYzAsEqD2Tt0gKbfw25xr1K+v9X0zXoz7CH25rTQd
Mj5zJBXaZzK/qs5dCfHf4PZZzbUuWWk7eZywIijiEL5EnbpWcDQNn2rHdip2J5xA
VMzXB7sKn76JmSkFcCRqqmscB7yGHEFWxN4A4Uzgw4AhJBHIkLI/Kt1xIqiy5c/G
CWrUTQ6pEt1cSTzv6v5mZkO6R3UGHM/DIEPHu3+F8v/nsmnbanyp4s5HFxhcy/yK
4g+hcGm47uEBD7fVJ4nrrZnEJmXIiF34yfSMBVL6u382M5iL8xt3//6JuP48v8Ev
5lQWGDaSc4TglSH/a1OCycCM0rfMC9Mg7VqEGwPF30mn16mlSDUX9kd7u20AyKAU
x9qTrNCjQr7yKVjCqBRz7lHsLda6VV/qpgPyaLH8O5LtVQgtiKEHhdjHPKXIvbh2
HdfpdAcBbBWYltOz0HdPOZjRaM/YxkjdRfWFRYkZbAlxanbAx9PnwmzWCj/PD51P
LbBvml3yVOwLsBlGrtqf9lk8OYWAhudcKJrpEQLEwQLXaWkNC7oLfUGp2vS9S7TT
N/pPWRkfk6nTC75NDkiVH9Aj1VmZs6hbNFmPm2MUuXyuXOxie/N0EBJG3AlMpOOF
Z2klK/6k0V1d+BAvzR3ze+GIlxGTjoyGkL5DnqWhB46/JlRh7yxLPWB9+lMj3VZg
TqfedC/gEDvKxnzMP4hkd6rjWOUIMzRFaNzmP5qCY8QUkIW1X5XKwtIn0Pu8vRk+
X513C4DUy8KXwM0Y74Tm8E+8lQRfwc1zWqcO0bKhiUV+H9tezL5YkpXLesfHzdmY
go5QbBxOatgsx6JvPEOe7KSXc4c6D9ZD25PYGBDfXtYVBI4kFLCXnTW5TG7wAtdR
rKzXJlpbKKXquf9GvjILDTrKImO8qJyizV9cSzq4j9tB88idaPTDwrUVfptF6Ifz
L3Pud3pB8eDPEC9SL/r3wArZajOihM6OzRbIgjXEBhVMYjkrAZk+2buo76VWbEMo
+XmFczSiosY9PlICdGMkJMUZJObCNm8uma5PRnlvliU+DtTB9UpRxpbBQ03ZXuLb
c9oBHGbap0a4nIXSPUURu+WHWeEizWE1bwCdQTj86uxzysqW1PP2OO8dGjjnpsfQ
mBD5zlb8Hy/4smm8T+NRdzp3Ybh6+ExbA1oPvZWRpZ9pwYNzWNImnv3AdvOVGwLB
EDA43OglzsIwc/R/z0KpHLhiGNY1maao+em6pJV2SXQdJ/Y1GV8zbVE2eswHjOHA
MdZ6MpqwHTY5fWA1JsPuS/DWEbYOA6wKhpEU4BOYqZ/b6vF++B7rAgHW4fzqOgRA
l9nhFFqRzImWJPc4JYEn2PVqSe0Esh9NeUNF9ZIDHR2YXeTf6vlLzj3yDzIYZIPv
Ig+jarsU4ZSKJR206dtwZNysVKaVvbgRu619HkfMMwL6jP2rzQk1ajqpACiUbsKS
qUDgSArgLPTWlbPhh0xd0/4CT7fFfu/jgIXhYN0pgKIheN6+mblE8yS2IhMfL+nG
oF+QWlyiNx6p8Z+K6NZ4P+CdbZQEChk1ZTJHeafyFVYD+GMPlGaB52JsF7Yp7FeD
5hm2jILN5aPQaiQ71htrOhI5+b/3VpCFpLSTPGklv/TMLGasyDxwnXy3GDHUAa3S
RCmDtKnpubpU0nGamijcEPqc3ETQAnxYqm1BXQs+ZB8xenQrJ/65EcnXToAOenLI
40IKPETIlaC7ZR9t/3jQXqlcSVHL6PeawBp5DO5lZ+gSePDlda7PY+uojH5BoSsn
WMb14Y/GliRh+pPz7unRfE2cYZM6PqBFAfA59DVA5x89vu2aMbYzsYfTfhxY6n6h
yp7iQn4rMY2JX18M0ob1pqOll8STTbvsNAjmp/ego/i0JdBbFpGnQVMUdIeLtnpX
jGtKRVzqxYCP8zpl3MfP3LEPo3tSpW+mF7LrT2t4bID758c2/yOJlE08saclxyCs
aa4MklASEFaI5aPRuQ4TA3FFKyCkSw4G8IC1vWi5QCXwhUrv+azZT++/WghT4jVI
AUDqWosgJpTCYklSEj99/VSWQdpukZ9/IpMiZqk4q2pB4oX4qHK/exqlKaWqi4wj
fYoyXc1PXGZxZpsDECmyjSIsszrXM8vC574pN2rGsfO6+jYF8Mba5WPAB6fqTn+1
moWR9NvHPOy4QNlUV2pdvmk7v60wgoNM8nAfuovVvdaZzS14/nNRtcnnOskFEVQt
SYd/o/6qeUQqgI0SnakSeOAgeUhywyI9+FB5osQLuDE+fitCwZLuGMVe5FuBL3sg
MfE6vB8HB6FFp1MZrF6QjD95I4ygFeTXJSR/vaYZSHTy4zwBANt46kdSy7nrI0IS
QQf2vNIem2tet5GZbFfiGmz3PNz+R2wjbCHboP9s3LQfJ+o2j+7wgMD3IgQFXCWX
nXJRr6Gkc0BWoqEiAG3C5MJjUxojOR3ldfXpZWpz1us9ZaLgtM3F+DTLesBiITGD
tX8rx9NAwBn9GsJ5od38e8ZLPSgSD5JDcGKaxnBWNcTFDYTb13cK20l2baLM4057
aeSMTA56NXj6ueFd90bUzyn5FuSvS16VOoUbl9yZHvxy2L0YgDLIieWbjlUuAbxV
5Qb9jzjPa1A2df+2Ilb9nqGsoEawKmqZcV16H/CUgCPT/G47fUatbAR59P5asaJE
42+DSsk07QyczYBJIZMvYK1US3zWUJU89/c6PlMN02yiYrT5jLF6R7JJoW4sfeU3
5ctyaq6AtYAwNJTKI14gw547McstzZXyCiaTYtDjYrV5iIBbOvNmMjuDWNo0+24B
RLvt6ikmRAIIohXOn4U7qIXHMSSr0c9Clbb6hGsum99rd1iQAstI507WQu/acyfB
2ufPpHbx2SBILJrFHlFUbhY0oZ7mebmbW8PK2UNNabqh0gjVaUN+q9Kv2TFd3Vis
8k14FAs7lLpQUEo0LnB1CE31OiOmmIazc6LbAlXFzXddjtlKOuwaiu23fD64RY1P
B12X6JWGuJoSQQQWny0v3AijDlOnbrzCfnZ7ayJjd/nGqLwymng/YQxd1WRKaxX4
MI+tKe8BMyOdq4k+hYsHRwvePHz5q4VW2DCor1z6NNejP9ueHULahxyP5qd9RMlb
lYsJOgxQYHGrTcwA0ARdEoRWdhSHU6vvp8i9zZw0Q+iQjwEvbg3aw4bRa0VHKiR3
KhTL+uK5J/PrZdQdTJyt0y04UzAoQCHXAPiXjUwC6jGKVXRnEOiNO2aTpqnZxvqH
Xpd28raF0HIhDAX9XWEscjYIm4a8bZS3hSOL3g+5hGtF8LK4XGuEZRlO13s+rY/Y
xIAzVpAIllhWNk2AzSeafe1XoXfNeQvhaS8nIMcWEgE3rRhedCQTsg9axGdRhvcw
JJtmrqaeEOzv4JAWizSCW3RHpdllNxcrAgGkoQNpmHkMhx/je+8A0heTsK8+ZFlG
8o+OBpuQXswDJuRTB+UB6b5VDaUUpG+D9NFXSgg2g19ZkUPmAJTbIVmdmX5SXtP2
U15M2Ko0jTwLfBDwKO7EK9jj5jbhxnIlfdvmeiBT1+hVTYEijuROpo+lplBj02PB
kK4QidVBbCUdpfOqcXIyPGjLV/stpZ/lZTpNoQz2Lk+n2fgpysk9UyAYZfSUF6b0
1Lm8maGS6DkeOd9c/BB/lpM58H5PbLWQ0SSBV6jX8KDG4n6Ck0ErnhqXJFlujfWa
m7RTnq7WwDa0y2bxBqR33KYpBWRbbpOHHbdeXVKJs65hl524PWHWkYchljvJ4RS6
1d+zV4Nd5PQrERvTQ2hFnBeBNH2YNRDucHiY7fbZH/nmzYs6vz8PGVtFp7Yzf9nP
lE3cj0MKHmTE+47NqJRWwjTqNttXNvWPzcPVBskQvUF8vg3iT56KCDf0E91WndMl
WVpoQQYGsnNkzAdWo6Nz9UlnuaOcSKnGMCUW5s/UB8F9GOWb1dnUEJI2FO/D1YvL
pqKh646xXd4gbNFZnERbZgHPB443B+OAQWaVUoQ/l6jkZm7GtS6a6rXD+zGCMEUo
JpolGaZHhKhhtLYEcp+Z2oFPEaPxt2kh0oPEn8I3PcBYmPepLORANu7hYJNq5Rin
sHamW+OgtUFAhjJI+rCJzpXOn6QwO1ICzwGyN8/0YqunH0mhbb2w1hvfatygIdub
hkHdlv+azJ8GPvLX1YH1OtXNEYKtSwDxpnaH3U95XfxettKK7/9JI7K0bbpJFlI5
jDTYu2WKZxCilgWv2r4eQJu3648yqU85MBIRiqaCWv4vpJ/XT/QiQya6nTyThYVc
3RPVLVefw24aieszh2N1Tfxk8ZejqxVGG+bLExnbGYbbYwQgtgDa2jCQjZsYT7Dk
yd6q7EIdeOM/WcAtULge0Gy9aPQ6kZZuRgR4ajMwaACfMeL20xs51BQ44zuIQ2oo
mthAzJFXOnv+1Cw43Lz4WJdPpHws1OnQPeasjGyw6gisx9iJxxRtvPywXcatVPJg
t9I1ItS3FredHJHtQ6A6C4RiLrQWl9pwANiPURd8dSGAJqVA/ktpF/7940zgNuKg
5ZUt2W9p+STKvHwPamOfnW/FH1QqrhasHoES1qKckQIBzJ5XXt8JBadrbdThYy07
6rHRPBcRU8phMCphoGcWmQIyncb8u5ydIBM3Qgzasma9+s5GPAzWNRB5WoMx0nGz
2lfn6ui3HDQK1rhuvDM0LO3XTvCZ4hfBVbkKRYckyD0OO4TJ9gXhtsd/wdm/T0r7
FLgaS7N2Y+Xkvraw5wm1WFVSYo+x8CfJEBUcVVNjSARzQ+pK042OYzMmZDwMuMio
R4/6NiuKUyYXPvdmfd/T4n2sN5j7NYbPsWhwzsSVzfANjaF1MtGb+INqipJUVA97
LhtFH2Djtlr49mrruj0snE1gW1iQdjbOlUjre0xBdmWDryExmdIGfzEI+zJCdjJs
TfTZkiKRueTHmbO+Yi3FOkACoArKizj9F8swYJ91UQPNnF7BxJoVAsLN8hSUq6kf
Mdp4XCvju7U3KG8CziyElBDXWA4Ds/hQ8nRUhcI3RBAdz17qzkbOo0tOc6XwuPPN
jZczSYMcF0HkMOtN3S6a9fojtiXd41ocO05s7MK6o5Y09Jc+RuEY+0A3kJsKyul2
AVkOmkXz383WRVH9InPs2fsvT7t06WYYDTPlisD4dhHwP1EdsrKXH44OkAAr8zSC
roJKmxvhp1gnvh+0t8EvEC5WFzCz61NIowWmwKi2o3gUOMbAFfiMPeX+K0cj/0hl
opZImqAVeAN6ecPVm5aN1un+mh3ZJ7rEAU9w1x0WFPfmbxpfOY0xlLoxXcLyLlaE
VRlBzJ3zoUmTS1AX6ZbgtU4F1S8qIrtg0LmBL1i/4NsfjA6/ukz7S2D2y7ZWwy64
/JF8vYKjqc4jexJwM47AJesT3MJIPg+a7rLd1rszMfPcOmrx/qJgxHQFM+5QMcIQ
MpJQepksgvbawoZGYkIqSQr8dBI30H0EJ7vrGvypwJ+PnLqHFhN3J0mDxdR1bAi8
1cvwgjuGCe1OmMRHvMNHmFHTujcAA8judbPvq7W8S+opSxtjAQu8zSNImncsNI35
s9qiegQgZsfdK3qUbHGUwpfBNaw0bcrTiwWxFW71z64+IUPjqDJmIGJMBIokmKVD
P4BThe8GF0inT2enh0Q+KqE2M6Fc6a+mGsuSgs1YEBwbWpPhe8tEmu/y2kW/z4fn
xeX4tk+o+1Cl0iduqnUbLxobx5AjokZg3SAF2isUM0Zh64OD/xqbT6A6BAJOH5Kd
OKlC1pIwZaM0dLn++e/kSOedYoaovE/tH7Cr8AYdA7MDjL/GgH+TlfZT0r5iY+ZX
yVk75sF+VrVFgqbvHIx1q9g1hSNtVdTfe4dGI5vx6MIpapmoocKOJ1LeP0GirjC6
w5U9wjfDMBwUVBRjWcbrVwoYdKp06GjvZm+czLOKYEqi9FRsD9j8abvRs5m6cINx
r7KENiM1EmHrv9cARNKTKROJSpKXs0nxe9YmATM8zNS6Ajdii9FEj9Hx7u1MY7xc
4l79JAbGzOOGqBdKyhdbaOP8Rj3t8pNK3FsaWbRjsVSm+E9Z59Ct6xpBmlTz1oL4
tgk5kz4vaPYmNBygfBVtgqCkw7BcqZqlTWRAaMDdfRmJ5pWE4kZ5iVA/ZuSeXKQc
Ki5l57cyuSJZ1vNe4Cxp9FX3S8AInV5pbIl1Z0dNT2TFE5XkaIf0cbTgIC7dXn73
a56/TfNjfZld9Rwwm4j2Wy0QsUjbCenyyX+Vb+xPySmrJDoB8KVV1dkNRIYjtquH
TodsYZ4MFw+/nD739+e+6i7oNqBFhEZ5MnFj28VOfyZ8ZclzJD2wygWbcs1s9tl6
CSml9AfmA9EAOw3sVygKTyloEry0Aijwm3TEj3+YzAyU8TjDMkeKSZt0btX87rIj
3qfvoK/KGGeHkPNiokp7vfPCvb9ENftHB4ysh0o/Q0LRJIVMASW3o5d+fyJihA9/
nUtaEAvJc0tvUqHRL7jPXKm8FBLy1Uc6V39+MuIJindAjjNiAndgsm+vyxDuvsFr
c9/mGI/BrIwVaa43WgiIXT+1R+BkWcU1/nY0G1LvGmQE75YfS7G4lh8A+4doUdHv
4GMVfQ5XSRhRu1jg/n6Fmec9p7j4lrB3mx9eOsS/VsQTsVfis5ejL9FiBmukUj+S
US+TYltm3FSaLbXM82XEiT7p1Nt0V+0Gpefmos/AGR/G8g+29s6wTDDlR7v0uego
sFbkSaJpY+1cchH46XsnEwnpWl92EsZfiYuyJcUGlRyiCkzt0WNw2d1+9Sx2JyYZ
48LaCqXen/LZVgjWmv2VTzgjNpjqRC+3TFZ8o8xFcpLJ+BF3sMcTxHj2ju9WErZg
3ty35Ogc6zze+waXwtp7Q4scs8pLitTIrGTmLZBU56TEab3s8v9MS4cHA6TR3GWV
4E6s0Dj2RKsnaAT0h5bG+Kao8evwzDJfvZ67u9mo3+GwN9uqiTt/TZNeCRx+JDqe
7DUjjxh1jNxnmDByMPo7fosPFV7qE62ss+qaOuXZwO3CPykor9HTKNH9Sxd8Qqcv
WO5o5WmVv2+O8OS9PnFfOzq/C6C6LRZHuJhFopr1BEEAgr9jl1q6xai82+mGY2N+
LGnQIE69SJFlws/lB4ZTlFZx6hPbRJLGe0KfnHGhKecm2vUVQnedIPg049FBYtGa
3lITgvTex234sPy2blT3hsNXhs3pGiRTuAFrNIjqQ1XQNNcw8Pe7OiHbmE95Q2Xw
UuOWvLnOA6Wj1C/ew2Xt2EWAJApsVD3+WM+wfYfjZ2uzGny+z0PK1jG2V/0gOj+V
HnNZ6TpYLN1tDaCz1f2+SgeSdu0sRwHOeG72LXb99bgkuhLKlfaJBVWAmIbRh+G/
koU6yFoEUJhSVwkH0SyZhche/3RKiSNcN+hjbGnhKxQRSR89Dc6I1mm/0t5uTwFP
TMo6PeHzbAZvwn4V1k4xvVArmINmv0ooBNCQNYX/4MpIduMHSXNFLWH8QQJ05U7P
U1mPTvN1WZcIBzgkPXeuV/MrpA/2UkO/4KJfo6Z0IlF4GTuJ5PjZM5mNXz9reA5B
+5ZdC233x51eHLeUePVg5n3c15MMQfacmpJP6i0EB6aBGGU/RepIBpOrKWXQsTpb
HQI1zNEnFlcYGDs8iClVn3ngPUhN6Upm0qvLBKDrb1bAyOqEuB/tdrsBiz/ZogrV
iA1JkT+YA9V6Xl2ZdLjo/F/zdOBLpLbAADj0NH6vsZSA+k/a5iw3OOzpH7SZ7jO+
RFxif9vUUFSrO6XVHoEhFbia7owPPHBF1mg5akI++/7JXj81sDS+fta5pl7nCMlj
MQpJ1etrFUia0EmkqGcHdQ1NoYRNMBabFw4ZbYET5JJxKzknSTgxN9dWVeuo6Fk9
quFOuE0E7ToBiLDDT3cemconhreQdOdjQUDwjbRfp6arRAq7MbHQzJN4S4o+UEH/
v9OaN3W/jOAp+Wz/BZo0XsmUckR1BTemLlecEz5ovUPtFTwWmTE602S/xUY60Lsv
zU5edITwCANJjQPqE2MRpbfk/xuzYDNDgk9ASB9iNiGcpNTaSFpnkmfN1nqaEqy9
+sdWeNsmW9JqN8fdgStblgmDLh347Btf1VQ/ETQ/tfoVGpY/2aBNr0Xv6bFMhOWc
1ma/UevsUnCh/yrHrCSt8Q/Zo+/bL85Ls5ScjofH0biDn4zLYOh1ao636mC6Y+SR
y/B1qfMD05O5vhNs30qnpeQAlkvXm5OjSTMfIojXB+gtlkDk9VMFP4pE1RQfGx/+
38CHr21JLP2oLJSmT7jM8iwCmHbJofbh/pyinkIZgaIwsBr1tEd8K21yNpfA2OsG
0JtXHPcCKlQuSCDv+QVFNV5jt9qvy/mES8twITWzQ11qjyofJHMqrU8cORKp/qHv
NZcLjr7ZUX1NIBLUrBwli2EZDz5QVFZZkbihYqDDDD3PdrM4Yj9osrBY35000Fcg
kLiEoGHdwXuf1plMvLoM1tyUPfBcMeHRXW1+mYrlCl3XaWxYbvQNuyvz7A4Szqzs
9PYyVsb/x/d8eE2+Gbvx+oMuX76SuppawIM7+XvT/ciMZn4nBOTKOQfIupIXQkDQ
JI8B9sVZstuagQT6+JdCOCZ080jZJnOYuQgWnVXByZcx7SJLxtDI09jHliU6eYO7
ON1SJyoo3FfHV04dRvElV279td37jO2QcoHmRoKaYPa1nzL0NHEh1n8aRf7k2gPp
yuZMJ7QxwAIZsfsNEpxD/BNPzdwzfY/6stpQEav8xfNB9GA5RhhFi/vpuU/9cZIF
8rVBpRML0HLtwXgVPUwihGCEorjqLogtXDHLEehMxDwF8AIkkj8hKKEdsH0fr3Pf
HFBiMf9RRkyLzvJmIWkWQeYbzOre4wBr/68BTET3fZ6qbDO7G3/DmgWiJ/+x/hcA
BQfYMJEONI02ICT0KD7CaWDnkUdloddCPafsxYRmz0g8LiL5sDUgteDAg7G9vQux
nCl3R7XIGYZWpX0XbX8aeF5YL/ihkAMn+IUqTy2T4h0w+JJ97ALAhtgMchGghiKV
aeHl7UOUBMT2yn1uLB66bDaNY95QpIWg9Dax934tGuM7mirjhpwNPzxd/jXPNmfI
JlrkqbLrz/+o+CRQWoO1HSfmwH0f+QRXYP8sEJspbAgA4tce7pkcP4HxLU1KfL3l
/hP2lIhcn9B6s++koWUb0V09krdSIq28VAFiDSHWgQb8HUXWNbQiIkGxYTp9zdDi
auYaxYfY5Wcfd/x2WNEpCSBntlBZjp0R+rxsfb5Mi8FaP8vXO4DiEVCFZ/PQl/vl
yj2nlAbrmJuUuY5yU+d6RykSKdtRFYcGs1oD9TcDMdT7fIJkIUHWJOv8YFTqEWzU
Uvi04003B5pAsIxdTQeTOH+TQtGk9EKQB/3rj+d8P5cKboBc8T6YVgVVXAR4tr57
wc+VzhfWQaKizCc4TvcB231HmUROxqHbTUqpHnGcNK/38Ypfc2lnQ1fQYlV8idSw
amMXvxivueKPlW2FaYa4NqBie0QRYUDg1oNbluYwybCUB+i/qr+8ytlnt9pdr2kd
x+B3B1HGf5nsuXHx8N8yj7rZfttOp4Lg9rG7RG+lNYz3mFSt0v1rR9r5HThg4ldi
LefSVsiZshxrS/aZZ85pyyY+iIVHfo+Gm4BgJ9Mld2L2w3aaNCW32bEZ3tBg9j8t
b8BqPT8LPM8QjCsAasTqNJAaWv9Y2ZPkMd2TYdzwcAuNXwQ8D/P3eqWjNd+rklLt
W9YVt4TGJUdh716q1VGicyNvdBxvp7EdrqCmnaZu4ZYC0Yfvm2H6ZVmc3IGvrHxX
VVvvyHziylvw7b3cG3noQrWdDJK3+VvRQWUHQwX9VBTxS1n/jUsa1P43k5WVRvp5
VW8DLGsYZxLLE1D/Z9XCgPoWYBhjlZKb+bNzbskN11pwrkWFG+6BejhhkM7Tl6pm
AmMOHXf/zCYNQmPZwy1clson+FpTPbCfXfkNLiLlKIO6OaIY0wfC3lGcQ69WLj6B
itt60DrV+DAnGmZx59abjgpm4DkYckvgrN3y7mGYK8FBCcgsulFcTZXt2Q4YaWuJ
vPUHjVjrXLirA+1W1iVD0r8Td8mCRGInMmPTmuH5TQkvAVm8H/c6bzY9zPSP6YeC
9YhELoHCXRB9vq6JjS43h2TRyJtAVTHfMJyWuaeH5Fk5KGG/VtzPIFRHNKrik93d
bB8Yl8aLFjojOOToQA0KxyyagWUTvtjbTR2f6O1aMTDjTTzBIDfrnMxOxo4V/vhP
XfZniTQpPnY2SeobfhjNC21JKsvIu3RR4xvJ5lzYgLMhPUhFiT1F9qnJ5FWW3xni
jjVTmoX6j4RFwCHeHMk+f0mcgXkwk37NEpENEXAo2bSzpi11y7iYOGCuV2OuXvXD
24w9pcFMc6yl/+sUkN4Ij+SEYoouw0BHyP6iX1zb8X2XjNLoTtmOzuVL8AK1kW7G
v/4tw7sjiGrX6Vub7hNxQFJUgI8U7tBLPiq+SkCn868bVTIYaR0H/L3BPjTclffV
pry+0KfBhvtzVGsE20hs0wHE7nDI5d64Eq0Lr8R+DgTR+KC1Jf/uGGaZqVQriLlW
5e2DgDmW3j8fsOtr+DPa1Pid8tAdfJ3z79ZC4GdBhL7DgJwyEx7zcL7gcHPLUwOv
/kX4FU6ajyUB5RnK4sBNCTHZ8Zk+faXXP++ss/m6J6wis8Ey4E95RfXwIVkPGYnL
8Ebd8EAUnGCZj+JsALRZkwUfKKu47AkmSrByMScn2TfGiyNE7PPb/Y95w9y3nZKA
nyh8FnSdnlqcjY+bnK9+Lmqtlj9Uh6ils9zTHBUuL9JUHvPbe+ZDD8evR1XIpE3X
yxJsCVeXUGb1SEIJQ3vsfrixrrOoRHdEbY9ebNcqLrxxXkVuManwY2h3OU8UkFml
VJ6n+LApZE2zqJejbcvmWnTMKWecbaup/YXpDwb5WeNoE86G5WVoo3YZyvLgnWk3
iX4l5wjAhkDNmmzJF1UKGkBAMih6KGL91iw+UAobT5QD5YlfwmixlF1VZtUKCAuz
7bcvS8g5Z8kVw3thQmYtSzU0XNwkEj5XGz5BTQ6kbWVnNbBTkpdyfnNM/05oifvb
Ntkl5YK0DgXXy9PXz1mVQqJomibznJvTDwXsJzhD2Qj+M4hwxeTDnscqVAWx0dtc
MyxzMKguRMHaYdBIVgBESGHyb545FuCB4OuH1NCgVP/LG+/g7acFJjRyXccQroQA
6cV5hVNXXxO59egcjKQWbT9odpv+0xsAT9x4jpm4S5/lUvs8BENb9E0isF9G8uHC
zkM1RSqPgu8L1LJLFrX11SU11dcwVe8eAG/nfCEyyL0f038HQklc6ScD42+geBGR
DhjJ5oc/bzVbQFS96F1sPu+owss5t4UNzlKAn7tY63pCzsmDhWhb53t4DefysHS6
zQx8V3h2wp40SUqur5VHJjo1mK8gWgcdcUrS1A8ekcnNdYAVaxxck4cjbNAGb2nw
zziSscCVO+bE0ujqplyGhZHEDMflGk2zYsclbVuAWqheTPtQA4JTkRK8LdrYaNiH
CYyM+Cx1O5aAxlnNP9omaklrlC5PKIOjoMmznF9SqQTfiCjUAtxwv77QGi+SGykF
pHKuPKcLkmG7zBr+2lzeqHHQGp2FrON4WgfmWO9PPBWCVS8FmMQRlnjf6AgnPjyT
1zHVibmqZ5R/oxNULhT2HdZo587mCjEGykL8vRR5MtT3RoFu05tTKl3ZlyXPfcqN
5KKoaqF5Fz7TJMyFJ52VUKldWxD1QU5sUpon+2ktPy5QL2zuiDHdVsqJ5cLgJHkL
UI7yu8REKI5FklXPlPr+CfkL12xs1ykc7QO3eVZxeUyQpFntkiGUEhXcU4wxAOBp
NOe4dr4ZK+2VHAEny+t7FQ664gvqWrTNELtB4V/lHbUj2kWBgTsT8Jk43MNUZYzQ
OLFg7w9U0BozwgvLLl5ml/AoNzlq7Hm2rCJbDIZ1xc/4qidfPV7x2K0V9/yHgowv
ynQIy/kps0fdnsoCWMSNQPLXZ+dDj0Gv1GdgI7R6mciQAKgYGEG9+xAIfQLlW0Z4
VNFp/WsF83cfih1ekqDb+BZv7VeVx4gYXfhdNpvodwKptn+imCN51TSoatsv0dAz
5N9RMVLB/wqwgRFQveCgeibv4ysZgl4XALS7Ilg7uhSaYXokzrV21KDfaEucQ2Gq
HO0+E7jBt5AUsVqqipuAAMcMcgGEARKbd3DyIi6O3RIJrl1QZoGppSCu86kyWZPv
Z3d5QQo+OmsdyrftnItw+qja458hmhqDHllY2A9AHn+HrrJ/KpsoGvh+z5XVsMZo
ymXeOsK2sBe3RKbiMFmAEfQ1XpIr0QYUIM2MRdZZIRW7TyAnQ/6g0o9KG99T7g/i
23OJywrjqN8NoyUvGrq2CMxi2G85kuG4fHyE8pKmQ4T9EjbyxTOpTtV0Rn4euWo4
rRaIBq7d/6ro4Cq9S1urf1i1ZMssWwH1ZeVNjRL9H7iR2Hr14Qwhp8kdCbCIno79
Ww9rcdWGSP/m13mDIF6xpRQm8UhdGYDXjpeAbqMUEePhOoigFJYkHqQDEQG9Cp6n
czF0iRkEvFr/vRco97/OA+4paV0IRahE5otZhM9YJcJfoyW90yXbmC/Su8jeJrw4
wYXFtsHYnzDxoRn3oMXh/vwWGOYzbYcsGwZHPLYHO3y/K+gW5NfnE14KMdeJ+/t2
yg7rhhfV81euq1gikI7bW1i3egGv6cZO0bSvzHnUMrXk6vzhu4Gopgsinnr/j18j
sT4weuJe6GvB4HJq6m+H4ITP2CidvzMxSMYKviqlzDjlzwVVmElrmDl77I+z/tor
pV4JYK9sFcR2WUTwOLO1zisIF5m53ICQN2VGFDW51aQFBMzuj2lhVQq9akf+bTeG
KP+IQx6m6E8vSniRwjQJeRfN5bSCnvJNGHz2w2lK4xoiL1JO5jliRZCyCQtcREKz
n1cy/21Evu3oImHciVwjGTOCs6QcsltzeVs2jCtrqmmuFzpFlRQeq1+ebJHR5vCD
3+HQb+khzqBrD7sHswHvCQ5s6eLrbb+1hQ2v95tKUx04rtOyeRD4boUKdJwXPInm
QpdyBjxwGWjUgsQG3Tfa1ZdN9JeFD/ms1myNLUMccwT4Q+PU0RiBZRty833AMRip
d2sbTWSLc9yrsYVAZhomO96xLnsInFoS+VcG3o2kX3H66/EYLZaMBmUL7CxL25vH
mb+yp7sW3sfopZxj2dB3ZmDWOtOy7+oPbZ1+8O6t63WiXSlxUBK/Mw/wACBWyVaL
fEHjM5HFUr9i/rOWWbz2lRZsqEbGWoFn+5f04McJ7LuefZ16CL65RgyzTE0sOqnG
AxP0ubKKJ5M0VLETXIk8KZLOtub6xaZwnV1mJZ6kpb06ZL5xpWXKPDmEG1T+bati
kyMH1/BPQ6f6DlGNXtuJmmKGxSBm8fS1kawRC9TupgfRFwWzbI22Xvtd5uiIGJAU
LYtOoM5Quym0aGz+8i76ACqtWIrQDT6cEZVQvO0rWZ+qR/9KSj5tnyO73+/Xv4v9
gLTkgLR3/wOLb8ak4b0LvO8gsXPaaz/T6/9785SRTZcZ1B4NgL5WTbRDgb9dwwfP
57LGYSy9Zu9KPS0tBupi6+Jg3DN94JD1OK2hdW+gTykXCaPZGN6ZJho6HvdCFu70
ut+NHv8vA8nVxxkJrNmbhQ==
`pragma protect end_protected
