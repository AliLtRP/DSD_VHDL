// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QvjEhdhon4qbe89WU+P3X4GpE9Uq6pkZhzLZddTX1TnF8f6EZ2cPMweL7K0y9rXC
ZywBpNHL20UlqCMNLbThSb0ORCQO20uYEtAZqElL6+HrN58PQjN9wPWtjHF3GvOT
fZW4MuKACCi/mOVc6dzATa4NuSRRATeF+3g/zm2gmOI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7296)
8VvaHsrPGFpFGX1urKZ+Hl4kzcVx+0MGwyuxvkTQUYi8nJ87JIgO8Tyg3XIJ4O1G
QvWWsPiE8X70wJrNHZKtHVvSNSUlIQtMm+4NZy8MDEfaJakIcGVYpbkKrx0j5tb0
GVoe22h6S5Z+QzdHQ+hVmda6YCdfGWYKU2CksXnfbZSf1GIlL8iwoxSiPtvU2rp5
lzTFufVfqzoknwADlXX5SgCtKGKXRA4aaKKA8sOVCeOrEVAyoZmyAW1mmIWyGG/a
FfZt5Sbmd0H/7rtUryqpegrO9n2sWYzrVhlREcSrP2FCUHwwAmPjABqkp/LpBBGC
snqd/CZ5yR1vozr/b6A+bZT5w9bxgM8Crn1UcPAaKII4MRgFt7SAM9nC8CyF10xa
+XW74lqF7ndwB0PGhCaI9kVN2SuehxiZYAqL8gRjP2eJSwQZ9YEf9lFT0lhOqSUU
fjyTlgFsPBzzoxlkvU3iGnCu8wTkJ5BSHkvx5BBfHdV3rjA+yuUcH3WhrR3dVGLG
/RTyXW0R1nN7r96EtuT9WRk2WP/3Ab4kkwMorfF1KFAwtu0JzKDt6/4fkQU8wl3T
iaDgiqvjQ5HpcnXcnriCaD9F5bLlkmp8Sql+hMIty8np1I9KpIT/pVfrzAtpgLtF
8oU9WIkxo5iu6mkVy6wPdnT5T5rbaNySQzGVpLfr727rTApWcNdEZ/JGh/FcyQSm
Kh8xiqy+5yx6HJX9Xtuodg/HN7DIt7Ld0/bTnI02Rnn2D2eny911Dh4Mn2fcNPu3
txQZa1n2T75I9ZzbnV1rNwtVVS8DTmk5FkWiMsm7RFsNMbFM6Y92BNYXMCUCZEO+
NO/hwCW9jX4tfPpGLbWqxOMDmDWsowzbUVTGlRQzT+cj7RIeA3w5v+iCbI8uiI/n
OQVtwIKkj4moW6IDMwpHa+tnGo2sK50S/Eoi0GjUqVq8F3EfawsndCYH2Q7Ijonh
5LB1V62vBtMeWRACDQIUtw7vvLo8EDHRAXxFq0S1z3MG9lIApeNWY4lx06y/56hj
qWATaTS+IUGYvrBCT0df2xuHrxIbuMc82OY8m7JbNdqptxyft7tFjgdRmEV6mmKX
rnEahaNDvssber9Xs43QNLtV3QYju1tpVP0IZ7RDADE8Ol/mhpZ013E976YD1UK1
HAXhhkBzf8z6xmlug4+qmBLgaVfdv9nW/unS+ThU5Oxcd/IonbE/HJfFEJdgvV3f
P5qvCPqTzVCClcGJMI95k8KIQ5uNU4HyibtkaDxEmGGl1paXorfGWN/15dGT8GGx
PVVvsghOjy0ogs3mUacMjBQVseBp8yYfPcZrla6c40upbObBJuJ8qBfJ/MhlzV7U
i6LWK6WDVOs2mlkocTa7sZ0wbq1CP8LxENkFYdEjk4CNg/9smF7JAZKN9xL4tNki
b/yBkki3wwBkc+fJ/4mreLUZY+YUc9mnJRWYSVV5GWZE415tmAGYwdyue29RY3DP
5IIC+Pu6KHsIy1z4Thakftdr/4sDSTlTfJHzXoZVs88MsFdnqOOXlsDgpR+AyEpm
JCgGFHrfTudBK9Kax4IwfAfszIieeiuWjKUG3+mvKD0Wc5P4vy+/k6zbb23JnMXC
QoY4Y23rLnJWknsJr2RJdMNxx8ObqQ/Ab4NDjS63URAJhinZ2DWq4qtfrQWIn2a/
oLkAGXMZsjuQ2v2t1xWjTtLPUFQw8D+V2NYLrP/2kzJbcznhymKPKa7j/iHh8pMj
hcNQT9Mgt9GoDyO8M+OuIn4OXR9t74OninaByBxuJXpI9P+AMGVuf4UeX2b6+NvM
GsQRPhUzRzcvPyuxfgAqLgumeBEVt1YQ1c4PM5+bZnWMZvo9hjjvaOCvPr5PfM9b
WMORd9NWdhjsl4nXiDITX5fZaAWkMD13RobEmpX9L3fq+gmwO5fjTPBDK5ovERSD
ZTMe1Vr7/+xPEfpqlSnxT8OMcmnZIVE2FVkcjzIW2gCG/+gThDLMy6R/hiU/MRTH
ZYps/rtOlp9LR/xq7X+yFzNCCCLjsQzdxGhe4f3HBJ5fOEGXqRouiO/9pShsc7WR
LNtiXfOJnr27AmjRAovVl/5sp4Ec6VKVfw39r34Bd4a804FaTEco9Hzuctl5y+Y4
ZlKanjQSEXdxIVxlNJPiUBAIw5OPJLvM6sjt+Ns8UVmtnY+IlQJ+4g8zKem3pEU1
6rc1ML320cTq7hWrwNsFyjzkDjHLUEbFq31mfNm8oiH1BV6hSz0BcX9JoScSqMLU
rAHv9LRTO5ktbj4LkGcZOLj1Bd8FDTSPn6voFUWXrotvhNiUpzzAax8B7dEl9TCJ
rXK7iDeZsrPBmDV/61IHW2TMIrvVrCquXwM+j7SL7I1CmdFfJUm25OgjPn3N/z5w
ZKWrwn4TO+XjHKRgc2mph07RnGg/BZA/MEEcXIaf22oi4ktMe+o858/PFWOY8O6D
HJ9hj3PxrliQH80JzVOGjAgS1WZzheoqW/4j8ZFuiC8QO6hX6/owpmdMAaGmFp4g
WGr60eLfMk08EH1PjMdWbrjpdIWYwl2E/csSVSZCKbLWLQ3HGTyWwQGKob9BKZWY
ytDVdT4SWHOA4x6jsvQdoS5hzDNY17j3X4eKPoiHkUOSpbdSqGunG9Cogf9z7S23
fC2E6Xzl9Sc2+geibNTQIuDdgHkOIOzPJzdjSc7E8mx6vHbEAD6KxDqvz+d00VF5
SdKmh/D8PtW+tAIOPwQ3Dv1DqbMfkqmhbps+X+zVCff2R+cphs81lK3w+oWs5Em5
gb42EQSrLq45g440ds3duVX46KB6zNo2dRWn7xH7rnAOTwmsgSetjvHVzQJnZR8M
jWpw1hAf+bfPM1+QzOCgz5CnKsqlco5eCVPGeGa1E8PijmW+FctG8K+SM/WQtp80
JXTXXlasTubrDngnoiMi1EB7IqpHgstgjtIa00JS6L9U3+LyJM9VapuQptsfhdhx
n3q2OvwHnl4KlctW4XrRaxxZQ/saUHivH+9co1AV05h/+h/X+zsPxW5id7taNZNb
TU9K3BzUpltBjoNWg+5t0l6WzhDmL4HnnETKBxshYQXs6z0vPSfml++3PQ9f2KCu
Jg5leqbjQrIpBw2skwDcRsvUeQfQJZs4cCwHiU+XvfBKDkFfE+/53GBSd/fkkjON
MZeL64mCrmO2WnRMG6kEiutf4oVIeKHwfIpbmSS8om9c54lNndUGIiwFxDsx6Ez4
CMgMOxrDSgcXFvy3TvXwh9DoPU05loEGNaX4Uek9/U3a4XZKiP46yz0PfGMDHoEc
ShjLbM1c0Li1dNQDkAjefq2uImv2QnQe5bBiRfO4BvFTbVWeT6R1YEipr8+ZYAoP
BAabRLSmf+RtTJ265+OqFTrjgO44mEY7Z9xn9SR9Kyn4rIo35pPOoVz9EKiSxvzN
r1kXHHWkVW9iGDFlirl+aQdeM86/bDAQSbNQo8dHgkmiF89bZQq0CArwWRivUsrE
vFcowKLgI1wpz/LVbwoWvdXyX6CmrginxWpdWodtrRWJOvs20Dh83msqPb2iyVfl
YDS/RO57WkFd4DnvUoObQAC/ibgzlTdj8KN+92jFwjJ6/CqjqPbDLUvstymqi0RP
Y09CQibQ2T+WxhApd6abKURtZlTdE6ksrkiBuZ8NGKtsyyic9I+qcV3sh1a/sFcO
LSW7TuVDlhjwHampvms7wtDAwgI8mt/fkNVARfFpkdumtWThBcezbo7qd9Xd/1bb
lfFQs42Z6UJhqQsPOFy9ZEbFT37bpqJncbx7qWD6klHJohVNb+OmsbZIR7o7nAJS
tYsnGduqZzMgilV+vTelmkregj7rnfH6GCnn8oiHuetmupgSu5SVlpfGr74RmRG5
533GW65mmeM27DJBRlGn1DMd0kPERhjUFKe3Wslu7ei3DsgNVmO/qMb4sgtS9K84
EpxmV892IWpL/2imsXsANY6zq/wpK6NpAsmplqqpY39wTdK7KKzlJdZ/N+O7PFZH
ElG6Sh72q1lxW+cXAp5xm7iUdBeyLPdmDlW6TOOZbQmfSWmnmApZPC5w3yuJnC/P
AguDhh5Jm8OBYrkZ2Dm608ss9Ofx1IkjRPr0koctq+bxXDhPTZfo1Jl1eiRwGbyE
lKeq96YMN+91cx41BFHku+JVeu6z8LQUg+dul4Wm2uiEBVczs6xm0bHiltsjhxfJ
6AJQ5iOnke1Aw4B53RdPUTvipGHde7B3QqRkgb6ruFFuapvNpdDIUkcoyIWe2FZq
E1u3amMvX2Aa88OvTxB3d0SYHSZPKwkAPNZDjDRvJy6/o5X8Ve/6NzayVrMjlJbZ
Ykd9yQK9+UVG7TBwiZ/dl0KKPjXL4dSgD2Wd9uQVzJZ4LFGflZTOpZrfhgk6PBzz
gTfNl0DcTqcnKmXuLfo45X/p6ZB5KKVzFp6r8UdYDT8oyQauGeR+VGqPZBlmeY6p
41bQyAY8QfPx5u1jEW+mi3tQGEUsGt7wvqMPtI6kaN824iBiekrGj4lr8R/d8zvu
m/I8aRTfQyc+BAr7Ah4ITMjpoQD+WZAZCFCzk57bMndLR51Ls3Zix4Qs2NKcUpo4
SvSVToWd6n6exds6RzVxNI8QXbOw6XJ7uBe8shX/Lua+8/xypmcntIU+KlK9jVTD
PxUF00r/CL/VGxhZB8ecAcQr0b77KYdq6uE7Xi4AddrCrB8emc8d5SzEZ3eeI5Qx
zxbpLJg0kKhYf85dg08twwpNon9yz/+/VJk6KB6wInEx8dHY6V4HQJ/G0QDuIpp8
7HIvZPGSFmPbJi88X+RukhrYKywkJphBojw0YamSJNEK4QGMsLAkBGoNjeZI7O/L
/dYI78571L5f4bCOln81NNLkZnarnl9ehOXvsM9BCoRMluQsqGcs0S03U3Q8cRO1
cPb4M3lHKZJSVB6k7idQ+rXNh6PFFw1cHpmmaMZG8h2b8xt1SFAnTtEE6W9s9t51
DR7F99a2gTV+ii6GMMgQfxnh2xvM26U08QNsNrHEVgg09/2F1EdbNaASRzkniU8K
Y8buBXPoXpPxfwH1shv+vg1MiObeX9e6wFGcxS9EH7WCdeP4fqnCz36cqH7X5RQC
Gw4r6kAlg9474nywNY9s4mSKDppgwfADaMmkLtPDQ0A0u1FwLAf5gAqxACg/a9Ul
kNSRYMD5yeIBpxQRVDiSbWVeoas0cI3tJE/K0yX6gTJYFCA7SaV8PkMk34bG1SFy
6duQGsRMeY1cuMyecNA4Ng9yqwKB73Mc/5Chh4d/aCNAnUd15ptPygKLCRmM6cJH
nqrYeiQznqNmB9HKJ7ha2jLEtDfTpiI7VZ6GnOhyvQjXDKMmSFlruvM9KtP8HNGa
b/+pFWeXcvlrJFFoeVHAyvyKABQN2rEQwsqRNlZ3aYbQ1XJSttZyrXTY2uHKgcyS
j0KlBQI8xIN1CDrr80AcvIxcuvViI+hXGn85pdXsRj0nE2iGSEb4Mx7WE1yMks4c
7EsVxjXaTnNtpzL+XYMktgn0/IpJUVWpgDgCfQcbwJyY2ODkBo/GJLSo+m6fWp+f
mfOxE6ikccrG1KRFIbPGwhPgTG/OdZXQ6iHDv+NnMzShiptRROqUTe08Bfaz74ow
7InQgoN1AZYk4yzE7wlFalZhpWUDQlwsqk/XiZ6CVKIYLdC0Aux+zxfF3OQankey
SA1sK+aVv/o+19k77ojulADbTBAJmT5GKqBGR4bkSOibxIknKfO5YhQNK3+TjDcT
+Q6l9zl6UKKSAIgifeEcpZNDz5lJ36TmgVoHXg8j6KU6h+51edxIzSJBwcDwYj/M
n64HmEwWI1If/nLz4xugIFN3tUjvXozjd1olKve3qOdqZLtdobxhkM5xP1NsPgGN
W96hpydWD/g7NC3w5mN/8DX5eBVDyMnf4a0MqArkYGiq0k4luPvC8pVnmrq03jVu
CzO309/Jh6K/Y+qUjiiw4MwnIpL4ueWw7CfoFhoAVvxba7m7M4OvdtudFEg/VWfU
JrskympALbx9UO2gWXlLBbFIMi5jpMAE5Zh5600el79ui+8jEZIfaBHKvMuqtA9Q
UEq2HUKlvUwcfJl3J4tF+uXLggPKzM2RKOPjJauO1F1zZB21xYi9zvAFYGJdS+dn
q6BOoTds85Uoy6RQEZjOBBkmA+JY5LUo5d3YYK7A5b2v3jTl9iTriO9dBPBi1loG
FCEH3xCgPrRih0cZgauTWx7BOEUVs/0i8xcO9Q4gDdcpuT+i9aBr5OMuyohjb1im
URZ9+wdueKmRTRmur1vu9dK6vXb7pSkb92anZTiI0Mr1La6MeWYZcvGuuH6Ad48p
fc23Gc9jK0OExozGOIbJrdq/ZlSbLowIMC9xb/FYo3MgkT0/+2tzKQmrFqmhQL2p
Iy0okuNsH6pmBRpYTsb6LlqvSYGOlo1bM1G8SiuhaviJUQkdkJoaP0uk/mfwqqBj
zF5ZRR2oE8g0p/v4RMHv41gifROeoDMlkV2nZ4tiFc7nU9KhltCpbooagNZD+RTk
WVA9yygr+BnblwrEIUT8N8qetedOmDmIqprmgh8KTrHeRot8svZDMTcthhqU2add
AnucV1ZD5PJhOBk77VpXnz+Nw45ovNgLywDCe37tv/7IjCcnL7cponZJpA2ZwuO8
8y8g152wHkGHU80ayBUlPyQw4ZrgED49Unm2Ae/CrZj37qZMwkoBzh3xVI8dy1Ma
jI2auZ7GWUkseyS1ORdwYuvWtyTPGADngYj7odk+r0PfiqlEgDow8zRSrtN6P6ll
awWTxeJILu4osuDqnpnHFHcfP1iqsKksK+bFGECALAD3JXzbWnqJDf6wgAWNml29
8O1qzqW9xxnQucZbIXeqZidbmJ9yM+Y0ZzyTWo7bVafuyfq+klZft0hE/G6BlSny
s7Y4ZIRnaTZ6f4ZTsOx6vrUPPwmkB36h779Yz5MlJvBwLqiOnvv/dCbqXq4ctP1S
pbszV+wRHgfEyXhazYe+Vw2tEVnwTVzVABbHBe/8XgSpY9ll/8w6wSyIcNuogl70
/6PmO0actmGO3nCdJvuFGHD8IeXKD2RoCdVexZJeo2hSYI0G0bx0XabftAJcG0ZV
Gn65mnY4wUdaVmOHQzuznm7or+r55QNK+KbJsR8l0SbnhFNsCg1KZVmOJHphJJ2v
Myev5oLcZHbRcyD4Rc49bCE4m6fb+5WdSpNJ8AQoZr56K6qyuYhLFQK1bNGw4kdk
2FsSV8Qxk5/7PTWqCvEZSwCeUHFLcd5VU5ZhRJR+3a8MCThu0YXBsZfZYRrN2spo
eNMMmrABpLe/QxnsUe72dL37GJot9Zmmi5f5v/uCXRyhVMLxiCpv+R1YEyGziAYI
dy04dnMie7WldzoiMG3MujU+C/mWAbgdY7ji+eBdnIP4cgfsNeGv8Uq7ThTTkkQj
ggtg2sG4lkY8yVzNvw/cEGHyA4wgkhq2rfQEUA2kw6NlA+M0RaCWUrCscG3P1+h5
z8tFaXfdixADzUiI4OSTXI3yqmHvHaJiRg/fVll+wpw1K4Jtxhgio+NaouxjHGC/
FIUfdkcqgtIAghaN6RuCA3hFtPw/vY0dDOUcmDc55bsP4DZvQ5YyX3nSDE+m9Zld
Ad5sVwMTMOvCF+zzeK1GfgzgwrwrrR9RU/ACS3LVSfgBr5dFlgr+JrwG/ZhAzuGi
b2sq+q2MLwyVPb5epEQxTyrb5JCYSaUGaqLS+ZuZBoXu/tUUhV6SCJxxu8bnA7aN
vkp5e/i1LO4wf0bLbHSPj/WUtWiGo40bcKKKLHTO3RKjIKEXXM6evILZLWOtYsOH
SimJwHrXmrHCHG7yHrk4Xpc1O5Iy0ex4O0LAaulL0vcpskU36Pt1izamN+pPH6y6
AlUrZ6dpU2bgaPCJ+5DRQXIE3Q+qXjoryNUFqasft2Y2YcRDcDNfLsP4pX5Re8O3
mW2T5UoOg0PWAQgZhjjcJg1P4S5gqL2UeC4M+T/LiiRG7NlwHbXsNctiFAxuLXvm
4BGCwxcTQ8ZyHXzglw1vTO2IfMrQHkr2SJ+Y3zTFP+HQHGeGMHXCBHkVub2+sOuO
wjICZyKDGgLQ+y8aLD4ggni7SKqAs0OmVnSHu7Z+gEqvA1xIiT8He+erXEzltYUZ
bfK+s/9jYYNueWHTBoAGDea29JqcqX6RiMfXH+hPyuQYcg4wV3O690sEycC5pisJ
vq73Zlv2JDOXi2R4ZzNIl55Hk0X3asMRVhuIxbK3JtHjfKUuSflIDsyBuK8shg1C
LBWzR1a/xz7+FphZLAUxN34v6HObgiXLnnJoMdPvvjeuL1E4VdQLCTS9GryFY3xA
YkiC7iVFk6StgQoRpgT5JxfJh7ZegvdcWWiY55g56+y4Ozwwb2+esxVNgXdvuYQq
8Qof+PMfi1RAFUuv1p2KFjBlgYDLZr81WdxAROhVfsL4S44lHzmlsxqQB7yYErOr
NDU8+i9VXf3NnOFm4nXHrU83r9PqZ4wpg6MXWgLh3jpAJuBz+ZaEvlNYB5+LYp9e
ZLO5ymad3YkjQn/3SxeCpUNaLbeSt/uFjYwocogn6uUgq7ZFwF2tk4+cgrfFRYlH
VxMErQG6gkk8H3+Bf2dWS+JYmT5XRVVnm8fDwUlD4tnr79Vc+0+hH0M5MXUxvE19
fQrSQtth/TzJZoJRtX7PDvzmJEt/fr1raC48G2p362aHadpEpqMqYVIX0E+8g/h6
6DQWE00s1nLEK6w775DIit4fhpNBOSdd74hbqfata+9d1Qtg+h9d7Uu4PYShmYlq
EnhaPBWQQXIIlIF6LUMyzLQREOYfTvu15K3bs3ZuG7H5J691EoLttPADf5Ju7DGc
DQmL+o6naT7bQdriz+TJCnQIifydvdGyG9VcMH6XAM3//EvFLjXvabiGqvPkc6Nz
7EBcF8RkTiXxTrWPvVROxIUgkKeZ9HLB+CRMMqgKr4HS0OE3Ca4uzG1roIRbCfma
TNzK7Pq4mso1Grs6H/VZLrDwpWsxGsaJDI4D/5GaofcEqCaKtdrxPvmzLfw1cIUi
0by2Em3EAnq0+BbwXWeKaqwuwPaKdza+1tIsUMhvaHiJVJYKyedqjS7ZSJsnOzln
1FKRm4d/Lm80QlTae1tjIwybxrd9uGAkyKAYWdtAS1IXPV2RBViBa7U4VAKG1WZ6
sy0JdNVn5W3kxCqgrTAiWTu1SxW/61TIud88c5W5FYdZIvx07YeQFjb8SZDdUD/P
Alhf5vvBfbJVF5mOFSOdEgURkLZCWYZvzLJxer5rtUC6N9Y4eitEIElcLEQN9iyp
TdCaOacyZ873nHYrpPKMxyLpwGGPTw2qcC0mHgCnk+rp81bTjD2Qa3NVaurui3OZ
60DJf3wAy2P5ab/lh9y6dVTbKMzYBiRyBoJqyebZE13elFZBJhyzvs02LWWShGW7
DR41wtHLGuN2uTkQfJyZMslN3ZZRnsxsDmiR628U8YbqIh2jizJB4WC8TRmWJbKu
GPk66Gaw5b1H+rM8V3XJhbblb1cD7AoHBYj50h5h3LNKR0wsXJAV7bhdxF6iGEC6
qFu52LGhz3rKQ7wtz80TbzOeQOR5hK4OybGtyNIZQ9ayb+jkD1ha9aTC0+0nhuYt
mx8WalkwElsixSwurth08Ucxs0zbhmV2TXCWRU8OTiKCDeH9CQJY5rDBCEGGxOYa
nqrR7/qPwSVZBUoljMDR1o9OgNuu4a5ow2KIUxb4SAk+A0jIC/OIGCYH4NRFMi4+
fLGvy0cReyMsMpaTTTuWqojnxJO5w85G57Zm8zfuTxXy+/PhT1t3DzD/eAVBFuZH
`pragma protect end_protected
