// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fa6epcKHGlFZVbxh7mg9OZ5qhRO58199TLYlTbBgxCq3eCTTlb9MJtnyzM5XGXoX
VSDahKe1hqYzu6ssuuvPUXgm2PjKb5Fz+go66MKZESMBAGhnjNxDQUAkt/RbI960
BEL6tm/mNq9wn48W7BrFlwVZFXJ10QLAO7PDRgnBxQg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7104)
xHwivIIP9CY71o+qy/kzbArXbXlO2GOZleSfD9T3hWA6lhlnMzV/Dg95Vc75dezA
/AY+JCJLMqN2iTxcvMHMYok8/U/zsHj09pKlODGTOZxsL9eR6ORzXkpDaCf+F1JG
zaUYNftU7pBcIL/8gMknCrNKGyLjYrLc1ZfTLlfT3U6SWpUG5b9Mh7VHkUEZO/vx
gFC9VK9x7Am/JExyzvoC1oOLMjO/2dLJaXyXnt4C4O02BGGDTQj3beGGlkVGSJvn
8uPQ1ISuF6Fm1BkA+rBmDeNFemqIuoEmQzoKhjUbPlbBYGF3w+xdbHLySJg3H1EW
gpXP0oPvn+ug5IQh5HJdpyX7dtxirOyZ2ouKw7reJGPWYutwq2Q56n8bkACqP8yI
LbUo/DvoyDZ+VMZ7OKi8TH6M48EWixjg1ZFVPocY6p0ME8dhdPd9PuWWXm2YwW7V
Hx8HvWF2BPu3Ux1GIg6AbyE/kxSUaUpDOi8vkPp8238cpWmjtrsYeON7GwJsv/Wf
jCbzqeTO1Vpv26x17TYeEwRO3DR6Nlux12nuDScDVxtNhxSN4Glk4xaaNb5O5RFW
YE9I7sRmaKqDU1CcwGuuf1vOFKHkKW5bshMRRIp0x155QjNRlQUMg3Feng7zZzrs
Wcv+P41LSIXGE1nPn13DGeoR/kH288dSY91Fcn7uysg5ZAmFdLkErUgJ9uBGHkqN
PFraspggs56M4V1rCZ46DW68RxTYtz2cvGWAPiZ3sv/Pg8Duv5W5jGzl9N3KMPJ+
XVWFTGYFaRnDKPCW0VaKOtcG9ozoUI3vb4KxjiTAeBh+C2hoGjWPu74jy59iaYP9
fPxDkGVAjtSgIIaElFg312Uafx/WoMVwQYsQ5HAfC7lKs3R85ap+NEcnAQ1dB5PU
gZtA44OqKlqsiGBfCYAu0S5YXymrylqbntCUetc7tlye3w+qmXypewaAeeU/wMlj
BUcvHJhNnKLW9eFfme8ZpRprKl7pNKBb/IJy8qx2ojUf3jJyaWiSmQeuLzC55K0B
j4EAqVe/O44MF0ntH8NBlG/9yrAqwValsL7IS1Im1Mo01CsfJFpJBrKtqcdEJb35
bYyselYuZ/ZoGeGnZ+uTUBsEdB74nJQm4ajW9LMHjzXTeCrmaDlM4UWW7hkKx9v0
JvL7Xag72xR7ahKl6XCKfczN87SyscoXKqz6RG4twwIQSqNIeYLdN/5bz+o//Anw
N2Ab72WfMIoQy27zVP+b2kDkFSqHJSc49aoS2rtH5UwhUX/bEl8j6XEGcN6B55r8
d56PyQS2Wd1hrCTiaNo47aERwqNygC2Zia/J2DVSIkfGnZhceK+WhovyO96M5cVQ
O/auf0/NkfnIYMXtvDsgdlL4RbycXTdPTVXMtaKwCMoAaAn6WLwTsSV7XxNs6AhZ
P9YrzkTrPyxEwyR8pNkcMeHLE7sAQ4qFw/ojZTCl/rYUl8njVOk1nbwri/4UaNvG
gLW9I0d223l4gJhJ5/8fRu1zuKO1wZgS5aZFCav3arAOMW6G8xcCYPJhoLE1Nr5E
9M7SD66wK9u7FSv9vI2UnlK44a17qUNT+dnKTouFpgsIw3deIEI5RVqmEs8dYH2R
Fsw6t9clE8Z7JobNXMvlnByIyAsN8iIZGK1EQPGuBn1oRPifiLXcGbfCvLKccH/4
UshuXCqb/EgIMSxBnLDFRnhbbcUAXtnDcUX1SOao+5KxQDBBGWRg7o2u36ht4xak
m77GW6YaoOfkW+WDa6Qz5qd3/FqMARt9yKjlg4wfZZEPUPniHTDt6IU7Bx0aUQqR
6Li1TEmDbKkdexqtiCd4EMc8xm/sqh17fwbNXg08nAni5/y+Y7iKc1QJrO9mRsMo
Fkxxh2ofNdIzEQl9LybLj9fe46f+c22Ds02DfLZlKDLOTNjeykdMtfC1sUiT8p/S
5PLQR160HZtKFQGhu+8fYaOXn+sJS/36Hq3jT/NLYKUFNA48NRUUfbOTICItcmm4
q8oh4zJcNf7z0MT1ji1MkLgKBI+zM6X5ppJI+Ri9pHrdl50vfeoSKsStZPmcy+uB
p1u/KnE08uAsaGVbWhH8MXbVAu1wGeBOPoIO+Umtfi9gnLgTBaHUx6TTdEF7b76m
VKNWJUI8Y+QgSbOPzYst5IXlhmudWEM+FaeB3Ws68F0ifhiTSrqP61XXrs7UFG7Y
HvFAIOsISgIYqXB2GjqAVOb/X/EAVUafZ0k1Gi1mgLZ4+jXCaUkocbMbMOTA1ZD8
qzTpQgbR7IgHpTRyWi95A5AvJBOel2mI8NAiqEQzx+cb6xQVCWty/Bd35RAljPfn
pAVed+i8uqqdsK96KVPORwNQic38IvB5xIS16q3oteC8NYh8U1xAICWZilYh3RYf
9kpbLvmkV35epGhd0HzOq1Tswjp3bgqtW7j3hiUf7EQOzRsPa/Kwg4iM/rNrJeWp
Zl6OsXPM/CYDri7oyEty0wDfJZhRANUWkE6edPVTAAQVPiqL1RU7+CEQUzHIlEne
K+yQKzpTXoM3XISf0OG1ScTnwH9DZPQWjebz8GfEbEEf4jCfHtKk03uyIcVFppy6
JsvmdN4ns9gVzReePFznxPUnM5hjYxShu1zpBNox+xD4A9BdEgF235Yd7HvgpD4w
ydRVhJA/bzzderr6v4sud1ohS/umcWwcoI87nJLv68GNOSFZ0a2F72Unnfbb99kN
YhT56dkyOxC73ZfMDHlfq4FCa1QUgy9Iif5/CxETn0ghxZRJzv4hr4im0tRT5n9N
Sc9cSrCkTh73Q2QylkZFmDK1BXet3bSjbWhkUMLTD6nRDW2GBHMpLBsxAdNjxpcJ
V570g1t9qUWbrz4oanaNXNtVKCnq9KdGLu8MqAYbptmmBb1qfGzKIV1te82ul91g
VCLbC8PGdmIFIDJXja6cIPI9R9vMHUPXFXk0CnORqxbdunfPCu8gwo2mNNgm5diz
jUJy9F/Qp6JUhPzoG8GqfiO2HTtqrf4Ry387HM2SXP3C3XEMqwoGilBzJCWubuWm
3iSBGKKDPbs5X5iM0nKH8r441oZBuk11Gp9PCeQYm0eI5xLNMZtUZIrpyrq2OSTr
/4XjZn8rXHZC7i49zXSWRY7jTvm/QV9ciOSUUc2/U1geFHoKaGoLljmgNjtMC6Bk
xZkgFCCrBYd4+ZHmKa9yJ7F0cCtZp/D3TM1ruJvE9upCiA68qexscXfRQruDGRHH
IjXK7b2JK/jbo5JuUJpY6SHXjrv0M/gKaJFovXL1N2U3F54cd/Hi2K2PfSThAH55
Bq4A/Ku1PHwlOjU70ShhOTCola1Aqjhu4zAjxQJFow8Yq9+I50q7OA0SOJA25C27
sRt7M5AQHWfEWRaI3PC7qSlLmlY9zb4u58tCFNFVezst3djgRm4ElNxIi+yC6deS
x+K1TEwDKlQOYvYitAKyPAgNcbEIYYC7Qo664sd21yajOZtrYsdxRahGBkb1qaTk
WEEpRp4yP1fRG2fxatuMrk7IJjbhc5D6b0Ix3fE1erTOBoYdL6f9NtIxPbm59zKM
fpdg3yk3soC6EKL30noSpGQ/7tjb2PyX6gaeB5uc8l4tjFSCiVcC4x8MHqBR3NdV
RClkz7+A9LlMjlhYkPGIFwvxyVLXUzkiYAnpD0ICCTWO3w1Zs+4HRE3wZSILtn0V
wlmX4fmWQ82P+kjf4aWvpns8GMupK4heTnMjx8KEDeisJlytTaz3kkH/rd4KTabl
skXUYDwqBrAy2NmW+NWxjdrCEzMXFjYyTIhunLHmqsaX3dK6ynWc5eeEy1erYFZB
23G3DBzOF2rmYvsuW/oKgHpz+savPnrZTl33h7GvdJkakgsYDFw51b2HVrqxEKyh
3V6T/1pOvjcHQMZ3vViMD3LPbTpRhKIlfkOXnBNCVEqsH6BRl3GKAkuSCk1tatq3
9xozlhTVHtYjv9wd00wXWvS5DN54T7sSZcvfKDLcgue0lvWGTNgvBjFz/JafhJFW
M295SLwVh9ryilop0fmpp7p0os+E9BruVlkWlh3d7+F5yKvNu+cmXay2Amvfi8NO
CfQxSNDTTqo6PSZt9ZmJH5IUZC89uQJ1FXsIvRaZq3+lNNtivzgeeDof79yPVtEy
cG+tfPVqUqVdjzya7zlQLgAqKKgYUM6WEBKC6X469Uec5tdRDjsnE78hW4JtCVuK
gxo2z9j470zdGiC9KPGJM8GhrWuh5zHBSOjZgtzSfqnOgGk0s17NCU3LsYfHOg2V
6EVphgZI6W/8Q/qZ/LRt1wQjkAK2yxMPlvdZ3YXuKqUZ9AFxICUy/Y/39QMiU3oV
cnU3AmHOP1kwE01qdszJ1xZ4ej4O7mJhNRpilsGffmi4qUgG45mO1vVjM0eSlpYp
//CxsK2yOA/hhDhJwT7zVcdRHrIA0gjbfPc4/SHsf5lFrnP7V7y4fr4E4Z+PLXUG
kmuyBbT6kiGn0UgXacE0ZyTzEX5F4ddOTFB6nSaTM3OzvWDMT9VUvu2p4pP0LTa9
5Kr0SWwKVZTLxWeKC4lD8a9+dNVq6HSr4v77k1fLWDPHlbq6jkMnKe9ErkeXx5WK
Z7llC+8wCfx8FcsVq1fFUuBTjQ6x/z0W4qwXflkUrSRwvmlpE7esZ3lNwiyizdbS
xuY8fo95qOHVYA81GIrs49IJUgkj2xiJO7hUKCay8Y5FraA4+ubir0A7c8R6Wg14
d2fi5CcRTYpz0xZO1F5hpRtbcNS0AsIEdRPZfX9FX2lMsTVs7SrlqAZkIt47YV8X
CTgxuqFD5zQNpT3DkfEgfJ7eUp1VpDP2Erj13O7rcLpm7jFpAA2d8UjmTCO/z2V9
S8QZg5xudLpNtyvH0DepaPG+Z9R1YaCD6/pAe/imZwgAGfQiQyIV3DZ3nWaR+Zmt
mr/l1I04TMWyYRID70/z0EWPvMvpD0To3cYCYwpNSlLOtYnYNFdVOf7G/+X0zk4o
VhTWUeeIrcBDEejbkCJL0DasAMW2O/V/quOHZLBVPQzIOY/y+06GdiNHLGc2j5gJ
6qT6gdQQxmK0ubh3xEFjIX6NS7NTavhidjCaW3rWgsOiManp1sZGXV0n/TjxBD9s
1GCdIcb52oeZr4TDuODsdBoX90jaW0o5hXvwxr3CZv7vewHogpbd2G3G+2WBSeDh
MmDDh8BP56MFx8XsVCNG0WotVbvUamdwAHZfkFv4BfKTdUx/OtnQVqDqDy87VdKq
FXrNkgsM5swCdAiVgurjl4mBPnE05ku37MQIfNw4126Wztkt2sqpP3esE2zru3ZJ
tedA0O27D/voTf+V8PUTQgGJ+QAEGZr+xNTYefdhIQgz5YxayOKBMOYHsJ738FWq
eFM4/q8L6oh+OddFoxez5iQYRPlvNpMuEQVaKrzTsUHh8xVCBwl9a6Xd8qoTDpG+
ECkCkuosiZizMoqeDaKqvjnpykFjTB4h6Q0svQWAykN+T5gLfRXZCI8wKsxahkKJ
8nx7MA639BProkp4OGEPLE+1BBT1hhp86Z5BtssB/0Dq5XxlOQvm6V9shS43xjoE
dhkyH+L3V3sK1SWSUPUs63WRUFs5cZDRvsj3YRq+dPcmTfp51G7fRIqbSVZgrx/i
9X4bvJlQzt3dyku84wbbzvy84FktilVjzQS3PefwmVb5ispKiRd1yOPiHT0qqWie
fRHnbGlZvTA+3hEv7jJSH3UH4BJYwHRtYAd7466CEMx3ZxxsdR8QCMQ7KG1hO73i
JNftVxrSQ7QmzXUVA4wMVKiw+sNT8/c1R312Jwf167EdrpJ3NCkesHgclRjLjzmp
0gsocI8xgWOIF6lkm71ucoM/aEF7HllpMz3YCR/U12ZGD8aUdmA/l0gcdYD/rUYf
XN0JEkesrhJf49Snj+mG4lFClacXvM5nwTCjQS/UXb6xm9THJ1d5ms1eoR7IXqhn
2VTn2LFr25wCKhOHod9UxSbTTD40J+zKMzTgqtlpvPxYdOFotE7WdOHpnphvLZ8/
3oNZeIXijLUEZRN/tyF/pk/JUG/1yv6HcGn+f6k26GpIIHAe/Iiw0w4Kx4LtG+9j
4q93vUL1BO7r+OMKDlJfa06IntqJbMIb7n6shcKPw1fKF5FEQ7WpLtn0GDoMeWPR
Qotpa/pYtq1LyTx3j4Ozv5igGRKmJYts2P9ZL3yBkdHu4PE0t/wF4DCWyQFV1EHD
LPxn8ZIc9PnsJA3bDBAVkfIdFnNq5TB9uuNqat+CpR+kWlbRaJtVPMI1RvwkIcRj
eW8oLzuJPeedEuegmhLi8yYT/xDDE0xh93jGqB9KYd/kH5H783Omg5QTFK7M7XgJ
JUUnW8bWPcqnZiTE1/6nAPp3/anwF0+nICWmE7fW1/tSGRLDPH4bpaYaIbzB/6Nj
WeknPt8GxRmYuqi++ixwWHi2mhfyEHCoDau0AXfwPDuZhB9cU5xvzJjgJA4PMrQQ
pt/2scTCSIzO5nYAdjfMNU60rFRKBiUWBfo66pQjEuKUPTzSjZtQARuvoKOhaUl2
890XHiriT0KCX9boJVFaPIm024nHPpI5o4BtVhn2axPVFVVoxqSwKke3dGOt++f3
p/AP3VwahRi8SIbc0u8pJDyOmMLB4VbsLEp8tLDG+gCae206FLp4ggpHb7uMzjPt
+e+jhN1SDc9pM2IAq8q1F/QIJgxNBvA4iwwniKr7xoEcrykwGE6jB71jH8+OhsvK
jJoSCTn8N9FRbKfJLEUy/6nfV4oeQ3An98j5ZkyAmhnX+XtN4zzgebSjC2eeh/A4
5Z9TZbja0oLILHwfdc8ZafSLMc+q8b3lGkUFu0syDO0ja+xbLYdUCtV1Wzr4yOnh
UA+9GApiQuMBp3Udgq6kJLpmgCL8pnH3yNnvS7t5JRl1NaE3FmhE/GMrZjU5zFbi
cjqtAku0rZYZm8yMJgPiNH3oC2SjXeYPF2t8JYT/WIxiL4ui6xJ24ouHpDxNe3z5
pqH8bXnV5+X1ci4uTqeX8J2WvibgdFjdy6iDLxT6SDEtg4TmM1hp42/iux+IEwFA
cWbi7r7EDLdYlCxNjkUFTYi/t68vMEwk+AjhrrJFvnl2Sbn4nq7lQTPvrzpepnEM
e/Ci8Jpyf/G0fS9ysYfTo9W6fzlqgWNLPS1RECDbfmkHeOtsxigP+5mVkjeAGxbT
kEsGqb9ccLDMx3aPO1UQE5YBWYywN7C3kLtoHHeavMDyE1pnQctMxtr5Waagq+36
UsPSmkPJY4JKt63MK1NOi8PnDGKhLaW6Gfg70jiSvfqa05d8shXVTCOZdea6uroF
xyl2LmSmd7v8sfxaac8L/MEr97w5I6keSBR4YzyhnwegcqE02s6s9iQ0dWtGJzTB
WGNjm8ftlgiX/5/XTMZwsQgoFsBeibrSOcVHEMQdMETJR9LTV4DqbYyjXIpCJcCl
SAhkWnsN8RHxveJo3JMusiY/xAd/8zVVEdxJsD/H9KGLB20lBoeBwODiUKNMRyYU
OmIX9TgnLUnM/2TKPKP0kHqHRnRbVwr/X97mF2jMkUlGUk+3BHJ7RP2h6XnEtXbP
KrZuU+cCJqxGa4sB5VY46/WXsG5PRXP+wDDkogFIOqq1OvITkVyfmplfQ6dzLlLg
u4wD9exxNYgryC+pw0FvcJHY1woZxYc4ZS1NkHVVfgi5S9FUllIOys/as41eXH+R
Mqbzlp/ED9KaJ5Wt8+pJV2Hs6FLAw4cBPe0i3XTjGMmchF1LK4HJZHv454W1kMAv
pVk3ZM0fZNXl4xsHjwqjb/zwxxa0Zi9l5dgXQbFDmsJQYrxBSz/56vIcbQjwvCgs
Muh6WOYqcvLh9H8YO697sgHuEkcKckmV2nSnPJTkYQrWG/eO+3LWzKDo7GAr/FxC
LLdK5qtCp11MSVBQm5FzFPKfpJgEEkzNPcxqDlCDcqjc8keOwZ9qFRELFe/2iW+i
ia7YVbr0w3VmRqF4eJn/O8ErTRXmsbXTKWEPXHouFh4rsPiuO8knujcXLWWeQrw4
Pvt+ilIGXch9sThOmVsIRFvH4eUhlix9PijF3mMQx1fmhBQMZQlguKy3LddLHgJ+
kaQL0Qsk6SR2k0xJpHfUYy1oPfM6VSsYlQ7w4RYYHEzNaqKxkslUJU56H3M75XmM
4sdQCtb6LdTFUKAiMTq4uVbKwVoxWw/4xK+v1YMuKt8Q+6LnDW4CmCmpc4iS91D8
PZHwL4ptSUldXlpkIWpuW5pcoHi27UnqorKRkl62x+oKWD6TXlRSwDVlCTQ2EHaQ
c5UqJGIyGvP1b/+6ZKBw8LmeH42WwRcd5360AnE2+hgs/T/oku1NZqRlf/vp3YgZ
sF/IvPWIacCm8rRJxWUiTwmCuoPdBSfev6hmKM/P9pxEz/wxYqglENw9i1JhFbNY
ftdNko3TlC/FgLWiW2hcA4uZbygK3PbHB7tYdyyv1UR0ajI2TOHJ35ZGCGFMOXy7
E+9V9zd9fswy5YkAheu9xTYezEkqmNmnmSChge4bfZjX8o7kaEFOMHar4suFW0vZ
IYXN7M6Zm6deurFrbvSaFEv+f7kZBGkGsO+Lh3Ur255jUypT+WeOL9g3XajeBQ7b
LFaWmWhWvjRuZrwuctRnt1yezd7a0Dc8QVzfI7wvNU7NTnbrG+M82Oiw7AfKgPbR
HybQj+2jrQPgRxtt0qLUC0e9rW+YZbzgF/CMmuYmbH+P8h7eBjrCYB8ULD2a3k34
YdtSw65CMsKCv5JgtYahAUBYvLWKJ8LlZw5KKbomwFy8ZQsJGWB/tSqWXEWyWqI+
b2PMOgzn3tITB/vfD1fHeFsDSMA513xUVfwg68rFZaRY7HXlDG74gsqlrP/gU4sW
ub8h1LIFwq1GPuooqgwtEtk9aL4UXakNdaXpn1RKW0oidBjJ12DI668deb+OWt96
D29h1rYcCxTFLsLeQF5NtB/0aXVNnb6ehZuJFskwzx7OgmJ+RaMVN7MGl82up888
Auhysr8SQVfEQ0bYV4TClfkW2wzKb7F/GGIU0I/kRpZezkZYHzQQ230hc2fGkDLF
/PPuo9ZR/pLUpLPSCae9kkDvbpozVIQI9qW0oW7JrMwU92Qh96G8WmO3utqDn46r
UwFl+RNrjVtH4YcbR92nuHNz9JVr5FBaSpETnshHXnHc6mFrQaqUNUYGvRfF1SJv
EVIlzi7LJeqoCP+k8Q223uzj3IPGBnM/jOcypHEm+xEuywps5aZCVsnpdMwYrgsQ
XVVU30YR2KtOGCMb94CxUgMStN31iSF3si3RCAwX0l7b2QRfJ6J3pRXQKp2edDWx
KnL3PfGVj8dr7Xz9pR702s1m5bjjNXgtUXRKObfvn72JNBBsSqgO76iPaMeybHiB
KnQhmEUeyuAeTVsF1sogid0IJkT9ifp+Md4inKvdamuKfgfwyD9YB/5ve0d1PRdF
aH5b53fEez6arbmWrTN9nVV4uEx4axcY+4rLDTE6caT9ck6JfPvxSLFePP3DNTKG
QPU8+VaoLe37adfzOuua8WCS5VSNTM+Lt5iz+dipW7g8sM8kisDpdpppifZeMeQv
`pragma protect end_protected
