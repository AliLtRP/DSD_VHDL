// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XLsOjAJvlhoGorkydQoCN+oyI8SsSaPrgXT8XjdikI4NpaGNustmEJf8e6R4CGHx
Jmh+/JrnzIUheY73nZD0LhvCzgEByN+mgbpf6rFv7rXSvHfF2Cf7UYcVRrvg4YPX
V9nWDj+3YHVBDfRk7m0Lqg3adKFxl3HmIXDJK1FieCM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3296)
qkVzm9NdWV7mehrOj4P3pp7Zvqea95Zz7+4WWBzKCyTNjUR9qcCHI+Yjwiv/Ykie
uKr1UZr/JzLNLUiWaWn2qdjPMB8L9d/cfLYJyfcQTEd2hbepzPnRQgXEQJVUsEC1
mIC+5xMm6kjJjmuO9eVSXUn6ti82OvhZkNZDkbdiUPu6JpWJXe59Itarb0CDX0H0
VdLsGszvhD0f8SoNX5j3JJpmYi5uKngcx/ZtHWWhdyrqBscrl7pHpqrwf7FmEv9Z
aqMfJi1tAoAclFPSVQDS+evdv4G5EsJdGJ68xAvVJe8ZnGO7qdIRceWhn9Qlb+iE
e0LqEbvWtjFrfn/oPKNLDvD2P1J7M0pTf0O7+RmiYQbdGJ3K8p5coaN+8c+Qe1XZ
Jie1DsoJL/F/Wh9Ij76Jnhh9g7is8Cl3Zx7p8PnY526VgZLz9McIl1XGNPv9ergW
CpxhGNL3lVmc2Ed8yDt0KD61AobHbRH9v7bDtt4lvmEvq0ZfWkprzosH739nZz9I
vuOKWoRNruxm9ozEgx+Sz74/R8YKMF0j5bNw+HrEV1iUnIUJg9LhknoWo0CMSXIu
PIfqvgpbOq9z6REKBL/GJBsLo10ioGzZaVJDPVhXpu1FA0oipsH7w95edCDnGwSW
wFHUD572YR+dg4sVCw2BGuN/tqMEIC4qCpA3AEKJglUvaIE0dJwzbXHKmo5Ujb5U
BadctRw9qybDxcNLvogXjYH3vytDNrmJBLBaD4mK4Bt6oz4BDI7yCR13CXavq8wT
AUtS2CwleF3m+57wx1R4JE//H3A/y4eo43t2ftpIexCmAbPR7wcyUYlY6uJfzb8V
jWXXaL/jQ4KDSKcBk6N9w4lp1OdfxhVx2qbRkNaJW5rRcLnqN7PmqWKScN1izBlg
RIbURNU2yaEOKZ3OTNsi3DZSyoEIAMrizLLGt1G4M24SI19EhLanjc+laGzurFlf
CLmpx2PSi0xUY8NGoHhbYiRxTykNKj2i5pHRMsj7Khy+ACB3DQWnOrqFQ27S2TRd
nHcQqlF4bWJFy8CgdwKZq+bNCBHbPSL/glIfBZE/DgRYInNcPYQe/+JHd3OnB0WN
kizCm6sMmtJJROL1aCNKJCF6ZbGEi1CPRNUGPZwP6FQ2Jawxdx+JGBAtZkejffCm
ZBB+KF0niBXZj3cC0WJ0f0JLQ9y2iIH814NFWGanFM8HHlzu9CXyqF7vryHlJ3ex
d0EPlPg2OfgiHsig0SzNAGfV1m3HDBtVdKbSv+fsbRmpzIaaUy4z9e6p67aoOsjQ
j94lh8FiKKONErHYxNFBEE8bS4FnyEr9uDZZvHR7foJ1TX6REswX8yqAMSQrn49y
4hYQ+2GU7fBhZOgjDPV14OnXfcnSl6gA8YfrXqe90h856VfpaGbZ7F505x7TKa9N
JrJcKHg2Tcj+QmDVK/HR+20eKzenqDMPJhvZz7so95fVXtEphoLMpBy4uzgzO82l
dfUp3Kn3rUhhpZv0AncOmsD0Wfc1aEsrR9oflBhm71UI6aZOZgItWPG+hHFDtNVT
pP+wZvaeDjNR5jgO4Cd29lH0EZLTCoLDFhplZN/P5+/NIvqUrjBmigEHDar4HtWh
SBfeQCl9PD2EkCQrWpt0eMojVcxXRnE06Ey+J/aN+XxVyISyamQlCBuiuWZLVjnJ
4Xit41+CsYXTX08LQ/Wq+b5+/RTQtRuZHVNrryO4ZlULYNX3YDOSvStw6Xwy8Nm6
7kLNg0WcCDPfOj5jkaAyjs7Tf0rWBjCFWNAA9DGcTeaupzWtKKICf7RCDEvei6hX
CYABZlxZUlO59iHcug9ThQdtYcEzgvP60zpJJQokjTt1YLUyvjdIs4Ifu0JaQpMb
0iarUDjDayDiU/XkNTExZrycZg2Ys1pz67+mws+7yj0Y3SRbPcSq2eXFpAoSX1OS
PrBRVcGqkL/DerNcw1xc1PQlcTB5TpqV2uo2GaccXZYvEV1XPQMpN22W8wXgTERq
V6MKINDugWoD+hQhgzthHMB76B43olgNpOzDa0bgkehgu6kzmWVj43je1r3ecd+x
CVbM4zGIgS8GlA4Wp3K+QkriF2XGOGjSikH925GR9C/IHze1mFIGRHqOGOP6GdFJ
bzb8aX5vpCJ2rwwIKpCnNViVoPCzFZjiBwGDk0NqGwzhVRsfYzLsjtLMontxwnEr
lh5QvTV4yWLQsF8ucBjErSFjl4g8isXmMq4/dVSKei5no5rHkbIiTYPdXbWm5RHd
EgckirqmZZviCMgQVIdbMlu5GOTxhFxx9lzzTg4eIBaeD+O1bv9ok4s0kq1YImwJ
9X5fL1o4CvT7YIEvpkapD2v6e0ldoCp1tTlN49hY5q7UizrBu1h+EdUUbc4rD9LV
Tx+oqum3/P/jf7Qttw8GIPHWL+ktbrtSkWaqZYXfDk53oial1JeOjKED6w/I7swV
XTf/+LesBieUkldb8Y6DqCP/qL7otoA01i5ikrbBPj/k2X22P14SddybHTodY9hS
kGoB8a3U5UfPtEz4W0DbCIu2PeitKgby66nb9I+VDuVxCaDsdf1H/MqY/nsben/S
61WcZ+pFD1MXWJv18Wxsqi+bv/0+ZTYoIrhSTWaB3EScjwiR6ifjrw+06vrHP+Ay
AvdXMRWJNVDMbdji/AQoldDecxTVhw3rRhNQMQKaAUJoev9rWvocMBm0PMLJ6fOi
8YIfRrWY2WAzFv+AOlB7t22AFvZvUY3e6B/HYpTva/jwSTvNCqUbkGBhbTY5Gt+M
Z0xUmJuEfHKfhqso4EN+Z/SzlYbiEnhtUaNQWQDoBYuYCDByPwOU/4zw7nP+LBYS
/dgrnZnWV2bVL+VcHfdyq4elYUl1o0H6IkDh4fi3I8+D8t1YVrMe9h9n8/DsoDQl
/EQvg381UEkpRhH4NmFXNNTpsbTE8F7m/Uhpdpq2Xgu1kHtsHP5Rk+VM8/LNfnXb
kCALTwxceOy3VOD+i8pjgFDQAx54JfGEVosJhYkjytpzBMzsJsl9SGacmXaRq7Nd
84f/pdhzFQNAlkfRQHm4Oj8ln1vtdDvjjMUd+0/lMXdpZ155dPweckMmSW0It8YS
VseSZyDi8YtgF1eRAfqWA2uyLofnrHTs1HTEpChEEcpdcADNnC6dB1qZ3GFBDBcg
rOLp+/wuHRvkYLsQgXkTu+KtF3SjNbvoY0DndZzb0Np2sWJljLD3SgeIn3MVIjTe
mwMT1RhxzSgGT7ML4Gqw+I7cJFD2qSuf2OJdhvAIb9saDWXYjGcCzK+0O62Z3MoD
99TmBgJH+1CW5thyr6xMX7EywRen5oaI09g2/YwBeodTgY+KFheHIVLG+vxiVfag
50az8gY5+zHX6XFmBRu6/ms2fTm+LevwFIwwcume3IjgkpiI7go0cAMvdrowmKPE
KabJ4b/NWR2CunpNZ3n3qGlFLd6NeoJWOzdtglxmO2OBJuJqDGjf1rGYvsYwhUvk
jxFFwqLnAr9AfKTJ0hhTNBApJavmdfZA+Io0NX/StOgnRDYnGp/s8ZEeBWjmgUvO
47Hfq4w3yrrfTMvVJop0hMv+lrGN783qIZo6dtPk/AijPHHg+hVf5Gf9FZwofEsh
u0FhyX+5INO2xYhYmdtYFSaY3YA8nNiAWbaK/52J6AQYRdtgciqnN5srPVKWsU/+
OmODJEGW2+EBNOsBwBxzsu0D5sJRWycmQfmN93UqIWtZKPiMPfitxcxQBNGi5+2l
GR8/gyMOVmT0tNa2zDoPazMtFb5DYF6on/xpJAYLlXwk4KVLWDxkeBFDegIHAOdZ
3YLM7W8Xom6uP5ZewgmiFT0uCMaE8N1ItNMeZtwkQbbuQZ3OZV5mI/KPqBvOp7yb
nzL2fikezkvzPxpvGGzcw1i0Xws3LnZdSS4YZTFmP1lbtze4BEWIdCthkdR2ic3g
vQsTN/w5mpz+pAKn6GrcFSVXvM4x9ltNVweAxlkBYajJraLlTqua5GZKzAaBfSmZ
hpwV0Q3ezfst+YJNFOfcFT4a37H+xwTMeObTJaq/UzbpRHTmVSzVnuJEMcUzz5Xb
Y4vdN/jUKpjJcYInaDWd2feD3b9AfV8qlej08lrVtOtNdZTs2AdQYWNZKxqHHWyJ
2Wp3lnu4JdLIdUDQbE3/h9wv2iTHWrmlHDOofZ5ty0PmwJGfSXm7OP3ojn/bArDW
l5qxiej6KCzq/qRe2ZtrcCfwVWCFJUXo3GaeGMLwDPrqyUi0zUVQdo8SXaAAl2CC
g2UPAEaItv5wDi1l6mg8Nlf1Na5L+uVLZ5756wmYlQVDnFIVi/cslynepziLIjs/
CdZHRTR9huAjbH/3BI4puRHHQPyhdVSiufBAeLxFBZ7jUwXFOX+2714ChEECTVWh
BFy7M4hCKSs43roeIX9Tzkk4kpcDuwzdvYdNnqdBRZ4=
`pragma protect end_protected
