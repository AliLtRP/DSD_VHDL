// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
m58/8tUmNmSQwEI0Fl3MrBhFeUnBW7DVeLKRYacEFHx5R73ffsfx7g4MEIBkvfWW
+/6Rf8RIepCf6IVlXDBLy619PsmKymZSef3Y9E+WMARNIcLARf4u4Gt4LPguAL69
SRdLqGJYlMiiym07YmaLmsvS/QO/gg+gME2XU5o82I8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 86208)
l8j9T2Lr6OIXDtvrIOxPa9nNA8PyJLA/+XFsu4JyOl4zTiqP9j9TrJeZ0JaNrgKK
4xwECQeTLqY87fMECR/dvDtWxwW2gvWWsiwlIvQfssd5uf03Zi/r8n7xvR4AWeTB
zwVMI5IjDkL05sxAcwKN9cytE3IBe3NlbFTeXsnsYNTJQwmd3ERYzq0ABvxLpIzl
FgONaisCfSOtw5NPs/9z6+ME1L6OmAGGBPOCRK7P75XZrMxOSLuE/dNO38Aq4NpD
+juQNtwso4sxWTszYyrnFl1Uc1kCkEwQqe1bpKqCu4zXm6qlaT+/oLcnDWKaJL7l
nN5UZo9ieTAo1MqEQePOb4X4zfyH3zomY+hAxG+agXCx4RCazBiGAbjIw1X2vvQi
cpMvGl4oY7SbLZkDGikNMF9vYbbLDWRbEzdAkP5iMfO+yz7FvNRpmSLY7LW8ToUF
iwqPNXNuWCjIxjyaAZeCPEq6exD25MyN8WYQne9lfiPGiI07r6l0vNv0iME2Q/fg
klqcpR2nWmS3/Pezs96F9Ywg4iNL09UM4q/v9F1GMvBVMJMvMiZ7L0h4+Ep3bzEy
pAyIQq5+wcn95dzz8w6xiGNEC1Dz/uMWhA5EPGaloVMaD6gQiO6I3ho1ikKOqplN
VOFM0blzEe0AreWdCZa12rLqk92sY2Cbtb6ZuDBrKG+JaE/7n1ctzs7eExRCtTVX
nv7qzvvGsjRMzAXwi8IWQhfoRMt0GiOo2w6OzZFoOXIzhbx0ildBVDsh3hlMWA6I
m7lwWZGiy2UTqV028sEDA1WWsjh2QirRmDQQucJDi3oCCJicu0jZZwDf0JteMGP9
p+tmD4cAbxuXfYRsLU9JzkiWKl3OPmhhndEN7CH2LSSpgA4r55IK+Au14g78lete
K1x4suKabwwY1DiwMBUW6hRvQp3F8DcsUHz7zqCdH/x8ChiIpgWhXNYSsKupmoEm
hq7QCUNakUI57c3bpyYjhKxF9vQUMhlZ4CTh3nbeN8rOYjoe+PsUhopFbGYbxXN9
Zs6oEKYEzqZbGPwrWi4tR1zqXxL+SuN4dbPzi9To2w1N75D+48W3+dEzJ0zzSPB5
xGnNiFdchIZaKWzHEA420UmONFUUJ/0u5E7qZxetqmub4H4/GBdRcMwSvOukvDGW
P5J62oCT3UTTK5QPWuVTlGi6vhvqrC2GeH5LUlQ0TtSkf1mDCY1LLaH6Uwf0RQFT
ZXX36OUVk14BQaH2qSTBNNGEgI1mux+GSwrp26lQg14rdflh5cNJEomFGjv9PwEu
6BICLtNjdRvy/s2K4YHiKDZPWR+D+kxHCpDBYCsnV2niQoH0tBkmPPDLipIwpkge
GUaxoucx6XRMpZfsVBorMNzV5f3sIw86KBE43PyQgHROsOSoPWUWoZc0DinDAuPL
ZwhdFVwFgL+kNvCtWcj8qP9hBBDdJg4d41D+ynf4RyZonL3GJcI4GZkp6r4yyrcI
0IoDUK35Y1V9NyzUc1dFYeqMoTYst2oO+JfS6PqzAO7MC9AJbDvbR/nGXSi8PNWI
aKE0Ni9MQhP21vGzJk2me0kwqfsEneP45SB/vUpUj4aNRilrTsKIlpKnGtVJi24H
EMejBUIMSECrIDOKcGwUKyQ7Yw9cn18QGgQTvHR6Yev1e1bASTO18Bmql9s/R3kr
ExsIJnEBQMS8tFQezDY+E60FyE784CRiZ+1FBsUbSInIWIbBNoZ3ov4AVbLgbPlA
UAUoDo4mguwjS9TarOEvzLM0yG5Y6Y5pHn/XrdC7ECHXrLdem7PTOLK4exVFYkns
sj6c7BVOW0/MznYM+uZpYnkUVQLtf0TlOa/0NLnbdAFhWGdwxywbzky5wLx6w2BS
Hi2VqEU64y4v9/NsKj3bYgsKejTU6qJcd+oxWgrgG+9eBAV+4fAEm/zDdOxQJulL
Av793Lv9GBJcX8/Wy/j8OCH9cjlc01XeNARheRejiviBhG9iAPRDakkQerrj9I3Y
J242SnWqgAyBy1ZzXjFkiD76w8EeHxLzdadxW7OT61zVoCITCpg4gL/FrYvbeE5a
sizXZjpLIA7VWd4uSiDnDTsNa9GSXXrEwqvM93UXS6U4PCo0ZzaHB2iUvMLB+7oe
iC6e+QttoiJ4J/x/7dfITIoWqGJnM2BEGLWPrjtndrXquQBaM9EVyuZ4KXABLauu
T/1opBwHjBHSFhhsaJeboqgT8WZRblm1Tqq9qIQ8v9K8EuSbedWnSMYbL9U3vWfY
nxtwaNblzevu7YNXDrtLfjVZ6tniVhKHeYh0bRxbUd1fTSSPeqh2EOclNF9sf8r8
td9kN3doyAlKSI6aGQDL57PNMxd7UmMwSJNLUWgXs94R72ftDD4kJHqlt6rbgexb
djrF4ZhxBFpC849VWOKZoc9Nt7xTF+6wEFDLfwJ/PZR8nqWE1ieELJg+Tr3ulXXD
thIah1x9S0TdY3bprXnzIj4ScGTiWttemJUSBhOXds/rdz87k30VYJ7mxH3gYyZt
MEj49+9yP+zCiPXDAHGm3LzoGUJp/qYKdMVza1Ebxbm2tZAiqENKR6+ebhuLn4ya
WVoeC0v+QSq2tvKyp5moPbHpQ6USSZ/yQSX4wYhYrIoc4LYQED2iGxOGvoCLjIzM
ElZsaA00WqS+2VEFmf55l8U0NnhrzVdUk1/DifAhu4haQQJhwO6dDCYLdQKXxkJR
/YyN5FIQGvha4Ng9nEzijDyxnE9ry+gv9pOJVdcRn9INYbGxeDl6P8HpBotLTR3g
NEea/R6KA2XBfeWTYg7w6uLq7/MC8Kf7oumkMK0hxixuOcIcipjHWYo/ucUFyUFk
BLXD6mZGYLkbudxqt1aP5VPc0Gev7SnN6BUJ/J4YUIMO1OhWVP+OYdhNhWwWbkKK
83WpD0Tes2WWT3oSS30enRgb5HpRLjpHUO0VEu277pEwXHog+XyV2FZP/ZKmJ7bV
vD+TITnWSvSAVHRFBL8T/7XBUVvjkhRGjiqeu6bQV02mWKaIYf/h1IWNDf10XgW8
GDVU6IMQVMe2p7sbZt5MYAw3PDkLw2aEkufBpcGUzBjGooVPiraa6uwuM1SmP9j4
sEG/lFWbhRbXG3QyBnPpNPvhpS2brNWPrXn4xsrUvwtcjrZeF5bkM1Hw6n1FI0s4
gg/8Ns64I1dvZ3EY1XAv+TDGera2M7cj65Dr6pGwxaNUvBeFKEEZGr5cgFpfUNUZ
5eGVrZuuCvFkae0xdu5CXiZJFlcdgOdT37d+XQDSKmUI7bJe3jvD8/XMPTxP2tdH
Xen5q4Nw1t2zax741eF/YB9SNtnK9ELtMltpZfgu6zvPjsh+AYz20hrK8O6WtMP0
GC6ENAqIld4PyZ/6wZbHz8Hkhn9WkJEiiVNVD0c1YI+1TRqdUrqtW0fDtnfjZeez
fFMLypoNtJJ9xyt75xV6WlG6ISSimSxFjTcloRsEbyd4m1KcqO2oanwuQ/WR25wY
C24gHUmVxo5b6vztjWO0cB3ODdAOnc11A1Q8wZr3somyj/V2Z1aNpHonM0tbiDVS
WLj3uoRMwxxCCR9LbY2rds4kIV29Dkic8Biv5RetxjMUHa8Uo93sa5o3wcrfWpo+
HEhT4XURyoWIaybsG6QRUnyVq2LQ6cP75aM3MmrzrpQQCLTleeGd/lYYsp+HP2W9
H7aIc3w8eRBD3Kofns3rfwtk8lqgU7GWuw4ZbnCIZZHIxC+KAUVo/yz41DCAAz01
Z8VBwOZKtA9KWBEFP121WwxWmBqGiK5z71ei2E3XAhw1RHXkZphaLrlfa+fuS3bk
zHwmWip7RLAhROs5pUcxldXmKrhr7cq+wI5ufoAN3OgfQYMy7GthSOCBiXnXE374
0AsGSqgrZ7uPbPJ5GLpRWhpmwQH1THmlm1lqa5NhHa7GlcnF+hHibS7WoPIhbT5M
6ylK0LgBpdtX8g8YEl7kQknm3pa38LJtUUIUzSuvZLT7YtkQgo9Rg5pPTS1cdgS8
LDIgL69xTi8n7x0giFphRPnOGS/tUgS0QsAcTTjOjXoDRRevLRn0BdpGUSABThRG
7H/bEsztceqa8iWSqX9vEXI7mjBtniHzSKUKX0iKK95hW/eUssPPA37Uw8uXAX43
g8XG/SElsVvL2fhuoumRR4VuKjAfeE7BX/rEcbtYohZDTxzQ/lp82719E8jgozRj
z4cKN6xuTk/TUszCcxoJc7XKLQ/r41y6iUjPMdo0lLw15Jb+TrzQn+yi5/uBB9lr
QBVayOgiHNXFcdmBQnQRArA8xJX0QHqvETx26fbiW1iWVBLtjoSzijPPTauOiuqZ
Te4TMpoOC/PwciEs9UsJ8HkBpmgCZrrv8nOzcERxXIDZ+OmuEAdzu3kO9caJj3jw
OM3vStlnHOyAY8CUuIj93zCT21ccjhvIYJzZQ1mFV3f5aHl557U0myO0ePac4SIl
ChqK2H1aep7JiuAg0SOAPPVe4emxW/Y4z8v1uoNnsI5XJCDKtp1sCQJxqcibSgqp
Ysz7OVm2hMwmJE6KYe5z/TNmw/AaCDnBuzEjnc2nPMqJi1kucSG4uIGhn6r/qbLh
YIUBhnl9dJhYKoVcAVEq4BaAqktPNEih4umJ41yvSOTRBgIXUe7C4HM7VVEUBnRh
z8jl5wQJazEXRxLDtplMWPc3TSFLxSVEJJsLUyY97BqFeZveRiucrpdiT4ay9ODB
UbyQfR9FKpNF3qSeT9bol8xtj3JyiWoay74TgOL3jBt213QWbJ0b+ZYWrw6trPEt
Q0uhYiks9ZF5dAPk211FP4F48v3nwMt18MWEo3U7Nd3zBIckMW0kT3dfW5efhdOV
s8lkvW30yU4u0IGqqGQqLnpik9YFRWLcIKUDlkFRawqQ5358DRqOFjBAhJVb1o/F
jJzZQsoM5SYYC8YD3P6x6yQwGMQn65uAsIUBhaxqf6BOjbSFgdkjnu7aN3LGiXz8
ldlt6cPnCDrRI2gMBKHQ2bJu5cwxxyZvQq+tw4Mh90fJR0kbCJmpTM+rLZoRZT5x
pvseKmM1aGhkOBvyM1eJ4fc45f2oNf+hWXmOQsOdDUoPGac+W2QumS+atJ6F/07l
jBsdIk2iYlMt5ooVOkgeTKGMs9C2R5vMPRClJpT6+k7f5yX262lsOeevIHzgLsiG
UOWaGNg0FRzDtHg+URiYKMI8N/Aw3Q+KF27pVJMuK39M7gB3ZWrYw2PXzKdFmLQL
GkUeJ5reelKm9t1HSQnYQub+jO3Qjm6SXqCZQc6XOFFgVfgz/BkKdu9qUmDK4MC2
dZNr6716pXVsw2hVyM05f3XHJouvEpr6zTkJ+pOEx7m5wy+XyH3syihK/lA/Z/WR
KNrdjABx931GWVf1LcqTSxXT8gFYruTesKBurgiAVPS4vqE5SaegVOQzUW6GfRrS
SgI28otka6ZDRqkjlD7AesYiBNExBKWd9/s8k5dILEYziSWx7cx1zloR3KhloMdG
GwR0Zr1BRhlNrsmtvocOyqAdT3ct0gMJNsC2z7aJlE/9Mgbzs/6ofd2zVtercR+q
bJyXTWK1UaRD6EHrIbNyOKeu/W6Lcly9KrfuK0O/kUh1U2yzlyTOtqs7RKV2cB/g
wyyiCHVIiICTrsQXOtl8bd3znfBADCHn4bOcjwLyQxwNNTaQ/XoLDRjHbSUfYVZn
n0KiTByWqwGJjSuqWSz4VJHRfosmLdXzTmoGev7s9ePdnxWwtqArzSc0ez6PC2l5
MJTTJtCuHpJUM6m707Jtab7AZMbIgbRaivhoHPB9UluMK16Y+zGYLT1PkVU373xm
kWd1qSpODx/i/sLn4NmgyY1ETBtQjDRaCo/TUcRo1S7Dqhmi3iHRQjIvltEh09kr
7tPB7slbtYvIKGsl96OLxEuDsjecGBXVfvBvNI0giMdooswaBjOoIPTRbTul5RK/
O4FfMwNWCokHMg5OPT5m1I1PCyMmUEacEMUA30SshFVzE3uKpwXHPHSLAbT7ldrm
MSN+CEi9yLBPxPyyx0E7nAk+0ZQwn0w5EBaYaK1fpSmGA7ledvrYx0BJ3DtnNBQm
W+DRlwMhg2/h3OMeHBoSr69+eYAgY9G2sVhcN0iwow+xouxvABD7aYisHhTX52ux
l14UxSwynXMPEm7Ov7XlOHUpkwrOjRWZmCUlbkIY3UCGYPsm9ftRqEkYoS617qHo
P1o/cfPv1xbhtJUUMDpHTK9rkukKgfo6hmiCG1bb+zmwv8hMbiDDnShwrOBUA/4y
ScBchBo/NDY/5VwG90h14sNtcuUo2IAU1oY09BmpxxKqAel8tqynKGvr2nIYfnzY
l/GqHVvybmklDaHArYuxKCmtRMxyBuMgI5g1goJDoQoJlz1LEUsa3CnUTZA0D/+Z
uPG6gmJVgHiY4u9xubreaZvBmkk5VtCErmwcoqpuMcSKX0E4+cYqXjOc9C+P4ERb
QeAQabDkhcckteaXaWwh6uI0nGivkcklUVHJfJIeaM91H8CsZt7ZMJaAiTXMDtS4
9qGG/TPgLCyJb01SGK/Rb41SbN2uVb5ITyuqVW8+9IMB4gKyyY4VBAfOYXEB5vxF
cCMTuvS7wrxOZJHE1hRT4YagI6ZvKQ9k+zKRxAaW4PCpzN2lxGbbHfBvQObtna2C
80bSos8wYwpIh+s3IVy993v+QWojikJuH3RJ5D3YTyzxNtHWVJL5GzwBlRSmith8
hYUS0D0mHviTViSL2zDRXI3gZVX8AglNTvleZEG67NKiQc9fl1bSDleKD0QemfQQ
dSBmvUWehKw8qiR3HYeYCFouYikSjUz6zkzbc9ioFIWQVXT22UhlAFb9WJIaIhCm
VDZGiveR/llqwpXf2RSoJo9F1kmdo+EyRO3E4Lw0E4sWizG9vYv/ZLNe0FXIg4Wo
BlNMgSXjVteLMPRdZz9vyxcdr0SIQCp2IWSvUzP+b4tDDCFtfrrFhI9+eD4TKJnW
ExP7Uc1VKuZeK8ymHYkKRAW3Yu/C1zk+ullxaUTA5qs5mbMkDHd/qWVDRpxMy+ro
iKLqimq/zDASR7ar5sz5d3uv+/s3+bzEsCw9BTKb1uvEB4KEXDmcq6wdGFb54ljg
oHjWLPovh+7dsb4H90UZBkowjhv0/dn3VIc1/vtswH4GH8GEhNOXTJyjF5bdNnko
5sGMqC+/uVvKxQB/4Lx3Y2ddPfoGwPrSGvH7nOeAcmdnM8q4rZhCqL0oVmbhQP7f
JN+FRf3pcpX4bK1qIlwqUmBD9kz0WTCyimtZ6QFb+tILt2TzDkVd+vWrbmX3tknj
EBlABJdfNxrIveJOusGW7CzO35yRQ2k8iPwkR1cytbg9/mzC3rLmgCFIqrbS77zQ
4OzP+CW1NA6YAdx+VUYPZh3IVeUrObM0+Wx6+A6sw5VFneP3CtBvYhyoXEaeqkvC
nbdG4siTF1FfEDwZibV7pQorVCXQNNI2ymG74dE6GKDUXqHiv3lWkRIP5lUn2e+w
4VJU6VjCkBW9bfqzjnE34Y5XQM+jJ9XW2iR+93XxMjsxSQTPg5GAX2H9cSYrlCPM
RqUfc67goxdcBHeoc9lGOJ/tbAooBi9Fu7DwpHcRd5Kp18kssCLdSXm1U5K2nOOp
gZZScLkrn62NEAAqBl8iLC7jREbVDJY2aP3FK22g5EHrHpvPSEbYBrzkgVwMWWW/
Urv55xshF19294LOJ49Fe1axQGWlsrLjGYrYZaa1zE1F2+9BsKk7xbKi0XnEqOhd
j9NCaZDVmUL+g+ogZwhplm0cBMgKZZTyNpuK7SPa9DpgPj8d6i04b5CpBtNRrKjL
EqLzVC6IijNWOqnPNR9S4TmfIGOC2V6ciTFO+S/urcSuGIgnVLiz+a864mGETYzR
MRSTIwQJvTrZTMw6DKq9vhaXWNXGVvfI6RxK/K8OojojdlqmnYRGZjdG3pcpIyry
XQ4XM7DwBlkviWXEjlJDBbSNA+XgNPXrav4Dx8mod6O4tRwZs4CihR/0h0U0rTEu
ehgkyJ4v2SfrWGkZyPJsxyPS8KTjMkJHib0U30VkH846mej1/xbjbImVXKKg+9QA
9/utdoR2kVj5n1IgWHSbldpuVZ+w2I1ftJxGwHnI1iTlX4FbME/fA2NY3wj1V8PA
BEPX3jDI1QxlWPjhAEN0Mv5UtDikPqnC7MWlNYc1SJPRYx2W6vmLieaqfRn7pyAH
772GdOfhM+56ojMG/GmBZhuouOpIK2rI/hEjGRv6MipO/168PGacPJo84e5ZfN5N
RqhGicNC4LsBuv/LD9oKKw1Pq1nJpnO8IdNcKYT6outRm9ukHipcRyxfNDGxU2Uw
elBXlhqRfpcL1QqYG72SBi5BtkcXkhzAPIriwHxcYZwtL4Cvj7ngxIWsFuHFQY4S
JND0WXyH9fkLnDHrJFxX8NdjLYACtpo/86vON7dhb/P2ydq/6uVRpVKoeZRc0iCI
ciNrgtANT+lSTrTiME1rxVcE9Na4dlfFyqJEJNIIyruy3OWfvdvuZf1K2yrfpC+z
qHW0ytsLDAZIfmiRzC7Snc52cGMXhdjWweJnE2JNnAy2OiVRr27U3DelMFxrFnmB
6MtmdjCDyNZI8KoJ5c9sfEypn2ZR0z5vkByvfPJluah4k34oaCm/j4oHiwbt4nSY
KDvbyPXhWYjOs3bJ5nCCGC41gLYWX7wEqceMgtRLe5jQ/aM2mfn4njTj5I0REBpj
Fg/eguf853QV6iRg6HHcIaHCkmKHBzSF2gaGwhua4t9wMvZbnTQ+nxD1SU+2IOhR
YHb1oT19VzmUN6zII4RW1rSLb+EGBqjIQqDKHfcGi2jLg9PJiHJjSWh2ka0323x7
ntz7/xBNMGJZ5p5cb11KuWGV+RdE6fm9sSOr+PtfFTJQ9C34za51krnWOGoF3VnI
/3pGq1ocpefc62fEWjzmbnw9lzDXQthy6EDC2wDVl610XN9Em5MDYqrqXenwVSit
axbKMkyuz/YrVdTkFd6e//wCItXUFvNoMoz7rUvDjWj7O6oxG8NJdVdOUX9DfAty
6RiPcpMB33iJjaCChk8NgJ1+O7hOXsvUPfhbExb+zfM2nVYvmPPrWqHMJziwbHF2
PHytYY8Iu5egjv9CzLsfdoQchXUsQyCXE9KSbYP4XB18aNNg78Or/+xXdLDUxAPk
WaFYcKXGrPgR3mFFOofj5al2NuPEaHOh9NVDB7irNTGwxYlHuyuEdY3KZUhxOSmu
MZqKG/frzdzyrl61vR+2N+nv59DIWr3YseBS19ycrEpoEy8Bcioe5c/UH/xQRkBs
nM/nZ62o7MSZf1zGTSt4wma/l5FDIv84lmQW5TZY+/TaJr6eOGgK1NVmxNGaJ/vj
qlU9F1TYE/k4ERzfAIgAu5UjT0s1wrhN7/2BJyv01lZDpYd0QuGvSwwAVTObE8TC
LMlBTym2v+da+mXm89VVQv4J4BVFVj65y9wGN5Lb0JT1ugFcT4nAOkfL/lzeVyap
KstWvXngBXaT4gkhLMbg2IJePqNiypyV2eSAmoO8U0Bqho/EeZEe2TOoN4OS1JBs
NGck+GWIUIpz7YuSX5BN3MWpkiiIifOv8iQtsF+JqVBDf9mPAiWGKP8KGDHEK/VY
6x31t2Em7YpYVf/uKjqzZXR9BdhcsmE/wpESaYKWJ2t9+8f01A465rKBkZxXqDmK
o5yBCRM/WEguF+sQlqqWpCVkjqYt4sesbqXjfqH3BjZXARiHp3pK39uKyVtAnwjq
Pe1/4afS+tvp3LhcTrbac6T4G1WdyuMsoD9mBbtv4JG0yMOutEbaKIarS3yTlKS5
NfoCvOQ5jwpO0BjpdFe3h6P1NdDMi6CXGxMhCONrFrJ4PMWjabf3hGDK5Mw6ECmO
GX7xGNCKaTt9pDTy6Wt6ziAMg1ifmVdJ3u3n+aqVOYIc0ivXzXVtXbo8SVGjAX1z
KYilkYThR2057ukmfGYr5qkzndrbfesOHbnoJvkGm+9gK6kHq/geZWgvn/r5icCQ
x/2COLx65DsM3YBl+IiEmoetIhpbEdmrI5GDBZ/yzM/pA1qkNrmImkBq+9vGXR2X
KFHSi4HayXRCzAwjaI+NCjokso3XbTw02VeizjKV/t93XORvSx29VcnQshjPo1cZ
EV+0Ai4CAyJpJhGrt03jg//GICj8ABNrOOPUd5Sk03gWtlRuqIO5yHLnODj0Zx8W
XwtAT+wPUxUVUJl9iNFk8BOUbH05Lr6K/TZhFBVsNimqglWNHJh/3vCDWsftGaCv
KFckh13AhPr+8Lvb+GnRTMoDvIM6GMqHzX0Khr5oBETxvSFHSom2NasA5Go/sAEw
a1GuQM/KLSmE5BW14Q577qLVGW18qDbfdVDPqPlDG/qHuKBVIr0rRhz7u6VO2DL0
9CyyWCxMUdXATMOmnuT9ElZLN7VJ5YJ0NLCs5jVheAAEZ2/OYbpbUH+Pw+kt0qEQ
01qzf/qmKLzH71L1hg7t4ws0aTClSxf6lkDTmXKfCTPNnUL+anL0aO8KwmTJ45c7
HeKeP0vUOvvq0ei0h07hPAOrfzWcN8VoRQFKt1i9oIqn8lVeSNFAJoOwBKwX/eH+
hShPqykef0LFNrlUpkzePP0C74pUfyzABV+8xaKGuBhzvcaclzEcGauCFZPe9D0y
6S8bAIJX34UFOqqpZL1xO9UmH7KyIQzm7lJj8WpDlvYHY6HEhx4koH4qw+HXiVdm
SlLFmeW+4t2zRKOmukg+pe5Ufws65ssIvfO15dAj99lvhemyC8CaVC8rxpglRFPf
sUMoRRbJD1j3v8EpT2vH+PS7PxfIrBaqOMMRaUzNx4FstjQEVR/BnC2+EnyyB7+2
u73aOdKHsAwPRzFDklOwrPQ1R6SyebTG2tZMZAulWZg9iVvIoxMVpTZNk5AQlgur
vTm5Eo89LAsvWBdFdut9EcJkrFKyDklw1AD9lGxX6/R07rHF5iIp8i4DbCcKA5Qv
7y7xEVQiDhZ0ijN6t5sW6trQ45r0dJP3idZtDvL9AmemgteZkZ//a4LHjRfhM0Xk
YXvZd/yjMO68412tK/T9uYXyjmEzitO8APcpBFAJOsLj2+LjXwgOTLiyEW9tl9k8
JJs9ZctQi7ZV1BJAQ1Od69/FwKaIH6WizD26E9JPeF9CLGxtqYIxBbs0xwQpCcOc
utLA5xP3j6GKqX/Zo//YBmVCzCuSRAMnQa1upkjuI8bBSEcXGFdsRseS3hBkjPUv
K2y30sX7GYsTahyE5HwwjlB5y0hZDdAx5R4fFN6dXW1k31Wp7lM3B45A8Y/h5yNR
Sej8uiFlqf/tDsSBHtTfonlTyFjMl5nM3wZYOJ/k9e3aFguP1dWMmBN6p12KsXZD
PPg2HZZTvddEq7wxNYIpy/ByIMMYBBMvHoaC8D8T12szE7f4rgGiudVAdY3VmLzf
UV+fHMsUsRF3I5KiFTtCuJLOzn6yL9FUv6uD/jQLDpQD5lc70tFOUyTi1aI0Z+OG
a5qJox+fEvVQ6oeUBKUVZlq2mD8NZ2AdghGtdoSH6xEgsdWFdGBdIOX12wmWGu9D
JslRJ5IMN0AM1n8y3gLcQFTG5IDTO8k9QH6FuBm2xaPRbN3QvS0ZTb2EegggYeoe
28i317HDe04CgQAvlXWGvFIcUTifoEzKOjYlFl4wTVguh+fQyU7vU77gm1Zx3tCl
OoT5aAzHxBn98EkCueW8COATpSYAuebLXckSM50qxzaMJlohQSB+IynCzvNwZJDj
Rhm19zG/99ZEt9xTdErGzOHsW9VeK1tEKSNNJLWfpDZqmuadgNTZIx3vwwPP5v7c
jGyewPg64iA+pr9zU/aREI1DMGt3HbgoWyenoMb/RKXPcX0D1AJk1+UCEjZ+qb/z
hDSJR8XBmnxNRT+nTe8PiLjxCN3mOr97s9DdGUSJyMlwY0o+9ZXvZ+fvxKlaCYcC
/+uQiiYchb4hmide0OnSjdekXnJTAb3HNR9PUB9Xf2f/ldtR1IGa6HsLpT7BVZpq
XFMVlsNiwA/p1aC3beMR8k4/4PdMHGnhcZCCjABMCoq1gr/z8O0PhrGj0HVbx4te
NZvhG22MZ/mxRueriy4e4rRo4kb8P8qox+co1tPJnTtAb9EHyWHkw/VKb+tpEN/U
INWPggOxk/zJOxGafYToHBG5ftVsNwqHl4KIiF4dLf635EhibcvHcKnG5ORPqZda
oxFMRc2ybxjLxWn2ZaujtrRObpRXvZWXXMHXtduUgMNw/pb7YQ6PBpcZm3T/QLew
GmOKQcWiVsplv7myrWwIEIxplnTGk6DGcGqyuPXHgZVxoB+vn0xgX1dW2Ps9ngEO
02nKA9/nxv3PXBZTUgXPYrAY8wN1yA2MTnupK/7+vc/N6bFgErCsicJgx/3TZ8mB
lAwPtNF2OYQC373b+zcrTFgxFnfN1M41IoTUNXGDDifjZghWddag2wwNttjUTjob
4ckL2LN+4wF6aiafSBoKzF7eBjUu0xoQwuvEmKCvNS8uRJ5BttweLFPK02UWb4FC
6DpflEbKfEvK6fvVPGGYAp9yDL/3EgbH16ZcOU9EzeK+XKw5e6IHuqL15bhPtP90
uJdpWMC8u3bL5S80zDhxCEYAJJcIT0zhTjnq4+LEZhKqCn+LT0itUa1dL8oImYoT
ZfUEJGCFb2lOiRzhiPkGDE0VkN79ORprWWfGzpk7NonpQi9RsIf+XHTIbYsi1vkF
8fR5mQBuKyCCB7RBDwTWGlshyVEiBRf0AB7PN78pVGDYVTZOK2g6WDlnhN1P6rsw
9yc6H1WNHm7mnREFtKMLGSEUbLPdsPiPCXJYLx3RaNpbdIJ50Kixqz0FlxDDO825
1HhFS8nHa9f52mEb+xOk2UgRBgi8ZPKKbjrv4maQnFzwzTMu4PzeaykzKA4Q/4eY
CjNYgU10npz+0yeqbo0Hj/9e2Dz5UZ7UmRaXscjD93vgVpcbcNehniaHViSF3tdy
PxSBqcpXs2oBzEawQfiRXQFoPRm/MgbvRPP7vdbDxW6Uyydwwz6tXalLJIbDA4Cu
34DkQsJpiHi/7ye3u0Fp4aLsIH/l5As0pb3GHOiizYae2uBDOeC7PyP9LAAtsmlX
8gLb0+ciqEskbKyOpAAVe+8xdjKjyiOHMM9yZj4GPTkcqTANCJUhZct44giVlr2j
yQEh2c50T/ChwDZ0CJyXO9rtnmRjiCCYJ2ZweREmSXo0yTLQWkzst2RBmjtwMssv
gBakvIGxEtz7ew0mPOgbrz7xepqVHNMSGjBSNbk9ZkY0Z/2xnywpqr8dmRhDfswe
qQV0+Jjwhe+lrTJlG80BrrHFQdfUI0o9L8Kti6DCarI338bVqT0qrPAa79D4FDFO
HqsHLZ+KGTmvU/XsmJOIAQSnCjY0mCOaKQkyfeSSap/x8tIATF1O+Zrw7kN0Oot+
GVYSLvaVdGBDln558KAmWXBtbRRZv9ZdrQZrM/8bVkeESv0agj/PTpgBY+ik4hHx
khAngSXDizE5e0VIDoI0ZwTEilRPis+4rMTUP1s4STZhg8bpOzC+7YNsSuLl2EPh
ShOPJOwNSEgrROYKfpCgXRQDThwJeCX3JtuTwzuodfnUCU2H25wfJa4HQAqZqb7d
Bgj64qCniUz4ghRgkImdCI7ycgCssutkXlyVFUTIspu4szpXOFra+OsLHzYYQUw7
qKnny63cSMThV29K1SQxFYKECwc38l4/55+i/9balEEO1D/BRJwcz2sZ5/wnh1mD
BOK8VFGWRvLDjtEWtRWpwd3e09ClTQ1XjAdz1dyatkLgrg/Pa9FW77hEXgs7H4//
hkIZ5ucjOUsoPrZFQnb2E1Q5UJbJhwiKZUZT6tyzhsCVBAVRZNADwdoou7G2Ujrl
SeUiSgsB5Re1AXhyKUv7PRoGwrfwuv42iggJ3uaEhW/fdO43A5emDnd4Og5KNUI5
TEXFhE9lGEUgL0MgwlUDKsiaRFrDMtAKBTeqf7csHc8olUXZ3DTiIS33yl2U4x2c
F4j17iCZxB5oJLs331ZyPj9RXmZu0/OreKLYNvAldOOw7MfK0m3cFS9x8HMqRHx5
y9HzK0X43nJFOIXPkPGvSS3mAvTVIrqgoBZf5OxmBHguOMGXy4X7ocImd/va9rAI
QPDCAkyZQpQRIFhvW8bgxYcfPCMTLXgi26c06m2S6yS4pYjAl7qvZdnQ5pKvOIaJ
tQkZa725oYv2/jq14B5FFJZ5Bfa1SPrpL/r2ZFo7FMsN51xHxzg4CMBY9iDZJ9Wj
mR9XRVKU7GjiRVsLvLdOyrTODk/19BIfQSiNkZL3OkDIkZoCCDvkg/mvZnGYnTck
B0urvudXUpRYdsYLV2XM0rmlQWWuuioMP8xgrYgdP20URfzjaogvK+yEL18gsgQW
R2IWz18/ksri0UIdQgvuey9Ov194+fyXpRuBG2I7CaOYzoKfqhwDhpCEKTaj3RA6
DPQopZoUJca6633nqON5c/ez2yLqbKV3Hd9j3jrsVkH5gHVSSmbAM029l5eHTnLY
lDYeojoqbAaQIHNqotLnMq5Jb6qHxAfz7hVfdjHuhTMZRhsFqDtCeqHW2sfLCjFy
+6dhWXACBd/FKuLiVvQOw++jt8txdjaLDrwpfQQfENS/t8QdxRYJHEXfvj5v3aPz
kmxeifbsTSW2RYf088QWNbn8leTzZAZJVJIaM3utIl9TuLSjQWu1LMQXGyxetIRU
lmfrDfUKsH+vO/rMVRj82oI0UH1B6Dw1pc9+CI8vCIZ5eIho/0iG/cRIgTY7oIjt
IKnKs76yv1hU+a6j0ozFAluPtRyiYQGUE5tLeRsXyllez6X3QZT6nDmwPfjWr9QR
deaeSNOdgmDp83oqApH3g8zjrmsGHZlkxeBRuPciBmChLRLvj3h3GFm7WSAhY5Ai
2PzDj7NXPiQfel3DlPEwaqs66izknP8J4dqLYdbKfoaX0QemOFzRvUT22/z8lcLH
pKweE0PEeXQ92cFz3kGf55D7fIPOSKNUr31UN5OSmZnHqnFBIDgDHv4VA9S2b2aB
bAPLbfMaq0Hu2vQSk742qEeXIr9SfPy+qGWB27fvxzMO65HfgJWU9DfN0Ge4jAca
zoH233zzP18DMIkxI8xdhZH6uX0mZmLXiIlMf3So4S5Lq4nuGnSqFShFjCXFAaau
62XbAr5M2N82IaiCfYIyWMoy1jus5aMKUO6IxTtW4fRZtyYcemEVWxeDPJvi+b7h
AzY8p7dMu89YTrvHv/LXXGnpG0e2L0GiXKjE+O2F8Td/QkWfq1Oj+7Fqn22o0BIh
D4nVnv3mMy21nYu01Ti+GYCN/QUhPsxJv38AQn6wYUK6fWJptq5lLJ2RLRzdvlsS
TPqWcEe+kag4XJXB4P15jYozDpFTai9c5rUOufRJn1qOPEFCEmkl1c78LSg99Y6M
/TKxZIj5rzG3XT9YQpaA8Z9asDIMOUjyJHaXAfH6uiwEXTlo7To4O+fASHlR+82d
zYQA/UYUYqzleAj7YHo+dNwX39PVlRCLoqiZOVWl1rv5yI6RU6Fkv5GdSZjESYcf
4C0V32R82SZVJltKkoeC1kj5H3bRrNJWe6I04tFvVNrQsleYLrcGwGQ1CIg8p0CO
kGBBaDFMiaSLNkWKJH+RF+AUY5q2MTW/FyNGial/Ks/2TaF2ny7jkVMvIm/XIBMS
ZQ38wWoQfFjuEEz1ITRilIL+MMt8azG61YW7n9Apvfb4Pja85iAN7sKc9mbkBQvo
731qqpMnHWIddvnTGlsevVZFTBAfKhqdhAZmf1umttMzr0rlJO+vqGeR7S3FbbbB
xdPYI6fQ5Ray+PO6FzVzZ5YTIgSoyX8udMsi3LgdhMcO2bYKS6jSilP392kFFliS
Z9dIbNQCsV9xVFqKpH778Mamm7+4zm6UPUFWvRnUkHQWTgW3+pC3rm3pYlkrioBJ
aSkVwdAbUIx3uVzbGbDN7kR3Q1xETU6VmWIlqbR9gNj1JCQWq4aFxjhpAKmY+b2D
L+4VO7YpIrajGuGT8O/RfZh42/H4cz/IFYqOVuuRgyJ+jhKFwEm2+6FNHFslJD+b
WzcK2LutRmJIv/Kyd4DBrocOo2YcDusV1jzi65RFKqta2muxk8W5feE62IG1Pyxf
/YOT0O10Dn8dK2mGrfX43Ml9/N4pgRLTO6H8PiF0rVTpfLkv4KADRJLE8KMJVPrm
ZgEAuB5He3kM2uRcHWIsOzeWn3C1DdxrIeHIYieipNAVkaDVpydhVz21g2wE077X
9KVSjRhLkhspgtaT1gratBJIZ0iOwtu/sQAxVP3xbRZKHXnEdrL4qaydodXdctek
6WD5Hk/3J9bR9fbUf4t00JBW4uYCbiXtspwlM4kHcC92fQFUcePT7iRYs0l0klv+
hHyetWzoILU6bzthHTUpNJjLhtTY/wlAIc8a4LXXLeZhBEqSW9NmyaG/ML43RpA+
Ka3PfikCchBdPJU4wPqE9rNBfQLvDWpuLZNJt31lxnwjn8RP1Umj32mc657AwVUR
kIQmrJzSgUSiALVhWjE8niWnCcorvdkiTdoLAi2r88Y95guiv//vK18TPWWuLCup
kqgUHGponAsQH39M+GR8lWn07b09vGhn924ENZ5rDZYXPIPCG4RmPIDJh1lPBNYY
XuWH+jkViNRdaZfxyjF1axpaa2NiqveyGxXyYSxWvojYsuJOuWfOfdjSfKWLgdDw
PK4UGNbbrBhf6TuY6H34xwBT82zp1Lsrd+ij7mKLpHf5f6kGh04Yo/rDctLlIOai
Ml05eJaVozA73YZYV0pS3mdA79b4oyf1GmdKBsQSZxJXDChteCy2eJc5UQ9vt0Pi
I84Vmy3AxilTCd9b1aZr3WNu5MwVOLB1BPXml/DMFoA4YpDBAO8p3MGzDXORVTAe
FSe9xnj8B6R2RwfoaOFLjpDZOK2TvUn0RUXuFLC881Sf7sy4qrBHeBegh0TfPOS9
yv67PKfzKfqzfcaBFEmgfiqw9BSa0qjIMCvqo0Y6HAKVVTnJGmX02NqIweGM7nfB
bJgiTbFlSzDNCBbnRHXMLEsZd5OIQcZwrz9qAYBAc2hpyx86PzdpWOotOsqVgn/T
nA63OaWIEaOzSt6xSMLj3N6nj3xtAIeh5/EFSXFDjPsmtS71H1/6jygkWLuEKLuN
oHr4PSZetZAG5lNtnnwq34el4aHupuH7Q0NpCtloR3swUW+4sheSWHPsIEMmAxax
Jp6Gvi4+5VvySb/9LdqmkQT9d4+2fwdRMjN9Pzgp/B67+VWqDU/DQI5kkHMDvjWl
mVQgimjzesSEONlnWGuUpIkdFE9xuUQvpCdVEr6H4eUu0T/MEmaKe3SvVfSSgZHn
Xbb0I/TkqnZB/MZaO4iAZw43DNMtH2qqmJHzWMPvV1Z4RGD48Snamvk9JLaiXrQV
EHG0ZhBulvX4HEDwlO2W+wWMYz8NGLw0yrM6rLC7bdv9X5phFyAghkFoL6fUwBfe
GHa7al0MdC9tzdL09/0dD4NFeYd9uvDUaHBOX7I3TfQXjWhYxsZFT8GboJiy+cp2
7/mAejlBKhJXdX2Sga+972/V8Qh7OUFMsENRbrDfAsYpB6B1j0/7xkG/5EDVhqYn
FAkD2XGak9afHCJ96YgPi2S5hrLQSdngeAE6vlclJOoL1QjfDH+KF/P4EZAvzNNw
zGDm/w7jdNOoHznIQZnyivVsihbQRUHE9HcTjlSQHs6PPqOodjMoMWt42ELMD/T7
ppin/+tSdtli0xrfjPBI0G0+2ehfGUaQHNaYYjsxn/CLMXHWchTLwa/VXnlKvrzi
sX0u9+iLh1DD6h95j7k3QbKkCvR/6cwp6EPbNUuwIP50NJlKs2Hic12A2HZ5ECPB
pgY3QdwgnpDFYuKmglGh86I/2oSsUt8CLtrgecBtS9amvTSByAHsShpJQnvq78H3
O/RVHSHbTHf3UqwNemBvbxZZB8nRd7MebpJbm4gMqcmFPiTQk31LuK+Y5m/cCtGm
nkYYcfEGSc0koFKl/kIljO4kN5ItiLB3po8z7VeQw4x7je4C2ngSxRDAkQGmbIhl
YXPegQ06Eyvk6+yAyvCD6VdrB2TUWgf8GP85MKNY0UMZ32/AWPcQM+wBpK8VJach
BUKUIQ4BpN0r6zEkKzvD24y84nv6p0OSmL6DsO65ggRvbig8ccP9t3BQgm++PykI
nCrWuvGYWrY3YvD0w5Fx4luS+KrI3/GEPnu6NZKf3u4spyaPHMmEgNJoNoCVu/M0
1dFehgvyzLJR21zzKhBfb3Nez0EZrvzh1tKdvDR7jlPpLfelBM/T4UMFQnqPGK/p
usGBYYtUtIq3JFPfpo5IOcqEfggx8OLc44mAap2O34DhWe+bh9AZAu7/sYeOxpLP
ypABX4hn+7wDTGG6oimZOSJ918JRQM0KSWWI7egW3nikaEMS6HoP325Y/M4ZY2TA
gR7PibZZ3gCFZZPMCteksgW3bx3QTzD15DVEcm3kuaOvmYQw8/1MK8RlIWbpfpz8
sUIPDu7uT9tZpP9NVrlY2Jzp57JOk8Q1YC0chxjcbnV7wpP1EYZg/IczjKHhzXsm
VDygBylmovpZWVNsZ03iwpEhKsXmCbyIQA+smleKNq824UoaZO4SJANntn7bgLV3
vfxnKMjcSW+9UAdfzZloyiYY02hawEQuvfgnaJSzN2cIEJw5j+hY/0AGHufVbbrC
YvrphtYkeO5bLC2FdE3N8W559FlwePtwK5ZnbIgnK7ArZ+K4k+iMLD+j/1Zf3/zK
ESLE6+3nOFz6GvzpP3wG/CK8+qL8/WIyZFdRo/CD6yL2vdtlsdLJRbnw3NjQMAHE
si0ydSINJZKWkRn3rQNNFfdDZI3coEQl4SYCnHpKTYIv45rYZUivM5ZssKQ/Gzq0
EoYVgy8j2EVIjA80JRtl4DPy8nc4N6t2mDlJlyvTGxk3vwR1p/k4NWf8GEohyEUd
GhGAfZEb85VZ7k7csJIfHtihCU09H3n7T1E0Zn6pHAIXlrBi/irzZWkIril0uEVO
Dvh3iw4S6UHfnnyHS2Ayer4eYyOtiovyX99pb6M2BwwwcWSpkW3JeyE2gTUWfBJd
qWwQT+NMYqau+HMBRW8Wx+wC186MLaj0s5NhbIhoelb2Va9lMZ8xF33ruR+P0WFI
5jG+LtdkqOUk96WGPROhEepPbP2Q8J+2I4NL13TF27EWfmKB0SpmaiHShBV9/PjF
dFa+gqoPcDYzF3Qd1yjyFBrS+5XiR23A5jHIks+OrLSa81ZVMAAg0tneg+Z2tVYs
1oFy4EEcA8zm83hs0sYLmBIUJtzIMj1x74MqJD8C4hdti9RJ1K8ww1yQ4QvBGJ7K
VIO3mer3NXkXh0xnXiIFkCoad6sqTfSoQgzzNqxVqw5q92l+ByUHU99fXRHV6rOd
MgGt5kkbzvI2qq6Gy8bZAJyLhJ+59qAo13Bw84dVyfGB8/yEvaOVIm24JJGi+x/B
XLI0DkF2gIOiqmeC37MBcKdHJSTAkgRCOj/cOvyXiOSFiRlX+fxePj38jjJ36BlB
hzFr22G9JiCEhO5rDE/BC/GFKtuuKW4QufNCSebKrJf1AjXEyaso9VIHSX8IxULc
1W3jyb0J/hBUYH0SF3DlZdrwqBVjKmqTTNoZfI1ZQdHmzKOiy0LJMOUqa6kiwM7L
nj6w4v3a3JAIG6T+hQJ8OvAVh0xmESjsIFMyMB1gPddX61xvKvb9ykhUhl6JGtL7
w8E4kivgy4U7XRt/TEL8AzFBNcv0qXnWLMQFhIG5UYvm6hmtJLKnh/iQhAog2BZy
O+Lxliy2d6ENhJDid6CPphP24syijoLLWQePLIvjuQJEkk5LstVjChrVLzGrbMyy
6nGYhGBehiODZfogDtboFuHydFoq4UA0H9+Oyouom8OGIRgZnNxC7Y1kQBVfA+re
oQu+eKYRICJ1xQL2biCapcmiTK9OTrc4jA6LuHTpbtc4drjegBPd6HIWu6m1JSbi
aPdASyP37y6mga9fFuCyDOtpj0XU0DgKW2qKtDvDUVlOa6zPoClz7vMBeC2om4UB
iCBdVfw7/ZbIVxxMDbVukeBU1f7+6ZU6sZQXhlnvi5Az/SVpHtKZjgln1V4AX0FN
c2TuGdPukGSpm8EsdPFZt1ZBYAoYhdzJ78jOFqv/95Fsq1MTO6b6YTjyjLlVCD0k
88jcDmUfkk3aAZVljccp1UsoQhGbyeh+IjPlBK2/3eyOBLvUPK2Ifr9+Ts8+8qz6
OoblnVFcsDivASaNfUJtB/Wg8Scgtm0ENXrvdGlsLQpPYAJ899uiQGfQpLOw1Y8s
cnjXYVLUfzQPYTQrzhdfgpE8iVUkX/u4oBsQqV6CEo3Nn4+ISKe8z37NIqWtq93Y
BeG4nplOW0/4Fc3vWOg2TSGti+BuZvB7ORoCwaqM3hZfv7HdehYb3I8lzAtD5Ugm
C7JIOHQebMuQRl9Gsr1HeKZITsWQr6WRr/PxL6/rm6qAmxpyqPTu2/RF69R0HBhB
zk5GzqO8TCGlE4jJCTmaTCBQxt5Cm6kXGmjREwct2EtcQW/MzKN8a36U5PRvFO7p
3D0s079RBEYUCS8Vj+FzjuV8tYbxidzJXc3W71oliSuga3gfAz+07EtwnV7fhRpV
/PKCTxcpNa2eM28l7lgktBQnj0mxoFAgTTg9cB4azj1YSRsqNaJDWZB6gIA4kV2w
T5/b47wAGQt2zfQMWXRdoJMKhtgVOXL7GjsFAEzxXi1i24yILqzYrC7MRt/ezmHP
eptaI2ZdWiuMmGA1qCFKyIVmOivIkefpq6uJo+CYMj3BXanFEZuxpHrZhIG4LnOF
/K4p8FVJqFG9p6G5r/w6hQ8Tu5ek+y1sNtInneRW/VLsWoGstpiMRkB5ldDyrLGO
UOj/yyQ/LOv7vSCqx9p3lCKbsVjW42wVzzLGZYIsqCW6hGYal2FpDbgw4vGfXgs6
yZm+tlbuqQ/pv5LkxcnDUlK91Szua6+SsiT54b648S81i+fZbKH0cSBSOonuXUGt
Uyiva/HAI+i0JiVX6RWmugtmkH6r3hliqYCwIrLdCvttrKNj3VEhZCm1TOzR4gWb
7NBpiTYRmmCGShiEjc0xdIxfVj3uMU3/veNQw/jB0in3Ecz2AHYdYTC14QRhxU4n
AWUVX0grmZ3FCokhJwoI2HTpaxfV/cSGoMWdPaDPmEvRCKwgLyhq3z6E+di4I69D
lZg5Bf9PC4aGWLW9mDBq2+7i1R9qk7DMZlwNO5fCV+i2huP4liLrae4d/R4KaCRY
bogjzzMCPxbcC8ng3m951JatmnuHUHsTcngygZ2hJfn7DwwUUJBDQ3xVRrG496bO
GchuClZkxOZ8eZWTw2gEm7dpXQcQg+N+b84hVBA9IiZwnJnfVWiK08tnltaoB/QM
9RHOamKhIU8JUMayLiHosAd4itBUrgXIVjA7Sx92bomaai6QQxvfqfkuvyBVAojM
I0DEaBW283YJd8xNCDsaTimlQA5Mk13nvGMcDlVYNFlEQBMXLAapOoSau41ctsOP
wI2e9htDlB8H1Pl92G/4GX/KuGBCxu8R5jVuqVSYPgW691h3WhqN6BEqxSrTKkkE
QIPpPsbz3KPoxDZtg5GWFoWalA2Y/JVlouXVshEfPEev9VNzqbTJ21i/JqD5espp
OAoymgOOVZQY2HwuGZwJ8u9cE1MICHpw42SKy/va8PM+qyM/OyPw5R5Pm8/4H3Yh
Evf12fpV5YuAxc0UAoN/IjJY23FpEJbkaV11//Djr0I+rg/M7wjixSBBvJ8Pz3kv
X0NLjKwGx2faAhtFzurzPH4pOhilIaF77fVEFpGiKIEab/u4r+fGcLs6zkONhsAH
lTAfwHHT/ojymeIGI9FWQQ84NF/RyAmw1VqQH+iQXx5zvgKys98S877ztspp2924
oIkXLUJRdjPkD/NGKe6NonNnUJq3vL+3+XrlUGyUHMXIp/uebQDoHRfmc6N0gmH1
W5RDRSOTqbtRsyZgicWFr4R2H+k4iGLAEFY7pFydA7tdwbqKzRQtXRO2T2dPGiz8
oXhWjOSy5jdtrlxXvoRcSfa66Juoh6Wp4zjE0nJI1T9AdrI1t/weq1gRizFLDZKk
0lwHOI43GSkgE404Qe35g77OkZ3GTxfbtJSYluyHw3VnEX7OW2NREwLW9gdqP3D2
bsFpM7ZEU3iT49dwl/pwKVN860cDxlPJagp4nwCPeBOjzQ5SvEg/H8lhEjzfjuYE
fa2M97a7A0+phr8nIt0h2le80udTzOi7+XLY0Fyvuu9zS2CXyo+NL6ziCrU4BLO9
NJQrHc7YcPNC8n2h5Ow/Mg836JWyg93mFTKzTWC3AK18BgHbZMSmQPWNpeGSnamX
iRqRS5+xBkupSWJ5AngpM/01x/Ui8W5UXPmWh5/Yqhzov3Be6KXGoU62OrRM9UGC
GrtjS88qxRwCPXIA9N2fNpJbxqmkIZqo8ZsCIDpZUo/szhOU2GE34KQOpEEUfMuA
K1SBuKzrwJnV/vvJh1BnDwxe1m/pqs5/Be3v/FeoxfO9NJPnzx1cxMLFWuLrjCOt
CmaWC+ZV+WUp4reiYAMPiqCavp/H0HXDviZcDw7jGlcNFF5jFrlM3skhRGQNSyIB
Eyz2ON5uKR8GsyIBckZvk7YS03p9OCHleJavWwUaFkB9WR2mCYzUg5pg3tTm+1w6
1w1nbhERws0vlqBUek8F19BooZQt8osatbhVXAEujR9CUH2d53n53gFZ3wv+tgXi
O0xibc0VKs8QgIo4wDoyB7o/CyJbqjaoUYwPcoXoT6hTlMfdGKlI7RZA4WvbHedd
zuOfRB8VJPi730AUF+K4gEN6TZM4RV6sFIUcsL9x+pC3hkhUkESyeXti6AIQW9X5
tHTglF93hov4/4eXD1nR+YfdllfuryDthIsmrQeX4a2aNbhhaU1SLUGEYipwu6hr
7taeBsThjZTKYoa40v8ZoxuufBBTKQGUHuer3rAfTH7QEB+eaKD+sZX9AcdGCyqT
8XVn/OJ0GYvQNnUT5CihV+Uln5Qn00IPXns4SVdpecpUUMJUZzubQxMT1V8DwJY9
pb773De7Zuj74BrZUx2EfZAVynzg0LMnbEPdLzmXljWSqc6vvjrnQYqG05q72wXV
qY167CW0nm4OgItSJxDWb0bsNc3p15SdfjpCxhrdNgYS843HgVSiSi3HqZonqFVG
MTQZzxhlOXwK0qVGGkiyFG9zLT++mQqBXM/LhfY//z5lSPmpMDD6xWZmuQ6IfITx
sC0qRD2JcoEUQrmWBcbbh99oRxs2jVFk6wsNIlBb3OVYG8QwRu2Bs0exD2yc0RqW
cADZUkqeDeOveK+rABTyumnfSAkTWrIdRaGpf78slSniTD6QXKgxhpmj1UFEG7jO
j1G5p8DmH/lYE7gSzOjOjV4WvXqC8M1NEd7XM3b3PwK2Uovmdv8ASq2EdcorrzBk
PgcAAu90NxfgJy/FMEeeXoZuE203hXJorMUtCEtg+NppvJOTK7TT8aNuIrmZYkEc
RT8MQJbQka7cToa5ODnaY/NV46SZ+tkk0DLaufqScJXHoxjXDg9MbgxXv5S+OvtP
JX9u8WB78aGE/nPtJMjZMGduUai3r8zM+pDzQTkfBQosfOlS52BV/xbYEWVOCltV
lfKoa/baMHBTLerbh9OwXm5pESLG6EDwuKh3HUzZP0Fcq3qOgIKtEOpt6p2jq79j
2Y8q5lykLk6IQQxirY5UbrdlPautlXbyKIXC31gHyLtTulDuB+IoUt97TIr35SQI
3tnrgbjYTFNQal25jH2LNs8qwUJmg+0vh3ogYJnxIaAPSMVHcBqX/VMEV7aJ0/TN
EK+GxxvE9+l8/YLAd+InxtoLy28AXo2KJe7LoTKvt2TzcXpq5TNfWqcWp5fXPfv2
P/P1J+b3jT4s2OMKYhns3aYUHv1MJquftcdl/CqdhzNzn9v5myXAEWH+J9WfR/fU
AreHMoA1oNNaHwyTsZox+xxM/I4BwIHctHl6b+zvRILHhGOo0BDMUAqUYlh5BJvg
7AEJXM4ZC2a/fb5F6DYQDM2M6sGv7Jtpm9MTiyF+7epzSlydU450gRBIbKOgyeeQ
ICo4+YHF/XYmXPK9Z98X7LwjTXDSCA9OfaQgh0thYRekV3SM5LSxS6OSocSEHP7e
Fooz6ogH8RNn50PO9YrOb9PmicncolCZFJ8BndVR1R/mNxz+tuPaY1F3WXyq8Kk/
6+nH4WQnjQSlvfPbBARP9hRwFIj2FdIxZJUVx/yOV9/CcD6be4l+bxPhfyUL9eY5
B//eYZXHje9cYMzKju1x0EpPTo77YvUFA9eJX1K0kZmPxYs1PIQ7YsWZ1942N7/J
HsxLc+z0P2hk7O76KkVXrPKRCxAazDa0Gr30+fd4WkYwUUAk5Aj+NKL1x4OMhHb3
x7fvY+gm2/1E9q7a7RWZAzgp2M3YdrstS1PL5cHbXI15gSkit5gcVO7K778Hp2/i
4vWW+62ybu+KSoG/2xq3/xn+366jySoOR3AgzF8I8PTytLIoabLqIFaKtiKclS3h
g9sfr19loRTclXpcsRCEaM/NyO8Eh+SM/wiZ+yuMWoLtq0Jwpg9jLR9DeoCmW7OO
8RDG3ZQ/rEm5dpOTe/6liJCq5kPcVsossc0a5B1gIqff8L21TRdUx7H4by8lLDs7
2o2L15bihTG8zELHeIvw/0cU/TX8vcoBw/d3EMyuEY5OaH7DR0DPleDCub6Ne3xg
nX6Mthe+VyYVaOKe38VhkH1BYBoJ4Q5eYgA10d7BPjSS2jo6Bllh/VvUweUVoKBq
hTLkxKzayUQYfJjmrg6fvqazdcVnHwNAu1CEi6rM8JvOByL6B3erYQ7zRbPTOf1V
YYGGV/Z689uvy69Tgf7sWRAIKX9Fct0zxZapEHNoz1fFrwZdAWukgJT2JXSVoT1g
vBcbDOVsxyFXHZ7B+1CqCbkU3bvcQUfQumovaKY+2SfFYIoK+rVpZrKEI8Xn+CZs
OVe7PxhFmtogcuyFET9LDYBnlD9/BZG73xKvfzIUCEH0JgOPCz8U0g4aPTvp2qLQ
awVYiy47fb+11GrYvM/mhTrQpfx1mvzcqRSp9R5+ovgavxkMwW4FvaQFJk/YeiII
2/qpk53g/WKBaeG5Ko6QpcRxhXtt5h0LfJQ+c7np+NLwG1t8QJCLeNOmMAaHWWo0
ZwOmEigyrhVl9SHKijk7fbdc/Ui6YmXT6HdsrGKlBjPUttaUpvSTmFXfT2rSBlrd
kZagIFF5MZIXwf0nQcLLjDbu4cXoSyWuoumpPzOgByMq1d7fzHZafjQ5zUDOtnPl
6MDtHjnJ1ZZKKz14fIUJT10cecDQi8H0f6GJH24jxU1vkJe91GImqIiVPP2y7EOQ
cacsw0pRkZVFNGmkD/rm3/Dl4LnQYdVc6UoRcEk+/kbg85WoGi2tqZ2OENXLaCmH
U067xs9Ge19MGss4bFVJurFeqDz5OODjnoiw8Y6KRho768HG+x73KwWH9qAMvi/H
K45Y80Ft1/wFIKNboWBjZQL4s1mUgzEPb5J9PiDL5r1lIZ1F7C+9qcyZdwrOMq11
cnwE54qI2nd6Mk1rVu0+SygIM+K6CvxUWelxryTTV8ARaNnsDEg0kyABoH+BpE6T
JC4KHftL/VUw06XJn5BxrMpj+j7xP7ggips6XyXoDDNc+Vsf7QgIBSw2pJtzrmx0
ksXDJG1QfI5Tld6yxDf7fO5KOLaj/LTJ3rjRxNZ0JIy/W1daiLyTAh5cKayUYMGX
lih18qIAs8vlse0VieE0pay3Q9uE4irQh2Qr9qIJNg+P/4DFYRzMeFBndqmPlGFQ
LDSE765MtcQPhPb8zZaAH8hAyADZztpjCw+fViX59AS+dxb3R2IGEf/gGRlsV9Bg
lyceKjzv60e7AjdWtJMlYUnRwilzpxGivCHRMN07/RttbCuU3Fidw6oTBaSKYEo3
L/eKg7Fhz7PWGA7/HeLXNBPOlBjdyIW/XyPpLIDva4N1/GK+kzSoFygyALmSSo5V
CdsA8BuuO+H2GeF4yr5KizYaz6/CHkBnZ9/Taw5i1VpP3V+g1q9+/vEZt8OT58Uh
kudF1auXLq2vh5QpykifKuFyiP/As4Mjvq5n1Z3bGWWQ0blAeyKbNu3Id3CegLc+
hc0TPsSqYuFX9JyDqkAGTHsQ1E2C/ZXbqVmFKYYnRzpwLsMmBKA5Ki3km2PmqmeO
b7HQTXjaZjSUdgSKa1nvVagUTpa9cDSPPKNbT0FEhmm39awwnVnkj0OzsthvKcyJ
ua+0yowq8a6fp6CW8iwSsE2wgJpLK3i9de78T9MMPvl8iw6T8B1mOWGIwHAONyQ3
b61+MqwOw3vbU9qydZ/IGnJwy98AD22mD6Ces/0v0zWQfzn7yeGn9uEust5LKglE
e4FZ1Wube2orQ/fruOx3rJ3Fx1FzfTWqgiqZbMYic3V6Cl7xojup3san2F1BmEwT
RVIiZpvn8XcQJPn9TYJQiwnoUWIq1ma7dlioESOu2nb/Eg0/V7awUSuoqs4UQaQg
GcoziDvSCZ9MJI1SlQiYz77vLboEHNFhPbq4LPDGxfQ5AWGUDtUyC3l6T7kNUbIT
NZnOzpoyhpnpV5w8nIDoan9eO3GoNoEorzkcQ7+Kg5vUrgX1j7k/2BnC/IP1m0ve
JxqBMLAg0zNSkR7PnJG/v7FwuM9Dkhgqx42zogWeqg48hcS4iijClv+TBCz1KWNr
h66M7zvoXZ93VAq2CljXKFrAQn3Kzotj1cPy1UT5vwQ1rcJ6PKBIkCoKVFabOU3g
uEt8P+BkNNUpgSglzFed+l7lvqZkYAKT/v5GVJyJd75v4L8AOLd6emoFeTIYQ8W+
9v8zMdPV3unTHe6v9uXn7s7ZVvxdbEq/dg4Dr8KEhG1+D75sUpooUvUoe3IaGoI6
zwFmxDBv7tr1I6T8OcE9bl0zCcXHXDz6HjF1SxXYiKGoeAcl+0xJRJvHWZi3FJPD
TNrt9wobq6wODFo9RofmIalEj/LwqRX9J4HgnjCvBGpaXlzPhNhpmLRK9Rp4l2XN
0OQUyQKN1qjYsfYfe3XQ8et6OU2tua+Ca17ONalNDuoLjnIwyNP56LTL4bqjwK7W
SJvjvmARQJQ8ySH8E/gP89C4rWhVBpi2k8Ys7X8S4szijVaX3cqDf7O0UYkEaQuR
ZP9pzOzKghX7oPJmdexEnxM+bZa1ThySbHj2ue/vfxrgVWNxJH+7Si8iReE0j4qC
3yKINVQ83ydLpK5M4Oi+sT/k82H9P5zMTmBFQTPLau+ZpSVywl8Kv41J9gEI9OuE
QmD8WjQScCv1mvhiW0o4T7Y08kjI8JMnekrCK8gIZTkt6XyRfTlulWlaQ/Psyx2d
Sl/up3mmXZ1+jD5sDkYItxEl8zvB35r6LXiG18HlX6HBtG9/XmumI/Uhcn2Vdjef
FvLebhvGrJMAXObLgqR/e6e/O7kw3muzYSz0ih19hl3WWB156JCElHMrOGaapAGZ
xfCxN9BNeyvxtWfCKtvhKKOAoy5gWOEIfCFm5B1m9ZORT18lAxFFUUF6oNMNUHfV
u+w6sX6xgR7f+l7oTyh00BIkG1jAWS7MlfJ+/klbWtQljsdYv/uNhVMxDhs01cuU
rc0c1XrntQVWhE2Wn1R5+R7byJelmbX26mvLMkyNAQ/EjV8eN6ZB/AcDBaWA0Lmv
i6VqRFplsaOY7UCb964QnrtWh30UrqY6XdRI5AIYMFsrkgrygi5Kx54GRxnZzElU
Q12KogLDRitjTDTXPR1bW1mSlaip/TdneLK9V0O//57IsCm936JcOexzuRQO3lNA
Mei9aQuowj1bwpO5PHKyEGHSbiaC+uMr5RSAxr8bPdcfQ4+pvDr7OvSLx024dAbj
XdkvCRJgf30NMlNr2IYz9EJnkI9lxQ+ZHNXyPmMN2H/2XwxzmNCY6oINXeCrBzsc
pBF5icz+R3TPt1FvsLLOy2SqAafTGSojnFQHlZcQu5KncOKdA/1GdXz1H05dIRZ0
srN2vzM2goOU47W66M9yEDTZkqOYl41k+4faqLpgtBsxEZbuy3VqfuorkijFsUAy
Tmw6f0Uozwv2A3dqmKpszzKKgDeYdKyEIErEQI5mRCqllPnoUVkwbWMs00jwnMZD
CMvJLBS4SXI2v/9M1QBOzHZ1oZoZloN+ULUziQ2sNj3JV9g6ZwNbTkPw3F7KZgF9
YFO1Y2nIFS7d+jSt0einrBYkXlNyJFNVRKIWuzgXvnvoKzy//kzS7fjCCavyq4Xj
YQujGjDk8C/68iR1Bb7oNKWnI5Wzurb9GCdg/oh+zh3s7ST3ch1h9Z5o6n1RDibA
Mwf53fKZyARlvo13XqDobnfR1ys4+jC+uXsj/EkeHZ7rE3B5IuuBXRMFc6OWAQ5n
ouOQ2wVdQSFsSAcGFgAxDOnTZ/oJrOkzQVJR6LjEH3IN4nITFK0rPeMJV11LGEIe
HeUJm2742K82z5z6CyV3sor/By6tICoFZo4ibyoGjXqKArkncSyJ26BXhjh6QkRZ
g3n9GX1EMa5VMEfSD1Lf+N/gpMvs8GjxRRGB4phMgU5uXW8ilATju0g3/GHrkeHG
h1pzD3lQrQt280OgmYxiXv564CNUu4bgT/rPzmqWUtzH5FVuFyVxKGrVqrM+aw9i
6hKG0JXTbBvhowQPrSugnjRWXJ26AW9lYiVHp+5UXE6vN0kAIZktfJon190RKvVB
NxUF8LxrlEc+q0bMmjJmTGaUwPTN9dKGGUas6c0OE7PEd7Eeokq+pV6eA/TbbfQq
83ctrCM7Uf6oLL2wyDyWo3OJKbFCODjX+2ZsKQL5jHgwAa3wrbptN0TYHgo12x/G
3ReB44rkyUHgQlXg2kC3IZA6zATrku2Ix+X9+XalNeCOr9BVxEz8GCRjf4Hi4jI8
nFGdwhiFlzwoDHaG/zFf7+ag0OZpX1lDX6DS7ETBLfTMc6b51qyhg6r1UcTGHVtr
Wmuydv5HzLXl1VDOhSn6kaSmQnw/W3fwa7wnD4Beik9BwEGrDYsOkmjQkMmb4x7S
GQFEylZIDKU2uvGzAG+XLyyW10hbSWkdb+922G0LkM7KOaKuMYfPlJEpknM4m2j2
INW+orJCHw8vfFYpaY6R8y4nIi18WIXoP9GzL+B4vGNpLb3MkImcXyN2aVHcsh7Y
fIgeGnnBNmGmJ6dpUdWrpfEM7Jc2uwy55q91j/TnkcDwXDAdHDXHkGsPfPQPq8Ub
78JKbYJQEd8rpctvlmBjcVm3ptwRhfZYawmADzVfRq5GBzfMMH2wF3MzcoK50vI4
Ty09OihBI02AGar8kyItJOPookM9SYlsWHAWJyhsn44S0cp3Q5l9Wmy9nBouOjw9
iYSH0DPzLwDP9cEBgMcryOqRDdBhy7o1TpOpDrHPiAitTB9rPe83692GOWSzPxgb
EIz5CYAbvZoRUJIGQaUJC8Ufq6UpPQlRBy02Jvszw7ROsOY5T9F8ro7NMLdwiSWt
2LeLR0i5p5c+rrtd1CJuGzu/1F/Ut4b2ROgo6MGMjnWlFRA0fLCA0pfAlcyDOhg3
DBqPdA7ttNQIYkluLs2MWTUT2gTh5VnMQftLE98OBJeRCWGllZRu4sL9BYeo3FL9
RgjVHq43uvUD14X6UnnfuqiVTtgcmNaZiiiAtVCIG2GE3M/fiA71TlPcMW+/Wb9n
cVi9OTr9CFaL2GN+4czyQgZYKAQfqpLNWAgRSWDCJoLvJZXSwr6qm2TSivuFw13S
cHHEVAYXLjzoHoV1lBUUD47GqUPQVE+gSlY7DE0P9hRbHZGFLQbVWjaDFDdXNK+4
yriEwGvjaRsb9fL64yh/Y1xbZtPXNkAEkvS5k6sIJlxDtFItuBY3omje1fgp6zPr
xYv5i9KC9h9IpBEZpNybEVcZj7WLYhLCw5seXZDPwaMFnzMrl6pXyexJxryelWZi
GH2JBFMm7jZXgN40dp5rjcBRGsOAag8X+VFroZCGG3Fj8Bdb3LQ/lXYrENQxT8sX
h7f6AVbgBHQ3QKZ6fmQkzcgPcOdY+gZfP2YPJNFA7SEY9PKV2jdCEHieT6yiHoE2
K/7OTqgqrqPY5QLt265IOGOAKaxM1nrt9t7MY6Z6RweAuDXYfWs6XS7g2zTdcKUs
nogzbKEsLJGk5nI3ioRS1ECOSqVdGNqWLZ/TonGN5nca1gBIthJlbLwy/3Kz0Dhq
Y9guHEu3LMHDcd7F+4NoXAuANwnRSjlrgBsS4J8jlOIQAmenIm+07A6q3c0OTP6H
PO8MBcl1coUyIaNxIOKRQsKEEIRGWv/L2ZfhhzfRvQ4Gjgkemgq2cEBZbjJOpGFp
vkfsfdNZzXjrcCaN4blNBv7XAtLkMTAXDAJ5INGno/6QYjGHpG+yh3CKySKsZuoZ
hF/k4PFr9NN0PNWs1LUMDF4xpkiZxTfj9W4gtsHHvLlM5odB/D2N9E3hEXojrnJf
jyLCZ5hdd6N9mFtPJiesTBD+6PSBzMoeFt/5jetpLx1w4d4xKzuQlAIy0V5RRl1Y
xeQXtQPi25chKvkbZW7uG/WRBW4Xxwv0gTfOMGevPyTJ/GSOeInqezXhqegnGqeA
rpHLf8fVwmp9Y8q2hHYtb1tbSsnstsiq/Hxc9SNWIssiPtYYxWjWvGHELMkb/ODw
DJxKNWiCKAtyIxj7W1X+ys2RnU+OWT5A/uH7PlJ1PRT45T0SnpimKj7L2mK4/PIH
N/VuymKupeeaIb0XUu3hZ8EwHn2zNRwRvOMYONp6SMilILoG1hhaeb9bEijUihc3
dIOX7pgfEgvTLWHJQRjmiZ3qmZJixSuI3+IodIAatzW9NlowI0QcvOJnNFEjGUgl
6f7TYRYsriVbE5k5CXFhaynacfMvteqqFIGJVIeAZENhponYdVTiw8Gwq1anRXDJ
JxgPuGE9qSxhryeUPRxTyzaiZ5TqDNMDWM8N8Yz0fEPM20WI4IXYCEWaIZdjzbLY
NX4ehgXbx+lfOMFm0Pn0VPaQcZ9NTNcm0suGCuEavRql+4la+cWRIiOlj70xqKX3
cXCk1fwqsyMXTo0Vd/sTFAjDrZD8JPB/HJITRf8Cx+BJ/0peRlwBNFNnA2OOzRd7
4DBLR7PuLgmqnaLVBhvvaQdeV9ZNdHRMfFyJmDdaAlLYSsgY2si5OumED8pF7SXi
Gyw8+jjvSZn53mOLYH4vnpB9I2dw+mE9lpxA2CFeSIMPOYIGuYSmFtqO7gy+Rtxf
mrlF93TVTdhPGGL5YRDV1mSrC4VrnKkbkNmMFBQM8u6Eo6XYC4tmJPFuvl/tbTDg
Q0YxH3ye7GvGS7rh5BgwPRcTFjhBev9Deh/It50jRb+u2OldZ7aEmkvyq4ym0LKb
8Jp8cvt42Z4tuCBeTWindYsvLAwu2zV99xTZgTZWMnIImz4X+puFSIeIvxIC/e/K
x+p3sZXUk5RwRVZJYuRibTx6E3TAMBVKxDZNdyfF/IsEa+YmcMPNqDitk0DEdB20
w1aK3K4q4QNrbmdoFtuBMGUGZOm57ZaSf4YhPGpbdvlDd+eVK+1LAo5KnJTUn2Jy
gFtCUS/Zzc3xuHLrdZ7zTJvyer1dOblX0n0e/if8D+9i2yCP5CeKwebUT+A+WPC8
gl6FULtbq5vgV+M4h9HxrrN9LBe0/pjDDTK4qcv6oE3yi2s011QH70XeTrw/Ma6j
mSp+JcONn2ndFUzW5RHVQds2IlVcYfRr/+FP2pbAh5qmqy6QuOqgBFrDDMY/n/L7
oX5gtepjjB1uBf32DKEJH2u/TqCgIaWSliQFv0KjHD9Oyoqb/4u09l+XqvoMQZgw
sYOqhThcgmzyT1zzIFR6BTmNZUK3ddljKoAq+/0z1P5D5CEm5IvDdndPjm57V0EI
yAkn4N1eJljZj4LNgF9PUSbOfwf+9rY7kHpAiFcW/oCrXkhc3GYGCPoxTsZ+inMF
6/p5r3haR8uX7F9QposS5PYMTs5mMe5t5PYL8EGVsDsufxIamdwhkLHUK3HVIlRn
XHm0o0NoVq+vdjKfsxq+d5+WAq7zxZveUG/TtOGs1OMpC0AbS6mESahj4dPXLveZ
5y7JrzK6e1/ZcJTOWGMqguvRwJGH7tDW1PB+X7oZaJD2FPP/RKrewGx9CBKXr2PV
robkJZXVcn3/JlFQ3wcj4iBzld5Amu2O4O4IWIutbuFivHt05A7X8/fuiTU9lyri
ZL38NXUxUHDKLTO8JaAa1Q4DIw1QP8wTYLIUf07ghhwB2hQgY4l33+53bFyr+tzr
RaBvX7c/XXMy0rTEbOb4Fak/oF3CoxMO/qP81YtBl5Vk86HzFWlZHYwmTV20NJEo
O0HVhLGu12K4Y/TLvaVIbiQeQEk11Rn5Ku3Je/1BN96dmQgAmo4aTcf+BpKMlkt2
uW1C671zMNd8jalFQe/FfSTO20y/NDLRCNiD4hQmf1wDmloaV719QBOLa5Gte3ZO
CTCrfd0eNwdSUbg2rqjQCc3zwpAy6EfoiQ7Zlnm4RkKt5vx7lIFbs+N0G131L5+p
DqNO6MKFZBOSc4FTVxSCkfjV7ysPOxeq1/Iyrn2vlqPHKucVvErdMF2TVhHL0m22
9gnUbsX/XauV6d6aQx9NLTareO1byuN8jigs8uNGz9IZMHU3wl9FpD69AIKVvq+D
vWc2tG4T0W3reuk7ZsMzOL4y9y/+BZRmelHNg32t4aJMHBgdW99uctt3bGLwnYoQ
+4KA73OkuitZwX/3MNI3Znmp1wAYoMRka4IMod2H/YEy4EmDBry3Oq5FxSTOuMaJ
B6jQDscFMBcwnVwSqUNWrV9hzmzfubQaLpulpKiRvOJ74VxrHGgwKq4717WL285i
XiQoc9dpsVRQCVwCpa6zLZFuh+koQuXVECvMH8ZcmMp9DP6IMDuYq2lRe/VGbOgY
QJx3qT7DX22dFDKzg1u0ZmTxyYXlXnVMfWoyH2pD4oTjVXBpeklW9FoLgaRDdW7L
aujZXuDYakgnZSgkmNpIpaXgyg0GUFt+yVqZEtCopL9HTR18ejIQD/SBisZmJ/M8
auLBvn3oaKVieX7R8C/E1dlNx1Eca0ILwQX7/xj85SaK9uxZN5PaAc2oBgTKKKMY
fHB+/8oE6MZgPChdleSPffWqgfuH8rSxIzeGd+FvxlYQGGwBFOXDfRPVDXfatD6D
twMUtSH1jtQCavRBICbPIFdTxvTc0w8xM6KOF9K9HePewDW5RnHPZg51EyvPT68P
/qarl42sW9yT2RSwivHswygvNXYcHJ/fLYda03vP7Rcgj5kAumUp2MlTHlQqkjPa
9xsrTOZad0NWEHDxrhAT5JFkUP73dpYPpSCjHok7KajdJBFFzds85KbmeWO/j7XS
cOTkkklbuZKaeWEw1muElmoG+YG5F/DHWBNoKR8ooddh5FXx42yqy3/IHzTwlTFs
gzsHgEvPlc+0W7mPqbYQ1Aa/HhbfredMM0k+FkUDvMp/E0NkOzPrjxjVU3Z3xtXL
ChbOWCeLYHUqdJfBNP/aIU6K5DGjU83+XBvCmf1UtNWjY0VZulRCglV7C/89wf7p
p9oo13c0WRENtlewB0RCqaZXx/GWdbFIVFD1Rr8ReS1t1uXT8QNVzfmnJItez/Sq
N1NOoOCa4VLkz18bKf0R9UMHHWkgKcOEnHLOlIst+J69c5QWU6KwOFdqJ1LWLvGk
d7GMMJGy7Zmh+SnEcx+2Mu+bqZBNFVK+24rFo2futMir8RSSFjqZuBTm59yXMg//
Q1A05c8e7L/kS7THDO7aWW977awMcO3UrvhJQb2JXWRBSQMJmPKsI1sKAORAj1zv
4vZOdiCV16bsR7BlaM9trCkuA5uc2E0kaBmH9h8PnGRlnsZXxEfeXAw34fLmKobW
vs79xLMUj9Ykg5qfHgD3ln++5nv29LY11+CZamptsk1/uNEBfQ6OtB8RFeBR6Ise
blaMZ23GP0SBtnOrwxbR0asHVnguvBeSBR9QCDy5OUtRCqjwwCa5rkTvwzQOHzNG
UJbA9Nv4Fkz6OsyTFDGZQTpntnLevrWqavxXY1yiWKrgNRt/IGi1/ywp/hwpWJSl
8ZbfSaaTU/ZgCjIP071rCxQpRbmLcbzQVBHkTGYEeXFryhCQZvKNgqd3Hk6HWc27
jlzta/Vqwp7v8Y4uMeu+YrqQmwcT/YAA/nwEZ5jS5EaBHY1/o7JXzM3b+OoWzAD2
ZMVUUa3tDkszMUhg/hJXueYo0VmvR5doIYQp3MVdYF9uJX6r2xZo5WdUaI959Q6G
LcJOm7WQLH41sjVyJfel3tyN4gceyh9gqt7nutLi5E0Bz6a+G+Am8cujhuyvJc3W
GRhmpV2FieXyjGwopD5RGL9hcqpkUBAHZayW3nYbo1ZiQz085wDdmv3Oo29HsggW
6YBDbicEZVtsETTn5SeNu/7GsUbxw/HSt54RFHLj4Rrj5FAQYRFY0xGzMMMGbNjD
48lT1K+ny0SV3HifNBESImKqRszUyC53V1Ynh0mqAV2Pwq99e7rR509bnkM+jH9h
1Mm5lhwpFkp4+czEhFLeUUjSKrkd7aNJNeCHa4x13WHboCT74qPpv47P7ri0SvhJ
0Jcg10JCrcnd/C1Nd2gWCT4WCdyg42Uvy6eKJsvO8u1XJclLryRcMVWvHmC8z8OP
kYqyKXselInti/GxXOlV6XNsKk/MmnSJ/fqwJ76dhIwnAo0xsT6Hyzj7xqW441Uf
rAtSJeZQwsZHTtvgoWUMLTq5war+Gu58M0BaJgGZUh848xBN/W/8DuN0T4yQpYJ3
1WnCKh/fuxXfR5TXHLKszTIhICj89W+w0TA2QGKq4+O7BkRd8/hz57wRzhMvu+pR
tlLCritqvDAS5/T9B34aH5C6AaU4evhfHFvg/vN+hE/Ho7bELm5g2p2k2NrQfjo9
/wxg/O7+0aoiRDkDlJgVF+b+61sX5MaLf5pVKkIWN2wneb3kfEeC2kzAo8G62WbW
dElSshnndOpsfgvzMDQICZD/up+oItnSeN9xMrxjwxcEwyljKKrVUUUjZyEtjX7V
As7b5Ro8blN+H0oEpz4r1dyjB6r1oBoR4EupP+sty1qGP66p+QmtmqEpuIKsDK6t
tfjujvv6gtGGfgm1aDcLZZx9uQ4XsREtD2d7/ywEs4DTKe0I7vKW8RunbkCEA3PY
AEiFLUOqT5tXFzVY7z9N0cXqEAG8yI4rKZ377sOgYQ686ruitazkVE9JQsFs+M+O
PI19Pt0Bp4VxVYnhbjwN8u/TEOjLaCD5lxgvMnDF3D51UyUUR86ElqbmCt6LhjQq
bUUlyo4JELz7Be/dHthJt80fRAMcFe//IKQgVp0jQYI4sREc+iHCz3nJXjbw/jrT
Cd6zg/z7HTVFCw++WKbGBX42TKvYzkfHzKHpmTc99g6i+nakyyATA4+1qVFUw5OJ
2nVTUaunJHwx+iSbbrIaXXBZn0RzPlSSUvYXORmO1ZfSQXc6NGDBr4KGF8ed9ukF
LOylhSkHkgIK4chEx44GymhI0vD/fVcwGid9KLOW5F78cIhCMQJacXKKrYdp9H52
3UgcUckziYxG3J3jTt2UprjpWmOQE7oo+XORn2qei7w1KKAVzgYK8pgjsYdczJU8
HS7NZpXmCG2oKsC/HZaydDUFrBgaYTTgpCfKqFXjoKRLjo8rAcaVFwgKf72BI8gE
mJ9mu+h3EdCjH7sjPV/+OP5TjjAbB92S/n7PLqQeqZyUWB95DxhHCGWmF5pz+mSt
LS9NpsNtUbd6IVxjg2ezHdvj416GZ0u3waww2imIGmvdThpM0q7s/ybCElNP5+WQ
R5+ywls/OaK/BvtwdY9zhCgIi2/tEtbKsV66KTu+eBFRQ9R5aGPXiXjBsKtSoJ5L
Oh/ztwjNM3JTcQln+zVVmkjpgLfgm+yoqbTM9REG7MSWmJnTsWA1KrDtp2R5mAtr
9RSg0XadYogjGmHy0q5jDBHXQquXJecXueNCM8bM8fAU9IUb4MBTdn9FJTfdaTtZ
Iq44mJSMS+KiwWQ2fg1g5QdyZxJAKVrooUcAs5Xp9Ptq4rvnsS0O0FfoJTHQna9i
N9sHFuqV7TO0k9IbFdPpcSrqXLpA6vV+2lgKShxLVyaX0LMt2uBLxHhJoIaDj3r5
845KfYhaqSyxaZmqAxOHK24gAwl/FYpI1d6UyLAMPMJoRUt9lz8kNCyf1FIk/H7j
N0VycCtg7hKdkDcC6tghxl5b234kzul80wp188lkKy/3o3stjiKXiu3Q5N4eFhCv
qdvEE5rzDgJ6wggwHzbQw9qY/aACCsihMzJrBMtClYpGEwi4G1aLAlo9sCvpgWmr
Qnc6oYQFgTBQz66fsuFeRP+cfNUy+FSbV7eNJrUbDYpKXu/QWH4tYtvGnSXx2/8h
pLBGyMZSe0834KYsSeCGYCdCo1RNMF/sQXnSo8dMb1L9P6H9a5RFcWHY45ph2LPE
R8NlqQY0XNOCOoXBAe5uy5Yy1YUobDX7dvhSmXy7KLui0aCuifbVliDNzPp5lZ7o
bQVv5eekkkluX/VbTRDac9n8mffDJFAqjYq4XPqrbEZ2ZvZy1Y6C8+PjnyffTmcW
YFjkhUOk+Yv7pX6uxXItajT9Zw8wZXpsTcbYI0uwdqophp7kBUxT+XrYen6pd/M0
Vdi3wnW80MHCEaccHX5yJ4pDazyibOtUK4BycPsnGU+BnmBr4QwbTGbCflezWs3U
Aw8NmgxqxdASWWrcQMYREQVVYehIuHcYEgSydz/FLhBft6N3NtSJsMylGm7JtCLH
eJx7AETIjFpAMRCAAweSo+e5vahia9Q5p1Kz7zZMeSfOg493duR6trMvcta2PxHk
AVLNNNpN21Kryye2MuCvy8TPB5sPJ8+pjTGc+zje82j/YNH+p+h2G5JThSJ2PFJC
obn5zvFBlW6xigGMp2i2Hs0v2c3Bm6gHfmbJeu1BEVLce37JS0eh/bokCDx3YR78
saRG35c5/VFVjiHi7I0Q3bMZlGFbohg4dmrqmCAgICPaIVWPQncQZq6UAF0RVBwp
Td7RoYgQbjJWYOu97znNp5D/4wcli392+BvtMeGDkwaQH1J0Sj3L7W5ZeTjhgSxU
Bqh8EmxlzYd4ulLKieM+iFA0Kwd/nj8YrKrAO3zAW6WhsuN2AoNOhMuyX1KP1QTZ
gsJIAcUvtesPxq2qa7oUC3bTpiH3bRLPh4dWtRH2YZok2awGNLwWxdjm01cKCoyZ
/pIl8io7W332ChsiLK4ty/XTew5PVQLSQrRrtunVwGsW97ddLVL0MSjre6qR/LFO
sJV35WH3WI4dsmvcuDm35lWsgfYlN+uzSrGt7FDKrnUaorXLqHRB52f4SLz10HaI
e2sZY8nH9E3rrBk3/KgVVtNazjAg5gnZh8DP0xDJ4wuVPbehd6g3ZpSF5HP9NOhv
abxGsFoOhjBjji6834uMdnulxMhKbXX0CCgqPczNW3g9jGHiXV6VcYrQBCA0GKRb
lLGctEk34QTqiFBba3p9gUF9VP05fWRJFqNVy1jvcV0fg5FqkgN69oeOA5Z8M8f5
gDb/2Sp0YQYwALiRIkBEvK83fhi1bkLKcOkjf13An1NUjm+zzVXBFKHhJ9kNOgJE
IraGPdX2ztFVm+mnz0u6iMQ9OAvELXDvXRkN5vThGDE8olVXp03XyLLFl06Y/56U
gFOWnpRuczzrU+EDmY1SUyMxe7lh7/sYnl/jYW5emz81FtkSyLxG7Q3hguts8+cf
uacinoi1psLsUixmYcIxZ6URtcy+vaaxVbhTUrPAEwsC8UPthaXM295yvLwHmp7o
TUIlMsvPrQPJaiDKcsnHXIF/U3uUHVk/UiAwdqz0vl3+4O2l9I9UcPZDCslc2xAr
NpIlRw4mhr6Kyq7XKcZAWNJpyEbwCTdwqdEqT1JGWYRNK6yPz2QFOn8bD9/TulAN
IbqMzGuHMPUT8lYEpQpKez+yplWY8Bdz1Mhxs395ou+aZcZfbGlDtWs1qIa0QiZO
NpjsIpNLH5ZihDxmsP9P6V6JplT8HqQV4h0JvV2H+1uqqo20yizNpE/0t8PueZRn
J3CRI9jI3a2ubVsSNQ1nU3wN0QC8g++IkAjQQC4v4+EiUiKnBk1b6XG4kOFIuZHz
VpgTN7LDTc/89XSV900p6w+HfcYMbL5jGwSRbSSyYEmJvL2xK6yw7akSoYfFGTE/
/ZdJMVJQaTbR+g1B6T8bx5JIDew6wOm0aRAsjgyAXHb7VVg37kXaYMZrKH0CMKmt
d9/ZoAMFxRkwgsFZPVvEKKKUX5RO0umG3mtCrsavv5Wcgw/nKrFWViXxBAW5ayEy
tTPQy81y+7LCWZMGLK9a3B5kbbBymHOhJMqyvTQ2opsJK/OELbymK5wAUxGZV/Br
H0fu9rsFAnM3POmAg8BWEKdWc6iID4EAY+7dSKbHRssw8oe84c18rGyz/bTRTe84
Hco8ZM0huSH273nu+QyQsY5TwvqBbVuWtIGYGvUdrvXQ6TRpYlVsZHCqT0dv/X2A
AEmaU7bQNfx0fnGMsjLMDRNANEfWxQ8BXFnRc6YrvHSmIkFNy6Ib7cRQdskAs+aX
TVhzKwYUOKFtKCUrEYYnWFIEbcdAkkYchDf/8MA/pmEwVY0pYPhv71JRTcwWj4Am
gRajAT7As1grxLsUWKGDeD1/nin32/7lCzBXtU6RypvPtbyy6BM6IgDVVQXoCQbi
cYGUUtqVO5L3hy974HU8VjBb3eYxrgyPSUqwlgQ1EUbfWOLD8ISpvrz1QBCRUDd5
0Ijr4kE1BYdmBIhZ7Um4FkVsDze32DwmcGMWivnOSTY0pCMq/7TYqO7V95K85l5v
Aj/pcuD2WDvGQYQsOwGqwQ84c+2r8Oa9uIl332XelHuDSAyp8nV9gJfrxx62Q+P9
gswnVMKthCUxT1yV602JftLMHvyZrJGYTpZpuK52kogLRweF/J4fXndAOBU80SO9
flJ6gDEa7/ChSyLMQb72AH57B3s+FzrFrHA2UYoDmLd5edn1ukfp9B/Zf2BglyCn
3frdsxsq4YPhQe6R5Xv16Fenk98/AS8vRY2Kge8nIiAYmRbXNEhyriI4o2hE2ov/
SINMFdME9RqLGncbv91PhdByLHPMmwaBFyOhuWqeBxM/GkQEiq5YSSkwy/VmIPsU
B4uou7AQaBoEidnxK2qqacmjYynvWZlcSzP3r7V8skjs0hJghr7hgIEAPtICqpHF
cD/QD1TKItcsqkahxCdMacYtoxKOLeqLOliuhdJ3gvnaB+ga8Zyi6IFqYefD6Oqy
F3u6/b2vqaL0vJ7H/BEZnjN91yykyRs2LUnpJVUYk1wm2RcgmItbF0zrRQAA/sf9
6ZWt1b6LVr/sqTZ75eQkvBupqVRMJwoFztcOpyK0uoOJVd6kNbpWm9EV0pnZOnoD
NTcAYgopumwHVHmMelEeDRfrP4k9id1Y+atlzNBDwXi9E7RapQWadAMh1iPYe+o2
0peJC35YEWjrFlK64PM6VNqTq1ChSNU9ADy2fx3cVWjKY9eQwAo8oLTapZ6z6eV0
iAb4Xd1WjG54nf3uYeT2Z2FpEi90+cPRtt+JyQl4Iebnf0A8e/xAg291DiX3HYfW
dM8dhApBGHE4Sa6wwQbYyRisojEM0Y5BgqiwV+x4wJVdFuVkq1Wdy8ww28x3gUY+
OK5TPaHf7ijTtzXdtCo7XbUDfkHc/TtBuYhuYmoaf9kSOryXha9l3MUevhhuEPPr
IzwQdXBpaj7PyypWP9T8s48A950afqkYRUq+SmW/pNksP0dY4OuPnxjmXQdvbM9i
X9rHGm1LHS/V9iZUCk9SuByYsLqtX0O3/bjjN5cGWhHenWrha/bK57xhoYnGJTBX
zG8pJ1++oh0Yp8/E5Ij/w2Xc1qMAVBV1IPumbdDYL+dVDNgadiYLiqSk8f6MWElq
7aByPkEAV/yF3uLd57lx2iNAnQyWUIT7a0yO8udYDczNcO5x/18e7zEGRzQJ+DSj
lDyQfam1b3PGjtOQur2Gk1BWTNBM5sO5dDtUdGUfpH2hjoGMMLq4sbV+OUdj/gi4
iwG5zRpQDhau1JgSN1n7J6tVgsjYIo3bLPanENSlf/m5qUodRveuQgLatkVlnHjl
YIHQLrgJoIo/m7tEOyw+gIBWaKXayl9rGDzGz03EQ4Cgl9XIaeiFhF6O9s8mA1QF
S8w1WPvmv4nUdVZ8zoOBDnxLJcbOGQeAbPRuDyoVX8Xivs0qDeK5XqH/bTHI8K3Z
tvVqx0dZi7K6+Pn/fxriAVLaUK2n6/KFZwex3zc1UY2i4bndMDiESklA4yJR1WNF
VQoUaltix+z+/oeER84nR+47V810VJstDNJRp4f4QtJLUQrhupPqjEPuHsW52Czh
Xr8t4kE4EbWL5lvaD7fFzXuYBgFj0BYMbS8FlfS4wlGsSWh0b9aZgemY7h+LBdik
d8c69pJmFOXlKyqTignjLvjf33b6Ba7b9nA3q+KqsDyLAaKIAYfNNm6fM6SKJbWN
TELwHJwb/ElzV0klvkj0qyX9k3ebH6XtKquvoi6LLws1lstfP3j+BLZouVdoTVsv
0bI2poa7h8vVL40dqH8S8WEGQQ8lbZJc0cMR0ewNQ9ZkTjgtdzC3lB5WcE6tDPIu
lZ2Y4ajbmCujqiB0t4XDpgc9MzdrLsLWo1sZFHy6BUVm/UKWbijcHV3fwWuiIaqM
S2Ff7N3iLL8zErtv5RiVRvziRXWXjTMA/gLfRLgU+PIVrMgS0rKhGJG/HF5+HnfN
7Vg/TLSRuQyq0clgHrx/Rwf/Cjls9qE8feIwosmD5YFwi0WSuIqu8cbUNbOoJL6u
N8thc5Dadn7OHB4rtbs5jLrHBRMgdzcoYHFgA5fVILXeAJJ+wXujKEcUoLgvEuPQ
4WWJpcMtF1EEgZ8gXw+AetgVKfvwRdUHodxXQ5x+zVKpzu9TsnHa0u8kQmIcpOcj
nAvUbeY0LWjdah9cHO+W7HaJpGCg1Ik3p5L9H1T0bozIXNdBSHYuNIbeeod3loN1
t/mkCa35I27/T0AbvAmvwJh4ErJeFAuwZ/oqALqUDM7hczHvRnwmVBhK2nEDE6Uh
xoIsCTmIKUniYFz/4+0lFs5gryg37iaQ+Uee584LWhsXUo4rvnoRUINXUO/0OH5r
BhmyLpyfyHEUPHkeBjNnW431GLSZyxHkjq9KFqJ+XWSM7AS2lDs0ffNR/tJyvJm8
Wk2+Jls7qjxjKBjtc8FbySn7NQmDKvtZMAqLEb80CPI3YNigKftCjR7JcVW3wxck
6JwR4MclhxcRwT5FD/1AAJub7Y6WR1Y1zV+DsKVXuqRyEW0FM/WKyRmx0Bsoma5d
OBsx/fttkdne3H1tyHZhLnlBS8EVix6uo01vqQS9nTCN0Yzp37vqydJrdfzGYOCK
03zci739FSE5gmMMSuV+gv2JChOa5HW5d2S2Hc2rHbCACqiseRnD0EtH8KXn18c1
cFdKHA37CpziHmJkALP6rVsRXg+OvaqtMZH1MHOa/yEMVSeVzvJlVBDKQlgSnHa7
YxiT5OTt3NliCVS59s4rIrajFB0T6XeJjcbroNmynsZRZxulsadzIXsYUKxeRx36
OxjwdBfbYhHQiSqNyGYWteZ40qutAMKdiKovqKvtLbZ1zhes9kqXtexU69xKZXFC
LiLdvFY7h0f5RRYR7EKBDwd9DWHfEhvwQxkG9+i1Sgsimknjheh1WMy6ZvsHI5dW
2YrvT1MaHPYjtBdQO8mFRzKo8tld7O/4hB55X+MboVYwLPJRrCSTeSNYCelgeECy
OPTq8fLktxDeroG5J+BZe9sHbTbtj61jg1IWLW0l2m4OsU6/SY9TPqdg9SaN/VJn
j0cjwc6PAmAIQVZFidbIlfd6eGe33kny4UMWOyr3CKjihW9O4EbYqywngpZenqi0
O85mbA/sizpXifERpV/CR+3QhPtxF9T9boT0zAlNsq6VTLe07sekWUwg+SQILXqL
bH4GBns89egbbKDs8KoNm8vq+asZxJNNAnN24tG7ld53rI/kc6ynHUoClP3CXeAS
2H36CUJ1EK8DbAL4QiI/DR92uzyFKMahy9y55Ka29jgYiS4msvbSsMrDW4N+J7uJ
TwyTDudXCFMw3l/+QQZ+UV7lxuZ/9gdmdCvJmZgu1Qb2S8avH1dNeA34rNpoHksG
kMJ1RgitBfx3U62PTZC8PPOWTIKh8kCPMHBPeJb6/W9o7flfZgT5g3w7TvE4x46R
JtUS4E7HJBv/uhB4gnbfO6KkjxwT6acnbNDgQVKiJYLrDhbd655ljvgWhtR4/Uy3
pO3tSHfExPINg5FrStmbdKCuEiGnXDucJuQKIY1syNGZbBuLl/D3RDvrx+kuPVAW
3bCH8AwzwARPl+ll5xF6qAVMyJfVIDqwN7jkQUZvJG20dj+EtfUgtbsjBXztnF2q
jMJiakd+yNR25zM61uqXvmSN1Y3cFYEwNEEWljTRCQIMKb+v38SjifAIwEYUSqUL
mT71qBs0sKqvhnTjCC4oweQC0P3RvS9r3pn8df+QEC1jfwztUn15yLnVzf+TtOoH
El50aGIB15Ud929VdOzv4PoK+Z8EnQZGZsLPRFT4/kMvHpiUA8GtW5veJ+Gpf3SP
zmSHgtJ/dysepp4eILx76ooM0PzVlTXemLnfmqzs4R9xlUddmgJjfzObK89z9cWM
NypME8Ifg9cDIpNmzLWFMCXGLKaDsQtCy0vKua77YO0Q9qI5RjH5E1e+BfDQMbJk
4W7uqoLrETxmQ/sC6cyxy8S35nbNg7/qCFwHmQNjfotHFDyf9cqQasTLB0D7epy5
QVZMXPdpCs32fP3kmipEJZDG3zkip8f2IL1SdbQhDwuyHTiJyay5bezLDJykX6uL
IXKxDF3U5f4w1xGDLua8i8NNlRs8t7ftda/UYzOmSov2LCpDXEKFG6KX20lvrh2d
RshWGQu0IbWB3o3vuKEjf+Rh9Kp060kKHiQVQ/B8Ujzv9rEKgLHRjkQTLB6w1hy4
gQjKlaoQjyG0X/jAbRTvTZqQi+noQS/LZsnW/I0BshLPBbhrGkm6jOdUW04pYSMh
DL4PB2EQTI139w81mEjCHn9qwDYNa6c57pfc8tCOxgi1gyARyqIKdgA4tpQYPwYC
wuSjsDbADf4Ch6TNeGv1y/jXXWx52+ERYcDxlJ5rBccWf/+XU49aD2Yp9cJzP7UN
rWwwTA2mqJI8UylBbeAqQ4qrKlxWBPqW3w6FtYQN/5Hc5iqoB4mYwRAn2SY5aLum
Q/rmqK1MB5AZSU45huQjDCm5L3MhRprUm54YflkYD1lMeQ9dUILT0U4nrJkC4LjY
lOQODcNgUKh6CADKP6+E5yhCruCC+MWsY67ZeM45Xsb5Yg5WBC9shCl75RtKW/aa
zwc7pC0TBCcgTBHvKSXNboET+TQaen30A6LT659JMPzNUt8ld8yQZ9aWLxqxG4om
Kup0GemJrJkhczqd5Wkb7okdottOOMj5AtUEz82BuQXFhvq9Z/TGoJcy3tHEOpyF
OfYRFF0mHjlOimFZ6bvnLEF6Bn5iK/UWDVcm/GwOm6nqzskNUoaPk6QONlJfH3Xu
I6a1RKg/2etgTeZT0hRXgHnJz5IFTqBEz9MfjPlOi8ngN6keMxhv2tViqAI8XGUa
1hDpdaYc3teL/NZc4jymJE3Y+gKcH7ua4qO604zPM67Nigpjp+Uw4YXFknBuGbfM
321xBsBMiTw43lz3hQSit8/lFTqThe9OLl3qjstZbH7lQEA2jA9p1qd+i4xmLzWb
BDUw3lkP8bOs7/I6xNrL28Wjzh9ilZaMhGIojwsWEQCGJtbLWR/rkY+06p5+blvW
YmOFkWjtUEFyJhnbds90MMI340T1HC1dOWx9wzP0idJI6iEtfJGDm59WIOy+O5/4
JatYo2My8UIEBLNIkOPdryDCqzLW1qoz/lGrHrS6PDSs9UHZbh36LOHnN1DdY4ur
IvIp+3TNN6GMYXokieXlKeFF77BG6DMwB3iXUT0yBqRWp20Vlq9o2pctZcRsV5NQ
EDaQT/S0zlc1vOAIJB4D3pv75ztiJWOunWuj29CjbtZBNKDCavGWnIkZYoFb7c+8
/Lv7L8sljlgBaApX1OYKzN6sffpPpTy8l1UBMGO2dLO7aRqRhMlhM0NfH63mjdJw
nXLIrjRmorsLhh2hcQJbsgwcuQAHIWREtiwxrOseD+GJIMLfkRg8NavypkYASEjg
3eSm3X9wURI51VtBmOFHDHbQIcOsVVE5aeqLQSImjQlM2e9MqCYnpnR8gPDLYIf6
xvcZgctqVuvrBRBX5m+A9wlfYbQc1kNyoTvCh7kLXTDHgHMkwOogOIcP2T5zf4+W
IJR6nj73Nm5VmX0HU7grxrZ+AbopRGdkduxxgChd2PiTRlatUL93twzQk7YXlFXF
vh3ica3VeOl8jCznoFzrBJpnuX793HXI8DxVpMZu6xLMM/7Njol/wlScy/g6KiTQ
S45xyViC2RklJXMpxSC1pSGTaPWXlIOFjlD5DKKwK2J4HVa67JrA+zliRJWXWDav
Os76zbu5r1SZa9e3g99Jn7yvVRxgneA+2fCNzy+3o8KL80aYKT7IyaFIIjLouHv0
buLqe6Hw7Fso1QEKi/uS7s8NxKXTRlHFiT2DmOT1oydfR/7knf7QZubWPhY9BON5
/qz892pEueXLylVx1t+7y2VaLljA75+6bpTWvp+uHLyj/9KfPUKFlUoxXZuZy3CV
fmX1v+CgpHjBQRxGncRiSjzdWKtF1QtiOgaC+Hw05mYJ1WszllSNSsd40RivGrX8
2hysiQR/lzDT5QQUWg70DQkyB8jK34ch460Aqc1oQQnasRJxkB99h+j4C4Tn6sD6
e7zG3UF6XeBG2TqOMg1V7dtIsh2Usuj2yNQGC+Hu/MJAEcgKM99Ys077Bl47vcFj
J5RqIZmaHWbn3Gp2Dm0pYF+GBWO2qtp7q5qOtZRQw+RSgiXkDa9txgrzSWzijqOC
hm8QgBoEZIAiwIJoToypP7guetfxCNPAn3CgvPz80gqx+/w5F6W8ONwN7q0PR2PX
nTNU1DniqjDQXpneVnKTmB5m8O5nZc8xxAEMM1mTeTCmmPYdiexETdIzgnbOjImQ
IifaeO7BLhYXluGDxKJj0nVmrn/q8i/48ka5Z+vuTZTG57X3v1T05d/zhgvSdPOM
EHiJ8aWOIa/l34roBp/9BY/hVpYOB0N7Ui5zDdbWnBI+2AI8JizxZ2aJZCD+fUnO
bQf2TZedNQWSbOqxvmR0E739OBK/5m3HRzM/MX36fV+emKMuR9jGheo//Xuuxj9X
1Te92MUMM/mgIWR7ZtwHHQ1Gr0WNtt79X+Q3dFIbCqLuEJsVOX2vo8UY2T9HDlro
gzlpXS6NI4BGk3eN3jPoW8opeXuPfeCeiZvmP9AUFpXDV/I59U6tvoriGrJE2U6E
4QnF92M4E28D/LvLce4yuMOJ9EutV6Dkym3FFrsI8HA+XTfKzqO92AQ9Qw4KBOmr
rkz9xyeQJT8wXwSxX7Yv7fSW+YNgWvFw6J+V+oizZuKvZKeO/0KCaC5ODbIpz/Sb
exbFGYxU44SQLjxsA7kDWRdpi7TBYjrtR2jVqWIkGuU6m6xO9+rSthD7ijOwJPL8
8P2IwuCuhOx6ZZtEHPgFZEAFRlvsCoC8WHwMDeDCvBlSljcHLSAClZlP0TvFtDfv
PGE5qcpJGtm/c21OSFsJbYR6jeONqxu9BYeMldLwh87Y/JJjH7EVXeRn0/9XcHIq
ZhhUVhn5cfIZGDhFA/mr5YdBGZa+W+v1reBFBI9M53/T4LxDsQLqhAFkDyqQHqXK
+GnferkazW0ZzyXFClz8Exq7W6aOm2EuTtTdeFKpKuMjlpfUHUtI8eD7EMPcojGx
igKpzex2+o8TXEuUS8D6TxN+kQ/qiml7ejRbTcvQ04ZOM2buW90uOeEseX92iVnW
fcUY2u87fxGbYWoXVd1ryPyE4YkigPLAvZX3uPaSXvpTgA4EzB29OpvJdnfyZbar
NvIf7IMkBFZWmQB8JEEVGXZcvnW4Jdf1Dzc1Fj4RixG/dSiPfK7G4+alQpo5x1he
cm0gKtQWYjTp0pYYu0UcOnICxHdl+Ia2U2yRFkvRokJxYGknmOqAkjwIPCFbGvNt
nL99uh6HAdVWRkmubBxW9C6KD6toNSivdK5ZY/PO7TK/6atb2PfK5p/ENf5X2ykY
eYzGT/RxQjr+N/I+sFK2FYnvXg4P/MPcZjQiN1zeC6XLXi4DKydOX5xz8aAonMV7
6X6eaM0Arz0FZDBhZ44Zj6LP/9w7fvT9kDwGnPy1Htmz742SP/QZgWcMfc8bX96+
EmgJyQmrq2VA3a5yikCni3rE91JR3WwRswoShLrZLDja017aUa3I/MCw/E2bMLAS
PVvsTA3Jq0wrySpBEzlaF2yBybMmtrCfkZX7p3umIcFg6GdgcTZPkujWXU21iXy/
qyWnrhpg1OZv7lgH6Ewle6X0mTk1MRB1rVPdCbiXOLu2kNHAvGSX8a9h4XZwk4yX
cO45yycHmSm8Ufd/ZWrH+hgX1W6WwwtIY6G4QGa2tUw4CcH/uemP4I756rUTzQgF
bBCPGeyfSnmyp4U2OwYCBv7MAcgys8TMJTHofAW0TsGijpQPEjnYanVmCy2MWW/d
N+YrwMoY9iijK5EvufDzasyYPLaGdGmckRC+adoIlykzxTmHrt9QS8BPJ9tqWQin
g3/q3D8CoFQH9PQi/R0O412Lndkpus7YdhdIxXfG+opS/6+Bgs56VOTwx/gQ7n2o
Qnn2vRaIv4dc6kIa6JGWebo6+ZUaadw+w6cwVkS4gSZE3BNnyaj6qzqVpGIhhOY9
VByt0Y4oF6vJ+y5dWLAcZNiqyrvozlO7/KHQSlXIOumQfGdCl5Db99Xh63siAhw1
uGrWc+xFdYRbH74gJefCBEc1IAjRKamQ4L2wh0AkPfAwdhEUAHWXwVRps/5jvayE
AIINq0gpasS7bTdl86m5czDELmPi8megZ+sUqU1sJzOoR6T4XDhRT0pox9t8CvIg
Qwj/FYHPJMfTVRPhAPtUQ/dSHcC/6KRQuiC3h/UWKwt2oT1VwguG6p2IyO3/6Hvd
aZj+YMpPjU1AI8JGY6Crjmvpz/GVZopbtOfM3nZjNLdvNi+F3oh0mv6W0qTR1Owg
8rG1MMMGPv4779azP18vV+YqXWCVk5bmbi7vtSFW4VpaWcVHUaCFD7UElNcrRfOc
vPusOYOI7pC6eboAn5YAv2AGdFcTPcodhPObJkzpyk+Lf7Gja4omwir4UCigK9sI
lS2/tmyB+kWKIFv2eOhEN4W4hqwWGvIvRdTUu8SEPbejYgrMmhDJRzfjDQTsI6F/
U0+yZV8FrRKH4IRTnYoexW31Y1ZuzJ3L+QHI8h14aEJPzYj9ZdXR5Gffpv0CfLBl
SRRMFCnItaiVXE9cTXnk9YqmTiDiobtCyCJevkoDpsLRSGbAxVWQz91ay0pFxWYW
HtAFDvxKIUefmhIofI4muwTfOdQwLyN+ck3eOmtXk3inlBMYk55c1FA5PuPDLtP8
WVT3hm6Pb8fNfgrlxXFrpL1dAa23zUdQz6yyWZIPxAdarhqtlfDEIeNwIuJKYVwz
9sVkgE+TRgzQARuLj0pulXTdQKoxcDmX5O5VrE6I0er9WV0ongMrlLzaoo+jmHoP
H7GfttUZh4I9NvOjKdDiB3pUA2zVatRMnb8oqWjfJCiJhFKkEdD0TAavRCtinBw0
CAxSj6eHyhTZOae8uDCbXkcXwsohLbZlDTnVCmcw3rrOdltppFjrkBjeSl21KJ2v
y5nEb90JJdgaCMOPDSqg6OrrOR/PV96pdt31RgV6liMbhNOw9cTXfIo1Wwb+h9mM
OgsWE1fiugtE8ctYhR0RitItJvm9elFapZev4C5AbHX2hl3+tN7LuzBAvxDswSL2
SFnErQhSMJnTKo/bgbbBXH2K0HgLO0MehF0k2oWG3gOu8NJNyTktqaI6DDOeTeoI
5CQlvV39SmVyRKxXQDL8cIwzYWuhD0GGQSTkuXE8YHmUWR0/YaD9NV4oayn1sIi0
Ive4yI3mnzxL5Iu3XxMEkwbrZnpG7rx7tFSIMCNgklJFwHMrL5fRMB0z+xcieGiD
DMCZdjC4oXPecYDVeB2s+hkmA0TbCupyBqEKvadwjR8oi3TcfVxNL8H8Ynkqr/gh
Mr+Oqm4JhW/+cOiShP+u2ofDmVOaFy/kbSKqvFvN2nqaoSrKItcPJfgwtQoQjGYr
zdYv5BdHAEA51kc4ayWqJHkoQfyPJ11F5F62huZkBKX5d8jViEopAa2Ag8m/VyyG
+Qmd9kioe7rHADWn6BslT9uY1A5vc7Lfr47ZMnbM+gsDFOqgzWtuKooCVcjdB2mX
V8RPv21Il0CZN5O8koFvsWjY+P8Gfq/Pbg+fEPydEKw3Gy/GFqAHkhO3Z7oqZnQC
63ibkQk3dmYCFcgBAzQQA9c0Mxq8fgo2tyc8GEkVhQuL0ltuTSyMaWchA+4/8x3E
rLByUv8YX9t+Pz1pV+Ru3vZYIue0aIKRcKgzNNgsIS8TcyuEfRd/trMNjxbnW5qH
vjI3Bt/FWeAODMWj29iFR96T7RLfQnaE8q0YAratfJ3Dj/cLoCGTGBIpyMszTY2U
MWWRGxgbYkD8UWpchY/bCZOjkbp8fheolmlnaJVO1G+x9Gh28q2HB9aiYs3aQOGx
AOYoAbzEtukobJ3cTGeVpUuBKeAj3/+FIz7NZOrieMUDuIkZESy+cNIeWJYE2KqK
jwN9oTYt5CZQ9CNFAMyC4qhjHDaI6fyNuIJYUV69NbSM0Lpzvb/aSBFesMcbMHJt
L6xjtE+SH36nsf5j0vXsKr6ORf/JvcqT/ge7DZRwstVZE71aMIkT/i4uWXuJQdPO
fMXcLMo417dORcVeMmtqOX2+zogcchhy5cfTZ8HsG7oPIqE/oXM+HEfmeJsKHa4V
YukuwMvAJv3QzWGTGtMSf7upmKip5A53uxhNgk99YDUbNYc5QFkeyVua5R/sAe0G
Yo1o0LeaPzEJ0bP2DSw3IQ/z7b17wxfv9FNK6PohKmz8PtQQa2cHb38Cr7VGlbna
BV/DNPEnN1juSZhKVM2DwB8+5QxGaA2UY1NfOTIzur/jXi9xEwHgavUd20UtIn/e
rtNW5ExFQLFybj+E1JMkZRhd0j83VA8+dM9FMox0XwX7iWbFQngdJD5JjB5WOg6+
7sPNt3U7Y74Sb34HEikeVwwMwMafabP5dHUIPdBr3m2MPvyIH75EnHPK5R0dzroz
K2M+oDncg6p26QRSCk4KqCTAnWP5WvrOpaBXmL/RH55tw1fr+Y0qHgZQx56nMRv8
aTgNkDe1fyxCz8c8TpJI8CtHzmA6pGwpyKbv51blEg1UOoaHhZfnUbtVlCrYdeai
g9pJotJyi2KeMzl1PoFy6PBYJAuRkF3J42plwZuuCve1bzNDm5sLGeDk6pA4xZqS
iwW69qhAN3a06uoOg7uy0q6+Gr9xDjfgjaTh7THlDy/ynMYJhqb2UkqhPTuyWmIO
p7dzzaQMxjlXOOJzjhoW3ATAxcVjscubbdKkbFoxUA3SZGF/+LKJuMbduGRyu6AQ
QR8U8aVoPNpYkFc7xEcQWqXoAs5Q3nXF9C2IMQOuxbd9/qKiLkNED60eiNuF2M9x
zrYpvyjWtZRejHDiQAF7+3PxXDYSefMVdMt42Nsw0WevRIoG2gf4iFSavB5c52TS
VxZDfkX+TRqXkweiKYUH5YOjHRCVCmFJsuY014+Xqdl8kygmAj5NvwB2p5jZ9tk3
Suf5JW2QC6io9rBVZn9r/vg2FeLbCzzWysaPHfn9XjC2bqxLWgBp7qN+4YbRxOsz
jiPSBMNTOcxMDHJw5Argc2s1lcSCkE1cUwNlWU8NsQyLfGdTQqSTsJNgx308R4+R
gxNWA6wVE3Z3McSQRtB32DYG32w3dYPOemWpKMJPJ7XtPQIclonUIrWAw4aMl1gU
yDO7HMo7FxFQzv/B+SiGBc6s2kC7+ITebe0xnLCqof1wMAW79gzDErgyltVU/69p
w5Juaz1QTjGjTMQa4PqBj8Tn3ZhM4rKgdElnp58SFrBcccZxbDbT7XKCsXaVWKld
HTzw66N58DnIcCZsCKdCSvJFBH4qKXuQTOpeEIQrzVOMbo1Va0nctGx6icvv8o5B
2zAoNaJmlXNxqxzRySQHanzS/UiflRyGN73if0GG5Td8MJRV2xGX/gR0nxJ/YTfF
fCP0rK3kz6cs6TbRUJVHigR9QQE+stDQrYRXiBkAIfxMg/ZCnzipmh749mGf/CFm
TzX8q52AOmYmmIiqwh+3iDClbTAiBUoywfylPQ4sYpSfXj4Q7Vb6FyuhTfqBdkWm
P/E84ojrgRs/qh4owXG5lE/Gj7ZzFGKD5QqOg43RpEMLQJ/HMTIhLIebX0Vbvpo0
nC4UiFqn4zZfQwsEETzTjFWQS+yV82Tq245eZOoRKGFF2y+xFbPpb6Dbf9OxiyhS
kwDx0kUosjzGxlajfehIIU9bcn43XXu3Vp75VLFeLOmuqBG+nxPdLTHlxmtJpKIp
f22akSatGe2XYMaCYknocrADrt8dpeopTcGY/GZEMm6xIHerQWt1LTS4jDRNG3tJ
qRtUm5fHv94BBv7hczVh+CwIB3LgtiI5SbnT3KPuQfbHgOrQMCiiz0izX+Wjktwa
+T5vgFbd+MhjnB5KY5E27SYidEZ7589oWHR/rigO6B6ojGJEa/nCismWSQooFqed
boi/hcDczygzKesr15UZs4J0FhQd5WUpXCwYOHxk6DqofxrJHzgbYzTCizH70vOP
jcTvp73EezaNGbP6QMAs9HZ4JTatxdwWj3m6XVHRi1CDP9wZ861pAOSxZPRsA3X3
CTaGls4915WdeKMST4bNrJok47Dj4WHrjeySIwQ7KVMS/m4LSr+MMqyv22IZPGgC
dtXp0FDpyjw/tIMh+nN3qw7ivDdAn9lKj/OMvf7wQaUJM+JfUoW1brlSFXS653sp
aqcJLQpX5X+N4ZZCdW4iy2MjPW7yb+RrFqVhppQJzfTV3S29mf3+o2pH0v0oK5Hu
7ygJ8QguxtruLUvzKrzHfhDeLyEbdTytkCOcBHWCFmvf8IbjzZZVKcqlEDdAF8qH
FzxKHTRq4GX0wYr70Wv7W1VoKTsex1XewehVUedZM9gnoWjr3Ov4Tcsl9Q8EwdWd
cbdi0ttPcepsvNne+EJvtNHFlxjuYshmPeVE8dVcjlpefYcNxTH3e+cUX8CypqbS
f1lLurtXikQY1KPpMu8GlZS8+FIJOxrSvNrvNLrKi8Ae3e9bOb9GnxN5CPTqs4nV
HmT0q5lZLIeuMDjeoQUgrC2KA/r8L7bzeWtMmr+mwhRf0AJ9hk58RSFMDREYO37K
9FPQRgxcdxzKqWAgRncDMIakTQH+9jlGw12v1YrL8wlkWpOmAFb0GHHJlUOzjH0e
MDdP0KovB4mOJUQ9/fggFFaXhSd/q0Dpy5+qgNDxwAI15Li7+ySTL6WUg8jvHPVw
0fOTLcq07L4RiqxAiGuKN7I5+xmk3BxoXNd6btTMjjN99raCjgUJOFr5abrlRQux
iy4qGyIO32XxnIrke8Tw0CVJXbVXHkk07oHEkMYxeBC/B32ltWaWlLd/pm9IqXvu
nMStQnsUeRYtDc2OCTItxFNy9KrRJkfGqVAR8PrekPATSiVH/Ofv+btXfvmhd8OV
vPSYUF7pfqwk4unWQpYjk8zfU53Dr8mNIrfOQP4WQfjVtl6U/2hcG+bC2zjnvjTH
n+ldBC/1LDfhcvZvrd1D6uiJk/rv95PTvaHvQoixg8lT6UIO/DPpYB3TCUV/QG0B
70rGi+7TlnNCa07hbWQyHBqgzClHBGhvmVnt6Q3mwxg1c7p7QZ3yE7fSMxeJ9TIa
H7A10vnU4LoJorJadBfbDlIP0xL8V54ZVw786bZlya6mIrWpxRLVmXX8NB4xmj1K
5ogw8Jg7VQsNUTiTyCtH6nw+WjdrBYPYpeSf50Wt1CHhoa9vA5AwYEMfj3Vi4T28
fpQ7Zn6E7sk+mdQym7bunyafN1207KchjMYMHLTwEPsFbU5GwF2ZD2WGoPPgqbI9
y7JpkVEWSYDoyO26+esL+XaX0/42VZaXGDtacyTSveZbDox59Tito0bMZudx9H3B
nAAmSQ0F6i31xO5n4lENMTdoZS2hqQLWfD+wXZK9sGzHGK/6km3PeMqEZBSni9e4
hFaAj1v3A90Whg5/gg29o3z8UWVwR5MFmZ88CfDd/dte1DFvEyqWF4IHY182tN1R
aUi4xyP9r+t8Etnvk4UVhs/5QwL2Tw/DyDOi11s1CVC1CVRjyny4tproBCQJmYBe
JMPx419LHRt1PVuaOSY71tptfatFvcLd9HmjuKcshwS3br4FDjVCv/+25DpQ5xAF
rt40vhhTTeEbJcUME5qzyysKsW8Dg5NmBc50spZF3ueJ1qCAA4iAwMCzFws+phEO
w01n9y8+BUVEGGoC7hvAKhZ3KlndJ05OpZJtAD49IdOQxvxsNXuj1vEXiEsDhdLp
RGUvI1tEIg//gOFf48qkMV5GhyWwT4J5dUf22FGV9t26kS8Nx/2rYV1Xi+PFzz0w
PbV10GbRIyTPoKxmtwwnas5wzTgoAboFFiRnC0PTn4XGP5wRSQ6S3mF588zIqtSk
3HtviL/ZoMFAbaTRU80gpzuC7YIgr6QsPEjyYg/0puFslHQV6OjtruG8tHXCrWoM
QojgLCeUbVRH73DQ/NYsXmqy7qmszoTqjQ8zIENKyqLF9is1VBtYAlv/VR5HfW9g
IiuJPWBLL4mlRofYSy8jR1bSa2TwgBg0tu3TaJl3AvX4RU2iYJ558bkCUDuO8w/X
EOv+Uxq4cFP80o6VZpts6ACGEcG9FozXf9t5OZnlA247nlfA9Gq8nXJSrk1LZqFc
Q4ZvpWm3THVDbamDgLaOL3Gp8Ro8Wl1NC7kMmP7y6xy+UOKhErtB8bUSYBAvxDlC
C1I+GprbdwjkGolCa5A+4Coe2Sbg/Zz2jOUyK9oBv0L71A+70FoV84i1UKXmpcak
p6FZ9B1PoqZ0DuvtaAzDNChUMvMXapzzqsHoMXSA7WqjKUD0rz7M4o4G3Soi9ULw
/34bNIR+mi+qwAHa4eVL+OX5IGRnPmUHAKQi197X5CPuPvMhQo6fYcbFkGISaZOy
nMAt6XSknujCzb1ocaCrHdk7ARSWVr4nbrHXeTRDxxaiY5QJytAo4fqqPfwzx2VO
pmL6ouPTw3UXGy4inMje7PhOYtgn5TfytluUEjzrRKJHRjBlM0W8D0a3M3xo55TE
7tuX0YgTNvdHlIj37Trh3iwJFuyaGxi7K/SXHPNpc1dzHHmOUirhRJdlOfTl6s5+
ziDxFVDFXRDb8NnMejmF4ny+RWV3EjxJFWANvABMIgG7jADn2JhB1GiNnSzBHrfL
5kHYTXxVHZtOSG7E7jFbtqKZg522VrMRL/zjkGQVnqc74T32BzE52CpEIwE4OcHL
XyVmp96gSFzOFI3g+K9RzEQDTAiovro5p+eWLhFd9qzz/xxSze/QsOidpgXWu7cG
I0Xmw9Dfnx+FCe4UHKrEtf7ZE7fKVjy+WbpG0NWZz6EZO+DQ1mQ0dA0vvomPMt+Q
WMKlMJS+Ucd9bXmAsvh0BbGGzb597KVQjRc+6amMMgIaI88ZqA3pEKOAULWCCXsY
sBzejh0+oTaWaGz1PUoGtafwHZkl1dzUxa0EmIAXSTZkBcJ8HQKL+5QVcgxwcFtJ
w19JuVkimX74TvRaRssWBLoIJJkPLfz+1uKF4oL0U5W0W6Id2dw25ZC9KUwU1fKP
UYtDwEk9RKceajFbUrMLgQRfxOwDHO/cAMA9Moj4nGxWjzDwO27AxQrA1GID7GnC
NO2Pa4qZSvhBdwhO1d2mC//8Hv8lElafMIZ2WnIN4aC+3eKSpWkRNoimIxefHOed
ELuyodPWGoGCMxGMSVjYaDhO7ydmjwmQv+fXqgmkmEwRIvRNdfDt2yfznV2vHG7x
Knc021KXTzaCQa9dbO3mQUl7CIjPEMuC+6u3Mk9ZJpgmm/XsoIlOh6DCi5nIw5IN
m7SY2E0a25zqQsOAsUhH79SudVAtPW/j6cpYSDo6M8vzPL/NwxHSHOBHMsnMVMK4
i7KkDsSAE+umyIoCBUWJ2AfMx2yEtBogQUm7a2ASBslRusTM8+ngsAXN4T2LR3FS
o6qrcnYafQwXdEOgHd9s3OFWVI5Te909UlezRdlM74OPVBHAFVGUsxlrBXmwQQ6A
67Gfus8PtqmKVYyXedSY+p8bBZpxuWYwt6rSJFa3CTCmtEAf2FY/HxWUjO0kBqD7
amHZOPoKU3nKc0oSengRjJhM0UC1WR7d/mgrmm8T7lu3UOlUUwl49z9OGhyk1FXY
qJSNk65zBX9cde4WGTf5fFnjPWnLvv6PtRJey9FMKOE+Xf98xZQt3UYVhtUnChVZ
pPxIov5NoQGqmg6b3IIVkmvsJOKZ5/w9O4MXU+W/HS4rwQPizUUXseX++zh+Kixo
gGaYAKdRbyL5GXIErHLGtv2O584qFz/k9KB3KjuorVNaqmyi29/BI6SmPGFBYyYJ
vg/1NhBAKQhBOymS3tL61x4+ethpVU6oXjbrftZEgGbsiqHYa7GVQJph+C7Ji/yX
PPWvJTsk+JqMt88mNuMT3pbicflDJgfN4F4KmiGSqk7wr6yw6OAgsram0uUmqWXk
KrDTHhSNKx/uWWwKglNAEZhiVErvnCS3DoX0vzTUQYGg+8kLT68SkpuQfPjN+6bU
iWjsfTAkOhI5VurRZvIUKPHGJtLWM8idE4QgtIsL/2laE+s2NvPeQoLw9GlXV49C
RcnnQMgFph+WKHo5Voz4zqCRD2hOT/c2tm5pnapxv4qyXsfhhNQUR8faSVhVK6ba
iWbgfTZQF906DHfj1cQ2+dcWxg6lgibhpwy/Qm0McTTXqTB8jZUQoQ2LFj1HpXuy
aPXYr9WZ0hYCAebDKQw0HboympzLKM0LiXh9/iusBg/MQ0wXOY6Rp2v5oM6SbVKq
IrWwOtch+3FRw0V2NM0Rrw0rPDo3//AXlL9LlZH1Cq6skgtIqVYvibxRyV5uobf9
0RWXUZA+8PZ8txI6bw7apZFGCRbXhrAkccHYOGPMcOopqzpaj8gPsHMbHX3RA7aW
JUxicjIoObTCTyRSynmlWqVB4sGn8/A+oMOXV2EiJ+nT1hLShWkUgTDrIGNUJUpv
4MrPvatem2815teTE1NRYJFE0jMq5RFk5XUo1YR9YiXY8mGO9zp+W/XfvjHqkNZ/
sxsd9MXg9pql7/BJkWTgL3jHa7C5lZNkyWXCdWg96Yp7Y4+Ofm7pOdlKtkqj3RBj
gamRkQDXIAqo+gKas/ITXe8kGSifb6DEQ3wdJYpolh/pF1+eHvco/4igjratPj5f
Qm2A7V3q/WT9Or2dDcZa5n9mgreGE7lg8n6zx/GA1EFI+SZYNqlI6o80ckJpgJG+
EckPRQfju3DlvtmbA3oF5hNgWth3EAmr28Rj88K196+h1SgV0Nb2eYxYG5oPThzu
g1CQJwA8Fz/tDOKp6Av9nWFqBTBjXl4k2JaEreqK/9jDz3yava1ILg3emIYathbw
hbu1cM/6hySPmOD1O59lN+uKfny+BgUnHoayvZz25jEyDOzf8YJtMUFGxygwYoqS
UFNJCvbaPTkTfGvQU2k0RBKDoHJmcXNbq9+aEEJJeJ526DHn2PWGIRQ0bJzQMWtl
pR130sQhk6wdHTSBe8A0YICxYTKMZzKfNcdSVBLpi2pv7yrM9kWq96rrIS64v2Ws
u+rf6apfl8b7p31lqokp5J07RCO4oOFrFf/EzhSs3LNV/rjmLPikcvhHwKVnIObv
MCIXfqckOyKUfVSKjO3kliGEoMqFm65K4fUfE2XplcP4NC7MXOXfpok1ZuFWFkQ+
BPRcn2DHo4diiWSoifFyeFoEfLbv9KRhYGAoZQD5oTAXTgCTd43uITIxlpyCsTNM
y7hgPZA4hBexQQA8EmErsNcS7H1dY+A81v/V01o19E/bIRd9W1Xvj573Nq2aC9UQ
RYYjk5/jAS93I/ZjZEDZHZaKQOK9lMhcW6caDh2E5z5hXPL4d/JTJnbEb5X+VM2u
NgiCySOeIP6PqdBr0DhqQI/HrCVk53kauDX9R0lNfUlxbJaHcX/+ttZvEznk0gzi
+Lq09KMLtZ4uS0+IUgEAGvZMlfKVLVbZJhHedK1rWjC58Beq3NGxaS4oWvL5pIm0
L+wA0x2ldffCjBdlBo/ECOifb/GZyyuHi5NeBOXCiRo9fcyCRNQ6eERLXYTQFksE
pEWbhWfgiRIbha3UFP6L+z5QTmBo0rdL8eGrxJK9Nhy1ACTTVQXKULtUWuQUe68d
6LuTewcD9J5XrCophQUQhyhQuUnj2/UiCXO5qp+ZFuPq0Ewk5RZcFGHQPCgzw5P0
39YDhldGWufvpKUTXN1m8rWifbxmrQlcStuIYkgvHiIFBWhDx3ASGiEqwl1T+Mob
fSwgNDvI9m1bHcEkZW1MJzz8jf2xdFxv/I9Cx1y3REDSF98Ew1m6KhJ+3JacsDUD
+wyAhAdBOBkx8Q5dv+m1HHOzB9zDfH60SHgdu4U9puRCAWF24D28d+hxvzvI/aLL
i9R1ebWQqgrAb5ZwiJlNpdY3fgrdurzGiMtHnAserS038muUUdRXVDKlH/nVSOap
F12lP2eTeoqX5mAy7I+nIPKH8o0SbAfWEsv68PKt7NIiTfYgfLigqKEWC3mk99nF
vNgypz2M+njPvq67zEyBj1ZBmrNzTsCYeQG/YDIu+kpE1vVNIZnT9UX5J2LUmVFG
R35txfc4qchnkXO1aT83SD8kJhqiIbDJLMzURSeT04aS8FMIRYUH3kY0uNdjeLlO
0YY0b9wc7ChjZ8e9GYXDFLiatswOwEbm/DoRIcpuyltEabLcVckM8WEo1vtX+qoO
baHiJ5LxZdrhBedZKTETVYnB5zTYRlFJrMFgKCwX0n5S0D4m+0qiHA4yQGGfiVTe
6j5xOWauxnYMx6lBgwJ7gtK5Rt/XbTzqnKG1felR1+It2oaneQaQ2R44cTcvCBgL
3iUPZxHGo2YF9dQGNjadIDrVqa8MrWoCfsnaPgFL2PcL+D2FtDBLJzHb8Hhp4I2e
AoV/Xieybc7oTq7lpjTF3ic7Bu8bRzocO0EtykvqUvsGDip7cXdam+cFhNqzYT1U
Ipd2BtF4sBz03vP11T6N2ZcV+DKMM+TMjhSpG5otWaV+1ACqenu9VAX98mek0nxg
Cgf0qA9g0i28ZQmJl68gkz/gBI1MCWrXhjBSypBSyDUeLaPu0Pq38QCN5USoJi6R
KyBF2B0O7UoicgoDkHWDHXkydRsN4gpeihdrfu0WyZ8Rx3PnHf6zAyfEtsLX5G8I
2WDdt9xydzNzqqgJQdFAj2uA9WcKGo7TYz5KcbCkaSt/o0WRBg1DwUuawYJ9btJb
Jk7bjKW2hxag2Qnl9uoxi5IxKU0WhSwVbGmS7GTlViVWNjIXAKWfnZVZuta4c+uk
IbV2E2uPDtZvo9kX6KNkC8kKHKOXKrQgwFUBQPbA+/gW7YF0DVfvZ8NnnK4uelVU
onz6kRSddCWrU9IPU1DCxGW16GNHLPmHI/VZC55Gjnbv55Eh6pHbL9HiToB6fd7Y
rxpO7k3CCeLqIQ/67wdOxyXsPoK6TR8n54fvA3woWk4rDMEyueXryT1S4gNXHtR5
MjZ9KRU2QL2pe/2RkaYqaGu6ImC3r1KZWztfkm9LqlmG5Bzto2U1wYpL7f1RmNTc
YjDCfiQIcGxURjeXCIa2IAcoGyQ+wyknXPy8mroRA1BSp7vdG+K4z+2yXDE20Ge9
6KXyMd1WN03dhq3sK/qpoy1C4pSReJhO/aLhHXd3ItOrhJKzXpbU2NoAiYnoPqwX
fZId9I7bxqunQej4TLAvlLLROsTbDe+nJCeJs7oo0IxntFoSqdsxvJJ3qk8vCq3Q
RKVd30wx13BzFQkZRezELGARuomQa+2LKiNmbO+W1gU3NfQjfyj1RKrgwHME/B6s
cACobIodHAEgd1N48uFx68S4q2c3PE3w663LQr0pU6znD8hPPQ4BZB2EtGJYBoFJ
BzCOle6ex1YtHTxTq2WimjHhhrJckptImEB1P4QPoWbbhwBE1WbjacHRl75dfa/c
04uLajanrayKQV2GoG4oOGZ9QPAmz5mJb4139o3LI4DO+VJZtUtfhruHePdWPQxQ
0jogFZT+i8/BMPpy4HX/xe1TPrlTh1OJCpIWIfIttrr1b3Rmx1kxtVKrwCnqR1KJ
pF1NeiOBd4oybC6B5X8dv/Quz308gFDa3esyA7J7xfghwNqiI+q10uwH3Y2TrpWN
Yu1FNC4TSuUlc2rXmQ1BUPlzJLhkj/EWZjH5zpfe8Z3lHZ0h8AWlnhJZR0BggDRp
OMqbGzECVwgK62kS9TfP7tNppN9YWXdQHkAxlBda1HRUdJnPpfaO281sRN/PogMO
2T92/Md1fdMUcvjASZIyqQKvSyq45rQc+/xA4CVMjCztpCW29qq6cxqMq+ZZLrqG
ywXFvg5GHdrOYg8lE2zpBGS/w/pkA8qTKpCucAJg9qa7BuHRI6HimuNMz+nLRb6W
7FhkH0tb76A6GUEZi+9W1iq1zfRDJDhOmRaHLkM/4QAjbUBtbxXR4t/QV/hL5/K+
nzwNyCA7INPX1V+yLXsRGItDakJJsF5nPQp7FQsQt7cUiLBAapubH4bGbuFrHrGS
490hnKxt5Pd4nwhXfdyc9abKclEb9Hq19TTWosLep6p7+M8sPLaoJrIScDgn9w17
zcrlIOTL9sPIjo0wZZ3pzD9e82FWjN3/QX32K1Z7VNRDBhciRvcFAXo5wJNXvlz+
Re7hfpIbDQlmXnVee8ikXVNI+0aw2yw9kDqWO4hzTbLkJT4q9RMVP8bzbMT+ho3C
GirRUduRjKxb6YrCzQFTBVbL4FtfnP7bbIOQx3jSsk9QHgSejfZqQ531eWcsfZYw
d0m7HDBwC1hufJ7Ysk0DlRQxvtE1/uAysFqthbMH2nFTkScFpVtPw3i1oppi3ktA
16h4CO+R9yyvAfGbzeQqiesZtC5B+kwnnJenDH9pe7cwe/24JR6Titpoj4uiCBgR
7Jjd9bd3Qjm8XZipMccVBqRYI7j7z0xxlmG606L7dC4fzVHCPFx3pwpRFBnNQ9yM
wEm+bjNR/JmLcteQMrrnRzzsj7TsKONw07EiJf0hyKihjYAMdV+71mJjxStqWAdx
/83krPLFvCjKfmD9IqIe/ZpeqcnfYT9aG+FcUA+V902UoMeW+U7oGUNN5jencZ42
9lpbs2g3ggsyR5TL8KIveamDqmE3QflOjwWwx1gViVImNa8gwQ6VDGX08nUnzZQi
/pXglFtWEYf/wOmU8uQDAXpxHuWR3kdT9jmXQBxnDmMdtxA+n8yvdNxmZT2YBnI7
Ao/21VA8bCVGPctbcC8OJiWm0VOXDrWJPkstqt7K5sBa239svgzYUHsomFEBaX6N
Txughsgc5pVz/tofoiWx50s6XizeJpvGy07GdtH7+FZCwlrdjz3BBTNaJULtWpVj
HCdxGsV02vpo1ScesV4xqW+hSRH95yW+Ew+xJanIKj5H8Obfz5tZA4S+3hH53YSG
wBPYDKd/1Ie0UjlsqLq6hAoGmfst9NnPJMP0FP+rU5OVhW5L2PGF50szJljz16ra
K3lWit2ufiFp2wf37IZAS+mgLkeB8j+K+YsEWSq6Owl70B8Ilko3WuGPkYZopcmM
rGUlpb+2Fln8Oa4ead+r1ilTMmJgRthoD9h/ihY/utqCmd9W4LX/cQQFQH8/ahgr
nkssLHqZ/u3hYcnLeJb0OaGh1TXrFlpSRZvQ4Q3LzBDCT4Vvl2H1WThF8WvvHuG7
lRdmC1kkfiOxTnQAGvwTE8XKCN7VsQZ2Uw7rMomArFXaJQ2JtlnAuGTwHJffYt7p
MVWL2ApVyKZOc4BePj36IKlDk37uiEmDQcZKuw45Bw/qA8/UyDWHYp9YvQnkxNQg
ZYBoY6oT1v+C5jK9Gvfgj2Flw4iVgs1po7+hvmyCHjrszGwUqL2O0/dEMvefygJi
lvK4UtTjHwHIU6Hyx2v4jd2wGcDeCliPN/Up2MWsKe2WjYgp44MUyZVo8vF3JGsY
R3/r9GnOWkTen93nboDyoqHtqiVb2XJZ0c5vqUBHK61Sy1M3DdkjyYpeuaEuCmRX
7CdStYjW7MGcS+TZt9vRu2UwKzNH0HRTCfbdJtshppi5yyPoCEkDygKd/piIFLIV
5XdNFBgiJlCrE5q5DpNIwQ8bzcgrbUAd/sTRFPeVDc8Vm/b3cxMwnE6jCjIJzXrb
PWesPGegwcjG9gzfGjQzgpvhcMY3M/i2xknu0FDpuFeIBFnT9GEfZu+QjYXnkUMm
KyUOUzAyR20fsUevQ27zbsRvuqS572T0mvYoLMgURGdb9u0sqGSguBNaKkOVi5fY
5TEYmogYVEZtgrtVYcxV19xXHxeS3NiQPAJ9oWhGfFuTTjYemOjIfjYmRQ5loigh
AuzWD3lFj1Z/pVLdrdIKobYBxsnl/dl+iQfXXmAKQpNZCE9Sv+COI5em4Xq8Bpya
jmPQtrZhX65PFN/01clzrMWDrrCyqsZzJEOlbheevY6verksp7YA6w7M0L6uNYd4
/UEGUsHzSGlSdw98jbplnczR+nC6A/Kq+WW+6IvZ6TnMPD5LNpsTo9fXfoVKaB7e
1AD9Axxnx4ENCcy1CTtoVQVaHVKpxK1w3iOVAp9gbrcR3tgRcbvf5/DGYdgqKBks
GA7/fsj797SjwzjvH1hgXxlignjFLKbT0F5EB7i4wbZACDnFFQ+hALflh4dMYhUe
XdWcg4mmycgrSwY4RIDx4NRRWtcGpLAjkkoZ3tLedcemLtgBz80yEdrrJEX0MvF+
Ezw4GtOk5MiQvrBP5lRwX/pcl9MT22gXLiooM1MkDOzL78Nz5s49ja52QCIh13IJ
WEhXn3So5VeaLRajoyOwFMAShCX01933Fd3RHx9e/8SM/wSj1f5+hKZTA0BH/KG+
D9wyUQHnqS4KEELx8S8YMLmH3TWBsNupCVcQO4+6jlgojSmaOqg/P1LwIoNwg3JD
e2FyNAUYNKmHiYY9K93SgDuPBrTyOMcipgx5QFwYxFFkgqPHsIjlgSHOXLhxDy3J
FN6U6bq+BHBGc2A0pyMvBRy4lAyuKo3/sJX0ms8bcMiErj4/h4sE990yUdldecPT
SJxASJ9/lAf1wJn/HjfzeHWfG2IwiAuAmC+y46q//435x2P8AQ9y+JpcKEvQpkk2
pN+zQPQE30SpYcqPItp3KxIrx0ywHidSPE99cNrULmNS2mY3zHgU0Amk8YvCA7ZW
NDDYyJDvNG9wTUBVwt093NEHG5PaAcGOdBGQG65jPSozXY7i0epXOwCxAApd+9/d
QneHZPapStnh4YVCxAEvuciqLdSSbKaiKwwwrxtiz2J44cw08GGsCoFaWAp/8Lqk
GOosGFIpnrFgGHdq1Wmp6013iXPQ5EqvtB3u/xGk/JxdvQwQqsOF1PgeVVJlUI9U
YcGEhT3axxAjE0rlhuZOtr9cczmAAwVXSQ1P9ooCS4jLqhTbKUkgLY4oGmcD5DP2
sPvPQAUF2sxTYCVruXQbJQhCoWCZwLNxugTqNIBRltwPz+YePSg0ButnlVdXOBqd
UxdhPD/oQwBQCe4MepxAfrCxf+ayn7ijBMgs4OAiP7NWL1AHpyBVo6rlbSfR0aQP
O+OcQUWsru9GfRJTerEVJqiBG7fCtTHLjZhQn/c/LB5GuU4Bx/4mnfHfng/A5vHx
GRhbNrZkKR0atQ+eQtN4JOeGIkmq1ydACfvYqCm4/YoKgaigJ1zgq6Ein2hkhAt3
kqPZWPUWk1GyUyUfdUJt1J6wzxT8cBY0zUH0n+Vy6oT7rtFlqIyup62S/bHJozfh
+dSykaWxdlJaNsMc5rFLSbL2PjmHtkRYC52hRVkAv6vxaig+Lv6iXh1Z8v6y0SaF
Y+MFdSJm+3+5+3SHbsrSFBddXWy5lih6Oq4r6J3Lsxane8u2BjnYTBAA/4wyEa6l
jiE/REA2p4fnayWn4NmMaN3gzAwkuetCpf6pErUlXnHiBKd3WW+BiFI0IMgwRMo2
Kj0rnSHln0W1sV0rpfxPJliw7nA8Seai5MVUjb1zi3RN5zyUEG1nocse0QOe2iYI
c60QFZcZOa5NGf0shlpvCGYnwWgSQ8+ZyCMhCrlsjxk7oZfdhC4lxqr3Xo+Gz64d
T0c28KMB7hpCmBJhHlRdLAQvMXmV03PVI6UlUab1rCMcd/MSBS+XOz1f12j5l8Jg
mLYZbN9k9O4uSTzGQ1yTA7+UkoctV12IhDlaHEipQrkFJqzRK/4J8Vc2lII6rHkJ
qR6O4ERSJU50xlgS5E1CgU81Oo9RV6qciG+Ugq7msR3TZ5V4vIUPkw6CSeRyqj4m
p3FvnvHWZfrLyM59FD8J23oACu8jTawrEKA89dTfVYyrtbh//BfQBKCWTmhjky1q
4dyjh8EfAoA8DN2nArCmD2RSUYojzi2leNbrJ0p+tzIRbPm8IdLAEP4Ddc3aQlBG
iXArasbugHOtEFZWO6cNM07aZReiNoskzWumm/LDv20O38TouKRm+5TKMER8fTnO
QVcKSsI98kJbfkjo5quDAJh5bpZ2zUiaas4rr1ymET8gB5UiJfD0upkCmg6a7+HD
mBk9DwCwRnX/zj+sbYII62Zhc+xQpKW864EBF1kTYlnpP983G+RUHw0g5F1mDpwL
Zn+FRTbCqQTNz/2kfjVh2s3UUv+Ocf5enK+a7H4kHl92K0XROLf+fUHuOrAVkroL
sf1xls8POWcDw00+aQJHk1nnDKSrsTa/jIsW2WEnH7CSThTXTO229dMhJNS17Mbd
r9DDLXsQovm/M3l9weg7pNeD/eob8ngCgja9ewhVVzwZSQZ6xEEDI5VH7SrJSp24
Txo2F3ELwl/GAFKWtKr7pvnT2c4o/rhT7+V409U0BSwWIqwPUsxwn5YjhRIK99Vw
BpakzhOjyUh1irZh2mpfX00jEzljG38cx3G/2IEgBMy19wj9jWnsOikTBcd2Vu48
pEtN7OLBjwRwgiufmf2F5rIfKQKpFUjU9oCQehlwtxDDxXQeJx1226FFh1fi+o/9
XzfYcHB75N2OKzWA5xEDc8pGPCDd+y3+9Qgsy6rbJOerODhjQU3eIC5/IRxZKtvc
li64YgsCBzYSoSFY+yLsYdP0CsN4JV1SAFzFRa70Pgm8azhYamgmQrtbPH4w7xWw
0pJY+kMY6OvcWZ3Rq3c723H7sAJvoJYNuPkd9hIydn5rrWGeQ+DgSVfg7DE6nSOx
1sQRyYnsAkl3DvHPBbsAlrBBY6oXRzqAPoEGYg0WcGl1Fo5zx9viI/G+c13LLHDV
wuhMhrXEtq+IY7NiA837irmazH2nqdo6HWWkj+V9cgfnPhzMGRsFRKO+TCi2YMk7
jON4rhOAq814muoM3gdKhT2mnoSZIFw62TR5l56K6oK6BtIK/incW/XNIdVyo77f
r81H9KFo2gnjmKlUf85HRwYZr4Xq5L3P1bPqw/v89bR6Veu/UFDpAH/hguHlbNpH
gpoMFxb4shcIOZp2UJPsT4hXTWoyoALQzAZarNB4gmW2jbEs/tyC0hnIf7X1VP2e
2s4ORTohnxxG0dp4cx/Hfb/Z77i1AOCpUDN2kCYab8Gn2QHLJYTZdYGR99ZZM04J
dTi/coN6azPnn41J/IDzBMsJm580ioA5bZ5IGwyOYuKp5KqcRrhnIqqwdnsfvwEO
sqCRpJ2+mkTK3XqRLebUW3mh9V2+icyaL1yBg7hNnESmSnNf/QxXnlZzOPcjxRbk
01v37AkpKLiAxDCDAW/NPZvafyzFcPux5cP0s8Jb/J8osG5D4YUqnpR68y8TkcBm
nrEhmxVfD40ddttSli6OMZGTPmARVZnNsqxK9mEWWslmyOGW22vn7MV6HGJDrYtM
kVRuJ8AZMvCRamwZnXV40Wu8uZapWbirAN8XVQVORdnhbwjIgkyVcqHRSpfHSz3f
820B2Xo6L6b1OQNKycMVxIv5uFb7MhlVobf7/1lgVwhSXwhBRFYZ9FxFhFk/vLMD
M4+EO8RnPlo8eaQbj12o5m5WCHzQavRv4tDZce5XiSwyYgu/fLyPPO3fYTB5wDxG
PlqOwVGP2ZdD5vlI9yZXcxKzHAstwJvF1PXg8+6D6cQlKCz0oul3ZgMRgER35uDF
y5DI0jUuoubDzMfuEwN6aGqlDDS5d0yuNzbLyeE04u6zq42gBAN32cDkZYXG05Rs
F+A6leM6qaTsKRzg3Wkm0lEkHJebiVyCaCcGnESTsLTDrWz35QMWtSjKTo7Nbn7x
R1Q7fwwERFiG0kH3Dg5FB+at5r8wqv0Xh/ldVbSNa0KF0rAxGMsm1HenTZ2zd3i4
gs2F+3Q/5jVag0+nkGhDerrMhfVrvtETLbQyH9QFKO5B58CvHxR9VVYJjnJp8KI3
8OjhHCPYRVYZSvaOWMoiG4pBC/UcQbY05UORshB3hBRbxXRIKA4mY9qXa3OTrr2J
Ce4DnVnVLcozC7mIrBClmQpSZJ7JL2DfmKamL+rsmpN8MzRSEfYvDfDL8vLSoa9O
h7/xUroCNcKdTycY/guhcxCqpluGR9MHeiWFkPiWVuPklwtQXyZLG4O1Do1J1wOh
IQTVzYxk8BtBIm6lDVSKf+RjpwQMUB2w31TogOg5mqF6eq6r2fCKxWdP+ReOtdKi
sjxpBn3z/gR7KvPU7MJXWSC9QaY5MesCl2080no5o9rf3hADwP64DLNEV0+xn5MX
mISM7bVx5FjMXHJg28whvhkjcx1UHk/BeYO8k6acfNPWHTQdCrG4Qu6n561Mf3lg
7DTIzFt7WBiC/KfozoYsfh+lfBhVBsqBZdnGXcxs4quYBH/TSV2dlZ+AhI+0Ay0U
lv6zKZF2yPQowI3i7ONg+40rI2Y7cIcMuVODix7aKmd+MTIduK3eW6t6i3il5SAp
Qd6ZSzI++6MYdpRS0y78OYgYbZIkCu00jN34Ja3wddabkMnE91aTjLITHQ/8C3RJ
9ZjdUf4uP2BAz5+rFs41/w7k4RSBerN3LmzovdEe1/hC0T9wCpYa3t+U3it0hd+a
tUgwe0NATBwF9L7M7dZT7QQcXeOO0fR3P2ZV4+ZOBm0xtxP2tLzD5uXvRqIPYAg9
Zi0aWdR7Bv1pAQT8uu4UzMTTj6gk6HRWYLt4uaTaCzPt+z3Qnh22tQdTdWPGty1X
65oFzhOr5hIEUSZbrKPEzxo+oQDVh0LcIH9DVA6UWEiNe9I49C3PZaK5OxbEC17a
qjOTiJfWk+PTXxegCJFGYqbTCod+imTGwE3Bzza63qXmbQOrW9t7gKJlKqeV6lqw
zReBvWbQs3BwbCb4DjTEEpGMpwjPRhRaeFVohzK8BrZOsOWcRgZWfTkSVNSBjiVx
U1ScMAF0xWv/sySvJvanmgpUHegjm2AgRUm2RRnKl0ghVIuBShbfnva26KAwMBGP
6UYDBhLgaWJDBqlgoMhJWIgaAmQMmNVQk/xzeirpzmfLCOXHwZF4+K6K0JUmgWIg
nw/oPBMdxRBQwv573BVeBR5PF3sL+6CY0Cl+UEC+xu4qEqvQ0C9ZtoO9YVLW9yuu
SALn3PEGw2Yi+xAwqRbobfOiqIDHJFsef0LF9RPQwggTCSehNgRJAnReyxc9Rr/t
T6ROHy01EfaLYx1EEdDZCFbqn4xyKSsDADV/7aTK/CtskAMIEvYbad66qDTnYF0o
4sk0TQBDCWkthmR5otYwWXfHwZ80lnHnpMXhJ51N3gwg8MlhpH2tajPzvU0MOtlu
BPfKLW0B92dX4gxnMTPKA/7/LkakGxJYqI90klXxHcBuZdFCTDdipu2U/vGsoLMO
8X3do9hdQRGs/4vd7AsdZh+5sbYaIhrIB8nfb/v0mR1fD1vkCt6wTh8NOS6W/Mjj
ObW1pDFCPWIN2BP8Y8LyMTc+HMHCVA9XF3HviAicZSSmPiLXWWk9cPVqfvrw41VG
IH4IQiKbH5WnxKuz125oTzgClSmBBkNXNxxpynDRll29QQiNuCj6WmkmI9Id6mAQ
tdwgAd+BgzHbJY75bddRSERJqDzeKh1Qdye10jyIDCtcR+CugEOMS5MamLZ1o9FP
fuJSkW9YQJAzCdAtzQ6uLkMIY7jJwHoBdkVhe1MdDvNSBt3A1+rg6RnSzD19n5vt
EuL+YvQWYcMePi8aXWAwvA2GUtRbOsZE6VWOyWE44DkiPS4H8zm2IpM7cAC68Wu5
7q7WuPOcKAJ1mWvIEvTKMcG1m87zxgLtIe3jEJ+RQHnLDtu/f2JPEB/cmmAhPTeJ
FlpBlCzVM+SmDBvNVGEgwc6lgEHJ1mXsFwmbaSHn3yth/0A9NGFORsRj9+Xa7mlt
i28lVCdCxqWb/+JHZjY/tQ9BG1Riug9KNB9mywHJXZnl6K+1HoluU8Ogslk7/xhe
MKUhCVdEm3GflUes/seOok9GixNV/xKGNA31/l9vfKS2LT++bsOOgcoLnuHk4ROf
QBEqYIIKq2wIYIu1FMtoNiK9eon4EI/5Tvt6n31r0Tbny1p/rOQwXTmayLkSB1ga
j9WoF9A2AS539wzLvVy3aZ6PWyZ/ZaBFqwbl7/aHe2q5qoAsKeUhP4x6/6GfSZTb
q3kbMTM9jpN4XCnRqSMgWQbWPTI4nAkfMGRGf+11V5i341fahNmuAlOr5cm89q52
Yt9bDt0K0EPhkesxRAQyxB2QxEPCL5XSy4CSHzmSyqO7qhJYuyjh/5vvUfVWuX9U
iCXXzSNaRkwLEBpAwydhgQSFhOjI7feNE5xvwMFNkISPL/v+izxZ5Kjos8GIZuXr
HKMma8IMBJ2DVPzsEf9NVyZl1h6SlXVnKtu717eYkXAxZV677ohmXpM29TGNO92T
hv+fAPaKXvB8/0Eyj+OsfBI4wZYGVZT7pjBkPNIdFSfaKPxWrNMfo4JascAaqnep
lFyTLx2hM8Ex6C0zrSf02V4fEyKErYcGuDqfiYcdyK9WRJJXUjRbi6G1pFv6nMX6
si/K+OfeO6BYoRxgMiPm3Q0xd2kOfMdZieMSL3D7eLPnldOObkwZ0NuoHXBl2I+w
7wvZt1If2WrvMao/pnOuPIQ9+5E2iCiNtAHcbzgEdedaevojALBMes/xspevFK7r
BinZWwMDsU3K/ndiQBEaf6QfGKStWsNP8Y1BizvH3lrSSoSlkYr2/2rUvq20emwi
OLcSRnMDO/DBQ49EGKfAmPGC/86qHqYbMbK/+tCpYy/SYhYWao0c3ztf8Zm7Dvu/
lOT7XnLrQo/U5g8ZoWuSarg1BDZKdg0GntoTUo/zOswKIzH1Q2LPBxOtO/veVktU
KOTHvtxG2qn/XYw5uTvMVJrcBuwORk0ILVC1zcZyNNOSLi5tkOR3uMK+iSOmUFIh
JGt3WG+AINPeDz1VTLTb/JxEM/CXYkYX14342a0bTQPycJ0ycG6J8Y/5EvwEawyZ
ycLF3XOK+ORnbm29BvcZoX226/4uBddNl54tT2vzV89SfH9MOMGL2uY0YJ5cL42m
DsjkqBZGbhDxL8LL/zmhjlZRMEZMyJDvhhaSMC84i2UHljANax18hUXG/YpGyfjx
WvxEA0qRoSvwUs3nebRy0FatNGdN5DPqdEu0UrutaPSOTGQUhLJAm1aAxdkjLHji
0/v6/ldjzVu/jVcVYLXwUM4oSCJjRQpbnoYorwlWPE55VaAf1bzxii61qdWlfLcc
CACggp5C5y4FhISnBOg2lr+wL7/ZiNSp8+VnDunM0pXHl9D2YClAb/Nr14cmonSg
DnCDa5qlbpD+PHm8wlMDWbpZXtmZQweym5xpKuAoI1SuQpl/SB5I0RRCevN+BgBo
re8eqrWlbaesmcwCUvLGbJowQImTD/SYp3GHB4eqqn8CA5c926FMQlnzPpfdg4Id
iSQ5L8qHju/N9vFS5a2A/uP89EgGut85QotaPvI6Tn118mTZ/z7xyFK+rbr4MHbe
/WLI3OFz3q6jjGbxv5QKHuIUCPMcsOe6gBb3UTduHl1IeQBg7aCGSh1V6MdHbH2d
UWwtWoHUMOFSZEH/xCp4GX1rMPCJTl7gRi3o5MqEt6OoPz8s/ubrIiuUVo2WpKWE
vW8HuqRXupfgl3dMSIzLKYylvZPVdw+OzdfY7HsTAFhviqVGBuZefbjYysryBbD3
nVr0grbBrSx1yCMKGFRlAa/HpbNPNE61mzHMxhPSPIlOdD7WXOSPHoLf+TfFKlyy
o8i7G2yMbTRhFKoSVBQplJsiXa0sX4MFtshofBuJcdT0rA2kRVcIdaPKrnB6gqYC
JB4J1J0c3cbZC/Dt0cvxMuWdkc0v7jGTAM/hGDuJguXUVP1s+Fyn9WSN0t8RVCiR
+oWzOU1lG/2ryR5Y0JqPrXC6hYtBvI50HXhj1uHpGnqeW8wpEO++0rxycKVPlJtX
/H62gVkojt+/5Weh355a6Sykc2qcpN77WqJsMeQl2+Qjn3waZFIrge317nigvYEC
GAujjnHogVS47cyGyfFV4gAyTP0QoCzBFxdTL8pczF1o2O5E//Nhfis3/qEpqIek
Y/G5kKCfCFrGs3HBPMsIexQTUc0VK0PsmwZrOv/iohUXNsPwnwqbG/Kqb1Whe+As
tV/R+XvZWUYAoQs6j/cHPnIKPfQN9mwzkMwVkGUSAFD8g0tuv7lLaWXwp5wDJuhM
qCNT2+3iw6MUKCXa6uuw+aJZwcRf8M2xJk9Qy93PQ3pE6gE9mJL9z7Hqzz43/9kU
NFQQf/UC4Ds28mY7ZKoEHlMgDgdlppT/mVv0+QeSvC3O2s3EcQ8zfTkCp3to8smQ
Y4ROGmKwIwJUO6N/qXQ5LaHFyLzG3U/HY43ETSHXVPAlOO4XribMYE7xt1+t0M1Y
2QzB3FKoW0yKIu3J0tEHTLdap4pRqoFKLzsFRZXwum9lTOx+pGi11rioofbLpA2s
Q8vBUD30X12Dbi79AUDhYrvnpCrHqz43w/Jn7sbTfNORKa7iXs0l+6rO/7Nbiuyp
rby2KBAGZeFiGlWr+asZCQKiwJyzv1cRPS83EQjO32oMhYkHKdfXTETOL8dhQvL2
RFkMkEidamJSRF2O6T7VQirTpYExIZ/xrsiwMGL1zgwVbiG7PlW7imDaZlk+XDbv
qbE8VMf/E4CxTi4yKr16QTFht2yrRz8Rh6GRNvAobbrrB2nGJdYwQJTDX1ZAK0uz
MS8/y++4Qtiz60S4TlFLLxjcQS+Nr3XkzXUAkoe7a7HN8dDUYIeGHIhKXI8C6Ltc
SxGu5U9tBXaGELRJ40fphKcJpWxu8YaZq27kH5hDeJgXiZ0vaRMGUXdnpZef4Wg8
Hu+WQPyCGH+MdoQYQrErZyUzUs9bD+8PsBYtXncoonb3M5SlqvWeYX96lJ6vlduz
LQ2zQn+z6dvZvpqPdNdJaIb/vwT0RAlP4fjQlAEULg0R73IBUwTFQQO6L3KzcJpm
aI63Zbz5vsr8xQFWX8KdTSbLOzXAroamVcywsCH+Q72fZJVd/v4GWoPsrxcRIZUY
tMxDZseRIHS00qKtx+SPG+ZdhiqGBfqEHQ4khabhP2bT2wqRy/m+OTcfkNexbGuT
6w6BDzsPuyyTDlKBHFyumyHn8tMxBUSVbPfTVx2UstmNCELY8abMvVaNiwnRI4lv
yDa4ecf2AKxi8NLdjpQO3d7VNMpjshbDnHc8tur3rxuszd94RNCOFMannnfwrM8d
Wt1IGqoFurIc7z5S7hsW9LjsDfS17MCVTDMfHQsyAf+7Gpf0ricYPKQ75gpTOYRd
oWqsopleetDCbjU9qYuC/9tyNyhcxLIE0k5ifJ1zt0j5p3vlBxayKSN1a3kEaK3c
KYBk4gRaj4DI48SX4zPAeJOrND76TXhr/prSZSH1Y5cXxuGuzPZ6o/26dEMoIFxu
pPaaK2vhVTLglDPZ/vl2cpfg1WOFwwGWtxDfXkHt5Z8Ze9xA6jsEPN6lRtqCLQoI
od9Jl4NHRvfg068D2AHGKaKEakqN1LUH8mu3gAEmAHvaKKMTLorAImpS8o8g5nVt
Tw7leddOy3YNIH5q70dNgraNxQ8zGJpQ40Uz+1CTiqbeW9L8rlreYdLyk6zH0ltF
ezQNlbLslwakmB8DkyTSIUJ4LBIVDe+olYZz+M0kUjLKRCHOhEAnkzbsb1bXtLRR
UbXq5NkC9R8lAW+PZjxUroQEFJGmzzpCyfHdJl1Ry880STUTAJXN4sri/UgRaab3
lc9daJbjbtHmt6bX64VZxXqSkvAFcMwN4eGSVXdREiiwvdnP614GJRuMpLUNwBEL
KWi+1xbj9enfCuWHY2Tw6c8NNYS+gU3sxcd+ckebUIrA5HjXPUg58HRBpGgtPkoj
C54RWu/pRsa2pshx2CCq6ZCx43xv5hyCWk7m+qvzjVEjaWJ2gEO3AIPHN4hG0Qeh
8c9pmLTIhr6YQEdhg2kcZaKKELZR53fW8mIgC6LvWcd1Xnjqr2Qc+TwmMCfVknLT
TebnoqdYBJP1MM+GpT4LXdc/KTTGgr3A671eTxORB8q7+S/6LiyW2QQwW3mkS3xI
1NcogUmE9ywZ8gEqNoaV5kPmVq70+OGVhM4eQvK4XBEPhtHNki4JJZGMqIt4BfFV
8F5/8f7o1vAXKj0avo7rf6C5+0cIMy8QxitIoslF2Xg6K84aopmHdTG9hPpPRPV+
YCSFRYR26nu8vfn1YV+E0rlU+8i+C3GxdXeYY5RNRXoY1WXKr6wMR9PYFBNLERHc
Vkw2JVEpIqswB+fihL/rb/BZZDshM7TgWr+yynO3MxyRlED/HdFV7XW/H8ITU6NQ
QP5FN8BQwQq7rmwKOYnXoVJdNdcqr+x4FgGfdBH4gvRKlmlFKd0UY/wavJlu1cBl
OzQtNEy0PGtQk4t9fylPcXlMx/gBo7DKHJ9sFdLEUtSYX79TnWeA4f0ejCrwMTt9
jF2LpFpD34Vhp5v0+caYn4K9oHby7JnoFjJrxBjTLhzdJQ16UlGEl08snahuyYUX
lkQIoJtVimT5s45c0LK6ODyxjBKMhEWm+ZmZOaVpYXXU2GaZ0XtGzpn+n0aq+6vq
12dvG6vzLRUsWFMjYz5zphOcWx/CPz3yAVmh6fBY/IEHkEvVihLUwydSaeXmwFZc
9hjX9FPC5kUb9IIN/9gmbYaxfupRUTInpVyAJ7paJ2LOjAKNlb60jDpoYOuSVNTt
w8MhzgF/hBqrDrfbAvJB1UL7jy2jYZGYFVaswi7bADhWKGbV1TLEn5lcDMjUfO57
10SbUT1smVPqNBL+6EX3jt9IU0xtiZrSGsR89/FJZ7ER8Q4oC1/OTl/yOWlbW0Ga
WMgflHQ5TRY80Qdp1WXPZmkdie6DFvfMS5uT5vDQwGIJCvwS9iz3jnSXrSJKkyhl
Qe8hIaHwuSbK3QTikM40s1pX+89Q8PSQ5pntcUJoNArSgAXWTIMwBEVqvze4cyaS
VMuNVA2Lvr5o52VCPf/G5KUBgYQijrEJofait7Si6pF9Zxco4rknJvaSjfLrEX2y
gCMwyGA+RsdhVvAqlSeJN1Gdjd1YRgiMcOjkedVlULMnQDwa2HHrsDoQ2/7AlGKK
TqKIv6ltsBJCGJnT0fion/ARzt67RfIMAG3jhJKJR4KnXCLTM+rpc/VSEKiI8AFA
wXBjXB20XWJbd5hedarXrELD7pWRT3XxPEvVFEJPqjBzOmJ+yppSCAHetvoLIenw
AT6tXzDkwBQvAV5r1sr3/aD7QdR9C2LPezEDkCtvD2TKrw+MGDKsc8RMCtXXphQP
yfwRG86NL/KFsGxwvniwnxzrkBZ6ofM3mi7P70QULg5NUp7rN/fwYEKd/cdA7gUr
6VgXKCTJluyOtsjTVGBefWaxWeAeKru3NWUtez769FfRIx31D5SbDOKqzFVxbF6N
4LcG8vjlZd9BS/TO4YrDiKAiP5FPUzIQZ2OioGr10PsijRXwE9GHB/2Ymzph1B1j
iADj19YqSxlfvTnoqVCin6JblPLx6iJ6bVktFJS3cqRDYrEIAsUI8DkPbGeufZL8
NxI+FCPel+afiUPfSwXftErUv84eLZC88nKVEz+HKrEq1+4kqDzQAU58Qhr769w4
5nLqAQyVxAo78xFYPyXx0y6E/Abb0zej3ic3zZ5f+iwW6wlUY+TDWRgf3k52NHk5
IEuExgAIhHjwkizVUqxBoxuFT5Nx3zTgwyBPuDePS1DPzMdZWOhKJPCbs+ezsDk4
LOAFfRyQLZsDjY3w8K3XXzCE4z6tLEsgqpTtVa/4++WnCIVhhUYlAIhFpJMMsKFO
KAHn2jqJvOJ0kZABK6rasQaimMVYxSoVaFMc/BBMpXc4TrQnZo5ly7zlAX/EkZV3
1OC29fXhU6sYNXLip1NauHQd6PiyuYrE7RTH/371O5ts5/9vyyUn5OFQ7M4acKPa
6J6c3e4DFbgS/hWozETr8in60NysPPleObOZ3uMlPC4JIzeG4XSwl/Ok51rIiuUV
zp6ddykqOogt1uI2Zagp1Oz+l7B4ZMMQ1RfwZOppPpJi8VeNPr3sFPmk5xdmYU62
tp67WxDmMkjkCG+tDmH8TWMQEqiUi+HiCn615Hc9wqy45pdowVsuXtYGNLigM5RO
yZks28BCnm17Q2r0byg11GaNltPz+rELKbx1WP5hA635nuAI8FJFhsAOmGgM7VTY
KQIEBmQ1W6PFlqcgbIxvo4rJzxPfHpsDchILGhcqHBlZgLCe/ddAU7xocZx+sDJf
wTx1JBHg30tW5T1ygmjwnMG0QMc+LF8A2IGJmT5rSia2cQiP5BZC/46DY7ae+2qu
iUAGbNDKlvdz3Cwf0CvAgZzWiynORQkKmLTv1Ntc87WsW91N/0P1MnO58noKLTtF
MTwbuiCKdkKP9iv3DapHUo3iOjRQA0ydugGTrY9jb9J0xx1PBM4XsjXhC5aqgBVf
3F75RdrPBO56xjvA9lflxZn7jUUbgd4gJc/TSez1J3W7vkoUAl3I0NtyYnVOehIu
7WsPnXz6r+mnwjUJ3vCmtsm3mdWCQJp2XK6bBmNsHbib+6VinsW1JxWxBHLhBkip
SmSJEH2+zOFyvKkv0PEyI1Qs9tFpeANDjsOastofkH5E8KIMbQGZe/mGegubpbhW
0NeAZbYfday40QxGrrDl/naijugvuMrO1iKF2P1HKlYHr7juC+BaUWDGicG6HYSD
+2cVtLArf0cxmub5Fus45lZtqsxZQnWT4RRX4iOcN1Cep6YU8K82slP8q7FJupe3
h3r1ehPFIN7ryzj8B+/fXDgcoYr2rmudmmR1bL7dZUcUz5hsR7+5PQo6sFWvIH9J
gTj939WW5wde18lhvKuV+Sqbe/mJhYfC6MFUmwX2AW8jjN66t/zTN8WGXK/fkHv8
CUmPooZHy3QvJY1f6euWz6QhzfNR7BCatSwWr+PimKhBjhpn33l8wjroWNop4GXK
P4SKxQCqX4wVZ5WjuRwp2O0tkgCJVduN1tu6gmYEd1K7OX+iC8ucOyROO3l2zY1x
0MtIEwP2iZ10YSMpCkn3ZwdiaqN2x5oTZIO6GLskeupqC/fKgGRziWhZk/jdV/j7
gctJ3/yb/tClltE1Zqd0tAs9POGdz9j6+JLyjnv64Zd9SFQhBaOfLtjo4zlv7UwR
FL12zBEc27suN7/lOyePyaXVz6+4eM0QnHKwHyos+zlZyLuHmQSMHQ+eo1ECjOVW
/XNNTNTh6Jz8iJlVRPKYzNcaywaVb0UGVy2KhPK+RcRv477ZGhph9pknU2VZfdK3
tH5GUIxGiXI/xTZL20EDykxHYRGmafPrzxbQLPWTwuHzs8LFU3HPswwouMe1EhJ8
YAhhWrlaf5rsNYaGm1NCjFv6V0xIKBsfoOkHPEA0XVemNhEGPP3bAFyF5+36pDVk
aXGG0q2L3TWoHkwdJxD7ZM2UwXZDt/jLXtAOU2jzI9mbBG6ZltqssowB2vPb2ROD
Oz+OupeJgKDV3oYNHianI34DMJC4lx1cykFCVOea+WhKL31UKbtsI+k41+y6wdXU
t8JfqLxoXDIz3Klaj39BQKsQDyxfn6jFeGCMtO8bFIlRyHSLqW3m6Z3pJbe3fmrb
kuahYP+hCism5A4muj7ANAk5TC8W2hc0YnqzgWix6SmTMRm+DOnK28/qkiknuqLT
QigYzkxZ7oDe8/c2W+c3T0DCZXpQB0VBvRv9lMBS7sdxLVo1rA8uBuhviML53V18
T9ypoU/QgMYXfBoTuDpSUGm3mu9hdUSnyTOy9fEAKSJPuxS+09z5BeIxwaO8go6z
1XpS6ZMP9dcVJ2/b1z2KTe8GzBzgOaEtJsXSTDb93H1/BQoeoFrcDxXDZLIF3zkC
XOUMgNentCqb8PncBEFNNXzewFemkwVOzFzgFGlW8D+NzSSU5niwkuyhCdlaRmWl
lxa0Ep3zkMBBZtcLboKEnk2uP+aFO0aZPiW9N61UFSrZPO0W/CKyCWtbha33UWro
9FxhNxUtBy4qvkbLl/1YJJKOcRyQ1ks3mR3HzopKj2KLRxa1wy9v96beJyC+6pQk
MdHcva7D6POC+EXVgL1cg/JlikHyGqSWnHojEtHV++eHkOoTurk14NXBIMLbV/H7
1l++dOMWZ9eAAocTGUVe191AMvWoGtVm5Nbv6SYEDr3/Phes+NZbYRmwdDJLN1gH
VAILtMfyydn33fw7Dn/GcbvefIiP+WeiiydnHFQ50ljJI79EIQyzP9i7xFIlzo3j
h1tloNOhOzczawsz3ZjstW6l1C0E0AZn9C5i2EHsVWjJMGGVwIp4y1GyZ4tcFvsn
z9ty/ndeYf7jVjl6ojDnOfRNA+Q3e3fAuMb2crzxfIM07mLRaKElGhbvvP7xd5u4
hR88o9XB1/avVZpyjWytMdHwT2vHhGcaXuntmW/i0aVbVzfcRMLbm8xePyeTuzGa
QhEwVwjDFCpyZ3izYSqwebdwHhIzU5C2k6Hh+U6uRww/UyWDR2XrZwuE9GUgqvzS
hE7O+Y6irCkEceEPoRjKJX2hXhNQZcAmRojw4c2jpWCErE/WvICINVmTqHeSslBo
U4pGqu1wqs21RHNF6c4/bCRSEgjw0KFEeo6p3zmCaLncsLBpqObv22PMiWKZ3xvk
rDjo6GnsEthPkpnr4z/YaE/yl8uwKYyJO4Umx7R3r/KizFuoAI7A3AWvETdmzzYO
eofJaWiqvq8sXWO6sBnzClc66+l3kXvBGJMAtoNiB2porey5Eg97cznqCfOjRbIO
UNYEIKi9JTPoTBpBMFK2PIBSHDdJseRdDHuyDdmbCV1XtBAm0cywdizkD1WeJRYQ
h0YLu4e9G7sc5WbsTnwgFRej+BHYKQ6JMIUbUtARzW128ypoJhU8EXZcbZCCZSkK
kj7WKZ1MNf6WjcHAQ5CZ4wOBOVgDuFg+7MpOwNYCPwlx6sPI899/9awpGQzn8Usu
3E3pCx2O2ZaLDc6yyDIXVn+ysv3452ii8AMrvklAODTpuumk2p1f2Ko9JqY/UsmC
ioYkTHrleJ62SUXhWeHb3ioE7TlFx05XbBA4Od70mJoEwbyt/nAEmCbvH0l3Yx+z
ieko+HoRBeBgBMI+y5d1U4f5omJ/5twpmfjN5mHqojsDToOKE4cN6iM5Ng71JVIR
7pq0UbPnoiN1rGhYbfJ4UMncr5RSd01TiweaOoGqwHVhHEKFGaty5Zq8E4hxyGtl
xG3niGoP+PPebiwA1xQsgzhT1BBEcBgqQ2CyOH2k4ATfl4RHdPKQkSm9Iiq6s+QL
OC94AhTrOFWJ4iqLXXLwx5sPyY9+PKt4QCPndV2eTS3COyBWcHKbE+uSahQgB8b/
eVNzyWmR74s6pt7bSkIhQ5N+D9ZXHTruZSy+nXTdQUPy136GKWy7J5VAHRQ9PdEn
RgTePoG7WOXiuPoRGXIpAB6yX+ehjBydmonweW/726sdq2NH79RxyAPQFEc2V07j
Rw+zUYf9vhlf0RmxjRQ3/tviynDMAHOhrl6f+TGmrLzSnlIJO72nSjJAx52r/z65
vNB3ECb5GtfIEXmpkMnSwShOQDUaTXnxdVPhd3B0FecOZYqhtqxqr7yy12iI7853
eTg4jI5Sm35+LUws29b371qRrshDjJZh4y5jbAlw93RIN2Ct3rHj3XXHNfChaChj
4dNFBuA1XbZIW5fEDRzcM/zg0FfJ3gpMVNm8hxPwcNYD90tltsEj4bwWjqq4ZjtB
DRDokyvsHdPW/mKOlkrwFhe5wQAa71H/mTsLXW9n21hZbM0mlgqkuNmFYaVR6QQ2
CU7XhRXAs03ssxx4zge14p7vn3nqSAro06NLHtX14JG2/87kUOKcEFfvWRR0Jn3s
U4MsWSTDZfhLxuWTjLxgV9pfsYZ6izYIPMLtKd6y9Xmmj+GZpK7lzvLnZ9Y+M9y+
yi96mmkrL1jsFSM9w5arELvXZWXtu5/+f75+AfdSdpkUBdMMF4hshGNtvyWbyu84
fPnuIrYAH6yxLBEs+P1aZ5UZB4XslNcypcgE9vngkkQo7Sg5pv+bnXdjfkZ9zIis
PV3LOmjnsEzUV2cxn1g/drXWkfJ9HZTvjOZT9BbkyRX32LF5LQ/DDqG5ufjYRW9q
FccLnu/Y+L4x46YXCi7jcNvtEpjQauKc7raMSyNaF49G0cuvxeLEtNCbaWqg2cOj
RDWVryc+J+FahnX/aZHz6h9RdDLovRr8KTXjD1sw06c3mCd5Nyy65tYHyvo0S87F
QE2teTTmnaaWI/nQ5YDd8wUKx8JYPWNdYwClBrz4ETyS30jCYYz0M0ltQVwOm04N
ANW5X5owBFOsdg22ev7O+5EBrVX18jonm6DS8QveePTQFW+DxZhqs1mqxRS1lQqT
/ho4qgzF+c7M7/nE7tNEKnPvEGp2gFhYNkKCiNi+GJr34QZ7nwH6gcgOiABSfU9Q
kdPLPyXr887ZeGv/sBcUSOYPMPmNMUdAUq0aF9e2qcpuOcrRzHxpM2KePkETOnO/
bw0Qla7fy37G0Bb4C2wCN7Gdwxl05uyukFilpvwJo324pbFajyq0n2pErkewM0oc
xYPeTn0JH36KPT0ucXaJys9B3dU4YvbvFvJiLDejBEEopynQOvlTfo45K/ZJuB70
0NQv8lk1ezCRZ/px8X8rf0PJk0xXIV95ITeA6+1xPxDo1xCoNuoH6dkZT5egaPZu
KTz8nFhtZ8Kg4eyg5ivcneDeP6N6gMSxUwaJtHduw+3hlOGXhrLZM9t4BqOe3aba
4en+Y2RbWuTLPP52SL0qslS/Yo1ziLcC6pNfLywgsqJ6hld2RsPiAH+WRzxnGrnG
1yVf8t6CdOBlPaZhYC23mWDHlfbAM13vmN/vIeVE/iLvEOWYrg/oh1OWbmO7iQLo
g/mTSStqd3Do8XeDjvLeOlPGgIzpkk41uhSj+xZ/gMWl9MGZ+tjcWgGT55c+sXrr
pa3uhkUW3GIkM0+2Jik1BjbjmBM+JojmKl/wj8/Uen5ccp6GMzA3WIH1gPRETyEk
2UFR9HxukXoiWzG/yCOfXYDEQaXJ2UiTfoIoEtgCI1+wVxAlZL+iUTwnGA8+4idJ
qGf24r8Hh0ifItxzdZS5xqclzl5pIvMKrDZx/HXRFE0Q38eH3Gz6QUf2n4lPehLh
zEWZSzi0mQwiD9mR1ap1N3Y0NLmA3Gj2+hrJDWxuzEtvd/TPYEcoqZlqhClNK9Te
BH2JOTYQdVfX50REZN6aaiXhpGy9J0SI8NoudJ5ftTOV5GUfTL7g8kJrEr2GgKPf
cbiUYE7xC8D9K88dC+RfcmKlL29u6Fy1NscugAOW9bMu+ZcauUhJb5Um8+6SZnnz
ptDD9xSIlwX8T9niOUm/qIpwFCtrZjL+B8q7H/2zispsqGgXNghX2j0O384TarMt
uypY62aTMo8ygMNe5GznSf9dLHs7SiysKtzbgbtLXGn1fWPpTyz8BrHnkqLCN7r8
bOXlgyUBXNO1A4zp0qk9Vpon0m2jrzNC7wuSd0J5qgvr2rbxBuLn+WOACKCwn4qm
moJedbtmjl29hid/m2M3CPTmmkFbVAcPubUVh9skPB9YsElSzkNlpjUCkoyKV5YW
UTtlTKU3kH4wPdfeyBgbo7nTMy3B0aphQZwKfJ5MdXGDAM61MrmBa4BEaSHYTbUi
dxcuWbTfPBSjTNZDHSb1Xzqqn/2O8bOJx1t66WlXPyfCdFbBsGl2nHFDEngMuGAu
EHVf4xoJHyrJ8iDkIsHsykkrgVkCOLMq4YhqMy0hynH1Lcs88gz9Msa7Q7mdu4d9
F/UJGDo/2ulWhMB0geZD2hvNGwVhr/WS6Qb9kGn/TfyWxBVMklkECXAQEWj+kqkh
3SdN2WjpKKEv7piYK3+KTgIm1cbMUiF4n7X2T3sZxRnMKSj5ogsMYey3Hx5er/YZ
hkBfVBjx8OajdQ/cmiSCspj4ImnjbOokKAiRtswNWXebn+USI1YxkWG6Q888MGLI
1T1sLtROqNWud9CXIz587eyRhWHMPIcR/dOXt3/x/9Eby+LJ0t4iEQctJyzmSQmh
4Cw7OXxIxBfVHgkOhyg2DG9eXdUj4oJm0D+t8QAk+hrKQSGy8SUcyYsnc9gRFF0d
n6wwKBi+yXZl5YftJMw+LDIir0xgN3DMFFAHdYnJy3wwNzN8viIGFE/3Dfzn60zu
DooY0nJUs4ywnklTTetvhiHL8OqAG7Kw0Ox/AtjwRgmN+h+DHVjFJdxFDiAZt8dp
zrC9pp9a4u+qupt+KCKJBzDooPKlpiRYfOqosCXE6/Gp+FAq6z9GYZUPM6WKdwvk
vhOmJ9Y1IijEIqrAxdCO+mb9RYQCQ57hscLLlLdxtk8MGpMlf3FV9W+dwdiDdvA4
O5C6Ofiq6huAoklbnVdx1AE/FHfAoJxGg8fEWuSyAgDZyN8fCTg7kJAvfBYVKcG0
ei2ATTGufFx5NdequBWCFn60O+JvkTUiN3ayLri+QTQ8b9okSrn7P0Q+16WN0xRf
eJTahTVr2ILr3BqXx4QDxcK2rt2CCL9FaTinq1pb2u5tzd6a/Am/rNw5nRJUhdmA
pDApJS/CU4adzME+vOhkPh0qxdv+0fKdJr1VcYaKYAd5vr3g691j6P86IgrBFhlb
ZuW6wwzb0Tn/u73IwA/SQu+Av8+AeHvkQThq1d/VTlLa4fGisNJ7z9iw+n9ZH+Sm
ijz4ioduou/YPaeaf3ZAZaqZxNWVcTxZj2C+zf0lj2p18dYw6smBPB0Q4SgKCHvH
Hogj3RpydKXx4il5c+hRU2RykWrQchOSCuarNep255H4TVmfIDeZxal0h3lqERJn
l3lEqavExno9O7BBewNF67B6hL5+SVrpGE1ze8cBOLfVmCz/piydn0mNo6f+h7/4
E+e4Mxve3N2iu+UXfSkA2NlBQvb8yKIiQMoPkKal52QEOIafEOXBYGmUKxFmTuAu
KSt2QXz+NamHBsjMO+tdJ7V44rv6yjQUh2koMOrYBdTrUXSOdEInA4YHmpAxNN26
qcNP2kO5RQ7Mu5McKZimhC9L0EGBwYAMQXjVaXGzsw0uNxJRZ+8ORPKpmVVzq8Pw
NkYLViYnWtD3qc5YYzC4BY+wP8uIBMbJZ4DX+yZ0VzAIckO1/NMkrNT/MEgw6wav
y9z2/zmi7OlwsYlUVUKSqqBe0eo08fZUWVhxEA5E8IDV5Yxy0RmxiWn5AwRLhgAL
tOhT1kj9tZWSImF2Rq7Bg+bhLYG34RQaYlWXBdh/F2FqiHtqepKSTQuxNrxHWE70
syIJF8SpgMacLCHo6NG8gMCO4jbFwDtjjzNXW4odJFwcWZhYMJens8dl5TfXxx50
js1Gj3h8CO8xNHMn8oZ/WgXMiQ//GsD7ZZQfKlFEcBUsq5ZE0/8/JwsIr+8DlfXG
/X4ZWyAv8jYHFKxLH69f2KgDXfb/Jflzv1hoQR2/nWoWw2V9JCmMZ8T8aOqe5pPe
/eW+F06dHDM2vWLir8UbjkvrSp0uB82tW6dUTyUTqT8uHazXbO4yJtpXokdztwU9
RMzgftHejGl8JTegjHmKaVlAz3dqz3+SgrLIe21icsB5/jY8tccVg8NMGPqeSz3V
HOQ5MpiujF2ov1BtDFS0rBv7C2v/ntVThjiV1wMa5avCxQwbVkWUhzy6fx6G3jn7
XrLAOXJHGRzyt0lQqdy44BFog35Z9Ci2B8C5zYyyJeer3wcyJw4Ybv3jRYSlstSS
p91ljkDAJv02YMKX/sLgLm/8U7wXabOHOnJWzNnwO7M10QZ7CIK7U59vCAIq2bMn
pKdBiJ1y+R+E/CUjDRL09F5bd/1oQkxmp0Ye+a4b0z5FahXXvmukSqEy8r0kw53m
ASw/AczljlPl0drMSWk2clqeWA87JD1L1+3SjG6HWpdY8DgueMwZm2uhE3HzSgQx
mU4Tei66I7VIKev6BeNJcmRHKztYaGmXNGDanFP0dHZ1V5OFXbv8/Svjq1m8yXRZ
HP4IpHgFIu42e343cLNGgYMoOBnga741ssJ/Ntzfr34fwAbWSgvuoPWlVLxqUAXJ
Tae+TZ07rd4iIFdxc5iKYYYMboMpuEb/GWqFT2ygqLa4DQcyj/VhJ7gakP+Nz+wJ
CFZpoQzjhUFY0NRMmx+pa8wrR8y8yS47pRqnrJafOPL56c4xXrhA7yYFo++bqKRB
wHL/X+nGChBOKAOJmLfeV4MTcAR2P43yUcc+GaYlFzuISCudu+i5u1XVE4xhAO/f
vXXZT4b4XEMmKxEHglVXESmpystVeVD4pCuVN9yeusu+HVO+uyy53WqdCSQGB9Ev
/GVqndm0BlYAdxFpSCtXfZXC+wihaJaxlHuoIC1Q8A+BQ85eghVtz5Sv9l6Za/f9
1yn8sDbfqNSvRqHDhjjtsWGYGSv2YVzQeYgWwYS15uBkAyiRQG4uyPFBoUNs+Y6p
eupyE0TFBm6WAMxio8PyKdv3oGmvWb5ahIsaIemQ/6R6O/1WhGZCRyGa3IrI7F2n
nwgEIvaGc0PyKliY8j+a3C28NizLAULkpqmpuggaPQ38Gm5+USAtgy/3FQIQ/wxN
a+8tCUDD5PAQEOE4xkNxkNAK96ANBm+yhlr3cdvwtnI7gP5SWdf2RyEd9z2yzFKk
apbo3oKPOOnV5hR8wY4Vf/otH/JVCnOg26cS0ZQ+R+PQORdDcNWXJBdzwYJPUmK2
MTD0K0etWM/o/tzfEsf82W8C6wBrjM4Zmwp205OoJeLnzT9XsxrDmb4blNn+mnlg
uMQ3P+YX8raKtHiZ5ZcLVu9PBPDfZ9pdL+DvuP70Om9kVmaRLlrTI9mctlC+L3BM
AvmezGA/xQK1pFKQE3+AD6FDs2y6xWHa8zBUyy/zQ0MhQsr2vzZ8+yVegIsRKEGl
1yStzQn72Td+OYRrxNTVQ4QdPOSTVimmWbq4Src9SRdfvNblDtQ8ooB9VRsvy06h
iWEQWPHNONR3/gWMwS9pOdOQ7F4lknXIxmFa+9WHeKqmTsfxliz1Af5F/0odSm9+
HY+mvdNdygrh8DqtEMJJEexg2oqh/1MIj2x2z5T7kQb1bOaU7Qb6etBIxAHg3V6y
NTDfe4/d3uUf5rhfS7TTtnpjSftr6YGEA2bp2GZPiEtr7L+PCSb4JjfFgY9YH/2S
5LiVJfbt3PVk40HB8bPGERe0xSQ3MFZmXlm/hCQjMA4MXUDSIg6HdXF9NA5832+B
M+f2BLznqPs8DdvBMWNN2QzlWLRkGV+UOaewt2ANSptERAu7yI/rNO8SDSFQZY68
D55udcslMXudKL/frxHNlUMuLyYVnPUFztNhrNDYY6CWE3rH9u2Dtc7OiBNZUJBi
ggiUVV+Pb7CGh0ZY81bhNTNdJ/xrVcBbB7y+Nhep8/KCv2vSfCSgoWYX7WGEswqz
Kfp6nfDjis/nqvMVwzUJYAmmXEpiq+lrQDvR/4IOmxFwEWeC4k2UVVqGYQLuNQPA
/2NhgUZ7aF6K7rFy/eOZfMbiEq+Mcvd/14yfD3RvJ8SsUIML8QP0H+BCEzwaqIQU
2RmMlMmS2wEi+ZBe81O1X/iRUjqbqIT+q2MrDKKRxOj3j+r3znVWjCb+wu37rogg
1Ugr99QiR2t1/UF5h+/VjP36ztCKNyfNZF90tSh4GHnxpoTEY3nwU7pS+uEJYRvI
yg9HfQWHO1qgyWbjF8bu9ebf5vv7Yik+RtFcFH3Vyy+QvoDRri+TNoaQ8wDodT+V
/vnJJbw+dNd7nKx9o5GRV6guLlCZUaqjUEy6GUGXTUIj3ujE871QvSNRVktQIy0a
ZXYCz9J0zbEA+7I3riOquxgA4vvibAh5wXpd5VrrZb/FYaS4Rg1g5ZYp3sqDOg2m
LwCZXpaNcuwKOrWUcjEDUEsJJXPE4/BtaDCzki86hAo6GiqzxyJqxVvXZLjyAzNF
nSLIRRU+UvogkGp/NMRgQEOdUT+wIFltFGOzlhLf81tZ8OKQD84BPUl09O0gc1hV
4yaGyitUe/5eYmfPNetHLEa3O3VbMNQpGpsTwNjkgI4rmHGXmBFC/VLa84xqd8ow
IsNfXYEHN+xwx4/hhzk/mYrydOoghzB0pTLP+UJ/qjaD4RE8t549G7IREientugN
xyedy3XUgoH5fvDQ3ysVSZ2CZp6kKvkVKRRAOCfn2LHfBtlXhpMaaVDiFBQBTTON
x8MwYCgls336GGV9a6urjfeZ5bQSI6tlFJ644CWpIg9nMkQpDfUtHMHRGgaNiYrc
YiVd8fBn1+NuQ4l/HkyzPaT+1v9ToockY/0bHG5fXtspdTxGgVDKtjwwKoa1l/O/
x1nXJ9NChEOUqpMVguMz2Yc4BCiDv8xg1dmlbsaRY6fD5HW5Q0uf0jsZt3yzQwpS
/nf5dqqaBfVTFPS5yHay/FhFbh/VRvqZlvrrDTui/6C8ZZa70c1dkgghfoVGhgR3
WeGLl6jcj73Rxktih+Zi8Zwh0TtlFQuPNXPkhy5OAYE5CgU8s9k/2clrjtfEAv2G
ftPqM0Og3LE7To4PbQTR7W3lDQ0iVYzrSqNjuRWiob79YMwmMd13DQ1G2dGvX3ri
gnToYWsM2dDTCabbgRbscKYPB3sSk4mJw64CZRSdInX1JAh7PPAc3TxxcjHC55+m
GbK7d4ezqND960Z8LoxsGiZfjZ7i6bg/JDXJC4ZBahWeEmtbvVnLozuCUdho3j7z
UC4scNyDn6+Eq8KHyxxpQvw/4qJfaraZ7scNMoSrNV7doWXmVlC7dA5osO8MXQVl
tFqIdcZ3yOwGLg6PLxCruAjD8M3SLpfd3R6PMBfpyxbkMP4XrakRSUc/1rRA1ens
QulceWtVtRQAynmEcEYbQuQ3rDzRp4ZuyUBajqK4vVkNCjgHDzgbsXzGCrSf4My+
eHVWqMWBMGic704+lpKZri3GbM5Dc/8gB696xfwLaBIG4H0cVi5Z9FApXmpx2CJm
6BXUQjGni/h2n+U5Md2NwOM5CurSCc0+DFN6h8dY0SP0fw4EzyiaAsu/jTDhcb+w
Q9mRvWjV3eTZqPfUE+BOFHuRv+72D2cLCfPfaolwH3P4XvenI+oFMMtPUCcwsi4p
YkD9uis+hesFS+bN2emO0KAB75q4huw+Hju3Te3j8FWdUtW8Bh0W9YJTP/+TAgy0
ooWQqGWdxCtNyfbTsdNML+SaeTpdgEg34b6oQ3Y/6Sp/Taq2lOO4xxDXCJ8NOIom
caBXNPrjhYjiNdyYTCx2Xuu1E5t/U+4xBBgfOiI+p4xZilGUjlKm+BFy+Zyu93zT
eUuxxrbby7H4Jv/+WCsVBMW19CDkZprthkaq+uKnETc1gyPYHgWBFiJ2DFIc4UXM
JE/CO/y5VOxo0P1CuVzw5VmWVK6A432xJ026hL5vurvfFoC3RpScIZIBghxaSgNH
EWRMwUUBh4zfdZkPSj6Ng0oPsC2o50I8iORKpyWmPyorBLL6HaEjhILsAA2oogPj
hqAI+vefOcjNB7QrQqI3aVU6vhUqSPV38ER8/jwQsMmZT087GYilWmIIJfH7e+TL
sJgRVPRUZGNYYSG8YppiDoFpiDdvvmY1mALWG6CFnxaaRzNRLW3ykPPCZYr9uUq1
f4p40lMnKeP7ulNDQnmEXfMvDAM84asa6A2yHFRTmzcjHTtVH6G7bybOzl04rXPk
gnbxzH+xmatYShcDc70fPupnl5zIhyK1yx75Ib8HCJ1D7rVfQQa327b/Q03EXvTn
SB5I1basRe4HYFPAFwoNBYAqSon1bL+eZkgYWbLDsPwO+v2I7HgZ8fjSZxPpP4N3
ZvRuHJdqESTwSy9DYXIia8zfLfuwUWPQUM6Aim4Yu30PoB2qQcHdC4kO3FTmpISY
S3C8d+AhRIN4vwTrLX4RzSCTE1HxRCyrkVvamxju/2EzP9RWh0hHdx1G7l5X/a3H
AK4qiQjRIu90Uv1ALhg+wqrw4gSboHMHZ48LkyxQfVZPTEbZKkd8F1yMk23iZU95
UPMwBfBXB4Ls0D18O7dgo+VbVeqhkZ8mgsXpkIbvBxcu3GuqN8XzirX7pCA0qyCz
7BT/EOnk4wYeTgdyHRO1SeHhPftvIyh67m1pMFI6ReRCH4yH5onxXJTxqGkhjDb8
KmMTBBkmT93pCkVhPoykkjMF9vs70Llwjm7anIvnfaXGv8QD+vo03/01ijxNwIo4
EFxigPsz4J+La81T/EkQzoBqQZORxQmWFIdVxAkS1wmNWwfVNY3EJeAfcJltyuq3
XjxK4mvq1tgjcfP15bEhlqrACjSu2QRsJzF4d++tA6O+b4kGIGFZovoJlWVegq1D
ALSdIm81u/wETLUA9If7KbT1rR7ZgnIQatZLHEYaFSPNIOnFsjaWyKfLH3rg0252
xx8FU+6M1A/yy2bjt0GDd41HEEJQRCPoT1z/E4BvZRdXTti3pYUMo7+bffpFfq0J
EEJwA1fIwDFPGD+bEf0glH5GGLyvfXTPxUq83IC/PW2/1KYvOdcD7OLSoZhBHOs5
5XkCKtD3+/eK0LY3RHnxyHUSXkpuv6TgJEyBOPK0rAQnxlZnYFujkR3bN4R+KAK4
QhYhFYDYbX/dQXYnYkvLhJ25IL9qejnfzQwPWJyHWRbXwCv6bMjruUCfsiAwH+eZ
RXMuyMZEa2/rHQ9ZWwtZQHL2agCNE89Sh5HZn78rGEvSaPyaW8eqCpJmuZY+dfzz
UPRSG1bCUT7Lyuc5dn5MP+qhNaCnxGMICJXrzsOEtlaUs0XzF+rD+5KfAFZ7MLFS
UI+C3vkt4ZitH3VbO+IFzas1oEZ3GpHB0ncA9vnf47JJbAzoUxGgdDdHUkgLJ9de
LhP17wZ+rK0fGhNv1zsygHI6Fb9kySr1BAabRutmRI/rDI8fA/vJMsPN99PBB1G9
tFuuMxnXG1n/tOaP+jevzYIv51cVMKm0k+EPzGy1AiZG0SqRk/opMQJIU0fhhMr2
V5z4tJjoMFcMWhJI/3VGyxLJmYsub/4ChPAhbZF/awn5cKMlDOeSv3GBkuvt/HVA
+lKM3so1wJsj/X9aAQ9bY8dNzhzTO+TX+3vY+YvcQbomZdrKU+h20QdxNfx5Nt9z
nSevwiyHD0YeyH2I6/4YM6w2eeUyvOvvsGpLF9192eEUZyTncLo34831TqhdiQM2
qoBzJEpcNh7eDn1Vwz07gO1/GnkJQVXcOHSdDb39DxYzfaV1KhjzsWhvS8tkhl0b
bqelfxmt8PCaCzoKiNUtrhNrN4+Ybfru2XmDGC35uEUH0WWBAQOsT2KXB2hHO0lI
mwO5ukZYEmLchGAYDeJGwSQnB5E5KVvs/zfBQNmQykiKhKVYcQErvTbqx/mKfGeM
qvU7GLdHYQJIqagoiGN+W8TPLjmx4nRgbEtWm/ORxPRj+ujeA9z3dRhXXP9eJXEb
fVyR8oIgsOIcoyi5jZxtesFTDpd5A5Dh41sSN6B4HTF9uxiY+XjLRRHZjGMZUI52
BmoXsJtbZkVfOltwKkRb/oM83IBdoE5BmUw1Mn3P9BfvAHZTAHrgLJIdOmLDVeMu
22tfjcIueBt+i9KREs1c2LDK78WJGPdxPzhN/SsGkJKancYUNLjiBrel+9TfJSqp
kpzrbW4XA57h0xMvwdoDsCrjl84x32ITxYwY0FCrVqIQzlLCLHiomWu8oQEXbCGH
Zz+ZWqrUaU+qG+ISoUjX5Q+91qM715ecdzn9r5KcDbhjaEYZwjBvf3hhyEkb6DNR
5FVzr2WEcqg0KewmvVjsx5SIUn48MPirBVeCyd7JX+b5WKxkqeVtJ+4Dje2inSga
MZXRCXmiS3C4BRVLnAtijp491AhhuERyLUhAatmhUMfgIxJ3dc4KDIWV38H5pVBK
gy/YbxDsabLdfATZx2QGlTohwVTFd1Y7tdLsyCu013rUsHtJ2yjDh2ZdyVzTl8TD
BVQC5V8VjUGoSxmZ2Re22cktsfxf7bMBAXEjDOxL58bpd8ATF5XqyJfRLNRboiRb
Dy7tv4R7l+740mH+jVC/u82RAjVl0qFZ6MKuNtspORcwj5fGIRw2cd7EGv3xcW51
QCa1uCU4GxPNdw6mvBYo1YNNUVBeINLfC28dIDiassY+pVgb2/6tGYXILmpPRn3r
WkWZK+eJUARkqtE0tR/iyjeYU464D9ypfnHOz73WQo33Ve0mr7odBRKv6xEOFe7x
5Hhr7GdFhfp/3MpF60YnES/Asp+LlfansKhPpFX8ezamV8P6AQYbzemWYiJ5jFsZ
lZK+7YFasR4qziAbfosTkyr4VIFaLkPxQ8r5SRBVHkjJvgKlmZOGLKa8rbxCnvzQ
gLh535UtcG42J82tz5VwyY03Tl9WgKvji96Jirxq0kbXmN3kcbF4dqPL2t5UuqCJ
ehZJBzskd5ub7mW9ObQHjts9i2wmxWxedXYiz/Y7vOe6L9oFtDwO6FLhHrIJOdU7
v/ybIVpaPfbrbwQsHRW/uOGGBHICeADxicdg2rCZlQcsKAKwPlSsJxVz917rL8zl
krWIAUZELvoQPrm8hL6XiHjF/JhzGfTlLutL9EPmrvgFTI/HsWIk7x1nhyLzqCA6
d4mkwqlII5J0rvz5j0LsFowlky8SKJe+PzGHHsMcy29zgmBvW4ls9iIVZA2V3PNV
X9Wi3Zpb678sFuYt98qrbroeJs/SK1z9mIe/Pp0MnhvgsR+JNBSY1fFrRaEtukV4
KuS5dhdkwISwG+8NDUq11fBadB1XyqlGz6/tYXzAI6/NlvPQAt1YuMM9huBuXOmQ
KSR5PUfigirkigc6TDUm7ce4MlFpfyxV4WmauhL9vnVs09icpVclVvSPYapTaDde
g97MpyTTqDf0uXTIiCSuuIzA4TbZ7i2KXKdu3kLBLmg+ck0OuqE2FoEO9et0IPBx
N2DkdiazUkenMIM+bNzue9Y3S3pXC2Fhjdbx1EVnXJzpMnZW7FNgsxHci4tNdLF3
vEGKMRvFQ6Y4cOocBogTA0fYT+2uxswq9nqhu9rVxDjRfuM8/4EkO3b96bAy/w78
S+bb3K1cSwizAcLBDx3D1lmiMT97+WT26Wrv8HAHPightLDP3EL356GYxBIT2yB4
mQpJJlYLR5q5PIxLX63BjQlOlDi9o1aJGq4nkQONTodasBE9mDEYh2dttUjTH/Qv
mfpmQa2vjAPzNv46k1ChBNUfledUGRLy+BLTC8R4LdJ2tQIzYyAPtECYYp6vodCE
orP+YsqZ41RbtzjdvKRpMRLDX3Tx5nsaz+SkKsHo3+2i/wvTjRVzck+VSohvBCVY
tuBdt2B4iLAzJiZSKTtDfvz9SzeSa5v9G6R5h74RJYHkPHcKmwshQ+xBdaaFZwZ0
QezEjr5dVrUavTU728xlPQVqC2uhZ9wAvF2fj2ecP27B/RurXRsbEqio73VIdJMm
X+B+Dvt6Ci3Wsce2ZvKJqnaXPSehC2aCWJTqm0gHu6oGyduLGCydq0WV4iRNNXmF
x8hnqrs2w74Tsc34tEHXQOnl+gaXu0b6ozA8lT2Mjo2ov1WBju6Qm/K0WEP/YWBv
Zl41oWIsUmpGVsZjyzsuA97Z7mxipVa9sUMfpeFXlUBPbyvnxz3qVUDyG6Z+SJsU
QtlzGZ/1cYZ8CUMQoW50IXnxlXLUUjm2AncLlW2MGfJCIRssO+2+n9f5Gxz4EGs8
AfApebO4JifXDc4gjwHZLwe9Gf8kwOiypcR3AWJa8RCkJKmR5Ufe2O7Me9LSRH03
6jPoEaN43+X4uBLLh1QL7odgkSdM1sVoGC8iV1AyHwWR7C4zOhl1p+rtcqhNBklX
8ATm0nbAhkPwNTSQKNmuo/xTMzQJ2l1pyZndmFdWWaO1uMgeX3k1EFU6TtEDe0y1
IpA5j70D7J30P3QYwglWXQrcF4ov+XGBDfVVvIxYN02+QxsbebJd5vuVoZJ1sg9d
7PxWJPy9LRveM2HFo4sL4psQ1/XG0uD6H4whfUA1B7Zmg5yW4mQBPruSj35+DyGo
1vUcBjUphUlUq5jWD/5abjB2QPYg21TqquSDZniyJACLzF8zhy6qFRteMj+5QzIO
ManoRCi6FsmF4JjrgpE9ZzAKRS2Rp9xwldfxpP2fwbcTg4hUlAp2f4po+2TkJSGY
UsUz2sZNrX0sUCNPZ3njjcdTYF9v7tf/i1otGnD3AzNAQsvLkoJCRO2Br9Uqnkof
AQr+W4AeaU4HSgK/wW9C2K2HcUAFocDCx0SI+1pnhr1d/ajVc8zvS4fnL4/KCZta
9yOrr8Mt0uZcFzIVdcWw5WDDeT0YAxZLv8sXE7uCp5gGShn3DkGf0+mja4L7pnh0
3YCIgdrQFP19aO3US7k67Xw0ef6QZjPzs6KWIEBelp8RyfeQEM1gnlWnQgCJQM9Q
AIoanraRGvJ5vBo0Z8z4a2KyPue97W/qaiSGVKqeZ2g75eHys6rbBXrzYss3tv8F
OKbi654XmyDHnyBJUIkT2XZ9zlV/luW9+gAIcF3cwt2cY1sKujLrzs2nlanSk/oE
ww9OxMVv1HddT45nZoYkXYtI5UR1vUWys6TCjBZmw0xgMbb8G1bItfR/P7Cu0ZJr
MVcdL23KWh2jG3kw3Tg2Yi+fKlPtG3ie78jGziJoBOl9ThIc9WWZ22XmY01GgX+t
Xz4pbwjGDqiCFQdWPNqGHKCDssIEDuuhQaOxyAf00dfVdpyIB6atAXWCVvhNcTJC
u3RctquIVLgu5PgCQe+ipfh7T4OGjmBkGFJ6DraM2vUwhPDARqUHv2TAeeTAUyjF
oA5GeYYZT8LP65vbeqfT0Bw1/XNEOIJAj+IEzB9Q/7UjM/qqzsNBdFAyp0YF4VGo
Ok38LbD6EXcn2vDbG14hc5uG88tQXglylawQamUDfyxkuuWCiej76sFnxMBdGQJw
fCvgRdG4NABccGZ7VHMEf6/E7uTf4i6NCJiOaJKB2Wwp+e//TYNOm+fDTVDaVe1s
2RtsMpgTTu1SaVZv2bRcF8YwlMCyJF4ZIhynFWy2kt0omeeWmIZBkdySJ4uWsWfc
MYmNYhPND16s+8Ocw4vwsP5CJCZnMZBm16A+9OSio8a1PMKeZHz/L7WYsVOKomnU
I4nEyBzTcnwOQGCszL6jkzT8niid2Oyv74a0AqG3D6VmiV1FBLn/k1wVbBoo1EyK
nCOsEpKkaZ0OoqhKzmZJSrTCERYcorz/rhnj/9xVF7c2z1ZLwzo7wZIkRqlvOlO1
zUuY7aFBv2AdIpu07tA8tvnZR+faWlMLVhu4pmA2kRWGkk6QThGxd90NtKI+ScSg
UtGl+N64zJ2AOLCTcqUth7FYIVsDuNcYXfBYZWb8ui+Nbign+uPmbr3kubT4MDcc
lOtZHyn5RBxujsAoQNyv0hx7iu59U4K9Da/BEQoBn2BwYm1XdmFL3P3TvtY8ZLDd
MLBjzjb1EVMwvnzcCq2Gm7Jwiqq/Z3k7a2pq71vLcxCp8DHyBIWlnkeqzC2JsoGx
5w40Qi4uAOCXRdQTxX1GnX9+qd7qxRT7fQJtxBTMfel3w4TKd5SGLBawSJ5IFJew
8/8MoJwdJVRr72a6//RGfx2Ytix5MpvH4HyVPOEaol0X3j8A8aD4on/oxgE5mgx1
7Sd2nx7kg5Iu3ojH0ASbAPdsz2q9iv2agylT0gKQQobq9gahxBIr2eUHQo22pIX4
1sG3+bbQkmfc/5IiIyxSoI5CwgClFXMj823nJ5b/9LqCN9T25kwDTkzLTQxTWXkI
oJjollgCGCgioHn9PJmV7DpeoR+I3l7Rb0xOpm7bejmpR933fGkkgbJpm3pELopx
L7NbZFnRQMofI//k9aw+iOUZZz6vBSELgUVEJ+00sD0pe8KImQJr74LqZlclxBWZ
/2LVPSiJJOuC5kMGUG4r5eunW3WNjMMhbTXXAl7d4jIketDfzTJWNNXDoPaE3PU7
6o+scm+10rgxk9qWdoxAMg4jkg9xQTObr4N5lSvEniKNPYgMg069PNGUUngnFQFP
+3JwyirU937KhPk9/G0FVUK1eXUEhA1aHklzAzJDiuS41yvlWS7C+N6qKj4bFyk4
5T3zrBS8oGZXPUa3gdtAhIi6Peha3LGAvbJsgijeda9sAgspBpazY0creKBrfnCt
8+BOjr5yvp51DRP8R7WI+YRyGBvoDIbiOtSOc04oVOmywuH3xqyuksQVGV6VrdOc
Tc8YIBgjUsh/2GDGvf2A+qyuGw2URLCsGjlobdWk7LCOXLTzcsvrX1dO5bsY+Jni
GOAPDXEUpCbxhhXTzTf1jjmnri4hMTQpYLhEm7CER3FZz9kKAafSW6jheOCOxTA/
8jvSzImwg2LZhumPN2VwvVn0eoY9DfWoQyTmorvIGhHXyEkjYLh7FJDRPI8NMxXy
3v04JcgyzNSJ/cy+4OED1Z6lXgw/IKHXlm0UfjIeWc+YoyG8AYDUM/keSwE1b6B5
NjczeTPAuLfVBGLJw746k9dEHUiZTTfzJQ0g5rooNg48Bw/AVPTHmZOwIPkQjGGf
OAy7VE9gAnC/VosPU+JRo7+35osfTNyfrzbfcKChXo+D/GXey8QvhQjUAMWvgGrO
a9RBj8U8SrpRCdU84truaUQpUhJSoUtesKd6mmi0OHnmyIwiQYAuFI7iLRk0/itl
/MZ2dGqWPxylS7QodYF8XrICwSO6fxdaH16Meobe8fYsCCjX5nrn47usJk6RYJZs
KjeHR7s087G8hi/Kk2TnxgciydIjj44Arsf0usjeS+dNvGw9h/40BpswbjTvElDv
743cMVev4P7lmnkjoGBES/hKbWE4dg4P/U9G5VQp3f6iguSLeudwDCcV1KZrJoOC
sU7WxU3Z/b/4HPvDuIKjjo1nHL1yjH2FnUu8q8QUw3+sTvbD31CNnPdBuaoDYKeW
0XrXae5aTaNXX1ZqhFnA3z3KRkfk4YnTkDfnQiA9t/NBygjswYpvKS0lewesS+Xv
l93LIxRyH1fPDOUXSqje/3DsVKSPe7coE55LwZyJkaFb3bNA1CoNc/f81AYIzZcC
HgSV1ANdaGgXeGe/kjbvW5k1Llyo7SDYS+ap4K9vPD8AP6d/piO64v9VACrdt0RJ
RbTBIUryLMS4XBBlFJe0Upy5z0RikbUyiELPDuq7l0RHiK1dEoHfHpSzEncXM0Jc
NLTy7hW6j6p1F8BCL79TWf4RxdIQ5GeCUZI/ZJE0lFPQTbpHpZBwCxzAtAn71kyJ
yjL6OcDXPJ59XnptCnadNi7xEHbIKu+JcAhF6LzReMKEv7g7WBwz+8afYlhfnSZB
IYLSeeHI6t9CGimcmtgKg+pjlbvKKdmoOty6COD4lAEGj6Ve3D79pTxKAkt9AYgy
Z3AK15EM8TE18jFHCFR32eru2JonT3i7Ocl/TrdqwzQuXw8lqCgK5ovDvm9r0VDN
EYFJhmz9blWIfdtbCy4wEe+eu/kMl15Pe9eB7idFaQZa+984/tIu6ebFX6YBIr/a
VMqsZsvGOAPmR7CqVt2i4SW7M9lPzFRjxM1G9FFHJfedn8an739n3+biBFUsQ5X5
PIws9Z+kQgW8dMEsdO2Ih3Y8KLnZS9R7AKAy/q/5xnGC/tiQnoWfLf69ka2rNah7
pqbbIpTlwS+vNRP8JErERMsBVUSxHTx0ldHzy+EC9ZqU/uy0KgC8jhAZddSi9eHg
TnBF7hSUMHl/9FxuwiE+iqPdF69uTjZawdUxubbR8mxEYbMjHJiPDXhl/b1Qxim9
EhQ0/9UoaEJJ3XZMIECPnWC4Kl1COtCZNNhw6oJ9DRPTeqvQh9czuSGROKEgeSlJ
aZeOPRxqZ2C9MWc0fgQaNd1KQEiX5G+xZIgMQaW20p46fkQaWVP0/mjcBPG8jiGA
9xzv5Lw320gAn2/OYUWu/Qo2Fmr1K3WNrY8noOuz+obrjbeU7jwk5gGL9skx7VSN
s6e1sAmjm0lMLRlNpem9scUJrTAME9zvxMl+wwbXLqmR6i3wTVL8rZFq4tbb4zsk
biQmm84RpPAJmMKWPnoLPjZHVmhk23+6N7rTRSRJ96Qi991og1mmAr1tWdd4z2qM
5hxA3lmpd+5rR1hLL7q+IPogh3EjIBjKexwxXYRbMNIdw54d+MyZAUwA+mtBUIW0
qAdjKu4xDqEhiqk3KbzgWAGq+p2mkFo/vTJCq7W3YuFLdxR8rHKzEuAqXz5yUMvE
tRsTRuC6zHtOdPZVconkDubQ1lyYzzI65aafk8cd3tQaAbcgYvqNf8QkZnQons0J
M9CQQXMPKkt02MYipVWQskzmV0PaCYHro6nTk8e0NiBqAtgHXDwxxNjl/R5c7HiI
28uWVR0ukiJKBIEiphJcb5o1G3fkGwcthDTE63+iYHuZInENxvTJaaoD8WNJYmAn
yNVJ4Pf4yFPqYgQzRhcsJUo93l58+OhOPYmZTKKc46JfdsCWd89RUdPNCrkikQd3
IEGgUsxBHgsp870eIlPxci6myUdsYatcdYoHHgN/5eko4oH96cXh0SD+9ThqurBt
dWljQ9/u4NIU0xBQjiWmydo0T31Mp4lMz9AwVzKMG3QNeGacQotzqpW29EAxoPXN
ydTjRu1swRngTmmtRoo8jxNNt05BVWcBw0LwtexBVnwmakJ5JXfIsQ2YZru60M6V
jspZFJPdsZ+NlVnQ9JXfD361XJH66Ct9sveEe/m/J756arQ3r8yzulka1WBk3Udv
O9vwBd+nz7BlMvsfOtS1TH02PvmjpS/2qMIZU2exbILwY+AxUbKz6yu5xN6GAS2z
hNSLQvbi/0/WRO/edQLmO82b5ICNWShh8PCCaij1KKokvdPojGGZrJ27PHcivSQ6
/UyiunjAxUifdCbjaRn3GuNSHGc6FlG40a0X252Dwzh502eg8Kio/Mca+gfpOJrc
6emhoFH7W/44VzaVETKw86K/D5eYlestfL40IoVtzR1mcqY7BgMyRGg0o233t0Fb
KrPi8mKL6Ot6lWSEHIne2MKbe8/Cgm6ipSUhOKBwwj1ViL33w15geGJnj+IfdeaD
AW0gZ2sx140CtAVrbp+J5djkeGELsR//usX2/A0b5i51JGXfZsqMWie/HS2513a1
xsgBqv9r+HmezaWDHRp7vWDxBUAqYJqj9GX8wbsjpAyhh4FuJ8DnTpZB3UKr/xLG
EyCV19012LAoqbHI3FqPjz2raERMZl24ojlI+0KYaCOEyyhzxjGund+JKDLtVJAk
pmqTnAwLd2b89xw9zruoTTij/9ZJRLgB5f1oj8YitHxfR7SaNjoHTotIE3YrunyU
X+W7BRELOZId1i52mJbob+DAOed9aBJ9xGWHYt1cnrJ0m/XRerpPN2DmvOaMGLTt
h6UGNgit9wMIv8nAvw2xbdx4dPbOWfl+84lO4RXLV2RA9vyfhV7qxwA5aoCVtXR1
fkT1JpIFmHEELkUtVyw3ukvJ04t/5t0gn0XByvREiDydouW7jlzCIBrKjopsgZBb
2tE7yX9D3QwzfNKPIHhQkW+kJFifJ8o1DC831/6QmAwyRTu9CUc2rjwxN2lYMP5q
qbB2ru3S/rjSMu2N67HLviQbIVtjzMS8+FsXyTKaM9T6027f6s7aV73G7lTw03hC
pe0VbT9Ly3AMF+yNb4WRTdYTzIKFbYcCOoIMwWgMKPQTze9mBHLJonBoPio/0yXo
j+PKQIjV5/+tJ9Sbo0yn41WjeDSmKll7mYbwx+JT9gbj+KeqtVvauw+dVZ6SXwOE
by020kLuDSjRCwOps0LrY0gP3qH+Sq1P2VQc5ohLEAlgbQkI0MSAJlgPNwlx+Oma
11r/IdOaupreKd6Gll8sYpXgbCzzx1zh2AqgKF+ROG+4H5btB2g+fMeLx0vbk3gy
K3vq+HAWlwysiXmVogpM+szpscT4+VW9aqjx/V7XDva/xR9WG/TVfZLxz3ATl1xG
VGbRSFgAsByO2mc0GJJxkW4wKaAKJpQ/KN5t0451dLWumqNeIGL5ufzID7ZsEgk3
10w59fENc1PMT8kMNxS85L78YCxPskcIreU7hbO+4RI+VaXb+U1Cer8HjUtSOH7V
/mfQfJvuclVlSHEqYyrEqtxBPFAVbHUt40j51BQPwqtmh7rHTewgjaDBweoOva7i
7ds9vKghMU8M7HhCfnQAXRRC4v3SscL1dClekJpbzI9wQkYdx2Aa3gxSOHOSUmMD
jAYoFievkegBg5/Nq0fkfAJkRFXA1pmP4TwbEm8fv9A9jGK3ANRnGRHoKH/Ijw/f
7/JQA7osxZROAObMHAu6Jmc0cwAKBIhlpSsO14v7cRAtD8fs/RBw14fzxdMmL+hG
yhckkcrkUIs9Uk0vSnD3sx1xbmkNC0425BWNrdow2U2dV9OwNvauWV3fgdnRw+Ci
Q4bBbdvin0TNdYLT1BZGe1bRZ6opcBDDsLt0iigSN1sY5rff3JM89J7YFenVrLOt
5ok+8V1xLSF5JAuizFIDTzRR5Jwzj1DIO7GZ5FIpCeXTsoMbgApuf0aE/jgrW5hf
I3N3lDC0LE7c4aufialVPWBJz4ZIZBwdli4o9koGJzkiV+L5x2DznoNPegjdUJgd
Yj9yaHHTwD/OLm0T5QRKbkb5koYksZJc47UWIHRauIpz+p5HxKU0PDTt3+Dh71Zg
GUC/3duqEuN4bVLHW2G5jhTz3qzwKuUU/mTZnVQsg3FxEQiBh0g40iVZMhL0fzl9
DAX+J/oGDE/yMQdWGTUQxtj3XgHzTvgtNUT4wvH90RRL4lqCcSKAvXuRnqn3xW1y
+OWLQdoHCppHZtPCMdRSyB/t4ZylO8dKllcoU4o0TX9l/v3ggliIe/g5kg5kMKVk
0yZymoWOxwy6ct+6a0Rf6vxjCsAiF6vUNU5t/Ny0uG1QArL0x+yofb2acIYJ4r3N
IdA63yXXRMMEJLFyyA+aekGWzBI91zd8AvNAc21NdpcRBALjzuBN/oh3okKL8V9Q
2YrOkzbV7DSmcn2PHC4+kF+Ee7iFHKSE0ID2fqXD64uCq+RIsHE4AZ1TGurxQUHv
kW5Qn8x+ZHqoLNOB8ZKl9mwGbdH8ETTSnK9cNws7eSQu/F8eRz4dH8UOjcqawpXB
SqsjvFJ5xb7PYuXqR472Ad8IntHFvMpEcMlZrQNtAtN0LGA5KUvt9ns+qj9t21gx
9LbuKbCB2uVAxFvfNQ5miqUsG0W7dJHOwCYcdDgR2PCN2jTmH2B9eSiaALafuHeW
GRmn0op2T3ckzAyBBTSsCAMdF2Y48FZjPe/yzHOW/XRrViPC/PYmVa/HwrLs6FpZ
62MXef4a4jaUI5ucCIe+OogCO1I2uaMAVnQnUobzL531hlFflkVb54/BNaoafTR8
sd/1gpLcJV5fF3yq6yO3ql5c+YDAGHW3JK1M1cfhyn09Y7XdAlPhJBU8dB/cieAz
MUCwl4+fSuAMXfWZA7JB+LdAB1qkX2ZZVzZDH0CS0VPjAC4ZBPcOMr6VVyBAwz2h
a38vda42n/hUNd4Uj2RZW1+4axDj8scIkup0GtsJZx39zieLVIEorbktDub1bjUL
KtRMwfXtt5gqlYGClMtlkF8MUeJnaKXtu0VNBcR+cVVAlBP9kCjF5VQ57HBBtIl/
un7agFwOrbMDwpZuZYbXOuu+kah16UkSseT6iJ6G8goebUi+6rhTeyDWlnvUFSEE
V63CkEAidrITi6jaPflaVEMnFeJA7CtvKBNKfVYjkW8DVTnnw/wg1uaH0//IiQFB
msa9dFi8pYrA3tu0xxg277gmYG6vTiB7HyCIegPFT/IGkzrUi5X8OamtpevIwv/F
cO1YfeSWXadvWegsaRz/ey2SAaM/qiQ4vHtOtdfHdHpmQPM0Pgnmxa4Y0Jqe9Gta
J7GAbyx90ga/yG2UYyJDTdcC7Hax2wHCpFR92220VHId4UMYdEZ/tL4b+Zs82DnT
+mbyjk/G2hPfgFbLRmk2edPss86N2a5nBOfQiltrJtESRjXCkUaIZ0hhTWdstuPC
uct4WWmwNghB3WWDyJwRfp9fJrODVCs8KLcPw1Xdlymh98myr98vwBzwHu0FtB8T
HolGvLr0c4Uf9cDsx6CYYniRvM7M/dt+pSKUyn00wT2QzJWfTep1BpMHatigwM3I
BE6e9vawjhb+NulXKm6UQtXVmKKPrkUS8Ev4Cmu1w7TnTc1ewJz50I8A4X670qXg
J4042yPzt9kUShP4Vsy8GK4udpvWfcg64bFKH8pEG6fsfsdjZhtWwX5BGtPR210V
udO/gHLj0LOC/EdjaGJHyrvgBQNXCbwbv81xuNY0HnSXl7K1H5Jnm5t4nQD+wPoh
HoDkktK8OIkDcmkxja+K7tIN8MaGtDy1h79Eguj5vZ6Coy/06Clvm37PE6zFnmPG
9L0nsVkZRrhZwj3t0Bs8WYztlMzTS0tEdzqwnYM6GFYiZmpa5jJrta+ruyy2DHeJ
zoI9+VKd4Fc1/ultPuMTT0gvUAZj9+Z1+C0XkY1l53mA7ynvx2Kfv2a441KGnFwK
yw75+uTsF3USYsQpnJJFoytkUoenXv3ojDkpWzQ2OOPoItbn1hUqUnIzYlf6R7mS
+B0ISlSQf1dECfZaZmJvjx5mXKimMrYdcLxwyEgzxbdpWJshX5AAFyrbUbtpuxnV
IsMMAGEkKpfcii/fsnopZUnodx65FNlOCoy9lTOvhijIKEoWLRQNkcjYTYq2+mZ1
x4ET6p4wl5R1ZwLRJprEDyoNQ24yRxg1b3qRR8xRTFDLMT1E21U1CZxv2ICGnK9P
q4veQygMwTw8cP/LjqM1Sjtz+w1UEImXtbzWZvbC8s1y+5yV/XJ/2NzfTmzSmVSy
FZjChJQNFkRI/sn7mlkRJSgKXj3xlSHWV7PMOXQTC/JqaX9uqu3I4rJyJn8+b+jQ
6ID8WqO/mFLbV8xjik7M1r3P7AjUVDdT+GvKcCiiUwwGBTJvLDPoKN/71wFp2trO
Baibz+9nSWnh58R5Y39CElReaIXI2qJ0D8ca/P0j6gwTI84ALrMjBnW79IaWf4mN
037/cgURN7TRrswwuInJheWy1dJmKmxEKcWraN23lj7y8bIxmJOuHSBnHf36kGne
pRgFoRj/dXFH3O9zxRxQenMIontlUgqBEHAexDMPEng8elZEgskMJkSgPFSN1L/y
o93s7qmfLZa8XrPiE6O5VOGCFul9rtUzokwulj+Da2me1oOcwEZDN52Lw2alZFtX
qqo2yjXFlzuiDAFe8x8KoDwX8+79sXXf2pypj/EZr4j8TWVnMrmPWZMmErsHNC+6
Tqek5dZyY2WPPj6HM1/5xMXqAH1k0vUOLTHAGQcNr7e5ioXu8sTN/6tQf0LF79dp
YxETxc06D/nk8MiGV0Vwae8DU/Fm2b9A352Cq+NwlKYIDUC5askcKWANvOIBj/I2
lAayD5jKTeUrnRHo4j3LSQg6ye4VgWoxWFhb0hncqbQN73GDHH1cUdBj35iStKVb
B6S5OEDdB5KRSMmzLHaCqDQt0n7VCQmYamLrZg6nlTkF3K3mPz1vizDlgzP007PE
QCXB8Wct6GzWkRmcam+3OuwOZfmc/5XXbwKltFIss2xgWbm3FeiXfK9EfSMbmngz
7rjbHQYjdPmhgrrl61LRmcdFzMnJkpjhDVpdzYXTfEmeQJ5r2eEy6++5PzZkSZA4
wdkRIwrllvwysIqt34Op8xxxgSaXkKjCI0bxZ8DUbKN4GAe1NLFUJDGbXEjyzDeW
eZTQda79/jhPHO8HlVCsFj7ZnUyqd9OQ8NEm8LKGkb9Mgiu107UQBRo1eDaVWbyT
kjvHuHGG71PjVLIDeIG3z0hDJqsWwj6KMEzdDzj3sJEYi1LbGW5tjrAfAhsu6BRu
iApc/MVJcwI0dtUEaC8GGSHeAHWssdJHLlF9EJCiMA3YByi/Yxi7VpKnKYE7VcuT
X954XsAFkR55eYjS/nZsLRGAzfCxqRtJYWHM4dS0PTitgupmyC4IjifCCYM64L6a
pFsSYnmoVY3Awr5x4Mfx9oyqvzeQf/WE4k8ayh7I7lrp8FvSu/j1jjvMpuBrzmXi
aNSGBCCsCxj3YY4w9kCctQw80R3vLs3aR/CoNkTGSkNrc3sYptNXZZTXkAl0phB8
NjM9AJPe6ZfmZ6gctQyZuOv0oDBzWdEdrjhrS9zXRTciw4I1CHAc1DZ0RnHx1pVo
WMRD1PPvDxbOotwo1YiyZl9LeHmClz/ERDt1Qd/UZzHsy13/gc7Fv5AR3NwHcQnC
BygdwBXSMffZfOuVm5KQFxm5qXxwU9bK0ApL36bOg8wnVlNYl/pRzcg3pMdY5SXX
dggTGqkL44Myh5MXYFEZxH65RidNcz4Ks89Hz2fySvcidrFZ/ycpNagRlAGTdlIx
7Fs/ey9e8NTujQQsZkqRSEcyyvzVEhrIHYzDdt1d9F5Upn6TRW1cvL6BwM3SuSGb
Lg/gCWqbsGM9BGaKO6UWptWfC+RPPPozz9017EISnohsPnY86t2FxrXkv8FVBXZf
OLci70DAQ6WTS35bPzqJbkikxNwRSFrDCuC99dtlGx51pwksS9sXDIy+6fjWwzun
FnCB6g2xer8rwB1BpDWQLisOnBM7s9L6hJbEF4BoBYfeSCk+vL0yRKTvuN7R+Tzw
+rJeBlHLenQE4VqMBIUu0+o3MPSmzrP8FXU+L7APd2Q6bqA42IPXJsTaOtG9jWl/
PRacSlRBACuA8xNVVcaZ5R87LTR2/+guBJlC2Uc03JjzAunxMF+yQhKAXmw1FHwA
PbMU8Cf1KVrplK8z/XhS31XOsXLULgfSnHRYlB0ebY2DYU/uqr5XDonz33TwZHC5
Q5SDGTdwQGbvl14/P+66YGYPVegEanfZ/BtwZMVHmInJDKINbCZrbUnHmsPwAhZd
1SN2HHCYjXvv1ykP8H7C4FETagKE2eUzPjm7gxt4n8fDR16SYHxH1dVdfGTJMpw+
AoptbKA6uJBN2IUzMY+UZ6BVNKunNPmSFbu5YH5pXS+WTotuh75mEfa53lm+IJ51
jNxbIAYNenigLfBIPxhTVPfHRmPwboet2wg5eZ7Twz/wJvmU5NTPXwUoAXKgaVPw
Sln1p4bXzP6eAADo4QGTDCqb8e0j5K3ILD8EDNq2geht5BdrHSHlUs8rbgjQxdxy
ussffMaX++MwhQquD2Owopc+IVTk0vAglk3QFfH7CbaaHs/WOc+MjcB0rMJFvbA/
dk1D+0wpYMvnQv36RT5I7nv+dN0jgDkbC+jKy+M4rdBxaWpbfHVSM1AIyVZHz31g
ljndOgmzHwcT7zAXjKHvGLYJjKVvfqGsdT81VQX9NXiFULn1qRIA9TEVtXvWX3NS
vkW4stYzQvt96bquuzk/0hzmVNncd/rx7cqhuGvkDihKj4Tj8W9TYuyJPQonDbue
UorcVq+n2nB5imueFtZT05VmYXYe0M6ltq8CFXxBfnkg4exMPxAZ07onLc+8wlT8
s4r/euBLWTcgxiCMKqgcVpAXJAqFnvf8jCR6aHrJi46GLGiNO+SbrT/Z+BrbAqGN
1CKQ0xzyz6agBHkobBIhbx+nGPRYUI2PQwmridNyG3gPgCmzWsl81fIluPQqT87t
LcuWlSejW+FvSeyMCT6bQvR5UM8NHyFaTumttIZV+Of6D9cAoPpCDYRLzbgec2+b
wG3RIa72aEpgtMtP/CnSTS6nQynHFuKaKgf1sdXq5ngtc2E/Ryr5Pafq7o2WPmlW
hxlgeKKLESVvJ2HUKCrFtRxMS7JSyY0IfR27Jib0gX2qCjwzuWCZEdRgGNLsxQ/H
qLQlRTj08wljLl7Xjyitpo6UEFUODb2gYgFiD+1Ro6NkpXtA3bMM2eADkrxE02px
ToxlRDbiu/I6p1s9fyHPcGnxDthHt/yQyVRrAq4d0Rgu5vBDR5UQYnxUkoLMOOay
dTGpMnZwo9W8X0tg47KrIO8+NMB0xfbDXYKlbggPpezAFGdqxeyusDpZs9HyujaZ
hsTfUb+efutgkPbnMrjT0bkF6EATv0xf8/lvp+ogB+slWWPPuESg9T7ZD2Egper7
c6jNZQ7L58usjLwpfYbO9ObOgp7XBKB8FEE4/KQr5EGGQKBORLDBuLDav/Fl3Lw3
phLyLEi8s3Tm6zFktobXJaMToONg8Sa+Lm2c9H0yOSDYSfScBJkaSTmLZkhZBYXD
LrtWOkjWS62/M175BhQ/B4ezmWAZmfcixTfT5IGQn0pT289wGXHrSqLJn6v4KXFJ
lSp0B8o7tlC+hhHa4SWwaRg9/tG86rtyc2ZhZxrC+pTCgk6RhZURwry0v/ZEbrgH
VExVwx02IuCfaz7OXnOrOwMcmqHMfyUEaolNyMEdj8Mfyq8qkocJP4saf7eDiP3j
CIU+6/ZV/PrVZcDcO4WnapsGzkqIR5VidoCZ480WdrI1XC00qS+Hgnz9ZLpD7Mlt
24s8yRayhBbTl6r0z7xGEYvTSndspGtgoqTVC96mfDilY4ihiXl8v3ANwzKSowi+
k7b/pmdXe7Vfo4XW63UkQ5cAVezVbEIuIBX2qqhTjZf6FjBYjP0vP5yK5Mr/mS9C
+pS6o2vmVkYpedhYZY9lUuhcPF/2JR3rJNl+wNjcljg7AmXUnny/lJOvjTGgLwHP
4bHzwhdLHZs7egC/ot1PLtE51QjIcMSY4zZ0yRCobAqyx2lQxQ8+yUN3xd9K3JVs
jy+ZxKPG37PFAF3piiL8LJ189ejFKitliwKFZjYzr7l6GgOhtHgVMUXJWjEHwYUd
yy0WbFWNTmZcda7+Ynxolsm0uwcPhVovHj6tFJNyZbYNQAL5kI/iaTaCnbzO1wB9
AOF51T2nxPp7fbbswsLIsha6cVGxqLoqgNDPPDl26HQu4MtjnrRYCGs/eqJf8dh7
JGowg/ROtAbd2Rneul/K4JyoK+7P/EMo8i2uVCY/r2AAyqXDIVtXe+yy+H7oFQJ6
o02uDDbUgCIuTlJwzDpZPnjOMTP2BM68cc1jFJxWfWt64xN34YdRpbxUwMn3DxgR
z3UF6lTQzY2bouXTyNI6jY3yku0/Su4o0C6pva/jbWkRMBs1WP8roL1nH3cOqDG9
dSspJKvjUdfjGL4lEEwvx/8/SCXRaXBbEjdUToJSSU8jZYmHkela0oLKySUFiRxJ
Ogspg+GD2kZisAGOUvnHjs9hDo7AR7XSQfLnuqo+eNRCAUyXDd09Kw94MwfUQZtL
2s/pYb2S30lNgYIuXXLnhL2iyB4lV0BTGe3YyZOO7m6p8dQCZszHpUjti7rrzZb5
nvubVfDRcO+cen/Zedy69tE4xJVrGzXcHDVHhM3jPblJIuHmM7KUVaPnL/Xi60tz
GGhfp0uif9lXBsQlpu5NBwS2jZstFX/mQ4O+HybcJWmMsBue+3yOf0TfL+cij1dM
6xiHzkRFq07N5C7zLSwytEotHnrlya1fibc/I0oj6s62Ey3lF7/vGtJMONWol80/
OcqEEy2xn+taz/3PkcOl9jMtc5hWURoF8um/unWFobAtADqkFkDwUYSatEIUg3JE
VIyMuk0Xc6zLIw3gvgDpNsCpeO8IMElDVQ6LZaMatq6eSpEkrO8X9Hp3ka4Is67R
1ayQyT3mxhCU35Tz9yOMT7qUR7k3U54MhyNGBFHfnf9SZvFg6Jk0TdhaTIjCFvht
/OW4vfdL9nNNzBQcnJlQTvXIP5Gh3Q+5hLystIIEqXump8cpir1QXfszeAQxNeaN
iDYEy9U7/ZH+zXZC3Y290O1IfsZdOzzreGc8DpkvmULP4bjKdyj/NoyNbX2f2edm
Uy7jYBYgQwirTw5xYnj+y9c9HFeUiKzj3CjjVw5Qj75xkzbj6pe4+oma3OpEErST
cFsC86aYUYqxsctIRbOMT/u59CBG3ZR5nSd1kLzpnwtdlntaMJd8I5AxAFhjnwaF
UKefZZDuZFfCFP2Znm+gyGNBKcwOkBtl3rp8Lqr5+ZbD+kI++S5d30qSRSurnDX5
fjOTGl5wjuz+o1xZb8KS8nbfejbLE6wiGwGFdng94x7WMbai/jd0CjnrpkAo73bD
3p12kM5d5lzJIQFJPRDdSQar9gQXSUT50E8fN6+ND9h0RPyv1Rm4OMmAnjgpBj9Y
ABxctTmRct5qnBWJkLcFTxKw9dbA1wpd2ZEWdH71nYLoFanfoqXE/NOKirnF4Yz1
lvsZ6Ooqvgnggnq4IzBUwQscGk8trSB5weIMhpNMS2yzassUvTUXtH9bBxsVPWRN
AKVEF1gDkH8XJ/+TZImgpY/cFBf6+lnEg5MnKuyYhyvmLTF+35sDLJIcLc5zhVeV
C2GrgoPj5wnUsu6EdrdGO6xxu7MB8ml2QQ3p5RbzO1gZh1z+NA/ZD9r0G0JpsuBc
3chnlEUsXVjkh6c9nrXS24yLZ1bOqApP36V8LA4UmGCLTFzeEfwzBE6vIPgoHJve
2qwJsMfM4SDnUz+fsmYcf7TqyZ+0yLNSaIL+sP0guRcRegnBOFo0KWyYMWa/dUTW
En4W6JOYu03zm0TIx6/lhyj4T9oc5IwadJ629DyQ7CZff451DARCWJhNihXkmmXq
a2lmUAb6h3f+bVWWcZWxy5znQwqWIiOzkIB+IDRxFxT6/oSxVgCuJ6hJjeO12Zx1
gbMfH6mzaYg0Q5qCaq97BKSUym/g2ZlV1pck7HzFU20aCryvZgISCCmpp5kvRSKQ
w2BUci3CuRH4lwkvm/gRbiwxCIv9UdrbsVVgferJHuG0HCvXh9x9Ul2E/HSqVJs0
KsNcdKSmpK9/o8EWBtkaRMGcDnxNiTkiY0xm54uA6aMeTl4uRJXvpokoCgwnKWRY
vWlNtdKeI7618K/QMvQGkNWkT3ouXXIQwtV0c7eni5hNFr5SnkEDK6at67rsJrXs
d9jjbwmuUI1LX+mjrZlqzeHqxXrrhI/mKlX3nY3J0T8t+vPaxAs8HMB7NY4xgBib
yfS7qhwVb6iMLBCZi5Tb7UK3FuvmLWsDzmEiicPjb+yG8FJcOKtg/GJzf8Wolv/c
7MQ6/KcziHB/v15u06OR5eQjuGUMmYUpMXor9e0EfdYu7bfIngaLlcYCN5ip2CRc
pFEJRe633zCXNXMbshosK9MdZgFayGgvkMU1GiSrOVGQkyXgVeH3ZjNJLfFiQJ0H
ZS3PDuSO2g05M6WbjhPfohayPWhR4ZTT0XcD3ldweV2nbT/Yhb+HH858pjpMB5kK
nTB0TU6+71IrBVLK2/6oWOAtmVrHKbumCM0gW94l1f9O12/AzQIHWDdaV02dQMY3
ryH9vnHyipfGHdB1icAQqFvGLU1k/ai0utk4XXHwdZoKir1e6GkrB0PLWIKPtQAn
yw5c39CAAJzJy71D4y8/TepPzR1Cr4fC9ia7eNkHPnJkNDUDIsKWXEd2UwFvK/ED
5ZqUqHjoVsf826GoBfbwXyO0wduT6hhlzEDfVUmHiu3xqbgMmBxkuL0PpUhkmYev
uosw3dnRbqAHq+zn3pU1cKbXufbbCk6sKP/4nI8pYmgrq25bdRBNF8D6Vwhp0ibA
FDYz0i7T3Tj7XqEagl3BImC4uJC4cD6ue68T0pNPV7g34Zv6nazPL+TMWvZZcK+m
RSDsH/tNto2hqs9o+YPd1LdC7tSbX4AJoMjWClFuAXt7kqK0bPchKZg5p9xzlFco
GfJvSBlYlFhGFX0BMWCUeMCEh/QaTt73WhZ9LRMzjmHTldIOH7GyPpBaXslUODU6
ITm9PlwdVnh+W270LtD2V5M+WaE7sREVB412fi3XrTXMssarDoSymV0cecMRJO9L
24AZ0S4g/Pf2SqA1+6RuHfa1STeNmH5OfZ3HZqjNtYnLucd3K2aMxWEnQAQ82TZt
0JD0FGjPnCYyCPC1W9ySFjQHe5lfQ2dHPUhCg/idGmMxG2boBYVzXpEcngzV89q/
NqzBjHPhIeEykVVumpBRvUesL3uYCFbXQuirIxdx5cx0popQ6e7Pon75mp1V7ByQ
rt/wmBBm8hrS1pHWKUcNJfWFmC9RuOLwsumZtq0GPJkyVq1v3an0hDQX3r8+/Ua2
GOZzK0oT6wurNgsrlVLyC7C0FiLDF7St6D7SdXLmUaYkL9XzWOAiPWAVpErZ2GDW
vUbkqv6cJiwXyXYINAiGyVXCSMadwFs00A4uYRE2T8y7Cx5fLUH4fojc7r02pknW
sQvfjwu7IgECumoUse4jhAxrXARVnOLMlwOVg7c3vpcNaPkLBZJXynhVVpfQM5Hn
B9OOPb3S9utBu+RuRQwejA+DBXQkk8dzl6r8Xa6RV2tz1gXhBeMkb10wtcpJGKeK
5ez5mH8tdTisprkgjA71dMGVrngYip4DFrDjbPf9Dg0Xhw4Fk8hGzxhvwiM4I+y4
e99kvcaiz7yyJrw8kcQXoiJwHNY50VPPWRn8Mq1X9JnGMpJAuoakVXO9Idp4m9xe
rU0/syW/DWs9CBqEwxPy1yxJF6anK/ny9o9tzFffZrEyL1KvEaUJtvbwaPuRcOl1
RZXuNh7RaquyvEkVCK69sOAE4ve+4tWPTo+blODQvuMabCVHC4TO+Hh6KgpMMoP/
9Io/KR2JrVLeS0I4l4Fl1gWmpu/6sGN0p0zsjhry+XlKn7IZS733dpKLqLdUdqDz
WEtqr9D+Z3HowMN71lwgMD8Hec+fOkPYi3mfSkuXnYkB65hRokuhNy5xxmNfUqGh
7J1sCZbc9yNoh7o4X/0k019sILzM8DQD3z54CcCPjmzjCq35yeTLl5zluWTGHBT2
e1dTw6yCgn5seW2tQ/r97Lc4vcwLmfvZqbBUPrX01JZugl3hVdDtnT2mSIy8nIR8
NHgGomHTh6pNuLxvvO13BoiL76FgdO6qOZul0fdNgFNmV1v2zJ3U/TEmJeZohMAC
IzTZM9dM4QptYqvSpH0Jl3ymvA/jFcFYMKw37srtf50Noc3pQTX2NBIPiT5GTsXl
Hn9megNDmvDOwse/o8pTO6NhnQy4k7DzSh1Gs6bilnZR7o0zvS1JF0kvsNppH6ot
JU3/S4W3k5GpQZAvPMvE5YfEA+A6luKERKaKhgIaflrGYJ4cP4wGiRxrKw4n3BpL
HGclFO8j/w5pWGqZQyrGyo4mK4WPWwfReskCPozCMlgQ7f8PLceqKXtKpFIcRYeu
KwyI4tnjIK5x+kPLxOqamd9gnIymbnM4sqEhXv/GdN7v7DTMAdT1C3Wn8VczDkfa
zYicKg3K/JdeCue99Y9tGpi+vFbUevokXf6rWghJN3aV+zVc+R4mUU5GgiT5Z+gd
VoDR7ssdk1CQcH8SKzgv0Nkr4s6+GjAntfh075Gv/gIg1r4fZkv+FDxpTuBT9BMH
31uUT78lU0LDdWoJFPZj80lUSH25d6RR29twM/ys2/Ej+8UcERhLiWfxXmYi/J7i
XhzC0GFOhF56vhskASHYORf60V9J6LsnKW+tksZVVBZKIj1NqE4sHBcskYo08nCb
3a0agMVzBCUAE0TZ+M9ZKdtVoKkvhlY6BUDJDlboLGyYxdV1kHTpXl6zcOCHgxg3
EIMqrcZKD/jLjy8Pn/QLTdk0yqF6ly2MfrC8uNE8fu2wxGb/Me4ue1+NT0YDc7Pp
hHZVe+uq0lR2QLjBqHhMJJ2KnjEY2gW+gSRnoNV8odqE8/NCU/DQbaKm5ZscMzdv
dr4TNiL2tzzwLJNLaRT4tzqMGazy9Vs7dV6+fGanG+ywYaC8H1o66SiPfRvE4ac9
QNjZ5VzXwO/H/ev/nWzI56ndR49qMoDFg1KGQ5tQIIAhYkXE4HxUs5oTY1ICQps9
TtBbhr1zj4p0mtjEvl90a96f5HIIeDCJtMSiiq3IqTQGcL7MfoaWc4kSgpjkZCwO
btR9oj33Acxxyka9zSU6Rnb/3qwZZqjYLUsH38Tu1STcS9yuuCcweaIefLN9Tdt5
VzXpPNiURVBlRld3RFxzxa8MNI8JdjxDqqmxY/4yYmlxTo+bMdqMs5/mfLVtwzh2
PEFaEDSXwsZWAkIgULuMTL9zdKxptyPpGqrpudj+4aOO1FM6/bnvO3kMI9ZRBLQc
hEx3LXS855uNVAZOKV4yQ75j08rXG6eLbKgdLTDwrwRG9gYNDfnHyjoWIfpjj5fT
NMtYufhKIFdkwtRgpW28EyKPoXb2XcwYxg+44Bb3zREe1tLAB9wjSQz4d2pJfV/X
3+ixm1fmEZIDtt80AF35GVBzhpKPzTtnzaTvnHzU99IH1ZFOrVUc3jDUF3lbNJMg
xFiPwPSdC5ySclnnNyp8vZm5g8T44GNkPX6jTc9Tg90iETwRaNbwyqjMoFMXn53q
MQnvr/CwkGqvfHg7HJvmtpX6C7jmbU5gZugosF19fyUYU9d3hPvuHSJfncGrj6gV
rYHO7PwKOdJyDEiLh3Nc0abjkKeZf9/R+rZIDKOuUEv5YL81kNuNkgyLYwkjesFn
n89mTeUqC6duDrB3dp1jy8QV/T5kiqr9tGOExf+gbur1uFTsW3DZB0o0PweeiMb0
1hM/QL48Tca09BDHsb9Dm9qUpmwNSWFo1H5cq6Kahem4t5NwZpBBOR4kA7DlDY4D
vSZuwSTEeUfm+yaKBfP6iofmtfo2j9L7JGbA2hAlTmPoefpnu9i7KGnlJj4O2yUn
HHk96TaTE6tZwLrA+Ntq6hZvoexREcelYT8zXiMifrPYoQCY69tP0ZXOZ575xUQt
UbieEcRAYoiZbZ8B90WRNaSAmHfhuT6r32SdDcPJt6yPiBCHZY/UK5V5lGqXS76J
R8r8qMq0Lr1vtoBPjnrhEuLDyRKMTfBT9zMA21gbyUoXXy0JPeUn1Hmnw2ulkgff
IaWYBMwNhphgkB+c/Zdomi9Y7FuUON5u8nOSg1PzsTZpzury4Tznmbi2Ix3rtu7W
SL5mGjKMefzN9F/oGrF88gTWbxoJ25r8FBI4x0l3d5+naQzexxpK1tR6DI2p/fdU
Xepgj+xXrlRlPjn0zNpMeUYXGi9HlX+ll6/7lK+2TgQK6n+IA8p4L5nQ4ScXgSQf
htCke3tKwcbnKLrekhW3wQqd+dD9LW2AG7lYiInwLsSPqn+x63pXTM5T7kZHG7g3
uJ+we90AQgy6BjeXfqVXyDaZGlLrTdsseu9r8t/3bgZwP/Ot9ZzqA8kvBoCgzlOb
XFa7+vgJx3wkYbxJnynqoD+kp33L3RXvUEU7WmnxgEXo9mFjuuOsqYzwOHRQUcuK
i2dCFzyYd727TsMS0h0pwqUUJr5LoBIFqZ/hdg27Ml4YvO4BUbuH5hs+roL+ic9/
aeKckC7VggmDLOyQ5rVm5oj2ccIzAKXATUKGF/vTSbwH8RUUpYPoYPcOMEpMzrxb
+ka3x4wK6OwKadGHwhH54wAyeDxRzCU0X5k2wUBPVMogyJUj13QiT7c7KFF7sAEA
wexfEGiMYYNokmcfH06U4XVD9sysEqwVJuuFCy54iBC/eCqQr+2JVC4zgRLsbHEy
+kvlgg0SA+yN95zrwWhS0l7c6OUkjPN7nD/0KxiArAUYfwioJbLfnzCa00fBbP5Q
9INWjkO1pDzNn497QEKNS0G1j+ajVwLj3bJNBMquOW9JrtL06XzX1UDOABafvL0x
amoV9L2ybB2l7FqULCbIn52ovf8U/qf+2wXLBQVkVeRhxK3L4ikCKkCzPzAHZWzJ
sd4qrOWvTWKOb6Tl8Mhm/1V6CgAmeYOlFcXHuJ7Dgqp1vWFM/tTUMdjXse0OdQML
sXpgUO7bksKtft7TXb6O21urkoaTy6rv0gf05G0FWjR4WbtjMR2vWHHc6Dfg/lqL
hlKEYnjTx5mQnX4s1UZ8USFqFa1BJjSdw+ehUWBcGVJrXOc/4CUFISXJIR8a7FhB
zu9yWMEacHnZ1gScLf6dbAQgJMkDFojZ+37Rdtymbo3F+QtfdxWRwvQg95NikfNF
e3YV2yKCsPFQxLFUTVbqaEpuKdpuvpx3IQtGTLhXcNyfhnNnEyHFzgkr3EMpbLEB
oIIuoD7fd045pXUVQN7LX2I1kDUA6doNiHOR7hU3awZDgNlPXUBguCuJ1q8m961A
MDubsyAL6mpbjbevKkSUxF/QKGKZlFscwmij68GkLYvCd+mjL3d2F/EpgAZo/e+b
8NjqJX/csfZj8zGr6QVSGjb5g8GhxRO42AiVrfU0nsBIP2bNVAw2FibsyM/xXXYO
4iIV3fm3LBD+jrj86m6WQGvp85F1xEPtJrI/yEG3MtFyrpwXjhTqIGTPhpO/pux4
HMuLwo6PN8XzAjjhCZSFgRF+8z5PDzRKJgp0o7rGkM2/tnE2FWj4dngkxIJXCoYe
+tCjsocKu2RZKiH0N4qw/uGvIp24ARbn38BAoiISRQWd8LqJIc6otR2UMvnzb422
UFwkT8lIbGjAgcmkQfl0Q9iB09NeYn349sH45IWyf7amH5mniQRcpjqDA461H4rq
NeGv3v9qX/EiCKXmbsSJKmVf2/ZBgfsgM7t4JNbdgaQBIj65KZTsGBQUDU7z2UCp
xdG+KMS0sBAy4SzM4O+PrpaASZUy1jciwJ1iGhe0kHqYILot+9NNF83oACfnUTjG
zZE9Q8juFsWjjq1UcMe4QwecXadWoMq7sVopw4eDH66b5kTJlNRQbi3NnrF9hUZx
cQvpS8L2LoJvoy40/1CJ9gAlckGPciIv8wAv7g4NO/35H5Iey3IsnG7GQT/cyWvS
yC20ysdXtOx8wvZCF8ZMn3n+AtfOJ9wBWtEa69o+Mi4w6kBZzt3emvrjwLewKcbY
hnMINm0Si701Na4zckes6D7cN+7QtmmHd6FSRe4WCszr5Wm/wOe48VQN0sxH5Lth
T2BKZr0UpV9tzxCHBEGNsvB60TtpX6YREJlCU56joqLxaKDouM1Bb//wccFmxFj0
bi4JbiDJ8H/Bqqx+6OshS8/pWT/WY+/zPpUG46gS60I0zCoLopuJNiAWBvYwvEhr
zJgiaMXbpHKdV7nt+nrY1HCZzgo7hj9/FrjyqUuyC8xZ4poJkWKbzq+yLa/aFQtN
5dLZnUEnpL6dAmtwO7sM8FZvJHkACCWUBXPpOl0Iss2uDx4qdw1CW+uUG2zp5At4
FKlpJ3H5hx9uw9ujLrAXK2c569W13OJe3wYRBa9wkj7NDxM58the2jGxsoVWRFpp
2NOdMtIdLcwTbLopHl9u9K+w+PYTcofQO3hyhMQ/RPUE13CeAb3dD0YxAC4fOJ6C
TjM2Y4QPm6uNUFT+9HcZ4H30B8kM4iIhrGXULHKYegiUFa0kw4owOeTvFwuNpWRW
xB5GwE8/HaU5C6Jw0PgZTb6FzoCZHVaUg1ryo9Zx2mMKfaGyGuB2DjWkqV5QYwLl
ddUqDeIxRXSHAiLBNcmmE7QhKmDqvyqRuVaeYGGPJqZnlI0N+SDFkQIoZD7InBUz
wwqXgS+ET+W5QIX9h+/UBAi4LTzff/ICYFiD/Byadu8v31BSUKqaI6CylIYMkUZ1
4tagtkfSPmftAjDPtphSRTL6puhBl3pGhIBSf05oFZeCPXFghuel5F0cmlvzZoya
XRR0FLZsy76Ai0Iuy9tpBvxuU44a+e43y64XcAkxhbBd7vPQQjDfhMMUj/eh7f7A
e6waIGyEOJgDTv0/oBhw8vG8e0vpk2Dj2bK+8F0HuwxgaIQ2FqLwgbnUKIE1why+
143+fDm6nxOh70SzY2aNtQa/949RLSS0AQCI+2w/oSo74/PfRyiaGbV2vrL0G4yz
t6PIDVBhwOkKLujGQQLgOT/ebZ+wCOAo3gJdKSNUgZzS0C2+P9LaDa22x/11Jsn2
s7PvudmnfSz+y0a4oFgNNtG8vR6L24EQ0Szt3OicYp8KRURYr9Iv50NbRM6XLSxO
4gT3kOtag5mZkYcMG+D5JFHYn+pGNfmhOzGe8cRZoGepeV37I2tknox+l/JHfLyQ
rAUjsP/brD6qMeeA+1iZNDfb+4PaPwEGUxQV0ORU/r2Q2FJ+L4uOfq562TS7TPf0
47hswUHtjAWM0bnNjm8sab71J8yy8xwe4oamhiO8W/jzW6GE6KTp+6gPjpICNJ7F
sI8/X8jzM/IsdRyYJMetJ1k0RB8Jp0Frs1QIbnCim3V7Q1LL9PrmWei27EmiQqRv
StI5ZAUpOaWZJxmLxhvvpmXzs2phTH/WOt4ZcYAyxpcgDL1JMiDDXemv4AC9kXIe
o1JTPe5fNusCQ534F8r45RbTgwvWMFPQISILJAUt9ZemHjE3Hcs7XkILEgnCrceE
CNO9b1SgpvNgN9ps7QUMoRoxOU6EbHRXbssiRnUtOtA5qK/TjW6HeuIu07bMsFpK
9Ceyp/8ytdoKlnI60DXXlDdD5QusT62haajZ/mm3q5BKQr6JEw0IfUC0qnZUplox
2d4JRNI94Ot8Q8n1dgyjoMFBZRO3GzXdk/Arx/OPQY8MSeVspes5CzMUThxnTh/C
/fgU3XGx0H3kKRbLpBm6yW3hmzOLQFeScbRhj+oe8xvUjL4adqgfQ27VoVvY7Imp
OXrpehF+1zR4WtgeYlMmswq6BVy19PZ88iUW6QKMrNlEic5sDrsGBGMz0Bp+3RT3
LJ8VpwMjB8Yzh/PFSHCvOy3f5rvqOaC+YCKUueX0qdLje5D0G9Co4C3+VyBFQoJ2
RvRz6X7/RsjmzCW/AQquH9YuArK7qsg0WMfskqv4gG/+3uq7n+UA46z3LIY4W3XJ
Pv/bStEVI1MK9fk01BGzxGmfxZxtuZW7sN0FrwDJqISqMlL+wXcJKhxtKjgBb9Go
KKx4/VZT496Y/Ft5H6si0Kz9AQiAYGIVvQqwdtXWW2UlLVs2w9mATn8UMNFYFZ4Z
UySecOQc5HGhaBiXnaScy+4SLEC9fztm0GT1bSGT8btqt8n4ucw6Cm4PsabF7m/m
gdX33/SNds+XgJjMGAJNVAGKxlBxoGJr0wwFiDWXLJKRktw29426CodtXj6DhB/t
oEjipv9n1ryz9UTZGTyPtMp+DKc5irXZWCrOI2JK3I/yF4dpU9osfXM+ww22HcWB
zzLVTlxWJY1rFkhPLezUNMgM80YUm7JKJubEdJD5tXebl8zNYp2X9oGViLf+hQr8
h/yeWpsI0cRNz1ak6bck0RLNRliGiqlN6MxiJTCNy5QOmiTaKlDbzdWRSE82bj5d
ZKOV4SvijzUJv8xRbCXhsi3MWTa7KIyT55dPFhP3+wqG1yx4miDpHFcYSPRnoS1s
sSLAt9kt3s1WTmcj158SVO/6TkQR9CBr6+j3zJ54VBaL7qoFWxCPekQpKUNUf738
Nn1dhZucdm8KyCgXhKdvpE0J+XxaoMkSixorLhfi/hKr5mXFkM+vwavnOBvQfo3t
ORZDRTY0oPJ3sEnJp5bQmIOhSa5ZS0Pwr2LFfDqeocj/RJ9Q+xDjPUSnccM92m35
Q38iUD9OGpJodEpc/4yYh/I+KlVCehL0r+wP3ZK29HhXgBwj4c0598Pdy1bAaMoN
9HAmkPKQgxdqIxSUaHGcuD+vgmJBjb7f7tSNwlcLgKyXXydHnEB5SfC2PyiICSuM
ZpvGrlK9GO0MVqyfJM1y9KqIUzmFAxn1M1TN2fj8D70iXoP1aExqWKPwV3xvdK4O
6SEnJiAK5GVGjvdpt3kxnOUd/GxiPZZw5/cFAmZ3qZNM1rKzTzTEMWJDEMWLQF9J
mSfW2QV/mpVpE+fUbOSJvs9Pu80aN/lKindkiy34vRMrw7i1osgto1nXxbLcR9Pf
xBjMkWFo1UktJJlgUocbQMkldh0thgMYvW5SN2M57+VWLO8+K7H7A4IDkeGJwWLZ
8joTt6wdkHtl2CBG/t9qSJplgGogO4pZyYlApQT0O92SLx7+Ap6gVLgc3bHQPJ6k
3q8ZTOnMBt1rzJRLiWTsI8dw33pTdVfCTfjcFB5gYuLdw3EXvtGUdJbZnILvvAcL
OR0Y58ybgBJA66MzVTdfDuffgXG7RxwIKByOwh3CaSysM5821O+5NozoiZX2w7ng
NQHY7HjRkZ6HNL4PLPvoX/AzpIWxD+Wy7+1344YfEVMZw11vz4o/UxidyI48nolq
8AEirJeY8Jk2DQoU23cF2/Ty+MGxJUNUsk4tlMikcTSZXMyu3/KQE5Q/7XewBv+f
3QB5xAJuHYjTsBT+Udt7W95nV5S8GF+nzscy452+Hb+RQd+UcKwExBX1/wE2iXU8
+L3j9PpkEw+9gEg/BTDNLwRoXIGVRSYtp1ryGA1ma7okqouYQWH7hj60h5qN8eRo
NQy3w79vfl1dr8Sag5rxksf4Th3kWqFviXmGngqqHRu2FdE+3K1kByZQ4uXoy+BS
4HWw/YZV9OFbA0gMQOQsOxdiVCrhg0RBH4uYsT1GCpIPn/9YI8LlfCuQNz9iiv25
+TGexM+zyFEWA0way71rLgKgGZlOKFyw3AoQqVS+pIoECy3yS0GLqNELb7dnUb0D
IPfBz4QSCcfe3V/4PFxDQVSIMrcCPsut5H5+2nOcSx+41oKGJB1fy3FzcDStSo/R
ziOPZrFPc7HoZHhL/bSUdcqSWgNRCehF5ryWrGRyapJ7FZ90e9lFLOkZGzxYLow1
Y0oXYhQLS4scYJWVJJ+WR58FcpsY+11MNObhAxa7GwMVpbH8zQyYSH0lh2ikfmDD
xiaQTryFjU0Ug8rXSUIDV8Nvvv99W6j5Dzpu0D9E97Cq32qsWKNeKIlOzpJsZBRK
z5aMelL5PJRGhx0Nibbs58sVCledb98NrWueY40Vh4oo11o12LnFkM0cpGMwhH28
+HlmvI/gvQMmRtjfsivgd5ryfpJwhNSK8AD7zccd86rnl7kt2kpiFtbXrx40MV/+
Gr1zKF9iS4Xews3srQq1Y5mbAlGzNLH3FNbMugZfMxZ1wpdUlBDAGsFey57OXJ3F
1CJNX4StG7VIGJscFlIapkw9gNXWvwdsZx/SxiZnhf6s6BIlUnl343P2tg2EV3jU
+NXLlEMXLoBRDm0PftV+hQyq3yzVcUIKjEsnqFNzC6OvzGUTxeFOwXUWwH15/hbm
X6e3OLvHbL/eDuTXNox2RSe36+YvRMeEAgLZDu6wfsIMJgHHs9EZW1QO4hZ2QvRr
scOmMyBwlJULSaxxmpLLpW4wV6PAfXf7uUDocE9Idu+DmUvRJFUIH0GTBaQOrLdu
77+FDt1hzQl1XmuajEAZ749C0GByaGbr1NhTppz2V143GS0G60Yr03Fgf2ynx4iY
xrEpcoH2kuz+XGlVaRF3shZSPGT4vsIzUFDNz9+bDindm3bwzM236JIyVocpHJjC
4WiZA8lDtUhDwxJqKL7ylIodVJQ+tqPRczV3W/xbYI3XNn1qsno8VtOgZ09FRFPb
DLpxpdgkd+yr/qs6dpp9LqR1iObYns9ANUA6Ep2Njy95FUV2ZK69Ge+wW5rzqDxH
OUCo6+aus+H/UVv8H4SZJ719LosXuLNA9wjb0kntgB6DyZMevMjwG/21B15OYaP2
8rio7ZiQj9u6DokMTsGob8dIJngGv56Idh0/BmEUwHP2sfirFPirJmClTYEVvIQp
fsBvTuwOZFiZtkZYuSp3rI2dcT3cCnzqUsBmdHHnAf+Ec/yogQa+lfEjQLoV8TOf
bYX4IB0jJmaLA5JXCFfo5EvcshpZoV9z97pLWSaT+ZMQLlOuZrJah5U2deRw4zL3
vJd/UPMAZNyhn04QgWmpnfvNIuV7eiaCPzcIudX8lO/PIEXH6GTHntP7Gdl3DA8t
tfBLHp7Koio4TqmmOq+HHKFaqci8OKuqPSbUTEQIKKGD1XsiWVeJA3QvHubON4Iv
Tyk2XEIz2RZxbgQYUsbbxuRihHw6ZhA/TEWMCoM/fTRQEhBYq+IPrkap9CRxWyaP
t1kbg+HZ5idmOAbOTu9ghV3upFS6VUjrqIN/nX2VfS4dfJuIscwDR/vyA7W4f1PR
6tc5y4na5ss2FCXUKzrzzFWNeumltecj1UGdDAcVhilNuLUW992y3gu+hiG3Ty7F
0AKTviSOmJ2ZsFQYzqtlsFoewi4VyduT4PSVTxMBdH8j93A1UKw+/hjo8YK9q7wJ
C9jAJEzheDmWwM+9RqQUDBtRy5nMB8FvWqPzF2lM2vVBSsIeV8ao9p704+L14+AE
E7EAzfK6nD4lL4ReCl6cHwAgBHvuY4/GWXSJDWf9QAczChSx5AA9f9X1s3Bfdxhy
py71H9HYhnHVhX/dMrlUnhWqJnVZbp82PhmXueJPtpWNiY1LY+dcM0djFhVix36C
GV3aPYJ1JGHyWTXmbFIO89bW7I+t8gcd5Yx86+GHtgrurgJexO1uWR+FSeERS+4/
S7hO4PaugpwyoJ5UJkioASvMPq6En8yBJH3xjAaXzBQPCuPMEJyK0qi+ogdDorTo
N8G+7yixAt4meNU/3C4PXNdM4vy2CgT65zgb+eLpE7ihj8TWvu2TUIEIGPCh2Obh
bTGIzwAodxmIMRq5CHg2xz9B5Jnyka25y7LzL9dmQ76AT/4NXI08bygCygQIK+d/
f5T9t+IIzq2jlyxjREMc/IVY4vJMeZadPCihnGBQKxh29bCJS/olQdEW3C7xO1Az
ACScDlB2NSAKALZewKcLSCykR7OEP69LVL7m1JcKL4KfWMrx+GSMmF1Ko2XLmoYP
czz+7LU1dnt9SljvR6O1RGruf5H4KfB+XMxOfIzudInD3g4xf6AMbxx0GZN3jnur
LAoQbIKsSDMNDbcxzz1B7W9mKsuvjLZeR4PWn9C1YoFrqU1jj4m8wR8jh4+sBnUD
HHRIRPTtGYZ+YQ8JCVThnsP93F/UUOc74eXX476p2if7Gh5IAUgxZe8RznZWKStW
c/sFt9csNCN85ZrrrvW+6N2MYpXmD9pEhGsZ9fn+VlptgNbh+hU4V6jqtjiTaKhA
9Um9sghEgrU0M3ItXw5eYDzTpaOxukOxphwHinK0A1zOzGNjVlmUtRAQhVPCMvJF
NPiq9I2kVeINQ26CVYwqgmv94bCYlZV9JhxNkq01O8ja6Intk8imMphELqZXWeD4
`pragma protect end_protected
