// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b47DAyJMQAERzQ8pPXvpoCnaEl2iWb2v0c/uD7+bR23M5y4jPNoNsV5vIgWG0+TK
6R2MDmlwUJ5JZX/9Nql8ZMInzJRK6Z0I+o6MaPdAkWGhv3gnhVkcOyuj8spcS1pr
5kHAo0QtcOpzgWoC4QETeSQafmnBIiPvRJld3UNq5eo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3312)
oSX1SLjr6sYzB/7niKKEFzoW9p+ba8YpR6CbmOjMmMxPazxNPfpVgGJ8QEqt9WCU
4prZV3aHGJOrMwQsWArwYSap+3rJ1cmZ6/h0nRjyIdPnnwwM6167hFz9Zn9xbqjK
nTcpDAzdi4rpLLTm559Px+S3r1/OjVipumoEfIEHeCktuYVvZnvmJZkydOmhCUp7
onxP8V/FHIVqVFIk3V3JkjefbjgFU/wvhxg1j79Lo61h9XDNGDTi3glxGa2oDMKY
LJeNLy+2Ot2ECXyAOlcxOVmCJFDNBbk4KwNYLbFOZ6RH58DSXQ2YRtOUiebP/q+M
icKz/MxjLrn/i1kwXXklzucPMLsGrI2YdjYMCqXS1ZUvEkqmYf4WKWq3jtk39gUc
KDdbly0uEQB9ZznTc3d0IiSCBjWRs7xeVe+k1NCLF5WqZcpwhmvTkqVWbo4wuPV0
sFxmeT+GRgm3vpxe6Tbn0pHqteBtgS6VFPFicAZ7YJliY1IYu2v8ojGkXA6v84ga
NipkfN9hOE/92Zj60wEeGRCqAj66jMXE2J3dY1gx/7EM34HsuqZOuEXM0Jr8MV2z
4/xEb604Z1ekyl4+UO4UyTgpaGWUBkYtrXSMSX/GhpMpyYoDe88kTp+aAEB4Z5lc
qvsXzzcB9bi42j+IhGqR67q1Spsnfnjn6GnsiERZHTGpOfFRSWn66pQrf8noOvrm
cFj4uInH5E6pLZrK6MC6SkeTqmnAMsmen0K5BolU8t5bH+s6UCP+W3ky5R9syCWX
mic5mVu/Eg9clXfqt7BP3UIwVZJv0qZ7nLjjeawXAOdXJ9zw+eUCHE6PcWUmnCN0
iYuFItl7B5SdESfnT8WiPLKxszVn6I58wf5au6qCOnc5VuZ1TIkh8gKXlBwQBrkO
s8p9tE7QVmkjN9I/kAVIGV9t8EO81wgumRjNwSdAynPUO2uN8mj4YI3ZAokzxber
HHQJ/wpoPFVCuCcpd0Zc2SLeR/7v1SmtdXXT2zJ1zzHtdyZGkhox0/L9IAGIZ20E
oTZaa51Qpab3kEzFiYNTPBdKYGEBDCYBtX8/oz3nneInnJN0asTS0OeFmjeNFmLm
xIjj4D+LpUxNKwyOBr/j75KagSpVqASw3x6lI4u6fom0tQgyxeKhzDzERgiDSkDh
NSnBkbF2/CfsMUg/FMdpsqeE/747/i/9y+7zCqFdigv2Xnq8qnqyJhi67niXPsnQ
EhVDgmRMZrggfNhgejHceDPUr3N6/KftxULOoqa0Gw60mQsaypTWq91Sgqprp55O
Yf+YB/H6IGka9iwodQDwxT9kVF6UseXpR3d3OagET63SZk0kZRqI9M2AyH5k5zJG
SugDpaCm74AnPDm/no7PRtlrQbgxNeBfkz2MKJ/vVSC5tuEUDph/O0fHDjfJH32s
Y8CdtCBxre2SEIg/HEBvXAvJCW5d+5Zw4tLK7cJR0eehFR3ApChX2VisJPk8H8o7
3hn12XYo/l0E6d/V+3wNHYDlNH5snAIvQJu+jnKa3FI4kUklIjQrhbdXAwRJtcrm
YiHf08ImScP7tWxKINEfkrXGaVOa0JF6ys+fT/tjEKphrVFiKfG4+7AGCrNFskFR
LPHoVVbqaIhjbHuybrzpD1hi4Da8MvOYyJca5FsJpsqSzDlWBCB3kiAd6fX1ciVw
duMuVV3qxHPHXDlk08aIvK/ldVgNWRB6XaWIsfr5YoSKsvvaToA0ZgzAytBhZoFH
zGxcg661dzlLeCgqqnDsjmwwv07IYMT5WvSApwG62Pbg17gipHm03tGVsnZWo23b
3lxBl8451C9T4kFiXTN37dLGntjmfcXwBM5RraV/odb6/C+dn+nFLUhhHqgj83Rd
XWTSrliU+xTNfATdg4yqcdyXw06GgUe5f9JVjFJweoqONL44NrYPPSh7W5h0X+iL
YLv8vfY8LIDhnKcrnW+PV4TirkNjUYV/AlWU67+zzJ04t+4TAcA2OfzxO/YV8aC4
9RJRQO60wthaJVYlRJJ0/0KVFp+VUAfn8R/7kRpstYFJTtH/qNwKb4PkDhA6TwPt
hc6Z+/6qbHWHbsTJXTimUxHbt1fkw47SsYXFeF+fyZ+ekjktCbjZw6AVz/EdY5ei
2UuPA/+k8V7wPq9unQSB3biq574TwUQMpRmo+q/lfFZbTV7Or6CkWkg8g/334YeY
U+YVUwjSoCphcXwCLALccLxP2O6EFhNmLdKqdHdViIAqlwKi+mI/MJ96cBofSM4G
HppfS7Z0BdNW4PjIQYiey9ESHfAmKjzZHKmJ4l5hjqcXVUqFO0XysQhQ5pXJNt61
hsbCTyrK7UHMWA7rzL9UgvrHkusy1uofzIlXpebOIiDjd++URJfFD4xd6r4gTtkj
Kk3ucgGCXwDyw0Mh4B5gyh8Iit1J/03STdBfxFv94gpyGXT39ivYw4RNAnl5Cxy7
sMvK4NRhFsC878lMLVckUbV7w4FGtv8+fDzlTto27yMpdYMzFPrTrYng9LWNtw+Q
ZPG8Ntl6PP+srKqWOtgxhHRPSdRbVGsqn5E7avngOUY9eSNYkk4FVl6SMyMzI2mO
XeBFkohtMp3OppdsiUtYfiksFAReNapgCkGAaH4ycTz8PS9y+zzW443MLRBuxe58
9qymBrYYTQj8x41zt1XzpU5czpzk3frJXspeunlCwNOKsqGjyrNHgUYNoieahqNu
FXpfuE3wTdovIQiHyEvSjgYOU2A0amqZ3H943fC/YIbr+do2bh4nMc3mQoXyz+x7
KDqPoZbl4KT/CCRFsouFqHlku2MCP5TSnlx8HUU06vvYBYUUYNdxwX3xO9nLyPQT
Uwnn1O0+8xKvm6zJ9Rz4qebaz2QuFnKIqWYrYk7YIXHva8fRq6L80Ukpw0Famw7B
+3cmQpQdnEv1mbCVcyuVLbFS6ZIl4x2w2KyN1ceJxYha4hNJcY+7KXm+E7wDCNPe
GL5i6qAxCkdfsoVVsweKy5imD2XZieuY64/RY+MrjgGT1FL3Ex/Hqwv9Q8g0p3jQ
TIMVGVGmujMLZ/VWhmMIlx5mWaf5rHCvImqcbRlvimiINiLkqLFn8kt4i0+9kS4j
RKxdkHhoPic6dR/6bHFlF1vlGS4rifKQrorkyKbCpFOeO3UegC4vO4NxKk3ahYPZ
xLFRCtkMc2U7xWYiQvlZb5tAENWF8cNvJJbsnUhf14RdITSe/u7mZgVTci48W2Zu
MSzL1tJEB/deWIfepTxmuYfYS596UlAful9Nn1ZVGS2ZNSKS5xAA70mgsyinQ3Ka
Fbxq43zZYVYBuQhzV0aC8yy+i2jEJpmtasx24ee8d+HSs7kM/xHPwMwWgFCxvIBN
mXZZQS9g3jVF65EOvxIPJFKwNUaog1+LMwF2sISF+ADAAfxNdgIaWTM4jcFZPrxC
0t31Q9Q2ZXjRgdCkQ4RFKxC3jj57oXqZcIaTpeKSTGKDqYcBPcv93DtCZDuQpXpa
Rq5TJl2gWsXM515qhAZx6ZumrJkvnqzcPIBdqeppPYAx+VE6rDBxiTV5etggWAmJ
3zop+R5/Eui0suiwsR2Z+BEFqkCf+weV0SV37o/wZ+6/PVKd/09EplAOmc4d0otg
D8s11zYJUon31dkqFQd6LXngiU35ci4yk4lEANGYO4tk+s7k7cMb/548gXihpZRM
2/mrasQblMGi9YnTq1GElJHXtokXfkBpRukkM54ORZ4jl3a6IV4h/8uy6breU13r
wg70kYjsw5r+pOAQzCETeP8KVpV/nuP+KD9Qdj9+9kB9S9qx3Ql5x9EgLfkBdcQc
ZQfel1mUk9NYnZpDT57EInqprrxmGyB+DJVpPP3Zyv74RDXJRKCIQp6E+npsloKJ
BjKuz1w7StNf+ApvssQdONjhGz4TIUaTnt/fyqBEfn01OMJTzTL09qKTNUj/qKc6
3gBCu1Q5jV9HAYCHN6VO5MPE+cAbb/e9Mk2IxgyPd0E0p2cfIEsSngYK2mTA7vVB
e9lQakxy8pBXRdrPpDEHsADf/5UB46tSQpa6DItz+u/tkTljJ8vMMX4HXAGnSJtV
e8ItU1Fw07yZ/iajb8yUJriWeIqh1V+YDN7kLmdYkZI9gnvvphnLHKIMQ9se9nJg
aMI8BGjtfPl+SbPYbDs2ubYFZRr3Rhq1nhh/jTqXgnY3cF2wBZyGCGTh9qzJyOOg
qWBdkmE6On5wNUz8fKJtN1Nkt6QHBk38Pc9tRZsaCF6zeJCC1C94/p023Y387y3+
vX4oOCcYfYHDopLwilq5h2PocU/rjgPWNUQQ6sFeH0+H57xxkSxDM7OTKc7J6hgH
dGIg3OdWX4zENxlr7CUTpoCtoarJ3mSXWqvoLqTP3STSXuK7se3yliobjLTvHcp0
nzhJrDo2atF9PDr6Wow0k0yanvX7L30DhRJZH/MJiOp/Sx321TAAnNnvP3oMoQW0
`pragma protect end_protected
