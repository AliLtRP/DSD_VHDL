// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Atbh4RLx4lOlOCBDAVvzyBPPjIOjkEq0w9yxmOOi6vGgmHiFr/OyG0v6OXDOuFgZ
riSPeS8MD0T3lRUiQmDhvfKX4xUYpkZyDWxLEwC0Ht0UwtyKzu/UWoYRWJcbZAwG
nIdYPvYbNBakSjihtbK5YWiBkVhVhe5aJOyEsxEptyw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 66432)
uwbbtpBj8kVMg/5t6y+BKautcS/GqeekxsQLcA1YHUQCKhzwD41FtANcVY4XbGkn
rxbrgPNzgoFweeLTyoaDNsdyztQnNNUs9uQvVeJeOIXWgFcwgFAp/LYpklNm+baA
mnL9Motorj7n/L55L8Kmr/ixXSImWelYwR5B/ufKdRfVXChxgx+3yITtUwxErFUS
9aq1vlLPmZKAQhMvpmxFObU5KI0sIypTr8U/4mRBaZ4IiHaU2NdYXN8lWHR9cfss
d3zm7NyofrzGz72u7RrJHWCcMa9WZyw1951C1pyTMAQt7n9XfGbqasExg1Y1kOx7
NkryOmv3pAz4qgGhGtI/tr1dYfGlqsmuFlrUgXU48F9RgJ0zMnJHDjEL24M84lP5
FCMOeJ4nxAnJCt4SVLHso7oDhZnCtKDwYjnxcgfR9uL81vz1AbfEnyIWzCQ6UJFo
r5MY2IvBDkqL1iWjPW6lASgXwojd0TBD2b7N3J47L7UdYwYCQRnHxOmvGXMCkPJG
2MLQUS7s4LuvFGe7Sd2iG8bVuPnszyJppiOaYBManSzeAuAdNsVAoKOnt/ZHKpoB
k0MdjspUtvC0Dw+rzFWFE324Gg1ffzhP+G4P/4K89kS5M1YfwCdJWsAjEmPAI7s3
dslz3e/+XfneJTknCvp+LmRZiclnF0HqjXEBNRiEKuxazgJ7SmGPM/2t7hERPh8X
fuHqrhIMkM2t43Y5unIrgg1nDlvq3VhV1BpM05KYXy2zF0NBOtlGfwaPzxpXfj27
XRhYQGVym+VvGHaJOo2zK53VjIKrlMYRzC/JO2+7Sjf2xLixfD2Be+LDgzqiTHIo
guM02hMyGsQsgV3ofPNB+jO/MOYMdXFq2PGegQqqVPj6g5zkDuHBWvj2cFvDaFCt
6FsOLIboCHOScpq5Upw3HtoBk7zy72Kt3j3eYukGZQORIwTqGZK5mf2Yshmqb73J
Of5leT+pbqnpW1BgXyvPY56yEykRjV6IRA3vFQYL6ftt3ZBmI/Olv1tBAi13EI6S
y6YoD2evdwEfwDSX8ZCeLbXLLaKn63fgsDAU+lgJanRUrojN+slfPSWAkOjLkNUv
8PdiLNLXE00QNBrSijYcNDR9pcxjCrX7aiLZmR9HbFDhRXBIxCnfjmjsTfPP2bqB
riASdE/XSn/uTeAut6ccNFnO5DgfgOFr3m2TA1U24j3EqbYn4eTvyA72h0zo4kdi
8jc/F6lIjmaO8lxD8Wl7YQtA2WCQLofOXLSS/1jwYZBDQB3uDiD5rNPuFnF9kWLS
/S+HCFd3YiSrIKgs9yU2/qgUzLfWGLXFMdcEW6bEWQ9EKAFRAkH2qEQlBSy0gB9k
m5N8oqPvssH1O7L80ha3nTn+N7vGDbCdNfvj6hFvo8aiUAY6wkZD75zRhpXPcoiG
lIrt3y+E7MZAO0Oqj8ZU294ZRFF0ESwwf+F4ifHwKoMT5DFCRlexmboGzlrKvk1T
iga10tkkAvsDnc7kp6gAbZM5VYe5OVHPzD2X2Bvi/9FonZSGOntaYGc7SwgXQtHW
ilGAHqbDB59EbUMwv9+k7xA/0vdrpfJ1U/c1WWIjJGxiggszUtHm/N2uN4qOpW1g
flcymV2DTFrJ6rNenOaGCtMsrAQ8CkqmVpbVe3czAYFrvAbDF52W4p8PWGDQ9hCi
iakoOngF69bzv9aTCIhKZJGCnRxu45t4Ca5q20EukHmdGjMPCBpzBCh5eDVqsJPK
OZ+JkK5sCGHeXwla9geit37WJQAaC6GQpbsJ3OAQSsu4H5rzj02tJF+BR0Hozsmm
3JCG6he8kvEHr1wnlI4Xhyt0Byf8qKPAhtjgESykaxor17NOgowwovZ0qed1vSmA
/xEcdS/FpB+qyT5RtEbgwNPPjvQAjRS1uDwW6Az5Rs7LT0Ea0xAhaqXgReM4iPb+
51R/iJCfCJe5LfY7acyB+dw1FJVol3V98eL+YtqY2cenVpQC8a2Q0P/t98sKud6h
1Jl6N/2og7MDAOp8eQ88KhlOqNb+UgaIbG3KhP5P1qhkXC040njJH1cou7vN5sSX
VWYza6oP/1S5wGV5+0M/C4oTyCTm45YvOlevRG1PqEYxKby1HRTKNdQ/Dwn1a5nt
5ZWvahCo3vbdKVtRoIyAptR8XK/RhzWDYLPVjQVeRwIUhjKPoMtY1/9HqntSZeh7
EWPvimaB63aHa3dRhDsJfStoUqNlE3Q8m4XP6uXDld7XuU8idv0eY+RStbaQETWA
4tdse0C1ER05Kbg+IYayw0H0GZr3U5GbiQs2EylKEb5jC+a8WD92H1toDk1sHMov
CzT+/TM9QAyaSYOYwm67qs3LsxbDjoma+HtWzg9lZPWHkBoYowiLnRko4vxgZ8Ow
WhJlhGGBd0iEnQRrmCNUbMO4ErAhajFWxc3PflXP33NcO4OXuzMQ3vtJcmVJh4NN
w+QcNlsOlokJ9OZ9lVYNypzLyMBfcYBIG81h2mJakkoZI7Ee/Sc89LJaV8gL9hT3
fFkSdee48gYjljNBSPEW/tvV8dqLEy+2sJbop956kuBVahyu8Nfw3//0Dik2Z88A
QNR5y66w8jeIMB9z3jwxCu22cEzBMGHk2htXKQBjKWLA9Uw7tsTZWjtE2K4jeOnG
d32sc0HNXOYkjTcHbdQPSJWwOw75dog3G+11Ql2m3482srMlg/hqRp7tCUZHvtHO
0yOLjjRjpMt11I0XrZt2LEbUv59a3K+H5JBQedFphQq9bUz+WD/6XIyBfUf8AmSj
xv4Y+xBKOKnDtl9yHuJu0bFHmp+ZGaCzt0+ZZYteQDcu1RdXzYbZRkCirxLWQ3aX
oXItxsUJlujnnpdqIwdHFW2Gov90axxrWibtozkS8lLf+FUfBubgZNJEo50jIWm3
/UXig1UAxelJiPPhZ9zU8euiJaGOecDRU/k7RmZJl4fbTLEW5z8y7175lUSUXCpT
EGrt02j1DE+VtBDoMkVfaKz6OAMa5gBCOw48icjHrDInz7YL+3D9gAIbim0nMU5J
9JiyKed+eGlJVogN1BXSr8OmDYVh89/87TWEbXmIJmzauojU98KrjCHq9Lv3DxbB
s9MNJE1i7FMzDzNV7JHyBeqfamqKPeBmaUB2jYH0IfPjfJBqniTp3bz917UzxTmr
O9RDRENmxqI8rB5W3I0+xOGTrbk1jfwxxKOVcClZ0gIYggj3RsNFmGe1V0rKTCzX
jGEzub4amta+sILellbTIhIBrsjos6Bydv/4MD3g4y3g6X2YtPiYOM2wZKBEG12S
pxDa2Z1jZf9KxZ40HfoHp8jjPBrpoWy9wttczzFSf2+ad+/SNxH1tgH68lT2nx7A
ZLEF5fsS+F+jsGefNfYNs8f0G/4QqdPTvREj6glhXvgN+omoBVHgYbTsibPAz+BJ
z8zxP3Ir2x+fa86vtBG8ft24YmiaJy0btA5IotSTP8GAn+D6ELUvKdKfJ3THx69q
p8cmfV1+TTg63sKUIHMy5WsifL9gr81guv/R2fplRNgqkY4L40SiSQ/nuDno1YGk
UTMo49JX5QhYivqXq/VvwWe7B4kD5IzAvmKZyWf+QZTbaSswst/SDH13kJ3RU2fv
sXY1RjChbZ6VDEVKkRJeadenb3gQje3/0ryFp3I5+Z69x1Drd7ZG2ofNYyQABFab
NV/EqpelIm44n+3+2zveSVgSLgF3BYDvZt0ubencJYnUy1I5aI9oRmdnKfvUeZiu
PfFmlyxCWjUHLNoTSzvfUEfRxwLFBOJYzYOghmVP4+B33QdNvgvArmOvD3ov4GnO
cK923DdM5ivv8MqbsMzG5N0EOgHHJCtu4QlTYgLc8y6oA+dr28GuGBPsH42Xjkf4
q0M+WJAhyFjTMj9Dzd73RRlOVi1VzGZVz1wiF3aX7RahrZR0wh3/s4lBbZZeRZ5F
7+DadGcNKfIh4+D/+xe5XV9ZZcnIEHKnzTvv6DgSrI/7h1MjXe2wefgvwy8xv+3P
xkzpDCLEsJvQ8cfw2jKvpKavlCkzUFi8TR/4ucPcwjjH1/lw1C2JQISlGgZcyCKl
1diOmYzQTRZg8Oyjwg2WYG2WCzbvAZ3cHsFmrqAyNjT4kagtZPiO+S2o/W/8zw57
t+v/DGLhqZjnVHD/qksOk08UnekZNiwPTGAOVH0RPaexSFIza94LIioIiimc++yR
JtA/GEvdKMilv7yhqBqIYHBpbfmtqCwH5g5rtIIf7bGwYzd2rw4+HnThr99TCxKj
FkH4hm4vo0pOrfxRf0NJed0w6L6397MNRfgozqB+6IMCiDxDqUdSqR7oJDEcfknc
/wbljJmTHDYoa/myQc+/ZgToa4IgPFqj9mqGiMTOHuJ+jk+2o4zeIKLKHdSPC4WJ
ozhz1DZqKQOktj+si1vOU4rr5PgYLvrqJfNSq6EqQ6rt8hG7tzkw/49mizKsX0Pq
VGn5pqdeUsaL8dIX5XH+JieMz9R88HhEOK08aNObb8Lhw606VKtXDisvVuDbuN1K
skxiZnMqZeICs3o/zalTc4oRT5hm7wn8aURATUEJ+KwWSdsTTbcdQmKKLt3IzdLI
am1zbLuKxvkoZn0cF2UAqh9gIhThhMeLPxxPC9LbM4rt2GqqqIixU+J5e6eHqKxb
r4ls5sQZM5j7/a3HaAgWfKJc/jmqRlzrp/saknaNyYicYgaLpXi67OzrH5c1fV57
l6a14NKHUMlWMe9/BfCHVY5UzG46vMnFZVHmlhHHg6z4CH4Fhf1MX9WwMwYfHSbR
7Ohm6Ar06Zbgx54KjgYahgM115uMIo89McLu70GrL0HVAMse1VAitIoagzbWg2l9
Cae50/ALtT+uSDQyNNV8pIFIocKaGoijgPc45sh+jzqcrN3Tm8tZPbP8j48flRUw
6zKd5tb9ADrd/4f72msGO9wNSYJ54juVM+fkC4+KHs4V7iuKQCGgQnGVS2D0IMCB
c3x7TwLgNObfgWoKtZLXCDCxCETN+q+8/TdZrdwkZn1dT+iYCuLsSpeSbQM9WZi8
s/+0u0kCjCiGAz2TbrNn9Kpvn4k8bw5qU3us/RWH8eE5YC7yGLOBEMPnzR1AbvYF
B7AdIV64+We5TOTgNesC8P1Edcqo4qTet+ECEBX1AwCCwPNW34Xdv/zB3AHBmX8L
KZz7oaUx/IYHjH1AoYJXpnl1+q1v6x/z/jClMs6m84EdA49u0PSA77UfVL+7zOjJ
aqV0XrMuhGm8dbPCKsSmo8sz6D20Tmb+XSL04H+sSqCBlcmJ2FdOCkQsJRn/Mqpu
eOLWiLJJoSxhJnl2kJmCQgp48HtYAj4leDmyOlYQ5tVerqRRv3Vj6gK6jv08VpGU
/MQ/YQuLSQSpcXRvERqzVw92WpiyK3hwVq5cgyJbZ4jrwmDVF4PQRQhZKogh01Mu
H3Fmd+XO2zQLkEi2TGXx/fqv2WeHiG5qTwfezLLx2scbJnVEAmiy7KYfdElKIWW/
stEC1feyOPtdu8hNNr2RcBwOOjcIMQfBOjl8jYthyaY1SOrojKm+MFzlEOV+s8Gi
Ik4Rnna8e1RVbB3/2PKby7IC1oa/RapR7ksi9c+Llb3D/iej1MiTiqjAY08BAjdJ
kVgk1k9W3qxEsIeMrloTU+5Ym2KQKc3dqIksx0q4NGeFd2tFQp5+7RlVTm7rlOFf
fTgxWqxAJ5P/sLgCZdGUyDcdGniKtcjAsRSYqBmLkzzYchQT4MmsZLjG2wD6nuwj
D0wvlGfXBMm4U9OoFFWNNJRNuE7iof2q2imn7NEzPR1PdkyuC3w/AV/TqCOohlrr
fqWgS+udXxMPBUE15mAgx1t8o/s3zkpAiR6St2ujpfY4KSBd/Vn9oNSpl6Wbl5s5
YJbT2NtjTxT/vkZm9sIndGBcdqMyMtVjC4XKefAr7Osn8RGxLRb8w9sccNB3oo42
AmBtmTCH0A6iskb6NhSp/r0twIHaUI8J9+tHw99ircq/ZqfMv/M12HQc+CIFkjFk
0ppKVeBfq0/k0S8Agw1Obt60lE6iQggAAt/mG4ZHxmExoUmnmkEKy8U7S+fTERnq
Mu6QmHXTjZRb9HR9Plxt9i0QWBrvIInkoY2I2trVZc+bcWokjis6//wCr6B2JB1r
1ADFmGYqISjI2wk44iGYb2tndZqN0zz2C7deOl7xeUBOY4oPD1FeET+FZq7Yyzkv
1Bb/eCeidae4Rq0I3LK9UbqrfNfwWmmz8kEPt5uSyik4pj3yvmg0+3mJ9EaIsKqM
Nw8DDNH3DYsZBelM7M+dxbCPG1oEtdcAA74zIuCT30TrmKy890bt+I6U9ztV/YcO
n67MjH5a/umgjxBOBTYElWGHmgkjYMtY6rWQBTy+02OD/LmBkeL2MIM0YfJ5Zurq
g7YyIr3ji9GWLO9UROQX1Sm+c5Wssg4u65WAGKAJgXWKzW0g9mNIo2MCF0ldkzkN
JwFzYJo3cizRHRGahmadZfhBtoKL3qIdLERexYO3DN3bB0Y2oI50mOhK+BZcd+QT
/Wy4YQL+qrOQcvdmVvyZDYnw1wjyyEUikpDL+1Coa47GL42BQhqExspzAxe1VPiM
fCGZV3cTwU9nw6MFdWu+oOmVKEsyy+gdnNDg5hbewuHbh9cccPQB90CBOQAxbD8g
g1h8PFsH3PCuRlq1L6hP1/p6K67Z2PQnAnfqsrhOJCsEU9DTfVZ69uCUBwwE2OYO
xLFZOvBqT/gPuueuQqsHkQiCTdB/AzUGZUJmSB9Xj9nxaxDx4p5Gx88xDjQO3QlE
OwC0q30UJ3B8vBbN4yqkdO+2DQYe7dIla3kKAwvTtrJ26nNfPpBEBItwuiGmNLCM
8Ua2NAIw2cEtXGRpooLDgWk/r6UD78NjQAM5/Y7fhtPng8+TPVZXr9NdnsMPxtJF
LRD4gFGpGPiqBD1kP/ZziziBBtRrO4dr2xOYKBOi8ld0NX7I7Jb4tjzyBpCDNvWD
/rHB57mPH1BZAyIzLiUcLBonvQD/DE74xQ5shod8AbgTpc3KoKCyWXT1YpWWMJtY
oEC3iFYj2XShnIuh/YoLEqnUniBxQv2qCbwWhRIszvfEuV7lWYvpS4637oT/ny4L
3nymgG9XGZQTzFMrbpS9IH81jo0LWPa46QlyeTwaCBvd4R+2ShncaCOgAtAVovSQ
8AUgYwf8vbZj+/XMDk3qXLgxfWyZwivmCvDdRZzeKS9QXqM3NxjFtXadTgmJz5I8
h/r/ogWHTRfoLLgBtLWD4XPZHg4wduZXDZYE6uF0ekypJ5RwRPaH1h0yq/aAWXP/
cfiy4hNZQ7Zm4R7ii40K7sVa5fOLPkbQuWeqaoOrrqOhGNx9GgfXRwqyi5HLNcVq
O2HTH/AQgwV0+YwFaA1gbJlHJZRDoi73UHK6RU3uV5Nz1WB1gWZu5m68OZBrxxH8
jgidfoYcvdPDFVrsLmncS1iEuKFJDPgKVaKXiFpXwZ0Li/1MfA2Bopz1v4eCu7jI
LnMeucRpj72rBbNJrLvQF/AmuuJWPLZ5j00q6xU+Fk09s3m7ahlq+H1CDB5g+2CX
o07F9JpkNuRDSzDt7m8jOUXGEx7XAm/clsallow55fTxk5ucrenxpuDg8OIEmlZ2
7/pcStKUYnWwJ5+XhXSn11bS4gdGEjTN/QiqRJIvyZM/5sNLoLRcZgfq6JehqTgL
WCZsZl+0HJuMmO19RaG5oLPHcSL5KXgsjKkU1R9HD0yl8fqGW+dGidtXj2kYJeAQ
Cd/QXT06Flk7f9mZ6NJE1lJ7p1uke2BgyKAA5mSsWN8j6hXBVSs9KRV+BmDCBLzx
h8z5FLPgn5+xLjpBno0wzp/WhwJtjLzTDtRTTQ/2wIEFjtNEU0dx0L0brPCgj9Es
Sb7Pg5Y0NKGRlKoLCiA8+KGyuyCMSRxvJ/zJ0h+arxP/SZjB8Hze6ZgNbVkBP6AX
Ov5ixSLfqoe1rc64Tl3EZmQHxYcaGnkiL+G2irMi0n/DezaUOO+CDW2hXBT0iGQm
dt7HrnOGSxhG86z7AfaFFX2QdGWNkkErbfgilzBeGU0oAQKkwuLYKAdtplnyJD1G
pfIDVokAnrhqmUA8qgza1mWHMaiR6C0BEhHCzPd5VyuCtl9B2YYRk9qEiQ1yMeB8
MwmIxirwkEraOLi4Jp9nvHH/MwYu/TdS9cywb3fAVRUw49WS5C4oECC1SMXn0Poa
6k6SP4dAcqT0VzgUZ5rybgEEqOo0qM0fT5PRBwUwyi3H1uSS3S8mpdrP+95/qXeQ
2fomJmucEiEfAWo1o4WuOU/leG4By0fIeftJ8IydP4kK56M4lpbrXnSFgsjVZHyc
h75Ii38ftk9tRE01YmBAqlgms87XqHmGbuekUtgyPcSytBwZ3wvuHOW2gMgfrQ0i
X1mPPLmHs0qLJwkxcKTpikjCguHohAQFwZjdBi4Hx7DmQa7HP6f9mCNec7W6oDcB
1cEeg0zwnfSfuChCvp+5D1qze91Ic4GtWFRGd803LQrAcQGE4SYt21g9EaQ3RxKG
Xha+RadLmcTk9O130Xsgs4knxIuOgXiAaQ22m7xhQMcuk+sGSxgRYDltSBMyJZis
2ZRIZ9TAMYZe0pQ936HKTHn8cX3AERT8lg+F97Gdr+QFCCe+bWsG8xsoGw7IWmSy
ZfDI/UoqIm8EV9MNu+JG5VKsNUEYPmkNNL2QIHVEwlHrbl0JM2VCZegjUyjgfjTE
zdt9wQkdJNWnoKmkRAYk70XdoBWmSTvhMwgZlbBcDeQ2T2TcLUhO5WA+LMvB7Yb3
Oqmd+xaUAX1k2/bzFoXkWK9+ttHNAeMvC2CHptYueXOQPsrAmOovGlWOfKIIa7+q
8badVB+ynsa76UHLrIalII5zeCgKzXlJsAd4YnXsXPohQLvL+BaaLK5kT6fdqU82
pxthKIPAN2E8yawRFZwe1aDF/lJQMRdaLiS5U+70fzn0Ou9b6dhM6d73MoTweJD8
RJIVkoSPOQuXUbGTiUEo83zA1zaUrobmLJ8TfOefQKmmDqFy+bsSraOHNDKkalvc
NzQjWKUa/1WneHHK3Kgr8IStC7B9Gpeu7UXOjPqc2WeKqxNhgxfZpRZI0+KYj8A1
oPhsjq98Y8kGSZDVQdpUL/HMuTGN7ScrUD/knIMxSZLoiioUJcN6B71OEfyiPxWI
9njZELDDW5j2dEihwxhbml+ZMuXxy1p/ukqYNbESN1cyMHTnYQzjWHBpYijerl0k
sM3BjFh5bA+xrwKGabmWQ+ahCg1iRQZLuUt9cQcE6NmCXtsDu42tmJ3qGUEIe90H
f1BpmlM3WtAQzXgzRE5W7Am0nUqsX39kPeAbKxW9VeqC5VgGMqenn61usgai5kGZ
lgmi/F70kY+ZUfy+a9xEpR82OcAABE4Fld3xkmJ4oIIRfQkEi32O9pWWtajc328L
nURKtuTiM9wDQMh7Jim0Uhb0KmyOI5Wr1GOMKvkgvoUC8hxBKOGGVvyMgg0lw0dv
4TJnFL8yJR3fP0Ej/tPPwjXbvcwr96iGSJrxIUB81jMlJsaTl3OOWJXqPd5pjxwq
nSSk8iNHRv6Z/mPmpCscFP2r9sVEgutrDDB4nu7FoRiWOc45dE1jD5X5GjBwIan1
YbpmjRW9WC/6rdlKE8QefLPvKAFnptckZXhfH9/3W+u160Ccg6MBjUHRQpSB7cRq
x+2NaEzIA11OBa54tLK3iI7rIBEz/L17Ou7JwhKb/oC0+wyCvtFhD1GUiIYB9bpf
87inPkysNMHi8K5RJkqFoyEt3pZrCnE+xSLtVgV2W603UGxuvSCFIlRBUtxUs685
bWAgXZoM4yUmoJ57kM2NsGM1jbeeQZpTrt1Rn3seVbZ/cYJ4OJUfohoAPxylsSWb
1Xi9cuwA6FoZZZekYYg6E+10UsVOL/DBnDxILYNLIG4B29HUd9h89zEm7x1o0xr+
CT8j9HI+0j1eHMeTMS7PZI0nimO44JXBj9+COGZz5eRax3OHB63r5IPj/p1kMAQ7
OOmQPa0kOvclGP4How8sJdqXNrDy7IxCXurrScp/p34CMu4NJeAttQbGHmaJIsrV
ua4O620Sdsnk9BeMS5ScYMIxmq2rTn0AIcXCcu6GZceNcyL33iCAZsaD7SHOgxbg
580w89wyNNcF8evoNWVPnGutUrI3VkxSAMBU6MHUD+C5zMagDai69qWZyPVJfArw
03HbhriIXBPrVKNYi7gN90anDLTdzqJiMo5iqOzNR3ZEGknGqUGeVPe9QDzKNmgy
s7R1ANEvHdhKdurwlFDkUtXXTdVrLp2kT5HHhBt4WKjiRxCRY9JQqczHpR2vIHIi
ry0epFE7yoU7sIzeafNQiekknuHusiJvO67wBzQycBSagMD4M7AfYM99GVZiIjZA
QvWswgRn5yV0IWlD9qrPJmoALhuhggJ91xOGhzieEoWPXG41REqTpMCeLUpLt1fR
hgzm+aoLZVvfhVLeZG8HGPi+laaS76izeZAoJ+/Wjzsf5EAmz9PKc1cmdnYK7YgL
30/ITwUh9ZWUjtJ17LlU6vd7j2suCIK0PF/hA8dHfdViUNstZjgB0HB+uZD9a6dP
GZYpfsT4A69wGA/DUrBpys6cSHtoy3HtfgDwx/uiM9FoNiDKJmS/rtIuHJAj4MwD
vtpibvRmlGvrCHgzst5LQfPo5HaVenCQ5BA7pRJENr9bqYcmm1Et3/lmduGEQ6Wt
dxSabwnyD+7wvwWSoCm2Ano8eQnXtmUq1WM9X43epOkyrO4bs15zw4z77D/+V0a2
MZtVoa99/XpuxjaIWVUYMiS1aX8GpzUISCAeBWt5sJijO+ZsLzll8wgsHJfLk9cm
J1ckdR9miPl5tuR5W1qI0+CGz4YYlvnC1v0FgW0RjZZG/JyakjaaLI3H0zqHVTNX
xGft0CMEM0SK6pOC1CF+hP2eKPsMgd33vqo4qC7Ok2H2cyQzNjO7Noxi2gu2YmV3
p6TEg1GsY/i9jBwOctVstT7o2NzUSSo/U7gNVtYafrUIB5io89pq6gBf30iS6u7K
qUBKLHPKColy5NMTrtWiUeuvBwrDblyzbo3ydepI3y/b1tGOWRBM9FkJ/8bg9M3q
0SS4CAqvpm62NiUSotkiOhaxsXSxI3gT6o/4Ihx1K//P073s38U4Hf+AvFVVO5ug
q7YkfV++dTHSDjoJkqhtWXzTXfMOZCehPS/vOI12fNr4a/JmukGgVL9VWbEPC9v6
cFFcNue5aGIkwQUNCxxqGVXa31T16SzbMckzDce3+aZPstheJ8sww04qchlEolBy
tYaQS09EhYVO6gf6TbZF1K41csarJoU+31F6aZWdxnAuuEVlynPh1UczSRYXWzmT
dfxMohlRUSHcrix9XK5DXmy/UHpcN/qZ3FELDD7SPPj5bSopFBe29dmgpQm2b5+S
5ZGznnFGtMi7BGuOHmN1TD64UCAFvKb+E3nyb4ijLYi6lgg7f6B3G8ns+eMcceF9
U3Zin7HRHxt964ifF6iEi/0YgYmu0GNMSiFUXnSQrbZxWXz66Lcz+2QawaZTv37e
GjmCDeVlfslKNZMRSsjTJKuX2BjJObxaq8nnVqf5VIpsRhbkEygMjJaLYUQyewKu
ijKcouUDgBEKeU1LLyDHQAe0LbM8bH5W3PG8Wn/5hluiMs6VdMVH+GZ1eaUuohNZ
kK4ovnkeApLMd1ycFqwb3OOlJ5Cojo8KL3emN7UOYEyY/IDYWTkqoVrVWJgykMXi
Mv+FQHj6EAGJ08YWICpWjUPhpgCMpnfWFV8Pyr59q+Tf9vzoMygSkmAVFYx1i3fI
Swo20/W2B16LdRbM3qYE8Sc0SbuMFELXU5GTi+NUX1vJTN4el74jKp77KbqbKWkJ
78/8BgA6KcxvFMKJtu7QFldcbsLa+kMls466RAK9opepeZFD9hLjQwUccV9wuLCN
PMtYhmn0qaTV3wOtnZvkFnTffNwnhJ+fgLwgA7kSgpo2pvlQ2jVDn9xjWHm6GUvT
7bCrZzaKQMfy+64jxPviyrgNAVyEH91WJlPDGVgwRYMUzZVdl8gza4fLIVfMC9fN
Lh/5Wc2+oDNB0nUP3ivwVmezErJpw4oXEiuo8OAGPsSTz5M+ml4a6MW9+khn2u9F
pg5jd0/YFNKVejbmR6HOSfG3Fwdhhjc2dCENrEFsgDSeriDzF5hRljf8tz17EyFD
wIrhsRygFqTgZYIqVAcOB6xO3C8h/9i9UrQKhaeCpJhunv6AZaVSJcHdw/3Pq44r
PoPO/JMyuAZvuYDZ3UkmbxVau1qkiwlzml3F9G3iIsiz8BLY+S/QRqYgoWZqpS7g
k8544v8SQs5JrijS2L41xmZ0K6W419+WC+Euzi6APHwpt3VrKdNlDpMw55GHzvT+
AU4jAv4OVPlAld2hsFhjy5fC5QJItz9ZWEbbqzINt6Z0KdVGD3qqjIFfRoXGUAqx
erMPVUNlBngOm6K05RcnW8yuha552S9w4JpbH8dMzW7Id6hesA9J+iGt0wfabvgx
eqK4I0lH9Qo1p5WwDTs/rRXOh1UOV39cHRyAjqT7AQgUWgB2PiD9a7Q2f/M+fNKS
9QSct34XLh8iRGdyM7k3OLxv7YLLvVPqM1VpdzjDskYjzDH5tFw7wbA6wYn02Ycp
RrLQkW9/1yx+sG8zRb0lCTbhX1sM2Gsw/blWdZ6FHszeNmP0JTDrlCDRYsy4zcp6
rQRD+0fBnfmuEuRZuQK3HaE2+86iZOh0kQsEXZ4QnyZXfkp/5q7kc2cFET+eCwMX
BCFoo+3Pmgt+W5eSnobaiLDTH0J1wyLjT/dErVO0ZneJIh5tddRDcEWfsdClFjUF
bzPwp8iZ+FACQ1qdfvgc+ewZJInRTAOk86tChNlEng/7vbkppf8YFG7g24Q6R8RK
/3Kw845PZ9har95YKE8sQo++QfVq4Wh4DBLocrqQuBB1E6CPirRGzCayW2hlQHdf
zK4AJNvF0msdGD7JLZT5wjFXZarM1cgIYIVngzwXJWXsn8AKik7ppfrXZxjvx0Sf
/4yFOehgaVfb9gNTsuLa7x4ULRGC9tY6NCkY0DDYBnr4Amr04jUrFWYQ1DXOyXnW
/bCHzLvX/xV6VlxnbhmtxUuCNqpj1VwGLs5JUPUHr7Nr7hZfkbXjgTIF/HSoP3xZ
/52XRSfELKycQxzkEbwZPMQrL/tIjuZ9rZxIss/hwkEm2F54k922ezSQddcg5Sra
IBiXMMeWaTnuhYI7TBsCEIFyTmB6jg6Jy9fnsXptT/BKI4q1G7AXNE0rJ4eUaIl4
1vhsGTj9zGjQJqiM/qciOBJn3YWaIBa5et5k7gtM8UGLYE3DnPyBx4KKU3HVSU1q
AJCHYL2whcnh7HXVX4dXyowKOv6LllM9tshJwWKuOwfHdVIP29wIA3WwKA37T7S+
53ct8HuPCqdWO0lUq4ixMxBlGGuQ7Y3AmM/cNNIebi6ivs4aLLeAWT4Efg6VA9Yi
hxOCTolI0BH5l6BTwmCc+Ne5wFVBhQ7qBshiS1tvseGkSpu3xer3wuuoCDSTcXa6
2UPSLHVHFzV3SxhSTxhEJeVBw9FM+6P+kTtD0rvqPucploY5jKHR+ME95ZrXQxD+
FA6aSboqTC4bgW0QCZ/UeMhKONTgIlAvIVQ2GX2gHVTl+/qmpAw7vK5Lj6T+8C3O
glEYIZp8VhX/vFnHBvVeZuHtp72j6IDxU/xyMO7P63Q7/6sZfEESjhm33d8UzDH8
Uv5xWQ61WmXCMBsINHaiB3CP/+WuXsbNTPNSSitWjJiBDLeCSZxmkzj81FC7XPXS
SkUPJ0/lFQJLj5NCpiKi0bS2o18wygnkxXysgBML4jaKOC7IuO6aCNHV/99iRJgC
SlBzkAeQOv9uJnZ39GNpnjIrFeyi9opJkJYtfMO4DIUEzChLeOIYpq/bMI8/hfLx
iJHezVKUFuXqHwy6WinL9IF0Ko0Y3IZkqyC5V/Su3bBqjLQ83nrp6OWxVEamxr7D
3MEwNqp0M7xRXV7KckTyYlqlQh7Y0cqOsYVYThnjnySa+ldPIq2IGbqErojdGBNW
oe4Pnd9f2opybgRghFT1cwBL0iFCIBwd6N6X8F0u/fLGgQf6ZVK7OyeKsllucT/Y
5VL+VHR6mnazMRXJVUqDAUwP5hXVccJi28sZrs7jIO5/amSW6G86zjokOqTvFwWU
yTnEKUPpXS+/Nb4KSdQyoNxBl7IdsicsjMkFiTW8Rokd/yN7Zo5+zO78f1D1Gt/Y
s02RY/GByJ+46HCvyNQMAddtVqdZxnlfOTkT04XJjeMiGy2I9ma/M6YzSNFGl+Qu
36vvJt8URcWFqXG1LOwefnyHOKEcQJF7HmsB/r+4Z01Q39xoDevYntSUP8QN6SKE
NUCiRD1pzWjlHzoC0RHPxFIdKlOGnt/gWASvtwD7h0RU2k1TPAYvCCQtO7a0rn4L
V3ZlA03mEbWt6NGaV/EKRFA6FhucKATjr5Rn5zvTHf4eyQKoN7ai+nbYlaTMcRlx
G+w98YnwU2D7MVPFihi3M2cvwLVUyqk+BEAShCQuxHcuJDTuIp+7+1ILnQ64FOod
g7oOdcxoWaY5HxBmIHlRi9y9jKQ/68kv2lW2EtroV8KsOmYZwXBaCypRPWZfiSbF
l1VsyBKXLAT4feALw7HSeJoQP0BoL4EwO7OmweHHhDjmWIs4kba6aLCnW+vmzCK1
4PGs76m3+G5z0txI2rEPPlbaFjSompeoIDM9zooaojq8MZUzdAvKHsYQLHsPdiDd
idg0AI+/e/38Xh9Vc4KB0ipYIIHAG/umLrYKFE3sP6FqRRBwEW/vPNrhPiWD/ez6
P22Unh5HmyLuvzZeYm+eaZmwHKCXdlRDtTpEQpX0gpqz0lJBQvqMLCxhK2ZCDgQx
nGMxXk3UhtJdWwn5rz4yRLdm8oNh6/oAFD94klqRpbWQ0NW3wf0XHDhWgRtqOPqo
65FCR6/v8bQAW1rZH7eA5CfnYtEEyYi3TqNyksSqz+PDE+Y92Kcdef4QxuCNxkNU
Q1LPtOafgmVLGMIfU6N5hpMCcztfCKnY6eF2JKdPXXxP0QoNG47W/hlg2dx0GNWS
WRJeueDMQkynbFVciVhasWsxvwMcvSyV8U4KlBrC7twQoyGwci6Dk0YDvH8VMSrZ
hmJ0RYF3FNU1tun7fyyiThgeG9x0povhbN5HGRqx7AfS7EaEBHyQLDQ/4JC8Fryk
eudZE/90hak14pxC89a1IvUt2akqJLw+zQcaZsoWpCTInhf2Z0SbgW1HqWUIUDX9
7xtSDhzK71KWNvBqQ7GrUP4AUT9Sq8do36Du23eFg5342HfLFN11cP/a3xF6Cm4I
+EgIVUmVBxBiLeiczNS9/u4BrAZLk6rxRoVDmQ98Ysq/D2q8PNyn7wZaujpJ8TAx
90n05WyhZDtE2w0KioqqclURB/jjATxtF2P5Fc8+AYxtrofcg54LYvN3phW3IFHA
i9maaS8xIuHbknSoKjRx2gbOcLe3cxdsn2I3DTHZQlMWyBgCPeFyHqH1sgrWaaFX
lO25UiVNPjImt8XGX+7rVLR/++JX5y1pBAlgPuG+CrONq1HDokkuk7p0yf6iD+XI
1ZazkES0WRt+QYEkh/Dx0qq98udSF8jQnaWkxPfous0ttZmkuLCG9y2Ib74EzRTv
BtilV6kVMwy0ZGqBzBrqicSgn8zuXWt6tHcBgpm+jn4SIe3Y32UDtpmyhVkx0vHd
4DKlDmIDkNYBDeL80ewruhd4jkKFXjd0l0Z/Zl2+XuZ/vrRVeyXlymbju3RYDZ/5
MfID8K7HUJ835GEZeGkHaFbTlpsThaBKwfBvH+rQLEQgkVfPUh/4YryASMUjNSTU
QHlMYiiyOUv3V0FYY5gLUN9ii2cEx/0vv0l10giBzPRY4OOlwTZkonacpy5Ji2Pu
NxFNK6eZdSRmqkfCPE6q32RAQZAj/lxrdsQbF+0Dv6Iw0Pc3jLuORq0xBYPG25HT
qJcWIs2MyUV1dT7M6V/3Y+r6uKym9fEISMAIaksjl3ZVceGLJNRhNmdYrcdzVJqL
S3BBnU8zhG0dTApS2GDwE0XuwOmze+j0VS9hZnpoa9vOiMGOA/6AbvOWQVTstE2X
fZVjTdIzJPezbLAO7QrI8CJcxh4o2ZsKcNLKhdBjoAlZ4hpw+jwbdSbGB2f+W46v
WndQLSloKRBDxsKaTwqnhPbQNent6u6mVHIpESmsHeN9IObSY2W2rgcmswrQq5Ok
o06oOxZDssakW7REeRMoaKmk4qPCQUxgVi1ch90G8GV912EeYTSV7vWl+1KIbSql
pXx09DT1RyFjoNoKZp0zGkbTgK5sasJOu48oWjmd5bMohiOfS63k78hT5rP8xPLs
ip1EQ/wRVXkNUCFGHyBNy/dnQnozIuZqHoqpARs3SDu+EkTxTmEEmd/YuUlgMaSS
HcQfU8OapsaEcqy++WLB1hsEsVVilILsIFNiEv4iiSa1y7GzL6DyvpfMh+I3Gn2j
JgxIsolbIGT9Lsur+68tsQzkuBkculCrcFz//2FrftDSMRtM+CbPDNuJJwd1WIHG
uqCMJklhvYz0/pzuT4/tbe11hkwcvtR+Bp1bLAjQa0DjHwjpg/3hVndEHgrwt3kn
NiXiH9kZjp5jbmrDVcs96/29vhHHnh8/P021tYcKEuEzP9g0fxyH8SgPLfOVr+V1
00h9Q+7ZQirMx4C+WaDKekR/IwjpWrn4efFJpK9mPZG/KCJ3qU+f6l00SgY6d95A
AJU0nzxe2gwbhg0eGWUXY8VD/rCMw/HxiFlhooaxiFxMlNDKxmiNsDLTIsQVnuSm
Cmyf5UPahofuUKwdOH8XNgPafm1z2J8ymT7gTTqkrE/JX00Ne6LSGr8tg50qVhS3
+2k42K81cSscBf7fWvbHqYybFLbCGI+tBz8GPDeseShM4QOIsu+qSchlfE+6dZTI
vdriAJnvk9bbNGdOpHXN0S3CfuUxtcexsWuGxAnEP+ODA/1XpZ0dZEVWk0uQdmBH
IEvyUPYQxRtngiEKz2NM1f3mQSH/Tr2DEI102usb++wy2lQvIeZbjancNaEyp2EG
pR0iUgVS1xEMqaL7jgipO5HmENztsNPzWOMjLjwkdvzFR0NRMMGdOtGk0VSKSDqd
1NGSzl52IvqYyXRxGs87gVi0SRKO0GezEuBgGI5L75Bubwl+A1BeKCG6SQpIYnIb
S29/2l11RJ5mCOlqsuuxOgHMNYHuLBUPWG0GoDm7AO7vtKvnlX+XOwV4ZIjp9pOa
cB3Llq5T3+VrSFZZmuAWMSjEIcnSeVvkW/TtYbVIJzx27B+NKKm5afVvpz1z3Gc2
mPdJ9KGWRnlIAZMrgrg41PGnJHRJc0Jch0RRK3hhdtJcpgSLxDI9HYCCq4HavAg0
YW935uskU5dEwUe5V/wt2MEtjTP2xx7/DhVvOkoIHQ5wcgR5mkGAf6W1Ojtgepg1
lX/JVZBzvvpMSjsKTAhld86gerLHDq01NxIxW4f3Lw3io+6SeyQSb9vESaDiDeyw
GWgRhxrJh4SNm7B3ciikSMfd2Pt+VPE9SQbpmhDwKSs0CJBBDN3JldDOUtGg3LgR
ObJvEu4yKJSIuMDi6H0CmGSSr+0AaJsc79PUrdGY+DzoHrFV9hyHv6cuPYcSgLh1
f/b2MZeIUiwdKr3aoTjvqFSSgJvF3i8zgnydDhfaLfkuG0IAStzDeJ8PJnQJuktM
cuw+clBGGZLcsUKgXRTmKBAYd2AlMB1gRp6WNTcJ5hvE5PG5DlKNeZ4vBJgaupwc
kC01MJLCZsWUJfLUKhoPdfNs4ZNJYWsrHSG1HfZdUSBJ8c7bVY/IVoevXQvtOZDp
vexMXL9Dzmc9hd2NctTn0YCxY2DhjgyJ/jVZhiyjDasHm53SHS8A9KX+kYvN7235
Aq/tJyo5fg8z2rD0hqYvZWRRlz0VfbidZeMQ5KNiXFAE3KbA7OtYhvMAhMTDDiV8
FpMy1gil+SwRQkXMHn5e52+b2yrX8yKdgDIIEiF8+p/TsA+rOGDFVJ3wS7GEA0UZ
4jLURfRFrI8FID+E7LYF8hYasGyaJ4Dpnuae8hobnv/LWDBXu/7fV/cqnFmPyL2A
cs/nnwgAACYor8ux+PhXmeX44hlYelJ0SxrPDBQAYztwMH0pcciybLKsN9+3WPpN
kz0kXO2FrJIoZ62bAekJwV0wgWa5U7J6ZEu/lFbEoQvuWHdoGLTM/XTwjyrrdibK
FdEZty5WzC0bZPGoeWfMq4IGxjU+DZpC5xZkkiNRjXzT/life80DTj69lIbJrQ9Z
TQwWBuwecEnrNlI0MW7dKxcfz25Ml69liREAUdoORGkJ6o3POdCJq/lX3nDLQYc5
6l5591OmeHcah0vtzzyojeOy3KuS33U/DFtnQiz3Kl0g1Irf272CNxSu/fMiJbIq
gdsyxIjFome2QraNNtVN5wn7/QYidI6aU3dmVL4RzWQSG7ItMVQI7qkvOPMnK1z9
8k9dRl3/0ZajE0Sbtm/r/Lhkj3JsFctqX3v+j6KjyrH0lNw3Pz86Y3V7pPUsC5GB
sG4TH78Vtdlry97GKEQ5ukajy+YQVB5AAmM9xQpdRxuB91rbxxSYY42vJZ32VslL
2XpV/jiVOpvX+kdZUFMJSRg5odQXcl4MC2cyPQbEDMi/5+vmtWI+57/XOefBMGhf
4cjvXjec/yVoFVaBVmpEPd2tj16X2OxESyLCqusWAWzLATBkzuvthTsB6UI8N5fc
vOwWZGjVvmy1YSbvu1MGyVMas8VRnYRucI9hr25xyvfstEnwF27kKTZmYOsgRNa4
aZNfDeyfqjgpWyGYy9W5dMqLo79K8NluZ2qX+OlO5JLPansJvvGszNGnuNcoE4tx
1+VSaMlQD04BvFC/L7cbpf+96/Jv0uGOGRaG3OYTFy+bK+l6zmuAujKJrab+yqwc
c+15uyAU7XmVubLbvfWknJkasVZ+smbYK6NNgMWyDV+CvR2IdSxGlhqfthl1sCt/
eLA/rD37gS0cDmP+FXUVz9O4qNTpQlh49iRpwDkj70u9u8JBnbGFs/twKB82UHce
PjlDtpyl1POBwxDNQxhpCUJT9XbekwqXVfxvlVyi8LMvWFj7r9O/aVM1EvSvWCHu
1bNZe0AJfZvqb7noZpa2jvorsKFkB2d1C9hJXXN25eT+9hpqdgAYtNQRWqOsOmot
l1wE4UDc/xFISrDbf/GMLrIkOCFim5jebVNzUNjngh33sC6ihwVNmmMXaD0nLU83
4F4BM6EsMTtrbKiHQry4t73kaT43sx6uOnBJ5PwbvnXLPcBMtna9roLFBqeVutVO
jNpNyvLoozzoFqIp7Qth6oZZJBVZ1h+CH+pvfrYOsm70D/1En5Ta3AZ0prvzygti
z/750jK2IG/alLThJgWhnxKTVsbzwDxcOk6JdGAxFBi4aFX+zMkNF2tjMOU18UE+
LA1HEIGmej9My3Y4zVacAM67xH2KLX8NnsCFeKIZwW9Uka7XIfMDeyCbJQk/vihh
KW1QY6ZGA2hw0UKBgIpdyFgrZtvFP4xgb0pRzNLfsQEnI9MTFz1uXo0ticPN46EY
YBhIB6ETk2xJiXF6JqyVOj4k8WBjJSUsNh9mbwdLmfYPb7TZw5aky1Ffnq5Dt+0v
jThFKbvVvCLe0euFmFTS/0hP2ng0fnyN7JcLqMnTMIJrvPypYfCldR+/FT3x8bny
3oVDKCMhBtZEzUw2WGY8fMR9tNdzGU45Yc9th2dnisz+gEemsst4DCQORnIhgkMx
tTVkEuk63l0OgyhmSVrVTMM5uhfrmUW7B7RVu/8tHL81QhWpHNazU+CSxeroUiNc
/5nmprNu04GqGovkqBJD0u2XHiusMRVIAwtaGbWrwBMzvWTZL2zlainC4Pa5bDZW
au5iJUg3kFaKf7MAVXVAt2IiM+LX3IsjuUTSOeY7Ns0qh9Tn2KAfrSmmz7Er2x/5
SQuYX1J4frZg4xzxjdzdSDWLU37h74vYgLY6MxYZd1jl4otT0hCruG7VdwvQWraF
kGqdsqr6Ndird6566hKLY0d/AHHF2XYxlL1nm+I13xfNElmSW9FTIJndj3Mn5oa0
MImtG3BAasMOgQejj+JeGywIBAsGZk2OAOkPVPapqCv+wkb7XjNWSOpoJIlX2zNP
mCc3X9AqOAVLiXNewUPdRsSPIIQ/ryOy9UesCjOGtdtMWjv/xlBTtQJSSdIYBQHu
Vmt6FE04Qp51Ml5w1ttOEprMROSpNbddOqMRBh8BGgSvg+CkATcz2wMZZTpI8mxU
8ALirGmsEzVOt4/YUiA2P6+OY2qNwZkmwpMM1aIlT5wfxIK9l1IX1m58f+lkFHSW
QUh4GqAY88GEqFKLY5B12C71o8hL2gNhDUiBA6zeDptvI+TN40MnZmCgHqeGgLcF
7hMXX7Jc4oUmd8pg/lCO4of5d+ydyeUq0DyuWo27za07+RHYWQu2HckjO+l12A2M
hAvehgDmQrdVa/eN5y7GxrI7Z/uAPB9nGKRw96VMik6Ks2hAZfhcGg4IWNti15S3
PTtWvv8BP4/npli0iBtocXlHCZ7/JhCVwOlxGFKonYAsxa1zrVL0impv8tWMO2rD
UTlemAYa9RufWk3ZizYCIaj4SNXZTG0u3dG/fySFDM1LoDd4VqMTD9Dt3y6FdcIh
wfIjnqqu8AgSznz72Ak2gKZoPztQJ758H0nmZUznax3cXKgNzxM5pQ0P5s2U2JE0
QeWZSDusLk9270E/sHDvpnraYASGAt5DqhHUjUuS6ymG2xpOcIWLrLNwBQAcXzBu
3MbOBatqIW9hy92JTWZR7hxuua5ovWiaklq1HiBOvHaFpMx8iWaq04XKESzPmqD7
+zrJioMiOuyy1/lPp/T6Y8ZYvJG76B3JiWfSBhPHt8N2Y9BEXbHO6TRfqDaMDd+r
mnNOeHsAH6XIgeVNMRDR0PS5ZeAL3RBZagsgI12aFJB6r6rzPM+sW5KEoRerarCD
mqJNMY4htEqqwz/Hjb5RS6/2YTxwJn6lGIwAsCKhbnVA2Lq5t5jWGRAC68kbUXJB
Xlkywka0t/GoZzCHngVZUYPp6Z85Lkk2NOGtwVd8cibX0ad66NcE7cvjTueUoP3w
IJprfG8W+KweVRxdYRddTgVPBse1yt/op1EbUKKqwQ1fEyExMoBOux3RFzKt61LO
l3wHluY7VqJQ98X6OxIN59KEcenIAHXm3RhPRBEOlRlxHrqJQkUwP/4bbXideoX3
gwawAnzb52Vf77DY1gVs+XPbe11F3BF7FxU82rkkYjbPQMFq4Cia2FewrPHX/6lW
PwDzBuhXEGL/QiJ+iY+OVQ4GzErOp6445ub6qtjz2XkkjLbRKtZKd9GTd7EPRzFD
P7ylPp6yOj48Uovwt9EGVQBdGZxKFyvVTBj6dytu+FhteSX9d1/i7qsMzHVZJFCN
Q9CJfILUynut6kv59TLiQPOMPPnFBUlvU9fW8UU2QAWrX9pYldHr4RzPYTLXA9Fd
PSLLUrEnu8qz7tY4UbQPFKM69mLKzBkEy/VVSx0RbEkg5omagfMc5exzze7xWGmV
ZfSgIdIx1c8OJB3E6ekb3b7MiwnvGYOpHNYhDSCToMWtgYJ2qm/UXu6szfevXoiK
9FIc54A2a4GxzbPaYBjo0UEadumWkfXKE+76oRWu8z5hC5xqiC8A8yhppqp506jA
Iw3Ak9LgJAJTozYv4gbnV5rAPYcD536y3drwrSnAdnrCD1N0GEzdzTvYSjgPP3Zf
Xno1xKZSlRhMf/zwLz0RBlwy9EMt1TESP7h5iPTu6QlGiUC2MYk2UjTLERc+rVaa
u6NElBqdsNkU79R0T31+dKhUqkOZUj9SNUR7yO7Zj0cnq+XgBnbZRN+angiqiOBX
Qm6ER6sZ1QKbuEq5LOqmy6e88okAg9NUFzjhujPOBTgTq1yLy3/ZgG/QwcSHGAxZ
1if8b8/wapekWiXFCpxFeH99GqJWZmdobZnObGCtQm8ypOFGn2BCD0Ad83aA/EL5
JUE3mIhCvOY+Zh2glcpm2x7PfqgYwsQ+w7VckH4rpF6N28OxgvufxQnXyQkZAVAb
rZLJDEa90D7ylYmeGWSfIhYf9T6lJdKXE7mUNwz6QgU2Ko5ywhgiolDBqZHm6GJi
oQTCGpFIRVasxjDoWNJ38O9isE9Bhvwb6SVZpRHRpfyxxP82zOQ42Tl6wZa6NLQe
MTD9ZtqkVrjRyA2Ht/sduFxOpIT4nWMeEGmkLBQsDfVutJkYI+qOUhG4GkOPcHY9
irUPASetHNLfeQXRhsLj53pzaFk9igUA2QlUwoIxvP5tR6G+wWuKKWPHtwk04x/B
5LruRlf86Crogpy3bqJu4LdORXrtY0ymV2DHzbZrOaicj81DXFq9ZgyeL8dRfcmd
cv0gNQbnUDeGJ1WDHvFtcqYatCEYf/cyoI4JpQqfIAtEZnCnFG52LyrGHJ5hVyye
06xclOBHz++IxmkN4R4TM41zk269gf9WgPke+NnVkww8PZGck1DTn+AWYWkTL9cR
e6XcTlhcdpy/DmUm23nhnDmvuadhHLHQXcgoomaOMZ8Lh0bRPi0X3JVxh6Em22mP
ZijLsoArL3+gj7pMeKKlcT4NRhTsnrbiwdGAy9MBpCt+8QJul0alLA9hRUW6Ei5/
4PysDo4PoKBLnxy58xFwiw+HVblqccM5O+UO591UQGo8xcmExZQySI3VvGj0t855
fgzZz7HoSjnGQhAgvlLqlen5bhGp3uFT7APPnPEBhqA+8FHEHfPDF1P+3hbCsPhA
ClFNJVL2kxtvd8Ksoc5wmpk9ejs2yYKqwaBbbX39ie/yG7oblZbEOGSZt2Fxd3DN
M73fzbmM6+mC1GD6evTMdRSWTiWzUmtkir75joX+imoSe/ioeT9CDlL3pyI6TsQ2
/QP2cYD3GdnfC9GUvB3MDTXbanssoL4+LREkRLRYENxHZF4hY7bkK76iTD1PWbpC
SUyXChlF0iMqdLeK5ZIoIWtPMux3tNkRTLZaEpwKB0iYwLPhmjbiISLkN4Of17Fh
Uas6DI9tanNqMpYMQdhnzKFgPVktUBJ4EWycutCva7TU6UaS90zLgQAOk5sHT1p6
/RQaq2Vo8jtih7XrlKJptljbjq3ekKl6kXSwD2njMYBnflbiTVIgC/PCgkeq0qdx
jZsBgtTWu8x2QaxOsyRGPe+o1Ecr4HJKvUnKCTqK4mSOKWD8vgIFHxodgc0OANUr
2q4W603jT7JF900+Trkq1yzCZ4hK48G44ixodr2ZqjhbY1oJ7UX7A4lwtcCHSpWx
tA5snKXRza0nl9s2NAheyBLmNDZIWEsxWwxGXPu6EwIYu6qZ9cIRdFDrRPVn/X09
IKwfi7LupCQOssaW3heucW4LxkVMfpM1O67b5vmI2dvlte7PBo9PwyuOLrgYbnUK
I+23sK6MT3K/eiNJzsj/UKSkhRciwM4lsyRO3QWgwKSNI5QpQreKI58/3bDYQrFm
MY2Wq6xmAXZrQ8rIKT2E02ELD3JNFA3cKVF7a9C+mNl29wQhpvjGQocuvfsLRmHG
XA6BfUsf4JgPOyVAUiXFJkM1vZo4+664qQ3eoIe6YD8xbY6qyz98DDpMfOPyO6Qx
u2DMoKWBwFWMmeMPMLiNPkZa1n8afQ3VWexd5nwmFU2mWQ+ZFwjXM3dUz/v4aJGd
GKaB+T2xJtPOVDCOEROtgT0sKzEjvRS881E+AW1Ww3uVOMhZy4seZl444H5kvQ90
22+LoBTDEzoHe9cG7UuGIW1SC0mOKLFQij73EuqtUIGYlCAFiwlEkLaLvG5NLf7K
AekQ1JhKvDpk89hDgsfXyf9vGSGCJna2RVb+P5xXo9CcWLnln7eQ29Um+gRFLDC6
AgvYiqaEqbwyxQ4r2aJimcExzVnlkZfjOK5GeEdjucCYYuHCASIlNInu3URcBqBm
krS+uhu8Vfus7/2rUIV+pdEaDWacE4nbWhpybzQ1WUOccC1a3kTz5+AQ1O7EzpbR
h67PiJ17Cqz7S8OaVQsBoBN1wUtj/d3EgNDrtS1XnPcZXekt6emou7F9oWKNU7nW
yCUpC7ZmujbD7defohKqiEurB0aGHQ3Qb570VaDE+AwN1Vhkc+OrKQq9cE9sJlM6
tK9WpTqjmCBKygnppNpJ9LjzbuFtN7MjFsWDTppdLj9Uh/0Qu0/ea7ZH+FPhLh50
2MR81QOjOycczaYi/Hm7WizLO/PslI68q+76uifPpJ2G9F/7nrg+gDkMG/oq0F6F
WYkAIIKXQOCxB4nvRSL67S22brXztUSVh8gzZl2GmfaHXmf6hIucnaIEDDIh38e0
vePZGmW9T6jk/TfFlwMKBiFdOgeHVrztQazETLI4vRSJgHm9uR3QqC0prRHlsCiG
XwWCoqMLglyZm/w0pxuMOJvji3oLbtfeVIBJMzCl6ZqhUtwLw01+VXSu68grbjHF
II0EBo+da8Ly7HSP53trVxxwiwbcNpsRhgsYbR9X31dVCveAboP2cBBSBquONp9Q
xwwyri8QfI+lZ7Ozjn9bCUMQwBMPf7NOm8Wff1mRwRx949TssVOWtS/q8Z/q7Wl+
AGyRzvw7wm5GOW+TeZNYix1pw/94ecoBbxFSgeucV+HEAaIt1p+UlxH6RTMA9WnO
xcOIhQ5Fj6pFz9lRdXePocaj65CRVGDvPfoi0F+3tw7SX7+y0cB3SSlFYvs0MZ/g
I1jDY7LHmmn+Vh/vhWPPTpZgOcmva0+8wpWmR/GxGYoFUPxFaf+a7aWkZ4kxOvGz
an/bIs+JVwYlijsTbZMqiG5T1a113BfpIXCjqaLIGbQlZ5IyZINpNx8r03VMifaQ
6jgYhqaOgCnVMYlrUn18JRmrMSzJ5iJQtunVhqlQlT/P7fmnkOgu2Sdk2/4IsX9W
6EapspBpLnZZeic6COamHDm2Du/WqA0YRc/1bUhOdslkhOSxrUuuiebbjLEOjvVS
4O0gE1tJLZDwPOwoFv/mbw7bSiE1etHdzqUzIPXYWfqfcqpl/fJsim0wRmgfJPXb
6f75zv4CxuB1CUSOYY714HaoMBospZdOHaDWR2uKyzlV2j/VY6ZG7dYpS74oftUU
nKBQZ91hpReE8rvGsa+jkWVoIII2J7wxUx+PNfWTJTzFeugStvEdl16kUn1pA5PH
fn808DSO9L9Rlb6FraSx5Ti/ey8n9QHBtg3NQBa3aS8GDIqt5tTO0BjfWlenKC37
1CG2CqRy5dD/ilkzTuhJjtj1PBQoXdykO2WHsuLcliOM+krQbhEzvDwvf1LdbOHG
wzL5M5PlwWHiGQew22751R5X4UVDf/h7ttRRN6lTnq9fm101wQKV+N3qs1HLux5g
hEDZVIvC+MDTFF19P47pc4elJ7l0CmU/l8uDcqfbmGAjD+GlHzjjbeMejeRqptvP
16vJePVfZnxyQ1g2BmPaklskdviT7aAuVv1FabY/b+wCWmuucm1tigGmd+RD3+2r
gGoA2DhcKrHY3LHhV4cjUz5Ig0rgnyTve6tMc979bhcGpaPbL3d71BCABydJfsxv
lpKjxnyXkr/00TMQjNfIgnuqbJBja2f1j+Bb3DIfybclpApjlLRnKBifnZbioZPe
tbfqoZH14Nnwg7Xsmc/0VzVt3xX+On/mqWXTZTE7l0Hj8gsIZfbTQWY4ffNdJXsq
c9jg6JWqJ/DcNdTcMNurOYY5Bz8lWysdkE/TXZKqRn+Q9UvsmAsjiyAWT2ZDpll0
PD2OzyyclwBkD2madhH3z1VUoczO25x+qVQaVbRrsxH2uXO9ze2t5Azv/KWnCobf
G0WzTV9SwZ2PBAAJEKI/S46PJpDecChcB/YmBevq7/YWzZP+tnK/y97m90d/9Cq3
dbi3pwVhvBJfvdA+nWcaRE9/cLJf/ZvYGeP5vPhzcap1QIyxwqa6uoxUkFYbPkai
j6cVg0AEi4nuLzaD1ehh6Ak9GSu0QyuZlqSOW0s2wnFcOedk+aUnSOLD/qwzroxN
N6NPE4suv5xZH7z1YCua2eMRpriPgPOc0xptf5e+TUKgc73oqY/ibM7+E+3F3yRQ
DYrLfNJv0CeicJdDf8VazSmRqgh2IHi7AR5cs/Ueuf46AH7OB25cFdcIsoAdoIap
R92alHHa9Q8KXAEh85MLGXtWYOeU2dr2QqTxOveTadEMEk0MGETGHE/FG419002c
Az2ayRTDQliA6sf99Zt/S30BazNLuKZYEaKJZxTxsxft7+Qgd0J42pW+s9vPKpaV
kvOR+ybzDvVmmSY6V3Fo2CtlW+HOt9wg2DEgvJeD/Wr9Xij1yFdnVVxso1ZkRTSq
Vaz0HUdNSLukX424S7OCuOh25yH6VpDLURyiP7J5y25VWpFeOe4u+wm5rII2uSUY
VM2C6KK9ffNa5MYjnd8KYRTfm8xuI6hAddddXeT/lVco9teicsLbTrMl85B7lpz1
9uO0ZrYv+V52af4cZxy4JbjMlGj8yL478ZtTX+WzJnEPcyWd9bLFklBgc1urM0za
3X7fVU+2TQ/dQG9YzwrHs4JBY4CXJ8AfF3cFN7EsOPZ7HHO+Ucm2TQ1D/n+E0W5H
xZPxkoVMCDVxNjmJAtKZ4rTWJ4i4R596mdSGBkij0U2D16W4H7+xsgE98SkvS3I7
+fbSBWxAm01l6hN3KpndKSNGevQDu+PbYQWoBqty5HVXt/s2hCW35TAcKx73+Lrt
bBrXY04eXPlqd/nFdDb1ACdhnBbUucEXfn+7AHXCUHMXx1aBV+Ufo68HggGYBkkJ
O0N3teiEN8Dm5F+EppOtDGG9+h3yVXHYpu5D2ZsNq7OhksVWzLrNCSW5eAF0J+2/
dafXGRRtM1aAzoDJ2xh6JldhMiuT4qVntaDH0ddPNKd5Pr9UIm4Emzktz4Dw/2BT
IfQPZ/vfQPkstJEGYWMEheHAf/2PyKno5ROoRqs7hBlUxgGynN8KBhdyud2Sxd12
0Zan34iyTWK8/t9f8FkCdhE8DZ1zsKfYZ7cAT4j58mmF9sNUIBZUiuYEbQqQ8sbN
2ccSdbmAVuDunoC545WZKrdRmI7CBMK6Srpf1jcv+21mGr5j48GEPU2w0qmV7d45
xFOTD80rNMr+IL4hMV09FJzOaaeNu4bbhFUpi+0+tGnjS5zVpNeY8Pnk3GEAAD/l
XkIC/XVQA9wndSU174hCAw1R6LBlmn/I3wO9W1Ax54D97GosqKZaBWdsL9HD9ZwH
qTIJ487xQBOYQ5vKVvX5qS07fiiqNwSVDWXS6TLyADGOjUHrS0qqpcWcJKQ0y7I9
7U5/w86zQVY+/Y4zMGZ1dtSRjhEn7DuyNdEBOrGsrmONlPcUW6LmSgpYsxbuDrn2
WmhfhXAbLYbLotvhyp+VoqU1YWlaNxibkgTHW9OHmQwHzGPEb0BAegl5xiBCZhc8
fqEYuhecR5j/ojxLzlvVxcCPbpqBsUCVzromOgYFkdSPjpGBPOGPHf7HfSGsWvRj
kpe+GwLyk/z1fShCyIf1J7Xp19ebuybl5i+iSrkAx+257PvQi+vEBSmUK1BM+cwl
Pfw75NvLDyyk8EFnNZMhPOcWJPwsALidzegg4Xg+MY98qstYysYrn2hHXlPdhyxr
ZahhBzaIGLqt3jHJavAUzxuY60fTHwSKSiCMxoimZ1XhTSDS+TJuR+rSgOb/Lc15
3SJBdYmxU7/AhILWBMy/SlYrd4HdQ8xqDQshX3zVAG5jO86ov/wE4BjdAv2C61/B
muRJRELCrkpQ1FTkf8+aCiM4DRBjq9KjOoGxWPOfP3t8+8A85QdX0QOjMiNskLPF
yu409NuVU+rb/pP50d89m6Ily/OfB+gb6sK+5337Asv8nK4MaAig/DiJk7Pq4TPE
2dBWu8wQFwbCv1j4AyEfA0XaM/HtVNOrWSIe8evOiyvmsJEAkWPJrk5fGWXb9xmd
f+iM1nKq6PSQfRfN9uqSJjNnm0QY8JmDvNKy7A8dIrMaHjPk8mI3nyEfxSpW6bNO
/RNenYsIXfCH/11Dimh5cx8WJkOPCqzTQa0j2ehpOojBh+LFeCV3UjeGFKSBu5FE
6iZYItiiESvwKjPY7rSvtc/3wYBBrK2GPK4jSvXZDnm+7iW+cVPob+EklG/al907
RpfLyCtyKiEb8NASOdZmqDFTp9bgPFyxIYXJv2dj6TROfa8SNeALdC8lqi4jR6Jw
C9aAF8z/JYs2jw1UtCY2zlAvCMH+cPYON1ZJBNkvfM3nvm3sYZs89k1WX5s/fEPe
89GpAdgtvEt3wvF6zwozCgFSSpNb+PhNIeFq9qNzJV4OFfOWX4gwtrqsab4q5Tmp
pdQy3uEMUUS3hJSEZe93vs3RCiO5tEkjBBUTplXQj9LFkQRDyBLazUhkm+l60uLr
SNABobZFfZ3/fAOOSDTTmBfNLBN9sgvoU9+YGx8xHc64Ln4fW0VnrYhEqU8CdlZa
kSpBmYjj8OxjCa0dWDDc8kIlIJRHaLdANg7W8C3JASihN+arYLhlq+nRXnmRe+GS
LxGxCEu4OoqBVl5WzpfbkSQd1nrlgjYpvqZNA1Ko7ZjwUemH5ku0HurqEaIkQaBv
620S9t2UBDn0MvQ+7/q+Hyb/JDqQwZgUqVglbTs4J665E02c0Pycb6wtuMHy2Iiw
DhyeaOybxHtZbG+1l23aihkjPqdO9fabOZR5gGcHjWGLLj9kl7CXiWGIlP4Q8WsF
J4V9ZuuN2ogvGssXEg9O7vJPJtp4QjeFy1bMxfG5jmUtsKDWybEn7jls2DXdfo42
67ZEEOK/0XVEpx5DjyLbc7GfX/fglsW89STdL7PEACDnv3gri/4tdhKhG5JIw2mR
xbd9DctmluMeHNbUJt2fGVOkYZsDdAw4WCuEn/4/ebP80a0MKP4iVeknr+4PjS4h
CW9V9BvVy02y7uWNEOSNjii0pv5OwTZqpXy3cYfxPTIllNBPjHQDKrUQRuC1Y6H3
A1PDMWW+gwMZIfnsXCgNFlY+t03JdDPQt4s3mSlyi7gShXHXRIuwOsrp/0A1XD1K
xyfrtG1S+YveQYezpriOkC5dwG/D3G4mZwROjRzI/MDk7s6/wDB0A3eij7/gCw4A
lPU9qWD4D2//Pzd2MQuShLtG1uIuIq72k70isfeUWkaaw9gCEOyGWy56mbMdoDHC
Fb5As8wsLp8QGu7CKa+LsWDIWqPMkdfxlqs3dxXOyqQl5OqZNLH+FMf5f2C0rNix
iTttC9qhvx+i7YiJm+2QPTFsNO179kG3orcVtFOVwmiRIsBh3yuUPVnpAMaHJHIY
0Gd3RCe4PBct7hmGZDMPGMW1nvJSp1xS/b7CIW4uMkfkEEASe8F0tUt8b+UlDoLt
l4mu1Mf++ZM15U2V3SxxQEEu9uEO5ajBnu2d85S7waYVQXakLHFwfjNZ3uNwSpeD
axqjcKxGFk1Wv/0l87IgciFbZ0ypWIfwGNKiUH+gkyjnOLy0p37VFcpP91LQ7tUj
3NDNYecUGjaMmkg2kym9ujIqx5GeCTcndeU0W0U3wJjNGNEAWKtNrOmj4ZAQ+bKV
hOUknLLBJT+KCEDfqIfVsIcnJRVxGiee4/7rflsi4sqOHe6RL71f9yl98JCsP7/c
i9FIt8C0Y/ayBwyVKd9EEPXzDxF3/xVWNGjgtFdJ3dkheiB6Lq9TcujGWNNPXc6U
b2lOO/Ms24lxs5hxCY2x3qjOMyoRC4i6+cHlkG/QJJIVLe6uuYdR23VsxZcedfvO
Y+2C7lak4+2Q0bgCVxJNoxscb5pvBVXaUtfQL6FV2XrCSEVqwB5Yrwe4kA4xEf4H
RY21Lxc7MWxzTFHfn0D21Q6HCIJzHv7WoamNHBpB5kd3/edAR6VjKdXAC9ld6vrB
0+tf02OmpY4RsR7TVMfKsQTwyaAvrSHoiqcSp7p9mYTlQt0n8j5zj0vTU1JWir/G
TRofKw+hdqIilkAbH/MIaJUYhrt9uTfctgxFoPITmT1uidmsd4JhxEEGVWEgFQuU
YZjIeV1W5wwiuQMrcxyfgLidUvbbnFlvydwiumZnrssauYeoZvldgWVbzKw4S681
thryNa4+xmFZYzmXm64lYir67fUodWJF4auZdlO/FI22hm72nsrIZrZpoO+ODl2a
bGjNHoe9fORvklFPJcNwztJjSL13tdgljZe5+NbZ3tpGgHEbEoPUnOvuSV8XePHq
pf1CWBCxYWCK3BJRCg/0DLZLKxe8nWbJoKPX0HT0txuNdI5sg4j1AL8pOUk9Fcpi
9vBE1yUOlelmq+m5OhAv4eLRARbKPZ8Z0j/dSKx+KDj0zJNSFsvKAl7S4TWOhhxK
5dJXKsb2OJEhJEGZ+KqrVSTklH/uiUUym4WsDI6uXLfYkKNWUVlsB2VzclKYH8CI
imdzfnME6IsikvuxfK5m6LtEaD8hBRCiEocWJzMeD7Ur5gRXQA3ulsnqzMCV8M7E
d2NcSfBCtO58bnvQedwKOsYgVscvfR8kaO5CdITC7d8jfSQhRjJ2S5TMA7U8nO8E
DJTQbnki9DP2aQEgE0+wZuh8m6sEJ0lA3iu/zihEHicCahh+m4gLl1Dgs7ZcGNsZ
SRU6t6kii+CG6BzFQwkidCrnLC1UopslcFHvoG79weQjEIGzUBUJm6GaOKqGhpNO
ANeO6ioLLIndp3QCSFHNbYNwakeb3O6OZ9MyhBavmhT0ip/CUp7OLy/VfXPy+bp+
/R4hIwwG5OPt3vcAu9UmgNokw5HKE6hWJ3NaOGIwgDKp5IeyUSoXXi0bAmWSoJBn
nwJnTAw03zcvXdtd1brxCQM3SgaYZ6V4EXAYof4ACHJ4a6JyY2fKpf0XyMlBqXS0
A4OULztpB++/OOFxozkcvvfXcBra04njpKX5ffxhctiQPbWD9SZwTTz+cNAiwp7A
upaz6nVcnt5lO2OHhehP6Nn5qNVKUzdw5UkVRfIqpBgMJd3XO2doQZmsnDFOUkll
7y7SXSnLndMHv0sqAnn8jevdK6WGSNKg44PE79J2maRQejLx38/6GITMMxmkimuu
y/Xw/pYGdwTVD+fICjsaLhDAByZoncDR3IXtyYVMo3s2XF3aLlFNgcvVrZDFFSph
ApOW4/fSOtCfHXynXNdM5o2ncncvaMjzfdaqqLN/5z8jEs+TZbNhnE23OlEmQeov
LfoHyRzzHaEpVSSs1gRGLxM/2hwDgxRI3uB7otNeQ0xaXumZefTuMROxtvBfYkEw
VXuCtEl797ajQtf7UYNrIv+dD7AV9ryN9tUefwnTwe9kwLlVrH+mOAQpXsQqSmZC
O9SGcMT31XftMhmJvuNxIg8w2RAPNE2SGOtSNz7NZhgnXtoiK6ZTLUo64WHj5ESD
AaDpCiogDqIjOzEmWVZzodUfWHkGckj4kexOGrVbQ/ehQpEOoUiJ0Cjb1Y6T+CRm
4ewsqizzBJ9rxtF3rCJOya9LE/gB8x6TuewAE85cXqQp/zg/3M/sIP1PtrN+bKRd
8hZ4hQfrW6TvCH9J97ODldGqUPtURVxUjy6D5TW850IG+Ow9bO0lEebR7oA0JxKj
LlFM9SoZm+UMcOAIH+moOCv/GvgeLp7jDGMMh6NebBSI3sesDSajPK/eXYzXGseo
EgUoLJo+uuJyHVvIbfJMmGgecsx0+d9zS2iyp+XLDA6wfVlmXF32EWQ0EiRPIe25
qqVwKSyz9jY83Xi2NRZ/RYll/HbnSPHeAvleMOuByxcreypxcpFe+BzLkLn0cNiV
K+r1ZDZ12DM5mHrsE5an45FPkvFkzmc5uFCvxV6NVm5OGIzHxY2sElrYrdfJxGsp
oydx+P4DL6cvb6kI7RLV/CJz5pW6OuAzWPpFzWFmHjz9YncubVilsMQPb/CoWstY
YoxZRkvxYAq7IFgl8WYDTAR2nS3a0FWaSXtIqGuOiJoxDN8eWWb2E/+aH9M2OGlK
cqvwSzE2IHyS+1IBtHsI1gufvfTac4EQ+yaL+aRZFrE8qqKtTWGRD8GJKqknNHxT
aJEY5zMQTkkL/cQxEyX+fvmlZugatgQUBPBkLQNAy5G0G3yOKqpT0qeJDSMVNReP
blpyxh34dWTr77hCMtz2IUEWQ5mrUTlIMmPQpG3W7JjdZXaZJw+gZdoibfAWlCMi
5uHevDuC97HrnoEVgCGmccdXpL0ZfNnE72s0SXTMDAqYNXCM4tpIBX5YUPIhvaPi
+PHUuVUNGq7ImWVXMsE5mbdL/L/adaRfszJr7vE+JgTivEvKe+JZvOIO9mc5kuZG
Axi1O8UKmNjBsqUZ8sk8JM1iIW+YST0qaZhxqgMdOSajEB8mt0IOa1HFzVVbLcb2
he1ILcJF2TTCzQuloFULwnc9Ul3dNUUlauvlDM6pA4mTWpgXbhenSiFqkDUxCuTt
MEYSOfteWEtGp5WhLnawPhDiWiwSbRTiqXYE7vZxuCldmazRC5WAxECU2Z31ahzL
AWFYRhAtiYLHFTHntk2ANAt+CVr5c+vjoJJE7PL14SL9ImD6OGMjx7lvsL6zYTy1
fjHzsAK4MBPqo6kFzUtPHIgW+tnVqOuhHNDULmDqImLvxSmcu1FBR2ssFg0cws9G
yGW884ulDqeKdfZrigKibL7899bgDNA+64tdcIKMcK07A3mqY/xAJaiJhShPsI2/
FpkHdJMCw+5gRtN7Oea3LAzrx04ZhIMejP6DbFCoS3TozlE+u2YUuvQzUl8NLnLV
/nWFmnwkUSmKxtdqgKpUnvW++ncZlwmKq3yKfGQgzFIYVO7PEQ7UrvU9fIjiu5mt
UX0WAedDG7ewI5qFik7Ljni3NlaUB5Sy9wlmTGmTQpOMItaoWNkjrSdgkuvBR5Fi
F3vcyVAsbrdSt7UY3RJUftjCP7h3LXsPdwBKBw+Vf+eWqfM3J39LBhMS4pTDHMwi
vb59WSwHhwqe6NyqRmmQ2hpuwMwwQV7LwrDKHvVCZJ5FBD3GYxxQ8AjG5cPUvvOm
y3DRUbXa6J1aFrnKaPc0fDXRVhZsSixJAUOIPQT7lFkOfMm2rUk3nI+VaPW96rt0
sTDhmXUZorf1ZrLORGFbIjDZwwq8F96EHwZCaPobd9pSFD7H5J+bnqmNNoZN79mv
2AsLzNWvaoiIfKltv9CTGUeXZjUw9JTCr4Fp8PY109G4y2k0GlK7lQcxnxBPhFVc
n0UPwqMYkHDfaCcr/ulAi1OMhhHQWd9VJDsMUcfQAd8rkyXNBfvIEhMQJy5VX4iW
oWuXOzEnIwHnO2aEh4W4M9t9qXJLSBLwSTLDZJvj3jWWWf4UxxSk78d3abiqNPm+
6GnMdSQR5RUvx1ZRceBJvL8SHdRgr0SrK2q7wqFKoSYB16QGJPsdlSL1Wv+u4Was
Y7KiygBE/P/zesepADz46Z439s71J82UC/U/47cuLWRT5Yib8U0p7CPFtZJh3AWu
2Bx6+nD8dCjGJwNVJaCQ360Zb+Kp3wIBAhnDYW7htZMXw4LMDp0XDAmJlQZN/n/E
8iz2ZXKn+1iSPD69QmrwLFPOd36C5XMY9hlMEkXzSDXZCR5WAqa0aXvPDrI8dUYc
qjA1ycfMeiOkzlPwG+oDnSiYwqksvut37rfmH5nIJZDhP053mMB6R0Jn1GrzNj0E
EHiapDqjZmvgC30eqzumb1pN23rt0YJJoSZcuSl/39vcMD5cNcJHLJTs7Z5LZZP5
eFFkDsJW2RXRrfhGm1jB1LYw1UeYsBOPwog8eIsH6LHe0O7GKxDP3UFFtFiI9pZc
cXy7VxGLpUfZPkwyXzO+Ex2ZmcKdMWNjOU9xsmsqgJ0SuEoe/qbIrk83/H95a/bl
Q+uQJKtvoviNM80iggsyTcLNSyKg9yMMicZDM/wS2853V7O6dTWApQEoDSHDGqRh
NMfacxpOSU/uCZGBoyGAAURZrQGXjl+fm+16cRonXFhUkUhLrZ74V4NcV2XAtP2Z
VFKKSHHlL1WHIthNOQErVmizsHF1CYjJDXsA0uuDy/SgnKnws7lEqgKb3T6uJif1
U/FzpKfIBSsAOJdNnxD7UCgNZW0JojxAQHJVvF5bvaHt5NJyBaSZ9F7NT0rWDarr
IMJurOBqwUpVZIsQZJzedLZ93OuMHH20RjKb7GROyVllnYYyHlE3u9A1S73OGgqV
yrJVPMPgnCHaQZlZl0iJTE2Dj6p5wUNnvzOelAvHG6MPtPPDcgtPQ6ZlZ8p0y8dK
jeeGphen6rvXeYoIIKWcTxqMI2/dqJOISShble4DJejBaCZPCa3SUBNpHh+9RIGA
chl351sMIM9BlVxvwlWGCNtrfXsHRIWFkOYUoGLh/yp5V5jH9jsllGqin0FvfSQ4
xkqlZjEwumTS//DBcyhbOHQ5x8AsvJ1I+8TSzrl3pFfQ1pbKLvYED3JWaCKru+IV
oBUSkg9PFEPeUcjBCjWHb/2ggi4qAQr3M+paLwH/BnVtMtlHvsUeeL6Nd0/gfXES
tMqQ6Z9MkAHBEUV/t/tNfGlpYEG5kaRq+fnmwY0AXWxkcy7ahyuQwIO3RcQc5bMk
iGhFd/YQz7yDCabin5KKk4FGQIkr92CMPgxFDoDOtQbLfCId15/jRvbNZ6RObrQM
Bkkb+wy+XEFyvvzUufI7i6msQP66bNRDNTNlgjERbXW9Bei6L7jv+jN93dUc5UbJ
ND8AjUDbhAcIgUuynCwxDFiHYTSfCD5eUWATANV3zWlP+Gpan5udwoGGjMFVKXM0
BxUwqEfmsyUgM0GVRwpAylH8feYgp9hwMNGBLie39fp3EvuS5jd8SvHfu0nKHUvF
BA9ruVh5xcQMztY5HEH+bXHdNv+n+eQ+qLlUmCDoK/kpt1IKR9Qf/PgYnVw29rdQ
Yw3B2sH/sxQWPMiH6KUTjHwCvAXtjjxiJDCBqBz0YaFmsXsBBUWZiHp934cWr5jD
YJVscdQdZM68bddnUBAaGH2Fvm/ftpMpy4PkJJCA83Sikx12EZSyr7QioxNKlK0U
kVc7/Lh4lyBa0+icBoGF9BW0kwqTMprEffI8+9fiOuBCXdy+JEXlH14otGUkJckN
c2Qb1UvqRy26MoCG2+xHg/nENt6gaJMOUAXWEj26naEaWwre8GIOmE9UYaUalFzu
ADf8OHA+WLWmYS/F6YjtGAuPBZ4KMmSCdRczt7hfrfhky4K12rm9bQBZ4BNLTcL1
M02WIzEHuaiGwwCVAFApKOwomj91L+rStLhEtubmvdUOmCVvKeJ4axXlloXqkaQ9
0gO9L0mtsFW05KkPacSHdJWLcu1MV2HDjLoIjJf3WiWSMYt2nngvAw+CpKLA1Hpc
vgnxcIkL43mY79tchfeoDgM51d22cocRccr26bJHvIqi3QDSDKWqTe0kiSyrmdNJ
zRkbc4cu1cTza90UFGYqHTiSDH27VEoioNjovqVz2SGx/0axFofkzOBgxxoJAXFH
Wfd5aCV4tFUuoJxk3UiQZPJss8LGvnQ8nhkHiNK++unxeRFStS5szbRPp6SnmPWT
NWP6aZnyHt7cPCX23CQYz52HX6NmzMZJhR9E9xfKJrttUriHKBTj7Feq9kdos6Rh
VivUyQfic9sfE9LPYwaUO7OzF1O4rFP7wuVhlQpvRnF5ggmt4AYvPpNax3/QEJ/K
wmn+rsMW8CUAfX8twks1mbHZx9tDABEfTtgZiZ8UWLbeHJ3bu3YZMA7Rg8GEUgkQ
Ai37NStMq9l3Lklyw2eOxrWVptNpI8NQ9mT1wPU265fYypKZH1YVDcI3m7cL08Gp
8vxVYm0aA6dSnp5eYzUmwMhJGUVntSrkEFt3QXuIaE2JINau8jAP8oVIEi852eDb
z+6obr7TPzReyRDRAAtf43bb7Kas91uFm0xiPtzjLlxm1ELx234RKZ8dqaeeyu47
ERWIhOyqZO9SqkNvwtzGRdlQsAzZ57bhlvJMBwHQFcrVHsl0OrFNPR4gk2pjo//g
eZ2L7Fglaxm7m2b5Vt/g+Jc/FYLSZG+CVWDW2c7NvwxxPgn7J8PYI91/4UJ3XIrZ
noU8eUXvPMvrWhyjlqaHoX8DIe9fr3dzkRZ4bPcbcTo6MtzLK6OJrv9Gil4jgCtS
mdKilBRr7+frW4Fn63QPTdAEpPeTiZW8C/cR8GtpJ32uGmvPZcY1ORrbiQzS8rqE
ZodqauiAfK5Kuc31mh0I6DOkPDxPf453OKC5NvanaDkrmtWwnJYhqI43KqebiiCC
g36rTm37vu8X/QgRwV3/9sGMEZfEYzRQEaHtgwf5fLlcU+5fu6CiO2CRu33Jo5Og
rnHphrjGN7S/vYo+7+Rb6eLMw5C9t5nbj9r99ASTBMNOuZKIizCAUnq2vNqabF81
U7T9PMA0Nt0Sp7v2K0x0wXqX231QdyyPOu2SWVY/VuLFvxp5H/aMserZ8GRbBmd1
hQoaM56lHGO3MCb8o9PhzVtpY+vU9erYs8buASIwPYI3v9gSg4VF4jZRDtCPKzCy
9M4Xdh71rTWLRVAlwp7yVDdjljQvspESrTPzG4EUPiZ6ZRAM1KmOn6Zw10vmyl3c
sOwd5DBASHWf5l5TJsrLH/Npv11GD4vknSIfQEvljnwT9oTd6z5CuCmcb00Cq8ne
Jnw1UxDZsU4V8i7y0Bd+0ZR8ZF5dhCwBj63ORSkUpk9AJ/ZigcihYvtKKDogPYX8
rDq/6HL7abyiScLShJj1YQ+7SaAZsK/4lQmxqNTV5qOZhcYijGye0xz8JbPbi99Q
uMcyonh4Fq9f9VQyIwP66Yq0wiAZnXib+fFAe0l64C7zxm5OC+9SdMb0/NH7ERog
SFg5y9SMt9hMN2yNQJAXvKgXaY5VqMCtlpfs+pJdlOeZBXYsTDHlAkNzYhHZ+nTB
6W5MRN7uOVvwayE9RCr/+QlcyjrQYlhpbROmg3u1JyCxLJ9RDYho9Aj81woz+vEB
wBhHub8MCEr5RzE5orr2ec/Aqk2oKpuFj+d/rr5aAmhzuC1LMhPe2O8MkCS6tdG0
RTTNue19CudmQ0l4Y4mNDmqzeIEYGkyqiWGZ/5QKhvZLHN9JUyrRd/V90pbwUTDH
hVU6Ol2uibW4ZYgou4KKQ1XtL/n+P1nRXE4W+9P8wI3IVlkNwEj9FOvaOAtJIWib
bQaVHOwTpWG0AreLfV3AQ2tbqt4p9wWw/69yW85VeY5r5CabEzs6UUuM1jlXFnRS
UVgcTfXWke1tDekNOyV7IICibuSXxdz3NHjJdQsCA81HdTJO/DFCMwmRXXqAZE+V
eIPPWZ5LuaIljd4OpVxXLQnt1H0LhPJ88hB78J8138CKRVWhFi7QEzUtIL30HjYC
YCEfPE25wMwcD4NJ8/l+vFiaOwLuCnVZOGKYRMF8Uy8x/L2TdRFCdnZmPfhJ32CD
9wgNar1UUNAPsCiKs0W+i6BLJau1PnUXI35meEwzO44BF6XUzfOg3GcdYODL7bna
1D3pELSSGKSDGiyZQrt9fsIbIzaBnBY90ekIPzTpxzZ+6VY3XLEy63m2VlnSVbe+
iRCcCm8k0+2rbvZx4GnoRFxWN89JSBhDf0SCxhAo+bW4J/htAz2H9lZcBCyL7Xgi
3YbCyFf71JsKDJ5FGBHsRIrjPAW1Pst1aeAwB46aKtJ/BTHVPv9jWbgtguuzxoEr
eIsRWc3axdM7jx3a22qIbou1znpNI8mWiDAZ3Qh1aIoOTzRmGe9ubl19H2UQ+4Tq
p2/iW3QgPoLyOYFDaaGW6qH5It9jjL5mLvYALUcExCvZhfoCHP53r3DaMIma0u4C
EpHLRr4O80mTIiQKqPHxYtM2ZT6qj3FJHOkrTurTP3INKgpS1DFU7M9KM68B/0t3
C/K1jbhL0wGNIa1e0bkRsu3R/MN9yekOmJvD6g1+ZBKHimiN9IhxoLNOcXgqG9Gf
JZjcA+XP7h6G4ha2UsM+PjX+IZG2OPSFUHhIomQ5/Asgjp1xuP1wutetlvHhtn6l
B+WdRQoj1VJTbkl1AV6RlAYOC36lWB6+rZO94tMKWmWFx+0ljh9W7KzkWUsJU55x
fTs/HJIjpQgCbki6zqWHPiTXuE6cCBJhaylzoigBmi5O5ZAvCcHTCG+aXbNLmdtD
Cr+4erjFZK/ClvS1fr/gVDc4FCvvBz584uoQdP0ppxfO6vUVg/cDwxOoH9Xw+Z2M
zLHae5OEan00/gVRFs+iZtFkO2EljvX9V/insRcLVhbzVuDgtf8QSdqdhpxNLKM+
dpW+fesvei8qjqYs6hKHZZvTcC/ubagkj1duutPktKFCenLXFQooIPMIK/gVWc0P
qdi/HMqtd7BcTnSOUhSKLDoQeB+qOuopOJ8tbuO9hjatJ05JDw9gkfg5VbzacEyk
yNTI4TctME0Iy4Shw7nuqox4hqTbybZHbL0Y2iRLej42nnVM9cG14llIhB+aQUTh
xUPK1XcXmMPe9fRxAafLI2B7EGTPZd/Tkdfp3snFWrbCkOCETEYsKy0fRsQ5f0bO
Ftg3+Wgc5VJbMc2im6GoWvTOtzZdbwbxemH0mx0ivDHTSxN+SZrRASNwhYLGb35V
YfELhY29UR/OKZpomwVH25SO2e7OJp34vaHr1vwnk7qL8JnvS5BJvQ4ucPsRjuvE
aRLF7ciM/FiNITHeQZ1Hk00omsQr2Tff0njyFoFtD2Pt0ktQQqij96xakOsNi0Ln
k/Ad+MSRHXXwOywzt/QWhKutDmDuKgcjlmlcQJRF4upYpziKyOkcqHEarODjRhVk
ZYFtsjAnqo8TZZedmq2uY/KgQeUtMV15Hw43oBxrLUdGXYjNQWHTZs3MwKg88EQi
AEiTQMuVl/ld7MflQx8Cc8mXWQdanUlntcKZAkqMT9XLPzXkknhMoDmb77YAuixZ
OHs9FyLgn1xrKwgFJISj8g/YObl6Et9d/hqsC7cFNwQLVPuTRE4SA5lspcdZn0p2
zI8dZxzeNcNjoZJOJnXyIoTFI08tM4ZFIUgGiZeCFgG5oSJHrL7AwsGjRSl4gyvE
nfQ2Nrb6fTK32c1aH0rqiJXPoT2qd67LGt8e7L04FH+s7Ahx/MC/a2Pqsyn/MeYQ
pBRecPFJ5dyB1zlnFt5PIXoHVtfqJvcBPUOD5cl9xsTYtVCNs38t1LY7fyA1RNfZ
eqdw+/oNBdZQk9d3ZhCId6BAcYgJD+PWHYEteXHM3tnJ4xpZ/R5s9sujZ+3ppcsF
O5aD2G5SSAtKc0hF1CBg/YesPi7vST4zPwB7tOeTuuufmsdpxMnTZpnk3YkvRBdp
FN9MW1hffNnWCV//q2C2R97WnJfNanmffIQ/xyFpy1yXNAZAZTMXuEbJV5PSjA8n
x7VPRKM8GN4N9WAU7qUGSOKYcrEkPB5ctuf314A9jOVsgZthfkPo/ABp2XOEJb14
oYPK5jYplyRU7pIBn30aphnSyg2osbo5PzQBt+QHhqESYdwMIjeNvx7tlVsHWXWN
yuqDy0yXEN8dkXbl7V8QJsqzQ1qFyzgT5+xDe2ecciUVRRf58EIS9Nc/Watbkh/Z
dCQhJYPKp9o8C6okZO8Uf0mdeSI2E7UsftMdf8fh/lCGwYMANkNv7Hj0J7cEi5zc
Y+KbK3LiZNPX00iPMq1tNwRWmOO+lAw2e+UO2uIH7Yr6oYv4eT3EIBQQ/ORMiaUl
5KXy01LfG1ldTiIaris12GsTUcsaGuZ/5oR3tj8DTumffANiDOjzc3LpPFONqb/Q
McO5iVP+cB3nomwqYeVTU0/41r6HIdAmT3hlx0J2Eb18UP7x3PzO7/77Pe1mMdSQ
lGxrxbuC8UGQWAEZ/r6fzhcaJRCo8QHUMVIMief5RnfKo35i6Su2U8GvzNFr5LBx
yPk/WVLjTJ/tI8hETsG13otpOdCXeylI9Z8LKKmJJ3lsyZt+DlGeUQiSJkCCF7h6
VgC0X8I7ujfX3RNCbD9G44CZPHfH+l5sGlpTT1EJkLx0pXo6fclup2Nmco6Ma0TZ
gwZ50BGp1ZprsxTmFQbOsfcD/nrhttNrhDW0nV6GAaPqYaXsvee5JWiU7Q/b5Pf2
n2vItNFRcyTYTAJem0dolQETDccHrjOsuxPTV/K9xkbw8F++4uumlPRyqdavC4WS
EuNyv3cxOm7gCCvG30ntC3jMm9WEE18yqPMNO9hDHGWIHb0A8mnRNYloPO5RBKq1
ILH36HRJ290OvJfx3BCEEmNV3Y08YlTdehtgWgEGx8Lpn3TJP9av136m4KJ4y9wT
Izt8X7P9q0FEurZLkf3m9f4VJcUWVdjzRUfIe/o6ujNeK5hG2XA2XYK6uvkXyitB
gTFNac9F95MkpBR0fVSmCg2K69Rgz6Umcn+335L6cok0LMN0iJffoAFE/Lo2HLSb
pAZIK2fIbXYgRNZT0/IObFc90n46wJLIuyQU5rILsv62cTKrZXZjWk9Iyti4hQfS
dSxdtIfSzQHj2GDj3bLTmCGIrzAIZ71PjoBc33px/A+TgfzV8phccWt+6w5cbfv7
t/KGenxVO0SZBO/9Cn2I34LGIUIpvOKakbu3smBVbBy8UBWFikJmznSdtPuotJF9
I7i8Om0BeqyD6jBH8EHW8pf60SycncPFtF8rkopPmT9OpAWX3/Af86wm2lRHTyKj
J3rRufGk9XzuudPaf7YcM3Rjmj+OsedZUI7T+EgBKBWY5FYhBQNVwTcpLyRDKa1q
2qqkRFQLgoLl+ugFGvJ+oRFaSRgXrZz62/ba4GsqRnP3NUSJQuLJfxuPsHcHogSU
/6U5gJeEOGEYkpRVTkquFZVNxYOEx7qX+UV0LL0agHBM1ryTv4F4hRLinTdwb1sK
cQhd+fgKGlvVga6RCasPC+zVUKMdUYiQZHZZllSDNnj9FNsSAI9Gp2JX4nCd1S+n
Frjo3y1TRkS4gXmyFeDdy8FZiEg2MiOv4j3izc1rJxO8xD0SmMHh2UEdHrj8uKmG
VU2xq6jwmzPKLSWsMlcuVk1UcFezDWRy/5jyjjlqn2mlY318O3JL2P/cAZeK+fYC
VIUG0erzC0sD1xzyA61y0wLfgJOWoIHt8LnwntFYW5xesmX42up5q0P8wL3BH1LZ
v6hhxLuwIeqU8aLT46mTP+OrPLq2ZpOyc3u177AFB4et6uJiJwQyExdO1udEuSyP
XVR+j6pxOoR/cd9uj0Esb9e+pzrlhVQcGsr741QL8i5oN2qS0tyPq4/xV7c8NARc
pNODpLjHiKL1JxLJv9PhqTbYxlROE36zZm2OettVlTczUptvtHIwISJsDwzKWTlq
kwsN3gRJo4VL4vtnZtldHqUvdeuJPnGvmL6/VBIkRdj08nN1vsSfehxBCu2WAOTV
XDAC3QBvtZppgCL6pNWxOvMpLpblwnROGbiN7WAbHlFx0wqMADT4b8JAqi7zI2Lu
VuzuxNoCYlvWRBT8tWhQKyYDqjaYkOn/8fCrNAarsgZCZpLqNr9O6V0IrJ+b5XjP
ZKlKC2CVyrZcxelZzWpvxgK+Fir1yyw4vPwO0YvWetxRN6tRLD54GV9uYAqWGxwp
dJQuGfieJIT0+yN6EEIeJxFd9NK6WRmexet+lxOeodS9JBu6NlqYmDczsdFbmH6T
iVLx7y77sxUo1klZhHrbDkS9J6gWXtdAGIOznHn562UU9MrkJFPecqd1t3FY+67l
1vB2D5qtPNFyhxXF9SS4LBIjZhppWbyZ5AcAv9LdZ8WNWjWm/Ag+rjUOkm4Nneb4
jZPVykS/oQ46C7yarre0AbetfYd6sI31G8D5gq7Uk15YLcMJThlSeBQVM7tvCZsi
VUbOGFbA2OEPYRMzSUHS2oHFR34B+y2XEYZ5U8a2gs6hyPaNhaUR+l93xkaFs6rl
sOq8H1BvgKyQ3vDLsOw1dN6BvpJoe/JZ72+MgrkucqOabIxBFcHlknsdPpYvlnp7
xTKRAmlv4ge/B+X/PQe6WomqTmtLlNdCDb0wgVzmO6/KZYELfuNA/fhc1fox+3ig
o2rrmHkbp/WB6Cs7rxyvdbc10w96+MZxvld8dXVn9OePSkwxtof4oYs5oIT7s0Yc
RUR/mhc9PvA3Iqd631Od2u+XkfgBupssOLS3LDhNyC8sdclZoV9ya0fs5+FKwMew
MzK9q/FgpRz6p0nm6ZCj3arnp7AG9sucx3PXd0NR6B5im5l+4lsePmend42WCH96
HsAhMS7iy2lpNPdusceDeKoc+qPrhEqzfkpGes8sioFTcPro0cu/JBhLtYfz6Sj7
46XuPzS9kiTh/rE3sDZmbMt0Z39RcDW5WBCORlhqhMurycpzkYOKr5B2GsOtc6vu
IVrOmCh3z9IhKlzZpVx5t4nPAaCa4fr9lSd2K6Lxsgfo/35CYPEqCd4O77B2MQbH
ZRXig4ZWVoVbBDNHsglseIqH28v25gBXXDyJPRoDQxJFSM8iR6mPAFRQoCtvB0Iu
7QDV1EUrJ13pD44dLXHdyAZJjmDiOWNdBTNpoiSppAOgA6LGaA1XnHrIZ2zoWwoj
TDTSP8rJOg8xc1pGOLnR/TwH/BmYeotRYKjfaThw779Oohd2SCRBYmkfl9+ov9US
+bHCX31aCKqTLpp3vE38viKD/rqliRAtvJpbcCacMlVeY3E2qnWqgC2VbU5eD2aL
d2eymzqPTAYvg5fE025Ajw9Pw5Tj29eOZ14DXH4ZKf+x4073U/7kuYjGvlOp4gvM
YdYHme5mCAsSeBQBl4i9SQusubbGV8FKpwFKCpR+KVbdN4sw8G2lkN4NdJKzWiPE
7Wq+HpA+xIhAFmIDjnoqU47oQ8S9mEGqS4V+ulEcnWtenI80r/u6giRBtHOdQr8O
F6GrE4A/B38sIAUr6W3eFM3AGYYj9F0bYIwtQuoa9fiS7sr3+jCN1UBXOaTZ4D2U
fb7I8SfcLoim1kIdPiFbk7SVvhT4rXjUci9SL7EwMBDfkypVNGOv6cw4lPBXZgIM
D8wlE7G3u6OLy8SjLaKVTBkoBaI7kFFPGPkDaa9bh1koKc0//a/1se2H/iQhIqNF
IFA4KOw9zSivDQ+ybXAEEi4dWzXEwu1J2FlayMiOwtv/hSzt5f8CeOJFOphd6BFu
ctX1iljFaM0U0wjPAoj8nN1XD2ISWWDx64sGhuwxIvqwItloYQe+o7tgNvR9k7/V
NznVrrZotgrTp3bU0dLonkFRRGrRQrQ43qmUcq7HsFJ97eYOuMVv7TUAIUdFQ3IS
9GFxpPhZ/tyVCR/Ir3qwFp5Tr1QZxiEzwa8tJTCASkZ8GwfuJ2tbRMbrGuCvhw75
QXpckNxGP9+G9V+4qyk7JkN4QTUz5UnOA42LTq11gUiBQHX9H8HmhdArZgmvzVLz
fFcQ/roENYhEpOhx/sKfXhfYC4kovn3XIb6P7NBjBeOk4MOPSNBkcOKfdxQ/TbzR
StK7X3Ix0SAUql1ITrbXBSWLSnd2IvQ3a7kFPod/YnAwb+wQmOC0s4fqCHne7YDl
57So9QTeRstSEZ3Ja6KZ47/UsarjRFeo6470fZTdjcgEd4W3lMbLE92b7FoSmyze
7DR2izHWUeaSL8/WGGfWbTE9balK8ksfAwFxfdCBbRmSzPa+B3BaRnJLTZY3hB5z
BvFx0NchRBtKEJXW43zRRJJyAMN6mZBu/Ac4ncaQPwYv/zKKfndbV74ObTrvdZyz
60TZuUdM2tZZuBOJXDpQmGuFYE1euQEv9pjLFZf91bhquqpfdxhkaWKOseGvSfoL
np3fiB8h/EvNraUXOZRYDRFhgGe1TX6VWvHJebp0yWg/lMpNJNyKfxKL5VqBoRcM
TxI9vhOqrH8CoEA+lGp+Dt3Fg2Fx4koyzX5EEgAmsBbjhhHlVsL9uO6T4EMWOKo4
AtWGuX19i0uN/FcgGpqdM5rQw6K95GTAGSlseQf+C4La+UNRL+r3WASse9XMQkfT
r30jps0Ffi6epY30c01OgKiL3RnUjL/u6oddHBVOIplpdlIbIQooR/jU7mKNriDC
2L9zEDPvsKANic7R1OGJUALtdvBmQRE+mf+3GSrW+xfcfPeMbW6VgJkotgavqudu
WZkvI/Jhz1edGt62rxfsTUbaYx0r/AswpMbgEfyw85SkOclMdz55w4DTSnGRBkvO
wI2LW0VhDBBIAFBi0qZozS5TZnkrrPR5HyRiY8pAZMMespx3qAJdL59IOE6H24LA
Z336uXa6j/xbPCab0G0bH/JI+ct8snjiSBQkiq9XFTYWfxfaJVzA8Xsfio7XjzQe
6Lbk5Cwe/9Y1VqlW0SeRYbFmWcQBw3ZvDtDjYbzPVd0d1eMBCeBN4PG3MC9PJfS9
56K3ouo0dcrqLlZJNdf+MbevzJJGkIKjEmDn0g9PiD2JJC/ya9MX1CeSAf9jhUQT
R/xLwwNKm2JxZKScnNqwVpIx5dEG5Y3uG768LUWSSjkDn2dRlhssUuoqxOCm3RG5
KVnxKn6ZfDHu3Ske/usUYj4vwpyGT0pNbenKCpQk9aqpLk23nAMJastGz8Scxf8m
zjcxAfo5F0rcpnQ11b3s0Ct/nDP9/HpG22mBGQ+HDDQmmMrSuw68jO7TNVfvyHHa
C+ABhE002hL0qS38eJSf8eXdj6cBSlxbB9zITTmrKOixEDxJpwHMkNYEJZqyLRyt
gFRO59f/4oIE2dImExAVLRzNNGyZm7M5CS+v2j1ZwI8I7yYlg5ETbSZ9xJB6rf4B
wY7esBL+ho4MDCXr7Z86EIc/bnD8+YY7cBjjV4Qch0OJ+Zy+3WuZApWEV7t907Cq
2FTGDqGDPesaakQbliG2LcpgFfKemLmTxK6zuZ4boTpjir45aXsgHTHBENPvb1qA
K20bwgt/V8d1BFXDfHcu2tU6EsXr5e7q5IZiRJKiS0Ys2Hz6IEXvGbSyBWGBtgz7
5ZBk0tKDBnUZaElP0F/xeIiX4Tj9qyZhhBhnrzJQ72/E6LCciSkDgplq38E6yZuL
c1Sl+xeShNxK1HnsSyLDciz7+6JPQVkfNn0vWdK1rB7/N74CLUdFPszBA3UhVKRm
dASso7sdmquK9qZrIQJ3AHWcZRk2kuFkeX+o783f8GD5qs8XC4prgWWDoKzNuJJn
vj5vM8dw1wG3lOnIzj0JAg9odeOiwSQD1V4n0NDz7X1x/yS1BS1ddq8hKxsznaCZ
mugCuviEyAdmBIBnAJslbjPj0fLXNIwjDP/8JwKH2CWKM9dfEnTSZCAUkt1S+G6d
h2jXgyBH+DgIAcgC6gB69qqyLHwAPVHXAMZlMQWlWGW2mhSqCfb5bxbgy6ocmi7Q
TcIGtqEbDwJvLRtkF9UWyhPhbCb/9RNSxrgwxKbwlMtbm/+saeNd4oKJA4F945PL
hrvpjkl1N+W7vuxLqvyJzfAGawYL0e3VK5upHGWsO9s7Hkvif0nFIbpBBG0mNSyQ
bUUCoRBcPQzFCJVhiJq5duCVqyE/IV9lYDZnHUKqq+ssakIiy0CY9aztT967icrv
a+Oo0i3gPmk6BxsvYBbgcfQs15Ek5Ibap3v1xKrVEaZZYZQ63fc1ciUnvmW2CohJ
Ao4/3vTxqzQiBWzPN5qa1HhQ/bQp927kDnUrHNW2pd8z9RUqrPoP4/PKqZOWtBIZ
V5UCj21NaXUgQAotQd2jQ0dfpvJy0Ba0YPz8DndMhcLU534OGHBgZGoO1QhmfmWW
0ASsoOU6PEobGLhRuxgbNOMeg+Z9w8QLixYWDNnG6c38j7lo1kLI48To50er1W5a
/qswbra2gsDDb3a7+5ib1cOIQqUAtsqgfXNCCoAYT37ZL+WwuQminq7nrdmjROMI
G+AvlYeBLouWcpey/9bBExmDQzRSSK6qrorcGQ0+fDNNzu74Fa+iXdIMvA2smM2G
uyJ4ZX3p+9mkF/3N9CztvbnVLYygQErOlH2ilZamaE8efZ47twnN7MW3Q8CH2w/X
QhflEU+nDCQjMDdQcWBqzYqX5DOvih7OPRyZ+YC55+1oZaktYpIS6A7wEdE4auYt
K9KgjYlgJtALU+K3VmQGCZ0kXMue7YCFOSOCoMtdnXk7Ew5ROz8qH7kJSNJKWz7E
dgH3nNDLixef9Ax7I+y45lZeNE7haPJlNNbIIkIphTRcS0Q2AlsWxcpDylgGfCy7
IJ1fAMSnvnPc2KriX3WnTLoqOhvkzlsQPf1t21xBrYdP8+sdB/RRiC/xCMecvam6
U5pn6L6LIvgskdSR5zIl9QMTXsMByl5bQSXFjE7oafZpc7VRHpERb79QK/bMfsFO
uOQ/6CihmY81KECPNsucUO481kVaXkCXISx84tKkgyW6AvnaHjtM44VtafxeuNwp
TwToZcwUzimoriAB7vZqLssiKLbqaYh9eLaBQYe4WbiH6K/E6MltYUXWJ/z/e7FQ
rO7KZayumEe1k2QtzbrUr532115VWDrOGhcGAUwSBFORJyE3OuVolmYlhWMKcmZP
rKI7cFxS07y+IYHoc08DCZVEnaN9tuH/MRLafWFjmX/r7NofAdTr3FYxRNIElVZL
q0m+vsYxnfJxheKE4LGhu/VmdB/RAQTZvMpjFh+Wjw9kT0dfGXotm16qYU9VYF7v
kAmY6oXDUCzRSsLEmfLFIorEpQdxcuULv45SD0NyV9f8bokXqagFCHKHGdXQML3s
WAofka/2N3h6ttsFF1f+QPFmTLylQLP3lcE8azEFYKzDsMfezX74Q1+/gPzVqThx
EkVmsXHDU6iLYrZ7TqarnqbV99TOAPnH6Wr3E2q4ZZIje3leVzdmnOUNYdrQkOmy
RpWG9HK0R/2pDHJg2LKJur1yKsBIDILahPPy7wLJevRzaXE7mQU7GwQh7ujeRcPD
cGYyVStozqmVL+Ou6g4fjdjQ7cCO+av4hMxyFhB8omp4ogUbn9tVEBZ9IMCIuqeE
xyPxTiCiYeMefhCQRyhFWXA+hG6CG1o3yHX1cfU8r3iO1gX/k9FpFEMGCBpQIUSW
FsPCAGsGMABCHdnOJdMAO3ptK2YGaHumTn+JqhXF2rh1sK+dXo34EAUUhWkjIKmG
hJ8xcQj9uyKwBmfXUo6rr/SzbSpiCkcIdIUm+GbWUDfodEBhaWbaU6mUcvhx/XCe
Z43Qal/TTzxL93jv8R9MiR8ZatG14FJ0aUMPQxKrqWXzsf1xov7bzybh1jeFEXxZ
bQHEubw1D4Ef3bIBzmb+2SfeRzQkHKF2buWkaCjIbzsw12NrOwRkhZvtN8tdjRLp
qAKoaG2TRVYBRJikw30RSZ7VKp2Sm24XYO2rVvnruzn4h5v4sS8QjAke4PyCyBCv
0+R8DC1AbNUzMgw7BEbAexEVlYF/G9slcQljO7aSm+v64+4r9pZJ5GMfc/SjMLE5
u0ewwZPJKYmkbQymMjqvwoABHIs8tI19U7MFhLvxIpfMYH7Wg+xM9Vu6kg355z5J
UPkGJXsJ6E+4+vD8PpTbrpLYDXc974Sb3a0wOuLHZFggB58Hi8XcfHSJMmVACr4x
hIggK5syJhuEHDAVw1e3uMMXRl3/itc7G3x7tnfH6DCG41GLTpnrDy+ZxexEKdtQ
oJUfWFUCbgqS9axBSBpxza+IHcxC9Ej+uAzTnkQI8DPYhQEspLcLAKqZxUd48Jlk
visMNL1FXeUzRXrKzXPSJPla8368R3TnSU5zoIIcfpto9isX1WVb30TpmzMYwXl3
INx0WCCzXV9gCthpjAFUMt19IUSMdyiJCGTZAPLVrotkGIkEnNOs7eG9RqfRhP2D
mSqe/4elkyrUFQlXz6aYYA0vuGHfjk+wUSKuX0BFDA3PjGEt5MnKTmTqIVzd7+pj
WrAl5eUeDHHtF9HN6cpDznM7RYeMVIcC6VDR6ft8AK58M+iVckGkBsdJZHx2FHAV
jv73qZ22c+Xh26jpHnG35Umh8YE7p2mX81P7WGVR9md2juBj0Hbh/mw1IAQZe6z8
fuAVvK1pEeWR23Nozl8Shnxpz6Qs9jGmvrdgc5peZs4Euoj5Zy9peMN6Ucqkp2I3
dOdYvmn0KiF2LOI6Ydhq3qgMR9ygFNpe6wAyqCtbtStJMYXSa855IOd4Hy2eA1nM
sKl+3yM30NHS3V/dI6/2IZBwni9FBDgMPAKdcP43mOt3e4pQFVNR6+EJg3oT5tUv
TEYzxuhTuAUStx5/ekvULMg0pF++kpdA/6lUhZjtZl2tqm2NqEjhEaitIFPnGG5m
aRNlKxoO6EdI6MRfxzT6bZT6nw+GI36OOoPnGQcJ80J2SCbaLci73L9AqdKVx/gT
FkjmL6oWOXKKils2a6ERsb7eoYAXFyfNur7AUmNyef5Kp2PlbsFDuFedt2fXaDJ9
vlyC2E8bpVu2ZUdRPnn8vdmq2TTyK41ONzkgixuzpZwxZWTKL6ytQ3kQ0pcfpUnn
FdS0AUDkwtAalXSOGPQ6P9VsQLhdgEA2h4iuY7ChSOjbnQXJBQj3rIi2wx4oxPjO
hhCdl9TYL7faRqfKrwwGN4gljCnYbEYyMHUpwWAhngQJWTX7fXB8g5yIOXZuMS81
gYyLZrRdlAGnrYrjD66zVdjHXovgq978JLX95r+sbUYoeyii3ei3ihqbkG7ZokdJ
2E6dZmvW+hD7+BDWBLchvPK6+XL4GPCdkqc6b4LsNsZqHRQiK/SOxYdTT3n7gFA+
QtSLq/al3+EcULC4IB4DJONKg6dOf+7IcrOYasFD6S8Iu3qxfK+pLj6rrXZmd77q
Yv0dqBwyH1sluZFV/SlvT6H1nCYkE/cvIRwoMJp8WwhX40xqhTCMjyGFqSw0T5/q
JBr0YEuQNX6dLzLG7YBAhJxU3p2JZebs/Jb3TiixFnvcldXnNRJGYwDkl31Graa+
Pyt2ynu4CKyFBmeCnHc0lVQeZuSWBnTwQ0smwA7XPXDGM3NToqKApHqTczM/+NIE
g8SUsoCF3OP0ZFYCTZgl2gJ9Q71P8YIPTQxyI2yrgD+QVennBIPwdN87hhTmCcqf
K58L6jAmr/24LLCK/xqA6LyEK4GSuZ1duzNQHIEI8pVBn9kR9W5+WM0fgcOJJwp5
l4Hz3s/PVBNSUClwkUVnRoet8BApMiFGSgmlNP3kGWVVzjYceueDypWcKG3VUZy6
llXALV3SbThpOOD07w56DoXWbQmDWHvNdCuazMuNZoTn4gCQA/N9qUx9/fAK09k5
VPfsot/MmjpMAmdUHMFZUXtdjLpkGMf/OvaNnZX4kxRdHjAWr8X8wymz87Jnuuix
qH6UCkjKpEJdheFxB46c9mP4A2Yue6Vm9poBDXvYK+1DhAa+RSqg9qJCYXvgwrlD
JnSbf2DL4D+jJUDDFqHKy7sbe0gj8vDADsi7LgKW/7MUWtGH4GzGFu0b7uIMlP7K
yBYXHhR9kltKhaS4QeTpq21d7VxmNs7ZrM0fb/N5K38x4tuKAE4JuGHecC+Z2h1F
fqoVcnPkbfS0J9iDazFBecO4TCyFyWw+ti7SOgJFCGvvTL1aQ7wrOMtj5bNUMLfK
spLe9f/0innSSoGHfPXtYpPyWFllzZkoytTxFKrZL6ZS68YIinACniw2pqF+TcQ7
ietWtuh5yLp4Ku/mjqVvWG/aCBeuVz4i7i+worrGrXzzOPrxtyZRgzBORt8geXVZ
QW6QnMC+iiDLC+212b18Vsp0m/tOyu/76aNYiH9/aw4kB4zDDsmNYLRx4slIXzrw
kc1gVUhnMkVMQfCyCKB5WERamH7QY+liDhokn6vhw2mPln/VvWsZ8FKvSKc3E5UL
RrKZRYTFJx4jxWMxMZ2cvkFip9IOAzPK14wwoDBWth8LyJhRvzPgiZ98Rf2vE1Rg
bfhdWX0/k+KYyLYIUjEIXiZo7W35FyYw+W7irer7w0j53nPl/UUQ1v7jpCQIGrz9
Dh+gFDmXSwXspGg3L00kfdF7SlTsacpQOgvKiYCLEgb1jTwA4ntpwGDlz86raaFG
sj02eEMSCXPm3MAAGmZdq4QgT6GKAqdLrlx7zZwrUGBiwOfP813Z0BmRzyc5kkjK
jIINzht4TVn0PoTUcDpVsrXZginPDK/k+dfxIS5LC49mPf6auKTqMEjanuwha/RQ
7grDlKA8f+RZD/lTQPrdt8ULe+cHK16In6VH26BrB0k3UZvtQsJZiLpF7rQQU3Bm
uJgpdpKQEobzklwhr1+PaDPN4GUeDi/rjisS9trSWEZH3Ig5jaoUNmTqZnQXQdbl
QQOSYPSCsL3uJSil9o6oTbJUkZpnLiLYrat+AEhuICIYyMtnzwqrzEbX0S35Oeqp
oH4lT9Y1bV+6+CUJFNMXwhZZB3bof9DmJA7Dnsad26DfJ/6in0ElKy0jx1gbQSzj
bBz5HPO5GRLjRUASRXIUuXdhKuOLosffXroTudXsz9OfzGb3sAjYefLL+4C09zkc
zAIyeq+d90MnTgcmzaOOYQAXNeCpB2GP+0hZj+DZNkt0nZMcmK65w0F8k6xl2vB1
5vSu4RtU6xE5v1XDTNsXfp++jTpHF6+5CPOGWFa4vfkq79ZsiB4ukSahFk1+FqA7
UOPZLdJNZ2MBkIl2KgbfVX+qeca+4dxdytpwcAWvcq+y1wBW2zR1waeD/gpMRIZm
KFLbKsTWoaupXMX6kqQpMPth1T5HOTpeqAXqwNkmsB6ABk/iO1OttCQsy6l/xZ9D
8l09qZwbHNAQCYMZYlb6SZibnPLuNIZrcZY5cynY3a/n4YdepsWmNP0rI5DmajTj
P3In0CLayewiiS2QLzuPsq062b5DTq0re3yqta2/ctF9jk5qOSkAhCO91HNkfstN
KfHKJECJhVpTIcLvl8pm2ES2PzNhtWBM3i+ehqvUK1iEWBxDZK3sXXwxBSjCImhD
2j7iZnVwX8VLT8BQ3Xz8j2wiio46Hha84plzEpOBQCXPTX7jcnUZdCjsw6mk2Cup
dDOsld3FY0NDOVWjFr86sbI0PzYTLyng8QGuhJB4wed6fMqaggXfWCIydJCgxIPq
RvEHcYquHjMQebBZFJRq1K8czd/Ek5acO8GJ4bgdEo99TIjenLXX9KE5FYpu5TTg
5yNYyS9Fs63DJtDOuyV+04mr5qQcPhSLGb5soW8Ib15wjqI6SpP4gN/c+VWYsB/V
irUBDBJFm61zsuiNtTUgCXZYE+HQavnApo/ae+gXRxpKBKfYpKkNoFphgNJVGfgJ
n17MR7dmI+EpfF2zJAhljiKMaQMEMhNEjGiggPeJxi+XZDAG0uFyA6wxlk0j3E0W
8zKyWxOwrb4b/w/JHfgooeeErKw/O1SlXfipa6HItb0sNeHDP3iafg7XOol4yRjm
5HqCoDDQR/KOvmWd4ZZmTAitRRozslS4vXS8Sv2HST5r0vd8TZSByR6QdYiUeheJ
RatCiluV4rgFHd1G/KyO1JpoTLcua8uIp1ilS3REfHX2Qe5hY/e1n0BzZ60UqEIY
uxS0N7i0UFVzDNiC9a/thHowEFso+S8sOYvDSnaE14C7D2qlDYh1QV4960TkDgvq
2Luj8eeVWxYJ3903cFcKSQhrm5I7kxt0iIHZptf1uQ/76BvCC/qTgfjagQMLqYFP
Mi8WB33tPKNbRsNBArICNLE407C3rGpEbLZ5K2uo2oYI6C3gNbv0nPeK+9aNK9hg
v51CVto56KRAFIgVidxxg6mwLOV5zIg8yyXRwNkVbjQk94+nnI+EkTcdLmeaAmYF
XuwK4jg87zofLEZzCF9WA2j/P7b/fHmBINLysZTljCsbg8C65yADPJnLLC7YBVby
0QOIwb6gx80t/FVxEUtda/flYrziRKFwuGiCbH8em97Lg8yLU9Lc6kGP2RV/HUmv
YimJ5i6okEasdInuT2FscJoKluwqZF9s9IwlmYeGE/KdAmZYq4UfqKNC/gocmbbI
iFbSpbaEne+n0sqnN2Qm/zWHCS1RL+fVBxWE44fiIpBWSUTLkeISq5CnQhZmAwfX
DCl8aPzlzjCi+MAf8FO2mcXCFrwO7AxKdZrP5g3G8Dmw5TLIGD5ehF1oTgtItatt
Ety3Kt+yTAsdg0MmUjVlsJvp74W2YwcnhBGgbzuYHw4tLUMC4trVUtZrCtR6Qewh
6cCSwj54LVx5XKjo77on9mOLvraGQ8uOekCLkXCCL/8zeIViYMWRUIZQy/5vEGuf
2IqDgq0Z86e6Q73iKH9ZciL+qBpq6lSbPXgKa8wK74OuUnaoRNlB0NxsNHfS1mRL
U29fzO/VaKQV/6aDDfx7fBimdOTM0EWP7BT24NoLnezMq8gX2JwvIeUJhtwml90A
csY5xid9ZBYFTsFSqB/333n6jVZBaYU0IdghnR2Pkm4PB85HxVMtAbKqDqGK/Pl4
tcQJrj3vaVVzMWx5wqGTHAcXmjbggDLTFDF47crLfB44y1ugqtLCutMQSjyZKJGr
ga3I/JQFfsMGT218BVmdRnzYxvbA70155I94end/2IcpPkpurM7TARRF7L/JwFiM
+8AgBZGi0emBLSRjIGyywvNoCSFRgBcoOfPObLdsANSp1J2y0ifIZ12UZ8PgrwnA
ZYbR1MtEeTGtRO3MfGK0bPSA96NH1PWgMTl47f5YJSkiVNmGWG+uhk3e/oaXN8aQ
9U4trjyIOP1iEqagX8rEGV1uDYH6IpgIGepnHsZh+SSXe/977dLEgsIOm4OKBHuM
GkEA65Qsyn+cOdzpIVki1aHIv62QhdwJLB0HrWQJia8b0IivD3POiqG7A3i1PRFD
S+NwgpIlWf/OBOFzDbFf0cZJUCPnjx0Tn1Eqn+SKC58Y2IUaZ8vV4hKy2ZKBNu/Z
NPXGP9ieAAladi1tkXpsH9yOBeBTMkiB9yd7bGJSIBR/TQG538eS3u1FnCdLKuZc
VqzBquOA+jmtf3SkPNt+El/tWBh3hvhkHTG6OWfxKPU/JXc2RX9Guk2Iz9K8BUtx
pAIqddLbBdRJqPBRsrb2Vjjn1EsYZ6+i0JQQFUjWQ6dkqPI+XS8eXEqS3fcrUK5+
MYfUiYS6yxdLIJ9ItyWCd99yn9+mB6219EtTGfGfGWpwlv1/JtSlsLhmxGzipuCH
tM/3M74/cBZovdc3K22q8GvQYbBOLN+fz2XlOIs3E3CktJ4iHbMRctMKRKTL+0Pt
+JFTwizg2NraQe1L27+ttJ9AU01lPMKJ+sHf1btOq1pTgjuCQa2t5dkYpcn30oYf
HTCbwEEbVe6WXg3OKtY9I2IcLMOVr/N2nlKOupm+Ip0fAsbUit3qxaThEhsarZFf
13lYNppL+nyIdExn9BS4vhfojTZ8sksZdXuZWcN7zzc8kQaqrKCe4MOYHUs8YBZG
YHpRwWbgUgGsqcCjNBLGJUZtUsVNBC5hre66o/Axi4xq+JRzwjUIVStPAWYyApJL
fq3AZpKbRu18IgnhO5sRN2Qi3H4JsqdjXh1H96b/Cut3rpwjv5f0cOPCV+1hwFNj
6BDnAufCmAV5s3ManwhCJ8JMAkoi5erqOrrlH6ixc+U4cj9gVqXVIYutAVtTm6UX
i8gqp/GoiQAKbz6bt7bwAE9P39eyjER5IWv5XqB5/HSqXAIFE8repz60c9uTbQLQ
Ax875X0xgeeRwU752PmFVHcv2H2nj6shhptJ0f7p+e3pHYiU61L4xoOb9LuPLH3w
nG+lYc+AASBuyMaeBtGLhpkdVu6LkNCuBROQttcKjwYzduJmS9BaPlza/X05E23E
FB6aski9Olv9JN6KdSUsoTsAxhQK6uq++VriquuWqWTNHn00ah+CeHFoGNCPT9Vh
afsY/1DI5EI7wqBM10tr9ZRcE2JcJ+7gdCf9rczl0JQ/Jp1n6fOgEsSELo2THUXt
0X9UEAIm+TcgFzibxHsCim4bhT3wxiN1NfUBa331tRJzmy/7CSY2vGroq3rI/pne
Gbd6qAnC+sMLntm9I+3yZYkxB+7cvAeviLUPpwLSGOYDct0YVGhjMsRGKRiG1QGE
AWmJDmEm0HNdgOWRhwm9tETvU0zZJtytwJWE6Liz6fs4Fdr8t8+1pBF4nJgn9i2s
q2QlMpUnCduNDvru6zdGr7xQUfYxQOpSerJ4U46TGDHHK8KaGxmVg6ajOraIwf1E
i6mZM/xVhe+mNc3KLmXPYpknIScB2zUb4vkkE5jvF+zoXIgV6DS4dnpQijR1Gum9
P5EJ5kCn09LbB4XkOBBjGti9nIIHGzGKpj9szKRkqNfQOjpQDStrzHJpOjqfdNZS
hHnXXjaBgvUKLGbNGBLQxX6ofB7jFqmVzjk+gfepWEq5xEKxmAXSmRJaoR8rYZsD
wEyZvxUG5TKG6e5C3t8xYIzPNDBToj9ob3pwc7trobKtF5Og7MlxeJOnDoNpsZA5
Y4S3Q9WQU1Y0e8kjoGaFEvvK7CPjlcH5VbiAxVkPpjEzNeuzGw4KJKWmxDBv7SKO
1LhKA52UBDuK/vGEC24tqqkIi4C7FDl3M4s9UcDnOINHjmMnRFHz1EJtJRoL9lHA
gE7yLZJdkTDEs/W4YsMRban5R1TpiI0zvVXEUZsYgZmqpL03BAElnJf4XYsdNfpY
Zd/1obpsVQgNQ4cv96oXxK3xHffI/PGCRjMcEFa4m24e2IZYUFycKRH3K/zo9bLM
un9ZX9g9EkZ3sU05Ur087vtDqjQH+sUOs2c37/FiiyYMqDm4NuoE8vX7pYLcekEX
dkRxqXSMAFQleC7912/jFP4pjeiiyeeLuvlnUK7bQN4WKUUMVCzZWBNO7CSslJg/
UaVx5fBC/jKsvAtWzJbe8VKuMnKubVbAWFRJ7HZIgF3cwMeAqZBRXAKncSegLYdZ
2Oyw9FllYdMpet02bFcfqxQkhS/wutGLhL8+hS8PE2vmNb1bOxDm9gb8D6sjHdvJ
acbYkIOtENELFuk2toCfGGwml6hOslm29Xdph4ChXLlAr8j2PK+LtNsnlHVjUdDX
+5MXTLXWZvPKY0x7vcZ+NLnijEkHWDkEG++PHiYQv3BjbwTntLcq8LPfzWlucXwH
3cFQ8d9K+x3pVQMSLhmYh3HrXX0nEUsSLqI7PKbyRqVFvQtdui8yXGC1DUF4xF1T
evfHyZeqdgS/3HrB5+R7ZFKN2aBd8cJL5mDhZ9j3WhRx0Us41OwXj+mPscLny74Z
BUKZ6+TNRidZM+R7zfqasgqiL/wGXcZKTm1tDm1Ztf2LGQmpLAtXiMwAXPf2KN1e
eSKh1dWsTxm+F2IGeQSXNLdAIev8cd9DuYkd82LbjZ2Fjl+wypADh5sBHXWVQQaW
MxGolu1mGJeQ9vBILF7yY/lsVOLxinqLm9oc25m89VXdFBteH6CWgyDIzSrLRGEt
xyeJ4O/69jvvB79u0NdDsTBs/AqreLFgtn/+1Lhth5HKp1vU8+674CfD6LcSz2Dh
+x8Q2QPcZTl+xv6AEEkBO8kJ5tRkGXNFBrxH4juyH96L9SsAIi8ceT+nq5wLxDOt
2IEzDGMSunH+0duFW30kFEsiyXIxBBZh5mTKJemMBZd5KVCYfuTupMWg5HgpdmIi
ycjljnpjZ6khSDodc/sxo1Bq26po7dNVQz9qk+aivDaq1FnPNbXKFAqFnHaOr60v
2Y2DnvrPgg+WF2kOH1rKr7IEMq+VoeetIKedj9WEioVchVR0Z1qhuceZ6z7wgexg
W5RijAxJquKcuLvEolRQL43jRyRWMTQL4f5XuMxSvSM7bIFCgreJUlpha0VGpCIU
dBkHhGr4H86GGjGRPNqtHGeNrEthfDlProQJCTf4Lmtay2ng1GGb0vTuxdCO+Ii0
b6QKCx0ovvxjiVGDltZXQTOGcM2V94KGmNRKi3OuW1MaN8wSywCPEf1t8YsRNcbB
CeGBXTHV2v76XjHCBR7dnl7Mi2PKOwZgqwZa07QpvX/MA8RS1jHyukz/BI/7Myn5
pGIt/ZHDwaoIDpxvAeWAhxmYz8E82qa6vRKJlxq5C39saXnO2H/FTj9Qzwva/kZS
Q3NHKnPKrfKhNYAPFrkHwVZ4Xr8KnnW2RmBpO7wmbScBtyYA3BywtMKYQPCxZCPc
v6hRUh0NTO6e/TASHgp/oaH3ajgKQR4G4wPhGorURUUKIiurp8edASX6x4ushrkM
0edqlh3EDlbndva5svKqJdSurDUqKlBtvWx4uauIbZty2aqihoEJt6tYsNoRDiUI
i8ZLDsV17R8luET8DsHtrqJusaxqqiKW5RYS04NAINgCbrTtxgnxCu0K5L7L7nuc
JW5+HJvKbSv7zwybGYnqWhe9sFOvrCqhLNN3yhnqtCJuyHtOm499MXK6CkJe1fO3
TS4DBWm+n0gxfQxIS3dC82O5P7qSxowbs5/3+BvXcmQtaikVRH4ziFckVUeradlf
p7RbFOvsSHes7JQZFWVjOtX/exth9xrum4V6dey0vICsSx5iXf/SAwCEAwdgmMKL
xygUTiVmDZEs+KtBp9s9CpjsZDRLAFadyiaHe522alUKfAiyXaQfkEFK/BfPF+Is
Xb3aSIKHiqXwJ/kvXrvkxdFD2ZtC2DiP4iPCVzvCdmcnNtZ7bQrejgmMKNaHH/lv
FGvN/+lPZCW7qukkhlIAdKI2gSbbxbH7UVEM3weZ+8l9jhlYHtApES3DaGxGoG2f
z9ITvKkR6pQ5jTlNQFO5+WqU9icysqWvdC/Gdfyn32JMIcYIEdhrbvzIR4FOTHMf
VyD3GQw5JnyZ+zlV3bXNuDdsTRmRNWVNIBLvR/+CmwaSU13BGnZe3R9bfIqqyhGz
9oWQ+BGoVm5Ohvj6rDcfirQN5eTMUyt8m4bCkjyI25Y21TDYfb9kb00/CcBJRagk
xz/CLABdPSb8lOvaM3xH/6B4mKtxp48MGV3DID4kZUcbFL4fIrKT8Z6vtWWMqJiU
GhB76+6yswwPjEGzGDy6E3WJDEGKnw7kdcv4bvGr9EjKEVLuyGuP+vAImVKNeKDz
HkMl7flD/TyJmiNjQvzIY5E88vnUMtriyPTYzOERyPU8HeRqHqnQuzcQxSv1OlPq
NGhL9fvLwZVfmIy+BGysMq/9vvONY+yfpOjicTLv/095u+HPkq8yyDLHckpBYlfb
myFJ2BC9spQ2x1fV8zblf58URtw5ustkedj55XEYdRlisNJpu+OsBGSEl+JT/VLd
lxRjFgyDFcmuq5O5Zk8KlQfK58DiAygKqdxJNt74nwOD59YpTE77Lg5yfpPmBgeF
YTGYeWBSxOlzN9Lvk+EUCVZd7Tp/c6etkQM+9opuB0HBMHopRt5itl5iWERme3C+
b4DI7J+RZx97oW4H4mWQ6x8HDByE7nbH1n5Cfg6PcD6k8APCLUhohWNR91/9Mdow
d5axZ/ZC7BTjzOAwpCmOs+dCVOq0n+pJiKcZHtAcO94pw2TSEP2A3vCHgMeeEmF8
MW3EjtqmlDNg5HjGgDS4jR6t/x26GWgzqwr6GO2ukqWhRMgZxyhj4juPKy3uz8et
1aCztK9qxt2b9jqeCBbLVxJT1bEQR8131nmBSKynFGJT8j7xMPEehts5r8GEzpkE
XhHE5jvqctbT8rooFmqqoaypqr25HfmdjPiWyXC7qfU4KZHPVte0GQ+kkYAe8ChO
VFATlAsdrH0ARLaDgRMTouJcff3I1l5Nipzm+HnbNajlKJV5tseSQPpYqOrqPvvw
kT0aVMochKv7AGFHELEPbexqImM5JQLUf0mv7M9Q/WgFjrzTRWa+Il4jccV6sM+t
GR9eN+mnaegXhLROn+liuxj4f87pij6FAYL7tKGOCCSrfuF7iLRm6Wl4/2lKAvfs
bB3X4drU5lkKEtBuwes6jlbjaUUZIH3wg7jvAqXceRdO3a8C2o7XJ79C1dSj6D6b
G4KX2Z2s6mAAuqeOAMGx9mV90HsJryMQPXPC4lx4RXGwxQT6+ol5lYZwQdN8tOTA
0GmjqieK9zDCaxaKt8jk1bBDl+tB6KdjHpzznrfzgOJkFDFUxh45U15wM1yxPAIh
GrvtYffQUCUGRihYwhMawXKffY55CW2Zb5AQqyiAFjHpRbqWw9Hi8shaBPvIFW+Q
HsxFGScUrUDk70NOwabGXx+fPnKFDgwyC2gBM0bVA8wTE4VbLQKmMmyfU8hzjUvZ
w5tpeuuU+uLq/y5jKYnxP5LJoVvyyFHa177GEJsvwGhUUKSVHYTFwTfgnxRywOWE
73mSEvtPFqoL2B+NbY/w5HxYM4XruhfTBXIe0nod1X5o/GEGTC4F6cH+H+Kkot1H
C+u4BzYMtF3v2vVG/+/X0oUhUyEyln5EwchcALw0kBBQllYBTFfukvdIaciFjO0O
zd3hfwbc27MdtGbFwIuNThAExQP5b78AoWkb46IsvY7hLHhfoidlqlITwmKBllkX
m5amuCnp8RX72SQ/BG7l4GzDuK2awBT0ldVMqVhd51OzVtt1icHXaBXlB60avndf
PWet5CA9MQdh9mKlWo5BKKYfSB37JKnQidAy/oi9KMTI0qnVlV3sCQN1E9aUaN36
PIKBKK6XkjbmLYpU5TBoO+PNPWvUI7wPkfDN/XTVzJhTMb7om4tGY23NdNusQ8Nc
zb2/redYFBHw+hICTYyw5voCw5Yy5sosUNA7c579l+VZkhrsKXt3xTCox1lkqhd9
JbSJhAyV5lIiQc0m80kLyWDsMIpALbYp98qjtZBTBXrdUokgdoXFkpQE/u5v8tLn
Q111SZOCBFuAb1P/1bLYra8AZVvCdGP/QlLc612HCEM2Bjf80NeJkJn7c615TVDB
P5Ka2YEZDJGP/vxOBslhz2C+bRF+b7L1XU+ppFSYfdVWS6MTwhta3xN6yBZJnil9
jvDXlb5zX6vUvyrfSVTlKnvIJmJteBW9/3Fwdwz4XWo4XdQ1ZjFI8LOwidlrsxeT
ypxaia0Ink75D/tjmi/EXqOVzQoBy6x27IsDb2Ylq5numNTALc4MRjvY7Nk2mMBG
Qd0tDoQYZe5ZJsXYNFWhyAElPDp5zezMd4eFcWCnyVMYe+r4SxqZP0UVAwiNwLI5
c0VViz89RCBLCwlCNy3AJnpvFMxSKmhyJn1i8NM6HN93lZB820AoMgJOnkOs7zsv
F+PNzrZVl0exeM+eY+V9An9MviZF6ezlli8B+5flZjH7dUa11kSIb5p8Q8nqp1dc
ZRluBsMnRIQRWaL1ON5ny38zOurvQKYkQv4nBz923Srczu2lfrcX6SCpb+v4OkLq
rxYQyDkthqXJ9Vh6GJItM7UZxs4lFMQfXe8k80Q9TbmT8hEOYvbCt+/m2tIgpRrw
JfiL5/7WjNks/5kPdkHx7tBWm8JhlO4m2PBYyUUuHCdf/QCy9Luds5ZMrKNOfZ4+
uD/qu4MS7UIIkPK9hSg2D28UBipMaqu/fWXr5TOprzuU54WUue+wxZJX4bLItgPG
vtH6tk3diEn53kTwwmlabCn4qt+VV1ze32AqwFKNjRr4FzCxkijzuG/DdiGBwdes
1Oy4vtx2QHhSFH5/xYSftYTzUoZadac1WYA4u2VVzGCYYZQnoDtDy8jPijhtwrJu
Yn/N0kplEZrHDnLwMJJZTZK+BZkJDIUsoe1mKOAYShQtTlLaT8BnnXfhOh6t8iTX
sCQ2znPRLz9MnKgJM7YMMSXIGNb+XixwNNmW7Cy8eR5ZwKitArb1vxm10FmqjnGW
zCmuhfWzjoIpd+hYrt4+I9VwLHBKoF4UXidjTDFfnzg6xJyonlEOKKWAGvgkOP+3
4la70Fo69MY7HyHy3VSFyo31Wh726BbhqZMv4z+IrFoRpbtqBX69h7UE4uOIwMS8
a90LKY+xd3Si+QiLCH/r1uZhkw353ySgO2RJkgmyhRCH4j/ZsHeHbkhM2Eg7jSd8
iqfZDbpIEwowxc8D+IcSLtOUwKGX/DcMTw0v1xyypwGrDGxKBAsay+Wi7+C9E9O0
OvAMwDdksE4euIp4JRNHcooyyL4CLvpz7JXSYFrfwU5SA0eo06vpjhtNMrAnEnq2
PxeJ30XH7d1zZ7we5NaG4yMc3DauNl4Urdq5GqRZXE6KlE5rD7GBWdlBc+73P8mP
JRAdlTimmsQrjZN5wBicnbwEEPOlutN/qBFTJaZk2ywZKsVrc+gQhXE67o8MaUji
ns/W8qo7i98du06rKqIMGrUz1S00tyHNTCEsSGT0iDPQuwxCAATxNjyOzW99KsrN
mVmJbQTLx/HblfG+RqCf4JDT1NCz6t/uY5AtEcBmXm1XKx8cZfq+5OemLC6+oOer
p2TSqAxXz+T9SvvEzitOIYElnEubq0uoshLVqHcPSN93lDssJDSVyF60jNwD55uk
3YJIG2ZI1DNCrbVwR2xsYsKHgGgE/3sbqVmFLU9o83AL0l91TAWyuzvaKe2ANhAk
LJJzfwLaXazJx7PQILB7BeqFNgaJSkQyNJdKUhMbNgqnoVBYNf5SLEf4s++16beO
tSn/5rvTrC9SxvLy9YEzw9BVhSU+t54V0jUkJT749BbQ99Ja3+MJNdnDZ3LNITEH
kISPDSZn0mnIDrjVWm8VGvcbddeYhBXVw27PinKtSPejC/Br64O6tdwp+P18EuIt
/bt1eP5HE5ao2HEb2DEuqJMp1QzQLPYF2N0kLJYosy78LyGn6rOU6X4gsuwjnpua
3FaYUo4T8MZzqLBBwz75C9JaqxMF86rDXTDO1/82woQR4w3EYawzRiBonis247pV
rbYEExvoqTAovabmZy74PqPtOdJxJIrwCtxaaJlGL68RvkooyjKXriNC0tvuC49/
L3lvoYwv1sZm4Mx+tPv8xRo4S0uV4r7lRSnwNkjAAYrPo9/HH3xqYbkujWhsZUqZ
6GtJi0gHUJSCYBJrK9xJbtvjddTVc3O3eyJFHCDDNpnefRIdQ/N5Yrjq+q4+MR6Y
YHhJ+mX9tgLkLKa2NHM3E0NmB1Q8Tfwzj96NEmuYnzBC5QBqwEtcJQ+dZE1udTXQ
jiJqay5oYQxiHT3x8AVTur7t9nWnE8D1aM5NuBvfaqtv0yCo6XV1rIfOITpyEJ9c
YBd19/zUD0Zt5IJwqxINGX9KKh2/Ru+pXudZvv696JDgzufuXzpKB+22/8Rnsx/b
L1Tdj53pfYfnNQp6EycUoQvyvzC4+QwsrGPXoV+w1wPSHOlhylr/Mp7ln5LY+AD1
/DyFILviNCXjLUldfoyDNpQKF+tOrrBDie+8jzBuHERF8tQi6xvJGp+CWH022P6C
9XF3EXeArL+h7gAdBlsivg+ncDioEBhm+X9POYl/A/1/E+4F/rDorpNNHthmVGhD
CbuqA4oTxC6nY18ICpEWUa8XCB9LiDtAzNVAlH4UiM1kNZ+tCJQFVU+ykBDnbYfu
omdo/lDqd/VYuU9qWuoL5I4F+w0TOPJ3tsBbKBQVmNMoiij4tm4h8m3219wIxMjN
Zoi3F8j3JZ1MzIB28wLR748mduDaaWAE7kRxk6WjpwD5mHI1P4EWjZMIR3p/LI00
lpferfFGMPdJZ1seK3NO8kfCN9a2nFjZp9W1hgMZ2yjBwrn1jHDPZKMrCjNvbDfZ
kmbZn/w2PgASK/s/GPNOH4vDAw+y19ggFuoJ7MkGPKEj5MljZosI6X4CxuKnR+JP
ZSo27bAUPGiqrrnGRMY6dCr5fR15tzEzSQ4dUS+4WdOKZYL1PvRb3Z79T8Twat3R
qazJNFKCyl+Se7WH8YAMFLLILIpd1v1O/3jcZyWYlOjVMyYOpgNYkMBYwuTITfTh
q4+YM2MCNjm2LRNrfmhQskLfraOOOI/jn2D69HbGkqAvw3jNzDSG+3WPAdmqLhtg
VgkG09hWLh55lOQQqdvkwdBco+BgwjJb527l4nAh/vxw8EkYYRqY3R26OpMpCkvf
j/6CqsB0L9vCqjTA1mI+kXpcDKWMzp9zRSsnMVF5iBK/EGiQItoF4ai3moS+/jQn
nfe6Pq4xFW4Subb7/vP+hYZdOlAnHTfvuJbYHG9rWwKvoDG4noUivjHL2szT4vpw
YjwUMbG5AtZxItCG5YxdMN9j5X1DnAfzhQyj/pv8dOWi7CC0YVhG/2iVkuBcfyWm
zwIvvuNsJg/ATa4jNUroZSWMVZsZM9QvsMNt3NwqLR2Z0T/FTWMRV4Y3uyV88YVW
DttIe2+BAUvptDsyW93s10TG9mooI/i1JMRISfDvGBX3AFEXqVCccUFl2RpJggq9
VaIVWU0tBACDb+Q4BAxZXpko0iCLZW1beBimqpsnlwVDFMG5hkGPOFsdpvSjKU+a
HN15a9XFMQ0Fb3xRwOtai0gtJF9c0awxqhiw3A0uOpmuetcfI4u+un91Uy3PtFC9
68fFD2gKBYQeMOcOt2ZF5tnW1dWJe0UOvOOpnfiSTE8I1Aw8uq7k8DQcEeF4HVFH
QYILjmCAsZjVwxXjnw83s5NQUrnhIpO+wbUKVsdBjwPe43iv4BMXr76k5HL0L7q8
+g193jMOW0vnq0mJ3sel1o1isZKvPcIWQAljtkyqB3O7UO4YyZYBv8Bq9Nx9Gm1z
difRuODGR1PEkPJYSWRCzv+dodYvSaCHQa2EyXBHXe6+nL9FfubZwYrl8BqLVTTk
V6oxwsr8oojALnSmUdyvCNHTf0avZ16Ye/ZkkHklKdNH0fwuLbLJf2HwkpXBXqYl
RACto9GwLRFvtsWRBNh4pDDixr9PPQ28Y5ulk7o3xZMXteWMHScg7tkMjv+Lsmq5
T8NSdaz5tv1HQRlpCOKpKhP81npy1SWsJ3qSRDPGsg8lVSSnW8cro9Z3D23EFeFU
mY6annyLCj+y6vfoVsTgfPnBn0tE5S7qoxBYKsFW1N3JFnFgSrn9sWmY2XBdywe1
K0mpcrjHOdHp6wH7OwOBCF0/F136nT+1+4CXteFFesAeuksFoje+8Xf88h6WbqPq
AqvyRzs/ABJ52XcbO9fxYY/OGpTYRNg00ynM8FtLRLXOoMya0g35kX1B64k5NVmq
z/J8F4IlRGIhPxNuvBYkN1DR4cVO5Ylyz7B7QP8KVtZN3BlfjzXt9/99rn5vIbUp
e2adVD8yNlDB/trFdnbbJB1gOF6pd47HWKNyWzLhHaV9deHOUiRaYuG/FYeKqs5w
325ks2iFS1xLrOfcc7+M3giogb5evk0YXCIuCOVVJIwPUz2FlwP9lb7aqx/fcGrM
TbXVVg0Vi5eiBI0vDGCjYZMYMj0mFpGbM4LKs8mC2N9XrbetQ3GJYgIaGkO/EIIE
+JN3oD5V45fCJ+hM9cfi68BDCeVbR1ft/HQGlAjM5U93TJryrvcqSHSFWH6uQ3VZ
l3ONFTlEzzFFG+BIUnbwR4VSR/wlgko3LBq4wgYjn407oWuY6ociEmWp3NJM6Cs0
pQJL6rcrEcN5bafqPcV/ulx3pLqL3Td3BmKNRsvlnSKId6WX6vz5DGezOP5LjSxr
UtOa6FVFxMbsK6Om0fHusxiBP02l+erv78Z306qyRt7dLALjtEBaZjm2bWTeRasn
LOAzQ+22cFgNvl+fsy0z3qGaXX/H4ME4IAnFHEcqEyKp/jdnHrU3LO1TzZFTgtRZ
O33rqlX104DSKsf2K21woCjReBK1phcO2Zi0sB1o5Q4qqaaQu1QDxZB5UWSwIjmc
UgXVcf+1ACG86e25op620P7yvwtVuabVScjsw0oHxuFnD0y9Po3bCVghHBOa0LPT
bKxKiBKEXLpX13NYGH2KXcyl6SXBMqmdf1XizyTiDdAReXaLsn9fUYS7LiMJEVM9
Cu1gZ3FIVGE9eDx2BKPadhzErISXIzsaLTEdJgYveWVak5bp7mLAgqNFfcYiuFdV
o5yv1u3DRXX5rE2kssFe74lG4HFwOrMHh8I/dp9CxXoQ4xsCSYnTxGkJB6fY+XMP
p18HqW7Hllwx50MZWQYZdehpiV+eYIMuNe6zqZNVLacnpCYUR59euaW0cLH9/3+T
6H/MnRV4vatZjDCmmh/4u2THsxI3+VohrHegeOsofwD/Yg+Heh3qO01c1fyuYCpU
OJ+1BVK57Fj3KN3ADGS82ecRKQEhk+8Tnyac3rIiU6LYnR+3YQ6td8T/5S//c8+c
pPU8u208GeojM6nmH8zUJ5o6jDeb8lTge6UyqFIpcSq6CYG1xMYankfpDYPgdrdC
tBy7hgVeKcCGSA+gnmHMJWlV7aGpg2QZ3ixLuchvZ25IEo7ZEFnHwfoZDSgux+ry
ynkcGNihoBonHCmwYDZ/Gc+8ofr5K18ed0jYOW5JLMiieptZUjXloySpDc8LcVYK
TgN27UKNjw+VA6e9klITMEjXeCZ3I5DA3VjBodrO5myLonmURzsa3LjaHfsz/KsR
DawKyaCzFYUeAR46/mn09GmHMDBL6FCNxtFgD0qQIGEqKajUlGNtSEead1nvgdop
O31DVdEv4W4vH8kg/5IEUeaD52lZyKMuhQ8iIpmOBmkO48/Cj3IMLGb9j+EGNUFn
Pjo1arjj9xc00bMEi0+ssaupWMQIbM53kbjdnNy4vECWpizIqE81zlwnaggHNEPC
IYXNldy5h9Mj6j7IkHyri/RksXSmLF6FCExnzIhqcR+d5oQ9GUDYhSQgiQ/XZB0C
ZKGnvUgDCpPuIhMzyH3gJju5pMtJisF0qWJIF6EBUoWohevlgNmbGP18wzC8Tqa/
Y2XwWIALQHZkz7ViOcl0RN1MLra3c6BBMaW2xr2+H/aX6Bl1aaFUAsUU3/wR2YPz
6M2yC+BHavMNwNQgiLU8GlL0wJu3apcYNfQMw4L0mtWtaZzvkDfte/wz3ix6kieg
GVosNaO3gZI3VhQLQKZzYlOZGM7VgRr4TnZtwVRk1QFdjVRZbEQvdaziB1b6OVmy
nAXmsI1cM8wwySIsfjaqyV+C1Wm2TIihxLZDTrM6UrC0xM01dulDhWUfKSE9RweC
1+Lc69DKYF9hsLXar6+blaHk45E9Qj3JkTPu/CLq2jI/XUNFrCecGsw2lyY1B7qO
fShWukivXmeonRlWNTcUN8C2fKGn/i73Hi8tOSGI0BPmsG60XAZ2hxFug3XWePAo
IzQ8HHbwlqQPHlfzKhZhOKoORIRruWV8R9NFff7rwKxXKlKyimM+oNnPehipQKIs
MzhavTlWNQiAghCnq12nfagvs0ShrHkSrd9U+4xiwutshKbV0r97w6/+kiWN4THp
lwQOo/u/VfeOilOdwWs0uiRgRRzgHxAv/buKiVGZs7qqs/ddgb0pMtTSpRCKctsg
VhiZFh6Q9AJVPTEZKauwUCdfdfa9A7F78qtQjNaFXS+s2X2SNIrO4xrBP8vnVFwh
ChsZ/RnJmNPH+DfQ/QGF5SgU9qaT38mGv7t3E0y1xAc1G0uP29xAnKKutKLo2wd3
9u217LVotCvV1KqyudvsZC3TdSNSQlLnXKxOd7K8nj3ht0/h28dkI03qnqRZGXvF
8pegLfNv5YI0f0ojAiJTN927wvdy9AATYUcJc4iUuCN/E+M2hyIbMydpnLH5CJ8P
tjE7JF8QgCuAH203nrOmTtowR9SBi9OUQMObiEs619wVrKSt/jixLFQ/ZNLYJB+h
hsOaDbtnzcukkSpfuua9K5RYmmxN5t1kAkKqK9v00XHfeHO7G4UE1pzSR3LEzXt+
1boy5KcPa/+eYPvxcMCC1zfQ796mpQVpthQTT/9s0vldedho+AESxkd7kNdC3N6h
+fm47OTmg/DRW3Thm85XMpoxR9BNruq2Ne1qMwVDFfISf+NA9VGeosk6ohzYWOmz
XT0ydrFgoQgP2kmJ+7dLQq99HdUShxihJfzn7yBy870CBENeEqeJAujImDHLzsT8
LBf0Lb3LgkFGM30IfL0XZ6j5MEcUFHMZHKo0IOVT4+HEHtB2oTsgezX/6obIbfCd
bHS6Hgqz2/xbXwuNMnUoweqirxfkuj1LDUa+lsoKRB24lDXZm8OT0ci8eP7JeXG0
WrfQwh3QcsKVr59v7oKz+aDkllrEgS/aaMk+aLpkuv2uU2I+IBDZKuho+F/X6XUm
l10xB7GkJs2SQMB9vWzrgmU9keMfuRB8eJbPd9H7DG+S5xDduhA7LaICG3TyzVZ9
HDOal5YZWKQoJVfgpMUHWoShEr0Rnyh1Jc+/segOiNSajz3qVnF0+d/c7d50e7+c
YntJa2YaKhmMlZ3xkflKqB/pUnoJq6icSN/MeKxl3XRqRnAryzFVeNe9/rh/7QQy
C/G5V8v1smzAnalw00gi9WvGh8840J2R4eKUd8xp/TYEpEyJrgvp60+dhLOdnvVo
uIOk65oF/JTyqWLU44u7F9a9so/EfoplIUBlcrLEydF3/G1xCAIn6NCySbsRDGas
BHLmq/alC5p9WN7S7Y2XGYTMPTj2l4JiF8rVx38qUKxQOb36Z7uPC/53HYyNEYIl
JBxFt3KgQouAET2vHaKJKcOvvXeOTu5k1bQcyFLSBYREKJcJrVFajlrz90mIkJ8M
xEDVXr9A54iUo1QAi+JEpa1TcR/qLE7p4bZe9DpRlOWm6YmToHiSBLeDNK4uvtPb
b/qvVKrvFmbxfV+cb1sX0Zjz6HTq+t7olPqybBBpL3Ksrud9hZ8MB7RDFwpaxODs
r84X3nu+koBnL3RrZKbeAEPpsiok9CTN3jDnauv1PVqio9LaY0RQiWMeM32DVgpM
XuI11ikMY0TEWfSttn0RHSMoxXF8XPUGiwjrwkRHaxwitWe2BDrQq0PueEUrjVJs
4ol9knZXPZIK0InkaxfHjLO2jMyDPoW7HMDguuMoky2619ISOTdC7Sq/+gR6PERN
OCV4tJjySAhLr/6YpsTH6I090WNQwjFkcWMLwdIU3FUtxBNZbB7TREec4YMUnTe4
vheI41nyI+73tNCsD1NzpziYLmzjg+FCZBraLk/7FkzS/VzGyWD7KDxarBDSjU/4
JOtZeiPnc8B03lz67FLKmD45BrgMQCSDSsxbcVokXHrFw1PmkKmUT86zh3zp78d3
Vw1iEQVJx1zqeSEwB5/iMueszV7Qs95FESZ1lHByf86LObfLKenxGLEgh2VhJtb8
BvPFWtsato0uZZ4J1H732loiNOsvraf4IBLZLTtdUm7TmFMEUJzTD3CNYPtx1phc
T92xx3R9WFfwkGkKmRC61fQKU2fsLINaXbxvIt0uu7eMnE460SWVjYqiKPO5zupl
aGfOmB+/bf8TPLIcg/GWYSuEfstA7qbb+qgsJV6KOHdMWQJN1vPVHlIlhMSt83iw
gnjpsbwyapshDh6KIVXCHpyDI2RS5PxWEs6X3QZzFX+BFHre8x0hjvSw8/xjMyUv
4UP04zzlQOL41xDscXOl4z9DiVg5d77yEs5/Z/DB0W9Ba97m8HZghRfLsKsxTDrW
n3A5Te3YQxxfgP7odaXTioi0OyaTl6SJAmHho7Kz2fgu+uL2VaEJoBzJ/uBm0JGB
SDPqKuHbbxFGx9CJEHd8U9vAaAnjSvCarFogsbYdZimyiYMjoeVV09c2D7NWJrkg
Z3YrNe+K40sOfrITyaOEvL5PFA2cedFUhizEIXeD9EB6/7Bx/rCxqaR2/7I1uiuV
UsWWWz7F/P4eMioLyuL8e7VKDC9VVADMoCgbVpJHlIoZ3vP/BjNJYy74WjG/oTVU
dygCW6MAxiIUEbo82fJmc9EwTi6R7U7tJBotk8xIDsab2QTUCK4ldIATwlCFGQgK
a6kax7cfAQBq5bvrqsd+nzw/p3e9vdi9DiQD+Gl//obrY6Xjxnbi3hS4IacwL3vU
XlnaPllmrBsfkGjz5deJK45wCbHFTqBuLsWtoX9xNe4qRpwmt1fKLqbo2Nt/0u+G
8Ou/z3AL8M3TvLIA1nsSMD2/FPjSjQALKZ7wFcai+yfk+zN7vl3+284MgPr64VPX
lnRy4tVFR6BJJs7+7kewFNVWyNPElK/9jkmbZiR6opi7+zcrdJ4tONZ5ZNhqv6V2
k2Pe0PhrG97q2+PvoNUMbq7BT0WPSx5svHndsiO0DhtGULifcbAIaQeIqYfR8Vgo
xO/ImAshdBpud8gq0atLWxcnC0yFnIOYDohIYxg2A4mFP6eGNq21Y4eFQuQ5s28l
ht9hv73L8WnBo+eNKjcZQX9M1FCO6og+C/avJ57XEXadqN/FXD4dAEOgAirRynOj
B15L3Xy/3LnnDZvtHR1N7Jm+OkL6uw+BCzshqj3+HWY2Zvt1oaYvjjk+L+eMDNIp
vQw6Zi8DhFEeBbHS3Y6aputnNTqc3r5musj7t+gJ+XgvutOGcDTru87g5TgamJ2r
6N5hKefrhz1HwGe7XDsqCPOhUocbzx6yA8lJlhvYp0UBbEccGG6z1H//azhoQvIJ
WlXN8MnIA4raInRnX1RMHUAiJ9NGHbmPV0ugBMd/Vt4dpki0KRQFX0eiQizlG6xS
MSZjGnd2WU+2oMmYE0vTpKWUBoa75EUyg2wtga7mSA8nX5ckOm2puALeFv1+XtMR
OH/rpAPaxEPev7txTrguka1uRmlLYcVwT/Fs9xxbPQxB6W5A+EDkwyPvO/j4TL1W
TqPjjsjw8WmCqJ3d9eWW0AMNauD2j1MJf6Hehb9tLZlBlWHpuBZsP9HLW85237oS
d7iJWKDiOXRHlxXtPe2To4hT8pTQujdcByVbchd2//AK0JQhtADu/0yu/GLUBUMu
tag3f0w5fb1HdWQ5aEgwabTULawyfsEO4ZX/LupxEyrRm0WDslHv4qmJPJ2M2sw3
Xr45AAXqpb+he0QYDvr8byACaLy3pGtiSWfo5gkUJcGoT7sPV+qnHuD7rbYrUZzv
kpspdGN7Ox9UrMwY+h4Z2eRMPMbJHmal3hnEfZ6BuAte9O1EVY7UiEJy+6mUXFd9
I3XkmOqT441z23bEASlMwwpLqz12xlHb7LrAwPW98l5lHjwqzy2UoGKPHOO72uYa
LHuXZnPc2CcbRohNyWZiqrAW3ESlUDPN833KOdzonwVAX8GdB3tPfJUnsgZuMDwx
gMlgf5AipSzXfZ5qifflRAjtbzMzwW27YpBQC88hBfkHbwvPZ5XZ/wmfweGJN2NM
c67nCXpcVdwnGsCsiytuxZSCZW54gSoBjr5XHAC0RTS7Rex+vl2xW/3Lu0wvic3e
IVmD7nrGc8V+E8q4rM0dLSwtVf8AsO4VuYyQmRTwLKDtuHmA3BQdkFAeVcNdW+iv
H8wMgJJlFzVOdlH4HmVflpEfHCCVxCZATCYbUmM/31iqUuaeIU4Jop2fxSOaxofE
kjRy2IZHJRT4cI+hKtyKP57sWPeZCXv1YoEXnaxyxMnytRDSVGVIMrZP8aQFlzaK
2a1d2llZN749AHSYlTCR069abQxOIHk1UnkFd1yPF9OXi3iXY/+rGVjKzsi9x2Cf
rr1mZZ3cUBVMBjqXJHkKyITPZ1JVmHBMM+3M5UlOeljRaTxbdCVbW2+tRyYxuEfr
huWkvDQaLRbgCzVtIWyLsePZFWqoGAH9Jy5ZIrQGhhATRGWqzS+GYt7rJUXu+CgG
3D0P1HOoepyMCIgvkmg54IADxTbToBd8SOq/wzDKBtlJu4Kh8iV73CY53W3uIrj8
IJR6t+JVbk0/wMkxBbkk3ZTcDTJWHe0O8k2OeFayJmRfG/GUrmwvNKb9s+CAT5q8
ofpHzEo2tlO2z/I5cy86wlNw4mfboOj8PlBaxQseMqoPiSvGdksshzFByhryijDF
FZgBI7VLJmKyQ6JKKsFH17XVT9+0VrsO+CW5xkMoDElJ2cChxQ4wm1BL5G7ZlLMo
do1s32NoFrO4OuagJYroqaZdSEu9ttRcPb7mysQHqIJUCio1xWS5yHHEJHN/RdgD
0vZAl5TyhG6bqKclOSQoXDWF5Rs4KUbHZdXu3IvH2AqTioigpvtHbwhrUgDYsvlk
HPpEBCinzxI7L6cZ3ldSZfgpvsVfrd8tLN74woBU2s2iDK/sWXdEu/bXwIzxI1sK
D9Zs+VDPxVHdKsibwK9llSqP6ZTCnhxbedzRty00Xi1+boJRxVgmqSwenJl+Pmf+
JWnhl9Iyp/DJN0Az3w17d3AYHILSzyboKGg0zh/o1TO2CYBfdF9ZvvJc7aE0SQxV
hk4vzwLQtqwM906B5/ULY3S+WJvOCJ7hITZ+dmM6u36iruQ21uTihTcbSxojWTem
5vfzYCkyMEhWXT1IJjOLON+PLIbAJUBqDHRszd79u3Jx383r6DgA+yMvMeUIViP+
dfG/tbcFlvHLBjjurd/OAhP7Nt/VstxVruQUzBTIdD331R71TxZKPAvH/FURpSIG
OMAVRNvWKEr/lzZVB9U7tZxKCO8B5cIqth1r3ItqEbt6XPFfsNdtfuyi+2L4EcWh
uEnl8bupLyHAvHDI4H0Rh2CkbUFe/39pvgRfODscr02/F1UNe64tOBN1OrsIz8XT
m+fCDEK+JZoz9ytrorWWCoD5QFwdSWpKkPb4OkdoSYIbnJ7Sibl7p1qoss0Cj8MK
9q/2WhN6MgNLZbXTFA8cyk0I1kUoHabJANeoknWEKmVJE0UoBctJLU3JAuPxTwar
bTkhp9z7jp8sMPMjhJmxMCcccH6iEzEBJhgv1M3B3N7nTjAz+hOCjPpE+y7Z7vOz
FjssZAqJ34dBWDdTbCIFIWj9+7jv475PfK2YM6QkCSxwY4yi5mDkfK4JzWsAj22v
LnpXQT9HtD99a43Av0zNw7wZELJvyPBPAEAoZ+3TmdohN5bUi/7tdjny/SgH0bKr
TReg/WM/ZVH1+frqNdBnUDd7ao2roWMYUxXSd6gvh9XJVXoSu/eq4iS3jQcsgqT7
jrwqKQbJ4demwDGpxRaQxkEbG2sktL/8iHW5mRBm1f7mA5OIXXFxnutzVcO8am6c
v377WbuOVE50bZXXDXKsYLrveUJYO6c9ZxtQEr1LEHwh61M+X7a6rwjTS4XHJY6/
H+eivR1gymEzCdb0GQ/LIgPytD6hssYbvcvSb/QUvj3/LbEcTp8nGUGSQtJ4Cksl
dppdIOABfwR3mlEHaf2Pvgb29ecaGOKIfWQGdUP3E01CFecvH5464EFGbNZjpZ8g
u7qq57AeLBo1rxuai1o9QMDfDr2FuqAJE0b6SVomzD+c5iQByTdIQ4Ul5AhTs/XO
rj4/yv/UxxIdJF4bsa+AYARpDqHa2sXoW2yrzpzNCbU1d/ZUfqlZRf6REZq5kX7J
pEGUTm1jmtvqFlxq6LvTQW8PjxmUn4Vj0ekGW317aiCbiXufFwF5Apbwlnbx2Tcz
QrlVRPxe0n02TYUgg0O7skGk6PmKYLzNeC58L9/QNtx49ED8Gq5f/bmA+kKWK3jo
PHnsxzN4IaKP3wCwfTnc57YnPqEsXS/ZclZ3VPzMJtwSXXxQTHM9wiQj1FER457U
CcC6I6PjFYXgJXcq9sH79a5kxLGlcE/zomHaGnQEdYjk+ObPyxUXGE3FDIfHJ3w1
8fuBuIcvLOIuJ9l0yp5hfdHZOVQeeAJWdZ7dCN3/bBhCgF727WaLoFrMWDLwt8yi
Uaao3lTEvkTOSB6CQM7R2k/r4QGzoJYdlZp4SrCsdAHBI/TEUx7atVCw8EpUvrYd
StauePPBZdMIMp0NoeKVnWnvInRCRyBQpKretu18R66Ir+E7mHa+CUVZjg9L1QOM
fFI7VkfKsK4Sg3IDJpr6EYJwFiExuKvQSwueWcWHaB93IAiqqH70c2v9mepm/YCv
Xfht/nerZ1MfRDerT/AbDU1jaEexNva2JdGNziygX+O5z2CrREtsl00NXPgZFnua
/4rg+Wm0RHiWf4qNz7kLhWNJbBf8JTMMXO5NNgEl9BRM8F4oHL0NsuIyJ9ApGJAj
2NPHd+3jjz6RfcmnxUe8qXyih8jE6iB190zfMjsh819toywM2/89rzoORRV2Ew0F
GKFYjfIpVs90OpUzOc99OcZwZ74jLf/Z0tTWb15cuBL7/je+w6+ehzAcVMhi5IZx
3vDqJieqQKI5Rw+QhbmE37PG+8mH8tSjGsqU9Ir0zZem5lEFcLliBWQQFpuB0ytM
IKgFalh8qyqknCoca2g1t80ILN14+L8nkj4ZLcipYVyARrb+4aUzICQs/exsq3bM
RLMVJX3XenUZyY3tYKx4wEg/tnCJJyBGuS3xpwci0Qm0XwA2/5iJCfNL/j1GEWot
RNrCFfne9piUnII27GPj5w+pBzvYeUcU/QGfJ5RGSV8AsiYWGyBVvYEqrIk5+Am6
ym2gEHFmiwfsWB3f8ZRo+kWTwjAbJUVhHbtoO3qHtjIpv/+lltJTjUhcLsQ6GD25
h5IxPoeNQe0u0P3Y1K9k5XqN+TAeiALYeDiF8r6UZ1oCUKBqgD5B3opxkXT1SP0X
m29o/gdclYFdGBwYx1SSLsxiNZCXHR+6WAlv5t/vm0Pg5KxAPdP4Ntjvgv31BZr4
8c3n1Oq5atvLobRa7IN3hpVunjWragvJAvq+yZ0L2GhMy5E2Dlj6dUbqshQ8eMEW
NkjPEPEeF4fj6A6CgNaJivaB2XC3c2naSEeVSNAMPl4YWwP+7fiYTk7jenGQumAu
bXJMAIxDuOfBboxps3uhdS7XndIsl/j42yBXR1ZDPRTM9HE044D3hiSAYm/gXJhh
9cEzdBRAfkqkjnGoMEVXB9dyNzPJTi7/if7X1GX/iEnLnOLfWWao1r3LoBNaRf2p
p6h2yFGD2I8qegWq/qHvmV/aG3IB+uG6Ygv7yJ4WphyTFmC3AHyFTbVcLGHv9PgD
vs6JAOc7JnV7TDb/5XKaR3PLQ4yOyS5ZF9sjJAfQxRanRq9SNxwycyJYtUAzPbiT
aCo//U+PcwUbNaDKS28bsrACvsqraIQst8mUgMCKD3cJ6ylyhovCu38gagaIo4eL
oCQmL1e8Xl7uJ543RKrodaF1j+qDaVX1Ad1xrou9l3M8l0hoxQvuLWhVmK3ZUp3k
SgLwMCmyXc/r78jd0E3bIQrc21t7n/uVki21D7q9LQAyCv9m9YtW8Cj3w3N25Rad
7bUP0aT5cYP7SmHXl5j3p6ixf76a2yYyHcjJ7P5fY0rD6XwXsYwO1IovdV5R7EH0
kZQ3bWgXGZ3A9y9V7NVUqNpwCOVZeOIqnIY9JU9B9hEI5XQ2vFeHZafHj1ElG8mm
UVaezELuWrf5vH7oNOGfBAPZsItCXgSwXH7BrMDmO6S9tUC+tIk4hYGrrVvyaBOF
c1c37x5dEFlmkIUeXYSSDvtRneWft08lwa9v2A8vtDgyBtduOKXR8EaPojZEggcL
5VnpFCGhdEiSQ28BDKHDkBq1r+MD3MTnQ2dGCEIEzR6LUNeY9MnY62ZEvo9ZDTvA
/Uf9DyqwkXNXETlwMseiUhATcbXsMAkBAmWQHqKHR5To2EffKPyLwZ6J1H4WIGbV
MdO06UHd0yep8GWZkPhrO7fo11uxcWmmOwNhnzx0EBUYwtyVNQTk8kSctjAvJ0Cf
jB2talYmrY84PfsBv197HTxJB7gjC5bR7fIjKdm5XrpJi85AK6BgmvUhOCeQxq4E
96Wr0e7bVAVoeMY6NFSzagXALsobpFqz2bT5R07pDy22sWO6CH2tTdWcmB4ANThe
p788MU38Wy8/eZ0AfinneMgbGsqMvh1QPR9MAsCjCmxu22PzXPQMXzNssZ5qeN+H
mbAJ8ns/v+g6ep0YfHoAjICIf7qJxjDtrnVb5xQ+UDW8a+T4IAjGR9oMNquRe17T
FpFqAdv5UQR4SQRcw5GU/rIPd/Nt2wN/F0UAw9akG3FqwAHCFMDGtfyFkQorc05d
esjzEMsS2y5f3KYt9CqBHXDORZ9YvUEsV7kW6YxyTPjVxopkZlpC2Hf0CrmTWKgV
rA/eFypFV5hW3lq8z5gVeKQSrXIhDtXKc5UxIhfhIYbNA0X2H6QyV8CUfnrLWNoT
oSxMe6nZH5bDALMZq7ee2jat8twZZhmxxiTCzkbQnuH2M6i6apqQSdxg84cntZeu
hs9n2PS1Uak1uXpHqdByIqpzXH+OPO/9G5bjlCdiW7K/KH8pZ6aAAJlin+LQRvNg
0OQc/rqqfUD5bbMHi7GDWY32cnCMMNUZngKG9jNOp7oRmP3k4wrszDgKl/Delwy7
pWJZfjmbHYHF4It9lOWbK94eTTRhxhi3S/O9XlP6FEOOjtkR8k1NJU9lvTVd7MV1
R4BW0GN6AoOHAALHM9gHERkrUnfoQWlSccBYhcP8LeMIZSfDSZAMgoR1DOrLN3an
dr7UHCeUN8wgk82n6hlHLsfzGQOJwbceeEj1mHAvTN9sLKgWa1pdei2AUfUiPn6j
V3B6Vf7r4mxURmgS4vkFCfQb2LM9kyAmex5whyR5onRsVnO5B0r8nBn5oP3d4de9
9jKVL7TuSxCv9DoaXJVnqPbp0yl5osxc8BNIDiEkaIqzdnHtvlihQUrCFaiDgd8A
kxrpozhhvB5k7T9+oTvu0/ilsQ5GN6Lk8C4MZwrt8/MAXrHhhHRmgj13Z5h6tSHj
uhO4KEBKcIc6+rd30l+i8dMgv7zhhEGN65iqNd9nSrppOTnTFcuKm1bBm5KV9yiC
S0Fsg+B8Nqs0RzV1BYXGSB/Y3ZFZSKSkPyauwy+5g8MiYFjU7wutaz/Qq/VXaFTd
aZAHGP7WZGdqIufg8am8kYCBIOT0OM3CraoUt89kbRNUJYDsnX5ZeYy39PdX0FEz
VUUp42oF+zuY/nwo7bknria7LyIQFnacSFAwh+ZJ2eEODSe1RrgsR4gMcpC+b/aY
7e2OYUrDH6wsS3xDkM1HGQ+T5PLokX7ZmD7eFMd2kBgTW1hSTaZMaiQBZQiaO2uS
v6ug35kIeRiVM/SHlb/s/yS8bBR1OXabrkJGkCesYgjlpVi6Gxlfexv+uCw3xiKp
06FIZoG0Clhyg9HYf+cctyDJSOUUrQN5Y3pM3GaYQ7tERaj7hVuxcyqEAKewJCx8
U8A8OU74aRUGGaKWXSKb1Pv2woXuhZcRVHwpAzriXbzCn+3IPPHgzdNkbKujLxNi
QJLrXrLHj6mzNR/FQBdcHo84QLBtotFrjzlmek66B/SPh4MyOuD+22jfyiEc1DOe
knlLCd2BCcgZPm+xGQpyZv3OYqWDBTIt8AKyeeBM7hS1CsnXsOzyh0Ii/DU5q7gp
3Cbx6sv1qLtm+p2K4uvPBjbyn3YZl369ykQCHZVd3r/Q85HMLrOVuTXleW/a4OS9
4uHwFyrDIkqyOTWa74LmZqdXIVyLb6i2WnlxKSNB+s62PIcrdDKlVWlDobZ/iOeN
tkI53GjTP3pfMlb58S+9FzFGhPVAPi5tj2wXgQ2cNSR5hD9+2QmdbRmeDyQ99ffv
wTSPHk30ISDzVXpDw4NJR+rs7MDGNzd9iycELGDEFl2OATbTGGYF/2LfsdNIGPX9
Naym1P9ONsChAxnmJbyAA5cypr9rxIX5GvHunM7WAQ7Vtjjgi/DaWQmgXJjxDslR
sMjII/2dxd3p6jSOgXYbER+9mIz/yailG5DQJe5B7b2FBuZba+KFx+foBXhwAEBx
42X3Nyqa/k4aLP9jHs0VyrAZtATrgmiFUdjMkSA3NEvPOhI94pB/3EDEZBZcV4ZT
ncbrCuEMPCn8rOOJHBde1mNR092Q6givh444EBih/eTJ0oxwv2U1reSOqC6LDS3z
64d6RqoNwA09sinaxsklEFJ845JRp9724a+ByzdK1moLCKQVK5ygbwOI3rVUxxPt
StbV8yw5A6n5SymwYIkC3vUzet3VFLa9GvuQLBIwFjQnljzqzkDBOq53TefeJxj2
np8DzLGrOVOfE0vPhV7ZLOb1DkTPBFNyY/2LJ97RGEKwTkdxkNAMxICxrJiTJgWf
W5spNb5avzpC9mz+A3kjygagykm3CbvWNS/xsSNRKvLk/OLrog0HWfBgVYjytdW3
sZVdaPLT7u0Ku6mTKvCRxNfOGqE+0hy7BV5C6DNYFiy1Z5sHOl1UuCSuYqZdgsFN
HVYTJCj0zaxnZQJBClZny1YeC9KZ32ugfVGkCtGGXEaqokuMcEmzKQ3WcLGKhoPg
ROuw97Zg9yjpoh2T6NNptavU1MdmkeM41fJ97UCAO0CtJ8l0fhYzmmoiYIamOlBZ
75zGsU6ySeIog11NoIb5SYjMVOaoj560oQ72UA3wWCuaMDqEaMqyh0SilujXZGtI
meqlVT0FysQlfpwYITUja1K4wR3QXp1u1EiUkXZbJTRmAGe5JKCLNmL4JItGwmd1
IkUgf4gHbK7hURtcUMblY/D9YuFPD6SEuQi9/ZBsk+4GTVH/r1jpsppp2KhnTk57
wqh8x91BsVLl5k5CJ+WWvDtzD/bGxeu9S/n9HuXjjPByBWA4qpUKFWhSHbIrisX1
RjNkRLE9Lf1PBKAB131sdmJjyB/p+qkKT1vwv66xp1B/XGDF4dRt4HMFTcWjly3V
js2OP+Km3qBkGDjqdQUTD/0LqdNgzhsQsIYwAXBWILq1+uKqFrPT50ZkVrUVhM96
1Pb8UC6wP9AHqTnLpelLGT9bRnX7Re/4zX10mKoDdL+qpNSr+qsExjIVLzy/RWJ6
miEXqdTOorb8QePWapd0L8gr0Rt6/S1/E5BBA75ck7uwPT5yrWJ8LUWfzvH5kdus
B5OvHxk1Usig/xVNlFnJzoqIVg2FmHixf9i+kn0skfOtCkqP+vf0C/o2bJOVm9Ak
VFL62uBF1JsHuwWhFZJKb0NgvHLz/lsxUNUySDPF2DGaiQDs9sKqU41CEsV0LK0a
SI0sAhnz/ovMPzXk28h+g5mcSwza8Fszri+BF9J1Hox9dBbqgaJvmpsZiQ3gYMmv
Eul824NLS0PO60Vc47oakwfm4I6HZDxAYjD5tUrlm1U1uWk2HUo/PjVL/lj4r2Oe
l3zocjmRIXFGIuTnn8X43dn+rfcePamFT5MDZ5zNY5ELIZYMaP96nWxM8RjBlL7W
epvvR3LHkdPhdPsEv+d5ZvM+zN5jEqHUiRCKSKjUgpXII3Uri8sejBvWR4v2oBHY
KxawUeBOYbMJoVJ/UD0Bd9iLHlYBFiPoMlA5GlzfYg6tnWqUWaHL2R7EzwD561Oi
QLu72E0c+zXLEN/I8ABIEWMT6pcT/mi4TADomJR1uxs0utwlGZW6cuqxa9m272lK
toSQW0Yb9pbt4e5lOfezKnf8qiYtB9/ZeDgRG9GjcMC9U453KgxWlE1EA6vEAMCz
1RlkuNJzw21BAz4JVXJrOaUcqqCnhgzGUiVcoPPbszALTjBntN7/bnB7FnlfBhrk
JdM1v6XeFBU+iVPZoei84e5g9JAZaVL1f0wvSTCJt1YwTC8En5lJDs11Wa8gAC7T
yTg0Gl+ZSaMA2d2jkZoQTN8xmxVU5QYzNbhWpJu5b6ErGU98mxvZUX/ycN2pWzoh
T8na02liLY30+ByQTUJcB6KBpeEBs9mbycPmxZBHNvVanFPiSEQ/XdTVVw68XSVe
vim1YKuPZj3ic7p0rux3g1ONaAeVwM8G852ZfNFkatlRirO0VpCl6bnnmssA1TTL
edurzqwm5P4kHKfRyjA4pmgEYjC3lx+IqpSQfDTl5E0E0LvisFHW0uJuKz3LVC4e
diUlK1dunEEFV8Y9zQB5q7L6FvtpxPppG4y8tZ/ixm999fI4gyW5aYIlXOQPZLQv
eFQ3v0yd0Yx1+IDIu9LQMmMNBI/Zgc1xDPio6T9vngH4Nji+zgZDX6u3dNA93tQV
l0DNQGvsdQvNiV3ZOM0fqmlQ5E9gmq9nfIOg+pm3ym8010GN1p9kOLpi5pNT4eB5
oFjTWRApZyPC4FyFqvhxcp2uRKGUiQWM1WDorwpmC/jHtuKkVV7AE0JS8ki+M//l
Y3EmwvuI2tsRgzwONgM0Vu0r6CT5GrB32QbpwQ8fLWj0ic2tenpVcBY8MeQ/fzkV
x9wRL2Br4aXBaqTATQ341LL6G1TJd3wGWKcq34WsJkAw3KFwLmePdJjlrHoHCeOO
QvzEcugDzwWmKBaEqFQ2UYTxd9esh4Ip+zD+xpkWeyw09cQ+lcv0hkyLLL5AzCUQ
thJyAikxk0ncvfalNzZNe4IeMEwrCe/uFufLBpYrFMEZIaTU2vq7srlg1KQdtNod
DDgfH0Bgq0uvR+vJbUIKNYCxStj6U9jQSueBjY6q8SF6LlHc5R7wzYPTtSK7i+YM
IgLhqpQyw8Y0jPkm19ThyW6Bb00OkT+bCmsbGD6lDmmAiXOE1D/q9Qeu2dnxmf7K
FMcA6g9xThrz3iCJCaTHi9numszBz+Ge1u7SqFE3stvjFGugvI0bCJFNrYqfEYJ9
8nYlxQRDUKQJfm2DKRFqu8CVd5usUiavCXRQhs61Zw1o87JYy+bY/tZfeAMMaqbp
dSCy6iMQsoUHD5/l7TVWPnQOrqbQsTPZTZqt360MSRUK+vYOWSUaeUbSbotkNMzw
FEQeuD/BI3HoHXfBdqy18E1DIBJ22kcxG1QHqeRZ/D0reGIdFrp9ldilIlp/kL0W
f/lwnMdu/DlWiJPyqkeA85EhuFodz26ZIxQ4/OStngYtBfYSl7/qT8gKn2LA6Qfv
v3rDQ8nEoCeReamRKph3Tn31ZmyPtCeleuu64dHwSz76uMIWwqWtFThVkAKk17Gh
Y0HGB3EE6PT0z1fDoISi1W3M+XrnlIljefD681H9A56+k321i596rCcM4BAZOfsj
giyrNtZsaELcsNaSGgM671/x7DA4qtJfcQuFy1qKMWCy+Y02iEM9MksC2EmJ4q3p
zt6QcME6sRtjGhIj2X7mNWxA07ONEeWeIipwAdkplJnJipOX8jEd+Bh2RkKRMvZ7
C/hr89PuSW9DskRBh/FGEi3f1ZIKczi/vhKnToYWdd+6xnfAMvS+34O638RQAbUs
x+u5DIlHsEeMgffj/u2/v1CZGS9EgZW4bwnIuJyYLaHr7ayRyZRgtHJyzCWpYbcd
VP2czeD5Df6qqYbtR+Z/rTUGDUY9+E0RN2CBn9gCXGF813Je0ZB/k9cd+xwALmSn
8ASu4X+WL6rh3SNDBWCNAbnFB8VKHjY7z+EqQfkPKYK2H87e3qzakfJiiz1ZGmsR
GoVofL8FW+MK/u+WTax6dFd8C53VNYnUYURwrj2HdsvWHoIo3kSPFsGmXuczY3o3
xRuKj5gcBNdEI9BPtGWO0Tl1XBymuD9VAJ1CJVGVM+xKetVBBiKOFf88LVXIed7e
YOMbvdBiTEJCq8lwC1Azu/0bhMYzkWIDLGK3Og2EV9TXd/QcC+v8BNN3eBoUvehB
CseJcrFdUKCM0qEmUFiuleCNmzj6LhrgchZyJ4/zYALujLzqP71E4RfTPhuGIIgJ
37Sxp4XR6MnThjsdoqh00LdPF5skitEWIsQjMVBPPTBLCx1x+D/wI1yRu0Uc7nN4
hFwliVUIYrNjR6zH6WNS1GTpiyU76hZBo1xr6rrrguPOW8Ly1t/llC8xFErzkSj8
fH2SOr8YpLfSRI0jM7V/upYsvJwsLxupDkmBk380reGMTK1HE1IeKCS9oykG8/bi
Mb+YMiQ+fKkJ2ey4tOF4zwkKjP88UEnmMvrWHfjFIyb6yRxPYt9aEigq0dxMgOdc
ebBlhG3/AEn5y07mE084zJHqshDHvMpEROKmL+X/kJRl/0aVzgt6BMApovhej1lW
3/sXmv64Y4ErjnDDQhjDqHzfUvRJbSyk8uXNgGot9+8cqqu3jPjYTBzUVRZTjqBi
eDqeMtXTUriopuMfPLFV28Wj59iUiemkiM3gM9CChW5wTFWEurmWNI+3cAu4CG5K
FnukJv5MMfSoCpHl6Qh7U178C3YZ4+VjMLaQ/zeZG7/aVSV85y4Jpa5dlxIu+rXV
GsM/PxKX7FZ4di0mBV5HGVFA45DLYy6TQ3cCTEP4mAff4JKLCCfbHFkNmcp5Tv3R
c6sxA0EJiN9ZedpPlLoFRsDXFXmUBPZ8kVV0/lB2Fd4JJXG/JdGg5WZyZJ2vQlYm
abO2NHyAqp/fN55QAeQI7ynbP5DrfUKqLwbX8lSAynQraY3UjprGfiLRHS4B//iV
ECN71C8MnwT5MThz5VWU0JxR7XRMjr3/eL/8AzMbgy/dtDHaAYKSFJHfJFfnRTLA
4ZGSw/RvkoFo60WwoKOr2XwDre9zslbkKAk/niZal4weXD5g0ks4dSabI/2MkX9H
I5dgH7x988Qx3u7ymCkU887JafXDDtDhMwF3WSGCdkJ6dxPCriWgcuhvJ6A0AA4G
CkLmp6v2cmyWqXXp35vFmEg0gg3aYLnBwDZ2sLpN0Pr4qYgmx+E0xE4ttaLdvU2a
wFjmkqeqy5bB0nMP3TnxlbEIl3AcOlUGN1TOvbd3/C3oIEEoQMcA6Uve+k7phW6K
qOB3c3zIWoLw9k4HxUv2vSaxPqRo8Zts1dkAQIH/Yz2Zrphw58rMQb4pmsb9MXQQ
nu6B1HcearqX8W8ka6HVDxVaLPi/CFXV5XI6Ok0LvJgPZ8emY9PABSCckQFJ4DLe
7+/C+tIn1OCLzHqntoZamxij/F4ANkcMstMa4ShtmMMJRW4xWTKVz+haVnKQq3j7
M30k71ASUWDPpbH/8khn5DBM2JOJNZKbr7v9eUR6eNzB/EfudBNE39J5fa09ORX8
p5yxFa0RJsBNh/Y5VUaysZoPMwIrQ+l8HP7vgpkBrbmgdzG0FIvwyjeu2e1abxHp
xJHNse/AS9/ezX7TPJjSBbM8mtXgzFD5R/YRBAKiCjbnY8U4dp5i+qEMJ4X/S6k3
E/JMf8jINSR4Z4CU7B/Cdofuft5fd6s/KBkwf8311EgkqYaL9m9FPFtFvvFvgbwm
52fj+lCZd/jlnbtDvX/fIhjpgr5DSGd12I36G/bOmd3jQY1qTIs1VGhDnq6dC3SE
cmZlJ+eQWy60kxdVVKXMfiZnflhllJs+DvdFrG3HyKBpWm99TAJmb2Ijk5UqE/7F
VKVaMQ2TkwWAhTQh+x76EdS28l5OKe3tXNcdltVkeuDhiEz3b2y1/paDmXbo4TdI
aDSi7DR9mtmtyaa7pNqeuh9C8+Jo+Vmy8iTTKfSiaflE0mNtNtO9on4QY4NSHkl7
8nKTVKjbl77Imz1VUKsZvzgukegocjOd7odzcjMiZa2y3q2aG8igZt+zMpgqiV+G
b4HYjhMZPGrDVu0GfmkTUziA681DmP5NNGK4+sSdumshBgbVgCsQIORE7b/YAftS
vC/aFYFdsbmpdpfeHF+GcSgr9ODSPtwECXmzOZ6FuqS5te5NXomQDWVl1KsLJElY
a8bzW9PivDyicbu46/ZEPgW51GnelJg3INpH7w9l5jECygLiDYhC3KhYY8XVSrjt
VzqE9tEDRAJ+f1bLJVzFZybIS1J0WALNjK0QRkA1mowICKmItntLlGlzb6VtnsK5
s7Uhjz4deyf2+WvaOrYU0rUtjO7kC02cmEyroj5jgRJtfmy1Pko9Pv9H+6KcJ60B
9Zhj53zYJv4ZIUOYgsOnasiinYTt+L8T+/ZcWt8VKwYXEo+8ArGwiDko1cSWsPYH
LdhCO9nhQftN91KzTL7H+ZaBZGWEGGtvI+envOZktGb/217XyBe74/npNnnTQizu
Kgif5WzjY630mYXy5sOPJpXnnsNSE84XBFovxPBz0kTils2AR/uiuqsgVehX4MbK
P2r0+IMp8fipiOJGpugmG6DZtoHMEj97jY777d3Z+8Fqm0r28q3emXsDi2TVrrUn
24W+MMfFniOshqGGmg8SKMG30ONCPG444yF3i3FKAeCqVr0nIX5hxC4+rBPH3oZm
IVSajzRaFewzQrS9D5eCUnWrx4WtoMaotLCh5LJig8+w+F6xchxfffK7fRq+Ksv1
UN3mjMaDJbMaxzuY5o6BqNDusIur39abHxfNx57C9F6IVTDo+3R8CR2lTfnpzZKa
6CNO8hcf1FxAGj31D1SHEIqqqdaIZ1uKVi3Dn/r6xxBEMkQvCrBUhPi1XpV5Yy60
fnPnunef2SDnCSthE21yB1VLCukJMSU7EjFSkbpw2MLC16DQ6DnbA2gLyuOiWZpA
ONfPt3EmfSDbJUL3e0yM5BEgH2ncJbZS9OJIDvqu3D85kGLv14mYXntdqPR9C9GS
LktVRwr+MopmE9czQmVCyz3anlZS+O77rLy6fXclWog9gD+z/TdOhqcSZT6wPhLI
TqskKRWSzTaPjw3Vjf5WLY+6aO8JRSV7An4ef75KuBpf8WF8s9P1BLwAHmwXWhlN
UCJTnaL/Ec3q09Xck8fwJohvcub4vr3QoCZpSNbETguyNdMdipp6ogJvvyTaQOZJ
zu64ifz4R4mfU3Ub1eriym3LFHAUgSAm+sS556ytw6O0ziAYcrDGIVkb0ukA/67U
kMbMpcirJX5qe0LwNSwszo5PI2JfdPxti+tGB2LhKT/1+SYQnUteIf8NRLV/jmGw
c5RLsOAaafx3zleZbMC9+PMyxGRrR5zMGA5m1xcKescouAZ9KL+uaWCAX7ST8vVU
VNRnAhXaMa68oiu/zknpyE37ETjHpvm0A6RGqVT5jV2FLR5Tr1sPHLgREBEZnVAi
KerPG/d3wmtBCIZynA7DnL9hoLCU9NsR7Ca7uYK2OXm6LHeZc8YXMMj01JFA62Fv
dLO2UdGtb0QxxXZgfUZhAoIlvZCCNh3bi+I7M+Xk3n8SEmOWVJu9K+nbMJ0WXkdH
OCOKylmBEzaHLGZgiLDaAPW66AfskR1RIk5vPRd93rSeyt1hcNXJwBd756HL99tU
5nINSDcrsbPiFD2M/A+54Mdle6spnSOgQsWDH+BQzw+Mu+g8clxdUuNHgGy2gone
YcTum9P/+b/Kx+WiYPGPH6Cz6XEHfXkhBXh3Cvjls8yeWjyVpnJa3ofAWdUFtKRy
Oyi/LD5aCyKvIWiV5/0Ns7abMAom1SGYOPnYop90ySfdiZCQdP52VJp/4KJzvfb7
7CiAqTO9ondLD6YuAAp3hF9yXPbBS2mMzVGoWd2CTXJFEO5Z1TdirKciaE4VNcAn
0IrPtcP1IVWgMZJY7F894CZpKvcbs84eVf56IdOBi+Oj5ITuwWAxjciMe1ueMD9C
HD5nsKeNKW5AbEL+ihAOL9vC0VCMPO/GD44oDc0s9OLzr2VGq6FQZ0IYRpo4u8gz
MroShfZh1wgP9rIE30zkKWEITUw+jnXqiQN3MQqcBTwGUaNdBgac1TITsrz9gsCk
BnnjXWHxV/IKkluBhpisEMxbW4rP78CPZDGNdJT95jknY3+0cShbekHUlrUfJOSd
vJXxq9L0/UlDx8lUdzjT4XUQluRBP2trPW0i+0YSoTdsh+Jn6phTX3ORGuDrM3Ks
KwdCPIOS/PB1Gjucivme+xj8smcoM9wuknzeFdeyBZt0nbGeFSItioRYldj0Uhf/
dLlvJ6txT+XIzlmNSSA4dLi+2diHJIp8+XyCIDunbN2lQIq5Zr+RkhT7G8QSSdXk
h1yCgMx2du7AowCNPryLmvXkr3ydxZgF5XQPz4sGTnVL/hsToz7aNPqVFzrL0QNy
vMntv3O1nDSl5pxNonHt+hMgkoQLPAHnGOxM+sT35k3Q9SMxlnJYvMrrrplgFSGs
JljqKooI6VDwfHBHAoDtdEo0m/CcAr0JjN0X61I3ELK/2SWTAoKl6XYtuoDbsDqP
Tgvqh1yY/JVlAprT6IXrwpmAoZl+Zd48I2TID0iRzpz2KugWLkGaaWBqmDzsUed6
Q5A3PqoDNbJXn4neXTAum4nAONPsl/UUluWXrQeQmPTojlGdV2TFIhTpNMvysnIP
fAXBN8v5K+mMRYelWsEZUZzW58JxyyV+fA0a9kNLraC8Ld1ft2IvjOuYzhKwPMHL
j0XvB4DEoT9c1XdFqIP8QQLXOy1McrYvPHzvic/arKKyTqw4mzkBH9HuyZRj75M3
UB3P+MVLwYgVAaZruPpDn2x06HFHzFwmWJIG+v8luybJBlaeuVt80nSWiuaPB6S+
mE1pihstc5eCiAT/EUJT+QKzq6MIv8wzNYLTBmGZTUZjKW3B5iq7zsoDICg/wer4
NmyNxKmsmyqtWMqVVkCiiPwBc+29758SdHT059r2mYRyg1JD0MDR+vmI8Lexrqa8
AcCeh0KuTZwTn1PbQckgvIlr3nly6FNYR0ESSIxWVkZOefMgR1+AKDgWkESjBAmF
MvjwpguQ1LyKEiklyGCvZONRni243kvacUImI9aDsa+bI4icwazhSeNjUtvKbzZJ
jGG4OSUK6pU6SgebbaEf1j5wUh7ZI8iF6KebiDufDMlOkKoCB6Utw4gYh6Tz1UN6
E/xlSKWPlsx2/7/6tXhhsu6l8GXHVBo4LwS+xGUPaLXYf74IXdd5XljtX9oBPLM7
QctPRy5MZ+olhobBDBqLg1C0u8q7aMfIWEQO9SZbpDAv7dFiNdNip6gXjuGJ0Cu9
OA+6e4BKFotylrDBW4MNliL8Y6M0BzE2duS6KgVWjfFvnQZtmiR9+tx+vyUdVq4F
IE4I/gkbkTUmiOxNpQMvlyb2sALAhoJFUGmZ656PQPN9xQXGiI2a/vKpFoa176t4
Mm1jK8dNgXA9l2IXfzlf+D+QvGOYVxcqJUoEDWjy4jKpJNt96EEhhD9iNv9R41BX
1xAHBYbbct6vb1tnZ3bnEKqHs8ykwnctzwit6PeBOrHImFSVG75DLsqlahhXUTpw
y/7UJMKvpzCC0Y8e9PQDh6p7gmkUjYeCB3u/wNGg0e3jbI0R5VKOZWPwKZBWCa57
c9G0ik/OKUmpuz2RJ1FNHKU1LFUrPygDZd72G35fQQ1oZCQQc9GJTfDuH4B15lhU
9pBSC4Uy+X8clD0zLghYwS0wOM1OcaAMoGu1KQMSahZkhEExA6zPUM/uANDhKLZB
KT6mmnX1fQfwlB1sAc6BLtPbAieIcrdc6phvVspy/mlHpFwyClCKKcH9sbRDySyp
WUkEeQ1HrfKMBYCseQNlDL6K7RumUuKRbbOSh+/dhnXQrhHZGyeZHMibgZvq68eQ
Ub8wG/eHDDIRxNDWDKHgS1D1SkabVxf3IbSPc+vJmcuryBhObD8ALvd52i5XWVhW
msL26YqWDvGve+wS4d9RAKL9eFB1mIKEwmSAu3TWmv8zJLr4dpy4LwePe8JR3QCZ
7mUFH5FeQPIZH0LgSDA1HjZAX+sqnC4dyMdhkFHMIXsCCGFgJC0xre+RCwVO4pgF
gy/2KqgLctSHEw0FSU8SkLBuGhYEVjZRZ919rV2+a5Gl/Xp45xuXcZI1KGdJbOR4
z8l7DcGz/ks4Xx1jcYQIxpkADaUwdoXG2ic5gDiW2wTDYUPD5bdlmyPc/8XAW+uW
MwsH15J1gMthGULnC+Yxeu/WtOmVN0YYtWvGXiLrVE+0kKjpsDVwNNQtVigPwN8D
v+3KASC+zBG+aSkKnywJp4LhUuYyre/UWpxLTDzOkEOgB44Wv6vktANi2HKrrOvK
zTPm34t0oMbAQt4QlaKA63V8d/qXtdgjH6yvQCljMkldFhlnqysHRJjR6sBsYxIt
Yemi9U5REJd7ArIT5Xh6xoy/e0xbhEEBfoNS1lYdLwiyMX7elApr0bbIE0+u1bnc
vIAUYaoYPyvlT0R0vfA/XDlc0IUQzg89QEs9a/CJJfp6TPOjI0dBNcNH5bqoIQrU
Lnkr5wQoEcLf7V5rOJmKutWmLFycQ/tdaTviCFTKaxsvKj+fJsOj0eJP9iiIMq2a
IFpOk8jxCBjf6+5N5k0UrOPpUAv6aqghOQcM9FDJuiTYwhUpZylj0kEMbQTRgpBF
m8Xr1AdK3e1k6AdChEt9amS9IOsZyGGadOeWzJX1Ie0BYd8uimL/vnilujJaDHRI
WBrcqTCaHMlPpGV3UtR4qIpfg2lWUhsE1Nl7WHAcilB+aF+TkeVkkys5XJjJBr5U
3JqJvqj8XnJnbm9cEI5oIE++dRX2wDFIkpMWu+qnpLe+ffVspAFI0pkAa25zd2rl
NbR+xVnSGdhPwvRLGXYKhTtG2+K3Kl5X5ohCjPOZVPRBfIzZ0wGnFWTqdItzJgeG
r2xlNpNRTm+NB4lmmrMBcSNIclzFjZexvhAE41lsMS1cU8TZgMNVAjlvLb3J2/l3
8pQwdVs2tdK+FZfMsLRztpDvdz8SFnMsLfyWyTP4z0yBWpeE14+kJj8F22OwH8fA
2PIsOUlvzLdKvNx82BMNwU8p0NOoew+vBuDv8zQJ2d2uDs6gQLRtgPLTqLPD8dQP
bct8Q5FFvSsSIm4Js/tulzBlzIrrJZu42ejBD+icOIinXHmESL1I9jcP3+ATLP5F
mRvN0W4qbSUSA81DM2i+dWheuGHa2OWuMje5mgqqROkkMmbUeQIyhGsRfQwawW4s
ek8BEraHy4OHNq5Sj9CXK8CGbDtMrS5HLsqi6XfaXZcd6HT+roFwgxNXIbIBqLd7
4BnRccHVDhS5DR+oU3nh1qKlmy1btOMrRqLcvJ/2RSwDpPtYuWZfuNPMAxUrbQmb
gjkmnChHosHZZY9FXkraRy7eFfOU937gFiRYmwiZWqsjdQyE4IO4Y8PYt0J+9dUw
NbcnyhGj9FQRuYaEh8uByIDp2yc/x7NMO/YYGwYyf+WtXxIw92SIE/IhxJQLvftR
ZksuKZ8DEq8qd9FrsaBDgeya03XOAqffR3FZPdDI7Zanqm6t3of5ZZb4gz7bO8Rw
HNaQR2Jp9T1BTrFA0i+K9Mqvv9HC8pHgBmDyd57/vaXMkJSHeKsWYRkC+tZMxKJo
rzABtuHCbjjynApRKr/Cc58kaDXn6QXI7E9vDW2rJq9z4DqzzPt/8f4wCiUZuFJc
Buf7QJU13cVlPPwj5UfFSWBo4A71I6/285QcWbp3Eb0ljUBBNQd9x23sUBQOASCQ
ej2Vp27tDqvGZmtc6iDjGDOlMckd5FYuQrcMapdFusQPp9OzXmtwwls+Kfih7MvE
PFR8PmiXfUTICHI4QYVwRGM+UvfT4DK7B8pqfcSo/dIyf0mf2NY4WAlq2cQnYWMS
gefEbOBLaHUB6GHh/0e0AdqNWd7wEs6uUeEfkl5FWW5WM+MWiC7QfpcwtfhaZzXP
IgvVoj/O329fYWTP31Kz0icoSgbOq5Aj052/peapw9KwyEvCoy1KRDvVLz8LjmbI
TTiF1drz+Pc8i/cj2qhSr323nqXcmf2eH2EsL0CREXabPPpnd549PQixDaEFaZKK
L0NZPeEsIKdIk98En0/0j9LtJYUG23ZQXaGMJ1DXUjEDF0tkbYS8npUxJE2MwmPU
DoR0RacHUh3IsJ6Ci5QvwJqWHhul9jRzl4eozeX+2Tw+IdUlrUTcKW0NmCDGkBc4
uQn6RWztc3tC+X21f/Qdy0rnAN0XUfnIKzbWfv0AlEijxo6vcYy79oW9mPT+NHiO
ZHk58qgnhxF8bwj+1PXSdbAu0ZVEGAveYZ5HquNqxS9JDFtQLnZGuGWS4O/K9rjx
BjLzjsyTgXrB3ImO6yhBM4A1bF80iDb0Cyb7B/LKLzz6AzVcz0NC03dl4U3QG8Rm
2TjK0eE2uduDctNs2OrS9YSslymRyDZVmtPHJHoqgTmYg5AwSAYDC5kuGVnnYYZy
pgXDv7107dumEIxOWpYHw7dYRBk4gu4OAzP/mwctV3o0VvB1ljbrxwlXQtPfb3mW
Q4G3bJv0vwM9+Go1+Vw5sqrdJcKCEBZOz1p/3O+f8zBQ8eIC/pbdmO1KyuwVW2+J
xwpqVEb4os6Uk8+I32ffBuclq02irCNG5r7bLfxUsBPwVsItuvuhOyNfcYhmhCn/
EmRQBjjf9gyXk5cRN27b9LOXk1UHrJcOiRRcI3c4nimx5iRTbRYyR2wFefw9qClY
fAWwT8H0iWxsI1CGTJP9FkmpHhh7gOdVzp26dI2bA2OtPi5f3W0ykSvqBodWbdH4
hOLKyyJpUXYjhmO4tMVzdLWfqLYrpUVJ5XpblaZIm5iHgdULWYA827suyRyntFDF
x3PshR1aIF79V+Mds24oWit8izZbtzj2f7hzTWJ3HY+WVi7RlRmMFjvRTXaAlPxu
9nPHscFMCoQ65AXj1MxSL746lJ33OAosUAPVItXP4UpoduLZ5dqgETnFPxhujz8P
SLsTfXFt1RSaIS8tsLZ8Mo7zFnQqex/vmrSKTz42AvPHvsHbW1qZpJ7fgzktAuB/
WxeYvFEbE4I0D8DT/gbjayz4IJKQ/TAGnIiB7ncEf/7jnYx6qFjg+pSdNvaDjFYw
8gctAnKHp1LGCVA4cStHZzIxS2MA6A1lY7P0kNALbawLYxmIDQ7lz5nkdprGeHer
BCTbXuROAc5bORNvGvxtEdMrxkoAVtCZxFSEtlTSnNjkpYsTUdUu7FGEYehV8OyT
1bTopgrPEttFjd7gqwowqduboao3liBfKGYNMxPgbf5JUxFlSpd7tkD0OzR/IaIs
YmRNq2DlLpAABNmES7az1yKd52sC1EbYA7ufBZlSFf5TMtLfY/CDncvQMzamF2Cb
txP/0Mv8YT7MMFKPqx+bIwPByCxdoM4rca2HGrcPvVMZ+FzITrVrKQHdALJWN6S7
DJcLzSp9QPNXI9NFbD7SOF3bXsyJZFhiooDu8NkX7n2hVkvkzf9WxlZj+Pgn0bBf
q3jGYBHuDXuD97Z03hMg6L7yd/LOZKfMNXlpH7e2LIJNkueA0Wxq3/yMu0+NdAMq
+mB61MFMUNSGnIQzBRuzfBs3OCwt72Q55MwA2Nho8UnnG6T2+VmlXisrzstRyjZc
3jcjMr2oz7MHO1YYTAVq8h7r/W9wnv5W/R4PEdDjLVm+3GZOIJwvBty3/uzhXw4M
y9O3/tiSf8XTomyis8WoJaBdmVxQYUX8i7isaZep5BKjrMyJKQUaT8EsG9LTYWn9
0p9srQmwmMU+pFEqo7W9pDPOg51yCUpwYK6rVorITSYCgRpVrAp4PgCzBB7SMOFK
txnKzMBsAILaR/vnp7WVmBy+qKKSHrvpcCcMm+KuBq9LpqhssQI2hIs2lNULs/uV
OGg5RI/0VND59B5W2Z/4nNz7cyo3jOK35KzHMubAdeh8MBgFLsGsit4m/d3HV3Tf
5S7YnEMaa3VmZVipdYhW2n6mOxd2lZbI8gaicoIk22QTG8QmOrDkihfZJul23X/e
woFt8nRTPM+4LY8Dwp6K5u4GwwOPetgQDLgXIqSMsN0UujkZmZVEqz8PmwO3lnQR
yzs7LQl6BAFO0VNcacgiMgtgnnV3EpzMIlMpcQYRjLqa/CeflFbS6E8HPP4yagaK
2WSsZ7NmHoYj58tB2RrmFw4jTdbXCnmBV27/1b2xk6nPt9R1thyhtisT4BePIrWr
3aOj/gs0ooL1PaMQXhImwd1IupE9gAirYVm2eSfDNLn2oCzEIiXocvb6SMHHVa8L
`pragma protect end_protected
