// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jXQm3BrKOThxZItjjH6ta96cIDuQfHLNPFPOCA/Jph8qpd4yCEsLCfLARINw4Ry4
K93qjmL2ge5X3LnXRcM+I0jvEUEQFmellA6qi0kPs4c8e1bCxuXU18ipYHMr3NMY
W1qrRtN9rCiUU6DhDYavGZ1D61NYsIwm8lDAAmkTxrY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48288)
0NOQnyMumCXE+5X+778Sn+w2ovjsh7fCgksYJUyiN4uRULdwObqfnQtAQ6l15wfQ
GbxO4vX4kYK0HS/ipwAZ6ifmXz6sygcA6q1GfGiOvmSg8ErTHgW08NNcBrWRuG07
oPoXK+40o60MuK7Ohaj+frWedICp8c5FD+xtndF1/aM8lj2pFbSJeP8UPp++n5Uh
xmhpeOPCTswxF00pdn9yKOPy8fzOwDBt85GY5Uvhlbn3c8QCuFGyEipgKqOI6bxF
bR+Lx2UWHSFD9rAROuRJxeD8hTwQhkQmZUEOVi2HwgR+MpsJzrShADANafgUfg6U
IgWPK49vZ9I9YMqqFvTM4sxaxGX+/hA33BpQWWlW5tEzF2A+TF5xK10uKEPRj6Mz
SL9acKRQKg1AeE1HZv4PPWA80EBiA2a01T9wcgd/DbFikZInjOKqQ1XEiuhyD6QI
vVAv8yTo1PAv+3YJmZkMxRFaGW9ThmrxVoa5wYQfMrTQMqrESsZQr9IFrXLcctK2
MZx9CPCWhVUGWDY2J06fjxlXHUqgijvkZcpgWwbbkjk0pzEGpI3ppb3X+0JJvtPL
OP6mWojF2xpwS7WuDE4KiQFQOeh/hq01LD9AkKSQLOPDsuO7RjN6XmN4NUF49cqC
zoAqpDGc/Nz8K0IlqT0TbnAZ3fiODh7MFGTNT9o8sEh4rryyfMhLvcivQh/6yZ/x
RpH9Ld5dhFMjy37+7rRkvY/CGGI1UglFkJ70HmAaXTqaPiFLhf57pteuKr1Nbgf4
4U8b78llAO2C7cUdROvGUMtgbWa4uMP/vuzt3eJbulZNTsCD9hvYRVXf8XqOFZ/O
jhRxfsqbA15EloGqrhfCrykAE4CcuLZg6OZp0fqKj1c89EQ7g7cNE7F1YZOFeq0o
5FwACr7vpVJ5WXBlHYB5eKMaZCgZm7kKtU4a594dUji7bEaKIsJPged1rsgEm/Li
tP//L2Te0mCcg1h9ZRGiFMINz9pnISBw8M1AS2RtZ16LjXbOITrhuBqWcaIwGSdt
zjyUjEjr87RK2Z5eZQN3pXjtrSrWBrokNPaURSUH0XG7VMFX5S6jarP9YSo6VAgU
3OIdMzOHqHnPaDEBjHBR3mEPneCu3KylzDafIlNoqsmCqF5Q8tXiC6g3ot1ZxW5H
dze/yHPOrC8dp3ppexwWpkV6yIf0+akqAeqehGwV9aEdUP0ZJSGw2pkwubZR3NdO
s1XuCfL6HT6DnryOq4pgfJFGhLxj/SkH4gxc2f3utyQaOlfFQJAuKm6I9jCz99le
tLJxMFMoRVMy6omYwViEM/eojn8m10RbhbZ/+7aBIBaW5zFBdlCm2PX/I2DsTynl
1+bv3aSoz66XgBTKBRH2w2aMoxWL7A9IRZY7ymQL9ZaZtRPEtab5U1XOki2CRvYv
t4HoyGLCvyb0YOoba9dSBGlL+L/4aHxYK8wENghn87NPmdM6bBiHXs4643H3+gEB
buDazMtKdqDKJRifclnOsylt/zhrQJ0VAlC6GVL2ZB1ON1pvNABcEqHsh+OLM0j/
kG+2uvTElnZS6Ale7bc+vgPFUx5x2ECVCLaI2hnxKbgKtgp7RBzVmlsjR4eYIvf3
5wD4H9V3xbM05KIQOEdpEe4182Tt05QyCxnBk1l6bIp/tUffBX+lrB8BAkdQR8cw
N9f7mvNKDIDhQTnM+ROGWKKH+ZCwM9J3ANMrJ85uBhop7vDwCd7GuA1QEhPcHHHy
+z5nNY11yfMHeM4VZ4syTK4sK60UAP7b0UCRnHl1gJe7Yc+Ouq1uFaKahu+4oFeu
EVodjhoQHHCJ3AnQyG2sJET96PraAflY3NLxD+oe+Ryp6jTBubmug6HPRns/6ufa
oDUnN+s75KDi/KqQJTulaKW0FRzodYCK4+Q63lpvQzKwBXxGSaM9fPqzpB3iceAe
9uo0ldFqaze0VMnuEA1VVbAxSm5dgwPN/R/ZS99rnAyEMuUBhigVf/4qAJuibzQ3
fDmQYAxXUC+fkvomzJBamWRXCb0s6eqBiUJn8sF8j7QCWO0FexQCrZ9LbSSNNeif
o9fOx7PDZoWs/HX6qGw5Z+vSlBozCPJR76UUd6L+ELVcEgc33rQ9rzGg3aee8cFF
INtLkYu/XdUG71M54RNFzQdctI82iqMX/e0CAnwrDsxjS7n2nhD766GyR3N5imqM
DOc7Jt4DgWCVVhMhVogD6VLh2gsDbSSPh4EOpjxLRlXGVFv9VxLFcUEQDcys5NSq
+1a5yZEo8fBMhiGkqMoZxI8AgIme+A9SM4nK7PRMO2Abz+eVSK+gityzOx50OUln
ZJn3SitV0OUwQg5iEN0H4MxIC+2uLS/rHVyz5jmoshv/YF8sCxRWAH0RTvOfIZ6W
R7ag1aFxKrOccTuJFVGq4VaCL+/8JRDpEkpzZEMV+iE1JNbMh6CyQVaD/V1su0hy
tyap9HSDnrOii4PVdkqDiKbIA9c3yDg19FBPZ5q/GNMM7NDGX4gedfPFg7OFy/nC
HqU4OocDJi4ihUrjaO7xRTKjV8aM+a4Bc2E68XRzwmOIFV7P53mWfQfMsKjsIU58
5rwV1faAOacbdS8AwWOlnCde079fJ1a3S7HlsClQVn2GA5xe+LmYox7zhWzsCW+t
iugjvGcslR3ZxwbbKgQ8xG+xYAYDjjNJ6n+bYr9fyZyUNxYi6HfKzNcbZz1bK/V+
yfpCLvK+D7yfXJqzz47hy34Eudg3Lv7DkUPLGwu80YY7/UPT7vogFxJNBPwHvsby
nXOnhIO9WZtog/jVCVL+dh+FvLKTvntHuhsVEH30hbOvx7qkWSQabyRJ6MJXsml2
cpyyTmgGnC5p3C6fre4/SuWqeTHwHo64SnW87OTGuha+CDalu5fr/UjUhn8A8eAr
M2hnmYX9xjHoRGQ8pwZmK6bUwvDcyrXAt0rHqbcXtio33evf0JhTreTkU2MKrLKA
62iZbwGpN/UOka3KalDt6vIuxgbI8jkU7LoYLl87x99y14DAwUZUPrfvNtXWlUws
GgPd+MZFrM5nJtRjJnNpmDdsJAgLwHM5ZmJbyy2HilYibemm4yq24BjGhWIOc/ix
IceU5WEl6B2eINX2k11/94k83ppNKSGYgLrUBD+o3TQWjC5lTPo1yr/5QxXQoPt1
HVmfTgaEvlzOs/RXq+uu2GlQLEEe+PYOaaLgnwAC1uVV03AMNFiVGeOty3KvvZJf
jMaMbzYtZIfXdHEoBymZFGMHIFjFp4oGx4ysXZ0jeei3GSegwOCOPoAsZDMpYvwh
VthyX3gHGNsprXI/s75Q5+fLtv4rxlQEnTtl5fmANP7M1uFJe8UfARUyHtNfdm+W
3au+sSABMQnplmeHp/UnUSSAZBkLUgGebDbo1vV6HfAQTbirzJUXveyhC38vOHmF
KoLfuYgDXC0veeUuaUek6KHYEAboIn8575ZFpxeC+gWn/rGebpyD97CsfVO746pL
myy3/Ov8GVsBPl971IPphW/Mqoa8QhTqjb5PUOL/SjDnSuiUCPPasklHeWgB2oxQ
KKoR2Xi6rkPwzbmsVg1tX53Vg68zUMnBUYq/bKG1gDrvrNBWLgFhGWfk4tHXExOy
+JTyC+J0fubMWN9C9xmUf2qc8USHENdNmckXHqdRK2aGa46ycI3OUiR/u2VO7ZOb
0tyec71ihdfsJyr0toFWByTRQBR0IzwpRTojJZlPl05R/kOCIyUVygjlxo4VJfHW
X+xHUL7LZ6Qk6d+ct5k6J12Q4XBKf+9iO0RvhnjG5NJfI4ICZYIEOmFwJKtKJhBG
oizgVPVYipuZ8h5NDoH1s8UZvgzQGKlj7+q9nF7Ib/74f4AcYBRojDwL+1Ay7WrN
+l94xSUTopiHGY4/TCCOIfGeuMU0mHVhC9rfT+c3xXPJkWoSdZrr94kYeUJ6CDgU
K9pbeYi0CyJlCnp57M02XB9N3RHx3M6iOyw4Dew6tr7KcpJvP8Ektmp6V0CFfqm+
05Aw2tHCzuEVsTcPYJPH8NWRcOYXwGTy2xpzcDgeZLrLveDhmEKATJ7Nf7nk691A
siuWpS3raOGpgfrT2fqbc8S6doEh8NyuDUK/5DCxUsgGI8VRFg94ffSuSIZh2C+5
AoVNL1GYDaPxdwY+bn53yOhvwaVOwPbt/T7wCeRDBT/qSNrUYAIFEfMQeD7Y3fE5
1rHumK5YkNWRWphgCeJltc29/q4iMkZii7bmqBO1io9SIqbyb5Zfo19khujBHhOj
qcxKHD7jFGlON00RV3mmNhX2W3PFKFnhHgp78ThrE51DbkMFpQeCE8UPWaS9epv7
/atK8Asi5Kf+GVMz9dSaty1oX5sU+BuGeIaM6tO+e0+f+AR4Eadl2z0/78q6A3hS
+XBpSWujExJcyTSAEyqvEMBep43Huv/ShLWmIIbzqs81XDJU6hjnoldOu8qUuaq5
V5q4/um6u82Ei/Ad6/UchHi01VJK5Nyb4gFCIKjm6Oq2NiOXHDW9GHBv/H70Ue+Y
AL8FHiyX1OwYlnchZT2fAsNyqicOQOZqj6CJn7XODnyXe6xQwJWUOP5qn8HjQBlS
JRr5Y8qY60x4z/ZFTN5m56Ks3qjQ+6lW+OGQLMUXcHLeKKcGxTc/0PguA4b/vJRe
NeYFQJR8eQOKvnZrgIu6HWvELXHcQPgZDSYn5khx6hue+YCke/+6lNDTw1hMQoH9
ZG1mJ4+pyT8BqLjdm3yR8eVAIox31aoe7vrI0n8oK2NzmMrNBYaTYkmsT70EmXy+
bbDnBE6WSS3HJuRo9Lk0tvjB+lytolMVWWPV55BkofSo+J5l3dKh3AApdCKVRNbP
b+BAsCWF14GgYL3wmoVpwjx47tjS5CTP5U6E9J/j/lUpK+lwJwjgXD492S00KxaR
vEhuqZTv/L2U+iWitQ9t/BXGIEdssvA/IXFQ7YAVUAz6d7oQw4dQpAUhSIRdlN2m
vWftcXXONeczBqcg1TLcJlfFlGCc4X2rw0WeVJR51FxQMoEYCX9PT7Z9GTkcmaof
gKE+3oqz+dVG6WL2FKhmHaVAFcdcwZ6HPA5du67dc3vUJcBV927WwQteRAJQR+QU
uDBiFbxzV+FK/Bbk43xOJrPt2p5bbff6YBhIrp0oVvXRw387bNwRSd6h/82WwnDu
38AocxrL00xUNYGRUhjbKqFQGTGpDSFtj6r1vHJ74TppCO18GhEAKerbB1RJAUPL
BooZm2ejKEakwxprB13IG1WI4Kq0RPrhbMDQpOZcHz127/n0xgwflqgjR9DTPfp1
jjBoTxfaGZJ2+oi3/4FU2UggjcT99yyXNjtPRiNB1BC2jgZdLmfnDRF/qO6VggmE
AutfioEjezNCZFRtQwcsQxa4fFsmR8wkTd1nHx7jKbOpru9tHSISJcVuBJRVKTIN
l7anJ3qFr+VLH5hikMPrMsRRcjkYcsLWsXeoZE8L4iDZyVgmtZDRr/yz8h4ipWC5
ecod1/e07aiShP5gxVXvUTfIcn7dmywzVAUmaB8t0y4GZ7OVm+zJzeJ1CoNAECFZ
k9AHETmwMNHZvZRZ8F6W7eAhqXOqUmFhH7sgnX1AFe4wgbyWaq7k1Z9EoSJb++NB
nM99RiEIA+l9h9gwTQAucSk4KKW8sm3EbdYIPV9Eb/G/9NkD8ad1UkOFcuo4rKw1
1T1jmTKzQwHqa2VGAI+J74FhiQ2b71IUOD0Waxb127adm/wzRr9Ms+5tzjwUVU5C
I8Aus+nJzIarp4Zh25D3ECSen/6ptGcQDn0PB4D2zKlAy6hH7zkAyi7FznKcHkbl
wZVati3oAsJQ/kDVz0mutpi53Uj92VQiNvZQgNcdDCTL3By1b6vEMRstXHoeV3Ub
upZH0weI4AZN2jWEalHAuURlPqSdRXu94kpf5KoNU43jc+p1lEUxBQeuZxvLbaMk
ExGy1xLOivQGClfvTBvaQgY74w2wbpzt32zr3UOzHt8frtGw73wJzCZdmiBMYPSi
8f0+PPA0Sr93U23scRQkq+WNwFdGat+GdJM3/Sna5QwEJxMaMAAjdBUslLlg6Jru
AwST51i1Nx9dmQG+psFLaC77HXI+oiP7q9UGSSzp1tRWxg3RgCUH3ViYkRbsNJZ/
X+wPsWONpfpc+zwgIXS/Lprqv3lSfqLCibseJ21sV3+FS9xOjkkUeWGXNdZAxhfA
1H0oce0asZB1kjUcERHew3EoDo6doQYbsRY9GDIe22pYTSG2T7nv8RkUdvY995oH
6MXpWumqhh3FU77yaUN6X6cA5v6UG3HfGA7TJxhjGmjGDci8b8VKaM6oRGfHj36e
pQKnT44P9P+wwB+sHCaDFDkvZsMZCp8povpcHprb7zWRsATrnhc9lGYYCDFFvNEE
HsqLQg0LlvmOk6S9wnl898m6ItcN6FGVVeDRzhZG+LHSeoC0dLnrH/qtagCJyW6d
Rwp0j1Sir6v0TZAs20xpMPO8WtNivT62Qpj+k0AFLrG0WI3Sio34jX52ghTLol4J
R9qDOC2rlsgxwh7KQpirduEPYv/fxyU2MWf6DCIrUrlLx/pi0TJAiZPr6+O/iMBC
POKtRpxBsTVItyzEMdglF0e2DjrTsiy5uv8XkjF6eOtUvMYGU0F2GSKMOfIisC4R
Dz/ooRRlcjjDkiDIFHKzlB1MU9sKZAt1w/d6czq2u3lPFH/tLUekEzSnkJ5CGzhb
wQRAFXsH/vsVhMPrJBP+YlY4kCP0L0eul6zGKg5rkTUj4BafBAITr6xTvVef5JUs
cI6OqWuhI1o9S8HEMkNj/c49LPAMrnSFo5HB7fsBDhTRpshLvrJPnGOyP6pb09ep
TL3TyNh1NHxv6cm0Vr212DY2xBE2CvT9qmBvsPKi6IgqP53dZc17Sq+JZyRzc8IC
XiICgKmSChhiwxtLVlYyxWeAr5TYfr5xYgpQ5DuTLxE9I3kUZNralhGGFihZ68JV
mzGQPdPDN01f4WW7ksHmIz51mRK9UvausYH8XnBAtn6V+z6w5mfko9TUE8MgRzOg
v5VEAiFjoCk4Rmc3VPk+jfBAQ42gLZXHq1HDjkL1uN2BPUXCGXYAf6/fZS5Max29
8Nvz53kJES3YCnsMx1O0NCoZHOUe8PFUWwrO0jD1ftAKWLXJIfXhMTG53rpx6QM9
ENEPAGSXF3C0bqE2CG6FtBIOpgyU5Ru6wWU5eK78VCTZwIcqbJ2dLZr9VttH4WLA
NrUDBgO/2+2lGPXnNesznBgBsdlAuidlz9vhozs6DPuAXswUmqu/mcIFikYKCtfT
kbJMajqTLfnj49Mvxy59Gvpa6svlr0qhIVW9gEw6GotqIm8BqUjZCbcGSUoYVihI
10a04B/OuI3UStzChgOQfi3eB5NxiMJrriY3TyI4OsgRUTa++JtnNxGpnTMdJ6NR
UuKDgj8PheSjZfy3mu6JlfQvrlKAWiqVjKfXDif36326lUL8CA8gO7cdbgRnGWLq
NoAfUBN0Ufdq8bSsO7z1pOAnZ4VH1y5hggsNmeuKl09N/YMIvHL+FB9WZim1qyHt
iDuCd5hSl9NQWSj0JjkhlRWI+f4plwqBzIC/SqKBzrLPLQHeP/jUxq9mborLhSYW
EJzZS9//17DtA3rF0MW6ycBkx1IR3Xujz4G+kRfqg1NeQ/p262ZUCGFBQ4e190j1
JqEU+ZaawlcYgD/jYNpNvY5cBS/h2obA9nXC+gALHwKKgLKH1BXENb/rtntQ4yEq
6OgQdmFkH8yWxjD5ts2BkJBo+zBuHanfhI3u6dmKJeGyl0wl+VM8eAP+7uJeCok4
xGKOQO4XQ1a8z94sa5MQf9scUMgPu6+Y9e9zs28G3vFuJiAZ4FQHkyQpOlE6BB9Z
h893+EkFOPz+Kpq8ycb7mspx7MyIl9JaB0v+bYOskhciKGIlv87UPP0kCnVfP0Wu
UqUd7/yOG+tuFMG8h1itI+h/DkmEU8JR225DHJEeOFDJr2AEfje80yy/gFifJZsn
jqT4NxH4rr7/+yRnc4MvV2ZdCxcGP06x1Z1tbQFYgsmpPmPmA72uJQApF4l557fK
6Ld/gFU3mJW1Rlklg1+Ps4tbSy03d7Rcr6Bnb6DgE6nWx4cxhPnMOJ/rQCKautXA
pWp5btO7NoUAH2jHlXpkxB7Bk7jukf0FXx2EoSe2TrhsGgcsevz1fwDfM8nH/4Wx
zXoFQ/lj9FB0OSt/n+3sp14RS7sMj55xQjqzadmGaSJGNrqX6VURc+E/0HTDyzJ3
epx5mv/qIoAhKVu4oqCWrZGEKzCieAoe6k2tacRuvrZqkfhCVfkYXU9idJW6sa2c
a9YuM6hY5MXdO99KXOLAYosC87HF+x/YrI39jSqOAnacWSTPS294qG4MuUHfMxRd
NlpSEZjbDu6KJcCVdm1vSwM6QPDRYoRl3lF8Yq8xbwfQMiw/wjEWUiXPpXaG9RrE
80xYBXXcYI/qNfhGG868q0iMw4XPW0IR0/gYMs3JsrLF7M5AwMwuheoTM3qXbFb/
RoX2cagJWId5hqO83yjJvqQK4OvXS6dX1Wjfnf3hXD6SOxbE1vHrO9fxWFV3R2uh
V4KwTL7WF0wB03Y4Q+k3VWEMFgXA9ADo2AgGsSKMOgFGziUB9e7nd3K/mQEU2876
86Z3oqg1a216WE9iHxvl6l3fa1e8NJVJH+qcsSGVqnX5ogRCJi0G1jSM0jybrTjR
XapnoX4y3/l46ZEoLY45qig8tGaeur1h5Q86aJWu7ezEZiAbo9tc660FI+vBG5/s
63N6+Pbw6fteDEnnBoQPZME5Xde61qI9r9iUtV6xq8+4v/1YC3zSUH6cAxjaOKfH
ER0egc1jBeGpuBUROe+3MVJ0DluQEDPJwJKNfYTMdQ2QCkNhkNUbZ6XgoeIzBr6B
8Pe+a0sHexgO4JdaUHHDBgc2pvvr1yYUwegSVIMhTgexPHxD9nynCDHyFvyNuDkf
MCRnh4+8ifcp2h2maXap4THT1AeFMy7ITFkbU8k8NsLUFGNp3ilc4JYmBDmOrbF5
iAL87GJdNGvr4b4iKhwdZddl+dXvtmWQZ7/hoQv4GEy8hT57UxV2OdjZg1jMDqc1
srslPKDlP793iFQFoETh8Fvb8wdZ66VGLNiP9PXIDC9hp3h7ArVU5nZe1WWjewxB
BCwDoyiBefLyOTo7npmx0qISqxllPVphVkwWdrhlPKe3E9Fc+YJ+4axkc2I3HjEh
SWrIwkTf/kbjE75QV1LkYG6J2Fk69upyfLhdIF7vvscmVvmC42V3UzNeg1PMv2Aw
hC+LKnXIREEMVZVRCjqsK+o4oRvgeeNp1Q91jwYwSo4EUigw17FK4xLkhbecRRPG
XgL48w8lRnM9jKAAnsYAlH5oxXWcnILvWw+EO8DkRz4nziS+l2u/06NJvmbPzUcl
ayRSLMRLXX3EdlRxPCwc+cDJZt/1MwLgxekJ7hgn4Y1VVPY7p8zo5aJk98Uudqas
Ih9wP+yxQItBURZO0fljg3wzHTi0OMdBciNdCVHl8lN88osdynR829MWlxgaq0Jq
PfZYuon0mJqmSWghtsup1nU2RBwUbFpCiSCeEon91zJ+VqBAHNwF7Hn2kpquAIux
3Ova1AbMFm1V84Ku7hqRRsE2M6lobbtsLEyF/ySd1H4RQhEdForL3K2JOdcF0sKV
sf3kCvBHZMHd6d6GLaG0Vbww2udm0NRc+YVLWSCFy5x7xBzpNqj4s8eGRioHOvew
cpD/njjOF5xa8s78opgLHgxdjI3h8xvYotd0LSYbAtgtbrnqh3Bn3+C76lmkGJb4
V+BYgIRajH50l6hnKutWIYpx+M4LkMRIYHM8BEdtXOBytSXGDtdefLqsRg6WMpc1
oEAOcTvKxt6ZlK/cZq1S+Z3pIDL1mxbJTOVlC3EsKDcbBYJI22EEBtu6rFNwGw1n
k1jwWuuZjtGX11/pu4RyiTp/waVNtNLXFKUPEc0hWNaCzYcTshkEm+7QWYDuzCZA
pa0q6XbzquWyEvd6tAqmfVvw4ID8PGSehEISatamOZ5hSU994BLgl6HLOhSf8TpW
PcwmPbQ9Wyb4tZqWltdsK9XCUerBbpA4HpllRkIVH47I0WT66tz8rl4sDuypyJXk
edMwxy77TKQqwU+KmT+/OxuopbQMpyRSXYYetAsa09RdPIANMMZ/G8ZbyeuBBjvz
hrWSo08RF9i8FpdVmszaPbWR6nD0vciVj921Fb87tSre34T20qXTWcJyNkKbaT23
zXBKM4x0/bzVG+ZKld6YOnfTH/UxbRL1URon7QhUhFELEyS/lb6RbBsOlqcmoGvx
k0eBKxSmxBAqpTsLDLZCL6zm0ft4hEQwLxSzgJImBkdE6Iv61JyZxkhv8AJHMBS2
4JqOrF21aY/iqY1V6BpccAfCPeHGTfWfYdfLGOrmvTgSmA+0Uajw+uAm+DmDVLCi
GAOJcsUMMoqfOqI3fAn6kMsABI68wA+bhM/Onkk/Uj8s3emV44YxkKgBzQshzQqT
v3CEZqHmWxMuV0y/bLiIHThHLd6lGNg+stUAVpEMBJsaNwUKJOWvJqDl4iamqMW9
lNXWPWTEUtRn65t7fzlGQW5BfeHF/4pTpSICkZTpJC3N9+aw/xXNZlZKjtPZeUkQ
og1nK0dKvWGv1ONOL2MYJm81V1kIlsQ9wsU7DO1f5zMEaVa1rujWeA5kjIpqX4s8
9GD6Rkcy4WDvZwvYhHBQjP+1TiLWsOATCTDs6q1swATggmkkT63p4hl4U3HUTDKT
lpTJgeyO0HlarlY2RzqBCuHnrdeLPvAyMIb/kIsrN1YoPmKTPQ7wYtToXw/OUeVX
pEpqlQUYC4eEKZIBzQ8vo0wkzOSUEEqkRcqsZt/CtRs3g3W2xzFJD7F5+jgk6o3s
baDm6VysbqishZ6feXtd7EMl9Q1eiO+ZJSNbPzuTGQlvq1O9YxnJYVQHuGdxLxbM
1jW0RAbhBPFhqNFHoBotMeY3uLQm0zu3NlGLoCPZKzeUi4h/SOcZt8scDSL/Cf7G
8/mA1w4UF8if2mGfqD8LKazQPg+LC3wTM5eGdvDiV8MNT4LIFE78LKAJudHltF4o
RTLn7Xxpumgd9nhtD7ZCzJ+i/XEfebIXj07KIhJ6ur933EpSnuv7b57X6hznW3pU
h0ejVOGUfBTsrBQNqJ+UiyU3llerz0cAQ2RLzvcbrPbhzYBLMaBWdsoA466xTLH0
M1sUO59yVjCPsVlMmPtsylu520hSYBZTcoCXdRZFgPsx7i/fKDU+7WsGVky/shXO
TMabHBuOWx3fa0d5igzlL2srnT2HowE4oyBgyFHN+0/l8qC4ULDyMPlkD+X65N9p
KqlWVaxk3YIJZKkfgAm2jUEKT3/RCIl7RIuUArlTZMiAUhatXK1SNkLDsmwXTsZE
T9Yh1lND39lxRIE9LPQKPEBhsm0htuY7gYnG6Rk/uvwhtWEUWpAJAiex1EqPg94+
boTOYzFSFxzMcIMMdZF2v7x/p59hDNZ5HBfzg7MOGoeo8GRDPSx8+HlRK3LPurHM
dOsKIFM7WPVRtADSfrDs1/B4iPuxXUJ5Xl5eG6faYFgW+MzEc+Q4lcIwHiIuT/3P
2oQc8q3LFHfoUKMHqLkpg/ILXethdVCwyqo7Hxih6HQeZVzV9ekaX4+SgvViP7be
X36BpXKOwVR+n6itBOKt9AQxm36bdQPhQi4V8FXliUGLZRUsNhOlb/BLL467V949
ILL8G8qB+YIPxqIAJD7lylA47O0YoLKO1giJR7fXjQBhZnw1HAE4EvgrVjomcMDX
UIewEuufs6xR0CG9fQB0cswJBvX9czuR8/mVpSiX5Hs4LTZJNsE95wTJu9j2Ah26
+HRfN5Q5r9IzGhqlD9bRszf56CaWoTnM8cea+//PTqylav9ajl9MBodzkv2xVPnm
Mr0JsZcSwj/UDyLMRO3Dfk6Eo2Ctgw/yPCybF2mJraMBBBCgOpvEAiOsAHbabcty
wedcCFXXwvBkj8rTvow1UnY4BEW874sm84K3Nr0CLCAPHK66D+QJhMaaU+9mdy3x
uXTkA+i+QwpixHk0gGj2SO/RHBGFwckUo8hy0P/PZ3A63JPTuXMqbHuR+rOmepMv
wYVgp+2CITNzieyCstIEed7m7HmimC4OgOxMfiIHHdaSjc65Ta6HbFlpbYgXUivk
qNygQkzkW77/+rpJSCsyyF4enkcgkVm0zn2g4Tl6mKT8PKV5e8lrwg0v4CKxcsBu
bP9Hdh+dO0mHCGqgAhCjLb+UvmhYow5eCOZWNiVQ/W/QHRJnq2qMVvVN9Hn+6fnG
iZULi2KESh56aNbriK/o3TYrAPZLOt7l9I27KTxDooiOCosX3kOYA6CLcQSnSJH2
15fcVau/w9pk3EwJz9NpZdKip1OALDEVgKCbAb4IxyFmMjtartZLEBZQBsy7HvR/
cdeJyzqTpGBWnGJCte2qL2qS1N7Z0Brgo0Pv3adHiKM2hJCov/utb4TWcgyOvr9R
yA/uw6CCzisqRcb52nTkwFH2GczCKeophTJWaF4iegiBZmoC25cANBDk0AH3fPhH
HR3FboO4Ooe/rpFJg4O6c7mT8aPsPecUf3cGx6Cpu7jILcWn/5qxaOX9rfQRu1d8
psivcKzmR0jx3vPMckeuYetjMmyuOdTOufud56tf77knj0PXmUSZRZlW6p2pmCps
cKmVNV6jhryuqeA+lwelhnhmv1lug6p8csyXNAOk7IZgTw7XVvV5+el0co2nZzLz
q1VhA/jk8qd2wNjbEiGzIjDTbfBUEaxx4w03Kz6VKWhXhLxzCeMghb2CJbt3A7ei
yydwa0NFyBNp+vh4BdfmSTiccBfv/ac+RF6m4OI8sWtEf7+zZPql/hmY+3XdRxYJ
NTuZ8MHKmSOw4t4j3dAIWpQ+SIFZYP/vFLhLEDUnnFk2yRAYoJ6wJwLvGNylY4Lo
/FQeyc+8bHoitRsaZJkdCkASwbsiqhdJ5kJ+7JHzy4Zt3UZf9da2+wGDCZ76eYBx
NhzhTc0ppWysB3DUmxzvl9mJACnlu+zAKjkIB8xWaIHXcBxGJA2jO29vkStUiBMn
sBBpYCUKjsOqN2MiN7FRGqgb431zrD6aVw63amaF2BXw1oU+YJX1fcVbGKuMiEB9
F1VhxYrC1kjUFVjsqsR6xaAZCemASG6eRuDtfjwgvbNXeBreIsN724aB0Mo5dP+x
buRUwmC+/ZD85DrqBjIIWMd1g6UMRfwlPraLmnolXNwf3fpNjExwuqslyiFUdUPY
G0LHo/AEEx6/VTp9LEQlyZo8SWfscWWSvhfraNhijyvXMW02+zl3HPQFtcOSa5Pe
KSWPmjq2e7xCHM6nshPC5sxsvzkPzGFQCU5Ka2ANfiqSVrrJjSUJY0FP1f6dYfAc
M2CyLpgLgd/l7WqGDUzPERY1eyPZbm/w/BqEK9v6Jq+ulmk2tb/W8mtLXHF6qCf3
IDFBlhB1cCKFgSDCnhnk0rkoTYb2nptP/hildhClT7ocYK/RCnbrM2xPGleSVvsJ
OO3nWShv9CA/0PQ/2Ut0kdoc5z7xgkkpcXFbN9Tz6Fg+OZVVJISXcHFQZsT4ffBj
01/wp9DyoyfHPi0byMmOhb7sUH/jyUJg/IGfF57TU7osnusF/zzOtJ84pnA6+HIe
YZjTOSL75/cF/jhQwYC1rdDzGCPMBocAocafjDVRdX8tI9DGaSwNBvipHqed8cUd
3BuBvxrV6p4Z5bE4NcBD4M8OGeDuN4DVj8K0fBRFa8j/EfEU5kE7jTJ3QZMpB8Nl
nw7dt/6QlRDxULZO+rcPvYgvoikIXvQo7qSpAJKU8WE9a1lOYCaegWgFXATjLAvK
mh8X0pTdeSU6w0d2/+c9ljd/w1IWzZNI3sHO9Eb253qQDVINgqgOQh05jJtrffUh
yF/InlrGl10xHkyAwbPBGqirlZyY2L73LeQPKhE6ELn25R9nw2SDVK5SoCMDRt90
jysoELC0PmEesslfDKiu8OaGARuGqi0R2vmf2xathWgRX1bwOo1abhAIvF/hoHOw
EdxMyKLFxEZO6IPC6nmDRSP2REXVIeOGtDXbKQGbcf5VEP5APbdFj0SGNcGXZOP6
wXUmnqlG6Fkp2XVmCozuIUYqGx8EUAghNFRmojn/1KpGTtFHOdF37gcDn9Rb6ZiJ
SIkdWnAaNhrAoPwDlGuUuAOWy1IUkyIjDTLlbVz9z93AoJ/mmgw+sbE0j7Jp6IPM
az8VKFbcmnLAfu+mb5ivwI/deEf8eJ9xucTVlYCBGhR10AQTVPGPXTNh5LEmt9WT
d7jRQga6cgr7THSfQDco9hWVvMVe1Q0+/xQQi0tyfdoIBb93KpB+IShdo78iGKZ8
6wNt4VnJPSz5I5jJRYorRwYmWH2jZ3ECXZQ5xIsL5N3+GE58O9OWlRI71UJ2uM1c
HQziW7z6NefCYCRjRYVSAFQnWYKScHbFLfW3XxxHrEnY9+SpZNTOG1TICiL0uKEA
Txo/I2scK7gDQEMeVj1OVuL67xLj9T8GqNOSJ+XEjDs+JVv/ZAmNE+Hce8zJ6dJY
NUsYl03dmLlSXYTgj73zyxWzQ3Z0C/x575UBMcLfm1lmqt+t0rcc0Qx2JpFN3tQT
BMo3USGrUiB1IeWS2/qnQLhrEhnaeE5jDX3qDGfTuk8o1RxACSv/MvZ8ryCCOmyz
IW3NhkIygFBrbGPtp7YtL46Hep/5ww9NjOhbWzMURthyOLpb2dVgvxaJ+vtTO7y/
bJcSnyfu2G4xxjFU92UX/dBZRD8MZS/Aslnf1IHjL03jcAfGJ3fkf44Ht9t06fU9
Pbm2T7vzlVIsqXRDHfKzvIy21vArlMkB0zE8ZCQYB7aTQarW3mWlKAdS21GMyefi
Y2vJ4zRwywCG3fiV2AoOoEPdyycukO/wWQkMvAPAOYKnJb8+SHidkB3RVu5a7F3M
N5NEL77+dxfT5vplUefYYcwxAz5viwBytGas5hkXwe9vpbzqYnuqIJClOsMi023z
YtcGHDh379YjsH+c61SWsQODLtrz0hRMymssrJ1yVHE2Wz+G4WPKlub2pf1hcpkh
RfBDgdS3ewOkgDtn2/GKngwgT7f8OG6xzYG0TiG/SPSWI8RWYD7mMNN3xU6akx6x
oAyW1diQvvYv9OizJWqu13EsXnHtz1GT0t55bcvGBGZhMEA0NgFbfPCEmL5re+if
yOWYQKhBh7vQXqFVhV/Ar/A858LbvmcsXi9m0SLEn/hVLpNVNLqmKPlKH3N7XwzZ
/SfS6VoyEmU5V2eOBE09vT2KuVU0HwTsoi+/0POiUcsUfY/B/e/vgSmIrZDYFl6a
yneMRlntEUp2LCrkRODk6sM4SSan0qoraiAD3CSfXp1SFFxlGIsRu6oISdgFwBMq
YqBKmCNXJ08fYvF9EfIohJZEmpm98Ty7qXPPku6/0LRB5eQwawCHGfNDGrZYV6Aa
bjwNE+7umcFNzQrlRwBeRdqacDEgRlsBxcRiotF++Lv/4ssJg/ciLWRrxkH8M4bD
DhLM2E1TZjhopSJFRrBpZmk3k6Zc+fiEgerCx8g5Nb02reUcXNj5ICqRCsCqzv3X
GHUiCKgn82GEpoVFbaNPpxLXPMP5kzynxakEyR9KPVEbddsHsdjs0pFaAE6And7/
GaVuNV5yYtj3T+0Z6xESaT97KMb5cFH0QmdwxGir05A5bPQWGSYw3K0+ApFqRNZC
RVmgN0JpjVofC3vYj/KaNA/8tLZJJbIHrpSJprGZ2D0hpYMuWZn4XX4v2n4Nsuih
nEVC/Cvg7vQ1aUk9zQNLb0LkXVtfL7/cHwoRwGeTQtAU7trnCqlZpF5Y28W6qFph
wK8RDazxPZycbF7Gv1G58Fh7Az/SEOaDjAZE6LhveE6h0xkMAw3d8mCstcplSw4h
10k9sLwvJysRN8DYEFMQrQY20PC2hFehLPjD2m/1kMCMf9z+krXQr0EryOdB5dcL
Eu+KjL6PlGMSH6oSjkFK/ZQKLwYfTEPL3yvtIcu/Pyjq6L8PtFJof4IzyujSdZ17
++NBLoOxhbYMoa9d5bZyZ8owG155hONyF6sLeaXt0gzX+nMx9R8kLkPuLQPNy0ZD
lOObWDpWehTo5Y7YSe/e78x4AO0Y08Ye178NzOyzMhes+SFq70nsPsvBhUZQdT8F
uFoHdzcJfvWlQcJA3pKk9J9hRf0PvsDJjP9iE9wsREFhs9mgRIIZkfNyLMIumXjU
T7zYtAnXFzIRLq4nsHuwtmgzwV8KVmFDY8wCqGVuOVySZFJpVqcFDNwZu+aeu3ix
CwFVS7oCBpx6SxRdFIwB3+mVSVIH+SP6VfGAWpQtPDOajUu4sJaT/CA3z7Uhv2so
GEfnmz5yDSzxfz4pMna78S2MrwN/PEcUjajTvZkHaFGwH1XlFibFJouTM6HDPjTd
V2WX6b440rg/XX8WODMys7PENvAY0u0TlaOEIvBOBdj57d8z327UgbdMwmcHbkBV
xYJdMrT9v/gvG8dCb9mxD3xB4BJU1jPO+tDg1kpUhUOskcGSZ9wRUPbEhydkdZfF
ttL5B2k0HSFUHk/z1U5Mk5TPNr5CDRpIJtK9BRLvTiP2urjajdE0ewFQcfG5dxcu
5x436SQTF7so4lfwrJHwJrL7S44hKE+YzSDRXMQA/Pg57nhlSYqLBSyD9qwi/0hs
NVRCVH7EA6L6QIx7sDp3DLtAhEavjtNgi3UVUrsS9WgY8ZrPUs23wo2aeGTHDw2M
o9df8CrqDGANqQ3xR/peY1dhS/QH/0RlmR1sOQ7tTKnKW+/YDBkoAsIE+wIuYums
6/15Qvo6uHwN5t9EaeguMcImJVELXVOMqgfLCYsz+VvyQ2F9TwniLBYCLsx8PFlR
sBq8NqThnRr1Z4em2TvrP/1hRclT9B05TLlzhRldJxstJUrfNK08VDZD+2HEmXxi
ezTR6s2qjN5/ycqxQBgBX0Gh3CgyzzcRtdYnBjDqF5ISpu+exLmIWcpXMpvJHZZf
ya71lWML4ScX8HrRSAyRT1c/3n2GPwFxqwWEG5PmosMZ6ujC58kk6h3PfwSq89Tn
JXwh7DyDisnZL86ugiL+ncxiefipSso2XCmkqGJEALAc9ZYQ1Ksmu0ph+C/AEF63
oQZDNZW4nxLreCLjXNcQzB07OtRWILwM9z8gz4xPZADgmNo+HJjo2C70gq2jiKn2
RMCOS5hAPNu+WkytjC+qooY/IzWEMNWAgvM/RQQmDoWL7fufRr6MUH2rz+lvWYju
OsBHo/mU4bSxWFM2GWHwY7o6UpeQ1NPwLUOgoU5BKSG8T/Rq/TYxMzCJZ8qbhf3D
Ifuf3HkjgQ5WqR/BZLbInRBbDybQpNKQDUuKUsbE0nvfAqATZQxTOTtMq1zmgMro
fEFpHJSAZ1AHlLGPxtoxtjwsJJxoi8fW6quUc+frKBWcaiJG1kF70JrfScZA91Ag
HBK9BpELMYlEmCWoCNGcWQrbiwccpufJCYT/VSbiHLsV//TVnXbBp2W93H+g01R1
chVD21JQZmZrAukQmZ3rFNEHD2/4WwAndmMkeiOrTlj+qW9MQyVsszjYrV4mC5gd
ZOzckBWgesYnCqtUeRsBHNzwssjYJqGmv5nheXN3CghxUP6CUc2Q/Yo2OsfWwHCO
QDALl53Kg49JWvA4ggLcXf91RpFsQCWh0DL5yoa/v/VGuytHerjBjHeXaNnVKjSR
0c5yTyV07Jpa54Qdx9AcTNvDSMpd5khSqhNn/oxe88y3Edyd6OA8Wz52WEXI8Zue
B0rCr6mT+Mons9yeBW0mcZrdJVoMXWCej2qtRLhr8gecxtdHDAwBzwY5NRWQQ39k
eNwLsNEWNRt2WQmWNC94F+qk79ItkJ/W6+BAuRLd/SMgAanPjJiqfL+vBP/cO7/K
QG1DLLa4ADlPpLq53bYwEQKJfaC0EylE2IiEblJ0zbwCjL64OpAt6WFRXZLQ3AeC
bNosvaZ/TkTlpl6yhIQZ3kwIGy5fX3l0tujc7fE/wIpTTjUvnBVr/xhCRE6cdaea
Lqew9mcH0O3PB7CQsQrWfXJ7zAp9EWqRdGGVN7aB/0o6fNXU17e5J+V8gnopQapH
YvRRnjmKFxfBD+kCBygfhkR7lyeiN+yaa5/JZZpccYIwSE8+R9fKgXVPz3LTlxTm
NfnGgWZv17nF6jVLxBxOAB4ngwaGwkEvEM0Qsfxyj8/ZtXbKB2NguhEQTIr24Nsn
xppK+pGadLJ/ksyDnOcSEBUFTIOXKf/ORDPTGXP8C9L+4yNhHEnBDwFqqGGpJpH+
qepiKpICvGl67G89DJH9XP06MuTSCawASsulq6eGk0TynrbcCzqHZ8F96CCUcx5y
YZnoA/W/g8UCibk08XviT9MhfFtMwjfgssFPmeI1gsghnBqct2EQICd7v6o7qRq5
9sWGJb088EAaygmwgui93EgMgXYKgH4CI+Zf6RkIcMIXMPIoPQS432VrSXyuPu4G
9jFoA3hHcqbAMvaCcNoWOfmWVDnxkZD87RsMeBzy/fdxjckitUdGF73NJ66A7xLu
wREcdnhJM3ShpFRIWchkR77e8ZBYTjUNhOKjsANjPfZykyM9GyqR1CDmgmfRQbPV
bUZXdir3H2nk2SHossLcPcMos+WBEAEyytrAt2Xjc/TML2iIO9flUPqHbq3vrVjK
yzuzTUfF0JcPwljxnwgE7bCdO1MTHq9G9FzcnfOgKNl0D6+XSaWJ7hQx1lpu8QbU
YRab2VMzws/cAiF0hpKOxJpOQ8/sSNTAD+DZAYDadrgFaQOFotrYKtQ2A+wRm6xr
YqCHAcWG40nZsJD60RLbabo0og3czsyxHlpZH4TUFyt84Xvu0LK8Eylw9cBMwOKv
I8MILxIzcI3k7c0da1hIc89w4Rd7Ehk/up7tYJ+YePIwmLcqgt8eaZWb3jCrSk3g
SY3iZb5GfRhy9Fi2xJPROph+9qyngJjfyxRqtcWuTb8MME3Y89ALlYLrI/4ToyTc
hlB3xnfQmNZ0ImymS2hdlLTuToa7PBAi0n5cdskovos8yf/+DXfCJbtJ/1qod1X8
DhJJzlb4TKY0QQbAAUQKPWLvc7xArDyoRAYVPa5/Fwl036tW1h6dfFh8vlUYl4Y1
GFXkpbGiEr1NRLiyUXTOIaaFh57pgoEZv1iUrlBNj38Sbf6cVM6ihNqRkCBO3BMQ
vClvfqcaNzMFdCrt+bLGU4KLlKZ8pvrjprVSkVBga/DHhv1OJEd4Rt/MfJLnZnqF
PnxlNGLjwXSo5QcsLIgYUYQ7jUZxvLBS9cC/tTQ8zZsD8kQA0hG+XL5qfNfF9yy+
pHI10Fcd6x70Vah0CeSOo5un2OK1XGy84f0qpTslgx30NQ9YmsHgz3zBC0tI85yo
ZE2zJ3FiWJTpAwipSr656a0iJ7sNixBoU2btY929DPiVzRHr0b84qCtoJwdSJOBD
gP514OBtLmhIO9/STL/hZR1YFMuJ0742kuSUxHYRXRPm1c8pC6Qvk4kOFT06dIxS
zFL6QlwRQql4cJDWPAkZrA3OiufEtD0G2pz6KKaCiQS4oH3RcvE4k1T46IQKakGI
rSBQ0KAD9DcteBZazOtaWaEtJMmXYAqCcMLHYvz525FRhtgjlxm6PoqoitiyBphY
m0CbUUcdLDGTp5lAkCYFMuD6R6phgtDmQeHNPXWhrg8TkS+qS6M24it9V9qHzTX6
/Mz1RLVnDkKA71FO3mCTHTh2Un5w5DXzKhOjxTqChIFEpdib5U8CefxCqeRlwf9l
giArdfIr86a59ja2hXpUqiVaVY67Xg/DqcsnMwLOHVN57TNuDcQY7LH978nJ/bMr
CW8mlcKTcdP8hPGRtPzj2IBqZDjLdR6mQKsle7iL+ym6kslkdMpSFOgMeKxt19j2
kUr9BCkTppctqeMp2sTaejpeD1JHN05OgF16aZc+LL2l01QQsFHwTQ9uhdGyPc3n
XKqlDzQAAJKT+/Pod5w3+jfpt8N5Tv8cgJberaHT4fZuxxI2bhb+3ItGCKwnqFXr
NhLmbv48gZpFGv+ta0CptsgM72fHWst332vhO5XHj9nBwKheleJ+jV0z2lTknflT
gvZ7HAUNHmW7kAgPFhcYem54oA+bZ/eCbY5ZtbFVfkjGPL2uUuAzrqRxzD0PgDMC
WNnu0FpZI7KrYykWELvq/3qOiSTXiu7d+7EdK7uBOF/kuIrL6zfEr4p9DGWn7elU
gl42elxj+hsovlMv0uiNW511nR0xX4cKotyFbvXYemW9edcgvWUCa3yWUY7pdh2s
W9zw0GHWjNJNqf4J/GESFgRcz+wT4X7OmTGR5rfxFAoj+LEZ1fkcAJBeHmaVzZlZ
bI79h8Li9R8GjhU2b8g5ryb7mY0b2oxq/U7Y0AtGyoWTST8wCD4PRMDJgD1nbKr2
LWb5kmTedrH8cwtYB73F7wjUkxTtzkQnPaFqv4Tx31CJ3QhV5WXdZZj4cCzcWbtu
EXgetgRLqsU3OnZ9bMqXOol6c9yd1iWwhZLHs+jNpmj0cNkA1bnRrmHWPjcFZc71
n6+d+ll8QzPR6y5fDmqw5eKiZkOmjHYK9k6WsLRBo/2wwDlapRuDTeW+AwW+GWWj
PlG6NX6q94nYtVBmHw9dD2oXpN5EHxAva4Vj4o8LchqzkoAMYopln3JSGp1tsp0w
81miR9Qj/p6BGM3k9Q9+YdFMxrg61RGIaGH4/m5f8kTUkIxCL6EicLZZaUZjHony
uMR0tIy1Zp8sBBn+5IJes8s1MvvTFBRomsSiGT0yyCnNgfBWjppm8jopAMKJo//k
kbOM1M7xQtmnwFXML9eyb9/Xy4sZyAPW9BSmvdSOK1hmkDushJ1jSvvYGQfjFAPT
tBUkkKCfU1d+j8x0Dsjj9SUn+YUv/S0z+NufzhEHg7fUufBqMjUg8tJJlthfPI63
HCetlMAP8/umpnwfh0jlt6bSL9H68C8XikvR7CPMu1v0UjzUvAKLePXuivdMud5p
i7Yox3WFk3Cw/clLW1iAJPhNaGrgTlKPajVX7wR1b2YSv9w+f4fOfMxVwHkN0QoT
c9IGeKO5SxzI4m8VlNPGcjjxIbXwXkXPdZaFGw5T5iW5q+y2JMzFhWlRcwH0pEG8
NcRdtGyDW3DtG4rWO3ZED1kmNpbt/JS2eTZezlMhQuhSYob6y5owAxEzQtuUCJ5n
iGX+kthw/uBiaxSbaCsZLaK4Kylqpl49wVF8R3/mTLv73rMhqt5clWXPsdkcSf0F
WvAJr5oGxHkAjBlIt6Y1cRbQ/JtbMPdAxPKCFdB8jDj8Aler56CwBjSOjIdYdsLq
XHZEKKHtOLI3v2jIQORacbDQoKTWR5T+tQNLCKQNTNsvvY269zsfbmgatozUgAJb
af82I5OypHNXcMWiw5IlTbOWtVo/sN8yOxkmzFE1XzagHqsJjTtWKfLSu2E+PzSF
IEq0NQjAcyll4R1RSmXSNi8fJ6kW8Ptl1pBHxD/xOktZSQ0OcZj4NFjajcPpS61R
cBk0IpWOLevWf6Nk210TD0suK+TeAiGoW3m0QZvWtlly97BqqmswrhdxUvuLv3vM
MdiPMPtDEh5D05uZ0Ajy91YXQL4rZcipLXm4egpEKkKmkgV7ptMr4rFFliAgmy5z
akzaCcY080Eol2sFhFQFPyPXHGhM9Yj6UT6NurrYF/q1nD01h2rNg2EPH1umZ2st
d0NFg9Zfql7VIemr62n+KN9rSnBiWZTK7yXlmFi+YF1f3MkH6iGkTPo2r6pqBhqn
XJ+VQjm9//FRkRAoSgFSpWDnH2LS49Jg+3TAjLLANFfyaB15eALIopkc1HWk3N4z
Ix1K2U3tMKpgAn1YrgL4m/cN3zqXcVAS7gzZUblJO6NDj126SjeNGfEXqHj9ikNm
U8VMh/VEOYEwAQrx+/+cHdQH/H4jwsdmCuL+4z9qZTdLB4BVf0cRS+6L/X3Yn59f
A3KPb9QnllN5v+sd1IvDQik0Ko+pjMb9jK/sMMfOFJby/ZTCVhBp581WwPPOmRA1
z3Y11rJpBmV9xoNHZOjmdRnumsOuMtRHMwil9WKR8e7s56NyPlidlOxC2fjM81MG
Csm3hc0Hxp8YvF0UOVH+wE5RJznUiG1Sj7oQG6MWwqx7gpG1aDjg7dhsehsghQwD
iZHrW193sCB2giI1/IjEfnaJguSzNKlkj9uws2I9FlTmcUpepW0s7rM/QVZc6GnG
+i95yvFjZqfGry9eBp0NDaIURGXulcolmk5VYcaG1S6drbfXBLcvG5ZCU2Cc5V5k
tEKdOlCMyfeg4lBhaDJhl53TwGNVvtUBbaBa1NEz5XNesUSZ9gSkgkiXQ6gnLhyL
BKhY79G3aeMwRWM+cxODe9hxNRZ/mgKoZMijSjYJ2WZfDLRtJr9QG+HxwoP+Yl9J
rJ6En8Hc/COnwZyQLi+vHO5QNiX6jx2SZH4Rxz7ExtXE+SNrSfmfpjqu84qWhtH/
Ce/JAijzAO0f0PxOH05nSW66nGdiMzR71UuBTz+/W5JaIZJR0vdrQ6itbGCbrZAU
vtMQ99AbH/5x3pInxokkcPac13ryapz0EVcteaow9wAlzB4rcYmPClYQT7vpHD95
I2EDH2nfzUK4/imub+dMbHaGprqfuiGhWAJv6j7wKfH9XBJRg65PMeU3CeblsL1y
2pbkTNn3BMRP8Lj23E5ZoDqSZDhnmE9jLPcizyfMYBbolN67GlRNnfuyQlAmYzLD
x5VoP+xRtR5Z//3jOPAYTTR3OxPwJ9vIGi8jXDoSkRJDhJgyOtccuiVbyeKUN8xh
h11SWANmOe0VGz9ip7DZO/lYFA+Agd+YVVEPSUmDaw3qxuY7/LtCJMFQukeYdQSq
TBxSxQsXBhZRQwU2SOkTlFiIypNS+xdCynOZ3oN2a7hyHmde5rwAZj/eovUWinFJ
M2Gp/TcX8cL73Fgmx8LTchZvJgr/Y8jwTqkUQcurgW73d58eL5L0drm5lBT5JM9U
Q9yq5AMkZ329d78I6B/6x3SmAg3XZD70LUV5+MMHScZ6+HCFi9jrrkOOyyuyKlK0
p6WVDYNacjsO6hD5d7XidpvuFzX62kpBf7REkWDX9jZf7s37AgfKKCFoT9n1Ogh1
ay8ZEakUrlWe7EjNovEOR12oQ5U2eeO5js9JiclILAPzEMRWVWV+l5PzeIE0CDV4
w/nrLwENq0ltgM2/349HasAxrccgakKE+hxHHDyvgRgsbeJqkmeQ78GWLbPycaE1
XrDR0xRHRWI3cygU3AhJX/LEKlS+gPs3XiOJtbQX5VK3pZ0yuCtFN92veqeD7yAI
Ds7+AVOyC0H5OqshzGt7Y9KrG6MSMC0GfxQMdFQQDbmJEKJod1JKfkh4iwb9sTFU
RJCANQHv5nftaUfr1SC8TeUBPEiG08rVpcmNuGLwhW9E2z+Q7++hNzZg5/CV4Hrj
WkIYvKANat5tukeVFY/jaStbYZ4/zOSsgm+nABIKzHEPcTLdGz7BjkNnNaYfmKOT
Kd5Vd+TiNo8S9nCpDQvkvEs4BupJNFIY2PLuBD6p0iAurFJmimNuKxwMOwcloQ67
5YkFeD+qWfQsbJkCUtuO2AqLUxEM9TD0MVX9kCw4NocPN7+IH4cXHf+ZKI1euTGQ
2HwoXtz/FaR+ButBW3UVT0sAAVSaAizNKQhir5OD/EzOOH51qy7LY+bTrYzqAHzd
5CKuX5fFcABJmNWvi0arWRjzEqzPxi5Tsksd5FNy1YsijHM8Efy21tGZOlatAjwI
HOgFXU7nSgK7R6bgxBq+jtY+WEST6ju/Zzk1NKGuK0AMWHNZrQL4FcibbIPFhhJ7
2pJz6J4YEo3Pst6Jb1RvbNHcM2WFKzvT17chVbTKQdGQd869h7KCJEy+QRkWyax7
SGUC6VJnelvGLW5rmihZxPPzwH0j8/hkjhk6GXes6MyHBOl2yLUWAndHuEnbQ25K
Nd8p48Di32Mk7T+ww7ZjbtMpkBPxt8Stg0/ybXTQMpl3aF21NwJd0lX+vU4jVU3A
Bl+r7WGfsTkxIZRpg0A8Lab0JMAQp/L/9vCBgHJPFOE+Mvb9XcPIUitjkcVevTQn
4kXWSlGokin6ya7jcWljB02jpzePH1BbZIfRk7iRXq6xrImfTN75E+88o+cf9rF4
w2Qlam22GPx6/aPOKLNP0rKHClFE0wDq3+wIVTtf+qsD1c8WuLjBJb5o1AC+x3pY
gUpJJP7FAgEbYSMKl+lwOeOE+i0sVfO3oruHe3uRH+Ew0JsPgj5SAu9mNS3bnqeW
GVGXoyt76IfgXLD0u7mxO0DEl0cwaVzNOWIO2kZ5bq8gjtKYroiurwhC/MrJwRpf
kAlHCSoY0VqkwINEMLJus12+dmSARD4OLbL5Xmu0Uz7QurZMPD9B8dS/jm1bDzqo
2BcXZBDlbjCWYYn/bwQPrx4sAq5D0yqnirqSO2mz9pezOEnCijbCGCdKICxmi+Y+
c9DSGLeKjwyxxeiNDzz0BMIjsROD53Y4J6aym65n/FR2tN0rcbWtPTHtVs4BwXCE
ZDBDo0UHWzS6lfI304iGA3drJckDcexBCxUqmlQmD7s0tdXMN8SbAkMjyIHe3og9
oJSIEyH304XUgB75XaFRzQk5ySZQp4vhrwM7KMjIL2ewNPHg9TK3+ML1jieSg+rL
0E3Fjwi4HuXY/jex80zMJNuV6eW2PGXz0x0CSaNcd9d/RVsxlez5SQZvGLqRm7JR
G+XZzmAmn6y6YkHg4HbX1ooA2hMJ8hUVIeG/F8E8oq8UYkDmQ1//e+hIj59GRPDa
pKZmYyD5Eatvh6mUvTDZd1F8t/bkYf+ENFMENk+bgwEnWLs8dVjTwu/+Sx98oL8G
xTMADChFsuv2VqCJXB0KPLMBm8x7M8ZjEyUopcS4ykpuF+xSgJkM66w7bxHSuIld
n7YDiiafg79J+FA8sUmk2YPjXvxqvmUrLttIILQlcMcwpayp0ZvKWgfsEHqS/4Rc
WOsHtuHZlvjh+iH2JYPB7mSgbOnKhCXivxTU6j6zrD8YRi8KGT7fb7zG7olc1JHP
pImPQbYbAolDk5Un+liWzh7uNffhnpU+pTHr2K/8OWiyuGJuZbIadUrhae0qRCBT
V1TnrSXGZIwgIlwHYkk5cpSjKavrbcaR/eCfuyaJY1duH+AugljA+YRBXehjLVOI
+ieBhIjXRY+nz2hs5yEQ14wsXBbW7KTJjqkikinHQX0uPIrej+BkHkt8CmFBSMEZ
Bb4ajeekzOT6NRxKcJeU5LmTix5ODIBLvqy0aMKlDCCtBNdGAmF7IfoO//kZAVqk
65JYEV2xq8YEljQDu9ptgrsrZnLxrV2TAWOdTJA9YTysum5MvMydjDklR9aoPTyx
d/ZGBRVLioueQfpH0qPlqwiS4rrnUDjixtpFbdagPw2040x4SWsurll/E+Wcr69T
XFsQYC/PSBuo/Q2tT6+OpfziuYvfai6otP1RrXNy8tK6UA8WcwHMeMV3VsUxpU03
tatRVQ30MaUrH5bw0i/uoVxamPD6c2+58E+z7OUy8ccWTiAyM2wvVS8v/eJMBRVf
CI5GxfnXsZtCVd0NImXIfuNU1UhN9iM8DcJX0PvSMS1+BDIQ/xtgDfQ6lbDSj4mJ
WTuRmsxlmxCgiWnjaG1zQwZrgWR7yTov+gKby5j8YMd/d7GYP0r5UPHgjkBpZnUG
oRHUwgO+Lh6+zvVOWJiCugcuDjhy4IQjrIV68WYzzMa2nPZQ3Otlkb2mDhWIKamE
nzyId6OY2ZQicSr9L0EZ3flTUDuxr9Uz19txlyq/uXbUiy9BQ90VQO+nlb8Ah9Q5
s3lGkc5R753opVgDisqiPLjx7BM4/pmR8Cm9T+0cjHazUmka4HkTJuQTCo18yzN5
v+dInL5brkIR2C53XRiVReyYplwsp3oEkMJkqDQyzy8ckoTyaugDBqbmARrR2SsT
74NGs4hvsfBhl/zXlQXX3u8cWde50AfWTBYnjb4aQ2llGLYPOgQ8Ci0qpQrKN+Ni
PKuWHxWhsuac6S+nlPvjfjcLwOhX2tcn/v3iIx+gqQ2Nt/nFDucHLDlIXaY0d+J9
vFEiF/kTL3HSWmWY2OgiG86H07uaOvT8ZT4k0NCgT6NFSC5Z7a8tLZW+4eyUhINu
fwPKJyv2WF4x5mgnismC13s19eG9t81oy7LCyD4e9GEPr9RNyTvvyZtRxVsmCt5d
lGWmWyq8+vzvBfs9wXn4m5I/6h0+Jh6EmR2Pt1kO2yTruBe71Zb+0Ra7x4nX76vU
hOs89MiSB3bIOxK9ceaL8ZO1Xe5KkgxElv6vTUk9gYOOoylLa4Dbltl4VFQNomLE
aLP8LEH5JFToH6ZotGWE5dLjo6pnJk03NeaTFc2AiR4XdhW8xXoAgs6n9aEz8d27
DAJ91TjlhYcRiOI3U3mfKVSv5ErBcWTpB9wFNNj4K2gmZ7fsQi2hzehG6gdJuYZ4
Ogkdl/6LYB/5huRdapSrSutXS4uh3y+iZr1WV1rWgV6AfVDwH02s+o0AEwuyq+cs
0yHO1Pdu3YX/M2h+vkMA1GefNX6wajTInOZEPbBTDutCjUPaWhzAaOB2cByg2LgN
puGSLDWp7+AhkKNpG13tRwW9wIpTqWFz2/b1fwExlFFUa3UNPEmdaNxbh+r0nU2q
2fDtwbLEs+pT44PLI98g/3hWQB2conjMs9P4w1HF9zajEgK+YcrYOznzEHKiONiQ
BY+criSwZCUWuvhgU6+jdPvrrDK3nYs9gSbm7vLVpqmfABIr2WkSLK0nl3GGG0z1
8AuIFuO1YqYzMwO64W4xRCukYcBQBRl22H42CTcges+LNBdSw1SXGZJBBAgQSJIU
lSBQG/i4YN/m65WmdnPcqRgcYZR/CQWMYlJHWNZh2KSrDRF+nlHBVf0fMwHpp0oZ
HMkOYzIKVCoAgiTsj2nzXMp07gwOPj93aIt607OUmJz5CB04zVpdAqirtA5aNdIi
HTL18ssIeVJZNpk6DH/PqxK/VVYg7f8vQlShiNW8vd7zhIUNr9hPeubdwHLfF+xj
zUyUKoBtByiv/giZhGGHJwfbj/dxB+XmUEmBi+ugrSerLwpqrpDr5s4dDvhfM85s
cjNu9OQL6QFFnc0iO0NysGjptqpD4tqaK79l6Uiz2ytNvYkgbo+nzvKf2UjKGeS9
Z1MYUJm5Tg8GP8UvBx/zaktjWtb/Fm0tgmAcc+JfhKbuu0zrh1TNs6I1XO8F1TJa
YKaDex5JbI00xCd6NiQZlrlB70BJ4xcgJPXmo3fITVfRo9dO9o+tdg5F4Gx3hH7B
zhY0Sy6TU6eiej6c5uOsMzEcLh4Ft/85U7QHppzuwbK8swj3ZJ+jY8vO7WjTgCaI
KHUguPz6SWScPFXbGedI6VRYvMJpcU/ctDUr6o7aKJfHPRstNNRLx0+4f9yvQ7ZG
DIi9RsA/Z1kBMS9zDQ84SXe7a5Rt59KBO3w3mMe0hT26apo6IQ1TB3QI4eunw0s8
GlGUu0UGTN3DS1tcOarAtuvItDATupCu10UcU1gGzzLCC2GrF4/3BZPiHyUw/xGK
0pC4CZfM+3pl6WDeTx2ZTmtEfF5geJ8CRq7+k6toG6sITQTWf1+M158J2FvhQEe+
3uZ0IXBcuRQ3N3jXrvnoDR5VQbFRvTzZS5H6wIse5Wlu5JxsGkLdyb/V4oWQgzL0
u1q3bVAAkSyVrh+LakYs2VZdYN+UqnRyE7L+kVxai/Uzze7UKPXWXsd8EjmBFQX3
RV/mjBXmGEz/AnUIndNJicHBGS8Ic2lszOGAPmOQs3qTTCTeV6FCKdCnfUBlkFuk
fDVuGG8TbNvESrwNAv4+VPuCapaDHRfxmRxzKkz9lYnBtUgJyMtc7Kj+sAIVWb7/
LK+o2RoWT0ORmUTZ2yIu08EJFC8kvY57ODs6sC0GLIAWG13VecN6VatH4+EmLmYt
e2leZcjUwoxk9J9SBJ9iFLEozhC6dcrw5UZQj0NtYDUsmmfW4efZSUl16PKcPEd/
GVJ401QQ/PLfbRG2hFj/aRGwYwXdjZs+FdunH9zVi3Suau8ctuUKpiQmAJSUondQ
rAG1lpSTdG12LpgJyMSYiQbDPBASbEtcyvmaEZMA78jNjt9WBu1ffKo114oEJ4Hq
CcR+l02Yhg3LTE4FMSDjz26x3uQ4PP10O95RBgTvqS/kCxXyIoO2I+2IWt3Qh+kM
loywtC3gGI6pU4kqPNO4Su7rtMjemZVeLFeOKq5Ce6ctwHnSFhbn4NkHp0P5sada
LM6Jf0fxhr4UCLtu36GZwmiRY8vjIjyRxLe7id4y2jrAvv9W1GD4NYszPJe67yRV
P78IVHQ2ttt8SRMFwJ/AaujCHPs8vgTPiwZkTYaI3EGanQMFexrB6w9vmMw8caje
R/Mo4Wlb9ZnVoQfbzka0yFFuo3sna7YxGzHHhGo5cv9mTXMRsoJm064YNKfEeHPo
UANGqKlpkQ7b/kr04UlKSdRFgknBLf0foTv2otOf8H4Ar8Twa/Y8ljUhpJeT+n6w
7Tvx6iq5XZCcT6g9DdUBNeBnM7gywYUsRx20+N43Ua70I79cStoyIC2No5smgP/5
6p25aaYuPsVwAqd/YLIoXZ7WOhhoDixlm1ze6NgeRU0WOhQiDSHnYj8Uu1a/w9eo
nQHa8ldBdILH4D0rWMj9zsUf6Y9WwD0f1wJPOmFQnbRAS0Q1ZRpAg0GksmnoEK5V
PuZEcwTlXvaKBL23bHAkxrPVTqMEB6a48TRmyba4HcmmuOmGB36CAwIvZXMfRQax
R4JsIr7ZSw7VLuNXgGBIqCi8O54uQNOP5TwT6DnVRzXdBU0NrNhrGME0b2aETtQE
0xQ9RECcMbd0W0i5vvaBxDKSnrbZ8S4g0ua1wGZnURnkr4ZV3W+KPCLfIhOm4n8d
4mZ3HV5C1yq/osYGUnizNWkPp6KwnxGzj9uTyRZWZ/U/mxZ/jTp/2v3RKGqSLRyn
DF1uj45q4U8XaqT3HjPkHxjB1R4WN7ZV5J9JLZYa8IDSwdmUPDugQMPUllkjNNm3
pDtsWu6KXRRzJXcjPVsN8Bs3+ssh63criL2xP3i+QA8cMES8XLhjdKgRz38YRP5q
1sIdBMBJQFsuxnmJFRwPs7QAlU4bggsZQY2z4RA+KADczIj9Sy7KatvLTbPyqD8a
ejw2MgiI3/Abazl1bcwnwu7WqK+LtR27mSoQA2YTQzJJ9CA0JUHWl+vdi2zq51i6
iwd404oXjpo0GnNYJ7wCB4jRaS6lu+S48gSzTqqNeXleXcJvPdBaS8I+1THXpX3d
tFXF2hU+kydStqYJjPZ3Edmhwja812QgaKZVlzxwwwZC7WV1K4CONW6eNkRE/Ac/
ssFV8MM3oyE7s4mjCgT6mIKVAEaQ/8I9tKxSUok2Z9gq71X29MS3CG51ZqU6ImYS
Q11KlvNVWGxaO7u55qJcsc0NTPU5SGCsdyn1btAUWpCiauJK4LydSc/uXBY0M5FF
rtxmpss1d1TAPl92hLURONMEHqsS0h3BoIxPrJFt9W+S2PpFR+yvvsVob8ZVtgq+
2FESPo+wR4kgfLIev15iTnpmC1NOKSpekItItt+uCMuhmZ+vuBYh3slgRDSjZvIo
AbCjvP/4y2t45Vjle+8RJA4fAsNHR837coIwu1gZEytfSQN3fk/VeWNKWRqx1dUb
2xcVEXVZuK6AePr5+nbkkQauSb2Q6No1THUyY2tIARdtr7wN3ywPWpcRZBxVv7PY
dK1ZXTPby2ExOQunkrxtZTZIvXcrS+69SnBC3BePINxhTEdUsy0MbhYe1ayssGFq
fNf8q7UcCBxepwfjWp7kQeIcr+1RF0yo746kFai/58uJPuVRqAULhYs+rSLcgkk0
1rDmkrmZor38cADQRiGhdxuYd+EKSJ9laMW21KGhbf7MSSXNLMkYHAAUKXWX8PdV
2RJ57zy2KxDo7YC+l5HPSh4ASHDV90by1XTAqPK+Vgb5inWVgebH5lY/zkORKVaC
zv7aht649HZ538r8fZfQ9+HfvaKe+vjOLu2vkQz1cQX21W3nWBBJq78QGgwDfTNH
TQ7rRet0grBuQ2jtmNrtNe1CCLtoMIRdXYLp6/viBytTPyY8rRThFd4utGUpnLqi
ZBPK1Rja6wcMRAsAcnThMsGdi+FAnpUqGiBqpF5iK/4Z3oO7SObjFWJYKvpXCkoV
wzp2k2Okhn2/dd1CfnmNGIoPC6/KSfA+jn0SARJyg/5vejKBMfOuWhPGeUxZ8Z96
pXwmkTBDzux1lc2e6pVQ0klrEmT0OhADbM12QggVJWVGXeEcS3cuczvyFruh9RJT
KaYFWzY5ezPAHrKZ5T65lIyTwaIAxb7WzXevUKzpNsXGWcM5T+lXNcoj1d+pH6hZ
ZN6+bfEJTIm37QjLoyiMYxwgj9uUfARnqIvWOLEcRHdiaF6rXRuiMquDGCuSBxCT
OiOOLu1XGjjX3teu8IdLHZ+17MKYBwehuW8dFQbdZFUhAYOglgcbqnJYmXmD4tG7
YF8Div0YNGTKaJ8WY1aayWq7UikYBlLPjwDELCswG3olE7lRO0TclGP4BjmgINe/
0h1a3K8V9HJLaI70C3vBHea4C83X12h4pAH+wgI0DOSpO1PQX039eunvNAsX0Qm9
vvhcdRApwzND8I0PaVYyxuIe409WUmJLT+fn9r/34OVjbXSgYprKw65kb26L9/1T
AAB9bAZmBBfMYws1qHYFRjZYB9f9ymIjtYZYt1TzwxDTM+eD3rxnQdk6zdWM7Sqn
cXGBZm7voPzUGa4obJzitPSl0U2q9n1LBtnddIHKupMJXxChkjBqoWMLFI3NKo9m
5Ot+Izdd5u52AuG6kTePPmB5MvUyhdHr2Ls7ZDv4mGgjLpM3zqVqa80Lsb1V7Jig
3LdnhwH+97FHNJMq/HZfkoAkGiLQ9Um1jV33+10qaOfioJTvGefZVQz0tlz29wo+
JyqmT6oVj8uhRxA0E/S5j9IFxLOx2pSgr9tj8N7oydiOvOF1QU+wjfwTsz6zTNB8
61TCer0jRtp1CDoeSiRNOMLQzDfWZj8C/17iikec33pZubMXiuMh2qWgUz539Z/O
30rjpujNMlRBFSFv7PhQOy9jNbkZzvPQCsrmTfKEelS2PLt7W8gkGT/SAOoJqpG5
6kjKO1kfXVkylG8H6dKzA5ZEGjmJ81qyEcdbbb/CB4QCT+3yS8skWRSrO7Gt9jTs
uup+VJM+jzNvhvSZRmKR2dP6A+ZLa2L1/Na3c1J0+OhAUXwjS4O4xDZmGrYtbBuK
tNQ5XlRqYXGLc0/ybclK6hZmXhxxU6xUuEyzJ71gHg+Rp+6SyhiqBFi+g+tpS1/5
FIGqJfgoe21rc0WaUJTn5Mc+H8L4pqfJEfUyG8/bv+vgdlZ2yz0yooBJr5b2XY5x
+CdH9amIcZxZmZiFWIKKvwuB1S78CPsH0f1GihZh25chAxq+qzCMpyu2FWPWcPbA
lTwNdM4ilIqyWmt2BUraGhuTovAom7cKhyAd5guaMci6ctf9Fge924RnA7aUetYK
IKPhyN2YV1pMoU3QlmZSwuh6z4lbGRLYRs+046wcHYG3F5F3P6D/UlEF1jsmVQ01
ciQ/dBM+IHve4cN0d0NlSFqpRuF/dNytgfy5ieXqAE+j2lTmUjRVGucVb0WaGXlT
zMFCp97kql3lFEicj79c2SEzI4hViyLmc5AeIemsr41hCbTge4zfGOw0YwtDi+Vk
4Cdl5F+uRtWe4GpfPn5yvW9z100/9FiXr3bSM39oUqLUknMCygPNz8f5IHjb2QpZ
igKT+XwBF4naexS+UtTPyOjj5EoX0pSfoCyaxIg3iDsbSeO3bZ9ReCnHHwFJyJLJ
LZSfZhBILe6GW7kFe1vxOqubyTKPko2HIRmbrVGi4QKoTyCmMGIrXBoUQPZWi6Wg
l4xXwOvpYMVe5PTy9xrERK2FKJt53AVCzb+XqRG7xcKd/N2yiM2r8icd7Xf6YYds
T8sFtcnlkaGRd+Qu4dkMgMNhq/8kWM1XnMeDQjQI+6jCMrXLVbysqrrHK/xxvWvc
M9eRw7Dh9nSZHlH4pYCbVMwWnKwOuR5AbBpAS4YemDEs3qBqRVgvJZNFWqNCaQ8v
5wTJ3dDGrBDBNwUAGEEHyrraKqfRl9t6l8CtGMt5DwjV+gGidLLuTWmHN50A7YRB
ius7hhowm24RBJ/rcB0jJQuuv316rjflIiK6V6cTUjmQIcMfpNvDZbrqRh2NS6Bk
2ALR3hh03hSphTcaDrXdnGulrqn5qMw1V/ShXarIZHJ44dMrE8Dy9/qyfTuF2qVG
5uhmmmC1gIsbkG44x/A4di/8JY81tNptbaisAZOVVclk17+yGx6i86EhPawcV1t4
tDnVPyaETeacwib4iMBz1IYIVaTQ5ExO10ztFKAvY8IlvBqFISa8OQpgt6dO1a3w
gJtoMt1BTQmXXjvkliD6lnZTBHzYOF/aistDRH7UFzBRFOtjNJkGDGJR0nUtKLxO
tA4IKjoDRs3kcjjkRyJBnTNec0EmASaqRSxo1xjCYlqOILcO/8KUQyGFMTaWOOBR
MReu11rS86OixgM37MgB6EgXPoESWevsW87F38mCI/LZ/RUWDAG5+7o7AA18UUyq
PdlRLpsyQGHoWt402fGx5iXr12d6nZM7+JLbAbDqEmdeApSbfJ/HGsabidRmBOcd
f+h35X3UhsOVtreYL+MNNtDIcGEeC6hHJClzUIEJpYo0kS+vMgGilh2jcisPnFLy
cR2nNoN54HeB5nzvFm90+rsffQAudwMQhiWDO8REeMgUB30Tx6BajcVE7xX104yL
lpf5OtEsC4epf7eYTppvuwLTL5xuSo7K5HTBUj4akgj3Y1ufyBnFxWg3KTqVvhSf
OLTq1/ALMbuSUN6ACgcopT2cAqkCTFOwXJLGJAZBHeU0Faz6IythDIP1fi36oB6h
Wk94e8zieGgW0CLy7HGPdjV1vxNmPVKd9VDSN0bAZ2JRT/3XtIhChbKEwvaS4YSt
oh56r3TI9PkWkfeGGejf1Dr5zO4udMMPH5+zamtiwzWgP0TrQjUVLP2F96NaoHJo
u8lMl5oXMuWgYWyYp+1skfTgKx58aD6JCB1L70p5urWmdoHfGGjjYfqBPOdT7bAt
UTUG/TlGTftXytLbTkB3FPSQCkbtYbYR6oyyQrNuVRPfM9cprVhI7JthEGrEZila
JQsMTpTw9eMkB6PhAo2w7BdyllSR3qGCXUUreoWfjac+AK1Dl5EExhn1kyHxWEWI
f1d1pqeZwUdeaOqTQtehSi0ijlcST6UYwTKkYdWE12zDDcPBhjq8vguTXKpwZ5OS
YHmXw8qZ+b+varqLNnGXXAah4DEOefkPkwxupYRzqqwgJ8VGohLy3KHT4tiuMY0f
4Q6iTVFo2MAjGEAu6wqZGM+kVW/7TJ6tqt5dgX6fCGRYqow3CYFagBGjx9/QwMC0
dHglXJ+LRulKg8kvbPeZa/gFd64MlNuKjwPOnkqKS1e6uE8JP4sR+ZJMVariGRnx
xErJEPYjwUn944cJF8OnqM2iS9lTZyAqxHFkKq5cLBtxL/zaWkMI9yYpoh1VsMyz
oUqFWbudfIoy0UoUWM1ZC4VWTRyztFuVzYvCgzO4atlPoeL1FHSsKgAgFg4UwZ2O
G8ySTC7DwRzKIh5eNb9swFc4RqCo2V9Uv9OCMg0pF9bO5UWHJacYNRGOkIu7IlzD
qkYXbqxxeRDXKDJs+/OiLxHx1ej+i7a/2k/O0tpyij+eBlpAzYHMYkHGhuJd/csY
pVYnpSmR94oR++FMgxDT9LWFYymtVWBVEudozmCSU6CyecLX8UfkaVLLcpz2pu+z
hnaEMWF1VDSiSqAszkcilDPO9EPEhUbY0U6jNf8+FYnptl+ZlPWPD4LATyFTWJE9
xgignfs/Dmo5IWQMFos0UAnoZNxeitg+9AtKPy+sHahT9kWBiuSEtVwggNPyJc4G
nxLBHj0Uay607NkH4WIEbzwpdeuoNWuRurtFve7MDjmuTiYDP/W2plCdzXhudKd6
HX9ABga5joMlB/cX8SI3XMimp45D9fS2zRMtUiV3ry7ZninQCD9skYBLA2mgQmqr
TBdYI4iI2rCwaX0tjm6/n7u18cpHshl9bLIUPYw4po9f6rl9zM+ljqqw8tHsrsIQ
93alLPF1a+3SULc+c3rcXqcA992OF8JftCnA2lQeXQ2QEUkq9Qg5k/RuVzsSFge1
yCBEzWIj4Ofl2eV9FKEUjrMTgKY5tEzyToTZBREngIm8K9rWgvZv/27z/LQZcnQd
GGmr1Zo0OHK4ZhNvBA6yVnW9mnk2Heu2OlIq+w0fE6DwVtzFWm6Cz5ON2EeRkF6p
z6LLHBfyT4vQv1il0uef6CoXhchuef/h3LIToe3ND6pj/X9OM/zWjC0P6xsR4Dus
q+/baSYf44ByTdnziqWqmgNtbGDvOmZGu96v+h61HP0/QdxmFUU45yqz8EizPw8M
S4iwqCxVev8bxfSiiN+J/ERQsJ2uOhYC6wGABOR8pFNhXkVoWD/0slhQThop5iUY
l3Xf3VbFGzEcKCvPckP4xpXLJLwXbRtShb9uV1RR17uFOhdCHdT2e/QhgePLIoew
7yHUkYUoD5D5if/ZOCqUV0Hqxyn+qQIK5dHzN3EzcpcrUC9BSXiRfJXstN0sT37K
0520J+9yoJ0RXDHc1VLh1Jc3VPHs8Q0pY15HLDnYm7/GRkO21DDSwIX9xpmlz0zb
hur++T7S/oVCsGEBWzpp8anDfSV6HOoeuFO+Gw+C7fHKXEE1cA/YBIOPF8jmP7u8
x1ldKROA3nPR5iBVVz/7gXuiaTJoDHqIQW78hzW0QBZZ59Y/kHgBzK+r64CJ1CJA
jRcgFRIiHAQ4f1Wlz6RaraxJd2pqqzQnXdUPkxtRqt9WjgbCsqSxs0nHRjp9kvUN
L5tOEVKPHyfg4BcBhnwncgQFgZlHpwVGTLr6iRF/H0+2Z7264sYmXyiIO4j85Yw/
MEe9R3hY1LRMZJmVrgrqaADgc0hUEuiMVrX5IJqsQ6ZTImabsLnj5kdl6ZMXsGtc
hQ+RDkWlFb2ENUPAK71U0kZJJnTU/bOokDQxmjg8zs5X2JYu9hM6R66dOgeor4Cx
VEDXm+i0gSnIgEuOrJFq8RSCzcHpF7vKySLEnq52aebHP2igfAJZzvtjckEta3tw
F7Gv9P4mQcV21U9YQpZVCmBhhD8DdTDE1Z21/JpXmLl2H2gXd1w37fS4Uj+KTUC4
BmZ4ogdWupF98+o4NpyR1BAgZrdnpp+psH1ki39ZE0EEKFhPubB8AF6L/I7mNcDF
8UeODYrMy9tLeQclvJ2q9I46lymu2v8YCpTWbBYRWOVvyFKaHy9QgNq36JrAtSYo
woBof28VFCGwxQ4qoy5mv3wDal6WFO+792OVZZk2XYoTkMzClD5LTx3HBu9pze05
aNYGmqn0A3ek7Gcv8AIu1nLlYLBdxM0gGKYOu5joUGmYMfxMPW7oJqaGaMB2H4Rf
i4DyjI3xWcinMAigmOT3dEBJLyJirqvEfQk0suR9V2qTW3lw7JEu3yz9w4pNgVT8
pu3B+vIwKe47UT+Eh4NyC37PEvr6Uuct7qcQQ0n5/jBi1JlmtZ3DjjtdY4kkrBa+
UxZZKvKoyXE1zF3odiQIIP+0VVx0ETuY3R0Kq+v3Ss+PJQxmygAz79cMI009rz07
PhIfO1AyrReD2l9Cz5qmfj6GK7P/bnADe4WcOW10NX6veeOu1i0HwiG5T7qHTfrp
Q24+A/GZ/nfoYoeJq465zYUU/ocZJm9B/xkHUUzZshI2GbE0PlGrADU36MQBCBuW
LYn/s1odWmh5W+U/u+Kxag8yfdyo4Tun/NDvXlY2qGHiiSLMda2H21AQ9uMPUteU
QZy7IgEh1UTVe4pjnu1Hymwq5cMbfIcajzGCTd7fhN8x3P2357b48pUsMzOoxaR6
62n+/ZPUUUFPcqSlrwGECleF67ps48mX8CY9g3+q7ThNBzDQoH5BUgxTldZB9r3T
l06v54SG0XwD0nM/GspnPwYk3be47TODYYsnj+A3K0WHattim4cuDa/o033N1Vt+
b4ri7vrm4uPzVdPmd0JjxonfgriVfznCwzeuullaq+fH5BAYDuSJ0JQVmuHrR3C0
7xKqVM3UCM6nrVQn6be1nSnqubYmecxhAnUzK1LFx9akpA1ZsDqAf5NTgiG/hYKz
HfS7C5cMRxFBJ8yj13Wnxjk55YGnJGinPlh6vfNKKBz2pE2xFdrNUKdU9lcQ5lyL
XraCaMRXGxwIR4uNjwGlnD8tD3ndYzkeqyuQXBkCdjVcAFov/LzWSH9n7cFgAJz8
SEG6/Tc/Y26t3QSTMMq20lE9lgHmJAN+xp7OectYm7UYzvq9OD5XFPR1rOrYJg2a
tj/4zC0xptRct8EQM0ChFJwrjB2R7gizujj1ZGZV3I4piR2zZRxR+9ZjwTyWiLCe
63tTm/ttGO3j19zN5nkkCMNsdKb3P/nRGSohhxYCu6+e2DPZV4ATgvDI3B5nqx2t
FIM4mBsZXOyHaN0O7BujUzlhS8YcNFIh3zm7+NasPkTNY9LPTp6I+/0LEyZFmkRM
Pommo1jfEjjOS8F7i7sXgsiOG4ihWN62nwHZlr++cmLs7zs651ygNg7C5QMgS6yL
nJFV+Viyfm0Mn0u4Q0mtcfSlcb7Ot04+bmI83tAcCqtTlEI0X7yfN2Tu7Ac6+ZbL
wEBrZ85mUBOMhTC3/ZnY0qzPvUjVaKtSupLo+n0+wf7ioyTETjXY0gKQ2jFtzgoy
OrcC6voR2Gb8KTOYo5S0NvF5xolGjBqvVl90NNDSU2hOgQUkCV+vB+1sUEcdOCC6
yjQtL5fCKkyFeVNPHqPNAZJz9lBL2j10UxunE/zfRl5tO41FdM2g+pOWGWIat9b3
ktdCpBw1s0+tlcz4y5AIiuWmEshpMIXZCe9pqfWdJ55MXR4hEUEZC4Y6aITNVWwH
uvI1NLdRpZHgxbQyMBoR14UvxB0qRibAEw1g422USOqXcGYaj++i5p/S4Cgu5/VL
bmysHc7oeiJue3ZW6coEVZ50XtWq6SD4nrTFIUH5QlKF864fkRJf2ndebscYKZNG
PdEC6UHYMwD/HflXhnCuw4iNm49BUWZCbus4Wdd+I5TzDT3sJBoCycrt/UZsZpP3
j9aoUl3XLw8GCJeNuOZd1vPzHmHZqH6V1ymfpNAccly3h72RcTMTCGS0gyFNYqM+
kEmvCDNmC+cAz0anPVU/Vyr+uBT8hFbM/p4O8JT9lijPKW34LiWVkw/VKIB68L5d
jEUDQnex3pn1au2uo7B5j53nPH6sPCwYgR8lrkJMG9Ww6hN4mqh63edwPADVmy3T
FmXG3RkkO9skoo2rsITCCpTeuRfQs65BKKD/ysLGYn/ZQEtnWLyZHRhZu8HID3JE
SLOFDryYBjhGKverOHNvxnlBINgMP9ehxDDHd4YQOdnPaCsQGZB7diVFH76C6m6c
KhU1e/od5gMEhnPy60E23DjnwDrtrIU/GemvmTleQw4/mxj7ND4/mkMQPTnjH0+B
z+KJljeUkLfwihQYLFDPM4SPceXWo+NRP3ichlV23PQrTzkA2+sb8uGYPo4oUFj1
cEEl0CDK9ce8jPeKG0fg0/al3De3hSxtLddMxv6iqc+DBQRt4XidT7B6cgSIWPgf
X4WU/xLbQ5qz6xLWqDNIs2JHBg7BTw2YFLg3jSLZBMibp05eUWeqvzBNBNRf2ine
F2L8Rt+Z7Cy3LxMo9+O5o8qQEsrEIF8tkdOPaFDS2enqwM9jUaTwGAb/berHHCXd
mycidax3edRsu3m54U2sTzgmkIlzlMoZMDpmA6v19CM5hO8yAdIu8t1BBlMCmVZB
J9O9NxjSjNQ+gKOiJVkPbk008RKOGLXsqPqaGQRZXE+GXrlQ4vOppDB8BB6zomU2
l2H1THy9rYp+YQZKrKx8B2mjoccyhEzKNcSA0ncuwoiQ7p2t44++InxMjPRr/Rfp
0tK8xTa8QqvIHbm2ezYcTvzEJ7b9nwCC++uxR+uQXVc+bBHB5AdO3CU1LxcBz/cX
Vi+gUhL3G8ld2iZ2Ms71Xa47PzacvG8T824hhCREz42h770imLcNu6gej1yJfHle
IRbLsq9OMn+4gwsL0gTVLzXhft8YcduqC+L1JhkE63Qa6Hldmo1WyuPERXhtngaF
TR6zOKC0bP5xsk1Sqs0WZWusJdxRFW1DraHpKcxwfDToC8K2KrEXsYwtX8sS7qF2
Kk2z+fupOlX+8WZKPO4CcwA/M293qDflSf69eseaKpensfU8fbdZXDtKwoTbSOLh
VGVLGjqau0VyH5UjEJ9goJf4TkdJg5hPXSLIkrUFPdZK7KSTW6u3LhfO5KR4brie
uJqWCE44zYeJdn/L9JVlZxPfVXapu0OHznrJIjg41v/giWtPCQmgkGzQOsG1G/vi
Q6+CtFGK0jcxA7PNdXEGxWsTihPLZZmce3kcaCOmxl+eo0NJL71d9mRxVbn7MFTz
aAj+7NcvZ4U8siBj/M5F53moPHBpTdts2HGaP7mutT/Uf73uAV5CQV6CMXkn21lx
KDjMiiNe+MawBgpgHDYTsXHRsEvGyB/bitgkoYYgr58C3ZfsET0zVupJOfAsaSqo
Pbn6vImqkXA4o+a6Wm3NDuTuQufJjDnRWGylT0zUgtYqDxrx4HW0K3Yr5bebotkC
wBBYwLvMBFXym4POnai0EUORTtH0q35UEALxki4FyqwdYdFNHwpAsGPeqUOWXnN7
qEqKWLbetUv4EVnrWXDfr0YXcdVgtGfxPY0e5FiZVKiELiXVr0h3YjdKx5g2D5HX
uO3KUItQCEXNZFndXfhOHQAgiZZ7BAlORrNYhVIsx4oj0QcXLn4Dpiwy4KXFs22/
HfEJgxU5X1j7ylAgR8pu5LjKC7YpgNnifQlCL5yhUWS/dh5RSKNQmBwwPBFFdo2q
r+/cN3R4ZfjNL6FRfJs0pQKdOMHEvxKHiV5E2xYZH+hyGP1ISJk7dUG8+zgBtzqQ
aFmVCLDf8d76H6inBYKoeVIoIq2ec3n38RTgthmFSvEIO2y+piAhWFGVIT2IFics
TQrzxWw898QKwi9mog3nhrUSlf40b7ST5ZrHG3fT9sjmP87lI9q8RKu0X+agaeUA
gpX9K33XvEhTr/JpjhNV1aFfSAxs9Omqnf5+bhDwqsBNTAiISpButa2iaGVSN3r6
4cE/k84aaX7nv9hWxWm1EmsiBN0Ul2wZGmFsBEGY10uEJ5cewYMVLh2qKpHEpycg
I/Q+Xv7UTfO7xvft4mzYS6YtYEQw/w5G0X3o7Ce6A25BqJ5r/vP+shts6+zcMvTE
Wt9OFWo1sXYu+5VynotHpN/s9YWJRPD46ct7KfBDGiAQZJc6yxgJxlWPff2eprre
BNG47iAeALApWH6NnBWosJJamUyvw5jdIqAc8P9MBVqZuGh522lzbPQCPDvo0WTB
AV0jdXhx27i7horve91hMxSBJZuchlJFL9sUUjO/JOVFb19oyP2lgzBHLUG3aPR/
i5A4LWtfPW1A8JTbfxBm3hZL2rG73/lBTVejuR8RiXO2UOaxCSU1EojhK2eNEYlT
AAZ7V91nxvFYnPZ+OPfn26MaZkmgsUIXvwCa0LZ5pLIWoSXyCoKTs+AM3tUa1rT5
5+QD5U9s0V25gGszPVPeA/2Retd31PtcmPjJHUqYCBmCI5nPKc2wuKpqik7Q74UD
6K6L6RbtcgPUh+4FKBgH1rWnCUkNj2CoR38fzvWCu6au4EcyuNhmaTWfic8CJa/q
XJN1Jzosid6O2oyYM/GlJiEu19vq23p1KCBU4hTWRmbYV6hiNV/Bjv6TuZCDCUpP
+jEBjUAqD3vFDln5F5Xk7lDrFgi/WpL9wtNx+hYxgAnRo4MQ8Zat/+6x69bl6Z98
m9H/kKUW0SmJx0LTl42v/U5zpBOWVQQSm41P+6yJxUfVDA4XysPlsSlG5bBc2wKF
VHV+O7v7emR+JWk/ZqCG02hetArsRyYmI8bd0Hn4O8IjwN90LoBydwEzYk82Sbll
dE2owy5vDuJ2lYVjwIxhdMUIvVOEyDEWOGPxoIIM3mfmLBFYYYJot9OP0Dih4oMM
aF7QZY2bDx5l9pyGnG3lHufzT1ouQRcWsrBzFU804PgmAUgHuBXWdFFUJ26FdvlA
VOTrx0gtW7Qq0lbSk7m7pTz+W44RF0EkCRk0mV2sUl3wylzPosU/1ARfSE2SZ8jG
QV+EUpV2J4KC+rm8+h4D6reih0IJY7MIjhDteNH1hIDPQnPK0+zAMz+jWq5ald1J
u907nCFza+uTEOk2Lb9qVJZ8iufwMa5ID0wqtdiW8hygvnJbWnL8H6PhMTAzGTET
ovusKfYKLZtDnzqr66vQ/qubJsLcqU6tLs5k5rHLDDl5+ylLVTe5s6aCaNpVj4cH
yvTlPhsdt+FL/XZMGPkmWT54Ar8FjtbyTTOMYWH87AW2ZACdw9FPakG7a5eEonKE
l+cn0la0E05nSFN2S9gr4EN2xwL1fM74OUVoxLB60XM/HPIOJiZY25UqbZhrTek7
KgXf2dn6KXloAJcafGyxoy9+/wKcoBbKoP5qr/hJujOc+wl5qpjiSQgl+JCfjnLg
j6y8ZyINIqajNNfpCssxuQ8AG9XAUc8+jvShNRVJJPuoQV4J/xCWGUan2TF8/Wld
apKyMT9ZyXorFLlOF46YWkASUqW1sdLvDLkXN+1HVHuVzkrLDBMOw8Cz0SBUZ5w2
850SJMmCEDuZmfmeOJNmA9k8pyIxXL8cfTCTnTMGl0/H+0ghSfKuC7rBpz1VQzXg
Xa9nhRMQ00GJ+v2NLaiad1gp0R/XIEY/MgvgBrb3aEvM4mcj1iYiyLvOCIrCHA3k
JBR4Hh78B2ySkqKXyK8iRU3JiN05zeo2lIyL8aoXKC1iEj/1ZKFanQYXV7ewzgXP
svnV4DG7oNLnt9NEKK2wQZqHnigLeIxtjFwyuyyEZwbxqtkcTUYBHyesppWyDPYZ
vGYJXeKnsFaMHGS07xSjNOO4uWe9+nJx27r/EJOktOMeQ7mBqniHjgfugzZjf1Kv
Qi/0kPUvyJc820HU4mLa+8ZR7aScOcA/kX0QsEGywlutThQpOTkguOcbzlyCL+wW
fSDKwkeRxUASM+6vDQDnUkmrfAWlH9E0rgvHF/OGJUdLzjMr0yJ7aUpUqYGgnAyu
X+3XO0IFd2IVcr/rcMPAw2d9OjT8JHtuag/AgO7JPfi5bhk914pRIDj1IJarYdgW
GG7ypZMr8TMn+7kJJwJRJHPowZhnXSF5eO1KeAWHGQ2LXlJRALipMExz1tD7DfE8
jpiNWgWRyu8MBtnz8wS5DacVL1bOPDTKPIdSgG1Y30jyLoLn+IfpEoljoML0+oUS
kM+Nj8gl52tcPrJnZug/5XzDX4O8tU157BKUOwnkvmUp4NB59KJyYDyp8jQHYi45
m65hc305O2tKZxUlfIlcNBLLI5YV6sSaPrIkKpQF51Yh4JiH4S+gJAibVVK+MOvJ
l8/vqUwYTht/CpecqV4vW8ov1rIXc2eo0fIDeGJ/uhIDT1cpxEe++9dTNae9172C
yKqRfbPeA30XVxnIJqajJu0XFZ5Jbyr3vWkBoFMCTTEEjtdCf8oiYf+upLJsUgeC
HTBENMYI+2h7rBxgKWITJGVqywVvclrfR9uGJ0rHVVX96xY29k5Vv75rwhud+/MT
pILmzsEPeuuiREtcxEXhtGytABzFKOyHDrMeqgzmGRtpnEf0TfMBjoEbf9RHGdZD
K44/TMSAcctgSUd+dei8wwDaTIXAQAnxyKkB+bdwMpfylKPWhvT9CqUGFsLZi40+
QNDSlsDmArDdxjtA3SzDOIjz0Utsca+9dCjx1+iVCVSu0U0/y+pLB8+MuePFpaNf
kvpRpTzrScM9pGmLMFAyfnA7vLH9ghiJrg5hUrsbIv6zYoIxVBcDAkjhx75JLpKA
ohgxsbm8CLuwucEQwkAGWaK5d/ES+LcmBBtdx51xftL5nr8EduswLoOJbIE7aM9C
NYYPLX2nnqRhkQ2Pd6vXdVwRCIaGEIHqQ+kFrUg5rWOcrEl67WSAIiQUemUAKt3P
7LDI+qjEfKdXwYPXgCFiIuiHu2holwae2YW3EjmvGGHW1dHdyjU6YfVoGkc5FUWu
QgIRPeYeb0HqZYKqfyDRGWAibNhxNAwMDvYsDEwPfas86cHGXCbunOqcKacFQzS3
WEGAUtKzdajK9/C1yLgzi1VMkHQ5WrGQbWxvB4Wr+6GYiG0cAR1FFLlbgdYs1f3c
Z1dZKP9paazYbqO65qSyemxZrKPoXvbqrKQJRRRVlrDCXXrpeUvWEPJkGnFb4jgm
Q/UnmYK6esr33A4Yt30b78FO/AanzAlDndoIR1UF/57ht4merA1M6ZjLIUL0lE+q
xgZOkuQe2b/GDvLFUuCDN5sE/JNSig59lEmGKiPliIYkSKgqYs2FYkfPah1c7f6d
m9vZdL2Cm14jthqfar54HpU1OK/u/TSaFBb3bTGkFTCcnhdFlI/2/Xz3cu0fLnab
2GHr7ap2QSMpQEFMYqEYjUC7stA0qW911pc3PbSguIqKSn1yoRboUlWwVNWDDJNO
Ov7HVvpoQ0hYqZ8q64fyWIgHQlhssQLH36dXjP9j877+tFY2voTJ9rWO5Zez4dP7
Mcfalap5lKWvfglwGPSyXo6Dba508W6z4cate54Iq6gfX2U45scM3bVKUwBZ2HZB
ijNtAbx4poP59y4Xzcm4L54WGFGEB8FgV8i/zuCguwjvQwhqMUo9TfcZdAbvsp0g
s5fueaCMB3YiU34JQRKG+K89NGNiZJofgeI95THq5TfiJZ2xsviRGmGy/MLqAJh/
H/42wMnZUg56aT2cQ5nkuliQG55DoHf+YhUwfkxOphhoREJErP86gjnIkQjmf+Vp
/a6DJ3Hmz9ldMWe7k+xXdQk7dBeeX2SeUAbtSlTUGLK0fLjmyZjG97VPjZW7PB+w
m0myF/t7eX6+Wf4KEuyuYiXSlnUA8QkNDFkE9kG2FVDhJvMKzJcGp6Rwobos6GNe
Ql/jtmweURs8ik3K0WVYaLUKPyXKOA17JyIJAkPsSot08rUPeB/IrujBu+O8lZFy
10PnJ0Dhj4HCS/snjS7QnUioZcxPaHaTVfZ5MMq5Lyt4OiX6gvN8FvFrwiupdPPG
gD1gDCHD4/wnzqzP3gp1rqXa2WtiYoYU3ETOZBjUkT2hBYu2PFA2Rdpr8tl0fexq
Hn5iWVvncKFDqsedxcuaWrgi1MfM/VnASg7X2WUnjVm/8uejL0VRY7FP4r48tqfV
furxY2Rl6nUIrkZYjA7d1lHN8TvHlA+nDlsMO3kRrgRDW3C6c21+67mXgjDr3NjP
KqzjURVpYhV0D80cXsA0qDNixn7P2FmEyUkyaSfhyeKN9U+sCmicqK3vwW4bcpVk
M6Wzm9nbJ4oSjY1Z0lEwIaySOpuYHCrm+tLmFxoYBlXd0/q5Ivpcsaa/XBTgE1Au
5/ghNdaOFEhj25I8G6IsFAxT2BX2PR/YSzESSMgZ9xBeIkPOLaGmZgKeSFObWG0M
VksOTXCng0d6RSTwfhC1c+xtnZ1xOzKda3d+4T+/j5YF+nEPWdT5w+Qdp4gLPkz3
7IWJ86o4oj1FyfhRE2ZewojZK1HKq+PPaVvUVsMS577cPwCt87KWKyWdln3Bl6Ay
ZK0mFD2js/viTAYiq/iguQTtmEH+R4vy5bUDSi5zhyKSOoNFdOh9o6Pc5L0O9uZQ
XW7Gtwe5aLf5BKf5kOHtcShibZKNh1t7HZIsiRT1IfRDQNouCt4WzFIQtrY/CUQ2
gahP2VeYA7IEnPJiaufMp/y2UyBIfXZypavT92WI6AEeUFU0h0sX0eZ0T4Vr6tmW
0VoYO4dfKGCIX4hF5k49kB+lv7OTmotdCaN7+3QG3zBqwYEle+saMGUz432MVd4q
Hj8+4dMfqR5tG7eiSE2Z+m2rUlIq1TseFxBo077904988ddFvjSoUTJohr7pIGQc
c0rvootfhIum6A0iGjMP7u6kuFgnQpZdTaYUCsYhClmmRZsdVKeWggxprFSmqJrK
5RAZUCCQB/X8ADsLjr8m/tqP+tKwFGky/wUFRd6JtYnDRiYQoQp0ScVHfV+b+xxb
VD/L4D+5KHNFAfHSy1zdDgq9d18sKzx1PFL/clMjvWFOooQwztalUh70EbLH8Wev
5IZSNHQ5KISKplObkjc+QnNzqDQLYKWlgbbdIj5h2Wjj1kIfb9ZO971cO7p6xcCj
/7z0eHyj0ZOXO9DhgJjcVLsXqs+VwXaX5C6aoNPd9WEBIyTL42OurmfmRaVSSUYx
M0oFp98Ev1BAqluS7YKblR9qLr90BS5Z6ws5p7o3b8FXdNgRTXTcuNdiQYDbZuWD
vene1jA0i2IJHZGhg2q/mclG53fzHtro3WCogjqu9EaIPljgF7pxhkzYQJHB/Ph/
puZ1gB3sF+ldUI3yQg1Xg68arxvTXoidmrEFwmLVWaWIgqvYHRFDkmIvMGHETuD0
uAF7a2l4zh9nSL8iCAsF+H2bZqq3YtKWSHK6Xt7GSPCCQgkSyj7fYYl9H2eBaAYN
VNg/0ax2kB6WtIEUwJRMzB+vh8UIu6a3LQkVda1k0AQHYR2puuX1Y/t/aW+EwqCP
AkeNkLaV6TQEBWIo87nzoG8B3SWB+nVmO2PcjIpI9KVrOusgCprr9ZS+oSrCMNwJ
7WdXH/ztAcxaUJXT2REzSSOFNFQZ17dWFgCHrW+w94rRa2s3c083+XDVJ3FjBrk+
0ud9Pm8SYChCmfJe5F3ohNg8ZBAYrU4Kd3qPlHNpqLwjyIrOpJmHJxRHCZ0kUIS4
pNWC7pHHJTyjSd2QBXg112EZGopORZo8ITX4HmTcmIN8JWiUKcog1Vnt3UffCv+4
QmBqwbkG3eALgNtyuTf4s85gxdBUrKVHX/mGY+jKEoEaVNKhVRpXcbg5mcyg7eS6
NvZizghOIO7960dMOKh+dz/4j98ZZGt9/iainY3wGkcUWsBfrGSp99xhK25Z0G6M
TWFsMjr9SdfGexU9ZkJjm9nlm5+ym62Df5D3DPS5p8u/T2zw/veZVB26Jy+9HsYm
QemN9L5eVYm1Yxv9pBDDM4apO0slNl/FhyLeMETp22lgD1TLeJzHy+ug7xCIYvyX
K3EK0ZMDONYPoTE/F1bp+MmXgjtknkNyvGLz7YnjdYWqI5/DJFUrj04t6cOwEANU
FxMxKRswKxlAGanRkvU1wpsIBhA8DMQr95YDBCTt5T+ajkzZGZJ65bWNxXEZhtMu
Vt240WSIZ+lmni0/jaikqwfejlBFUdFYu+flVqGAcsU9URiglFH0L+Cu5vT8fl2d
xtBVOOt7NFANCaF7DgCmmjBF5EIoHvcZyARCArtA0j0L/jDy6DLtdY3Sx09jwzCi
Me4f/BU5AHbm9t97ffrjcSzGFO1TjVtQCPuU1MwwT4Y/iwq2K4F3bOm0VOKwcr58
Uq7fvW5hSXW0Wx0ZbljGzgz5ZowllYzbmV4Le6XCdWa7K01/4olBlDCUZelPiFgW
MXmvgndTc5PTD5Iiv0NmrWlhmMm5vtEOilBzEK1EJi7sQKiU6VzVOw2yflrogsf3
KcWu86Ajxz0GdJCIY6bj9SBvy0Zq+5yQ0VeEtEaek8STH/fqXPUHmaE2YwzRj/CB
OpzYtmmx07qvRh7YIUu/aSzkadgLw/kW/mS3dyo0gWDLYMp4GpyhNYw2RJCypo6J
HoHLjyoR8/g6I08xCbRpsYMhTt0a2dWcUUJy3S3BlkNd0k18g4NZks6MZ3bRG9iO
UD0elmrnTdfMZRjwoe0ufmPF0O/zfqiy6BDx76I3ttJPnl6qSL8wXuGYL+vsyqJJ
49bkxRXBbCgpZvcP582H3BDaNZ94kUUm2yQW826V+0MdDDXDvv0Jyw5VGlNcTU7q
BYvDMApqR6hoJoJENHI/ru0Xn/fSRJq/KkVDP27Lwjelh5SOId1mPIq6CUdu7gDl
v9+azNKZ7WdxmmdMuJarE/PhS3ydyqVwPUDQhHLyIS3dW8YK28pbPpo+g3A+ut8q
qVZ1HvR030UIbgkAa/bxFUBGy2sVev9R9gl4N01eR5rlbZgAvPtEzfJk4l06aZY8
4davODkmVh9fibJj4qu99OMm3G28ilelxjrT+87j1Mc1EkbfdZiGpxU1Rp92hqqS
qZiaRRdCpcY1fNUw3IXEDrVaNi73h4mSWjvcgdTdPu13TegZLNFILUEnRyfe/iiK
5a7EN07tbdTCmSNjOCD+Si4hn+phDOxKfkqoOfGoZbmA0LhDwYRUQXXtSTT+OBay
rk4fkoo3PQmDtgFAcNbWHG1JKg5uys5/Mkm0g4y9fitOMCrDtGC0GGwUrQ2XkY5Z
7XdT/1M176mrb60ZKS0Bhga2tEuTTcvItiBV0GipIdamKkQ9tdhnOC4IdbaVS5+q
X7aJHQhnIcUZ5TSaD+03TqCJYVlld73/NUstCE5/eQDsVE9cC1KtA6Ls1lj++pWf
n/ryQts65v4yz9IZAVUMxEIlI+FK0BDMjUpf5pVMEawtbi8Ue5X3vW8/g4GYo1HB
TirC1CD/INTZSchu/+UDkeZfemt77LkNBytNwOHnSDFDREnCllwJauDczPu1S4Ht
lz362q5UsAoQA04OLvKdrCAH2Tlivftt+XYuxuM7KvFnQYw+VzTNuOg9pVt5a1iW
TIzFvVaXTp78g3C7FZ4L3urtdHmUVuv82eHBSj0Y8CgZn+c1P8SNGfFfDlKGThjB
ad80oSIorh5pCHXDZMbkBrbyiZ7b2Fd3b8TF+1j2JuZ9NuJpJ7SY3fgYt1/gC0NN
za4FfEVmRNJveTD81XSRE6N1TO1A8q2QJU09Mnq8wz9O36te0B0vwHwFOwKmJUN2
nRRCnas/WFYwWjZnzV6Gs74Oa5x3jC5sEtW5CNP3+1rPkFTkYVxXqe1eCGbGdgvg
+rflVWIU9FJJTyClIjCY+EJY/iCctjXnjYUgKF5rgsycBhFW2lJgsDTwFG7DmlhX
5HUdmL3yCWaYti3iWyn/roPOtLzgb5GgI6CwO/vP4eOzt5tkzcNRE6R0FznPs+UB
zzBKs6luFbvcybzdqceAAFOi3s5bKZ6jXhWMPNsoUjjx/FSQDSQR9npPNym4R+NX
ebpkPcFksDcTbWmER6hPV7vC6icuaaMTL0oYSKHbwgKVs7J2TEprfqrH30B9qNwM
cBB6wRgvl0YjzaZH5eYs1x60SrM533DiOGk/hMXZbYy/Hp+Q6U1QDG1OuJzEW7KG
2hgc45FxyZwaLxiTNOunJ18goGEZr1IQEjuwyUU7l5MAaTbWjS7MKfjHi3Foj9bo
wgccIfUQs2FWed32/bfHMciNiOvvOGQYPHKPi5Cs8eDII4NTKHfNu+FmvHOJ0Baj
pCaiOuBSWCdmi78Hf5WHG29RJ6ZJ5wKmVqbpAsJq/HJWqS06YkiVi2tt3XPMzh3d
MQLm9zTc4Cg8mY+LrM0cLvkBWY8hzLAHOWm6ciSZD+cgWVhS3WAQaSdcspjMMn7F
rZkVBEE7Pmg2geilT0V08aMX5wEx5zur6RZfJ7vycAgWg206J9umZhaPvLKNS/Ir
nuadAlyuqAVNN3fKOnACk8gVEkBHzZKzkmKl5sy5/nwimg9R51f3cwv699k8zVPE
+iZn57oTZBucbgnXrRtEeC/72/4NBYJeVlKur9hc0k/cJ+lhlaBHyv0BEntihjsy
ZhYh5+4u/PoavYutGXjP0+UKr3Ty0Hki9Oc/wMPYXEAmOFehgzrsyGDj04ssulsp
oA2rv3I+I+y4yEaIrLq3lOeJKTnFnenDHT2oXbhVfAGxqHDvpx/0Nxis0Hs+ea2e
cEuYg3YnKW6pqTWt+VVzYYug112hvSGWSHiDyrtnd6ivRmOvz3ZLUV+hsSEUJcWU
Pd6E7FLf2tZiJpkJtUeBu0MtB4kUSQKA6UY+vvQWfs6i/xlz9iNzPaWpDaRyH9VO
kbrSZtFCVXqr7iR6+g+k/HFtgtYy9duXZ+xSBop8X9hx6CIHwFuYJy3g1AlJbBF1
kbVEfPmCCgmZ0LV4bZqu6hbUW8iqw9t9HE2WHz11UQRR3lnhUq3KW0ML/g2yDjf2
HdEb5jqFYXO4CDMmjKTBYwpmXymNXU5t1+ES4cp14GPKlnSlMAri6CK6DcEyl2XT
g4p2N+tdnpkTpCmFXF3ejC4ww1HyVjADpP/DYys10ZCmrl89Gm9BMZ27cnM8vHeh
UCyZ0T/lnxVigm7UABRzBpBrtwDiKjirepKFSoSUsqnnjcxUGwH/m5YUmF6lxqdW
ANIKpq7jXXcQpf/NCviVCAlhX/x/JFD9bDP0P6APZg1xIaf5CTqiM8LrLbm4Xh6V
4psfWWehCOrK/m3u227dxbTh6YX4JXjdkWSNqmupsdBFMYpAB43ErTxmLttEmce7
7+VpVi24U/cP7eJBrkEyC/eZw9pnLZc35SEb1d40YjvSzOT6aZ8qrmjo3vZZk4ta
Azm5MRPc4ovQHHQ5BGTHJ70ihY43WeOC8/GmN1wY0aKkBK4FOzw2Yp/S2iqUTg0M
P4QvYyX+9XnU7DobwVfP/bQTlj54tpLeKCz7DdJ69H7DuZ+Q1+4fsXGJV9yS6Unq
z3B7tmSMxhSnZzc7nd6JcmRqSKfpOHKZXjK6HezsBPDu7L0587JSDrZNSlEpK1w/
LeeEHujwP0uRdpDtNbo1/sp5FKSe35sSoQ3PWfZkeqJAKynU1UK99iumsrC+vK5s
zYVEnVVcJQlavqQlxOZml/epfEnpo3Kgvv1LxIr70PSyXkLgrrM+t9naBffruA9h
ougIfSGvPzvT5B1/SvKeEQArZxW10l38cFcVZXM4QjXcc3tcG6SGNszNRie3/Qt/
vtHHJ17FMBa4p0ga6Oi7uQXAKnaJIiFNcLsweVILUIVUR0JEW03CcTGMrCGt6E92
A89ANQi16rLhHLnBLyeGGaSAHne9qFXBxNvIAEcJ/ksmMYH/p6tdH498WwtIl7c6
e0eAm5VPPnip7rfU0KZYIdrUUuxk0G4Ilj9oonhhmslQ+xyrFGByWqaKEE7Hjhzp
GM6YdDAv+8SWhV3UAyVahoKodL2tRF8R5AjGBLP21YxNwyQtXiauoLp5GLTNc9AB
Zh7qFjpT6HgsqgyGpWotzHiyA/ZKioTeMhkjsQUb+qpnsahARpMx4dafgKM+sq7p
p+TjLlxcZoqVMzt+NaWzkF5l9YC82cND5nqcUt2cnb6+kYyZHQ5vGHvU+fjVJ/yA
nsiEHqgQ6skhorwfUWDUJRA0yXeKx9OZ0GxrTxb8SNX0hITCcqlZHu9XVJbhCe43
NJPfP14L3n1V9a0dj+9MuM8rdRvgQun4oc9On+ZtlbKXmMYlDf4aBePUX8ZER3A7
IF5mra9VEH2TJuy9lrbZhlORJjUTdGvcwQHySh7h4TQkdM2WeAM4yPtIN0ubtgIt
Lfk5cdIRTR53aUGWdKAmC8N2p08fJtu/TG1Dvan4qMpqa3RsZKgUBoleJnp4yM44
WvX1txBhSOuBgtsbr32LFhFWtG3R+SXh1CY+hBEIkb5tdjs8BE0CHasiilfXk7BR
mkO1UZhYVro+SFKFZGuu9iX95IypvdyPV2XWRAUHCwV8jE9Sz3tS2nuT3D4F8vI8
qaIA2zfERZRaGCWwKdNjvYGo31VxDrfQyf1aHV9W3o8qKZ/SnA01o2huN88UPgBg
7HNbiRxGbvgJzTO3tYTBt7tzG9BpDPLEiHb1Ya5wlcOOMKvTZ0m4ET9iTbVGJg91
t1MuVIfaBYLapuv7N6NHq1rX6Gfh7TusMrpXgKZmR7DVxEdHH930GUQA8OQFERXf
uFUIWNUq3GnGChP8Dl8PJtfYqdO59bNZ22O3JeCmDY80hpAmBhcpe+LF4DR54LYv
4vLc0a7O99Pk+EVwxVPiLwSn6dHXMaTMM3oWVZIUmHMS6W067IlSDMtrvc/jpRqj
NCA52bCbWPGLiEgDbljHLHqmYNs9NXJMy98fg4ZC5DPy5xq8GqIe90Rh2NBTT/HX
fUb6KaW0csVpCt7ktbwOQdAHOi+qbFVR06kxnVjI6u+vwz5SWA+PN5gyP9qvfJo+
NZQJcTKlznp0Jd15JcuS7AetBQxKAB3EWVzWeJt6R9EVzG3AQpyYcQbXpK+8C6oQ
6hlfzZgm71ka1Yv4G8GB7PpCMcG6fgJclwTBUNKFAKmKZiQ/GPABZt1c1ak00nZI
JYSnZoxQBf6pdPjf92aHwa16AT+isU1ArZJmVs+CivhamFKFlRbUp+dN4FQizoim
MWvMYDLS5tCz9byjspKJB11/FScPSnJQ7Pu10ZvUHi6CrU4M9hMS18ejU/owQggc
8OUTeJhW4+NGAItRRfzj+bVU+pBxejzHrP63Z+c1lkC/6cJ7rwogz0gCsmZs/EJ/
hi2mjNNSWxDyEGVl1Qq446zTPgRahzBsMHVeEFF7yg6UPBAWR65k7caT1RPm0XA0
FUfAyQTWBBxMDVfR+6JEWa1eHUYXvyYH4UPXGYDH8PwPZ1eYUJmBhZME2irdNwWR
8Y7AHFai4oyDAt97/xvo0n7bWqLj/lv9+TuKmNQBVAB08++S6eAeRmC7F+eALyGN
RAQXgLB9i6e05ABF6/R3NkWt8qyvgsXgB77qxUPexC8na93GqivqhvHllJQ7P9NG
pOllCYY8+jxW6J4TdW4V2rLFjKXOsEuBjYRvT71RuZrFPNlEmOYSeV09buiJwnOf
vyz7IWstQyk4w9mF02T3s7BdKhDW/1cYE9omwoUXSyIr+M1GVD4oK3BE/Y5QQ5vz
bn3faMSIJDqUEYlQpgHIlTone9H8gf1dWgjFDEb2mp/pARq0HEowlunyM8UHv3oZ
cahAgTz8VjHL58RFEWnqTCo6jlB4Ur5lphScuJ1xXhGBSHwKqnl7wBda9zo7CV0b
wOwL3nuKNxGSNjGHEBo7AbcJN4c+Pg9mm0D/yUgD2gwXfd5VwJOUyNdibgDwInwk
nab9UvFMCtQWcFyUbRjHYIYRCw4pZYVN7lozDN1YZgkW+6Kk3XLCohoUyGCCGeA4
AKxbe1acaxoaS31PK8D65s6VhSE8QTpbQIUnpVjH+jcqvz/GdFfL3iIWIV+den2z
0cyV3/jaVU+cTNfZT/YyJ0c830fBMLUD3uBZRuIxxCHrBWQa+P8CM0TLCdrhqmpu
E/obJRLdHgcWLLvgDpJ+vGp0I3k8NzmieEwjOyIs1+56PYhrtfjo0RgABRLNHv/8
6w7A76CuI+4xu9Cz5lh9EeOgc1D2vB+Ig9M8L8sxdGlGpOKXjKD8xkRt1GL+FAwS
vDjpjOTvr+6rHsjuUVFon0rCNYox0IxK8E2pJI4Qvxua2xfehOuq0qfWOW7fG0hu
pxROlrtZtAZOCE4APSaP4NC6FLCj3XrbzeG+eZNyjWFMxJ06+KGG7oZl5EplOJhV
REqQ2NvrNjaS7Jv+rBidHZjkwIv8L5lOKg05vJ1ypuaB2l1lWARpHx2FSsXR6I5o
P/TYXBO8D8d91GGWMeDEKLi7szj0fTQ92ZXolPQSxrB6Yzcl6zbEjmUegBOncf7G
RDGgWB/fTCMSWOi3tlkKReX91Btl1vJZgZ9cagLu+/yYSPe398uc6tAYD4GGdSjG
MJgLodqlaapWAf6U0lAyhp3rdOflTAgE6Rku8KT1NUZcEvo4FHKyhg1gfYRDHP3u
i9nfZrZ3Gv4gazoxMoXDClUwGu9Wty+WoYWkkDPIrpjiDdWnQQx+1aCJbQmCv0yr
mC8OfqopaEFTELdp8++2Hx01wSopu+Hv/FUs44wpobY8Md6fhx/6ycNieKAZMoZI
GUhKBAlrqiz0vqnrBaDTyJ0OCBjDqxGEX7reMn5W1iCcXaU8NX3dw3KWQDgVTweZ
y3vPaZHaZLM7iBRNYdcAbPBJJkmq4EWdKoUm1YH/lK845iaQixEbj7Zv8p+oGdu7
Os03/gGbjjl8HaCJ2E/UOZOW1qI4V0LRklYJHwTux+8aRNdOaaHPunOyIKeXLA5p
ltzJPmVZYZjHhoCxAxocI383Hr3pS3moiEuwTuYoH8kx7e6uGUH1bNI/Y7lGfTgA
MbYFrYOvgjZqC+i93Rl1wNq8XTGs3emU2wzqc+wAA9ZTxVx/bPRmTsf47Os7DnrU
pWswxVdZq4jFTnVEg8HLY1cFQ2IfYHVJZ0nD5SNRIe2jMcPBRYQYQvg2MxanRREy
rju6XFwoR2N/uwsRbPBFt20DJYFpP8hY6tKqP6P4hGVNCvuLeJWzl6p3TFGMPAgg
Viy/lf+to2AwvD2C/3vh7kCKS++EAFSAnRNe3iqZvst+Hz8kxOJcE5izdcGYwIA3
3nPfQCzDVQ0BagIWwNDVod0vM9gL7cSFWieV23GD1nEkdw7XmlkLNuaqRYdEROpe
gVyDZmTXIX4edz+TghmafdSMwNiH3zGqQtmc7VQYO2r5TqwCRlj+0CFPr7ERaVsC
/+ZlmXJavrEP7Kg8AagLh+Ca6FbKPovIgfkKqed6jv3mKLftzG5IwjWjwcZCwfxa
hCEXbXe23czqcMqvQPV30aomLb2SNAFR2MgL9cWtN2VTjWCYpuOwf2jSu+/oHzgk
Z7iI6aoo9q9aNDn5ShiuV85ZapUFKo4A1eeMX6oEvpf6wRmVDx/xqNZ02fB1Auqn
QmfMkK7dWHTA7s8NqP6KqDTuv5iUYBcQjLxvqaAT9l4eUJnSkILd11baKd1PE8W5
iMNv+dQQzRgE1LObaPrgySjdTrYMrvLDhY2MkGN2ZxcJt5zMVzL+ZvSt2Di5ynVZ
DT3KRBnx/Qwit3t6XLZilJfjNVK+MJfu/+OBqqHz8plDPXJvR2JpmdKz+YU7HclD
pyrDddypgjjthF6dDrR31hUq2eAdd4UUBOBiMt8dye/XAn+jODBHiyVdBadPqokl
GMZikEfKRoCD7ehHCJ61LbetSUV1Z4t5oXPfeLPc1fsrDunBLAEfR0QOzqH2xZsz
m4Mtz3LF/i5S+1La1pZiZTPNZTho6SeuNqGlcyKEatMsNxhD+gkWSBL1oYBd7UEb
/C78TNGySaqyfjHi/rZRAgIF4vAORqTjdlZrpWhnuYLV7mEUkNXt+jH5Y0nWk4Hp
kwMywsqtO+vh3zwmnfL97xTOUE+nyP5TTcoqkR0NSe6j4UdvmbfLrtK/I5RETeQG
TX2zSp+L9Ruh+WLOA8MRKDkghiTmE+2brExMK3ul5HfQ9R28fQE+ZqRFE2CsOQ2i
NnFck4kI2kjsWkS1dmRZHJMrm9AUWHIwucsM8QgEWJ1Q0J2Y+ZhkrIETvoUIVKY9
LTZDOn0ve2PUdEcxPcwf+GRQQmuHC9MUpYdozafztBPV3JU1peJ8ruVrOfI7w0lw
zLin9DGpoKvZYnx9GzAatD3Z2xW+6gCzl8rMJo4F6wS3R8ALrIjQ3rZu9pRGSqJW
Xh5x+DTQ3YPIwh6ZMhqiqA7s1JBkHGLXJap/hD701YTS2aEK85Piwlsj3iTbMcRZ
aSYuYJfPmrmPJUQQIU9nL9apYEJxJLzQJO1Z0UrKsJ0I6mmcGN87cVOsQrc+FOdi
yS6M0Ajsqavq4BNRA6iPDHxBKCIwbiTOgCji261K3D8zs9cO3SIZyTzup693789C
UMMNqMD0qnxyWqskJTc5KKxPoCXZrOmztjQuCoYWSuI1XqRA1HYgcavjDq2fnRTr
RgYpFA9p9pivoos6Cn497m2eLLj1yP/bL3JY4S1d7hqC4g07rslXm7Fi/bcPrWEW
dIGRoH/STJRTmAW6YvtpmoQRPTwyDXYYqGlQA4Ax3wrbc/XFHJppum0nKNdZVFiF
TeFSeGHC3leLZ/cYQQJVjT7ra/GCr4Ya0E22xdvN/t6tYctJOosALqw6rWOvWxDa
gw7OSfDPiRcMWgZvVqy5CPkGtuwzieoGsUWFC1av+RmH2AC5/9ymluNNyz9tBssl
dDmV0IJVX+fxjeK6Y0tsSPxCobpNR840KjuY4kOkD2btO3a68eBbZfMKZ7BP+Qg6
aiJejVz55VhwjQaSaqyGl1HjnlWR/S0M60i6IwyehqEHixiaWgf9btwNFp/8rSSW
MAfkvbH10kfxT8cdVHNJSG1t4AOlUXjp5PBPPaCBo2usTf5XyFbYORIWiPlwGR80
smpNyu0wk1mxQh1uOMS/N/ODQwESKlqG+uiN87JGWATF8wsWKkCgQlclyvdXDJdW
1V0HUR8kbeQWYEGC8ImKJ+gHDZU1ssg11eyDIzIX4pJSBTLKbge4Qh2jI05BHVqF
ifYUDOyb/DRg/XsVieoW+oT9Al3ojiTxDt1svvKbCZfLI+TRwomRf7UIMNVfa0pN
qQ6v3QeGMDDc/qjkQ5+zDo6+kLuexoAL1k4EyjpiVi8bs2qQXuLeYQ3X7xwHNgdm
r1Bb84Z9kIUAi7EEMqburw4UJWR/bS2I62iE6TCBxdgnPEB5rNXe/rHw/TrZdkj2
RfYP7A63MTGRN1pL3B3nH3khiWQy+sT4DGYXipWH5KkCPWFWkWIS9s2arkyUstVG
6+GZVvECsUS6Hbqmcx1h04KmcMtcTkZ6RnOELhhb7cNCpDRpXNo2wvoMj7iJ+cSz
McNpXxCjFLqYgVRq4MqF6h8AW6Z6ZMjG4PDpiIzTGBkojCgynWEh1iu1ZrxLHKjM
7ddrH3DWzbNsA+qectxszVxSffp7AtTSVOecinct4efkQ+ePqOdl5f573EUBCAJk
7e/8LCVRiolBR0jizzfDJvHfsQS5EKtHyG/l84GLhWb9QHVKcpJlpFXrrqEKcjog
Zs7c/qNUdBty/fP4RKel4AeYEnEi33wPktMp5CBy7/WcWY9Iin7sh+sov8sSTQJ7
XRBY7xxLjFhKycKGYEqsdfza4nIrPNMEGIyM5Z7vYltbbgj3qfogKrBXMWr2ZMcR
e7v5/4wX/8Yp3BWHne/Gs++SjTuBP40Q4wsVsn6tlZ8q3kzhD9VdAgohx6E1Jugx
uS0vLE9JxarEdnuNi6en4vNnvUMfDBlHIoYdEAnutLArnCHXcKnPEEePymL276gA
s5+mZ0RIyt0I12Y5X+t6Msh08nGGYRljffFPCqiDAKYKxkYln/8uGuW99spXvxzm
ahGt6MRAcTZ2IP7e0xSSGi087jrr997R4Bujw1RoEMMhcwehg5CGRCQX5BzebuDu
coqgWxAQSACZdgHR3FPzYS4lpd5LTcZpwsbNF/gS2Ww4cas9Nxonpd9XwWrHOa9g
qy+mZbou1KMYNNvwiGPF8cUt3bEIi8C4oxDWPxtErwnuCg9d4K75Ma+2jEmeoCdA
O5u/yyujr4jXJjE30kwz9F9rLlMlVsF3aGZa+BomY8K2Oz6leL6xp1vaCZNa32ym
6LSWbTOkPsi9yeB1hGdXvRK/RLNyfRpHB8ReP5wnI172Nk4Qqd0gkx6LSRObMFOo
cbNo9x3kWr2AgYJ3P2QMRL4OSiAh/WYsTDUkzvu0sNDoxGiXIBnMqKaUNGXGF5uq
d7OgvOzJRZyjADFtR6dgUcD+AbwF4m0l8wZedHSKYhU4xguLgND7vmJFCtG5X8ir
JnVAM7cAqgXwCKoylkHsUs4G3i1OBGIds+M0NHP49oE/II2xxEi0ZLKdb4A246Nm
alXDxss5bjaHGjOO47NZR8WHQ2JzD69P9egnirFbKeZTTQPhKEaZiINADBMiZaCd
4kcSVB2tZDYmTTQbaGV/X3hm1dgmygbJHBHMzyMPcfIbsMSYjN8dF4nFncm/mawD
jGmbUfm6fom1BRRhfLPpicHJ04/sscxR1CWi1/yfryaWYurQtX0roOCYy8SeB+MH
w8ElE5FpJD9n3NivnkLVj10uIMA3V13T3LQxNdqSoX0iYA8hDs7bmHozRqO/s5Lq
2jKu9nYc5Pqt3u/+Y9uAnU/G+6l+gp+EGvfhdXa5YdpuKE+Zgj/KpXweqUqqS8BS
E9zpYC/TpzZOFGsk/iyBD71UaRZweupTku6rQqEm2bzg6v8g6pOJcp2eCE6lMlrQ
lpzJdBPslOuz2Vxp36ycEiLgmyzL1EO79WBf3hFDXgzGK0GnbEX9H96wCfXqb5IX
ywIsrfBjBLp95teZrPz993CrvVEtkD0HTZPUpdbGMzVM8+kjDYws+Xy2BWkRJbE5
Zz5DjhuYQCUeNrgEj7RFNdC3c7sDf3V3+nsIkB9h34ZlmgJW2mqkL94ECMUFURb/
3FjrnG3dvixQGNIw8XUrAxH238gAeq0TvOZOQDK2r7aX2mgumOYsI7iPC7bX9MA8
eKRQF3MXfCuiYQPnw9kBaVEFeBr63z7K74++6uvwLp2+AT3hmqT5F905O2JLHwXP
DhUTaENprxFG5CMq/a4jhyCr6rIIfNmRyY4COWTdaEyTjU8aQbZrb3Fs9Bpklwi0
p7hUoauvI/paO7CA8/+wwBeuc5+o6QA5KTHzKz4lZKlKjWRfxIz6VLAhSlLPPHSh
9bjJLRRH4UPkF3FzEe1lIHFbFAxZ7CmrRM9mr76XFrCn8YBbqklJdcxeSei5q7Bx
ZFYfJ5DYd4w61n2aydVjXsV8jviOur98mCPlRaq6XPd2G1XBg/HU9t6zfjWzq7ni
n1dq0aZIrcKzogzgNvwitWeYhymdF47c6wCeYYiD196MPLSgaIYw5FAOSR/gZ20b
Xd6uRo9TF5+yS9GCwwuxbMPTn/XMQ1sWlNdjbvFtUzOeJER/x7+/EOnQoOPy9ObZ
ssFQeQlGz3769I5wMuKZqWtk+1xcPBjd3oqgHfkaZRe+xb9J5kuCS/Dbx2caHhW9
UGxT/r5zzmYni6/h7zuXK1mSbSq2D7TEGWFcSfc33q1mkU52o9mRsC71c/NiP2Xi
EhQIf0zAYgVU2UPNecPWGuS8uvv+SkaE+yPmtdBOHwNChpoMIvkjOaq0Kcl35XCz
ls2+dX1V0Q+1vTWGuFBvloh/3o+HJNO9clXnc2DYi8kvwWXTYVoVsTlru7qaqg5Y
M9HsYcyXP3Xwb67Cs1/YCVhttLc3KJlwzGJgR6b0GXWxS6eCgSIrzBlOeLYxeEE+
DuSylG7kpChCS6xcniWUn8TmjIDWbzAjC+mRYR2ZLf/ZXMJVHJEFp+XSOTARf1SJ
IgTlJ9T8ibBNQKF/HDDhvsttHyk7W+uxjPYekgfs/tj0XLAhKg+pUeuEHdxwtgz0
MUum2huZ228Xd+NTaPcfiIWLrlzrF0unRtJcMWlbQcCwMX2iPXGAiYCOLtKQeiKC
0u9AtI7dUEVZpP1lh9eCaame+TI1hJn0dFJqNwEZRFBuJiQv3itl8Y/UmncDSBTp
Xp5Yl+wjyJ7v8a4uw4GZNW8dsB8n/+p2/KvDUpyV9DUuv3UySG1X9mnhVUryD8DC
VJ7mrnYYy5eIN5G2N7/xYe0cmQ3/bSZfgRVASTJIk35zY7WiFAPLhjpB43TngOWF
LeKo5jd8J0zm/SWJb17Pf5bPktYU0EtfyBybjqAA3ltAsV8WioN81cmlgzUSYRxy
SLMtjVDfek09VrNqWBSF3AZAqZx+0mAgisSL2IekYAoOKUn+kN+LmTTM1QW0I2+N
YFw/DlZ8VE0DUm9l0anSNEvssWNvcSsjmPEmH+4CMtgPisY7OJTgRMppOBz+r0yP
xhXrZQvsr2e2ZQ3wq/gPJWmxuowGdu7xxS7B2EdodnWFcnHQAFKmeYnipLn0dd2w
rv7JZdiDoNTrNDKCGs6u+5a5b5IzhW1WBihmirJavdFNEm/rHausmEXber6v9ZFL
6wq95x9duDWCPuf56jE+BRqhiXIPt7m1gyGtqbBpCH0wylGCBC1qzcM55W8yQC+E
IenN35fqAD2PVULddC5c0VofgtDp2l8JL0JD9wwK9TE+Aw+QrORdNBh5OyQRF3SM
dbPjKRTJ0s0k/Sx6itxbuwkGdeb+v5CZIsmqBUbSIgWnUqW+DsMpq8O+NoV6xNQ2
e4h8HQDbyM3NVoHPZ3KIx3dNEMS5opGtG9VB5ZZ1u/DGswCDkO7uNKXxa6I/lR/k
yeBkqtWzD7SvpGS9NPrelaj0a3mKeqSg1DXCHq5AWwP5tcs58fddSjRP6hPeCar/
xjtOfcR/0l9A9rCv1IWnK8d+j0KuM0iMEhYHWYjvIYWWDLJ2K3RtlNUipGxhAFbN
SY8Gw3WuBELeDDLxT9iG0aHknXIZJZlEc8f6K+9RbozYshM9oaG2zff6XUaMU1JU
5QkDiYHPG7kCaTNBHPtiwCVoq3l1sroAGdDRCaEiLciFHdwgnUl9Ze8B128JrUzn
9jcb3RDUlLthQje9cyq5MSqqGQlrDziYRKEBH9SndCVe/m9tNSXh6omleDursbnr
ROqPi2wpQFYMda/XXRO51ZFJkVW8R2nZvKpmQinwkYhvBoUAy9nvy5p2Fd7HA3tm
eee2uhLoBHfNkf4pfaQ3TrJmHt+qlUS4qP4wXnKnivxRHYpbKqH7acRaP7+7h4j9
6JUSE3jTFmmGCcDNRx7nm32X5K9ZFsLQc7U25oTbuZA9uOamqGp8H75sO2d8odb/
bM7k3BPua4+J3Jzrvpu3BKWY5hkqBaXloTlmxhuBBCcidjesbx22a8/a96q0Rlkc
B0Fw1NBLuafA6kHmYVXD4u6la70qfG52fcdm+yecL0H+cz97o6MzcTW3NxgaxY2m
lCYlIvsJQ9XfEUMkUbOFSv2j/maBrzTLYgIczCTZ0RM9NEtaeWPn9B0KB1ftLc29
+HIqsH0dWNqSbn+JDQcpCllk2CWsk64oMJA732fS8syKrAkvyh/FrHksbYFSYGdN
NBbFzh6jrQ9K2gV4OFLMOfPwgtJ3v7MZNqnsv7YiUB7DRNFYj8iwaH9Ls95Jgcyq
+6o37FeDWf5wBz0vI+YYs7iFrloCfSr0fWfJAECLYbKaLTbgHk6FJ7W6qlYVFnd2
aPa2HFJEkfW1ok7mTkNjTX5euIDewznaW3aX/VN7CMph9L2MXJ/+v3eYqcBFmWWc
XbbGRGJr76M/q0YPs6WtAVrcwnYJDLNKOlRJSTAdX5XXg1CtGkfk6SiVfLjjIMjV
YzO0nPvW1F9teTZKAih3xD761X/42G49AbyewsXft/U5RLuZ46HBuMWJIg5c0fL6
VR525WVCaSIsw5zvpFbvYdX2XagOTkcQZehD0gZtm7NBBI3SC83Xsf53mSvqlCxL
4lfeG5nlWV2Jn80vTt3gF4qAg/EwWhQmck/0dRJ2XA8nhI4Yh7MeiyFZDtOa58pR
wi1h0y0uQ7TSrNlMYUkp7BJNdMLMTiJlmkxvfoAf79oHuzBOQKRlwjRy/VsonHFo
9yMxWyiPj2Q49Fd80SQvEpcdipa1FrtxYaZLo7AjorVQdeAW1eo7g9Vxm2ICOciJ
WPd21MGEtm9xKsfXBihbFfHHJPGxe2Towah3KoFO0PTs5fbs9FBJuINy/KdwJjW+
o3GHnwhrxrrtvQ9MKC9TMsnHqAJZkwPMagSqx8VUJ9dxLtHIirAkcwzwxb3TXMWI
JjWTkJkADdWm8dh49TmTd0XHV2EOcWqMewUOm9OQgDjio5dzBjRWCiLa7okMl1/w
XI1qWoocbvggPpVv8lijhdknSGwgivkIbEwAV1zB5E9zdF6UIf7YdHjTvkVGZ/k/
fn65Z5hxmbXOe8Z8G1O11Fprah23hFXraQIz4pOBCgD2enDCo5HZhEur/vn1iCH7
vDdlDhFjaoj6RgZEfi1VQvtr2xuBS2DvS/j5UKArcLhDz9d+X0UoSqp5oD3zyiGi
UCQgZmoz71H/SxaQOyOI1gxB07J8yYInqjAQM4ON7x8Kc1IgMXhWDaPGKdq+6G7a
614EOnXUYecfI2ZUn76fCe1DgyHse4MCZkBvy/s0iZRnYVbND67BkdJjnX33uVD1
//ducH5tI8GKVmRh6pnhysFCYm3b3ERUaeW59cxDfpj3iAsUlP4BsWIloAqNj7g+
uhR77wx+dTBWKPgF47m+NiHhCFG27cbc6tdMBE0dFOpsT/1bruAcTTwVbrVphZWI
wRj5Fum2wHJHON/4DX27LAqfBxWgS9AifWnSo4o2mifQwVzIuSNsTu3BC3WhDfI1
PXF5kaQ+IPZCs1cNkgTtybznilz9Rm+mD7vpCWrTGaXGZ2rw1g85JwtZ6BivtBCf
WuLnyuQuswNgqMWfWhketEoULjY98oHuSkCpH3+NUE3ZUsuiebKzGh4zsjvKJz/8
lYbAufhh2TiOcFPh7A9QMJlngbW3Nz1eNMube/4zLLTXRe0twudZjwLU7AIZGCmb
FEGC0SR+6R9wdxh0MKDak8onDX/+jC631wLljHy3rv2Cl+w3fWd01emlRR8Du0oG
RIBocWxmuRF63hzUIDv/jwKplRdHCtgRYxZIB50Y3cNt4VkFsQahe0vLHRQbBsao
begRQK7kW99ORbyWJlws5uUDXeCsypvWLHMVEvJCtbOgwFqNvWNZZwaOqZ59+ehC
pCAhM6gypIIDYNJ1y6OEmy32875UNsp0viaGXfjdvmEaLuCbfC4TuzpUzLDYIsct
5zRMHZWkWWI5GNJtV+RMeAoUjxjizfzDUOrtp2yBz6m3rHw4GfzMpirqZrqphpK2
jmP8efjboOynm7qXYhv7NF+VT7LV+c04biobEGwSVLK/Ee/X6bLREmZvbv68HzCE
pIz2Q8xnIRrQTwdjd+eN+cYik4+kAQTnWhimnGID3Mg/5tfD04Q7Dtdx9MMuJNdy
m9+w3v794ZD4EUID2z4TaxQTJ27ijEeyeoE9jQQkypHTdv/BkzB4TbXCmKplHE43
FeJLyrHkfrMKlIc9bru8iXUl50MajjbzdR1P4tHYD5eRW0c9At9kXrlpbHtADICw
AARa405Yer4XatkSrY1ad9e9zMoU59M3hI51W7/h84reAHBcD6U6OOLGzqkwZftZ
hsAWrhrhRza5LLn8pJMXJbVo6I6xQtJ9xuFrCN/IyplJRxUOk2g2ldrNWHEr24Ix
XBKDael1dkS/taT0Dl8KE/JRnNzIRUsVMbzSnfuf+W1rANLYXcrO8QbdctdiOCSa
hnWySzgQ1M3WOpxM7IHeUqVB7lRE/T+LDraVBYbFdXK9L6+MopnSsj246CriEDCm
jZZvyytGeV9AgmsTIMr+Uyqcxsmtkvws28lSe1Rtqf9G1R7leTfTw1JXtVTfuaIk
AIyB878d6LsV/yYnxvBVeO8jEhw35YEKS/SsSUBkegLIDV1jP/Hzf1uW7YeKYsW7
qqrKP/ADnbMWerSPKJQmSCs1ceQMRua3/SobriK2DUCG8ngN8gGk5txfloVNTccI
UkZURx2QEk16l12mZEdn/yZTLrfoJvTUwkNQ1a97efvOVujh62U3s1MkR/byvYRU
O3MgdeY87v+01Be2rQsm6opfeLR88gfrCp+m+PUOFRldX9Nt9Xc8rZRQjoqfwa1L
7X/0aw+yn7/kGGYUSbZzoxvU2DI3sFJ/glDu/8vfD9pnEHMacrJunO/sBSiexr8V
FKc6PsmSDqim3xbWNEosdRaCf84l9RbC0sPMVlOWYBSw8OuYqYx4x45hme/zOgDK
+m/RFyhHhZgPU74fCXBB1kjzwc9mwWZB8oki4WtM4RXY4+gIRNqnE5FUw9jBuha4
ZsEDNUQIPA3WyEf2QBTwfjwGgLRP83I0zsuO5Xp7xGZjmH+ZhMYNNNncseEKEqdX
FUvq5HksCh/+JasNk5zhiHhKW9YxjCNuIBwCud8KvOXRGrtyP4c51RJd8JNbEHLy
FmnH2q2XQKvWE6VNn8afosIJqGs8MdOuZpED7r1kzt+fld6W/0I3LckRAP1s6tzo
kpXHL6Jq+keKVWvf3OcwzxjjjVn6Tade9p0drA16kjdbkBCTbyHYqo2do+0M0ozE
kai5KrukkNClITYOtK3VWxXW++FsVNHZoBY8z+yP6S10nQiL6Q6ZRMZBKOqdeFcK
Um9VlNGAToJFy94UwOm2BXmC2RJZdiF3jm6sY7gpSzeoRpQaGvDp6JHuYSM7vBMT
6RUqL0wET0W49m9mO25LD4bsADiWjU45wbJth11og+fLLw+Qnb7r5kE9p8hcm0Un
BKoxSyK3DrEz21o58zQa58h1ssF91xJSbTvmmU21Y24ZmMT9rZNvROi09VccUCyl
wDb9wl1UxvkrfTA9DDxexxL626hmMvvyCrRoRyD1CmzSkGkMvpqVtTkDphUHZthH
DFFwYk+u9Ar1v5oXasvQLUNOlj155PYgt2+UKRH4t9pUvLuaYUgwMbtCt2hcSKOP
mEXY9geLqR6BdI3y7q4jlVzFyoznJDLdIdmzUr8I8g9NdPwTrTNwhTyVVPscSqr1
mNW77MvQsXj3SO6NYFMHgpUkWJaj28FpaA0bVyxPuQwSBHuPRhTtrb9YeUgTFCss
kLDQYCjMkuIoDoQNnAxShWR7KZ9xvI5vSfZC9jOdhyQWJp8JAzHEufmtS5Dq/hgx
P1FtsECB0A/tbytZh1q91Y/aT1y5QRpMkHJNbpoROQp45uy0fLSDXLAJLDowG7qz
O51h8tIIpo4MX/iU/1tVFseJhdOEaFJayMpxAsO3YBM+hj7Dq1elbL5TMZvkT7U8
lwaVupfKzhUbqs8ZCr3u808nDov9gFPu+tgQQIBwgCoyS5M0P5WzCHiuV87bDsU+
eCUSiJj6hMZQiM1+DQbk3UUkkBVNRjUng7ROhc43M4n/MXbPBHjun3ePxrgOGSXq
tpX8CRF4j2kuhG+9qbixRXScz5N/dEJl1KzrtTjWU+zoBACWBjbsBLXrGPVi1pqE
iGpymeGNhiLx6n/GTulgDfBwRibnrTNRmRAbvQbG4zAMX783BcYb5JfGSL8T4DAQ
NyUWx1PSyRN8Ir3aUYbUW4tdB9m5CTfA/IQHf98hvYGOoP0CrW4QePsO8z7Jrtdb
rFRvMIIm3cMzD7E2RmGCQcXaRSLyDznT/58FKF8uVdLHE5pZvv1F48HyjEBJAYBI
1U+rmmj00Ka48rgdvqIciWbryxmfjL4/c6Fyzc6zVknm7KAr+4C4rF4jQs4zyp7T
3O5GH/ULB/hJoCrq9zGUcT4mWHhnInY6zrJpsf1yt/+Gyb7JW+qaQ8xpIFo9Ouqn
6ZJgnBRZONf1J4w7rlmJg25aKZjM/ElKGOdMvX96ifIIEVh+UgRC7Fr4odEWBiBr
ASbJlDdOCeSKIUsA4ZmA5OJPumLHkRJLtVVQiQ+qOqbeu00Ov2kG5onVMvoLZ9im
SUrm+PAAkuvEFt59eoO2RnRrgJdvpvEh8DML1m/CvlrhoTujAEfQZClUlEbyjf6f
qPnTvyo2gE7I1r+ihyOCE5+jHQ2AnhglivSKLbLc8jc1/8ulLoBep6Svow7Na1+o
us/U2+PZQX4r43Es9eyP9MD+tbFq/fa+ZdPDNe9BNpKhtUgHv4Y+f2ZrDe0YKeNu
H+4QbpdEMRSw229G1lbU/K9xtg0D8xvdZVDwnNqfAG0OOJu3kShOthkwV4u2zanY
a4Sl33RV1A01cGofwa3rekm5tpN5ZF1+9Psjn+DP2W4Dy7PtCLFAr0A712B09SQP
GKCeEMilIYlcmKNQ7+5tEMPgZO7EclguCaOFxQu7vs2rUWTJdzOiw904Wf1xCcAC
2QZwoHoK95nYwPhrjpnDPRO55JNj5sN2v7pF/S5d0lxYVb4dZyXwCMAt9vOz/HmO
tiL8+T9jEeLSWaBBO5P3iehsmMkdnEUCH6fYJ9kjwJMBvfOGbENCoY+SE57sEQ12
W+PMxgF5OdYP8mYWJjGvOgkI471573XWqujukn4W9I77Evx3VqBqepHDBqz4rGk3
8GAEV7ARIj/V7XiUVdUcl6eQ9wKJ9GDn29qPgm1fKSXdh/zlm9B/g4+bi+TnrPNV
KnTB5NgR1KkM9sDoRaoP8hdS9kkdD5YJfZ3HMah6AIH8oG/ZiKiaimnh5wTmwvlH
Lkj/rEKaI9SvGlzaLkdhN1f2zwGH7F02KsQLJZ07OUjkCwtoUhmPiU4Zu0bGiBOX
BF8IAwFRNAQu7lo7pWdNcNWdmymR1TUsWatt6uqHQocB63UjWYI/t6luWC/zSX7a
GqCpQxiAAmAD9LqFtZ4CfW8XWVHl1yhdPLfW3ItYwWAkS6RwLn8Gxt9v0BYaiCgd
H/DUWpexi7BbV0wrEQvoANIxowzO/2pKTo8j1vdAfAWB7hi4igfmGrur+uLBbaYt
N+WpxbeOEL6IO82Vu8zqD6lmYsztGg6YlEfXPGjCbJNrNgj51GaRMiU0LkCYIaeu
JOYsa4ecfkzbPRSC14ffpAePMcK1K5vndFt6oW8PRee2PMpIbpTxaP7Jbg3Y3bQo
pwRzLK08UNl/+s6uO8dKL7IMVes72/Qor+qYFIaafm/EiwQmzRpBJHQQtS0ar2yf
wZ6h1edkks3b1Q7TmKR6tnXgQMmwxqHGflkJAZhr7XfWwHTNEbATcgU/mmGMy6Ic
baHpmOzATFzpNXgD22y7dyAXj1TNiD51M+z/CdE65oGAYWt4DN3tzUv/+PEzdwxN
bEAessRr5qA6WddbVaFRIYHmBM3i7kSc5w8ewp7sqmX1UeZAWEkNalZ1DC/5fBZ/
2jeJTcoSAFVWKCmxrJwlEOBnaWmf9mgP/wu2M9rWjqBXP8BtecROKCZUX0TXreAd
`pragma protect end_protected
