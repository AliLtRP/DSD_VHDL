// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Eu93kzgsKeat1Uc9O2Kd7JQMF+KhBL3zLd+/APPajSrjCqiWU4vX1lcuh+72y3db
G8Nrja4/rE6uBieFwBy0Pflqg6YvnSDINq8c6zWKhHoenjQ+c5Df2vBQnbCxXmsb
f5LpqHaJbIBNMQG6xY8J3wFOTfw8CvttEyFXwUsuSu0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29056)
30g+rFS2zUY5EVohcSvA73+awHrDsardm1qZcE5zBBO7166L3xbemRyA016QFifx
dwIkSv21uO/XWH6EeCYHa8E01qQN+SvSdg1hbQVWauiqZsvyZk6D9ff6/3hohw1k
npiY9Jfd6IHfYIU7I4/jtX386V1nexdKflaKrFMPnFHj2+XoPqASzuyfQfUJdctO
WgALJmozOeoOKckLbaVpVHhbISqz1rGt5TCHcSWN7N0VS0TUJOhDLt5vlmEZTSME
dzxUWFEXIqu6v/zHBIpanLFpderFnPNnp3gRupySFuoHMOKfSknJkAhx3S2xrZLQ
MUOAxrq69ZiH6Z0N7cGRCKUE3ituJyAGQU+BLcwct3z7Ck/5T3uRmNEYkrvbSfJA
be2hgEeP678xboJLDmpypTiv6ClLj2nWBy1ddxJpEZ4gNBfmDBGfpAZc+tAd1XVO
O/2g1r5B/b2a94XnIr6ncO/q2CYDnV9T/g2IKMPnXNdWBfI7Wpm6HwTr2qQ6yiC+
oQduTki/k7DH3J83E7qbCcEOhmcisFQXz7arEphhtYxGlC6210KTzo6f7/uhkDMW
eeAwJTpYe0d9HZ8cILNwtsbct/De52sbCKYyQaiSJxDaRU2ySGeolQCJx5jwhr11
0+lMQ6db2c2O9y3QOlSNCZvSidZPhPUcqFpUr3aQFD69xgBHkiUBVNd5gJZaLf6C
B+yekhN9LvLI/fTIIbffFgGvMHG4993IQE1GbNL/VBqurhrHuICIgBajBOcA5XX7
b4IHxPLXni/Tv9uSn8uIxXKPAPXI70TIL0H+KUvCbjJv8vaIoRbANaWcpOvbwrX1
MVDUThiTprthnVvwm80L1SS6CrE6CYMR/itV9lZKNjot95InlTJbPQzLA8lRGf9X
JuwU+wQ8A9WpJicSNdJCZPKSZFebjN1zYV7oAMhFmhzNEGohZ86IzFtNImReiVDk
X+yDyyhy/JXJr6vCaYsmkY/4pacf3j9GbXm6T1Cnr7qAs4RsaeJFMMNz/K84cqdd
EC/sZtx5DKF3WS0jcgDc2b0SR8JqgDuufnOWAb1TnYYKdHyzJM9Fz3tCaobL2edO
t0HOQR2uRQO7ebR4wvrKgscf1Apy6eudnDK+IdYj0cBxS5QhTV/PpEkXknxlom2E
v2T6U9qlLfDAg2F89PWgggplkWsVHaB2K+tu3X0VVR/oFLbHykcVpLt5lM2vlH+U
6B2VvSeODj6K4LZNeZMVMN8l1uXLJ3OwtiLb8oBPMJ97UxMgr8OId0iMgos3bspn
SNoO8hi37WWyCgchpGolRm9mXe8IYdomJ0pQw/NrxAaQwHwO/Sw/CUEbgMs5quW1
p87ppsbO3U6LdWcBVsLqd4+7OUwQQ6D2BMOO+AnCdR2y84NndFonUG8RMvd8O7f+
U39758V91icIyegEjmeyhqlSKQ5I4NsGa/YRwDhp0zfsnJ+UGaeem+a8Okw45MN3
Dhscq+uk11MSC/FYjKz6KITbXoPzn/3u/WJMyoHw9dEomiJho3nt2AhOVuZTP/hc
SotCV2EIYxXa9oyZnF7OJ5z7B4VDBVHbE0aoaE3wyrhXs0dzodGp96BYw1c6G5QM
+mZMDli7VPx8bKNeXqv409QBJ9zAEeOc7sK8pcNQ/DGA0meQziESp0RSOy0URtTU
TxE8XZ9qoRFjlMmF8MJO8s87PI8c9SkXThDDHNqYLP08YxnUTMqAc3Lu9wOjpM0A
qDqaBJwQ2Uxhm5Xn0GjHkmHfUV6H/1l7PZZ6jLMXRnGY7JmuyfZins9v+UBzn0P2
WbxBNLGUt/xhZJZ79kMvk1UyzYajvbQgAeYP+ATQ2ad4oik2GlldWgi/Z64o2KYv
uI8ptMIdqqEaHJavHFe0viDwDNCWkP68RR5rOUNTxUiP7JZs+a+CUf2tzeWcdm3P
d6PQ2lWsVXn7d0gU+abycigwY6F34ZY6gw2ZjeJ9Jn6i+eL5DlFAkma7BvsnFzEB
bV8RMJSJPoqIeCAO+UT7XMEZmicFM6U+B1/8VvG4tXd5rfLtF0zMInVQ2esUk5GC
HVzgmKKvkUrcdGcyPbgKFq9LblKHAPowj93ljW6VdDMCCCVitvvwV5W3Pdlvl1qu
zQsfO9wvvjEVHnnj1764w07/wXUffCOocU3lVS68tfVJEUbxV6AjSsQdMuXTMcVl
WXMKsNRDBfmZmra/M0FLi4ygyHk38b4dxR6BlAn7FNfe7zT0aQgeFTWA2m0a2qN5
CUDH8866+o4ZZpOFjMZczNvv7dagM1GyV6J0WraOmeoxNxm/sbx5hwqTYsrQOf0N
tYEJAnvxgPcFBQt3F23PH8r0Gwd7SWFE6nw6E0U3K4x63jiAZ+5OKwa35g9rlBPC
SnQGqALc7EduVgAZ6x1ds/Q5d39d7XSR1wb2udPnLKOE42uEonso4Iew2Nto23ly
wM0DLg2apXFsSRF3b/DmYKLHmUVcJQvGjP7XmhElgFWGwD01UGsypdKlhy1lNsR0
JhBvVGtZT9HDNXtGg2UOE/M4j3oxh5pSR2Dx8NXRVGNeM1QP6d3zhGSrAIXwTbYU
Id6p0e1yDN+/nZBMW8MLUHfYpOofh8dHQhkGDfGzLpXyvXjhTI5qjedls7INDZkL
Id8QYtyX2kytIVVgNC3K0Z79j9iVD62URxKPixA6sfPp/rUb/ZXktkIyANnme0bR
Ou0bjXrwsN/i2fFYHDGE2k1QbQzSOew99Wfj4JVqr/oYPo/uyF8jpbbk7cQfxBjo
ohiA7MWIQy8z4WM/mVoiM4dGsRUp9DVgf/hjNyxletF6XKqwGIT4rocNleEtXh43
abwOrTxNBxB1RzJMlIIF1kAmHQ9oXe7SAoLPQDjuNUfA7yaV46oyrEf8ahfswRlH
iqgIv8I7YhWWuxXf7U2sB89L5W2YpHpRBZhmzsEErFfEXTjZXuZLoN6C23zRDNai
Jl1rP3xhLpt0lgMfHp7YK4Z6OHdC45VEd1XsdMfYjR9PPNH2IlLtpv83kkJOj9Pu
YHgl6zoFl8Z4OC0SvcwKWqSLk2icnvz+qHgyxXJnwXa/oouvkxuc8bpV8lvfzYgx
bCGkldP9piNyg7kEjxHQWOhsaxRQLDeCfT7LZXRb1F9geOvKy9LiYKBPJ4eWQnLF
S4rDEPe1qnj1DR2vt1Oue5ABYSYTrDRYLkorYRxF0A6spi8sojMUnOs4x3DyDg7m
hxtGmAFlkbD6rrIVIeU7O1z+nuFhQo6TkTaBmm7GAuHW+S0KAQnKmVlt26TkydUr
Njj3U1vYih/9L+Tnta6NfHCiPeuJbRD9mIiFULofC3wUStHBsn9WY6rh5R2q/xni
Grfls5ZuF/1RclTE74FSgTdsG+gz5iMO7rrJrXKCyg+2dceGLxn6Ay9tbzpVilvx
L7GlVA5VHJxhOz3HiQASBB7p0IpoAGAAYCtA1E6u6fGzQLwQKpMOz9KG5tLfoC0N
48dU653JkjEl82l+i9g8cZKe4dq+8WbvwvUXrC6u3zZQPKA1BnVkwLKCYWSAv4Ms
+Mhtts9dS/gtUp8DNAv+QCxVME9uCQSTDLYhUwlHzbJhn2HqRzi4OSj00y0AYLPi
pLhhwzv9ue25xZxvbTEPmkIaxTYMkd+EGGbT1G4WmmJWduYlsCSGvWufyvjuj0zM
RC8CPxXsF2pveHRTuHnY6yRSHDfg6xmgeCsbmqcXhA6xDiNlhBx5dvKOS48/MomY
D220GHfgTmDjbVTdxrEVnPJ1eifJaLMKTvvHQKrcW7NX/KKW1Cb8o3zNnNldqJZx
XgPh7oe6uilvoLYJGPSExRFRHsNHwFibJQ3StjxWUtB5bO0+6h5vShBlzxlp+AQl
7j5cnwdzTOuqJOW7qSzTZylUN/fVyfma+Db0EUAyL6Yo0Gymo4dnMPODjXdLJBzo
8INZdia97tMeJgxZuS7mWu7aLMrU5GrHG8KZJYO0/PGkBfo/c8iZw2fYt2A2ENG2
9fd6ZLEuM8CWLYWI53kXsY6EWmWKOol2glcl0EdcvIW8s/N0aTLE05zlZRC5mVlJ
aTa3cpw4whsDNTOImlWJrOgVkKV2Rmq9OURm/ZCaiF7X2b2Dm2yhKP+fIxYREbzC
6tGxS5omHZjoNKmhjwb2n5ynIopHa0vnk27ByXxGStP/cldGKg1aq6JPL+auCnbz
MGU9fZrkynUdnXOos9Tq9WW8ChJQKNZY78Q3HEQgGTinwDI2jSVbiGya6i9vPMgo
O2IJzmzuiC/5jimghc2uXEM6oW7TS3ZGB0brwJcD+PldxhW5r2YI3qVy4OPLtmne
KY8Ba5i2MUsevWEjeVYaOeJGuhZlIUkh1a1RDM3jbj19oMf3LZyjiUNAJtlfDYUW
xf1wXdGeIezoAjF5uJYk7uw0GllN5O7f/53jHN6g8etG5nlTOrZFJ6HSE9OAF1QF
u1XmG+ycgyWHrYxuOoKpzoSset8irOkgzI3rjyynCtFQ3ArFJdXxoEsPXK5IIW4R
0HejgSFvqYxx02H2wdqiyco8G/WgbeVATFFf8c5nN5LOOOKieLnAN2RPCNaeoMvI
3oigncWaAYXas/1UdA5YGUtQE8lro9DOlOjJydR5/WPmg5UxksDvqMMLBdioTOSN
LTf5VvkViwqJxpJOYlNmcjxb61Pf4ZGcjtGbFhaXXKZqmbkJkMzf61S+gw7I56Jk
WlXsYJA5mUozLMXGda7jG7YUIvXYy8ttOsCholPVKOmbbZf0LlIdmZGOKqc33zqS
jE9OW7Htw5GQJN0CS/+tK6w40RBUJPBzWxlfah7blw53jHxUlAvdUnVB9OWyzYx8
LWVMW3g9TJnOlu6vHU3u1kglJbM3tN3DTXsJiQjyENbXa3aqXe99ZMQhmaLvd38f
h2hSv0U9UXnJ2kEG7gFfMo+VIffoZRtBgbRWfnUq40tYZXd/mrtCOTb66CkZEQq1
ip+g3t4VkcVmrQlYyllBt4o2i63b8paNMGRqviFNcCTBfZkvHFISxr6olLK7McnF
a0XRiVGPRpqa1Z8F0VVPV8GJZcwsRtwiGzi5pQnUendrpzRsYgTBhsUeR8ocVZqy
GYsnxsbxA9eMZKrx0/FI599IYK1rGsww8dgXDUvmnH8sXNc2mMNKqMo7Cg3s4ZUH
oVCfIi1dD6MgLH1H4b9q882kMKR1p5XVUORbxNnK8SrPA5m8HUROkTMFJVGoUMMF
GiergtEQ+NclpD+IrCg558g+ROAwVPX6JFLphUtS886bravKFrmquHJDGcnPCLaL
u3jimz+X8gWfJkHK05VicgLcKUcXfJoQBoH3zriWV3gICG+cM1txcybb0NAYR6fi
EWokjZxiB93Fh3X47JS43Rv1/Mr0fEpkCBTBRiCjswmE1/gA2eoxNKsOObZKwGdO
d6/ZxMPSFUQ6AQE0HIs/iKIn1q+2MHog3DCpQSurYktCSiSVWp1QA0mXKOn39m+l
Z9kuajhwseG4RXnO4Vfm/1WEmDHWbUQb7YuWqhWzCIrALPNUi7Z8/w4wfGsou6YM
JXP7TnN2FaqU7UwXkuxpgNAFyrVH5fj4PdZkz5mJvf2wkv5AGuRmGq8lVqsVHUR2
7XnpLqL8pwhT6ZBB3Um7pM9M5zBHw8Q50mjSXNc9XJ4L8m3CUOiMTtBkJs4Lk9Yx
jBeru4zNRGpfxgDW0rxqJiBnDUgdjkMqDSKBFbmn59bYiST3eIKTwEfeJ2Rb9vBo
GoLDYRC755PdB2+q75Aj09iOYdXB7cEKleY8CFEvlEu5+FwFC65pk/ywuC7ssAEi
awsaq9k7FDX2mN1MuYtrRNowlK3L6QTJ7ZXZiHraQuUyHIgL9oTGgVEFKzFd+QxP
lWN0L4buX3Z5zP/f2+SPgADUyfmFOYPUNA8uWEWU2moOu5H1z6EXvo8ITfM8KzP3
IcAKmDLTNrZmpVxTnIoEu7jQAkDsqdK+fxUftyouMhjuH8fRdEquRPivFlotIZUk
n9N6nLQ6+tjp0MjkTAqBraZ1exzrULW/8Scg1yof0BUTb3qfdtIm4Vk18+g/nyHt
AQZ/9fA8JwjCHLJhEst7gC/nNTk574Xj+7Js7sUTYZJWzzzhtfdylFQNhkg8/Upm
pdptaVb3r3paBsK+SYiCjD3oCZxgyl//DxwZsNqoSq74bLrjWppkAVfpU4GNvbM7
4E6Bjbl2hXo5zTeW4RV0nycqa+XDdGctmhwBrxHlIxsxRlSgvmFNlEEA3InBtkyo
mGJv2Q8igf8MgvFFMCi6C7IzKZaeqHhQseBmQlUId71/fSu5W1Ko5zXc8TPTIqgC
QwlBtY5H9UsgZ2jiW/Mbp0uDMs6r8xvOn+Gp4qA5776pyoUWnTB/HWeh2LsuPi3L
wgDAuuwzPGXNKVZzCgzLFqxowGBLZSEUv9EHk90iHanRySOVEwOuKwuYVTxB/rJA
hqOuSpwt7FEiCfQrNSPX6B4rhwM5quNqk//YCsAsTB9+X3QOHuuabL02/A6RwOuu
O2j1LUgWq8aJdA9Yv2uSo4SAm3Y4i8Tg4jcP7XMBCKPA/Iu0hlrg044y2aQ6RQiF
lu/mrXL+tO+HiWasSq/es/x33Ug0/dK78nk0R14xWMEUahtGRVQm+7imvz7DFLck
dr2OjL9TzCuHXO3T+qw+Mp6DOdogFRLpInYHLDwEAUT1L44RjESOGcTuyymK96un
/k6mY7AmY/eaFqTEMS/2N57wmdxD5mZpZT8IeS51GXfw8Zd2yZzBr3IVuX/w0y1P
fCftKEfCxRdvEmrp5obl7/nlQnKKjKHe8fxoVKcVzk84O4Z+gNdAhIUusRC+MNQy
yMPgE0nxuVDvWI1B34dX4nFKpKelJPknXHR0JwCj5jDYIvgKLXVZVO/MuXllMP5k
bRAIETjk4bosmYM90LTBmzGPvZGEE1oVRY4Qtlbye4q/Rwh9giMJt7MtYMyP19Kp
OKhT0RkgrMU4Xl93ObhOvQiaV9MidhhnSxqHMCe5dukO8AUwSBfF/vw053/DqAsf
b8CjRQldx/Oxikqlwcbm0uJ/jeXoRuJa7yZcpdiFfqJAw7tjrilKkpnuR1bYECdQ
dkMrFNYK2hxknwSwr7BkuWWuiRJt4Ii0lvmTL5RZFfiypF0nju9IFFmdlsS1l2H7
/KM2E2r29Y5K06/TS0OkGVtyGkScrELP/JeA+sOx19VrX4IUbbq2WHcnCTfzL1+B
ilIz53P0EK6NHvEVrBsAaH5qLUdSoXrFeQLqI/17OHJz2s1qohZYtIygXzXb/QVU
LUSgUsAzuR1e2Ky4VKSbENGb8N3Pu2bwd2chl1dUzFZKvBJoX7HzyUBE2T3nufMu
lyE4eRKChUFfvHz/kxTU/2nc67N4rpuoZF/D7AoinSG3a6P3yOW3zw+TWBN6Dwht
+EIFE0wZcx2eiYzJlom2hw2NqRE92/NNRXzNK0+tWP6k0fssc3bVs/1V+zh4CRwn
OI70pZjiH4p/fC4934MTMKg2o63XDlyuGfWPx2lHysb4aD3HwvzHX/wlcHBUB1JE
rrSIZOIGxorRicqVrK+pJcKMpc+c9H+VRgLwpgUeApEYPVDJVDo4BOxlbihN3OBy
zgYvVFI+e02SWraD03+R19ZFTsxXkcuN53yDhQtMiZZpfNNpJSnRQvsvRc3GMNxo
oCgYuJsnFnokFtDSaEm8PEtsCzuEqM3RzjJge9Xn2jY+NXwvQGhqJ/l27w7g9mSl
hh7+Ai+vBEKV1q49hWzHcsynwfw2z/4tj40qZytigVU9Jc25pVjZ04y2sTSx36JJ
Y8j55NSFLudX7iQctDXsKHPvgByEQRq4fDh59XiHAVXmrq9ujycR8qn7MLnysnlV
NplDbqdziJQRXS3pZwC5ulcSvq+ilx+iv4xhbSLRk+Um9kjcV+QC1UTUOWWfHZlJ
/mOx1UfaOEhq2szogns0Rq5y7+GVv02PbhFnaGwkuUIJnszJbiKqIIj+jxabm8QL
hrH2IEvy1EWPahOQrakvLuTIC0EOJYD72BUmjj3HKG1ziZgTvszX88ue+6R6f/VN
ApGtOkSrOPbv2Hzkt+q1wfvGEU/Glo73GvnKrsVd526h5W78BtPXriuJUz0Owjln
50/Qh/DtbOWgXR3WXcyTVEyoynejjkRMBvy4ErOvlQGUQZ1nSffEqbE+wCTY4vOb
xnGaa1BIp7pH6EUtbMxtj+pcY3l5qpeLpFwaXIb1S9qzbHAR0nLNiuqnfvq/acLF
pfZiIcdTPf96QV6j9V2JS2NDMEAFEgVob1q9Gx7hV2qX+CJhtgkoyReVRIG0DycQ
N90w0AVhabqIf1BB4M9fLENPHinb38EUP5RDSa2w2Vwm9H20LCqhWh0EqYu7FhjE
Z320gs45x7i60cVs7THq6tZCzXnZi25c7pGiJbUwUE0cwt21SVO5RAidtPsmTB2z
B3tzWlrc9KCHYzLJFBZUhFC28tyiE9xOO1DlJENLFb2KhLLQrXAYCaUCTEhgg9oL
lB7k+n+obzClfiBa6hg9YPnmpkQk+niLxNBClZNd7GOx4WOJaluLca/DaNhH668X
UuQ4tpoD+4RF3xjaOreB4nF1ceySCGRxP4dIQKEk3owQzNurswsPhQtUchcd4yAn
RD9yGz+b2TJ3QlyKGAX3NMTjUPMj4YGQ5vVfNYuV91+8d4Vpd12diA4Ngl9qJdMH
4CgnjD/wq5q5ii1/NPgPdYEYHgKd3oDRDqpsm0hAWfH1zltY1kDwfVTs96298pp/
I0/qNPwc4RIlwwM+29wQh0Rt6pa0brTqlMlUEq4cCQR3l0vFb/mEE3nPPXB49ADM
JptyyienMK7FDrhXu2O2hgo4rG/5tvEZ/Osb1+974cltK7U/niwvFzMiXsv5IpDT
vvW4WG1eIOAkuQAYeT8PYqzw6SpVErpb7ExILHKskmRLaoaQjXPDBYeGXhgdytKw
J4HZ+CmP46rLUES+frVMxRNmJBLTgLOlWwPuEsIJd6d7aye/BdSp+yCoQepIG2Js
od8ar2bL/n3Ig3kw5njUYsP78WhYZyQ68tlSSafIKukwGTO4po8cIEvbOaTA2xlH
pTc1jZypfTavtQ+JlxnIlZ90RcNZz2reuJrkPlAWcsAHQt7XkflDb7sEqBf9N7De
8kT7Su749JmFC+grEb+0MEq2UyyWh7Eef1GEJpKXKRdztqZf5/XSsJMFPfh07eSz
f0LugqKuh15PlL+cSdyZHTq2v6uc4TMyQ4SdwzRCESf4x0ldlj5FZfE3XjcLtiIi
D56s3N+Z38x3Y9QmBu9eRAz38p4u0acs5tXw6a3S3JxrdZZD2aY2WN/OPPR7H872
gd+nUqamvpejjAMpWfpgG9raN1eyLYIn4Bnjos6P9IYW1H8wHy/D6VmvI5Ahfy22
iZCRlUiwaAje5MIdU5WN2SaScRvzUJagR2s40yLKYOv+TyOYxdFpcHXAhgF2YVby
GrN6TzF7O/RX9mIkaZc2BZ1nBK3GvnvXiksYuzuki4ZXEuYBkXMgUrvz2/sBnw49
L2tyBkJIru4NBR5sXqN6Qpc1t43Dl/ZfLuMICPCBkX0Vkf7xVXv1ylnxAQfiVkCH
V3HQgI423a+4LkpMBH5nmh92dPYoOQoLifcObCNVmtco2aOyQWSJDic2k3Cli/5h
8bT9fEpzPkS6KbGvP9P/zAXmMenIR/vcNsgrNtlPX7+xW/YNG8sMXTKkP8s5F1+v
5gpKNI7zkKRuWNBoymYtTEXzM3hs7MtSkeqqiF91lolJaiKBkp41RYHG8Qiat9Pu
GXi54H+1SE0QQJjxD4iBGQiSve5sA68traVG1GWFQd3Fy+xO3VXedqgNfjgI2JP8
y6S1ziX0UJWR5x3596QgKlgrYQOn5/obgNsAH8d2dDEpFD+t24s2Xb9kdHjY1fC3
DGISQ/GR+Ybo5Q7RZJbnF9bsegDXdlo3PVuIwFyd9A4TC2C6CSwmzkzmh2gjAs9v
U4qAXktSWUJBpZwpVDD0t3g0cm5rhz4gIGjdft27ecBaOZW6IpPKqkKw4eAnNYlZ
BYhzmEVna0WpNBjjhEY5/3KfO42ajY1XLjU/lVSXvqP0AARllY7Ua3D1Mbtp9OR5
6bgiQwzufjFX08Dgbahs6utn/ZGNlmJQPS3Ce8rCiHFIp82ibt0+6O4KHcgWxm3c
3k+4twHoCppAzi0lmkGvTVdtFUHxgZLocknoVq4K/dTrDHWBY4xURiFOg+CnGEyD
yHwpmu/F5VjJRk4JrBxgj/wKnwi2gjiZ6cTafELMLXvq72E44dWq8Ll/svyW61dQ
9ZBuC56q+qnMB4FzJcSY8FIdIda4CVwSmx7kRPzz5W3YVaxxljjCtVjx9LlStyb6
6SZshw3xdbQg6RQq6iCjeVm6+hJpmfi9TW36S8UAZhNFDUZD5JO+wvt9M1qcgNzm
fpXzmJ2Qsi70cECGK7B7y0Wcuj+cf8ChhfcddMbjDCjZh/etudPi0a1arOYUXfAF
k3UqVosui7xsFY7wmAoA0S7zEmrwzwm39Ai5jiGGoKfhR77uy/erxkaCJ1SISTAM
loxalkCQTTEPMRkiM/JmFCqaFOihjxqu+1frTkzms47vnAGFRH5LbqkIHsvO947p
GLfvov9031olrO9cCTJjMzDXUY71k/Fsdd7m9uiPZZQFInx5K+fHOPHXD+G5Q4t9
OopeZ0jM+Pz531J+OB2XNUs6607HrhylmfYz0+MILz/jSOR1mFdP96qrnxxvamlA
2mIam+LEOht0V+4hnfPcfWhPJki8ChsF1ts+/oNj5t1u0k7V1xn1mLdLRo6/wPTV
PZ5H+F4WPptLG9ht80Pr/WoxP+iV5bYBFzZJ5s6HghkZ/AVPvebVNmQ+yK3RSEHM
FL37dqR24kvTck2FTdVforUzecbwYSJ8n1mumoeK012obR3/ikMetvuqAgab9aVB
rrsFp0XvupLlSPSNzurREy/0tpaHousYPddfJwlZSF+dSczIaZk29c7uRfVBCuxW
s7/Vf5lTjuuayiiKgkvplo4n7OEMS5GgXHZItIuX/EM3AbECrKR7NzG61QVDXneO
eNEeWRAeiprdgD79SBN06Ogs2LGciqUMRHOrrXi0JOFraAZ83B1fHlR/LG1T5QuL
0TvdXE0qsE+9sZ+r61C1lDb58++bxZ+fLBjTGObB9FcOI4Uu+8QZY3fB3D9wa6VW
9V4FZDmMaNH9u8u0XAMsgUN67xN8DsTD0sX6o6oS7ry3M3AWfWFFP0CqrgQ3ZFS0
RfvDTDuylAguHjZpKKiMVbrlQMZIp234lQfZGIzaxNXHZo01htUZJy3apE+5cOXO
s//8FZ7d5WSETwBd5sFD32462zNbtCbK4jCMuGs/UPGKr3WMcDHq8HZrdIjpzT/2
rC6obdC8EGfa6xE/re9UNN9BHlWF6Jc40Q7YuiMu7utGnY9Ml6CIJIy9ocxWO/0n
kKVNeNd2TLXwHpkdvkIXfX8erDQsJeMWujJxy+/cUTTyuRDdKcv8DiLzCTGLtjlL
M3AlTRUvnMVH/8ylQzt/vc09NhgrfPALeQGW1XMomEiL7J7odZEBzfGSL0mb4WpQ
x0K/SQMdb1EJ7BS26oYBcfs8cPIoaozoORh43aGer3WQNFLRN5LHsc/Vh+9QKGKG
USp9ZMtRjyU3My9h/ekD+g7K1Sf6+gQhJ92SB2grPEF5D7YQugQqr/txAO/ujUnX
Ko3oVuIV57WOeNDLviCUxkA5gWFd+wrQ7PhzMvn1sYIcjT/F5UhktvfzdmakIH0A
Rl829EE8uedNjaCi2OTOYJFc+kHZ94C0HD/RbnMaq4iVpcB7afXDgTUpnTR2jTPm
/CHzSaykjzMRbJ3PDkPIMcMl5V1LRYx+vY9QS+x3I/0JYFjPO28alV6xq6UpmtSt
SNhM95moeOLKvGzD6N9dPtLhf3xb+e/bLD1BrKpwP3przPKf0AXdIZO4/P0rrRHP
+2i9XGNoI9y/B4B9mGQ9ASGm6pVuZEzyas5Y7gmi9lG+mFNMoOEwtiBOt6DBRcve
aGhXxX07FU/Zbn7jtN42yemkFk8ksz6fLZx2pYvdqVWL7aCZEKeFC4IOVOAoPAsc
rAwGNj14hO4huYvDMFXNvQGhGX++Ad/QQrLF585N04OH8mi9cNOdx/JXCIaXgJTF
p3MuEAvCTnu2asl9YSigfMpLVbUzZy1VFRKMn7bvhXK1Cgoj8ue/qo7c23j5l3Cf
QiG0p+10YGR0I718nh1ROs+gMds8baBaQxcxgq3LdYGc+INHrFtSKqijQWZWW0ug
b95mzQpFEnZq2FZwmpPblgRCaR+tnWEEybchgEW2sK8bBqcwLCxQaSqbNyIEH1iT
Fi3xbsUua4BgWzgKsb0I1XKWaJp9fY8duC2L1graIzDuEMbZ4y786Z5/Z5ZGt4MW
LTgtudok/xdwPz8X3NbKRC1ba8H1JycYZuTZpf8okeyz13lmpf+FtcStX+PPZTYp
NulY5x8G4pkj6EcbzGXl6RjLvVAWho6C+gQkYBScpHHabcSw2chyIrq9Zr8UPTBA
wJvdOX5D7gHu5p8bgArS+3zhTIoaNFa8uEWFF6t+K4tpB9h8u0EaFNZXDqgO+7I4
Vx//a3osRS1pyIm3QJnvdS5KfVBbKgg4viAUwO+xNJDC7CO2ZVOkZ7nvZOmbKfoT
4mXPF3H7sse4uULzpNgmnEbbQfxxKpbfoIw3LvobRvhy5QV4QhFn+Lk5S94whOUH
UsJ+j9mqn6TUUHxRL9/OPFFYRY0+m7IbcU7aG6JZgT6dJZrMADsrs4MyfuLuJtVS
3HqcMhPuZdAHSa6kh/2E/gjkczXEG02RUCu9P3Tx3MZQPB/qoZlRClZOO2Ikoxva
k5bwTWAi++sz7YURp1qF3YKhrgBJY+ehf4tAIKj4b3Oa6OTVdtksEkXanwaVTBrI
FwyKWuNonhu8WEcmR1csAcKV/oI7yJoFyh+7wCQn3CXTmUhLTU88bGlB6QMDV8zZ
NtJD3WlGYHRhCQ4s5mLSgxJBwpnUNrRoolX9JSr5fA2sVDSFFqICwAiCk3s1qYlC
Ig4xZFF4XO4st1pcv2JAO+03fJl3+jvANavSp9b0+OXRhgXB3NCgLnd5ByxOXOm0
KLeE5acSrX8H/mkVasMxmvNHZsHcrIFDRk312512tg3uRjc17DoLQQ+poc2uvIY1
OcP/4TK7agsN0RLlAZ9bQLyDiqp2sKVqSPhb2rT0FDEfwSyq5tfXGNSVCSHCW5zl
NIx1++PTPEinrNKPxOWJas1NbhdBVji/uQ8ViYZexmrCDoZDtYBI6RbQtra4pImD
R9xC645VSY1Sqf+f4E4Iyq9hqjIc5i8fWanL0/ZLF6XHnpVXhIGGVG7VNyaaJxbu
r+sYZipc4jhCYUv7Gxil83U9pPIeuN8zVa9QRwq4w/Ebj82WtdlBfuDsuPCQEn2B
ha8xL4dXzNTzHYwUcxR3somCzjF9LuQxUOkRXsDHbu5tnTfrq6AqY1dzdKaJK923
FhIiOe2nRa6Zddq4Ghm3L759W7rHllFklNck2prQIH3spBccK1KOxlGLwa1/9H1X
Pb2stJeM32oHpwtwsr7os1nHxOwme+uHRzC3xMnRzeTFiEZxevSYXZFFORtYFmf+
i3vNfQnHNRS25lcFFfYigJw0Y2qpQnFyqXfTSic4El8TpClGSPY+Wx3T2U5bAWE2
kAsQEwseSsc4FWAGwuiInYFyb3t1PzMx1NCxXtUjl6kqyK0whYbQcW/ir+jzQDNG
6TJYaHoB9qBehU/V1g3LPw6jbD0lUC2vrzYlx89ZXrmrYBUqTrooqvDUyTRJDJtS
D2Y5YOtPdv4PSzFd+eXGGWb5Lvy9W6kpxZL/aaOjjeQCUp7yeIs3ChlqP/LMe0we
ngUgNycQjrpCpHo1acWyhbCu9alFq8In776K7DoAPoXXAilQVPl83ZBNq0MgiftN
UHKhyvt1cYO3Cfub7NI6zp9aVBMywjGkJNagCj7GmjuG/E51r/tY8R0q23qSkQxh
xmH1GUGvaKyNLIDDvrijpTOJWaQEp2MdkqwI+L9NzrKzGutohqXUh5uMvlUhJdNQ
eQd09nSVxw/SRes68qnEAZbf1QIFCV+fTm9GOJvMroTF1mddQvJU2p/nOgdk/0v9
Y05o8r/HU7GTVeNaQ4w0FyZPIuQb26hqVX0YYp4i1SmhQeimYxfNq8Am7YlypCzO
jWPWbq1f3t+brw02rqAVZA+B2p3lk1fzsSY9+4OaGzFP+Y8gfn8Kigsanc3v8WCa
7FIhvgpI+5dg4k9JtEHHn7YtUsH4LrE7/K7K1GEaQwV2b2VkBGSLobdrOY9ibZfr
mj0x33ZqyUin4rGbsPp5wXivqz2dcyrWmyca4Lo84HbPsWSz3a73pdqiSs6M0sp5
UqxOp+qGxVsHcLt7dF6JztGt7xy4AS8G+I2wAAhHnbdSpW1pedFDssSwSOWNwaPp
kcvCvmAPPTKeJkxU0ZtVQifjSDVIhMp4jPYvV3CC2PzAra8DNssGNoH8bilBhQTr
cyOG4NgghquhJcwANIAj5GjqCwsmRuHdk0TUXgWX6bTVivwKK0VWwWkt70VbAZCY
zsnqZ9puXgSxhJGD9WYwzy+lQMRhhjy62fa3t4/dIZkGVBUE9E0O7D5ws8saEwIn
m6BGgkshl2IjGFYKjovZaSwIsygqaP0lPfmJ5/91v3+qgJIj5wYLVp/bLIThK/aL
W8It25ko0FZvYKgj7z1mgMbHbiMEFoMZ0gF5T6KI96ZSXq9gJsgaY5WK3lFe5EQ+
/FihKwOPQnU0ePqQu5FstwSdZeKP9r/fUpODkt0zGKGOxvyGnYm7qA9yBN/ejqHD
6qKVzXKzKpr4qx0dgzd/I2bUv9Rm3jEj+3AFgJsIH3BdHpK6MzSFrthoUVjpm4GA
4aK0jvrHd+Dq7VjtAxyCzTvoV1zsgP520yoLggCaijEiDYj8UXtEZX3wMWCcCpIP
VzM0QcgTFxRmpdY+Q3/vrllg0lgcEnkhJpMoq+qu6+OMWwLL5qbtjNG5BL2u4MoE
PkuEL3tKs6bzA5f+d3cj5AxWez8Qa+g46HI7pXAyjVGahFqHgqmH0pjPykWcgFrt
FkCiVH33VazIDpsB/wfQyEOSZcVokjIccQ/Lk9TtQ8jQaWVPJgQ1cAMXKbkWCJdu
W+0rfNJIlkExhluPS5vPi/lYXSco+1uExgLmRtxrmIJJqO+FOxoJWDonZS8ME66g
ivXN/4pj1/DpEP2AuVsJOk9lYvWPFAhxk2qoCS77RT1qHzq8kwgxe/eueIG57aJi
mozqKlvq3+QgiHQNkgN9T2nJZjljkng1XuMHqHfzXZ1Q8rvYSAt8SrNJrITabwnK
aQct6yzPoP/zo24GTz4STWhxOGL9WjVh4tkizO/YAVnkSnlxacgw5jpJUrNq2KKF
3HcFSDrhC3lStSNdvNIbPFp6lI0KUr1JgmgmRdyt+/N1r4UKeDnKNbOUKxU0NNcf
R30NSRNoV5cpAKODTVbz63asHJMCqgN2iipADBzW95XUJ8UMJxjx8hp0JprE8ANr
9U2Nly+MgEEmJTjDbAa3FDVAwtCh3zz7XSXPcanySrZr4Xt632MSSNxi1w0F6mP3
IlB/2W+5dF4BEMEp18dZO5bqFM3GY5DdieVt13mqA0QDjBxt35UuEHfYGhBshjnp
VkZghLAa67e1aSia2A34vRtIuV+qqTmLOV+QAq5tb+71SlB3fyRRT0MTyySDmlvF
kGArZH11ECYjh0DP9UzyiIaQyAydfuZO9L1umFBuP5uZcp22LOtp5ZHp0/uY9sHh
IwbH49ufW14bb4fLZwxL+OiJMPBRxMvEQhETKGMj4RYinQ8bV7Ur82Ftz1D7TLyu
zbDWwbbY3mPv1ikBoOxU4YfHevh/PtRcFMszwgMht/kOyaML3X/p17JDQ0mYmYG7
Fa56erC6PSU0w80hyeJUb9tyvWlKq9VPxVlqQP4iE6myimDRYD92ZiDgTMlFFi/h
LuTUqNygJbE+3FcpUIKck24WbOYcn2/6Mk7bgEJ4gtlYqTLXfia3CMgkqrnVwtuM
lYmASr/VQyIsQA0QyV8LqUaGZyWEs6nD3zIo9r3cLOYDR9vMPke5/jJmaI4OnMTs
fwkTJ8kspY57Fnwhu/kr5B7jXBjxkm5jHMjDn5OaOZWthm68X3F4/BQUKVoU2s3o
okOzyvIgEaIEyCMPSinT5YKzQeoMiJIiOQat5C6XqsG88cZU2l59uJn3I08dI4P9
lBEP2jD/4QpWJEuBUnqgyx6o/53qNWLbR2vbkJ7Nz7bHnYXIByDw8Dc/m389S4OU
TY2qO6lXZBlsLvo0vZnW0cRBUgtkt41HOmQgjvGkDPW1f9unwv6X4TZKGlxixcyl
c+38ZrbmjUPWOU2CkxGwWn5YaWy0NwZjJcCImd59MBvE+WObC5Zdd/UaK7VKeuib
feQQyfuCYgG0aWIxKuqz7Cq0BKraLnA+M6nJR24CAcbiqz/a4TcU9EJpgwo+WWlc
77bnaFDlyYHOT+0rRAJC313gqlVc2+Y21F2D4qVNtM75S0LN0H706z/tAjd6jkH4
OMhvcpKPUZVsDNuc6uzxnV5IXW6mB516FcaqCuWHd9I1Iz5ojSVL+o/wjddNHjLF
9/ED+c7+DnIX2sfVV6qMoy50miww0LliSeDMeA8cgnCG7bOHCyvsFgwXTNraqEts
X5Weyre9EsXW/gmwnmfTSjl6zuHHn+F99c0NwSpTJg/t0Ara3crgLe9wQpD6vagk
SC/Xmvs5x8XgGlpBwg7gmASQPLtuTerI6ijjeAhulgdcuZjpazQ+txjG2tleqbP1
g5keOLsedHbRLSGY7ghrJpUuRIYNKHKfBXw8YwaUJhFgcU83jfxB5w20ID1R73ON
NnO/67YBa5o2cuAwxEXxBe8g+AWWzXE8fqbmyqdFTXvPrX/DPVXj9wbQYjJwys7w
AJ/MyBk6y1ODh/Wlspc9nYKilQGhezvpqkBJVjDVlCJeRvAMEkXBFm/Ob/IALw+C
vSbVXzzMdNpnR3fP2VzZrTlwmg2rcqohnQ57WGyRWiFluG1nr3fYW4L4I+wFT/MO
6OM/B7EdUXCcri+FwyzlKeYdfzdzjNf6TO0trrxLXz7mpGy98mAvDU66W27uO6zf
o1Nf13XfSgSiutqU2DPAyUnNrROErFc2//BSskhaCcoJMlzcsBON8WLPw5s1zTry
gYo8SGq91lI7cigSsZA01ULMxli9sdmbxEd9La/RqUzyz6UTjTXf5Cyc1dhETFqO
tM6+vgEA6LD4z6B0WP9PmGVKgEZO07++VEeC0ykpgRQXSGPljXmQmbh/tewz2Toi
GTl30NM/TG8mckUUShN+JUO2j6uSteQPvwJXO3mxx+smeenAMTc3pvgTLkFhvywz
0butHWtZzAbYt0C2WFaqna1qN0pABW8HYe2Z2Q7VoJ4uf7dtkFvpOwb2bVIK9Heh
mEFPNCsikgeZk/HMQ942BTFNi5UAIksm5/W6hdkHqhfB9q9YOZtgOS4mVJMqyzPP
Z6HoGkDtVcRzEvA2tgX98gDieXewBgXYWcSGMwc/n9NU4i2Vn4Jgondh5NZSuTnS
V6nf1Jkb/09Bu/BI7iGKcMTBWJHvX8uGiKcybDAcGJnkGR0+yE6T5Xx269PGcvgj
Lj4/qG+vjjquNjp7RTL+FzDmiTKaU1o39EJ+OMYsEVR6GNNgpDs22Syf6Ei6PrpH
BpcDs1tVaYLqsGL9+ylNmtisCqNqkUDHEOIxFXGzgSYAfctrfZBjjIsiLdyLpuBz
63KIS2eB+7HV323ICVl2g5EHQyYBkoX6CXGvkSkQeKaUdsm/il2XVN2Il2mZ7Imi
DT8ulVHkvo2GX8kHo/CXCVv7VcElkfk9bBhJL5I0MJNWZ4weYuNMbg9fzzWmdX3I
2+q5S5beVRILmYxCfpZ+P469nkDNqca4zMJ94IYDtcJqUeVnCuJuaeyqZ557DTZt
IyJNTXWG+ADfZGeJsPkzTe7rL2x6O812dZclerdADk9QCBn5qkoHeW4vXlCx8W2r
+AVxvdmQGGi+zYRUaSioHKO6v1nocF9AMyGuuRgV2dvrjzlPQjgAHPZTcc/etSVN
wifCnQk/vIntkrBBMZG+ZLAk+5rJbsi7gwf4M+3fiNaEXcUNZZACBoW7+4mHbNFd
BVnkvwpuU/5ySVC2shQI/uQ8vpVvOmFerwwp5M4/Ag2lboxpokSdKS7ED5amg6YS
DX1XGP32fYbkyJpllnrP6xa4Q5BwB2Jm6wj1c6hbbQi4dIZbiLj9dyD6P5myW40Y
SRCQKqrbXN25dUloxuhJGNyY3GO4lh4eiJeuF6oBPGWY5xCkInkIh/qXGF+DbEfR
oX13Gd2l63Vta/4GiOjVkZe9FNRXnuC2dgzR4KRopIGzsyQs5U6KSCCXNFz2oAQu
gQ0XQTaRQjH5CpBZCsFAh5oWsnHxj0tkYjVrrxbW9emeXIqVjM+su8YcPzKeWTXh
DfeYb0CWS3Sb57PF0Fv0LrMnF1V+CusXqOPwnWjtqd3/GBTHJ40UpUN2LRVCssCN
QB8XNo6Z1Z33li5qonx0eMbzkTVQrxd4me4FK5wfn0y/svwVqkSARMfxQRE7kFtZ
aIxjyk3rim32uJsXkcVhmVRiyHhG8jvVWIDhnPfepShSzrlhLw8uvlFGKZzTMmFv
BXvowLu78REoCYyxDaN9OJcYN6YCUfAFaBI/85OGVQ4C5eorgK7aQA9iI8/X0CTd
1t4A/e8klBZYYMUxCHOYtS5xCn1PhOswGwD4Q4htuFOdtYD/TaSiQMd5hDiKmmHD
EjqUv7bDcZ697avtKL9AuKVneJ5Zkkj8GcGx6J2LOqOZk7FA4xsFDwkh/RA1vz9I
LRk+w5RqaGbawAEXlcjbH0IQ06XMdFSJfznxiAU4kVcTKlcT12e4nh94mEsYytOX
Ub/iEiIyB+9cjvXEzQv+HhZzlJUtpCwKdADXBLS4W61vgJnza9l56tw5Zk4xALW9
uAGG/GCn5TjTzH1sCmllRPky9B638N0x4Q+HKp63MkcRDOubPLJbCTMFUFY/Pdcy
2voI190m40ucSJkrO/8bsOFuB8ZyVkzYkvVAK3nw2k2gTull2SYnI/E055GNTPcT
3UPjOCTYTfiYGH0DD5mWKD15KUYN31kolcwRETPcOSxxkuHXpq0puNOUWVxL0IEp
4Awpi+Sk6/FROAvfb/UXDVhek/KqiendquUxFYCEHp+p5b4QIaFpVqSZjKr36KeC
XGV8ahD8Mz7KGMb9EEBevYi/hGNpw7ILGpFXE4pAPo7Gna7uGK/PNgmlt6AvkZp9
FWRlJqma/OCdbn0Yk4A1ljruvTvLbLq5SMyxUoppODfR+WpduJJ9pGLN0IpZ5M6v
+6Ax094X/3AMjwPZBVEMHupaYvtvua3zI6Mc9wIXatRJMI4UgdjsUjFmQ7zIHTNU
TD/LAgQGKpPnNO1ONr6ukKyy/bFuIHh+4z8wRMH8Ysr4u9nob2n2blMzlTsaxKWB
fQoC53YYUUwFMEDvbxBEyzWfaVSvNaSXNcGOq2iH/Lqu6sGu/yhLJF/xs84LboeY
gt0BVZKlDmNjIBcwvs5gkq0cltjGo7QM4Rx1BSKWlU9Dd+O/fo4xbaRd3+L8+hS6
8ZEySo8fZF8RnvMis/Dw3J5pWbNZgo6WRxO//GuPvtkyLx3pY1DbOtuWZuOvzAs1
Cx5+IAfXmeV7AjvkvvXK9l3yJBcz2bB8KG8Ygqkn1fo2VH6eMWNsTsOe5tOVMyP3
OMsQGs+OhK60qDNM4tVQ65OQlfgKx17d9atDfZacIv/4900DXuzTd/ug4JSMIHRe
V9CXT98MKoZdPWWoHLYZwonVfNDDytxnbQjIU4hsDj2KYfRPT0BwocZTjnuAmGIo
nh64CHoS8MfRyuep7gjGe0vDd7P6OTd80XXsfMeUVDS6sqSjX6bWrwp0+LrvBMJ9
/cEYPmg2XRBdbnSpsqIq5600YIm6A9ZN11bkP7WF9kss2lCy1mnTInB2dN8H0z6a
g1uCEsVNrQ6pVF+TV0T8GeYLoHub9onph+b9uiVX0g4oAZvU97+Utn/P59XU4K1T
Db3atBppB+NSAFPNRJzRO6WKrvokk9ID6I2XWgjceNXK7xXXZvciatujN+SHE5GJ
cWzBFJtzn4HTKsNzst3QGy/ei2yESq6Y8F7R5aMEa5j0FbYmWDP93IZdkdU4Hxkr
o3zje73y1oMSba8AbUA0v4Lav0sYlhisVffPPpcn64s17Ww3husXCt0wq57VnoUZ
GVcTGMlCevx4eKbcnBKa1gLfWMOCe7Ilr/+0lU+3c5MJqRW3TwBf7RpScQ/+wemQ
BYrl2/PL5Q2hLo3jBXxuxRdAs6BSo1ETQm8C6daMFaf6ovN1iaDmwJeeWUqPh49s
e06gz1FulkdNtT1rbcby3PzVIu8fZWX0/HOZ8DX3NViCMNi8+vnAGbCh3F3omWqR
kR6EQf7lFfNNzLvWqEc67nIidhJW+1F/vXcfc7r1U96PxcC1SMOI5Rw5Npi6rUg1
bd8Dl0zWaack7CmenhgZ5kSPjqiK1lejbTzPAffLoIrv9dqfvAsExS85Gi7ntV4V
k+otS25BYYUGAJtwh6yx/4t8d2H64hrFAh/YsKd8EzigDdsl9X0MegF/TD347rJ2
Bz9S4eiU87TvllEZwjePnv9z5n8zzmfyj5fb4cLIYDGastj9W6acxy/xntl7KdDa
MJrGWOB453fqjOeT68nlJJF/MOAkdeUlytsBNNhC1koLJIaSSi4k7ilD6AyYkavM
nvDbnW43xqbgUhDG21+1Em9XxtM/6BdGvSpjLIM+LuFTInsscbPTIIvFsrTaKIo8
QHedGhE2b1dQ+pcDlEc0J2uPqtH188ovBZyHnbU5aEzGjfNbzJDcVDmdWd+RTDcz
oAr1tlHKc8rYgU96vBpXn31zqn1JimAsvvoob2D0uGGv4/7jX/LIztUzG+f1pov7
xX6kMAuerizeuZGLLHbU/1Ay/uxicAnKftbXN6JILZPVZ/my2td6fcWFNX9uTC2S
IoplVm6j1Eag6Wlca4O2wEtHfUaSfIetO+Nd7Ic7EeW8T4ZpZ+0EBys8N4WFzVQR
IvI3sXSI1g5Y0MUEyAOLHjT4vt6oqIG86eUOcYQBYLHGbFStP1nPKh42EAlpPWWJ
r+34aHyhbK2VmfZi88eyLYqiCRmL99oJeKebpi0X1WQgOT7nVOIbrXh0vItiYRxM
u7UytbFh6I5e+TcT91WlhcreJ9reOkYmlA7QKlPTtkbysS/dkLYrQxDd0CE03JZU
glWnCjGZQPVQ/d4yACLLi95YBXIro8BklN+Upz/0Q2NecLXhncFVbulSe+JzwJgj
M3DofAQSSJszetL65y6XBkf+9CbNI0jeKiQhgW+Bo7/F+bgiVKFYlEtt76mv/OPe
P6Hf3T0YZd2T0wJHRlRWtepkRt/qT6F4GI8oM5Tsxbt9K6jOylUwXEPCQUgOTXum
aSSeKcyheh1iyiqe3uXHVrrzBooApmZzQ7AfQ8j2b8L1xqYixPDmxAU1OYswop96
eTZB8dMeBVeNY8NxwOVFVEwWGmdrgG0eOxXPxpjOdoyVQ6C8pnbaywHx2h1PbbEZ
6c0WO5bjV0TXrjyZlciqTj1o3Kiki7u2F7UDLn6UJ96tj4hX0+aAydRcbXHyjPOG
stXYJgbb9T6TPnUjtMeXxhcdztsAZzzVWwfSXU56dge9qWgBdawXAjWjFbSh7vLw
Gk9f6maubJvJO9bapvWDWi4d9lX9fqpBJjSOB5DzY7MJiv/uIl6fO9pEyBYT6hAA
3GLwhqbsjWV0JqDiv1OMK0yk/LMGreIZxGuCP5/AP0h7iVkBExFMNibpDqDKGeyg
yWLwwRwxJEC4FdISpHR4rOjTR7XZksKrkAIbyLLm63fh2LlQ/f4Dka/nFNbqkNFZ
NPHjvao2Ff3Qch9BQL1tMdXNaXOvTAPSEGtvZJ1sybyqyLKD9yFrGqfF6cUgWBo8
5V/Jwr+4SziAQxhp6AvYW4qvfHZpmKYmOGx57ZFUnuc9UcmVLtMSqjUkQXOu4ly8
CQ4Y87hh85lZGDDY36E4q3GUHj1LltRt01sBEiLUgIPSXCclyfM3C9abv3QJFSgg
qyS9MLzR2A6tn4Zhg54cP6NP5w4/BtnzapY3wKdH9i5Ksx7SxCbxYzSILaFfa3N5
cf7FdHZVk54KYnLKrpSvnnoh8/pkvIo3CogUwG3uVBhk2l9q4paSjkWUMumgRLix
9Uw/xY5NpgzyeAEMQY5jFLg3Ty6PvZj912p0wB0l/oxo0ZRmpqDfnr1YGDN1QjmJ
+uFrOb/efIpM1/HFhm5bgvH4vGuCnt8H1+OXUkg2J82ckJSMUXPnLS1HSmOMPUkS
u2t4J4fa/TVVdhN8VUIuIm66pQqX/RGQjWYpCrU1qUdjFV39FsKBUA9yhKojreGJ
R1f0OXujbKHNSOco3clZeozgRL1mCkhrkVnDUvU2EiZA6L8EMROi8B+858BN2poN
aWw6q+nOrgZBjQy+ARAk6S7Sq22dTDPvMkkOFrh+pbYB6JJpeNSHrMVpCjU5Kbg3
xPvsPqg8jfiG+fvFACbVfqZ3QHu6WaRmJUM3UfBHZRLaRwKipoOX8DPuCXUwXV0B
1lk/8H5IHm/iVNaDVWCrS5GmbRK+ua2eyMi0ORpeV7Km9hmT7TFcoG8Ytxq1SEOy
7bFXHK7X09GFezAxl5OcK2aaLd2wO1ikC1x6MfI8B+gtGRhXZA8lYZAE00bYJWKn
c+TijHY5Z8kLlJci9M53bOzwGqspomlZ7OQWXfjCIIHFDiB26wPYBicYJlpIlYuE
q1n3zrQgNK5phM7RRrIL9FRn1OGldYGLSR+D0wLtezooGpz/Bnjgh9qQQYXiHFLS
8lXa0o+j3kHXssFo0P0aSurZ8dvOjDtDJ1VS2GcpBynOhctodwzkOIFrlk2nmvaX
wmZfnNOFJ1bpQpCsrIcA/Sb8VDv7pXaYMjzf1x29ncAfkEJcZccpn+mdZ0/cOP9P
sAcA4qOrts8DaBeDGhScw0YqByMgeK5Yc+enwTe0HDMO1zA76JQPhCzxC/c8EHNl
vBK9oO/4WVgpfq+835vPkwSLHNqT+fvy7vMv1rCd4u51tUyXKtsKztuE37ruq8Yc
oV22OpYAdEAxWgNlizXGV8wSI3Z/DnAgN2Diz0gtdrHpGa+Khio54DUddKXYqGaO
KJadLaZp97j1JAFstOgipM3Yhvfo+AGsa500K124bK27CfWHLg5qCIh5ocZCrTk+
vDJVC783HMmCnnsDUjNTt6rpthZOxsi+pW8vkEKEFE1bYeeqsQSdS9h+qpwseRFT
VBMHLqRNEQPgRGQa3kES1yz11DW6pC6H6S+XlM3o0LRDRXnESjdIOuYhqnKCIdVS
N10QjmaWwADHhyDjCBI5xwvGl3mAy1QjJ6foijfcaDWBQIPEb37TE0TUJ2yx3dJt
V/SrXkj0FVamHxgvBMP4LXrpUPBj9dYUU8/8i77dm/J/dOc5aqK6LnihfAOwzPNh
pNs/5Xf7HVEC414Dk8sNxkh0EMEGC+wCUf3EkEDphtQhYnB6mArEeQT04wM5JSSr
PU/BahmeU+520QNSBe9M617gsbc21z1ImLJsaDzXpTSIQ2t62XzZVLRH6GYINKRL
X327fcOO4kvSE5KivEx9EBjjMsCnR3L2lSqm+dbVP8WiHQTkvTF2cWMFDwi7olqE
o3+ISYNZg/JCauUkgbRx5XQHvmT+9yNJ2LwBhLY7XyN1bN0OuTDthJ+Qrk4GXUYP
eW+/mzrA2AsE36RUl2Un4g+oXsJPyU5AxDWvEgqntvYD2P90LmdO76AazW1SX2Cb
LsMg8QHwsHY4RCL+mox9wFIp4LrQQgYZr7OjsNm3jjZtqc/F1A/gFOiOJ+nXU3cm
tXATKnSBtxx0eE7CXpeSnwqMd6rlNt0/Ik+HrXS3i5Mklkm1TnDlCRLRu8o+eRjG
7jHiH8CMtPe/+q7xddxwm+wXHXeg4DLJE016F14UDUd18An8MQRBiFr+cDsbxERy
Eo3uPZPjy6QXfIeBcKQJyn7YI1XFjF9vXyAUQptAfF6yj5yAS1Pby39Ij/GIKK4n
MAiiuoNGAuFaPXWGUvudfgMhqdjlGEVY4F9bdv/2h4kXzgs1ktICLAJvSGef4WdT
XDNnbwAiLIJPivcM3zAAQ9OrPLAy+b9YKRjr8AbozmM0ezrHQHXo8i1+WpFUVvXT
7iUzhpxoViYjn0Nki1WfqGK2JBKXq0sMA3Qbr2j1y7+2Wf+TAneRFkL6O3EOmLbY
lxhMkM8M4HPfEeXE3fXaCNM236ZKNI9iJKDZWi3Fb303Fae6NyKeJIps2sH4SIoi
yKGi4gyLxfU77PAQp1U4xy2pfhxXZG9znb5igqJt4nwZvxHvdUdnbaTQsoRilAm8
IcugIIf3t6fysrJO6nMzvQGsSJJXcSsLyqCuVG96fRWnZieJQPY2IATPKgbpAL0W
WtvboYhEgvOZazW/jI8tYAufdXOTjPnRv2S7NgGKJrinHU14nFA95CTG646Cyihr
bmT9jFdOqEE1Xw57pbnqCGpTJ5MAobHbvUmdbEbZgIT5ekVEtJqLe5tONeeroPdH
t0xzFwJ/rpvLqbSn+feoYbuYXmpXaw+/bSMc9qADjVlIYH8ot14UkzjvkHHTrpsi
oOawToPITtyuU8QAORIKR2NSaeMfb9ee0zeh0aWtEcI79luxmUGD1t0uXvUd3KPp
4UxKX3hHgmk0zwl9dz5hQyZqIWColEoRRUUy4SS3ibHMSRJF9TKTB69h5iuVFKIR
1ODobAQ6OCkqWVAHPj3Dfb6C5Cjvo1CR3YxqFnBYJESruVjB3fuSmnLvzWEYvl7p
9AMmyferbXCOz3/mjzzwgX//CsjvaRutXbnjRW/k0gryqT0DH+1qntvE3q0hWo5X
FGkIKnFxUv5WfPLeprAw8VFXQaBaqTIkb+ilGTbaVZgg5fNF1grLyT6ePNMAW5aE
b7jer52DBqwkN5n0p/jm2y3S9oG7XyoTD/xNObkj9vZ8AicZwiT8x/2YsA0N8KsI
jAJ6cyxIWuw/PkeEIUF9jTCWI2Nk+34xHVX+L91JHm+h8RDmb6+rbHLblkSTyo6e
EgbF+3EZDCTjAzJmkwjPiB6wOHlmbypcG3kmfHlTFot8VcwqcSw4UxEcZy39PJ3R
pdmqh00xT9vaK9OUK0rB3tYuD4Lm8I4i/K9hUTmSpzul6r9IO3D4HAp86PNUrmFT
RdhCxhdJs2IV+Gb2PAdt/ElXPhPdulkGc247UkBKcw9E8VQFELf8cSp4nN/+fbfo
iMdAhNP/+OFzhFDJfb8WtP4qTFRUDMT6ilSlEw5rwMJiwT8p3Rhk6u3DCtXHtbsM
WLBW40o4bte3hfsuFxpR3RlZJWJc9jOCWrbpVEj/X7nU2Y/eRJDkkBlqtWNKrQjz
1MiaHZJhxpVMmzZfzYRrwZQFIBML4PGEwmRztNTFlNcH5aIs+hrvL7c0Pos/7O4G
XW9VTcoca/Em3ENt2fS57CkFhzo43sRGXHSo9ubr/k//pleo5R73ytMdK7BCdh59
emblilgzhuW6FZoWj3V3EqHYSo+Vk90ArYsNsRPdiZY6Xc8gioLIm4i10jpp9xWc
Fks7k9P2dKCtdrmus30Tr1lfUhWPd2WAR/f4iyIBYR6bEgP7Y2OwBL3C4PdLNIzh
7GqRB4BSL60ZOlaIjAZ0qc31KwIyoMMbqLjrQseV51MzG/X2HN3hJG2TZ/ZPvjuj
T7Cy2RaiJtQnpT8UsaOejviePGrKTyUPuwWQsVbtiUc/nScDZo7K5AvWhASIueRt
gJX1u5cYvHh+RL7rlk0yzLu+bUsG8hAv/4RSJkd7ObB/OJHi9CMpxXYJOhw9K4jn
+Z2PO8ydGLGezRLMJbodIYcEgVMF1qFYpiiX56O5q5oJBTH6CwlBh8kKSQAMU6fo
xdK9vaihfEvFTTOsPxaURmb1dS6it/bL4dyDqrVswyLt23snqrjYNdoZycTX76Y5
XnZCJS1cT30DoWqY3k2eHP8TYUfA5FYO03cp1JhZ5venhds1ykkObUc9ra8y2G4d
GDOVqWDIZpTxzNBuYbDuNqsZh0d2/03x4vzp0Tj6tfQjEw7RfpcfcVEvFKDGLmqI
2fhh9HIOVONf8iK2nGAdCiX/swwZ66CSnurSKF3J5v+vbNiBOyGOWFoPNNdB9MYn
le24rf93uxDkqm3owcvY3VfE3Mt9VFK4tos+BzpZcTqPrHSP7wq/ukHmix24N43A
XX9nf560kLZhQXmkBjGja4KVCTUBb5GZ5VOLhEbjH2hmlF0jAcJLxj+SAB4qkWf7
LZzQI/gAUpqyhJhX06od//GpqW9bP1aYlhK7dmTF+WUeKJc2xvZr9VkWxydse7us
Yt9wRZqgt/ZSR/BDfhAnJqVoWv6o9CaPN8iYDpsbLEeLfO76jjFejvW9Bb7ChRO2
7nXk9tkGpfU4YkF8pEhZyHdEEI1CFmuIHxSoNgfLv1jxz5rHLZf60RY1MrkFiALX
xGdMP1cZSqdzGWTbS+UDe3pVdnvqnYzkvMlWXyLfHa9GAfXJBJlvPJOoUrezd3Om
xoStodTyGu8KHhC8m5YGomQ0QwKmLT8SxWeUPr9Acfy6G2dAtWFeOjCTDd53WbHV
Za23CI8LAGS0wozf29N4Hm4SqZPLX/SvLYSaN413o+pYOwdmMhksvz1dEtHHnRWv
nTCgT2m6k32I9QQCJRXCIWp+ziEf7KYE0eTpX/wZO1ZNpGqmsVff/C4iz/V0CAO0
uxhecJQBZAyWR9fWHjkJdO57Bo8Efsoss/SMwh7AxyzotxDdYahxCFFqWtHk+ouO
o+rfulwG9KLUs0219vpZ9q5eJ2cFVvs2q9ySJVLPHsstYkm0B7X0HW2d08QlddNh
inSHWwvzDdxvcDloqrg/IJCCrsIx0I9oejImeicWPBIZmD1PTDnlHNEgSa8yDq0I
Lo/5+eYUgSXSS3OwFP8WXJTzklgdzkM9w9KqRi6BW1a1eSkMYQEMgjPebGyoY410
rWVR8qLIN9AsMu+/EEYKhbVZoR3ttG9LGGu58X+m7EhfICen/E8Rnu5+wNoLXDa6
UdKFUZzR89HGR3fHmXTbShgnNGbFHqBRSJ8tpPXpWoj3lGg1kaz45XMT6xeW8wzQ
bAfXgJUpL0AVuTLachITjnOmcgm7SPmRPdUNHyUmFMn05ZATJ0RBldu/dVgNCBvE
EwpjIgoRwGYLAwPzLTnxJC3HlFImaSTm/RQbbwQ2YddVrGjINkqb/LpC3eDqYdvZ
mmzq/jZVqh91Ldr65/x3PfNHNcym645hx95FIJPZWrHgGBBEM1OkUwvnqtpd7nBI
vgmYOUScClP4f/xD7SCT6iYUCNYJR7JJ14ld2IfNgSSI10e8alK/WInf8x5CBGnE
sBcoBNCVf6EJa4hM9ql0KNL44ZFHdyjJ1kM0rswNdsPMCkl690XN6YMUz4Oog1je
AbgTn7Mz7d4SZKD4V1DdAXZkgIqX1Wa3aVLn1unvpgOCUNUU1Z0j3OLt2dS770E/
pKJM5/qbcc+CSKByWxHBwmU3SQO1/kahcV86MGbsgsSUkCQEUNCPds81B+OwGnuj
276c1M6FZm6JWcbnnaB7xjhO6iQoPaenv7LPTfYfyIDK/qGs1MzDP6aZvrHSRa8h
+wydbglD0bNcFOx0L7UyjylndCJmhHNagNGtL7wmUgTopca7t5mk3I1K7N0lklTR
fzrrt3J39IJK9QNG/0+mh+B89vzAcBSBngL0Wc6zf+ge+z/WKUT4pFDcXVqDf+9k
4siuKYkVn5gYJqfojjO0FEPRmAu2Q6S9gIGmje6dXqTdPgh3cZHO5/uFFmcOfoQQ
wIcUfsUxXwXNqGEWwG7U6XTd0U36lN3h+u3Rc/SC0q4mSDJNq+yIzx05D7Crxyjt
IbNbFiDZlNWFSQfghdpFy0jJzt01JWTzTixniRukXrzdD6WqqYrAtKpEjj6Xu7HN
NWPFY7Dks66pBw71YJNVCugC/ItxO2Zl5MRTa8/ssvJxffXFgtBBfLnDCDJWDjqh
nPKwvLntW3ftgaCPq3az2Ir92vpXPTQXtG1/tn3ZaMR4pZLhfpfBmh4TKTCkqFpg
k0CozFr97ayusDPq8xQSMr4X4RIBTi2Ntzv8QY4+xV4gRpI6c2z9zxfbuSj9Mb8y
gWUWAJkVrfti6loau7M3G/NMSWqpTZWvnoh5D3LPO/KLAzff2l2b94eiOWaPqRkT
S2NNYEjOuM5zbQRSLpsr93yw2i5dOTfL9eXsXBwhDcJrHn/k7XJl6pf0iYWc0J3D
43knqR9/6+J58OuOTuKopEoUYg92s7dwdVIVUCj/VtFbJAa7Xi0nfUm/17+Of7cN
bBCqFhlNfYrzdv3CPIIKkL0hTWeP0r8V1LwGunkkxkplj8cAKK6z5i79iZeYxl/D
kWaLelMIedAY6AmbcUw1e25ExDE/REgFDAvvL5JqpZ+WbIh42u1KT/hLaz8EZVlV
Bl3ov0zAMvYFUUa1Vtybeel3ztRAcB9CYz+Mw/hjMxltm/LFQwwzsJ/bOVjOZxoo
ET8wQyKBzzzKfE/9x2tyk+eFcYznKqBgoapqJugPiANQESAb0cWnV5weYmg8Cmbc
0sxMalfpFYQ1Ez6Cjx7nLx/eHloN3GKzzd53f28QbbTV5hKuh92IRDutyFiYKpxE
OJAA7I+eLdfeFs5nCuEglFBF9RHUBLVwXgMmutgKCN7SkiaUMmavDzS2bmv1Q2Jm
G2IgvHF2aK+AaIwFA1q9D3zTFc9uLWr57ijN8yf3A7SukltfHFA2vhIfxnZZUPRr
gPVxod9TuhO+8tWq+I5fIB0jdRonNFG2KQm0OwcttrFyJj/Rjxs59Hxtu3GQnZRN
V1HvfIESV/z3VNUO3Fc5XbJ9nffIH6pqpqBNpYzNYH39eOv74A/Pe4nFFlj1DzCV
8JjNrvCTYUrvtwOnJtNZ+E56AvDWilmZ9aHRAhf0bFtNu9OFlX15thr7S8q9NEu5
ZK47avGNV2z37DevyOlWsoZynmUPGfJTEqjDprvLL/g8OcbMve7PQNhmzvH5dBLn
vOlpUJ+cIua+bvBIWT1O40isqClNHXDwY4tU7OFSmA7tzW91ZCtW2Ia9NM06Mhkm
RgBoVZweHmERoDrZTAmT6lN4FEVRlwaR3RQ9fIW7+gNdP+D7WCZPKADBf4L3ekGQ
bsmOXb0ByW2K6VRXxSxyedpvWD2UL5jj1nXk1ooHhtXW1AucdxTSebM7XRutdL41
A5MmCSgxYCJJU+LizCuwcsPI5BAb0mXkFQBogSROv7HCPcKa8xJMGSoMxAAKQfj3
JGOWA7BV9c30ngBktQaG9Z2VsZ91GWN0Bg12cqEFrrkgTX16PUu6oaQC2chdKEam
OctkNSRL0dfnAjkWUO9uW8hpPbNFlQnICFQZWrTiduMjwY/coSaCB0aVAsDMKqpb
uAu2/3XigdXesVTObkqqzvTFnUNqyeETWo/gppvPYPEHCQjWpP/1NeW8vDW7r27M
nV0ue9lNsla7JW++Ryc0GeT4Re7JcLdw1ISAMgd1Rl01hZp4GwqRF7XPDS+Twosk
l+dqL3Sly/Psnijhrzs+ldlj6JZjkyEktkNj0Z3AKDwKS+CvMKAEDVlSg0eg9mTZ
78MubMeC5BQxA3tfMBxBJ2oXZALbwkyt+Xj8WeIBEqRWsfnHRFjNAox4m5OckvgA
fqzKrJpKhRcLJyjmF+ShZFIoNAzgvLQR5gQCBBcqVk4v9Fac+FG/0N5Fc+bQmFFp
b7/rEMjZeZApfMDcDNfNOyWTmGMBEZKpiI94ppPqhtOFdoirkS7WHW2av5Ll3c5n
+cN8FKixDBdvRPQ+lxA30BfIjil6eTG1zrvNnvDG9+7fSdFMBPtflQ44qBzLW86T
/jW0Jd4dgS+6QLymjeR+PlMF9EKsNfJf5v89ScwesO6Rv4aR8CvPpDf4GvTBwh4U
ofr7LaV5Wo/wwoLdOj5iZ/tp+V5N7to29AQx/s5zsJawQPQbqa0SyQXQxJPLDBzh
jPKpX5hCFuxLcdf8jmmSYgZ9bKQ/Zp4IO7/RHcUDtuaVr40FZLHOSE2JvJDenX3F
XjIJubbx6MGirQmM6DeiLf2vIAbLKYobvW60LB1Nl58wZMVL1S9ioFP/lQEJMXhf
AqIo7kTNzWFbvgO6XWQc5c1/S/8W4hSDsNB3vfNvGT1wjbYsMPT4iVRG6W9/gSn/
mJZ5cXI4JOi/Qni/WRCR+1R4RL5eC7iK2qg2nkIMMXAYe1TT2tte5Z6EM562jbpQ
XsO9vY8aupD6TFyMG+XJTYV6UWSLBr/JZgv8/qcXZMX7UVa5oYlcnPccKSAFm3B1
TfsnBUIwLmiN6k54AIWhAAfG9u50osoiwTmE3DyQg1UevDoXQ/sPfaT/lyiWfUzR
cAXDPKy/cCud9KNRafrQbIJSE32s3Th5kG41t6TnBZr4g4cDjdI0muF/KDHMrvIz
z8CkDaIBtCALQj5A4WNl9dWv2XOUl60jLGNyfpqGJLEK3Jm43QkLosGdJNnoxmfn
HnkSBSvixuGJHr3IxOY3vAP1MW1h9b4hCi1KgDtd/a/nWNUpqjcTSmD2AbfCcfxv
Xh1xgEinoYaEwV5EBCMTnbrcuOmLp3uEBq8PrxZG0MuWXHAi4gOs9m1K4LLQJhl0
eb4Gb/Z5DZeILxosOj5TbtTvsF5kG3w22wxEHHovIDJT4uA0XlvEQFgoWq6d/8qj
WPIwPFXKrxRAK7HRr6kpgIjUCrDHk8eYSc2KoA2BTyeybFMxqH4y95paWcB83JNv
xMjC4ujqLJ4BkfFZZBWgrCHutRK2uc5o+qSYCub1YY4lNkUoM0XTXxLTCvBqx2oi
9jOgFh82l8KbngRqDQHEeFkd0g6j9Zh02RnqkfuM5JNxFno7QSRiyLIBXNEzvHuf
9Sr0uSNc2DJgZQhHm72sMdDsuOcJPPdv/9DEEp2WHq5yzy/yW4K9U7KLMZyk8+ZM
Lauo78lTOrt6/gAkWJVFC0pi3MYC+FD127F1Rx9d61FV0IoNzKVwYjlL6S4CXDdc
MvWEpfSzaTVdL2bHZL9UF4a/WAumFltUsRWBswx4YHT/IuIQKe1kY5Ox6tBCVqKM
+bp/3bIBLHBor+Sr+zdpaIKcY4AMyUke0IflppqIHJZJ4mBbJmgaTLj+KqY2/qgf
n3q2zX8NMeEdL5GcMMOQCdn3V8cRvBJkTF4Pko1Vrp0w1/2Q31ig4jcdpX4n11zU
MjEh0muIurIWDIFjvhmeZ1RX1lzYaKnygOhKvJYaWUBBdHc1DIOsA6FAIA2WJpPN
N5Mw7s5HuLHJqKkLECs4MgHiRXsLMVVvNg02issMLgIYY468Xv3LWOaBUeUtusEK
xQWYXtsMuBfZwLhmopFD+juwTmLrCyFLmVo94wtX3wWnjnORKYruHlKuabePKrlu
05SsxSsHUdUGcx0Urpu2yWT+WPqQfkvTM3yY0JLc24H8w2e+vlJsIBEiRK/NmY77
C/tJTkbpVYWzdS0ImQd8E5zg7YdOPTuD9FUSHtf+KdRRzSdiezOOP/ECKH16mknV
l2pXI0EhnPldDSNBMd5tWFWEPT97T3EKlB10OC0OLQf+wzhBGDtLfgGacEr4/Lsg
In85EYCGHUBsiNi7n/fkwPFJXFCy7kF/0yNusNmiNVbwIQMPSLPQOqyYiNKhGZ56
8boYqln9w/FTjgfXzGSBxDuj6hAzbzmC+zuQOccwThsuUq4vRBban3BENRCTp7LE
XR3ySv0NPVPZ5aWBpMHy2UzKeVrmdBKWfFTBsAMn2lbkuQ3gt115XHLvP3+t0yYs
QHo6wQn7OJU7KfV8Nzjtpb/z+fnJmOItlRRxqUH8oAP6A/qLtJkXn8Oa/Bgvf9Kn
8irintYJL1J7XKzbBrFaPqdCVp5fc5dxtH4HWaxtivEOWWD3j6mlVT9Rm0RG6bJ0
l95iezHh93D3EaoKxJu8oH1R2yiKYHfuximiA+GKZgIMJsvl40dAozdxdG0fXGGN
m2d4pALsPbO8IBnat2djseYDuEMgfValM5EoWOJjL8J20GJ3V+RAZVqAlN8KbMGV
rz2OP/yC01+DWkPOCNyCPU3zbyoKi3HxvKxtl+JvINDT/pOU6CZ/c5WI4W7Tz5Ft
kj82NVY+2TmocZXwYvoo8qCq3B7j+/lJT1WUa0kvWQQn6uuFjA+RG7NWhmomwEfC
PgCP5Rb83bf8SwVBNLYpfb9RJVPu/26LVDpGWBKP4hri5RYFkmhkDmkh518aaLEQ
a8VzXzTu305Cd41ZzFkWJAoryg+ghei3Bog9/ohs3NWdFfmsJWELpJGHFD9KnNHz
y6Tohs3SL4+QKdoHzQfMNB+8xDxCQTGe8s2+VW1h9pi5wtJuLUE8ws/WhufNqqCP
rHdji5IhyzNpWBMF3u7ify5kzGPJpmH4TOzeFVrpdqdQcbs7ayCA96R0tdbxCTRY
r95Bo3xl+uJgv5oFi9HK1LWQ/7Y6Pky9iSgtz9my8VMied4KAdJ/6aE464c4gRLC
og7m/x64hzMbqskGyDldMfwHT1przqJ61trCyWH7uNsNvk97mibf1n0rYXQlMOVL
a5gmenBtSMGR4kO30k8wYrTVGAun6iotqXgCSb1e3PLRkVi/Kx0b5+D7MTgY2i1P
+zA4ZE3Dg1Ve4g0okO0JWxF/H6I7IAn4QAK/Kd7e5+Vtm/sGs+oGrz/wBTLW8wJr
3U0mraZCYXDz7n0jfC3+Qy0O3fhlvUcHkjUUP5B8q9nOlKroKJiIAK1i7casJpPj
xLq/nmn8xs0VC6ptbGM4aNDyLDo9dOaSh857I5U6Gqwuanyo7hckMS9Oeql//MVa
3P6WKCeb5SOH846XMaFAPaNgWRwya3+iK2Ao/ogdAI48RIwdr/vbKZQbdiT/zrvA
X+ADgH9BX7xunFWYVgQAa2AVgD3aHLR89Th052SdGkGpGdFePrDunGArpxN8jlES
9I30kCVpmarFAjVY+vwy8msjSjLT1PIph0MR7nv5UzOqDGyTgTi6NKCWzaAAIvnt
3CKPPF0IM0RLg9V1RkzVzA9B4fbfNpgBM9EcPcW6iFrwJzRz1SMdE6knGZQF9jN5
G+PFdEN8OoXfazR2c4v2CXPFm0ik9CWd8hgRD3qXqN5W4I/dBJZgj98/Te92ZshM
xpy2alsU5OR5oBabL6x99xN5aiZcxA4Bx6crInB2tY1rUjijK1hRqxDf9Y8DgeP3
oOiJhKDMrvy7X94mOzM7Xr6KyDZtigNBJ+oRRJfKQZgLWBbFbsHlFTl3vKuqdHaR
KBAQadIDiJFOA6UfiIb9Y7XP909SYC/iSZTESsIOV1DglPDVTpn+iVjpaWnG/4j1
6JMN+TVW17ZmW3qOyMkprIV8hSdNGfITyRHZFkroCk5FNGNbfzV4wGRS4sl03eQJ
jatLbaA3RPJ7FnarXCjV2TldKqUq4PXCas5n/gyCE67V+XjawyKJO+6oX67KN6TE
4mjci3AFYkrl/JPWYawDGpPJkZjVtqYwE/Mbmi1vGgcBgRfhKlhkqmKSZvHsJUDV
RilsdzjNB89Z0e39IRhT1Hzfpux1V8dj+Vh4yM5tQKIqGnQjSTBeV/UllHXPJen6
CYV2djYQTwF3voJ6WrL7ZcNypqlqHGWnS19+5RBteQ75lVUr8qj2/B0FbCf1DvLM
xXAPTJ7s1oOnSA2ENAV6fKKsJ0yUWrIXW6iF+iXDGicXRfmQY2OK+vITA6gd9Ubf
KgtUaS4bwkaoFHNS9gvpFuivgrtg19RQMAmTgnn/kwR+Csop/B+Eat+ge7f8of1N
vJSNcGLywataHtFJhnc82SV7D1fDBDvGDPZuxU/4a07muTJEK9UnkiSiCLTcN8BO
XAiMOE8r3lbAyANKhRoRjiiFlCDthqRwiZlXutU36B9Mzy+uAPpPyp23Nr4z9Frr
d6YcfRc+ys0/wyFxBigO6M2v3er2NHu1M41l8YjWaFCI/+SQFw+bmkS2i4Qsyg3A
gBr2VEX+HDAxqVPlo2SVaSQHX5Qeck2g6iiBHsVnAU3PGzHw4PRvyBAFVReu6xBk
74jLAU3xqSHMHHkwnKSCLaynryww+ySh577ENBjl39WrAhG0FV4JuCIvTcwyrSQJ
9KUEVZRfbGBBohLbvsfBGvyMXHSaxqMp7NsiIePZrKej8Ijbfs5hD1a5T/NS+WpE
CzpsKJYwNBFFJ1pRKyY2h8nShi72dgNB/EzY+VGVtZYsB3FrU+8zx7a9WJYKen/y
D93aYVEVBtlgc9WJtkXBoRCNh9Uvgzl21VP+XYygkyZR9OcEBTPbbp7cEbLyVV9Y
fCGIdv7TtiDydwPfBsOyzq0jrnu8beA/gjt5RbWWIcfDPEqCehBGVwuzBMho6GuM
drxLA4zAByBg0tx6UkjzPDgErHyn2LxkA1sYRwqrXmzaANjmSNbplPvU2Oa2JCLz
CBbyxSmf7JKjLsOCSGWOia3uVneiftyt6ZUlejifqfWZ6AVzs0dNpj2FLi1Delvh
65T0YYwJao2ZvJQzapvyHisGtzXxixDt5VruxiKwMMo+RY5htwqDNqYSj4zK5XC+
slSWMUWcne7vTuxfPeoSOYpWbG4/k4kLiglt5+CAZKqgmrnvR3aY0EpiiaZUskjI
RrKKkYN6q500vWQLiSJtmr5lGt1xSggrA2hOWWdeIB8537YAe5RVxjWGcmvugWkX
PJW1P0+USf5yKMNOVFCjF2AJVg4rDC/B5Dg5h9dap8RuHoD+zk1TuhpwFc/i8rau
WGB+STfJdqJSiFtnTDSxWB64AH8hKm+UTwdtdXkio/0FCttI0l1+0KSgiP+v0bPR
uHedqGhO2b4dlt4e8wUn2gUcTERuRdFl1imSYyrPxEjDu9uxHSffH72GJGcrL9Qc
naVxQWdzwI61ZtlIBMWv+7x4iRLOM8AhTXwCQBL0kf5sZm/Z5SqCUu3joduEqyLA
UWU+BL2CLoq33KyVVItGwWNGmbyaSaiKRwJnSmmfETQm5BOOi+i+H3pxdAxyajTr
uYsoCgwPP4aeZJ5NfE5Vs+YPO2EFU/raZT3GWdjsmS98JleolNxJg9hQbIxtMz9u
TE3rxbyQo+OG4HPAxPMQkNPta2uWHdq4JJ2LgoKvmWutVwLAB7zrluf21Wme8y6g
1KrleUSKSZ9jV4eUmZxgguhZYuOutoVKaT62SX14ffA6ikLr8K80hEdNjtle1a9U
W6h8ShJ7PcyHPKhJ01PDAr7W6SAiyWpt1/Sv+zf6XCvM0ZZ7ML9lNB+sT3Yyw2hM
1OgCn0Ai0pHf1bmpEwh+r78Zl3Q5BjNQr5PJc9wXqBRrkmyJo7bx94NePSzPXbJK
JQ9wmUvXkyInGqHOjXWc0vPMZehbE6xK90VoGDRYOy0qggD7JYPzIdRtiHPXrL40
3fDJSu81ZsnqwRCof7yIYs9pPa1YyxPM7GV0zhyAJPny5SmrMNvNYiR60Axe/slP
Ik4ISBdHq6UjeFBnOufP8j2ZgZF/QePx1ZQWFXbScKDUa0/M54QxoSfgNx2cu6he
Wv8ZgMAQ139NTA5f9y1tCDgqWpbcqzM4nHSVXtUAQ/UuOQCfqRMHQ//p6lHzENrS
lG+GxoV3N2pYycf16Kugdh+vvblJRHPy4fso5FoCkmIbKJAvEaL7e4g8ec8QKxyv
+oQLwi+rgqGtPZOSoYQHOiKjateoYAobqZZIW0OV2dbWUYIEjidgSckh5ACHKwr6
WVcP1uZuNjvkIqyL9bmw3VXwgiXI1lp2V/ZIJdzmvuslFbqKiMsD24h3Vot/6Tdj
z1jjZ/+toTDFyDvOArF3kqK5n/rYRClq+ROyAn5QYQ6u4BzUCp2qJv2Cu+0Cefjs
y3SLW0ksx773Nzl4TQGT5SQt3q+zPapf+uoXKfdWxSp5yPN+trH9admt6VO77rxp
2Il4d12TStyFDdLzXHJ9Cq6zNKiy5XlqRhzzFeIXKz0N+hwfJ+bpgExmFC+HLfW7
H6W0Vrg10bfTeCyIDyKIrSC9e+pldtkOz7+kAI+OeDW78L5Dz1QizQhEec8FQCmc
M2HfisF/IrMoh37hHp59B/KUt8raFtQGaHUDHoA/2WcYktUHW+12KJlY0uzX3xud
sYXNK+5fr08oUZkBaxlaJMHXCP3zh3ynxtpcoKPvyRtXCOmHZNxU/b5S0RcJWTbk
UXRgVoNcm/n5oY7NdQOE3jP44F7xrGnuaOdOx1RDLgAT7trpsJ48UMUhF5d1oxqu
CRL9gL+MkOqSpLOslfVoWYb3JvvrwfFm15jOU1CrTuX36wx0REY3PucSWUixaIRr
RTES+XSI7oVt/lflfRPoVL8jwG4YG2jcNaXk7sEApuqESK55F8us3hHeToCAzWNv
AzJ1WrHMLv532b0pMIBJwRu2egyo5bThZcebCy6Ft4Kd8wMKt9tP3UXJssb9egyo
LptgVJ+C31GMMk3reJxr5zSBzzXjfft9+xIBb2wViXMOapWPiYR5tNXoexNWWurW
UFoISgcV/82VQX6zn+Xt3xJBH4dVjhaCJVLdmMK5XnWm9o2U4DaRaf4kGqdeOMDQ
jokfL48FvzigfNAnop7L2iQ5PKTKom9GjHejgYNiD2J3nSys3PLH7q7GQP3vU+8B
/gwisTxWNUMwDo+xTUwYmCwsLwDf2E1GH1lQmpCHovTuw/TzGm9GDx4ZiNVScBD8
JBPIowJ7HO4mzfdLb1e7Uhl/qlSbTctfs3RwoNeE0V2ZUjMq3QsEUUanN3lz1b8B
iAIUowIC0fMOHFaL05PDscJOHtPAd/RC7/0agsfJk/bStHIe59Ff80Esd4O+wQn5
Z89d3Zrojcoz8cvCIApizy6mO8JsVjuPiiyz+AFnH+FoKgyfkJKorm/qB/qnrfXD
0qtlg9h6+N/fpz/ahuaIcyChCcsoQnrWbbjvvg6NcwfdGns8n3xPma5/b2fN9+tQ
5UhVtbu4Is5V2bLGjrKd3gPAR5oTZw6/c61jgdIP+BWKOQtI1j7Jiy4V4hAowNJ6
PoYOKUy2h5ApuR+/gvYAU8Xwcb/5XuqhA1uca7v1P/BZNu1JHh/D4DpgnrrGLfvr
hJVXQAqLN/sVvpTXF4vTFIMilbL5QFS/Mza63eSqZ0j7C8W+y0D2fW12bcdMS3+F
3f0k9pknKYXghP8YE/rNc0dtOnOZ6XMtfZ1OYnVrAJ0kcXnzcszXuDT8SfV1yIZ1
zepCGkQga2JSKeFkB2+9G/Ry211owfDcF2gu4BYZvO/Q6EshXnF04By1hgzntNfn
JB4F2Tu7RbTKHzq+i6eN1vsv8tawVMkC99zn3I8h8WLVI//b7auaN4VASNi7rpRG
rK7U/tA8jM9Qt8dH9X/+Q3zzWvR3lwnGX00ftTsb9dPh9aRZGEkkPsd+2waNSQG2
wxJFRIwS8DmyoVg3C1cqNt2fJ0Nnvw6WwWwYY3Lt5xwjNeGMxSSKYyfzerAoq+HS
mAEZR5HkEJXNXg8+g1lfq39p6SiBctGDzZ0Xo1rxqJB2rCGyqN/tPxSCIw6nrjCI
UF//RCIgmFSSSxd9cyADmYqPP0z/8Ru9GlP6JhDIsiapJC5SsUfUUeewFI3nAKW9
pDE8lU1/USQSwW2b2Ex3TTdVzBdESTFvY9t36p7/G+4Wk+QxnoEJqcfhRzQXAePi
34Krx2F17NWB2RAeXNBMgG1B8jzoecz9EV1a3YjnUJIhVatEEXx2uiQBCXaULbAJ
DvDAAX6e8TaBEZgHO8idNOOkZ12YaV6jE7KFfnNH0LEqEkTjW0crSciWHO68MxIx
v/8u0j45ui1NaChON+ig4+vF5H+5Wq1+2vfJcCoULgnfpe2Lt6XXkUp7GgP8XfG/
FKy4w9AlLawFc36sU1M+nqTp7Y7qF5PKkcqlEgJDZZ4aIsvTLeykaSA2RhxH4FFV
1W/ZDyoIzC+HgOf7qisyn6yihw9I2slLRv5sdDCzgxUcsRdYYOXb6RPg/hfm5F8i
dMIUBYvO1M4MEwlYjqZSUUwDvg0JDhql1iWZmkEHTjJt3vYMpa/mxtUeCT9Jqh0Z
Rngo6I08l0S1yIgahesqjCkRLUt/wEKSKYeZUaqwoo8GkJzfRZI+orx/Pw2/gJ5+
OsJyUzeuXKtvOFK7Jzzy984do2nn6DbERaiJ6XO4W9ogDVTpH8J82ZAGWb/ZMIok
bGdP0sAMbOxUObexIFaTe9J+kLuda39rudktePtSHOeTFZtNz5D0nZBl/T1/kve2
8vv1I7haddVpuFrHJd2e+PkT9kyAyxEihixV4M7J8tM2uq6o+YnRIaHfoaQct4zI
3fYVIrAG+meg0dBP1HLF+g/maK2dJYS3wk8aWq4RmMGV7IsH9hpvc2eJvXMCdESx
mShmUlLR4Fm1u7I5TzSywT6tcOtlHFQjx+EOGpemFuRZX4o7r16IaYOl9UTfEvyn
Dzv13eCnH64blGbdRKQaCqoVTR+LiOgYYzzcAjS/g1Q44QnWfPpnwXFkJR+p6XM2
So2qEhMsycu5i2y8vi6NUmPrrsbmOmopT0Lb6UPSqgKX9VlvWNpCwbSvBJ2D17B7
u9oLebQIQjSvYm4HntQ9nV/KPewo1nB5L5d97rb+B0Ch/BsMgGJEkPuyc1uCe8Fr
j9it5Hp+S9nzzUbnzfI43C9FjwdR8Y++bVLTA9f37IiTvJkjj1TBON3Ux+ar16iA
WCrANfvY5uejZ06zF9xc7b82ntxRYgdWfX8XSBqpYipeQTsGa50NZweLpRRzwGEG
jahtwlLre5MvLCgQUeV2bg==
`pragma protect end_protected
