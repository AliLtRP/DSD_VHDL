library verilog;
use verilog.vl_types.all;
entity or_4_vlg_vec_tst is
end or_4_vlg_vec_tst;
