// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pkmVV+StNl1bChtwUuzvFIkthvcoeB6Sf46nYQ52nu4jWQvHBkgkyiFX32VN9YUt
RDkALdZ88d2QMX6pTXRRewAQ6V9QTG/vzGkSonL1n2Y5C34hmC2yJ5OlEo7dgmja
SBmFYAi2KpA9BbOG+G3WC4pfewW9446j8J/aGWGwaTk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6432)
wnKA3QdgP19Ve2EAt2Oc1mvB3EHc1iwmVYV3GBcYLvTbbPwi9iz5hUDTV6y8X7uu
+0pngHb3x2LzxQKFUHZA6eJp9YYPz4ihbOCpXkbtet4l0ZaGLi83IX0QYAw1KY62
DGKYRWFUAJu/8AA8qqOStMIyhSyvctPD7RDvYcMhy/cRPDakT/FdbNy4z2fBndqd
sQ+YQXrjMT6XrrpgV4W+Mub47VpoEe4xjrm/Kap/Y3g/irBX1AfZ+91AQiypT5Py
hfPIc4EAgACtys/Ks3DCafzMdar9steRtyva12b1x4REN2LE/hUvsJZLuRfPVJty
vj02nFOwV6NPulfSp6A3Nq3buc3xC7rEgL80zD/hL74+d0d1wv8tHde/1RxluYVx
NQH3LvE6pTBFWGG49D/GzJliHOUy4EEsbBy31IYRj0XnkZwXNsRipdVBV5jbSLbd
R41TjQgeWbmkowBFRQ7e9ZN8jNk9jRAJ9lhWwb27TIidbyl3SMhVdxYW4/RUPN5e
Mv885aJK2b1k/HpwrXLcLDw1Rb7UjzY06qm4zEN8tP9kVEPD2L4A/CJRko05QqLX
quagWHRg7op4cB8PE/DgYxpu+x9lQREfXVfDcnw5R9xsQI0oNdCUj4sKSoUgtueo
Qm4JzVx4o6kFVLGakeYmphbIanMK7V9dKnNmrOow4AUz4ktSS1HH+edSt2UpHm3s
MLKB5oqzhnpPo56p1Q9AjEHLe+pO0cuGuh45zpNgI7HVQ0bm5AMLuQp3fODvQo1x
QMhNf6whzI20CNQNztpIMy+0OeSE9R9nhR8CTibZlOtfbqapjijX5BXc3DWmXHVP
4gp/g+OIgRWn1curOFP0rYOQlOrIiucFvhBowXBsNARKpFmOyyd3lHE0wN5bWw7W
Um6ZhzozR56YMWEkYCM7ik9Go+I/5oVOdLpA6qqn0z29XXqJXAyzLlNghDIrv1P5
mszj5x5CcsShovic4Y5xtDNQNCnFsvcXz2BtHtEgPxFaO/Rx+EEM71KKyW2oOcmg
yQC+6Oy/HJAxcUmI8gAUtYFXIiTxgbXd0C5ZX6OJNBUzvTOpxZtPAkDuvr8PzEV6
Lukxjgfvxk0/4GMSzEMW7BBURu2BSZa1UOzDUdSiQds6LsNKcU1NwnLpyPyE2giB
hzaE9oI7PrxSi5ujjMpPmqflwriwYv9Rpta9iv2uPYAHQv4cAgVl7lR1uO62fXNT
H+3ss0omzIe5cx8/8BCMNdwlj/Z0Jp9KNskDt2oSp0hTcMPmLoiuMmQEfGeabqUF
aQMSnWZkZsGJ8uGDT6IYQHNu3Hzu7ekhAyQfZO69peAd6bTQmjeCiCHWsCMcc5Ld
McZbZKKXgq89oNdP52TZrxHfV4yPGZyDN9SkKtF8H7HoQ2e/hJ3UrfIcl5XSEFBb
4HxPSMCjftvW+v2uZ9h/2/I+CTg44AyIieN9cB0Ugv04kBRBkUDfxe/UWnPYcI5f
wdnO/+RhUxaGoAEjLtfTBlVT9U8E/aLg6ElW4d1tJ2run3anJ3eHL9iNf8xQVtYT
pF7mTEG3gCnHtpJ1xJcHGG2nHlsAhfEWbGkr119sMQXbtPbcktZC04p20J61YL8M
qhWXCI5FKQYMKlquk32YL2eRd0+i0feMkKr/Ei0hDlr2gerCGwI461tLxNpWoS2b
hBH+fojl58JxSzLsjZHYSrj7X0DKZNXqzwdRILDB3gTxNqUVJZCAbHdDZfMtoXzM
l7jWWXfvPg0+01VoPNWD7XFA0eF0KbDgTLig+23UiTTR04TKJ3aaK8OQUmPmhip1
8wZ1Xkz11L1v2lKGFB4NF2C236KswR+SLXngZ7jEJtsXtjZL6UmiVMHnwVB4FddJ
HKDIAuzMxeKh4MFYFDjzzuh43kjtdx2UMBKtUyBluwGC6CZ3NNEUCe5pIw0y9QBx
1Ii+3v96G5mPJ4Bj4RD2x23Pnsxf2beM+1wzZpJaLjJipc6Tm+sOHzkOuO6s9BNa
XjXas9JP6jg3qWrrA4f+7I0hnm0ykyEC+rKcrd/9IJ3BCMMRhID/FPSVbeYrS4Mr
aVwLk6LIcnh/AKqpFHxdi2Sz0StU4+SA0i3OzhLtm+EsN5P45wtwZBUjVmWuK1Om
4O02lsp3y79nSGhzhEDe4sd9ZNSfKUJvePN4WSC8199Br4WFrRbHMtzbq3bjuzUB
j7yTRSI+UhV+sPryEPvrfzUSNS09o/rRUuX47iqP7j6tl0Ta8f74+OectsZwE1pV
Sfo0lkAoKPVOYYllAACU9GBdCksl+Y7faf7mX/HpXz2In4A3HkpnCQKsL2UAAMRU
GD3Laz8vFPeLKGNFg69w4S6TfamVQce29ze5uOWgPXiUw1054hziXWJWCF0ZHbbG
zykxKB+lkkJdIA597qUgLmVhld7qiGBY/AQvk7L4Q0IgKiUI8giIvK99GFCVCBj8
lyNl0EPNHTHYLm8y6ZRG7COKYSGFwJQ4dzBBQ52nW/6Cje5CmIR5DLWKqxQEaCId
04FstsTrPEa5LeLEjm1YewCzz1aCufRXXY2adivHam7hTlnAXehYyI9tnJhLdD8M
I2qPtJpYHnZD+7gkpaAASfCNa8258woJ0do3aNsk6ZPggwvvLeHWdFlY5Ux6OnfE
mTnX3ijzBPMGGoCoyHOaLXKsEmmgkg5qzeqUvDAVWqZuNZ4p5JV/+jbS8Krc76yo
Vl+GDTFOXx0wDY53K+QrvQR8PUYGiGa5W4noof+f0N3XUBsDJaSLQep4LcNRKSmj
NVcouj5sNGt/a9KSw6utnPzQ2Agnx56IuerkRyxyc9XgjB9pE5UplPM+xYSokKZN
Al8yIe98FXc+5mlXJbW0KktKKWMBuMHUqFV/WPD1NOeP1KZHLsIIUsLQk8JxNeUk
srxj5BA0QwY1LDmHklqsbirbInww69kYNW8Bt2fXofRz29VO6SoYT7+SLLGFt0vD
v60FZmPuVcwOX1UjkXSu9dqeGha1bNFSK10DRlKxEt9rl5/R1+zw7esBmJABAAAG
RcX0KJeww5zFik5ZN2cLWbETD3d92m2r77WMRgIiWuEzauUbB1jsOeGWBGLWnQ6B
TZwhe5lq6RLisWnJnx7WkwqjIyz1I2ZZuB891OFGyuLiu8XbF3e9E1oPQRf46yNd
zLn09JDC7FhHu2h/4lpM8gAbQzsMDdK/tAvsO2A/TJ6dp2g5rnxnO40XTyh1w3VC
QDBIZ0D2DYNAjHf24I1vjdQIMK9y6Vbw4qfGrQ7wtjj7OVW/sN7QsbZw8oRiMOPA
ypzZKFSIC+Ymic0WRqMcPy2HrKI3iY6asJLb7SOXYy1JhaHULTnxqq+BJEsd6aUp
8s25zCgEVaWJjbiW2Jtc8AwExAFiGe6R85UzkvwwPxoN4LL4ZUdGA9DRgf4oZyn/
PjNUlgvk6bJJ1t92vGGAwBP654RRRmwkR4NeFyfsjGik2ConznRy5PyL3psciJ5p
2fg9tq4Ph/opErKR1yjUmsDcfjHRVXXKcSNF2v3Bf6J+CrSNOVim1eEC8kgC77GY
JdHgDv4RVHFoMLkM7EY/1sDXpwE1ay2e2LYh5OMpqMyW2oCTW2zfqm8VegHH08Ui
r0RK2PpNm6z9bKL59ObMHgxvHEGoUC0Qr2jx51D7sfhNX3gvgwHykt99g3yklNmH
g5xKaajAPkBg8POL+35JIi0DoD7lDTYURuoH7He2KtYlOkMyuG2b+BRRQUkoBCBG
CB3DLY4xLICvGzOR+LRf+pFOzWOeEi4mjbCcZmhp3x/+wygkN8LXmXCbFkBZMIIW
cDWnrryxpAHxtEHyx6rnNnPL66XC3Pcegx2+r3k8Lbqi3OjIXUSgEodDbbMh9B3K
W+HZ5d6anXAyItvovaZIhWgPMA2g5+uTJz7NN+pzPa7cF61LclnaTIIsHHhZXSXo
zEzaKSEYOScLTlLsVmAHfl7Xc3CkTVfIR2ABHH2499FbOCV8vKhKB+HoFcAFjE/M
gvDqE4UCNFE1mYi8vUmjDXuDY0I+oFm2Xi3j8lyN/ulA9pa5w9+yb6ltf54pgbtP
9X/gI1HwNoomqcodBuxRrIOylb5VDSYl6sDuUt3GfR2rbq5M/GEssl90fX+GlB0p
VMy33p9gIJywdoxqKa2jlcReHA0nXnyxq8n8fclRgY5NzpDLrqeSU6weWkZAatNQ
4R58hK/YkW44CkyFVn2RkIaLbzUCYQKYzI0JOiPQrAApjoMQR94gRSsZ30tbeGlx
262yE96S9Ok7UQqu7ZPdahiIg8OHcYdaOrP/L6EH2X3l68ufyvufMSMcN1dgrAqX
v5MfMPDJVVAU2MAEixdf05snkLXL2CPLd9iyjjilBdsWWnJXy4qDxdviT1JpjluE
KBN9noZj+jgk37LTJMqSiwoZcrcqvRTerH4kNPN/y/k/55GEqpdBi2rlBNnLrWUr
fIQhM8Y6ifEd5vGmgXGUlSPlyQvO0EjsKllNa7C4yXabQ6FHkzSQAX0NWGkJcpXA
bJKjgnb90B8LbB9sRondqx+xgOhwiBd3cZUie6XMgqCFyPwf5YZhD09ycpWWakVq
+TRoVfreEJOntFeh8q6AGwOuZ1WWYoEu7UJXZwO8vouEwmF4reGP9PlO8L3MxVTz
+Cr8SyChXmkK6V3VxiFUANSAcidm9028cxKa+4DKZQuUecHIaFUGZlacAoGtdQ+9
wVVwFRC2lzriBSiJcxnx2eSxqvchjJ23F/RGFEDcXVFPsY2nM6bQ7mVOc5izUK8M
PpD81+JIxHcKgRAD3Agrpl7xTqI5n93yxIeUegaw+oVzWUZQAQBvAeJZz1GIQ7fv
qSPAGghedFXJYvgcYmMrlShUcbYPQ2ev7NrzzAzXo8XZ9fqxwIOagfi12wSn2hFg
Ct90+NmKI7nFm0YfZ3JgOJXse2QCsLP/QiOfXMMPH96tLbnbAWDEShP4I8hrOCFn
K224OSGfTC1PhUhQdhv8h8QTh2cFwWR/Wf2wkwjJZYlLGmlg/Ddfoe6ENWzOAQX0
lsI85yMx5+Vv2xZ6TyxbZhKIzNQklDEOedFuzZXflAGXvudC9nYs1RGv1N9FMrnB
RNfMVn5kN68w4C66OxQx+83UlYCjKMVUFWBvgo4tboQezQxwv9OnizDrwMDMY9Qz
LTIODOlqmI1PijCJDFKE6MyrC43sQ+MDfb/ntejeg9CLbrUb9SFrVMckHamOIK3/
Y2g6mIlatLJWj2APKSlKNLIoWi9eO3cesdjrxnFldxnVQ9X+dMNiAjDEnmqZ8F3S
RiOsLeDSdLGgRNrNUkbgB6JXcI3+UE6YxaRMjWlyKhGg9SEiFlG+k2rO0UnJ4YGN
AWRXT+sE7/yl2lTyC0GZgF09PhpmhtHPfoVv4abo3O0EYNV90Lfi/DAB8wqQbA5i
GYKIC2zbXuLlmYvNGnv2mSCQoMBNDQCdTO9dbC9dMU4aKGLZDL+un2+loyLxuuKv
s6IM5S+45zRfKpxdzYxy8+d/nbhBXgNnD45ZV0x+qtxXX8E4zA6L9jhHCasRNWbB
jSa0j9oNenebHXqmPUtmNXZ6d7MrAoTPcdp41VCUzPMscspWuDBZkI/3BLSdttDH
p/qVyHWPrl/cXYuC29XoBmTfiDc8Bv5VHj894CQfOyRZ1lDyqM8SxFpKHy68nzeX
QfjAkVeFlC1cE0S6IroeRS4A5OcS8dT6LDVpMMrVSDyMgNLdnenDUmSbYrG6NtWg
qz8mn2Qnwfr5ALCpyGjJYewRfBGzUPrdewt58QQsIiCNwuEdtxBGTsXwH1pqxnzJ
oNK3Phx+MkeFHdOOkPKDeZSplnhELdqCjAzDmR4Jga4rmgxe3BxsNmIgJCPuLOPL
YHGUAmDZWs1KqQpyU1APAOGD/eHJxDNXp5slqXjs77CH9YwA9DMd9khXLCs5cA3x
2PQC5KcVF0e3fzENgZmBZkJKQQObzu/58CyBvMxEvYhTm6+m+QA6RjIwtX5C1A/R
pGRKGm/Q78Jy01hVJr9AtupTBw2z06U2w6/EDR/s2C+sCrJArzUQlMtd5am5NvoW
940R9Pj+Thgp+JGna0M66ssrPRcIqD4rUpOgU+hQ1rCbItgW3unPNkGp5PNzWsFN
FATArAOSAqfve5ONIZlaAf2gcFMR1ovy7vUcOL5YTXiY7TGBu3mFxhSv3EHtV8Kk
m/nWYpSXHnkW9eEPLpKPyX/0FZtSiuPNZLPGCWBUCF79rPlR78+RogpV4DBenq4v
oAVdCsPGTm03UzsgrnSRrAoC8ZcdixnUy2g4F8S4CwSGLnnkerH63FsN7JLQxeHS
a2iAID7rlfw1TrOzaRG2HyoAWppkLWDWuVy3WjhEZNPqI3kMe3pmoya779WNScA5
dvkLazc8/eDCr7Lb4kq/bHjsfodLnSIZXhuSGWrnvJAIE2CIyDWi5qRP89qJSs/w
PLcFIDEQJFHnoIbQDdwMd7AZMSSdixGlhnVB0hnWYJip5ztma6mzjLHvZVdyKASH
HpBmH4U4BqSbdUFiwggwnNuhBkRnNrKSHw+wnJRK+dQUlPn3gl1+gxehHz78HcmK
ZRwxGs1V0j8Q0xUwj1fm7xzkI0rsOQPzWdGpfuFg2kUuekVmN6BS+tUeEb7m9iOZ
AGdyEErA1PT1gt/nP3SfaluRYczoM9sHysHpvsTkxuB/D9MIzGuajbKy2hoErQsF
jM7nBOG1zruUG+XZGsUHeMu3WxxTzC1oUDXoD2IxhQw4zSd5cJojyIoVJpZpLgr8
v/T+1n5u5sRWRvI78hNGmCxBweDQ+VUMoGLQxnDi59Zsb01vinjfx1TG4ZzKpLkr
eqbCAvEAVNPp/55VEODkrBn2mQFaEGh6YJWPSRbGJ3xuyRqt/s96tfkR382PT89b
A3ZpL79xSKz3ZJM28LJShBlRe6KKWmSrZFo4mD+QMl5V81culO+2r8TCzLL+1Xlz
sog92Z5XrGJ+SgtGSb3rhxjGCo0pao0oddaPTZDlk+t7vI3yIWNWyBiokMhBPfK6
kZ8ovsPCR4AcNbdNdV8sRxQaXj1A/eWcJUsEUE5vDCnzL18KbteLlv1+kOAo71jd
n/oUftpqRXvTDo3Eu5Xs7MO1k/Ds75/T+QoWHIfaq9EJn9GWA8X25Bf2GH30mELd
WtKaoFeqySiLvJjutuv/PEko9CjNPo7zwKPR0+mQOTgmyrZPdgKuLA3tCFox+wB4
bjWetEFdypYz4dcfRSJYWxyuXkTwcH/JLH5WfadNkslUAspO/vjQXBhSAG5Ni5t/
9G0n4Cg2w8/BtWrPVvhks98CZquOYOGBJkzVNd9ZZZrMgpI0pDng+cE0R6XTOFuM
/c37DUw1FtFZGH5OfkEuLICx68epajGG/waeUT3YvvOLFAMhBMTyHq4urE/37VlX
fZNtRXNGueLm1ke1Brfdm+rzd/0d1Age+G1DWEtJrvIOvxWfq7SLDOZDHQnzV1dc
+037BGz+xWJQkJjzNPt6c4tZbaWjWOGC0faY+bgYtgSZs4CkUr3eKLW4DoKQ2pAm
yrMCgtqDQlA0bD3mDleN37Kle9IqYZf2I9ZlkSWBZipWDTVkWn/yLs9+cORePiMe
5MO8U+JLJDGYLw1pztdfdFmN/gfOVias6TTKQ+wq0RhJfM+832YU4IQlCVnm+1Hb
EwTcv+3dY1zMIcmIAGm17Y/hN60uG+lUwBHAwSz3i/xaVK5auTODlDgOnEl/xl8V
oOZr/5VhNCWf/xxwx3IhiD3Fk/xAhRdhsTqfKQfrE8ekymDJt+kks1Y99GDQKZYS
MFG53/B1/UldohsoyN/hrprd+PGWtS1YZRN2ONzxAhhGODklDp5wQisLsbTpFJzB
cW/VztYnOH4vTxXS0HaiT9sUuqVolxLEqsN4Qm1DbNPe8o1V50jFyEkBH1vt+P/T
IqOsV0900LZX9nFAeVi9MHjd1nzgmtuBCLe1MHgucWAEUZjFA20wj3GFG72uegmu
sDhhz+OOkn0VKz/SXa3pLv+ekmZbINUsOIYHzYh/3pvBlLc7un+xr+edlmDlfDl2
Mq1zG9SbOrMfwGfziFTrGf9ExLVCgm6XeUK1MgHYkwEJC7Zcs6Q1H1owkVZvTGDq
YsXZ/Qd0EriQ4/BS5KGETaK8hx+OMnZzbhs6/wZfQYTUOMg877/7YpvhZRWu7ibE
nNcSESPKph3yHb4dQCB/vKD28XChYbkbJY69NT2OKyv9U5aIAIwtGavndm2bWplz
XcM8Q+XV8F8Jy337MIyU40Z0Prsud2zMG+NyoqZZIdvLhQa3M7x7I0/4i8h2jixc
iXEOog+Z6CXAO82AkM2v1AeY+QTwYFwYAkmCd3sWUNoxFU8i+oIxeId3/xUO3ZQl
6uQAD0iOq/UMco+zl833Hn7OcFhemaJWi1v1LFqSIWmCMMSf6ZOp++dhn1Ak8DpK
5PVupuqk6aM1S72yyCIAOfObfshP9I3x+f2+CGxVv81vXjmY5JnmmbQ5JvWt64Ap
uf9vNJAwVSDsOm+kiES/i99GfN8K5YaSPQzyxsD9bEDUJ78YJMXSKe7PtTl6mDb9
hB4Ry4sDKPnkXPvSK37eOlF4a9dd2n0HpDCb+ZHWTyrBKSpv5oTS3BSkp7LoxL/v
`pragma protect end_protected
