// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qhhQopZkrV2h9puegl3CfA4yGLNyQJ1jqQgJMAw728RBPXre7qBmus9O8//0SOew
mm7OVSf8SYViUTodIPBf59qgD1yDehgpWECztQXSGOKA4DReFHuX4e3eRaVDQGhi
5o6NVFakhZhKf5pu/M2uckBMNuhismGfMvTjUpIC1Qk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29056)
R3wsPmy1XkftS0CixCkNLYN/87xLrgHJURw9IhpCP0b3iyfWxhs4cFul6shZcKN/
deMy4Qk2GU0U1dFSj4Z2DUJdheRmjl/3Ms9eqhmLvj3FleE08UwbQle8/DGc6QpI
IeDLoEV2G1iNjv1RCPvJbsuwPUJq/r4EAyVUWUjxOF0sIu4BydvsOKNTDno3yeYz
Zeq5eubK6NCXL73l7nsk234jG6JBe2ZJcDe/UP7lHRLE7K9L3FnjR6iz8lSXvGNF
iQLEIkf1KF7XgR/nJGSisJWwMgdFVmXPIEVW40Ra694gTdcNs3Dpso50aiP3EReu
kMUmSfkIB51baD+AyGEAD+QKENBZV+ynj08BT+TKXi00IGwGgp219YmYADxEejHT
+gjxssUxUD8KM2rR0v+hV7R7LT4nHS3Nr8mIW3KyFWgyiFnTVeRp7pF1OjVWDoe/
XDyzTKOCADv9puL+46YiPi26g787xPxHDigskGyHqgLFfVsxWd82JvWteYjcQGqC
CriWzTCzsDAtrtqhS8ZzfCSTc8wsjY1QKKA903R26vmJNj8GdB2oz6q7nWOdWDCe
1aYZEon1tipFPsgyySoyV7WjUzzgvHEOmUQYRx56ZhLVEqZ/soDUqiUeJcqd3Ohf
wVNKgu9taLoc/69Vah0mD72mCajARI54oQZMxiE0WdM/P/Fa7TLAtMisvt9y13lk
qrEaIAWPi7jku4iq8x65hSdrGMzE8XdxHd3oPTrEJEd9h36b/6ljrRTGTIwfbH5o
ncET0QpUEYC5HKirXwnTA/nC2s+5oin2waynNQHaJaqJ9n00eTfUeYj+9zt+yf0J
OkYAIkRG6Z4Sww0S9SPtApT17v2PExZCYTDwlZOEScokMhv0EO2XEFnsmbE5tjiL
A7ooq3VV2ZK3lmEjcceSEDwjcwUc2+bA+ed9MPcK1sRjMmOTSndLi2AeJtWrQSYg
ZZ0yzyUgKR38pTgrhhw23DL6vozZ+V9hO9zTXkWE7wAxoWLq5RH6j29wqIRxoX9b
B/EOptZd7+WmwFpVap0qNYJ8kaA8X1hxmuKtXGartK/2arT65BkyAidlGpMPcuGb
N8kEwv8b20ePwsa3/crgcKP19QIPw4F2djCUUJtGpky/1vEdji9wmYYtToamyjdl
khYDUeDKzsbZCLan5PmhaeVH680vccy2CUYwP1Re+GPYN2bWBWibWIq/O0K9YbQd
rFSVtDRNBmLijSujYPZkDFLUG5nSsWMK2+3DtqJK55JQNI9xMlz47bieiltve74Y
Z8o9nqAEL1ASo1A/YRRMY+eGkvBr7QIicEImQcstfZoLsPmVl/Am+e/3cEQvt1sh
UV7BF4j14k5S95IOMWlRfeP/gkbjihib+3KVAmoiIN7BmNZdfqtwupQR+z7Iz/gg
By9QHbTHMBU1fSiqcb5dWs/beVEQ4LHPxU2pAsK74ub794IRZa/DQFMBA5c7qnFz
fnJfxvaT68ROzcypChfcRQH1TDs4ei3MhN4TPJPRKAupVKF5BX88iEOfuLx18a3b
TJjRZke0aqJX/w7lvbB2OTXyiQQxPAIpEx+4J+pCHPBZ91m6hDg0WM5vrH0MZMAe
wIj0y1HDRUZz8ubGSWC+OiAqvxy98V0+8vRbDVssExGuheQBn5iWGz64V6w+70+k
xV3HRKCSCqZ7Hc68RJ2UIzXoD92loXJOWb8GjoK59mlmPaLDOyNDIEPfZdRGhvP4
jpU/JR2/H13BM4Oo+p8raZLdRdXfIW9TaTMLeayDiGEVEisFu/EydMtKboQg/8cy
PflmPSmJnlRdOGOfZ2c+K9+2NF3pkkGyi7W2jKcTHcFuaIiR2gvrqpSPwNt2srMK
I+/d88UoHAc4wYJwbRu80OB7EqOgeP5aWlGnJlbldnOMnxDlh0+jSaniK4kheCFf
/Vaud43a137yOp/FBGa03TStTB3Nc2s+Ff8PQiZ+Rp9gH7jJg5O9TSQo4hPChoG4
3jHhIWEpKVHDvJmk3dgXf6PfpxzVzXIJh4Kp5vgo1AWHUPoK9ampLhJTnx2ev9SV
dNbu1N5M3AEe8okFpJwytR1kcnIEyFf9V7EgCb1M5couJinZ+6wo4eMuCfjXKlVX
Kd8YWq693PozH0exMk2BxLsylyts52Ld3ylvtLPijulQnNkg1Jz2bHf73uGihvSZ
OuTvCEZIKhxE9VVV7+VBaWQ8OSCJ+IYqgcA+GveOn1XQF6vpvQP6HIA30i1Y1tRQ
6nRe/cAD21tPDczi0zJz5WChIeLjxF8St9v9U4svuWA2Ru0XYE9k9FhBS8kQ1nj6
O1vH4rbdLCPmRr/BamFeDpBWpEwYk/MpfvvAaIDyaIbigOmGxS1FYRiHGrvQsKlv
/wskSV4E+M/OmPZ7nZkFRcFzszCZ9+GY+0lPZTprfuKbohy7dZhdkHoiwMo0cFSy
4XcCZPcpoDClsJgQ65BRk4j3QNe/toDrYccFLN7G+efV+tVxoPU7M3JY0MowUSm8
jYlAp863JfRXBhHn8K1Pi6+DY6HWRaONjRV9thLefTH9EkA4096M/BzAN4ecLceo
YJu2PZnE8M92qCuBeopUCaiYRQPru9qnNkIh2sKAEk9mkgE688Y5Z2Nmny15R2By
80EuuAS03rm6bibZN60b1+Pk5iDRutu9grNbnp2niTYsSrJETf6K4ZB7zmu8S29w
9GOHDEH4VixZfQIWdz8/VQsdebi5MQ/p+XqD9assbG3YRxvaWn9qISo00fbO3Mm3
ye0Dnc+1ajZQNQoc8jsx85TKfyY+atrsW8OpFXDHRnr+dxiGZISt6/k6mmnK/rcQ
7d1epiXMSRhTAO2lm+tzLfU/05T7J0JICoXKIXmyOpRa/xqmkplYIWFVL+2NP9hJ
mXEHBv2LD69cjatV2yOR/BMtQ8vrnW3CBRVGtl0pdsQNZJLl0pjO8yNq89DeLdBH
RpsXy8SfiCzp7A9kF3Rga8PVEOafjH8hfgV9s/t57M7RuTbcMs6QwPy42DbV/ifm
eodCafFBcOYSCg9ajw9+q2h3Gc2kIrbfoP3+dXrG4eNF+Xjv8/GEYk23UkAtVZad
Nt7/liSjxKxHJA3Y6wuhx3MRa3dMEoNjd+XHW+IauA+2FRtrfsQuqONi9DdrAopS
aU+CEWBHlJnPwM9JwpxWVcewWQvrEWzvnJujOE+RlzI77ro9mnbJUubbR8kVM+tj
2Q4A/diY6jvLrOPiyVlimYmwtu74pRvMBgGMnqeKUuJZWZnVzFPhisxTToNTnj+v
HB+bl6QjlEMeTHDmDT+AZmcU5gpuHHAWWTyFpgYH3EzrGl22WBO7VImFZOrRgsEl
9zE0a+Krx4ZIyzCEB+NVzzXSttpiUtvBx3c6b07Ec8axwLnwmXf5/I6WLBU+IFv7
5TrI2x8XcknvFXrCBeOnrtK7BKVZYwH6eYTcJpVQwpO3RI6tg2YNVNsfaqko+WNv
jtm5bI61u1LJcHPGeKeC6JfZylO47oSX7v2Jcn7CFZq+j2YEPqfPPGCKGyCADkRy
ngrDuLS0eWcQgLpZpsAWY/rTUYA3EOh88Wn+SiSW6WsDLAsE++AvnN59jV0e9tc0
pd+yup71luTxAkxZ2ySTu1GkWWcsJQ8EoHIwpZsqaybTfZ4f1I/kX/ufOVaDem7K
vE477yUzdhgO7rwOR+zYCJtAi/tKbxNBS8llMnDpT4FHma4dzboa22cp4lJV1v+/
apFdNpZAgHblWmQ7Xm9wYQzVeH6X23ZhmtAaW5gK75YKPN1gIXxfMN0mWX4aDb1K
vCAu393rYrBB6nGQeMI9YzZg6bLDY/3v0huHqxZYfxliRQhwaHp2XsJytDeW2qKf
F4qL32GvwyI2dq1E24yu+/seKYiTVvYqYbsw5OcclYosQAb1x2rqGmfMGXRoU8NL
ezc8f4P5aaZg+FU2fUcFd0L3Fe9eMahBXzbxqNhib3Ot5yydSgRGK4WWeBSL+7Mo
anF2V7p84+hAB8ExzhMEdY/lTbOljYZRp/+DeeIYibOSlhHTQSro4giJ6Xp5SteP
VVfyix6ZOSbj4hEAi8n3zwM07YI4zkxSJ37QKley5jIsLOXa/V38ojJNXAOL+ncf
THV/kRathzxazg2GyBWezNMdoHmJNtcyFFvWtHA9jO0EgHl9srTnxY6vNlR7FaOh
Iih9qGbwbBH6VjybFJNY0a33iShSb3bIE+16KmrF2MHJP4MinAgghUhRifCrcyUn
K4Uy9u1+WBCtwhR5diYCwR4qvECxby/x3KORLhS/noyraObGngrIe2RsliFLSwrJ
PKUPjkLx+GESbNKYQwEYG+cZL+5HLrgdbSnVPOQumlColhB2rzSz98H1SKHr49EF
IFkS2/2wamChPjp9onNkzIy48Px2DSvu9xUOXa3gMFPjGB6ekiV/ql3vCrNNKH65
M/7N7qQqWvkaDG+De7ja8TonRb0G70AP49uCYaIw6c3TjXJop2x7veCWYe5NiZHJ
jfSC1/CwdzCXRvpHpqjyNIJMA4/Lej4aoPw8lOqMlVdqz0/lovyWUT3p/TzCHdJi
DBZicJPXaKXfe2B5okYe6oCQjp3P61rqNxyGCybAGvUlYUrXtufw5Zs40Tk8j/8A
9KJiX1hU+6xTYl6NDmux3SHep/wKy2NHssEhtaCR92r5bXgZFCPxlLHbsRZbC7Fs
DqzMHPQC57w4OVV8AYxuKknbx7QSHxq9Z6ZZ3I7mwzWGQSuNxSKJTJLG7UREP7yB
3nYPpufXXesgV+eT227JoDfy+A/s8tAioezH3YXHlCLV6nAyAw+bLb2fAFXQp/Pp
WEQ11eOeQsaidrAEfiqlKdnq7cKKGqw9iP1+1aJAtOV4MRNVssF8XmUrAVocrGb4
g6Wt7OR0wxeTqjdtTact2fpnriTi+JNghPREqsNYPxumTxoyOaOyh/harJ2D59Jj
T9ELz2hdfrBjYYBKtzalGRS0rZAPi2qFaHk2BpxPxbIAWWuvO6HHiXMWW27beUjx
Or/Hs1JBcMlrGRVymLnc3gaPNde/q8pJZAuXGZf0gayGOaVlfI0tHPKw5fikaOxb
cbhSe7LQNByNPWobRXK6Lo53dSQLsVQ5bHvkNOVzYXFgulGFNuH++5R9lYOZTB3R
0s4QTcC/oyG1BmM4dAXh+p3Z0j+hQDk/4H+xeoaWZ0EkC2F9EskAIea1INBjLQUM
+w5CRoDWvC/zcXj7QESOBPlxm32deQYvNSJUe8du54aIpVUUwFiF2zY6LpqRQ5Yx
uEr1Kx8HC7AHsU8YaQ9IUVux2oYg/KJoSOc8bAMTNBPviWH3gO+y3fkKls3T9Qv8
VepdpmWvIs4+cf2Lr29x1a6kRan/qi+5uuWwIx+VgKXO028Sobb0YNW/tiYXe38M
3I2FPCxC8q+Ysn0bD3JRukmKOhUXp2W7sEIHo9sfkrfEQVw0KWbqNJNPBsrxCD6G
kb9/boPO4qmcpL4wMqGFVQqAQEugiWs+fKysjAza0o7lcXtTmU8w8yn1hmrG/QKA
Jhup/zTC8f0JhtHekXlmaaVznoH+MmUhs+k+G09BHqIZ9I1vToXJsFvqpRz1TCVp
iQOqxiuklevw34HNomaqZ56Wt2mc3aGMNOdtCrl8TPxpDOLCWYHbL9i4Z4lZtrBv
TarXmQx+rxx6oEpd/1Vga7gAsTl1yYrIcIddi6FsRs+OuYbI1floK6gb0cwjjqoz
u6LosfF+WvvQduA5dL12lWqvrKqbctd6avlpwcGLMF2jrXLGYHEmmXN6XMc6xwDC
IiAHM/kYluLZ2zStecF2KpoX7cYgQzv1WfCJYNwlO5Def08R/q0fyULgifWIDWht
l0kS+E2W5b8wqK6G/3Tbk7drLiydeWMn20Xp+R6cfzs27qrhYWgpnJ+MGbaUVlAC
WDIy21c+3992vTGyEp9vAuxUUy4UQNASkwvyT4H858UiW3HH+Sz10M4GV3g4Mqfy
G/0BkWoXX/oJ+G8Hl95rd+YYWVJUzgICsojQ+4St9Z+SfkEZK2Gb/2XYHuxdY/db
S4wx5Q0laA3uJ4HYGwaN/pQbAFetD++BH/t5iGJz36leEnYFzxgLnNbPLHDxNLkw
caYitpFlobwm+hDpEe6a5nE7LOdpk7EzelQiDdrP54aft8eRbkWq0lg8w3aAAhL/
mjUBY/w5hMvY0sc5VkIX85v6YkNTf3OgMAgo/iSoqP8JOB21p0h8JeAr+0ou1vME
yyPfF/bMNtOPWqMgM0fGnmqlZJN/l7Zpa4utoSUEgkvp+R0yf4Bg/GD1hv6SJKhO
LFIx6tqGnZA5UCQ/3AmHVYM9D3FqrdHwZUAwt3z5iEodmnsZ8dksC2UlVCO/mD3j
ZlT7Jse3j8xigzElEXqBcCSrSw9C0X2lmvDpu+QgYCrRC4i1meTZoJfcH6RqYemD
eeYUCbLgPYCavxwId6Uwc9Zum6/vWp5xtaclzH8iKRIJj9ZbPobcUpRg0GMdt/XK
ioU3B90ewOSPKEJuQqzXVI8FugiyCg0aDe6XmEQQeMM42MBrqv4Iq6FXs6ivvE+j
xGGpjznTR6TjZkKmPdDtSoa8xzmhj5bjDTIqeYMLhnM3WXyZBMFkdlyZPhP/wiPh
9oqwI3lAwH5+V1UfEJif6PJJy0icZzTRpkvYsj8dAHhfq8/0M4P8PzGyyYFno+hj
7eBE6aYPeosumeSq3+3OxXBIdQhfJfBn6IGMgdF4u7rckOVb/s3v0f92iwhLf8jp
QYJyLlqL/qRbuW+yq8u+dhFnp2rLIj/B6H0D6v6UHA7gMRkCIC/6SHc/CvNgas9C
bfRR5s/KRavlC2wYOcKoFbcQnlqaxAWQ8652HF68JOiTbFU/1qNawhDbDJlcq+5s
TLD4jwSC9ljjuDLIlN0RzrWFibUDMdyR7D7Xy4mzMQAxH6K1VopGSXBI4zO/7t0C
5+HbCc3HKhEFnmMUb53lHvMgYN1ESdPSSCkFnICpp3aRmOKONE4pYKlicDlQlGnS
wIXLkyQebQJz48sEUPWd6PEsqysId9uvkjQBPn698Tgf2e+l1RdPYYDOMowyeWqs
b3UHPc7O9BJl17534+gM5VeFiXjIVBdoM/L57qCyND8l8L9qWxP0LN16nenKXcp8
2yPnBmP5SxDfevY+QcXtN1dGLr9jc4b9swmI7yxZoyxBG+wz7yvQRrgAyjoqucbr
jNyJj/8f5XIeqIE5g6pjfeUdD9h+HFvYjuusiJkSAamBcgJZblJufy4t9H5Pi5iU
gscJoxJ+9rzw1i66eDx4KqYAZA5tgTJ7oOfbpqkIEuYe2Rq+vANWJqrp2sLKzig+
DY9qektBMW1osd9z54JvYnh0MwQdyBPt+ah54PgI2HyPBUA8euTPEPIc+yHcLgrq
7EU3n4xJjcitGSy4vnQHmXKPAxVEJ6jDGSSUkrob2jQRAzE2h7XlM5RDO5kIyrCe
m2gTxpPnhkR9H4hz38qmlvwUeUCXTuGnET0eAFPMfJMEFbC/ebp9A2fTny/lDMCZ
XtjArRtJq2MP8B2EhloqZMTHmsJcQwuvKPpKAAtOSl6OGKWrtiELqHRq4qlCluQu
gmbD8iCiFV/RgWamQ19EASW1smYMDWqvrqR20bnJTn6VPjhj/pDwPRNWPCMoD5u9
prLCg47PAnv960lKA266cgCl2go33ypgID8hr0CELOd/j59/6b18FzQM7vXU6TkR
VT1YVpUyz+2yigrCe/OhBal3lYmAvGie2jtg+wSmP9EY88hIpO8cG2FYULe2YY5X
chllalBO3OApianUYDVy7xPJgnBwBXTpqmaSW1w3pWnJjkylg/In7s++c13pc+as
zLdZlFPs6hctxBBlGLP6DrFWu1uKJkDYOrM7f++4AhONM1jqipc9xgbe+oerTR+t
zkv4ftRpDEkqIs25wrupbgtpZ3emg+0Hd+yLCLmPoFzrWcSx/s26jyPZHBQ25imu
0F+CZYtRwKXyC4M+kYE2pQ1FpcGre00+tRKxyW5bW8VW3R4CgIlyjwwBjb7gQEOn
G5PjwFMTQlVd0VQotAv7zdmYhAtkG84ipIEJehytK5gCglUUr8u+vxTeMPVFnnu0
wVihyav1QmChBJp4CJ6OZZTc7sLzERTDi2bfATTiIc1u2Ex9iKAdUnQAeO0nc5t9
p89bhiaXpNe6uY4akrpA7xy8MU6Qsvja4Con0gTB9kWflgMe7VyOlu8+xqsvowDS
TTQxIYRixop0jRy/MBw1n5bJgOHx6p/hZseYQZrwqkoG7RMiRYqwezwUB0A+JCbj
Ah9VY35XB7QcBJNaGevAOdORMZANxB4schyLtHIALMI5fGhruDiEySQTpfjr7hGw
5Kde3hirv9KNc+sxYV8hxLy23Ir9R08iYvVh75Z5D4ji9YblOpBCJQIE1wxTFwSF
N8/UKPX8xpdvneiAvKcw5LlnDkF44iKP0WD+IC2J1V/kLV2ZPHs6J+MIedQnKvV2
f1F0BVu6ix2eqGBJ/CyfwnVSRw6iisuZaKaypsjh8HafPF5l9/ewFFdJNTGMexLm
/zOcDVXc9n62aw4vC3G+nRLmW18fOXrF12dAquLloSUsA7brIL0zb6YSwZhzqpDz
eu2PI1YnO8Zbr2rdEui+a5YNBmN/AXN9q9+B8VnCKbQSyluLCAAQQzj7skhAISET
XFyGiSJ2tpllIInik+1aWS7ZnrCkpfHu7hsye/FZyW/Q1kRVFAmfdakuQVT3VDsZ
OHgbL9PXgO26LD/FyhZoaBLNmiZPkx2C+1TyRi71KhiZw2ajcrhV6wk+teHXiCRW
kb9rt/E6d09i8Xe6pHEiQqImrB2SOUbZfM2PSqy4lpAQ3d4lED6cTO7FZK7N+Loi
n35A5X7J6M7e6hJBpz8h37iXweHUcInBGZyLbZeNraQ2JacnyO5fXShStgxGERy7
2gDdfqP8Xmxgf2TnCFt9u9oGFnZek4YNYpliGYd3Cl4mWAwbfAUiQE+nLU7wcdJr
Yv/GNHWklt70J4H20TeBPFZ/iYRcCnPbKLcQkoaWqGVbolzYxw45/cUcrn4b4lsu
a7fhy2+f9PDeKDb37Tttl8QTvkveWoGl7fsqrBQlhW8zpsTmDpN9GzjfcbjC2SI+
LAF4Q2YD3FF5FxPPeTp7UnRclXeXuTAeG34X9+P2J646eJnUwrtlRbD65n1oX5pp
9Jqiqq40M3Ycyuss4XlNLJIEnAPPz61TGRHEPbvhr+n5DSrDva/RcBQkQ8KLUsSO
ASj3VRUC7xd163AoLr8afpsNwonmYW0OpgHxNZcscRFAFvO6FCEp8ljOd9bQAabZ
rBsxxcwszOEPPn9HTdcg5tw/g/bORMn9YeT5oEFB3fX8KMbDZXs5/K3yElXw60/f
/IKRtq8T/d24mg+EltUI1znPvx/poKknf1OAm6Pv0xCyB671QoyDwO+iGjPOMm9t
0yoAuN5S8tCMQeSYfB1fSS8Yjh8jSV5meDq4Ycdbdysbxb4AQH6KVaG+KPKkPFQe
qxa/89xZlqywbsNzaVZXf7Kgz9kD1bayKBV4O9VVnF0YkwyPeByahwEL7ZgGIBav
kcS8wjNIBYt4ec8bXTYzB4xN9DKHj71OBf18QF5DyxdKXrnepVeYc502yhKnSE15
fORoAcLmXGwyw0K5VCDDUxhCXsEJ29g1GPB3jTo1jILQFTaZsvVN4LL0NS0lxGch
uRpI3K1Fjkfm3bfEibfpvZ5vRA8/7jSMTSHgzCO4Z5/TaDiDz0GRVAmepM1vTIW5
RuyB5HX+Wl1SQcV/l+rbuuA1oEHxIBYvZEpOmLRqxTaIAwFpgA1T43ez2+kHX8PP
KTxkh+gtvdhioDeZfJfUsnegF0SF038SL/sWi8WrSNHnNn7EMmp6F55mvzwE+CA6
ciRLjuAFJGXvIE7zTiHAJw6cPG0gQZ1FdKVi1Df5PpWZNtKZePTOpJvmh6q2XWNE
2VEEufDPDUeHjWDoBxVhoMG4joCqXfEtXmUbzf/deaQ5+d4Lr3tEcTTfJNuHAZVz
b4KuKKkW4Jwt55Kw1h+WKyNVpX/Ist1OYMe+l6BQTIqK3yasQ5iND+nZ9MGaHhfM
E3+GeLmwfJjgjBLZ5L8vyFqjMOedLzxymkm/nj3tpzExQbjdfrFFQV9Q985A6r73
osOarnAej6gZYL6Q6sEWDoD5mjo8y9GzFBUO5jSSHoeydOQRJ984onmVD7gITLqc
mSR5xyFZ53nuWxNdRh7pVcU9vylRceNhuO+aEDciE3qmGP38Aa01hT4aKIP6pv4K
mvfNHBAl1xaFFymyx9I84IttR0ct0fZsbGHfzZ2hTJq5wob/UEbaF8nnAr5pkXvZ
+X2Rb6S1eV8fecfYXy2yU18irlrdFucDgKlQPQPFuLd1ZezbqW7QqaVPVt/bs3By
digxPEfLWwrCGLpFXdva81Ou0XISN5CBRy/6aXHAdPVLg4Va6t4qUsd+GaE2EsIf
A2TIrRhC58edhWusnafjQLVIQ2iur7g6CySErBQmC1vF5cE4pgLuvy70ziQGovv6
tEhTDZcgEndzYXeDF9PQqN8aBtR0oRu3dKvR5JGSjHPOAYhQnmFsKYKvPViMlhiI
fm0nxvoChYxdzf5+WiMEv4h21AuLvSSIMHljEKYp6aJm/TH8ZCe9X0YwhLvt5lkr
MCD+hrjzSRjL0TElHdSB1jqBdqoGNGn3TOfRbjJ+tI1EXVEawoU+VRV3KyhaB1Ue
EYUreNbUxzlkuH7p+6qtCe8oejBewSHZf0vlbDh4/adjuaWDr75XQ3HfZrEh4aEv
E7LmgxkPIWBBfWSxlBHChsM6aY7owM0hYc5LnSqzFameVz31XaEIvcSpKCGitAzw
l9Y63Axz0oVp5R/C8Urp1N1JFaZdmN0ii8gtpXiqe6nojLA+xxrkK28URHw3WOMk
C3PBCyJ2iRXyDKz/Dx86IIjTEUa5ItN+4OGsR9OWXaYc5hlBkyN7hqE6uXCZH38L
sF3j0SRZqyjlDgcpCDtdyVWV7fSDkgqrSlqxKRSOq7CNVk61LYCEI1ozYdAcygDy
gzSOSWu755SSXaidN9Ucfjl8QeoI88IJ3IvxCeHaZSFIxxOuJv0A+N5mUf4v2G2q
Pmu6RpiGHLTmGBO+xpUKMpSuBagPIWjL02r5QWDwVafpET5+M2y1FvNh/+OzJrxU
zjiOX89TDSZxEwPV1ZjdlMSKteh9lKbmKj9QIcODsv6XYnuYilqh3NtX0whCoC2u
qIebnvVmm/v7M1e0O68iUDTVnPLl7Y6/TQPvsYaBCNj3JZ4wOOXC3pkziRrA9l6Q
a/ZE1yCIlzXMxyKmaLpJZD8BHBD/jz3S+2cuXNdczMdjIY71WzvU69Qry2weeqd7
ewAu8xhI2aU1NCkLoNAMtOPu22+38XT3YzHho0QXPMZhNUVKR8eFJJHkymqWLmdt
XMCs6mLhMPD6z6+vcaA08F3IXiqvAjz1zKY+N6dVvrrcOrKFAGpBDUHpfhVlX/8Z
u+3Y80HnK4ofp5yoMCiY+xkJXOwV5JTARHuENGTEVWcTaEhL+Gv5Xzvum9a1ZX2F
lpIRHoiF4kTu6fGiy6VQlG4o6MsmRBEWfOlCZB5q4BnIWd04vLjE1QVD+obaerkX
iqiL+j0c+S7W2BKgwpUeLjqk43iYGv+8sTpKxCCMUdKI1tmQDdkEhlAUTSvEZ4N0
21UDiGRF5yVmVbQH+fs0swDfMRd2RiANN9xvb4YqVrNHf04FcqD4wVh10XJYgds9
vBvbJAOQUPVYE1Pz/cbjWWXzK94qiaNUzBfJCRhxKlpxYWWGQCs+F9MzM/WWvUip
zWWRCnvi3ClHskJdnwlce6z/SpnzVKInOUZcMs8d1q+l6nvGc2oM+vw4pqgiTuQs
Gv6kDJ0cm4T0Ix5Y+fvNoTidX61yYi09XJh3Vm08meGXmTMst6kqEAzkWhQfKcKZ
YZvOsbzd1V2hMzTXdUCUqvY0fIO5R8Xw2NjTYkdNCKgx/v5lpqRn+xQ8pGV6i/Oy
Z0RJx22AjOuI39EJnRszYG9a4Izg3XGk2grn3VrLJw/U0JOU3G6anS0GMvt1CSjI
LjmQ5uhRryKgdZmmVuf+HGfpHW2yp45vjPderna/jH2Qs6RrvorPXfemhfAfDGsT
iQ5VgeCnuMcfs5pyFz4C94dNy/Eg1c3wb4+1Q/Ws1FWXtUSkftHfTK8G/Ypzsrgk
YIWHAWho1m84zqfJuVWdIQJGRaGcyyiV1jA5XT+9cldrObekijQOGI4DSrEmjIgl
IX6/aG1hGdRvx/diqGK/UJ+Xk/j83TL2dlvSVip2RIv7noHjPN1I3oR6hmt6TH2Z
STxSfHOem0m6LP0MYwRsn04yXOizSP8hvW+cLEqA0FgjR2t1TAxOovBFcO9eZ3PO
KjOKm63gPwhH3CSwvNPAduYRTxkL47KP2GYWdg+2g9UYzcbOe0oKz0oLA3Km+sDy
pbukeI2Cl2oeFSIVtdoCLa28kXAe6tLl9WQC/EiROx7UUg4nMT6Z/2RIry/6CnJS
ohsau8kirZJFfo1JsZtffvAViHw5HxqS09ONK6eNMYLZf7n6GtrUJ4MC9ts9bfrX
caIkOUFICd2sQE078zmONIeIIzx04A91FrzW5N45lz3JBbMgCsw+cN9UGEPYe/vU
HQosQ7oLyubZ4pQNmji8G4awnb9efIQ1H8KPWCklQF27a30vom9p6WERawkW3MBa
pLYEKZNe1sYAoAJkVzR5/YekzrdWLge1p36dknLVnnKGPv0+H2Jb2MXUlETaHaAt
G0esDkQFnl9Pt6lOUqzrusCw5bPqCZjnl3VAtNnNBjS+r48rKBdEOvnQXfxUbdns
Cd9REOm5LkR6cfnd66MmZel3RQ3y3aNiQ1auqHPTKuxOh9sHX1VDRwHmvzwbYZhc
EyyUhN2yrA0I7H2lfjyb7zsNct/g8vN0E4HoJ9/4dW1nmnQyiN2bqJzYZWxNOZ/q
nF6xRV/kFELmg4DkJud2YoS2CP1mAvrtHK0+3VSRGOT+8vzfCCoTOYfzAbyyeGwD
6+eH5LZaC4kQNbsfbS7kNUnWQ6Rs+MoDjgrR+CzIIsoSPqLvVU4gQCzw387Jeftx
SVZzpzgOm74ogRRMPxAG/cD93gzohwoP5Q5Sxcgil6oOEcxmnHdLqjuNvfDTWIEI
DK98/iYvSu3sZGRmzvmKG+GDazrSyVFYtovONxGMC3NL8AiUolrvAJqkUgC0yJxj
GBMx5+aPYNIYJJC9j6neq5QdJzOjW6tjoYMo6K4vL2ykEHN7zYm5zEeSl+6yaI2X
25VoTEZoGVa6OPF/NzMjOJAUKsk781XdLDGyoK7x+6HCg0+jxaD5Y9floU1sI0LN
pLIiihMJAkFOQhYF7d6UYVxRJG+3ZfuMIAHRxdtr0KLpdF8OLosAfkYb99l4sSVl
Kf9BKPGOQKEkjDlwD+jbql0QEHbYlqcAkYMFsjH9l/ZtVH8543o6VpFjHlg/BSDK
7ncW5jCj5m4ex9QlKYlJjz558GGuqogpj4BZZkJzchTW0gVF5SsR3t5Wkgg224Aw
CrzbuF5lw/KoQ/weEZszrUuKEKun2FgOU7RgfSrFqERNjTvwX8+6PG2DceaxQwMp
pvfWAZ3ULDobpScJzqVdgTYOyf1Lug2Y4cFxxMXv5lWtDEYqIt4oV71XFNRPmGbl
+SkqzfOiDxrr1fR0ABQqrg8bnrJX8Bueq0IKF5rMt2jZC6iVRn3baLh2l2H0Bv8n
ctkvFYGOo3jADJyRvv4HRwLKSgv+/WNv8Q3gcWmPGviodZRqvwfVX0kdw2nm7N2J
nW44jexst365bvLG4GIcQGlQ0BdW3RerawQ0etxzrHV/2z/p9JZjWddv/wqcFtNe
1TKJ4GDbSrtTS/MQr8E6JtHiGNb9e79Ot2IJIgfPh3aBzbpVZ9qROaJxKDrLWhf2
0mDPQ005cMISf465IxF/frD9K/mu9Nsy6hz54WQu+e1JEcMnphHI45G2jpxl0CYG
5Ka0Dp69lsWKJGmzDZY6/jc1bUJhJzgthcU+R71BfKBAnsjb930kSgWOFZQucP16
tcKFPunaG2rw5sAoHtnmr4v8f3rMkPOqe/3+9ey9U8CqOFecQFzPjRwCeJYdcFLk
J4N9LFz5DioVohIXcgEfKHrK6jq3gx2nGJf6YYHIR7/A9ClqK1uCvvoT1OU/x2CU
mPrWUDzHwah2Lxu22AAONJT122WgYg+iVwRJxaaXpZvCBGRDNO6eyTXXFjtSK8M7
bKwd9/SLfZf5WZluRB4QNTZLgZro7Z0i+DdF3g7VhkTI3f/mcG4NK6VbLy0wL4Ks
KxhzqdOSJS3oBuBvS3LhmP7JRaTnTwoVdrv4uOAGJM/4pvv+W5wb3amhKcGvwSti
saLo8B0HCEsJsv5k8gEFkE1dIm7dmf9mfe+wk9M5yvFyH9T3FkSdpjF/F7eAMfB+
0lQpj5sbOdVaFHuqqsTsBgIKDvO4gKh9KoYdmZFbxFR46ojK/nt6U1aBksy1KJXO
MtvOSEOrTutHwleA7IAqNXBw2flLEhKbAYNFprkKMI2bazdfp9VQD5Y4afnUkzzb
gG2H/jCJXab30cUF4qH/Yn6HDYn+U7hFLHOuYcKSZXpt+Opq7Sh2UJVfKI5ym5kn
1P4pfMR/ni6GwS2+UNfEnmEstZ+G7BwQN2cKPkyBngnQOkXs8dqcnA15bdj8ghBT
5W/wtkl4IaiZ2S54pRWncE1fb2kD4944oiPzXaw3IrEuR7KlecWNq/CyH1LQpvx3
byt28ZpbVi7r05yvMCj4s1H8huo2bFJqigLI8hNSy/lcDF6GGgJJg6CL56F9QkKY
/AKvyZOjzx894HR2l6VuFQBvDQJQDOnrDvrVazMUpjxqrRwZVJGQc9RwIbml48AJ
3oTeePfaGuXt4gy+PmyI0OvVdwUd/En8oARJj2oxNqlxQ+KURNY3utZVK3WfpJt1
0VcNmgnverw0CRd/a80zSKLXXJBmJ182bBL1LvfVhgI8B6alZAWyWWwAD/PpPujb
39QT7j+IFHQ+DY7iVES3qPh1E0KeFRevmpm3rKTjz10K6SNZEOjJjM/eX4/xr1wY
TkU64FC3OIWmPtBwQ0e/UaKN8nvNz+CIqlnV6k/87zrqk2xNuz/KmJ6mSlgp1s2k
j7Myhghxvdc+jNYuUwf/R1Ptjd13+9KylkpXXJh8h3JDnwfQeg3BjSkyvWMap+rO
riVQ0G34v8O84ask1MUz2NX72DJnxl7ulCsFAODOJJSgE/HG/Kl8b9us5DVXLDfx
nBkXhdS5wvFyfykktTPoAvV9OP2K/lblP8FW+vltCE2dOBXozJEcNoSdkkjubkUl
3Vzi/WqvhxSxPJSykQBi8QBln+rQJggWpk1+JRAEyTqnnADRPrim+hYas5aw+w8L
xmVC/JtO8eIwAzJsunMTpyITV0C4Wj4S9zk/mMnHGuG5xefgr9zvEUu86eauqaAW
b7Pw9BK3PcLIdX4v0348MVEcRc3srV6PU47K1AJ1EnV838TZnyWpsJCNVoFw7tAN
L16plYpnnUFo/bGC5drawEFZ4RgvXeKlGn6IW6QGb2QCmeNsphjAVnkLYPKj84dF
q/0LxdS/cTkxbDXZWDA6xqTSA3SZfKkvLNFjhZ1GsU4hxVswNA58t0Wyk2V1dAvu
2ZKSqt7RK/a9yogUsYzYr1+DfQiMcpre0qWozidsfTZpKc6OIEEHUL3EjnJfFy1V
hg7fMHz426gkYsipZahK3bXZSo4OzN3LEF93gXYgqZNscjE6l0VRS8XLFfRbtifa
+WEODFiRQLZO5xUKjnOcedhNl6JwtQWwtBv+VN13bBO0sHTW0JWz3lUtfV+mIFRK
rhtM1bn3mFWY3W0lDf/qMW3x83x4gX+Z797C5JoYEKxU8a4GyoivAkuDrV19DQe4
qNzHQ3EqX3Cl2bmaU20LIOrH3swdlZg9h9f2jg/fexfbD/RHkURZdy+OgyJ7aeyp
s0bsOqfW7mnvkMp+W6tDilb4eg4asKKiU4byf87Dnh/MDNDKd8LoLaZqAZ3KYT/n
TkgXsTh1u/hLsaF74YaWYA17H5nGzojL+pUn3OalwV7J+ODpxZHiyFfzlzMviAFb
aqoKKzjYVCgPRHRbOmi7P0PrqWyNTRgQ15BLukbi80AvsCSFmj36bvQy6ncZal88
VwKID/x7lwVm/gkwv2Wmr7lzp1ze8n+XRsGf+jDkC6AJBrZtWb6bXjoZyaN5KX7c
4n5USe4MewnlBFpRtAwATMCl922kPWqRScLi6N2Exe3bOuq0OxXK4G1kdEYglgaQ
sOgAMSca/qr57GDxbJon7QKElZ04vLoVSpJrqgKrdU19bgsOgfGaR4yr6w5h7ACP
ISaZ7E9gyYQiXsbibT/1+/UNY10fM4DUfA0FYv5Beyv6KiycNvPiJgmqv5anSEZD
MrVPvj9lf02qcbfNDZo2jaNtOW1qqwatHnEErkEokv0WEjJ698Qn/saB2L4Cg8mc
TAGRHOHDbGCmqTYEtaitQyMavotTy93HvIeg+sE9Eroad9rYfZ3T+JhEHsz6m6PN
0AjyVzurKsQRvp5yFxvZ232dZ/8GiS7haOwaUIvKTwtuQcmJA4lYTyqlELn5PIm+
X0GYVnuYDH+hdVyCeaRpVOnqBOMuSOLgeSkxkni7G07VrT2pugdX0OXohrVduexn
XAV1RcC25RasNtmWf0JgiIWdXO1VrE7uccwDpyVGDCWbq8ji9ZVMjK6ktZLhE72E
ZTdiXUXN65LxJ1XXpuk95Jp4fNiZ8iq9uNBy42fc06YM27Wyd0tEfmzPo+eoPrtl
jd/ykynNQwnClmOkyu1ZpyhsVCfF/LU6xpfxfGyaZ9IzB+MV+QETO6wOt3cfSEWh
CRi8yI+oew1V0SRyQY998M/8p7xe+yVnJUeBo7G6oRg6+oArOGvcsx+HvZ4Eg3Ot
2N4kzLWvUTranOAIQD/0+i0wZopnPxfgCDL276EOc3Ll1OzUIgeumbMlYwDOxo/z
DLdGCWU36Onc7P8GpUkLYissh/R1IaRwEC+OTasD+7b9ckWnsmHclm6lrd+I+TIn
Zc6cS7bX4MzgttclIl5VvAOJBsaCBjPQZ1b5wGlBnp+C3nY7oHq95iPwgzoKEMn/
B0fs+664D3VcDFd11LJ87HmxwI8AiF+TugUfx+IjwoJOTABUAjKS6hEijmIMVgFy
0bTb/Ds4vCY9DC4cvfShwv8xIYXpeUN9pLqA+Hg00TGzu9e7BvQ8Vp2n444qqc/j
Z+kabBCesUzYGmooqHrZGPhKs4ZpMWs/4pFAmhk5IbF/gP08Yr54qv8gZa3vPS7Y
KwfZvVOa4aClMPwDHS6Q06QI4RjIYcdXB81f9djLAc6ghgsNkfJ9Ren0Hoz9ou6J
9t+AnKIGopqmeLQ0PGxdOnbq1PxgGySpHQXG7BdkLc3a0cxa25Elshn6riZHyhv9
GhPe+RfgZMHbHlYnoTqa8+rn1AtzZ5W9aL16gNYLpMRb8OP9njnqzfZmAXmZtnqT
mAGpakIe4qrS0qUcqpv5rvNGO8/NNkZ3NXhxVn4iM8L5JdSJPBQ6XLBuONCt/6LT
Mc3tSC6+VavVLmSFzPD0GXsB5SBCZJ8o/LbdcbX1BvLxrPljUMTARcoVlEnp/+3T
MEjDdLKHt4DCy++hBHDXEuRUJnHb9UWY3dYT85MMprSZxetV8syNwJ7N0ndi01Oi
nluqgYvMmcNAH5LsSJJpQkHnsyMok2LODlRiq6nV7F60ej9Z2458KvhjpX4Du/uQ
jyWa7dtMSCzcwbwPQlwhr5HVo15WTjFLjb8iGJYrrNWVU1Bum1fKjE8krzsMHvZ8
1kRMCWymu7nfRJclqcYfq2Z5wo3NiHdgOqbeFXwq3w3jJKj9ShqhrWqTmtj5xPbM
CtAh9LIMAXPAnitVqSQC+TmLpW4sFXJORaIqQ0JN9v80+aVKoXSeYz7COZaweqWc
4wzlkEnLFw1rx46hDGhqjfWI8IYMoyxVpD2FJnypqLo4xZpvayrTNNbjtaB154GG
na9dXFw/DSqYQrxZC9tCgG3mwTcotj4zz8ah+wj3oJXywQLhTtcfqoXLcZymusVf
iW4huCNXNv4AtUSvlAGhVhfZ099v4ZXepPKLIyA2o82FEEXulz9nkz6rUPhUlJNi
3DbYmTMmIfZNLtv94WY961trDmn7BFSgjMENuem2M8md1LZnUz/dDhplVfOK1Oxe
X8HH4IPBJnAboO6CM786Zw1iSGzsDMkjj8cplmKNXpa4LVIktePJ4hjFjJJHxMed
OaLFTeuYXc6vLzwTZJHydj7j2fDqh/PzYzVMT2YBIGL5rnDT0gWNxH+tyF3fsfcA
ka0y9WHPQC3+8G4Jq9eHi5Ab/W7oJoIAESQE4EXka53uT382ApN2hbqTRZDIF/2K
L3Y966RDTUiIYUwc+XIivBAtHb0r0pzkazSQh0LbZiP1fIGsVFhUAHj7KePYC0gd
wMqNjb4AJiacHgA+YmawcHMeVOEBlCPMiHQL3kFwT7s+EaqwbQ13Gn3MNsBRIDK9
jQYFit1xQIPXAiOGcGQIvvW1SqSLE71PGEYvuIZ6HXf9we8nopEgSMHaHbWTjBwp
EKiySHVFsgs90wp+nv4V0yGnse7Cvmctgo4Sz9Px/OCvB2F5aCFzxPA0M2Yi9rVE
yEiE/xNBk/c4X20iO/zpWOwnGSgu408XfrvK3mNqh2ETrTcLhc07WAZNTOQI7e/V
yrt6YHFPaM67MzacPpYqZ9hs16Eljf3M2KMnQAxD1Csa16osX8Umo9cr5PLrlGb1
ix5w2ZL4Jbod7I/UQaLO0jQItepkwDsk6kdGyqQga55js/qJ06AgFTyUljjRyHOD
YhVt+h0+K1D7c0L/IZJrc4suxada3+/16Jk/RWJkAxrY8SNhf+LCx/OLWsKMVztY
fwv0cRj++E4MCLiVsPDoKw3pr9V0u3TInR7fWUc0fw7iXhIbJO4rMH2r9+6zTVs5
b1x1zXM65AZatvCpt6GxA3FXJA1JauiV/igsw73b+Tq03kO9yr4z90xb4p/zC6Rf
RxPJpXb1hoZgefjTEGfTCf2Mfd4JTAgP3tAmgtLgyU3ZaxW24DXkI8saBIA8M26i
LTi5+cm9IAF+oxQnUndRhjrVuYvkkJdN7NGimxQT2zxj22czhecT4P+ZN6CccNVN
WQvem+dnO+RcKPEowDDHjNl72GJ+L/u6KogoW9kv0tYxCTYnTbME2pDozuQtNbrA
rMLqocdhYR1CxokShpwTEw2T3hzLdNykMOOJGeENqF4uBfAkNZcna7+f4DaL1SNK
xcK6rGp8G65Ujkeel5N5ro8ihEKNaDGeogtCa1xGs/FFPxpQu8GhwMU1q6wFSNVx
dY+mdkfzFOfzOcKaiCkdNKmEdnQG49JFBmXa4jw7Mm9bv0R2UF2H3/XzeabxhsTn
ai0xzwjUP4WdwybZsz7OipEV5k9nCN8sYLZm2a81fGmhz4WclwtB9H6NoNErXpQQ
0yvGrMtbcaaNQwg/pbBaTl97De2NgcQSp8zYbtCPaDXFugK1YpMsjoKf+STv8GbZ
12j5yfi9ET7934gwfdWYeve5ijDHsQD9GF0jir/2A8Hl/fCnm581mNS0UNSw7WtU
9jsPaYZLpLVSvZUfwO6GD8pKObPR97N/+WQ0oSHAgASUIkYcwALyK+lyRkj6gBxV
MlJsoPurdEW1+FXIFrZLYMvvvRVHjR0UxS0uLtpvatqj1fB+cyZLObnsM0uvLW/u
yEqYBkcZ0Tjh/VqHAQK2AmzBso9Hnbn1zUINIV8IUJBrAG2K6BBd0og4t1IMsEph
lNvVc24exq/Rr8261QU443DcRqEVFxPLIswPZi2YeDeSzetVPPMkhohszwdTGnFO
0O5OJRMMbYzOp5FLQiw6W4J4FCSjcfv91c7z+bs7Ke1xLJKFTbV+ml9nYfuiHIyX
zLO0O0b3n1GAbYTwKpLExMdOmN9KN/2DMdZEg+jSBkQuy514F2+PGfII6g5krEn7
qEpiXd+eXIrVZiegh4PdS9Ej/qv2BTli+21pE0GcnzLRt12NA0JZA9YLvh0fXGg0
nTh4Y8hBmRsis+ocnmkQSyE0bZBOiv3AJ3Vq1Ap3E9sLwyj0ejN4XbBmewXkajSb
CfH/d1INAFUHe1CP11+6ErCK/29DOe6nncMYAN2XRMoNetsSyPyfdiCqTjFx07o/
2TA4p3d26nTM1qlDJHvXVDOp6eaUIfyHUJAFi1xY31Kv4U5MlhDt9PjqTM5xJBzx
uR1nWYOo14LLGF2DDv6ST1PUpbjOJ9P7iRwoc3YOxK4sVo7PEHRxj+pZD6dlkHxV
MbuIT8+zbHrygLLFW77FNiLBL3aqci6O+T6tAZ9zxrrqBj4ALr1Qqpfrc/qr8dOP
oBCXDUzFfPN7XEV6r5o89hR6gc7Jws5725yeoaw9nYmJtudTQmNaj5i/dL9rF7f7
Y/M5xg0ikCMd3hl6Op6aR4R6Os7OwBk91aOA7HxfVslhS8Qs07q1ac5PD/fZuxcF
vZcOUHNBqZ6/Ew+qW3W6xTyIjxZU9VBNKR8NnXz7JbBeM6snd3KAsEda1NHvLB59
f+8DwcbhaW6qY7vVSGmmsy5REqHnhD00N7Mea/LIQrArlIiAKfVwIwryD7nP9o0r
LgXuapADF1u9fTX1QNYoRkV/4PwrWLfhSQB24z4yDxpvxMbTixXqjZUUnfNilf1v
0HXrLjiE8OhLGZUTrJqpiO2RQIrq6qBaIW11T7yGQyDeBq9hxXNf7rQfU9yXLz5E
SyMMhQvH4nTx2jaZl6i84fomAXZ3irh5YXkAvZpu+hnRHaqe6lJDxfpkAjN5XqWc
7OzOuh5Pmgp0KHBtkIIkBG+GflhJYK/lm+QDHe9tuSdr4SfWk5payywawEUwdaDs
ggRhCMWeKOxzgDBDkh129iHZxpzAY/NyMJIBWyAOeNX5uKDLEI26XKRY6Yk8Oiyw
ER3GyCuezUCjOi1bH00CXRGj/sKW7QHGA/ThDW6y4/X/ouDebpRUOyyozhALiOZc
sDuQdabFxNWNV8efRGKegBevzoovbFO4DdV+gLVVJxTNQF0VG2AjKGa4Naj7yvjc
YwnJm18i1jodWjLRPkvsGWESTeUTemzgYXJL+B3Qfu9p7whs1uE9BcmBVuCFEYcQ
k0OD0lH6HMfXpOLGFdpKa56vGg+rcTZt5JCrG/7fJzlMvEbGEcuEqQ69wn1BiEpE
saV67FCVk5sF+YDRwmPDrTDMtsnhhyX2MHsNBJZ8JSp994sXgp+4G5Z94fKxCNk6
nIOzJdCWrW/cePR1JQctuMv63NOAF9nnHXGR29e1ttVF+gchSFHCD3U4D7/Qi3Mh
pBg1JEXu05145VBylY/xE7rfpWd4JM4ALmfFmIgitO4QpDvjPd6EN3Uon8OP1xAi
ak/KdVjRr39RLkI+k6YMeAjl21DbpaKMEKkVcJp/X8I/OETdtuhh8G4mOq/n0myV
vtUZDPiRmFYKc/lsnxR4PsZof54BJedpHzYSO2gBWmsFHovIs1vO0fNF76apuXny
GcgmSoz6x+7k4vqenkUiL2E7UpUmiZMfy6SwcDDJbj8R65dKEnMAMjbOuvZifWwg
q4z4azNZj4wf+co+lRYJ9EQECkAYgwlK0PQA7H4hbSEoEN7WzW9ZMbAUoY7b5IoS
sBSA6czOEz4nVP9lMAGJg7VZlGOTWrI5HgVfVciqdxqMcpnRX0vK9B+VZ0xab972
Cme23YzSHixlM2e92ty3H2l1b5pQuN2XFvadBJ3mH5+T2HOXWEvIo1a3Oo+NGZ26
8ubETIcyAk5Px66rCM1yhGom3GPclA/tOHGOLScZymgdxu+BsfZCg4T902zEDfq8
zACyAuuLqIQDe+in3C7lNsT89iJ+wSyeSwwPOFVK/fc3wNW1Oxf3BvNf1eCBwmsP
dAs/12WCEjiihHdHahsQ9T3R5WnYpXfhGcWocVYUGGBeSUPyn6t+i5WnikpTIEAq
MabgGtu/YRQE8MPmfxU1SlbCzpE5QENmlmMawDYeGrv8TD8KCx+JmdMSa+MeXj1E
lpOmXpTVB6c2iytkzyRZwp6OI2Lgk1StH5sbSTDR2SzdHMZ4lyfc1HqyidCu3iAH
kKYbbHKasDn2+zP2q8jLaB8GFMA2mstWR5j9D1cbMM8X1wCPHZFVycgnaCQ19+j0
GHdWgQ9Gf3/tl6YE2QAWO1DO9zZf6SdDSSToU0cKpLPdeqIB3WcTEg7O07Vaib97
7IC/+RTPR0x/8XYUT4eOXwmN5SyR0Z2+ZBiv2swQHwrHVclpd0RZZaZGNj49uV1K
iLYQ2yFzc1XJfTwPTqy8GeJZVo98UZnWMlC5vq3Kf5XF12YQDp6vTtSHxDJ+h7pD
1hs6MxHuwALKl9ci+3CooJKwgAz+V3+PgR55bz9ChOah5WOtGRBeXScZa1JEygtl
uuQ8sFdV4x5oqN5K4y1SH59YGyKNl1kOr9n1BQW/nc+v2Zr/75zeLKAPcO23y3bR
TlDucZ04xFHJ0IQlhzozgWdpk7fAaOoSwvI/anMVlTvbxkiQlyfEJrbTIKUP6KzG
lcqIytRIt++7HVbT0h4sRyGdgOcbPc+PRE9iQgDGswODPh17nQslCwvijQwocGcS
hBJMJ71js4JBYSpeh8dIKYiiBdx338tVVhaWrO8nGXqDrWOCPMyFnGrUGCIsVoFe
L9KxUKuL7aeXcQUMM/PR6ZIbW+DZIRPZdEy4UahY5zEbn+PGgWeIT5I3AjUAFQnV
SDhAenEvrBeZmQ+d3G8c5s+hOm4z8jvVrMQOu68dOZOgfuUoRFlcXXKRITK9w6b4
TTmHFsz+Yhb5vkTltvWw7p1+DFHcNH7GVcWA2D+9K5us1HLyKl8Cy/RLfVSFTqHe
HZ6q6OMmQavhIWuR0EfmrckuNc/neD7vluYV010bCtOvE3j6aJfC7mjg+aISDQOM
F+VZ1ioQ/RBHl9IJARiMoCf3fzcIOE+qwfB+XcegUS5vZb7VJ5EtB7VVGkDTlgMa
JxKXC6DXqGKl66G2GkRwrRcNW4rYmF/ClvD0RdbDDOZDsHxSmxGBGVo/9OXoBIsM
x1S0+VskfLf85y7U8/Jc03ZA67DP4uMLxCXJiu770viKyYA2uy4mYlv63QxeOpzt
WlNVB30p0rI5AEUxO3l6UfSt2f/t0sC72Ium54MYgRwRFg7yimehtIbhfanMM1Vr
je3uUtFSQSiI77e2qDcEct0ek3kvpM96GOsoLllzjNzZ/VEj1v7sZF3+SeaZ4StV
ung6J/kadvoxcUlGwp/QyNpSvQDxgbG5UZaFLqlNuxcyysXJAjc1/GRQG5UvryCS
yDMHpAKkj4xIcR1GXcunERuVdWjjBo3kH7qvoycXlQK7pQcCMdT5x1yEm62gnQjI
kf08QzBAsaL3FcjZOnvnKWzJJNR6eYZcSbvFJCjrJbj71ovUVkbjSgJl8X5DcjsZ
HW8CgPDZ86masIJD7OTNHs8A0LPJ3/1mNXlJWsSW6j2ySUzzTSRJ/aHGyWdsccv6
zoKzFUglc5upMFcnKQm434j2stRSJj4HsL7geadGJquLFI8bQWT0uexBSX+20dya
UNmV3Q7iAfmto5RJILKq8e3waYw5Lt/KG+KdkuAv1S8qQRu9tfG6EKediWOvAHbZ
wK9fVnn/hcuFwk3JdGKMEZQJRZd7G32+ZLAfw7thOAYzDtgJV1JJN/Jav6pXW3zV
N9+fDOxXp0sN8K3KOiD9/wDzwisFTODQ08wnP3lTgpq7H23b0OOs22L38RZvhLnd
bqe2NW/3IJCftIF0VEb9ymJi+A52Gj7hTG4RmmNDbZ2GMzMz3mFc7nHI2PuJrmZY
DidO3ZPxYN0oBH+jbfST8vI8k8mvA+yBB7QYbUTZg0IvSZJWGNYghy2B9KyR13nb
bFAYcL0hGF4jZbsvEaiRaF4YaaEHjM1s6BwIDyhQNu4PgGPyA0KvS5DHjgvHvScq
SG5M3/gXhTfowQori2RLqiD7M9jcVcvnrl5vfNWVdelBVkLAXzyGnP8Umyn0nGha
tPrq/5zFZo/rBP0MFs9DP9GVyFMqiYfbDncr/+85Qo4QC3vjFiw4DX1C4w9ikdOS
yRazY4AueFU1j+062ijGQ+k+4Kct4CAZ2Ln8KDBlDwbJCBT66fPMoEg3s3e+FzXQ
A/eshzgsU9dXBi2mJ878lXRQI5YyWiLrnHmamtqMVoPfcK3112NeDtcbsorn9Q+r
bi9rhnV8kohPi32hooK5XoyrZwN2wAX2InqeFGdXJtNpBd6je83CwxkjRy6ZQpyn
eaeg932dD0HxK+dCPtbZbrbGc5M0IjYA8eIOPmSuxRjoqty/hnReZIWLRr6sLZ16
gLDBZCAxrngqLG92jakx8P9SNF4c/lZJpZqKksfjs1dkOEXOyrIsxains8tGSnx4
USENo/CDpIamNbH9aIX5S3yFlIRrobbreRSvuCjGUbTJrptXzww4HpE39ZCpWzmi
6Iqf+OJxfq+Ayp3Dco4pMbN3bvh+OXbqu9XvJ2Xcg6fNltX4+yutXYnLfdrkS3o2
uowqRpOfXV8fP9avj+7bYOLUYEZQ1TgTFD8Z630I6mXLHiYm60Z/NgkrEAmPuXI8
YUPt6rPLzXvirzsC3cPAyvdqh1xNeJKGQmTMKYhDrLPB2O9D3cgPYya9P5nOGqIF
B1DODYaCD+zgT/jtH2cTsKcx7KfkYBaS9XJPJZ/15yIfAYuFYDPJPkssdrDGZN/n
knuJAWDp6agJMzZTA3ewOUh2B1vKqCsYX38NSY/80qnxgg8OvRUZSssYGm9hVNox
GpkW7cQHDfHeolqaED6Asg3HoR2gJ059K598khNFAgKhMDnNtDRQOLUTaHEvwng3
ShV8vk1wpahbsPGwwolb/zBkxub50EJeBTUwf6JI7MDUjlyKZvQmw/wyumeHItih
5MWC99/c8iG99WgitchUDMHteNLXHuay2TZMI0G2VxJ293JPv/pzWH5Ml6LE9Eph
1NIYKViolukM3cJnEVgseBnq8a5g8j6DBlPROHGenf+pU71/HzDNCHxlAGd2m6Ao
FqA7SMuRxtAC6gvJwkmxxTjpocutxzuSDJ+AP+LMifL7+eSSS62tSgfeSrFpGtEe
qeKenV0QzlQDyEw5AS+g3YUclyRGFE0rXwyrPsetgCOmxN8xRKBiOIesy1M8C0rS
JBR6ZRSBcj/SB6g6f+HpxBvABruIAyeQ4I1OKmRL1qHeD2y+ptoROD0OGPDAK2eE
S/oP1PwRew1fmqqRjXMJLJg6PeSx/HVbVctZmf6IYfbh5Pe5uu2OsKYgA4t48ve6
0e+C3vkCLgU2g8pepmqiCIdkSVr5AG+yj3TVrAd1TPQMJ4V+6NdYkorlIyklq9ie
hdoeYxRUo2TtNQ84fhx7BOiQd6hNVUlSmbUzoWA4LfRVRf697hl1m3HTdfQt9zNt
kU+b2ic3+t8tLNWzP27GKexZ9VN2bcs8i1oCJtku5+BJz+UMt3MaEUWe5ILyqnCs
HqOabDdsa5XiefPlkCTh3QGOdU8gk6kduOU725kWP8W7POUy6miCW8L0+dgxlerT
kNRuPUbl4X3K+JsSdi7cNdlaaVwNJeT7zenXefn7HQHZVj8AvsRbbexsmUdeRcnO
H2fqQ5gJwMnLtIDfNNCL9YnOBcH1kblfrE4N2Q9oKuNvN55rBmLHzBMVXulJPWTb
MNUzPNggD4uzzFvard1IyFvu0JSii+b2k57iSmIfTFvafJfanlJ5khcABacOM8OF
uI3VnGiCSSV351kwg98EBtoheT7N9YSt0mY0ixkRTg3ZYMEZ9DG2/GN/4TX1hjUx
GPDUBLFsCoZxn8baHA8vKzW2Vpj1Noi/jiwJNAPxGMNmsfFrOLvYTQFSAI5/x+o8
86URS17H1bIn1RfCVmP53F188f2JSBEBd55y2BLRXW1FTAXHEu78mmumE0KOTLDL
eApIlPHDk5KbOd8ZdZN99Lq/wtaMZ1linmKpsbN1rWg3egXqf7MkYGgUO6ntMS/X
S1PJsOlVioe95e32cu6UfPS6JuzHpLYt9W34VgriPQP4HGQmny6pmBRNBdNTuNFE
/MSlbLEfprbgYrHkZSsEiKPyuMg90dYav3CIUz/UC0CzQI0yGaO3W9wvPBcMmnCN
ASpbzfQTuxYw98P/kbbhNI5ui3xZ7nkzlbRHr4ZLcbDy2YZPx8xPcdi0vY1sZa+n
e8V3cdrizzZX0Q0sPySpkhWgratNAAwUTVYFgSmn+gA8UiLJ4D39diCCaVaN2kaj
fBqaPMPw17CY5Ep1MtaDvUGnTSleIcc1XnaGl8x9t7Le689J+zWOgNHgIIaPWXgf
qVdKVZUHkG0UqLFaXrwovHNZ/t4SeEUlQTTilT1IawrBr/eldTRZeNz/gn7yTUh1
Sw1eEOzsu0X+V+Zr0H1EBZ9y72tp9+nAsMh6YeaUA1PgPb7VSuPd3UFBR3FR3ibo
qN4FU8vXM+PN9cbaVISgOSDpwNlvvc5VlHdeXlUp63WeRpgd15uulv7M9tRnJSoj
FfWt0yZi0oY014cZCfGfPZrrXekfDDpBFUZDJbWSkQ7y8lhHgnF3wUFtY+ogMS4D
R9tWKJ9Ww9pinw/bWmNV/nWAaUWsZv6YbHjr+oeEBdlqRGzotojlclerqaxue6Dn
GQ0IqlOmUAsLdXDqItKYQkVLtYJRWeD3Mk3sIjKw8d/roGzboIAXIS6lJ/iE6bsK
Pc2IEctOt6rEjXr2SeK7e2QERteuBddh311Z33wRKUBoD8jmFVOeluCRlAAAXuJf
k+thCo7NX9bUjI/LsvvrvWhVEZBxKm3sjQyQ72cB1vRd+2y03sDIXrwdPfocn6iV
ASacSxVm26v0x4P8qXb1zpLdw+xVossmE2m8AXxihimfuAW0dPX+XkZkFZT8gk/j
M8djZoO+9TsbnXm9bel0Clllb9cmwTBqwWDZ4vdo5GWzH/n205GNRTh7vONJPgwq
gRScuE1AoT61/5yAc4ufXN9B/M5zEWPkbt8qNxbQnBIWTEo8kjGXoCGjmkh0u+df
gdqNxJIhmtl0u6gXAjPAZR66NhyoUvjmiip3BjB+arlZZ3lxm1saThXbtfkAjDHn
6bCjkRgYYb68QtK9xc2F0qA+LAjtCjgIvP8jocwQj0axe5Y+Mr2U6VV1KdD9V0lQ
zEvPOr2NKsNEHmgs8g7EQ3i0fFMFziqJ+/qVRq+AMSgz2e2xYU/IKCg7QyIyYl7Y
XsxQOgpf/nHj3MyZFdoU8a5MgrSPARBu1K8165lPsS2yGHyDMAs529SG9JIrQobL
Qa86LCNpL7ZaEmzsgzmrPL0owmZcDSGEqGvUVnXDM9FPWzFDNKVr4ypH97Kx48pn
3/GWAHdzZ7/g3ttCxi6PtiAGfXD/MjSBKHKufN+yEj3jndUeVsmwQ2QywC1/1Mty
wAXz9PhD7IH6DUK/PJH52ZmFKswb/ZfIJurRxKNcl6HrIzL7FXwbpFjYdy5IHe0V
J7rBANmhiBOel0EQYQeBHOJ4A0KqxEIWAqGbQIWi9ynNt7Lr9KK1OJ29t7IJlRv4
tusKXOwiqSFJi3VNi1X4PhetXFmE1D3okYQeKCJp0E71Ors0PJgpUXzUb7gYy901
+rH3B226Ozpu9oNZbgo0FgMIJePsaiAvV8zBEOJjHCJCNeICvhn653Bz6ZbwP8PA
DfA0OOlmtMxbRMGu2RfzdAxS4F6usKTffxqgFUSHAyq/X+0RbJPn6PgJa6lPLRKq
HNd97XZUV8NYxbCtxmrHoB2X8Uxrtt4Ld4xg6Y9fPLhHtzRkp7WmLcfGI1AHUSFq
zEbv8YHpvyf5G9skZffg2gij8OyuTSs4cNAk7h/Yh/gtlYu28oXim8IbUp1dbBRX
opyF0Sir3Wixxu5AOCmGGVQ8GHejsfbCXmytnO+kFnNflv25aGxrYlGNnEFgpPUr
uTThxHhyU+kbwmRRbL7n3D9E/7P79tYoizD7FtQDsOh52tPZlzE5h/URmxRlPwBu
G7aT2IOUow9k2+E6Ac3mZ6TEUg1aZ4rEDRxZam8K+aQE3i2JMRmKdvecCJgaQTmd
F+d7Mg4XAkZMo9GXJI4t5fW3EF05ICpJtMXSaOqEL/J34C5YlPGtElF6qcQmpCZ4
ZWE+wRb6rDuKafv7qpHTOiLH9+mxivk2mt2+drpruGTHZLgAKcwrdxrzaPqrvSkG
SQBcJWTuNCEY4AWROtkg2Mw1H5iyi0k9L9hLoS2VjzRkjfwU2RUsRUecjWeHA2/F
Q2qpgQPjKVorjAZ8XgJSq0bcAu9Hx88ywe3VubrVxbWvssH6WyQsgCWd8GL8cYLD
QgWYXyOucR1v86qvWSr0LhiWdAG910yBzx/pu0mken6+0KmcBW+JsCL0GBXqfGoM
Bm365IIUHn+nd+CmHCSRV7kwCH6NWvVXdavXMokfUb5Gu1QqGrOUtQWLW0Z4k3hu
K7OI/Vlem89eQIUQ8DwqjWfM9m6TD0b4Zn+0zCjnjcPz1AEV0wcI8yrvOqBhkMTD
I5BIKflg5RMgf2m698TQJ5hKUsMJsVPI59l2nDbeR5svg6++EJjuBLJUtxpfShE3
cUSHDsbRWaMmXKTeROqxCIM7mw9YhAXOtRJ4XLdjL8wDpdLQvPNM7FL2BlcmPPJq
0EyvF2BW+XgnzT5FPU15pl2sExIGCctSFDSl3IKYPRcFyvCxny3/Izye1JggyJWK
4fPWjr65PDuG4N8CHeCxsbGuJAYHBkEQSTgwh7ke1pWTj6n7mC+MfbX2Utxu+b/f
owOQIeacugYRaMDSrJbC268e7lKQIaH3U9HtsGsHIdPh2uteCp0nhGe/EZ/Yx3Bc
DzSZfLQGKXSrn6labtGPgarexyzzOZ/LujPgAytAurfRjPg81l+P1xzl5PTsFUWH
LqKF3Hsp5/uBsDM7E9CL8tVXRybSKZy4Gy1KZhgJpe4ke3ZbgV4Yb+smjvI2y5tg
ua6O1q3SyFPRdQnjitRUjrlsa35U6/+j5+QxOz8szGUdg5AODfJUdcOwXnHb3gET
Nk7M+VlxNNCJD2pjbVAU1O40+VxamHvyG9AJ06U1OF1Uy2zr+wkupJqQoKPZuLAc
R9734PvPJgOZMShmFx3qLELaX5NNOmXiFcKJ6tN0WUQVqReYxI+ypJ1PEdbFIvLX
GF6Jl2kIqBMQ0Lh9tWJk531KpA2fA8W2sW3j8o9x1+00uiGg+QQf0tqK5dL/YltL
s8BaWajDo4Xvw4a9FjV5rN1Zmy4UAAPjOqzkd9f7vuhumzHnLtoqIdoeL5ay08dE
QcLuG0MGpZ7P2kOp+rGdbvYl8YFkSWfBzFrOG5EbpAKqLVATcGQbIG/PLvZC73oQ
MGxDSP14v+spzBfEVvyeEP9zfPOW0onV9s7gHclnjaHXq4cwyPZkBygPRycm3ZLK
QmlgSpzwd5OqJzPDc0MJVRR0oBWBFV/4qL8Nf4qgeaN9YpSmzz+YucONrrKVxrMv
56Z1VVUi6QCO9EvMc9Fu0dkuXVFbdQhPKDZWFQc6xJb5NluSZzvzMczUGBwHPP//
C7Hpxa+vfOEvPtANB5ibyqPXOt+PiZfCeRX4xIZyCGzJpJgnTG1XVl+cFw3MUa7O
r+/iDpF11h9hV5TbRSncNzZan36/chjiKCsuFNMdMHSY6TTw2VQCv/sBcy5gEtbT
7kSzX9z912em38FgO8xxBhEHWd2AGWBz+9zwmsdgC4cIRpzH7sScKHGLqMMAgZg/
LROMthM67Hy0TF59QjxCZuPatl0NLShsP2zVXd47VL3IFAh7Yu70bHJdDoGDV1b6
Ri02lrxUzUzT71Xm5nm98BocEmCf82bFLMtcLFpm0BPO0oxYaZniSxj5i1nLkc+D
axbrJ7XQYTYfAdOaB6Ypy20AfavU3HWTjiZ0NY53rODE4zUOJYuKGR6gnVd5XeG1
8uPBGsZCkYNvZAuYVkHCN2Aj6Pqm/8rIPCNsshcMR2jzu7THAT2KEFIcp33jgTGe
sCsUtm01D0+sKlceupWNsMizuoDZWSWHx4IdX+nTRyPaZHWzI02oU2NPnxJqVjeH
ghR30dQPpGt/Zi1I7vQc36g1TAyxTA2783hZEl8LXD38IrO4uQh6i6mHwGXmOcvf
W0rHjhxk1sTNv5vuzqfmy+E1sIKWcttblrmBDFL74QRq2dtFdlgjnXQlZijQzeJd
6rr9fS2fKwlQMr5vAONIvoW5Bm9Y3BplMP8uTmfSzcI1F9WfCyATbVEAGL9D47fw
3Bu+kcQ1lfWn+elIpoSY6YptKxGjU0bplL6L/LeDbdeOAWrNIXYv+tcPF5wk7x24
CGpUVMYHN8zzfjluEjrGlmViiucBbjliG1koi3Qju2VwIzmCAB2fRVHUJmieGSld
/Q0bsgvirfvr/DHNGlKcNy/+4CFVCJ9fT2IHujlvOlzYhmtnyVLKA/mFMOQj552O
SohSdTSEl4R5ffcwCqOfInouKxDZTgTxMbXdh0TT1+FTJ4EYvBiwe8R7xMmhGjP6
Gwd/j18ZTnKMwBl7D31or/+2hxdHqI/E5FfIntgX4ahjoBeK0wVJ1xJPWj7Bk97Z
Tc51WJ3pGgP6T9NM2+ljarkQiHPhW9jTxts24E/PihQdg8spsJyJ4G62vJWZGBXS
UbpeyTd4lASY7dbH8q+H2fOGAAxoz/zFkN+oVbB56l2l3+14a9rvyuRWWkqr9tbU
+BlNVEsmcp69YuN3DhgCo+ou302GmdEvom+NU/zvrGSW1UBPOkimhZkjcAMgEOsD
eg2TwzjO6HvkWpV8DlGZxcBbZc9WrnvN2vOwu8s4izlpFVu7ti0QHszbMG/xO/Ef
XHxTouD24Df2oNQh5f6vtPd3b293mNJzMqrdWlrlP8qZ5k5gs4WxSDHJt+EkfiDz
qCIECGkjYu2MomuHd8qKYptl7ia8mHI2jkcaop00FUWl6xRv3NgaFjuZ+tacUu6J
Ln5/NvZ3XsnJpW7guIk3sPsuh8zGLYGz0ef6vWM6CgvV//LNDddpCObJZsMZVhDu
Gzm6w3O2dV4Dk1kvsI+Gm5vtBnXAiXtwG7rbVrFqoaz/ToIOoJgmNY8aMVfOLBCM
mrGmEdGXaPHUWObLmohhUz4lPJZzEc11G4K97aquijpIkxIfScdrcCwYMv2H9Rmx
959X3VVEbQOdmR4I23ZGEEwkKKq+ivFsu4MAYMQqOMkflYhNxxQwr7JZmu1O+jNk
L4u40lgUpT8ekgAyzrDw7PCns9s9SeST+fyslwP5pXkW2TIPVCqHl06U7tR/5Qjk
dHQfCEHuIOoGFXD8Tlb/pGxJIiJvjDv/fHGqa6GeIXa1OgruDcYoC2xJpexMEpCN
RB0cJ6JYks1crWFCkmXMLC28QeImAP2XTqiSP+wIlkUZzES89z7DrazFKO2dNBtT
zv8bDt1w5rStEZeeoOIkyLHjGeWr6J8ZKtO/rqV4tvCjpb66UmDKA84d/yQnrnN0
6Li1I6OPLUn2EIqmyaArG5UCfu4b2KxghkEHHCyrrx2wPcSeKf0oerZmyAGsQWVN
txvyD+EGYe3+oUEViGygGzJGFH5D9OcS8gIR6QY3ough4UciAs/QLPQcS8VcI/5h
xPR5Q3uao8JupaFd8Y9p3Ego1i5t8JMCea6pm3QBvm/cW6OwZRefUeb6bapG0r6k
O4vfIIoPCzNEJSgfP6GkVfWvSy8jGfemkgHTNbRwyy2LVFiVpubbFVzrOzCiQqMf
oyn3Y6Fn9gcV8hwg8HPSIAw73n9T3+tCwBwCBodf9XNHs7cQVU2aI03bHqLwhwKe
KJnwY06jvLs2lompnjH5Wc7gEGG8R2TKm1JXdZEfOp3iwUWFFwDyZOJa+T0fWcyi
GQF35j2VLq+IK7z8D6KLXm0ag7qMxKTbY9Yv3kjnGWNA9nU/x1O2DI7IC3ntu9W3
XoKzu0+CqoY+f955ksf7mxtLP2y/08AJ8yh+NnFQnSTxSEdg5jeZNCXHGtomiard
X8Ju4zIvvtfGCK+emh/qe5qey8M50fNAnQz9+bwaqAY7Oc+bASFXtqwiSfPBWu4P
W4bGAPzoc0FOSSbsRiZVocmxoVSTqVdc2DAwYmtf+ud5rd0u2ZwArnLgSaEyqWhB
/aeARX7jElnn3+zqSGUKuc4rWCFOA65/ieHp/l/6W4jTDMsQRlzsBsjIHWnXyoKm
7Vr75Sa1+8J3QrBH2f80qtBRnqk/MAG/L7rOfdGFUUUrFXultbVw23vqJzhC63Jo
3KQgjTYbB8O5l2W7hIV1x/1dwfnc8Zbi2e/IiBYVbQOsERVP+FeE+8IPGdlSPcK9
s/G4km2Ff+MIK7GhynYj126U3hYTTkd0bZQjFvVlZDVbw6epmmA8MDstsTsWTO/I
2FgA0NukTyHK9eAHDWBEhIv0NvjnUpAwG6ygxjGHHjTuw6XPO79cLXGVrIowwUif
0opWXwO3GFz9+nGQYrgj4+/89GBO69QEaddP5TGme3LwaacOjUGPPhulMQoOC9vM
ikTYY7bzdcBTS80akTTq1AefXZ3fMlhUZqA7u7EPScIXvv2Iqahc5OpzNI6lGKAJ
sGH+7BXhlkL+YXK08KQ+NkDln/dMZmP0uLSF8wfeg5vtjnwRcegO+j1clK1ZLxB4
s8s+/0JEyKNVXfaLfZPVvTT13aE72MA8gR6+/LEeICwQNe96PRklN8mKDS0xzhJ0
XmB5oSgGkN1r3RK2zsspW2fKZvxO0HqbCpWFw54HLXXi49e3GxYnCFM+kJipabGq
rRVzhTc3k9RW+weqNZYh/1nZaQX/7pJXNCXpS56o6hByTuxD1SN3Edm5I5t/gSUp
SRW0OReNinElez+R8CA1GHyhKez98MejDA5lTBoJuFZNDuPdrzci+hwtOu3PCMsm
O0Poc6ydqWQaE/k0VJVvIoZtmh1kaIiq7ETzLenjx6PM16ljq3CQd+yheykvGmst
jRMRSRBnyBD7fbNMQVsGGAWqBwAW9ouYD7vsR2pyuaofAdUIPGG4g/4AAUQq8W+c
0q1OJhVGMiWED7PahJJjQB5A5Xmh+hg94ffoS/vsNjsjb52o7WQ6SiMw//LqT6O+
TXO8Cjh3Ykr2d6WtuivQJIt6DM6obFq9FmO6B6Y59OWxAfoYrVDnHhgeEi3/rNKJ
S8BbXJDK4HfqH/cXEg/x9rxKnN20Ku/8eUcEFtFa2hJJhx8DE228EBZP9ZreXEpc
ifl4RngvrD70J046QbcIGPonjpvi9BMS2Z9MThYcaPVtH23jBa63F4QCe92YD3sO
RBlCDAUAPzHYnwqksngKdMcPz2je+7XQb2wfaOp4CeOng7DYxx2x0jr9OzUmGElQ
CK4v4v1pLOhsUct0fUopx65xRb0b+9maA+eYHo8w//10F/Dz/sQgR/6iDlcggIGZ
wB0IoyRTwTABCLNhHNTS2H81xkJY4wkbs3DtkL2q+OuInqttOwtt+2JG2x8v9xkn
uf5Jm+CPBhVRKaujnpjmXzv8QiNzdSxTtch0Y+6PDX6Dn1BqZm3OLHNbWirFzal7
D/VYyB0D8wI0LrJVGsUTeXvkLNjwPJYfAvN7vATw/ZXVEMcNRJ3WU0orSypMwDTl
4kNDhLd8qiALgMgb3qnaUzzFuJeS7BD1sOYBEZe3Gb66E0K0G+qjwSFwjZG03VXg
aM8LE4OrQ8p6oOIjWrHrf4o2IKUtYdNyKINmHPgNPCmUyj9TxFXEVwAKrF2Aj8T9
yq+dWLbDtvHDDgO3IlQXBftXVQgi4pCn7dVHP6p1L6a03T+ANxLx/5r9YS3vB9jF
T1GbBShiFRrY5/Xus5oaFbMLPgTOZEIGCp5DyO64Mx+CTHMjt903OsEX4TrN0sUF
f+tcu9y6Nb33DTCGx0iDJdYsWJ5KfuwGhCA/rElCRaLTfsSrM3lyyFjYBuv7lbzm
ZWHWi3LBXSSp8Krj33+TOFkVDgQYA72NAQ3tYOITTAC/obroZhVG9N4F1ELLYRZn
tAy734cb3Sd4l4tq1jza7UDVGMA5+jIHPiDPmuxT2oV1gSirsZhYJ2TIGqmo9qSd
PrADlIhRJ1ngwxzhb6JB+651aMV6lrTBBV3KGXtEAhrho+5+813RroLz6HEaPBfB
vd92Gygl/0f+ljFMrgQP1xoeSatSy1w6Ise5ITMjY6MgLbaclCIpG3Z+pjf4dYf8
/WHL7zBBTvmigH+pig4Zq2ub6COyq4BR2Wz3jjjxuVzqscbugCIQkoJ6OwVRlcP3
OZOa9NOKJMh4vhbosybk3zc77jZ+qTrsZvBrCN9fp9r2yLc/tg7iofM6xU+gF2Fm
BY9Btk7KCWW8OFiaCKvxtOzlUTq3OOrM0paPMjXWtyzgbbiY2UEgVLOWFsyrHLmD
gl0pUS9tj2NpXges3It6pwa0dBuCVaqAm0kETO/F+hEJVmyAsRhJXqwrpY0zRftU
SQEeYFYQc4qkp6gf3h2Kqb4gFmbhZ0ielTSD0VorCAttZriEOBh+ISIVThaosDoZ
KiCqNjGRoSHpZtK03+Ts4FMIUZflHWvc8IgQm6c0DXkLkIXLQd+y9SmvB5KejwOc
3Lk9dZ4ttDFQbxnATA2bxS8lY5j46CYNraEwebj4u20jjEeTbx37ok27KOVPHiq9
qNvY7810bPq6823doxy2TtdF/BZ1p1AYpJoPD8Y+NWtMLZGHjQdVJdC4c4KhTevS
vxbmXu1SP9LKTALeSk/cBp1epmZVdeGyU6Gr5oE1SJ+Gly3w6firanRngYm6yIOd
99fzjIusenFVFBtllloEUcNDR6NpzTu+IvEyynQT+Mvsr3HL+kL6Mf8wir8HRWUn
kSgNhIe4iJ0YV9sTwz4jK3AAgE1gwJq8P22yJZEXV3N8paML5t7tE6azhoUlKAzZ
QpQurWG72Dp9jE6lB35wgzp4VMfPK5dA9dLwjQc1R3RLjSlBmzqQG4ek1A50mE8Q
vSqWe06p78KrlRaO0jWYAijh+27AfYGMygmJbMV25zC7iiUxnTc0p8O09/p8cdpW
xOYzQen9rHRc6bAJCOu//HxEtXWFxnzB/U08rcDqnCARhMPBLiHGmz1EHQslMtlO
2b6+hHVaQ4VMOSSgM/0u/AWuNwIqEHmNSq2ifoOABPGP39xAo8b8xc/OI0cth4qP
K3K8GaVbAF0FOU3d61y9iHSUgTH/Io81sJeuBJEsr2cXOulKMQGpX5AjTK97rSyt
9uM2QD7CENBaMq/VjjZnwuFRRGK95V2p6dhotlOGj9N+JvefyV/fd/nz+67cdrUE
XtXB4dT+luCOkOvjdn8bXHhsGwneTPxZpusae/L9q2qppaYKjdBXGlaJDJCEXI78
NwhcEhxzstowlWkaDNeVPTNsGELjyNedB0q+gIkx6NKHbculZkcd+TQTgjOwkw/h
DfIBvo4k0g2kSTtHtS9iYbbmhnpd/rhm1qSm3ToEtGgIRqrqXMxqYPqu7T9O+owH
0HcIuHkAH3XxO+5+ueBQSWnV2qdCdV10edMMyioLidE8X3sWgmFxTKtwbIJmh14O
WNlOIHWVm6Khwl/GF1RExwUhRrNZ1UWT7ixYBc8CKA/HNAa60gxE3ld/juPEn0/T
mlm1aQ92oF/A8Nh+7DgML1GqejIJOwdyWHahSZsvNv9OTtefBgydOLFVaTM1YNrv
Pl0hVy7+xrwxYPwNOHCOef3aYfshZgpVbnY46VaXR93ymu7OBKGws41KEMgB+J8+
yTO4wpmizD3+WPqR17tUDiiV7ZHmt4ysZpcF5w6f9lydDjgf/1gCQE+S8UfWhPqx
QJKY8rNdsMHep/aFH6o2dsgK8BQ8kcPOmfZIbMTyBCZRHqGJqjhuuXswp6uqmNfE
xH+hYz33BbKDWr3sorZatOgVU32Ps/LEYpSVpykVYfcvyjstBs4yIw3oaCsHIey3
b9BssBLOIjJ79e8UzaYzas/LtCS2WhF5F525+FCLJIoqsyzmvnHPW9G5KFz7esOH
WUewp6qLvWk0CQsv+fHF5bd+8gN3i1BaN1SOwm7j2h/OFi7tgRuYlvcHGmtIuzE7
peg2ZaSg3YFRXb9IN+ByhvnvNdS/+0fnI3U4IeCw1qDJ7osZvG/Z+EO3y8fYmgaC
LvzWPrwLciJWgJ8M1zsocdyaq1AP2QmrMt8bdUzqC/njBkd4B9Z3dlEmmdefN9xu
XFVodCbLMk3A5IT/mI5XMbYb+Omr67+KoxopkydHIcn+fqjhMxRwtYcV13wLtPzO
kpdCdVT4MAarxqNcuWDyxoBy6NNxe53di7I2rz+RRG3KYwU2wtr4ZHmpYbhukiX8
oXsEFBONEIMfXEwXidp36oM46bpWUFeaVD0vjdvVcNc/UbT1w1SUtUiFgdjIcqaY
DTCTBxE6NgPZDfEZAbcy/s+OT4GRY5SbfU2jSfZib9oji4d5IgPZdjD7YRI6U7Wf
JOZqUTD+5BKBpzz/i6UJicOqds/xcm6BXm7lthAJBuX3eZcI9sMc313ts80sMzsA
DAfHNyIQ3DcXwBgup8+k1VDAl+NPD4mp7BHf6ncWFC7R6VoKJL/ihNDj4tOEEwqt
vP8/W3o837OZ8CzqQOP0YJu4lYdTiowG6PPzBysGflcQPJBM56ex+l+7+16JZctF
f0/uVFH7qqC6FA4YWCKrq3lmkFSDj1OUlzRWdnoSlp+mcilW8td7mZyDMt4PB9yv
Ul57ji5y7zNoBWGIvpO+HQGXI3wUtKzWjDK/2OeQ+Q4qwr2AlPqt2nfOvGtn/kQD
aRR4VQY7db0xX9S59kpdZLODMxvStkotGCM2BV6EVyBSYcLs5POi0QOtAv4H5zfe
xtizWI9393v33RFYDTBbXL6XRg/31OYAw6WgEtRTkRdbg2V+EUxItDH36Kj/JJOB
MxdWqNcCmLCT1O9gHConvyqONrdnG470XIaSsL44PkE5iJu/LVL+dgOzGJd/DvS6
W3uGLWA1x8cZD0IdBzlElcWgwQiTXTPcWZBl0BOjbmVisgw4R2vfyH2AxSFIU3xr
YCdEUBEp1/cULOMr2daSeHvlH92szRwY8I0wjC43Sc7RjxID6lf5+1PsRkMQ4hNg
jbtVLiWnrg37KxtYegiM/14txfAOITdoIG72WXFky383d/hFWfU4Qg11a3RAugKI
9zvTmrPel9RWhZN+4NY6N+kv6GtCjt3ELbMxl6BSBCauGrW208gzPWKGd9Y1edJy
xI+MQXoA5sJtxvlkvmEriI+pE3LI9K02GmVuTsdLEX+UsqEOa4CKv92OpkZmutzc
paQpQpTmLIyhZUEFi2Vtz/QjAQjJ/euRPZmTha+6e1zHM2zotOxp6k2Gm2r1Abos
gtVzucQNbPP38ftCz8+MY39E0bLmIQdAnir/3spvhBgVMCIE3mlesZSLtPzCiQ8S
J+X04wA2idda621UVpEV5Q+QVrM104SCN/C8p6k1+o7HKsV0RgbBa1PyUAICDpJn
ch75uuTVIaQSVetjZWTcJVr+khFFe9+IuFbqC7loomSyh1l/LIYvBS+WHypm6obV
nad95hUVUrX7FOYGcWSP/s1PYEZBOFAyZxkgGAR/ltCpPScAkvCRvfJDIw1mkdR2
0U+clfEYJXyLQd+KRzdrGJW++l52uBCCj8MU5qPEHSgov/VIgDAlrvQAiW5vhrCQ
tHSwYgCLRh+dHCvHeF73zTUJbsiHJIkiMntuOQF04HPBdZCxDmy/g2nm6ytlNOT2
BUfR5oMIWD3X/jHieoMsfhkSmFGG7SYo5EPnFyBw1Gy3MN1IPCQaiLgEXix9ZQxW
H/xW92uqGFvhdz7X0VFy8L8uFIs6cC7TdQ1Tu7sa4S7JTjTdsznjRsGXaIWR3m8Z
QUBv+9L3Qdyv7yNzVhBwEtkAHzR0ALO6kublzt4n36/LDvcX7cVJ/AcLS+IXPBKl
Mer3RnGsAbsZxVThN1felLJjXexuxdm+2waYy5nIoQsBkIMmLe4rXJU+1Ph9stEj
4flAHkLXabiy9uTivxRrK6cyeuxYeHrVyEe+plYAGRLk7UfUyTnK1anpmn6gO0D2
yNfYaJOyt8POKRwHg049Y+4CjU4XX5wIPOZq1e/Xk0cNinZWdoDCkvUk180vCAqn
5CtPKCjKdDx9vHCegf8GWcOAT/4ih+Uzo7qDTbgIdd/RG/9cJ0KGOO81OhoMGiTR
Xd737FJi1vh8Id3+6Pws1QibMLSIxxuol86EvsoSRoNbkdPxMpR9d001roq17GiG
Q7MB/QholWBtH3cpV/SqzY+oBKHtS6/hQjBAvnlkCqIkD4XTTgT+zzeFgqfU49Dh
4lZn67DeU675W3W8AYTLNvqCubmXbdUuLtW0Y5JFtJUx8RkDXonzP/7ZwLpYNaI8
aEd02yUgBry/XtZkP3g3Oyfp1Yw3eIO9i87nvRAkHIuDgRriAKPn0dB5iwdp9tMk
fgZjV0aVzYMxRFXvatLKbODyPTlv2XQioeKJKtGhtlPvjlJRt9qJay+PJlm+TWz3
Arok7GmVVvoaArX9drS1fHKLVWfvMVtWiAL5RktmSG/wlq7SJqpf+15bw/SZyG29
3570KYpbbSzk7D2QmIkYS5kUn1QadWMXAZKoyV7HfFsi/jbjrdbesKY+Spi0Mtyn
X0kc1OnT6eG8sO4vmY2+Iom0wvzMpiO+ef2IEw+ZJ+FkmvUeRfE0CeCuNmJNroBl
xuC2ncm2dV+Si9nOSabl4rcys7hl/X9AEhymBvIzHIRCYq69d7mtu06sTITTfF1r
crcLoQF81THFxG0ioYDiu36YV1G/Id9MauTlC/R699t27MIFW94r8YRMcl006ss8
q3Rg9zTJaGeko2ligeaY1A==
`pragma protect end_protected
