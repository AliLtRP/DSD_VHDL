// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zh+LkwRGqmUEU+KCOo3CYrb1ZWl6fyswQ1hmiJ788XOCDNzv8G5IPfMEtdNhJoBE
HLxL7WJCWlWpWyNsMrAnL6p29Cm98OOWjxOAXGPQnuSgC2f+uZ5nyoqOlipI8sFl
e9NI6ozbPjwXdeNWon8fcW5/bMqUeRa3oXOIXUc7Xjo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21008)
p82oL5xup4wfaJJO/jqXEDOOso566yyksW6pbqL0zZlYXmqwguh3D+f2jWAkVxwj
bwNYyqpsXwVYFpO1PeJS2Spr8wHlh29Ulh97v+Otq6XQZRWMoAQb+pHQ4rTzmZxb
LkVoZ2v1+wVjzhkb9N+LOx7bQNpnca9YviRxU6r0+HXsUjRXCucpeFTbuTdCxAB/
3ntaNq9NMIwLoXQ3xPJRorplKUHpMNrf1hRE6AOTfAK6AWGuxbLeDve1Vgf4da/d
igPTAAZWH9jl8nIKY8Rw4s14D89UG1s9I//oVbw4dOmg0JaiSoUNbAKcsx3FSfGd
RfPznWXiuJmAo16Col+MUsO8mLTp3gJ8/OEqNRIeU6fyXY82ID9ibBmdYH/O2TX6
lkuNtgP+qYqq7PFc86cxpnCo0IA8b7kK2qgQtr6ZL/93YXX7h+lyl/j3d4V2mfPx
sbESF5RxChfGdG2m9oOTlXUZNU+2KffFroIHSeDIwqW8Ttnoe/Vc/ye9JYlc0+bJ
1+nkMTNYseTeKJswM91s5p3PPrT78dAbXxYIMbEmtt+TCxxD9X//AYGPlYpYNhE2
mr31d96YO+hfvbJ+NdX9UrH6txojLqSxQ8mvxWK8iGSJutHwRe16rwmJxlFRwD0T
waW5l242QKqG2AZiwSAVTr7Gmln3gKUUe3JpFo3++EIk5YjTH/XWgfhjNZkpWfiR
rZ+yOe1Er4Xfo+cHTlpiwIVF49Dt2i3AHTViG0sRM8k6xbJJArZVLQrbF44p630w
Ab9IuNNC3ix1OyLD/IwCKfpV6FzLBcno+ec0tWXcu1I5XwIUV7etry0++LVJFh49
NbWWEZ1C2ddbS5Mboa1TECp3FnB5emgCr2412oDWSjHE55jAADr1i+KecaARjOOB
xVl5fbf/RyjIrfuL5v97LtLteod8ZD2xkfRVQ3YIMN+mPWkdLvhGKH4Kh7us7U/K
F8MrY3CDlxMxkQcO88gU+cjc65bD3lLyx5RCQCLNYlbKNrRHd986J3AphMbTKbi4
p7jLY0eoDfN3c3ipz8XmkuVHe79yqrE5KSFmG9UcQWMDM0qyeUmalJQ1rRaqcJe7
XBZbt3C5xRsplBv29KnMl0xOT44SwI9JnkN2pFEo89mzCsGLoS2BhHrGrD0pm9yL
IYoBJv5kQa9f5dTrkZKPD84Kjj/rxQj2a9sXZtAnr0951vLtHNmkbfblXpER2ARB
/PZcQI4Mk0u6L3GDqAXZksOnO56VgipGAj2/KEjo7MafwG7iG2dLuQDmXfl8hCXN
z0aThrz0p3E+MQ9wq84flzC/ZYvchJWzULIV9gc9SbyjJMHJQ8t3Zt8WTrud0rp5
NduhbhWluE3GfaafbDR2nm9IyJQX4kyYFZlIuklWxVY3P03Bj2OTANTDdwIWG6Dz
vpKCiXSwVBmQzDtQUGRMY0rQce9JWiWM5RHltg5zkb4VB2AHSBimdFaN+DBL/RWr
xdl7rHCLKdfM+0XvoR4EbEP/tzqBybim2g/XpFAJVnK2849JPHZHVaFTmrezI2Px
tJgqnC3xBdvfkzO5nxz8biTsnqX5QZFok/DcqYqrqrNHbvZ19OAJSPLWKECswG4+
txQ6kFDK27ir/wJqhwFxkEOgDFTCIa21baZroRiVbFMVTBMvoUiFRTD3IBR0JakK
XK7z4Zr0E/2VFteceukSQUFf2kJjTjUofyqsXSTSMSVz94HpvWwF/hdVtzdShHjz
9J68hwWrHvmJ7iewBM9Wakeboj2w1XeguLQt3A9zDcF9vAV41auGfL3BRTL2+a9y
dEnM6t36XmqBFh+wUkYHKFlpJnmaxmQsGAuGY9MjaQyBlf2WHYdKxMZb+eUqoFGU
7/UglVwzQ5QQQEJOvg9B3F9DtWYFFglp7aLzWJ89E0N/Fo3ShEzuX51CIhjlYE+G
bRvOPt4Hj79ndUpE99cMnLyfOmNpn99RNEs38+PqEuMMWy10/BoDtKiB1kYpdN0w
m0a1sgguqvKvXTyQ2UBmPM4D4Sc6C0JjndUb7Y/hmYFWrI59PMIhFMCFHPXIhy/9
cDllTWHGh+QiFfkq+wVdGX3GZzS4ME/SatC0q1BCjydHyieu/i3glARCnDvmdGrI
QwBOP4f9nmnkiljg/ktU+eF29FURcYgvEQKjoXe46kHKUQj+sD0LqyWAkiPST6iq
bvDhr7AaZiGm6H9b3Ikb7dBtCUiH0gP+Le2CPJCxRr6Qv8nBE3wgj7KhN3eqVeGG
15WEBal0lE7WbUyMbbYxASnKccYWP2EYCcDQV/DJIX+MmH5gC4/1HBX6J2/ckMkk
2LrDWXh+UmCFXrPEHoi4f9m4ALvHMI2cF3/jfBz7AkGeyHyhyS8zzZTcC+sLR5ug
K4onaKY3m9BNuI/VMaxtLcKgvInn1nfjV1DWy5AjNJonzSydbwfQNcvuAFsTSO3D
mTERYwywhN0UPXIIdT52wr8R6/ksPAH5ddxlCOQBm/tpHmpiHn0k4eQAmSrtfdve
K7mPBqmR1BDstDG7l2p0V8XA3tZrmzH+2Kkeh81/JKB6ALsgIHpsGnOKEYGkJvYF
vnWmTeljfuCwSk1Q0KdJoYqytTSwAruk3NyCdzljJL2ndZ0jBtWeKEw7dtKDsh6v
izVGi1KWmNRU9m1vQSn8GIaTOWJ4oV96suS5kVkZG4uD9AOlzXpPEfz3tf8uw779
WDzmCHdc2U7nuH8B+0W1zXiBcJeXMTpe2lHCie1/B9nWKMa1OKIQXyfliUZg14Nr
HuGdpeFc1O8YWlgcQEXoCVeEi4vL6NWpcvaEde1KqsmkouUFX7TRiJiH1W4xv9Od
P3k7e2ddIy4OZ/FgjQurZnhaobfZhXRYNiede10e4TAkoYsGzkixXfklj2/Yi7It
PU7F5o87E6+eDdXUCGYCtSaWKodgeGSJfvBxd6BJuSko/74xDgh8j4J+yPTO+UQn
qapu9fs89KvNh0f5f2UJY0jAgC7qiyh6T0yZtdLaeFL2vnY4HDv6ntZvm/QtWqa3
sK3qpoUa1xMMVg1qJZ6UbEPIzRSkvlSY4HM/3Rm3h6zAw7a2peAUhdnahG5Zd8Zk
qrBzsTPWDJY4y4cy14+OpIXv1NrEvErtsYAyRInR3J62Kpcon3CCLg8XETeyTjce
JtVqEYANRFMkWTh4pAZBm2m2cjy+MGHrQoIxZYoXBC25WHXV9NfvwzBgE910kZoa
Jqp3dFy1AcBrI0qILIoaywl6B+zjoxLPsDHBYrkYjyOL15ro57P8kW9SPuCltDbA
CCRJR8xJVKm793z2c+ZTggujcemMzGg80jAOY0e7QzxPXm1quJb6fRUh3mGOWQEV
wfB36ZZ4G2lG3N4IJ1Z/Y73VZrxEYsuQIa80PcDx1U/hAhUZGI3rnjTEMaPOlzMd
rlFkPdC1GgC+S4mFZymHA53jhZdqRu3IMHh0SsLvhhHT4y+DViz75rotTHr4xVqO
UqzAxV0ra66qtt/ALiW+99cpQ/KsR36m6I+ulE4wQScyU3wh83aM2Hb9M4BsQLti
1y1mZhbsjiOa8ZVcURl16fI+O0TPDmzMsYbsQhDtoAP1nY8IAakTSQNbCsrx470E
BFPBE8fk5CjlZ78SQVphDZr2QSjKq/2VrwDkGSXn83/ybEgZSkhB6YEgHezatbe1
A0dl4kbXOPzxLXj5ONByuV8STMuzBuTVpRcRR4nTmKTIfW+QUJjNg0lVf7cktoz1
muwKKYAIlKj2JFHBY3mBwk6pXYaQ1Rutf/4QO1tIGQjXe5/MG7iyMGS7p/siNxk/
FJttaDGWaLDJMVi9N5jn7TfpblDk/1PCaXU1ocURybNYgknHbOrth84fKXgRWL7v
uFcGpAxp8NAse5O4J6z5y3B4jnR0vDt+cCYcMnuAXTdtIvn6zlZBsJbRrguTKHRA
Qp/4ddvVy8BH71aio5rjaQytNE3r/3jNaGRVi580dAETVX6NxpRhrsDKCcBPXC99
IzNdnyHmGmZYjaRS05faG0Efp/JrNwR1gaHcD0DFopsf9Pz2VkBWV/JF+0wuVYFL
BVMBRtgL449ti6tlttnHgAcf/WZBGKqGNwh4MOrPxaUnGlkgbq/LDWzIp2yz5yeI
sg8M9nNx2Ng9WOkZeKbTGpvq/gC4Pyx16L2oXpXT8o6xPhJTtA+JNpemGpkKbOLA
fz9l6ywCReE45GQn9JWFDtWSx4RVw1dtBkNHqm2QmqttiJGgXy0smLWr9lzZ2bgX
Qdr/Lu6q+o+FJScC2y+FC6FxHLc4sNJ4fyBa2uXaCMXaJO33I/aZlCEEZGxNmuZC
8gjozEKVjc4T/CuTUChKz1vgpE1X5po7PiUMfoA07WR3ZpXipwOKv3nxDIzMDUqF
BNIxA/kYpD6OCGFKRlytlu20IvZhCspbIkpIthyw1VGMT1CAqCO0q9gd+wmBgNR/
C0ome/tA2sDVmfCmN7Hahy3CUtwqRgTuC4ogGPaKu5rfPO7go17oN164nFC0xvLx
Lc8XlgwlXU56h1WOoRVk2etHL8CXUtcTeFg3zvhNZTO2CycdhxQZB2jfep2tW3G0
6SjJLmxGWzW1SGTgRw5+M7jvfPNnF1hVULQVJXQzHRbFqT9yoQrYlT+xZHo0voxI
+z9Z1/W0GQf+0AX1GGywif6olZ+cz/Eg1gpq4qWrXNihxae1/7KTKUi5wv8fdTyU
uqVeNo2NhbloXuP1uDWwRp5tj5nzR/iGNpqI+m/Jjqex7Rj35aFg6rBFGn0VhO3C
SLpYlOyz1wX//jjxM5MB5HTzYX1fULmiGAxqBIH65zUC+jRDsDzq0K6YOK3QDRCl
/+2f9bI+xQKpJ4B+e56QuFwIzEGfv1KPW9c1+UUk+oa5eja2vDW7FpLFsadK8WHV
2IbhMtDfTWz8v6BgHUXo7nH2dGPBGAhTcDYd6KrWZ+E5u4DOASHDxOZrialxZa30
fOemtPoIN6Expv3PaOh8LdEw8qs4xNLMk7IuN99Ms9RASr9xvdAkHs8ProVgNJKw
pOBAxm3y23lbqZyUBfeHLCGE4nE7IqY3fylq+qoGPaTEt1Zn3YuRj8ZT7Z5014LC
Kz1+mugOT42bhHw7N7g2bDBij0gfsKfgrqvOhqFJ5RDnYELg+Lm6tjsd+N6x1TB9
6CgM3ouTJVmGVgT4rZk92iuhKIVPvvoInMtcEW7Pr0ofCy0xRnVh2BMG1R2YiGgy
0PsRCUOElmjaFENqRRHB3WZfpDJl80vnNwW4radN+I7oGdsrxqDNYBNg+k2bojMy
Eg3kjRP9mLZFPbJyl52s8oN6+xbgCJss0d6Wx/S7MkHL9H5d/ALpi2prLyfwvxut
+uZyA4X5cCwaJ7EAgRDCySPAn6hCnaq3q+6xfUCQXI9tImreYPuR9UxQRUyPMsXc
KVZB6geq/14/28q+2cvf350H3FOkjN7ylm6AL/3L/VA3h/j2DKsuZ2rQyAxohDHZ
VoUlKDIETrfxlsH2lC0gwJISTqc5mvMRZT07rKMNFHebo6z3fdhQdXy7sEnYetzg
x8badx5S5o67qNWrwUKiBiAbnOnw/GFusad33V6gffSMbpfUKQ9ibAUQAcQVqvdR
tIklM+L7OJkAewYfadJP08ahcUhu5qdt0s+To9dQ0YijFbL8GBxJtnNA98QBztzl
3hL11ufTduF/T1XTNBGnT9kwVtMx5NsxMX5eoz2dOOuvMTIA/qlMaeQ5/k9DKagv
plvqnJEXqB7o5lBL3VMM6/0QYfDQMCAkB646Ish34+8qAGHXMpKjvyJNu3r04fyJ
dqi6Ldp9ZsV8XLJWJKAPfCIZMx3pfPuQhTgml62ym3wMlWS5obZ1xx9P25NF6yJ+
NxkIUMvhGSdJsR64G2yyysK4/hMS+wQVERO62gzM58+jrX58qBDS7xLIlIfnyR2S
acm7aO0pf5VoF1p1kv5ePBsRAiEWeZYN/YL97EnyqhJBjYZr6HukvyLhVVptmj6P
3S8HJPQ64yW2gVsx1KdBbl10YCd4K+ZWeOdQ49euCxpfqIoUC4O8NYKdaLT2QC2d
sWaYXXsiRtFx7odIwtrGtj6rKhcR7JffrHfaqvTdeWp9WdOi8/KpJhXGZUyC+wPy
HhXvrQcCu5JcGJ3WM8iiZFa5wk1Pha2/vi+vA5bLTLSyYyrIf04TdB5I7fIiYdxr
ZEbopsFrwBDUosU8yoDcVTDwmtJRM1rSY4MkYLOioHFs8qKDmRasy+YoN5PIFiwG
uGz6BfIMUAiBfhimHiWU2fQufilMAJjrJq7rF5zU5o5O4A0iXvzSTmqyponWxwfh
1rB3t7Q1OvPg9Nh205WEGq1LrrTypTZih1giB3jgn1pNqZiothuRw1M+mhyu+OJC
qeXmz78h2/y2RBFx2SOSvwvunZZxxtdDV8Eqjs8wtuqBq4erZYSZMcN32sgET3FI
ePTpyEaCJj9CmwLqSxsDD3ievds27EbDwEfFS/4deR3Qmgfi+Pgx6BLQpGPV4jcj
Ws+vfc+r4hWI2POCL4ULbRQskJ2X2SjnNE81HP51aGRSzmpdgm9XnMnfp+D4SU5F
lxpfiJgDFQY50Dc3U7+hsMfiX6Y+XIEh4MuGAmP6BfQA9B/H8lERm9nuznd5QiD9
FyIQ3nQDlLM4lK7C9B++/BBe6WKCX4dPtb9fN6uswQKqwmETbggqTLWxa4CPJx84
CbU+D+oM7nfgxusaGtg8UTbR/AHS6se/sWsNNT3qycAMfqkM7xZT3VvikQO6uosw
zYqr2F9TvQkccjIW7Ogap8i2S1d1RWnmOaIOowDJ994Gl7Cb87/P+SLGO1cjPp1G
maXgduYndweUnaBoa2z8xB96gNkbp/rI1xdKGaY2DlaZaW2t8zhPuTiqS0lTgrZC
/tOLB+2q39x4Ir4XJJV6d3G9wqX4XhilgIxdSd14QcKlnu93NnvlJh98oQvNfo1C
L23gtXXDgJ+4M/0M2yROoNrEjTd+dnr3/Lqf/rmkHjn0q3HvM5AaZql3i7IrDU3a
AE5+BVjRLWw28YVAKAVUKD/gHVtJCStGwi/0WWk7DFQH6f3GvGEXZWsiqlOaSNRk
DVd97OrNDgp2ydAnZGa0udGkrh16Vy+IPsL5Nnc1Kje/SMUIqH2SDGmVp8iR2UaK
s5HGf+nBRA+rOV6fg9szluptH0Iry55v8UKSyCUsouC55AGUuwxgZ1ck6bM5xRka
AH5SDzxM32ogvZmwLOtaCXRJaB8XKQEeHNJftlI/QxKn/cxr5cjHO5gHh/QmJ1nZ
NN0/PFuUDKpeLRugJPJANuzrafiZIfmN03EMB/D6JvmiGV9uK7IFVCkKeb2fGLyX
dvnrz92B+R/ShdPu4aMznWz/RqaZO1cb+aPO4GFeY5re7RvwWHQKYzRY+YbKx3yr
Fb5mP8tb0wP79oCm7pCiMvZvbqoB8qAOoRbUAugu1lEg2bhTuEoMj9lcxZ1zKGfm
ymsFiIPu+0342hRhnR028FoIRA6cEs73j91gPGfbWMRILVZI4V5t8oD/0tLwRQRV
//bpm03iZD7B+zd9+gXbCRePEUa3iY4+F5UejBKGCJooBa2s7Ds/t2wC2nkQ6AaB
7kcs0c64unqpMD8E4JQxGfYj0L2lHEFT+BwIsM5PzrWLCbimtkS33Yre6UuHDreu
nkOhY2NTlSKDaXKnY8vLHXMBCYjYOzBAN8Ib65oFG5MZn5N8XqhvoEcm4lQ5Fhb7
aj1DzknvNz0ZJC/A92/yHEsRYNz1+L8yj2Y+Ut3f04U0Ij1oYf+MRnJb8pT0U+Tj
zKKykmEyu6rGEU3KPKLBtDSGHekY5cA7zPbkPd4RlajPINFoRwBdjqg4U8XXVAlC
QxxTwwQEqLQkX6VSaTtiyNtieZx0KjWCmDvIiIQG0z30xaW7j6TTjMq0sM76LFqB
gEYGbjrsmrTN6XI3oV560wRjHpvYj+0D8F5l2uxvZ2Zyc5S0ZZyUAiq6sNLf+6n8
cr6k6EGvj7e2YWm99YBMceXO/MKjKUu1OixKt5TTZFwWNZFkTY1BxKH4OkIx72pN
2t9I+zjT2vvzbTXKXDHuV1Xy2SQsflDnPXDm+50SctBBZFUxY6fwZdOMl0U0MxH9
Go7Rhm/4+t19d6kKLhbSswJVdwGPx1XEIYhGh11G03r/DdqzxX7dZlSFTcpUgfFJ
YgCgJrl70L6zFhyfZtE8OnNcnY4KKjrI6esCU7lQhdlgVPyDjd88f5we2CDFo0rw
uQVQho0I0hTMLRtjVsz+AhSnUa3kofrYdldFUoOYY+1p8l6dyQpeikryF9SQPMAN
+QSNbwTI4VhU9JUZ/3FbIw20fn3I9Dl1p9a6hJlsy58LpVnfcj8NhK10cjf5tI5X
YE1Xkd3HXuub48bFHhzXUXXzFshsAobqFgPgG5Gblhwg15Lf6wCeoFdkP7dAZyej
IiDhZsPygelL/UoXtHu4KJxRAo4SuTA98JrUJSdQ3XRbvCLqnAeO85E436HfEOky
mG/BV2T0JQ/fwkPxQjhpi1bJJM4OQjoGHU4dDvAXwzW5xLp8OAUxCyCGRSbXkeft
52Q7lN9qbVObs1ahDX6oldbrHNslLx9IH7IzM999xrQp5cFXC26ziIgeHSXzEukz
CifGL905J4qKa2MjysS3JXheOR+kj6c/GWfMj9miUa9aYIEt3qN9/kpqWasI4R9d
JNnyW7sgSEscJRTPCfa5vjWeGlbMLGEcZXwVgrlEA6iQj/F3vsvRylI/HI7vckTO
mPjdOuUFMw7hoXhsxkbJRoxTMw43xjik5WSb6enMqrZ5vjJFwUhtAeZ+zkI5hvpF
zR8I7YdTln6OXqKaCS7iFmJtdbGCW1giTZtAbitW2QfOr3jhMO6BeqI/bU9xti9c
hFnB+AEReIxm39pBHKB/ASGS8twnUl4N98mnJUKa0N1fHpHACf/QSEOqfB1ryQ75
uUS/Y4ffiffgg9rP/BBuCC83VDbl7yvwwHBtzj9KWpug2ntftj9GKHu9tzUyZ0Zq
ypveDe4vK/BxlMP6dS4HHfC3cjPbtu8uWfv/Ktreqwhb0LCLNfRxHS7Gaj9LQSWE
B1UIOpNrfTTlKrGjK4Br2I9lWnk5n1mrKK7gn/2ZgGXZ8y+y1mC2pAJfsZ5aXjc8
If4Obg9yZM9zW2UTDLsNUeep0+KS7cS8INAiCSBkIRGTyNnln3iVYIhcj4mpOs74
RbmXs18us1woUroy6G1UzGZFYnc2bm+XvAEScBx9zWWRw5vbixUw5gJ5b3eNOVBr
qH5xj7bM378saJGY1zKJCW5kAA3VDl6eL691YgMxQ/b5AZiuQ+Us+P26m/EE140+
qmV7VBVLuU3/w9NHRVeuNNskKZHbFY+jULiBpUR8cME9W8vOJnZP7ZrZbrSbF1Mo
hj2pBZ5PG1HYA1W1C8SLbBd0cZPEQxfKV9/6mzcj8GYi4bmnIeYiPM6urX1Qb3LM
nHjzGO2QqJBVqm+fLsGY2CPe7y1Il49xArvcyvpo7Zi1JK9ngI+N2Zw+nzAohfvN
3BMGvYyQoJNathQFMaf7HDHw3sVDO5kqRHDsLN6B3Uk3RrzQVutLpMfy/OeWas9Y
44R2afqFwVA+nlfjO3j82gzFunAg06K/yuFmLDPcUD7vwR0KmKchQwgCXCemeDeS
qDBjLAu6bja5j8EghLPsivrUZvxb3MVO41QYKVeY8ZamYoLrIRTEfwGrLal93N8s
SJYdze7iKmlFg4DrlPi0YsBlGgApdCGczUWJRv0bC7eoXasKhmq3TgPfPTB+pVgJ
dKvuvsGzzGjI81JSB60JHRwLiKGTwgffg1xOabQXoE/vyF1HAQDSX0Xf1xmfqqxr
AJwP1o5LYDOMySqbZ073wP3wvARdjX1lHEkWWrD56lx1EClpTJMcU7dF1ofKURCX
mhiq6fuR0SEMnueQdUo8whSBggsSYzfu9hRBUEWVo/SwOX/JLJsgptL3htr9I8Wy
IcjVELDD04D/SgPA0u1qCetKPYPGcwnJefwrXiMOGL3HT5g95ygzzs5nh+zr0eAS
iWGPCCJ4jXb3gSSOasZ+oJ391KaP9YeXKq1kLiEJ6CjffnsUuNd53y1YPSQKTgUG
cRl9OBQZbkh2dLBO3AyZZeSE8rCBfsm9nhloHDDPq7BxPgwOP1cJk2gacuqhLl6/
FEn0h/+51qoW7Bzgkpay28Rgpg3RgjYmxpzpNfcRQA8LAZwacINpNTOY7xa3ijTZ
jdAZg45p8hllEhAzf65hGLHJg7+uijHezXLgUnLauMtZ9Z9qk8TG4yl0aMoyYvMD
JAqYfoglwfH5vhspd7X3rJZCP3ZjrkVptj3pPKzO1CBJUsZkBXhE2CDDcHlMQZCv
Qfe0Z+RHXIGshZeOZjRt1u7FpeVQ6ex49/2QR82I/iNPjWHGRHigmLw/hSbOfdsZ
vOIiBCEbu+I64Kxhxzqo382O53HFue7mYZQM+D0oUul0IhnQiFRAs5sjTDsFekOt
9lRRZfbyeI+eKXZUv3eL6mE42R7464mr5k73+3CAdwLRaheQZ9xGHwbd1RmvPsdH
oBGURfxu/qPL1KvJa9elpWl1aiA3crpiJVHIpOO8C2Tn2JBLPr+f10z/9keChp/v
C/w5F24m5JM5hrrPSz0KmVzty64/3PTYJiRyCT1Wl2KaMmZ+i9dwJXk94JCRfN+l
UQtK5TfmeXtzh6is0CSKdxSnFr+qlmuR7TsAy5UxUVxWNN8GPFlRRCEY7M6Qw8VG
/UEaeOi7wczsWR1hkEEap47fhEBrbPO2kjF44qdmnn9RHEzsoKRXQCkQVyOmmng6
anF7UKCJbn9liivvRukVTvCLxzia0mTIsKtreRapj4QUJnySG+NgTULhNQfxtp9f
BhuPjHYbstXxT9CM+sd15wBEGJaEXR0yc3f1hZqcMv9FuJyX/gaudwCMn/KDGcOj
OSEGCZCaB1my6WdwzEv8hNKF5w5k1fJPeGcD+0781QuMuH2EHV4rUY3AZ8ckdALC
DrGxJAqGpPAUY6gYYcAUiXi288gRV2eXKPzbkZBvVXcK7ndHMOHj46iUVDmzhPAf
VVVYDZPf9Dhlgm/qXupDUNCFdEnJWzqKQrLp9zw+eocesdxpj+j6lWyknVYRAEAO
zVqdJ+/Q0tZqnuFx1yHXcIeFOrIfiQTCUlQyc5OsZpceUNJLFeX3vyp3F3rnVZST
5vvcwlE8O71Kp4uHmX6DWSP0cWxxy7maRgpnFwfW3uQtbeLkCyLOAypLZ0xsiJNp
DiX3ZYDiHePiRT0Axa/s54MnUNWp+bNttdSTW9a6UnE29+bQw+7fjEokQlDyY92H
M0SwDoGCJuNkJr4iVNVuLdDa1f2CnanFfsfK6XByAoiCf3S/dwvu0cJS5zNM8GEI
+fE8tXyg4RZFi2e2DdRE8alxdpBGUfDOpqDHKlr+yHnpYraP4YL0aS/XcIBjJ/ZA
GFkjiyg6/OFmn1zFMJZwTtuPozC76SO5pMlRBzKZ8uy6vtA+4W5aedLZju8Ae5Oa
5Ax/osubMOuvj1obDmeP+VAhfkV8SomAtfnrGQx3jjq0zC7yMzOvTIjW1F3Y3Hwp
nCpkR8i4/4d5Ox9MKJm+QX1X7aizdQNuUv5Dl5lZBKA9IyBhY1CS8H9UWBsEiHHg
sd/zhsnw3et4wFPaDZgLxUHBBeg9QCNfL4qv6oxZb/L8uuEI3XtXFFOCvHFVLkGt
aqqmTAZApQ+5Y8Uvq2m+Z9b8lyMhwFmgUX7+el63twyb5r4otsTLqrtJ4ohiPK7Z
mlTR/AIsLQPrgOP5aCfnAU0vnl7CSm4LXz7HWkQXZrXFM6wAqbiUvGX5I3v4t2ir
bYzIFhPZ1XE6R5ImX/LxytdP3MbgsFhW4OsR9bbLTFoC9yS+t1NTIeORUChxrDaB
fSfmgkhTPU5OOgVtfaiPaIeOvrMYGFJn/6hkGqOC/mQfjpknHjyw9WM2XH2wwu6f
skR0rtjGE+K/xrERf9EwHuxQ4h4CSBBQyoV46I2ueTjCew34+Uf9aF29PEReorWE
RbdS6/vT17ojqY42l7u9begS55EuXbpoMY1LxXzawcnCbuXspln8LBiKuXFGhotJ
/ZYSBiTfwiwdirjgEjZ8zCl/WSLdefDnbZCa6n7rXQgJ6OTMdyxhiDbTMrdQuMkG
lmRR90LCe4RCdRW0xuCUPJ3spkcXNQQ6E9lkcxrIyib/1bYzQ6Prz137TQ8psf70
5u3wtbDmyWBf5JoBuqjb7A958UB+zfv+cbKtsbHdOI50oCMMaPIjr7OzoHGtG+sx
Dtb0Ip+9xfzRgmhRdGzDzVY4iTLl8HXXI1A/Tjg72SitCi54HteulI68O9wcOq6g
PO7ypkH0aiONami+qq7e/USsjLmC2WFvx/Xa/m4Q8p8D0NKF3caOLeWwB7BE0GwL
j9P/hLk3OGdoMuweTopiCABCMh4PkyB+huf/gMmQIUOoo2eomIoYXQsIIM+OU/yF
NkndRJKDyb5jNQIwLRpS9Nsrt9a8h8O2MBkS0YB4vtXfb8kJhfd1c4caKTMm9aTV
cviskKiWALpPR6wk/A1EeJs5DRjf5SCTIy8iHBjs+L1/HBI4Att5KD7qOxy/22S+
sM2aHiTv5YpI+2WbT951cT29SAdx7yZwaM1ad523qh8Bhp60eo38NpLzX9i/8JaL
lGFy/GlizmBY0mHQ3uG6wmtQaCe+vtl80/niHuq6a2rr+EAJUVxhFmCNY54RlogP
jvISK0sIdAdSHvH5OYKUW3YTIvpq6bFt+iy/m06QH7tViy5F5wIo99Sr+IPSyk6S
G2QUXw7XeKww+4bWU4d48vEmfb4lNR6wxQEaezzRqfaq4Fo2aGVh/1JDtEFz3AdH
f0KMKXLlxe1k+OugK9t3pzOLoPZ874+6sbGS6IqR3+muXlV43recv4TKMlixGYpQ
rLKCfLLl7RM/8shkmguyOOM5SUsoyYF9du60tH/A2kicBY/juUXe/Tpi/3eV0lNL
YoqtIsHuLA/N1we7kyX721rHpW91PMMRLioF2xRvHRmxIKLUhChyM2GChcGj/W7c
+fzy/psKvGKZn1wcKFy0/TLEO6iopg2rhBPehIwMr2u5FrkFoc2azvwM+QuiNAf1
0+hE/0iWOaTk7/Vx+llaRug0TmMYgqk4Tyb7gPO0jWY18wXHh0KeinOueoMfQSxi
Q+qsIhPgS9UhG764fy5wHf/iSYKnoMoPtwbBm5wmjnFe/0B9oFvdFbmuB08Fq+LQ
t+ZOX8z4mVixoVRYDZUs/6iBeA8/t/1pqGHkfUF1JjeaxapogvGP62baeHwwl7oy
4JstnCD5rYsXOfI1O83JfwCVgq/1PXwkZ/E07qBjfcdDtpWpKD+VR/qZDpExwDAA
fnOh1d7HPnzwBI0rKxKfqBuNn3SJjQOGyNEcyFygEwPKl85MbEGwhmitGDRmzhIS
5p75XOTMJ2DxQbgUi0pDEnMnxzDjp6w4tqP9ywi7Sda0cPSNLNbqmRJCpz79CIWf
JGvAQ2D9nSDX5WWLz4WobgQ0kVbQAMsNmWUuqHQPVrP+pmMqBIgnQZf2mVqd/9GX
pQikGz2TeI3udS1rSePROJRbuQC8OkFuG0nYTeGiI6VjmsIudi30muF4dFIxm1RO
z0UShFNZMGMNVdMf4tXRLu3Dn7/5qurpP5MSYXbWqR7IXmlo8UggpdPorMbTFYOp
v5Pan+z4Y0q49pQ7sTeY8EzsirssN6zdhsqdRaFTKQkpvJlZqAHjum92FvRtksZI
21FSRBWEfJ4mzuQ2Jz9oYs6A/Ry2ND8D228LUZ8ZSjuR5loGxOajj8m6Hy4XBmBw
Z6nSH0EdFHAejj7Jzc2kiz0v4OvcRUD0QHS8guueyFGOS1qh3oQbgFFUIMYfPZ52
Wr4PB1zKacWuKF9ylYZOSp7zHxJCsx6Ofbq+y39ldGcwVpP37xxb7SusSRi9wJUn
iOWeEUBOrE/yMJCI9b19s1Dl2Fc/narC9v1gkjeCZAJgSJ33M7T1Q4aNuzbzd/Nl
9s8vqnBxROVjm98ihvMLXq3HnJPB3HH7gCjFBdPczplZU6SKaHvSC1Sq5jFSkF3C
EgDn0Wc1IsywVTQDmjfsPmJKDBVKyOrcxMRhthwR/W1mQxn6y/b2d50R/pKQ8ii+
ylNLcgWXX76xiclsrej5jnrpb9ycCgnHfMJKcHoFyY4v7DTnjGGBrvomDKHPCGwo
wmFAr9NN362skQbqvE3QfQWrR4YDIf4KpjxVJedTqxCm5533x+Ey94r4RSKxZvlX
LWzN4Q3rPjdXGxioZElgQaACvUMmdVyybZ7JsN8EOnXFv8kzYIDBUuax+jmrRxje
91mp9KGYmp1X33dMNlZAa2tDGBr4SxOrxxoDZTzPdsSQafZun26duaOCQ5nBJ/B4
4hKp9OGVljX2bFPRBDooJ/I1zEjZ7G/To+r7iHvNZDgk6iI4OqLPsr+dd/O6NtJ3
lvY/LfiNhvhPc3kg6x4+WJNFPZQB2fBAC25T7fFeP3fJLacnDmvM0i6T4qlLjCSk
0BwHLPAf3vKc2EdunIJvdiClNFxy5E+HuLR7d9oA3IATxA1Z6gpyUvcOkUs1ZiKF
hJWgXzKLcZj9Wqkx5klS0IRFGGqTnptE2oqFPu/g3HQS1WD+BrFkxiiJ7mDJ54xT
TICxcjra7DU1GC1LVfywAy/vtwU/wjL1wisPsZOk5Loi5WWa/KpmvXw//DBLZ1Fc
ThmG8/tz0OAH4XQ7SpkXx0lYoN7d3OL1PHwMf+GW/Ofj2+cSL2icy6zcGjNHk87W
NPauBe3JSwgyrgKqHTGpJhwP/jcr3eSe8M8Lg37RF28iwGt4yBPAQffEi+bWKMUF
jCo7g2lKnjTUZp/4xOxiHGlgpX3wKM8K2SREEkso/pnu4XYQ6j+KpjXSegnJYRGy
YXnVnjlir9WYsth890T0JIqVJMxhbLPCoO9CJMwxOlNBDFyF4xos9T5xOV2yAKXw
RFBVJ2Z5tv+devIBPFCsogJAbkXRO8i6MimBgmqUWTYIwuZ7hghTDy6me0nKlEbY
nChRvgoXeGcivneyG4Bw6DHiIH16lPWJjVwore6PLxJsBlSN58CTHu7/I4OQHZUK
JAEmgoSjPhpwWbBqlBTap/xmngXXLXMHFOkfC1eQVa4qHh+D6BMb9SXQnu4Jucou
isqVmi3GppXwiOHiWjQy2BwQ18N3nE+noRGxLS9mI1ZKZOyR+a33x8SCXyDlch0z
NfZT9MlDoOkZ4VbW4wB3qsJ+iLcYiWKOVMp8weiDSjJKcKz67ew5SKvZhgqvbKpp
WubFurD308IcGBoNm1rNz6Hz627OvvBXmZTr6HXqsenfC1NTFw8fnHs1KbXClSPL
6vAiLbY2oQcq/PXDPIqypLQoW1VWq5seLGuFCA2J4QnTlEno1972zyWhcJVDrdlM
r6HUiHevDjUonPX9SY9Rl4y02r14bQmBYOCOU9G4XHL5S/p1HFntZ3P8XiaT99bK
K8RUAaoHXZrFmjePnJKD7lPFb8ZROxZJVxWtJEKuZywvtWxFLpK/ZbReg4tw2dcd
9sx+JoESricqIT+bm3rzT3ozGqIkh78/kFPx+jJNjPGqUbphbV9IVfik/Mo/3fNq
L7lYjpZJjFPr/q8cWAu1LHqN1wC1Y5BRzvEqcsrHzg6eo0kOq4FvdSQZM18g1cte
RQnPSVYBhBfS6wCJbCYfZ1fFeXTuRHJPARfmUxX2se5KvGiqUTNCdo8+TZ5lGj7P
qaqkKMFWpB1zQXpEzC4M//VFljJyR13gcV9y+oMAiX/KN2RVnml1erI6kl48F/S6
w8RjIHDnob7rKiOXkuECrtbzRJrW8CyecXIIXTybtoUsEAm0K4juNJbXcpnaoIkN
6zGrHZyYLOtA1C/jVuSM3ubv2apXKlyBICPBoCy22XZY5HREXeSgz/iX11MPkiIm
myxLdQGvhMag5Bd9IodRzsflRW+1r+rLQgLErW4HyCO8Ohabb+6l3iuKUQi+NYcU
I7pwNZAth34iDb0Xtu1MWBcgBPqG+WScnytgq5TxlOkDKU5kIh7Aze6ZZl40b0x4
m+1fnq1WNEYbQV4xRtKBwr9abRrd1VBmwrlvSSBrfbrJykvDyhy7IGAcAnqHjXOL
LwdHDDDHTHb4/XxpAoAk2oVcZmXRl/pN34cZhhNJB84lCpxgHvvqSxD1qlwboP8f
sm7S8Cgff5WUSu0U19JvUHQDFnNuIIXAjFgiimXTbvmncMYrD2tWVcMv5vj0Q1S0
GMnvuDP8MAhnyCsz7TokuYeKqHUuDw7xTnk/JoQMy+DOL8QYiF1BKmaZ9LHdgeI/
Vn0dvGQn5t+T1DT9lkYTdYBXbHLxIhgErqKCLzbckDwOj6R29OkOURBo3NnFI3W1
gidwxEvwNOEkBmkhS5UQ0fV8thTHfONke67iGDZQ8iKaPF/0EZ76bsM5n0q7Dvma
cUTcu4fPTZTDFjPPPZKZrAZlOYh6m/Bjz1EIrbWudF8Hq1RxBLDjoSd7uwXVdGc9
4jdlFUuA0mE6uTK/ZHH5YhXwzIUDRNqM8CE8UVDDdskBqWx7rJKnglOLZPTRQ8wW
HzULygwkD3yXS0NBcmdO5TMw43fa4jL+Is1YYJBeJ0rdTCrCXCgn16ZTMPjqilTS
OHqqVbBmIBFCsJmOIv8qu3WM+e61QhjzEEwy08IZkA8zQGvoj7J2b7+TnDGBEHRL
spz6EfhCbFcUbwqPtZHiNYobNgeYFWkFDjqiwbWAAmj8cpUGlpwvUJqTYSz/lKXj
pBHROvtQM/5bDQtzl9FhIzb2gBcWA3XBSjjKA57k+rqJipoRBejrK9gDPdy1muYA
g365LjwbYVxIPvUHK4L+c+1o0LAAbqH1oeIX2dFbj/2YKKz5tcFhVSUBqMJU8Tzd
4/jya0yxRe8l+QYKRWtp6pDo1KWboYWY1AQOJdnJT4/XYOrXXPEicBsuRg7Nl+Ss
ABLRMhJfUcUFzpjvx0akeGy348J8VxYJnpuMwt1XxWtom7cxE+6GAGFz1B5QtyC6
IusqN3Giif8b04fH5LTcNpPlV1hZyilqPCEnemnIq2B2J/HL10yqwqY2eHabNwcv
trJk6qkuSj9SdMQNb6kFGQxdVd1yBdt66gK+m/53JaxWxmmFlQeZIzJ3ezqC/ELR
YTJqRfwOF3QmKCclz1QcXJtpguMuYoJtTBZYoukL567qi4lWeZVb8xgMk+/bbhHc
Lq6dsL3ktgnwOSMj5K6LgGjiDMBn/whixAugNK10q4HTNhFBnB+hxA3EcPB9Dqsv
rhfMH6lYFIMwsifFeWvfgIWHqM37cMRnOVRtiETq2qrwi4bUFF6lXM4XNqYzsZas
NBJ6j3J/WDNa7m9BZShPS1Hv5PdBSiAzv+O2sRrzo8QDSX02iVamSzo3UBfPfFqz
rOrtznlRLtrLlSoBgHh8yhOet18PJcSi5mU7skM8YIVKHzdQAFPb+aKD+3bXJFE5
0UQ6XL9IzUQlrDCP3xPrwpnUqP0QA/gWDsN6ptr/oaRiI3gsW+N3FQnVqLQVyL22
PY2M9ff2FS/5c7/dkcWsVogZWY6HuwTil74DXlvxWWAZXVz6od6qduRx37s0DSsY
8zlL1qdkv9JqoHdUOLFU6/YhdcqRtUO68j1QdKGT6SSvWdY3vdO/zt+udUaFPFFL
evFJYnG2EQ+QGSrAJgALEYP9VA7Y4w/ctcz9WBD6OmuEu+73bqJc91AHoJ3NbiO+
y+B8muuy+F9bNiZv5CyTEVQM1MsNwXdJEgDnjlhHey/qKP8w+ORZ7299DWkCawVb
WTyC5WuzyegscWZq8EtgSfPtZj4tX4QaJ69YjgUri2COx7YKKRussczk1VpFK+Q8
ioGGiYNVKGVP1VQ0OulNSblbkf9Ol86xtpE3vwN2RghrSpwRvcJ6eo/wUW85pv5k
NT1i8zbXEPTQnhVZ4zax9v9HwByNV6LZ/bBE0eXwdRAMWsw2kB6Ovy8LLyK2h0As
z5H/7M8b0vOEu2J2Q2gOP6fy3tBOtAtQx5nUxIg86Nk236WY3E7hhIZNnk1nxtw4
ISPNjWB5bNXZNxC9zDKpIuOpGhcW+Us1Zt0HKG5IzwKBmkDxOalmRVXmlif27ILZ
QukdBZeSNgHmxzRAObgCX+CrrmPT+lLjU79Z6MLJi3N3BHCyv9HbVsa1ZctGKKR6
1/Lj8e7G2451CHo1nPfGqeBV2lNj2M3jMHo4oIomcpESJbHpOFDqv5Gj6BG9qZFX
YhjXu/Z5OacFTCPWF+5sGZWZI4/21MptUSq5oguTQkah+fFhlMWwLVID57bDxL5b
vLw57YdcEGy2cco3kqU66yDik1neQ/qX7EYxGl/U9hmoZqwUj+YQyBMhwcb6bNnD
tT4lAuJgYNteDeCkNv9XHLPUM0KA5jxn8t1+P4MpV7YLU1gE3rHrTJRf0FqnCjdp
GIzq+QKt11Tro53s8yPx1hxEcwDAFSO7Qe20XhT5fyE2ZUa61EqdpBDaKzMvekJt
kNkTqq2mb+bKFQxi2al+zkUJcYjakcElpa/OnATZKsTpD1yqSbXzSOtd+hH9VPIr
S3+9kAcKoLQBHnJiZTHfV82ll21+XmbUP0KPDNUyxnp3PyycuvDDYK66SaNLhmck
c2mYCU6cHeeHDYfFga9WCYKAHyn43gANzikmkAITDCnm5avFhiPm2U1asUf6Fme/
7nCGgniEndtXQIz6ZECom6cftsmi+jPduWeEB/FpqiE/JaZsHmUr+QkeMlPeeW3z
Mp5QK8PDeZcyjpgxqEp7CFMnZ8kTG3FpEMZHSPB6Awqt5SGMVzdHCfTKEAOqQvmb
b2RHm4b4H9K7LgZefDnuPc6mo+UQkvAvUskW5TGVZ0G0QuHRhml31cFnudK2wNTw
f+u7ftYgjZsHbz1VbmUDEKMAPZgS0UT9C6gRKjH1zN8zEn41H6r1Fyuk5W9w4vTP
h4jSinaMEWDoNY2b6o/YThnpXRcvTe38y+n4gNc80s0Bs4tWeNPN6cBNa0OwdWkE
vQvICzFKm6GGyAW6O1s7DA41P8nQgWt1XsLRp3ZBqpvSUnxE2INqz7d4OBkyuvc1
Br7FmVKo9hvKaLi4qFHAtrpPqb2AOtcZ96kvWylflX/Isj6GTjjX8TT4cWysxbAK
t5M5O+lAsUVx00p4bNCgj1mBrrQbqj6Q5/sB02rP7goSeO3hCASiIN4a8QgGCRu3
OiOOUqiuXHDpOVr+Ux2SHiSn/TXvLVgiwK+/M7HlH1X/ATcGTM7t75yGd+l1YcIQ
0Qzz1nrRu03n2b2JarF7NrLGJGa1qwab0z1yIZ+1vbf2pBPZ82lTtqiqhS3njxOs
eGw5zjSRzSDwQkc2hkwqYbkyP1pzekFWBGP2zOMK6eY4hFLd/O9k0FAb4FsfGmUO
6gnek7OPK6vh1wsoFCcgobcSfvV+/5yoL7VIQXWG3MsHmG5lk7fMkv1M8pTbzCUI
jPyjUINRGCRZ8mFMa462MpnOyqwrz0KC0h/Gh7s2mkz1sZeH8JU30fOKaVu9XwQD
skUEXb//pm1lxmwL8P9pYAqgQmpF4yYxW0n4+lYHJEvG9nL+WNtG/4DGy//rBqPD
9/ZXhNo/9L3dbetcDS4XdVk2o0mgTK496SNHu5H6Z8bArvXySaeQqIUrjA2lNMWB
lCNp5MckHHEBOPh7WoOWOkeesFhYXK0+6fwzBV5Q8CxovTty/fmwxFYaY+TTHqzl
Aro6wHpR6G9cv9ct8ZTtwf4DuG+lLEhenbbrrUhUL1F+S7dcSrwJaPWyYaW4WGI7
45ctctzL+YMyBxP8/iMePLZr863aJDBk/AD+CG35GarT4XjWizJI3QttAEw0amQ5
diQlC/ZR7A3rXfFGq6YGL7xw1ZuhHF2c3YzvcepgB6kdeRiNdpjmDSnRaAppGgKy
q2GZF44mA7UEmj1XiFFnP21HN1CW66ft6VR3Lu/aHKPxGBnBWttFmCBsudqwkaVt
hyubx79UefRAKac54OKk+t3YHmrCXA+iAAJK8NdVXod8AwoRDcFjv919u00EqUYO
BiPgvb5XnhkxuTIFowYeXBJZQorvWGjLBywIGaR0GeBq23x2UOoiCk+0mvnd+fPF
xX34a/YITTqYl+OGaqFCB4uovSxoyuW5vcCAv05uEDa9i9i/n/vBFWktAAI94i8N
2rC4T7v9JMJv7YY61J0DBpqYZUCL0wUn2mjrWjJ0TW/5db8Vr9z4QKgIl6SO9x1j
zSDFCx8ILbNmyTIN1ht0TF8Gn2UuHye54jk8/GZ3lKzCJteJZC79usP8i25RjR+U
tOOHihGAHi0npu19eZF+j4R+ZNmoWlD4IEHC/25L5ahzkSNdf8FysUat/3KQEHaz
4o5XuAub2bkP0PJbYJHmW0jF9Qap1naGjpxmoCJKpc74y87vy5V1UneIN9+9/OqN
vJNtZ/mXVweCjU9dUJ7Q7PKh96za7aY+ARJ6peTRz/lqenJSBxuJfhfi3Wksqc+y
2Ok/jmUI+Go6j/GREtHHVP/7RHsSZblIp/aP8IcSY2ZGujIEdp5TgECaqfw5cCjV
P5bPBKm+NPdRVMeFw7jzKRxt+DtKBDcrJyEpMsZcMlmNqrw33769ZKC4NTKECRDh
iNgBhaWLE4846HpF0nfbzG7eRa/47RpuDUrzxvBcrwqzTVS4fMxGR4MgyZRQ3ipr
1u7HnuYVol/+lhHwCTkJEO1+g8zo1EZU5LGHEuzpGRqJ9Pwt/xhuBtHTedRxngxJ
eNprwxlGhjqpYW6N7L9+n9+PagFG7s2bS2efkDjMG3SNSrTIl1h5fmM3ymSCLIge
VGv5274Mnf/30jEscuxMt46Vw/FfsPCnp8s2BeK3xDT3wPrJyrYUkBCI28DRzuaQ
f8tGJivQIUZZaTBxI5QYj0oo2d8PSUef5tblFdZpQ08HyeHtr/3VTA8MhHCNnmDD
a8uXPyl920v9F6WswME5KR8h6wCdQEJr3wHvsuNuRim2tCINSFM9MDVWYDLoerMs
7pSZ4Vt3g4TPIID84/vQ8rPBUDglljD5nuOEr4PwTLitERzxwO+Tg4DtxfhZROF6
mebnT5LA9nXlCR++1a5l9KExQxpfCFW78pGuhwkdM1qYH9uS0Upf22YtuaOlHz0P
BWMVNUarLqajP07IWXUvtalTVKMXhXtaD/6xtNDGn0avTK5UD6sVC6UeqbCpa7Da
ULsi08zJnv5QvxW6sd9d1uKM8Z4jjB69tBug23/H9V5iI+2tlaGeQds4qk3YXvLh
zFIjvX3kjzv6O+Q3SXs8ASXGtXUXp5FKP1BVw7RHjxpItmNT+KqFGR5h0tX4BqAo
FdX7OXfiwbsHQWo8a/N+/Kk1RVOwwWZQaD8++aaneQyIvOkMYTnmJwCPsa+JHW/h
2gScUnYN0GgXEhj/aZpLIUig32fXEKYGj5DEyn0EAco5sFmBxt3BMNcLmcKIrH8r
EYVzd9HpF0qjTpotSCNdDNDWRMqXdQKi3YWfBG0wYO/ySH828ppeYi40I4LsMyMW
8znl2HOAMmlxkn6zZS8Uw6+ijOb/c35o5MBxpnAnEV1et4fi+o9WahTrqZrrJkB2
U+AOknFciRl/5PHdoKiiC2CT1nal8OBMepu1vSaI8NX8UnbZotS1bSY9GvdTutNm
jt7pom8r70+M3RUfTbVfQ7zYUjeis/+NPZlzX/uKE29TcCei9LV60dAtHjaBBCk8
GLPBy1KqFTlVID/1OPMERj+ZXbQPR8OAR1h/RIf+1nJ4xL1FuqL7K20Y9knsPLNG
cNmwQOgbb/JLBJcgGxGd9u9zniOOKK7U8/VrPBuJleHv/0apzMhnu13ZvntDUUD9
rstkFdLj/dDq+SgwtrsdZwboN6MpV2rIFMAoL5JA1IdgBNf5mRT2+H7sKmJyjfb9
mbBmDppxLed2uqtN8lZzaBIwMMTLWef0nKoeqtwfn/gt8GZZJ7KbUZxBvwPJ1w1r
kOxMkmIY82NdBv+xfSzwYUyI8HOYySWcjN8+qKwNl+a3+dqIF2lux1PJ7gh6rL7N
ZRrKNvuzJXSnF4Rux3sGo5hpZzn5hJfapu54LsynCZ8w1OMX7iTff4yY7I8QjGv5
F/+SRw7ht3zpqPFkUfYa4Io+Ad+ZV8siwoUKmcxQm7H4Om/mMdAGXlJmB/yXUB3l
BzlJqbQBhmL8sPlRfvtONspq/8YJa1IvDc3IDCIloJZ6p48CekKJ/E/tF8Iox2fR
scEboOxkle6DF6hjkb8yqdKPWSBPlsURTawtzP0RTQag7bNWb/UJGEoIpqsdIc/j
BAiE/hiN03PfTapvURcPh+CLO+FbiOGYHbW2o5vFzn+U84cTfWjSi4b5lWokVQiE
PqXmyfF5YUyFHTa90AxwgOdmMyfNDqsQtDAO/LHk2Lf5Ylth30onuFeiJRroMwEn
aOXjFZN/YHyt9xPgzABB8bX4BMr4GGr/WshDvjCFXLcV61nrZYCV2vbl3Ch2f6+9
qkZxG1M7R/TemKGcex8iqbKNiZmLi+lSCWJKriOxHyPqX+t8ADKuYtPW06pRu5EG
Lhog6nu+AyG4nju/1GnZvqPV0np5fNM1Kn/m9iFTTVGFpr/wXo0KLD5za0Kwsiro
T1lrtM/1QzWzJEkG+TTJtRaENGKDckv6FoeIVNw12+vsDvND6i1bi3t2GXb4/FVS
0b4MBRu+vrD4birTEigld1+7tqiFTPRxPpkrp7Gr1s73pSw/2+kYdgNw/Crsr92K
SsaVhUTvLWBqp4YBzUgiDVl0qJUnU8JVARBCek8EVbk+xXBfrKGzzj5KE2FxqqKN
rAVUBziEqWilC0xqjRX7nRe9M9JuHl5AwCWUBhCM207QtheUeo+fFtB1S2s7A3dU
xLEWwRaCBkDPWrya0UBBUWfn+I3eZa6Uq1K9S5roNM9iUNBl/jRWc85t6zF8VwNq
rUG3jzGOc2ZhrEP8lRMZct96dhbj4aQ1k5WUKSm1zgNnIDd1rx8iF5Y+y9+aN51I
Efn/bV5A480GBgH/gjUx+O7w/Ma3ku/QpIrnb9c52jb/VlyAp0c8HDvWsLEaOv2N
mqiEiThlJvdPKxQN5AcSAoFuMXM0K3ptA7Xc5F6PhV+ZsTKhtHALpaYVH5ajdCfm
b7aPaP3kocPKz1uaAN7EL/3F54jmternswlyBlcNMRal6pouu46I7PsEUMYAN8DZ
YaenU1d31IV2csEnuGYm4newBVgdNcwYnrM0nEKEkIfb3iAAShtcEOawpQ0bR56b
FOvOEHOCHYesuub1jaHCBtP++amCcPzMTkBJcSK9Felvx/CfEpaZdbmM7TtKtQfI
JmOeTzCwUDh/6pzUct8+DdsWbbkzhrAZqpno6gv0Q7dP2Yx2h3utvm9IdtZSJcPi
yMnGdwXai4jKM10bQ2kDPCLX/DjL/Sg/uHpgyrcX0e/rcI+mDOv/iaOwKy5VMHBC
FqF433YPrVmrz7p3/GoxdbGUH1cMfoIcQAOFXHLhYVc+Zndf/GoLoaw+xpfItO3s
DTMOYIg4wuTJifK8J6KYJcKtaxgdYD8Ag1DUlljEO2xXdtop4dqkVD+vlo82GzWh
2dri/P4vDQweLkz7SkgfDJXRTFk5d2mp+mCT5RvY8qnazN6mOsrM0o3kNcydHRau
LNiccM2h7wEOshe4eLNNOoaBockpQQ0FRpRcpvtk+rY846l9BPSwyLqYHLt/5w2v
6SH/lj2jJECX2ITB6nsbt3eCTFJbMfX47OeCHmN7ClhCY9NVagjBjIt9xBWoPlSa
xNPegKK1Yc8y/WgwkSMtz/DT3i9XZNNpfjRV8cIEuE4FnsG8WieFR21XT8hDpyMA
LH639Xc6ymskJjXdw7ZeiBbygDpbt/ovlcdXjqDvTDDawKpJEetriXNX8ktx+/Oy
4mFJ9WjZ2YIc7QMakBkydSnR5DWTu1t2qHEm1jMtNBtimLaER4BCW4jHy/bdm5Qx
E8xfEwTaxM3qqZy/mZQCK6CFvaqSp88aO72ffWu35SZECzQ6zpcptx81d4jxSZAF
Rmdy0zhP/R44yxKnEOmNZXY7VeF0I+W2ia52C1I9mix0VbKETBhKmHCgPx7wGxk9
9B+uBgEWqInleGRO/t/orKDlBDorkYsULU5nrHnpFDBKuGPBWRMIB4ctTU/daCbY
vrM2FYhm52IUsZWGu92ychz5ay8ncaOgU9+bMfUCWgZ+n7T4jA9KI0iBktGkdBCd
nUquaVmLCZeZW0LWaAIcLaj9TLy7cxzPMytELxQmuOS5Yele1CF1axnu1ZxKo4UZ
kGuvmAh8in5DsrhMIf9j698tKzRmKTQcEPR+AF/3NB7euafFtu8fBmpxUvsI1WQB
Ftx2wiByhxPV4vvZejAT5ZB2Ji6kEOBZkOS4SZmtLzD75zcvAQGX2Mr8x4aNr3oH
0Wq/v2i8izCPWgHG2ZcNbOEVTuwz1F8RLWAYspCDQRT+BanPmVp0S+kDhSNMf0uF
pi5/BZUff0lAdcQmkTD1As43pFhg46U6CKH8AIKs4jvgJ+/5DEq/uPRCBrGjZJjr
Wun/7CmHBCz+3Pd0OoqVj/EPQH2ZY5JEkiw+0JYyd+c4UBkrukdK0Kge9rHSH55a
iAzCOYJM33f0DFlH/QbyfATiOnIkooNYb2HDpZizCysrRxS3aFwCbGYH+DB36VC7
3i291iWc3MXsU1VGZ96Bsk/rmwsiRughIM4F0SGFPIDIrLI3IRqqowv0YnQc8PMI
Xr82kyrdgwdLwM3mXd+rlXRyuVmFdQ6Qk/b3h0SbR8jGtVR6kP49PeHgXMuMrZjH
ah9q9wtiOCBupeUswXZFm3oCvi8S5xMcjaplNjIPdT5fRyleeuOW9I1O74BXd6Mj
2CezorL4lKdVr5h5dpuNLeC3MgkQJdGihFs/IXdCQhFRTjMeMVIuyvlGutsuUA08
Q+mSq/Cbrq6RiyGZzxzU6G2NgZoWOBVJ0SiNJdX7emy4kq/UDIq74dpmqD4d88Hg
rfYBWAl2DgdWBi6URX7ve/ih9F8jpYV0WStiIBqU6CojPuwER4EfrnHzcG7FN44R
sU68jde7X81HL066uY6kRRTNGn4KvrGiudK868DN3juRMkI5JnOS+SmC6eyPNd0r
JG2jTgWH/av0o9q77SAlIUWY+NuyXAb7X3RQT5CO6Va1rCN0Q4PMASmmy9LZt+LS
IBsEu3yTBeiGLqXGnm9kHUdYM25bOvLO0ks0/8VVuJDXm1592HxNYlQfvj15bpGl
onWKf6RLu+gwmBrt9GYTfJeYJ2324+tILe9AA/oQfdj1p2yxknK2ZoZRnF9pDIc6
hl4vmO/mdJsiyL6PUHHhcVYAUhguDV1PYyy189trPidUBHZTSkJCe7ygw0Do2YyG
VC3sFGWsF4RzbP8YkmwQY6C1QybSgyR0dLqCexSXIApO/5eqfBwfGIV3/vh+oQTO
lL0+kLrKE6QrbL7dE6BlanxQI5Na5EEihiDA0UEYHbqw/p1chctiA48gSLY0xSbb
vqUkIdiLToYSUDIP3ZlADF/hjNkf1hd2NoQHnvgLEVQ1pCm+HoZ+DK7FrXGTqLX+
/pmk41tm21iabRTO4VvsHNgOdzUxOzumxHiXeOJ7/fUiHzn26k63mr86mMJnT85L
UmaOklTG/fjCXdhoEigBZQVBz3CqHsBP36OEPkPq2o3L9dS48a6XJaTeY4HXdZzd
gp0Xt6XYNpDmOIbWaughLgjWF7yPlsiI6jT8ULCw4VXjBR51GJ1cI6Utm0JqSazO
leUySPt2HTfyeMSONtbOvwpDisoVAMz9zJaGf6oOPMreTogK63EivZwXtqCWpPh8
c3Uv0E4QUZM86hZ+Yo60dPJWhSHuIDBY0t5gmNyJbKo3U4F/JajK3sSZSrJuB7UP
oxRILA+ATJCHC4tAKRtva8AW6nRJ7P0vG0H/7mcubG8mEiHQxRit2Wb7SoKHDMqd
IgJJJqhR3G0gcCJnBTBN4593PAY+Cd3dsYYpRfYLB/ejwPRpFTWau7ONW9Z60lNU
bk9qgywn4AXRHJZtrktxhbeRgdaXCEV98hyuFYHTiScpvnw+1TEGcXC7w64Ayev5
1XsK2VFsh1bjStfCHMdyT8RkoMKmyracTQjz8k3LXLK1GXJ7UJYATW4p8CpplN8H
YzJGzDLT1ef92zzHNvlmfQmyuPhshsu+sxRBui21h8n1iMKJ1fr4o0PECHLNBgDC
iGBm9OeP5MIOHUvWuZK8QOsdZGN28tzXX8Xg5MTCslssTwL3DkSFiwD38I1HouaR
tRKM53UvFIs5DDumcGuROYeayNLYtPnG7WjnLJ7S6QEqVelIz8/Jw+rUxkTpiNlo
jb2OeRDHdkRU2nDFNAGbqOgfSdrhlBTETtw/emsri39OWSLAfUTcwrqd2sQqbhUZ
LBIxtQbTIm3RLl5mNzmyEbwWEaJcRtNS9ihPA7xhSZJtjpaY9IErzrFK5VOeIhWB
3Ef1OtgRW4rdbH+Sd5EVfJRt8fw4ukkCUDm4kZZsBTlN3O5XIwVB7B62BZuvc7R5
HG5fH3VOBURrnKnN7UaddgATWLyvzdz5KvBimt2Ig0oWpF+ile/0fHu18Za7Hz5C
oar9CLiMPZmaVB5zCHiJCJaUueJKV16/9IKMzak0DkVjzxP2RbRHpTU/PWNNePZo
cEGHszmW+otmQjf6SGWOyeh7QdQ0etZ23KBuLMWZVIFEXPmmPKNjOWD+gb3yaeVU
RF4l4R9IzFgnl0h/9PReVdz8iZDtHE3tIO/3HCqtIL0iiRxgzJBt8GsrL8K+9YOv
fOumGmcv8c2ds28EpwGLCT1/orL/y9lPAtnq3fEsjlfG/uv1ObIYEcOy9sojUtEf
6zplyBg3oeoYt4hlimxxvCg8VBb/PisTIx3R8jPhnnmNHRsUaIobXbmaS8TnL939
VtFTdSxjkw7voEdzNtVnLTHyWf+Pl2C5h180MKDqvFeSbo6Syniu+aAbY7ineBR+
RteIkr+ySb01IFWSW8o0V5VvpAQWRX5xaAkgYo8GOXljW7PlYYpO7SDBtSQDvYZ6
lDv1GDSxKmpdBWnhmDYk8v2A2tjo8RI3IndBZeGXW46WO7D0h5mVYJQCy2Cj+kQH
pzVjW/8r6s6cqQxcIypk46W7ODgO4KP2Dfo5bZju0v81B/vxAwHDE9ez3kMhgaPa
iY17QB1Q4qfzrlDAnZl2DxMVUDYrlXMOCcEKRsq9j3tmDe92BH6yBFKYLHYDymgB
evsyatJx8KgaN35jOiRDbny6BdhybyN+PlCx/6Dmox65rYQ4M2d+XFjqWbQNArxV
xjV+/yvlxOPD14WUk7Vg9FHmJzb61o5eiLi8V1ue04cbwDP4dz1XY2ZAL57YPza1
qEygRNfuvX1S+oyVtmrY3gUeHU/zD7JfFF61hBpnM8dKEmMMqx1KuEsqrbKku4LI
s706prhltJfkxda61shsdDZnDkDiJ+gpnoe1WLUaN4MRtrYh9qAnS6ay2zY4Rn2g
efdyhUEELMFVokRYF7li+9Y5i6/9vM0H4M+UfF9guNwzvI/OrXDVDwtXGQjV3jgf
EY4x34C77GIqQNM1MSRYzKkis/W5jXzTkal5Ao5lFW123FP3fHu4w+V+WpQTCN2j
9OX6ho6y8R4lPhHCLFfiteBPxscJwtWfYLYWXa/YTzb0VCN2COOQN9UbbUg/iUJ4
HEO7o2IvBAJKaYTwKxzAxxuO2oaWLa0fxvVKrNBHvgPkwE154eP+xY682Oqj07tY
7jf/I1HyQebv2qq/AB3jm/Hs1PF/jZUuP43iD/KIwAfSHL3NiZ8XOppMwnukyy0p
oJ+P+OKu6aouwEvkiYJ348bQfOsuCjAGsF07KIpvyt/d6FbOdfge+aRCaNdV81ME
IXgT3ukAOpp63A3lHYb3DBV36OPPYgSOoik6H9iPsV/FzeZ/RTZaNV9N5AvufMdA
Puf6y0JznxdwLlbwGdPP3kzN17FyFBrSLKalI8N3M+ysIUO0Q2ufx5J826kbPEyn
BVofOofJOtQjwfkHbz4ZeViaZLAHUIugyeNOvnI4l+D9QozMyvWVlOCm4qFYsK5P
y6Nj/S4sJx33cQpxN9owGMC3SnbwkYBtHGjZZ49XhjM=
`pragma protect end_protected
