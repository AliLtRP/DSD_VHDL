// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Fh8zZDh5kg+FmWgec8Vi9QeMadvHNjHuQC547XU97M8ifYLIJgvxZtfQuX+SbqjvVo65d+ZcPX5v
IrAqveKGORqEwJzw3ieu93MNiRJTSY+w7HefIOj9WzYyl9WA+AkIfNQTagXiw8yXTAANf3yEgywi
17Owh+Zfq2ysWIpVGp5cHeyP/C38AyK/JWSRNCkCyUHYI6MkIs2dj+CMsHGDnESE1b8ySX9ycNyA
KjkYH82hPiWzsE9poB4ZwMc07KX/zN9yJXK/RdFs36TjO0zsvDNkT86rQZq8STZqUDscIXrAmlnA
kDmlV5p+GSViUslEgeoP9ofxJ5lfw47d5Zui4w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
rE1Qh+kzsJoFJfAeekt44OcsiLN8puetTP07+Wa+YcFoNrrDirwhCd4v0PJ4Yk7K/C2Pk0c+7hod
pFn+8Ji/mmupjwWXuAqYKoPs6lEwIfaDYeuAcCp4kS1AtD8c8PH8HWaq8L/8GWTQo0RLy9eBKElj
rGHYBd6aH+OVSZxndHC1IDASVa0YbZk72CHqdXrXNzk6ELwfY82GUrlGSJ0z3wRA1Hx4sN/e89X7
kw8f7EG01kFA4/x3E1foRddg37TN9Uncp4fEZ6l4pO2Na2fITa4SGqa3WYEKUGdtTD/EUbRmydMb
Pzid4kMQizhcjJCfkvmdF4jrpUg5NZG26NQb8v9J09H2OE+Y2uen1cD11ldasGtDTY1IEefjivsS
b2NDt+Cff48dJPSAmZaEw2I8o4Tsr22ceyFNL6tx8cQ9Yl1bh5PcxuvlI7ect5azbKuZYTGZk6Ks
ALvXsK/P15VNs/28MZwsStoWZNJTTKZ0ehBehw/z+M3spSH5JOlTp7qfNy+ReV10roDtJ2v6f+3M
tiWXR041h0aiBNrxL2+kLY5rfaGM/f/qi/FDk5SsG0x5qGuR7YFjyhaT5OVFNn10I6ng32fGdix/
lur2gUThaujEi4HpjuQVeyDu4BHMIEBtSA1NdODGOuasZXHc1drA7/YN7YCMq0ivA6O46dveabLs
65JE2hWRqSrHNBwDIjZZzDfYKOSFUcDTs6hbxLaxejU3RKdqKTVrlfOLmwXq3Trd46sk59+e0Gku
hDh1IyPCt1PgYxh86YlcyoKFX4J04kyj7BgwualUGn9gfA8TvH5kMkUidjxy/nmhGjaZTqp9Y4GM
TQ+sYZTI0aLNOgVazuBPwB181vsbhb34EhClmv0y+3X72yI03pZ7ZN/AGk95rC346Zk28WJBOm+f
t6mEEtznINk6aG0SHFD1fa4bE3Fal8uJ2T9VeQt3qGFaFKSeDAzUwGuhRBCjuWAlc1LefqmYz6z+
sAW3nvevEMuqPEFWnZwgwhPm2VKHwjYIfr8AXiCxY3kQ0V6x0saNg+E+kJU/WpS5GzGFSJFNV3rr
tqmxHfASB9w9H0SX3aHi1gbdSLPYBwdwvCG2tB6cNp67SAkrnOcGWtM8hI+KbBPs3ILWbbH8lO6c
rN7tSJ193/BSF8Y9ynx1uXcDmBXvZGLcIU/FzLAweWitNBKvxBjrBc7c5sdFyaOgY6CONGJF7OqQ
6yeY5kfNGwP525YTxW2G+i7mVudzsotjaS3ycDNcMYD3VzLhmqXpBShO/NYJAgrCMF+h9ZymzcCv
zReOlleZ2B0HbkZCRoYAVAk0yi9Xze6yNFODwCy+qpb1Gj84zNVuVs+senwOuqtogXn0dRkq1N7e
h9EMSs2AMR6AElQpDNWSATvt4/SFooxry8pW7+HGxCc0Nn2stSFqpQawlVpr2imq0bzYsOPVWtxU
whAWBz03RwQ/vzW0PKxfRceYsUiDICrRfQhAv47V0EwEDOT2T344mYum94h5I4nrHps9/WeWDMeF
krfrrF2VG5zdMjBWD1oqbQXW3NVxnAjUMQE0rcms6pLZXFZ2AwdSzt8T0qc6s1hfTbRf8SsxrH/4
qZsXuvuA30edlmk11HkOsOFCmoX/PC38ACfi5b57mEUe3TOS+8ei3E2YDk92YbCQWjHd35vLXqYF
v+kWyM3mMfSCa7oZTOWDXWS1utVsZn/BwkzhkMkJD1J85ZorB+RpXnU+tgVoe8lI+UsXlI3LXRNJ
mVbc5eJ1NcHczKf1wORJNeDHYESlrH2QlXIeG6X/20OKeEE1KvRGq7uuWhSavWpUfLGCbJM8lLZ0
ZvITcVpmFiib57u3ROGOPC4HNSanarwwWOlb6q5TnAuFmhwnBneEaN86t5njrTQDrujI3VFl3qea
ToFRh2UIlGFeM27SR2sT1dG6okJYzbI8WN5A2kVttjxkrmJRuMX3aHpBEfrH1vJrZmBQxDpP251w
XRgw3d1+rydt11TioMeaE6ww38tV7dKFV40RI1SLmQMDcVDUAqUvR1dzB+Ln2O67U480qfrDBh9+
/r2NVmP8pdD5GdaRuEjlPSUSRCzm1IqdxnnqiklatmWFZvmzpcqJrH8hl+gN26dZokoHvRlSPjRo
UIUJuDlf1Sq4vtn7TSnmBS9v56FMXQmqtiEKyZrVg6VxxOw1nNcl5jjHsucJaEgXlBZTs+/1ouVi
h43Eano2Lyqx7qcVabV/PB0TOJr5OAlvfS40c6mqVHHSXtikarSh9xf/gt1AB+nmKzF+qEIWoJ0+
gRrTrQoktSOA8nbA4bcGehTErIfYrdVH5GY5WCPcHM/Niq3jC24CSLl/dBkg6UD5V+BIP3DMLcjz
M0HfawBpUL3bjxRsrpBhR0HICehmoiblVvYJgYZn/Ik4GoQwCC6xyF1+lwV2uZKs+VV26vBPmwWz
3b/tFpOgrKAcI1G9CFiqEdhWanvgFXeC0zaewunTu2B+ReHA5DeH5hshIB2kqoUKF3/a8hIZTI4N
WcdRVIttdDNiZV2wYdOkIx3q3x1QDJbC35asISI3FxsvBpxPq10UMBR9neOA39WxEaf8OXRdorh9
SJmMJ8B0woSVc9rWTURFOg12ouKTpi2Tj2ctbedYLS6hzfpyCaXgN9WD6mGWsak99MuG7nWL+n4T
NFExMjv+Y6x4i/d6VRj0yeBAp58uGdNLtawS+M3yFIjAYe724FY3rFSILI1NRuiSEWIUD1hf+37n
UXPE55pvaa6WkXeTOxC1iQ2HlilFI1hnLXzlhSVXDwq7MtPQYCG6R96Z3tXLqHP5ELl2rP4HjoRh
MWjSurgKbfbVY2AXsYvNpjvs0lEkp36mK6Mrh2n8IhRtbAsek2Ec830JjSA5virCuoJc8/qkulN3
9YC2dFlHR9z8pdr2l16S/2L6+lfy2V9Kbo4+AoTQ4umhicRqsaQdXCcRAaB11Z/itdot8fpQS05r
zol1S42OTv0q+VkexuMJ93ZwWBB2KFzZfrUM3ZE8XYLZ
`pragma protect end_protected
