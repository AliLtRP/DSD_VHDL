// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eodQhfgVNyjmi0mpl9pXYGmUEtZxGAlXJmUPktynUar2/i5la5O/TgEaom9Wf4jc
GRhKwSBccGJvLGWgE26vLyJXS2a6XpMwvBaGsRpsf+jDj40HNtwC0UU+8CKlgsgV
BEy2rdVWsPFiIfQahcBL7/Z+HRJqzI48RcugCZ4ee8c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16960)
DNkfGBunr/VjM6BeLKqTj2BWW//zKakWQ4byaMxUar5ZyALC+hkW4+lDOIZoO17J
eoE9I+sQBg2gGxw1+0WE/wU8Y9vX/S6KIL0OEodxxYF00mnRbT+mfkOtWpPPSJIu
iQPsJPlaLv5NjjQOBCvcYlhuPJ7Mt1Kc5Oa6b5l7hHWnT8ajrbaB2rID7LkVG+Gu
QmgtnFkh87TBpSH3xmdbhE+IUHmc2WFAyNmAC43GC3DDsPoW12oxAs3CBu6bfZWZ
Uek0J9yTFGwRz5ru3zjzt+hx8NiC2xcDoY9FvCwjeG0XmU5fVkMgIVhF65bu01Ie
4h9fgCXcLB1yJD/ROd5V9Gx47y0z0AuBCsV9rkt9kGwCCoNIvncpKnbKgBWAttGU
nPB2GcmHRL0sB15QwUONvm5SldpQjiyahNdiMxKG9W17o7r1FMYonsvGhUus2VE4
/7+pFePF1tBxnyrxxlkfkACbgaftOyzG8hL/DZ2hp7fa06M84sgKHKU36nca5wjP
sS1Jl3LUEAEg/JGi135xdA0dw6fEvHngo/FJxN5RSvoUbncgLDQ22EMVag0Ov5SA
N6o5ZlH2NTECL8joE5h0uW5Gf0NK1/tRXm1QA0qwkPh9FhYc7NP09ucbwrsAM+Gj
uU6r+LVuFso9ZpKWHgNCQS07dHtdH3m9PkXAiFv6lGO4y5GdFlxT1gJIurRqT+F+
nA2wP0QwbBmxROhnLUhzD8m2Mk9kTmcYYo29gbTlxcqOJUVTgITpoAWDMqvzVA0j
LUU29gwKvBiq7tKnkfQGN2EI8AUy25r+a11GalxdWbGe8aNV5T4k92hP3SIlCEpT
g54zXNO0lkKs0hTMijsEpssvIZ7UGSBA4u5O1sx77q8Ls3n6xivqZSvlzcb2hbCo
o6Eh54b7he96TIQDdlmitcJ4h1ro5J0WL/FS9G7nkICdVj8kj2VW7nnpuSDam28+
K1Wfk7z7moEpDdSbvsDsxwd2F49OcHphURZExf5MjtzprJPcpXjGDv4CheYPeGsN
NBS7wTC5oe6peYfDsrZ+aPIXjVhAlWKA8vvmbQF6SoWx3fmeSn7EckxSEEqfc18e
JJJnpvtfDEiXVR+WJ/78gYkRLHZ1C9bzk8bbUtBOXrjp3u6as+qGaHTChuYGtY36
XZFFJYfR6/5cvDJkWpGfe2eiUCUD2MKd2vq4P4LCiQOEhY2bCdZgRpU0na4bUxs9
FWbC3GA/DSK0EOoAQe7DxDsWWxruyFFAyaLVZhyTia6APw5A5Lr4ML0r/hGUVEGT
NOCFCe09h7waci3fe5+MfbDm4TXoPRPN8ghxP+e14Ljq6Pq6aTB3BU0jlcYjNJ1F
t1PpQpmPVIXhCYyTbBPFERQk2BUvk5Y0UD3cUJjv+/6BIkfl+O9gYpJMsOrzKPJr
Zs3hrtA1NBKNygGG5jrRApYNyhW4Y3JGaoY2VJPU+hUrjzzrNNcs9MAsKCE5QLf2
LYj8FE3I16jT/2GwVsK58OceDZBmgvQAP7dFugqRbwqe23iTXwB44ubKE2CGLbeg
NA09ZSCqH+oidLF1lCuHW24UPXTuJsyhOnHOo/N27eJxDEukMjIhM7ggt1C12CL4
mMnMAiAx8iECnZZtW1im1lAsU321TjEzhFgBOcFwUewe1ecLE6DEm8VUO1aASUZj
yp6un9MtBKDRYeXlbdnG0BZsdkvub41xV77Zd96vwZFotYtvHhothnrv4HejfOZ0
a1707yUm3/Pbyb54OZ2/o1wijQYVUBtPZtigTv8eWT1oKPvPxh1HXAwn1Px58Pd0
9pOPaq0jGBuveuSRQRWDL4PxQ2JzG6GoZgMfHyj6XBCb2IMhFV2Ba62Jhl4kjiCI
nRwxF1wrlv+roYnYzPKnZt5qbmtl5sqhZD/iNxj13fr7FI9K4O7KRqIDGUX6ZXzh
G4Dv9cZvbBrpDpFNo8vhaRRv8zJ1vmaB9bo/VMVkjUQ2oI7QkQoB9gfyYdevXpOJ
WQOYjZpPFfGi4XklZylV8UZFmNhHGFK5zQb391xHbIRxB4FQmyJ/GQnz4mS2WYtj
XNAYhBCnTXNnH9rw3lXXnecQyoJf0uJjtVxXLDcnQekp8qrhlUNzDcJjrrnlF0+K
a39gpAinNLH+Cfmtz7lepoAthQ94quh0+aWa4wgjVLQCXv8RXaqwf44Iou3QRmwq
Zy78ICFh0Go/LeMwtrpZPO+yZ39MnWEaiUWpBOtt99pDy4NL+VvanXm+T2/eymbV
i1wuD1vq4ofgU2A4q20o2fSycAKbMq4mTOdH9hwUfFGOoXszunKgDh8OZdJYzPiA
IDOViQiYQJ5QcLO3vr/NYpLetdxHZAbmmM9MZ1euejM+lZngnGoYpukNUE8yI3LE
BbyUlm2OMmST58iqXQdq/hJWpa8CIfUR7z00K1wcWW0icAbs9j2gohV0g+sVNNH0
Q83amfNa2ApO/cAKC0+TNHOg/wr8bTkuj/hFXTbf+IEkgsWlQWs4LMrNuqxuOzET
U2g2pawdi2pUNWN8STSegMahG5r9kVu0JOf1xYRgFCGERGVtLlKxit1y2I0cllDY
4dmXmmecK+KmnbWvDCsxShbK/74v0XO22UHq2/08GpDdF8JYCTTH1fX98VxrIP35
Cd3vnZ3EKVd7wb8xceybjSub42SceoTvW6vEaoXqAtikpIiTZsYkDXdzqFt2o4kI
AMBl0eFkPktzpqk2erkDgEcvf2+p5zVlA+n6S7eEIY8j1UrO/paJIpGToyo4Ezil
4iCEaw3XrXLT8HfDc+WFNf53tvvu3adGXnv7PWG2vkkVE29lTQvR3a5WyqVRzlEc
gJdIWRFw2Zf+OpinWxMauKBFcb7syxNAFimCgnzQ255zLEFZlhQ/SlHg5/B+lnKI
joqjUZb3ejgnbt4FZu7hNC3ZdZDmgrylZV+YI8ICLsxCUC+9+gyZ+LBKpqA/7n1u
3oDK8A0C21GL3rZohrsKUUiMXY6gplCWy01kxMp4N7vbgQYfEoGrKz3CeZck9n6V
8DT1VAVu+ZJik4PaHZvPR5ipT/gOfme6CE/z+nF3DKLkZLxzdtRaklND/xSePpg+
FMiQ7Hx1aPGb8Nwp1jb9RNdcP9eGIPVXBnPQdEN3uOl/smPBhbi+x6faQsWeo2nK
BDikiXJijuWMdRm7vy7qmxVTOYXwgTQ0GCg6W3VEcv1BbmozjGt6TdEwtvO6ZiEr
ZFvIIQoT5dvfYVta+HcUFo/s43IsGPIpS6+pwTfZRhYr4Us35J5vzFCyXma/XHhf
W7Cd5ejZt4jkZThttBq1leq7TBK9iwCOuxSHdxh4Pj7K5oZHi4f2IZ6FAGiVZKRp
FJOUZLDc/xQSSNLL9k7AaPgwi4koqEWpEtAdZxRlaIyrnrfXuY5q+/qzCopnhBoZ
F1xDFJFIaR19foSjozBa6Z+cuPj5gCdhg+Le2A/s2zKGJenavMraSCZdEqHaaXjT
p+NUF6QSYYX3pJUlOKcsLP8gctnZ3ZEnf5r4QRidNGlXPGTtWA3xImfAM3Z3EHFg
xiL2e+nsL7Kf/z51OviyDkplNN1KvWNRkHKzPq87s2PELJ+HK5uZ/mNxqLiySwFk
AbSJoJVM9fukhq284N4N++uanYMaUPq/Z5k6ODdh8/TPHM1I3OayyVoJZQDYh7o8
kZkJwnxmMVJeiHj3JYBaR0L9rKpMxEa80OKroQS4RHhkIZCHHYHtr59CnR9BGJsV
xvhm5n7R17nQz7Usxeyz5J8WzY21I2bENWYC9NZnc1oe2PCJuNv7VH/DVq0xKkD/
oPl+aBp1Qw7B3w8eHLsYSt8ARH0Px39lgBT5xgxZ6XjVQvZbiCRMahXkaGeF+87f
UAbKzIShueMukM98X9/iXMfYzO9ta/4lsDPUokmS2w/oE2cXSsm1jisJN/LJjx2S
+6mdCe5/E+21xywR54GHtcw2U70l6WH51lWbGMHX6xIsbXs9lQalbpm1n/g6z/o5
dnYLmtyMEKI8oOAfCMmOLb0aQZFA6meZkjw+GZGuItMLoUzUtKf1CdjCpIx3gMk6
r0f+Mv/lqBRME7jAoxZV/cHz8sH2R2EovTBc+wlW+luJy0uC+xRBz6XTAWBqDVie
m/mLPF9sFR6fnCE9ex5LHvfxZACg2nWDGNMLjGbSxEtnaQhQ7GKhmtlyiAzNk1WO
yQ2TWDMaeh5GBKY8WOz0IFAQTHYCkDveB+EjxkekybW6PEbEkqd77LEYAgecKVXx
f993sem5aWjHPK/zzTl1cBi/wJ+0B5bMyN7z7i65/7Mgsv70E/X2Detwt9L/VDwx
GcETIDfBATwgYW+quOHOnBCwfGEsyp1kB9PJlflK2q/SzrzUhOXUZ1wS9GYMXgiX
zoJnz9aERxP7AUIDF7vM4fDE5yBW2z20SYOnkHkCPKb2w74HuogA50Ne7PqICwsc
p/Gd0cJ8EbnCrD/2Y5xewu1MDbdKCnSLj4jvfwP6E2MbpSj5wDsD8UlKC49irp2H
fJBmtLCfrwr+z3XUNFCScjozyF0cIHIxBD+U4oEfLM8ZxO0kNNhLhTZFvjBKM4IN
03dwUbH7Y6cDZFYitLP+AI5Ry0AXXE8LeBQyhvTzGkDT/RqOHJkCqdxK+VXqR5My
tE35vYAqVHPJJoTqHBVABXoENGDep/w4lLZTy917/+9W+jjRATip2iGq3zVwNhzi
46FFmHZhieo6u8gadgXQvgPm6vWgSvUSQpcO7OD2k9XQiQoZMDOPvRRHRXD9YHEj
dn1BjFX9fvEvz5IH2L1017dZjciQk2DgpXOov2aFKxrnIyFkP+7e5B6500kqgGho
4OZ4KQtBj0A9C1noe4YQLBBPXag2xcV1ALar+VOKU9jasKq5955Yt8w4Jviog8Zc
UJfSArL4UzB7hYLeItztescSBTvSuvEWg69UfeTXnSishj7+4eI24tpSeZ1zkNWK
M1ERcZeBerJ9R3Qk6VETkWeYFZQ6nIWuG2MwKAkrcM5+v2GFSAkWxp6OnJI29jfD
pgXVG64JRjVTkZnM4U7lWyDtQC1KdiBSBhdij+Wh1R5xEkDwGKo3XiL/v7Gcf7Ru
GHU/QyHsHmiljrbMtdL4PfDtspdG5tnPNbM4GdHa3nCqjhzptcN+kc0KSAxR7/GI
XMuuq+H/V0EMr7qiocispEYvgN4567iEuyd5itvKAQ8KpJ8IrTgJBmuLU6uzU7Sr
VrPV4zqZmo1Bb4jWaYodCGyYuHnbjMmoL2/vn0iqHusBj+HQ9vf1587UGclx3m7S
wSyxl3m7BnnF0YIekbIQlGoTpwok6jv4UZ7WEN7N2LXFRgE3Yr5dj85uCH41Ei7e
dJyIiFoGcYIoj/rA4ttjCmd385JVGf13+qEEi/mTJ+vOkXKav1vza0e/5EAfXkdC
3QzIiU+eIoNW442Wh6U9VbVhtPEQb5te6MjxBgVcxORlrsmraJrZH7RArjPPbu9N
kpMnQkRNrAjHUyfQpAsmh3D/NKkxgcA+JOCqK/otqtM1m4Wil/BLMwHmnVcQQHqZ
CKbvCY71b7UDrSU8kc2D3IcCR2jUMfEhK9y/kaLGd1hkor6OKTvXyKckUQ43qTl2
X/7Y2z/QVCZqD1Ny1NW1UOOgwA0MXb5uVINxKLzwXBZdJnMdefyfh3eUQueTiz/O
AAN0V91red+ES86BX7whTEMm5hMbgcRTpLwSHJDWgrTUazjdvfi6zinl2z6eHcpM
9Q6QpilEM5AyTrCC/uNAZoTIdr93GHlq86pbiql4FibyyEniexXMpV2uYhpdROop
kblaG5zRei+XjpLy8UMNI3EG781Q+qlnb26rmssX2us1WsJlUcTnlAqDlHjyeMGW
ywMJhTupfaKpwdT9QYLocmWVT8AEs2HKP2ZFGVESabyOdfW2XsjrSvD49Wm/bekh
96Qe6eK5fFWjdvZL0LPyju2YB5X0DUf3KY0Rr3cRuTA0sy7SdoK891sIv52UCB/m
aUuhWwnrs7P0E0bOYUy+KP9PfzIw8oBNGTrSAQLLtCl/Z2OfLJCY7B59kXhd4rv1
An8vxxljvawQyZjHsVYaTfd8cNpMRiwCsrww6sZnMAviHGuhDVXi+Rhs8S69rVms
jC+MfDzkcmvdUotwZHRXrmZwuqsyPLykp5FtXB9fcmyyuigyXvrpOTCEKFrX+PyK
+Iqg8WstIRQLyHFDwMVEqM4JbGHZungqK0/i82QIZE5Swi/nd5AhvC/okTC8szCB
2IReBAhI0KV9Hp7NBAQHFV+oWwgUwFvO57i9nyqNFlHpIQ/vV2aREHf0HGveNRfM
90qgk+wQ/izH8yxrz0Z3STKJPFSef0LAhSLmAPL53gMnRsJolCXT3uiX/DO54H0n
Sn0WlYhAMwHPCixC0TFizTRuphpMFC8VpOFiem1BYCZiRVqjk0GPsHPAjqjgzYAw
xgmEcj7jpj2n5gfV07//R/5JIslQ3Ls17b6s+jU04eVxtsnbPWY61iNKdkzjAl9V
G67bC4T2Rh2XswWQuFWakiIY5o48ap/8drf5isbLztj60N03QucaL52TJwb31OVk
3SwsuU1/Xio24cOMFRgwV/qK4UvBGytN63jIPrq9afnOVNem3AOAXegcR3Vn30AJ
VALh9+Pk6TFt1Sc7h9RS9FqES4+LI/hsfc9TgKjX3DcS8/67gdvu41Je291veJVF
zx9miIjxGKFTgqqBhU59R7PboSTZLOZSvm+4gAM1Saa9Fxp9R74Fko5MoEl7OmWK
BrMFws9pqh38LAbJQS6St+QA6SFm198hx1aZI7VnvBOfMWQ9CPDqvkfjy/uTAl3+
b2NpgoqQ1Sx4TBoiuThWFEDSIN6QRuXZy/UpQHFH77XTTZVRJ/pok5ARpHCznyhI
iViaTxoLnlzQ9KWl2oW7pxptuWZPRBeicOswjUj7Hj9J49KnsFP0+vmZAT4rWLsT
YOPuxpck3ry4WuasDh2/QLXggs1YMj+zh2ZlGf9QenKM7JmxxLDA9caCoZq4Y4Hw
ZgkKppT5PZnmnZ0S34N1iBaXTk1DMq0OU6EUDEViYlY7ogJF53N4L6mDb7pH/cL0
erG50zmHbl3YFqw+mYMTIk4fPuLEuQfM1VhT7VBMyTDPx5GWvcXCMeSJgVAE2v0H
qhGFSKRDARGNIT5FA083ykDkNRGL36aJm5hdhjNGCrUgcXPjBIXwGvkg5sjst68u
Esst5pAJoknOe8kVPNyvyKsqd7Zk0jQGetkiKDQ/3HeBqjcjLaTIWWOE5VGznM8t
fWVpd0bn/N+zvJH2GxYgtnGMvy9crm05X4nhXH2BTOJnIWSJz5QUTeb0izT9ji65
8oy630njL5rwr5lULKcG36fh0JvYIj9739eGaMM92364RA2/KRTYQOq954jB/SJT
fNoY+sj7+C9YHNsBwk7+kkeFseDfbVmsSYtRmNQQqTTFFOwDRZTRZTb6W8mp7KWl
/PCV3syoU7P0GTDoJuKBB3EjrrcCkXIwTTN88TFDT2tMVZfWOlDVtn1i//r8nYrv
D2KR88LQkJEzerUyCPlBpYVzpTs6O+5dV557OgCkpLZ7eDhbghPwlnyiTZ7ApMAc
oZFKxv3/qSDYNS66CLHLMFG33odVuTCIGhM591TVsJbv/x9naJYHD9suBzDA/IXs
ylgmG282a19th0MYSFD+yy73crHRGDnmLQBPY3Fm9UAQMU4DiMu6s1I+XoRketqh
WAFNHyHDEBfXZMr0PPe1WcfsU/RfSOHDXiq6ZkadL7qwtAqQvmoFYB3YINMaNDRu
F0CkonNada+jgIWVVQZsDmyHfX2uYvm+eAv6KcVg1Fh8Sin+dnVkm8RypoRPBUVJ
/tPUXOMBWaDs/ljWh3UDIvWxBWAX01wkx3qwCFlMjQVGS7Ol0Mb4tJRBRZ1GgZo4
WAJcNWcl5WKEw/9DSnJPfog6WqqhbUpkWSGP2PaOKg9FOka4Gm2QWTodWbQksDXA
n90DiDiZChg3mY5kiE5kdwVLs7GWwNEx2q5iLtEfldrR0ZfNlJ3e1AsbmOUkj/GF
FTZ4mfSsjhQJSJNQTAQrpwvcGcD6PSIQhqUP5jFOEej/G8HNK8TO+wEYBEB/n5Mm
EH/njWs434sD33I0Xz9BgRwZIS3/WAW1Xpveo0DNUodUW5j8t/uWygPH31fs0ji3
pzTFyI1QAu71vWvtXxcJUxNzSv5vze/pMgg3Agw7bUZ2Ypw7LbEM+vDlLXrL1FlB
mdZV5/4mv58TjSXkS6elRvtW8B8w2FFYUnDHYpZB8J/tH28ieIDIVV+nadp4atN8
QGampUK31lyUsT9cLscbJk+QpFQ69f7o+nWDnPcoZhzaNdPqgB1qb4GCztn211g7
F0h55hlsDPmJahpmvyvzYhvS1jx9O2ARgkuzDvdzof9vzms6gdxvmlNjKoubGqya
oeyrukZ2OvdcSSvTtKifl12Xjv+cN22eCBBG0ni8ciVEQgZTIsur8/ftLUlKNVXd
SjDQQoX2yS9W/kZiG4wsB02XV5L7N1+nSs1WRxqIQwdm97e8tEQYZbum/fKhbWPW
xYEnLu5lruasO4huIF6ZhbEN5Kw+qH7MJ8FgeHhkjgmmjiVGC6dK90enp/BNqpiZ
ybqbOCQTsYCGRSljIPhEjVLm0JZ0oxeoiN+9mBzVDDyxUJkTnXFZCxw0mU8RRriM
4Xvm31YrJQIwiuPaXlh2HvGg3SFmAZP9cE8uB7OP3bFcKf7gcBKck3MnyBuNeRJF
zOPilg9LjQwqNbgJPwUmMx+M/4fcpuspdMXHUnjumHonnvNGAKllGCOnaOSzCKPN
JO+5r69I4m+h9e9RbRNOIzFowPckaF5AhhirGV5+92jeUNAyrmDq7XOquO6lve9+
M5IbfqJeCt69ApMDpPLc6KAtszzLEo0Bs1MHrOMoBQdmbHAgR2N+l67KgjlbjNyo
OFLsHSuz35/n5yD8jH+9bRa0Tpi3DZJqzFyZcbyLM2BGqJvtvcHYhaFdQiokyn/X
kzrUMG+LReYw5bXhteaBFDWOqhlGjMuSL6WOlf0SdZTc/cfIzzkX6/wwM9KZ8AQK
FrsI+Vqfnpbk2LwcBaXeFIYpgWgE0wuvgsWMECb+adYr05b196BeU8WJRyPGmZHs
Csl5YDu5DYNcerhaw8e8gvIycXREuEI5m/LyrPVWlv6dJWhEFnUd3vP+R0+VX/Um
lzzy6XyB0n+Z2AWY1CtBDi9IHOKLksSHW3qgmLhPSt3r+sctlfnOOAtDmmm6G2h4
ww1j3mD7U+J+pO1w/gj7223TXYxPxAhRYpBTr0FY2jNx5IzXC9w3BKOwLKn9nPkN
hkzYQTZLh8GWkjQArYNOxX9H27dkwLxrKcWWCKaOU8tJV3I/s1f4St0/OzyF7Cxu
f88+EGY1A+wPeTuJAf+roBd+cAG8HnXUiXYpZSrnWljhZiH/EDn8YYNCz6AWiTCZ
kmNqGkffmLB77PyYDofGhWtcvjo5MA7qIOEcvKpIAwaqgp14tfD/nhehztPIXgvi
OKVfEkHI6NJMft3Uwgzfd9r51ZEPaWlL4lU88cj14tBfexLrWK6sxcLM9bAibw2o
IsQ6SlwzA0tcPkO0RYTs3iRAiOnDC0rRSB8qYiIPcHsAwWHxOOpP/u+g3+LZivCc
EhneO51XTLlCEEGXjjgwUjenG4m0aT3Y7Ujh+LQlIPmm8RAIbHvO+TMi6d5pJanU
HhcoujJFS7u6IWFwh8ujyWXteJvgAwHvrxRxd/OsM/E4qRoWI7uDIm0FniBAL4F4
1bFDokmnzt6h+NDPBTo9X+Q5KricBgOGQxIxrDbNKQwqOumQ5wz7FHsXv9uegI5m
KWUx2In5zuRJQLiEu984GoXaQdpXHviWExIdgwho8wPDQd97v6tVhDxzr0dQySos
d7WcvFJRSMGmburFSNso15IjRBXkuki0TQnfaULg11eyv+Ksrv7+h+tgYHoMdfoc
xx0UZzONviH7V0BHngBQsuYh/ViiGj/Ff4IStpxRNrmU6K9H4d4kTsBcuRR2lTjE
JdzPe8v51ymjBC9wcei/8DlDU0DDDajsLrpXz0TDHAyv06MZKitjZdPxCRHI3lSx
vsHCf9kMSRWcWPl3YMGrM2ibzFLC6cTIl2eYU3hvZ+agLbqbh07ZCR+i1YDZlUHu
XTRG2/cKkiF2fztV8Rcbot7DBErSwdaOPp/stmED9tbuFRVy0n1VdhI3rI0lKruT
tkFGXREEzVKV+IiknUfHtF733xqsfaSd5od3SeM0VWHzOBg5hCyexH3j3cn7lbyy
SpWLKmelq8KqIkERSus7aF4NOboF6j4Tt17as3MD3zdsds2jke4TKVR3iiqNGYwI
64IfgUFs2mBPfXh2mVmO0YdUO9UVYPPF3CUXjWxKP5aajDXadPYjrpeXfT2GGcOb
p3nVFZtcR8yVPTqW5BmEOXi+W3H41tG3TQA3TockrWTCgzxsIT/B8TlysZgr35IL
ZjOyT0jOl66wbAdNJrpFZuM7SwqR/AdgTJ+FFDJ2FfZVB5AA/lIRVut5V5YXIZUU
w7j2TQ2bquON9/yj0h9sGiohFxSdbc/+V7V0vzp99JIOm+RiTD+G8SHPp/nq4W9a
RUWrR+bYFr1PKxS4xozOvcA/7JpnuPxP95peOlAmJ+cFSfqZdnkgdlfMz92o/y1m
jFoI4Xg10WBhE3Y1k0D94KGyo1DrzLIx+79s9zYMCk1kjpqXuV0M8CCd+9dDsOoH
LruBy/+gw4uj0W+Q9IMqAHoY8tpZgwKyWUVyx0Y1G0+661fCleOqKLCZ1fHEQ/30
sPPqZ9pBEFkufDSzqLxeyOnQeFgUJc+lemAz1AH5jGnl3v5Yk6N8AqF8uRXGfmaJ
trsh9vTsaTZAWSdW3JOet3gT7siHiq23gAJPIx6+hWvJ4vw0j8aPs+iXJcJoZ1R6
voEMKA34ASUIt+8TJLNBGpG94mAIEfbpjqtW+rC5rFBLcYTIxKHCUI7rE41TFX1Q
fPuppUVRDztgQQapXr76UMcxts7rOZPpT3N8T8V6lWLfVsVl44OjUpYaUT6o3jDO
hBwQDTrrrhsUqEwxzuSAU665VKj/JRQaxNFa3u2bFI+rWM7cD1dFbMnQ3D+nqHGb
9MjWcz4nCq5vubtq6Uvs4iZDZg2hx3B7nXFhZ69oCSHUHf+JdlTIdwUzSCX3gufN
S57eKnfPjyBW832ehYo2qPUSvQB0etvoKvFV8ueqPFffjRjbRaKhCzTHCzFP6fE5
Qn9J85TTqhoU9zNmWxi0ZKLy/9+r5ooiAFChUo8kqjTyyZx5J0I9qIg7llSVxC8/
tRqftTjKwyIbDDbyGDPLHjQWfLfoyqHW55toBdmmw8IA26fk7ez1gzjxKJdh+bUX
3iuzYl3vkxzELZW9Lszc03aVdCOEuS8cv7A7SaDXt8cGdxGWlPFDKpk+vt1w2MWS
uNgbeGc+yIAzBWfSkuCzcVpZGPlZLrftvfruhfyh+RNQXX6oxB1GuEgWZf/WJEL2
7PmmYYCH0KPVEXyKcOTDluSVl28bUYfTIGl3GXOVf/OiQzG61U54E8oDgatuLA1K
ffrPpn3u4kN36VnYrA9J+CwlM94z4rnUqyKgyYToIHT99FBi8LcmcB4pn4dzDiD8
RcuwdnzcSQKX8+JRhTjv0z+zpf0DHnhrkK9ypZOO6l2KGSdUy752x8vSXI27OWf2
fzb+o00sOzRA5GrTygC2MbDtFWFtD6S6iQnRIZlBu9MB/06cwKYs0MCJFCCc/Rpm
rBnj3ppWm6KjNE28KB/mDGzDxSX7ht3XuCDFCUez7tKoIuZ+9HDtuL0JLL4zhUO8
8R1W1kWIDEvQichEks1M6dNFJxKxvihb8nKFEDE4F4Wx7D6HuBsX9W78peJnavih
COwYZkzuWK4h/eTwe03Wpvp6iRiLSrG4LS5nnTachXlkN7t+laprUMq1o301DKvE
0hqQWmPJYPrIBAIIL/BIVIAdc/fviiDx3IzUSTFa54SamLnsToosj9RKCbnPApqR
rbaaQXhxPhrLDrSeyzUW3Femu276Y7CYqXADl8VgVUwehzuZPtuBprXySUhvGroy
t0JVL92K3u7hT7q2oJrBwuL3QGWH4qeV1KhVrsn9hn0QquNwgYOxYulN73FtZhs4
evrQbfMzz+eh/1BdGutbQC9bOLS33jLKMstMBKg+z+TKJUIN9BQgUjK6RW0XmshV
VStVNvs5NuNPySILB6CnzlwIC6+nmoo+trnLVCfXbSWnWF8bg8NIVpm0zYBsnhCI
8nZgIn6bSE96u38/xYyGJr04qzS4+X2/KUGDad37D1pdL7aC00J26q2eXTRu7K4/
Ub7rAUier5xT9yiOQvVzTVoPkGWgOZoKmwtdP7Tm2C4PIpXeRpzvFfasCmPaTFBZ
6Ayq0E3shHOHJGdmGGyyyjQBnCPHUEVCZ7vnFn2E9ouPpgLYrm8y7s1fU7twqse1
Gm35dWMYNF/RtQUKrN6Wd1aOMZz+vnWlkrHTvPI3QNWsScWL5IsLIGROcMgCPCpa
mQNplj8JeQ2EzZssIYtyYTNkSck9HAQddafU9Az6VnCs1bXVWN4PrKcH0n3KTvvP
rerxRt62yXTkhOXjkDHvAbOhO/u0gS/F3i7GlfFL12acBuXSAKL3dOw38NX3eIzY
0+y69zr+lmb4n/YRvaMZTvySOcaVK2+VBi3OdnRp/vSYuJEAl7qbL/kNG8f2vSUS
e+jeT6NJkamDQrvCT/lpNjcQRFnwqyawWVZ22Uw4EXLQoiDXIGeuzylDk/Ay5NQ7
GVi3ieqxilME8hgRbu8NI/AtZr4IPjiBDAPXW8qTUDXwSm3vgZLKzZy4V83FQLcj
vF0+F74nVr3+mD44Fvfxuxg1jnwKpF4GXMLdHRDRPMLh0Q1XzSEMYh70fRefGx1N
+QTsiOeDQBJhnJPAnxt7GIweETyLaZMjVp794A4wdZeISC1CKtkYKoDjUYyURSKO
GDOcof1D6XbmwlMfvwPtvNl8Y5PR1dKrXdDAqPTxznM4+/8Eq4l5n6OCbUZgTCY1
Lh2CdD2KO1WRc67fOQq8R8eCy2p712GjosKWfWHuS40RldTvERucTJrceiMKuxEw
lhLf1zkywHAAMulayhy41WCqeuS2zK0ucuNn6cJDJUWN0Rz+k3H2g6321y2XBIxm
FAl1U8Pi8oYKC2x1uefRuwRnbsO9gNtcukMM5lpdxRUDQ/EI1XJt5IIRCTNi5cvz
29+2+h3WqDc7p+/CsvIFAqCJ0gC0ehpM/uAS3bSRUqJWQYRW6WgMgwP6pSajfKj5
NZZyvdgVUq8KDzIpo/7dMJhonxm2rpo7Ed29A+bGxFsbcUGPMv1chRiv88jk8uRk
RZQ8V6MzdxgUR0HZv9+Ws8G6YiIBe0mgDQU64B7NpVHrF5FasnMId6r7ZH9h54Qa
hTTF55FToT96f7DrgwLj1mUIV3l/HuRZI1Z10BX+DKU++r2mycTfw9K7z+idpU6h
I/+ILhs/ZXbY51mZgM0/dNpfxwzuwaWn86fouZ3uE4g7yK1+WIZ7L7y8TNlgVPCs
mScHKEBKxwmEybtC4YfrEWwFKwIbS7b5tMb2GZSGq2u1d36Avws8KArxzqtA8Qgq
oAUs6hnmri8MaQJF4MPBa002/5BBtT2jbXm76uKPRyYotIJTG66DiiobHkSJAtY0
iAR3sGQKqiDm9uA048zKrV6BIgwT0/ItozduqlKvC/qANGqIYjhK3mPrBIGgQmEH
QjFiYxZgB78wTleyHlD3xmPzzKHos8eReh4aCj2+tm+ZYNJNGlyX+6zH9Q2iGaHK
rg0yAUaW81bAMUJO0njpUNgrKXLUose7fCjQ85NW47MUjQB02nsx3lbmHPddh4r5
SwZsuZVCez1FzZFvlRHUyBJ1j+r1WzyGi7ZLniP6HJnB0fekrBS5QBMtCJViNM+0
O8FLouL+oUuPozw77cW+kzq4/6/YFWDE0DwUaWPESmZ85paVItrv5qNs/MyGgEqF
H586xpQddtR/2tZ3uk0317J4FWvNYSYrQ/DS+rxUOLf0t/gcfL8rME4ptqqQiz8b
llUlMwmG8J/uMWLoCApd0AwI7Cvp1PqhxPDo4xMnggsK287P+QX2FQ+XMmEcbqrh
mX3QHexVuNdxH6671UNPkY3Zn3MWIg45ICWsV2GV9b0rTqz5J4RmiVNNR1XhrmkV
RckJOn6nLOzpCaqV/bQMA1asqUz/psZ6yUAay6bNRNjoQJfJMUYqcVty5PE49Njx
UqJiLYBktdvbX3F4K9YStp75ehmuKB2F5ItTCmz23RdtnaX5pRMtZ5ETLUhJI2Ko
pSVNasZedreY3bWtpJ7DiuyUfyciDKrvnUAIMwiTIE2xQ9KErXXcQ12dtcY8fKWN
fXv84HFR1IWacLs2018d0S9nRwHHOVineGHriQhAa5VcFyAhfXYrvB+/+cJIfzQG
1Hjnmb//MUMEPoRxdSeuV3xhFrmXffi3sYqYs1wlXlcAmzOmVhFyzsHBig+PDF1b
y5RjkCGEB7G8PwK9WD+mdPpsJg7Vd3p9D4Zf9AAAw/AFYc4cWNH3zW2SBnutrIYw
fjx3HDMwqMrRQ9xI7/jGkmnIuRhEnzksbvODPRA9Y5CoMLZX0YFrO5dLa4KhEFVn
MKTQfIy1KAZdFwivjbaCeeEv0VThuYUGLebMCjKf+MbeYgJ7u/6MbOpIveB8jh7p
k3g5OiBHcFGhT6O3ZFWn5r+OZsPLGYlmsxM1A6UCatFmThvoxlMpzTLWr5bKDSWH
eZUa7cppBbF2sokblrhVnsq/t6RCZxWsZpNI7oe/xL3ooi20Gt4/E60fnCACTtvM
NbJS9bG34vHGGyd43UGXWDeixKF0EinMQB/qiQEbdWBYKV0Dk5EyK5LiUBVo+EMm
e6oBejKSlyWUPSykl1vVYtCJ6aZ+G93oeRnL/mo011wvvHY8B5n9Sy41R9qW0HVs
7Jj3ROoDQtvmfAbrLf6I2Il86O2b+vMSU5AOOfvI6AOSOautLjGrmUTlO1DTfgz4
9CHag3vkEnYoTUxYeYPVYewz/O3qpxF2NApAUzuBCEk+opADxC2smzLyeDnR/mjW
o8wNHl/ULlSmyEv4kVGudnJ6mzoH4tV62XkEx56rEXuIAmHQgZyYq+uzgSBasrmg
5dQ5hGfb66mhIfVwn2AU9EKIe0Dmq/5AVA1Eq3qIoORWOeX/3u8LPcLRc8U8/H6c
BxjDCKdjJlw3gsDiDu1sgGOYq+X5NPNTu/UB86qqH51lG9bCwgmYNY+08tp2sZIp
ZyylLTjox+xwr9OyV/+wqj0PY+WA1hTqIJelKmlMeEt5u0KKB50DtELRiruWKUkl
52gcQ0rAZvS1dJ2kxI3he/Ykv1uk+vswYiyDlR1khI+6D42Fvk45ubSGtlXqjWLw
UXBY/+M8/FNB79xteyfJ3s8/4Pmmyf78g3o6v0Ed8cWKL3dNeTgqugpra6Fu3oNR
GoU0elIigTEfpTy6SAICJuG3eIy0s3+sRQjPJ8nRmmCMCVoZsktQ6gDF38GhwQP3
Y+qaFkh0j1Goa/EZB0udOO6Flym8gKnsGpIuj5zQqaN3q+8KLNNK4OqGmaoI7esl
8xO4Svr9w/aIRI/2quLdNYaOKLShVAOc+4ux7GF1gx9kfnKjMV3vfbzHYUs+GNQC
yaDTlqkzaVGaQWklBo3bOHH9zuJI2Rkiwue/4PMjVPyt/HthaPTdH7LJ1lwfmDYL
7gzCK3iO7hpmcXC6MUg5avMBomNNf++qGS0Rw+r/s3o/a3OkJuNBg9sutKkFh3Or
tSABEYqaSts79VpmObs3v1GgzwrKK8mqt7tBeZ2kqum3+CQeFNNZCaWAxN2MOnlC
oY3FgCEaJJkzuQWrNNQH5ao1dfaKX/amnLwjYX7AZfGph7wTKQN0VZOKcjoIUtQE
xvJEs2axJaj9NMgcDlScyPtPLpRortAKtXuza4YZfMp0BqrPF6DuzvOpeNrRqsfe
ydGzpXHtLhR6qFU8AhvyCwAjSwmlB9OXU5tOLZgw5trssiP+crvDGbIl06oerMbY
mFDibKt55B/g/+zEezMg7GmAgoO8+UiLWoR5Qz8e64rw+UPm+7Whq7GVaGjLwHYW
aP1qRl9gSoU0EmXP9qIVEFIN48m1nxUkD8WIlof9YtyS4JqfHUdvpiR69ve6inqS
uWQMeJMMieTQ0AR6Fdxw2chmmZW+iWJsxbLuoyvV8/ihWMabYdMxyqWIfOxqCfb4
z0BT1K1yiZ6rKLc2amemBFQ1g0yyDPTyKfuuEWwsQX4YipKjNtoUlfcZhOdEmrsB
ALcB74VoEdgdWzwQRyLf89XPMrwbKQ+tL6tewd0w6nvVxXfndp8gabOnr79hil9S
Xs6Yc+LFiD3EtUxqfKElpEOHSmWuw8nz0VOIk1bB7e+xpCLDfic3jMO8epkHGGj2
/7BZ/tIJar6nYsL3jP/bleke0Mh/SLcRuDOa6tUBuW3Lgh/NGUBCWBhnfPSiTyAi
hRDJ4xU6gGMblrQua9Z+tMEFZQzzij7RFuZp4uygvSPm6JUS5Aeq2dK+pQ1+9wZa
tcgQ7YJZH0wm2nkfJVZQ8W8nzm4QLBMpIjub87AZXtnUcLx6Ttx9YXLbGQH0ezOP
GzMLComz5urUBzIlAOzkpDoaP66JUCrnBrpPrlh6cc3ReQ7NKnOXDpIlbhEx52NG
OqP6aBjTDu8yG02+4EMuDeLctQtq9jovVd3rQag4s9x71HgUOcBbcILFfIt4HU1t
/UZngxCrwqsIGoO1YGtUxZSevFPAPB9TEcjpumRU65WawvK7P9tEQIqkJhJM/B+E
zd0ggkDZRB56/E6v5SBnk1/IM9/Za7TMAREGvowPFAilDWskexjlWIFMhhLkNdCq
rTcx0BymAHO2xhP5QHl88gMEvFweWaJbS6Xwf7aL+Kfz6bmHKkeEm8RbdEECIuTu
YwKc/xNhHBUBSPtflBuofwR6cQuX3wL+q13y4KCnoT8oIYdx1kcpwh9USR03Rm6z
W+Dne5utmrkse9mJYbg+eELsUFat8bL6UR8qPk783RkQTRSaKrPa1VHI1fDgZuCH
w3jz3xx6XP/qalq/u11/LiEikqeFmxcKnRZfKR79f86jlWJGKnCyWRZpuBwEuSO6
323bJq4cDcXuKr+hq9/zMpvmmZL0u2QPCsLwtaM6Te77E8HhEFAf9AUSmh4W4pOn
Uw3orXrKIhwm6a2bOlP6toRPgbuAObjySUbicgWRsPTTeYpRsydQAun/ozD4czoU
+z1bBH+XRnvMDxJlZNHYcpYAcL4lmcGYfxAfnncrH4AR5IyVSeqhUI5P10IH0DsF
h5hF2Mc8nfUEdFJuw6JodV/LxgC9LgU2XdcBAEflzgzBcfRKwMM9SQ0H/uHPM0Op
1ZQODB9+qcXcL3tK83w712K7Kr1L8DeWYcYSCmjqLQShp635+NJW/OC6UTyRUdKL
rnrcSI7kg7bHvXHwXrunGqUIltHncC6xMt0mA3ayZ/Vmhniqih4KCBHImRZw+vqv
Tk3bzRbidGKLmQwbJtyYuaZHxXT0jJFw/PvMcZYAk722AnDlDXD3468Nd1d/hPtz
gTQn5n6tXn9OBOvjS2Rey2lPgefIl30QBq90yKhV9RUazhlV+2CDIjFgC68wIeQS
m/8/+YEd3urSZVL5HsWpWgcDw9bIwl0mxwsFwgTGF5t9spO040G7Od8EFdJaYlUm
D/7jHzJsT8WgF2kr4jw7Z1GlGi5fXQh6oH89b/NIWhQofMZLzKyB4ihVYeiSFc5Z
j63NAre+lv0vPM99tPjxFzLEXOSovuKdi4Z0f+e+bJIoUFqdxRK5667RTKNa4J9G
2CqB4R+fu5b7ETKQPgYExzqF2knOZhzAaxQiWUP1vjJ8+VocxEiUO7Z3hpFZKGIQ
z0IghhEJvEkn6YiXqvwaWXgixxn0OGIMSdOuwrR+qbbLOtP0upCQT6wUUZ+Y/3o/
py4fTC/4Y9OE3ylp96VDXS761Kxtu848a+Qik8pd/inx72q8SVXlA+H2cdzuNVdJ
iZ3BP2hXIdHpQOhsCSuiVqxZldbxX4rsvfpo/nUTJvJ39HixXHVUig0655zGSHn+
abNwyhTMG5u07QOMrQTjzV7SYV0wTr0bBSH7Hf/mN3uqXEPEINsnfrJecmHkAD7U
TkUtnikmDBh4rgcMY4Os/WphJACpIowV1gYfHC1ODsYeDRUAzPBKWXkq0cWOB+TB
ASaUBpQ2wy7qQQ4aSBVkHnrbhNHHQ/OsxAs3axQhDYRVqbNmTTlzA4xQhfdW4Xwp
2Cftig/29r9TIH+s1B0RNbJrijw+c3TlTbhNrVo1p37gMq1lq/DQf7Vkcll0U/1G
F//kmVDHEs5nC2J+S7E0CF0bYkocNXnrip5YmwwI0ifXdMnJ0KmEa086ts37nhnC
uuEnYCxolkJzWgIJmfiGgacmroipOieR5QWCX9aaIy6RrTmRyZ8QV5WMWQKxL2D5
MbKK60k3R1Jrift/mrxBiK1AjwWKtuCMh8qNajqkICg6aO1A7QOZIpAb5rr7CsnQ
XflUunvzfIM3LqhaXmpmVsGduArmkb0Qi3w1vXiIQF+8XBtUGJVz7aAETGU/x7J1
U/l1KPfA9BHfVcm6sEsCNu9rOF1nv01McJO4bY34fo0ItoVK4+hTNYASgc8kJwiZ
y4sBbKuXKb/GFAVcZoj2AautpVPkhd3ffWT+Va4y8dZvBsf3si6YBhMwU4KUaVhC
6VwfHr3bXcKVmKgTVvTOYAQvk1jxOs4gW5tomu5ffCSfqqAiaUPHCQ/TzKSmIF2b
d+bLx/2UGMx5nQbOv+Z/4hgSbJjAdpPWda33nx2AGREDzGEtvPOYduw/HRko/fsS
zF+pKbMP2sEtNEVNa90UF6+d+vVXmH1RDiLIaVW1tb54kobPfuaJf7eSlwgz6jmz
EwCzxL7C2SrXDlX9VRS7lS3qbJzt85iM5NlIk/d301pfpmjGQBYObWk3DdWLy9qH
CLVTVGpxIBUePkvOcx/qh6YBPAo3hfTTGtqlrRJqY6s0cNE+7yvXNeSR6eSO+kd+
LOgJvRDDktSVsXHyJC4Xr+z5n5d6PxOhDfN806wRxMXk1mNVeYJ8sdFGys/8EVUg
G03hp/FcXc/YipHZNf6Qsf9UxVYMHeQvS0y8Q0+n7ZGi0aQWsDkQhrClnqHCIhtm
QcwwWJaRM72Lcdh2G/hQPC2Y2sqFN2s4+Rvkij11/68b++0PY4jLuZh4a0rlrzoG
gpzIU1WzBexf1P+onTLIsYWw2MAsOup9DSv+YXNSU3SOxhPvynuz4LLEhcSQOZds
wHwWiaw2TLM8R5pixXxW+z3j07iS6zwsrvPza7ZFg9RBi3xtscbMYOm4nMLDrBGq
xBiVZhyzoJgPWmncqbPok/a7zhPytqjagF7YPF92KjI1/bGKxnkyXKbO3dux8x38
N5fAOi+t29xqq7rM/Cy023CGtAPsBpw30xbj3K2S7WhnMBPSAKda/LW7D8ZdnFaL
fEg/seSL2yC8H1eZmcgScILcK7PQp28l3X/Ab9Z5yLFlK2N/lmlzgj5lRgukP6SL
m6Zr5ZNv/TssBq7iWyNuzYnUulaNeFYXcYMIRgDcXj6OE8y+s/Lni11c3FLlxGKY
EC3NI7lmbtpoucLGk2JCDPAHCu/S662ONy+qKUEpUNCOw1kUB4gr3rjDF0OmTMHA
z6PadXWB0rhRD0SrmetKbpJcODZrExppQHWaI8U6OrN34V+ol/Yv8zT/GVehSZ0J
oXYxEluc9rST/yOaUd3olxLjrwJWf5q5zoV3QxLSlJ9weFBGNih9Ca2X3Exk18sp
VU08DgeW28a3TNJxriBtK+qpfhebXZ40HVch5hait+hTNu/CGJm7NxkA74qg6SAs
0F2nG/XcBjlRRfwWBH4q/iCR5DAtb+FXsSsblOxcjrbxT4e/HihvsTPauWg7GYnr
/gDLYJZRHqrrOfe2GTfxNaonQ8L69EVxcFEC3uMEcVEBzM7vLTPCow7GvSftrnrO
bixNQLsFFfisYN7r0kXFAzUn7GaFOpcXvmWmX7zqBC/Fhtg0Sb85YtpE0lbunq6e
Uz0w1z5ZvVUPzqJhE9GlxPDzcfZxjlbX2y7VNue+xNPXPfQO6kLVH439+sAtphXW
yF/+jg0yOjJdMw9WIKD4X04CozToPTY2KGv6zt2ii+jeaw2+mdDgvYMxQDqj/d09
+EZuCpOPbNdFDnvuyog992OQISGlG8QqcDF+iR9XTgebYbTLpbL5DniCzUb1mMFL
l+4kVQt2wmhLg/8HjUaaZNWE+ADukj2tA3FXX8qQfJevS9h4wmPBHeP/36UE/qd4
A+eLNuBZeaRAS2JWT5ymJT22twRMsh8Lw915/lpyNmddm79eID+2Gdgrny/3BfDC
TaY3ATIiJJ4zGcIuQwb+9JV0cKvLSmBHKvhU4fii8NtSdkrTDiVH31w48YI0Y34O
Pv2lr4e+RWlu6rXO0zy3B5zlmjEgHPCjEtWF+cOI6ygu1MhYej9CXYhpltimi6NG
rWAMcSafdrVCqsyWfeXsQMRmAuvYpkxjRCy4m8wdyyXwuCNi2QXBGaDZrC2gGFQD
ptoLrZ/lYrA4L9R80Q5G2f4AH74W0v1nCuh8s4mtYcZ8/MQ8r01MJz+yyukreYSB
BN5KkVOqvuGsxjNeF+H2IEY9g+NByPomhIBsBhVtUh2pTUsmkfAT3wOpAEfA6PP0
E3B84vbeGDPLy6Njle8UP9yTKR5LvU78gCffrw6dISPul8e+MllTU+pcuW+TZM40
zVlzPOkAWzpRkhcXAGRQ+217wuDy/OsHKWHaseVYpcs5bfWnXR5zPSjg8LEAwlQd
qXN4nE0shO9Mwy5ZjvnH1Aq2Play07/k0Vkp7QN+Z4x6r8hV7vkE3hwm6K/wkH9j
bUs7QpzUKz1n6aOsImU/xiEGyRitvZ1Pb2BLSxZyRfrj75NjfppYhymSrqT1rSm8
OQJH+UIhv/HnRZBiMgihuy1EbiioOWfEfhCoVCadbd7jEqMoiqR6fIT+o9GCJ3pa
n1TMUu0e3BQ4Gm/PiAW6rOlmnn1AawvYjKPjoKae0hEdnarI+UdsU08DSM2K/K0h
itM9aO80VeC0dofBax/1zznRAzbLA1iSDREXh1z5xuQiUjNkPO8XvRdO6E7OWQ4H
OSLjoUlrhv1XLXYvkVUt0FMhPxEcuutJYBPiYwlBhf6PaPwAebv4btq/oKJz3itj
w7l4XKjV0fdv9GUYC+cqdcOvp+jV6LhMbGmXPQ9KlG3KupuEy3WvvuYJpNv3McVn
e8DMpZum2t0d+zTEPdLofPK0KKOAeJvOzpz2CG5hXfx5m9vOsAc/daoA+qd5Y8QH
HVTYu+RSsVbgd64OQqelZ8ieZXqqZ3A0kg84sf1ulXw19EkYq1DeTJoV4DkVAHbX
wD5oa3zgl8PFywlMNE8bV252sA1dOniQQtooBkQa0yF3BubBq6/KAiv6fVosE828
gsl2eeFfl542duxMSwCGmlcAETPj9zmnpvjG4TkcXZxLT02ExkuNJc5g83swp6p6
PxpuWNh0U+UVglf4EpYNRNh1njT5WgL9I52ptWDKxDaXzih1hsypVse0Fj1n2aOl
BYPR/REwa3wvC2m6xm+4ecUYJEkKnb/cushngQ1x68kzpr1hqO4/2JBrYzLGAlDr
2nr7JrqSaXj2yrc53yUFLELDiqEBHZ5tefL1bHIlQCjDvbOLXc53+G5X+DIRWvGi
hkXDbLsmplq48EUbtMQmE8DQ9fwGbDfY7R3FBKvPA9Y84evBWImzSgdvo/x7jfxW
nzFYWK2tkr5gcGwtHGJn9pPUjDzJshPjqH5wbN3qn7evYa08KvncLSY60oPd3XAj
IXTnM2+X+d2cB1Xuvz2K2ZOnF/8IJcV57E3nWNnr4YHdcE6OnpmmWqRCtw/f3CGp
/s6Udi5+IMsEOFfEReTG3XG2YTRRp8x/RX9iKfDsQSHNEg35kWbSnYAXIsS4YBLM
T7fzRVU/UnzBrba3f5ReiZArIVp3hsRb2hKsQg6Dh2GsSBLdwn1g9mbGVs8IkDxd
zButG7XolDaeMnZzFXd1mzr/iuKdB4wmL5T05nTgXHvrm+foOBPDPylV35fQiXts
3I9J8te8npbjT/BWiAwu0b+XDabGtKad1TxB+CCz4QIPOGwpv+fCk9PAvVmM7uxy
aV1kYwwhWujYDYgEUb+8Mbtc/cxhuoC8ZGaUNiT8yzPw6XTn+EK4TRZqgRTOO+W6
zH8vuOwaER/wv9NeO1qoZb/5jL9sch6V4qYUDlLNx3j1gg8N3LrNy/r7rcq1mVql
PP+oohJ5BI45G5DlcPCUuKSXHubJbUONAW9EWq0cvNQOdWsY4R635ASGsXSUVbX2
Q8ATu879LXjofYgL5N473OpcgHHRUibjGu+e6NeNykqnk5cN3dBW77PzgcGOvH8h
LzYviazECrsyTDAmvP0N09N8k2c4Y/D8NrDnozo2cPkzeTeM/y2UoOs0rJs9Ozdx
D+Ap77B1q53QnRtqh0a482R+y8LhEqy+oC+xVu/YhLG1OgBEFN3+3vxihUGfb93B
Xfjz+uelQK9L8/IIsR37DIxZ/kGr+cSszKQPZ3AMZc02bMkY4wIlX06q11gPHv9M
DpsvwbFAFZrRIANqHPaRTQ==
`pragma protect end_protected
