// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JXtOHM4IyCsUpM0T1HtQyh0kSdT+A8dDZr/GpvRUK1C45rqHAloYzGCUSpPu1pca
bc95Sij5F7t5Fi85/ulJMbLVOqifgCHDcVSn3XiC9n8ES7yVtICdE27tND7DI0OE
4jOJrHB0aSF06eqAyw7Pn/YxfRyhZWvBPHSVZ3RzI7I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22816)
cPvfznoLv32kLnlosrR3VitPcC8XJBle+mDVIbHACMd6wLg79sDaeHvX8w2ZThVA
1x8COEm/4scuj5+HiPCrDqhMBXiGE2ysgMXI3T4kJS/+1oiezWzSX7FpRJWndw7f
BcddwEPnkCgu9JxVjChJKVPBHF2cDv+9A8BCKnhzs06TK9MgfA4NPsem9OD5SxYE
YV6XO0o7ZsCQgvZTWFiQwfINL6IvOe1SGezZ9/57EgIl9OfwnFnc//2bm2xHNxDV
Gx+exWTOW29j+d75DoWgr2jKg3laH38D2Tg3kc+Vt3SyFn6CDMKUqGekYEkpAgB/
KwTCyGHxNmnTx1ydDQpt8xGDxfWBR62K1Q/cGNH4tOczhhwIB+U1K+QRmk+mzRx3
JJspoH13wAwWAwKke+8w0wsXNaxAn78Pm2M+UzFy2rd8lkY0J23UdeAP62k6GW0k
K105Xi8eYS6QW8su8gV91t4NVMCbipr2ivFLKdCjmum5DvTQhRLLxpHTmudONIk1
2wx3h1V9hJokTrlAdNC1n5loc4/mv8GJh/gjXptXde7cXYjzPSEz8wt+J5DNZA5O
HM13e58DSCqooH8IgY2WBuXNRh8kuzXy0fsvtB+HLaJsti/1V7RMyGqFOdKifyTs
VP6MuDepCKrCVNc/SesiINOTLO/UHBkZo+qcbEEGGbgs7liaGpz0nTRU4AMQMPQu
B2JpJ+AW0BMvDspND/+TLpkZoDZXGtOJ+0ahEe2g1MupyHRzssGvtNUYdWHcOj/x
ED7ouXyCdXq9GDXQXpsniHvMX0R/BmfSmzEwY9zGUNZBb05fLrOSnwIBmyPLISn2
fSDPR4Jxahck7gwPHOGIijRSGD8KOYqXBpuqEO1hBB/+kDVzH9VrFSZtJS5oikiB
CWNrVzBTISjfOlZctHdclLrk4SN0q58DZva4oy77eVLrak5ETONxxRzbdKtegjsw
3HBxKxp8lMzTxxcx0JifQ0yc2suubpTVs8BKaH7r7K3rMMF8MxYGc2kDv8wt2tWD
IVuIepQva5+20oSWLHiflYwHd3rpJIm/1+dDGqNCxEwwZDqAqXExCCiLfhZOr88Q
Bb/J98QtFUiBWMSG59tGe4xYNO07oooJJB4jNGGl7SHg4QABWqTlTx6Gl1Q7yALu
dQsAPM2EpK5v7BiVte+UkTtiVsHqyaizC/rvZxN3csXxY+2602gL4vA7tKgi5+BH
1rEfdRXnBNEsfWpoSIlO1z5LIYOmS1KNW7mMPchRZxxKGaQe3z5cwZoQ0BQsz3k2
5akWPMy4enZxLL2POGEyW93KXSBpNSkdbVefFeNRzkuPsLdtSQEiy3j8X2v090y8
/sIEgejUQYfADnwMYKULP6nU9GkLYZnTfxu+JesrTGLFfEWqYsxnDE4bRMJY9y+w
bp5Horv3EqDidWrhM8n7wEjRju942rztPfiAFoq+nBok+O5/XNK7nub4FjLY1kmk
U4i6tztz/CLjuMn3+Qyx9qEVYKMBVunEmv4f8UMl3kyqzaqWCjnpvk1cEffxoeBK
Pq4sdyojOgCFEwnV7EcKfvilWgYmZr0KJw6Y+8xA6+whdt69e+v033+dn814doWh
/0S+/JMxBSahs18ZZyX0upbJB6o9912UmiOeAu0WPuGpdFNpkGVvOBIQIgLyv6zo
GzSgs5ss0ThDD6qP3n0xdqxPT+pVTYT8RP+N6h0cefr4TVGbkflrDd03nO6OIrZ8
yV2ag/oG2n0lzXDaF9wCiNZDfz168/13mVnw8x0wroQ5EisMwhZwEtc0vGScDfy8
Eb/YHFd1V/ECNJvDK4lEXcqrYMwyL5WAgRCLMC8O8LgK9UAF89XPqJO4QvaEN86/
g2U1ou8KoKyvfhQ4kpnm423UYRNHERNAPPmWCpGwEOHDB/wXMB3b2h5/n0boSETw
M5kldRZFWpojGSWN4aUaVAYHDSlRg2SnKVdiLhiCs5SBKQgL3NKmDGF8YkdW28yy
pXQ+GwdxWqEqs4+f/v6KmZuGXgLo0Mq2rRaJvywbVbSS9X1mLPk92qzYGWEI81aZ
sVRaMC0rUz3ZEsfFvLsLRtA+OE2QojYSlYBjVHWrqCOczhvXe2GKqBj/BZ4xsmG/
uZsTX/qHGzCGIVSNG8caO7T36D1ADs3Y1mBVt2hvkQqxN1valKEKqkJ3YL/E5W0j
nwzrlrdPKc6xqZ7YPpDeoeabH75g3WL4GdRw2dKvnhrhFoX5/emyw1bKHvwXoQcU
8qUYuH4Njz0TFt0NF3/e1FEOgbbywd5vs8xgBKTW63NCY8Kn/P9vkFz8VoCN89Ov
fupq1/2dVQ+iWgLFdwPwCWjxcf0fEghtfwyg93cUGgpSDXPBopSLanJ/7nZ/MTUE
oFI85U4GfLAPCXAg9fT4WmrJhU1K05WJgzK1o+k6tad9yILWd0v5Hj/RthMgf8dh
mpeKLPO2reMof4MIJIXUMLxOjQR1PAdmvCJWos5sG4+CIVJw2isgMDOWqufB6z39
0n3h+sNMg12g4ggqO3yhdsK0WMaP4hSpC6tjkZfApieBAHfjyed07MDN9j7EJ89U
lrGIJ5edJQ0q/Of11e+rZ12ciLO98CCLMMzhuqpQp0RKEgY5MzXzdysKPb2Prbcf
5vAtRXopz7a3psMFT+qKcilUe3kMjYJ5+lhAOfSeuxPlR84nUgPzrWGw6P9qjuAO
nSXdceJFOF7teWg/8UyNOFYhYwJC+G/SZpQmXVZXYK8NUZGUNFylO5QJZhzCLRy9
zFBtE75XKTBqOoleBBLrPEFGBuIcH7WoXnyBFqrVv/fd4S0FvR0ss6Dk0xbkL890
OkEfVmwt3ULL8d6Tx1CYde3apy7+I+MJdfFEH78eMfasioEwQx6C7FS1REm8wYUs
yxzcdGcTCjInWRNPJ2rGYwmIGaUlYx9qQkgiIuNDH906+lOYcqxHIbs8Du01lueW
VFGcia6F1NTekaPY3uV1nGporRT+8jMLC0mcN4HcQlWnItXiVFeRB1Hjl/KovtBW
+rSHvB3okM5kTX9/40r+wOXaxVCJRBPFTsbTaMft8+ks463tsoTBgdjCKqK0zBy2
OeBO/zxRRcrTQpI7Bl4DdM7lKtGInITS/VHQC9AthwDN2inAsS7J2kNjI6QARjqr
cS2oHz2HVoF18QKkVnkvkoy/3EeNABF/yoremv0d/rdGrPmIoMIfFzK8tefq30fV
xwWDsYWFiARD/uD64GKurnR9iPAkcOmOzScPWh1UFhG0vGYRgszD/bpFMNHdljp6
x9QRRatZ2fFx4qs0Vwb3qJMZXaLKjvWj9qL0Jp91UyBxBJwgwb2cbE9hFl5a86QA
evIZhRGLg86RKJwcHn5xe1OaOAl5Zq+JxpBbfkxt8ZxkgHGJYmS7c9pnmUD7mnnV
dPrN1GgZQ85p7x8gBVblVjXglPbVhtNX8BvIQ69dtdGcMgVcCnngQDehurwtIMJn
txrNHBG20W7+QG8HshkYMc9Ka/zpqxC3+cTDY/bdk2asdiaDqjD/4dEm4vkOMnRM
3cDyctjE+vXSzMLnmvmB+ANLYK5aFHz1OWZJoOb6jOspyT0SqWmiXjJcJVVXxCC+
6FEfSwK4MpSZU9dEXo9J7PfmxmetL0/CF3AiKIZujwFFhL8ExWahm/HRN9KN8aJZ
P7H1OaCjM3m7/HZrILskQ1yNVgVMgZrOAJ7NXn1Reh//vUDyUnTdQdZzJNlWCFZV
pb7V00bO7tYzwPXmxrOlmZGDm3zKiLBc2U66mexm0V3bC7npTIgSvBVv1t+hJ99v
+kY9dooNEuI+Pbhz34u4uEAwfeiWjx0iHa6kB1jpebb6dPhDgq9eHtyXOyd0KJc5
04diEYKPSFILKikjD+B10rDEhIkXUOlR1QQxkddNq+jAnwTIOBjxBE71DkRjPa72
E4v9TJlsJG0jUJ/C2iHh3HxR6nP0tcr5PKG12V9uw4pjFYg4RR6s7TKGM4cmfojj
qsAXgL3fEWrgssrKUqbPVm6eDhPAwlDH2q5z85mW4JUvtYQLaPbO49snAMTQopUc
L/sFs5CIDK77vfn+ejHnwKEKz/kns8lDRLweCPyafYDF0jHDCapVXU/acbqa278W
Ufur3fmXqM9rSC6UWZp/YjWekJCPp4owZ34ZZ94kKdaStrJjP5NWrrG145Dbu2tA
o2Rgw5vEz3NbIiRyWcGGxMbPVyNOtqgZQbzIS3YjX8ebAfqW4RtPCjq8Wu/vOrAV
2RV4tm1K1CzqOmHvl+2eo4c06Hlr9HDTnVHrqbuRnMyOyezykkFaGjMeorFLOhWU
vqBb01RmlZ3LXYLlHba9aoFoxM1LJeqLltG4BeqKGU1rd/tCHIitSFhZqTzbR97j
XbTs7kBne0zq+4h2rZO+qMHgla6jYjE75WUJ87uOgLC4tt/6sQewSwXpOiTSVLZx
apB3ze0DXPY+kKtdc2jgK/vSEi7zl5pzGt6wFtv/AprM/8LKrJuqYSqcqpx6Bzop
ZhOfVLPX6BLh7jM8oNcb7NOBPx1mVxEWgm9aP2N5SiOiVtYn8Gk1yxsbPnsZIKDy
0HgzsHNTihzJIz+H8cTIK2saITLPxtbqCotzN4yt3c9m9ygC/iD9LR0POoTWACoO
TlSc/iPxRIk/+ZxT15sjoLdh16qOSHxkxlbsg/8o0mTtZNJchOne3a3GckRXTShl
G6uYTe/8zkYsxgtLjveQootOadUhaHTBDkXZmfDEkbkI1redc7m5kIzN7prRZ0uI
VexGAniQDdhjyEiJAzLCgCkOQU1+D1MY/L7vfJKvrcenD8u9asKsyBwszsJFnz2B
t775Tj3f+Tv1Kg4Jbl33lQucinUnmGrfxIaCforeDq3899mFwTLBqAut3MmUBmGb
/m5u5ikHgHm3dVogJhlHENpvH8FpHZSPnWhx4ilfaW1XxOMmA6bKdq8sar6Rs42f
/RnyMclE9cNQ1z0SGvj8SpovB6THTcAKpc3dXuE5FUgSpCJC5YqPQV4V7cplRfot
bMHO3Zuna8hVh+VeD6ryhQLytwgTM7q592sXlfMzJcSmpUs2wAE+Qf0G6EFJakJo
2yLe/minjY/NzF/YEP7bBnvZbjOrIDS+DfsmDiHXNPyomyf4g9jWJhjN0DqeF/4w
dQJH4FS/jxSbSx/Xqc7OfZRqioNdb7YHd5WAQFdjJit6tR8oR7j5D9/gQxprsx+e
6UwrPnQeApdPIPDsHJS/sXSiLtGt1MemiCQ7ypGZ6ZSwcubFkjl/s+ltsGZdtIim
QZZtuZIFM0J0A45VjybA9Bv6gMv3yYyZSP0VXOrvYutjA5U8K5cXZEpwvRktNpGT
h7cWJCYL6+pgyG2FAtabdCTv07yzVDcuWu7ykfLMX2IYxZTrwXKUte3s6NKqHY/q
LMm3NyEucC00kOdpQ23YOPfmtOrPchuR4RCQoPfISxEgVmcb2u8RN2plA6aQBC0O
fR1hg9HkTzYOozrbi9Dw1w6iL8iOEm0YoX+GtscaoAkUq6Tb4XRgfC8ZWZ5nOt0o
mgAAa3gr5qx4waHEZEAFAfPMaMD1Z/nKacmeUgmTgGsWvobRqsYxD+KgYD/dvpzL
tj2yOn8UD1TPLYTz8Tl6YzQ9ddM3xnNrOevzn93iU/66IRMFehpQJEjwdD2URW9O
q+lDMa8EiLJgoY2XTrimHNYN4kKUDdwy8Kld/G05WviEaqk0IuV/ZVThCoTbAKNf
p3LWPtUx5JaudNbx8AEj53jfBqs30zzGus1YHfHQ5sfSedHAVSTNM/6ylO4mfVFw
swGKxfPIprOPEL7F6GgEa1ybSJ8eqZWhzNgoSKfccW2tEjYWL/ZcM3RMpXjD+0cz
y7vV6ZExQDQybbCozIEl9SLK9OdzqZoRgwMCCDbB5n3Pf/UnlNxbCso5DkXxfPOa
XLGrlQkUtODGZZYb/lm0vU8k23MsYHpItte69hHAfjuLvR45+0HVg9n3E/dx3x8R
+gotlUz18SKSKT4UCRKHXIPdAwpGP+M28j94nVrPYaDmsWfEHONiCLNPyvJotGh6
OpJmJbx7vQgyowtNKoiEw+mzhW7J4XqrfR+xOPsc+y6ro1ZzrQdlPASbsf3FUe1E
5jMyiiw248V0ePBPeWzpFua47vtcp05TNS4O0MUI8qK/GTlZ3ebQtHWFcFqLMI4e
1Fjyi4bL30H++77TKARsjHEayJCobGGYjgFExPh9fIw1wnlP51U99iZqXMmCtgMi
vfZ3HucclG2uVaoVIqgfIlDpfWo66W6sErfu7387kYwlwUsOgZpN/HRJJSbh+SAq
yolxcHxtyR7mFP4XbZoWXIdTD6qrgaGHKzX4CgV6Wj7NeZgfJbqlyWNnpU69wOzH
4JG/RUkG64EJkFtZAIJPAh2vQAaZwEs+gRO4dlyUglFrz9SJ41ND3XGRD9nKLKGu
vkZ17zeNFz8oPuPRrKWcEdDvcAp06Nib56bt5MHAfoC9RvDQ6cvVtlpE/ZpXtHcg
8UE/ICnBGItHqwFd1beEHOkRoLBpK+aST5PZ2AzDIXr5uNXl0oXlmeaoxwvMHr55
TUE5Z5igeYHBM1Q8MIXsCD9mHtdakBnwwufGYj/0qi2DHrBNFdGVWDo68Dtselz1
wTJSEk7RFI+ob+OL9Gr9wL8ZB1BeStmKt9soy66qwDmYyve58PDHpYcAeoFfR/w3
Aroxgi8rQm7j9FkAdSnI9nfKXoN2yfM9f6q0bsF7V/bcAwZQ+ltZIl3M/Y53DUF6
WelX9JWfrbBG0z+QlYNsIABMkWTi5L8WRmV6moM7COgKFjeu7rqCT0ua+4V5PPsH
GZQ9ngY/4YexH6KYHaZ3dJYsrXo3DidwHQJvUXQFyfLBe5YIVmOrjfHpNkIby3cQ
hIUxbXQAF9QKNXsW87H3dAzuoIpdqRLWb08AL1gleAyeAoKf/VRoZuY9RxaM8kL4
G7hmGHlIFEs43I1WfTfpJeuLz3xecULpLV2ieK4IFFYzZJpVGbCEmDWSHyywr3ni
Vpz7YH+KCRLn6bjUwAVR9Dd0pQfTLYrEEuZi4/hYr+kzkZsx9biKKhubJwwxV5GY
rL3ycrWgXnkPgvf3bGBR1F+5YKnv30rAry0TuGLZgShRllISsNw1+04okLkfq9i6
zv7CrEZrAzB1vF5kdDqnrYBHJxSEKwN7zW2Etd1QrL2+SgGDXEFRA8LGlFj+BwFl
II9WbL/MCzMJ/63KBtDTgsmb3ydbgOGCiegaBhvKu9AubLvdjwTyXMwKPW4fYHuB
KDRlWFeEwXCOQLXFx30kWJqVmZc3rdxQ1gzk/Gp1/LPrp2dB6K/wKU9KAlih6Z3Q
SWAH+VatmiAHBSG+oHiTAPiU7WZzNXtLSumAHbUHc4shkUTZSWQpkGFoPXzkA1st
P86l+TaxsaTJ6ZyYwfBCMuE8n58nIGRX+XmXU9uP++ShfURxuuzHLqfzq2RdHrLC
pGv09NUvAFh5X8Vw8Eyof2ODqUPAzMilpXH8uRLA/bAjtUmQNJ+v4w8qt59lVqVG
gHEUn4UxFsqe4aW2d7GloN/uvSVYr6egooYafum97V7lsjKOJ1F2OK7XvyPhbhLR
FlJm8cMTL64YUfZdai5nBQHt7BIPlGrw9YBGQMDMDAGiENWf6RRf8c34an6QkEml
YPcqz67W5bKv4tlK7nyx/3nTDm5IJI48bhav/CrhFg/GgLd44K5yyev/2usZDSSZ
gjCVdojHuROhtZvAKLO4+1OI6eVw8hXhs1+ActI+1yLCwipLsNCm+eihBrXuxKyr
829BwTHkiDsYxmfMBRXUWuGBbrqD8BoV3Bndt/gsSz3JaC3PHBMhpVkVhzdArcOm
q68prdrPQZP3cLxkJhmJt7DHv3AKIbB530+hXvQpbR3ODriI00gL3Qr0T4sk9C3f
uvPbHOrJrXLM40gWCh1gpD8liLxOMIAUIFg+AQEiCqbtbFGHcOsfOwZi1XnvcbWe
nqcQzYgYUBlj1UWFbgTFMxcGtypE3/FHjHOuGHH0sp/Xhisvmj17sZWjcO/oI72g
tse27r/f8zcFiVVTcqPxMJrjFgutaLEwWFsA09I3XhHV2NO9zXWXeYXIq9swwYG2
gfiBMKjuJsS36i+RPOuTQxfljZQGAux8XPJPRy9mDXy32fEKVnhTws5iT445FByY
1wYLv9VMvddiiLjbZu1vY5QHh2YisdszPXgyyJEulrU0KmaSsMse4jRcWH3Bj6LM
NYAxhIhLIco1zXr7tKJWQ4PmXeU6bHjZx8eB131bH94hd+pYZDPN2Eh9DOKO0hia
NAeXjwApagn5xysf8wd0c8YJNQ+2XHcztPXICyCfYGQ5uHekf31vQkrfF79M9ziN
xolwltoXIR8E32pClP39uYLNsWzpbZDH1YFAh2guUCow2OLHwmRgKIoGS1qiFyXP
VTMDH5bIJKTCoHtqKPvobTz3Zeyj00K7Zh/exoEPtM/dej4rQyRz5M4UzXLa+3ED
3pSpbBEzZHVFxFadvbvSEKoJYczTtJqDpdbUxqiitxAuxLKDqN08M7MOIO98VdrU
f3eb53EtqFAcG3ERTpFmXaBA59AMfuN52zVvVQcr2NpB9wF9jmFSoIjIrWYepjik
refVR7PWPBJ+5zJJnlPPU3TMF8lF5Ag0Sxhjxbbbca5Dk51I9F42Rxa6wVLpDi25
VVyZ4jzyxW1xzCCptKvEPuRfXuoH61splHwaOw2HFAs6NARkucFDOgXJLtmtT6rm
qHah9nEVgw4/iom4pN9o5AvqWfPFU2YNdezP3/Z2+QUYeaqXtR9X1DFd3dI62l2X
dihcWGdssYr1w0sR4wI/OAilHsvxm0BX9C8LTvoLZosr4aBajIR83pDkubnHUTqk
tmKTAKXh5pHvikBeH701ffDQ+3Os5SHc2Ck2lQNc1pjHORaYRYQ9k0gzAFVTAsdH
ys1ujFgwgMNxkp0EPlqjoklTNt3NusbRvifhdzycBO+MMpPDQk1vDQTC46romAgb
ebGLK9VZ59TklpgGTEzh75WRMuTUUXFII/ecWZ5ys/5AIw8j2Kl1esEBG6jPhEUP
aPYDrUlsHyStFHlBzvGPIbhWQFBFAVelHHOdzhQkAnFLY4OeVJcJeUALI0e6xvsL
/8hCpqNf05/sd7H0GqF+TPFc8AGqa0Amkj7dZGhvhwhGDiB2Ar/k5N0MfEEOrCa3
UvxEJ9evFsinbQ7ucGzahpNYGAtCUiKvI0rHR/vXEBU4jvZr5KKDaDmlMRbBimBb
TGVe8TNvlUzy3q2dmKUPMMM1WQp97mgY5Cve8jPg4L+exKNVe5MvZo4mhpNmc7OQ
uzj+XuN4xOMO4Wu0iO/gb8CStuYezt564t4vJw0IykbHI4B1pZ4Ezha/67PtXfSL
Ia9wJS+V0acrDqdZ5U2Q9jUF1CSANSF3D/UiIo9HHMlhTSrDqEMx3CP1+HH1QV4g
CUOpfUFdBqzq9RQWVrADW+y3Y+zCMedRUu1prSY+s63pxsBCMEUo06fnyNWbPxQ8
wjx+DGvaHGfmPvhYN0ry+CkhKp/mYBQAGkaDTumv0aC7+iHHguYgUtTCDjYaB/y0
upBI0ZgOioXfRa+OB9HSv4w6P9jogqiwOVCtiRq/nBN7PqbI2d+LQdPIZyDPUQhl
5H5KPbTNLVfXrki8LSJXxZsjHeeXiLcm2QSzuwafCxZoisMojNmf4VjgKPdMkTte
qsiq9q8RQld7ILje1X0tMr0HB2RyA0OU6oKPFfGCrPl7LSNChatGmQyIhh2WARol
OIj4rgVW2mLkaEGJk8jC4HwyoFHJgYjtAnsLCfLFn/LX6Q+EOaaTKgRK3dHo4wqs
wnkFTXk+s52Yvc5hM2r7u2twGwcqb8JDT0rzWdmPsmTGyLuD7+BMyWBQbT5rmhuR
xVvzwL46uM/k9An7VnRGNrQ3pIyU83DF8K4wuD4Qh04YW/DGGcxzZudo7vqZCxyU
zBA/TOTdG9ImFwbT753SBJLluILQS9DY3A9zRTLPhX25HXvV9rvmEf2JNLCl4/jd
5JCa3Zax//t3qYTE9c9xiencM8X7NFR/dYcfbxCwTp7w2wjwKcstaPUG4ktpNn00
cYZoAyJ6n/z6HTfguwT89+OTCiPT5DRYBrjahG6nZLlZeSEJHRXH2XywBekVpZp3
7rQNFPs3XzkwoTOrMUL1cJ3gvpceoxVU0r8zdyF5NxrYG4Yt4BF25Mubsh+yMljn
yeetUB9PL/Y+madJVK7QQ1uCmTf9FbebiNIxImcoMXgp1NoHRfv1nVyIVPdwRnBw
o86qo4BeBB19/m5Z+iTvsn9+c26rxxrNTenYlfAiAqel1xYKMaNLr8kFgP9JjPcj
At44fCNeltSXt7xHHiEwe5SWCMPD4rHYDo08rrgcilZNSrm/MYGQeLaeap5pLQP3
E3xSpPY4fNtWCWoozPHTGcEBVpWs18oeD1abue/fpPUBF89uryYDcGhuu4cVMPIE
8969/M5qxNOXYoQDBIULSCRIKriunpGiarqVsT7IJg/7+PBy8tsUYAZ0VoZ5NOPJ
GofkGraFDgjEX8MhScQtJt+AQmdR6GoUciqZ81rDszXX2fDftGTs8Ppp3IIy6iBn
kznj4TG/BTSbUhZSwg2ugh4mdHvEqVzI/mUqta+Jqk6R9TLDvopBTOxTIqrRKDGO
EBFhxuFqA37gz/DzLhnGReCPvPZVxBHMPIABwFADthaSjy0XOVm6gOXMbxeatDb3
Gfx3WJ7STSdEJH0k/juLfLy5059NoT5wYVim/L6Mo24uVtaDnHcmmwUY4fjMwXWl
eKMgfwNf6tANUdPCcIRuUhs/IhQ8Uw0ms1snawDZJthAoGbJ945dUt4BQde8hLgF
kG9NdGN0TqqNd5Lr6ASJU8gKxn1WgnyzrqpWgdKGaxK4z20cHMKmyIHK2tOYsovj
2uIF5yFl440ZLBBbyETjVag8qNzaZRuDZvZsLGZ88iiki02s46rOX1MAX+V5tcgU
JkqBujLDVGY4zNvew6HrclXvRuTj39l+ZXRd3wwbKUKuL2gKCxOFyYAMLWZcLip9
rzA314bVoWexWF/LZ2mB/r5Fw4sWL9vd8tcXEs/v/t7SzGDUqYHQI0ub9GFgdvuq
Sa/2xkS4h3tE+2wgRtjayrjWCNQr3v5Y/1rcWSESOj2xs+Wo108KapYIFXKQMaGC
+mCPNSLzN96XFsGwLZ1rD6TvRFKT9dAzIu/IgnR/BParoqmN4cLvhqgyT3vrFhEh
n22klN2ZVbQMr+wUnUPbGDu8aQlW7PbDBAXzIKRv+fB7zVtAmKM0W3+qyBR8vJiw
g+vHZJK5bkuEyXLPF9f25t+l3v1288t6HgeAztN8dSog8ZW4JV5VKzsD2pOY/p62
kzJfUs1qCYU9zBV8vY87r+9H8/Jl3QcsbuBJfAQgfOU5ZybXW+ovOBkGnH1XhPX7
5k+UCCh9cWv2deMhT0dCDKQI3lvnka6/ivprc7qkpEKMhKp/IVVWh8yQaH3eBy70
Wu1npmYz1UzVQ+xWByefwvu15jBrUfsA8fZzm1DOf9I8S0RUsmIA2ZFeme9Vpz1+
XVbybaj/W7hvFoiInvH6gmHbhg00Y2O7DK8hA52pbiVZ8zu7N2I7zd2CNnDiRthi
eSzxLWLYot/QnJhKMSUoIEIZpds03qLcNcQekh17EebB9nGCOnzR6Lt87TucBptr
aW6KStLOVt1F8ht8OrGLqx+5mz12l3Xv+jxUAcOlv2GhRR8wk1rHdSDtMJL24i3m
d9lM8B++IIbUklmrWZu7WsMAlSp2sHNwNuXWwfr7BKtQGKu2kxoO2Ib2FeLkzlRc
XUC6DrZdtXZcbvohE4oUDlLkm62PfBUc+An2nHPhnEb0f3OQ2W5KcVeOHVJuzY/+
MnEP2LnSE42zUMknKj58CJVCjnsNiwc/BNrB1I9oLJlWvSMISmmr2heKJjiRPUDP
zIkcpMmoPiet1qm/YBQS1BSHmRfgBqYCSh+nlOk2tK2KXpSlvOXzikZ0rChJzfKG
h63glvz+jxu8Hvr/s42+u3rm5SietyOwoCsOpHY1BvVp4unndbT+vVbIqlRtc3d6
A0bkGh7TbSsm7Z58AB/YgtOHCPgman/1ld7meIsWRA3PvJUpcOBLbXGo4MENUfT/
JoFjsU6Xj86HbqarYGrLBXpVDu3eb60cfZUMmsn1PdtHcjmKz7RtjEaN21V7grhC
OECfgTwWaCX82Dw3JAob3FoDQDNNEHblGNF8WslMBRrW3w97VXFlGz3wZqSsxf4b
AaaM8Wm1vLBJSIv4sJUHyCZOjE+COffJ07JqQLs3x0++E7YRfv2C+/U1SejA8s21
2vjfjRJoCJ14vS/WORkrz14RxsU6AGDM5o0BxqbefDEBthNkk/AFZw/aAD4P2ui1
BQiI86ASiIbaqe9QKASYUWBLQIfGyb5mdMqOutBxjXoclHFZ21Lae832qyiskIQc
wKuIqGgL9coWb6TXkTsUVNwbNbdcjkVrD79NWW+v3WNhbbmaFykSkjOuAp0w/7J4
i5mN4a53NhlKcy4N4bP1c0ah0EebcVjLqMxY+CxBtO9LLqzBRvkYxfmsEdfAkAFl
0QBt2UpPITcf2gDBv2hBD7WTCJbXtg0OxzXGIDVWe0blt5MwtJOd9CJVvS+zArMp
wukflD6PKd/RbZIGnEqfYharh4xko5LFuDiCFDjLw43d+sSh1i54uPXHQZsUkt7h
Vs+0TdfLPsfcTeRWFz7TL+qbIesCd+AesXgmK7UiP0DeA0o5VmBfrWkaWETBLAa5
UWawEhiFtdT5IrJ8aU3Vr1qpsNe8jc3dv/B57E3dT2Fe0GzEC3St1mwq+dUVBMrq
KrWoRIkOPJQrrsMTDgkWHx3q6qrZxgprauQgiTo3juYnDKEb0dEApIdsgfSF5nnu
TgU24b4v0RpeGqR2U0pzYyNbvBAntjQ/AjSlLZ6CIFfrkP9BiiOUzH1teFtSz+Dt
KTPYf8P66orDDnL8ig22Y86uKXXeGNyzcOOZfHhRRFhjYljLuNxmc0xPhVKcxgvY
RQj4lpy3mWNWgo/vKPZDJHS1X7alwd/XGQlURUfKdio5gLzkjiRmW4r0rXmEor3X
6Ovs+eJ8v2r7AVag0/9z0+fb1I/BKlY76XEiyr0V6HMYqWzXpslDmzsyFY2dnkYk
F0Bbs5kHNX0SCf9/0e5M7n2/5UQTWl/ZtONEBP44+VymIGdEoJGVCqMSzgNuo/F7
CwhMWZCTk6gwcWz6LN7M3JqraNhnhLy4ViedgNkmm7OIHmttlz/0hyWOgN2m48A6
foFARPE7ohs9yUGSm1QisWRFn3ecXD/vBj1VHFz1jOhx60ncGWTYeNmiqaZFqBVs
i+NSKRbo5JIrGiJoAlS1o55AWz51PCtkC1+1qa6YwdEmTPtl7bJc4bjkjall22OI
j5koNW+0KPU/+KjfSN6AEizoB3p1LmwvgLDSvPs66dxOOGqls9GY8h0gZ0ZoTV7k
BfkNaq1Bsa32d72IWyqV0xFm1S9B5R9XMwbHOXZeq1FCfD9gVhT8JA6u/FLmsTPe
cj2ZhORTf66arCU9MKiTs+33JkQKB5THHEGONq3UZKTnM14bccoqHurXstBu14/3
1IvRAoJkV6p6CRkTNb10P8wYwVTfy9+d9etKEzHNmyUqIEOLa9qDY3k0W77anY0w
/zNb8OhdMkJiTmKxObXadGz+a+b6TqhZTKay1obFgd5DwKTozJvTUaV0W26r1h8u
e5SZu3J4epyaOA6LpJtHSvq9wLeT4QBS53pAkbyqFhKWKqjkCXJapUUHlCrGdeYX
B8vJPJjymOPcTuizeAHwJuH2XPxGZ1UlXdteuUs/Xf0DEN6ildqlYrLbh7AXEsSg
Ze1sNTN0wlILk6X6I74VfBq0FXa7fkL9i/WOKR9UvV9EIDasO7iBWqU0aqDldD4y
e/cNZG1DfLnf3K0vDTuuEIsICSqGui2ng7dp9n773nobyYyK05UyMrgo090tn98R
Wi/U/qDts7UUqb6L/qIu4NxDdAR/5s9SrfLefyAO8onY6UjYsnpGXVrA2gMSTk7H
yD22JlTjOYgjtqAQ2oYUeNq/9VAFJtmxOXwTVo9RSvtagRUaeW/teEJDZF6A1xDs
x49r+8lJkUyqTKts/SgQTybQxhS5sovPVisvldLDkPs2mOyURS6d18tZW3+0zNrw
vHRPpLxv3oLTLcuHqS2BMRZyxOZdblpbyE0+iyL1SRYhV2Qf+6J9F/567O1Fcrxk
hO+4ZOUGMnxgyrLbf5XU8WSH6TtJVpl6lIEC+4xX/V/ETNFnWVg5qimtmSZXlbFk
b8ALm/kEC1W+6UkKT2h9DVUYAMtr6S935+1V9RSc0CxdTgE2j4nqylsclSr6yuAp
/wvkcHRfCmJUGTnesOadCIraCfcKpxjPIb+GSYxffzuiGcJeSt+3lO+9RLUEl24x
YG5pO0C4XWldYwJjEi/lNZY4KGZJwHyDoJYvPWie4JuaRkhwAO0FmmaR7+NCxg+j
+HnQ/KyNtZ5+Sra7dlEJR7Dy5rzTYMGhw/c8aQpdkC0YOYLCZeA2QMyXorHX3qaG
FdxOxso0kPADTSwzKuKR3vQUCtww33Y5RnsLBUykrH/lU8oQCJN89ij0U4rFCORv
HtIriXRFNLTnRBCg2Rfm9r8WvTpviDQMIKOslHqFTYHoLmgxA4YBinT+p21uxmlt
E2cJea4Eu22xy8M2Fp+QzGWhwUya5adC+vCJ1atdHm3+JzUeF3/Ih+xhE3sM8342
utjhb477WK0fr9vB2RvExqFat0Dz64CCMC98Qu0oKPvNyetrYLZ/NHtNkS5CsFNq
77PjwGAKURq40e04dMG7rl5Cw2lqy+LNe1S66ZSit8vE7l0Jdh3FK+JykfStSZjf
g87pJjZEmkJoM6xZAf12vFVcac8WAlzFPJMCRZ7v4lDYG72oEAXPPufs3NOV7Y9E
z2wqo54kGRgUePXxRo4xEvjvh13FgUxbV1vjh353rDbQqYwFo6BTEPDODiOenpH0
7+08eXftC3Z+VcP9abPAqpvvCQh2WTAADNwzTdgJSwn3LxhmZTkgsg9JO7AgqQ8m
Nn4YdwB5cN52ZIh0yE/qYQxR7wyEMOz6BVHyc1bSZEeD+RYm7chFaW/hRLJCKYRd
Ui4G6ydfQ3tD4ASSBq1jQUPi4T+KxVtsV76ljvKAuLrMj8YOFjc/X1VE270R8ukB
2iRKNJxcTV+VvHaCokJIrbYoojX8Uoa+f6UAGXxwpilvPQPuowBcMFwi56f70qAy
e21Tgi0gmb7DRcoibGfO+RboD0m+jWRIoPExI13MhT7jC3TO/1aS+v/8GhJXBMta
oQx+qSpRyRFTYNLbJx/eE+tVEI2r6mx4jqQJV6OzMnF4OKZ7qL6AwkRvc3vpgfAl
Z5yfthhQOxxZi4sSnVclvVsacm3rWnSZVuE79V/cfds8xzdgoPIap+opCDQmgTHx
DCoCVnFNGxvGCXfmbmF7P9N6ag6Rz0cBQ601kYaITk7KtIkclK0B3vYjia8c3ox6
8wRV5Y2s5ZjvUSg9jhD+4YoSoV2MlHTb+37KxyjmDFVrGEo3Tb/IzyAiMWkVdbNd
tcWOM9EkaI0rY7fZHdG60d5UQITAfOOThApJPeCLC5Zo3pQ+vOmfaiKdnm65+D4K
JUlhJmHTRNPk8zUMd+kzLTrl/bO1tsvU36TagxGmNRAv9VaBynYhnH6GzWTXLYnX
73fWD5BTOrjQc8zfJXYf08IFjFvy8y3Ext5YSiKGfo0s3sI8JjdsXmqJouf5VOAj
yK3Zr1A9XeZN6IRDJfbAXtAuY0lMYibGKBDdvgKNtNke0HY5PiXxE8jxOKjwF1IH
GiHCPwMjExQ6ZuSWoENLdAOycC5csK0YF6dwZTFTl1/tOcWRZpc3gLwsBzRs8A11
fdVsfmRxNj77XgEDEM1fAAI+kB9ZwlBRchLE55b0MkWrqW3JwnLskjqH6JUktnnO
roX5LnCcFBruRQgFL2L5bWUr5LpFHZoQDAiTzP9+QciOK9sP6c6v6xPQUHsl0ABu
MVIUzOeMxe8zEFvF86ec8BqqQLwJ4rrHai1Pwa/PQbkkpaBqmsB6MjhDtEySeFu8
IVX4oAON9m/OQL9vRuk2cNtMt4EOVXBUvlU7GCLzWGYiLArFrewUM9AEJCu9Hw+F
xybgdHubb2xX+C1EvMVScMlVpapG9CN/UzHWXqcyb3WkiwUD8LT9xZw8+apXfpKO
zfO5n2Qdst9cQ+zIwJlBhpKaUvOArzngFxo6xqkkZ+A7pctDUgfToHbNjiT4n/88
rO/gy23z1PudRLzSTks1D4U5LI4H6mEIZBwdaOXi8iXtZUT575oXuh2DD9iCq7Ii
jtQ9iM10jE6etjcBz3JzocKZmeeI8cFem+B+QMGbiMoqBXfMf46jFr8BcgbX52qR
J4lWPBSOt4DIeXub88FqazUcIZ91OlSmGXfZwHTlXTHOTiRKWsmbKMll+XnqSlVp
1v5rllV4FtAVxU4e443sCWbB+v8IpGC9uvCfWfQ8NG8F7ASglsV1JkjuqK5Ajqhj
KbXmDS1UbiLsK/f7UPxZRdKnTnaceGgtiBgiGO5DMRBuMeZ1N8s1gGUDjMOn539k
2OLxS1eFYLrAEIuXTmgqi2XOjteOTZaha3iqGuhkaM3SatRIYCZcsMcGCGNVTO0X
+SpElygmehAPNKxMCXQDbftQzCyS6m85qxTEsM90anFV77/ghi7xuTGm7XMwnbo0
vOCSW1THV6MXGqAwHO0kIixas0w3WfYeqWKUBlDoOnLiB7YsNqeKyQcdg2RT817P
iTAn0sS8SYVGfnQ7n3GA8p/CpXhRIMUdcgwIr+UqFdFm2FsetkamCOQX9VApyWTG
rbA9ThM6B8Vvyskp+gD3BtrU4sOVN0pNNpY826nOWhISZmPhd4/b0Eo6GQOz3oF1
mqN1kWCXbEDPh0fjudFzya8iSaw+IB4MsgI98Lmkj8DBho6hTMS358eAAwGHFeNO
jgDYNgo5JnqMYfJWxeNYemk5sWoERvtgPXi43erZGENTvlbIXbSCsDHYo7e7pycW
pQxomIlqBtb1FO9RANSxf0K1V6Sse7M4hmFX9BmYNf4KyZffhOOygfn8SMMskV69
MY9CteAqXZb8zpN4ogr6YhRXiIgOgVBmd0WA4bG5KJl7QVgU1u4WvtWuvsrQcrcP
/RrrB6tWgcCIyNRFqyEmjT8tG8sctYVC59yG0P0I3YAuW2+nJTsD8HDbg6juPJtD
rnQbejRRKkjScrATZQahGBok+nTcMYyTZFn01IEBrE9gvDsmQsLkq4KRn4oxiJD/
6IeUUjqlW4CDF6UBa8xYzS1Lqi9KoGNztRSAXsLc3/+8ExbH6T+/B27VsWM0fjKO
0mbYSBrV5KJ+ec48FKYjVfYnkzkUSUIQwhisDW3prHjU0Pv48oben06qnWJLuXZz
ik84i86gdv25pdt9sJj0VjPd/BRq8IJGcvEYdZri/5cLhXPTSdak4F4CuKKmXzr7
X894R/27nAFsK62OnWDw92+TqSb/+FgBuw09XMXLnib6mm7iU71QbuQ4ISD2fWzc
174Ub9+jfddAh3bw8Ij+lPEEFd9JnkmlM/Z8T87xcfSxfuGm16sMNZONQQYl0+7h
AjiCrNiP8qEUWWZpqbkF2uwGfz/vOKFbrPhD7+JZsEQ4n81ACSnvXZYDkXwXBRsK
Acsd9tX0lKo3W3dM3RHhfyGnHzye5zALUFfGgFU2dqvobIWrS4PTUL/MoHQIOfH6
Vvq+r9qkwCzUingRs2EnIYa0vmfckqhCBe8q38yJN+u62dR/I37BIZlVy3A4/xTj
cp7sa5WlYetyUz4y1Wetuq79YyX41icbkNwbw638XHYIS+rDOXGv//OlMcTcnwJz
ret7FocpLhmfzzSOUkhlVKtzMyFfjC2NXQtEqlfHXEYgZuY3ae/zFFMbEZ2Hf5GY
+dACxuBacqhY/xsRdy+GNbvDR5TXQgx1RVaLM2aRmrbPfjJYvkyaQGGPfaisHd8F
cmGKxIrOCR9660whXP+bSi39WnivfUu/0uwJtaxrA1u97e7NJOpmwIrI+auR7tn4
wGnhRzzMZkph2DEqRAu3ghxpnxqG6Bdjtc/Kv94GYOYJieNDrc7N3wcpgiflhYh3
oRkgEHM15FRqTsQE4ljsd/1MRjpc8qo8KN2WnxeB/tUqO6hU0ca5cAphqc8AK5wt
HCuVba4bMfWYPcrB2eUwLKABpC1qUu7xvqACXqUGn4/rfUZneRJ/ZUnHkVIXnWSm
QRubJL6af3VxEGSn3s6umNB2vBpcxHO/SK4R3EwdYO/AOmVsFVuKeNMhpJAbB1ly
9vrCUuJL/Xd/Z+6oGzoh2Q1Sh4BTjQPyln5bPJFIQRv9N2ISjweZeIY/tfomM5XY
naJU6YcCO/oLWCb7YxZc00Kcazxkj0V9dowAYCTDVnTMjccYzlpJphI8zM/0AAdR
Pm4V5EHEfKs63piZfujer+Bbg4u9s5KvVCnsw7nYN+A2c5vjcalljJ1Ar3I+NFBO
nGJB5GxEZrnBHMTXfP/os/WEBJts9gQSfvkaEC1uOfAXpoARNLM/IDlhAjvL0nik
GYrq3uyCaFS6CT5cqHHVSqc8zKAdR8DwG4pobNjP3a0XRvHjCgGavWbIW94GKGYV
0VIn/mokvot+/IUl5FL9cs3zEmgbd5QgY5v+Et/JKPiEsdxxPzhyXBMwnzukeS2F
kGpOCVNZLCIqDfClqLkaJMqfxFZkP7WgHM8Oxu3QaDmPC0GiA3xCKHfUhGzkXCt6
02RsRsdrEfWODvQc5t7ADelLM8ASjt9AV4V0HbkXeEdp7mQVINYW/RcW4MknkBMS
5s8AwRkw2u+rFFi4QqnWdjBdt8D3iHAeaGpkgs2zdC1xFXUAQB8WB6ftjsAEsTaC
awUzUFROpFqaUy+AQSLNwBDlCwZOhGXglwj3zTM3B26U33BpaenY3fe5Nfl+jC/1
KkXz3McRmvtw8IqMam0cNKJFfLxikvpJaV+pleDAUHDhJMrl8zE6ozEbZvJwiEkY
5NGv3j3afJjzgQ2XtFIfpDeBcoT9Q9qDr2GiXLEr55Fi+hCKDBGOU/P23rHje/L/
WMpCdx2XILnvKgqojK3bFNpnXY8BQFC02Am2HY78Fca9MUKHxRi0sR85B5G4jj/I
oNKbHDMJlCSF9VS8ZHfY15TOrv//9Ny0FnpOiO/zzrd2x6qNjS3T5mGg4Is6/gQU
/mw7PM7atO4rJI2/opmihmgyiOjkEY7vj0kwLbHsMMi3F932UQMUFFKcya/sZrWC
MJN4uz1lcwuIkTiaPuhHG0IS3uxv5DXMtH1JT7yLiRAjGf0GzYb92vdr/4tTkFye
NmNmas77yp3MSnmwAGZBZUUxAYN+0yF1YpUUIAUzbDxFQ8xPyZ6csTlFCJHxHjj0
ozZuVwQVRixQg/a/2k5k5S9CZKwKoMRcDoOfYRM1joA8oj7SlqqFE/jT8579YMEo
D7ZrWyPW5NG9GClNk9cHb2Mw76EKWn5NnZ5ypt2642q67F0eabFnnrc4nObWuRXL
erRG9A1q28qq5bnAuvJZMTmCQvCRGpjyu/7ZkcbnnX9shZ3LIqzVL+PPjkm46iyX
ujnWgVZZ8tLjqsvprJ44v93KrvubLYASskhkU+fhhMmaOuU/SbdQKnpa48eLm4QN
QkaF5JooSceO904D8NiH7Xtt69w5zSkvRkoaeWJbzmSbmtV3z8TF0fe3n9/AVatg
+4q0jkauVPxja80Q4WZCfoFd03nj44DPoM1kVPbzUnQEvUR87CVrpW3Iuqu2a3nJ
mlL4YX1ekZm1++3pMFo/tITyVe/L0wAdeuFLfdnzGinaGxa+PhFo02lDWVMhyFbq
F+Hqg4wZPBY+DBLQ+xkYKIkv7zbNgg7RK4m7AZho6Yhkak3gPVZ20ucgeDT0flzi
YOI6e42McyTNxqPAJGPxqcpnKnSG6rVnGoXllWTe7bcZgG5vsnPs+keEQGimIcF9
x1qcbBZ0XxcpID0hKVHkCfwCxu4EcXMlACuC0mDJ2/8yAhAeTeSeriqDdrJpWgpw
d/DYOupX8c+4DCZY/AxC2sme08HPn7n1rrEIQZPMd21rYcfPA06gyrQ5Nf3Q/aha
B81y7xYncaSSBmD/lgdCC9alWkRQh5fwU1rNXsVNhwgvZm/56OmPriqCGyZKBNC9
CgEhHFVZkk2Awy6GMIF73d4UQTn2u/nbSC+tBeAElc7EHKVdEMFwNxobJQIRQqyq
3XnRk8C+iO3kqH/vBG/feKhN02D1SDSDyoUYbMCS5EPgKWmSuNaQ2DuHb+UaixKL
wh+Ik48ijXfV8A51dnGWvhc0EXT4bYXsepaMqnAw2euVaSYWZcydTpFidxn9GWlB
z7iy5q3PPRkUoUYdWXfncaEEwb9YJ24smXMsuGqpEsgwiD5dBMG7+axLer9i+o/u
CoeHzpfkXG6//N+rqI1MTZbFYCYkJBp3nO/dTgO8ajHCtOUEJfH6lsKVmJJTGOkL
h1AXcGbrtNBgTln+lnpHeuE4uLL7qY4g3RZlDgCv08nm7ve5X7v2OuxgMIa9/pnD
DDGIy3lbS51lrt3xmIIp7m6qukkL89DBsJ5JAuDvcdABv6BRIw+bhB3LT90FG0sn
IeW9o1jSUqzobUFVLcEe9yEvojgmgfsbHdGT8tN7my6xc2DXPrQDitbsbOkm68ao
ded11nXp1kCIoD6oPsEEsrA2aDkE/kFb0CnfQp503Gq4L3abG4zSs8sqR80+qOkw
RhhaSPV5c7cDnrpHTyICCJoi1ICHfH/ar363W2jdz+f4ryuFKzyLjrPDtgy4yfoG
UMmbogKBsZ/h3BIMzIg0md1ZfgC/Dl2mwF7XLZwLLWwFAC64evzEhFwKDJlhm5EJ
Nm+DIgPSMcKm3D9BLffBQ9Lj2ooppDT6gH34thbDOLmZjQ/Sn/V6Ji9HKUE+4XLv
yHJxDWxO8V3f0NRh1hT3VPI43T9Wxnut/AaEKsvibPQ1N80piI+bnWRitozmeICL
g1DXjFlQb3GaonGQbirtiD3kXfaGR5QMD8OiR8q6d9fW8I+Bl3RJL34bCx9+28Te
njCJQWB1skPsjuRFdeL2a47CSpUd9pCQra20zi0OJ1RG353zeeN3gx7dqRgV1YFT
BiDrEKqRu5CX4nLIjW3Lc0mraurrQBqp6XN0PH3e3NjgYRx/ZMFJEFxm/xiUE7I5
lqDKvhUlwCa6FFWNzUVGptikz8NyoJq4tIFOkw4HjRxbsG59lxqfMPy3K3uUTQP5
jjd5VRIqrapnV4sHdIm7WodG6MJXto5cjgNE7ACStkiZps8fDkO6fhvFOMXSB6D5
NgWWVdynjHEodT7Pc6rNlAcKMZKe6L5pByDNRd/0spttjz1ni32AlT7AfJONAT0c
3Uje/ixaqq7fhGAaPp9bDodGqwlo69vfjP7KIT3idaQ8ylzEtDiuTP8aFLrA1BIy
FWphVZSwvP5/b4lZd+95EJOYWmUqtOqZsnbRkOtlzSP7Hpjue2b9WSSoGi8ZocT4
cQF/r19prmIZs3x7ndsgQu0f2Kq4/DW4MKLc6igaspgOBSr2eTsSLY/pHAiyTMGh
jMXMgsxUaeGVfoh9/JYWFCCulyzZTQTuIYsCM8VikjOQEfIrZhPmH8Rl5esDF2P0
/W7hi/MTPlBsh8oDLz+rFu0OEBdammN46yPSfTlMJ0JCBCYLF9+wWbg9JNQ5fYq0
DfgRhhZNyRdA5oEKE6qZAJD1VVgr+AQZ9Kt4dBrMbUFpR21IeFBt7iGlJ2WE2Cru
+S3n2vmI4Pwql6J16W/5pteXKN8CU2zSpY9dNdGWXllV28aZJXoB4SwRR9H01o6G
L4ml48WDwiNuPFVX+cbGI1XK5snfWOJZweZZ4m+V5XwmVAH2llvcB29BVERv8DYZ
GyKB9CD0igDxZzwlQ8ujHMxarxf0PHJPytbFdEshvLmnXzRyoAfpzM96byT5dE2r
3stPtKX5uW9jevQsOa12fsNC4FBNnqpn4dxufjDE8Ozd3KOgCXK+xgqC+/iIypx3
VARzQzJiDotQCkdxxTei7E/VvxxrpkDoKRkQHr/QFidHMubMqPP+RKZj/AJZPJnN
sZLxFFJEwHpF+J+ZR9axam2GaVTk/5qBSOJEE1fHStTqdzoHwEpY0+SqgN1NO7QS
RwtzNidTo69PJLRGBz+PftEKCFSUb7zLDXFSLiG+SF8maQnn8+8PjOs/zUcLQMO0
QYg4ua1+wCMMZesWwgCxFpUSoa7i1CHsDN0RPef73NvX8uNlv9DAGbqYzDgEUSXc
tmgcYbZe6HqGhsXkoqmyBQm8tBEoSY0TPSIUrDnJGXrpLLj9232laxJlNqLwK/8b
cPgnt73FIt2zztfo4otjNWZMALogfKLEMz35Ak9oNf2HyiV9wovpPhDgT43mevg+
T1VA1juK6RTJaWij69GzC8xR9R9/7TEuLxS6B0Mf3gBIwYb7VmMqy1vCXn7duHqi
/BXROtp1/pVP4dj8DjBjTEyV+diPNjoKOuUdWvzsIquYuIObUjDhmpE8+za3K51y
CkLM0+W+RGjqJykYdNDnPDWiSnD2EkE4dlIEiTZaKkzy/NJy+9C2GE2dt5C55Mti
TUm9t7UDRAdp7sjCBMEzrmIL65VPUlEbtDwOCjBYWeCP6JNYB0l4pUmsMspdBxKe
R+ybBWEqgRKGA9Kd7d8+6msASKPQEoIeIL8ZWo4t3Q63i/n2stV1DV+2qfdnDi7S
vAq8v9yS+RChhfPjHR9ZIn7Kz8JOGzu2w1YLyuejF7lZ2rHgIPniOPERGpFhsgL1
4GaAyEZnUxiHBonRGk0wW7k3CLGH7nadqIrbSicW5V4nuZbfgD6tSB8eROaZ4yRk
+VDcWSvatMDb/k1AiQzTA2626P8dv8po1n8ORLK4jgD9nBxa556CG49srXo+uTLF
+b5mkxkXt50CGr74vWFu0BlUJtHUEcNAUDZ02mYKLafYo+yY+N2NknzPm1gtJFJo
GJPvxJkZ6bnBPWkeW6JxCMoaYSnPP4YrkX/8CyY64KWvoOTHxvMqbrlHXBYSbOsy
W6cMoW1w5KgVBDbPa4dpXLnPnEGd2AXwzDfd4Pi6RCuxC8oGke7yp/60kywNOFg0
Dhm34ZrpEMzxHI38qX82kAit8xSM57EHsJMw39En9iv6UA92Hxg/SRvPwVzfAv4D
zoXkpYtBnUkJ9gb2m/lkkwB1QoRM0Cfg5l59mS3G6szpIQj56LpLasnn16zDw2gi
41VOq+KV8QTaG1RL1B5yYIGjEG4oSlVhptt2j/OEHxC9b0NRIuAv2hF+hJpG0NPc
0ZqtvRcljnucLz6D23evhw0Ud4yl5KedD1P4hdGUnoYEn9oKE8kCUlQANjwEEWB2
F2dzciZ3AQaIc3T0guZJ6Ey2z/S57AA+tQCsgScGgx0Feiqoi1YqW5iMBPezL7WC
BUYHkzoijLkj/emttG+15B8p4zliPG/bLXxnvLtCRtNveGeibAgmutOBmhR4DtS8
GxTMqPFDOmzurAa54VNDYCL/MgpHIYO10Wg4j5Al9n3Y5jbHJ03KUD+4Zrf123SD
HdXbR/Y6ZJdpuBwV97YuGNGrfoqZqKo9Hwdl4PykaeQuo7LAU5mnupAJ0noXGicJ
5lmR1LL+ftIjauF0RCQovk15Wq/UE9/T73/1qXFeWO1IeYEv5hAh1BkWIE1UljWT
jTCBc9DiWXD+HZxGRrmzi6Pqx+oS7JhqYJY2aRdRMtHLGbfetJO3oQML8uhPDYmL
69StPs2mBMnEDTDgcKEY6T0SOzqMtzPMN0y+K69JuCXkl3SiPBvtAY/ODLUcC+/M
IqnhcUWHC11RhCG4T/8kfk3rAMFhjdJaX69IokQPx4JS2ZdF5yXVXd9h4/wldYRn
ICPb5wdFfH5yGjsJWjpuEba7qUTQhpR/R58edvWme1M+34iS4NOnL9XKuuY8AtRy
6syg4ApUOayF2gLWq3AfLhM2i/W6Es0/9lhv3FpSAaP93eWrqsv16TUIEqtTgJgF
GWi1+LJJgZVQV4rzTf++NzUljFD0yR7VemQknaHQfo3Zs747swqr8qghZkcBOaOT
SV376kOPezp3tJa4gZyBXYr0EYzEUSjpsdQCQH4wXVj0NxN3O2K5xIdA8z8hYqU6
mAI0H/kFZ9WNUQT4oY79oQ9vS8DItxJKrT65kuuhsa2NQyD5BpICU1stBIZTcGm7
6GiQFAy3O6Q5Fw6GeLWtfDR0AxdOEOjl69vKZLbqiyS5edL90QunFh2c+a1t0DGZ
7Ot/JVzejwsXNOumduGYips4Pp7nFoiJZMpjfLvumW8OGXCNqRr0hGrFjP/GsPvl
+k0rYb4z/IvQaz17qrWQ5KoygjaDqGVwHLJdczz/N9Cr26u2xRYxcQ8ZFnuO6r/l
o+hDbweIf8eIYftT8LAqwqW6I0wyKbZGguQFelqV+H7Cw6DkjjnHcQNN/NGsLfHs
HCbrF0k3A4M+bK5qkgTow5TaQ5cqd9biAiXkchBDnD61ZNck0z1AMZot+aA8y0dh
2ID8rcKJyhwHTuSOgSM50sgT+PUSwIcf3hpmO/XeaNoRJ/0VBPmeNdqMWr/FNHDY
M6IX2Ss5cuhnaj49dOLjhVS49+VMa759itT6AetWZf99s/TqqWsi9Cs1PjfRz3Vq
DPQvXTKn5sYCZsZ1QDE1iiVd44a/Lsy8+mAFs3JmZGSkaP93wENwIO5Nf7+0KQDm
FUnOLi2cfSpQ9Sr1wkiCbYQ+7PSykcEhHl8O/fl/HU+/0BpDbOyT/9kQNPIRLB2W
GrD3n3mSOPzA58+WJR/rjHuDnJXctVJ2QWw7pz5piOHH9wwXiSbzfO7abm9us3we
H4a21Yj+7FeMrMYxeZ1uJ0F59hk2AxGCcYyKbIijdEJfrvG36BSMP1WO6IlkdwKc
XG6Vj+2lWtqfbC/LCbmrJZpSMhSlAXBgY+jcngJAWVdA9Xi023ybB9uM+Ds5aF3B
iLI1oUnqPH7PHyYsLWyhZyXwLtA9hsUHAp/wqBnyeqA/LD5Vjh75zJ8ss4yRsudo
G3OPcuckO7YbeGRDXwGIR1wX/MbrubiwQUd9znHpJY1jG1uHzy4Xx7hjFJUkW5fF
GYoqlnYUrE4f10ZNpC1JXUWpdvhuDRc8Y4hbsvNj2wnzU0fWW+i/dvpu6G3A8yJY
h0q4ZF0fGm8FGbPyraJEScTiA2ovk7mqwFfyMYy8wknnsfEJOROrLLCPpnZyePEN
fo46G2pG/tyPJnSnLKcyD9gFWekF/Ac520wGQpGjVDzFrNcqz/BXz7cE4pReh5Qs
Ra8o7fzm308uwSBHZx09+jpUAIO5NC1neD5N8UiO/ccmszg78Sn873refYDEJvvH
F9CLwLbthDjNy4CYO3Fi8eid/HRd6GENFHopXtPq2zHOdAMybuD5c48I6VwaTck1
HrGDbGoq+UOtZnfV2B8hYK6qkQbIkdeO1SDRrUYcQIcqlVqJ4CsMkdPWJLcSGA2N
ECcD/3IrVoSRuOS0cgN8ICDXrmy9KEUe9zcevqhVi4wrgrv4cB2rEVVXJpSntLhE
gXh4mLgdxq0QtHehT+rxK26fP/kLNqIKnf3aBMM79RIj19FXcEYsIgl9hQTRL0v2
CGW1qbRK+1F+YYeIjPfLtiwi3jFpjaBmt7FrVV/oHublnI2jf4nAopiYGLJ2BwaV
t6OaR6rHVjY0LXKebVZOM0ktW0c52k+fkhqnBJpQDym6O1t+MFMjwEXPQPQ5hF8A
/L/PsGmDHkFwwMWTz/QwnooSBCKrTcB87KDmO9eU3anOHWmY76+4d42rhIRdrQ3N
YQ90M0PNgLTNPkP3fxeQVzMj05iBMPdHzMLJQu1sIhTJJKc9bIoQrXgQl34Qfg5k
mANDcYZjwd7d3OVR5mcFA4BXiyyJ6QH1v93C8CoBBWm/DlOz5DWQBU8K5IrzeYnh
WZLLrgZYOSaHnFgQp6aHC4XtrflbQWHSwwL1hyFxIC3RuC8/4+kwEIeAQ0iJlu6J
xIsVNVymM0OP1Wa8DpMu9w433gRmUo7QA9eJHt8a7HIN9NyT4Zxkqae/SLVoclD7
cuAAHhPSWSVES2uWXvQHEB2THijQc+8qQBBBOWpm6Kpl0NbcE5r6uhkY2HUxy8QR
ZxAHpa9Gvs5NVJdEjnmcfcl148q4UNGeh1TDxd3m+sMkDt5DrrNe/ZTeS/uCy+/x
XAq+iWF243McfP6n9uAiFLUbW8FaJeOR1sw7thDgNam0UnflXcYtjytBkyNqdodM
robH+X2+GzOtGhOBcZQgmEmIzd4LxpOshwZHvksEdKhQUCa78F4b4Dj/cY1UdzQY
4sguU06oChs+Bh4hXrEKlo0XanmxR4pyo0chp42EWmLoj9HuoM6QwKc8iTQ+1H2C
73Rcp/MhYHA59WXjgBZMfhTj+0PFxkQXSXRqE2z+aH3mzD1RiP8eQMv5uB4qw3LS
Ydp1ZYNrEG0mmjDXVwg572cIX9Sye75ODai9XIFf0kROUsEixnQ6kwFgF+cFc7sE
+YyotXMSi/JR2xv9TRrkY3cGZzTCwkFFWGbyE3EZTJ3yuGOs8THkD70wYxB2zqiN
J8g0n/WEThgqrrX53mQuq2kFhkscSrBn62/cstNdCgBwVpBER49G3p2RBCZq3Jk2
bdEXDeyVx/AfyP2U54SkqgZh89pySTOVbhOElDleInXvYsMUEZDNI8RkJNZY9a5+
9DGG/OuwK1PLX/cj/wpoMGnSfZNqwv5E1RPtQAEHZnsVjrlLQ8w+9173tgY1/zeN
kIl1PLYb7z125kLqEJ4zajwERTV6gSmLKhw7tCCkAeQfmq1UezdtGe8pjHA24J+K
UaNaTPRAdeJO5PHVczYGW6CEkYUU3SN4ya0ZjEr1gj+kQXqZJORg9IBCJOcEDzi6
+TC0ZvkFRlUaQfnRHQdCdLTWTYthzhPSJTMjaCi/V4HA3s2Qi+xxg2Q1OtGzXTuI
MFHYh80DWqwJbc58L9h2L/f1j6xFQY46bcQDgQh6LwZ/4gmMdIqFrd6zvc1DMmvn
jDOi+hz6aQPOCyMnk39sau219jnuv7m3N0KxYvdezxL6v50MXbt3bbeQuGbec7n3
O5jPj5/sJGfZgl647EfM3J4UULyvFZHIs/cDM4hJcDUlaUK5nFk9RAO726lsJT18
cxo48OS+BkzqZ46FHTimFImRfxLikLmJwtDW3OzZwFvwV8Aizw/RO1M5MoJNljBB
x5oaovyIEqHAs83IKEMYEKAxDME+RgaOFXOu8nGpL9vaBb9mTmtTvzPsFHAbEk9q
1ckJCpiPqnBH0LJMD7fDcjBN0PIj1tpzPar5iLtD+R9ejYTGP9csd3qJKbQVy0UM
NGdGfkihpvqR84q1dTWAzdq3uHfx5hcAVgBg/d4EqL8r94UxQQWFVg7hMvPlc0vp
ZUcPjRBF6xtQpkL0+irFCwQT5Aetj5JqbNO2bFo4B2b032+SY/uA+exp2t/Xo/Dr
4e8sWpc3jhblsaR2NZzuvA5g6PxPlLI7d/C08zNS9++R6/QlV2Zc/8W2FnrBvW8H
go10AvN02yTDvRgl26uQXE7alHnHNkOdBlqDgtFk/+DLIABOVQnOeQK9HCjEHGM8
zxWqnsoisgJ6BfAHoHPBBTobvRVRXDqlM9wkErjebwsfSAj0xFmhlWJHUd0bGRlF
Z1VQNi6Nwf/0QoGBx0NnUFI3C1b0mBSzkHcRpfWbr6p8EEAmCv1VBh7Yzez/nfQ9
v++s7CuJEQrEk4P9c8ZOUYnmaE+jyoW3RIOlIGHChDZURm6XsdsijCeBvnxWL/v3
hALqcauqgVzRWC4LyVy+bqMG10angy9grK9EoQuGrwTHLqRvbRw2PDu06op3YTMK
9yn+s02G1TbW1As8Imrf/GnQg4rSY7oJZSCLFkKCZE3O8X6NHowD6SgIAnEpiTdw
PzHm6thEprTFypTqQ/THIe6Q2Obe8Zdlh+we6IjZs0pRLpjopxCMGqgkFaxVV8MZ
Uk4iLxLaOTOA1gFxDpdFutff/w8i3zYI13Kqk5A8ZBBKPQQ2JwzfTTmq61Qbnla2
PCP8ub+p+sLNABk0mYpPlrGnfXp/nr/S4nrIio/1diIyduQz41niV78JKa+iGmlQ
lD0tWr1eU8MiKTAGamDiILocts1D6+grHZJplUOpTIjarIExIxXvHbWQ+FSxcbto
P81S3m2PS9trHX9qpN+LQq9iqQPVCdmxO/oemyfi5hQEEf4Z+f4gCcGaqr7KR+GY
jkjujKFiMgHf4SFDydA1sR7ufEf68futfC9M+zYiKUPVta6hkRhtPnFwSHQC7b0f
xw6hWuPLlMAiIvSB6S9veVjDzdps0c3bMxMz8A+mFMHjyhFfslyOxLXpP1sObW0j
DvnhcqTXrN2Ipqe+8GUDAwEBqNvYImFrEr15+SAkcDaWBf4dIn0T09Og2XhGLvRS
5Gsa98dHeASDpySTIQMtqrsetCea+6uzo9avRtrj7CGbbBlQe6zdwbpfazluV8jW
4cqrjXRdM1RHoDTUUbiQmZHK46m0lKYES5MOzIofcVKZ4XJ9ogVXcpNJpuiu848l
S0IURpzYFQe1i9JiuFTnwwM3B4DkcH61vZRlXOc/Buv1ek0nHuBGEHhQPg7MCH1Z
Eab3V/EUo9nK9+1EtM2PRCVFJMvKWYzJqROKMGfHwtempbH32PP4ppZ4+Ddh5Inf
EZoMw4p2HmlWS+jb5bUKV2m5aly6K2+O/mX8ocAr5yF3a+L/ZhR8LKzay/nttNEN
J8yDSdaKX/rryGGqWbb07BAFD9X9D/0XVDZ+Ch6uUHpvlSzIcF9FlkY9vWA6dkhx
tlDUtm7V9ct2cfeUH2/tPAa1BDkqZdh7PwqQfIroJRaoSYpBM8LVlvpyQ8eVhFod
G67BEglxvgEhHIr33An0KuWybgAXdlf55PHU2SmOvKlNtvkGbGbnBDXCUicfQ/nM
ReR4bQ7eLYPxzqAPEYlZT0TyuFHJqciDM4Mr29FV+IvJA8ClOjP1ywsYGcgHmXaz
NyH8pA1JncotBDeh2vET3PsHhzxk9z3E7EzQ8+l1Mu4yZ4AYdpU+VvHWbQcxMB2S
90+pVxRAf4Chbqop6E/Rnzd+Vw+3kpkWhkzX/svE2Lrn+yWHe8+ePrDlDHopu+bt
RvmH6Va5rsjHsImJuFlBxODO5ElwZs1bt92uHfspS+g82jgqD8xb0R5SA8QletRw
SVKAxuCsw0w5ZNeortVtMW+8ugDF8Wnh7X86k/o9IfCvX6qYdQP5te6PeGgGOWqn
eiisFdsK4ORm0ThnF5Z6U2nCLGilQvx1gn8WEvz+KGZH5h5zW3JeFRwmsaEfNuPp
EwjLkHrNuNPnKW6krX4fwN1UJn7XJExGHYLEoXB7AebkfPG2vDCOIsc4RswSyn3n
TiFFZHOz9lsPM4zE3j/CjpfQiTcC/3Hb6sEwamyHZIjGDjhJOuhCKsTopKCaew8n
NXkV+N+NF7+JQ8ol8HMtYyrOvZLEcWPMkDnO4RYqPjgQ51eKAtcyVy7msPEs1DQo
uZNUHZHB9hp6ThIAN46b4sMKY5HtYXUObAQ9URejeZpj/hZPNQ1bsnjyM2L7/xul
9wq6MlfVGvkAb4wA4Q9DqLg6f94E984qXpqFBA5+cwwlX/4zLqvDM4X8vHrYlHmG
110UmsWGESSchi9G5f/yFY2A/lC0OiSz30+UiZR0rHYLhL8F/ugad5dVAX7YR4PB
0N8vdVTymLyQ2uDpdfAKdUBEYrcAJxpWBlNSq44/o+ja3c1HZlUumDaSmtsQblb/
lohtT8A7QO+FsL/MWtZVOEyJAPeTwQ4ZLtDJVnC1iG9f0MQKM9vafdqiLANm/m+U
V+w70cLCUpVjxV2FVz5X26B4PdFjIhGR93dSuu74TndFln2KMc6w9WG4YVluTxuc
H7l0AFwjC4n9tu26v5r2v2MLFAqgI92/DflZsXtfH3Fn1y9yZkN2YKqRe1o8l/v8
+OUVrhS+cJna5FYt9hRlQYW6fDPwr0pV76iGDVY/SE69Hd+eaTGb1+etifHuNAY9
q3P3WL6YRh/YP4Im0870j2HqlJCPPx42dp4NqWlhLbqsfG47smZOk9+/XTckTPez
G1ak9soj2Oni9YA7yYGzFMnEajZb8IOoTkuojpnwBW1zRmTuuBv8eEPtI6U1L3nJ
JDPrU8TPUjJRm4dtl1iRgozFjTKa4gW1494EwyhAMcEMKtOL9oo8HsdA7/uUEPP9
XZ5/41WMxfmpB4BimYFYvYH1zqziV8Lgl873SnfvGlunA2oWCEC5b1TXGjD3OzUu
Q9HefTySsDfDtkkCFq3YVTS03hgfefF3hA/b8VA+heZMLmoYJk77db90Sp4/0z3Y
riOo5A7NHtWD54Y7z6y2bgkydQsmSqKZ0gCyL9s0daHSKu6N0GjmgFXXrXRJAEVb
PNQAH1mJjuHqIuP9vfjs5A==
`pragma protect end_protected
