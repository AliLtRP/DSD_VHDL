// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A187Ti4CdQm4lZvaa65bKDVQSRGk3hDUXYwMFQuJwTcpc5lE9Buj27FOZpcVgxUj
Pn3nxH3U0igL9CEFWFcYZ5LPb1Laoyv/trztILFT5qXl8WFkavECWjFMZFqOUlxg
IDvfoDX17nZVII66wRJPSMmbL0Z8vPvke9d6ZUl0zEI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24624)
n9loskkPa4ofdfJiMxMQzAnzPOtW+utc4w2UuUuyfzkZkaZ4UeVn0HlR8H6+mGEp
V4UxAY0GyDZgyzcL+x422IDYB27Sdjw5KCbLiFQMhwnTQedJUu6rb5pLJO3gdqao
ix0y155y3aINupH+PeTdFDeZwvb/kOCFwd1/u+3Y+34mTZdZngyCHUHbckjg44OB
KFtWZ6zgFGOhMsRRAgIQHFsfKB8Dh4Fx/Z62ehPrSj8rAL43Se8WBQ1bmKyy5AUd
iVQhqbdVbv9sW6dsi/OzHx8xAOT0pAymDGnwCrgni27XkJNLeg44WV3mXdI1XZeo
cmUes34aP7ddZzLQ1prlVh2lDmpMlopjx/HyzGB+KGpv1SQ9VepdVdCPD/lI82dm
FW8m8pR/7GipLIr6DnrLfX1tUrcIYbTBcgMxk4pbfpL8mt2FnB7jespprKOwuzln
aEBOxsGqzj1Xo3sFQUv2+CUJirWJo1Ja8sC+3EBcC7YqJmZe6kuRftdzwJhmNkSM
qL3EdmzrYdoF9h/25p2+wehOtHRc2WsNrreI6wWyo3oi21skS2grwPDZpwXfjUMH
GJ7GKSpP7b7TPQpW+x2wWkvrMBQzZl84U6n0xmIfTP/rW0Daq5F5MDY/OypB8GoM
0zOItfyEolxiJOeFh6j791Dcbfttt9ktfLmFK7E7HYix5pccLArmgsC/JeES9sDe
4judbd7EHYIx5sn+WQ99gpGjLKFZNd/pye8IaOUasEsMBMi0exIvZNPXAqsTD99l
WDfm2Yzmpc2BnBWpN5tFtUMTWObcfmt7RpQxdUSpWnsyju5YDUj1BNvLvgpoKOKo
hGWsyyi8+hxvqpUnWZZJw7pkKhRCjvlUMM8VWaTUk1fIrCKDgWfpfkLmoh50n5Qn
sNAH6cop9QUaHKdMQsP774MnLdpH5nOEJYdFXh6o1xJaCVa6wuncOyY0pdMmeyfN
G3s2S/XRCr9bX39oaa4qcZqswQEvw7h03RpVEJisAlHPLsYBrIPGbtNYFxuszjyG
JukAUDMbCQkS6SFrAZy4zMKZlgPTgPA6bIlMOStNa2l2fA7AZyhNyADFgIo26mrU
gfbQefwXZzuC81B6EZQCAvGRmJidM3Wj+y+REIt4Law91M7NR2eWSY77Z9isKwE7
N6lNercgKMImsYSnQSLTyOucFKObEzURSo6icZcq37darTk56k77PnUfg2aBmn4F
adYZT0qGSlqaQEn1n683I72KVTHKXJT4zwK9M0A1seFmvWZwBVdyb33kO6nszzzw
aXWtSR0vCgbLOB1xxHzjN2/iPmXwgj8UOih/G3THC99K7hUXp/Pll7Fym6gp8xWp
fDRExDfwXY9tz/kwjhJxwCmBLcetb93ZnfPuMpNYpWLRWGRbG1GWEmx3ELUhFFRp
WLVS7xjrHLurxr51RgVEZQO+7CFyRHAU8ggaqEds4ZK50L741J00D2u+hJz8F9dH
4d5WFJ9CFS63ZBfc2SStcwkSOw+ux0IDssJejSiAEeZzLMyhlMdB0NNi+yhnDfj3
pi/wsUsPUfdz692UF9MG9hjkkd1eJ29/6veZ6/0G9+ajtVFLBE9jiFaB3hsjhNcJ
U1ekZh6yJXTg3DvAOkUKWSfzJBsIkK9KsGeozDxiL2LQlpnEiIihwIxPYIr5I/o/
iphN2/sZwhiwj2IgmHH8VLRalsHEMFQdqsQQZEAzMhQ2/II+kGLFd5o1yZxy/W3E
y7ZOhWXTqHqcTZqfSvFMqjzJ/y6IfNLwEMx1NOxI1/hsOukMFAmbqfZVRoSeLxhj
EsNszt0EpD/3fG4CcHIlLDMC6q8OrWrb/fsRnE62DuTiTu9omjumEJTOQQhGDBQP
xTEDn3KUKgm29B8ahWtAyMueAcY4R5jRgQMyGuOiUk7P+HGnRaKGPYu+mJjP4Rff
xHXYZEihCv0BkFoykfBGScZFigYuCjGWRL0MzLJxyX8KogH59jNQ0aW1IKdpTPbU
Gk58GlzR/ljWyuq3dWOU/0f3zJK/1DVbJt9OC4Ie1wtfP1qZjNYw6RehvdkN9HOC
qWVA3jPXIEYuKFo6EGq2YYzSfXEyvli4/qoXoDLje4sJtj3/oZGNlotdAXr+or4E
rGjpbpfB8xldbh2RnQ1VCvNcD8Q7u+81N60iRt9wDCofN4iQvsvengOe/DRwLpAn
dWoCUaE8GVjEszsU4kiN8Ay3KOziVWIJSNICu+PvRdXRlGpLXAhAcRZ6AcTbE1xu
bvfLw4Td0EUK5fdjN9jAPiC3PA3uCze6pWqBJlfaOL7Cc5rxdgBVZFP3FADz3AJt
Xm+TiiDMe19dod8l75p+t1oqJ/gv82E7F/QVRxTQnYhAcT/FkTkDrqTToJfj7irC
cPxlJxROQwslGWlnsFt8X3bo7gxIWORAvZCWF1TCmCoRGeDws+iKUDUdAoM3MPf1
WHGAV9zBu7h1Lp5hzl6ecpWBL8mcvAq7g3iIT1jQJHBZf3I1kTNq6LOONaBIz4CI
U/wv7ZH46UyV6G5Z6VENOV9PPjw0MP8Ww07hZAXTnMegx7dQGeM2SEiEajR8N7he
QIf2BkBCp6hCH3LXZxS0VzyLfiNnpfY0b+5YzIyIQU99Lly3NkFSOMdOnY64EpkU
XC6IePJlFuVgmgMmT0qZ5jisRFDxcMLIiJMqTioe4FBR5LrObJi9Lr/1SiIlfMKi
+awY/i9YvZeUWS1vtwr9En6MugqpOFUus8Pi1OA+ySiF6Me11zEOxKng5iRZkbyB
qPpfgR3E2zV0t8i/heuVysuiiicOw+JKHkQm4sYUoujjBVbuQ24UNDXm6AglUwp+
IOdnLsfcGRvyOv9gOBsIN+NPbPS3iFXw5Ln6tpPG4Jx69ZDFgWh89Xv9UgytJlDY
Bgv2yaXZ0n9nMoTFL/Gxr9ItjiDRqo5N+i3zUiR6zDcMpoEwXB0gtbeRjFwsOOPc
zJxEO07oeeK2uwfSoo3Px0zXuGpBAkjsHpwttlAncYWY/eHhIQKHP5nG7kA915tR
VK6ZJ33R9Bg5pN6sx3I8uWP4G6cDW+XNNQLXLEFvMWOcabUXjKGCbSSAEPojQugw
fqlzMrwOPmbucnUrFkEj2PasDL/z+V315aGG3Ss/JtCB7z21roan1L3TeDogHPre
g2c7cxTnrIInaXultOfw95GzEVRm+S0dTo6AwcseneqaMQgV3Aq+QQ1akXjmb/OB
GWKh2ZhIXeEFaGs+1e5HOK97CPZY0Pa4ZHm88n7fCtYO7uuJGA0idxcpKKFrz5QK
bd5/sIMS0bjn+ioCQIy8RSya5YANb7oJYwKteq29xOjbOjLJ4y3Z4nOJ87LGKWKg
iRcQGCeCWuJyrDWJWpvC6r7J7EloweEp8GLbR1B8TVq96+tDshohNBGs+strlsQo
DpOABKIDunfL8x/g6qt3fCwhj6UmIWeEGtrtiDWvbhxkA0eqWokTTRR5q7OBoaP/
pzyVzRNYpLP3A5v97IrvrEKI5dw9DtFPo72DCX/a/xffoq3tVW44Z2IS/OkAWg8q
8YfIZhtD61+B6EHJZjQCKficIUWY7slilIpvUI7ceHAs55fwFLb1DQ7BDg0ibQtU
MhZYnJe1/dfk8egnthbkPnxgxgGLGtGRL8fvWJMdftRfemFKic96ojE2nUNOJxif
XOfJ4vO0TyxQwVBU4MmMZ/pPJVYvz04/tb+d10rOukYaRESJb/RLUx5gxvcRtZFj
sR2uN7bhiZ5ZG1wSBgj8PJSDMH+I5XB4S+Zg7EjVV6YVWLqITLXsZ6GpGn6SG9WH
zKNbAvkJqfgO7SxN4CJnD1tCy6uH0yEUq2fH4wbrYHPTlnN4tNO/ofUBjwkNd64m
JUyJM6DONw0PLr0h3hAcbXjC4mqd/2DcZFcg7HMYQo6pPPrdlumch03oCBqtgKh2
RTwFAxWNo+rhTXoREP/gCn8CZRY15FgYWzNmJBwIvaPY2pq3si6vCE/lfZQTQ/Jb
dDQAGgWB+STaGRQiK7NSGy+a/UKyOiEShv7NpwOcPjJrm4VLiRiUuWMQtEpO+SxH
9/pbK8jIucwPzSZenZ2Ejy04qa/9uYPR9+ofUk0jGDwr3wAeauMO/MKAV/rUDTcq
Z/QqydxmLNJReDQroyindhXC4uDgh+el0rV9Ahqy6xbfgEkhuyU+3UwI/PxV4VTN
yDv5qdLbdXMAjApX8fAURitycyAeZAmHHkwYUr+GdW4bQjafK1b0yxVSDikpcbVJ
sCaNkHh2D74ovI28AFirq6u9HHwiRZfqGzNSd8YNqWXknyby5bIwb+duaWGbjnJM
8L9t9xtnBl5J+DoUQBEHiDzco8kq/Pv5MgCDdVcADvfUtxxHkJPUvrwozSwy8v0V
0FemrfAfwY5NfCmJ7tgVIqSeaUolaHOzpCKFQmOyfv4tlf5kLSAUPkCltv/0pxQ7
/OZrQHrEdcLhs9VW2p4jNpnxgB/u0Qlf+J5GtMPH6oDgc4ZYlHrVjLc5VTDKuOKC
L4CXAHVkRgjzr1iUnc1ZfkHyaksm/XcJjGtZW92xFZ3Vc4yIBaGAh89AmxE0FYXj
1ia+ExInqpKpC30vrPwqSSBL7GpgMTqWRVnXXvO4lvjoT83UvHbn5rbJM4d9PA3H
wdjjxHf8h8syzXY8js/8s+YsD1swVJ4kY9eC+t2eOnLf/MSf/VEh7Dx2zNoJ0ABZ
JD4kLSRf+39F2CjMC4/6T0ILY2nCKBReZ7/sEXZAfqyzkESmR8UwbxwF71KquNZG
d1UifbhNqJl4pt4UH1n13MCeMros2UlJHg+DyiRN8Tf0Ttm4rw3VljcBu4wsLRJs
2u3RpZYZDAWtoodK6RpxDAfTHJePV5eup25QtVpfsy4v+1HRfJNcZGMfJd3i+4v7
GjMddXERnHn6EnQqW4bAS+Yh+SWcvhNGI49RKrYIr9rHLwGI0QbNVcWNg3CU2GeR
QePKBq3dTHEZnT1+WhONUK/31R7hZNdeIzUvXcO/HxEAXOWfOKs/02D/Kb4091L4
V5M5GUkPV1gywqLEJrUgKISz+vnWhgXv+D17jMYZkVFrqKEaNHyPP4SHXpXyINyO
Rt3fU+YZUyaFvCPoLlOMOoIDxjJDSac+rQPZDLSfaCGesaJsY+l6oKj9yp8pzO6d
X/0Hu9OgG4m9BAwk76rUoZsuafoldYWWnmaZOyNKNsyxaulUgRR2TzJrpK+st8vv
uMo/PwGG8Tcc4Vp8Vg3ezWnUQQW3jFqQDePJC5jrJSiKZx5oNxD7yZHj1RTcGWjI
qG0WaX9iaaETnezHUeBHefCoFysVEyOQXIsFyH/AdxID8K9WPSvYxLsUrRcMJUwN
G/QwELw1isLW2bBsu2ikxhl0WU177YRC1eS0xPIbP921GnEPiuqdMZqwrAtxkLTI
JnvK3mRAtRXt62DgWjerT5MuTir6nyZTxYNJxfl4/qUBtqb5tTEuMcxTLtNl2jNc
tmODXuF+hW7V1jfih8FTdIJTYGMu0d1oCIDPwwJRDmdj0bhMf3/jvxekGynZu6vi
HDCgDO7Bw4YS1d/yjrd+NgIDH8ShTIBTH/8fCGShsQD/sDHQIGW4mDOLUkFvUM1k
Hblqsyb1A+sn3xp6Ge8KbrGYUDeAmod4Cr0r9U5dczUiurCIliGWu+B+AUj75Bmu
YQNXYEMOhirinTZgjH5LOebdOoSlV0Ja3/CaOasBm4I72LtPREn4zMoJXSXWsNEi
frNJ8LOaVkWKDL7FEY8JbxrHA5q0CoMLI5Eyylv3Gj/z5rK1FU+PCLLZbQ8IQK83
zuD9+gI2wYepPX6m9uAx3ZnO1aAb2xBgG9FYt8de2QvlCMO+dfIdCNo4rozuUgrU
hcTx/qr4qiVkVlnkhAXUkwHNziRsO8BXEcVCfDupZ0OomDS4nn2lLxnn7Nbg+0Em
St4LNQV7CqUG2zVojIwUGT2KpeDOWr5PRm0DJTLZXq06CHoarA4v1NHDFgQNoVgk
NNRpTdE0zlUpAGM16cxBduzM5AM9RtAr3vc7shh/O25RPu5h3VpwiXonY31/PCnT
ERvcaLP9lpnAy4vMfbxP9KfzWNPlf3GtL0iFj1HSt4Qe1oZQscJH+6LKr2LWr/s/
pks9Py3LkNtwR1Gr7gTMFDQYwxqwlgJ5n4LZECz2YqnSfHA52UBmrj5wTuwf82Am
JYVFn2LafcZifk6AAVfi/82ECBWVlLgnuQ4w8yY2/1bwWJEDOHvbfOfJ1WXgyCiH
nbw218itNKHHusOTVERvqy5PVTyKpODEECFf+3Co980AXdQNrLGxp7R489IV5HKY
4/M8J37x7Hp2DUop/3ASEbuJEtrQxuGPpZyy/wW64kkSwMEPBnPEIEGuAvFYJ1wt
CClKzM3wzgT/mgO6gBHO47HohqwVD4LDW7+C3k+MzPNK1QyM/668ZdLZqrWEkBg7
3M4/qF/zLQcNKGphOQaZfspJpmRRgHNhRSGHO7Y5vnfOdvhUka5PCY18NtLUVlA5
VpR1ifvOIa5fPgoeyRgN+clpMwTL6de1stm/oXmrijEznwX/DSY7v4DqGIljeceD
3El/slzNFPfahfYz6ZFFXzWSmyQMxrBwO6qCkRWyEadqT4aU3lEKFVA5FmH1EC8C
L55O5T9FGi47poBfN/I5HpkxVfCXA1xhF5dzBhRySsdfg/CQKA/XEIgvsDCylleW
7TOCcfPfm+M3b583EaaM/QcByZ7wbguyaWAHA0QoB8Iy5U63o8Td9J3sSeBpG2V1
DMn5jZTM+IHGK2XLVK8H2udiDeh6MkXsBia2QHnaLsq6qYHbGyZx7N6LDCL/fRO6
CG8CJBXet8/GJ0shSoTfDSnxpFtMfo6VvldLbme3EpTokQpoxDtEm7Dtyy2hB60f
6V/BO8QmZZTdq228ruWPiX+PtKU8HdvyCB68b7Z5XDDTA3seVwOQmrbqEzNjRI4k
XSfG6cd8haiw9xHtGPTEjzW8Az707J23IumOJ3D6800rBa6lGC3CItd38hvGapEW
JwPWJ44Yi7kFccJWRMdq6zue/q/lSlVV9J1yMscRmzSGC/+0Jt1PbK/sRHVCcbDf
mlkGwOlMXK5F8GKIKFrCq4Uc6IaQ2d+4la/vh9ugVLgZLNyFnCaPS/vq5sc64TU2
XKuT4fXA5aw0gWJhzEw831yfMTNRiszH7sIzXrQPec5DpF+nY6mrMqYVWYJD+BSt
mA1rZnwg0YHD8sFEd5UijBezcwd+IyGigzslQOneUNmZvk0SHUCerY+Ut0ZJCaSV
fSS4LurTJRmcc6uClD70DXnJ8rTN0vtbO7MIw2PqLhSkwbPE4p/clk6u6G5FW47f
+WTkBAkIkLVL3SUkH1Ocd81taplWqPTur5K9hIeLrYqZGjQa6lWxaER8GFHrbHdC
tiPx575sHyvdpaKzcaJYwFyxN2gdUD35jTAw4pTYBFsDXGvMWUtI1jiSj6DnBsP4
Sqb72eAL8lC2xR26OyphUxAY0zQZ/UsOaEUx8CJ6JTTVieSV3NaY1NF6LBirMLHf
XkvDyDhg2C+d7NeYyfuCj8vvvWpB31n9ILyC5TrjfwlesuAzz+uEf6cIUL/F0cXk
2pEJcVJyNCFWJ5pAcR7Ln0NAzkTLuP8oqukYjThF2lhWE7EVjy0EBH1arAFmQFhq
4MvHQaPGGv7fuNhFbmaKHKYONLaL+8O1M4naO+N73GRmkTSyU2I1epWzmM42tY+V
Nv91TEo1EcJrxg8BRRAGNnSYpAXme8szi9BLF5Jtu9r/wkdfk15xR0sniT/GoKE8
NW9zOGDjxvblGwhgBAlOzur1QPy24oUN7cvibEFzbp/bEXKfBSG/zReVfnG63BDD
nfuiT5FCAhGNfk68UftJwYnrVrKGQ2W+roiD483ST4E3tA3DwOO3fvWHRLtGp8bs
181U/glx7GCG2skSB3dIpadT2ONOxkWL9hOpB+LxaWWlJO1yOo7tHVq4UgmsLdnh
ekXHUWL9ySjecz/ID//Mu0PpxO+q3bdYlE8OeepXIpXlgDmn7IY6G3Y7jJehoHin
9Jc2NyeDpAz/0nf+t03ofzFlFqRcbLlTpefIUJS+xe1PDJRzZyJSp1STkfJsN0BU
OFF01BkaDZje1R0y7RP9sK84W7cqo9iJ902NlT+V5ukJMVdN5W5GbH37PQOHpIw0
OyNlcp6OwxdKiV61DFm3UUbid/aypprGSzGlIlRu5K1y446daHJZS5KTjQblIMQw
e8PeAugcNSDzlaCuE26q1Gxpdlmnf97MG16tfvtTCfcXUk3MBQOkup31AHvrqEE0
u5K8U0PCGAxOoQxFE5RVhMd4K+UxPPzm8mzIvP7R3/qi0A6X8wJkrqCk/1kjIxfc
KCXQtMoB0ve7u+az9WvfdYhQC8/m50PowkXnbNViIOkZT/zGNxS71VCA+XzTZmjd
ua1qg0KEeE4Bqay/iPwzbkuIwH8QyIcYTc1M35mY+PDCoT6r6aWNJBCZKUZfaejf
q61QadvtMXqWc1qAQg6dhfEmUYN3246k6oW846NEkVc2uMHNpIrRYmuv8OSK9qg/
wx8xR2Sxd/fHwrgXW2+ObEPnSfy6UIZf7f/v9OlB1s14e9On8KZomiuOBPnrQhOU
JDztdirNbRHhzy0ugPRq6FhXWYloGizY1+Sr0pgAjPUV9qzaHj83S9rANt2yCxK3
SQ05QLlHEJncqL7GXFsyEW1ldPYEOhwxFa6oFIa+ryOgFFR0Jo587HcjmH2kk6kg
/gjxn6mI7cjnw8kdtQfAerjHTArDsK4oghj+2YaId3AoRNY1zObThEaiJvN7aZF4
/+GLp2ebP1ceRcV2GuC5UT8lV5P9tqCWZw0hTnsjorCyDfjdROgiN5y6pA3iL4qg
9EAk8/lFr3P8zrqCrJtFIpDQjg3mDC0QGFW7DXInCYYM0NAVszTYFChJdCvebvPd
vWTdpSBjcDVQgjxWALAsjiNypbB+P/MQjMLsIcYL/DPGJkocMd0K1JzcmrAgE5U3
8tcWiBchu5EnNbJygSAhqbAaA8jX4xYRQssx5nCoyotyrwv1sApPCKSP0eStR+lo
3oMIehPipqztZjGN3wn342L9O1YBjoCdHUBnngn5/vLZ3nmV9I/PQSYrampvO2WP
kPy9P3BNxaimnAZj9QWGQShC2lVj9OrCqZI2pWXz/+TRK19f/rbL8ISfqDRCL9fz
7ykd6jVaxNhm8MyfdioFPaUbbF0T+2xOJaovf8OD/lzbHHGK838NTa5jHX73VOgk
RFRoXaWAM3mgszsSseV6yXTDxeZsfmGJVeMcNadDdg+yBkDLCkdjM5W2FQRBA22x
LBtLara1ko7YlomEbi7TT2xolzMjjQaBI0qGvstDrsrLkq7VSPvvJUuXohI2wpD2
fYRDuZ4/8VTnzva9ln9K4DGq7R60Z913KIZQ6B0c0EC5x9WNkzuTe49RZaZ8hINE
ncoMRa/UIHHIEt6kSZi62yQn2eDrT29jPjLU2hxNdYAHrcm/umtl04KEa8AxEV+4
UkBRLvVcwzj+HuCDKR+4UIIkMpsNnDT1ZsqMq8yoocbYFCYwm/v+fMAE+IiOi7sy
iU/1GVvjWp6yvR12oCdC5v+F8sJrPOXrwDjMQx+0pjbVNjoCho94P4RrGg/ptISk
XWwwu6RprulZh2LcHvywdiFt/N7KvWwg03ULLoaKl/YKnO5GCia2aILOERTLOxH7
06YQGM4IFqNIFa+KYiMLF/0ok0cBZ1aLMVqTtzYfcNPsvZyqCkczjaJjZANLb3xU
3Jn3qBSIFLplBPI8dZe/cMP7C4Hs7oc3uOOBet+JrzQ4a9sJKunjKoJ5zG4fQ8N7
kM4MqKqJQsNbel6WH9p/3oVBRXfQLhAcQeH9PclpxRWEcQVh1bPMsZSd+11al9da
pKkPCZMKU5gacgqiIG2cZ64o5EB3ekxKIm5cU9dT3hTAho3jFLDguop9DPxe+UmG
HXCxOT15TlRMeO5GWF/TsCPRa8/MfOJm9T506XLP7vvpYrL95k7Ucrpdevo2mzR0
bmzj/yL1hRIOizdssFe25SDYxlP0UO2yh3HqjgUEMFh0XkKKq/GWf8qhVINOuJj4
ECg/+S95ebmeEaxSYzpt1bYYPSvjlBgxngcVbBfmROBBnfOq2/tqw8yrM1u/2VMu
Beto/h49LB9fkA/AniTA77LAXEPt0m286jSzkxeTjGOVHHhywoGbpsQuwTm4IiUU
KTPDPYVvbewo58PcXVP7b1VtuaxqFdM0ks1/69/bvmMu/ZcZ8E88rz584uJ0+zty
ONRF5TWi6t73TjcOShO7uMRmWW251T9sxDiXztaWhz+fQJk283JhvuD+GbfYl6lF
2HRdRjiyuT7nIQ2a2Em1oJwN9+y65pmxFZLpWx6iiivGDws82jOKv2fAbX9rU1ht
V9nSQxmdsT0GBx2Rlgwm0bjRA4jOceZRLOGggUUfelbwvoo8AS72YI1ajlVkQBX5
+cMHfLTrjqh+FWcTxUs45SUmrIFhAHFlCCN2skl5Qd/4acWXoiv3CP4ZloqQadaj
gTqGtsrY8DeWB9vjxC15jwQSWc2pk5tc0YeHAgO1dmHCmapLZSNUyHFZ7CyCNOHV
kqaa7ZVqZt3dHovceG9maA0GBql8Q1BbVJ5AGLiJk9+8EcwdCgqYAZyBif8q7ieh
sbmcByQ3rGEpB7C6DiSKB+zlgfzDgY6R16fCsrkg87jhcnhOJKzqsPKRy5CxdCng
UbWHOh/P4GaJayQ1mnUcQJ/m/mQB3Q73pidUwI/meC3G2VL8i9+wuMj+qsb0Q8dw
7Rgxzib9CthCROmkT6xt4LYu2dJvM5dulP5M1U768Bs3gyWwBs9G2qCCH+u1XR/O
8Z1Jt+RoryIGIW+lYJKX9L7y8Wtorqs+claS+9rV+oZZY2nou7ZcrEd5RSWIiXux
juKVTFh/IhQZA1l6pkPJS7GbXZPbLXPHS/llSRLDqWCfwYZXLDNyY2ZH0xNYimzJ
Ks+XMacXgwMwU4SePz5IPZwQLbPwaa2TUgpABoPNppL2PCUxj/7/8IC9idWKre9y
yYCaaIDTQjvMvnAMRjNHDdOwNjzPgCAzS6FzeNf5vUc5n1sSk0do+C/UnjJyzQjQ
gMqmshSGh1OjIAWKVPJaR0Esd7Yp2QYuv/iGiNQL3oGB8REP5pQl6TXrjbY7rzDb
d4UIl9cS1xCx9bWeMrkN0b4/b4e51e5sfW6/agXcEPzbUg9P9DZxUMiL1c+qNsFd
cPfSDkCteNlKSXRzxryNyiNFXV/WQpvLJTas1eql4zn3BZrpmvkEOWI3WXietqY1
isfY8EkYrx2NQsvHlIJ2YEPDqmZqWoId7NT48Nq34K/tIj2bw/0WuKH4kKBIlWeR
2bKDP0oBRB0aReZSNuB/2CyOaCJN+aJRKzCqs9qOdduOCSFCr/JbmGrbRfMLBugV
WufMK0FFvJ0402alrgcPjyCxYjeoHhfsTFbPbV2UeSpYhVPL0BMTXQItNN8rBORs
Qymvm/G2ZUPDEFQc2J3ih+QdyVxwzel6gIvq9Rm6RSedgH9JwIjp1mEVuNQSFmnO
HGdFfmGzhQTj/by4WdC6tOLD/yKmE1ECkHcOryQzdd/JC1M8Ul2qJo23Hpaibu/N
32cXUIKZE+Hki1vUyLfuUFhnTCqr88i/ec3MNoA/Kdb1SCD5iKogsLC5FvILU04+
KnAEjbbgf7zRM9oZeQQrltuEQgm84l1bp5YLF3/t3Q7G/EgpvtIoF9+X1R+MqOe3
UwAU8jVk7ZF5UM1DSU/ZLrSvPXSiXKaKLmIZC5GUuHMhFFnNRxFjH1qDklzQSTQD
bZZZE8KK1VCdT4JpB13Ndd+FAadexeuDvENw9vyQ1wH8knI5DJY1tdg+cm7F6fyK
pPkJrePQYETpwtLmN9BQPb1XuRpcp6h4Gr3m7fNq9/rLheFr/DrDpj2Zsrte54I6
Qt51gzJu2OgzllK6g/dmDHZR4H901GTvA6QmNvG+TQ4L+fBj+QTBjMJIA11cH549
vSWFxuPoGZajxZ74EoShm/FJZZtUNvg5WvuIocyxsjhtQNqdXdjWUpizNf1No9Ur
cQgPOXdLpPXNy9g3vLbvqNFZJBE5OZikS1U1jbEnkvO6rjTuKx1jjGEhfscu41+q
pL8Lfm0dZWwhMglS7Ospui5H2RsD96fswEUL6t0v3Lh5YpVDqFnq6tfO8dl42PuD
I+HLAYSOHXM6+FFCggZjTk9LQjumG2e+R4YBShC9u9eFFGco3d8Sp737mb0LKsO4
zU6FJh3Da7IULcCvb6FThx3Pqshf2PtZ0uOsdfK4XQOj6+6wSPSj8C8g5gPYfXQy
TvNoKRmGkgFuhgQHtBLhxBOZjAYd7kw2ZvKyfsybq6/7WKkBN7LzampbeEYw4bxJ
v9FaU5tZa+sNO3vDY+FaW3NhCeYhYHYQClm3fi6K9UZqtyJPGoUoyvk7qq+94ItP
p1uBQOPN2szN5agBWyEoXAN3o/3wZz3WbPPLUibmjJDJ5YWkgDQVlv9m4pOjVLAU
QPTRN+5hZIxSW4uiGXybGt1G9mLo+ZawG4x4jt0iVN9MxEL362I0/+l+zg6m6nOd
Q1UeS24ywV0yl3JBjVZBwWm1bdGYT9kldrbPQH0G1fAj+jlMxFVlRuGAxjO6G97J
DCWeIiWdnLVq0N5hsrV1lt/MHkcpHqRGH9DTUS5q+Q5vLeXSgiKY50Tw+/sV3haW
leQHOXYvtO2NWRaszN/LAvoYbguurkl6YPcnQrnpaV3srN+DXaj2b+tELyC1u8MS
VFmznqolurC2wH3w6FoxVO0Z0uPg4Ym8zzU3Aa+HQ2onsSpcO4TJecjy5dcxsYSS
ArMW/RKLfG8Iega+N5Ua4YrFSmiR4a6BxEypxjWtwtP2a2PESEGm5C2hx5nT2c8f
YJpYPBJdBuevjBVfqUzoERGKrzHnAycK7WrjNebemj4KypIMxqSApuLMvc8DKYq6
xxiVeHcga+dTUuC0AtFzIIl8ci7wdcxmZ9QmMqCLTKuyaL9WaSCPPYJCzajudzlB
3FN5BjFT+VDObVtBOmAPI9IoM4OMWDF/t4uGtomaJlFqmpBnwklNR17yUCjJcOKV
FBlkIAfh9jBKx+ZHEKOOnwK8SzY134YqLqkKtCLqdjz8xx2oM0WRXEUrJ6OFoUdH
ok3b2YQPjQV1GyKMLApHOkE7iTMrZ9LSU8RYtvop/oKaBlcpPBhMTJWnrOJsufMd
wbcB29FF+rBI+quCeKOrFsmJdVNcqAR8OeSU95pfr+LyTb+X6sUKaaTumRyd9as4
LWlW/htoR3K2nbTrkiPo8K2JoIIPxIcmEiwwYYo/N/XinAZMj9cg8Xff2QjtE3dQ
wcjmv4WOWCLiby76mN3rtUsVPLzhwpw9mijokNh0W8al9qYx/YHIQOJb58ymyQdC
SVhw5QUxomWInIwTS0gIp2x4C+yr1jO14MQtMU0HQ7ejQ+5Pk/hB8ZgeDtivbRGu
mGwNg0LnS/PVVM+wQGG5ZCQr2k9/VJfYQogg4MzvKRQTP1dMkCDW0BjhWWfWpf1O
TaRzqfbBOyt0ehs2oA61+1FqK4YZmjhvnDPJ/64kFO5PhJ3bWzT70NABVhk8H2hp
VrDzWWqLgW9NbtAt3AHI/JFJZPKBEQXr3b+xmccT+QOlL7pUzayKyCKByqjPl+EK
FUNiHkDmEcTVkf5qvJmHQ3mcEodxefZ1CsphRISEB/OMz3513dwgJ2l/iEDnR+w8
zCRCIVhtJ0pCDiFDuo/61lGWiHL0OI1yMpzQ5DR1NGRFcdSEjD0oO4PlvHrKZZGi
Idlz933shFY4asxVjJ0AVbfHxgkSuBh1G/n0nu08LZFeK3bypynkLZWOTfI+Htr6
evm5GxNnxHT2tAQ63pVgNsUXjwQv4t9sPFH6IBSboLUWQ0+vjVagRuJ+LWLj3n4J
VHWwSgKl/uxSai0x8wcA+s2it9cXC1MR47iLJeadMDuKwsYGssD+O/aEcmT3UM33
cgAin8GKQSu6+sQGhTjwsULPbuRnf9Ugij0xqzS9ZDZ4lm0iI4hdZezFCTrYd9vk
dyL8TcBCGU9m97FaNw7cSIKAOq68ysXxHRsogByZsO3gmUXaMLVZWLYzSdYLLPG0
JSLZExWX4zngniWRDC1Z5QASDL6VDAEe3hJ3H94IkTsYPDm2Aso3Ode88hO+kVxJ
xko8ktbR5jACQEXf5nefqX9hWS63oShwUYxnXQB9QZHbEx167Pwkb6zzg6Fzujqk
A8Sfnzm+HgwY4aEGHn+Pp3i8pfF4bBLQxdCaJvtBUz6HqbJ76bQ62x6iQr1zaGI0
aFJJ/reLmdtN6qiIQJsbi+AkTF1NOZio4pqwvzM8RGfXGZfE2ZxN/Jojmwjyv+vk
4fPuQXptvnvJQ6mO62aBiPorVBh9Lw7czQ5gyyiS6YsE7nSgQd4yJbs1UW9p+xVf
E7NYUmObWdXF4wyFAdDXydH2XWXYE/uT0gy9yKI3IsccT45sZpLbLbcrLRCCjlEi
grhXS8/pc0usBTsKqQQ0EuUwy3UGLO2z4DZAo0xDwQlEVMXXwKwc9SJoJTO2iGZt
SmHGI3Z9Igw72iCl87PvRD9PfBrb/SpSmB5ZMVyapZYbDklq6h1HE+h8lOP2n8Xj
uhD4VYsdLpbN0bIQJMMa+sUjzwsorO/LvccBcIlFzXSmPvi3Q55fuBcvjW3QLC+z
/FQJMpk6VgC4w4NoWufOyG9dl2EoG3zDi5q8/TTS7wi/WJqUJIUYRr8NSvnF/JEP
EMcqxVSGwXoqSTZsIshguA9M7O0SlOMVCwR4auaJN2OtFCg3qIPfa414ozJKddDT
LEynoqzb380BDuIFXD2S5Cn7ktR160z/gTe5HfVHzQAKt97nlRQyH1DXs3S5FuCW
BZTyLjN+CigmkpU3vbiJsSkZBM3aRBGNnSmWbOn6Or9QkY8Xpc+9duk7TRCWf79X
l77WQGZ2UBfE83bVXgBZNX4BTiKxPW3LDwej1TnLgRI+NrT0VxT8pLRzDmLySFx9
SDz2TS9KpAWsyGQG+s0c6eBdIFd31cvoPwWDYFikb4p2lp51WXNlWDW2qc4fxMgq
wKvTb4fk3aSDsOvxzOl3G7/rbQu7TKLUbaza1q0fSE97TNpugmBmf9JkpNXRT3pq
SSPdLyVpD89kniuzRA6GboxtMgwFI4GRPMH+FoEooUMH2e4f2uQitpNc5K+dAwxC
kIjj0pzt3WvwP4EkAUyrzldYvmXHh4iOd6Wg5BOyKtsho+UR3/e/zOoD00PrBAId
8shaqr89oSdZcoEmN2hVdmy6T95QlnlqcVYsMQ6bNRGfaB7MQQeykeA+RfbcJpaJ
a+C8id6QX9yiOKxKc6c80ZrUHUENTnfoDaYqsHeIostgn9iiwXxnRJ0UHR4ocIdA
k4epdrt+lBMd4OzWrFo/9iuoa4C95nHkhdWYhtZXno8K1AiqVRO2Al3SOi0zW+aC
Z09TZxwLaMXI1+V7QeTHHo7ShIVjYAa3ABoZhGFHdx3nlSs4tRJcXr9b70f8LwZx
R4EZH/M9ULIiZmV0Uu9WlbAETJaHZLbW/beNBP9iD73yzBlLXRzPCjVTYebTFwit
DacsIzip6IzMJBQEGY6HgHFhkaTvkz5wpNkKWX215Et0wOa3yGHX2MjRwfR72Fh1
ygTNVy3A7oRC4t8lEVdCJXb6LbfHl1CHg65vxcqFeTwJsXtQSk7e7ai30EYf9icy
mo1xdhyy1im/l0M8zfYW1iZDL7/ZEk4FmebrU7EYxbOrlgcE1GmrVuDtocIAdpT/
P6VCGG0L3sZIG5Htdf2Fztjyu3S1zY10RCU9S1Qm8DzFykg7fTx0AF2XdY8XNcOh
AaQiVNi6vAbouFOiG+odKOHX5jMBlMAD5dY1qiH7i8JXnktvcxyBTkSRjwNzIuYx
2rOVadEs6+ddOa4PaJO/l+DRqQY5c8arRTheAc3oY0vKVjFufnTFgafxmsbuevi7
EHoWOySPud1U7mJoWMLrVvUrv0UX+UWluSmCPQt+8oM7CN2L+Uu7n9EFUYUuDsk+
wyzJ5YBnuq6EHWaBHrOlhg9R9KQ+lriABmHiQ7l0WpVSul5zPLZBTd5Yi2qKBGV5
6Wbz4V6b70L/dch9DbDzQvW07PFMXYDtI3UmxeEZQ+4sgUNehLOADFIR6mCuTbax
NL9tXbxik9Vh89hxDA0/uT2huDCLR0mYWTLZXx5SYuuTg6xUG9GgIunFQ7wH4JTh
nR2OG03KJh2YSwjZFSHDA0ml+vKds2cGpxjyh0VYpt3WNyseYX1Il/2MSejSLfHm
HdoKdCrE/7Ufc5vM/XbeNWc/8eSY1lLWUPnlQLKCa4zdJ8r2zIk2Hv/L3ctOuPx3
LlFIWsF5bhOuTays2m08mT155VxDNyl5ihpwzV7xtgUP4q1EscyQbQqDXoQ0fAqu
U/f4vpKzPhMGHCrwlalOBZKR30HFWvSTIuz2vaX106dP6durk96tzMO+iRy0CrAp
lZ8xbi3HIMdwnk9GNLmQ/3Pzz1zR0Kemr6lme2mGTyAR9zD4DUl+DKWOzpvzm3gn
JznaD5R44Ei2UmACVr/bk1EcxwxizxJGpjWXy2QF7kLmyP/fEFT56DauMcrl1oSs
ZUQ06veQoIhrvGz7TCHIX/w9dbwxJ+UlRWLJHE4JwMf2wnWD1EZlGnQaSNnmGrcI
FHb+20IvZRzAG1GyFqh9BCfeh/rktnqs94jJUWv97098HAkIONOseh/55V6+J/gh
RESyRuHjkEMFl2fGTy+rA5yZKI6mtbBh2QTOjIqlcTmaqcIp7FzxPTB4StN+7yoI
ZmHAZnj3WcK2tTJnvAOGPENMK+Bvs+DkpLU9TMIXva6IaatKWbdxH3/zfQ14Q1ba
+VkDBmgJtv8oljWdjPOaMjX1A7UPz+KU5FOKVZRPvkdSwrC8h9P3kJEOoXTRVRXs
g5fg/c9AZ8/SgX8WH6RD2N5uv/Z0QpsxTkb3LC3l8IvfDt+x0qvVrHr6/wLApDQ9
RJ3KjeRNSmpuCWP7kE3vYFBL+7P9yiL10Y4u6QFM53ni7CzKabgXdSztzhGeqNi7
755fx05MFqeaIFKIeo99VQCGJvtFXQpuFbYSpF38SjJjfDzL85iCm30zetgbKPDM
bOVSYJmeYiCBL8Mm9rbYMnvx3nKX8fatFXuIt3jLmanBgsUC2dFQ7mrAN6sVB9Ed
13Yt4Y5WT5oSavcxY6WkxRmoBymI0OrmsbAs9aq/AZQBh5M0NOX+KuNp266Ld/We
w5hPLlYLeDpEupYdA0V0JXtbA88oOJgW3oO4ZAzDQLj3ejpWOMG1dum4W9MgURTA
nR6OV8Y2Xo6X1ddILqEvmb7rcIxtahBvO5V+TjWosPL64GFFqHOnQffYolEaw7g6
FclM7lrWKa+lFlpfD15LYaqrS52riLIjOAxs95ycdPaiVQMC2Z+OYQLmiBzAbh5g
ITDCrWbe/tjLT9RTmfsNG9m9/4tc5LvrEnSnYkSJHgISOagdtQijDMoiTFuVR8Ho
MReCGmsSrbh712F39fSPDu5rTjTsHQCRgx5ePKVOI/s1LntzFKK7/WtcqeW7n3gQ
/cK/7HrQv+dGochFKUD7LnL0YFqTZzjiFPyB55e8HbInqurRanS7Q+FMb0cRF1cw
n4sHCnTJlsX8QcYefvgBbnSjBf2u33CqfSPh50gW9RJ1aIrYrgRlOblmMPbqDFIB
U+xesgEYezLyNKbIMapqp2DJZvJzY/EgAOpzUZ6xS8hmxOR5zarD/8lMhshOgoec
CP6ZGGgbEnwxOphrxl5DZmTXqIAWFvdIwTVBb8CksSccB86UZUAazYNGNON4Jfwe
o2O53SRJknhVqVPIoL8dFqgQhrCkZxBIK6paXTFv6eVhekZ5H6o+rOJmRGjxZ7N8
DPB4pGPRT9dXUo7Si4u6Htq9rq3rhmyfiMSg7Ll8q/Ftsxa3RgHDt4ptje43G2P1
MRDwuAvSNo9iSUShlxMytzf82kT1WwXA1fsaQsIY5oYCJoFV5sJWdeQ4Hhf6lMi7
P9NvE1HrfCPOCfUVW0jPvXv2LpWtEwFJoA+h6ZO8EHc1B6fnrC2XLkDLOQIuPQ9F
rbaZV6LYfgdMu3C6MegFS2+tQhp42xSccW0gH7UsGr6EvRIDVh1jclDVohjla8Y2
HgEthL5UiD5UA7mrgUH+ch/NPvStge1AENcbncm0XKFaaWuv0iE2rxFbOi/D0D1r
p8fhihzm22u4m3vTQRNnNr2l4Zv3RHBsLcynLX5Yg8L9DMbT9EluqAfCQ87B2K66
NYYEvgsfBBcHOWe8kui9VOxBwxUjbhH5Zvev8Z9luHEYuX2kCnW19KBz5dBZ69iA
CKAJcFUbrK3h4hxxR8v1VfN40EKj1fR+QhSaA9KaNXSOFM+Lz2yS9rm2+fZzA0cn
y0qGz4ASV1SajgCvGQ5m5rodFgINvdFfJhOP0xdTYofpcbV9mACcLVyG/ueEVgz6
wHUjqyQt9wSpidgpm016AKDz0lyirmsFSqIwiIfVc6C2EPOc4lg/emU2y1yGcMQi
l5v4gHQbKiUQBtptua7bAFy2rdOLh2K9B4o95Ky/r6vRHitlaivxbGdXkOxSGsKm
2j+nlHQ9OxVzvNXF9c2Qyqsn8kyiIfHno7bQzc7ippxMCZPK+hVlMMyvtpMUttv8
uNQOpxRr9Q45/iZOR8XxvkRvtPELnw7BYrL6jON8qlM1u3NR55FPnvTuA/JeCGy8
5ARzmGJosbhJBXPukAfTo7NZd/0/ysS/Pq05SJQXLYbOWY/X23tW8qbqS5NjjNgD
z31doikXDCRlLXn6+RwhWeUI/oOtvpEyxPMh7+eII4tFo4B9kMAhJ1ZzCwHAWJdX
j0EIxoHPIxmBVRLlhNhoEm//T8CWOScLarR5rYaVBbgUqfDA/ybVKhkRqUWQDmzx
HXICJLSCOA5wS1qmr0xKkvzPXk7W4aV0stvQsg88yjdSJM4UvFM5zGLGnmNpwPx0
/yUCBK4DFW3r48rVtsULK6Hxo6zCmKmsMamepmbcZSv2WPJqDAmSD2YMWh6F+I3Q
dUTzGomo1w1IgE+vXjFEPaohtz6JZuGm0cpXhYJe99ZIvhtxNJQ6uHgFXzaG/0n7
lvLrnX8mC4umIqnj+wG7wm5Okbummhcp7eyTPLpAS/N9voVRclciEz5qdJNnLDp3
JRJEZt81PYk/jIG5pnK0X8Vr7qLU3VMhnb0CYHhxhvGkdoZiyLtlHi4DYLhgwSWR
VSyZrxCNTZPoVLLK4pj0qEwSQL+DQGrYDAoMyvJOtU447mmlkOxQCmKix3WkMMAg
DgUahb0V3Qo11PGzI4291aFN0Rdo/Gt6f8XBnDTbRerCN6nu3zoOAwWmWJbNGTbX
kZIR0LUzIY78MiS0Zg/r0BUTrSKUrDOMCnNiRFJA/jmzhpOFpoprcMrMHxmEDaJU
fm+JkGkBcDB8aum/bwXWXfytZGVKjRtLZrA2CPYNrk0SKsQTBT4D/yNcnFAEtaAt
C/J33kG13sqVEs2axxRXqTqI9CCIxxN5HEmf+DM0IQKNFEKRMwr0bWYljcIrdkRG
qU3gnnmmhzdeg8iJnKu14auR1ENMYcpL7pRuxCg9ecAz76RmX4WkgvySN+OSJVwN
g+a8l98IiCDr3qAuYwtGsBdltyL9RChLVqUUSWCqwJ50wrJ7eioFhHIpIZaztrSG
gW3ksukJ86weH9nr3bfWMOgK+0JHHYgB6S7UBL5sDqEeNj/3ivJU++C7+gL65ano
uITgFrjN0PbpuTEP7dMOxvXFQdDt0eY1Q4i9ka3f8dbZe+uf2+FfcNPXATk3AEE6
FntVl1mwp5uViqhzlNZzUJ2fnsriEr07f5YwB1TLcdQipnSd+4AnfZgjsm8VqJcd
7um+AVcYAg+mcPwqdg7PXY74vA8aZSBfQSz6Qf25IzPqTTp50Y3/Y8mkrWuFwSvU
XvpqWFeG6abvRz3/5bKSbvlOATZvdWC91XReMjcCFzoqlzwN780xhfXv+DxOmYeM
VEOY4ekveONdLLXYFTRurAqrVpoOrpmq6++xsimEoOhJ8WxMTmm/DXPoH+dvpROJ
8fNHmRLprwIMHZjyNqOLPycNxXcP89K4Ib72S0vspi1YlyJw+6xXVM55aBBQjD3p
HTcV2YjNAi5SywBuJLymD+FotCpCQRLjVy38QLhterYMJT2866HrOkpCJAhlPaeZ
Auxiy98aFYc2LkM+jieFe5OzfCX49C/K731NPhS6D54sfwr5kCjXGxS07w/XTn99
YMfvCAtkv2GFwcDgTfufAKdZuIy3Bme93iTH8nhlFJVXak7a/xkzNZ8J8yJcYOOD
KNR//YMla/5tjEYn7cRCxvBhSnhncOTT/tuUBMwy+gkY7FVcP296Dw0iMsbYlQq9
jgn7R302CtOTZRBubOLJbwDIfhekv+gKTfdyMQuPI7y+AzOUFjJOTNzyXWs74Ned
N7PVbO6ej2y941y/TblQuEG4rTn2sdggUJmMqOE/wZmaXPpCUVKfPyJ0XEZAXYw/
AwKtxqqruLeHqxEU8FZDI7OWIkO2ueG7bPrKq9wxBPi40V3fY1sZMmn5NK69g+7D
ldNrE/B3BU2ZOpL5ElizGXHAAqaaN5hyE+puTtz3f1utpecQ4tv6d54RKPd2X59N
rUHsNBREBL+S0z6cZJIQYVbD3cuSOrewuFZJRym7iJrfA49gHqWe7NIkFNJeJQWh
GV4rZsydqij7qSpvVil6LsZYFUSR7n57lp1y94ScCczKvN5VHhLdDRrolVCxILdK
SBbHVmYLxho6sJvPmFR7EFpcB4/6Bo9tGQEERvtpwnl8fvRFF+xII1FIhFKNcaCu
e1I5PNFlEc/wNg/yJhSZeZUPlUSSPsqk5CHE9HX/U4YJ+DXMAooAYnhnNV4EMXlF
vT26gH1zebf7nLFJiDGi0yBGY2dljz8xFpJS8s+citgg2WaFloMlR4pgDz2EXiVS
AL7MOvgv0AD1tfIP57V5YWe6vfMYW5GC+l6U0hcp3ZC76J1I0Z6aYVI+NzdcaYNk
jSeSnF5r28w66brpyRkbsYjr3qdDZTcN5oL83OITPJrJJTaVGvG5dhXbdgEwbGTb
GNP4HOqdGHVUTcTSkHpmQoS9s3Q+5HR/w/Z4tAkcbzPsHg78egbWTI8q0uip8IbI
T81cIdoEwsb5tKE5CTKM/7zwr+Sn+/i02tWiHjRoEK2FridkCDGGm1kkINY9m5OR
WZghnRYFclqkgniuVWcnC7yXuNw6rEtRK/A60WKNl9tcvXomLUG141QzbI0xK4Jj
a1qVR4BMMdKWocuyo02sDhM6fTpJqaD4lzrZPkA8n+Vm9Gl4ltao86ssyjTbXNhu
bFMFDsG8LKEV/DNpHKRjNWZLkCDkZ3eGcIyb//hXkDXLFfEFeDHDSl6Rr5NYiYBv
Hq4PKoN6pO46sOVHt8coUZ4JA7KZwTLCOg9XuJ/2QBaGsaPaPIrOcCVW4s22bLCu
dIy9yi5CI4kcB1v38LTmqgpf8ymOwfWSc/zxui6LoJs0aYbUwQtmb/Jk7X0iV6Jl
dtvc876nQTo5dW4FqaCo+aTVhXukI6tDuidOjOmxgXb8oMM/nXrjpqwqMxrguKzs
8c6bfL6V2J2ZQtfSug3cApCN6A5eHSmJtex8+jzDgDSceXZN6McF5TGl7Q9PGBor
ESg3GQBDwtAkzscnkm6hbWqAvo6XXYOHKi8VjD+KoN4MTlqVxHNsS8nYsId1RpvJ
8oNfzq97d1LVVzr0o17ccoi1m57e5cDMPo4NOPwvfLZF3NK0ysGaZxqX8DiOOf6R
WUm+Lyh6XFc8KmMGoTGSjzcw4a6UETVfC+JJME2z59HyKdYLSsRPYPPLHdpVczJ3
ecWJ33aMnnwUgHVLBGdX+sgiq9uO/QtENhVE5zGi4YBXLQoHtNcQ6ri84e4zw3aE
Wr4IWFNYeSd7RCzzY53pdyKVsCbwNJo+/Pk1Pq0lxJzsnBL5v9OpRc9s+zLjWaHG
RW5XB+4kY/B1XekQvpxwcpQsrumgtZ3M2Zyf8wOAIqCYI8pBeYo8lXupetVNhE4T
BP8l361xTOTHep2RPnXIGnnUSriLREEihVvMgkzQ7tb2z0K95J8CM3ar0QooSRsN
tmOqYjgWCKvN6EydyFyXzqk/Y0AfzyVP4gpaErvbm/d1LeVCaf2AGMjaEnrlJDlu
46eQ62wgGdAink0+UAUcVIb3x7KMPA3egmLvfW9l5up1wkr+X0wssvHHJbowHw25
7kF+o8iUTDEUXAOCoz7cIvAfF0PF5bCm0f6ztlb/2Rct4zhyS8KkyW5hDWTclKx4
opThNvhKDS3aNwghHTqJWGmYtA9ykGPNyc/TNPPR0YLeoWpRxEb2ZsHj+Kf+sfMd
KFWHprA2zUWdwhQlGHJ5ZG+ApWFmttbqzp3+3PnDMl2vKoqPsoohN8R4DzQ6tnXN
1TmxnFI4dJB60K1mBlCLDvayeJIC91kuuXVH+8WFtrMfgw9pChlacmSLY6uW9tmY
73Biwp5MmwRibjbRb0TRH+hnCn9HKiY71o3JXIiGVCGRnnUIwh+ZLtfyO3BbbMwb
XTzd/ubIof8J+MV6TeAgjT5F9ataWnUeZ8XvlVKJjGb0RjKVEsCkxju35JuydQGp
TOID5WAY6SOAXsMrIeWjIjf2zeoYY8FPsxw/0NdYzzLDaKlrvfbRXbwNoCnpCOAA
DjmXXSDHOJmX9Owmt4yzj5GyEsgvk8NTAgpnn+MBgRPpyK09jOuBdqESOmS2+hJs
fPB9uBytnMCoDProSfFB4ZMXLRUfzRyJcFUtm0xH19R2n0+uvI4BoRpbKo6ylQoM
T/NTSSQ1DmD7DeuGl1m0RVBoxU1Nrg5/ssCxDH+ZiSZJ9THO/72jqNZ/bbyMidNx
cfXFxs05XmFVV7nwFDVce117bUGRbq9cifiZSILxnYRuxLesFtinxnJti6zTOx8o
XJRzSN5Z54Nx+/GEnHLK7+FXOhcp4HRgcx1WLX9Cs9Q15uYhIn1ENPtibGyl2TIm
nz6ESTORNHpGl0G0/bZQtcAuLh0/jL+N0bCPjaA6EcF77p8e3E2eYZkB6CD8H9NB
u+VLo8qbH119Ki+0RSoaqZ1cicgxCGgDJnROsieIDhrC95dxa7w399m1c2XUzpxH
HXp0o/9nfkOf+0bO7NnrHVP8qHSqNJF6L0Lrg7rmxLzqauOmWm+u30Gn9XrW+4Sz
SDpko3Vc1YEz65plfKJ2jITPNfsllIad2XC/h2a0w3jtgZHaxFBC3pOuwacsFuTk
c4pMGc50WJtaSik4vSpISCvVWdp9NTLCgBG7I/+Us1IpfiBMLRQ+DfOWkjnSp9I8
L6p5EAZZQnBPt1nObkuRJFfAj4u5tsfTIbLqYAkgXhCzbYISrC7RsKGjFv3IYlFH
X+P2a3HjpiRBt50yOlWI2By/FryMsdZrUvD+noBQxnHwk9/u0y7MpRs1UpHVi3jG
+T8xCz65bw1NnWiabpdgUdl1Ih8fGp3KsgJfk0HiNMNpacm387kYIhLMoC7FM/0B
g+C1UabtuyHd9jg6MCBxz27av7FofmXv+BaDav6m9qnyOEus/56FdwZ0MLkuHbOM
PjjNAparNezXVCLDP+ccTyunwtCmZW0S79dhRDNUY7YXPclJ6o/ZKs21JYVkJ2Su
Y3B75le+f1Ty5xeOzdtgH6lcjvoZJ+mOZkqMdgL+7x1vu05vtom1x4Z0GfVxEH0L
fFmoRCFatnThlVKLKt9/ViMvJAEAgLW0oEpx0WoOZIBel5xn43bBt3xfOAx5pw/g
ru4pwW+qaYGbWLU4KrxgYV8WmsFqJSvk8GKR4EUF1MIUl+OCBDXadvAoR/fw8VXD
4NysloQYA/EJtT5ePINrynAGXoK6CG0CtQfvqH0DFCmvaE3TKJnYSMdtb0mFRHgS
mngmgWOys7+lRyXFJxe2rRzKgQY97362AKjkYWY+KSoN9lu6WfOsNl9gy+G1pD2L
vuxDsJHbLr2DULkDz30q1CV6C+YQnkmI/DP/7/RkHOO33PwuQXQ3k4bcuFAE1lSa
wXCOHnsO9sHenLIlUB683ilo1w0yk0TFgDaQjPRv1FGW80lQAy4k05xRCy6xZRde
dha3HLLv4qBaPrVrd5ziLHUT7GY0/1SpcoP8SEg1dfAdes9NGH5ac9CxQVONI5CI
XPCaaKxMvsllAQU0JDdlk8edmtf2qCj+FFWNPpexAbcFTPXkDImc9a3xB3HlVJ0I
9U9BKGlJVv8OmhjBdZLJAkTUzsEpYYAprRUNVm5VSdgGbUC9VQjl7tfVaMZvuibI
VPe4bRT78pXKR+GYdRL8wNytWsMpUqSMXY+wmsN0pEgSDeASgUSleTJBw2wzb5Z+
pIUdzk+S4s0kEb35AEgJ9rJUVxja/O972ztA4WpZzoChj+MKs00/2PkVOZDiPHD3
9yIMEOYcRW8AUHMzemMuWYazs9+9UxPI3quwg5HaJYWvYdMNcrUA3S0LBuiUmkvf
+33yddmc+BQ58dzna8m1hakN16BFE1/hrINWZSuo5S40nBfm63GTnFHPqJyKcNet
LCZ2SBuYw1/fuelrBzO4vwMK13w2MNEWCJrz8Z92Et1cOOEHhHRtiFADEOaAOD7V
fe25phbbwqWxHu2ep9HqVFphcihkCiT9kpfkPUywiAAjvcLfIX88biLXlZkF185s
C9+PSl/iPdSixRckSniYFHUgKMyZBzJA48PFBN0PoiOwWqt0F8vidFNzzQYfjfqR
Y5PU6TYqpqz5tQrAFk9r8cLXZUZviXTkiu3au6QxMjdCaD7XCjWJkAQsqaLcyIcA
QGsz84SrwWGRrkICyxG+f1y0JjQ4uHtczFOVrvBgzf2jDozkSlz+OgRNfkcZdE5u
AHrvy5FFiIHSiIi1K6a+uS9j1OcoezbKKIBzIQfwQEEiHBRMf68TVzzYPoK8O2c9
iZhRaDwfsUdP8P3Kr0M/y7u5PhoyD0l1nU79yMNZpFv1KgnNsoR53jILhGiDd0/p
hwH5XQ6OAc20O+HcaKchq/cmqRZHLLU+OzhE+4jryJAu2y2r5xmLR2b8FISH/zKF
6BPGHlXk8XGUMfvAWulay74ae+F90vDbE7PRPORpBj6bkfBQZ4OJWqbWmcNbu7UI
NvchxFFZKaoeIx6UFTXkNpRSztXbihSBC0wqDK4FFmp8PJI6RFpNJCIrBZ21qbhk
Kib37b0jWEgp4lDrilnCBXF6yy3RSr/9/GAVEHQqRTc9+RA8pv097lo5qmwT1QVf
cfBoosVBK6nW1rvUyFo0lLt+Zw7FzfCMvOJ/VZjtjGn8R/RloZ4hGPilPoyXMD0X
za4iz2S15YRXr0Rb6r7TrbMaCJjRurEdd5sFOsUezZBUPrQfHqHBSUoCUoI+/IdA
NjNz8SMKfZ0+OAXiziqjs4lJEsDAI9yh/wVPM+0or8f+xbvIIBhX/PAI4GKGZAHM
oecEMJIT3MDPvXDB+I8TKcP0NzX2otWagaG8Y6JT9ntlmbto2PNub1sOpiMB7olB
PmvW7BTZ8/7AYA4jvozwwWonqQpALJkird4TS7xgsp0eBSnI46vYM9uvcQQ6mInP
lmmFLHjO49Cb4ow6AiS28D4fguqvuzJ95KbdRz+do9KeLh0L4A2TvX8ISmmV7fu/
GheSnozbqr19Txs3y9fxp2GDPS93/15Y9MTTIPM7Hufudb8KxK8C1fqH3yNxv5ez
Dc0wMtgoLnCPih8ccdNKtHvNEL8kwwjKvJ+m+VVuj9sPiJiq5GHMmHgGAhA5vMfe
mS89Jukb8YcnsGu7xLGlgITMRVMVNI6cBAU/D3pBC3X/pHqbF9N95rwEnp1GvF9r
7ugfaGiR3YUY69cOOMJ2ADuyTFsjaDv1OfzeANLG3QrgHnyXtI/kJdGIFbT2SsM4
FYXMts/E1hOiKXICtlv36iQnj0WCWh7rsiR/j5hjO5DBZo47GibtHoQ/UtyIk0wM
d4DYZnVPEivUdkeKBsYntI8TVmiXlLeSR/ySXFL1jJfaERzZP2BsUWJQk5TBu7uo
8OU+RlbT0k3/nka+SgZ/mmhofinU6FvJan8oxpsv+NJ7KNZbw8hAt67CxK353HQZ
tzhSfFiTPpAnrvjLvbGmpX/zw6hfD6Y296iDDHXqK02+VUzDjYtXWuifZxRiG7Gn
yc4prGS5ASaXaEXf+hyAV0ivQ1tMvnsEcZp83/+zRIwD/uFR2SznSip4kS2KiXPf
iXeuGXZX8ZNFzVnOsZQZt/v9dfbNb1BIFuQBU+zJSzJBMQ6Qj7hxxoSj8nzhJcj9
zNf2NHrR3QtU4g4qqH9CGf0wrMrSXCGjm/rVodcfb1gOINu2IyQUKhXVdL2Qgls7
VbBDP06tdfiUuimftOkDQMmFndIU06WwP+qyLo7bH9za8nGZmwFqqwPazqK9VEU1
OEr92IgCBwYsDC2WlHKzCVS5ESI5Hf/pTz6yHPPxnAZPKxBmQws7dwyKTxttDrjQ
Q+GAGneuy+3sf25pyYSDJ5TNThd0QofgRK19mshRqoHlWJBSXY+ezT9VZB7iEqhG
TntmB76VvPAZJD4aftB1xAADcwpJwgRLOrPQta56Jp9FkA+hvQG14ki+gixfS+IU
baPxRhiot+5iZ4zgQzhF/LgBpbC54129VODQnym/Nn65fMaVOYuGEfUkxIfP3Q7g
KiMBU1HjEWINdeAQ7F1dtdTcPDRKR42vmzcc8j3GllShefytPGzbowvRWShcygcJ
jvfcTvkNtV3bQ2P1Sjzy6emdCb23ehJfc+2+0GJzJgq25tZVyW5K0denUk0a8GX6
fznl+CND0edsCup7stGmT3X+98WI68aMxn6c/1M4STY6UR/gd8g35B6fblNlZXAX
e6N1fL8hX6CFQpbVsGAFg1NIDU7Qn63k7cWM/eDXtd7rqLip39ehYQGH6LESIKQ9
ah6O/cjk6PqgLEkguewFxQRUM4aY/rU5Ip8sDvIf2UZnDg98kZ5K+pit4u7itrtL
ryUbnqwde5oS+VrjvA0RL0W6CnHiHy4oBrJ35xS0TWzeJ5pdafL2qusCyGej4GFT
GFw6sRKr5iB/S+nUHYmVu7LSez+uRxXxAU+PHhhWYFvTeYwfeJDTA2AXdp9/cf2t
FCWwUyktE6m6M2sjILTFCi9QjrOwY4vE2QMGooLgj6rcTSmZTcGg1fWWbGraTKNb
I+W1IVvYZU5l9y/itVR6bJ6HVNUoDayL0FVpvMCV0SQVWjj9c/wI6IY7+f5sW4mX
b9aTJ5YoQRPsH+IXrjrIiXGbhdbZPfzL5gX6AvP6bseUu9df61n4SO6+j0sYdv0E
OXijXrFwp7CN5DuS9W2My/uwgv3PLg9WuEQ7LjFpqqXLrQwd3A6za8wqFXY62QsQ
9WehMtgCn5gnCGm42p+nhBR9rRI3zhSc9R/1nWiZVjXVfQwrvhuLESwnPaSLvEy7
I3pdjDa/VrinZ/lSoIPxbHjljJcL9dlNQESA0/HnEddQnEWoRaujRCAadrsgUJNT
c1XTBeHkjgpYnjuELJBdG1L6yE0CqNgkOxv4+mE5tQMk/LKCPnF+KW0SBfZ8G5JB
I9Qop6eXOutcD0cnfIYbVutfB8+Or5/HEZV3G0fmB8V2Uaf23EQdcp8ubh28JGHv
4Tbx1AmQRNX5m5HIuUZqlVNhE8AW1D9yzQPsYRGa5sQV889EF4FRzj40OeDjUd3A
hGnwoA+mAewCTjnu8iCL3ckwgRVInmvzWsZm5iEZAu6EaS/CNhtQfKNV1873mmYh
Em8mUntzEn1G2F3zAf+XixdkMoFOY6XF6/8bsbnqDZvkFfYp/lTJMj3CjHqwIrL7
a6J63JJTNySK4C6m7ff7CJYUCrANpYq+unAxpJCjQhKqpM8xawEjcGJUwpXRJlN/
XNab99WEy1+l410bISj7F1nV2QhWXkxXFfp7WxAe2EcxTR3cYVkwQyPFq06S/Qx3
BslT6I2Ur91+MD+SDIhOCrxC0SzXvPwVyk0vem6vbHVBFGu0HNOHHOMt1+qvqLud
BQsggprEzcz73W4tHr8Kg+Xj9LK0aXhqs3Oz+PzchPDZvSCzpPhNGcIosj9nM50F
kuusxTN40oJvImyddlUN4AKnV6iVfT9/IUZtxojr9vjzBnZ09CY78m00baZJtV1T
mqrirh35ojkN9DiqVRxwaQUpACyt9lHWXqR0WNLsAr742+91Z5n6PxdQc+WTdgNJ
3uC1dvOih8OJ770J5nlyxrF8yqeWA94Rt2dzUwntgaogs0Rn3BSM7/kq4ymh7R07
RWM1VeI+OA5vCia5kogOoi8rIF3aGEnHgCyDsZkI39n/VsBcbNIz66oDHzTYut/9
ojKDQ1+IRq1Z4b+OduwoEuJKxvfOKSyqxf9MeAbHQRCF7aY/6OHjpD1LXGa/92M+
j2hgClOPqwh8BBChJtAmdiogm91ndEY8LWTVosM/ZxRkrxC7JOMCccq0wEJMrjqm
tQSKQjjYvV06ZclSr0cEt4wCxk/WywMWS03g+tBNm2yrYdXpiorJ92u7WdP0fvNQ
Y9bj8+2Qtits+ENcykiLr30by7ff/swtIm/K2R0NPeoNwLC0bKMdN2oVMWAIaApU
K67TJKlhWlZZN7tLurQYc/AYgOI+ZYy4cpRUQqkIWNNPBRcQHlOoOUwpjILD7B8n
3F0BI4g8TVC0nYMCqxORyvVFS6lq0b22WvN/+BPaFWgz5moyMiEvW/5LpZaBsEMM
7Msa/yl98gVOs8M8zh0WJv/yZOmbIydnhHL9iFD/WerYFMybLXZPyve0dp3kDDpv
xleeNPsDC8Nwvt+AHDWS40+Cu+X7UNiWJUmde9V/MqvLZ++w7MlScc24qDkttglT
hYa/VxqcK7m9VstaTdIzW6IYRjWZKLMMe+s8dRydL9pQEeW64kDKKhE6S73N2ACl
qK6toJojQ98ckRdFmXNEobt2m+/9y4FMm1A6hv+kknjybMwMujI4YEbBWqgo5jhh
4taa8gs3OIe8cXOpmvFWFdHwINBdkehM1zHOxHtVsP5ep+jblZD8wlL4RVImSTln
ZbQyzw+ngMZmsq/dpteoJgw02BvmPZ0RDKdbxrHiwXiisPuQSgPiWstEroEYfru3
LtU47cvAoIUShzhwOwqy/ydKaMZdFoPsMhqyd1Tha4AsrlQSHykC1gTNl1Iex2oA
Yf4gQuW5h5bDY1Jp40m5xfH7W3EHQuekFBENJcxT9B74xCzoTPIUslXIXH66odAd
0lPPgcNFI7vbJiX3wmg9RN5cNWj3iL967RA7BxG42Yn1p68x+mWT0GXqXD0zxyeA
d1OZlf7Gp8ZQ2H3WQtZOQiY9tEd+gF12Jzzm7ctFQ6u1apaX/0gJrmxR+1CZWh5z
fd7c+LL6QkhpZ1vufbpkTHQl06c0YoYRevX0VzHUai/MqCUcYaW2B/ckNvRdh4F5
xbb8n3uzzsmvfrDJwn5vbPd//f629/KvDsZ85Hpu/UQPql8eyseTlg1HtlvcKa5l
CUp0yrIeq+2qz1ohI6Y46fck7XFqWU8NHs9LFI2QUICATpYhK7i/prOB9i1cDotl
slT2YWwEfuNq7FU2GRhov9plcZ/juc0GqSefkaPK5svOsQ6pxyZh0x4KFDVMWHpZ
kgdShIIzik9iu+SDCcNADdK7tkIV8Zrxj8CEDy5D5V2NxdOvqTphxphBwT/8YU+5
FMUN6Gmbnn6J7n2nettekD7IZi2QR1C7uBJA5O+sPydIk6QReq6/AEjrbQ8YnD4C
qsybOUzRRzJ0hhUZPQ6xeC9yAjbScXEC2m11xbiyZLVJC8iZ/MBmd0hAcCNvleSd
h3fFgdKutkyU+w1dwWhlpB8GXgstOaOjBOmMvTxLD0SnBCYm/ClNYjqD/6kpdCJX
gp4hB66UpelWwwgx/Xl6IcWKAYDMEMVktFF00x30xk+scnPnwmKk93a5PYiwqIGf
EkBy+0+Mvo5rzkCnX5DjSk528lAXm+GKnVB+8VjYtQ2ww1uNB2VdZazqspK+DTQd
PocDFIcNkhIBSc9tqpx3sXemmmL5mVOFJyzrmvB57geDXNguwD1tubf03zCidPan
/Puq8iM65hVsC1OKeIUGzIn2HQh1Nb29mJc89BQWmJGD0iRdQ4/50VjTrepLzXk5
VipjpjSKhvqSzK/ygAN2+ZbJfC7ISHphYU6I/z3ojqCY9+bcEYyBLpX2o8uWFy/+
KUNlyRxsMpKbRmMGevQIjmBcj/+TnZSRTsMYnJtChyZmN/9VYc+LRYkNXd4GSQT4
wU5iCXz8xxjovN14s0u7JPS41tfT8EQIc7eL2sAT+ovVTrbkpLjTXBZ4ESGipuhh
fjbD2lLxqu83+C40zQrlxj0xtS/CbExcWkTRQh/o8ub3J2zCP6KW3cXGjhcQy5E5
n7Q/efZ96v1CZ0qNEdwdmVFXaExJqlxksQ/8y4stDF4RzLlII6YmevpGqfRfdVNq
jpSPyeHMyet6Jfj4AI/D776YU5lUXnhWYo0SK6VT5ofsLCGWLyCESvNOARG2uLiN
W2ZeH0qlkdde0eb6qktzwE0BoAUm8722W3jc899g8pNm7T+AJsDZgKac1GWx6WeL
dMqKnw7hKnGgsuJw1hvx2tFoq6z6LdRrY+tfUL98aificbI+RqJQ4kF6ZNv3jyeW
yVAObeU9E2AVMyA7ilGUb327t1AhuGBaqpPqBMqIIsYwfarPOB7O050o6bbas8hi
mTm92gbdem8vZD/mvGOSVdphcw+hAd+Na4ulHA4qIw2Lk+FhoYPWLTM00IbLfONL
3q1zCdnKXYJtUMZJA3e+w4OWXtThrZsJIxiahP9TtQlH83Es1OjGCGHanX6VaMXt
VWIMvGKdVt7tE+9aQoGXRqCnFD1REvTgECzbW16lboJBRZXIICtUosRpeUjXjGAH
HHsLwLZUoqkMr36RKjrzj2s9r9tWAHq/JlRhbHDoX/czh6pWL1vdcelER+4BnOm+
JX6etP9w7GGvwuIpIO5oUu2OygHPWhXdCPDfyMMTCmoO5gHYRU+2WLx3uzZmXwID
xw+KisOljd1lg9J1qmpeKhbBHdrG7Mk8TLPLRTgjsyhu4tJR4526ywJeToGZuWLS
9nvdVdcvX2JR9RoEZ3i+4ZUGFe76FpOK1ANqzGxv9WFPFXlPFqtAHRwLUBhQhAgl
NUCe/B54phNVTgg9MEFbULzs49H4vzNreZNiTjywmbcbRuzPtZRj0K2BAy8OVakI
vYNFgxCuS98RjTJLkj8AJklSG7ZeRyqnKUylYFOx5SQv/+jkRUwajVnjUgSyafjI
LEyUpttekqvQABujQ4+y8B7zh2zFZl8DhyO079iRw4dGNNu8sdUu9jOtsIKrEjue
6/j0W82mVQ2yjuJ1D/Ijtlr01JzLOJoAu4Wzp6ATLVnTaC4ydAU5X1xIF0qK9xvM
w4wI6aVgLgy3xpiKxIVbjVgxYV8m+Vzhh4/BOa1Ox/vgnHug0+uYH1OX34bjUgUW
O2/HL63ETxCvZqpBEwXzW46iRlXaiHAm5IEcTbqmVwwKYQDySVuTDFrwys1P2GpZ
5S1sLHT+jmSmc5hywzd5A5Oo+sH9JqrdLU36YlXhy1sY+UgDt8IO3jowbtKArIua
FEleyqLwxFfOVjmLsolMwU8v4VtGWNfxN2NLu+gZA6yYfUGdQBdT09MMPwDAo2Dw
7RZtZivCE+U9YAiEWtbiYfdJgAG0WbOCeYA4eRH86Vgn7N8icoKhbBxRsybXtprm
izKmdzGEIK4AbYfh5n2YAmBNj6/DyzmTNpOSDJafR/F3+Qqkm+BtYSeZ0jICjKGA
8g1fFJOuzw3MhXWPhGVOLdrug5igdxJmEdM68fGJ1bkHkYbRXnblZZ5Z/ZcWZ0fz
q09U7rXImjYOP9/sEaHB/kd6gGAi13X+EeW/8Y+E+bfZISbdYyY+mpBcq286uos3
/Kdtw5kMP8s+Y0PcD4dh3rm9MtqCgAaueKqWOcl7qxvAgAa7mhO7xNABn0+j3Ahm
GziSHI9bA52V5G5FpF9g7hfR1hv9UBw1mACRMWiOBmMZdeCg44ddHeoOgqNWQ319
QKK8aV+/b9U6NV8ECDtC9YTzSM1AtrHhQhB+UXN7gc95DYbMHCvsvvT2w3QOiQKX
LMbtlvpM3U63eTaIq5nuIWocbwR7v1b3txuz09BrPdzWg9Aq23sebMCldFgM6nIy
CCzX5dUP7fuWG7AzB3jdqtkzNPYe8RKhHp3945xrgIRFPe/DEoJMfomh8ljwssZz
PTNtCZiebHEc8o42PKZKTd+DN/lhi1r0v9TVD6ZqmHP0eC0WfAicf6s9u3U365r9
0O4bDVmSZMZTT99zEQL/kONrwB8nHNPg7QdV5mqvb3y4ES3IjfDrRqOv35MMY5wi
GAEU+Q7u15ImBdY2hHjHVq/YN0fEkVtlOvvhoHEAFqzd9/FdCG2DvFC8tS8DVy+y
WJmgFTPv71VuRyARck8aq5RsyZsj+SL/TA3kMyqbO6sTR6ph5MqmnD/8/ozCX9Ud
vMAhqzFAsoyHHP7KLAVkg2Sy9ZVf5ntpYBvvFrgDrbIPDOh464bCojHkCYmT5e36
DZzc7CkjQyp4UQRrWxmXE30BsneXKfY0zBnmFXxJPsmHWxsvbhLGJceLcuYnMc0W
PbypCQ3VHUAjKFfhUWMl2HRjyFh29Q8ws5bQOQDa57gPuGeYEHbdZWn6M6vdV8Ii
3gmJna0XZ7qjXjz2+oTOC0j6nuzKWbrXaU4eeBAljPi1Y0KmHdXAZUpD46w5uhQr
PpOGrDI2Cp+VGRuVp2Yi0dz7PPMmEKb7U+sTmrXoBCflZIpOcvoWhaGMRnb37/ei
+qDSallL3eM2ua1TBfcbOAJAn1cwv9Sgfpjc/adfwGRB5iX8bttns0QoMpf37mGJ
`pragma protect end_protected
