// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ecti2jeyJ6nbeS7a2mfTr4GOKZ7SI2RtO83w2EjgRPYMOJwxg6bpBQGNWquWUsXq
BuSQoDWduazyxc1aGLi7ABdymqkBOmgxARjVmzGXucKPJOuXrfeDqtToy2E0RZ9Y
c5QnWsDPQsX/oCYIx95gNcBzCTZwjWxzOvmBDNu1zTg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29184)
uEfUfWXhKMXk9FoH9rKeLdThMA0Np4/tRwWWb7tQ00RKFA5baacoUWTHmLE1fOzE
eBMdVJNAuKszSbSmGTQ4y+/5JLRfSWagkf4UW83O5UCgfY5JHnKSOq5O0Jxtuazk
wVJhOfEcNzrs0m6va/iM5UYif2FAdmhvmd5S8Xxq7D/UHjx0MOfMYtoQ6ITTyspm
8GU8ytftBt11z2FPschJ3cPlRD0qbA6v37Tncu4PoUAVY+bFjaq/fcdnuXYimlJp
trtgu7PKxGiO/igTBDDa5esXfXzzegF5AICLKGNWJB44oA0VtkWe1BgXZmUfb0fk
QhEaePfJJ1sdmj7UqHTxH4p4h+jCiTaWceU49EZWKA/6unimljdtEUL7V95JcS4H
isC3epIeucCnUDd4U+6FUDhmX7EO4btd46WmuS+t7W4BaMUvFW0FnlbLsEnfOYWJ
r/kMhFISfd01xKf6u8kNtXT3qfBXcnD0o7h/AZIvGP/G2KnSP4JbbIGkYwNrPhk/
L/lUV97z0VhTx7WbvvLMFIhkcnIG3Jx7bM+sgwYZsDqnxK2cCh2sgI5aW9F2jvYk
F33wl9sVM+5n3wE1QddsFzWOpoxzCQofa5KRrcNFYko0jecZ05pIFvmUSmEQBDOd
hlF+SQhvRkc0h8/KT+uPT/8XOuj8idy5YlSOu1PJgZruaPeK2iSsOguV4E9+4ObT
g9ZWFF7A/cR/x8JiPrjb1lQt/JHy2N9k35TaSwWiqyHxa6u3qidd/6iisepMW6jB
eX12dup5l/SGTlYtI80wbev7SjpCsddJNLDJaAEY4Te6iHQkre2pSYBYOO6CJ3/q
1l+nbQiDzOWJgMOqExVoc+u955U5iF36c7O3uK7DuX5yogeKUNs38SYwTzwPRr9F
1qcAuFrLxIhUpacpWi+8UCYEJDY8sffnzCJLsNqRXbW2X/DjMwO8LRtmUNeXhP/2
yfgAzD7bSIbkYZXJtUDjjl60p8wvzb15IpHirSRPJ+2c18edsyMj0TZsv+v797N+
r6UZPFbAK8rdlEerLXikjSDu3VAki4gkHixV+8RI10q19PvNUaO8qUb3DAcfhR9k
0S4X1Z+G+uL8cUGeZzSwahBNjVG66rhM0mIPuU2zqqr2fTkura5VPnkIoTNTO/hq
ucghwE3Svh7NGzHlKwaraSGFNJdRRl+5PI6eoLwG32+dBGBII1EyGbPZzX6A4TKt
rwpm2bT0xE4COyMBnbPgF/DCbaZbZR1VLuGYUwg/RBnTvBOcf+YIHu7EMvq7uO/R
xrl8jxt/IcIAcAa/UF7tmPf5bp1Ytk/YyzoAACnRkOSLmpxbkZRT8/EDS2LCkndu
5WI1FKYRmXTJ0E9MsG6Sei3vvsNzA+yLL/t60uYowGcRMAb1clKZ8A6+mfK9GHN3
S/2HIqTxSED3IAjFWbR0XAcKMUmN3JK8IDwErfZhYt9CHLcRxfYeinbN5xKMLNgI
TA4YZ2e76DpIEg2Dt+WpDKHSdIpENZjlXD6me3wbqtJuiNhPgKDu3NQLsmcg+KSC
TW1h5aM0eX80gCvKd5SqYVsI2mx6rJzGwe5T6ciGATGVy9UphgiAfJx4shhp9IZg
aXH+p8XnG5bxdrCreeUp34XiD0ixkDPOFUConO/fy9vI7ORieE0FZaQZOPJfdOot
BhZk9gr9f732VHX0APAWwzpQ+NoDDnmBnoGEt3qMFj1bDbqPotfygKHS7klbdz6x
bAIR6CZU9Li22+40G3f90N7MbEzfG+lTdOx6I417HVAPKZDwk60n8lRIcAi0q5gf
qLfbfJtrAzjoGpQfxoeEEhRNK6YKi+WSQ90OWSihzRAjP2Nx9e7C5QpYUJl3yp5T
7Rzrvva4hTTs+WQMROL98izF2LzDUqgHY4dySqHiep23xlO4Bde7bld5LlSGzz/b
GGtbIjPxv+iE2b6RYi0Q6LBMMyayDcykuuFP2e0feuQw8HTL6DYikQGt1oWthLFh
4zGFg6TG5c5ruL8OhVCKd4VA5B5do4nLgSPzii62YhsmxKxAZnkDcTDQP0DXwVxD
rkK4aiIwnnpU7SW7rK2OvjPAg1/qe5UmQb4ds7dTMuBx6sy9ui0is9OjKYlAtaKB
EHbKCCkB+84MByPHob2O3mryl+TSzsR8LGINlIomCTPb/p6OsAZB7f0bCf66HO/i
hKCUJUOPWsZ9bciaeKolFnx6U/03e0F7+dEJgRNFkeEzgNsjJhzICkX3WA5iXVwF
kZvlzFKwdd6tE/hKmTzRP3OXLpdtheKH+xtuHvExjdxnzVjJBAzLdG5ynThXZV27
W2skJwBzRprHvpMv1GU3dsZVe/EaYnRHPOCCu5b0yGkQbByrUup8gFOsVfaui65H
oVJA6+je5nQPmX9U9Z7HMsGSB05EOiHiwoi0mJEFNJPw6fZeW0+kV0IWVwsSlHq/
vGyMVT93qpDU2p9l96vtoUN4hSo7Rg+ZFdkkWXUiZ6mDhluoBlM2lKHZbRC4QqVP
U+XetwpPyb4v1keMuqBLPgr8Jiim2HRqSq1RT9YtH5eUFfdFvxy6urOofOFQmM21
Ac7k2wGxaxaEwHejtCyMJFK1aYrM63PPB6bcY6TltlfvpEQwHV8QJMOmqgWczOSi
dnrWmLi2W7KKU0Aj8nKzJmgRE0VpYufHa2xNkgNmGEIzXxfEutzbWQQUEKuYXuFm
MtcetB6ErZCCP0iujGrVJvXNiya0ifatPn89ccJkOLtWuMZRCenyT+lAPl5niWvq
mrz3TfFU3jYDT/Vt14/QH5D2ZQ+LhK4jCZV1y3mHmezAmS5zqm0CTKOkTfo6o6nU
zto6lsFbSTKchGshyMSE1Nyc5DF5yDq3GHSjHbeK+Bp18ro4i1gY61P9QM17RwJO
eWmfTBcNsSbjAAZRZS10/HiVxQ509ZvutAKBjBQgbYXlXs64XRIYaIFW6IKKu+Yf
UseXvstnsPTm1IM0MJq0PVO1afSa/Z8vDOVV13J2yzOoQvw2Z+h/r9JPk3lmy9Sj
kXg2ov734vQx+pXth7fa2TmIYRIDl19JHjZ3lGUsFEzKAahK7AY4g03Ov6f2vfPP
FaPuoP1L4tK+9YrOrLgJA2QxkUifcVTFE0XVZcKOYmpeJ9HTal7E0BlJ3hB2H/Zn
W58CVSnOylW8aoesOm0GfgXiosqdyAWaKjHs3FUPfO2/TwVnZnv2m9HodN2nN1Hg
tq48beCPP0HFy6g9UfATfusJAZNcFXPZX+ETWcC5yOl1U/qHPZAG+Tm1Mzgnr69H
4p5NCbjd53m+dyZWe0MzxvZngyOFfwwBXjHih9IDwMmsjfueKpBpytVVvTu9t97R
DYdgbvhgo85pQKWwYGFL3U9qHslMfDKwA4eF723/vw0WF28qpxyhlpppVq2O1dKh
9thfV0TayoeEXM2+IuhQ41cSy26ILmUf/+0Bl7P4c3j27AZ1FHJgWlaxVjJDteCv
bezhZdEnJNKeUbFAoi8aE7vmwoR5hBpcNNer/+8C6kgSGOngd/aOZ38SZP5QQ2ko
88s/vRBbY+0fVJMsSR7OrxElQUZfT00B+zjMlPmbset4EGMSuRVzkhL3VJ8ZDc7L
zp684es9kkwoab8h7P9x78HREXOizp7oxjwdf5hxyuyQDCVrRrX0n5rptalBiCks
4rPgSxor+uHQ4+m4/0bnWq8iwCTDyfsXQRduq1WBdz78CAaS6HTLfeaLJ6KMuq/4
73O1aIfjyEA1OS1WzvL4a6RqZSNyPWnr+Waj1WTDOwxBl+Zvdz5YWTC5xuxAIaax
ZkqCwzDSca4aAWisJCe0KnfUvgc7TS5aLMeiJxsy2pFHRr6F2lcxVv428EGFW/y8
gmzArOQ3ItjrQTD+5NyFh1nPFCXjMeUJWaK5FvxIixs4+Y8tQyorTeP0uAtNUS7h
siXe6inrh+9WM21ljKdCAp0bRYHwNGQLtaCCoNc94RXxh+F3fsE230rgMnroHEXL
13GZYNCVHPfu8VPsHRqA2GtfDYcb95G2DRgVuvRWhmXVaSbminU7IxBWi6NOgpCY
FhVtqdCs1maaKmf2tMD3nZoX7p34HPIGMtASbIcOaKGhyXTZdolYJGeC1MGpoboK
aPFslAyUf63F4Bzw7gMJ6wtsGxd1v4DvHwYYNPxTzAmmkov9ndHuHX4MZTDIYNEW
DQmDiKTxOfkx25/E4U2aRcTs1MPxSsgAenzSueVovJwbYXrCjEIa8OYuJegM9GR8
LcRjrXNyUOl4xV7HwYU3HjwQEFBuEh19k9ksgoUaZknkap8otyMZo9rUe2u+SBQe
eLAsD+kGmD/oFiDGPrjgEGKPqDKWAI8jQdmc/HMRan99/phAPKqt1A7c86vb/G8f
TMHln28iydBP4MdnSCIuBXiNdFs7nCXFKoNQK02moQM+RKgtqgsei/dbvac3wqEy
MrrIBwgSgNIMNhYDew0zMboaJbN7JxvAcVmJjqnIvP5AP5aAXzZ1cW9JLH80eGT7
h91UhsMh7biFD/QTV0r6AxuXOpOK+c/UZ48Y2xhe04tFqv+yjXoTf/zAQ6uxepLK
4K1l36DQzOclJ89qSBrSOX6cqFSEOTq4n1MP+dQTzlmT6eML7Hq+qPQgCpRuQG7t
h49qSAov4CDn+to+Ix1YQkUkNhPSTAJq9uYy3H6R0ksqsIZkB64Y0inOjijBkNpC
vrhWmmWX+2EhTVPNx+wf7jrwi8RR4AaztPDJp+it57t2O8nRC/M55TOWR3L99+zg
WlocuYLEcnCWDzbNJqw9Qti+ctCTa/7MR2h36kIiw/9rHWODirSZtLAtcW4TkauG
W5yoQTo1fvsuBYGu9bmIDNLy0w8cA9hNy66wX8GX6v6iMhRmwKtkLJ8DHOUSh0PV
u+p64ingch2SFmwqUTxmtfP70sZBn9dwYXkGy/EDsFpPVBm2mokmnelPHz66S4aT
KcLiUaoy9e9gvfwZZD3MCUZCi2hNKbXJzHvgc3wC4Q6ETITevx8KKhSNy3KSO0YR
1T8aM+URLKNloTz08JdEz4XSs8hv0QwRkdzv45KH6SGmyaJuQgUBcCOXBG6fVZCu
sdByArZ18JJsvob8/TOUph5Ir29xbMJqxVrgtyAS/bAaED7Qp9Rnz+G63Cpf/DNw
bsfBr0+BDLAFvYnHVJmvF+iMz3gKM9tUAq4ZJfXl7Sy4E4cWs2WKnFuVYIUTo0+3
bdJYkQZzwJ2isCgUi4H3zw7W25cS/yOziChw5/PwUdvtHoQHroSk9HK+hbvKlmEh
KQeIrem7gpQGXYxkxVLOHi4xZNwnGWwaCPrx3ykbxnePXQjpjTDDgW+OlOidLdZo
YAtUf+1evtzi4ceMfZF+N7w7V+vQX8/jdFw1zdinnfI/FLswi9K9PpB+CUji8qOm
3omWvhi7MiKbnC+p/dvz3gke/ZyrtCayhuJ7ka2I3gPZki+OZ24Hb9krFzHwyJfh
T4muZkwD7LLoN7eSIQ0zEEnTsOB4j2ML9SBsFwqwP67Su4sI2sgRvCAaPh/a3SJi
gFRG7UBdc71urz72VK7B4FMnue+P4gt9MyJfYQa+nC9HOPWRsL8MB6574ue4gnM4
jGT/UdM11r2fwnt/8m49pUuE3NzjSqyKhgrtKjOAdbz/+tWhs8r8HP3laWYhhaOJ
H2DJi6ctuquhdAT6okD+PqeraR8XckyySrDH3Fif8E8NNTwtAFQnSTrqnZ5ozT2z
tVABqvXLSbdPR1R9WNYt7gaNnghl3nAV0V3Wj6N/WDC9cp7cXZrH6lzeuXuD87Nw
lbpTStJXYOWvRP0SD1Eihh4lAYDqxvw88+OF3pRejabhJuiWnklNdMiZslMXSquX
kXiwu3/yLg4sPPVuliTFk96O2GuuIlQEqYYFZxbiBAfAUW/rfSlbxnabq13L4v7Q
1UBNbma/AmDu0fFjwoeSWW25djzAQi3RTmwU2xsTPxHddlVnNZg3TWZXaV00wozk
2kdXn6X8R3W0ImXAVCgJazSYJl/ZuiRAQ/6y540/CJGE+aymOPIY/FngfP40jef2
H90y+W6Q5kSjdM5/EgXEmdUTxq1pND31+g16GqaljXRbOWz7S13vtn77tZOIU9Hk
bV8y0n9Jp/ypXoYNyayItjX0U3HxHuM2hTu2pGFo0FU/09WM+m9AelZyX7dd7dcO
dx0Quupkmdkk5RgHBDjJlZVCf4nj8wTAgiuG7nvAkunllzPs5DWyRW4EJE9UL9J3
FN8kOKifhwI71sNgwdtazl4oa5mYLqfTBCaCXKFsyqNOWh37QSbDRJBS8FcPbnRP
NWtfYaRrgl7pTdZDahJ/RE3GyeC7j9x06FJ3G4PMfxaaobMCRypV+J4bgwCH/pkA
QsDn10Pb4nMlyk7awlVmLOAo/G874GT494ze4OZIwDkUXkkAyQCXDU6SzxyfN+po
pumMTgrMEyQHpCxQkpIoeoOooHIAkkFh/APW4w8p3wqFMjwgRJhz+kXDm/ejQJsf
Z5mRe2STmPAoqyzl/Z22kO/30d2tVDzZRcyFCarKMC9ECzujr//YXfGVflDLNxXa
O4FJXl7cGq2KJt0CE/R3dEnmz4ipvHVqgjXS4okUTC66JbIhZG+TUDiwe5ok0rBI
FIKbvxkcSv9pKGmyt1NuAi4uLZOf2VBE+iBKQYOxc/rHx8kGg9OUpgloBSc7EpZm
82CXlBjd5z2WugGb8XSnkMONUspyg3bFn/DFQbpgxTDw+LBavxwdhWt4UVSzR3uu
L4atHA1nAobqoe+hWPr8Tt/GmgMDsPtKsbWVghJ7Vj18F/xLovAsvT6QRRzHn0gJ
3sly6laT3VZQjlmzre4hOEscGroiqf/P7ahDYoa1BFgcPts4cK8nK/yxN2sdJ//C
YjpV0rXDXLZP4+QxPcrEfNuYhKpnJ99srnMwnTMwFaLP9my35g3UamP1zK3v6kxa
thSXpQa/IqWVcYjbRG/DyEXiNKFKQZOpDCOv3tu4iQIgynJbXYZy1t+7LF4PI2GO
nziJRGfksB9PHegHu/o1hx4sW23u/Jy+8+Z/gPny1fgEj0tlqh3IIo1MgsurdwLJ
1DpodF9fXca6diUHOVEJ1LZydFa5QYMGa3J6nEUc3QG8na9Zq+ZToG9otrC6yZjH
awlGGrUGsA9i26BQzB8KDvO7ntzLvY1zVqK29XZHalZoWKGSRbGL531gQBm8NxqT
qmNfOQq5YmkIKn8+3WJFh3GE1R8dDDF836Kb1aYBgM5xcbHl4qlcfEZgswwr/Cox
82Pciq7IHeEHzHhYIZ73hmiE4vVfIKEvcUCy31Z613jXJzAfY0Kktk/sL24r7lV+
ZtGkZDtsQr8Vqv8i+lRIhU1u2zsrOjlP4R91TmXqFTljSPs49wXrHZ9J503d2Pgg
Qe5y69+9CSTUeJVOderMr/YHtl9kJakgJy43XZJViUfF78R7klnCBRic0fqQx8uZ
KpNvdX4LNg448IYWH4rHHczl33yt5qByQd10MsYWkH2jIZSKioUQoX4/xilT2GLQ
T+VXwmNU+Ii3cW+JIPASvTYAmgaAIc2SRNkP3hqIMdoNlmTwPUe6hnjixgmyGEll
ffYoeEim1rALNtohOfq+HCtsdziBNPA53xRGRx40iurMJ0fGrnGiqx9loQ5LSriR
Zwc65Nq7cV2441WoRsRpwL1ycfQYScI+ziUmqa/Z5IkFozyw6vLjVl2OpCz9xHMo
Kge1vWSY6tEcd8fO91t2076OdvQeDmxjzw2922Ll8cfOF5RAm9j9fkMAIrnhkZ04
/kFn4/rypDfccoC5gfvBY9ynTNHwI730lxriS2QDDoRNyRrwi79HA2VS7o00g9E4
Q07WbVzed3EXtgpkTr7se/Bwbdm4Nc0WsQgkl8iBpM8sHKznwDme7wO3bT6fdiAB
0wHKkbejyf64att46/YK02h9kxEce0bJfQ5qsti+iLBVtrnETOcDRywWs62VcptZ
GqnTYx07yBJlekrb/Nex8pxKSGvsC60xqjDmMrYvc8MDFhgPmvCYrQlVSY1n31yq
Z93pbJa94NOXyU5/OWOyUIHAWAqsn2nUnHVxYoIzoyuphwiCRCOhCiIvDHdgFByI
Spajk2RUlX+cftOssNAm4HBPoX1QcaPru5eVnZXpv7ZP51xv5ZUwc0A7lDgBO8ey
iBI1b3JNwqiIV8VsOy8Tv1xX1BNiR/GQOviF3iqEFqolFJWqQHogli48I+gKHPyL
m9LDlY8mploWikoirfGsG5V1adOC0wsJ3lQ+jhESsDpifn8tmmuW4Pf64wr/KY+3
hkNX6v1QhAJWqFIbwtg6M8AC3dAHEYiiwMb6hSsSUlRQp9br9+SxzvpzNyaXWIqO
oRW+J4WiRVFcygH1YExVa6NhgQb2H4HM46fZq9Oy4DV+qCRAkeCFQ/buAoWwFrQZ
VVCosObyvYOd8uKZJC5w1zm6SkjjfTBHkhrXDPXorKNUB/vwdsQEyxOK0vHUlBme
oDnyopKAgDN0Ku+jOpx6j8jItbJcl6XllqolpE9LbrcnCENU5V6fGJ6LJfc0dBA0
IU8sXkzgp6ndPnR06bbB9Bz72Rk4Pw4Ejv9Hzq9UcxFEeYGhxiFG8nssP/08UVh9
rdipNp2vSDT7JSHFLKD6/llHCG95Z3IRQjC4EStLPquXSjrttd51UFSg0rLbnE0b
YzuuTOkvrA5Sdtj4imIf67BcdslBSE9iX7hZlMMSE62NW+Csduh5Ld3q3LVytaF1
OaCV7y4YRMPUGZatZEHeR6/Um7Jv+/vjLbhMuadHvh6rqQR15EfbcnKUWzi79h2g
FwtsapphbWHM4hqaag1GMvPT5D2nAXy5Qoh+WaYrudZa8miLCEG9aRi474YwIZ0H
Wfd7lA/6uTfv9ot73W7gBvzMglxxzjjzl8yW5WCwP1T1yMz31RBcsN727YaRZfvU
YNscnpxlAVe2MNLZoCSGrTL1nbWaQKBCOro17+g2wan6nJ7atGSCHWJV2vph907K
WS5Df3gz++AJK6y6+zdcfbtOjfZds0sIYyQ7LSCINdjzpGpKKHmAcvpBDqZElbju
6gXobfTRBIoGJADHzTJbTZxS+0Z3OhDb3RZKljJUGQLp6gDQ1EksUzlxE0a3IyN4
OwDPAKYuYdPnKG+ZQDQj9ZnDsTvvufqwfLl6sBGoB+Ijkq7Vldd3gpE8xioKlGps
UvtcXOl+x6lC8crkWyJJzK1ox/Idx1tzZY0D7KR3bda5YJkm/uMmxii5KaUJ4789
vkAs59l2kUBpGUY3LBh2TpO4/V/o7GY0TWu+dJi//q0qWnp88J+HuqseICkCnUB3
UU4GQP3qU4IHO/AlOH+A29nbz3gknPvUdOM5Ap0A9vl/QYtm7yTLHJdV9jyVCzNh
nRn/mDQx8xjQFpdK4WAkba/NTDPANfRvJouhzJ1DH8veDmlSic0/KhlZABsHGr7X
ssgS2jSb4Bq9yuLm2r8wC7X/rWP1sfOG+cv5UFKZ7fQYPW4MS6e57jy14gmZt4hz
ftLIkX/m8TaOp2yRBHd93smEBJYFgEBu4Xn44Mj5mqIY8q1cvYSktpw8/HnnUdec
m4t9xEzaqzAVxtxTp6CUfytFbE3rtvSCc9N9JmYo+BBACnmVT5G1NZJ/gZGtV5+5
lreR4Ol9/m5u2aLdL2vax+uELuCYcsJ2QeDpP+u2aADAjghcowSai6TCJ2lCcUuV
xxY87NM/op2M2H6i6WrvIO8OPVDbqscr+hks7l3hauhsNMnv+hUlo2YqVyGER/4V
2ANIniH4vNl74SccETcp7m1xQmmps1YYWw63BY/c8IcdSpPhQb24TN2j/9CCQqEu
biAIaJpUa7LCYVGFTrgZZBQaOnf7TUimzVdQyJP3pbwyMN0pVAwpHGUMcArJTY2b
eXa8RYluVgtHM3K5MhH92UEvQuBDLN2RQ81sYwSdONT9V0vly6xgKXI2b0H8iihi
F6mJQp2mD+RHXqxt0CSfyiTXGmNgQ7Pil39GkxRD69URVQCkDi3AsIwh3myLPPYi
YatS8qseX3OH1bU97lZ/T7OnXeikKsumXyOhPIxbdjClx+F5TrVvfPaIaYPcw/Ei
nwc3U8Nrk4qpZkQinCipgOzwph0SQiLUQ+JalyK1HBmqGrzJsVsLLrsPd/Zo1jri
+m3dW7p2KzILBV8k22GsOF7Q4WN0bJzm3vHhZTIiYRhfcscNKQQls0ZV8z7FBdRI
MIiurVwOHvUr3Fxtle2uuiIbbf8BiuNH2FUvVMPlYCYs9C1K2GlXOnVNFLtH9MoO
hHu3IGf3sJg4u1tuwMwqAlWIebzfw+z5Qmy+s6sWZOgWGEZkzggTDq53Qlbo+Cp/
ABm/pe8hYZ58cCjCwvwWknecqyJnV+frtpiGcG3oIbH64WMpKguBDVTlhLSKUvu5
CW0kh8Lu737tS+KbgCNWBbvTE1b/iE8xuk5/8Ay68EyltfAOliYKcWdFLfS4sOEe
KbrHERfyOuA0CRg9zWOUoS0QQPVmdachxezXYX1eGz1JUEqink75NKf5OdSx8yyi
2ARGra1m7oA1RS+e+PxVJvTocpvyFFr7n0twrm/YFcwISjNqByUDGKD4MV3H+bgB
N8iOfeAjmk6Nmp5Hig6Df/ngRza0zhN4n44t1xmjkwUf89K0yUGKfVuO4HgyZtYc
RPYrqDyjSGZwgAdRvSqBinXeXlKvrnkyRin/5efc0nYuwQXOmWfSNvE6Ac1uajY+
RQjhxBBm85aJOuWh677X1YJoxY0u2fKG9Nyy4FVTcpnyXHq8/cy5wqT6kIBjAPTq
Vjil8g7ghyFY2zhfgG0QkT8xgRh27DfdntX6IGyW/Bp3h9xmsmit3zUpC9Fhwz6H
I+TcmMxGQ+07kR5OjF/iCeuqRJZtT+xZ5Mx8R0098ufyF4iON/HvQFWp9UvzA8B4
xuhkiw69RtPo3q4ca6XTRDYyF9N1yTPVYPesaynAOBS/FIIuyKDBANp6IM9cDNv5
zwp5D40LhrWojTz5nY29sPl/18iJ2jftuche+pWT7VbZPsayrsGAKLnPW+cpHnO8
SC953SHQgJkL6cY4Otmx00k5+fukUw0F7t0PfSi/UDisCeUjqKO+zfOAr8UUyzV1
zHcWTyTKsPv/i/U/RdDgWq38nw7Rl235YIiQXMobHcIp0TGq6S0DBtBzlnZ0NHrS
5EDdm7WI1CDugmentDbgSVB8spnJWcc4gbEXN4L3lxaJheGaePhsX4wJrmW5b5wX
MbqN/1H7V2g/1ve6tHGnvA4u57xg166ndMdn2mHCGTAO7Im/7aqaZEv5J7erxtLC
gftXrSrwbX7/5QUpEWsM3x/QwTy7aYFvs/56J+VvYO7a7iXIVfaIfcOrykVwahCR
syxBkD+03VkOiIxK9pAYm+e1Cu0M/yFnWCP5OhILOvYG84PGkekvJ6lTM12oIvNP
tsOqYwtCabpcVrOgTfKPngqs4YAVGUOjaT7zMJf0tcNANA3X5dd5OSRqENI+sgvz
p8Sao4M9ZrlOq2zSs4nm8Q9Ie7OYJuZ3ZTEHGS17mifO5tFAcum0+QU9HkYbW7YF
0roz8PB44f+IxMdP2WkZy7XUO2zdpoYSh21JF27D2ZsRdTCrFDv3zBfQvQgutfKz
n5wX8bZ6NjwVZOiuJf42v2Ew5hX+abru8QYAUQaUebtfCKUhg+ZlikO+lB8mRF6h
v41J+pNFv4wnsEwQfp6OLMqM4yOfyBf4VJwHaKnNwoxLasbNf31KK+MSPJS/7igk
zLIYVjpRX39FYQGyeQC5xOAQOSSqWsXu92oK3Tgvyg18A2ZCbGI3we+bW6vvQ6oO
aJKzU2kL2BCWe85A+It8YLhJ+X4/uieVVQkefO5bvLIpIcg9Vl/Y88UbeaLPbgoR
WREl8Vlq0qq/yUqsynv47VwXKpLQhtJ7U3xXmZCCONdimpJEZ4OsvXaarNPz9xvF
SPJRqbdM6wsw53sfzun/wgBECmUDJzbi2hSNjO647repF5ybqK0fVy4SbmRiyllB
HsB8JQ1QUY7KCUhoWOT4SeGlGYnQCj7I/GuP8DVmwTJ3dYMn2V1kPnqzyYjaTxCm
Bgj/pPEalZo1cqlAr/1Xr3zxFbqeL4/7QepICqOJDT6TaBID6zVzQluTWoFXfbCt
xanUwufitAvJsDWbN7rN2Xww01UpEoCqUR/ZMcawdNuc8K3/DCBbFNCGYgA6RI1M
OlCcAnV/SmwDxGmUp/QF/kxmZJZUEafPaGEx1ovAlnUwEYavO5yZsEZBYFfj4Kle
PC49mp4uy6dexhne2nYqLHKPBVXqATYD9YCCiW+o3hLiwqkLB/z/myXU2/KLCr+R
4AXGMlBiZszFEyihV8P7qU/MJiQU7fLaKeWkdC0neOV8OFP0FbRrw8zFCksyXbqQ
Srd2xzxz1g/hoWq79c2vs230EtFgDkOaq7vELjHBMSlnzyAMfjTNCUjOMdOd/Fq6
CxO49QMtzw82KAU9VAhdm0Czy/YMWV37cdKDJCPK4wPnTkJH41vZHKDF2zxvLJdi
zmldRlgKKaMzQo3yPjLs+r5fP4KpLoirZHwGj9rgbqaubbxDYpkO+i5NUUB+wxTr
4ncguVqYu0LtW95Z7auvm4/MXFoGP8Vnh8fXAhQrTUA8qlXnXwefzef/6oXP2NOe
Fyk1J/MESFcxNlNnBNl1e63zeAJ9XQCdeFMhlrv4aIuqBS+UFUS2jl4UjKcWSE6L
xpASk5gtZfGZRoq/DME5Jg/EtgEWGftmiBpx6Ql9EkEl1cs87tCjjJc8HDEGIdl4
mFRQtnP1z1Ku/7z/BQUD/OndvcAYbYJHIVUVNJfPVRcVbI5V5qtlkOyxsn9JUnCj
yFnPhGVZ1NfgVaXFot4uunj6OqviXokQ4huUJBk6wOdaiVBINr3kW8jo+YOCbxsb
9cjI3DAqW+X49L9fGbvJytUgYz90fB5UnXutb6rAmJErZ5z8UatQOo9/Q51rqyBN
s382Qg3T5hWqEvd34nfReihNsXdL8ED2x2EnVxMuSk1Sxamu28ZfurVMhn28fQmH
t1WCGnIzbTwseJZaTs6yflmj5T4Bo8fj0/A8qlL2c3V86zsJB8y6RALpqXEF2PkP
PvzVGbqAoszXdXtF/DBgE+2Oi54XGngbJQvDChVlnPyQV32WKq+rYoqY1u4JmG1d
ccH8F/ajm38lqiBIDHiTaVIn4xzLXwBgyC317+epDsfM8LYBaWdFWXfnbWF7W6/t
iAbDKs3fpy63ozlLMaaAsGBsSWVEHd9PUniEjGkhfYOp/mQT3eD1krKcnBj9NaJ8
swLZJRIKTdKkKRjH2zlKPAVO1avNRwzKiMqeSqdYW3TA2TZmMzGeeKL9xvgwr4ZR
TGGclC/b3yDeDomXsWCJv7rchiQNobx4TcO3yLW3CEzDodQlGbObGz+/TOsta5ao
nh9tDsh/toXEz5lW7v6gues3oV4eqTp8EDRZ2DRpohVjrure8L6meiTHSkkoUGnw
YVfnbAEPMNM5+3Lz7gTA13VOD3GlQVRcUii0I4QAIzAhwE66ntLsjYzgVt94RFOr
x5Xl93pA8J1mM9HTl1ixG+AekYi87grxVYIR7TWYxxL2vboWRTk9C/Havns2m3/1
ZnTV4Zsq2aFQp2Dvv3Q4sKTrmQSugBUzCS3Oxz2nwYm1/Ryn6+AFL7okEd/vPbRV
JDvtJ8WCGy+wHC51Bfet1+OfpMxfQbayETf7F8ipCNofk9djWiSoNPy/goUINcQP
ZlTFLCfkiy8qkM1sRWHyVlEVi8WcQTuZ7bL/P+kY7cyUVPW0KjIzbZHFa702pdqr
foRKH5aMeZ7F0S8pjl78QMlHSDG6BwKXeYo62D8nBSjpCcCYAEtUNiphCK+Ww3IF
euyO961V8srOdGYyqHORwfYUioM7kMh0UFECmKO4JU4J/P3UtG5PXSP/367mRf93
EFVKYmKUvNSOvnV94DyBD7BJt053eBXspHphuf7k+MJZ7p4pG70kgb/BKiV5lw0g
sXwZuyqt/OtbKLembOQlHZqf1QyJmsLxJxvIe2MlhBWHEIRuvoOsaEhshN+FZ3ki
0U91p1lS3HafvzcSyycOWBU+TS61Cwur7gZ0ufJP96KIuBmq+nsdadPEUl9Q8Zrh
PDWTY4pqmqNHOHxRNGf74VhijxChBxbcnrDDHC9E7XjY4hBnWfBi1qjf6rm4nssy
TLae/VgIxFedAqLAQ8sYcc5HvFgE2j5uTimieR7NMokwKSYwVSdRgBVendAIJG11
AHm6YvOtpM3GmW86UZH1AHl07JBaPEvqwNQ9qHMlmaHrKpceaMsLxeCEG2U4Wskg
49fvUkL22+3k8BgCBMLN9Dgu7eGfIKR0nnOCRh774aFtIq0/deSvSE+V+NOuDL5U
5ZXVuWPQhO1aKXLYFlS251Sv9E/1xWCUq3wQa7oQixZIA3yQApxFKMAFyXuLTPx7
VrCcb4BEmyTzvc1LbuZew0K/+ptK+lRTikOUgcGQbZLCRNQhTOGmMLbVn0VAerKg
qDeHiH/C4qO0IZv2TIFUSFNgFBDhofwBQ64Vo+SF4mzzhvr3pDPOe10LgeJu2Z+W
SBC4YDPDJmIU+l3GLZEzrKT1WwJ52IhCo34U4NBI8XTXCGKFDFb2vqY/b6OkV9tB
gKgfEn6Y53uGyhV2EYQ3z78dSlY026gnHCLSCUQBcuOxrI0R8cvZBHyu39FoxBCl
mHYoTrsmZYCkC3brb+qxb0bOPDE5wwM+zK/H+IwVXRjOu3wML0hj03IfDj1N6R0h
D0em2KqqLIYkfEM/DwhONz59omwQxezHrz2tcLyTwlwDDPQLCRFeWZrqUTcGoF5q
FJd6NI22mj6YhBw4Roer1s8Dds45vW/lFXUJ+QeOw+Nmsy14KgasPnAXI57HvLWa
/rFAP1cB+s8RhSQoOwOytjY5WEqtlfDEMzJa34qLyQ5cqd5bbV2i0qzbav2NHm2k
OeKZ+dKoRPMLRKdq5EBDir5sLLG1lkECt8T9sLq8WkKv/IHwlGAvVAIOO4eQ+jS0
Jj3po3bZUNdTvkpzb37IqlPlyVoORFddD3Cx0l4bsmdoj5IHNBraquwsiSbcPWGD
R6fqhy5MaA0qPNrBqmA2gNUm8hfhnceMVaHdwHGzheBOag2IGlNh+9VOdZm7hVn8
H4uj2tPXHElSBStOW2UWJJBIv8Htxz6n3oLo/cqN7mT0deLkqIsuFtS/IMlxtzvo
XnXVrNQ7/BXNpj7VtomZwMb/mt1/iYzfSMJ9x3Iy8LgpwJIxzHy4pltrxHToSvcI
I2xxb23joL3RZnnQbRL0VekZA67cwuBZXWvVP790alZPwuWt20MrorTzYycwOQoI
ceV2e4jRcohiyjEkf9FkHTablg/Grr0wSLrSvvauH93/odQKR8Li3vN7XrWgmfAq
mTxHTxJYpDMDCp3Fz8dj+oyl8COaTWluMzI3BYg30+NNtE5tyXnnpeZrWHa3q+fh
1GHUIjjBUP28SYtHcrG+R3vq1BQVjGzW7JCKwaNBQT9vQLE1IMT5d4+Ji2GRX5Aq
9/9Mxdr2OHoruVFOHKHaN042mwiCRF8Dps9hZg9mNDOYEqgHvtA7UTbSI7ltSicB
KPt5nvADVOHwnFMn6mjkqHS+n5fIbg6XHZOPug5zVCb0dKAFR1odhtU3jQvwpLuE
AZmLYfytpRAzwy7Sh1xVLCxkzgwy6G0Q/12NGmSKTc9xLzrPKVYnrDmmRcV9a/30
xvrrWIaY7losqgngFNL5ja3XTJYN8kWiZtr31iuAe+tuUu2eXNaDPV/DHV/kVZSd
9kxg8Omb9rvmVtxyfG4hFu33SBxXtQv4N24dErJcXXKTE8ApsLPnaBT48siMSi7f
4cWvJxkLt1K7hi/oKfe5skGLaIjP28ZckkZJWux/v2aZAKnoi0kYb5JRGZ19QLUM
riuL3tLXXl+tsrig67aAerAuqMVfc9gp5Gwf/36tRbNHs8ot6v6aQ5hbIuA4smXa
O7LCa+YnYF84OFazvcoEmttYzp1r9hrHuwPQqBQjaP/Fstm3HNQKFhnp9fv/vzYD
hgMUPTdbbu/LpwERPR5k5OkV+dfoKHC0ShttgZGz2GAf/ESsFqhPxme+ussV3lNA
rXo0R5xC7/JUKklpFuiAA9ic5hSub8hgSR69qkgDAHVhMRb7NC8MqlHjIf3bjtH6
AvfwUCysZC0JrhFnJV8Wn+CeE7oeackBdKAw0MQk4EZAMjhIYbwIPJbApMREgZ9s
eWB074+lyhbQa6vA6vSnYwyXfOFHAGvNBnOVnI/Y2UiN817wI9A/T2E39KDXsD5/
bzS86oyZc+JT7wUdcIgugoTN80xSzY07PQZLXKUSXpjG/EocYB7esQwTfQNBUQ2F
DijZRQgKSlvYLyTZ147OFY5DHUO0ooKAUDs/HnngbTi6BAn1j/1yPS/C/NNdgyUh
WGfHfr+X5WujyhGz2NIRsW5mmlAz1kQnYp55bHgjDVbrJ1ZuspLCMmdKy3FDMZCt
60wkCKnhayfery+dSq4u5uh/IgiANO9xMPXrQ9RHUtP4P2p1tzbsd+RSoGLN7LeO
GR4+j1R4uSSK1wBxyaq4VgIYRSt6IC8iZ3XSjbmp4/x+IM/gmlj3YZQDc0I3TM1o
bfDIn9KDMMCEw0G1Y6U/QlHhLdAYcaL/UEy2+/IETx3cG+ykRI5/c6bfNr10FYK1
XoPvc/x/A81mGoAxBqz/C1W43ORtb0hUd8oVXn5PpXjm/1fAjD2PxVlFuJEEWXqm
9OmgFSK4whd5p8sCCbj47xkbOgIb8/Z2w+jrXP/cFIUB2dZTqQeXMmkhhjRMRxzi
2n2hP3KUoybMLesyA2b0ojhddYW/kFGDZCndzN/wZHPtLvBlkY0rG6jAGGFb/lp8
9B4c9WFy4FkVnZLKtmR1y1psCJpR3qAcDxFusBh0G6pNnJauUooVJM0kB4uzhYGE
PIv+/Vu7azJgIfbKSy5uSt/mFURfHBhdRBopWZ/EA8AL21X8s19POd7fR1ZBSGtz
foUwo1xMTT94LItF6bqF36OUImhSHb9MqePsoC49WQOTgQ9kFO6MQZ9de0gNJ2dT
x2SUAWMSisaRP6cJ7HUYxaynTpxdu93rexDuOedQPJJZg/B4mGOCgq8gwAN5F0lC
Azi2av0FtqnZxTLVsgLATMZrJETLOBAL/ZE+tkN9O8kowhdvrLyr6Fxk9Tcla57/
H9H894SymgIp5iiGw2bq+9xXTaPv7zQha3vaImNFABF01Nr0i4XCZZxv+N634QzW
2KvZPSdJQcecdQbKY0VmJXqplW1FgggE+/TBsbKwaILCvvntBXX6Do2Zxt+OBxyL
v9/bo79Jlhh7AntdS0L1pboU3BI8F1JT5jVoAZ1bvZERk7h0RWzFhFANjNk2CRxe
zM7S6QYfamS1ydsbLhEbLtc4vaFx9AVCJOdNKI2XB57j+cfjJIr+27V0J7g1noQB
RZo2ClObY+4Ha5SdbWhmzySwA27sT4IgKC4aROmEfiy0cfFnZEM6cMACHb4wdnJn
oNkZWho1VnKedKcmhBp8cybSuLZZCjTfbh6Gw6PwsTYrdZ9Z00plF3FfBpdDc2M4
IkxLHpSod7pyxdMJfSNjpvzcKUTbY2aIrqGfgE21cvFOBd6lgSWFMKIqD82i6xzu
JgIpxwLITDc64QnW8FN5VYfb2cr/skdAbi6FXcm5wyZf9nPrDkfaKNpc6V2UQS8K
37nngUyTVq0qef6F88VwXbaXrD5bIPEjcZ1P54ikUstyhrkGIuaEkE+/eXJKl6KR
asK4m60yl6VdRrHUMFSWkjh+qdONogdPQE+4LU8TAMo8CQyQdePq5WdxPQtVbxaq
BpEsditHFtmniSBfQ1+CU/mnenfZaXYkqI1UHiwneFvJMJHgspsMjEUblk9FOpCb
NGbYFpbx0eZn0wtLSKbQxXXTTMWn+w9F4JCkMzhiyGRH/Imf20Y++EXZGgDaiGwR
qQCW6v4ipO90F3u+jjImBLd4xo5aKB8L4jT2c7LceEBOTGpD7y5/WFBAImx9lSnV
uFlFwx3hcofryySKn/UBNYAhc3612rca/Oz72flqqed1tFP+qrHZtt7PAHs9Dc/h
Bm5AwdL35KvAy3I+YYGm3kbt31DISrE+TxRV/NRpkxzj1484oDmxNfuMNCja5aRM
oZZTtrZwUwKHOgyFxaoxRGeSLOdATcY6NfY760Roil72iN9Ife2FFlckuJLNqdvJ
h56tV43kLlGKZky/8JbFt/7gbFmx7DWCUyqJWRfoulo3YCj/gHtMEOocJqvcEPkF
Q/VlttfK3Gxu1eJ0A+3neh8QnBBSQsOZyWaObgS5/7B2ujja3NA5LdOvfL4iIfLE
73nSFM/c1stfuaT2GzG61qVzB8AMG49r2WleVjeGOx3MwspuLtT67Wz2uplXn5Sf
RosgtwlAm550BcDY7jXQZLc6vmOUJfD6NfQNPMIWyOZQydA/I6BG/L97eDn2CAT5
Nt8mzM562uSdr10Eyjs96SJpakDwtEnYhtn6rPoZvWHQM9I4Cc+W2CmqnRinZ1js
CSM+iuZNmws+lbCA56fllNRJv1ttmsuszGHfaI/4dyCYIQurXjxijT7LY0Rrn/xe
dShsap8jZRkkWEzPdbuso2qREGE3oNZdGBRXjWOiC5NGy3rVO0zsxQbBx0eftofF
unOastvcqjyC0uhxc8iNrnUb1d+LQnWGWyYItMzZv+9Vh8WNo7KI7Fusz6Xm0fUT
DGF6digRE4zJKLDDJ3ZHwcjknLsnDlMqxB0MOTfwByaHmNItSd6O7wvQ89tU6zjf
eoS+Uf/K4Ta5fHfUj7mIY8mk0MwTpJPDbFD91EHJDedsDsDU43ywegLgot63Fa2h
W+S2Awg6vdOoCXanHyv92E/5oO1g9l9/WKJTXEXf0a9n1At3RWfpFMCGMIv8SMAu
M3/gor+bW0plzPIVXyaB2pGRXKHgSGdbcolxzUFektBDEXZwF5MIQV7eFsd+kk/l
KAQAY/G5ZjVChaerIFJG6U1Ae/P6ubzx9oe2BYnE1Vi6jUrLEKFw2nwKfjCAPOiS
yqEsPoymDJI4fwBZc1JR02UsN7kXsFfiVFxuYverUSd1eSXY1+la+eG1+6VXmN9i
ImXjhX/SGXB64ZRqYI9kHjiRQTh0UioTb6XWADp0QQd5tsNGw0cT/TX1mpuPm1ec
PfR5dd5ICJLwKXHh0E4nhoAnxqzFh51GdZV7rbwU3ksRicIoX12hUNwFpxzsnsRY
crkI+LAENRSk1g0mUh80azFNlovNlhYY4KlBWeC9BRBWLlv4LvK91MrJtVISPy1s
TeMxHmGyk8lD9DKLnnYEU9zHNHT+SUcCE+LKZLGrG/yjfX4CjH1aVn/VSBJyplyz
elSFAZZ+EgSu0O+5Itf2EI48EiMH29KRwuoZd9RAo/03tJwjgxCvlf+kV0t36z75
KJeXpKF+IRGU3gBacDFSmZouJko+hLLxRdiRX4EFu2eI5zrvdQjVvezTNPUCeqTr
kOR6o4mAWeH6QxAHrlmAMDN7rvg+v+/w6zwCxSb/jTu4hyogOaZgk1094cHRWR9l
1tZK7ytTyLx4A5xLaO9KNtjukAFo3p0d//yC2hGYQKnFpqCeIdXNasGCG0Z8kSun
n8nlV8Hv+KAKcuPwRSkySdqHyqtA7wRG0YuiupFEpQK9whJZVn6la/XT4F3qnUvv
/dXkLilXqkiWtq0idJtpfHxk9E7N+/GCVMYgpANpRclEJXkGdv52vNTOWvxFQJaI
CQEeznKw3tp0nWnJXGplvtDeeZ2wXFGu/Y9pXpKDtqqBqYGkKGYxLy+xk1nmCh0O
S33UNccb/AZ9sj5BHoTXKvXFu3UmpMsy1tsozR0Shw86HODSbQhOOQYYvBZvgC9z
wJamTGVWsUniwxRi4Udv1tll/crF2b/fk30jUyb5F/AAZpTAvU9O1qoJ49snSeX9
c+Av6DielUSrVM19wRSkrBjZ7QfI4M4cuuKw5FSYCw4EdOK5v9xLKu95ZCTwaz+p
2qzBP/c3DZ1bKlT9SiaKHVUS04T8RtD+8YgUTap0tb65oTsZ886bJxdfm0aE3tKx
rkXaWUvf1gzlfK4lE6SgxkCqHkMLbdJpxBdiWKnmJlNOu+t01U1jWzczgIfKCOGd
7vwnwg8pA5C742I+r4MkSAJgBTp0UGz1GmFEz7QZDUxupPIsEyJ36i5572GW7N9j
DoVJNq1wuFVG6nLKfyeqQv9BS7ygI/FIkXzYYeX3iD/K8lkuVvMYIqy49Qi5UQZ5
9NaTVnh7nh0IhO5nUzeX+HlwKjcSowxz2iFaHzIYahwKT5EVxXlQ+APpUyudxGXv
0YA9tXks7cDZBANfbhHmvhF/Xu9Gc6RPq2ZKPCBVafYeb3L7ucBuv3+8JqnXAKDR
kGrKYunOCU1cWZKu02Pl4uvhVhhgw2N/AkC9m3HSMreMjJduJhqvvzQ3MutazzBc
KcHhb2SQT0dfjEunl6jR+x4IAWUkB8hyj8pUz5BOChuxkHjFF2HobsameBEUvaZU
XyXafGC8bZmmg3LkHCad8Ztvi68E3JM5jrductx/PUb+VXO1vTO5GJctvEs67e9x
W7GM9uZEseOqB1jwD06jOSHxOdQjLDhtFnolTlDNm5JR9v/yaRpdWsgulf5TCl2+
XV99so2MMEQqfDuO/slb2SvbYhX9wsnnYdvZaDVltqeuKz635Ipj8J4f6JGq5/It
mBlbrfuZT5PbWfuA4P/bP/90ikxIwaULrTtxhz2gl916FJLCpWemWfb3Tbo+4amB
J/SN5Qs1e0M+5ibhaMj24Af3cMUckkeRlQi2VrnAl4K2Snw3FhDBhP4gWW1tArd0
cBVAfTe70NBRU7kVberjznhQaYRkN7JcdbT5y0yEzygs+kexR9OdSQN6nV8VNuUw
CI44MV9KiBf2NWdcWrmR7ouSxPurInqzBSKLNIkPlsp5u7CRwkXqSoCNaYsqox6v
veqizI2DAaKgTvFyUD9UMAi99oqlY/4SoPMu9Z5q4/D9fpKyvy+nIgH29oonSChq
ZQz3XWktUqVSAn3pSeZOtuTjtqyR7x8uuKG/60gRV/+gR8XS80ijJ4Dxe/n4zrQM
TQQnxPrPffDDum+xa/JcVhZJbI02Ex+gKpZckjy/yiXRzVyQfWFBz1oZPgrkrstC
+edxa9wrqQ7NZsAevoAhycEae2uz61k+A50jTKqbIrBcXQiFqq7zzUCROV1UlNBO
h2FNyen1ab8S/f//KFAsGkkldfol/op9Oa5LLxvcRSRaSllJBEulsLR9KkEMP8Ez
ztbzqsQ0G+JViu0fjcc/+IjeJNG5W46K4PlgtXxM2WlQLRwKkl5o8OYAEWwimwC6
0/Iq1weoNRY4kIDR8ZL0eOUXvU/mOCnjduMNR6N9azSoNjAlRQTAisai/mHQHyoB
fYplra3GW5U0PJLfBGCBYb/EQ3y6RHChfhk+tiIViKBpG7MTIVg+YbMmBdZPsz+o
XImyhfnuqJ7SqIrsWNA9vXYHoHpqw5sOMa3lAJLSiDXFzaozQgeyjonAQ3X0eoQ+
HULIlw+47GHFBMhQ+MxMSWU0ylBnC0qAU8nWT4q/El/pBGDCKK6W4ouYFNS//NED
24q5Qnj7OcxyQGTqoSZzaifRYgH7DPRAkFPDUo5DYDqqKEDaLel+mxEsaJh8FiXB
v+ZiC5eHF3qP/3dLEu9LiqA3uME+UeSf9gQ0IyaSEMx9eET4CefmA7iNRgTh3sT7
eqt/1GAr/uVbS3PlWMonlA2FmqpM5Y+n7rj89NMj/mmHk1j1xaoOsNDsZoxkphMG
fgOwKhE4FZlsyBLEMKffZoTMsPv4JVV2ArvLaKSDzd3S7avQiySB86f02mNv2HaE
jfPI06BVo46w/b7F04JVDAqo5qQ7jI1I+UZUN3rf06BsQ42mLzUkt5onnJRAUso3
h3g7gOpMGHSfArT1GpiwPhaqhVILj9F/Ho/FTNSuN4DTWk9bR6b4YaEqK5mQSXMn
1Pz6GtoWxE4HvMWAtpLSNbS01555G34INej8zcBCYhs07CFDHiShQBbnTZmGDG2C
rWE8latp6IOMhRyCGz8fO7xKQOFe12kKfj6iRJwMCH847kZOVrqKnTQakBNNzjje
WxJzZKuriIdFlATwrGxUYY1avd8P628OeUwc4/vcB8mxPT8XUYHZCwIpeLbevDnQ
Ob307WNEQ/TpjcRAl2uspdi3aatep+lHSoq3zLC/ngUCt913SwChgLBV+NoOqCW/
7VD0Ufa0KLDL7af+xNUT7+dbMr+1qIy3rgOn8QY0uXN3QORUwe8uze1kmPJ3aByg
vZuz0sb7e42kO6UozuXffOrMBICTgSYJFxXRHKgivF3e+IypUwkpwCof0cOn5Rm/
zZ567NDq+y7kE8vQ6LWE5RxSecHptStnXsvnI8++3tFmgO4/btQLYfLb/sHAOtil
4VGJ3pM185w8iGBIFCeo0hA0SDiUZLHzXLo9mBYPuwdAP7hhhD6jooiYqkFLMsvo
hduLw2o+vqepPuIQ6Tm4/Pz7HnG3qJ5enk0X0WlUPL6K2Ns282y2g7mCLCddcxak
yiuGyqLs1sGu8oA3SERiLFgoanDsgTytq7C1bk5UhNFmnk/Bo98mTdxTHtebf2+Z
pJ+PykUWwzrqi1Jq0Y+bYT0JcNPtbo+4juqIX3b6L7D1TS/NvLjlDxzTO55gSf6R
2rlr2c0FNK8cS7RCo6jGKSCOytompqFUg2JT+ydUtdUto9pJBv+GJ4PHRZ75g+Qu
fu3kHuTHYU/N52nvjCgtEZuTICYxkDwlo6Y67e1SPsPyG64vFK1+fING2YSZ7HYS
IpGqQzerp8OFeJJ3AfG5Md6BbK5xNq6vqumWtVqUuxx1tMn7ILed7bBOnrpexgiy
a4Wyvdb9rnC7RhoGfa0hhIw1fCxZ75nggRrWKNBHNrlzj5+3nEtJ7tVqbw1Butui
N1YqaO2R80hfuhhTdg1aY4TY4iKyU+JJFxo2rwxpSViaRRJX7q5SHHDaii/BzKPS
Xzb2Sqxmj6tdeblal8NEzweUO3Nmb9XzJeHgohaMLuA4i3Kz2YyfRZGxFkbB6QGV
JwG9ku4GPEukDRtEJGaWQRy79CFS0zjo67h0gifnQej4PW5nIDOboqDsrocHfTOy
OvEcoOujmUj5V0a1R6pZRHhhsfp/sjJYVDtoqoRWmG0BuqOWKYfHZR8EaRLC+XUk
Ep0vAOvsaKQoRFKl4k1qQH9QWhNVWqMFmTWmqy9EWqxM0ITt7OjyOjuZAvFf8elt
9TiPhzOfLX/5FbTUXvIhElyo6E994hIKlVg+YzQbuwbmu/VcmYaGiLoDiDBdX9NZ
vD5Gi2DqIIG36kcQ6QmTyWZ8OKP9Tu8hUHIOrwaGX5DLCnGVwlDZfKf8sqt+P69X
2y3wKCureAv+Owgkb5K2pYB5GBQ9M0NVUolJhNj6+yh1k3TNBpUR9u08VeEk87RA
GBhX8C2N3lnU7zZjYLKXga/898tyeWtWsUgIdwkRrBsyBxDHEGDttJsqFo6IarlD
Dlc/4uS1UvQ7sewj0guqkry2WSZunpbMmuIfZV56vYEst4zcbB1aiPjRFhyEdRDa
K3qscO3IjlaD8XJFvmJW3WlNous7dCxtJd798Flh9Shl5dTjVGLGS0eL3YKy8cQQ
fSTjBMZJK/c5fSu5BBSxMerl2U3GQkgkOTnH5l3pvIbQ43VsY1C0QafmL8wrnt9U
8K3bBCZAQlPHPDX8Ny3YvQKZyKHFojK36E/EOBD+EfuEZh5J0K0WfSqcFjE8eNWc
bJ7T1APoL5496i/VMY84bs2IpnQyY8+BmYRKvAj/dD7Nw36odTUep6+xq7o3Yjp7
UuHIk7qS5oSe8pR8Z/itNrBaNM2mzeXCOxdd0xWEXdYl92UrsKGcSxrHeLDhLuLC
prGFvq+Y7qAEnXJxPuFTq4GLZLWytYlDxjmKbHxLpftQMuZtQhF4q8hYVYcOCmTT
XsVM9Y8nyd+fFT0+F2gT5Yx9Uenyq8LTN5n/ajAp1oG/4o+6r3tEzsQ/HGayvC3+
wv2wMXHxJ3Ws/cFKzsaTIvs+Knvtj0agdQqnVGZhIua6mexP5CVG/Fir8UDdzAcN
ijYb06PNZe14zDx0U7l8+qTJLsfZSbwutxHFuDPwwKdgzMYtKbZJT/egg5sF1TqK
q1y1P+kYIyzGkMUgm/1OpQ2SQg8ubekrM+NCDObDmbZcKCdBaWECYxUBsp/Q5LVX
yCReZ8QdMShEVRZyXARR9rlVBlUlOUoCvxX1Bazum21Mmmqwklu7vuPLG4ln0OlH
wvGg/JpdvZuQTs7fiwtspIu6K9KSvWnpunv0jevaA4snu7ZrlBO7vsE8E0jnL9mv
mrOesMprRliCXOcTxrw/KUchlDB3EosdgbwQpx+OST5UJ/JZ0wmLSKKdeLUbGxmu
cw7QLFggtj2WVvVWwmYEaeCUjzlNEMYZOQqaaP56hMvqXpM1WpcbcSJ8bUb4QL0b
qVU4bQvZzSeMmyrZRcw6KbpTosUO5aqQYc8c9skqP+NHrIYgm77CmGputCcuzVAI
9FrLajSYbyHca6w3rWZ6WI+LuxBCPJcLEjjRptAsV87qE3eXxJfgniBxzi1edljr
Km+qqbuQQi10bzO8qdxA6U8SP2uF0u+B80U+fJO9dXIyk0oJbQ6e3fvkQpoABGAF
dYgBa5oSSZJyNTQ6D7DxDdGP/uTh5/vPTKGVfpDpkIp3me46CAFjN0f71wpp/1va
zY6wYcMr5hnEifCimkB0n8pV1+thNkqYOtQHe6mFc6x3cA6L/09FPbhmzkGmRMfH
FjkDcl1LvZhiwCrXUo64noKclsG//CITiXD4igMo9IZuMqi/zPp7hUfI4g1AvM6c
KQc9Jy3ytGOLp8KdK8WmiTVrt0jgbgDF7Q9QJi79E8V3Hy7HYfUeXe9vDYOyW73Y
rRbGaWsV/w4XMpCr5HB8UjNkvkVhHMubIunaHCu8GgbJciy27eYehBlcv8ew7UiC
/HNl81WNcRHdwPZiFLrUWmaLMZPIcSaFcTkAaEaxENH2hcfu+LRCFcWBh79UtmlB
1Xf0ze85Yd0yUcGCRFNX9+Yc8bd91+D2mHIAHy1JPwAWbq0xcAWWm5WelsoyOWmR
TLn6yeBoKP6/HotjW2/Uk904EZ09DjoaC0UVtuNLKNxdMAVCcYhsqJhxQfTv95lc
3pkq85cLocjtA9cIuIypxk/Cxo1tC+zQq7ECXnMPZgI+9WaFVgnvyR5nFI6R+9FG
DagcQ/RfF4oKef5yMgegeNrw/hGJYW+jU0vEiBd73iNw9TivX31d9L2jacQasiHD
krhfQyjXFi6E1HwReqLG2NbRFaDG0QOcPCAcIOk8UDW/MfqXic495heBXqnpA+dB
iUfLOxYsdVdQ64fmlkRlBDdm0rpYgSkpD0vxaSv+DZOnpbl4BPswVh6MWvy3mb5c
U9ALzEcGrFMsR/KrdwZjkhLniWhKMfjRWvO5btM8tzpA16/yAPPHRwWr7yGIRBl1
E6jISJTWLL4CMqmahpHsu6pWzEumgfGBN1M4aZsX71EfmFF/UnUORBSwfFh/XAcz
PtRZo4nyiqn7TSI1WMuDuG3dyFcXlN4Z4B8j7U99caSXdkpzNEsCACQPCK6ir0gM
5LVP6380XgTn4yfplKQcHy8wHs7ep18wqoY3vuRnYBXtEokbPAlnZPGGP/xwPRA9
48QwQXfX4dWdPSY9lnEFgNGDQ4n4fWt2HxLbvpLrJSSPnFTMYQb8XvQa3WHVl4xV
pMDrG8xWfl53YwZwJri2kwHM7LJSJmR/Rr6KO+z3aqshTdAfGfM6axBXZmhLo+pn
MLP+6SPXUnfPduSI1DhiCoKx2E3SWiLecANrckwRJ5lo9MxF/wQzdLHcaEO0ctsL
GRlZoJMdbCl/DnYxz2WUFdv2RYX2akE+9OD7rk1wtpfYZ4FA8JY/lNkadpAdam68
lbX/38TkZ7BCCqN4igiYVHMf/MBMsnOAUdk385dTlZ8/6N/NZ2fgMH7td+B7s1bm
A40jvsGWuX95U52DgisTc84gJY2MiDfrAjCKybCqM4quDD2AkbRZ23QHIisAB/JX
fYG6Co2aGa74CX0Gwrqs5gaJBrdYUhms/m+hIh96Lffbb3atJj6Eq7O0DuNPglcJ
srj09fuf3+sV0d3ViSef5qpxFw1SFl/OvJxS0Bh8FqkcaiGYtMDBOYNvaBGQd1hi
1d0n1iXvAXwIkNr/ygx0IvPmU44Hyox368mbk4pMsO2GWP6DA/fFxb/WZrnWF7es
gDaxORUW3hfPadrI0keysPvdrdwpgG9cvWNxRuQsrUF7Cpl/eRbPXbVm7ksd8uSj
BrpxB7tp0qnCr/MrdsJDzJCnyr30BiIlyw/7Gn085gyZfxiL4CRYSSGl4JPMy9US
rec/finPwiKBWo1PJXbSph2CSTN2HG8ewpgVMHgZzItgXZg/jEit47xVsVku1O6D
SzIIlQLGL/4QYqx9qD8dj+283/diVMGRaCx2P7tulZMBv1VVpX/NN0lu3VIUOulj
8RraUtn5gVlH/wsj//FCX1YpwAkDTLlaxHV5iA2PpTWgBBSemSAT3Ux7Cy+f5LvU
+oAIYVnuk7HSPD5PSJtZlhlk1BpCBjQ1olJINegbgqbPKy31XzmrXmO/UtXj+IeN
GzLAN2FXaSgOX3uaTzqJInsqbZ5VOOwuLuEmCwJQYbYBHxg/nUN4YansVl0OJUi8
+YJt1Dy0mw22QFJHk0MqYP5m6WeaR25BE2vVzKhvumnD3t6IsjOev8HUKa96VzJ9
lisftTw9gRMC+ThCmY4EnBVfwnTK4yFeA4hUlhkxzX5MueGjaswjZG8vXtOYVnUi
FU7nkPk5a8y86ZMEC5dxb58Y9OjxTdkYEXnUzUim8ILMXAOt3aoYCAGeuQfhqKdr
9T/TyzZf/k1cr89Dxg6wuKiw6VpdxKSHB4sCherOV9MYp8opc7A/BQaHJdgoo4WT
qRwINJLzvhRamDiMf9mPesx44f3eNRwmftOQrNlfEsaQKnezDZU6musGw16xiZ66
mSl2VdoLev6I68wLQzi8TbvjkxZn7JLQFn4WRG9nQcnqUu9DEeCTEg2qJFfxY3v8
nc+Q1klsbXRxWBPOTLNi4FWJYhAT5eBatA4TT1Jc7qDcWJMNRWT9H+30/UC89AmV
a+SLxxmRNHEqG4GWhL3r6GRzjckjgyClzku8ddtwYnSjU9809HaUUytbKmSD1vnb
T8h/Y5C5c1thGpTGqYX2j4wKTYSmylwi/xJfk5iUIj8zEIGspWYwz2KE5BtDdY55
g7vUnZSCVvWe4E0ulLd6vZyTH3QsqSWQ8woRBINRJK8t6jlmykRU88bkROAJdKiY
t73cWTI38Sa5TieIH55jtqoNUOV1zjQecrGt3VfKuZ7GZhToAzjIkZrWSiMVCxY5
j+r+3P5C2hXiaTJL2wdgzCeeXTv43DxSf1gu4Ivs2CD2dpRKss6xaGaDntrrvDBB
SC6ve8PAul0To8NbCTDpb9bLx/zyxH3985s7Ux5UbIMbRXq3ahl+ubi9bPAFkF/K
3PsTlBUxgC4ZDH8am+HsLU2XJV+iva6q2WcMrX99spFwPPm++54kb51E7fGlSkVk
g60vJ0UdLvt3qkFUFD+Jdn5dlDxkPEZjouH5wTffO7lEIL/55CR6VJEck96s2/ZO
tj/qTyNdq73SSfIplILq0kMc0dZncAuWJc4i+vaMAAA46U7BYp9LOxsGtB9vq6X2
akNbyp4ZBJ5HBkcE1cTZlwrG5zwuKPbW0ldxfbOrf/Fk65vN65mrxqtIqHKZP0jI
GdKBSD9lmC3ulQPHDX9RwmRZ1ZAsDBtP5XEjayoGYYRsSuefpBpE1fOmzOcFWqSq
0gsjPWbJSFsmuZyyhG/sZfANiZR3BSqz0sAITaEEKBZePf4CzX+mY5BmBnvwm9cU
CzYMD1zgXCAChFxHWVja2CT5vGa36dSjMraK8PUScr703BxUXiBJPgTSe5jAnurt
hLVuddfHMl8cZN1uAsCwQzxQ+hQ7rsXfRjwDPrLkXgWxJ/V2bZpQDRjzRQeuCpMm
jhTJFJkmo5spr+FBWcbpEufprOkx8hQ+CotyZiaEd3G7MfGbi5lCQX9P5d4OlfFq
jmu4uaKa0sdimd39jPFdeUQ1iatl+QQKZtMFgxKH1GM8TyZ/AtMGzhQ47EWh0q9e
bivCMxZ4EPBV6TU//ybK2vX38217/zhwKZA93kyf84EEKiCJpzyL/2uITinx0CpW
sMDu0nN1zYiz01BfAMoh737Bo5B4Y1g+lF5mKm5NqNUWXbIgq92g0RkpvdYKCbrz
gXtmeSdkfFvarBo0uh70NVC21akYJ6KKhBV7Ad8ncVDgTY/kl+jzKTjxxU6+1ws8
vQ63YEU0xTwg5bzbPA0d6U+uSmGw3V/nyhuHLfUWdvOOvavrYU+2cpBnR/UKga5H
A8rAn8JLstZEF2LbSmK8BcxWOB8qG+m8dMWgBuM48UWxgMc73BwoCqfqHbGhCwQE
ibiYrBksjtO2N8eWxzd9uHJOdLq6k/XQBh743x8644lp0w5da0luiGIjhQuopqi+
POUS6qtHpL++tdnZZdzUBCr/KfckxL8SlSng5d8SDC8d1uh1l49a8JVm4DfJMGJQ
B8edWSjg/EfiW6a3phD+Q0Oqbd9CtyoZJYWytqCcqDurZg5BOaTgQIobmJwwfuMi
xnSAwXglr4CIunZ6YrDf1Z9ZVNvYWl4gZTGX5Rce4LxJn/+98zf+YEYL1CytcMlg
PZo/xRClUhjSZDi9cUbirYQPRJVFak0pdXXlJTnN8DDIaKHNVtB7LaOpgeCMSA3D
Cr2HQGCr64ttiKCfVOg4sflJSO6gjwvM8LwLqlc+wNu3N3aaP7x4ju6ZH4y3MSUd
B9qxL4DFolj8eXqGFiWNWhkNVrgqt2mgj7UB/wRfopy+tYhVTZ9qQ3VS7XY5/hD6
ktvwYAIOhhwygluzl3ygeVrqAdF0CLknKsW2aejH/8pRgTu0bYoRom/Qq7B6Bubu
Cb+bQY6UCt9KZuaI6caAYohgFKLAzGIhcBlm2y0WI4S6xFzG+nkP/wJLSu1+oXR8
88xDGXbwjZgfgaV3isXAIcJJg32vmwDIATnPFlnZIqilL0VhsvPz0gkJ07LDCwlJ
ImE62kAQHIPaEAh6x5NrrviIwJ6SgmFvqmR32ADqg7gFLciKdq+DcIwza2uq5KoG
KFnRkVTmZseIgdjJwGFZA74seJReGkYvD2EgoAirPLUe7hX7un3LUWLB5jSWDNpP
FxqRVYO+CZ+0M8eNa56QwzSUbu1zoGYc6Y1FABtznc+jJDzazb5g4dUCDFLInUz1
Gw/ok2pOnyCXAE0ApbvrNlS44nqzvFnasm62u/fsOyq4Jxrv7CXjDd3q+FqQuKW9
uyoL/QW9d8jpd5nYrR3y0ylsh3F8zhGmmRUyHmXi/O+NPZ+3EK5txLoqNISQ8ZlE
QvYIPDTvXwqziiyV663h3O5vvA6Z94YRQMPG1ZMYx2GmAq5GqLvz2o5Ln1ILLRDL
+84ZTbH77yFmQjLrolWekk7qYVB0Wy13W3CCS/b/vIfEp9mdWLrxj6StRJMn1BaD
PLHGJ3atAu49+St5KXYsssM9eJ+3NoeGIEZQj9lSO2cKBKwbSl/aB3/UNgZ4kFCq
58AOXVkqsU2ZaxAJePlI9O8p23W7cSNrQS0bfiLN4gdDmII/2j3OQtuk6/yDa/Gf
Kg7zo/9KuLd7S+Jv1Z3C3C2JoCCKexvE8/NULnZPucNvPjCu5kAuPEw/pUWAKRSP
pCuxdCFArOnXbtZNJPoiQuOSiYp5aT2tn25KRgD06DJLtkPQMF3x9914ZwcpSm6x
5SwPZN6vPlM9V2ZIC8SREpTADn39jASXTJ9Jd0PK4uVJOhMuKRr+OECkh0kCS7cj
WpQyJA0WeNyBMMbebd5UO68FJmZWI1evE1P5NDBGCofUySi/2Cz/FPgE+D8DvFQW
v/2O+Uj/PVWh6E1VnS8iRt4C0zNjhBv2Lp/Esso45lYGhWfSXY4sSyGBrOIS3a52
a9rJtMdAuy9cnblKIg7zlQJn2xGGedW8Ux9oKCLqP494HbueYCubutN0JUExrxOZ
15/LHRhF0OGd1KaKxCBsXh/E5Ett3/nHmDZDjjmEeIOnOcKaI2ODNr7sUC6Fm3qX
Nxyc6N7hHRPJSvYDNmrtUzhgKUaBsH3KoCBFz7WSq3kp53CsH3hjdtmhPowgcNin
REkTSG7k415zAQ1EJi+j4NE5lyBq49SDv1wm4KdRlyVjz/knkWLfBD+mDwDNI6i5
Wj6oT0XASChlrkRE29Nn2G7+dKlASowXPBaYE3YR04P7Gf4LwjOFJuV/oS/Xshym
Y6xsCo0nCJ811vyLzGfs/nllVT5zvpyhbGS9nQHkhGbvIHMD4Zo5yukb+VaEPt6B
d2GUhan4ORiy2570YSm53WNCm/8WHmoAxMZw0qINjo1LHXlBpRuWUQ7guRFXc5l/
/bg0PwUy50lTrrCVwQwqy8HXsShjQO9IdBaK6OAtt0V9n9XwxSdk+H/UUhMpSN3S
b5iIvzxCurYXipCJCGYwv8xZZLpVi+eZ2d2VM0mzHjDwZ6hAd16tBLaeq+p/Ik38
gUZyNM9LNbvqw30IQJDVr3Y3WcGnwx12tfbv4cStk5NDVosOMTjP/TSdsF/9UyUa
Xn44bW1+/kn93kbvg87ba71MJl9QQih8RxnC4DWnISc/quwhRVCkGFBXonLC8hHy
L/tWea1j527WbOgFpgsslLL0NlLs/cCSEas4k8dYxs9fEtFxByYhcsGZLRbbhGyL
Vznw19qRPwKD9E7ZlJ16IuXw4uFjsRlavND9ZcPQ9FzXHGWyrMAvAcdl4OYCd+Av
pXJfOQ+Lb1IWARWifSzgdFuj3KvujzfcP1T0WZKWdFigx8Wq+J9Y6QIREYYYrIT5
7viGmimhOS2UP3ohdEfF0VBQ6u1/qymhFcfF2gsbNXlEEXO/dAUMeOpDU42LIB+o
SIvAN5LeD3rK9zWGhaxN/gwAmY2H8ZIAepGFNW6YZ1F7QshjG3k0CdrHIbg9/ovx
lYcGXfXRKa6HGhiwi+N0uminXdLz5e0t7jGcg/CbdQUNwnWvjnqK7PzkYaAXp9NA
k6gpwyHMaEFs/utbD0o3euAAIEIBCmCux7RVTbYq0+FdTnD887U/6swGnjQUorMZ
ArRL2+CBA+/dtJrK6hRI4m8Z6zRAOPsdQqjVlfr5fIX9gHLlHzvFYqD7BkeALl9Y
TPSOr2jzNEnjSQFNcaV/rp0buN2t4hpNQNgz95kqcgFb7zKJgPF+k1G5UhETRibi
6Kf260F1G7jeOtRmIpuVS1zMvna5npDxdkbF0ofodZIXDe7Z6Y3LulOQk4NeL/um
2orMsPC+eb7YUD+0ZUfp2Z4yfFZBJatbcOktdo3JYNFxA2A6MyeJlEXCiGzwyME8
liI+cUTUnr147zyArF6TKWvUD/J3nW9x9SUNrHqsyx+vP/gqgSATIrUbkx6hZbf2
lSA3t9kF4W2/nuvuf9mMEE1SrSicXHm9uwU8bTjwOHDXiYWUMKYBAbJsZPNshOni
oCJEz0UwzA78NDx+uIFhlzw9bqG6s88jH0AHoynIwFynaDaYss5xfQJiA4sFen3k
T7KtUJxxOSrEp2kVXoRU/5HH+oJfrt3hV6IjdWUOENqRwCE1ePHMsIBlLknkOkhX
JBq7wC2MmV4Sfoupwhkib/plNEMvpEMfVqc0GPazFV364CMbHpyk63LIFVYJOd4w
uSFQVyRLH2I4fVwpIHTIlSmno4tkupr4bdox6UI+0U7s/TUzURUtIoK6dcqf6Nnh
dYUSLgxnhaze6JmSLXpfjbMzDrSBB1TTt8BQNWjtxtfsz9hqnRfJFBH+qqv/wySe
k1HyvdsKQ9pEOrkigtN97hzi23zBm0KdFGLKVpURhB+gm2QvnTz/jkzD2Q6rz/mj
wIgh53TOBX0+pRj8DRy0odbaqvZPg6H9KgLUsQvuPegohJKZR4NQcuJCSf3BC2bZ
FzLBmv6doN5YPSvuhWxXB9211to6nz+DKhjnOmkva0YWuNBXok6vtf2diBRutvV+
4FiW9sNd8wPi5Dy88SmRSVQ6qw895WbKNZr0p0+uQXObDGMbFy7xoiUj2zPNsLOA
ZcXZeqefVhxf0tnUWb+nSM0SGC5/JIaB3iT4w7HUacMGyRmJlHjW6qhCq6RDFfK9
WijV1WMCVQVTuX9lqrguNAnNZJXjSbNminUxa68pb5jOhdllz1hEYeFNFEC48YA7
JD4d9JKcmJZrCj0Shx0kc6xetvvJtelRFinQma/SXzKZQOFyHNdYBkqSjXHLZYZu
Zi86PRw+Bui6lgRtBxZ5j/ZHR4/EySLBiqzPb8YmwsfruyMk98zSXZFTvmhqxsqC
fMEt6ZGbPgACWu//VZve+3zHIaBGWkNJP4xwLp+pdQA48jb3nzj7hPQ4lXsJJpRq
K/QzK05n62qnq9H8VtS9K/qOWEwA3D49kxG2vvkrbLgt9YELGKPjHIymo47B8j6X
kcicwayAj7qo4DRVvjm+sd3oMqjNI4ZLc5qedkLqqeMFEliMadO/o30Eg1yWDKdM
5tkH8E7OT1mXnsyhxDYNUO/tT+DZw+HkVRKulxs10CODWW/HQ6LJ5RIEcOp/CwSO
qpMY1O3Uw40Z7OywVMPxUQKo49nj/MckVzhc8v0UpkwtEuEtzLyJUIofoFC+waZv
9lqWqBQbQG3mXw9S4nLkXVIWRVQyCSiD8rOKD8kqWYfxSRdY2mHnoyFByJEs+RNL
kGaw09B/4bce8U10wvH7XtHhUSpLy48xJuDHhFC5T3LR4myFJbQ+IrLMU3tFxFZQ
1+Lf/9M3ISVqBPnHXgxIZSMPYN2Yd5SCzqFX5K3vGkzELK7UbaQ8gLBfuOnJo1Ey
Ds3QXAUKLn1hhIe1fRPYDKx7ZukqDZZtGwJo0xgiNsiuWhHsjg9hKr2vg2Ip2Xxf
orVFhm7V2hhq1oIJXwT91Pbkf1a0bVt2Dj1o/uQmC9x/rDSirF8byw9zsAZelmQ1
CEci7hASFzaP1vxDqyfuyiFV6sZ6Kf/c/+ORA4zgEKlVcQoiuVpqLHwyOkrzT6N1
zUGwy0wONssxdEV7iVC5RyfqiCVW52v6u0yfMCtp7I/8p4ARLxcz6zp+aQ1684wx
qbnT4bFsZ0mNDjjayYsRw5sRfoctafzz07aVJtD9ksFTrZdWBYoMSACqlcYqBq4K
jxi4VeGHXQVRiSnHusvkVTcFnmUXGvyniBhF6AVmZ8Yz/fqxTwmvPTRra48hdCxd
FcGTmte/gM3bDVU+Ds6vTTqFQnh9T49yeYX0zbYhcExwSKwa/Kq1VzXjWgxXNpQm
3xGNobBw+qautJ9lzWCIaLNN6Cfy0J55/s7HNGBwuGWJHnDm/qNHb0IoFC4RCgPb
vbGz6PZFLYocEJDdiSdiklwQXIbRkYGQTn/TutaAIRWMRTHy9+lUgEvSqrAEzSdQ
qMwepNFzAYcyE4KWGDxVVf9xLq4dRcX3uACx3Z8FGxrcE5xC4FCXxxhd4i3CAlwQ
R1H0xQX7yR35Nyob9DiOjpn+csgQN7NKBGEXgyL9YnuuILR0KGB7K4yk+zhguehD
xC1nmDxjfmajdRPLqTMn9zSEYE3bIhcNKTCY+sy3ansjD2dLPt3ZVDDDTsDSs12R
D9Ggk5dUcVpM1XcXtEF7YdZNw/zL/lFTYlWq0CLWkQ4j2Ras5lovLa0keoAFay3j
n+13QGR43EmBrHjL/+C0rHuUnIuQuJDFuTYqIebwEK7SPF7fqB9StH4oAsYKiMs0
EnwTBMVpODcEoU+W8YmD0FEAY2lk64/EASsHQRte1O1/zOpXp7Il2c3o+UZNLr5N
YLmT6WV8UADizlwpNNeglVOASxiJNvAVaWHHCjJW3pFGf2oIharbf46wU7T3WcNo
0/JRUw5oZbwdco6k5iakySvN3jZ+rbTKbcF7TnMvSO5RNYgWkIgOrite+bRryi7h
95ZNLirOqw473b8HQkygYZREfxREi9+NbWgkDZIvyWRdBxcPzHZmXCtUAZ8OXMAf
eMcIpINpUtojoRwbrbguM2EdXjJUqLFAeQMj12OoEhgartbv26M6buVwRC+u2cn1
rX2MUti5CpverbyB9RZdLG+qgkU8MRy8O0ljXyjrxR595KzrAXDZ1vYyVvZN5XLk
e+8hs6/i66t+P/QRoRjo88lFq5jgc1PmRSuh9XOX5GoF1HeZSmRB63AlDosZYo9+
FDpT/cmYIPUSkXBnJaSdeG0WNRpjb/HtDk4CiHCcw4K9Eb7f8BtNtcIO5EJPmbEw
Ow/ZqIuXQVLXvVjcPE6cgUImcKJSwJUiww5G9LpyyNaokqG0+2T3LmJsLGttt2qu
ZhXJvVvZ+hN+OfHIfo25iOqWA/vhtjHIaPuw93w8C7PsLz/bRHP60bLsZPL1w8Ao
ijjmQz+NnvrWHisb5uxgHTc9ERhB6CJKp6RPffEqrsPlsdfXkb2qdXacKYJq9GMO
t58gvPdIQL/r1JtQnPrX75KrTqJnATkg7K5tWGIjlMGSji5VSvquG6nL4ag67Afv
yON2DLdBQfU84sLHGQkoZuU9l4TZHijyGKhA9Tan0DhutNnPeZAKQSx4zTsB86Mr
7Vzd5X/8/oDh5RaRSn7DwiW5JnMItdYwwrfNr2cQUzNPmaEb8wczBL/e+ZcvIp+m
IwJCG3Y5CeNPo6QejTf6q6Cd/YHZargGuUHJbnygtXC8MXWuHjvvpF0Do3q3NzwH
H8jRt7XMfc3BISi/W9CIVJ23gNpbyBSs4mv2wjYqfqlDVHCMxQw9UVz0cIUREgxg
WSvhrTCa5DRCFmW4UAlXTWcwSn09KT19AefiQ/6psl0XfCXVevcsJEhGmJbQZR9a
tkGy/KfUNAaLBFkXlN+DP/G1SW9UuAl87Nuivj4yarapkj1WzRkshoxR4G3IGv7u
RwUJbYhHlSMUqowhgVSuCBd+CMUQaohtUhJgZULfBkXSeR/flfK+R8OQoK2BCdke
ybh+yEojUeuz5z0OzL21WynUSEVuZwQ21376ApOk5FSGdd/o2+1xIzY458tsiJFA
UQKDB31Pr8nRl4xsEz+qX+i+Tuxv6X14GC6hyXb8dlFnExGgcKoT+1g01vJKoR7g
RU7TwFUAshrnqj6llbmTucBIRpXqP2JtRL19gVi7LDy1HSoe7D2vRqns7wJDohPr
SBM09UxlaxKD3dC1u8fcCUKAFsN1SCoAetDZcWJksXChRZldshP7PEPi7Q9sNLWX
6IwEIbN7FRLBDeeCF3XTjrRALARlOKnxE3xux767V3+ti26N5RYKNMTmV17mm3Gj
6iI6mXI6fgD4aDM33+C57mSSzUf4lbVR8eXU9ZyI8n7c9VLu1kmP1tqY6m7hgz44
1G1cvnaxC5SoPPp5FULltMclzhtFhbkP8jPVGcwv/tBAbHgLQB06ZRBoDr9PneC/
PHrBao2BOQ6Mh5Y9WfyiupvCCRWomBAwv9oSdLbZlZB9nVs2u57JJXaeKKZ4j7W4
MV1EPqWj08fiV9UI150ftVAxwczIYYqZrBgEnppbXCGyJbBmdlydVCzRL9FLidbs
DwobJzLr7fUBAg4s6Svj0Qi7hV7yzf5Ay5Kxdo4VwdoHZH8aFf233IB+fS2eOlk/
xaXWN6CHHPcAKB6WPMtYJ3YVTtlah3Adqle3EM/8PPpyZqsqjTcVf/DJgYo3insE
J4pzI7C9F8Bti7scHYTzct3zfVI6IvVq2Arh90+S7lK29Oua+o89lYwosCdd6TO1
XfpkyPxICrjjhCGXrIsmzqRcIEJLGQhCbIHDBheKl+A06DhDnbEauZKKt4s0RDx+
go7ho+qCDhI4L+lSy2pDTM/j4n0d3WDfJJy1jxIx++IYZyqmcwlqxvX73MahTCnd
I2AS9RbkSJcNIFl25zEapLhHv8QujlCQg69hgT4PXB5fnNqo+JlNPJnQt+kZ3KfZ
Gp/tNecCHWySkgqnr0fVJhXSwwadal1SuD+xZN8Rd7HiaKtnVDo6DNgGnKfOw1sG
WrMOuqZwuHkaUpTXD2dVCb/uXn8wpDlOPeGRw6A3O/Ri5X3MLII6hhF+iEcVS2nn
FXNrWu2g+wSuhLcCl82g2HSz0hDajIkdEuDOzCLFcpcXOFUUcT6DvbszCkrhkRph
o8qc75/JC99lCFlKLxLiosv01Po95Hfz3g5LZSCbQ1WxLekSa3NuEkGaZUcKrpV8
33aLEbDENsX4P41t691R72ZKa82jfDL5zVzT+RpPSb8R0zDxoWDw8OQG0ZG05ccc
0qtHSc62oeaqbkkLjK8qaPwOLOz4b5BuGbCDWUXgJPn9uRjE2PqLGj6MzmbENnxV
mpdxktsolEUhbbLT/ncBbtJyf30ivQuKCVFVFtEqrdreb6hg6dgdwVqFPXunFn2X
3uTzfzGVeAuxKg4Jnenps8e7oGC0Yi02fNKwUnYMFqL8/yxP7HLWWdmBnlN7Q0Kp
m49WC16ciT9x7VEdMhbmClEhOP+Ii6q+oEeoqHwwcWAYzfp1UdKnbQE4C/aMmpwT
3nn90eyAwgYT6fnsbXJDOAs2jiy5ueWPccNkBUFJiS9wx13yMnYqeoD3JUg3/lAR
Qnwy1ElwKjQnsb5hUAeI/K9bMgPSC74ZcHxqGPb9cktim0KMlY7MX5h7rVNnyCl5
cxa95YGftjbbmkttEUB1t7HTHo49HcbWlZHUFR52OR8M+6dsVafPvMrPEHC35VPS
oegOsZWPYtdpwvrCh0KgrNJ5t/nXDgUF1c9JjJiapIKG/k/6iiuEbdkc0AX6Z1zj
FOAnFPZk06yoXT7/N0rIjUCxdD/OHxhYrCery/AownnihvqJK7P6wWJ25D1+qZPU
jiJM0s3ViMutDdyPrwucd+pnpo+vHPjoM387MnxTEYSlBZwzC7bCt+jn85mLGMAn
GGqbfCiCkPwEB4sYEQ1pC+IZUHhtCIzmxf//krgV+t65/xTPN99jkHL1GfDm7veW
YF/yiYlUQ73y0pYXzQG9h7b421KBCCBC4s5ZU6NDIoSK+WiNpKLhJlAvA5EL3lyA
iTN0e6ye4KAQWKWOMyJNcp6Lk0WZnCnVKpmmh3GYmYaG1/6JWj6Dsiel2ncpmqS1
8slt/fZV/4knHwAK58r94ElqkPfTFQ413uhOC70Ly2fDfUR/7JmdjXhPQSg8zJfK
lNBgAs7LDxqJNkR1xsOGPYbfy8LPjPLysT/YZiLrTMUYxB9KWw46HXH/lOrLAlIA
0qhoHeOVpb36Bc2esdnrtNj4AQx7tmwcm/AwGRoEss1oXZVQmw4D+LlLYF8mlE+Y
Yj+b/kfGfODieF2RwBhdB6Q3ZKmIzjb7NXGLfDEOP8W1Faz53QkrKABPs0o0Z4ES
8xH4EvVX9WVYvPsSPF8Umotnl+90uKQ79woa7LuJbVQTbfCNynMxhlIoCaY1si7u
kjHRcoRHheywTiw0HSa8tiF3gBWxsQB5cwCFt8x7fomtdC7dHTcvTinl6rs7X9Dy
iBUxTN9Rilw8oiQgjfuFh9oy2pOePQW8u9t6TbSA8KaeMZLjztaQ2St1I82f04BU
onwv/oQdFmQZl97G56yYvzf8lPpb5gqGedHsER4mBsCIAPkwqwuU4q+YdWMqP07O
LnW9OBjiWMBhg7W5JChP8qPmruuEkQVkwV2q/pbOeMFN1joZ/sx9Pb3XqclCuDzV
lj33OO1qoG9ujgwnBgDA7LPsfk+KqwJHyYNPySmFZr/l+GuqgQUm5G7nWggjrL+J
9KSXtgdi20N24Dd9QRYVqEtxZwnjHqcQLB6qvdUy4TzY0UoSVWeQenbDGVlOZTxt
u+L6n8noQHgI8kvFGj0+g03YIhkxh6enAuAOg7rCH40QmLUQk0ggJjDnzn5EUTFe
sq9Cs4PLPkAshA9JKCQSYoJm8JE5ay80ddUzQ0WJrq9Xj237DZw7qfTAAH4tmKPw
uV+Z35njwypfRBjlYIiogX2VuRCZj9AvDAcfB4c+bdifOaXnJuCFnhs8b0tt+au/
ipXMkKWw59IWA4sXsMDy8K7TI7Il0yA6ymB+nUBiQPLOHfLDX5p+oZe59l2XpO6g
g68mTb7mbEvG0IpvItGitkX01W9aLsy6VDrJjktdi+/6d0Cnn8KIwhzg5rRiKYlm
q+Q5W2fHrAW1DUaesLduU8iRASLLq6xWoHpJvRBlDkb8QjzimkKO9cJGak7YKCpf
Q9haVDhe6GAcMVajvicup7yWwhhwT8qsjT4Amy8ZxBR8aurjkxz02oVsfuestl7R
lTBaSE6uY8HGvAq5dGkmcvNyIpqq3cd2OIuBBkr3xonBonnvAMXiAVKtXwkwpVSv
/kMHqFj6JDDNoIubFAKjUk3vDWr1E1F3W6X8JiD753bzZk6LQbxUYxwlZ9WGOLeA
pS3rFuPq3Uv9yEONma7ANoQbxaxA101JeuvwK2YHjdJrR8dOHyraBhjQjbrCFP9N
+U1AZ+qFYoMTIai1++7UjKN7B6EXNggYVeK8C0xb2+Sgg+E8MG/qK64W+TLtZop5
6CXS/Fs5IrwF0S9Xx+lnxOo8wylVf29acDOqDAg5MjfvUnhJD3FEE+PdWIuSzHeM
IwEN0k2+E+jsZiAVy1wJ/Yem4h5psJA2Jz60VJoj7BFRbGlcT+tCknqGflqK5cLR
S5W9hrgLsc7K9nvDf5EaE/2sQRFt3Q7UrXwhkCzmwW0tPM7GBr4p4QOIy5nV5bO8
vGyszwJfF3r99NuAg4NJ11XvrrtW5CpNKhbNr9qcRCYaBmPnRj4uK10YlAFI3NKx
UxJvi50q5a6oMqfKW2Fw6dnPpINuGF+s4HEq/2V0bvyBX/ucUwuizTfetH1qy7fi
T4PLSAzsgUXixM8PH5KaNgsrd6pgzngtIIkCLr0EQ5AH+1sFjsziOJaxKnluu87+
`pragma protect end_protected
