// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
izXi5AmlRAdK7eJt7LFsrailjkhzjKRt6YLJmjJpH5pj5QvqtTTKbEcwByMOVfUX
wfp19qqGcrwpmniZOqxRLAAZDWRSjzCeZ1gkK+J9/LCFaJeGkv90rjXk2oGaov5+
1khUuEw8qJ59v3fXdZtil9gEmbnx8u98xa+GP06sFMQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62064)
iPxCl9blfNkYUN3e2UrFdK7ExhvAlrB4RDDM8kl0OEoH0sO126YnIirgjMFL9oG8
n7gSszTMueP2nmo50TONN/cH19yhGHDll2V1Py3ClZhTcOjjqY3HPK8rh6CH+IKs
SzZM2RXuXsTV3YJYi/ag2XieyPJz44O3nkTd7VUP8XXlhXZX8DfPzxj13PjN3E0o
95znymrbIJIMQ8/elws3Z/hwVa9I4zx5Rl8wgLZ4HXJ0VeamNW9cntJqrVX6JvJ9
hC+Uy2Lh8JH9WQ0Ty69ojoiKwVhMLb7cgQ5NyTS6/6hXGTxqbLRVrsmfxgv8wt25
9KUWhgg/d96ZauDyFKRKdPyKWgSClRgS72fqbXhWqjWjy49TQaleIyiEWaIgJ9pY
7UwSYnna3pW6l9D18cBGYmAWFjlEKW0s3IEZ7QVIdBQGcrFcOCDgiWbK2GUi68y3
aKrBJSxy0xP54A1Td/dA/Ha+VxWOB+AXxepYYqw6AkaTMHnfbXzCZdpiQDLLDgYz
SsYieZOUQ3H++1N/4+YJmn1W6amt+YL6KY/M/5QYdCimnFuGC6Px/XJ3AwsehA1T
0GG7dFFTp78RSn1zJtuyjqN0j6zovkBOCdJ/ZN22jEsHjJmiAFceM4eRbYsoV3t8
Usabz4WOqviFfrgmj44CYD/14FBlsMrAnEJb1akjXykjPybbvH+kuprAUHCF+QKG
18FTeO2QLV3mSIhEVGR1bHyXAp1vng7zIMhv0mDMACF5GGIU3Mp3xY1mArYUpCbI
pw3LUZrzNuhpakCXbQKZya+GJV3HMQZYprooqMtydYv1kv5PQ/yv+kE3EP6HtvSf
agcIcazqgzdhmqzh3YOaBpqq7yWX2RARKayy/Tob620VlWmdVWteQHhI9eZUeP+V
NOV5wLYWjqkNk1NVyMb8PChjunYWrAgkm7oGLjWc2jZ6JZfYp8AepuNodYajl1UH
NbonZGvwfrW8xSgfls8BUnSDv8swPGMq10+YYIK7UqN3cgtyZwv6wlRkjCGItaPN
WAN/HfaORtYNtRxQ+9OaLNLHRw0iuLN7GfcYoqXlwRT7o10U+MxuKkRBfzgsR59C
XBs/+VfOEhiPKLzvXB60dVjuMeKr7k9R/Wqtf5iOcZ1d4DWEQahKPBBv++I9OIwh
cQPS/8EF0f1YaRqBpKcTAgEoZs1osfAm6PE0amS+G86yYBRIu+bOuJj57WtKZ7gy
LSsHvOmYMFENG9+bA/nYeGgw/ABosIw8llawg4RAqGDOLckXFyUuUi3xqNCil4oC
T7N5KFi6Se5TUbb3SmpoVgXy+NwKTlxAPla72ULsZHq1XVL9W16r7rsJ8ZD9UAx4
w6Qb2kFwTzBVvPF9L3bwludON45sDMSfrrrW5c8+dEacQgDf1UBYIFvH7Snke4L5
pPRuzK5ZOnXWRT1aVnPBWZEo8byhwYARwJJrLLvoMxUZnbkhwDKAlnBAcvNYGSlt
iqYMGB29WHA1m/mk8qGsedLHWigTir1K9uRpr6FlNvJibxzDNoblFEXKlTZEfSO+
UIvNwY22TZl2x93MH5dxl84nUJX/Z7zmH6VsbdDPii815523vU4TbRFc0nezrpcG
h3ZiHVuP80tP4K+hIZUHbkUyca/Nd/D/iGf7zEoWk3u5haLEkUwYBSPvu0Y/10BY
34fJnajvWdHBxKIU1eVft79BfmrZc41I9yHiWzpTpVfKuRc5jfmGfrYwE/YanTIf
fpXKDMcJ5tGbzljIlP/FOti3lB7omGE3DiVGW+r/52RRiHuqUtTX/9g54RFQkxyq
FaYNvr9/rwNVS9Lzi8ts0vSf7WoT9Ye4rOxM0+sU04NymPmlNiDdVGf0vxy6nfVW
kXajd9wfxxzsnwN/sJxnAjk3x/ItS0B9jafDnn1O1P6Upg95haWoPq/WomWRJERB
fS4kk2O6W6g0HZ1uBS3ao4rWZSl70Jm6qxR3pe9+2p/z69LpABFHhA2jgrDyNSKo
KlL5oL8Gp/m3Z7/39p6o8JHzC3qA8piUDPO4aIV/T05ZjuPVndC/2SqGnupeIK7g
aBdNReweawmbm65ZIAkKWHdae9a+wN0Y/gC202jxdx+f4Jg8AA5GBr1lH8Kj1YWl
K0ozZzLjJrMRooUE9LIMX6edAMAA381BLWCTdxQ9lMwvi+lCAuW00apnMA8uA2nv
XbE46Cqeeqjd12OWj1bmjMornxBoWZJxlhtqetoBQDmJHWMtBLxjkUZuoiA+w6l5
073hCaqHgvdGgoccmFPxdSYhby+2blVvq7zzPkxaRGt2zrqHMEQd1d2a2q8eczuQ
vajrYzK96Zm/hyA4JyaSGhjlXpteBpbiq9VXLgqKdTH+un9WYQiuaAwM9pwTWPbx
3Y9upKs/CSAe3tvnpSbTZGpqTdOqW6W51cPTD6fv7hkaxJPBfjxkd9DgfQvFHj4+
/ZZucjkFH4+OUWtM448BXuFAwoCo+TxeY7VIjD3Bm1jngprauH3Mi+SZSovdOs5q
gnQbxyNSwEn3JFNy8uFUlzn/Nf92Vq9hfGww/SFEnH1xGW0xKYO9b/AC36l/CJgk
h9/zOq3ay/bm8EVxaBuTdovaruTR1nMO/yscoTS13xZOf9twFumYzFFjoA/770P7
ApHH5+8sNaba3P5uQJx48J5F4U/hfY/kHlFZYOnBsIY2BhizcGAvHOLpni3o3D0H
xEo2yzCeVQvKP1LiPofaWykcXiDPjeBMxp6JOK9vSWjMTFTeJ4JoYEPrwG6Bd4eW
3VrDR3NWkFeHbovbUZTWdRXZqvLWnS22biaa4MzX4+cyz9NRqmn+s5D2Nc0xm926
TzrKx63BAGuCpAEODZI3kjBz70RiTyn0cJsT1Z1zXwsvuSsae1ehVL5x6RUIcfcy
Ro3dyDnKmxq0cSh8qMEpcXor2C5XFiYD/9Qxm2sxueidaPj6zDRTCaHciY/2lkhw
xuJ/UO2pSng2AFlolkVejyJaFz+9A3pRYRmSB0mqdnwXnwIOrfhGcTjjIUf7p7Hf
da1aGNnhZYuMz2oXJwlfO7hmTdm7Oh7+lY46jJPuUUbj0oPA8ZVCCG3i963HVZdo
skDhFq74HrpSUN773fhLQE1286pYMONGQJA+q0Zlc8t2jSFP6u+6hKBYH/hgxSQ3
9M29tWeR1jr2qcJq5pHU7xmIgaLOIV2pO6tROeq26/8q1sM4OIO+F6Lo65Qr9bKJ
I82ZPjXGxGcw3hKlwyJsHbZ3B9MnIlIgPPpu5lXhfTBW6qOQZUmfyt8xvTfwKi9n
27pdYYChjeeky5QWWMhKbMilF/LVCgqTvq2c9xp4k7h2STMRNPXMKu7XO9S9I2R8
ayY5v7seA3n2o85mfgGw31NwC3RSCkwvHGd71Ml6oZwAByZl0ujVLgSroBMR7949
pAXVggQW/ZUKoEX4cB3b0FgdEz+JyR+M0FW3nydLXKzU1H+SFSIWwntTjqLQXuqX
juHYpti0+n6KQMpJMBYa9tCTNsnFMNJLZ+Mu/ONSmN4umPhqyWIAmmB5+qp/Jwt7
7fS9fnOuA2l+Rv8dedklRoKHD3QRV7TJq1V0zUTJkqEirEsLyE5444SZpbg2eiqq
xFyOMOgIZF1t3r5ReMX0suxBUP3ojyPi+zkvE/pb5/WnriwI9xjdkxo+wae3+1/W
N1YU7xzZbGImGadyEBiSH8IOjcUTaUuN7+dd55ws87zpmOTdJBYX5n71XfheSFmU
cnNnTLVBIoVqihxbZR7gvEK6MUTNiSI1pCkoGnAPmkhyQjrbTMuK9ZTjXnE50ppJ
CK7kjvCZGyFEKZMNvKZyE0f16ItgNdmTWq6yiA8WI4VGHAjCUDjP1rMqdU7K49RC
fHYRxJgflPpEgD5XqOL/B+PJX5wvHUG1ZGcMEyL1e2gZqH5dpesGddvnCRg+ZH1y
cCxoR4xN/doNNEZ9jq/IvIqGk2Ayfbm46/+9iqhJ1teihQgzftcn+2ur2TS9UGWE
sGo4v8PSXWcyZpcv027Kb3JZnFsnleW6qYHO3ZkTheqZuzXGp//b3JVFZ+CoUgS7
FVte8CCH03vYZGuu9kopnT2yEObACxIphelklKWgSxvh1LCJLxBkmSarah4SnSxp
Dw/lTYip6m9mKe1uU+A9RfXxZ1JH8aozBzPoVR7ziinXvzH/jd4uClkpV0eXPU4k
r8BXhYWtLkqqshbpIUb0EosALwTYWADaVgw8Hz1brN+5sOA+qApuO7FXt/tjCyXv
PTjeWvhoodYtizsN9bKnQJhDdA68NTHvTTv+eZ6HWaZE/39FfUjGWXNCBpusWhFo
76nxolsdswGA7hxujd7lMtEt7NaEJ+9RtIYf1MwcpcUAepdgt3TBt8qgtEVLH6yG
F3brG1J2KLzUGAgq2BDeMM8LM2RIZVT4VYjACBie3/28J7u3q4fuDK25wiNCudTQ
rxANRAKHzL3w3VdjWrV9NiAhXks72LiUvM8XyTZm+lJAc2dH5+gOsaBTxiCbcoxv
DqFGqasoJN+eMpe1l0N+oMGxotXDTjfCN3JbAMO4tfBaV4Vnd/JegzeFSbksTXiT
kW9U72wbKPCosiDAOSHEVzwUYHeluMwNwGyIMxDS4ORlPhchHo+sukNqV8zrxBVe
omcqndIUV9V2LQAATChrJz6dubjNwhba3NkTNwQlNnwo04hxfu0mFkoXcconxHLa
nawR1nnTEUqn3ZAq1N3VmqYUUAuDe1NG+W5Ea50HxjMwxNKVolt8h8ke2s7mpxIF
mu8DidDfpIwhflbtJtTY4Xo3PUrWlHl2Lo96Zf7AoJsNm3fx20c171GeaN29lCcV
a0a258MfeM/cZTj57PPDt2d46B+S4Sp4+SSrYME6tg1U9hfaHanDEaz/5HfeYk1z
jieatACfBbW3gKBpaElsBs0I/l4U6rt60KHu+IqRR9cEZH7jsjz5zjrofcck8fU0
0ZkzBfno3PE8KMoANYjAAGP43yfiJCrqyDUNwllJ7CDFDPpc1DznfnLA1s1HGa+I
rX1UKDem+LbhAaAMn74o0YGpbghEQv2FNd8l2XKD+l3X+l7Hz3kHzcYzfOhRiH9V
6wHzNyFCGD40rNgLpngnVW7pVFjOW80LvYR6py1axpe9UbF+xQ4efofI8D+t/SrX
VhnbPBo7rgA6LBNpSEnwOWnC221a9K32Z9VpRWRBB1xowrN8RwZ3CAIsHy9IMEPq
5T9c9bVZ1ke7/1f93UC1MB1rRM/KGK/7IWenKDj+OEGjIX8mnCQz2x8rI2k7Uhyj
bCmVqnUvuaTDYH+ZZLzJeS+faP+8pbXrsusZNM08MetU7E0hFzmz9PL9IGKf7NVz
qTtTAbPnXoMhGyb7vL2WK2GA1VedQA0xe2iylvJLLg/YC+QV2g5+351vyKtSGnA2
vw+dUQ82ETj15S0s5xxsOHbWvX7NoM5YZcN3E8fW8HcmWcVIBil5XsrWcU1on39N
AUdsyiYdVb1vcNBrk99tnzz/NCJ2vyHZkhSnzuFRL7eRboXkbTIGeeZMWndUw+VJ
IEyah9Y9Slsu4gUEPZ3ZxGLHC/vbb0CzcuK6K5kOjdOGDux5mVrtH6MnfuTeuwwH
2ZfECfj4ANhyUm5gmmXXkHPql+1I1Mg7UHZAkM36Rl+THgJhsvyPdHaLbQ3STvdL
lT3CnpbBDVIybFUTKCK4xV0NvNls4Oi1e088YPOs01hRrGJEOX3Avx3y/rbLstSH
vSvLcnEaCet7H2Ifgr44O06QyZMHYTCiE1KtK+zKFSyXUQZ1IJAqWwm12obCD9rY
5X35MbZ1dugOZxOMee4MB0YgOxmvxq+cF8Lr4IB2ulheZ4hsno8bIacwc3NaK64a
Y0t4Ax6kgsDmVzmZ4z+YX/AJE1bnyfg0yQLBuQ5WzkCcK7OsMlOfJc0tF8+mWi40
Uu/ngjsS7+vuTGOGi6rux6rNjX73jKY3I+SaSjT10Ae7pajg5e6YIUrolZ7eEOrz
mwVNX03AJWl5/H53V/25xMkf7e8EQ4b/7+cGGWTPuEO4zZ7W6kpbrxYQ/aaOLEwI
COxCqEIaBhInmXAq+9FXzRUC7s4ORmy16XRCCWRk6pimQ/WULTf4P5GSTv16Uxei
Gd4EM1gy22WfFTXNmtocW/Tq3J9JLz+u0XfXYWI86sTFJ/DjbALh44rYEnJo6OsA
jMc7W+UZ6lpHxyt7JourLATY7AjRAKWLR99tI4eDZj0Qz8bRbLXsRehDIQ0p5jrz
3EThDfQGGRLQzSzNSfON3hB6N91TNtU4JDxn4wMRIQ8GWtYKeJbb4uhYDmeZlRuU
frQPkzW3kf222ix57Gn/sASnmjmfAZeiC1NL1GeyONqG47NWLxwx6+DVptmk1fY+
dinenHQZLHxnAUIyP9Aq6wGQ9Q9+mBPGx2kzVJhv5JTCsia8+yOi79J2nbhoBdlk
5zEIx2LzQ0D10XEUmXXIpvTbm7uJX/GtX1aTsMhUCPFwjMr3GFl6oPyfX97zd7KG
LX9iDOk6pnaLDhSZzQnG678M31hQdVHMy3iXbD0b0DBP9UWNueOEuokf5b0rciKs
+R1fX5om/wzS71zwj4VF0F09LoESF4PbRd1I+hbPJalBxkj/ZfVgoZggiVktVkNm
ZX6Y8658/NAu5wwUvkh9/vNHW+onjWNcIGh4hn7cr1tfwbiKA2ffqkmXS4ae6+ro
IxhASEOEYjJSNcOtiIz2BCibVCA5o2a0dTbcX3DbhcNtPlvI04Z4JryOk++T8D0R
1k4EDtJGT5WXQMZvJhpeMnZ8ltYbfA4v8e9VPa6usJGxrUGOHboKCyMfUz9lvkRa
/Rh7A0Qebd0h0zWh7o6M/bnX41/Rx8VXevLWsIBSByicACmoBeIDJzckibsxVPez
d3rvp7z32j/QJEYp28xupizLwg+snwhSiG3q5EjYMXI+VpX2GUnmHzYl6WN1+n9R
Dv+5B3B/D6w2efh0jkpv7YbdyqhJA81vK70qi+rrNkVE9QqmfsFOLAY4cuMQO3td
4qY+ckfLmzLoG7XKHH4wy4DuGyHD9h/obA6wwAXF2/kxEsap4oZSjN/mtsa9hE8j
mQ1awZrs5jhbYzKu7EzyWzfTcPYCvuH2vZTJqSREv9MXtsUnyJvFWUDa57oBJgIu
bnsPs5r56MZ+TFDBNV+AWTzHC3eLuZ8IaOKXpsvWlzaq5brd272Dkif6KBsuQBW7
1Qb2h4FPacj9AY3lXQKPM25PnJuoKuinmaqvsJsufX/bvPavEKUiPt5IhsjwoL/x
SXd+aCWTvBpCCT5WD7fNXx9ZDBN80bRI/QQUjPkcuVfIn98t7WBiP7NvrbLiVo00
/J9J2t9dyueujhJJPUo/swLidN75qmUER6MK5GOU+d5hnl/EdQlBV6XhcQOPP1NM
U/uNPu3STJYm9crAVUjr9BwFNjLhkwnJdFM+dZkZvtCADihzstIlH9GCN19YZxyr
+h5RoAxsct/JTwEwMQAFVF7LaCdgDeUvMjb5I6JS/Tb6WGAuG/4k1brgvnQKsItX
NrtUxhtXLDgaH0e8uHSj3NxIurs5Ng83GoK/PuM4Il1VzwxT9uyps4fApyRrYXEr
Va7qRjR/brOQtVfl0uOe0jQ9Ii+pSwbG9AiOmqAdlhxoNVdohpCiEENtleSmBfTo
tDBksuYbNscFj8zJIW7UC79N0eETBO9M2Z4BrgFF8n+gwCQR+yZttuQFwyesEPME
YYpNujBl+U0lBXznXf0pHbp/rfLzn43oVGHibOrpikbjd0PmDiGzRad/xss0hhJ7
hvwuOA9X0P6cuQlDOVRMjuHGoxEU1JyYigPKjFsnZXFAs2F/hlx0rElJuoT3DWjb
VBYAi2nrclPCoIOPMv0mHY4otVP7E+C1jgKxCLWtyiMPlFWDrA3xWLu47FyL7e2z
M+eZq61dBeZnGKL6Is0Yso2icpz3hjetKM4cU8rBIh/E9xzYGpFMAVfkYrf2SDTh
GxSVosDxl8m34LIZcm91VVqfrAUAwvzFsNOuM8QorazVS/kXIxbN6yWQhh9LRk2V
w6R9zW83ITvqSCM8SmboPY/hVm3eO0bwFsWN6xksYYBQ9XaJzLkRYxoQ/cPXd+3u
G0HjuFrQLgIpX4vvsusYTfMGjrGruuMCYo0WPIFQMISdQh4loxYiUKQ297+17cAA
xEsIbWDV7duzF0b0qVI1THDO7PKJrHFQiD/WbCzTcGV1V7WKdjArtyEdTZgBh5uE
CUwYB2wERVXkH2HMd4gAvHpM72YLzZcur1/lyNTQ3dGeIuq7wbo6bu+Z/WjrQX6x
znQE9ZYonvRa/A6UwMmWY0S/huFvEj2qSX4HHVvDgtYDbr3lG/Lkrfgr/Nz2EG0E
13NBfz1C650EPEIrAdbATpLt/fxriPqJ4+hYe4YYvav63sxutXK8p+rc3pQGJooY
C1nuZihaWUaGkEbX6554Yp9jED9DsLWOyXDN31hZbmI9TmF5x9jMxMOfJZPhX+Sn
8HdR74m+T2q8DFq6WVfiD3XxNK9nwqmWuMh0wMEKiJe0NaUEPbeTvwxx9ogZqH8u
aUo01ZjWJA3BfuFV/SPExRq9eeq/m0gZSNloF+Kc8li5T0goR5xLhDkH08o/COAJ
aqgtBy9MZrBf3e0t3hNU5z4SIUFoYdms0Qih5J1mFV6dXSWd5TtuRUkxDz0H9+nI
kEKUHJY57y8x9i1F9B61Sbpl26M/oCDWLjtELWC5jmPr8HUkRbp35kd4VlPIvhFE
Zm3XAXrAUxtQzbZUaonJ3l3WcjJb+TT/2IgidGA4B15EZCHir9YObWk/vdNiiZwg
LKznI8u5Tcks+mCGs9rui5NlPs49IXJjKZA7lFgkMuQrEsMKfslifEA4MlLUO1+J
QhWjYTe59SghWhwnf2w6ZK296diOchvkubUJvAyjm3aJkDsz1atg/T1pD1UPOyvL
wSwRRtzfNzzG7q/NcMUwSMaOsfAdv7ljfKYc5XLnD/pUughH6htwdTvZBOok46Np
aa24gFSpQPZVBeDebH429OFCcqdMnVyNPT9yReCQdwBk7A7uUck3yCCC+3dWaWYw
xY9LRtBRb5qTsTeUwX9ts04gtS7UKESPWcVikU67+2apyO0OQy5uomsvOt9MokzY
0HOtljOGqb8O8/dc/twPf04McP87mO4M7TqFMZHYZGTY2iSoXueJNYwFpdKtNQ18
JwXEdUExWc76rZtKnOpusV3Xra53DJR4mvPSkmTHASgMKm8csJvLnIQ2ELsEf6jG
LP/u6jJ0g2klac8/Rf34hgDlb0ZzvE5iUsqu4hPoC/jUyRjVRD6hWNDnDV/QbkIS
oF/2L0RRohRiYMIqlG370tHnL4YFDDi/yOx0RZ6fZDEFXjsgJSwXwYQW9KXPayCX
vnEa+XKJpR362/pBBHDoEndsxP57CjBBTUemXQ0lAtdS9riNGivMeIl3YHO9uM2P
6YgJ2uWquIViY1agXeJ6ez71KwIhAuPVcY5fOoFT/or64GJ1v4QUxS4+FkjkOY5W
A8vsVTOH6WquoOkrrVjdJchsbephYD8c7KhasE5RSUoEzz4sKka99z+HTEKxZiom
G/qg/WX/UNCxBWH73Z970x0d9JTBLskQcz7p95bxHj+i2mirbMC8Hyg/WgdoGhrl
YLrIqww4L0MZMjd+2ns5Vq5oydwu67tTWMce3OUIYfHKudIwnV9ARQYFBRmLNUv5
FRppPs1DRRKj7g9BTi6rMzPNgjy1/PlwrSOnzWs052vkFY451kE4OsxxJ9MbAYDu
xnJ80OO3ta+4SyIxVDEg+TYOMcddFpib09t50YiQRg5ZP3QW82WjCKU2KLWtXO2/
oTSn7ZNYMuLReC0WwHS56vZKkfApmMyPagD84zOSAuRyyPmy8jgjvacwxZNvbHzg
kOFkjbTNvQHQt+ZCP8Z+L8qpeVNes3DDCgmT0JnYRXAcBe7KluFIpKWGmOZafckK
eSppDQiOQ3Mz9sH9T9VpQ6gkX7LLw2yNTY/UyIr9Nck/pbD1JUIwVCUQQtKUuYkP
TpErjHoQ0qgeNG/byEiHYQQ12lq9qh5L6KP4a/VtSPClEsMvEcmGSpM7+yOeXG3J
4B5j7ITZqZBc6TBfjFxc8CEZ4VZvtX8XHcls/77NFNITpx9m0bYj7j1n2PhQ37t1
Uik0VG0wKRgVhgXT/V4wPR2zuAPpjjufjtnyExp9Razus31HxzPTrX5S93S5X3Y2
4kFnkOP+L1Ah+aIiKvAA+KN6Qm6Vlj+SKwf8iEEJNE/k9Jmf0AS485z0/vgWUg0A
KNDWdNQmylgxiNbEhZP4cFK7ESg3KTL8AFniKPazd7EFCR4I1TRKm4gbjE5wX5Ao
eobeD3mwWPwZLGz7lhH6DcQQYbl92W+vA89yQpfEjXuCNuh8SvFReWUZciAlrT/+
4icPDHwITYXxV66MiAIU4Hat4mMucpCs4/Nud9waqpOVrekY7TGyh1uYVFDUJmGx
fHpp8CHDbYn12HiX1vUe1d1/QQqh/9Fd3vfcs9n5sMTFBAhHvyizRKGhSa7QS3Nr
DfGOtq4/6mPwA4Afb08ZjQfEqD281xaP4A4NZwOKA+SkQQvLDvW6e7F2Gnx0dbS2
2P3IkZGVMxZRUBh8JSzPulZBlgqI9sUfWngIWiIiqcs/1QwvxGqqQDFxBPJ1OFTw
iocarcGFEJazRbRX3IUYaJ1/A3HCbpvc3wh+y8BJrFpWVSNgDPQplzCKJJ89Nyw+
NSQ16iYTejoZWe4GLN7rlTHuqP1oA3tmTo/z/JdFaqu3+hpaS2Gu1TzYKEFxO02P
ZpB++Qy6l8fcEqdJGvy/6iSOlDfZQivPDMGUokdX3XbqdH2wIJfjJXOqhNDxtvii
bNVLR3LYTHBXBV2GjoVIwMbsEh91ax9+ZxxjdjHy4GOvg5njxtDPggrhRM8fgC2v
k8bTRz42Eu2UAfXcaNkfxmDPT6gAg0QKDMMt2sOXs9QQAfFXjKzTQqaUHUGOThAg
JejMXoxRuHKNqw3iYgmpoeKt3+EgmiSOhmQXshis5FYeSZIl+GoMtdJ9vtHvHm2j
lEm9fJM3sIEauI4SAvJ1xZ+npGJtaRAm4kakV0bj2hALWcY35eVw3vuVq7+9zbxA
m5srWoXQ+IoOTzirLc4D034mPRaFsiYOrNtFawFvzhosn2fG69nxQq2RtyF3PNCO
8htRFgDOa/murQJcvSiSSVjvuRD0OIcRLDHIaiwgWMxjBqqc5s28gJdlUILx/YhN
l/JnyWWiWNIlfsVWZfvCTPwmu+In+IHBGcIGNQ6u145PgZ4cO1/+1Yx520YDyB2C
slOtnPUq5GV3BTAwKBcBg30GgiXJPS32W8Y4nrVdlGX7jmZhx1yt2+3koBAe+RvX
abDOLFlOdj2ZJ1lKdwx0n8ckSp1offYxKbKAIwfAHH5Q95NU6FQRu+n8cmlknjiz
zl9/JKYICmwbpxJP8AUzm2Y060vkSqIzMd9CtBzXu3IkepInGNFhsdEpi+DWwKj+
s/GauvDoi+ZaUXLMr4tb7akRTWQNGZRlhcMeeeW/wRx8S9OeInQ+l46Y6+u3pl0u
Wj0npLa5DoVTvgzNodNvZV2VOrTp7LtgOkrZmOZzQztM9K8zFll8qDPG8xOgt6Rr
VqxCRkt232INfnfkXZ+V6jfirtUzejPVZ7XvA8+Yn0z04W4pWeLVmpEmTleR/6dJ
wu1U9TCUzkm5guFwzfL4FttTWzpCHP8JpvQT8WnTR1aGYx4F3UxjRNgB/BOVfzK0
m5zZpYhywMn9Ud4V4idh4Bksni1npEGTU29aBRx4A2AobKhCuJWPmzwvPgXnWnl/
EV9Dfe/Jplf5VCsVmiy2rjUlUhjXEdzIhslWePJiyUG3i7DU2pfBfPx4jjnJUEtf
PrxjXBLFcp8yAEc3O3Cxk5ULxXy64yEOpuzrvrhg35URsIelm+f4PHCPcGq0f+Ue
X1LlkRoO+658baKLa56p6vQR/SEXiV+1zhN86xSIn/N/aiD1Cr+WgmqQGFW6/qsK
WPKD3LB+Ch25klG8kimbuJoaTBuUIUA+fNNwEXAeSGJqVmfT5BZ2dMrq+0qGe6+J
vEVw46Qvmw6yhT44iZTIgdRJFAlQG7A0DvkI7mLW4ozLNdkdQOWfn5GUKqk+0ZkA
ryJN1losYFXFO3i4MEiOxmTsVL0hZKTXQfa9/CQTbaOuXEWsS3Bv5l7jUkBScGfJ
IhGEoVHPEYDnVDT16OSzuTbAZz6HGk+laRjdnR03f35A47OZzyXzkZOt0G9r/LkV
Fh/GYgRZC3/eup+Z4aAgoUV4MphsplpbrOKsFL5Hi+yGGYH7KOHqj+PHCaz2p6+2
cZu/7qUzM2VmtVFrlRB+3AEN6Oqj1QNRS+H9XlSnpoVzSWueDPoFOTOtW5Hy/lpA
NmRR3upSSL7yDbkTPTzkHvtn9JVdFLWzcvEP7WlzOZfT3XXwodktpTB082UpF5he
MI+3kysr3t61ctJlokjUM7YcSxGd16GsRGzt7vPY/I5mn8GivkRdHlJSutAy3XFJ
BzDa0VKriA5JkFfZBXnRM0Kygdj/BAMkOy3b6FhLFHt0StieT7yfql7zLcAW+Mkm
WbcbXIeoqhMxWwZmW4gvYqoqf+TQAjI8q6r1bbyhiBpz5sxclIaS/ll9VmOTMqwK
wyaalbtbT2JfijXLcfZDrT0MgQDvXfOIbeNgrJzHeR6eCZA0i7C/nPqwtksTtbA6
1k56GVFyHL2BIrQh4Qh9cLUf2Up8fwMq7Xl3vRAh+0ga7c8IJ8v+Z6li1sYCNoEy
EsBRQAVMG9wWKIMjYWhOiQKb5yY9q7HQZk47sGLeCf2TRkEe3H/jBfxRzKgZaY9P
AzZoiPxMAUOaZSlwxBaQXXU2OOIuy1qi+cGNGibXAbpm7BOdqxgUlGHy4ulS7kup
2pyOtKKhLHg08mxbjmYM/caW9Sp4c2x0mSyDpG3RXxUH7o7Tjaz8l5K3OipeNPr4
cca3TU2LgF/fG61Ux6SIg0Ew8JD95DfU+97FrGcDVqpF6WaPCFCZdDEFF5WoKB5V
Q28QiWjfWMQuaB+N+e3t0tHqfFtby/sAxd8RBOUxaGtvUtW5ONhexuNPYm5nrvzL
yp9pMMobMwCCy06l7VaC/3CJ2r/w7u3m4UCYxnAVnzQm1yu3sTcaOTxm/3/yM7pZ
lpYKvVMh+6/+s2qZFyDxKm8G6RotXH0KDV8d9khoC787weuyoxu2VneCiWTdoIw3
eC8NP5Ps329ecN78NrmubD0QkbHNi9Qu8ymtZ4THF1aLH3/1U1fATLxI4oOGTmUz
uZTjeR9MRSU79zOzTNf4j6E6UFgdkpcKCyoM17tbmuXvJ6Fjmjux8r1o2HLvNkD0
2j7cIqYzF9MydEjuxIuJcMba+sWLYd7TfOV1HWmm9g1Y80j9gwaC13pxei2EAhOB
rIo2Z/fL7gL2EEFpvB3d26yshLqsqLHo7hyh/jPxEe85bnSwGDYZPymEMRqC1d2k
hM4C+zY7A8YhghXXLe3F2Lgm9+wjBPX9PTEaAsFcdkC06JB5DaBs6TILpCX9HPit
VqDhbji8ByDd3a/NdEhbPb+TGMhjw+esvPqo5PNdOeNo2rHLEhbLI63+0q3GXyHu
A4mqrT4HbxrY8c5yiIfm2WaMZFY3BIzWK4+/NDNqEcFxpuLOeebxL/cFFEh3w8lY
IHTduIoWzZ/vi8L3kQgxNc/DHRtOty4ZVF+YUsVVhTSpE07CXnz7S5DEoHZ/M/b9
cl+TYTl1/Cd+1JOJaqdnq6l8A/rPluFxpZxQx+1Ldur/Otao6s4kQOqxkT9j6isk
S5rIrNRWnTqUr9TRFnBe9onziggpDv9vrxG+VUHDbyt0OupFrKKOAB2I3gNBLgu/
MsEf8EZYXfDRtm5yv5q9MNReG9aEeUSToey6R+OAJbSIQwhtuBGUICnqfI9t4ziU
hHQxqZ8ucziCGmiTKqtigpnPC7Rrn33dDyANaxNoFeio6h//jfu/DX8Z0LqrBeM5
XCFfqAaCsUfKAbiYJHq0HHvkC8Do4elDL6iYL6VdlyavZaurTHtnASFAQz8aenMS
m1CKo0T2xDea8VSO4OekxXCza4D2ZTuUGhzVZ2QuWvY5kz84y8ATOCQKJvPKiDa4
sli4s3RVguFI1JM4Fvm0sPwLOoE1y7oqqyoFJwGvjscNjMKOemhBh/kd12xNFG+r
muTlSo3rjLhIg35sYekiDKdoYixvt78SfF0aL3ZfQKONtww9ASZ003uzSOy+NHZm
g7zGQcBKL0G2EjviV9yNVPYxFFkY07n6KdhlgtvhNIgmBpT16iVdOkRFJTWeGIl1
oOMWwy2VWTTnoo4MkRTclPbrpjOnY3Ml4F33kBAt5/C2qfHIzLEl8Fs90UzRHvzr
gyUcSGC6IpwnOU8qA0xXAziKfuFlkMvgiEWtluBHt/tF+tRUi68S56e9h3kKMwA0
lGeWYYodMXi47rzR0KbZS4TzuLc0LYuUOFt1H4iqfsI4GSah6ibhOgeFdjcCJDsu
AV23VQr4trgwX7XSzp8DdcKu5TIle1ovUNnBEh9l9IqAqUKxRgNuYOlmhvEAmr/o
tDFkC1NXT9pLpZOft9rib5ywRwegbSmH6r5k4kIa35tBdw2D7O/uUBx7Ctf7FUuR
FyPFb7kZO9wLzBqnBHs/evgFLiY6EUKo0GLAGEIWw+9eY06RJkXmUEBN44DkX5Eu
rm32iwNUnbbgK6BQGlDKDlBiVCkKsyhyx8IhusbuNEKc/3/G29E5EVsh6XFwk1gP
By5icI4+ayAXjODgYI3tinyROouUmscAAhPQ1FHHd9BtyGsKEefMGlRmUEnPGLcK
slrDyE3BR5sTVzQnVuJ+i24Lo9EakNf1KA0yqyZMCfefuB37Xh7ttcdvSLBBPB1y
SC9LqXPvXK7KMmPmSwUUevQeC5CnzC8kIXYdcI3r1+e+tVNjEiJVQDFFSPC+sHHl
7opjT3fJe4tyVfg3Jkc1TTDXVLzhOz0KVlo3lvBy9p5zay2timImPULuJ4qf3Gxr
/3oDrVYpOPzpYXAM2PqhN6Vd1OTJAj3Qx4IS5HNgrasQpDa37jmFxipV5IlrkRtJ
a+AhI4dHgwUuuLkC9MMuHsh2tEV3cf/Wn3oByv8j54GdFP33UmY+HufaJHVBC27H
1faAT5VoAOg1xwdrEBSHzeNcrJglLQ60Zl6ZhIrVxXXO3usfKOkx/U4Otz6G4T9V
WzySBvUEi/MNXnewWb0nGhuWktXAj0tQQTWCtM73bVWd6B7mVjM9N2LQqNnBNg5T
0H3AnyRVmUhv8jGVFX4lR+rCAUd+okIf7vNcoUrnDxyN3WoQ306LjqhBn+kEnT9M
J46mNd2gXI04EwXbzZuQzCT20xIKG/ucXndhqppInDkBGhiQ/cIBvWLHiEhE+Qdc
nAUy9wI8XaFbZN4jszR+wqq0ET93MamVJyhM4u1qt9x4fvKo3lV/PlZmAfbDosBV
hSg67P/HVyikER9t3/Db74CrJzmGqJpI5YSHeVo66nUNNSeKwC+G3n7z7K2QHYot
6Kb4oAAZB3GGNPRGjR2YVZd6O+8aQe5Uwx25oZ71ZNmz/yGAF/BfZwvSXDaBkv5A
oCF8+8eGJDBCQFpJkpD6keuS+sMrWJPRppuMsxeD6z9/Qz2U5juGYiaNGqrIgAY5
XmQHKHbDBr/yvT0kUI24/WdeHwwLNa+YloA1x9qHWO1Uq73pMzxdZFfJdi+lydaW
eB0pwyWYv8om9LAFHtF69S9GaYQ8gRlKBrVRq9ovEtsSA+Q0VPmNpLw9iZNVDAyL
hPqbjEmTt4ITHMjCkmiukZcV59+y0nCzjlUZBGuZ/lKluR8zfeG3jZGZhj1Bw8rA
3VUqnqvEynK5ksNc8x98oxNS3Io8m/spEBdm0NIVCTzlmIlFIBykrQ6xEcs6xDqk
cA3FH99+Neu7stQTbcxvUDyX6DwB1I/2T8RvdfPAHLxWlThxwhghBl8wjO+FmhMK
aA/IDVBcS6XONC/G6z/jUBSfOj4j4YkjdiNpcYbSMWOC3kuoy30WjZe8ckgmoguP
hXugUFIkgUtECBOECeal85diRWP8Qfjaf/EF0j797ajbljHzOIyr9SxvBKCffCyR
odJ7uBBRqxwz6vhh6L+lUZM9484POd5zQDFt8V/woPhZ4BM1LJ4dT3HM16T+9rsS
Ca5QKR1rMpjK0NUUAD6/MCOolmLVfM2xUDIgBXnhmGrM20kbh2P1dIfbJRSl2UPy
/ERmDEdgi9mhrPX7EoyXJaXOZphgXMGse6V/U73W0U4oYHsNl+RxORfa+7SJbpjb
64lB5iqa6OFrQ0U05sct+qRrMn4YlOTPxFFfXLqdPWHu1QdAuXxtbZ5+ZsC1QmMl
0+fqYBzpjO5u+W8gSupmRo+Okk082KLUxwsm5kQx1IuVgff6vqY6znGWdpvJ012X
OiED99a9135ACe0wEuzzCt42RVYZOZlIHlqtZS+blj3M18gYe7YRR+xESEHytA47
+w0dOg2TcpIfdPWEt0ZR4eSudrDo4i8O/qf7PwoQnLvFajdWQcbISIu2Sb3Z+cQh
qHlZKi7qbrCavnf/AnIGoHvph2uKizSp5Kx/DTz7AXs1b9WzdVCTHhWDcIp6+MoK
VL6iEgqh/llQG3XiSiBFOoTZyczTHBg5SsHYJV9tU1MWcukIHVrfscTQXz7sN3qT
ubrOZ/OPmR+ql/eH1H2aU1gyrE/GWJ+doyjNV7eE19/QFT46JsbuM4wyyrwq3nP8
8PltVBQXydkamPmfPb7ZqEZqBiXX0kHbfWqOz+nTIZE4zLt7ez6S/IEz/Rk+BMnU
HoJueXwfXhxabboA0w2GIOuHyOEBlKPI0hVkO5n6sJSa6waOuuELR/oj686soSqG
AKS5dlsWq2PNtN8iiV6rfi3CJhCLryBNPAlNH+qcYZsas4l/cla/MtVlDC88clJ6
CLytufZZx0qPWhYmlTzsX8Q4eS8ioVJN4aYnsenHZu2sQZkVC7B7Vw88p/0ljKSU
Df7hd1rvxkC6UEDFzsrPBV8w+/9Gq7iVeCJSVkZrxy851z0rMEgwHJRQ3NGt1eYF
gIeBlL28SZcvap6R6hCKA+/RtCCXBhL4aL8eCvhNX4ECkQLBZsTC4ao2cUPNslbi
T82g+yMg9NJ9+Jp5HX2VQi5GQwZUpkU7voRdLvTYiKorc9SNZ6ldBqN7A3SA8r7y
oZgLa83isS/d2UMrqgQBgv4nEEqFyQj4XNqon8oRcF3CtKwZeaABrBSvKvFLZgyW
CZIngrVxlQy0Zt18OzjwO0B8wSXnw1/qp7CVHym7AOxEMiMnWkZlcaDuCnLHF+uO
Mddf8rc3H3BIev/d4FG7scj1hfSj9OFWzr526qlmoZvQP1tq1eNFAtWetIbF2Jbb
NM/WNjcGtmaLmbC2e+qL72uMkFgp2JZOWQHUqHwFzSSz16boOhaHFR/y/drQggGh
+D7uj7rX/GhOaUHrSudAoxURS5qskvgcEdQYIBy07kTsmIwr+o7UCG7AFgvsKERW
mOEzF6oPx6bFEqhZaqmLXquIGctWGerZv4aJOZ5iJsGPhQERXxmUon0sE2hUkHkT
pMTluIxmxLEjYU/kgbICGJKJOuT/6nP2KIGhkpiqTqV/SGdAVOMlnxCZloHPGcc1
wgJEwEw8MSDwf8f3xPOmDqhBXTjaideMWfjX7DvzDr/tQKMH1QUsmXtroYEfVfbB
zjU/DO6YyBXtl6S8OlCwoG/mUKNu+oLOWpOpgsTMNo0BD4nBCpKmaXLgndUuPJDY
AiXOVXyDJpYvp2FHLIjQivD8yH1x8JRSJ6GC+aBFhSEjQmoiY33l2+iHVwp/EBbI
c3QktiLCsdWZ1V+m6Okj0W1jdOI+QVeDrWw6tCc1e52KXUPBKxk0A8CRW/FTmlDG
/IZSo0ZgDm7D82jFyd6J6+/KKkFyzGRhXNlWB00Oc3NJEMS/NtiAiztA1dh7j+Kb
2Yw200PwnVJqy4SUg9fMm38I6AXEwgSGJ9fqps223YCgHMWk/nsZLc/DMiqIvfG/
F+dvUfLGLjiBfsnROhTlzAWwB8SrzjTaH9aKNqg6znJTXiyaHRtNKt0aQsn+G57z
6tNqVrQo5HsFGtCw5dOKPl5HGivnj7HrBXvmxClC67L7dd0h4FC78aIa3/ErjeFd
8cFTZXr0c0JUgUb6ITzzcKjRX5aCReWPMY1af5/vN+Q4tqA1M1D0gl3Ch1TTSSr1
UpD3RB/4F7ASFVjrN/i9Xoe2MpLjFtb47gjaF3y0rpix1B6qTjq2JKotLlzMqPIL
gAJyFm4ltFB2Zrv4n7M6/Dw1xTO3YvaP4IiljDtLGD1nZn8OODW529lf0Q95+Em7
Czf9Q5jwklDh18IQDNz2eeaCewkXJm6j4fWRSzNrusKeNRMoIfJwI05SY/DRwvnV
bWntNB9fNi0aFHnUNNFHI/LU/HxTLXO65vL+02DplPl/Kmj63V9u5ZOw/14o1w3X
bJQvV3W+ajR8SW4v9Hx/pUJ4p1LaN8wfk8sY2iSGGwZKAXlGBBjNF9T/wKwhYyKh
Z5mEW7NCw+zZSR/z0i+E0KtT8UytkJntlDpWHqCrC/uQpwLLgEgQ0l624wF/vZCw
GMBblCRhNjjgVOJeggXS3h/OuGoOUtfNwlOZUtxiXipDMGCW+uTnCRMfbBKx66fp
1XDigAnv07PAgeIP4Nib1ikXQu6MUzjkJg6emDUVl0YVRqjx3lvLEdGq95a95wrh
h8SqUKHpG97G0FoE8j4vdlrBBJr3KIpPvlIzVLCuOQp74Cr9+TY1VqYQyVg0IFep
GsUgxUsqg2qQmq8laq46wPbJEhVq835xLEzxsj7a/w+shOJFa90RgGMRRth2S7cq
CEzLsCyCVDPTaqTq6Hyz/bMVJdjpBJxwDU+yiSOF35fsohYC/igWBgTkRKi5MRko
xV+K/K0op5GFgJiIxj0wuUTcDtAY6zPqfCZoRzbcG+s99992DNmtQ06cGE67bVUF
Hle7VcJMUG5JoLxyptlxtph+uIVda/smtENc8L7cn7A5TjQaFUe50YEfkv4/tEUK
ww8Ym1t7DA90eB2hFcZJxQ1hdwVpen0/fb9x1k2azPHKBzi/jPTj5s7vb9mcYGxB
c8qbevkxJPDeRy0yha0PElSOBCk69C/ZQQl8liX+0B4nQK3+irfTQ3GiWw+8yWCR
ntgaL/Z4GjnqmsrFom4ln96zHENWoAfVKS416ZkoaBNN0rtErhCSKgO/KimRcTie
Fp4/VjlyZ/kE07fpQOHahPAfnc0E0EtaVvYYXoMAmUh7YAhE7lbQ4KnLIXw9a50k
atDg5S8yBSTuMtZsrDx8uBh2uAM/ROoh4dZCDaFOdBQA1Z07iIiPSqKUNrTDth1n
l62wllGrAt70q6lsWS20TvdVu7a+2Z++dKonRN3pk/brVYTCucTAS8KQ+5iz1fz7
nLNE0QrrgtRiO/ybVbZkAIfQUdU9IDNz/NMGe38afQ3hBVuffcoagtD1G86v98Py
S91cLl55DZPSxl9oKJdJeVXMEJY+NizNMmN3F2qUdIeFC079Y8LTLNGJ53KgkJOZ
aX9e0xT+jsRLeJhvQ3TQICwtpXtk0f699RIN377hiRBwMzg3K0SOT9GAiEWrUE5g
8QxPgLoGk1vT73jVg5oT+aM5aGYJ5BO6edfMiQ12A3MF2a8qhh6kx3ACVpbvmPon
mhw9w+WBKW48fx7/ehcWgNwl6he3I13DJC1ffxc6sC9u25xMIQFHwbwZP1ORpfdx
YFRmfYj/jgJV3xyjkjNZI5xTz1pAS+WG68A0MYDI21lIptsXJTCmB4/5iffwJpvI
CVs0ycCSIZBJ+XO+h42MJpH+cOYQp73k+QaBdG0DpDPY7yuXOItF4G6zgM6wjqG2
1/0e9YkDZOZ4NxANptAdzxWhViVPLLeSJuJHeIKATB80sH1LIUQN+Et8sLIjeHy7
ZJEvRBWm6uof+Nkn3Yn55Q/RiDRbLHVeDfmgSx5bvBvYzuLPbe5R2gcJQZ/GUVT0
vHZFzeX/d4KmGFXGDbDLd02Qk10V/LZnU2e92XRUT5W5GUe8GZPPgVhjfzRNGeKh
0uQ8auhgQO5/N118ZZuYQI1UDHSTRNKNdcpMQyYIB0LBxHrYU0SUtOmp4K8I0Ucg
lYmi+VlQrtiJ2KbKYrBclDDJl2uBJVol/nscwUZntukAZHn2MXphr9UJqKgbXDcf
7iqUoLeN4vuJKA3wH1N6J/ao5Ogq+UbTl8W6b+NX+zPlR4Jo8zSQzVnvY1rfVqI+
bgLvulnOCBTBHHN5v/jIo9RfbY5oHEqWg19TOgy6jGvmu7j4NAEHxt3GIyXVmO/D
3YOTf5GZtpt0jUX5p5ChtZ2jvvai2pQZ5EgGf1CQL3LLrsKZgbDrs7/kyO739ka8
fUhnkhyCghfB5xYqO86tNHSt7UHfeI7or479XIyyxrBoJjWFiTlEsEt/7J3REYvF
9QSXeBU/W0I3PrtNK8lROZFmaq87z3BMds7VaWkzZQdS0kvHpw+p+bMEyVpEBN/9
PG6tYcZXlvw1JgXmsufzLcLc+KA3JbAwM8gYxIPhBVik3eBkfphMYkVlwmHJwVs+
pjcF6qxdP/vCUCY8z9at4kIAW0c7y53WrjRefcN4IqH5gZqbF4WvLOrCpatdRKxU
KzUPEt/zCUGExBEtuL2r754ehbJcGeCqvMOUbnBZmE9tbjtdIVib7mlirrwS2wcy
duvF4KPRQSEal2DjDCUfGKkIh3Bm474q8e6v4DCI+DDQ9j4UxccRCAaP6kkJ92LW
gVO8BV6Lm2MX9K/n3i/2DJZVlgGUfQdAJhwm+cO2VzifHVOS0CnMRfdDB7V5hTA9
pWTT9mkR32h1ePsRw/9ngq6+LGpJ11IR9AVQnY50WrhGU5YJnRTWBa97Ii2d1YvQ
e9JLo+n465humg2eoUIKyWJWRUCR9JZ0x+HuLR6ajsL/gkSGXc6+JxDslx13/Ze6
px5EkEaMSupacvRPTEippaoXOHLWqGTl9W767PJIZ/YrbtPARRn5LjlR4cZ8YTUk
0rETP8xIyiHDKiVLNR13Dt5Q84wzDhtZM/A5p1GE/+i5h+4Q1+WEPpm1l/kOcRiY
XwPc5UBL49vueX0+5/L04657O3cIDKq3sUMwXxQDTzP6kumybylAA7BXGFa8mNjW
fQvDBmS1dnjQgkVL3LSJmUg0Muh8juK8xqhHDbRz6cnX+z6kLMJlWx5l2EkggACY
ZI/vY3cCPyHOKfDH+hEFrjKT2NCm3YhFe3Pl4QQnCEanhGxMvvelJlGBHHVSDzLp
46L03YCPk7IVm+VSz3PUSag8iBWUg5E+5ieEtxGj6XavauaFot4VQEmhb2l+jgAM
WEoAW2QPy47LbGVcorV2NJl0fWTY/z/7ShdljjvI1tyaJx7BOxOcD9v4N5ZfvpxB
cVKznUQ+HRyWD3XrM0W+oSbN2mVL7dtwSNNQBBLuR4/NmHZaxKhE2NPlG9x/RO+W
GvN+z5YGUlqPWZfm8ax4TRDEHOc6HbFj0r3RxIb+Zc9cgJeSaPS3VANBujRWCIr8
VZ2n0oTG1Y0E7+RpCPLl/MwTs3r3T+X7nSh/5VfRbFpCI3dR1WpR4XaDlHNP7w7Q
5gQ+MkH/4vDxB15DmjeNAS0AUQpBb7EUNEr1s0lCEcda1PslO/zvdw270qP2iJDR
lNjRXvmrIkw5TpJJ0zyXv7FF/cLXjPcphyRk8JSO1j9/meOf1Jo8HkODY4aZ3xX1
beOIoyXEQEzsRszoMKTNNuhtjjCkzRkket+sgDKhzEQJkz9g75U4MfOR1ngLTgrE
HE8iA8jeTGmwhbqjUZAqQcYYa1RVfhzHUL/c9TkNHPMo596SpN1uiZrv0ezED8vN
ecUYbXswFMDU+AoHfCaaf5WB+vsxadpkr36L1YOhftbbUbKkXWYXINdvgd+PvJUp
EyIfbeUsf+A38zpKEAztYlc7qvHyEBr70JIEraVcUjgmyL+VRri68hnFJAus33lY
1naEhdDawvEjbXomRu+iNbSHnf+aXBkKFFEdp4mtaqOgvM7QMv6Gqs2x/pr7BhjD
4eHhoCiVWZhSDvVsZ0B6Zp9srANyu15BHnaAp3v0FGWyyIgMOhghqNRKCITrsTyR
zQOzAD2apkVBgCCpMr8Gs+unskoZu02Dj0j8dZAn7UauUJR7lyO0Pwawo7U6FmE0
feSzjfC077C3X27g037YIPoYty+Hd7MN/M0kgsvxP3lkPHJYzWREevgnqOQ9qjvQ
mFFIOSr4trwPTIcd8mLTnEX+sIWCINUbr8BDIdBqdb+RcBC8CC5fBtcuvM+G58Yj
a6L17B6rE9jXVm21yT8Fn0Ez3LSyINYmsRmI5WXpFSl/RzNQxwrNKXHWERm745ov
hgBL7O9KlshyObnfqV+XNCShEfi46Z+RdI/jOXdoODnXJvk57SV76059VzYzT0gy
i5HPLfBJ7sa/xEHud1hcNWymQfedeWI3Ro6uqaqKXcA33oNRgU5F5oTocPMO0tjl
6v8vPRh0ZOhv+j/JoqPLnzOEYB3UCBUHkJxNx9vpeoc+XUVSr1U+dzm9pkhOMIQB
6VoTyd3ueosCG0PLIV2nFVsI+ZL7xzvqv7IChPsGbU+yfsmNGlvhB7CFZA4T9uYL
erqGucis4yVRU4tVTgMgIWe1VeJRs6+jtHQbI5H1T8WL5+YiQszXzRwSv7G5VHuC
xI8dvg6bOxVdyFfA4BZI60tyECpLsalJ5MzohcKb87iQG9JYg7Dwnt42m963iY4U
oENxqZG+gyhdp5Sn86UQJJmTyLYJ58yVF3dcvTcXGI7kmclLbe7au1CSsuVOcZxM
/Fsyv0r9DGJGLw5v80bPvkcTueTNdPNixvANVZsaX+yjJRKFJpt5vbhZtq5/8a9J
2w/uptSpWS/ZtUPAcdyP5B4mdzXD2JDWScl5zpOd7cm1JdGP9hzf4cbVYK4Kj0u+
IR9zpp4f9w0swv9lAhxvR3CxgNy4Rd3t9BuCsX6tilDG8eN0Ud6Bg4Vd46cXwBmN
Je5hgB20Mx2OxHMrkyDM2VZ4V7I1XRyRf5z+6s+XmMtC/cFqKf+6DxTwswcys9So
zEH+/B68PKhnxJ2f2P4/z+3FJdE1QFHnABfSCiay1ZCWT2VPIcxH4t6MdksI0l/Z
k8wca+s5QA4IOm7rH80tKh/vTVjzhAvjaVAXvsioOVPw0BpSetHa5GA9MkepBo60
R85rQ2dZWqbHc5HyuriiiMPMzI8FTXQOp0iSwFEAX304pQ8y1zv+h0CS52JN2iW2
S2NbwTufA52FyUbmn105ZTY5fWvyB+g2HUzXM7IDvkY9MrCisMIfrrFZlsUfiecG
z99HqgNB4plOUJ0bVksg754q2Olr2+aJa9mdY3t+qQAewS8uPAlC0nie3XEZaArS
gT/XwAuLd6MkzK0zjoZcQTuxrlUA8Iis7nUElrkILKktuAp8PjWagWUYMvCXB4Kb
hFm5pvlI+dr+kws4sqI5KQZo3V83yl4P7lQdO4Op9naw88ZDGVShhpgfeSCSCm8k
nYCvlB3C40TP9W9hyzbxu4IMasPVv8LjSjXbros8x2dZJVzmCE7CHE0mvcJULnzw
TnhSCWd1BfZxM8BUQBFhWPpgJNTpfbBosgSUv0ZLbscMfSMIZknTvTkzr5K661rp
auCxh1qBWT2qCqO2wBvFXQcXPyXG8NLr/Eeq7eKuOofQXlQnxiEYtMyYNMJQRz3m
uomBfLj80IjpOztON2FB/MZpXfgxThBGJp2BcDvj5HRUqHRJcn6/RoV6R9f+eJc9
UOr0vd6Ps9YNmnHoc08aHOIeyJeGON4/mIZstRV57Yu8AhH3RdgVMs5Wz1+X9Q/d
WcOFH3M8vnzAPcmdULbQu3PcCdbu7Na4tz6jzNkI/e4FLfZ1OHY0RQ+soegmsOrt
P6a9A3+3uunDnHukymzzpV6zrorf+RygqNcoVK76+x/851xC0UAwxakRe3ieVrnM
otDeeZU/ENdq2oTvn9isPs+JuRg7dHOW5QqoT3JDSARQTeTfJHljgDl08qWr9AzZ
l3l8PZpGH2fvLmR7s0ugwkn+eq9bZdQSQZYNZ+2e3t+ssfY9IPFd7cTRpylqAvMz
XLUHRj3cvvMw3zll2fLuyYzAOsA/HuopF7g0oERxtKPtclK36CKcfyTCKUss2NpR
2pLYtGZP0Iy/2dMR+S6VcEbic+6t1FGL+r5zupdtx9tQD0efKYzPR+3XYEANBoM+
p+x1kz435g949ii3A3f7tucxoBJkUhbLfnL4G4vNVy4MqWQKROQBoWMHVwI85bME
ZU7GhRZBXmz+esXfmmC1WSIOca+GlHkVO93IHVQGtDy5z6oSSCCNhShoMhFcZ1c+
mUcc9jOzQhY9QNBxhFaial8954WMTKULnn957vIi4JxKXoDT4+j/0Wqf+xu476t5
kqzxJwEMA/QswFdp0jsmW26lknNzDYM47tdLuOXXlL0ON4mkNKPsBdS4oL3v/+xS
ibMiYVNGJkgDDyzWidEqFFEmnazr2r0s+mWXTWB3lAse+r2Ap3S4mFw79P6ZaVck
1J73LJgxxDkQeeWZjduOPO5NnzPYGfCD4GVOZXQCkXJGBqveAC3KzpgxBpnd2b8m
7su84dsfJRfaGGJ13HZRx86WSlhwAyQ08Le7l6Ih3qUnslJtJymYi7+RK3mF//wV
v2iRwG02V1oDDXLfG7rz6Z7IJKmdHz8wZv58o7lRi2XHXxPsF7piXl1JSRYWpqig
Y7Lg8FWHrwjueGYRUtZuH2AfmjjBrYq8h6X3xDrNXhop4FpwG+IuPt9Hfjy3OWp7
aOMIR7gXdMl2ERRvEkPPgqf1oX29Wc+RGEH6FG+n/J9GICWMODGGJMs/r0aCOvmG
NB8nuo5snR6qUPWSDmZiPqWxg5IBB16zl6otIysH41M0iZwJKXsedvRgmD7AhfoO
nvWOh8oehav1jgj8x/XxsPv05yAfqzEeLImuETCXirsPDR5Q+CA10L/5drmf+959
iY5cu7Esqo0fL2hEmRyZP2S/E8GHsk6v8W7dWyVuQwuHaD3IPRnle5d0dvbnB5yE
dGIlX726YSZr0+VHh0E7A9FKNxGXbAiJ0jiLr+7INjwxbzFshVteRoaLupqX7FbR
kb9t3oSqFOj10M8N4FvfdcnXjApRH38I48uM4vSS3q28vBizk2izlVqrj9Sv0dNB
dvChu8U7Rgc9Y1UHKvoxgeUziqrfnaruy3DaBn5C2TymKZYxYBmwImdcXx1PhSGg
rgy+72UbQwV112r5YMR8+m01LbXXgn3rvy+71Y8KeqeEAqCrLDXUWomjpLbBGV9x
0ULJ4FFPDwTK+CaCdme2QqI5SUZ0DHVjThi4uQO17iJ/bRG3FA+1/9sVFP1Jpa2z
xSuhdh5FQtacvD7s05iM3L3sAMqKTDR39DJmoneoFwWPWsoJ7nOo0P2rQJFVZlPj
eGCIihdOdVaGn8+BxzuYpfHjoWsJro0FQZJprJzpshc1wdTJtR4N2Y4p9zLMk3Cb
dVTh3zaTS/RQnrT95v3iEzvPCkGgW4zspY+xI+1CdGbXwUOYiC9eUvK+xsXj1sLH
nOryKGBxAOqZGITYW9HND+xVroO9Q4h1wWzRu1eKWcH+C5RoLsulBQlPxU298ILz
+0TXrFgPHNi6w1r1kkhcpIqWyZOEl9iLnOfj0a58LftHSPw8xakQgMwCKXGM2Pnp
SbVBRWFRcRUHeM3tFgcYFjcbTZkvk5QcOVIiXAS80wfPMrfVOz1rCWhcJhDDwQQh
bzI/TggnNjdUNuBps6kdL4yHzaChGzQ0rtD4FWEAymFoqRW4jFmtdszCXPvE/sVX
zssdjWvy8ySoxT4sXeybwnB5sxTp0nibJ6XiaElvSa9n/1FMEyB7xF/DgBcVgSK7
5yvw8oMTq60SOeGRbEIi49hJ8qhxQkUhrbddyGEPB1GtKnOauLSnT51nhulNHRuL
KApDfqlXk7YR01sb2GXJq1QMFaUGECu5bxohy+KOIRfPT6Fzql5ojx9Q2gvoPS++
QiRFI1HJZQInxLNIYvAaLRs/iHZYAs4+G1L3OFdHP566Wrgeuz9Mw50So7sanYjC
Mn8fuxB22hIOPNA+oy6NQx5WDb+7VqV3bL7/FxdULLZkXua28dB12IoC8s/EV3Vd
CtHF17JgRiip9uQDPiijqHwvRZboRP/eWtBO/iZtkdH0FfKqUYGiuu59hqQP0NP4
LlSIh7U/VZyHvnwUf4H+ibA0Vu+anM4/yw6/oykVFvmK5KphNeRjBR5VeR3HTU5m
T3qZVAmQ+Je85upIbGfYw2pU1Rq4a3VfFoSCb3IMsoJeYw1HkypvciLfW8Hy08nR
YqoK8lW8L6HngZC6cFrroDSVBR6vnA8QIugcIiPSnBLjQFFI9zv1rA5NOL6enPY9
mEk5SJZHE1XJyK5mF43wiuygIy8rSKX6PMVd0AExNuLV0o38ljiyvB7e0r7TJiH1
bA+8IITxfglSIYavnRbhiHuOFmg+5H6TGDlM0c2pvzbm/LeuVh9J+0vAa0P13Jc7
KILB1V5fhm7XBtkY4ZgiOoH3jLt5v++J4CtxFJZuoYx+SHL6ev4ZRXKZVAOqp3lv
1KmJrAYg6B4Lomw8OSPyHmEbkPFB1IWvpnWs4iQRmE16lmZ5NqI+cb3ZS8/e9RHx
fb6aknaAUE12+fY3WEN5/SbFWNUMlkzRYw1RNlzCnFSms+mvDJEjxJVW9qsoirp+
bYpizpekGPXzfVRofMpYVOP9t4FVIMyJI9hdc5XpHhKfOYGKyIACJdYGjPc/jkKM
gPqVWDmKN7MQ3RhV9rQXwN93qMDpLvakh7S7ebSAhpmwefZp0me7Zs8IrNWhS75u
SAAJ8xESKLW8FfQ0wLOL0DvQXKpDostkKOFQtBTE7cGRCYHOa1e+fWxvSLUJAmT5
ifFbc5E8qa2Dd9pqC883jtfsF03e+g3lEUIG/NDd/IrVr4ru9DPwsa12uG/UIUWl
pwqIGX4CmBhA7DNjEf3FKN010Gf/9Jcze5oORoA1CEmn+v1mQaVpYZSaMXuHz12h
8ldpoURpw90+lKFiquW53qBlcWTv/kS3+E9i5amh42rz/E8m4nDMGaaxUCR4i/1i
P2CA/JIO12vj3UtDHIVyhjGhyM7Gylxh4EJTxz379925scVzyEpKD5FqGrUFdpM/
c4WNAQtmsq+R4HTTi6ew81TX0k/E7NN7DuF7KEboErQmSPsXp5SeTVl9jtXarE0l
SYoX/66K5AvHMyGWLZn1fIcANgZeX7v60mKiLuETgzvu8+TOrUGCufM1H58/sVot
hUplFsZ7PvgWJChMIJAHiNQu8Hyq0GHxC2iAC0DxqCo066zfz+56eGz7++C6PvkI
0D0sj+7oYy//15wHFpofiEatPPbEGyZ1rr4e21oj4N28N/56BQ7NhoRlVKvbhe0F
RqI6doOEG6XRNU9L1GuV3NBxYYsee5Cv3ycDUSV02a+KSwunF0PeZV1U+mdF2A9K
zYrin2TEKdT0tA5usfmZhxf6rAuHNzOEOeaRN1i0tWpYb/0F/cbDfBTethCLpBnX
Qwv0+sC2I94iBqF0f5X662XrCrjqI6HVjQIWqPT4e6cp8XeLxhoymeurNkjMuyVB
jdrThWM0Vz4PtgDAlNCL86066xhsiBSL94m5RPIv+vOojv3d7DUFzQqDO+vy1t8K
04OO8elC3CRTeQ7UspKUX8XYB0ofG7NI/cXZG9LE1ABcA2266gKsym09BhLk7Aob
wTdLLoK64CnSoY1zLf4A/n3ETIfHzzSwSmN0CgJbA+n/J3lBd+iiTTUiRRFekzwj
iOF2nrSyUvYIpDvXq4uv2xKyEd2KUrTO4J8JJp2pMaRDPnuT00fCjBN82ntL0Xdt
Iz4g6lf5rMbjEBWLQFeti/HfkGUs2e3qt5FwRq5eW7iwlt0UhDEKvhRXFhPC9U9b
tbJB3ckr8A2a4arJyeF/2RTGfevu117UHL/zx5ubPyuAHl3bpGzeiX4GQnX7rLyO
xzJGMGyFu7qqPwdQwUwqmBS2KRw7+9cqkpldHoe1jYjQY4BWCHDDPJy6g7kQnr5X
VVDvW1gNJGAexVF0kds6mz8ZbwhnUpmT+s1YYx7Jf+B6mbn5fRLaK2DbsH7rTuM7
70xwn2HUfPmHAtwYXjvhfVhhM0/oYRdW6lLqsoX0yFybJiu8ouhnfUnerVvCieoo
aSuOAJC6A+8VxO8g3f4Vsj3mtAPQxD9/hpshn4AhmSgwHQ7/IIl+x8XD7/Sl8xth
2GNuS3MNDTdiJGUIxzDL+pLlPIbNmDrm2nia8wmLQxj3T6BPwnkXNuNOwwZwwj6F
S4j3Z6o/HDQeXGEme92upo2EABK2qAdOI69/pXOrH+b+kSQzU89ZMYdGl9cycsNb
qDn0lmgauMP0fh5b9VFaT7WfD5QFEGzWd+IYc1XQ9HJC3DHh31HV0VO68HHm9bW5
1ycUvSeRadVd+NWXHuE/gtcsoczhvdB7SL/MRjyeKKtP5iU7Mc7vOV8bl8XApmn0
c6t8XujyNkWVXCo+IaIc51nyqu0CEfB7GEGF0LGzqUpMcNB6KImXMIrZJ/bwu7BA
QQtK3mP7BwN9zUrzT90l/U8e2ODm7huk5dLgesEZhui5/eBo1SLmLZ7PlfJpcc/f
eHuFE/WyxSbWcSJGcNForPHAhRMT6VnijChK3rbTy5gX1nqGFdPHvoN6McXYaww1
hcgddIyupDxx1qAE/rCqLtvQO4EDzF0qnz/qmFKAzYTdQ8z0dsPeIWaUy620JQ3D
OR17ieg5fTzObBmlxocO59yBTrhlTgXmdEF3y344Gz8d5qk56dqawSmfvSGzz77K
04vbjIgRS3Ngl/ZC5Ay4gql46p/6BuRNro4jWBj47xbEH74aMn04KsdqJ7cUtcQP
J0wDLAhprcA2ewq0xOuhtiPNnGvCkXji4CpOkbZYYQX0K8Sr6S6tC5fxxwmlcKt2
n9ZUwq/MT9GJSOMNRPHYnXfq9zwI4D8Qr1zndmo66FewYEFkZe1OgBAJjuRiw3qJ
7JQs7NBOeRNpf8pB4Xnrf98kvtq+N36lHFGxFmrJXbI3mXMMzL5SZFu956vM2fKB
yh6HL3ikL/bkIZ8oR+zbw6pdccgIlIoLcac024mIEKMMTXGlyh+f9cTWX+okCVRB
CAR9izqdfpALvVEL7Q2GT1fO5PpftBNjEljS6k7ESSquyutLx1EUe0HNpumYdJVm
nVSWPeTvQY24PpM8sPim5tpcXnP3KMdrHdN1/tuME/cySoyY4TimGbjBUurmOAwq
Uu/6WLmsu8krMPso6MjscsMvffDDAuDzQ7PQa72I+FoLuGA9oSIw8x8C4KKSf2rd
Ieja6eWz6vicGHF4sTfp35vUWkd3gMjIUvkk7TXCxpSGzW4MW4qUzVHr6JFFF1jV
a3VZ9QnbQjAjUqcmMg7iGZGiYhifTYTnFtwQdgBUFV6TmqrZ3R1v5BCejAOeTd71
srbxgjGvP2OyTGp4cfTUruaiROW6qhHYN3DYLJGfO14eOc3jccDVLhVCBuIOEShR
k8W0JG9mYwntB3oNfcagUIhynXuBaDsXVEtN12IHOGXObn/5cUakBTRFEIhEIT03
Zx0n0EQkMZ5XyWAgFDFd76u8Xg2R8muTbCbwmyiH6GIJ0YSvZ5T70SWZOSoilA40
/Zfj9RlOmvuapQ6hoqUBHLXyOGQyAfh3HOy5sLI0RRpw2lGBEigxJx1GaYNQIN0l
NUyMt855T7kxwkoObbSlF/ZzIDEvJyUsuQixVYNIQv/jZ+GiMbhZ4CE1aRDUIfiJ
LuVgoVYpwMIb2SPErbxHnKLIugcpJSGXECDZ03fGW18sIGaEGKIFug+QIVAi77QN
eZi8hb9iekp6NijPxQzrLJxaUoGIGuEB1TdBfVKCe25nVJhyW1WrV6udKDT8bL7q
zhaG3Ml3JGJvG5dX5OtWE+1q3kgcScUeGX109uXrZonr6UTCc40l1LV9cHNn4rLf
U6/XOlLWbbkw0FZXgM8odCQQLMCtIeVHM88yr9Oeke//QJbbO0EkvAtt6n5blcYl
aXtRFnyXGgl+PvBgkMrAcMwDlz227Y4mN9rZRyZEEQbwPVeZVN9W0AJyP6qgi4be
mEih/RCOonnC5tMF/5Pg+5wEJfVCHjAAM68aimlKVglltfipXnuVRXX/vHILIhr4
F9muUxmDchMDkMw06zW/414dMg2sBjk1CEWULMKZ+nvKaepxc8VuLni9OIR2FrjF
Y2Ub5JzKbChiPAu3xkPckibg2jtTv4UfEkO1OP7VJY4Ym5sp82eQpnbiGVEnihnO
p7LWy+QbpiRtobFYe9QBN2Zj698FrqtQny1Rcz2u4vpusnUbgs2Qcx2RF7NerSbw
HHp3fq5rwqT7X9XhEL7TRrQFHEaea61u75Eno+qwKfdR1rnwkmwi/mIbj4BfaPYt
EAaxbMmFgjHwNfV+33mEWHGVDOQ6h3HmYqTbWJn2HErThEXntn5pI4pTzpjJOmog
JkA7FZH+HAwkxMrf5BHyLhYLuctUUet1J0NW7i5RkF5k8U49jxl4RFhlcKmDXeSk
AsMma8fgYYNnk1mAIpv1W5QeqP4EPogXlDlHFDX4AtkayUEAEzdHIo/hx+MGm8nP
/WsHWcwhtRHx4JMe0mB0ahcJxHKPL6NCoMJNcFg5fXZCeawaXCPzHZ0w5g4t6tHP
DOoe+7k0y62Izk43DZ/scf5xQtISfP8OMxZKCBFT/OJmJFah65uBrLKESoqtvoCe
NcChKWpzmacn64HN46iK5IGiA8ZKkLFxxCc70e2xALMkPpeygh6O1ax51WoSxhNl
uDPLcqpM5ClvDRfIjWbKZh2W7/lZbtH1sxhKVxQYfMm8KGyBoGV83Lkc2C6i3JYu
oE8D7sWqDVBufitxM42cyoeeHhw40ndKskxzO/ZxxN5atuSYsYbzDGWbGBFWKZ12
YCSeV6FvcW6J+PGDya8fxbNY0SftII4hXiypxaqd2FR6LXDaQClTWj56OgAbd6Bk
Cyhhizvjb2D3SCa3g4gWjWeuedS9CNRXZAnwSfz+HILOzhae83EXH2ps/wEpM25l
fUgVWay98KjWam4+xwQbhvHhrtP5pS/OvZq/PvgpKGKvIZohTy6fR+G5I2ynU24Y
UduMJgSdYCWCuzc+Nxae/0ZFxTxpyTv9tCNGUrvl1Rg5RkT+kdHLScKTMWrG445A
d5Ove5gtin8G4tm0SUv8mqsMby0Gd3I3qXtsxGg5EfqQAqvorDK5S8WRl3GW7Nmh
2gw2n/rrLCWepbBl/OEOela7tplvm4+eVAymi6L49KUw1o1xkmv1kfN9bFlCNeyU
frubTurJqv15avgCGzxLNkoER166n8tcwIWwFkfTa26H53FbviyUNhYTLLuTIoHF
RYiwUuQXU9s5QNEwNBpKosz3Z8wy3dTWAvplWDRhhXu1ZLaiMywIa+qL/3dK/8CK
+BqwUNq9LPA436TXAln3pupEC7rF4zmSH+macCMczBkwSiZJSLEunJhYuXWAT3tP
bnP286jaBlj+apXWAipKFVCqr6rwQT6Y+kYj1s+GIlkAX5OOSNFzUTEehvPYMsf5
tUkGnA4/J4w/WfTkBWFLKlMA1dvLmsAFqF+K2r8/7kqSNuRXXs2P5Voomn7LuEnT
sbi+c5Y4BVLG2/89A+KwlKxK/XBdkvDfWfUsY1TrbDnLH6+rCCQpua88vcc4bmjp
gzB0Jwr2jO3r/jFQRPN4wy3qYvUAosCZ3qNVvPnYtJPbBTl4KUA6n9Phy9jhcYPe
jXH+fN3fp7U3pIDfx6Zx+6RjYa5FsE+RiOETi5kIa/t/ioYUm6sktXjF9M4m62++
oO39p4Ojd9OT2KGibciZQgzFowRGrHenMt/qymIaaZ6ykRzUbTsXYP8LGMDQdycN
9f1/N6+kjHlE9ls8H6qvOupsM4Ei7q+py2mRgTqUBFOAY7dBagIrml3UZsviKAUk
0biO5Cv+Xyj3seE3p3IjiuKTYzeLVuSwKAPOeIZozVtOJ1uqoHx5un2vD3G2fGdx
fhUx0oxtMy/HDltRXm1lC3KxYbxkFNGAQ0NoAn/nD+U+GpbATxd8jbxpMTPYsj3m
CXdWyLmz7LSplkq+8xGan9ODZlEeiQkHYA3/8g7q8bHgWLmDJqV2j6/GEZIqksVZ
BK7Js+SXHNKfSwxJ1wYGZkEjx6VBasDiWQumA+cp2D9laX0JxLFxStg4yNJPAGSV
5FFLRpoqd/XBj+wqxjBZUOnEmj3MPI4nywsU98XSXYgJl/0nVZyr5iG2XPR0uVSJ
OBpRKO2dTNbpJY+ACSx5ExgwkCGoenYxB4f8a7e7gQxQ0YJqTBGFDC7CAQzgCkgx
GTWnbkuVBSIh7e4AufPWI+4ifXt+2MSXeZAT3yZs4HH0ujJEEPsDmDkEeW2cX9il
llio7VfzZGhUyD3S3/asTVuLfWwKZF7OOPh38Z2NKJj5ma0ZVQcG4u5U/4j/ww6d
iNFGnL0yDIkuWrpPll4rnHvHqdd3cPJLn4wZFEgs3KDNwkrn9FXnYVM9/V6UI2a5
cc50J1Pw0dszq7RFOOyzSs1sMnV6HAuUIsWe9DuYOQagmP0AD2QF/8Wm0Cq4yFvM
QXZvw47F+YnWyl2zOBZr5BCZ3rTlzp4lBd4D1RxYOUrQXSzRgfuC3+ucYy3uwmqT
Qh/1zgMEMg3luzLgiqOC4zR3MnKBweaduf8mONQyid8oJpaRxTLbpdlVq1QLLD+k
o5Aw966TBgB1fCXr/49PDY3qh0CsLGaRXdXs6NpeFQDmDgAJnZqW7NVcjc0MlrO0
QdbPazfQu6s+GS4X5DL9wpF96WqzosO83R+tlhRGiMVUov9mgbdB0FZHn0OLXKnx
ZR7dAvosRTJRs7QZgJuGBWJtykRtXbrMzXpNGwcHT5+6/6f9x/1JjPgpnyVQA/ua
v4LZ8beqPCKtuZVgC5sXlTJ3oV9v9vKbz5ITqFnKBPMfyUBxTWfJIhgvejjQ/VWR
FuiC+92186vUS6lLhHi/goeEUccisq2KjIAEMFafxMHmowCtumJr9TcPAuvuLllt
kSTiVVOhd0sgP0sUu3YoVwmq08XRrYpba/ce2+G0MD5IeZGrkNqTHrmtUtxkaKQG
Eog4+NQHIBDcB/dnN7xHQ9+rJMN18sL8FPCElo0yfe13cPri3EETDbBD+tt4CqxY
h35XzGsrQRmsjh2mfL6V7FTr15AtkVbv2grxVZjPt2tz339bY7d6qvFoJhIVstUA
4mmrf5hDPjTT5owek10AQEjx2gOtL00mU3EmcA3yb7ltYBOvlcM3xjyTNNkiqVfL
4KQTfvck9cEpyw4Z3qyy2ilRyU8BzIzTdGHgNb1tF5O6EOlMqM5F4jcB7vAdVB+f
ZKIYBSWXWknGdgOAtKJxU+rAIFNPih7RhnBDbhpZDD+YT0guShmLvdh/D4/5+sXI
5Lhr4QuNuCaObEmFPRhlQB8Ym9+YhUmtWlxqo9z/EQDd13qvwqHpiXXqCb+P/e0Q
3Oxlzf3M2eSvKRL1US9N3D4SAvEwEjZcZXQ9sMeTVdmy+RWF+3utaYVF2nfdqLWo
TGVp7QHA5MfQwGZKdf3dBTqXEoLQ9OTYMwuf5O/+5B2wWAoKjRxjXLSXEcZKB3kI
k1r1N2fvVGZhYsfSC5ExGSfz0DOyoMdpZCyNYEtlKYxsr50whzg2HjBviCpufVI4
aN/2CTx9Qkd/nUi8AxR5GLQaVJR6VRPpjgMplPZVFgevqKnavk2uzBc2ArWkXE16
7jwOoXMTIelFK7Xg+eWLh0sKohipyAbSWxwyo3JkpPvjFXYHyQgEJ7QJx53uH8y9
wFiCWwXGxO8DPmBBVQMmPttz62GFWgr7D8bhhTkdHjsDJD58ok9sKio2PBNyo/+R
Q2F9ux3Mv07YYLPX3Fg9HkOdDJ6C/w8BWLUybg4hTnJxdRBsP65Fnn1+ec7DH5DR
mYrD8qGY1MhUdTY7No+aNkfTnqQ7U3+oaxrlWHlOXeqf2gWqpL62GHt1xLILHRMX
3XBEuFSqwH47kzzrDL0OqAYMMRp0ACL4MK5DprJhvc/ljtZatS6DxxYk5sJzkXgn
tdHMUNxL28ouM2JU5Dsv/OIuOGM7lzr8bqDCJhbgDxwKtwc9+wQDZ5lqEigsWdWU
9ALRBDGk2+WRzqbbJTFcal+nJml++jX7KffU+hcaDYxGMYDHQxtuh7i6FBiYr089
zClvfATiodvZUg0y9fpexCMeIrOyGr+Lyl36y3b/vLiP2Xf+am/NGoOBkbzTFJqQ
TTG7F9wNNxdM1pxk/Vwoo3d5cCHmYFwf6ep8vwd5wJRk4VVdheLxLY4UZKlujLdv
8qk1HMoOKkPuRU95WWiUVODn3edCcpxQ4rFGPqRXUjctmnhnrq0KCrmNX4+bCIOA
GRL6gHCj8+kj0d/yTiQ+W3hXFIWBOce086FMjKzwkV9Pv2TCv0T0sSHEzDpw/LQ4
KUYLrBMW+Cm9KO3QLotX+irP3jV46GHOLoz7rXgAF4VFlzSfTy0k64gS1221TUwk
lL3jv5jThjw8eN99M/aijfSCre/YN+3n5PqvbwDdBS3TXexLO8C7U2fexhk1W2Bi
dxameK2SBn4Isou5cBSt5et9hw//pE2OmvXiCoDHFLSBTn0k/wBjobt34t1wOUht
tXyCMtc+EJtFAnYTwupUn/C2YmenqmUf5RAhrmmI9W0G+6a3PpY/oHbuFVl7DKdn
whrNxaoR6pHL4IQsMIo+s+jSZMw+pYM9xbC+I3u/ps9YCRhB6Lc2D0Sf/ueFHzWh
RL+EcjotJ8QLjBzPeF5JamcQpxDEk/3fIOnxG7+s94vzf1vTCuBhx0WOgpE8pEI9
/6wzUqaaj9XTW1yYUhKLbZPZLhFHYB8qgGI2qqEDuPuTIHyJcc80Q+81YMzbxx7E
PgkwNFH5NFXzDJCX78n1gxcvCyBz4uxcM5s6KqhigiRc7Jqx4zGGwzjEvh3p4h4L
/snWDHYL/Wzv1jhIZC11QvzFtyhjN91uDeLWMV5AP0qCWdErIXZQUkGK0r2TEsyq
dTB/NQ+L8uxW0R2L2RoJ7ebwBHsemyXPQdfPzcSaXeZXA8ZP+m3YSP18d9TE13PO
nRa863KpPreOLsEfPMEG+prlSX2vg+jogVzgTaJuJXf2Pvu+OmoVScFvVUKXw7pn
gYuxsvu+BiHDEGD85JYJXWBW1Xez21wENvwNzrYlREeibkFEGUSNNCDHpEexsu1/
AVKRWt0FVxgTM8kUAgVmcHJTgXP63ZVB/Q7I03/0ZszPogPN7Uly74wLE1VtYqmX
g5Yx4FL2c9ltfrPDAkZjtrvyTJV7fTrlV6NpV8vsucafVkTOYYIiuRRCfZfPHhcl
ymBIbhfi0U53h3D/g5oxad79TRe8DLXNeTSJowvRqLKaewlTzIIU9kJ0mRqzoKsY
R1h2zWpAhgfNngYorViuYXLDcLKPpni3gvxwBiEbjgRz9VLxssBUztyW6gqrILPT
Pu20HtZALtqTHELsXL/KBxxXCScmL6d36TDfsnOPlr70yjBlsXqv7ECZpsUqdet8
tRLiqMTIiJTIDAlDn6dYOSSpXYg3EgukbKOKNdlPrkb9IYW6WceaaGTn1zvu1eKm
+GZxGv3XAnqYr2LrRMQbeuEMpd81JwI+FGW5qGhL/xS4NkA2P69HhBv8t5hExSbD
DxMAI4DHhjuh7fgcM+5ftwQtHn71AxZQQwnn9KWY9EjjgEOnoneeEt7+tpoqgBAq
4ZHpBNr9+bu1UWs0RYN5moO1/1zx6+ez1olNZRjzjmB7sIX/KEPfz0xW5YkoW3d2
/2N1cQCKQEw0UdeSPTHKVyL3PRfFMFRGQIsgcYQvkJW1RRhk0S1XhcEqQ2bH6TQo
HBw184xvQSSLX6jdm4zcznNiRLnBbEpuAaKNu72xvPx+3V8PvbB74l1kMxN7AL6p
7OvF2NIQ1/XPl6qZr22qW9ZYNTiBtRqJrVe9zdVpnAOqoN3MrwGC/8BkeRgmDRPS
Q/SVp+u8rAZj/VY8XAgjIJtA04jfGvB5KVUEUnIf4v0BVG0bxjjK7fZtbJUm1QP3
XvI6otdA5sNapA9Kepnk+7Htp/JUwdqQyma96Mw1wh3SI03f7pafRn5lc1buBrK3
MbCeX0UnDRqGvWe/jp53DjLfLJmJFjZWi47/TfbBnQxOtjNfjVls01lKG3YBH2i2
qk3fQYr5+bhXJ2glzzwybWYChJPL44Lq7CMLvA4xiJfn5k/TQwzfcW0vD7Ga/70c
yaubOvYhZfO29dRbhOS1uSx7URV9n6ZZyH6nmQz0sJFXljUxzqyWjRk6euEcIaUr
dduyvN21UWCV5GoJK+YPBHbTH66c2+SWRnpT/F7/ek5BIkYWSoGzDTwIF6aNXNxL
6jG5LAVrSSn/RTuP2RHzWlEIJIyjGGJ3xslQi/fID08tUeUnOmHz9XpN0zs8Jdy0
tV9AhJL4tk0CNDvr7amUvOb/J4PVLlgqdUGxzrnsiH0q5iuqcLskNyMCNnnIORAW
3Ur6KeErCAbxpBEgs56I/GDp4bEnVMZOA6fSPUexPKwiQz7Kg8Ki4AYHEWrjJAuf
0cnDqTEEnMva+uo+G02Vc/7ktY3aLOTO0W7+BNPttkugtH5Pjp1X/fI0iCIgRDKH
InLmNgiIJfIsM8vMxjiyJU0G/NPjo/vw0RecauZ+tqdhetLxpGwLXf1oIfk3v55N
sDJCErsHeycw10pPnFcoxA8kEC/0dli2iywtOPUdPH/Nx9taZ5L0yt0+1MgjCqI/
/njXqfmq48dJ0dYQOwaBeL85DgyKl3uaDL7ArJmDm7dUA30VWc9nU+8gIMQn5uuH
/0k+64SUtcXUz9BAa37JIJJdhzJ8IcVbE7tC4GOmj+Twsl2sR6bwPl2OWZF+iP3T
yTtLySH/Pu+0wActrsOyEnOW0eIEvPxrpOmPCF0i40m3zieai99srBVT3D/FtZUp
B7HMAxfQqMC/zMqTXOR9eliLxYMfO4OmYK7ELWiGc+21Z9Cl8n9JmpK0luvKTQdj
tDU1P5OW6a5/eCIlerH6SR9PotcnpAs0FFvsEGNXrm4qdOZpnoxj93IHjPOFOXO/
Kj1d/2NYkQsWAP1dEmObNBKz7dyUEa8iYrVeAEbWzLZfL8SWsZLqD/STasEzjeSc
ZAQSTpXGSer8AdEkt/mYolm8nke+1VwMBLTg++Aw9z5DpvLb77MKlZTJOo4OxkDa
9JRwohQapls2oe2zcoPP+OsX38bemSICfcirpS6jQeEY8FZ5MUUrZvpgzHX2jpLI
LFp0xDI/bxfHP+M1WzhQrrPQpjm32QXkoc2+UXMN0NIJVVmqva7cb5uBQV4rqFqH
lIXgTVBARoMSZXi3CcR4wdJuSPBQcIgL5qVtw+A7H3HH3EN/w0KfUHT/qjYMdwoE
I4I32qTcZz6BpORmL8FjeNYEEMdE6/0qb3/EVfkZ0/cIxq70YDlSUAvbRDxFaCSt
/1erZ1H3/NHE0ZWvSdnDpprlzAnr63jnfncypO/9ql/axX7CKonNqzdiRAorY+90
notpnKiNFmoGsgtDknp/KgE6Q3hoxYR8bpALXqeY0MdJJ7mWMRV5jm3YeG7sYlYg
vIurtaNPVNJYq+dEgT2XXM+PxykOHtVu3xAMpf54qSGGhbVTgUKwXpgspPYmf1dh
9gpvPazkSuB1mpM+3X1X/4gbqlVJlJrdLssOisPPpCD0JMlqofXKTOJS5SzZx9K6
dP4RjOsI/9y6yZqaCG3WAgLqNCVx36QS+/lPwaxCA416WQJIpENN/oc+qWj50Qj8
slExF19FHucuWo2QLnSa3ti//fxCzs/4Dw36ygMMVxh25c7Y8LyslhQqpzMPROCA
l5ESxakDB6OIbDaaBFVuIG1XhTIhZP1Zz7ot0adQ12VlpPABTHqOQMXlPghbLJlB
3qbdtuI3gOkd11LDjkcmhPAv1YPehc17D6LrwFxQS0crRw0ar9giMEBG1DDCm2kb
mWmwVzm++HNb/lDqyz/IQVwCngZ3vSBMr+1FIKlESbGLNxlohsYiQhimEtvu3Js7
HI91EIWJwtIriRoX4Ag1O84+UfL4Qm4KNW6rP2m6qGk/fTalK6tOZilyy9oVmRnJ
b6ojU3EcO4v3rMXs4Jjqes8wzOmdjQlfXFLR94b+XaYQZBBYAsPKZ0xRLPKynW5u
ft1Lme7kpMfaUCX82N3jAPsCsBost7jHOWQuzAZyVHoAnl4+MwPcwEAE5WNmd9yr
CZMNbc+dUbkUKXrz87XaoT/Sf1OspHLQaQhIozD6H6dV+FxRtHeO4h0R7qNBT4Sj
y+KeIs05mSMxw4RO8sY9JK3U2MUaurNQHdAx9I90cdLvReJQmQ52CVuJYMx95SiJ
gxiFEmLQpmCbXbaQFSva5gpSVBVAysC76MNGcu4BwZoXHagauPpiEIUTJxaouIQ0
rZNwnhaNcaY2ww8gzy4B9RbNyOEgQlR2s4w/v49DkMxGVukXO2HzPJ8y9e5QwQVK
PEy5ODqA6ibmdpt8tqAqCRpF2uQHMT3+wbyteV0tNGqyyWi7+IBnXXTcAg6vlRNA
BHrZw189ncE7ONkmKWgQPXjbEWMlRXUtn7lCcW8XNvFrfRx4hi6qu8W9+MMkXSm/
9heQ4JYD3WNU18fQuY4LiraNgIPZ4NCnaWqnsJgij502KxttIpZJs10yVIrrJ2sN
r9Q5aYVBDbRE8w43RMEG8zbQiRmFEg188HndSewNGfpeFPyaLH/hPaN/e790m+wr
Y5/cbwEvI/ln5f//opKIT7FRr0UJIYChuuqJViens5Sh8TYB+bWxUsp0i20SEh54
OZcWPRuPinOs6vfDq5niDp8xl9u3B3hvJjiz07Mkl6aGlvxLiw672YOqbzPRaxjE
b4HNrnO3mhkMAwQWW8bfeTrB/CIe95gc+OT+6mYwKAKNCoeoMsBOgEavFRqdocya
UIlTbngPLypRvvNDCjrXJJNZQHhpGu+i0JnC8dspYXnoO9SNCD+nPTWA/nKGRjUJ
/u5gUdElwqseo9DcJlZiGlPmkxorGDnsfCu5cjwe3vnOp1dMOopcHoCqm5yk234I
y85kCv0AL9o2eCS8NAARMEc+JYZzGZFDafYNIFE9BR0gxkvxB6j2CR1boOSOpJfh
rancwdyBYBwgBSwzBNX38rEWLO7qF1CY2F1+NmL0h/5Bn0C4L7gy+TfFNeGvI7Xm
x8n9AVWZW6cgW3NjwcHhfkBPliYXiS9RS7NP1mX6aFKiEJ2qaXxqqvuL9iHpzKzb
J4G68M/RWVHAcHsWSGk7pWNOQM7kcB1J3gfSCk9qNVWp253jgKlBtAHlwcO1g9X+
B5O+hHhQyrUwvfELxUkiWlQKMIsZy5Ticcnb7fX2nl+BfRSxvurkynVWocjYDc0H
UNcfeh8blkXTmrVE7C/7NMpHEwgTEezelaabiLXVQdE4ULeQ2ARqyI4DABftgr/4
bgPVOlLRKfJ46HH1SlGp0gCByhmvsJZ/lYFJ/TRs8MJ0+ilmtST+Vxfqsb4ZB21d
NFGUZ43X2Ewdx9GbFiEYL53hpQ7uGNlov6kXCyPPfFrnxG6CONH6o9qEoKnc5fhA
VRLkvLkJrdfPQBi1/Cgx6cT8fGN6PZp/QMqwxgXV6VycausohrCebS64oNU6IfsW
gUY4cDMrcsWN2ItjDsqflVsE1pbdM3N73zGo3Z+ef4TX8ry0ufE5PZQbWLiOH1TE
+fEGfQ6sW4m4mIoPL4fO6Qq4ZnZz1+CLh8Ev2eI3ZvPxYe8VZrcVXWr0rz5J9zje
FeDIb2sSH11K7h2cs+ImDLK/nbS7eqV2vBlzYSsMyq7sSYp9ibMvCu2q0688uthV
uR8lHwMo6u6bMnz8Y6cXKUI+VMHU2t7XUfCKKa2x924SqsU8lLatSIjdemgLKvSf
ZH4HTxI1hXrztsQ6nrHB3weYOMrMPDjm8Zb9e4viOF4xB4roFvTqj4J4C35Wm7nu
HonS6Jogg9iZSShEp5t67k0wRkQumBvoIeCqMKW+6hwu4QR/CAS4SvarFrWeZg1g
85XLEVFF0TZNSnwnmeJkc1aUX+hJ5SNK2T/kIs7lhehD/lqnawIAOeqJ5EvJEXbo
nsLcPpMrrDakmBZEGKbwplI3o66Li+knPeOFp+ow3MgP1gsM4FG4sOb+opqoFm9V
RpmQRuAlIqjyhcr2U7OYXSm1lVApvQKP/dXB6u5/kob+u46do0Cr3pLQc7BUPfFP
I1AnNS5ouSTAEgp6yot1BRouAZOQa3XZQnxm1Zz4odvepW8F5AXuZbhCaiH1YhnD
UY3pagR/tj6iD7ryEYv1KRJujuQRbId8pZ72WXDfTqwf1dsR5DW6+reNKHuhptMm
wI02X9M3i69iDVYXPQRsM/HmapoBsDzoe8IFJSPj4PlptJMsg2/hagBpLZ6oMKH4
wX1cYBd6LG/g6hUA6W+ud8QwSVJDQmphq2IRuAafCvByTeocS24ZZ0nFOrAjNnkI
AMkqwzCttEWAPfBAw22MFqfNAN+EJdS3iTJ4Z53d6g30keYU7B8eZDawSg3J2hWH
yOo26eDqlLhW+St7O9T5hVuDG1DlKDYoPvJPpZkLCQQbfVY8Lu1DJrApyKPexXKy
uBlxa2w01/mfRW+UGZCGI+z2B1bM1QLPVXClTIka8zvD6Z5Pw99nEFiT8FG2eGR4
bVqQuiT9/wJW2VxoZX3zarkzxI7avjjg8+uVH0i93u/cpQeyHm2f5FN722WyktHA
aG7VcjWLMKV796H7MM12NDD5I0TSZOCYhKfwuz71RvCVHcJ8Pxe3HcWG6aYmINVA
7d03U3n8sZk6ovCvyuERZQMpt8Q9lgGOqAOwW0Yr71pa8FSw1KQjGI1vaN7fgih3
g7w0uvC1vfzykHmtNIaksmixs3Uj0ZfGk/hKv652dHOTYXsAxrwjY12p7JIA3NY/
LI3Q9tt4G10piStQ6YoLf7kFZsdSInriIwFiioTR0T8A+Wq8L7i0jpTPt2iJsQzI
3tGtA9Rjczzw1XS94qV8NMpapYhCBgfW3wbcLt5wC/fawFQuKK3D/p59gn6B7QYx
Dz193w3OlWM30X4qqWJ7DtTKCo2MvTDNWtenZVe36rSduYqfgJYCa8kA5j5XZ2UP
sXVsMHZy2nb3WDz+DAv5WyyC1XOvKEdMmOd9CymkoR65jRfhEGut8I6uj6o8TLHJ
lNzuLBHEoR+g2bCC2oJgelmtWxDdMlyWFXN91rgg0x24DL/zA7X3gb90mBGDKq9V
+U8aqtvXNk0hdNJuBA3NKMfCnQof8jwfIUPzQah33RjOZIzVBZ8W9pOXol4oSL57
tkSpoIJxqOnC7cE5s04Vfc6eEHm+E48/2m5bd+qConNh0Kd4gfgXBnAFxYmlhYLJ
d50Gw92Yxp+TuyPj23ME/mnH25cMqHh0arClKAKKYlM0/CevtvKKldvZkxictHVD
b0hcopJKp5gqYGG34ewMY+2VGagRywtWmc2GRnxjY92D4WiCir29my4FMFQoDlE+
9BzB4V/8/1/TxpgzrKZ2WIXnW3Ui7KJg5eqr6k+4djzpKEeKMU2zjOsGnN15WALe
3osURBLzr7o+zy/WKK+q6Y0p6xsECrCa4Nx0MKqZP6ks2Q2HB15qmoacAj2j4beE
bhlk4w+adsZCwVE37BBy0rCUJ/PUYc+7jRDWlWZEapDqpU2EAGk2R+wvmk1Ah+o2
CS7pWG0TTAZ+0VXceB2LzSt7E35lCg/qSiHCGesk8WxNxSBseAVwnw0iKF/RstWF
fVO92TAWG42qiOowTks8wgZYJ17bUu4lBfjATpt640xrS/UItLvXLGPRTB3h97/Z
A8cOYX0xuF2o3gOjazAfHog3t9Ui5Hm0aqg+WCdyytQPsFfxwtDkP6Fjn1Amd4Vv
k7hDP24pI9vekBr7KMJQ0K70ji0UrFwQFDCSAjRE/9r0tHRvfKLY6eQF9J7MXgVb
SBsP1Zeavmn1kBSPmF2iafwcmbOXiNGPZDLuTwPth50JF/AipbcXRAwHG2mmeLT+
ChSEvpWGblXWnWnCaqk5FK/9x80jFIc5HtZrDA2bbaxFMTYvTzllCZw1bYmhH+hD
rWLig29Ud02GLri62RLnQHYulK4Mg6Desayt1YSU1hhynEmExDjWEfV/y3bNT9Tt
TZnaREn962tHyPTYKVgMtz0c92P+QhuD7mesfZe8E4/PrnY/Sy8jSorKK7DxK3dT
eOUO71EjAniXIgAU5MxIjatorxDQYJYmmAqmIncnWC9MWVMPdGkxiq+OyYHDAi1g
Rq0KGdkAyi8Psp+w6hUNgl/0oFjZEGb/JoWKXm/cTrZxzM6eqIr3c0P36myxq55R
XhCoQo+2nxYDzMRjBgya32NCEsScT4eCrALQmnwrfeDn0MhLT3Oycrt81QEXYuli
F/93a/mAZGLHyaFoU2anjLFgtXLcm35DuYo2rWJ9nnK7q5IQMrGqsTQKKVlBC2Ou
tpdXED8RxBDIyobIemZXkpQMTSjm9YI/a3hEmbqfiCI2aKSscZJkrtyx4fmcszeN
EG8wky4yh/V9N83gZzkUfSz2DxLhvgMQaXDQ11+k28wV3FA0y+QEV2nDY7OcB6mH
nolGG84eKM6JiMa6UNNaQTrZbuTVUMzbk6zLS3iufScmAZgTsbn5H5KNZlE0/++7
XmPa7fmvYBCj5F/7ZLg5p2ZHc80/NGcMn28n8yjbZiwqN+xUntQ8p24mPDQRC2RW
PH60byLKAdypJePTXZkMhDI4boj22t9PDTLDsbjhSMOKMq8G249xOB3slR7GQKiV
pRnKU53YGc6XxTA/NlXNyfvFNXy3OP4/qFyVGpWvHZexpWRQH/VrsF8TLewAYNk5
374IKkHHviyCxmvVtMNyQmPzgh1VzAltCdBmIP55Cgy9tNfZSy3KB5sLsH0SBYnC
TEwvq3tzj9snM8UJPbgnqlVK5WzaDZEwBw1PAw3EfUjKveyTj3CZxqi/n1h0ompk
SJFYw7o5x7nKLfBUw7lfhBDmDVoY2992KtjKIBeX4hhuE3n2pcdBKAktm4ZXjGP5
fj89acOO57PCq/h8oL1tkKxVpmWKUvmCUuqmQJ7/Um+DZ+WxgO2mErQL4U8T0xbv
fPAjYUGImDWxnighPpxz9uFi4smzH4WGuZUD/cn0PuRijeki2RypV2NT1Awedcjg
VLY8kqZwEcNdR0JuW39p16Ltka/Is4pc4h2SWvloFAgpci5jR4UHvO7ApaGY9n1P
8z01r/WFTtywFbleNr7iZcdS9s55dbsvrQILRtiaBgyxZ5k8yyHMpd0usw/Hx9bh
ghOaHAsP+EjsZNT4NflclJY0kdnITIFIOyqHOvBJMaQJODUXF0aT2GXy5kSYwYbC
4laPMLg3Uvd/jBSI3mL/I9aYDfYHH4jDGKMppI5aKVdlAvG5p2Id3sUET8D/yb/R
Og3GC04zCO0A1GNbNr0h4SwXiZJjOjl2LJM8n4aGZTQ6r82y6+/C6CAEIj2htEvZ
3U3s7JdY55QSTwgt3phNa8CHp0N/afgUVQOupzpbZi4sXInVJpVYKok9JnVmYX9S
xddq6fKvAiWSxTSr1LFr/1xUu1lrYzT1sQ2lvTQemxSDXqg5SVrO+UfZllg0dCpz
ur/0YNmzV+zbLCB1oIxZSF8YBgPiUgXV5mRS7sZ4JV3xtZc9cccvvgpsOVFCAkUj
dbGdVC2eBiCSAXND6r8bs61t697pICV7PDWBEd5Q9slI3pV9ijmg1P5SrmXpDS5o
Y6wCbalpTWXi81Q1BFT8sOM66Gu98rK3XGrSvhng+5AcHk0znpVCodVD+f325b1D
uPkEFzr8SVInMHDmJrqwqFu/J/1K13Mgvcf4JrhZwwe7nzsNnJo5N4flDaKvz1/N
aFDK/RDtAv9kBDs599+tAqsiYx9oxVaNPwih8CR/GHut2fGhvO0/0C1EZRSxtcAc
eCNhXsBCpkPLJpqujtzFbrleRE62jF3FAtiYYHol3evGy9AYQgk3EAYa4FQUKDH7
6+ZES6GUUgTP/EhYzoKMBaOh+OOKZdjQiIjpwiYLrnBLA1iwgSgb0ASdTzbL1517
wPsI/qOyAjc/ZuD6BSGGXHsEJ7nR7DntBAjo23NxabChVagPNlQKkP6uEw+7vB6F
pf3S8EeLZ5gWYVGrFCr37stYHgrcla6Y36A/CST1zrzl6qpq8c4x740Q7TShQKhK
ilQSKEEp5KuO2fHRppST3mJBIrB+ohZhN6tCREyROY+ye35xd3X/UY06lmGWBAbr
cknDMM2kn3Mg2WLxNro1UemBxzP7K+Ia9GTQpmjlGAsQKDLJQDSAfgRk5nDhGsCB
62MZ+O8gZoNMUt09eeJaJSBvg4AkpSV/aZxHs1oZ4x8ogfsafR98pMHU9GqYaPFd
BpZ+yr40JQaPKATKSUHEhNUh/TtOMsS+Z4Uqv/yidzTANwLWQ8uY8f3IMJGiR6dI
EZ/IZvpqRN9myqkhTE8tUD9p0G8XwbcPWTNly1zgfJh4e9gg4q+ETS7stzoMDUBg
nD1h6hns6MsTyoF50U11AadACTg6IRAsVjnDF27Ykxb/LcuNgtt0AFuUDmK/s+RE
XiJ06edpYuZ62D7zOaqRxUtrpd80Jyowb8uttgspF1qFWzKHCorxDo0gq9e8MwiK
ng/bfL1I3hXrg0+1oM40I2BIOFewPpTmiphXRqf8l/82QmDS0vPRg+RNehKog6+y
y4enq5gpNreiiSNaJHZzNvtiVzXT30gDHqSbvGbbhMy0kREHhDpl+YJZtCXYor7K
awfpt0RH1sVXnGMxoF+xQ7N8TvZcB7Dyim7EDR8pt6YfYmB7CgpeCD2oPT6SdAtE
mcq0nwpzSCld3a6xsQ2A5bKnZ+jgmEw2RiFInDpOPWnevFznZmycMLX+bQ0UzOMP
Ab359ga8iWH7BvMc/qOwk7x/ieHO5E4c1TrDTnMn96yfLGG7ZxXUBrjD5XBzYXFM
HtQif5mJOODh5rM85mT1mlNoaJH4h0/K2abshcf6sO9kDUFRji8X8ljwyvroREoK
P4mdaIgSUruZctiMC9cJLPoENfWkgcM9ycWByKeT4vxL5Z8SBqmCurlm7jCuF6KN
jEwDL6y3d10gJqeaaCXX9/fuJEHfw+j12h9L21Lisufd/dhPyBp80x0d4diO2GNS
NqB616wjX+Lo1sNEo8COp2ASwW74SaBlyV2C7J/eFd5a1j6Ljv/a+Cdjy68o8IRC
L5JMDyeqjyjY39QrLHnG+YOrSw1SuYCzFUGJUYxg2NJj5WyCkPFwxdjj0zOPzmEp
6TxSCLO491Uby9+GnnVfKJ91PvqFdbZ5yGbNcyaaeavVgp0O8l5P32OtlHqs1EVA
pl6P2FTjmquM5T8e5nDMZfHyAnWsxDVyl0HJNw8iRaLJz5jlKCIG68LRFq64GUT7
VYibQjGYtXG8DlWMJHR2kqXj1+/aybjYCQrBneiNsGFIyeoeL0YLvQNwAxNGRaML
/t9d2/Z/FRi0ENiOgrnYa9pM6M5RHi4Ur3lLrIo28ov0n96WmWOLjbAhNdyfuKrR
BI12VSd2ciYsfN7yEHCgzyq2YasLCFPSMjgYeF/iM4rYvtR0YS9f5Z7nAomqE4VM
mpSCsOkP8kSjO4w/ulHHc9ivz/G9XjiNlLFavi5RLa0HuleN/kgZ1+4PsNgRw5sG
HSjJaW1jhT1IMZyGeTDaJ8B2ZB+v2YD+h4q0/HhcqeZXKgkZZ59hKuJ6HVCYRo6i
xfGAjegR7wHzLFxR6r6SvkIFZQU1XO5zrgwk8JPU0QHyAfKSzJbKIibRUKOQGYTs
gU5X41y4ds4KUWwQxmWOyLVvqrdpKf9RMtUu/r4g0bNpvEpvkMVwZLXRZ/5xn9MO
y6+CPZ/XMyrkBB7q3yti0NVbuGJDjAayLkBYgVHg7uh8vuEzWX+7K++ewpUbw4G1
X1MzP8U/SvqVEfO/e2j/7YKvd5Xhok1ma0Dn0AlcqvsBBojQHwq6zNt4WvYQMULR
yOZfZyU/Z9yave3JdF/OBZzaZVMXoh5Q4t2nCsBE/vcyp6Ma6zjSrvElo2DFVMsN
WVKCvllHIkSwQavg7RSO1nxYsARvHsSidGyE+rTL9ddkl5hd3eW8hiatDOxhsjjI
UKsfg5Ldx79JmzFxsvA7FGBqhcMobzhy+bfpWL6jbPTCYDvJD4rVzurHk1d5hgZh
0JkKNtEJdGv7Ca55O/PuFVKLF4GS2fxgOkc+4OzlnUWP1KTZ1RIMK4E/3T12R1Ms
O4twOn2bK/cxMijkUa9mtGX2opWpbW/M17V5FgeuWU5zY484Sl3aw6EZmdg3OkHk
ORCJr/BN4rL893BxACkHCmMV3Rk6iAvszSNjbRwrKpAPZwFhjsr40qfkp+Ia1/Cu
LsPFZBumAVkIeTiMd0ugAoS7t+tTTsO8NYS84abl611TL+6xZIQVZnUZz4XypCo0
KQgTWtuQQtV7Zcv5vlH6UDxH7xLyZ33jBJg8iyUQQz6ypVcaGrdBHoqwsDLAj4ax
DHWkYbB5GTFFPM5EG6dhxCU1PrnlOAeV6ntcBNrW8cB6jSfJkEwhuHFh5a03DGFo
M0tgh36tHXwCzl0h4xzvI4EecVKND3wJITC4RbNLSGMABGmP3VSDGUKInWc8j4oy
OyyHwc1vGAJ4HMcI3NB2Bx02MvCIjEki9XY4gPxY09mh14wbJnpLMKV9JTdR0ZAe
20O8139ezkTlJkGmp87xEtevj36vIWxNe1et25vEVNarXPPrKVMjONdoIFZYmfkR
A46Nwyc/kaJ83GmesTBGmonnUm5iRYb4SlFH3Q1YOJUCs1CVyOgt1Ztqdcw6Y58b
+J3DMUFInlDMIs/evgtwVyuzPPdGJogpHyWouYbOt6gTSlQQyUYYNmpqUGuXq1V/
H69P0tvEWqXz/55ZbTc24jaLeK6N0tmnhoz9SA/QMohmxo2Nj987Tlrbg8CmrKNB
6mKfp4FSBoljG1HUYpLhbu9uIAedO+sit215M7xyaprlROkk+r2f0bggZo6/waWm
VpfKb391ROXc14cBH9IMMrmfiUjsG7kluzdi34dDkrVByFf3ZChJ9td9iwKlYPDs
BZqpXg+OyhJmiuogF1Wzjzqr0MHAOeMfYhTFFvmlmAhvh7w3ZjG2g2qSJdQ38dy7
dFYHVz97pmsw+Jz/hcwuJkYS5/RKvx5iVpMGKNkI12stq6m022WJsrx08zMcb+lu
oVyl7KfxcWKeJPA3crn6eQcNx9yE4gSwCiZW8IU0MPd8Rv4ugs3hA+PSzlqrWdrY
2vCXAD+bh2QUwk8KpYKfmQHBPAmAVri47an9pjT6cXQ3ikzvPzZ8xEhlLoS/YV2c
WXbyd6R3OSQT4qpeclbecrOC6jD8P0An45sXYY1EFw30KbvRIzAdycKnV74E5Gg1
C3WMBWlfdf+xj6IcJ8u9aqZuCpn8FE5RTVWkTaHBeAwAEaQ4X2Glkp8TkdE70h3U
OPe1enFM5n+K8+TdGSuc33PJAl6Fc4uD5cxzn7QXlJ89tO7WHBKISlKlTqai+Gzr
TzrKo4VARVzgMi+Rxdk//ZyTqu/5IVo9mgzwmth2c2h+N0s4wiIf0Z5qEaYndQTY
EySCZg4P8f9bgqkdQrPIfh0+/fhSZG2wM/UEiwtsNRkqFdbtpI1A+wsowgWKzCMQ
aqZ3I8YUQdogLTwePy3M7QGBTemx2g+F7g2xyDWqsp2dnNhxkzaaUhi9BB7wJbbA
1uUL96ADK086BTKrJ7rqbE7NGVncDnFoDQvJSmXUd9GrudSEPKRIEcM9+Zk/spV1
RDu0Pz3xfkUS747wo2ePei4s1AFZ7hd2Ca0cDApq3kXY5+aAJsKSstNgzbZMjV0E
l1MgSTmcPZjbr7YGKME8JcSEYc/m8pQrRszHBDNeYoZYCaMVa6WUD1vHoVOfaRib
SbERRDg2QhXY1TNx3XKg/Roka32h0M5iJA2jm+F3hk6lmEI2R0JpKr78hF8sNrJc
hiTurJPhmRBUEOHpL9by6Es4CNhNlbGrqIvb/TqUEBWchvvU5I/weYZQhpRC5285
KzU4kAVznvLjFqpTo0UO3cZaggLkvPwkbSzQxopHHdPNAGABkNcPOJc6FCMMPGPa
kuJfwbEAojRMWFdAL1JNVInfHdjACM9db/Y9XStMZfuitwOqxHjaJjwMe2yTrMHI
IKSfGZlXqmc2gfrJoeQrIF5FeIVG6vYuHTP//GVDp9JoDq9yzD4hZCUtu38Zs4nq
teNEPgkJYcXEcBYiQaa0eEdi73la07Sw+DDLJZc3NrH0LvHi/ReGj3h+DdR2l78B
cNw5Z8KOF1YkuRqxfhuSF6yQflFk9oxTsYn2w4LEfluFg+nvgrsnxu43dc9rN3kI
w6Q4k2Dk4phmGC7G9TlloSjTuI9mRawxBuj3n9cPt7aII+9EacRpY5ZuZk+jLgaB
Q7vLsRBzzvdnCEpRB05KEAEP04AfxCOM3EbgPMqy/pr0g9wA3E4jYM2qCzgFCy5w
o6VV9CaMOU2Ex90ecv/IjQm6yhDzzVqe7+7QBlD1etuJrYYr39lyD+Vqxw7EsS6Q
acmR9u6jne2haqK69P6Ik9T8KNZp8fHMxrapAxLnjX6INiLmTJm3Oi72ZSwiIORX
it4L3qPmdwkT/TOdkVrGLt2C/JqY3k5Xy7u/J+rX58U5aTvKC4Seu8UY45KP/wsQ
eaEFVD5ANej/6JtvZFBpvujEBYzZCNvtphShz2QUGMRcTwwRYicAwR12s6RR0I34
Y2Dtez1nXxTwMmPKFgPqGTGj5X77QUaMZrWp1nR0n6jSrntGkj9yobpydhM98Es2
xVgZBJA8P1EoCAdoHTNh5TBbfZn/Tyj/FfnKzakJH3ZrCySuGgR1IoJGKy6XnVJS
Bz/qYmc+B8edmH019TRJ0+RqnDEg9pf3Fz62sUXUaYQJ/0EjLRCHNuSfRF7lASWg
G5ZKX5J/hY1I0TVYhXS0C0HM3Vk6nGc4dEb6Tpa9L9zdVJqrlaMInegthCFOAML8
gz2f4y45aC9pES50Z9HBBSZL6dRA9dfweylXDUWLonW4rZ+r/g4SaGJTQXfFoUy+
4atHCt2aPSZaZWDCafV0XmQ3LopA+yMBTWcm05xRGfwNynPk2/mttcaNVF7DsC86
iaIftWBhCS5UNpcVKzJ1hJpKkZEMzgRMgsZxSrfg/ObbJlOE4oXRqcKqCYRRHoMr
QIkfKLoNiF27cFPMct7i7NQt3USkTPovwgPSPu4a/svwXUsiHOm6GmcZUI8wGfIT
X578iN64LKERO8W4xMt/WWuLZbvpRWkia3HMduxavDhJjdXmFQOiXWhGEy7mz/Fn
HV6meLHCaeaR0gozP0jayaIHfnQAcf1Otv/Is8UVsKjxsxUP1hZfcxNxrzOlIilB
Pq+6bHhjvOIPqsyFhTm4jtoo0M0jjAVxJKt/VOl4RB3RJswxNd0mzsmEaSIC9YI/
oaBHmDqEg5/pNbg9H1zWm8NCay8p6lGrESIvA8MQ+o+HSjLyY9V3hPq/M/7QeQDg
qTRDrNitcg68IBPze/SfKUd/MrUqOzLqNpnOPwG3g7U5cjZFo/mMCVoil5QEb+x6
ZP1AoVLPNd4Dv4cW2J4nkyVrUUOd1zJVas13i1a1+Rq5EECwujvRwQ+oJGX6eEVU
Yn1ZHmjVwMMVnm7HzecxfK/MS9f7XFUgMSLD6ixwXmpXzJovz8RwSAjUAf+Rs6t2
2QXqehM5BZaQdKWagJQpA3Q/YxDyIj3HKtmTOwIZZk4WR3xtnHGFC5Hsw+CIehn0
ldaj+V45wWN/VjbmtYFOjDrZ/PI0eIxNvehHKSe5R6Q94AHOWYTEWwBI95lF/XPX
sW8and1eJML33we5Go7WIPA63T+pcnCyRIfg/5EjfSTr79kanh+iynwM3j82U9ww
e42zusH2poLzmXdOuYUkqxGHtCSPxl5y0HjnRTur09EqVquL0CRov5cw9Dgg639m
i6iix1RyhUcfQIh6VvG7PrDsUNBZzRbcQZi3jhblRCMKG8R8QC6FSQ+QJuWNzXJ0
r1n93aErJNdf946f/qOXY5QVNA79m6UEz6OsxXCzNp5M2YxOXVppj0YUALs4opwX
/PSZcpc1GgSGPxbezjwb0y5qlVG8FBdvIKUK/fVFg5BWVM6V+pMlfwDumGCJEx/7
+/yJmi0WcCysGHsmEiZo2pDlPT9I/LdiD8KuVrbmqQ+YvdhP1COgmARhJ+dh2iP1
jaUFyDAxYMyBxNhRoGuSNqA3IsmI41FM4vFV8JPqY1/3JNyOT9i+kKNGtO7OyQY6
+54fb+qNRPBVbkQoLjZ/Pz/uvSq3zzjJ7Dtjp4GzTxEPqbVnujlO+KKSJwlpHwOn
6u7c6sNtvemAMWmrYIqtdbK8tLUdQdugh5D174kx+e9D4ircwX3KilImaAnGh8/M
+sqUp5tmECRdx0ZEA320nytFQlQH87+KmD8y/rOeCu7U09z0GjVe8JLIDvn3SJ/l
5Xtr5CHuGvu1EHM7uGSh4tvU22wszzsmQEG+sdUVJ3Uvc9IRYzjFlXITYVhFpAWK
RgK0lYn7d+7ulFfai1TxJRxnVJ8J26qthmOrcu3EXGKZ6s/K+RZUERwVfr8saf67
WeYcjDVIc9wgoB9jTe6oeuxZM8HWc+BNb6fmy/0EFYaPXolmC9TwufvLW2vYhmnW
lKMTzbyNNC2Yj8zEHOFC1Q/hH8UCT3XbrqWq0sHs71lLNOHqdozHViX4AbMUbV2E
Wdnhqa72zATJSk1mjDB0p/1QBg/QlzhX6QTOkp1O1rFGBiL2wVprVKF0LyNarqRe
nUZy26wNdtD6BhLAi5SKXX+HqN0rsBO6WfPBbH8PPxlYNh3nhSIbewmFGoZsg8ni
je79lHyvvZvthkYzTKeo2HhTQznWAfdQBy5WSxmoqkzYrX+qlvusgehSQKG8sV4G
fjde5n46pPcL3pIv1YkschTOwJFMF0JBb2uP16owzIziqARnh+U+1WCYHghTHoXH
mqIboG7P188Ukaq13bKAZ16NIFdPyhnaFOAuQbserswcSaAAWmOtiJDgwmciZ5bC
aN7WHR1NvX/UfpZyPpJZjuRCQVm7MLiOqaWBpILsWSyOjbJ15fdgUVBkHrv0cMMa
kuVohYP0R3z/dFKSTdnP2AIUogn6SgDXJUt2J+XQUP+SljhfcP96srr+5MSfaGz3
mP1UtR2VUNljf5qOTz5ZSizo27S6tHfmB+DWxTKC2ic57TtJcW1rwTrlhaTpudRs
IylhDfeVCTaHbAI3ZHj+YdAzw+Z2eHcw6YExz1LQ2wptepeKXCYCM2VcAVw92wMr
BvsZvyWOLOo8e/UDU8geggqbtY793lnDHiohpd0SyiYqtZZj+9LmykvLkPDYv71m
XU/duCz0BLOjLS0eBNcBJNX7ZrmeWKOh6HqxuqNa/zFydMkbs1cgcFm1rEBWnY+T
6Z8WJUoBl/RonsKav7Eg8dcNHTSTLVVBBNPB4+ZwQke99b0yZyUEuz+RCc5f+4ZJ
Deqah0z7heDxLC5SWH9EoQUDr9i7OKZT2Ii0SE4cuMUMNDQgMolwfpt8WXPkCf4F
pso8mc2rylM0cIPii3CqajoHu/MDWpmlRVeb/tM00i12mvc/9b/Ab70IfVji0a+C
3NBW2qdefHCabWc4KDOPbQJtkY3JAQW/lD69oWWAs5ojK3IiEU+PVvtOHu1HUpmC
l1vAvLs62SFytu7afl0C3pL7ZIIR+Xxk93L5gLz0eB9vedeOvUVl7t/mm8PMtVB7
cpaaBX1OeybKokvwK7eRBVxLuvlxRpcH7otnyfIilKs9V4ZhQLlwLqw64HjY4Yzj
3ByAwhGPgiUUOAyXNABLBKGXXEQxDRoypMhG/3oKgMk6X2S35+asc+LtR5jyAE2k
ESpX+Xy34f9700EF6h0FlxxZ4bsWjUm6zYthqj5wyLP8DaTV6EsEQKiLWpw2uFIE
pqNZHrSD4OAr8RJArydr/MuLETkJUxD1w73/bE/OmPPPRqPc0xdwdk/pvcP7LqBu
JuOhkkY2qIjNhOyvD1UrXmPNEN6pWUPxChP6ChgnIyhcKnvnz9J0QGcznLbImKM9
xR4ihKQ5HCktc908U/WdhIekiKa1IG5+F0poKtyMMZkrXKwnYXBIXfbUCEPNw3+7
92ZOwL8CcIkuuF832rcnrJJfAL1rv/nVDJ7fnKC6eIVfXIjlxJC1kwa+SdhhcPWz
TJ95T/QvF8jbqyosqfKrzXosghQpw7iYpAgDFnaZKhz25m1x3R48jG4LoumcO4Y7
2BYwHF/4+X5nqkhccDy01LJD6ypngZreCGNYWNbbZehyUHaFytM1nbvl+8uaK+HK
BfgVPFijLsCatJ1u7LMDHomQ9KKOTEz92rNvT8ZnmZIfGSembCEaGr3+RxjH8psl
xHdoTCDGVnFVR+8ntJyTYVXl1W1GGFcV3lixoELsdGDcH8+dzi/SEnj0IyVNLSQe
beoMHa/HvrcJo2ODGbIcZuMJRirnzBNzkVQbqOGIOIovguz4eempcTzYa7dke7HJ
Bk6uEO5MflC6WXFA8Vby3TrNYocGr3RcvRviZioj2HPAAqQrLQF7enTJLqGjhWDW
EwT39ALyNXXJ4wfHBKgE5cli4weXvSbAbJzqDsHjZ1bv8JZoIw3T+z5J+efNmr1p
AVR1HWhOLs9HQReVirzCV6y4G7Pux1FOAgFXzrB+h35gOZTZjMJHXXzZGxod0arP
Ilxsi2iPjbpsGNSQ8EjsFj21Xl3kRRvmoa1efZ9rKgK2yIniP+kFX3JJ56hTk8A5
sYZ6peYEY/yEJx1cugmO+/DUUBr5spsAPen4OTzQcq2D8G5vwTbLy5/vBLVMN92Y
BxyvLHVSSx/DuWbDSvkl/o+jf822FihwccfEvqWBvz2lfLPqk4fm1LbeeQg9a4FQ
oj/FpIlWjdF8WB0EAW42sfpe8nnlCyaxt1GA0v5TjGnSD2XJdWmLJ6fB0tuX3RXO
9qK9HgG4m/VgymGWpQ0PxhABg63nMcRJjzvP4yBXyFERvY65kn5ID+NvoebJKnYE
IRJCGKpP5oCeMKCyYDo+SXg7COke4Rl8M7xoxRggE2eySqKTZwjvy++Rwh8LIDwj
h/oQiYHiLUTpHGLM/0T5iCwccQ3WdD8P5e1SSCefiqzjDLpFtKa/DISAd4N1AsBD
7R9t/zO4kRxteMwLxYm5PMM5wkwr8vm/HTUUoRYLA2RA4ZcYxVRg/ByUruCv6HtL
t63eucxOGiSBxmE+LVHjxdSqbfxZhuDfO4+XoTjCOkH99j0g83F+0ggv8tcmg5X3
+iNihJgL9Cxs7bSx31AL6hM0pq4nGtEfT3x1NVCn9iRxPq1Smhd1pGblPhHPfPMh
jsobF/t2SP4RxhUTW+6HhOPZOy6jprji/D0+QXHkQ5BaDaWfaU0EQrmkut6a1fVy
EO3fWtKkHVJyy+62MR9IxlvQUZFT+tl/LvZ8XzLujz38MQhDwvUd7Zk3lYAR5qKL
zHMRh6caGZBgkWMTOQTAZHDjQ2mXyoHu3TJb1o8SggdfNl7oISGtllwFy5vszUnc
K1zD25fbdk3RwqkUWAgJIx7eyVzrfgc0XYuhneI7umW/izjf8wRoaTIrihuKj1uy
YU4RxVXfCDDOZKHHcGYHibCoPk2QoFIc8NFM4Rg4r4iksANcGFq3mATh6yr7rwZo
B26vlt7KqI3xP61etylUeBn03i0liNZsen5wmMYq/SP4+skYMTiq4SziDHhne5Hh
3zjeJuIRbNdij1ILu7twYf1clmreqmO8MlCe/MyAAnXst29d3oO4TSv3Ni0bwyQX
qSvbljLFc8jLt2P5JoN0vdrYYfVoWcmTV8CMr93/peDA9FNJt0LykRJh0MJfg9P3
Os0KkjxLMxaGYtVeuk6qARUo4xT6/DWOvsA82flhtxN1QsKKwtDYnMbkImKZvKLY
btnm6JWYTbRNhJsUshHtK1hsvDocJc4h+q2Xko4oJU6UnjV3NCRRmboKBPGBaQfB
0JPwJtpl1xdg1BGGeeZBgF6/kJFThHrCvErJXg4b53B0X1ssZ1exlWO4Ahsn7rDa
uDeQbqNF2dzOkHbMrKIWbcqWuDlTPzWfFzI/FfdWOPbn661qqEIBBAXFX+HZRdm8
GwIA6cG2qRQCD8b2v/li2Wng1Fm2Rfk2GHXlfi+nG1gQXBm3VrSRsRmX7TubECv8
wzDH7/GpAyTO/RlQYlTP7OL7up9FyT5HoP1OejCGB89dU6NbI90Sge2JU5CcIU4j
3UR+QZVZSe3wmiikVy4/dGc+HC0GZusKa+O2dPiUNVK+iFdlsQzP2NjoXeuZX7fh
1lEmCNBAlhZUO4uq8Fhg8R/KOfdG+OG9lHzdQIoHXNFeseHwibwLj8zRYfMcLiuA
ZSeEOr9odiyPYULhEY0eT/DQsuEhz8bo1D6aLczhhHpEN5PHJLgDXvbQRFR1Qevw
ySICLFwToWT5MFyGhHkkVKGCSwg7VQGmmazoNS+0G0CvHylI5bYIcnohMgtE7mnS
NExFUNuqwnZ9t/HUAIIcDf+u4Dw99M/cxIVduMweglpXSHxiCgwKypgF+40u6nLI
edHTCzgAE0KzIPjQ7IMNwJta4gO9v6owQQWPJq5OhyAvmcOZ/FIFjUo/3aNIBSqb
vYcM3LJ6hRAKjiu6fVScH6AIhGmyvQcQgvc4mZkrTtqqlGK6yMFnyi8L7Gp5yd4m
0QDnvHQ8dwss57XGacbep8B2mYIbvPB6sdytEfyNk1FgW2BEAx/zBk3CuR1K7FiK
6nBChppyH9ZFRWjjiU//VPUxaeb0Qw5jz2THOLiHJc0lq+R230450WKJMUpIKiAq
gq5vlx8P3jDQZcdznI2iyuuic+K0v2C/KtVDWQd6kj1cVL9VHKLNKLm3fDnfz1oq
l5NtQwveqmEl4cHE6Vdm+Cdv0chXaBPKFym6fc4yJPqXMKms23wXWc7JMzyyoYPZ
0FdZSAnJ2yIz5akj4+Mxi25AZjaP2GmVffIfSkzwSh9KUW0GE0oWmvTYIJI2pjRt
2JQq+pt4gfIOPsATykZyWGCvI8cCTd4V+2DTHRMv+4HE6bz4LvMVxxXwtAOsekvq
l4wJKiK8CNd3rHBffUIOPSRd5u+vzxqlIDss9nj2v5zHEM1OYVX6Kd7yYomSxL7T
9HMUAiRcqAcWpDg82MXfNGOmL2Gm1xixCHO4LiG6WcqOBSp+IIdmLb8LaHSs3lNP
dFXpudRa+d6faloMgV8L75tqXd3svED3/5KAHFEfXtuK6GWjk+lS/Ko0D2NJJ9GT
zOgvhjdFXvB7itA1fPXe4l/MpIaltKBtyqnXHaKSoiAZ0eiE3OtP4Qbl5Bo7qj2v
UhmIJ/3HyyQ9imFAdpt8knAm1xVuoyKOWZY1PZ7Wi1ih8gGFDkcAe6ezFO1PYYJF
Raroh73QWGfy233nqxqDkADtsdS3Eps5nRANztQwTzBMT8gHriAGcIXUYDsTbEX2
lH4/Zv9oRuosEWtCnsEq9RYQNxIxfc1S+KFd4tTf+oozM25HLDTvMmypL+f1eR62
BHWaSOzGTZgd9BWm7j3mJVWqV9tomgmGEFZU/bhxYERlDTVWYcLvrNNtLXPHs9Vn
CwEHkEEoC6U1gJG0GdL0FvDj1v0Uju+2sRilMTkYtOxPz5qJPaoq/2ME3Y4wK2nB
6b8+kxstWzApyD4NrfYPSAjMTH8KXi0lKEVVW7173unQLAnWvyL3kmtFK8G0qKF0
ZwuRv9YlR4CcFrcdIthThdPiL9/Q1P7qU3g5V2+XZHONHcRFhMQ4alUsye6EU4OH
2hjxLmFyb0Vq+fjBoFr1QOmErSPhvZJQtoYTeoNdxltPvSOsRVKg/F2RFQglo1ve
XpXBgUyRRW9J62Ff60yqoaK4GTSC5ToGO9gVeiAF+CyYn0SrF0T/jLseDkCTQHgU
CJ9xX7p7GKIk5tYpVREikV6XbpNw8J/ZreKsxWcQiKnckKDHnLnrMYsPLJP0hOo3
1kCtn+wO+JCuG9NEiwQUfbkr2ufX2v2gQ8Fb2pGqYVW3fG0Ib3iueoMlkoZ7kBYL
DEz8+oKd7wIRC1b4j3+ZAxn8KKRJwJsI6MIdwAv8l1Iv/GZZRFxPqs3R213B8BIC
/B2tYjQghSzjiheC2H5ZBWtIGIUCukJ5luRIbUI9TO+RMdR4hjCQ+IyQj6jtBy9v
J2fUNPf5knNp9Q6Ki2BmkArBW6i5CLvf2qxe/cyV4a5BUG2gKPpXpAhI1SIyDIuK
RWEW02UHn/HRLo+ViNZL2oT8UArkOr25LIrFUMoBo+iDZe5O0fSXdd/iO5vlmhHs
d11bt+2NZBu/ClJM7+4L4GJtdHDQeVdGB2VdLHn41c2C7ebdr5Ehic8GPhT+UbDp
ie/eiohN7buoSWHNbovj0XpDlMmFRCqhBhx9WpYoOHh4gntSjQ+EFl2xhW3hlFgT
MdQeQ6P9Cr9Dz+XotgLrfE/n9qYTcphzl8lxqflEBmj3jVJjYNS3e9MIb4VeD+3j
418QFkzLLvOdyRXAXOgSTH93gDfJ57s3VPHSaS/LnQykKEqLMKhgvaCkByTHgyJq
swwNVhNn4RSSm65o/HsZIaTtHiG3TqsW9cxGxucqT0VUcrvcVHIYSXnFd5MmCtzk
Oyye17i4FZM13IuVRz4brhAnId1D+l6f1uIlgX4XyjBUmPr+1lhdqumwL9lAHhva
mCwuKOO4x7iijbqN5NX9NZRHH454ZE2frz0JDkWplB//fayE2KyYs+wHx3S7hGPZ
NMULS3Sc0i8Y5blx9+wAnbAS+s2V9kFbHETON+WDcgDiOGR06aWBhFr/AET/Jegf
I8kkuPBZAFe14myeWSiXe6mwqe8wimTlr0lEl1Y+9DR2TW1zWI3zxJljBm7GO6rO
yre/xIIbdBOd18knlQuB99QjyG2yygmu+5/ldZFbKJc6NFHZzikHU62CLTVhH9kO
SqRCVWmnfD3jqWqCPcsPe+iKbBTQcl0006bpJTo7ZlrQg7xZOfHl56LOvcTtcGdN
Pr0SiBDo1vzbq+xkdD8ZWuXI0oQmx8nKvcA/Evt/1CVO5/VtfC9HUgIj+Matk57C
gTKYmDj+EiW9kZxF2dqmY3nURdMGHh/Lj1kUvu5vyL7YkLyqc/HjeLTPuuAva7ZX
pgfMTMRFuKf6M7p5fFxRXqOk+4Z/MnDvRT3DE/kqicWPvqKExg9N46p3iAtXrBOZ
ywCUPksLmvAzLP4RKW+BmHwwpfy/Yx2NZ5VZVl1dLW1FJjWd9rRpgfuPzHsa2R9r
6kXoa9fRZzjWkZyr3NJOhvhlNAKv6IqXMTKKyarGwAQmmSKDBbpB6+guCbDddQiZ
WFmmDLAA33mFXJSmcl/+RoqhPT17pHovAHva3sGa+xry1MD++zGZ63cqFkZLUWJ9
vOZ4RAmNDEijPFCrzZnTISVWUQJMk25E//t18PEO1cv3BJAJgN43r2uE06/6178O
XA+YB2W6iRi3ur+DV4lOT0iWodtqGNiVotFz2FGD8ld3sEX5i1ysgs21xCGbvfGu
rDqlMjuQKralHXI1inkzavq8fAHxSs75LBvym3it1HYXpHvJm2mR8DitXl56nSbj
r21wU5qE/7IsxjlyXbmQ1k1cAX3MqYwbmecJmtlq1OW+qTxwJFtAd77WGL9ciwpe
bdsFYHf419vTjBe5fsf+XMyT1nK+tn/quRZxS+EJd5UssL3T7jjUTTsAeSirRko+
5FCSGXycRZXZwZ+PuNpeApMJ6MFKctDzF0HYT7N/wTl+Cq7HIHmckDDbbAeGboWd
HNX+M/wyqA7kPMIzLUVx+3ob8eY6Ew1zaDc0PbEyxyLUg0cKjaGBrossZD6X7g7W
jkG6DI4InZWjs+vHD1UJqxGJICPO2nNnWXCFI3yue8tML22WkVP4ORJI3fOoR6YK
kyActIgAYfDIYVfA5Bzahj2ozY4fdw1/xyMEgi71iDQ09YPte48I7fGjd6sJc0Dh
wCd2l+GhnQzt3IHJyQKCBvWTzt+83dnndSvuz2Sm7bVcfC46e2sAHzeTKF5W1scL
G7j1vjj1nr3SLi1Flvd++HksfLWNpqw/5KAsKlmOJMG4lSbyvPhLKpV4w+3Znt9O
ML9/ePmbuifpkAPdTyG65o8uslwUbMek4AP3JtvCmjsiHu6wR3cnM0UXs7rY2KF5
hIfpVflU3OWTvtM80TGkJEaY7xwz9bwq/jriLAYTKb3jm4dKGPBJ934E37Q0NdYV
EJlx9CARpbhmRQDuPiXnwj6tt2CLmhoHUcqMZon53tDcXrQRa/XNQDFMXA8N04N3
oKhZsLu6NcObdLBGjqEGTcfWCgH8a22WI/zF8nRroOu4Ie1hKN/dv3kDy9vx1sry
GiTwEXidAzWvFcUe3jvFwFKoviazQEjz1TR7lxOF9dePsDl5HwEf7YIKno909IZ7
hLS/Rl9sdfvwOpn0pv+2MJrjhK1p68lTEkKgdNPY9jC5RbE145uIV1oQchgmybRY
hbYdBOqy6OueM4/CjhxyE2Q3aRo3eaMozmWffgrizCndCh/GZ9ZnMNp8/mBYidli
2Z+GenAKIGJOOANVQ0oO7NllrvOPxFbHLgFQcb8FqtSCA97U3LSszxc3o0u02Qyo
g0Z6UyBIaV1MAkc8HdJumHhcdbztvDUQzn2KJiXVsmCBAVU/zy3Zv41tlFDRYUBq
y1gYfDejO/fTPN3y1voKbuW7RsyU8CeVOgZ+iE0MDslcSk0cZLECdgK9cW7rj8R6
1J8h4WXUVQpaSY9pmWjJiT9qNm7quhXcGTviqPH0OZNeICUiFtcxIIncCObC3iTA
Q9TqflgVklosHGq3RZegSg2pCZKgXuAhiGoOBLUgpcxBS8MuxVhT7VLAHYubiuFa
LVaOM/LCnt/wEZ3C7lhCK3Bcv0h0BaX8QRvrao+NQcqfpRD9wKJQSsqRccRnr7b4
4jT4jqgZ3b2poHOHXpK7UnkwHsYTxmji9yMlAeDYbRNyW4ah+j2g6b74FIUJesiq
RUZtJFiaKOQlH6/cBTP6HIgL6dcQeB0h+zx08DQusuR7wpOndh1lF6HB44L22/1E
n63TbK8OAtLfq7T4psBX8X8JJvaJPpcSGpVRg3oVEzzJwZCG8MZNUBV+kJ1WvZZ5
kNrQTgo5Z8fay9iDtgi9oW9EXcmI9D+vVs7KERRbw5lT7iQctmabwhX4LU0ZFzBV
wR5XlKyFVV6SZngoDHmjrUxUZmkc2Qj3TCjeQi0McwfM6k2uW4p+F9Lb772fTEk4
wR1up3iqrAbNL8noFn1jVDx1EQHNtCMgLYtwJwU33cBhWyyLZfLX7bfE/ElCXLGZ
FtBvvCTg8ZCfiRlJyseXHh3M0jXAUVnF0zObIYoWIy9JDMEaB/vTGi/ZzBxurD1d
HI/mz68WaiBUtGlnQ9pkvS8e3E8x3NbQvS/wiEE+bnUxGi8gD3yBAk9PY6G0gIBi
1AAVXGs6ubIIRr58utNPzxY2Vzk9ZeFIO4uklTnwxB2MT98zSSzTcDaL+s6HSXTT
Xr5f1Pna59ulCZzt/rlBg+hXTgUM/l0y+s2YONw6l8CN+G4Fa7vVe4Drj2PDcUJc
rB/XJg9Dzl+LZcS2L+unzPFI2g3q9ZEQI1Nt22upfUJ24tMoeSgBzCPMVze652cT
8Pj9SA5MWaaPSLmh4MUhZ8lVO0CVcY9HVYrfc3vEvFDUT4M4RrfRSPDL6mFuIYPW
y05LR9ur7pN4yY+0ozwrB00DmLlUmLaG9h13uvuGux0+CiwdqLOLxjKII93b408V
EWY4JPJ/LpXBpOAP49Rzrvv/kaAaaZQOmiAwVyYgbr0NtfKCOwKYiVnIK9W/2e+s
8X+3dmmmh+os7mj54rZBA5eKNtyJCVgMJEg1AM0QkoixtDLkTovLBMrz98kSDGh3
Llc1d+RyhfVTAER5Bw0yEC34mDjFr4QWZB3SLxkAL4eLjGkohffHQj9akVDUFmcB
97xt0FRQttmc0bhwgvqEhEXz7QoHHHuVzq4M7LiWwHKWbLyiOWDObL18XwXdyFFL
SZ2dLL5NwXSHCGkQriNHVTA+2BYViNt/Y/+qB2XTlgpko+3siLPIb9e7GoItZEUy
ue5maQXGaIcg+7NINFkSy8rGdFb8Deutk7bPVCMBZlUvroRC7oEYO9EkQqAyhJwX
25LFqFm63qM+dVp25tbdmxx1ZMEmYABujPHqA4LcAbmt68s6TwkP1Gx36hk3gQLD
RJi3ObQgvlww7wCMTX0486nf91RnyuHwCMYnqK7NsdpOehaC6eTLPjNURSDxgHp/
6sUztzPdTEEdHgk0lqthoeNqUSnu5pqC+rInv3cS/mDDbJh1RDAMMTvc8nJs7uZK
Ot3ItgAZyAVZjp7K+xxE9f9M8p8bmaqIrQFyNsT47x+yyjkVbkr+iCDAG8/bcW0S
/B8gRPDKGB4sdiVwVlD6CA05nLAOWUei+IhtDEw3WHIqQ8nPkI0yPyxQHJ4F91t0
CfV6KFNwsabe+D/i8VZGepGKrZc3I0KIF3vmrJoXBYmCw4s9huCFlxMH0ngcjW/U
WF5luRBlrTYQLbrmjU8t2LUJ3rhTaTanXpxrcDwZxFGoQQMiaairVw82ha7XwHh2
CqYJpZPwhk97AFRiQsK0ITi7NvKjXgklqbo5ntMith+sNvecVj4iTtK7v9VEWtG8
/E9d1JnzzqEJDEKvAeJoLihK/pXU5JgD2CaN5iX/h3rUrg1GPnLmzBuTyxLAAkUe
a4Sien5pVJSR3oK8YBAl5e0+8N0ZWD87mIwJyNT43lstQ+iZHRrj61rhCWrOzz2Y
kfACXw/XHB4lzVbnS/brnM+UQawRfOL6w1QTe6kWWck5t3xfc/uaenjqRMfIhRdg
5BqeWcwpLWSe4SfKLqgKMXJaapMHAkQxXLGBUZiQUiq0DpTiGwh3kA1S8PXg6YMC
JD5oZvhOrqSyFftRVky8t7/XRnrgigQCi8gqpKMsVQO/6/F5PWH86JrLqPxFTy/S
u3rmcGDV1WzqewaNrkezsXux8MRc3FTmlXi4hBppDWxLflKiVbPrA3tvMdWFvMoh
S+JX0UUmA1GGM+7LmmsGPw4SZQG23Vdo+EUtgXQMfICDmGTQm6Ah4J6oHvvMyeTO
IcR58BvQEVFpqF6gITqitX5T9rTa0bpSjRDnDwsjIn+PdW+RiQ2gmOMIUr20gVXm
OJT1prO6QfugnBivbXAWH8hpWou/qjU3Fn5QNhaynTAYYzYrwmBAZr17lYePRd0y
fZmQNxxztIA//gLHc45F5oamWFdsFhJMx7XA3KnPfu35zfrkZcXZqsMf951tHjf7
BlpwWyQZvRyAqhWEe6L2biaKqxYUr0p1udmfdmjNmHecRzhPVwAzzFVpDzkV3/TG
2ZhoLpJ1U9LpWlAss1tbpWhfgoy8oVIYOMJrer6UpkomL9vYwahVYXPU0iS9z4z4
Qdhn7twJqrBz4TUdSrnGx2CoffT/okxiscXlWEIZe4hur2uHYfuHryWxEdF+Jape
Tz8uI8hMLOIog47z1X+2aFhtfot2l5ZlVl8glVyzae8VUqqXKiRh6PdlHKdZ0TXA
6SHjQV0TvRtc4X+1ICtHfDJ+fb6s9nY88GMZXrd0yjHn68POOvx/aI8dGti8PxuU
/McvcDWtKHTqkQ4psoIdN3Zvo9HFPO/sYTlPiyJA5AJuLijlicovfTeBir6bZLND
Y0AuqklgX8USnTRk7uCBQg8Y+J1NcO7w/npPemd7q30kTQoaMvs7MxCJqSZ6FvH/
1ntmOPHjGJc3OBUq57wB+c6o1cCOq+BBzKnBT+V1vqSJu02ZsebTlffqRwPJAabx
Bk/y7xhmGX7BpnEPiEIZwzgOhhXbxnElGoOaJYlmhEDfZ1INFl1hCkBbiMzWr6LY
ek2Q5wb4JSJgmfP/rzoAfiI9MuUJ/f9If/iAefKesFiwHdJwj/VQ94pb3XOAbucZ
qun8PFQRcauHb1yRMWMX+z2ZSun4Cdehc7DEZ50ZFF1qxRhq3WV+WkC63qtfg9sN
vznPD85vpF4u4TwdT2LQOotvkYPCfWjA1mwnXL9iCoxxisDG5/aZeSL10B24TMZ+
oBwMaGZFOvMktFcOqbTI/hH5HQ7sz3/kYtVNGiZL1kgkFh4ycMrpSRqadXom+ZcB
RXVR3qobTtEUOiuryPKo7C+g1fp0MSSL7PEYYOKOEPeWUST77rrDuKATJKeNUFpX
cvjEcubCcYnvvGxy5InJ7fI9MS0dDXAb7iS03wgK4iERTgLqu1YWd+94l2O8Paym
ynX5J3CivB3lqQmCGxQycfnSh+57GMYRNIciPENpH6K9SzNhfOMvTPz6/YgFROHL
hNAmeTQuktBOYNDj1MLFaDqS5b46qhMTCmvhfNPCAg7j0b57oDwG/vo/c9WiNzAE
yYmuErNrk2Y/mWeaH1BBhOm5ukGCFVGZ/7c2H31SQp1wD5gqy1WNnNQ1jw9zchxr
2dgkCY8W8ZbC2U7YX9yFbh+WTIhciFTgVxOaI0RV+fZ2w53r2p7AwDNGOMdJpuoK
KjdcS7B+V/+4qGqiLVZjjU1190GtQDTCxgGPrD8CcaFJbKQetlWLyC83MUmxVvfD
iHCBfMPGet69taKAhfTCDBpRtFqnoYqheTzyFITwmYt2AXhlpMrRY6AtoFq0KF4T
E1WFQEXRG4w2/gNHLkVijgHWkyvct2KM/rY92cXWu6SOQJHCafwg0lxUEyz3rozj
GPAgrOBCRBgsAWSfqS7DOUSnq2+DL3y8B6es9xk1op9RQ3Ly+EDf+oZcwkR1uH8K
WC0FOIVUoVMjWjtuQxJUQITPtNmNcnAPaSwjTD9rypAGwnn2mLLeJWsMlZUuwwST
zwXhhQ5Mt/kibVwUtcNsy75OAt3uDQhF2C0SlijGKyTU/9ha0niYcBwduhTN02rJ
3LntNzubeKyb1fmf3tObA4tLl/gTEhD4s+gHe1oW7Sa6HDwQRA6PyCPyuLnLVPSl
0g5b8CFeURpXifmdJ5R1lxW3qygxlplEs2AtQeqXmvX0ySsGNLks3gXE1rpW0d95
0aVARTHI5D/64Uju01gftvwqTX5Qi2F4jtgFkKV1XdOXifLBqtQDUCVIP9+nWnzV
nY+RiOz9QvEQ3N15oN9XAgy9P5KE9gVJtg9AdsaquzAekUjDNPU4GnQvdvvFXn10
TKEHXVwKcpPDHfaPOjCLoD0pUYtHRNWCzWXJcEsNraWaXxrJVAmSyQmK7qqVOemX
ikonKf8dJj7JoO3Tpe6/VSkwtzOLQ/YCJBV9AwrzZyy5+IUNyKDxWM6tQ0MI5u3B
2mXYuXPfpuHTIZZqE+7tJ4WF1bgE4zeqL9cOn1WDRAAR0Ww+/jgl/TqpqBDIITWk
0Dwc0h1Pdd37HW7pkhQ1yRgf+9MCl0RPTuve5HWqShEG+QPn912J8pHBcPsttq9q
Wk9pPGbkDS2nIbVGWU9G5nu7DH0N4pSS2m4NZeMldNLYmSv1tqnOFeKz2oTklMbe
9VqhSNtzfWTC716GscG7DpbWEZ9ARcdwgwWxv1zrAa4PwfV15/4vl+2SWhLM+mgJ
UVb3/sWG4tXpXtUsgaPUc8t2ktPzJIa0r7Y8HWD17GfWprvl1HJy3VBDaSn49t8R
U6/9Q5hHFw+4O9iPghxWi8EiJlY13SpyDjphrDPKG6MV67xhEmK1V5gNxmtfrRU+
yhDzq11DnjOiczv2YcG8Q/SQn/kB6JAZToHBvmAy7z2131iLtThIeaEvbfQ6wgHg
UBwhaPkgVpBzKSqJvBLisleicXhncoMligaRYufz6WwFldpmKPVDs+AMqtGZv8wm
dFRT7MR4F2xMuBS/O8iGYDeFL46gpRYRDIBzzuwoI1ERoAdsHPJFBsPQA3Y0bOpJ
bVHiSX3CRR2qdv+o8FZZ7ZvD3N3tzxo5viWfBF/HLCGO8hW6Q2ktHLETvlkWcmnv
38GsaDNDYSnGiwDh9QDrjZVlnEgau3pvMing6sBqQdkpLpy7TmZAtWtMzTvZ3zOj
04Yeyft6FdQuBIBGFjilqpFMMSVVbyTIyDqz0aTzaS0KUYxIBt4G5yMZUd3jsQGl
FXo5P73P7S2M2DM2FV2SR7z0PPZXDyrmdiMRqFJk+en3eZhjNKX/8IKYddSfXIpe
hBLY3jC5jO8IZvb/oHQXDhR7qk4Fqp8nHbDTBjiBlAKHUK7O5B/vBRcETlfVqIpT
GCCvfejqqLNGN2HhqP+o3Snm3QOrx1zBpjAlI14NpWteUsmenVBAPkcNjUBK4gAL
rdVB5VfZHT7IBKxa5rvB+J2raGhKHJV4RBceUfu+KVwu33Aj7nVY0JWvqZTphb2B
mo5GS/50IaKLCLxRdbFBkoMx0MVo1mng6OyE9g9IFVw7ryhEPxiBrFyYW2qwDsNF
oFg6UaLpi4Qn0LI2yXC5IIdgtmT5s9pp8HmOxASC3Dt6Bsbn9eVzOc+wp6peoKxL
esnfR9c0xFS2hQWOHMccR7BBF7KMaJwgrQIAMIj5YFOyvcXREbTU5USLnqGkPian
VN3DI552EZFIE/eTRetO84JG2RdbWP22wMZB2Rzn1CXLtheczEP1EHr8J1ZHMDoN
trFQ0a5GMn+wqd37tWcSnfF1gJ97YabAI4EvVfBqhKuXN0dJIVAhRzOt1vGy3nex
J6Pq0qbMrvR4W3kfnzFTcxmFktmmHwGPNyEa2iw3tAeOSSiCsAiGlyU1J/Joh4IM
xL99nC3KEAzmggCYPEa5EsFQf+kdUBQqPb1UXyJg18bPlHnx13HwuoPPq3EIiar/
8o2PKH5F0rIhz81t7EphV/yCjDXi2CelRRWafnHppzjfjk5+50wce95eR1VG8SJi
wjnpGEFG9MsKGk4CFVS4dYDtyjsyRZi2SFZHWMoR8xFI2bAQ5+r7OcIUi1sL9Lkg
7pm8SrRHpwPRMqJvzFRuQ7W6EiuS1ewRNYwNRBWJhVYdhyYqbAe3W+61sRaUumkM
x5tix2w5E+BDSAWgolUw8Bmv508cmI9exGPvI7Kac9zt6CQ2Dp2nFmVzckQvBJNd
ifys+jt6MMHSEbbrRH18XOT1Ilx2oZgvomPJhRrEYNQiVLb6no6I33UJ+xVJJQed
cpW+HKFMxMuHXyaHW35rSY3tU4rYYKlOwxB6YrzruROgTcNFm1833wCT/qsto7ub
aUwpSHCSK8nFqTRoDxk2EcsLy4kdcjdD6mijQ/gub3VqfRFERAN9R+BCk90HOuQv
tesiGDI1eNrqplhcMJPd+0P2Wc+3VCOPezpli4NHfv72JVCcuLGqF8xg4bRi0yTH
iFR2SIAa5ppdqV40pF5d0NynCjtk2EfUhhU6vS5M4OFofs2K1aeZ0JQM25TT8rX8
ZsFAyPDKjJf1ZO2dxABkgQEYmnKe02ND9xGFfzZIxB41SzC7Gx3JsKrA95nCCNtj
pmSHlYJ40hHXVz0vqqbu0w2QXPJgynTETDNlyBhLDc1KTHeJUI8KzQqr45aFCiHq
lgAgyaSqYkaKchkgu+mvAQ2PM3sKFjv6gZcoywboaHuBhzVQqfaopaUhqyNBHioI
sc+4JyG4d3MlVzjH5amrOAd9EWyydm1gKix4+hEOBuiqh80b6IAxN5tGz3NyR9vl
odNN5AJrAPW7qNnkuCL8lYZ1l6uzqxEEKNaKvhfkWcEnLpejoBNiP6T2NvGTP7GX
nxEodv6zNoyOdSqXESR26SjmEy/iaHnUvXarEiXWWZsNqqOaJnX9XFCLqPl29myM
y0irZ1lIll9R0VzLlh3tOceb6UsaCwQ4D3Xh3uBO0txhFH4KKHa2CZ9CgA7vGkZa
9qx8Kg3MXcItAGSl/U0nj/iTNXlwzV8tJD9VqmuTFQMCBTfbfzLEV7WTr55c7mN3
KYipG1vnAgCJTXXuh6DigeiWQhckcGkPBbjVxSXgzWE4oG0R6jGHxso599x1FvtD
vsqEon4bVXsnzfcJTNn4IX42a2QomQAGW1yu6vxMAKKMR7FEupxdgiy7yLOgeIyc
l6sfxnswKU+zUCDpnvSEoG8FpSWpIdLUYA2ckFXIRN1Btg1gyDxH+jIOJWFETmuv
XfPWDdo8I3MBUk2zp00VlbJH4IwdVJ/J7kzv3AOWvlkqBcfEVpsaCXcO5sVeF1Qw
HVHHAtcDPsama0LxnuuzXUHhI6VDUAdiVGpW+EIWTkoaNfW/qZms71AIk8voQ4Nk
yh3z2XFUl0DsHy68IR/Mkh44/7Ww8o05L6A1SQSEBd5RYnqE9jrRvLhJZiOc1+1/
Mg0n8JbKYWIwxMaoc0vfS8405gGFANTrJ0qI2s2OE5mZYqbzp388he864iYhvtPt
2k2WJXgZVShFsSLtZICs2msNBC8LoR4QFkdntObF8yKX64HEURl75A9e1bhqekoj
6NTvRyoiYUkeW9yXoBJV7qdppNwci/FpdCnFlH2wpmS4zJgS+W2fspC/GUWivIlU
8UwSL3sP55sZSvvsk3sLcZuR+ShReVcrAS7vBbSzZK29eQFyln4Hk26R/vY4cym5
qpwsD5DxhHfrVRpst65C6lGKYv8sL0eCK2829p5NxzI+fKnraAyn6kL861odqFcq
Cp942Y2rGR7xLNU58YI0BwnsjW4PXra6FY8BmJ4huHs1OC26qzAw3s62llPr13qn
yn4FWem9YrIft5ZUdTFaKPx0k6WVGcTfZzS51LMIjKPsT5ib+0R/cEoVqfpptr8q
HtjkiE92+g36U1q71vJgHmSzKLpRWV+WXBzYnL2f+7q1Akf54qaa2cyRwIgGVnws
QuqtXalYhVZGtSLMs7D7C2UWdpVioijStRfiQKole9/jHUyRTh+oUvXk5LkMha81
J4qxhqw8nq/s7kjJZXUxTgWxm4cQMHk2QKizL5w7ALyt24G2IgJsGDslIZ+ueEun
8qcga3ZZVJmLSoNoyJElD4sRGKeI14bHM4BxLbbQYvFXRLmhCy2s8qkLWoWzTJQz
ukLe48TWRV+8Ko0Sqd+ckpPN6H+ZD3exflmAWBTRCbciXRFEwDAPlmjj/x6G1chO
dISTQg/x7ODHlI8z06vazV++sGMDYK7vKAS0jqANbk73Zs5ewWcOEO07mmy8I0XU
41hS9XtKdfVZLTJT/Ez1pltkCeq1qOgfUHvgidnB2xVNNnFK2gGD5Kb9P4NsvJMR
QAAbkWclfpYZrBIhlikA4fDrPJJvcahzHkBePN/hPS2hx02ROlnIHxDo10ezS0xh
qW20hY/MEL/8QFgnXF9fyVuMudGdLe/z6CDVCHqqiGFXdmUhVZUL0urLrc5gU72f
yLT4p50dne9lEnGfqFe18wQR87Z++2uHQfpWI47wCbDxpvfcOlBpC9QnbyWZ2lqe
R4wUfBmjNum4SHkJ8pnCtojEih6s9uE0704AELdgVXEK1MD6wj33M5YiODhX8PYw
eadKEhQu08jyHzkluFP4ljqeWwkkv70piiJeqg/cKJuwy3UQX1G6jL/MX1PbUskD
6sPqtY+Tc8pqnGfmh3T5qXCl5ZQV33vrcqkOm8EH/Y4nHaJzKKY7JMgsxzPYCc+w
SYce8rTzN+2aOweln61vvFU77c/UkbfpTDDoo0/edPly4gqr0PG6KYqy+EhcaqlK
R0E7Xj1EUtNaFyOtsFc2h69JR0UE1bOM6bYSWuXoII8pYfQQjYTJiU8EzaHLIqh/
rSLeQW3lODAs7IN33hHh4DZuchRq/uHv/Mv6eoqQ8Uc/qaOuBCYaVR0/auqfIY4c
gbIuFWA+z1BK6ZqR2lkhlcm5FmeRdkAyFRJofC6vZ64p5xEH6RSoyssEPv/a17gr
cgHeEEyc5N3Ry0uWRxmYf54tqkaVHYOWv/VWcNf0S09gez+F1TwBGarGQJcrVvb3
ZCV/VZVD8kymkfw+BihP56d9q5PHBb+7yJfoEEtyBG9Lt+AiQSkE3+Yy+tQ0RmLr
tEXqLyjNfbD8MSQa6fnZgcpkSKonkS1l18X45jG8YeyXIiTqFx+Bg/wuQnR3DvdI
IvaQVSuZS/LH/Y1YIktYR5eVBVnYKY1x0fO+4MZl5m9h6JSgCUPbV4+Aad4WqwVO
oC0W9sDN/Lm6+cMu6htsi34GSUY0h2MzqaJBPnK7Hj51qtwwoK4FgV1aXOVig8p6
rjwtoHV8HaXoADly0o9h2Dd7dOKHhobi6mdwgutYXQrslFXR1TOCpP0ZKdPuT84l
BikHmBIJf11b9WbreQbnMaDy/7Gj64LvSF57YKE3kyhyMkhcuILpdWAI1A7YinsZ
CCeTT7MzVnoEkDXUKwkTQeyd95Qi/S9Z2sqzde6KgVTrwZnmDFvizoDlBjAF7Yfv
fWilWC34xxQlRHMd2Wu0CVkj3ryzbemU4j5W2WHDhtxyrLA1yuFo12/Y/ECy9N3+
PWzywqnf8uVubefrJMzNSy48pM6mp09noWbURNshchjqhDAed3+7P/eyGWpLl63i
ho8pZowPvo1T7Ei0X6DAvSYyvHacKSQMG5lpxS9aqI05qCqZrQeKB+21ei6c6EhB
nU6klV3oEf+kkPcqiv7oFxeWbAF0kXQMUsDtR8qL9LRwYSKTRo91esEwvT4FAnNb
002MnBu1peW0Kq5GoTeqt6AMwhLJ5irLgtn5lMp3RPEcC2mxQoKkm1hBRPILkLoR
94DAk9LySX3ZCoQC5dIZdvFGuC01D5q+OpwZRUtXh/VHDzHuRgv6X3Lw5fpKqPG2
GNXX23JQ4cd9hz7UnTmzW16fkVjXyY5e95XZ8mLUDakLsiUJvWURVpyB9IX9FT5I
UDgbaGk0H50FxG5ic+BYxG593RnP+/kdm/hy9aKFtAdzix2LQf1NWgecKn+H2d9D
ZW6hCGN/fn2DG8xHwIx3oV14T6XwfEHOKjStz7BFdbfHmLDedTmF2ncFCWfpMnQ1
+S9jX+2iGL2q/CriIXV/ZzWxV3aad+FT9qiwwOkNpUHJiRwn35c8d07R6DYT+m/o
L4haXAZ2Twpap543BSQq0n8ajEiCzwpoyGpiB5cOJbk2sNNviPC79UbavpSKA9qt
ekwV6vHygJMNuAEnTmpwwbIFNFy4iJOVRH8qnhOTpU5RNhlIvbMgim1S7e5oDcL7
yqJrWeRsjJI/ww17UaiyGLQSuytDk1vpnV1/1ePXPJOZG/Z9VyuISzjFKtlCI8B3
RK2fXDXm06pkZD8xQ0Iw6XemLZWtkokt0ghEFeLbOIOtv+Ra+IwVKthuRiigN7Xv
bUhwQ0WT2Tuz/XLgloVryyLAUDBXIMKxKEVHZYJLGSkyOMirqCtQZ5BpdrFpuvUt
gIR3yr5hfWVULiTHOmzUQ7DbqU3+np2PsOUuqU4ZWSUK+Lfgelc6fF4iq3GeFm7T
8MzOb3SLzRm+kqdMXaGrQPeCQKWYayA6A55b79tF4TgNXZz5ocf3Asu4dHCJlavR
pSsapoyM1Nkum9I2sr/9XWdjdVY9QBEoHPnwDZpbViCiA4medK07rpbv4e+6v0Va
PDZ7GCHOvdQxCtydk+pGMaufGVKJ06YiSG8h64bav+xnJQbmkavqJWcGlg0soU+U
WAD+pYJnjDZ/29wOikMbP+Cigl3vnopjb588qhV6ldP6ivOERPULPbVCXtrvwprY
QU84bxqNDbnUEWebqCnodQalsVIULaaSyK/DdANPD+HiagdR7miGDjSrglPG1Dsm
YeQ3NVDB58l0fBy57yS5oLzOeCtXU9qSl90w3SnKH0fS4jx5Z0tL2P6iZKwljgV3
WJmeJwlv60uZamGVaCoNRNanjrOzp6DXVcdHpI0EWbUXLPHqbBZVfswnp2MCujc6
vKtrZVFggctpePCe/2a2M+Ka3meVsbF3qVgcBFzFMApMDTZZXg8QE1jOOqxxcJTr
u/jSuXkOR8uALoTbh8cXpz6sRYInoPwyHLaeah5Nfm+jGhVmChVSbcpKQ4kdlb2M
NymrW47Lfy0IspSQMktqhXqCOa/06YlglB8y+1iWBE0nSkurVdVrpx3CKEdXF84r
bl4tamdvPCWKahWi7jsZAX0UaPFLLJIzKcAhlH55TLmqhh/Am5xaoeVavqupewUR
wQQ90dPMDtWekhgSH+OM2a1XdYSA0HwifZdmGNAWgUF0PVRKsWfRqIhJxZy2kA5c
1DrIeQVDSvHDg5nG7Xk2wkaZLBwRmI+/rhIcDKMxDIKbImjbPs2I0tuFOnG9+rls
0FxzqK6vWmyOiuTTnaCxlKkyTpJs9WWTpa87NCZL4TOrl4Zdq4rY0lwZAxrQRBOL
cpeMnTmyo7hHbpcEw0t85+G2elmWiiUYLGZPJq3pabuR+h2Ys1O5bdTR1jm/zLtd
Kak39oho3+XPMfH3VfaGwYAyRqgB0T5Fez7vrlg8+7+1nvapqY+gezsynUv3sTvQ
KGc5TtIwc8IP6ABCSz363t8HLCKuAF55nKTojpY+DmnS8TStRdc0q5QLswOKCtsr
8fNKaFrfNNB9QxLsa4eUH106CNUHEcFqoC9HJ6137YB2H4JsUFJ2jiIZpGDkmZL0
LcA2L+sKTVZuCj4AZUAQr1866NTxh0dfOtAPBJIJW2zLPRrpAvUAc+a9Tjq29/MG
Yhu494/2hUUBY5HQzMkHeR/CPvODXzwpUaB4Owo09XjkASQy12mi5g40c/Bv4pqF
M41O1FL2+P6P7ZErYbfe4fxlEe6fi4CyuqYpLxdtXXPkvwV9iFXwPveAT3elIxf1
GlYgW0carYO/K2r431WHPeMt/lYYJ/T6SHZUXOOCuglWfpwxq/HphLKhgq4tfJX4
f5a52lHDGtAYWptJGG7Oa8mVNu3bdJyGy3uJe8ytuLFxntlmJ32lQFf8ibyR5EXh
IZIaNJUu4PYt+B0sA3WDt80/Km3aADAfRqjbrJgdffzD2kbo4vybjpVJVf5uEkii
aRspNbjsjVIqYBoIC7RGAE392c2bi4Q1HeFA9qFjGHRQaAMYMIn4XoUg3jAjAE2u
eXccpl/TXmdvjr7hUMVytaoKJI5qmT08Xo4MHasqOP7VVbXOgDZXgSol0qvV0FXn
nwrn2F1XFWu+0652HPIjtFd2e6TjVIL6M71LWCtQmb/wD5Mpo8IMq1596Uwz8Ouo
fIIFneu19neqhZE9bnBEDTmqSnp2zKKcyth1AF1FDTKQ2N8CWPjDApCuJESWOfqE
ILK2PKUL4/fHaUDWKPdqP0jtt/2NfSqgsvIkpAeCXccOFDIRnVAsDlI360qQz54d
jcbD/d9B/1I9IY9Sg3HYumc02O91p7fA8ABy5QeaHSp+nyIhOPZQNRkbF6EP8rJ0
NnjOgmCwv6FqUpzw1RfG/a4paW23Z20m822fkoU3+7Y68Nt4VxEEGXUl11wWPQZR
8tbRzG8opWg5bD4wR/t2aoGgrTsePxRcN+NdtBTZpbIG6+IUrPToxpDEJNFWMbh8
aUpJgBYHjEg6e/sVhAl50Rc/RmwzkcVJko5zaw8s3dtQLQTqTlmblcWnzbrEDtJ9
GVY+jHT+VE952tuycbyNggAxaUe5TlU14HosVoZ5DSjiX5h1FBP2SOQ5N7r6uThJ
oeZ41u636mD80lXxHsqBpJAOviUiIUgOYni11/7RrXptEAuxn4AJEM8312dhAVoX
6Q9hBD3/aVdiVTV87oZkrWXAzRqraMqy+Fbici9mJe3AuXwdO2r2ZjE204BjAO6O
IjGwgi7zw8Yvju+G4k4ExTI5qAuFkDxN5W0TB/0rH08qnUWJwRghDXGc4m7r2ui8
BS3mejQvr8RcedMSEoh6l//dU69tHsKdHlw5AdRPHHikG3i+5Kjpn2DXSkWedcVQ
uRV/n3TYcz71P+R3th2fLQekZXgiA+Zwg91UWEUQCj+RQo4vmrDtps9XhYhiUnrZ
ipJT/16s3HoAR8bSMI2l9P37aXzUGvce0V6DpoHjdzvV2xUWcx3IZ2wmQiNjiDua
AlprlF/hhHaC1DI8LuHibNMQZ0rGzAdGqEbkDKBoBQVz+6yBtAUp5uajJAAYgW28
HcdraowvmklTJ2zaOXpnoHYzsglMaEokIorI+bKQ12YVWSF+8r8HSlzJGNbqoe8G
PKkMccg/XLrHXcsfBMHoz6yr44VFtomOGneMkOeYzIuGhLQA1TiMsItD32OkIAUQ
7pszLL+Lyz2urd17X21D0dCEVk0443WFGnWTy69jpwfftIlgDO2vKUAaBF0TbGmV
HBN6V8t4Lkh06Y+Rqr8qwF0n3lA7SKklv4NKyZW3/0AKpeNOzGorhtN0yxj9scbH
9RVHDlE+7WjZ/fcCfXYIyzqsD7FOuC8LHHrrxecXXywXohavU2eS2sxLdYvD+0Sr
nxCdJaF4foNO2OiQlFdnImkcVVAWazZVQ5FDZAxDk/zNsPH/Vz7WmfGcsRRjThst
lVJJOP8vu1d0Hb9K88SeVppAXeZnaGSCB5xFdkd/FsXieE14clxPvAH8Ycsq5P1+
H317oTpt3NIp20CVEQmBHSrQyuysp+9VyuAclPZfwFOu/a7fcJH1yscNbclceYDn
Dvj2W9Vd9YbgPiSS7fjqn0F4p9cvs68PbVbgOMQDH0OvVOXky5PZT2ZonhHISLr4
dQXQPgtzFfkFMbanMDlNwSoiqQHd7tvpxrZrGLk6QFzWglf3zE0D3CRm6F6oZNkN
Z8cOGuAzP8uWYP8G/xLSpDe/OYzmgCIXVqq2/U29ceM5tQA6wddX2aPZ43gh6V/+
WsucPSBYMSxsY5B3a+Erd40n/RQKW8VlsyeQxl/o58IhIUT8wMisYcLSpXsIpMCZ
afJv3KfY8VGGRv693ub9pOGknicSgoS0hUwVXPXcuRvAfzVVUYHqCQU6pkDsXRW6
TBSY5fxJhqST8KMNEFqU9hPV1kXHmlcH5AJeD+EdSkA7GWWVm1DuoHQbQx5tPQe4
FM2FL076P6uvxAwK7CzvoXMsPp9V7Nn4pMz6J8p4TSd1K1kdz+XQlU6pQphZACC9
HvHp20zQvSTgLx+vNzpxIGSZzS3mSz5107+ktK4L7mhcBK1Q0+Gr3KmanPjvltw0
iDdByTEEbGLj7prv2NOXFWlSI9HQB12Y06IoZTVRT4IBUVpO+TiGCt0qfZvlld8t
sHwfgq7DsVq1M7oQUHAnybHNSsU1tae/QLE4Alt3qXauozegfMm7rFkwmYx1zptL
IbleZQa/f53Cm6ZEEV7FTcSndMUV4xw2YvayGAxrhCpl8bsHQvszyQk9Qxnxz7SZ
Bcpnh4mbgxWs51tFwLxIvr7/MWXTBM9x9krla8MVN6w3BJP56z+oWX0uF03TOW/c
R+Ns3r30bGp00eBYHxbljrLvB8j5QcfUK0isOUVI8UFbFGicBcqIFeYsDTESc2YD
VY5ijAoZIyJf80mnqCXzH72T/VKFTGGwUxCv/HX7OzvVoaGh94kRiNnD0q8xBYiC
J8UixDNF2/6seSvIF8a3R1ojcCoFQNcaw236uqO55p/Y08zCBwl6Tp1JktrW5sPa
Y7Y8aWuXSbY6T+WYE4hRtdO+3f4767s8NMKg9VVInsMMwHXIDniSbwcZA/4sLXNU
uncvH2K4TTpqtTFqRNzZPIvalVzryvJ30D0W4XfDeYjN8jEGbCElwCmsqhy8Msx4
4pWEfGT0tmXuoGehnmfABCQhtIEH33Xx9wIvjEtQKuexfSL+LoGa6zrbVwTmCA8u
/4v9ZiYfriJ9dFWI63TSbxfVxGexh1mj/wrvvAROw87AQWh5y1/e+oann2QCpbwT
B7VO5LeDFoQRaaGClfXaLjTprE9qIe5eLPFlk6BngJeVB6qB8CFm2lHUUoTekeo9
zoEE6Y3raIJeWLQP8Eakj16rxmkIql3fJjgnI13C/l9hhvcr+LYbJ26GURC9tGrO
9XZ2mXZojzdiskVRNtdekmDeJlBg2qPRW9e+g0NuHO6lKKFMNcD+Us2yr+4B6BiE
ZFGB+UlHbXuAoPln7XrN6Q0rlFi1913qbPDPUaADGTtCMEsPknLoVc1bqP/jyhgl
gunHIRR7+/ZsFUhqYRo7CXwIcaKc5+WsZfcK0MFkr0laj4E9lxULRSJLYby6kp9H
nzRreoCFkXFXZrFxJHaC/vh5ssM6VooQawaI4DE/hafarAvT4Od6jU9/020HxL0B
6CqGjugKrUeTYZ+2XwlVSph237eEING1XRw68r+VD5qsrq/LxMByHsqLvDjBomKm
WZfl7CJd3CzAeELY/AoHn2g/NILbAVW8Lk8teOxnr+xUT549L1mXrl069SB50/3r
D7jsg4Pg80TjH57OB5lp+A1TibXDivWTmkAQXUXylGFobPwj+gfdBy+tdVZMO+Lg
uO0NMD2Ek6d+itX2cba7cdrfEyCZwmjimk0tNLrTAeQi5EKkoBJPT2UIWLm1+tc6
/YfS3qeoBaMIKRIDim5ucjw85gnPrjkqVf2MOrJcmrPeiFRX+23AolB7Ky3Ikfvz
8PuEdQPRK6kiaGQ84ZHTN+H5Hx/BOZFEcpEJTuJX4jiqlvyN3aSjosvi+D2pm3vj
BU1Ymsz7mBboQivzjbW/ADzg1ZuPhb2Ot7cGDPk3XM7oQGZ3j5k0cLNmgpLR7Ox1
Vp1vz+E7IViPSD4WZqFFrZ5HkPYBqVuhvSoGxv2OEBqfCQPgnGkuTv5bBWjvX2FR
Hn6vta4MXcfiljrNMaZiWVyWd1dRF1lU4fWqPAlrKarCdVUBisvQUWghLOO6VDqO
hURn7ON8UtBIwRjt8ivRpBGx/a1jkP/KVfA7c7R2kUGYz702BlrNG7wDsdKu4ahw
6yMkFm+CdQb2k/LUOkp+N9x0nTUyj9nPcMk3WjbL3Z+oqPWzx2ImTMxmUiPvX0/8
Xstn/XZyEu/Th7whhj13r58TfTMqi2s7YQNk1yZM4E7YNhrJPYS0dcsMdVPIXKZ6
uJY+6X+P3nS5cvPFG/l+R+S29pbvulv4Qg0UGu42WkNKGNyMOfCloS8dJs9uL8Nf
pigsGqyIbKYQ7b5ZeC3OnxmzHtbO6sxcfm/qnsaOgnZfdsB7/hiouje2Gt6+/S2N
dzdZWFfuwd3txtigAU3dvKkXByTIFlBGpqFjYeKHKpcx4paTb3TwQmxxek7TmRhx
LVpRnL1HhT2Hhf+HhPeQhHO7DCrt/djSTf4QEFOjBEg2twzMjPFCR7fbzsk+N3ot
5GYuOLUrB+I5RoiVyWZxmWdXRCnwCRrno6ExQFOz2wMhgcjHrSd5LCQTtsx8Q+br
NCxqvJiImF/OVRv/2HEjAIRtC78k4oUobi+nco5aahy37Car9DgBw5PBunW8AcO9
VuakCuHlE32e9KQXERX5XjgWruphYb6+K5LuonU6G79ldBnHluRjTXr01Pl3TK6u
B/0QH/AQF8toGvgRmw0mNJrAzn8txygG6r5alpJ30uaeR5AMIwU3vJRyZfZW9ZKj
JOiyU/BPbbTGyZVanocYnL+9ZiqumplISN+TDxiblQ9Wp0KQ83XvZiM5zUNXIL0T
0smNUk8ayV6yW1PuMYMzTNtiJ+EvjZTx+4eTfHp3VsetfRNR6o+wzJwZZPBKcsx1
l2JgbraxEcNGeVOi5qBSiMWWnoHbq4N51vqe2S+W7MZ4iG0OYIkAVZsTw9EYgnfP
QR7+LF6w7MUNq4rof1m5qAgvfVOP4cEhL5fT3eo91Tqzsw7miYro7Pj4G2RYteSo
cF7ySEbvZ0i/IE/5lAE/FKtSUzD6HdXVv2ziYzxklzumyEjy/h/30lVu+4qZEBWY
mrG6LNfTeimidsB4PYzPXBGEkqgtcvNLA/6RW8YJSYtPoHxoTP8qrHE52lP0nO80
p1i/uvTxdfiobQmLoClgmj4kJiiJ2nUExoCrXFwgeH2CwPGALGZUrXKPUy5NBY9+
Dju0+5jsik3YquiYiytxF+bvLfksmE+e5WWXYh4XOXFeSkkdAZ8WfyTWtIW5qeep
VrmKpyCasDGH8ZhEdFTlSAqCziF6YPEqvIzZHAlA1cJI0wi2bLVFSEdgnuqV7Wwd
OZ4L3HpYRPX6/z69VYV7NwOzfT1FhNb5kekXk5clt8F1id/+Y2G+slo3Cv37m6p8
EStKz4ySo9gUEyD0f6XQXtLSsiim5rgP5UlG0OH31CNYi3dl0lE8l2oqSaR8kH94
5vQa0LwtHT4nIW1xnfNcfocPiKUR4qhVREqkjfc7dSuDdHtNqCxvvTs62QN7X79Q
HYhyFQNiE5cSa2UzGlCUNhaSq17KkbzqOd4AcxdYKZ30+LkrlvlGdRGTLj1CrmTa
ZwxCuqei2OV6D/vMmN5gWucWgi6bVYu2fnC+WmqFA/b5NEBTBSWLl69tP2HloMeq
pvXL8R4ZxBogQhOmz8t6YT5eXq5JKFxRauvKOSdmtKst6nYUkJSlgVu+r456z6pw
r1XW1cw0pLXwwktEieQ5/q2OivCj4qWQn9gMhk3/W7BDNPQhM5n3/OBEZjaH6FQ0
AViThqOoGdP3+7mJbiDfPBce1cRoj9W5RfPl4PVwm072r9WzIP7jPDSO1eItxrt/
UG+2e6FIyQxe9m4V0pAW9p8Z1szoD4OrsFWiA7jOkx4j8M8TY2T6ppkfHrkMGqSJ
AXKz4dPwEP0xCs5l8Slx4UT6Ku21vy5cwsNYtmlX/n8NtwAjM5q+NA/NwYXaqmqX
lt1P2UXafy2Y4HeLFsCJZOb84A5cyFkCqi0ub53+lh2tnL5XxVsN5LzrF54UmFGn
n9xfyreYjMG0DWdh+80RkCqz+usA9NoIaD5F/U7cMFolDowFqMsp5edD3fg87JTb
C+x6+uEhw/E5nGpfQLHQA1QtNv+TU1ZDTIdfEqcE7lBXIK9AWi1ssW43+Dm7KuMC
yTcAPdl2DxsP05SahexZUqm2J7HO2DLlfK1TC8QX9rsyot985ZBHjbQ/RBWf9K2t
1oSrqHaJOBJRA30uyuO5dGZ1NjsFTWXf8clPGs1zKa+RZsfSg2USlH+1XEQPRxIi
OsiZ1enI9OBI9uz0xobnlDNB4chYlUC4lmcF9G2I0irnCos8caA5UIk351aAje2c
aO1mBSOC7RtUjWUpfFu4s/MxiPlEbKgA5fyiJXHXQbUfR8IdXxhsOCY43dd2Yb9n
lIYghBycHWZcQsnxtCR+w5wdnY1sjEkS9h3G8yWYt/8JtA9fwU2scxtiTkaLilZI
uLJZRlpfR9nDK0qyjuN2X9DBSRArJSGie93OJXwk2XN9piyxARGCXH0Brf/1Ozha
t7f7QRFbg56f9mEQwOPsTX94cGlKP04SGGNr5cYMNIqNNJNMFIg5i8qv7/4EUkzf
hTmANh631lY+0zy/9SDkdoDz9Mfdc3Qs8eLIyVJz1l0hsMWdm6k84whkCGTBpyKi
G8F3Bk3Y+LAt6yZofUr4OeXVxiRBu5oU5zn7Osp4IkCY513hzihxdMuEWF4TKBgt
jWKARNjdyz/k5RRwfB2DS+60J+O01TiQ08ZIOsSpPS6JRzK65DSN9EfFDNRlTo59
lysU29H++oZNXqzQMpWzOKPnl8bVtcUbZOdAC35MBscWHmDIK79iQLpoBBo59bJK
fNfsTD5sEqFhNvGM+F7Iv+wiIhphc75S1ZJceYmjx38HsbsiEvKKhwPgUosk1XAE
1fvNoUNB+z42x3QVhJ8AP8Vd8VJocJAFOCi8DqclgZ5JlDoBpMPPHQ/dECO2A4Mo
kRyI7h63P0V/iRrFvoDuuu1vnRjES/8MXvHT9FTwXz6yPMGCz72kuoYYSQHtNee8
UleOS/VY20Ligz/QiFcTjf26rS3yGL8rJejMksrekADiN3ME/S5JKnRsZoG9ZgTP
u7OI7IQD4lAx7MwW9Ossj2zLqDyIFceddtWlw7FnLZ74WfKVSIcuuHr6mhmwIDT6
Kuhz4zCiPOoMzojSb6pSv8w2EedeTRTMuxVrADX8tZGvkqIGB8JeFtA82QO2bCgw
ItPm1T8Omq65Gf2OFCnhQkRCnHXQ4XvSBA7j/l84SKp7C2pMjnUJYKlM0WO2j2Ug
X8i+XN/yu/kck/6lvNBAK/w2cPxdi/aeVp5nfAFRFDkolNMTJw9pYImi9a9xRIF/
DaJi1QCEZtnwT0Jlroa7FZdDgseYs3s9ta18rjB7Xe87OhTsZTXv7kaoyONeOH9z
is5mazbyyVZbx6ilx/zrtBw8W6xYW28yfKBY7Aqje0+SSHkYR7gvkkcdYl2u2o/l
YPqmw56hG8GD3BZtdMy6xQI6Fa9sjeRBJggBA/DImoiJjE2JinBadJcb/bRXtlph
91h+cgTe2cgd2eWNM2ddI/1t2uI+0/7iK4urz//c2QvA/smf1W/F3A6p4WiyuYYu
tDNEx02svo6WWQlcdWmGklK8fWcaHf7YjGwigxvmPAhdR2gLySLFItfup23nMiNz
ZB2PWaxyNwr7Nu/yskC4bJfbliOC0zrwfoQCjxrnitSl8PIvbxRb14dT0lRSs3Rz
SLwJb8gv/1nZzbPhV5xo5N9DtKEDlTgiJ390/hS5RNfI1V1gZhfpEECmkCIgXH9u
lhSBWwtdCbX8rEnsbc5ulwRg61q38OYl3yI2y9lYNwSQhVBKRqMJ3fYZ+4XhW4Yq
G8nfOrbpuPa9KFDVCcrtk4/a0xxZO6LzPBS6AZK42FqUKCtL4EYBHHt7q4XX/QwK
nq50B3qqEf3sHv98s30SdQ7Y+MdcKH58oWMcBRzOPPSui5biVoVzWSsagDgGAH49
jXlb9vodl74ml36Boega5ZptXAXAjDrObuEQ72HotXC4Yd0VXtfvcfV1M4LPMDpP
uP0rssiRfI9l1OtkLLYvZkZgAsbYBx5vnDzBgmSUVYkfkdN9VsmmhiegXNuHs+Dl
GmlPDUycUq3OrDS6B8YZ1P1Klul4XwKOr4ekQjpa5tj5Z9u2AjPcb30ja+44O3Ln
H2pJ+KVT7UKBHSqC2GUKrJkaDJQD6Hd8jJIJsQvJSR1f3F9X3Cg0Fv3I+pnDhmjc
Dxq205P5ZfI5Z9Hs7AL1QjjpTmvV1MQcBOZ09hbGoikCIGx9DErsHK8CLx0vo7MT
hFytVry3SG5Oc2ka+sYG7CwkjzK2HkkTmntZToMbOiOKrscLsBbhaEvnk+j/28jO
sQuLh52dW+B9ep43gmFEm2/aI4W8IxxBCw9j22RW8QdYiBs7jB2fDfy23kuR5R1Z
yatdhgP7vZYX96LuvyGSFvwWNurITrNm63Iw+VvERjAqbSopp+j4jG0U2mNPoHom
eUYzFBCHbsdfXLKs59rPZ/8Y3jFqrjCVON6JCDrFxJuRMps+o3aB262+YXEw3czA
bl/MmjYkDv8WDcjLgYo3sO31q7gZzLrLr0i2I7NAPFWJE4MO9JIDINSSmj6Z1viu
bQ0RE1+5lvyYjQx8T9pwcX072Bmfv9fMvtTpK41OQz4RKCuIL61TJYOhd2p9OsB7
gK2pmP/oc118hAPjfFA55zcUnwj8cafkGyaa/8UPjvQu04KV4jBV7nfDhizjBdml
CEAznxCkvBCHNQP+YVW4zJPjqmV33vOat/xotWUUJWL0W7A7mX82Q0cwR2+kJMzf
E0NjHrqDPBVdINO7W48WDkSjX/fTDNNET0ohGQHqH4OSpAQqaEaKTp9iu6hArbIq
ODD3dpeAaXz/cYoGwcN0+Qf34gXLvkSTbqAshkzlyBj4Mb7dvoynnZj5tWl9dolu
wWTrLrRmTkaur2ju1SWVsjO01IfP+WTNW/H1dxiBuHjjilB7nh2Qe4cZJ98YdGVS
sDo//ezT4JpNjKomBYfGGbrRDnmyXvDW17m6AamFefrhcn7fwhxwDLn5hge3IpeO
yJTBS/r+fFx/dTFPTpEtZKxPbStRbCh51ww4UPQvg0waGoiMIMhVPWi6dZBn/xei
QdKQ+MbwKiqn/yqNR1hq05B4n2pFe3K4KLo+BDc7Esz0ECywpkSpqeuG02RPbn5n
OXZOkE2dgxd/9xY3ajRSO9PNDBt4YCFGVJZkOXcRghVHHMreNRlkdiKW6wHhYecJ
+dq1P62f3Ns05Pj73YaUsFceyvUjq+Ltd6jr28FCW+R1wD8DQoKXMP6x8/JQgmXu
oouDR8Wtopoxw6MT5zCnVEdjJeKahvJwxCcXDLOj1Vh4IObPGog4gDuhSOzPYNsU
tyF2EnbRaDJtWW/oaON24PHVVFTvgTqgG9V6x++HjIo4fOM4sgbCHIUnjppI3tTL
25BWE/2o8g6H6iBNf4uU0j8fXcf2M0Iq69W8ADMq5m85rCXyyzRQbCYAVSRt6m7Y
kYNe6ChX0Ufgq+gMdZaE7GPen4If6+95KgO1xDirzdCP4U/d3Uii5XtA0FfJA0gF
vDlTK3aBaBQeyO/OQlrKPzRKoRvj6gncd99jzKETEpBG/FoGkbMSdEhejzs9KlSJ
Xjmxb6jP49SieJ0LJsSKqpNEkFpqKTNddtdBeOODbP+vK78K60qK1Bl+vlMW6D2H
9xDlcPgTaX3wtTUYu7OVf3v7rBaL4++EygC4v4u61NsdGbGKIDnwuTyQyHDoIiD3
O9jqpmLxqmSS9Sn3T2Bze6YIZQj7jVS9csANFJDWgsRX+tAZTlFH8s9azwu3p72z
pyevWbRl4P5/kT5CGNDzjRXlYeEbgKszs3T/gVn+AuLac1KjdWhw0GYD3CKizz0G
5h9HK5oOFZcloTe2mLImGbGWcx6XOJL09HI4OHi0DOWEhTzftENQGoXBgcy/eV6+
dSSfJlZ7q1BXuOmylx+Ill4D/Xt3zQ5rh5cUJzts86UxmT9z0lV0jYlHw87PP8ff
k/6Coo0/LTspygXJyAzmxuvSpQq1ne24IC0LTjZuN7blxopul6+UkYrfDrN81bW5
khFpYQo5FBO1SDeATf2obS9F22Zgiccd9tprMeCjD2/Mzv4EY3/GbWOYT6rRLalu
n4WXm8B7SX/negHa1dFSp3vTqsliZT7e/tH512DRwBNVz/ImRpEax2k5dmMBf36u
BCGRUef/jL6Z3M4v+a+kQWTKlpg2gpPeSZMNKd0fmNpDZ92F+b6Jeb+EKdhEXd7u
kUveJ2m6z+MwJNeoR5du8n3bqRHlu2qMOnyAwcecrb48A28KOXPYy3NdCsMrURco
nTG2KzhewDZ3owdHsOEY2wiNhbsD24aqgg7iiW93tEyFkK0tmDzqmn600/U+MA/V
Cq4rxrMthoDC/TZqbr5Cyqb36CK5za5JkawbwfZrttd5RxiYto4qz1O1adzxgsJ9
GKLgpuiVuBEfqV20VAlLuJJAS7mCw+rWSxjB8v18Fm7Jb9tNvbzbKU/QEsRQXzme
aDb79UssTiFDfHn12F8xpt1WqGI9ZkrkDFvu3o42I0IfL+g6jV3bGY5SNO1q63UL
OebFQcSkR1Pmz2czpzx/pBdG3lqbD2FrIW4+ofRRDzFbnIEEQoYlziTfGwmnDk3l
J6Ymli66gu4IxKvuF9v19oAtOF4lab26QhSWlfMKuLcOMiveqrIqoIXRwFAJ0Vet
PqrguaCFaCXFfQDAt99Ud+Gu167le2UPTA60MqIgyXVdZyI1iyvSiiUhLT7tAruT
UFP+LCP3cYjz33zOWds34YRFt2jxhV7U5p2GwN9QhK0PNA6UkPhDCuYLm/nq67+U
a3a0OHfaxY+b8D2TltJmOUdtgntl/9c7GKHH0p/Br9XHgo4rCdn/YmL4louVh7mq
aKKB+1A/SRikF9+cJuqbM7kGbVLvtRlOPI0rdbOeB9yHAuMtqhSEofZBjHpF7e4B
53jb9horJDYW2SrM9d05LIporswACd5ed5YC0aZFHD9cemG0duXRkfNIFlLTmfIB
ZTMAF4KwVPhWikANdN3Xxv0n4gbkTGKFS5GJhfOYsWKcSba6zAUTqOhIZZ1joBoE
duy5RX1LwVqkak2IiffTNn4Lu84zhfn6YXyQ0YB/jCKKg8KD22JBl2X4ECpet5a+
3VJH7clW+cjHMcv9rESjqZ/RTxZaCzP/v/6kbCNq1Fep/CTqeXN26xO8G6jToEYI
dCvoKAMIMtbkTnv2wvfHVua2JyASF+vJrQ3utUWWAce06Var03oZUfVDRpjOvDN8
qcRfSdATcbAGw8wK6UOGR1zdYJRpoHRFhWZ1OmUMr4aiWiRyLgPRtZzEo6yyil7m
fqxBodYCc8RoKJx18+h2l7drhDOG/2uQlXJgdHmgfEVR6e/enuFod/fgje6UQDjG
BYxCQY6ocfSS50X7XpQ+MirNBHZl0so4wZk3zpHw7WtEbB8nrtGYm/J6R2bkYg2G
Pzx7n5mUPnMpnATVmM85nEU8gy3q6uKOHwIu7inUHGx7uBdWL63IMlVTpk30xGxE
F+6GMwTxuZp5PFwWNwK6RLYiToaNIhtlqI20a2AH5iggQ35LjLFISfep45pAKUr+
Jh9lzxI3S1WnrgxfKUZMPPOzgdioebGGig4UaRlAJhhT5FSPhex2xHhpK8j4Go7U
iSK89qEYkc0/Tce4w+DmvZ66bCfVSHCcN3RDoSxlAI/ktu1NjcEcfjMAVdE1Lqjv
i5wB5jHBt0aLzwIKGXDoEL7zbeNax4ofWhZ91JfPVD2JvLSt+pzOLC5aL8V28CGj
3H4RQ2SKmax1LDPkG31AVnyS/UmPUeKqqTFw0PDQAoiQKLGwjTGULqzACtaoJfSY
15o+V3IFp89cgKkXWun3SEBDO0HYjuSYRxzw6G4WdQXyx6RMChiKsQCFTAa+PnZD
mEtxRBGAqBzSsi/YgwABqeXatnDMBMOcUZ08oQxz7phk9KC1frhWzABJNXr91YTB
GPgQpCpHkFDMzTwnTKo1PFKUYoI24XIgflCbCxh8TIfGVR9Xqub57JPB+fKQrGLw
EhuBzc9Wryqzvu7/XMK3gZkIDK5V1lK1H+6Ybt5ZmRrFBQHAhrfVM+p6u1fbOjcW
SQHoQSQ5UdLhyQaw7v86XUN03VpAyt0fG4cu77k99yHIekT7VPLoKzvExBNke0Dt
`pragma protect end_protected
