// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
cH+MWoAzRZR3cXkVmFlsWVHq7g8oFtkaHH+V0tFiRxa23KJUQpHl1TDOn66ZzRwR3izePjnP0fVN
IdDtzwTdRIfcysiBHCDXDcMUXDFxb/hN1/TXMxdSf5ZiRX5D6sZjgnEQmT4jVTBdNckQURLS4LBK
z90C/3ERRIqfSiOTa44P2JF1qy7LRPdO5lD6YhggkCTvIzC9jd2MD4ct3zxZo3DHkUEJ4mWNI3bz
HkHI9XOkg8ogwVM2keTG4G/b4lWZ7gI7ch1G1H5zoPZQh9aTH5t9haQu1eFidoAmzy7H3SZul7/q
G5nfUPDYA/7+shXWS4fS/Tf8nF60wLYtUz+29w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
63l5vng/oZASMijDUJL1ny3DQMMSV8++IIG0y1PgpWuHun9+FO0819huQ+tnknOJv9U/undvk41Z
A+WCDDIe3RPv54jVBQ5RapMl6+sAJTH5AvvhWPK2Ha6izyI8H8bXHxFC3DdRThNZ/Aoj+ATJQA8g
fwTkVq2jN0FcxUKdl0t0258wyzJDU7YmZe0M13eWEYPaahddZtxCBt5Gumq43QGriIs7AQoHxD/y
8tBv0mxR17fHisO6OwlC+tG1ZiDz24j7ifNLDRl4+RYcaCpMVWTXHBZDqxA+bWi6Vc/IWCkqs89s
Nm3u7lolADCI2pgY51n3NCxg1YGGh0euq2GOMuwfIdxCLE77wTGVRrZb7o87yg9SYDXpv1elOcSh
iZS74eo/4PzDl//1HL8iJ1dCt5Yh5wOQv4slAOROAm4/68ZtQwVNTFU+UmVWby1aNl6vw7XpF2hb
YiyDNDL+vvJe6BIKnZl2bFGgt3xv8KNAuDziYyVPlhG7REwPeEvvvbjKaGT/vRKFb7HG3KakxC6z
HIS6MduWv48lax4cNDEh8jCVjcawk/NoLJLnfcDIIL1rUGntZ4mWw1eMD4t20GT5Xy8/7j/KnlnJ
ZISgr4aPKeyZYsBTR7eJ+wDCQc9TFQiEb4jordJJi+laxg4LLSi6NvGdeCjPOfXrsZu5EkZfmeFG
ecpgx0VpoputPXS2TjoboRjC7w9LG310JQxKY07LBxX2N3egErJ898jWIGsUR38yN+BY9cfQnKLs
PA3vpo4xdQSBwVzihLRvJ9Gfg+rWte0ZAJQsGoSAP8DBM2XB7k+wn9otR45CQiXTqeJts1BfC6Se
ySyiKA0hq6jq8PuQyZdjeo2VkCfoR8kVjdLjD2iZZ90YS/dLUiySAGpL7eUBTzVk7UFbapoOLSW1
EX74qhb37sSbkTrAXvd3fywp2GqJFok3wDNG6XmmH3HrYnguGZavwR9+dGr4bDowkPJoS71w0GTa
z88kQQO62HJf9mcX2KJEZQh6O/Fq23R+vMu/reC3CYsgpBhJ9OoQRxw2bYAV0AWQo+eKzoNg7bBv
GWqmqOL8gcLZ5a79gIVpbwGxyqq6ouUaaGYVRjgYjXvLSvc3SajN4cf2uUoYX5lvrynmxFMIKHyT
rNyr+53e9Mi142VWvpzE8RkF6RR8zA66Z6t6mul0VhzK9e0i5sl29uSpRFIT7RFhERwOLMlJR4wE
79CEjyQ0KuOMqDORqdxKkujG1qTLg+DSWwwelTjg4M9jmLHASUe5uAJCKLCgRalx0mwEuoKxyjwe
9QJg2w7t9/Qrblv7D+DyLR8q+yI/yx+0CuzYB7b0Fiz/c+bg+87isn0YQ5d56kxkjU+HNt6MealX
scsmwwwlXh0fnNJuWCCpBAIE8NUq+jdxFDKargRgkDTpcHEpaT5j1K1j5/1mpe6ClsWdZSssfYM5
BhR1rL+mGkBywCwBOpnx/GRlFhuFmE553uFjOVBeDs87jJkqRy37O5LvGHCFukvD6JFXu9aLxQnG
+sXPEKmHNk61z9y8+94QNm2KLT8ZZILBfFxDCfW+cuTd6htB5C62zRPFgoR84Ck51iMKU28+TmDy
1wOI1LtQYVkxK/9EBhNgnQpbxoHGtbX+1O1enjgH9+RXAPfxH8SMTcpld97ybfQWQJurFIaX6r3q
ZQKaWtsSbQCJfRijBZKf/Hydb/m5mf6F8z8AOFWaV4rvsNcZlr453tHBHj2WgJ/SZ7E1gBcZKhG5
SSqg9lp891ahHN3RjWBvQ3zYLVjztB94PYZYCmF2jvonlzA5uwqH36Z64fGG93P0aQCbk1WDuSR4
XtVN3P7ry098GwUth5Ull5SvPUoWlEJqt6dW9pbJvM4sEtVSX/1uLN7snBXj4XKqWPNV88bnkZql
rnXVTBtAqbXR7CtLlXdRFhc2Z5HzyR6Oi4wGPZvw/NchiN7/oJakymLkZsvk15SHTx2pUea1fpfg
JCGHiL0aU85HycVffrVCtP1dvZSjkiIMumrKozYtH1TD/SJjmBGSmCIf8kdFWsnYQjJik0l57xfs
x6FJJxjGW5gc4c/kVaJE+txaM0BHjh3+iXg5RLtIBRpajEyzsZoIt9Na4sfR+La+7QSomk4tmLcx
WB9WaROI/QpFvskGlDDRhyaFBfPPspuQlNwxxifOgXcB/SN+nZ/1JQm3XLkEan4JBsZ2y2rZeTOP
D017PsqhiwqsSkIHfJhOzq8HsPxEW4oK3Z/TTE4KFJFp/bC3nch5wVGj1Hyg3RsPC69EceC/2+zs
V8aEWvgrBuheg1e/tyPjw+FlKBSvu+kgdUc/4DgrE0/6wb1PcUjBdR8XugehiUgdqg/gv/wmZFOp
Ky+vF/WhDI2h9XehibGq0HGGEDD+TXTwLh+Xf0oG3QpnHboBy4LuSv/cyf7d7L0xh8GGr+zr7FZC
VjVu/XKiWthNfHnZrv3qijZMOGs+NYs0/++yrNGvNIUzC6JE49c/ohSWmjn+72p9svicNR67FUJ9
IdfFLvoM0OaLc45ujGxDg4NpjkYGgzKz1qk3pCo2bXVXncBGoBSRyeFYT5N7ofdsLGDQefz8s05S
BgPv+Q2fipmyLoz17SSSmQY7ucdTh009yijveA05WSzmeVIvw4u+JbAPeqGq6EekCD9zg6j/F3hq
4uOOZpevYIObQejd9HkI+2Hce4rxFp7w0ocyJSsA6qPUGTcsC9u5OD9b1lNJjwt28CTflqAAedLj
Isf0EBHclz0ujA+Bo8Bx/VDj0sNjTZp6Tw3PQLDeyEWCirM2sVImz6UTdK7cJwHsyQlrltu1iOoj
mqYbWc3p+MFfUZYp0edjqnTQFw04mNxWvqtBU4OxvTZ8Go+SfD50V45k8J6jWiaQYW5PGZRs2ti9
ERoE6WSNMyecm1d9qt2WFt3T1cLt10GM5W2HBQNb0YKvudERmtI+GkBMJ3OZlVjDRp4uO2uYHpkf
N3Ms13w5MjjqTIwIQCyzblR6qFoq5uHkC4xb1RdOYjZgfF+oO32h0x12lZWVyH9VwmgFEEIYrF1t
QFft5wjjQ5OehIDURvCeEjhvrXZs6DGx/V7zmlHR14icbG57bIvHBhLXH0UtW+jwSGcF/uWNdcik
7hrTEnUyUxRIFgZotKgNfBUmXBWkY1Vx7M/6jAVthxXAiJR2O9zdBzqNs0eEtPqfWd6JvUd+tsvU
NXaG3s2XnkXzgWHmC+pjDZr61xb0p333w0nY0vcEJnX3bOL6q77y81m25EQJmJklcZIbscDjxL+M
mJoQkawXXylgOP+yw/UR3tHcrYbW3vTHdGM39wkY6qfLBcWQVqkzzDPVzDzBQR4aQrotCITc+ARR
VOrSM88vRF/GwvjOSgMG36M2VFb4or59FMOvGPPP3ONPxu3eLVhUduwnc9s2oDRfDA8JlcU7EoaK
/Ko5lAS6COxaXkCyAr7V/lr/4DIu39FgUoyLsWoYwVxYDYCjNYkqrSKnzpLdYhMAW8ijpPJKolan
LEozmDXlhS6KMzqmNL0XaRpVfyoxD5H9kL4ut9X85TM/IS8N3ED/qzzuPXbcuL3D1hw1lClUFQlO
wDanGSX1VXhxHz674uZIt1DljjpsOg6bcy/u78+BrpBUiC5U83I6GmmvziYxq3xLxe3UV0dPkTPT
+yna9NGvMnd9Mek4LXLJkQ+KcroANTUyv0i2Nvhx1hDg15AxQVM87HzK8kVrGBG6Wds+1V5q010J
6zBI3EwFA8vR/biALMNg9hDC/3IgjN72QDlD3paNMWSKrJLnwGbqgQY0jo5N2m/4xCRfupv50NsU
mLTeJJoeOG5mfMhaJarLG8gqr93x6sw3bEdDQ8assZ3bLhnh+zHzv3IbCgYzo4GdII+zTNfobsPf
tPNbei/FNGwC7czbjuehoNpRqlbik01RKb4lcOlcY/FilF+3+CKM8IzkR3IAZIpLv9Dx1iAHvDS2
4O2aJm/PTOoU4GW3FQcRiw9nY4QIETSMb5hCRJ3jQed79zLNZR8POSvNl0GA6hzx7sGnU83+ucuy
trDXjUCOiunNBy4fGCLRKzLMlbOtJNHM1uOE+f+hwtRDkWxICMZSJ9WBVMyRj9eG2dzrJqiYVbg9
o4FxmQCAOsDhsZTbZOYAoasCd+z/nAvrfiBVOkcfuY2UUN/l5NcEe+TABZRmBFIZdIUxIY2PNJAs
Tzbiqksxk6XRd2azpJcF+5bW/d+dyJ0StYFmW6izViIKoquyoNwDZ9d8DKX8tJeoXk42EieofuGY
Qxamh9HF7LEJvlgH4LKU6I1lWxxMnnLCcWZN22wo9s6bGpBc3CHt4fWRFaTiznqotpOyBWKmHAzZ
aoI2yl4103WkVhfhu56fV2/LE7x94yFqylJg62IeU8yJhMd1UVW0VkHArV4BvTBnZ36QVznD7U0V
z3xShCbubk/Y3pDBA/T7pXvSFggoQGt7hgKagOh3EOLF/6pPAHPpNUKnhA4rzS3QWrl7yy932WvE
mV9AMu6ET7CjR3gOorVr6Pvt+w+0phgurMeoREf94HDe3abV7drcKs8C8WYT7bWFSm+kNKBdSLVM
S2A+DpJPMG9zv1jmNS4yNjaq64SP9EOtU92fBMNtyyxSi9kfld5qWCdo9U0ZkNz6X8YTm53D/U+g
aYSbXTFnP0Y7fqlv6gu2tCQhJ2WbG+I4BGl/hoAtn7HcYWbFHv2EEVplmgpdu1NSqgTC9NVBsoiE
vC8IG8d8LZZ66EYPKPVInCQXxNdAi4aEuvRKMeDa00qXUK8udk10dw4hLhu4TRan0mZpCENzhsrA
f6K5uWgFt8pNAZyJf/2xGhvR0FDMyvX6Fs9kQOVW6xPSg2tV5tyQf0efqxe/rI5owo55wisAPm3Z
ZB78TB/L5sW8lo9vI4NWmCJea9GSpksWpa9x9a2ruLc8lELov3p2NhpCma9ipYQ6kEq3nGwQyPml
T/JMbPs+IT14PE5nt/XeDSAzdckbxQmh0kAya6xWFYUncYBa61LckQHlJUN2+kqDe9UHBKVrvFxc
S12j+Xtc+5Uh+iBYZdx4+sET9HK/92bVou/0zNzQ7KD2GNS6Ge4T5Z57bVXfrcj01LCIW9rhE/AB
DQ/Z6tLHbZMkI73fb8Xzh+u6MDp0uFlxC17+8DbVQlLO7cm3QrnmC92TGhCtOTyGH27TwPzpfRh3
8bzoVvVXcp4EDLmIohoB3a+BfPeZujQecCf/5fM4lqxChX8qT+7yvogSCCybtxEx77aWq9+ZKikf
Nho5dnRbxWyonOmWyM+Joc2Ko9VqHEHhn3VyrgRtLiGmXSn+5UEWJZofUlrifzXMD+Nv9vwjN+hC
lrUyWsUlZJHKmCOegp2g3TUASuz+1NQnDP/vRJd0aZNaytLIHdUaa8iKQ3XUvlh3+6Nqdogtu85H
XrGmmah6WxGUWK0B4QoH4ZHXTne5NSqW7n84+p18qLd1Xkv/RJzFxcAhxmev6sk/tNoVGBkuOWte
7l4NYvxwZk/BiYlqZiIql7v/Vcuu71E4P4n2Uzm7zpdO6h3KRC/1sKrfUK9LhlLHo6Zwb2uBj4NR
I7D989TJuqS0nYql3CxUnhdx1DKhBuqJXKx9GO7y2opy1kMbC6cr+nd9fHfHs2QJoQB+JGrQHkVY
wSJDnRtDxsq/OY1V9vhK3CrQTktPwEsTZDw7/ykaYVJGELFAfk6BCiNiShajKcHYP2ZsI1FJsOO9
jq0hqGd7E62L1Mcl97VasGZiYGa6JBOCoDsQGX3sSVj3S+GUhWz1hOuIyiYBXEHiM0mQ09VJqDi3
i6G+6odIg28DcbKAvsw5dgyxzpSUIhX+0o2Qj/KvU9C8t24gbxrHegNyyh1KjSjMpo8U7g6x+NuR
qehjWB1lPLJ/zdmoWvdsLVyjhbLkhNNnYDBisdud3TP0Uh+/xex/Gw+0tO2bYgBll274kuH1nvQt
pjGLdT0Ie3CXVRwXeBYNbcse01U4PpVSKlLe9BRC6RrP6aYzgt5SAOixdQOK/CdpxweTV5KwDn5Z
8l/hcZB7VFWeI/8VRqNgQ5qXuZt17YADt3dbjrZcz4Rwh0d5wU3d4xeOArChTpnAD2dx5Bh9cxFI
l0eHcAchfeqo9jz+lu/EG/6GM7iIYaVHlWTj9XO4RACyX9+KLFpyLq83hY5oLWVW/KF6dCLKTlNW
5ZNH9YnxO75WEz6jOcGbRbqoT61CjFonayH1+CXmSwJJ+HPI2S8orHbuukB/j61uJbCIxM4L58kb
YbNM3Uj+Rab80pnTflMcYWyumkNZGSBSs8jG8mxI4XQFG4jcth5K9+hoOEOAE8u1z8rMLYqVx5u9
YdpkXBpi6mOSiVh+dFm978WUDxticVybJ4xDzUglDRaO0fXEIo8P1oYwMEprXfkK94re4uTNoElq
XGou3ZamAhs+sApcmEZgLknwT7m6rilXl1veijnW4GOffKaMWpFXZLWI/E6PJjJUntVB7qhru+v4
HOF9TeBFiJa+pMOdmR6XPARG4sKi+XNvcfhLN8ZcnT65ubhm5imgotqoooO7H6EIN6iYMkH3hgkp
+8M8Drw4Oe4PDW9uF+VN7bu/S8Bxw2bb/5+Se7mHawiouYZev1CXJ6GPmENKq+QELFc0TKEOEQPS
gV71sJqID3PKuImlg7yyZD1cZNuHmSKUVQcV6Cm51D7bwMY2Muq4ZUIN844LVBrEFOYXgzpFUFa4
CmBVpLIl9gwV5m3eDACRC6VR7fDBZbOdPBGhwY02YjcXVQeWmUL2P2qkOrVBx1nSzne7HTpznX7P
7kIb72YPeCtBr7dVI9EV9A2SnYum2OcC+63QuGI07Hfw57gM98S3Oc2E2QlLPvNBUn6aQEy8ZoVY
V6NtDkgTERZcRxbBfXJfi/qXYETM6zLr8o2pbUuYrMEgQ0mh7im3YfjeSDx259oOWVW6YGU3V3s/
L8fPjxuEo++WDv7WQPZ8EZQK0fHYEoCuXP1yX0XrY2bH7CNTG+MSipsZu3CKo6ICWlOy9fuJL4Hi
4yayOw8z50eMEvmM6f8Vj9ordmK8uQ9Ar+vitC/KFX+zKB3uTr3nuzoZlMFcnyH3Q+peu8ueYA2V
wNB0EZmVhqPcZXhjpol1bDWVQqAHD8UfjVXRNu0PId9u4ruelbtSLjqilyUwv7Dqvr4fZUEayqGY
h0O3OaXtTOq/NHZBtYWJULpQFgfBbw60bWjnarNeZCBUBirQpge0rXHnyDzL6sDLidCibT+Pz+qU
I1wVdjyWNkWtoLbneYvwmSKBz+sXz7/aAP0gS6dbrrLKV9f0cSG3dwUNcSHsQy4KmtKGkz42MOJc
EIuYfB40BiQGLdCQmw4cL9IH0LZS88kw1oyRdDm15+i4DbwQuiXJrTBcBwLd/R2DH2VOAeiOaYXh
tGYh0kBfYWn7cs7TXr9o5J6YFUbYWbWHJlEElNqJ0bWxc1mBHsNUgj/imQbgf7F8bsTrgFkzfgWi
05PdGkod92FEMDB1FTfVhxZf+oOn3Hgeu8sJwQ2NSQHdJfuzv5Y89sITzl1gEXcHx00oiaKemg1u
6JbLFq7rOPs+iW93hIm5T9QEG7HjDtNgmvE3XY3shrvAte3w3/jElAN2/xiFPQRU5TiAhuuUzk/i
ziUzrDFs1SnIdajBbY4mQoULfTLQodHgLcNgCowbZ49jor+U+bhlc44BioW9+LLQr0Oe6RvY0WVt
0oV5lk91zNu2l1le77uKV7wRmtBgcYk2X1b2PXD5wUoY602yRhIlvYgwAsQMsaUNTl1Aj2j8w+9m
XK0rbCe4OS+FFW6TnNRzfSiTeFKr+kgQvumiy6Xw0lsdGIeVaEeKfAWfGKulrkSP8nJYBYV+7tCO
4nEow3fYrMinmHsFLebeWQEvNhao03BxHbxCj6FHUyOAHUyZ1Jo/4CInDIC3kJ97w2WlOzwwSEUI
2c+duluR03zq0lEbRLOkAqGzHIMUoMu+q6GYcf+MuEahb1PSuNb14Okljbl2uHnoc9DGbT3bqzi9
ukW4vBGYhzSn3T1RNJzBoDQh9SOnQVQZDNvBYqAZlXoj+7zJp9W+6E2OOG79RPJJtndkQzHqj783
/INO2a59Y8r9kP8/zfIT8D7KLDv/04zJKSF437pat4OWvYilk0/xxGZtar9aDyFnJh87ehDBotx4
pKiieuBbKlpqTFJei/aOrWlvj59m53xri8AZiZDf6dGlI1muXW+H5l4lNxmiYpav1agUFVhdYN3y
aMH1SOUghTeo6ZO52CaBZ6+dccErW4ZZEfw1GQb59WVxPaQapSK24GOlqn/EGqx+4oz0xgjJc9Fn
V0oTxE0ck7KWSllE35uX8/dMEPknvO7OaGhwC24+MNwWkL3Pn/6LldC6U3hwBUdZKXR7JSKSiGar
2RFKW6oablKb4SwRUes5GZGJOhDMuqgnNqwRaf840V8i0fIIxL5u1UWPQfv2RUWCZohXmLr2oTQn
379froG2yR/4i1O7l+mahCEvIEw+LGktUSJ0t2SYYKkQldpzi7dzFrV/rwdI+U3rtquf4fgf0+us
c8dZOBvbOy1pvlU9dsoxCvexKvTqaaWrrjFA1lE+vlkIktG1s2u4b0qNHbhgrybzzioH53+SElu5
JZzdUY3rPIwZF7nhsQfoGa1jnI9Ga8QuwCqHr8k6UbmUn9zgjXGM2HkEQmKqdc8tk5gkQFLdKQXl
nQABdEfCMoZKjZl5I4YXTw8TG1vV5KA60Y44JGNSxFPj6G/ikYaEe2sGl1UPOwh91sHfC5cZ06Ch
FXXzhToX0jAIsBpXKvE4Wm2+1JdRpogCg5sJoxWTJ5w+km1azMFf1AXwCV5xF9Mg4wqR88oOdM1m
rylB5X7HNmn4JkxFuW/q+zLs81yqZzUvdSEnMD5/dAC0gCFwpPovKWezknsp72ZWdkzYFcZqgvLy
SReOojkxh/kxcKGLc6w8SMcim0L95hkGo2phubZ3W+nQzwshjlK7Nfg8Gp9FmRgHYirNuLjgcYLc
xjQMtg8HSeKG6SXwvTdv9x5lZYMXoMuRYYeNPNFrouOXQiQoYUa7+SMpn2cpTzccgIw/73wfzwHP
yJr2JPxxSu3c6iH5I65mtoBIMPF8Hxit0f0IikCbSnOs0g2+DczzcyBeY3Mt1RlEW/lMeLHKXiuJ
sWdSYFffuW3KVcEn4sxt9p6JV5L89V62oGyW3WqBFfKt5vQmzAMRKpzbr6Rr0ZAZKpQFZPxUdKcg
tRBwRO/uh0fVcJ+9OnNZ4MtCSDgImUFcjQfEcDBDL/Qm39kl6u2FvIdFjfRQSBS59VJx/B1S7Cbw
ZrIeS0Zlj5oboJtAB9uw4/kaLO2Noxq8vQJVDVQSjUpLXJc0SFqabYuTzSIX5+m5UQOLv4WBpcKe
b31KnpHtTNrRVoiwK28jwamX3cqEqFvlqpzXKIcGQtX3HgwnQPPPZKxEBfncvxhr6RrLCqbvcfJv
hRA14GBirab/MlRU6gJAyExTdRgLaINyErtkJ+6x7xM0yPXchRDqAdm6FPCGAiQkBONPvPx7IYde
6HbRpvMurTveC4is3kWxPCDHj8KlYv0pxyAmWbD4EcYpAygUlkTYBA6Tzj+g/IbYgXDXZUzahoE2
k4yrZCT6z0NKYxvGq9CTtAhDbaDxOHQjcTlhp0E17yqEFCCF7yR+j2BIcZPedrGmTfs/BJD3lanf
GKYQaTWmpdVh+Cz8UrHdlpu5VGz5wx0kpIdzH9Y86NopAAGQPymb3Y0OokOx3iI5fnnUtPJhYdRw
OjSC6XNbfbdemEf/WBe/fjJjj6bwhh7eJca983iYYxBQf9FeCsCwUjySHRwmdqOtxrQD63Z3xVjn
Z6sXp8JmrrxoZ72EcrcesOUsb8N9ogtSqU45kURBYUpOPqJZmvNB2/wJ0NFvKYwZ0/TqzI/DQBjY
PKtIegJIwsDy+EXI6yM4sHm0XDen7Ny4w92eavUFWfVC16yH8GSJGRPX8X7qBKDlADMdQMNbO3Mt
qPSFjHJj0EHEL1ptuy+rB7vhInBDOvsyQISyW7CMzFJkcIkpvxCtlqP8rjg3hyREXnxYcIqHWHb+
GfmPU374zr6mS8fl5i9x+d5abu5Rgqkw1D8Df3jbgCRngTwr3vqozI4vKfi8Qx/IkJOSwX/96NUD
Nv1/9GfGFHHC4dIbJf2y885tymTcH4kNjYm8FsFIO/yagDdnETW0FTzPArtqSlNwniQs7LCPiaH6
mD+Bt+uEQVm8OlLaE7XksezfniJiSDz0VHYR+csxShGlYd36RGinY1B66CmXc3mW+2iXYI/rjZ6t
r8pBBZe83C3/LCxgTZuS/qddtnCBKBiMKAoP4lZzUntGMFa3cM81b+oU+i7UUMOPiZddPOLa3PEB
s6RKY/Fd6YCyWwGOXNKIoQraDcFKxRKwaQR1Llj+ExHTcIru9acAZT1ipQin3yv2995Id5RLe6Kq
v9ryt57qVSK+x3DAcLR1bxnYxKAvVj/xSrAXTZErGa3NIQ1vO4BSr2Fl/X7Fs0NqxbOmpOC7yntn
xO+BpxPbHmXfd6L5Gasb5M3ZOQZyKQpC28tGFnA2rNTmfn1f+BDRq3qVD9PAvPxETg1jzigLkm55
rkpLM/e272+o9ST8KNrtV4l2dFi5FwaeFOqVz20jTRO19YS4tLjFSSdEH7+dpvKKtSxy3UAiUJe1
zqnPZOPbFBfqxZNDq5YMo64WG8I/92V0A0rIcJjy2ldbpHzdlBsZs51EXYAS+RO9V9iyLKjzdITS
WE5NyXeiAJgcRw1d3rBEGbMpOAHMs0mLXr8NsjfYRFzS9glfNTDTKlO2vhn0NUhi5N0khDldJ5yK
L/5nTq3CDvkRSq+t0REAsCbvurmUJCUSMXvA2QQDgPO39Rmx2hA2BkCT+E06ahw2pAgBnBJzGVkM
nUoS1porHCDdrvemtByIGA2l4PAQwdyd7/CHXw4lLxAp6Dht2Z7sIy2LOQ7QugmjtN3mqraEKklM
RxCihK3C+633v+tBefDwnKilMMjiXebvuZlPJRY1+x5InTgOUJ+PtRi8EsbYMFU/xlbL3GFNPC4T
LgX8zNIUGoStU4CcpdmnW/Wa/HmfqYYKEU9y44HPPHdeB6VLHnpOr0Vj3HOG0bGqpEiHDMCoMWzV
kBbuVCl+t9mxUxxry5k4ofuytv1iK1j8om84o9e5NUjq2YRtVc8Ni5Fz3dNU9gqLQAfeOEeCkr0G
rAbfYnUcw2tu8L41t0amhKRVI7if+Wm8AJMGhXQHO/yC9ejSt89n9VYMQmlH1+pClNeSfAp2cUEo
qDwWOjgB8gz22ORmRzdPBalDIRvcVgIy3+nyJOFQVpwhb6kyrFk+pPMniwCVa4JH9R/91JsnbGQ7
+AtwELDL2GIrGfnTjzrX1litaE+IMPmgZo6eTF2W1KWbpIYhBL7NrqwFo7fdvksQadLvxCAPVod4
KUsBRs0yPbjs3DAnRAToTTNIorCguyofB9i9MCygMO8WjuiEFCvdn51OcvuIHeBux4KapSqpr2mm
chCQlPS46J9/ysy4JH8eC2pOnRWGZ5EDXtNfXCO4Y7VMU6Z9jo08VIcOZbUZg26H0wkjSU1ZTXo6
rmB9HtLiRNL+KHecQATlFfmza16+4G653cc4QSgH5xADGHOYL2P80IAzmWqnghFjI2aIbNwu4zWw
1rXP/OcvYHIT6lAuY2ygFth/kA3Dnz5FWLgGou76XqYslWb28Jutw4rzVNQ13r/6x96qwIoPCJNO
IlKoZb1qMlhKBtJw2C0RCV7GzPUxhLeYSMx7dT2gyQ0jA3hUQYa0UJZv4yqG89ltSlKEyVsuRCdg
EEQrit+Yo91HjEJdx+1ACOqpRpo45Q6iHcZljGfIkOnRoblaBfdFGErqal3zCbuMuFcRcXl0AQYk
+K6RhkM3WZ1dDgGYz7AdDbvKVbutgLL358pZHve2VzWkzEXMJjbdGu31Gy/VZasayIR3vKe0S1aX
BWfscIFalGJCMTG6EHUEPPPcRZgaxhdkXru0pC94aylOwtOK9bmiaOZjTJ18oPXBkwgpVO+LDBrS
soWGAaPfKZrFNXvNgqGYsDAMKSUATXI1Srp/6Gf4t2OI0bVG2N+tXBh9k1nkAuanHP2YUv7zJhFR
nsPAPgOUGGkkc9URlARQ9Yk6GXgWuQPJ7MFh8qKD56mmThmgMhG4CurDdYKDkD5ccNIrEDITWDzm
nIAFAXlLr/oVP0xjYgWShkLgW7NHGv0gNsNQUnoGDCWROEEKFqf7TCDDY+hG5IpuCrIPvJ97saaQ
fxorz3gsQZhpzbmiNL18iUqgqgASz4/BQyzGmuokvJTEyQf8oGcVokJUjkKzu9V5TIpGOFmS+sdh
H20KWxj44beXEbdV/0tJNF3KY1ifhOJmT4lX1fCmsCr7ph7LQsU6AjhRlsOnKXgWBhqpBE8S6oez
fRjxqr6cJVm8TxE0ZIAha7dQXCVsOb1SHnvSQ5TvCgAjnO4tyezx2PGuwpidVeRcZ7x+6SKwyxP/
iDDZeA4k10oNBAgurnR8HgmI259Z1V/1Xse/9uJPiKgbaYyw0IfXYaRuGBiTAlM073IeppZD8C/O
ga/rfyqSBWzh1D8vkolDmA7rR7c0olSDMOugT0KrRcr3UflQl8aLig2Wam+v6vpHnsTYMEDL3huV
3SusL5YlcvGGQm3IDIvW+KjS2fzDJyQxFWhxa/Ch8+daNPS/9JGS+hDAns3jsvtHgQ2pQjUSlS9l
omw50iyn830zP7kVYt9ULyq0VNjjFlBgGll5hvCj+AQuM0HKLpYnNB+0J8DKQCi+OfJEeQveu8HV
//jymsrBrp8tKU4+4ew+ihpwnwocTKZdsFFEekWsOLqmW7UorzvTJ+ACUjKr1OZtSL5BoJfT2Fga
1D2tnS79j6ezl58Ku7PiKXo6hKXkTBcc6Grf4Quy53eLjbHQq2x6n1EGcPKiSJIxViVVlC4iVCGG
Jw1yXg2Mw457G97fKslzjj7gMLt1URIw/hJL1bS0oYV9FF0CbjTde7Y2nAzK9xpPDh1pLhOVCLgH
KF451DTg47vpeLEGtlh0JKrWR3ateTvk7fW6+H21nAQYcYcxN/7FWShmS8HMWw6mo5wekC60+i4o
dTHLfLKQnBmWLK2HvnkdhLquH+K4Ja/ue95Hki2B+7KOefTPL5ULLbnlSeN8qIi/1ljGYFBTQD1i
rK25EFOABlHAcTv+0a6wwAXphKBoIkibmzAb2W48yAtk/nJnm7Y20kCL2K0DAa+d7AOGsQ9WePqF
CGU55zx1k3aAbYuCffhX6gKC4in1EZQUtwnFJqvGtXfJYV5NIyQmF/NsN6Me5vqnElp9kJvUzdrU
VKNruJvP+342RsK8BhTh3h+LQFwp70pA7c24tpVDJpsRbaF5PsXIV5+ilOwui7aHFTrTq3/NkfmL
bGkTzThffkONgzUtX5jPKwdefLGzy9rf40WNfh81+qb6HPeIjOO9uqlP+ldpvVUZhvF50Pu5Jcob
tC7YiC/8VZPPWz4YYAqwUevsSsbTDCRL7rW99e30uKrdEvxa81L9HpiMsG+hdJMAh8eWrgQ38dr9
IP0Yh6HAbO/sbcFIptdVmXaP0s2Jll0xtzSnqzv5ixmQSMAw5H929igVYNwnGHO0uUi/43M738N6
q/dIcNlzqOwo1fWSMBCw1GwWqpS6F9YR0KIUCfWQUpTMIUzDQ4r2uGjMq3u8m4woGoMfnX2Tx1sS
GhQoJZ3OqmLJxu2nC2mcvyc6Fkh8kEgFmN0BU9IeZ4sZindoEm/tHFo9yQDkJNzFfYRK31wswoem
GGUNNcfekNVDegD3VfhpFCRQnqCmfe1kXk8FXsBSTZL7CUnhYnHegpWYlxQjyKBvG5vGwvBnv72v
XUWlAtByUJeyUwnpoe6fDt6fXo9ECbe5iQhFXZMLsDrjTI/kKBqc4Ps/RNJz478KjDz/N9YT8geG
WN1nLKHiuXRbox+RBbE6B8L4XpRzYLTNwJqSsYtFrAkMnQ+hQBd1mtJlHCQZEU9OO9IcI+Xe4Q0z
sqy32UreSYaky5b/imG0bcfjV09TG+yh8Yl3hr+JlePwLKaBV7SlIloiu4KLYbyQ4Bz8uYhtA8mJ
bsAvhAHT9pJ4p2ujLgSDTzNvjZaZZn0Dqqepetxb1HKy8BVgT7GYKTuGsmvo7vdl7gbP0yxiTncX
lyIBXJ5u7N2A7iRqmWJ2YbVttK/KQ5BSOrrkDCmTq74g5Puz/F6JanmPyNt7Bqs4hlThOb4dB3kQ
1qHTKkqPpA6HJp9KSetX2MuHZqsO3eQo9rO4ifUqp3DOqhWiKK0Js8mWqBg8GHjoYDDVU9O0R+hS
mMtDzHpIF08WLppOXCKflWJVSKJ0+PZyB3KZi1Ry3PFN3qT3dH5hq/fNi52rctMsAxAo4m7fbcZN
Fvn5UtCF8wopfyfc+D7bDh4J3XNReXoOP//ytKpQbsQmp5oGzgVeHdtIzTdlfljjeT++G2Q5nAgq
w+uMAnVl1XMxkU0djERPO7vW2z8Sar9bEaRMc5dOudF2XLtLayFjTBPsjCLqu9Gdi7uFSFfspR0y
EKeQI/l5FQ7cEHTnITiEpVkkr2a3YB8JvS9g0hrSkWVhjMR5ReUON01KR5ODT9G+WYU28I+XTDoj
QEh2/8UU/S7qbkC3FhUPVDN2EguEV2H5O4c4VNs9kXD4+yy7h2DEBaT+Lmoe8RbNUJLSkGhHU34Z
fxWqoP06KtFqfAh+VYBLqBAfe+LQ/cFElCcrJO3sz0NkGh4yfjmZhe6pUoKArEXz0Z5DFgehnrMx
vefsc/Zhp1vf6WTRlaOjRRhMoedkcDVNI7MoFqhr2XGDhy2wxk3emc/p1YoIubwPpEwzlRcJZJyE
H/HekSam0LodOT+amR76WufMs60AFNTnpyemde4BbRe5rd66WSMr9ZnlWnuZ8EDhMWtkzQdHkkJZ
MLnXneQLk8PTSZ9/nCjmAvhF7funjoQSF/5ptaCe5BeO2OLnyo+bwCXbYlI8YRpIL5XQ/QMa9m2Q
xFAmW8YxhwbtLyqsmHeBWqEJizRGFZqcNPcfkcDQmfvh8l+gh78jnS5SnP/lXCXCwUEMmdc62pT4
n6gKj8kqhL9cKqG8dE9nVEnNP4eD5GiLC+lhKQhOLUD+RZHWWgoChuWcAtPU/NgUsoEUE2Jdu1J9
xPdTd5Vjj32uA+yHMv7T2QU9in8Bo06IJwmJu/H+3ypFqWKVr1gTk/c8fgNHQ0ucfus6gWohtnCx
JLgkAJZDxDswJCl8FHAzbsRkkIl3TkU61hkl5FGFfu44t2yU13Keaj1yVEC5y3SjWNWuTydyp1OW
oktTIVPBs2gPEWNQ+DJHhIs9T6wuc2+P6Dsp7IMvQPRteFwt0P0sOyx+G3bzXd7IPMHAVvj3N0hz
518o5EJdXCa8gY88EllQ1xYdR7jbQNSAaKGijRwxaV0M/Sbpv5HYNhBWl/AsD3pMWzghyQCYlff9
YSpSbUBqbvwSoKgOHvZ7p6baCRGF+gsxoKP8fykvlSDEsTOoYhOM5RRod/ZEQU6kxogx8x9cqkTh
7vcxAAYhzPISMBLcus+AT1qjMC5kE7P0L0iGCn7VwH8mWlQdwfclsMEkoiIm5jQZ+EIhO2y7Esxu
VAFDzJc+lXutnBOghT7/VfaxOkkTkGds2m3Gb7Yf3qsIvSd3K5gn23TVB/iGuTiWzK3PriWahuSP
Qy8xIrkUCyT6L3VrA2wAsnwcpQyxBWdgXMVHEtJSYwAEVkhrv6MaetQM2tfBjET4MGF3n/MkuYiB
uw83TVLSqpfFz488vJHvAsWmHLTGDncxQFO2kG9Nu6jsfyg3WVxODCh8lPCw3XgK0svBT0/LwxsY
9ufDhTZygAJO2nM4M3vT7pMOwgjpRMekU7Zoz4vEPlAyPYv97wNLBnLcdPZcRCPjKsjzdNnn87vJ
wyVLjPd3UJ133BZMJqrgRFKTLQctKcYm9LrcvAcaOxjZcYE1ZQ+IHQb4zdjnG8T1hjYBv7tIipWf
PzqS/PM5nlDKdrzZoHDUmRar66Ga9gexkZtsyL0hrRDfz3/UaqYq2CHEw0/qOuH5RHkeNd6+Z15H
oGd0GGIYFXEpSDbM0PAA70FmiB6Uq89YyvT4SxwE5xC41pAv3kYddIwF4h7EEGPiLSMqcB75pbAP
MKUsRbUWOcNd2s8T2NSuy1nUjfEKx5sbh+bZXESIKxLXJ0JlGoiBueOVhkh0ySdaxpNxtGnj2UKg
imxbpieoSupzsidP43GVADmr2Xu26NDd83wFEa2JnVhA2SKM3MY16Zb8ExNTvFWBg3+rNczXA41o
QHM6qeRGGA9AOutAB99GhTngF9s7rXKsdyuwTAS2fkQbVfEXU7iwBztnF51kUqBuH9MebQ+xrhYR
oS6yjf0M/t7Fn5jsCbCki1iyK4zrl9r0GpWD8c1GDCCLKtYIiZo/5Ew74Nj5pKqJSkZeDQyWzS23
+G/Itwnu0wQBTQW5LNJkyAPtoG86H+f883Gi9iW4thKT3d7FnMe7XkRC7Q7Ye5K33VLxnfeLffnP
srZ4XKxQiP5jnllYJrLC8eQ0tRArGDm5QWsO+tFBc3qwEy0z0S/pcGseaSCnM+fqPc5d5ZhkcyMx
MIqt0WNHW/+O+tXL2xJPR3Zm0HjvpoGjX1lPVzLfBz1uXMOoGU6FYCqH8lcQwni7UC6N8fufceAx
hx+n+CYcVxPMyPZM1MATmYd7wXVh15x77RxoYjrd0L1okDaFvt3AO05y7Uh9HGm1sS88CDN9KXbQ
pxtF8KSBHFrp2frzrZIwGlodTnp2rzvIAQNsUAJwpxEjRXsseThAK2LjmP7TBq82U5mCspXj9lc0
vfaiv1W8hObzKeYgFZHOyI7XNkzZrLe7K+eZvQv7i8/DHKPK0oIOSIGDZ3CfzLMZeNW2H2i7+caE
MB2A5LnL41Sdnhy7KB0IzmghXKbtx7XToq3NnarhDBh/x+krapVbeumpIGa9AEs/GCpfF9zRqXDk
I+4q25vlmiyBXCmvvNdAMnomBkCQdJ63JljqtB4oRdEQCVAfxkdbbXhriLWZnA7G1gAx4hsm7E5s
L3PpBsnJktPb+R+0GekZXBHgvblpD/EwNVYPqEp/zcszLBqryj49ncf0CD04TEVi+UZO3ByE3BWT
283DGicgMbFaA4YXKwdLCYz3NM9fgnRJ3sD1YVLd27o4BgJ4jaRlGpj1rXbdrhTBC1UZtr3twpST
vMHPcRa5PcX2i3REmLOgLSPUt9xANMWaq2m4/aDmS5tfavR3g8GIOtX8ys4FUthtWv0orWDCvXN0
4nRrno1dAFIkOjkRYJlyWpFmE5VNBp+D+mc0QFrKyIzRPP5dTpFClUeCHVx2MaAEd9dfuhfyTyZV
B7boSILKz9mnkNmdHTBgN9gF7/525FVjWIlPf4nloKM2Y6thYyAVKh0e6aMqrT1yAjLvRJIpP6dT
rBPy8FG/OKwOwSf4Il+0cF6h5oDSiQh0WTs5zX2X7nm+BvhDPEMAXR8eapBqLasD+0BE8l7BOArP
xtIVzUxuUNCY+XxLlaRHutecIHx0xoOKtT7cGKmlyVEYHSl238VX1dooP627WmBvJB3oBPtkQkPB
ySEZORWWPHJeWBn+F8DmgT6rKP7IZ4XhE2bHM3ak5+9PJWE+o4ZElYWMVF5sHWtd3c9cTaqdWEC8
P7wiPvyCz+Lfngi68suVUuzzJcYHaoQDV8oAighkCi8/6E8ZZFV+q0yuUKfViXNEwRfeyMyh/AbA
zp9PrkCzVfNFnrzjKyMZ6r4zyzrAG5LDE+C0PwKfEr+L3yBglbaLaFYUEoZprOmhy6l91inrH9tg
8U3I9vhyNYYXfuUXdY3JcVcc1RY/zOcEdBzC7XcIS6Sd33+mBjBjTWQslPSIFWvmA5fabniqhnyq
pHCp+1U2tU2lQVwOJWL+uHRJH2ReJGggjoQMOvv5QT61uEhfgHkun9r/1lx5dQJjP/rJgiNd8m77
H2LejKGlFjzlfgoApV0gIoZfAwPH8JQvm+EXNUeHb8THkQmw2r379ET0y3mkvIaGnttYVvIkmhOs
XwslodPAzHpr4u+9zk9T3tESx4BWEJLsTKjC4ozd3PO6ku6UBZRpVsQvK2+IZBNwOg2vyWx+iZ0d
5Pt4wprowGtV4gyouwVEibNYFcjf+ZGugypsjG5jlCRH59aoZ2VZSsQcekY7aRJEx7PK2vkz4FWI
r4SPMPYamDnpcGwQPtGuiUgwg/0w3y+Tp4Pf+MNwYZvRmBG8ZoBwx4PIYMQWspr6/ZGhenKdMS5y
fk6GNI1ugxnHJMDXaSxcgwYfddLxieGcoS+NkLWixGI+3aU3z4QvJZzwhW0xB2s7ODptdb/m77fp
6Id81bPzYD4GNeHQOSMGEtq5bk9HU09QUP/yRydlCNhJG7fxyze3RsAAbwb5ujsK0i7uETOZ5O+y
qw4nYjUuVeW6y1wkAbiUQPrHsAoL8beOUqDwcvyemfwwQ0ual+Bi535+u8breKzIXes4SikVMSCG
57ndAakrG9V4huWCtkVbaRwnZ5gPU6nEOXSKQM009xoWJ2u6S4zloIh1Uw+JiNeQxfCnnzKX9jZB
mpudOuS0k/TLx/WuYE6roRpdnwgVSzGASLr5qkTgma67YSAGk3TXCgYBMHHP4irnjSkNLW9F42V3
MNMW4I5GgwJHJHk62iZ62zNdTc7d7qTSMaMxcrE9vGkEdUb+hRhTY5Brb2s7PDZqScgk8PtQzWrS
QYsjMSI3yqlr9CsTPVvfzr9pHBoDcICtQg0yte79jl0shVpErgP+yn7nQ578hOmuss/e6jfLzzUd
EN886M2LGVgPVlnqWbcfbNMHpDLgQWPQ3amiAoxznvPB1OSvVfO7WnP5j+1ayrHezDqOLPbMKdN8
d61u1e+5KS880LjFf1kU3wq5p2Et+qw3D8vaGh6al1TRv4wuGwMwp7C2XRLJU1jIsxK45MtIkcdN
m5ImJOkbuCeuyEMmGCyxyUeT4CjHyHIByJonl4AEuY0o/q2+A1VNNnvfrNHPuitHuNw7WwYHSPfA
itjz2ePdRE1PJWTGPJO5gZUruzOOKlbkQQ+u2iwYz0ogTci0N5tS7SQIoxi2uVTUutBHbNOvjwTP
WpYyUE0Y9S4ln4rz0uw1jq2wVqabKDaCFvOVYXt5BC/wT0w+NAk+E57HoYSgF+NhfVjiPFXE9+0m
kLXmkJowWSaI5CAMX1OpI/9i5HLKXqkZwr+dbzDJnEKTyGjpBhBO0LDCfJSTbHMDoPxjKcGoUZu9
QJ3TsWnlVOCrn5OSdY2xyJ6EonxzfUEBXVs5LnmtJz+QKluER0+AcL7sDjVIw4BM+FKYQiNs4Aqr
kt9nSuYOWKpILlZkch4XZ7SIK4jvZdsF8+ZPkIW3RZz0OFLpuuIRhb18++epTNPZljg7T09DR+u+
QLXivDlbXuYvoD4fEvAXrBFUalIY9fDf3ljaqjyFyegEYWl/GNFy5QrSEORszfoRHwd19bu/2MxI
LWEFaS0Vf5yye0Y+i7FnOji0lAwhCE15UOZgAlv9Llxxqc2m/RYUF0U5WhChPKqmYetuHrdwQQ2K
RfgW/eLAwyuw8fkcExVEWAqv6VXYPj41cQOpYT7p3Dbi5Yxgf2lk2n9cjcMaI6hJg/oC/6Uqhjsv
4krrmrSj9Ema8jTHDKeEdKGWPAyyUJwEw7YVtf/bL4VhPeudsVj6E70EC4wQ3s1+H7txvSFSyNLG
8yCYlWdAiBQaTAZhbGlvBHFtf9x/m8QZe7GRYmQ9Qu4J+rxjm5JMcrF/caDNpjdedeHNOgJZX5Z3
qTWCbeDNHUHUhZa9XOZKs0Pf8x8fUlNYHnZ3gax+A1WEtsRA28YXdCc8Dhlaw+MsIefusGvc840k
VamaijvOOBdSxWujLoWMm/8JI/+tApQLiKftgKSxBdvRmnkO9PZTVznEMpk14eHHf0+ZMi8KsEMr
X3VEC1X3r9XD46Giy3hw8gmSRTw07qO91c4SbEeAje51vtTjd8SRhyzV7NNo8mujPbYTUPyjk+yV
zDrblXM+L5tfoEzrxf3J68jFnCqHdwCz/ZhHRPNJ2adWSIFb50hXN3KHQXVDCLKRwUFrveedH//4
lp12icEXMmlv2zJ7Nv5eaogOhxM5lLMjIM4RMEipfBD9oRKNlIZZ4wI1waq3bMGYD0je6p4pwwSS
5DqZsTGvBqtlXcvl+gNxSVphEeBn7/6rvcFYZjsF4Ki3zU5EspXYg8Puf14VqNdldNrOPE/CtWQf
BasxZSwFu/e5xTOwwZfADSJCKJjboSNAAVG81CaAGkGS3h548uvdsmo0ZOx2x7DGylcdKH55/hfc
M05zwldT8YBgvxEH4UIDM8C+LuIjTcby2BsMs4/2Khh2IcqX88tIR3ZJVNSOpEcTLY7y2eSAcHtv
5Bd288+mVkHrxivJHQz4XpgiNFXZ+XXFjxgaSxaGBhWZGAxGAAa2V4PKxxFvC0ZqltFxkIlIwRM1
p0WN4T72rKL+YhrcY+DDS5o/j1qtP2fhHxZ0GUnxIqhjbnhA5CRPVqh6Hhy/XTAYy4y9KTFmNXyR
97OCZ6s0eMWlki0TF4+clTqooHgnV2e/VOkKf5Yhd+Nd73aVMSFLOc1kAM1v3Z1rCpxKvvVanXfw
oTP0MuIyf6Lw7MyCvqpryqDdm/OR5oqspL9qP7lkwJXJX66v/ppg3jX+d9ICrrfXV2v+UXUCwcQT
lv4HU9mpIV4hdUw6yTjfTBIoTLNMpfdHUMSa5sQsPRrh1WmZEgPDzgEU55Ve3lHV2oEG8pFXA12a
G7rG+WNzg1UHZQl63vuVCRQfAgJZzIkuUNeskcTjxk/6dC/nXxmjgVrLAS93wrw79VV1rz1KEsUl
PuzBUniIfobgvdUBRWw2L94OJuzVUDO+nx0fgoZnwx3AMPTk1Kc2yci5FLB2T9Eh8IpCpbRRT0hR
SnsFyHZ17w7Vq2LBKDbeTWtZspMSfKoOD63y9NIa2m9DgMbQKmOf1DQsyaIzkB7fu6rJFHzss2/Z
1mAZFEDadUtom8mtonqKgpxJXjBGbq3fArGDKFGSejLhBCM0enx+h8YYC8qw3o40Hc7pSqFeVraG
ncIblY/L3bnxaY8/awou7yvCNfzP5kK07/qvGvcB3xWekvX9l3k4nJstsK56Re6+cr0Zuomjuj1n
wAQqXfDZMOeAiMlZD3fm026OryG247D2OoS4Cojl0LymdEmL3DPEwt2w1n4fMO0IUx0+Y+H3xqK2
tP3gc4H8SwoPJIHhRuIMmIMsw5FG1khLhVj3EwOmpaF3NRN3QDlu+wZgKPBZGEBGUrkeAK+EIkCs
Q2i/DNkfqGoySuZM9GIaweXuIz2CUKhkA+XrOnk0wFG6TV1iYWLSrqEky7Fi0XECDWW0emNZLPtB
Ju4+WytZuqTjWBL1rquS2NntIgzxCR6UDSDmfFdFu8TBN02PnVwYFSI1tTWWk7WYk4/i6NO/EPw1
7MuG2EGUwi+X4T6RD6CWzCy+lwxLV/7CvOqeL8sjNaZNoiEIm4tzAokx88ApSIuxjTMpgth/Xn3l
9LoDExaLIToyLPNkeNmWmoz8GL9UJtzqIBu60Gi+vsMd9ygrz39eXveyPpeE5lDqU5gMA1+3awH8
qrSzcfFTZvDJ5kPKguTt9DnxlC5w2C+sxeCt6mo+9MrsLnJfPfyvtYZRt5FlWCovkBM8fynisYVB
KssGEwjYSH9a3OV9f74hynpa1Q2ahA4jnQRSYn4evXt0JfnD7gWEyHbvuxxH9/CuUu3LzDyafEIN
S4gNbUEi4xFQGx3kmpPbAsR4TL+ojFLumXXnPn/fOvkBrFCFuAk0WPGzOe+dHGsIUAdwskSGATTi
3gUisto0pyqVjNJXUjqLeniEgyvxy+Do+lici1NmgjLmBqHgjSSgtm4lTAB71nu+V4zmYPrVXW+3
QVzZSkSyVctQQ7+E0i6tNRVr/Yc+uBXVmPqMUm4gVZeA9MiL0mslbKQWThbWoVoyy8eBiwBqgJxB
Zjm8bY08c0dvPnKsOQQXali2+gtLolnxMca3SfmR3mfcSCY+KX1fPRIvk55J5so8wdqWEIfHOD29
UOtNxhWSaWyi+ay6ddWZUT+mIxhRtookEOdXzBJPRdPBpeOvZUOEXquLHkTrCYJMbHScpwk9UbSE
WM3HEU6Uoedjj8VInhxJnU2w7ZBAf5NL9urMsXAF0pjvWmw9pSr++HEPmkdyjp6IiU3GkQ5NcM2w
kUuVDyH7JuiM4EKBeXAjejQtGuhB0Jew3Lmk2mKyq8P9qlHxN9VjR240C+B5AKgFqckA1EbGzHpd
hBdNJqnNnCewI+M2MFiN+mU/33a3HmpIRj7v7jRWUEjMHdd8KEMIDi1VJoD2sCDTVG+NO6k2vPzS
VeQpLW23J/07hHMhgQMc9PqQB/NPsxLrGLX++JtvAbeSa4PvH9CxCy9vOfrGUOivp/u3s0AV429G
LaodErJKdKVjxd9HcIBrEB8bgjgfMXwg6E48p5od8oK1eHLugzOLhECAJ5bMZHEoPiXpF8e7HV3p
CLjQd14DhfeS9JFBvgGk8dxxRggkiUSmB8q8EJUWAJhgB4GBkXVsEGuvpBeAWvmvkB2svHN62nvj
FJM6jJMrxvAZ3Ki0zBWyIJOrQRB0Z2AA08BcouIpbf5D1fIfbV+eDear1cTA+7IfaWf63SQQg5IY
ls3TjIQpa6sQ/3OdQU6lVYqUAEgLVhqFSOwtL4d4lZn4xO4OUgA/W9z1h5DKoANURgx+1z+/B31r
vwHmkC1OsglAFmth5IoT4KLY/mIVXDeji5MV/IheU2UlhEyTRQC4Ybt/ctGNcIDLN3u2r2dCS1Xu
LsJ7g1iKBlRQdLHNrXH9/Nq30yc/r7uhTYODzDGf5rZAtT65X4BrrZMZk2ECdOQNcAngl6uT6pdS
yalFlL/bk7pjD2PUHFPMzpFnM+mkmLnLDFKzVst2oijCxNE+n+H/ndRCaEwq0ubBBtlXDTHGsZU5
s6UbU5/Ca9lLMq0eo5BQGALKxbPwMSf6ImEcY8WmBUCsIHJ2GPS4y4WlRp17bbB7Iom2U4Pz3qwn
rR4Ho5o+qSJfAXpESTpViMYeVsMHTVPFIQPIMJ5dR6SqYzLINh1WDsuYBErRVFJABq4VLCpc8ZSo
9MoLi/DRT8yDALZTFTxcnnJ+b9Ix0O6ItMJsA/O/rqHuLJy6fue3pxe6QBhgAkkSEXsYEVrV9iVX
uO8trfRUB9mGT5HxiHmqg9kSorjQ/2oRAxaNdxx6Ut1dcGBjSH8olEdU//qYJtI5vrwAGR6e2gZn
fPy5DbaYnVMPl70iYLfWVEd8amljoJemXTP9Sgz5NC9UG/QYw8TX3FN7DxPD8a+jeC/nKvGXzfYK
K45P/78M2ILpt27w/ttezet6VexOuRAUboWAMsh8PIzuWTJlSazIQQ+0Alj43+plMHdACFswwUUS
6Q9Gc0+Y855JAasvbvD6yn2XUrKPqkyorJmpugDfMW0keXi0E7vCBIHbNSDYhVCKyCqX8dufIqil
vRlVR/NwzPH/zokGlRm0E51Ek/B5S5GvPHO0u/gGGe3tuKvj3W0DHhONvDFTAr8P2Rdzye/H8jZC
cuX3RJG9CdZH0+R2TQzPTyzj52xUTUOIsC7oCw/C9/V8ghvAruBMYyQP/itBkndDdSVTADcKf65B
fyxlZxmDxMCwpQjE5oXOk1rHmYRG7TgeUxMOg9uUW/fjJ52PTUYBJ96c13dUn68WHs/ycWC1xVaa
tABEQkGVre4Abu/RVadADYSSDhjoUQ6d3IKQc9+fhNTMXhW1L3WWM54/iGh/DaeACZuSGw6W0JD1
oDSic1e6UgmNQV0ZtKeFqDAn80RWTVNbDSAgY9YauazgsA/w6HFpAXriqSTCgGmO4WSWTuYjJ5XZ
dxEPBUtFERPHUg3su5lMd1g1iMBLSV5LCWW1/0AR00Tne+BqyrPc6CE/IijqEy4duUpre6Mx+afu
kXR04Hhn2XMY/LGEN5368MDpLYgweIsVAACOUKMzrlP0q/QpTsAuVFGUC2AdyFIhNgJp/MSjTi3Z
BsevhVOoeOxpWm0+lMWDyHDKgKKElnZ+koo50oQ9rnk7Ilk0SXXLnoMQBNMLU+uW3sc0InPvlLcG
KNV7mBL9BdXbMNcdFOYGo/las3o/MYZvk9w1ozPzw0TgAK0jgHIIUDZH/6OpQ6yB6N3tbDGjbmdC
68vhgUW51TbW+4EwDGiLkkbJ6zd5RmMIuFYMrwKky/4aoPgeLIGCO2MTyg89HpZHaRY3a4Ff33R0
1nMyYcvhsNEChtww61F7hh7XYKVCtCP3ueCwpXdqj62Ij+5MzzN4G7aM3pGUhZUgiQqfYSoMVmfW
Dn3ArzHPGGzo7au6oCh8eJXJ/A1JvmtMEc1pwnXHSJm9+/mm+88CZfwxyIAyOJAmP1d0AFOr/AL6
68qXdj2EHpJP3l2Jf+uskEmdqgknu1lFU1al6/NIlcrQneY+sNH1NgHwspl0F0VHeJ0K6N7tSwcr
Uao8ZYG6d10wtOfOyab7RyyopjGkzJZiNpD3zc4Q1tY7qNNilAx0F5rzBp7JUz0FbK5o3AuhsF7Q
qYT35M7j4Vq/Q3INnXSFZM0WLfp26aM2ltZ4u2vpe4tAGGLkEsJXNf31sYpA31n6M/AGD1elpCFD
Kt26U0RmOcCWQXmtx5l+f1ZuEA9x1c9sD0na1wnqbl/L3itBGAfZu3ldTZLBWQZm+uK7Yo+YY9zR
UwWmzxXKAT3+P44slhuymEtNyfdCQi8+dbvqTNLfzbqKXjChFuXW3ebUUp4HeZhppUh444Rso0aH
MQelvEPsl1aeuKo26kSnuT7i5Cx871XgMsv8q8e9cz5WbKT5xgHbkVXLBqoo0ZRh3ssTMkImTEcS
JMehCfFdDra6zIkAlgktnRh4pYAUpBXxGMoXu5uXI0oOjm7lBF9Nf95gxps5DCL0JQ==
`pragma protect end_protected
