// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jGnoth16plap0EJALYj6vJyPJjAXkZEwIWea0bbF6gQn7zVWaY39qOUNs68tdDTx
7a1Jt875nIO7ezPKq0VMg3AXphfeUoyQPf1MyU1ZYDEDgbNXBoRJlsqiWSDYkoYU
0dluwH3/9xI7Uj/kGgE1ME9C/G8ZN4QnhJ8DyqNTo3c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34336)
Ynr3g0WX4IIIS41yoLG7MfREcGdI0IJgHlshvPjBBWUscOdAK5UFqYeALyibhWew
iZ4LBhCr50ppMh28tLuxAznEeWI5vUrzjvrHdO4yLVNMPY3DEK7cFY6FNUlGxrzj
knKK41YXBTWLXSPru0V8qFvdmhaKynd/zq/PCR15y1Po0CvjyA+3NYw2axhjOPsJ
1LgRYPLRtnFyPna1TZRU7wj5ivDs4KJCsxegLnJ3oNTX8GGg1nAzx+UJsdn2FXBH
NvVqigm3VwEBl3++8EQAw3GvDmVGGCRYH+I890wcNfuaoZnJQUJMLgPOTMDA6e3z
qsMT1RK0+knTGXJ1DYQebe1h3DFck83QPQh6e1Zou8WZp9M6xM5cc32ExGgKGf3B
HSjyfC5cpd3mtYBZqS0Yn3V992O7WAcCszboRrAZ00fIps3uxkzMrfxKU6LBv9xJ
l5mi+dthTsO00uzyVj+1lkqBAKYs5XPIRG89JdEPjcB8NxjvtYo7kh0tre9ftDC8
K+hRbW2MFHNDShO/5d4LCNdYta2ZfbK0pD06mO5GUXmlT29Ijk52hl4JTfAYgJ4R
KYx8Ytnlq8ZJknG3og7snSobG0cdgLG6oIvW5+o4c0lMIKQrerDZzjaaQONfiU9g
NZzDzXwTk9a8418YrnscRh6yDrqVuAykoTBMciXPhm9tHsRYDyCpTsNqKjGfFmXx
n4TgCT3NF7WKYdKO6z2K/WD7yYmMmT508pZ8CUcMBPTgHeB29FuHiak245yyMxxE
rP8pU+2Zs43u+0/6zERVxR+i/oU5d74SvWUZgoKKk5vSatWjMkoyBtKjcd0jN6Nh
wkyGu6dFOjNMQq9RgZy3tmERr0vsefoo56y8APcLPBixXhHR9wF3Y/7yZiXAtxXW
0uxR4ZJ5POTlT/DYvu/6fclbaz/W0eL8dQRWvRzuBRvzpDtAkZk5kPeIl64Xo0/b
poH1CUYxpxye2H4Srxt7AClxvuB0MK6drF7WB0BC+a8ttmatMln19nBZFiZw+htV
COf3FFbayn/ZK+ktlKwA9Ag2BEOkp7ZkcfLQYC2BowUB6aCjRUhQyNSGr2UMOzRY
HuCOQ7gXb+GHLJR52sBurGjqtImwNEJUdQflVxiQl5rggfNeY9Fko8UjQMksf+In
IZLEZ6frRw6Y04c+Yfs0FDcGdrtqGgmC8Uj/hfcN2O0P5nMrJ9NBJIvU4hLf4LlI
8TzhFN89Z0PUVQfVaLZM7o8tiTZV1FWZAj0L9HFdhgpAVv0wJUoujf+AEWxNFFmM
V84zkQXMIAsc2eHkyUCm03h85DWxrfkWK/g8Xa+6Gv0DH0a5ukTSw/7/gpb19xTD
Du5UIxvesMNecG08GB5/loIQeCIHNjfBUlO9GX1BMCZ/KO0lHDS0lMX5HDnAEF+9
W19i7avd/oFHrwqgRuNTnWa3TXrgcufNxmvwL+LCuugt9h+mkh3C94qkan9rZBZW
cyzBsJWsl5fTielFdyWtjy5fiOOtPyxdut3VdqoM/w+BTrrX4X7vc2vCDM9biex2
wOAgMVvxx5n4JkaXHmHH9rLeGUB6FbCC3LlRvoOrdqWbrs5MV/EjDjNpEkDdpdMJ
NYjldfnxvKDmNmyjugDfodtUmaYo84EoX8P31HMcjpXKEIN6ZtAUGS0aTNrklqEH
hHWVD4rOKEloGFPFbGxKs5w+KwMB0buK+z3tom6B3ZAwd/ZybMlb32rOHajVn/Sq
KEODLgTavqapVwwdEJIKP71oKCdcz9YtqJhA2tbJCD0eqYc0y9hn1K7qkWsBNgaj
BLpMBlBcGums1pMq9kB9NDzxroQvOLd9AVMgI1kmRrGsqPvvxspdG8QL/HMxTQoZ
NwH3Xpsx0h+UyL7LlDqZIMFDlKbDtI+TkNjyjTggj9ouyhJLI79UZdwEZTBPqCAQ
3EFid6uHsJlPNKtL6o40m886s2jz+WCu85C9ibmcgjODpUueg14YBZpACaV1Mp13
TPYBlKgxjq8avjPHXkF907mr4VHuPOO7Rl9CDVl5NfSE3jjfS3DuMZbxwPVmgCMk
uyScRJb96AOucwwt6ivIpxUo55Y3mW0y7Elg8BdILax4Vnqsbkwj2zYMtP3x9CMC
F9t78SciCgr5wS4VuakMB31Pl+0Cs4IAQ0lXhAQlcC8hek5suvwNE0RZcIyWEqbx
yuCiBZQuSpajpyFpo0np3fNZ99YXwh55OBkA236uCXJMOQd7tL7g+KSH3+s8onIg
PM3dqoFPGTj7/lWdF1ZJaICXqeR20ZId2JKisYxfz/rxK8DaSaYR9PW2eKFcAW2x
tYKpJ0A9K1dUioVEZSakSP/YCaZ+DHo1GKKmJdGKJ59W7964BAFr1nPwzegFiXhL
WNuDHAT5hhiQokxJ4V0q30ZtCettlCXFHtBS7sf4YMrANXpGZPP/WVBo5HyGBvQ0
i2pKGVJ84VhpX2scctLHL9inwjWeNQ6so3JIxJR3fpJlydRMlyyZhbecL/kUZ0W5
M864gLOTztKL+bGVaKR624+hYyjEonSJDxK5ycocbWTnyQVSPn3fpoHO3KX7kbEs
YRhYg19Sb89DBt8lyzcT5YqKV8I48zsShro6pVey2852qTgWEgHMRvS2/07EBZNA
1ywnGh3kghK2i3qymMdWfi3mEnZc+7YS7CHSM7jgH41Oa5wDNtm4nFo5pFh4OU+M
BhftJB5sTnBoA9Fmwmu/hP1eJrOb1NvNama/5ZrY97WEm73FCtwzRlKaMkzJuFbC
mZmAMvYjgSPifejsnzVunSTINfeoFWa11ERJ+3+VmGGsZgK4UgRaWO1TsauIkEMI
BTTBQVyJdk2qBms43bmsWgRFtsK2oI2GPm7dOwUTU46nAAwhb/YMTOzh2CRpX93P
DsGJp76X1HXKiJ9wJkyvl8QL/DmB31YRoXT7tRgRAqmfTBz3ZRuFVvGhtpTg1tgm
wI2bx4plI92sYAauHUoaV3AJUtS1uuoQXNIwKtzBK+IijTdNLZPOeiwAjMyex0Hi
UU2XXani3XvZBWns/WKwRXQsLA5m0BR9Ft/ElE7Lv+yAzpALd46wfuJ2niaEY2CV
KAbXL1+2CN0mss2txhD75GugBgcdZlSZMtoylAb7KAtgkebFocABLdlZaluqWNZl
gZuCP6bxhs5YFTDFi18K5Q5sXJ5Xp1cmpWX5yhRO7ieO4LDc3galk2G9znnT3ws5
auiZYNrMa7Yb9GDSEnxnj4EkzJIdTnThI97PPGkTY/8uuyThNkbR1AWv4GsFjMNm
urSY7wMSJ5berGYPW+izxvX0iL9bcmNwRd2i47JYlOyvjGrNLgmMIiFoevO1xxwH
YDwQiW7YFRMlua1IaYmwbP2ib7P9t2ukeZBvmsVxL0++gQzQxaGQFNzFMFqGgCv2
/YygomrsXThxaqnen00bCAH11UenjuLMx2MJjmj+CMuWT8487opc/M75zXfB2MSG
CdNuJe0Inn7ZmyfTsgH+v5jvjl6EQFL8Kv3xZJihGlZmvErF5Y5jS6z5Kq7t1wbu
W/LQF6Vl5eelf1AsBYuEpyA+rGpkcaO1reb6qhGkXz3JsWZgmeB77Nfm6SEqbpWS
ETjCy7S2k9Mty9f+mpIi0sTYlmPXNrfYss1IbOIY9//rjqeWBDrfnROfK1Psvike
meTaV8STDczHbcg71aXyN4A5bx5Q1ERCN7rJFdY6NyYjtziKp1HK4GbPuoWUNi21
TvwtjwFDdQmRoeB0jvuW2kZ9PWG4vfELf6Yw3rrz33SCM86454nBVmQZZCipjJK9
aJyIDxjuv3rAT9QLwNzLxfI0Sy3HzFjLksVzv5oP45BpwuFS1F8uRqSpgmujZ0Ut
4OMdU8YmJxxfsJolKYEhsbtdl+4zuwhiglnQVTq8CvaXwai3NVK/sTSqjBppJBNc
Za7WEt0f9i7uPvGYFu7jNMireThE84dMf3EOUH1tPHs5NuqRQTZdzRqQ1gPTNxoT
MgA+SyebyBCieq+IQIXjgmYGFP1+Fqjxtv39o7rGWCyilt9ST21q4wOv7sBptoOK
GaN37Mpi1rhGoS2RzROChRm8hEo56YEY0d/l9ZcNqtm4mzXaRL8b7GIfGa+E8vwy
nR4eobcfrbf431ZLHqXTIGu5XQGWwIxmbFUaEQi6Pv0x0ynwmVNflGYCwc7HI4lM
iffhudzgDDIQ1wOqeF60fWBruB54hhcRfXFRkQSiqK5WxB6zMNik5IuxLHUDzvx4
I9xkXZHIj3VK1qpodO05MCHgwQoSAS8RZ82/MK0Etc0ISqvKVGpy8YOcfe5TE5kW
XAfI50SQ79/Yy2oqbnWcrXa3X0+1jLGHXM7ABhfdcPF4JGhOoddVG6K/6HKzfw9W
562Y0XXgoCL6KjdvyoUPtnkQT4NBqhC6sRtRg4eTp64mO65VATbbzJ3YIpT94GmG
yhD6WNpQ+MejyL5HvARUJya/iVFD6md1fyt6qlLt7di1GR2S76rSvKifWFH4RHx1
XPzlXLGA2alypmYmMn8wz1xBcv4R+/QZUV5lLQUKh2f46FsMG6osl/iHn3TiU2Ul
CZHkyNYRzwa/tQs6GSwVf9OKtVMowTXxEsRuxAUjUJAUQ/wETMTYpAyzOACFK7Y5
GyrgbxUJFZLr1s0Y3GCPJuszaHDPfoAvv3DIyGU19XpAtpTMFG0tmJhy5n7OvGqJ
uzfUuw1SEhKgpYsJN/W+heV68UBGJsW1RsiTN4sAZgeju7fvz75eKwKXJYfcYHtC
hXX6OsNmUTnzU7Dx30R7j0dYBc4vwDosYBae/gLiMXtpxlEFRQsiiDb2cHEzRppu
tU00HUeUANPOOH4y4Kqcxd2UjrEBkXce7NDhZeErt6I0U4NE2beUAohcN3Gf6EcP
UzVxAsWHU1zXc3QUV2gqFusSwi77H2JTUSW/sH9SnYoKz4Bv14JHALgxELKemqyN
b48HsA95zTHLtKcHgTQKgd98ZH61xMGtjaBV56CsJZ+EUTdo2QB25jdu4VVoFWAx
89Abl9blYVRCGNmZqANj0ud7B3mbNsXgUD/x5abtX+YknYP43ZZ9evOLoes3aDdx
4OG0rzEgyDlwdHCemYalHUHcafvpIXY8IG5uNduVRpX9opk/sSBa7qkoQQwLg8zE
3FprlJJnioKKuCUXf5tOfhgYNxeUo21E6cWMcSAeWPC2q1UKzAO9AqaBZAn2E9IA
Z18kttcSV6+FjuzzXDGGtAVsg+bcRrQSZfhNGZywKSafdhbmHGF/lEPpVbXzsznj
1XY4BsbVZWAn7gPMIitIzh1dC0XYPLONUUGWXKojPthwCFhpQrk1FVeJkPh4ps8M
9PGByON97El4jr8zM+awit2cz2yJvhNppTuaznVhZ99mGAeqFt1Nn89WL6L+HAj7
kRGZ8Mu6IOsgI5rcNl44KF8Vg2jz5UsE5KxjE7wyTWaDsOuSs0h4hSd2/+bTaa0N
fkUNfaAg6jmBHz+o66EpLoH5nRd2DbHg/PlErokGdPuPzIzBl7Rsu4ksce/UO1a7
0Y2pNRLxjY+n9AyL5hFSoRfvh23QPi56NRDgfiXjolykouKLRtWdDWRC624IsLSD
zyeJ8bptQ6qCDJmEAFzdOlXKMBA03L47+odenh/l0Ws4mO9MFEuhkd55e9drfAJg
KCTs5o6zhlrqI/+srrGfFJBZEixfnK/wDc0LtpgKhBqjt5dLoAx5wnlAeeBBKCsY
wDStLfWW1SJjCC9QFwfVNcdLGomX73tQnew5brA3MSaJV3mWi8agCUsRB9aHZ5v+
sE/AzS2s3jcGD5Ib9UoEU6fntIQymawGujCap0AcUJQ01UNCQzc2gWnETc8tCY1N
Uc5z5/FqAYZdvzq/PZZ7tLKu8I0FuEeFLtAcP7k3Iv4+IjLOR/+EdhxRdAPds36l
+5nYEoLAw0vmZY9ImNkEf0Jq4xDJMNhRJxShon8/CLrfQB9EddWjHhKWCO8k2F4z
Ep07mAaJE4rvR+VXqqH4ndx/Iqmlb/iiZsyF+yw3hLmlKZwkq4mT396GUIficdJg
rXpqC29DZl9gg0t1cBIe8IgaZuqzlYfONjlTKs1UH1ClhgFS1otohuc/sV4PvEVT
G6AIzjDQSIctfOoXdBo5pl4s33mijxMazkLxxIhdelcCjpj5ItvQxWVJIrNRi+0v
ieZC55fffA9zyo2vXak93U/gXUYK0MZOzwpMYxC42+TPLsfXieN3xEMo8F6SzDTb
vlKBmMZ0dUceNLcVTWTzVNHr67EJ9i0Im7/7jzT1yJdl0MWdPD669pJaZUSb2CI7
E1d13yDcHK5SStOl46RNgq1nAqse1T+6u1yBZCxsYQ+ApMUs87UI0xKNUIcxdPGE
LnjRzouBlfYK4h22FcGVGHXMJvid/FWrzmflZnXNUlRvnusb8Q3/WYp1+DvaIdsx
ONibwPKyhy9Bbi5Xomie8JLgtX7JguAi01W1J2qMBgg7Ua5p6/IifZpHdfVKBfK4
n226jR2bO6idOY9LMRA5imM1AaKXFUh9k7F9+tYUyWfGvKNm5PKk41y8EyuRrjtl
YVBKExx6nWW7z2qr1++6TIJrTYSgQVChch6Ibv/+FbMxFesXnU0B6ace/lAaVpiK
K4VIIZyipz8z0UkVqG/GMm2m2h27BeHZJfF/EP9VsI9Hj56KwDF4xmYYQXhcxokq
GJm1zED1IQYja3I0MXJr6z6HR7+FSEoN3BDvTCDlzsdFU0JJpDYBytCye3mXyUon
YKJjcnrj37p9TPqWbe3FHq4VhmkMt4YG0D5H3XgfSUOQZnN3NPfpdnRATFokEbEl
V6O699+3CUjL5ctBMG0chA0jN5HlFjdNXJkqrmeWIafGzUbsb5rPdSkdl0HJRFL4
iQ514vLuUUF4rpxWRvJL/xLMlsJDwZ5y6DFAT+GJk0aeBLAwI2siFMAg+iu4JKal
YBr00i+v/yICP7vdEAHuUS0ShkvBxjlmwCCz4jiyGbW/1jq/ckrwIo0uSv3KNiEn
Wju+jQzm1M/s4PxHYX3zYxPGopnEccRmp0+ExLXPH9nHNL+AllrcWFtRT0gQz4iG
CvmhIpm/QuExrL9ooX1bEywac+KdcY7W/Yk1NWC5gk1WV9c2X7x21QqZAk0fjNJd
as2bQvId+Y2RO8FcTnkurRSEuQ131tyHVuEj1WRp08J3C/ZX1UmNKFXGpjbPt5kE
JprNPtJXROtHT0oE5VIxx7xXSal6UvkIPqo+ntY1gSBt8UB3DNUTPy5nYW0qQH6z
OGLCT7g3yaY2r7yvDpBYtWqHSHt0rVBTGgUlCEyUjRLWl3hx1nNqwf5rP1j0YoXl
p5NMhP92TA8FQ87AJg+c+BDTc2lyUlF+3VElBMS+y6/79woulGTJMks4VvWtrEnb
ygcrXBOA72Ail3uQSKwk75euVw0t7h9LdtQjsaNKXAumabrKO/hpvsszrMz1pJlP
OrhsWga4vvP/weDwjBwWG7jHivr20f4CPEjqDfs6q0l4t/jBSPQPYMMfkDLYsdy/
54892QWNbwnMXESgykfzezGEFAByWKnJwDsXiCNveJCDfhEtPWLn16jqJJZv52jK
tkAC2y899rpLNtxQfLkrwtE4Fdg5xGDsAaIPHy0LsYMTzr8TyXYGJDJxU5ODb1vy
hBNFy9X48bvEwkEt+I9Z4LrCqRo37LNlu4DkgsUfLsR4r3PHtrCr6y9Ugp+c7ZCZ
wdbW6SiB7Sxp/YVeUqZlPPgCkdaAYPtEsc3sV8vNPDHQ2EU63qFw5sLY44H2H4ux
fs2dfML1ASCtQwBkTHX9reC/lIzmsrFabPDJeX/0AdKQSOMkufmOVkol/ITSPo+q
HDAITtM4btKk9ggRQfNxxAinY7oTqANKHOPnK1YqNezipxasUcwSDTPWkjKdZ3Tf
1oS2jsSJdSzlu/VaYiX1afFgxZ8VTHklCiJ5UMlAbOooAPjHNOQeiwHNjvBMil58
moxzZVLRc7xO3YYgVeoVtaQca0OoVvsSqJIUC/9AhXvsc2bLKdFKNTzTw8+1fYFL
HAv4WMZsgOSpuRNwQctdvGqYgWhtTNr02xGIYI6oP0IAux+GrO45RyvwT7KL2TLV
2Tjxb+bFMYXE8qEEfzw3UqebCfaz7zdm8T1lbuYZWxYS5VQGTe/S1fvkHnC50z9S
W8e1uHNjuLO/O/5h2o93anZlTyeSHzDgLytiIluS1EYps9pgJBsr7UY0ZfxQnXny
m0sAMbZYdBjke1V5M/GWzLMzPns8Q4inYhRM7l16mBfhm1Di5gM7VCXUD1jkfXzc
nOx2ObGmXoFdtsguIPh2lY8DLMqwABy9UDbKNsLt38WbG4/0B8ftloDm810JDIc0
/T4XgvqKRj6dh0Oo5id7wI62oC0Eeshsp007M3XYr/B1YM32RX9wE5VZWkomlA95
3keMVUEbWEhg/Xj+dc4spwlaW+vePzujj3XmOt/qF+FMWpGPI5xPfTarilxThdUD
Tuf6ZEX/HK5nAKgtHeOxmupMceAp6U5ZNc7K3i6XEClLnMp/jaakB5yMd6YUrPlx
7PPQ9C62lqR1gLyntjmp9ukqqoV4KXxqKlrVxQu3s5l04Gi+OwSnpfpTHsztDzI6
P5Vwn8w0kYvUtJMd1DjaDRPICR+MtpB5RFlOx7PtgjA9M76Evu9AJlrMz8vVruut
FjDParLUSxavVt5TZk7bIyPHLfG/Celr4YMZvN9fliwSl6Fey06b61KcuIfGUGHK
ab0jRjPQFx582uBuOCHzUiqJUImGuJcXRi21S/QM9Jid6RKVxLtfuLyDXASIM0jv
80qNyrmIQrLbQOit1u3FjVZFj3Yhrj2mEoGQneVgPDsSa1IFEVCbPXfBVNSab5+W
luoSS2Itmaxy9LbqFyAX3oLuB9cUwZkyzkVugW9m9OMgj5jjSYcXQgkqR4gYgv+e
+R8HWFhFT53ydPatHDpoRdhmSgl+VdEMQld/OhHfVWwKW+RkVCvkG0J73/1ERYp1
QKPq/rlZg3uErlQjGXnEAwMtxbuKdrv8BXZCdMxr/JxkaIh3W7yiMylSx8Tdth2Q
zOhd68tAR10LnLU0Kk46fMBmkG9qkd2ZyjZY55Q9JSD1tZGuXbbli189bt98FF2y
1zAr0Mgq85J2Q4LSTcqckXQDLFQtwL7pIZSi0n7GAmacrISE5mp84DcIt27re7X1
c0Tfgly46C40b6CpmRT31f56HgpiVCdqlhYJlhVjPey8ByA2XvOQEPT4pqEKnFOD
hvc8FCg5LtaUipWr2DmuMXhLLguUsbG35k7OLn0ZwRvWrfLCNHX+2tRG618tG0h9
5uBT3tPEC90YojTaQoL3FjHGX1Yrl9hUH8rR6QyLlTlfmbsmoTOVEKh4sNid1OCT
K7PQdZLEHAambxu1Y8vGaiEzIHxoVCuIO4kY1+8Kq/J9gGtAsqEn/a7TgbbVcwfI
CzSeeMWReBhwwyFxrBx3s/5325Dru1MMNHvRRyylLGWAyDgTt+0wlBuD5DQivDjs
Pr7LV3ANWaZxThQjDTvDetADIWD0s39wzj7CfmsyejNwyZtKH5PENRHrJzfF7HAJ
Cq6BOHxGYNq0rB5pFSHEen5lflam+wvvZ5SRaaR+cGe6O1mZ/CDQtGYnVlqI0xb2
Mf4/FFuz/kVym8zqfCbux0YjDPzfHZrIy3fiMmWNDp3z6KQooLUNjR3jiyYsYGtW
M6DHLS82Uy3C2YOpFRZ1Pe/Ww94JkS7MmtedXQvSfdSpKOsxDOubTIYhh0Zk/rsC
+co8sg1kg7zjkxC1h5g1ykBSCou5wrhr3vHGMh3UFF/DfCEqqqHINAjetCmLcbHm
RrIZaLlMVf8Iocoz+xUsINfLtEZ2L1i4fGK+3BmN7lddKh6OtCWCNxHZK3KKjA+w
zRWPR6AwHo2Z8GNJRD4DrfcwiyUCk5BJdQ39yetXK5DBtBc4kEPOIrHEv/ee32MQ
3BeOBME8bHWdlLuCcWIjvbf96hwb4uyo55z5eMRTqzfLRfqtlrK6WIN/fKJfzTsY
cd732TU24nBnFPGfKHoZVzI3pKFZOGfdKxdLcJbl1y16hgBVXJjTv9HIyv5PNoqJ
zg6/amhMOcdOJHGy0k1XMQlTQ8RnTVD06cUCJABHVsPXyAL1rP9jVeppEZ2wk+Dh
JwaAhxuUavR1hT6VH9Dpx08RXSw4BGAldBiLqWiQb6BpiNiEaxPxq3g7xr/DZoPQ
fqy659bTrqnYvZQVtyu8LyE5redRKZhPZaqLZ4H67TxnEqg9MDQJ+GNZ3Fc2EyP6
BIq6pnWKmjbx+JQPuCcsm07kMWXH89BZARPlqO8wZ/DCv1Zd6I4XpGeiREiIww0M
bl8u6l9PxugMNmdfqc/k0dor1GYi32WPWO3yNQqH0Hy15/23a6aXnXJu1vzMLAPO
SB6lOM76+M4IQ/WPCMXJ192hbdxDSxvlYsWjdX6yNL0diBpTDgggQBvvnpohB8Y6
2eoTLUsPFpNxTgYLe75a6GFoAV7HQ4sPVO/auoR5v3sX+TSrUdSIlxSReT75M/3P
2fJmqiUNyDPbOOXTzBj2GG74IN2iSzriNyT+H+vTrfQz0u9+MFppbs+KIFTEmDBn
p96ON62X/fjoyc/ea5jJ76PbH0ER9TzE/k+VV7MX/DVmWIkhd7udddG8HB6WNEdM
nuw3l4DCh0z9EiT6Sh/BLEhB3IzdJeyeVU5xaNab2y4ay69fXmhBAFSa7WerpvAY
eJilrHcd8jioVYg6DGL1FURfee/tjhiSKiKL9QOQ8O/60NslpsXJjFLG3tZ3JBRc
e4he4rntngIAtl8PACk2pVODyHVOMzNSrR8nE/SRYtGfgTdapQM6ytJGm2JLApr0
dppQTccDlfgjFvJTDw64q2XP7BLr+xdvdkny/Oy76j/fqlxtcLJNJo3B+KT0gMrG
rBA84mgqP0TVBfAi4vfbh/LOHKMlwrLCSgj8jc2UWUTUfYf7/JX4OorGF01cqnmd
I2sxVqK3yVCPdjozO0d590dObtscqMjmGB9hELa0GUSq9P96zgQrjojh9QMGqaje
RtVvBofQtXJeJMAZI6NUnAWeNY5RDi1yt5SZGPb49ZwPcY/Dy1QstvWDO1dr3UjD
dn+/uGo0SqysQ4N6h9pZTWqZzsA6OwQBx6faqUiUcjCCBmiu16bDx+By5N52/YVw
mFfulEM08fxXjkgyI42WcsoPhyBZcTSa3pWwTntC7vkVwYXXiZJ58CXdH9nVyIDl
O4PQrg7Eg+C3L2Un5c6g1LF6kdBj9SZJjT0rjga3rqfqbqWN4LQW09UXSO79avKy
5iWYyZvKiuf1weKizeM4QchwKrT8O48aJeLWlXsD7VxxubWNbKWppxyj0+swIhvu
E48RZNCgjuksZqtGAsM2RS8pGl0Po2cMbvxd+FNb7woEau3uw2Hy3Dd23y+CZogj
ZLHIzBDnvQZ+rMcA7nU4BDOfpEuE1T+YnBZDik6ENGKIr85CBlU3o8wl/Hc/N09V
SEVwIF368Pql6TazVOGOTco9Bx+8ecKYpFupFScUvb192dA1b6fAr2DsZtIx+Ycd
LyK1245PFjMXPzbhc3qrwlutAvtiRmEfAoyCFdm+w9SCJN6hqymOxJvYiFsxV7av
Q5Wn1dMXzFTiR9x9GGvz/T5jO6b+kBHbolCFc9KidOnGFhn1E9znxRNWsC/xYmuc
YOxF5SmQNfw9TU1hht9qhFbx07vF82qrWWMOoEZ55bnkOWltaJoltkzykNdzCEJN
C8n5fKrkt/wCcO8E8oIBsNQ44AVgo68WDEDKLzxMEPUPhVlOD3sCsbOpuIpzQkba
UCJgvbXweFpXaRILVx9zZqJg49nnLhR+FcWsp0I7YRzo/YWMQP6XsojpFA5nRq1T
+QokZo/5h2pXepFpf2nOG3Or6Nr5HJ6MhfTeMzdfPD+DL5gvhZrJg7QAh9fFtRDo
rlNyxe4LCEz42UeKvL1ItavbkA20wIfAFuTutgU0x7xRCtHB2hrb5pOBD8rqaJOP
r0lkSLVSV+RCmXFHHrDDhZaTac+GA6/wxuixFHNa/jMaPJfbpDsnpLX51x+GTbI3
sOM5fooI1j9QFUAXRV0PG7JmqPu/moRm5+gpVgJHVqpudJGLegC+/hYwoXI9NrOL
9qz/4aCMk+jwbyEBeyHZl8r77sklMyeJP0C/JxTfHp6BW2NUeCLrEbU7t5sbk0SF
ZTFBsdGLXLYWDIavU26MVGV8n/2DWdmkf/RPBb4MxrCHS7Y+Z8qJy5vBjvjuunh+
iu7zjjP33nNu6XFPnJ0kGyPvtkrB3CMjs2A1H3tL8VAklglczfr9NRW7CuK86Fx0
/gRbDrpHZGwTgcaljNjrG9MskjoDpw7TsoCeV6B1WpEckROeaizXtKNjxGBmGpkR
9KXHSg0MLeRoQGZeyA2YXu+7AYLznNIHceZfq3LxvUkYrj2Fi5tomzI+rOLuJxHb
9x3VVz9Kkang9UOR2c46bDTJJcxrL2I42tuu0iaXjzwJ8XWGd5xR9luo1nfW7RiS
AmcqSzBaoZZOmK0oTCe6bDRo2mFaLOQmQK/gVPUpH1kiVp/v5ll1xufyEuQAl3te
JalapHuDRwSeGIsrdRwIzn4BKfLOy16DXvzWGo+wI621tTM2FE3kfXSpR9tGu3T5
hHXMYpHsX2cqiEUZpdLXqh1RDNgBmMwfpfEOMRFtHV6qkAH6hhdrjc4kxx8ifURK
tF1bBmSe/NF9wKINtVsqGWnTh7Le9OUkGhHsatEnjK/2SxkukAOUW5u26CXID8jr
6Zcynxh0+PwgHwUoldaNK7NTXgYSQRuFmlr71xBr83Jo/GTp7RvuwR+rVzE5roAn
cpq8wMdCfiRlnWPznU07WE+AzC2u69BiA+pO5NzbQr0Nl/CylUN7oi2gpOAFwocT
IQzvyHDDgd6adiskr8eBiQzED7lwCQsSxUppTgCdoSjNr6zicqkwEsu5tDuaMFjN
B5d0vTdUjck2cOuqzLV1pgqqEk+KA8P7yvnPfAvDBi7WD75gOfl8HLMpbhaXJMEj
WKte5UGxEoCOamqhX2pGQ7n9gP2VO7xJ1uYIapZiMvpA7bHUXaNjsxMhK4tNArNT
r3xJUSZt8R04NmKdO2fpqkl0HS51Pj4mez0LxAvzbMgxhrSk+TzMiHnC+uymZ5eO
PWYtFsT9YKyNYzG2EfgaXl5GAk5cIr6U1FxeR98DbPNwis2NEUP2NsMTQP7bXyha
dGrPgWAodrBQabKf1bEUcyUO2DrbYtuVkF/6cUWVr0S77mx8MijGn6o/QIb9YiI5
X1gtGOj/oy0wDqoniTm2oT7tkDQhEea1o5eXLVSB6dSje0UFkKW13UL0YmfZn1xc
kHhuKcrXXUHDLXPMFaYS3tXan1TSb9FWPCxMxObvJQTldNDAqWzfDGkNRBwuvYmo
XQq3tlWue+YdYoex8cREzxQK/l8NYLhgayF3v1Ekgv4WzDFUH0yfRkA6f62UiSRl
jz1mYoS5grra8lyOat7kot3kl/7KJyLRlJvmzv9xkcA/+hIfxonwJGlJ3rInTRdp
qizSFxcPc4hbES/FLuEDDM/61p20pfkxnE4RhbHPSyOZbATHeLqVpA0ZaUKwnVbB
RA47EsZAxhXNET/UNLQAwBI8wSbOr1BRoIT9WFGStjk/ZlFBbsGRDWU5jVB0llgY
7ZpflHhyH8WlZv38rDcFczmDVRXW6WH5IKaopDRiAo8lu2I2XeAdQYrIYqD3fC/X
20+FfPSJ4oZBzDBLTw0aY6a5DoryjF8h+e3dJRWmOF1eU0Vb8E/hEk4N0gZQQc0a
lyiFNBMKeRLwvKY14D4bgRRsfvHesl92atajXYwl2iEG6PXwmGz77EMhq+/TSdEd
dwNfvtbQbrTS8LR8P4bE7Ildl9SZ3w3Rzqxwmavlp55T2LUHQgkBcZER2YdsgtSp
eHuugD3V+ZV6xO+zaygToBSxJriN5EEuJ4QaTM/L/fWun7yJaJsds7A8MiGk0Zln
/T6Iem8JGyzOg5O+uhe6hbI2OdvrjWgNuSgOHqWrCVgy/vskoeaSixdA6l16SRkw
4awWZaE9ldQ8STgs14bTscXcS22ulKHsKGPD/bf/SCxnDeXDv99NSs05RuB/aSYi
wqGB8PLKskaJKmYaDZ0lRfoYCqV/rvCxXWePD2ZkTWKn1TvpoyvOAYYepzw7kSXH
P+wMOL34u+lSk/jJWkL3bXTY/FS37B1pziwrnx0/kaUNDMD3Yb/wmlmDcCvusU9x
f4Ds7sERROBCkRe3NuwLazJu7VkTjLtzZEmIzJTN0QRIiwWbYfAmtywKfiIyEuYr
oy2XojoHbzQUhp2nGMJh663t4/BruuK82zvHIJx1vpU3fL9sLnkjOxmBbJqzEtZ4
jR7CgXCqntFoTEOWiW5yGDJGWhF8OETkYgm31fLehIPphRTph8RSffPnUGhiI7/H
KqYh/kLWsjv0QGWG5vcQPWG3hFDUbW3r6hI2w68376y/dxXbY9zB/eSU+eBByQ40
urinQZfuYfzTMNjrhevpVV04+HoMBmrXPEdjHEpGdgbS/ub97rBo2QHx1CxrOuGi
rWzpDLGHStWF2KU2t9+jBB2rVy6P4kpD2GnFaHmYScPvK2bUg7kngKcaD87WU9e6
qMtr1QKy8f/c6W3DLU6VkblsyNb0llboXbJGr+rbbmdMPgz1mMW/vSdqjL2KgaDI
6f/1FmalKNCeEs6PVtk4LGTFyoPzTqU5+To6IzNGGME8R70tqgJwtQDcZFHnt4fW
KDXQL4AbYHqgKzSLdOoj0SLN4Hfzun82MaINKeVdQlMxqffATYULRU8WhOTh/tVv
iuescO5XrJlPvPn3uKfPaAxd1sHb0PfFTraWS0xsJOuZLD32ol991Cs6YeNbE/YX
Jrcl2t5R9HetE5Qh7rFVrwN6mS2lTwDtpRgxAb+mTASajmEhPf0KrtIcOO2C1SOE
6IG79YShbw6tvJXWfuGed0hLNEoeSTwAeci+AFj/64mIN+OaEr/0kQ6wlKQ0KGtx
0eu23OcttR9abAVdA3PtKBfl2PBUDshMEjnia+7cxLJ7l2KYwH9faQNCdfn/toWw
xQEYKqunBaKjHV2Ttc4wTgx+7DuMIPSiorzhA+y4tkuG0FihUJLMVqPpLmR1bjXo
zmIGcf3PxkA+yGHE6iCOgKcPZBVzwtGREjiefB0qWBv+46OjaoIscKKWGqmD+O88
WTvcp/If6zGMPbcy1BPEMfnwlsNKpsRiSq5XHp0eRZL6+hpnCkrf2JBpTlL+3y9m
mkFcVw7z+4yKsoE2TvU2IDHICdExpMDuXvyBB/PcmFwM1BN0jrvR4bef1dvdIaxG
BJ81TCmIX5CV13ZOVa1E9fAcppkVPZlibyEms5SCOcbgsrllRFHP0hFiJ5/uAgDY
Q3JiXs13OjdajVOTD1mOI0hrfpzfcpjFvPpo2HAIzp1guDf0CpQgVpZi7ScYE0+a
uO1dt2m9o/luJuJH0t9Ex4Zlg18SOAkeel1nANvx4nqHvfNRx/5qctmE4RUca9CA
VyUfC3QmvRP82YTnq3QV5mN5+Ld64cWjMkUpXYyVLEDrLx99nzESdFp/nryx4p4+
akBtq8sVSbdldvD7yGTJIzMe6OUhHJGSl31BYGytdT0K1ziw1+saGgixqtCXPGtd
55tTbennUYYQaJLpDiVwWlU0ZN6NBBlhKh05dPs4zkTKbFFtZsytww1BUQ3n6ZzO
9VawFe69uAGJ9fwDZUkbvljm8hp8iWB/+yloOz12kVfcRMvDc4MznMjo00Zk+oi5
ZVtVybBNp8SnmV8AJO/qJF6xQei0DJLqMj4zv/4K3uEbuKZHgz7OkenMDp+BA6Lb
eGXQqztWxYSgdUDKhyj6fzYNcSVFOFlGPom71/Uxo7hOnDWky6Lbx1eLwxeXhu3I
GZSZa/txiWO25vD4pfQGj67pbBjhXI1+Tpt8xiBZqcXYz0r9YB7gd38N/rCjsnem
kuX/+v0569GKf7AW7n8XwSdCjuY+cXvMHXlEzCsuuXLxjRPGwx9FGXSXFSw6zZ9S
WdWJxKvPQAO7tHaEjkKpNsUeZDfkGMZQFz94q6jG3s64Z766jZKzX/BwpDQ4/xF4
c5SCTytflZERyd6vGz6zEouI0rmdus74yzRL+mzMmqESTJCKMePOB5BUGzwrTp7E
yEb/crDBQqA4sXKrrbnNB0muDoNx7N0VqrEPHkomPP4dvuUtzUVWI0Qn8EZzaQqv
0D9sxC+Kxs/ZDYtWA8Texu8CtP2x59usujDgupTd+EVEwblNhmsd0aJ9R/aMSVzJ
0pXea1e1Al9jfrHD8LsxLsT5OExMVHcVOQruFOO7I1e7bsELUP8jyC/J+w5Wqpcp
Sd69avjR7C0ypw8X/mGWZ+ZAS9nwA/oIDW3+FmyxIUpGDckuIMediLRrgY5V8W3G
QEBTuK26N9myEE/vWfnU27z9J2d4rsg0JhTxvtdLhxZarATpIQv43VXDNq2sHUEy
zNyGSbsEd9g0mzJyZUV2SmyyvLLLLBVhWC1Cn3QZMCZGTZMZYT0z1FBZxPutG0eg
jqC25OLTEZIjAlrR6NEQTcqJFQraa6pGFILIzUMzA0tP2sjPgtUEGI0qIte/l8Qn
WlU6fPAMXTgrk0Ej6OxRU7NozLvI5cnri9kf3wE6k511sfmZHTma6WWtkk6yiuXQ
D6VDGbO1KHq/eBdrqf1w9d7DGhi/IgMZv3hRdUQ93JL6FVcr+uV6PqlDH/O8EbN8
1MunggEqu0+IABNSgCQqL9KhArKo1R7427WUPJZVcufmvcDmvinmezdRCYKfT+vj
2AqjGPuKdAjghijbS45qopvjjS326l4DfltbAIj6k4/x+zEBwmN7muRiBHdjkaZW
JG5Y5yKPCqqGUHf/coKravtsUkUhb32xGLmkjgKIBkHht6PqtpCOSYpZBb1C1Qn3
6f97elonH47/LQRB3D5/4FFXZJn4Gp/mFLyLUvW1w/cx2+x+TMkkS6VAI7FpDvoO
Q61NM92zLB2M+4BLM97z9j1numiYKvR/BX4kn12YO9ArRCT14OifWRidvKp7Rkft
xpj0SEHaLxuEA5PaQSHn4yoKnljaaRYhgNiGpg12E+wY7j3p4R2MHe5wpY5OhZvz
aut77BxJ2rfPvub1tyOEK1E5ZCGnoWyGj6lwlKMN1mIhWvQJi2nBunIlPhj7y2+E
jL6XBbXvHPyHuZa5e9oCznaOSIwRbdl1P3B7KDfFZ11kFnhcd6uX3ARr8woDfKFX
LFI2KI8NFpqK42Hjy5Y4tsk50FYPpVPWcE1ZxPwkiBenhxe9sE4p3UZSehCcIIX5
2kG7xM4EILwx3nsNsc9tnBqUaPafUAKCKhwYI19IDHqeiHhBCdlSq/SzUvudu8dk
H773AggUAZ/JW/ocviPGgRjoTi7BOU6JyP7p27i7htcYgGZJwjNd1KPxtVccvIkT
kprYavQEAc8Dkyy0Pz8LmuyY5AaRp9Hf/6YUcZJ+NZ4iBatgi7/V7GzYg4jgS9mQ
Ri0X+MeFcokwpkgTZlzZrc5cc5B94wRTXEwGyBu5HoN2szBHZKLpYyEsD8JMEyKG
HpuXfxuC2JBDGgka/GnlZJOlg1Y4Iue0myZPPdiIdSBI+ah1rD1cVGKyWlZ8+1Jf
KnxkwIJm9yKOdH2Nla9VgCrJ/JDQVQMHOVtyGrqe5FCd/iZDjxsqzFYHpB5x+rXL
04MeZ6JM7gIocqrQ/XMe7kVMWJvZOkoCP8DDTsKsNu2fNChUAlEBAqnIgqnwWwsl
cWhB4UYmlO6fBP+i+pR7uOG9SKPbTaMT8jBKHm73JJCBttvojA1uvKgHE1mVKr8y
hBxMx+dG4+hN5IXsByF5aGkjtmJbFfwT2m+NGX+rsAyTFoA6hirkaBHJduG7SitE
Rc1Ri84h3KaRBuF/z71FWolwTm0AxGFC3reTYknGRXEFULmUhWt7eSETDKGNi1Aw
If7o0l4893wQHemrnhjP0ms25YEIPRVIBgoDm2W5L3UBkVayYlzyvs+IeuBI58S3
KMXaRlM75rp3zfiPDcMe62nwlbGKiHqJCXBf2Kt1GfFqKmFaTAV8pVwaupajpVgH
OYJUZonzrqi8gw+9RLtxUbErS0teJwl/ziJEGvYFDB3L/a7GV+WXjJ2OqTIaJlAN
U/clrp+Xtoaygm8CDn7U+SlPfjMfit+35ShGDhYyTxZdJSi0NHDWbL52UzpZdsUD
CLkjjRY5Kh9WK4SUHeQTZYRmMgHalpeU/qHWaLi8b3xWGFv61VutzGUdCBjZD9U6
QSHhjV/kYu1jUgwGXjq9i+nKKqzYVPDW7Bf8Ps6IVURg1BPSHXkNxEEGSzrBpCHR
jIsDTm75ozxYhOdNCYvIuPt5EuKMF38A/j9BZvmCR4QutXODH/5nBKo5E7G+ww9t
knybg/o6fceYQJnSUzf6j5islYpbMAl/OJWMgSI+3v8varAa2U27TOS7H9k82S7c
dptQaWpv2cfO9plLd7nPG3s3ZITs3lXbHrOHBG1wmOdVz0cDUG/u7seKN0EAlyeM
NfnxN8Ktc/EfhBlr7qc1NpqHREcWF+EDjuWbN+7llEWq1a2dS7m978rwzSAduSmD
nggGuJyGQh0e7De0Pz+VRtdmDkpgRGNKDQU+01cBmdBzAHuMwOe7m7pfCirLvEwo
rjSm1SN44P6NZ4Z6A8Y+zE8fR5vlCfZUXQvn3/D+zS8zEZpKRQsVn9r578d9mmON
XCtQIYtfjHRx6x1EI5eShv3tNWZN3b4pF8+nDO7wQAALrNv+Nm0dXBedVKhB0ZFg
1kIsXE9MJzDIGaO7oUfHA4DjZ7SHiSEFkQ6qxYHetsGFZRLACTp6wGkuFLRBmWFg
bGqTQvmPzlf5bOojVqa3pbJEtzUnVG5PsqND9EvS2ZA/Fw4GmU+arc/c7bENNv0u
bfR+qI3uOpRZIDu9+rQ8kV0nBsqj94S5BGcEcb+vprBP997HHTJdUfVs7ELC3qU2
+X1oMhnPKbHdarlsp/x6Gyfss2gz9i2SDM6vngOor6f8YqoUc/sr3HtFsCq+BSAd
nNIoRvtuFqDFw50F/3MuLHy+tCEWS0r/20tFhSw0neYqbMzoUgAnqOPIsWpzE5nw
yBYq2z+nlMjh0z+7AnLO2FK9OONBGMTyr2Y1WODLU4VJUL/bGWIlvkL50gqdxpdd
CuNS7aDVjtVZ/MwpcC1eShMhRCO9SsdJ23DYVbjP/QUTT8VF71pH2EIZNi1o061z
VI2UrH5nARzCloYCU3yElb4Kp3JEBvTh3Yw6N2PXbvvJos84d9tgLsvzxvezC859
DINrYFsnfmDhavd0KGzYakxg84MPjv4Z3PS3F0P5H/Wv73MqugUKBGsIMAwaYL/L
OlqqLYYIhJ6UMArNPnfpDHGsXDx/0NgA+R/k6BtKHVVAI5FEv98gC3zJg2RtYzTr
nRraoeVInEYs+ZfUiiwy+wimL8tDlVzyN88dNfE1yPiU8PsmzuXd4IeTtzFBVTKj
wUlTwdEbI6t/4AlQ4xS2tpdgcQ98lnm37HIm+y4xgueEQbCrsUWALn6AmPfeJHhn
fxUlVGCiMsqmT3OV9uGkGfwoTVnxzlxWH7cn7FiQ07F2WJUe2G7II6/10rSYDt7J
IRzvj4S+5FYlKidtcO6vJ/WhxxUABp1/+QPwre9kDrOj7NAw/0JgXJhCL6El5fvQ
7RJShXd3IACr4SYMGq21cvPOzBOhg5lLc9vXjxgZoykXCqC/AtiOxlCGIbeCij9f
ASZqSNtvw4/r0Xaby0g5U1lvXkAWMLiYCrNNKie01//3NoFO+Hqa/nrUOOk+Kath
AfmllByXpNKA2Zk2MgXHFZoX9TgzQxrB0eMmZO43W5/SkmUUmKilZ/n3e1InpfYu
b0UJB8ucy9zdkg6G1K6LVEHgU4RKJOR2UV43FJ9XD77cOd3yQQyufAtA4UW1Vt99
Zmp5oH2zf9JMRK23jrr8zhnHleEv8TjnMXSoawvyl6zFAEtshen5odH1qrrP9Y6C
tSqCuz9KZGhQdBsSW0CrD2dS+0Qqvn/JXSfejbZJOmHfU7Adj5TT+OrY3+kolNy3
iYPvQlM2A79Ge3QQhBjZGWskfglLSF+Z9zlSCy2FOPvkgXDiNQvHLnrZiK9vdhK0
WH3HFcFg8w/Uufjp6SuyOmCEDAB1AEqgeQhmqqaRcPJ8ZDDyixa2AE69VnijR1D/
6464g0QSqaMKE9lyGsvEuNqcf2ggMH0oLL2YgNi+PFjQ/2n36A6MQfAI2s6VV/XR
z52LxFN309BPKUaeYNrSbcFx5oleXKy2dwJFlsQjFlx3rYmk9PskEOpWo2gMeJVj
y8TIM+zwpeVjI6dlBgufd2u60aXAfwa1O913pdqPNZsTvkAVqNkXQMCu4g+R52Wy
O/yBJ9sVJf9WY5enXdVgEu5pSXqjw1LV4v1oIi7ifHYFzbCKjRAJFKeGKCK0qrnh
9znX1+2lq8Y6yh0W250qMGARSs1WkbQyGIbTdG3cqn6tsoN2vyLymfvrzYKST/Th
0REH9pqLxasOkJHKoF022/AggvAGxMtR/Kjsf1W7zXIzYdOpo//kPGDOMCmjIVKP
mBZoWxNga2YCt49Nn9z/fY4YM4Yxjp51GFs80jM6/sE8sYg5pbyn6GvVrFwrtQLt
OMp0KIqyl07C+kOfOrguz2HN4utE7nuI+4JGW824jvmSaRJNjIhPk5r3zEg8OY3+
LDxeaW7it8Opgg2AZPC+csWaYPeTJQjCAfvhlSA6O4jGpnuQlQ6dgr3IpLnEmgbl
blla0lCY1f+yjnrPRoMlL1H1Nnd3STlE/1rUtPPWNDG6oDnM5PhQgOD3JMdUP32D
/eYjaIFGbFyKqHi/GbaEAXE7KDEWDmybM5w9giFdSPJRHf39hbTrr9v/7c25+oPb
iSU81bWq2gpxy/RG8XsQDSbn6fNzOcO7ycEULABnZx1WnslkUneomqk3Z7f6WO8o
E4BIddP7Do80ofxrxRXR5tQWaskdjoDunYJsXQTSmOEyzg/pHC0SihGILDHapHji
OZr1exc2y4pwVcrUWknketB+rZXicgrjSIzPURXRbzz1ppVRiHHsms6IB9RbSBN2
2DYMJONxHG/AO1cNtH570sG3ytWRlatiZSqsSFUcoM4UiFfTIH9+EIHAZYvfob37
F1h8LdystbZvkJssdXQeagQpXW1n47nzO2PqN8EIhrzC9Bg50UF/XO+PJt1WO4c2
bpByBWRfNC00pz113gqJgMBYIaPpAwAMW6GXiCRDAELI9/8HtCAuhhIM8dNv7e1K
Lg27ej2BIiua8Zd6uUvSS1Mz2h7x+k6gDjSaOOLobz+bpgQPyJtqPeLQIBrkOPoE
fCRhv5fMcgE7g4BqlLatOl86BW9NfjUJcg+29ptAQX7BREtF6d0e2AkKvDkZEHg7
/AjzGHoDWzyCbx3T6cs/s+GZrHM56xMW4O18/zUeExcvIIVITd+jcVjB4zB6cp4P
bCdsfd8N6vpoifrxiECYetcZ8g6II4XWITku0wuLYDdbmhpBMsB0CkhGtFBeeEzu
Jd2r2rf9pTh6OxrxA+/9xB/R7PKLSXtIJKyRWfaFgYPqm12NIhydboSPT9ZvDNH7
c0+wFquFFYC3ZqT4soeebeLKoxNC9b9PaVSeqZA38IhSRUuxlr+ocY1bolE1oN0s
Z7rzVANIsDPT3g0XICXxqtCHM/k+G/k9qjBYqpnQOWWm+4K8YRrpYuT5EWyW/uf2
k8s2E5u5LZP+oDfEwraclg55yYJ4K2+U+q/l6rKLnTKS1NICa9sdaUUzt3VVw1Gp
0tspnJSg3XQ/c8GLvSRVEqq5owmXWGzmeYYIRgr1fc7PgE0N0+TKIwMPhj0T3bwz
qJhj7b2ZVmSMuLtF8gOeCOElBuR7pi/HnnSqiGTlnjekmC7umT3C7CMyBzZfkEpq
psN5GrnsdC+4IOWkdjTP+N+8Pl+5PfArrV15zEfKlX1cHS1aVOJuoor/4js0j3qK
e0VuB+jSk/96Uh1Xiv+CiYURRK0OEw7zNiKkVTeoepFggaN3dnp5BnaXh8s+GfRd
G2suIdTkON6qj0PhX8nfm0h3h+e96ltEWV2HOqaXaxTVUWzXP4T3//p4ehn1/ucy
2eb0H/yBMfeA9VfAo+PEe3tsj5+dlioEF7dOVU4Y6jumo3V0GCs0SmF6KAWxNGdY
4013Ii2/BM4xIDn6A8QwW882Ub5i9+TNE0865p4vJSBzmV4JtFP0P1t7LDxBVbBZ
OPBJlVFCnFvkQuOqoZK7YHE2BC2VpwGQjM8MBPHoOuS8pCDGLIRaMfaTrNBERlmM
CN0NLlCXr13aCm33a9ch3HTPZzyfg/vhPru3Mpu6+dpV6RhHvPmkKQ9KDksIulbD
15dDDk+Vo2P4Qc9Z0oYm1s4/7MVEszY+lkDLRawVCqAFG6046LufcyJO86Xtno/u
b7L+mRdizm8PCNAf1Z+2j/iGhUeaDTCFhgO0JYLRBZpOEjC+aXB5l1blr9mLlSGY
RinylhCDcXvfrn8xgHnZsWS+HrxNhFaPFABXF6pIRM11Ftf8PCzeh3DxM9cdGQU0
NoNJbUYt4pNpNYNJq/P2XL1Bdc/LmwbdjwZyIiKFWSg2LrVFya2WklULitQvNl+0
ff7HbwGlJdd8wubGkz9AKaIxdsTW/WakLfColXh0orVfDiRYpWKhh50I34nXTibr
p1z8iuxCwOwwjULbOQFvRGomduz36PCz3zLnSXbM6NjGyobbxW+hCLf2rnTreawR
60OzN/ufodWyLwk7Yj3HtEoxjG4LPAtTwiGV6rEf24sA3rOiltMyegLB4/zuemSf
c64oSsohfC7gLqjFzkvC0t84lUHKnvL3Rr+PppOlG/zlsPQO51pKlcK86HDhidXL
HdO2NPY96ZozAtgdRCByhkyjx1nzpYOQaW0fvNf1D8kantEApKhSpf0vVkJHZPEu
52tnj0THDauJtGmKx0ozpUmYwG5/KatnzydyAUuFnamQ8zdMbi+nNBwm+H1Thj7z
9TPhDZYZ0S/zOzrxyA5XQQTWhtK864WxX5heIDdz94ZKb+RWIbi3388NX0rsLE8A
g249EVdWMZSUlKdCqp5aolVVoejgt7aOXWtk1fepaQCB1LFkmVPNBHBekRFAJ767
5v/K/13DBfmDCSHmBbIzLTrm6suvQgpxt79djWk555Go6APgCC0lK3BBScycc2Pn
ZaNRi4Y14Me0OxVMZugtbm1t9hWOFr3eRAwPDnWSdVXxtk5VdoiLPywA/ZgAHkf7
YDEZ+hT1svGy/RCbt6Px0OzYRQjswa+dTUf50k0KvPNsZzEpKb4W/wSbAiTZpTJp
as/XRZNn856Hon6LfrM6IQ8fK3YlQXSKG6U+SsLBli3zh316a7JGaj4GODzqW//E
ITnoMymNTGp33WGghaoERIFNiGvn7yRAx6iVfgTGJMc0NZ4qI/mpNSeOlGzdvj3w
SIBREqR0mU/jx+S37K5ddxK/svrRnPne8SShyZZyPsCy7RrSoYzkySsbF+DxzMzh
lWFlQW24CmUoixyKwNxGXCluBjzBu6tKTQJMrDA9rrMB6wDCs0n6MCa9T+/QsT2q
2xddCxAlE57HZoHHaTs5YdAeko5qLYKo7a8+nAmK/dBFtU9EdwE8AwPSSwvDT/vc
DhEwahNZYYNeHzKpgatrvic5XXCYH/YpC4oHKV2oSV+JnGQaaUNgx5JhMGllUQPH
1+zFie6Ay+POVbsifiStC7ZjpbzsXsxX/fsxI/6LQJB6wEmuLPZ3pefwKzCVYKt/
Kw1XofqvURul2BXFi2Mruj8FhYpzBmqGLIp6I5MklS0zXASs24ZbG7J50nomTnBN
DED8Y3mDDHqP4BXUSFvAuxMSra7BfR0XeJQhXGpCEBNJ++ed4wQWEppg3/FYeZsD
C8DX+YxfdLW3PvLajPwpsmSLdp/pzSaPHINsM3UGKeYiNOt2sBuYQA9EP6EB32AX
S6er58wex/n+jLZNNuQ3uwHPlQobHxuaf+MD8A+siS/9oNUakGv6Z2wA0Bu37Wnh
RhDnFH/E24+3MzYtDPi6zNata729QZ284HPNMnGaKnQyphJSPhrQGgInkC5dh1i7
8fdw1fw3SsKETxcyVRoZk0U9LR6lBL2Sc4ui6tMSNSHit/tGbjDg8n2hIAKArDsg
MY8YCzaXdlQlJqYJshvsKDBO/7i3bH/ubE6NVBe3h+1fSN4qaMKZh6JsxxM3VYfE
Uy37ldMTbRsUQtTOfb4HuvpXkaOpXNZCwMaZqDEC42mwhjRtB3F+aEqGVIrr5irD
CaZDAL0cHViEhwYgl6wemF/3rwfEEkmLS7hbI+KdOnESY06AmfWA80+1/AT04c+T
bfUjXq91tz7UCiCoU5M+nfP9s41CXrMUacB1LzMGkKRRg+4Ycx3fiwtFelGEiLNF
Wy5Gbh56euttSeLu1c3Q6nCR7i8miS4qm6LYU10etlbrqxlE+UGADpsRp+Rnj8lN
2F0G36P4itlp9rFrBvIefCaV6PgpTy+hiT3fWM9ibVILFHf8cOSCOsUeBxg9RaGK
Goq+XV/0KXpPZ5RLvjQTjuI3VAOGqWywpFlD364j9T4UXYpgQe8VU1TZLtC2zQUl
uZjz/4alQEGNUhofTV6KJLGe2ssxn8V7O43iySDzW7uVoc6ZcZYysBKmBDi69N2X
IqgWGYjvAMBd2dmhr4NS+ra9x18xqoccFOzOsyIlcqWboDCqWqggcvV8bjompcqQ
f9av2AByGUk8+3ZWwwBDljHWUYu1FEoYcQsEPBQ2lgleP4tIeMnA+QxR/mIhtsby
apl+lB5JZnf2nEH2/gIFB+Ykuy0qIjayZBVPf0xxrzjHcJBvbo6Bf3DVbM7Nle+b
Oa4uVcE+gHMkZ2ip9Ljxl+ze/7d8Y1RpxNvCtT9pO4VboLwWDc7RiKSur7lO8von
nc//D+86EUIPwM3PzKVQVWHYYj5uLHGK2mTgoMip/PC4Pr/GvdW1Fcka/6LpmaID
h49568oMNcvyXdlilvXU5SgyWgeOdii19sBr20TtracPZOWl98YRRFXvGZplIWfb
0hpkZgJAg+Phy0NbniZFFBvHKKna3n7RHMLNCerHj1XbGoa60BqkBc3Lkh4fRJxc
KYFBGUW7qSjNUPuxqafO4qYlx1LGOFUBRMoGqYiiYVwvzrw8sTWIe9oQ+CXP4dJZ
dyURyuqau/5qRTgB0sPwpk+KHygjU5gc73R1LPrjEj2THuYCgrfo1DF5leY0iPbh
jcGY6zTQVXeab8ejro/gyxzvYtc+PhUsoxKzIaaIbOGF3dfYmlfejU+NSJkpgImE
EBFHeHxoBwQjkAPbMU42pXk/pBW2p9beidF8F1LgLqE4azlOQWRZCYo6wcCIw83L
jBFjMR8l8w9RY8I1vVMzvk7HKknm4HTfTRHdE/QJExpLFU9XoCbJPaa767UsT2mi
XDV0yKzCHnUy3gpYoqoxB6s6XqMwkggoVEg5fbwEj2+L+k6hfAivq6N3Yybh4bn0
X7eDhrMcK4XqCHNFKVm+59FSAvhB7LBGbqN6F/jMf1X2HsIMdfxaQKNsRtuP/1oK
KVtXLJQTlcAuAKAdrNVPDFM+zEzUvrIK+0qmWJd0qCAzuGINtdwz8WJhu8GjaFD4
EySwja8VypppQO/OF6Db92Ajn8O5rLfKzvfG0jiBp7tzMzkbdvyA357V3ZSrU+AS
6J82NtEqii1clVkUF3I8Yxz7XcSaRR5+ecFmB8QdTIGcn0+Eh+Q6mfKJCa9wu9zx
xOSIEfas4hGwR2MEV4xM1CzWyJ9xFTbjWk9ZvAHrKULkao+3VJ9DKfXH1aCPkmZN
ucf95lKIMA9q4vqw7JPjJ6l0RkGyssDbVMrMBAqM0fQ3xoDzxSn+CamSt43R+83W
Fjn0PnWvigl2hCp7s0kM4FRADGmoUzaRD0g11LgRz7lqQ7v6XLLFx/pFHiPgW9om
1+h1xbVQXHFgBmh2ErdYIDceBZMJin2nYLf0odfaE21+FHzhH0whs6KUyh7K5RpF
/22lATS0EQaXP5xEBjhip3N8l1dmvTFt6UFBU3S04ab+rUCiQsCrDkd1uqNZ4o1Q
79jzZoIsgw+FvzdBKaGZin1UksS+4eTM75DCzt8ttnluMhKAWdjlPBevlWfIriQE
TR8WTGHJ1l5qta7+9fl2G1sFzC22jB46F604SKPMMwkfoSvv7Om6Q6hj084qjM8q
SM12kAhtlpiIzKuwm8aFbP/zR2eCrqxn2cdAEGeG27vUDb/Pqy2GM7rbCkUEOJxv
56c5yZ/2aLwBlu2FJZKxH5Lyo60BW+acEd7ltOzE4u+F5XH0k+VFp3tli08aqHfr
OeySRMtKt5Q+dc2DgKUFYFgnQvu9YYC5eoSIwgDXO+cLrm/J0C5EjLA8mUzWQkFN
ZMngYZcWX4jF5e/ywUQOFpYRHDqQRQmBH+RgsJYBAZbHlh/1maMDssfF7aIthQc9
6OO7kxGSdXKSSYVZQXFEfdCX2BFsaKmh4J79BmWXEJKWKRRakHM3uFB3tWqj9gwh
2fQ6fs/OWTtOSii/AbfyN67tcjkhK4ly04tP5QT1irh07r0CwuVVJzsTf1tCQhCd
o9eY+zYlzAAGf/oLkJUnlXJZZLytK7CCPALeb56C6NfnQdb3tUD3Eing5f/Vcv+T
OdlFXKygedFIO5KE3tgmucLmfEfa91H94dm24hPB50sHiiX/fNhTwIT13K17dNRy
D5b5ooH/XpHNGe5bwVAhkfJpf/u7I3zRJ5+HZwWVlO7VP3b7KVYBVYuDgH54XWb8
L4bd4unqe6XnO1Do1jwFtjQy1xMQRqWwfBZf0SESW0kpiTnHUfnXfnXa5doO8afc
/WiS0fWy34toesS2o7RvpfSRAljuEvozU0Rj02p382t3bnb3C3bFgyeaZsgH4oHb
9yzl8uEn11OLmYvEqMPPy610hm1yHSaw0Ck8Ahka35B2lxosxFy7jroycM1QgdcT
fRhewDfX03Mn7d9dzvV0rSnwNnuAPC3xyXWP72j9OdtTnkFFxSjDJlJjmiyyBuh1
Ur+EOcNjO4IDlZkYoFv4vdeuhXZwgwtAkM25WsA4dQf6KEx116dZhJRufldwgAxT
79G3KmrK9lcVdriSNFr2drX3iF8QPB51ermwyVNOnUCQeeJEIhz0emSiop173mDO
fZWDwOMP2dHUyfDOiU9Wdqe3NY7cDjIWES6yi7ZyI3BYBpBKlTTrQYf3iDZXI3OC
2cEY33Hp1am8mDUirp8O/51T/5PAU1iqEL8edWGgRc3TDkX0Zo63djEBHHS9eCB4
vBtNPRmWL/zq2/5rxIldTg0WKCb8k4OwocR3ic/FF7nJoJMdLOnFm9jLInpOL+m7
Mt/vMhb8ORfrI4aFRUPYLIjf4SEKiFT8uP1FeS8+/9/Ccpe97fYy3U3HSzYoThjY
3QPjU8x2gif31SLJFt++9bXkZucfgy0T7PaB21Bhn9LJ8Nka1z9tQUnIb7YJ3ORV
8b0gsNLWtcEseLaEFiGka3CepdXjmALzbabYmQfFohygN1Z3W9PN60+TpMFB6yqC
oq71VKX80GE5hpIg178YXYgObtfiR8jZQColZIBt+hi2e2VwEzaOrCSYGCKDbE95
5zQr1bJb+Lph3uXuUhF04Y//vc7juRIfyd3ohLa2tWwacp9eVDqkJyaHyGIoe5tG
C5NDZSyu0Odt8ajBq6HP4jMqR3gt6nOCOrbqxnfgNXQbXPR5hPt+m85AnjWiZus9
C+tCH14dBsOjESWzkVOtapwZ9Bzk+mP8qcL+oncCcBfuQtiHLuQmsDJqM17O1Dz+
vJHmrX22m5jOZ8KdKbAr1PcfT0exYRRC10aUlpOzFFQjp+YotiSnApGkx+nC8R63
RMowv6NJAhs2c5+nkhAbyb9HPItOBPC2PvyTdxKBOdv4CViD7iwX6w+hjom8gaWS
XA8l1Og5//8A8Aa4kfIQPRdbfW3BgKWaaUdcUTyw6Bjd7zMU0FJ8tDQ7Ke6fhCvi
asWwiwA1VOwXU3DY6P1JX8pz+puY4rgVM/bZYfpYNMEc8NKO/nSFvEYNSXTYQPfG
sSrBZfbGHJtnUd2bS9O6vneuW0VeQot0K8X+2C8gvyPZbEj650rsuj4ieY57s52S
bgDV5xpaDXBgxKHbxcTd4JPeJA/1G4nZzM3MPbpGeaRPp9YH+s+FdDxR68UFrDB4
OqaZSUEwLlmCPwJWvkNNxYfoxWl15ROTbZMYHEp0eiOd4e2ciJOs9IoHuwfNn6pn
8wzw7LtdHHyb51kwmxWQSFyk7FGk65OtDv1K4H+0aJvuWGsWj5l5lsdNRd3uvORN
J+zZRZWG/Tl70eoDiM18qvWFRxVQ1TQLA5Z7MtVANMn4lRgHpPyKVyfSdF9U4Wdy
DOp1OHikVCrCn3j5sH3ijpQ8ajyNSP9uKWzqxKpZyNJZbQxBLzcG4VX+9PniWh0k
RS9M4YrJHz5oFwq+eeybOTOOI7v2GSw0Yibq0yFrOBE7yZ6fsG0bsyv+iv0FKeH0
XlGQB3rvMoH8VR3n1OfbRk/HmQQDUGf+bQLiBPe5wuiFDGlFXPxWMtzKD7eeZX2b
Vo5PNPeT4/llc8hcj7kJzSRGyTNESI6npySq49liW4UZaQ3hODKVu6uUnF61gWJk
gmjEKsvS4e38YhpYsQZ/IVy+YVO6n/LNn+mRo6+D3LafQ2C79+TsyGX3uSoIlnaP
fNiYNvm+BTU7tr2gfxsSslBt/9hTtlcynfccpr8t17oRr02UPVtsT3l6Hot5rTKv
IPwEqwyCnNOQ7C2P6cfzecD9XMO3Dh2/MLAOe05mrq8fRofxh7AGoz2S5qIqYRne
hPGBrklc5U+YgBDeafAUob1BOE81of44KlovOv22KSdhPxYmZQTNZNGKd0U/563H
D6rO3s3I3Hzd77mo2yk6+HUe9hBNjgZ2AFXhrDsPeh8O0+WX4Z2GKz+ifBc2tCKF
cbstVpftODp2XMXU2PxGpXosd8Uoj1p9tkw7qaMsv4VFDTgIylpQmcSAdTv4AcAN
9cWMpNuv9996JFkBcHfXA3ca3q3xZsOpzBOmjGGNxIp6/n0Bv8WgFUbFylPjmn7k
cYfiryGqpE/uJ88RUnLEqHj7AYGjNTP22i443ExYg6DYKVl49rdswiFKobUqrhyx
gv1yYzJYat+ut2by1a81kPpaBUqHmuRDmyjnKNXWFuwHj+DIJU6RHVU9idxx2Il3
n06IZmpG4HZdBMaYPK8f8UU3dRayek8TVzm+wXojTfS4cHDTZ62wh9SgVLA31G9D
LWyVO2O3PWA0lnkoBn3Et4PA3RmbVr3Mogo+HcpNbQtBAT+t8nqFd5FCTw344EAu
MD4e/2+OnWUGrIJWatl3cA1VSbYTEemIG5vm7R5jgpXtqJEY5foSsz1d+ZcnUH8U
AfIUO6qnVs+k2p3PafHMyCkzjLpEnaANnr8JcgQoFcAaS6FkUeVdsVlTfiWlcCsH
pMQDoQ6ehQ63wq8LGrRJrGTpqDZjzi/ayxCcOnN89gnHVEoowulfsnO8xfx9Lgfd
qcxMcjV2aBs4jTP100a5NZ6IafyyweToL6ub9mxX2NEBaeLNzVA9gyMpXn5KUb/m
BkxKdO/yvdUJK+bb/yIvA40Gq6GZP6rk4kEFEhPwc9kIVaP2cSp3IKEaOyQzzoQ/
6o8K8w4U5+U057VIXcciPI0aIaZuSA6xm88vETdPsyBRUTMnrff8CCHTFOdnbl6R
9OFKlD9jwcyAU144paOkoXAkyN1DuSSBJXs4YWTkLAlU/8ex58nvU0e9Okoq4QVJ
B4yCz50lfUHFV11z+9IXtmFkey8C8qVByzs5Y0qhaYMreDWxM79nB0kcz3OVDJA0
8ebbBo48/3+kigFbreLJUzDZCjAyDyFbVLOtx7NRRjcBIp0M+g1pW5xzIZvydTqg
NjbCi3ox8zGEgXRjBB7JCZlpzcBrqCTxF+RT/uLC3McRe00YF0NYJUFefrq8gzBC
p13rNpKvamf9u5YgLGVIX85JDPdsYx8J9/8lFeVHDLxRJNYsV+SX0bwkz9oZyJps
WEAStwb8VmgC0zRE1tHAQUOzfVxWCWnL4UDCoetfM/TxuHbWdLXVIrbBbZxrz4yQ
IHIj5nXW30opQwGv1qLvvUFAJIWjZasR2xw+Sf68X4gRquSiXSeXh2aIBjDYEjdQ
Dz2wWUyfD5SoXHUKLj+uVG+3HsX1z04AGbMVkhYObrXFHJ0+IIb/MQ3LKNhtwgCk
y5UmQmyFmSSPcMuyiQop27lGw4YbdrWslxEYt1HWMivVwX1iKcenemk62RiqOWea
ZWoGYVpb6wEeSLnyyNYS+LFuRH3YRcluj8xmcu1RxGZXMyy85T1bz05GZMiYDaaJ
Co/14+Igcg53YDY4kTM8X31qAtFWYUMItmzzH5CIP0boPYGMaQ0iDHSZLanWYo4a
MNkzaBYKQaCRFwRBl/PC64LSlhu8qZykqdIY0mJichh609TMhwIUAXhQTVF5FMMs
3xW6Nem6S+pFOhgJATvLS97wXQk96DRxrqXuL7dT0m+LrmN/nGgyRwUH94Swtv+o
fVDVYOT5uxC5W10nu4MJ45uKFc3hHBp3IwgQKCs88kiOEHnBckPmbWW+m4TidWOg
cZVmlNEr03PmwO2mua7VaVdtDTUROTmk2taGNK+h4CDzDHUxqpezImKxN6br82oF
i4uY3ZknYW400tK7qku9bWjBaJ/VsgilftuLFGRsIiIsCCjQvbnjAmWEXDtH0aZk
uHsN2jWiUxZFcDEDlrbzf5VbKmc36JeWYuWyt5/ZPCFajDnf+Km9DgceM/WTgi1f
ne4rhNirYE7za3Yk6WeHdQG0+8LWms/SZVkt9Kj7GGkAlRYH8d3iincz0Bb4A6lo
KFO9VJA4Ubldino3kVucfiZJew2+AoFi49ttUwWgk+pM8oOUUmHbOhuwg4T1ZDmW
r+dMehKi1IwO3pxYMTmm9qE9gnZlZKGKTrvPHCSUCIRF7owpuJvMpRTX5a8S10bg
7Ym5zeyXY9uJtMMOL5ZqKKbzwR3M3IQs6ZIpUgLiF0r/RWXOZfHSfhhhZSpi+RJU
yFCNuZl8YFSjrzI+kQvz4hiZQp/UNzUQP38li86ZsS4Uqo8Ti55yufuooA8BKMKE
0gN8QVjk8/lEa9Lmjk/IlsRLTo4Scr+QKEGjdkPRE4ZsSjz48tzmcLLicDi26WED
BBLsPcR6PVdY8roXX3QAgjYlydeprADS8bnIVyZ5PM/FAaR+HLuv5ksK+qQCqq1e
+MrpXD20FtJfRRPauKuUMaUn7dB+p9AMSf2BDzixcK1a0S0pVX9ZsUNoiiKt18xD
JaSe8V3K7LTgnNKE9hOavkyK9q64WP/4gnE7Cpr5McMBjcO561O5kUcU+pV7HQqu
oabrrhc4xN3rAHfrZXjGhQr+CPVMKIFicq2h95T6AUCHHonzaGT/eX5kCf2ha2ps
6VACHmn9h5X5sZFD+NDJp7p3hfEVA/FYa0pV6clSgkiaBPXczxZPs5+rNItr0Tbz
2qKTH3hmqmWMVGaktbcJL8pCCu6qprdTHZNnFFr2W8AYIgoP/2GO2cs9upkM0qnk
x407R/v4msV+/4qLFqkn7WTSfqhxius9cabc1YXtOvkq4/k/t+o4Fn9uSDB8g9Ti
rReNc1zO9rtZf4FhitIUjkZdwvJp/punC5w3/WVqzhhDOhPClsYj7hKCQoUPJ010
vd9BM0SvMF2k3XKzIxwnB+HPIWJ8q0j4BMe7jHxBTu37+k4ysyoNuP00iiGS7JmW
AVqGXwwwfyi+tjy9Hm0B6fZVvVTsJwIwbKR5oq4Pxq1obN7kKcpIEGiWmM/AESPA
GmOl5xU7GdGd9/t4E2gCNlfu7LO9bWWnCT+HhtP9YOwb0AoLFMO754dO5HaK8ckB
/tQISBdDc49qi9bsfPqtV1i5RwNpwflhg2KIswjClEVgaC9sKshGvedLahfDUXY9
nzgb+Zh6Yw3fGk3rpzm6JQ0xHZ8bEu3yV4g3ubLZAZ9iROdzvTMCDhTS2LapKZ4d
cgYmPPyZXEYgV2s/T4OkbUiSS9xr8aQ4F50mv5BaFKCaKTc5NoKvFBWeVFocNahw
KP30y9h0uozoNdC5I93pXA84qwc+CYR0Pp2COsSgZtHkoJFlWPmGO/91StEOBQAX
KL19vYKkDlGDZKFJBe39R/4mlJ/Pdm8fbYmqa4ao/Zhh7SNldh08K/CfMQW+cKJr
ZQqGBDgHzZPJt3f4Ny6AycBcvJgmLLDeTeiHG+SC667f9/62lwRV3Czez2TVLmmt
eKKDQESiY3RbVpJ4tXwjClWsT7nY1rk0rDsv1zcSNxjiS+mOwPbZUCVZSo8GDfiQ
PPRW00WVsuI085iT8se/3TFrnQL02G3G0Gh2WglMGY0dn2x1ULBbR+yfZpdrNMCe
S0PQ7ADpKzR0GW3Qb49AxpvKDWNSxC4mh1Ds0twxwJ/jqSMwwPMLyA3j/o15TiWQ
ZzbFunquZm5ruiNcTwCcrq+FOpeYn25O/8xYWdrCvShVUx27iGgxlR3mK4HGJjXE
6+J8L0pYjQYSpUuBgBtBljSU1oC/Y3xiGaIHh2aA1j6+Zrq+Q2ofDzolfHgLP71/
YbMIoAoeb/TZKzVkh385sPqTvgNeaTiOyN4BNLkScNF9d3WdUxWmPQVuWVFBTs0S
W5gbcrTR0VUkJtLS8WhnnMedr3vQoc9OXAwGSolmY3+aSQRVwxakremQ8CjChA4w
k1+k7R8bhXXiDh3ip9QOyDmWSro2Dfkwl+y7VunRXAvhMiEKrizgAZGt12HYF+bg
wrGlJb+W+v5jJvuKd7ENxHd8mYp2no2+oGYWQh1pEXUYrVVx0MfGTAikmMx71dmP
VoN+hSFuIQPEcvQxd0CTfkHWsW65x3luQ+dldH2HTw/0WgnTrpQwZXu+2WwN5bsu
3l8INJcbHX9XkEtvDxNPGqvpZVPNdFHWtL8UfL6Xrh3wPECyH646zYY/DcamhRLa
fsXeITbncltaQZHNYxDetX6h8pEt8wTwH2Urly2RAQDFmPkkK4NT9vH4u/Q0UoY2
ZfgsiOzsFHNQlsEboVlhSzvBbxRDVgY/8oPnVROas0DpVr41pFTxBpylZymtV1tD
Fn6JFBryMIETK8hcrp1tdO/mZq0yFPqDKJbD07esp2lQyb6VztWFYCUfbxUXKSW6
Q13u7Ni3FfmK9uJL0YmSmQCsji/i7mrLdV9jgtbKjHRvxeVgUqCBn1ecCo+ZwEcs
1HcD4YzZoNpBPwAwl80d8fpp1xbc2OQfDQRH1TB4/DUTAMabBTZsESlEJVuuyD6m
qtqT1jHU4l/E5U2HgRKQCQ8nH3c7rCFVIflA3MBqkmNtDTGtttjM8TK59cCJ4XoA
62g7SjKz/mQZUNXQ5SijTZCypVDch4VPL6tlEVDDOVTUu60BtPhCtAfqG5wR8Rzy
xP2Ipd7On7YzVTos8OUHx3HgQAhHXDFHrCTh/kc4qdvJzhdCKRYd1pX/zaintCBP
305rINVTnhzPz1MUribe9hyEB7hUPDWgzG8kGEju/e2qbUr6xqStRrAZyddcnDrP
3ux5/gubLKPes4l9QK+T+r4rv0phiqR6XBXSOQPRpzQRrUl2Or6oa1nR+RNCoEk6
l7Z/I6LN8hr4yi1FYKMwqpdBxYQroFIhiDmSZ1PZ1nrgn40IoYUdGB/b/RP0uGZ2
6XKOCtA+lVTEmRFuH8geofIrkZ7inMZOMKJHJV1VhaxLeoC0y8FnCtWGexWJJ1fb
r6C3ouP8lvwHpL3paIlWL0lfWuX64Ea3idHWw/VgGFiLRJtcv9Gf4tXdLIT01FSf
I0ZlBjxzHqiZ4pTn2g6pqWeJXRwnweUaByOIWrqVICviwIUx8Zf+BXhs3MjYawyr
onaS0GOOq3tvxo2pzHBpiwA+WUFFIgFrwMV/CCAZZa8oBG8Ivzsm1X/NVNLlq1fV
FZu/On5Jj/50eohyLMYo4vaMm1YrhkEoDogAusggO8MAIUssZI9vn2SHafqxW/TI
xuq0mr70Qc9R/ROacAQAmewUKnlwKHQY+8zMP/dEyq/Fu+bCv+asU8coH6OO8s+2
DFdcmCPBkv9mj8EJqOqPqLMAsRO4IEFyIC3PslewEanY4syqRKhx+n2xtdIcqmd2
3QcwMvEAAaNLA78jZmoZxbUfOCoNsdRin2n8CwykkpCaERhCBrDFP0pRFXLO8lQh
JSXCT5xL901ZA2iIjWJMCWb501ft9SOyahG6C03lZPObFFaLrGUKb4AEX9t/SWdS
roBWY1KehfoYVVaOJkQWj0oqh9sO5xDAtIqJ46UulXy5+RD0cuVuvMfVx3Gr7MIo
a47OF6dMMbrUacBWXhaASc83ilvISixipZBxDQOvNeL2IB/vkbFCsGWAi8kf6qqS
xvJ1dcWRIaupmLLVj99KI4iPPfV6gws/Wzo41PTbVeqPmXfvIY8dMnB1qzQkqqgC
kDcpcHR3ClfqV4HOqQQVLbs5MvmtiILXw931QkfwubHRpmMWMMy1PhVeaMMBhz1o
746uf6k4hsXrFXEWjOMiw36W8RVtxLgIwBcLj5j5Ibi5N30A3pWPo7PYkQwvCIh9
kEbGDht0Vebc1j79CB1lIaDA3gwKZkKcC2c5tLrpMNcRT+UNRYN+Y7sQ7Td1ePUd
Un4QUmD9pj9jOC1mDxG8l3zjnlMVEqhDiOOnZT1FPJsPrOh+8I9dUsTv6lIUKw1z
4yOvzjOrekGQFcYaZj28bysw1BtemkaRmj1gzdg/VfysCZpFgHdQ0UwzgLlUmXkf
4VyJdJs/fzcF4RNg0HSQqMR0wvKYBvryTYmvAeN9AS5HL6h1Nh9+4gjFTTaQTejr
dZEXsjc31wPfsZGaD0RZOm6F/77AeTvc8BjtOoJHYfi9I6Ar3FmEfZm5f9KFAHqN
GhpA7hTy72oZTH7y+4OrLZh9BCBXTXqyBiKfQqwfLrLzOc11ozvBvBhDvvzNqUIA
f5ZJuYTfXLOgEPI1BiTt8MApnU+wM2kfljFwjdceg72Uc3wTfkVI99Bzesd4SvHK
Qq53cYiw4W8ezxSBUNs5PMyAiRcZ3VsnTBKkqSo6j8HDceJpuAQ05PoF8FMvAxzn
yKMMWxyjYm0kyamC7hG+AUnN1xB2VhH5DiUKlq0tN5lbZC72g0E73CN1YWGnJVpw
sZDfR7NaKcZwPWzDxguwW9A22GFEMwI+jbeRGXfqVRdN/TV3fOi91XyKTJOpe190
u86jrmm4S6AMhmXrZRBPkE9wpfI9LjM7RYogRc+QXaiyWscS6V7UO/N/yLrh2Pvr
f2SHj9Tf4F3RuoX1GNDMrrtMD7hXnvy8HfsJ1K7vGZxlChYNFz/qzGJUwusl8t3k
SoKnMQasdsXO9BAJdIh9N9QriA4/kXid9CR7TKxHi/G4bXtE+KMWsPp5+Tr/uiUG
69f+jB5MuS2kON0QjQ7BynDAdxepqWXrKDHllGujz0Sqp8EAFIpS5GuOY9R/sfJC
EKfT9Ruh+9zOKO+WBmFcQAdT097D4PJ5/W+bf6Ngm8gclr7BmBjIaWb5XzyDIDxN
kczocdDq8IMOU6dEceJjSpBsb30mx0YOUewv6SRYk/8KFAmpgNJgKhkzXdotpSPG
2BE/ahx7RgQlsza+aW1At3wu6ISjSp+DitkmZ4mS0lslb760MMw8UMqfZuKMPIyZ
gGhbhnbxXB+ZmByirb+4X8YC+vsCUaFipo+trkNgoP92DDygFWHcZTDfR1lez1+W
EoCXpMCLb2QDCJmDxfT0w/uxd5FzDc6MHeF5xCSfM4niFq4jqK20A2FSRqqHNXIW
9wcYRMzwHLnIKeFzyHuRkjsIZBSZTMgSYEpWPkc1GitRAyL5LYq6zR/sioQZleY4
KfEpQYiw6Dhpdt12k4ZyioZ2PpVLBBQ6ggkAdOq7DpbiyMjkOnf6hZFsqXQmOO4W
dpcQomN3BLAh9bGl/5r4G2y58KKH1/MrTD7J6JcVRsK/QSvjKiqz1JCz9Quf3NrP
tpWspisRiinILOp/WlxcSw7MPMmPqSF3OFJR4xL25Bq0bXjyZGk3NAznZQywCm6A
xjJuR57Qw5+Uj+9ozOnD9BQ4YIxC13NWOPu32x+BnH6tSfYSZGKHKnNVLGDp5xHy
v5mqQaS8bzbkB/aKlAcW22O2DueLyb01yaWVIsF4d9fypY4mg6dasztO8KyPWkVz
K4Eh0GJPM4TqVFMPjlm2mRuheQ5t/6FYADt6GFESyTHM5a3GyKwYmkhS1aXvqxgy
/iLXlWTqAoSmycgwmRgywIJgEfJhHNkjo0rEg9daeZMhfOaLalnQX7Kp05v55GGu
b7McV04RzjSDwI+2EeaF1oPCGLNWn3B7hHfI2WCgijTNvjWXlZXzzkp4NN6l07cK
TDwDz+I9c8y7Xcd7BTvX6UUyFE4agfg8BfB6Q+5CazI2E3G78KoFLwBM+C6yOQDe
pKFJDidnBSytgAXMoh/kqYz3gbf6DNJH79rt9vcDOrC8QqjPLy6IgyVYV/r+HkrL
x3INCmxo+3Ouv1NnLOuDzShS4ProBOla9kUzhVqrKg2hl/sp2ArRnKKI6hGFqPsg
l4Wr4dL66zPUADdElPc/veuECUrX61lH6eVT4C8LZRt84ZnoD+jukVTnfta3DQiL
XD13PI/yIoS4+5iwA6ty7lx/lXlHATHkTkamXG1exquQlRe/19C90jPHCjYXhfkn
4JHvICSBKR5A2PPzB7QcdOUmIGq4epZMMM1vqcLyyTeW3HrKNGp4bbgkrfsRs7/S
9ZiQxMFW7nNn93LMM34YAujhTbwEn3Gez5EJidk4nUkhjnOIrjQvBKXOJECdJjPk
3GBBBr2KBDsqLh4VNhowcBuwFBQcp4SBqJ7OVVY+3rgzIUgbIRqT2UWuQFT0EjU/
ejPLzi/fUNmdnW4u50CCeF75//PEgaCN23eO3npgjqo6UBv+CpWMqITP8GUIgeyV
ek8aTGCpPfXYVpqFvZDgyHfpA5Rjz7m5+PY/S4JRS24ArZaDdjATTMNTHqIram0U
wnSvtGgAMEvTRi0qT7F0N/QHh7ZqlNNew3AQmd9fYLRByJ582rZlo5Z7fAHTUiZC
5wZwkDDEq0FDVOnnemE2Y6Lm9FuVZQsxWrtHL6dSW/CWtqyEQ1o+e7hApqQ/a6TJ
6/En0Ng1iMZ4P4r0t6cu/mVWkSKAgr88MXp5EgF+bnAJ0ejanDQd+vRODmgs8Ctl
Kz5up+fQR1ISxdEZ9Zfpzl8mF84b4nhXQVGcW2aH1hgv5M1z6KnyNHhXFNMkqpMH
opMj6XEZFTPkX/BujqCH3lpRQwU6Nl8/XPB5rrjJ5Nm87vVBSJMFvZ0ES3rLt1Rw
VcuJ07AkzJfYUk8leAIQeClWsTOYnYYb4RlYtUtGkd24ZvvjhcW0Ws0b5ipRGIVt
X0gWnVRRu5tydxgnPs/aJNZdVMTqpu9xtTzYPh3i0yEhwixTCf46wOXLFLN904RC
FgHI6SQhWDyZ6sp9LIYLefJAYjmAu+KWAdZVurjW3XfTSPJMfLqCOHr+JHoCaj6e
fmh6dY6BYOGneUkyMzetCcbx3TV1LTDGWKG8xEeu3NUvsgS7cOS9cZd3jLQ4APEg
Z60ZLVK/U2+zLMm0I55rJdBYGjppjP9kdzWwfLqkxfAH3voYsCwbXyTp1jJ15KNb
/MefbxBBdqe51PnxZVTNJzWQQIERN55l/oC3vgcwDYjy3RhPs2FteoLurOjXQmAd
jxfKScJJ2G6rHYQLabVWDeImFX15hW7aHrA+rwkGnwE59eQEzq39l4j5Y1/lAzrd
yLlRZOp5jauRsmAmQBQLN3gAUy7FHJkge1e2Oud5LsnpSe0TMxbhhcsvkqS+FDSr
5suIfJa0U56SwOGLi7puLwUpqFSsFII/6wa3YNZsqCU0R698qR8Ib4agbOwaoWSm
N/VOBLNtAmmTs6HCXZgYCo0abiR1czOJaSS4HCxX4YgleaPa5OWYhqA38MG3x0WU
o8OG1irlMufyBR+2N/j3/MkrOMDVHkRXFIz0uspqFqNHmq0mfOSxmuEXwMnjb0LQ
LvTHFqE0igxqC+VFc+62xwnsNmgE9zM1SmeGXUFqImXLLaSQRk0qDBJTxJtTI4+l
u0zMN7lT8cvFocIdm3UW8rOG2VBGsV/shhwyv/zd/uB9ysbCmmx/tM2qHFvck4L0
lxlDaeSxhypDR8go2xwZ+cFQAkPj9lsqD8oRmgIydcxoorbSAKcl89PrQJv93J+n
/A67faV+UH+od/lgBWfFnLotycW1Tw3lIY8jGZZfwdybpM6edJU/n/IuDgaAifSi
TBgg5c8acSU63xISXRWaGo/yEQCQr9GFBeirJpC3UbIjHzXvLYTnudi3GLSVPiQ9
nveCZZwmtqchf+Zr3jFy99z2ybuZXKmuQjExcXIeXmCo03lkmzwyH52JOyaoMvUX
XFLwKHRxMu3U4v7XP+7kBsYeIxN3YoAJJkn+3N0gN05N57d3hJmXzxc9f84iwLoH
fVNy2XxiVD8hTNPVtj+GfbwPgCPMZmYGjB9LTtXRxW3NHYuXVCMn5LnG09QiVsnK
IfWhdR4k3mFLFc55agi9UeYN6tLlJtbYOqVlog43NHduyhPt+LLLM8jePna0Fs+Q
l1HSjnzjT0fIPbY+aPhw2B8nPai3kDEgP6j3CP91ZexHmL7RA0aGpl8b7Zgy59+Z
3Plw5OPqW9dy+q8fKLvGFfqHndokJMF2He7T8UO82T6wm5HUP5tUsRDG56ozmhz0
vb5K78rKYctvpsdhX/K7K4pFVtcmXd/veJasjmUrbammwhJzAvp7ANuu6KHeSGe0
3GChpA5RJFXLrLxGPa1o6s5Y0pcjJ6W+hEEzRS/07EyBWx7taipSVnYQWLHyRGDZ
Jmh5DGS1Thfo8XyNxJQV4v7okUTbscVTbIHcP4hv+8qjzHStRns5j0xsFVizfJ5+
LyhWQmzii0CIIkVJNU7/5AVwAx1acVS2Y3ozI/baJ8dudHW720w3+PSswNUf0mZQ
AWr55LoWrZHwEkRkjI6Mdtq1Jlywb62jZmp/5eVQjNPjO52CwhyJRCgivKvmS0tL
QyHyfjVaJfkghfifeACxHcuPYd/i9YwYMZIsKtf86p4/6dlatBgcsbG/WRWvckW+
MlGO3FZ0TzL+lGzMYLFeVJiXvdPGNa8grkDdzQkzGpE0Naf3AuN3sybedjF9aRFE
w1tnEInX2H3AT90E4Vw1umx+hZEpwO50ajVVNTdhn7q1tfHYfOcNTBhoG8CXZZXo
Ctvf8mttfb/U3MslEEbdpwXnJJMKvw3a5+Eec/17V3urgiSlgivZMLHprou4DI5U
gG6XUunVU58HfTsWvg7vh58wZB3qcBIHkUb3aVeD5u6C96z2fxcdaCqX8LtpW3sW
XpNZUCjYy2N3E6abh7GhkyVY/5owrC6iEI2PtLaf9tUJN+NAiMYkd2EjZOXcYF+X
3InZkqdaGOguQgNekvLs4LLNiIrURTQ2pkzOCMUZtQCGPENd2l4gDIAhQJXlSwNr
8Nu/l3gZbZAhPu6vlogUyHo1banj49YocRN4MB/I+9ztf2ToV2Tn7o6dlI+9S7ml
MMwN3m+CZHu29/qigwxWkeTWL5JSpDkXSyo2XnxmGJVr54lWzaDeSbg+s5/w/kZX
MDnOS2ct114Aq2RUMEICljWLbEYOHEIcq5SUIuK1YlRpiopyUHJ/AwBexh67vvkT
pf+Glmbp5Xz/iUMs6aicGtyFussoFoxkxmhxIw+LXTaNiyZlL1E0Sh8Ut9rvkr6r
pI8SDpYjThk5QBFP43iW6oGWbWGQI1g0pb5fbIffPASmQ374IrV5x0ATNRUnewlv
179GTDNOh/y3UN0q3NbkzuC8jVAYihQz5KC4YPspw3mJ7t2iBi1+E50T/mImbCgD
aSEDWAque/5a5Rgd1hO5fD2sk0QpSVu2AV/8rr8DxFYipbM+Oq48v60k/6ZfNH47
SAH1oO4k/NuImkcnqNw0d0qSnNvM1Ds0A7ek9wVaLkOeGqM9EWOceDuynM9JZwVc
OksMFvsst3SGxHTim2T/fWDqxdHsRshBd9gKEmXhdHInKE6OEmXZBQOvZXHUmbxi
xTZYOzHKMCrgdC5kHPmRbwGojj49fhmExV9eXt1hy8Tt/bSwQVd2BSXexGQDMLAL
KAubEec7dAR4nRhiKezoVkCeauJLv0UVOgmtZ9Dn5n1vrqcbaIavVvR22E9HLvjZ
q38rzERnUyBtgOj3aCc1MAPn4m5alCas8foDU1P4fCUkCgSsVn0pHyQw5sXT0h/e
9PXZyMHBFUx+a1FOX7AEiOLnfaMfCvDn8RmvoCJV0TxqAt6QZ8ImMKpvf7yCoTI3
mIDxbI4MS9BSi7iZIWT+b4GVzJBihv0l0LAQcf80YPiXt2e/47gVlF2sSwTPKSaU
iTEMyvL4JtAAeFWKn4AnYCDfkmqcvl6jbIO+UNswUpavXz8quAyCYxCweubFtFSA
oLx9iFx30DpuO+nDXJ0zuC/5JvaRS9Y3rucF6kKEREzLNoRSxhK7KOFyVBiXqkRj
chXXoVvuAHFbfzm5PqE9oRKQrOogZZy2nI2Qt6TphM3GXmYnWpguiMUq0IbfKuKb
TIDGmNKhKA+SK28bJujUcNE0OxLITv+0+LokVgxydlgjg1qd3HtN60JayJZdnYhL
FXioZ4mVeUknB42HeVz4DTvTioccRByTqovwEw/h8614FzkU+UIMfx8bu52ukuLJ
fA/s7ErRAWKMv4Ef/6V/txOrDBqekARbqC9epwYUeHf+RpgN3I4c2VwiD/rpgR6B
yDszyjMS/wZz5/KuWTOtUYuvUuNRWQUEM+aq+kZvXeLPG3wER2Lp1091olc49MlO
ZpA45ABOTblHlEGF+/AWTPgn0elZ64nLVUanwWQDZutnO0RUgJ3N6c1j4LbDS/S6
F0WXrbcnrbdsawA8K44GqNtYfiMRk+/ymLfcjQHbuvmtDbem6uY9RVxKu8l7s96Y
YwlV1aoshqT7BUFFXOImbzKUosY1VYtKvI82BY3GIF8R917I1pvn7kPm9lrpCZyG
tHlBLUMsUXUh7lly4ZlkYGRP4+zhbVIXHvwEuVo4ss5UbU0fzOl9MjK9dxyIwudo
sAc1FS9Ob8GOopQmAruo2ZqQNBUWqiLrV9uJZyZzVE7sNaCI7qZUfDK1NkPgTvw7
rnkxEAnGKDiLMC3mR65tlbbbcycryuRKy4oaQMCJ2e40VuQyDfavKalrOg6z9LuX
NIZVb96kWS/015x9UY2+CuoUqduZ41b4Da9+lNwuIhROfbOOiJoF4FTkiyMokQIX
MBqlSpC1cQDT1zO7Gwi/M5uScIvxO1lRTf3bZ2cHqmrh9N3ty+k6a0xkRNcigP4G
43T3/OFzgStOsk0mhQWXlv7M60iwfDFISejjCNi3tpbaNk/YIUrKIPB6V07sVqAw
csJVgm+Avwmlb1JhGc2O6m65gztCbMj9BTffZImL8b5jsMAKs69pUUPnDCwepJzJ
r3kyRpDQrJ+Mw4paQMxy+yuExua6W9cHm7MgHvWg32Iw7fIuNaqpF2Dz+k1aesb6
wmj5q85ZnGB6k69CcNeN/J++fgH+UPAO7L6FMrLp9CPbBxQ9d5V3hSwKlpG0QK58
P/eTgofv5C2j8RqO7oCjIh+wbLOP63KnILUsa/U8+FfE+EoFacTamOmRWBKhXXiH
D8KgIjniN2/5jK0XRUucur2MAASo15vrVM3jxehLUMdfyW+brewTW+D6a6sdcCgC
OGtzyc+oamhAWD9sC/fSfUa0HFaHfNxMTU7jHYlMb0cDTzS2rH34aKbIw1K+KLYk
SCtVVg++vMihz6mUyRv0sahq8XzE7FWhGWFbqMORUy4PfR9eeutYooDPS6y93wIo
u+LEwFXPqrDwmihVckCYdQzREsuDYfgezbpR53qZKpg63QVoG/5J+YEyUPYSeNpW
Fpmyri9KdtR9Px8OL57v3qet8T0GapUXuj5xXLZFvc+UAZvLxhTV74AB83Mo0zip
YumK/goicj6TTP7RnJ/TCAFDoL8AWFyEFYooFzlkx2o9Uvu0NbD1Ur+7xCrDu7jR
Ibalkhc+LDl0KZIdgoYjPgazjSoFZNLt3+mK7Ug35t6Ou8xl+Gcu9TkfgPZdO3Ez
w3a7RRqLFi8EY98gVurYsuUmoJa4Cm9HpjrffF5YuQGbsqw5v2iXbij4KWpgeDl5
Cwx0Yh98TJnNKivK9KVb+Kv2czueWPkeWlnsBmoyGuRf8fOA9vmrI9DM+t86eoP/
ife0OG6jSusiEATBkpvCBnrKEzFYP60ma8b9WwGt2IwI0nNzsJ6PY8UA89M9Xv//
vPF7qihpSjzZxfT0hQmlQA53EDQl2UnVvUC8pjl/W4ACWS4xkPhzjcAnrNwY0KVL
nor87/8Nh1u7ogCj+6Ire0qqFDN0lmyQfS2t1ykJI7T9mcghgL/jxMJmXfoQN6uv
DjYsgUpMvpFkQPHhoZAp0vf2wxtTZw3Eftt40X2V18vwe51U4UgfM1cYiSjBP0Jp
gJv4A86Klk/FX8Moz96GSJeS+KW99QD98uH6/tuq4mI43Hz99eqpjvFJnvNT34IK
wiSkkgPWOk2t3aZFuCI69n0ioOyof9o9+V+HUlWhjH9ArzmylQqPXU7X2nlJ73fr
r0dZs8Hvd0IHU0hZZoFOEQQKYocnuEiDhaE5/YyErB4HZmE8B7u2Ylg4rGKUcPa2
LVSeXLbOEzmnpiqE+DPBSioN7Sa6lVSPqV5vGlV1fQCZ4a4GLwTtUpqUUw5XxS2G
7GzvTWlFD//pV6kneBqaEv5sRYe8pDIduRX47ESQ2Xo47etBROsvFt90JDf++0ka
+RPQ2O8vckhdjEdXz2NSdPxguFrPKYkM89sNgyH4O2cQ5ql0/J8eFhtu8VmF9FGJ
D9TPkferdB3xOhmMDPUBxaDEub33P2bVuxsfqafwqINjUi5jZ3/ziImWa0Jw3LNv
lz6ilsz+7ySDQK3reqiUKnoChnK88AZCcsH18Txzj7l5O6qQVIOwwogFycNaF0H6
XhPEV7tRHKKR+teIDIt3L3b8q6vq4arOcHVh6nAHZMZTNa77Vwe7aITtfhYT2Dic
YSnrCZlxHyhkkKqU4eWuAmOAXuIrkv0DfJ9yUw/Y0wMVbcV8TJQyte1kA4E6EzZv
3JZKvldt63Du1/xjPTGB5MiV6ZDu3+jC5PJll9IYVL7e1L4m+IPxTfFQRFFB53LT
P7R7JrClKX5m1FnxheWIQtffg1dhDc2sv/IZtRJKc+S7qeyOMffER8XEQtPkrZ6O
/86TONZ5Dmh1e3jDsT/pcW9flPN3pJYZaj+UBDykUn/Xwmkvb76CG7AYohOwx5HF
LQRiq1xm7SSq9Ks4dHvebhoXtJeCaefN18S1F9rhKhggFbSQSysfKOG+1mc3VGkq
QbvEu7/LjVgEhwDwrLv34BLGWADu74Ub7H5hi9u4nBGUorf7vR+1SLq3waMQ82UY
vK5vmEEECMOfl9YT1JGnY+XdyupegQtDn4U9YyFykyFe/FrgtC0+u/jYjAbSFIz+
SpmZIB9Dm3+0XSQ20PN1gdmuWmIAeXeV1KCVSKD/4Z7SEqf4IzORnZnoWRnZbyMa
hAdGQH3a9otFfV4P3S5wlZUuUxfrwtJ3LQ9RXUt03B/vV2Kj/PJ4tbUnz+MMYL67
+fOpoMPf42JrqCE2jiAZSspOYy7LOh7SW0jnDVg39AnKY5gsbaZaWpxe8PxV6sND
f6LV70n758RhHizYpgm/ATwBXIv1Aoy5g5X9ZsFVUWFiP8yEngc2OFYlzlW2dijP
vX79d0jD4zfCD55mNBCDICOL8RP96e3JVFDBg3gK6W/Oyf7ezxy+oZ8RVWbsULKH
tBlMjpqQ1bm0g08LYni13gOWD5CsBV031AVDp9tu7NvBye8rl5RxU6ue6WagJ50Y
JCGw92V6ViSitTD+oC6TcgHohxt5sQC4YuBhtgYUZdcQg/XNQWREG2DFeH2MsUy5
wuN1my4z15dlVYo/7YyRaqHN81lbyxQ5ej3D+tf1sh7kOe8mquadH+cW4WDF1+Ts
gnhJFEheppzCsiBYdsmEkPQ4gQLidazs7uzvMCgziFrnbsgn2ELNSHVLLaQjZBnY
UW6jRNSZGzHVPDT6IMUd7LAufS3H1umdkbmUgtPrfljmsCFpv3jRSxkYkGihgpQW
vZqP3vn9QgQt/e2tuNbdBlzXEvxGNbIUVrD6w+HDVfSJQRSunyGLBld33eLATjSG
WmDUhqdkL4Fxvy7QVHYz1A56NkUx8EVUnV/ursVhoK04V0K+XNE9DHhPZ9hRfV8p
JALgtVLNMO6H9MTCsdVQsJt/Y3yWwq/Pbxguay6l8m5OwTr1QhmRs0YGOiVh6l7s
ww3j6m0sUQPLRCakZxXM+nxJ5QX5zkw89o/5mSy3azKF6wSEg8X0KvO6/gyJV29a
3Q/z3w9UlmnYKBoc7nvBWCCnyySpemXXWk2EJ2YN1UT9xv72Hc6FdX2iVEF/7grM
4q01Tx4WmlbpUpXE+XQA+xolinIuHevH+o2ikS5FIoBu/1vsRcGfpUoSJLbu8Q1O
hOhpsGMjsQL1EVT9aWlW6/iaeDZGQ/SXKGprXOxv518e/CE0rSrwzZtO8H3tqG9S
VAy/JgsEOGMh3mViPhbaAB59rnMqVtj3hSa09vI369ZEOOkR/C5yDk7adK+9SDCn
PFw7Uzt2XMvBFjIzg9cs0itRjI1MOJAvZWCpMkAN9YL8pOQklybqS0rg5+n8z2B4
ejKlVfwE4ufP08PR+5nbToZpC6CAKCxSoOKjUiPjy6S/tR1fMk4qc68XdZJ26n5p
MBLvTYXSNstdM4y3dyykLrmhWJdGcY0QYGiDbfxwq/zkh3/xomfga5G/NmixzF+N
YUjyYTY0NwTrBcbzyQb/UbW3Dffzr0Sg3CYx+y/ph5y8LVgbLpU8kPbNLXAmRDeZ
wy37iNGqGxOjrW6Qg6XUdNDcQSwY1WJr8f0KuoRBK/WreJdOO2YgIAIeiN2luqLA
PRzQHDOiTF+RgG5jcDKSKkadLgyaiWUcIk70r8iwxBr1+RwmbM3hBXOVBFMZnkYo
M6Ssnyc6GP5ow+zwqwSIaOuXShbqNn+7LAj7N2lDB/9JtusJyHAJRt6a4MJpWvs9
SV2wcm4KijEMsB+A0S1+sIhApPW575WEn6iDB1QkAndkPdTEi5VfwNaTHYx/E5ho
Aw0FKf10OEz/oteEC1ca3w2Gxvm+cH1j9xuLKAMJ3fKsyYZnU46jwDxGUfb4QqNh
rtJZTqIGOuVdNsecHWo87P8oH4quszXff+CNARTwMg66DIvy4q1rTcQaV1MEvbH/
u/gZe+95u+NwGSYf2CbsFFMPwg7QKI9FH7x5YBRlQ5bUprZTmZkmxFwsLa9e/tqq
Ezg07qu7IjiN84EuyrDsqtutUhbjLcTFW5EZcjUaWy1cCE1xnlXlFMvx2TDrn47K
d728+wGuFJoXbD6AZNJbRcAVCX6qPeWxEdu0KzQrwZdYEgf2vBvjJMOT3I7r9hSl
cE3CfmVCJ45uKUs1rA5ZNQi1zC/bzguN0yT6jfxjftOr324N7KOFNA0K36w3fYXv
qWrjxYGRMEnBJtezMvYe2/EkxCuoGgmsJyo45IIA85LmEieggHMmEnzp599T5pQu
UXgf5CnQSFDTS8FIih2JqjebZCs8leDXdNdEO1TPCwaHYHOmac8J85Na62f6bZlQ
xWhVsawP2rmm2S8S+mCuZiiZBdCgP1qx4QZVsIGXUYRZoojwR/3Acpj+kcl6p+au
BUU48uzc3bKlWEb1oGm0pg==
`pragma protect end_protected
