// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HV7HDYbUhugl4nvaMRfAG34XyWxN8Pf4J3vpwghWS0vLiGkHLxLm0XpAfGT60AUl
AHD6QwmPGakA6soU/rHHJmehsMQo31v10MrVaavPrCE6GN0NXMrITcOsaVeeGLN1
gVbr9Bj3zWsIsnqIaB8taeXGtkn/1IlB4ZhYHGGVGtc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34560)
DYAJkrgZoulNudUXZITSPkH6gHfUTq8RnkQD6Dwn201RWV+MATzSis4yj6M1QWk9
PRtXVzZ5SfOuLMD1XB4gMl43nrtrarEIFW9Si1GXPV/Ig1dI2nNKzb1ZzbBtB91b
lVYdEMRAZK0BTxr/ZKeut3/c20fIfXp2Z/XNRrOxNc7/Yl7cYt2K3gDRGwhhNjdt
+4SAuSpm3ywqvZ6J0SisgrRIrsRgwTDdpn3LXMx+qhY8P2KaZawrH52dWG4KJueZ
jX2X4ZKTKOye7dc93epD2L20GaIYgkM2lQpD3qP67gUQgZQqh1CSTYtkfcIMI4ip
QtmZjJ3hAcB9n9SB0FS52TALHJk8yWEl8o7nS/ooW08IrEovceKshSZE1EejsnWm
Ja57wBDMU4VV1r3ocKwpEZMQC6MLTvpHgKc1fsKMIXLJabzt1Cko++G5ni0dVNkF
Qj5dWWWiAwYocKokBI/vT2eGj+DIaU3NMG9lVsogTienJJBJTpqbGnCHX52ZuezF
hhAG2RSFvar3297wkUdMyaFhgqwKlhNdd8/EtcjGrwJECOab63bOuuI2czjdmLTu
zkDzLNOwufvgEfKNhgZlcf/z6SgzQ7CKFtk82uUhDW0ZUKNS04MHjseA79enlCAM
ZOsZL0tSm4Fu2i3VMEmnECTs/Rtuk3uyibXJXCE+mT49iJHRrDHXrl/jEu8HpsZI
s4C0dJQDvz3+E74wDDu88iCaR08UZHFWSxvSgiROGtmAIGmCmIkb/seyxOREMCe3
JJfBBEKV0pr+H9EBFKDlVcgsbOGjmil3iXMSkiBAYcp+5GBQWbHBE0SpLUe4WDmp
2fH57i+7Wfl/xB47sY/eFMyo8PnVJbVRF9/izpLe+t4jkosCWkV30KuuSYAjFF8M
pyXXIXIpBK9XE7Vha/fv0legPO1imvVtNaN3UCl6bYjXTssin2aoQbHhcmcWTlJj
959PspTj426Ml90an/AZggGLfDTGUs3R/8gELbqa+Rk8mmTs5HF1tF+QMOeGqrqt
xKK74BOhGzze8Mi20kQpCgoFjRy6hOBqgrXS6SlsPF29CU0QICuctlMDdIkQJEL+
C7EL7ApQYdZCdX8ZPcfhoYxNxhZpEQkPizBMX/zohG72wXnbZtzyzhRkB7cxds9P
Et1QGUySiQiR6H283hdmSN31qeJ8MQj0fe5AZ4rdmOqHziknY0qn7KJhakQqFANp
RXqllEooUkTSTb2x3TFP8UqljW5+18cywj3tGtEBgftYsWMQ9yX2mQoPMoRi/pSB
CZguPv+zn8xXuWPHsGj72hhZfyMa8Mq7TSzEDlG+sA6WbZ2y5xVdLE5AI9cDunMB
47YFQqInGvSQW5LwAJipTqVrtQgKZTAE+YAUB2SwJ4SXZGsQ620buQSe1pDkwz2R
mBrLHegH+xdndOqYN/dRPplfCEQrhPiGhkZxYcHf+7ygy2GxttQtTA+paDNquPEA
LQWDYYbSCnUZDuMIAWp8XLialfI94lM2i24QUZjgCV65j+Kq3VL7lvB9i9p9DGY8
CwtKcs1ZpCtIrUOH4UoOUjrZLlOI++3Ohuyzah/1ZbkEiwpc7K8d4Od2NfWGTiA2
jf3ujlkUBb/J1y8XOGcaPktzW5aFTfmTul3c4MjPiPK6/yPVXmwi32mC3ah+rKwx
nf8SHgkmxlK/5JruyMgH9+aQpcfSZWMXgKv5tn08UKD05SxPYAFTuKeuXvOGvNjt
viQpT0C315f7JHh9deLVtkf++zW/MVEnIlXPeCh4dC5aK2CV7RBUoZAFOeAtRiku
HQdhVTbjLiNO7XHYc0U1nBSWFVjNUOjxxQ+gvzq6cNe8m1K+WJRAMIZj/jF1J9ol
0eomcV7GVIIzH1pJvolKNfmf/m/2rMpHXjzJ7I9ZibX6+zf6fECnympY/0iEfeA9
PRNBgMzfl4ru9ANqzkIPsTdiOcqEg91NqmklHvLglJOUxEVC4uXL6aBEV6ldeKXw
6WNWvQvIeaJVgqHBe11E6yhvmZ9Zo84AWUiyPsD0tLl1G3Pp1D9+ZONRr5DYxpu+
HN0u0cyDaLa5c+SCr037QySjEZ+QVzSBcaLOIyB8nXmUe+vmO1/HlrHndWFmc5p6
YEOE9kXarpQCj5dx7vVT5CYHZamF/mhRnfAb/h719O2UYdJ1oijaXqZH7GRG2lNa
Vwdz1XAUG74SPbhlnGnpKH36XuaVCuNFEgTliRALiyaruYlrANNcTRPyoQS+pQAW
NeM6/Pr/gCjNXtnG+sgyRjRA5P4xr5D7U1Y+XFFbNls9eMb85hO0M3Ck9+hMHbO1
WFN9k23MeIx87e8OOh4Ml6kwqeAClQFltEMf3zOFV06BVQBvLm39RiSJ1bDfwbGg
Mz5arR3PA0japrTSKNT9zP4KdmaAMDIvvVUmQqZek/kBV/ydeEBxK/v3HXTLy3u8
Jo7HA4bn/0CgxMf0zXzUhRcBk8gadqPhD/LNTi8vYswd+XNm8kM8o9rK4yCvENWt
QHsYWxyZLosv6dpKaRJlu9i+eHbuOSuTGSzDmYc02gRpb5PWif4z+ApLjkOtoLAQ
kShOk2xRUTt9taRA0NFIwa8+0MG4XgK5zI+5jTk/SI4nwvHRvTD1zdq1xxF+rnSi
gGWR8b6LQsVeE/63Nl+nRGbpKe8DjCIV5x39hXCITt+Eb7bm9wQOzOc64jSfkBgz
0iyoU6eDxLcSPKGlA7b6iWM8Rb07bhbX4lka1gGXgVAaQZFv3QBuKe/NfojGfo5x
QVhtewR+OtiRlMSkd4z5iTB1NlPDMjtIRB7rVFx0AEaYMOcaSfLTIKedtTUkzvMc
Ak14yWhPKYjVYVtHagPUB2iUpXPC45vq7yVEf/mNSoZ5PxkKAkU81DJ/jFe028W3
9u6fJx3SMNrPmmI/trnjEr19Sjol5dRSyuDNEJYJH84D3t9BzJx1eJB8UhEwEqMX
zQN7c+yzn5RlKOeBYJV5XsJKedTHD/JpeFb17Rq1M58lpKyRzZ2csPzO32rxW4hn
vwK6ESIJDm3rdJtw3rTcDlC79DY+UNE6o6lU7p8sVdzfyzcx6BPwgVZ27sXaxR7H
YtmY3Zn8g5udFa1YufDOIkE1a+T1rN7Zh5tH9WiiXiOZWUJzHLZMfVxoxwa5bDfa
cMJ1jHENkSYj3Bvc645nXIcOq/cRpbOQX18jThe/twLL8LV70JS7SOWPOvTMA1xA
Q4mwvDCcEgJBYyj8wNjPCB/WaasTxSP81V5PBugOi+SQQnp0D14AxitmbZ7N1JHL
k6wm6J39p3yHAUoWUDkNPlpX5KIvMzaSFzBI+1mskaQMgjhYbpHVHRkj0+kqONq3
I0UW4w90Gp6fPRPwwf8td/W6i+sOYYgoknDY3s1lJPojT7nWxImoTy0Mop93drL1
OggmQaSNEgMKb+ypmKh3MkNW1H/7ufiOuMsPOdyohyw5vVqO8ri4va4xZWcAHA4W
rBdO3CvB+T1nn+YAnlCsgRKeuAMTOTpRzHGRtVQcwXmpcDOQ9sHXrwxUwoOn4Kr3
/LtoOxgSZHTawAEjupNB1zrpqFTrK5TCWO/zuUh8fTn0HJfJpCtWG5WYw2yJeNUs
+zOWoEh7nocbkzzy1q4Xy+5y5Bchsyiufa0KE4fiyFYsn/BJ/8pAHkeEtfygKRZR
y0ETLy9RuliXrfjW+rW27QWhszRfb7GidaKEM1kCPn85G6tFAjdvg1L+FqxJzRiC
lrmLB0Nj49m+4kAbxeusKjWCQ1zNYpXPfsSlVKnyH+EZtGaCxKfouzwCNvE+58ex
ivlFS+s8qz2e9pJVyL1Rl/hFoIff9nxb5jIV1EGu6iqNRKtcMBhJN4pkFJ2hnLBX
DigQvlwefvoyrhaKQCx8ExWa0+/qyo81Jh8d82MooV1fAh4ESC4LaAhP71Y0TsHc
s1rAHo77xSx24g0qRTHFWMQX8nOmf88rym599rki5cK6bJnDpJ8yYslCRlS5N0cK
btVvEaTUBCwgsVyMuhy1yMC7A4ZYGTipyFHk2UquPdWfNHOyFk6qbeOQgPCzRYW9
s0uaVhsCIYdGwljWrUeUYr6gz9XQRmNQNjtXfjtvsdVPp63qVTQdb3oN8k30qCKL
BM3T/yQiunpgJtHDhJ9zG+FRMJVkwz9LgqBTYRbViUVPN0rSn7Jm53ya+6N6Oznb
K+7sBnNSWieZmvYwiERZET6pJSaRkszzRFhilr0qIiloRm6qLiuqQysyi7G4kuKJ
UXO/RzP64wbRerPDtYK0w5E49jwiZEnlbeq7RTdgNGuLUn8p63CVmag4RU8hRxUE
KydnjAMzi3ERY55xYuvNh6nKJupMP3TUd85Jjpo4dASWkQy2cj3yUokeNlsYPyJO
3M9yLdbZBaphVAoPKgXspdrs7+1v/7qTTSN1MRahapBzT7Kob6R8gD301Pi8edJR
JOZFK/A6fRP8rtXKmvKOvh7KVvSGcqoZiqoW2XrmbElJdg4nX9mJbfntvBOs2/a1
RRgvN3wNhROQtLDCzB1XWzHPJB+dHf5ur3cqP8aJ5piagU2d040Bg08sR+srWPsW
YXazCucxG3sF3TtQ0InflIRMtf8+gHM0CdkDPW9l0CBXcmCJqaPtLK74hlQa9J3z
nsDC2KwiOwk4nGP20cwOG7aFpx9jNivLzxviRv8y8mMOy0H9axZt5+S43+JadXQh
oC9qocwKai15WuGfTvJMc73HWSqWvumJYr3miy89tXOSz/dsP05rH5dF9MV0X+xm
hPikZ7m/+wor7m6E0sU3mr3LgWyoUSocDZaOJZ+yMnXmG+HQQgwUpfNzMZ9ALp63
jwaLwmkzBjDpdb1L+8txb+3eoO+hWc14aMOc7RDndAs3Xn+gC3+vTPpZ/U2n1SYY
zcxeXMkJEBUyRJrAZsxULoI3WnpYg/5g/u/YI7cA1hODPR1PipETfRMrbIVdr7vi
c3VZOkYHSScyW94Qn6kYKgtM16vp9TicFwOPJNSCh5S2p9xhdHDpr3Qiqo4AO2b5
unmGBUtZZBLgT2ksbwIUtWwowvqr9gaQ3vNaDpmidV+jAXtShMFWHsgqReuSmis6
ni7g/8fM5LbvrtyOTh2rRegMcTsuGU4ra2u6zYeDXyu8B/Umkks9S7ZQOLrCkTz7
Fy57oSZoTw4YBLN55KAQi3UqNpeb5eTJXcUV2DdPO5yDwtuqmneh2IAsfmdblMIk
VBoYNO20UeMKw5miJ4Yp/d5yGJ3EA7PQYl+b8ZQnPMr1MuTE79CBtzUghKO03ZMV
IKoh6mOsvsNsuvzMaZtiKcTJomAfwCuyVe/f9jURWCveAsG/pieY+rVO3lkkKLLV
dYPNfwb2ItVvbHLC1gFjJf8leIDc/zXPj0WTcb4ROXtn6GSST0qdyUJx6zkH8SVX
ZbY4V+GwXAdzyjrioQ7uhT6g1CtImyjeqqQ+hjeT8gjuMLYrzJLe0ZQ81l07FDrd
V2fwrZ6t5+9YpfmL67GTl1xwEQoJkwrjPaSsMWxc74iCUR147TXomOc6xehWuZoG
qi4+daIAgzxsy5R9/9qnBfyTnTdPPyQo5PBN4eJZq/ne02arYUgp/akwpHb66h8/
SYExDDRIk4py6cskUQnAHvXZe75QgYkkMyAKoE/M/hHrAFFifh4ZGU7oE/ETYwwX
l3cQDFLoqj0bj590FgtneXzQA2UZxMR2o+YAUj20ultAFkQfnxOpo2kE/QLRrAMS
5tgY4GRaQ0N65J4CVkpKMvBH/334dsy0z1U8nBwND6S/3Af8qPTvL3OdFTvv6yhD
IIV4EAC2nT3gCpCRA9iI7u5ugcZU1Ii7MlkumxfgSOifgNIKjMZDKwfDypUZdiz/
4s7JcfVRlQpt7gMZ9iAL6ctLBYTJw1e7Uc8RHcJbHJm/AP10WEBZgtXromTZr5jI
JJs+e9Sb2APnFfPj9pd6ZkJ412W2e/2Ev1IiG+Llzgwcy+xXAEjSxqFe3AE5Vh59
sMJeLV40UKkL/C83NLfmpEKWwBEkOB3BsyE1nPXbcniy0ell6nLgD3vz+bjmzaT3
PtDySjUUTNTMVR6ob828TgqdALowj9/orgK9M3cKE4gl3ZXBMvskMImPD1RK3Pnf
t+pnpvzsgJC0lrmZT4WlT8GqdHbobFcvSE52siYIg1QyjCKRV0rE6FNIL2ZureI4
gMnpPAKZci/udkUsSJOanqHfkp7EYimRmQqQYXdte8Xb2WuskaBBI6z79QHQWr11
Tr4b7limOQvLEYhPm/7HPLh2tN2pyduHvdFDCz6G2WVgvTWCsZm1x7BgpEFot8GO
hMPfij2IiPq54Dc/u/b4I14/xtnS9AzOKX7yfQNhv80AbPPNJDs/S9EQq8U1Ghk2
I181iqrt4Ag9k1RqhEgcj5UzqXo0wZF1riHbaSpX5ghiPKLVzbb3Nesqy3O3eVJF
S0w3He1hdPKsZH12Hlwxiiga6mPtXxhxwtKSDy0uFsMkFTWXk9S4rfu6XYE1gYhi
pO8+3Lkfjme+V9v8SNFarl3+2CaPpJzk0o9XtMKiuBpXkNSrDBKGARBQgnF39iVd
khsPGnObOvk4qop0Uz43PHAQQrDLG+8myJO/dCiw/Amno5pAfRizg/zPAJC0Y1lo
qTOhOTmvBMDb+Eh+jAUeA5LvD4L8/TjiFrAtqUNgd2TjRnvlxHmH3iG6B8I6Q62c
3yIuY2Rw52jPntAgD7FS/BvjKZ0iHQ+yqSAUROJNTjpQETTv87/yaXy4ZXanv5lK
TUeIAOV2n+e7GYiBmFpD8y5DLIIW9tUfF3k/sioTVK37AT0yPvCXAsFU6NvS/QYR
coE7XDa0BrJx8IITVroAshW6sBO5idO6BG5XpgJ1ifAM6kqLI9nokGQ0kzTbmibX
n2Jh/YZXp3Rso1xppq25GjpfL/ovsAmZXlYkF5hyWpcb2gg7kTSxnWJWc/McRpav
X/nQBd0pKZ8CJG0rcPcT8TAFIE6ICIyQPkWT2D2ARl+d0rD7DqEwnWB3Cm1TR74u
9TGBpMREUFgNPIvJlwP74D7ahH05TOjAYMMkICVFwUsaD01os5wtpwXQD9ouutjg
h8J49Vtj6h6EKBulyaM4KUrGLwR6qDu8Ab81XNLkUOb250zoZy5rjPBdgk8lmGkc
cWsUwH5Fubg/4BF5gaFf6Sb9syPQLJOARWkjP85OUe+VcCZg+dtZ/khHTyrC+RTn
ciPNm9AbLRJv5wG9OY+lh3APwewTnLgIa7H88rYE+FyL0MW74kqSnOAyqUh966C4
5U0b8CGdQPoO4VNubhWQA5er28/Mbb5kudapaymdpays6y0Sn1DXVKI4Q7V8JQTe
UU1OzLAoNQuqt2AiUYDg6ZAdjjbB7qgo/+GDbZrjv/1xQtIE/dWYDaupBPGqheUu
gdU/OKoN3cQH6B4N07VRP3D0lcX0uZuSG1+NdYq5/lV3m/osZ/fSzZE09tPPQgwK
Hsi+Grtjk/ZaXbImdX9rcRfDgNqyCJGSb+9sBtGe3EVSMZvEcUBDE7gf1+d77eio
MjLANvFv14aXsZWddaOzM64TbpY8/1Ge18H0Ec/xVsBNBfUEGBBDkjULWDiBqBSV
YaIIB/iZ9z+WnBj6lP7INn2k3V0PJJ3VYnJB7s2QnvmeKKK5QoZqgMjEjkr3sy93
+uMiYynxK1WkwaA4pzoCcpAiU4XjnRI3LCCNWZJ0V2xNydMn1/8uoAc9hesYeEN4
ZLEdXTADljHCc2CyTfxwnoBujvRFaMtMg6p6HW5hDHtTHJ4kyUJl86FmY8X6iqyU
sVr12yntiyFl46Fp9paGSx6QqLHZyek9aId9eHEYcIVKaT8KYxCrpIjgMqtpupcS
DJfR/EM8CBmIsn4qL8yMO83O821HnDMg7Tw7R16VExNoNhu/Q3AjybzJjH4Eke5G
QE4vHroS44m/F7g/GYaKfAUrc4Lca7vOot1JYOXt4JEBJGE4Mx267o8tnc1CXC2m
ibmBHI424xwtBQK80UN6Fe8iQQqo/HRkraXLzQn1DPEBAhBArqnYVR1+p1aiFKDF
JgHXMY2bhAtwT8M1GfTmwHtFkpt1Q4zkpuzl0mKc+Nr7tzwPKqHF6eCD8cy1XWha
iVa86kpwYcLMOI3g/gZQVH3U7ezr+B3opc025mvRTR5zDTQ3NqndMHYVzkxIXfTL
e4k30FYIcrj7lGmj26Ka28CIUhaFmBizgHomEQ/YvX8X0MTZIVDovrd5CvhyKI6P
30S6cweBZDnU0th6zcXBac/plCSOMPMr28zpcQGREUBYWZ3CDwg6BZa0Sz1ttIPa
kvAiTc3igAlKihZhtEQXDubZ7r7aeboWumLFLEJdPwjqcv/x0HZnxA5+6o3RASj1
HxSb6o/tvPCeEisrphjTrJp04ryQDSoDDw3d87yBMGYY1x9hb0QKUeEWsMSrdwRT
ZrBWnw1QUNh+74+2AE2WQHGTiQ2QmZGDuUUnxpRdS97SV/3rzb8miP/fSXi8UlYy
MfQ93B2beRH9xdwqsGSCAjmTr/KwfhGUyhXR1yetdeR3F6djrtLZcjV0w0LrvGyO
EAps4/CKkskk5cgJNBGtvuBB+M4bTfk8Stalwh1tueEc2R6kt43UMmcKJhaVUzfb
0jmFdZrws7TbgueL2X5pOEUhWGnUjmaZ1UCipK1n5vNPIWonM2u3b8xIf13C1RKg
Cc6om9Dn3Ieutba+Cf9Z627X1UagoYGFHRva8fmHmRbrY/DPT1KaKDdH3yHyd/yp
0Z/mKbOmaj3bMQSeCYVs4jxrSpLfxukwLyPRxEXs5Ez9bzka7htcO40PCYxuc3Eo
2DJbjKk7KEzNWAaYFmqeXC7qXgiACooUd9ieTLlyDXy9fZ52NckSQlAtfBS6T0Np
VeB/0f/y/dJGB+uQTyPOaStkQe/2PJRJo13TicrIbqTdbU2W4BJpfPLzJFx5BB+5
BcJbg4eDX8FDVlpmo3mWL7lm6NLwXKNE25AVh9a4hWqnMOURH2pF60EKFJM6mGaw
j9WBC0cjDfuXUpmtqqwpQVeAaBRxIF8HMc+Nr8Tvk/vIJ1bKEpUfSu4hH27kyrgu
EVEdXju59Pbond1pi7Ig1aL02kpTbiJ10IoyjEx50wpuO0uqecc152R3yZv2/6dt
RkzIkba9Gzwdwb2baPLYGTRhBN6a9xkSu5fn4xHVPDPRWGNT+tZ5ql0e06nmd0RW
hvS+xPhv9foHTK+f0pRAnsJlkDDpjN3cKBm05gluBZrVvCBYtMdw+FiuslLmAB/1
AjYz3W/YaqooWi6eduE2BUVheTC4VdZnitHez/4XUedKUX6CDxZCQ9znHJknfmuP
0McBQ1TzR8WgJMmbgeWXRzXaUd/mifvvXnUgmz3sCSE69kFLIL5x3Hkq+p5billO
0qwLT+BotoeOEfMQ6ERwqaFfB6NgR+Xjr155h6uTL58wptgdidDw9SIvj/UH7JYp
rOIquJUMMu0PjIt158btxKfYRaNf/XZAWabMqIWsRr1ql5HBZLXmoiq0IzG6A/ws
KAobBdYLMIP+rku2hRFTGSMAOXoMwtcmFelqfhXNL6zn8dTUj8C1V3CPnP1Og8OU
xZDhYv/BORaB1WrBOGPw8wc4/rqfylUGyW7/j/NxZvWT4M2VF/upu13PfUylpYfq
DcWA5ZwMJEh6uDXN/ba6EBnrFZU/xQ/+buWGlb1KtxMFcnZM9/YxdkkRttPnma2N
DqDKMlcDICl3xFDvR4cAEqcOoyWerbwJ4WYq99G92Eg1DPMHgiwREYNWu7eW4Hsj
5N6P2sfzHGvH/p3qxu7FU9WY2M80Ie72i4iPwXnNKrD6T9PgowJS2DNRc8OFx3LU
MPSgweuM1pMHmqTcdq0VjiF6XdlO6WEMFi2jvRizOpQBzi5TYG16o2WmAG0cEkcJ
vTouvU98bRtg1Xjr02eeiWvh/WOyyFOETlSHq0oPnWOlkcTmU0UI/UmUkicIb7Yb
z/JUJESoVKHF7J5zNpW9/lDQgT553JI1P+kr3MF9CITDBcoeXypNNXjpX5hilapY
wDQ+f3x1+rTPU304FJ7b+6pMUOuV+GP9M8q7vgM2vgrDk20GC2dbrXqci09lcXBy
iUSrlfJ/C7z5pgCuqueYVulKYPb1TIUXjRWcse3YBQspxwNBxXQ0isxRRcuK85k+
FWnPYK5kiji+Xyv9jSdKjrJmZctzCPVi3XsfBGSbp+p0E4HYm4r8lYYQBdTBR73I
bfbjBiQFbdTk48Q6oFBEA8tIav8IfpzClv9z/b72vtbaioTOXxoFdgIvyoM4et8N
bA+n6fyQqj/VwU4n//te0mUtfFykimSUkHPzuGjarGlnOxGw7dYBBniQwgwNhadZ
43dWJJvTHk9bAIrtkeSTdx30a414Cs1aFzJrSj2q4XlRXvWOcVtWjB8xVRXMrc4U
ip83RixmYKnr4moZds5K6v+kJWfH60rG3zBAw4fVsRprwWKsgcLhsVKn8XWhn655
cLoGzG5CaGE7LPD7Q1SQUrlE+Zj9vhiEzdiIsy20c6P/7U9N29F10ilQiEsynVwY
h345dCDv7GAvW9hXycMwAiMkNUMQ4Jw8n+WZmVcklVJvzf/Wq1SXVaEDytWApv8y
bouZtG6+X4gQuZIqlL+c4mQ+MMt1dfXox9XlKbkZeWRV2IyY4XtnZW0OIG6BGBBw
coE5hKRC+OwRnlo6oeVgfSY5YRY+k71gis9Sz1cID0aQ7CuE9Df8WvIi7fP3GMw1
Kf9MAqHXMSx20dV4gV3CITAKtwDeN9w24/1Ezu5kDh0WpbGW8K5RUwfnaidZE98x
HGo6uJRvnZDNMNKrWvtOKkSTq4YIqmkXAncmOTcSkIWp5jeb1HdpZgwxJA7d0n1e
5YjF3TSdIxYzticVsgIRhrDGTbV4sBuUEZKtV9xcpNCAo2syWwfABbwiaezR0D33
Cj1veC90E4CZkS2NTDG+NIrxNQGwsdEJwSB408pEpzM+DLShJ6THq9U99zW8XARw
dX7bWSOWXBL84aN6vVY4dawA7FQiPvIptMekmrn4IFSFn24QLqkaiiYfMEJ4Q++s
R+Helz2tGjCqX4YcmsT+1Cd//qB1Yathz34SKppLlEgljnBRNRXUJKIGTAZhdSnS
P13SEsJIyTd8m3nuw+xqc0a064j0kSsKC6AGwUHCmAExpofsedElQgeV3f9N1xkt
+BArZxVlhZ8ccWu4yet4KxiVQo2FuClUqzbmHE2XWGCgmZE34Xu+TI6VS6DLOJLc
s9/a+JTC1fxvrigkZoAXQBSa9jgAWlOSQdKfbTz+22h6xF4Mm+Ge/o9UepM/v5IM
zIYU2az7tVDbTQB+SMsUS8vsxHHnLiN2G9B6y1h4VMau3yuEsfRSfRK+oaOURW9v
h2UFywjNs1GSDBDd91PACWUaDYNKiiWSNg6OfmzEaYKTCVWYnWACJLxJkTL3+1eI
CkhlgdsP4rvmJGHoGwtgFcahVEJNtP4dIIZ79YcEOYJdJMiv/yNU4+aQ5P2YFrih
QRC8eJ9tPgN2POxjfLvHTfrExW6nJ2awybsF+VWwQNNsJBvJDtf5xO1aMsNEr5zQ
0d0mIWzVzIKjNRigx74TgG52/XwCFXRe1XZTEvRLp1FOKrp/r+B7kzYMqtmhEcYt
sgdvsW5q5HVqmNrHqGz7o1H4v6mzAHh97UNHkQbXjEZ+onihhCEVpqQq+C3yfW5u
o0CCCR/SGS/Jkp0z8TE7cWaFVIbZu7uT/UIEaCFyT2/sGLcbIhQHzI5eUVE68Rzr
9Qs8owrUiuoQ5ssFT2jQgFSAMdV9S7W2W/Q2c0xnXUhwoFQ4hbr5UFp5DYhlEOjh
DU8TN7AqNqT98WtQ+5/kP1QiszwDN+ZfsQ2j+mcdmejLXDQN6plsLOO1upL/iDj3
CSzQpP+p3NBiRfBOWoUAht42Pd990m1p3nML9Q/tiVfnWnSUpuwTSneHwB9P4ArR
NV+0D51teWUQrhiAkioxhclo/8DGklEy7oCkuJkWgwVa0JnHGNtErIJSMYdxDLmz
4S7Lj155tFR5auQDI7Hq0DxAcELlSfa0kwBQJGbf6rNNkety8zf/R8Lu/ol7Fx7T
9TG2BPtkxtrgC+xK3umbSYdsxziIn0pCcM9Xc7HFwy9Kksday9yrSYIjQ5ENvzaW
zCClhmQGDmFIztT3YtLdcBmoTphTNElT6qdAgcw+w4kf7srUDQ+Dug27wsXfW8GZ
iIEA4Vpdx0nRHwq41kjBHHSijyhR/JXbRwDIX0OUkzu1ieRtdgcUAJHfq32wYgNM
lQ3QFiS3ftF3YjvEbAO7tyBJvj4Bvm3u+RTYyKGixMvAa5JnmFXrv3OZF2qtacpo
7GGH0C/vXrFkUmETlqAvMD+snrDjn0YsJK17bbRnGQMUGg4WzPsA28KsA7naBa+K
iomWgslqQhEC5awd3Vaqj3tKKJ/qe3f40O4xpNkQ8CcmEMgBkMK+cedxwcofVoR7
cwWZNoFoaNa0mflCJzu5L2zBtIDz/Qj5yqDxIX2mezwYGljMjxQuQUdcxARiAXOM
nN+yI+VwuSVv2hQYQMKOt17GGnMg/2tHSJgjM0M/L0pXjBgaV5c22IBFMvrjHttY
+lqtXT/MOkizEp3HduN0/wtWdajjK2S9rjfuXejPn99p5/CTaHgn2/4Q5pZI1s0C
RlvwYCXXZ/hegsTJLTMe2OkIVJrWj31J6+jiAOr98dfTU6lhaS14fQixbqrJ5GWM
2r02rpLAaOnuOJvPPCXBASkS6WI+Uu79fIz8uTSu/l/fN27LuZPPU6RhPyKfAWsa
ikWtuZkRGXVGJ6503c1yVjdGJeKy07EQN+/6e0tFVNPI6LaMx6hj4BichPnqPKb8
RfMzwx4lq6C6aeiXMmZU9o1j9rK9gBxAjTfELINm7Dhgvw9wzQpzs9pUXIZSz5/Z
HdfPq3SlI7YLW3SF2TEQUObVzf7+MCEqrYs6Czxb3QfayNSJHVOrdkls4q0o9maQ
A91GxdaDHILn+sYjhRUvD2W1XiMMXTjOo2lrGQbP3i78eOHx+bRW6j57LLLFZiKb
6+MUZJe9Rh8xVFbudLFHx6uBuIydGYNJPp6yKz95lK0SKJ0E6t6zdcTg+c9KGHkP
dQ+peI60rtBrE1oc1J6eTmhGZk5yYzTjZf61gi3CXMz8Uc++XhVzWKsD3k+98LqP
VA0nFaj+6+8pfzyEhaUTB9ss+JR8++nZR82nRUrK0S+cZNgqZGfRmUyf+n1QWtPt
lp2q8em+th7p8u7xTmcWqmi2YlYUoCaNYILeaD8Ziil9U0YP8sgKZfXHUEyqG3/3
yjvOYVcvlj53rYlSb7Rg9TVmPVNWW9GdTn5/KQ2kJ+78MRY3QtlwiTGslZpx9Zl0
2JwKql3maJECozofFARG8GImoIWIfG7IU3AQ0Dw8+BmZC+O7gbt75mxGdR3392me
kpt8yBZsv76+11KQWvmwS9x6Js/V51AvJvrobgpqq6GZlkgpMv3ZoLv3JAD2DNy2
YKtGthqJ1FNItEP7iQ/eAdGkNwOffDGTMzh2yn47gpt6fbkqsMHJ3GJz9KcGp69L
JXguU7Y9PXK1cTkY2sltnnQJiwV91sCTX/1zmSFjqZwiJDST8fQ6u2tTkCZUNiCR
3oCfqIYOZ4ZZTuBI8IgFU+Dd6s4vKa0WmoyHr/MK6F2awHR6h1CQTdQlN7KF1iP9
rCl1KNNN5wfF+GQK3YLSedyBtyckhihw9dTaD62nOYR6F6i7VwHNSF+bJpKnMZaG
RgeqwHR8vc6VawxSU3OeDCrqXwl4vMnj9WfnX89Y4/hy/J7aG+o+7RtS3/YYe+zO
iHeOju+u3R9hXm5PqUDNx+rKN7cPBXSj6/v9JoatsEzZirnidljBZq+NttAp9Gn1
mDW0rYMPXYNKgwFOt+jckG44mJmmzWSiHzVoJunEaMTdhBglB1B9TX5Bqr4WXBWI
D1Pnps5drsv82EpN5cn9J97Np3NV7WVAnQ7PofrGSs+eogqhMrpo/wcQruQj6cb7
TLZwC2bkoqiwW6I094Ra1cOkyqqlV6fBFD1RrV5ozWC8HnicUxMQcxCuohwLuGNH
nxw/1WVQNbpC1NBNKcs/JkpvwYGmACVdYU7QECVV+I6aX1TDZFSEpXqKvK8h2DvM
JMiAhxcrEMFrUczxrPNozbowiTJHU4+dARloZoArwf6jRTTMXnvj3apTY2e3LzV6
3Ho1ysk22gw5PYvJVW1ql38+vwd7PHIVd7ifJK5GqCnGanP2vU/hzS3tmRL9FP1M
o6S5tOu9c5fNqoBMk8ko1Q3SAskPIzyhsb0U42LfO4C0kgLngjxYbOePXDFJKy/w
FCyA4OCWIA/aK7nO+XMzNLSDLxJF4dkOxWU6kLj2Sr5cbun6bGIlwz3/5uqqoiWY
ckLglLqm6bwoAuyyet376cjnRTnGWjU1+HhIRU4KCopHmDNYs1I4jFcKadgxb8eK
CtvYX3B9FGACiTEKD0P7FlloMRf/Py8+XW7mZOk+ZgG+g5fN3Et/rMYRSUGDUnzE
un6ymeFcMwy32Jn75In1T/IIWSBM3L8ypgH+cFoP4ER8gzWbkVVyy3kLCSMFYVUC
LNVZPopAI60VBEmcmXe1lL9EoWVMqEW4dJRQQXg4+8jvxyzpmt3HocSZTqRENk35
5zaQTJfRQCiFN4PJfGyVr1LRb65aZoUSJLLs67cGrQLeaanzF4gN69u4J6bt+kv3
ukNh755yxiu8PYsjozv/YS1k/mlN+NG3mBiGuUktv2ZHb7n0Ofc7+OTbc5PfULSa
TZejpO86DvmvLvxynRGISpABIP/dvRe259B6+bJZYvl4GIBnSJois3V2wsGq4cYn
9mKqQdFPdh7B2X3QYiMQf3gMyJxaCi7FXRpZ0AwzAXAtb/nKFNizZNuYSr+Ydd/A
MhUClGNpUmtQYwv3FfJpDempIJxmiYLwti6zpFQ7q7s3Nv6vMpJQl6XL92ALmfAQ
baOby/e9hVsYP/EcTCa00LD13nVIconUyL5QIFs38kgnDOjfn86Igv6PDiO2AIMY
q0zvehoYMdCXtzVnsBb0y4QBKzQzDycAuyFy64kKjnNrXp73UdGb59t6quKZA0c1
WpAnV89CBvZoHoSKLmv/IdEv16pmAU7VtLymSS/HH0fjslF6rf4wNi33pz0GD2/L
yy9LXN1SpGKeUk1RYuBXLo3KIIujc3GXq74zPSWRwN39QHdhUfOLcmNm4JE1QW+y
QzwEZIJXe1zqZ2aNuDhKld/Ca20goL1kKe5KZlRjg3n3RgK4tnO51DblkAMRQ2md
u/tkh2Pgg2E3Zlmo4totNeOgkHw7JdZ952tswYnIhc6yels09noGfLQ4jUhJ5+YB
ErPoXFjqt6VL74CTHESKp+yYz2nPMxrOBMgV3t8DvvIqoMUbwIgF9kXFH2QIQuUN
ftrDazQzM5aAkhK4KnLHrFAPaWcwyy2AvJjOmMbulQY51KPGwZAVyAPoZKrLO5pk
djCggOhTD+QBNsKs5REtiWygQkyRLqi4ZicaaNsa7QyXu8wjUS8iHuwPT/SBfUq7
9iqX1Xm9VjG+QYZaIi/QJc0I9MaCfbOmP2s81onVjjHHi252cLe5MuKGwWiu1AU/
wDKY2Bc6jXhEbotZtDaKFNOCUbqIpnz3Tj00sLhL+ZVL1z80MmCly5Y0qsDh16+d
qbzAMIYT2TJOYIs5aypG/a+kFMPKCJ1OeHN6kMPE57iYF14r4a5IsOVOHj+8eV+s
/s6Dlzzf/lFAMYiBCWpzaK9ZiSbCthoIw+5GQdm/oTl09zGHFtQ+xtXjMa1sbbeT
aPIYHWHkeU5bXRVUU9uHQzvCShrGqdk1xiJ9THL27ratBcXyBBpS1GzfF3ng0OM1
nlzNuTm4r4dSg1W1fEO4PQaG3sFYcp7Mt05+OWnxWNL7oEjEYY5XJtmA3MCCmiC8
NGN1dDJJIQxqBm/IEDCjKg4buwfXCP5oMUTIGzqBjAB2Hg7SWjU3ydSo1DwckyNu
GWj0hmKmkM1bHdzScf9dX2MPn/mPik1vnU8LJvG2rLxp+rc2IV7bPLnrfxmGX8pq
Q0rIk1ukm5Oz5ePAXITz6bF2Or8/6cJrdVWXEvpYjutR7VSgEYbs9u3nz422JK+g
v7TQymYku4q4966G+rftCUxTh5XzdCsqczy5Vudb9RyWjWnIPFM3b5Z60/cichri
oBXKM0NrAuj8Z9as5k/PRiGOD1S8n4Tg1+OAc/lFoCmE4e5BIs+2CGBArSaAczv5
21NyVhSjRpQHhXao5BzVaRiJQyjv9qTyRHiE56wzjuw75859XfxEPzKiwV6i+Ivi
67cfeOcaqSBFFgkxV90Sh8pcemoN9IPgbrK+mPSyBQeeqmJ+6AivfDalvYq3+0AA
/rJnVUYCbKSUZCdUQuiEEblRsQZFoIsuqg2vpzrStaPgMZBRU8vwpO2gqZWFxz2v
hhbPsZ790MSc2YOcv7Km/ENTHuLjQ6txi05dbo61/CmXwv4qdfeJdX/B7x0WZpSB
9C8fnJQXdkcZiQIjtaH96q/4qtZerXYANKa7hEnEVeYzKq/bmVOQLSF2nKKu+Qk7
J/JIVTspe2zyV+VYJIffjHwq8U0pYKbS064nF+k3TopFjiG0YqKJPcc8eVvKiWUc
m0LoThk7NQ4VZnxDCeSF1d9eQIR21dtsbi6Kz3/muLVCyxVTdrbYul7y6DavrU8n
btfKBBydVssQmkAw/WLGNpkyYa9MrFM+YzrgFtDP9iKtczLg/P7E1ImT2/3tkh9j
dsxjSc5Uo5ZzuSGNNOPpfQKv0lc/Er16scMeUA4h/loqduGQntcr1Ciw9xgZgS7N
+cAYZLRCpQ3jt+QpCMsIIgBKdidDOHGiwm41iOqwvj8TNIfWzqsuXsuZXjX913S9
HV4ylq5X0mz0lU6+m5vFWGRp7QcDepL6wpI2bNPFrkqgepBxsR4ApmTlTmEkNo1O
j4V8TOT6tPkurcHdETjJPHK8IGS0gvPasu1Cshfndr8/n2hdtgnFozWUCmzUJrhO
b52lyg/QZgu/5TXmGFjeNgmGT0qvXqNmsB9l0vYkMLNIrep+86pkyGPSTs+7E4dh
FWOnuSI7uwbZRc774G6fBMAG1HVr9C6dxF+qSUHDc6Cj6QygPaebEQAcV9UeCo5J
AQi8wxHccPo3ab4q2IEfNNO0Y+yh3Tt3cnEI6HC+aN4ZXwxSrOgkec1VmP9zWEFu
pU3Q634NoYEihrYpmP60yd4Bs0aPlWkFMU70+x7o/cI/WiYrx3YHCeut+5NibgXu
SRxbUtEHRJ4c462whE1Rjv/EZA/svAp/4kIECc4KJ7H9u/5mxnLyZawx/95b48B4
r+Y9r+z1OE/iKycKh7I3pnfHN89RxGm+LuDiIrLJmmqg1awofjVt/AHBcpwwAc2b
0O3dPbJlP+d7Uxu6SYG7+bmsLHH8Kw//4fTqTjUZpHx7QKbh9fOZtfXGd68IkyHe
PZDAdYNn0jxgWvVGMtax1q570IvKCjXHsRhyZnoAigmtEVYeWroceNYt0qgUVSLj
3FWifGuNwPgImIvg6TaNYGHl6jFu43hHfezztGBAXcJYJWFtNHTi/b8G8QQtj3Hf
E/OavAmrwU6PW3HF26lk/x5FNfl8KNb83aL+c14IPuNCFXYo9yoCxgX+DetWuyCj
GTBIWj+8ETPSRN2ezpQ3XIYQrB2y8mfEgfNVvDXfMU3eKTJAY8arA/zg7X+ZLR5t
+AomqODslc38lz73yaqC6GpPyFXmeV4m1CnF+VehAObfHGGNJmvj2707Fb85YppU
FMlkHsp8i47AplVWeAcYM7LgMsDmPO/IqQTUYefnZjUpUjCyVzOUHeWKgSMksDCz
KTiefDJh8nDGaicH6CooGJ4Dxv3nt/reILhlj68Fb+2fH1Wh06010JOg+GBX0mQd
AUUnAN1AU0vG9clSOT5Uslsz+L8NzsIc9GQoSf8WgwWflrrfrvn06NMmjAbj3XoM
5ClRqyTO/o6f22nTY/+ZhsaDjMl011oAHgWZvy/I8hGd0GLaSbWfuiRwI4DhNHYn
HoDlpCYutIJ3X0l3uxm5LaCd4zVMv6CwrrqNGJ3Z41fSusd+inBZIVPGAChRvF8r
tFjPGQpZqW9cHGpbe0A6QmFVo0ZyXHrdTUx1npcaaW+RCAtTdQBDzlvXsMV2irYx
0vhJghkqTkQ/lLbJOT+X3hL1wrAXZ9YN9wX0N2vt3dtj7tmgP6KPQarsC45zR0IT
lnNs3nU+R79pLBrLDFaZLxC9fduYrp3iZQqX9/kRlLzNL8CXbDe7HTXqONWgLhNa
t0touK3s+3AxadihH1hHouD/u3GD8k61nR2lhIPK39pfpjpiL2sbIgzOVZPcRx0+
x4GhtfkTaajeIu+iHyo5fLrvw5n/rU4gDw5Wu5woIRa/wLgZM1hFVkLPUwvPU9/Q
+uUSAdoJKgn8I6ehqjDyispk4tJtdTVStJO+3gc6QoGKAL5wlBD2YN/GEjBo0UPW
BJEr0mExasXhyRNU2osdAEZN9krmJ6Gu1ozQ+gQ4UK8+9HULP5g0Q14U1Li08DDK
2Km08HOJn9GvkWrb9cYbhU0rXsrQ0o4/4kcdEOx6nIDO5MPlkim3EXgxhV4qoS5U
idy8wVOSZyEU59KqbapjUPpQVK0DBTDMCu87+IxO+d1z+l+lQVsu9DI2+2RopFwY
o4sIm70zwNJd91PluX2rXLrv9YMIv7gomM/DSfCB6FfzujAy1jY8cXBaAGiNePQB
c/Xk70lIZPOy/UstnPAPqqzMyC9M859V6JuYzird38JmW04IjGB5BeRbLYykqUlc
J9uccz+TqTugnQmUyKX6Ys1PUNNFkibc/gATqhPkdU1594YtgBnfIPt5jdu/VHr+
mHJhL58b9+Hh3zqyo2iT2NbIHtiQ7uPH0NX7wgnZvX2Fjhy7o/H+dHkaOYoDb7Fv
5wrQ4erdxvpUe68wLPzuXo5+tj6WHU0uJYRP3UHLWLp0pLIwwFRILKSQSQIsS/Mv
he9xu2Tnm9kjgW9MTNyQpwPLVICnMSOAmiAmoZNVwo3qFPWtyzJM0Fl2JIQLJVyl
qKIIUe//pNuBEcUog+yArTp+z8F2iAcK5nC2lDRcoOQhYrcDO2i8zDO+UhWgH0GO
azbtQbxp9/0+4EFYmYqSsGypjX7vEs0gyyAmvvvw04gmoz1Vx/VnPxICR+CthW93
cRG0pGHkGBCPXR0w4J/+u3hAj7HlHq+w6JZ5R0WakLJXXwKXGaS8+FUPMlFu5P76
fLK6tce9mHS+pBoUiWuAs0Zmlfco7/EWAzsKkgF49Vm7BTdskQJVZWN827IlfJ5V
yj33s0QOnlplbSNWb/3QJOkbigAqzc6dbaGzOGe4GS4Kagu8WLrUsFaGdcbSdWF0
OQwj/hpSt35EU3j+yg/TDRWvPo58UqHViC6c9raICTko761434L8zn/oySs+GoAg
CV+fSVdCl8FneybNfMQ8u8zBa9//4nOdpTUyv3a7cJ8vEFGalKdsyeBPqFr+z5E4
6cGFdix6Q70uk7rqZLdm+ni4yQUYA8zWf8oSbbPFETpB5onx+Vy8fkVDnfcffXfK
ouGINjqQWQZrfV8EJdSXzqxTFHdNn2FIier6E1+NOZdOOtut9lrLAXNedoSKRSAm
AN7QihwkIKfgnGGhGFux1P7uxxA0v43mJCL0p79V6Y8uTJUOslwIOP/11qAawU5A
8DOiar2EUUxOwpOUtkqAL7auo6FqSwAoGIiYTtp6gezoNJgsdsLozk4aFFiTzH9q
7Vh54XvMmQZsndeRb8iluTfrF9yVW8Mw3NAHkmWz9YnZzso4I6yE9dw8ZFHLQxB6
EthY8Q6FtRmtAbQgSokRxbobkY6VuiZrQ7Lu48IH5F1wkzNhXD/CSRKbkxWQ9ZgH
gheHrodLMYXdwZRr9VgYQ13rp1+PvcxBx6Y20mEUi5rLpQFHDv4zmx7luN/ksexY
SxekyxtrGptvtEldb1/XY+Ps9EC0C8lTtXklaPNbo38qBg7ccPOuO3BpTkJYeDyv
IafU6o4CtemwWoftBvW+bMkvcnQQNr6b+y02LHylVOpbNKGd4V8PwJ37muB/KM3q
KpII9mZ/YJez3LV+CL2KW1rGIONNvuGKF7Jg3LkqVmab/w5wznnCLeoHk790cks6
FscWMnUZpXXUeFSsehg5rOHWnIZU+O7N2a5zmcAO65dO6CLSf/2jSCCmzRHUsNxG
vNMtUy6T3LEq1d18HC/ciyL5AgrhZejCtYMo8DoFlDmGdnN0O+6mI/FtdfxOMxng
OG+s4yuNz457lE+vzT9Pu2mDsdz/i14tOZVMkeiPPXPNaLdveL4QYfuRUNA1aUyj
uP27RUD5tXeHQfZ2KznyVlAmuWBxI6Aq/zd6ioA9D0BRyLI7zr1BrRkrNQbDeJ7U
a7lLgvlljYg+cJoXezYOCPIGbZydxvSYsya1cwuToKl3+OXBzgD04gMLyllZ1Bt9
zgABKfVBI3c2MStVJNdCQuUIcgu76vcSE3GNxLHoOlNiSMVzsmku15+2Z+gsrunK
iJLzAE9j0CLvvDqlP8uxOXPfCCpEC6wIOb9YiHHkMnu3+HfGUjDyAbCfbzTGbbSm
URv+g+r+hb1reflko/KYAT0OPtYqf2vU9E3He5zoEPFd5j83Pg9ahM83fNfgdwEP
/f4P1/QtK0YNaJ/C5KMuflz0IIpEkoxy3Dj6gn0XTa1wLBpG0CGaeaj4IbOaGeLA
LUK5cCwY98Kt2L4RNGtvKTNhpKS8wZd9d1gfm+inQqRAl9Hm9tDtiKXbofPDUQWr
gpHGmvcyk6IeFB+7AA1dshj+KV3tuJH8+1dU1t1bdTGvdsB8/EDPOqsuY1el36Nt
Iq29qXcuur3H34djWPqmdk/JsiwTb2NlZgJmqkpn+481ubKFdGZkksIxOvPxcU2W
R7LwzKZdejD7ogjvSVP9HiH63goul/aQg/Hszk27xLgWAsZdg6nczIGF1xkRbAnf
/G6PvLU1FGCmPwdiPeSPEmLNWohsxGdxdOmg4Oo95LWMNANVbHwEpIr4jskSd4cD
v1VD0oAEL9O8krL6pwpXo3qS+CNcD/5Yo+8EuGFH3ZejZA5wJRRQoOq9A9ewqZEe
fJQpdjF16kq+oWum9Fl+iWjsJoYWG2ZJxKTlWc5u3YqXKrOIE766kDr8972Wdy/M
VHE3V6Bz3+iHMGkma6kxXnBupA24a/1rhQsqsfk+Msk2wIKSKI7uAJWf7ibnZRI0
0d4YzeDalP4s2UVHf47jti7p7FTy6c/Jm9VaU327oEtwovj8zRaJ8mL0AX/cbfJp
JF0sB74RyY/SgyUL7NTtS0CYrjyLTOmK3SbkzkoHr796WptcDRCk/obKjRywpznP
6pt3yxIVsqlnDHELncWtSAn4F0glCS7p/HjIlTpgXsAxE4nEPTR+Nj6FNsv8L1jD
J9HD5z5ufmyfNLzSxI+jGFj9daAAokbzNbyUvEIW/augy2veSRethga5DpMmIVZV
sXNDC+gHSNfyLJ4R388jQoJiFIH0K5nMOWrwUQZc3IsLCjT2IXZ+h/5jHi75C5yN
8q/u9vKnuYDgZQMToKHxarJLNQMTozFsv1nrinRdZ989Te84GilesRwiF1LuWp4m
RIwfg8sL7KHLI7M/+9d/UBogN0qDGFgSLUNs5coGB81xKWrxFPUZPe6E7uiGcxKy
cium5jprtrF/FTX1AGj6CjEZh484Gli4PWA1MA5lBAEMp+BEXfqO2bHH8giCbkoZ
f7maPIjhtBvQr6Q4BW1y+oe9XGfWJJQ3RD2DR6YEt8BqGHGCX+0YjAgkKwiudCFQ
1JV2QhHu0NnKzonJYJxxl6nKjJr3h32jmPjCfht0kpVPAUWTO54tYODfDbIbm4eL
rNRfA3TzAoU+iHcH0xg4SBIKlJHWagzxE8Bes71Oa3gHHYwTjHmGbh7xf+VjUckj
DZVa8zJfufdSP7Un3yRgp4J5aLR1j1MUsDXwB78xT9KfSY6nr8Yyce48Z3VZY4K4
/uvJxGPf/ZQX7gaqIZVzUL0tfoS/uvYenQuYLKcjnO2/iR/aYaYhVvGq1T6aFPKi
/MSUgFALL+iyG6K2r1rN9IOTr5AfQF2HOd5Ko/8yAaopafzt4kLUGXorrG/y0DAe
jbkAi8hILnpHva2jiZfqbBtvXjWsCEMJNkZ5DKsSOXF80AFUKGc77VMpJOZPiTxu
VxlAyXyqgbSrrpYvRl6JhgHhlXBzUWpo4WrDI5O+W0ZzxzusxwjzZg8Z+QijOysD
bZyxs3zuGmH9N5wl8i6/f4szgCOWkXH9u8JhZbaW7TrGmyk6mFi8dCLOqO9jMDNG
+C0W7qJvqNwf6oON/bmD+wetpcHJJu74gONqO10hi5ziE3WJ7PxE0+vwrEzjmPbw
yEIcfzmR8VYBcYUZ3W/S4TFBlFcQYmYydz58zTdY9Dajgzz+8k8nNuvuLsiDZEHo
ZZZKo0osl6f78tufp4JWL9Kqp6R6tTsuQQyijcmViu1S4Y2fklJZ9uUIq4ylZOU0
tXuXYLKy3JcQNyclu6pNv5FtkXUBQjLQp395mmF3znWvE6fDxKko4q543c3MyTYJ
vkTzXoQkZ9QbPI7khekZSCGWJ+Y82qIrY74Ogl2POD+wClh4ADFeM0xlt+QDjRFA
/HzcPe6gICjLTfLG+h3u4qb8R8LYXyJUDlOFSrv4m2mOKMYrDXyp/pBhVhMAtnLg
Ayl9DaY0BWvyqQQfYjJdzyS8+M5T0TkJe9fuEHhKS8mdG5M+tl/IO3G0o7FsZjVE
5zfVR4PaoL0vReWkaoFWfM9LZ6O2sspf0EZst5J3snY6kyv5QkHcKwn5h0UeYCq5
RX262O+iZfWPWlpyETSfyYFNvhubhLmoS9LUUtHXkWoYQQnM6d6gRf/7tz3loqpy
4xogvY4TsUyoAaqPMtS+dUwRhumoBeA3xnYslrrzw5Js3/U9CFpLEoF5c/gpEeYw
cIQP824eLzQw70ykBuCH6102qbUcvJ+pdpkRUmoJgWjqtLy3VdGidiwDU50ZyqTi
PI0fWtz2SydrShhViNN0cNMSFQrlbLuZTkMPl9zxIZ1yJd632kcnU4V8DnKAaByd
gSigvvufweESkYd6AoIYn4SF6YJi7YmsXtRpjpEDexFznLY0loNAi1IQaJgl7TUT
y7swM6HpMAenHE4ybpvofLQNQegJESL1nMjwTmJCDwpXF7W8uDaTAeeCyiDbxR8e
rxhNxPDJx6IOwtmHpmuZd7zBNZqH2CE9puinVypSTXnrOa7ufgCjDG10wSoBL0qv
WiOFZCK+QtNfZ1/C/ET8Rhq3Am38hVtmFrbWwLjufvzNCA2u5OVuKuCCqNCLb5Gy
6DIGH5O6j6V3sxrOMHB7P/pCL0ZoQS93Alz9O/8I4ymYQgJScipZPscWgspMbts/
BMU7tY403Y/8L3m2nJjpnVdDNo0gEnmlaNlkGW1Z4WbXzp8izT2iruFJTreEUVjE
VVab2L9qOumlGrWg5vrE9qF4fjDgDWe3gcRCIiFBtGyvYyDZQx5ncpCkmDpHqg1+
g2PLgi8nGABwi5r0auR7zVZja/+WydizL6T8FSnZQa8LOPC6YDbtlBUohjpx5ItO
FkMz+30Osf260aFQAqe5J/IOaqNik4MWFLCQJnhmsLzFnHk8weSgS3eU+gxNco+5
VsNkZ/lh0YtHzARN7UOqvlAcLNK6zRsD7VcKro7v6hxcgvSosZbVbR1AWCEzivLW
gJksd/s1BWFA7jLfzM3dsF2Mt5ssyY8v5udId6ezcG2VBwZ0iBpkkb6fx+y2AXoQ
wFGBc5vO/yX41ngNTCEaMiTn3i3UI/8noONN56AVOSvawYMzzDt86uw4zPVyFeBa
1lZnRBAFHi+pDR6F2IJYJUniJRrO1wWY9QRysSo9D1BYmMWvlvjNuFTYJyvnC89P
xDkz2L9CjGXrC43ScCv8lWAYtJviukDOSTlnkHbgrLmFH3Xdd7k/DoHzB3vV8inV
Z3n3mx8bkYi+PQzbfcZVjz/LOB5tQhtRC2bK2NW9hImfiHnppusGcfnsswK3JVSS
LWaoKtLejRNa+QLB+JmQKvfd17hbLI9EYk9/xA8DRNHuPPOWCcAemTcDuBkBFMXx
ZtJXfFbcJt+RYgMuhzAVcZemJVz5sZY37vk2CfutL4ET3AAm1KvwvAK6/NoxLbJN
HWrXMHXa3PIigTSY6FCNcn2NF/s4/2NN2Sezo/uzjj0RgpIzzjKpDQ5qRXoWDzML
wHrYKXWyzAO5O6OOp62rj4toWOwXGprYH5/IWPqhOxjCFUVgLaDmhcSHtXeLepWP
nsmYraeSn6WSkZTwAiDJ2fyMm/TsmM4sCRfcjRT1p+XsPHvpjs5Ph+KpNIYdlthX
omqOy8wFjFbimenbiRJPnRG5s9Dh31B4W94IO0xjKq+S+R5IPQ8IjXP863Ezl8Fq
q/wRTr+t6Pld3do3aRL9+W+aA3bF1IO/9vAkBA9wz8VsW1x9mZlvgu/TLWYpeVZc
QUdQmfFLqL5N/04Xe97QF/0p6zMjATPchDiNh1/uXpp3HY/zbwj4AKpva/edFmdB
0s+LDFspQtClGSyeStdstd8sF4BgqFVf7gtZB751VgEgDyTsAcpNaOj0bRS9YUci
LR+ih4m57z33SMNGlXWPta7MPFKpODO7utC4mHZR6PhlwW8eth/QXZ84NJpvfSgR
zTRz4X5HoIXqaa/CmkfK/RI09wqZGkiO1JzQsbUzz7rkF41hlbSavtYsG+rTgbpD
e67xH7zVJ12RpcL+ZdpW1QpnYsVAAWtLOZ/IUimMaSBVhs3DzXmMSO3jlzli9nes
UFF+wFZcW33f74NTN1mVImFbbbdAUifY2lsBKJwdjYKDlurf/f6EzAPCdeL4fsgA
4LA0Ok4wW1mOQNtLEqlgsDigfajbLhzikuWhEypCn3ylO9/1mP178Ncp5ZbPeh9l
K9mzSSAcrRh9pvoJK6jils4WXSBTy0XPiKqp8Csw/bYNeSBdaiB3Q2H/hgvfc9aB
8ucRKJAnDzu9jvs4/v1C48yBB8Lz67wGslq3+qzSdq9fk64rjYkyPh6KqDG+flRP
3ld96gv5C5ZFPVgcrg/qpywqkGwdlUtDfMsJ0eaIWV3g0uOS9nZUb4FWCQYBBZuG
0uAJPQw6zim2NYAI0Kl7O6xwY6KjdGKw+t1y9uY+mbF2MnPjdtwAxpelgi/F6Ym6
AjcagHFiCGgBd5+NFjM3L6KLAtUu3xZ3PsGQChrSxivc7X4Uv5o4r3nfwttfO0Xm
AAGZozYkqfQ99A4Nx3QjkN60RRxyaFM22AucQN+rVcVFOPi4ZshabI2ZT76irz1g
Af6mHkYs6uGZcw6hJ0pwTzWBYAV+5WWUjlV+AkLHRUwaEyBkp+LkOeSVjON/bkVu
K4x3ls+EgMA3jyrNg0aA0W7nUQHaNAUyWmNSFUyZISm9qmdgeasmTUPZ7nTU0jYP
A86bKa/EIv0mZDvUj+vVZdao22EN4NWI07+iQ3E1Q0hmrtMMOCf+vfByovWYWZnj
eEeIyvf4LVjVdW88IAwZjc63wf7HklegQ3gaJOllRWfJa0R+uVY6Q6dsoKLluffm
HF1317vyDJZt6AIMncbo0lRLLwdr2yVLHVJDEqtueEIBHwm2KmLkSR5rUD2x3Nos
1UDTzNYKQrxwsDamC2WfI1O9YZCWyxSPGUnBynzyPRbqcE1Ti6hIwfpidSJB0iyG
L4LkmZrdsoMOrCbGGohlASEpB9svW6mYs2TIt9hXnOcRV9hfGmgOtY4g/PldmY1P
3gMAv2/8jNE7lFFFut4lUTfB+kaaezHdayq8GGW0ECtFrBUwO85YsOlJ5n0iErsx
x6oNs9VgwryC0ltT5YqcOGLdxvSuEsPsOdfJUFZjNooWnKFpmeZfTWDaX5R2CcRQ
2PzIwa7h56rN0MBQM7RffYAOXpfYjIvc6bE/B116VY2qbWii9KHHx9u9K20ChGsH
TyMw0Fi+tmD2xVeS3otiZd7DpJsxA+I6ldI3YGevJRn2iSWn9qCBoHJ0zvoUb2zj
w5SMt3zX1TWTiUkfv5wukbR7IqYMxGxklADb6XP/DUa+IOdJshvpkhcAqxOu5fTh
/GZoZBcwMTIKnRV7WVC9qT04WdZ8Giykho7PrvkXlP1+RG3y76VXJw2///9R3rE5
zXqkiajsoORppIDujxO8mqZqdZJINrBi3hrY0+xOCGsE7gDQhHe1jQEfxcTbtYsz
m0WRViTDikbL5O2LkmQCLNLLldDQeyNyGxMmvxoNlKAmsOwQoCrwQg+xNlQrh3d0
oII6FZ1G9dV0Bqvcrc4Efah9zKzfnI4zquaIsyyJoqvaBDroHJEdhhGBGKEZUcpD
8sSUhlh4iauvLZDqPM/O7SRH1j8OM3PQlw+BFcOkfdTSEQDU5jqVfVcvTAjED14I
mV4D7QVoNju+OuTuNTX/yBmIzpXRCrmN4bw6iqgmZ7DzGO0OiMXmwRVT1TZxsH2o
zQmYNxHJYx2ZWtzOozV9Am86IKS4GQGB6uRQRAZ0ejcHfpmi+qD3MwdD3FR7og+F
QU7mChO3MOVEwAPxO1BXfYhIRYaRq84L/P7x97drae6DIqFrHfn6jcYhJ+gKIptE
dmR0qGfAYPt+tQ6WnJ7L7H+PdrtH/FZbaaIfcbeQBufG3hzQUkBFealrLAUmO3SC
rG4P3o7OGxpDRsFlbpS331i1edSfduJOChE/C4ZuGOqOeTS/fLa2265fClH6c1jq
I9l4PLUEx8WjdkhoM7pdXRE7w92EEu2Jgjew/wTDIld6gC1ADVcY7S7ZF9A8KgDh
MbTXh1jn889kLqwELc7hT77VR0sb0xAC5BRKbo/vRCWogXzGR+etozAJ3Zpl3GJA
a4mef96mQuwxmTFmZTDFTsxfY3ENbt2nhqURmQEWLkkEKrngd1+fGdA1LraAZiN0
+tLrqWwCz89E/wGYX5Gtfs+deHnSkDfbfmmv5Sov0qbATvcfFJX7syyjGm09YumW
ahKTMuSlO2GZCV9QpIJPaDU6ap7tV4gPRGkKVsE9Un0ZsvuIouF2ydRunXDv8Pha
JlTMMIbQBvA8KIzukFIsdXZSnRCNBcVJENMWo1/5r9sFtYxdbFmn75iKfeKQx6Yd
6ypbjY7UC2A4/SiPzL5Hx/SkSQzdXCTzaISEp+Y/wDKdUbMv4W7JhiEIxc4T3rs7
+9v5HCT9w7AVirM04Edv57D6EhNglyfzxm3vMlJyBwc7O0klkCqrgefYmgY9BkXT
IQsCjjNkfQskeu11ZZBBIcuqOwwqpD0+lsHxlZJHiyz7ai4qN6aUAKTstNEGXzqc
h0/k/61cTLamTUnDNM/1o1ldeOTBv6sKQjnGXRRl32iXwMKNouCTxcqqlwDX2RHP
Mr9Hikk2bZjCoZP1diSo25rwT5+PxkEJxO9z5XmXnKESTkyv8Wkyqfwa5q19vpl/
wJYeoLJeS4OjlyXQXK6xI2F2eK2loAPO7j9UovXOnPfQIInZFsEg7wYEC9dMfNNS
gY0sIFPvr3FZ6lUbn0Ox5U2N/VO+ZBIF7JXRj4JsfZ85AiEfAL2eVIT5vtwR0PYP
irPGpg+K/S98fgFEwFX//V/6xCqHy7JLE2qWXrEqHcZraISyRrg7S4qSJtrB45qn
n+sWaASMkcHO6s7pTnc3T2mIVGyIDMAPl+3fx1S0e5m7sQjRhNDP+V2LHZ6YV0Ij
qoHWumDyeSrzOxPaYjkIUZTL2gvnoiMP0RHGHQB+6YyQcYV4l5eZiuwj7Vf3VI3b
scA9IAU2XPQ9x4g6wSALJw8qxTySV+EN/Gneffv0qify7Fl8N5WKLgx+sNrivU9v
bIGYd7FHAMk3jVOOu2Yc/C8YuLoMB45E9/Wd4OwGBko7Dyin+arz1gYjgIj9q8EF
jpOGIBzfcbQ1GxUQp1z/m3XoNBBACIR0Du1/MxSmCB3NRD9Jq6ktrNbEOeQJgMjL
qKSaZbO4kwAbEPnm8hF1WooFMAa/S41HTj/E/rewUgTLLZBDPq0SOQbVcZHFE1zW
bogjgnmwSWRlgKYlFepW0gSz2U4lRNnx2tQj6rD/q0GZInRgJlgvANsGh1KvwoJi
fKtVAYqzj/TV2mgFvngG8i+jEa6hw/hWVicIbuk4BGxt+N0YVdyz+jnLHfY4XR8t
4/Iqu9bT6I6MZ5BYyrZVJF9tegAkKtz8HbLXW3Jouft20GjDP4TusQ19QvtxMYAy
CtJNfGNVfpfi5OJLZG2NqT/wQhXwq/+Mk9nYiQwh2wQ61xza9Aa47wN27D4HJ0jC
DroD/B/2ABmLuVYq0PzDaEADKGRFRxn9Dlr9ymy1oKpJXRUM4zZN9L5a7lEgiuFj
Sul4kIiERUVnlJCqN7dVCMUHKGrg6vTxnJPwx0U1+77Oyb2mzw+BON/qiT3Q/J5S
CM1k523Gb1hMViKyp85MAZe+b1Byo6/lDYStYGeq5BwE2/9IkBcTBT+HaCUNUMGf
s8wX3J8+JcX2FZFiIhL1/DMg/vDtt6gXlfolQ8ug/ejj2/LRBLv5SkF4SZJxE+oe
4DqcIke0MoGaQ2I9qyCNWDQ3Lj/fMdkMCDXqCHl9KLqYUFd5BH6fgvbQQLg7ekQm
ok7VVh409VEL9JHRDpJu/W3nUODVqK0Tiy+7jVsLvzta2n+7ajcAIYAEi/FA4WIX
1U7WY8qfmIzbn3r7e9paKzXSjcnPUdnOWEEtzg9rqNdA3N4s/pc6ZDEuil9kweTO
cxfNDl0cEahstLE1/EgctGvRBoab68io6GvFQB+xOSQNQ2bzkN9DvGTyNkaf3aTh
F0/6xK1yT1pzGW+1V+dmCu85yDRl42WJGKtBWx5ljbxWZs40oTXUe28lprfEddry
WkKp6GmLrRGy2eUtrLoLAC+gVbNTGBgAditXoX86Z9dX07n7Nh3/C8IDwfsSwLJ5
OjGFH9P8yK9cFhHpngC9gKdPKQks1kokkKVBU7HOyUDr5NljiI+JGmMqhUKqLoSj
sa7PQA4BqJkDo2QZMBbXfaHJCNO7HPs4JWgmPRhZrLqmHgIT9AqOcNU9kG330sG7
T3oL4YDkMWpezdr3M5s80ckAn6655ifNhO8CQpIVre0U7u6Bp8l9iOaNctiLNkm8
1mvz9c14xJB5cEH5BqYC26pIjJqMKNgyPfkZ/ECPFO0a/QTO6rIDHwFRFgrBjmwo
t2+pbWlO0ZPuMzuLO/S6I3anVMsDbZ033k65HlODLizdjahgRZtHz3kH4rKud9+/
s7GPc2xeJ5NzyVk/yJWJWPV0TIs2eaXciVsQcCNJGytozrNqUWGtP00gpwsndlSO
nTrrT2oSCD+AbrSCMriTVqh3ppsVJRNAMs/3BLX0wmG0tBXLWm1IFaxztUI4HrBk
ThThkaAF3O1Pyloe6M8RTafMvBZIizPWf9FuGVKNMeZmwKASCwACgrtcjNq3/FAx
dmTrpebDpanfENcMXtHZDALuA3jEUKyYgVAzjY2+4gaWrCp91BVcULmy+laOstBE
057mDzOLtGUKBNq0Rf/QpL+Btkr2Wz/Uf7WxN1T2PcQxWgKVFrlaEXqyKUUCu3E6
sV/W/M/gbp3RrS8xVPcRcfCw4e6RLdRF2UY4EoDJYaGVokRZnHBTV5tGU3upEF+X
2Z+TfUK1mgK0qsAJtqy6LnkedCu13RCw5tBQ56rFf6j05gvXz6/vratqd3dGdZUy
sAZpVF7KW9WBARKIOMA6TAET1LwZbd9l75NevetcIy/MGxBd9rB/v7y0FBORZOjL
wc3cfPIPRO/vmX1PoeALRjgYLDWQZ4JFX4xZuOjiaj5WZlyc2e5Kf9bZSOoz41Pb
QzfXb8qc9sLODg2WUQHgY0TlutKC/G9uQh9a8F4dubpm5coOk1aft1m7Fwi9Gzn3
8CK/jWmJyiJI9mPMiZK9Krb+mlkB1/N2RT5mu+xtieAbzY0wSsCdR/jhqQsgF3zA
HG/dqCKD5Jf7+RdGskOEDJZOcanDaG0ggAiXkvZrEwqCETjkndb1ByRiv4wxd5r5
O9TrNtfGaFTRnHMCi8q3Jygo2+NiM99k4mUPZVkeZANRWq0atT6JcetW8eIbPRqV
wUMmKI+OXJRxc28rXaDj7hYX7cyrxGdP4dM0leCPTPKBJz/ebJMhBBWg9Xzpwk3y
4j5eSSB5Q1om1uQ9V9vzr+9E/eepdcIxIxuhWV74PZnibnHZLp1R780if7i+M8qP
ssBiY6TbWyTT1rix+gSK1Eux1LPZJ61jt9ts9LOFlykUeiT1XezNWtdB1tHY0FrK
nKLME+nwvat+n4fgd1QEGkUZq+kcPAqZgr4B/rKF8Wp6AhH02LeZixz7swkhe8wd
2PCSyShYX/b+lrMtfHeBKMvtHzZhD9xnRzmAmaI9yekzkv6eJFCdJWoPBLdCAS70
vkgB067vUW+BeXD+bakjAm9jjXgaTOgqpDzpbcrjyEIa/RLq8inE4gLJegPl2NhJ
lyImy8Annz/xRFh4WJO+7LxBuoFiK7BxC4qaAHRb2HmqZC2Zk6WOkpdwHU+IDTna
i42IRl/rjlIFVQKFXMm0SG0818FvTsABtx39fq3Lc6b1YLGR1sHhY1cS+tO3zLzl
UJRRtOcAh1tDH4tJ7UuOFUyqtrgykctWHDuNUTIJIMtuuHQeW+4jRlhUlJKDL/pM
lem9yc0Rs4LKtd+QHz9xV+MLFfZT4LpU3kaNc4m0GLA9xKthB23jdAR5u6+k3yC7
n5rkoHKIuPzSw8MMafErL6Io8hzFIxGvHQHFWf0lHtdDUIDfZH/qrmz/7IAy2lCh
dp2E/p3D+mm98sAPqmC17tQHqAaKLm+IwLYcITT9TRSE4kpDSnUFDkSMI4Gv+ECe
K7RGxLYUYh7RIGsc1JfKeJxMyBTIqfwWcQ1kGXvVsEoJ5O8i6V2FqrqISpBjVEj0
yLfa4iDJt7kS49JmG8UniaD+jgUM9XJOoTrNW6Ickssn1sDyINcbM4ddCuuH5fLa
2QcyVcxOrHHV5y1bITIEjj87Ty5M6ZfPHvCGL8xXMGYh51X3suQwTVELY0MQwzqQ
GGgqAtL6asT+zoPAYr/7PA9FCRqsKuE8tuBv2qlkvXXNj4NJPGxFqseaw7p7ErID
XRecD6eeE4KYRiPeBq9YtiimQ5PB8mO/2at/DO5vVDZkJc/DsJAQmhDiabxz0C9Q
NgVuNochU9Rn06nXbbrLY4SuzTixkb6l1/f0Hjl9S+PKOw/QvA1sgdwtSPGWApTp
WZ6DJ7RyJgkY8fsW65IbKGRNh1K5a1K3cJtkBW8kSLg/Q6AndbbmmTK+Fxhbq8or
Mh3/I1Na/BLWvT731jsh4Vw07Bzq2HzmSQWR8HfhsX++XTPt1bBB3F9pbg1NOYqT
DrFYByf5htgulAxEaEC+iclV4ZEoYmRGB9MbYwxDvMJmzwE60F85rnSu1iUZxyVk
DtvwMIu58D4kpNyuIPOpzk9DAuM8qIUbHblBTYN4vsxU+y/+MxM1HfploPZ846xh
Z3+ewTDhBl8Kos8/f6Ykyhucx8ONE07n4+DoSmIFy5XSR3Q1BfO7yrnffI5xdJ0x
BtqoI0qrx+c2b0MxYPRe3mi6hrPUMHcQiDWUUp/ZO+WXlO42Sz7cevLb2aNHupEf
8vVgbsgtrogpqjB+Uy1mUtiw7kn16Si5thkp4PuQ8zGbGf8NAffJn7RjN7vOYUPu
K8Mh7SJPFwgIs+QP60OjFNZJDRviCDDt2UteWmXOTMIB+HLuMjcxMDiu0wJGsxil
XxnHms0BKc7wmOkflx5V2SLMG4kiPxq0OnEXQY0N0m8nLZsBxYyq54CqFo4deeDp
G5jdkLWQbwCuMEQrCOP4mwHrqmkW3vef6TBuzfAqd5dKkvV8B3bHX+D0LwCWj3NF
dDyaBzyJYYx1uB1qp/IghqROJdqDzMd1Jg0Ti189kX5IDGS43qCAGFE4RXk+liRU
h7l+uCQIhP8W4T7JMgcYTqM05BLlerSCTqICHWcLpxvVUA8nh+n0YV2g0ovhEVf/
fwDqyE7ejAaKrQLiTos+0zM2wfavYPktn9DtV2TIumYrRqRM0J5aZS9yOEtIS7U5
ccgWykHHWDQdEgn9cPMIkLljvsh1HUnhzFt9E7rd03933uLul5+kYObP0JKgZQXK
RGkXDy5J4d5opz7rMbcNQQmAY0aCjHeXaoQZ5uSW7j0aC8NG8IMi9Yd5nD89XDsL
7fpo4U47YV/4jw/sUW+ocA+Sh7/0jZzawL1iIedO7lxXMVuryyt88m7FA+9i3t9q
JMDDZVltnLtfYtVPMy9EzsLvRJEDv1cjIDdxfikBFjAxU/CzAOk1CG39n9aHR5tU
yZKS5fphzjIiYeuK8tIoQznQ02l3wkztV2FkNOgZ5rzibPSgxaQIBdovU8s96MRZ
h5YW5y5WrAoiX0SZookMRRlGWylcPM6/+p2qbCA+4z9BUSWMIkUr+nl9K+Ck3R8n
mARDov4FUFoJaSISY06ktGPrafxEmjPHdP8aKVwfqbrjZfiQk4oeIKjPycOe5+Os
zxplxG9gYgo2KTC5Y11tAEjAsEMNS9/MdhGKr1X9aoUVNrCn4HeKPWzrIlWh9sDS
MPk730Mecx9kBb+b6xOCnFIMx+ce9OvzZ3eAd50xU9DfmO01opwjF2LH/17f/93Q
mhjuX7bohSy2Xw+PGaotW6CKO2PfBNxrjCbnh2DAZ4TLChwhdx5pbZMGs0jpkzpq
OSIFCYd/CFA+YVA8QB4Xeaj4grYtcAbXjnqO/1m766iYOAVP6TeqTYyPtfqkpoi2
abv9mdX+l8KO467Y7lGKLOUGG1KJTdAeSW01AVdDdeLvwTDcBiNVW6V3yFFv2TYF
8rXGqqKSWp4NGH+FEWSLwqfZbVgB2zueiuLgZfIMdDO5jlJgLmvU34c/KvzWhbwN
YeZYW/bYEdsWbHb+BnDtWkDJ4IhKHEfaqXoP8tEef9XJ8bUPr8c4GYC9OZKetw/o
7vXdGUDn29nFiyTcnfS74luFhz4RtKRpPuOfON+A19RHDqoAUZftoHE6dpPKtmSo
jva242E0XAD0lwOGt/p+ehgwTdaIgLCkIc9mpK+B9k0hvGOsmRxyNmkTlK8vZdXD
QQrQIiTWAbq9YjJPhrqdT91yUbadFM84+8ofZA7XzfyGzIZRVKBjXXQf07b6U1bz
x5OOUo2UKsymcZjSL7ahTXKh0+cY/jGv07WRsG5paI3/6/HR+sW42OCdLLLfMS3Y
7onLGDFTw73VYxbdfIyiSWU84k3MvOeSv7dkc0wn6HnZBh0rZhc1rMa0QlXf7zv+
syTKVrBsbVwcLwcMFZIplLjjK4yw1c5n5Jhia03/ih0UnUrTloGj8f+9K3YFLVeI
yDp4rT9+E/Y6FkaMt7kiJNOTqyxFEziFrkjKS0ejr1NXa4F+5g5KeG5p8WLEbLtd
MMlC/TcqypbKY+RlqoGpPlIzoB4Ef6LpxnYx5Wtb4xF2ToMvpvKGcTTFkkX8++td
DoT7xjYmshVAnyg+ov2h9c6aElmKb63dtMu47fBVZEHV27oXGujBnYd8GRjGdjbM
t5YYNYSKvK1UYqMkFTZrCajQoJ+zZAzahtxX0C4Gxs7LWWHNXwMsY5E4RALnW5ie
veS+Ra+q+KsZNuF8sIZpkfA5HGAx5FzCLjcttnbGBs/js/oj8t1AmVPUmrQC2NU2
mNc0dYGpcctPMCayqCQH8N+ePiEjkwBmjt5h19dCWDKJ57c2g2WLseCLPYAwftu7
DyGWJQqgS3qSJzDBn8C0v+bZfmR64UDmAosojyQt4chWMhGK1f1Y1PPExR+BqLMd
Q6/1F0H/ldiG0VX8qTVm3jTZfzgcO1RvsYUKBWwWnsg7gDCCCCPRI3tGgDtbRC0X
ZA6y9/LgNJ3f4q6i5P5xFmbqrFTAjk+1Ers6NwVQ/+0gbuBefKCrZnZ8BT/4akaT
DtiuujIujpctEtpcsMYRY4+xkWzZ2GmVLQeyCw+VPR8koeIXFpRV5qyQGfGUlP9C
2DaB4Y4H8eAJFTn7iuYWL2Geu7dQLoOpmPsCM15XOMcRgeQmCPUii/Rdikh/u2q/
410t3gLVB+lP2A68NzEKgfZ2Dkz3of8vy9ol1H/AeG4dAIEnLE0ZjlNWpntIGCj9
GZNuVdYT3+k8Hp+YphiEyU6THK4KXiOB69SjfA13aXGwgP9BS4KH7c1YDUiiIHfD
c+Nk4QoU8uGG41lM8mpUkUeSLVbKLUZARogPOI2eidrwv4kiPixfAR8WH0JAY7Jy
WiZ7AiZJcD6EIBmzsIzQQA6+egXA7NjtaNOjwnMgIGqp9VJf47cJ8SsiuItT/5PQ
uzU7bFfu1eXxUM0YtFAweZzyrz1DIyi3Jzyl88kfM77gfSXssQwLKDtNmELGGMxU
nCHDv4hJ6luQhelhozlm63xJWFB60Kwe7dgAquiM1/lCq84XPwCMRhoR/gLzir8e
tlZl23o5DYU9oWSJ4laupvt9TiwBuCKDYp8hViLbOAgCJunpBtkMrWYIwYxRp/Ko
2QAjcrzOcwBmSUqFrWsI5rqtCDv5RjvaOTB54vPtYXzEejeoD7UCn7WQuF8TwnG2
Rgfyrw7HNtlATFAgOyjOFMWQ5bs99UrMYTXY4txOu5vxa3bOExYiFA/AgMI4dflx
rwqRNNTRASnNLDOrnbWNmFB1mwM5ejQ1xhZyemhCHhj6ZcaRh7VSniouM2ye+PdQ
zeTHHuEB1kKACZEqNgmjOOrIhdUiyGpv7PzZUBDClzWBriRRpa2TvBmO09KdjaXn
v/dvGmJCzCO0M7SrlEntyCt5WpmzQHebis43vY8cvPUArXe3LuSuUxTY+388lC2+
ocP4GWacqHLSzvfLJmqQvZbX3v3CigCx9BoU3jDcGHD2OBeF0PeRKeYG284uPgxO
dPC/rlX+uk11ukaiQZODsdY9u54Ct6MW2i2UnuHE3Cr811i+Wu4jUQA3ejE28y0V
QmS7cr+r/OeIlrgxq5lL2aU0I8XljPuX378h9u+hdfbGhHM6YXvNgii0AH0GvE69
JMWVEbWvz7jE4kFnTJt8ZQK9piNQN01xb731n1+NGOC1jTzNnRl5lGBskkFpC3d3
eCZ1KdP181IV2cfV7PLUBDXZjo4nIOtpGgzmZbBvb4dF2I022x5GIEBceCEAz77S
1X1Cpa4IDNbNtK0MSxe4uZKaT2ZCYFt6GqtQq3y0v1LuQHnU4FbScw9PoOxhvcDM
VOAn59tj4PQbZWkUnGX3PjegSznQgnOtMY5/vx/fP/Zok0S2F4LcmLJXAYQVqvsK
9VW65dM3RRrqJ3aYEHUFsFyNftVtEv4Hn3/0ZmGpIMCODUKI5zcUpuxenpuOrmtm
WRu5GrvKVv7XfIgP+b4AsEPRmJuIyUlbMpq5ZWLyd2hw5z6i5Mcm5w8I2iKlFIUv
ZBIq+6oBIQM8vYNrXM0B9pwv+niwlWNpLLfmL5uTY+xlWD2jXleckTCZ0B3osn4U
3+5Q57+4ZU1ALRnadU1JrWaFE/WcbmkjUfctmZJHs7bopj31CoaMi76bzEtqPMMw
sWFxJlacOfRkLMdXir7kphCtrnay+Kz65RCOFmQKFJguKKmFTwxtRG7deWCbHcTN
AdRdyvsvMb/2zgoZele038UoQ7tLChCFXE82e8+lvCfERKUccGItjSnqAgN9JQ1K
o5uKq1qwfnuqM6xC/NpGWgstp90GlGfl3kAwo0hxyfY2nS7cw90wZu5H4FSrz8l1
mfhmqzjqP5iE4KkS9uvhi0/OfPFQTiioPXJx8Tli0G6jtLoDIF/9O1ka/94iNVjr
+Y9WwOMV4ApOn2nN+Z1fMu/TCN0hRiTJsCrPquVNBARcKvzcHwrPfrPEAagYPG0H
qcLMPUWOUGXbnBC8mR1mM7y/qAjOu+L44lSnuMHCCrI9u2S9JzseotrIoiqma1+G
porTT41eELOt11768PZKXdk2uszu5hYM5CWDV8hIq3K8w1hk0XhNjPPFaHRdOS7I
fciSpXMxgpJQ7H2o4xZCY9EX6yCmzv7/KwHguWriksy/El39xV4mLl40bevZerrh
7FEE+dy9i/h/OV46nG/vjViCkvRtXl9J1napSt13HLlNPMNyEjOKJZoPCNSYDAF1
c50glFukQZOvTIdkmt228ofsGxFJsPeO5jzeI+unZkiLPTEPFnHuTR08Fy/unVvn
rX2SWm040ymt8BgEg5IA0Iz0wJNShfNgomS9wpczp/KSm+Gti3CSCf4JCjjjqTBd
G39sydkXQch7EJ7idvJ4yTqcPY9kk71pjMc3oNClfxStWWSetUqMGeTL4oT1IhxB
iwZM7iW8habETtVGTJm2btaXs2fJ2PdCNoKmvDNHQB+A0AvYUF25f0eRr3BTYXRO
DfdNuVdoiqkvZouGpUoRIsSptl8ckG95287F4a0s1tnfhEDvnmZ6CoEUoMrXW3dX
5k5mQ72oAtJhsT0qno0q6ED1o1sGYiKK6bwICn9hKuE6Hkp1w3HRnvxWe1UjrN1z
GHtAdPx4HkOQPjvsgfZ9AjHJupAsrqHH1Fn9u5Mb8pYPsM4TLtr3gKBaWrPD9W+1
6O7TkJb1GWswQOJ+ZjpShJLC0Azmwb2Io/aFl4D/P2R/QEQR/2pcts8s/1s62jg9
eifN4n9idi6T2gAnRDNEJK/eubFFCGfNgTPE/DoYmhL3GB9kj8XzHiVzTIDFbnnN
2wDfxVgrRzr09E3NtrISww1BSDcxynmG8O2E0L92j0eTzbvKkO/KpVWPTfFZtx4G
ULKZ7HgFl4WJ6Nn1QBXF6zb+/BEmBhbkDLk+7TQVSRF2tpour2psiuiNzkPY0/0F
NrU+h0gbpcCEjCvDAERwFzfxfn6re0IZgFv+lxSAtiS1EPrHk5qMmq1SndlDqT6m
DUNrwLJ9QrSLSYA36bueuJfwj/61xy40IXgMMPKDB5vLloH8MfLLNF0a1bhvtJ0r
MVDQt+VQW3veOJvQiY1e7RcsOeAJEUtYjL2C7AGg+mJF43Iwt+H/RkEL6aLwEYj4
nP8XYsPiZ2YiaToOQ1+QL2DsPu8CdC3nESYXxv+xaxLC2+wuFCpyNnuNGF2idfXQ
BY8t3hQd/UVYtC/HhEs0gUg2lzNPGB03uTdrDXk+oq/HHbF3uEjlXd/83ejwPEBE
ZTKlDMO7Gq+hlCMPFznzVCd5mqHHzwnWO8OtOiKyWWegHwjQOAfFdTqsqUytGyy/
POj4tS7k41zaAahRe2ZeGaEuy7QKq9Orf2fKRbeZOcgbBPOktJuJ2UdoqOxC92KH
rt9KW9lknNSpNYvSyVHpliygXTClt1dzT/D0e1hZP6Zc340gDkHXNK/X9Y/6EFf7
tB5aR3CPav9UdhxlB3qDac9uM0IQqF1LnyfGqgvGYKyA8LeKfUH4rQ8fYlAp+JCx
o5lIZeV7bGm+Dqvvy+32nyLFZlrsNwsBmqtqyP0sNUQipOQz/RKAjwPOLZO5brox
BDTxN5YQCfKYzIQ4Trhb9lwTjSbxj2NBZRGojHzUeI6Fk4gWon0CMJ1Hmqbl9lIC
m9gNITlh1WdlvH/upempD54uHegyhdQUOfND9LTTO2VPJcvAgmCVx3Bo0ZLVC8la
A8gkaEkeSh2Mv/DNu/yPWv8895hcJ8vhWSUQKcIJBHMtMEX+jRl9ftwSB5I8GEcQ
Lt272W9LOLwaz6xuAUpCtzTDfDsx4GhZ8DoSZuq2l7fsxD5YocaajZATdXiijh8u
KOdZVVI2lkts9Fj8FBBv5yOIzz6MEQX7WH7sn4h803qM/KS6cMZ1JyVLMws7oDQr
uxUsaiH3n2CeBvLoQRYSI5/x2ON9FVjSDP2W0QxJXAr0GYpL2yermWuI7vvt//YW
NVnI5MP7yCdAT06N4a2HFS4reIHcRkfCPWksOrsjSrVfBxJWmoTl9JtP+7L+Pol6
3GhFtapYlPHzKtn2qZ4VILCw4IAHA8YX0qnX5LGG2Nk3KvR4izqWgkYuLYOYNlcV
SvXFv6abIUcl9cdASK33gHaPZ59EqYIRtYsJwjXPfEjWw1wO92YQjo8kcvYgBAxN
LNJV+JnhxW3fk+z74bng3owgwwOt1bsbcg600PKtOMNOQdp/eCLB13BgENVbfhMq
lm758aK+SBXdRQriFDWXMGTY+3SkvinBm3i/xYybLEgXLM/t7igH7ya8LoxUSVNh
aHmisroSXKKsNhAtgP6XsH/gBCfi1bjzZ1idetvlv/8HItj3UDeSf4oo+CYuxwt7
oGNbl4IeXIfkGrG0bJBtB/w2jgWxrFEp5E8ShvbptstMD8kTlLfyoWiYhP7omF73
HBIopEx8gJBAB7SWQIMmTVY1PIzEB0H7bpFawV/CBdekR4n7XswyU69JqUCCKJaf
Omi/qhsvw6hKkOGVjxeeNg45mGoWV8KRELkMS8MeyVzu+WC5V1+L38+3cpfAF63r
ngj3mO9u9/bB5YURL5ofqzCsWfFvYgwuC/I4/3V7KVZFsVUnM9r/coUTCDVFEXB9
DgVpvOp6cxyuj2bc4iaUc9A3KIODgT3AvkAnBiEqUfMV9yJNCOROMUZnpGD7RA0l
seUg24ajORpUBZvul5O1O+Zq9+XhClPcMHIOwhLdL80O04/tcpHMb8+7kbxuYL7G
5aN9Az/IFLrifYafJnnVLJ1f6ftBnRYfPIE2/JcmGw1LQzcOeCunsQBrjpEm/CLb
fx5aQC7+BezmgBDbC56FhChl6evC59FcLNl4q/k2OK5Vz/ptwemkxt80BJblxH3e
GEkuw4rl0z4sk5l/abxGpI+s7veek+j2bVLasyt5nY0bwctAu45vQod5PtqwWFf0
LYxk1MBGZHPa1f/GubfS3v3gx8FN7NeJIKdZ+0vCmq2ym90n7TYg6hSc4A7ui7YG
hhCAW0yIFdrZiKm/w+GMV8fQKPZ8deGrxnSDG5PNQRaQ94q3r6a5VHpQlnKLWSoD
hxAKi+teOu/ZxzBbSOgFhGnR/i/MUFY+EGbQ+KAL/tYzA1TgzWgYHgOjk05RLuOt
K2nhpuxHa25cDTeYzo6L/s2XIikG4BBu0lljZsujbmMMo8Ud1fC8y2wiLSyBQZW4
9d2LGclUd0DImfk7rCfOtmRcGqhkvS6sZ3GoNmcO7K0dBgwtbe+vH7g1Rn/GVEer
L76JFgnpZKJMxYXCXOrfwW9zOTMAYRbzXAZQgQaPLpge2+fayZnPmA6lBhh6i9pq
EEw5ojGcPNXjIIL31nFpQskcuYrtP2DmFoKstW3vUZnt3BKWHGYDmPTDP5Rw/c5J
+KujJrFLudi7BNa9wccO8Dwm3YOL2ZoGcCR9oiz15bTPy66JGLIZheZALODB/Sbk
NrFLryazJfDXQWbiHqLmT3Y5DjNwx2jjf0V7pMAX1mrbMR8ZIhEFAbDkcSO4j5mY
28enURxF+0DOAyvUj/mFxCa2h/y9dufj7HogcF5m47T6o4O7LS1O6bStGsLiKgrD
+VT2ymbSg40MRON4jcT11BEpnXV/TVCsjssEObV/zyLDMWoSTUuF8xJYA/x9f6QU
6R7412N8zv8Io6xLFMIkbIQkcPa28raVSJH3DTsXIOSSpWBp6UVnkYv2VNKAfqke
V3HQdGz7eYs3P9iy/W7IRzO0oOGoBOn5HUYMDMtrXwO8SgRRZEOqCoUI4e6DxylT
wmgA49BiitZPDR8u3SANJs+ckkog5AQdfQd3O7nqy+KdjEzwEWS6pfSReJcEUrPn
K0y+vyPZdTmHtRcGrhzk5JnSComhAizXR5oCvwiRD0v/Skv5UhdfZQsG+ZMKadQY
R4CM/Jz/3XvBeHwvPxym48vYZf3C/IVtTHFIBocC7C7ED5x2bvyB1EQ8eA6Jsx9C
OoPxm7e13b4Ewr6Az4PCBRoSKXIKrurCZQ2/UHiwcyto0wmoAESFdBtrXxStZkIB
Jyv8Ug3TgD+rZCrqr96pYbtBcYRb0L4VGW6xpCvSaCBjuzLOY8kdSwSFVeKBKFi3
6uW/9cUrC1oYyrQ2KuTGBNHqEXa9LANsBm1K8BSEbrjuKl7Psm7R5JfCJGmsjH5h
cbxR3DqtQJpZykyuL31WeZWnaetHpf5eXeJ1V5lpgctHpR581r/HZA8dKUXFbVTa
SmeqoKJH4XPQrU6X3g7oUIRg6Nt4FIkUQ6fy8R1v9/Bm2R4RfdGetBE3kbJ4FT4V
mNMFbDEvUACetYclPiKCl29kVwWlKUMCXZgMXNwHgD8vPLLZgwmHHMXlhVeSRG5c
sjCb1Jhfc0CzJnXya49BZdEFDneHreVISYjb6X+3AxUQtn3/jgD2937F0sYpWB05
0ckcKcs0KO6sVrPYAlS1LUmyeZVBK5c06ARIkFKnfP/++Y4Q8n1rRTK3ShS+ugqh
C1L4/Qq68MNYkOlFeB2APcMAmGbi0eAC55Kdem3mk9H/er0fTZhB/YPkhE0vQo9x
g0rVFM924xCX5g7IcSg1L/kzQCpsjctxeYo+Oaw7/PxfKMLUoZ6jbmChAOC9Uvxa
bvF9IfmUzMYgs5rl9T+rd2CzAQp5o20g02MBo7SNZCyqLrl+QiMLyrs2dDtlBomq
CesoTrbf/mFOX/MFecdPg5KhoU5ebkJdmob04t9+N1rSVGmdLiC+ovfr1xuGI+dY
bykaQLY+mkxEMIF9/nlGy1dQXyN1yEmd9nRoxRuU5cGw+Gfxosx3EtSJpl71oDyV
fKhUxBepMScpj0mXAZGGxEnxa/QS37cTVnWT5Nkvm0GsaB4hfinViUBdbTgtKfku
wYA1JZGS7KycSW7TI1swS9DVK5tFd9x35ooMlnEKpV8C6q8NIfMm4hnfJZ56Dfm0
4ODjLAvnyFUjHm0Mi8ktiHBfIsLykZ6IjNCB3pmVRUEhGgqtC86E8rt7awM/70l5
ibyJ0DE9w7gA0rSBDJp6GyZIjqwDf/x9YiGcmyae8aXDN/qS/qJxBtNfN5UY2ovp
vV3j+4UU8uCzQiGL/ApNs4bpdlvNUlNVN0JJDGMkhZJkEbmIan6rqLSN/w0thz42
OI3ZbEsNf8kUvEJqk9KAceThrwmfhzTHqRlj4Qwbt2F+rbbPEHySD72Q+NPNBdyN
j9PPayVhR1GMilLQ067P6WlzdM1pf05LI3TntPslhSDdkYDXLwtMVWaq1nbFSnYn
S6pXERg39bJ2t7vO2ZJJ3Wtcy4mXAPPe3Pi0nm4orifZUYUlPO1JIbOy5O+CD56v
o1aaVRkiz7GhYr5Z3oRGoIVGcJnvHpNi4bSkRZmYIe2CvhYP+JKzcyU0EmOUJMHG
LrBpJFWxt5utgWjs599WqOcJnrtB4FKLEc/p+o/bwBjXgvk9xJHoULk9UllXY9oV
yoREWoPszf3KwhUEBRb2sL7Zo/HPWKIr+KMCWy72DuW2i7f+KhQPNDaH/Dd1ROTT
ehb5hLlFOpSBeztwnBeJwD1B0z0UYkbs7kFNVsmJV0wpBWx8NrtaP8aX362MImqR
hVFYYNvRvVhVi3PVI31WDeCPpSpnDRinh/R4yPiWz3rNOiBKO5d/CuURU3Zojnjh
vwW5SW4ctKHQGhogtdS9xCZspb9M/TNULAlbb9OGvDGxlguxkadBlXqAmQcTA18G
5qMHKT0ZSydayOktNGyhMIkELFeBScJeHkq63HiSMLV7Prod5UbJBK0aB3cPQb7D
rHXFUdDZgNv0bhFYdPaVjDsNVKXmTZD22j5tM7UUN9ADJ+otXZEfDQ0Agwk66G7j
57/Rv6JubX8YaT3qkGZz2pw7m+qfcif7lEkqdkUbR2q/mRy8ke6CqQxBvqMTVTkT
ucGE8fWEqVGgmvrzEObvjrg0L+hnIaHdatsYwCB+lmN67KDlBkxo4PG+26A8sxWZ
6Np9rpmMPjIRwIsw0G5PZFMt8uZDTUdniUyXfBt0w7R5zS2sbsadv8+hk6vTqGu4
fT2HL+DnT8UcV6B1xEMDmR4j/0gkrgZAEBHi8Nv6t+wIodNXz9lbb0DmWnZcf+J2
NvdfLOO/wijTTb3UOfN6ZXIk90xBiCehJRdzVA7MBsR61u2zR4aI9yqq7L2ixVoH
w12N+xSuR6DuvVhdX8nW+lX0yf+tL7A7ebXVYb5E0rggAGDoOXug3Cr8YAYqU+3s
to8xaYzTK4/dN48L2VWZPp9RnqsAvVNq0lgdnHPt3rSL+yBjpyaHJuc0tmvA0v1L
eVB+REKbgoPx+pUEw0iQDu2Ptld75x8uEsvaVc5MxHLU5KFv9BSsKW+sfcMR9tZP
QnQqFO3CVAa87WwNNh5gx/LuaZhBXBYknjcZdKR/kGmNnPhhs5vSU54mSC9qbkUT
T4YntVoJtsFqFjsgJVblQU0dCrSHXtJOo9MznyNSQ9+El0jWqoRzCYxb6uiNkDx+
L+uBUvuMMfIJ1jHv3HLGHIEVeeCjlvQNuKoXobnd5M/MYB3UnRNzlentPI1VINKr
ZqtPz22Zeww99Vg0xkNQOim2zzajK2myZ8ITTIC7oIxUvgl4qNiuBqX47PoHS7HH
ANlwldnjG+I7beUX3BHZlcGhi91ELww4GiG4yEFzWW7nUJhKAydMj3nBmS12X3Yx
ZjhyFOlzXWiSuUdAAKGlivTCe6uDicRyl+VR2knK3hpIGzhoVLz2Fg0AMV0pzIFz
GLjQLeKgFOcOTsxHwgeLczi8qIXcUYr6C35eJIqIAW7L3OlT0+Nbt8y13oNBCNki
NazUdxQuUBjEzFvpz3rmrOpVfBLuiGtkD84jjPfFweu8sOlRPwjXtmAC3bfMyAIT
FLPMIEExcPAx9hr+0YezPsX3iLwu8xkg/6wPILxmrQ/30CWQJad/ob+vmYjuJFAa
PAe8xHyaJGhIensciABQ8L7loX2dJIn7kKcG2sguQwqv83P7SmnORe0GWn2GZbXw
vrYbC3AZayn6XdUc+ReFIrWQauh+S13jybJjbmAHC2gbQYcygsR8ZkRtZmIvnZYa
kPfDHpI6+nMrPRkOBGfeHwfsmxyIlOEkYCQ7NAp6yS1sOtjv1raopL6pbFzDMzlI
5uVsn8ahgjCSosRD/GyQnIOSYpM9mU+8b4/irloCHPorCGHyXshlZG9hYZahISEz
gONtVOcDWmfV65TOMQeE4Y71caV9iD8PuZcpEiTr+LwK3uuBHUYdvtYfdRchX31f
65GsH1C3XxI+SnimY2ykKHOEHuoqgvE1WjVxD4KwSKn/yjN9ZrYWBdvq+4JoiX2+
yZqKnrKqJ9U6J3nN0r7Fp6wkKw2/l0H71x2PqUm3WrYN9xYrrDSlTPWHq04PN/YL
Dm8qGLOI+xwpOcovnX1JXYWLgtan6bZQneZ8tmIzI2X0ug5AEhJZyywTtpfKfgWm
Leuf5YNMGNRRprB5C99wds3JUhtAMvj4WgjwKCl/XovUaDvmPBQB+3nyaHCQeO6h
Qh5PZujb2OMZHfn9GDccBEzaOH2w+wzQ3qHsDowLGovE7iW3hOFLEnfSfXOwwg69
WUEu6ZuhS3RGMnRn5VBlFhLV48+bIPwiAu5qpOKLlq4zCorZ8j+Iz0Z8SuHTdP0S
d3ijeXifdeA3fLPqZrS3rxRAPleAUKiO5Go2h1xl3uxGs6xcjLGxX6s3SONAqND8
zLKBy2Uu8nfEXgttXu3Hh7/dLaq1/lXtwIJ6KPapPXOjxQVzayQqmFWa4z5Xxe14
NLpcXWb3LaKaRCaCExTikr8J+w53jG4X2ir4qvIPSIGbOrOJoVLR7ciGo8ain8cA
BmWBqgoHYwpwCB+Wqr1PcYiVx3A8my69Q1d+4xI3zwCsbvhx0E4I4RkNR+8l7VRF
Fs6bEmB7OP8gRwH0w57DWgpXfhRgyhkeyM5+CRMIfV2tNZ6jIlNeFPQwy0jwK/F/
bDz6rh8wub04F6VhA3De//6lPPiOmg2Rgb+g0+kDC9QTgvSzJB6FiVsvsF42xPjz
ayV9z5pWNTqXyxSllVy3vK9pOmK7m4RIVGDchJYZYTzkrj2KrW7iwCRS87WPbDHg
jC3i5p83oHR7Ha8pXh1XVs6lCVEY9poJ5SfI20uBh0AzaqOwb5bIiky+02cw7gaM
ZT4KkyWFdA63i9FY35Nl7EWGHI9oz2izQjnHKl+yIBhyVcGg8AWfjs44hJpkEfEt
wwJobYJ1GCd2OzYdkxffoW2p41daPVZQuQx4BLgEgdMTqYjf88EtH57TmRwWlGtU
NwyN47NWpxAX3tpP6xrRLEbkkYE618KC8eGXPXzUa4BpkeL8i4snYM9PMuak4RtE
RUzZ/W0/7twzSX0NA/Gj/KASzYI5Af9sfmm4d8XqGAPh6fxHeA+xYE2FfuWDIheA
gTBgE7AtAvJlBRp33PD0VHsJT5wZC38X7a1BYk30BQdfamk0ELl2QVJ4uu3q1g6y
sMXot3kzktq/alVhWrjXiojUCgT+X39FFymscsY1fr7EcfprrcvY1cXZvF7NzMjx
7Knv0+t4Q7zISCpvkAbmiUroAyQrZVK9lpH14Up0fvUREpKQIY4lIEUcPwW5cFAX
kSzqXZ6HTzKsjlrfgCuR4IAou+ilCgvVk/GeJQ3GPE43l9JeU+ReH9n5RuFT0gxP
rUXGYyBye0JtmylQkPBiVkwOyFo8ubhRQnODiCdX5vtk7gWCwGA1jT/LUjXW0ASq
l50KkZwV+8UfZdJtNCzWxl0tVaHdieCAf4XjCpXfG2mdRglmsSXv1MuAVvsLyTOl
M26+PUr9ofUflL6BSe/iwEKlBrDRuJ8/iLc3R1QJ+3hSZcqIcjnrtMtrDdbvqaJ2
I6XUBr2X68DmBNk1NYl12cpj1U1NHj63+R0ilgZj+Wrh2K94eZOWh+9BsaJ+36A7
sDwuPVTf/gWTw+2+PHXeTIlI3k3k4mTs+8CTjzn457j7yIXvP+1u5ublUJeDhxhw
HpRvFzTZ5PktHQpp7CKtQ3BpFy0MIxhvT3YBzPB73XpdwL9IWfLBrwx0k3SYdEMF
dF0h7oMoqIFwtNlu8cVdkLQKc6pNRHCV3TGnmBXAgKyVdYfgtjPVU6dzILg2Qdo0
AZWv1ORbKIgisGogqPTLR2qnB8419jzcfWFymLqauN+zSKRft8m9TnDzM3e1F2kk
OJ1QmAxvU5TRzJErStGGPis2JT7wPtg2R47zsAkYOQJIVk7cYXLtXTClPslyalBV
V3JEWh3O9Sy/58RQBJhxOlHy+bzXdCkeGbW1ZsY4hLbDyexvkkh/B1eYXoTWejUf
WS1dsHqF2RTJioMEbKrvikOBCRXJ/ALc9JAY2rV0i7I7JeRPN26YtVJ68TOn+kb/
9tZaFBpZTdvkBhd/zOIrs4F2CTw3nNHHk+9G5L0oFIH7Wmu18vyR9mty/DDs+P4Z
4kBmOSQPkx5Fgqhs2n3nr9dzMLxVMcugcb52yydCFiBTHrHMKsbgXjPGVQ+XuOwU
vaKVnwghOSvjOXNIxPbIKZBeozjgmO/R5ABxTAWmfWMFaEOVsOSOi5OvB/JZJmB8
WhXY81wxV1KVvT1zB9/1LYPbhmTUbwi0Y5o22HUK3rHPOayk1YJiSjZJaP8IX83W
PD7Yf2lOsQfiGG1ESno0yKqrqzgODEJeGuWovxzy08jL9s4lebGItwmpnUNPnVNd
lken9A/xsKKER1DXm0lZghzoVnPbXpYLmBbbYxfnou5pv5jYRs4dHSTk8Ug4OAW+
wj22sMlrnnYyfnVleyoVn+t8rpTCcNCAElw406B/yR6ADdErKY6Va8Yk8LOpGWMY
IHO81wkprdsMmxfrzZScRPstKNFw28TmHcLI595y3eImumb9tKR34ep2PLa81rp2
ThhZv6CSOYkbuNbOhAh6cg5zh3J4GAMX3XNQcxd18i150VHNaB5tZBwbZCnxvnda
ax4NZPhv5CmNeVy/9WxkPNi8hOQyQPkjyA4VTQycO1lB8Dq1U5TUdg4PyhN9UlMc
VoY19F+yTFP50PMUdRBon7lVpPWFKRBFxV0N8Vi2syOVTwdwGaA+TSBNBs9PGeBo
ogf5zqY+UQxuhM0ErNWZG3sw2oTpDAwVcD3aePnW8E1W9JZvECZ3Q+4sUWBuXMyG
H5DakRfOaZss8pXAcfyeZjXemHZn6S1LFEC7Zv4GOpHGhiY+UoiAQkaTrwV9PTft
BZpUW+rmr7+Oxbzz1NQ7al3hRTlDkMTqYDw6n/mSEGAj9aWa9LffY8gIjasG+a8J
7yuZ9A8AqottSpnoZtBP+aDdrtejyHV6PDIVZSEBW/8PZGkfhSugIoFPDtxr7hQF
`pragma protect end_protected
