// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hJmcmIEoJSzYzBydUn9TEltSt9icXl/MfSV2RSZKps7+MVcH9CbGzT7BvQfRDdPU
MRBSwIy41HIXu+rjhYL8kbNJC5vUf6I3VxVQcnmFB63SB2OdyYaC0YMJtx5Y+xJL
Ib6WF4D57id0ClTmW54+3QRtDw1yq7rvVmBdUQ3++qs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4880)
/6Of7L3RtdQno1bcVwEMMjzxsHW+g1VcrfHbIUOt1XJetLf0dN1HBcw85ntxOa16
HmIT7Inkk4+XuI2FWV2bDdYvvDJxPBb4TFJVkSa4axrYpXiprmxN+bn/UczQycDg
guKdae8h6VMnsXl4Z+voVCp2vy8EGnnNi3FoHOHsBniFwQugiRbzfnhHuyw3Hvrj
97xNgmuBh8anurrSUTVm1iAn4Hud12H8hhYGTQVI8i1iXwyjQfvePY8xHdd1qIRN
gsD+/6mu+6vtgbdgSowMGlGuv/7zvkLFVgZip1IfZgORDsEnwLp/fTL+MZuCpiCf
KXgmldBiDPbPf2YUBPpsHjY4Ra+VK0kjF8IG501UBXMaWYpfS2elnTjYnWoBM08x
xdfVTSk/AO70/kOlNVG0lijZWidlsE4GFTJAW+ECfPlkjEkw8z+wNgQRfgNKOjRd
ea/cq0V+jcc/quz2KB3w9LTle3obDNETwcILWZFoiI8c1tfAYIHyY06wpJmWx59+
yyqLBcJg0ePM6VhqyNsbKjFSfyTmukHclYv7ImIG+/dpJuwNFsGZlKfi0yc5vTD5
0qjlIdElcZaRYappliEYroyYqFgKfU5lbjQVyIjLUlhWnfFKIfZnotkdCUqZM36o
XEy0MnPBI2RWgZ4UMlyYaTDNCPmmaRUZd6X4b3I5AmMh/T0usSDk3UqO2oNh0n7l
YnwAN/FYrtP7i8QroseWim4JYE2SlJZS9ulVC3uAVs+om4pZ6ltbe1NedDCv7UHr
4QcehQsntftxzwgQ4AkKJAwzn6IE93FYno6Dwn8PBFfNfTmC+hpAQ0tQD/7wWPxk
glN79H+MkHV095h1/GVCe/8gyZY8fQc4/BAbJxbWnKu1ugaBEhHY0YH15tBX5XYN
A9w/AgBwQna4GJsmH0DuDLfja4rqcbkUyawYVxYTnaEzzlOBJR5CbPhyzd3JkERX
qVV19DN8eoH4ZBEmmtmlZMJsN+7uFpUPuCc0WcYI1cln2DB4w4uVJlWYN+ZVzh2L
+pVap6Y8qFcD1vuDJxnPJ/EE0n5Nst9tUG5coqq81/iV5VOKuDsETiHgZkwplVE2
7NnKmtl9nheDyAvq7odIRrpVSQp2B15or1fQYHVd7XXWVTNxlDL5mWL4W+WdFAXA
JqmFhhJsCJ8cKf8C4erpQ9ma+LktxFp2H7+LWxBui+8MpqPWSTpgkvtswnqx5pE4
IJaL3zj6K4tnJKFCAbqTwP2Zb3g09+hv4hbB/f/CddM4yQl70SL2gyeiOYqqA0Mn
mk9rrmCNgCLiwzZreTmpUt7DY/6CUSQGnnIsOKZgR6CKUBwjPNSTdye+g6vgG+W2
rNhgwNmpHH9hoHvlFsRtDCaZdEq5tHiCj3Ghzba8Xi0aXJ+Wm4s0v1RE1J1uSwFa
dtASm4/0zwfJ0B8mc8EibdriiYz6xGRxNsNX52/A8tX8s4NUKLTN/t3KFue0wVNo
BbLqI+ny68c3ZuVbtxPXXtEj+cuQbUwzyssCGT+v5H1HExOC6mZnr1fByNPzVx19
gWF67Rhycr9AYrnbaQtxWxL2VYTHorpOUAd8oA0yr7fKvb/cKu1cz2kQwDwP+FJk
Qw/2ENFYE7W4FJv0UQDrkWg1P43tbBZqUAHvnSPT83Gd1e9yxHQi/K+6k3YN2DL3
UlgYBA+yV893alY9XjrPN7Hk1PlSaoMcfkB3E9xI/6Nr3ifsHk4ET09HK6wFSwTa
gnlbO7b8mVRz85oJZbudSA/gm2QyuADgCGKnnSPE3KV73HnNTVjNLBk9w22iGJBC
qZO9g2PUTa7kzxHVtH80u9Xvl4KaFDy5JYzTFfIqXDO//Jrluut41x+MzVQBC3vL
hGdKprqg3eQ0zjg3bHFmD1j4hrauLy8mkVYnaug+y38MAu9HHwb/cX9bDn7L0ad9
Bp7Bic8zq0IXy7aOKDARB2i9+KDtE6AGo6Momuu3vf9Eh1RVYVpDWj5faJQSSlDB
kil7YTX3uHsFohIIbrZAiUqgdaeDnMCc5n6RNZ+hYF2hBmWVcOmiQ6uF58Z6OVTE
cA3L4WzVc+yyf2bYzmj0uDAN7l+VzwhwBifmiGpeG9UtYMC++GnH7Y6MXX1tzjGU
h6sd6cWPu6+Nf8tI2Hu/95KMRpmjQRWaBRZR+R2A5F3iXy9jJ4EKSZY/5mRwvi6V
OBwr9K60CgS7mXH2H5zzDhE8JruRZVerlUHk8sR1ZMBz/hdXx1Tayff1xeSJRkL+
klMhYMQ+zUUQqhetYaZa1y6GEpdAx4UYZuLWX2hVWBtmM7RgiCs57sunmQ5o4pi5
uCkEQZ+NLqS8HHkYrPFZfe1O1TCH5vWx85mo12ZfOW6U232GMtnf6DILeG7+S22D
AVMqD3RP4SEsKDvC4Zs4Kwf/hSQIusVVkM9l27VtZYSGtOPMosIrMahALVc1QEmP
7xhkstOp9ZJRQYLMqCJJ/H+D41h8F1X7TwJ6Op8OVVbVpsrFLYg0iiyPkbyJpvYr
NFkpu50N+VW2vTXJyrP5PamZsTMYPGBM/GAfOEesOIBy2ElkDN2SN+N+wW1cuPB1
jzRnlyRkut6jMQJ3u6h6QdmBS4TE/EMcYG++DFl1UsEB1mYZfDP9yS2+ulAp4s26
2dRueWE8wXudFf3tXGJuYC9xPj0ZC1sS9eP8VrIMY2NW3SNJDYWJampje/nDoPHh
7jGD4zD7LykU042aXKikCG+gGj9veL8bKfgW6g19FeAVMEWS0Sn1Xrq6Mvbl9dj3
tFcJ2YTZ7zAJPpdVowo5yQgU+5g6t+/F7JbyQGg/v6GuVyzGaf+6ltb4BJlaKK77
WZrY43eMm8k0+WcplICWTNk/hJZsQFoeYHk5cjIkdftRe2NMETitA8fqtGMh2mYu
v1cQcSGfBqW+NR3WCkSS31pSBaVhiXUx0TDE7bhfIxFLLlAMvtsS/WyRxpbYvtZI
Qfs+l5NzrP7bBqUDjOY0MNNwPuMwI0OkOJe0atpx5e1KtFoCiFZBc7jkxPEnhVX/
HuBC1jrULTmMsZ2Dl7ZeHByqqxIFM9Jj0U4/c2xNrcYDhe5TkKSUZ69yvsXGWVOd
EVg5MKLYoKhQtvkGXe5BR1JeZIMQAPO8MHWgvXWxh2t0mC/k2BVT0R4B6qWfNjPJ
0jehRyFYjP7+6wgt1J4g01h46hsiRs3CCVoP6RYYqTpQu9IANXL20lqqKldbBMRT
/WfFhTe8Ee4vRskB7RzRDAfzI2ID+C4LuIqgSyFzcVmRLVuryCOwSb1mmEOCrvsF
IXP3rHoTGjnjdeAIqL8MGPQwKNXS8LGYB4d/awY8sSrm0nZJcDNhOGVRU4emM3Dw
KRpoIEnd+PpvAVxBwgQnfBy/yhaw9AWvuSobt4X0AUW3d2EFW45thUvKCLqGmn6N
fO5+R0rENmwQluP4Wuy+MkIM7xSHzkotOPUQj9WOijzAUW1Wag02CfwxgTUBeZWv
towZl1kETlGCy6O/B25wgSthDrUVH2do+TWPomkHXUQH2rXhOIBsNz1QWD6uU7fb
bQXhUpaHEUslogXPZ1ERVbIzhCNx7HM9JePNzsUBE4dHkD2tMrYsx7bSO7Rx5SS1
rGI82OBarBbbjFdkU7hLZaOTbKMbBkkKfmGqda42rGqll6gJ+2EXANCP8/awAvq/
gdPkSBZwHrgKK6M1Nt4i7v/DTHvgurlwSeHOBBUdwlJ5je1t5L5aUVhDABI2kdjs
zHtDXfdlROlpbPE2fKJny9W4y0EIuwVjFdLQhmNHH/y/pJJgmt9Fo3u+Nq5rZDmq
keNCjB6LVtPGdW/nl6BZewXyZeeyeg+faoA0cb71EvPzvkNWrcnZqF7/yKo7iIw5
L/m+qRELZ4NnDm7ETjfNmtTB+h6iYjObS2egbs+I4rxeSOJXD3I1/rbZwrhaAUpY
Cmbblf6hC84sfWPbF6VrwxbyifavcS0nFcqTyEyeQP0NmtFo5JSrAN8rYoRmYjyW
WoQU4ssxFvttl5k6a00irdWqP+bZxKFzfJu0+ZmErKnshMK0FGl4ZknHNstU4/Ln
FNqbxtmlF/kGLV0vq5B0RhbB7/rHH4nAM4WTJWiATXLm2pkdne1fWHNsYwaCQgkM
KzfYhKZpOHJuEF5kgOLcJUheMqyvsBnjL7h9SeNWUti2yjQ2z/cxdrAEx4h8VMIj
IUbPuClLDMHPIahpMizCMb+qSJAXWCqIMa0L1P6FMk8bQvJHnlIlZEVTorZcoJ0u
xc7yk1VKlOnNpBVv08obfMe5oM/WDrHA/1jookF6aj7pi2Ag0VlHUfO670+XHwla
8N9/azGWkH3cspmyao+4o73ju3gyZ5crbhA+zNcyenOzCoQ5gFM5tFlVnlJPbabj
VV45NAybv1Gk4HcOEjHgAuSAmRJVIOt2UgIzyMhk9CluMGEV9wWuX6TzZnOToNuR
mjFnpK6EE4VH+GaGs0vROl8MY4DG8AUa0zBAeNXM+bblsVYg6/J4RTgajYcxVU7L
A/p8/XdSmrtVinzb57gTz5GQSn7SZoNqG+egDO56oHK+LutbcZPu0kd86LeQH/tk
9/GKAi2Gf09YXLSbpEbb+5acnzTqM09/r97qD4KvWJLdeXWoEvRvXbV2S6cp+sSN
AE6H7Ysp48NhrZyetIRZayyl1uH12y5z9xjtUAyfeRfX9JFhBhUs3NUbN3Ehvs1J
cCmrkspvJNJaEQBR8PO39710JVW+6vq2Yv83WnDBp663n1HehgGLheGdqXt1osZs
XrXyqUNLTGT1JtDsKIsJiu7QYu0LsshXDVa+GI9jR0ywb5BsaBQSNrYXBhbTHS7W
JcUDpj97kJmTYwM5JFLHokGB4jYRuEKTN+o8tWFKFe/L/mPr46jtLxCT8dim/R/7
fyAIz8V3S/TMPB9rWdvq2/0ESkV0/qaCCwlz4D2rObA2JTGd0UkSpC+pSfN/i+nO
kat3R0XaZLCHDi8gt7H5iFIMTP2aFQTrAQvuOEhDvtKZi4vMj1zQYzCa4YufUte3
RkRgKnp7/VWNcm7ssHHiGrs54rb4meMtOBbq2jBLcCFpT+GM5soaLjGfc62iYw3h
RTJwD4zpyz5ejhufxh+j+ggPfs/TEz2cWxMKAH+xG/nHwtDS7K0QDThNqU2nJjDA
ltnDXuYM6qY/LoeZqgCy6bei23zjvnXyCkHajp5qaJuZrLQ6JwaCjhzLAopwmNtz
+Cr5UnAQWSZe6oLZ+DbvI8sw6Lu2S71KFAagLDMu4nPchGyjRNWH4woEtQQRldc2
nqbmtbc1lAEMK55zVCm3tlNe2yK8nefd9Rn3pKigWSJmtEznt4UJxXHnLrrZTS7+
1R8W35NY+6i18gUTTtDpYDzcJ+JjltzjAJ43O3/JO3hb4mJMeh+CTONM+/bpYz4K
b2wUTMJY2W1xk5kGcKSt+iSs6gPfBYYUpahjSphS9CNpYmZsUdwcjA53BHwLj+KL
GJrQDSMyLTLaoCFErc7tn9wEL3FPpKMHedkT7meMIgI9dJL0+wti05bzCcSVHz6I
vIFwT8QodMakEUWoFEWDQgeXaWEB9Q1wlPzKlKQ25RH2DlloLcoP8QGR0bHY0oIl
8QkCNY/+SMtweKdIQoaYolW9350zl1iXWp6PjmwUhp3XTPu9clOqns5FSy4Dyz2S
PAo5TkEBUXEMim58BE18ZmqMCFcgALr/9XXX5+CmHBad1VC0sHzOHLHWuIadc2VU
w3RZC5aLx2HkkOEQBTa2LeH3jk9Z+IZ/pVerItVUwZTMIZxVVGt3aWYNx80NKUDK
aGep2pUB7sLebjmhiHQl4p7y8RSEL7+OdxsT/L+93VRVWrrupR1X/LlnT+cQvBMd
F0q3wA7yKUe5BrZRwRRbM65NgzaWqXSdOqGusMNfwOKsKaLvEcAEjee9diGLchtP
JStoWqVJ5TwrQpEMF3hnSGw5UR0CRKFmTKo7MAVg9Bw5k5AAo+msi22g+uKKrqIj
ccY5gUHDJoXPUMINKJBzKHiEFZTeB9w7ydG57ezMo6m2uOep94faCkjGZwJbmRLd
ykjDrRLMg66JuPnvGSfOnPdPb23uM56p7o/Uq2vK+EVWAt0pcZYwSqTIsBb+vJwx
9QWa7DIWQBCpby95bwQ7ahJ7lIpZU60Tk2eCe6hPYa4IiAGVcL1tYPp2bRxquRsf
1ZyiCRNkZFi+Bk5zYpJP7fReAblsmSmjuwQ1PeuxRkLudWL2y+Rtv2lxDhZjXOHu
0Hil85/fnjI9tRjWI+VyoJAtE1GbmJjrSugCETb/i405C5yD3ZbxjiyxMGI7ympv
BQ+4Fb4bnTVwQpBZJVx+WlWjRZRd0Lor0BlB1EkLFpnZAT2Vv6tU/04tetWckJkn
MKUDUp9kFA61MUIrZMcYDuTbpnnI4GUmmMzQLleFpFlzx+DreKEh7FijpKj+eWwP
eQ3IbSgIp9HiOAvLxidS265/R5UaFgAFIBgRbwZV8kSaj9WAT4ItuPw3QWAcJVUI
gXdwum04loY1AlNNL5miHzFLuw4xOgQ8ChEshEBF9zs=
`pragma protect end_protected
