// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e+qNfmIzDJQs1EECihWMCa6oq3YGFUxfxM/BuCHVvJXUjxGstjQS5wP76S8Czm3+
PoKavnM03vi4xgCwQRjN39/pBlSLZcFcqYVkad3ntlLPSRceGrXkNLAPJmeLSFUC
3ItiZWt+GJ5ey7QBaUiWnTTpayLwYDxFF7666/P8qbk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31312)
JVh7rGfaIBRCYFrTFDerQ9UL+l0jo+e4Vd2YajKdMZEoivkov2gpkxrhcb0lVvN3
txT4UlynLRibQdI57DDdz565UKAVPh3w4/APDlAbmyTNGbh2nRGNaGp2LhmpNbXQ
5KbGuaNsbUFzdX97C3WF1tnAXRqMMayCNUtmWmb1WnXbINi+W7TlQeXnzX7S9uoF
5CwKZOj6xfkBMIzL+m5slaOu9o5KwA8vBdLzoonirSvdscNbV4v6ypkrJSti2x9f
gRtId4IWusLsWO/g8YuanvP1pQY0wFqDZxfAkO4McW7ggxVxY7vJdQ9yZj1b1GT1
Tnze9lZ7mmcdvAf2CG+yauJi1Yvs9R/0q3TcAoPr8Big90Cs+VqhNXnPBA0n9yg1
crZB/wEzrQjRzoQ/OFH30gK2XACbG82CbJoSCWxHB24RDyCTKnTFZ9VOZ0IUDDlo
71iTlGLzTqaXfg6vqbARhfqKNARUbLDZoVb1ATdEOtBZKDrIuJ8SqUCCMBo0CAiW
Ntu0vJUuIZVAGn6GENFrI3ga8coyNBFAvAaZNgC4SG41KESg5TC04A5+3K/94DHV
Sq2RsVFBF42qgvrKMuJQZLyjFlbI45CidvUExkS2/n8maZeLFRISPO0A4GeLpgcr
VTejQSGMAnLRGqaZ5KXp9jnC+uTaDcL8jcyvZMKdxayjJF0tOIgc5Sx86iP0hgQa
eQN/8aN2kIdcmqApTK4OaMS8MQlXGrOqJnCCcWY3NMAshTAu7Yu75PlqywEZytlJ
m58ZM7n+oFeSGAIh3ic/FyYeDUopAojh6ZAtLMvq6PD4bKLKdEsW4jPnPMsDd65d
X7OYNH7lx94I02m2YlFN2QSW2BEciM6fiiIZQC56R5VnfPsJLtJIMH+CWsaia4Sd
TXiT0jepYExAS6Zf9vBh2MhxVv1OqwlzAhl1IHpCX9pSlnsNN8mZXii/qoQQKjmW
hxx3i2MJePEb7bhZNFdSF77kQyuKL1p4hMCeWh2vjWSMWO8CdHrobct2r7VmOStY
bcTKlSKbH+RuZB6Hcc0jFNiWiM4SY+lG+iZI4fhxSphtcT3GgKvSp+nlkJzWWMFh
Yj8Nne6exjb4gf8nmFVV/rNSHjQgtsfgDN/mQAJoVwIsOeRVv+/iIJB/hXOc5gcP
cjsO7DzFHVreLyZfu0E4LGXlNOpbd6iXRnhdsgdtcmpgTAN+X0naVGZlCKExdv77
BuRTWn2amFE7JvKXTBaK5UUaAKbLuwieXcyUHcCTan2LVhykGRDASvxD1RIqWZS1
gd2oVRv0nyRidmEURwjKHyq9FD9tQ4j4HUQzPMTTwhtIwCD3qJhP+VDhjhp2V/ba
Y+xO7fsOpukbeCDlQ79q4SN83M6Ye7gVqFV4ol4OhApFTUbnjtbMoJAavm5alCfe
LwdruzKAyG6KD6sFRxGuL+9+OYK9NU3TyU5bi/eIAP0OGtYAunFlp9KRimRzf5JR
bqbBP0pLWLq2Clpfg2T7oBspbmPy7YYfqPR9OJhsm+Hv6cJA2bcKqNSjCRJ994jN
JD/Xat6s0+3c7lhdN+09XuAqwkjulo2jXGaK9QsCcpuBe3bmLkmJNFFD15i83UgS
JXb+hL5YWrUWnnGUSQcZPrazWLbl8PTc1r01IZ6l0CTShHsbb83CCY1xy+efeKiM
FF7LmDifUAFUzhTMnAxWxPAzqZ28TSj0R1bJQq+Jxa4Ae974D6DpZ1Elub+yc5Aw
70r9tKMiJ1cXJqdg6POVEwC7eeU5YGD1GqNNUQjRdjhtKVH6U00Df14wWlbMTgjp
NnzE7yWQ4szn+IDPNrw7kyasjTa0JT7m6eJbwN0/Zh5paO7zWTOAvL8RNN/JrkhG
DDhDULF82a2XOBfwq1jgObg72hW409SyWH/v7CMAepYdi33rMfg7NCb/d9VoCyMZ
B8iorp6w5zvlG2am91POpctiYiWmvD8s01xeb5+jNxfDJEv4ED1VFq5xoeGvUPvd
Uf3ETSOZj5fn/KsBK17+JD6JH5p3xcOb47DGj80tHVb+/wvKBXT+QLTwHI5XlJeZ
PpzpfcBPo0HaEnk3mePoRQ556WEnFjQeTGm4KgxayaR8rJy6tG63IDNwnvjCgKwa
I6/hGpXsWpcoCrXlNWzSUhUg6XHSI3NKDVwerAbG1OIIiHI5PoreU4oqMgmGM7rj
p/19WI7EBqrACjCfPVMoWIzNDCqWCq8NvoKqAZ7NwkvQr/DZXiRpjEiyaKcAWznQ
gNd2pCzan0nvo86QfMyW1sHOgQE6JNDq9I6y/pNDUPDzUkOq/OVnw2tejm4GCgiW
QQbIx5QlvvgkMxXy3GihTD3kCX6q6+PAmo0Gfu+7S57g98YtpHbzdRB+LdHXn0Jf
VoNxHiFal+k7mAJitKw5GiMJiPL7GhJ1EzyLqifLvahpEsDZBM5EAuePqh38MRGO
iR5xFQTc283l4YARqzeHyI0nEjxNBk2IBR/d8ZF4GZWkM5dIDQiBdpwctEWdZyqt
mkW7lQLDfTgZJbX3JYDDDjhrcli/pMoSUTQogytW/gFCdtFvcfTudTPuT7zoUk78
SHcyZWWDsAIyo6yZku4XaVlnUcLNRMRCXTM1nsP0NKH/Px1K83qDeodlgaKUv6/0
qTtMoGWR3wHc0Opn8+7NFq2hVAnJRlw8Ks7SVGePof5ZJEGtU1u80hjl4UbzZOH0
W53Tcp7enjFFi5ERfuJVVgGCotO4MlJwGC7yDf+CF1NVpL0ALzsYQ4LD+DZkv1XI
YJ7fdpu0vRFYAMbMu+p3hzdU936RWr3GWZlDEVN47DO0TGPgiSsUNNpP6ZXNIvr6
/aeJ31OkyImsIgxqji9Zq1RphdbbM6CCX9JAbxrvxQoV/hnkQVbJuuZWnmjwVRd9
HaLln/oyFZA4kM1TH3ZdzU//hEM81rHNYx7U431GdrXkLrjRlORRIB9Fik2aY0kr
fZbVTbN9CAQpGFPB9rBPoBIX5KTcOcHbTNoearX0xiOqaWp2XZG4qJtzf69GdzB1
ebVkiCCChLQhPZmgxcpJzIP91Pvwknb3TxHz/YWphYkcT7Ww7NPQCRZBoOxNUUdD
1MzgXoUEQCEIevh9OEBuy+PAo8YY0iarY5AtxSFA6mdMcacGSZy6ZJrJ5BSPL+s2
2a8dQ4CAq6oNRcseYD5dgXIZwTA4Cl15cJBVFQmF2qucDHPyahpj1na6nCvOXzGy
bo0l985kIfMc49qvY/ux6/UPO0TYT5tyxGox+N/fHV/0HlLOmT23YqByKSLrqdyC
YvkEe5nJINFKWYlDFZhKPQG19WZ+UF2xLTgl0yCdEULP+FnCTyKSN5JGitnTs0vi
j71Ux18zC7hShTQUnXlCGt3YfvFFSw7lG2NPYZQRz34WYoJ5cQnc+CsOjfOgyoCN
9PE8v2/ltVKGfuPTZd9aS3bw+iHInDPt6fdKcSGu2kvd7QCjuvvkgMxApC8bMxHQ
0IZMFLEIByFr+r43kAs6uQOIgpNGYZ/MMsH02e6rR6tgG8JbFDkAGbzW/kry56ds
RMCwkQ0mSgxhUJmC0tA8q6KaG5groaE/yAcI1kCg1d20jP33ftRO//oLZK0x1LW/
VOFHpH9HfBabU6urkhwoAC9w3fZjWx/aXKot3gqAinP3PSqalpVChX//E8hmf/yP
rn5EpcwdAH8Vtk4icHZDAJn2XXprmtMqmOiECG0aXhnq+1GjL/KioluQqdrZqzit
8sssjxwaY/BzE6V9R5e+Tw7Dm9J5bB1UgRHL0xiF1tGv8RB2DHXtxLl5B9cMhOmB
JF/a3nIzZcZVJ2zn6uCvjbdhJYnwALatiIwTNj4NwSYIr1JxhwzsR9GVHp14CfXr
QYdapGx50NqVDOCcxinUdjjOyMZVPovdOX8PsL08rXXZHZs22oum6wTYI6n7CeRo
PCdCexwRVZn2oFfKEHw8eM/phO5B7Qc4BIiH36BiH888Ou13ioa6qXyZV/Pv5HYF
pxM2KDjJXsFHLYvCysdehVcqpkN4r+8J+lRVc6A7yer+9vaFBikjXmjrZzBRczcy
zMcKOkuRyOzRkhvzOSShYSUPVlF2NpETWB72VD9sR62JgJVEbXUSRoJuiXsjSG2H
V2U3qdKtAMbH/p1P+0/G8Q+Pmd07VOVz1poTp5+FhU8sbxmRjm328RbZ5402hBNn
+Y/NvCeV8LjMrhtvmnQg30GMiLoHMWGLV+5SjA2Z7mD1gGk/uonTTGCTUZCNmJB4
OInpWRWLLthvIeY77EM93xgezGkxjhL16p4AtNu7urExNzyRtguwcif7GT6V3z8J
lFkmaV2nvuVF9rtUvzlJZ+NHgn3btgFNeOENU2vCLiALaka9PJ8CCkbiApuFVCH0
dHmqjt1u+VCNoAZ7f6KgtwIlhGTHcVtysR+ICG1RhGKvJ7MNqM5PVeVLQsp/pe6o
hkpHrTS1WlIVo2UJaLAj/HVenTTCrto5DgaS6jXZCajsca9G1xPI54dNtb9Hucbn
3HCZgK9FHBTNdc6v573pkJfN/yDw3scudm1vkAfpVNHbDkXnv5YI1Xn8rd0plG7N
0isJfdgUrxz4AM5ReKN+WoNvpZiZZ5roxjsoHCchCdeGzcNWQCXsdpCkoEbos4RU
I5TfohDjnySMPZudAT0fj0lapPDMUfIQ98142S+LpSNTIW4zVGJmG2EAgfxfUACJ
2CE1mfImL6l7/6LbEmQq/QHymy5Dogril/72xZG7zx47wD7b3GCI/6KjybgpgePe
tGAa0OA+N1STQI4MPz15HcxWHw0c1Pi9osYVLOybVf/et39hNUV4OswR07oLvuZ+
NMfSBI2Es7j0b4vEqfRdipxm1R9pRg9ZmeDn3mWtQQi2A/LWK34KKva29OasgUcQ
Pa+fqqtTo6QTQFHfyjMNZhxg09v6CvzPVZBNYUuARx4oqedefYut+hSC5Nb4zqS0
Uq5XTiG2bhHzx29nZAqcPK+q7FpLJhriVhbf7adi/z8FCMAfJYu/SnNLkYU6hQVf
sn9pv1l39Y4KEMe/CHnOeewTWZS7FtdPpIhBnyHyiBsSoG70Glz6qCTSblVR0CGJ
OwHN2WjoIxLFASdZ9vKPjMQ/cvzlJJ8unDqH73vK21Rzr68vEIYlV4csAeSWxuF4
3gNuAGej9RdY2VUhX4JT3qnvUDXt8DEOHxAdz84YPyZjkzFp3FwbLZ5m/Sh2aVjM
DKAzgbGxq7gCfyqqRWzEbYSUc7Ohyf4gNuGZsYF9aGuAT4WEKO+vmBooKEKezvCn
SmlRsfmIIRnoxynnNVnKKl3tdze1BdMB5TTm8ZfaOy+L1rSLyLN8C144qL3X5c0C
KPWlbyKtiI7lljlx/xtIJiasmLfBBHtmWy/2boPJZ8LI53KdIy3yTSQbgp9Er8/2
9Oo6TkVI7JIrw/JfJ/t4vBDrgRtREO4SYMDMhE6sckgms9EJnQ1Ycx3ZuwLGPRWC
lgM6INq5SmxBPlohk/+pEiaqPuokY2SHPjlC/p6sbfv1XumnuuNPXB7sgnYzYnns
91OHCeX6YznDyGfHlbN6nn8plF6A7hFWMGW03AIKW6sQo61wGgFK8q7TOO4WreOD
EODSBMBGv453+Xi12TF0EAJQvf2IolJODR9DecG7NgoxeQFEpe26/7jE/fixAKUk
AhxHt1q6rnv/ZYGRaHB7JYZfExr38EmLlyPrzxZRn1c/Awtm/GKuDvCI/LDMYG9B
yyCaa0/F5pKdAXT7hKgYciFSMF28AZpJHug4hG+avhxbiiPSpJUwlPINA4OFOscl
olkaxM03+GEYWinrXJKCVBHi+W5f6IOKp8hdNJAChHRftENsOnvIQ9HtDko+decM
7l7nRW1brs+5XaI8XBbRPmill/YTgGmw8H2W8nu/cyOa0z09DUGworUUWcWQwbrA
nxE8BIz8FnJ0rUZKH7xogJifUKcYLLfrFgepXcCokkh4jBd/5pyxfKoAXDmb+l6s
ElfOWFHHZ1hoMnHR7hbJPSP8CRWxHlq5KHupxv9XrZVZs+8fpgf+H/4LsNEibQWG
3/wvjzhSBIAqxSCUu1YPRgyjRxXMNq+7QaXprtjVeznl7Q432nREb7HVv50iIQNB
dxkfgfuqx1AOy7WuNze/ipij9wKp9SmZIMl01nCp5eEdc2Vjr5D6n36Gg53Rfaw7
V6ENYVx/3ytz9h092Y3BIspk9FbruEf0W45dg18FoSNxrYE+JpuIFxCexbjqWoKE
Z6Bhr23/8MgSVD7ekH8iIg+txiughsTImpDYhGQ1QCt4+ArYkCIs86MZqiQA+8+K
Lb3r1Y+zRvbLhIwvbJ14Y7kL6ENMHmTaAAnbgRVCAvOoyQvM3Z9az4kJu/Bq9ktu
EN73vdDYc4hBHPV8C8hPCa7Z92cRtX4P8YRZM31HVxmK+3S07noZylqez5MshnJi
IPeRNLjBQ+9JQmIeMvcXt4FWfJGMpT43P/5iSJciuMAPboasN/IqP023jpyDuHGe
llx8vTAd/wQMxIkO6i4rvSZ9EzlZsabTxwQfIMjGCdeSiV3tSVAj0RXIL3EZd9s/
Q1v3hRu7gMmR11qmHd4j9ZfZ/svXJeY4sX/863TqGDVy2jY9cdQIDLEtmcZedN+9
FwCxKu+QhhUbTKSZuFUdH3l+9euYN2P6vANjLJB+zq54XKmMpOnH3wXS83F1YLKk
Bdfo5rP9RxCLurdr5taVgsx026iC4RwLGyzDogRUrFJXrFj0eK2cr1bfuP5hbKqj
qyVOntITYNt7QLie3KPA9sW+iF2xpQ2gUDt5+17ecpgnl+TAhgYVrouydzBow05v
Rt+w3kuxv6Wuz1cToUTWzhkSqnzYpOiUayJpDNXsge1MjsynJD2fzWhEN83APJwV
tVeFRqUI9UZp8sO0GJUPdf+uhK5iPS1SaPrKHIhbLxUKXoMrLjxx6L/1XxLiz3yq
R7uwIIdvnqem5rY2S7yGztD2/1CFDVRvrg999ZxES7uaKUoraUkVZaK7jlpkXKuT
f8w5DMZk2GLaE8YHGh9sjgPzIe+xP2FFKt0JJSLx/Mob5o6ZJ9vBShrPhrjdR34u
YN25PORNatVBPxwJpjCOCHhL9CtUu4ovJ+DZWkAzD76wTl7hqVCD+uN5UOZfqTAW
bFPpTFemQ7NGZ19bkzMqgpdEtbUzuBX2eykr1lGCbozbr3rHqTCzUYfT5sgNjb8C
lKWXF6MUjhyKg264VuqThsS5Ah26WPrI5gHDL0Lm5axUd/qN1iIlAu0/CGrb5UUt
iZ3Fu8DEofFRWczGv6lRPHABJNoADOmeiywCMxub1FHVkz5AZeN873teSFrN1Don
TQnLVfovtWpgDi5QBOdajHbCAbx7OHeBBZr+lObDkAxywrZDvCEl1Bc2dQwVBTfs
fy+Hc5URMNDz4oFi8c2L7a3pSD6trAROzT2R8k7Tbew0uU8QLpp966QapZCYxfAn
AHrV47yl5A+ypWJVpFA0oa+SW6g+LQeoTiiTL9QJLvZPSEReC9XvV4oGWmsNOBJL
/QWGiScmx0l3Luo3iqLKT95ST1NLzItGYW8PziZEHrOuYiMBOrH+vJTIZRrMl/gm
+KFC7VeleVxrZlWN/4twAqCgPFSQWqxY/VjIVjNYHd44CuRPQJI/U0kKOqhYzl3x
SoMgFlhLUhd9bbpLA8Yo+pxi79qjjM9W19IvHBMBoFcncaKuvZfwbaU3xviGze5x
zxRB+ltH5Vob3arSK6GcfDYZZ3y3pbWW4XFVFoomJOP66FhPAbZAYyZiIuO1WQ84
lE6u0Rgns6ZPacleZ7hrNiywRLuY32ulD9T0pBE3Umw9Z8ncfwBfmG6RZmKeQ3Xy
/nYzQnGLC4F4n1nnHKaWmLDVuYVe7v9yOPaeP+A6vDbYnUKd3ttDGKTjqoD6tEil
hwPgxzmay2i7vO4jO9zr1dGEGrkuAwutiZW8G9LfpySDCV9rGgEIIUqHjpk0neTT
lTzHifJB7GLp+Y4ye2PyEdejNn4QxGLAqT+oNCKWOqxGNcl2SmQQ4QDj3G7To+rX
69cSEg6cdgwAEIxaLc+PFhLiT/1JQoATtLKTqb9BxhTmDhjRMWSdkIekuMtsJqBx
jAFSP2mFcCd+wDCW+4X/OJQphoepjmRikxJJlZFoQpnzNRfz573+9w0R2a2MuQlV
jpBSwJ5Kdd4wownjq+04qlPUZxPUsjaNndjenrmc9qVFyQXpqSIzmpKlCWm0+kO6
Ojm421GDiM6jr/nHF0bZrnXpvn4oay737YlMUkwDSzEeuX9+QyawuFs5+IF9CP0R
Jjx09BrSJE/HZ9+HtrtcnLBcE5n+F9rKKe9fH03Dd6Oi77St0rqV36wDY6br52W3
MRYzIQ+RnaLmvK5A5F+owOxGgDIb3iu3FFUSLvpMZKoXGSZSWvitwiQ5wtqjJGNW
5t1tw1Lo5tqGJEuZqusQ0546gRD+wE/EU61FBfLBLWs1KGJE8tNem07JV+vx7LFR
AhIK88ZvFxRSSGGulfH++I9b7MhvCi3VchN7kK6xt6Z/COXaJ7+BSGR0+Ox83dfZ
vZnOtJhOXcfglYfQDM3/gQn1+8Nq3WsopoiiIfm7nzO3VbIcCAoWhxPFW54Jg04Q
YGh73Msy95A4xNaVzsTFo8A/aa+6oaBvqhpY0n/VW3pK4kznQ4vc06I1w3LEuZw9
fmfOGe9wgWAwZjrIBPjUcCUOisxifnIzSDu/GHYF6GpP2RaKI6luyWgy9Jmuu0wO
MQQwMwYZKJvZZaD4NfPE2M2R87gmbt0u1dlD0yyJktrjIMsUzkiGn/LAgcxI8zhE
XTlNwssDBbT9JlIn1fnCHgdnobn5D//qY8D+cNXj9wpAygNQGczgUUjeyApfDIE2
6c34y795BmjGYM9hMOM7J10uO3kQkOB2uSyXZ+rNOx1Qu65p7UI0c89VNiTz4Vnc
emDhpLBIPlie66xvFqPBCCYn2LT7Xu4wio117f218ZaGb5zuKZQb7AaoDhm4es25
Tv+kNk8+AcV/NMrwZYEV2UbUuJMHasALex6WBOEGVA9V7KHp/WM+8R0GThRfJf/8
fEnM9cHv0FdUdj4deYpXOM25BKK55Tquqs6VhpxrDR2OM0B5lQVE4X1egL9/Nrcq
pCMqqH93lVo1LHiugqnW3n0bciXS9Z4CkDXFA7nJp+HAhxl6540r4nZu+nEjmC3X
quu8gB/vJ69KANgiqKQJTFvl4WIh54+fudzwwG4XbM8xfidjIm9KJKpw7/+i1Bs9
zlq4zAu+fUZqW2lMuDXhFnRuCyFqZtqUXjeyaaHjRo7DIlnnPNFMKHX3lyArixe+
0l6HnWEgPoyFcRNV0q1M/FIhc0OqslmoLboP6//H49IkT74ciGDlA1yf2lFCTUue
TCaDsWgEVmZzIEUVG7e18TpoHQf66y40m07NJeS1IftN+qTw6/bFsNTsC/cVVVXg
R15OnTHXn84GBb5ir0F4+lI3kx1Dn072daHRNkilW0qfOuBkUFQlFrVU4+b9wf6m
nMiuTneT1IaIBsTb1ztTjA4cQMgX+Q2sWv/dIVKKg6cncHOZz2oMD5ediXmb7Vt5
iF3RT1X3xauq9Q0mDQNhu+MAG7jWt2les5LfUVQMGgLxAJc41iDYAJgqQQyP0/S1
Iaim754FMNVOw6oCRWcGJjdJHf3979vkll9pItv2W2t/cS5+OX4tzNO5IbbO0kLY
CfdVvrPKK0iAkHpYLaLpVXAYQoqZS2Ec3pw+DJBsruCz4RGWYmh1NkZIoHeess4M
aK4CN79nvlyI5H2uKx6OasoGXXjxzop++9mJKNGbKQN0+e2pzR1rUoWpOhnzLlTb
+HqHQySSS+cP7hLXOvPH1yd4kRuu/vbqMo58TpF/CNFiHxc1PM3DjrWRP2I1bQam
lvkP+R4CBCmYL1ZAsCrXXGNz2yTdjykgrIZuGhsYsIIhyCbzOUjnDKA/k6HnXBWc
PVa85NMMrFdSpjwHGy9AGqpvpTvHk8f+dD/nxy6CacTI1bm6ZqnS/Vg3azc3Yo/J
9XkW68pj6p+qzF+Ct94abXfbzbBp+p0d3GRoV5OrBrs2ANnykSN6lIkDosye/2s0
8qdRlxuwZg0XcA6AnwkaQcLCy5X2GbJjVuJZ7G08vZLE99P1P0heDjIK68NqLjpe
XshhggUsmmtf6hjamucQzJ8rkTTXFulZ6CtHhxz9ea5lpO+B3ADNXbEvtckeTGax
Uao+AnK0+AI9tt1fwRDpqXOnfyYSkqVFqhg85H9Q2u1EK1tKPaQNr6nlszmNvEku
pxtrjMwWXChl//Jij1qDy/Llcq7yrPA+mfT8urfZATSpFavBl7aLi6SuIj7CnYRf
uVTPXNSsHcO4tXx+xeCm9eW0/iPmo5R2smeLxR7xDeIvn3W1S0VHI2no/BpW7s7q
1UBU7DPJ9sPKDHFs9M0JXSs3s7D2mwt40auARqY21bfLModPeJNgvmtJzdsxzuRs
kZJ/hEOFs4TwuGLgJnwbRJIs9YL1oRGr+xLpyTZhQR0tL+wE5LknC4AYLHQK1bAR
L5jcX4XuS9Eeh9w+W4+S88G0499mVLUkN7oEhXjRKEPTFsG0Is1Py82r+kydWE42
fqH5Y0RDm55yQvcmZqPxIHJYzahztY5HwPth4Uq9yW41yvBWdUji9azq/7n1/25m
G1ASaUuByuQnzIfyCAYU2PDqsxaren97gsucBFzxi/BFx36hDDWfoO+eE3bPQCKG
rqVqnWAQaJu6TDy7tVvBPeRXFwof0dfDNmajc5ZuJEL7VAeCBaqHxfYUexY6aevB
ikY51ehCGtwueLP1Q6BLkxAxcLqzRAKSzu/H9vGJGcwjVtkllm6Yvf8ymNJK4Y8W
MKowxk4FVYVwTQ2yDPsBWiOYPB3ZAciMt160NJUhu/fDlTAKDng73tFe6BfowbVi
pVU86EVo49NtWuLzl3gfX4RF4kiTJhfD9rwUFF5p46cQdpPpABu15F8tJybWJmys
LzYM1lko90Z02CxcPMfdqZ/uP6jv50MA3POwJhPQAmBd6keoY1kTDylc2O4Iuzp3
8d5+BFo5M7cMnrf8FHCPYO5Rbl8+kyUgZQHL6JODfna9Y3YsHGfeqq4wnWfnw2aP
fBq6omPvgel0VVi+M/pHsd+ztOCIeb+Nvd4ZJcwfK7htNRr7fvTVULjNLacMUZtk
KfoymZZAr2XLbkdNQT3ckWj8rjAR7s6mOXMJDw6VdJcRqcJaQCqCi408gREe7Ez5
JOre9dPPu10urhIDSPxp6ERLeqQsPv0C+BNG7Y4xb6s2CNk66IOP6Pzm0h3U52vb
nBnNP84GalOXVxQSBm/eAf9kuToy3hAc0fn1DRO7fl6IY2ERE6LJmBpM8W3+Yig3
StLrD5FFhAhF4qrQEWIr9mGDQV6wBNIUJxrS/29+eFZIVjtTX0H3p2b1kevZfju2
G46RtnPQz2Sm2nP5r85yq9IKKda19yccUT9+OFukv/jh/WaQIxGIKtUdIvWHt9cZ
Fm05fJwfHub0umYDVqF78CQqWPYAw3Ncfm2bTgalrrEktW8F/V/Xg7IS2Iu805MZ
WGZpGwOAAYiqwlS3K3R1r2frCnniyp3YBuzXq8qh9TiHIgfRdn+MfPQ3yhEeQKfB
mWMKl9YxogbPwAXDLBpSaKx7htDkYkG8Y0HqqjUrpAjXcnqdYeMvke3Z279ty7YN
iUjCAiP/nEYjJnxuNQCsZnd+jkBlGTMdN1p/WyHVaXkQzv19OBTrzU7ytepQ72gd
/5MTFnt4ZKOWi/oYdo3qx52n5jwHuzZeHsiKdLWLr0h1Y6i/xHfcN9Dkqvs67rcC
T1VwGUNPrfCG3zYZJL6PKPHM75ed02U8vENfGGTWs2ZNA74FGEgmKJWshjmdi2K+
hATrlF2iwT03AIwhbMexxKVYWbFn3vHm1cMQPcaRHmexFU4yqig0Mq/FCFfjt722
1u3LNfPoXAgGNLKWGg21OscfLnWauAJIRvGjiDJbZAopfPuxxAt0zsNzgaylD3Fk
O195TJLgZ8zlP5E9Cy0G2JzDJeyC7iLnvZRnx+Dml2+aatnu/wsCHJhZmCVroEaQ
nCsiofa1JVmFfyIDKEyl+Mzxm4n6teduMGBy5/xtxzI9E/ClDGREB2MLCknDmie8
llaE3hNr1gpw6Hl0AoAR652psoc/TxZEQuf3KVdrqm2LT0O61SQ9tAj709NTl0q4
UklWNP+UHuliFnzLCiQjC92G9OAUbM+UzZV1j5ssPhvPS0eOE42TPhdRwNgkMBRa
DmhyPdDrPb4rWYVhOgBI93U1OO9v39HUDYPZSYL/zcE3RI2zZAEOnfnEmMph71k4
EokxkrYAKb4fp7jPTQan746TO4M6RMyVzbAhiPA32z8oVPPeJowyDDjPkYNam8g8
qkTTb1L9JOaw59rfMjLfzzoRzIuLTUkwBRN4+FCVfvSr07rqgYSrnT421j22doyh
z9RNwNjYwEITfJgs3ZjuKKpfSGtR6yDSWdsMYFLZtBs5bdLWEfNLvVbh/oGTk80O
ps5fwPgSy3uJbjcGP3K+OsfQ26l/+ASJ5lGsUf5dPn/7RNZgN8jwWJHtkI9+YqD4
RgrcS8tihkD25Tn9U1Koc32491/c2r071UEG6++/IjUQ7DdNoHx48MpBA4pzMlUf
y6S47x2mOofxeqNeH1rkAV25siQlppH6Rhg+FeE+c0xaW4mVhrUnVaGM0kn67saA
GOs7Lc8MBKJTIzIxJhUBVdcBpBxVHUGQ0eC0GznpNC+6WOpoihB5CR05Jph9SDtL
B+CSyQMXewgPB9DgacU3ncRKb3/I3YaGD4kVztGDU+h+WxOs89B4DZQFoSRnf34K
wTS5nHBjIDeqgnwQUK3FANpS0Ghl6CmE+3IQ1pHEQ4wqrgROwsP1WT5Jp7l1qLzo
3A7ZqIQWDjq1EtJ4PYX+oSWP6H7JfYf1EkCjQbXxSsI7mx4svO+7l7RXKAUUsPYA
pzDSwDdtoih8dhEoY7zIPO9FxsAEqDYlpXnXi5yDNTla4363WCKRf+pIQKbL0+wL
QmVhx4KuPHCeKbgAdObzEhJNlL/aOiHKRruE01ojaVnLiXgpuydx2vZpP0/MQ11D
B8eAwobB3/XW4lQxyZrYwFR1u3Pcfi8XKJq7CIrYbqbZJJR2gfwjh6YBnjcU5cWe
8xXkb7sJN/4DoUBNszEPtFbMwWgWeytjJbV4LrzpdCFTBSOlmVwI0W0mNPbvObU2
kPI5kIxWkp8GBAtHbyRSDGjQeC995hxYCSMY0Obw6wildUpZBbMl9nhRvj66JRji
83iLaGhYT8JyadQgfvbM0mnsdf5qa+IbTlbfGXu0nmf1n9r4ZiLm1jMT41RrFec1
VFKzWWKVcg81xi2BSUG0IO/T3gWoVmzwh8GqJlTeK2jDQ563Al1/j/ggQ6s5Lvk9
vyCNdCIS5s/CSYFZfMQZklDBGEdX+jBC1U/NdelwSpxs/wCrPX4NgvkjXbuUPL3X
PjM1cUq1NgsYjLokHx/QA1sgnhUqGCa3cxv/KDCK8WSmWNDxO0eyfKuJL6kaVcY+
amIUYUVOqY0kDwVIzmUYqpylRkU1LL1TvAu4RiJd/8jND+XsaT5Dleg22P4ThuCI
RF+txP/ujxQbQIdj/vXNWn8Pkg2GXoUeyzfPrANh+wyp9dC1C43KhuFJp5CxKX88
N/gshYP6ob2xjfLctatSiYXXEza2beHeBYttEhlFL1mltRSK8rZbW8xDNO7yzeYB
/yToMjOOdH7BOfiYeBfqPmWx8ND5FASX3froIuU48VzMZidy5zzolH3s4kQgOJLx
tY99Q81gfdp/sIEUhyUKoGghiOPL52F0dwB7JvwTk3DpOvB1VDJu11+bBYxG4MNb
WRqSHzt0giJDgOd5iaF/PlekK8HLVD3K8ziLkSNiYeXbhzhpEKRXzs2cog4j265m
kRrj1ZMKNcFsXP+TRZqO/cnks2Zbzc73MnE+vfIilq52kuYKs3fL7OBwmT4uAR7e
n/vMXfB9QB/ouTtJdCb1IRGKmRKcu5AhdbH8F4Itp7DbB2MhGfhjfMkOr0GoJYIH
KhpFl+RsoaXJJjilMj/FKd+Lw0HumvsSedTniNXrvKySuCFlxBf6vVLJRoghIIII
T4GrWjy0KMrjPIDomaoAZ2WeTOQMo4c+ZUFMtakIR9d2/ofRYcTUIMevft1sy5zi
DRA0GFMGWUODijKJYUkwH/cxkApkPPQv+W0pp9yVVfyzZ/KLcmVCQgfAKz7BV6L1
eFMjMesW2GSvwJdAUUt9/csjMIYVB74OaTkkv1nlgeao0/3fLoumUkKUfyhWMUIF
1uRbsrSh5Fj5nsKEZTcbCz8m+StHgQyywF79dVKMU7ztSTYK56OqCGIdcjsHb+HO
8AlSsgJuAxtytQN8AZFE4Wq9xG/CojKtGm27gXnWFdpjAfiLMfykh3ZN8/TORAC+
0+xiRJGFY55c7FBlXUFqTvUIJRxLfJ0Hsqk3aHtVfAxi/KaZronCzHrZo891M533
OKRDW4VNQgZf8exsvaquVydKeqrlJf4rW4JwL5joqymXap9C+u5XyR5fWO56Xpxd
96wlcq0D0dE+Y78t6HKcHhtUk0x3oSq2PQfAQrjACnCrSXKNbyuOcC21DXg4wpVh
5689p26wM0c/akTj6a121crzRkOjSZ80Cc3s9ginQVtAZQrB0FD5jBQP5JyS6lx/
bu26F9rzAchqFqCYO4N6og2DzN++/aGVGrRrMbQZ2ga/9rAfGy3tbyYoBnyyeSf6
BRleJUniPACK2fE4+mNrbzsbMSxJMf1GQ7JepYwd9xJxFbblZYLmORerJUJABQfa
XlfB84/zh1+9piWzAkrkRt405AH2lS247iONlOXu1QJjMG1+oi0rUmmGbUR1CVJX
pameA/fmenKyl8pzUnGe9zPc9siaK24tYMkP5sfeK7hCSAzLdUS9qpkP0+GyBYqh
zCbEW1oJtkWc9Sku9X7IJN8QwRZKqwisS04SsH0lfdjrNfmXweG+HypWHLBA7/gl
NNbEwq8seAzkNFnb+lvVJ6MgLNPxaxlBv4tCbZ2aKJIYbF2jKvOnhEd0zd4gVyrQ
A8YB1I8v9tubb5K9dbPxXE6bYSFdPYZrbp7u14Jnp8JK8ixBPH8DbhyjQxb1npIx
jhLlyzMx8WAo5g/h9wc1RI3jxp3y7rgNcsrsxlLxbfbG20+E5ybHvVpKMrO1flhI
2d4AQ8WSaiVSTbVK0AsupSVJBvGbKo3Rg/VvgekBn0dMgoiGCcVnfSCN4SD0qYM2
0Zk6C4D2Qb07JrPxOVZX9QQL15LboVM0Xma47T9u/qMLZkXj2df/nnZQqplUsiFP
uTHWB0LfzfjEV1uJYvRqK4VU+VJwQVUVp766z3saMhd4DyyxoKTVLIvN963MyQdU
vsmBx/lSMJNRACMLDHe6KveJR5MpQBzQnYMAwlbsuxcT3hgBwCxQUoIYUcRUE+sW
C84XWhU/p2ts1SQ3mpl//18Vr60lk5tvi5M3qBZe8jDIa2DF6P8NII81ohz58+aL
r/fetg5fTgGKVf5cy/3WO6IuV0KQhJcbsFEFTRAdjMooBCfIvpP3Mj5un9wZSMfN
gevgfmTUUQnYIWAzgDo5SOpnfSKYnM3yfXUdmfeL+MNEz781bgp8MREMc+PIEuP7
OHCMyYfCE4wdcir6h+dl84Zkh2AUUeHAmc+G9sg3WiS5jAWKtFBOKtnHQ4a6+tVt
ka0HVYD6j+9YwNPBKzsZUz37h5u01koExITAD+utRxS0yBI4NHrB8X49XxYhyfuA
PpNaEZ67uGFnNpwVkiWKlmv2AzNkY4bex7pbWF5uEq51oBxEulGO7EXhIKVFmOiz
V64PGpeS//H+JZAopPgbrQvhPpeG5aWtMTG5futI+Def8lwRMeKacBzubMNbGMs9
RS7bFfgQDEzYuSssdplYjKY9twUxxrZfxJYuWjRlW37YqarqgJO3JZXxokAzTfC1
X8WZAbKKZxXScT36YhzUVj0dZ8VNrm7H8IH8i4XUHg4NtNj3ywvEQVeETQWWCx/J
58ea/a+9Bo5qLUXuJkFSSMhfbI7a5aelH7njd5ukZRFCgRDxMScTg88un+9OIFri
VBItwwasBMkuZokT7BT1ww7sYSK8mjprkDeqnL/sAnods0zFN/9WkZv8HvYmshhQ
q00JRo+DLxHeUzzb/TWXj2pUBUyu0zzasMt5esmv+1ynshUY3mORSjCmji2k6viX
iGG7s3Revt0IrRfNvoryeLgVGCvlKAfXt7ZimbKSdEWjVaUnJay7su992fQqg1le
uV9pucZ7AVjKBGMj4cxpWc8XqN9T8Av7BZK+jhatyraCYbr6VzOIhFuua+YmsCNk
oLa8e70JxD1TVjp7wJf+H7DqCbmRypnKq3QrXmEdp+4lhU5ivBH8mYw14M3CpD1b
THp7RKHYZtwkTwz2Vt6d8PiRVyUKJO6Y0njX4rZP0GOsF5HJrcAO3UghVWiGT6qi
LJY4Z1AHUNFIqVi+vpYC8CvKj15hbPKvQpxsIQvKYPMKbSUjJg17v1Tgxr4vwfQN
Gy3Di0yMZWhxCNiNBwBD1iQJuza1KJ1h2w1EX3d4jWZXc2TnGL5w/X3na4kgywtf
2PK9btnaCSni7UVnW6d2PyxI1wPqzgPXBxU8b5cIAoSN+7gllzzp8iqSFfO+DIwD
/dmmI2ZpLKKO+Yzm8QafZITUPk0KO6+8RQ/NHnbSZVPo+srH3IJ+YgHHBVBTGR48
1X+J4mQQAJoo8LAW3BB1hctPKSPzuKJIdXVY6Pf8SABLZKktkmDdtqpSgZbzeBvf
Ri2YwjNqkGlN2Fc4BTk/7ZhXSgXqyJxIJKG35RjNwb1I9Z3UsxcuRWqHDzkrCGBg
B8akmE/Oj/dBia60yGd0XmZ4DWSteQ8JZJdeS83EYLJnCi8S+fSHVGSFp0CzbfNL
iUYeQB1AIb5LqUC0RH+s2NazmYflkGyTduMP1Ya2qhiqTyiHhlmccPexmbwHnwhE
Z62BYMo0pgqRjs5jnol2BwJntPINvRCrVWgIPslKAf6EPX2N5y3pB1ayzNLkEhXA
e9r+9O1obfCBxqOS8oSpH4AxsksZ4YjtWLvBaCd9niaZds4CPlYdsAE5Hlb8Rat0
SNMEXEYbCv5+tc1xCe/9sl8V5IE28kvV7V6r98tV//CdT2sJp63V8zTKKdAw0spm
WIzjs2hhY0oHSF1RZETVAPnIpDormfIzya4p5tNUtXNYD+lvaZ3CwuUhTb0DDvZ4
oID6f+fD+6hFny5tfr5f15oleottl0N1k+aslXcArKxhb3kQ+/L97PDfMzw71B0x
3Y+ZxccnQ0aDSOR5Rx9plR4fnPi/jAUS2xcA4DXc0XBIQ9CUljd/tkbWiOhE1DBy
4Mgf9vCOq8m1zcQTvzL6Z3vW+vUA1OzcMzNImloO+T529nUlYkbQ3j1bJH/nEudz
b3VxpGfIClB57cjt2Rr4CBhrryAzqyy9VH2ATjIxHECpghCyqJ7NdkUKjW/NVm7j
nBLStjvVYAnMh8RwNpFgNwXS7xMy5dvOyXsdHPKq+u7fb4ljt2yIN1CxBelU7MJF
ep9nCMOkMB5wGaEyqbFioEQowpyd7ZjYzv4cvL4uehBuozIMaO3Fsoy51DpjFzTT
HVvfqPQpGPYcStLap/dY0XAsWxQaCmVgf5l9ebXhrKQqD6gjAWSj0a9tdTSkjHTt
Kk93SjRuPOK9aBNzMRAbCVfyIS6euCRVEg2EZs1Cr7eguK4NRMyPPqthW4K1Fc5r
ey3/jPQXetpGD6q0+zuubqD2pJrobmSZCI17yjBgtocAL6tISReVQlHxFi4CC3Pi
x6HAeAnLMYQe3prTzD0fB6hShFUC+UHN1ZtD7zRm7gQDFEpxLoTh62tCMysNZHZl
C3BXAyr2acHaWip0g9Fp+PetcmnpC5syRxMxyojJDo9RSob1/SS3/DRyUk7Utr8j
WOagTeOOqhSxglhKHaSKphxhm/h7g3udtM6LnCHqEFWj3y3+wjzBckm7GNn4Eume
M4X/ijA6QoZnonae0cnoEHcxoJGwPt/INKC4AY7Jq1BmhatFtth4+GUgG7bDTOam
WJBja7q+gFXDTKL0TeF4+1CoC3GbdP6sBZQpBpX2CvZxYS4jOdpoldFkhhSp69mR
mI9xdf9K1EN1FdqFW900N50wwZ9VUJo/gPCmM0sBhtLSuJH0olxpydJ6THVkt7jb
ZpPowQzfWBs8X821ayZxtxUv9nQG9ospez8oYBkj9RMFO7jpFai5C3ztBroesvGz
NcWRo2lyemFg0U1X2A44fcEd5mj1M/ors6XTWk+8iLcB4vrZOP+7yaN1J8mu9FfF
pEWtN/lf4Kt9r0/oq2WaysTOW0hIpdfG83hEvEuyQGbnHC2R/qDcoWUWqpN6adlp
cUSP6yTybWgeYVLcrA6GNh2EAZrn6qIvuDL1wbYe6oa+r1Lc1QMW0APs/k/KH366
BMO83biPeywUAaapaBSccMapPxO+Gw/skIZeMkejMaUeP8Y8vRX/3lQPLBCxHJGa
rB9cQBVG1GkH9SEFpYLVhBgY/5FuDFrkQMXdV6xAPvX0ey7kr+5P5vJywOZZ0Ptn
CRopXQT7nck1zEq39rEHgP6LWyPSEGETI8mdir86boupo2GDgYxjL34bMDYIYlLS
6ETwu2jEng1UEe8SQLrp/DKLTkOYDRWOz+MDyYqV1WL9Dhs3i4S/qX0eJU3XS4EU
v9MHx1a+x5WLpmfFWdlaVZTo0xwJ1L1xO11F+WMp5qEXH0wbT77kOzCt81LJ+P36
Wtr7WlbAw6IczE6NJtDyVrOyKskIE5cGQwFxJp0x3vFusX5Tgde3X9jV1KBM6b/K
kuGKsQxRIo+c11zSMvfEP/koBMnB/FCq56Jh7tnhQ3cdYZHkHOGMsWftY8fj0mS+
CM+BI4iuDd8MpfvtwqXsNnxRujHNLe6Zm8xkaUlAPcqHhnoGSF5x00AixGlfyHYc
2ob9rNsmKT3/TcCgeJWcVQkz/bZJq5FmZi7cbJm+jsMJ3htauT+jR9H5MTXWQc6Y
cSfO3HHtuAvh2SRh97ARu85lA6pOBHlsUoB17x918T6kr3+FoFdDfQVaJYSk+XGL
03dVryJmsfsmIdjx6BqccuTXS2J14amIj18o8suHUcDTNAa7Vt4c2RLMNjm0rJhg
Dnof6QFCJ0ZSJ+GV0Bky8fP0OHAZ2sjMu8HZ3zoCeql9Tai5StOAx18Y2dBZGwEn
DFAnN+cc1ameSuu6aY3nbRF0JDvY7CSOYCiDSIp6FnS+b+//MAuPkGJq8IzblUwd
H0GbSUwlZyDosiI2wEptky8AixGlg/V2AzQuHXc00g1VBheez16gSNvaYmRqRKWt
N+QDVekkpKwsMSJfrFa/HfcNr4Wv/SdoM5uNyWbRs30rnjw0wYgfiwpL0yl1DGhg
siwGDXCcX5AlUjqwHOQgZwcGQsPeSLBDgy0+VSmPjlZSZFpcVlwWFYHPKPXF8NiX
mMjHCNxj1/+m1p8fMEnfHNE1cahVmGQpAyXGHCRE+KwzR2JkIGik12eBqwzVRpUF
ri1If/LIgOTenH+mT4XMe+cuCI1lSnNE+LrSfWvr48sJ5qFvNhvGbFfOdsan9e/i
oWgkAy/LYVVuNQ6K7nO5V1DoXrHFG1tQlo/L/Do15W6fgqvXDecRim2gbpAxmU/S
ClRitzI8T5fXCE7nAnU1bNX1JQeBqi7o6T1TJSIDF1J6n+OQ2gRY1wVxpaXci/SJ
Hp1FDoMtsaT8sdAuSC+41R+mMBQtUxFFqWM51zus+Ztu4PTWZQk1HuiT+6UAvtrM
ozvIjnNcGqtLoLYpeg9K558uibvR2U+bArFPgjJTIJqSJ1jo6kwewPX0zZpCGx47
GVOJAu5DhVfxCUF7FKRP2GT2Pe7EkKdRW/MosXz8FdiD8P/y7IidV2ZRjc7oC6hl
R1KO0RTWhrYmVPC6KssHz/xDGgzbc/ErUs9pMlW8UGrcSXw6YPIwE7e/Ey823D/o
45pXQkZq3nQvoBuDHBMdtJweSsrEXo5ecw5pMv13fGYPVA8Ki6l1EKuMLmONLEZz
AlDg6rDSvbPmAomI2pKz6IQ/6ShQJe9cniozOuruKQ6+lL1zIqMvezwjatyo2qzf
5GeB2Lt3ikYxKepIcnbJNcjN1+mjCZZKGPTiwBc5Ob9I3+cfax8SV055LBGHPz1T
KA0Xru1GPrm51k7W9t+bBqxifq3L0do1mVRIJnKkZYGu99YlY6BLXZQNglMJYLO3
/Ed3DjKGk/EJsmBy0JEHgzt/wqRoxC+gkcr4kB2dKikAc0JIH/oz6KYLnDE+ZKHZ
uZUt5Mg1LM60qEWFGeWYjgUyoT5UMEbTTDKOv7E0MbyH15advCNWCu0MUwjZK353
2KIfleS1RM18Zj9lwkT3YRDZCC7UQLbQKUzpQklGmrfTMq/Hpfv3BpV3Q4YGUZwq
lTZY4qtMd+YYaDj53B4UxRL1NDkGRvN87D81RTz+RiPHH6B7FYIbKY79njdK4hMh
X9ru6N2bLjNj0Auh9B1aiEkPGTy723bv4FF66l8XhY5CgDCsOif9IHZxvgwpqHt+
FoKrmZPfBGZCF4zK13WIzlm56/+sEbdFA/ftXCoW7IlB55oQVnffGhFbSMoqWbVh
KVw0b6AR5q9IDlhG8SvBn8h1u7wX1nR3gAO5ciuWf+nEnTcxdPG20hVRFXEA0xcL
DxiWOKjodneVewHxuwJJ7/JaKH0ie6pSVr+8u9kQoYc1dAwZqrK2CKkejKUCQEOr
sP/DvFQEW+Vq+o0hOnzyTqbwHbOjMMNHk8w8wyZ+/eZnrDEhpwdCyVMCg7F0fdy1
UjlmkZOYb7Hib+Gih5OuraOeDVoKXS1f4IAlPw7px2CC60fRYZwtNVWsD0zW0cdF
vKfybtkuO4J7bth7Zska3EfTpQ7waOI/+aGqLPyQEUK1uRx/x2anHThly4/fGvzH
CUknR8hChouky/XAnQ6lm3Zh6UI/A+/d2ZbI1fSog1maDwVXnLu5n17JPwOKu25+
DWInaoLmzksgRLSmYc1QoNb7AtNLA654GjwDRluydP6gnEbfcde4YAsYQo8QdMYg
SgaL3rqQacfQO6kehdgjddnD5b+z1zZFlqRt8Z72O5BC7vfjayVAuclpWryIldeC
GMl3kh2Dk22YB3YOnMtEorZO1zqjHOFN/BQeawD+aZ+FsGqT6HkW9EDi2LUCkA0R
0FJnuqLnnGb0MHMu17lklnz21Uo33/r41DTa8gV1HOVROa9WL4TvLy37Tj/ny1mL
Hd3iK3Vciyu0kpPyT/pamsusZrFLYgw/J8NF99jQATan91E83Z/kz9ZCd/Zf6kHK
ckyXH+tHiC2X2bQS1KV/X7KmQBWEnors3TUknWFtxOBdnxREdcQkYmxxw9/mz1Vx
IStiLLR09oEyZE0WkCrhBAzX0FjxdEZQ2mPAN4+hppCI6dKzNTT75hMQu5UvdHCp
95uK80oV/sDhDy8MD51EKxVJtcLmwuTF3FrVeqheQj9oGYooN1kbC+cN2Jy7zw9v
FNVot8G7S6Oyq0Ewviy3nsRA8UME3zyR9ZhkjqteLlhIr9ApPIQPVcEa2ZuGKrIO
P2cYBln2uaDwRHsdZdY8vplGQ1nkSbwtUwdpZ3kDd9k4X7wMwlFIC046UbFctrux
GlISgVzKc4P/g3GsQVKC9gWckuZisqqB3AqAOpO5e08hjJS6NHS160JF8ks1A6sZ
X+ElMZ7CR6FEQMQ/+SKl3K8hF+QmrH22ABtYMnGcHY8W1qhMFXFZUJksKxFWV7Tz
o5S3rUZnT/PepodavLV3pfaKX+0DaVQgI7nND9lCGo1ExaV9G7/qChiZHrv5/YBF
4mMkFaFD6WkLH1l19GFmxGty6d5Wj2O81JaxYGuCsUBS4xAYZil6yKz20vJiSi3m
c7GkDMmW8wXc8Oj8CdiKovx2e81b3+waisrg+hmHug9bTiUPkTI10RkJPezBPJ14
KilLFvtAYbhoIXBefrV1K2MkciVkloIwTdfUt1s3avORd+kGJK8LCHhfY6QDs9+/
ZUvktk4472pr9MzTc/rnpmGL6uU6c9+JAKlncF8CD9m+qz1AY0B2fZ0DzeOBtueA
EJen09BTsnJ2nu8qsGaBWUYUcxRJn6d3D9uCuvpEjrqmHn4OPAVODLJGPpcs8Ehk
WYr6SuhuONbWoQd7Zw2sTGGbvonc8cZge7W0PFZlk+5DbGS7oAi1TU55xyqIWya/
zrygMg143QavQ5Y3LaoFfYlJREO0quUb7yZWFCFhCjQZes2p0qhXTFAPCQKla55S
vGXT0Da7N5+17LHQElpXHjBSnzXnQgZ4XU+HEnOQCx/zx4TC2WfekNBKOfGeps+d
zNW7fOQKgvxiAwAxQMAzifv04EC7DM0SeXv/IXuKB8YwD9uE5A5JnHstp4ludBd4
Y+18cRnGPgKBiUlukIC2UOXM3k96BGcf4gpEBpMPtU+1nybR+p/wFMiY1CONDLz3
u/pZtP8pCKxpRSlAuISkpYdpRS1hFI00J9PknjNpo+Q63XiUBSt9AK9Lu7w14y1/
keqD4A8QHanyooeiEaXQfpZpl0vMsA8wIUuHO5YcJUY6MTLtqDqK0aLD7O7IJtqT
+xq8JXpIJQ0txy31BGp28iUPzWn3qUP0JVxlf6FRFKjdEDi431WPc+oWHQnIuXdU
3PQNwkZ3KjgXPTrPBfqangxLXsuWaZMlqIpTNnWTBYSTcaGxZnhVOYHJN9tQTCSs
d5LYyVhDwJHQDuLJhiueSQpXWkmSX5sghvab3XBW4GPuQeQnUuJM8qamjcHkHUTV
FDY+cWCtMm9NelSpFoIAkId6VlsBEfwHm+U9V0NpNEO7J999YRt0T8r5XnyAuA5c
fsUScZayXm1M3xDC48DkCuN9RFDrou4onqWEOxmP9h9hdU08mWzQuokT2uCrCGbR
yY27WWrPnTznWiUqmXqqpcxoQHzBD+6Wk37jfa7D6BrfoHDwaBnIvze/0GP3aJ2w
DedoRbeBK99z5c9YQKwrYwMPgXJ61/as+eghf2VV0LT89YIkL4DLboWMGSLZBbMO
JUv6LybwVo/2pPO9MQGagarNld8erEXoctACoRmrXlJa6gbyMaXOU+9h3iNzaUri
/8fW678mA5lWZK+xzsmqzpQFrXX/IxKwz4OL+E0MRuL4ofjdaMzBV9+99EelYDcI
ndNPom1rSLMxhaAeCgtygpIpRZZWtDoyXFdKzN7IRc7309bxTkHlu/91xe6AUQRn
IlRXrMEFJm7wa8ZqSUa+v3Xh7wBukpjgzJBFjxOawB5S8G4js4FVbZeYSr7/8eZX
cciyVm0C862ba+TTr6o6v6VccK7CdFW76TiX/A9SGv3hE95m8U6DPnEHjj61ZR5L
I3fhbm3/KREhwwbYBbwaEejgztUDMXxIAtK25bn6W+ewVeXnwfxc9qEAQFMNmO2p
3Umk4i9JBYV4BnLtRN9MPHWoVmXt+8/E2Ge2vSvqszAevDxX13xRVy6408CZQ4D9
w46Yk7gsU8fEREzyrEmFbDu4DVO2gF3Yzv/cTM+vMNwgXtQTGjBeqUiT6Xvi7ijW
39C/SZmTF6O8RvfNaaF5qwB8qPs6pYNtwtfv1csZ6YWg2HakGX/aKVNe9nLOelsL
s5gK9G/XJUNo2gSrouTPYqCA5qM3qWKQHLe74IUvVm1tDJiHE1L52MrwBkWroOtA
efnnOXsS8QdMh2Gngj5liU8eR+UfCs5G0Bxvu7WPzIYzLdVzYmK6AXvvFUWQD87q
LwZFgSM6/tCen5vztTuvNMB7jbYDHrI50n0pi0IkqASX6+ugN4gqjPmw+v7vtct5
vcDo6J/Izxn3OWjIjs8ynIbvNigomZRZ4koKxKiSdAxv6oH7GW9Z/GyMw+x619dl
urUXeuLH7aOoqKOzLBhv970NTlsYP88rQO+gwV07niZBClluKhvg/13YTCdRkHfE
cc+h8V6aQ0PkWzisL6TwV4brxsPjpPhcRW2CyXjHwjwBRE1jCbYlqRNOX+7TZ3ff
EFFxnkXDhAT8n7OL90HDCAakBTip0LTmv9R1Porb+jYOxurpnjrymIakd4iR8cP/
6DgrLmue2zjrJ4NEAd9pqylHOnSv0V4TJPKs2Kz7Amqa9rjI6V80UbuOyRTTl7dl
/XswJMPBPgDRCKI2IDWInbBAW/bnoQ6wgnbIkb1o2GHcRLcpDApoomZJz+y4X2/c
svvP5OxJUnnu8Bvsks8KwOFI8TbDF9GtViUGjcEY8nlZMMnvU/jJZuJf8nsJwPL2
byYjYPVLQQ924H6unlEOHOoVrp7FgUz0SBm2G68DiB+RTLcciW+0d7+0qzMAvbAE
PBecltkcQHJPn7xmCU7o9d8ZFvi4XUAjmbJZyatfXL8mEVgex1vGixE7J2Ng+XP9
/eNAiXd9iQhJCFB2H8sAhSgGs3gpFXNvjrO26uGu+0PohOI2bNlrxCdwwY0lbRR3
6ZIk6sEv0Wwa92kCHID5Eb0L0hiH8anNwcmewQyb391qk/MnaZI/P9H7E9WMs27C
kpaOwHdJRn8d5xuzyY6jSiiXluj1CsDNZiinuXzpnMQVIwRoDPlhpQZq1JeWSpiV
oy27MIbFWGTG5o9J5DelWeoQ5gZNcXp+x1wQz1+3vVg16/InqlwkpAICoMUlTWb/
svOBrF3lQAOlHx/xwFGonrgYPENgr+MJjUjgKjWOj0OIK9mo/xG8bDzk0ZUFbf2R
yjNCLfWC1UiQ99l1aw+uM3s665Mrvy0X8SI4w8S7gvsBFr1MW6RhZLUf2d346Uux
HUFwr0CLUUGAmlLWuA2DXfW878P7+dRNCtvEQgywINy7pAaV38EVAKSiyA/beztH
SDcv0+p/ouQ+ZMVGyXTbqq4pbQH2wdjjToVeZYb8gDYFUkd96hfN/2zhozJDBhNP
Cyr/g65tSvu0O6SVZ5J+agbQ96JfxWCE7dHtU568ALOMukfwY4Qz6IAQrzo41EGY
+OSq5fl7EFsSoKS4nFBxqww1rImexcpPFs59VxSmRnZpTUbR8DtVybVYnijvwzo/
80MvbMipwiybeht63wv/RnhpbytVYa7g0hU3qZzHAdCfLJsirrz92EfU3U5a5qpK
A/jS6YxXM5BXVpsPuVVLeKO/iAMUiSI40ADQ1k456VQ8SZGkAbdmb8J5d1XtlBHP
QOd9lxy9DrqzXKl1I47ToGsxp5CAHxRcOriS6YrQummr/dWHDbweDOFy/kJFrFGD
INqzyiT/6TtFOC/aTDtCOuWET/F/hUUuW03NguUJ52n7Nc5jfCDW2l00LcksKSya
j8z8kNc57QqL5sZ8+SB9HlEb0KVn5FqkUYvY1NRd1oqyO2tSB7IxI90EiJcWxshS
TGnY7gTKUkXRNjctw3wf+r7TBjuc3lEGSSlJ1gp76tCyJ5D4gWa0gUBsRz7N2RYD
x+1+fdY/KR8ZX8awpYFJwKKSKxuhCz9LK4iNY9kRD/x84nUoqKKwuDuxp2DX84My
gBqvyTq8nN5Vbi3EuyQayQ/p6/uiRvOaDcB7KBMyUADe9NUkOiybQVBWER4AoguG
jZmfKVkk5XrDANCeSulxab7g021TecWGJUGTCJhVZSubmkbYhswBPv30GoloRlhx
YYUAI7cNtv2uE73nRJBMR1cRbk5y0NLPcFFhZUDlDMnT3p7dKRx/X8ft6irFpd4r
i++LymLRxkzxIggHTja5pKeGY+IsQ6RJ5iNLOzmUPeXo3WWGEaV+sMQ98LcnvGzd
MzbTcZCab1J6aBWZZcmPDYS0Sq5BIvGUtkKe6/rJX7WX+u0VTIh06FlDav4Hu+30
I+YxFep3KRG4ebThPWuVPerBaH50mLOS18irDQC+AOQ9kvct66PoE4uX1XSPggdS
BqO4lA06ZBgtlyWmD2T9YC8WYeTFAQew3CvmjgGzJRbU7+4d/szoy9XlVCDVzucU
dW2VTieflVniPG1/hQQllqNtv0+npqOFFbMK1+bwC+vPr4js5DfsSAW95p2ZW2xB
qTOrav49Zf+fjDiEhFSMaMragGBiITwsRzBWbtllbOg9cWLuEslzRwOjRse49kQq
3JTzhButrNePIx/qtUTXAuoF/sC8V+Sy9J0RGqUmUuAtJDH15lOAQHOnC9t0VLkR
+8I28QojsCgk9QYIvEy38YehWA1Dyn+rqsQ/xaeLHbgYaCd+K8aHVa8E1LnjiLrY
4+41PXQmAeVND7ON7sfCPFoYwhRfW2gFUEbe6khUBVqdeu+eWls4oyEK8g7BHgQI
xP0yP7Hr8i5skibvtRmDg5UJUrdmb5Y16Pk0jWCGuNZkxA/6TeEHQwVClBHV7DDk
8TJf5wKXlPPP3+KED3UAWwqJQubbMwCa91n4QmQ1dQ7cG6FjmgyuHXcE46hTekjl
NNk8y+qpwpzp+Aazkkgu8N6bwTNvrc5lIsygdo8uq6CsvgUopLcHfCkORsc4cpqp
l+AOdpaFxd0IijdC+OCLaRONmTAPxBceZis8kEY4zOZhsl4LEFzv5gikfE0a4IV0
BG5+BdFDFw1u/q9u0n8eg02M8iY0dVVFcHTSndimygvvUk/0VmSHLZtjaJlJZlBP
TIwGEo231Hq0U4OFXMYu+i2EbC+8a9hi0QxQrPl3Qv9yBMcAReDOgOoDGRVLLaTE
IxGcfXJ7kft7V9cqPfOcycMo6NY0aTbR1rXMDQhgAuMvImgKbN6037l7mDMxeExi
1Dkeq20SPi4dRHFTqJljJuSCGvJEkTpSD/MilPBrR+QceVNCAJpbu3DXRonVVp7q
DZ9vmF3fgQs9Cf+qDh32b7+nNgDrsPzKQUIZY5SfWLbaAY7XYR2WeWSfQQ4WGtWl
xK7DbV9lLjPAuamqP5bsAFCsKvDNwldvPwS3WlsqPYCiyGoZhhbbDKa8yqMCjveS
CeZ5BIzgq1KNhk4o4paar9Fcf6vD028R1hQ1qjiNz2VRzQmqnTOH2aYtFM4bbtzh
f+e1t5Bkdlmcek6xHBeCAlHVyG4UG2TjzIdSnBAoz8Ecg86M17fDYQiQDq/ZN8in
X42ptpL4dWrIuNfpx/8s/n63kEMMhXkl54m81wTvL9A9Ek2dVnzUiJWHbsJmlkJ1
fVMKBfxhv/wa81MbHJH+Ow02L80Z+1FZAhfXK7XoZkpDnCKZql9nJ1UJabkDdoXA
6AxOCH5S/8ldSoCry2divEzSCDJEM6Z7sWqrMmJZqnas0+fIFWvuWHU2A1njkKR3
aZ3FFyKgfaAQmSjFxb7ILDAAkDJfq8ZXCeylDLuLWXLC9+mM64IiQUogJHiTrkNb
RXZWy4SUUos/zGTh6vhSKVt5ljqQsepGeZSwFAKCLcR8q0EsDtGTTxv0L2aZGeLZ
Hx7Xc/+bzKBL/NaUMdVmMNR/mREc5FybvE3txiEQI0jTRx2E9MmkV3YX+LhaXQgQ
7GpHFxH5/v4M/Cu6wsirD0Sz83dgPS8s946LfQSLhVOSijZ/6wYJ1FcxZGuoHlbF
MIprkoZeQ947nGJeUYMpSdvqN8iILC/T1Wnpwnr4FW73bzseDKUBC7kets7Q/VA2
ij9CFvdY1un/uI2XxHBQ5WpKZpgERuvyaZv2XbrOabQ8TQ2woHzjg2SIoSAfXgT1
1vtSSYpoeTGfz5cbLlwty2djBdq6FusWP7ctZD0qI2sR5jlPNCpW+y0fdzwcVtoD
KzVyuyFcMJhZdW1naOkv0kCIj2ezOdKT3Mo+aCDSyYuFTm+k0LOnqHboHGzih8nA
YuzIorqUK6m/aJhucvyAU+5Kpk3MwCuZvpmFxoBwCkWdNbfs/lHWeycIXlp76Vun
HD9KRqnXKYLxKkcHG4Rp0HUZ1r8s6jmce5XN5Q61x2MOKsOvb9b/vXhugATm+J38
GJpcDTNeeDhtHyIusHQLYNRLR/4pW6AMyRoCbP6fWfv9GzdMk5Ez4InR8c0UID9S
os3sTERaHQd0d27wa6XoF1OUv8vpdVsh4BfcImFa38fZRU3KWAI9eZo60gBkJd4S
LPVvr7mThVGTn8G2fYyLBOhGNI5dDz2gBvV8TuxkJ6z/M5lzSr/vPEpWBx9DwPgl
S6euvPa1BrRG5Jf0FUBTTre6Ayk7bw0X8vyTfzeCrDCrHWP+cniP1Pfhp0IjSO35
Jlp/qK2p2ufi/6p6l1nL5uTKAGhk/VtU1///tM9j/B3FTTuIdc61flce3zxm8lv7
FCp59Qyjc5D4WYRGRvNfF6iRxf5ZJn9S9Fk/3QbXxS+CqJNnVwwaHwLpyce/258C
29e+c6GZ976Hfyp+ivowDlaVxnPmnkJ/ty+fTXN9XM3efA9LRZlfxetxu9pwxM2x
grXxLGTkogMUDr5E/GPQuVUychViPqQfu5XzNTNp+AuvOg4Js0ujc6QzV9jX43po
HlFZy/TPCaud25iROwAPyktF+zFMlDnl38TEuzwDw5RTrbhgruMl24Y6d/NFCt0X
PhMMgEG1mwscguOEDEmvTYwGashkNFQajZXHjj+Ft3BnMcIYsFpM8Cf+SXLsMeHh
5Yo8tf6MPKXqtgNAI3a1Q5uGnte6wWq6DQSxvCh2j5kKBvwi2Z+s4XU5ATThfnFn
Wg6INP7kgMbRmX9t3uypeanqHlvsgZJlGO8FKR3H9qeKGwWvVAHTiYTvTq+AXJCt
UrMwrSYEDsO4OxPZuHo6q5l/2AXagxnRsD2Ne4XFAguLYI9vkHN5fvrct7yi4rNt
ZHLbWriK9hwwxfa4MC7TYgHPu4dL0PQB0Dq93DVCROUZnUPWF24HZgWQC1U6uVra
1zYQaQOQ0lQLDQU4XlO30AoJy2mzR6Fe1hPf1nNlZT9/iHmvVmMOoz7leWBqby+k
yxGmW1ghB63o2xhSy7RGLwnsBh3yIl2j9iJFOdBTV/ChaPhgjxu/ala/w0bjtIkX
+vgXAj4ZP1vV5EYSJ9ZEkuev/LGx55faIzb/LgJ+UmA+V5nWq/E2tF+7rv1b3WlP
drp0xkrog734CNGC3fDEY46qXgngxdotu3h//LgYX9OTghvDyfGi2Pd8nV2DlUSr
JYSW0wStHOe0VEsUVr93HcUjNgRHGQYuLfFQ0GTxshzbgYKZkoi80JlwvQ8/isV8
mfO9K4lhCUnOH0VtGJc+2vrX1rV0T0Cjm+7wI0mkZteCF7mfpP1P59WL6/Ysc56l
QMjDLKkb6/ukTwQZLTwfbCY3gqGVVCcbibctq7kScFKBv4Ln90BsIBxuhNGcKsjM
FRQguHdnMlwf9QTsyL6X+g4XhyEvU7L6DM89AlrMLOv5dFUi1062J7e/610HUMPz
Xuwnq9UchAmXHW4J1uFwGU8AqLCwqWrbnwmWm+p12kip63uauwX81szGrY3EJ4/x
Njodectzzz8wLNbkiQW68MB1F81zVG1MQBxZPiG+cjng3EzARF36XSUAQkddymKh
5y0bk/df3evB12accC6P+GggYMOZm0Zf2dAxQ+Qm8Hh3cbj+keljEobTjmhK60VJ
89NbPXxsLTKPtHTiQa5tUYF4PhxuF/lMvTTKtdgtFxdwxIvusSXHS0Ug7V+S3gin
5pQSK9uYk6vwFsq22AP71EEJ5ai+QCP3mpR+pA4Ju30L3g526OJjOxavyrG6gf9o
RDOlQLpbaB9EVu6ckOo99Km5KQm1wbxmUJmO1JBBHCT08CIqFBTap2RpA2IUmaPo
28IgXhuW/v+xXZ0/+b9dl3KBJxLy1hKHVzrmFqxvGdI5Y5RSXZt2lDXIC/+9ElGm
Pf5lWoHkprolEvgP4tv+ivjUCHB/HsZMgcELaUcRtNs7NjO6Gx2hL5S15r09X9rX
2W2x7sRY8MI5BB+GCwHOSCjkrJnZI+fCdF4z6HM0oPJB0WQkGcUXgj2ZbZ0vlCPJ
PhlRJKRC1PhKWVXbYjllO55P6LfxCkU5ChiaIadJOeyQSE5jJAmEWyydBRvqXl3q
gWichcPQsYF7VtxBVXnCBjDgK93/A4F3IYZM4gvDu3AhaSn2O01CzO71vTEJihZb
O7vDgR2y8AmP8ksA0/L89RSvwEE/MOS2S+RjtqIPiu4m9/v558zJFVBnbSVcgIjU
R03rSG8I0RWh2F59T4wVKUyd/IosjlLTGF9IhG5QXuea458VSkiemjr5YREa76DC
IydfYFWRFnANRAIppJU4iTJFhixc60ZE2zYJP5vN7aVaYKMQ5DN+qhM6E/1/uPy8
RQnxNtnujbgaWJi59CBJVv3Kjj11cfLbP2mQLFMpObH6FiH/IV6KbDKtY6wVvjY5
XG6p1gRbz+Z8ark7260HztaHay9J2BlX6v2cVrWcWwDabVZZfcwSj87SS1pvCfpc
wX+DEigGREI2O9WqkPqS+5JZtSmm9sSz/cz+v24i+VRHFENlIPuCYG/+F7mppFji
QfbWOy4LPoCDxZ+DdGhqRI+0newDx/gdUVvUGY1iGY//YEpq8QKdyU9j8oLOaQ7T
oDLo+xMnzW10MstDXaTd4zxyfzta/qgo3szLUVHNu1rSQpSu7SL83N9TAGWF/ffM
Xz5Enx5bqMCn+2cOaYF8oMy43kyIVXRL+LhkMH2iSNlmV7i7bEBJOVq5Z2sws39/
VSoWK2KVvplxEHUGnfU8qxl/OrfMhd/M89mgcsq7YEmHe0Pi4y+DtB0R+vne4mQS
UNfh0PcoyqOXXxJXEF/CSdTFwWHz6KBerXGE5wxzCx7Xp9qml1e127fL8+pNNGOx
mjNQXVWIXG1BCM76GZ4ZuVDRRDJmjPEKhDNDUbWi4bqkzfpgZmC9yK33vuxb5cXd
WhWSERkWNko80zxJr1wDdkTOdBPTYNrV3tH+5e1y0m46AdRSLYw/YqE895dDLXpg
YBXlDbpnGsxHJf0FEQTcfV8xnqokvUkpGCwm2L5zYCJK0gbjT7cSrGiLX6QDo3xn
HOZ9Fu3Zi4cubfAffpUof3bj9T8mlfu1+NTSkubUsqcfTuDU7j1KtSydxoEmhwxU
EdVrtRbMgbqEBu+6SpXgRRhSo+yk/J9fHEL6/GLVQMnGFeowcg5YSTRkWcUm7bC1
1TVX9wswapIkqHGHSYsBfEhIAfJFj8zoMzdW2GF79vKV4vCOg2sDM/kdaTUber42
phbA8LQbGIBL3tSuciBnU5s86lU8h8TUOKD2+QcS4C2yz5pPOeSOrgaE5DaoiWPS
WW+/araIxcQSZ8N9Qr3aLQ7Ubw5484Wc0dh17fso99JyIg5VdTGDug2hlKfultBO
lHbTTHhUJNEmQMSRLRBI/OvMFVP1H3fNyKS1fCXRn+RkLGTN7aZa//gwXp9A0SJa
Cc4wx0SSlX6AQ2o9XVnMqU19mFMZPem11dbxAFiPP5CKYj9oyB/9JYoti6cyyaAu
BbjmsU7FOQeRR5DzGTfMldes6HOJTG8ZzIAXWeMV0DsJepekeY8APlN5bE/DkzKv
A3cZFxuJktbAqyNS/CCoKKF0wxc7LxP9CnO13Kmsos5zi17hG4Vcmhg10Tm+YhIN
2QFDryxLcsCQnTH6bLIdmyc3MwS3Hh47y2K9M9UdYX5iqKZ/UQvjfaxZij72MnKC
KJag3oXB80+eUtbUN/aTrzL3j0MSSFuzW3csXIGgkaoQo5VXLXIexv3Fo/qX7/zU
vTR67HFJ2tNgT8JlfnmDipJ57xpCwO/0As4I3eIDwNaHHuVNjIegrE3nJOhr+dPe
hPhdiIpwIGbW+POLBK7/oTxogmx9cE38HW50Iz85rHvQ3dvQ68X8pl8QXqCz9dva
K2ZsaBEZ7aTXnivUcYH3WL19n7JQxaZ5l2DZ65Uo/i0qal2kvqA1+K5XciZmYbkx
w8kPaIVDwZmmwTi36xRnU86YBHVqDQ4L55J84RLdrrAH370Ebe3aqLeThlGhKxxx
0O/2xWiKXP8eoZ20uMNuZ0Tv0cSikBZIWyRSUv1VCck6Ul36+8/xjZGJyMNJUQSd
v8NwPPnxn1XxO2XlSFZYvNIOOp7gwvjtq301I7Bo1N1zS/8RjAYLb3acvQ37y8qy
katsiY74b2n3maCmUr2IbcGQa3U4tME9cmeIK8XWTxWM6B3DAPlw9fj2WXQ1BVX4
KIJJC5g0WwgY6k1LvBOmOrZKH2T9rlxLxyqvhFk9y8XXgB6LfDIPB8SAPxaqIzHa
gMoJc1wURxxQ1XYWmo1NoJhouqN6TkYmz97wKBvbb1qT4Qj4zrFpVhtqlQx9aPs1
vsrMkgjtGZP1FLXU2eI9OIRLZeSUNpQtN0l34KNq/UNp6M0Xl/VVgMePVsei2ZSr
21XLg8is1WqshBfQY0WtVs0Gdh9KLD2Z9R1I+YaWJED/bCUG0tDN2jn37g0PoOUP
gunXGAtIU/H0MzuuhBsyEZhSjeoKhWJhpZOfnN34e/pe75h2NLROn/1rYp66MntD
FqO4KKdK3GbQpt/RTZrUfMbS9iThbb3v/wNE+WqPE6ZgeA+QoVgTcE9zxxhayiSm
y9Bia5qFhaGlFn1UQbV79PsjaTDLnQOYnISlG9CKkfR+6kxJpM2SDpKLws20PQuh
+B2ZXD3XQM0/CaUbLkAm5KB2ZUDEMEu4XMAHH0mJZ+0j/xo45va8AyglULAJiiUN
6KQOT7H45OkgAWu04N0GEpYOijCFz520GaIcjEjjvQoi8Sk79GSMr47FapRSvkvi
bQGrh1SKKKnaOTsI9jzZT24/00rZjXhx9ymbTDut+zVXEFF/tOkJqw05HJDdBH/q
2Zzj7JiaQ54pFdTfgqi1ByqmYZyqv/5ly6rdWG++0qVFd06gOQaCD3dEDNxveFB3
IxS2JS1VpAFETb7+acE195DPQFvdO+uI06VJAdglAsHmrOD5I+FUL136MH+kpIQT
VYXVSZ3pbjn9wxoTtoaV971KQ7lSgZUCZ2XqK0a5aJ6lXR+1gMoavLrqP/UGckc/
kcLkgtZVaZcmSIzIXOy7MavVNfAUslr00VUHHZqBdk9/mvcTYv6c4lggcpf8W2S9
24Vj2l4UpDN29Q4OMooNmU36rgiZe4stEOTSXw/yLCHPWSK1qnkc9KOgOMNTf/Wz
95HeBczYhWGZZ4G3xkPwgh6ekGQBKqHHlKRjfS7p5Cd7JjZKxg/CWle7nC5yS2x7
nBNp7IWP5jj77v1jGVVbDOWi7jR/8URwamQ+5XpGa/elZl0LZ3+ubZw1yDg4palI
yfwv50Jr0hxFhYdN0CfDkQR4iM6Ghz17PmREzIMn4Jw6YmYOaddm+YiR6S4y6ML9
x6UsnqBQgp75USD26sr1DGhT4MxMxHAaTW34qYydyy2EoW4KSeUuG/E+LQk9jOr+
vyIH5HNr05cHEAnefL4FZn4jNC3b9GTBWtxmRh32qAMQlqxqXABVaY9XsDeAx2Ta
1flfBrZ7uFqttxb5EE/ls2s73Te2A69Pehnjb/6FE58HNqvOX9GthdfAeC0uB7Ld
+xKbb0t3a9JZ15912aAHnujfDORqjPZVMIaG1ELt3+jsdN1bnubaTFCnG/vTRpQm
m6vk4m5bNnrN9mcdncrjMYm1QGSsJvi3mpaRnuR4lbNCygt5bw/ONAvIAYEojYGD
R7kPMpnwjenVYXK5CAzDzrj5l5qK2039ijf2lX15bd+P0b4W4gxUcmohrS+F6Sdy
NLtIqdGTE9Ts2RDK14EsTxRSVsLtVHaNkO63gLMKbKY20ccCNvIn+eWZ7UmNxFfw
42LzAz6eQf7MZyxRKAPtRsLP06JRFkTnxltCmK7E8tbBqky5OZ9OP0p84UY3nGfe
1/aqzywB7o+Ebns1/HPv+NQng5Ma0fl5fau3/4CVhd4hlrMiZ4Erh8NFYurh1kbF
y2QTQy+W2TdalosnAnndNxPemGCWbHL1yGIY3zDd9O/m4/41pwmyjSA+EqJn30g9
xFXrBkGmqiwmn5yiTGyJp572Pw9jcmabK0zsisxnPyVDaycfI+8QwMIen7x1MN86
+txsL4zyMzWBPDqvtQF39Z4EC2ehhwsqQWFyTN2ZeCvO6v39UznTZCvXGRScUeYi
uANmh3/DkUAOJhXbfoYyQoPkIAMml1l3hBrdvRz0AdzgPxpyKdLSTwcGeTJeb7WJ
yhMhdwten5nkUGeKdW8RnyiPKZ0cAKsb+Hj800TcC2OaNHLyCTeth3iBxqelt0SW
54haZ8H4wPpnVDubt/hz2RKcZwKFwTSi/ehuo8KhmYRHuUenCrY25KalZBKBzo6W
3jknPqG9Z9ucTSJrEwPuc+LlKuaAHAR9/VmkiZQm3+mN9X9myIK+/sRT7RqkHiKm
e/jUoHtJ3dZJbt9KR5ZsQyruoRnY0qwM7e5S37K0XP9n3Gi2rrbfRqQI/I4pUqEX
SFsUkcq641gZaw29XQZAnonKLuBGxddTxSD+jT85GnoqzMhDnIarSJ0lZBCzhgah
3bqcy9FIxLL2nRzuLpT5DnitfaJxAC2t9951mdCLr7wRzWGAKHFh8zoR/ayGadhf
iFl4QVw7VHO9F8ykboCO7Q4l4ho2qyylqO1Sco6HkybBxzA9kOReqjOeNXGRThha
4bg2Xhg5UMVbzQuxNMeA5lJFRXMt9yfpCyaNDWIVSDkxW3LEpsNteMQCNN55xREq
/GKDuFUXQbcDpdXL9fgTQXMJ+dm8RiKqovxEHVS17znzjLECnKGD2hfqeU2/Kfyy
0Hw6/2QUdZLP+JLQMD/nXcLmsO9HYMnDwwVcZUh+yXMcxV0iq16WvCoe9sPwtpqG
UjH4WO+i3/OZfV1ZEgBRz9iw8UIFoD1t1lfuIcrGSGhoquz9j7KfZ0v3YwX1Fcww
LarA6NjBJDjsUciqPl18F/HfSBTo1Ed8hvSqF9gWc94OgZqlKDeQngzYuqE5oIAJ
zl9p4OiJQkdaK05rREnJujbtKc3prv3E4lkr83RKoh+RsZcWiNilQU/ArGDi3JuP
vYu26kEnPrLiupQuFm6TwL2sjQFSa3XUy1+MoMyhcWWBE6tQ9DP1QoLrQjt83ZQK
NvVbn4UZblVcsXq8LZfp7cMzMQQXV6tx6RBLcKUeeT1r2kCQWtul+j8fB2wDjXPZ
88c3xosidgSLtPjj0YyVxSeQoCWGxnC2tPxyJokYD3Th4A50Al1MJhvVx2HnPvL3
BsXp/sA5hO6i1475otHTLJHmw5I2QbE5HyZ+inxpq0kPv/aSpNFZ6HfeLA7SNTaf
3Nz60vEbWGtZ5ko3T8JYz2A/jdPCGN092fq2k6sTUnnorGLdmXq44RedxFx2TfMP
4FQiUSk8RScSJwGpHwsUeYclIj3v5GAzbsCdaMXOkv8qMtCJl0nWq8KXPvYcPsxR
+eJKGYNY5fqlzs+l+2eE7C2KnRmeQCgySVvcYw0cLyl3UkRGVW2uUc+YcgK3dccj
6fqu42HYpewm402wAsSbKwCH6tKNlbyX2iLZhhLlDdCSD8O4bCCNarXZDv0NzilQ
sc7FPAZeWz4Ab67CgwDAsG4MjGD1imZ6u/ayVxwbH6/NBb8NV09kRek/bHIaRbqF
luZbwJ9Gd5P9ehnBUekccNOrkcvSFBx371Nl0mCAv/PD/VwY1S/yiAglxYX0Lwzy
aWqQZ0TfaCR+onhEPzkSyRCzQFY9FeDvUxYd0l+tds3GIO5pg802SiJO2ZqCXzxP
WxjeFrNSl1MB4yNFhM4hbbuWxbysaMKI7JnrnUYoee4AvnZUvqOHscLJkdtdSOhC
G/v61Y1gjMNE9OinXEIKdCa5BUVEh5mHB99g/lKYcRc8ONpV57bkuPbR+IfN5XfE
0/sKdC9jYmhC2QE4BgF9b14f/Z+YEs9xv6dyQOZqzS99D6W/gRiBdWG5YiL6fd7F
pYTMadVync3gBx2/zUuhlU7OXeqxnE25mTIixHlyAiic5tAlkmlwad5KEKjFib0C
pWvWpnXCrSyYL6bXeLq5Rk0UdcYPQpWoS1KIBzGHyt8fVVwlH8QNK2/h09U6dxFA
QyJDL3iT68KXswActOgXU9+vaDBG8YPGmLTCU32/ZAdLlhFHisy0PPp6zGNo8B/a
rbx9R7AkJIQZpl0Ae5WoSbI6DLNYpCVLmOjLXpjuFPvfO3UHzZG3sU/3HoUg/LhZ
rMWCFJAPfM7p/ObqoF9JQN8BD300i0/9CB/tcPMlGSqvPII08dPwYm4FufIdVZCK
Z0qTZQIPc5xWwVOZ2rrkY+B5NtGYjR8hWCgFcRGeLiwrCMVoKO36mfGdZ3VeobYc
4bBmzngL5rehvqqOaptDgljWpq7Vf2772aun8vF78B+AdeE7VfqG5I28XmYipSBh
SC+Y2bRoNYJrBXcMjGnducl+HbzFsqO7Vz8xYW8dA9rdTGPquZbg0P14QWjFoOJ6
kqgvZbW1m7QQc/dqWvi0tUsREP+UOoCMRixg3pUM+jkwtx3f4JR1Opm4jOG/xOJh
CoxRSDzhMDHLkKxrHpiQ7QCRqlPHCSlUyc6DVaunx/EKDSFnV+XHBPoLvkqcPSnu
JUglhoxnBGayFzniHDNuZ8YeNiT+gPZjt56d2OhZt8TLIIPpgwANY80aDfbclTeb
tWLI7iHpjR9bioQ857yU18OGeKNMD+fnytkcB/8sFR2UcUvQADE1TfSlwiI1RV05
dUOlFscVFWRc/Bm/LHYPdDltlvlIFbtVhfbZer8+8hvkwkR0/Uk9r9+Vf4YdJ1Wv
WMU79AM4bJR3YxqI6QDLxA+VUPPpjHeebgEDgEqnJKaJ48+lYBfBAvtJ0LkIABzj
PGAXTEBIbgosSTClNYLTJf+6oHs+s43lUsk1JdxcoPOGvf8FANN5D6nbyiFCECAB
jb2/DfYnveRa5IX5Uf1PLvHTmsyFtGXKUtCL1SnOzcI6jPELX3+ikrXmP6T/FnED
LDHCfAuMzVYzfW7G3ucIrUuQbllmyltCZrOmKsYiH9vZEMo8guYUx8wTdrlDSkH7
py9XJX1MJbFD2RSlsGgNBios4bMRiKRXppiN6dSqhEnw95UzZ7UK6gPp1sLrysBL
hKsLtO/K+jWSl+uqQx2ZuNyz3q4iNP7im5t6UnBcEk/3953293WgTLKuXYd4dO3v
xPKG0a9AEYjE0CRpwii0cnpOkKRbG6pmpRHK8VElnjs8P4qT4Npp17ILOiE+DdH+
6rKaRCY0rrG8qqI5iRhnkvZMvSOi8P7acsq9jq/BpPhuRiuI32tSOKPMubMvCq6v
201S+GgJO3/Rkcr6nk8xoHrOhSTA10bnpPbvUtvtTqKQjElO5tmUBvJajg6dMrmP
JF4wAafvB0Sn/RoY6evLXBpG+l2jyZHTYpvrIx4GCa2NY6JbnR+EDuGTXdhXHbrd
Dwog9RkIj8msYK0gDkObzex5ZeXhh8pxIhubXgDkcbnZEY22563UE6gLH4xIxbNZ
EX2PYEiYUVdp22l9qFXWhymMZaqP/i60IYUw5ca6RUt472NgwbDLu0CCD6slUuU9
eJPQIS/I528o+zDmabXtHYcrx1AyMvLuj3V05tUmbzHv7up/paCKyyNQY9cHxGNP
YsR1Tw8OHe69XnS1vxYrsUPnQOlsfUSNxjMnAzTz589phpNVDR4ZoPnldq2nd+CW
tWyZH7HLmtbZhIqr/xfTiu5n7y5C9+uCd77J5QO5mXvmPwZ+wvLMecjj93nmuzrd
jH1A/CLw3EQLkmWTthcJ57Sx4/l848n323OCszRM4zuuAUU0DgYRuOktvbfA0ZUx
j67hdR/HU2ONBgU95r8IusKtgQovvrCXKdJ6C1jOZqHxmaBJmkBn4xKJrhuZOp0M
0YZWi5UG09Tfk6oqq3L2Tvntboi/q1k16pdas1PFdjGYBRg7RkAibwi4EzFEcYQs
6t8eIKEU45cynsoXJCiUKiz8VaMm4/k1c/u033fdIHAqQzuG3OV69Rf0iffMbmlF
hyoK8cX87ygWo1LqccDMEtMoVycJThw8wgKk0KzYtDiPTp9UtJcQLGN2KA8WVERs
j7R/Gl+NnUKi9ry8xrMogBSvyInsAuBtJVhT4sl+44/84ZzqKYQ8mi67tpS0cY2h
vq/dgVe2GSLJPx2qg59f9jjhQizlHQ5BIh6HX07dRlsqDkaSDp5UFHMCmiJDu/MC
X9+WrYMIe1bQUYehRU4uNiNTc9M69W6/h6EOisMcdCPjBRN8RwR0HIkM1qotRVby
i95wEIugUPEGXZMucNgBhf6pU/EOmvD0+qDFI4eEkfa3fwUICqhsLWbL1Y274vtV
cs6ulR4zm7iay79D7hML/2UXOYlHtXJ5+x2hqkqSjxQjwRx1SbV9zdiCKJBJpgid
ZuaS+glBwxuge5CLzqDBs8SYDS/OPFu8be47lbitwxLieFEL8OX6Z+ZEzlKr6gup
bU1skxJiySVDUGEZ7jHwPM+r/oWjIWPlB6keDxg6a6Z566+uzsAqQdKl2aGZJW9j
O+SIp9c3V0LXRNRI1S99mQAnMs5z+eWZvhi/FhGaiRj8+lX1QYSZ/u6klTkJI4y7
HHKEeTsMnbZZVvJX+SX/sZuPF+hgsTBy75fzbWdZyvdhtjAipG/AqxGGGkyowA5T
ZA9MO0JEgdPukoYtiq8O654UzJ4UF1ooCl/bWZj50Fb1fi/IYyppEIJ3WjNXW0qx
EosRcWPtfShmIQ7hFV1EpSrbLeQxZqEXufEMgcRnHUzXbket8gF+IqwrEpx9sLMy
4/RCfhHCfqtxVRzfY+rtGXwCuxKoFSpKlN6MMS1z8hP+e7Tks/MkQcbfsX5/J+h7
6++w2p3gqiuAwY3a/QT0tgoC3bGlUzF3iPDY97/HKe3hbB9FEcugt1PRQh0h9mae
jtdOB7D3yu06IzU4dwZn+z59/Xn1bKptFANtP7zQoZKyppdRvHLWT8r9+n9AC7ct
YE7cf5Pgxgb+lSv57F3QcnVW9tFji7m3ZQE5ColICNXsjsXgjqsBftkiJR28G6IY
Bee8iiKd+xvYtZNhbU/LZ6EqSfJWcr1XA0o9j5451/HElCFpSc6SW19b+2fkOwxx
TxqkBvrjdmO6jR2h21qMuL5kNlbIsxWTKHHYS4bgUcVSyQ6zzWWB8xpSqfQk2QWG
kmBk9pcBBCCUCAPzxoAyoKwFL9cL7Z0xoF78HVfoefWYoJoC1fYrOCYtWNhBoG0B
pVs6S6ohLTSttGuBnkJnHygJ52EDnMgnqsX2ZpvoPk4AVADRbuOhULNWk3uW5tO7
XyHaefgEoG/FuB2XPCbJhy76nV3anxjIDCmUSTTCKMEp1Z8h4LF5ECI3n0I/pOku
o0qNP1YQcsGQ4LXrQnXn9rhHTM7dAomF67gK1hpTDS4RlMuirR/2ppCVOfd7L7iC
P9NfYTfLv34BTAx6dTD+DtZujdEJVwlEBLaGAmwH+5JZa4Qkj4LehLDohqHaJ1dg
EtmCV5s22+hTfRR9iSmJZN36kUtlRhl19tJ4rTlPqb9pm5yJE7px3D9eYlRU2Tcr
TgoojMZYF+DjJjhhsFKv2nFyMZ3F6xX7bPQ8iQBpyqW3I6pqR2hpm7LTtecr5js3
0900JZkf8AgPsbrRLRTafxZLTl2HHx64VcKz7PvA9kZNlPqP0z+bWb+7KeXS/6fg
KRw7U2adJLTTgpWDfHJY7c1cg639LFd7ceA5zVWtwVh86srEr7RjN9vdnTKftV1v
OmX38YsXH9G1nywp+FelmG3lJQ/KzuGdiWTUo0vpY2x7p5pZMId3w5lFrQy2xAQR
3hRDUGnEk4oNujeO6T+gw2tfzc/mGbbbaOUfq+jO2D9iDF5COVINmYmSqmI0rugX
k197N2oeCRlLBTsbi5DShFYI2ahF/u/b0hsy2jtSwNdx2QoNJcprgOk8U5FKGAtz
sV/b2lTtwQL2KPFT+wlLIoyZPhDyDm/teQltsFsn5dLb0YIReRw3uXYquX2ZB48k
eMYM6P0ED/TCWpMMnROiaPw8aLcLhPepK5sWdhWuEv0HtCZ9RXADmH3+O/JnWA/+
x3RqT0OfxkBBIy+DdKb/npu+0uj+LSzk/i2OPe5I4A3NrWouTia63wOfYuumz9nm
L57DiVZNZunCNrT7Kivt2vhmbKFIjIepA7BTlUl2/BrD6EUavXwWf/gdHKNjI53w
FacItbSRWSTI/iFcZ5+1pjW3wlAlpsHqnbEd7vbJShz3WBdEarSBXCOmqh/b0m0g
TUNOu8LFuDh3m5YV0VDpeLY4StDKUu3Q9OGFRPFaGRgIbDW3+Ukt4uKLQr1jIirw
r27GotrBF0xemnHKR0qlB5eQb95Ncm5I/r5P3EbkpyqNlyMuQr21TYzy2b8Qee/i
umnPd1icSLVVuZKkXF8LuwWpcL3ovVt5HOpiWJhJShNuzaVWdyR6xGim7mUSKr1L
xd8bMdS8u44dPWACBIAV84+n7R1VTUUbcf84mhEXKeV2hqJOlswx8tYQKKJtb2JX
OIpwkqeV6ZML6QbAyBpZ0mei8yI+Gg9T3kznZjQiZfo3a2TvJlFtdNfBZFqUYri7
ICrq31OJ7/jMEvz2ftxLJnvOCXquLYS9XCIFZyPEU+l3DAfFZb6XAIU5pDIA0piF
IzOFQuU0naQb+Q+0QAGELlcgeivmmGU48WLzY+GWD24aUsWMonygkHkN19I6T5+b
zYkssEORfq5iW4JpjUR6hZvApyChVHFShAMD8ZxOCTEFaS5Lmq1Fw4zAxgsXJz4j
QIMJ88bT9v89dGtUiQ4Cw4ls+FQFuJX2SuZ8LbawyhC92HUxM7NtYYvjGPB7EAfr
5IzSkaNRy73s0LfkQLKmWbwJDR63BBlT/EwTObhtO7JwXqlix01WmRLL2p2w9RHT
TTUvCdHotwaWn3MydzSRktX4cvnyErVc/BNlBXaF/RFKJV7fCt8SQiJ/tVB1ZAiB
xM/IICrvDT4lPhWv4QE1NaVo4TpoTsTr6qKEUkpBRzAg0opDhgaDlSMPcJB18/jK
1gksJLeMnHNFi9i/hAGd5ixUZzzdiHxfXVVpVuRusG8MdOjODw7JWAryjZjgrHJq
fIBQteHh+bHfMc5ZNe7pq7wZ69o5Op8VH8nXgi/+BO4UeaT9fechB9ieUGNOOE35
7za7IeMZGwG+8/BWROBeO9ltJZjHj5NZsxtitFzYNDnjB0bXiPRtdnvU9bHYuRS1
lztMB1Yn+X0IAM8Y5IXcxM3Tfy/hVSxKIsPoRnqFQbHy56ADAD0A3FTaHZjUZ2LA
Af9kW4lHl4o4rw+LbhyGGtQyqQnylvKlbcCrVq806Zi6QAxQa2MWFuWaF+KXRT4Z
lHo8vj3mrcFGOoCRWX1G+30+ObwsvlwBvyhHpgbHiEiAiCiiM80MRKpKrGxdx1Rf
fBOi3bS3hRon+HhIknEhi3kEVQL6znAkF+yLpArDDIcWOR7GYQ9+yjTdqEpm128o
at5r2QN/BjOhNYqidOdYYVtOj87GAzMPHwYzBDd8X+FRKGegQwcYCflIxlsUXMgq
JuYl+pS17K1YB9XgXWL2ICxRxNU2NQLon7vb5YfdGodE1JsZ2MjIi8UXGHzmVML7
0R1czA0ETKNazrPRgIaQrlvVinKbYLIiyf44HrHBmTAbhvsVuMd47YIiF5HOmfrX
3oVImXQv6ldZUdSXfdh8hNtbInudH1d5EFmkcp9dZE1ViNqTflfOPgQpwJME+bfV
7Ey3Sj4hbrOIs6Jr/tEFRaYbD7zXpM5HEc2hK2tSnjv65MD07noXgnJW6s/Ue4Vw
aESCUc42Rd/UZeNs+BKFYfrAAHPPxtnfIqNtxjFgJfK/CZoi/GBczIhRMNrlzjCj
EwKHbzE25rvkec+gG+52KLbAZAoPQB2OiPBeaymDryDYy6pXjGdzLKpLwgDha4YU
E/g4csvjbaMKL6Y0NB/21UxQyNCw0npjWETGR3Zv2JQ3YPIMR4Pff5WqsI/Fh74v
jg+f+a6lGZ4mgnczOzhaig==
`pragma protect end_protected
