// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lrWAIWYwFrnUe093tPiWZx1bFiLe2jgsfMch12VaQV8RQrbbb+PIdhkUoDpz2TTj
0Ebu4InuWbPekj/fnbxhX+dBB0XAqomTM8A2Jtdp3fkWmJIFmOxKsE5GyGJyD5SY
wuK9myg4KPQO3mF1+/drm50bW4nXXT6id1PFt0enfd8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9760)
vG4L8hkKvkhfQcQQuQPhJU6NwO8/PRcJZfzpsUFaqOPYAhDrejnd9hYlKCvFPJ4r
yDukVG3wWTcJDliKZ+nuA4BT9A+ytyKSgx948Lx8Q1Kmq26hnzhfsw4WXM36mK1t
Q6oMfgb+pm2yRq4eXuEGdG3Yt2XCVMhNnQnZe4nHOKcEzlegFEDJAwvwuCqVY7C9
vNX9yW0RvMv3qEq1j6keRdyOpqw6VWFEsoqixhTjU06SYBZECyPzLH7MEOvFnYk3
eSn+dO05cqqK1gxplem9+A2VH0zU1QOt48tQ1B3wi8KVrczZfHZSM2g6s5lwhdZn
ZE1fpE28wpnAQYqb86yHaqdqSF8NUVSdtJfQoOCtyb+f66Wkk/l4u72TJ8r9P1oY
1FKL+lPlK5NTrEDWr4mfbF5ipY3hFT13GoGPg6Kis/wtHVYlbivekLWhku5xxpHw
oIUcJ2hvKF6Ko8JXWA9T31phmTe7jJ/saqOkuJAiAm3qqqzZIn/YgOqFywJvn45f
0TbUoW4O5dWGkTef6rV8F8z4XzEPINabTrbJpYUQyo8XwX/v/hIfuZs3IuZFVhPp
BK+vF1OuOfQG+JNsyPogxSXmSZ7hA0N1YM4yzSeJ7mIBsEy58caox0KtKurI69tw
/y7uJ364Cb0xODeMWJfbJAqVY3KIPBd+uONyaFFrxs7BN+xGnuSKmB+nJFg+dAS+
wDZfpBQQrGevnSOaElUXnLFV60siu6wqSukp/jwBlIZovz9lPfVU4FNpc78UF223
WY6FH/JHzL5Quvh10X6RZlOznP5WY1lyNDx2acQCBH3PZu1nHLvzAeNgjWbbo3pV
vn4c9ndtcWbV+TLuwVlARq8WtFGopR+A3WeHxDA9OlyG+H4ZbIi0a/Y+VD71BJ9Q
g62o0oeaSBSLA2xAdc4ZSQ/QVgTkf7SNIJwRnNxjqapPMLoLWpmQPLXysPEIzo7p
1L7xS2gkvG/60mPG/0YPzhDkFSzOU1BCKi4KrbCx0tm825yiq+muU9LHvw3xvQ+y
1C1z2Yj4ZwI1oIixqVHyHHrrxdddy/BHGjH0xZuJUqQqBpnAbnp8atoPciMwtcXO
H8/NQDeAbfarxKb+wUAF2Agx5rl8kjDE6bDj1zMOKmvIIrOicWPWo/r3+qVip6wL
yX4qvNgholSR388enjnWtsQBP751GP6M/weRUiDkCQ1+mZvM5YIWP/WCEBQU1vNB
7Pxvbdxwe9IegTBVHg/9hGnRdFyJ8+WIIat7CtbxkZdy1UJTtDFjWPsvuBniyVNF
ovBVG95uZetPbHQVwhqCugCRdx5t78bDYBvbMpFIN2+/mX0cLo0/bUmzNAiCZMRx
NlDxbpC8/65tOp7do+iXFVXIwtSE3RBLZbGAvtVJoWicd4tWYIrC+/MLZvkknh6d
7NW7XxBwrSr0x6DuXbSbuw+9qrDiSlKNTkCMoY7Wez+h0uUIjZDwL29uNpgtRvXc
H2SnRsnts1noOa5Ejcl8/bE85tv5pEegBlFFei2CQjkXheyQ9USXQKpvxNnMEFgD
2NSs8K6WhOQag4wE+7KsXR8fB4RH7hcnfiFeNPCnz8PWLNF6Sa0w3Y44XUFFkm7M
VI6CiJDkEKdEMcHkmc+bAXx99rR8iJlFVntX6SJv9WayjYuqEJJKSEMM+2yRTMWr
n65+X3+UsjFFih6fk/M6N1jS35Syjt5ibnNxuePFdXRoMXEMpEBHlsEHS8woETI0
y7vURmMnfeSpyvLM9X2hT2P69YHYyR1c1+3jwJripv37l28b10KnKOACR4dr3oQY
phkCczza0/+G2c0vYfV6NxUiJ7NPK3ZKb2hZCnRT/yo6xVmnjSxFQn2Aaei0/OMo
+D/V6jQp2r7OxtyLpHThaEZQyZ07Rz9H7tHhqxl1ABlXLVt/qMsidg8mm5M44v2g
ThQP3cgdzPpiGhkCSs7DgIr7m/0jgmkV99h7un5//LXj+ca8Xkyb/tLSnYDkFPEh
RDzTy258kgDnX5M0DQn/lvhNqNxVtfwp6Dyu6gC4nNzuPdD60+BOCQiYinsZn3wC
e7sIovs0qNvkGC/63DLBz3lK3Fmk/wkZVwyHe/jAHySde+Yo0Cq1uIf+kijqjdii
yCO18UqlW6ATCg2fo7Lh4d8P+XNo77ja66Ifd0/PaR4pgVj/f6cHpL0PN6lrGEy1
BBrtnu7uT841pF1aZGoAiyK2717vjOIx9/y37Yf6yvnULNaZaQCR12I7vNovjaaM
qeVZggTs6YyEmQ7zEjoftYfdvMFRRSNfFuAthAZtM2uNlz6Rjr9qHLYo1+j2tk6G
3LemJ3T2U+cKPc4CQT9X4FzFczTzQU7cUYjE+hDABlPSzo+aydgyI70ADdAQQIpk
q0LQo6hTufmbIZTbIj4ZuhJPXYJtyYwSWVK0/VLGlFqLKoKYCPsvfoOcXpe8nd63
A/jXRc4P1FFhoe4QxtDFbN7VZz4AISfBczRPTRhN2mgG586Hf2GdWhYctNV365f/
ptNaaT+Hxw5v/gL2MeglNTrMSFvsuauDRnmGccOzfECgTz35vfFjBm2j+kPS2jDd
IJqbBO/KrqKvf5DkP/7XSzo1ZMRqUbNlTV6pXhdY+1YK2GKaZzrNC8zOm2BZcbE9
WHMoPLH30v3oiC3A1RdKyo2Ae4NTcq7xfXyO8m8nj3yNviT4RcPovdf8jh6YuVFQ
S649wfWmHnkelfYgEi+lJqucRzATLr4Y31+f+yHNirCOhs661zrsrV9Z5ZjtstZK
MOjd6MD7AC1xhuqOjUjuDIpqk/Taec7TnJJSTKpfVxVEx0Z3zA20ENKFMpxmTPvx
CbPixhGR/myEsrHo+1Zm35uCn1Xli3374Laj7JOiI9dDh5/yhhzE2gDBALf61gIs
zqV+z/4k3InULQnsEz2GgVlbCJymO2ZLnlCQUnOzSXqQ3bIzEl91q6NLGHzL5jRV
z8cpTH/dXyL8qkle7MdqUOoBp+yl7aAutjNJQnu9f2ICMbPTFMVg5Vz+q/TbOgKn
Xx2M7Sjk5bdtpB8md5dEXtEBX4e+y9V122rEXDzZRhOm4VHBYLxVfP+bwKuFe3VC
76mjpq00QTwHIrFsx0rc3ulCOkUswfPb7ZwGc82EPUMTTLAF7WB/xZireTnOxAMx
LJPgdi/9aG8oRJdpaixV6C0Rm/l0L0h6x+olWg56zTHDkNZQjHGl9LNvrF4WrEC2
YLVIXcYIVQoSH0kY4NZjUyRvYGCcUV8BzInG1+EEGVhYYsDp5pQ54blyKU1zGhZk
4Y/Y4P1oUshRCniy71wx0xBySkoA41ZRU8GGEXz7IRe3o47MAFRE2i+a++wznYqZ
384KO7yzV//Oi9skHejd5OKHvOtdZHeLms6dY5s4TuLhUO59H2Hwm6YW/p1m3wW0
YRQI55n+4ww6Escw3BdCJZmM5V1+/MRuEM/sooUDKFN0lIQtlEYzd2VvBHShydbj
fMsOmOcH49K5VBEa3/amKMVKFQeRZ1XbNe/OHqQhZIiVKydzOJKPvYzPiC611Z1H
nCNYwBlXPh4b1pN7WLIY2UhWp759WXmFQ2LhXc9K3XkfXR0uVfUBL7kQ1o/fOvbW
6ZrwG4k1JN1weTLTHFGd3uQVnCqt5dy3JcXt67wJkLLAhaH8QB8gl2jm7rSDDRnE
VhQqhoXVaXgsngHvve3HRgx+Sk8pvGYKzCFg6/4isW6DvGZ+qmCUySvd4svPR2iF
Q3wd/6p7FsigdRTQ+cal/npRmocmeQv1wk/Tr1tB9PL/824JuSQf3rvIRoMcTsWq
/Vg3pUBwDsiAHFHBCYw5HNpU0zHWRXNVFr2ucWTuAclmUhsDddEInZjtSTSlWlR+
hQotaqf5DdyJ0rumxQLBGbQ3uCsLVn6hNIBlVoqCedsMI8/ak1gCNGXi7nyVxVfg
ZQVPdxDmV4RW2QpC2t3SGzMkuUEDF45tly28rhDUb/vVMkti3pT1+71Mm5SofOzw
hmglLV5PeIgfLj6nlrGuu05eM8XCtlWLOEIskcKU/mR+X+TrcWZlrKDvKmAwduq9
rtEOvbVMVwSfaO07VrLGL1fL+ReyqEul4Gy8c0C0+Dw/Lie7Tcpoy9qf15HwKn6G
u+l6QR1yn+N3r5RNHr7yaXoKuMV26iS7284bKqnLoTgF+azr24GSHWw57qr6r8+R
JC0KnrmxzfbvoGbi91WAoGW8NRKnS0LPotOJiZX/jAB3AWXXdHYTaxxDPNQAs5oS
aJOXdx1TOzXD0vDefPEaE/gM+C40KqIMSe2KAH9y6vO9rxlXXlELOeKp0Zg0G8ty
eHxrRNgFKMebWdhAN1G9oAsjSsDstOps9bXop7FXWhx5kT0ZsCuPAg61WXhi155e
Ek/s2BncV3oCVtHSL8WzxHRxcvCnukpTrFGzrMWxzdXgPS6Vkzme6PklHtqG12dA
g7gLYPkpVmGeDYJqO33gYrQpNHKIpnoRu0yPABucSmT0kXVmmEiZlU29uM1zfkVz
bR1PRWxD63avNdENpFR5MXXrTbUj4SGgMs8oT2EAx1Y64zw369rnFnjgnB85IVJ6
StJaUAyzPugBL0k2gwJzA/fh2lTnegtPDN9LTjZvkzZFxHoV4klKerpkz/vkPu1Z
B/lOf8c4b6phPIZoxQZbyyuzMZ9oyAAAocCRfBfU25yKWZ9bf8pBtFt8d9WDXKU0
45PyEHFT7uAv/kY8MbWMR8xqdPsn0CL/AbHJMM6gCrxOYqb0pWnWRvMd58pDerJt
ksMXpiNWjG1P7dN695c1A0NNmLUUNebfkMZ0rb674kyOsWW8IzKvUxnGHv/fkxbe
jVvEU1DUrZi2AnZi+++o+Zp2nMSRUJN3s2ycxHZf3UyNRoWNnqzgvdYeUf6moO3L
bEXITjI1Ajp+YqrdHbGy0b78DQ18Ta8nqTiQeGWI8CbrFV1toRw5/UoqbvkK8CMu
aOxrLgD7dDSAJe7kpgtUGHDwCeVBCo7aOtY9UNt5xqq8pGvEXIyur6IvVt82Lg1v
rLELekPxf2wA7L90Zr4/arSxwRfmnIL4YNs4sw7u/Qlgl3y6rwhD+PigunP7od0S
EebVtZ9RkcXlq1na40lYDoU21mEqYIwr5mmFeObS0+a5orshK7wmPXNC/Ludlq7K
kIJkGB9XtqWtLfJ9Iq1iLAtfuqjSZD6Buh5tzZ8K5fyUe6zIZ6aKxnAsK8JHRBIV
i1k8s3DKqUZF5nso95NKuNmcJ5KLNPjoo4WGN1cCOuuofXJlKTJQya0MP7u+y6Ce
zUn7aNWluFXz4RKj2LyDFUOtjzuvaJb58FLk//ZwUuU0IXvX1MnRcN1it+JJl6F0
R7CDz7rajEBe+9qKKpPMb3ft2BL6At6kXfzgSRL/GZR6+gTjZNLHAHmU5FiANzqE
0jp6lF29JtoAdeeygfY2YoxFjtStfNTxGrltFHzjFAMMXqrjpDVMIm4IpAR8LoUd
bOQlnsCcGtAF17eRisxY7CTz4X5htwFMgMHo7/7ga+uBu1vZZcJ9HSuNHFinIrD4
4cJtDxi9r34sfexV8OLkvQRiJrDUdSatzGmqERetOg6tZHdlTo17QNGsOKcsXIzk
D0f4I+RFg0104q5fIYcYj+Tu5SDPPY+hZ+VnkeJq4Xy9SQWtmfWg34M1I2vqtz35
u3pYwodriwUcxtYxwQo8fljKiuMnurvkylyxQA1hXV/WatG0rWzqjmogIXEOkpei
qNJMz0qdQhFX63fYFF0yvTKhAGDpuRUZSxz8ICcsgiFX8eYF/dzTwB0RjTBIdO9k
Se0xM0V1qgL2DALaDMFPkp7Q7WdVu873shMYRrpaE0mM4yXtVvbAjxuhDAofGWLX
PYz18yfar7Pgf9ws90rNvz1XNds4FLU50pAtd+iVbFkFG+h/nhSaB5kpZ6YtcXNp
CHOT3bcAaKQJJy0yjmXyJWiD1NDcookF0E6YXxltEXzd1ew/FIbnWrvOHrrf0r7Z
ZAy0fr8El2XpIPLFhmc6dgTUrofoWdgRKZEZf4GOeTLojevXkeQ8jxflJnw2Ut6/
HRa9VZxhB6UjaL9UV92AcuqOmh9zGg8BTSdHVqaCx8qJlTWE7cVPq2OTrM01rcQl
xQF1+R+4iPIAlsqdHYKiXLLtqqd71Wxwk7xGrvl/RZGmRaAM13ZmUpJY2HvRYB1s
dGCiCyLC+tZh5C5HhWFMgqP6gAEmXAASOZNYWSGqtMuzshLAtSf/lioGu27BZ8qd
XLWyD+96vJ+O0jjWijV2SP6EI+yQIjfFpRT8jCvDgTXExgMx0K+oGh1XrVOlRLh6
J5IAn+4CyW+AJ+0/BXcGLu7kcZlBPeiDAdGz19J66Qo/nk1/q/wUaZu5enRFU0VA
umojf395x9c+a6kr5gy2CMDI3V9EsJ3uYUrWh7/F73/I9H5iDocc+0iPxeBrXVRH
SmcQ9fKRB84qFlF/WjOX1lT5cHa4Qbsu57RsRd29936Iort50OHZltlL9NOsH/xa
5rKjbCFg1bcUPCFsVUcqKbvS6pVfFJ0cgIOtcNe54MhqtZqVb+33mOKfI5jgz6dL
yQOoDBqyaO0QRKfI80NWhlWAv9VltEj8KsYp8kB5rsJJzj4VhgQzyW0qHqoWe8AS
ROTOx5EELYLb2mWXKebjQl01bQcL9m2CSMFZQxA6Pq7V3OFYiCT0zorHPQOIlkfB
x8jMm6Nt2c0HEo1/rEghJVrE8Ns/lYcun1ZFh+rq1m/mMTc61Wr8IhzmhSX4Jbuc
+LOg7o6QFE788ZL606DxvaIYVfXkYlmodedFQ8EgAmU6RWVuu+R0X2b5Gyujpujw
bMg0+yRSIAeLFeqLyoJVu6/1du2Nq5h5ltqn0eXT6eMADv5wYdZlIM4NQajJaqpu
08PXzIEJWO0cjKJV+n4wfRo2kxt8Gm5Zd0E24fZYCDx830Hajw+wK0nz2dmNUSHX
VV0uHJMFXWYR2HlEhK/baC5rH1aQjUA5BHn22zjBJQrmZb887b+3jm9yX+0FbYhp
d/AlGZ442nqW36V6q4GcpUuWLC8tX0VmooyJknuVmNi3tfKSs4j+/d47am40VMbz
ILMruDB9ePfnSay3lR3c0NKnYmdJLnqjbskhXOsSFLz9FcfKg3CM0SPjU5fRZ9nM
y1Kbs2xGAP46kbdpLP4nu+QMCiTBcCTL5xkFhz8TR9QQ08lSZT9ZTsPf+i/5zTh2
pQQCPWUDGPjc8hRwMwyhUhfs0/zixOs5uZ5nlDanKkDzTkw1atEGLMJVP7l6yjGD
u1Bvt1UFg9IfEcaW9obMy9UJjuB1VH8iWNKlglBXSmOCplFoul0XC+aXZt7Y1C9N
I/tzDfF4AYA6QfJOEBQQndVXlhwSBUFRZ/BZqIIKkJYa5+UtRbHL0JpQmFM3ATdr
xQNA6MDq34+mMTtl7cFHsCmwx/o8iEz+xPqORpV9i/t1/60Yh+9hCNuNO05RoWVp
gQX9sK7xB7edaQ6sadaPoha2dEYz9lGw+KsSG1GCzcXOtypiqcGBWFeHN+ThWvmr
yGuP71PhItaEyzgrigRj//v8/gf1sk07+kL6gciTLlpi0B1t87PjqWJfVvChb0m1
PZG9Ozqaly2a13YxGT+2zyep1UEQeQFg3G5L3Hp6yKeMFTD/8Ij7Gz66EVLg81QU
0qIIeEqYQU9CF5wjk6F8dZoH3CEhcuf2q8cxnU3jJYyxG8fSjh+QIYBH3szNUqca
aRMHOY4IUFIDgaGOBW1+WVVGy1SOAwVwTd0NAbGIMeEKess5vtG5jE7aPnXdBm/c
7JA+QuWaZP7+WBfWGRBQdJvau8zCE6A8Ft7k8/fJHz3rYI4Jghu8IQsR2dWK0uMO
iwxhHsQx6/2K8uI3z/2gBdP7hD6rL3TqM3BmAi6czNyT7PNdOF5O5ExnpqqhgJOW
U20d4gxpkjn/WP1uhEzOTYEa1Ryk7oqMFDKenjPqqh+Rbl9CXWIGWCSi37+b/+Dl
LCst62KJ+vfWFd7M7KloEQ53bR1AhaIe0pObAqbSs9xZ4GXo0WmrxMKCbZrPPEcW
jsNm80etZcPcw9hVmzc/WZ0vJnSfFJMZYMQCxY9ac7RH9sP2e7Jik3O6FNBP4uFm
1o3nsdge6y2vTsDY0eJDTwZbjcx5D/ntifc3iXAvo9bG2fhBdbc6ofbegpa6/h/x
geMoJZeZau7lygv5jbIfk4y+q8HSeHSwqq5J4osyLpLqNsHLifHnDmSco08wwUah
Nt/uDPBe4tvt1dUqHRjSunnjzSRVikpc6mecN+f6XpzFdmBehvOkYtT81YA0TP30
Ogc2nu5cMhasGROKGGhih1cscs1g8RCODHBFDFuvLnlZLDh8N3Wx7rW4+CjiLKGc
0sclx9z/wsvNV90V4uUPn8G84ZxyQa46iuOXGrXWj0+XQkBV9nPtlZqxN0mQGKTZ
F8JdIxCzLTkEb7OorQS+Lv4rGm7UEHq7ueGT8HxDk1lJ6U/d09GZ2OErmU6az4+N
sQ1kd4Gkv4wQhsxSx4A13OVyBUFKUGcUFY2bvLFGwfjPVatbwK0D8J+rE1pgMcAd
F3pCWqxJwiy1cD24BIjlpX7KxfqGkb9Yv0GfnPv9x5XRy3GrUeWV/oLaE9bmAnXQ
ixVcZvQ+9jdGSlEynyr8+iMS7QxWyakM0BZXKbgDNIr6WNd8dl2OpAkCgQyIsc5/
z6m760iw6k21n10KNw3NyxNdnLludizUXh4aA11ApKDGBp50YKqusKgzz1KlMDib
0DgI7lQUFPqyfgeePbZ7woMWerbLOuVrmLa2GccAiUBM3DoA5D5kN3gZ62bmEaG7
1720S9urTpIzDrR4Mi3Apj5+dH/rZ8MYB6mY362htAE51+TrgALa5xMWivjvfzwE
S95vJvVn4eTLkWHMX7b21gjl19utmZ0XSHTBlmBpVwdYFGelKeHBbfQqd6M64dfc
m4rTa3giZDRmH3ciH2BQ+u+NR61QXCc9HLEIqP+7ZlD0GGcvcDN/X+YJ0kLex7TC
9Pgs1CrBTgw0wkIi5KbKze5Ch2ZxItBnRCydcBdOc/+hpHnkUiZ0/O6xHaPhYOkN
Ik+ip5EJopiGR8N44rgLidwsYCspjVN/QA+5Klja5o70G3ctAWYYvpfKmzByWcfP
t10x1SkDySDKI/J3xuFsX2TIhJU+u1FDljKk1gxTAO2ipdIekwsL/AbDpeMLwKDk
bC4ZKHnA79QW324EyOUcnZ8W0mumAnOgTyUzNB/FDv6Hz9Kw3xvoca7HliOdALhY
5gzLKyggcUqVN2krpbm7CIqdES8zlifCagLwCo9KFEgtBJoNkkhEo5oku2mnP9jf
7DF8M8hoFZeeNyN/7xxOxn1lcVvUp7tNAoEuFv5enCDdCm6MK7LC3pXzbqVKKYOc
FyZdJwOHSJaSLFE7Tp31zDfR82nR9eD6qHvYeOEk4o5a7ZSWICRwaGJa4uuX4m6H
lbZrfSFIT6qkQdx7yzGOuWIOLdPV2wFCv0xhYpBGxb1PV+PgXpQ9vsTVLp8V3mIg
ShdxAajmeKQRqnwafPSRddKE9sGohFz10Aau0WQ0NAQ9WdnBtVXVhiVl1l5KPKoZ
f66QzpwEtRIIVghO4SXQqIImx56Ej7IUh0uNm37ORzsiO8vA/83n8sWJr3+C0Jg0
+KGAlnXdjdkpCq2Jno2cSw4dQ2PJgqhWiqAINFzw+FAkRdeYs43t7uII2U/AtSns
O5SmCO7TGfAaj7Ax5po2vJEcYcpwSZMikoDpUbJ7gpXgqdAFABpHS4gwIOxQ0Tmu
rp0OmDHDhWn1zPQluv575nCgtX3hG6sMEmZLS9IDNYvnS5lQPPp/Cm/mjclkurdL
MC/3mNNckFkQFtZO/ULcO2olER9P1dNVsgJpnVdJy3CihANgT9RVQurpqrVfj6PD
SuOlVDdDeMR5GWBZMj9Bks5y/YTLZ9s9lOaqSPAARhhzQnpHOzcllEHwn5MwwBNt
5GL0+tQZEFo9U2Z8F00eHxBX7NGnu5sMmGffeDlDgAiHVbpNSVUzNIfpW5BIt3Bn
v/6RuAAGyMeRv/PLuFMvX3zYTuT+EknPOL8kTn+h2khOTMB85CxD3REjEe1arquX
aLspVK+LZRNNxp+qo5h1rUGBas9tN3/oMRTdks2pez+tZq1JirPQYfcxw6U/ONRU
IPAGGUp14oMYotxSBuAzgx6i8Vwi9iRfNhLtPPLqUm3+aGJdx8sHux+uLcYIKE6H
o7GkqYkoSkl8XtMTM9MuGzNFR3pkc8Nk7nO4Cab/bw8+nyTWThcaDjqmpNt/0fbB
R7QenIbPb71H962H0od3Woj7HkfuZOPqEwBppY1XisdFP7vUlEdv2brxjTUBkboM
GNb/8rHB/jjNu2a7Bkp+2aadjVpuknL7Z6dWGC6vNrM+/NmH/bTuxnOjrrMbZYMI
D9ZIi2Cc9XPJyliG+GA7U2GxA9au1Y7jjn0cwkE8TKQfJBUd0q9h8wR/HetLsm1Q
GBJA13Y+zVtElRIzik1zE43GdEmctwhVPqnmKRCpFasp51laQaKO6u/zdAHVnGjM
aV2l0d0AbYZWMc+KvuPFLqE5unslYHpLf8uWzuAYgKSJs50/t3qaQ0C3pgAHxxBq
/0ysfSoOw8G9HMwe1bHrsUjfJtRImuRfO3K1EntR9UPAziCbY8K8vyzYrlsHhdg8
KrMOGHVDJdrmSigwVfD8TvvJiXn9yb/rHBah/dm5zLht+MkrR5mQU12su6FFbNHd
81Q0SNxCJRS05vDJvpjZXFzB4pdxQqngF02sxql4XOOejF40d3oomwwaVgCUscJL
anCifwXOxm2H7575zJuWMoaud8muTpBBh4zY+63h9YzBSAPR6I/E0DqwYOIJXX7p
idf0N/gvCqOTg0ESgRA1USyg3ufaiGk5PEEkusUK7PubJUvY5nIdAqW3urxEM1LA
K32pQOQkArE6byj0chNLgYu0Z43M2+39gOiswV40ZdWtJpZMe18DR3Rs0MNG76r3
9wgjRdL9YdRN3y1ssaCpqaRMXQ32b6Mcm/LWJwNBYGuLS77toeItj+wBh6nJMJ4G
vvf5XlG9hwu7g8Ms7shk2Kh6tJnMnMo5DkfrO8zobIOBEa5aSzhAf3aeOh/mQGCu
vb3uKGw5IdV35tZICdctHQT19Tjfg7C+JJKHDEa4IJG1K/zkb6qXSn2pifBe5njC
q/HrAxst2qs4TVMf2aDSC6rQr/mK01F+BjqNtHhTQtI4mGN89j7G8psVZtujKFtz
JclOc39Fn/5GK8891WHkYkMTCAgxJinJ2R18mNCdRWmiYSRzNn/lQltOrfARx8AW
CILva+ZUguYfPQ4r2hcHn4aeoMKBeaQRxGrkTBloprqDQM1hMXrdQsfSz1c3sAo+
e7NL/aBcmMdXcfU7w7ulc1mzL/AiNw8mdnZ7HR5VM8wIKdOnOqfqzAaGYzJqdKZ1
yowj+i4C7xXgEcOjfRvJ+lVr3xrA8cmDMdGE7gcX7bopatUhI+CSUWwXqT3pPq9G
xg93p/BlA4ZtB0mbtX4D1L3oeKg5Pnv8I55CAwc0KBrOSRIlSrsODgxsDeFy6yiU
vXQ/pSVPrYn2eOqFNJYWKtcB4B+/BziHBJ5mlEEjLa5FopsxKtaED1CdZkz6NdNt
YOiKL5fH3whKKIEKwaRBRbJimARfgFW8XYuWtAnEG2LKXHN795GHBYzCpeJRWPL4
eA0myMQNNsOtvjWqQd691vAEHxtDeBrNFv04wCUIzd6PLC7UfjyzA/qXcIVNUX6g
gksBSWmZ/KDk6VJjbSmJnTpbGvNwLog7xuvH3EaTkx/n8O44QuYutW1Ngv5Enq9s
p68J4iofl3dRY/usDCzOTC/KSJStXo/eSWyyE12FBF2LsZ4bQdeccxj2Be5QTqZB
O/G9w+ZHrOibzRCJxQgV5RYFZcYkZb4d5iHTWZIKJwwJjSJsDgp2viR5j34354y+
3eNYKfsywRHvzBcyOgCOVoQiAwAk1JoUNzwvxo/0a3PZjdXkiZ5bwnrTmWU0f4tB
o4bmSUQ9vtf+WmY5ZOuCpnA4X7Iui/4TKOsWRkywqLeVtV4TOpX8b7fpM4XHaNNT
mNDa/1HmD/nKDgXsrlPH5LbRxyLsxQ6YiYSVD1XlWk9UZX1dgLmCSoX/OYKtTiUp
RwaAr7+TJH6ZXdJ/KS90E/ammnKuMiagxLp4NxQ+t+rkaF175KoJeD3BnXXHG/Up
ZBL2yoWiDElBBCSxNZaOvtXFwRUzgv+vBKwQtW4RbI/WNVxdcU0CePqUCMsmVjB2
51a1IWAp7AcJhkAgnjWghg+2glwDJ8CMfQtUCktKM2hAVCrlPiyJtaB+NOQgTsFz
dyyTm7TTr2xZthgEfMMOgve5mPHB1SRhQ6xoldpOqa9W4N1A1lD95XvEI0QMXX6w
Txqj7QfNvTw4EtvQBQtJlT6B6AR/FNRvHXOQEBMzAQOuS2U4xo5CFj7aD1GzqZ1/
6lOfytS1B5gSufbh3g3fM3xMpw+bRwWDw7tl4HUn8DGkllSH3/fsXsHkCwLj1lYf
2OqFmN+mbQE94lnsobFy+C4VqprHqqg6stM8sqOQUl5dDxNguRhwBD7NRpZQ94ZT
4lj16weyrKXFet6/e1Zu9P0Qnxn4A+ZKcK3YKY1oMCmW6bS0gfjlO415wv0lQp91
5e14udHdtX6KAJCHclVghvvLA6OyuUgg6nJJl0J1E/BqOJFOmDO+iHXDHmIRGrQo
HKxmp3rtxckfYuQWUoIn5xQ1HqVND6F9rkILsoJD8SJkTjfupx0CEEOOfnzKQvoD
zhVQ2g0pEJs5ZUnTQ4tMvj8CyZpO/s9PRZKb5m/Xif/iDWzG7nQAeYS4IojKBh9z
4NNneyBc+1TBly0SrYmiYzatRvp2E3Gk6g49ABjJAJ2UlM05eqmQfzm0MEmWUnlH
MN0gXcZLn2pnmvE03oXTZQJm3RulEUa0N4kw79AH8+2cDJL7g3ZDzui4x33Vfq+I
X4XLZw45mv+6A/rP583baUrEMtVElqFblbP0xgZ+J3VBwQR1L83btCxHw4s15rgf
hO07vbqCm0GPKZiN7sBWuQ==
`pragma protect end_protected
