// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bZ3bALUAD4WNn6nulZjFd/uVHmJLTeyh1tlCoQazpseK2tlG+Vkr+nJrRxT7wFD4tiqT8m60Q4Mp
tE1H1WHStV5GxRSvA3VbeGrM+d3ROo9WFbO46xU9tQH+TFK4LcTYTv/CH/Lp1/1gkrPtCHGNlZr9
jhSKVRdY7Ix/9CWl5v508xUGJ1pMkbKwgm0XU2jRNOAjnYfTcKLYtIm5hYg1LWuSk4CTn7FqU9mH
LeClllukV4EwWC4pVKeBvZyigqN+TTzBRjoeXbAERz+h8yLUAn4YHlFRBaT5jujI+cm4GxJ/MMpJ
z73pmpie10rTUjwWFMzNdpctA4lyqH24up+h8w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
RUh810OhJMVOO8MUqP1yao1SlTQUCZPMh6SAO64mB4x5uelwMVP1Xm37osE8iuHYA00m2dnxGf1F
QHolA3X4Z5t6gzotk7qeBo6DCazHD/M48TS8nmp6n4oJG9bidFK4Dvb52d5NXf8iXXPqt/48dmcP
9fGnsx9B0391ZsOO9ClVNOwetRvc6aviaM7u0KNzv7p+ABDNKMPQa0gxiY7H73arpLoMGUqrbGOY
QjWJG39AdSY5YxHE8vwVSLVEZHWn6u7lL8Y8V+4+wQth98f7e92Etge+hgaZIStQQmOgW9RFDKJa
PPABBz3qS0Qfzjaj24KosK6sQ5oPif8PTmEI1Q/qiaAOtGvdDmJMMv1rQQ6V8FcrTUAL8tcaIq4m
jBzhIpGYbL1kEOD+uG+iPPCBZHZdbEhZZvJf43MfqQH3EoYmVA85vozhbu9TLMOJwtxAU8DzcfRS
uJf8rgO9mLTz3g6pEPwvpvvkwqk7OS49yRPpYyfdOPHWez8Pf0hrFQ+2wzXyd7uDrg7wXkQCtiAv
kcPq80BzhB2p6/tkcnuZ/A8LzSFIIOu7DffayJ6sj0PmR/dbrX7RCYfWOrFdwbwPfRyHDCtxeqM2
htxleNQx4dNcW9s8akU+n05sxmkAs3Jk0Tu6Rv4EKm+BVO+LY1aiLdXYtyxwKAsGR8K7m1e3zpSE
gTlGFafsZUbN6if6WOBP+mCKKRZvuxLTobkoxTBUnj6+yCouXT9ctYzLMch3p5P/TNS0W6dJrvoE
hxAXiNrrza6ICJRa2W9zv5jU049i8W8P4mrZtMSteONwQNVpr4wbESC87teaXsyN0HE0RB8/xroM
ekBHfcLmrAK8/5iffE6FmUqA6GR79xj9/gaYPDhO+v2wEn2grHCPdRX96IyvpRtXiQig9T35Y6BU
XkBabG7oKrN3gTPgBuTwTEVNT9iXP/CQVU6tLM5jUIBtyq22R45nQPFQTHVM4OkOISS6VpW74NKW
22GjvHr30c52DhwzbA7g77woDE7tqrefcnUVpwqnAww6KyH3hpOWrDQu8nMN9gNlSXpflPF5zT7V
LvmQDJlBBiUcQm5vmTOKi1ZNPbab1R01OH7vAwDWxG5q4afnet6EY07nMkpfbpz6g2KEMjbhWKfX
huGUs9iUGkN8+2EWLZW4sCPx1sGvPv6EsVLvS5GJPsWPGrG6czlgGGYsvTpPvzTVLinTA6VzFnyl
4SZpdw8XlI7kMMBt6AJ4+xcx5DJ+nJXoFr7gv0CEOKP1ufyYUshrKum4dLHONO8u5KPDzvik0Ihu
LgVy0Dd0lRM1a70aRnnyCdGeiJwmiA1KsEXEj6Q+vNTIiW8efsTDo4g4l5ZCTRZZJZnYnarWShWE
s9CkmR55HAwAu5Hq9U4LEFKmT7kPQ+B/UnCa8gkxjA9feDmI1v4KVRjavM+AMds060DFtD4ypXCS
w+fQuhGTs1avQZQ0syn7XmaB1kOkUo8l3Sj565Jj+DtxAqGPnSmXMkt15ahJDwNNNoYzmuQE+2OZ
JZDd2rhacSRgsIjn7TzhpNKMZqKsM5h9OIA/SwEtKMpP1HYOlu9LA9j1utYLlIJq38N0znFNYP1k
R0cYS1WkcGI43Qd1G0VmfjyuNBmeFA8u0ZSrk8OGmXEaMxMiSP1KRkhFgwvlwZXhYN7mQidsU3md
5kb18HwkZSHHL5tkJkTW7dNuUo+kNQXnMrhHOa18H9NIQ/pDqVKhHn5kL8Tm9eFELA9SSIOce7t0
T1dOEr7UOQ/I8NtN6YTNePf7Zz9gvP16yh4z3JNkegOnUAG3DioQ4tqbxxrX665yVt7pjpWnWj7L
O2aPxYiNhUp6dzZ3FCk4PNYZ4vSnb5HWGlFjUKPrVwlVQeX521WO9Q8stPDLdmavF+WDIxoWtLB/
RPAdllYdoCThxygNR60wQ8+k+KrJ/HVNGX03nf14vkFeeHQmx/+LRyhvmSgELjBs/LMRxlW/dTD4
itjej5KuRHlfgSKKePNHO+fNXZ8GC90AhzMS7jem4tl9jZxQmMLsNY70l2HxrSgDBvX0k8klmPd9
s6jkJZUxU4CLGMlMv1T4KAUMmaSFpYDdhb2HLBUUD0TOIKU2goAgA0/bVFx7uICmZ9u3b6Y96vyG
1aOagGoQv8matiYM3IH7fGAL7QxnpxMQ2HZm07mE6a42t2JcUD1qHdxqUUnwhePCK6D2+M8UBIop
Fy1gwgcOD2RZhpxFwYmf5+AHdU87RMDrEw7mmns5EqEpvKhc9MKW3JiFhYSG9tZzRf4IBdlaMTNd
dTqhqYsW8zfcTQ3OsZaPDzvY3BIQT7xOs15SbhtS9owWyxXW5zk0DiSj7YEg3Bxx8PPz/8iQyNyF
JRXCNMDjzM6SwwHG/l+7t8l57W+wYqtaU95A7RtZtb0cMa70iKV3jRh4eiVBBSgnHMzX2ddkvPZ5
TmOH36lX80xAgmplMNSETFoMhojBUqFRpzgA5laWGpgpY9OyUQuJWeUUyvIQdY1NK6n81DU4Oyan
L3r553QYG9Jl9NcvxmKenG0POGhJZ90JNdUdNsB1oTlGi5V6hAI7tN9+wsZJi8AEpq+H/R5mLZQ+
iywomTO/sSyjp+48zT2+b0YBqJIj3ygAv6UOhPSCzx6CWUepGTJWHYGYCzZiwzzcPKfwWqJLVv4m
1zMdeZtZnuZsRqpvt9/FQE0egV17AiGTkPcsFPUGZvMeieXG/79nzFfImqXwAidpgL0xXBd+H7+9
w3wGYDxLIFjOsoAEnbtL2C0RHs11Bm3Aef1jeo5VSvJvAw2/oYNa0iFCJ7nCP7mhJNQtTNqIqho2
YhHSPcrXfiMgjgLcbx/VC53XhWSpz5Tm4daz+MOCK1pT/Ge7YCQQtnssnRrRbyPNFtSDOfG3bNYg
tQ3JZX+bDCe3HkvEquXWOdk192oCbziJ79TIf7UnWLuuEK+I5MkfmYpFig/HoNwAQ7frIxBQN8WU
XU8tJcpOgHYpd8j5Ztw3ItsJYWS8j5Q7N6rZ31aYcHtgWL+6oX3WjKBdRrAJlxEvZ4h7AL6XDJsU
XrOyvEUKsbjHz5kSeknZxAiBOEmudRaeTJ6nh/hX26DDGNqgDbRLfYRkbfiOnzBs09Pvpxzyl9/y
VObKB7ORcMCtTk8YpIlpPMOMVcJN38f9gCxxMBYnx260PZT1FaHVwpkzoH359tObxL8NOSDriluv
TO4FRF04guSnZr0HljgVTbW2jn6yNu040S5QRh2Vma7zI0GBzmG2jYsvxhcwU2rQMMXtg6Vcf/Cz
KfWAwDxIgKJPyFpbk7OyMB9qZYVM3Fs2zCBLFJ3nAVuJLua+fT2phnkTztVLCmwvf0p5dT3xpK6V
eQOFQ5R0vTWvjdoe2sm1oqTqPRHhljC2IlMiJVCbQogprz7AqAnE9QtP0PGEP/aC2imVimCdFFQV
DjJjiw2HcgEBnBFCRu/bpXUrYdaGQBS7ZUQmTDDhY1weI/ROuut0Pusu8xots5qWSMFo17aOqx8S
Hdd8UpEQyTgR54o8sVTUm7/KYZL5+Us8sSAi7iIb1VrFq5vrs6roqMV9iilM8iePZZtFkCoJwSpS
0hHj75ksTXNUpeFiE1NRFgaEr7YhLtMC95RiXKHjTHV+w/iNPWM1F7VmvBjL+pSf3+BuIjgWy9dk
m7clpOH+SQIedMfyh/Z5ODic90LvgnIKKmsx86Gkn0OI8F0hleptvgXqarRQTBTh9Kz6CTyRaIQJ
Hj6Q3/vIW2bDNz9+/BQ5B6XwQ4J+yrxZDZ1MY5RJ7vcg4NeogAcYQ8K7vcofGGRnFYxWqP+vBoY0
a9145mC6kwRUz+a+Ep0d7llkLcQbIZ2CySHKcHD/3r8tXg0Bre4ht46BeD294QXKOSLFSw5uYDmE
ZqAm42FmgHnykUmgZVdmDw87ARuVMF/4ZbriTP6GNh2cRSAcVu2NzCd6wxOD0zFutXM+q96jtQdJ
GUIYQmaF6OrksdMt0KO4ElUjxLn5EApLGjrubRVH6aOApudb099rVHGwELwL+qr946OP/B7K4F2+
xYCv0gXL1XYnp5WEzxDMrtVFT44jp4vfeSQ+QSI+HkkVe4BauGXGUUQa/wT+PHVO2sMFo2qy7CQV
AjklQUf0YDIbFCjTIYy7HwWWLVOcQIUC8ojMbt/kQFgBgexqcYDZ8STT6+PtuottslykF8A2HsuR
IJHfW3RKOwKEPvyvebTTIkg6GNNiTL1ioNwMRVowpgTWTWVGrGDnm64/PlTRuada57Otdw/A2+uI
LJ/m0f9JIxANd/MecDJPuwhxF9e6UxdF0hhUP4fqQR76ax6npErxnkm1m8k0MtoBfeRqTJzJUtu1
7Qy8a98dlv5DfVaX4HCvdar5ZvSeUw4P8ErnR+m9JGUFVTmSkG0Od/ExApsQERfFxhllcUWjQU2j
dhXQFEgGhfpNFnxno+rB6jTkly9Hmd9GuxClWia49i/LiCAyw9GTeKP5dPrvphRJR64b0q+5kKr6
nSJbnLhH3I6R8oqNy3vYsRRn1Rkhb24dr1hOpCNprr3KGU12HBZYTFW39Ct4Ksyz+PHhGswc6G+B
FzKflDRtcp9xOArsP+uEIJHHv/ur1UT7ONNwjnCIRH3VR4ARnByvpH7S44cuWgSuGe6urQNaB9sJ
hJ+lrrJbPKv223HT9zi+mKEfhgo2mBP36iU1NF4aCCIpxtemI2d8dD6b6yaNNyP22odbGpb6j1k9
6OaZfAMrHLEMZ9OKzXOLMgDwvy2kskrNO8c1lhcHr6Vj3iPRemxzdZ0fadwL/8m6zGHP5wontfdE
wIFfDWTQS4c4/ixoBuSLuzC6nUbGy5IBe9h68ntoV9BwcjI5SRqeHoyMTfkZwW4Ong6Egp0sxPvX
maIYpHGcDpBMLMegEPt4CgPpO9eBcNELH/W6pYeYqyh4BOXzazszqcjOdobMDz7INDUwtoOU4gkd
or5/wNW4a9uzTp3rjcCMkY9LDlrtTxZAn3H5h2xW72N66tWei66zodvQXq4YZl2GzgL3DkhBr1Zn
hOZB2DDQ8+AmaUajDJ2/hR3vrP/1eBMEso6KKyVgGPf5cTAJWbtE7LQHz9E20NrgOfxJ7Cngy+cW
GwGvj7bsjMNaWWsW9TRIIFZ87ROWcxMQ02m+OlKd7ELi02aGjgmkawgeGyDMUK4MT9szyDoHnsZE
aPC8F5AoUMCdXzb6JV3tTx8/EteV4io8XwcHnmxEkjfjnFmTznnCmpwpElwAVVklqgwV9WL3Pldy
8HvPQSfZB3mUlwQyxZ3DuvINeYrEtqAVjpA1+kQmza72XkJ4ALu0UJ7/p8joJH/90dbihXO9edHf
kXuhiXZyArrcDqFiaPL7aJthHZtB5xF4GrZByl8ENJ/Be+nBD6O+MXIyVtEmnWfbgDEHsAHucEQo
oZ4bBubv6qx0uil7DQ7iNVFsZi9oLarU789CulHzCwV6UNZyZSqDvczJoqp+2e2EUoJVnUFUJh/w
1c3UCNo+jNs8GnyqrmugkiclabwU1iMX+f9aP/f/3QJhXFJhEVENMZEbBrC7yR+pbjYXmJ5cxLak
gGgEoRtWRMehhyfr+IEepyOk7lM+6xtIFmVPNYrySUGUqzU6gks9EiKBHbVLKDtBNHUZBytbsuwg
w2j/5Yh6izkMs0AdQHfwIvjZEh8ZZyt7ea1uW+xqEKxGF2GwDpKgekFQ4Gmvfji9RdRqFy6QGEKd
UA4AYysFlr8vsQp+QqgxD0Bv8ilVXKC9iyffLT4aYUJ55CcARkFkJmMbVNs7rchTtPlM7PJnJdME
oa68j00ItvCvILn4sDAdtbEDbGP1upBuoctjoiUUTnCTPB3fMKZmYJGQhVhH2gXNHsx6VwC7Fb+p
GeTbg5aHxz3BNfsSXXfwiQD25aoOF+hL6qBh3n7Xd4OY9GkSYCi9fBusSZYwEbJlpm6wTvkK+ngW
5vq8ptCMBat3NUjhVvXYiPJiH5OuquAwR3Yl/CORnYVYZTAQ3aUchlizcb7QgUrOrf86p4NqNVE+
o0byKt8KPwtIpVYhNQukGlfzqngSWUosv+ieog6YXWnaDKQlz9tqC+LP/WVa8opFWhhl5W153DgJ
9qAPVX3jPiNfMivHx7Qm+QkQUeyDdq/QOkAVzV3xZd6nCFDX4Fa/JGr5wDEa9sotDuuyZ41gh18i
ISg8cHEAi567o8W+yF+OyCaxa/MEx+q0NHXT4QdzTbD21H3gEfuvoXt3fo+xqtaxJaLEc5I7cUEp
DlDfMoScEzAviGnfL61s66eXcFPai4QI+20de2WV4rWglqPYaCDuymugunXD41FCoPCQnudVkA1y
zurSyz1RwkwWUelbmNVDeO+Sb3kHEQAJWjlAFXuMjvxVh+vAqaV6rotSi12uyzZub63X2vdYfYb+
ZgjO8hixpIRcspPIKBe3EnOjx/rHHKDaJCdVXHgrZz6t+IAy3knE8H1gECS98ZcejqU9jtZtAxEL
ztV2V7QLKNr7g4JfoQvV1KrYyFTjAcP8Wm2mkeMZyVUN8jsvT/NbevIdmee+2QjfXyE04I0RtLGb
3Cy7CHyqYiHXU3uUwHiUyG2cteVknfVTDm9Yik8Dd8XqjtAHzNxWSZJ59/601Ntt8XRCqMbALyar
5jSuGM+GlvjF4Y1zu7ir5w9tg91zjlB8YPKstFMtWiFNGNZXyeGYnJzYHqnSSJbYv4P1ntoc6qao
qNhTG9Cv3KYy52Q1X0YQO6NM+SxxkAnfPsdnG2ibYLC8xK+Q4zMcSRlXDLTBdK+U2HYDE3iJ5op6
WaDOgdAlKNjDXPM+pvpJjQeZT3TGP+ASjZ+cAHS7Wu7L/TWY1tELEp87YPROarm58dsKT50bM31f
oeVANpanqRz+Xq3qkzT5MGi2dmpHpMdmlYzc+l6Sg81+LlTImXeiXjhVKk/yID6oZL/tHPixXAO4
bwtzhuGxa/a+nJ7ZsUAwS+sc/ba3P5CeDGQbmjYfXCiGlbbHCqgUxFpqkpEFBC/YQgR4IrgNg9AL
wILCYs1mQ2NRl22baKdDl0pLuwccfpoLoQuIZQ4ERHGQUe6qndJZix7jgoAHickRn7gev8XSv+Kb
I3/AKelZnf1UPtZk7IhIpmOf6ldWWOhmylkbcVBL9wbOGQo/UDVEZAqIf+nS1Yx/wvWKB1CHh0JV
0RgxnsYb8/CowPPJfiOjHvtXrmYfDiYSWtH5qkOz1WWaGu9w2xLlDilsWUoXw0HBHhjetJp/i+q9
ZI9dUyiKuKj7w2pdUW83fi73EqApChnzTc4bg2FFmxsbXynFlUjXzbl/utpn7fKxD4x6j/oF1Ghi
KD+HnK118TnVRxiQFfltMm/WVSbz+Z+kL49PnfHTNN7Gc94oWu7Px7k6i3oxbhzRL5gk0izbpIVp
BVGQRF7zS2J6ZFveQJqLgAiJI+VD1S8HDqj7u5urgCDQNSwDPW/O9MRiKgvhdxe7YcH17U7QRBNA
rLkTRsbVPAXohVtZLKKgAN5hny/zQlUSW0PRt65yJwH/ROmURr90kRc+ihh3AMivXm8RCSyYGElc
3oTj8C34StpGmYyADv3FQcooftwSo2XpXDJ+BzpmQ6NwPcjNFBsEptS0gQCksUELut/UGuoY129s
9OjxUsHzqc2JJqgKxaFps6LULak1GfC5rkRDFuNNeVX7ZWESw+uuN00jlPJg3qFWMXfKJyErS5GG
jT2ZmwCdnxlCKm/4sm1/a33JeA0RJaS8deQN60ETuJPcNBNHOH5PQ1P2/LoXbnhP069DdRSyz/0a
EEaT8PQuXlH7SwQSA0UIMHqk5d5KpiKIhCClF8jgzMqX3RLtA13T6PznZMLPyQS6c6MYPFz+XLaE
//wnO041uCG8qW2RPdYgjUuQA6Re+EdT0QULQXVlz+0GpA2Eu7McGJvgB6tF4PJvvGWKAOJYa4YI
aRuN3115NAWrZ9R41XSJiM3kpQkZQjjPUkBoi0jHGMKeOj+JLl27MydzAwRgaSB4vpImC1M9T0xg
YcYkpeSM2tpm5PfTZk/2jdbqq8eC7/Gnpn7pESK4gF3+ImDDxzt30VbwUbcqJyvXtTjPGb82Qvt3
tdhNVzxenXB0n3Ik1ohs700fkbwLZiQj08Tzx7R9ax56iiQSbiRg+0izPynhFlNpDexstkH7bW2g
4+yp6uPPlLKSpo2/65udBk0clHE6PnrDc7UnmMxwG74MDh92QsqoWEAdc0WcRT47XXwH/fXd0YSl
p9VZN/i+Oc2TyfY854JkWDPRsa15Uu6i0/0tSu4IAGIe/fQYPAvac0zKW2GbbzGJTl0fRZx6TYER
yP0bMK25EgOv8R0sZ+nV2HHsVsCneTPB+454bzVvVSKPZbEK0HcrizD4+XFk+luRqyHsVsmvYumZ
JkKvl6r+XOV7QKjZTW4RRHrz4FcIo0t4hGKetSQZ+1qaD1+U6bPefsnoSlfz3SIMA/7UA691v2Fc
rP+hn8WdiNPKqHSMI6MUsCvLAIzBpTG0ZyWFmDvQnzSVzNk7Nsp14wWMjTEL6Z0uGZ9g7GUT8zda
e21wzzoE3DgrzEQgYlBKkAanImWonVvNKhLHPjkHZUdd+dOlgHoE5Y5IKrv65cZmZaPzks+x4ex/
OOmjxyEzYz5fBFcN1cTOjiGdri4H+OOKpHhb9M4nPY1HbxNKQqyXHrWLTND+XZxkfft4yWvPlJi/
GvM30c/4JNtX9voR5tqH2t7/SrqW1EqcORQR1fEuyDhYDeHcdRHWGF5zVAuh8NZvdlL/O1HLN7Bu
f2iFkKE5H9ny2kA6Z5d2oce4d9PYnLEBdRrD34RIg4ZQM3hmEQuQuBt3qSGNlCu6rrJk/TGgM4tq
HjHuqgmNsjD9U5+ky6vWRfaIAJuTLjLIgk3ih7iXkTHnfdXqpmYj4964QOT5H6abHGcl7LwzZP4o
w4D7618N5pYQFpv/w7Z3VdRZF+75vyq6JhYDxcLVcf/xiWON3zBBW+IVOaJRNq6nShQk33MuV98E
XdUus3DoCs/9msPjK7fK3b77y34eG8i5W5dEj8uxkF0XuTvx01YcKSGd7pBPXER7YfOU0TUwi06f
4yqjmhBHF4OMlMjEtvEE9vpofPIMZym2v/y1xXtANAa396ML05urb6YKzh5u1EhA9okwQvcphJkm
rWQs+AouFXXVAOlEZO3hMQZe/vPjZhzwfTNTJDCib/f0poSbHGQkuqLgN8jS/NDDGmO8yrI50f+B
CUpLOxpN/dR73PNj5OOfK2f+2pd4jXxN3G4OPu9wn1Ev7d9w00GqnRaQgD6zCeVrgTNx7VREdATb
WNhbE0Zujuwk7aDo9CIcp8PqGp6Kr+XlkO4r10yrdeBAAiUMxyQeASHW33wlDjaIVtCYUVEhtyjP
yMHWYt7Geqqb61wizLhtBtQX+X0UYXwUzpLa0OXWNU5eUjruldwM+kcM/TDfqgji/8D477BzKK4L
k8nBfYm2Dj/WAyusax2mgbiVIK0BhElx6y1JeL2K95vTp2DBWJfgf6HLtsipCR1bsnPpUff+My0i
oL5eFST37XZBTGTjJsQicr7CUPQJ4tOLiXukXWsPm2N7cwaUmWZ5r/XN+DqndVwYbNr8+3Tx9U1p
uvjttih7cFDAgku8jrCRfdIPfdcWG4l+7wKPmo2KOQy8IWA69CG3wmwCkeEWVwDQsPzzA9GKpoU7
1lA1BQuaQMe2iBnBMynqW5tuws8CnsP6vdbARn9D0dgPY/9fdJTPiO9nHyLAwWX6zYGg2hd7hbqB
uR5+tM/Tm+uY/bJT7rXL8AQIBSZaOqbw4etBr0h/+ohlFxhPWgaYHk37kzReLu/jT25JsdiWlHpH
zPFZ+RQzceVsThJPS5Y6HNoa0TlonQlYVcx9uCWZ0qVg5W1shQLjUnqZAZk7AO2/27EDx2jbkYQu
oyKP8zRlHzQ+Eg5V5brOEjtEHaljrImYzr00sX5vFhi8ImwsDxxc5joqtqI9Un+4hgupi+L2zglR
ZS1Ul2vgChfpkPh0Z/m1+9uMPeHocLw39GPn4sS5oBCcoOW4ORwm1F2PNc73eSmnnOgjv8VGF90i
u9x09PVkDzuUTX/ii+LnZPdHe/VC1muOr3AtRYm/IoQoA/I3HoZ2NF/bdTPNC4IotSkA3S4R7D7f
fA/dH7RnX8AhYQY7GXclhIsJctPCtN7YdlAW+09U0njS4W5064/VkCE+h4w10klEUJKpKsEiEDhE
7ynGyUDOa/Ti0gnzK8n4G6O3y4taev/SbGm95HwNHkWkeJExVYj/M2WF6Lc+YCoOn0bBUNc3CTKA
NQMMUl4usuNBA+UDeXxAxAniU9f3I3azVpAPf87rhSGeQBS32OFPbet/P3QuoSRtwP0iQYpX9K2w
hp9Xuo2X0jfvaCLwLOhyUcD8tikblnNceiwrteQUAzpu1BvumhlqHlocZpYVWxVDNirNtl27tFh6
Q5+WbMRViJFcnAbINezxeDtmM7NRKiRjzc57qDO50QJ0j4zne3GBMqEY1A0ZEumOfN2/HImWNqMp
PL0BRHb7lW6kqh08Bu3faIsseG31gz4MNCfulFwOFQSQQ6g/ZPEOM20RG+T1ANiPVOoRhSKbXB4S
Oa10Y7F+DwTuDbYeQTq6OPuKH9+FoVx7VkMf8Tldnc0S9ETnjZ5f/OKwnFMW0VzUasywcMAW+78p
0N4SkUh5SnJpq2yYQd2X83gp2WsrfpzQcJCb3gS0kRS4pOpgtpqdqrU+9Gw+2EP+ur5MYFfJBt30
aAoN0cicNJOhP3cN//1SRn8OLYPxZFnzi+TeDMwsor507OJIO4o82Yru0ur2B8W0Qw4GVhJDXgSK
mF+3o0L1pGNMEgFZqir2P26UkHlsdOix38zB3V181xNfnc+wTSsyTX7YcYQ/WnduwvGuMQM1S8cH
CdP06Ucf4onwXBE3kCiU/FSLzbZWfZ4WlMaFM5YZqhO/iPmEaiaZONMUAs7kxAhlvOSBFwoOFXH9
`pragma protect end_protected
