// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tT2pPnx5SIoltdu8+tUJ3cZjqvdRwwyF1JUrl6pPzpovm6gwodilOxVWBv+R7gnE
JykAuhgv+2aoqammU+k4zpdUDE6GTVgEexG4cyhPCC1jDvf3HkbxiThYhbjr309/
cr3YTmAxMTtIp69FdKNahehgdoNvGGqbAFVQgQe19rk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4720)
o8yITwyLnF3bw3YNb0VIyXQLM5WOEfQFHpNBEVZejx+nwEX6/9TmJ0WCBiAEymi0
t2p7k/npJgSDsSJcaz+tEPtmLidyoHn486klADLzlQPtz7ZQ5BGz//cSiC6hkcI7
AD+IGmw0ED96NLKUSCccat15QrK6hRa6wlJkHoZaU5gMLtgHs3nkKAtT3/0v4owe
b3jtwfqyWQH+QVJ+Zj1sO8MEjWUFEWeyqaJsRCIv95qxvgNuFmUSLASUMCLGNZT/
cq7NB/uODDCtlSqjsWrjPhPoxPLZ1qNXt7ilO7okvMi3aLmYyxxspJmdF2QiqnhB
axNgqXzZi0Jbo8pAwIp0g5CHUt/whbH+JaBKP0uU5IIfo99V5ynT6f509CsU+LGM
FPvJLrxOV/hzignOcvsYV0EeWwXLmqYIEBpv/gCFn9bTPp8BX08QPC6Qkxg2OoFD
gdOQLBIXwBgauOks8EKdXOxhlB9KUgVMGISTsR62E07ukyxeLgdDvzyncXFQ4cwb
UgwCWViSv5DZqJNZJ8fF9U6DGOPKC8C0aAnL/wzbmivxBoYpVr9B5BKgr/+ohXxr
Y9R++ndG1luONadMz69XhCHmTHRZjVIVycNEZRPjchnfXRyN5cV7Z1jwlYpIiXmJ
2pmwqEgIxYZH0Z/HWtCpi2mQtFT10okGo/11FxyTvKOjMjCHSPUFg86LvfhgbghZ
nQr/Rgc6SdjWKFkmkd5stmu6mHfM7tpfbq+EwxinoBNrp+o05pqEZ+JH7SuKHEPN
On6cfJCxpecs4vimtl8MzHucfBhDw9z5tRmSbCoHpQsTJA70bSSzFdsfUFqnbZd1
DMHWYIndnzWpQenpKWibUWe26t65Bv2Kq3X1G2scQ58d+G5W+19Dxe9HTbGB/d9C
qVJ7Oikw9gYLG/aiNO9r8W/yRoZLNoXGWQwNURpZloHjYWrsEJwGeODRJq8vsksF
Lg4HQ1MRdGPJZovgjkX4PGyh7EXDCoJN3YESAlSCgp1SQvDOKxjNjX3b12rBdXEx
QU/l+ydA18+qluUMVUpIMRDzcdNCSlXn5IfiVzxa5q09zSexZIp2l/Qr5pGx5QxC
P3w+d7926a+0sejQoODHyW2lvkMlRQpO4mK72+QtMD0ucAFSt4IOjoEjhhm1VPOe
rShiMu/ZT9g3hYfQqL8ML5ptGu+gJ7uBQVuUqpRac+TZHekT6M67yUHIEU3EyTTu
EwW7wuxNwfTzy/A17qu31lFkeotlnVFR7YLoBuFQoyQ3zSUsZ/3+XrP78RqV2HJ5
C4mykwh3Ypj1UbXwiaaiMROoLj9ViLmJQxoiKzMRlTKyeXdOeTAid8oIU9i41hmk
jVSAGUICpbdaaqzUJtE25SioAcXvZjvZmw5Qst5sMYvwqWx5KxaBFLZPBlt6UPdE
hITIQv4CJ0CVi34cgYv+d68Af867hiopVM/i5PAFvWPxh9ZJ3C3xRIx5NpvCMa06
ukAk8dhTgjBHYvMVPFweq8hPj2nEECwGOIIqRQCPEWymhdUCf/3OvFPTXuayJdHY
IZM5CRnWvG4SLY9oXYhLDkzaKp6QYfSCWborO5epEu2D6sCnC7s+M6hU/fPZlfcs
2UjAyTG2lpcuuuzUvimMAggWqD6hleO/375gj+A15kSUZfoRt8uYulb+ZenTXio4
gI4JFIubJx4IFPyvsXYdoKPkNTzPzbswlrOVMhKl0RV0ulc0eCAubxpdeMdoozg8
hgJYfNIUqVMp4ouTAxUHksQeSQw9Z1teo17mdp3Zy8qhnh76cunbxRKy2ZNd29Rj
cCCLsBi5S1eRKDAc2Yy1KX8fhf7sYnfeBjVmh2su0NBnSePidjSHYZqbbXPbkro8
i5TW2ZzUfjEe3elCZLCqorJ+VWQv8c6xdRTk7w+mT6e/FYSOn2lKdN2MlEqzN5C+
CXM2/kQLq+spCrW7xiTusPuHA6DMvrT7+P1QiakPbM3I35Sr+ygrB7pen1izOUJ/
NPy+FkkTi9o9feycd9lLE5y3V3joTVkdoavg80cTFESeBPg3XVcgyITsx2A5V9m/
d5nEyDDh8Y8qeTEfTO53nheX5dDHamt3f4JmlvjK0w3gWEHzRkBBgnymiYJfYeoV
hD2FUb2lOX+tnlESA63OodG03vuWZymShAUB7kgkpY1uliUZB9/me61Qyq4CMVjV
2OUjeBFa5PhT9Jee+EtBi72JYmBhFANSgIg791QpoZTQl4quRmzvZ8KtPYAzIAg0
2eK4kBPV5j5kRuQ/Kpqa/lh6AVwbDd97litYzlHp5Hv2y8GaxShKPsPZ06s6f51P
2Xcc+p4Ou1SDy+vJbyWxB0k/vkjyGuPkGntYsM7KqkeNBeTnrR0sjDnLzGJASybO
AmzJAf6+/YIFERhH0V6uLuzWzBTJuNgDblAyTf7w/ZNbegeGI85EMoiEB9WmEAd3
OiWb0rjmTGRm4C33wVjshl9UFgbiczo0rFJbzZHVDst7mFH8i3U0u9dxsWwiG0U4
oR9gtUP2kOIwTYmhsMTADqQwVRYbQIs1jJXWpHsZn7K4U5WmVSFPb4QtokF9sakp
dJpfwfRi5yeb5+YQsf/nWCz0vZO50T6xqN8Dv542CtZoIGQhGPPw5QzQY9fP+GZg
2TfcPe+1rH4DwfyT1u4GpJlLgGToaYQp/6f4Ed3qNTdNgGE4oZVGHvuLD7zl20rl
6wkrZyIwNxgu9U4YiNWYnBzZTzpdWWt6dYe9VJq1VdNDT8bhv9ucP69y//Pmtx1l
DWUrpMiL63udxrkMZ0J+/JRSR6EmbWTXEhiNqpgR+0nHeOCsRs3upF3TozhsbcAf
pVxDO8YAGHV6wu3r2/iTTxWv+4XbHBCCtM6Cao5meTr3TvltbzCRBBNV340Y8qVH
sFBS0/c6n7fvjT6GBy6jNLokujwcCbDU2/JculznMzCxvy/v6YMGk5wTOaLAM/ev
lsSM68ZUcA+mdyy/XWByoaT+1bc+dPYDvoYguEpou3IU2yzE6lsvzHm+wnlt3eQm
+GqNt5nB5HhZAG1skgrI7eTLlnDUiX9fU6Agcj5DSeRT9pA9sDc3lAOAFRfMolJF
dt4JpGG2w8x6tZ1rqJWufJG47Pa17W429mYIea28rUDIYlj0Z09QLwcXswtJ+/SA
a8UaL70mYrxI77WUHDKIzDbAZ7/bUuKK5Lmkeyw9Rf0O+ibzuHlkC8lyzml6iVON
nGQww1kwECLe+0GrUyLUk/g7X6ozEM8KXzuUv4YsolYvO+qD44nRc4MK3E6zcSDT
/dhPCBhTqk8v/idfVel5tw7v3IeNVSJfHHCpzCYluB6Kxc9jHIkCeAKaiSTeGFtK
zYIpNQYjcNvWuYTNQctjkGPLuf2NNRPpqS9Fv/NAtgkB/2pAHOLCcoXyjf8M8/rN
nsVPv9AVae0tmBRnsQS34Xy9HbbRJrdCurpP2aovLH4BgOpPQqZ9cpaxsGCrHYpX
IxiFP+Lu52rTWtatKRGlfRUkBXIc4R4WLID0q8y+f2c2K3AbGoj5EvAIDDaJMXdf
74pBa7tTHe2tf2M7hahirpuw8DSgKdjbBxO+ZXnsOOlrSQc919b4wsoFotUhFsKZ
57c/C99yDGsGDmfE+cFKp+7PEiOdLcGCeah2q/BUbZ9RqngrNqfRH0PpX1oXgax1
+eT+6TdTLK8Db/Ss3bygu2y5I/G399Je0r9ijL1Ki7Rts07lcZv136nI19hj7Yfk
vkbbB+AEbuc8A+6PwOy4UsuNmQ81UuUwVuIrqIJwG8nZWjD8Mo/9iCREn0iDs5tA
C2YDmQBEZGHPc/+yJxqemxoUBft7hb/cD351bTZ73tjuZTF7ZcIPH/thXDhjgjI4
HVsu/qr4woBWNUH3A0kEDUgZtH/i280S+jGA3UFVTu45xN2RfWPQKjPEnrJ6DtxJ
pDfs3QX1tXUtP/PILs/g/QAl+OYJWybLpVN/xxKFW5nOXyeEm4dS1eH/FIdD2kFa
e2TAHihnwin30VHmPIdvO0PX39aUlHQipMUJB5uJXFv8M0MqmTMaqfZZ2PZGkrwC
setS5/KZWawQkcOd2uOuLgSCG0sZcmHTfkbGENrWCFY+NpgHmGMEexMUjdUb5SNh
AtV7IgJSsbCFeJBuHvx0p0xqUC5XahG5kYi0t4K0a7YfrQc4AA9+hdQjUGkV7vYE
P93SoE//Bx7oqoLMZnQ5ACIdzVpybr7XHTDIkNZjUnmGNFPnA8ze7AQ6dOuv8pRs
cuxVNrpT2/7IKdNyFuNPrvfvHuiuBgIgvS/5M3pdTOzV7mOO0koS7gLMmj2zfzJ8
HcNP9QBhsXHTXyPHXZkacsTJyBGxE6FvLzpAnKZq5sp9Nw3sFJBt74UhXtZAnbB5
1lCmI4S+3TNyuqizkdv9yaTK5SiuDXmb/oOnJQ6evEtdf/ChJzR6EYXQr46MOBEB
a5If01vOYHFhNtpGRvWAQzDatBNu/VoQkSUVhUS+J2V5Fq1AuiNmw+340M2Eh+lZ
qMjJeUEcO8bnsv1JbRjlbs1UaTUMBw54pH71P9z2btxcs7LbAzrxJdKzYlYFRRWT
YJhbFkoonstBNJGSPJ5OVdNhKIFYuTFadVe1uQfvwvCj27i2ywS6Tf1R1GcUd8aH
Jp7rYIwmIzBV/26eCZeC1NFLcBMTgtO+4UVny4nI91CWO75i389ekHvGBsxjIR0e
8Sh5YIVmA4mbbpmDB8cc6pwapucQbZnU+Cyrgq/ElsvNh1g4KL67ZqQDcOuTW1fA
eN3xg4Szz7orCSGJYNgvVAuymFOt3mqSkP32hO4lIFjJlSGEPFIT/nuP8sqdczLY
B+ifYD3Evi4V4GYFPPGrfykyJl8TT5GhQ1+ZD7erU0f++DKxXX+Z6TQ0AEmPHPG8
2Ny4Zrq0+ek0VX2fFLMDlHmJ3plKSZjL5Emq8w17K3h0HJJXFBUrIhMBrIvl1Tr/
dZBpkw9hU+ysPLRIzen7cezZV5Rtew7imjFuXZudUT8FCmI15c7/KUh4tTCwKbpX
AzPlUZLTEXKogTID4yG9T+f6G3v8Ss4jLDLmZk2AA59fX72g8zC4j+q0OaqfJLuU
2WTUnS1qwrwjcoIDTKAwCu7RVcbDBpkVX2VUkX4f+Sg+WLhz5OWjQnaJ0r4L28ML
gMong8oiygYy9s4O073G6hLhULi7rM/p6S3ZUp5tmH066GkrVjTH/2Zu3rxebQ0C
EpoFC09+Z8sloIY/MVkvlVWPsObaVBL/2NquSm1CaMBhE9YJoM7Uu2VXCS1VBkcC
2q2Lk7UbXLD7tDfUZkAJvHQKeepl6ZQ7mQiIHEKi83xM8TwC5YPa6flLMW8ZftQz
Ku+ddShYcc4HTkxIgF4eQI4F3Wn3e70YIg8l+A5xNrDnQrRKluPE10Im2zHbL8yd
4TkhK3ePyONCFOaRFnYUXPAjIFC/tm1kfp7uxnH0AKGTEuybbBH5/2fe/O7X7uqY
bfHwT46rq/PWYpJwOuwTmIeD9ZVBfetW4wCUFjejHYqr6ScQ0VlwJoRD9/geexAO
C8NwTb9xFBQSP2lyXBUhJXKjmauHlsC00d3zsAHqTpvxXXPh1wpxLQDyqOP3LOLX
zapfejvxxCT5Sr3bHQzo2w1pJeTAFmynOOvTcvC3vdyPcN67PWt9RfuhmpClyEWD
EbO1qpgo7F3KeBHQkIXqdclMwLM/gwRRyMes6IzAe5oY+LjS8yaSm0fVHd1dkPBK
xA9RbBJm9lw1xAbPALKjWZU/uuHPrms4bs6aUISUUjvJy6Jpgxn1M2I/aWkZpMUe
14fBs5650rfO3027V94U/WeWMa9A0L5CF/i1887mIRDxHZpIn9hLr0eBVLYyf7kp
ZuhNB9I9VzIawhac67wkteBPg3sXZYaLYSQtfsf3FOxlvErt5rCVrF/SWngUe55c
HID0ZTBq7N5ghn2bAQHsiXgor4D53yaelnkT3sUQrElbrsEXmiH5ah4JeseYj9Pp
q4pFD0p23WP11bc4CL+g/vTCGJCmJ4gqh2o1CBgekS4vNy9cKJqZqMomVH8f9qIy
4GT5i+uWl53zxuwXNCMWcEXNIZxY3+yygrvixwSIQ4ftXIAk0tgAn7ADqQOtI7Wg
39wTNt9bItPooWoI9WCT5p7/pSkual0/vFJ6xiF0+7ZOYONdVYCi3ZPISmzd4A7w
1zRkRJog4nN6g6LFSpziWgIQK/WOt+DIBA6M5HPmRVzbOm0de3BUde0UOt8mxLTk
3zDz55kKkCZeWiAZoU7H/vRGvEWEFPjx+L0OlSQtzL4L9CEoxUwgJGVeS5aDcGfN
fYfYqmu6MpbXPd4VmY9kug==
`pragma protect end_protected
