// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kuU84W44yWZ9fqzyEWPiBHvuSbZte5BJ9rhSmUrgql4BWoJ20Ij0XPyT/Yi7siwp
tLqp92+K22kmq5QpBKusJDwpQTWxYlIeLAeabDtigGTtXcuyTQD1tpdy0PzChodg
alADfvhSovKq9TnkAJ6GvTo0ux5wlPz5p0PMQc4Ikus=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3152)
PIwfIve6jWmily3ZAAzksHfkPUOnRJ7AuXT2y8bTts2+/bM2UjAauhpppD74EKGf
IfNgtmyYBCpPz7kUdaccA2bwAMfmezX8R4oM/dlkIdL572sQBxhlnbEIkhoMgEjS
aGYOVWDDCTLEi9WBBF9Cqkw6fkENcQItZmpZ9/fOX6bcw1MKNMlJTjtkYZbF0y5m
yYTawnu4HFrghP2/YeUWcMrQwm9YrmLqE1DaYaUeVM+58wJkC+El3lPKm9McT6uZ
ZleorHxkSZfkqH3XWISjU4da6NQzgAfvPINMhh3Ro+BowLQyGUOI1Mo9h/CX/aOi
pCzk/A7Uq4yw32bSmQ9Y5hKTFUw8eACXUT6Vn1LTuXxyFUCSqnwLGDqVfQ28j+g/
4aLuuLpm1iuTHTrYXjna27pBLa5voOWyTK+LktEqR8DfiZ7Bwmg0+aePEWK9bz7V
q3nNfslL56ocMuI8Ke6xbp0f2tRXdu62VCAxCtO3T9BQA/sU6IiHBzU3HWrv0S2O
fnQQX6kfXhg8AHJufomWtlLvikSaPY+R3N++QMCQghMJ6LDqtVm0Xfwe2nloULKJ
plZEPTgZvkQ9r8pjqbUeO3cMdTp2BhH2fHk1OAvXbZ3GRz0yyi4Jd48h2juOWVVn
IWuJG0zkkG+FWbNOz3ybZBwbx/aBgQMmhqZ7Jm38GwiIAtpPjIE3M2u8dzxFL38Z
G0i92Ig388pml9vrot9OHJ0NhtjzDV1+fRJdx+uBaRLtVwezmRx2XwNMkihtH26T
Qwg6e/fq/SBpvk/InGHKj67U4L0665t4L3KyUSSXhzVKYTYinJJ3gZ5nbU8WLCwb
7T9jZ+t6/fXOgPJcoJ/gnz4/iu8mP99I+lDHpjIZ3M6YKdgX2VYrbuuwHRe/RM4s
2NBuhHC+6c2o2MMePk5MgktHo4d1+z9paW6emfdE1I6u85/+jmKRF1GJKi1TjlER
0sX9F6KOysimnXNbRvlAZIlqJQbmz0nD0Nf7Y6qCGIInU1EZVou0XwoU8cELHgiH
ytM8awxzZjK24ZD/JPxNZe+V50LBAQIRYKFNhssju8PkGarDqTRKNc/kzS4HcXXf
bfN/NOw+91z5+Yno9xqd4RrImd70vVnK6uquybSVoRwqPutM1wRceowcvdNXf3hQ
C2fmAj2XBszhWNVMdhL4EtQfOJCUBy7uUyaOQPYq1BvdeuJfqYLeNvKMfDr2ksoV
xAaUhWWy88nYlb0itStEP5/gV4xzneaUmC34tRsfodpicGbg+JAXLNqf9rTeExeL
/WWSUn8y2vz5vALtO3SZEEFz+rMzo9nzHX8e+XZ4cjKftV218a65R50GFriMdv4E
JkRKIohQhBDsWtNNCZhIPpPW3CFrZsUddpCDlxisahRQqcmZhDXRVu9kFmXxcrte
0UU28idCIwCS3KBR/5tuz933IT5bZw+UA0tq4S0IiqB7+Hr09JGNtazECa2w9+j4
GJ0vak2Pnr9xIivX8JAfZIKZgeS/kSu27tGk0KCBOS7YKUzqnmbZJr7H8i+NBGIw
R2O3dNROyex74mu87iL6B7zVysDJAkNr9/PMu8ScseEtuZ324QsPPSs25/Gzbh6r
5OJw1x7fAf41EM5Gd/jSpnZNBv0N5QVNBLXTkKO9v9V7Chc/79AS+Jutd2YutNAV
7X9vYmS01KuhbbdaK+y2W4rFr3TJu0CiYVoDKPlc+p7e10ELU5B4JoII2JkWAznU
6Px2DomEMZsNLoaqjYtwMAB0Su0asJUYc17rvReR1WZ7d2ILL89+6MAYKzy5vKS7
LS+TMq8hrMYQ0VlXRodFx42pqAwKgiWv131tVC6/GziOqe7vZVdME0mbSVKXV1cp
4d88gm7F6jRybssn4uOSmNf7yvF01KLU4WUn0nSxl7JvHo/7tfdYQgSU6Ym4n8fj
60XEHPf3OQeF398qB6wjAilkkpHYNBZJgS1k1McL08QJFU2+RLAFpCw2+ToJ9xgG
XSDcYBqZ+XJ07uMl2MgbcmQn/b3yKxj35ocgfQmfumMudKKWBmipGuayB42AMrOi
1bkQSTN0BnPehfc3TzIceDcDQgkecGZze/zCMvOIO3dTk1AxHgxo2UNd4quQXH1l
zPTKUOcQJK8kr8C379JPKdSwEAa1qRbWdKn5FMByO4+EYn7nFUB3FQ/XC66fTs9A
JBBZBjmH7bC1s4CHw6P58ILbEuZKczzP4ktCxfZEleboRFXmnpCBi3Qm9OhVyB57
IWa6EMEJFXlQDzMloUL9mPlV46Tz2wiVHNOMAGyEqjwWRIOM94wI9VfnGDN1n6t4
/fKd27MwIUEnjxTAyWA0QHhnx1fH7D7Q43P/ILHv8sxGIS+0j6pc0tDmYSJbty22
P3MlNmWql8Hv/BqCZJbVpqS7sdCtF/qFYam9AH8JKTPO26GSl1Y693+Dkiam8AAs
t2Vs5n1mXSq/IjSPeBqO48j49Y1K6TEJrfttM6JfpO0Q3Bk50k3YLblA9H2cDVwQ
j+J3yRaDvYbH8T9JCtiwagW08qKjxJQVzYX1Lz5w/y23Ry2WejVSRW+h6gEGqbvy
yPcjXFxQMrAB4K5ZdyemBlbZw1xCzMXK8hJguY6Dpy9ghW9MefRA8wKlSaZo8UTV
iIaBeChAAN9ZsS7Fy/FcC6Y4oiq4U78/dK2Up5gl0CxwAPmxXirwtZKzfY8Ncmza
41Udoe4eY+D8EKok8cEHmyFTRovVkDQnUFd9Z3rQltOAY+l3W0kzVZe/JA5xOHiZ
DaSIjyhy8DIX4RcgYfereXJLoAO54AAqb8F9Xn5imdGfOZzJk3ekIgksysK3Ljke
0WJfT0AuKOd2gTp4cXeHUPla2Bjl2h5CeGTLz7S1wk0Hq45wa54kOdqWTim8QpVx
K8TimSjUl3zEGGYwPurfJ1CXVt2SSJRNwzOvHo94+KXkPBg22uad7ZacDLsCIrkD
O31X7wZC0ylSskUY4DR1AwWALhUt8PRjEOTPrOUp0Bwn3BhejOtPwAbMn8+aQhpp
TIJjfm+Jewal/GbzCwUNjrNSixC1zmzd1dBavHLNU8KsOixFAKdd6b83qjqtX90I
d/YbH2AY8GGGPb4cBFWO1D6dAbM9OpeNS9T+NUc28xgjlh8lPQtkjCa6Eg6QRTRG
rz7avIB0pc0ZshHmctRT+IesLl0ruIMeK4ufRrbczUxvE65iM3ilFA3wI6t6JXny
F9+wg7Ep67WMkeLgtkkaIKxW0FxsrhKoMgLcQoXynkmUprvyuYx5IASAsV1HIjdA
EjN4/3ArrzhBvGueupBohDEBsb8kUvbUsZqTv24P70pplHf80u5AgLB8hKXcEjFe
R4ZTV/kNEe3DrA4+xLpGW8T3RfWxqTz9SpxsS7Xxa5eDkJ3gGYxrTeiW64bU7L0f
iRKM2EDBelFL7zEyT9aiCAMeAWiztGU49hmhPrpjHc1ZSkx8AojaDHWbZFVhcPQW
qqgoH2EQ5j+xcJEmJQgYIKps0uqxQGj9EDKHNGf+KukLYabNN3Is3hMV60n6Q5Wx
4airu2/4OyfuvNt7nc3G4syvVGzC8SLam7Q0Xpww2JFGt3icyDNdRNL08GgqlKft
S2tN9iMsIUnwh7ImchPgI2nyG3hVve9PP5I1/rS/HZ8K1Nt5TOQPHTfH+enipm9b
uBZkfhpSbsqZrftkeZkmAhB2O6lcZy+IWe6RemhxXsrZDKSfW00fjVivGAc3GCdm
dwJVcKw75635A1eS3DJ97kY6OsPg0pGYaRopSENSujjJt0gHpA50fplWZ+KYvsF0
J7psFkbW5U4nYIBBpTc77whqnN33Jfj3mP+Pv43YFK68m7bHYvRvg9l5UIuLPnej
4pO8gdogyh1xJxzN5Ebu6daplgglqB7U8BRXHwQc9LM7sE5PLjbCSUbHBZeFLbKZ
uw+rQUxDwQ6vyiywKRcuyEkvlYpEUl43J78e+XiE5vrQ1wulwJ4kH6JbVyXYUOPR
UaSAd0ruKI4jdqFBqPQe6MTeC0aNsCm92xKlolN5CT1YT45N2i82YY/YjU1AfugY
Wid4zucg2R6ynIbu5iWpx4wUCoazfSH6e4c4zukOAJXI2Fac63+GTA7NKjCfo91Y
ZGbI1SU5zl3oyvAGFt+JrXS8nZnrqP3lddo/tJ8ZC7QqS4XqHodHEuORXaSDtnXv
yEl8oM1p+P9wubdyeHS7BbSWbozSVPxbnuiq64TgK6k=
`pragma protect end_protected
