// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
X5tkLngpeONgfUZG4cbqahQLx89ZWPiP19nCdDGc6zzguHmb6pxVacEYyOhYwB6ror3HoiZu05oC
BzdLMP4lsEuhwPDjixExFa1C/2+dOMFqOVv12aPp2AwaQCVJEidTCjkqsz7BP80jiyQfpAcyGwS6
SA8XsIRofLnTetY3QOLtv9eADnL4nmg0BkgrXWKHldxMHiEHYI3t/kee1fDORfrQjExIBP5maXc3
brWGIlgsW23VCTNyg72Jaip5oYPj3KLXoAx9GO40ZMYWVWeVO5aLdq1BJsD0EGoF4ksSmDCdbyco
9qJrd4KzqLg7dbFWve/1EZ32XsdM4kaG41Kwow==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
kYGSel0ZAoNb0EkIcpOaQaLLFyFS/Xnc6q2W3Deuvrri8SaNOA7eshLOOcbduFMi+xEcdJAjIoCv
jjiL+Y5bFNlOFsY0k8VkOtxWdrWd480NN0p5mDiSqM3kVDmZzZgOJAsa8DBCLjadlXa0iEXImhDt
Gc/QtKvmlS6RaZf+Ax28Cacf0uotq6xyT8ck7VmvGy3vSwdaHlTWqPkequpibPY2Q6SkZ7oED5zr
N1CluuIXe936z7hcRIGVA+BIStg7XLah37q+ZzSuJ5ZKe+wc21w+6CaC6fdgXvWpWQ9t4wGW6O49
BLq79God+NJNJjEdFuSFINSAhBVOLLV2U0x1Y10MPB+r+YM9aECR6oNmtV79RR2b3See923Vk8H4
u3VSlx+VKWIvzuox348rZ8A+tSt+9tHkdsFkCfBE8aHMMShGm2kijD30l8BC5aTvIoiu2es+PheO
GQkQHhXWZXCo7LI1fa+dBtoVmlIr9InV1Va6x9iGa183R2cdLf7QaiaCyvGwpb1OJ5hCGYlNd1GA
D/6zsP1Aos6++v4yC3IxCePM84pPzxJEW7RCqhmIJ1ld7Ad5JqgIv96KohlbDWj5t2bKJr7RpG/m
tEabMx7Lzgr7svrmV3DbzbvY6AnGDhSJs/hykbCk6rwskZ7a4fC6E5DefCeej7TX4sdN0nYjpLIl
mAVejZSZaFNi35eWOlpk9CaiAk4shcXV2inR2+Q7YQZcyv2IWZIoUkPsJW9s/xwFAr6bXI06jA0o
L+QGfRXpJVJs5EiwYSxYoKyA9kEPkps/G6FAgxElnAhtQI8avoLPaLAlWbYy8RHPr+0G6mCsfEhh
pX459EYb+ii9xvUCMRr3axcX75GIo7JkJVYkPpT+GsyYxH6nVE7Sl43xEfkpWO1CwkMeqcbI8w6k
g4UmdjvwAW1kN5Sd+Ha+H1bTsl3BGIpjnTVCtDwTcvQc2ZVZX2oV5/3OZEuvmPcZvZW5rFYM3GFi
KaqWvKXL8T0HB5qrUKX7WwIqMK1L7siH8QVyyHkRv8LqzPixvfg1BN8jKHXEIpcy5pN3JSug6uj6
E2dQ2GxzQGX8hDooK6uQ8hdjxHGkok8nYQeSSRgPu1++KK8uJGOBUHA9qJDp4YmA3agY7+fg7q1J
Tasof5ahQEp1kaF43lmx10vImhfK8C1sNTHlVhY4RyUcwBCca1qpOt12VaveVDFb3KwsCfT5YIE3
ys/Ontvf/KHRhqs+LIIz+9YDRSMyfYk3bJivop6z8nf0rT9OYjZLoc2XOfcpz0YWJA3VgZyB8glz
8GQ21kfJDHO/lR3FIEnjfRmnCAMAlu97vAOUiAHCpHL+Zs22w6j4TS301K1GGhwSW7orwNb+5UIR
pKXPDzqJXi3GV/3b4wQiyI3WmmSQSjpV2at+khd0TnBAUyIwja3gY5kj3i2itPE7lAQQreuorGvl
PEQF6/Yw8rHIFwy6nzjEk0Kdi/tiOjpg85lz5UTfKtAGaGS+cIPVdoWRNqm8YrAXYbJiobZtjtSy
EzTIqhZl3zBMBpycADgcvF7Ymt5RpnKnUNMAXwWU4Wkc8wjsR1OSr9n7yY/Pl32xG7tjbpnKUu7G
mcYEZUQG09lmHEWoVUZAwSBlAaEUC66y0a5/4QsJC81fkYXGrl3doC6gAhZ2k8z5H8gGcR+Pos5J
VARru1+YgaMNMNXyutavzURNToGEI32qFfEAAPTfbw52AdEqkCO7mKeewDFM2S77jZ5l+iaeacKe
nn54TRREdClwyy+x6cVe2kfE3+InbK1V+r0+4bfA7fgw8cMiMmi7S+U9RmgqEH6A7ikct/llBUnQ
i3gtoX4FmBDNjzmyPcIIGqTmFPXCo4Lg70Gexk/bZsMaySBUzC21wg6Hqpm1GA7unEfL1a1pFi6R
OUfiybT7JIdW4hrnhZPJ1W7Bki/tGIPmqP/T7g2xsdlPo5UdIBkV+n/yefQSUgfRa5SrZq2LcnCa
X7gNKEpufM1mzH+RfCgLa/KAhaLesGKqb0cmBC0LvmDzTn8n9t0fRARmz7N5dni4Bu6fYxmqxDTA
E5bx7Gn8WjNn6oQUnQXDbVL6nA0MGhJ2ltSdTALQjqEv3EueAB0LypOnnbhxDLumSqMNkYfrdH0c
n9JoBrhR6DeY7AOHrhb0rTs/GpWG3gbMJFS+qXTeGicb7JRZfz20+AnG4OzmFv4ukkiKArCiPlGg
Nwmok8CQnONJpMcazqHmaluOo3FzJOoe9EgL+jOWKCJGvHFVYhkAGwsmuEvT1PJbQ4RZaeEFcWDB
b3/eAImBVeq2u8N+tQoZ38B3D/U3AD5gSmYoR8stLBuDbTe4xLNIgNOrHhseE4uJBw1deSAbFFBQ
0EJozCB+hgmND/OAgcquCnhhmS7jxJ1grG+9n+W5c8HuWdRHS+38tfWzPaUgF59Ilk//MOnDZiLs
wJCndCtgmwRgMvDF76CixQ1Pg75WYdisQA+9K3CH1fBMJmHsxHJ7C3Wss3IjU57tgXov1aKzQntC
n3hVZnISGCE9BghpsEf5arPy5OiTE1dfOO1tGvnxA/kjhhEFTqVYNbVkgd90zKT+KCKZQFOhD/ez
SQ8U0V3DcMbgYu3T8pw2qo7neDTpE9gz30BIqb+Gbi4aq6cUAgAvIPsK3JsOuKlBAZsIdwWUv5bb
DxutjkzkTZo9Q4CBJG+YyeU+U9uZrYlpu/Jv1Kv64tV2h7Wrr4pefvSM/HliJh3g/NdYKuJNAJ3u
myly2il7apLUFtpAp/Bz1J2FSZKWYVe7Llj1QoMvEkYLy/lCIyNAnwVOIw8EBBFZn1GeOQLCp4yv
VzGIU8KeYuD3YU2c5CBwu0M8oiqOYyjXk1GstX+IECNdzF62xTGslJJPp0/Y5unyuLjno+Sf8cJt
cUujbBzqtLMxRNGWWooKjm2Jpr3ombVMAvO/ybEYNjwNCQEpBqTGdJPx/D3SwpD1K6gBw1FS2RuC
Ut7wCKJX9U+Dzwz57E/fZJ7P0lgA1YU48LWx9YXSw0501AW5ltG7IP5lbn6CekOUYHR6OOZXqWRK
mW3uqM6nT9nQt9KdYkWGytx2Wl3G1ZwN5Lb4KqnXnuj2ERIielLWP0+1K0dQhbs8PnArS4Aif2UT
DMGWVZvoMqwXuPZy4Se4V9BRvq5xM4NqnaA1sDKpz8hhHh99bJlmQZ6CwchFiloQKZ+3Q1O/98RF
sx0ZJtNpwmR733nCkgzAuHNf9jytlCeYW5fvy9lGCd9JpiKQzRHTrWrrTNbAMvJJmPrnf3gNwcNe
P4Sl87wrxXwjnULg/5Wh5ydlZB9X1oKuB6sUZxuzJDxxG/6qLaVAeVkZN0TfqRmhajs5BjV2Z5wt
fFWho3gIklG+KFsPQvPJ+UpALTRioRzbFLhXlqlKw1qPiwOScouug/Xja9o5oVxK/vF3DsbFh1wY
bsTfzxOX5/Bg2RaasG+vYpUymE/dhNQClYS5KAGaycQMRjRFRLloEPRB4Z1QgDizlYU7UysX6v2u
64v/E5P+G0iyPiAjaTmTjg+JCOtFWAGNzDnNMa8gsBS4VpyGFt5Mc3p1JybgjVc0KcseLAc9l5+/
KQ0dcg1qbxsAek/3XR4dKtd6RxxwZwaA3hTSmd71jEPg8gwRWx+s+j2MjRtjC4z6izPbunRUa8PU
Z25NU5WsQfvhC/Jrd8V1yrNL9HydnXvkvgAyznikl/shNp8p8dfRjdiWN4VAHPTWgc4Ac5ANcvAz
Jm1fCDyuMO0LuUR5WHKRmWxTV9NLM0KJ6iJ9ndSbMVwsxUNFATr5C/xhbx4MBKVeexfLgaH6HUAO
XWislYxoRQR0boTg6wN7ubdHCCxzvBvwJ+PiInyNAbGZKQoUfXDSkC8wPW53BRC153Ta2ixKa5H5
C3LlNADm0tb23HqQGsGSU7WZ8EsUhCNmDjAP9SiLGYpTZ8B7JQQYxQaaD3n9vvRAjk7XiEdPWzA1
6U+0Nmi17Om/fQjw1JQSQ12U1oeiLIuB1iX7xsgo3GA4fN2riiSmhIZQtmSrx0wrMNhW7AkxJ8xf
LV7lRqUG5L3ivYM5XhXYXQy/o8E39SNXNcFPQKYHJOehgEzenrYDp6rGcbykLYajBdLJ1dFpSFaF
rEoBYTPofl3A6KLXEm4iJnsX8lJPatB3TGaO3P8w/aNiQ9oJW4iEfTwfeyIGxuyMSXoteRhCaobl
E9rDBpczNUwcUnAokNOdh1o/tMyy8Sj+N/b7xTrjIY/jt1tG7nGPvWl1CrSbib+CMVzIMkZe4o9M
23UWsRLSZeI/o7w4Z1sdoXdjTfu333kyAfs/MhSrS5HwcTw96ZVlRWBG0uX0+mYc+9qS+41aXQP7
ChIfQhd/0vAJw8iJCVX0/Cl8yEmAVr+lyWAcskIulsarLEBN/CxHqJ5rArJKvkdk+63GxWpv0cV/
PExtlZG46UeowIW2B/aP2bhPo9Yt7j0eB8ycNSLZ6j7Z05gYJc9uHsSVRE98qaARP61OKgboYD/J
Pko2AGGbokK7Bs9hfuEgURjg94YZ33Iw+H6UvksGahUkvrdihSGddQ/zQfqcWiXAZKGr9eIdGyW7
AuvPGKwQr8j6AE0+Bsm8CrW1TU1+xF3YqHD/vHGK0BkstkJt14kdW8eUdcVrDaNzATrxho/JvqwN
69yXKrcIclqIiWz6J2TjojiPc+jlkH7fx9Zn5tbxqOz1dw/y/IGBQKh8ZyXbGBBJVy1nHdG5wxtz
hvw8a1Ns09YG/jH5+ywMHh5sRbJWOvPcjfpXTH4V82PACGQjpA+pn/9g0JSqedovUixH3Slwjxhk
xQ5SSLzkKvjpbzUmEynyE9BN91BcSaRV3pPN13pcxkEbzybwmWnuVGuhQvh3gYUgOVjL+xnBKOGJ
i08/2mY/5EExr8uEnk6bfyi1bDebxSXqmKG8yd9gkPNSFEd2qTyQUo7PdxRtxeR6TPR9eRLdEAu7
NwB+t9JhMAtFM5T98cPSiEQ8nEEEWe1xLmKd1G/X+oWvvZVTzola9QAsVhzvGFz0U1+T29aVxFp5
ROVsjdoFrMvyrMrM/VgUj2VI4au+vrJu42pkPFBvTvqQbxwCxE2+3sujBv/4uncWwkdGzcIinF4g
Ex14OwtmTAUucRSlqv4h7ppTec35aWzH7m4zvOdVKERcTjCnx6SO3QrMz9uynqEmhrx5kZVCT8SM
M7FCjxlQx38aSsSy1RtELi83WO++P1ZoKDR9zl3pB/POb9fOmk46KweBcejHMx67KKtD5dtw5Qox
ttj3FLRY9kkyDW2G/cvPcScNHwqTEjPOE2iq4arVjDlKBrpwv9aDToqR2/6xD3wZk/L/c/hNDzkS
3mCZxQGxnqJrbkQrEfEQvvQle4NWxqD62sVZsWzY3plcqqoUrXcJMjmY09RiTOp81CX5Bw36DxGE
e2GKN6a3AHrNsWTcRKsEn+NQvS1mEu5ol0R8+RoaGXfJKHMp15i+ZlsJ9sWxgkEqJoLKZ9Z+S33y
r81jNIqSvQBtXCM58INHUTUNGkdzN8XVB/kF2+soppsnuQQWGkDOxFGB6V/ZkMSs9X3ohWXCeswY
C+OJrEUY9A9mLEpI+eUTJS2gxte2CfPToWDLzkkBHyzJ1qjwxFuHwX7wjbqBK7EVHZz1seSGV6cB
nGi2dVYu77DT3UVNjRwZfwpvENZfcoAfcKv89/AzAljUj19FA+JWqF5sAT3jlKHWjtWXaBSEnpQW
wU6s/UsiR2CGJRzZ/fNJLxTh4EwuFDYm/CASHoJgHjwdgTmgVVTTFBpH4J2Xel5Fv0eKijob3s1e
Y9F0glGMhFT62dyyBb4ovEYJH8uuna8doZ8L3o14d+JRhfJfRSk/HeiF/cNwh7zCK5Vfs362ieWc
qYYdDx8SFMwZm1hbFxW7tOgu7TsNDeAy7XfVPRJH1Db28knYiTuTF1uxcyz9k0jYcTRG6q+z/f2j
PlRkCfWP7RA1Jgq/1SyanWpsR3S0l0qU+RE9pCDdMuEPRzG4DwIky9RvT1LAlHvOUjpmO5KD9W+q
Wr0fKs3MqIvG9z63IEpbF0wRyd1L3g1ZPWpdSoi8uA5oaByqLLAFIBBQrr8jwMpcQFyWw5IPY06A
8dD+usLTNybVFEn08R3jnJA3vrKWoQkBfbUPlRaNJxSddjMne8MnTpRXsF++q06dnzvHt1AuziYs
IiNwPemyYVxTvR0+zh9x0ZcfO36QQRcB5I+ccF0omsSecHuBZnuY41X1gFCwbd/rTmPAr0k0agh0
Xsl7YrzAtJLEz9/BA93BMUZ/VKrs8AWZH7mFrWsguVMUuvmV1ywljBKDh/uUi8dkcskkMMKogR/A
VKx8KXHxdqLJC3v7ol1dI/i3AkKByR8dBpdzUOAnKCHhTOsiShe/uAXsJE5NlQmifeTl0Y+x/iKd
x4cHCVYrmGvpE05qX+NhjDMIEJThzf2LiMIBEWYqTkof7G0zIsHhsPUPHb5sqBQSDXGFaW5BBFmU
6+aa2pudJKywPDZfQKfoRq50X4tSZn/+B+cI+Rzs36qss6OfdCDKxiLmRJN3/uSkwYGfilGOcjA4
AkkFQCbYt9bSoZ/GE/laZU9Ugolwpn1O+axnjsWxZzK1CiK2wr5imjPENjBb5SE6sumIlsCnvGKJ
BZ/wkXbHeIn9OmhzXbJ5Ia9uqG1MRileoJBhhUPHOrsVh6IaV6OzIFCFvokP5SOjthGx7i9zbPk7
psa7Ujh7iJjh4xibpUXWoaTZS2203tOTc/dZMI91YPV3LWvDx5Cwv+1vdH1ilpvcJm7lL4/WCxub
5hkHwp3RxLBIQNLqPC2IB9uuo5ODZ1CbPTJDyqPp/Kb/hVahC2Js1YCZVKWNGG3b9+gVlRSMTHIH
KPSGYsMb/OogzkCoG49zuaJb9dlzIND3/A5ALw8p4WYCAExnw0tfyTxXRBNwyHxdyCZhEwPTaMyb
+Wkey3toXKDQ336F1Ed1KGFkArrlwAaidrAj82JfCJcWzGSYO82xDcZ1fc3iX5l73RcYLPHlHhNK
BeharHXPYHLPpjSHzcF+sAktmvUBYXNWgTdHkc8Szkv/5SjdCzYTYuXnGOfKrnmVr5Y5tsK0lJc9
BjN6Ik4Ng5p+4lV1zU16KVbUDPLzYZ+seBewq19JvtRRwhLgAXX2mhPYFBiyG4IYCv9De+OJmIMo
lNK4/hRetS2iFyiOfCdaGCKL1lHno9eBMHcxZiVwiWE3nSX0/0BbhMZUkeYrHhaWWn0bKS0SrtSx
nZbLhDC0Z9lbAS+NdW4e1taCrWu5GJpghE1roLdmoKXinTyOxPl1X6agiQTe11G40YSrd+rCTYiG
7FDbIOCkVOfsC/Bs/d3da4SVzkcP+KBUP3q3euCJOUCrhcFSzFy8Ckxv1zql1zmf3kOiU9S9JU47
HcEyPCBYufzaxc8ZOxQ4yuH6Bku2Cc1Ygq5ncYeHiOdkVZbPnigtbySFhgjadnGsJ2Xvidl/x3I7
NJyzCcTUwFOmA8MvMurG/+4z0VHxy9fIiPlmXHVR5yLjGEn+bli96G6dm+bM4PPXdD36ZSxS0y8S
/3cfbyeY1rrjAwxo1DeU77Gkf01f3HBg31iIjCAsIBe60vag0VCwKqDCeykTNbXyTelGIdoPlXmz
4SJK4Zsar/4tvBQJMS27R24tgIOr70Ue20/nUW/4RyM3GfcQ+5H+3VCSWdWI6RRBMJlr53oBo7cE
SLWtP8CivLcnozCRKOb0do1XMMjBc00KKAVHumC32MbO/S7pcQccQAVlDAIbNLBqdtygKGLg/t7h
hNPRF5LbkbQwc+rabafteQZ9+a0uz1eDGQf8uH753UfbnUa/OcHQYDq0uxbZD7iBPPqmxNcVmpl5
DolhFwIvXJ63Spo611KJKHDmTpiuTk9/sGOHXTheAgUdbSHeALYY0P1v0jfwRqhNJLaZROi4+5Y9
4c/FjEaDRbFIhbx/esTXeavbWCZeFb0bP8/FJCXTWXY5bPnVRssBgn93w7pIUxcu0MtGR7VaU+1/
4wwrErkvEcoSMuWKSxJIuPq9Y7JslZWHgmN9DMJLcgNikJpyTydiRIjogDKs6VsPgmrRcdtmBzD/
9QqdBnFXhUstTxFRA7NFAU32Gq2iL/h9loFgwy/8fGPJ+ggdDfBNZ6GAI78IEaTbwLsvy2GP273d
+W2BiyZeobyKBhHlgx+rDRGW2gV9+3i/z3LSNN3QQifRWu1IukWwsMP67T8e3GsFqzp9QwNRMD32
qE3i8y7uBjhgHq7pTp0JgVoigmKkoQUg3jkKAFqKBaI6+LKsYGnXC3XfnBpcVV+mMjCILuGmGnnV
4BUescfBaXbdImMFQpo/roV5k5FCsd7jOSSKVuljpIDOnmtgXYsa8MIUyOmpxJHyFX/Y6v8pj7Cn
ZVbK8FfFdNIX2piuLOWJpz0VCl7KRzB7VXGVr/E203YOsMmkbCWTPbvz0XgoZmjsFq5H3B0BVEzy
eZoUj5adVVGUbXAl9hXgDV42L2t4VRcCOJ1+BzDVU3rh+qNY0KTiTL35RIDglwxvPI/cLP1Y543A
oRSge4DtaQLlo44qiik0jbuQjToXaeECFW7RySjWd1bs05hIfOzsgMx07TY83fC939UUpfm9FsT3
njS6dHzDYOTRbtxTYA9TRyuZY0E03et+drJi+C6CxLe32DusYeLZUC9KKhhFerdqn8t73LAuBzui
UWGqycA0vaQY6bTeKnlqqMKKTYQ827n/Za197mNXJeOPQcbmKbuq1JvQTsGvmLz0Ouvyo6N2kcs0
eSzoW2hinnkezD6VI1m1XBRDg0u4Vh4VJZzk1JMCQ5QNM7l3G2aPnJom7/uOzthANKWvt07kyYGT
nlyCnJVttM1LR8K//u2Wd6bdDDodNZff31fNZaOdfmU8PP9lyygQM6VSQvn/xgTWdnuh5ZsJ0dEv
EFW0+Nu4XW+t5x39gA9D8HNvNiTv1a1u9Jgh6PRZlbLKsIYUW2wRquwlh/xnjCnMzTRdYx+SnwRk
2QcuQWuqpg1uXICrmGFvkjqDJ2n+H12eMJYJ9xCq2UadKx5ve6sq2RBdrc0MTaH9KmgiuOj0200t
84LelHNyj/YT/VlvVkOjcSIcrxZz2Eev78kNn2XcjfQkuNMzjwiL0MHqQ1/ihWHs69M5y+BfvFiI
RPyr8qqXnSfoRIfwMuc3+SpQrGfXmCZT/3nQTL4DqBi2UOgjiaYqwJMhNqGQot1m4LBGKOgP7qo6
j6NoT/yR5PJiqCF++sdYsYhJisndVBk3VMBLLsPROEs65lYHbCHef8bOCp9SAYejds50XXS76F9c
8roMJaju0OBxOXON6CK63rilOKWGm1XoMO0osBEVd0+uq4AqZApJ8+LqvyHqfURKAhKERYH7DqBC
i3qK96jQJw8tKOgybAaZFWxGZbD6dArts+Q0sm6TPfAJPOlELTo8afNmeIGo6FImxhvKeMJkYgC5
WmULxlIgPpJUv+RRg+1qRPXZMxb6SFZL/gfFASwhBEKHsgZS+N4hyQh4dwUrdwEwBoLhyz02ZjG3
tgW4wT4F4FTqyHgX5eGHY5bopaTv4FvsiB3QZ74I0ahybfiJA+/NA5rj7sfH/dTdvpcQ5WF/qQAT
kiDNbtEqJoxUYSndaHU+XqQhbWJnbXxsQ2tUhrR9qEAsXmw1aAkv766xXkjQGTixfA4CtIVrZl++
msgluOpGpaydjb47I54Xpf9hEKJGrh8aVMxaY0VAIlbjhnHrCrexDydk4Qt1GYF5em79dleCtXJz
8RFpfsy/Gl170qFCd8eyTFbeJWT6PTB+vCani3/LTJ+k3VsMHaozW/iSr7/5/7ZrnCv4kRozyGAb
YU4hpeWSFLqrv2OJaaY2stEgVlk3xKfsSyorT7ajtkUrBnLwRSNB9Um5U+hpOoeg4KLLAb+O5/Xq
mQ2YuhXyHRDSj3AzdQI5TOuoa+7BU32ZZS0HBCN8Bq5qigoAo9CZQP1SMZNDGI+ZgBu7+dh83nYL
aXp9xqtztZ3/RzoNK5qGyd73UJZLPRFUDqQGiUgulrSPOVieU8drqeSY3240+D9n34Gl4tnZ04Yv
wEsSvTXXDtrXWbOto9nSntPyaUcnpRj9YtNccfqB+5R/fGpkr3P72kgmOGpBMIzbJRVieJmvwAhR
EUt21haDUI0N9qufwZF1CKVyna1iN4QptgGTWd5pOnUHiFayOTUZ+tJoGQ/o7ojIARVeDYESEco0
8LHbkCv2PyjirHpFCqlGF4a2JpxvSEYB26uAsv6/owf0PmDEIuuYHMj5A8X271+PP9iFA7ahB03R
msHdjr8tzzPHWVrns5mePONXJNS6meue0JLDyilcwFlAk8kgz3IaK8LsUamnGM4aSIFt3IWuCXjB
qlWg/umP7VMhfIMZ71OLJOinvNPOCTO958S06rkOrj57dvIM6ANTVoWpHybOgQ9nnuFKAleu+bUJ
pKsIhIEn26NHQRiSyt1Rr+PXHnPMimL4a9LnUFFc9vg1Yd01OWnzlWHuZyY1iTjtx3ttbEHfziXt
l2QP0s1+uqW5rv5awCQHin4Xa/X6817bxcZ0c9d8IEWvmn8Q9J4njo3VuJVikWOKEFwloTi5UJ07
LGoZs4NcvwTH7jkSjKiaRr133L0x7Z0tU3s/tb+TNzJ28kdCeWYRtzsHKixLIAOGuAs6iJMF+r57
moKEr8G0qUNQgtzl6Z4svvfOEFVh3sCRYHVAd9V5MlofPHynPxN0Jn/d3vVmXJfioyNAUKNpEoUS
s3rCdZeU/DHkkgqOZrWDdaNPVjWiCJbIyJd71FxAHrW4cq8EFlVMS/7HeaqSOk7sSJexpp5VPLlL
dIsfRUEgjVbWPcCN/Fnl1l8bIwrddVnq6TvlnJWb59P3MG/q6XV3pTCfBbgjwF1SNG9q3TPRENpW
TQJMbmVORvYWyq19TyHjUtShRkQKq/PQxJ49VhkfPSAtKsHC2ksEablmzhgJNcLwYUbk25UHHYmo
A/vyV5399VktNIANJldQqeAC2bk+WsCH+fESrRzrsttIfzNSXZP6/Twn1773PR5wgPdmnb5Iy95P
YEJkJFZm6eSiHBHFXOyaWnwYsTWIbVdaHynEajIZJ9fNwJBTDjRYB5ee3/4KSeuu6wNWGh/wXhDG
2aSs7myh0l+XH0/71bNwSjpN0XkEyGkQpox1jExLfWx3mBHbB+qIQ89Zn/XplQMPdagYn8ht1RRZ
Bn96xK90IsW624qyr3VijGvMnGKJZJsfOPWJxT6uBmmXmjHu8vOwQR1tAG1PGPCR9UDD8MIU2Ucy
zrQN8MRGGC2yIccazJBeWQLI+7BDa8cFAQ+gr2dZDebnQyjM1khOK3kYtUhopILedh5mVOE9tMWd
ecoNEzioZPWOEp8UZ7FC0FdWMJfjmBhv4A43ip0R4P/GKbeVPGnXfgha1q2pZ/cKOFDx/ywS19EL
SFYxsXHXKdS5buK3Ibv8fTnAp3ShtJAbT/Qto1vAyglIim7q4zmIFPThCtEeE5WIx7K636i+NMyC
sQsiqHkK/Pui4phsfycWU2oMBZtvKQf7DlV5PAdt6GMltBaDZtKfKSCKTLhKjWwFQtuOUAb3v1zq
54hpO8+bdMoVtxgRSuRP/5l6th1aIqGjYUp2Kz0HXJ6JpDfS7CNh747GMeLuDMmEoU0vYITrUP6q
b2Bsk7dnBBCBzQ0fAZsxNhSTVczjNX0HGUj9WkM8nITNh3zNcOhaEj7ce2h4iQs6eo/Onk72sv75
sh+GLHyLl7xonpSMhBgwQ1aUk/alg/0stR0Hv7QIubOfIdPObVUDiudXzousItpNLAVp/iQ45kc8
gBpNOOwKcnGmtwGY7ZHwl/C3RE0aYytdQskQFyJ64LMz+WoF1fDSKdLo863HKG6wO+YJI+1JsmkI
1k4TnQ7uHMkeYAznbwltzsXRScw4nlxE+K2p85KzbtkD0wR5l/U9jcjAlk/uGOoDk75NJVkd/sln
vBuePj3UU/P7+VQS+j78cDtn1wLu0+o1VHXMxVEZrx2ONW7WkQPIbfVPd4NaHhP1yDfj6kVUfNjl
YLxICN/bIxlagP4wFPu479CXTsLJan7Df8M7Frm7TIVJaqLo5J4ME7JLkmgymP8+C8e6BLTgYyI7
/Fe3mRK5UvHe/6pTOKy3kGyJfuZd7DX+bZXQvfMEL2fs6KQwP5wNz8RIZiLEh7LKBy1RkZ3SyH8n
RNGxMS473+zU1umloaAITjM5NEPal5FzVn7fxgTv2tIx5yPLheMqfq1lAQ30Qn67u0k1uY4+EGR1
JrUNAFw6ZyuXKfu5slPAJw7f389FEVx5UClN6oBYejr/qV21tukOQb1edzBCLIzCSAg1O5eqFW+e
mMBvWKkCnl1/1X2U8TsXLcaJUx3/9lDEsu451Lu8F2aR45wTLwL9iBBkF8MBUN4TMKwuommwuOqX
gOFsjfLsV8m8o7KDproHpikE8Fq99GtU+Vz625WaFFGRmSaO6urcKnVEafTPoQeCyYGl0w77Id/S
2TUlw4b70VJ4yk5R9i/Og3y5kyLSHcvVTH9kB9x5jVvyDfkk8jIrKjid+UdMTtvYKa6zVfVSJlzY
joI/cTVDdHsfLeDevIgL8cNYx/d038iMf36JqHwPPywLKTI0xvaV78aa5SJLitUJVt6WP27Qo9UX
ESnNnRh6UlTHl4bBGHBq59zJBigBbhc0rGmHzZ4af7s6ln55skM5mt1ygVJVPw98OLoAIy9cLcQK
N1+ZkQGjsm1YxQh5mTl4CTTbSsWybllE9kDSGBpOLL0ndXowPhqyuluxs/mrFUl5tcD91G+PvrGQ
VDiLVcdsa/C0c0gvwn955d1j0GKQLiUv4ShQ0Q5QQoIdqwPV9kRV2XBLe4McvcvekoWVQhR5Pn5o
gkePl/+N9W4TxTVbNp3jnuPfTttEg3KGyfWj6ZqqYjFw5nJJelSoU4r9OgNYedhT4H+qFo/lPPdE
rkiIepFcP+C7j/pPngPwrFhDQncmVeEkGgxOUA4xafn5811ap6CiWE2WSfrR+vAlg1YcroUbufke
13jCGkQGC30XhoD3TtMfiKXyXmxyBZXnwEPfufmskq7ES1ROpUuZApfeMtgfO0SRhlh9oYVjNDL7
Qemhv/reTl7ZDzi7sfOkUZamJ63t9b3qKtx90WoMEduj/ZbKieJglBXd3D7wFVSjRI1sh7c+TvvN
R6zofknKlgNNBXXOVHadeVaIpsA71ZttupbcVOkl8yCAyFYkeakhjvbvKTcn2ZpOyaJxy1WeuNrV
BsWtrjje9F97jVBjHxcF5Z3ERT5D6RarTQNIyQUVic7/y8VWppbWU/6tNr6Mke+Jf+ZxdBme7+8b
9vy+Ea08K+KP6Ah4euZGCIxN5DldRf+Vg/lIdQdJ7vteU1XJgnnVnZGUVmPrJeJ7ljxV97GAg51Z
ylKhBkA5N0yRS5Y3hf5RAHwwEO1oaozZIYcasuLuFdVAmEZ29J8uX1rNzaAUPGk3OimGJk2VnfHH
su0xQx/pPPUlljDGWe1X2K4DmK4Ohe3/ITFAAnJdsKBn4r5d/UTCj569YStQKBoHYZgsORkE6avs
gH03cz0t2Sw35gPlJbOUXTsnPZHhsd8WJ9qWOTTTpwQ/4Q9699gTyNnZOsMJnVYcoHUaZFXIF+Bm
ff1OusrkebT7K8ZeRrYQadJQNX2b11H1xA6L2lnNtqHdA6f4UvEfSVTLENPYfJ2G+b4VxWPQHwXA
6SfH/pqTa2gKQaTB3MyFtfzjhxH/PVMsDWfi5zG9PDm11qnOiONNtk+due/uoTZZnZROz1c54+sd
dfutH6Kz+8Prw2zBJjDoUqTywoCx24roNult8YqZUoj4PTw6CGOMl3nFD+k6FeYOVi4QM+sdE2vY
hRe21aKTDNy3lcvo4wzIMDbXiTl90R2ZiesovvIu6m267c/DStZVc6LmQnscsK+MgN3JT8SdNDCI
izqbJUeTwZyO1Pw8CFZXDUPh7M6u2CAgWbnkE7D8Aqu+WMfSLMr8p9JefVxCAnqBiMCc2UNrfmsa
HuiyRGurtFmQvItdD19jdTqLVDnpnfd6BlcVAFYJbOdDqcM4qdMfJO1xG5eJAC5xtG6wabKs0EoZ
oZPotBor3IK8pn8xxHUCzZ/RuIiVMrbFtYuDqxLU+vIUZoYIdQFxwp0ZvKFMdzq7iqumibbJfT7m
e/IVU3JE6+H9n/haAEnapfZifV9AcL4u5BEAlSDZX30AdZHICbyNaeC5iLB4R8atHad8RoEjPe3o
b5eHNUBvsOkkwTJKn1opk6CJHokZp8EH291C3J46zFxcsWat3mcEa6qA3L2YOI2XX6Shs252LvK5
IQ9u12NRUBQVdGYkj7ud4KAbpeUQxV6+Z/LMMRbhAIvQTyEXfSURNH1jeTSPHLaSELZv1ZGZjx99
4A2eSfSj1cMBrECB27XPKVt7K0PbUj/uHmASyZWks8wPUTTViphEr2F6IkfZn2w+Yu/v92OhrN/8
+GZijgx+lPqJ5upLpqm9B6BHwKj4KPfPSMxFHIcYcdb9QnwHZ+e5TAh3zTxnodp0491Bf9TkQ4Ri
bgiT72vlx0CbW1OD89SBFeryAplaVSKIYXWAhwM6XCX08MU6oVnsbKCFfUBQJWRabe0i96wPQiak
N3unRtaE60enqzmbcyS8SVKMKEi1k3iS/jIVywhvVO3uBHRFEgM8Mj0IZP/DUctYxQ4Ux6kxK9xt
34EMe58GvQ6ATPoimMYydQRwgsOKJhsg2QTfH3UX+BcqSHxp7LCFmzuFHESAjVMQrQcFeNdlZtRR
bj7lN1V3PGZIYe5Mz+v13tN0RuokCMulUcbQGSkp9j9Y7CU4ZCzjaRJna1c/OpezcN1OO2xduKyb
IHCrwD2P5UmI138VJ8NwGEuCGOZiI6PFekg4qJsjC2BC4rE0LlDJFi6H66cklfTJYp5NISUUlz0r
fAe/Rne0daNeJUfpIux1GbPlE9opi6CE5vuMpoeu4V6SMh02Y3VPcU41rDYbd5Dp8w+8VNKRxXjq
Hzti/1QILWG9+zbuOnHq3Q1cW98kF1tzz6TTk2+JsHVz5SnylJGWKdhEqK5xWcOsf7T71j7MvVZy
kwZypR/7J4OPceOEjujS5GVa80iqAoa0OkWJ6SlZzx7dsUXPFHUnRbTTpMIQ6L64lMzITB58PWvI
fVYHa93tidjfSUaB7dQrJQSegra+1I6wKtT1ZwW6g2lDLI4nqr7kwx4h5EO7SOdxkRnzzT9IsxpN
3Cp2bgPiiOTpQmev2eilAK3fh3+LThhaKZf60/yGLFVeuTHy+lR+hdlcc9BW+hBPPyjvgTsZHLkU
h4s0O54NJr7qZvS9cqWmv52dj5oith7hzKuwK7bOdiRLfG6YZq+2FHXrBpvkua1GaMhRrIHBIfPO
Q72Udi6UxFyHD2wezYnDfcSqNXmSs1zP7yvynWYv6Vxo8reIizWZSo9WM0WWZTQrHuFCTzu6FY6e
SPSEsQbnJNsrWa6hjRdeFR4xCZwiDg7Pfr04BNYvBkaZX21hF/O/MHTQaZVKjsDbYQGdNt89XTXq
oBOrYywGWQJ0l/Rvnz9gPNLfw1eL/E/fGYsjycYzhKBPwSPh3PB9vf/nOa7DiVeVTrBUug==
`pragma protect end_protected
