// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OrUmfqZi6xYZyfqlYdRK0Pv8Np2MvMrj6RBCqhL34KNeF3YA39tCb2u9OsYl+Y/5
lNwFtiVVoQBA73cL6kcaJ4kuaSzR2Sct5VVqKzYVYpRq0tgcBrI1FOFS/VySFdpk
vI02Qm7Wo1jmwxNCm0GBHMVlbZ4WFLPOZslIDJCXbnQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10256)
+29lPFnWAznpKoHfTQWZD3HlwsnDL7LAxF+HEyntTKH0P1sGkKI8462gAybHP/Cw
4BgsBARawpA620CUHgsx4a1GjOJCNVUGB5i9QqCOjqUZgR1s6OKqMsjmsZwgsPo5
TVGbmn8fgVqRIznLORmoCUJW8ZTjQFGiMnfI6MoBb6KV7EiUna70LumrI/s2006e
Bdow7/9BXU7bO33BJRQmRATTyEYHmiBPnUDQtBaD4OxZljJ7f+YDwjL2nJu5bGgn
hqvL5VHPq1R0ujByxp9FopLXXKWhj3FFVjx8ZNAutDgdzYjM/5lG/+BsDvI1aOuC
Yt6xYhuCBKliLa4TrASxbvI4XzeJA6DPdTuMtGqsQ7xrDNkTeub6jq8joPqhriMQ
OdWmQ6B+jy4X+qDDdWpiGLiyOStpfBgMvGypKtjLenhahMb+ztXJyZ3KjNOoXg/j
gPYQ9aQRQ7qqCD2t0ys9pnbXUhvmHrsnKokAvh5jBUEmwRL1RKFDz/obkgcVmsJH
pk8JgMlcHO6dMC4B5rOAtqQOI3lHUTqRqDj3qvjvoXf1kIddHHJEw1bm+fUG9FQx
ZPypmcGvevwRCfYtNBUDzj3SjlfAs6uQKUYnJ8v94zkMvWeG8vM2lSuusoxVaCLu
jG7Ayr2IQezfZdhSXeuyuYDfUf6tQq7BWyKhMgOR2cCtFWp0SQn8eTMI8j8F0gG/
ZikZFCeGrL/gxPmb0H+0WgqPtA2okZKSVYeLkPBwdLeuZ/EyNxNqSdO6U2OlebIX
/rd5BOjt3Wlx63HTjNvRv+NUvP1FK5oVYo3w00wIK7fvzBnMg95hAsj6iKec6cqo
Atibew9ANd3ddI5ZVXSRlGQK6c1acE6wm6SaF/04DNsDRZBDSUJtr2aWReualWsd
09mVd9GmPvzctS4S3HxgWOe6tmDD/wUjpAsex4pCNx1pz0WLFS2EjdbK/c0d7uWC
NamRWHCQxLz3j6XKm5s4XOTJmwmXmnfcNvAH2E4bNXBADsYC9mf0dALFQgVhrQ7B
/7jIV9Qwx4MwBZmj+mi2JeqJ82X2ZgbNRN0X+3OjW5K1z4sIy70LUhlpfN/qfDVB
+aMiSvxfr7z6MAUZMJg7EjILdmh+fwueEQmRaTaO++j2a11FNPJ+Pibg4a2i1Wiq
iB7WE2cLt5OIuJnUgYoqmTWQsdLT0P5qwnUXhotiCX7ut/wK6cwuXwoaQwSkaj3Z
DCAeOaNiLYzGAVXPsZKTrCL3bVAf4zrv80EV7HXpmviQoOHWZYqxsKhhJXRT02kf
S13yFuOqMrWQNNxGPMEFDChAiDJQjy6YMjNDO/YTqoHnW4ENKO3uiOWAHG3nUl/M
wb8zPhq+BKfowXIa4yyZ9XU+0F5xW+Q5BkprpHbYWcExch6Q0fCeFki7deJDWRYr
3R5Y8WEssAVJAHFHklenmK48lCPzNAMsBNw0+VyGSpc/RvW2BnjpU36DtCKiT595
ibdbmIHw3j5Mb8wC6/aXKwNs/Wlk68/xUNTobTK45DWztSM/Ao5wYflPZ5W2cj+l
oWPVZ5VGkAQgRhcLrDxZ+upmRha1WLcAbiDD50zO6KCQuunmGappwghchj4cztni
OHt2x9p+1dLA8SKaVcbW5AZ466jtrvY5KV1JLjTEl9MAiq4hnDUBDng2W5acSFED
RiJich0cFDS6qrpLtDXlNWbAXjbPoQKHUj7RbroWsSeDmkkyJxCO3y/UpLwNJc7E
+xckWIN0ygMOe23ZD0Ogeb+GtayWx17+pYbTuhyF7nIHD04b+f6NRtsZB1o1xM5m
QjEl6YJQDbP18zBCrRlZI9q1eLpEWKeGvhQs3vZc2iWrs0f01kKqkoYaJl+RuZ6h
YGGAw1vyS8XEaOQa43qyO4alp401INoxhV7lo1XBs2ULVU93q1KwHLp58iYRr8Y2
xTLvI2AbrPZRTcRZK2adQg9jGD9YfK1nCrqtFYtW+dwgrmkaKd4dcCKopWvS6APJ
bI1sbW/EA/QmDWVtVbU10c6SGv/lD+0RXGFFLp1ViUrJmRnM0sVxMYxS8u6FhPCl
jAcTsIe6Umlznn+Nu/17VnXbQZ7tMKaUegWVDAqrlr2hGvQJ6jIJodLSZLhHU7mM
E1KQrmAdOTJCuHQv4+Plidgg54kMTixZ8tGPHHVv3mwJSBax5EqNS0uGkLQ3V3JI
Ejp8hLuv/6MxyCPi9WM7jSMwvexhfmD2Hp3nvOjo2W6Z7jXxZ5PIKAzIFmLyBSTJ
h1Y7YitDOUlrgL0McWi2F5IwPOlvMY2nEdU/d8arz7jlLCO1o32aa4vVkZmwSed5
saWzB2w9jSbjuHwv17SBIMSVXNrLNzU/jPVSWKSb5FHx2AfklROEhZeXszo3JPBu
IGotO3i/I2Bfzod39Jd8lNg21/PasF5nGpls90HG4Y+z5kUgd6bkQNdefAkXBrzw
jHhRortW2aXa2vJN5ho6D1NfMBbGS6wG6ryCgQM+5gwn4PCh/7YiZT04PExt39Ju
CK5t6+gQWKQKg8LsKJ+KYnJZm4xIp1xO99vdPtquvtC0o2qGTBwK5d80LqsnGLxq
gfTE8s3/Gg8q44VdDmKWpiF/HR5JU/y9WSAEBfW56ugD2UXRY0MTS4TYa2ljwLuw
rpk+KkLy8xUffW92bUfbRwi/vb4BnVfiFeUq7MGahKLrRp5s51+WobM2AYjAkEqX
j5UpJ5BkPRUtMKW4qTHjlNUU+80qzadbNmihbBDxMUlT6RdKwKrSQXT8Sx0msXht
BiGToocAWElz7CW4ueFJsxDIRUgtH9xZ2+lVDwkBcetNtWWyvlv0STFUwKz1rYh9
ZpppTrgEAd/9jQd55YUhDJ9nnWthJII8vtQijwZLymnBkiIMWfywglnRQkrMnpzY
ky4l1gXUNL6XNIlNGf7N4m9MPmHL4jadBMvADG7TnysUaLPL4So33uJWiti7LoZU
La1NtjbnFeDMdrPTQHGZm56QYSlA1l2OvBp5U74ZeA8yDqQQZ1rrvq/kf8k1q0Fk
h3h39H1zoHq4In6UG4NJ/6rDQrfv1E/GK/ikeuH5by4YrcQdwEXkND7dSDZ7eR52
smJiAlQlXsbvvtmYsRucCKB6NODuHQrK9fRd+9x2UyGrpnnyFgtXI/Ub4J7asP1T
WB1eWxdd1qFH5/cgt97DGduKB117jIi8RFdZNwc3QbMM7399sYmE+Bh/aDCDlnsy
eRYP8ijLxTX+oCfk101b6GQKx6WMPL3L8AqmN9I0VSL+oVI+mFQoFzgTT8ZSz0Of
hwrlPIJLcZcqf6DYzwNXxkwTTBlgfXfH0CTq49QYRdDcRjXbg0BnKWytO4xcOepW
3Oth3Np9G8D1D1ScDDaPT3A/DaWPSewmRRHWruK3dBsQV3MjnVM81efJbm4uaLUZ
rXZ1KE0Xn/56XJcVc/cBPjB21mPbqFeKgz6Vbzz/opRn00NTADoynDqLrn1nnfGh
QojLh3V39wIxu6Zu6nDbjFjSNw+8PR8fqmRWnQphmdGL+IyUFQsV8P7/4KRk+Vd8
GUopvGQDRi0FWhv52TSxMsBoh9ia3UO7kfCX5t91QtF1kLAgjOU1tYkJnHdapxyN
fcJTSDgSklPXx2HVCQOhbKmHoUe2vNlMworstK0tG2rUmEjW8/+FEhsSZ/rwSl6L
+mEyS7fVdXDXavFenN7hCFNoDRx5iRZSBN9UeVtISg01vmnHUynMIDd9KGige2OD
3v5vTo7EVfF84TmK/4pjZRW7S40p3g/lbrf0wT384uV0wGNZAZJFiMLSD6Rnb4XV
NAQd363NhbD+Gwur/tHkXJbbwzF8fpmJFFAiL09UxpNdv7H7+qMy1GE97kyl0Yls
IinMm592oQivUV/4EUD1aicIuXStlGgJ26OYxXas/f2y1sldQee9jxifszxktMo4
n5KEaOJT5MWJN+WuEXT3ci28D+3aWo2FuI/+jjFqWIihzlTHPEvLm9TkmV15k6Da
dOZ7cd8Fe4vbdzKINpT8ZVinAFARdKYotT9U5LmYspSVzMRkqX2i3KHidsBww1tc
OOwc9C9mGMA+xpc1/xEg9fc8P8Q5VQ5B/jekMj9LMCXVJQ593SUkosnTX8eHPyzA
RG5ojD702uTmJPC5xD7q8bQPiFj5xRUvF1+f1CXsVNUFJeaLWJGc6H+VKMWZC+4j
MKmTKCZYvcowo+EWLVbFbjdvLi7XynTmzUz6kOXYzfPWbBsWRDzJVth0bTfg0vNl
tkROE/VyPQ+Ol8RpAKUK9YEvg6lDjHC7RRXmgN7q/3mYFXJgxEIvn74Hi+eHDEmr
e/TGny80CUTIil9gVyRx9VzNs4vAIBfMEmtr4bVaFFVGyH5nb8hPKIgSmcNfsVP9
SO3KHvCQVR8yK5lJr/AnUIil15Fnpr4a7O5eriW9nsszgR99RWI5HgwqF80k8qCr
imtwgylYMKn5V4v+rVYjJJ7mfHP7c2fKPN/8tpvbkqBbFfKJgUuV2s3KeAq5XnSy
9HCCfq4hIrH6q9kKGYU+Ev4MnmGJ6BbuOBOq5ocMNgdXDIqarGvG08jH9nQx0v1+
GM6ww19BpbgwnnCrW5ENw0BLZnBOu264vKCo0OdnYpmkHq+rms/8bAj8FaCvRo1K
fr97/ZYkX5VS9JPOni2gAPBtNDxS5+CtpYHNG//R77dSNt1ZaPhEXgs9diky+yxr
nxtN+L5NRPSibMfhjSWT4ESgrwOKlhWYo1aegdkI04iwjr2G1sXAPiG22WJhL4uK
zbIZKavJA5+Nhem29C5FoIPoXMcIGIf0v08WKlJPMdRPCo0jSFmJlSjQZ23jPQ5M
DUFetLJHU6UHg5u6TxGM6Z2zmMxz3nQQK3cJ3if72soU+UNDhvqjlmAUvae6yIE9
ok0AdpBZXjqINMTdQiETkCqCFZeYuivy6kPJ8vUGuRBs0DHNvf1o9GUl0ivHgRCV
CSRJ9VVnEs1ne37jz7886Aunb9lri4mIhvexafVllUJweSvj5DOo4jSw/CwqBg8r
FGucUOYp9yvMvfpEJG+Lbh0hw9Q1SD1qZKxRBqVi9mQaVduAhqaGI+LJw7lHFZuS
XMo98TkKvtzQ8czyp5dGc2L7bBgI8RmmDvgyGbjLylvmj8Ldxpd5f+0rd+2NE4UN
U+yNZqZKZx1337LjA3xVelFccX8bVmH/l7JrVUb8p96Zyeng7aCIaXC5/Dpj6sWX
8j6QDe/ipkI2C7L+VfmQLnU/qFBxzun98ITThiH/K2mXqxExr0Zl3S0vYx+T20r6
BOuJG4VlPrbpgOEA+n1FXcEKFVgf/Vexzv1Kj1tBjv1CDBnqPhModEyVwp/45+Z9
C7lCidf890ll7m+6TjsvLD4FfRmws/cVSOAVbXKPbMEuXMr8PymiktQbuxhaKvgq
BB/TaHlNMhJuc8OJKqduHOL2GXtIZSUeA0zfrOH8xh7DuaUeffMUilgbclIsjyUu
Lb6dry/wF7xJgteW0Js/IYd+JAmEWdzY6IVQ7uLw//VevQHmsBNysNmTBoyjzdo1
d0TTLuo/EiEW3AHe1GMTnRGSCpkVAZi2pbN2VjC/peYwPW7E7Xty16VxrH400An3
ceo9Hngbh6ZqTFU08foboqPQS5biOxe/iTNvx4QH5jtwWvzf22e+Lv4GSukR4437
sBFmLeKdkvKTTmMDnL0bQLWE88ZQH7uNNf0apAdNQId7cHD+KIBmHB+4KLvFjg0V
RRTNvZWr5YyJ9yrmKOa64vaUvq3JN0dlNxWfzuhkGqk7y5DKyy8g5+LFWJl+8YrY
vd75Yi5wbrvwCGdDhgjpBiey0gdkyg9uejLrPCFWWjt3/G1u7QfXiV5lCsB2+Khn
JaOckdRSdxijJpu8sbXVgTKt4/H6al9XXj9lPSS+Mm9N71x2bVaJgoZHzfda/zcG
rPXeE72iVC210Qi33xmXd8kydhjq1vMGxD7O8OBArwcoiWQCBI3nOFbd45iAEduy
8IhulIEwt0M5R4lCNLPBGPgmiVjenePul9zomV0tNa+T59HFC6BpSE0/z30AN62o
bSqqvkVtKymzJj2Two7+DTkb6ZKCiLNYfUDwnc3q68IEcyD+txS3A0zCzwFkNI6o
NFt7A6gazozFU4tUY54vMQDsHJt5XTeQmeHidLf1ZavtByzLdBhh+E3oWZ2T1JUP
/YcShhfOXnXyBJRkMjg6/yWEBwvRlHCpcX3/wmHQs2Zl6ydyB80H7BkBFYA88w30
IJ3Pw2Zgcj12WvxAB9EJXAYTSCGlk9+02PeHIFbRSTVMmJM1sl0fU+kcV0EnVB/J
ZE8bQ/zU43QWrfj8de/4FBA7UFzQo9eTaHmMCuRYjVdlEsvlZ4vrMKp75ELntMkh
JrUQw+VbuzTevY4nY8iK8nI0zFYJBorQDsfUKeg725a6WIivHLczOX9MOsJ7khek
v4b0ISrkuvQcMktwakNHOB7zzKd/pTR++VmHGR4niAi5OlHsbMzDMTLPu7edOpnC
i2hSwoaL+Y3VSl9v7sjSfk2viOAJgspGIFwNTXRvgKm0TdVMFmoED8uNUgPhqrkX
+QLJY6PJbcQsoLm0WUBKy80xdLyz4R5pXQfuHtXnYdsUmLeF7GTeq+Tvjkgc6AWD
9ATVN3nZM43jKyxJF4V69qi6RXijxPg30zp4R3HAFSHKNNyobMV8NZ6U2JlumFfQ
4Grs7xH7TXNgdhXezafK28btPMS5qgwCU1sQGK5TI79kxEAS9n3/AbOPVkUCKmiw
G27uiRYriEFqPL1NvxMcyEcrry7fg9eS6QCXiOT3YNZJVcIHV0s6LDjOq4VAK/w0
LaZuhGQJ2PNSdN+yGOYGE7vT43WdQ/2F8fhSWotRKWovWiQY8WVDhLGrxpRjkLV6
yuYW3bENjFQ0ZnSz6Po0e5oSfDWz+1GtM81sYUDEjf8leUslDnnmw3Qw3R/zijDS
NcQKQ42+pM/TopqO6o0wZK50/09XAJSx97nAaF0cBV5uFIyeWVEHS37QbC2Y/oWL
C9xr01yrWc3N2oijGtIZXPwycrau2zzzdmK01J1T0AQ24BsvHa8kscikkL017kcc
NG+UctZFIFcNhza8AnJ877VAKuem9AbIYYZ4L2Itm8vvzUfsSjcARjDwXZynQUmQ
Qah5mpO3oGhxf+crAYhzVQNd9CyLIXP2/ErFYxIlB0Zspsu4E4hrOR/j/zpcp3iN
f9JhybKVOTuQbzdICHx00fi53KpxxptJLeWbzbvHxyZTOD4XrZgKne0BkNHBoiMu
X6bVau5/B4qlBAhQhjrqyD7CRz9zq0Qvf3+2sYjPfV4M0CinKqx6Bn3qaLI5kMP0
m3QJV6lAaxPigQ7/s5l7QPWEU3UnFrG0zyKANDwruskjFu3621W009kFSSPR0E8l
iv4VXQCK6waZdzapQykkJHSimLb9P/w/3O5EjqjLBFtUBLuJ5MhbyKoWWyuO0mXy
heX69FDDQ+wWrPosA+95IoAbyvTI2gqYb9lW9wJabxRwuV+TQ9TVMnhs5OkB8ur6
9UuIcd92Q3zKzq2JDBoZ9ZjmT4IQ2qwtROBhrwyFgyzmjQUqsVu86E3Jzt+zIX2x
CmWNpMv3remtpaMRNPWgdQDucOIhHpXw38q8VVHzawfOw7EC/vnDV09wHHdKxUbW
xSmAMX5T11pUUL3pFRbdu0JvuYrWX0rA6yV1jCUgNBNreOp/A2ux5SvIMgTN0Nr2
UX64Vf3OKLpQs63qGvmUJw7SzoZVOfpozDOV3DJA7CRc2o9WaTdiFKSmKiK+d1dE
dpsrYI2vPtNU2e58GJbx/V5KxPlfBMQ+Nq3H16h1zMVTKGfhCg8CAjI6O5U6+d2n
VSf14a0GbuwL6LZCwrJ225i8JtkDrQ4bDXaEx6/3MxY4mPi8BuxNhgTBgN8zOUQk
l/nAuypWd4j1G/LIecudLZ4InbqBaoOQ8Qvxt2PlKJflrp1Em2gtuuCRiarC1Xms
9jIW9kbkWyVQHQRw4nKQ6GiGvisDEwkPVm+m7Rh6GkOzCyQYmtsGHgPZHt359zU7
Qt4ta6qqExfvBWmnex5e/M8CnxFKchbOC4YyuHkUJWrgY4dkLF/HYk8CvDNGP9cm
S0nd0Dt91mtcS9e7CHy5L3Lxp9ipuDRDbEOkNZWlzgfEPO9zxm8RRpiXYJbrRPPl
bPZUm7AZRMHgawkoWQel1spvLKDETA8TXOAW9KAmgfTNPNF8VqA79Z09rLuOIb1H
XA640zyYh3WjWUDEibqiVDkqhwehdlR/yuK4xNOSb9MY/jDrEhFGl7Urckn40urn
CxsnLez45kwDVIm0zAtuoWrmCTKRmRJ7JN+EXEJcqU06AcJqE38DD/GAIn0d//Ah
pbPKjA9AyplTtqoVNUzyzd6mBb1t2ZNe4sT4RutlFEe4JPSqIVNuYzJtN9oDhcPk
6OhNrEdJAuo31P7rBy0fV/8qVfpmdmHaDR1SPPNrJSP7uBX26a18us6odFqWsfB1
7ywwctlsSk5eigSHHu3xNS6aYKDQqi7XtEIjrZJ6q2yuuoMMoFU+zrJhfWnjsFw/
5dKudFSee4QiAANzVseBvJI2pYDLGL8x7gs2oyyeUkbfYwEN9p77SKkkvhsG/4+W
uDLyzjInesdsY12/ASu8eT+zMwKJrCuuMxKH4m3w3s5gWvD0oF3gcLovG81OA4tk
piuYiEabsfCjsWAJx64IrFEWobB9Ws5D1oxAG+1paaMMbyBULWoDd6UeYzWTyiVl
E1Lf+77XWIzWJQtNRkf9zWu6lbGABvb62tcKaVJIPy0OiVBzzU0aFvwQqbSpg5yI
1h5wkPOv6mhQCKtVLEg2Naj3kmxDWDaDEA4NAWLgo7fSBeRoh70Igkc6URk5cOKL
PzvHZET3ypRhEv+R4TZJAhaTATah/G0pjysZxnPhaqKG5NIADaVp54p8PoRVk+dZ
N4LKd8oizAStFgl1UBXkZgPmQzfbZYuQ3rjN6IY+los+BKWSHNHvSR7kW3r9yzp8
bVvq9Viwf4EFI+WQwRn5CfJhS/MOhZvQ1j6cdBC07u2XtLQmyaF7BeDapHC3t5TY
bjKTnQXfUSt5c4ZweAKvY+fpNcMv/Zh2QynBG5yr2A+N64ZAt+8j+mDlcNSFJlIY
PuUsVlKTWOk62bMCjBfA5X1eqeT7XgvxQltDoaxYnVllFoapKsIY0ZSGpwBg5mSH
eDaS4a+H92jfrBKP8wODse9w9vPxfUxElsC33ZB4VWUda6m7YY0uPv1uzC0IUitq
G0Si2lxnM00GX3rQJ9VwAVwX9QHpBsWvXBgX02JzyAWsbSsoPkNoBFiKoCTdW3Cw
7wDXeIZreNdkASOPpXuDmSCDCJ2XVrmQp7Zl3qoSfUBI6cK/PboAL5NYs7kutoOq
IbPWyOCvrPj1sA+Nw1ds807jtvOIfqRvrBTzFrhErS3y6bNdzXdMBT02J40Tgz94
82oj75vDxJ9TmBbTP8fxo4TP4E/mgoiHX281GhYUsyxTVzQjaaCLYv4Cz4CF3VeJ
7nE1qrkDemc11nEK0ZUpXouwRfLSGbh8tM3d/R8FoVf2NsetKZxJbUSLQmxXwVy2
WJ31cOF7p7+BC4IvmCglhlXYGCxnAWclOrW3FtpQK1XcEeAbV5Sklm/Y9cOWlVpH
LmmMmbmjYI6eeRHHydpmbqOrcQldfIKd2gw128edVj0zuIevUTZKgLN8DgwOlCGD
6VVMBMSCFFBEECACf4KzilLIYJaAM6yqsshqj2GfmndxXZ8YtTkcvusQS08wTPdH
TJ8A9dmiKccfN8mezrHz35CYRYRk6CDUAzFSGgWj+5rYZcRv3r+SjvLas9yeYWCb
auoEktz7MXIt4ndv8cievA/8R62Vw5y0sEvqfnJMTnDkxdcYMpaekMmueH77MsM2
FzltnnsMlJ3uMzhPPX4bk8yOkyhl82qb0kc8hKOypPYBUXSnh4SKhWkC0somXyhQ
2Tvs4i3DCpVeBTwB7M3cDOTyaNwlh7NH+PF2dzr9C6GOTWyirpwunMwv66y16Ndz
flDFeUa270mkmvXiJ6UvsbpYCJU7wlFUgNdiNm145iGJrst7zEiD211Nih+Hb8fa
+QZoNkxw+FIKJxl3ExhDiVkW0h+vSvMzBWOv59E/bMKR8mrWtyfMkgO09mCp0YeB
MHcyE4YPb51NDamN8sai/QtulBNpfvAMvHlAWkbmtVkBfvtvbc4iqKEEpq0EmJpr
P4td+CSC0RD7KSnquFunQ0NXBbYO3M4KiW3MzU6qssF26sLx1Lcs2RWe6HdIlss1
hE8PK4Kyp0wgJUMS4TdOVLnTV2lFvn7Cvy1oxnUC6oW74OItRb00MOdQQ2N7AbKF
qpAolGX+xatEQlhsSAjD2qUjC2L7rKGRaoMVgJy3+uwhr8GbjTmPHgKmdkR+4CDQ
NJw4B8ZUakpnpEtOXZaNRFXvbKwU1VJ4RV3TOD3UmQXlv3KCmfN9OV8GqBIEA9Nr
7da5l/3aPDcPNJsLlreNfcO/IznZVnux36UQuNC/Z4I9v113PSie83oBpHjqTbi3
4AdwFC6+UiNkOWlvetuzA/vevDvkv5E5qAyFpG8O2KaqcLC0tA4oHGMWZzOX9rTX
Yvo53dmEMMcNyq4Si714PWQkAUJJl3QSqJIVECiYF4qqTO6zLCPu8YHGGP8LeuwR
/2QAsVTEDO7yYxUu2S7kj71qy9bl55VPCN1UQ+Et8TIY//VopxOpvevBfOSNA92U
IiTB7EzsNkdgVahR6+fTHVWEHumVAihFxWNIk4qfbIKcEjHjWHeIdvhtfZgsb5m6
CkuodYtsoNTfZQCJTP1887fhXAUK10p2nOb6yTPGgZkelsjJUupn/gDyqX3GsfkV
2zWA9s9Hxxv59Rs1No+0hT52gFlDtVdZyKgXnKkWCi+5HVu/CycPt+4EQ9pjCYsS
0vcKJhqG45s/XpDhdSUZb0ENjfp/qUMIWKTHH3VynmTcVoiL0eRSvUjwIybuFSU0
I+v7d3qq7273wG/qMI+JgyUmU7dU6HOKDY87pzWKL8chHluU8lw6N0tZDRc0FCjm
FjzFf4We6Z9qC3Q2rkKiN4bbnyy8uY2150Y2oQeOu3XmTSOIboiJPCVPCVDMZtvZ
KedxB7NWS2UwnP+4BvdhamwoI1gf4E6r5mH+1tzqxomiYOPTwuxDujWgH/cMYjQC
3qeBYszfbQrzyytjAHT58uQH6OSqgTBhWGvV0cScO6AlRr95ycXpm+hntwqiw1wf
J4M5dz1qQ4ufFHrhOchrjKrcUnmYFFQOVhLVjr1S0CEfpjxgAXgMInCA6VkV6WBl
/2SWIeWugilmZ64XXb3al+WM20N1oPqP1IdXMgqsq3md2GVmwQ6Rx3vUZtrcGlMW
NURzjxSGsrVF07xg4TYXL1kiPDwPC4/nVJ8ReFkhT2tX9sC1bCf9WAYrC76ndRWu
Z1ifagzYHHyakEyGFq49mqktNqSPw2xfcdh97xQqd5JY21s5UATCQZAZGsw13BME
MiEE5BEVoc18KiddkaNuHQ4nR35DGZETPixXZVoTeBUrh5Lcx2OsK/BB151XsFkm
UIvpqct5WZ57KLIWaKCLLzgs9vKlGJosmKQVT4Nu1WDKo177Cto3WDjWUrVWfffY
++aFliGPIWubNOBl/hYfN00tj3CMyuR/RISh7K5XBsZl/jxYa9COhlIZ87VMRheZ
O89NlLVgVL89eI1YDipzcpJbg0m407WMTfXCBviVMH4uOpoPgjZHqVClvExZ6Wzp
Y998penLTRIgfb3iAoROvgX6o+CETKmO56lVUbOe0OJib3JlMgreO1/1nVD1HXH9
HgNe/XMmehCAnOuOWfM6RoC8iL9eIh9shQ0aa60QhuV5sciKkK0ZM8R+jrRINEed
c8mD06RZGgLQg/mO3zwWqgCGi8vgtqEWtRD5GGr1BPCSGLZUesKQq5Pnl/ZkRVPt
ge7g8psJggohcLrvprPN4QVbeP3KAxytpS4vLlzLq0W7C99b3Xp/UFUw5GRHLWpT
rKokRcE5dez6i5bgyNExNF/300HM4umMMFmqIsOUrJH579sXROcVlzbbP2IbkS45
esTjl+Zzd2kU8VkwRNJD/J7FMUR8HoCl8s4a3CBQ5wj4sQXPBbHjJD5OB9j8xJbA
EOY7u9B9ig7O4wZ+796rqFxvGWDUUzLt7LSRNp34E1A9FJyHxuAKTSA83H+gfD/d
gnkb9wcIFzDMZ19KN7qSgqn8BekBeyFNPssOcB9UhmKp5AI4DaxPHYmMtIIWW6mR
s1QSCmKoFdvS0kdRPKAmTaQIEyIZnM7mAmZrQ1xioEQqUWhD14pfwRYilQMF2E8I
KZvC87DL9s8yd+LUnHAS3DzYP1v5ntWy+cxHLDI8Ajgn+tZ9ANw7nUFwZQ/xvRO+
XM6pASrft0KtaXgHeEBHK+l1yavI/o8F/RZ/fXTrmw9/eWrtsOwa91FA4w2YSy9q
kUkJdeXj25lZR71GKs1NrsGKrsFgdVAOrV/4w/p/UkGkeOa88hWEYV/7kIQSXWQO
mHxt3cAPuwuzifgxe12MrTAjoCcIpJUbLJOBnw+BpMaEroBsV0ybuCKxTCUnzOxy
rQ6z52w8KfBwpemQS3xpYbVfvIqnHpiNgP7JJ80zq++VqaZZxgMhwpuADUril3aI
ddhyGkgYpJ1g3nGKnF+hYRzzNMx4xzJQ87yWUhcSfpPjITXdMOB+FmDPNAP6y/QC
W4sN9xqIWjvWbV5M+mqAByGqfirI3hUsiSIe0h5hRQYn5Xxj4vf1FSLXnEVCnMjV
GBt/RVNS7EjfrkKZzsSCkG+aYjtI0aE73zPvEmufW4dtRe4GztyDiWmGcN5Fq6so
WY13GaMSa0dU5tX350mQLvJS3nNEjZlroDLiOxxDgy14KykvduUTTxnSKauCwV0L
ZxjtsiwPhXjT8fMqyDT9m/bMBBYGvJuXKWespTHgNSHdrpHN1Ldu2a3ACger8goq
Sy65qpsq/ann/RX71S+x7EabF8YIz++3Nnm3AjWB9sUiEZOEaiUCkUt0HdEgWRyR
d1fOcVNM77Qbhj16+EF257LN9C5A83mprc/E1Zc3m2OIJ7XRKk/9RCMkO0NFUjCS
zYv5+x0PQJmu86t+TGyuqSycCtsf8HTx77oYPUS+GUEaZgP9AFeDmN+js0Zx1x2b
TOsc0LD6guv2DVr1b7eFpbajmoolHw9H0Oz8azihuBk6vnQaYUGiEvUiCkjHNbu9
odyedJeybDkkHcBypycah9WH1xVj6g62CtcVwJF5aZo6Ew8QfdaeOWBJFhdsh0co
FovhFTKq45wqaTETEUZLkxXxy61Nj18HkDFqHncwtAMsLmrjluiCf/8aoeKwaD9O
H8PddJkEy39ymviaKJEXoyXIGf6paiEyHfaC62yt+ajsiyFP/A0o9LXQkRoH0ieT
sDZLh55dAjwMpeVL65AQ+YA7Q/+ymLfbejSrp0GpK/XXtqgPeti7sWiafwtZkgdZ
3fivh04Lu+14+r2v4yby12AXvuyrS0GnBElhuCmKyEDbWYGhk3iDHj9NzOunfZi/
YrVXUb5nFv7BvxhEhqPdJIgZo6oHnGMgk245EAZLCsfvBrhx5DkxO3/jjhVap4Bm
ID7RMUq/teul9Dgf7xYgbWjL0LyjnfnATAWK/kuRG7rt1HmeZz/wB/pHYIgEabcS
8/KLldLlZGTgHrTEuve3DTrbn90KqRIE+soC+gnfAb8=
`pragma protect end_protected
