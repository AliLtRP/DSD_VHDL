// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q0ICFBxn0Ev4BHB2IPHbQpynUWHFzNWZ6bp/T47Mtd6ie7sRmUCvhfoe91oPV2CW
LKC69X5/H0o6K7gYkRfEW+Fi6QPfXg6xow0UZi/wY2/sLL/ugUEDEuXcndVjTvVs
3iSWp6/st5KWHqyR1yLUKjZ0D2/WKj9HL7DJ5p71Pac=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18544)
s++oRAzhCg+sPmfYRb4GT18uPr5AYy4Bb0vSy37vEZZkSPfBI14qti4B3qyLeCVC
PzY3sqfKgq1tLAMf2IpliOauYxqaBInGGrk+97mZwP+rA1bsZD1SqMuFEsCBkpdL
5KiUPxKZJQR0As5QsgO2aktTXo7SCyzqcFtWIuEUukyPvjVIylcEZR1XkIjr/+fk
l58VLVfQYvBdsSZdjrrkzQjJVu1s27zU9yn+0J28H6bhlq/2FSVovlvMgqQ5S/EP
LQzjsrnzoOQNtPNjzbclS5vpZ/grLEb7p5TAXBVlc0LagARXvJSSntG6cNBb99f0
Qx4eYJ0AghrTvG69iEK0eBcRF3kxyj30cnc3NBB7jz2ib3ar7zXTYsjQJ91y9qAz
FwtyErU92ALCjx+8JEXcQmeVIO8pYhyNwxzVmrb2dsoPGg7qovbO+aBdIK23shs9
Mz6PbPxMUpkJhcha01Cwjs74+c3mhIwsqkjTe391U1SbTfxr+X94XOBnLp5xu1Ng
H0ah3WuKw21GjH4xBi8MtEriz5U+LY1pu+5RYXFGcVuC5lsafiPjlWSsUlDLY+Rv
qv1v6ERFLGzq1EtDtq1LVKzrfJ2vZbpDDdPR9DRIblEWKj0GrpXmwqlcKth1PHzT
shVfd3/lkWVwrBiBaYikGWLLEmrz5aY4mnpmHrmT1ntpIVnuZXMEkIgdn9K3VWkF
1g+8v6qywqcFhPRFaGq/dzD2qsOsxI79EEApqFg8/ACAoQN+9gee0fBxm2MVxp4k
z248y1xumg4RHzmrq78AaWnsFyUoyC5pTEhXvnkBTt1eJbqMzo9fG4xE0HfofUDM
ovjjCLKle9oeGB8BdW+qeO3rDY5Ro8cJ8NXRSZpK0TOKsS0Lqfhp1n7PJq6Xt1hb
VkHqDP7feY4J+4AGfaF462Ozq64DERF/fFfGIS364ngxdT69CX8/LEtrGcRqxF40
yQxdSjwAdxwwurLhKb0FzGdFnKOdmRDHnbbPCvkgIDazAUyzExPCoxfFJJqu05bF
zt+sFgxXVQqL8ZD0mZ5zW+Hx8gGVkNsTZqFvJMM9OwE0Js04V33Jes9vfnvzxP6P
Mk2FnxYVYDvYmGLb98UR13RQ9HH+jKp3CJ4sgdO+1Ak4Wv+qF/YyEpMTSa6w7LiP
kfD4+H/TsgSjGrKwagYLSvVhHl2ovA3OIthf6wIw5v5GARVqUYFmGpG8V2r2RPS8
x13OOiTsKmMiX1hK3Q+W2kmVc5FgIeYBLnNcJHKIFdy0AJC1BpXMZ9/9U3LbuZjH
bgGrZaNO/+YTHnOY8AZygblx+vTdedSfHRMOe4DYLNc+jLmOj3/3hYTo8JDIdJbV
TLowSYIvypcVZjiyQnirPbz83qjTdCPvgFbPk1jgqpw1AZx7vvrB7+DN4ph0MBLG
89wzmXf65wKXckdwRaAc44Xfo5JWkRqUNTsvfLLyLPheBo224cHcbA4D/VvRVjEh
bSv/4cVFQuApXcow2gLJBiMpzatdu43j07yGmQV6FYl4SXRcaBUbGQQXyKfwMGXk
BYKo8+/27c6PyjDlf/GolAgE8ihskBZf+jYs3bQLemkVB3e13uCt2n5wZSUnsIsh
ir0TM9EP/LOAWHFDO2LMRf9KtZYJR9Uo/yBJAM7fGL7nxocfv9FGtLVKYhPFK/P9
VKtHGwM6J7QAbcfOYGecefijNc/C/RflqJDcMLV7lj8BGYNT4zqpQKY3SPG82mYq
CSB8/p57mHMqomkVWBqQvF5bi9JbOwDf7HDNd77p3MscyotnlZYhORTxLeKAKRkB
yearJVT32/935nRKeY8XHuBlVZRwA3B1nGJPeXXlInrny/+448SqaDpZmHOefG5d
xLvj0dZdH1z45i4aX/lE7/a0YdLejT6sbbrD8gJcOkiVeN6kT7d9Ka2Lf3eN869t
kVOHZ6uGc7tbUrrE2ZK6rSFdEtNjkwxbsgu4FyBJNQFpxejei+6LULiu6PHW2pnr
YzTrjalhHCB8jT2RRkM33PYZQ9bt0rdMMhRxRgz0IWgbKTSjo+zvC0WgZen0RY40
Adg7PP8aQ2u/yYYpn7fxkV79LDtphRB0Rs38H+Ol7UaubbixLh6zoNl1si0eIjGF
OeLOC8uBx0ihGFROY3vkjMQ+c0bR7xc4D2Sg01IxcZRUVITbqEki9j3iAH17Ilhs
5h+KkWoaNzRY2JcDFBPqup7ZKvgd88E0np31xgcaImJuclkwmVrzxtrb56g0x170
o6Kx+aHYz5aH90CBb7RDyX1i4RBscbGVc8LB2IrU1X4re8UQIyRcOu4Q2Sn7Njbr
qk6JjRkOtu5ZQqLYaKT9Gda8eFNQjuKIWzlvhvcw+aSgZ0XY2/1kt32F+0x4LAaz
37oydhFSJ3RXvUEaZKvItI6VI2yC2WP5to/Z7lvglgkFJvbmXx1231KyJEJD02VO
DtM1QqKNUoAndWzhYN3YFVdoOkK7YJzUAJojN3RPgfgJ2BN1EZc/VePMoo/v7hbm
i9N5gQLTlXKm7VM4yC1gidhxdAmImXkc8bXAIAKANFY4w5Ee10Tahbo08q2eP/P3
EL4gI255MSd51M7Unb+9wtSBIXwkuhqGsSeQ5n2KkkeJZk1TEancdLO6B8c4kZ+9
JDy9vJcsRBFfeQHTAs/SMe1CPDYWwcyOQqyj1UK7F+zNORPyfAgH/q8RUAbWyvRp
DqJPLP1+bI71S5ryKC8tV9JbF1vjkOhzIS6zO5cvdFi8ci8Dbk1RFoj5W3MtTD0u
5J5yFOlT+2tPm3HPIw7a9Ga+hDXAWt/ChIIBVkf72vurC9TGVBYpS0mFjujoE1sY
zbUhfOVIiyk+dVGkezdQDvhLq8oIkWcOtS/nL4jBZtuBKvXmvwOn+N2FWqrwPR0F
qi1tsswjw8SjeM+xEtzOwOEuVzH2mQdUqvq+ZT6QSvReT57CbiqIlzoBo/RNlxbu
p9eaiqGIdmX9KQPRr5kTyferV6PnudTflqUZWVvbTOnFNFl1/73teJb1Y0HeYSPY
AL68XOO44B4PS9cnOHie1h2mU40LdXs6TjsqEjiunOn6WZJOfROiHmp+psvwsPJm
BBKZzJpDj5Kg0DHsPiuSP9xDA2KVcF+EIOxQn6DpvmEYqzDlJ4D7jnOnlhmqA5rC
PeLXxWgOx8RZewcrzNYakqcQ5DkLLe0+Eqq3vAMifj0fQJcxbI2KIjgGipJ0Kb/5
QUP5Ft8psXEoGj/Qfr9s6gvJgJd9wgt28SBVsGmWVHL9hJlOrxHLP6B1E1yvyzUR
WAuH3nsbCQoZ/tv0JqR34GszDGK4nwaa2F2vVWq9k3fTB6S9b6sjUipCaxNeBmUJ
jUaCMkhu0HgWPPLOUyt3VddzHW+G1WdPouaneIC+FMhiSnAQfAp/DZ+YPWDiBa36
BayVQF44ab6KKUZHNk4USM+VavAvVtPaSFYp1fqs8PHdwjdV8+tudpw9O7ZQVOfG
ctwX8qWkLBrAsuzVZIHLyX29xJt+ApMY+q5ASJ5bK5M0yDA4/u/U999XhmMQnk65
C+FqC2WX0KUj067WernqYBkj/e0Smi/Zj6OB1Ema3Esz6w4jKVcxhpGXwjnADOQJ
pb/ObYRP/vFyXC27NY9ZwrMHff4VCT93Y/Xnerelkn94Gh072kGzMKVT3huoaeUx
9vmFuKxHbZghLJfyciTax8/Xz8QnVLxZDKxRQjCnBX6TlR/D4RZWisJEbO9cnRkc
1BudBnfxrYiAUylwwgnm/4sCUxjBMU8EW0Rob77fRIjIeJotCi/ZRb58OsZVrwfN
RKuSm6/Mc//wWVoK0v19gsiZIycZkjhWfUxTbHSuSpP6lWZZVn8doBYOjfkDHnAf
/D9ejRjVeBdscHpjSWKxgKPP2Fr7XYyWZzp/bBpDORPAxHsttGGHjCVwptS/PeA3
ly5aTTVIBkcSr8hPioQtJXOu5Po+R2CT4pX+acgRamVab6g+G4hai9ArjT3FTFBi
1wKisxUW1F9+58ZqonsRvYzZtXOPfeeGUnvG4U1RDMw3dKVMsPRdo4Zf/vccJHa1
V7kNS6XVXs7zS1BFeFj8x7MxfsXV/x00G0lOOedtiJIOrVjim4gbkwB4osY2fa0w
oCUpfU/Bn+cG0dKESqyT3V+ZF97z41yqUahqugDhOqnmx4fllWPk0okhJDHUXT8g
AlIiQoGV2z+dfQysD6ywvlRUJWM5vbhoxWdLJ/fX7whK7hgTySFbWDhetUNWBHat
muVdCI35yk93fTtoGcgRb9fJ9lbkKtufK/+eJDrxYu78HSzatD97CIrtQIqVhH/r
cTLMgHgJzTmuuvn5VSA4Cqv1ILOP31qk6MvS4TBGcgMV+5Zht+ZIbHLL+7kQTM0L
X4vAC9Y8CjVbx6UEiyPT9Olhks0y7CoSz/p04mx3AsWZe4apfCqyioGCDT327LJ+
tVgPmzIG4cN8ENd0xWIMoOn1yCtfsY6RrNVVB75YgZ0SNWvOt+ES1YPbBItcOaPt
utkLM9kGnSnH5AF1Q6Xs88niyRhDew2T8/zRgrS5xhLeqRQnluybObC8Q0uRMdcM
g7uxmesRTifyg8MGwla64cWvM4mbwZFWd82x2bf2/kAWwSPCE62EEAPS39J1X21Y
1kyOeTufg+805XUxC+1DTYvHlcAwt9z0Iw47G2xfrsA1ZQmuQSN/V4QlfVFZ49TE
qzxfp41HnH+p0MrTk0bKWDWe9GIsjLQ6XfctNmkNIy8JH/9CT3Vkh8ZPYpLy4JTI
pNrYxTRH6FwhmF2m2x1uDJRcNBi46O77Kbibd5PaTIxTWLbJmXKwaxVXQkGNl088
iYiQmsMn5q/iWZaHvEi2dK+wl8LGxgbbmQG2MqQPAxhA0Snnxq4DqRGfO/XnIZyQ
if/Ay9lLksLn6KZa9qdyMPb97K0eOn2FvrXv+Jqs6BxpJb8MORhPrPDheo6z/UJF
sKPaY7uXKNdtLy7m8HzpBRNWN+sqX1lHl++vooi91/ewRvJo8keaQGj4w+eXI+w6
RQ5ClYlro/uNOGlukV7aAAS3J+WONN9JSfp6hn/6fnoDT2Y44lMRA/Sicb+W0WES
bJ+vyP4R9PRZqySioOGul9qIIVdm5n1Pxn15885lQEGTmggJFAiElQUacjRX6Xn2
H0nnWirL1GVl3HkDn/0hS+xTsyoQeswEUlL+oJ82PyJhk5KbKcyhZEcUn7FJKJmQ
msA2jFFL2CIGbQqfdToxyXGNIZ+qDlzrVuGjRhypToMw9bAUU8IFsymeY8RxPq9Q
eb9n8A4eC7R7uw1xXtWzogq/3u3IMeVgrUQK+iNlWPgSCa8JwKP0xZ2NbTWzao4F
U1Rsl5guN3WOaYAsRHXn2x5YXrITVUU6DQ0LxNSfvXiykTRF/oMyS9goqCGGKdHd
lFQi6xw+F58Du1B5ExX86W0IZ1YVB24rtbLqd/ngjnTSPDCTrMfSbtxJYoT/bd0l
etV6ryPAWObj2r5/dQcql02i3jaAqykLPIqIfPnYRhnEL70m4ts2NROFGjOZZZMU
AFsQHq0FB1Myf0+tRZIzQ/TAfsCWRvfX9I17stWb4j4WMWtiW+lSop0shNRSjLPm
2/WkrfH/SVBDJ4v8bDSp76VnvS7xEP1W0YPtyXDrn5aQ0FgjXC8MehxjBc15+xuu
9j01F6NLAQO+eea70SrkQ4vh6Eqgzs5OfcZVsvLT+W2Ds2aYnSFzEx74h5zEO4h9
3RL9piExCS66LVM92wEjZqPgWzbCp9ykIw6u5dvXOQJgkL/VDhojTaxQy2z/emPq
EAosXpK9l/eV7+4RQqvTfu4LdYG8bx3AEXQrVim7bHWOxdhL2rqy7DtTJ14FeoSj
VewA9c6kv4YW7lYqF4q8Mue3sUIjHuHwn7YrJzaY1fP8U2koPKYntbn/WcpDxytr
EazTQZdJ4x/Wd9kEM/Uo/OkqDcPXY98YrSegyEUtN/VDd+7HJZQJsE05+jFnXsjE
rspRNCexLQaH8edv0uURD9JpEt7MKHBdz7oPiz1RKKnONfa+cj+uefHrDtg/9oDu
k+IL946GRmcPMMeE6uq2fYqFSZnGUKaPIOZp7Ux7/xQr3/5Eq4k0wWaBzKHUrnsC
nGRzJuQGH5egImqvtCOhme/dqglQFxuEcH19eFDzOiBb4NdtFMlvvk3yAwd67SRR
zubWHTCNR0KCkh9FoWERtNiqf4hVC6FT6h0kMmliDNyVaAlv4yM0fMG5lcnFqvvb
0pMZSGXrUQREQa4GTJBVB/+YX6U0kOu5M701JKcwvDXIX6NPXTPu/HQuPmwh14OE
xt8oxeTUE6KSSbKxyzCG/QQKvoULI4S+uU+T5WErlpcxzLsBGps0jFtgliNxrHBq
7tu+aW2aB1C5I+TQ3vjG68Y7DBNzv6g1CabZSZQPHVWfbxqDyL60ylckzH0ul6Y7
9ihI/2sqXH4PdYjREiXybwcemvGxwqSiYSC9m3bQCzGUdzw75ruir/71jVqcFwom
W5egqE2/+Om2UEv9lWwfaocUhplgWoIKMkK6+i0qpIjH8y7sIvAqh04iyijvhJRf
Q1t32WNPS4peNyp2GUQtPHrYVeEWSDHc0aMGP0RIkV1fe7EY1AInyyo4vBtD6cKH
gT9NSvAzdygbhxhVtrup5GdYEgMu0/mkAxjoY1FOK/DGN2p7ihw//xEXVmQYQkKu
fvGFNRFFJkbsMIE4ia8RfhcAD6VX3u6LvGndUxNTU7hEbSOYN0za1Da1Ng33w362
s2TXVq9hvUThjmXoZ2WS77arRCpih0Qw6RqYu3OOeH9LlGQ/u59lW7geiH1yIx61
B9IRU8Fdhousxvz0lRJb682XNCILp/16dzxdimriMzJew1W5eA2fhTT0ta1G4Wa8
DEqgQuhDhspbVgLWUf60kOLTup42+hpF/86KB71jSzH0uHhBHl/1Q9kctiz6i6kW
oMJQjWr6g3rF3HI7bPIvluyliti4xZhGkbSLp1jcLoynR1Fg1OBueHHvjlXwEs11
UoKeJ7WgpYBYGRUGxtMHJ9+f13lgQ5IQdAhfG/TOwDO9HUg5qPQLlafWMWuv+EXD
iQmwiCd+DnLPk5GBQCst84VC6NLgBq/ko+lQhrj+ua6PlBP+b0u5kxHgiYrGJzkw
BsmKLsaLxp1bzpqNJERibsIn6W2QlKXOnGgsyqRiLWtLZm6b2fXryG6Mbk83VpNs
4ElDFsqmrvqZSjb48q95cBxh1hxTafPjgvdBRytWcIM6mlPfvLYTCn1+NbNI/zs0
jvIu1qyxf7urbgnDaOnjzonl+j95w1XEAojm8Za1qgXPAFaxGJ4UVZjdm9O77qUe
1QVPAtHb60f+J50ZLkVehHFiwT94mupjSZTCyR2236Gx+jfbbJ46a6qRyS2QppKl
AaqFzNZRKTiGsPHsKl+r0BCPXSc9EWS5ARYObJQQa77CA5kPgK4bvu+AjxsCVGaC
ZjSlR7nnbofqLZhzVRmU/KUz72PrJt9KIStOfJ1MsFOXSsR0rHKqDMqipwzWLiji
yGi0wRTyzUug2mOEgJjz2eyI3RNyLnliYckLOnF8qzWN6mfskyHqHfJ/1a6wRYgo
PGafQE6MocJ4dA5I0O7kF2ZiAJMFxLR488RDtN7a/Tm4kR5sK8lkI97lCaUHPCf7
UFtXf4NPmRmpe+a5rluUXwkXojD7D8GBywelXsKBiVluqCTQb6Gv7RKAddwpVd8o
lWaBfYURPF+4APeoCmbigw0zZ6eKQAvKXG7NBUzh2o/TOPmZbATVdsfDSimfZlvR
GIJQwNkVf4wV7Hm4Xf4NcbQFVPUS0k/B8PpK4syQuhGo1SqtlM/+oZBlcM6y1/yy
3gPzHwqy0G7VGKf6IsDE7VkAPjRn2KPZZAxpAZSlyCKbNF2bg4SuQNG0RquYfccl
jmvuWpDwED05H7ERa0JHi6Lt9jm2Enp7TJivAUtuIDac3CIjo36j59pAoP5E+nYX
E1tvewzp5uoXt3q1HNgsC9EMgjeySXkznRotcj6xHgF4Mg8sGPQT8D/2vWM/A4mF
f5OXZCi1jRJWY83LKkVGvbPp46X4gPQLsmd26uPPFLI8JCI4pS3+N7FoQx0Oe3g3
RJBPmcHwKuSELhI+QAG9sP2tHRS1ujnhEtc0+3D5FYJ1L0sjQWP2d9rm8KPoCKBu
6SUHZ1f2LOwjvTDGSYfk+jvVEW/xdorqxOyzRWRuhAA/YcYftopX0Ew12QzzXawy
xdUZ+VnD6yUsld/JznqNEsMwyGH4FIScRTCqc2zK4pkWyMdB3BYrgNu8LYjOuFmq
HIEwkDprxxOfZFk8SE6ogwqcRWhfCUgnL3IgmZGAx8xP74aWdFuqChG6vOj41Mdo
O9wdo/O/VQ2R1Cke2KnhR/ijv7Km7XMmarX2Js3DzQNBMQLeg4UWMgjyG6Nc/5cV
ZfTRJ6SW1XA9kRpS2G5vM258oIEXVB8hN2N+u0Q2VYBSsNraEVbv71u0kUFnhkGs
uknFo0W0b0kzxLXiWk1Bd48Mgn/DwBWIBO/ULh1yp4Y2nvBsrld6FJcaFKwiTMlq
LZ+fsh75FnCZmikuVfQabANHZ07Hmg17S/DzyL2EZ6aUsYK4r91I0+xHax9/qxbP
TQ4GtMh9palTAwYEUHZiT5ZOAGNoMP8iSLW+Es3Hukb4e6ITuFo6otS+9uWajp9m
KPTG8gt6hN1gTd6SqWtd1ttByMXe0E6WeSwVc3EVBaQsvHBR/EJ/s34nvz1Gppbv
TiYoH39YkoaDdcDWgXyTuJvr/qtD4VeyQ2MlnXsPhdy3GTr/BRI+brc6k5LIhVKJ
P61sPOobFiSVwUWCBL3s2tdyPITJc+so7WWAUYJ3r0wNa9Nyu9RSiSbQmd7DYnnB
ev/kGNZPwta9ytq1efRpjKlOCwqHCkCK0gVY6dbGLS4PQNqMi4IisUiwmUVZr5LC
yccrLZpBzuOXnZeChEDb4Ld47MF1XSQUVWgnBqvgDKvl1UYrtEtqPaC+Xqcc3OOZ
QoEShxz29m7jfqH3Aw8CJ0JZiGACOxyj7JTMxq41eWYEss/vuabKAuLaEk5SR1Ua
7uYl0MYsAcd+aARMopIqGuK4+t5yaLN4m0XD6+2b8JF577D466WqUYcTFmi8XzkK
BlcXWmrYfPcMNYTcVA6HuEfAgTtoDJychgsf5skaCdfv9ielywEsMKNbPmLfSt90
Jk89MfsMX9/aufpatl0UkhVOfGkRpbbt4zWbXMP3UARCPECC4iXWwrA470RrJSet
QJJYVbH2sEZVje5fKo0nar2bPDumHvBN21H2wycAATKdPB32BeJaGIfWb7gvbleX
nIo4SV9kmIdo0FJ+xfQJCSQ1KvZ0DmEsqVaj86GERjsWgOyH9N7ySmPXAik1XZZI
UWCAXBMQwwO5uv6cEcsuXc+oPP8x5KwMqTZbNnCpSy4RhSHBoAq/4IMPYZXCws1Q
IzAK/sSz8CYdsU1bIOCZnewTTyJ3xSipFRw/PkcnH17PJozTQdaJ6OwzytIItHS4
v70OV+Ox4AXTHmC2pqWFf/4kdz0kLH8wbgGUlqISG7vwD11Q1uEGJj0mgJ2qFUDU
JRUGEzf7yYt3rjXqzymLRLMJzIuCqQkMhV25Ecqsds5YTd/rjK0IoAo/G/E2L+Yk
utHi6k5Tjf5O8t/cANfkuzG0V31q5Y+O8Nfbtp+YOcIyTgcmU4SeLhACX9JoIhfZ
TtaFcPjJW24eBI3oxbb9LttuDkcx6tuG0sbHrKJWmwWHSxitvxCCkI/vsld/voAz
H54YXD9v3zDkLyy6Fb/ck4DsTKpBY2dNLiLgs8kO6Bd9frMhgk8sHQUw6HVmUcCG
jWHmPXjLgXS+jTTHU2Vu0dRHjNDC/ERWg1Vas5uhDG1BwIIbHLK6dIJ4qaCBCbbG
FfK1p56lSYdpKxkDDPtCvaOmgxF/on5NQcfqKOAfts6ZvyaANLbymGi2nIG6Hmgb
KB7dNYsQbubpTBbXax4Kim7jANKnoaAEmYVxHGb4VS3rLFQovqzHhbyU6xdA82tZ
CjRwJY4MaDQvej9fyQkY+C5MvP1bUDiY+ByR9ZljIsT3C0udo7zqBcqkBh9k+t3Z
sNL3CefXpDER7qi/ju9TwcwB1JRt1A31PyjfnclpqiqZ4co+hZ5JDCyeAs87DqlA
j29DBMSbMv+UP2kEepVh6tH2yZBymMdDYGZDYlBnA+VZQeDyjRp0Z0Zrz1xR1pJ5
5XiqOd6KU+XqbG2cUZWTYqqPIMwWgTZ3ns9eWdBQMPujwrlh63GZfO10MNNlt6Ex
SHrDXaTghEhM4LkFbh3EA5YMDBFh1vifVbEOTfjqVfMIMGayjuTri1Er2qnD96Lt
wqNrXoS2zfjNZ65XWHiCb67Ev0hHY5HwD5Ha8my9ti5uA0rtZeWlJ0e01NnCsQQ/
fzebPEX+7tLWcWAmL2jMY4f0KQ6vrGSm5UYDwMSGZeIkDbAKxXczZGF58DAaMlfq
bHeWLLAw9aetnYHISvWl+oV5LV/kBVJXNc7kbD7+fH3YQvSRolNbl2KYbkFg7TsM
ceottWw6cRyBEPyuhVBcgAlJtjfAmy3oZHrq7g2/D1PTjjZ6vvFYi+1zg6kWMfQw
/RpGaheOmuMVkGopBCiiPFwVMWBh80SXO45u5sS67MZiiK/SQJDmoAqIUMRZq3vJ
A2hLu6YfWb3ysvOZhlobxpCL6hKWY9GycBCbt83387g7b9g05bXdyhkgYnCRe+Kj
LHStfO3l8TqjEn48EXLKgxlWGpHLtniIo6+Pp3mcdkJrfE6uR+xvWnbzxFOAAt4p
naszN1/SveIZARsyX1Ioz/sPD1bxv4DFxXcyN65Pw2gSZFFtAJnfEEE4wZ412d4Q
kijy92hEjGnGUy3pjCl2yxhn3vBizROReUUQN3Ji8pqDRSeC7SvkAVHn4kCEbBzL
Qi/6uM3YF9MkU/o5jxumwKcnHYzHG2aj66RJ1JREhXCwK39DKLiyO8f2j0VwqYJo
3rUOvmJVmAslKeF1WH9nCSEvedmTaL7hlB0zEDTXG738T+UogN8AduV5Cv0GSJxE
ugBiN40qtN7Pxl+UG642jCy4Fj9nMLi3g2VwLAMGzoOZzJBeZCl9QoARsFuD4DCb
sxvH8aCT2l22/f5G31Mo5NFCafqgstDYoxAHVq5KBGLe1zTUMwV6hNk3KE9EV2UB
F8UjqmY6iWjiX1GVFm1DK+l1Vc5WbWuLcnr/Ih+Cbr1KREazfvKzM1rvuePjTwwX
1+pg5dcjkxX4R4poiwtCq4/HzzX9pgX28xky+ajgsWsWCAslDeqWRJbCHwUrW2Tl
MTqVDvJKHi41Ce2oV23vvrsL69Cmz4tUe/q71/WXAMK4gnWGfrZTjIZk/wTWyc0a
+om1GWObkuXQXnfvWyRYWofpG1xmLi+e0cvAcQUydsXUDAMoIgwejDiePYnLDE/S
sf9eulsHlhEXXy5RmtB+4hXNmJzO1WCIWsGSZKKWzYxSN3E/AcaioqSbKRY69AOn
2LeRQfFYEsTshoWTTxCkFaKCQYgOPVXnewccGRdW6I7Xm3gB342cdCCDvnAzEN3u
L7+z+W9pwgNfT4IRas0T3lsxSYiyrVPCRRE+th31Nm6c7xQVvAqHXQvlKzyN3Bnm
MGsJ549kZ6LmUOGVnI8JXEfeKwi0sL6PcvYfVAx+mLHe22KnZGZq3uqbqSEKqvcc
Ijo6S8CNwQOBZNA33qA4asrFB0pQgGEV7zyL1CbqE0MUQ9c1h7KeYPuQbmN8zMxX
sMKmvayDrxbDBNE4U+M4rrW4+2C0j6UN/67ve1iRKKCBh5DU9XiYKgEW9Pu74pdn
548iUq2DZT+bMPK6k0VTBZXkOzAf7Z3mInDEdxHlPW9JAN3ztDLJg7+IQZd5zZvQ
dIe6IZ+avpCxDBia0kPWlwsJOtYraWLhJDP56Cd4aq1yGtBWOr7pOq+8gnz7TyWq
3rpP+AZAuTUHqgzvGyL6G1ruAKBCTKD2OyCwnlLbyCbYLuUP3pHkXlamDyoZ5rnt
Bf8GeZ0pAm7y743x5IpKj/qt4vjZZylXU4R5BujTA28Wfk8ChsLW86MqE1VIbfkn
RdlV7NkY47VrCph09QybURbwttxHRFCgsT578h1JefN3QPHNkc6IOMsiRF8iz1Hg
3LOKQYqcqaD6TY5RyWV7453jnInx9dUmdnasV0rjPWrUTkJ9l5C30bsKV5GUX/FN
net/s8UsuRUxUWetIHpEr3y6Cm4EgKdz9/K3Ji16ldOjkeKG1DLVhEbxalfFMoIz
1TYR/X+0QS4z9HeisNZzoTiGMfKWkgU5WktCThjFQfeUnk3eaBNRemkuP2eswO6b
jRJasHU7n3tx8cUI83ydwVxmuvS4nFzjoRzJ14YkGWDXS3MZneuZTq3dfdltYEKk
9c3PfbKGGEz4w1hUZ+JDXgM5/Rg+lWByHHhkigNzUZuMUGXNCeoAC3ONzt5686Ox
fLnEU3IgByYzIEBKsYdWfGyy2zTRe6LHn+vPbRoO149I+2PsOzkr4frEdc5qAj+i
daLBotSyqc7UDaNZjeVdJ4UCVW3pmHetGJSWMdMhx8bUmW9B86qtS/Xk7ksVb7OK
leSLrCsnNvE0KdHvEteRPnn+Tke4JAEUaUSmuaQVE347//UyN8NAW206ecg3HFfM
2AnFdqhWanErLPaW3StHmQjCBbBlcNCXbC0B09uSxQ7C7YUQRtXJSs1RUHrduICf
hW/3ddsinVEj9MEJ4mphI/ixw0ZwV62jv1De6kzx5t7hr0lyJlhST/ONoaMDmji7
lSpFiMbmDmo7hPAEgHSsP6pIeU39wrm1SbO9Fqjg7GOxN4J3I3wH8b/ASrt/BlTM
prwJef+1G45uY6KvIjkBbi5PVu4+HXgJ80GBb4kAdwu4MAUjlD9z1XCIgtgWsHcR
NGlMur9HPeSRWiPll2dXZRbcaL9vlgd9nE9x0852pFlxtySyKsnH7q3AOXCC5juG
WC+cmXiBl3/4YEEeZywpzHxetOZXzSvP6Vwn7zbucQ4T/v6ef1+1WECu289fnG4T
/b+YcykTZy5kt7xmvGn831l6FfuB3WNHAR+VIVPMtMDSLn/R0q2771k9wxvv8Ia2
Xb/jedtMZ11aOrve19oBtRjykrg3eu8hnWACRhWFN45y6SrfILEq26MSw6jWlkNa
b//y/Sq3QSws82OODeAyIbsUFe+b0mgKXPOYiM8nJzmFZXmQZ1zZZ7Cx9HnVCKx1
hRKWRBtzbYpkadQeSn5B8FHaW/rIC56MDgc1FCFbOAEnu0qaQmEpj59IaqA3z5we
TJh7xHeZSY86cxIkCPXj1sLVtNccQ/hZRvGyqqMVI5RVnUzGAhxJxkHl/P5V9HeI
bAPEICMHgTUQisfuFu6tkLSbmjNkWaumY6Im2Le35I2QegSq+ES+OWzNPQ1x93Yw
96ELt+orXLABPlPf3kfsxGoKuikRwPLnxsZ0s1IqewW/XQ3N+LoVmK+cBwu3oXBB
W/fQSZF3Vt+T1v/ygSiUgfR9ZoBCyfmMcnqG/U1YUfBGqLw+hC6ULwQ9GT+qbm2F
ySCLVns6BywCW0pIV+Q4uTgcDyIMdSjJ/i3n+aeYEcQTyFlDmJZphR1vvzyBPt3M
HDZsnL27eFmpL55zYYrysl1t+L0VEpvGnR01XxJsDTsouu81mEpI5X+eYugoTUNu
RTScEUGpG7vHVOnbSTkkF5bzMwUdhaIelQBp02yqAkN4I9YbpcEXjxJd298ne9b2
5Xn0D4wvHyqnAQmy3FMI8zsvFQr8jwzXeXEPzIWVStXfcKQfzd57JKudx9I0XZQh
sENy504EZno6Y8TvH4kzxebq7CcNUH4gQqeDkkiNgaLpnqer8k51d+nO6zyksnGB
7U4ZFejGuHPa/7avGni5whBSaPHbgSejFIejfTfb2ERh8xn3t0H0OtIWMot5akHd
ablxZQF7rc3Je7FfqRqCJbTmpH3c+cKRIyvdxqRGYWWTjJZEo3fUtIhRRr9Dn5rB
a5a0PhDS5eU829SHGE1SPO/Z3Wxj9OqJMUy9zc/UC4hIG/yU7FJRUfJQn8nMBBHs
RnpnMynENNBzQkDj4+2u732xhkmODfYUdQZBn/snAkWN7dD5V0qm3liOgMpr2i/x
C0pRL3C+8Q512DCyqPxDo0bWTsDxoxzLbLrsRRwVpCHkpnAtNBmwDlAQrMS5LAzX
a/ibypW49eQ5Gn+o8ywN0prU1GCmbWZnjKKRnB+ddEoPMeLspOqZebpTMNole482
vpaA6ylNsIVmi5g0tNKLx0fkeKIkaDF7kzAeArVOS0EYvsewxddPujpsdYq+DuRj
+hpVfyp+1qCxiHfCXoyu5q4u2u2kD5PiaR50X3iRmhqoRRYHBBw0K1AoPqumh6EM
2AAEaDHcZWmo+6Mqxja5EOEih/FrxtQjApuZkfg47UOvYlG4e6wEmOfYLhN4HN4J
zGgLTqrDbtqooCjxdGHlFzzkL4cJd+U7yoBNDTZ6B4ZlayfOCdGh1qA5SkN4dZXK
4GSxSdqXlwy2oM/OLyoqWYm+SqZkQmT3oIZwD50XZWDjpRVJu21bbhwhDrkI47Vq
MoSBBqzgaz71wFmQs4z4ph964jDQCNaCMmBXwv4N6nSHlI38EyV+658gjxkzZ65K
1osDF+49sd//TBvxaTTL1AvozT7BlGghwKoPH/I7aM/Sy8cJY/BhbOapKx0qUJVM
1LtFsvdYxzc5BrFoZop70Sp8f7DjTmCTOp7pJOqlzcrSDBroTp2/gEEhOT92bpmF
3Cs2DStv8SKMCxOKSMR9utqsCo5DWJz2kGUw75zM6iJ0ge/keZG5WdMfPiCcIXcX
aCAIce4KJV6wop368MerZM4JMXxUiStVa1jKmLEZIP5jWzF3NnxLJ9RINDNb5+3e
Rz0LpOS5VoxTvJ03REBzk1ZZ5Bc+urOT+KVfmgCrswSO+lQw9nKzUy22dPhcPvzJ
tL3sriSVURHvJGogehi02HbNPCmBMxsTL2/jCpJmQn7zYnK/ET6GW0nYopViMz3r
Ee1QqWCHZEr+ptyRdm9gOumc1JqdW3VoUSNhoCtC6XD/yndXGLW2bfV4Mx76V9c2
PfPit98CFCi9h+yWbiQYMdJkOulIbYCubYsRLMGTBQCXIsmLv0CD2eUfq2Tj83vz
IBd+BeeToYQ+bMiZccfRsxJiBq8EtdSL8MRfVrwJuwEOt2d4EwPDlPupnT2tbxUW
E9KWAv/1sbjCeg44wIFWiqZpJAaA8hFtKAQyh6sWIUmaVu1k9TvkIsI9ihiFAp8E
XbbO8fSAqdcq3fyJxexqzPPAKpF9qmtBD15GvCiq/DEdPs57M1Lu0nkCgGWT3gjh
TFoYIUXsH0ZiS4tW6Z+oQWZ/jepIRILncj7WiKx9z2Wj5JJnXh9iTNoNg2YfSGnw
ddTUgsSCPpPzOupjUutWTw5ETGM2bYYzcuE1/IqhU3yfrxn7Bhs/to4NAi77EMUB
3Y2oIiIDtK+HF3wfu+9LwrLbPiqfFRSuOAccE6S06kbkWhWBDsoV5rpeYFy5vI3Q
vO5irkgwOHpaZkFsZSQDiWxbsFVHBR54Xlw52iuhOqhRj2df0M2CT9IVa56Z5T4S
aumI0XajeFyIJQehd4BAHXonny4ETMX2m6EexONsIWMYN2iNykN5hDNiIuuYT9IZ
M6iNa6C4JC7pOzQ5bg4kEgbIGtiBswzyqn7T8AO/k4HPZYnQWuvJmzFy6LB8rHdX
5JdY20VB8uFpQzTa3ewMsuBOKI1ewAziHUbFmzCPJFNpR8WIThf21gIszz/j8Jpz
fXKcD9gx8+YcAyTTyK1F1CAyvwSx3wqaCedhLI2Sqh0H03yAlo+WRffuctF9DUSO
pXauS+NZRkj9RPIf0vuwI9RwuCNuIu+HCvZlwdFy4LafM/IW8r03UPgAgwB/a5N7
vvb+TgQ5qUiCHFa46Nn1DqhDB/VAMWGf0/InVlv2qaXAAaP9Z33g/dUDdYIP5dxH
48ItGRYQd4wb63kfWOeumkaqP0ZLAg8hb+NLz2JdJpe3PAe83qOCancsdf6fqPR1
EMAZZOpig2sZtGvvAw4HJqEKEJtR0xR90Zg9wMeFqRNZFUcTLzxds6FudgKAZKXP
4SQqrraiwGWcfnnMRhawLkBgLchlOMyqn+hK81VQLD3CZr8ilTkhTO3rTczM6YIY
poJJM2Rho+hm8CZ9RQtXnHi35YQnnqmpIlmwlfC8ge1VhCR4AvRp4xn92MV9Ixg1
Q+zGn52uT6Z0aI50njlZy326qB9++f0sSBAuvXUy6hl6eL5ui2Mo3Ng4FUyyVeSS
IFe+DPUWeWsS6NRyDLvJJCkXKFL7Meuh9nt8YX9D9T/TQaEcaTBSjyd+77ux6UFK
BWwLRkLFdE+NWqN1lQ9RJKB02CGxKDh/XT/3yYhzRSdVTQ/KyDB4uo6XbJgTwSZk
QZfsm+CaZK6KEgTR1trJn9OOuk8rDQrTUqczOSH8uljaQDkc6ZHhJu1zlbMeb50e
YWLktPGwlLUaickub6iH4QQyTCPdGym67b6Z9+AO+htFLqqsTwchnQC7bTLYm983
au4AStrI8QzERtfleRs0uGIFkSIo0BSCbMm0wszzBQMpjlqZUtPN82NfGxQAuCp/
6Yjg4kJJ3zXt06c5SAagf4gx0c6oY3E2YkPWY1JKq9cFo1voGJgdD820kOkceIYB
W72fCuF8VVmjRwzC1DoIut2Bw6GxD6fC7c80Kv/k5QyM9jj6wER6ivc0ZKBD1qh0
E/cSGw8HF0Pu++iM3K6DYIZLl2O4+ShzpHU2+h2MxXymYF2G7PKcWJ12o2uI5NYT
1KduZ17G3DzI49fwnsJ2CNRDjnziRYaL3m7fqnPsK0L5npmdSf4oGMN3AlZ017Yu
QR2SYxcnYALK6wfSDxw9T7RVlZ6CjIv/zx8701Fq4OZdwAvweGOPeZt/YxBdlQuF
FfMT/bS38Ua/Y1kBHUbhHgDNQZPnE1wi/VeGBhHj3mCCvZYtO1RC+mhk3v7S4cxF
5aLkGlEo+vD1YMIH3Ro3fxCNapmDIqo2GmBvBtwE4uVLi+hg566HyuqW1cY779FO
peGQyvH07OG6AJR7CMPpUvB9nqZYePBT9ZvR2GJ9FrCyrqQ/qqSrzyeYbXXZ0n6I
zJfoIKvD51zhW0WRw5XfLpkU1f+Cr+GXMaxJw9cUyTjxEDoJufe9j+Mx+sfwX4Gx
prDidXtH0xnwpSF+lcCirh5/UoXjISoQMML2sL3LlV0gW5fw3rHKiuWezOiLawQT
YdItaJScx9nHhLSSQWgKodfWyhVQosnCrgUc1821xqhjxzaMrXjo40bBW+dvD4Hk
cfWsYg5KIvfI8N7KoSN4WyIoT3ZsXFzUWpQKqVofyePqii2rPujYQih4T8W08H9X
RPRVj1hytHpdRkljBS6WCSZmltboa0mFUdatKC1qgnELLAIn5XuEAtJ3ZqrbS/eK
ayjJj/c53CUYw1J/YHHbXv5iGcMlHRMWyoA8sjsHiKhA9qSPcYAtbxR/h4qL/5QD
akQ+IuaDkdflSWb+k1nWFO5i93QVrWCuUunBjcbAbyYJL34niwi0jdjpRE3k65Ul
G8kL08dVzLl6z9YjanDn1zn5ZqmbMIuFAbtT2d2q0Fa7ljgpAm8C2u7d9jUwgWEA
jSjv10zWv7Yvx20SpCmgqRA7bfF01txln2vsnKxTPR/2yiRuWgVMRxA6I5c3EPpa
UO7JK8yIgZskc3K4A3ZopXMN1PTwvCMdTGiEVikKgPErMLTbqrAJ6hM3f0+sisMe
7uyPs40y+GljzLzznUkeWyWTL9J61kyiPf+f7yNITSnaTPFFAb/5aZjVhwzT0Vze
4cg1qQhJGIAl8/0ZS7Qx1F33WGkOVDKVAT9lcYziS+RHlFmD9d4DxR8qzCSgt3pB
zSTBIIiz6FrsSrrnzaGUXCc0sJTevuTey3QIkbY/JDw7NfMKGDPFm+LT4Agzzpk9
qbfPZYlg1cw2ylEAJkPssYWw6us8pjdIBHruNetsa9JGYfsCrCEyQXOqDL1KFiva
7y/n1AuV6IkIQ38frq0ccls9ZVclXZdydXFFYuOKJbtk7cdFWf63XXUBFWmc9MMu
0lKHDpYX3hYTzL3PnUA+Y9nFcCLzJsfHbBi+ttyThG64xzGEmwJslUp/qL7N0KFP
beceh3cX+bXjwSh/w+S2T85H4zFmZ7LRP8kgrSwodiQ6gmTLemwL8zl+VHjPbtTz
ObWPR88lyLZ2rV6CpETfFv/dR2Ezi7qo2kzxiBcaxcEnvAvBpLO1Aba6B1s/NexL
MA1FSfNq+L9F06BUMQVxzp9SObZZE1wXrs9OlEvcWp5IHmpRn57JhyyrpEl+sqvN
EHDUdUeH3Sk94oH6JLCpkW4uvkVEcV0szS//ATj+tdh+AGv5ITA0uxn7Vk80WDBp
qT70RzUO+f9vf/ZughmASyGpNuikO9wxYGXdoS1BS/Lu/mFtOLRPG3o56w/YWWEK
rnpJlHKnGtDsW1XjhUMw+STHR4CstVqFIeY33bUrQxkSKsTynmlyibvDqcjS0rgq
MPHcwr+WsMWjfCpZcWtcvnpzqV59drSMRiwJwfHNFImOr+3nZQco3tj6RhYU+MCa
dOWbv6IuO7X205/J7JzOCR8VDBSgcynbb2k6/q4dzubk4WZtrh8vf5Pf08bFeuP6
PRAt+DEXrTh7C8tY0ahN7+iePQnMQorF5/6oWgmuqFqwSXQfrCEPx51wIJRv0jOH
ulZihrS/0EuSPeTz/GJS1dAiRwcWkGBfiZu3ZRMow7xUWP3yoZ583wnEvVsD34D4
SjVSE437xaYTbeppv4rBMqJQz4cpPnuZl+PrO4n+ygH7U6iXtgIzXbcrI4N11bZn
5UfwspRbiz23YV9dAyRALDmPBposaomXkDynDkP8quu2OON87qumDkW+bujKoYU2
4yfS1aklwdRn04vjjOvKzWidJc3QumjH2hu1JXr/vWqxTtLG1jvT3QP26TkskhQi
KE+xM7HX14h/EGcWkpun3jNuac4phwMCneetWpahI6OH3XuHlUG2R1oYYxgPqZLG
EOcTlbr2hWixpQSUN0gIJW4nuNgH2Bik0MM+AlRKhGK7qetWWx84IumQR0Thy8Hm
hVqXMS5Us7fnamDMkUbHT+iftE/dOLx7BC6xCdszZt41kYf36RNC7+7XJSS235rM
uUvLvx9goZs6g/9VD9y0DzzpfSHj3UM1GnetQgyuBo/fWh09tRaccfiLFWJk49h+
cIhDnGC4zD9SR+iVJGatP8L0kSIhSRplyPK0xRL6kx7nI7P/ZPUKIRDr85GXlMKG
O1xJ60qS0p9TAlF5Xuez7sChltqB9oMDiyjh13293fR17inzwCBmSMHjidYsYB7+
piGiHvW97ye56EvhuLqJNmwDkOPRowxmo4Xwat1xkR3680ALV6MHirVAN7TNSjFC
lrVvvNOMJpzd60TIgK8f370w5igyC6/PUreRrTN0/GgskdTWIVdq/yHro+cZYZrC
uiQke4938W0qRX/uIoUECB3P26FihgEi0H7HJhdqJBgenC6m3yorWKEbxAUMr7aK
3AobooKymkpazmgbeLsudPClVuAG1hz/bKlxaJEnPuhgrqnvXYfCI5yBQjfDZbh2
tnf8gMXkbmdqqgHMqwkDAajbdpSzdWMj/M+/ONnSOc2sRL1FpnlZeYvZMut0NTGV
1/nID24C/hc8/dn1J0TUvwaM20LoC+RAD6kN0DeEguG1oS1GctFIM/izic6mgF3s
V18zlBjOyFDoVdJ7ngMfKJ8CGkq6itJE7zIZ0td6a5KCE6gTQjueabHOqYJcAWDa
nX+c520XRsQUVTEGspPLZo0wS2PO5loEK2OpHF0Nsbn/LU8PXiRvbHtwUKBrxcop
unjVzPyaGbFHmFBk4m1rJv+zpzaSG4lPJdlQ32Xv2fvGpcYmvnWWHOsEEqdLpotv
tZRjkSeVzDOjd1eZ3MCuS4t+pegzXSi6ZOvPM4gbfgbTA+2xi9b7ZoH3ZHgBctcR
doGvQhcv+Ou+uB3bCG8q477cc0S/4AQ2rhXnYwKoSaMDXoK13BqrjkoSlAZPDrUD
wrnMF7ua9c/Kc0jEXasaUo2lreOGBICPMVTC6vkC+Y6+4nOQELrr0AEYBKS3Uyh2
68YR5ieIAZ35dUwnff76kv3qJHY+0RS9lAzRRLfYlzybdKw08YcGeV2jhggpgclm
Qs/bAXUFU21QicVSJbmgJgGSSzb25ltbn2oFNpiFFMxVAny7dOFA/n+/UrSMZpfw
NRlrjSI1Bd4QI61TRiFr59mCJ6lIXqv1J3hl68T2bQaysUn9Diz+pejKcvlIL1xh
JJeF68D0v0unElNOUljtZAsJdrGqU2DMxFd2qyRO+c+yyL7ZprIVY8OYQTaRTVa+
GSH4qSNtxmKeQeiCnXRx3MLHxRXg2/U/wfNIRNF31KoAeL1dn7pd+w9m27sWXou0
QI2/XBYcqoP+AthCc0t9CK7w/D/XqelRfKTWs1iJWm45FHnn9BTCt7f82xShZynh
Qn2uDTySm/MgTarJEJuX/faJl0D/xP6991NVJjJ6rIFL+5BHTwgbmUT7yhfUW93D
FTX0BuPfDknjZvIpyhVDY54FZm+4IuaVypDQt6dHKhtAaglscJ/bNsVPM0/O7Kia
LaAs5zuAELwwoROhOdwAl7wgzc9aTe6r6q54bP6/gEDNq2C4Ci2490l98NZ4RX2I
8Omw3GRsdbKPeR6GaqD9OMYALE+3q/55xGlhuS1KcRQOaFP8jYr4WKOHFuHA6FS2
CARl59OVpAQ8aQXh118ErNUq4SjdsupBk5JNdGdtcKyWFckRY8VGx2t9vfkD7EO0
AZdgEncCc3MZgFMkKy2wpDdqzB2euK4xjqYZEgM+841IOfdT/LwMCzRwfiA+noDj
uUDKJmRM9emNAf8RcOAaBHCR/45xrRIvxK3R43/a/LBXrwOle545PA6U82N9nBwg
h9KSuhNDRMjL12/lxWapVMlMUaz7fky/rWAhHTaCuwvoz+qocPFrfqdj+cIJnPS7
6Kp3e5356NiF5c1PXy+rPll/rnrrAu1RmZooCrMqv2oF2HXw1ouVv9DtF1AhTL1E
C+eXHuFgzU6itFr42nGWltE9MGzYUtGgZ9plB0N7jOxTQDHeRnNMgmpY9TzmSjLt
jSPdekeBU8Z/1jQXKfro2zrlo0RDTcY7+N6TbhTdZ1V+GrqcpBQQRaNGf3stVByf
RQYV6FEtTOPlZoFrTI8cyHcd//Pmi00xRClGy15YvBlpAXaLV9gAYNOzTmuHpdJW
4deyMuB3T0Yuaz11mMP53dnXaLkoVbqvf2pKHUn2MXZqyPYvEN4JmoU7Mk5WKJGY
mr0S8KsjIgJ3W2JY+KGIsbeMYLQVwK7cNBXQK3/zyCEdKv8HBhdPQxPcJY8aknsM
QmUjAk09jdBZlbyWxzHZnv5KMJiYQSZBMzVwwNxyeG9rIlQdOUrQPjd1mf/OEviJ
MfbKGlwcIosfz0zBoysANPZwdCP7LNwzMuBBRmoqeZhs1b+mGRSrNQfkAd2P58Fm
t2m8fAfvzn/FZiQvXMABhIUcPaSFOc3TaxdWSlbcF3nGaq0CII+PZQuau5azSNfU
xaW13T2JMF75DzLta2CvN5mwOeZNxvwQWYD+9/k6ezTnRy0+pTLysSbAlKVi3gzZ
zVcHAb9lAhzNcexdeW3g3Fc80mP/UHTVyNAFagfgnpiSk52XyuCQLAU5DOtxOHdr
f7FBWYCWmpDD8Ci4bDSuV+I453hILMKWLbw0MyvAnW5exAAoHXqT5bcCfWkwU4Uf
9YY57w7UCz1jQBCD94yKBRydUsW5XYrekuNoFMm2EzzGZACdR70WKJUHeIUQdYKb
AKKFTk+KHB+X4hobO7yNQ15NaZnhb58qDGanhwuHitL4ZukvQhmHTAnRXAPQwwqk
fR3Vc/PwzMHSl3Q2rReoGxET8GXfyuLXJ1UQch7riJE43JxjDMEuHk+yLlNCnZJP
LC1qpZ/eMSHcEi0B7P6m5InnymGYCJW6nZzp54P6p3Kiq5Iby+Yamw9i5BNxwQK7
44T7Kq13UQmlPp77HfK9fQi0CduF0cRTpzzhwmCEYeXcCEj1/nW7F7YM18ErG/Em
QCLmk81UGxHL3K0r2xV5ark1wVm+5BSMBxNBzfmAQSiN14wCLmx+PjPzEy8OGiQ4
HnTRV0v8K6YBfhT3BSS0SaQGHhFfXGeS+DzFK12wYCpL4bMM6uU9PcaH7TDKJ3bl
kaifzCoMqBe48bAaem2CdPA0ecSuejfG0mHNbyFydw6pDPRQ6BbtCH0ViUSOqGx7
aJiMuntLY6PyWaRiKptTshl/zLP4hlgdjruUk2g+cvUTHz0WFCeG5ubXoRY/Eqco
610lZmD/vky5/vD3uWFMZ8njJYgKC8/jh+ZvASFY0zTICMmVuMBnEpS7MMVx9qQb
EQ2Ei5+qR/2q2ck8plmJg0c/aZ3KGpdAdHdGLSCERodygucd0pIyUCHk8+6aODFK
YxTDAqjbmqWGK21eYebYjbKqG8D+pxpjrur3qQKf8iK0MS3tRJ5U+GLwbRCu7W1q
Gau9amLB8BgnByGLH3iBZRk+uSG2FhQoPsbszJanF9D1c+omSxlxOT9c9k17QUzG
LLYEzmA+l0DvMTwcHFrdQOf31g6h+MFdnYxneDXKjXhfJ/IhkjdmZvRQdiASvnf9
1ffaE+vvvkbHEkK9xa/aZ/OE1woHMQB5Jk5Z0u1CwaZP/EOSHum+FiSCyyCX7Ti2
4/JzxulqhMB/FZK9iUUm1TGFPPnAf9NbmAnObIAUBfmGYucnb2oIKjlQ2pRTh4B5
SiMapCGTP9uZPMtsMzUEm5juKoLoTnECp79r4SVHlfNKZpq1xEQKH24QvwXLBuwG
sLX7S298rstLOrRvCvNCIncsebsSwZNblGKgViA0lk9twUmiCRv8VeyggO1GQBTC
JkdSSSp0M8ADosjI7bX5jMv8FPnfoMa6NmKPu+fup+ndkI5quTIkW5olDSINtzHm
K23csYx2YRKo+FbsI37FXB4xPB7KKWnNJqIHj/6ZRQ8C9nVUsLiHm5Tjym9fvQxz
4HaOee1JSdIvl+LNqAxgEcaXU9pOF/Gmokrl1bO0xpHMD3V+n0fvbc9DwbGfAWEC
6+cpSLToOwHuSWiYLmEutMgJxHXxjOmfUvhKDj9RIG/7agz90JgbByP4ST645flB
brETg1CzquDRjmk+yYKc093j5e7TLT4dg292piaQvlhncV69vPitQdP+aFcswo75
2Cg+5LbVJJn+3GxtM9QjSnUMVcITINlB7o23EyBle3T5HiEyloroILvOt5YJSLrq
LCeJALW8isapITtBR1YpVxloHtSHwtpqtptkz8Hzrv2Po2WtVFJ1JnyVDnJxn2Wn
vYs3TIY1cQlutQQvCey0K67vpcvCgYpDPKwg3r8yTAQHcApBn0bbzRjfhACrUcS/
QQlbmqQCHL/O6BbdcEFYz785eX2XG3iLtgpx4t1LN7J9esHgMtBEpDzymfHt3yhy
xxyf6xTUJK/4TQuqGB8SXecAwHlmasFHouPVPubZeb0NGRfaOcm++7D/mmvTb5uB
Q4WI4H8XRgxr5o/Raj5Nfv2QdW4+FoYGcgG3L8+YdVbP5PT4E8IKHbsY89wsW1Fm
50PuCaBmqSHGpu2h4bgts+r0P2hMC2N/nV3pA/maYtSv5n/joqRauwM2FD7Hzfoj
vSdQtNpQc8pvYmsMxQhvFpovgggRpwUo5z6dmzs3AQVOQvP47Mbgn5u4mVycEOUK
Lspwx8KjFrqtYvIGkaFPcK6MmR5a6gs0gJluDeAIjT++3nmXXc8VAzR2s0r5umfs
pgRhX7CP5krcRFog6Cms4y4LfjiMeA7K1FcJZuJ/6kv+xhyfgAO8rw/Hn5u2M5MF
D8MwnE/2Yy0Dav5XbUAyC7RNrRXnfLlw2DfzAfYAVzW0xF8+2wnV58TzVzTrca0b
L3//Y6tKd+tT7F5sGPKB3ttdj+flCtz/MMp553a4lf/TJuuiv52uXP+mum9wQ6Yx
9h3l7YiQGZBRbkeapoenahggzvc4OJsjXz94JRX4NHOrDiAUG3V/tF2KTRNXpOy5
WPou0DI9ie+6oeEPqS2EbPTBaNnKUpzTvqKYP4sW2Jvn7ZUCsV1lGwhpjoyVaxTg
m9WFrMGowgmuoF7v3Gh3cFot76/gfX5VMKcd3ZFU2yZBNkDG7sMwR46X//L6WBbV
93yEHeAcdJFYQTkyaWRTgEdJa2jYady2PXqIEASzfqewDMabruPmBumjrg3RFKaB
TXdR1X2zTk2D2+7NTx8tQsNXKEjoM7DOoacvghrY1795fjfZC+F7J9/P3sVQo7zS
0Xp42ar4hEMK/BAk0iuFMmiyUNmpihUZXPXyunH9EIX/Hop6hIrvNz+qNhXR96/X
HrjbsQBp6amX/cgeEvtbQWs6jNHhXDM7FOY+91YU8ilsz7vEilsmGj/smJbzg1cO
+HblH/6BPd19YSffbEiATwPvSf+zzFCutsVDhlzi1zsUFw2B3BR277YDeiWrl6HZ
CwEGqE4WfBz42N06U+BmrRNRdrWmCCfnLCSCgagZux3Kj+iw4IObI0W9FvODMe5T
I/rJpdVykQdpOzwHcvHhrebcOxszJSQ+BdJo5YTdKHgcr9qqWczLVIcjwB25fwDU
ypq3FbnzqJ+BacnY9rlWdGwaatApvuviEoI23C7BZvFSpy6ngUnc2eiTGytOnQwb
hQUmGq5jZGWquhrR3GO3AA==
`pragma protect end_protected
