// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YUdM3yYr3WfZ19QRsGvM7BAfnjf3RKUAmpX2FaGmCLEDwTDR5Ra630BiE4FnojKQ
fn0xB0765ydAvEpDtrvTprKgY6gIbH3uF+EV1Hde4exe+7CLw9NecS5nFbRnhhfF
wTBrRX1N3XQ9VuKq1ygBcZ3lYAYNkg5GgbOQLZFZfK4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1552)
9+yeslS9yWK1QPMTygm2HCXTSj8LX6QjdB02aUDb0m32ar/oK7iZbicIKzBpyK9n
dBv3IaSucl8lawcMt2FkohiDXU9XntuupgDHCAeUIrXLgmeZqmxo4iNFKeLtwQR3
tKjAeaaVKl7awEjCmiIQoZFVSW0zyLUBc5eAOMX5SFPluMj4IEVNRwWXzFsr4jzX
5iIoznqY7ugldzK4rQqmC1llkChCoyvKkAt5jnt8NYK3ROMbbcTWUIQwBzm2/RRD
EXkWjZ7NpSotswJaUmRLEV3mIyrxMWDcpyi3sXqVDWtw+3xklC1pfv5wTsk/iGi6
KYr2NFEPq1BmrMyAZsrkJkuMnrvk0dKE05w1fMKo25FJA/cLcKixCCzYQtMikKww
B0oiLPT19gUNTcRHjHD0QV1QLzHj34REIOtjmZbwUK+3CJK1NmFDD9e075h+rJ/C
x7iMB+6pc3WJImeB8uZG+fRwAEdaTfZsLQWi4HZO1fijeoxx44UniQ0W5EaoPw0H
NQjMiImCrTLVijyI6LqWP1JoGC4gNI9Xe4H2JivcIMxV5f7e7+HCaur+pSHPzjy+
BhodZb0Q9aBb7E+bq9trCy3dXa2PIKI5ijIQlQqEXQGey2sHz7fHuoOsHzNnJsmp
u/453SRKTFVUXuuMvNS5n8kJQlHwxezJwNFbdlwpRXr8mgscSbp//M0mCrgy77U3
hydROn8Vabj9C7w6piUM1nAvOzQjauCb+8zoI3jD+WWOsKyZf22mZijJWgccg3Le
gQZ3jDpXHdiirIqxxR5LBKCyP/2+l4IYfkk2+Rhov5eJ743xpZwL/rhKHJE0ljvQ
T1Rj1c68VD6z11Ba8UUDWRbxCE05qDSwSRtNMzStDDROCSLgSsCOVxHgz4elOs7R
79E2HDAr36g3Xk8JKD31JcyXIioljH92xSfEsLDyIOb3PM+AEv0x4DWbWwPyeTtz
nn8eTro0ySNiCTbqbuYIK82xKvxfhQeL6oIjdAVnB9r8mdLNxiwBnlKFT1oTvQ68
YQqNpGbMSoTKCCnneR9PwCK1ReW0wLDYvu5xgPI6JdHvbrNu/OxtcGobTAzkWTAV
r55Og0qev80X+ue37lEXAuRcv1p9dSV70+9Mwv+nFtlAvvn5rE++sxfZ4nHqTtGx
/ElJlagh8pU9yi8879dsMRKQj9OeFQ0C8kCU4xFd8qCQH8/KZVsr68wMFZB08fHY
CokXINnhI8tNxXj83zM04OKT04X0C9sXP95+3NpArQiazZFHgkK5/QzFHNuQCTnE
AwEoiG53viyrI5F7SX0+//+MN/xdwtgIGjqfMOPHjX97RYJKVIhJ/HWDduCirSSN
X7a5gvQ4IywQYOOU7jshUTSx6XmLKgMFbgNgTVfqKXde1YkyeATe94AiSBGwdxCQ
76FTbLSqX7od5r9/zYbaP/ojxMFsVE209miixJIEeLnbh1ZqcP3MmQ1EoqzEK8fR
sCptCVxgSvYarJxdod6ka8tlurNDcUBoGTXap9FcU83YYBnFmseMQcYGtlgFjXkn
Mw8BZpx1TVUrTg+RWIoIMN+QrhdY4/5BYgfEsBAbJz/hZWq2hxTrq2COcyuEFS3w
fRdxMEJeGme7Z1cPJLmGRTnYFpy9huKrwsQdwguxeseU3HjC5+NSFNMa4RRWVP6C
Tf+lhyXHGFF/5jnyyXyoOEduDVUEgKA4QA7lXibkXydm4FXTkn1gRL9GQhgCvUNr
yQudd8fFOCBjYIdHJgIVeKhg6Q78xyu82pkPJsWDD+RkmHXR/Hma8YuVAfQfrE4F
EEeNmL2VsfRJB1b27ZOC/e865IuX1BDIhFi/XfrQcS/oTMUxJ+rHRlLLeTAi12Fe
dWOzF4p1nkdkpPxASmKxXr1EeiWiSjIbgO8lP3Btn4cy4RWwl4G6+ooGscwh5WlG
brYBTaid3EccOS9SdPRYWR4F1o5FhYriib7VAx9zg4IaWYpRK/m/Sxj5EFVaDBdH
huX/wUa4KxZyFdsfDsy9uXTeuTmG7wWWj8p65yPMrGDQcl5KNV1xxUa8rAkdDzDg
NVuQ4QhjD7su7GwebS4OPw==
`pragma protect end_protected
