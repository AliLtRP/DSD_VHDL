// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fejEVRrDha5/7Z4q2y79GIV4Mu6AAbNMy6djjbFepoXlgzcS+XbhyRlkxE+/JcJy
jqy77/OUOkmsvY/gb1Wx5+3H7LV7wwo0yuGOZ/NdGZmhheZiChWqDsPLnmWhq5J6
wkgMDMU2RN+K6NGDSvn5ySKPpPAo8sLl43uD+YaoQQo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27920)
aR5jYeb59v2fQlb6c35+FQbt5RbkGFP82aZ32fClIbr22EqbxU6p3JwxP1KSFpdn
7R2jLvTeoWgdMA32tWvCvIAkMtDh500JdFwjBJSiDDiocT7Dpmx0/Z4hWx7JszC0
D/Rb0lsdSeLyUgI4y6KRrleYUco7VwvpGGk3b2wn+mHBt31YCd5yUUsveXy0pcR1
ofrYW9ePakDGj1ronf6cL+xezZk3RVWuI7VEBbEZlOCXx7O4wK/XUHf7TRuNk1fU
XrRqdJEoeRGWBhrYi7EDwe90R+hOrG+HAsu/OHAGWPTol12gSchyHJ0ML5PxcjDm
Uwfy1dbVdDf1pPUie9dISGjqM7qGy1JEBustg+GCpahdiMUlG2JeoPjwRcWQSSbi
6/ySblbRtNFk8H3vUQB23xNyuKexf+V6/bfMDGShORJio5fav3hxuS0Sn6Kp8+8V
53vVXUndl7j922KkrJEMZNQYm9MbIz//pzfqBSZZ8EhJLXT+qMHuOwivoN34tmEg
ETMJJgr0n7nO4lVCABpp1OAkhsdDrxPuporsNLF4dR69xNv1QtnUT2l0o6CSUGwx
73QegziOue+2xBYnNRMyoIOuKLa351Nulg2lm/FxAIJzjjbIBkkW+2gr9rxErd+N
PEHEuk3R3kKliAcwcTb+vHkTg6T+Aj/Tbji8ZnwQquuIS/lix8uIdUrfC+SjQDwO
fF4LHvhOqH7cyVgodkKcQEVazrNMM6ZLdgTKXgZEq69C95qpfFpUUdt5BeC39Ag6
oHIAv+K9nDtGLQcP5nuWmbTyDy/SEJkxX7p7SzHkSS0uX4M6e67s4D5/8doixVaa
9QXcVAIeufDdN3nJKd8YBbSM+UDTk+mkb+zdgwI+3gbBhTke5nOnwN2haYJ7YAkT
hEq6O0QDdroQnehGAWsBkC0QM6Y6VvdmuuxFYpr+VX2h1VgR+OtTTlpibdf3XzBJ
A6BSmaHWWTQXaAh+6bxp2KWZLsIUH3AWzG/2SXERQGDwHs5AfeXU0iGv2QA1dU6n
D5thX+lZ+5sB7ZUIV88TxRfkJB/U82+Bwp9WDKT2YQNeLfrYyh3m4PltH5z55XaR
3bFQwFdWTpOwG12EJMOQvk72UxQVYPa9lmsRGM0G5T0tFEjfDM3w9UhjFSKamXpw
bnG3+J455+QV8GMPjHSgNnALMomIwxROoJJ0ZtXlvrCNBR3LCXvJCd8YeBUNDbpc
mxPwngiwVEyWHfTX3MYwsb9pfJacTnIfdi/L8/m405eB1xQ2oU0wOaVmngpU5nRM
n+qMnvJEc9ERNrpTe3k7aRKrKKflB2P3WH2BCJBLA/ljn4tOYd7xqoDBr3USJ2UR
7WtGiz6H+Wh84j+sOzHhEc3VdLnn0/YM4QcGna1Hdjq4WT2HTTg5cqlPF7xhXXbn
4Ez9EfpyI80j3eqrPTotb9Wc55wApeeTt2SzG9ld7b6k0onD+8Vy2/hFhs2wIglI
q7KATpkDKxEl1aucyUc5EdlPUclD/9vNDGENEZhy90baZHHPMxUA+cLXMx+AnA0F
9PVSUXvSdOeCQR/Xz9rajJFtyxyh/k+t4AxLbT2PHYJyMxCBn5Q8lh7PG5/e0yps
mosXgICdgB5eln4FWVP7H7GFACrndpF3BnGfGUrX492ZXY+rzYXwquooNVCZWnSa
OeMl54/QNpXeYixi46Y/2UQaYXvEyrUblJW9zOfWAN0KDjNjAjtng3LYkzNnEqqd
36O2QA165e7LwcQ2+f03g1NrBgeD2UHlo+gH/GKQlOPd49HlGGHV5Z8ZQr8BBLXI
sbz5Xpw+884wXznIs4ABjQuQaJFEy40V3q2nzz7rwDrHMvx6deE1OzFINJ0a3RvE
IIWmJuWu78D8m8+CPmpp/8XA7Ds9+2aBr8XhV96fyV1CVGyXYajcfm3/ZnASKHaX
sK3TiukuSgpd6UO6JTaSW//CFtSrkbx/ki75VkBwYT7GX62E2GWjRox+EaTFH9Nt
G4A8LOQv8XGQrrNjcniUKREV93M5+QH7YjqL3QFHHacA71Q9Dr5gfGDknvOhVQ0R
UEpcmRh5rTYkpzG78IOecDk6Krciw6KvQ3weVooMCu2q39NCEgo83ECZlta7vjQM
ZglIy2QU79JdfrJwKekYvrR/HCNobZ+lgzf7CD0OIA3sp8O8heD69/nQvardViVO
UNLqVLyR395Me+QlxHJ+hi5LpYplWta8IWO4Ivqmjh4wI98wOWmv2KYepSaLJkTD
+h0HJUTf3MY7DNy1iZXTbz6D+9JphgdRfOxoiShkDz6mK3HPTJvfyFIzpl3aN+wl
pBbuVUzWWgJiO/9AH/NIYzCRGtH4hNDpk6YirLjHJy4dcfMgk7DJJvDEoooDH8Rq
ADEKoYLwmJOVVll2DKlgpK1HtjCweIldZUKz8RZZY891w/IYEGdXfY+l8hqsdOAb
TJKAOPQKv376sBhYbgzgKIYKazPHTJiRz0+JYdzO3v3njMKUobLJl8k7MCu1YLAa
7wHmxrqF9PTZm4+QrJmEhDuSxLItJiy+mpMgmrpdMtw7U/R5cxPimfLJzzRdICUX
WFjVI6jOh90Th2bbkrVCmCkKGMQaSpsPjDzYopokckF+vTIrUHDeiIMlEJTUgcxs
CMwNIVvolwE6L13h/1a6D5WE1JQ311x4I+aWU9ySJMV1yWGjdmvfcIyro5hEY//7
Adn2Z8PG5iAu9nocg326PbCPFdVfRwxsA2t9Gbp8lFzNwnoogadt1b4V/A8Dd315
4r1010O+AA2AcrOk08sazx+fLKV2wBSCEiYddsb81BOfquQ+fPTOdTql+dSXyErV
HKCMisq5p+NvmvJ6XQLri/j6/lqafMKrpWxMpL5aZS0lVeV8Fbs9Cd/3/4QJfchk
rO2Jg39b4I1hUTVW2RbgmRvSdWrH5Cfjf+jzS8K7YaL+bwMmJmS8G6nwBpBqL5g5
aYI7Z7lxhN+4+Xn3psGEqfN5eX00pPOmRDi5XBs8AWkwMvg7E+8cKpv0Qt3cEw40
4vwOAUFy3vtyIgXVmfAcYpUamL+yZYFW2ZXLtXcqb2d6YfT1telJckMD8USbTK8P
femAl7WfolaXS808yiUvhk9+tV2mvcAZurToGenjQitcwFTOPp60KRmGnLzYgH/x
d8DXBVfe8eCVQoxxWbNTdSRHRHLcpPFsO7F0fznBgflR6D9YBLT4vLQuAAkP1anQ
mBfdjp+kWJtaEtSpyWcqhp+f4cNasiGawgFvIj8+beMPD+HHjb7p6r91pL4WsYi6
6G6/DxkYL35LFz2d5i5QLa0DX22ZSSY/uogW4w6MlwNckqKa8zXwMDRBrSpmlyYb
RNDxkNoaX7n+muZr8BHXWnLzkwrji3v+XOTwwaHhfGD9WNlwfyqbEvqExcE3PMdT
P386ArrM9c07I6tVfyA+U+XSmeqfCFUjYLT8Fvt8mQ7PcRQ38/FXcVMtgfC3Axsk
yyf3u45aJbnlsn8e3SWQd8kLiq5kfi+bx25s3MtKgUBs2RaxcxJXvAVusfpuck2v
pWckHDSKBQzH5jg5B+QyC7gnQslLuNSLbHB1WzdDJMArGLtUyo8am/Fs7YbNAF1A
wtXnLDDlsfdPn9wDga8ddMEQrWv4uqNwnZKEkHf32I3avwMgwj4UmZkCNjZEAKBw
JXluW5wjAWId8R2Zf10gUK7smjf/Er4IFoHSjuIUUAIZo0uMyWn0/lOKlwQZSHKz
ICgCw6o9wwakRKPAnEldMUo+tAS9XTS74vNaqyOrRKATQ9YpI8xRzLAiq0en4SM4
le0cSPVM5ZPk63Ne+oj3SXChdUYeFSyWl16C7QB6+N3EegmLHNao2fTNKCHCyCTD
T5gzXf5XxMTkuBSsUxfOxi8XqNxOO75YI0y0qEpHjbSrCyq9saMIpUh0KctAJv0F
Zs7CZQj/WF6HiYNPORXn7vV7LAT4opcf2GvxYYWb3Ee/Ny4oxTZeoI9rC1VT36PF
ZY01dL+qxhOTe6mrxZxTDqBQrBRb62Q0pPEwK5D8yzr0ksPN1reZwdMCixOF1Xbz
5VPUTATbY4VQ+jVyyjlQbttCytvQhPPcVj+kG0u+EHkxY9lYibja8u38DL8+HhtV
HH7FN7hB3378e8xQB9kXrAsnrNEVEnv6sgzg/49/2jPPahUUXAcs8zigNxOcCYcj
sibkRTX8cG0yisfJOSw6WLR+xpQbBmJ9D6rSpsB7qZQ5/dVXRSPwZZmn+5o/vsji
63lJoxyhJO0lLRiRgCn7aXsaVc1t/6nvIR++/bW1XtBzqO8JFhZUcEuqg2rSNmiL
p7JG2s58/S3z/BydimJ+tJfZTbGsEVRrG3IB5foIUPCRtH4LHvT78hIgvnmAk35h
KUcMljVGw94N6RVkgKLx33kf87EA85OBMPH41RykT7/UV5ZIDMNCsxD0BHJxkWbX
P5B8G82/JZCgo2RglR0ZiNUjxrnQJ5nz1A0ZkHKvDE35NotaA3C1bO/YmEsSXzn7
cpm43RhTlvR01ppXpFVLy+lFme4WRb0JZ9uva4nP4BMCK0qvIJWj0+sn3wOK4iDr
bblqUDmYwtnz4sG/gbm/1463mAKaPn//9bUXngMwlnD7Jetx29hRK/bmefle9NTd
WgJ2C+0oQyXjPwiwH59iu5+pmUxq6YdLNnOSVKTYLGO4SKZBJ9FMQ1UNv6ExgiRn
RSxQmQ5qk7a6kawabKmjRk9fP06uS43WE0nksMHyr43DSjfy7p6+lQBy1MMAAiTT
thIlINld63JmKDkQJyZLU0jxDgGUMBikLI9sfIdaWWOcatMkC1rQ4Mp6qV4TnCfp
zJcQrsJUs81wAWE6FEoeyXW4RmxgGsZYzvFEVs894vaV/dinZhU5xeszMm4yhbYw
g/28gTwpCDjw+UQBaMp9/IO0oiENulcnhe2f6IBcXbJSfHW5YWisThuHlNtfkW/H
XJQLhJHrwC3l53TredQntKHOhb/P3s3RcpDWaGFbJ75+wm5qCCP/+vR/F3IZMkjb
sJtap83OiDlRT73aUD322fGuQrYidX8Ah2TgH2XBvL2tz2goZ02PQXNUBX9+g609
vDELA04J7HGHYPqdv4hx2eyCZEBEOwcKd2SUDhQUyLkeEk15b2vk9u4v+8WmeXAe
nyH7QoPvpHG1DYCNu92WoTp2wY/+tLzc6xVCE7e3W391FXo9j3sovEY+v6BjBn2O
TKQf615Y/Vdol7UnEibKrGln+JI6u+3jCfKM09EuDXeVGTN3eI410JD5jj/NUTyi
3d+wCzt/QRjsmiAxl5dZxpdTR5ywWcaSYUYmRkQPl5LAIl1Y6cltIF2MYi6lcBsJ
yykkc0qJuX8Yz/SMtjnQSc80Gkuk96rA8NQ8nIEZzQomZ8xMoXMWOc+hKzVEoa1Q
qDihIS1ltnSW17xptCiEvgMrRiQrMnJQrpETRjQtP75Ly+s4IqtRNjULOqMS+RhC
MPG44Ho+ZUHtfldkTn99xBeUxyeBS+WBbDOJ7Gb69HT7V1J4uMj2EbeZ6R2qzZmR
ADgXYgii3czcLQFJw6j+JBf4YCDrcBFu4iXT2nNsZPUCRhw85CaW8fseuMq4qj5N
bbhhuFQl+MsMiZeDDSVo1ENTSdr4LJ9QVyTiwrQNy7g8BBFacfSbDnq2qPVjghGO
3KrgaC0nXe7WdofaLNhLo5gyxiwgbL5x1LUPm9yB2zQkrb0SsW1LMnzlwEkS0vW3
nS0BDmEBKqftK7z562b5TojcU5V5g2IR7qucen10BxHNPONbuOalVePwsT8VLw1b
CIezFXgJFI6+bgQw7VD+uYTWOoskzi5vt07EUVs0o6sgjqX6ufU+dKi6YgvK1UhU
lnVe+53EEFs6WaPmRADYg7cZCQgN6V+Tmr7l2SIa3cygdT3X68czkIiYHsAw18eF
UMVqSo6nX8bjjCFY9e+HSo1oiuR3q38Z3dbtcm6y1V475BKJOCG6gPvFhKnvA234
hd0R1eVutaJ5fmaJfiZQXhpXKWBHlgiuaEEioR91XQRhn53CHF1S3ju5cDdQ2bn6
oK1IfrgNXqrdwN/SUB3rhccwn4de0cOAgc7qSiBj7H11My4xXZaJ4c4pd9Or7oeh
Ace6jVmkvX5U8BHIaJONQ2Fbqj5/s+u+I9XMm4tfM4A2vpMctcfCOhrQ8axWHg5d
RNujWgbj/7PQpeT8yXZZZJxzgTomCd71Q/ZGMvwFWfPqM/KVE7cLcYr/9Ctfl90/
mVlM3hBV/Cb1M0ri0Fi6QIeqsJzQ/Xfiwg3B0bUtnkDWmVZw8G07/uW29Fb63KOF
esxy71CAkD5aR4oUr4SK5ZvkVOvC8KdYY2Oq+wHmh9/b4ztL5owfD8cdLT8JdSZm
aPG0r+m5qFZtvRqtQJja7EGkxU4CsWY2DLKq7elBGulIrbn/O3sB7zKyDx6gmdZm
kCfi55FlXH5T4smoIT4Zca0Pg84RftF58/xCRPVneShmCkWLe1WICclbm5RMt4Lv
ZxQFzwDFfmYztv/uQfmGVMzo/vWB13fK+Z7+0E1BSrsdiQPrqSLRKPiaVbVksjRW
eXTRMTIS5WKJBWZyr/fipza+N4bywdBzdk6gXBsbWc1VzZ9FOXzfoGepchod9lTI
LHXEWneiEVpJ49D8in8lqyl44neRI56B3xeISMJDlQ0Y9C26OQL/YUX/4ppYBmFY
2kae9654+cHI4qPOGMrXK5jTDOG6r2A1WSar3MZtUu9+uYeozMZNP6N2P6G8aUkt
orJEH9fqix1cL7uRQ/ikFXbGiU4+KMFa4MX4sPrJfVqZRi3k6q/rQk4byfaCGXcP
gvTFcjxjYHeA5mRdK8jrpQRRevsR1RoBiHfvzrsFQrRBls9pVwm1nwpQwLS5t4MD
5lOtQ1mU/4gYQqokHdnEiVeUli5zj+fmxAniK7IgznAYDb4pdhzSiKI7SVZNhxq8
MAAqNu0oeA7a4Fsbd4cEomQev3Mhu1O+wOQl2xPdi4YvTDFZM8c+Zi/ErSD858au
DOUPkT39C1vSQB15VBi8+jPwv6dSwlqsHbYPjqend8CIQ+M8cB7F2J1VjND3ckrT
x+/AKd1/GwZtpARpmCfk7N1yRHC3QaZFy4tIGlEaqjZlmaC5+w5YgzgCEzalHWW0
zD3ItypHJcz4CbQ7203CZVZsBkHUHbnw2/8HeaSdYfQ12zUKXMTl767boJbaKxYd
GWkv3pRtrGOkrYrR4sG95XocsUziRSTzIUE/z0cO6VVNIBJeKZKJWayKg1jAaFuG
lWgciXshH+RX5Vy+x9OL9SV9h7NbNIZDLbm93Noze+D47m0p2Tpg3pPLj+P8IaUE
zb1eKDD4Htk3bGDuw7es2w+D37P//YpTTOyIOhqoVrV4J0yGjq/yEIqUmvkAoOCj
rbD/f9VjOV20BO79WmzMs0gD7aP8NgsA0BoOYlC95ofTnC1dMG7Nmse72k5w0q4p
bYbe15V/8F4bK2IdteajU3yOz3/64/+Leu7PcoE7VBHj32Tk/gjGlfQWvCmDOsxw
vNz9jArr2zyXge/Pgut+jfm+vFd4NwzOI4gtyuwseLvbdEc7y5TYQGBeg+6Cz/9t
y20+SETA/X7LZkR7PSgup+hf35OSad1DoJ623aCyzIO5ByUCIJ3LmHUH9cg5R15a
NsuanGM0bF/TXGXxfqmT2br/L4GpnXaGR/KVtlAjvoYta0sqr4rkgSnsfWhP/MOI
JBfiZr169v5i+ag3TfBhRqod7RIO9Ss6HdQZ10E/Da00mnq01B+IJXrf8O+PiVBz
4IVh/ErpDevP5RNQkCCcUFXw1F87O6bxI3wAEotEJooYE3AxWLObo9i4V1igLNvD
tPKYtTKeFP4IVzMBi6sdx32tURBSKTge97AnqBPHG7OD+eGV9nwe1SOkOLLJk7ED
z1IzQnhfig7cU6724Hp0kOvWbYtzWUwBom9j5zafbVJZKDDy2TlZ/MM4Z6rJmg4g
1e0CEupZ75MXTint5e+z9B0b7wZhq9O34Q6r5BmwcNn+VqjJOQmGliFVf5VyNF56
bfhs7IZNEvDXD27Olg+CGemTxa/4AwS1++90WAA4+eCkloCrPbIsCQC4mhoNBIU3
wRrGBS9b+/B6IrFt/v22RCw0s6Z2k6cJW+NilnqkQDKVfb2D8bZX5YClL7kjW/J9
yBX3JczLm/Snim3vhIJiQVplBBVmRCayFRPV4HBY1OUaVIgdskLMGIzlm9Faxrua
J6SdZDbxP1DhsXNG8oGy6EX3jfHZbrhq23qGF/tT6dDtzOPzuH6lI8hUa+ltLkPa
vFujlAuvG/Q8/GSQxo5iBVK53L9skop+IvRsEDAcybffoo5uF8uTHodr9vtA1Oac
fh6tpYtARqWxKCjbMGA5KhzyJ1xPaKYQgTUyFoetfrDbzgZl/gotiBRsLIzktxPp
uLvM02rca4HD7EVPBjIhGmY1s8YWH7YHBPW3L6/XvlpML1ZHXzrbvV2XOe3Y4ncz
/WUwdMkPIBUFaqYDW6lpAGaCTJZPIWq12nqZC0LA0IHfmQoYPyooxNhTWM8X0hLS
ZjkKYrGY9q12R7Il9PlktAjjYcU/G7hL13lx27q84khrMURyqp1UjMCJ/YuN6kT8
XxFPV2qFdeOyS74N1MUDN/28U43jUJzvC3xT6Nd5CVzsKbXdO7a3niLvskxEwR3v
jcf4wiHmVVr1oE7PqvslzYLPcq777AERFE4WSSjb7B3benEAls51H/JA42fHt929
rHEWqi1Zn0cMXvrDS4wQxuTuokR4kAQQPRX4/qpM00KpzuLOY9Le1KEZIkk9XVSF
WKwxLGDuYjgs0yPYyFt7LPqWzjvx/T+CSg1Lt9SD6GGgYpcswNQN/+0QCPVOIqPC
D9nFcNh0t64sNP+9W1YoplT/UmMWrp6URVqg/6f3GVULYNeiaKnx4yWKTEhMM0ep
Pggrr2ziDcgIkZCu8lRNJbo517P5QizFT7NUGVcu5gAE3QuHSiF25n9WWv7vtGlL
7mIoz7Wn9YlCdu0pbk9qXaEqlzE2i8c0GXE+TBimzQoeZcrZQz54TRtFvANbJekO
q+/uUkMSEINKc2b1m4dGI5ZjR3wnWVDVcH+FddOQM/IILx99d8yNHMJvhKRdSre6
LDBO62Wbx42/kC94wmHGCGg/6TYjd+NXvVOGYne1/SJCIQ0Kuzq7P51ekcy3ImBi
CipsLtrWtW7oIlzEoiQBlUOQv/OKTwrb2nVZ+LdAjt2QT9+BUI0b44M4bFHWMjKb
QRtJP9Sh/FcslQ+m9Oj2uYxdHT78zj7hO+7RRRgX7xpNd031ZX9F8nl4turDE8qI
+VuSKHmsS4+TKsPUnsn4jaZavuYXyQrsGJFIcpRUgsNYB3BXz1Hf3JPR2ItDORcd
inTFccagkMQKNYOM3SEkZvGfLHmqJk2Q7GyToEe668Fb11ClFjsZ0INRp6YaoMi+
KfBy3YoJt7eemRi/7dhyMbYaJhV5YAS5bVWwHAuJxDrToaNpgFyVCrx4zOdfn40X
FUYYwHq7GA79Vihceqi1hKeQW2+vE4GfmqMHzfh6xG316e2ulYeb9casujvxSIKZ
BcK0AhSkxwBMO9F5yggsCvcyRRa5er+ro5hfTqQv8StYD3EVlzf2BUWBnso0apWn
mHzimi5JrAd4K3AOV18Cot8Blg1VaWhc52NAjPM2BqIUke/nrA2eRFiIm/idPa9J
XPP5GcdBXptPUQFbVq9yavXiKYaqnIQHWXlhihENR/WEloCNiOtPn4FTlm0qQA+m
W3gS6jiBbCQZJV0nGQy1jwSUKoQHQJwMTYcc3LMtdbBOHvro7iunaHzL4L7ipQnH
d3E70Qfa8fHzI08l4ghImCtkgt1Wq349za9BqRw/7ZmmdRvRi7y2MRMYiUmQrYFD
nqstlLGHtOnmnIMN4/b+VFZ8gEugbJTeqtqPJG2K5tNMe4YCJI6h8RoeXBU/sJPe
2St3cpLp2vV9qFQ0Zz97uM8Cxty8DCzqb2U2R87yYuDV1WvvwXzkvlZk0JPifoBN
Pg3ww76u2qIfhzhTx8ri2R2FoOO+DvBl3W/OjRgVPkAtTIDoRs9/YXu/5sBJALIq
sroD9SOVSEvZZmUAcnZNBr6tTBZC4Mu/ykZ++WTLOt+G6gXyEAtW2h9Qc589pww4
wDGnMaSw9svd3lDWMGZ0YocSrW9GFb6jgdwaKPSJNEk9RI77M4gKSB1S9SU+8Eku
lHWwn+svhsXp+e3jZHpAQA8Cg7PR3RVOXZhqQqLEW8hIUity9BzDt0F+35cZ/peX
TDX4pZCDUXgOIy2kIbo2SM0kKd+qOlSebkL12uaKMLTrne/J5oxsSfYS1MUdrY6D
DEqpnp/hrCvmuLOSOujVb74wFU5PwmIqLHC0DLIdf9pcbzde7YQcmEAuYZxl6aZT
y/kVZoNIpArDV1rcdktvNpa+aVuQpGJeR9BtK3VB89Q1Lk3tSLUXcbgDbN2iv826
CuH3om5I253ajYZxpd6K/wjqEITMu9GFcZwwo862D5bRbTNo+FXBRWw9H0FcTD9g
F6yzyRgtxC0LhmxteH7ltnt6qqApme4KRAGHp4NXt6PCyxfVWCZZHq0ZJB3dgUYO
ViIZe9Aqhhf3jZntwidIaW38XYRJjhZ+X3XTOilWejru5lYRE0qjZ3Fq+GCxLVr+
nKobgcH/wSCLcw7ncRb5fKOqkAbZtPnIJc5tKCcemyiRpOT1ybfk9BijIuuhAxNT
mtWES57614zshqtb2D1b9TWob/H0yPKblAp+sr5ttFaDbqNVQY/gzaSNewixnusE
KsgigRH8lLWVST3U5wM1k/eHHMnFMqNdgy1o3M2j9dP9xNLR6I5Mgm5s0fMZrOvu
TNuISlNJzsTLE/2/ApFmDtaLbwf7Osv2ZkxzCgBcvxO0+gMhA9/nQ7IAmXQbGHOm
ouSlS4ccYHiAmqcxEemFsC7YY0+Hdni3lIavbAckorJjgDryQ666An6XeyGkBrGi
sc+85joPYqSpK2hm2OKykFrH6WTEsHNSDOdNLBeXfcohFQmD0JMEMmwTd7jPCahI
IrbLrpbqGGCNjgn6ZFdBUmhn4XNUAM/47GstNJXH7h4id96vOdV0zZuF7VifEVY1
6P9TMy3oNGVyZ4y4dMu5DT6TrqIicBU5XS2wnWo1khHi4wT2lsQYvDJ3eiGEyKkd
Bw3OWD7vxhBaSqluM+vwItuGZq85ahkspqfi6hTMuDLq6CFAxpQqZPHOlsX6U9xC
QC9QImQbW1PaShOvy3aSUd3qq5XfdKAbJ/V9iiWrItlrL47dfB6oGyj8b84S+Xuv
ddK7ZcFVYG8HfJ04Lxu/YwWOx1FZVL2PH6rIjbviz8e2pIKOBYFjOZd4L4R98D5k
ufgVQeTGkaJQCNtYQtYvBlyBsGUNIaeEH1jPJYxED1Y0yQHjgu1FrJjQwrbpT1lX
Pb2MmVnU8Ct3WcdbK9Ojb4HIKgMvO+gNrQmtspg8Eo/sQYMb6N2x/8fHxOPqCL8l
PlGmeoFhqDV2WHMUPu44Kzl0kjWN0l6v66OkDTPBdNX8LgOrAYAGLluRYLgXzOMG
2xhlBGTbRVkpjstCALovB1pAMEh8JmnOkig5+Yegfdp/Mj7Zyq4c1VKty70nZP60
aZ+k9ScTIh7ftpkiJzC7un+WN3b9e+QU3mjz37Lli+Ct1EU6grFw+0y29bgFSd2n
XUL5KD78ytC5/Mb/LC5MD2wErxiFm7uvCFw1JXRXFyZEBX0vrGGxK5lytdNfjoBY
gGbzlsndF7pLdiPUADwRZ1I1xGM9jlEDwR1Nynb3lNs15jNES3nHtqLOmK3exyO3
G8hLEwUjVIPI/m8Eb01kASEjVG9eCgsrk9En6qu9LEm+cUNri2JjIW16k94rl7Vz
TMsL0WNF1bDqFoFyqutO/0ub6g3R0KH5goAqAaIFYvQ+5UdBW+TI9FQND+kRT7x+
w2qG2cltDk9EGO4ehGrh2/6o5OnGHFOe1kezFvYZ/M/YFhWnjB+axec2C/+gZj1J
NkXhI1kJa9C3NiV+IbHbQLkcWns3DBYtGIRnEAQYOY/iBMDXP5fdMnOao7czyW3+
+t8UakjU0yR3IZf9HSvy2R/3+YyIwq7QNibq4+k5ogynM0M8Q/y8qqifkTwptEDY
zDGUYneDBDyJMjnBDHerD9l541A/YoiAvlWSPzeV8vTkXiD5VicFMNIr2/jRiCbx
1SZB5h0i38XHqUCmx6HAmSfedAzol/yrn68LuaeKC0PMIBbG7i+8/apDqSfZq51d
bsKZwfLwwWsXjxP8oUS911eun/Q0EQbQOiL/TQhiABOGDwoEmHAXbPxMZQLB3JIH
1uBsmIafpvcQQoH31Yja5kqAtDk0hny3fk6otdEKz7F4LAff3HEGybqC6zQ1LqYw
EETTohsmpbRc/hIv1Tmlq4smMXkwWlHRK6cT02VGXTzafdKBVjsGrYueO/NPgCBP
Wsc3f38cTX2Ihe0HW+y7+GpWUT3AavjQODqAQJkgGnVpr2Dvk8XlVGePH2eO1cMy
T2CnmWcGjHhO6EMV5L1mYrBKCtuLR+tOyonTX1xX1OpmW4f7URlnKS1rwNlNVHAS
OZyzEqr3cB94TlZp6AzerM4o10ixmC+sdVWjdY2CfIwoWpt2dhxrJFnUhLUd8OnE
xEDyqrIHnQW/y+MBWjlNbKunWaxFDdBIjNU7/EMt+KSji5jaB7avZQXXC7O7cPBL
EVQTcLUzTfWLztH9g3MYHi3dPXolmT729Zv9+VZqGuIlTNLQmToXJitFG1P1DSFs
kfRJYH2suTBZWX35t3RSjk5WazLHXlE9YLZ61avGXP4nCMqZ85PI0hmPG3wx0tSb
OUTJpXJfLdB1ZuMXeiHh937InSEJk0LepHSbZ2osCPIjCGQsj/B9ExPOn2XwpyZU
5FbHEFUpgaNV9n/xUARJ6NKNtdoNsKNAC2Qmx/fOY2Gqj4S61kOhTpLe5qCJLbdY
Dmv0UUTtoyp17ALOeIeo+xQrtBYQaoMwzg1LdTitb98rd8gBHimLDxKkB2IbZ4ZE
OaWHO6EjMf7HnEuMRwDF60m3uCbx0PfnzBvAAB1xozfKpc6cG6UXk/YOVK7NUb3x
RPqd73SOKsnndTyci2DFCuQfcSWww/U+JtU+Wqz54Gb/Ln3x3kEeoSU9fMNdvwKg
NICYntq0DALyiwrcu6TOYT5RhrSMLR6GZSnmbWBfd21qWg1UtHjUWNS4WHhyFsAw
q8QT8szFMZrPLjAf7BNMLDMI9/uwhW+ZhMFxQUhr0ofvSb+4DUF4YrMwcPo4YxCz
chjlQboKyYWKVflimD0i0rvUSCHCvx1sRskU/jo+R/39Jp5eRlLy74fgmGwU/y5+
btC71YP6jC7ZKIv0haBaYd9AoTZLZl9ReVeu6KEqVS7AMIVZoOe201JCBqLfTogY
V1XFZU7C8IvnDHdNt+VHDZutKwBFpNw2rWi9IhoxCvDkRP+AHwFdCeJTzMxPfZvb
XdgfFUi41rYguf2xkY7Ob5VRnDhwUid1Dayi6IYHiI3CEalr5ExcCuj2R1ZAgPiO
7QWUiRaS2XyfiduqMqmUcYruY+2BdS0IlnLWBiW6d3KLOxGziRa5c9Y58oiIxt6P
+V36ScZSEAlE6G+Iof1dbqP9wBRWKf0dxyBKRfK+VU2k4M8w1QSeNb4MebfeNCFo
Br5aMi83MEu++xo4P+Z0xVUXm46Ojl9IRIAYb1wIQXxy+WyEYMdYTm8FwvBU2Ne5
W2IxkAdNO4ijXvFlM2HHbdl80E0it+gz/7Qy1IULYmxNlLNRCE1QHAVkwOcohbg2
w1aGxrHYB28VziWGocQXoPusXE2ES3+IJluVRChTHMVjdThm6YBwMgCm3o/0VvBp
BuSyr30ZaxKtRjB4ZFte+2YeY+dTCSYEbzNLxSElamfxhJ/QN3dhLSMPi85jCgf6
ICOr8BJMom5zAEHzSfepUFc2MPsVYK2fgL1TWSFEK0ZmGFuUKpA1Njk/tqUQU9YJ
d8U6Xmb3QeKCIgWAvOTTtKdJBDI9z6Ee56pnupeGHSR8K+JoUQmrwy6tJ7fmdL/d
6zROOSzy4SEO9Gc4/QLaDgIbDNDoaeJcXDnzjM5njYkgoeyNMx5jN/u6YwdAUyJh
ZALdNfkqc16sZe4289UB40/kU1TydpNHAyNmVOW5ER+CaV5MkDovXARVqH5saNqx
sMsDf6IqaQpQaMvpXgmSuSM3AdftwoMzWOR/E8MRMFss2tc+vtxHMk6p7Pr2fH6A
U2DeX8NhjskwtS4D9HAjPD77zw2SIr4fnuebn8qLwNP4wbS7TZAYPoWqSBU0BMjg
z/kjReYSYpQua2hungPMnMAvlPnBxq20bHdU/jk4iXCGQYu4uC3TznwYJFK6Ng+S
Z2ymBuR5cwoErarWY2iAG3AiqaPUqxWvbzn65qTzi5TlZ/glt+aap5VLhS+7pIRI
/y+usXIS0y1HrpN7gD7sLIFzVc10cB3oOYc0dvp2WKvF2EqWPybqCRXWL/XrWk4O
K4aaWb3SOx9870+6dyIeK07o6hEv09vs6k/RrTw4wsQ4mQyrpqIt/1SpEXrFjNkc
RsKZVv8bLuyo8hPulbK/H9kClcD9WD7PrXmJDeUGQdMPQVbucCmc/R8IZG/6BFn7
2BbIWh9Z5yYMycWHBtPPbaPOtzmAwjxW968SSPoQLdN6tC8Ckag7gwiAzJI+n9pN
PsdhGKrRE1DvO0ZkjU11TtOyDc4t2KjhMD0oiVGCUW88x7ewTmxcGyju1mBIq6H3
ldmKEWhMWgD5rMK/djIBjwuZiMBwc3QppiQERlnMoSjyI4/J11SurKy2Jq0vDrxT
ZHZZict78OVrPGBVvtee7SK58UsOcQNoo0qiW8Qka+AJphwcNh4EBW71hgv2TRUO
3kpZxrSc6JHVZYom7M7SpZeglUV6eqBQky/26jVNseswkzW/7VhhlSlQZjPgI/AV
ObtsBYMuv+aLZOek5934BOwWdufgjNw43gnS86WN8zB+KXy9STC1T4lqObqDraig
8eluHIVML9m6YnueQr7WHroluQ8srUAdFnZHOqsyrITAqZddvA4369aqnLXfQ7/k
HPfn3oduz+jBn80v9mLdf9Za08WYNLLfeeGM2ebge4ZeCMyMBKEYwdBoDWXyNEUA
t/zOoJN7fHgb+VcIgdYBgBJTIO2JsY/axXtLj53sE27G3rAIx0+qw6eGw/gSc4IE
YRfXjIkIz80GFlyOH5UQ3Yairk0GYA/ulwcugTKTHeUcvRqWduOST4U3/P7cyrib
OFM/hbl0SMdSii84g8vUAKtvKWgsDxmQNpy//ZSh8zwag7+p6HfNCPFoLrEn+45u
rCGGwYTUW5TySmld5Xq+X1yZOHlZiK+5vmdhplypmJX3Gfl++75+ONrfPXHeQj/D
6Foibt3d6ytjaTZ8Pv9oUQJmd8QvYiWYDwJWWQd7u6k0Yn1x6MVLctuzz6JXcrJK
OQyeRjiRXXNEoD0Rsr7Y0P5+/MR9Q/pR5sM9p/byiAjfnxJE9prKOXIGEPvWV4tV
5uLaHJQ42FzAC2qk8bipPvZJvc4HDJRbCuf1dht7q6FWx3zOHiZXw8XPfxkxWlxO
P+Lt0Dg1NWNGYNjBjzphDlV8OiE4eIDE8EUGMMRGyjn7Ht5K1zGqAFB0JW25QR4V
O82rko4TuGIb/j6HvRy0mGkxv9BDL7pnAr8CE+ykYZTSk32/RUUBp0NDJIHkV/E0
GFkC0+fjJQrbOaITWDxdS7N5miOvjYP0zlkO1Ynl0eN2MkqahiZ3oK521Ad2KsOD
ELJn/xBSkcyM/Quubdfe8U779tXO3DWVZLHG5/5bHt6hIJOneR/iUQ0rVwunVtdr
o9jvr9ArOKzcakGHakV+O6jIH5yPYNIRmm3pOPOWZIsyLmS0W3I/zxgp1WoGIui/
kW47AH9hliG/3kClvt7ce3NYeumgbX7DaEI/jf5M19m0d4IqGn1MfcHN82I6ZAWZ
+ORJJpzZ+vJiOJt8wXpKiSKWHfptvPZISjcug6o5FGd1eyyVgkgiLggx/xAiheeg
5UKnhoTNOl+KtUxhqpixVANLCaPELiDTseokBVIOyRVQ28YbEVNqoY33wk8uVDUe
20g+NKT4nMM3oY3TFpYVAGq7LpVF8gpDol/sVzoNrhMFGZVHbcHexSQYLXB8YaQR
lJK4oAs9lY7UVbm7D6JdsidvnPGao8pHuqNjFlVaHyNIJwIWAAjYUmExVqiew/n3
TQcm8zLVaIMAxGhNCR3P22dc+wxU3PBtXUtqizr7Fkn4NNOXEhpqXRXVt9VKi/5X
KFRjrkRu2YeTsftY0ydtbp+wxlWtSscGPfA7QBOR3ZGd39vPC4vnNfuV7G9FuefH
pLi6LCQNab3B+pCMzI2zaa1Y+6PKKGRUZ8gSCXaVAL00IhKayc+5moRVi+fvt91d
Ad/NX2f3fEwTdINfW0phKXk+62v+Nqrl5NoZcyIHmbrrn0xTwuLSoep/jUPGbp1T
eSio0icd5L0+eXxAl85ZvD4dP6Tycq9y+4eLTcLAvSpb9ryUpIwrUBm6yUAuHUDq
wIiwLNlalr79H3JzXmGDMirf4F41Tvo7SB8q0aDLzH5XICfQWmcJMQzOon+BMRaG
kBKUvkFg7n0XBgowoV1FMnWwCrW05zoLMQJjod1QnAYrsPmPBNYl6gI1KSuTrF0p
zoJ1q3l5jlx/m/i9Wf8j9l6y6f1BQrbxQXmhAXARthWZPkrGx1f9/Nwyn2oYppQy
QVDGVbeqJsDE0r5WKWYC4Cnw5AGu1c+I9ZliOj7vLac4lfGVaY1q21GnCXNlJj/f
ErA8h6eUdmLbdlCZkJiihWvhjmi3KLPRckbulWPVgpc6qrF7iEKXsyRDKRoLPJyG
qbcFM3/iJLfjijZ+bazcUxBcGqgy58nQ+6ONr9JkivsXeqNyOla4yjVoxXz7BmCe
FI9HxCLYGdfE4Zq/fbyqUQiB9B6PU0MpsYlyXGpKmfP+1MAZ+Ok69cg4IV9JJp4F
wLEPm4VMGRiappkjEYfK/9Cq9dv1JlfjIARgOwiFcNXeM8AQr6DuCLByd/OkHavj
42tjTg25N9Rx10aNDNmRm2aJZ4xAIvcmVKbKPfDyGk/fTyuSSBu4MKqNvkarzkRu
lgodW4fhFwHgEZrdvS/vRuXqUVsBov2wbohy1IIehzeznX3z/rL0hQOdY7/yXB8J
ycNjeOP62MdMyixt3kze3FF3lTICliKRjUXqJHdwD09qLmA/TqulReJFIeJAG3mq
FC8hHwBAHr9LHc6oKQJQdAOYMLnMk75KduhFYj+kRFzuT2xLAiPu4R44PguFL9oH
l48ZaxOJ3nhD1GRfcQ62UQ+jcdAsEfXO+V4pdBKrLGae8CExAHb8WB3PB5oM4aGl
l9MKwBrjoRJsa6vYbNx13+NZg0qJviWa3Ds/D9YUzCupRrQ2502x4ZZNv9YByXuc
rLq4cdbG0bkbMlC4Kzm70mL12gx0ySO+Y7BeES972FsyZJWGNjmYpSCuHfg01vIv
Nt1/6hz7LV4q1+hl3mWe7qL8YjmzHSbf0C3f5Ry7wg8e4wIMNJ0WrhBbhbSK2ceX
JFZbOjWXjtk9XZ9goMRrOs+Jujdv5G6T59eaYvztnSns3v1XS2BGHubwGXTnuizN
/ZAJk8I5PNYREWA3ieYVwxuWAPJAEatIwzaQWolAZ6RGD9V2p6zhH7S32VkNKW0m
jm39N8TzXeG4PLQg9fxeEkwh3+SElX8J9HTmA+DlmxRggjJ+BLGHT+nhXClMhEre
89BcLie1mQtMDJwLFvbsR33qVjgdITgD6XLLeQD7Ti8CTr1MpkTpivaoxnVsuVbt
2F1c5PMOHts4I8MVF3eNHjT6j2VGO890ksXo+5VLIEDKYHYlPgevcE1+NRRQkJZQ
JaZ3bK0z4u5X3OBDi9JDNCW0qzDFrKLyF0iYZsrS9tUbrrGXB95TdLwx33+p3q1E
G3keiChW0KSX8Jd8XJKkKurGFNBUgEB7B0YBkQsz6VBNBZt98RS/USgoPBDEAbZT
Y9iCC4UQQyYbeN8dPdubXuG2X52i2lrlMnbl+toF4pTvG+1HW1PeLHzEWBN4dg3s
PzI1T6tE1Otr9FGDmqQy/3CDbmSV8ipRPysDvz0HO36r/t/8R0ZJ+fGCpUwG281Z
WImMBBvCMWFyWY6CypPZx00r7US90/G/TD4Tv9SUwalMn4dPPFYO4n5a+586m7lW
oU3Fbvjdg5TYJ89wzZ0uJg+2YKsuu+WzSBFJjiDTh54qtLz83RpPuA3aiR4coWkl
UhS+amOykSFqz1zLg/UzBF5BhMKb3+o/NHSRHMKVG2UOfgohiSsyUd1nPQ+51Lcs
W10YN3RJGZFlT8MB+5PsfE1KAKYWXSRvE4h29L8seFo4Th4jlrJZIr2fSlKb+da/
KOW+d0Dcrvx8IaUDo6LwH/FsqfuYQEpR4CbLj80JLTmky2diFfjNz6EjH7bwGcQw
xgGNa2AfOozYqON8LapVMNwEpxk4NsvzQb816s7ntMA2NpeetFk0M9LHKNgMMi3f
1Ivylp4x1DNczctLzkX1Gy0au0gqslVMSp6P+YVTejknOcOFYmUj3sIkQS2kVzbz
NZ4+mQfreJvCMeE/WkjPoYJpGNduaq4wDsaMgIGWJ4MpM6bFzZkenAckGzLG2GVt
Bs7WeLLYF/e7BE1MxD5E6xa4OfIX5FCt8nBO+7B7cXGJSsv/BLwejEAqaSV8X6Qy
CW5fiiANreUjNgYtgxEHgqpwEcLhBcYIH2KC1diANQ9m8nWXSaPhTKgQdkeLEC8t
7SpoTREOMLQBjKTNDD4qDuLs/LFD5cB/6WPnuiG29jN4DcYryYiaZuAi0nUZmyyS
w0/ZxlQChRkYXK/z9+VMHqWC1BhxIHbfnABlDuhzuSXyCvDjw5/gdfHz1f14V6dZ
+MtN2QJ8f7s8YLSWtQmxKxNdGWonEBn+SV+Cgn5i9EcZ6O59IN/qbY1uxvZDnaSY
0pelLqadnPI5qbCN3FUtTKlauExPXdq6/iUuqA3Th8phQzidbcXdd8ks6P4aLkzf
g2p9IjXHJhECyfNqXOXB2ANkz5LuBQrPUEz8XOXezhlnbx+hc0c8YOBMbvo/Ng+1
q8CrOd/vta/n9mkRF0JmEjQsKtWCJeYJByvhP+lxsH0ebVBHYB5s5UUe/PwGCbdl
AU4lHxB+Orh1zYG2I8LCXbD5lKzZX/fSYqrSBUMyZYKew+mVrfMrOyAwdaGQMSxz
yZgQ9aFMcNX4qykz11rAybAh9MUsKH8pXobE00kxoQ7nhQjxwoFNsIP+qvKoyFm1
n5LQRvBbVBhWTp2B8E8ZCn3r0M8QNsPsXccnV3fDUxmVivlgRqXMR1175mnzPvP9
2EjSLUl+ZAugYQAFrP2BEBVRz7qZda0FzaI9f2eyzwvTYuYdCLm4TM06It/j/ni1
GviJ1iUyezRrh3c4myNgD3vsHMj+PecDL4fBjoj5NeohAVyRnMd/Y4fnX75vINgb
4/rmxQRWerRRW+t9ayQppJ0qxo1CfEp2VzWsu462WiQvJ01eF0cqZR6Ff+MAmnTt
xiuLrbVa7i3bW5PKrxV4VZC00BknVKKcg803wUabljDRGdYiZYHfQhYuBAnCi5cl
bonQTvqhhg94kNosscns0ER60gMVVxrlQyvr3csOX2eNBsDHI/vZoOujl4ygwYYT
owQ+tXAsmQyJSF8+op2IWGc0ktnUIxH2bSK0aqwdVifN20xUaX263PI33u768Djl
SHSjzDVkVHKgLKmuz2LBUAMVZyOk+TrwHSkzLeWTLQMtwKZJTC7GdsazKlb9X8Gy
IvC6tYDG4OwRQ4Lf0z+IhIolnYRrey5hH9ZugZ3+dm0sVJiLTQMmsI8qHEAcdfDz
cGnUYBK6/oEX33ig83DeEK7FhRdz3fRpHfLr51gMIQtAvdnZNm5CMdJ3kAdg76NX
hIXvxsVknQ8qp6CnchU+/ujBajr8fK19ZcPADMoEZsV04IBclGsSQOyvYapsJEj8
v5jjXaEdZPG/IC4M6BeizAbwmSJL1LHqwmIqgGKizMHc9p1mm1dMl+Mr3GJKhKO9
/BHecwPIqaRiFgZCAHWy2pMb9HEDC2hKl94nreDM0PdzFvPJLmZBxiw0xLY2euMX
RGUlL3t90Ktq/Ox6nQ5D5/x2krWjnIorMANXVUcmZ3piM+uZL2Xv1UeZSEzfnqeA
S1+K6uSb7Wl0laMSi7+bJqhgLLbSMzkyR0EhLg9c2arPtiiv0jIkpc1oewuZzqd9
+hYvXfxqehF1nOzp4G1i/g9A2po/RknCONKdCLg7cxln8+7EtliWdZ8iTcoq7UnW
3SEsNTZY0FCX6NivCNpvazd4oadis4zO6tB4dtYj8nq/ks395B/SU9Rf6mdC8ir3
D07MHwzNLgyGWcQfXlgHZ0L+ZoDdhP9cpUr7fdUdjcDhPvt6ie3OaFrKhdGMULfr
8Asku0Tl7SGtekLTyQE1hPJGmwMpqHgHLw3loWIH1OU3mAsEzGqzPOc5PQcKtI/A
ejjLv+0gvsfFgbznKAiamnoX7VAGYQFVJ9hohLZ9EaHqsTWDkEHmvVorR7nKzfjI
igih8gynAd36dYvCFmwKnc6rVGpxmjie+epN6XFzRrH/+F5fGXXJlEVZkxWdmUd3
Kbw5ltKrldlqUbKGygxskJj7MkMgcWDffbxahMaGQLlaiIiLCD4Q4i0wXKLbA9WC
oYyK2cZ36sDNTp9QEn7ESY5IAd4HsWTOQoMWU6nye113N4ZubFmKGjrSwdNEQyH5
RUOYWigYDgV99SzkQ2c7Sujr8gbO9FY4zIGzFHG1Jksf2/+sAVYJlwM/8aOizcV9
pWAF411r55b3erFikv1wSC3ZgMft89MaeG/dz2YMdETkeehwJVsyZxU8jx3zuheF
GeTJkvmCnGTmnmLwyuGmlmRyMKPqrTQ71l+S9qQ8E3lyQMPMXfFUJ6yMyGw6Emyl
jFpJnaMQX0smq5i6OljqPDfCj7BgfYhjEJyWg+oZS9hbPbi3ql5W4S26GzFJBLAa
ZRnhI9Qm9ZfLJB/woJ7oyO3ZazNKWqlpDgT+G7yspxYNTgCBQYBOIlaKE8C6XDE8
9MHPzNL6J9IOvvMmFwR7wttE7YzUxFP5XBiMAg0tnCrqEE+n1ld/ifdDKKgu+kCF
uTRQr3QEvZjwSJjDM8M99QOB8AoamYaLte2t8ZdCsqcXDWv5Cuwd2Rs7waMNV0a1
WM2xhs0j1kYmijuJ1JUEcTNY7zgt/srIH3fICU4PTR9kTlAyCNQtQ2Aeqr5lXzta
6nvq6giLCQ1PlfnGT8vQjIjMOvCZCVwhz/RNqnyCLorIxbyJQQZjWJ+gnucvNJrT
14eaSKAXE+8NrITn7a8SYlFuOv7LyQ5SM3UzwN2TUIxjmC7NbS49VjbKYC3f+09K
WSvWbYSFNeh8Yktlp3Rk/tNpbvTawDG1bPZ452p5sshkATNALL2+eOXq15UCF+fv
oJ9AoylVeTU48aQfbHUtVtzgUK8li23mvKYTFPhVLK/rDTOCEvx+ahRVQsakHyRg
9JwBnatd1ycGrfj2hvB/l+BQoN8W/OiRUePxM+iTu4GJLorck9BOqCf2jxC+nIXV
CiRPMmxadQmFgJuU6nHDuYuGiAutjeAMnMFlv4b1Svd5OjHoNctwAxfLbUvRNBBs
eB8z7lTTC3DOu5ezUnyAAhRtG7raTRkNJP0Ej50H2pNVT3wcgL78oF6DGNSI+DZx
41aRAr67C34C6ALmnPa10ogKDywr8YFm13H3+cab947KJpt/izQZZPqnDxyFp/qg
UibWNAO5uqdd/OAER+tj/DQXIrtZgBeYaaXBcUlo43vVF9FHYq/CzxPit3phrxYV
J7qxIbe8ZHkUJ2jtji8RHZGSNjzjZnQ/Lmm6lzL3UjME63JJGqesxA0sZkAjzVNV
n1zUPrU62kVAOK04IudB1WDohlrGB7hMIjlctgrb0BRFUmpXPWIFY6mR2ZcUnnRg
1GghoCpn3UQ52jQCqg6mM+ldhPRNWi1n+fwzl6VDQWIzqWyGQ1Dpr1l3XRrok7vF
wzCarP46WBEYWEOjqJdFu1Ki7iMdHQ4hV6XdMfYCCYyoraJ0q4MzTMVYD395PBLW
OQLTGXXBY3YcxNmzL+CWAt4F6R/D7CAnrgKkAQpN3lpFmmIBMz2/+baHcgmtxahK
wwf8ZvH19fOj3/N7QpHZGTuFf16L8nA+bNnLueWDt+UJi8wki9oqElkcffG5H5l+
twMlR42VrpxXfhx7fkBB4unaiirzreTUmNQNzxeZqnc7exq0KQ47QCOtxLoq7ye6
LsHp1EFKdCk9NJ1ftlmelWKVIbFGfLiiGm9OgTrblP27SUqwawhGsh03LKGF53ru
f3v+ISimRDhfnQZrYlR7Jt9mA0N7E7EObEKwIou4Rlxy4L+/KRqVKNXoVb3t/ykB
7gX+nKd1pu7/xPfcHQuS9nsCwdhHq+LmFY/qxuW/NzGDK6i3ocaUd81Y4mUvo2pd
xiuRDsYZLbmI/FWLQaqQxoZLwkOdo5+jOQMyHSx4/ueobf/yvYknTz9HQspXP7nF
pdbC2vBhqKHTigsVnS9QDDKDRvrUMQf5aCuo7K0Ccs9icjOGq92aFV5mG6vlZLAU
nrg8N5nH9apxoxBRM7MzOCqSUaTfW6hcehFYZM7283e5gRbvghd3VY+DcNvfkLEU
s8TG0dDEY24dBCr3kBSFSVQADWNAs1RZjqMcsG4phGgukXKdgADRASz9Uc/B1UTk
Gv/ZZBba/RkPE2YOoZsbRGy5jC3FRphhIc3HYnvF2KhL6tpcc56P21PnNRS5aEID
x5DrdOsMsd3W/YuLmxYWa9Ah64Vn/JYXaqpGp1FLJAd+wJ06I8gCXphtQ/+A4f6J
RewY9Wj0WbX4+ztJMdL1wMaWU9+tVEUSYBNRfIC3XX5vy8hEUXqn8eUc6CKNZbVx
IeH/GyrZYg89CDn3jU1JZccDDY2gmS6r6zC3/E2Wv6XF9R7y2u3bgu0tBtxEmEWh
9XXaH//R/9Cw+h7Gf6B567NEHpnc/I3f+WFdw0ZfUWZTElia+9bNn1lDyln7nPie
f+4c2zQw7C+1viic7t9seg6lWY5MNLM+L+Fx9rs+sjz+Mg2W2PFO32b8whtPU0IL
uOloSde88kUQ0VXci/O4J7m5AO/5ijmLTfd546YZjEjCqsnY1rOTTQeAlpJdd532
neQpI9tU9jJWXKq+04rq3gdrfin/3eLMGGsLkP/61hGEAG4GnuYFoD02tfUeUX/M
udQshXcMMcrqu00ehWjoFc4NAaMLcmdixq2CsT+r6Pkeym8epTQDw94OxrSailjH
w3rXCMD8ktWQkBCd7XXZ3Z2/lWbLk9+rV38co+O790VAyYjs5gNLEv39/VuzCBKH
n0c/YZvrkp0NBG/ggScMsCu/r5CHOMSr4Ktq+Tu3Rv4odMj970I5J/vwbXSe1hUI
qb93hkvXY3+wq1pfvUoQkXfd53b2vdWxV9M97PdDaZeZz9XRsKdNqT0UD1Bzppuu
AyYKLpt25ovNpHg9hPX/HRQabQMrFYctZsMQciktItVXCe8Ekspv/BahR1FDzrPJ
rEiODO227n28VMnyKmRfQZKR1tok7N4dAjrSo9Seha7NrjEUDiDsLQXk1x1tmSH4
QWrF0ezz21OF1maLQGvUvgH7L90K1QvNMj20oHO4e0FU0M7iBjuTE91e3LPbhLMo
NBw4IDYHR0ToJ6Y5pec2H5bZe5Q9EkCAftR7KmK77JNpMD+3XIXiSzp4a2iQRBsO
XQHgOm7fhJBiFOxDHLcgm90r1wsuEkHg9y3vnvGAVBIEkI8Y5Hwra0N5xNLGVtu8
q0xAO6ALVtNBe1HprbsGsD1lvl+zFg4HYlkDfStHEFIh6cyedDQJcqLX7AtfXSu7
+3nR1BMwF948BnPH2l9y3hmRSfqnNT5P+PV18aZuaYNJOX7zQYo0O4YRevJE9ej4
97QVUAQcgFRQk5eXcA1cGID95ZFZcQmmdgV5DbITSeN80TrcJRQhaFHvgXzmvZL8
YxutW1fDd9xtrF33Gbb8N7wtkE8suEqNuf74ww7FQQUOBEQyScz+5r7vzwA5PtG0
UUmciXNcNYYEBqufHwMLn7kdZGAbtB+w7Rbi6qdfwk9+XbMljxkZTONUhnEkIj42
2WKwnTQYJohjniPm5ikW2gqSTeT1J6D09WEZ9w5piSLBzsHinL4ld+E+je5RoUY+
gD1RARtvP2W0rBhuginE76ikbYbBhZaKEJNZPp/Vwyjpmoj1WKq395EFDs7L56Oy
gHGA96rDfcGXnWOVAsmKNJW4p4y9tYYWJ8CdDCECiYIMVoNNWgYlJDNkcu9dBzoQ
6KpOzssR9qFaORNBhfPmDli0TGb5sDxw7+wufsCbEX76h8qP7egmlE+GhWNnrlhi
4PyYfsKCPr/YkNjlQLOYJIKcFD3mInSetoAEYKpwYUHugNwAqMHxZJy2eiJRZkBm
rLxu+KtftcvUSve/DV6aBlezYmwmasw+YDiJYBwDH/xdK66PP8aclhLR33+pShO/
ymx4mdq26tBQLjKAGN+xNogDRUFFB1CMvbMovYmb9FHZohxnfAGUjvTkXc/P4i9W
g+9oDV9TKXtKipjl0pE6YvBhIfjUAlSjqsQtbbA3jBt9bY2IB73RQwbx298koKQx
C+/rMWKQFMBjLlKiAVrNa8zUr1VPrrtmkBijOO9RF72/tOkJmUNNZuAyNADdwcvM
Tqrz5emyByPdbAxaBsFYnvGBfbz//h92nQzA5IVMfVN3Ga0M0BITrL00WreYRoS9
nJG/gMNB35gzHIJ9BGvs/RZKHS3DJmaS6x7eyxfIjwQjDXfxVCGnQaQ8immmvlGm
6n9cWkPJpcZIpD1Qf1TFws1YLaaPO8fxGTVbO7eunc4hBoT2pKbMeNfAQbPmkT9j
y+nzsB5M7LYc2QQfFEFh5huv5hjAoymy2bcVcLHzz80bkrUq/DIrgh+p4cb1emBX
IMhMdTjZxB1HdB2gjdWTeDQ3AAmKXSEcaPjZ2B4aw8ufwetJZLcMCEV+bQsd9rsA
5yDSZ+EpkOpgjW3UZxbAYKGNkoqPp4j/GrLAi9pSQPbzAYyJKl31uUC23NC1l0ho
tm6Hb+zTXMZ62Zcc6hbnTlnDIgAaXqgzCymFedQPjvF3ZPwaSJ+9T7yxS9bPD3gx
dwibRHWvgxUJ9u9ocbGMQG/Vy1I2S7UYCa9nvYW66eR8HDx3vWMPtR+dSWTBXS/G
hNAAIZKv56kpyAnSrSlC2sJcfB07ii8TfAEIvwWBTTrtXHAI4nVYNuxF1tdPDaVO
XsYC/phRuAPvjQweKXghUOdklYNW+Fw1VUsVi238l8idIG9sgNko1g3huosAvcsL
ZEiMptnd+q9aAZC6GhOEy5kMOiV3leopX1idpWYwUM0XobFiDE24Ustyys8vDx6K
Qm+atvGdrHIThv5Yp/PzNWi+QZN/0Ss96CnVuaOmoO8O63UGsAbd4GnLICwkfGM/
bs9HIl22izKqeubc7Q1KcHvie1xGX3CgdJTHCwIUiudCFPTiv20oodmhwJBStSgu
XeyXjQ7TEhJyVlZbe5dU4tPFgD6LSOfhVYdESz+c0patGMdh4et1uWBxNT1r89OY
rXmYRl61KWj/2Ezv4A2aLoy2dhRDRYRik4RG2bqq+rgZDsWzJGt+sUfbCFGFmBLD
0Y3G7yjcfN+V0dWbNaAh65J33K2RYAbUBsJEoiVtfbOS6ryBUfEEEgTng4R2/wGD
pJjguskcO8cu62NbXqWnBVI7Wzpc1OO6dFGJjMl9+aqqb3gvrvJMYavd8+dMt151
gKSIotMT5GeTRcfVcaNiajWOEwAQ27RWAexnhYd57GAL7WsiTlldtnFMJAdbPFOx
k03cfzdM7soxTWNwMWFIHKbJMpSD9tJoMR/Y+1D9Wk6rlNbrp0u3V1goJ7jUsGf+
20jkRnj5vhIMqZvyY0/VX6p99HzfhlG8O56M0YEGtdB6izAfMhtL2XpP1frh2aGu
luslYXPB1pDILs7/bw74JKFSLxi80XG6AG8H5xcZcBNFxL5G//TlXT9xvAjyi4Ek
E8qyT3FMErJQqT4/7Hu3ARZuzza+3cNQ6qyltS/kh4KZl6+WF52HWXQmNGu/zgoB
x9Yp95BOp/VnN7MS6dAjj81W8Sjen0LdHtsfCdlNUBtxIfy5H+qleez0+6pPp0i3
CI7opkWIdAbpaMCqGOx/4Qj10G5FRD7IwLQMt9DI8CyDvt8yYFWWdvYMQdbpn79h
OTT2eqgceuKQnGFmPZKssB52YvnpPvTMF9MRxu07971FaGMHavaQvG058thbMqMm
DCtjmHa7y7JxgAnRjVyaB6578WplPu30ie3DUlNG04DC+3aVauc0Y+MNA6yo9y+K
8ZWAEaVAPogt8DQylTYfG92XJnEHNoG8wG3Z2NxYQAVXhHcJ++Vh1w48lTOgqCbq
wp8cqDEMNku40f5iZl9nfHo1UQQDJOQw0k8JoytyW6wKMUJaEK/9LqomCxo7W76s
CFBTeFh3gm1WtmN7DBhmVyWbcpHxlkn95BfbqVZcy+JhkyCYEZt/Xz3ervie+dBv
eqoJZIMAgMMutFrwVSXMyR6H6hMGZh5x64v/nDDT1jqMx349UJA/sabfq6cKzE4r
EoAqPQY6xW81yRUXlRn/35fcotJdOlbPWYmI6pHCkt+vGklzeAQ/5+ZEw1xmJCxO
ByRQ8e8AVYtN1zLUAoE/PSCsFfn9LbWPN1bci/BbZxlguaup5eSFNQGso/XxfAbU
tU77VbaK2wMhOADXpW7yRZPRF6q5JKGDnliBcmtgQj0DCkhN9K3v+WFKHB/aljrN
JatkLT3VNLcZ2drZKAjx6hou/DdJQ3tXY+7PbhsKkK3KNFS880i9V06GU4htfhzN
/Rh+G+WIe0TKBWgNAD1uR4ukzQw1+NqkAYCVciUqgx+ib9B5FZcKLAMfq6QcbkUf
Zl2hZOueawwTesWfETnQNUmDLvTo92uMDTm6YgBqXXHocfOXXgwK0fCuFTlzAXg8
yNcyJT4/8u1VhKpK9s7f+H1as7cxb8pEJ85lgY/STmWeSdKkwi+5PqoFq4BgRkGE
/fgtXsZ24cMAgEkmYWF5OCwWEbbYz8o8O4Ebc+0zWOJcZDL7HLbWK0xUFpXF/QZZ
4DScgqt1aCeugudnVVSz57CR9rmJlecnqYadfD6U5uoBUM2tU0ags4OVgaHrJcJS
XitkbVymYg9p8LQt/jF1N81kk/iWoCzU9UX6EQQeldK5rjmvrHSOSKQuEmXZBXXT
TRQ8BJVPHjTg3iCcVXxO+SSCWNPAuvIzbGyXyzKIpAXLyzL7zY5zYVKpG6BG8n/h
Qga8FQ56IoFmSeBzwGYRNYJiqKJ2Qi9njOiHYXppwgYnt6fJgQn4vJhaugJGY22u
A7hw/3GrnQcFVDNpFIGyiPFJv2yP2Ig8P+5ID26Qgwm3+DGHKadVkf7Vhqa2Um1k
kDqg08PGB+ZNGXQjhpvhN0MPzKbcD6LkHWl5Il3T4ROpxRw1hzVPCVvMPvRE7Zv4
gVITo/7Qa55l4uFmbdUJJs1BocHdPkSPPt+Xdg2kHEcuzdmO6334PnRkXotI8ji5
TICt1Srrx4tGBpETwz9CgIus4XUiS79RUHjABk1UJUfTk6xbMt1RMZCyuZ3tW94s
4v60bEx7b785Qf98JUzQR42ymbW594fwAvDlGRARx6695XotyERC/AXWjYq4KO3z
5tmy4Td2JD77Vu0IWXuLd7rxEwaW7Wdkz6RUXDbC547Uvn3f9I9bS83DLEPy/JoZ
HuZdEX1UPXaI3SCPBCD819eHIlXpoL8dGCv3rYSf3jOGE7GXqJWFnPwC+fiAVQ55
/5bgaUBtdVV9ckLN4khQYqU0A2bpVp90MQLVaGy5q3Bog+VKcC3ruU2uBdrCiDbo
Umr9NBraKFavQibz12BzaLjtpklRZPnPYzrGHeenb/IgGFqTT+lpYufw/pTBpJnS
jOP+vMK29eJVPgF7Fqd9PTocX5DG8x70xIWRkiXee3twff3RpupwDn/TTO5OLL15
zNivM3O1kVVDwg7ejW4nU5To+gcxvilqZ88z3dCOkT/j/AUYMpjQNUNSMGWEzU3F
dq1TCmF7uY0fpYsil09EfCeJokfA+VnKpoasw9ae2hLIK24X7Z7xOMuFpfv+MmJP
8GUa0zKdFmFi/iOF1/pdT/u6ss2aIHcjlgU4acOgb4dpP/DrVg1XqHkgFDzMprNJ
o7ODdNN4zI0eiDGLU8g9hEA7+3HbdoP/08pU3TtJfwXDexmEyyZAF5BgKZISqIo2
nZ4eP+/A0GV3nMMFqSFduoDkkQ3zbWSzzHBagBjJEmn88abnxN05bVBjHSXmF2C3
awHG62Y6drnioxZqazOdiEBRy9xxrZHjdBbORDLFb+9r+/E7WnOBkeB3XIZ2CTV4
dkUfb3zBtPvxx5+3+b7IsTHdirNtNTbilGu5dyajGtxrG0w2OarXJ3YSaFW/yxkA
Qm4US91WVVpApyLOZ7LvhgaO2vGGnic51tXRcFIdHCi+LuMFM2NPrXSsXXUsajt1
zdCnkf5a+xVbOSY1GcIi2lgE+vqb7NgkDvF1MkCIYw1rfGKORnWzaMj16NrAPSh9
Yp0jbzQQGoETAZFQG9M6YA8bcNoZjKrIvSb++e8lqOxo+JRqYFOsZbMy49AN9nC/
QAaVntwpzYTrDWYdGUOWCwT/4BV6aOn+JBbnNwLiM0FYFeghh4TOgwfMkFlqOKl0
0gMqfXMznCXQUzEmqcKfmfcTavvfHVCwDmQ0CW6NqNaBk5deLUUb3+s8eFwv5dZf
wQuG7Z7U1m1lvzVTuZTLDLm2VMIYF8wy1YAw89W61dA6GtBRyYgx6bs8poqO6roR
PlgrjN2H+p1MVmlY3j8clRg6hIttC9TpY+ZgH9sfKK4CrueU+QNayssttIZitxB/
lq/r6osJkt8hSUTUk1tNV7mLKX5znv7L4hGOfPOoRitYqSf+UOlsaB0/74j2pPuF
i2y1wU6m/OCsxij4NtQ+0oG5Q+0hDj8SfS//Idm/RPbCH+6Xu0hbPvzhjSoZvHZH
F75V3EprsZLlnMoLLxyNNXQ8DK9TSQj4LWvyxP8acSVqQCdFjdpe3KLS1shGKzrZ
99QqPyhBEEiOdOM4bZSSWuqZPtENuqf96K7C3Tt3oYAbIJK0Jr0y18kTYGajAGD8
9fz/ZWHNdlQ+2DfuLGKUvc81yZ8U9eERt0DMnF1M/CFneOc5a7NNjzpYUipxdblr
iLg5KaQyDZJbBDtkWwoInW6kKUjNfeRNQq4Y4TbkSLNTyHe54/WxYHMjKBR0LvhX
8zwzNLvpfA4W4rRT2/HKBF0nTG9yR5oEcGexDEX2H45GpRQW3c9+BxLw9VPL+xy4
oczLa5uVzG/k9yz7IznHdTqaAx5T1J51253zaM1My23iRLE13dNpzqrhEj5hAdfX
ZDlC9cVZvbqxKdKVInDzynqIo/OZV46UAGs3jtZe2uJJKRPvwl1CMxVrLw3mDwRi
J/kfezfwDz9GdH4DU+5RQK8x7PLRpoRTnef2/8RXWFm0l9iXchkNW01fMMgLMSvM
tG1ZR0oGO7ggPcBq2KUA/yDQUoiAviVptfLrOXg7XlwIflteUub1zvsj8DGEY/lr
KQZQyZlojI9Crwhu2W5rKq5tI/sDCII/kXw05Z1ubWRGeogBWyw0YS6rhILY7X57
I45ktAj7acbbqfD7xzqhbnSsAJugFHSPYYaw876JcG4hhntMZGa5JueWHC1jJ621
Z5MidsyrQU5qRmNIij2M/S5nbwN3aDydUQK5S2mR1HWCESgEGNoF4cCA2AaKddKS
2/ptj4n/NLhty08BwMRS77Ove7rfwJxHnmHfjq/GFLFSrZfRYPYHElWlxyrNIj1W
n2LImImDXGloRlQgnArBP3yi9FxZKq/MhlxmhbWTxOp9vnGmgbfiFWzzCttsn6QT
sqmA7KFWxnMNH0SBtPRvlKRzE92SL+Zce06OiFS0+R8OqOzPiYrQr8pE2WA74Tea
DMatmQ/j20KuKOm4Fw8G0PeQKRmwNZVTzTR//YjViHdxna22cC8UbPIkK7eHmStY
Zgxfvtbw6fySU+VfM7qtvnADjuMZ9NVWamp3kj5ewXM9xVgYwXqpn+GW3b0zK8b/
TxIzOKS9KBCxmm3xY4Rbs1gqcZgFzQ+WXYCj6HNbQ/C/ZTzfNv8i2TMqGtfKqwzF
4SMWQCxK49E5WlUqqFTnvR7LdTUU6Mx5IMCVANrQ5J+mXCejmoO2Nd002Ge248/c
9JDI3x0NnX+qlsZbu7k0aNi55oe6OUqkWiy8MQmVb8bENBxdHz9mId/nC1EAgofa
1lAc+0sT3TCXccvj0Fgi+fSpgjtbzYjZEEO2BWwh3UAF2buRV93rNA4/L3VDtxgf
POIPWx8CrIgWZtWN+I/x6J5bgHo9QsH4lQfyi9/9G5r6LCYb5aH3/sNDIz+63EOz
ukC6yTGW73IiHjgQMNPwlrYi5YDeONvhv59Sg3gc9d3Z8LWHy9D6GEXwP/nfEGeM
ocs2KlxoLJoNzAO8ZsFkOT0Kf62lAnImFjyBg6mMRQHVa5oONme3y1IYc5E5s4EF
HmXj09gRIW0JY9/5iKZwVICwlmVlDMI7aHK8AzQeNAxiPomks87f96MdtvxRi9lq
YPnAutVQxYCD1v0iVI5u/n4lIJb9Sp/O1r69MIQhnlB+9SkpQQbn76wo6m80DY0W
MMibDYgmLaI9d4w/ZnEnVWTU1FBVtlGtY6eGuIrjPMctS/OUCr528ccDwnVY7ODH
TOvMlVUfQjo/DKSm2SJuG7/Jmd3g0owud6Xc8hwtGgwuBjJ5iy6cpGtJJiRDveD7
LpH0SRZZv1YGTfOAog91N23FgOVaDFDYYNcMor8idkiLZEVFCWPtc2+05rxzogOj
gqo6mEOmrc9auSNN6DkFKEBaseHvSE6to7rJ8By9p4726O3QXXb73E4KRk2w/Xdt
FVfEdPgKDrwCB1choEJLzCU4LRqE40pcyOwxLZEfkCucZ8tDUrE0GEAfsV0yazcQ
yBbkFPlyz9lNcyS/jmV2cnZUzlEfaGr/5En11tsZ4tJkFPlpBW6XlD5TgRMMblTC
lxks7evQUjR8HfbXJ8xBGmXnPr0OaTzfifEr/F//HREtd+pz9iUVv9tC4luLysUu
S87cuUvx+Pir48R14lay4K+OUgBK4zgXucZrHjxT0GS20sbQYiGvJckjonXiBmSr
x2i9/AmjHvggEmq0DLgYpK85VbBs6p9lsWK3C0l7vQsdPb2L/g/AZVtGeWcaiDw9
2pKpx1vprhxFddLLld/YAZkLuNqoDBt2QRoAowGcsBXwhdBa3beNf7MFgEzEvrjg
oxe05ylFOgN2QxXS8Ew3Chy17u9GIQ+bklR88IvwKl4SHCci4vzeqJDCGSwhnfHT
albcxTGdXMRSghqByC0N4fOt7lbXX2z4fE8sRcjaA1v39k3rK5m3vXf7ST1RpuUg
gcLiajEjvNijpfX0SOP0u5g0WSqYUbHdNKxv4E+b5VcMYOnpn7YC/iBGk1PKN1pA
5MtzoZn1AEghQcGymaifLnGCrmFTu5GkXRQCqgcUuFwpdaoeR+UO+QEc7uYU/LMj
y8ASBOPQrPpNtJNf5PHYOSPC4Tu0EjSSC5AtKATMF7PT4K3fkKNQJVYox4Gco0l4
ipANmtAL530h5z0zrOuHpE/zf6W1fWVxgJQYAA/yZWSicGJ0g6e0BGc7XE3y3Cec
aD2eLvSZAWPj/HNLGMrF3eAPnRrlN23aIvmVXdGiERhzlJI0V/mMgEihQnetyDRS
ym+PAzIMbw5XAqvebQCbTJp+o83kbqRAchVAmeQFe1fsIXT9VAF6lg4zjHGVYxpW
ZLf1XFDgDDeJjjkLDQQkkDtSc7d+k/ZHQwRfuG0gL6EL0Jpu9usxCDNzW0omz5r5
GVJwiAqgb9Z6/8DcRstQ9d94YgKM0k1iBiPJDfpyQuYawjSsOUIDQT0Yk/aCL6SZ
sZpTCoUEMdnfJ6/awtFewBNYini9Nff2/RJydZ7KlVjLzf+YQ1bMZhy6UaTAMe4j
CFFzcgvi3s5H46xAFArBs939Idv+0d4/XZdNrMGJ+i24DPmRDbpjqwWmWC8G7Tjg
nXyAROEuAIGzCHnJNV7ReqUUWzHFVJ9JNlfMBKQ9DpCSCh/De73BA1t0LDZwITwi
6Nj5ae077M/piITmqa8OmcNWYwAHXjYMGIDIJMUg69qks75ZEctGhMeFYeRP6HnL
Xn27YbH5OOMvsX53mbgSE3cpiR8EK0oC65XFKgsVL2iHQWUuNncvJR+HLvgJjAPG
2El9EJpCfU595SsfDHLuJvAos/xWGSnu+PznFjO/NfhJPFGaM6pF7hAOpXxdzXVc
xgGoerV4Fs8krGRAjLYBE1OTk/3w6SCpLOnL0qsWsYXO+kBc7c3h3dLx/EOnem8V
GaUxwIyJ9fy+Zd3rPZHBxXd79JAAHQ2nvMz0h8n7p8nUHn0hnQC3XKhPF1YBINZz
Dbh1EDaa74KDmhj3Z7oO2ARnEt9/FLcOoFN5OZB6VsniJZjIueuiS2lVe+aDmgx+
AvMxt3Tk2MXtgVINIXlIXh/lm+/qzU5RJkT3lwvNkOUwuGQhEuOOezKuhLyqfpqA
f7qehUU7xbrN6nDhSFAa2AJUVg7B7NmESqQDTpwcpQ2bVei+BrAD9GqMBUqjV66H
FSBij8NRx3iN6/y30b4gHpbJNLwiKEVF3r0OEqhw3p1PgGBF8VR9IwJhbZHccdS9
OraYhlaSRHN2YarigLQD7apD5Vtc+K/ruMJhoO7DVhFZIXzBTqpgEF+QWQ4CaqcY
4DncGuxQmvJSHhJUIxHsL4dlCMajPh0hwY30/9QFU2uS7aUIoNlqtT+gtCy8RVOA
XQqB7yNSGWnQebyQvM1KgQaUQ9p+kvC/40PGZWBPxL35mly56DL/VAAjHAfB/5Hm
6DZ7x7pdxkNkD0p3v2j7k68gcTTzywiwbR4JYvsaVLleOTaPKifZLs89eXa5a+56
ZxrqcAeA0MEwKEzKOT6gjOEYq1FXXqjZW6H8qp219YjxK6UAcoTuLLmjinbYMUFG
/VWYn6aLqpoMaNUi14LbDJMYJiOu11ano8Vnk0952sY0oEBxvLkRniDlM1YsyuTT
7ebovbC6UmldYVeOmN0m2X7J+L2peY4G1YzpiQlxxcfY+YANEy8ES9sN5sx8ZVnP
zLH0GPXik6lDFm4EscGDAJGLJeOREKC00eUDiCw0/WN/bKNgIf+z11pGVKaiSAyZ
atILxm9j1HZmn8vlaGJLpR1JCLqppHinbkYc5buPZ+bFZfg/5pL9GyfoBp2ukuTB
/OZehi03BbmbQYo4LV3rMF9FT/pD00xTmT5HZRn32lTrMeQlI3NIERf6t4fxPGjW
3Kc3BdFM3FTbajhZDT6o3eAxxMYQSaS24CMsmaLi5ihOS4DCwCL1dbuqCLC/Okxc
3STMJQapNXyNvaFl31Q++f6PxcSu9yyN/U1h6y5q3TJDcocDXndX852g3lN3PWjw
nL8uWe54HFABYe6df/2+apeWa0CnxdMzSZXK88jahoONVYB9EOLJaUI8jHiQIbQX
QC0OSWshrPL6lvhwhCLNSXh99ARLbOupou8OKWjjt2ev+K3BquaEvw9OofiHwCm6
ZIYVXI1lqwWp6CGiMTomFkO0dMIAU05eM/px7fbEwtzuJk/MJ3rtuYZ4jA7nwnH2
GVNda2zWd7OCrQ/wZ1rBOEgm67nlc2M2v+l1irFiwnUQvHAiRRGPmCv/XFWBGIUf
JpTCIErdHf5Ddfra19FGNRH6UpvRod/yrX38k6EwevEi7VF5aqnkFh+9I5ePShM1
+K1oH2ivVGzBMuW0hu8q3oDTjobDB2wsqSt/QoRG2kmD8crVXas88rtOdTgSNChe
FT/iFn7m9oVmTYHfQtKGEYwaXTEZj7TCwjEys8blj0q2ES8pNBCnxZCTKyYyFTt0
GJyj9Js2Q6DWGVCuDX6D64lXs1izcotqP3xy2JMKVdtu7rgB7r422PxvHtIHBhfa
T3OjIRzzeldlJkbu8hk6AxOGFrwAMULN/uGdFhu7RftsQHRHaH9idByl1oWdBoXP
g8NQZlp62Kdfb0dvVSWfEF/eWwFLXYE9eErsvpKL4HClAocF21DibUJfvH5QmVz8
/62sLp8MT2riFv7TOxyZkoePKi4t6v0mza5BClTbuu60oIIgRIRTrVkqGyBovyrs
J4Y2zJ1vd6vHP4pffbuVsBw7ajYvJx8ezC9F0q/q6nJl3pmwzyPJTX1VM/dV7bw4
CW4nfv4DuOdICkK7AVCyu3P5yKsr6W/ifd6IvZZepMXbBHegPpOCTcOM9UzzdX/F
Ik7EAFrHq927QkySZGeNLmRdqRQx/ErV2yUQsotyfP2BP20gP1GGuK4fd/NIOMo4
Ye1OvNt7dai8sfDS2jr7eSNPV6GM7mjBHoONcqwh60XvG3/X+M//CCfW07m6C/AB
FEWSKZyksvtNJphVnjqptBaM6vtvI07NoXALRE1auQlXCb9KqjQ87jDY6JfT0P8C
x3XsqzS7XShicNnugRrswv37qlT+sLCh2tjQbR8g7xBJbJTDCCVZFbnSa2KuCLNL
fzlxBE51WnlrweDVNfJSr6GkHbmjUfCVux2cMIKZx2z5J8zJhiWqKfLHG/XsGhey
Owu4ukpLZ2zoFMgRquUOYw7HTAKZ+MAP/gdlhDw8L7qCFN+grF2IoJEOfzJRsnkh
Xqj7ZVmWxUHkW6kMCdygvbJNyGm7TDDKYJ29AQFPHfXyUMavl/L45hNoSVOkKwDn
8md1ohW51ChzF3LrigO3bVgPN6oNE9+BicLUiIfTj7459rXDgDzIlMZrZrgd1Yc8
d5bsdywrY4yZ9Hvp9fQqFp0eFnagomU0gQMd9nDxH8qEGVQ2gJhWGPWOcU6Pfpxc
RVuI6PgEqwTA+m/D9uPwzKK+7fkeL18zGQ5V3lDCqiqfpETjn/4FyQb+S6s28M1C
4xlKssBaGefW8c4vBQ4BPLPtmvRKcfNi+WyJZC2J7g2Y6pdG0QqljT3lyR+N71Cw
/K3X8T2gW880RrIvvAgrGzHMe5Ib5VmRVrAp/+kM5dFg48i7pK+kRmJ0VKC4600h
1E55zuadciO2Ja0jw73b/Nu2b+EuCZZIZHpkVnhGcOESWoUQfuSQXCdEqfppiwI7
MD8mysBvkldQfgzZo49Osvr3Z1oQY8rhM97XpSqsbdGboHtVwT83tKQqFY4H1+fu
yvNC549Np8Vxf/Ic/wmkHIrDIsy3EdjKiFq7DR0vnnziSUocObsKR7qUuGim1nkr
3pq3xawD2pzUlShKbeBIrvsRmFFQofLZNv+nomG84O1oUd/et8UdYE7PrLyCdi76
gQ33Vn1GbOy5lEV7Ek3iAR9vJLOlqQG1/42rhZ6en06s9hGVzvZquP4RqWqrhrj7
56EuW4cVDTXA/MocdPI6jnnXwV4uYmHEyEHRwTYKlpsMlRb6e26gp48lsMEDvODC
v7uWWutD1bxNFcCNitW1nGG1Lof3y8kEZbfWvSctCmTXrU6EPlyGuFG1pI/I+1n9
4tL4EC5e+CDS5i1STmzZkaUtxwnQEKeqjBSJconBTaFRlSz4Ng+xfaNmrPFT+1UL
0leW30nsqWz0QFArD6wVhymYjuomSqup4HXkP6CcbaY5cbfUOJVWr/muS5iXVguM
4EIX8gzhoBYoGBPs4TjM376Vb2evbeh17VYYHEkqyUZ52vj73XnQmWGL6l5GvJna
kp/Tv/BqnUBAG+qzN06EoPXtsnv2ASTmX3USc+aVqjDR0TQ99YBepXsL+MmUt5aJ
nYuMHrzDiiU3IOP21+uJClT14ECS30Kgr805B11Vi4dAaB1kZnNB+iRiwtqEr6QL
FS3U7xA2Qu2tJV2QCQYN06hDqYUdMg7IxfpQXuUEY0Q20ZHYTGA7HHnYzjvDCgSn
oEgHDfqMneReR56ZPNkdZ+SpJogQvL8YKSsTS4LlaIhzuqBXBoSdUk7fZ5p2uJfm
PH8ZFX8l/TZZF8/NlKA1wkS9ZQo7YI35qtCtHRwTcIP78XdjzrRmsKXAGiUT40vZ
kqddp3ENKhHvwLMviL6ia4pEXZA7Q5K3YCaeQrZCyGR3wrc3WABijHWbbJwdxJCk
Kp7lG8bVy1+BMO+9zrV6+KPyCM6H4Xs6edgMiZD687Y/PGygyGfTcSWDXSXiUceF
iICI7x36sg3+NCyRuNPizuycDp2gd1AAnmhMYFTNsJLXkWvJ7U5Nv1kqJrNRREUp
1Bnw58L/7NXHubf/tehc+lRa79TmPYYQYdKUU4X/LXTA2HfVZvh2GucROzkz+AxT
08Rs6FlRSdM4dqmHNeFoW0sCuTTeeIJfaTXA/frxppBjrp9uBwJTK9fvRaWanIeK
1FGakcg0HMWdeLIE9Ae6FbuCfXY4neBUbUus+bZVP++MwU//qQzu9c39tmy0pe/8
C0Pwxbhc6lYJ4P9qbgjmNendLyxsjgy1UA2MlbPwLJO7Za6g1OmI43LjwxXixbD8
7UHED1+uh1sufuJN6QOXa3yc7NSqouofRjb4QHfyfJdi2XCNcnE9m9tOD17QsgIj
PUbAnAxd8q7RwySkGZ90OSaUx5ScR0rkS3yjqngrleT303FhXIXTCedU7ISRrgE9
5MzRvNmPaQ26ohRwQv7AR2O5ryqUl7jmUnZq0PbrrxT1w6DeaMm6RS64ypFWgof7
T46A/z9V7+ROl2un0YT7TMpJxPTamydTgngP7muls7JmFfGphajJ9PVmCSSG+x6G
3Ai83tWGafxIK5rJ2psFPHiiVGz955H2sDQbHjwnW5JBza26bjAMd+T73skYD2dc
aoO79ZBrKZRG8GDxjTLbXb/AI5k6kRxXYXj+ri08VDqYD3jJ0vZTPcaolLlR+1hy
nH8hS5egoqyx/KZGk+qvp7NGIZrXo6lTwaw1OHVt08oucn4aId1rrfq3e6P2UtGW
dNEg5nGPel9+n/K5lnzcokJ2LpRoUqRxu9ZFTa9koq95ZEJoUnkvn56wCZYyk/nC
a3M+NvbbzOuSSfa0HR0ZZvxKSYXB2Lw6FW/G+zAJTEKlFj8GnozsswdogdeA8lSi
mRaHti26gSIznJCRewGzLjnZscO5DqcQiHeHD9W3N4tW2wpDMzLxCn3Wiix/hj/e
lpcLiQtrtUYS+CDTSUnMM47fPK2L8AEeAqR3k0cyeOo=
`pragma protect end_protected
