// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
nzjVMLKUwvMiRHayRW9XlB3/YXCM/7z4lEDrYJGPLyCClCxCWVrLlNpFPNSzXlrWDooZq5JGvU0A
8VjZXmJMMmzXWSrqZRuFVUVm1l+J34d8CiFYChLYv3tztP0IKCG/yCapBuiFedGuDOWKZlNIld0t
CU5bHvRLBtwQiZPyuARrTT07OUjiAv7xK2zacKpFV2vms6P7cnkK4HyFUHy8IG+I+kcciFFgFaxp
LvkcHG1WodxoiDdhcKuZr4b6IWOHzf7vxRKIZvuu4WDwdPEkXDRRoSCONAutoxuhjFzof1RnROyl
scL+3F3m2qRqG1GrGji0DD4J8zcipH4BY9bTDQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
IaN55wMQ+2cnALAX8s6cHqEAjbGYnvjUM/Kua5OwdCS3O0mqO1bHMmFBqp69SAD+3aSO0yJWHFuq
sTDtIDDXXXLNIZa34MVlSubeC6PTTOt1jrmvj27mqJO3GSHi3/MdVJCLnZc3XgpXFgYDJK+tQow/
BFdvW/fkaeYisVXDqo7/jy5XRLBqXHOCbS8Z94ZEqbgywBj8C6vQhFQtTkAV8FTdwovz+k6BEJZ8
OW2oHuaCPZSniqR9zd3O8Jh/9PwTgEdhzjnLJODHutkbc9/mZx85nNYN2e3EBYekkO6JBJh154u2
PMwXjb4LARi9DD4BLJ7iFqkwl4Z7og0TSpKte/1XIp5QAjUnAXPgvPA4//AL4xzjj+HXl3MieRrT
n7rACovT9eqCDjDffQ0flN0CmOeMWV2FE82CL4XtK5feEbDfZpMBN3WQ91Vwkb/oVNiM2N82Cufg
7jr7sSrlSJVehrClk2W4z301wC++cDBTYWVnVydcLmA7DmzSYbtZN02CYhIv4Q9ZslgmRHvYg5nj
/LooWG7ECOkl7OP+hJSakoS68nDz6nqyK+7elr1EzGupoPag282s87JmKLcU7XnDJP02gdr0Zr0T
G2iO4e39quj946C1YXBierb6yeNhMcE2wzBkKycP8qpWoijLnh3rN2n02mmWBH6F/vRYbDUTL8Rp
I/5tju2tTVrF1QecD8WK5plB+31lxQvR+XGC/4kHNYkRwHindVphNRzpwT9y+BHHaq1FyHvYW1b6
ra9IHRjH6sMV7WFhSSBRjGWCm2HleUy/diZ1wa7dtb4A2HTBJ5vUCq7AzvQHNHoBmrxI9vSSOIiA
MIBq7bQtsFraNdfip3fvV6E8/kiR+JizUvVNtvks402qBTS7oksleHqqOzel34uYdCnRISEiOJV5
9r62PDgID1vkNBTAkexz7XHyoB6EzKGs69faPkUrwQab+/g2SYWhu7R/sYPF2kFiXSrzPnu1VgHV
emyMqumpqC/+fSag8UXS+d746hEZrEXnWthXR0wjY/3iivg92HqRDmj12imVz+0fB3te/bzTgJCS
msjTa+tHZV6FAKnWfc0VvjgWkgnDzfEpTs5eS05YB5UiY4xvd2faYe3IsM36SjByaV7dkALQz5hK
QD5+8Ubbl9cnHy+ll85XwS6jOxwsthpC4MzYaaJ+tNlP5mFHNFVkZ1oCZFo5kMnmfPiNjPgw/iV5
+wOfyE8NMxP69+shxgCr80PjE1S/3CBjKNuhv0lB0EIjoVxg49NhKjZcabQFBlutke0icWNBdhpT
cklNPoQEaGmkWLaTuBORENKAz+M4zuIBMbxiyMcgiKEiWHAOHGq+7xF6AVWmVRuaHE+tYOQ3wR+G
U61BtKBkl2LTzPXVUoVP7i8JIJYHSf1tR7Jln8lLSXzOhYe5jK/VKZEJ8Yg9/VUbiaBGniRzS9Kd
FNjr/hJKdf/RZCpB4oh/rWTtKltzRiPnwukNsR/1bftiks91lQ17g2uTCV9tH3dhIVcyszRqNnvQ
xfoWriKZLGp6aWBz8zlaKJaiY4laAyJiJGqNac4z8Nxp6Vxq3AKapNiVzB5bajv/CVVemUD5X8LA
IbdBztKFtJKyt9+lMM5Ts/zWLnjtvP7Rr+wIMX5+sTQs6kwFW1F4WUMYAsT6aLM9m9gIvBNrUBvy
eqyz67P2ENfxVtqDm3I4oximBn7SPONMCdsXdc/FpLxj7ZzBw/Lv+XlBm4X9m2fX1jZzQRE1vBTD
f3DNptkdtfqRajX9AwGoCUF0P0GOvv6YlrBVxquLim1tYPonWgmBZT+ta4HVg/lLboMBtYBh6o2X
njbpwWy261b0i0KwobMOIHA6VM6VKYDyL0G2k9DJja15rsmxogunOwxxV3rEh9RIRK/+4Ywi0rCS
dr9fKwXsaD3Gtec6/bx2LQJflkv1l/UrBA7EXQPhlyE1Hrl+8WOVI11A/f6BEGW7vsA7jEeHm3in
qmhZb4duDnh68wJXvZSGjQJV0yx4vwjeOtKbnvqpxpOLu1Ku1RWn4WeFF0rTWgjPSrYVQTn5BSB1
jFgAFaJR+lWVLrwBthWCv9kcuoMAQEV+Nai7hX72pmrZomwAoRgCC+vMCrjQp4QhtTH0CuG57lLb
cXR9iON2HAW8uHCVPBOiv6vLkKNbj8qZf2eX0EWmUMWnoU70AWnMcIzlLr5jGavXb+nyX1c3TYEo
Fs8I9f/Qd5iluNKwUZU+gmUJ0Og0oISA5YVgnKjrA1JJltmE+dBH5UpuoqR3aVUC8STfdvsL78a/
3wMHChJ8RPu3As0Syr0AqYZNzurXAtfNXmQ2uc9pyCwfkqxye8y1L3kUyuxVnGrsnAfFIwHxKpO1
H8/uD7pYd7+ojg0dN7fDVcklMlwkRheYYMC9xQYmM9wWz/423yvbG3cXNGa1TsUSgOjkAiALdU5z
GEOZ/ttZu+gisAenuv0pIdiIItnW7qa8dbfBlt3eWkMcuAn647PkvG7Zg7gaihTCzehCoN1nYC3c
C0LIPLLtBmVJlQUDZaSDWfuKUaw5f8jSJVly7XmX6yLiDneKO/wbVYKRGtoIJ+l910+ZfZykH+54
bprNUC13Keqpwzo8VxD5P75BUXo34K7HP28GTVgbMzJ5CyUhkvz3wxh68Eow6c4S22ZQHsgxc97c
fcKXTgeeoAY4Z7qCtWwbZ3d+jD+NxG5Ak/a6I0IZ11oYOkU+gZ3oUMiNIVMxOXf+V4hZizCuoGPa
6YA7354MDF6T+4m6FavofxXHwaeAaY0Ph7ZLbR51n2XcNbq0CVpSi0rO0akcyUm4Onvu1mRWiV2A
8HRIrKCIBAO3fGOnqYpBVDkstkLpL39dqNtmKWw7Yt+UOQ8rLbF7oz7p9PBttxi1zCoIaJoW5+ec
hK4xQLnU/95tdw5gJIOwjR0feHLnWYEFM325sFwa/tjzM1n2aloStPU5wJVM969FFEOrL9e/oOuo
k8llcjNk1vTQhmESwavO8UUfy02EcCfRNAwfewaX6/ptsMGotRkVCWPuLH/isTukV01WYK/xjnZ7
/7xzKxE4sApcqVc2L+IoGBay4KhROJOOmQbEHQhcnqFmBOpFEkFFPNSOS8lmyEucVaXOX++8Mjjt
TztUjF5/SSami6jo+USzXSrI/vdGkAwLVXIVB1WRmukZC8ZY06BWPy1NMKIKQKvG5PV67iiRVKRL
/wwPQWZf6FLvP83u3RAak8g5pK6dHmacQWQZ1UiYsZ5hgn1K0M5mbl9J9RgJxwiN/xrQiR6xl54H
1vp3Bfc1UoFy4wJpNbyOye1BCstTGResNMfnsYKdnurCxVvciDl5r63vhC/iqhCHIz77/58D0+/6
BaVzmaPAkaaZdeHnD95532Ym1+uPv7t2rD2X+fUqjV/c5vf9IESPBTLRYDT58VkUoMNgYprcIUAN
xjRvmJahHoZ5P1QGwVFJ2KrgEXqCSvyyPr/7ZkQVkwVqjsSCMYLjniI6KST+4knt25hsM88Woq+R
Y1ck5FM6pK+5//omy1uXxljOSXyH1chWfJ2PiT4/2LtfjVDFlnU3x2dNAm2O0tQQAe1riHpymLLY
6aqrPcS09IrqcD2blLJXmuXrE5QJfAy+EuNEpcX6g0c6kNnE2LYdjEr3OKCyMeiT1RXcQPK+TE97
Oh0q4Lqj9QpPHzCmUwP4fh9vwhzu+HVEFjXnARp5VUZYdu4o/L14RdUKYNjMVG0T0Q9VVdAqJ1I3
pjwiSAuDr9DR7L0F+I7YxOVkuUUVxlai8viyQC1oALD5XJr2nB9qOoIQxlmn7DFuBETT06+ChV0E
9C0vD/eJ8SB91r3Lb3QFkDnqWhxmbZ+YM+AWDwDihx1OYronVfLtzMOBPA0IU3ZEP+AjTqWzDDE7
bxc8ZhSmeKbmHKApRe3wNUgUChvy9+9XsitxMEDVU61kN3q3bKWyLHZXJ61OdeQG2UhifJS2tcwM
aPHMy2MGvmbt+M5ALbYRVe+4Y2zY+DniD4uzt2RYxKJ5KHMeOTl4CyVNTSrM7gVOQCh6aDtslSdX
61ADkI/6Ncj6THC1dLTg6qqEsvlPUapEDOe//byVlWodIvXrqe82dieg/vEaB45vJlU3eC5FJZqg
AqxoM/wCyOak2t1IVaEnYRZDHCp/DMaGXRI03P5UmCXqwNfYt+Tlczs7oBQV/seMWHPt5pEBOCgQ
XPrJmC368UohmlSbdfBOMhBhEuZnpPrrUAj6lgtHNHmVysL9cG5KyZpxnAC6YzNkzhKpaSY6P4yy
Z9LL30LIGJf6g8Aw9FtB8ekTGVba0RF3t7nRW/K0GQqv61dV/fo/tORfR3q7+o2TPEtxp8e1a4m2
4Qo2e2+FmMjgMtqOgaDgqbXW93SIhu3dlNNZ7Zqrz2EezBxzLVBz1t/b6JWQ4XfdbltuECAHkx0u
cTNGy7HZK6HljHd/U806BUsK+bYqPEh89iECxF+iHv1qweEC1IErUNdA7urFxZQw5S7roZ6+HnYn
mO/hUMvitSCHtjdhF+7yibVPOhAzmznN997v9Tzr4DCO1qMpr1Q69suyJaGegumQcSiK2soxgc6p
w95m/jNYxPwqQB6/r4fSlkFAXZOI1O0RZiz59foeSNAd101mMGAnphZDJo4lEpkv3m8OAW5g4ytw
XBz+E8Z7pnMKtGO02w/I16K2GH4y+IgnS/MI8/mg7L8gygq8NbCK3seshiQaMDIvOcYH/MuDCpYj
uJ9czAW+66RMf7c4q9RIkc+MLFJ0Tddrn7a5731GUp9M6UZGO7cGPgKpR5tj6qva0CKO0r1A6HV5
RDq8Rpf0y4TPJ6Ep5NB9GkmvGbAw91yQJD94Ca3Gve73MKhEG8q02ffeEXujBz1KRGb/XoutHoTE
i6D03jh8bR9kKD3xC3Dg61VOPCTUO+/F/kfxFytwjF6ywn1P9MEleLGkmU4xRVKHQIjqtFvWdsUa
viOvZOw4CCwCT14DzFsBZ0JoFLPUgfq5xC+wg6wcxIKogARaOEmZVHvEYS2xaEiDhICIhrI51Oz9
xbQhg7FjkG+Nun+KvJUKQhwhnyDkzTFxl5VZhN4MjxUKfDaAc+FYTY/cYOVGEjS7Rf3B8Pjq6Fyn
brAeMrPW+R+z7mtzg6SVVVgcLdVrPumxtPg5v2ctV5wLf+QAVvBC51Azp5SSeSM6zY36rNQHS/G8
WOZcuaE6MhXhTukR1YMHnNdv0vpFUY6IgODeeVel1rn1CklTCOsEnh/Ol+poVzrWu3pUTuiiBNWL
1TlFjJzvtaYCKYAJ3oUiWyM+ioXjUuw3UA+kvZysiOIEQAou3VJ8y56mTyBZq5HkDWXgFNHEN1V+
76xDlQy5dNqkwNv1OOtsEInd96kaD0NmERhrRSTAtBXJ7w+pTwQ/nI/MJPhRLS0eN8JQOkA9qmxs
GVpLhBksjMeajfARU+/KkMQuQ0g4uY3CEYlEucBXkTU5fybr+AhvXb7zq3v380wToyGSFsnz3OwE
LJp+wjfL18kroEotZEy2m/uChOPzcAB50J0N5qlND3Tg+elBqhz+cbIq5mh2qmJXHOVz8cjUr+d7
FSj1xBYMxZt8M8Oka4yHgSjIk5cBE1DVsEfJ6V7S6wJtYQ1dlS0yr/t0c24s21b60cUlxgXC9Ape
9RIonisV4iFOFOE9elAlc65whjSi39VqqCqfClGGkPVtf+Oo2baD4ePTDrBcgYHTA/CkDC1FiZdK
goAsmmjeOV/cLpc3cL5pwn34IW628QP4g0vNZ+H9JzeXDK/WhscqZD6mcHf+xGchDGrrXQ3ZCYnO
6t0X0hbTmElFH4Grwxi321cbuNZ3ZsFvq0C8wExu6TPtntjkO0kFb2+E8APeMOQg/rrKRiONSIHe
turZBB52YOOd187B3hHv7dGgA8J/MMCviY25x5hMfRAaCnFx86EnjIRdF2fXp25ks7smyz+LNhrs
EG11WwGszB0g1R6/Lm87+EhezinxjJVKbTcszU9WtY/2ui7LkXuRMKDZd2uCkJtH0LxzuoJda42B
t4Tcw8VPcxpFV6w+/7pEPQW2qN1WRTLxZekEK4GUVyJXdvhsn4HhhzLVoZPcCWtvzlEON3mcaR4P
cSFoMOUIzayhGQJC/Vm3JJmQrVfxvwA3PiWHOqc8ZOoD0/0+DxzYFM28mswaW+QrJj1oRPVu/wCD
rYxBG1R7xNZh8kMeekRvDakDILa1SoSDdIOjIFIITvt1Q8omMMmcjWVCIAhbEVeHJtY131Kg5JD5
rw22scnawxwuiDRHqvfdFR3T9JKkVUFnS8KjMK4laTEPE6gmw0CDb/O8g87DNSs1lN/VeGdgdoZV
O5ZgPBg5ql4/A7kql7tIp6SpSk36jJeTy7PsJGlwk9Gcxj2BOSQH4txd/cJ9OtBZn+RLqG4wTfOg
FIQg4sFsCIC/jQ/V1UFPykBanMxN5doz0jNngxi2dczVGD3K8WhK0KxmkuV1hm3E3B5B9jbWTUl7
lavU2PAEK51KYhdMgxrgO5HvBMG4slH8gd7ZkmZIrDTyX4VkdwcX65+skjf667Iz4FoSvdes2FsN
DZJZ9he4ATM3KL+FSplvafePkMePZK00/FlN44Qw/KU6iSn0POY9iP4osnLkJJET0GpZTtbK5b0z
7A7Xo+lMcmQHdE7zFAuduhMeg9PeYWUhiXkgMJLzI09DYmE0stW7QlwXJVhpYIyu6+CDIDxdza97
Ic5XNR1/K2swW9+OVRY2n8TxoEbTZj2KEBvn7YtAbV52X0VYSRnkw8l7Agws27kDN35iX6TSHUO4
h3kikpK6MEttWtqt9fN0N56IPgb0aAFvSwEb2q5hO7rRTCArEnzhaqsJLV651rcn1635rFAawu2C
KvbqbSsbuZgdZzdb6CCtoE90N/oHAZWB311BfSrfmgeBRQREOXYfiQ2gHUmqUA3FK4x4I/YOTNkN
DIlFUqNP0WquBaRonH3zfHjovx1SPQePo6kMs3oG8lhbCS55o3tSHIHywt4C1htgySa6uD+DWrGr
pEB1pUFQqrWbDDMa4hpTgPzs81qb8/vquKGvn37g2KrAl6ShpU1epkvV5RrV3NE0sHf/Q7aYjEAc
WGjTSKOEwEYm1bzysCUGVHW+EMiNYLnQnRzHcTdnMcZ+u09MAeUHkOmFuZ/qjxsg0OAig6BzVU9H
2N198eGQEDUPhDCc01kPzwi5dzjgekEmnDhzLKtUFYH/f0ui8yHlUYtUsBLwt7HBKgTZ+FRLSEZn
TwS55QtkX7IklaBU9fDx8LrUt6Muq0eQN8XWgWpr+qMJxVp6opxAuJd29jnlZYb2SUDi4xW4YQTu
WtJVUHqZfgrRBY7IqI+Oj1Oqzm6pjWBPRyiTixhgMVOsKI5qpXeWq0ntII83kuc8jLz3KsNOWH85
KboFUswgsUVCRrSm+3Wm5cEjBUSV6dt4y+ls8fkSzFqtVEXuUcom1c4diKaGcw9gKRlLZLVg3lBN
5q3nV1whqE4TA6IERqKOdrdcV7ic6su3XC69i88FL+iNxDsA+vDVmE4hA9Huitzf9Zry4i+xofJw
Rmo6eHnN/z5USwFnL8+JTOUhIvkdUbOPdbxGpl057aqdBJaxTILhDz3rPfL229Gmb9/H43DLTLa6
dAwfbSg+XZhb8Rvqq8IH5JuXOfLO+j5OmBqXvR8heXK3OyADQaojSs7Onkikqi0us58DI3TW0whB
QSudWFoof4TY+vXPKL237Vaz6z5mVmIwfLkWmDy12rIrIVKP+x8PgjVeQAxBagY05yNymoczDQyz
qU9qr6cc6h2zfuqMU1X7JcAXR5Nwr3bU0rnh0s13vTOwV82F8XsONK8y2voeAOQnxfpE2xRkNPIR
FwnzjoXhQyPCf57tmDGM6VkSfpI+6pu7cmCKlYGuCH/t8HogB/FPc+SNhsON9h84cIKjJMH5HVtw
vDKBtSxSSxZrNf4R/xyrpAS7YI/hK6z/7WfxBauVU8AyWWHYlK6yoczgO+bdHlblcFoikD8r1t0n
aA9ugIHq4dhXdQnxyZeUbAIml9jNg6l17s1x3AOXOeS9YN6ZBmD5rF9znyYwi3nYnTZ21Sv4v7Xi
Cf2XuX+0/6Tac0C1JrbXITDwgvf0GQ9J1PtiITlZlFyYLPy/gSGwjCij9LP4P543/RUCkBXFuU79
M8w67DIoO6XtMaWBe8RpeyV44lQ5IDJVKEc7Vu9dE8a+jbOw4x2gyYEz5XXAeVKbedZZxlcw8TFE
WvmhiNt7DvsgChDABmnlBU08RNfTqRR/rnZp15x9w94iK/F0hf1n2Ps4ayPozn2J8dZ6XLaHZOdU
7CX8bRgTQDhtFG5cZt7RbOFR+x6sSfYe2aZhixeksZLGifQ6IdXJx6K+Iu6ABZZh6S6aizFu3H0C
oY7frAG6gg3YX6BiXFCDOBkoS+JJrH8ppFtM9nUjrwktjwvupRASsGhxZdmzHHRmk/1DRtfPnhcY
r0ha/hlXU+2qYBx1pEmC5zHFEV1V56FiAsdQ3vBUAoOO+F7i4VEH0uGAUN78E7+6T45ZBhmRYS+B
F7SSJxWWMvMbWM00cxYMq1/FH6aUxiIZ8PafcM83dE4n4P7d2OBjh5XUlRHx7Wy6NfXV1DaQHXzg
dzVkf9YUj2wszHRgSF8zKaSMQBd+sxnr6NplOKu6iy+pUgglwjuQlupPmalBfplUvhJbHfRWtX9B
22du7hplSBW6MXV4u/XLXdF3RB4y//RYAVVBl9D++OlOrPVnflDQIfqBU2WM4aehWDAS7QiMBxKA
FluV7F8D3kQNsDXxlJPXvmRKVhKq99uEDU/W+fSdMVsSMuGV+gOILj8erfm0pnAiTfUhgm133DMU
Cpy8kAAaG9lpgcyUk0PwevRK2JhLVMPX8w6DlbvY30Fj7Xf7PRVGzKo6bDNV3h6ZqL+6DAqgux4T
zF6FAubA8kXP7IBOdZhiZJojxH9yofod1TmGZ7MxlVdvJW886TAcqAHfwRcMMGksp0SbxT1LcGth
9xGUz8rqu1krH2axFECdge+w1Ele203qFx1PRZ0rnAzmZ2P/tX2fzNsPJtOsCLTuyVgDzO1mqKMu
/tPveerVwG4zlh09BIFEWxVSR2pdmJ1FUC+1Ej7p5GLSl4iTHP2Qm9t7v8FLAhswZK1xntgMYJNV
FVl0y8uufZwOP7kHZ8CPb+whD6PggBb5ZbQZQ9FBci+8tw0E6fncXh4K90FLH1aL/kwPANAMYrvk
wmdiTPC8fXG5y45GSt86Z5CN99JAKTwHN4Ymtx7rZaVJLHXBoEF1rDYyKU860uN/FGiv3to0ZQdX
XXDlkvQn7iig+7Vcyvmdx3kHI7NqCbStd/txABl30R8iBgSBv5bA+/ofCxNpnOK2heXibZVvfHwl
71xh/0odUhbPmdtHqVqZEIL/ChEbZ/Eau6gLzeAVay6Zn3O7/8FyOdoBiS93SX2ninevG4TORFTg
WjiWOT/GcHaAvQfY6xXqkN5CwLitOy5jy9DlBMmFrEtbu4w6SG5KWJRz0gJzJH9Ylx0n0FsyJuzT
e4uD09pKuVjSu5tfv29hYraMsfiYqKe20DWMBT3ElASlxXDRwBQMFUPyqWCJ4f48LjQ8Z8/J59Mn
QMJkzsuowhuur96mFBYzRy6zHXH2jyZE8qcWrj7WCuoWLBG7XVZZZWhqqaoTNRu33OCjUw2oDVuJ
OHEBzVijskoEKdp56o3K6FiCabQf6Ok7O7avBgdVtm04wb6qfE5hgWhoi4DJjDF47bLiZdzf6NY7
Gr6GaSHWu0VlJfUDw/UO+ZqthmGIbDwMVEvFpFfgZ6GJ9ATQFkt0RM3LnOv7G5eSFIInlYQWxNuE
xIYUxh7ouzqT4j/bE5NLNhcBtesEWNJ1XzumlJs5sIQIyafGYUbzYjVdBk8Vt0jTUFvBPhx7brPj
cmSsWnbvRQj4tnHBP8CHF7lJ5ZeZ6y1iGGHwaSl/tY4eZHUmwxLvt/OeLNoSs2n+uHUPYv++rdq0
jN5AUMnhVAGIg8L0p5mb+Pm86K4o5NlfXY0dhA4oR/Lt/tLCnADBeHGa31ThWcel8vJOjdAbda0Z
gb+j/gDfHJ4P/o/OPb/8FFAj8PzvPg3CZ6+eqqPkvLn2cxtN0aMTXmEbTQwnlbakUDiDDeLID6mU
/9xeDazEvVl8kWtGxTFuqM+Vj1bJOGjAhyYEIXmh2j8y90oba0mci0gC1PJxy+OW5lsi7zddwfjp
2sEv9Jc4bVgFTvoGfGrHyCTxTfpZsslAYeujhsTQ/Pcuwtu47xyWYDAYz0fnLY4pTJ/pY5Cfq0As
BCf642kuvAK9NPCgiG5XXA7EMqNSCn87mzl0+9DGM2jJPKPHYW0qhgDT+pF1aWo8cGITM18qy3GB
pGVzgect2/Wgb4v0HYFWDF0w7+x4IRZutZK15JbBzDlN1Z9dTtpBbzFdezWlAKHypmcx5Nsnq2RC
Ap/+O4cceXcSk7y6oXP+TPltSBPjsTBvuAEQZ6YNp4tk2fSkmrHmdyW2FrI7y79l/iadiuZd2wPW
TiEN6QuzM54cyvlFJSC7WCubqg6mqUYJfrdbOIJea+sxVl/xodewaUl7rtLL1PhXk15zJApH3RiR
sgC9I+IzV/xgx1zrnIY7aoK4pOGlgF5Hf8Y0neGGj0EUQIEwvwubStLjv0lF9YHRtrTnkmlC+Voi
lyh6xWlI9O6+d0W3YF/B2G2Jq4SMmADUi5k5PtF20qAYo/JY88vvDdAhA6Mkdqj0Umwrlqsgw4eC
yDQfA7kh3qLnJC7+Fey1K96j56q15hH6We2lZd5Y91LLWwrjs9i0/yziId+A2h29+JAGRD0WDiN3
0pdUHP0KxYtAbZ9uLiKSHhu1ONIe3WA7+Ptm5JyYG25WscVKD/EsIvcyAonBlhHFrL4AE0Laz9v0
YG7AAynMhqDRF3yBe8IrOxgeIVcAAVclWbRmCKma9NW+5WyRjF7We6AMvdntTNb7XXgA6RQqARzO
42+/vvEc99jF+UgEPiXjN7w8fZpL7nIC4bA9LM4AZqU5BA6JIC4Nqx4sHquHvdzoBhrXuJ8lOO8o
kEHz9BYOONzLcEAOH7Jate3OaiHAMyzq1xIS/7rIWBSwvjAEE9Xv539irx7cTDjEZmgdI43GmyRL
TialcxgDC4XY9DJhtcuB4vcchztxFIa2NtIOh8SMBQKAlfEYgMa1WDbuK82uZ4ICpueU7gocxDyp
xMJmzCB4l5oywrJDF+oomSvRwR/nVqLNZZvut2zJbfu2GN6qe/EowVIrl5XPKmCvZCZDfqy9U44m
8pwcYsO8toSyUxEcMgI8s9QsXssnSZfzmWAk2io/uoDEIG4/kgeHn8Afgd/2VSfjqkFPvZmzT7Uz
Q04i1RyBE7v+iUrYm/AM76yjD3qZttw0WXIj7HyeCem2pNMoslVoK0LxSJmCwwbT6xj0DA2x0g/c
HImoDGbrfOI0lKI/bZhhLiGHIR96htfmYOA3NgVxx+/dNNuBlTw0xi7QYJbRzWYOvmPcPaCwb1Ds
0fdXCAbSV43f7N+6VQg9r3sAS63J7SPbnoswJQOzIggFz8cveET9sCUatPwfpRAptKJQGmhFz0kL
UwILWpKxZF2meh40FUNgXIX42ssBLwJ/NijK3zv7lZQLrjz5xXJPqK2IetTHuTC2lMASp7ZDtWvg
qTTl9MKuYYumqRXslDXKWGI+BPTUtldr9ejeweZuWAiBokXqfcLuBs80DF0xPuBUFa/M184L8K2F
4HzcJSY4eHQ02RFlnQ1DY7v5c7lVobK1mKlkTxmZpNgqdpbPLIFgZQLfiJ6xYpeOhbzggE7wsybM
/khV9uSO3A0KbqVgLiyxlpt/wmMvtzB0KeJNlSZRc99U3He7CTIwXLYc7I24/5374J5WMZbgsHn/
kCzuNfnlyxGI2396FHJ4n6Ei2gPBXpPFoyS4yx3qPjfN1gslna5G7cIluS1VoEWbCreOKwEJohLr
AKOI248+yYJx+SU6NjMixyuO3ogIY5mxiwrOkgXX16n/1FtiN52k5bJ4QZ+1D4rad0f9P1jxKMH2
Ba9YOZoIzLKy3vIGaNsF+2hFvN7UYV+053JhdZt7oGtrG0SkMEdP20UlcGg+Kg7jojjWuXIk5AQY
4+TZM9QoXMrtcbY8yH3OQrM/sdyTfQRy1wbbzhz4tcHKR+NWITGfKGUz1hUH17nCPehU6K/jFPU3
3RGSu/Am1y/KBL9A1mnYSa5L1/fAluMGU4c4V6IJFwIE7s98tqcECCgAm6KOo9+fsDJMAo67/OSF
hxb1vQUTxwfoEMJzcjWQBNjpHcAcFv763WAiOzj/UYHoETsQyDCFgovmdWfFBQaeXIL9aQDVrCAa
DajOE1Su5lWXmQlxcWc7QTShgmunrTsNU4LFbpV+uteIJPKC14E+RVQelWX6qpxk8S4Fd+XS+kV3
ONOznW16ZqJq0K529vcQ3n/CPtVURqKeuPNizuudKOlarKL5Xr2SpXm0wycfiANqSPqiSEsR+EJ5
cbPSEJsAnFXmxcIzl/kPdOZ/1sxJRxX2i+3/54stRK9P2PoNUtJaXoQyxwBIDoB0XB5hv1Zrb38L
rp0RRpbcQfG1JaIgFi/W9cjKMlEVH+BOwNtez+6hC89BAv5diEn6sweJp6SIyyjdHLU51HHYdt2g
GK9/2lorfCNZqvvk4Fzz3TqnwYNKVkhQzrfciZFemtmtAHYgK5VvGK+wWDK9aj0ek+n8pJ2UEu32
4xQLYP2dsJm5khFNurjpUoI/RLNcPeo6SK8hMRIRajb226yI1BiE8qLEZT8K0fOw4AN2xKBiJT1U
WvKnpuCXF5vM+vsdhLm2lQVR4flAQAOHPFp41pdhUEJGTvH8yo5+IpFGuKgcfENkjc/w9R1l3Qf4
/Jx4pU63jgn8CEabhR3L4iyQChets0bqbGebGywcsLp1cmTpJ19VGgvDUnlLoASQ7Nts/Tn8M6T9
ycJT2lbUuzKcr9tL1UBdIyoC42svWQ+DAeACbMnsnmDXJY+RKCpcZBqeQTD4EhC52HvRwHffLi6W
RZmS3nZbMZ9yKHJRmOMUYDtxbEQsSGQTzarg9ZZH4CVS3qM1b/3CDi+mZ+7tBi4PmeKl/DmWMbnd
cEmjoNYb+r0wcZg21GcCDDxOnUwbs2Ng4tLbanoC234Lm7l5Amft584OvpS2c02sLA2YlFnUttPZ
33yvRXzp+Y/Wt18JIeO0E6H9SE3TfPy5imDXcC3AraYA87yQhocPTICz/rVXkT6ebV6fCBFxjG36
ynIQLefeHdKg3zDH5gphvbAQPiEP+Vx763rhg2pLzCuFScbonZA3o/B9i5EhZaMQeGchFVDYe6C/
/Ui/P32YDOPNBq3Q6SQExABhWoTed47R59iPN/qe1M1MNFbbXMDGbPVxUOCBBj+zFNVgTrUpaiYL
iMVNtZbcl4PHnII77ov76V/1A74gAOtc2OedACxTB8k5BcKynZ469fydKU44lJDDr5awe21qYqQ9
g7uN5SwSDsosktnUEXknXzON+jl3q9EtkTCrPoxQig+pjtNUnGCROqvP2gjLRiC1kQVNyEb2GSUj
7g7OveDBNeJJvd3jz/SgWR938XgRmZbeqd3LbZJvG35p0hqk7bHItMDnxRXc2nQERXUTh0iSYHqO
qc2Ce3aubak8XBdqZD5nM09Y6Pwag7GYdrNFIN9AGYzeuT2chu/+QHd3NfvUDXkEIOUkGLKR6dgp
D15IhuB8uSHlfuWzsEkoCIGmNZ+PDqs5aSHKTQL3CbGRX3yZU4KgB/eElu6YcA7FhI+OVzRm+Qmr
YEfqKeaXu4Vj4P2nc6Ns+Vo6lQ1kZZlN1rxYVFMoOLnmqdR5Xyj0O5XJ2Dly19X29/zo6u/HOHvN
Z/KIRs1A7/YbWc1r0b6afFLdgJ6SfvpyHN0MY8wO5eC8EvtIPy1G/SRR4RVhyNdHSZLBERBFqcDl
fELfjUvVgoHDugjneF1GEXt+SRr3Od27HMszihg8j5tWghAkgDNfBlW/fTWyevZGvs9QDEVV+uoC
SZEK4GwvugFDkvd30HBSM0a3JsCLhdQwnBu0ImTKg35jHzfImBodneU6eTSQPtuquG1svkF432wN
dFwRIEPYgvQcVHAoWIUIBoFww18Es2iyHNOctUBTx18ZV4KxVeItJk9Ucxe+ZJRzqacQy8B6M8XT
BvCfFaSmBKnKod673aIu1gJiOrrO7J0cAoaC9t72o6BNCQr5krQWR9g+tOv+xO/sf65iuIzNI8L0
GnY6TI19DEtamGXnFyYu/14D4nXnF/HCjhjxJ+mppp6H59XScO3eZNLd/aBdO2aBhAiWHnbZJe5R
ihrIyjfp+WB14eEXObZjvWK6pY1+dkYDQ2p27ZXny43dzLABa+IMrfek2pgqJgTRxVzUBtiIq4JN
duQiYBQUyYmQmkudpzOEdros3DSfyk383RAmluPBCaoaFkuYDGJKTSmKMOL/GkwbpF/OOyNTmrFy
EO9n2LceEOTE5CJngg7Z1VJPrZ4N9Uo4yuoJNEILhy0coZuOxvT77AONwbaAb0GjsPcz4AIQrGuK
sMgddQaS95w4/foqVT6oT+XdwfZI+KL9/G00wHqYyzv/m/+0SlWlTzAlJO7HzGDTbmDn9o2VaTVk
Eiec+c4rZZ0ykdXmYPVfrmpBz2FwCh71AfUljyX8y60L3CDSADtMTybtj+D4c99UN3kq7d/1co+o
9/CMpGxWu/DzRrGf3s/JYpkRw+uYLr0GpCLKND3GyV7jwy2ujyesnGIM/uchfI3q5A17gD16CgQ1
KmmUVRKvlD06xCaiqgjzTxIGB+ByTRhQhnumeLmewigjPv3Bz/g7s7zNxcIhUOn1KhOlNURJ9WrV
xfpmyzt7E3NAICTMywAc32ghCDLpuH5yUdHWP+IBdMn+c//VNyfR5Wi9DHEMnowOP0N6nhxJFS7d
Yok40XFlhDH5AX1F6RD4iIa0YUqqVCE3LuLkU1uP49zO0Sijo9uw/S/SIITvoTI4IFo8BgcquJCL
/lOxL+nDv6lW3wWMcwxVMLeAEFkhu8Y53kaw8vofIcbXl4O/F7lGBxh95qzS0SiDgFZW3fI7VmgN
k8AwgK+5f2GJtAu5l8s9vftDsJyzoDnIoV0fL53yi50XWiKMTenhI/nrBlPtcLA1SSEHS+JdrUkk
TxixL8cgFJdKkXJILFBW963iHm5bAs2g+slSoMvzWFKul5kIgv2r8icrhjTM0co4AYf4nigz7YMd
jpio6q4UpwE9qxiLR9gjOOBxxrQylANAu3EeH0fOytgN35A7i/eEPO0jOoS7uYGWmcXar9NnabYx
q6LqCrBFpK16Hd7Ud0F0SyvWKfYLHEXUW2PeLizRXvKUagIemzbWZbAlUdHVewR67kHyDlxbEFdi
ls0cllOlmZgt6Kd9oU4T7KVSjVj7Pss2dLBiXCZRRBGcH8YEk6EgRsV0XS+sxkI2zFdxVNQaRmkS
uoHmpFT+YpoYfdlN4f5aG76nz30tE+YDlIlc7k/V94fDG//eBeaZzwXNIhZwGbzjiyF4VeT9gVQ2
wxWvkVF/E8eJ/jh4hVbfNwOcuab+eLaOC6zveWjzE6yM8DXUDmBrL4Z5DjJq1IDHkPMuleK7TUib
cQSOkNcWjBHbAymvN6mCjcug2Wqrah5ERT0o/D3SrPPsPuMFj9ZRF/OOuQNxholunup7vxTVGfAz
ZducDpWiFQoJkshfiN4+YWj7hgOqhYWVKffXt1h+dVIVgL8UU0Ggfi97Av+J32dhjjYzU9Qv1dA0
/dPEOorHO9/t9MQrfv46r4uBIBWgpm/fdc2cAWJ0qTCZSiFkgqU2IHAoHOJ0NUL9hbCxI4xPMbQy
IVWfVftS9ShhYAaXAHWxM5JCex+rxLOyHC1/SMpLjgOGfoyYHwbapImCGDEgVeCSiHrS0qZ6O8gH
lUpEnZI0NmzxnQyBusKiOrdBkp58plxAqvZM5SFNuKqT6wc2keGAXd55i6/teece6uBTxXygZfV4
VdbymbkNilMBA/4XhWuz8IB+r4aP3nEiw+/lbu2G0L+tezLvcSGFat1nL4wH2e3B9QeOAi6XhU4I
cwyxNerasj4oEYTCS6qTE+rlshlBLpCyl8sLQ1YckpjuCkEdJMGIyPmso6RZB8kVE+e7O9BaJgAC
INQ44HGhG2x/mJhA77sssAdd9JVzKntDavc9BgRyp3mEtNiuT79I/UBBcAPPO1ctu8RwSGRo7kVF
QnBPKAbR3bdcLXcGAKynS45C62QvghWiCjpNnyqaRAsASirg3lFJHhU8eJiOyGwELRMHES2WaHrX
rlBoRsaTW3t2o+VvvfNdmfWJdK4Jwt3obL2a4QjRrgqn8jb3eI5xUe8JkZyH/02+ro4/Szt1pcA5
UQxQe2n/IXyxABGqSsqJ0BgY52NxSgDw1hlwQ4BCujZZ/0AXIaLnJTQSW7BlBiESPOrj1gyyGtxO
LiE1/iT99HsHk5svq1Qjj0emEWAuEISG+Up+nDsOQDG1c8PbUNZKVkV/DgbzukJAHTxs/wXLNbQy
di1kwTzk8NyFESOClmMJFQvxsc51wV36h4aY+li0ZX4m/sG1jJjH25vVCYD6PkM0M1jsigMqEHm1
W6RGqi7b8mxO7LnKAZ90Z9XCnKEaTu5ut9CPbPbKghmfn9pw8JsSHZPlbi0+0mfg2PgDLioKMtWt
0sC8uxXRE55cGrWVyVOAssyTq4aV8Bx15g5re8DvFQ4qKcT8vjcFPS5gBK5TPjqy75PXaYQj3RZU
63vOjtupiNSiiVcpArc2uxdCaRiKDXHS0FcLAs8B1ZYS2IomxhTnJ9txIBAJg+eL8/9xSgC+WzKc
hVD2PseFZBEvls+bB9qhzwBbn/EofgMJqWLiNA+P1dJbOk6EhMXNgHJOrLs7jFmntmhG4ZP4lQQS
nANgJmYXvWIgGEER3yjP+WaRDLXh3YULzTfhm1fAMLtUUrWEOsyQsTzhIgayfjfQUQ+vqabDVFjn
uuqBaHPGrhF/Zd4WKD88LLZfX/L/1XFu9KZ/nMCJyiad3NjG6rF+2YmOomuPNN/xluDNS/yOeHdW
Z5Bfh0hvxvVlIugDSPvY0tSZesI0go1ZqEMDALwTKwisV52ZoLjeKv33oWminCPzo3j+ldWvhDWf
3nm4HwBI8YZYWNpL4XW0kVm99FGn68D1+Cipd0vjgdtuG0SI1yWGXYsLCac1e6/R0wmO+Qrajd7Z
4Qgxe+74YQ61Uq7LcdFaPjzV0leL9vEewVqe0FwUpJY5C/zD2sDvlj5hqRR0OLhfBJL40GVlX3PR
m0tGdVr9iMw3rfMYHimpKtt3RA+3t1z2UfbLe1Nuw6w2pal0VeCsEXM6mjClrRg9lTgKyex3OqZl
hN0Hw/set/jTzxdUGbtZb2ohBRe6Q44t6mxj04mqw/7bBOS76XmeyQKC6A/bzswxJ93QqarEjnPt
lbXxjTTAVMk5/Tnl4lgQwtAQZxfjDh9EcjSjlJqcQ2fKb24NI4UIxeGtvL9QdC3UYe9suFa6OPGO
KPwZubJExtMi4qpD75VmJe5kHn+oetgNkZgdSJRbPxj9pRbFuYH003buiS9RQZMeCSF+z3buGwfr
liiRHl1BFnBOBqYVF+pHHpO4BeUxZkPEdYmksdmpRpfKM2ZFX916pU9K2yKsXPHW6YbpzhHhXOpd
l8QgFqBsnH+oe/kO5Y5vIqaRKT8kPn/nxPo0TcATvIZdGZuH2od74iEDIC+jpGrqBebpeObSyq/z
V7uJlPDwbCKw/y36WiRxk1lDpy959owKXe1WNTB934clj94+HkwYgIBjjYFuO4Q19dyshv9tGCiz
Wvz1crSwYVIsWTE2i3Go6dO1PVk0eY2xPRaZy0oiojsB3oXfnNUC+o9oYWFhBh0F9EybmRJbrzno
VPvzV6PAkdESDGxnhfuVJQOjfWUh205zCj7/THjyHI2cY2M5XERJxqTY520WlfkLkH4kKPPvZdKq
QRp5n5fC9F3KznIZkklC6Vq3guAQAzBWAjpvi9kXO2fvMNSaesdwElq4d4BTe8OvR3fm2DgjdoZi
aWxK/CNkHgu5/MCBAfGND/p9+vQZF6N26idQSY6fqyGh5LtK6Qa9E0vBt99thJJAvv7n9BsLvNwS
os7Oc2YJqH6qlC04eCed5Oxa7D3MocM/BbiKH0rZeeaKpy/hxgx6QK2e86dOTbsyRd+KYEDRZ72b
yVXF9xscSk4XyIXl0SaszhWJCQRq621ZYeNZotO5R3Jfw4pgRPKG2RBeLbhUh1GBjdW1n+NSAZyq
3hMUd5jFBvQnn1OEVUA+kLyn1F9MKqhp1xKWP+7OR+25vgPe87Zx8zZ3BAv55XVJVq9634ScIUIJ
6TZfjdJq6edU4S9G40G30vvGASdKUFfBOQor7l7+lsuKY4NOIu1cEhEmmAjXgEEZThffXjHfRyGK
dMQOUbYbxKy83dT613VjxUGoF3McoPyg663NsfnJnDIpRBIdt/c0Ri8X0ThJJxnHUBPKyKr/odx0
+XKYyWJT6hl+YeLSvn5+2S5Z4p/jytJj11yu7DtwlkOoY3yuylMl4QFeV1g36/XabhXOfzUw+5dM
gurPUajupaZ3C9B+T6TBGnr0xmSXavaHUtDszPZfwD+eEYKGuid1F5yrfhGURgHmNkEN/45ZiKQ4
FFbz17LMRARJB6DLJj0i5/n4Od216hx8SoGVSguhxLsdwpEs8aTsg38mLnRlQu2ifAP209v0WHDe
bqPNlsKl8eHEJDSN+PaaHsVJr9sAYytxs10q8pTEwqf5bx+H2Ja//mVitaIAKQ6nO3a985sZEIiZ
yYCfgRusNhfbbKL4w7uyCX4KKBJgf6AdO6nHiqiszn/Ip7GEN+NW86YaKi7lLPBUOVFcwb/AtVVW
oECF2g4X+olrIyMR9QAs0b3uzMS8kE7Gg2wW4eyxoGLtHRmconxCjDjtOUVLF2odbvMXZ2Uwu2nA
W4FGEWqSwaizlCjVRWLVLlE+QSZUfWndC/Mqkxj4QAkpvCb33BjwdygPj/N52ZzollKunohNh/q4
KYjdAIhS/sAkrqjO8qJ9VvUhrV6p2rn9k8KzoTstOJbg/pSRfSxMfCfqopYeXL+7p2qJCmyGGSr0
/b3S3+PVxUbYeXswtufHmG6T03nNaErG6J53INOZ9meAMvmfhhOhKQ1ivsSmZ/W0kB+N81JhVxvq
muwJiTyUV6RzlRCv+ZAkNvvkLpAMd5UJ9ppkdz/Ny/mFg4RvJaFILscqbv+aYIHfp6rjssGouyP/
uQPAoHbsp7bdSsrZK0H74wL1vdhMr9BE4XmN0A65bfRSYwk2OktljXX6h/T82r9OqV4csvg4i0UU
tkcwQ4iT3d6LVKbs2LLaRx3nCNER33rqesX78a5v+bTsLJzwDzs46IU7ZkH8aUjY90PTSr214LDm
bXaESwItjxSIvdq40C+Zxltm470Dj4P6U5ftja6HHvXTymc6imUJJL26q25GpOzVdeSQ7Em3G1Y/
1EndqM7mFTtcDvhuBxkgZzixoG4jT4V6XfTEezRsGtGcNVZdceoEqytLLXLXiGpa7kbNwrbqdhQn
ceTFVPgNF9oOKJAv9AM6h6i+jBV5v/nR63KAhzUQxqw2PlYQKlYYAvEs6JMnkhkQjgZ84I/uEq/d
NMZIm8/3eIJoCttESRoM0ovhK+PQkprAw8QhiqhJdxYMsNRiT6DjCVEZYSFvJMpzONI1V1sufqqx
QUPkZc2ycLOliVNtFwiUhasPlqBZD+HqZWNhy1XlvEnD1xfgh59oej4ocK1k5dQggzOZC+vKnAQz
SOKVEu6JQfn2xL4fbP9e3hiBLGEg4703O8kDlGtp19xX/RjSvMqeuO/wv2jFiecRgfmR/F3q5jQt
jJqjlRVFnIm6Fd9cpCK6HwP6cGHbGETwFK+TNMI6pQCybPwB7kjoBDMwdHc8xQgavPWNVkx1X/1x
G7X3DDx20OQ2zNJlxEzEYrOZ+fq+zDgOR3Rw2hVhMEkP1ozhzHhus0T/F/HC6ffmddE35SfokjkF
RK2ullF+bwwW/LJ/Z5FFSBbupDV260l4VIkwDXCYHJ0c8VNGzVmdGudnYykqXWcz847Dk0bX7zFg
/8gyQ14Dx5kDmsXXhb9U6Emaety+HqJ0/2efMh34ybPlIj+AJb8zgdvblW7pDw/NvOZPiOggEzmM
aisbCDPWdEpHaQPk4XvW2szFeEY5IK0NHZ+QLAYrRz6fcXP5kfin3/VTI1nyMgxFiIMft4mpHKmy
vm5/4TSgoFY42+7+xZdhHjUFvcWyRwMHWUVyXEf5Rwb2Rv3422pjKWjlGsoiiLoZ8j+zDek+oGDs
S8SmqY+/PivMIwsinjRU+881mGDZ8bjUlO735wU6toizdCiKwNK4cyxc4aubOrefVQ3hLkgwZlF4
Q9+h2SBTH8kigSx/V4IYN4XMKG8IIrxvkK1Qp/XVcvS0npaGiOLZdSy8OEk//Ff1lG2TzdAO9tSq
uDn8Yqdlqmf2TH67X19oU04LgQauTKShqx2+aMLnPPJrXwDuFqFAtUm+L+6HuWnLKU6W7UvbuOvO
s4nHJt2wv18hNpcCID7rDkv5zMM612QwzFyEWt6WpzNI+ptr9v8LXnaI1l0L+7NFsGhZFmkyMiTN
mxqxKWgwiA5fGQbGAWAyKeKFVwBT4mewgo/H8obx3kPCezj8Dl79zw/jl1/CNeebcgzwWd68s7OW
BpRbdi5GxqSYfWIannN+s1j9nROes7Y5btjV4OF6eWM8/XbXF46afNE91EsR9hdCi+UgCYBm8pFN
HWagoigJVVXCdea8302Zp5uNduehaYBz1ahUZ3dqOUnl3EVHso3vaIwnAm/8GzG/wubsmwdW1OfN
7IG/DL2DJDFrbdlmBjG8ExbaeJSxZsnLTx71teQZo5LluUPDXg0DyB8HJMldAK9YNghtmtpFRfP1
PzjakNsUsQBowlN4f/NfGkZH2il0XFqfKnkF4MejfrFqS8oavx7aTUryvFfQQXFb3MKaCaFEeid3
aPG6Ty9YMubQRiVK21CMZxO27Ri7fKf+5RpFJpC3es2vXu/P8FlNMbNgG8zMKIPeTtaSnhQNlDM7
PVwR/Of8xGcNM5ZfFO5fmQEA2mT5bKobH8f5peJKlWTZjT5OjoKY4nhGsftXADAvE7LTEPbAW/yE
Y/gFY/mKcgZ71/96UN0nPElsPdl7T5orhCm5DqI4D7DDzEnSHOg9fMT3c7xGNpaINwLqH5htgALF
eUM/jdlDLzKgK9FyUh0cXL12xknUmoOSOb4gL1HvffCG8vbk6O9KeJHhhs67LbmWg9+6wU3nVHEG
gQnVwJRiHPVfNX79adoGXzhC3mX0FN/WTfZ0oo1JE36OSff5X7eExoIDCwHWoPb8+K3MZja8tz7+
zEH/XBoKBx9jy+jxFtVIBS5yNZbLslgswOo6cc8e8jYchSF/3fW3bEYCvEFrDJe5wGUAx1qNCXyz
KFSfWoCuOa+jm8wNNKvkHw5B8YUko7/UY8iEf6tp3ve11dHrUlphWVZOvksz0Kib6ZHGHdg9WdkD
GUvFjMJv8V0PUmnvBZLwCS+9bCCyUW+P+43g70h+ZiOgBbGFY6eybGC4rGrEp9gGruynqIH5Po6I
GBtWmKGGVnhY6/buimM0dk1PpE4vSm3Y1ITTx66frSBODg1xE4uddIRgD70G80ueX3NYwnzYBDNv
UDNf87ac3o0RzN1LNgqvqjF2Zn5W0kYlOhQHUzWydIqlPgfPzNfnvqjkumiZgTlvNZaOeXFeZ1z3
/Jfn5P+JifoQ3mYXhSQevpL3DopTcB6cV+ceRnTE9P1hUhLhxmciBGvu1u0ajKJG4WXoqvk5i8Wx
nARhayQ3q3AW9C9eCeRsF667s38a5oGlV7wK/2STIY7IB5Faqers0grDee7h5E5OIzsE6NIUkLMx
RKpHawJJHuRd7MynH0CTp1tYhsB0/fqmkEiEgFX6ViGI0/WzMwB5Zh6wZkNiYXVMe2h6EvUvjZGm
nfYr0fTN7DGjhpmLTTGgo4w/E4hOE7j4CJdjr0k4h5wjs+baylrfdNpJmnl7YULwbdXAgBZiAOVG
mH2HORDMGD2eo5kTWddjbkCrE+0YSI4xO7DZkHe8HCuTOrV7crb11BOl1kB0Rom1GmtjvCVfwkJ1
eUEhW1Sqo9UGFF0R+c7oZ/0oz0bDA/WVBrc0znIhvcfxPCoFKDwSnEyFO6dD6tvirbS84e/y0oGT
kErXDoBQ0hiFrfQlS6+QJ6xdAZjnAPt7UQy5BL65fLkitKafibzWdyBThneQvr+8kvRzUmJDqUyE
BVeRV9JuPiYjTLxlSnXfGVwbWA8BuSp1qufzCHRVA6BaZFCZGxCAgOUNpph3ZfHkCoNPfhLmaqDV
ll8MWcNnYQqyQ/qHfBsQb5bnDEEwzfmj/PXeTkO+u0HjvQWb1nY0TtzKCo0pI9bV5LHzRTVHnXXQ
3qpPHyiHUYUrBZ1BkyzDNhDaMybnep9ew5d5i8sF2P1eTUM+K4Ghg4LnEXryLTsxNfN0g5NksIml
oaRjCQtT5CId0Jjj9h2Z0k0Dkgu1DStze1td1508sOiuB13L1//yUIj6FMh5Ob/98fQSGwXCaJIQ
RJWbxHErHWuoifjyVsOHXBmDzyzAwEALEwckcU6Vxn59L85FE5UoOkqs7APXS8BUc1arSfWxhfqg
J5LU5Uwkc77GkuRGDXyG635/YKqSWB4fz7ec4E/aMIQjWiOtzsONaxZyeIEyzQW+6i2TAEEHGeiF
1LOhIu/vEBmTIf3vOfq8vkFOeWGaxUjylzUbkm2YxP3sQBuTxJup+HuO5MQiPjQhCSLiHt/vI5H1
gdZXuLpLjlUnmn9A676LsuHAgpJ+gaOSL3mJRWTs88k/olOayETSzM0ohoWva1IBSiKywnLsMQvY
jJ9IFO+Ua/OojdrLX5UWNCbJpM3yjX91X2gizHwQIj7OXiV1ZVKUe7rAIZlXsDCnG1PrEG+/XJon
9wzS/OCDN0VCHRtDgrfO1pCe6ja+y1zjcHDXw60HUSwII8auyL/uV/8033uimJqOGOVxu21hQzHs
YywpAQ0fK0w+lFqWLns4wVN2IRInoMhyP+ntFNo8oTFta6h8+1ZmpBGhI+3sqrVFWKcMQbkpAhyX
P7/6hJu4T9ycPsMJ8M23vlmPqIBbhRkbs0dYKfLGv3enTS3RhovuPhhjqG0ymZ1Mo6DHwavsvFts
6QThTmiBBPaneONTqCeCLtLEVKP1qhmcmW/yRl1R4AehfEuknXz/yIraPQU+V2FTbeJs8UPMzEiv
/+PckdqOdWN3k+R5qaWPQQ6sbSSd74XsOua7YR7J8oFr58nJ2igaYYVG7+sqbbKYLA3Ux1Qlur9Z
UMLmJ/onCtBrOzprT1QeWmiy3/dT7LQcC75xPP1jr8D16Xn/uExZvbuTuyXKY19gz/lyqk2+JRU7
RJAlt4FLDYQ2fO5zILZSB06aKpHe/CGKOJwXzt4AsGvviSNVl18icQJCL6KxQOEQUB7pOJqiCv+c
I8pOdpyIvvSzRV9IhDTE1NIg0dqvyzGRD20gNEeyoU5SM4nRxFgC0+8iWZwaitb/W+gNlHsGu8w7
P2i0zcS3wiQ/AO5JO/4WET4XfpjiDDPgisx89z/B1wWAWacFqkLHiXzz8ubgc4m3YjXjdD80flEU
BeSN+wDMPa5rQ9/FQ4UJUrGG9WRGcgrY45tqo963xk4gBKNqadmsM5MjceWTbFrpV3TK/9dyW0cA
MlN099dGgriIPJOVKnpr0RwqHZKLzHnO8aPxZnBJHLiEqnREsqcJK4NhsEmlkwMa3/ljNsBvyVbv
5IQrFZnFj9JJi502FHItwqjm4uqJsDeMtTKxBOzlTPvxU5eiuLPYR6ItWd1trnxtbpoduSDvoI3d
ywxu9rsML8YApjVQ3u+gIUJYf4k7yTZTBK3ocafC6/RAViGs/D4MdkbyzyXwJhb2qw9pJDyRcZQ5
mjmoWvAFXHlMTm3nrqy1UT5Jn2nj7Kij+A8D4F4qMWfJ0xkp+VN6pZL430f44UjQLG7K8GYPH/lY
W/bawWCi0b2MVRZGuBdBcsu6OeVZJpmsjgUclT6DTZZ/gw5qCbbC4CXfhPq5+/XHNTtybAliu0PD
lpBf0I/iGyjl7vtyghuQ4QaDHoNUPygs5bU4HtM6PwV85mfNgspo+N+z4HKyRKJGYYTlwHB9f0d8
SlVa94My7v+DOqTa2PKQIX0E12ke3Dof+8NArAionCSPPuQJvrPKu0FxFyvChC2tzsWgByG70R9l
x+2hdmU+khLMEVfKuem4iRUtOuHwN/n90rq8v/J25P5auFZ7lPUri5g4WUwNTUe59/uu5762i5W+
3ZwssgrMKhBDlC+6NZR2fQ0Ux395LDWULVKRF4fhdY+QStOomHbUne08zK5ia1Aj03bE7hjM5KxB
lpjraN/OngQzCJl3HCwNT3AsbmC9fsBybJ/etKdEczHm7cOWnNShwMX5hOz+HBe3LVq1cFRMJFII
DCEyxxQ1u8qEwfXNFYtEW9vMDnsdBbn2AKIB2tQOIlqiPv37y32ZrGRQatCgVm7TMZjBJ75cG6qU
iMTPX2IaQiQdyAVirPArmj9h2VBiOcLWLPXOo+TzFnyWHPa3eMXA+4Ho7NSBOPDm+WqxQPSrA/ke
lNsBNlyFnhIdU2jgOh77KCUJTrqgO3D5cZ6RYzwWcXjJArw3nI+4MTQLvFbBEMFE/Bh6hkkqVZVz
SH9VZ+a7ghRBGHaezGklluFqjNkguvNRd3n/G5NKRt0dOZfhMTBkjCtR7V72Ro9uXj9bI6f6EzdR
HsE8HE4+89Y2JdGcjy67fGkQw+Om4aNFGAz5yGkCsuGRttcu62uGp8MebwXK/c09d2kllM3Rcpg5
ByLjwrNBR66V5NDQ5GnuutW1hJXbldhBkAWnjgvSNU9LGU9D951jJEVuYQpC86p/c/ZHtEHijImu
74MvB76G+CvOADm4mXbWuLhqEz6ATrjQjBYkKJRVPZEHzdihv4K9mdq29gW5+S9niw6I2mbKErBt
wgALX8W4d0859iRptWcIgTlqZ5yjJ0lIPcOVvwyO5roZaKMIJYMVybw3YBIiwfEaOZ2baTHNCzGf
jwyQMIMjy1zPi0v7X3A/v+PWppu9K/EF64iTg83mcW+izvfNgLtSdhjJ00b//u4+X8rRkmT0UbIw
sqQ+CtJKs5fRQ4sdFaDI8xZYO3JEU7/q0LEaKDv6tvAHJhCbe9KU2iQovsG5+Qs5GU2LIki3TWrS
QBO8Bq04WqElcqg/LMVvmFZuAi9LlU10U+XNYx7jpmlSLAdoIoQD09TTAocT+D8+LxtufV7ZhTgm
OBw1ZSuP2N+3YOgkG0qEYEJGZh+THSA19JLYdfr5XGl4wD0/gX7OaqdJ7XInkhdpj6TZLjQ4FyLz
QVPyyeWY9XVzwiW43nEdYcB3z6F5dygqsD45z5kP4TJ3exzpgycbgvTTbRACUAfVgwJXN/yYZ0hD
vpN2yGKBY4XJ+pWRQE8OJ+8KgpXUNCyR5OZQhako0EZ7MRYLyUb6uJbX4szQoI1M8Em5HNDFIFr1
9BJZ5t97T9sjyUZ5Yrk8U8Xp6Lnic0gCwBL+5EXR6cyCPddAmI9Y27ZzrNe4ofrcuxDXMdMK60iD
Qdh5EjWEFyIWcPaATmbPZ6vmjzgLFP1GxHvJm9LXos4pM3WP3Va1K+T7A7se4za1irwiOIvIQuLB
s3/2jKOEQ8eahPY+huWCrd2KUoDLkUPUMBedjTvpE3MsEKGcilTETR6fnlQ92TvtiOvxuL7+YXYL
juDj/YdeVzQ6ekFbQigWJx/s5hS5cuEPd8yBk9VZKnslB1GtembI2XceyBLt86ojd3PS2koEYgCf
lapirJWe80NSZImiXgVsWmzjH/z1QScZFsBlGGqECytdz57e/KGGhSeW0zOo/WKDMQt5DymXUlLX
P2dJTttr0gTLlr5S34cNMK0T53ozBzVIb/fB8TXgabZV4Ti+iODN71woZfMSLK8oEI13zj3MkLly
oeehGJO321FtbfjniUw+Ux7mrJb1OjZZDIFCvbwxHCwzySJgCXRoYbO+vdxNBQ4dDFqQ/ltJ16Cd
S7wYHTon5kGkWhM+Zp6cbW7ufacWUwN+K8xhjtQmh/Mp/WiYIdq4Ih7k5JKhISuPjlICuvZCsc/b
YFmQsh1hKjRRPZFlQ3YWPEkdfiRH4O2EuidK70KnSMTm39bhZa3NPTFwkL8B0CfTvtQrEZyf7O7y
4OIfscok6RbOx2T+Q/N7UFB/6PMAOLxC9cPBNRn2LIEepPueG/mQW3hXSPUdNzCJoMbETF4TpaXM
6+k3/V2P5SSyntV92wBKwNPGmieTLhxuoiTHR1H6zVj5yg0XdcakMqngasovkM5/vHA5tj+Km7XT
zhr/6+5PfP7sfxwpRLqn+DKi7QACwUymGHGVgO7SuzA3SBLfaLyNUFAb6cD1hGK8c3eaRIZ4MMKr
45RwI+AG5r0jI+yjcKvjrXPGqB7DqvhgSin537y3TphqCdkO+bnvJO7M/DsdH8vqbnnLNiCZ6nYS
gKgnbf2591wbaPQizxm8ptphfFZgnO7+xGPdDxG/wfyUugAlaVffoMLc+4giOTG3kgqDrtFoPFLq
hz7CXwaY2Y29A03Lw34CNbyJLtsYHnGx4DWGeEdtR40jpEyYb4ZANGWYJA2M4opAtk05sIwlR7nO
60PHixIAmKmgNTQHkuqtpeycCu5ndBiUYqnHY3agVaosLNYGS3UT42vXe0R2Xn15ObZRrjp4o2wE
yAqgRl8wDOSYVJfP79SYPW4ez/soiHe3WOXAE0qFZyx46oVAZczIZLMKPrtgyhiR5P577SW4f6cd
d7WMBYGwM7bdIruhf8TI7jlh8XP9dADuEAyHdCiaVzdr8ybn/E9HnjbLCIn4a+KNbLFMQZXcDVxP
wlOAs5sphsMNG88btPj6yom/vxurrCZ1+dSmNj6/sptYfxJBr/V0XEO3M68S/OgtF+rqCcoAXUxv
tM9ank0hw3u6tR43Wl+ac6qWa4tQyp2jn5po6leLY34Oko1Wc9ypOSY4kLxIkwskk2PO1BLjgbLp
NIIWSF5lnaF1IJQg2vtzuInVrlYbsQeZZPqnlwEmLmL5H+psbMxFbQDFxslEJJcSViJk7PfZOrvk
ARaBe2DAUOejIH1XpWZI3h7rGEcDvo6BOttk1xUwe0lXr3AQcVj8CsNAmuZqoyblvT0xmiLqzxVu
Vq7LYjggomxkNDNWkcv0zqpMSP6S1dHZo6Lsgw04zcpytTenzhXB926AJ8VKGRyfvGX1ARVbwKnJ
iJR2ivmBGA+291fiCf1FqDNHPSrTYG9QAiXzanuyd4nZCjg3+LEpZvMmpnDgsa9wYHya25mzim2w
GFSeK7DFgTQWXZpR9rtjhjypf/dPpdkjzuPvewL1XPsUH0ZvGd2GXV5dRimET9kog9E/Ob1W8HQv
qsMnaVWLcPeEtBvQBQ6Q9VrHbrVnBLvx1SNpqNiLUUkCNeSf7dy2PwZudjJJuuIWQxQUrpcC8znt
CUZzm2lcL2xJW7iCHj61kfO8AcRSNKsUcNFgLa1UIGPr/nexOBbqXr+nA3M2aIgNc0dYN41UZBpM
JH04Rfdb9KzNoSaAwo3Fv9VFzXxAjYVC0ZYjQPF7G2ToCLz2hMHdTx6L98xwlvqW9Rq48QAAap7F
DP3PaQa4vqtE/wJw1HYM3elUvCRZR73er+pAnwVhgQIUvd5DO9sCjPL/RkyqPvnJduLN4dzQSbPx
nGGWRXhkgbLJlDOjyZgsQCVpRolNGqRF+vIzEFH4l2mzXg0C5B2txQpdxSjQ8YiSoCbrg3F2npNE
UDeyvc2hw/2hgFeAE0zZWrbdCeqUjuTvqwxSVE3M9KD7wF1k/rN2kcs7ZsGbU+ONHFUEhOqFtEpa
f4eVoxkW1j9q44M/DxNZK4FdjxyPpMb08FasCWL2thW1TPuRN6Be78lsSd4ldZWK9TyLQLv+DlAs
6w4g+DdD4FCxiUWa0YgQxcWFsN4QjSuDh+ERgXL8bVnVere1++zD2RAG9B0y71PUczmISNqmVbHS
P2bH9rWp5yVt2ITS6ZmzcZG3RIOdMWuvd9WyKK1yplwhZ8gFibDkNngBRkiZD+p8W1se5tDcs2uL
ge0729RmzxIttR2SoeqoWlq5b9Rg7Il6w7JaXRzvz1HkiQu+z9qWraQAUtt/mMji0bbfzu+DQwzK
L+7q0PUeJiiI/r7hsxmvznAym9bsFKqJY8o4hpJCPAM/b4UyL3Bq85a8Ng6BdPhTCc7En0DZkiLt
9NUmiUTsJyI53kR0/rv3W/6Ko2ClblFvdc/r8lRPwKsgu18/7vBL2URn2asnaocZwQXRguUrY7N3
cR4f69TN1NkGIz0qDQ2rgMOF4FVTI1OPBdHkK/q68J/jL5Trh/+kR8oETVPR7gWM9a9H+tK9zCmI
OzBc/PvgZRVZ7MMU/Mgbrz17DX0YuxPx8hOxiM6jJvIHdWiP1nsYti9OsS2gTyuNeAKGLQhjjCB7
WLuRcARLtIQu98mmitce/5V+CbSUFNtdrrW/Hr8K1Ydof6AY6xxABZkY0jvDnds92u4eHaqv3TS9
ZoDPrILESBYMdWFYHnfIsKAyPyeMTHhMkCeqL3ALdSBlRGkt0MakZQkx1fbFCLHGZ7nIQiH5t4iX
iGSEKT6oiUjMlr1sN/R8yTKtdceRiF01v7p6r3RUpoXEsdfVBAyjtJcrxpVLGZm2wSTbM9hp9+cY
OwFfTujj+Qm1W+YHZrNAWzmeW4gDsGHJ2dncafkeSlsSo6PpJljkbOJ63yjxn4T2Jy9p2M7J9JE+
nxE9ECrqfgnhaRh8CUUET6M+sZeZCd2q5ryGY802R5H8IkhTpPoolmCvLZZZVw/iQ2j3+A1J/1Hv
3qmxlrWa9XuqX++pIQKjGkQBCK7p3SOVnma4WdZLezpprr5Rcv+8OLGgSymsW6TSdLQ7nBI8ginx
wQcsvm2xuV+/XXVVunpeU3wR9mEQeN01OSOehVnO73XzaiIjo2oBhvqW96ePC9k6TYaXYdhkeCEh
nwJ8qxIkbdn/XryrqQHt/h7sBedBZBDX1PFgXxvDO5Q2wsHSCtAMb6pYU7hH4JKCj7iItLkbvV8r
pyAlGq2iJi9CwVbmkCgJQ4XP3Aqbc++0+ia3WynQGS4B7FcBIUiOfVWgPQDx1NI4SHciZju7eAU5
bQ6JXkiu8RuM6EP1OBz/8AmBdYBDilrqXPH86YSYy23J37CI68XlYLnrTbPhh39gi34/Hy3MX5RG
b9QzIHI2DgNP75As3XDehvkdD7ePcMieifz5DOo61FrGbdz8g58pTk9OxNBm8s33OzZyAd7Z8/xF
cX7+JyVa3ruy+E3gHm5SsZZVzdXj47IrawRan6JwJV6NLooqmUuSbCMAHXFJIWd15XTcCsDnztAE
0M9KCpb+PqxYI2tox+iK9zJujMAmGp92eGKH47XiXLCOzhKW72ldkHolreGoIHIE85GKmvKt2Utj
FhYPIx5KZDmUFeXIxUPhm2TYxBgo+qBqIlcKABRXXMrSbF8HIetVgRDBZGCVqe+YtZwwk3nlwmDX
t89A/MIgQfvJ4zJ4/UQTxgbqrbqhLze1YSR78XQ1JvzMeJ8eT8jyPHWhQxfcLPXyrBm3SbMyEjSv
pdDcR17piAyQW8yIDWDBYTFVPvRNA/AfoDL4TwgGu9iUb2wSd8tE0KRDAvcPBjXardmGv6P3BtMz
UAOOEVqdOdheLsFz1CbsboR30YBxO6cpvTJaCDGuccKrJdSrSMGqBKe1ciHzM09Blo/ChBltlFn4
O7uN/uT6P5U=
`pragma protect end_protected
