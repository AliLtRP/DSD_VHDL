// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g279JlsyHELGmtXY2JysM31KUSFND2CQKJ/GSq7UqrGhPyUExK2Px36giyPJ7ZKY
aeM98H7rPH+WC5PAB1+Txnkp5O7OTyn8No835XRotOPmIacODzHT+zoXgkxtwRW5
AuoLm3Dzj6leegRXnPeiRbA5ohC2yaWfF+kOSijsmGI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7760)
pr9bqVbq9TwTgJGWwyDTPXY0PlCDqsvCaVAV2Rxjujvjh03yeCfPn1BdKoPJzbaf
/SfdJ1bTgX59h/LuQcuiyOXTwpQaBMWDvaNSAu0Rp0tfS9kehW2bt/7LqZvShdx8
XoFTK3AU/BiAIuL0wbS8yI0qcfuugSloStOS7U5ny9xrUN73+WmEm0IEO2WWmJ04
D90i9O26ueCXRbISdMQjldNcdekGqruC8u1kuJQ5DFjTowQdSWEMRqbo2m9DYn35
YvV8N2T6vpSnrQWyDQHBZsKIrMrL3xjl9N/aRl7w0lKkxsYlr29HbLXiHL1q0wgD
Z6Gv2YXA2q2OZ7I+n5qtRjTI/daH20GuX4T5T+86tOvqxeq/zszpCkbjzxw6DObw
GF5dIGHHP59PBwTczhkubCdBwMXLGSpFt0+0ZBV+tzzLiKRnRa1d358bwnGk/3FX
iOi096n7cKD4ezqP/X/UJrAhKZogidO+EqJq2AIw/b/oJPMdUy9i1R3Jcgs6eDRV
EXLHPgaLyshTzfWnHedvpTMR+ue0teJPovYPTBhe2/1s74BiEuiEIECS9XLHkYYU
fh19oldC7BSVd2fdkbPBKGcHpw2xQ5iUwdHdeWLNGtRnfGe3Mh4W42jrFvzj6aeb
Us5KwE0y01kFOQM/kXHGaPKie1PnVxYvxZkH7ivjvcO3xstCy++OO+ISPtqaYtJF
3KwTWYvrDmIlBSY5KiPHAKYg+ap3PaXNeY8GlcR2xbnWydZpMdeO7Fbx7d4J0ulv
hP+mevQugmMQbyqsdVnAp+dk7hI3sAQz9chnxjJHwEtWBVBWuQfu65zMGkAPg+/k
fGQG6+fOEZyk1Rx9K1JsS9d1IHjljNqMIUE4v452xT8ghGo+ttlgJ30k150JAmuU
f/bFKYfnXV9fAiDAXPSx6g6vykmgFWfEWUEyILWEM7TD3nfQ+lfBmYJI3P5VsSpw
Or4H1rbPbE3cbg4G7GEQoe/AF9i/5b8NJ9cuQHrys4W53iUmq0sUTTF+eyzXrEMw
7CzyWd4t+v5s7hc7YGdE9mp8NFz5GDQj4iBHqJrv7J3ej8C1pEDNXSCF8+Hfrhur
EIRKt38p37kgfJR5MhZWFKBKPLEVXRygZY6sZds0uQO4GTP+4EvOPSQ2Gyv4NKQH
uuUZ4e9JC2mjBTggiMeu9U5esJ4sVPu6pTJ83yD1ETQgv13uSTqPxZUCS3Hmw4lC
20ngUPE4AMfWKd6wy1ExEhxfxIbOpmDBl2DbUB4Q5loQ3M8ZPX7dJxNFJkTiPa2R
OraycvjfDCuLzgoq52Yd325rqmfXtA74UCoyVvQ1UvNe/Fm0rj1SkZIsWa+RPnTb
IYu5iqjbRiGLRCvQldshTalbhseM8TPORgqhpqmaO0EQEAfjOizMBhK4P5ExYy4G
2SxshgrI4UD4bxXFf20RwVP/459hw4/arBblrMmrzZF3oZAu60trAAzIwcfoE15g
qDtlrA21t82oLStqCRKr8WQCdPCeKeGNV7jmTK1ksG2xssB0uVO6LoThlnkxdkrP
M0DBc8YoK5ko4oJOLrrTVeAnj67bf7ymfevzri5mdKvdwg1W5xo0cnoQZdVEa5+0
dFQnY5iqEw90KrZply4E9oAFugYoVmkOS9iWBQt4LLzBu6z6mQoo8rJcjVvnssMS
AIipiCubxy/h1TrrqfKJxU3mr9mzMQf7iD1a/aOKEEKX+L2G8kcvuz+saCKivVq+
KRRLVaWmvYJwJuoqLr+HkOUyOdSUl68b1S8ehsgzpl26mSkUeW4Z5lsYKa9zOHWG
4pGzoCCOB/xnnxqqitPuOBVP+wDZtXEvt0uyCmk89veEzL4KHBImRet9vxppQ90Y
t0qpm02Egg/qnY86PQuhetUfCe2GIyezzeskhdkXjNpb0SomFeXqieABNJizOfeb
pi/GOiOffpVL5kv5Aqujd7K3zMChdi0RRVfTm/5dngFixDY9NkzbVp9/HCer3oE7
jakt0WNWsTvZWEOq+UaESM0gPEKKCp2Nv/12E79bUwUl/7MwOlKfF53FaLpagGuT
2p5o2bv2uqGJfPU3JZOC2epsGPI5M5BXwqWvhc3gcH3u8UOVy3nlA9sOclehgsoP
ecDCptxe9nB85/MT7b/+NddrMgXSWjWjG45Mj8WDt6BY7hq1tht26bAAHwfbWvX3
lXPflfbOE6+tL3pteQSShVY9SWiYbj0T1WnnWV3obej0znMC1R9DiAQ+ODQt5TRO
lck6+wIwZpsKeQMBRHUFJTdw362Si7fwoKHDYlGG/yBfwhUynZwwVeW99YSSfXcn
woJJ3+iOAG9s94SJdwa9fZp3CYwvN/7v8sY5g3wk26nDpsn4OpQ76A/EMPOjFz2K
HJNv+Nib8zQASNdzheYTOaxNQRUYPRyTML47UGS60rTL7q6Vd3dFxRJumvw8CApo
4HKmnmFlIt7CYuSng0KxC6YmiAl1IB9XPe5kmu5G325mtjW0ZpahSo6aAraTqiQt
s1EnZK0QkZIdsR+gRDDJhbVL02/A0kyTsqqEC7WsKFomAM6LpGXZqRdNtPIjRoYq
mThLlTROdRJmBfB0y4ajGzm30Yk1Ru37JClyhmvRcI6NDh9rsKE0bxNOOW4z0YJ7
W1inoARPF1/Uwrp/C4ReeC2KNt6zqc7pVGOj7dnDmH7DiPvrJFozFeiccYKX55XQ
+P/xZHfDq0piZcmOS3HEfoJLzJxJ9ZIMV6XoowXzKSGzbVvljPG0EvY6yzUUuH65
fTr6SHEbsZQWu5YdPuRvBCl4fqRBs0YfBZCNAoVpXNjW2G/DH/xg2eC9DECmfZpD
j/YbCjjX3wWqLvZyG7Jw7oRtU1SSHpwkqxjveuP3oW/MU/zeGb2GH1IgYZXKBH1Y
9RR32l1LeCAxfY6cBhDRF31vnu7ib7s+JCf7Zo5ckB6baqZa6UA7c19q/Kv6uG3c
7t189xyXas0m5qrDiMUxxImSqTWVX0+/6APqXRaFwPerQoQ0KvAPpRPUTOzQOHWG
5QpPYO6trECpA/VmK8mOOe3NtU12kLmTQstDHu8Fkk3QfSoyfHm+XuijYIBcgqFE
mG5oaeaMqE0NYVQmW3PLuoOcN9GSMV0nMJxrNJZN2Km9H+yTR2yzmelJt7bmwwCa
V8XMHWPHXnmVoOjviULJOFrj8vhhMHTdhLoA646+x7U/XWj9GSNVCg+6bPOK4KqD
hyf9XhmbYsjppVwY/L+1vBvizOPqSbb1+ADiCIFfvCHnNSFeG4RqwG26OakUxx8S
CwkFkyUD5qfBvS0n1OaQ6avl8h63jyI+IRL3i8bp6/CJGcB4EVHhTpuLm305Chic
qTJJx/UKitw+Xl9ZuK7J7LrT043mmR7qYap56haRQN3zXNWWw7EOJ42q52Wss9Lo
IggJrTf7uu6u96Uok4LRvRZBjqL1KoqSPwZxfABEJbUj7viJbPTeyTSr9QoiaX/C
6eWpAYXD6t2OgEOo08IgiQ3VBV4GjkUMxvFNowdJurWYFvbZTO4t1t+qel18trRb
lKuBdFHzZHHJAnZcN4N1e194wUTHiH15adKYR37ByTn1/Pgh/IWu83N+5VgHdWRT
veIlMBg4JJdCxGogGiSjQIgCCVtUSOay4MEF1YFlZkUbokh+eszL86IdO0HQrGkB
QNO+ThWHHVsmSAYi/lD2cKVtF6JEH4ATNBm6XZRDdXv51iV6Xc1hQpkl102njurP
/HbsS6gkWq3J5t0+yR0omYWVvJ+DDfbJLAQqDDVKTEkbb8IFPxXfjBTvIIYrgbIU
oJpw3pLBg769QSNQ093c77FO0hDXkMoy5gtF9AHLzKkfc6lFw9LIuC3e4+nNwBhd
DTeK+iqE1ceFM//Jxvqa1g90mcPqoSSSxN8m1cD9mSKoWzWbUhtcXFQc09EbukO5
qqMiYVEL/k3K79NPiUAZSnBrsSIOR6UXiahzmVCZ0ZMWgq0anm1fZHz9OgplZU+9
eJ8JElKIAK/ljUgbqWvXRD7TH092GWHKKdxd7dC+UrD3zxxa464+dn9WoEdRfNmQ
aFcXpL8ArtiVzXEm+l8ZsuUkUihB5PiSappB6J1T+4Y8zvDzUFQ2JPCqxAEsFEt9
QVlLr9aYNsIueST/CitZ5yzmRw4VAu11XtDHBxa93WBB6b0C3rmfHtEtC4+wI2Km
fZ+hPN07aAk8SU3KSPpTtVbSsEnON+HLcxvQ1tbgdbdOf4wRq6ZMH8hl9hUVPsrG
VVeKfzuBKY28CKJf6YmOSa5YBwt+owqocgl1iscCM7yifM9K99/llZalVhs2caxk
ZogohICG8+3y+jwBg4l8frt1OpjX+m3dnShXwpD+IFSrnQACL7doVf9guxNnPfvl
XHdHUoZsHp6xGUMt+ju53lSmeLMNQfIkYES1bKAuwEgn5RtQ8s5bUwYKfFs6fqvC
M7vAnIudKciVgjcmhEhCHenee4US2l34GX0izFHcr9tfguBdgTaWG0OG+MnKz5Qq
DaVowX0hCFdGepbdCL6AONANZXS+fO1ZJnu6fGrs1GphaFdwX+TjcgrqQOzRqYmf
iw1JI1xzWtrC3YIPy2mmJXS2G/DwvhH62KhdiQiJ24I45uSinnb/7Sko1JLPWMLZ
xoCxZX0tP+ANJtocAmEicZj4FQnuXDl619G+R3plfG8MP8zkgdvuFbWnSPAezFF9
P/qPLsRUlgnlEwdypS3gX4dBOic9Um+h+VPlSTFkpiXLF4Hl6FskyOu6r3wi7uVQ
JRc7E6jtG8y7u21zLsrPJNLaa6yJQFK7Vh6IjGG4v83xpslUXb9S0a70aoS5puWR
P6ceqtwJ0J3R7e+L8tvkYixdx1zek2/Fhc7tvK73SuNhICm5YdDEb+/6wulgcVjv
b23n4d0wy2KBLKUnwP8uQXEl7NDojrShtdSiTtBHLhmbBatzKGKimgOJ7IUX0h06
OGsNn4OM89HuskEzPNR+Nyi+7IK3nicxf4Zp8oTEeNaNRxdYzH16ig1xWA2bhrSv
e5M71tYXpLrTA4sltbKkmcUyn4VoI4ID6bqOA4w7jl+18yCYyK3IsxOuBfsWt3VQ
oYIa7EVq5O/Yypiq24vVVTg9R/qxZDcrCxd/GKeG7KaR6AS1zoOY5vWRS/zT+LAg
jqZHRqURZrsBu0uaKrfExATrvhJ7cMIW7k8ARFNOaub2DOzUMYvJ8TZNqUjp20tX
nw0SYCzbeNvvpyn2n9rLsHBB0Mfu0xb5ganRu5lctuJjVkJOUP87QQTcHKobC/fz
YSEKl9LJsIaOxAt/30K2m6/a9752rAY2F5DV1Yo7ER6CNetu2rjSoJq8IcBsD/cj
wlYAbPSnqG4BB+pJHdFbIxSlqTnS7NnFbfrFogkPcpNKBVUWwFs0w//Rgt/1wnxo
0VnTBO3XwWTTa83AMyqDx0Ne6YV4VDBwbqg+Rlls1Czr9l4mWLmFsszRf5lrApZ0
wQcjxz8ojXbliT+dDk3qw/0EEWJ7NSZx7NycP9wtWOg1DqtrYYnyFcY3czOMZadV
NGY/1A3uPy3U3zeN8k1nmZfa+fWt3AZ45ZxxFq9S0JZ9wtUbGXE01I4hBMyGlTaz
fAkeDMzY/w1bzM/L/ajrvNowgTQoxm/bAQFud61xyBTno51QUmK10mnEzdnPMKfp
+DioqU8fXm9oEuJtE2m1vxFY43uxFc+8A7ll+WwJwgFaa5yCf7scuu+v996ZKTeI
27m8tK+3D/eKBFEIHPXcQSNBTtB26i3wkoqcTiTaej7rpjeF+4+r+G4mZh1IOLhK
o8nN2pWcIpBFo82fTKX3BwZ644jT1NypvIN+zS+7Pmy0nyu57YitJjK0wvIHs7uh
zeRTJ2HastyyqvDvW1tCOWaX2fkLzjn9XuOXqNa67ck3YAW5GNAitJT5hTZsZYUb
TAjve1aH8r+E3imXZS2fNlU4Ml13quOOx4rN4QMQFlLyCqU73KkT4VtX/40VWQzH
ePyM+JIKvdtTfBCVHboy0+6OWVTDI2jcFsDy/AJgCXUnCFISOuAuj4I9VCW3qErA
1WaIfiR2QsZgmUjdIU1WUwCD71xBOc/lxMi2x5X0KduD2/jjk61n2VdPGo2AklCj
kIriH7ok1YBWxdGFATOPqvG458IiQsBoJ+IdvtLpENACJDAT2DvGE9ZCXn2QWy1y
97RBaRqux2s3SaSyxIYUGrbtl9O18agDLmhJ/oBQFE8ZPi6i6tHMeLYBegyIjT/s
94lW0QnfmKpd/ifG/WA5k+b8wgaDcJU6yzw0uPL3H4yklyubNkpSMfm6DbNSosfk
LCe9ZJTd/t3ouXrEkiM3bKJLl6EjWVT34cxljMfCNANUqF009NHz1xfFF4dWMMI1
FHF5If7Bcir/GHKgBvJS+MeWhyLQbIDtXl+Ix3f4cWqjCWgPty/7EgF15iqkcAHg
HtuIydMMF0TuxVOlguxzIaZQUunFmZ6ZJ93+SDpF2/+ErGPd2lL2NRyDXIICvVT0
SQor7RV9o6gZjLGaIxgHY0i8/Z2rUQ7X6Ubm2ljy+53L37xog9b78KFRElwYbhw6
SappwifxMtENqzxfrsn5lrwJYlUT+gWn2YeGgE6KkzBMmnFrXpaOaW6H+kagD0Bv
1lxVGkEZUBEIG9Sl+Ov0YDe9eHZb00qqJNtKY9nIB2BbNQ28kPckicSd+VpP4alv
k1+3SVvBR2LTo+8SFv9BMq1eqXfFrHY+bq+8stu3iqRqR7gXNE/2Slym6am0V/Dm
zp2IVTdHeG5pN88OR0zwGDYUtwwkIdDAw5z9kUn6IGIfe7qu48U2a9PS3AMA5gBk
/Vd2UudqGDVP479YJVuZhb2dNJ6K9/ngb6CPrWY9B7FM5v/tJ5sLwTGSEm0AYafm
oPKmBfDMRiq81yCCW1cZ0MTdRRKICa0FOwPi3Lq8nGesuu0OilbvqXhKEVxXRkK2
6TvhmgQJXD3xndmnjDuD7T20lq1JUl3u+7IRmf/wqHlZwNVIpUh+LHIwKWwcbgL6
zP6nb8rwGU4N6OO2GbUVC9lLpbQMLgzCTk/v6MB4LEdsJOeCuTViKVespWob4OB4
avA9xXhlsuuzOfEI9MNwW0ZPoTvnbKwUWefJPre3BEPVAWNr+YMVo5/fBJR2tiAu
p9iwwA9Lu3E0u+exJGdGSCz08FXuPK0A5q9DDwd0Lq5TRN9Db2auh5nzPR0ilUGb
MvhB1Mu0s45BBFBYB9weJTQEPdnszp/K6UBa02a9XbNDQaLxtvuAc4wCj4xVWOHH
5aYxxP0sghk+0CsE6Iod7Pu8R9pz53mr7TbgZnKi70Pv8lvQ+EJm18YVQLPPLL1L
h6oqEbo9otyq9R5k2LdlywKbjixMnB/cXcu6koD6zmn3j2zExz+YLc9YXbTMcQyi
0h2CwEXXu6qZGi9yd7hh9T8CkrMTy584igqP4Rb7R/JK2GuLxLiHmoHaASU6tU6B
rZ4nFEVNxBsbImkkJJeVJhZhWpQYoxyI1OqSWLAV6yrsiCuEiCnvAuYY2C4ni0a2
TOy1RdIFm94YmtAcQUeLCkxP1CuR/AS0rHOtDVmJydfGjF9+zCGdOJj2imL3WRs0
k6IK+BoSWERRLIZPZGg4WNPCPbR1CVxdYLpWuCovaqi+KKbdJuBvMsNwkB3H01rd
J68dohUgI+V0U+sOWROPg9vIzhqL7VGsWNwgxuR/vZ/kCtIFR9tJE6dL/M89b+0R
tsgki73c6fy/c/gxwjigTAnZaDuApF+Lu3N+yfcTPXgymMTbtNkxSi6UTTk7LmQf
nGozHPmc46CiIjuOAgIr8roV2pFpRzyLBFMPMuzP2seH0dH/N8wJUXdEOz3aYYPT
/ZJB+GUrSulnujrejx38KAUmWAATQLA4FVsobFHyDDXuJrRj4+ZuQzgyQoaIUNbD
reksXUWlId3J2gaCuEM2CIvVwPRooxi/i6JkHeQ1Yla/UCG+Hduy7TVAScn2xT82
G7GerGCMaRxq3n0Z2vchMcXkhv+Eor8yQwNpaoPzWolnrqsXQ1dB79Hhu/yxR8MG
mhNyIv6r1P+nr2vrCV0aFec5YIKqM1iZnVjHGSn2GBlqH869eatR7WiENZcFNxBo
bF8RguT9kjhMXU6UkQQ1YzDO8y13FQ/tckq8KFQrECPqbhxbBVUDc2NNyEZSOZ8a
LIklIXOGMj3RhcWInfF1D85Z7t+h06lj0cIUbcElmcBUrMt8FtbAw8mfl34ASpy/
t098ZluXmcb3sWmuOfSTb6dCvc+zdrvjoSveALANDYbVXeIMMdBkkDpy/8vtE9sH
AdeUwnkBxbAZXCV1ufkGPT8sEyohKMvYlaKuCH3mSR/ixastJOoW7xxFHfdgk0PP
oohOFsuAfwDFj9WSJkAB8kQm5VSLBrzOCgsEt841b6HzFTNkzyXvnshltmcm2uef
GCg8FBnaqrrVSVhTEnuF3cGpKl1AQgbqleO9WEVTBXlYbcsg/S3S/UHWbI4zc4gT
99fxJZ7XUo2REX2vJiXyMCY0Gx5T8Cr2ckNT3DHEEoHWHcT9VOX2FsFjH3YV/JKK
QCX2dgGYtryfPS4RGN0B2QrYgdZIS+MfHq7mvlnKhSwGE0Wg6dhGV0RztJMOH/d/
muEU+uLeq6p6CusISaLIi29zsc/6O/rC/bl87rSJYOZib4indLfnB1BsGSXlZBqy
OZyiadVwZ0HPtqq9U1eeDr46lSX0dMJftC2yviRxR6RKCxi9DapnY1VhqbdbO4jA
2HX03VrcaR2H8qSrqTJikuiMswhePfWIVjgMqAIKaFEoy4BMqUOatJfGtGb2p93m
Wk6WXwv5fKvSCdNuJ4vP0hNk9LuzPSBaG/IiFKddHwSLHuWhGPBOf3ZUYvMUfIPM
mxuqy8zSLBT5oN5mgyB4/hp8yHmxf22Qd0n5lW9RgFK9Vzmg5mGfmg1UKcZqCmcm
8UuEvCvCgEFvRU8EMR6EWq2ZA/+TJJSopsOmcGwgEbyWoHx1jeXW6g5tzZEm/PoR
8qx+0ykinjd9T/LkjY6hBmzpTnNfHmtBBgOW+9PgI6cZ8x5fTynmo5gJPUsm+IoM
wJur57IUvhV2sMHhyAJ797fjf3YDp1NZRx20H4KhYL5di2xtuc0jny1XEkU60Zlu
bCP/0RAOiHdkyL+HJB6aWorvACwDTRYvM64iCrpUsznvslNbX8zTdvHRMwLMFl+U
/9veGXvRgE3A2c0r7zsM0cxw2m3SBTPVsT0+MPZIFy4BL6IrMkP0aI8uYy51Mqy1
OKv3uAVi+tz9N3nO+W/h3mPClNjR0THpd0QG1Xd8CNu2Auug17SLiHJstTzelDcE
rukPuPGR9OcufFkjs1Jy99XJ+iIvrdttmZ8jz2zL7Z890mItk82Ywu1ZT7sntxhN
Q1FCSREWuBmYNW5mTyx4d6eIGkTQWn33UrUaHOxJ0aJRJKTe91jfqSTPThmGKMqj
Km8fZp7GeVB33DW/u/j/sbVgrj2tDru04UAToIKuRgMcnG4g2cb+VbCgmgQe87aH
xK9Mkd1kii+AfEfNC9T1OFFv4sbzt/exBaeIgFkuR+EQnR788zQwHBocE5YvKcd2
i+GW4OGWMnsvPwrEqmAnxQz8fzGjny4X7gFVmdCkdPDA/rmAmd43A5boxPMsQOyd
xx8ThmWvxjs0AD6gRMsEYRuaShGTWe543Krvau6iF8mxlybCYntBu7Y9H6bdmopr
bcGEqeXn28G78DNlGnQaK95hAQg03ktBNwurUX3EJLjgfRZCbnq0eM0zHsK+5Q45
w0F2nGGucJpZ97VS8zm3cjlnje34l6eF8yXCAjmZLM3wuwz2WUs5yreBa5X5d/Yq
slTFrs8htKXl/kCJRlPuG5QVSYhaNjsqEn6ugf+w16gSUf9YYQg8+3rC61xhBSEk
8s9gM7atciBkiwgXr99Hw3XIPLZy0E0Btt3tsdbW5AdBILEos79G9aprLEwjYEaj
jv7DT6bNmf8zcVpDvF/RBI/hZAbu3zsqzqPshGA1U3ukS5y4ve4v/AjsKffxffs1
T148pyJlh2CmBDIwSMPH283tnHbYMe1XgYqynijnYrK0gkXhwTEsP9L1JktgHhOU
KZ0IEA5uKprOjnBOUSLrJiDLMxAvCjMXCwYZoet4fO+y1PkRURCRPeAkws19U4iP
migpq6s1armBrOfPhIphJXgL4E59Eq4ubDia8hbiohmEyl+lpWbrA8vxtd4gykxm
JThMg3OshumsdSUx1NhwtMLXNBdHaDX7jTm1rF+it3pmUNmszoBFpKa2807BUl95
sX6TdZLOO+Jy0I/b/e0Ydf0YHjm+2BLzXvLWYwdtnq6HsRI2q8bKFFtGh3Gj4c/u
3sDefYMG3RKQJeafaK1lchb5hHIkFmAjtlnsfRwnhmk=
`pragma protect end_protected
