// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A1L8YTdlH6HAdvtRMNpeTMC64vigP0X1vF8GA4QncGRZBZRaWff0aA9YGf5PGMJ4
hSr5JSG4XvkwDulI171vO8xxDEMMWd1npup5sW1rBauGHc51nY97ZbwIRytPA9Fj
nUwEajxNkD62waqoDYAOhQgeNPAOfK7My6fKsNMXUws=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 68176)
HseSQO/4WIyufxGFB1msrODT1yDgZREJDtixkJ7u70AOUI3vvbXkuS1MkIT/4R13
/+ffsM9DednrDus9Ut1qoqbvE1gkN2obZKTxX+WYSDyC4jBOP9CcZ9nLryryXwsi
w7cTv9TW3prxith3Ftqbvc9foVJPEpjkvEL1TPeJgMC0Q+kkfvq7qGkGhVdyVFkI
DfzSZbl4RRhYYTjJFJju9SwvCd1NSuHlq4MWXV0ULkBWz5MTVSb4aHPpTApls18q
nKpgacsMlbAc4TgPephv0l/VHPDqmtykqAsczLgWnLOXAtah9tboZnJa6Hr7BGX/
I7f6/CjRzP9tPmit1LCiJ32jbSQheAi+N49nokIs5mtr6qwTDM0z+XDx6fIDsQ4l
EU1ayajEQ5SbMVEupUb6Ek79VFqmcU8dcTC2E6lGPDvHGIkZbFrLteX3ZGznGuhc
z2KQvY0r2HmhB+GquLFcuDwhmo7wJPggwXAa85B4X3X9S6844ZyFpd07RA/0W7S5
BgdL51kTYMaTuLWKeOpI7oRLAjeMOXGgLC2kahmlerszRTELNpCI/G/UDkOHs8f4
m0/I3bWNwZSd1avHc6AJB3YgQY+AGuN+BrwiWTFox2TthGc3yYR4vse86bxHtZcC
klQ3nVNDMZUG/FFnWkC6k9UcIVIOhjN/iONTXd/j0gPMhH1wEzx/DikRxb/bQgGJ
lUne7oG6PGnl5CPD9zC1uAnfatbUZ8naMYpt0i0h50eR9H/m4prclj5my/KIejRs
dhNttXlSbNqQLUrO++czVkiEkXAiBoL4x7Ap6rHLlX7IxWB9v5DDi2SOSeH58WnG
cVdam2p1jXXdMw3lP44+m77L1fqsRWpHhOvs+4CHzHemYVi0A25Snsywt7yLN2yw
79BM6HtLHNWbaT/ADGVJXmoo2x3ix4DfESfkXyrfZoFihq+3wNSqTYM8wHIXnsX0
7MzxjWVO/W62O5xcv8GH57UK4+W6+XHFWucVRoqp7jiSPB99fzd5NlLqbQLUmULX
LVVXP3MOh+b6nuZ6SQSglC4xYLsiD2vscy42wAM2csArml3yO08Y4ri1IdU98ccL
wym9ZRhKsY/QRsvXcfSpkzz2zXeRS0NWsg8fhyBLJnHD1ZsN1XkAapFmiyM2WMDe
9eETkQnKraO4hxeDZaOEyQhy7h6st4lHPEiT6BMGq/uzvrKafrjP+2r+1aEiKN7p
jVW9gF5wCVkAW34PkYTdZVzYDJ9l+zZ1iLUEhbl72fVM8krvlCk8svSRNgkw5lxW
5PqQJxbQVgKekScJRwhNnyXo7kmZk21lyH1HPPHnFw80xewkwR9NiGk1kUAX77l0
kJV0Ed61caDn+s5uMZ88482zWXCWURGWgilMTYH7tlXmpuEOm749q4/9G8h7G5g5
GcSSZwfD3xvUoZe27WDToZU9a1ed1b4J1loggSoEzV2v58L8t7XvbskeP8O2u6SF
U64VlfUil+4FpXci3s0W+Tq1NOi4DSFkLPfWtzVVoYWK8avglbwHpE5Pa5/9K7K8
qEcb5D/t2+FkWojrfw3Xj2veSRPPLnRLkrzPSN5yDmnfVmJktdwwuTseNMzJ5Jd4
ET0WdVhxNVHKdn9r22+dfmpDlZKnHeYI1L1xGUys+mtipJ9XJ27Z4P4tpRevjr9g
11DgxD+uiSOJIXtoR/mq09MrHrsUgX2sPj3ISU2HGRyHocrR/zh4BJEwjpsZLuPn
QwlkfP9Gp/l2Oel5lDHxvwVigMzefmkru5o+0ZXYmSb2lAXxxr/kP7/fhK9NGTlz
6FQoTGXsmvVtRK26K5pMQ9JZ+gkCeqoMKX0MkL0pvkYcTQqKnQi9I6GSQw+RZWH3
EfzudSsqxCRN135vEjJLIpV/9ExSrDk4RM3PrHL8aEI1d5+i7JrdG+1J8/HpQGb8
xsbWKiujPmFWso209PBxtCge3+Rk6OGG8Y89FkzndzHvbmQuIDAXUYp/wdjN0EG5
xrckgcZ/zox994S7cYoeMaPStyb26HjmQl+cAOtDnY3kdKKVYVNBgqYsQQQPQFCr
1IKKj1nt5T1lM6GuJrClpQa3wBN0maHIpwEMlJGWQo2CYpIcR0TNR5rophG1c0gW
vfF3jrbZbCVLc2M22l+WUW/f28kbHtrpfZQ1q5BxuFq1IONimDxZX4Xz67QxIhjq
yk++N2SRMJu1O/16/lQECssnXJh55bzwdu8fyulWJzmJUWAB3yRg3Zl6Bz2s35F6
sqs/e+H7BsmyWb89hb4ivHR4bj6Dl/oyViEUPjiA3JiF7TbLV1mu2kHoFBILO0CG
qBz1HKAPUsGowtXlwL+RTo2Iv0N5WWtU394gdUK7VBIOadk+Kf/XCG9efnq328ZI
fDYq5oDr/1rr/NOOpz020jDF70Xu8gNnSQUKjTEX1vFYp/eeV2PbUbIZ05Hc75l7
Gz43hJlEj/YY/AIFbZXJ9acKiHXgvF1M0i+B+wyre3hqpycmwlxasr52eXXt62rQ
vVCg8VTd8FPKQ+EQN2IIm3rBuoSDskBLSLvAGcYCy+RhRydAGd154AiReIZdp0da
PZD6JwUJghQOKxwTcBgtnRV4eI5Mmme0FyU315+o34hbKnOgO0MmKyQj/fe0SBo9
e7DYgUOdZxwaKQykEHYzjQEMWMNewA8kF63cWkBxz5ax1I3UplyMUZNI2wQWpa22
KdPfEgSKrsgoi0iwatVlpOS9YpEL2ykk+3RzkjmDJDMjsaYihytZ3fz1JbsmUu4W
YnZkwFrtVT1CnjFx55CI9AwuGUbXNPfHSBsc/uRYka+euSv3Mowceo4L8IEPtej2
R7n9JnvEXjEsCuZsJW8QNecfK17skNdETVAbcC+pxGOk+cVYriXskb5fnR/G5zdG
gGNg7gBfbU+akSOLzg66AJoNdjzkcZ2HsIw7LMz3pr6ziJhJUBffgRcBlfegc6Lw
7md5StDoAcA1LchiP/BqNCOCDS3GcGiWYkW2ZZ3ErJ8li0ahCYZCn/axpo1+kYLQ
UWsu1oY+oVGJT0cuNBLLYtLw6CDCwUU41mp1t/zvySUg3W0LI8LymBtGl8AJdEDZ
FfPH8Vqgk8kCVzIT/4tPBRVwgT5sDPXvnzVErzKM5GvZ79ibC+dlOQ8q0HNxQuPL
MQdZbyUbLCtYZRSz4viulwIJYFn6HImrnGakveYO0ah3vvnIZ2f/rOC6ox10ljFu
lLNXnd6K/qPiE4ssH3ctggDcWif1H7aOUEILePwtlTHozCK+im/bb2fUWXBuN0bo
n8qTY0e6d4oZPI9+NyBLdbkUxutwH62HQDeO4mBxoYKNpHBfnMN6vNhloQPqcqkc
+3b532+sJwKaMWuMeSUeGKfDZgMv7qwZALTGZdEcLCAsvoo9OGo7xR5d6nyWDmMc
EVtnth6+6nM/5727eG73m65p1egwmgIVvZ5TGTwioV3oSdt/8DbxrTxorXH4GLGj
b/9VGFsFswkBFDAllRwNtLWHfIrLGc/aBtR/5OHZ4sEp88nnUsbKto3UKBaeImeQ
7q/N8u7RvoHL7GgYIvCrPdA0QiABfHn+qjPfY0T9kNIvsliRFHibrCNECmBsLkBc
jJwcw2df4x233bimpZEJRb8GY+2bZaU3VLC5LOuMJ9PXjXxbDzYFjdVZjM/mLmFV
Mt6pgQ5NArkrnZT259AOguXqdZe6rAoXuK1qjr3O+LcUNJJgU2Ltdm1WJbMlcxOu
kttwOQhJm+CC1yV1VGJvleshMDiV3cDPlG1wMqonzpYUuOiC5p0n/PpXmStIJ690
aYJ+81AK/4EypUyhIpFL4CuT3pjyU4ImcF4pdJHyCTUMwl35FQLY9Wu7pazwAJCS
Grp8XcdYeUkA/lW4UCMPZwscQyfgO9HoVrryAlKMdYtAE1MhfB/ZDhCFNmgn7IpP
PEOtd8XU1MzFgmM4cRm9u8GAcOhDr3i2zg5Kwg115tP8YCMFQr5lbB8+FxfXQ4s1
y9wTZaImERtc5jNLAKgxHdjibi7vqevxYglCvIzjGCAgKeI/vAmygGQBK8Gq7p83
ddrDoaN+UJKrE/9O49vNuRlIpizOCh7fc45JAeU+Z66/f+pUt0qxMmt+yKsvhSmg
bqC9adkkZ/f1H2cj4c5s8DCHW/mGjjnqA/SSAjAGmjNPCl6WAISFtkuVj4a6Xpxr
z3QzM58cyy+XySIN8CwCMdOfACCYKMbgMXshDNmju5nSJLqunYmtQVttoIfvP9pW
+t8mZLnLu8yi6pj9q1Nwe3m7J9SNsrscKzy7G47cLNTtgIED7KngY3V/S8Kg8eK9
4q976fXiREAWAqo/0gzQU11A9dyZITcbbgCWskPpWrBTNMIaP3jHyaAN0togBDz2
R6c+0R2dqGgTzQfgOM7rjfJbhvoycHlLqVHz3KeRBtgB6z0WkHigMkzwADRZESG+
YZl0QpwPgB9Z9vqMXb9VEwnPtoSOok9lDoIByRgSDRGDLZvUT447J5NyAWl1OOjP
QUdHlHaC71tXPpUpDdtgJjqqhBxlUd2HUmO34dbFBvCFxyfY2vx/jEv/7NvPfrIJ
XeOk3QuyPVHydY0BxLklWxeS5A/zOYvdZHnGpryLlUeBpPBN7WjzSfJAZYbJouSs
/P/QF9ZZEUIEUjz6BlESbg6PItJflENpR1ZZt0IppjF406H9UT5Kc+SzJ/lQb368
Pp+0KstmaaFhpcAf/hNCtTdR8W8FjYPkoOiMvz3YUPMoMH7Hi0ZHYcmFPQDH8VJS
17cu5QweWQPMArBCku5vTWtJK3yfKFOkqGnh8MF5tfCNRpPDQ3rjhXWZrrLdqvXG
vvYr9qHCYe20pWtbWP9vMhFp07lokTzAeHCgIohn8ltLuTrnspW1cODoWloMlM28
phgVtnPpYaI5ixM2TOrhKPSIdY3m6OUyARujWl2auOHJs+BRyQhF9igMfuGmqPEF
1DYsynNvrciAgyfv+mtkOeYUDXLuyU0Lx1qNKkz+jRP1EM/8Q45qCf9cOQBpldQa
ViysiiuY8/QPAYdWcwyjr6wSOCtowOfY1fgTUCPjq4xdIHDQ/rhWMqObUngNepDV
1CXz7p4ifjAdi7bDNS0ICBwxVxHAZzfaVVJTv3gQLSS9gvD3D4+bRz2B6mpe4lbO
PvhAKnfK8+8Gv4+f/cryGxtVEV5xxtQIgvQ1ArKJuFkKFIS7Hs5ga+F/d9/LIiGK
V+0PXGR+NrJntguh/QOmOcmaMEDM+EKSotjFK9BMlFRqi4WY6cFhqWFf2mH7YaEy
vUCNI6cv+HebW6s1iDkGEqqW1CBw2ROqZAYcTKVbJhQUoMP7R4sdO+tIkK3caT2d
FkjroJgbS6Mn+i038XEHDHnfn5/0Lh5o5P/qPb3ZTuE9sSCNN3Se13VbdUIpNlQn
E2T8q5apwWGttxHBdwWno2VCjsFnM5GfBpI38EUTGhPbXo2J9XcwVwrXozxoubHT
BRCPUiLE/jsQdOhi3yRkRdvFPqQ1y9RVxC9zmBJL943pG6tWxnh93FijmHSA78is
q1U5Y4ZiHsnoA5cqdVLfIo89IeEOCYA6trAZaWtavUHCOnd1H9TaQ36HM0GgPSJF
tH7oBhLh3W59lBrk0Z51QVBh1uIq5KgYjEv9Ik8GFwGGXqN5huZqy5Wz0M0rvJXo
r4M4AVEyxB1t2cmTlaojyE5h5pKbqxDOR3JNTOXVITnmS2kKecFxmoc+MUEpyocX
fp5u3NxQ1ZvDYBcdLi3FHWXGGgEgYnkTWTrUgiIWarHYnpWkre73L2wgx6DPTq0K
Xm6OXf3J8JRphGFKNkhVmjrLi+WPZZ4kbo8IprUvyff6Rz5Uh0Isioc+jsxNwqJQ
Wbo8m2kPWPO/AbJtB7AUc6CEUZyaGOmhxYdfek5Oo5IfQKjyNtdeuJHuIzHbq0fs
HFJZr0ov9VbMrnrBGdbRlzl55JN2hYBiBho1CdOTY3ch9aO0gPlIRTIC4gRJcxMt
Iat946AgF09t0LpNfjvjoQ5LXNTiQk2EM4lZNFsrPmraivBY38RDdwEWKOsmtXfi
AY63rDw3OBs9t2ziNMIZqv6yPz3phJ5qCc+I8MGKHwo3W5oXqhShuIaMk3B7nuXb
cneeh/AYAIB86j7KZHG44EqHdNSmjcopI09VWiro69P2cyzeOGIKRr6Aqt13kKKx
cvWxoD857JK9MFpKHhNqmgM0MoY/CU0hq4SdAnhoQpKJY0H/Bvir62sXkIjghUbR
R6vyNqZ1eCi/EBtaMkLM79WPWcqR1dK3/0rKjKICwhXtyfqaoj4V6sGUvYSDlTTe
dEmbpS02O6w6FGMLUz0lWNu6sKAoi01C9+SydaqdkovGoVGTC7rgEysVAYqetjuw
x9/lnzep4dud/TFjlDdRyg3vQFxrx1aFoXiFyjucIZbx1o+DWCm/uSYsAXVOQp8t
6PN7dk92AVo/cpM+XPwSimeJap3Ebtz3g//0IUKaw7y3LEmgZPpnsWQLm3hURvr4
jQSkGhkjhkdcQVCDA1FDtW6eJ8g+X54h0htbbLW6o+zsDn1+S67SXOhuz2nVzQ4B
u+zKQ6bsOtfXHmNlpeRGTfL944F+YrEsIc9q1C1mMwbJqq0u2MhBWDBebiAg0awV
nYArAkkkPPeXeXyW5ZVsY91bV0YvRutvikp8l8WPeefBuTK+M8m8TZAu0FOS67Vv
K4AUuu+nY8SkpKOWSdZBd/x1+kFoey34+MzR/HZvVyHItSU76MbG2Sf6cbCg9ZB4
L2eAhgR+bhpTYeNOcM08qpSXFjF1ERf/Ngi2zMjoo9GgkHer6Sh1CnLcl7TUqNGR
JBq5x49mZx0h5JlvJ6XXmaoDdjhwLmZCpGTacrScKidhsjposEBKsMembOjIRrol
wy/vgcRuIarPcxnJ2o+wzbNXgVGrrBAHUdCd7/u6awE6y83/EXkb0z4wuVQlyLVC
yzyZpLaNgwLKn1KxAvrGNw7sQNXT9UdA9xy+8HMtU+e4lIx0lVuG/gMyjwVmisCN
JSKDf61tZAhx7sZXlUvzw2uP9avZAlgmAxkhQ6fENtFYtSZIolBNb1NIXpxDWX7G
tb8nkAxUzH27rXfSWG3Qr10Vzh0N1Cyx3W5ZWP1qsJUDmy71HS/9t8Nem0P3NUVG
Hjk9uVEbJSVc47TdZCsfVUYkeqAKIPWFfZVnSWOePoGm2LJHjwK8mUCJQWVDb/0h
bjHycuCuorcuzm7iIhaUuG9t+iA4S0jB+9vYgszda1bP6yxrrSP4HPvtCUKqDOYN
Es5/pK2BjRtHw4RnowCcc5rEslAIxFaQCKrnm/nDafvb7S3uUOATnMjtp4nckk3f
8QqPTcXj+fdr1+0McFYd+Omuon/lELvl8SOtiMqeYeQWlIFyKtzp2BSrFFTMMay9
NY1+6CbpfZiHZHbMuoybtmMmO5wMCthMC7Jxn5YueTS9E3Tg3D7iuycwQp2RxDtx
NccUaht2yUB53+bXP4F6Z6BHCMYsNHn+PUjhMCwdZvc3DRqTh9WNO/E9Q/AhjNTo
YxEWpaqeQQtKmhaz/AaDw7M5ZhvsFAXsESOdsDCuYUcRT3eZSHI8YwhZPJzzK3ha
Q8M57e7ujjcag8h05A1BclSgwH9PVa9kyfyO1xvLT4WRndLLTKbaWNUSPgUoloid
TOx5XSo5VpazSat0clRALPtuaKbWdidB+xJtnYwTf4UqIONqfBHqYpAnozCF5MUe
TAaSnw1nZbr63RYzth8LZtVNhaZ2PnZc4r8019K9z8Z+onZG1ZT3/b+/nUnvEgy8
kKdVcYYji1zZN4G+brWhvbeOa6h5nwYS8a7yfOfzFa7zBpt43MuCGg7TDZK92atv
785KVK0Ffv4vVNS6O7SxQq4qCER/uqF6uEvd0/K/77iq6CdsumLy1BGwsscDCg6z
kWa7xZ8GdYtS4godfj19miEZEI17ieVL8c31tSgCxIXUC8jk+hZfdrt0ofbYcW7U
S4zkpKWbTPPqf4T+retPF1zDHAu1jNwOxZEGkDjgNKk5N7N2qmZqDdgtAXv0rNTo
n4+waMsQSc75hiztvOLIKpNJ7yrW80tJqCQif7cINDyFdT+hRyGnGNtp8Flzr2ea
ixT3lEreerP7yXSekfYbNz2C6tBASxgqU9zLhXjsN/aQPNV7SEuDvpswV22kZ9T/
Ch3jk6dMgaOt4cy7Aju8SIID9WY1xYlLjS99zCezjMADDTeUuiud/B+FpZx9ZcjX
8lYyXT90SOHIQtoVaTBrzK4C64QsvXRwh8IGGhEqq2/sCOZkL/ltwO38ua6l4yvr
WDlMIk9BMIqG35Zw4O2bTNg9QKyGTGhwU1MeZdO01pNomyIN3DmCOplHKFbWqlsk
ixtx4WddXIrRj325ovqlinPHez4dMcAtmwSLQPDFS9ePJP1g+mqG70Q3hK5O/h/c
kNZrJoGGLon9SEkZjfSe924IC1N18+FeowekASyk3mzHksOM0OC+6NHLZUcQTZxy
gnleLt48M8N60nsRVFwnzxXH5/dUEhLTFu6JX8QvAF0F4K0PuyX/cO4hyl4Nu9Cu
zesTnoJXxKS2Ko3ler1DksGDf5VGOANF/Gk4SXQJTFNInYdzljaa1VGatmAQ9m0T
34yM91xgMzlN4UWUmxsmWI0qqr17brh8NGGYzZPn7zINKkLqWt0C2534taFQg9sy
teoVPde+IOYJO3/q6f+IloibfTgu4S1UOt43/jCXLd7ChTfSiFJh2RvEq9072K/z
y1JJKgoTFFHf3dl109Acoy8Ie4J9FoVkKR8AArHzf4spg5KCQLz8uY5+ZjkEO6DT
e/lS4DTZ9ukkzpRFDthAhSU42XP9dEYVCLu57ZpPrt/BcTjE2/TvLJWEtHihigtg
J3n2zXvj5McQipXjm9H0OjWQaiuotFgYgOjnFSJH0ER1o9rTgGCdGZWxEJk/mU/V
7+YSj/diL1niKYsd/AVGvOELLwQ+hIM4Iba1U9tMqrFEI+RuIJ74sJ4Zcculfj2+
2W3GvfvlEf7dgilbmCVncbGUDxvIjow/TnP+1WKNg9Zl9I0HGnn1+uruHyARRjHr
x/HriC8Rji3fDfnreZ+fom02MYUK4j0Ju7ZFcNfmDbAmjC/+x35bzQIb0s8pHsvb
XyNDJ2d8n3/E/tBcKX/1aHQ4AIT3ghbnt/gaNVB5lcI/e1ETUUB7DDLitXhTQeXj
7xddO/7/a/iCHqj8sYmhBJ+1LmbbdZNhsQUL0/XY98gvXYuh1n0FPaf4G5OfC5P5
sX1xUO/q+qj1TRn6I94R17GAafYQrSTnatfG9pBE/Tc94bdxOg/Wrf9IEMBM2ZLz
Psk0XdvI92e81Rg7geV3DyrIomjShrVqWwL7Xt81hRaINJUGlZWQY7MyCL0w6R81
qQQps68q1fYW5p3ApXbIfhOKZqXAh/SQPBTA3wQzx6nYiWQOdLt55UUehLTpHmn/
ViFCEhJuWkQerf7M0juFNUjxJfCtBGndPHLeUXrxs19dJ2xQhl4ZxhFaYvIPowhs
2OOLaRVvvLTpHLgUGxVxFeuleBelpWwcBog2/jSQ5PPVRTmCPWPZ1n06qeRZ3SnS
Qlp6eG8CIhj6nr5tcgljs589LN/ZnnNBi43LH1qi9i9JrqNJqBv0RnG+EcGrkLgz
6YbuPoNPgY3XYTNj/WIypEcGHDa034Y1FoiWlcg1w7hSGOSiJe8xW34SLJw8nTTh
BqOIjyeg9I8L/B7ye3G9y5bG5bLB+JVrb59L1/vv4shTJR12FZoUme3ru645IAyz
NqKJ2W8C1/3Iugr0OoPrZdPnQRib4+7R7A60YMJP8bqQHKSWxA3zuikFyJVZQNDD
Zz1VV+nCjwZstIJbw+i+3DcngFWRDqCkPK7du8uruv/2uIdlpulPjPcr8ewvcigi
nl1luFSm7b5HAQqC57FJ5ug4H88DeBYcl7JhyGanIMXvR9vKflRXODrqblBjQIU6
86qr53azq5XIB3nwfw6pq0l69840xzrtxiO8exIp0JP3Yb7VDWIR0tebI4arNytk
xZlLu4D2nVTcj0lihFRN9rvv37DXG2iqOm6EfPWr7F2SI9Faeaf67BHb79uK8nuD
mBOd+j9PW6rUA9y+/d/LdiWdcXbnlDMpWusKynZ4NNj9XBWfChiwv7xgceIUujva
hbmdBLZbyfWDixAdnkIfsX/MKTFBbgJ9ycWTzTKYlQ4IPFBdZbof0xrevoUixAcb
Mnu5wijXuhzM1eyt8UZbEGQWJskdosFbWuETRbkg+C49YcceYVZSNifcCbeEOuBO
hKhoM4z9ZkgUQ3BoO4Ebl3WED9AurQ17Q4rNsTTRkO0RQ2+icoahUe/PBRRj7c/8
qILBqbfEQMFXfXqNizg09zIrCbLiSqrzsSMY5BSK5MNV7gy3PYkBm2wmkADJgApf
+OQKsrVfDQZ8NqAbRZIsc0ZCZ/R0eQ4cyREHbgIJNHEwYCrdIAP/kwwVG+/MS6f9
Uw5/M2UnDKkRFWCE8vVpQwRsbR11FrizQRNhs9OGWOcVh5RXFYdK3RQgn7hLa0ot
OEEZz31NxM4/2DJ7/VjQdPtKyKF/JT9U1hDw/R4M79NxqFFjAmvoJ0q3M8CDzRs4
RthuPNt6DxJL4QPXZMu2uYyHQDsM1LVX+qm9UODpnWHNALpzMCg0tINmKmZjIZBd
j6GDb3+AZUZpqIXpSAVVPM8eLQuIdREz9v3mlw8DMGS1uGervGmKUDpfR5yfiGd5
WEi5eUqGDhIQ/sifYCmzpx7lCdHAJcMpHWNbMth+rau/yP+kLUgmFPknS3u4Dx1Z
qZE52WKKgVFiii4rqaoAuybB3S5aRQ5PzXgeDYG+d8F/bBainuMXWJPUyesALshH
jevTHla3nZNuK5TKoJOPiQSirEa0U5xLWrPe+rrGlRwTUFnb5HIdSrA5eRSFYvzS
VRGT17xUtItzPV6ZM2GBoZX7IZs5lTPR5PQJjTr05IkgpWG/13baayYrAKrKf+tY
kli72B7+JwCO6qtYyaUpX3Ixg4CLSqwOgEMyrEIvIRPDEKbAgJlICSduU469cIho
KEjtRG1GKCa/15akFSfVpbEue+kxhNfuUyrM5sYXmETbeVGcVknZV5Z+1kubeDbc
lcjv+PniKPl6ePweFko4aCUvt/fuQ7IcdkEe2se4TTM6BJ2Grewg50eGYpJdtf2I
YeBGgGpG9tGP6d5Rr83pzVanZpa1urRE1YQIt0nT799TwiOZzv3m6790EXRjT18u
wfS9EA4becdrsPWorqCnHOhkAu8bZKml8Rkom7qOlnLVRj1x3KLlkoy+3jDW8Wbf
iCByjic1BwDCmKXx3AJT/ZQ2o9r34WXvSnKBsqbE0R6TqrYwuK3FxrQaj3hnC+1y
lC7ECmmo3s1XFa6cH84kn53Pwi7QzWh95k9/7Uj85kdDBbTCHnJxkCvdBNnUxvwx
MuI5v9+m5lL2lP21lgaTT718j0Xq2BnLijDvXE93OVlbQCDGTtWJBp6GD0+GI8BJ
YUBsssJgNpCWqnM43ICd2XX867ymQEfIhuiG90MmJcplimlkdSY+iSus8Gh/7R3w
fQ/6VvowKqFAYadj8zLLJNLMIQTffkC+Bf01+qAjV2m0F3TByhLV2+pslo5pFIaI
8enQGcN0vjjPXGeeVHioVBuA0FJHehke8lx5hs5fGXAtUBPOHUR6ZNf26LNrRJ/n
r85nlo3o/OSaGR0+GJn3C22AWidRzFJUxXSQyVE2gnqYfp9kUh7mLNwg0Me7BvdI
mG2dK3nxlLlekmoxImB9Yp8Wfv3ssnKTlW+ygyvYFr8jCe/+2qTbxjipGMFYQqi3
4QdeTzz5drDPE6JFoe2atM9XfMAxVpjEuLbNWpeJNh8f06b03z+uAEMEoDtqrHTS
4FUA3LhDg+0cHNYh/HwBUUzNdnB+CmcXYhO64+YnHMBDfAaxcgEBpzAwn1uzTbJT
nn6Zs0aldlEhvO2Yeqy1YNLxWLbhq6G22wPFUBfWruWaJxzfQ7v9h6pVZomcuOEw
VdvvJ6SJtvgokBGkbZnAugvhGdQK2SMQp7jOdANsEUumfEdUAdO+MXRSlRcf71LW
5tnCzKzXjQdOX964VMiFU3bBrFkMQVQt2G0Q5vj8t+8+XkFTAP++JSNweMFq85rk
2FL8g9ndnBMSoxWQZTx3Af2sIBCd7wV8PeLViLwwn8cn2nWELFVj4obFqHXaCOb1
O3bDuktJ57A0EKrYWfPbcYOq7S5BYYeXc+inigV09lO/UJe4XMjkinTDbH7CBuMI
5mDU2uQrRM4UkWiRdnwPSZZYlLIwVFWq7KlYKS+PqVtN7EcN47tNqvOz5Ihl6d9N
cZ1zn7SJVzpJYerxScyzU5DCBhVhaEzkdv0Iw8WefMBCpS07L8HenaJkpbd9Bcu8
xIz7slbF7GVEopUv/GWqOkVai9BxB7FZZd36JdWnUJkRRjwcPrvWutxCjtW5ijXx
NO3v+rIn4ilUKAixTPo7rSDvpEHt4eluL1p2d4J0Z4P/KyQ4wzyJ02PCdR631y8+
MnrJV7bvkc91s6s1Zo9XPAW/tkdi3f5n3dsJkh47s6KRnt/mYjy945q4AYpRzw+/
RJwPjtf+Ox4lsufCvsleGY+qiZfy4EfOJ0qnUcuNbrcLwgmYzjM5nV11Dkzk1lAp
Vibb0JFVL3Xdv0lH3OI5gJI2NT/FMwgJIW6C8xNnQOZjlpPDFY7LbEGUsU3BSVeq
oSurCuzQP4yphHxo8zdb4t/oPTkxW6aXOsQwQYntw0iKFiQzSPCQsDNoFdSr72m5
M6Kcsp8hIuBkmpO0PWID36543givD2vkZN2SqKRKLTFvTB3MNxzINRC1j3ssvToi
nsRtYYsyNE5s2vZyw7ELdRcwNbNOOEStFww4/tHoKEMMRSSxFicoaVETcFfVQHc4
ldbRENq7E3WhKKEPNh7ArtxtOaFgpT16bnGCylKJS5Qep6jLYP9WQGcQuacbdnJi
YRlVVFVIhAE0+tZ70Zm10Pe958z6mDXeoiIDDbMDOyVKz4MYXE2thJmiKtziV57S
74seVtf2u+R1IdZfPyuHhvtNf5jknBc1ascp0n73h2OWZTQHfdmAqKFb2qOJT1z5
u+Pt4CGpN8PLQr1iR0cTK+vBdKGhfYdDYy6s8CikTjEGAR8Irdc1VbNNDaiwaR/5
GUbYKF0UjibXt9Ri5EaCXODRLB5jDIXsLcHTYd9imCrIYaL4AZAx/HcJLBu0bueg
+GRFNsbD5sifE0JEXIhsnZV/cMR0iebKqZiBkV15M78sNuSUXYGeiKcMCMdUsJMr
J3of1TmZfH9fRA0m5QfrpMQiYqC+qOBygcCenbTzINbqRqZY6jLgEGq+j7zoIS0T
7brgmfjELrGqFcbx/Xwt+eKeK5noMA5DOjPi8YXCsncAhFMsjgh+ZtPRI+9UIgkZ
FjnpFqSahxSQQpOeKobOV7w7g91Ofjndhs5tjn9V15t6J4ADUEHm5M7XBxUGYm1j
cNYhwKBSm1HqCJ1a1syeYnu91PPGvV49DtKi9ymK2Ev81VxwBqHjP6+juZFmSbzt
GOgNhEtDopxy6SDtYnf9i4wnBiqLyeGr8qaVWyAIs+wYSWEFR77kXPdvpnvy865T
67yVpdkKj1ZZanjE+nkHCOk9RuLjY7AHOEuVXobH2vMdM9CyevDgOIMmfh+g3rvZ
oFEFYotxk/HEb9qESEY6EYUAmxuK2Ofr5MuFaT/G6p7IS3LJ22NICuiavujgM/67
f+NCQ8jKmCf0Cm250WZHc/CSCmu2rLOM4C4FmtFl2PaVvRO438S+gYTpW3JF/R+l
XIH2sxmEHYAv+EBlhyjqwbtox77XzQrr/uhzziJRsDLzRsppsd3Ev9stNguDznDd
9Icr5ikkHQjKJkukp51OuyazSlB5ctzknLb0vdMXqDUsaLJSIIHkPv+o7Rs5UXws
FU6Qyw6GcIatYReBzJ3l2YujztGIw9UCcnEO8ltEBPQ2t89EG4ghffcwEG80KDb1
jNxB3RqGNw3AVigkJFy0Hb8tLb9R0qqFBDkqSlLoJQNi1/nkxT/SceAMYuAOZzNi
uprrNkw73lZCWkQ7MT9ueOs4eWcG6GToa+mgRG0HJucUFnyksZdQ9/MYsq5IjN1V
4bmfH7vbxr2DV4+xh5hjZR82MKiNU7paK7dW71dAOxIJU9tCF/nv8R1OzgTTIKCS
YvZ0Kc+FQNmJb0891n3IkEDbQfVN20uwgihL3+TZFWdeQPbuqRP+7tzG4C/QdRtp
iLNcWo23vxlEm43L8cgL6JB617owjEZgP14jvGVdwo5y3DaLDjmxHXVEZxk/+qtb
Aa6v/NjzYdwRRh7lVA+rwo1QCfLQ4ZfeTgLxvwaDoujunC1fIf4LaDRYtqomI8pX
28804BJ5AE+OlTgyb2l8KZF6RO5JY4HtqwS/an60a/iw2X68kY5nMWtSbskWBYgY
KS1hnEE8F2cccyr87lGvGwJKZ44xCyWAbdmfU1+XZZ+F6q8aYCyyqAphlATXuqhn
o4r84uS3prhiGkkl0i2c7omzIZFJPMUHBaM8kW3EDwIA5dmZNv6/CLTSUCqGyxHx
wjiguQJXjDM4I+T5O5ClnuZC3T7tNnfyIxH39sff09TKCg9+R2plNNZwLeLZ3/6H
nbjGDiFMKxAJI67+cjAAcBWuEj/KdsP77xn1RTl4jwWmSybZND2aO+DxGgdKejnz
a25rtLPLfc1IXnLEqoRrsfELby3oROWLKJn1ZX2S2VcqkfQYm5neVZxzQpH5ezS3
cFxMQcgJxsxFHAEIY90Hu0Uf1s3r0ULQIPNrOOXZWTnoPJyR0ubnwdDTyXyurVsS
zw7iVld7W+1WAC/3VIbN/LC7WkYGawRiy+gc+Tx8kYtBtCSpN9gyZQaucLbzDnf8
pVbv4tvJ3t4VChw5L7KIu+PW+yTMm3oJgD8ziT1US0mT4rYWw319QXVlcS9vwXNf
cwePtXMRlOW5Ed+71nACfXhI+pq2Um/IfJ+eEHdzmzdUbYmZrNmJvIlHGy3PwHmC
gz91oxWxL6pXln/A4Dfy1dhEf/jA/ZJBvAeNvMjlkkyW/oYkgGYPcAWTYk7MByWL
iJYNTeGldOp2aS5IWIarrmEKNfPXOqJAtwWkK/z99Xv9X9jFi9Xq/+rvK+rWZkCC
yWOEdetDXVM46WoRlJuRJ1ejH6gkjFcgDn6WIelPaKOqIOeYWpWsUPB72fcJMYZJ
xVHFKUh2wURWixh0wRoC41kAz4C2Z+oU+095GP/kiAKwBYEr80mpZLX+bF2u9hPC
pvMtXJOt4BhJYtaHTV+DK14GM5GVpSsSsQL5yvHLFuIhw+kw/Nhq1xyM2hDpYt5A
5xt535+OOTFB/scGevg9Yvz3vun5704VXyIvq/WtNzx9QcdUhx0Css97nNNNt/XD
zGZBk7FMVnM8xavfycJpAyk16dEmLt+DSf2skCCuvtlTu6AFo0QyjjY38L3Vo3Qs
aQLLxWahqdbT+tVPJfsE1yhObcksGPTbPutzbqRtbGxrB8ybzrKYFrKXX/S/9Mj+
JzNUb44w51KhiBraTwfE3hnZsYZKWZ89ixs87QkJDGHbjfafAwxDkiEhL4LUslJt
c5UkWSCTJKNtTQsNQjN34ODF/MfdrqUXSSCBWikJxK75P++aiR8cXwbj4uE8D8sq
V2p66/GM9Ftlc1r/1TsNfBDvCDDnP1bYOaiX762hVUnYyw3lqPCGilwxGj3V/qtZ
oD6TOiubgbHb8BPSeK4a5JZW5pyWHOUy+eJs3dAI7X+T4N3AWBXD21wxAzn4yww0
h9YW5H36PEsJD1Mvf30zP8KWGR9iikK68hnWR9+wUI4fMKHzOTJf+6QmhtMvI7XU
ULQQsX+LsU321SwkV1xSF7izob7AUf+yQhQIp0eLq6Yn0nXEUFY7YxqASqdUkN1e
kli62kpFE0KzqJxs6N/Q5TPixDyhYfBTFKanMsuWhbtCHI0SxqI93NJTTOTeuN9K
hnLsKJ1QWI2wN2+3rySgVQ70WBzVrHxyZaVdB7e1RTC+h2XODub2X8NmtHFLJbaf
oDbsEOL3H1m0oX7EJWioiTy89jDZ49kWxZgscS7+joS8WQ6R/22lHkMOYIOCylFx
T9Ijj7DifYB6kEEWEMcEUebnKAOef2/ua5129XDhh1uGte2OxoL/Scky4j8ofcN6
OU/y4uxTGWUHs5wiI9vzCMuQnKL1aWuKKt9qZFeg91rE1OcI/Za5+0Ni6mlLa3io
xdG4qx3m+zOozAm+39lrgiZ1ZcdK0ENnxZqn8EvS+9imelkK03mGRCIaEpJZW2wL
+EGBrNjFPbW2hB6g9FqxhSoFb0MgOjFtyfk22UUjGEWQ6Hh3WH4RVYGm88rsLHaA
eKj1szIpUQgA6OSbR0XauqbNMoNDcffiTgl5nqQlwW8aXl6PYJbQ6sqDhOEPRRql
8v9PZdPqiJTrDYOtpX04ousKuo8pdKo2MmsU1WUMQCS2DU5o/R7sGqb1IEaRXY+E
yjAnSI3otKlLL1lk8LMT3NFGj/3XDZCNT+lLkXrKmldnXEwA8yFhxlOThvMRlaWM
l59ceCCfDEWcXHIfWF9GHnjnKM/0VY5467DE8Kb16hyn9AIxHvDwakDNR19x8hWL
xyViBT+gamnwZ8aHZ9BlPJX4yxSQqoMKwuufmHm6sUwaYGjnQeB5RGF5VtTiFHDv
p1nds8Gb0dw9rTAf4HjJJk0X8LhP7fAKEjZvq28t47lgGi6UHFyrdJ8Rgu1YhIaz
l1yM0qvBzKG40AmJfoH94trW19uW6PlM614DAWT/YSH4QUDQP0KVQhaJsD/IlyNF
SJ/KZnZQ60rHuluTCXjp01rVh5t+KdPFkmWPp+mmGEGfy61M35nr6KkQtiVnZOmX
DNcXn3AMKMDCOAME3rhTxruVFnbUUswGUO2bM9QIALQq5QTHNwmUR3GEFCJJ2b75
hlpGlS2X9XOmqNjZfsz1rNV35x1dbx0Aw/pvUs1D0EVbYRB+5llXf8aSOaQ+Ywsp
dIkVA1+B46E8uM/SK5gN3t36erILhnrpmDaR9wTK6Z4DgeRgj9l1yw7xH36490aE
kFwbcg5e7Hgsx5NPfk3WEze7N0Kdc1ZpPr/EaF9ABL/sFeFKdqwfEzMOrogB6HBK
BiMo0vPXugENrAGZYYH3qxWxavFx3oyZqmO6OxP3yHco/DTnBfActexGNeXSHGOC
Vng0/fEpFU3SoK36EAIr1QzLK1FEEhl5D8pi95xTckihrKxeV7HQLqVnHndfm/PJ
zMgSAL+PoLUIxoAsc1uJzwmG3UeYE09+Fh7bpqRoK1/Hg5APKiPtM/C/8nnbuikp
Zkb1bbFtiSQRp04QYPqvTZTKBdvNq5/cpVqiD1dFeeqCdX7Npn8ysS8pTSLqy3t3
oDz7Cmd8QNpfVE7sJ80b9Jynuc6DqdWuJq5OHwW2dCIpDToUtrWpyvp3Z86YK8Gk
dCUOpRwnrDxe6jLvRBqQ7crJEITcH5E8KPb8lZphcKWp6732zmVojBtqWQmn2qNS
+yXWhuUjbQTRBN3fvaSNS6P5Et/lKsnSFNj6EClXJutLYiuqhjPDcqMh28L5osgc
p/LRT7ybtiBE6K3phoKEyOg8J0b6awYTFhHAtiwwGdLakZ02B62/Ckl7Nzm+HMBT
jbIMcO1eQNhazOQxi9ed66WVEouBCb9kZigiEo8Q1DuVR646EMSH2c5lbOKuoivw
8CW7m2qjOh7MXDSFQ6FI1+oH+iXJrnJuwZL1RWBwkurSjs+g3n1NRTH5rU0FYFKd
ods49l8o5NJ1Qw7Nd+3uGAYZMdXL3ROqCIo+f/pknhxxL05h4xxNo1lEqkI0w+JB
MFahf5cSd5PyJ191jO9Zbjw/hHz7WsrEQzGWwlFwwgzGCzgJRcE7wx6tlMQbn9d3
L+fFMxZsDV5nYlg5Tx9FxInKKe0gIXp/jxY/WywmQVGuWYRKzxjWDhMOICiLsu7h
DcG8zTXEMCn7TzedmbdykvaysZDqke2qXRlJ8vqLXb/tvL/IsE3HieVqTaZE51EW
yG4VeKnQsRYTVmnhlXwXSwuygFVI8diLE/0D1JFwzFs4wItca8abXCwuDuWNeUtY
Vv1FOyuTqetxQXZsVE88CyMP4M+G4woN9RI3Qkzo2mO/V4nZ2cu0UYWWL1cHEwRg
kV3xgFniC8LyD6teySTxJ4BYRD+tkLnllHC8G3de0tfUGUGsvam7Hd+u7Lxp1a+8
hp3JL0ZeOjncVMW22SlWRc/0XyDUVbh2+my7apAylP7y2GoKAnSD2PV2fIBzJeye
hw4TYGnjsiCX+2DU73V+xB4VFrz0OfyFtFEAPY5ZV2yRZMnglfpJytWNbLrEjcOL
t9jVjCAufYpFvFQqiGwIY6SNwAtyOzucYe2/dp/wU5XMkHCORCSc3ylL4X46vguz
TvyrC0ovcQH5vlVwpM3nbQdFC7wD5S6OfiLV7xcJseZe/yD2bSpPzu/tbHUGJMT3
XfoK3mj4Mfl34gXJ0Gs1bL0yUoLJIJeO7PzjorH1SFk29K86LQ65CeJPmwNFPgGS
S/f5bt4SMsy7OrkkXn52Dxvmws5XKSGr5u/zKVIWLPT7hRIpOhaM5DSN9F+2231A
qh8w0UT+YOewDkiqNQd8XyjhX3ESsLvdBsE8fkQ2lf9ApyffLL646oJZQ/qYFT/P
nGQB9M8sai1aBu6IcwotA9T3okuh79jCD9O/pcG0FXGtMYRz/FkP3ZQ3ZDdk8fjt
ESswPk39D9NihWwQU3m82/gphhC6WN+hK0VOIx23ilDSfNYxlQeJKis+diQWM0kt
caTl+a2imCSDJ292mahPT0VcvCfq5rt7IRlK8d6VxgqWwW1rv8/OuhWIuKkEABnC
6OswMvroTD1Pn+8huEwILxVXyaSAl5DDhaoM7RQXxv2pUWyl2u+m51ghw0YI3cG4
k48eRQ3BOALgC0nTnVLkqigVW6IeiMhJNqTHvLfzf5LEEgy3t062Z2w7tHPRt86H
XG6RakrNe87DD10SQD0pljpxpInTeiM4/XBpSWrlX16VoTXqAV/4IoNX4mFBNvTg
tVA/4rnpX+I9TowA3A4yGyim0OYzR55hsvYY/jjVo6GeL7JjmGQCtzjSmXIdoaAm
kDB7PFtEDr0GBYkB+MJuo7K0oxrNjtrpzKBMQo0kHEEelsKfgkTDA3GtzQLVErCb
ELCOU/RpSG/RRLr+Ovnh1cNs8oSTspspKz72nFGGnRy//NWgpadMw4xDnG9cDTHt
b8K6sq1Yw0Q6NRfmrvXOF32pvKmhCuVY01tiJKdmWOgEyBWlmVv07NYoeaJc22yN
TWFbBcISb+wQNLZbJrYPmgsKtBypwqKFLOPydDOZp6iiNUwZ6Z++LAdVFPDLhflL
Ym1ZWfvbE0BH6ceHgDYMVYEMZvwUt31tnNnmZchEQbs7eQoafk2iHLJlLTJ7a+bu
aatkjfkuviLvG7TOih27tGeW4UR6sJKboTx85kX8pj0ZURj8y8OFye2/y70aNv7S
5ADZbtNM1KbAfjM7mR8NQNd758v7yTlula9soQO6jZJ6PoUXhlaDTG8DEjxjCKz2
27BpbEnPb13j38wXBpeAHzusu8ONbldIwXzyPGS7cnAjZHxpyKLRv8CBT05FV9EB
vjpaIWvMiNkWr5Lmtyax2XkrHMW1VgzNUZCkZOLjSrVYkwAgTceq9UXqYw9IH2K4
PyuXYCfFcxF4kIgo+P/PJJzrEoAHNkErt3s70onuKut/lGhNP360CNTiLKnXIKAN
1ZyiToRMadGEqao91/+gAYvdZv59/w+t9Vb2sMhN1RPnwRYxYddbq/Rqhq2zIv5X
uBnjQPzA4V/En56xMe1ar0cTJ53uSNCcsCBFALDm1bljFWk19MJn7UEE6DdqZ4Sn
DKzM6qvdG6VBDVufpvXxxYcc78F18TAMFIcduD5aDMZby8ldS8hNuQVOpDyZh9ta
Q3vnt6Pxv82ac72ajJEdSEj0SGBNcXXd0umOkON9OXpT8d28IAqz1jgV2uZdkWfu
hf5xGVaAnG/vkQ1GQgLgzxbUwVEqSq2Dnr0v6oqIPFVlnSTwLkIpUobfK4mdydyK
BWZH3GJ7VkHJuj7onJ1+xDzjGU25n2lNGc3trdJkmY6HWLM5EBRcXz8RRA4a+GB/
MqS9VyQUF0fS1Pax2w83f9sypvBX14WVATtbmUJ8O67n/ZPtKzxZyxKBiaoYcP6D
mPilRpJCTKLvfx0plJ/LqOcUi+SZ5q6L7ydsifHjIk8NIhzRIxEzneheMi3uO8gP
mwwloCSfYU1FvUNKU9Yo3OoacDzayh9aoIDwMyUf4eHITs1AF5FVr0QfXYcfiRNj
18hsuXSoV954xfEBhjjUM+3zejvWM6M/m/cwzIX0ahLgN7niiUklCh9qGP1/JIIx
gCGMEKwU/CFiRLPxUYrAo025dihH/Agykc5B4D3L05lwT8nK+CQz3muoTSJaa69T
0xl+Mic9aCKHzgAOrhoilql4NXJqAbRwD6MQfq6IaOHAOOgucsIPOuj9ZkkwdS5/
Qs02gQbhnYrZ6Vjk6hbr0qL6HUGJiP1fvV9Ryqk95bpp/BbKCZSRrNmyX9PLcAqP
p5jSZ3iVuLp+rc9jW4hRai6AK8oIPsoom5QCVbYNRAVKqggbstjwAdbm4IJAFQ9J
8EniT6A/iaoCwR3ewJJ1Bl/RqWg7kOKF/xeKu6QJZRucRB6vI+9hNf2xi075mo3L
ADnZvZ6CtX52KGt8JHQ82AZO0iBfWac3QDnBmmKPGSCkJgaXEECTe+G1guLgYIMJ
xPtzsMoL/5bqiF5q2Vnj6HPwzS8NF/Os9HMADOrWpTJm28KkmFwOpMEIfYnWkR6S
GgjfJ+EIKSibDreCgbaXBRDxFDOcunZlT53vpWot7dAonCY++xLRanGNnxgIxf5Z
izHekgIc3owPcEHPb686UyVJDog5CrErSTa8+TpF0xChlAyDfQclqNGyx5FtF3Bb
F48rLzIasw1epCvHDBhY7j1ypfXiVVtTaYjmzfp3Sa6EBGv+TlHshOdM3nTm3Bvu
xApc+ubeH7x4pn93CYuv5vDxmxNu4etw1AAsXK1Y6XCoM4Iv9rFSnjungEpyYH5x
97ER4xECn7EmaZUNN1MYl7IF+ycS51xmElnB0Na0Y8uXo8QP9kpivFXVn+en5rUx
C/lemD9vvp3GxIY1qzKQ+7rpFZF9DzRzsPLv/LPZzBm3lcNqYLceGAE7iWAXnTzs
wW8glJ8xzjR3bGMXL4WsBIEEPBY7eEJcWygdLPOuzh9p+3xThpaXkasxq890k4Jy
al2huK/K5uFqMgRgyd+I7hMhx670VPxv6gh75w4cvC/3eCY6zD0nD3pgu7cx7Dkq
EzXNKenW91wL1prA6vicnbPpNHve4oHI65t0FwUJNbrfCBIkHRxUuvGcuwMJxjxu
TaQOQ4vNcXtmcbiNB3syCwlPnzxSDNeoE4XzpB3CofBGFu2zLmQP4aAbHFRE7HyN
1d41zXE2FizP6Tjo9lnATGq+Z/cGr/pWmnuriJnc0symMIwG8fS9fQ45JnW3lLLk
GTbasbqBTGpSNWIZj4pOzZxnI1d1/y6qlZDhT0NJQ3jd01SDkBkz5EwNqA15Awzg
Lc9VmSU3lIKyPzqSg3INgN1sIlI/sqsbKwPzToIVFsp6+VnC3X0khpSCCi/YDbu8
B96RwCUgGJFQSV9rqDsNPVlF97/D1vdMFrRirsJLe1S5VaokzUl6K58SioJUL9cU
hoATWXLUQ3mpNF6pi4e1mhZWl/spEPQFnEDBdgpgejuDvUQOSd47ZUSFyQNuTf6J
dMpCNnOTslDpARH4M/LIjr4qB10ofd9I66HCubV22iwKCd5mqW7K2O7uiUF75V2w
4m55e5bj3oavwtmjhakByGVe1Qmqn4t6t19fZZWDCWYh2e7S9t2tPg2gHNZF76eV
P60YR9BfUonlXtNPNzrcY29W16wGs4sVIH1y61uGUgGKSJ1wY+ohKuI+at/dksiA
6U6ISkyxK7Y1M5Y6gyvm+onrYEQiEtTfyUZkN+v7cf2L9kCkEDUaR4qXMjICq7Pj
kNGSJKsHs28ce9IZpc5MBFRPialho8x5BVX6GZAttjAl4vW/uxzxZB/jaaw9hVPM
AsAVq6YII/6/PRaEeQAsp1wIh2vFvHpw8HUjoLbYoMGSs6ApeedRtCczDm+NaTHS
1CSV9qvmbBT07L5YAwy42v3/G2mAmMtxAuW7wToDDwOeIDLtZqYS6hJiKPiEBa9P
d0lCYbE6FswlaEanizD1SlmSK8bdzRjvBlb6QEwQk1LaEBAo37gFbAanAqDnqb5d
SNdsDOk+KgEW8y6NhpBuaUT5Tlv4xWCr+Mbh5qlWWSV8SwSYjNRa4zTFNYPi1xdy
1y2w5JXZXHKUHORNDHIqe3bL3OP2dGCoIoXDwIClBO+ZKgUD2qh7ZHjipa9Emh67
BSIPWs0y4EQ2D9WS0z/doj5eVwcfHy2tdatEmXh5zB0X5/wzISkqI1QHkju0Wlha
g6A/xyJ7k8Qgnv+QSBA8FSROb3xBbhvIr85dN7/arvZulW1nRcMnidGA2pAt8Sjc
FT8RZBu7DCagL1ORXrhD9qyOnY4LJZOZsYrxW2o7O1Bjt3kUXAzxm9x9pW5W/0RZ
ns1r1kTG0l4J2AVqtAiaM1OHzqUL79sQqFgmMC1EuD+KQvbd+Ln4tqv6GufjRH6P
CFVvbOOeOAms7V1cow17GTjAQxNHzMNaNvJoApbUp2RGGDL2U/3GGpJCKNxsJgEZ
sJ9FMeDu3IeeWZQLUk9dJte+vOFAS/3NrVm9varv98Yt9p0R2siFjF64meranD+T
arFtUi2jjz0cAD8RuMiFeC5bqvxalirndiR9sh5XXw47cik8xohLNTuOw8BP5Hu8
0uoz9frGNvNsOcm/mIIkdb62qV21LMQYc6tTgVgqIXrKTeNvNpxjY0UJ7qQ2PaTr
JNceAfqF+r2O/pg+zLM4JfICC8jLNd1NCjDZE+jVV/3/oB9vXFBtyCcfyMH3GmQS
mSIfjSWmvm4kz2k/NmfjaOcjeV23jiC8LhqooXm6TLME99dTNV0Vh5A65r46zCl3
9GUvoBOPz6YB0Z5JxOD3ZNqXP3GuXUWGbTJkTw6Zxf8pCqvbUAOrIevpFXJ+WHCe
fuFyQSLnJ8AS0XLsdEXsKZ2pPEjSVOHlhs4NRKRhlTegrIwOMU2Xa2kXS83ZHzBe
qyVHVvr/AtIVRenYOz2Q7EYiBwqsQ5LtQs2amI8azk52HO21BkTBfmxwFIKYoOZ0
oYH/EZZ47uRjohd7ubEt+x0jL5mffjBHn9fXxJH2lI+eN6ge71/yYu4FbqmP+IqD
UkY9gBzu8XiF+eobyriYKCwxZnlu4HVQOA45WH2Zvklo5I3eT6Hu4diVLwZ44iRX
6OFzZ/GlDvjO9c6l7jGaGvskXZYXL0MuqTO6FXDjJaBFGtYUTrUQGarHrepGIu0k
7/G0rqYMxvk42lin2JzCuZXPuKF9dKChSGHjs3tPWWVkIxYI0dikpO91MnffdYqD
ds8rpXFJM/Kpt8egJkTpDP7z9l/k4zRZEvZlA/bdtkIw2J/WMaDgVjN6ekPkGhj3
F2W3AVxNceIlfJPIvmOzV/q0s2T9/6T8JA2/4+XfFm7bEi1meD4W02PG+sA+NPWY
uHCPxYNxLCZ2R1vvAslyyz1rFD9m7MOPLVxbCTbK3ruJTFf2JhFcDR8PXg26K6qk
3jFaYH+0bMS1TpUiZ7HrozgCscEE/2k60Gvaw0KjyPPDVvSg/OelM7kueLlGw/A4
fOhDAV4XimLO4q2gKRqwOW2ywN2T4mhDWUzQZEULfwLySZsfzIvyPsLxbzxPaXBk
GoE/w9xTNYAdhk6D+oSs0U6hSzlRliREmETkiret5D56dKrx3NkeuHPR7E6ZPA7n
l5NZB1ZccaquMoLaslX/Je5CqqpS42DL2K/dOZQAZ95k0tOARuYGnblLw9dsPyfV
0vPS9YTVEDeIqv+1WC9yLz2vOowyBoEFX0l3cQClqcqBQ7e9IUrNiu/3bl0vvrHH
/zqX+iXiRYkAwiXFYjZSkSfBwp9xEWq7rVRsC8Li7sjBm0pxQ2Z/0gDdKJTdFyHY
IOyTpKbn2SlWERtcx3qAwyLLc35EbtLrzlVX+5zfHD47/PWs2vv6NabU180pCYOc
KXkDJBRli1QCYFZU/v8e0X0RMkzNmkVixss238jXSyRsqrnBWllHsfr3iAseV5Bz
Xro8SXB81lCjm3sYSv6w03sLBRrZSF5ul/kHd7uYkjduf3icrD9b5sabnMCfIcUR
DthhCewAVGr1etBNGyRVXECWRVW2uSFmcFg8wBD9JoQlQa3fgKDk102km36MTX+2
tiJZnt13EWEch15GeGRG1dPj2ISdFfsj3ltOwd4C3EQrdGsKfL/tzS6jRTUWy/Vp
6TGTT3EBTQ7GLwazm46w9wcEOiM4I3h0/V1koV8wtBXWT778aMT9jVJDV5orIGbd
Ff7EypAX0AZyx3CF4lPWPQ5NxJhxykuGyw3oZC5Z3X/oMVw6Kwaz/OwA5XL4sihd
RZ8K9L/mz97SLi0odlKmMxTmOV1rGOLMwILUjoiLhTzQnrPq+zaTjTkR/c3Wd4EB
vIo0n2qtgNqtTvgzVFqeo1nWePSuUnnbXGLkssLogUcplVSzF8syItcJ3yL2mjYv
yoP8Zpa1qs5Q5zVZ/WgbPPGpzRl2M0J6g8XFBQTxX35DKi5fMdPPm3RyUuRYLh1c
gqdJHOWSis+juUmdms0MDI38HbZqJ9/czR/VFzrGtv2ZvL3horHAssw3h2CPiasq
mjWtY3is/yIYiA7ZaV/xoUea1UZnExtLVGDwdtonWuWGir+Gj+AmsgXYLtjBcX6r
MCMueYaubufD+YXh/JM7wlr8rSSILqaj9CAaazAVNcT5zqP1XHp39FTJUYJmKR1E
vPV+ruQEIa582+uFLrjHWGOrAKsMiNdFS53I0jL8oRmP36q6EDmkosnpR41ITSDu
MVTrxERBPlGpdVY0GGalGiz8W0rU4QnZgu5Fa4q9ChFn4CJeOpaPi/M/dqfTog/N
aqxMx+stwePYrvmcfNHviTjvGDZjMr8Zs91qLllEcdqikjHR7mhd6s+eqBCud53Y
X5OKDDVRLUBQba3cwjyXseQHvygsE20H6dWgvrwpBpJabDja/l0hOthj/ePofh9w
g5nQKKoqlIIdbRi+AhO9w5neAyL3CC4HU6RK2vQLTPa45QZFE/JwwRLg1Wj5kHjT
BwGtetyg3i5Fq6rve+7GDkICS0Mv2nL1Jo7teY9cNLtdQICTM2YLBQqLDtwuveUg
4bPU5BCnJFyr0w8qmv44ohW7y4JQgpOONXmcqImxqInmzKfTn4RLg89kFteFlrot
b6pxAC/jcnXwXMEmoqBYhNyBjtVO+MqLiBpFWNahGwYLWI1xp2HeJOhNnH6ifNXZ
xoAKvrXVm3R0XMMxAj5Uxr/EejyS/oX0McuOGlVaFTHcYiETt35or9iyOKz4CWFq
jZmtE01TD7Oo+XaSAVeEV/fa1sh0bxrbIQ5p0fuzEripLHiKNLqBoVCwgpBoFxHh
5o2Eor7zvMC30QOPYPCb5Q2fnYvdmybPgDobDHaD46jOmviFPz2Xct0qA48HycKG
XW52CZX2cnYH0X0zjXwBjizUCIYsPomQF6V57KZ2QGhvXVar3dCWNq6CYyHPbEWc
4cSjrAlYLHYAIR4Zag9s+rph/G1agQn7flHDF8v9ZmiCyDderrVKGHsDbRUZH6Pi
ch9SvJKGsfuvyDpZvy4NmVWK9h8y1s6jb3DOQCgk86hVQ8M6J4CQxevHqexJvY44
BznS1mzwS7t9LxQTIU2J/CBdfHfYIA7Fpvz7JrwzjeYt2Fw9zSMYWt1er3lh+9CD
wpsm3gorDmPX3vQN7GvRdHcQkQV08LICNOPaUxukYwFYKCeViICIqD0yhj9ySYiP
i/4qmIHZ2IikEdotPG4IebNOx22deuOrlddf51S0C8roNgeEW6czowHwpPiq8rbp
bpMntHvCBk1oMw9ttr/kkdRiHTudsE/Fre2KTOKtVbLRDQFVx7J5z+xZViJR+dkQ
DoTt0rVGrwD1fjI7XJc/vLir8syi2UjuR24jAtyvfCuXwHaRym/eAp2T4L5LoiF5
y/gfaV3nsUQhOHsoZS8tpRMHvyctVz7pl1/D1V5566JUPG/sTFQN4DrE0sHUZRR0
Gpb6WlyEHLNueNgl6B+Arfj22NX/qWzodsF06gxg0pd1bOsOiA8mVwPSzoKNvgdv
0HoWysLG9Zbeyd+aJcqL+eHjeCrqGVNS0iHENDAhCwJKhg8V/IO92C6nY7E9s4UN
YfvsUHASbF/+ZK7RKoeUD8iU/3DGNyqHVZ8B2GWI3MH/RF+OaoilIfcp6eBDSnmv
DTHesaLhvhNaKXw2LQCcpw9ttc9VqoNRr3JYwPQ2jXlYipK8BAnJ5OsjX6IaK/7W
yQUEEuTFxY81VaXpZAkpI29YYQb0nrmQNzI3tNbD9gXppavijAPsrZi1sUfAIxM5
NrqoorXV2dF0K5ZK+v9pZZzstqWE+BZoTMIPLYE7JlDvlrWDREf32RtPjv4aDX63
w4VhZvN5JQobc9D+JUsF9MZwfqE962dwjVPMdsW2lMGkxV6n09aFkjm0YmnXV2VI
vVq6wSvGWUoVDcJdsNuGOQYOMOhbiHdXtS/qT7tfGGmgGqkTurqBWg73ST0NqlyC
et14i/DM3aGG5BuOyTx3Ed7bXRzQg2riMWcXfQJUA6EhEGrtxhBMbLLRyQ6GiDhu
3Z0fq8EfcIKGUoBJZWwmgfBH4DZYs9q98QZbvk3AKqVq6L1eodqF6VDOYlE3u2dq
OU+CRfBzDCpHFX7Oe0PVfSZ6Ed4LfomSXwIPs54vWRVqT+p3mFI+3Gaxr/saIadO
L1vC55ZbXOozWqn4wQNhe+U+mXeVSX9Sl5lbBubgVXDUNsDYcQLFUUpvi4T9OczA
OmiFtwWmAYgeqW5vMORjo8UFw6Rqp+XGO3s/gcsFQbN2YmnS3bbp8q+33xgevm8c
DzwwLAU/1z4Kv8oafNfTCjR+57OACv5GecOYcwwfScqMrALf1Gk80eOK0vghNE+B
c/Pp/Mpb43BB+9mbR9uMzC1Ilq2sPLxORpMWB5AVi3BOnDv+g2SUtl/BFyZHK95E
zGYEATAb84mbEdy3k232nXEX/gznua6K+hKZym8a0c01PECvywD25X5zmqFYxiHU
DHZUwsJITWBOasDf9I11ecauIMmULxeWkm78ShHPJYbdF91Psq3bpfH0cQOozh8w
0+SopDOAWssuBBJ7H6c8sdEV8+u9IEPEJztskUi1GgRJxr9CcD6ToMJGtXw8aQCM
ViDDRNSpMNHewelqfE5O/cyt1xG57MNtfxwBcKsKcDBj/UpaHbdY8/DgqrYwX2WM
NuxHuYxXfNEtwUHhuKr7x18i9JHGticS55d94pUTEhWmC7kmbsAs2zjJcG7vGH1V
dItukwEqhWQrC/T3LrnV2tIIttflEbwkrDqWJlJeFxEu7gCwv0+buY9GAjxsFeZv
natzINdKMs/wzDbQDk2dXXA9bN1ncjf9oeX8sNo6Qpqdr+AIG4GEdAB5f4WbftSZ
5S1rnL1aiIuknowBI3l5NS1SWu5C+YNClKTKV7ErvIFBZwBd3R7jtmYJEtCanK1E
PrhJuH05g7ovA7HwGCjVs4lDyZHAbbKlFO1LjpEjg3H/JjZdxo85FtgDZQh+pMVe
D9bhIyog9UQzWt3Lm5Rjlc6kFm/Y+uP4SCL1yosx3JrAoUnEpYk92Et/YSrHLO4E
nZdSJBLEFjFOQvcQIiZc8xqjapHJVHKtpp0lQvg+DBO/W8Bff3iMmWh5FsqBITxa
iFkBetr+MHuipfnq2PZvF+V+l7DApuN0O3BZRFSVWkISilgV9o4//vg+b1wwPwX2
PjRynlslzyhmieHnbxEI7Gi2JsYunS7JOofczJod0fd/X5FXH9PI6XdcvruEMbYq
CooCgNFNuSKw7MGEQow1MuPcvV15VdwoIn3QHhCpzR3gU7oVf9p89/6Kpsmm/IO7
PfqM00AA84YOA9fumJdbQ7WHZxNzwoGpMPIIlOJiCVIY78jM16RGduFZPBZ98AaF
4rcmpI4s1pBJDbShOCzewQoKiVadBKGC+xI0tEcnau7JJRoC2sAnbkGlrJS5uJl1
Kh+Hoa9zto9zZDXVCTy47txHKbskuRWZcpOgbNwjFDoVXn7Edu6bf8UcJ8Db90uw
FhljmLNqNKQSx16AAoE4L8I7oDTSI1I44pSCv6L/XrOfRvQaqcKnOPmejHDyIOcI
9AvlkrEUAHae6tsgtgfF9RiwtxEvEzA32YhRI7hANFIcXU/XuaowCGt9815h+D05
vaBx+jFZM1Ek37kd1nZLFc/OONPdGShj6Yg5uw2HivGQO2k9Hnj7OToRc2w/W/8X
t/pylQEgTGuAcZ8ODUX2J4iRB/U6EVSkboIYeuLQlIvhoI7BLKIsKofNN45fq9rj
5miWCP/M6yacZRZouCH6s6HaPqUkfb+nVY2tHNPPZ0w5UcVPlr9pK9zRYfz+HxX6
k6X1PniYPvFJGQT2j6yIoLHZqbCPHEsojlaXdFmp9j3uvr3YsQf6vOnz6/A7gzcF
gtcgVCAlx4mLtd0N02B/lA7kFkx6UbEqebMrdE1lM125p0bkJDWuz6bfCoEuO1M+
Q0o1mpCtJ2ETCCWe2VxXO8eELkOeXekpgLTmXFnplMw7nv5hXe+OCtz6xhyBPna/
oI0kwR7Ue7gNq9unxQbTsC/hrP+d3AuqkAl8kMKYYM0X7bnj2oFHd40Rg8jdor9T
8m7sMyKAPDEgnNURTk6qZsvAwjUdXyZFOjBecZgwmIfmFDFiVqiUtxItYyRYX60l
kYDmuuu2sWk4iMYLUabU257cS8xWTvBpabCxDuTeJi1bapV29uCE1zLHUYn2pZxt
5zX0oJpBYWJjDzdnkO2PYvIx0WsZoD6MDZGYabUCzqUkVs8gOpnHL2WbBpGDaMJe
ioWmliTouzGsBAl2xjUnDvOgPKlH7eZ9HB9Dg/F2lSc8bOzYCGbqK55vEA9KzN6+
o13B6etwP82bnfbgbpLm6aUwPK721Qd9UAHwVy8qeCRgKvAe3DCNlTdRwIdUhZU/
uJLJFjvCtQSbHHMKJeYyjNukxIndlqDeiHDqIShz9RBY49SGu/RGWVsy6uSZXAxd
C66HxOo+MZOXV44QFcNOYL7+adUuNkRwxNyL/+Kndfca+qx6++FQc5Kxvda9wW0C
INHPZ8/VVOkB5qHcsUCr8O6TR0R0Z1obtV4f7fvC1pt5cOFCqgSJSp1YsvXhCkWU
eWO2RPg7KUD3KM/fqYgBKH9ImlUVQy8TRO9NAyfCMsn1K/tU9muBsl69286p5fbN
cmZRP5zX6pyM3CO47Ex0L3ozTDYiErzdJg+pgx8a+/2KCuxJnI4zPapxdEVp7gvj
wJ8XCJtVhCcYvSQ1Qq+zMHtOw+RJqCcN5cpat/SnH5BvR8O/b0vbtcuvyOH9I9/W
4j+eTtLaDSzRwfvT3EU9Ykh/HVmXL/sbY6mUnR10Zy3cYev0xbGlES8CsWyGZ3fi
tHvvA4UfeVCLz1duTqAtheV8hCqHPR0jjkgnX8lJG5y9Ce3Tich0ZtjETjoKlwF4
vGJCfhzNQnwuZCnxtHq8uNg0jVMx9mJIvl8PGWTKD9mQTXsQFn6Y1vCAtGHLxvpV
Qc4cpfMg73lXMd9zDVr8qGq2MxuTA+2KBD9pHH5z8/UrlGRvocQZA+zrZbinNh2c
cFXZLImByQCh7YDo6v7aXsZPQ5fFhgB6yBrdin4JZKblcwrIinkPy+psa5Mbj9aQ
/LlmtZ+316DAGbOxfCcP6dCrszr1YNqPQNxx77BfmQ4H2WMCz2+fXcZfyUr40KP+
P/nksu3pJjhkZxnwFObAmfPgl31uExQ168jU3juFKYrNUrSXaJ2RlsrTaOjge60I
FnhlEUMfXc/FdgmDU5EH/o1KIMKt/FU5+dcMG9CuofXWoSb6cv4HIJV9SJRQFLZO
e8hp4CCJ3gVLfa3DTO7tEbD9hm0sKOmgNM0JD7PDvbmG9yGkq4kybGxt4qOs1qwH
+l1abZajvm1tU5LeHTZIchm/r9QPpalAGlVDkzezcYjJPK4dNKNqjeOd69YvCkOh
rrmFVE58rP8D3dZf5IGUlg71L0QkySbiQXC8I4IiHi62VLEO0FOCGQ8vkNHR8daV
o3YAPagvP3+IHSry7drQXxCg7oIG1IUl9rvAgDmuSD4YgFCCoEO0/ito0+5hbtPX
zFbRMd0TWK/Q0IjwrEbVaN4BGb2u6fRVhDrzfOWp67mWAMNGUxbRDJnYJKR7KZ8+
fqxV5UMq0Cz80zWeB0HgioQr3lxwWpGJpCz178tmIRD9WRcBdMdml8j73FZEpCwS
NBkWyXItI6fbiLUgQOYPclqGItQH1RQf43nHDIjOBYv23J7ee8Ep0w4fzVN/adhh
z2ZA1sgp4K+H8FTQJJ/xKgmN00f4+hlH+N6PmK9+Eke9sQxDuxtkjX84+nFgllYi
8Q0evOs1H5DqQME5eb1jVBe7pLo7toLDfDw5T30CopyNsbEWc+The2dndowT39dL
xHSdk67A1Z6ju/GKphX0ghfpORe1+G30CFVdssaLiagT2ZLZnpV20NL+HhIVZLb4
CMerrLaFZxiIQgAB+D2t4gVvPBz7iXeyStlyCRTWTGG6BFfOnSPf+BKijxYy2j20
Pz0zZH+qy2JlYSrTLS+Y7wGD2hDx9eM50friC503p4A1d0zTdbtUGHOoxA3xehkd
Eh5S4fT8aCGfzRIEzH4U8xfKvWxf595zrtmZNMQfizGqJYXj5A8U6ZPZDzzWdCTv
Zs2nk6Ydcn+eGXQIqV9aH85HRY3pQDtQT1/omAJS8eFZldYc49WUQlj6kHWDMUUS
HP5H9GnAk5EG8TItTmNhlB7dPQrz7ohq9RyOMwJVTYvtBS4rew67bNLe0P+uD8O5
WyZhy4gl5njdSAbo50xcCXa0t+yRCKas/tQHN/loQnfcPn0MQhYqrscXNJxrbY2H
MAxaZ1m9/Be3jS0FsuHPkyvnJgvIg1VA23LgCF8+wIeliatE+0PFTaAmUsWyElrd
OALZpE51BSomJHDx2TLmJQhp4FCyShX/dUxpDkiRX3sPN29Knsr/VpPZsUFgIduZ
p1Y5DW40LM7gWBunz2x+7YHqs706N4YB6Qxfs2xI8TpxtW1zxuvSqo7oGLhgdndt
ADXU4Z0v4PXe8e5H9BryNescWKZDfask8qNldBMNrHHhR49Q/g/Qn8tk3tHFEf5x
q8Z1lYlgg+PdXwzGiP+YN/OzWLnY/pRUYmdqNrErD6CiQFLJD6S+H715NHbLcrTV
cJfzClnoz0b1lU2WjgkVpZFWkOCV7eboLRMspvr0DFjXnjT3kaX6mhDOtvPXb2bO
eHw3Ieft8WiOkQXkNiBDYIYJsIuarhtg8kgke8un5nqnWG4qPU27kLGP7Dp6fTzw
Xzlpyxtrbc7C9yQWb718l+8jA9TIhS57tDjcKJscL3UW4vPix62uvvRrrKy/9gzk
0zLf2IxyyjS0IcyLgmU5LrnU5UqSYZJhR6tcB03Tv94t+94p2KkV1BVSYHK2J+FQ
2EmydxUpexrJ9bI/oGMbgu1tEB+IUeiJyWK7CKpnb+37ZHfcQmWe/GtpPQ5t0ObI
2RkAtYSCDrZQP3+0wuQ0V1ETFem0kuceaTgwKFbhcg3og6LUQ/0QeeBHfteD+wyX
H+v94w8epJ9dApuQnzaU+751BE7+S1mAwFF0jHv9ihIi+q0PRGx7fwoiin+WGTo/
j/fZR5Z5r6xmEpS3ShGukF+dlAsykuO8wQYTlyle5adYI5dkKhRqbJC/KQktAY7G
z5r71QS7FP05aWEcVD2VianwCoCdxCuSDqSZKNsAILek+3/3PYQ6IlaWcROD5k4y
7b2KZkM1IzjLBYw6WIWRpcS7osQCYiCsWCM+Gib9G/jtylUwKl80CYTScNmuafdk
9Iz1e6tUh2x+/HaWyu7YXgNA+vYhumZBdL9at0PQxApNWsOW377hncs0X8kfZN8s
ffZoB+uSrHBqwBfSO1RZTUTC6F7h8IEF7lgyepEtL5dEui44CMyEN+ikUdWGAO0V
MFDb6rbI1ycqbzrq3L+umRByi7S1f62IGdPOC4CghVHdvBIAavMuXa/+BcQQlqHO
1RwmdkOSP9dj+CEk6PJVXKbAI9AnGZqOjCr2sRaNCgDBtapmoxYu5MadHfwkjPIF
dmdA/DqhL76+kMu+k0K7+GjBIKLc5MTFMAcZXlNW4tqWseYY1Ub48rqOSuJGvNzK
qwCF3O1ooBmDElt2jAbnHX5uxvfPUW8tfuo74j7+uPf/bEEKeNh166wsvisWaOqc
I07nUz6sQQZtSKE4p02OuRPVJx+XBZzy1b1eSNPSWawzc1ljBExFvrZT3X9W31P8
tHqiyw0CWKiJjxgtsaQg4kK79KtwzjrkpdZbYTXKVgd8wNy2A6WsQ3Bo8jIR8O2D
yvWY/ItMYsQe4TRN9/BDO0CYe5xMhgNchyJKtQABtl81O3lurto8RfbcZkDGJQ12
1r0ZttYN2gtk+8yOgJQWW6TEcebQpAroaQaa/xVvKEHVCbKK5bFdZPYS+EXWj15w
ErXO+bEs2DC+8brgEUgoUIfmPHVX1eEzH4/CFcX2T2t0QODOfLozw2wYDdwngQHy
5sbxT+2/NCInAxCmL7jUS5ui3bLopi0jmHRNRB4yZ/288wA/r5n/gq7BKnJJ0VCT
hw7ie/0QDvr268YfIC3qjDS4d5vw+YOctUdHDpO+GXHgun6Hrl+F+xWgdpikOnbf
0FaVbA017Fw3Jp++gPtwG9Uvyt3KuuXdDhiasb5AdEnjCeDu65yyKpEHYxgK8Qsb
ctx4Mst3Q2svkJDrLCATvw/ghUfOkIizIDwr2dPlTcGpBHQKVUV+rEFHfJigO8r5
N1YFMqKOkLih1IY5N5WSSMiixCjQmpbpjqxn7C8BG4npzhJr036aDPx8EqgZ9N0a
I3IQp6yLkkCBzwXslrs5jzBlkyfegxCzZRyX10Wjd+JVHtt9pRg8VnO6VcrG8gWF
rVQ5+DTjh+ys3o4ROnhJhfwv93ytTXia7dvITA/9xa3H7L2SQoUYQVPMNfmI1Bdw
7y58Q9jZZ9e05SZZFMaYYW4AcJbLPJgMBQFuYiuoT2MgixdXcgudwV8w0vEgN69T
JZanO0u8NGKTUxsxqZsvRdPfPvab8TLoR3Al914zoeZODX78OuoMGINvuamelk9z
3g8KOTRMvoCcq3OiYnzOTMEqB6Jzq81qKQ9oBCFSVqyfQEQPL/3e6JL4VYPYErXn
qLnWgwG3DkCfgkeigb3JpExi6+xIXI+xSx2fRkBgfNUvby0BnOgMGluLL0pytQsF
UcbJUdWR5Fcz4TLUhCbggFHHZhqk1bbhbnoCEaj8zou601PgBpfogSOGMl7KPwBH
fh+B5lftRpEI6NpOrC3XNchVZ1TYACew+TWgKFWL5J6rKyf2HCh0AwjI7j7Osy5X
gtqtHwLRGZ+nP9NksMqc1s4Ir6c59/4zYqtQjqE+QJgs+Sd7LhOKl9J6831Rd6Ix
8THzQPBG67CHFaIxFPvXyimlzOZ7d66aRdmHdk7P5ZuB5GoZ3jfEdQ3PdeVb+4kx
3j3xQaBfPK7RDgb0ESYmxwf9ekizeN7x7a4AZ3RjHCfpc55QCBTriRqSCCHV+pKu
C9hlWLUX+WBm2kb/u4dkDWXiVL8aww6LLZQVEBrEh7Wh6fSRo0O1Afuu4EsC9xVC
MThfMpZOsIMaUMfL76Xse13kds6tA6AVeVUC/7dFIlEn2pRmkSQeFAHrcJLRFdeO
40DA3B+j9+TtvDjtK59PxI7bNDqzcjLMW+DiJt1rsQmSEG35UqqqNmouiVsyGU1/
GimUQF/fyeavt1hdDREFvEFoNo+K4D7/1JemJlImo7dPjOppth60SfQLmMDs2L9Z
YvA91GihUdNd5VM2+TgxKgIc6OC93Iz3N5c+bg2paun9ZqSpv2RPidB8GUbzWZaE
un399nX8QGAYkUXi68ycog0p/y1jC+7lxwFtQ6ge3XFc6xkbD/4tkRKQ8TaoQugM
pO7p1/ZfPgRX8CMJihCj4AlUNmMwzAIBqHGC1H9jiDBAa6ZFdOvG1PHXNAqrLRBO
wLC3nOfusRcjqY7+Jj8pQwMtI//KM8B1y1v5C2FZIwgRIrHp50zU8UHbvuumh/st
Q05Y8qtHh0zZLudUq8m4mrX/XDpyQ4nCAXsEtzzZGU2iJ+zxXbdKU+AvHYw330ur
6qWaaz43neN4cmU/k8KBMdQlA/XlkE4k5S9zzEP6z6oM+NDoR9GxhLCGYFQJIpLw
F7nCckq4vdjUn6J8w7jwCGNxxviqqeehn8qfy5GTHIB6Oh7MMOkcXfURjtu8055k
A8YjbcbX5Y0cs/gqyijTu57e2y0rOjl298PlHnNgUSNFa5P/1VjIr7DUnZLzQIC3
HkraN4CNF1zd/GRjzZfyVaWruw6l9GcCTUSerZuuJxuh9A78JfYQ/OUlvlQ2S+xw
sAx+uNbk2H0bLcGEOiaJAaTo6Z/zm4LT+rR0lSY7H7/g3MlBfYwzotYAgoAck/Mo
7Lmht9MebAOphcPWWnEuLAEbI6fTmNwDuTOgw5fHyVcf88jm721A1WyKp4s9QBZk
lKDWk17yalHDMXC2xxsVbmgG2yy2GUot9fMHQ9BBrW+w0xVLHGdRwCZ/8YVX3OUe
Rt9mBUkxye/fjTFLEFoQPQkgfPriyJiCl0MW7SDogVCHogglWNJ+pbB/HPWCre/X
6p1o7KEvud6mwKbli21vMive9Hyom2B0vb5NCzBhMQ9q6hD46MT99qhHL62SYUJS
MYDliGnpG0OL3PKmSJRyHlWhfPbmJUpHFsuSnKXQACYm10vPcI5U3WD5b0iCDlSY
g4bw3uRNgbQQXE5uZIvWIENJf2e0XZ1iZuBWylJfcqvgOtaYl7n3T5cck5SdlltT
5FPzRvLaCcp1oR29hxRawrnnT0bTqQcu5S/8FHdsH7AAipbL8ul4boAlTX+je2mX
f6uOeI92SsRZq7HDuTkSZ0pYooxLj1F3zfmAdnPsB5VGmO5/yzd3BbHam9+EpBC8
GqoR+XkA2janxDK5lU18UIxTFbHAJ3Txx8bIhtn/TLaYrCWi5dIgpIl3xsi/9hWi
dNbWJ88a8bhPrposcTlxFY9ZHbFkC+/pBSGLL5sDQ6N0qFwCeWK7kO8tMqPvV6SG
b+Kgm6lWMxviBU/kajYpoTAZxSTq34nBEc1JE5ih7hfHb9TJT8+saW9qjfENt41l
T0uozs54RZSUH5/5iHZD1h3Jvj7qIek0jSe+lo/kLq2Lbtzbz0brLTKoNNbqI1il
7JCEBL3Gz1to4YbxGafHMgj9BYeUNSxKPkIudutvovCZV5B1InCL6Jx1qtz34DXj
qnUPuLLPZsmgdRP1NaJF9poMqhf7au02hAr5Fs5PcJi99MCGpoqVbK4C8edNr4EC
tV3zfZjBpyooXsZgZKqgbxQPINioGToWc2jJrZMIbq4PWOBuLGFZFp9Kw2dI0dU0
vmHar35ZQvxqzoT7gPDUxl26p82vg5LjZ0OVXNdXsst9yiobWagwVlEvp4Y3K0Ti
gNnhM8RyU4gO3Y9P9VJDuGwYysdXPpBYIIh7Sx3nlKdmQ79VG5l3OTUw2kSegGzd
JNw2cvfLEsLJ4VoJMuHewFWEsAtKQzoJPtIMeWmWIb15+jJ2Y2KlBMvdzdiVljRv
3C7zawfw4uH1ghl+q8USk6a+fDt+/rOkreiF9sMd5lAEHxzjTdOzLp0GW/E7PtDb
aAV9fL2SWnl4wjjXvDygwdMrIRutLpLCt1JnziQp6dj5N2NKkpclFLN+2Pli1bfi
tVOhkq+UoxAZqaFBBMFf09jyZ58yjHAXaj/VZnCRL8+AAahSQrUiwE/F3MB2f0G4
O4HujgUhAHmeXx30SQnQtJ4QsZ14ccj1CyaWbbZlDf9KXCQPlTw8dWK3vKze3dqt
Ua6Y4RTM5F0yQRvoQHU2bMOP1AHYEUeJB8yD5tuPiq58debWRCvwHBUgTigL/O42
2OC17Z8YU9XR9HC3LRZddfU7+ACmimkjZvu+9/M7rhiiMkhd8eYYyOGxhCHKpelR
OrFwHcYimBj3N7S0FzRc5LGk9nGEIe8jJW+myU0La7812o4XQUHaPr0y1wR/474T
E7451taDgAOFGpXFgP8zztVJplevuebJZy4Xjt3oWw6x+rMY0lKX39WtaVwqB8yc
FYhIMCxZu9Fy2MaEq2tvnMCM5D6HKakq6XPQE70APjqKyUJynrOmpdCGQ1WDEh4R
MsbfxjcYsmSkrYy3RPTndn4sNJm4q2scLe2eAz+30iav2nYAKx2M8yLQLR9aC1VQ
XMl++6ajHiRmM3wrLKOR0e/Le4uCVuUvXlRtG/kSdyFJ3EbwuHJjEH5CTZ4lQXbX
arKtZONHhNyY/H0uaweqbcE9sEzJh1Ob+ZfzHujVUBYxnmf2pPv9D7RLO9VYpoQ4
4rknkEPQ0tHvFVPIzmal+BpHAqOTGaBwtdvDW1MJINc5Te3Mi3leeBdOedfkX6M7
96cMZp/szqD4/gyB1ERYX9qazyAawtIhGyd6JKwRYqa1biEu5WcD/RH4FR23+i+D
A2TtPhHoFs8vHjTzIOJFZSyoOQRJUPdkLgrvy+H0xe7mSLZ/zhRh7JMWshJzFZfQ
XwudRaYrJ09o/qEXnCsO03bRMM8qsTnCZrL3qJOj2X+Y5lNCDCjGo6cSx1hnt45c
MwjBEQb0hN+BU3ph3AgraX0xuI1XD+RDY2X7SsCqrvbCVCjlVXtMZ7TX/ihBfL+B
41nbtMLPCexu/D3pTMDskeJm4TyC/pJvo5xw5979y6pw64pTKXpRaLvnwajIRx3i
VCi3ANP1a9fMKgpWQSrDPiWENMfMk8Fnoh2H0IAc3/l3vgTIK1h+1Fi7APKciIPH
uXdjnUvi+riL14OM0t9l6uoDtJeCR40FagVr70TuqDfyH7MLJ1DeD6qdR3hpC+HJ
a8cg9wx/Tcklnw5OKh8U/j4Dd0kZrmcf53OcJ4aGeTM8ttb/3Ljm5CytAnVzoTRi
+4p5jdsqGU3FA4D0qEELUeVHeL3t9b11r9QmNR9abrIts9OU2fSheiFc8UkthkyI
PkSV6WnqOXso5/IOKHD7rpQ9YzWnq2hyAF7DADDgf3eMw+QoFpKgOXWd/DCSK9YR
SofyS/3pLI/H+hzbzhTrwYm1Ni5Ihc2o/5BNOliHpHnTLpmEFY88xEzrB3nMpKAK
pQo/dm/LSwERTm8f7KSDPUyV3eMY9DPHG3fAVHi1OrF6QCTFM26G2Sr7w2DhKEbd
zL/+nk+ILGkwbseUjInoJP7NMRuvNEfhQbUtMBFIdhW8ORiRsT0RBXT4j3FSVzaR
W0bIXAA7B5aeYtHh73o96qiOCPfmQblRYpxxkvL6KXYSgg8yD5Qp+B9P4PJRFsf5
6iyoDi39muKpPJ7c40w3Ut7OfBly7by84Z5aGobchPWF4Hrsqvh4kBJxUShbnEoH
Q5zyozEk/O+H12Mn1XrVHHwZTXT5TLXQAPz7qMt8vbcZEQbVWOeVkSqanQUY6Ca1
zGXd0+MckT80+qjIzFJCjoyx0fLEEbXdzAQalmiMvoB/wZnDNut0V+SACdprF2EJ
yYAKygCvEooaCDNCWAhiUzTG2Z3d2R2tIEo+AmFb7PsJYA6PtAiC1Oze3Us8GcS+
O2rJ3PYT8Z5PQuyOkBAJOZksN+mZaaZGZGFU6VxG1R/QSH8/GRNqgKBB8T7rP3I5
qfBUed/C5+IcwtkEu6ojz5nL5EqnCDVMgzjNsKh6nfdBh/U9L9BRsy1//HQPFVfd
eSemNpR4hPaql5o+DMNXp/fEqSsLjPrru7cqgRuX4BZny20e7FR/9XH4PbpEzNO+
AMk3rf7Py72n+Mcg1NPWqgxAOMAvwWpoezfIUl3Sa/NGPWMnaciA1LKzADLQnKpS
QlJ6wrjMan9VTYXPu+97Svy+t3dkbnNFzCSChbun06GXGYaJ2otFLuzQIvhj0hkG
2zq+6e9jhRxdVKeCrT10bQ+bKpddc102XZWEGQ5xqQF4NSXa0tYvgD7GM4ek49zV
yi+4XFQbSz9w9oLEo8nOBOtca/GjRmXae2WHT0IUqe+uE/Qq+mTftfjwWDKi9Gjh
r+ZooRmNT1nQbpZxqqGFhi/XFEWtzP+kllOI63lKP0pbjnT7oTVvJj7DCeL8uqfb
3okmNKee2Ij2ylGxMkaLeusO2tYkrnMjbGEKDIJUoTfSE2kYOwsaNtKmLk+OXyw0
X3KUDHu+ire4sfHyuaKE9b2tj66QhxHgmhbJuLxpgiOnNog/UA5yntECXDkjz9yX
jjBxo1WY2n7grDG9Lxz6oXjLFAN7XbTk2zMkBrqVvUGUQQSfvnk5+TmOLv66U7ws
l2yxYaa7o+RK7vHdGLoT9R7kdAZM6tN8sl2m/bqExNS1EP1zx8EebiUohVpCMBqW
6mfLlj/krvM1tr4XI4ArlVm8LZ35IzX7pMHEaAgKxoynEXUv46NJIzRUaZHtpbZd
q/vPYLoRC94mkHnEZxCz4eOGnppv4hiLZioIhtuAYc3xltGJrzbydlW1L8G1HrDC
Smdos+CA4JhQEUYq8eekv19Co77MbbIFTVWsUmzQA/aqJlW6s4KwlgMmnJAg2GjV
OVFAYJfS6o6NWiIr9mu9Cqdy1OL+5sYYf+vWMzQLZBznAk7gwR67Yu3AxjoNa180
NQU77ipMT1Ebjt/ig0RgjDII58pDfOb7jGJTRUL30/p6v7CHRr6DcuhVlMNwyxO6
W52iQoxwzRRraL17azSSncK6UVzkejax6i56QCR7rIk+/gRNtd0FvlWhRksJj4+e
FT64Bf5TvtCAWxFTSdQsXhXyVt35wvTgCLlKIN4FborGBtZJQSOaLFg3XRUAEI5Y
vqwJBehufmlOYNlCb4zIeXDewHwE7ds+cKguxFxor5d/0epchuS6k0NhCNa5m2iI
x5aND536SKR/TVDxjr9inilWmgjhbccYi44zt2SF/CJdDCUBNJoYKBuxcU61+Prs
IBJ575p5e4LXaovfs29KxF9DUQUxJKdVm0VJEAtO6fCa591d3ahGx3Z8aTZ+UU/f
2ZW/lFtfC80d0qhbFMYFiBYDvMoR7zU8oenjIwL4180UfcJFR7+H1kKtNdc0kJL5
2CvqWV4eolv21FshP0gtWq3udOLM7yRVAPkCo7hX8C5CoroeWpga0NiIMZWbWR9c
/IBvtPGTrPAB8hvuBmzLtxpRh3Gqt6ht6jgmM5yo8ZCxCRZHuHUipuKMkSHh/jo8
ZEKGayrIV+/bnN5PsALDm7ZGKPPGAtu2KHQXaxVaUjZ8y3VtAtUPFTRgYVqNkuq4
Uap+jxDImV10J+MCvDHT0s6CfvSbMsiMdy+b7w2b/2nnSMjZ6xc00rg0j2myYyHq
tXhEoil3OjbimnANdfvNtyEaEM0F1VBq8MJ2HwmoU1TbQzyV65DBTEC+XqyfEYth
QTDUNWO0jgSHvJAxq/qhp5ltX7hVXEVmtvuIxEkP+C/621oR2GFrtBKowyh0TiCU
lwoHE5fs2Ez2ZfkLgi8XokFbGXAGa6xt7vu2UbvKw3m8oszDjUwNuZXFFNGMgQ9D
MCLKrvv5AXXwi9W1YFGeeMhMdEESBbbsWx0DQI4Ew4sB129nx2LNoDjmqfj7iqhp
F3eIjAZZXARkudefcTGx4QqoIYbX29sv0+wU6obYkaVcCkJsVkjtovcaRuRlJTgl
i2WMN+Yq/pVQ215S0bKGafytmYFEF+WHvZjlmQiFq4raUY80Ve6D2Y07dv7ulyRh
1lh11jrwzcK3lGeC+1hN1ybWaLY46M3/7YsxU75JJRtmEs1iXWEou4peuq1Ml+Ys
h3dnUtx8BYWkmTtt0TFyum6jxIC0ZrpU8hx+WAvqKFBDNpVLGKFiqrugEXzNZLpd
bFlHgd/BUbYwNsqvoks4mL9iu4epGdFW1SWtUV7ZGVTkoJR2tXUehdl61iRcCMAN
yblytpN9BTupSCMIr6JdZjVIva+AtpArEs6fp4Q+l+uB1CxitCPMPTc18kgre8uX
echLm+AlUk/294zdTtW7VbBwzADdkpKqbLAJu/bkazwYLEmdGMYuGNQ27nakuFhQ
vLLogGtRtRlISq3Ej9hfld+4zaG/IJ29U0iBMa9kpawF7dgGuSIDXvtjnnP/CvUP
oarttsH0r7Cn/toW7/Z4/suX3Z6aLO1sNBTmpk/K8ZvDIPYC2qMDq8HNKTvqVAp1
SIJSvl7zCoXreZYHfjmx6UxHl7Eyd4cy+XKGVfd1rtpYH91KM7HkcS67z3MzQFRA
LV6ymnJkKWx/g2/sn1TzKnRuuMmpfMgyIGSTJlgQl9x8H26pmkOplKUM+C9pbUwY
6ZaQ9inhuxqyu8ASm6PFNwt7zzFVrNKydTPNqWhgxTEh8vnGEcZ+CJMf18CDJW+Z
KMgLuMyGgT58ALOGnpMFjiCtS9Nz0cXgBShukgKfChsbF+Lj2rQcDjYytH9jyL+x
f2KyOZbZ32W5UCVPLaZj2gKKZV5daUgLpa2gdPVFxzjOY+rfgNp8Ai3aJKTX5o1H
7//ncDZdVtDYhc+ab1m56MWvnUn8e/ljiVQh89IWuGCtXME7fCPJ0c1Fw4xeqcNM
k8XHhewDeUOUVuZ1y/wBTqSbS59icjX3/sDr4MapfuWLMQ1S7mip7pTfn/t8Psqd
XR8DBbw60Xuy4zIh7+WDvQkSBHAjLyXgycC8Umq4Epl/8cqD6n2TLgKpjW3NXLZ/
I1zRcS5wKYqb4mkro6VP+uibGS0k4U0lpNdodUdBCVWRO7MTgnNJlCx6C4DxZDZ0
t+GTgBnL3jqple1qa5u2acP38vf4/IKRwl+ZEfXxdlYu7mjtc1NTQJRxpYovuerY
6aT3N4nbG6VXZF92axXOCHzYbaGdn0PRNKkGTnIZDzgWqAsKsTMQhiVwOImzvwET
CTHseeFt0qPYxVrQeszCYsJsTaC3hF8UuDZTecbzhATSjMnu/Gba6oIQmy95xU9I
XxGBNUcCzuKbc3lVf/pmzLNuR5adYCupnCBuozvRXGFCEUr5cuMTSarnukfEQO6X
ExoM+nz+07bfPsZJ1Rp8hV5pByIBCCv9qxtCMMcz66GQMk2JNCe04mWt40Wl4y8p
KYuETlat/MHqXsze/ZgkxlIclrfRWy+npXZ1sL2h97/t4dhT/dGadRUdTvsR+SKd
qCHR9fNrf8iT0wKgYzXbjx4jVqNSBOP661SA0Y1hTlCddxb0S9h9gz7WZ4XYlCOd
DtTW9iOxnUWpLdamPkill8tJWW5in8u8W7NdB1cxhs4kb85z+V7/UY9/WIL1TeSJ
JwyWhwpQp8q/na18rGPmRnhxevcRIQiEAaODjGygAi+rl5v3dIgSsBj1SpBOVVdd
zDWIH2dU8jHkN9VsLyhPpXSeT+bi9OA2k2wPSggpg+8MkhIvfs2nvSrqmJyOlJ6P
gi0wVvFH8AUTD0fBCtQvKKBgBpOzEeM/rxENGHcz64iqmQ+bV2npzCDOPDr2b/vD
f7Bh2nAyQ2b6PCddk2b1OWmMtq+v/XK7bdO/DPKo5LO+yEauJ0VYrEgBPyGuSotY
XXRnXfbNb+TmAc0PzYtgyMnfpgmJ14rAYkXlI0M+d2jKKDo1r23Llrjfr/+KRzLl
y3/IVQwH97fih5PQNTNA+WKw9sQv2FKy2PhgneHnK9NwLuKx1/F381k5ioEkntc3
zCdj1CpsAmFq8ALqlZXKpRFiQtDzmvVf70uAgY6Sf1AQG56LjGiecHK9C4xYWvM7
7HI13Ytu/x7bMigVebFg9HRqHNwK6TFHhJx4n+70TpSbDzhGI8QxgKG+Qc0ow8Yj
8X3G2yXNMrWeXe7GsypxqVAUOjD4uB2C3t1tidNgVHYI6+yeHB/FhGj4h2jv6goU
mWRL5Ao7Yjd/XkkrMza3D0d3ttWEB/HbjCCtl0+0hmZM/epxgeadNKT/pYyE8GSl
L3x6mRPGpi3eMyGZpBuWDpb2MQbIOVZUfYixZHUWG95xg023+zSMhRtMC6DoimTw
WpIwIHI5etcPPIR/KSwX00PDctiTHoCXSzCtWp1gbhxjfifpANcXYLznsPKKUtM9
s5hnzvZEf7Avf0OSOBElMwH9NPTWhwCuFtN/BDyHeTji0z7lVLyp6tvazk2cXioh
mNpZmftoLRFQ2xNzt0RaqsMHovtMbx2CYRAeiEi2uxdhaS63ewDPXZdGVtyKqb8T
EgJaWDgxhA6DlA7bnJbJpXM5FDcHQH/VBmaB1w8LftGwHlCiu7Fmc9Rdg4b164nT
IUwfP0ZKPCuiPePmFHGMeJaJMl8jYRmsSu10C6QxZy1U7J/Qk6CrmyVkvo5raYRh
/M8Lxv+o5LHUqNGHoPPzcfJZxlSagUGRBP2O5IcWY98c5HHETLS0rT8jKCB919g9
wWRlWiAPncZIz+rpfgk76oC8BH/GlFia5lZYadQyo5Vbo1lWBElF3PhgfIHc9n9Q
FV68q1AvqURC6K+VGrBaF+CGkRpUgmdZKDYczClusinKAWHjbhj2irXVhymcSI11
xMpBXX/Idcqpwucz842McKZ3jojxUsRhi0OEi7Z8zloetxoGi1V8a10h3QWHMCFI
fGbzSNISgE+nBJIFWtSL3kJIu7UtTJQ0ckG02K/HOe6nB2ejR+N+m5hqAoYcfsTH
maLmtqnNGEdSfKgWFin2OdRJyn2R4y0KwigQeeQ+XrowJmSY5ewofUkQqyM8Ezr6
GgQmVlz1nDKljOT+kOlxTcXoK2PRo8s2cpYSXDRBzNQtxUqgdgOgW6gk6OEETvF0
vWfpa2mMHMqB+rjwfLVXgNzsYP8zSlQnwv/SolqTKyHfDqeGOhnYJvnWWVGeAp1c
4WuZHqE9PiHoKFOcoZ4Y+sKhY9ArCeQ40faakpUHpc/K/kz34MR0nEJWHUB8hoZ6
vNCIWxheb3IgXttqrcDkabTciYFN09hcfMG9E5UwcK7AadYH7wKDtR0Rb+Njqo1J
xwo7YAqyb7bVTCdxveCK06uv89qCA90JYagbcG95pyP2QYBVf3uVV8COsrASlkVu
TciGAOuDvRQM+YiDKOWHnrU+f/9IYJNT2tdiege2qosBosNa+3ispco7i52ga1AV
G3hL+oxMXLuRLDTEPcjBQjYvNikeSm14oLjrM12+Cu2/+GI0DdAA392nbyq45qmo
CYt3bDqHP58wjCFq1jP4QNw1oDEV9eT6ALcLlItP+ZHBgDxltcVe1WkylF4CwKv6
aGnC1IZf9e2QdFExoZBPwykB/5aWlA6bs0Cal0TpkTg4N6mQtyRzUgnW57hiYtwD
SwRo+jqyR+KT6x2M0YEdUA7se28QgGVoRq9i+rfKqZuSvq8kzIb9cLo6D+wKT44z
YcYA5lsjWwYFYkF+tWGPUanQ2NjlqeSnDVQy0yLunsCaqn1uvLKdmXwNSE5xTc12
UtvS+ibe/oHHwpqrTvQK5rptfD+6EdLSCLIqDkKoHaXTxFyWMpPoWAYbanJ6ycRI
Nu4olD6NDa8bupxDLuNr12AfPBNDWLDerNHfqFYx+ASRdC7aibXjkDeQWPCJgyGz
Go5c4dTaBA86CKYKFd26w5HpZ46RBmoJt6g3CjdqfMNC/nmNLytuwwa2KxYwtl0R
oxdAys2MW2fq6ASZ5dI8xuIu520uCwIzr50xAkQMsWEtmOKX2UdMrrpx0m1vOT9n
wnmgAU0+SLpoN87pHkibkVa86j5r1QAAoI1gYTTQyFUBCltHxDnmfQoA6nLiz0f7
KAj+Sq5Ku6kC10ENlD9hPwHKVoBQ3iU33ePy/OCydH5BgT4QxExYaFSJTRGpehqC
o2m6BevbndtV9hwolxkXXvlZzShDlYFZAs12MOE4BnHN5jmQvk/sOvTE18mo5R4E
dSy3SiVoXNQS6cxuqUFhZLkUGg82bOYd4KcNgfKcN0/pnz8awtFKBKTV5PJgrVNH
5YR2RnVe6GHefDd+hpAgcWSHkTU8C2jXLGx47+JQ0FqcRSmtCT99Rsz9ZW74Wxzx
RTaoS5ui/LvP4ddYYgQrxUpxPTof5cRi20bDAIHDA5DLOTY+xCtDeOwHsgafqYFq
jsb+ja/2SfNUMQdLdyi0+WSBGuOVNOzGh37QJX2QvDubYNB3GzQTS7iuTq6xkQ2d
f1B0o1Nl7lraBOCfwew600trsNpKyBJZ85/v9z2QvMT9kEFHwbbzhJPCFT2bfh9z
PJ4Zm68V5zS+J+nW3fKJJEc3D/bVR6dGglz8/TtIMSLF2r1GFqNlkMn3anOyvotO
fP9RgLee7Gi6suVCUf5ZtZeAlGCWnSBWkcrgjzQMzzCpbLpp4/3DpCgyaM31wS6u
6hZXPRMT05a+YzDdg7rFngpu5khmuXZRAKvbjF9Un13kWnyoYrwgwDTBY+O3VCkx
lcuuI89FlHgnebliURrQNo3Zs2Q7S1q21N+ILlwKWSBvWKbY8JQo+ClPVGl7Q12l
ZhjrIRv0W+MAUU/5Tttl4POa9VZH4XzoZmWqmlAnAAYTfeONxSBU5EFdcYruhsAz
GB0v4a0u6twFr6pS/WchxXk8z9UDs/fEZwcQWOa1aTex53ItV7L/n1779FS3FI/3
Ar7lpsGWs/ufHda0FptYfGDfJXq+pIV5MwoCF+67uSxeIA5Wxkj5Uwz8Jzb7HmEB
rsZbCh6wvdywSB4xcoRIWkKtEkDs2SsmmgJ61QcCes+Bi+Hr9Rwk3qCt96F1Nz5a
0QVAXmp1j5sCE7HkwWu3iYrkm/UKEgpLnepnMCFs6+fIZcI+3/gK7WD9UXaScw/8
Bg6lDfYyAf+zjv9YB7xOM9u6I4QWfMoXvx0GLbKpt8o1bNVi79Xbwr2sBz5Ta4hf
G+tjCaCnOx9NJDo+xSDBvL98MbCcDbOnvoTsGYopRPfd7YlMshtuS2ddR9Ql0PPD
0+z7g/P55N6fCKmJp13NeoxftMkMkMhUDbgLtc79OOmkz01ZeaqGPQSjTKzuSaYV
/DRTwTj8u3DiBjRDxpUhOKGF0Li21d7pAQDaxPbeikKnZMPG/MppshVRoT68XmYe
6FgCXKB5NcpNZ92OBedLiffnjDFM+lcMTPtOFRafpwmytnicTGdvUNU9fhUrrJ3o
Hh+qcgcR3sdZ+JWJLg+Es6nCANV66SgDf+lbReH6sga6nPHkHZS2t11ZnGMkQ8ER
5p62d+QFwWc70YniqQk48SEvUj4gqiWeGhVxvtbAz+7/6NI90AVR6zbk/EJdQsJS
v3qmAfQk2ZJzl378fClXQZhqSrBKokEVWq824hCSg8hB9qMrqk+AjEDi6DgzPwwk
c98BrYyz3YzYs/D/2x0QXE8YB1ts5kra/r1/6dtyVE9K1Ck21wEknAQ/+aiYY6+r
7NHr96v/BU6RD11mK9Wh3cT6zrilnEFZh7+/pxiFFByVwkgHwJBsfOCa/Zk6CWsF
9DzOZO9vMzrTPkzF9KTWCBeSFX1K0YL5o5PwLDDV+hd2VMYpibV5HEa56aunZDEv
hivdp5G5SVzverCsPBZ7KTrlyzgpapoWZCpLOa7N86jTagLkgw/v13aMNv85Eqak
UXvfa5iv4gAtvNQbJnYabRrd4EfKOhtRVYRuu8QSiVT2DFYHZP6zvwIXywcp7eon
k7FMjN5sSig9kt6zyiN8MZ5/E4cfPu9y65j76eb/v+Wt6UrIConp+9b9ipA1VimO
GbQD+k1NpM4l7NTNkbNFtsInEz20xbFlZOphPblpmClQhwzrQARCc1CxE3/2y7XB
KEnr2SkDhpBTn6fEOPQWyB2J+saYAzni0VhvrcEljrK2DKPCvdyhJNcCr+UBDk0b
YbmunBdHpomlVM5RPsyPrA74QctykXWLtmWDhGEiPvBs3Xhom4raoWDM3uIgOt5U
NBgieWVifkjinWHMppSsWz+rL6xnMxNWbFJetMWOLI2AZHkVP88f63owrfVbDSht
hb2xUJWJrvjVCLd8SXfv/gVO/3bWhTcBzVsJBIrOc3dAp/cWo+0YIOB2c/p1VsLj
cyOsAsWTXfjjnCzAyxhKdYrcgrdGOosCgaYDr/lWw4yDv18gz/jfsM6wlfI1sTWN
o2ZUFWT/9fxJ7U9nZnXP28xfKqH0lo2hXpBJZAdNYATajhEplwB7eAOEzXTdwUlq
Kc9Dg54Nm7FzVPSFzPjcXDrlgznF9C+6kms+xDchQqw0ZhJ8hVdmf6XVfAfGpcj4
xycM1hkW0CF0WB9bPODpCGcxEwPgAGlR9xdHbzanUSu5Y5vLl1mXWoJ5Z/RJzd1i
Wl6kLmFbANQDSJDDhLXJ9vl70W3T3cIhX6L9iaAKaNmI7LVZEXrdpjqJjzEK8rUd
Ohzu2b5wBt/B8r7x2eYxcLnu4LnplVchSX1L0i9/qLNSTk2kpnZnQN0JsX24RPy2
lF5NsR/vr5ui6BsWZ0Vy9RuYvoVMVZSpGNHphe2vUzmBVpRhJmL9AJXYrlOahEdi
MEnSuoY2XBFULOzasYMfUk4VxbNFXJ7Pj7nzGDDyiw2t94irnWh01/z3XRJiDwit
ynhTSF6uRRR5A/znbgTeyQlOaavgfEm3RDcEIAdCJ84+2komDLulUDMeF7UD/TOe
QXUWM7C0uoiIdCOQ9zz5M+4Jhco3CAICbeKBF0eh/4FwPlsxZZy6GKGxjWd03wOK
i8PMqlVFj6LJ0cFCJk2o1T1TVA4N4M3Z6/467pUS05RTT4V0IyQIzri8Ew6cjTPS
wuNcLUnoIOkaULoQUftUG0xmInH+L6VsTQlVrmXBeC4mdS0RzdlPvViAwdjaSiNr
Y3do2P7AzxdECammNl3G4o0+um5XwaReQCEdIfLZ2NhWqfIt3ZT/DUVaiDdSW3LK
P79bx0VsAtmNMCCwQz65FeYFSA7VpP56XXv72iXWAPoNUh3CHKdqvqfJUrZmMi47
JlOgbuNYA/cXsMBnquPm93Z6FXtkcTZNfkm1j1dlERq7CXW4EiOvPJSerI2aYe+w
CBXD7OUstwUuozktl1kh3MScFKCzDFMBXFDAflUNg0Z2zGH6oiSdHNw6qzPSCZai
FVUHLQdhskttlMXov2rX/UrHxT9S0k4y9NulKZtAj2J6yxwomLg7PeyuDlnw1jV2
DuOF4g4qo1oMsjAom6FZ9yHtDOBxPhruji25yGmt0MN59vJGZI9nPrB8aIGSoDsU
zl6xQqWQH5HoJbqtlDZxkDz2jKI5vKXk/tqGklSH196uO7vTan3F3VhilekjCUrN
MT3Iv/3aAPki0y9A346yvEeEFSWiQmLwCE5jAdgu1dL6EtTfYaH7ZXuEZvJmDXq4
3pWVsv9AjgmQxm2NxgdluJgl3RXFiAGpf+eHRTvqW0j985b6EdWNAzrUGpf29sJ9
ntr482bc4vJXZta1sdtp02luj4hwy0F/yN+0O9FtajEkWwyBQs6pTUZvKw1mGaOT
M8XCtXZ0g8zxGV/P/QTNJ/kkiHRx3fq0AI0Wi8MFO7hrj67vL3yAuiFUkqf0zlJs
nUJAsfaMSoYIjGeFYi44mj1rKl3vct8CXCQEHsYwLNCjesiC9hAwV/sH2qq2i4L2
DcjWbK//cw8VfhxrmInyUUl+CzvFW4iOkYKP6B7ou8HEG08Q9TfZkg7f5wIaLHVO
we0tLPnhzozOEiHloldLLX3XqADOyEjT7QXvk/CW37bQyouETsNKQLCbAu4+iS0E
9bwd7WebZjFY8s64kBTmW06UcXDla4sq4ksdkjArs9VnqicBpoLYUjSr7CzX+mzh
ehoN3A2H2G4ahmdq05O6onFbIwQvY+Nf5W6HsI4iWF7nJ9GR7Y/Lkt42rbS30vfd
HMqvXQraTPk9zQLpx1rVA7N0RfyrmDwggpvl8sPV6GQWHI8o1rNSsLXhy7ACyHo7
3Z2Ug1zGC505anUQltY9h+FIZY20PElIOsip9uguomTqCwhjAcuijGN5PF89KlAD
vQ2xPM5D4OnomeaDlDDiQr3YonALdX6c54MfOqyTici/nNGqyCBvm60/9iYw9IbU
+l9+EEnN55Wyoq/3XDwyl+cW2qyQd/pINltVTse7qeVZLWMKshWy5SnVj+zqAO3q
5HJaizTmXkfR0vKpT9n8fQjMxrcAptCKnyW2jjwwBxILDnBkyUxkKnzBM2/tgTVV
6blrec3mEqkEJ7qg5cQBNBwmlIw6g539ILcVW9AGPnAjH36GaS1/qrxWkF3txKVx
s5oTlVvqa8u8qbsi2V5UnevFoJ/vkAjwOFDMQib8aL6zo9fAN0tg05Vk5KXk9zt6
lX/AnHXZD9GYgVo9PX1GgqZfgB8xr01iFzR3eqeJWkMNzW4s2AusDA8/4VmGypQY
nioaXZfDtxtRqatvZJoHHcQtwzxMlatMGZVg/UOr7eG++N1y19rznKWKaAJx0Q1I
VHMwgB3HisCKvlYaHebi6rfDRD1ikYi2n4fpacfWQdY7nfSHq0WLblw3B4gnwftu
UuPqTtxX2eqylBMQkDc0VjJBzbHNUjofKdQplNyehYeyONZuekFXcoExSyG4xE4E
ImX9CARJZFVLYwEvvscaxqJQ8lf/K+PkEfXf/gUatT0oIue+W5iX6w3A/MWpgWz6
Ph9bhC2azwhv7ZszwLsR9EdC5ARn/C5rpE5zHieRo7vCbv8AD1EfAvo6uK8WiEET
uEcWaLeGgwgW1tztNsbgsF/WhIXzdLRtW2E58avQmJwfCpqs9cYIcMPk02Mt0d7P
FbijyDg7fIgHjLJvdBYEzgzkc9KRW+pzOLVl9M5RXnKbNbnfY3hPt6+OaeRKAGDc
onF9LuchseRktlNjI1VoWECeyk3R3JGp2oPKM4ti39JThG3kIMiKCIOn2CDDsEyX
iy9rh5bIrIA/3t3dzPX60SbYB+Gf1pJZhAOXOUEBuI/aBaOY4G3ZcDOAX7dd/OVG
Po5Y7C9KA6OvjpszoBuam9hzS6de1MbNUoscwN2E5NjmaHZsWaV3KxA9xM1/GCAs
yARxeZ+9LyX5qUAcJBuUtFddt1VfZVYTzUiYJikb8LeEYOnjQ2M2lbl5BdrH0OZI
zBNoMseyICHFeDzxpZ8UnfWYQNJZzl0wJsy3bCkx1c82LREVoBO9e/Eysf//plHn
MDBjpSl2awWJCEpn7iYIMpZb9io4BJ0zZr2mC8FKsR4UKJdH6j9NfLtSMM9kxVlU
w3VQFsO6AaXCN//HZ0YFBrzGJQ0eO60nQG9gNP7XzXLrq2Vj9S3pZ8u82+JpYCin
70A2ZpkDZGQtyjVkF021ZDEk/w9MUasnwRq+EeLGByN4WAB5crapj/Lb7thZNIlF
6Q4KpSO34oCa6m48z/Bh00OOntRv8l0PuFF8ROvU+49hUTEzVlHpMWt4MWpjicQz
LQrEPbj9U8KoYpndLehvXB37Pqq3Tak2MfliXKYU/1XMTFCs9w0kGX2PsobWWdyI
4wC4QewwhR/GX5dNUXTjdRUUV/ElbAnhoa+N+xwM0ka5xW5NiGecLDQVWmbK+VVD
5dQ+4R24JLYh6ZZ+Kcz9el/t9xC/vcakXuVIApseOoDEA3MUbRqyQ5esKWUQ+kVF
JdjUgAYTSe+4loLVCV5wIWvc6JMJnjGvC4CB7w5FlWgHyNtwgmjuKCnjBN/xhJAl
irUAHDCDAvDxiWtz5+CDOPuU+MfEa7qVUjN0sWZfPW+OpksvYSjvvTQDemleM4Gn
vF+uSpVydxFF/Ktn5AIwqtrt3pWMYr01mp59FroyOyJaZ3PPdCnx5MbO9MSjXIzN
dRNafe2SsRYGF94lyyd5+Npz6UhX7jjUhxG3KuS5oD57wk45A+r+1rLNsdyOt4e/
tzJ6N/z4jpboP+Gr4ICYHoxw3+sw8AeCWtOR3kfqBpdgkSGnscsDeqDQ+jNNaQg4
o2y1FtTMpwXE5eygwtIMzYHrb2vjmxNZWoCz6LKsF7gWkJN1u0B2JHBESkkucYkb
1mQaDGO+SHj0Bt7IpFOoSofhSpnEmw6Z1d+c9b4j1FM9DcvbFSpaDlpwrqIRJ6mt
/ge5+fSZgJZe6KAudzrQgioJ4t07e9YVz6hy4nniaOtIhJc88Ig44ki4rrmQUyrB
ox4SVBXTC7+qSQ68AMVKPz2YfRLAgDANeWCgtRC3cq8Q9TBFVMuRc8vPAa/155Lj
Zie8GppG0Duq/dkPgUxWBMWbbURK8XhxXSycEMNGPIEJlwUkuOv68wdLq965PnqZ
59oyEzGfDoOzYt59POmVrGJfQcqwlrEDWZ68wgAWI8RsN29fiTGfnfbIN9E86hz3
WJwUDiyCbTCGXVJgkDmFjUCw2GgwAx8y8PrrKxYTwGHjVszcwZb3CcwXcHWP0C1k
C62jB8LIuuk3YzedhDchHloQRKKbVL5XXR0UuUFmGTNHcg8g0DdJ6HrBe23wpb6U
9ThNN5KZ4WhnryCcOvJmQTJEk6WUI03raWX3kpGysWu/x4MNnetjfDZikfpvCAQf
IOfQXY4ugBT6e9oaAHEjEPXTFEsw9JajUy0iAK0wziSzToM+2WPgXmm7sTkXHCys
dla/i7X/739WwWgzfXHG0zW2ULMYVdGQX5J/qj5E7nevtp4SY816XeLB7LK7N9P2
bFl1Bl7NB/S5FVrXWJDTcE8IlF1j4ETumBv2ys7ZQ1oELKGrI4DDl3cm/SuKIZJa
DqAcSr4e7o5jiqhoaBS1eNRncArgGUK3sj3CDf/V3A+X3KItehzb8qA50bW8qSMy
4VBNFoiXyYtOy5xaoZYr+u82NveLSJUC931Np5+4jYgd3L2IB9bkmfJq0fqAmov+
WbToR4wbdBUj1NKUaXoBcLj5sCwGKjOTL7eEnO64MuS3kZN9urXKg2W1n+GSo05m
KWIQ3pHWLUEOjWSGnIz6iF6EvkD3okr2NNXDFJBp3k2Avcd4YMuIzmnzbT8YlDQI
AYniGSuKWcGckjYKeBtsRPBBWrvIM26vIf7fh+uyoxppALX1+cLDd/eXLeVYh/ad
jDHpozSmQu6u64y/TUnwfB5YHFOx+dEvF6A3aINXddjN54RiiFJkLf2k6CmslyvF
hPNWeiC30P2FNCrlP6d7SE+FJ3QGGZEZA7eNghkHB6gkU0Yx9+Vxif7pqz9+0s3a
eJZevq3UkCiBgRSCpAQur0ZUDA1Wvk1qy39yfOfHpqKQjpA+9FhMO7i6L92T90f3
RxfNtBMuvQBrL7julsxqzplDuC1hAMY2YjnQ5xmftcWNUbD7N5sjcj0ttSEpkgNo
uxvP+pZe9csLLTc9KjQ+dgfCHHFhRJ6fQ7j9fCnyadQFkvmkpqnHiPr5T8QanuYI
Kh7jKE6xx/I46FTU/nate9QGUQNxJnu98SiocbCLOTJ2XCswsCzJwQCu/Fscph1e
6rlVfYNnu6JYI8KhwNCL5pdpWAPW5I+x8tJrSHEjknuUob7Yo/9n9ouNXIIckyjh
c7IkLRBzUpayxsWVKnxPaMFSOX9HYOw4Cf0MKNXCy4VLm7UQntG0mgE+ZneSaKg/
Q63H66DM2K0kFmVyhHNev3khusNl3qnre2XEucTcZAfqQr9WWpcsYwMd2n2tXuY0
EVYLKDtzcxJJoCxxADAKHjaxhMMdVt+TFauucSmdf1/553YBQcGeP1w9t6xAVOn7
IZn5EuB4qXW9FuwALO/rTbUqKgKPwEl83Xiw6sWlTo3fwNJN3kpgsNxyLTddTwvg
WkWBdYOE6RdHV1sD7IvYwr9sA5BOOamOOgBh9M+yuR1uKE4vm2iT1XUZ5cRtgOl9
mar6QMlgiwLcL8KcMxQNdraEF/23bQoJOfic4HupqpvFykFyX0NErwDm9DvRC2pw
1FYxlOega66Fi7fmIjc908gN4QAbxBPkzxKGECtIZjT5LEa/g3afmA7/SooLqdje
ifAbaL9gO7kb5OQbPkjZdTZFGEZDWCP9ACjd2i48ftfbOTdzgoKlI51jz2g7kRpI
Xj5/yxy9VFd0bu+dvAaPQfQ7NkQldp56Y/XspaQk8sliGxQquYGgA5A0w79DziG3
3cM3gJMGZ4kbIJ8EP8af3hUgnVxvEkOKBhgENbkUiktVjWtipKRZwBlQL9GrCTTM
L/ONsuiYsthIwanLxAqCi8nUkun1Sehnx2M2um18ccW/PNeTQ9RbUzYX5LqXQ2il
GUdNCoNVYf4Em39UIhYP8w/D565Gi45Gm3QuEKYzI1R6XJIlRHnJb/LRVQbr/p05
htqWz8PiDDx/zaV2TtxzLBiEsncTl9PrP1fJthYg3DRIpWaZhbFZ59Xg5NDGhEef
PE38ALeoeVsRqBSZTwAaJ2kJbC+/BlW8gs/oCA3s9RcFE5/FU7sq3MYHX4SbweQ4
jkH+z7uu00CX6RoD7PrwHKDlGtq1Fy73yPL7hHqeppNObKXmUfZPvqgE3eeTmVoz
07DmdD69PVK6v+Mb53/mdTlyjrp6b0USpbsRXjaoggLZQHTWkEMz6C05M6v4+TTy
HjwDbqzbGySVSo/jpQy3Knb3GoIDjRUZOjzvgpOtDvg3DPzasmRtwnGRa2vQrKQM
6lcLDibPjLZyIShMvOJtqRF4XD4VEh4m787TZRyEXkRl0/S+QLVkb7h4u3NyTX9m
15V1HiNM08w061WsQBdGqhZfVa1UFxtwGuhGWahrM1MlT5YnHne6ToPLBJ4sojXi
5YD9QjGIJg3OiSqCNLbMou4us3LGQwbeptOjG7TlffdITNSAMCvGk/cVthpe7n+K
w2s/a3kJsmEbgt4eWF4x1M4vCmUsd/qgOHK9aSU5wcT4Wz9dv2kI0E9ZDtK6G3G8
urPUQEYDDM+WtFeDX3savx6opSJhF2o2eQHle5pyjmHyKzB9UkgaWRoXCFpSTPms
U/3jEwqtM/FGwge22IFVW7xkO5kKrNFsWQnv+WZb486ZA3LnIAVrwXUD5Q9dWxUk
RESLWfnGUnZCnYlmi9CDRXJCCUVYmo2Bfg1X0EHysk9T30jWbun2qlJCO25XfKke
P5c6KIWqOsaEe0PgbQoi3bphzTYQLvBsr5zdybfjwuixcCm3o2OQYvNEreNuLxoh
F5NWVknFvudz8D/5KiWu3cOMbW8sLR3+awADiiVZ6ahicJSifwuHgjOsTo8wQdMO
ZsNM5iEDmmf+9dr8CA5TfD+KZt2Yq98K0/xw/Yf2ETbVF4j99mER34mpPRX7Iee5
H5hfJcvT1dD15mpzRCMhY1Wsewe5C8jWXk8FlTQGtYYZ0wVA+NmWAnJqA5/YmTof
O3UcZ6ZIH0GtIasxYfpGJ28DV4zQAmPzarbqh0IjWoR+uCf9j5IYBbR8+yRLSF0C
NLi2eS+X+R1I5Qh6BF5IE3lMM4DTgxirw8txaN1gJS5r+Vl5yN5K4LxdjBST2TJX
qcX7RwTODcEymT3jn4DFDyCQaDv53l3LtmZ5Y8T7+t0HcIZpK+efTyefaAY3b2gg
7QSCruqDXwuPH0oAxJ28r+Xbpm04u8WAXWtGMq+nLkUjOdkb2P2FmX/EoZ/+ctR0
/WrTJPxPa3LCa5x7fm3xpzwjkz7Ykk7aghmzE9l1gxO9A5I/0PiSqBt+b6Wy2oFG
k9UGaNiAztEW7BB/serFVNwou6wL8LFmFHgt2/8u8kwgQnhMqlLSGoYl/2bn8LtA
QhZ/RYqhLWiEVjXI8GPmjv+W8ipu0UKCa5XSt3mVHaA2DGR5GvSkhFAq5jGbqP99
xylr0yYP4fr5rLZP6j8+EYaVgdUmCCzYf0pn6gDcnP6Bbf4J+mjDntaMlNVTsJNf
D5X4z1cqCOZLc+N2MEgYev55dBqPTi9Wtxs9R1c4O/1xPH7ih0SqtWjUjCIzIxMs
c+7FXDEoxpfut+ySm6KdLA5UzexY/3NGxKDAfmY3ERstdiH9KxbB+Iv3O3a1yZQF
tc7s3r4j3txPiCV6lXiZWPChNCx9yUpcBl23ZZ2FkncQNNU1n9I29MbDZ1doZNXk
OqVNxlAXcRX8mn7p0KLMfQhbmChSSM57NFFyhmkRIjMG6UN/cLDbkIDTSSFnldag
Z10Bmu2OH/6nXk6zj4UB9d/Nwj3m2ryXuDdzDogG/jd6k4T0xYoKqq2WMuobonbn
1ZZ1YRmxBNBIFIkkv6Tj/LDgrcFvrX/8GGyWnBbPlcwU5DeFZWVg4NC6H2Dx4tc2
tV/wi93d/lfZl94k1ngPX0lkHaXnHoi1JWC4gY9yoTPZVjWh51UDvUAUvaCbvzRy
qljamkHiGGyhUIQQS0/vDLYHD/bzPKk5Ebe49a42KEx36mZXUzSWmbBR1LuAUYsS
jaC4Y/jMsQoSJVqyuVzvfZSMgiRpwUbQ5sdodmGgokhzVzpWIycNhs1djZtKrm2p
VizEF44ItHJHAFdGoCRPsuKb9FHKhhgXmaMWX6NbGBzJOPlJGy9/qgRF1PNHQDMk
Yc2ATP8pNNrGUOwmtznQy2eFrZ1ElJ2gmcH2tZaaYcZ/tYq8qP1DycRwRIRid8j5
atRTD6i5eFVMNTm0K8yqOBASKQV5qwbYWAdz73j9JDzPUz/7VuT/Fzl3L0K8ePXo
yLe1js+63xBIazQdqJ1Hy76eWM5RjEmy3fHlDbL8PsjAJbxpFzVy0zmHnKKSL5kk
6XM6zDvPaCuoWKJW2V6SlvlpJ0ZOY1FERzX/nfrZ3FpCsoeKpVsAIoC5MyylbszF
v61QTWZyqcY/Ws0f2ZVnjh7xkHn30rpps0xKQGJVL099DF7p4hi4N3GE9JOhFED1
LWRwuledIJvlsIdf0sOVxb7uaqvUbwlBIs3FKRg6eGnvUNFUjUkCQWlTOf6/c4aH
QxCSQmGlLxvV6vdmM8ZhZZBpzOhYT2ORJrB6dR7gZcljxiIg/33eLAkO0Zz8KF+l
dk8k81J6nyzE4S+1xUFftBa2JbjsMEBNyLY+WkftrLzWNp6t+Vy0iZ9/4P2S2jlP
pY1J3qkymiP9JGC+J7dL2tz/L+5JX329ngj+wdkQXmuaWT5BwqJnAquSU638XVQZ
NEwKP0XHwdLLUaJBHkQon/kZyCA2CL5Wy9q71mx+8H7YNJmZWK8MfaLtvrn+jyaB
ywbXq0sReudntQOsQ+nAnIZHFMMrqQr7nIz0NjciKRmKfvbvQt56Tg8ifpJcR5xy
e4LXZc9kiw5Dy4MyjVUKDdsy2NKK7rGaF6ZvcESZwr8JpcxgiyGn0iKwR3O2ozYM
1Ztq7unNjse6ya+kQr6QvzoqR0qifYJ0fEYepgZX4v7N0a2XbJZDrVI9JEzN23l8
+KyKraDo755OBOOca1spfiGDwFnCYLBv5MLQZh+DINA/8QvVsz1i2tQaEElzdHrd
z5L/nYXmL8xZWQWZTZ7WX5klmlEm8TqN9srqZrLr7VDdlhTAHDtIaI8TdmLd8N0r
3PFpCOdnLLKajYAEssAVJEsoHyo4FLs9VV2/6C49P6jaZfSNNa1pxT0RtSku/q8a
Gwt2yjIytBYhB8nh74Y6vds2b/Aom7YeIyQUd3+ZqbHPhOfMPp+68sPVmdJjVx1s
B0W5kpdCeT0lPMbd6VGqAmpCNm8PZygB23QEAdoqz88yRvMEevuijWeBxJd32Ma0
SpVxJjBCHSLsyeCg2fPSxamULqEfeqHs0o3vjs/ZZySj8/w5hcyb0k9vZgmTrHBO
4s9m0orGDu5JQdOHBx0uv1/eUNxpeQAeyaQ951ZB++vExaMekmlb+U/XRVqmoJLM
jb/9b+EE64GTZSHrWucTEI6nppoDIGbEzq2EyhCLroHhPLD8iN8gCzszasnM4RkC
vYM+rlZBCikBtJK+1Wb2wpYQuRnbPbd36/fb7xCLOTskDwDZP4Y+j+zEPN2vU6ay
dUkeZq6nrA6fikaM3MGNPPBdK00EBkPu0kRxNYi3JXSP5QT1R0RMdBdWYjZhpNMJ
OYt+lJ5OJU0SdY0WP8Zqljmgjf1VuFeiREaFFGBhPXhsXUDtxbiidUQlJdnso9r2
8JyMtQCS6SdK1ig/GhJM9C6z6OncnV9XLIXMpcwAX06i0S3SsShLYFU7b3yMDFYB
5g9gbYfdVuHRWpnZt8GC7xyQ3N1klZsx5ce91uT7qIf2Bhcv0+eSQU14IJuz/fZB
UI+vlOP2f3s9JoK7r7QtkFJIYA8MVRj++dA/peQy8iOcpOAL6GUjRXas4sMxddkG
Uc/ao1YFf1JqxQcK4afE+MU7A+NOoXeZEJQuY4xHDt690ZZBEAto7cu9AO44/YRO
hR6GSBONrsidjyJzAcJtrr5aOzndZisu/eEShy0I1YMhZ5fXvVCfPYdFA8Lb3Ore
8DTQUgOhwDeQvDpl6UNKspIJancBmGYA+MkNikvj4VwcDw0VwUTiHXeAt1OlKAbu
74uvwOy2jR9hoQUr1fiFrb9XCpqtKEA39L5qrIMb9lfil039axdeD7oTAoKBtSGf
EJXmuh6tBgqmrZzQVvQ81skNJmC/KimaCr7ihNaZXqH0TH9lly4upxxR133JEtl0
oqKmXNwSi9sFKyFOHL4hASnqRs7CfncdtmIamfpAOD3NArrSKXTxOnSjoJI71zyY
PHFLL74Mzjz+b88IlGRvus9DP6dDN8juHO1K+JMthG5t0qT7VJPRFW2deACOKMye
70dobfBpIqnvKaRITkHG+j9h2VsaftJvr4in5ll5DYeAEfJ3FJpucj+yH+Wm+u9v
LbBIiOLsgQwK6HUWziw+EzaHxMsdxVk1HtJW30nccRz+MaKYHkWPN7nzzBE3+4fr
J9bRjKq4ZXYcc1bKzQcgqh4kkuFHnMXvyTbvCA3HlHhI7B6qcxLFkpybT9qfIK+U
lD0Rb8TRlrG1WWxob7s0GtgC0ptiOPtT5P4Jj0A5ChTZ0Mm1++k/dZTXVHCLbohJ
B1R5tLsI/saZwe7ABCtezK1M+PninVGHOSiRyG71eUK11P+/aMD+HRCctl9P3Vyd
OhijBws5M3Wi5NOgOQgkKnhieKmSiPDExnQxkBto6Cy7xX6fWbBWCB2cO6Rz2TZJ
Zvhk8JvCwWVaFM7V4RFailqQEsoWqwtzO1PxHen1xla3q0AdlY0yWBs9+Y9dXZXS
t+aw35YahUMbzQSkiBNyg4bgTeOxiZS6fsWFTvjwi24xZz/+j52r6BKFUgiKuGX0
MiGX/7Y1OMcS/WGGMvnYslaHkXWkwN/GurseAROsJ7niE+S2MtBbWI+J5Y2MGhw1
ngt3y/KXesPeeE+7xntnEsaqOrgf/3sG2P3YhZeRKJ0TJNedDzQJ+7S1Xaeh9gDX
npDiB4HH5KxVZZ0L3b+X2hJyNpmGal36PSmZeKIPqE41muR8G9NzI6PIXipFbJ3n
0+/I1NZNU9rE7lUPuACz22il/FUnTYOWDDvlUTKNhHHKx6lG6NEZz5jJftSEIFOn
0jmJyD2jKq11EpdYtO/3PdZDKcdD9M8GUMrma+efjPUG4EReD9ToZlMkQD5lcB4d
QVvbxLfLMwHObXqrUblPNX7623w28WNjOIir2bEW+pWTfJrrj0k+YKhkeUSaKi+f
uTmexbSZiUB2gmZkt4GoT7YER66bOxXJ9ho45OmBxgC6OfPnlH/O3QN9u17m/HP/
oQMFi4io9auW11ezWMlYkMXPjSb9Z35X4CzFbUbZJtLUtyinGDOEjWTF2dY7GXub
YzP7Vy2eg8YKR4fGN+Tu6kZbU+dVNKfpoI8tL1yP7KFcvdGyJLyb0psN6BMb7Acr
uM6pOiJ1R1ez/ib9+4ZIdrg1LluhJvlBzdc5AcIq1zED75tIrHPLXhRWr91QXhf9
9xj6LkFxon8VZo4JTvsxd7kSBASLzz/3YqQknrwexnTu6xHHugFcWsxoL7hw96d4
sRPstt8Af6X2gOv0oDxeGTg59+GhTMUehuMc8I/3gzVWN36FIrQVXTd40NGBWMaL
3IoytY7yowZ7q3k8O2+Er2TxpAixFkD/YKaaMinBad+D/cbilvclnMwMZG8QirEf
rF/IQEWbgtTZdMiNx3VHScPlhbfQ+NCtfQufAvgCi+MJae47CWCUBpxbNpN+mdvH
77OvX+oRwRvOuaBScAyCdW84rrjp+zovbrnWFIKfcH+KQsmwSd6WLbZumwpyQBtA
rz1jBJxnH3+7kFAKzHi4AN6NShIUbBkpwmQdXiKltrh0PjhbJgh4ln2HAWskvoBS
VazMWtOXwtrxdm8PaB40LBOqPtTgLJPZiFVIoEk/K13jfg+2l4wtbtvhqPjnlDuQ
2AL5m/6uDtjxTlRCfhEp7xLpDH0CZMwWLf1EXmzHfNm88r5XJosgMjgiIWjNR0+z
D7jg/QbfiWX25OmsXnU1uzFR0ykM8wyy6d/3Utlpqpflidt1O7B5X59go6BChjGB
YnP5KqSvO3WhRubOhOSvIW3AYmlDu4lyvDGRo6RqQrAnKgAi76Pvs9tAU0g3xPea
aqn0UutSkx28S1rZA1ep3rv3viEKBYVf+ssrlMqg/add6EynmvPwxeYwR7MkcEY6
8JoGpt8A5Zs63QmAWe+PFSAr8OCiFdwjaqNaxCML43NWMyAkiROQpWuxMG9LRSrz
ZOCeDkmriO5N/Vkzu8FkRvyHBORQ9xtS28yr1sKIufodvqVtTp7lhjBRqC5whNYS
v88WjFpQULBTzosPy65Gh4tt8nd5DGu5BBvVLl2N+KlXoDhkLWnKpofQ/DiPBuyQ
fIRIWjuRdraQVOt7xTU+JiDnAEnuuyMcdIYG501YUAci6/fVHVdfkF38yYfm2Nny
oaZST97B7ItOZ4COkf3x0FVKy4wgpQw3YshhhXxjM7DKdL10iiqeLLM53wWtUIY+
UKrVzTM70bOCRnmYxchOgNoQgFXKEx9HsDadPmhkqf9WFOuY75EBYuCvLBy0MsPY
kUe4v7GzC5S/rFNsPYQoEpBVEg8pAIXERLubTK0Aot9ZkWnxnaUJhWXq/mnOzsjp
zrVhJ6wFrYU6+tApBfMbeGjqm42XuP7FGOIp05Ep+wMRVUMBrbd5JZ3rxWHmWe7s
MHXig5o2fMmKcxRYlaAChPgH/i0FckJhtvqz0bsA0wKO2mjv4RylD9Yp1S8qCjiN
lf5SgOCaCu8YVyfOP3k1Q3/bM21GR1n4KrCFfS83RVJZQj1z35Q2/wtCzzI+q5yC
oS7nGwZ1JQrnoFWk6Bht4VHc/z4mB/NhGgjnThyZOCWF/cUzhgwQ7fNIIv8EaRX7
EjyK13XtdCgZ8oVeTlM5kqeOyHO0TXVbZFt1vesqjVP6dUaAMhV+cjleOhhyoHOM
Vz4hRHsVMNMWpxb40bUDohOb925VhwUnkb92736H4s12Qx7FgdJ7RJFSvcXwqStU
XOHENV3LdkZZnhqAYShO7zTK1BzQbBPfKzLcPpj/X7wUOhv/V2orE/aZpF2jkSe1
/gCD43VUvtFdbLD3xTaqugjv4hiOf1brvhtzV8ylxOtBP4GT5/ld3VoDqlMnuirG
1+x9G0+vX1sUDWhaI5FrMYHw3m5H1Aa4ymsieqLLl59ujSugxFW3MeZ5lq48QFdx
7ycv4NuMOL9OeNZEcmEhcKSSQb/bCWMMh5DFDJ/S7s5PpeZLT3z7HDFqs+vnlXkY
XlfM8lWK6vdd4yBPNWYKRZtDnkCUiWbQgqnc1yc1xhYRBHRBED/ntrgDq4hFZIx3
crjIEBnhuE3YMtLN5k/cbsxAx0ha+qDHFZWutcdAjN3l72N/EFJJB7uQmC+duNnJ
gpEV9IJWpqu9trD8++GKpRxW279vraRUUaKOZw9Z4M4qp5V7YImqQNZB2TvSA7RV
uuQXfqYHzEZt+NmytqPV2EOEFZsgje36lOozeUrf4j1v9z3SdZkp93+6rjeCOdWi
knKOyAfhTx9PKWYAin+j4cxmjyQmtB/Q5OlxxasVLLKzeY+hH9VuIEVu/cHlMEHi
DUHcn3JLK03EaD6axub2ALLCoY020zFQ688gsxYjll1cE/IQXizyOzFZ8rD/19kp
Ko5St5WGyH/jLNapokZI/mjFZ89tLkZ70DjC1eunoUMWicZvIz1YgBGnnPrdNHYI
VHWdgul+qPdS2yi6BHDzWl5Oss0nEqESZNUTfZUOR5nFOLWm/FMIp2Y55vSE678s
OcVLf9W5W70NXIJrxOWCcBzkjf2pDboA8QSdL32QwLnRMvykvkZkjoDXcR1d8dna
w3DuwlGPbRUeRjJZlFvNVT9ZvYD7mPnnULR9+5eVFpSMz0c5kPY4m0S9uwNih19I
h2xzmw4legfwfZwxZZUza2fOHwaUix63yCXyRM3QDKUYHjEfdILiAPaS866EadlJ
NlJEelBd9s6IJ8hslp72e9m3eMeflaH+7xWn2PbFHgu7/ZxTuTCRlhTEgzrbOMp9
jrePUZ4j6tDCbz+kc6YU7sCVJ1zBxJyzmcLZyjQ+bw4DyRUcE/mbnv4PQtq/UTNQ
DtNOY4tkyZh3/flMcyIN7rrFXnWMbBiZr2j+BbjOdGM1AD/zaW+EKDDmK0qbq05d
Sp502ct5xhz/avd3JrkRBz0oAF/Mn04ZauhTXEhOOTE3dpnc8cTuz2eoCkl0Qatk
BUiepWfyyUpmJl4AacW6ju7PWocuQt6seAH5f8UoEKrJ53JIiZHFo315oNU4BVgJ
svCX1E4VwogK2IiJ18Wt2g2E8w0UzMAaOeT84eKX/esTCwrFBTnTbawp83QgcWco
UzsQuNfg2i7qfUhNHRkhIVDhlX5JRD2Xf8ydD9m+qx2CkHeDJypa3tPzCGhsK3Ga
ib9qBVOSt1o9lkmyo/v88BfnIwhx6wu53E1K3yoIc2xwLrW5y/pCECRvIMbYTx1p
HPiAqtDIN5mGQrWybH7SiWW4y8YndqDWdnjuDhY21ap4rxjowZPuvdQ3Th7gpbHd
ao2ae4huohvcmL5kwirk89Sl5q3Kz2ziUFftf/Bj287OpSwZl6gUhBOIOIdQZWNu
cgPFxaY1Iausm95zmvwHAUqdRNbD5vXidCg8/+h3wi0L+AQWGwgJ3wjET7Qmanj0
DzjPk1QWuvNifK8+qXl64FAxOigwGRuOuC8DRJWzI8c0Uw1sUXWyuviIaIPPgJ/d
EGDjgFZrsw7eHEZqS0phd8iUC2oY1TH2M2+VUrgIYd/ulDpvY9wSuzeiK8rNiIQ8
WFoo7xgOW72xj3AWDPrWrvL1a3zHk/sPN3RCrDZHQWc7uBueeahcJUfiLxuFKxO+
7WSneOECzzarGA+PCF3Elz4gT4HrLNpnH8U6/A9m1JJ7pm+RMp+C1du8ON3KPpPt
lbyfTVrfYLbfzFUfRoTIvUJFUPLcZfmWQ858zSkPyUUzVydJ3h9Yl6PHjtGcBKK5
Na6KHBq1modl1UuQLSK3JUgI0ImNwehKd0iTAMPxw3tKVuzLwB61sxZG60KnZBnj
K85KYcFIp57HuKQ/3uSVNpopZEK8pOtBuomuMX1L//gqXlIw7SZ/qyO5A+hQO/qI
pDPxz12oICCFOUDnhgL4IjtkvifFDWk2OdqPjQwXRoY+EbOMFG/+f/tq51MgCMde
ozkC0zdl3LhQBZrbwZ7HKznYVp6HzR6bhxfPU1z2u37c96ZF4k/PgVhNc65ooVrn
J1qI6zNgzkD/feTuCDj6/acP4cIeVIY0linATRe2L/JSTx20AuVhJteCyNdi4VT8
xKN0VNXTIFZqMQnRcqP1fp6G7y9/65RqJiRDB5F6TRguPRo7+S2FxA4QArAh4Iib
PDCcxle5qW+/88uE9Ol4u6t4CApC25tkAIo1uAJMZAjN8m7Pk3FBXpIXePdtAEOa
onmKv+v5unGcWdric78ZokggEi2rH9+WDy6n8KA/muhtFc0WqrNyYbo3arBC+ZCp
Hc782ytsi8rWGRnTZIG8URCWXZLroTYyxFx/dhV/qLzBi7MoCfRpIPrMHNgRmxXf
sOK35erBtQQlzoEL9j50AOWTjcA0FqBvU596RwEh84kqKo0QbaiS/nlHtUHUnRME
mJZpEvIRVWv4ypAZhW4vir0DAHblgPsLa9uOQ2qtWHDRPALDznXDHVhvR/TbptsN
AEp9OfbFH3mQkQHhaFK2BaY6pwwyCL8ZaVp9pqfeJWbFUjSWcJAdQLzL9zht2T3T
Focfj+KskttxrBosakTSimzeebmmaMF7Qu84ex0W483WlHajKrjapllkfslIFGMi
qwOBbj+kqVpmdntHYnTjxul4bMzaHfisTqMVCSQg3H2+yVI3m8CbH02VuLVY+gqx
gessJmwSpDrm2gGsjZbMFgSE+3UWeAFLhWA86D/JH6kJYROKZFzh/nBRQO47sWLS
tPwp6ZAuEOFmm7gyu4C+IQzTucZj1Wu1l1yj6X8+8oN7VOWrsLoUgtoVI7tStnHD
Q8KnxouYxp27UBIG4Dkv8kvc+rgb70s7FX3Yzzi4dqVmBeftvnGaFDRL/PgcOnUy
SxpicJu5QaVP0+ZDrM5o/EntDZ2QJc1PxK8Bgr6We3z7fvfSQF3tcU9aVkl6K1Tj
HLv0CK9j4kvsuIvlmx79GSuSp62lq9dBe8RXCHS77yFwJfQwp3SkmeMSYkIXpG3M
/yhGB+yqFo1JK5OCIlVpAY57bjNtzFrlhEmBPyDmYG1v5QcftAmz57PPXlg7MOpE
tCMKwk1lKjjkYzDgqgHJutiSAN1JEzGHUKCeNJBmklprTa7jHDpL4w1zlX80zfSj
EkXdRvp0gcL+IAIp+UerJJt/7WmqtYJg/AS0m0Ii2iTVbHn5n+ShLPlqhULRJZfu
4famV9l36cbfbW1RFJ80gFi+wuIi6ChpmKK0CXZMR/TU4xMUk3+i66FWuZa2FXcM
ku8+jUDqOVghNA4lf97NnOj3MZf15Bwrg4JoCmWuNdr39xS3QG/JKokvjbGChmvP
YrZLVZdXsDROCMakIV/z5W6s3wEYp9K0vkAuCb8JVUIhYsyZGVfAm4s8GLms/EOX
pi2+fWqArKWqSbU15Uul9Es+LDa7M+wAgVqmdhLo1ylI7/odT+yYEZlrVO1QifRS
gFJJyyOjfZugbSe3qSws2ZAdY0AWNB5WDcINofgDsFlkDFQh9Kcn2epmwF5755Ma
l651jwuTy47zbhDL+StR/qDl6jm6l4oejh3w8ozoP9bjOID+Jh0fRlQDT6vgZWaT
3TVtFaCGliCxjyg7Ep7w0zbC8IN+zzcyfhvXb2cW6XZnI349TxC3p+b4Bei83iGd
sYnSXF/ay4gfy7tHkrUzGPykTwgJdtzr4Ar0DxXvCVUzrnFYLgzAqAMCI+XmTdLL
l/jkiYrfFCz4cSpFBuQ4la6U6ufpr+07PiEGGxWqx9VxBNfWpdfBzk07hBVX1f24
0EzST//8lJLnBASinKQdlmrTwAilbz3sQ4ZVmIdvQ82CC1PThVE49/PVi8hTx87J
ezMqCCoQQqEo0uBcYP97IvScg9DDn2DRQcxaankfQ3lo9mNMYvxKfd87cmRCagv8
XjUpNf5g0GPrzdBzeL48m5iVLk14iPOEgFvTBHxHbd5KWyZhbNzC+o0BBhKLpMLL
jqJWqiPijqR//Z7CZBayHtG0KigJPStLz2MCOrFTN2CEiIJlCCc/gc+xTVNltlkJ
6K3JEMH8eoCiKV75OphuCjkBAyU2gfVBoNuMIDUdsbiwqpeMFPSnApmlQNb4jrdg
WTz3WLh2c0aQTBoCmrI1PEbn7Tdz5lof3RnYW8cW+zzOQ3tRZjiVHImRctxOz7wv
soxHxwTSdxWbrrEH41/GGd2dioyn1K4LHYaP/jfXvJkJKgoVp+vlyQ5x/rDkTpL7
bQRnhCgXvsMfdfABU8ZmzD6OvZC1IrOdyhd4IS3MWhZN628Kbtnt+80i8ONITAq7
h6Z3VI/OBAG3cMWzgcD3Z2OuLbrztkl0zOqZaCujzPcnwjagPAerJMzBC0n/XzNA
WNn3W/RBPEOJbvdczt8+AZpFTNz39CoTP16mtnM13M7Wnr6kaDz/1YbEYZSiHaQd
YPZoRzMTy0F8evJD+vZH2x7KWar867t9op/2rdVsQiPKJQcsmOPlrdvIiAS1QYpO
Qgngk4ZsJ6JeZzqG7I4FBM8VVgmSFZNH5SOGiY1NPk/sypRnEikk3oYJa4y9QVqc
S/FWRy1N/nvYtPFGOTzA4LvfUQGvtsucPGaUtxp+8qFdhmOiAxjN20pVQTfWqUh+
SPQKGLfTMEZ7+mbRanGIPNLhqmwceYo2bVAPg0phtz9o5ZS0n5lf7zYZg1wfhDQw
VKfMyvM4sAKOqCwWBTn2Tn4YmB94FH8jAkf3FmhP5kUjZCBM4Wk3ubQSNAjXDB3Y
2QOIGz7RI7HwUSXwIhQNDkBgzbMyjkKvEzn+Ug3vabsj/ArNw43tPaBKIol2IGHn
SxKJGR6dlSheRIu58mOYF7OHyGac9WfqyZ4tKjw82MeH4UhROBTPMaUxBoEEFT49
vHUTQPG8ak//FdmhgSZ99x5kbb6HqlrEdjezt6KMYkw2tTu9PyKPk1gb8ODz6hoc
aNYy2KS4isAc99jlnga+cThnxLGENJzCpN0crZ6WqaO4dlQlaMM9EjuLBBAhClJv
QkH1UisFM9p1j0L/wcBid5SykR7LD41P84nT0JunaZx6YzifJVT2StYIRlkGzvgX
KtaeuM6vwVOSo+ZAXpWgv8T8yDHYaXvFnmSkGL4D1rWyCRg/iOmmGQ6YWcuWxaq9
UBgWejHO5HltxKIoWMUHOeJ0+knrSjjn6HiH+skmBRvq+nCyBgYJvKKAnpOV/wiF
FebtaXTPhlsE/syOycTmYTn1icnFRI/lpg6Dkl/79UMxVgxYboDCrENhAihGO1Ix
uooEZsZPe4DyVo53FPGJC4IS1VsLl3Iu8433dC7ILej+lBxCmQ1RrUif3yZdkcgU
jEEEsAxqRZGMkWEnEMBWgW5gPMoPF5Oaay7MnupkOKKjxZdpCoZMST7Uy/beBmt1
49ppBms3IOmKspyUBIi7ytuyKyWBMvHmSbRr25kw2B/2kTab924e1NWJsjxmjeIH
O5OHAjj4WDp2nmma0PaG77DcR2wJNCx2R9VHJlHMKdnPlK1VAD+LutkV7Umw3dYU
Th6c/XkJsYEgRfQnzDIOLOqkW5AbrUR5xsAr+GaQ2/viffFMIzgl89PyD8WYqBsF
1YaSQi6iK79zetqQZmlffVa2pHuqvhzsxdu7wd9FBShgWaxn8BLiKfvIG9y72mum
9mDyjkJXy6BgGXRmjy8TaULKJc3kJlZncLI40+3yy4PjJKOo4hXuhJeyLmsLdcHw
dhXwrZ012NbpXtokiNd1jzKMYZ00zfIpXtV7RO4RDrvdhQ67kvEEejCKicyfy9SS
eaqCFq0mA36P8CRPV4ruzRLoGwMxDDCVJa9/Wh5R+MTteRuD69w7J6Ed73UKCwZk
MhpcUKpl6TZ1dyMxilXE85QsfT7WdkZYggxKUx9IVYGSsp+LsUk4Zr+tC9MYNgdz
HTvjZM6Y5R1T+CHAHL4oFZFqtVEL/N0KgTu8a30B6+ui/2PXvkOvE3cnkN37J8j7
3+QpWenHSczU85LCgykpO57MTh4H4bSLYtB/zBwO88ACvvl+z799NhIIWIYx09dM
6ME9uCXYyhmnVtW4wzRwajBY0gGJar+m1nxRI+cGYTwIAQ2MGZegWYJG9vJHnq0/
6P1ctbI3jk906ePSXywlDP8td/mblVOJXxoASOUv8A5LDaqs6GiRyrlPRW8+F9sx
QIgODTq75RT0ZTcyHVqfODZAJ7DX9b4ruxLEH1CEdqAZ7o5plxCubm2DSOhU3wzO
arlnhVAkATQ3zVWNdYuUh6zYebvD1zsm8rWDN2PIeqBLTscdIEQ2woSG7CXu5dNG
9tsMei6u/3kQYQwu+T6IqjktvJgVc2VfX2ZS/T04PbvNkFJw8omVDtzjrSC5VjMF
f4mqKSUS34TpB8zjIYavoGijAJBXYpCXZsOghyO2kC12WbZrOrKcBF4oSLgiRFtG
0IQW+byRMVj+6LFTUw+OyLxvCtjerhFoYUNxG0GALjUHWUVTx+TvSJo+8JsrvYZX
9UcH916nA2fo8HKFSHn2DUEvIhCm+3EydypfFlcDWU2Rc2M1RuJwUCI2OoxwNdUc
9LMJZgp3JC5tbeHMchRK8X4Myb0JR/VDgOjWgG6ZcjQgQdpBocaAWUPFia7Lc0P/
v67Dn+xklxE6ZXaE1dUwcdAUzY7RtHKU9GaUJ82wqfvf/Bg7pWq8NR411wV3zwuy
iSM7KwM5TRqW1Au9Nbs5zNwy5ZlnfzwUjoo7Bkm+IWipmpRUPee3BVDok5YSpvS8
qvpbZYT/OsJ7bCeROodCzi7CrGAsYxnZLweyD5H4dO07j2fSEI2p7pFrQorO8iOT
993X+69l9sYd1XFNkLj0Ox/2roadCIAQU5AID5OtH0ogDGC4GuwRslv5CTgL5gx2
tPX8b0INvKY1+D9b4I9aSwhQn8wnFmjaItAhNdFFk2hxeJJBruCX4g3VHcELV/U5
RxSCOc8b3oSg54YB3Th1cZdGwObtwQzS8A5NrVFk7FRK4SHDkkVAyuFSmzfXqXI2
VVTdURMXSW4IEldFCkpdwQSAFzbhtcQ+GG2B3ffNULQnORF0D9ZsWx9/8QM+3ExI
uDi01+K3D7P7sVjE+/aGvz6zB68yCNkR1++9ysCDQuhkxEd54dGPAtzi67A3RSxi
sljq0H4/9o2I0ISIqLXBgGR8iONUg/ueAttZaGnQZcgZWa69f8eGYRKkD/ynkLLl
bsPq2rD4iOlgP21aXbHHklhRS8/OLxeyRjcNvnZn8F9O86+u3yRo9hUS0ooMJZTQ
rK9vbdG8dVU+UJvzjo85RW6EIsXR22CiOpKgf4kCnQFbCmYJaVwfmUHPguo4XmMh
yfaXEpIklyPlWAmV847hrMNTglylfObIczN3cuaLj35FzsDJVczDL8GaLvS4CoSC
griqs+qEJJsTY8kRqzvdoH25grLUm/u4mzozdXNIL66EOtoiWps3GjTQpiekP1eN
3WZohzTNNU0/b771hSmi6MQc9mc0aXTp4x0aP2qnoF6jYUUmzRCP3BfmMFC/MSiR
hxKHyJXTw1kwXaFucDgOMfhXNcH57XjdcLJO3ZELlu5wSVRrN15SnR0fIjJVW0xJ
am+RObFJhyyVHQDbd7HfP37E+tyA2PioUOzu95C7PIKxO95W0VhkP6CuPIbNhGRr
Qr64stnc7FXgMy3nemfZGMD4ZnQV0CscusLtm1hyUefB9XTgfPDW9SwjYMH1cSqE
s/GMXSntkJ9Vax8n4/C/qeROAUOQCgyo4uykYhgTHThqtbTnNCL/brVAo3l/Sn9B
T1YPLepPk4CIAjGjbYe3jk3Q9k5PCudlQ11UHd4ZGQEjt00PhVo7I/sDOYlR/L3+
0Z9HYr5HO+4/m87pAGXUHdTa3JEMKtAFfegGxFQNwkIHi2XLNd8h5nr8z58Uw2K1
+z7vlB2R29J4IrAyfxsKOjifXxIMnJgkWMcmmmxiDXOq4lXC597J4/qxvYHccCZK
k8ul9B6yDoOMh4yZXDzzk8VhN0DfEN01/yHXRxQhlFOfjIYzVQRO2xBXYqahHdBS
hXGuO1MV4zqLqFGgm7uTlLkKY33NcOiiHytkocMZERwO4Ej+Yxh59ZVPm20AB/jU
wQXBtNVYU/N3mIF6fJenQgzbA4W9oFPyg0hCduxMifAwdliX9I3QwBf4YJvWsLqF
ptlK872pGhUqJicIwRDn5kadrmJHYyg0A77O0BwjGWNMd8LnbvYiugnJyiE/YQPu
xTPFN1PF8BZZp/OlT32nOib9FkxyUeywjMCda0m2nGvMHKa4aYrAG0RSqMv+YHFb
iItl/i9IECC4PuCjjgpzzjyjHvmYdV4V+pEpPXgcBzJw2PTCEc6s8FMNJCERaxNN
g+YzFOK4xew5ZYKxD2tATPrQKvWV102BJ5g1sB77lxX9Xq/CGvfVcdCccHLWR+RY
kj0aiwSlFnJ4pUnCBEWk6NdXN2ZSo7DM0VT+IZn7ClhpusfYaE6BKhJhMEfllwJu
hcW+2KG/R16UWCWWjPDkZmQmLJmKxqW+R+qtVt+3riLJni5h591nhlL8+2j6NliT
w9BL8mipk48Af41gDVi15B3a7QKQcYMlr0XR7TRnZ3QVXB+D/ka40zceKAQbcTfG
Xd3OUT7epiasIP4wr+Mngc2aQIjT2919QpUTa/7ASDXuAjF0LlP5cm2S7R++qAXW
nicYJtOC35ZBl43RRWTr1JvbuxZGR0q/fUDOTsqUqfbCgiAOWbhJ+uWy3ZxWLYWT
4kNC3rCkeT6Ft1pPPQFbYTQ5E0qwtq4RBy74tdPMV0gFKx8pFoW3YM0tj8bwvS/b
TsKRQjGWEAshTYgT2zSrfVYLbrtxYFQ7OMGiukhFyQyCj0Ktl4KwiYy4vi8yKOkI
JxLcJcPWWd+BANsVCIFr4kOru7VHpmwNgI3hbKpQyJBlTLbRy4MAcjor9ERHeDBv
B9om+xVIc8+AA4ZqiywBgGElyEpodc30WuHN40cV1eh5YuV5MCIm6xmw9q9kQ05Z
ngEYi6rbUFfwoYHFISFEhG0kix/KyjtUHP8Q8j139Ky/gRALJ8VPFc1AmMyU3ie2
G7pEOGazAtyLFsebzduIIo93Xlsqf+leG9xjHP0AG8B7MYNWrUjnJvR0JlumfR2V
UEmm6prf+/eYyRY293fMRQcwk5LtJ7hC9PRYmFZIX7ecpU0FxAq/N2TdgcJjn/mQ
0dQVENAv+xhB7/G3OoKS/ozfsceu4tdHiljXxkVIo4YmCuLTrcYCIH0JfbBIzmuz
exE6n4Vshw7O4x1lxMT6kaSYejx/Yy905QURyFiPXlBtSlewZm9PJyzBv3rvdU15
aY5/oHQNDgfVTEPlp95jmENo61MNSB0pbzmHuaGn0ETo5Bl3kq+mXpqQRU/40VSK
qGwFtUMuv2r03qN6ZRRl4Xn579ZJshvWtpix/GrdCcWB7YZoOBr8zhNLywEhPKCx
g3LD2W8OwKbvVM6NMlcqs8zetvwMQCRgNgqg/EnsH6SzSMXUXvxN3KcbFsoKSV0Q
SKEMrA0Kbc6NNRh+Bj5voTramVRLwh9iUJXiIlW26EToQZlnVGpt5AcuCwYRgtTs
TbAmk+fvjEJ5ar5YaXOtOI+hdTtOyT86imPGVNi3QSHHCXAG74+q88/0sgwEFnNo
8mDTgIJgCkoNO+0+ap/RnAd1r8VJseQJudRsa1lMeeNbmP301pyBBCdgalQCHy/5
y8v7npnqExEWXWK6lZlmceybYQ85Xl1GpgKFe1KKKbVMh3f5Gl3MAnjGce9oK/Fs
iQaB82dBIIFR++yyvWKSTjpQUjK52Fp5qG7drQNt1OoZq7hW2pmGc4TPEqIxdCZB
eln0Z/M8hblKyYt+W2+S4+pkPZgPtgxD7kdSW0qrlW04kRDe2DgsCUL2Mjf1X8mU
C7jDLtSyVxd3ZlQhi6XpiVgj7x2nEvg4Q/F5hoGADrUObLQaoqq+WJyyT0MNas7k
rIqKLTSeIMSH+mDOJyBFmiaKKIl/RSwo/4WD+bihCE8T/egI30nNrtwnHSQea0AO
0EiT8QTCgaPK1+30x24wUAtODct6cv4UgLtHt9cDIrxfZWoz8wDkndfsPMMTnYk4
J4kDrCvttx83+7uqhEsO630lmBcnNlpctbZcTRG8+vBMAdTtPm6OFyPDf0xMIxJr
BvCXpWmo207rZIHJkb8ALajPP6P5oMtRhzwN+xMo4BdcBbPdCaI7wI6zRi6DFzCc
4fJn2Lr0U2V1/s272CQat+KhMGpbRdp1D4hGnVIES/n7E6Wni12kdYhPAkdp02nw
6i4asB2is6dh94L92Tmf4PfrdTgPiq3m3l5jiJHQiGWvKMHIMI71wUIEme/PB6Zl
cFvE1wpb2QuhIGAjRBDbikOoNc5JCoPgqibcDMk8VQnbivuietidJN335yIiLXTu
wxDWwOzzTdGXQR/Kg99c3iCLPDJO/APkVv3pBvkN0dH2vcuQpYWqxmP47zelX/cE
kXvNHN5lrtvKa1y+kY4UjmlYFzACEm3SdjnmpeC6KsgiB/H2cx0EnPtb6ZBOMqyP
wF6NQ44YrwveIBa1FiFBUXIzJ3S/bXBRgW+Jpjs/TXXKii/+eiiaz4BYPMsR2ePe
q/WDR8P9LcpbNUEBXjlcUTZk+KICBwVfYBYtgty8y1BTKkSmrXtChuOJeORQkG5n
1i3y9AGYfYaCeCaiFdngM9BgoB+Qbh+aRkSeI6HjtmQjLiZDn07p5usFeK0PaWyg
/kRG3uNQED7cR7ashWefZ6c/rHJYoRNLrW3IzSF+wI1tETgyCbKA0aVUEbrjaA3L
0qtG2z/kHZGP3zmEooSUidfu3AmU47NXLbQzIpTZGJahHt/+Uox9w3FCRP5bwrEh
nUOOjS9+nrUXB0DbNdvXGj2tYRGsv+anvpZGQFYG821CchornxLIEhGVsc0SCI11
j+4prQTTk2+1D/9aKLKzEDnGphVlky4RZnq0pSuws7/Nc52vmQFU4y8W/5sfgFYt
+xEqRZYqn7VGRUqy97jNqsLkVdSmzOXZVjjUAhIh1doIfGCgoyr59jiLCj2jgi6z
jspY7kkzUa9X/fEE1m/IYRlWmOyPUIg50XMiC0YD6XjdJaE3XTh0vxofgkhVqVat
2ti9+dApGgQYTanJz59VjpLkHYr5ydsmZqw/tqJdBEdyicdcxctd5eGfQ1xarQNA
D6pmVx/wddmJEuKEmsIHSjWKlnScQlGWjlNoYIKgVJG1g7/ye9ERTaJAmfDU8rd6
fFHDHcQ1D2UuFPT9iLShhFx4VdIo0HyYTXdsOauVL9YKMnNdag6vOlb5YqbLlyCf
XAg6qdEpfgfmN6mylOMn+E11GrwUu5Mg9oVQILPoqkf1FkZ59NDK2UydiAJVixjS
yWgp1h51g4MR4zyvDwqCbIOmwoECaoX4y9zUvRMpZ6JWRkxAEtELTNc0Oox8wbAY
1x7MrKZ80K7OCSSmCDg+Jiv+40GFozPt7+fIBZ14wEY47ZpRtcTiSOBYG4lpfzrI
rs+p/07mfpf+QcJi0xUV2fdZExtFflOYxoLmEMtvQ8yed5MehWYbS95o2EdccKTB
UBIHk1pg1SP1n6tjbIqvU1Orz7XBS0lsF0YwO+0hAVP3FI+RqQCiSwTATKwrQoLq
xqp0OV1FFkHKy6Dvl1KCQga5xCtgjaEE85DvRueCv4ik7QB3AYslgevd2qMP7W+i
cBx9eGsg3XVimk3Xd2LbBwXTNlw/RELbkikLg4ZVMVqycPIrZUt+CpYW+m5vbrop
/1MsU8jOhiKsa7VfqvG6t4rJkrhSB8lq36qO/MUCKkSmBxNeaFWaalTJg7QrRe5V
EiO1m3H1RmwWNJBOsFLwYfnsA3H5i3llHhcjUUwc2p1AB7H8WHdlsqM0H76cp0AH
ADZDBxwaBVN5TalZaaUcxmr4cS8awKVs5ssj7eNwQ2dLLVSmi5ujCZG9+lUkt3V2
c08nWqOKl+IY0ZqN8WabqwRoyTi0Cc0mXM58xBbq98oqicELuUAHQeYYSd6BNl3I
8es4KlyhcJCK2Skr/lvF/kWAVOFNTtudCZs7R7xCP77q6eOyliy53Ado4fihIVzM
yrxgTrv+KfuASlvIL+XbFJV+xC8ElBkD0xJ2qmkqkd9Tz4CGSn7YV3M9eSWO70Kt
4xyhHbonoP61R1Hi6wEXZ3Jm7HuGUZk7Qnr5f0D//7tHFg9ocqMfwXMNsZjK2NB+
1n0Q3UM4NDnPP7Qawc7Tb77BTXj5n4E1LEkTIYp7OyiCAkltvltVOfvTRePok0xQ
nGU4M16BiiHJcIFV1hNZSHjWzojOIFD8C7kbIA8T8DRdPs6Lnu/uGXJbD+DUzvHq
izecc+JYHTDF6p31jgEWqKz/Y1YYVxfjkN5yAfaLJq5hsEIJ7bbYdutCpCcGE2Nn
SPSMyeLSvI4ZiEfg0p2Mnlgq6xDCTP403gOL4paFyPiceHvwjaZ/q8wN4Q8m4pT+
SIX4Lz0lcfEPS7lL6agDXeqoQF7LQg4TheC6ysY+caFA/AZkfSy10sfd9ANCB6TQ
1545Onlb2djLG6do2FsBc2Q/YwbHHWl/qUzcHY7DdawpUyXx3SwNWMQUcD82f8lD
CDzVvpJXGoPTs+RL1Cy4NN6yDuZlOD6s7VGEV8+hVFTqho17NauePrjsGRzjEpga
0hdasoYZ6KQHwU3poy2x6oSgvBVLKmmwr03hWPtOSoa9i8UwsuD2adG0giZFmU/2
gJglboNFBaNWi+0TGf8APa990NwQvynvB6J+NMkgP+5s/TBqik9NLlavDCwiD0pt
1Pg18CFd6xe0LygGa7fg3/CJmYl/rI4TQnMk1BETWIuTtuRYkdmuQ9GTMNEuNEs0
K2VLLaHgN4T1rtiiL7DCcEKwG70f9E9JWd5j505ZCSvOExNwILhpYqmEYOuSxiSO
UHZ6bWrZmuTGwxaXPgd+NAEjg47Iq+ub1hPWkTQ5u+OpURvKfcwEVJqLK5Hs656n
fxEtBnkaqZK7A89A+NBmCZ+Zp9QxFTuutGq1NDXTASeM3F/C7OqS35v/6IuKky3+
CZztffRHK6TQn4WYpq48ZZttaKKrgwYk10Z/QP/Sd+AIExzznnYsByu12o9qDQJU
PgVFztwtK4vnttS8aRcYE2BS7psM0Fnrsg5N6wpvqRQykcn1P4YtiyhUSMr1CVrD
OLiwIo31QptEgAnY4kP4EpM1vQzAOsp8D90kguwL2xrpZjzp4yD+Y9M+K9aXzFx5
+EjykUJY7p6XlahpcZlsDw92FuCg2uxgLzSI4Dt87Dq7PpH+xd/uq2HIk4vlz32y
dnfJskb2934THwQwdqNiSWPBSWop9iBsZwqO/SN3IPfHX98i8V3ni1CBzcCvGupa
CGNmD4l4S3Wi4B25Ee/E2/Iv7uXZQq7+mpzfg26EBd2VHhNqaLvo8SeF94UIBthq
/WzFHW073AplGsD6ROLRyuPEBYh8laHsAg0oDJ4RtDZkY/HpXi/P9eiQ0xIUuD+A
uezWfg+ihVKJLedIbjj1hO8DFmD38/a8ylafdlthLM49YBer7wd3RRkWCACpA9Pi
x4K6KQeUBjpWXcKz6T39xvyJxAbxP4MwhSFyq51K/HgKnl1T481MdmpHV42xjQAo
8dxPSyFnY+yLGXP2+NM0XecGM6R47mbG/WxZgXrFYWl5HCCeP0lJPwj0dZAh5ALr
oR6xTAE+aWGsQmxaTLhCEj1pxkBCU+qONWT3UZJSq90DqT9AGLXO5MODVtmbcE9z
ppERzE4UHyLkbfoH26lZsbTCoNZusC0cgOb8pb5dWQRgRRGeGkf1/VNs8KoAe9m6
cUMNDpG8uTX7WiuYPunQsRPW8m4S79at9XEDm7+KqmXd6LLjhj+hwFdW2/ZUET4/
NSz0rWeCU8tLcRDydlyrPSeRQ6c4NgpRHS+8smogH0zo91F7AoGiycocPdvEjDHc
FqL88K/IBUz/ewODafaBijq8URhb1oaFfsTCvev/FYABsUrltMTKOFjG1tx4gYN3
CiMCiOU5Kjvi0kTRZ1ytlyN5oObWaoS8HWsrwb/raMSg52t6yVfDjQrz0MjCanz6
l9XWmm9joB1DeckmA42p643m6mhSfB4ZkfIF+KXXyzSa6yGpmLfrBU5Yvxe+I9O3
2nFitbYgl8Qyljz0xwo6wC6Rg8cLa4fidoLx+9NVDcy4eF3AUlDhXyLSqMjpFLAY
DDIKLpzYTPrQXjQwHHrEM6ABwopf9lXG740QkD68SqWaFaVVJ45wAfkPPDqkUQ1W
B0vyLgpzeLtaTOi/WdG5+kUQK89u+lUP5YkM3Pfn6iJCYyypEJ3UIA1ie8USoinr
1+ixFDIAM9uwVSGq5RqFK5hc3BBOiANVSkLcPH/gI/liUPFzMdN3JmI6ibf6bTcP
uJ3n7VlPbxduPso6QRQ3jzU8chK+mIAsA7qaUZ1v3L1JCNvx2S6ow4/1lwwJxFky
ARve8KEAwmbG2xnLiqiWGb+sTWLjPxxvim8YOBu+UuVGbPxtgL3Ri8W09kLFLT6l
wPWPL8SMuzV7kmWdG+Z9NONZkbufkfDWlShnkE8jOZyLm3yXILPi865SNgg9f4ao
vWqst0wYDwhMU1p2RcLNq2UsrsYOz0YI/R9cxUnJu/GUluVruOd6HaOi8fEIr4bH
Q7exgs/Nvio/V8CKiFa+Dsh8QqhJaQw6nUqtaSZwbB8x66QnhR/g1dEf09nyYmoc
dp7ZoMVuxKTneWNzpGOrRkKOLgPSHqQ+jNI24aLSLMNJ245gxS6VR20QG+61V0Wq
K4houKRUgseSlx5Y3nd8aruss+M1GGvNIKrcbiYplGWWUA+M7YlpbtU1yh+ibvXk
ROmvA85QiADTLDEj1t7X+DT5kNXlD29k2kmPGI3r0YZt636gIIt4u7yShbYqdYPj
r8hx64kHNibL4FNibKX2GMYEgH2KSrJmL0CAJ0WahENqfIUVSrVRQX+68Qdj4Kw6
gh+SsUKDvAelOdIfceIFmKS7yqyIOOWf1m6LTGEzscQ4mxWP8H94N8jpaCYfKqK6
GJYwAAVm6YyBNONTcoFF8iFk3XeTu9Aa23iDJefHUtJ1+J59dBXtl6Ct4wHz3p2d
NAXzmtAx037w4mTiy4ZfwIMcJ2JKs1LLQuye8ls6OBYHdGyAyI56uX6/w5q8qTuy
7dYVte8EgkRVXrc+dzFk8YJncrJ1NhA7SPczJGqGtOBjKHYZlAvx4dfbqjuMO9dU
VTb7FWXRFTNnO5cQWpUD/96RvqWQnoaJ7kV0QOkemXP3Mfq/DTzf+x9BJjvY6R+Z
M5mBkAIWxz0JTjGv97Re+lFwQPWap6KDHpcY3tfPzB69AlHzGj5iSk6bwQ525ZZZ
tRLWA6M29MRlDJIV05wXqgYjhIxL9DBjz1mNHqmOIRunlCpYMn4KVTK1+l+hX1h7
CMvxA2P1loAbo/YufnJl4TIYLt7RQz62u3ZYpFpE7JgwbZHn+AppvQhq6tMb/mgO
aIEXQGFILNEEDD+l6+myM/fHQdZy6dLS6cDlKcVUTH8QPHH8zYKX6YgaB3NYayW8
KagTdhupOeDeCrTEEv990Hki/875nnWjYTpJ/VdS/folaooHJ+HP7UAVKkBp4kTo
vtaKfwGAtq9LCTpo0ckDNsxJKJsDajHTyNF1VYxy3Ere0mjazWUvl2iR4BhbY5od
ywqMY+fqFHHfMZpHaQVouYLHAeWE36y2W0LLikVfmZflVYC1YP/mevsUwc6w1Xlt
gevhm9F9ZAeQnk8NvMJBb4CzX/nkhQ9JJDUivPM1Xa5BafALmNG5ZpGuwZT5v+fU
7te5VXEiJgcd3dcKXw/inmdexqYbD8Itrfi00MDFzpXajTf9qYVKUv2xBq4mHYGz
4LCzhq55Fg85P6g51zzRssOnCtdC5WbTMOnEHI2ZU8n1cbxyqeTyphYtsUs1a18U
m7NvtbGLPxhV2WH2AiLHOOqOpe7rDJTgoJhDgIEdtptBO78sTLRef2JdOHHHqv4v
TFtA3WTWfVmlfZM1AkvKBAgVmCmvv1YA3U/OnED344jAx53lCkcxgOPgog608Ex1
0Vs5v3pRJNZLGlBJ8obVUeTBuNrdz8bwGs4BF2+PCBr37gQMY2ZoWa6Fy+2uHLU5
oH1gD2mSiUY3QOg9Hkrhvji3zgcuedUF52xkIcS41TUwR24/UgJsFoE+dHb8dw5M
YyW8BjBL5zyr5kPnYIbrxUpxGlKsa/HPuOM6h2OWGM7Wul4WVyxwE8ypbrJnBSDk
X06BaU7kZz1C5W1JzN+PyOASJqaw29bCZ1GZ60RlpA2fIcJ3BAdDlkOSjUnyGnsK
yRwYRzJbLX7lQLmdbRT38STruRZm8ZzYXfL6g/IDz4Zgih+P1j38zBVNo+ZlrhIc
OvBnd96n04Z2Hr+R+P82oz+4+6pKzi3zYweE9R/QCFh9+ImQHrjz1NewAZxCCku1
zJYg8pNL8FtGdp8yQre8rJNl5OePt2srEyK0jzrg2m/Re+XtFdedElbpaqanF556
klqGhAnsSUcImbNlpXpMzQ4XICFLv+HqEzebxz9WCWuoUpeDJeV61RjRlhbKtb0T
HfH3BZ1kY7ih6mFumnDfNMKinR8rISKQkcU0Lx9QTbwAz/Nn/osduUVLrsvrkq6W
WQJm/QnNLrHyq8xabUtDK9tUCxjleqYgrXX3Kp8QS1KSRO91F5V6seA0S+TSScjI
uZ+dfcb1bnYnFm8TxINPsk12wzBGGMSUXY87bJzZguQsaltfh4ywuBkYPBxo8wCM
kh2rf/rS9Fmg56lxM37cXSoR54ZA3ESiXR6cogWHGII5qsL3oW9TJxtOXlJQeFoB
ywG2mni41+sNygKS3x6j00xI3bg8I2l+taWsjEOkP+gc25nR2h3fp3pF8Hg0QLcx
Rvx1dBgIfW+MaJgO6fARwgZxxjdBE/RcXD+ppDMGOpki3ooXKkQHf8pGvnXN3RPP
Rez1/LCN6MW/xKZiT3QqkLDMGj53aONwHz/lKfrrk7k4oj4kua1Mww9LH+h0Hx59
XGG7iRVMIRR365GCQvszfqKYdUK7YJbIbk6muwqxCgt4wX7twIiYO089ZtXj4qmo
VWHjkNpx82ft5esuOH5fLuZwIBaql5IyhlUWYK7/tEhhkEC6gHpJ9N/9HvWhB1jC
feRUsnP+PO2coTsteR3d0j998j/oRihs2+2QUVACzvp1dqw8xsu6XMi+Xb3Gk4wM
khBA21CiuUqYPtt72lOyVivlfzx/PTM7Bbq1qKsz1FPufT/HeMcnt+uC7fPZiZDm
eBgh1tpBAtFc/3oB/ACuT64UtdeHMg9GZWTNO6ISzxdaIQrY5YWuwfaJUCMmIBiC
B/IJHJgat1KZTsfhGmFW+tU6qVGaHVHgg44pkyE8JBhlO8wSL1yc3v65ygX9B7Xs
nW8G+j4JKsnq1WWz5JO57bHIDA+Ynw4msFJVaZ+JTcLkFtgIW2GczKqjTd9nPVwP
6dzKLQE3/n+vSsS+PoPYb3uXmtKeIqXTseJwv4Lo53t7DT4jibMbT/KjYpHYCLU7
6yLHV62WyTuQ4/QtmJ/cvdlIIYgp4hYkDWrcSWMyzagOAtVqBYoNI6b7676B7vK+
AT5xRGPFwLkQtEJp/Onyl2DR+DizgmpMnk73yHw84ZhzUFltscU3TP+7zRsX39Bh
0eZhzeoWqIfdot15xhlpjkdRANKPquvv+XZmLWswoJd4NF/vjbvDkP9TYLMlNxyP
FFQcgpdA/H0cw0Td1MMZsdFpPnCFxPTjY/zY1rrSwQZI9ShoP6YhPvjrkez1ARJY
+0b3gM4We9XGpMYq8sFAZgyUR/Lmg2vZhG4NNYmIHlNtNVk+fSv8jp+Nw5ezJ6fY
YIYlxD2QgMLWjBozJaZahUIoQhwI8awX2ZPM6oVFP+CkqzOcUsBN0++qW09z9DIg
j2jdvXW9+gFU7UlK0vftG+pZ4Ue0U3+gVNX90gQBNBCe47CycnFM21jzGII+6wIy
p1rOS7cqA3DBr4vefSqeHQk19gcbPkd7HMs6L+xYfutUV7FZ0L53TUrJ9g4ygWnH
U/Uf0gkQ9YWVVaO3DXmlfzDXbbM5bx7iZMyNgJk1YBDJ1seu5WyiKAL6ll/6g+32
CfLtSiTEyr7T5yAPb7Re3A2GnBVyiKgqsfAg5Vd12bYpE/XbZd/TQDRwb1/3xxGY
Dcwo/MxC1P/5dyaYJyr1JkDqcBnlDOTpUtxy+fs2mf3nAknMx0hPqEUqW//uj+JV
RarkYARk60BnnKDejhaPzqATwDBtKeQTGiSz/t7/boyr1EJohzN7Pt+NnXK4VOWZ
nQ+4+fXLEhr0b5Sl5FsxHW1Rmb+Pz9ckwbJlTlwx3Aw4hQuuNVWs5uyqj8HDkCxz
fO+tR3xHaLfvb4cJ7o1MMwNunMe+MjMgQYMuPyIz1Wmf7TJardKfsoUPG+JzFeUD
98rquFhFxlnGvP9lgc8HJx3T4FRxQD4I8yAJcxxakVdICNKOEc6kIn8R8uS1l5wB
+fF3L0XiTKDGZuRHNqX6ED8Vqfs2WRn7kUziiJmj4v0x4Vnd27qV8ZWQAPWoq/jb
zrrjflQDzPgFtfnOrPkjLTxM+vQ0F18ZIzxREZVbJb3V5px/08iaX7TQOjp3nU7C
1enRXcXi08EZLro7qPiLRVl6m6C/Tl9xXk59YuELgmUHMlmeM6Hbic4oPOjYK3W1
FVnE6HuYqYWdj57GrfEcqlYKHJstUxhMetdQsrFd+JsONXBP6uoITjOABeXWNFbq
hby5nsY+tIemMFJq2TzNOP7Nf3j/aCjh4QMi8zL5cCDpr61M3fwztnInEMLZNWL8
lhdiWprXM3YTP9fuMakhAWuSSSYxMGEFBDwMkKw3g7C1fjKW2XYHzdKnJmQ3FiEB
3THVqj9D70OqD9Eb5LKzI7eriuhQXpu+LQY/MSLgjEVhSe0Or4/zRHhJykxu7KAI
56hdRJo4E+alNwMTAFhUQLM66jTKjBFJqOTuNz842X/KcR61lOcWJGC8K5LNMNKP
mFfdf/AFJLQJ0TH0H3asatxHcqvnTG+Sp+QeOLANPN1SvUB44fqq2DzfKhPI5/d+
mWryttTPtYYpZXaq8Q3/XcjvTObperOGYoM8Ck4JcH9mVqV2nXvKqE4kIzKaK03U
GircWKZCD4+mtNbTV4vBMmXy8x1Z95g0ptCa/3uNHl+wUuIFR39n6AjKjNbvMnZJ
5JQN8JoPO0lfqw5dCq4DOlRsIWF36GYP9+YO6IlU/+1iHsnpHTxxNrDq9Jgn89rv
V83Ozym8GTF3DV6r21nq3klM1iNtnz4foTlZ3XAWymRBVF99Qsvcn34belVT5BX6
HaryvqKfaMkAk53PfFmgMUAhfeBlcKh7iauctyKF3FRD3LOTVaviwEb+OYDO8tVq
TR7AOrH/rRx40Lq0dOyK+0JxWX7tsRUUkjF5qygBojESzgLIpC0Rv5k+HW6g5eHe
RqZo7OPd5zqg18T/iA1FcHlCpAGgXvxPs2OqI3lprwhdBr35thJk+UN81GEv/rYm
8oCDskZX3c1ZdMBM6e54ueWPh5N6p6LQ6PMI3ZZglyG5HaOjPtb6HhXjfXo4gz0C
gaIuDif+d6Os1WyFKIx2PW4t/7q0A1R2oOZLeVPK5noDfZkvrCKIebfz2CrsSmQX
kSVwyE9XkpRtSkbC81sUPDx2DNKEhtZH5XhW2Lt4/kqU3rzS+IjdxROacHnLC83Q
Tbc14g52zJAEuONJhDRCc/RE8+mKcC1z+B7rO/V3UWhYfDsn9ydi8LVlO6sqeyON
jlFhT9bDeuTuLf6ZFJMBuD+JrdmynuOXuWQSSf8CfwgQpc6IhbonTQrOoqEETTey
oaC9U0zjMu4YIpnRaHjlY7oaWWSHbTzKbkw6U7FkDUNomPpH0GbumwcmY6r08Mob
vjWy3J1GJXMNBsqSht3FP+bxe6fE3ADqP3DbJW6ofHoggPuTSvvUca2vgd3ez3Bp
Sl2kFWaEbORJpySUtMXxnWfTdqrg9BINGfvOSaQB3Q5dIV5Ya6xLHGz8A2OjoaoE
KyCO83MToEwLWe9CNB9IXZsajXYN1+gXBt/wihcMPosIgvJDTg2EABKbp6Xwua5P
BrrLiWbcC8zXsxLjAMeygur/iODmXoTbqRynHuvKuk+N75dsbVkSjaG5Kxsc5m8N
QKJkphNUYiyUlReGUbkO10DboLGmDMqEn5eIN2ciKWeCLc/13bV8n6MJu6jLvM4f
MnjrmS2hvL7FDYKpdRVc7zgl+3kEtgDiuzlMhuAvK72z9d3CwNgwQ/1WIOPFnazF
3YLRxh8oKlaoG76K5/HXDK7NCMICxBZ1BvJ4cF1znvBT2bpwb1Flym5vEz+wtZC0
17hY5ZkEJpgLDr0J0fylLdc56VcsXovE3KP0O23wsBpyhlEmI4q1rQdxg1hTNhSm
/ZoVTy4JUGWSbTd4MT6bSa+VxsIXptKJBzMpeQPkXFmRTEbjrD0RB2Fn5dlxH5Xi
4q53+tu5rNoasN7GamP6paRiGOHbRQYa7EGYR5t7spolR619NouVJAF7hmU71cXr
oztCzAUe3WLwptMYH1BTzBYPdeOj3RNIOoO3Jw5p2DMOzqxHfTM6T73U/4XL5YcV
A82y6/dOIwcxLefmTCZpM85vjEO0k6Pxe+f5Row8DglVcnnF1MlQrfHxoHiWY9KS
n6a8IFT+cJJODjHvYK2/93BJqwfD4TZUe2lT27xpCCJseeKsSSDhTqZ5Wja+xsiq
jksfxV/KPDZr++/suB6gJAVgXWHfobNwOdIm9W3fyGKEUN2kv042IRutUzGG6pLN
pMHCVkuFHTBgDDtKWSxYhRU64SqVA5OUqhbwO5n1/UW+3iHjAOz3iObCrvvN3IOR
V2Q8OA5jsTzHgzxs7mvn2ecnWj+hhuCyZ9ONGyRYvPXOfxccoOrOEdUbARy92PAt
QT7TdxAOUkDSLxmLPs81su2R0z12v8Tq65v6YfnNM+gdi9JGQYz1515wB7G6UF6X
O1JQHSjeav2MvUh7+BA995LNRf0+2rp8mAY4SdEoX6h89dbdYzK4uCCwGldmuRTs
ufFD8yV3Zl48fcyvBz9s8xV4T3gy5kb0vgrFwD1H+K1fcMXMAR3BngVNaygAe5kj
FS+PECxaEHEmRVZyDgJmWodw04ASmLs7Y+sbj/riIlb12eqV6WdsLN5c4fXFunhk
VDXcRRYGRZQbEODD7wyMFm8yMQuLRPj1y9gQeH+T4sjAVSY2TvVBtrmmeHHd5vKY
bFoTNSXndEvZEIPOAp8oXMDcnYF+nnrZOzAHv32YxpcdMVtZzoYBcq+KMHhUZxjv
n+HMtgK1PKxFEtSLjTUQWtOXrsASNabzHvL4fW/1PgXALaYG+CTYX5eVoL4/jH0u
d4eFBKdy1v6Kd4DVOw0u7H62SYTo2kXkXvThRw6uTx3Jw3o7oF1VFNL5KIx5Qlkg
c9DndeaDdl/LVXxNOJhp2mzYHscbHP9fca39WTBPuvtMd74JN6TdrQiNToi+j0pk
uTXTAbNjV5drwB2ntSUAm3ZkoICBiwf9D+2B4AVMWZiTkD8j9Mx/sk7r+f10zcGR
qrXpu5b75FvZ8uvRknJ6irDUT7Qn04xkEC+Ogksbg+zkZVlkD16zam1TuC45e98b
tqFrS6YDQC8HUtvoCpqR2MVA/QLnAXlsX1tNK0nkx7M5UShrJhH3XC8jxsNmgjPU
sqkexynHGgrvX04S9G7XfFiFwY13hS2QSt5YpFdiUwtWFP2gQ4WsyBbV4ZXuFQVK
Ff4reuVP03f2semDAKHPz+i+RpF7Mgd+ixZn7sPMQNb5UQHdDOt+PQsmBVgTixfG
fKPQFgJTjkaibES47fSBVgoRdXaXw/yhGQOI6EzmtLnN0BhJcNRI0MsNvjUEAjaV
HqEpwesLzf0xn4v968QsxHWaPLcWjEiK/pe8nPCq00RPd3MiKXKK9pIXvM08LqHC
cHdLLJuym4hiTpAztGapoeJDkK/MzWhR2J0dUGBviSnSaN932vb09osePyG6fMR0
UMAD7wvXWQ26BXQzE1938Jkf0xkjZ6ObK1t+ycyEQiZKCndK8YikU6gTTeMSd3nZ
f9a2YK9RYlGzTTkVOgV//dVjBftKFkPTA7y51HOqzvK15Z/QKfx93xxa7yBuCZNT
1jD3Jks1tPci4udmBQe0Rx+nNhwCTCoyQ82tCUVxAC8thR9PiAZHk25PQiB5LmCb
WT2UZJ9IgvsyYoE4YQskzLZPUIoZayqVo5PacLB2/6bGMV6NAEBWLViSQgtW9bep
PkaxzM4FUEx3/D2Lk4CG3vtNljiLe0+izE7kLgTsQWcVvB/3Tv98Ruz7qUB03TCp
rexuM5ipS+4XGzpDTPlBZJpBPoBxhqykGwt2K0lB/d5tO0etrBNSKIpFQ4wqelhZ
i3jqr/cytJ0mTGT5Ms86tlRotJrKG/QgFVUlWSnOvDHVzRENo9rHVBGo/BaqRt/h
PJZyeN4r6whKyT4Qg3DVxoRN89bzZwPfj1F80c0iU9IrRSRHf+KrC6JOtBQBiKHA
fSNlRLVMjLqMABZ9R/MMqsKpSEgWOYkh6dtTKXq07N/ybEb02l6/bekBUIYu37hA
iltAPp61HHxP4apwDyuVhwDW9taWyJA2peHrLfDknrblmCuj3wH0BYkp/z+yYNoh
Xukd+cpWfR40VrUaJ/mBbMgcxEVvV8lNdUszOpscGqUex5KT1RAxH0D1/3zfbYKA
NcwoJm5IZ9SEnF/g8A1s5sVmx2jhPSDELpnEv9H6l5ChvGsI87t24ICSoyZlSV8e
0pkdnmQJS5fm7KvBoif9h/1ygUYWJoA1c/bVvzAZ/C7Re8rvVSaOR2Q4TmFK7UI0
ZAzOCeExzlBtCjtbuiU3s757GZSZDC3LVn+5PofFB4J4MbgKTj2u2x/PyaeRZGlD
vlPDKl/boiDQFK1AJqha97qotegkFUJ1ZIKpW1XqE2qzs2jjvYcxfr4Ex+rVUl5M
rLaMabQN3nfe55B/94SqcQSkHTt9mCXhI4B6msOSgf9KO0LqRfZEAXskfNhWPrEr
dbrnnGVb2GQvZjJTQmuHPaaYWMSJUlOIRd7rso60kMOo+k9TWABLvJ9p9y2y3MIR
IiqDo4EujYZT8CCIXmNukBM8SDbJKQat4ust7LVuIhUNsOqnqAiJyVPYQZh85N1G
Ol2TzYb9hyNrL3NXBRvjSgiCfZLSG6BUNrlSNh0XCPIduMkrwLzIkrrn8/u6Cy/7
0u2ypNCqcS/B2AA6HqgBu/kFL8pqmm/kOkKFfD/BgeJ31RA7oOwOLKIDszNijK1p
XxgW0q68GeNy1K4yVP1f9d6sRtBuFqRnwZXBNyrLGWq812BYgj/bsa61WTCNSX/Z
3BPpYW4V8RmhhWB7ke+npPl/Woxc3Um1EfiFlVU8F8hOMduqGwJG7GhSXKde1Wgd
aI3Fn6HZkXctjgTaRnOcvbgFb3VF5PHjTw4rSFG2G7Zh+QcsGUw1eJalmjtTYYcY
lMO/kWB7OB3lhsY85YWx0POjb/+Dv2Pf06ihwFXLJp+4m+yYEMUTfP9cgydzDDN4
brkg7H6+qTsGVQyJE89LCRMT1C95BfCHp9F85nu/OBbG5oZKkv5eWkFeUH3NHQlt
qu9EMKtaOTm+myaR2irpx6bykchDXONS4SXIjdCYK4LjTd18ix7BoocJc7A6zq3a
xHBpdqRDZHY2PoisYCQzI1vK7Ky7BS8k1kkld8ry2is8q0jHPuzMwexjnpQ40ymx
A9WysZ4m1/z4SyLzystGdlZKyLISiHPQGqi0tBT+0QLrjEec3fWZ89BgiE7bnV6f
QSyPRpVvIWm2Z27ZUf85KHHZrCXdwbD2uEgOU2PJVN0QGyfrifNyg6M4dGBjDoLC
3d0KiiWB69kXuclNnzkgOeltNUGKRyv8DHj+fcA59oIkluIZow3FZX7eVnHPZYqF
bkuKnVHB9M4n6wSw9qW62kkTb+xzZKv/SpICLUJ6t6qiCn4JPN9WK39OiaXI26xg
led5aix3ZAVaxxqQhM0/sYuzFnVLMu6fnWJOb2IVxgU7YTpe+CBv8Obeyy4aOf0g
Qnt29mRrJ/7n2omRMpgXpcLz4/kbrjdCoU/c+REwBzWSB+LN6qI054pi2TW6Hh7j
J/yCeVnqi7pBMD482fnpmIhHVNNjTf6SoH4P0RgAv9IiApmMC+gp3zCtY/xbdUu5
up7J5bLhn8qYBrTLKbBqZjZJzMh/oTshYT/wfCDYLLLQVzC2E1lCYNLaSOA5KB6o
uBigtY6UGyg6xPMugjrA4dUN3JTbA9J/Eeifa7BF1oRqKMRB0TYNYfaMJeqqB38P
PjRkOqVWtuvhYcPfCXlUzfNpc+gDbtmF2oOJcFIgj1KIn83DN/F3gBqAIrrQG3E6
QFkbG/dJh88cys8QojOtb8ojFMx0arPHKgB4WGjq8pcTIw5fpM8AnhoK6WCjUXdw
iRnWz0wDSbxDGaQ/RxkBtGf7ZGzMa4X08Q+C6VtX7brbE3F7VizozRCcg+IGHK7R
k7D7sOOVhOQKc2vdGmjfMQ4qhi99TkXtSboLOOSOwlr/mQqQejfuiwUBipe/7fEr
6N3A8uU2el7EgoFcG3vnDHnUuN4hIuc+awy5zdbxq8z9d7tD8C5Ltd9WT7AsN3SS
WxaTDn+p+rID4zGw+HNRrbh9IB469IgWhUkmsXH+fKChpWsh8Ahn0TCNJT+JdSbS
JwB2oCw8DVwDZ1KDovCYKHaghN5F9VW7x5iYokyuNdqvZVGAwUpsgFMWO7YJf5G2
UKd0PdoZMB8SNL0caa/4UvoH9Po2t8Bg8yBiSCtYGtnNKbvA99+dMEUmLbTY4jLs
RS3p4+xyJeCKc5M7Q9SWmRJwmA/JAfDdN8TXpzpsOLiUMNJzRudjr6RADhFuTr1a
z+1kPMuUfv5mTWdXNAnzXQEruIU1IimFtYGLlMJ4cj1J2hG2c2N//Vk9L3JnL0rl
tehpSEXDxSNYuZboUelzlQQCBMJHDXaZAHkMOPoMQUFSr0U4NxOgxUZUPiHgaM8l
KJ/No/zIZRWmshIT5qq/gVo8aX/yalwqOUhWrS5ipG8IUwA5+Z7BIWw0o8TKqUDM
y6ks7ESyBVU1kVt1mza4gmt5iieUoaxfi82cTWUhwzRgxxvFaypFZGsFgpdzVVrZ
K5IO/EsSeUFJohGTl1HR76uinDTgZluktINg4/Y21XveQQmzjhpL/U/AY0mPbM89
dsn39seaA1sc+ID+H2MV6AYRadVdiQixE2ZaqW/L5FS0WI8TupSFvumu82qhi/b6
OJ3aB1bje9SIXF1U7uWZWGhyI03VNV04gyUfmyTKHozKCTfNkV8J55nlVbZrRqYs
ygH6BLVUcoAyXfaBVyX8pozrrs54QBSvjRKm8lrAXoxG4mR3fEYmjL74ReM3/Iyo
fO4lPhSBl7VpT17bSif4/Y0gNEOukAbaprzjfAnFlCImkgej84Rc2WB8z8DU/ouQ
oNWA+9FWHLuiLKCcMzE6T5uhhTo2If9pJADTkGWNs9DZJfH1VzZaHR/wABovFnkC
luohbW1fmKb8sftrESzSVxU/dhBRCuYhtiY4bcZzWeoC91EIE3YaKWZKB24eSB9I
267kUsGzkf9rm78vbpVW5X/Os0W2box0jN1Eb1UM2XC3H8tBpBRDOHxlQNmvnjiQ
bhdThSMP66LY5jQaI7dCGgH2NyOMMWlG5pKmuw6I5B+cRQmRJcor7vhVnOeyxp+1
EetzzGuEMsZwQ/4+SbwuXB1rBqOFTwpTdkduOy1S0arHFH44TOjGhqbhyWH4OU+L
V+/PxBoYCoBm+1RSvgwszY6w+0IvcXhL4xznkydtrkYR7sW/QulHt8/ywS+ZnOJS
aSfWHxMXIAnLApLlN0l8aHObTreBbKb4PDLN/B/hB8ZJt3pSDol83WDvvy0UlptJ
RTspDr/IpD5MScEv9skpebSN5aem1PSNtBwYcVS5g2jEjVR8oOEldehmOhTSdl3L
4z778k14qoSDGh3ORF82K9QDu6h2c7HBHnw/+EOWa4HNw5fg+INsmDRwSYCKws8j
X7qZ1NcLzV0xk5UzAuvfFMxEzrZUpbaTwTGA31KCKMnQEMnbuds8Ee5Qu1jk6W9c
fuoO1WKz2Q2CNAtg0iywX03/8S5IN6s+lc+pJUKJ/SG81mY/9H+wR37rnf9oiO0c
jCnVBe6grwKkI4yInKBFQveo/SLhpoKTBlsPNddf/1QEjVRJhw8jWBoB9th9C7p8
D39WzbiwG4hcmR4B60TBK+9NbcDLz5ffIokjEnGFkaJO8XOvVeJZnWk2joHL1pea
UQSm4EIowJznxla8wRFx45eq+ioZK6GDpyoUSjF9jNGDw7u43zNiPc5QhPd/2OPV
zqODsNeF85whb82thHZEHcyCn1+1O+5ZkN3QyGYQ0UJfG1DSNtjgB3b4kmHJQMQ/
Ff90hcI4jqtNzq6mM+ihVsuLBy9i93R2D5xq46QYo+1Bp63zC7n+fhkvibA9d0R7
gb50J0OByqbzX34MwvnQ9F3neLcJYFaP7zNWAzWrDqFa/lmOmWIa/BrGt5YkglxI
CYwfmaY6D4DvNXdgujcBq2+oZ6z0ByzXn9ll+9cnHDEMWVeq0tgZMewjIAixX58D
NU4W30wtAZzqDbS/9fkpEN+XVbPhizjrAssFkOIdyOJnMBdeppEGJTh9cN/qYk7x
6WjaRjudFvmF3NFfSbCiCrB+Lat+x0+GPCXOKjq0x/rJAG4k/jZLnOfR3Bo1xxwB
UTUdzRxyvftDw7tgNsxZ4LOzs4RPesA7yJIf2c+Q4RWAwfoYwWQxqdqdE/zx0X/2
D0KVkGY7Qi9CG1ooyycwIAQTkNjDrCLjr9BNs9Cqat2o+uU9RdzYIHc7ARf38L0Z
dnoG/L8HDIIGnVLIdHAYZR2F6F5NmAhgNx2oAIDm+aJk093mImMgclMv763k9PP0
7tzYK/w9rbL3nt3wcwkSKogCDn9r5Z2dAnZYNhHOXnAxCYpgLnhe5lf8LaHSdxuu
WXeYET/bCs+0Gw4hjSqHjftBhby+1eOs1CurHE85FXWatkA5J5f0OCSVYOEYmjyI
1lWBgx13Wcomb4qNnuIq+EMgC+1Eo1a7vONiOke4N7IbdvIeMfyku3gjkWQZYhEu
iG1VDg8ateTWHKvTIaI+jZ9HVjyM2JRpYvqoANycBJyPxh+MkJsQGlIfiI7+75DR
BJnXfU2NW4DzAX/QA0OoSJNMeooLbIkRumd66etu/9yP4MMnpjiNWd2Rn5WVksDr
+hHLDiPg7fKahtAaudzvOZkN1sDCCXKjylCl/aOGx7tLNe1Ji/ZYfQQmKBFEL48M
enWp2m3U/UOP0ys96YJEJoZAcfot+U4YpFN+MEr7eorEvTW+HHMZTKtKYTiRyJJU
1cq5jqw2afHk1ZMQMoW2zGX3JcicLRlqadxBQaSTsRdeBXZxw214Su3SjaLfjUGP
o47p5RP6EwgDwxsHtY0v2vr0F6keXOgyvEH7z5TeAsYs7wWS9ZK/42BNhDfC1A+6
+NX7IRezJmT/FkavI/S8hf0PJPH2hJ2vVHkcFuODpiw5yLRuFPzuSKXjQlK6JYqS
akCYgaGF7YIyAWMfJvxMq6gRrIigH46c8sMRQ6sKLXE1ITI9qJkR/vG9lZANWpr4
GYyHCZF/KGZ74a+C0+8WSjqHqcbKQe5FO5ogUH3irhu8236JKTf8aaa68rRtBKkC
nzQ4fVgmvP0bgpI1XXYYO+LUygKgpdAjLeAxPTis4+9X/KFJ5ygCDH2xCFc1mN9o
MHbWcmPWNFPPgy94JTlLPm02asBkV1SZxmmeOKwiKgLiOX5ESz/RM9a6F+Lx3XP/
D5uGSptWeUizZprqFdGWcGaRH1+p0Xn1qDmPq8VTWVdS5zFcMknsqCvSLeC+HCXX
g0UpOiPiJvDP1gbDBImvBX+N6kfa4t/HjJByZWu/1jVsPJ0D1U2G7O2y+rjo8Fp/
09BdnYLS8IrekPWuRAtzOuNx8zK0FSsZ0h/qw77ZVT9peNaWjGNMpiRVgTfYzcXU
TUFX+3qJE+zMxnUkoaPgzHKvu5zDAd4zNfpjOM9rEOfIS7TvbWsJTPPHW5mR94a8
RBwQlHmz6Fwqv7u/jiysvl9KvPovyI1boGgyzdApMGv+UB3MxbSC2BOQ7DACuI8W
3ng4EbEdPXvkIzh2x86UqY1SRfK3sAlayhmDEXw9ofQaC+gbtd9lhccRvNK7mEoU
AHa0EFxWkRUJznSoBJIQZpXg0NrrPiAvVvcsicB8Vvf6dBlrkNaFGDvBuMRyfRuG
zJvaN568kzwC+ShRIB9KI5dfacmiwjUeRt1o26MvIGxN5gEHNOc+BFXNdyU/nPh0
Ane+Yr6Wr0txDBuPUX2ggjMTc49ln9TXjnW/K13g7qLfmx8IRi64cB+KB7uWmpvf
Hm7vzB2FXktI2oHfWU2Dpm6uiniopi0YBdz4lF0OcRMZQCAjBrQ2VYG6iohiL2no
uoI4WIpJmvE4fWmYv7MlWsy4/bqr26zrIkKhy3MG4YyX+cBxDXGLdZOTtvCr9rlM
dPGnL4j0fpgNiWHk8UbJrY9NPKHxelTx35EUGqaAIFHdyMSdLxQKnZOwfRLclehC
hiPJ5+d4DxoGx/j7wiOeh2yVm4nC6GAZ4sBE/X9UqilgvmgrBe9Pz6GoLNoUN2s9
HQsRVXaakbY/w5fGOzbVbSyJcRq/pG3sy14lWnbeH5L+VHPOAguMr42eCD8/GWZz
UFJcZGgyfFmiC2BXcZ+w8xHHUTByXY2QXQ0EJHBVCb8elPMTbb0nr1F3wts5aQ9F
WOjV416jS1DGk55bkdMIT7fmh2iwof1pu52I12JV4AEqGS7rVhdPzv3v9n3sqoxR
D4HnukedQiyCDz/PTyJBIHIIRKbwUtyM8+wzrn0mtz5tjjVOn4kbNbIiAixWUFsU
/v+xWoasyIDAeHci5mu1OkrWr/ZcdK6GYvJfskWOJvg9lzFd+Dx4D6ZQ77EP2ze+
FK1z1LyqP2c/yqPsr7zp55BCD0EJMuZSFqtlHVKyzRJMg6Yev6Hjylj/Y+NXTTSE
WtzQ5wEXTrBfw6YJsiiV+uiaubKglWrwQVlqDAPF0Ss9ScYGc0oNgnNzPwI5X3Zs
1yAl4zhmhGWtMEMHhYLMGIqyXBbBf909NQTXfoF+RL4ORBNdm6nsYoUI3l01536U
6BMXRK72rNR4+5sD/iPBtgKW5AD4TpcVlG8xTOE/7RtCqEuFdZ6REGSJ0QF0hMmX
hJBqLxHxV3RqF2yrQLce7Mw4nuuUxls90HQd/pFFD53xMXsLSilm+1VIYj9C1pMf
3lytTwLxA2jkLFWm1lRpMowgvRJMTcy70jCv+ahynfyjBa/s5BOQeq3rUOgog6Ee
E1yI5I1F3+om47YzsZYU9NM0EDxRSc+V/8yJRhffNhxYIW5ocGfS01Ps/rfmEpxJ
JENq0nkdMKh43OXYV0nwwMUq0jl/Gu01Gqbxbi/unwFa3wyJnMafXGVMU9hs1/V4
xukuqduptLr8NoDbHCA+vVE9kzTW4HMrRw6Q8En3JJQDJWkm2pfeOR0/TV68I4UZ
yghfPD5y4zOK/N8JqJW8U/JiDZppbqPa4asmhFQ78AYv0hlmNclXuzAUnpwuLVE/
384EGk2hObfovg5Qjm9rvfiznwgxfNa/p1EBxajqwJdG9XjUp8XacGSlwr5GflbK
thKpP/YGwv1XicxmvEJF0IC5QHsENpv7vZ5LCvJ+F+hsqHDIcfeWgL9gi88f3hXR
Un9ErqugrG/hVsBP63nFtRZwJcwI7lPZA2QLeveuZ7LkpvPjpdbrHwRSlfmmj3y1
wbqLX3QeTJxjlatEbnFK5bR0ETUlgba0cOZfxN0AbvAhXmmBvn03WFInTJiCB8lL
B3bsv02a836VE2GwCfSQWMTH+R4rBlrTWW6CH/FnfUh6sRqU8G+4D7c3U5I0ZVC2
MKWCk6qsorMae5Rn29LEoJP3hJqCEHcXYHF4dUSyhXG2CWLr1h6mvBlIgZ4yRmLj
EKXcQNiQx0Pb3IDhyvhHA9rKfMPTuhCaxMKtwYddZMnKsnIZ8oNj5TltX+endklo
Cu207XT7hSISjgDTRySvyjJd3i+ALXFnGRHpH/YGL7LL/W2UPlWIzCg2WHMKqCXP
idgUF0i0E3XIL9xWHtgo+Pma1N3JM0vCnHRjC+ayPQBVIex63EEkG+dHwqi+WVIf
KP1PeudG41W6LKsUN0pMzGXQ/RZYv67vNKSh31FAOoBjlgPoACsv/UWG1vPT5S1m
QtzE4fYXbWH2S2poLEaKpTFE+6YDxxt2HwW+dhQcm/O0cItUHDygIds6gmmK/Dfc
DJJcwgz0eJKVT8w9HNZngFG0j51fpnn11iubXMRDxWKa9tre0FRF6PRRYzeBTXiK
N2MdL/5hq8i5W1m5NCwOuOZlAUK0BH5lLwiyBoKm2HRtklHhZZjw6swBwZosLJNz
JBpR3RH9dIoadauZKCQn6kS3L9cjq5k77lS7z87UHLu9QFxBbiH0Vbns5ftN3p1c
M/34OanWY67csPUykjhRuRAEQs+MggM5zdDtg2H87N21aHayAT+4/lSCeiBIgjXt
OPqkpg/sQijNnWciGEeKJBynZ6e5Z8pe77LoWynp/6NMGy0VwixWkAzkMeHIgBNu
yIVrWIO2MOnmpc5dgLA8DDN1Kbas0zWzYf7ss9Vl0+2YOgLhpF82LDTC3Mi/i5bq
5Bq5IfExHOEr3QL9WJhHgUOmBbaI65r2xqplCt92YIDczAz8h0xHYHrxVGK2EA5t
OG+N200wXLdrQ9JC6LenruBPCGav0NOXrk6ITYHJv8QWwPkROfrGMczRdMG2ZQCD
B3ekPz8Ci7xOTTiS0u7fMgR7yARVWwNprpEvc+6CXDVLu7xHLpSVvF+0SqMovbN1
iJ0WCSrUF512CYy27w2C228BUNDFr9tgEbExb+nA4ckMVwabDk8agpXQS9tRQW1D
klr03ZdFRUsXhP/CKQ3oTpik6PdVNJbK/1S++V6xfUkzRwoSWwOHARBVfLkDGQ3p
NQRLs0QgX2DhO2FsGs/UZchpPbjU87O3EK4PJMrTBbNrWF/+RVTH3RX94qfW7DwF
c4zhYlwjt8sfvU+AgWAGRlPv24fkykLjtu/K2gVt0A8Rr0Qgkpyw9K7l1SCISK1c
MbuHaBrFuFFbKNXSMCgnUZZOHvvYwGRj5tuHRlD3gCHrlHm4ItdVj/vBkU+FCHIC
H1N9A8eB6odYYI83n8ozfp0ru/CfjAa+tm+n8kxwXHRuMhccCxgYSgRb/EiCcHt5
2CAl6rh7h+iVXYIUL6HmKcF47PMGHMOLHLfcbr0LpSMGkBS4ZxZbZK9JEcfSsSWh
Dt36dyjmAPDvYvhEbHy6dK7kll8QsMlEp6LX1OJYYYYDsbQCS6mnwENlcYmKEbY5
LhE8S862iSIqcxf8DE+9ZgEDVNw3iDByRlkypMphPHFY40aH2NOXap0B5uN8U1W3
+0EDrr++6r1KqZEKo+txCQ==
`pragma protect end_protected
