// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jgQpLyyz5kJ/y59We6xRjw8tSktPg1iZH6J65bVzkl9EIu93qzlseZcbdwfoJsaV
pusUe0hZZ4gC5cLjye1SBg5aqcwLoJB2U9JZu5qSmORjZN0Z7TLFfbt1ClY3Mnkn
C5M/0WEhdI4L/elOgzIxxD89AYUCCNIFo20kXbO7Puk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7360)
edget2eq8ZS7L/5ESmXaO6to9ANAAPqX2Odkv6Rvlc7Sbi8BBnNfGtWcDeYZOsjL
5Bp0BMtOKcGtwT/bhTwmm0RrNFPGMkO1IOWuownR0bYQ/kDXKJpzpD3RMg/x8U8F
CQ4ys42/d6v40beQnj3uAXn9eY0j0rZUnnW8e6XGAg0Z58THWwFH0NUDSAKftUfj
e0VpcUlYQ4uNaH+wxMuTQAtOEwa1Wlay/cN2pFXZNsW2i8d9eGh3sGqI82ltBndk
L0BeQsP/s15HC0943kej+kLtllMILgYUDXsppFHbZAh3R4uv4qDyd4jL0BTOe8+N
sd3dsUjh3Pg0LAPuLPcrNS/dxjLpub55njOok5PYExPSjS3zT7Jt6RJIxB1f6aDy
MxKw88xuDwjynwdUwUzVeYSm1j3o1VDRmkzhLJ66PasB11aF4GtovJNC0rt4o6wl
oNwJpRE3ssh+Eet9ztcpJRndFjthO3uhRPUw3DvY2/vf9LVeAofbHoc8Y6Cepepb
P9aR4YQ+vsGvm+qYXvLodhelfcczqxL0JffYtErsBCDlvf77FZfmfZAUMO5f5Bbe
pkWffDZMEkSDGIavuUcTndxyvBlcIxY0nBa2HzyQSTUMK/i5bmivzvhb80wROLLe
M6JAsqE2TVJi+GUGWznCBTACPJsewh3LnKBif/pUVJL11iwcA7eC9EW+CMijATD8
D2xgAc7qn1mrQ66rHHyY8wXzFeogwIMFN4EHjlXSMdEyVeAHRSKNKoYy39GKm9ws
JV7+yJE+D5P39qIfOP13YzLtmDGMO+LPpnV9yuMdc+SdT7bwKidwIU2SI0WUKWvt
RBPDyZz2uv79v+mpmD4umAsBqu19xsXmk6+LjVmyNEBra+ebVJoy6S0/Fz4P5DqS
ZFJmemxrIRg4lCTg1p0k8ttQ76jkBiFzokTXkmxf/Jqu7173aiytwmedDPVXLDly
22QPlcNwQ2KjoCJWV1FXgfgiZR0cnFNy7KokdT7/oq8pQPnaN4H8ifw/wkvwGnnz
WQCUMIi9rovbIBJ0Dsh07T6/Dr1fD1q8/TdY2RGwnREIjoT/fv0khM+L9hlb96fH
XVZ1tV+mzCN7gUdjdM7fq6jhztVmmZn8WmyjBZOHxrqAHjtwwmDtBFxcPjd/CQWk
JMuUhaZrSLOuTAMnhi1kKvv1Ak1gdwbxOrAUY8dnRwBB0qCOA17OKoTOLo9WTcBr
s9w7WB6F8XEbKuuvymaB5DF68lOkZDDyT9l9fj76RWWSWWIQsCn+3FOrYJC1uWS5
/RIYFaZN919VBjAj44E14GycZLsEVwDCy4k+mzewnQDCUZsfx01TJML6VFtbvTf9
JADMkl85ukoW/SwYX2R1/nI7BNZPME+rJIhZqiCwC82DqUNB+DSe6sNzO4uy98nx
TE2xcs2zpaWHOLGd7KseeFwA3I7pQuCoPabQyWiiH9Hv2eSClP4LPfyQVq6YRAqO
ttAXEIA5nxtQDDxD//ViRxqK2cVFYaQWmag1EbJVGByv4xAAvHOoe3ySwqO+a54t
5iYHy00SfPc/fhe9AKfFT0MoLQqq5SmDZQnZkuQXyinYPwi3a6KHplP/VTGaBPA6
Sgddu27am80VQ6BIO4+GrzH1DIVi3SqvH4JP1tjXCiqPEAPnv11E3fXMF7E6O8bx
Hanuba7yVIKWc1+d+qKh+L8ci+dGnRflHUqscyrqq6IekSpVP1ufRf52vO969KBw
NyhrtHecV4hmodjWBtpKwhw3zgpqvTZpf/ndPn0daraTEoUnVtmYgcFJuGAhCYvz
fGwMLX2N0uViHt3Xa/WjqdzGxIJpIcvbdblFVm4d3d3E9+R3+TujUsqssMXFlg8o
NfcyOzjmlfRCnWLAtC9ktkv52R9RW+10xAbMpcsrUMHIPZ04tA5alcAPv0Rl4Diw
n8vNCYiwZYOCTGqiFsfOxxlj1MOCUb1Xd1ymiD6zetKB7GSe1Sxdb9nUA1bmjKfY
qVYTESpbpafYqjc+FxYduQs99b20Rut7Z+CPn7f0XqavQ9YJTsAgPClc8F46wRwV
Wi+w1dLw5zKQjhyVDo+W+TJBTFusOxwBB0+m00ZRphGvdLPca/TIDaHSpnZ1Qqtc
vH3V50MuDb2G5KPJ/bvyd+hwU7hEJDJyBR9ElKW+dViDlk+3G05SnZQwviN5or6n
402jqcKK7ZYGkLr/b/28mdxf5gLIVr5h2M1iy17C38/zrAbyToq0pOSRBhQCXORo
dT5Q8UsuHwEFVDZr164RIhm1Ag+rBcN6LQD7ysQWBoJnok+k12BfX9nrP6bX9liu
pH5P3mh3/Q4A49G/DOonLSoBWHv8hGLruTXzszFlwnnk7Wc+4IegNFgv6g7g520h
a/0YGdj50OfgzALdn7epiLwnJcIcPc13rwjKuw5u4yh9rDAqHQEihWC89fAEZEwk
hbJjUijM26yxdWiAO849cvFxcKIT/7QPJ9sWPXkUBj7KGEvrUm50SrvWizyNK85W
IEgdqjn4HzxHzibj8Kb0NXRUGC0MTsaLTgq8z7J2/GY7GHs6uEJjdWPwPIszLglK
c6do7D4qiBYaEadh1Ri2XthCiwFdac7ucKddXS5pCFsUv/qN8VRxJlHZlwirL9xn
94fgb5HrS2dCKuhJ3Yk2XmC+ZoCNTJMIwM2P48h2dtu9l8bP2Eu2ALoS6jgKf13+
IyXCHRmOxVDG39zNZThlcy3iOeqU3MXPIzb+ywWjVSefmvM+ia6D5+5ZDKWMuNLb
T2z5dQy+nbEAHzyP3DhJ/0LT1egSYW9WHqrmmzAH4No6K3LYeC2LVRJDUL87srmw
UEnz+zky+Pde0W0sjPzm3qgXg7MrPP3u5jPjZ7oIe3G2ocKjqYJnHq6vPWh71Ys3
uGK5esQ/B4Ig3c/deLvTf/3qT22wsGHCDoDN8xf694B0A0oB0FXbjt6dVExmm1DI
ypIj2bN+4cqqRA6QQgDe/7rEPdCo4Wxr/X+LBG2B2AOr4KSalpo3XRhznAI+5Awn
/g5gjsGiKBGtQ9om3SoRAtMiPIpuSxcBDYn0A2SYNhbQ/iK7sFhDjg6I34BcjUJQ
K9oLIj1Uk8UWxSS3ctTOaR76jjIsny29EYWh68BXyms80WV9p1F6GBn2Gdnxxd9r
XnC9HQ82MB1ossI5pY9EMEeZpJxRtAZ6zCVGVkl+np08WbWOM4wOBovOuV2DNDV6
ncRCZyxmeKJ9UGzm86FUboJni3Dyl6AlUW4Hb2YtNZAmp5cft30qnLEUZegYBeKA
2Q4xxNPO3I5jxg3nqp9LEMONOjUv+783bE270GUT2v4MYIO97QTe/J7TFXeXtja8
bB0rUTd+S270edFF96kJKJYEXmsM62Xa1Rh3V2a57tQchFV4TjPJE+ulkv427at2
4X5/Lme4Kw4XAqKzv8Wgo1yBeYL+MuGMA4Wo1+OdXge+vjljr1qMkjO2RsbRbx/l
kLwBSTN0E28LXE+UZp7m98gTiUBQUdw0VS+k3zgoozE0Y7PFaZRR7RCGkPBAFcY6
UBB/YInKAt9/UfQi1VM6pUxcg2XFdmIOMFyxQ7Ll40VbJXS0veyaI6OrBWzxUt/K
URYC8eb5UPTERTbYEzSb/zivHIPzirseTHLcPo2/g1sDW/1Jvo1Gi9tyGrOAbuAE
bEg6hY91GzucyuZTnvzSzOOK64caQX9dv5LJFPNSHWIwRL+s6oJpCbLtkywvPnzA
4X0f3dBUh6cG2hMDyXit4xsvektlsoZhOi0aoeKthlmGRFPXC3ObTTn/ZZNpr0sy
rgJ2d6MIwKyMr9VUVuoiC2eXtPiUx0XgfGXuqC+mVG4F61qvUDF8ypkZ/x3h5VFK
Rs7JXKUThlcykE6IT9WetL2QhimR4S/Dx6nlvH+7m2xNdMjJD5yLg4rNcHIoqucZ
WlbLAVI3WH/GocIAnD7l3nymAdng+vysGsSzF7DxIVO0Jf+CR4FV32e20e7gZlTm
zDkvYdLNs0TMb7iUTRoSH6qglTHlV/yMB+5Ko7WKFfzwehJL+AenrdSJU7n2bkXS
/Z8L1D5nULx2EjizV+nsR7LPP/glj5nu7extCYtVCLb3ampnnYj2UHeWOTRw7qGR
X96erWyPidFDxvA8shfqXW3j7TMoNWi+uXDY8SE/l+bpKYE9/61nuQQJIsRc7rQi
kX3+6afVLevZlxFNZOeBQuor77W9+7JzrXD0Wtp+9e+0RGTvVN+VpTjukOzqSgVI
mbyBukTBRUyX0o0TQzXxYrW7FIvxLLMzBVyPf9MgpyXphQZMG5ZgxBfU+/u5ZGzF
UghYxvYqXjVk1zRcYlmB1Mm1Tbx9w95zSeznE0YwndPNZNH5WM6faWc3TX0VmJon
QGAIHAnGK7HX+ejI8X55fiWKgWKuUExgwPmLLz0MO5sxMQAcrU9gLypL+Zfcb/o5
g072oYA2VXsTb4ld2MlhZNstQUSYCDrG4umCrCBLNtBEp+85FTts6azxAqacknip
YY4Mpf/choK6f7ZYmlkTfcpQqdA7Ernk+j7vTB+ChcUArMNupdwVdbOXpVcT8edH
942PUG3nUyG+FGoDW75uknAuRAXLGsP9py1HBgGm2CMFvd+R9YXD+dWPM0odM1qX
c+ysg4VelDdif6fkuQrGAM04iKBwUP4agGOGL/vsuAsXqGVeTgr1X4dENKX22j/j
/Viiq2BOD3hdLYnaEFOEUHQzmz1mwjhcw/vKFV7DsYMB+7qqMBAk31RullLOs5fF
f7qtdIsJV8zCK4DwrTF8PkKBMiwfGVHMBdSvsNc0bdj8bTr2vq7/orJ5VK9X7JEz
sF5kb2GhBhJAR2uFvpxr7OIcmV0ljc5bLw0RTKLJUhghrmYeFMGYIHaE0HUG2tQZ
LpMrmEGtd4MU3eJsX78PtkCadYIjW4cIqwgvzPa7FAC/gt0NQldYKyjXA6Oan64W
ZFD3HbCK8qTRoKEnpbir52pAeEr56bcMGetir79cvzz5bJLUEfIrfDf3VzJZ+sso
qYnak+bhSX7LAo1lHrl/Hlz/TKwUmrrrrDPlc7jOEdYTsWJu1d9DLiSOc64bGBBZ
zmkdC8Wov6eo8fA5zrCCFRV2AaDirDipce7+cJxybWS2/9QHeBtVvHawwH8UDwWj
0CrtDO8EdPfIpI6wWj32hDIsoCPF4OD9cmlC4+jHKY8aOBKqHsyLkjHGMEhrlx0F
bf04WN7bLVsMGxMZ1BZLbxZQ9cCXaVzg4gGrs12bgOaZ5uTkiJkzMuHsUVbRCIGM
PEljU+9+2bYtawlz1N+JlegOKQKqBufTSFldheTRwJcjqIPL1JVnBoJK+nlluL0O
738hc0kSCt/P79frLq0078UB36JMTt/ZRG3cwy18DFqAyxZ2iQDN2R2vCUgA8UJm
H0SbhqsUrTgaUdfeEn5yExFfCwZ39xjZlFRj9ncB44ucXCugWEHivejb94Ng0Cxq
GR4yRvPRe2ChM4fr4C31GG2/YioRMfzW9bKN57f9Kw+MwK6H4HpHBKhchllEfUy4
TwAcsRW9EP25Uf2WwqpfaVG/lJd2/ox7K5DWDckD36y5YKWf4pxC913naJxQI/eD
v/98SzzfG+LHOIrWOxsGLMsmkJNjE2oZaQMuJs2Os7dRkO8Z730yMDQxncW8LuoP
LWMMvxBz+mgq6w3poN+P90Web6bJ+OoQP7LxoqZKRR1fy13Wj3yYL0YHc6uq4OKT
KjgB6zWcGVtT/bIj5Ij45mvEOq2GvVlenKbmbQFquiZq4StVSbYILzTzWrf4kWJq
l/T9cT0Uixa3a+7lWD6HZ1ymkRpRkOLwlayE60+VMZGR767XnuU+xs1WrQAj2LqX
aMXmSn2JM4xA0oKG5dQJuU2ORaZXNDgAh9XKyuJBOYs/jXja3/X+bYwr4nbX/g6i
razX46eIFGqXXcYUkxDsH0+4X6F6Wg7N6+tlCsPGjfIFalT7bRBgxfQsJIfuTvGk
iSqhrpK1TdFclbKx98TVOxKv8LeVJ4T4JJkBKATstTT5gT+YZXnEF/qyzlrlHHiN
Zh7MNABBCMOVu3vVMn6w+9IPCOVneIYHJSjLq6uAYkO2lWsLXNgvGWt5xJNRU26W
fYLCKznWIaGRCINmOwHCpZcbjJy10uIBwqcOXzY7IAnROiaSk67thv/0l1TM9+yJ
QU/ezvxFwT0ZnzFttQ45T6+k1tcPIwPlrurYambTCvoavMIXz5C3riHwh+Xul3Ma
16YbWp3jBLGVnwQ/TTcx9OYUZvIyjAFX/uwO8+XptKb3v7kV8RBTAoOfigG7lFXE
HJOS6wD/E4GJJ7RXyRqKvYeu5ejb/OqpSmUAj2UgWIkvYMtDgYmXTv6m3wBXUT2w
wv0TKNQvCnD9KXT1wfyzVQQ7tTLM/EGE5/ZhNk+SdMpkiNnb4Jr0Thpz9FVvapGI
T58dyxPkMgr33itlrpJFsNTNXQGSrLCT+q1Yoqv1kTEN1yDQklKx1OtUEaby99kj
IVd9cv9zfOSEELdPLv17t6sJiK0TUNeVK43lcrpidOYA6Sgd9ha7LhTPWtYCWjKz
H/RO3CJZ47XBkXJI5dq8Ty9yZvJ8oE+RxkxWIq2Z4c12I2jxn4o65Ig4xC5gYTcR
fklH9P0kqegOGgfjlGaJkm++XieqtUgRPfzUKWpJwHFInY7MFAA+7mBum/L+0JvN
uAi2WQGIeNpXvznEjrt0UPmSSkvR+OTmOzpqvSpQwUaLVVAKjKzvTUJAli+hFxEo
LzHx0WhhDwNwql+d9CB82XB2Ri3cPVG7fawlV3KaFfsHCYaGnhNpE0Oh1L4yJzaf
RbaPUkZ7eppRNSviibSjK+MmjDP6AAyhXTL+JT61zk3+VJAVglfNAOKoaJhNCQwa
Qkx4xpFn1m7Pw0nf85z381/eIhvvNvdc/LcVTvfskRcaJYbthHFwQoplT4m82Ou1
a33W+PaMuxm68dgSPwoIOFmOpzdfoS4Nl1sy55DJrn8W20QXpm7rNChBDeHj+OKL
luvZ8XQNLj09TulrzcjgkFhXWmesQw1GKs7dBeMrlOQuBsaqRRd9aZCMfchjwYhm
oM/nteOSNGH55Kz46BEg8WBtVI83ouQ8sx/iHYM7j3Od8YwTrXpVy6mOjq6/ymSO
R2ZDlfpymMdsLvsYe7q76bbniI8mJIdUf144+WmHK4h/sTszJgB17JHyPQ02GbI+
jb9gIPnzjIRlrfztNPSWvKTwsFHYVUuEPCHmkVqit3Jjdifdn5NeygkJfis8xI57
k991bUwI2Ker9fxUW2nSEDfqbLfnknL7DLsaV1Kj3xASDti08extXdxjqwP6p2YW
rvNFjwQ+W1g57/bT6AsXNL8/204bke+W1GazgRMRYU+qWyu8SGYI0r9NAXio2+6v
CwCT3TbmAQWSkdEh35EwJ6ISfWTVnfgmThjUtYrvr8Paf9q9V979DEHqjQFv/3Eq
NpR1icRwLL2RbKSwQl9LYvNGcC7pE8OYnWichV7wjuBcn9Rb8MbgZ7ZY8D6kkaCX
Y+XmSKLM7aXC8rr+BKeKztSgkpT/cqLLt27qcaFc2GFellSqSiD/wwpyzdQknTQJ
YQ5syC59rclX7GnMyDIbzxYFHkUualirwkibCUoCUYrlSBcCVffEW7GA2h61dJ3I
zg4TGp+9ORCwToZ6fbi4Yrf7Sunr29aK7wX99dyp2DIHGng3JjyvIvd1N6Ik1z5X
UEe5T+BNKyVqpW8/7VIhPcYizNnXhJ7NBxI2AWXm8MHGsV9MvVH93fQ7/TFfzY1o
XdtdDqBGOHmGs87vn2H4hDQ+0m+PM7vycK/b90K+lTuQnszvLDbzSn1qOdx+dq3F
F20Ky0jbHlaF66Ue099DdOG1Z60NBvI1jBsCnFVJUQlxGw3CTgLIlqQTEKySLP1o
wVMi8zx42r4ccvndGw5/OpX+2x63PsD2nTN8BibiA7BiLLUQDta2ja7HcgYygnKd
8JLY2HXU/3hSIUZcK5vCpSEi50Lp4qNim18JQWvRenU5GZLSG8ZSZDHDkTmMf+iA
Gr2bLpXqgUgU5Amv2CM/jyn4ubXK79PnO/W/6KyYW/aKvFAg0yY3nxrgxJp1P4Fp
6BTBuYBuntd5VExY1mvxtn4zuQBQlqKIRUw6kkfi8jJtfFZ4PEw17EvuO8i9yAFo
qNJTd3dV98PJGWGL5Pc668K98anNE/zXOgWjTM2RKG5mD6GG9T/TnA9ucK25xrH9
RHVee8CFJgWU88LbIQm5i6nJhN53z7LCr0Sug0Y9qSgYxwzU0dacHnbHgI+qBaz8
IEFLLVjp+2Eirw8RJIFqeH0yTChzkzPDnvzmrsl8Cks6dc7zYJG0YMxUsrpjuYGo
I9tZ6L+byRhphknd+lJsOkKlTqdeqtwc+QGZK403v/zlAIXi58R0V34XnGp71Odi
R0iOYpVtkqhhRMEMowwkeKlgLaroQBnmysgQ9WndSrmVRoyxPgYKZoDW3iDTZMJN
WP+fxpI19tmLEGPs5neBjDKRv1ERkWoRQunqwUVjBMG2YFzW+wCfkORtSlsFv0H2
wsSYJcjz5SDdRvMYSnQR/+DytfvFZbAtrxjqIjBD+om8CAVG3mYOlhphjRSwz4Fp
WMre7x0uCK+f36SGwvED25Cw6zYRUyhhjHxd57Zh9sTO1UN1p7W5iU/F8cuOXKin
Cbtt+7nXEFjvig6+4BF2GVRx+b2AFOB9d3zFbFJJ+z1q0qXBkYXa/+oSPV/aGsk1
lrxlqVWr5vAR4ETZxobt7ps884iAZfl2Ai3OW895gylsNPZGybpbie3woFDeuZz8
BGZPGovlCFY014ESSoTzx6fsb0xCb4G2gDD/Y4fZ4CJZ5AO2jM21ltWO9jtYwsQI
kY93eLoCgEDtDlnUhza4mbX9NZYmNL0ewNORjDOpQj0b5031vcqjAf/ni3ARkWcd
R42NAdklCiNNuu+Ipimv5sJYqnYQSm4DyKDziULLtD7WVXqZPXeNPOnDGIYPLtxO
4wjSRa2n0FN99l1zia5zqMsg5mMYD+S68xHWyX6wyN2JRKqN2vA/JgICbvM17z7F
GXYGtpkqJstX1P9dKt8OduXBZuNedkgG7p5KxHQvoomdEvL/8r/vwSUMJk+KhP27
gDK55sQ1GbZzqU6XZ9A3iclTryHOuDCw5hFPKot5Uav8ZVmWrruELEqWhFRO4E00
MljjmyYRcVDUVh0ZsEcwaCYZL/9fnqezzADYF23tdcpc1+ZFjR/G0WpABlJ+ttwE
23EqcmG9yxl3yACKoR56tLNpnDdtxTCnjgTnkdpAfBaT4Y6BNX8JZMntj+oasnLh
2MJxICxlEcqULTLnxAx6tbBwHjQ17fRk0Jjsv1Cb0Ig22eylAH02sx8EtXhOXy/z
/gHTTJYUryyGkPrwn6whBAnTx4vGqhFGktLrPmy1YorJkzoW004s8jlydfOEAtTs
gEEWqOxS6vTbOzQZbub0M6ry1HbPqJnb4+KMG5cBcb4n9843qcP7yrYdd+5ecMIc
KsWQks/2sCNjyNfRA1E4WR0pc1p+/Ub+6DmVniLcsvoB6vOlWYjFxBk8/80TW7wg
s9GLjcgzqQpnue137eT1J/lXL9C8b0Rtv4vO84HS61eX5xUzy/VW0IMQY8PXKyfy
5Ng6S86avkmZlRa4L3XTaJGPGRUGkfmiD3V3CS0E27GyvrUwkr+caaYFbfwq0HZU
AwNr1EaZ8EY7UQkgy+a4PPt6jv3whW5Tolc/VprxUJGeNOKj/rPwZEVaRVBbKUgW
3jv2FUa50A0FRCkpSruPyIt7AF4bm8RCNEBqooqIsKZIF9iu0mw3v7wvMUUD1pBT
s39MY7f4ytAA+iKh+oJBng==
`pragma protect end_protected
