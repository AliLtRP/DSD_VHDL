// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MP0IYC/C5hgjA+NJMxGz57h9BmWqZivZzmchsHA7VRo11PSEVbIuKij3bsU7A8X1
h2cinm9XySIoQVEg8LS3wOBILS/ZvhtSWDjArUvhMsBjndCnnQHLPtaHmmovrI/c
OybzpF+KD264xvLcHTZOJNvuOeyvZQSOg8LJRyyMrFc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
Ke95sTpFBUORghSZXP2OzYK0AGD8W1VZ5kr2z+mi8ul28wZh9w5OGlwrDvkRj6S5
ecRf7yVXvmOOlBOd0SkGO2O8ckaLm30zsxp5hnsLuOGhVNK0vd0YcPUEWpIYrFSp
3/GdI2oogpb9GUDkHYt6tsJxi1bFBj4JBCJUE1cC0SfrH/TO9y3GY6hKSn9bIyqb
9YzJ4iBd3sJ4DkWgk0KBVKIOMC/9JTpgO0e7W25PCp78QHlD1fgVe7A1Qi20Dei/
iVgxLcRowHdpnVb5z4vuhn2CwGg4zdbQQMFpKrt287KZpJ2nJUX53uj1SKbLJQQ2
amP5i8g20QQQhOpWDgDF1Aa/V6mlDac/mouddeTHYYDpMdrmCF6qw9TK4y9uWaBF
F1MnylwAt6bwL8G55fdHyvRtVgwjFhIKkKliuEB7Pqehg/L8iijmXrrMRipHVmXB
hK2KresnJTCCJESHif6IzOSLY3wdIsVEJA2MqjOJbi4mnhAnCL3kAAHUj6YqTaO0
CsAWGEZ4oDDl7fudZkLgaHrAyq6QOh39kOmOB1oirGfWrIZcsvtB4QxJcwyfSaUV
VDY8qxZ7mTgpDwuIDthZsWJDuq71rfxTygbkGIlTBe0viQK92DKzPCosHA6jdQTC
ij24k48CAegQtTdVowJq/o3TWGbDjNWxN+yo/SR+C7M9D+IIfR4CDEGxPENrIKod
AU0fJgYAreUULoBsnyWEFSbZ6gVuj9MKoC0A2YSWKfCroAJ/eoSGYXrzM/fQuDjN
3ajm6TW5ZOkoNfhT3fagc8FXimFpXXHCQn/n8OX58FVt45Lgpj0H5Q/U2VOvJsf3
/gZEYwxudgRL83dUAFAnF+pe0YrxwcIeyKTApbRVBHONRD2okEzMhxyLUgrNLSqj
jr4A/CoI6/HF8AeZZDps3nMP4lDAUi+aJ1F6BhEqDym90FzGTvdivbJeNR6K+zOY
1p78DBaefAb7DXMjljUL7pGL/LpYJ9U5CTFN4qwlGoJBP44kqWtuaLjIf9VdH9hR
IcFT1gP6qtSHyEjJvI0rvxC5RVMJr1ymogitxokp4ECiknyzyyA5c3lCB0owptah
+rSY1/YgUzgxWyLwo7gBUuZ7FHWJWXl+D4L7uTIpylsTS3gPVZQ5gZtyqiJIQuph
FZHDfkan6n6079Kv5E3s/k1LPRiLcxFEicQCVIzLW1lzHsH9rucoRl/5bFWutkYp
rg2xxvWOloQsCPbBUgmHtVnyQboWGTTdD7WRoA0sxILG4h2orhj6arG1Vx/Mc38h
C4tAqvn2hXUw1VtDBWevPCDY/Rm3gR7US4a0YbJns4xNlPVKFPrrpoA37AGeebGT
VNwPPFG6rSlgSWDsdPBz7jErkG1ELz4h9ABgjmWdwX3t4YSGIWRx+yE7KVgy5+gu
ej5iq/MW0ZNhRAOD3Sm+0PNJvAaln/pNd5XyaY42bSq9whEqUIhhYaByU0Ck9Mag
t02uPo4fCdF4eQApWbVT5KsNTXaf21DDOYnyHnGESPcppOX84viaiL/Kney9RAQO
zjWuONGbewvtrj/s6sDUYfTR1o1m+XcvWyERqVj37X2R5x9qn/MgMjk7V8ClXpMg
hsDWB75Mm8uV3ZP/Yj5z1nZCRvXzLCKslQC+5D+K9wK+HycSeu8wV6kVsO8Jef90
6IHAFM6u30/6G+Vlhw8RXjUzJuwdELsTugkc9wM73X3zvPp+ybRPwG0UFF208OLP
HIcObXye6vtYR1VrpsWVsVtycQ9gZoXg3L8JfHdXctMfWuBbbpkMAIVP6wTX0m0H
LWN6Wp4I/4mu9driOdmN+EPhMPEYNodgcaKAejJqehr5qsTjsNQMVy29xd/ng2d5
AVcQAH116zmAxuDcBvIrlB4KnzsPfQ4RgGX39uqOR5LUOEyc54gl2uX23wPa0mRP
FSWABpNARuGOBO5qaU7YJf7/O6QApo2U/c2Sf3DJ0xcF1o9lSElRwTSYXq7BC8qM
rSqGUNiJB3f+IMC0XNq+5X8ziRNWeRfkpdTXDKIS3aq74/RCcK2NtYAiDbxkPScI
SLK1hpQvluj43Zum7I9T/iDg/K2zNtgcO6Rq42GZXBDQnW3wzRPD0kNn3P2dotkg
4DllQR8mvDltt/AajXa2fNZdN+eA7cAOQ1/9DMp37j0GMnQp9uxATKlp/jAzWQ7Z
DLzbm5lhaAZupBHuteZUxt3yzF4EU5TD+xeqQHjmUDbm57BneX4n3NmW7+aDsiKp
YeGzq8wmWEE3x6LecMXePopOLP7AAlksw9UWm1l92d0+FCLgK1JfwjMbSAFRZnrX
udMAwgjkk1EybxLdnn2eZklK72Y1gjIz0flutaZm+0JaEN50OVChKzUWJ90fFbQ5
+uYYqJhBavpYpac1Cj9efIPJxOKcX86alv1n4+mGkfzMLD9sWo5Pc8DkVD32o7jh
1Ks0pZWiLDplRWNG8Y/xrV2FfTxm8eUyr8Xis1bbXNVY4kq5SOXumYjwb8NHHsou
7Vse21whrqagTV6AgLrXsHS3T+1j1uwP+GVj13TKm9RCLTi6a9F6t2hAw28DkB1c
ZB+1pa17aP1OshXITK80EcWPbSEDnwLwTDZ5m80ATPxHYd8h2JQzUltBbrIqF7rS
mNegOmLIDLfxvMebFSufV7HiPURQNk8U8sy5ElIpkQhsdP4pHfHAQKEbbZcbjc7T
HzA1UP1mQU74Yifpu/QaPIz0BhPpJXfKLD0QD78Admu9zV89ABI+6PYSMQfNavHq
VGHtdYD/dA/6Z/szFgNsgjgC0y0SJRJYoQbzGzJOddzR7sEtUz6MhJosCRyw9Du3
+VZ+0MflXkrJosdr1fXZZ2EQ4j9uD/m9sPaYV9Jf9odEjHpvsYxeVzRsZoCLxYF/
OpcnVAxJIufkGobRZgr7NyaqkKOpTJLmBD0JENj40j4XK6ZA2b0ZyRWzuZ/tZjgB
veyVaNQb69RSaaozF7PQYHLBMcXbwRvIYHWW7+ZOyWGp1RMjG8JZJ/lISn0poNio
SHlB4vufs5g2olJjgkSwTKU69MRJGGbk9WIW9q9/3m3WZNm4f7LGVEq5SBxzNUs3
2Rz1anEf7duZ0Rt3JW/5KP8zk/fRMnj7YFW9M+RI048NvUC1JNwxkuw9PKvXN6XV
pBKa7bfyE1l3kkP8a1T2ZdfRD1FfPdBfMcRvXoHLXoDtH3cXmU05AL+fBSlN0gul
Y+hAAod6KXOO10s4D/qpGh5dBV4927nyOFLpgLD5c0ivfqQUF3lNoL/AnLEgDYGH
02IpOjlBLZ94sT8uKngD4Me5jO8ANMIVEE7Ihf5kpbs0kZgPXPByZzL3s68DxLYJ
/N9S8vtrLQWlSCoEusSDpqoWgmuBJRVWMKAs++b1U3JaCicxUnz0UvnTo8YrAzju
u1gF8A/+1dlicEkqp1jXccbeAvL6epGIDr6ck9EnCa4GqDJNmysZPMXk4w7vH9b+
GHSFNbjWQaB1Z4vrDKiKKw1m9cCVAk0VAYMiNG+7F8UrDrM65VszmTCzlB0G8Qd6
GrRWRBsNpOz+zgwiR5pb+EeTjxjRaqfC/XLLFjzs0o7QjjBy9d4qrZsUVBuAyfJK
z/yp0+xjZGnrxWZS3SokgU3W3XAYw1vOL7MegaN5XeoHMzNBo5Mgh6GJymAQFhQB
Qauj0dQ6KubaW+1aOsIN2/rrSlGJP9/CVTZcBjqD69uSuuos8b+TNp6BVrOQSV2B
QTStyCCPQSzto220OVu4He0IbqnOAGTsoinLpMPzk4dKBiKfTayd5dGWjCXZh5Ka
j6++BdhdXQehLCG6Po5fwWGSWLtxkoAhQw6k7fVT3R1RQisfUfYj8k0TY0WItiH4
nho83aP1zJ/2g39PKvX4g1bmFimOQBWY0ZU+hqZY2qknBPHs4to/IpuDfOT+gvpc
4qaIVKt2LzhkyF8vXkofkmcK4IXrxI7oThIhJRbSjdwfrlZ/BKN9irmEuL0wm7qB
EpKst1vT4l7i+UG0J10VfLNSjSctGLYF3FBJuRMslyKKPsIrr5NB3IAVGmlUVIwp
P4vGTWdRQlFor/e+X+yAZAGlBjsERVTMLcDCZ+1UzQvNnpQWG928yv4n2TrZ3CQE
FPbgv51UA4SMjcljjmQeGHArCVbxYE4NGb+KLFSNY89l20/Xv+lVirZoB4HXt64+
f+cWeatKpvbCzY8M2phACLwKDjsk3V9SqFoI90iiJvg/a7Zzc620Oq5FjJq0t+HU
uXzcmLboz6fRPLVV/GemiLHP+jNJNug+HWGEQCD0kRi3Lnb71iORypAofqHEy5w8
7HuG0I0CoozLbIAf4xQxKbG2iQm9Z0Tz70IFHSOSCkOqSJywwfHqmvcCet+MFF1p
rLybRXBpfQzlaedMN29s1jLNQJupmUDO9/Z96tXhjr6amlWsQL9XpGezVNQMcubu
I0ZG+NZyg2AoeGCsKsUM49YQ8kXq35MnSuXTcjUmQO99Nir6H15X77PZhnv6Sj+t
8dDcWdkE1tdiFsMpNjUIRvcgHJiO9EsvVqYIMP8M2a6ntHNXdclLqeR4bgf//wok
IBRuvqN2Uy+gy45fMe+Te8IJwEQePA/PWyPVK+Zxi4O9cNgXIlc6hRH/qRD1v8lz
TF26IVtlwDv0zuARbyY3K1RpEBM97d1U2c21iSQHUlzBDIQRjBcRrPHURFjE9NHE
hfB3xs5n8UkgmNIxkaiQyWMuIVYcVlcFnGLDN/gHdHJebtUKf2BsDVtJKBZYWxKx
oiVZMJvZ5Fc0WbGk3guvXwzfzItaU/QA9lwYV3Zv8t4m4clyG/WA/9UBsuZxka7U
IbBi0chjRnoLhqSpvEbBxXCj2s3TJFzV/niTftfu3FIxgl1x1Jm4IAdG+nJqhFwL
i+MayzJY81noe2a//axOVPrg8+RfnI26ble2VYq//+K942rZq0wDXqoCw9TijcH3
Bkz8owVVqs3eHa/HQ/0/+5byGAQCLpRW/+qvvBgi6F8olrtVQhAQcg8OL8o9aFa8
sBNi+G82tm/jmMA/IWkyGcTxL3UeXicJJNDOf3fQj69eckHDUJvAkpK9i18gqYEG
VMEKLHFrdofU6X1VsFfoFiz4tGxUe6bO4qLOzyIIqQjvFioZoxMIcwdfJmhTcc7x
LujpsTFNzvLkjlcjrAxGsHCSWuBYQwhLABU5cEnwo2BZtLBo+jRZAW9o7rjDyLP8
kHOYWVj9XAhOaTK3DWEWs/8JU3BhoaBGFW9Dy99WCO4KxCnZMN3g1Tj652S2kQbn
HwghumBrRQwEaOoPdHp/z3omZNw4J18oJFRbvdlX5ze4Lx4xzb2nNWluTQr1KssE
gnWTwej84Hia5eAGMa6YdxR7YW/E7vwGFFvUA5E19f3EljyKMuhTk0m/TpcMcD+w
jHXlEpmbKIZE6HIzvX0bs5koaYAiHjO9gbgzS9GxswdjRQ8MgrLXH2Tfcb6Gi6dn
AqEOQ3Fs0cdly4GqTTnYgQOW/ZrNOiK/nV129NrazavCpYHD4CPWqMdoFS5YTXpv
ySW9pC4WJ3PnzdQKxI20/gND1yqpx1m0TfMiYeHSrOOz+AEs1mhgVFpit5Lz+aue
47aAkPeaHmnJWWZf4WU5fKA5fQpb756LdIwlCjUeHo/v5JbNc7pWczD+nXl3JN9r
XkZU0L0OSWuHkQlfOVrAb3eNl0J8xsqI4fslX+S+60GYtCu3ESsBnJ0A+X7hhM18
t/16k4iSYB7OYrEpGsiMQQjzQ8/YsAdicfCcuyVhynOPDbYfxmpAGb0PF4F4Gf7k
or6PcoFMpqNwipz+XiX8mQZyilXYheZuhCooZn42zK9+ELPJKW7oDMFmXT87PTzN
sUI7yURiWW1Mn5/6YUSh2z8mF4t+AkDUgyCiLoQY33ul1lLTvL0lOEydbi/2ZYhQ
vM6HvJcraAL6fDggFLg1kpYrGXg9V4SJIbTdVy9l4tY84zKhPAmott3wrWKUZJLK
hVCev20x/lpHOs6Y95+RyaxDm6yORI8KSa+PHbNLMsoEbY/ulXqeo4VskWIrtpCg
TIy99A7fAuH8xxF1+D0Da1XJapYhWdfq6PEVbDn8GCmaAqgLZTpCWs3gJXkeR7Z/
zuGdl3DnQ04Nhh48ARo5vMav0zLk8pFa4/Q+FZClUKZwg2X1s0X/C+hEWSNzwBDB
zcHuJD7x7JceQ204ACdY8Z/Hdc+OJJRU96IZg88tDykkWAj0pH6cAIFULMdBhGi3
diJPngqzb/YnFcOS4FqJfjd08sWigwfZNvfQ2llXiYsgkyEZwjOfGL1ru9CyAuSH
07q0ze1577D7FHUWDoEgALmw0s9VZMcrWhJOdWw+NJoV0xZ620+PA4KmKgNsSHjs
s6PuCtKwwueBqobYmWH2znv1oxMggk+7Yif/OFUWBHBbKDKyTUlaYDWOf8ylJQY3
HLGLzn8r/cTPNtx819TYPN5MENvyRwai8lVAD2mekVIWoTsTFn2y4xZZ8OzYmd+k
LAyRlH+urplyDYXQHCDTJH9vvI4reorUgWXzxPcqQKXmRGyRsDnJKzz7omLZQIpS
WjemkHVQIRnubtALaFv+IaUwhsXkUEIiNtKQDopC6KcAOs5rlHylw5TUYj5n2ZZR
W5YgSe04DQlfYRYvC9Ra9wNyOCB3O3t8OML/ne2SaMYlh42fEEbNgSXS7QzGPe/Y
SZM/gfZfAa5/BBLb2drBd4lRnzMxqs+wWepLpAerpDjEWgQyupQMGKXp3svNuW67
8lrI1SSOgmbWBg5ysQulJfLvqouhF3IMnKjhGr2To8bsSnu53qbKuSmxWOMK3vle
ilDDKU5eouwr51GhHCh+YFt7LE9rtilG1tS26Ohj273OyTfvHSgdP686DhroRLyH
5igXipgPsi3ofVKKfPUyYx5Ddq0RFXVdL0twOdfMhi8P+lgaPWyvlPV8/HGaD/S8
u1NpGV4fy8El5/6rDmcGkMxVLx0qk867IGObon1uXUllPE9TQQ+u0aSwaIFTZbbG
v6SpYUiIyds+qx1LY37CP4wYBiib265l5FAwCaNuAtRppFtnekoEMMFuCZpRML7R
3xVWQm1n0PtZzASD+y/lluspML4iH4KWYUn0ME9Z6bGrZv8RUoRrzZrPnAH6GDsU
3nyEmMZ6LgC5S6J2y+2rHGjqFLxJNq3z53SCH3DXEwtrzHCdNQ1x6de/3ZtbvRM5
vr5Q30ZIXxaurs/Mnq276ceQXZo8qAtFwmIYMRTtk2QHmm2uzLrcMVwQOEB+xuye
cdUYQR81Hr8jyI6ZMd7d3yJlFnqWJXCixBHh5DVay++F6ps+mIhrCXikA33Ac2mO
xFjXGWWNTIyXxiaV7GuQYGtUNgnHNGzXmTwO43q5GLlnTkpBPVpNmIqpMtfSwtY4
FThtEzi0Dm317eY2NtDUBAWf7PxybadZ2YCJC1/eyAHAdAIzHlF83WUr4zJxdLGg
34v9xrlNwrbVGKeNgi181GZ60GSreo6pW5xA32IoQ92GpcmUB2k8fWx2dguEPDK9
BQ8vCbS6MfZViMdWWo2N8chFykU2mclKHq60EpvGc5+8/Nhf+E+4JBRPiPiXV1mZ
tnW5sQtcYTriWVTeDGWiWmukkq6Jdd0ipHuVjQ2L0I+81ojGBUAltZXhtVvaAtCL
K7ra0ukLP4ascMUt7CKhCdnbUUFdLYe1HUs+28G5W/bUaSdwUhL7TUjS/BPvH9YG
yIhI7wKoud5U8b7Y4vV2W/bTfGI5PSta3ijbY3UwifXIG88TY9dHQMiKxBHZEHct
9N7TsrYN2cED8LiMRrqf3gqFw4iC57IFnoBvCbtvItQ=
`pragma protect end_protected
