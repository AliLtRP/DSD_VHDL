// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ltlA1rYmjU6fJ4eZvTRSEouOBZfGCpxeHVGCkgel9weB1QGMbwXhmAkdHjKl57ak
X79xClYV+0whcgNt7TxaS659g7u/+BnqQIOuY9OmJBUk9U6wEF4eohHIaM271RaC
2hDLmZjNzbFEkPDP8gDsEVegfI4sc6Rs+qqwbG01TRE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
vVDNippFN9x83oiQaYgDK+vaYdM8kvydAMXxHBEGpkLDBPGzwWzMNW1xBGa3vD8m
eIKnYuqIMxtV5qusiGH0yurYxRozsW48ANUCr/UbT80rJW9BUW1Zg5eabZxYD7M2
33vVnXHRsksFEe/Rwe8oS20YBcIf8O7a6bfVpWvHXfmcSGUR0RcEZg9y/GdQxgnt
zbZRl9yQpUkoh2gs2ZMhfzdrxTnPv2DSGic1allk2V5sgbJquzSWCEL7597EDEkz
aJpQZbni6LAjnNlntGuLRt97AHmxaB9Dg/kqmjkJe4SnoR/FeQh24GHqGCHSo0Pg
ykfpWD4j6qKjRnAo8MD0WckBXxzrQ6nnTC6de/MTjfl7cWnXX4q3eW8zWihRbtya
s3UDDoOzx1q8xLuz6r5DsdpmBC0Ml1+i3AS2A3FT3dKPZSAkBI8ud7nalYx1dAfX
3YoCw99WRwciWr4LmLqMVitVYNcZSvoKlw9saZTnxiiW2jZ5DQ1CJchXH+HHK2MI
bmMSYwhYyhUcyzU2JKztdun7j68DezzVWh/J1PCA3FWItWuepMKfnKxmHjKoiPC2
Hb2WM/A4lNzPQFE7opMpHHipwyDIraCaVXEEmScj87UGrJb3wtdl1FyJmA67umbL
fQ2IpSF7ymjjJ/GvWQA1DyScVui7VHnyrp7YHVpNomUCevPlUCWLSonWvIKrsCB+
6rpqJMTe1Uaj2BVoA9Fjj+GlGRErgtNbt7gU5iH9uig1wSDzHbOqQn+A+3i6e0AL
D8vYpJ2v4NGBPFvssrIDYjt3bbfICQVsj4KlSaJRqqGrIZ1uDhr/pXuFk3uEQYA5
g+uz/pjyEqrV2z1aIfJiaNDCWNidamfXLpit1niwYEsoK5577bzZpkJMZXUpmWlc
rpagDDnsrM+VJFinPLP5n/EMIj1UGEs4JYJUECp/QlbtR+RSRH1umjd5M78WR7sT
vDT2Ixfgy5boWWvarAj6sdHInrNsON9B5w0Pkh4ki+6e1X3/Es+MP+OQKpz7Z5/7
TFkF/Nbu3oQfigM9SsZylmD9vIOBU32pOnDKwFz4MGn6E335hWM7yBbwLgla+tos
fPKs2QvvmQDB2kHRu9KXnOagowevHp6PwGenotnimbb7wPScd2rqGoO+uMjbftA7
L+ovvCbUH5asx5VAcab/zyyICsD9ZVAi+7HLGsinmEDvcuBAj4hbB2lcfUmIdgNS
yvb6FeAfTGugJMMr5mQ4SGJhk4H4SCwxuvOAgMMVpdntFT4OHt+XcFwW3iwKVtwk
MXWk+zzt+7jI5GkZ9TCQH7UO/owfHTYjK3xKz/5wOv0FSJlf8op8RvPkdYm6Qe5j
8XNLuk1HJjJngWfsVteqT/Y46EPvULLfXavg8Jxx5oMHoWWyDN2pjeZp0K8WE3gD
RWzvqDULjv/NWjSiwaTpmmHGYyI2Fwac9zaB2heKxLV/SJ1+UbUl+UU1k/kAn5ry
W21vmMB1ihjQNb9LacmwD0kJH1UyE92xDfhfoWYNOOBxaeh1nT9yfgtunx9UyB0a
+D+REpxXIfUxzlPTObfTk9JmKUIGabZlf5shSGbJIDv0Bz9GsWHwWLfsUYSBNSvI
iU65C+yvaNbdT5xaop83MJ/5Ypxw5Rk8d70LMFI5yKbWwOBW/KFyxlcV9nJnIvpk
plL7arUjuAK7a0X22FiPGniVFjeByBT5YmVvj5v050980DTB9XiL/FaoUArGcKHn
eiFvvF7j2FbMAJnohca632Z69PykEhwv3Q+5T5oolJxv1YVh1f3l23NLaQuMDDVT
GnvNTxSmFnsVh5dABaW1aHSgFlH40ztPZ11mEKl9nq1ldWl3NfjexiCyOEa1Qcz6
NMj2mck+Snjb3Rb0qLOoR+KH+gGuiL0oduk5u+HAY6GS4l2XOA7E0ksGmpTkMNMK
Iz7O6Og8oZVLisygWwK57AjTVXVXaqlyVFMbK/7KiMfkiRdLoKui7keUtF8SaTQ4
Je4WLPxjT8EXGTf6npzm89+Dx76fJNVwcG6K8u19PbZlJFNUowZAnfqyT0sJ6EmO
RxqMQkQQncfgx4DeJsK1gdhzqQj5sk3JLH0Kaq2gFbJzjEVk8fYyu8jm85j+sxpd
2qouKNtHpWsqW2U9xkmZkD8fnJHzF1W01pgTzU+YEWU6Lkrn9tF3IlBjZo1bIZ70
KztJdKFIzUFdnq5xwqfvM6F/HPXc6bh7zr1YRU0Puve1rAjDBuEyeC5ZyHion+Xv
URj1gTy9/sO2RzmLCbf8XHNDrwzk+wWP9sHm24/Bgn9U7d1+vFlBb+geqhzVLak2
fSrvD1bRpfjuSAaw+WYIqMQqV5h9Pz0h0oy/Ep5CqrY1oEz4Y6psYEiFQWHstJr3
NMJmWVRG3vk/UVJq72gDMHjI+8mQVsUsBZBY8fP4Q0EOhvkMDQ6LAnNjmWxaOomZ
MpejxsoDrHe+9kvbz7IOr+zIJ2jpM5TPTKu2xD/AK0Y9dPKWPk3JMRSAQe2P+yR3
YSGoPH8uF6i+IVyXfWBn40QlZPnmhNwgf1SSeKQ75tcJhzuH/BcZG1OisMByN9nZ
ocr1V2rAATF/3nuZ4uot9UdV+4zGRHHUG/tFl6t1dp6Zl4vs8tvXr6hdBmGvQ1mB
RvgnlVtOibaqL2LMjzGU91JThq4aueECkoIbS8lofmQxPciX0ePm5kIIlai4uVV4
+y6y3uUERac5uGCyAkpFbY8bN3NQdHTahA+PoBRs1sWu8qJYG2c77YOrX1i9+Twj
lSDnZDjjab96MmRS49tkqL3eJOESD/Y/9ssywqjSStO/HARwCd29Iov1eJ/UGWOv
2XDkHMPg7SpBUl3Yc4xPTNriFxbuXzqaDA24nsN/WDU980jPHj467JKx7bwYu8zs
1dy4qYRjttOLI0phIRvnN/iVI6PUR4hsNGh4AXdDvnuNgdYxA+/24ugNFtEwOfX5
IGxI4fM6fBFPSDZ76D/DC3SO2gDN2E2FwC8rZ2i3nkvPzu+jjr6JltkZGAB9Xpbr
7kYptK3kxGpYHy3e/hEjNi4R2Rlvnesaxzx3RsMBI5Rqy53WLC/nX6A+kLDeTPq3
7qfXiKUBBumVxMvzXjeD1lnuMg+Es4u4VOni5FabJKP72mBuXXyTq61J0LpCNyZQ
D9sg+6UFySMzZ/Kge6+82dUBE1BRMrNRcttIyRHS2aCdK/6r88FWNCL4Vjo1gwqH
e8LqE50Cfsjn7f2mnRF4wHHJ82Wqg+u/dEERvR6gm109qVi1Nl77NcTEkpYS7PhI
9046URX+Y7+fu+FKo+WHgUfWYpoxAe7Oyjp6WhuXoCyLBxYp7TqVTQJz5l/FXizM
MpjMf5FULbnPDet6JrrHYaSlRWZUBngypXPz2WUKnxEaeEyiopa7SGdjH8h9Po/t
b/xmuLRLlJM/tLYqg8+lIg+61hsQjJZi2FnQpeVCe3Zsv/SL/3lyVvaKCStYCJ/6
AFUqLrDtoCrkNBZxEoNtboRliIxTH9k8kJfIz5uTTWfKJ+cTaapqYuyfrbeFqyDS
USFRsm6BQN2RtVF7vb8VSRMCFlhljd1gV7aexLBn9wD+M1ARimC5SZitwRvHkMQA
sCK/HmuS0YDKip1JqFnr7v3WnG9qD7g6eJvd58EXGWj9VFrMUdUoqtbmR+7cp00X
6p6OVMz8RdpBnJUPYo3QieGbdKTvklq2q51/NY4KP5/e8ZSKN7MfwWb6hndUcpV5
qO4EK//W9FVBtRVf2kKdgRdLRRB5+rtwYabvaK6AOBVqTzBiFBKsQ7goQCr/L2fX
8WvnZ2Dx9NA8kf+6qL2QCf2E4ZvyTcBUpBhN4ihvYw726Y8BQUS31yYPWLbBBLv9
v517hfgEmcnLbYmRmSKvLbYGIPwHWewvRx8aaD+lC1aNMIiYT7k3CRjL1Wyrle73
4zs5j6aevacduGSjayGA0LGkbBEGvsi/KkbdBeHOYxN1XfVmt/oFJZE+QDQmgtNM
zGDNc5Td5Vd1nseyGVH+67y/kPMnR6sGoJGW0C4uQROXDGpdkfijwK7YXmGookfz
rAmZJGpWMcTUq5lPnWFiIXq0+VnvnnhCccMacL4ZUfifrM+WdMg9xFO9c6KedA34
dCNWOLcEsl9Uuq+RFB3HAIAeBh9ZyiAPWKDFpwna3hHCRCArbf5wCn/YvhdsQyWx
O71VH1n94qdNUrHJ7wIvUXaMO3hSXUrVqx+iIf4W51KPdpfIQQvv6MidzqIYcie7
9uxubZdLnWb40iLM8+SEnMXonCvcN9ALUrGBFEBfzORWeWX2cWAASvhsEMvzjYnE
cFBcntDe7J6ZhVQXqkxZ/WNXzUOVoNzIkVUYOvIAHpnDHfJKph8fsRAKTUo0qMvs
7riyXmis1n8jn1ygtabdKTuDTGncjUzFsrw2pO6e8OfJq+ClrxCzjWYebVkhvKwW
gu1khvOyaY9WPBNsI1dItclSa+tVORf9gGEZIjsi4ub2fSbOHDuWFnk1dgNn8YYy
pS0JD90RQJOmpXBxGqG6J9OaNDrumatEHptsExN2tT28q0XHWJXh/86sX80QeFrS
muLr36Yj7SH+Q8Rx7uLFDNEze7V2rxglrENrGewSLR2bIYFGeZwsSiNhVbiqHHua
Jxrto6CbW8hJ1x4q8u9j8xCuIR0ylsM2K5uERj26xhIAW/9c4NcFyFTi+N78xk34
BZTCodkGdpAzn3/8Z3tEf9LtDrcBl4+dvXrKreqUr8ewyQTePX/b/5EdnDn4npVi
+d2/PICa372AJipSQB5/wP+WaVgBD/vuzsgYVly/37LlVpv9cGxDMfIN8CeYGVq1
/j/lnXv6+8VDtYn+1o8N0x77XmiyhfLUjDDmYl2dSqxjhcM3vrXwxXAPhW2S4wqi
9PIr9jbAb4igG+XVDan1Ighg/+dXtB4QUDpBTQYLE7OMLbRzdvVQWKjr5F1A61Jm
8F+tnJihBrETJIeW5O/lc7wLvG2cCWZPKz9UeU4NTwyiYLFFJfJDcPClZwEpmKGr
Na+azUaQ/vxzwdMm7O+nk96XdgeqeDhnYmH0rWU5oc1LYwAuUrXOosGNel8m0Nii
6AB5UHnsE75r+JUhtDiOU05fgdtuQfTbGCypUFlIuOgnWcBR/CTtOclLARadvxHh
IXh5mpZqn62t7CGZ/2ukII2NkNYfglQFRVRYry1wdmL4L/YI20uqeex7GXegg0tm
GUYqABzv1AnlO6NKppKLEYub1iSI+6qsD2fMM7hnqYzQ0FIIOCrHXqFdEXtOVC9d
lGGlDaFFbYA7P/iCwusY0XUV9Y2ZGjxp6WbqKmH53BB8SeWu01rabhJAYjNrbIu5
ZDpOx8pNGEvaVRRGatLKyaGlTC0CH3TgTIWjMsFICaRxz7kt2tyr6fi41kDwMTd5
CIcv2r++o04VpjeY5hmkf8c8kAcqfWGSHeCUKVeuP/LGw1ocClZ4Wz8wAE/e2N05
MUIiztUDz2UMJUkYWQVPCvTXmPBODBvsxR/EXfg7+nIYYhSz7LV3d5LRMGPq0L7R
MPmfM5f8FXf7KcGEy79NDnr9xhVT7/0F8lRpH0DuA8peHYItIFKqBLN1SJfMtOoH
MFP6r7PvIckzl3JBRx8mGUYavchn6zBwvuklldhHr7XgzPGiauAdSx1uExMhxK4m
AOwDc9YnsNvIplKcKRGpAdredsUUfweU+f/KjtkBDwgediqbLCL+Urmgkg7Kk3h8
bJ7Mr0h0j4cpjfNe3VU73eXYp2sOmBjDwcwlNf+HArGZjJlkYbVMLCZBpE8S/36P
SXZX2+eL4s7Aoe+h3ZTcnk0XlEVFP1u8ro+ha69zzYQQhXWVetV3uxeGfwVeNGZ5
+uOj9rEWa1Kq9NwyWaPWULusIoP8dqxWTHgpzsUrM73xp5mlbYhfmFHW8UZwPL+j
oGjSV5LUel4qYoCpcThyxTN7OOOYfz+RKL9x2Dkgtfdyk9o4flzFr0lGDcx7b9Pk
Vqc1BZ9+vL221RrNq3PoZsswZuagz2MVHUqMC29hCugV52l15V0hwjSsZVwk5p/l
yL3fNw4d684QlQpsEpVgsy5KwzSiZY9OmZ9sp//K4onx1kFMICu59ujn6Le5fpdI
y0hF6iSrnLW9dlWsOwhPVyfwYZAK7sCUOJlsjIl224ctN+TwfNBFjamGEMlSE7w8
7hyFMAo8VcUGyC1J0KXTLTubn8yr/0L9Q7nLlE+XPzSmcH5OMKAQtVuMHNCoZqm4
6PO2XkjPWZmBwBhaYHHwMn5ekrpiaIAMoFQ0hYXhqfM/zjwQ8HrDfJpWj8zmTZG3
NJK0JaycEX2QYWQSpTSizX5Y0p8zxRLKxGWZhpL9ci9telviO8LgZM7VehUZnbpu
gE1y4A+ptwIXybgj1ecYtiHxznidcpQmbJKPsygE4shSxr6AmVS5rxALC4KsALoa
GxrNBuoMxp5RCB80nunLZmJVw3EJeuv2PdN8xGgLHJzUGBU4xQeWGpUS/0jwHSq9
2M2bvOlQ2ZFUru/oBj/cEphjzpI/iIamHD5LOAfAfBVVD8vkiRN2kycbRquHrq9U
pDsA7X3d4Z72A6yAwqUhhHtNc5WWPIbaoABQYt2b4ghh2hMlMf25da1x8+f+HpFX
U3cEns/oQWCjhT7Eef+SdFdm6Wb37/E9blOUzRJYap0+HU7B8+e8vabxldPwwShI
SbFE4JAnFtVnUtMMf1vACLP1mEsDRmXox0Uv7C4SZUIV/BfhVlhmve0L8DKxtU1/
Y1g8I+jt4pI+Z6tEwefiJzKKlb93SNMYt/ndhKGRfcEissLH6scDDyM47VvN1EO7
LgHW5uD9/Wrwqjj01Qlz5r25SiePKHYfWD/b4jTDviMtSS/wb9TpBFeoaTXDnCod
fhJRDK8w052HH1kxh1hyN+JQyAg3avJqoc13oxQG91WK9e4ZO+vAO3u+IQpZWjl/
smkWBBf9c2gizfQvVxNXnlCho+7tGw9qMtDPgXVLGhIyXte42Z/8m1o604EKKb0z
YmRoiaLdkN2yRRdV/yLP++p3eDhA+mnIj+jswRy167T0ZaeO3mEgKob8FawAQ9S8
aVUxmsNozAw5noWM3Go2YhxbLFzbdLNA9fHYgff8knwcJIEID6astHDBA0UJ/Xlq
pp9SEfHHPN9J+SfpC2Es346/vMikjuA4OqUiFp9UsI+hNhMynrKYoN4sICydUIth
67K9sw9nJiz7MYcVbxDxAFnUptkBshtzpGG5rvnpfF5GHd4m41EWZ0uBB0iKRYHu
2CTx2m/lbU3HVTYsRA1+aAQwU1eaX2cBcTOOYTksUBmKuCp7Gsv4uKDRNgMVXGXt
48oXKv8lG2uBPYjmkNrnwr6OBb0U7uDaq4/YddkgmOHoJL8J4prUrJU7ONJzD02J
mvp6ac6ukYxDJYutRkqvJI9htBaf13MCoXU3b5iSI0Dio3fGF5zFxkaTT0jKXN0n
sF6Kz93ihh1/zLi8cZXzZjWbXC9IzjReAUv7D45qcIlbvogNu29VrMriTdVVhgKe
STZ7RfakYSRizAyj2p16rl4lPQR7MhGVrp2zZZuxePLXCkhtiYgJbUYAMWbf2COv
wg1S36yPWo06zpUfVZ6aFpxxFDp34uz61A/Vy4BSStjwcr8hU3wzMMZOhbf9k4ph
cdhT5B08ishWRVs3GXs9V4qvdWBewwbonm3mLd6TLUUegQXDfO5lwO/vBDCVdgIG
5zC4J2XPEA5zhl5Iw1iE/w==
`pragma protect end_protected
