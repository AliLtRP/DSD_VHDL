// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
uAyaCTdcdJlV+04SBIcI60jCBDnbEF7mbI0TfpE36UMoyXZRCdnfnt5V3HW7DIQIY8XxHxcTAMeQ
1d/aTt9CQf2QczecXfja97uWuxx/S1yyYNNP7LbHWwNC7XVxUAslid5J+deojtYZJFtQtkhF/vOj
Q58dQ1Lzs2hIMPK58t1hxdNvcq1IsD+ViwrwH/rtlblv2aDWvKEy4M2ht2vYsMfJjk4cpQJLFZ6K
Wz4B0q2ZIp9U8E4kS5gkABDBa8+xDZL+8uQI30tXMNs8yBoKtQfiasaFw4OFEjbA0qruAYcIgjZa
HYfmEtXHAmcYpFGw2YKY0+r4SwdQ9Lrb/mzI3A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
qinO00+AipXM2wO5EOYk38YWqfjYxmnYxBJgdbcXOJe7cI8CGgpdmULXMmlBNV5mLX7XpMrlHENz
Ib1ne89hWPldLVKGivN/Hf8KkePTG1g9r1Wq3h6v3oXVfyUE/ncmVatwr8h2ZioJE2cXFSA3ExfA
SNcGMMmNVe+mH16hpn6rQld0MdTTAs2VopWzhggjM3I6sB3FKp3XOiBNVtOFM6qigBZu8OssZlVY
AKbFlBD/7teh7oqtcqQ/PR+G3ApaPgZQ80kFQ5bz3DlUsQdYc4e7fEabA4H6Uw9aAokumb4NjcAD
pi2W67kn8tXIMv8+Sl35WZPz+CjdTZKcEtOyOj5IFSvUzze2Hgm4JfP/fUbuUZe7BBKNezDygkU5
5Toh2BVuC0dJFpQkvjhfPBa3zro+j9nY2wgryK+xNazwO6PgxTmWpTAJM+TTvKRfi477BhghocY6
YEf1OY+X2CwizLGEKUt+DqBZgmqvHmuG017wE+1ig7pK61KpXb5d6AZ1Kd1I7XYCGyRmW3OHnRp3
l54kA3naOFIpYtfqLwlMLnA1xa0P+7ZhGqfsm/2ZGMQqVsG5frtr8QaHqWXJAHarS3YwRwI1yVaK
m2mZtrrjjKuKSR9xjbVFCP4dcnRK5LyTR3kNGON+4un4FKwRWOqeaXKSn9EzhcY1fmiSAW1Kq3An
jOeXvRBtw/6XP7wnyvMK59WKyeDTTJb+fo/EVbrIitQnv8BrwvWgYlftFeT8NsiZoKo1c/OgVSuX
RoP5KsW8jtZNQLxfMIOp+A4iH386PuBxmTvPCoYqdiqr0rHK7tpRaEwu8hUTBWt55SwRFUvOkGmR
GTv5aknAMb7jmIegNeJGoPs5mg9fj2JDJbexzjpJ7A5Rw0YR1bpD1Qa0wLo1eTZZiaGhbEh65miM
h7NR7TE/YGiSaKaiNSKikmtF26o164WeDIqBODxLEFEF0rhL0ZDwwDVUAWIsQuo1so4A5cSiRaCe
YrtzUzxreFi0mw3kBmnG2mmq345YEcBuIoL/kUXLVU8ZfDezpzfiPpVfD0bbuiTB0ySFWc4V/Z0s
RVlKsyQZ1bzEHSZWwq40qRrJmfZ9A+AOCPcoUFgQc6114Mp5UiAW4uCkMCOi8vkbBi/w4i+XeImO
TeAbWZ+AYsyT2sHnWY8rgWkfXkGswB73qwxrP0BMGu7z72NfIGOHUGVuU7ns15HECkttLtNmwrPh
NJd6xSOKGKwiEPjbNR5K03uWRFmQR7pxfcjMJLMTcisU7pfZ8UsvgserwD5ccT38JRuG9VvJGkH7
eAekoCoV13PXHUNangoDRS/Xagwbj6CohzqD+HaBUNr/pGU+m9WYe3i9ToJTz6Zj3GtSg7FlLQci
t2yHdJIAMyozitZStOwxaRFF3AwrAIyAlndJLPp46AGLg8+6eXGmHMbFDFqNiipl9tOdEiRudZZO
etGVjLr3Kti2JzXjcE9gzW2Tep10i6dUpj8RhQWlhRuEmGeuMPo5FqCVa0RALsy2XkHw7yEnZTaN
y/fe+ynQ/bS1O1xgjDvm0cjNLa0e1ClFSOHuEzvtg0WlNZG1gd/yU7E2h9AcUCtU4YTZmr//DD74
cF+c0bDKa//EanlxuvpcjXrNKvT/MDqBepNtLECxIcceu5lfYK0kx4/+Rb2/bIwMRP2MAQPUdAzo
TWO+iksyl5Ho/wrn3nUZqgDpCrub8/kzMNI8I7lfdTmSEjoLLbc0HgdLgi/Mx1M74IJ+z923vCUs
C3GHszGFRLvRD90Ob+bmTuregd6dHf4FTpV54lnEKaQIScMDIChVO4lw7ThiVz8te+VR6K/3fur8
oRQ4yKRyHyTgBf4v8YbiNkTWMvvB1/H4x7IuY11kCFVEvkcmysX8T1j285kSMpPwUbYPlRknSZNd
BGnzh3nsPUSLQx3dt4ja9d5/M2syr6InYK9s/sKP+BxJJ6HjBs+thWMXDWi78Ixo7pk1Iq82wfuu
VulzoWx0QJkYkj6RrkydVBhE1rSbIwoF7hZ+6jDyRBm2HIkXM20fQacLs6xpGmH9raDCeAS5Sw0Y
aszoDWJpHh+wEX8k99/VijkeUgYxJaz3axkHMAIHN+F5XCuNoRSS3t3oo+hGeQJ9TUsX/JfAepKO
GAfiL0LEZtJZXii+k1AZhm0v6bnD5lnKUZl7P9s3WpFA+jVvJQU6KsYh2uER37JS9fC8MomIVX3e
uo/okJM1TekgkWHEAgc94ctH/aSrDVbDL7qFAlwg3s48oLs5L1FXAgM7fXxx1U95gJMHRoFnv4Mw
BF0YvWyxYiyN8BGW03J46SDcZ4gdj0zYDRe7DCHggkLNLYtU1mIQdzweH8DZHjQDJd8/2jM5ipU7
u6qU73x6KpUbn0BxpgYVqrEwHXURnROR8LY//ShitnGOVzsGXCNBrnkrL13b/0QPZSASgyZocgje
AQW20tAWKyxLn3afvaFamvf8l0Md0ZW+ujnCsbBE7CygR90ULrQszWcgpUBOptC9hhHFyh5inyYe
Ra6/SjXvFO7lt86ZdmEswYhaLx1wAgZSF5Lmbb/aZnwIOicjwHzVPT6p+I3sMCRykUpzES/2l4Kv
iLZjlAUBULFs4Q7u8qm/2lXZ3PuPhWsUIBW9CLWPrhsXnpZ5P3mDGVUbyQ2XGc4zCopWOI95Dt3P
WO5Jy03Qpzmq6CtKB1mtLEHyeQa9I8H507FmlgT8JQ9N+etCZ0AVBAtwpvlESpxuD1mQodqj7c5v
xmrFnKLqNuPzUa/CBMG1bX9JnTYuYa1UHdf344548k3dluWLyHITMNi8Do6i8kB+DuuCBGBs0AEc
DBVALWPwLq4ZogwFNZSTVnB1Qc+CV8S1tcm+7MZeNf/4RGWDGuKTGgl1GO4aHUKJD71v6dJBTk0q
Uq7E6wW2+lBSJjY7yrOI/pvc/mXdatv8mBskFRTsKC41UKead0U8/kapaoZ2DP61aEpcOGU2xO40
mzcQFp9pOCCnyFiQqKf4oTvvTa245HlGWO9Ytz9VJFj4J0GWxtGDtgfjrJsRcShc/peS/l601V4o
RVJaWOHbnKA3H7QnnDVkuTsF5qYG0Ra2jKUXSSirKEAjdPj8dDJpdLNzIN/56+c6GZbC219owfBo
DXLsPUbp0UgRbgnK0JL4+dlnrtQ4q1exGtnflFCiQ8tbVSbnYsYjamE4OS00FrLVCdL6f9W/5eOP
AYXqyFP+Ny0Sz8KMG+lN7jVHDoZHj96bCAqDs+kjjwo17OIvk0RdjZF7ETzBvkKbZT6f5zHWD3Gx
d2YgbNIFAb70egzI2taqKujgBc1R7U7xbLVjXaVcos07XFFFuyR6wHSy0F5w8cUsbGitBvy0oRke
jMFFD0VZmdVjkalNv21kotwVr2n9RinsEyLYk9YWKAe5YHVhv8pJPFBOTXPquANVUBiRgWpCAbTD
R0HN9AzMDTrfxG3J2qe1NiIaJNhD15CTNuBakQ0N0rxNha3/Dky+J7b86d6E/nM2BXQCtPbYigu9
WekzJgG3nlBSQf+u7w/dIJjakn+JoZglEV4cPEevafiOb69doKlpgGrIRd6p3chqlYH2owJTAcA+
VOR35ZSwUPdaBkh0YHsoOyPl3+Wdy2kY5m0Na16bUsOUgsgpNiy/vRWMJ1UNAD93JKcwTxwo6Y6a
ciThceNFL1EY2nFZaIen4Bct4ABRBgE/yBCPSJLAKiXF3s+ZePe5pxjSnEDkiZ65vxdqbsYUKaaB
OuoSC19OyhUWM2Lo/PnX81ZAHPI5CMmK+p9aBfMfuLRB0jC6khOZvJgGJokxj5NvVVjoJ7SQJJ6p
PuLI9Q+mz3m5RViUrOvy90JTvqJTXrCZFJYiFcCxKuEljLaq7DP6MdFgm8l4DL+VH5sBWEVqy+92
Djn6z+royPpG8Zab0sUhdLfyhNcJ67F/GQs5JuVgspdzv4DiortPk2BKDr3JkEWsq7mnESGLC3+i
qkDND51d3NNrJvXrCKYcFQ2fq6tjeEoKkKIVYQLftnbOqtKi3hakkb7MbOMucwcLSmTNfyPkt7nx
nNP1QUuxCsbFFV91c4GBM0AfysQFCp9agRQOS95IAjSLBwrzi8Ay3pI3trmkShJFxLiNe8a/WdrO
4yVT8H+tTolKuu+86qDPoHQLBHPktI9uC+jn+/VbN+Z947an7SjQnKjo3ogB1+ArOwyveOxnNH3K
ECdgR8ARJ4O20Bi2am3JDWkq550wqzqXaCo4/lQSWXZvnqqosF7IhPyfkAs+DMD9I50EF+Nwbg1w
dXp2NxA6PLBijtHa+YtgJzh+/c8fpNBgB2wjGHy07uT73qrF4yhJ1YeFe8Ydh5h3avnpnP71H7io
ZnQIFyZ1TvuK78mAzFsq/Yt/pPBrRFH8a2SMFZESPkaRUh8TgSz76e7TKNXSmd2NnGNQH/DHBfNp
EDB7JNa6UJYGeQiUB5FVkE71St9ONQvZHk075Q1NL2Pm1hmQoqlXkvLdTIQPTNFR/rk0TUd/2YSn
87CFoiVFaOrHOhZc5UH1VP+GA3IqBOYBV22cj43Ffuijx6gbBr8YjlVR830kITRU/y/Wdsm582XP
oTi9kS0xz16P4ecI9Ej4gpdW9TVi49vckPpq5Ts5Z3nZdoiLsPCfscU0L2tPZvDfv33nwzg+p0I+
cvDu4fYhljn5rRoa73fxre1G3Rxrw4/PXX1TwgMII1rVnIYOFRoqRlTNpv1P/UAoAgkIUg9MDNmS
1psuhRLGWOtQjeaaeyiynR7BjkGBhy+WMsl6cNpUyAjftR6s50RMVaVWlG8cMrh22PWCMF/Jz7Vt
Zo39zeqRW2U1gajchV/RS/FE/DRn6F2/9BRzCmzToiJ/JKXAmwrTi+E7lsCXSFF7NHXrt9JpZoBz
7TUBupl09fyaR1OaWTdX1SCIwvqx82wdt/m0dUNWTUqzCnjSBrZDQAX1eKpSyba50jYLKS2b3eY0
QRwF2s2Q1b5AAlUX/sCLXeKwtVaOfQX15rMuqlwYj1z4prfkYdp51xGxfwlsus4hFPGYFpBb7BE6
yUFyz013s56W7IvfvyT0vcylCwAmhoVpJ5qkX8IvJueKlf7FbFN48hqCveRXNTKRgJz7a6KZxd4G
210EORWv7I2SsbWzPEiKAREJwaTeo+NHdtwSbQF/fGFmEdAAmTDAEA/HI0tFH8alzEqwUuJwHJOr
hW7a9yBeqJFIU7/X0XPv/cckYs2kxyPfBvEHa7jfqNflIgHVCmEcpj3h4Fvnft8JQDYhVLuQt9O4
ny5hbvtGgxNjMnqU5PylH6BrgmkbSzySKIwVKsLzOe2zczHQBhxHkskGNEGN75slRU2di6vJUpDX
L9S2D37DZwWKZfNNgc2TEATnrXVrjLjzpvq8y5YoHRy9Qg3pg9of/WzXTVTcy5oGWYjA/WVDgUYP
gf606H0RSnyILzYNUDPtM8p+LWMfauDqfIsIcikPjLW9u8T65W7fcNqXwtgWALs1LmCKiHD+gges
N8scnXRVI797ff2pMM7zSG0lnCku4bXZ9I8Uk7yqaliN/b1CbQNKbpboGWiPjgPNz4kT6t+XA8eL
ye9FXJJT+VCGM1I2mbBfT49cJlg8WUVTYQLGpqaxIOj+NrGLucEzKv4fREGQ7TnYHadFU998l31j
sJWc4Lzg5GWjoTgjJhhF3gPk6gQXGhqahO/nWs3DTL/HHt0s5dCcmN5rxlPoMxt49/uCCVBzWkBo
mMimFz9/f8qb5fHzqUqTs/NvJYbrZdj7Y2Db0uHvtRd40wrop6IWwO2spx3wRYrfCf74q2tBq9nU
CMPhu5HgtHfRFmYjBGTkPTCN/yh9GlXLfNijUpdQLiK6ytifvKvZ1Ey640WY4sbd4pIPUCWziERW
/8W/++Ly8OTbFuzzLz0/OhZVP2jIsDnz2OsZKFOUTXbaYdNBEybg1Dgaa/QDOxA7yckoIos/AXQa
HUjGIDmcC/Vgn3gpbxJ12uIWpC1mVncLnSioSAxvlh6mWAbtQfudSFgvhXGWRoq6WnDnSec/bU42
bwmAEGcmOB1lQ76uWF54Ntaows7JScy+vF+/Any9lBzA6mdOH0x8+0gFA8LxTWQmBcZEPY0hwfQ+
QZtnsQEbZPez3NHGhqvKBI+eVIPDz0vXOFQD8LVvlXkUqatZFJo/6cJHMaUufd/8Wqde4k8uX7gi
PvskITNkFwFpj7FpYw/P0MWpCMl+qllV7QEswmGycpS2IhsND4uWXz/QrAseJGbrVOOKYXD2wVy+
f6EpE004sF4w2gvW3ta+LnYA4knF1i+iCR0cpnDbDBiTJA2PX1wfAXfI+3GSDvDWV9MCrsEJC8Hk
1xyF1bvt21tIqvRjMlbXKNMhPefjQQhtg2a2iYc8nThRHJlOFYr1mAUJU9WW4tOR57X2H45FdBMb
l8R50gTdA2kd6plrBwnk8Ga6Ggozf8T30oJtME/1jLSP8sJHm4jfNabzou2ralleqfVrPvybzUKn
zeJg0ZdAdywr67+3W+Oar0iYnpNldTFCvD/kknd8Br4jzgux8htt4uACgetq1MmNTLCH6p5Wel1+
PTPkPq2awu8QfmKz6lIY29etY9fjuDoGy7mGeZpqVfoEo57XQ7BsxQjq857s90RrHTXy75JcJi89
C0hazc5wBUn4Fxw2KXvhkUEkT/YKzga59mndNC8BWgQYi937lUUIQOx2fNsnqOh8aNu0sPtH3982
54kX6UfK6GjQ7L3UR5bukXdYcB689hLBwbdLtArX1FjHw7NbQwTUloa0C4CHU3IkrWY3Nl+/y1/I
6BuTBTBdi5gXPH9W+DkXmrJr75cEgxLO+0psoKShZNgyGEjL23exKDbypnMdQVfkBJqEgPv0mimY
QnyLe+3w2JUjDxTiEpQKZeIVriT3asGJCPyHsPpGxOJ6vW7WmklJiVzNPQb8P6li7Z7nOMcN837q
Qz6I1C2UUSEsHkpr1UIIgaklpUUwwGFijwPDuWwzHmn/fNjraGAleY2Ovu/R2lsxo72+Ac1FQ/Tl
FLrAHvIT+emTNiC0TMeP252y0flbTWtX0ki00ZLWsEyYE83/wSd55gqdw/ps5mTmeeQ7B0Qj+33V
C2BzBTnqMJ/eUzOxcH6ILpL7R1VX5dNAGViCqzpkgoJm1jJQi22WHu1TMMKSFvxkGmRSDJsuaXIh
ClOUtfU8iHdinG+0T5IznxCrEhDlATMUH6so9cVT7GQUh4g1+ZW7NwCuyd99shDc0X4YTnfznsaU
kbR++U5GagZvof9r9QrTJWRB+CjdJtVGz8RNxU5u0KQw6rWjN6lWqK4BfpAcxiuXzBiPRGB+VXIM
u/1ZXWf4jNMbyb3GKgWwKzgDoQWNtrkIpKHDlrbNpUNxWcbSjF9WlmKZMuwPepdLVZe/WQuWnvH1
28Ipvou2CAVo8PrmkUYNx8++caBCjOcBnCrhAYeinkYJNPU9ppH6GptcX8qMbTaevd+l+9ZP34e/
xCEEAbPZz4v4l/erFOrVPMo5qGrOJdi9ktiWHtxd2zPtJYsBTRkS2QJtEiruDXPQJbmhsl0y7Yq+
yuzmmQ9c6O3ZhwtIQQytBQdjnsrt0686Rz7UEaN2Qt0tUban1DM+IAJvAv8W2b5qyGlsD2hTX9pl
cXQ1UMMtoM33lEIm4DdVwpB62fv3dw3NTV7F7mlEGE132BVDsyS9ftV5Wo4BKEHt+sUwS/SeSwP6
3cQB8Tpbq7y/KgzpLI5ggLRbmFP3my4b0q2AoYVUp5ZmWYSd+TOWDje8IUILvGZDnsnOw3KehCj/
HCMf27RcfaQyBfa25lp9ZBF/mGFq4BAWNqBIvXrlMRvIV0sKuBwemdWdUkLaOC/f5gMsTZ3TZ3Dn
O0SjeN91q+fHU+OKnJxh+l5Kh4GAlFNEBgaitqX3DHNwht6x12DsFQ1Eb49GLCXy20QaQqcs6j32
edfYF6Lff8OI01gLi73VNUXiXQXZmImV6pcC6im1Vxx95Q8qqxrr2M5MkyCDmXwZBocO3My0BO0R
fmEwjB7Ju90KyY50duif31NAxiyhIv+1G7pXU7lmzmsJLWS9eEsp2Xb6TchIzm18MZZprvRRnKmP
2HOkb6dz8GX7iOvdwYKv5uoScRT2enkbQEyqNL/NZubJ6mbbiB81/KOg0uP465msGMXbLKzJpab8
yNyHnahRD+3AP5BJ8kir9WzjzQj0sdsXkE0rUKRJYHcxtyj+QWV5Ae9x3TXIwdVGYi7RvNFP7uJ7
qlODjcVCyu1U5HZJBjx1/PCjeYq9IwN5rRkSbb0nUtKzxnoXqTwEbae7o7uKU/XyK8sGIlJwwpTb
qnByp+4tPz+/5/CGpEcG3DbBPaE2V2jz8Md4Hk5MqBDJRztVo+HapXOXVZzXrLgs6IkkUj4PNa44
dHz7Nj4C/MZlKuutympNuy+9v4E0hGn35mhDdXSPhuh0A9BLveDFH/bplSul0C+OKCNHD1JZvhfM
O0kYY1YV1OCOw6/H2jYhzTmEXRiquQa3lehVW9Ny5PTOmaQbRcNgN/YNqIlPAJmKlpwFgltmU4YM
c3mg49hyl7oZzSrwCEBtwaqnrKIi0gFYEDbZaU+K50whYLO6n0u0Gd+xCvGDtaldtnhZ+svkRyaE
bPZ1gQF0n5662kNdjhEIThS3KpUkTJH5dukAnoWz3WxwwXA9iVQmWZGFS13fcMjj/G37Rw0YUyqp
QWBmwb3m5c3Zs7fkL+byB2ieTSaiLwY/ICUv3zVNkcMOW9OOiTLQz6doQvZNL1YiS0My835cxYxF
cZAvf79D2CjDTb/hB37tCZGOxCnXaZKdBVmjLFlC8mCThw4v2m17Mx0gjajPZuZBu7+G7bSEclut
lWRnNgo4IDeEGE4Evcq1xGXoEFbEklzvRAnVnvjxkRI/Wr+RDlC/BfDA4zLQFW1bW9XEsIqD6op3
0XId0Oya3bgZOB3WFWlJc8kfduQOaGs+sa/unRRWlxXzYWvHcYMfiNBfb8D6cF5FfvUrNvJTXH4B
+VJbe/CeTEikdRJT1HHDE1gxa6cvutW4TJtybtscqzDzSknqyrf/AlYMMUKNx0GCROwF+y8hv2GH
nrR3/0VH0QF9CK5gS5mgis5vB7y+yEkB3QDFZyuuYPERz6rDf90dOIlzoComZV50rJcdyNbkbAc+
/GobYfMJSQtVH6/KOJO+jge6VQxQdJepNkX1rutbe6sxnDFRGTNpkeVf2j88CVl3Zj/coKWDsUSl
3VNoCnGnd0D6nKz5EuMHUReZXom9p59NLvJ8e31w5FIER4zlg7stYQAel/IVb5e2WVdeLBJKtjLZ
EQmwTviQn8ZcMfU6KLiMH1UfBhXsshXHAy8cpcH7/Y28xve8FEWQ37tYSP7L/lJgdT4066ZR4Lzj
LeANUN0zN4zXPbjg7PVB0x/0c89+/2CmfP8coiEpogvoT6Zjpc1Zrt6VBx0VOCPCS0pzqMVctrJS
n6t6rxPjgsnN64XdAtQtPfq2R1M2dwxLaogBQ1Y+uw7HQUGjvhzhGjkc2Dnagrse/TJ+Jw1o9JWp
VRufMkiolTOhR0BU1ZWoerDtlVifak6m1d0ZZRhTtlV+QoHNTUC5FcJl99dFJXRYf3jII6ch6V4U
9vmOUBGlumVjShwZD/IHdqp8fKRJvpmm6bHKgOUs4aZbyy8FMoZuYP3dP7PNeTqbr7pUZXlhAUfz
Y6JFpFBXPpaU7ICcE3acif3xVL7y6ejXMvQj3/1QE8wFzK3Q1AkxN7UB5U2Vdbbu84JLLNqasj2g
Vsum+pvkMW9d6DlygvLW2TAuq1dVI+Ymdc1PK4q0THdFAgQWM4UvrudB2pUAQayGNr1orDB5ORiW
Ox85kYwGB0f66NKBNXk3vVIkPMI6hfgfTwXCyOiaP2YIPsTkaEhfb+8+PcX5v8zzyVfCsK41jk3O
YRj/PjfH33owINJE84uoHJgdw6J/tDnILQy8aSXVZhY3RV5grIie0WV9gNlz+tK2vo3OXiAfH7En
jmagzNGdNkU93zdgZvx9GCLqulXED0TD5hQByU/d+9wqwkFRjRhWUh3ZtP6FhZLS1s024ZJ9L3sy
JKAvFC9mpryqJDY7yUFtUqjpQvKjK3rhC7xBmtkzofH7F7QzHzjZ8EONwkrl/JDIgnE0OAZxC03p
OfQuPX33bQ3V23mWN19cqdRd5wcQi5D/GgOUB93Ccvv3DHgFWJw7XhiZ/V8jow7x/oqD66nH8hrY
BVqopz/CpKIGzKiZDs+AwEqJi41AJJLMvOeVAzLoZVhJhkycnQndnUc5mc8mH9eG+q5PZTX+AQaZ
fsZmmoGFD/S6BMlOx8KPQ4KK2vDTRRD08uatJDcKvrU1lZictXX2uvJHPp8AiXHVLN124tFqJDoP
z7V56pO9+og5FNlmoNS88HjAB9+A+TFnDKzjI3NWI7ngPHugRCNPvN0MorJA14BVG3/RhF4/1i+S
TL97OACZTHQm6Ze+gmvCb544tkgU78ApYVrBI0BcAydtr2NWuqE3lsPr+Nxj4m2zy2sBmzhLHFwb
PfAdfO6tCadlG5Ksyc6SHdPyGdb/wRUfmrCBU9ghW4IPsxBABuszAILrbne/aOJaFNjLiRDDdbTi
0GBbGLnBUzcO5mIoztRTYIhZRNzYNAPrrdCfYV52JR2/zzVEeEl3fMw+k8Uivp83/9h/NBPTqC4t
dECxNOqsw/1k8FgLTU5lkK5CATyU43JsuWFb4fNJX+4fZUx5Xr8luVyQy3L20GTZxoQYVfvKVTdW
omKn3vEjQy6v/I9wT0pJlqxyDtbCHmMcuFvwjDg5VMfMZ81yPNLpoQxhA7BWWD7TFgzG+MHYrKEF
Kqmm/+4sZSMo6dUC/DiiD+MYiTRdRLw0QPyZ4C36Ck14Bs7nkpZfLi1dZo0+YFJFI3iT2vVj50Qt
Tvk/BWI2gQgxScyas+4fzJlw5tLuR2kpdd+ham41FUHd10rI1Ct5q41bSXOrM+puNLkt013pKuez
FVIlJ8hjx8BpeOjXHV05kBACh3xkgYklSDgt2CkKqFHqKmDgL/P2dK/esjRcTQOlrmhlHpOgVz/C
6EhBSS6OuqoTe6qDvi/RKPuhArkE3hH9pyQWv2tVDGXCZUYvm2wluy05djsDpvFgaGD+zSEgpy2/
cpIrz2sB1CDrIYDiLRAh/yLbPRKv7+4Q4cev/ucrIb6j/gQ8huqjvdLIfzSizrZVbPeFwL+DkOFj
yPx2XOQR7Z4o9yCU08p2zXWIAt8bQKXG3uOMy8Y3DArT2O8jBYjPy4kTtdzOUY5P1sxcnm3sLLPb
BLfqnaCU5HfaeCn61fqXywL9wEjQm/ktXOK+AKoFviuB+NtB737XytaxwFX+FUHX0xIXvy/P/kEY
FQ77ZMjXuW5tU32oRm2mW0qbnLEC0jACkyubG7kZlVKKN5DisIhQBXYGSPebmgH5P3fQlw65l1HD
w5PVqhoscxD6p+mNyR8xb3vK2Zw5K5IbVSbY3XgmqE/mcxwfImLHfVweIhGVDPiHfHb9fryvu9jl
ZzdIKW+qu3CHaZMfHPNlH7C+cJX5pEHzjTJFiiwkhrwnKuHp4m3RQa5vFnP+pDC3I7WQ8HUvjbGZ
uoremxFRYumnXIcxT1qqG5L7wQ0VVtAVc5auHFgMwXn+pWX6YnK5Gc3NY9EZo+ysc+1m0k5DlX3A
1D4Ttyo1fa9GAqQQ3jELGt03sDQscTA4zmnEejakL+mdze3ilERHh7pTSSKAxWmrEFyrQ+XYH5WY
jxvNkvacfK20Des94JHAlnp63SVd1JmL3jiJbmeAnLLKZi0JORRBLbyvrYGfq5syIq33wPQ1qKcq
i2Bdv4KSzpUldwqadN7fLTyi6dE1hnRldU/RFXVkEw8hzEI1MAkXU3bUEzADG/hD+bM9sTtMd8cA
Y2KN83Kx5QwQr1lLnCiTriXSQ2KUed2UzDqr+blQwDiokRXKoLDgahlNPpQvM3gZQI+tw6e2e3hY
ZnNk3HtLNrieaMJhSw6m43syNU0sy39CpJPCjubv7xE7c7A03JJOWP+VD/DgE/TIvmtJycaBFo12
tHQ6eV0eSu26/RPX9zJUbHpnKj2hSKDY0EveDQJz1AVxEt9K2N3mnhrj3FPFeHIq8EFhp1HBqsTO
QL+6ynbtogWtv+z6H77rIH8/B/kkmAFj2oSZLNqSBkrS5P8T74fFTGeD+BhLGWeqv2JWMhDhFKgW
vHygga94fw7Lim651nPwM67uBK2eNVsKeNYBeO8euhZIxFbRt0mptOp4w6zi9ejTNvPO3MOsPYpt
r64ikAYdjty55+WToLXuv11wA3DGClR2UsLKhKUqg1+vLRPlbxD5ikfXmvEGP0ylNqQ+dP6gVPm5
Y2J5wVs9zm18wZNgMrVifjqnti0UyIKZ1NAiB8pBkm8/8I79tbarwE3C+kA7qFmVpfm6tKJTnLS/
UGXbmedGYU86bnYsNNE+YpdQc76uSRr43Cwn/gz3MHZkvFgXt7pyYZQ6sUY4DWuXXZCLTHqpz54g
tqQm/E+HBm8y1qZPer0P3r3kRzCT5zIkxCzKzLqHkWYMP4JPZ+LOZQ8WWbjsJyBFxKGHO/15QNMS
0MpdIWT4VMZgeoP9V7w6zHKLEw8C/0NCiEuln930iWVxNnz4nDfTjtnGSkXCkLxW5hlkKJ7qrB4d
oC+CyjW36vYU85k7+3RsvUwz7EcqzjgJ2Y5tBgVM4aJvJuP+0TPJFe9kDlx3n3qoSPddbgSeMZHS
GX0812bYOM9mf73RAnx2hLddyRKl5tT7gZdxTpGAlxmSPRT5/pcUA/mdCewdhiHQwJdSStdpWEnq
e1/TqJBtc6wQseAU94TQvs5iZSKbMcZ0F8FRF3LdmyZvu+d0sa3y8pKlmiAvpHXjHgerumBm6HaQ
9jUEj9zoK/YaqN9gQbkiaeviAxkyzLC3N5Vgd9/4xD+PNb6RiDpNZ+yyHfid2cOaXMOlK9DcUlg7
YXF4iQQDIZTErh9oZy9WML+mtZM4X/xWy64od4wESOhLbyV7ZD5/ytsl4pv9JHwCKn5w7U8XMQi4
DQj4G2zu3su1BMC3GC+aW2jamgQf/v+pw4ugahWFCVKs+DOp28iVSvd25JfeNCwfTJ6qcamQSsbK
cvbmqiuLCHX2fKNVM9m/zBw3rZqWjD68Iv1gOwhIWJZArVFHdyft58LidDOeItkYoK0g/HGO2ukQ
UrQfhOmsztNQ4VA+nkQJVt+ob+LPNABkQk0znLoRtmOkruFIYfYGJMNes1cAgJ4wM1CqnHQr5/LN
vET0vA4n+hv6Bi/qmnwR5mrUOZkkKNMNMmTu/2QelS8+wMOMr6c5aEYxXbpyBh7A0PynYUTGGh0a
U9UEm4hveqzmMHS9SRF/FEZHDmtepCNs7oa8yfsHkGFlSJFm6NKarVjAIDul3+G21MEUq4+DMFvl
016i3dV40BQiwH/CLc7jW4CTJzsSm2LvFRUEs+WyET0RuPEKCmmyAi2Qanbt/CrFTT+wUGpIk+GP
dGI5cHAikm7JEOa+U7FnUEUjqXdMvlONFinv0sv/Q/pqSoqEl2zdwdIb9T6zuw6VdPR1DB6IgQYq
9hmwalGWud6OwCd0nGAC5A6YidUa/DVXvHW6bz710Efx+JSmml4TqjfsVSVZ8XdDphGCAvLdfLO/
1XhyAG/eXtBgUmDcxyyKomeys3jFGYJaetox8psH9usueU9HvEEVc1g3odsTnrKIcvVRe/cGEVUG
Fi80Lm66GipHiQ/lT5sQkNYrbjN0mIGIBdMjvi14UaeXYFOKeeB4sPpQgKUQSelKOMe9yvMgebFp
mClqTVaNqR4yAK7euUdaoFKivxR7wmoJ2ATji6jeqglxHbznW7CkcgJeN8P8otVSJuXavQ44YlDr
ju7J5heFu3m4p73n8BIRg4QtlawSxGsWRtyKtQDJ1fFChYPAwgtOepuonUtMl85XKVRNymkV+Uix
YUb/NBjLesRad4IaWwMdUtHpcdhJqrE93pFLylTV9HK4SvGxR5xdsr+GtE1q+Kwz4k5XGL2oGUhV
FD/x5OIiaQyJ1YRQDuG8nvtpFC5uX14ZtixeqPgSE4mOSH6JRFPbtZYTbhhn8xze991pckospEJu
/kq4jqj+fRfB+mpKUBBxDkmWo3z/kbEnQ5hLnoXvvyg5wAmk/8oJgqo9cfcu9IT4m3d2Dv14QOeM
kCiIL6/JypSzpPUTkeY3WeoNyE9rGbdgvGaHjXA0pX9updq5Dji49f19LBub+RJ7XeWc2nDmHoRe
qGg2aHwGH9hcVO4rD8JVGw2OJkavo5HcPkdyWq1aCWy4ymjkjLS+PDKU6+XvJN7ePI3jvV4fBkow
RzQ+0irjK9FWCeKe8S9GyPPAks0co5rXGOOzrXfikmXmBSHNuX6beHH/IppYDrlJo5cTSeO/Wn7x
minUVIGVokQ/M5NAeQFDCz5CG4Q0a5VaPyXfp1Ny3DbEERptsJVb+icxniIFxx3NcSO0BGNgZe9o
/upT5Hs0MmgC68ImLpA7bc1oN9YgoMzkzwF0aJhIYdIv/4fOhZ3xTgyR75QuzKNiv4daFxFG53Mp
mckIciSnlcx133HLGA4DpdB0KF6UP5+V7HVmd2iQOcBACj1Z+D/cAhOHUqeuddZgQ/2yQHqlrN+o
NiGPYEtJRnWewHyZwgms39EU4WmTEAHcwC5CltQZbznSMtAo7m5OcQj3xpJBRUBMnYUF0Kwwgpa/
RXepvXZOxdAGWZkMiOABAX5d7dcOb6qaxYZGQqy12NOTu14we6MHdz+OY/ROVSS+025Ho/nlCRc1
nfqNdlFOIrQvOaipiNhArEh8BCOnaedB4iGWXDO9VAtYZ2yH9wRMjtkYECGF6r8PrGHZjjwBW57s
wKyyboDMVWofM3pSJ8PLO4kMmjq7C/Wj4/pr7CUa+5Lh7JHbQkh3F4yNNZ2jEPDJy6zpJCjvXi8O
K096JfHgGwbxy48qRjxyvVDf9gZa/NCA+0p7FCHBWMR6hHIfePS/sb9ZqZJSbw1+50FHOoEcAg9c
60pPGJX0mL4s+cSe9AkEz6N47ktxEhl0EtjwAcnzt/7QxjwWq1P+dAp3dzztslh6wofD+YqlL0xd
j8vgjM9A2HqFw/KJAmToKddmf2Q4t/3oP/wHNYToDzY5R4t+tYGlK8dis+h0y9jUl0KA4ff4/9EO
wgQjZsmNy1YDhG6mVboeK0HJE2efMytpqwtyMWxCpibElzif7T10JP50HEJ7UJkMgvFdZx63y4NR
TB8cCkaXVKCK9BKShYj7nQiPBD81lyMOG9uB1Min4o+4MV/OmPHHKB77wKGEZGgFBF1/E1zidGdn
ExZCVrxh4c7hjDVYzAklFmf2EIPrnesTD/k9995MPg51gd+ANTl1MK+C47GxqZSx4e3mPCeHOOi0
cW8E/524pBT/9uzPKRMF1Xhh6B9jEYagt8wB/hZfjXZWQ1lp6SYhfHTkCx812D7Icn6j7odHzRC8
xlQD8wUVHRB7BU+mOqFOFq45hvu04c7lBYN7bb9uKFtsk65mf3jrdEVlB3wA5GOlAnWW2BckuQTC
OgoE6lM+sY1xpahJxRNBa053+bHZqHpEqNbLBTSpyKYHxv4Y1d7Dm3+cs9M7y9wZ6LqM/xhWFgJS
LpcpMnR6C/NFcqzTCqZ80AnsNUXV19E16XIsmReT3J6rDcWFPX7Z+BeZNATuiArjlTZWsup2iWlG
rAAotsn93MPYRo3QpX5nUHLgtadOmKJZPDIcC+eD4gVbsl6Yc4dYjzWnUQ4eYZi5kT71EevbbkwO
dr08LFkUMBbgC2VUaizHYR/9ByHMogm/viUrW2MxxL1Dx4gD4+vZGxHKOlSs0jho0NlHSLrVUClA
csHK1vUHf4NBEmMW4WQ5vrUOnd9Qh+DHiFQpxlZ8tIp1pbp2l0rraWApEmDusJ2iJVkKlncMsKi6
DEkmgSE9SI3WqPe8TNfIGS+jHNXyfTDM2dTpM9IS6j4h8OvN8SLtZn0xvgldB0zi8595OSkjzsnn
WRT9iJdyKhFDpPkkxQ3FVt8ub9SMQKT95eg21rXFkFo7EsHgAI7bXTanZmy81tQbS0e3HomJ6jA0
sDhCY8z72mlMyot/lZAEfZHaOStu0/GZprm6c8bF424MtyPSGC6kC+ENfDsXcYcf34sDuTLXSN8i
PXR9ObHqaKazBoyguy3RFMbtxaEIobCC/oZCrxOALAqcwy/rbKuecPvuFMLoJKMnZlzEr7oVmfFr
23j0YWJ8OfhTKoVmeATGdwHLMZo+Rn9V/IbY2RbCDAy7UGkfXKczB376himHFuiMToczFE5Vu01m
wqoOwpjimbQwZ/ELlXn2JDAsw6QZMrxbWGzW15A4HQfHlo++GOvG4gNuQ6KiPhhsutAOUI22EMsZ
7T22q+CtQokVLaQDmxdWaHZEwitL4xDM9V7zC0KXk1/pHKyy8UQuSko7H0zgT9iYhXvVwPAz18/E
TaBx0/l6o+g/aZHAM9sftGiQ+ocEQJbCPBrwcpGMl4/IOCRGFmaVCpgm44jQRluecGmpQq12Lc5p
WvL9HJ2sWxOKyIyNiNns/NjbfXS73bqkrji+01qaQlU+CvJWhY/6iPnMFinXqjge7jJ+T+bs3jdB
k3KmOvX3w6OlHpj4zhsBoP91pmmIy97d/3OglYACswR1Xa37QWafF/mZ9mBSEfkfDInfd8nzSmRk
lU26DS/UEzSp4bJYau4inRmWVs2FOsv+qq2kpku7QIUljrWgoQLHjyH9K/616S7VcAqZ+0yb3c6/
sWC2sBQzRxVGurNXNsDpWbIfyxDtmkgaLIk36xhZGgeMgrOBczxiIAWpC5asMGc6VOGmkdUqNAUj
MtNg6LzyDyhXpcf0k1bh1foeLSxzK2WEF9KWllUcBKt0Kxnhu6zKm2BirH25Ki6sknTcVZttIsJK
HvhlILLwCaS8/x7ZHHQf4Gi0UG0oHeZ9wxj2oU+WQ6LqQ4H1lr0AUsFcqurC4XGSiOp/th5Qgx9a
R1GT6T5QcpP82M4cRZU9KOP+7rdF46QXJe30EVH6pQAnbMGDwDlNTvE4BaJ6Fj4HrpFA1COO92Ov
i+u/8z6PxekuDALeECA9S2Zd29kj4L6NMTqcnX6SWOBDCBeuo6YVVeP6QnufwD4fzcqPU8xqfjar
EENocN32+fEvsbOHyDT7yZd33SvCG8uSL/75XD3D+nzsk1UdtkF3UsBUIXFVUKkJpp2EP22iht7v
cx3vi1/vmjqZuCJOEhrObAEc6BzJ4kYufsnvZOgh2Axc9JhVAh7lfJmbfAsiFWhsl85QCYhmwfbh
aHMSkWK0o3rXbX3MDpsfyx7vXmj8zQYreTZG49RlStIjLUcSPbxt+bJepuYAosgY6EAmNNu7NaTg
UeiqVCCCxMe7wfL/iAbZsGniK2CTgOlF6kjsMtvmNbhwJHMxRWdfHPgBbeWvQsfiZ9TkU224/7fg
pM3sVdtJOjGSHmKpTdGDQs5Aon4wvLp6QLQ4NwlNnAl9/0Be+C+sytxp5ymoLNe0tyhLzsHuXbdC
kksuC55IC6a+QHnnxelCtrMDBjYjEZNZWsEN0ornNMc4QgrgoodKl5Q8oGoguqLp/YMd3QvNr6wf
VYNvyiPIAgKebVhp0Raqi5PbxcNkg3ArfkuvKvPwNa4XRxzxv8gT5hJgg2DN/SkSvB8q2222P2Gq
nD4LRBuNXLejqVpF5uNmXdbD/CxxnzeTt0eUBvDBfLCHMENEy3VdxDGjAUw6r71zHQrlx+5BTs/2
N4Rrlva6InnEdYgZgUDMk+81UvCgj9gljmFGkF4ykAJsX5RUDl3jpVPmUWJoOuYUsm/4b/hwDb/P
eFtWQoMBpiSP0vi2VzjIhqTNWeURi8Km6KYAszeCkUbqe6fg7clikxQ8fkad2gMjsWBDgftgr6Vl
ZNY/6dB/cf2AcggU0DyWEHlmMSl0Y4ZAk7yNIiUUC4do/RNARLs6E12ih24k6G1Jd5d+QezP6wwY
wd9rThPLYcu+5wv+Iw6kXhAPGP+2dro7NvHsOCaW2+Nqfo80b1Z48uCyGeWYEwyUmn4bZg/el7wg
32wATBfD9jOLYvXJTd+V0V2EVyOzzvHCPtlQ+pqwfcMnb/CRpilsGewUUWQbgsBweLrRJ2KJa/Jf
jOvjR+fc4KqxQo3n9lvwvNukynLG15Jy+SbZIM7G/GZ3QIHD4asr0G0SDpMKbSu6gRgzXTRv8zZe
eiuWhVr6tzSzC6OVLYelY3wJ8Ti4sbtTtHQun6U6Ch6jwVcFM0prsDIp8bw7L9lJZ8k9a6y6cWjb
GPzNenOfIeG65pKfrd1ZgQQKchigxGCDOR6DVl0torUQ70YphnJNY7loQpqwED8fy10vd5lV/ksc
MkJea8JzyxDSd0kwJaOviDfEXqlpBnoj8B+u95rTd80qlrS83PWbSAQQ0JdIut771YmGbei+rXBD
aWv7362hCUSDrwIma/EBwye3ubAC9476RlPhtYD1+oyI8xG47ZeQ5Vcs+Xu+uiV2F/LNz3YrlFfO
AkBNrzX3nl18gxb+rqzXnfS7bQAcJ4JXyhghdcReH8440Svjao3bYX/ZdxpDtO2XRQnBZ645oaoH
LwzZnqau70vVUYIEaBcj0m8XQmKqAu3oqFd5nF/F9Y9UY17pbnf7v9vkPr/IMpLycvSLrOAlCIuy
XkUAvS9DlZ5J6rk8gBdUs0ZPi3AGihfrweyYXJm/Kvuvr4eItCso3IQ75Mu6B6+Q0IIYob8ERR4J
8Vca4Mk6bnrYklqweRhy0uhD9uKRbHECamITe/ecUoldGE2yrvq84zAGhH8p211Hl9cNqd2Ub/YO
BFyzrqVhPeIqx8fgccF0JKgGsbD5mdaxW9mACbcAVSxLybdEUZHJOcNdRPp2TNxxDeOGYimD6b+w
HIedKvdHwgMyN5HDZvlPzcHeVqGAamozeRx8HIayOv9wKeUKSIQIKTChEaayyqUmS/hxNoVRTYPZ
qyCMNKueE35/EX+sLmQVDohk8JwoWLnix0yNoefxVFd3gu3Xq6aF+L9ZaA6jOVaZZ0BoVv1i1YcV
8knJYJxGGdpVE3BILVImfFSl4PPByVKyUfEK3GvkXnsAFxZwXUqSaHu6gBk/73POmTWTrOBdPzM8
c+FszofAYD9Ch3FbgEhmjMw1lm8UanSuqOcjcu4FzmJ+UlOhk28qTHuvcYEqswbj5e0JyHNsXFa4
d/vsyQIdM3VYTpDgWYGd1LDA/1dUK08qilmgDmJStGjTFt4EUpNWLGUkXQ4YhnYy/4/poc2imOVB
kS9mFf/bVGblWI5Op74rP1+g+v0Isep8IzZyLWAOPKDdHW/dfKNaGibJ5MAtL75O3LRn7w97apb3
/BL/3xClqpr5ij6RoVlosocKkYp22jRckZ8F7KX3GBrYd/vxyb+q17oeoJS5JJ2qbJra6ucpijvs
XC2d+af4aWnVHccv2wq/II5NbutzQK27ok8fAWLOg1VeisM/bcfC8Cr4yG9gWfeIaq/aUQHENTtJ
FiK/0045fVr22kJG2UXLwqwsrrCUcWbtYYYRy5glkpdPiPOrlj29IpY9nTfQJOS0hy0n5TBSmGfO
HVENWb5+WAhr8KBc75N7d9tEGkCiNlc9dOyRrVSIl9PP22iUmpjCCFjJ62PZ1o2jnq16/mU5I6y2
LdRAL7kAKr3LTSgrl0wYjcgDSW5CzkHePFBDh07DpC3lDIc3lQB4ZGHtcAHKA/B5GLYiGEz+lSZl
y15+pEw3au/U/7JfHBc1XIHswtK8ljNwJNrsMOI7Td0hhM3Mcp7UXRZxg4YKE8eTsw8YkRqqHLIi
8cvuT5nDUYIKl99Xr6/vPyrbpiLe/GEW6opMavabB9DguVCFWJdWSVnUXY3mgJTMaklbkhznvREU
qdgAl8OVBSZPH7rJxO0KJ72Zz93aY5kvAIPEyhXpKstADp+V/0U+ptu2BqSiDwqo7PiZxCZ+Yw+j
nwVsXLhbAVR/8GxXI7wluo/N9NJQ6if6xV2jYk3JCKZ9NHnPLbmuC0CDcxSb2cYtcgK8rv5/5oc4
3kwEcZM6AGLUm0RI9WLGbyE1vezkNxNnQ4m8kNLafy/w4YK+ECPBk07irLikBJlRG10pi4R3+qzX
lEvlif6PwdjND5+K08I89KmsngKBMSsc4qn7O/QcZQ35G8KGTP7RkmhOBmzuiQj1SodEbkvJuefT
pAtdDkDkdBJCtFtU5pwi1JJAMj+b8Dx5EltQ3pH7HNpjW3DPPE5h1geHj20lA0fx9grAInV/ir/L
ksr+IcmTMwpF0+h37F+pJYEp1w1uIlhNdwxQk3tzfKVRZuN4XqJOar/Rphf8+iFle5ibso9akSB0
Mk0x+Igh5Jh5W5OAMaXMFuepN++aafCFEbWbbGBdZThWRD60IOw9Z8pHHS2vwf/mjM5oZlJesWXk
jR4ksD9SfDqN38TCw4oP3Tc/ZtuM9hgWUL6PR897XeSedEF3jZhSax6Z46JhYnWOw4991IaNjHhH
Z6BwG/Ho0YRLEp9iCk2iObJzDH4JmnivHVBhUZ/e3Vcp158V/geGxkqhbz8k/DQIooG6AzKj3z/d
NssOJHMJQ2q/x1ya9EL2KMmx6cdgQxmq30q1jN+k8y5Zwp+1cyQ7zfdX5sV5GNn/wlU/muD0ohWN
BgUktnN16rCQzQ06R7kncNYRpHEobDhATo/b+CUVqPX2pocTtotfwqJ5Q3jn4z5rdyH56WSSBgks
htue0idR0EO+lNsh8TjWSy86hB2YqI5fCxilm91+7yrz5kyi4jhrTNxJNwbXiPqavk+d9p3EKrxw
3Vros8BAysB17T8UVB8v2p+4QGszyHXUmsyCgvXQQR54XdmsPqK0tF09m6mjNKJDHO3ORfq8NMHB
x3Eq8tDWX3CWZTYV6tISvJCvbO7BzrRnQVh07w64M16DTy60NHyiw4Au3m9ETFEWkreNtbmfaHDQ
NGsbkQveXapx1fNfBWdVSP5YpkWIyTBMzJQKjujVnce5zR0jMDPqVAHO8qND0D+p1HZHU8SK+P6M
k6D6Bjuhf7ztWo8w5u7XacwS4tZw9qffnXZDaqxlq4l/6jgeSguI4mnkNhAU+gj2l7c6YktVgvMj
6/UJ8S3PUM+wUy51pkYC0HAofJmO4DD1FrLket025PWH9dzq3n4L2kEidzZqcjcv0pI8leBfuhTj
BfHS+HU4qkB1C4UaHdZiiiuHp1q9a3TzPqQA2LuHanmC39SHx7N6ST9kaAFyEZykXKENvjWD4tLz
HNSkvtDoSutEqrkNhttIMLtPGJxNxQ5M/8asu5h3DcM7ZAOHhuIa9VTSztn+GYSjMiUsyFN7WyxS
BfLlEktGV1SdPxGwNl26LaZsOXQBv4aWdR1OSqS4ACYB2lNbOM9bxszsYt99At0WTseLqLRHOUCN
CO7xKFacEvLLv0ZFgjx/QN67B7uIO69GxiltrwPj34Zx3J6wOHQnj1T8bPETdaB+5p8dVoOzdS5w
AskTZr7WjTUdJrfGFIxB+DOar6b3cbxk5VyyK/Av48BbuIRFpWi6rjC+0YvFtJyupTy5yGakYBrz
7DBx4ATCqtAwRZXA3QpqnNn66fg/coOftWJtMYRkMgSoc5zCJfR56tzp10OdgqdMnZcmZFToSce8
yvupgARputo46/gBJBkpAuCMK2/ij98OSNoqzC5ytky2fGHRTe6BkzkE/c4icyQS0sOwgxy7fyHr
fecLxXs41UdrdGa/5NiQnUO3aPb8ec10hcY8gnRCHJfG9HffJSx//CAPHwWgpPiNN/RGilm2Uni0
xOfZWMeOOAWgKSwR4+6bh/4YXeXqTPv4FrfQdL+SU/U+MusHrSrk5DE5oc+brsLrqlza4GZecciH
S25Bf5na/NMTul25b5+2bsCRBO4nmdZ29EWmXIRYcy5hxH8v6UPmbgLFlhG3mhF8faXiRZRkzGD5
E3dOi0iQprV5ypFXyaUHLU1bdPzrStK55dpnebDblsQDUjOP9NmaUUd1m1ccCgSQ1Pm96ACxBsTt
+93T2mL26UTXyQ+U/YRi3GFDIFTI4PddbwKt9wBOD2Evbclox+3hnbYiHEe0zJ1vTOBxxAV4OmLK
jIxGzsRa0tmWIs4UMz2wAGw8EmdugqNq9Ql/VRlK1+sZt4Lzicg9El4y/KlHCH4vFlXFIV9vSzEL
M1tiJ5nYUZLZDYOy8hloqU0fxbxqb6NPY/gGR0aSWWWUz1NKthuqKPLdZH1H7FZvZ32nlo++GTPs
mPOW0/InBj11i2UmPjZqyyc9a4kZv1JbmjiIwCB9tVg9yngRxwUAa7QL/2t3K3nKweLSaWJlY9g7
V3zNwNTGc9l0ttQtKUhXlwAW7MQxe7UnOEVNrEGEDP+3+He3HN5Jxg4nciProUnrt9i8GrCxMVTk
Zo2DcC7y3W/zAOf3A8IjI2oy2AhAFsxM5S6kFD6FTjqyKJVoB0mZAbcTzng8XgdzAiEkJPSMOQhU
Nz45P+73p+7/F4X44rMr8Z8t4l6/PaOxT17sgecQaysmSTENOfGOBZzK0qVrNmIIc0rsgCZeyRgM
HsG7DwgsIt87YHgKNZ5eFSP6cNeurasfAeRdLSTMIIHpL/tCUNOJiUKrGIALVyFcq5maEN/1BMME
ExcfEeppLfCcurCPcyfXC59bQF1yVLC0onjnZKVmxuOOAn1aJLz7mkCmy599aXwIU44DurCxkuYD
5kmaaixzJO+AvqnpGGGtjR0zghRR6jd/89Sxn7nTJohc9TxY4ln2QDJYI0KLOM+klNzzqBAo7ZZx
5WKiCbkiOLBbmc7W2KBVFZihIB74iOp5fNZDhp5jZYRO6MNwcI+Wr3sSPtKwu06pHE0YXhjJ2B6Y
ALizHRNFjvwo44+J/v3WnC2rqcJslvyUUvwhprXm6XuH13i47dV0ijyUZhRgCmifbbNnjOVEa6WM
U+wYxp8aPawL5i2t71OraDeRPdQzeVC+2HTL5D0gcbvPla0IXuBA9MvIAtk1uDI6MSEjfVYPXEKT
M24IULbEFCKu7HkdTsNiYLhYGvjP6rldrkYmARpE0uAE71HCUn0ZGdOjswnFAkJl58gZfMwWnRXO
+Hoen5FatKeSAPu5v+j+KX8FDyuTmUpcQ+xm50W6TYv0pST0lQEc5gC7NGTQE9A8z+Bgc8poXIMw
4oefqlUhrxYWjavjW9PnqTCol3JlbKUyi9O7wAE7U16ryELCWTWophxVGfPmYXs9SBDOwKaOoAy6
r0GfGv+ApKKRv2zq46BamS1nmvsfaqk62SeX2vIdKQhUp6B9P3lQuhy9CWdl3SBxqnUKk885CsnP
dSUXeiWoIDNfFxabTm0S7+lHhMWuCrtU7q23DUX9MjFltWO4G9yn6JZjtaIPwX7BgnJ0kWPfK9C8
p1M0cMcxAzl9MwWFNI0rCVw9quysGENebnzskmnqtDVatyaz9OxI2jMD0Hjr5hrdKM0LFioS9VUb
JeaAdk6MNh8jTjEXRb8ndC9WjeDSaMpKwfLE2d2JP4Ch6m+mClXDVGJcwhB3GwNBOHSCWLwr7HNk
4ikl50WfZfXntLCrLu+WOps7EBV16fUTKgrfUlBrmAS2bfyJhThtsJiO4biXJc6ILrlF5tNHCr2k
Nn/2pcD0WmRPYZ6iqqTOSW3HqRV5uRt0cVhVZeofrWpJHXTWwMZpyoCJvzMG+X6RmJ3U+lUjGtPQ
4Mp57D1QVhFAKWSSrgjePHpKcaQO1I4IeL4v3a06YCZu2XybVnmrD/tZdzd5L62FYvaNhHDbcaBh
A7leGHIY66Ar/jrt38SdSIYtsP3VBAKF50Mck/bZjdD+Wc7QXRFB+jpPx+pAaCyLXQiW457Vvgx+
fj/cwJJq+xQ8EuZYVmkWO5sdv/ZcL2CZUvDvpsfZqTrvFAN9PRCJ2TUbZ+zYgAn/sG27wspGoON4
r1fx001+XEEJODTnaO2ElIyD9oCJgFdW30Asu1FZKqyZVwmFGjLMos6UNf3NBfAdRk4lzSFjKnMk
rxsGZR3m4LVKhPwe6yvxiSrwL8ojD8o6zF9bACnnmw2AF9PRAbOoG2A2BEa+iLtuin0pGzVplWQX
jteTxUnagRJdszSx65kHGVUys2Da3tqVFx1+sZrh17fNeLMkp12rkSxn4WkX8fCQGGqCQubn2i42
xsi0UAcu7d0o/TqOSr3EgwRCJ4eBPXHPJG2YE62PRntiOr5is+21OJeaFq0RrHTXosjrJSmtqkdr
MySbSq05kMrdzvbQuyeRzOTabYgBMnWoisdGLZ09mNB10KCArWL9oVd8Pwsu40uYnvzKDy29wJht
+VVPJSSMPOe2idgU7KAnmyZGPJ6OsIc07IDxZAm7eUUraxW+AGFDy5F6AHSRJyIoInWZULewf1pP
XWNaO8MufrMOYlb6lsk9GrW1kmut7MjC6ySSujpmqTlVNX5LzQ+uCY1fWuzPLoQ0UjitdjLLzu9T
eQZGfly5ukzO94kbTUwaPzhCLnIbsm+vyzfLeRR44zH5Nhp4aXh4YtyvIWHvdi6pwApj5oo72VAG
G5BzAMYVVe4XgGlI2r78gfl0y2hs+O9Tj7EQnCy3vPAlw3ZOCRwVRPcSoumQZ1SY1cao9vM9jokw
zk2a1Ymge3/d69LmTxKCo+zukmUSz6vWah1kfVqruV61Rf0kHP8TdrwQzAL0eSWDKE+Ri9fXE0s1
MOFE4MEPmIh6yysET/LRYONYcgU828puPmrdAh11woVoGXsJDjZmq+uRUEHoxBcERcSCHOQRoO7y
rdVZ+TjGP4qBErfEG459uSs44qSrgXxy01Rmv0q0SsQaAd5ly2ElpY2DPCXBAQNpSlZURlBB3PCC
Czwo5H8Yz7E+aH2YhxRZ9foAi9Zr5s0VrHKr6k2cWQfaFsbyXAI4RhQHgeIRQR1bHl3iNJa0ZqII
ob8Fc7ZJ5fRBBRo7pNtp0tpBFk5wtTWydRzO2oRKXvp2cKiEPYn+v3vHNSnRr2yuV2ZCgdXtWGjL
VOJyMRFFxXqhzlMO2dBbEf/qN5MHxTn/MCwljQlr0gwvTRWppuKT3B2sWrC0ttW0najN/6eWCrF8
Kf3qmybAEaKtPzfklkoDwn8LnXjIgOLD+rfsN+qvX2MDHbI4mAecZETBQ9zu8Bmwy7LbOlNYgy6+
IQ7F2OpjZt8HET2oU+TbOPteFtJ0J+EXQ4YI9rfxtCH1/utMPjmw1Dwq0IzX3AjZdBG+eDSCSWnM
s+KZluB5Se8yb4duWb/xbUr0xYy3CKnXlf3J0CMX+QYaMyzxsukDdc2kBhNZnxqpqt2Zf8HCy26l
4vZTFibr4CO2iNYTZ0v52/mMY4Z3akzP0ULqKS9n6fK2gTWUs7xA8q6dJdnNNLGA/5EpCL40yR3k
2bH8Tv9ruBi90/Lim4J9rkRpcsgZbKmlwZpK+nBCZ7fJsXERPfqvOqjbbF5kgYQSfDms4IywipDX
D5nYHe3vcZ8+/DJeJA2TpudeNH/w4aBFvsyJ5C0rsMZObsiaVBNgYbv80hLMDv0v6yZQ4j6TTKKo
XEK6aT4sWnjLuvo4+vKvFL3lg6+Boct2vfsHNgVsB4fEllgSjDUz6G+394B2jTJU2LDcSR6SZETI
FulO7/y8C8piPrsnM7v6w5AWJ4rc139byJ6R0Fh548cBM3ZEgrunOtxaw7EmciW++Cn94Si0CVVo
iSNGNJvF0YDYJXOM4UgjMBXOqs/JrKPAO/cNdlTGMYDjXegBDDF0ylCuNIu1c1VvQqVR9NMR+NqJ
5LE+uXAcDuu1NWPv06Q1fYtaC48ld2OyGnJDxIW+bPRmmPJxLSIwaaD3RqsLaOhnjVN72F0iR88q
7n1OrtopMMl+2lnfTZglfxsEUBOS4T51KGQSlIZ1ALRSKUmFXgZuWr9AbqnlaN6LR+iN5ICFVXoY
KgIp/rVvSoxyenvhE2yeWz67Rw6RHAzgx1XqbgvXCUZzt8WNhacmxv0AQRy6yDPBkUPwcuoq57jQ
8I+8foBCMA25xZ7pcvbqfTkuqHwVNAFyy8oe9it1ryet2XnpRMgCIVnBGhzL4m/qv/ZFOw4jByBl
16oQRQqX2TJX6iDO2VZgQpOQ0FAVsnXc2awFrELeM7aivZ/J63bMWYddrtaWuUha042QRuxqZswT
dL+I4NojqX9jvajJWbv9MJQEvTl1mBwVtMYDfVsQ7yHbaPEW8QWrYmop65nlaGPpDJgySPF9pS3c
zfIKAbf8YFkyQKPyC3AEc94Wj4+e95Ps8NEGfKorR5WlTWCURtHfKQoyslke8Va7n5RbUFn4vi6X
tHw3rTxBPYCd4P9fHrq848Sg5Syy9ztW4+3EB7EsnLobHxFMwDw98iBsqGJ2cKd/Aqlr0fpOWm6t
fqbJtC8HJ6ePW+fAQXIcOoGmNuZNDNAzHkEq+A4lZb2aVyB6IUv8tTKTum1V9dFm7Aa/j1DuOD4O
9yL3LIDo96WDVw+RN9i7OWTLIZwnP6XkSUyPbbuCXozeobCHy1zPGLib5idGqKnQhoATZvayyl0T
Ms5xk80tyRUH3xrrfpLsF9nJoc7JKpcIw8anorXIX/cpPXzJRnqdTm7fNr8ijXHRgqTCI+k/r6cP
yyOqrf+UodCCJSp4z2Q37zmTPpYJRZBfBYPMRJJseVPxw+r+HlICLxOStR5SMfo4viVd7oPf7ZBP
U/iI+IHJaztNibg4GZds6e9nl/4sctgbzzO0xSc8Heae/2pAJQ5joMFjwjrdmKz5nY2X6HaXfpvA
Ch9TWKxl1TgGCRgJ1bGLrRSR/pi0A+Dm8dlFz23Hb7BXen5q//fDkN36V89vCQ+Tdez/05tk1/FC
w35fX7ahF+QoPVP7uf+CBYBRSLhlrQMHHehsPZ83xjQJYl2JY9kPKdLbJc9E+Qjw83P+/iOwLWfd
5bSeq89Bwsg0rbyOJ4HO8lhwgtZ6mURjmV4Aqdn59ruP1hyxr584inMVIuO6BvdVdyrLWtbVag9J
7BZYwjEOvBDiM5hCscB1gnpAwTCdqeP74kcCY5O3c4f84Fu47pwjv6+uhqJ2KEbvGtZ7qWAcDFYJ
I+FYfQMcyXr8cLu+bPWnj66Z8TCCpYVS88zCDtcEY6WTEq76kDTsaQHnBSESw46X/H4lSHVGiTfY
bKuZHv/dWslreYXktdb9vPGz2PSyPqUmGqY5WWfbPndKB9zhW0nRFOrH5G2YC2YpWM8RsfCsXwDc
DfLkdU/Losfy6vOJkco/cjiiR+Hvc6ZbJvw5RErUY/4dPTdE6kHN8Gokzi+stKyiCZX/9BTthAA5
lpIH7EUilw3do+vPCy1YCrwJ20MpsnDPp1ychYY6WMpVQk5Z7i2DAgAUGagVyYYQ8O0VrXnoM5u3
Qk73df1K5ZuUH5S/9XEvH2afF8K5+WRBNU95VvuTsrAoTsN+hYtqqd/NqwIByC4az0R7t9dB1Neh
2l6b4ND2P61dWMBao5xKjjIpsHLhvxO3cXIIRw3bvypPCANrU+rVIARQWiSD9PmMjF6Zj54+rMuK
DxoBoYeEYXXqfvTpYK2opEfy3fcyM0aL7eIy02c7iCLbQsumIdGs0bHz+nCZwxPKSWpBo51oXr6S
KiOkGDR22osrRIc9pRR92VEzik7PP47QCJTqf/c/xd9DHCFq7AleFxj8kK3GA4gXZyL4oQXXhXaE
/I0Pj3sS3jlOVHs5xMLS+1KzHLmNG+G/nFf5eu5hhehE6clK5PsRVPkCVPXD+D9TODOIoCph3xTI
R+njqVCyD0Rj1TjOHn6DKjooekNSQBDZP+2x7OQFMPhgeVfCGf48C4D9SrkvvYucwP4JLarBL6GL
ZKq5RFMke6TwQtFdyAMJMJ55IejHYbNj+rBHoZ6V42X6J5rfmUCJZm/KsxBLyQtAvRc2ENUczM+E
M1JvYNphlK11cFTLGj6vixMuOvyfY3ZQJsPZDrQdAGnE4PwOFOaV6Nhqx31+HxPuvKzKpp/m4Oux
86WuaR//DgaYhzfumjIOixi4Z9O7H3fcqRqfSeRdhUYE7NlCwj85APx7Fmt+PVxlLiIbonJxXuCS
GRJuwgG7hFQhHXlUfjTN5/MEw7tYpKoC3fXBBp3uAEqscyMuzVO7qgSJFW2aylRLrJfkVSukc2E8
EGyjWhh40hUTb98LbvHi4arOjGtDt6axfsFacsn44CU7TakVaj5bFh3ZlPSVnOmZlIQ2XTJqIRz2
arXl9NAaLvXjnRlzpxDQSOsS8oYLpp60Ple5Sd++tKkCFKHOZzpxun2I8JTAkH3PZ61C18pPv3+W
7gtEeHXhGx7PO3HhCGoB7DZGoLgIAbYYMQ3G2n/A8CfEXnRLyf/KHfeVrYXcT1o2jhoPGgj9y5Kl
gSTei/QYaOVkeZdI4PcszbiI6akBv/dBO4Z8kSA26QVBXv46MetxUa6FGv30PFnxYTl/zrOHAuzp
OVCPAHVvtEmNPVTwWKwJd1DJqzWv8k6ddc7+kxO6GvKly18BLol5RAx2df79ysyr90ZjZrQyNdzU
IvoE+TkJh0qunPC3MwWyN0nOzJvHTeYNiORd7gxESwS8116soBavB91S6pFp05nV80wT0J0xVgEq
CXiBQB0daQplRnSIU1NdngnW+7xk0NIXpDe9gZBTO6EKeqMc6ooyKv1pkjy2p5QVezoCbqJLT6rz
tqCfTNjNSoBfB3T/A8ubR/EZ61AoslX/3Gk+1ThIiI6DsPwM5QUpwbsA4Hycjoh9EA74bNaexKp4
fl/ndBfYC55ql+m43FWMH0iBdQ+55zNJt7O7ETZ7MsYudM13BN5HddyYaUPMBv40PV7TWda/1cXh
d9DGGXevCIdon9WF2jN39YNP0j8BG4RLjsNMTlqZnuC/9HRxCq7YVuBGwxXPJROj6O0a4JSXfoKa
PX8pHg01JJ5HiMh1yr60osjIv9RtTEvyeFL1nF4kdD86nBvFw/mue4T5jkxlc/XJS4bGphwfK0AU
po6jf1ObO45YMJhu+NRFpzheKHnzQMWtnzo1JhB6UOotdyMIAe6zBgsHbwCf/4YfJYxf9fza/QfB
/Y5hAN+7sd43uftugz7TRhETi4bg/3WxXTOJS/ye+nGdGz6Kr8dDXGPTmbPnRv/4+QWed/fiLXxs
AVuKbZklWsiavIGmt52o9kcJSC3WmekW3UzSIdvDMDaigFPcvzwD7Vmg1d6NvQP5CaQ+uM9QUf+q
JeJysFAOvOG8cMq3h4ArLB4Z3EEcRw6EATUOUMqdGSFcUhTapUdD9GgQ7aeW/0nIguUfqavySgsK
Tvhosnb+/UYHUYjgwPFSGAX9MmK1xk4upmj+DlDjtbswHIEnrhXnzKgLw6X9zHrI9NOFEobh6ni1
Iu5c3PvDmAwzzGSqke7EOmVKtooyA1q/QxsF8z4tkiEdHR73HoWLWUtZTNaW2tpIfbl2PVht2BMD
euERTWIMwmU6NVUGW7Ho4wcOcWRPQ3v6c6Wb2lOybGOFCgqdyIAaMLz4lnB9yBh5OQtvkxgCt1Z5
giUaIhzSFcHU3kqTGz2x/tTRhtkUboPWagdcB3Jp6JkLjtxR7ARUUIm3nleEB6fQE9s0YnUuvzj+
HxKQ87+18t92nsN03V7w5FoUEi0IY9cemUCCczXm3mihh9PsjlT/ejlW+uLQxxoY2/UrYGNQFwuM
vbdJZaiUI9xkmAJeOkxh/qjuSZlUwPE50RolF0GHesnM4RUvqyD4rPBA0/ZtIZkMx0BLV5OQvntB
WY32/x7jDWpTx86kv6RieSetwnrlc2csAXnYslCWV2H3HnFczkbbslWuD03gFqp95i927JH9GA5W
9oopk+a2ubHilirRZbMQDiWnvUc2Hee+0CU3J2dNvNRbVNyyotkLo5LsOVLah2q3q0z0bG/Lxddw
4XZSaEeBWPk+ltqQIkCa46L7BmC21cSQ0mTeS8OG1ArTuN2YgKB3bDpIJmrNht1F/sRXelJXXzsd
ihj2P6j2NWuodXxsSGpuMDlVMDb4SWH5iIOJijhHdRCl7l9G9C728iAoeclWkpj7vH5o2YJWQ3Ra
IrVSLf8x7X7Flfr6KZYIKFyc27LEJe33EVjY1YWOkv7beQEEVVHwwyaULSGQU+0RAyuSkSN8/vIT
2H3Q7aZ+AnZJ39sYwxdULTFNMFy/g3IAkYBTtfLsE02hZ+b6KAaih2fTuQ5nFgky4cafZxNLaDnd
kgUm3MbDqV6717LIxwJle7W6Gr2/McQdqrv+LaYZBnDbbfh4dEt3f40AnEEn4afaujvbkdedddAK
Yvw4aJphHc8E9eUVLDxk1NQW8p1edl+/O7935BhLuaMebqX0h8xD9BFM+9CNhan2UPVko3ssXGy8
2FtWX7ilaPzmIENlnLBtZ7zpJG/RLxtGDAi1YO0P4lrvZgFGoQfJ6AH5aDli+Af3JILTGuZRJbcq
I5WCwrzsjuQhmyWCuz/fYxm8l4uR0OpJefdix9l4jLQ2I31UDMTRVNpXZnAWz7DFOt8fuWx3T/sm
0F44fV1rS1OAIpwWjYKCJDsVE0OIwqmhu7JjQiKo5WwSu1gn3FfSwfHCoo3d9LaQt7A+tbOgdZiO
sqpvRCQFA4JAt+/4ADrH5ICC05sseqkMSWVYzYZJJT/+q1RMDNH5mvlTO7Hk6DCC1cnMb67Kspjb
vX9Jd2Y3v6ZeYoh+/8e8wxNLlkEFhSNDjx6xqw2ufvXSosMHrQbffioArgM9i4dsf3OEfO3TLGpn
j10xfSojgvaRTl0/E2h4YNRqHFKjKpVAgnIAXSkoS2OJQFlS/pJ3qGtmj1TcdhiKqTBplsh1CcI0
xdHXLkDuXstUH1A7ab4knmDnAzX6p4X1PD7pCvi0ZqAzCWXtjto+hckboM0PoSQam1Q2SltH3i+K
MIAN+IeglANv14OxmkcsnFevu4jM1LK56DxfxZgtFitEtnWlxd5Nemy1ALDVQmvslQK11l7J4im1
1OxjptrEMCSsuhrBME0sFHhJJ5IhA7mfyPaL3cP36IHBV+bF3g+mXqHPtS++C8v30qSmc2ly7HPW
I+/mzbU8Dg5d8AE33NnuW9D4QnWKfFitllmuEV2IdSUzTA8sHkQS+pBxzuajNEyqve4P30VgYT8p
yTVv715Ctc06/GKBO6Ofm7sV4kdnqSUJSYeI3N+L0W1KTLDBUBzXHZ7+oLmAO4yq2NslGQQsKffW
FU1TN8cdDA6C/k6MbM1soEY+aiJLrNoj/q682JyEvfFirbuIUraoqSFWmvy0+f5ALL9ewYBqeEME
bF+MXNL2eqrxkuQdV5Ajc/DFuGQ1/EhouOt7EmCGh3suAlXILqk7y6YZVXLXJKP/pZWaTgfICegY
+cmNc5g8owHpSK6kO1OIF26Mij8uyEvFrqGSkOJJipCuMKq+1zmQPEIHdpj/aJmvTyczw+3DvLNS
/6zczmLOADajB9UOJvjMG4G5hA4jAWaEhizD9OpbAawFwrv7ggSsGXU7nb/lNBuNBLzT1b2OpVdB
gbaDR8NjiZ06X6SIRqb+V+1I/hQ6tevSk5raRywdiN86vjScjLbnhlqgcJZnW7UMpnmmUBvPALCE
5eFYHrSBiIicB8dmPeAw8ivpyI99gOIEyIf5yVLt7JXJbRO92Db6SXiV1J3NcqK4b8ghmaO3Jbsr
wOnHv17Hbswvp29JdzkiJGB7xbgpi5HbL/gYUDaJWq1J2Aqjm0l4YUuG7/f9cqiMsuhGRbs/3o1l
4Vyi2cRgvd48/cxMwCJzTlPfRDNEoh3+4JjWTJIyMwUfTYoTUzNiKlb9sO5AW5ezXDmdeokuA/cy
sXTKu3IOcxH6LneU5rYzTovXRvD0loOZK/85OujD1xjBejmj+vfzSbJUlCtgsVIqiso04x9zs6nk
JcQdYxCWE3fkF0xoWnoz8uIXsUoVXwdgptGdiNKgC53OMtYyvwqEb9U4oh+mtB4ogitbfNYuLT/z
iYwfPJ5Pc9EfrX0lL+dIA7ZAIqt3VHtJdXWfPqH5wXkfo4tvMq5nrBHNOdEZ9Yo52/0wxBTu8JuE
uzgKGQ8KPbI/NJ9MhXxQ22D8yPkcvkAu4J/wXo8a7zJ1iPcPyxUh4b/Qv9ZKLM0dXIRBg6LsV+sx
5TxkQlsRrRsiLsK25nj7Z+hX30BuWUONM0kf0vJAV9AE1udgECSaKq6jlONKBEd8XVIuQfj7SzDK
XAOaaREOyQxFmyJcVgfLdg5PoFoxRgPP9lcBhQYt1KidUUO/dSRk8b+8dJ8gdxbwc0S50zM1FJWV
1X7DbLQQaR+z5Rio9+SuHqtKvdX6sLUgnVn468otqHcSWLuBIfSWf/oojpFgSm7o806Z7f9FwtJ/
vAKiOAMAhdjxOJCGp4ONkM+PXydGmK5dvFVYoIRj+N58AFuoCTT0UjsYFoNfQ0xAPf/9kaaH42au
hhpJh8n+IowpBxvUGXxZU1scBpWh+JD0CiEisqNuoS/7W0ofrFWQK0Tzwze3l6SHKwHnaZcL3X4s
bCk3ZrCYTiZNRVpQZpzDvrbB9G0jf8Jf8onre++/P0SDg+hOERCgES9Y5ChUDOdzKE0kDgP1pwu+
FLawmDuMUTK5vTy1Q0rrYpELw+DKKyLrkWeW6Uq2MV9ttsylyldDMAqo1IUeFbq8W6Q2ykZep3bq
Ha6Xe8soWHVlXtsYW+EKRYA+aHXYikkR3cPfcPM7YZ+B6BII0NSeXWnWfEOMubhh7+tVY5kVcv5w
8N2rXKSBTr9mIgs9xdZLv1rZhCopMrb/HiB7917Xp+txuYptH40CgbMdGdeeMFXY+VVVMF846zel
UhZ5V5xtEr3OE8kiO2xoumYrsVz0qQZAqvooG+EpiKOhU7BTo0C9o6Cm8kvZ4uvL4HF5PkGN56Sm
zj2rrSpA367+YWzlTMuN1EGRBvOUQAGue92dS+gD+P0LNnU/Mh96NJs90IjR1R+GMONK26tHXrP4
R4SPhiI+fYHGwHATXvv95Np6Icuvgfl16MiPWjtv6vRxwNzv+AB0tAymiDi8O7Bmu22uTWCTh1qf
74k2d6OMhzHinhN8I72igQob1Vwowm7fOE6k5zogeWQjeqZPxx0A
`pragma protect end_protected
