// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XazMDBZHX9McnWbNB7ZkHaxNrcQIQ5Syip8HNIk2V9XwEoCcJhyy4CjSNmDogkNH
zdDn8PrlvxHh0nfp+5uVOuIaXMOFY8+a+R3nNvw7BtHA7rZszbbMW1/b0Hw8gbes
T17TM+X63NHQX+cG6YCxo95KS0EkWMZMb9vhtsCrQvM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3440)
UQYpsvmC9rojabiHBMdj62f0+jHFPC1tc1bw5M7Oms6wbLfYY9dRS28YI1o4ISr6
BOPZWMWO3GYZXfvuGCZVYhYxTPRkfmAUnvWBWIUxoizRC6iFT5s265x1HAn02FpV
fKzGv52dt+jn4Kou13atr5TghF8OtJ01q2lOdRLLYBAFjo1LFyOtCu3BUORi5vSE
mx4ZbWHPWqqBSuxFhgb9qUBjfKRnvMr6dOOZIA9B2SVJuftU55Ip9BwzOzpsBf3P
NE7Sy1YpSpHhIteHVFIo/zngYFcLeiBfwnJNoweOswhCf14WZGfbGQm9fRBqptlW
h3NRl4lxsuyGGRXph+D9LPprX4KhbFYt2Icg4Rluy3Oeh1Wq+gbAfbXE7+ebL6Rm
8+R8OrXfEGvqVL8Y9642nvanoYAH407NzZvQzvBc5ZgIg5bVrD3FrzjWCRiymphA
RGMX68t44d1t8BUjjlaf4FaI588pMcs6fEuGJrNHb9whr9jcL84W5irET3qb6NnE
GKEf53cYc561XUyAqXNIl1eiO9CmURHsSNC1nUxG/sqepJcpJLBrx8SnXowHxT8p
b1eOhxXUYrRM+4NhUCXHRRts+z6BDZ+zLnxO29hIqQJQX8mEPaYMeyiiS8Y7TA01
iK4wnxtOf3mug6UaBI36v9bA0gA3Iytz6D3wlvvpp8nlBfZAo9Q/+vSi0/7OCMSn
xoV2Y1O7Mv4cisfzPMX+zmCZyM8NN5oVemvP+FgOP0gfbAJc48VWbeN7McFxq0tP
Z01EWDJHbzpGgPqO19fMFFjaK35GsbqdUEQ5cUHiD4MT8BRtAQMYsLhRwsJ/EGTm
Wcg1N2bUqtLiQaa7MXwIEJLD3Yz9A3KW8UQB1kEytXMxvMVEAdk5KRTPVXu7czKe
TQ+0vc700MhZDpP7jbe+H5lX53tx1NOHm/0r0vzR5rUy/FZVS9gKTYD2a3xlEqXh
flDwRLkgA3otTNDSxek4cfTPHUKkE22WYF2ovfe6OUbsLUReRtwdccn6r6SrAexf
vn9ANPzNrugZjB/YXOJ48gixPuYwktqYXHBhY+6RB885gRV1GNaWOOdqQ+OYkL3i
ZbhdrXSKDdprYmn4u8EBhu1cMYXFz300vPEH/vCEmSw4ff5w1Maujl8w+uJDqi60
UjDmEH5JK/9EL3DIE55fL/t6mknxckKaqIcWgGSYFA1+Fham7iA6Y2M5E58wcVLl
mIchjjT+l3+sf3Ykq+49Abbz56G508yjL687Ze4hWd35/KrYCQ1c3Xaxn3ryiD6Q
/TlgfGPPiDmP5zBQA+BpE7JT3IkNeFABC5nWMdIFlsFvEW81uFOSFhXNt4C8CDkO
mzFBB1hXsiR+o4LEhMK0cUCFbp9voM5moVLbqTVPxeVX4ccA9O0lYD+5OS2G6D0p
813qS6+wgzFcZteT/P7LLmfE1FYsTYiJj2OYwJvedhLeUK2F/yNNbkzzzkCoGigD
8uOi8VvYnDvqpBuZVkYhjoedaRFW24+sOlmO107KyeDpRWfWgG7N9x7RF2yr0jbK
6Y/j9IEz8SXqDEefQjhJjy3aQlJs69gF1nj2lk2NPOlLZTgJPg8w7S8CDwiqrIdv
JuoXskyDddhVG8wBB9HMFXw/x82zGPBlnbsZzxrTdbOdPGmOfqJrUt4afOYHwP9G
3V6zdxzj2N6JB92aLodVbCEQUPT4m5nrgG5HVDYe5jgQbKz7D141cP2B6fXkKs3i
qpi0jEontmYvuXbF5m5Q53Pv5cNDziZ79QXN0T7/0+RhhtzPVA++ncMbhJBw1lzx
D5FcP1aIauQMfzUw76gzc4jOXZ3NguIvmrN1cSroA5V1gHdFKwn9DIykhkMqmK8t
nfasAHbZLfofvLBZ5q1aZVXEQT9RI8JEzMoIW4KbcIY7dOVtm2OMeGTR08hn4IYO
VN8LcbA4ElMhmQAONYCzQrjeuCmlFx8uEjdmOFkvwpdRA/R8jiotSOA81Gh0lQP1
y426k7SeobkPf9P1Um7HGv7wBRn2+t9HGFJ/CqE3O+0wQxpVMA2JzllLkhWxhSOb
euQgI1ypOw2H0/bSbnIJnDQgjCqkoZm/G2DHGTuHcJXrIX3Tt7+7fUVrghk0osxg
KHhuyn1nPU7xvsZC0MTsCuXNOMM0/lxqpfgdFPUEEdfnMqociNrliuZ1fAYP5asZ
xKeqAyJ/gAMnUXK92VxJekBQ75cbRXeU/QcEaywwLGSgNlvGuYsC5MyZM4MwUAg0
ws01lQrWpNvDf99a17TJSq6E2DH5lw2XPjnr4nMxLfKKj9gCyvCFWHMQ0CLo6zZt
MwC4Lf0TnZ8pk66No2FHILifiB+//0nfajCoAISOuJ40S404fivfGlWEmbcMH4A3
fLXJr4gJ3/4Y/bZD0J+i9nJ9QnjLnYINXRjM9KZmHSo5Rb89JJ4DVbHffgGw2KiJ
AD55nDhfRW7bR6+UmAxjns2G8Ql8+v3fbzSQUGfzIWxiAWq4BPO15Al5YEgH/thL
Dx4GIhjuUJLDBwbVN2TUSLbhArC8f+UHutAubUM+CCn/wmDiPeWSKV3mxWgwOUPr
kbbWcO2SDMMPB1UWii6zY2/ZNB61LVFkDJlCbXqu9fLffsp5O5SpkISIx9Oh7XnB
+poiX5rvmSRxfpW/AG7V6oUeFBQq5upQd9Mv3KnzC2OO/OgyihyxiJyVi9ET6mjj
R7kINq0fQcDHttoeHIuPJb1bHoQMmJA1RELJA0iq2XNp3uzVr96lIRlbh3suQ3ou
bfdU2iAVF9H1PL04uoCyFTtWCHAi6xinkU5+E20UtTWZvcz72LWUeLO7SudT7JZ7
vV4y2hV1COB4oSwJ25fOd9px1xaDjVa/1jJS4jcs88aLW0RqA/Jl8wWvO9crS9hv
La+5YbTwUxyou754Y7c9nCvuDx1QTq8BalFhZeVBT+uthRjZId4hprytsyHtpmHW
GGkOqdfMYrFfEgEeCO6MulnhgRdfFEhNnUzy3gBNCH/67+b1gs1KR68xu4eakEsO
gOVGDlPN+Jl4d+P0h7Xr+/1+qMjlcphL1k784neslcT2/XWuZd88Rsy8WGvdPcEH
AlSCGhmauk+5uK6hx7vz3cfOVZ17hYqoMXbjX9iayRafl+AmTft/rDcv4kDcyJ32
358zQiKH+lZZlGEP6r8BgM1YvEy/lyZk/3t6pfCRk9uVx+s/1ti9lKInRwZI6uK6
KtWFLIc4I0rvSesstwvlN7zDCMrfmOLH4LpIROBHIqXrobd5aijrkEIhhDQK2soF
z3ZGgYAJiba5YKJ1Y7DNn1bsZIwwe+gBVDUZSxHjBruvKOB9/MQwb34wuJ3ltPcF
ZjkWfgCMQOz4Ms9CYBHQZxOP6BCgn3R9fmoWZ0iqaq7n0EwgaVsk086Ruxt02+PC
deCdyMl24i5ItcOdAMEti52WX1DT+t0e303vUZS9H+TVXPP0rzAVvwJqTozfb1aN
zUV74uH6UTxXs7Twop2w7ARljlbVL7sVLnA1SLrx5WwoXQniweVXGglLw1Qk07oW
gMthnRp5n5ui4sbDH+5bVkZKRgq3e0xpWRJ+bVYcMU3bTpCqI/wuNQ9dTx7+sBM4
FG9sMTcVpCoLXwYf8GD/19aMBGYEMp4EEsXp/ch73UrMYUMbNNv5seMdPy2NyOY/
uitZupp2NGAueQtA11iQDIZRxEhuySzb4DmENSZShyJU+AGfwixeA2OfprYDuCrZ
Mmm59D0tHnBgrZxAHqQ9aj4oUjb7BeiKeLeg/BpzuXWQOX1fNjcQ81Z/+7lrbbC/
ZPxvr9janlrQdYa0CDaj8suq5OdZDwoLxmCpszkJPMl7tDQ26r35mOfxqs74zMqI
95ivnWwRxS1VmYqrV5/5gC5KQ6rGWBUekXAfIpjy4iehwEB7z/e+6N3PN+pUZIrY
b9ekQ3oIizvTIvd2c5fKhJQQsE/PR9sBK29Nl5l4PTQCZzaJzNcHYiCfcXxOKusl
9ePVn2O87miLZ28xhgoG6cE6ax9LwIWA33NxJilYUYzYwq8gXDLIgbXlAFi17nP/
q/VSLXgQsHROScK42jed5e5BnJm9rDV7veUUBD9GDdzgiiyAt3gzDDsKiBum0ZS8
WPOkkfQEmcQSFUsh/eKFi5CN2PmTIOvdUNZSk4vHwXVPytzRwQj8Tu40pDq+mAut
s9FbcC6SoAG3vhJtg+HD+X0Q6hp0Iy4Xfw6c8NMR6tyUXJWlE4KPDAmspmrfc9JM
X8v0ZwxtNjfxCvGf/v9l2wqMZ62GvYrmQglaXBZRw2f0EucUGghJ5X6O3OjfsaqG
G8ZZGXFIlZ0il4Is0nSjncmQSr/5Sn1lN856+dbVRCuVgWBUzPAMokkk4mPacpqG
vmNcmsUTzrfKC8GGhzXgrONLQg9nm0aBsWxX9xICKFTVy6tb07KQbrqagaFw2jDU
H7ZEmafagBjBZEMYCjybaHOUL6BCGIgnOnBKK5O3GJv0tdTOAK9qV2RGrDK9giPI
rWVY1+EQSXn6LVKl6nWtpEqQGyHtIHOqtZJ3PClM8fRiN4RnxJMlmYHa8CnJNV8V
ES9vqDytfNvPyB7oXrGP+CKIHdpJmGR1hLHM9HFFUWg=
`pragma protect end_protected
