// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YB96czu7nOrS/s5o86QqDVJ/Nyrz44+lFLXM9xObqq/dvTC8e4Thyzkf1hwezn1F
MYOY0PcUzAjT2AchylcccPXurgu+w5JeTdMDj6W19fIa6lRD1BUqeexgKpI4qlDj
A2Z7cNJS3uQ4vp2GRHRaq+DdASUeqbGA8l3CUYbT7Q0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61776)
w21jBsfcushmPIkfw1Jr6YHRNiIqaxMbDoqqM/W6hvXZMgjNzn587A5QICXHikar
0oJGMAtKA0UQOcJDGi2UojQfsnJCkf9FnI+oCUkcxlj5GMt71UZoLz4J9jCj+mt4
FMOWUODgzdxvtG6X512M832T9upLFVKQJaP2hSK12IS+0AjJbs7JzISVlIpIbZON
FDAomDS/zKIaewz9bnkykFTLbfLRluQA0w/aDpFPOyNi7pgwOvwDMiiuDUASNpzE
/+i1iKXwGbr9VFGp69yp7fplHUW7ce+QOVfIbGYKQQHhq8X/VRUE+e0SUvamtA7M
sPYeYn1JIkF0ihJNVMjSNUdSwO2sdWF+Ss3bhgKAkuVNKZRTRFYP0ANo/3VeBs01
g9cy7RGHw56iVZdm32WGuXqqraOVQPO4LkHVOG/nRq0/HkWFkYbc99Rorml3fDL8
t1CgFexLjQO6/uL3nGICc0wu+ZWjb7ubCIs7c0fnYAnirCXF4NZegAVFQko4BIe5
Ncrzo7TtAev6AIdoTo/bzDwW683d+S0orFbyFqqLhNPBxM2vg2UVxHicIOtYQccc
yj4I/MzaOJ8XRyeYVtf8c2tToPEZZflNGJhBbbzQz4SRMpPbFeENZ1mcKzspZKUc
2gx9W9Ywl+W5Rup4VNZn/TRnemIwWDb+6Rvts37H8gxKw8BjfWWUx9BVScvuN4Cq
dFYo3ojKHSpohASe6IjY0F5FL5GXJHoTUqvhYzLxb973P+qhhpQsIbPShrWvPb+d
fYG6iL/veSwpEZweGSUFUpebCj1tY8wtQZQOiBUejgtj8/airI77AY/RbIjU27VS
hJo3Cb6zdWPW5Y+8hyMYh9w+01dCRQgMudivbQPJHah5XnHLNCIkXOBNNr0I/6iw
oDq8UxDcLhLpR6z8YTuJaeRYDG/Ep1FYChDB+M3c8QhBbm59Nd/cSe6IEa+Q0ptb
G1y9IjM8u+JAUXOtDB0kD82ui6BlZCJz146pcwdpPabhDMqJX+VlVk4EqXlG9Yhr
HmAyHvTwwACjAQKZtFSlUXjUPDN7oN5uOIORElqrAywpSq3rnH4R87BtcJKbeNJP
cwH/h8iWxHSDKNXdYqAkvoskQzTyR8XVKv5DcsZX8wTWriAzEPAO4oVCmZF8KT7S
A9gOkQt6hcqSADXE4LeuyXWA1m0NrQE5rP8wdA2prhPByXs3jFTLJMOzaDnsYfa0
A6bWI3cogB3hq0aX2XuW177h1sOZ3yTqXKQpBt/gnxK/u6mwWsDmWgCeZIigxaGI
tLWKDugLWF6xaMOk0oHtyPpDxuHw7dyazxMX7XBud6C9vStnchgTb1pqZ2meYYM/
EHt9IS1pgqzJhfPSs+O+dgY1kirQSIrttn58oSWllHM3pEA97tfATmLj2tAfI2o1
XWApPYaH4O8gR40MXrxF4k+8vs/I3PGfrydNg1TQ9YKfFJLe1Lv7JoRlhDZ7p6MY
+Uc59jLmVPSv5VwRo1INaztY40070/ivbncAIzcbHzmonQEBsjP2OejLB49R/nWs
lV/GYe10jnH3DM6cA+pxgZne01M2PfpqhadUbIuhyRyLY29Ib+lFV6cH0WY9mXF6
hWPVblJXHwtDWrre9p5Ki1cICUV9Rxltbamp15MVCL92HQs7fZxo7RCXUnvcOHTp
KXc/F1MQVuQwO+HkbUkRxnyOzsTFNiXPWci/9j6gmRrgtrwpMBGof2oLRG4JU6Va
mj7KBK1rBsFHT1ycF/MB3JleLn3lK4OopfOomUglsY+/frOH3xncu4pn0Yz0DW8e
vUOR3+jhyiV8ky3LIyCRiOme6Yz0uw+1jPTxtQsW6Rd5sjl6UoegACDYVh+bNg3Z
7e/jh1X3Khi2M/oVHT73Zn8LX1NvW8EwYacSldceVY9rX/a11IfceCpzNLRqJFOX
tWqGm/OGmC1cNfx0ucES/z0+Kq9cm5EMT6gUbBSo5JZNfpHmnJbCj5ckckl5H8Sr
zqW9y0RPouNUnoYlin6jKwONhI+F9ZWQ8jOlF+NbZA02a3lOOF6xfTHb1OcmhjF8
Pl+6iXHqEXvHvNrQ6XXWFIHoTDI152WohN3gYuyOpJrYlxywdqpFdVtutLLkLzEv
zvxzXEOr6Pm2Z50W2g1iPmfku6nu85O5zqah++c41s41TyrD1z5/7PP5Ud+jhbml
EzEMbOLEQeEckG8li1DGDPy+9n+hpngHvDzWWUQjYzHckWFnjTGoRqtwGF+esbSU
5Am3ybXJQ2Aji37qQewblVqh9BDUwwQ17N6cDYfUEDLQEKcZsjTIkdnbQUQxbCAp
WImzPzXAjbVYwhtRVrLalDaJqhyitp8CrqMXEkGOwUH3CdLoboQDZ2kzt/eDxzIQ
4mXqjRy1LHTjw6AQMWJm9f43M5Mj+9zyxfBfRRaIj3+ztv48/Q0Hzvk4iV1Sn4mU
G/qkPFUebPC/0vbev72sDQErGwdBRooO0NlDBoGwCoirQ7/OZ7aKDCY2+TERNk6g
RHutMEKvbCGxEsBOAwwngcY9kVjxZxLp4AnjESR/Q0kQe8rP8VGAIUkkAFWrrbof
ETVkYyu+77B90Avo3ep5petiVhHUxmqU0EZYqCcIgPgql3p/vY0v41MNO/ifD7rU
TkiTMIy6XXjWr2Xuo88TlYOK5YzyNEbgL+OB59KqHJhGqAD9tV/sWLpntlk/IPno
XZwZQzF59DbKkhCZlS1NK5abK1xmjDQesaaC4VztIwK88dd4kA9AiEqvFLM7Q+Oj
epS7BC7QLJrSqMggx1Rr5/g5vHpnHgZGQP2In8sKpviaXDJVy9fGUrixUJa2GBNc
FmPZOPrFQRMMVSHuvkUGegDHZclZyOE3dWhZO/AZaBw/8h+mEHWite92/CSgzLyY
ecMjc2v9smFdGZdG6dr587lI+eLkG7xrHHUTQiVc8zlp3+AWsQHAMZptbU9U3nKZ
E59HGs54NEDM7heF0pQ0DNfU3VDEEUG6jsKQY0m5ZQuDekoGStFkWHJJhdFU30vu
WLMRomr0TvU97TcEtdwC4JFf9Eh0hqfatzyW8dPk8xcH+ByATxh3xWg/UNp7vDL0
gzB1aXbp475GQdMGN2ZfiTwvqC1N6FpIHbk3HbXgwoULcBP+aibS34FF7/Hb8FhP
he/i4cZL9vVALV6+08d3roVOgUVlGIxNzeA+Ed1rEcqwLCRoOukexCcdjhY2sGJP
YsLZc7v9olSEJ2wxObe4TKXpr2FZ3P5yP6PYSrfZQdHsUEERhVuc7EleBcNjAok6
3XjKrZGOM2lVJpruRGLd3w+DY2Qj9tFv/h5FBquUQYRTQWESpnnul9Z5nSbt5oSo
Xt5+liekmZKGQXXI38EAb51916DFE8Q4R761C4phquU0xhryVo7jAagHCY94J0/K
5EI+6JYskg4igExcwI9bSv+/Vxk2uMd/DPiD2YgVk6kh9QzYW+Mi2GWfVWTD+Wy3
pzji7oORGFIr3O55HG0c18eAc3uhLfCzopxB1gQnASjm9LE9bua3gkdE8FhrVloS
9C+jCN9PjaKWaXRJhc3cgCuGrKsXVaJvADw25EMpIy8YxW3SCJ+KGfu6zX40yMi+
Et/XtRd1EdFE7BhPIT8dV4nNveng//5KyZmvukN2iYNKfT1EqXRu2BgEK6fEwhRa
/F3XBGm35zBeR0raq/TA8qZUtxRj0d8g5AnHNc3HUrUnSpbmgwwCcL5LavIrE2KL
F8ZYgztNkpNR1LbgGvECOJB9cz9sTxTYpOsim/CcvDiRy5GTuGwh9F1lAeuBMxhn
fQf/rwrdjuof/UpuQjhPp8l+B0zfYAF4y1bB6VNiDo0MSVMh0G0xMOrLbNZLdJbw
Jbbq5boWcbo1eU0IsVAdXBjpNsAd66c50oIWhZqdXgQZv1rzPKnD0z5Q/bhMc7YO
VSwvBNVWUGiBtmg1mHmUZIzHEzEui1zeAvTny6OazCu3z94faX0TlWOlVj+6M5t4
furj9NUMMBR7aVy/OtRQ81Vq2s1U162PfLfq84JnoXXGvQ0TZHGg0pQ0yrgX3aT+
YJX6cK0hR4lPzHfWfg1CY705JXqfaO9U1sm1ZjbDMGEaZ9dvAn6aFUAMxJ5rB7i6
CsRIcgwo3VVGD5sNJFNQjTNu+DyunZSkuByRHTSJF44eWuHCSRqepuJoIt0fr+sd
hYvv0VHysB+pjyHn6dK3ZM1IEOihKIzVLNKY7IuwLdd/L31PIkc+8rus45ouvPw1
1mA+Z/8NqMSFRFNrefeVYAt1z1gXkAvZhIuhfyofZ4Orts7YNe0HFukFPwRQRKKG
oyH+M2IrHy4nui2KpHF79xE18gCuMcDZb4JKRNs75AlIVCmjjZm/PyEQAKGnm0E5
iFdSbq7Lz2EyA/DDChdjlcDte+DTo+xLs3PnKbySkuLea54HxfWgiB59I2Yqg4rm
xmcUS0PnHP9gAKhp72UETPMcCmTMr4j0YdRFYsOkiqesqrP1MXRDUtopS5ETO2ct
+KJzryUV5wpQpDrFLe+dr75cIYBlPyGalHhUChvsBcIB70tt4dhzkKdG/fBUNvDo
RkhO0mthrEEaSa6o/xb/OOI/U8TNTX+cutIcSaur0fct0mNatSwRbgCvTT+B92Ab
IWidZ34jrCvSVBpjOtgq106GIDfRGJxkdlawnaCCk4WzZYT4vabpZuoJKK6Ciru7
uqqsxa9u8qjkMQnymRRVIbb6p4fkWHoJC6k7MF7UPf7tpMVJPLNgz0P/GjDQnTAT
iZk04+VoDSLiwtSAgCCKyVTt54XJBQR8QH2iYUBTqI4TsYD8O1gHlRHAyE+WyGGG
jaI7YewIYDfiVET414JqBnkn4+avRMPmNvFKlhepI2pCueL4CoMR+vUAFReVBbJH
pkK6zna5bhmj5rHA6xA4p3gptjC8ZPpAQgne14EpTpvBXg5YnSw5Lxr2MZmot00i
pwCqeuybVUhbssSC75SaKcrhHaA7Xq4cozhU5NcTzkZq4aKoDRBZcNJjBSpuBF8L
B8m/oqc0AAzAROytG+uo0vh2lEWYE3rIuioQGO4vfANOkSN8n9AALt8hXIcbXYcf
CKLReyuPvvPnmE+7qKZyR5HLRP0cjvkIFUawNGYYgTHw9pMIC6ecUbXi34CZL/NW
/yCSbj2dz2T00fNNAorAgNaLluTIP4Sqbcc1A80XMkeo4odbA9kx21cFJJsAkEcI
2vltoeMvKMuRSVXUuZEEo9CLy34IcMMVxc0IbB8HZ87wzqfgQXLxSKeoZH9lcdr7
rpKsuj1dDvCT6REiguFQpbE/zSXIiKqxDGQO/O+pknqNQMM2oqz9d58Xv8/wOAJn
4L36nSM6agr6KoXSiRz1CEQ+kyXyXOo6nmyDGnUy61jdIe+i+vE9rjqKh48QquVR
Nai4o60/V0OiyQ3adK5lhS1pzSbJ0vsXHMhpMwH9dEw09NMf7O89BmsswLdtfDD3
fvK9nKMR7qnfkDkjurwo8Ob48fO1mygTafI9jiSi8dH1ghdtgnaiye8806VMELaJ
7O0qzM1j0MYntHdVtpc/nzLitX/O/ajLjhz+scC+gyiKSWkgquhfe/u1WNHi5Jld
3xfrAXruOEosv72TUfnI6Nv1aTnfGVKmAErmrvDxSf8rp10HyPUf68qAIYEZggsY
yOZwfstRoE3cYIMYiy8NEni+7y7SNiwESIvn6VG76RHWeK6jzgzLGy5XsXvD7k5w
esR7edTa+xcsB5bPqYtLdEOqVXqNLmf3eCRNISZ4nlzOK8mtOWTD4fxzfO4C6lJ1
A4dl5gubHzgKCKdwjvQGkUc6bPBQKdA5sRr1I+xxvrTa2vT/RO5rgImuHxeezHgM
oy85FyTPn8sYf0TkwHpqAjaNck237KfoPXX1kSDOfqT22zMT95rPO5jeFIyZbUx5
XSdAZa78l/zurB/l8L2o0hVx0WMR0HtbA1ZXLavxzqfYeCgKrOwqZvDUrPmvQtNK
9yToWySNTfIYEBxFcSh+uqwEzveFlWrVo+I2oqBUTw9ZnmdQix8fxaalprfaiHPC
nSA4gD7b7nqk75xvWgmg+fdB5hhSa0fk5RmtJgOXFJNQqo3tF0pNBYJ8P7Gmd6SF
wSQt6+iUgxQW8JC+2Z2Rfezevazk2n133BY9TuRc+RK3U6kUVB5S8Jb52dowZ7sn
A3Tzx61/aDBFuWETEL763pfVBWeKOMhgtMny6CDfcVsX5E4MReEE2tGSfZK2kW9x
YlHSj+AvWmKfxFbsYzzLep+syTB4wqeFNvuycqiFpSxpSbI06BCdzuILaXYYpgi7
ebaFvfQNVyei7mqcw62Wr8H9eeAvofkk+Pj6pTmf34gwTol+XfEOacADJ/8PYHsO
1VIMhyv4NRgKNDBIkai5N9Fm+f2eEiZJkjuv6titjBklNgAfRpo8Ysg3Xfk8v6zF
nvdmiwM8p9tsZZWoxoCxu0RMKEiK/4QfVlqIu1KxeMjF+TGfC4WwDaR/zqhosZ4s
zj7RqCF5y3CnTO5GIaLfSXo08OIRMyj6FYf8cFvRELwOCk59wKSZkWAniVgZOpPB
36Anui2A03kE9Mb0ucPlv6PG3Cdf0llmUjOIYo97aR+gHD0xGflUGAJ8c26KTp9S
cpK5yrTiri+KVu+/PHGUUA/CC5oxRCNvFN64RFuMFeX0IwRfKbNlHPU5Az4zjZ7T
WDwTXAimb14sjetuSz7BKYaWUKr1yODfwxEjzMIsHpMSm2bUTykuLbahFhD8p0rT
6HQNVrKEAHwKeGeRxpmpahkAgE8QtABrkSmgWHB9zGuxuQeO+pfE8PUpQHAEe2Qt
pSRDtmCiAhgXLaNExcdEpsBhIziRg2HKrK6tqb4YTd1ZVYjTXgM4ltOswGGqADjK
C47iQTIM7spsx4lr2/V2jn27LAJPGV17/LOJHIqpnl6EBbVDLqS+OddwpLxcAyTE
MtbpJ/nL2mVAc6PzvmA/Z0UVjwobI9/6YvnNHMZuUKHz5Pzv8F9IIfvbm1NqD1Ez
MPkzGb2RxG3gWeJ48FQxlyETn75Sl2Iht84fyeRjTBgp6Ibr/McSs941fB8uNRme
JJiOoHZX1hJHjRArwyMKC5+9Ew6CFGseFPwJQhz0uuXOmsNNLXk4DkIOjBudOJyq
+vSZ9uhe07Avp0UM+Z0j+WD1LH/Vl55grWeQB03+uJbh6BdeXEPE65Vzqmf3d3I4
h9yXdbJkqUZUmue8MB6HpScTu4xELTUx1HHyy9fN0zu8erQv672ebfLQiV8k9F6P
GAW94dhMXQn0kq2oaESi2vkMXwJ8cEwCOiyq+PZNknfnRdfkgDvTdZ8EcUMgZjFc
d6onY7nVFizMek83qTixTqN6BtvI3ezfTu1l479q9Ny+5jHyWSPrs7sr+ib4V0i5
3sWqosswvtGzmo9rxMwHLyqkCAykXk6CWnFZfeh6RQaDxZg7QvUn5zX8eBrZP6P5
Ieln7ydPITXslJXGMtcwVYZXCdtpquVBVkIAjdEPkf986A6L36qABKqqapdWNCpr
qq3LaOqZNK6X2y919Gc7ythEkIWJCid4XLo2stMoYyi/O/KdJN11k6fbumbd7tcI
87JqLteWKAN7GlBdcKfkHy2ibujRD4nxCshWaPCBQY23fwfdgKG0q6Xv0atS62fX
iR1TDNjR7n0W8VdPRMPkCGLkbNF4sgBD81VOXpxT2+LfMAWskYkh3/dZ7xWc5lQ6
rp0KiVWv5tfjXYLtGJ69W6IQGC5HVfX2vDJgJGkfnD6Q3Pu8shp+nmMYjtDNpZIS
lVtOZUcybUkM8QCpS+3TPkrReN3x2yiuF1xp7n6Wc1KKSXOlDCMaHGu2Lefb3NPr
DQnfylVbCaSOtp0ZhxCpWsVZ/GZ60qlFIXqLwohUDnu9+VgTvAiIrokxzFU6Xzyy
YLTbJYYRQBd8tqcTyT/y+LYYx7UwO6OC+tUeT30K2bgHSIcqe2/hE/hP3myzj39z
/l3x8gr3l+GyhvWv975tO6np3Cv/mHuTr9L1jzi4tIUqjEhZLMsg4FItRNm+0yRB
4glA5Zy6BSjQxS3+u/kE+qUlEehqRGEFkr8o9GCEMHfzTuXIZ+6VDOWHG03q3bs3
yqRyhPfhMXz0724M5XKwRnG/vByjqTYSbURe+VYnB3ufk6Q4fQ6nyk6TBaU0X2Xa
+J4HSfLOMJp9RctfZ0LwKWqVfSFuIKP7uHd6fYIt4Tg0MYuRVyzikMMBXauPhxEy
e+P3OY0m9AQxo/CaqjYwxapvfulJv4qCEhLSYCXkPJEI7fQ0qbzlhG26Wxe3zhrM
D5BX1ATYl7MB+sLSNKB2dxmriBGsXbq6xBaC1VrEuIoc7AqFhYHHa1HKUBVx9JNd
5+B7D/bDgoK2+lF1fVEvfUaBW30ukoP0oBrywYeB6qGRSVa/v2xkNJ4Sdr6G6N/I
bp8IV1DSfu9kNKE68y9ZaRjOEWYjyn0SmpXnU2VMO8r5UuR8FvspVwashCJaKaml
hC7fz2wgDa+ZaKbxsbySTKMOdzKVIttgBSvhjmCpfAtbemd3P3UGtjIdQ/ukT/Vc
QznxWns92RKk//xU3kylLISa+tQQFHb5wYLv6hVjb8YmD6rSpx9W6ztiDcQ/npqD
dWw8CD2wXPl1qa4uR1MqPd/uVMnyl8viKznoyu1Ikk3kNjTL9v0BORDGmb5aDBIv
bSfu6KlbS1RtUnZScVoBjxRoQyICXWj9v7c0kAYFeuKBciFmtPS9WuFz3rIPlNkQ
CBup2RA9lbwUiqh8YhSAr5ER1Zfg5cnoZsCErMMuc6qwXXuFsqtKWNfMosI9Bobj
6fl+WxJMFDgxuapc3UDuZcpnw4Y4z/2An7huWmLXAPbhMTnem4Bs8MMx4KbzHEFk
APy3piY4zkpNidjA6dtBCVf6ZD5R9nF0svtjYeY7yveQ26Fgg02CJgkPX6Z27ADJ
JkbDtfbxEAJ+eM75XaSyROcI/8p+tlx7VHPjuTl6MK2a5gNfSx7Snar+TwVN5J1g
GQfzMsQgBwu7RrfVkSZGULqdFAE0m+9hacct4jypTbdhEp5KsvwMcpOrmR9dktL2
6qX6+h3/L3IR5OawxVjJ5CElPaaFuqEfPNUziHw32n271sv7arlQCDA+rw9kT4uK
x1APPDBJO3DkddK545U+jvh9bNkE2K3k0JCSWr9+aaOdow0u7qd5v5ffntECbMzQ
XLwG44caV25GyUt3jP/N9WwxNvSiu3yE1o2PX3HTO9zTdPId/8qGkhPJ9aQWwh8v
PsA/YpfjeV2SeR0UDv5gBVAZ13gvyvucBIfDHAFNCVtUOsRXiL83ncw9BGqJ5z9f
Mr+bwOG5L0/zRgMMxbSQ4NBL4eArVW9dcKDiQ1X54kAOUkG0ceMsS3OqVATeqtZc
R5F9gnOSNDZRqOjT+szv/9UF5WRLmhYSP/9/JrR+CDoB6giKytrcgjSkDpjApWoc
wSdS5c71xFJ4YxfvLGGGdiMYGyO2Fwvx5ayS9WQ2V1jQ3zHOIwD1AWIZh57TNCaJ
DCHfgkZ2mcO3hvVAJGzPnVqWOilCLh73P6YC6gm7hbq5iQ9Dmeq9Jo8Qg0+Ltwda
Od3jTCZ0uoPimyk3aQAdhOa//qc6XueH698cccB5j7xfQAHM6oshTFxi+pUTn3CI
UWsMNq8tIwOohUaTe7eGkoMpQVMt/3BahvgttcjsBeQlqNGODV9qb2PVywyKDOrv
uV0qikitNBCLO/kCE7AFvG2olMZCxOXcvsgBaxL4C7OTeZnjIHWaJ5NfhSY+18pA
6YjDNo+FlInFxzP//ZuA8Ny2wxgxYX+ZunbEXi0uYN8J2kT7+AguEr0LZU/LrYPo
25LgZnQ6fCNb62g8l8g/Ib5hVSl8/e0l/pW8EN2h1wvJecD57Qs/98KXd+2Fskf1
3wRcZGxwpdpDeZjEQvHF3oVDTIv0zyqxQh0HeNCzXwBBg6UZ3SdNBhvxmxbt7nvP
Np/LTBE9CNdBZ5ygDRI7V9+4O/zqR2/QVpSnPXYy8RaxGs5NmjGsagDFNMk8absp
1gm8wsSlb5Ug2Ve1cr+5ag6h6DYA+cqaVx+iP0mmu9p7+Z6SDvQhNLvJAiCiUPuJ
d7rWrQ0Q4fYezPkok9VgerRYiqu3yZjx6RmvePcmj5IjqlLkoVAxLdodj12ytwTV
wIEjs1XEpY/wW9wAUyewCuLx8MSZ8tocjap0LNgNYWDz0Xx0DV6Ym84mARpbTtXR
hsJy67hdo2Q3gCzcJrrcvLUCpDjQHnMkZxb0QAYSqeFI4c4L2ZLNBuxOh1RXdX7H
htR9detQLtGnnn8pAIpDQSWbxsY6RAoXHQoWRwy0C5PUwn1PgqnTEKgImqUXkf0t
4OVnoXrDWJOU2mQMcWZR5ya5t94Fcrmgf3vnSYCZnd1/dKSV3+LIh38rkyx1unBr
4EyDEJ9GfcTGYsa1VDHy8RohuD9PwoUZtvWfssgpg3aNMVRPe6acjOax29byYKM0
4FVOExas2pbkZ4SD3aL3u2l9VGjlUPGJo0MDL/UaM2cHljDdsC6hpsBBoGpGt63u
Aq3eBBS6B24hnqNHIhaHfvwgbwxzqyeU0mZ5Jc7OFRk743SWjtFzBCrOKWLb9Iwl
4oVPdzjzWms87VYmhZICh+nRA8s/5AI58HTgdWSJHC+oFQCV5Yd7HCYIiYjPnCgW
DHtJBjQGpytN374MuipX6WU9+cwvOYICxaUQMCHXwxNwPS7vm6fYjup47RjZd2vL
aySAMvEx0LKB3nadzQtqe/aW/yW7e0rsV91uzvnf7Dmz6t01Cgs+u19SVsdRgxp2
bdKsQ4apFVzo7fchEEfMb5qOWaNqwngFUEw34458mNDOmtvdBPA05TZmpNat50NJ
HwzV2rXHdqxA2ycljrMcCwhdMjzM8MVi6IeFk7eRjrVwpwvqrEc3qKEA5MPs5yjc
p+TKTxIqsJQ0Km/6fdFGarCxoRJq3kELO2eAQ7c/CMHx7+ilz7GQMQ+BE1l2VDiC
bbeNfhIbR8qqLJsLJnuEt7eQ9xfm41vKXBivVNjvtq487b+fEJN2qQwsFF2l+jig
Kc1heWZIbfRonF/DZY01nOQN2MHV76zlWXTnhYKw8ggi+cNsQRnkeYudVqA/fML1
m8tQ/TGPpw0D15yBjSsuHqyr9ctiYJghRt0WDGf/gOSibkH/U9Srjkw1rEWW3RZc
6yGfkUkxTi4duH2ZztNlRN4TdIYkfoY8hPeF481Q6GBWGdCCvSIg8jFUadFjzOPv
yvv9PyHVCwL7zJWMaKSsUEC1iBuQXsN8I2KJkp5EcokiDtGe9v6W9ShHhFKCuJgz
R1pUMwRznlFgPTI2vzpUHNamyy5OoDLYqWGC579lJPSkJF61KhU69xV+NZI0KUtM
6C0nWTmgWhVkNx35/yG9DsnGf1xsB3TEWQmWCVHWm9nu3bzLp8vzeukLJBZ+zq/p
03RZfjVrUrHmdPAT9fqa8e8wRGPmyYT9hpteC+9gK+fPX2+2GvuFReXuSOIhE5YW
+o30O5SC8hhBwcw99RqejyBPoXuAv7qeVYjGQTq/J0pCtLPLf/qE9BZG/HC80r6y
C+RWsr1RJnbNHgVIWze0GwCCMTSMZ4VQvVMsZGswEoeTFoFzMq2WN1BLgZrgG3YT
JncZ5DGFTOZWTyZNvdvR7MjzJrVwWU2Ueh8P1bX8RWeq2dfqb0gA9jTFrpBEB0FZ
zwsojRgQ6oiY0WKFYlpshCHEPr5elwrXLO1VWZ6y1wiyPEpKsdEvP1CVcULbH/Xc
YE0sND102PZOLdasotAUnFZFZYcex7OlGSAWDR4xGtapH/9by66xb8nLVro7Wqe6
nhgeXQUTdTVyMejAHjxR30tmGOM2gdkBTbcsVbCP/XwzDFe/Wj+ZwntljzjxAxRU
wJPlDupKlmF0noLMXOarQUjMugTnPiladlLzBpOZELxZsFddZmLF78F3fvOYPfhd
Ewuva71Qt/8TI5NVL8KXJMjhqRMd9J+B8hIyRXEuvG/9qLLucdU/jq9XTWAyqSfN
gj/xQEFajZaTPwRyy1/LVcupmkwjUvBmN+giRSzfqBy4syLGCZN80YXciLrL+dLl
GrBD8yUEMEMaM7Qtq00fXwcfs3ftn00sllga9mL0/MTwInUnCM0XVAEbjGuVsevY
oBunfpwi4YwttWq4G77WJgKbKQ3wN7CFMT3iaHoQIFv/uLLbrLAT0iL/KJ4PBrc9
O14bXs0LqdiMQBQ6fcYQMN89qo1BFmyqByXj23I49/81VFwRH1vfhNDwtjM6IxVc
vjuX8P3dM9QfE4pnGAcD3KN7GgRhDYKmGX5+Nq7c9CsnW3TsJ2XrgDlKrdqWtb/e
BNIEX/RTem95EW0OIgI1qgCWitr0XzV7tTN4cp5qcSPdYNCGzo5X3gzevqtiRL3O
zdKK7pIyjfI6v6J/Ft6fPCgbWSmQ0eUo6NXpTHfG8PW5gb75ynkcHB4Dtky9ZXJA
VkLSCwwhhWDVwKr4MycpXsmii8TKAZupN5ZwwcCb4ZHAa6YxBZpCphAHB6n6m6QA
uTZL4mdt1xXDF6D9jh0kKp6Xsv2USxDJt34qpWr0zhvXImbK7Lsbu/WjVjuar+1/
1I7OsdIz4trCMk9Lw5JmNOonwcG89NVBQ/XYVJ29FR6JIjL3ATi4yG7dU1ivcy2k
ON3knbDstTERGqDncpp0uYh4TDDEk+15iA6pVONTfsPbsYalNGC6OiE89RvAHnGo
dN3OPY1wytMwsy5pZhGFgnl2HbwZQR0PYW3Ge85SrWvHk+EJ/+bivkvbZSSpshPs
8H0ghn/fbSoFdQjK3s4437m3KYE6ibI4NBBvAEAof29gXJiYYQoBEOEWccf4LCJq
YeyhxARfJEjTUasHZap3U3HAaBj6HWWuY2myMMxO6LFBl1gjPw3/G7IY7S09Et+3
cdQDLuZv5ble5zRaQybYdxcadNnBIL3Z7MwETxg650PfI1+QNovT9wrg3Oo5MlU4
Alr4lWSYVrc20viya10kqZASyDgGJVqHm/hV8HJoQe7fT3BgfOibo8QqNEHM8+Tw
5QZYTXu1rySOC2m8ZtrqsWWLKegkTglACiMUYQAe+8BFb+nhIi02lJkIvmDfQwo8
WUdsJ2iIIzKffaq+0J4M0+mW7CCqQgcxuPLHH8JELB90ee8x92wLZsLb7JTFBFKx
D4DgKMCt10Brf3DJuG+wPSLRshBFPmFUW+q6WLItKZiB8f79ci+os/z5cmf89Llf
l7uMp3njD4xdl9AcZ1MJdXrjL6epUYMEeW5D5a4qepaffUBYrUWEAngXuK3Xyj8+
NlugV8BUaPDfafHjFi/etDaR1Xj5MtLYui1ySIM6gY75kPOKg6JHrpA2agd/zvB6
LDCC6h2NqNiOlVxUyGiF+kbfm/mYtadlFQ3tB24DYY8r5TFIxHhgxiDlJjbKFio2
7TcPNdiJqogU7JBdgENtAK/PDOyyQNJxEG9D8qMONVr+pNgv9pzZLPSpZ0h3Nd/s
Grt/FP/1JeEjnAoiyTCu9sYOLsxbYOR6p15hKZGRwX6aiPqctchZS7tP9x11LFpP
MSPIT/Uqyua91WcFgATImN+CQgBxyXwaPpxxh8lYTUmFPouzbXqe7aHb/6+IdjcC
Yhs5T1pTiAhuNn1P5+1HtE7fdZMPCJOdL/dRptKOIe0MF+tdWGjCN1Sp2wppud8u
pB7BL3qBSSzEJeLpoKx3MfcnpUaHUHUve7uW3eOkOQkIuEJJF4qexxrnVzXbJgEd
wYTjZcS2SDn/7IjFs6Xbs2sGJgngXGrdhJVT2FMelNATeQhTsLLLt/aee8RcOx1Z
137ntP0jJsCWyQ/RcQB1mEPGXbBSBPBnZUaZZ0uRaY1zNvcf6ntO2WjO9CQHytGh
vUqB7e8sYB4bFnFEZpib7/hUNqYrNzJVsX+Yp3fpJZsai0kdf8fSiWd53ktxpNUJ
cUHw5fFde2XqsNYwZmI+Y0KOlkDqPxKfjZiGS/dUiYBqw8V4wYwtmisM1NUS8UIY
aCfTAhdI1FYGlEzPCsAmRVrC/RQSnoG4iiqCCjaCpn76htOAlGdugn1xbI+XJ9ob
wBXe1UzDCx+zx6kTJZm/+aB9tEI7SpVxgHxO8HXTxkgCNImOSOaSSES36VXoBL/U
3FR0sFIDuKSxiywEg922WkFrptfQigILbrVa1tK9+QAMdBqeZTXcF3RIRU+6c/pr
Er5xZGM2vNo4fuMbz8f/Wx+dc0GLA3Vcaa+vRBb0b5O7idStPvrzlAo7P/ZgMvPy
n6GdE3EZAxzqNUF7yKB0K+busf5nDuHVqlX5pnwFRk3AM6ReJkmRYnAW8x9DKNTP
0NNOV/khQQJSsg2+XusjzbyXteXnv5eX4dq1gGVfSdQVemoN/7+4InCqa56JpUVm
pCAM2ac4pTBw657lV5jqY3WpgqppOY4tY/pZeCJ1rZEtCuV+kTMzP1YvCr/HVWdT
16+lMiitgya/eYqR2HAk9/aSYGl5d/eaaEDSln4NW36xqkx5qIDTYkez2jjcA4pH
gZHEYPBCZTudMsy6m6PgmoXLvXGPQOv8FIehw7oDMfy8lnRaKClS0XpEfbvXyvtm
jJc40Jw13nz4J4CTqb58zo2yvzL9yHBkFNCBpI1YBqJumABC2MppoCX0PnpZdpRM
TN2LIsg/mLur8G9lmsyDnY1CrI9Qk00w9+M8TLVU309KpHwaKgbx9cl/4lKRNNG4
Ciix6e9AW6ANAXOxvHktD50RvQP3OUNhl1KQKZfqJLB8gBMRgR+5XdEtl+GflyIR
fbOCOsnTtrF0qrMNBm25H4W4Xfxaxci5dvvFUkcxXyuwzDYYIHVOn9ZU9JiToTqJ
soxT0fh+jfvzXBkFloF9R4CvXUTF0PhPLKoXqmhzje42J0e3qYOAPav4Mf0xYsPT
DG/KrzQVTm2f+Dd4b0RZKhvf0FYbuibRk7GFVh2rV9W+U/HamCFr8zF/g4citpSK
PnIlIM92DP67IHjm/OyeqihNxCxBtAKYMFqzUtRjNi34d5cn9DK19sGwV7fRBhoT
/FqTSqZ/3TI2MKFFfyVhI/MpkcYEe6sCsbECpkv2oxshrOKuQiXw6gALhJvhuzYA
7aca/NNaqC8LoeGT2lN7Mx1p8QzbnPdMdwQhRyEpv26DC45z1WTOCbFdoijUG7ls
5AsnJUnyiKVktCnVBaXkCwqUkUXjemAnjk3esvqwM9ET7VI/dlqCdHvRtBSdAiIw
F3CnP9dNIDGwX7SNan8e2oKZvoFFg2+OaEf5n9Pwv4i54VHqPN9dELzmMveCA25I
Y39Md+KKW6eD/83Q0rR8Xli+6izeUqHnuweyCTHjqZfKlwVhrGtiOdezIcNyPA//
4/uZxJiT63Gd9M10xFKoAr1B28QaqpuSNGDGWmIf/jFFo3s5CCrsEerlvM8+54UX
RRRI8HNPWXOT3sKk25atSBA+c82QMyQv0QH43NcjKEmRlE2OB+YEYnpw1/2Vn9h9
p2v2w2urFKyL1Dd6AMYJTE0Yj5iMvdWE//BHQAJn5CzjYXXSCXqM1ORGXW3ugHom
CrbsXnr3hdP9RWDoR47wwXcGh4b16D/RjvMGQ+5ZRFlAMAVjV1dl455CzZrncJsp
LjcrUPj80404/3lQEQhYfFCcJlZyvLkeAYqMToX+dA6ZddCHwcnUANvcujNX8vQ+
vAFu6Pb3PZR7HR73GzvYbMnahyGXuQtiopvKkceFp+0KUwGNrS2RF6Z5MPTz1Hy5
j+YEpjOZIkNRyiyhWr47eAZwdouEF0DaLVIf46pl+ov7i09Hkg3osGiwxozmvitl
PAddQ7dv1VSJR4+P8LKui1ZA+GOiYFQ44TYO8CWD7UJ6oaO/7hhAwZrWgZOnU/tF
4WXTI7hO7wfGT0hrujVqzISefM8Wa9w5ZJX/LqMPuSuwIFqKCQlE0VdqvkOBGqbH
ZFR/5hJWMpdSGLfcTKoDkiIK3Jrq8FHknQRUIvz79u6YWwU0YbEw0CQVQO6qdfUq
wZdazZhhXdxUW1atclKdfj4T0YRdewEMRpqD0R2i+8OCkfw4FmdbBzaMmQncbxV+
NCFLAHl1gJDdwnxkVGl49tRyP8rad/qR+91ig2+mggljadz6JCgbMyb+eFULisOX
48fsRoQvjHlee8vuafXeKDKfFivx2l1bd/Z3pRA9tuyOnr6bBbI2qRT6Bh4IwqBM
1uoU2hWAG348oo8t/6mPm6MxdYKG4bgNzbH+jl0LWPXLmm+JRjMgFRGf1FyUHA7j
YV7eAoh39Jq0oDTrNt9R4mq4Fb9pNB96EDEU7oyMvujwevGOH9WTr15r89d95pEW
xJ0tdf3YxCR+c5xzRK0u6vpXpb1on7ZKRh9MlLLxLKCH4QJWqUhjXmXg9eJXl0WU
jR/N1adKrZIs6xBnyw+vGv5VuZPNK4Q5Qx2YYMF8F+Cr8V/BcgBja7XTA2PQbLtQ
lUlFZmG45st4NchvXCyyhI58B3LdAche3R3CEuLn/ux11gtS1Wl71bUpu0Da3c6h
ZlsE6Ag3uP7/Gzd1yYYEdiV9iFAuWmOLXTRzmafrqKmhMoxkUg79+cGxiOauGI/x
p24Z7NDKBBTRNOfYfdQj0rCi49Z98Pj7Eiy/jErwnQQhj79sZfjeQj0kOKou9aC3
/BoOatRKCmRxATjbl0AZ2+qOnDvR96zlQKz6L7/lWcGB6yuOyunV/6EDwExkspZX
WVOaRgO0SGZMnzV5Fu3lEm1Frtl1bU6FrXGr3cHmwVHv7WIXISrKfmQAc4UrRFHz
dKOoK9vbj/zPI9om5cYls3VgFMVRzXhdIS+7WcW+lObfKNHli5A6NZvredNUxjD4
6DUjo4czxWra2sY1ej6gWAjEQeUSVsi+X5PKGL5Ldd3d7RJ58VFkSF2NxJ/XVawu
7EMVlHrYXBFOn03UljkC4MxGksSBRf51ALlACphEYXHyxjqZiz9pz3cQXqlgTla6
6xvQGn5J/IMANItVdqG+FrJzWjOOXxRm6jAPEaTJbEx1xHqBGIpAu66tDkcGVf8b
S/25WIXULymefEuuwwWnxYMPqwxsS4WdNIBh7Jiuc8NkRtVmNZ+yCfC6xp3Em8RL
hGEFx76ibgu+zQZuBr7YXBwIavpWdK65g/pEi2KMbfcsLf8sNBz3YAyAfxT5y1ef
L5FptQoSTE5mh/Sh2IgelTcWTuuvuVKaC0tkTUrSMpjHE9FdVWZjKYIEmfkvEUtR
bSaQsLGcRylcjXMQWXyEpWi2S5raznffhJ6pmw+3Z4ZJUoj/LOfLQUFV6nEQMt9G
2HoeZmZq92keU1FuExIewURgiw81Ur2uYZpAf3+yrcEdxRn7+Os9eys/ZFOIPdMv
cwO6HWxrjAaQUZ/YNcWB8YLrmFCvjNUFpFJzsy3vfz2WJSrmLDZ129zZHoQkRrgV
a0SX3DNM6Hlbg54uzxSKOvavjmxmByG/7U1694m/WyxR0YqzH/iqRIs9MYQULYcb
3RINNGKf57zs/p+BU/Y1P1Q9DUCui5oowhdcb/+xyFOo3XZKjBlnqCM5WBIqZRzL
14hdnx7e9V/RacAnX8v6RmRAA1Zl/2wCtbXuvQZVMVzhHQMuGsfXynLNAsNtJLgY
f+UbvxybvtkRvNRRu0/BO7OqibYvVb3Jm/xj5zrKlwPc/0l3YgqTx4yfhvbOLe5M
uFCyB7vfbIAuuZd7VOYT9IbuZuyKUA3BeNRhZjfqj7lBIkZ+0mJxIad8ATfPUZgI
xWrD3qYLA2P+pta8hGfwfLpBH76lMqzfEK7I1NdU7vqwmRGglELBm/4E4qgQPcmg
X5PnfHyTAKuFaTtwowqb1L4i8ec6/PSJZl5tjk1O7x7s+l0H73G9GNrN/rY3dNHa
CvQ9uG9aYms37DWVFW1x3AwQMWjT9AY8SAReQH8/miHmooeaYbsXp0ugot2L3z+H
nfBU2Sg/TEu2LhfWdn/G3y7aJTjwfBCSA4GKpMFoowxmg4Hns5tUOfT/LgdYjeVu
nTxRiEIDyZWWEB+6rX9upQhPVw/ptkFvf8SOvxsvDwSZg8+URBy0HkVq896wJqAU
plPVCPjAMcFA/x3ACiJkLIT987WuIGkWeInIJy1Yjae0RZuAZtHImA/JoLfzcLj+
F9lzTJ5JXajp4mdrq1WfrTbbkwMxnYu6SKpyDAZwNhzbdpB3m1EpvA1BmpR//ZBp
EF7rNaJclWCzsHwUmfEvUNTOoUfRVTfG8oDR/3vp70kbCkEqJxBdC7Sqd9jI2tDS
3hnFyKOHy5kFmBBd1oLfBuNsORmX5hVItq6ee0h/SBCRnDKP45h4jpnP58DsVIEx
ct+skOTZjrKSHKRQC9InfroREMVUGL4xkyuJj0AJ+rNtwM93BhSqjXouuwPXGsGH
459TXQ78/ZGwq9uo4tUGAGfRsWNyjZS+SWKHPYpXB6HG/VY/8dhCAw8mU1hWY+sb
CpdWINT3PKyMO5elsSlgGUHFW5W2ibClTpoxoJb8TC2vrZsBW16lF0Ja0TRAxb3a
coPu1mlKaLrJWIQuTfJ3SXNx7FhA+B9R1GnZyfV4Sdpz4GJHtKVaojCea5GRMZGj
zymSM0xxPn01ZJ/n/W8AQ2Z4NrLLJX8+C75+90Q0LqlJquredHIT3h5/IXRdRr3I
uCXQfO8Gs7k37NQyBKD8KeVmlCt9kbQA43kJMkHXXo+NKxzhfnn4dHxNM7qAF+gp
4zbjOT9X9Im9yT3lwrNOdGyXFMVxTNUgrr5h+SKPEPvxWF9QdaUi7KG/B3CMWaSI
V9jrJ934JG9aFJNNw5Y8XcOXm7Ra2MIdOGZse5sWCSYgJW7V7i3TVZltWPndmc0l
ryWmSIZt36i+WyV8cNkLxiFeznqvOy0JegQWAcYFhZfiQpNf3DCh8869ybVeDew5
ttVhBpGHvJh6iHXsYnN3KmNs2dbx8NwPDIvPTYh6fLE3J9puY9Dc0tnpx6S/p3mV
IczZmo6K1cHUVyZU1D7PH+6xmRkDlifDpfFj9idR4123xSdfb2i0nDHE/Ps6p5AY
43Jlhgp5In0sVJh/pf7/lmtW2ms98cTbRYGkaYsWzjRPI4tk+VGsLttZi3vLt+Lj
BWUIo/KXOEwQf74Yngz63b5U7BcnT4fsuCqGfj69ICu33V9oeXHMQr7EsFP75a1f
bK4vZtZ5mLhA6tgVn2HhloomQVKMe4ATQOoYEMkjSM6kZvb9YNj5s1F+s5Hczofd
gxL0QXnlS4TpFydm5twKOD3qMK6nK3ENpTWjyxsvRzsruuNmcdoPYzdWxdp0di3i
0TnUM3wt6yI8J0pootjqju1o3JQSl7CckOSW/LEJv66NU1tzaV5aj+qe1dVXHiba
XwtprINNM48tsQaxoUW/E3suofHrODPP+UvFTf0ICNrA1iyOfkYghFtPRV2AkhcD
+b/1hlLP0Jc7VSQ2+YClSWssZeLG6/cGj9S/PK163bRWrWwixcb5dYwDlNLAw9H4
LmwDaJF8cET7YYUafw5qlDiPnZpEg3Cx55j/7JoLrQS51JGzqF8lAkYl9Vqy/uj+
7+OrckuIjl8d0QKrEdgMuYkQUebKJ69ma9HXXllAGR3OJAr9Y4V1qHi5qFiVg9uv
kC7ulckGoamFBAH9jrr0nzCXtUIimPMKzWJJNWa4LEKfAN7gtMn/jcDKXxkoIK6F
ziU48yP9J0JnGn+QvXXlbP42WNFGlL5+Lo+hf8N8iA/Jdr8fAM+Txj/AIdkMter1
dZE5nkqjNpfUcxmzikGYCNVZ/3pXRoz6XcK6y8UtK8on4Gpo6o9hJjOWkRwtY+Sd
OozGmgbcbLyDVyE0dUEb+pj+D3xhbSVIClYPlIGKDfgJP8XKD7W48HDvoePC375g
KI4AQlcrRWQN3yX4cUOzcFPvu32tvgh3rl7Z98USTQH8GthMNQFVG+tAk7HYXPub
2yMV1/uVjBSyPjBpfmTSR3CgVcSYRhVBwQk/XyA460typxRkl6kvr5FDhYDL0cby
hCOhg/Fi3LzMbneUsGW/FxdbKIT1+/zwCU3HV21ujzh54I8OblVtiiFo/okZZtXX
vlksTML2+66kkAUDhhWQeY9VVY3SYG+0SHr2v2WIHkWkip0/EbdGTOVSEPidriot
UQwakZtcilhvdgx6Z71oUfydFZqrUPvuIyakL/x+1ckKjDD9+9362SDm/I7NK0rq
rcdIUS1X48jgymQakMBhQCXjFGQQvAEtWq9O43asEwvTRICRAfy7ToyCpstHGeeO
hzQNDSW07RDWdbMO70Lfc+ulmfZp8VIO/YRSoEGizZkmqU3NriIOEoExXukMGCFN
7abHOBwiTxvV0/XmyJBRsOl6hamG4+eJ/dQOdxXo3BjHn3ZgQQwWAxT5m+DekZxX
LbKb0yukSh1iiTRe1CA8hhrVeMU4NdMfzRgZBe3XCtbKOLr7ynqMAT6uSBF9BciM
C1qe3/3qKygWVhq8umfTTOXbPjBOKEMC3KBI5Ac3XWPg7lSwn1njblslymM0RLjN
JHxwkRyn/3FUrHdo98k7cZcEX81rLNAU1kWnkDnY3DhHCr73Wr5bUQepFEDewMAc
860+b0XLov5MnyhUoq+iWVVGwgEzQBAaJ49pnIUTcxxn6bWr/Rkg7w2LEmU3hFBf
//6Vfza74TZkLOHWVxmWGOkyWZqsKM5nTbVcfkLKV+1E6mqKDBoVu5uOV3xAkCRb
b10H/qVtGPiz99sUfHFClJkTVTSqdHKzGGoPz9ZHGZzn6y+3IpOeGS5JZQBHE1Zc
cQTlyoWS1cXfxoIRrn6tUS4rU0Jn7TjxJH0NAZTQ8JjS9U2j8wOb2n6LSB9gluxO
4Rmiug8JVTza9MMcDsO4OElGcVav9QhsmR7OZPjnod9wAt3KG9iflwrkCOS3WKDB
s2G4xYiGRR+F7vM/bj9gmOR5QaAE+uDtrdjjZkhwfqMps1HURHwNw36b8I20bppW
o5qlW2DrmSagbG/cZavptmbCATQwG1m8m7RZoZZ0KhpkLC5mXwhduDPynnnunoyV
iMA5J23THN91ai1pzEucH+zt/7fCHfiEZaAQ09TYCP4M78BL6UVgrh2gDDao/iJo
m93BQI+Yphe5BvA/nQKeQpru1sTnbZHUZwYHgnFi/enPxpunQRDExMcBLNhpMrkv
hWLdPKIb//8+vYm77z+jf7fXoG7Je6gYvTiSQwmwdQJScE0n63tYrCyvAteIN/GD
RxYo0FeFV23DcPkXw5weLO6NEQvl61N8FKSPvvPBkGPo0hv6cwf2HT41XgP6AAeB
JEeBU22oU1s+WMJt+1wpsFzuVHqzIfK2JFwzzoUW4PiqcibrV0zby0SKu76rjOEh
fPUxG1PUC/cYu/DNS6tkXDUkT81VE1zAZfuSav2AkYy4xDbIrDBZwStJUO0WXOoE
EQ2bwOuhbFomhOJabxv0/3XJcBSsvjYf9ZadR1qffiUtGFXXMs/Pdh7LpjOj53+0
/joluMLxRlbAddaymf65LiqMoR0/ll9NzVCGkG0bZtEfw3RF7WDxAjYrI+blxpEp
om1EUopP2aP8yvkDHYtbje94IFFZ1HTl+yKbrmkSS5UQ3xt/C1TQ6+ojTIkBCar3
1l+OdmEAUj57OVWg2jk2WbSTfoVY+AzjU8at1FHsxY+3nsxQju8CfQE7YH51yeUs
TImYfgzwiJ+f2CG0lmft6dixHviihpY6pGtYdWbqMeDVk+bHVsileSb7rM++8XmW
xmrZ9LnOu3SAN+nZMGSFBbZ37qFH/r+MVlh9YOJiRBe07rXxArwsdLPRaAudX8cd
0zxHJtX5W+vrJlyFcyjZd8mmQh2eAtkOsN0y6cvJTsYEjBPe51XWxpbNuEnhZJwX
g8ZfO4jwv3q11eG9JzB3o2wyFxcUruCDXLmlPKBIvG7+RjAfZViKeH7jyxsRbcJa
+QdrvFfmp4AltGax+JO+oQmkrxKTqIEcZTyy2sTf0+Nez09qT1kLQZht8afQqbLt
BgrfGI8cfctki12fJ8ARbW8VYTaLyRRHhEdRdi0cxrljpqQtK2xy8GGVFtX5G59G
08EAf4wgK6IQx0CC7b7qbzYt+aH6OMBbHUmUIKOLC/iTc6pe2g9AYNzBxF6k7UT1
i9uZmc0TleXBMaEiLB75TjZYzH2iXpCMe0s95WQ5QsNozWYUMjzDTTwS6igvsGYs
wwTG5/hh17HR0VPDC/geW5EzAoz1jJXLKlt7XENhDcbHpmI7V1lxRyChJuxVQElL
h/N3A9mL7tSsZ8uTgl282GpI8ui7LQMdEgcacztLCAx/+5GFgorD1yqP99+jmESv
Vmbb/bFMmWFeZQGmLCOExjHEHOg+FByNEA29KJYjRVz+6XxnowTmrFum8xgPpJyT
kF/cXmlGufXgup8YvsKVk7qyeWvaThaz64dpIYSLq2ibdpvEwoL9ggEbNXRLJ7/a
wIjWq/FXjjaaO03vlLZsAvBqMMYH5zaI2MlVivIO3snBxmdi3O1PZd1CJPSuL1SW
PEkvCpNpp6b3SnT1IkvcCYWGh9tfLQSr0RhjUx6424ALmS6HgS5OwZm+2kJNvmAe
lqQtPecZi7Jncqpta3EiA/kXEvuZk+aXoJNPEzDdAw8cJAPJ4ZGfA4M/Ynp3XAKc
/liL2nGJnLwZpfcS4HZC30+0FGztsP9Fklv5LKB5bIlE3WJ4xL/MQdRRGvzJMqoS
7yVmpWfB/to6wJ7tYqVpVjJK8RxRfcMTqh4Ky9SH5YNc0ltqBau9n393tXOHeK/F
wvPuSVMSgyOpngL3TqlKqYjcIBSHbnIj7BP5WxGCSo2SP8gunBkM5faF1fRWyLUd
zDWr7Yqg+dF7pcePR8o5T90Xw9p7/AsifNmzduasRNjYZhwi4K+uGZ4tNHC5gGUY
NlswmchpWnEIIpmOlEZh5LviQDFQvHKnL/5Kk7hxIbgB6VJIf9zyrwJScKwW7Iea
/bvagXRr/jiJ6vtTfB6llCbnJ6FNBjtKPruE1tL4IEm6VuovJoaDE716JHC3d8mX
p7SGG/Sx+5ESa8NrknpGSAAQ09riQqpW8KRxMJN+61xmg5uZeioEGDQIxjWeCD6H
DwESwhgUgF+SRkNtU+UXSFR68RilJ4Z9I+M9a9yiOxpKY7aVUJMRJsaEQP3hoxfz
B9RiX2v57lDF6QHG+14bzU0TR4HxKRUxOBNQKC2rx94oDklsXfIpFEgcBnCJ2HDu
N4lw4EM/cDuAUiC/NdLgvKqWMsY27c5CXcqXa8yjqgXUyiuSRufGNgwXzw45C0+V
LRCLLGBujgBvS3lIlJC2MasckWejoiemMZBbIIwogWWkF3IsTob7eclse4yB1FRI
AzZwTtVPkwzltW7DjRcDo3RYfcdRHRAs9fZdo8/df2NMfZknHsF+1/J+1PcmCHte
8bgJzwrE20Q4IGMl00wNc/szRY3fff2nlXVl9RrOcOr3VgX3WW9fWC0aOhZ/RhdZ
5+nqTuUyjpAUPBZ9kG4d4TrPNDNYJP8UQhtagfpRcfLm7b/2w8YDAIt0nOjh5JBb
ssBVp44n6n8bLpguwNWzlh8h5FISJEjaLjXg7YyNH1GzxXNndxq4Oj1AZRSoVdQe
GGOmuRg3FY9Qhpqy4q+uxZMygca7JOGirk5ju54Knzn2ZdY+i0XOgCcaSX81om/9
0S8yOUaZcTkCiuI3cwtdMWO/2BlBO2pLBxtZpbUBPeJbR1H9L9dGE1Sn5wmYvUgv
8P9idswXVMLlqWWr1szUfQWPDve05+1LbTSqLO9a0JZpMDCudyvIqGnPUOh9esCp
gRCNHhf6xKYuY1+BtI9P5BuIKh9ih9Tdc6G/jpNRN8eB2Ue0dx1YXGaY+2kOVUNu
ZYJVE4pqPPGGDNVDMkWL2sQJv0h8GPEKWUa8MVxl29IEO9EeS1hf52KkLrZYTPEQ
SgSR12/2JTqRVD6rt04PHNPerbnX2O2ktE92uGt/wRmb4O+1MrymcIb5zisDGm41
zBef7fzTdRrKDpkzy19p+6UeeIea1xKF0qLl3/8wmxn6gmg7LeqxX+viWxGp3TRP
q8N6Sfxj5sXdrrumiWYk+2mva1MDyG7JEKzd/7Of60U6f5mXbK5U1FReioxahuK/
W2VKEdoDF7Ldu86SJdjyCzuf9dBtPWoOZz4i+pLHsJr3W7nxTuAJg0C6QA7wyEFq
k1egtlpdC6ConvHWKTF4Mt7QtiWSuUdPmTwenumGrbjO3Q//4p/hSLz3/9bpFH/2
RNCuVoy7V3lUeh6C9HGDFYIemOH3PzZo/zXQmyrrsIr54423kzJstWWum27bDhE/
Angin6CnnQv3gZ/oxNqfiJ0u+V4JbD/mn3kZgb2T9nAKvo+9I3y2wDspNi85SGzd
bYGHRUlQ6Loix9fWrMHPdcs0FCx5vyW9/kzrmfboUydOdX2UQbpGxhbIKpUtGRdy
5nkkq4RhxpJXn79q9fXOWNU4gWz3vUAYbc1wVlVYJ5BIbyBGbQKyoqEknP93BcwN
bKYKm512pOXNeJfEmqqEX9KtNnOB0oXHR3hJrXMbrQKgSEXme7TYarm2+beozPzA
Gf8sT3EPVrWTwD0Uo7/2pc4o2FpFvIjw28Rn6WpV5Jy5NsIvXXBcZncduxbXCtwU
djxhahshZJPlmHgV+8+0hZ+Wz3oeID/4YGTn2LfhUXbu9Vu6+4Ri0xQQ2nFCsniE
A83DyVoFaZEDYQ59Vz0DFupg8G9pFa4nDnidu0pRHd+gYkrOHTU65vTHon3QDdw0
9HmSZTU180ag0aWvDuitSAFfXfP3P+ca8MDl2pydDb04s4pT+8RPugzujSNXytmh
IkB50aG9WoYxgjw+9e29cVdt8qphfLd5vt9o380gnWJe/7S+zZPo7wfRscSZ1mdm
Qf980kpMFtfIUPj4QS0Cs0mPDmMySV1Ps9lhL/UGOBoiqcHjBIsIXwG1hn3dVqHT
g68Z5DnbT4EQZpRvWvKJVEtCfTIiqNoG4zapjveEfhlBRvWIhYo6wI4V83/o3i+Q
UshCVXwqyw6kXkRARFckPAvSzLcK39Cwfpzt6AYI2iUzM7Ury+Oq3YPsxzTMQCgK
Zqqr4LiOD+zy5U/jjxrBuqQ8bki1DQ3Hz8Aa5A9+TnkCGyGx3jN3qYHqo7HLJhCD
mfQ9xgye7fzR69R+FR+2Lxlx/sjvb2B9qqg7VYA46CqSYWgn+PhMMcdstOk4yQdH
ItPgPtGjNVE1oKX/nm6vpeU5pkKXt0UTZ/zw4jsSLF/cFYpOKtvQ+ULlW3kx2Zo6
mar6vQFGorD93nQ5wn7I2N7jF705LJQoRizbcmJvv2P5hCwcIY0Fk3i0gEyg0qHA
jmej34DnQ0Ep+/qyNMGMzS3XbBXlMrZsWs+NY0YHOeCC3OpVgsHS4mZb2XIDSaAB
/uiNwBAV2328L1bzt3hX2zUD4iKMob6eWgSiuNHNQN2a++o9NgYrpFX0ItxEWl4r
hx0aIajo/2f6DtNbtU8kZQcbbjDJn7YaYrUY2/8ugeknyB6nJuVGckTJfDiujCrl
vI1jU2GLuGKaB82vg+iFDh7XO3lkxvinbPirtAQL3VZbyCs72Tq7XBNLLVPB7XWi
MvWN1NsU2ZIqtbA21QI1O94ghRLtCmODqRNnDFwb1bYYpXxjtDY+wbmD2hMmQFgx
rmndA85m83dJmau/kNP0dhdCs9zc8qhszJnrisNa6DY6c/PdNPf8LnRgU5fIxxns
sPzwik37V/wQhl8RoAHk28UnSmuhik0K4y3VRDtlQFupwtfsf8et6Jio9EomLzeW
d1THHh8wffV/7FmGcA4ScTjGcgpuPNPsQCJvE5RytFr+nDgrffFQ64h53YaCPOdz
g7ckrGxSJFDrNXgRbe+eSIR6tgJI0tpuJD/Rdncce86Lz4lKGVgcKE7eTaKfDdol
QIuSCWTZH0M/qVzK2ZXNE2aCbwLBKZ+By14OFWIKZ+oA/jn+/k5GP5n7yf0EkMtD
qUNtCylo/n83wOSsw2nm2aSWRhHx+V+eemT2Jq6Dr6syjWAXfcFDx0XYznhoVQ0r
zFNOjn8jT06u3jecWhjf+HP7TTGTSOVpJOeezAqkF8G8sOsK/RX28MifF+hpmuDR
ougxGWM3XWYr0gzOLKjheA2KsJSpMw2RoBBWf7nGUUsey3UQ138BFojqOjbEj3bE
mhKIG3xwC7QldLVUMkuwvaE1Rpq1dQ9ia2Gf6QhNPdO7Wwdktaox3CsiSLNA2gx6
DnftimUMSBPANQKZclX2nrAfwqVr2kleB4HfRbJ5InnvpJoU1fguylVWIZEpDzdC
xXJ0pSGca8EeH1iMunlXsvjoVJanPv0k0Y+El4mqbHN+o3h6GTJMKep1eNyJ8Q2A
VBc39oCGuE5ICX5NKfa4W8aqB9Lv/HlTgLoJ8IxveerIf8JsCulUTWBP5JkHQfe9
d2FwaCAPa4Z/e5o0FSE1ZcZyilTejrIOW6R2w8IBSCFnPxP3a3Z4onF/ow/WuS9H
puaokjOcHQ4TQoO7KJJrrt7CSVEhP0s/eHppuNsRHTYYSs5yuwFE/qtqSQlfG3mC
cT+4CVIu09mGHrFcL5pqXgM/3pW0GQ7RUdM4QhYjc13AG+ehhRrPynqFz1GYhhhX
IdetUnzkvrU/+O79fMpvCYC12tlr35ltdhxkh6D59VfIbtSRvcMdoGe+D0b4IMDn
+uz9GZ6CV1MQDEpgwdReQJ4lToC9IQIRNBIIk5A6CKZDTh4+4urGlZxbOlkbzQoU
snu2JrC2EVpKJi7LSpy0NEV9EJ/aj7MHGH7yGrmWXTw4eFBR7pAXCqpH9bdX52eG
UliVdWmCrAMgRwV/RaMZAi4o597L4wgo9SBYVW9bUgY8jHsnH/2ROJTMvfpkaKAe
J1xS5vBac8+vd1F/4t1VL2GQhCYXqrNDRx3C0Vw40pzQFAdHStWhkoO+j714EJeN
8FJMZJLbK1rREQkCVCLn9ANPnPzQdm5LKt6sn9R7+h4KyinBlUBJgKciRIwkWdMz
7jS5n/whrR+lPXCQEv973xAR24eS/K2+1oiW5zCnHBLfgpZJZ0x+g8JbgXfv5OsW
6IJf8DBx2Sdpb1U0+rnqGCrRSH7tSwXaU4tf1kzE5lSftaxfFYNOxzOC6AFbZeUI
tkbxKghw1bvaGpYfDp1VIaMpSO9TJo45yMelB2z/pOqN5XIlrnC/zyTq2nhzPUBb
VSxfna1Gs/cvacTZarxlCt8eBu/dhhrX3V3dUSWIbDmqiaSO/qoQIDHT3AAPoJ9W
smbFAhoVZcfb+KrqDoqixFqqrgg9coGni6nFaLi37DmPIN3LGtqNH74TxuUBLqNi
1hCADEYmi32PJirIKNoDpTrl7Z26lkajFSFvLfgR0+gcXdXq9RNZKdcCouZIR3y0
IbyPLPab5DRQJEaHEjdEscx+vkSL4ff3xZqcn5rSG7DmXC1Eg1vowCfT6vyBg+Yy
bBnwz8oAYRs74b/WEXaIER3JGqXZCaZW9/2Yrld6xnZMbOCGyVZgeSMOfrdUaIgH
IlhO3pMPAQgkL2clbpBYdMl1lJTULyI2TJ8D8ZYxwKbbgdCP+HBc5vh0Ong3IKEz
/mRSq5Tsc5Txbfc+O497drusV87vPwqYdmBePhummyZTOvJZFymsmvPiJ0eVKfQ0
EhIkvutFJyBZtdU1awXif29JcUlfayAIPYBwexIvnG5hwJhC7lKW2OEM0DhYKqNT
fj/8Yh+sLNGguy592F7j2YKX1ttlXqJQ8VchuNHcWvNPaPYY3Z1yf/xqNnrz3jCY
caw+3Mc5cD6nsNH3/fJCX5o1k21+inqseOsTeIZJFXYFOxY1L0W6oI1QXWXCa9Gk
wvcpSyLkvV9QbHMne4c8Rw2PBw8q9Ko2nwexS5TBz9IRV6Q5CjOAuvdsawDJtMzz
lMq6lWB0/4SyJVfvd/9efuaeDoxHvUMUUxfDoIIaVifSPFDtGJZVehALJUMsXJ17
ygLV+S63ln9lrEFfWZ7w3vzEZORkf4FUTzr6yzZhZ2GhL7TnYhyii/yBKSoIV7Sv
VLIxhFtlNnFXhIb7f1jJhCAepXUzDlILECyJdLKU6Zr3pkx4c1/lAZ73UPhefG+b
guSZUPY510//1JHutM399/tQRxypWK+d48se1kahsqYH37KATt0UY4FojXJ8I7b0
hYnvhVJ8SdnxKcIjXqCHGK5GGJxtMtw+VIuoR9scNjRvZas8Bn2tsi/6RZyI67Wk
I+9JDMFeofKH3k04Q7UKehek8h0HYunG5kRF1Tl0DRLZLihxuJt7JD4kXZfoXy0J
rYoSj+ygWLEn7CdIK3llUd2aQqBOYIwGP+Fv5uQEsHItkXlhfeoYbyJM2ekohOey
uzcgx79ld+2jXG5gXBjG3v0EGe5lcHC4FwbvdwRUhheKxhFuEVtTcULKN5YciDa/
ToI7gIjV6Qz2fnfx/ZwOATR+PguvIkgzJoqFNWAJP2x6e/7XykniDkBtGPmoZygY
X6xOzJVmsk8OEOk/I8/l9i2FdFhWdkF2vpQ773IKa5TQRVktGJGH3Lp4SCi64BMW
SwBV4w53bdddqH7tIxVEheHCiOdwyL3qKKP8BQIxAfOjeuM22OHPhDBc4GZFTFUH
t2Jq7f0P2LGn+cLfa+5AVLTM7cpv2FT6Mw3IKAo6My5kw7f4UMCEsFCwFFvQ0pUD
4vu3Km7SD210LPHsmetURal11+lLM26BulhPpXDajJzS0y1hwFezDek0raBgTUzO
dxst15LUTkdJ3MuUfvWi3B716SPhbNxY5/0SiAJwlafypAZS8UCgGR9P7jl9o5UA
6QQW8ELs30zkKXPBYIFtYTovah0wbcZd8sgXe7hkKYGJx+d1lIRZNO5IpGwHNPoi
m5xK4tUea3uSiRUPsVxtfU3KvvtusC7lbMCJXb+Yl0UETAxOtx7l9LtPSnIZFnBm
wHK0uLbe031uXgUIpaiZrATUXFPOvUQCKJrlk2uhhwaHw3GhWDIsOHWuptuH6J37
jr+IuxXgWBFd4+FyPoFp+3TfM7rHI02cyE5+zWgZ7Zq8ubwQOImBWhVVrpMSHDW3
eXY7dnjzZU4zxJTdiw0PFEoNm+XV4nljjybptFb2Soj65MXmstvrNJ6zZGVVNV8H
aOqfk+npgyutuE6hJIIQP0hHIy6MQnKgzFrf/0Ozp2K5rd9WoYMpjcQlUmn2cIp1
vEj3fVdhdbatTRuzC5asAPKKITdY0lQvrTAn+PMSfwAIQ2EHoMKzf574Z+LfIKmT
PbYVpshh3IozC7UV5Znjd4bdKwvxXxeyRQgExo4qBTa+kSNw3805foxr9/IsD6Ga
H4l26QR2p/Bd+mtqcTdmDkicBbI2f+1epOL3U/zK/Kollu+FJ+W42i1QM1TMJv7h
eD7OQtthOvflMeqW5958wyk1E5o/sA82YK73M4vs9YlN9a8WtScgPSkh93exDVIe
Rhh3ZZSighB6+Se0iGkdhoWS67JifOpy6aHPS/C1o6Hqvgk7/5cdxf8+TBiSJMJS
xyl9jtbKSdmetaQH49jNSfRbiD1lNiN08i1P45ofo0OtKBFKj1UJWOwDMHKXQo00
h1q7o0E3Ed1MxOg8L4rcULubWFM475Q0AQ/Ro4WtEGDdG/KbQmTs3+AlTtruuEPm
IJk/XBeTW+zZbUVys1GT2dXx8H/aDKi4l4nN4vrTHiGZn0vSsLjQIYph6wkf6lyv
EDTSN1Xt4kwBaIxpY5i2+KxILRN25oWaF3/XC/o6xAV5h9UxGOVf9lfIM2c7Xq6y
eeklAo2H75spVYrNTueN2RSoYBbEAPdC/rxxx7hyYduu9uTCFy0X6rxOONuCtC5q
RdUekX87N+a5OrFFJWc0z5iKmHfnrhh66M+iPdqIRrGnThGDcctIzP039T9CZqFQ
2KNSUZ7bcPhJTX4BzK/+nsh3TCjafRK8G5OJHxvldOOevoABsiPG2egr4q6BEdor
3JXFAmjzOl056ZxrqqudgNxKcaixF/2vTAjERWjLSpxDy1K4tqTTmcPS7Y1DjB3O
XYaAw4AwSvxoaWJLKjdycNhbfdha8uCdkNcqMSYHnekXPcy0dQht5ByKCp4///SE
YMbW7h/6Y1Zhb5UHCAwj1JmeEmlzZZ3ZdPDmppv9PYS0Ly30HIRFtHMOGyekjmA+
0RxUliahnjd9pKMbGZRGt6Wy5E0PGMRtm4VYG5pgOvoMw22ajF79LyPl3xBc6T5M
3c/NLV6Yli9XPh+utkPY/3A71OMHXcdGpyqLbe/ZYJSttnIC41LioODNqSrsdb0P
yUbmjzzpk58AQ5MuPUeGbyyU2OUrm0lVcOCnpvC9+YEM5RtYC2nzFw99CwGaVDSL
2iFWdcOdtW5rTBt1la999Ozr1HQPDEAt1o4134oeCA+w+C/RNdlVX3arc8mUBIPv
QK/QP2rG9EPvlXn3IoWSlLoWJnyDl30RYd7teCPWVYTBCC3PPKun9beBTp7YZtwH
xnXtR8GPe0spMcohKkcw6GzLcm1iXg4gKSr2axKEz5q6of52VPU389VmZBp9rgRx
pS1AnVtE9FGNTvAYcPfnPZwrtrJzbZHp9NQUHkaEK8ZBa8bMCtvXTUBzFgVxWGr1
nYNebrTpyi+nduKhsfRZze52cb5bTcNnHR7GMyG97XYYRHleaHDyUjdo6ucd3bui
wT/oQn+DiB3SSiRd+N1GbCIzpKI+97GrnvpYrl+Nu+5ZgBI3VgW4fqw7elkwTf94
ZXuh9McFGFBmM+6rfajac02bbZE9GNfGdJx+1NCb/xr8+4uN4lYJncQpROqsc4Rx
KpiXtez62Owtj6VYM2w3W2R8IjX2hN6KFgAb9LJ0fqLKL+X4hoBqvGonWJr/3G5n
piwg01Am43KJOJ8l3kz94/K3iItZ3yH9cAJqrVaaZgDMR/fjHt8e6BzKaSFr9UJW
zURDEMCzU7CndpuUYlwIclEH4ffnHMUD0bb8V9pwRRkdrQNCWl6BAT55c41stylQ
KnfadJGOWs9E8quiw2OvSYI/52vSCTys+Gi6SykkZe53/TUiQAnUpbvIBqsEiHr3
APdGkzzxIhACBtHTblVkafR7xxD50Nmu9jxcNSaoIbb7Nj9kntUCuvq2LoHmQ5hK
OZzxBCXIq+pNou+aC0N2/dRT3pMjbD7d2p4yWfxf72S2ujwGePUrnRhA4ingHTOi
ogtbBUgtbbysc0gT1hXs2YJM6Do2j642KaU4ToxNlLbGvFD6EFqd1i6pCdM4zXn2
Mv18bbhYITkgKDC1orAbJzBKgy8l8sEbMX3UOnPq0sbob84zBq2Ic1KQP+R2FOKG
sWRXWXp4NxSarbkRYN/NvLTI14Ox73k4o4wuf4ac6n/yOvjBFEBNCLwVH6g8TYDF
GZYmlHoaFKTpkJfX/Z3d4INEwCU9BrfXttPotSd/AI1ZFq0hAssMO4inatpRNzib
SkTm8/YsGamduSBjl3QnW5Hn0P8A6Kk7L2Iy4ORYrU9DxbfstHZepDIDKImcqAjC
sragQsn19dFIsqhx6FpUo87GrLGfUT3oXmfvCRkrqFqKZjhSvIhcC7x0sBypLB4O
M51qnP27dp6P4yoKtku+pEGmxBCLtz1EnS8WM99f824MxZsAmUrNFo9CUIGV34ee
1i0Y9VYqENXNU8CzvBT3KE4pg0E8HWfzTjAib5VWk8AsnNBgsH+quUyrCOwFsvEO
78nuaB6V1bnhyDBlsXDdVsq1UCfuh/2vey42mOWXmOAWOFk/ooSnXwe2srGsCv6f
g6hsOz6Qy8XFbLTvw8Q0JUrwTiNE5ZKxNDUo7hqYNmURST7UKYQePgRqTloMG1s8
b1SmCWEsfTz6TXvZln6spzk4dzCG7eqADu95pJ2a3v+P9XmtbSB/zmhd7L5t2qxx
N1DtEFjgWc/k3qwDp1b9O3CaEQ73iz41vXu3206fgODHE+Q1hpcnk/Gi6XSz8xvV
Fbrv7dR+J3aDAzXt4ztqKUkl3uJMAlle9pG+Bk+WSkHEowXxLU0EBWnyZtfMQoJe
GymJYmpa6KYmG3mc0C8TNLAYD19Lxqw/Agdlu6e2v3Pno7uPloQlTW2bfTAsl44q
qjBMHWo4UfKbklDx+cxFQJ2+Va8UQOUwmQIOL0jJnOUNXpnYrZKKniwGD5UESmsH
z7GQGL82SBg8Ngeq/ydSNv5NAsshDmBWSSvIg/dRfx7qsHeA4KlSBgCpy7PFa+WC
CelI/YqNWHuoK+1BfNqeU4L8XERHUOVW/acMm+zyqYMy7r90xm52atJx/jG9f4fF
vTn+ME25BrFf8JBAD20M9/Hqg0edYzpT8NlmcDode08qD2r0UrzUMLtA/zzk5v0w
Fm7Y4CHUAxXWtViOKv/iS4V4jdtject6oSWfBObg6sWViqFx7CPcsbHHbtAwJCdI
/n2m5fg9P7rdpgVixiO8PGhQ1SSxp5cbdZV5kdY82Dvr118KGJS7PPXTvFGPqQfn
svf3f+wgEMKd9t+j9rKu4rXRuWK+2m30W7MptAfhWGb4gaC10pswJLCTKONmmGUs
YEs6F2aIYR7F+BBMCPUdnfkSHI/A1SAN8xfCdESAVKVhvpWEGGAoabl+hVcQIRPy
z8GSnkJK9jU3p6L0f97eOHS98sv7aPSUbXje/m9tp7MRVfCnwIVQDfA4QOUQmAKs
cZC1ybWYLDUrxv46osPjvy3Z2GSUMQtnB1giD+RHes2kCgFEaVgee3lU14+IUOK4
Ps+nofvZTDz/VIHMOR87LWKioF9KbadpYM6WPAboEQIdXjdioFRHRG+knk8qyuxe
oieFnre+gq0qfMD3AkzaVLa8JtlnyKPN+2kpQ1832rN0C3zHY2BW4VvMNlyFjNy2
ntx9J3tNXadWPZBLVrDfDKsSMTIQnVKE7+19aLUzdawarYwbxaW3O+B8EHBPtR38
vSO9bt3k+54dkIp5NNTaUt1hn8SI73u0EUzgmLbxuWn2X3RHv/aWAAW7CyWgx1Bv
tWQkRFABag2iGXTLDGT3O5DRV3pB/C3MMRoEXq4mctbO+ozp4rmuioH3Hj6b2aiU
TuU12fgCR4wF+/Cky2FptaCuoaclX34WFuBu8A/0qBsEykqXRblPrvJmAl9aCJRy
h+AjWEII8FryctqFiTTQswSreUa4HEV0XuNO9JNh6qgtdxvfT5GXTLFucDrD8doG
N4TTkPGyZpLKq2dHpnKEbW2CpfrQmBRAiSBZBMZ1KWcGhaBgjO10LzkHenydqx0c
oAgAgf1cBzZg1n+QCEk9ZQpaFDH/75C9pSekNZq+aOiEmcupNHuJFYRdS/6jcBxz
cSuC/99nq1yxPr6BPO51rlUXSPlZvw3jnHFscGEkcCCEAWmTNSfdiKaEjogcrVzW
cccJdhkzid5jPK3MErH6uytXtyN8Zqn0s4Q0vs041CN8Q4qgmK7SrgQ1cV1ckTA3
5CQuPDOJ0/Yxf1BucoOsjSp9tL+mJBR2NYzsxAkBrtYlEIHK3s7KHDXyElUPxtVl
ZllUCxm0xBYkptUJDIHrw/POiAJxpIkBg6MpD0QBNlXw4fjWokAeWBUEZ6Qh/F2q
ZbEAoB9D2oecM330MFpDfksyyyZOjixxwVUIEOH8Oca5wctTFIgCk9ETKd72/PU/
cYB5k3lNo7S4f9HdhdLPVqMnb45e4TR7+1FvPNok44KOSso0pGnNHJRHhrUGlQ9r
Tt1r24n891A5f3SsM1vVmhslfxPvuun9YAoEELd+8tt3uBZP6IcVbuGt88+Po5r1
GQ2SSrmwpI12zLjcipLNe5ytEf5EPwpbMvHMshG3y4Ea7S56DYNm4UEpk3Je0J55
SWMVVBOSbNQcWsAbIB+aiG1TgNbjEpVDkG+9VSrwXkndH66ryxklvBtpBAocZq4w
tK6UHQTlz8ms4rM52V47xlQ9G2aB68Pqn7yEGYdTzJ2Q9vKvr3Sa3SwmD4cJTu0t
/aWnDrZ1M2OrUt/yEK3rPeP3CocAJxQ6lXTID1CTWR71uxVVOYe7gKpf1AdD4nQn
+hcw0/Ii3IsJqWr0K+ojQjN1p2lNwQ4mkZ6Ksd4vmq7+6i2xk1v45D3lZ5is0kA3
fmbvbk+MtQ3RA3JcS7gscRicnJESz3c+jnp+n961L9E2nDhgf5VZ4gakcBXaQeg6
GDiI+Io0exGuJHmgVwzAHM0GQJ9kZyzGrZ5UwIMzHEcohDN6k1k6asy4xTjmjGQX
pC+kbygVUO7IJdBeH19I/4Ye6vMNeNdj7XXCNPgO3SPgk+idfGu+GqgjwzVcJjy/
8UbKnmjFJ+0FcFIH3WtfeBMYUD/+ZgEJgNwbEdNg3BLI3QeIjxJOOgVEakREnKQs
itfUBy+bsb/t1f6bWOyAAsjhoR9bfAEupMnAIRzyxHIt4X+XGpsIQIPxhFKLdyE8
lgWDuM6iCC1fwjxOlmpEiOi3sOPI5RXBvnAgyhcPnvAQitMKKJN8dtkx2tRXLmcM
lv//aGOZa6cXpUCpyFkh3Czj6xRuYBJA7yzhYU+lbU6Pfyd0WKn/VDTuDcBfadfr
5nV3teIgQN59e5o66+S6l2xBqhUAmKN0P4jPt9JmXsqlyGybNXB+PDY2WVHAZHaE
3TFk8pMq3P0cSvwxh/DT/VKYyvgmYjJxgpUFesahpaOnhvxGzt7O5WPoXYW16ynP
COJc8BjcMM/c9JWGH6wIoFkJUTWYE6f+vVz66neSvVtTMQiB6CfeHUl1OZ094BG0
bLyhTeWA8jWoPe4ICWNKrRQ4ax7SYsnWWKQP2StG0Gd+RlxlRrJAQ48LWPgEGokN
XCfL6XILpavx+e49BSTAOyUwVuV89xDNbP+OZsyrjsFU5xirbhfJ+2TvE9wvu/kD
wdSKEJYBC9jkV+0f67GbxpESgCPybPgBvHMDM3Sd9Ddc6FsBlC9S+rImd1UVmh53
AlUa/KR9Dl98JPZeXNiBYeMI8OG0HPn55M1RSKEwF2Syq4E543cBaD4Q8TujG4aZ
3hw440kRbuGYJzkpMoPg0RkdhEXdiSQbMFpWnxUKlCerEYnzy/jwBS6dsAGwXxAj
VQTXdYGZVU/Lg+uY72qPZaC2sf9rxsOHPv8jDyPFF/Mw0j1dfZBOcXUDYmYtdytg
DxHiZWAwuYyVu9b6gnQqpILEGWJ0p52dJ3xEulIZoGncFutFomLHTIOSucA2G/So
HZxWwr4jixkN5ShtrQ9p08fsv5al25AXfZnsCij81PjnqTKt96u16xFpNWOAEI59
BgOEOuEeJafN5+TlvNesUexHaxvU2oJtkEMOS0NzVZj9yKXOrjTOicX0A6X5I7Ci
dduCX5TF42Yj5vQM6NTY20kEeSQO/+zE9uTIGV0kd7xdcC+I6YsB1rJxHm746ItE
tZauPjkYC9UvcT5ANpSr6koYqwSCwAaDBkX9lp+QbJWq608eaNVY3X/8AhAk3c6Z
4yaAdLp01OZA/ekkNmFuuRGyWB8VYFM5LPSe4ODVQ4myS8zAnJfGWaONje7Y/OHR
nw7h06j5aVchnIjelkQEWzIL/0A1OMqLBiS5ewozFjnO38hgAhFjYgijalNGT8oH
zM9Yjia48KTs5tZOp2xaXPL64t3bMVmAenCoeco8CCMZonYy4GGHu8Dd0InVWeML
P17TlYhZlDZ07ustFuuPzBmLSHdUsJiI/KXqxaki3YBhh2vSHCD/15ALryo1R2wV
2VaTar/chyUmUk1JO0hEJpH8JwrpBNh+TR0YYYBtGhJ1wKJ+unSjiTe12btlcTjz
XhQvc5T39aaqAtTu0KBG6b30yn83OHkIyHdOBCsHIhpQNsWbvaCnyqc3HLQ7U4Ic
K/MIHAl2dNzkJ7L7n+LQ394AF8vZea7Eu0hLRdvZfLV0wg8Wv9U9YNzjRfCcIq8D
dtoa5k16t9WhkUtth4jVUSyr2Atmbi9VixZgNPx5vogs5a05NfaKqXCQHRcAY32x
YJvlcoQ5sq8jVJJbMy7l5rzDpFJTvkPVYQBu66YJzFkNZvp5jpsJF1o1TNITyzIy
rD9e+oLiFmAbuJIZYy339Hy+hPEmJflQImQkIGXhxP46khODOtEBrKM9/wM0YZIR
pI+whROVG4/trs+s5Qkwf3tzW8zrlk/nCux2ubBsyLDX4WjxLql+YyQ2eKGeToMa
s3t+/C1NXi0oc6KIHeQlEzgyrEYmk2hhlAFI2tcYy2WCwzQtj2HhpOAQA0Wfyp+k
98s8KOleI4J6rAsVZEhl3HAdhst/MuU5JhxFo2vKEQQ9o/EmjDeR+Kl88W3tmHKU
0j7W5YkNR8jrwFkxV3F7IQrJTnN80ADXiPHW7RD8gm3CeHNWe0zpm/m3SVneD4RR
myMbT6z7SMyHO1moZbkGn5P0Wjp7tCZZdCmvic9bcsLjxJO6EAyCI4DzEpZMwYnm
p+arwd84WKt0uZ150iockXid9wM0wejVXQWdxaJQDMU2o/hMH3odIKOBzB+4UO5y
8G9thBJY3db4rkVFQKDJTIxkkqCdgFDn6MjX6/W+2ovmK6q/PvI1F/WayPluqA8Q
G0Gh5uIg0A7FrNMhGYvFYhOAfTsVWapB39SwNuw5t3hYFsjG2+slQd33LdhPz2gE
qJEC95oF0HeqKyos+CgQM6LFDW5TvgEHW9trJRp/rFHomtANUPuFEYMf4jqCm6lb
PWRJwOCeRA0ibCjlkFc2GAzMjqqEyIvahewCGeHZM6r1Od+UbfM4GAmiNtleZBMw
6uiakqbmpb3cz1qJBFaUN2RkKYHjm8Q/T/XTN0PT0zuxtoObC8wbSWYvYnWmermb
h1+FJohce81uOf2nh8fVjMxg6L73IcDIKOzcA0fK3kKV2IYabXZ5+TgfnyufhiOQ
2PsIBidWPrS/h47SAr/x1ZVKQx46eqL5G+XqfJyEQAzDLr0QxZ6K/ngA/+z/txQ+
MwlLE1ggc670GLLSesMMjLIh0+4W5gIi+3HEAO81AdKpVwDmRIRSFj5G/jQiOZ8R
J9HpEdRvrFlD3H+THNCAoh1Yi4dVRmfj79sztaqBS2CQEW8L1BejOKEb9YSjlrut
XUZ5AxRyiQfJEhm+r8tJc29AXz6dP5J3C/9hR6jutSodelGLTOzGAuytEL20NujD
BHdApt6i1gSknWEjjpPEDXWVXAqTwDP/2l9wHDRiuSpN6/28gk64j31HGQwaW6z5
wancpVx5OfY66OlY4TuU8k3TccmFG42AJDKKYHBZOGtqa50aVMZ3nGeskp6zxeWE
ZFtDiKXJgaxPwiC5I7o26t2LuXHYX5G/Av2c816wcvDFp02MXt82f95k0GvAe3C1
yok2/RodHePYShvM94RjX0+OSIj+A8f1EE5Mnrf5Fp/98Fsb2F0GKnU/gU96+lFt
QxrX6FnStn2mspQnbJyyJmOLGPvT4rv7Wj8I2tLrfMX2zzMSBFcY5aQX1xgSbDAR
kn3+B1GPhlKxQfo4prbO5ItbJogPOqPvqlMDOpCIe0f9mq0CAqI9lCxumXkxD/yb
Dpkll6KXYypY4vDcb83xexNoaI61wTeOuRRhgsBVaXDhvWYU8h6rhl/1FnA8m/ek
YTXcQP7T4vhC50sUS7psgwo973mru/OnGQav3L2U50UZeGKWEZIbg+W9k3PL5w8Z
fkdK5qiforO+571lhh7+lTM/n3QIapoJUabLSPkfwEZ8t9rXoiUdTGn4Cjn1kHQY
kEk1Ss/GOkPFRoqh5l37NpxQ6xwMWGRTDCmq6cTQnjVbQOMljYjwnHmL7E7gpI4S
qdH27bnGFP5s26hm+kahyHUFk5I77kXcD3CqMjsfu4ZuQnuO1NpITwvnFHG8MRYY
aM0seiu52KyvtnjULd99CV6iy2gt8vCtPa7i0WFyPbJ9DKTsleAvdHYD9Hgx3Iw5
jLRkrCQWXY8CfnZptoKKAZFYnRwh5DM4xq/SRMg+d/a8M1xgf1G9fJE8/h688LxJ
vFuMRe/N3NNwF8HbQ3HDU+w+EobqWxJdbfnj21HWntDzlVb0Y9ON0MlBF29BmyQu
CxfhYhUvB8YQLx3yTX/1TsmW+2LK2H7+rXv41scKiaJW1/4gj4lXoe567ZhF0uq6
15KpqCiOGUeDLi8bG5CI10NyL0UQA+bjnlT46h3Gd+H9kKoKNXaTGJdMjZWs7V2c
HZWjfmSdrfAI3pG9o9qBhjXZMko12Kw/PObCKFvGL1M0t9YiYxj/xYGpsw4XnH+y
ZlcwSMdgSUeUOaa8IKkp8U5+juWAiC54AXmVmettIotdiZwmg/D02h2fpcQ4e37H
hs9Lbr6j19XLVWDPhwyvJK/4U1rorakU2/LpLuBii5kPVhlzRoG1qf2EzKK66ZQG
S89QIAOamQLiG+AuPPnlf6QYBESPwugs0u6dnsIU2pWh79Ss3MqEqJLx+LNKG+f/
F+11pMYyivGWCJXrAU2c5A+41lhjuXkIhbiBG6G+DoCzZzp7jjDadm3JKl88gcda
A4Kl528eW9C2HNqQU0hGE6Fv5dC1exnTvQJzPuLGvNJPYgfsg6BisgCMpgtsxB9u
bpkYqhBtZg/igpaA0+CPhUSvWahV9J7m8+A1mNAaYuRcwujLlUFlPb1xph+S0wcD
BW9tENp2FixiZB7Y28j414CbhYCqiJaACRe1woy9nRLIBAq5cRN3kFNbwH0y4m2B
u3L0Dy7a930+uEXyOFKo/9FiCcO3z6BAVxxYzKUQ79HRn04GV8V1yFhVQQkfEfc5
lk4WFGmFMH97z74UirtVaaQBLSm5AY5jIW8x3cYd+0Z1G8y5UoyDo6esXZ66W6f6
s2b1GKPxvOP6mzj+eOZ3BUHDi76JxIADwETOzx6viwZKWWxUe2umZ2oaPhPfPTSQ
rYfXZqUX6rpRq2NgwWF+l9/aGaFZXg15nV9pXubL3uV50r0Xx2mIPJ/5+RZ32ySJ
Sd1d3N19ar6c7mxoPoi5qXvVDkr/IegP4AA+ntKpGiF46usUMvqMsPz/ZWmNjQN9
jfBdUUplXGEuyzGurkK804eG49p0YvtQ8/IurywOsisuzieSvDLkfRaBXQMMYm4o
mDptswLtCF75HyuWzFBES1VX/z3SISJtrVDvtk6gINLrwOUdBkMZs05O7lwZoIAU
sasyJgTStkz3N9XROVnQq9yhsF/WLi+844tVt9Wb89Zqg2noji7KdhzV3b6tIjf4
1i9nVjmLeYyP7yPJtG3YU195cAy1AotK4yhaZlmBWdYhb/qXy3HLoGGidnVLOw5L
CR8zhBbmfd8eoAKkuS1V2uuqRTzexDLlqucoVszWywISnoMjBTZUNqvDK/FXh3Kc
Ngf9585JpLe0K+uMtTnle68edA766MN1OuZCSpVcWbj3DnF3jyhRX22usfd1ztc6
YzXjl5nBEbHRsHj8/U2aI5vCRdhpM17L4jFKK0wtO7s0+H88hdCBMQXmSEb7eiXR
N/5IYcAW/B2gi5nfbqgKlU3f08EowNzvskX1fAjUqgMrZE6p99IpbsjSB5iiOVuh
ZmgPc1jcZukl12camNWjlOd/vyGWm2b9RNnHdjMmAU7z9KK44OnzoZxvfdFB//Fa
pyUx8esXyBmDI1ovNYsixXZG4DxqPDUHVjeOj74OYOfEg9BGiqGmfzymWZc6DoYH
ZGYe5r8CqPMkyz+Z2/DNKO8lmHj7t0GfgTTWgb0BRHrNzBn+KaZt0k8xzUXYIy+i
/p2+KsTW5I25M0H/h7u+GdiFAgcdEghNIOpHui24krs/wXaM0ay+3xW5XYHqmhQS
v215jdXV/A4Pi4s+g8NW9Y2JG1c2ESQpAjFqV8YpLCsaieOfxfKc0Md6bu5MRfc7
N1JhMceWl3h3db9Abk9X7e6/qsUgaDIgjospfSnJVbIwax/cQXkb2QlLuN5PJhjR
sdHxV2ctA+4iNdpcEF/alzVbzkhCs+QApOv295UVrlgX20Zq06qmmhpe1LJz4Qwj
4E/G4JfU3chDzi8OLplF+DkJc9A1BrWL3h+UXFRcq+xVHRLhsRxc+aV/RkbWkxse
KFNWOfTTetn7OiECxry1jddirXsnfflWT4usD3xs3rHKaKjq4f8afjXDGrGQ9z2/
YiOu4Fr6FoO7vhh/Zy7iZWTb/uRabsSrOQBPgJUxQswpn+ZZCMP3N6FiRz6oNVx4
cWbCiFPafU0tr/zuqjn18vqP3uNDW/Dm7K6VXJv0pTUEAJLMVGTqhor//VKmg6FR
KG9bUanq7PgkaPc9860xfSPSegt0YumAA+WlSxcVZThU576Pu/CoTyid9NRro0au
iCdDs02gDrsz+kVsXg6CidHfnTlsahdqT2qayHjXIQncxdC7tl7y1GCskRWe/3R8
iMn4w1VaeaQEkBwj//oQVVbN/TtQnMsjB4pTVeLSG7zvI6vTX5CbyUsrmmXrVUq9
lA9Ec86xG83XvOAytWyFLGJenmKvJXY3dqWc16sg4WdHHiWbGj/mYyBGg4nEJiJb
rqdIQgheBHjGGzpiMppGkcsoUYg9TPF/jwKguKDiTsh9e9oFcPbsai9Ewjza3CFF
6A7vQmc2/Y1JiYjz31C3wHiHQndDe6GD3O6vv0lqUa1moygKkHSXMEMMotTiNR2Y
6RcGRmR2pwTDjIn3D/5vOLFAbjz1Dg1YWqb3/iWZvkQ1kt9fG0l999lrgpWcm2tL
ayDJPzI7hvLBHvUmRXkt4V6DkH9E3pqelD4gY9R0Smz6TznlRzWf0O2lCnqBwZ5R
kMHRqGSeODtnwoqpvM8Du2XznG8MdwEEm/JIq6h4NCVUkYSpdNvHCfOMA4QWwzze
XfZjZxMXWvBKVveDeUTb3WTcF1HJpFT4Q2DXcN9T9TVmQzrQBamXRVF+j5EI3qFl
ImN3dgR9E5J3G3KyL8gZK8bX8S6cw51Aj4RrCXp+PQ8sgkp6hvCK+9OMOrVwEWhk
I2y6PYuNs/ht7w6MYsFlU3Ij/EkdpotwMIisz56Qtci/sYOLATDYC/LzTJ3JTAZL
VCCtrme7Oh+EeiYhfYbT9DenlU8dwNQnQTu03TQBopjo6Q4IPL3nUklULkVFo8AD
MNPruUxoE5kIU0KzHY2HzB16TDG/gwHhVaUo1w22ua4/VzQ2HCBRVWykClSVfktE
ZUC60FG5vuZ+VXUsssNcGk/JnMzJakbAVxq0GEZYLV/g74SCfgm9IOWgGUCjwR8x
v7Sg11thVFtYMzglnsiMro8u9rbbu8aM0mM83T+7Nb8GR3GD2aaeYQeIBwLHrdg/
wbw34BkRoz8diPIy7POUrLMub+aLX9KVL7YEw7PgJD7NT/9C9aAtITHgtzAHs718
idL6dlcvdsIyhfTF+G86HsDEi5qxdc8zs0AecJdkMpKyGD81MEmO9RTfDOcRTNDz
UGcCra1qwQ9767r4CZc7HUP1skTHK82qNT1EoalK9xMd+yVIwI9V9g4DOMdjhVIH
27VkY6E0/SxU2P9gCdnx/43u2YWrlNMZDJ8K+M7bQDM3hT651UwZwQ/vH5ZyQhbC
EYAhhN1gT08E2vIcHEBdMa18jXkNtceXxkOwxMVb4lUOxBxMwvC6opFfDX+tGdI8
Gj3nmpGJp9BdV3fMFDElIhAn6yJbYebrbyVM2KM6t0J01jd6WSyxuF8qgkcXog9G
Sd6hCpQPoJeJWTnbYDjH5OYSgPN63i7133eOYlkGvjE/6PVk9APap36nQ7G+wL76
AhgMoWEx+MMutKRqdfrXbYre1J51FoHS/iLVzuwz6w5uVkMzqnA3396BAOwSFAw8
S++Apr4RIn5LhVYsWXc/CpKa5XpFU8EDsKzQhW/5mQl7drrCXi4Zg+vZ6L8oJQhX
U0W8q78aiDVPHJaiyToIXzP24eBVrxTDGLYKQs8E8uDjkVIQvCjTbwKSPR7CcCLa
QmZ01v40oRNQ1sWEM3J7zk3XTmav/cqGZ36SQt3W8WafTk6sxJyHSnsLjMFmTpc/
FlBy3o5hKUKxCi5WJOUNGFuoIZ+R5VSdLMvH+5kjRiVOXBN2LiWUb/pmeBg9Ob6f
O4CbJ2GaL2XVHO3BBuhAJyvpWxdtnrDaEIFFQUYZR6FV6XMH9QitBpMMYHSDT+V7
hSxEVUssZX88iDjvEw7O5B59GGYckcTvi9qoM0yOa1t1TJg/UZIJLXGFCA0BA8n4
YJT7lqXuRDUr3Oi4rAtqhnQ/eJMu20+eeufjtDOR/MjToLhkDL1PNCFlbzb+qWe8
sC4oiJxidI45kk714JJ281mHuiS7fgsd6Ih99xVXiGTmHEIs3NvFxFc89Le+nyZ8
+3+ycF26trSqha4F9s/ZvavfJzTjU2XWzmv4R3Cq4wQ0FRwheBf5XOXhmcI11xS7
J9lMr+X7os83ri1uMkko2IgThzZaw39ZxOvrxfqhn8nLitsmrqtywgZ0dl4sW7MO
+EHnIe3r/rviQfnNAVyUaHWXlPOnobyQ/U9n6HrTfEmD1sYc8JXnWxI3u92kKbxU
VZ5cO3x/T/RByvUIcGCb3mvAKeO7ptTuoONS3gloOIrqq1vw9yy3eUwSboXj2zrp
4nn48BOaJn8tqgZNOMAa/STMQGPWmwHvMHFJIiWnjWIdSbqqERkG7o+ndAZH8qBX
A0/qKe0/4w8rLnhlJ41t90Golnc0mbeu2GNoAv7fiSkEz4kbwoOTv7DrWVvPJyTk
opTMqx+6piuegUWLuKwQzDPl8j7vATPqSYD6Bd0ZGGYo/JDyJNhAnFViUaS0VPeo
DZIwqecs4j5qGkliuRRpVr/R+fl7CM3A8FFMTbIvzIMTNVc+mebpHfgGuJrX3//3
XahDnml9/CU/LcNlcmjcV7n6SwhQvXJbIEfOT/FQ7c9IU9+oiTboUkNJoQejuYRO
OfrptQon/F64jmeHES2MjwtIJVQvmDmPRJ2D76n9UdDrY9sxOwAQr/bPPCW5Oudu
Apq++J5rIhw08/k+3q08XugOJbz/7x9WuEqymbXHrbBnVosCiNncNVGNhHAO+xT/
cdsMT6mTlERpe6L4ZOa9NHpBHQFbWclvy2UMJQRU4QeXCuKofmZ+60x25mJZ9ylq
W6HLxVQ4jfu/mppKSa+4vQBfrmVw2LLrh6bznNllQjcJbR/dyo57R7iHFHYhqTsF
4fSQf0OPN6CiilJtVpbsNRZRWHY5CuHWHt0/zyUizoCh6nFiQLNzXwNGWNosAKD6
HkIb35kCaeSz6bwiS/g/Z8KTvCcDJc7bnSecgCHi3ni+d02NjJydlaWefNCFIM+/
K83ypAhhblCJctQn6zGbI21sYHvHfrS1XpLNlpEU0tppSFnoZ54kXmAqCRURZkAp
J/zy3Gh1MtpAC0K549FOJH2qIcp2/y7iWTgP2s5u7UKESFVeHMLiVw7Z9qeAuqNw
diZp1BDENDl21P3R9Toxi55hAHOPXL84ZuSo9aL9YYea1dRU1w8ZXOFSaE6R9EUV
13vHJhYGAd//y6k9xDQTheXd3SkMxHmddcVNveUdKBUrYkePYcMAOdCBAaoTwZiV
yeJS5Y7ISLhqtYPRO6BQNKeRrXRIWc1tAruA1xB3mH1vEuM/+daAEDpXOvirZvPY
ju6PECQJBMR+pfGdzSm8KX5uBq5KR2l59pmgGrTnJ//b4yAQH2gqedFeY+7150kV
6k5Mk7/hnn4asEZ5aKLmM2cDWwJaCw2kYZmZR0ves65I+LPvfHtpkpCmhUgiJ4Ur
PvJdnebZiau0uVp6BVG/2huOuhjRqZI1c1Jg9Bb/DCqKVJNd13Du2DYtTD/AIFEK
jxqjq93J7BwUmzAVchD6jZtfi83wsPJ6ZuppAD5YyfW6KGHccZPeNf43f2H1jyjN
Q7JnFQHpmdHoJRI/460aoxrpy690nBkG+Iq9mKTtt+vPcPqD9RFy/r/mhvCwvhSc
lcGqm4GqDu6yXgoduG3QNmFYT1LB+FfDpdDEyzisVgafHEPYqG0IaDiqKiCJSRor
oy21FDgLa1nLIVduCHv+cFzjqvn7NOaLLQudeHyKMtVkvKyuIxvWa0Eg8THuH150
52H7Sn50TClZ17zvbHebuY8+cD3miJEUrrCX4NbcNZHFn7Dk4OnSUx3Y1v7yMopn
pwf2dyr6jgx9guUDnULW3Vl9p5s9U+5U3LbJcqfHF9PaVmh901TvYAYpSMdf7bB7
9ljF3zVkq05Yz3hqVq6sBYbaugseujRWWVpci3S/Xxbb6V4v/qkV2douJkvAxmfJ
L0oI+kLxkCAfxAU/UiuOFrSd7AUVxk6hOV54WrOA+pQ5h7YMY9eUgsfKyUscngA5
2Fc6CpwxXzWa7eP2x8hTo7QuDp9CpcGUJQaLVHGG/xWZTootGDtz15JK/HPL1l6Q
2pIqfD8m04G752+P4sDOswag5W5lsooOhOXeDGMXrVIs/++4RtCV9KwFkYSjrh4V
Q8vkxGsYieZstsOujFGWfnbnZlifQdapOgIkttI4+kOS8DC0bEXYfS6FSIqe29/r
2bZ6rJWEKlKFlvrEgIwWkN08Sq+pL91IawvFOm7YwYgIFEf90VLVVy1hLlp8PteC
TzRubtFrZZFDX2KcYYHGPqNF5E7t8HmOSuVfQYGGjcRdgPzcPq3AlFgHkYmctOWL
LotDgWtcbRC0th1Lcn5MUnYMeLG5S6blZaF49NZp9zQPOdJBdaRsrjxGW/D7BRSS
QtSJgAlSlJr9Szg9Ss0M6ryMhEGgYzRHTLDxK01IFDmfrhlxeSGGgz7olHcBtvKF
AEukXL7A5NzxugV48k22Hb9B1ENltnoIjjFq1YebbDZ0iMNosnziJmzn8GmKudss
g3DxnYtIUAZWyXmMZpBc5fdrh28nKqNhfge3ZhlFsyMnJK8Z495Tt/D4jsG7LBHm
18FJkbtygc0C2FdjX1EFT8QSUew/36DXgjsfB0otx9dxu67rbv9HcWoYuezA4tkd
OePBqMqS2dyCG2ygQMIYcMoZXGbf00HpklmXfMOUHVxYkcSMKEBBZTpj3gqgjyK3
QdNuRHbRy2OW/OxxryCKx3PImmn5H8XXcsQAgHdIkZfAZ2thz1xrbf9HY3ZjCs3Y
oJqsOW9UgO9o6dNgPwDOdzQGrk2IeZmJweKVexgAU5e37YqVAqYjFaSBLxdFDwwN
NH/ihyQ/n1P+SOGsU/E4ffh2rPS8zgt35WlHYnhpELOeRmJm0lFsgDQzLabWpp4U
TZCU5EgaojmKiBYxIkIT20KFSHraB12iHRyW2/Vs1s8jR/Jmd4MyjZAxhQym9M/i
a0D1VvZ/DjW6XuSVB02UZDsP+JuoHGpzCTw0yTo9i6ah9wIGvchZAUGYBj8iX3/p
ePa8oV6WgfJ2Gm7SD/iDw9nD3OTm4Vnkvw8jsnBAIth68F+IWsZ5ez2e+JyNN88M
skTGKbUVflUvO69Dc6TWAiuZsEL/mMYyid/XLkQUe8D+dJhCZI0Y3+CwxXOIRN3s
DjAgVkQe9F5dvEkImJC47OZKbg62eNvwzWAkN9Pv9FLpDDwph3hhZ9g4FMXOEf4i
m4wEwnqGlDCoQ08BVcuJVr+57dxBQnRwD1C9ZiqQ3I3Ox/MUMKMb7wp6wFHsouAz
yYCBuaGUBaZjDOlAv1Y1X0YFEuXJEBfy5q/zueN6qLBRypnkwJiSRzAh24DRgv2T
3sIKHurMmMAmYoa33Ex0Js1wPx1EClPAMx+/lytBY5rSOMQCNunvlzrskBhSN29x
tqhJaQPEuSygE5xPK8AWDMMf4XR4Uj9Z70vV7K6KUwz0xdINWlwuc8IiykAEe4dp
QPwlcACGCYOiTyX6bf/0ewUcq1dMsCuN0btyTMVJTwuddsETmwA4SeB56WKJbPOd
u2F+JwI2+rNdQ3rdyVYxsf+XjKQUDExcZz3u/fzVgIUj5BFBrsifVNvbKd7OFsfS
uDAQosBH1Z3bv18O1e8/sUXOpz5YqO0qXDCHsQEULR/WaUGBiUNgIjUEnwY7JR7O
8nwtEYkyneCP99Ew+qtL/nUGE61pqHg5y8v6IM6ccEq2Mo45FONVQO7SbjqP/2ha
QU3WPxkKQ+m7qbnTt1sePUtHhOzcGoHTKoNnq0oSMf0x+QZvKbLy2oI9VcT6Vllj
UBI+Ft8thEB4CCsSQi2RLgOQUrtRcvlUMLVrorb+w/heSCnAAoEKc5IIB+XbpnVI
auWy9WCFwRjW/Eeg7AV4DGr9CzUKzymuLlx4rlOfxybJPqYbsFE5EXWHtpe2KgMr
r2yc4N5fiJSUCXA3IwXa4mHSJrIKLkb43teRt+5iAKf+x9Yf/YbA0fJxzta8XQC+
nLgyYCyQXK17uUSaEUPUZcVYzhciNE5DJJl+Zs5m7b8ZVtZkngJ9G4SG9RRfL0nD
vc1fVe5H6faeM3/62cwrY6G6Y9qnMtLOen5dR6buzMvw/dxAztMldrMJ4hNRpPAh
EsNbNtcv3tyUdVedht9u8+0bDYx9ZS3ia0EHamqRhPwNXkbQ/5pSy5mShGTZwOBp
c2du4FrRqLMGHhPMvuazXhhcsR3XQ5m0IiInbtTDLpfrnnXKL57EUYgk3Tdx4u9M
HcUlpswUkAt1QZJme4+GIvbQBfj+aOFPHIP2KXv4PNlxU+Qlrp1edlnSmCY6T+Zt
QfV/vjqymrPZKpeuPp53Z7ZBS97+fFOH1Ruzehow7czw6E6To2V56ANpNLuMjqo7
s6QJa+7RqO5NHhwnEKOOrEZhzGFf6a0Q/Lxihjnz3omWqgFmCRJDmESCdfN6AJr2
GBaYd/d05EupWfArN/liH5aLA98c4AjCljjAQ+50NbdjpTfpxbobLEGEunS+qo0q
UdJljOmZv18dBSIpeTSu+ZK79tZ+wdxV4BuuMYgZW7bLngUam1XXySSa463f38Gy
tNhL5UGg2nR72gYLKjDaDtw9qGJfmmTVHH16XN0WBJoqbSjRRKeym4Y+VfoY/usU
aWTQI7K2dK1X4EfgUjfm3NEzHaet6UXdbmHW6r8Cw2I90G66iVw7F/TQoBJtyp47
5cDub9wgyz62QV8uNk/nQVatuqOgaCSBsqwRze2yw8hHpR9g/lsPwdvgspR6Kt98
NS3Tb61HmLp2/WLK7NNOOHOI7XxC05rntE58K9PXog6vGwTOm8wPoMAD+OTOmM6Q
n2PJd6fVXcHQDQ6C+XBx0KnVUEYZwWzHx0bsfjgjIV5Db77JtKnjESb6CTTN2spy
ZFvor6720x134JJwnQRbnxsxf8iGILLUOXoXg8CVUr5kXluZbHjUoQCXXGVOaFSa
0g3fhEBUHDf76N/UqKld2pl5WEqnAyAV2eZdRDfy3cs/AjRwbcBIG25HQhoe28XG
DCZrV68MxcVtyRvJt90C3aN+L5murGpidTs3z8EQg1Ubr2UcJ/aVs4DWM5vB8nVR
4vGiffyZvGbzaFCo8pNBJJ258+QQL9VKfEkwQ54isIUj3cAT4IjaXf8fth/3Lue6
ZWrGNiNRlTXSXiLnvebRE+oFJRqu2AHlS3W3FRy9onEqtpm7fyT7aPpGTvJ5hSWT
JTWQTJWbuEbR94M5eMpVP2I1DoVKnBuMck1fLGVJIsD7DoIvYNLRchXdDigeGrup
/QWWhIle3eHLB0OfO4JzNzBS2TT5WcNv6W+eLMhjpMDElaGe4Muau6GPelNTx0oD
AV28ueVHxdTE3hX91wAv6dk6Vb0Pm+MvJP4fqh2XctfMQoyh4201zCPZqK4Btylm
9iAlWhZzYTHGKOQ6rS4L5ub5Ytzg1SlGLeKfNPlRZ7WEm0Zs9ugfflCI6kq/OmTX
6emOzgrVfh+1Np0l/u3cyCkfie6GbT/X8fkMezGiNpy2DBOiwULdLUOQYPqOCN8N
WY1Sxxu1rHwRq5C65rH5tPqIqzP+NY4NEkHXajjbeGR+ZcjbaiZ+/fEI05Hkk5gp
J9N2WVDxxnHbOv82AgfT9Xn7JyLrzDpV42EcxJGtuLOIBAkBgzs9qNDQIe+fQMIu
aCgXZ7iM2XJ44M7/dCYTJKIFcFQyzeNbVC4JSlIUPhvI9aLoMkxWC+E9J6TMO2GT
HyMZXwptt87j0wVc7fIKyGhSr+O6Im9ByhbIpnJc1FEwqgqUn/u39U79+/yq3UL2
G+6PLdLE72nQDdQ7UHUgowW99b4XVAn4abOlWqOhju5gM35ii0cP2frVgBQ8awBT
+69mrQPrruJ7Nc7WeE9mAd4S+aDlbwjXDamYnUOXq0xVjOdg8PYZEZpUkXCjQ2BQ
6ogfwHreNrJQuNxCoH5tW8kZfhvUzkzRYdm6WUwYHA9w93EY9u3y4SXzXD42feLl
sJOdBYnm7Mm2Bz3j0FavjvU/+WWRvj+9V4qivR6Ix2wg0Rd8tqk9iZW5tB/ORkoL
hNEMVXL7X2fkdZbuPVrQgXaMS+oeEQMcIfaskUs8czSeYwPvX2oAhLBay1wAlPlM
3oKFNjtK1Se5kFa56WtP1yFYodn4dkTf/cTJnESqMmxu0FX7NBGR/BlMyO7q17pk
EchkrNcVWfSzamX6yG8RoTXVhg7TA8YcHkqM/d0B+It1qfC42e7IjlrRax+0QDza
saYo/arsR2ag2jC0l0rltZDzYqzLkfQcXbCfP9HkOvPxhpsde8CnmOuSV6HJizqJ
hLKe/3TVb5kMMhIflngH/TrizzqMHrc8rzcD2jBpakXO9oMSKiBQS5FI65Rl1X5/
+Gd1to/oH0dneLR+RvEZw0hM03/7QgvjBbA5PjrgMSinJgodZvDWagMHkH3V0Nib
SdMOXqmfFxukp+cLJqYFLYwsBYWqXndthMCLNeUG2nZgRzPfVbDp0SBnKzKczXZg
aMULTcEo56ZcmqDijdP3OEusorPsn0PTyDxtCcetn8Sr1COob/kihYVxryJsn+YT
91pnyeXFm9TnHYONVYKR6nw7rZdpx8EiZYpW/n65okYaEVWu6yvwG4tnsHSC6kE0
Bd9hoXm3M9u4Q7uQwuD89d2FPrfEb5+vfOjH4oZHy4gv5QlU7pnDCzykE9nOaR33
LbivWDU2tVP9k4ZHJZwLMkIT7EbaFlaisoKFoGGBO99W7Jl89e+dvvrn9g3VpAhe
DB/Ad/gW+Rxt9EkqUH68lVo+iOcTIrIx3jNpeTMZtOx3Cf/BHULT1l1QjTfL3Qw9
vXsZh4AVqr+l2RdM2aC/Ao+YESeEoGy2w9kwNHjmavaBP7SSp7f4hEsA+7YwdUYU
N5zDZ5r7vdMGTPDl2Pkex9s7H0N19ZYKnZLhs0IEDeqLjrKm4AAKj6mtPWpyhitC
12UgPCAxxeHOVBFXPHFM01cB66DYv+Z8hxaa4toSRDm+LSfYPrjinLhAfO6NASS8
e/ala8KaIrOOeg041uptRM3TnW21fTFxPfQS11pLOvkR/owD3Zi9q+w8mp5sMq6f
XDK5N/GWXQiK5aIFgI3dBZVxzyxEPwZmZAF8DMHYp96MRalxJJtD16OywU8bHHgO
oezABbQPijgWV/fbA8SOaAs7jz5NNN+gwol2XcAd7C2yDpMTLmvMf3xMJxE+qwZc
0m5lYDuS0zJ95NaSVLffLARI2U3vTbZh+hB28+5D/KyTXf8W+ACthQEA7sqO8eR0
3NcYxpG43c3nGQ7L7lElAdJfwnbcok0RYG2woaKJX8T0odSLzSm7ZgCdJ7cRODXA
7ithMcd0wH0SXSkjovqUnz5LbRo/TBZ0w354LIPPrNmC44aDxTLEoGEUJZcnqm9e
iGIeVzryOuoqnkqQNVB09W1ynDie7HxhrZCChpyyRVycvSN1jMPYfQdLDJgLRbg7
39qjVOXbH2QbVkGWu8FwyU97wgZdEOKJ6JK+lGKwDAG5V/yBFQNbX2sP27YW9o9p
OxGW3DkwnIzMDroyD3NH+cYetOWOoxrErE2fEx+Jsj3/1u2b+DTX34GkrrREUwrK
FUTwEqmDY+Dg6EAJs0iF9qYRg3fZT3mC+af0Am6dU4WC/liXVK/bOpA2Ths095MI
2jfKxY8r83oAw3e8i3VAJysTJrmRRJ+ymfoz8yhwtqpBteAiKoRtH/m4G8OuAmvk
D07xqOysyt3wotF1Rnpfxsr7ySAzoSJifhH2u8Rbiwh/fRtSMjXuNlgmP7a0JmP3
7EYz8/W/vuExTmi3FblLwF6S/NS6+QnB80Hr4fRbNlUUV/Acvek5QhUMkkmdpeZJ
W+ViJSzx298quF9yWu1NAdzUYmuinJIjwzuG2qWzdPSA6NfA7MeEl99dFZE3+bPQ
I5NLdFMxyHdCoyg9RLqdGiwIiTlBfTv3M0E93jwAZZGGbWmczogPNOnvlUTg9O0P
zDZdrazz9adCGH5ajoWvKbj++SV960MQ15EI8YbMVaMV3dNLSp5dG7R8m3De3j2l
hzMN+EMVfqrWU7cQgPxH26tbCO50LAXaWZ3q7tpNwFrp0Omvie6UKvvR4MRSSanV
v+DWdOwC0D54/JXuGP3klCZ/tqmyij0eDH8plDbmnZQRV4Xr8Jj41s1NsX46L9gh
OTkxyKsif02N3q+S/htEZ2R/2+Ncy0Ao16vD9A0pNAyS1/FaffUjTSmw86rqbiHW
w201V6iXU8t5kdBvwhn1oC+p6vdQy9kyJj+kB0v2YMIlIXICy87UIcnErp8SVo8b
fnx0YXAMgLOVLGmlnf2tmJOSY01vLE9phLOgn+v4+B98sJuF85ZuMk1CJNN0IISw
FgvhxbEDYulMZqOGZMXul6/xNaO47nXuZe2kfHwNQNxitvUC7u1gHPvVwclWIB1G
W/rty0JRWltL6me+iqrbfHCqVV/R+j3xgAXjD0zw2yUnZ1WpM8LA3jAyhul1fTWF
MMrVWp6PLPG72xD21a4VCg0vNVesHBJLA88L2r7xZJC9PCoSKpQi0ZjHpI+rm9pU
EEiNUEkYQSlvJm0qpHaWuQ3gFXNM9bJSe24hlOEFGaOGqQiPvBYubZFQehakfvdf
/5/hF10MzrPshTUq5nZJVsc+Wq27XzSTQrZPzQnATVLTON5V5DbFKhv9lYsQ9ArA
ckwpp1r/n6NsMbFkpfpuphkVbT2EvhC/71ddK6syYX+rgx5Q2/Q6JktmMDhq8630
RNv/k4h6HMSkEZrVsEKBZrEVgWWx4qhS73Y80Vt/hOwPpx0KzXIOhKUKvGR1aH0B
KYWpRyuMJXi/Atl0VBkLC8ZwYh7G7o/TNRk+fCLXiSyDEBeWw1bIIjh5N6OBMQGs
+4r6kaBTfm7n342DZWkiIqRl6lP62RYrMfg5mJMyisZJxx4dzUPLLhgJ6US9cLC2
RbVJy7MXnFE0FcuGAMG7ueRBxjCVApJKXm6p/hRhcrk+UyuesbH1EKlfOVCFR5qW
BghTUntL3+zqhafwViX2BU3uBrK/OcgeqoACAukp7kXLYtO13Xo0bFz63NLHPRtX
xr3G5ySYJh72SdQ0Ldyh8DngWHls05dATOG3gwNG5ao0/RMSXiwIJGxALl4gzgEV
KbMnKKoe6tEX91FuHYZeiLlW8XwiMA3lchHqmz3jX0QL7ifaUD7Z25nHLz3x0XtO
hR1fMGBQ6xDKPb/MNWrDT9NhRdFHlbmG0friuG/3xmAF4onzgKtzBLxcsDQuuPed
+bUi8Bqcqj3zrA6LEgVVRnysTSpDSku8A0FVSXTIfNKvyM7lJmJrawQoPrX763ef
ahXDKbE3iimATK54eJlBiYYoTnVfimCQa9H8+oXmeFCjynkODY9G2qFyJQRVRZk4
pxLXRysStO1g1ur/cC8ksfRNtS152BODJAFqrH17j3i9gzB1SNCIM6x3aJelPJKi
1goLfZ1E3Vyr9JSA5SLw6PHjQIb//tQ1xAtib2Qrjwrpt8zLg5swW6EmaRgeXl2s
5Jra2/YvcTkzrA15CshBBLZ3kS8TwPAno+O8mwUSbQNIcY+veWu3NkuVITtnSGbE
ZdweC0HCV8xkpRcOWTKqBq+db9bhtKo2nkf+prpIMIXnpWyOmi1MIVE9Of46HtB/
Ir39I1UOkiqh2FKV0Hb9Hq1t+4iUxxIjMWncPf3bl2F26pCZsI4yJtP6seMYoX3L
8UNaF59QBHgDhog4gNNHz7oSRzJTxZKnjrWg+qkTVj1Tvs72YdYn1d4XjuGOz0Wd
uJCZh5u/d+bp3HUMfmxB/U3HtvsYJKvfWYq5x8SOpeSJUtIkm+f5wrqDL6OtzpG+
0neFJmHMXMVBrfP12xnQ1ggsKRLenWk7lY9L0fL8CD0D6Hwqx9LHSmKwg1bvAayW
jv+bldeVLD/PLtrCtOwmpwsZRX75bT2pulAiNuh8FtXS4j4ocNeSrjIpvguh1OSo
B7XjJT/jUiZgWX0egHbF4P4kYbhKRfG3N66PhOWD3KCDJjPauBFTJS+KD1A4KlUQ
wVpIrSvcH9+xIZqCt0z9fBsdcDHBmZkwuB5541U7jqoKl90NvDTE7snLYxJx7mcf
Kdbvgvij+OXhfJ0sq5lj12eB2Y2YgmRJgUACJM+V9Y9HQSLjv51w/u7Z2TkdoIRn
SAV2jc0grTg8VcoA7MrPYmSS+QC1gmY3dcdNRxeheUbSCdtFEG4b+OChd9f4IitP
ukuSwB21h+MNfBq9vZot1A4WYpQhgboSBk8H/3oAlImgXgtJi5FPpa6tWEEw+k/Q
gwieLy1J8uUpY1C7Ic0R7Jy3Qab3mOadHtjfkQLjlOsglX6tdG5dFQCzJEY8S8S7
mnOr+yIBhCzxAoc216kI09AQCJPDNjvRAtB6gpu2a/MNyyQWieTWmAGbIW4fi8Xx
uVd880TA1UOOmvt4nvV90DB/3tDqAN3q294RNi03/U1MCeP37FAmNg1Homz/fBl3
VRzz9Iv6vVJFOrSm8b9qi+wo3cTVgsyP+RwJtNoKtBiz2mJ2f4tZGAcMsnSw5Kwj
xLikk6X6+s1Rl23ljuauD3bVhPyDoM1qksMtJuUPJYHxZvc5eaq6qkeugCLAInRp
x51nyTISMf0jJ/vyjV38z+vnrPE5r81fNR9G4zus/0vMgqgMsrJgSefZduvYcsrA
EAoGI+MM2sUiPOsVTBXopoO5sALt/FXTkIKF4GgHNtcfkIIeUJflQ4qbW/cnJZHf
UOrxSGqHKxWFicX4QZ+4cp8zm6KrD4er+lQQNe866EINnztJpm/6gEVdRAHlsmpN
d+2p/w1v3TJbSedCia5mexllR5WHngDcaDFD8gWTfX5qZs2LVBoIRNRyc25sFR4e
8FWqsLEeZqX00usz4xdjXqK3aVih+lIUNNxhH+QxnPfj0XDs7qCRq/dmYiYGkEeO
ZRBD/2JXHEViFnfHX03wnJloYXz8cwIyjWb30TIKh8NrkupgvyF8fdClg7qAKLob
K1ffFOUTHfCeYaAcFZ97AlZEnk+Ij8jVqQoFiX4VQ8X2zQk0SkL771cW5GqIVjGY
5Soxl1m5hR3WESKcBWChv8ubFflyy3bj44jYlLP4OZzlwjBCFH7t39Kot8V5epuz
G9wNjzDeVLxbMrBjEO5hPer2hjPaeOvOiKArcBMJgae7wQ7uXqtmo5a0fvDNBAdj
JxQdJFI4CvhaM/buZPZ8KTQ/QtnTY5Cwfy/ED0B8//RjNqmgBbyVBLTrthfWjn4U
nNVkMSioku26YAKmSsZTQqRt83apAwe9IqILgpFgvM+INaLEQ1tENIXPwlrmKL9A
T1i8zXWG6DClOT6nz6fMom0TtfV8Q7a4P+JmVJ4XohRPmumHjAlQR8i8Qzkzhi+t
LBm3u1XXct7t/KrycqLoyXTV2KtPO6ZD7/zv4hh4/daENYSmQESrTdf9VVq+cUsm
ANdblqk0xALbE4t4uDCIQKJHYZIWHRc70+IhFKncWi1nWigCNp2bz1QCWh/aB4R4
nUB40mxRVUqb7mMZU4840SK0VYiEWWtJivsdQiXOdiPTpzdW2BGoUJZmkMmWsnon
2L/DksSALK4WjdGPmwV/wFegCE/AnLF0nCDPg9nNQ9/SZu8aYCr+ImvPkyMPIK0W
Y4nL6TapHTgmI3NG7kn9mPhu3NxOqTUgfm08XCejThO3EStRXza+wsB0enJXPE9W
Dg1J+taSx26X7Twnz4MiJfSSGI1s5NBURSl+q6EGDgR7j4ughvwEOlKCgA5PQYtA
snsXdUgGiEBjJcFKoyhIvI9g19vMXyGYu9Nvzp//nveSgSiKlcnFQTsBEjuGbUoq
lWYqF5rgSX/IggnvrII5Seex6tTgztqpkhbzoivsVDaR60BCBvJFz6BC34Vb6gvk
tefuHbyO+eDmkTrASsTbyJTCDwhw5KlPbXIc8hvypBm8BKuEim2se4H6p+nImcLK
nDPzE0gUw7jh4vZAPiQto6TYkQZUqay56i37uZ14bgqYMroY/qK2xjoP2NVkElc/
s1Vtz0nA7ukmRRCEkVXng4HHYyGT1PgXYo3a9WSmWkLoAZwFqy/NjsNeRWZGHZRq
38jWBYyOVodxyZSg4eANNsmZH5H+SQmsozIr/BUPUHWCR1uCLKs7VVeNVamQnIS1
vpo4Rg/aLll5AciuJiNT1C5OvwxIxNbhCzMgRH6huWZr71xZwBQwv2IwPHZ5zk//
5QibE8trB7RD6m0IJ/AdRPRC6581AGbCgakKB4Yft6sZW+VkjnnBpnbGUZmiHxaw
P+c6KxEl8Dc0gpVEt8aEwoC0/8nNta1x66gwiNPO6GjlB47WA5aNUYKdM5Y/p0fD
jzD8ET2VI5JfTQ7kOCWWBxYjmLY+2HmqihsWKjJb+6qJyn4/P9hq5dMhySpa85BU
URds36fSwLOMvyN8ycOX/TOHTDydppxk2WUNI8P0yUBZWvlP4mGA4Bv1MDeILscb
ZPDNGz1kcSYDGSZyIH9+mwOd//ZPv9GIRlQb200PI8aSb6nS6xZxwWnq1iW0od7T
FKAKPgSww9kOBOvKtZg05icKTFHgnDDbTxwuW+XYsP8dPVE7R5ZEOOoHFtC01Cku
PSze2mmBw8bxm5Tv+V6rQKA96m9FV8yVfAK81XEXktmj3CChLa4h14pQJs64A2ls
MD/Ko3B6AyFeZHWt+ibeGu+5hTVWzKpKm2Vvzbfzrk3alf4rVvDRXEcMrnq7mstK
YEFefW3tGnyxTlD0I1lSYbWT2PD8kY9JPbb/sqWXmKghXL9qj5UwYPplSvQieVEx
GVsS1Nk+pycA8WPkqPyaIs8dX291xFscWblC/FzYFtuUMC5/G+S7aWOWH7/QAzsX
+g+/h0y2wM9hx6HB/eiHgJJ4N1GZ37w0a9UjdnESGEXD5OjLk/LC2ZHGbRvKkeqh
3fqsYlP0sVjT00qXnIHDF7XD2uwPYqqpmU6oC7j9NYVpfWrLcoKzSvShIrulieGb
6vFOgLhSR4MlTyGFrHhNOr3xzVIY4U5ImJkasuVy/xL9GKlCRX0oLp3ihW5xI/9F
36SzwxlcYmZe52BgGimiFXQp2cZiQ4EGaXAEUAwIqq9Vhn+VmnMnlrEfkBzlj7P9
82A/xvK01rQqjW7BDBrbe7/9Tjan/X6OzFzXMDb9NaLc//JP5zxYz2WG6/oorJD3
RvEy48yWaQ00/4f8k1nRa9A8hgSLGRT0IdwHUz/i0lAg0HZbgyoM0yJuE7Q3MExc
atT/YP/zB9bVN+ebfzmW9iT3eAuRkvz27nRbmKT+8YQzSPO3qHHICqDPOFlANvL/
0sJd8uUIgJRov8GYzCvWT6Cu3qWO7lnFZldbK+70DnNzq84CF61MXQOZgv9XFU9x
stnG8eLnnGT96xXRJR38wobunZBRvYqZvJtW/+9E9rm5BU3AB8A9Gt3KsI5A75Sq
Irul6Pr6zYWh7Rdq4gzxFY7pnkFBR5P0P0BZREXI1ytiLLyghb5g4sNrj7wvr6xQ
1I/DMRC2kwZCDSQ0qCADwfDBSiUy0/qZ7rya7JYl92lgqhHcyXGZxv2MDcSMZHM2
LNddOa+JBR66pZnbWtjK2PzU+BxEfPRlhTzpTqaof787gwJNSgJpmTBODTegR2xf
4OXWZWUvq5d4NbThuNFWUygLMlbLuk5UgN8cHCvS8PdJUQrRaAadYS6MR5cz7cTx
stUNR6+Vh0pQKySMiaUNdRHZYK7boewuLcMXZHtZ7Yjn5bmMoOPFCY9LKYLqeWBN
iCZRBHx37Y2eT4xotwvf06PcHJxnKBalRrCCk1C5BwVxrikdlcCQGDKOer4Pz0JM
q5AjTkNJVQdXh010qz6UrnutXrW82hVpItELKx8bEBdovPgF16cD7DJKr2MZRnDF
Liebd3NXAz483GgWd5QT8NkpH49hBRVu0UzmUW18eNurc0seR9y3v/hyAX1V865x
hIiuTpAQZRko/9EcSJSzy60Zzp0t8SELDNdNZmbNZQ0UoTVQbULgTCoctuZm7c5V
0jDpOmu2Fq9EUL+JID2IUa9b6jMSFRdxfFWM6av6hhF0H5i79KnpqH8ws4pypl6d
oDqI6spfA2if/52Mgt5VE20XK8bKWddVk1ja52O7/3oxt47+RhBypbUugur6KP6E
ja7qv1e5/7JC2UqxyTTudh8HFlV9N1m28cvqIlDqMNUE/0a0l8LOG4EXUBwIuoS1
WTEUjx/YWextvemQ2/F3MUrLXAZfRAp/e8r8DjWpPYjZw8clawqeOfpJ3saAB9F8
j+noLSBHdvTKI8yv4tkFC+c25ehXC6qKkv0Du/1+YBjZPKShVeDFTLFIWJl6UfEK
k9Gi/HWcyXIWGLPuAYCXXqjoqedjBPZZY0TVxadFLOQENjreLiB/WvC3FlAAdk6G
6eJ/SU2JaY2a5ok1cAt/iSaKnBttFpLuW6ucSBfBmN4FAuxRkr0NNt17Gy0/VDzl
YRbez7ReFaDLuwCsTW8qUbiSOx5mXTZC1bfe1ZDgewy3AKdSVnZTgFFOfFaQsjOp
brENLjYszoql4HpGEiHasM/J+ktSIASfOB5ywZ7vky3l8dYjA2YBzmMyy5LkKdkI
+mw/sqetW3MHgXbOZgFmmSl6VUudDvGWdYLbZxeqNdAdyp4rrdQdh8a/vpnvqY0u
Y9Pz6tJ4c4JAhEOosfauho0DhwWiATog3maHNF6vH35v4NJB9442I7iTM8PiC2ad
MDc7UhaUHRIkMBXrwVu3w0o3wxiVUwCh7elUpRQpXJyybOQhUqb1vwkz/66rD3SD
3uDzTf1Edurzm3FNme+xq7MyrB8VEv8Ut08l9WvhDk5GqPQVoO4lcBjoAHzVfWfN
YImuA1upl3AQjmc9MX5hYLBH9TITuK5hmkci3K7F23B0DmWylCM23YeG2nPA5NuG
+WVlDxsid7729038bNJxsblfVQj0/xII3i0M24VZlytcBfz0PzkqoQOVorRTqy2Q
HjJmNS6dSSCd1eaLaUy5ffY95lVNnIbSIDlxIxD0tcLVYBMDzocuMfatGeTDF7jP
/128FKiiK1H5kuKM+0ycRvvzim8JIXnysStzeDRe1MPs+DqkA1a+3GNNMlGpRlpU
gGGal0Ln00vvk0iXnSGMYLMQZjpZEqua3uhfQiuj4DI5f5wy3sCP978s9nGay+Xx
IQ63U/xrlWxMsqRK7iC3G4SOLClOXgnDQjrGoAka4gRWe+hY3eNzpSrPOwjvi9W0
KLW+o57GtTsLF2zXnDHg/p/rBIvG37HDhz+ix3j9XKQ518QNuAIz5WFB1jfc7VWU
T9YtRrcNgGGGOGO8MRQgUHbknt9EvkqhrMtOE7KyrYWUHVLM6DsagIKmcYjL30sH
lMaeCXDhqjSiinM5sTO/eTnLCtJ/IpQbCmhMFoDM2TUO5yWNKNKMHzQML57vFGt5
MsZTU5ybYdvxsPinoaVbcP5gbe1n4c3bSX8DXmnFoCLvAq+Tho3Vv6uVFp+/fRUp
Yat9i4LOx9yo+P+2kh7Mym3U15KpVyK0LmqkOOvjRP2u9z8/Yuy3njDX2HWgbqK6
W9rfeQEaoMP2bNh3YLJm2lFdkZogLRBGA9Q9mbezkXogT8ohmcjMrcBSlwJM/kwn
LxjcF9uvZJkKBxOU7bhWtbWjx2653xYnA5i5m+mLDY7PVvtvUexCTCVX714Z7Rwa
2JGAqlo634c0WJqVNea07cXNmOcieaz8R8sC0iHxbjFiBlPOdQwDqCkowp5PDV7j
gGbYtdNKBNoyqbH1/klRACqKqK4y5RslNQiHnOzZlVjgpTUU5dR+Rp1dYxUukY7W
XnwhQ4Cysp+7jSaNtmIpByOeOQOpZHfa6I+StJ8UsP9Lnnc1aeqCChWfE7Z53x9y
uEL9ohAZfddSwS6tMQXkgTFuWJKjz9dXc7H0PeZ9Iv2T74lyd67yZkwV4OMNk8Lm
eevKs4e49PCOtMlZxsAfkIrFCq53nej1z6St1TRE+UOzxhKMZNj8nAzZnQrPFl4c
+KmnjUnH7JFhq00Kw1iOcB7MJhRKnjmT4Tm5XZD9rIi1Y2P51FYAhiPuqDYhhXDn
4eLywveDWtf2Eq6DlSogviG8WBiEKvJlvfVzYcEG/haCtJjUH8yFtuRsPil5cYyR
hkSTRVopp9Jb8kXOZkbG66miT69ZmEJQ1D7kWHipxEZHMAlfENep2BKjq5YzZ4p5
Nc0cUJVpqrsHJ37v8+oBwO+Fw0j21c/uehJdP2q0NkRQXMoYQPUGeTWbGRypLviZ
CsPe17rYVxXzfZwGuDAUwi5uv5Bzt1WT5JOnpzFXlemGuGGZnn+mbzb8i69oY2Bp
/msRz5oe+9TFkg2OGwORU0/Bg07xgJFpq5KQpvqD5LpUHvdiEQtICSmbdvsRgCVl
Bxm5Pteg/MSYu0y+xIxj3JqSSGUOHKAsH96AUO8dUHyERP/nD+dWjPQakKu6m7BV
vi1G6RQqOJw8Q5DUNxXl5hKX/cpl0hllRsG3QH8ZSURDyoF9Pgglhl3uC8U6MFFJ
z6HPcS3cD3zuf52VSrClkSbUPXvwaxAKazfEI0WoFOkmfPr4V1DumAW7f6Q55FPB
LJdmMDCVvX9y/Us1KWFAd3jF/4fM3eva362Qs9QBaAofpuDujo0eMGcCjQKd/AE5
la6XYbx7W196zIeSJZjdpTlZAIMSftepIaVOOkYB3FEwAKkl8nVj1Iq7RDCAn9wk
RWZ3VpcPgP0u10eDtfvgAQQXFbpUIIY4o1swsDAJ3yCaITm3O0p8ee1NT6buHmdg
G85GkQ8I/LSoz6D3b6wtlwUWpDFghdouv3nNda54WbVFUrO+IvRiQpPCezOL0IfW
wewG3vob5GrNTB9zL3PbQ4JcmcKxkTciQg9fM96yYtjFniRtTeIoIyNWF3CVdQ9W
+fwGhiCeQBFtL6ngCmPbxkWyZjPR/TPrBrlOiWEYdD4GIEM1if15IyzZYlAM9AwK
73nSyPrP5TC3VBqW8J6z7MfwI0vJJokeUwyJ8QpM8OKHvgFGSxgRyguzu0yJMZGH
OBe/Bd8FVlA8mzk75/zfyyAkhEArLgW0cMWEPc/DNjtluJl63me+LDEJPmghbQJr
cK5QcgVDgFf/QyfB63qQ0RNKUQgX9m0phx9oJ5EfFtFLsa44Qz2k8Oe2rQMQG8Aj
sB9rv3p+2e26TMNjBmeB4DxFO7mNgEvz9pL7k3Caj2PsQvx3gj4JXZu07Zfbp+AU
uSXmk3hjQkV5/zqDuLsheMnT02b688yqDU4WNbd1SzDwNCkhQMNZAXjafJOQIdZ3
S4xiTYTI1teVSX57XsCvoJHiEWPoxL6LCjrWGicpFSGzuditYO7PC+OllHFQpU5U
4YftzkxsLbYWrjWgwBMpXB7UQwIg3aITs/Z43GvVPd1HNz1sEllboHhFQmAoC7aG
fg5AoqjdL1MnSS1hZOnil+o5R+HKIAZmhhg1DQp7NzVsWs4UICU4JY32Lwd2A2wb
xWLAxYzcTrrym4bA7DP21Mp3uDGZdEOPORUG3Lg3r5vojPp/woB6LPaw0b3PxoGC
Ifn0cAR3/mjlevlZ0yNU0G8wVa4GDy0hDDtNmrMKO3bLv2U9W3X/Nf1bxhHRejnR
mOs6VV/bHy+wHM1aU73Y3RxJTTaJRGLbrqFCeN5iwTDtjPV34cpV34EWGuYwI46H
Lj5k+3VGGDYnNPdPulEdvMIrk1Uetft78wD/HMxqoZxhci66Hp+8TTqmm84nQlxa
zL3PRS/d9Tmb0b3XJR4qPTkzs3NXETrE1VpWi3PW7z+StJA1Dx0Kj/izThPNIg6/
tMEp7c7jQQOpad5ozA0CaF4icEHLMHjpzxuBmAVolabYjjqJQRBaXLwEZPTZJvpD
gdDabR3oiAr2wMyGpdYjfkwseXRjmBweQyHqKUJW+Fk57qVIoeJbUT4bfXvJ8+oZ
DLwJM4U/tSqgeqo21gxmELF926ekbVu3dvmyj8DF2PxjKFmlq7ij5X8p3qvb1bf4
NpKRFq09MiRUfcoL9dYGpRU633VRSps8j0lc2SV+2hSLS3bHTdklXs6Q/MAVMVk0
XhavNqmRlqcWAgDkGUfKmnIOnBsbr0nLQvIv3ExT5TeuVeRciXriLe+7GNr1v//C
Q0owepTH2i0R95eK4dTFO0ZkbJht+WaF56I1m0IXkMgksX7yzTkfvqWl/AHVWVdU
ZtqZ9kk2s94qIRsfGAsijMGq2Kq7Rm08oLXFGfH8zH5EhvQGMNOC7Qp82kFGXq2L
Qo+eoiYDNn+gszMW/guaz0sGV4P+ZWhweMTigyfMAsSOjlSJgggfX+OZ7tn/GIf2
ybv5qJPvPKm0vvYoVMVCJi6PzW/+PQV70SZG257KMexqKZIap2jDWbHTe5HBkZmw
VxYJdc6TXEeG32jVUpdOkbq4hl2cIPUI/rXTf3yhP/4DeiBw12+aFNzP/sojXzqn
EzZCfMEvFrjV1dpPhOMxIwar4FAtl5oe+YV8WYZrNF0zg5aVWTXCCTGLFE4VXIEK
22NcWqrkA/dauyTIr1WE5fDgj6ULBMNzHaSUCyi/tyyxFNNS20/KgtmZDPlHIhPO
iUPiOcZ1rI8HLvEu++dAm9LVu22zX63UW10czghzvuMot+Y7ZkxCwPKdC3yIYLiT
Sz+80wZxkmkwf0eixasTOjYA7bRvItlxsBokfeX9XU7LRyod8SL/liwlUNr34sfl
17ITsOt8TZ4b3bPsTXOc/JCgvd3Y3JWinrNsRRcn+TIrQ6r+7g+YJoz/bngoNByj
tjdEFNz2zlfM1W6UDs7gUIsDSX/iTYsG0F4Ig+etJNsPg3x0mQcrZ7Nfoi6eV8t7
0fFhPFXscXdMs6rH3BxS98qzlCW+6I0tUYfAm4Vk2uNnBMSI8EzhDXF5PNXBzITa
RrDAkt4OnWGsaJ1EEig2mu3c2ZK7LPtHyS5sCY5dDCkofcY2lE2XAE5tmKjeDak1
pIoHIzmDJh8Z+8gLk7LP9q9jlCWZ2dwEL7z8L4BHcQelGXAIudwU74X2WiYKDAQX
St4kyrZp4lJkr6gwftBDM6jbfBycQW2q+mPPOWMsZAYi74tYpb+2BBtq79XaXfiw
ZQ4+tlyQB+T5/glxmQVXl5CB2wJjRwxf8QTPPkMbZJIgibdWCDKuzQU8a4MB8YhI
KamMXkZ/It9nfkWZ3whcFhnE/mrBRV+HfTvobkmxbKv4T/O4k4IGdTM+xVcZYqHN
KaUeI2ZTy570XUxvqDNEa9JOkVhZ4Ss0d8c/G/IjiPHxSQsVFduVlr0M7ZS3bC67
H/Ty3ExjPBaCJeykqTO/TNLgcHVg0aIwXLREXPQ9tS7FUaaFVJDBann75EhFXX3q
4KBqo4Aa3f2cZ5NABBftsapDWlefc+/41FdIF9Ce4eKFRZXZj6kgyHxlPCnC8cxj
tpu6KdiYo5DKcPU6HC8DHG5ILThxfGOv3XWGtnPn6RDXXgiXlb0mDLPgPytwH5+j
n2NBZakdXO4aym8G9hClfjwUYjNvPcR1cXs/DoKnd98SfFSMwZdcY9wMj7vchFMJ
SriYEhZ41nlIiGRFjq95wRzTQGtOsOurCs2bfInUn6v4H3er6HnawejnZ++KqkVL
OPlpyUoE+Yf/B/Pjv+xWsidrzt1qSXQFLZTGieZcLQn9KtdECVZJzYvoGGLCL/au
AI6beEiWEVcIeiaERvl44vd7NXJJUv9I6ayUfYhYmJD1pwI56UpQWXzLeeihSOcS
Oh1nsKJDvDITWvkvsaR7WBbmc7iE2YcObIw30+e4AwuyrQkCTlRsT45VZKqM4sTV
+0L9F4rdXJ2AIp1o2H9f+2J345GJhBCLDwPkq1rrONIUoq2HdNAARM8upJ5G9vUq
URwlfP5BHKrmrLU2+mfukp6vH+CZXx8q1Dxg5KLn6mnd2YZRvdcr7WL+z3WPlqmp
1AT4+5DignQ5G/4AdTG4yhWDZplrlp9DEotp+0VzoTvTILM3v2w8bh7Juk8i/z4I
GJZ0WJhsOnEzJyl5o5byzPeSLz92U8EjuCiJ+dSh+vs1el3vEpL1d8ZuIkCgShgE
qmTe/DHGq0o3SiyWKPneN4Lsl/hNaSs3vqHRMJRUCaq7q8VHuzSSKrrJhTIhJOSU
uZBs4LCMzIrAkfT+K7tfDrRBeWaBteXCLjLC6RxAEf7efFFd+W1hzbdx729lvXzJ
FUb7RwAsAdTUBGc1clVOjlCZgIDNboVRuWYF7FG0Ps1BCRbPO/dufkfT37RlfGF7
1h42rLDVPlEau1aAJJZQKauzChq4OpTNjMttjQCyS0k2ohxhzknYyQOszOJykcZU
WkZrDFr+gAsvSkAZXb4gW085OYgxMbu98HPuxgxcNJBniPI2gXoifaj+Gq//IpiU
YoFeDVPduc9QTprtd6jxuhMl+wACJTUlfjgsReq1XGFsjGXE3k4W/vUdFM8op7vm
RUeZILlcJ4Q2hUiKRJ1MjWcdvGu8OsrjnOUMS71zwkwOkp7YWZhhA4a1dDcttpKH
evpjejXC+bBhID+l1HgPpxw/qtBOlOVhh7hxPXVdv1r22yVMuHiAxuHVu0HlJdyg
r4xthbLr4abu103BFZ8v7fY0c81HG3stuilzVHqaAIzI+MkfdvBKtz9YIJGvPso0
bCCIKo40/sQupyB+caAR6bD4yACD5drHdkTSeMkrnnpLdA/I6TB/b78YGT263+5C
43yDX90551T4V6QCxwxY6OH9TU/hHOsKWmzm8QGLT9iRtKl30jm+DZfbptI4k1mT
zNxy8qkjkdeWHYiOzzqwTteyOLqaVYxhT4Vv4KDSpaAjhMc2cA8Qj7xPQW+DqtcQ
qJmkt1ZtoHfA8B+TSLzbrpxkY2YInIJS5mXFmwuc2TcBCCp6awsrdMj3hUljyC34
n7fz5HW0FRxNzgnhZqgz8NcR+LYjKIrzoK+dL9Q7C2WWK/1yw/qHZdYGV0XH2Y3M
Vca+UXyig+bb+gyO0y4pnbAMCBEDgEu2w6rSXVYZb8k6vw/nbaAA6J0mBvCJ67pd
OhywI5cH33VJOdS6RLj58vLgz6OYI0FS6LqkYmhGm4y9veYREb43+UMmd1PdSZi/
Zw4+J16Tw5nn3ZAqMVSb6Ogo6UeUUvKF9NYqWkkmGUmD53/DAQ9q/IX07YtYKOV8
LgMvqj64dPb2B2eXtAYZ85Wwhtl/4VKb9H1o082DBjusJZC68Na8aal7yWiL8qpD
AIuU5iyrMqu0ql6HvijO2Wm7wxGsXnx2c60WjxTWNeWF9YtUzli//3jHG5MiaqVn
DXlhuxSXugmWVC/RMmG735s1dvyZKblBE/U+gaelw7Zv3/AERkO7voAMHAKYvDZ4
ACxnNTXmoDVFk6MVfS0ylePpthUO3YVJAnksCpOs0JUBnBv60/ASwfaNgA9WWQ6Z
/s4a5NZqCsjDqaLMKkMcuofZZqBZDoC7Pom4MmADdByOpH5fUTPI/F63tl9BgXop
8vyy9k1UKYva++H8B9/kKgqtrbIJn0AMeU19aavjOr9uG1hPXMmIVPSItUhxb6Qi
/Pet6ajr2znS7u5XLkBj/ETr17CG8xXU2bTMbDZPylwd5VPhjOPGseYj12i9UrFP
IgbvEbyh0Aq8sUZtUT625MF8SEZ//Q7B8P+nBSjLle1hIQtt+SvixlnN4JlmCU4o
uUWvFzFjtILhE8wQwkuY3eFzpMvCChNbzA/C/wLSQUkJ3S6T9g0WIW0TUQWGOmNd
PqGZ5tFxNbKUZhcYN2YKEc3kCpLDlvZ/4jBUJgWruiazQOtvaMI7NIQY5m4/D42o
DQ3OY4FaD9/rsBSTX5fGs7QRX8lRS68remnoXSBqFlVvAkY1k0xWCp5DeniCEtr2
sSaiyLPutlxO1DwyTBtJsRhCIBDSKgTrOL85I7rDZyk8c8JH+ZMaye9BN8pcK0Kf
9xD8SnduLMk85VibtnbLX3TJICVhfXnAy+YRINnn7BuoUvwGp8ZYCK2CMQrB1r7i
KFrNJbbp3EVGFXikvTYulniTf9RWXVth2nIxw1i0olHu7IiI89M5vNyfakO/1yvx
XyjkLwGwtLAEbAy0QjRH2wydStsGmEKbc0Lf6fDqhCTe00JRsd6JQx27Koym+e1t
DktsGW22pQQvxZ8EjLxS+9TqKQI7hCe4gPvKSFtc3LHtyifG4Y8aDOwGaX/uTZiY
mf1qsa7CkOXiwP0RoBxtAJnJ9wqDYAAK3D4+d3DHL042GCH1wWAQiyPiCq88+/KR
gFsPryV/oZQjwMX1sLxmKvRKTlA/fS1gJD7DJasM2m8ZCOM2j0Y+vzf2M7K224XJ
xNnVi96HaTOT2jGyfVKhCrcCuHD4mxHi0+DaTbbRwdKet3/8zruJyUJJpJDUrXov
t3Fy6yb8W6A/dinpEI89+fEth4fddlnqHzMlILorqqsUkn92X3F4INboybkWMiU0
9+12JTGrPVaqhGGn+JmfR2CmLiglZF7ySiWTQrHV3XOCBBV8hwQMnmvFAeNbGCQ7
anjXPu62w6CROK3Fw1LLbxZ0P6tAKMFnsKrsEC6glYJ9TjzCx4t82Yle4/2BeVXQ
faK/dDSp7HhcFLoPefxklrhKoktPdCVpTdYafFSjsctXUTrjRDY6ptSvLfHD8TlB
5akPU+7UhA5aC26eT2anrULRkpVGIzYzxd+2GmghayMYiOoC1y7FtsEdyDyxoW1o
c55ek71rBGtildfj3LXTYdE64CXXRtmH5D5qYHc1kpbkUaiF4ssHbLJMZ66EZQ8N
G95FhMx0OXZ3ZZqNWaGi8RVOMqRoFVd/7ejD1Jhx5WAQs2/Jigz7alicFim+Pp9z
KQnuvgx2m5B2F2eRfq+5/BLecOVv+Qkybo/P/6+HBTTAFFiX+3qOERbllJDCBHZr
2x+C0GS7O3IWFf7wcqdJiJ3FB7mJwaiHvy/jmThMg7vyn3KCKjU5IXD5guaaCIVd
mBMyxavUPPpM8YsAM5dOlTlcfiGpJZcgIcTG6o3e15ZT5oPQMqOq6XdTieLGbh7P
RBnpOK55LM7JRke9dolACyXVac7oX1iqtdNNkTG4OT/ss47yiy21RtLeE4Y7BSxL
Cw8nUDl6mrDZylYsoSkVVHBsiDTBfWi/L5jbqS1aOtlfheyr+LoWVagzE+C8Ow+U
eOftEHgHxLXBPBtzlquxrPQLpfOLQNwYkiu0ytVkrFHqzwq5Sb+xPcVuMF8MJgfp
Dt6vpFXTUhZ3loI+VWVA2CigwpVwWAiL8r2xSAYdmUkbLsFL5h5lW/JlCTdhCcXU
H79nEFc9qPT3NEe/TR7ympF/akAMNPN8YmoijaFzlMTLj1DCr1CWEUUmmlzS+cCW
eaqddLSEQr96yTCPXOmoDF1qfLkpkisan9znHlu5cmC9vSY3Whp35EP/3v6JTakR
6Js0UVRV4b+S0h6XrG/x49OWDtWCR7D3f03QjuMu4rOWS4vyzkKzMVeRLdM2DeDQ
RL2FyXyBp3uZGIa4ff9MjBNcKdrlqFhNUBskHpmn1d2wtvbhvt1dg9ybhp0VbH9Q
6sz46pr6gkbC7mb+lC7rB2MDg7v4KAf8AWNM46nD9t7JDxzJOX3IwrQuOfhc5K91
PCpEDGI9OVZCTAmzOdXLO84fe9UHoq8I243iBvwtc30D+01j4/2OF32RS+jtSNWz
ARGBtzsknOUvwZc8uPNl6kV9ZdF00+J05JhNghnyCCbXwZ13tjM92kDkuR4WAvAu
zkZh5M3SlaIZJ1D4ELKy4ks0/of81/dq4sWeMA7/YBBvzM87KqY9tL5IoDL9ExG9
5W3wka03GenT5nCutgynswlmtt+ND2oH+MBA7ih0uwoja8rMx7zmAV6IdpsTWLdT
TxExTGyDjFMslTgGlVXkqtX7teS3nh4Hpj2MSBmffk/x35GHoQRITA9huew7bNXu
149SWOiuljiiQBXBCbS7yKOPSYAYcLQOry7pDFYM62t+mdOv6BkE43dpmgUiIWRr
CNdm7mkoLrTDmYSa4NMWXq/dSnCb9BsVMzgOZV7pBwmhfs5+atUvLtqswBQL0ZfC
XQd8xiemBQAQHLvSZo9CIwhUnkk2/jxCO4pqiyp7ZyLtVtzxhZwoKxk/yIGatCNm
sFS9Fo3uG+o6WwXAIAOdKblI7uZBvKp3ZWfFV/Q5HEUnkgJveEc20QNZnRoRUuPR
fjg4sUgc2irZagWgC+q/uBLAcy2jcFBTfWs++7d9icD8yOzH60VijMvpSB2P9sXA
AQPmR0PfEXu8p9ZneXRypgbF3mKfUlO3EQXw9RxYpndFOBkJ+ZvyYRKIC1imZbmH
wKfgFCMHsndndR+Dor4B58cnDR0x0I4kUySS06WttbSI/6TNLyugzDTGHABvClG6
ZXgY1PykFwRlg8vVFkeEFV6l3WDhHMTY4UoReASSarQA1l5T87u5Jrd+XFo6Gy0F
MN4kpdVeNuiNl3EKQl6qVlqgeRh0zGpl9ZZBGYumHxHMrcgphkUgvNUp/0xrUknJ
aLnnX+2CEWyzEYPh86T4+i9N432/rSrsp2KQwCmkgrZYZnriPUQGClPksX76bObC
Xl3vhiDjUvVMPjGiyAxJjzFHPQT3UmVHZD/mD/j5dMWMHFy4Kq3ILsGZwr9K6cfP
zJZzw+3fNgcRKCjuJo33v99VoeUiT5BwnJn7xp/dwASePbh14UAGat/EhbXL7YaN
Y7QOzrA5kVS7u6hXQwThJT9Q3zyhCXHMGCOKf3DGt9iB3x+DROHJFFx/X9ZVA8KD
0BUP061jzPOATsDuCyqAVXF4+IjoKuDfRda7DAH3p3kDlnMg7Vk7sCG2KEP1SWBa
canRvAphvzjg59vatZgsUPgFFSkaoUVzpcEdCIQ7DiDX/5Fs513yh0geHm8+BB5J
8HF3Ejhyny9hKC72nUDVzBnpQpoyZ0Q+0G4eKJwhiOqNn8Dc5941IXZ9V2OHKQe0
md8U+a+wPTSlS7s9s5nFqRBR1aGvql5uUdKnc81jlKVxzLHWuC9sYvp5tWmG3Hts
h4iqOkCjbNtyq6aYcHewH0aq7zHlcoHmmsdefo4Rom6HW2qebr9M8fDfK4UO+bMO
bBRxEIN8HaPCItduVsgW8MbRqg/LOjIFWDVkj6W2fKuw5PkjUh7WhrgB63lWX8Bg
YpseIKCYT6odO8y5VfcLnl6vZ3SvTua6QOEb+17UHVyeWSS13ImYhko88PqENPrA
nMLqynB3U7gDm/4koEgG/ZQ5kzaG/CHXt5wccy6FVyu/J9kUWjYG/9A8GkuPpZxh
79ZBCFOrWWDi6yEZf8pyUDl4H8hn9jdgR7QkGcGbMxjTqTsmHntJBotf5vhBwY8m
kgBsSbbrjy0T/ZmpCdEM6NUm/7o4/Uwd4ApGz9bDCCloCHAxYDpYQLNftEZFZBEl
J11eGrH6PRiQpBA9jxtHcYqSsISFGj7SUVI06Sm/oxk5Tgn//40mj7pt0OibQX0x
BDakNhFmJTAcJqpm7HaXOu/t8FDek+WxSV8yXgaakYvplzeRJXKqvzjso3u2TWmY
BrSTc4yUrz9+FLxGPRfHkgMZVakQHNZNe02spBezWFz0iHtaYHtvTe/kjebwQXUx
7TFGxReIu4eQMO94T7mFdaWXLKjkOGPc1ZcIxjW95fpjY9CmFVau/e7V7cjQIre9
aQjhpsOKxnNAEhPF2LMYDydJCR+iqLLDZEGrSQHIHSldSqyTccXFNH9xER/rbLH9
laS3aUx2cuJGqw6BmrhmlP/ofxs3I7MinN51irIV+dV3si1C+Uzve6C3ppM2JsnW
8TzL7SO8XiKURYywLt8ghbZnP2SBhJOkkZ1qxQYIVn8jq7RmHb7FIkjaGb0Zd2jR
coKkZN5cumaHWAEijDIqa0tuTWI68rnITGlg1msrR5U46BXFeJrP9MPr5QnR0Tbc
KDwD4G/f/yIXKMUHf7GJG6FKCF8uR2KRWlZvuAEjzkbplJgMdjcCHjOexTV5iIsY
hlIQUVUWDkRkD9oBq/EQiQ4icVP2AxKFS5TyeyrHQTg1U25f7mTgt7TAxkQREocG
d2u6nBQcBFGrQV+La8/Gibu9o2bAYYQ8YFP4x/EROkS8iDB9uRQSnMa4XBqHvV+Z
Xqrwyuanurx3pb3O7+/wWn/9dC/hvD0t9egY++MS2nkAwRrPw1PpBFDz3jwrISjl
yZuXLBkkImDYLmy1PoZ8ilGEBlcq7w32Jg/CM1MEg4UK9esSjshdWBbfZKqwbJOs
mo0E0pM9fELbFt/oGqChFpuVcypEqnATDIGS+iESopfZc17hUteuURkMv2uUDlY/
Wg0UcXm4laC3NmkMPwxeS0VHX4YDlvNA/40WzRLtXt0LwohNA9zsdOuBjrAnkyvD
pC/to6qNmMRalkn2o3fMuRzwFlENCfoCcjf/rs+1bp/EXYBz4DI3A367VaxUHO8+
D/7G9QFD6xCa0KH35mYtp7h62CeaB3tZm0OLi7vUyf0Brve+WuyH8y98GKxBFqVc
AYyZPaSzoIi0GOwpnV1M8bRP70VvUjQdebTsrHnqvksP9qc7TY/xakOshKJtkU8J
kyHVb9SmRKGE5a0RDmt4pkEb4H/Og45asMaX/UayRiwIWksLHKOP39WAYO5wyzef
x+dxse2+mNB0JRcyXTmTFvaAGuQ4dIrz4q5lw5oOzi9n7M6eM/odrg8C7tGBlfMH
vupUopJ62q1X7CxLh7ZIgqn+fheLiSGfP703EmDDTEkorjK5gogS9lJVJo2QvKPY
f1pf1Xp29YkaI2bH5XY+1WyPxKhm54z1qF9jI46yuvzxZppaD/2Invyg6xjEpl56
yvMWBAT1cf54qQ3Gw9jA2CTGCj3yo6wIE2ttimFI5OPvYye3+fEvh+6pX9ZTXOeU
y7cECucEpi/r4NldVEq9ntmH7GhR4jPf8WtlfEtLeTXKIraV523Z6lwAUOnRfdh2
zaS8dqIK+ujtpObA7pO9gLCe8S15IbdiwMGZsIOEwI5M5P4c+tr0cS1Wrg9GpKoS
XcLWRRe4UMEsTyo/idoEGW5XC9dAH1PLtfxKxSoYiByM0/9oerKmFl99N0R3iuEy
VATew8sP/M5/H1M/dHioa/o5FldVCN7b3MJS8oLT+kyd0FB0vCV28Bz8pPFNeJhd
iAMhgvPTvrBNo5xdhXjJCG7/MuDL3KHLVMlsOSdiykdlw/LR4h8aCMwA6UBtvIwC
XLOGwh3ZL0aa82DoeKc4sjgVwueguHLaGRtbMls9+UHtVT4ZLhTPJ1DuPrxDMW1i
ptfqOw6tBGjI+C+3qEP27Fz/6NkVM2b02ZkeTJK4eN/8DkNQHVzuLt/H6TRY6sef
vnuFcA29QFxwPBV0rT2J9DrPcSgG0VPlDY+dx0XfpRDPde5WiouX6UyrHYql6L2e
G6mVfFlcvo2lScAV+Si+/12jt4AOYx5CZgZ9j4Yawc/jTnmEyH1AOJVrBESh5jkY
ROQr7nEAaxBJ/Zmf1lZ+zl+2qvssPBe9+O6VL/cJkvY9wCD1g8wt2/W7XSr0d/zz
acEIFKvS0WzbQmdEiB6L4xVuBpBf8AuKpzljN+7zDi3hPscevI16Vm1PUXuEk1QS
TxIpiH9tOIywUKDuXDTWQTNUygMIuq5KFFU3RPtmXlbUz41MxvcIBRfzTnfdFVtg
d2FWZsSDnUvmQBXsPWsphFNd69gbo7thv5+tyUo+Bkw7dmOW3gaH6h0np76hLhPu
NrmaIVADjEoU5BNRPuPI1QAk3w48l23FRTBn4rud4A6Oh7+fWAruM0igywgZT0Q5
H+GMomaPSASJscn6uo7/Bl3IrQobwU/OukMoX0k34e4JISGxsF1nV1XXzovT45hA
QhFNtamHaT5KMs/fr8zZQM43Y75wXNLlCKw3C2BBjLZ3U2WyE8VIvlvlRLi9xU4j
LR76OWbPidOndi042DbL0moVogCAjwfis1vdJJ5pg0AKTK6OMOFPDaN3W5gbSUTc
twQCctK7dYW4OA7mtl69nUTUe07XX9q88nlCNAJ4AwGHCcGJU1XCUqb3G/oz6IJ7
XbMtZjnrjIGgjWGUiEcjBlSi8aEVujG62M/UIaxYivfm0s5M1B88JLhFgjVWkHF+
elHbhAv9kJpyPwu7xUcwMXk2qE1vbz81JNs4q7Qph8qan9FRZ9KRpL3lPow7Vwwr
fOAGdu6yeKY7eVkbfqd1kLwPWyxuNjFSbJ3Zm/dhREhwZJPHXHEeVLYGrurFiWOa
OzDSxmxTkXyiWeBCsUDql4ozsIM/fqx/bHdbPLwvabcd58A5RYCwzcTzzhUzG50h
3l6qd3nwrUyHXiDVlPGGteCAR1LuInrekDzBZOAVeH3g9BdY3sU2yI5cE/aY8lgM
o27Oo/2L5aWMh0OMNBU2u9nE+F7IAXirPmKZ2ndqhHKelNlBvNy6mChOsJ4ufz8e
6opKN5inPQJ7z9jhsmZ6vKRm7+w8d0qZ6AezK+Rizm/KPyqICXROfUZ8GQwgQ3m/
FKm8iIjTPpyISKTS+gJ0/v19jDSF7IKG3iRxneVU/ITUy7ydIhtqFwEuXaULimHB
k6nvqF077U5LHiRUjTaig9Cm6XRXMosQ3kYoCdh3LEAonZTCMOAcqVR/45e80kmi
TzH3Hzzz4qNw2WYsanyDRI8edW/bXvoD7ljg9Q6P3Ruep1CCxjtk+6DPmaIXlY9X
W0FzSczun1c59x/BIHKhjGMbxyY6mRUuQnMU9wacoFhqJVkN48X+PAdm8GVnf1P0
t2d9g0EyxmlnuTQVEqrkTi9RPrlDAQZ11oEXdZ6/Hy5MeWa0PegwtJ2+XqmUxxYi
mt15fymECtuQExo6cyUsc0ZRleavJKEx93V000z74YIFUUaHtJ1x5xupNOshco2h
IbnJOa/XV3MtgSeJ3Zi9cNgbuEiCqmHDBLEYoMkaQAxdzAjS6/v+8uXbDNkjnqQl
39dSXtEpEKjNQ+03jd7p0WmFVmh7zIVx9ag45VSxyxWD3ZMCVzK5S25aFxk95T77
MNIT9mWak++WqourIg/KD5uvV8VyrpEYaGYYztsa3e1x5q08oqHstVsFcmff/R9O
0l8veTozV/htowwDcfaSkxzkZod0v9rmCXmOBQOZzIt0pOdhrLtRfVbHuIjsW5J0
uiDrX9t2JpNfSRy2PkBGhIuFnTCbmRSMkKB8Wnk8uICAgzhLzxjy8nkQw0cpw6fF
ISYiFmRcO7zw2nFMX1R5Fxb6lUwFehXj3zseeddgOEkHUL2Ju8+covQdtLTu8T64
9/6KUOgyIWp/Cs0TBdYlETV3WRosebOJIcXrjM7DdWp/whA6dsbkP3MTVH4ykdDS
X5xsoOL6lFcmVPlINHp7xhudAPqUrDGsoN4FAdGnbGywgrAQ2wM39BaKeUgzzWe2
CrTkukLart0gnZ5WmldkEBaYch+sTuWSWZDuytLw32mG0onfue626MwOSOcYKRMe
q3lOiiGSQaoVUPF/ttOLO4bnGkkqJZWFYAD8BFvE7m5K9wU8VeW2guQl4eUr04AO
4InSTUX6MG+PqGdVx/b3DgvEcj5+6kWwx136u/I5x/lyn5B48a5VsPUgSJ8dmN+n
eKwM52bq8yG7GJcCeFIsi5rJwpGmhlUn1E7MfoxqhEDZljOmv2NBCrvc6pFRvxaN
bCKOyktwY1vyRASykHM2zSaEyHN1otGaD3fWH2309qOhmSrEbfOfBy3izpeT0Jbj
ouT+bNpkDWjxN3XnzckSNdnOF8a8eH8T6RIXxY99pDcT5HL6oQGA6ouLbb/DGcPa
B/PZzrZYHs2F7fb6ZY/2RDSha8SJo6Im+OpppficIA/nO9QuuChncYbJIwkHGqOw
fX+trLqQrBfO7IkwzfPfgg6EPZUxxLpX5PqyGegPTYVWDL8LS0EW2mkJY9eKUXpv
jt5Sw/hAPhYPBlmitqPe9P7SiEQ/IP6V3kBTShOY87yudUXjHeNNCrKQM/M3i2Al
IlN5NOR1WNCCMGALj2Hocs11J9uyiGVLPiEENZqcmKqtIdHljiApsP6DW5OHN/oZ
QgzoC2C/+BooiC7wxC8Z8cUmjGtAiQabB4nk7HUptOhSkWM0cS8QXKPE6sYSCy9R
4zPOxLHx9eSI9MMy9S+Y+/UTGLDe4lYAOKaIOcmf4jQlcnFcVUk3Quf16F7jvZv/
DmDj+2owevMkkTxR7OV6jj9HYsvcreS5bKzfqjsNisixOnRj38WjocCa1lCsC86i
ndA0FG3At+i8LR1YeCuQx2VB0VSiMHz8FQh+7oV5ohHpKqCJwMHGUtDDQDtUKUod
BEa0wW9dVSGCAREhUhSm1tCFe2gOf/VTrYPSyxN14f5zb7qBg1xQHBmxUjfk6wsx
Wqe06JK11LcjOX6evz6t5MM4SbLq17pbciWxPmJtkrCZ0ufln3Xozo3RqYP91br6
ms3kvysllpxqPOEW2F1ds39Qf6zAWELyVQGmlwtuv/tR2ubOGQaX4wXAPNUhsPY3
WJpEVWOX2Z5uBuoMDcW2yiUQbWomDLoCTOSzBagoFpC9PLbWqqFDHLSA1NtGiX8Z
ZnALofeYT7+UywSKZgmSByUl7BxhBelj23H6GkJWvBWxdMlR+bHET4zWaUqFntSK
WY1t/21jkMoFsrr9x0hNBMDDHOJDK3cxYweofR6mH26I/uEN0MhLW631Jd5ZoB//
ITzio0Mvs03cLoJ6JwhlkThCi7CrVQxLphFDcfiJ62MRV8NJhc++yKfD+3iNezcE
j4O2XCWWA/rp02wFkLKer43+oiu8oXpZ6vFV6topbypr6WkNLjHXZfA6sJo+pkaQ
TWbhCZbdxrtl9pcBGrCZhhiOvrNnrHoZcr86kAQNRWcOQ89MvBOkNB/ZeE04wasZ
Tr090oQtP8c9QC4QeDPoZZ5hPyd+5yE61vtUDb8QqBW+XDfLysnJOaQ1TTmeFMAT
Hyy8laCyuuZD4tGIwFUq2xSLmIqTUW8CGA7t5CIU9GGLPrPzah9QKnzL5n38Iv9M
Z5gG5wzhIT6KmQIPPxglq+a4M13Zbt+5+xXQf/jyfEfxy1uDMQJRVOu/w7pmQ3Kx
9kOeNSoyuksZnOBj9iywsKXiDuVrTjxmdueWiJJDDAAA1oJ2C4e7JQO60b1JPEoz
o5lN0oBFF1z8rODc7asYxoBrdm/zYDPWT55yaGjScs1qmH63cZN0Nz/euX9AXDpP
xLI85OH66Tm0AitIkMtN/zAmcWNT+noycD5lJ3AJoIXZyjpfMiRil2L9Rj1cnqjC
tEW70sSLLY2gjOWtEu56cNvhKdfqe3dwXqOJsA5Z6ypIOxXVMkDX4HfDpQ7js5OV
e8sQSP6hcjsNFpqVQ4hRTrzB6Nfiyu8waZ3Ks4Bl7rC8WNp67XC4ufMeqdrkR3OO
CaREpG1c2QHLX5BERb3OtvCX0TGGHyfDbE3irrGXwmUpkn7uLVmt3Ubx8IUG5Mmv
qjpDnM5MjZJyGtfTCdNYUSLybOgzkpFx4msfqDewMZGoCfulBXCckLsloFkfzLql
qltcocIim6cfYIF6DV3wZXGuf9EYKl8VAMveqBKvaI6iTRwyPtG2NxZf9QUoTNdF
FhG8Kz/RStkfhjbl3o/Ds6++afAJaqbFFen9/W3B02LaGP+rikAuxIcgBzKZPGEQ
Zo5Jh1ws14HSskuUYa1gQbR9oPyCcPVx2TAtFXxYPxcZmOiH8KQy+Qa7AOIeCjFM
kYjuE1Em//Y5Xd2FhWjfnnrVu4G81WKKmgrEntGuRS1YfMFh1EXZPz0B/YJPGq33
0HyuT4XEMGeVfmJ9WuEmyshe73hrePoROFY0eTzYxPmshC+23ESGYsoYhdsvKDux
P1PaC14Cg4AUnVaFicubN1imyFjvAebK65LVpgbZS/G03/5ECIawdqhG4Q+6kAD1
RrP80pbX809RIt4N5ZAl9tPlTSVU6VGlT6nzZRlLMVe8Rd6sHplRKMo8qPbCqTMX
jMPp4wPgkXlfsqyopG7iF3IUsxeefyWlX2zLzl4yAg97mWcHq7rF4qa1gRjXWG1x
bjo/tsFhI/oI0VHVkQT9PlpclALwGX/Khv7Vd18WUVRoW6WQqsr5ZVy0YFIuB5Up
JewleuwjgvIXr1DcNuYqdR3UxppaFTGuBI45pchFX8wLUWYbYaOU8U4ruOtQd4wN
Dh/Qjd0RNUesga/jyZTFKPrQ+5B/s8eIiwYy9/3HFigawWrmWAruMTn2Gk+PvgEc
Oy1N6dlq0w6JuNppyfkzIu36hhC8MXs9yAaId+CbPuOigwACkE4IZNbEs+6WPzV5
2lSSydSXi2OHVkJl0z1BgKIApLnxi7htp1DV8owU5odfxAvlCiMjQb+ZRqahtYmt
//fwcGz5dEhSDZIk0blrBBAwkr25zOkcmJNpRwXq9DrUVKOGOCLKFyg+EkOQHTyl
JqcYD/HE9A6L9NNOMEzuRXj5pDLEBDWFx5DIOw8zX4qh41lISVClDYfHEUvn5v/y
JwIRN3iihGcrLQWWMwM7UTbhqmB8QVKkmXP6c4VeYqgTZZveufEh9HTHSwuO56oq
/0LA+mTIac7sH/iYiEurlOLtSAdimGSr4xJfLaXy4QuddOVJEPo+vjq4EMdx8mRV
Z19VW4ulnyMYNBKDzirU6qPTx0RreKxNgqer8qUjSRpklJHscChqkl1NTwLbozAF
9hCUY9/RRfMh35CvjMQ670QXnAE1XWQ1RJfulD+pwxxGft5z8QsMFnohuS1OLt7c
EOo19uSUwhX3+owjcbMKiOiD0m2QqJm7YIP/EpaxSPOww+fOdG02c5GMPq8FYjwU
w4X9c9aPaWAoJj75QS2jcA5pTwoMgwftg9u0rRq5CtVyrFzjJDvtRXTBFZA97eUb
HzNT7lH7E498j3qyzkX0Dmabt8b1ycGSjFn8aE+mx+8ejLOHxCbyVe9w997v0XgT
+zPmVo7OqlUzci79o2rhzU58CdjcCtUbGJrFT19hIO5bxmGlRKyDPupgULjtXKkk
3SKj5d0m+75vb3oIJA6sRql0YnPY5chP83Y7Inu51LXR9w7kBJltdLHYFscIQqNb
hwz+B1xOtv9R1XRfYgKluK0xB6f0DHd+pcYZiyZdoYUKlrI0S/ySr37Op4vd0Uvz
7A4HpIfoIm8qoQQdkkj/b0W/Yy0gOPgPXV9tAHZ5S7NeGD1hwFh7NHFcWW2GaN4S
CJpYROSogG80BcmA5tZznkXLFLTwwxoQC77/xW0UmAuBaWkrLzvh6S4yBr8fZB4G
3ydkWHAUjAMOmR0lvWmlPR9F3SRJx6EyO/ABR68aNk/nxlYE3zuveo+kB8Snyvxl
CYXzqhiGRdqtPSUtZnrTz/rv3drfcVFmUbTPbxFQPJab9eJ6x9yWbVQYB88dr/FU
lrbUflMTMO2nkziZ61FDberhyEUaYj4qJMH3vDd02xQoDydGcDK7+GyJRnzgRJ+d
XO5Y8GziSFVTEx94q4zRGLlJD+SjWH3Tqqz+IC+QxVRK9J+Cz+WK97ltA+eLxXJm
bWVt8baaEdcT5cUi7dQw5spc2YycPXYFPeIcBRLvc7PmuB0F8CdTXgE3Sz4EYgPW
L+qmw8IwYzZ95PA8hn/qB/fnY2FBGoPuUUH4rJzvQxXGF8TgEpxLYc9zR6ETF+VL
bk4FEOsLKto3+gk+Ps880nfZqlEgeOqJeugr6WDcfuYrO0EBJFuKO12n/7z40k4M
2ZbY3eVxAAHVbfluTL+rYS/jDcL8LGcIEgaPtfSXmm7WYiq3cPTbfH1fwE/kLNyg
4MvODqpr+C7ijU6AOhk8C6F1pNBG4SNRLFa21maByMla223uccXWaLdQHe6jA66t
AscqOt4hiww5v2mBojDCdQQ0dK8oCn4XYi5WQuKUyYQYHrix93KFMSSJpRW8InAG
Cc1SORk/fA+kKUtKY92SK8f4zTGQr/+1i9NTvdV7LMO63PHMByCBvHh7LVD+X8W/
83nwQVPbN72n4PipJY1MIJIqEN98X+XSDpRnrM1sZF+xQxQQFmGlqUDYTFZf0/ZM
dbwXeRCY9+wrZGbflufACufx8HKwpEs+wBRJDG+vK1U7EwuUf5OQVo+3j4szdymV
E7sdo9+w7t9N5OAadHkThB34GSyOzzaqSAJjs0MzFHoM9RA3YmzkTfTs+gWV9JCZ
z5DRgngI0SdVyWJqt+tdbisj5AYnpQaQxfDqW8oPW/z9latYsPp+seG1rJxSgvvt
Ym01KgQr0tJ6jo61qEnYfkteT1SUEYTVfA1n1md5iJ+BYnO7a6mQeaTkeyvd512J
WsK49V5J8QD2KVvj9ldknWfvl8kSieQQvwN1TJO+uQo7EJA86ta9gnrfp6+gFIwf
dAt9iLWwBpflCtNyZ2O533CVbQRNxpZKgVcf71KS+h4PbXHOZh1SDb5KU6DWoAPJ
2Y8wIc0cbWAOY2BXujIOteaUSHK7A4uc1lZTRzJorQ1VrVyf5Hjm1VOJ8DguBPnc
5FFU+hSYgnpzLikQLuIyBOzkl7DaUkynnKw2IOxJHTwO3fAe8L3j4Zz6xp6Enp0e
+BO+edebDeXBc7b/k1izhDhu0K1qvwEs/7bW/abRX2sNjeXS9gnCgneJpbc0etgo
njPmyXxxbgobR9Pj+6BKd0ao9jePmNm1kHaNOewygukyN7JrOJvdChD9s3Stld6v
vHiicfxoEgSIOrxJdICle2mqVBOlCt0MSkqM85CNgnJ6b9g5lJYdzbHKFJa+L05H
tIM2+q+4Wzbypaoisghqgo7yuNxxN2a9pxYiJhgtvePxZjIHxGRj7lXKD6u89AxR
vtYs8+R6U/1WeUGmUPhpU5iZX83BLBiK2PEfhxDmXcHjlpsh7G8nBl7/ecC3639Y
VZZ0fDD6hvcLznusR2EZ8PPRM9EPfWaJN48zWaPeX4WfEKOJhMDow2bdnW8esGux
h8S8gt+lSb0vEU+CCnmetdlVG3X0oPqVr0rU0c6/FgddYNWmIDTqqweyW8kXc1lE
WX5ZaWdmnvr53y2u8kf36RhcD/V/R7gTqoJVsHp4W4vy9BgK/CfrqsVW6N/ulT41
ATOp194r55K4ijtYIeiwAoWzthWqIDShherutq+WcRXxpc+F5bOOTTu5BvQk7b7G
htqpTrqsJFKRc+G0VO51AZBHP5j2P9rD59+pLxbJe0UAtvHFwuxKnCFdbO8lEtml
qJrOktkCayfPV7x9goi+rE50ajXdE2yAsnCz9GdvUbWJzIzL+MDoKhCIiuQc2gS3
TMDDyVcJnS7Hs2rnsRJ0M0lGpuzbV9PKvp2Je9uMG7HkZSWHSueNU8/ynA2sfghr
PtC6k3eC/92/wFsm5lhuhbOojp33fNcVM+Daxf+ZZ5NEADpdKilflwozM6jdStC3
WzcH+B8omGrfYqwtHxaw3D1qVQWGgYNy2qS9dLhBltdfegelKry9bNhJ43dECYme
v3yw8DC6caHLOS1oHBtOzZU52D+BQSw4Ns/ey/ZZkuG52H9Z2JOpOSgi3CjxbkRG
5N/O+hrkrOsDy0sohYj+drMrpgrOOoS5ya4UWb6CZmTXBFyP+ws9e6ifgf1chcij
W3jKClPbsbQxwua17XnrGbhw1R+DjY3pw13dSmixpuCP/CD38uldp8herArNi8Zo
YRQNYAoU5pVxYdYXx5Wppxpxqvsg9+DCYmol/c4b1JXPAw+dNQTO3kTkWTBskx7I
l67YQeopLa51Wl4KxOYdkE4FXURxrZMfPB3IwFtHXaerVh0zbGqw8CRSJz8x1iaf
vodl/qwz3hK/kaSGqoVIzD21gW8/x68yTXEDIbbArkb/HunGJ1YF2Np+578ruMUM
RYD8suUR5GOHV4RlJLmnRwW8rTki23HymEHsisVqP8X/S3AlYjb5WaDNvOjJ0w5t
G9xOxNXBgEkxNRNaIiz8pF2DklSqpXMccCPjKxKhLcEurUEz+10ANOqz9R5TKhmh
U4lbB7N9feFSutI5PR5FPkX+r4YHvuR8Wh3CK4uP524/dA8xYJQCyYIIpdESmIOr
8KTioWQSDkcYZKcc4RjIUoamryXzpLTKmzV7DZNdwNAp3ZFiuqWZhM/kAfSUFgf0
Ram06EoZ3Vi9aQLmqA3X3YLiLoeiQkyL/8ddnjaHKDp74iwXu/2acKf1dVWpqgCT
HRTHzSCZnP5SV7CmOtrXSQUPI1DzjIzRDpo7U7589bfBvgZBB07pmFrd8OajKg8Q
sYnu3YRXyqT6dD3HaLADLMJueTfjmJNStanWFwuayhmZFmZXDcmU+YzMVTVuRuab
X8wGrl7BPAQELxWP30z9mwtPm/4k/5U6ayEj5Q94N0gXW70z57N/Tc861nScS3Ne
9gMtZ20acaYiDXJtCgtvjD0qvWquOqS9yLdya4j3oNF4FSoGsVjfPcts1F2D7c9g
HFykt+rCbikcEosCVyV3fhgN7v0hhVwec2D8JAQBzSk/xlWxXt3AFs78Mi9NkTew
pNg+qaCJ+RKBO0hubyvHP0ZeAbZFyF4drlwVFJglGxzd3fvYb0s8/7uI65mVdTq+
id0woYdNn0kzeYBeYMdbpwEHirWkHSnjlJR4AB/4CDnngeFRFZheiNCnUY9BJb94
Km6kiVvkP+L/se/AUEfhL3dW1aPE8jinxhixgfn/MjtoVE0vZE9X3QxFEQAJcaHl
ABaqla6rMMu+AYqCQ3MQbr0uq0/LmG+llXnpV79QLAFu9ZcDdDSeqc/VQMPcSGXq
Hw0Tyh/CJpliaQRKzaaSc3fB5dhdD8Kz7bUIM9tnGWfCI6+mPmOhJ3Sp1ZkkNeLV
JFHstXUh8D7p4UhlcYxY3iDpI6tJ7XpfkRo1JVtULR4Yaxud881pmF5uMcrBKAun
66p6ELYPsQJDxNBBn2cbsaM4nyL0z2/6/5Sp//V05rzIjav2Pm/w8il9syMXf9Cd
ZgI2ktQ+L9OvEiNDxtP3WCYO+AIz5mhPaMMJCTRPF+X82qw9g8h+LfDUChEHSBtT
xixu/YVCY+DcsTkEaHGjuS2kxggNtbIhBFSKvQu8QPNX7j7e1lnSbndYK3All5np
1FD+i21x4SZS4Jug1BzzhR7sWJ/U8tcNpUdXk1IPGO8zl9wS1nyZDo1L1ySqRUUf
l03M4CrsEtOTDVRfjpngtoMVWUEKbjFa0XC1qdPpeNwB2+8OpJxohZoaZhmEPdNb
mpamgLOsopuMLO/9rRSAW23y9e+SmFRjEvbQCpdpW/P2k4e49oJ3Tq/99wgFh22c
dP5oxhEZ6km0kDl20vIjol2SsO5TMBln8iGecb6qjAzNhXxBksn4phYiCRUOqqIo
gdaojY5aiO2Vj+ZgHrlemNHUmSLArCCJo6ZyNqYGDQnhjRHxfXuwrHeJT48coH9x
13Tlo68NugfNRsegmBJwGYfLZIzw6O29elu0WDzlFQLwXXt3CPln4geOOrqdWkku
62igrz1OhOsfFYQWFJsHuXVN2A1p0wYsSYVxl6Cf99rboepyWT/A5cY3k9kSSXVa
iHO+xMz/IKpmPKSC8RGUZlCF0WbSzcMgk8E778a3N6U9X1+W9OtaU1Wykq9qu1Uu
TLAItNpebNOICwyC3f59DslBAVvfIlzCmFScqpIvwKfNyzGDRKQdBdEohSQ8b5ob
HK6UxI1rO3mhm3hVKj9H4snbFlFSAAKnECTLxTdKXiiB8j2jePPUYpC8+PL/5TI/
uy6O5J5Tgtri3+hl5nK71CW7SXnjFkT3i35R/3akwDxn/YJrZsBLRfcN9chGoyNx
5aAKeomX1mAA03nol5ZHtVTK65mDQC2IE0qiMU7GRW9RZ7yjXm4+X+fIPrxpYLIv
ahXUhUN4bfvaRt2/OQ6nGM6wGFkFp5X06tuDKeVhvUS4UjGdgzWD0PBu8zS19DHt
sRg8Mp+BiWTz161/7+KfwsVzg1gKkIK9e+/PKOtks2bjbDa4B0KR54EQz1WeUp6a
WYNUJ9obO6sUIxGmt8iOAxuuxghU4+f+KHzZR4bcMAEODJkrZIGyE/Hw1CZopfIR
FlazkWl2NNe2dFP399NNzq1VnyfVIPtV+tnuX/5l60zStAPppI0EbLD46RZj4Ozs
+MbJO5Oh4s7/7xq2IgcwrGc5pn3HcxRDdUN3wYjRvkfxR06Q9TEuv7ITBMF37zLy
infIUVA6zLIQQSaC2Q//FE9NUXJG0NVZqQESxHdOv0oozaYWWbuiOkYnEpsRN/cf
KOMpvXC9w6F5gMHc1f12to5Nngvn3PGzHNlatRjgv40WyzpKuzfkhpb1kf/Ejeg5
DLY0aiajRE6X173gy0YO0/svi3BaNf68aldrGbPXs2nzheuVeHyaDqceUtm0wObP
W6yt+EcUlCx2CPx04lEalTrOruUf37a73+ag5LEDF2kxGYfaXW3CYBmXEcX4QUff
ot6GbR5gSzxBBuljMH5McU458qH9QJUdw/vZevdbqia38dOXXFIFPKgpdkWeZohX
CT3oVUH9xKJP0iiuF5T3+vQ6SCx1qYvxIqc3RUGWO6NFZCJIlbmLKqWHRTMjRaPN
fMyiLCdeZ+ppZ7suKzWT9yLyF9N3UPa0eQ1hg3RA2D3zAOGOPsnlAw0cFdrW3whD
XFizc/fyre4osVCOXFKcJVCByaQBSNN73EDy4sBw60qN9InVqNP907Q8Iz3FGANB
BvA73jaFEssGWp21xJA7IRILl/o97qUKFqMDeIcLQIp8EuBwYutR3rjcOvyM3SPh
nW6mIh1q1jlnJ7ncifJYdb6oMwOowqYgz0Gtomot7xc6w8a3XHUptIpJVm2IydQ6
CvzYM98H9gutV2x+wTmSy7Bqwj58AESGdRgIbNPK287SVbUqoo+lltBFa3pgqBxs
opbMDxqfRQbVvGgTVdpd6IFlU3KEdq7YrgkoqU3/bFa+ydEXHNKEoisjfbz1SEKX
zC5FMEb7IsR3fRfRoCg+3h/oHZov+FmuaE/inzN/Y2t6jiVsjDaP0UnaGAPmQO05
/1L7vHDmbhvhNUZNKwKtfu7/uUsoIVjjyeCGs0niFULz8VOsNeXDY+0AlhiDgZmo
TzFPPYvduzdgUWv1YmErRL58CSx++sEjGGG0STdxh0dt0SbonBD/DznW3EfErXk6
QbD7elb2GFlEnFicd2gS7OHRVpU93QttA7mnkDjwyQJJ9o+Fa/cA0GcFmYLt1EPD
3gQV2ticMn7DHgULO4qwEnBX3mBK03T/RkCcJoP/G1XV+yCsqhS2zsaLj8BF4FDh
f8gwLVaDIpQYKPeCkf+qTSq4rt5Y6OrNkD1z4EROXJ/GrKrIUzE9/rAi6ibfOkBQ
yX3J1YHcTotwCFTze6ZzENhxciIm3jJDQYCFfFwXEtN6SwnebEPVqN1HBF/H6sMC
69JVMDchveVAi4drLVyvU50KZDrg/ae3HcleErxvALZah9dBuQYY4QIwWE6yXAR1
59Ckzg7j1LD+pqD9ig01Hft8bfNhHKcf2Pmq7fb1kyHfDNl+3gbRiXqwYsTWOQ5e
qBdr6usrr/99EXiRbISNmtndQwR6uLCcv9iT426w0eYI8GLlDOUOONfh9EDDE2tJ
NDYRFIUp9B0253vfMXbjncpGlBlrQagQiUXeENVQIM7NHvnZg1w2BxPyxtevAr9H
qpnRVsuk9qVnk0trGvVAu95U8NBvaDqe4JhxQZOl0KSBb+vkC8FAhhtxPnUoS6yJ
VDqR6J75srZE1gJTBhJA4E8E6j+O17Std+DSad+DY68fMbpXwk3iDxPvaM1updx6
eMh00Q4p3zXm/bSjJw24m9G1WknDpCcbDrdH7R/E7e3gVueSrWS/LcFZ6Z5vtgvS
h5pfI/ck7Q/0A5QrX05RqViTAvWbWTjxcetmqO4A3DShrct4PvAYDRHgo7XGBzIU
n8uCjT7FWgl0nIADt4aO9vh+V0oKeU0zrWwrhPgXzJGT1sQMKVqfL5eAiksyc3y+
W5dUGaM0RRWYIth+SZoinLeOw1DoWvvGfhHLfGTgaSzyVr4JkoCEJmqyAbWr7iaO
1yfGNARzFRrFT0LVt3Y405FQzQRUceY6jierEVpSZeplov+7Xamywe3ZN9fHcaqn
KZJOljykRyHw9aYHNwDXOSAo8/u3U39fd+RrkLZLhi/3LdbyfkB7gLYklbgqDD2x
qQmWtDjyda7oAmksrB8CgBYIDB097g+hbnaiFqeo7Q9F719fHII9K5RiRin+8NZB
i2WUMr5TryILP/HwR03lLitdpvMR/HffjYhV2NUOCO9qefRZEu7lbzJgxhgalU/o
ReJeHWC3EiOJi1/zaNTEMG85dh4BBE/TZmyGjXIFaG6ft8frATkib2nuDQ77POf0
1AzY5pwdANAFtE6HjuUBCUleO4BKHh96pNL+TqGlDGkBD0zc10Zfhoy8p+pFAZms
ztRPx2VvdAg/wk6LfT7vhEPhh2wuT94CRartqHOYbhd0ALMNisG+ERl500w20lZA
BUrGdF1Te4c96T2KEnQguWCUmulfyV819aa/xhBpnX5gzD8DFuLfbauzeP41s1I0
`pragma protect end_protected
