// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
S/C8PH6JXjbvE2duBiYiFwb0jFTD8ubk0BmVXf7GgHFQyCCrZTbqpNK9dKBaJLhj
l5//03hGkDrRKb0fGsyICZJETa2tKCywyJ7SoCLUadUdevSB7tzqmJdD2RWpE5Sn
x2BoTbISTHihInazk936sgOCrNsqaisRF04Dv39KyYo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2576)
FNJ5Bps3FRVA68NLJXhuTIfW2PFMhxiZu9lEdMoNVS9ctrF3IDbgPby1jaePvPLt
mD8PZr6JhpmFp5xTQWiedAxWOCFxgtM63UaT6GSHN/04yVU9M4XC4a0lVxRYZBzU
qlP2izcTwU9ZU7hOQ832Qzoyj+/GiVVRHZtAzUy4dPEYNNvy12uocQ1KLIcnAbOi
h2Yi5R6z4/T7oexAvZZPEwptw68ME9tYCMwndj1QEzNPBfA3Qzj6Ykn2ctuXIgyE
WGahXostLg1C4SC6qM+ULfDKBA+j/iz/GnbJwU/wYR5RUY1GchMrtPum4/CvOveb
Qc9kll4xXQFM9ELdKkbA6XpQgEYGNQ0YOydDVV9MrxTAzJhGtTgJNet0SXJKiFUi
rGduyjfWIiy6hRVdZ625yPRgrqEVMeRgWOkfeG6FHxhBklMfyYefbQE1/E/yCGFe
Z1FTTHzuVYtwAfTmEyX0LEgb1sCEd7GIkTVpLD/ZLF/Reiy08UW6f5jVc0RSQURT
YWUaA4YHhkNwobOT3Jh/y8wHTwZfrQWLt29Her4mjy7CRcqIQxmSB7SHsxYybivo
0Eh3briTS/+u+G7UTx34/ppVm7U7av5Ad0arrvXb3PZkL6bHy5ySIJ8iUkbzvt+n
00GsXaoRdWkJ8jRE98gCZdyqsd6hZ9zTUQp3ak7nUE2tPqPogxNEebnUB6I5UNvj
mK/0HtDph3lD2mUZZhh0WUJR2zzRFZfWMDUTs92JEZMMtnhmZv7ZlRO+0A83ETjI
ZiwnEGw0NYLL8FvDBmYvBQ96GWO7sP4GNsltjFHqiClGd8Y5JJvgo2R138xIgc1K
r8fqDFtNsQ5+MnSH612DZGQy6R+SX9VcmGN3byBQRrQtE12rWPYWJKdK44ycofML
gYTxMNfHDR9jxMG2mFzv6r6E8BkX9zWUBoVKALyz/JFih6cVNI7IXrMnelfH0a6O
V54gJHzQDQvGo85ZBrdjhG6eXXNDmGg3neWO41H3+zGYsXMiPEHrWcNAx5kBCIVz
+hzXs2NPfH2OLHUCxXe0WOzi6d6t3Ozzgh+cR9f9UtkUIATjXfSxZuRTVDhssdzG
6Z3cZh7zsy8ay3eATsoCZ1hk+yImq7gwpr5C+U+oTbrtYKeVqW+JGh+g0jy8CeyU
vyEl4AZ4iWeyevr+8FcQa6dYufU97KLaPThBXWnjPcMPiYf4wdJBIKzupi2dmTLf
3hyp8kMrBXeQwi8CEDyjpg9GemJIRM8vmaXW8OW5wiryOFmKQJ7//7lkF57I+VOP
QswJWkac0frkNBCY28V2CqO1HvYHW2nNwxlQFhLV1G4ajswZS7x18E+yLJnyg6qx
Kzjan4wYYZmMB0TT43yiEIh7fV19jZdQuRPHaleN/7vvEN4zvcuivl1QlSGlC0tN
3+cG6l2li/VgBDznogAtkedidX1YIL8x09VJ0bjrEm0DQ28h5KuWVKTjBEm/ELZV
uPdODD4Ac3RCcZpv2T+Qsztr6VVhpsFbXOhm0bbU3oMcRBP4jVoM+kmDSEjOcT8V
KR8QgYvsthPuTl1p8W6Qy5+RlWZg5mDCnHJ/Vz/k8u+NxmzRtqeTX/EIDHsJqKlj
VH9zGiAPVwX+1zn6pzaTG7ABVRYXNnm3Gcf9hSGYpVFIe+6UWr/vpFKKctDfNoht
Qmtb4hGoNxm+i8XVNqeBG2nDdCLnZCLxe05V3reETYMPUL7k1LDIThweibgJaKXo
vc07iSABezRZzCxKCGb4cJ0IQ3LH3vH44o6dxaWh26bnaGMUm1E22vq5UPVT202D
DQm2YIz2mNvYumenLsOWzn7idB9NL1IN3cZgN1qfEuf4LqcBiki91x8g50c9KaiN
hVKqOV64zNYGubfJoqMdWN+29LLKbV7m6W94BAHIQyXr4jLejYiypynPUdtkTnEe
uEohilWYiUtsdzf0ij/NJ9O/UzIxvJrmPSmNn1eT4hesnfhTs0LleYmpsz3j7ti1
EnsFIkfsUcJP/F1GrysnBPjehIMnmxgwRWAJFzhRfwxc3s+xgYyfOM1m0XmCAG2Y
oeznSJ2QgawxldMWNcmomvNXSU/v5JX1/KaNOgYkxEY/64IQBtpDE17IMVxPimm5
ymadSYNFiGg0wy2hjNhyoDtNOPM60VFoGxKFEur57IVOC1Fntvzz1XmBsI7C9teo
7nZTco3MJNim/pXi6KKEEZnvVlwz+Ml3od8jnQn3RnwLbkTHipAVG0WFZXCxNOfW
VwlFS978HlIRcoR2affxF5zl5qoCPGnfGREdBgpIuYpjkChWHrUCeZERNy61KP+W
82sPX3pMznF8VJo7IET/Y0gsrWhxh6AdrOXnORhjlpMABPzk9Jk+zm7bgZB9njfY
hAuCDL7BImV8Bt+EukZWeLfdYn/T474EFy6SmX2Y6lxUHpBhkMGzOEtwZCwDuZRQ
J8FGNfTb2/WRC8lGURiXr8z6ZbvLOAR6MLwjn1uS2QT4ewjj2k/mQN1H9tOZyK2U
8+LHz+ziPC/JQlO/LxwGd07LsIWVDRoDVkADsXXyD7f73W4IWa+WS4905YVBraUc
IseN+iSSSft+Bns5u8/xbYoTnUlasMW/OSEkHulVm/ZTSG7OknMksEAIhe/qZbwg
acuQniy5+xXa9xkFi3prE2eznJmiuNnKJc6D5MmU8Vahh1j0AaKGe8GUrVd7o4kw
vdhUBBH79o7Grt68BWqC5r3O9o6fhh4tZYKr9hvHN7qKA5LxW6gOXfvzGvdpwVqs
XUBuDcF07PBzhOL8dBJCgdHAnBhrfmuhs6vRbRpd7fwjB7Un5ifDju7ukiUsAEtk
jBdnnRvYEiNNssonmovG6dPaeMqy0rmR/ABZpyv9122XXmXYvYafRDo3kigEyfPg
e8YHR8b5iy7NiQ9Ik7f3EnGmpA4JKWJmNhDGrq38fDLHxPX3J0oy8nE/ZzQ1V6mj
EQAudWcx7lCDN4tYtM5mDNxI/90K8mtZpeAeOdd/NJxNP6BAgGTnVWKwquVyBBMQ
OPH/XFzgwuzKKnVxZi5XzQASbfxB2tohVP1iefAs5yeE0e6dCLlhm7U1XJ0GMuPM
WgaEZZZOiNRNSOA88pcEgJXHoLfwtBgFGmicUS/E0yGjBL+iTJjCzIvwUvuXY66v
xy3qPirvoltBY3b0kL4P01ffTaimiUejew9/+7Bv5IeGlsmGRIXwi8Zug2wo4PqE
RsoopjPXIdlbxnaGr0L2DDc7sNJwdmKAFsz0Vd65oDN3n5SE+Zsst2hehGhw+Zxv
228tHoDwiMQ8JnIRymiQkBr1R6+na3bEusnTkTUmbEm/k9iSJcOmAvcgUCqEXFXJ
caXwHNhc+WI0ww96bPiAo0J6b14dXcQ7iCzFXP5AyahEgFEEuKa8JnNy4C4gkUWS
lBj8DBxmpgONx1Crl3NWK9H9F7Qh6IrKOHGhuLTClkk=
`pragma protect end_protected
