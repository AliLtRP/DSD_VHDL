// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
XNM5j05/oN11jqfKm//AWT4iyAb+hkQ/cdd2wDq4eb4Zl7vOg1wU0DH3Logm9LU935HYIE/QXGKU
TGmoi1xgQ/pXgVyVtF0D+yFtJo3edvzHWZc+abXu1o8uXYpuLNQ/QhWu50sxLUYtJPD51aGMCA/C
2HSqlXCfdO4NRs0eMf5sSDh89U7OXl8wfzM9ikVv2HTcsA+3OFVqgSRCfcp/oxryacEMy0leWAN9
tNtzI+j7QLguxoxJP2MI9j1FEbYUqhZ1yTdwu3NjWtQ6oLo29eA9qjUTfditDcpzeicCuFXRZt14
b5H4izxLTOfWnbAIvBj7zQDk6UE3gddHTwO9qw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
fvd//HbbvSi77585lfDbXDTOXZ98YsfCrxcLg69CR7SFN6uFv0eft4E7NBlBDDF+cF/CBeT0fbB+
2s2Pojwk5mbLoMancTC3RMZt/38XOSH1bcJlq6pFS9Oybnqh9612A4qqAPFkLBOvH+OuuTOF2MOY
yosYYlkAr+CLcED7Du3KP1/Nha6G6+bfwzD7XQPg4RK598m2M++dgJvhq8nC7xaPZAwLlGih8qLu
k2c+6Di2d8R6E/G4fgHKdDgv9ZD8QtcK1/YJDaYvd1fQbjOjS76VSoMco1Uj3VOPsQb7xA5VHgOK
tZfDpiBJrR10LIux+7RhLys82wif+qNjNiLYrXGHV1Gwl5xmDy1zS7pnkYh7OJ9uAJDZp4e1GPf2
xZ5OiJGxOnvCiUNbJR0IzSpmKQW+EO/EdJo1VpPha6jPRwow2Y/Z07OrKMr4dKG9trGUE8FlhuGZ
PG8mbIEAIP+1/8zjNs/BaiR5Kr6Mt7WJM4KgDwPOvc/FrKdhCgrqN+NHAnjLBWqgAf3GepyJqxkc
YzGpEpDu7tEwXWiHyyRG/Vh25p/kb9QA2MXEVClxgQXcAKi35PUtgLXbzjuzzEjfzMSaXY9hJeTR
z21dJ5DkXuAitI+nxoTbfqAlee8DIe+NJlXTNcqYJR8UOhNfQmsjsololoXI8N4sbw1D3rycgTld
hL9qoi9QjoC+1T5BnKIbXRIZnMtt/l4wyVEZvVoMUCdpeAoDfIULJBbMI8wu9Rn9yDnSyHd2utZM
ojzIJ7DvdNOSkH47uJ5+rUCunx7WBw/W544ALBGo7Q0Vq7VNfEcAteejd5j3Jo8hRTo8J/rxK2/h
AWBtBg6boNvaeLAjtwJoCwYhMD5DqD1eZas1/tIeSPQDJsoQMYI84LlOhBLrwi32SIlU1FKUItZl
mdanYpPkgjSpA/02xUP3BN69t2sG9uhblqGYkCD5S8e/i0cTW9p+rxZCc5B8lTISRjMkDx8Nsa1t
W9rBJyA1LidseJLBcckTugg3Fa2Y/hXAiFv3zpY5DzG3a07YLspsRTLZXFGccNWnpXHwX9JrZUgS
KLRjwkG/1qGU70QJZbzIJjQUc/I+IVnX8KFbjuM/5OjELkLZ/RVmtmCljrEcx4Stv+9x4MgvYYB+
u7bpLIG8xRlDK3woPDvxuKQUFNVWP4qkKjowsG37YZ4edHjjLlyyC3mdlcjTz/uwmCcehzEtRGXX
KA1d4tfZs8fYTsKAC4eMBkm4ce2EcP28032nw7wVIpsVT9Eqnd3HKKh/sX4ycgNc8ZoXSkPOmiTt
TycYXFkLWl/wtF4FZImIdiek4ZlgSW/F95x3NpKmDivVGCkRSrcSNltTe0qhzoB0WgcaOBb/lEQt
iVob28fcE7uRpyC+Gb8WKAFB+3ku200ZFZvN3N0zCT7jzsHz6ts4+TzS+7ukn2pHUKTuTw3mnQ0A
QCQzGa/SHwRZIo7C17tCHvQJ4f98RM61AAG0pr9Q8ezVr8nI2iL9ud30dPYaCf6ZfHYHsBQvR8yN
Scxz7UrTSW5lnlIeD5pkrLHS21losqYy2/IWnaXCANX1+ff4BtyasNdeevSP+5cHs0ZJjxfidGok
+JTK3gnF0ejqBOFZADeGQUPAs4M4lJMws/j5CSGszStbIG6xJlsw56a7Z3M2AaD4vzFRJbibiP+i
JvsmFndzLlSIznQK1Bu0EoKPk4VaAQ4fPJMcNq90am2ev1eKBUsMPg1ZfAB993keahfzM/gcUbBY
pVnQu7ov+HxTRDhuO1sLcCUWwieL339COOqw4sYaOH3SNSaIFGECuvXXMFAOdJ+2b9s5kwNQRmLy
1gWEGeXAVYFEm38MElXfgEZFjBzhAEnp9r1ssAPZTdxI9sG22c0WpwUmVaK75XsBFCt8epC4QOXZ
JZzHtQNpR09mlkTQuLLIoqL/LXLZs9fpruN6xr14ccQ1J4VqnwOGDOZuD11hurZls6zN+FLsPHZU
VSQMHdkz1AEJbHsLfsEwolvuyW+NyT5IddqQly/sSmnYVf54CmUL1s3toqyWE8qMaGQ1/xwLZWed
vWc+PtnFyBBT/9hAgHyvsuUfPB/hg8vvWHCUK1yrF6EauTltbbsgWOm0BCnOPMKCkc3/vpQzLAVW
JDIOEinhPvE/VkQIW3FimaBiIWcJgFZNwMMBXHg7lzY84X5O6OHP9ZGXPRY5ctpvL5OFyyvuLHCn
dSPPW810NWsY43fPAqgcW5UvbTzNJealI6+VJqUjE3Xu/s952LVXZtLHFCY1ztWKYUy5nL7Ai57H
weDOAu+6x1nn4bo32LvhnDRaxsFdo+BvBaoL2UryPgy+Benntz1mXHCKG67c3S0NxzICbUIMzh0c
t5LIBlwqG7Q6Eei+4m9xYqdcCSVwujm7vDa2bE58/0d5Nk895/EbEmbwl2z4RZomPBR+1mGO/Rgw
DzV+WtaE4IHn7OyQSLgsPc2xGWOcSAaR6XCmBzC3H4Cnz0f2Mfq4bRpASUHPRynlxuhge3XxFHT9
vOUrtBryUAluSV7tIAp+i9xp70wkvyRGzzO3mnqubb+6FhWGAvMjRyKAXEBKJTZvHce8HdmokR07
Nn0YW0d83YblfWOqX9+UgvVuCRZMQYkPJXMaeLXslm/pwQrhAuInUso+5B1rxzZEY8nbERCr/b1L
LIxLYHjcWcFWEBQUoXGP+9H/2jkoq6G4h39Yg1D4Icgojbx7Wr0acWYXzbeHDMO1maiPS8PYl2ug
5/NTqNz+bbOyKO/+uSqaqUZ0kqzyudKVB/5BNdcVdJ3lpElGlqEg59lfLCPttDF2iIaaaqbvtXBg
QlgXY844r5QDd3Fix5TrrTr3QDKksvUjRWafpw8nwzhsNTgRHRkxf3UoOO99+oS0J6MBr5nHwM2P
2NnINV1ZV1Sfx90EtTNq/MDw+8yL0UwnUmEwx6Jxhc5mekWRbkHbyUAdZBQes5lBB4nOG04/NuTS
DaBqHN4KvW4j8egn8aY6trNSYR33Wo/VlSxayLvb7w5teISUr7awrjlECHPiV4g8DibrGM9YVPOr
bs8PCjguHyCsOca7g6p0LbB6h4rpkcmBiPPa8XqEXrHjHYHFcNjcUz5TaeqjciBf5eZLXOf4dYi6
7UXa2wQcqCcHCqUl8G1lRPmVqs6FpQshkxiqwg4DtzVx5sa8p8P7qhhiyS0HwuAGhOHhb4xLfu4+
AUL6omMSvlX2PyV8neY2YtAXmiWeAPicR6RQoFPI0mHqkYVGWjEbrnsTEwos7oduB0kSm1O4nfy1
erCartGvYILmQPdnTmn6lrRn+avydRJAAXCW5H5xP8dNPBtJvEFDTlyR0xSFMNLiHUp84XyrZ53E
6nsopX5h+suFJdAv7ze72iwhlVw6iKGgXYbQLFn40SYseUxCZewUSfDjBbYHmU9SOL+jZDMVAwqs
JURUZTB/XKsT4aK7OzA8DkpFnmLXO+2LEvF4zqWy6S4pVT4vQOh/pFMmyYesi13nnOhVmgII8yzt
uJKb+1P3cDkWYAlcds4zUsN+dzYcG4vGGEzcv16wIeT/4tiidEQ6TENi03fQk4zqcUebQYlOf8Fq
GhQu+pOPkZwCCZieM5AzC+Bz+0oe165+f+6kR1nerF0rbsTTGz0pRkK2XJ7BjmgRDyLv1u23zoff
jjIRjx8GeK3ZBcYU/IHrgsPt5v4lFut6Ffgu6c6dSupQOtOF6oJy/OL1D5iVizLJIx8cS9kmubfP
9gmJTDe6RlKYc1rE5D5CMmFvwM0ymjK3VDPa/OJAY5CeErRWnn5k3jMCf7y+2+lrcrkui4MpmdSj
nUJChOuW8TdUwhj0DvFZ8krK2t6/pe2TthD2EzHWciMnNJG6/brYR0oMTBsTDrX5MrUEcnztfATX
HiIDrp64JTjzZL6uo+IL4yihA03mCnsOwjA4qcyyJx4wfCZEU6s3qu2wfexoxkyGDnbNZg9dD999
6v/2ZLkN2nCDdrC9YY4XhBgN2J6slEiXa9yEky7BCmtVlZtk2dTEZ5DHpl3+VxKffxtrhGOKEKxu
1z7mL12k53DpO69zqiWVhjXEtlG15fMyUz+gMTo2lUFceKy7vke04YGiCW0VStY2tF9kJ6GZqCRl
AHw/w8xOurf8eLY68bS60R702mGo004tZp7/QJfhP2PKecTjPln7lXk7l3rhjiowDTegoPo30v3x
FcXd9S7zKXGCteGx3yYLbifbvZXGGb86pl83OPbUfSBM
`pragma protect end_protected
