// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
C47B2UNjcjeW/qBeCcK0PAdYaQ228JB79V2xY+HSQvC0H1n39p43Ln1oW0VcO9Ur3pDaGxm95BrK
Q599THAkM5TLISvSPGJeeJ9LaXPHzqiuwCa5vhAKcnBM+XjlhU1BwjE6TSGirc2439pGYB3+PMgt
2hPJSNMduu+7TIoraFkTqCdtODUm9gkvMioRrMaAQojKYB5dfWA9eAZGO53xFpPq+dt7Tkvs/drH
D/SnSguLVahTq0d1wQp+0drM7baS89Oqb96IY7SdxG4n5uYFwd8epptktPNKyP5hzV24oFTfKo1s
w26dOrlCiogb6tVqA+B2LQPvEUH0tkIwrhIwhQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
YqoMQfzICipNt0AX19AXN0CzM6MhZyW+yHVx2kdQnoAjmxAxG/GvW5qgCJ5/FrVkEvtByXke7Aqm
dHSlgYD09+fzlOtLN7F8yo45mCGYaBF+SsFQUYafR8YvFCc+elWa/euHY2fpquVwp12xT5rM9kLW
IRiYquKCpEBavcQHaZQUGE9awQAk4O/Ses68TpHZ/Gu7a3+zVPEowPhipUmBHALpnwtu51WMkRcp
qVi6StagQlMuRBsSCsBBkuHffY5odvpkLbFANbw5GkEEl9iTtM3F8fdBj/6rELJrUIs9G53Q8N/Z
MViDnITejwNdL++nRXdBSriJXsCWEQs3GELVOQ2R+Pa/L645mUDpLHFA9aq+zPgsvfaBb6wOigTH
sDJYfvUZW6u5ZFokmBdCAiqV2mSaJW56mInFXulMrEhxSBrCoq97l3EspRFgHihPvEZkRcITIAPc
gbnq0mEBg8yq9zJU73NT5v4Zyk9ey+ytUJNzU5OdxAWA+N4ltX9Twd+4cwTWf4d0GEHMqZssezut
t1jm9S4GQkG7Tbt3CdJbP3JeRGNRyGKslZp5SLXKs5GRYFjSIEv8x0pvpwUKA2LgIfzMyc06EEkU
jkHnalg0UnQyoCJM6YVR5VzxG4GTFM5zQAznhS9x9vDMelWiYYkGgaxP3l7GhI1mV9sVsneiLRWU
5PukAFE1/Dz6sG9kdvL6/6SXUwO9ku4udzbVro94MbqtjFobwAO3cQ4V7y+5nm7QRXP3KXW2/Ct8
YiGn9em//wSFUgmFqtkGCl66D8i94wQ3LW9l3wbpJIVqYcKVDFxcZzkTcvciiHFC45LdAxwtW5ZC
zDUepI7aT0KKyAlHQmM/8yz9cV5hjMAhydSTq/hdZmLPdEm98MEuZpboXxE/2AYhSywvIzB5qsTs
D1ievdWJQ2rLcNG8WKNIMAxFWh2Dbt3qhR4Z0VaR4KnLAv1VJAThcu7Tf50DQ2Kb1BeDR/OF963c
YuG2k6AleFGi7Vhisq95bEtMvLiIL7MQp6VSot3XkFP2ZOy2+ogKN1U9PK/41AOGLjH7zdZMOsue
p0ThzT/88E7gv1PibqXpiz2PP9IiBCGXmn5AojYd7aWuPIeAnCNm2EiQXmqvoom6/vXInFboNx6r
mazFotmSjrEWMWwQTgskEU+UoH4ukIopFOBdIoV1ro0kZn5qIzzL8tapxtCrrfGCPOJmheZjtfS0
yQ3egkJIkG/R48Yn6JUJBoc94XhV4EnqQ0zPTKpVnlWa2zqfQliZI5E42IYpaZXmo79oSC8WOm7B
1h2qfF8vj+A1feXk4VvBEJaAnLOuVReHpZECm2WTWKHpeSb0HV38zegQ+SDRPiaM0jFDpKuW5I4S
/xG8Pyiohf/I0h75fBer+RG+nmPnpCJcceAoK4viFm97gL0iTGxDr0Hg0JhnuBvdoAZG0Od6PQ1N
p53mC47t/HZEWyrVcVlsMqlc3/y+7BqRnWaHGCtG7iDW20vtI36skgd9lGG8oe3Ulkg91Exhiih1
zF7Fpm2AHzWQlkeV6jfISQ5VL2JnP2zWcHeTqhS7Ck7B8snkik1auFbCCl+YdAH6CH0xqmCdFxG0
rSO6XFB8Wo4UQXzmRn1W3yu31Jn8yJ0ltxWKdlBwgGkOx2kQ39ZihDlXa27NwVmicYCWIIv1xhso
iyziaxc5Tc3iUke5aFmfEd/cWQ9gC+YoBU+bXbjLTM/l/udVHBZPoofmQ7XI1kWXBPf1cb6iSDGf
C+kZLbaToPK/WtPTWoR5izzJE414O/AZCwUJb7/fOK6pALhK+QiFtAmmMDYVjo45rzY1PSslxaie
nvcW2Otk5Rju9dm9Pse5H0XffwhSIwGwrY0RddTENk1EOxqKiQguoH5cajK0jG4VyWqvTPw53qTu
E4I1fQoTtp4fDoGVbb0+Tpsh4sxPm3j9x/hPwR/D0Ru84KzK5AO4LfaRAqUHS9KfeZLY1U+xlY85
wtvIFVFOhJUd9Z0/4prRamhXkk5Lb77qhNYQ8dgzTQsFlxp8s5Idg89KfkbSZSJAumzsmJ1JLuUv
GBkCbSp1RsTYkNT2S1LFPFqYZC5lDXuBcovQsfzUBLPgBYlsjVtBzqE3AyEN9Jl7xBoFJgWd5p1H
5qHloDVrnPZik8hDB+qBCUQPwiI2nZgJvpa6mivHJh0mnDdYn06aCY2L6jId/ybhwLq7+q5x6y0Y
nhYmbQ1hUOiOkOw2Q8fgzb8cRHXqbbv+80MG8mlnvuWvtozihv9ATRP/RUvJydUmaGYinveWAfJ7
OfBIlK5ya+NPN80J1CvoBZiRKu50HoGTaNks6kjfSSXXaLMyVunSMbcGoERarS0ieX4/iEcZ7deC
B0d9F7+OBxcqEMDjHRPL3QpRYCGeUxS+4qCjiiCFbKBQ4IUqgIjvxJksc5ioA2ItOti/yIA8gz+L
/l4m/NIx55kMRGjrb0ZAAaLRKdTDAuIJJl3fPV3kGWYxFneZ5TSm3nhDH3PExmiMZnTHKe1zFm+t
PycoSeDsVxRM3ocGe6OfrxyV8hRhroLJFsTfz7UBntTDBgi4fo8dqdHalIC+D088E5bbl/gRVdV9
WQb/3MO6bczR1eAMok55zMTqy/eM3bk6E0JxIqaGUbLCjCefR/tf971VjYeW2mhKc06fIIuS9T8S
asTt9huz+QHEOsHpHx7Mws+MVMVCtabhf6mavJvOhU9+NYBrKE27VQHvJ5yJyzI3dmJBWQqqqLSI
n8w46bS5Hdi2cA/8lmuI44EbSkil/iQMhUrZvZKUgvaMqouXD9yjUtWyB4xKemtQNatuXx3ZgoMl
KwRybiKvZOlgTU90pVU2Kj8w6cvYrYg8sfmJWAVf+6g7ZRMKToNI5nlemD0BKJzJPChFl9RjhQQB
z+Ah/dKOts0ZEFBhvsBA9w+r35YcVwvWRWeh5PI/5CxRdm45JSCErkeUEOTYXmmJfPY/6Oama3ku
hzzYoiK2lTE3k1Om/QuVFyEKMYs1SPX4kbf9geBwyOicJQ2Goh9MlhCBHsjvWHNtAQn8CpuOsd00
BTXMpUkwmra+81Afi8mbxNmuqZE1/FCZyZxtuZp45ng51iyrgBv2G1UKL4KsfoFi7lxNaURjaxxD
NqLpq8P0CbVBge53FLmrSFSsU2YWItaxur+5VFSVWHupwZKAhaMYa/H17yR2AQQHFt/ZUn75SxNU
T22O7ZU/2+TIXJ9ikOqXuZTJKf1ZlJqm4xal1LVCeH7TPz84DkC5DcrH1OaGRyIV0B7iAwaCBOqQ
4gTrnWC7kTBDG4xoaUP8kxrNXmib2IJfYBodvjHCT2SfOGANqa3tNLf8C5G+lOeSBgApANd4ylpV
eXuYzjU1PTrW0Sp2L+ZXtLgisXpYu9cZ51nbETSsbZLLv+2R0vkbI2BiJiGPkTrrj90BBgCISGcQ
J9Xboz7sTOwpxJc6O/MgNHsjgUI9vAMtFvVWDLCd+RbcGhnQH7B+NeA+UImJiOpooxZwOBTpmdUV
PZBLfuFgZwFvh0kIw0FuM9NSLYPIRQvYJPjKAnE5WyctcnG7d66TSy47TzQKlQHsYEvJ8KsInRJX
NfbF0+pNl90rsq/oZnMQdHxtXhQAeKlD7zr2rcE92pyIB0dbMoeSJfCjpG61Wx4GpFGJbtWmQ9yU
K6UHl5gyBax8xRBCNaiAtQTAUv9+AksC5V4URY0qI17Dp0quepUn6F1V8V7WsspxkODqtwMGXeiG
3QjBbTv8GtZqKwCmaHiGW/8UQMb94cLl+bEW9wPq750KtSysUuJZUA0O5eW1IUmSK7vlBBdm5ndB
JVs1iIRpBhve/2iIVSwo/9LFTMfeLbe7D9s+xIhJoLgwhz77A5XJQx8EJKEZDSto5NGedS5Vlaiy
WcuzwxwRd+lAwmDsmyrNUiObumL0OVr5lSR/zWsMIifuURISjlxJTQoyqtrrm/S9D/DqyeUDv1KZ
ZvMANZ3bfd/Haljgh6WFQp6Zi98SnJZCtqGMWPTyVcGsJfRw+CrDM4YyfzVLtRRYXcldLCQNbxtv
lGHFyyP6PXhsdpBKxtTDN+BCQUAhyXIXYBBkpqkm+8FBTT9w2fL21e2QG/5Kq/rk59X09LIZHHYG
qALbkvydUnZ1HWxIxW9GhLW5koalQaMRkst1VW9CxXi+ELXBvmKQ/nbrZwUnJY77WTYhLGHsyc8b
XrLmBA2lkrKLbmyLZFzZL8zZOJs6+KBS10pk6RXAXgxFtbq0GepXSEjMEeO1VvkzSQaievLxMyvq
dG7guR3DBWkg3ZTx80v4KEn+p5UeFiYoQjYrSNmypITcJ1r5wRnZGxeOmdIFwd5RCApjthY4frcq
bKRjI/RD25O0EwxWOaORwA5PKIV0SSY5gEwxDE+C+oxuBt/Ph72Z0bEbEA1wSSYjLwPCt3Xp6zvI
pwtVUAlgfqNtZ9QjLOg187ETsF4O66C4oE6MjBsL84VnXh5LzourXoOdiK/ylfqWtNINn60guiTy
RSSYmO+tBgiLPVBz2cS/OLqiEeSNEC23IDxTz5uen7C4WIeCSHxkzkYp18eqrsScOrz8n7CtbpkE
u4a897vsDgpkRVY7LSxxSCJkeXiCTwP2aU714tvhgaBIgtD5QFtfew8JPbHR3Pq7JLi63pz6VFG4
r6/VRkTKFbhlMPV7QTU7bE/C16YJ7bg1XXpds94EGysLf6x+Kj7s3U/2257o3ZxK2rdqe/UNuq/X
yh5n/etlUKS2UP/6fqZMAplHhNZfwp7FJQiHpwjB86P6MXgBjAjpkFmgPZoJ14qdBtrLzzVhS5t2
i3ji0Go8ynOGFiYrQFUqOeFsR/hQm8VK626IoKLTZFjscCA+fEDx1egUITnUgT/4ZXjF+0fyeC8V
SknE9iW4zDB7y5D6v8Bw4PeKeRIAYKfU6aHCvraVN5Dol7wCaVHxgqFnG46IGqf3RY0PdI9mJsR9
vUJRpdWDF3LxwjQ5CCgfjeh0AaorpDzdVOmhmE16E+AtkpvvrRFqcnWp+8G9Bl5OvNtMFT89p27B
s70gO4wWtw1Cf0mBt4LK3RTDj/fjQecFILTS2pY+sEixFzncSmTfC1KZc+JL6U7FaGJmlM4km3UT
xGVdGAljlDv31DBJLB+tfTVdA5/klxVfh8NAfxcHtatJ2qauJ7OMMU7lpEqkjHtLC2VDWNj2RBJ1
xDLNvsFGjmgm1rsEcptxVfTFcTpAosrimdXk/BapecbTFXxk+6rRkCB0jGmH9r/aeW2Vp8IIWTCp
pNLG5GPg0CVHXDkLt7UNQdcBCBDBLPg00BlPlN5hRy7irlRO0KxyHr7AosdLzTq7nhKWGvSxEaYk
LJHeX1jcRTrJuYpFXYacrqtu88SMk5k/6EXMc3tx3wTEsMnkoB1BwTWll57L6X21oxrhakt0Gtrm
w1M6wog+KiC2ND7qNCABHA1knGgC1JQGcssmm5UXa7Fs4cBQpncNZp6pZ03YiWuQrQbz/xRB6NGM
zXQ1rBMwU1sOXXN2Fqw9pHLBElVbT6aGeRD8vjND5YvZbbSbIIpoKLJJE1q5dyfJt20cKsoRbIZJ
z8m7b2wMRTbeHS2PRK8HCBsrqtkFWieJyARfmCqW6KRbVtoNJCJBU4Bnw9huKR1Y0atgK+wTJ1/T
FCBvkYQokQNYKefZM1tj2wy6wq4BvoKXlOPLNj8EnFC3Q/o1OD9+JvphBKQOEhIVcgZ6V26ljXFc
UBXvJSvsuoB2xomM29oCCmUDe6W1jWoj9YXu8C4eHRFwSrKDBZlp+3sh/uWIk8ySIkQJRD0sQHNR
XfWd28eP8/l/HnVWZ1KwLYtkFgeUFWoJLYlcXLNcy9N/AXOPyQkGgOIIaGUxd/E3wyNkt/zVJh6x
cvdcp+3FC5IxmvOCISQziEZKa9Qn+KgP7mnXHwxJbLaS5yJ9vBbfJwqE+QKjUfUDzNC8RmfK0+ue
MPFOeGJRfBgZEaO8afgNvICio/RyONHjLA86aMzPS1mGvkfEmcQIuEwp3zkBalwef9Z/o+YjxtF7
F24y/0oxIj9Nvs7HmoWyjQnfnv9alHrUaX8J4vsUHWhr5sqX2J+NZswQaDV28JjhCQn5c2OHvWAI
mB4I3tVbUFiqyDw5hI3KYVNF/S+01GdWwLyljMEKhJ75y9KiRimozwCCZ0i6xAPDMTlkYDAh8TlW
wjz5buLcefyDXe7+BzFiHMVDCRSt7LocPYrwPjD5eWq1i/OyNtw3ANn5/fIhqdq5St4PoBVJy15y
FZslF2y+LMzqjebn+0pcdjaxLwc1IYhsqcSZP4hVWVmSiGDDofj9qc4Rx5C0FVgPE87sr8sdkY/b
wPUtOvG6wnEIM01+ZqGlI7TcFMRm7hQnRLAsTZNixwvPcjZEt4PZktIjIudcECRH4aODUduZnrzo
whD91xQiHEgq+qw+/24xVScvCRxazyx3Z+Uo0wPnBuzLLqcsA5n7bQC1374mkooWPT59vYePcfsz
YwKoW25SUQ/SfF3O5wn8YDJQNMdu87jOQJqT0W5nWpYs06FI5Wd/hA2IdmYUzDWTn8sXJalj4U8A
aEooFOe44V8w1rYBt2EwXptXwF41a20n0WvoNiRylB39Ti1SQ+M6smtE0wETAz4wFeuotzNPRM3m
5/J9ws/gIcl/mzZa4sgQjNZu3vD7rwmNpHazPHFvDKr/Y3I0A3fR3dfRbqBo0sADeQMMGDEWQNjJ
tL8kS9wDZIpFvM0JdKKFsh7qgMcxk1vPVIiXiDCpQpUUuRcPG4pkXl9zX281sFpkl9K5vATR09rY
D/Fd9kMAchnSKIrhOgvuapn4sRfwEtAa17L8dsnSdq6ZHZ9gRY7c0yh2aK50Aw0CprO+fCK46ooF
oiuUeUfNufAX0Q4CsSdvEndRhszzwshb/JurEdKTdeFxNmgbRIV2sCIrQ5IoHuJtjj26SwAwDblY
fGWMzDgjDTH2vAUUThrcnG+tk1+KubVHqkFlYCuKyPQXlS1T18e684/Y7zpO5nOuo2L/9uHkXj8O
FJFpsUuJFG/e/7fXG2JJQjQ1cDIIUZgrWnogb85agiJcvb1UdGV/d47ywzi46P7zkmY56vcP0KgE
EIyFwJ5ZUdAzPUDyvZUB5KFCwuhsU0jjmfC7RnxB2vJf4x1uHxFOfVgDI4cJEkGoD3xNV4hCtQwy
cZOGYdbKRI7i7KUPia5ZAN/CUFgqD6rIkzACPdbggXY3hDLAjQ1ps0JZdwiLBCw9CXzBrmtn58xk
cTwB7GGIvORggareGpKLADHn3mb5qSvuoBuB71M0KJvC/Ntaw58/ha8Qco3iqlDHKapFlpKPH6Vn
IbEmhfq4xPGPchaASCMWpcYEJn5A/vhgjyTpe2kvPAU3o8oI38llj12Ynl48VtiTLoCywnnao2Kk
x1Qi507Ep2Vb0aP8rG6QdM2oVYO4hY6hBq4tUOK20jO8tv8bRCEUbKBrLnxaCt7HVHqGI3QwxQA3
KtY3n/6myvnX9luDzZVt8MK47UBUFYyrh32QuxVcXOGFgDnXRaIgEpN9sOEEUasItRzUN8trK981
Nf0v+ncwD4wsbKfbroNUepas6Iu2XDt6L/qwM8A9ak9IEZi4r4kGqJrVaEIlpQYLXT0z6MD/oyiA
ZfHBdIgh8jkGTfLMRf+GDPmCSvM/WeeSxXnMrM6hoUqPKGDJMDRzTawyKM0veRUMMr+YU5b1cxGM
Qi8gKGw6CzxGdPBxugdY8xRVX17yxsbLDZPDEcDJlBhxW40yLufv9NSuqF+1ZNv5XZkSBXrY+bay
+RNaOzWBn4P7Fvy3+4Fnow/y5mOjyjDC8C/h2V/u5VpT8eBEwA+8/elTluPY7+S3q+lkD9SWs0M1
u7AwMVE6hwiadWaUDysrdCiZod6iMp23swUPETtRoVFblNUg32Nuo6Nb+5TGWqiT/T+Tyz9ckSea
YO2mPA3VMfSboAp7+hEmOgCevqtDZysSmBkwwHXWM/1hvXvX03cKl1sgk2uphdyMcx7aMaMHjkxF
SSydP4ANuJxeNuLpamdItziP+cN+VTLuP57AvlP+ygbu7CvLhOht9gZWpFAc5wbByfFihEyzHts0
N522T2+klx+zgxgd6EO8rlTmXp9Yf8UEe1OVUpm00CGw7sK81THSUtGCpM/t0eGQ0TzqTHhCU/pP
ost3GJRExf5/rDDh24MQLrGYOZdZbVzpnTw6nnQqfKsZLRYdZndgTK0QcWpQ0xhARm/6OQ7yfc3t
AnpDHaFs+DvTD3AvS/uep3J7vAoESki7RQuI3xxCpsg4wVWU5Yokk6NlPLzm5vd7Cw5mG682WzUT
FcGylSNQFB8Av/jTb9BRp09qF0RlTNVzPylZenqEny1UZIJEMegWjtkZZXwH632vh3yUn8EJurDo
sof7hE7cOU7kFMR7f9snqui1x5aCac/ieHHLwseVBkfakPJLRsGy8VOd5j2I5owL68AeSaGEiVe1
GzZjHV3y6WKVM9XeslOwAsceFGnGDhdaR9QIdB5h8eIWU/Yfccn/XFbyIsnuO6J7Hiiw+mbKb8e7
rHd6fQWl8i/NbCHVWo/iMd1VGRG6Oj4RIKvCSA9LeYEFaVcFhNE7vNo8tE13+9NP4OTiIKfTkrTy
jaqBtpewryYNHWsRfMOjORqa/GylE8hcfH/Yr1ZFW0DrDScakLm1rzIb5f4/a1Fh0lEl65vNOasP
Ij98Edo87J6k3mMsq4xUIS14fpaRqW62bKjerKvgoNxzYqhtG71ZTVp/XEYmlKNveq0KHA/SDjOD
GCFJCu9hKU8a5QKBQpcbkN8RiNX4ERzOhLJ0oh263+kciQpVXd42/oQk1Zmy1dJTfTZcG0nyU+Lz
Lo+pPI97xgPZze0PfY3jkw9grBR76b1aemWuzqXEQf7TrLEj1PLJ1KttAqT0RmCd/XsNz4JjGx6/
0vjdALnLR+EzyRAo3ieW8BLz/aHtLK9QGxWxy1b+ABMvCJ52Ob4XxWZ9MoDNSgaJcGk/rrseCBEk
RNj0Yv/0cL+bw0iGop3ytCk27dVaUGZnJcgA4oOG1ZXl69zQursD0hjT0HPl6RqSNm4LvEiaW36q
JYyfqQyP2pUyPWNi3kbZKdDVxv1kBcPOoh3VYuww4fjo1iNG11vuaJy57/rXHH1qcyOaLqL/FTk0
Sc6GkCn+dwCSpekebY4TyoyCYp2CkG5V92gGtUTcWwGtx7yinr4APFilJ3zJVvQONqEbX8u2KC+L
uB1Md0P6OfSklNsDHYRcZ9vA1yn8QP3aqPNM1LoPbzpqrnM8vngJ1dXa81MiKl+USdKhoFjH8a/b
caSvUAVgcIyUItm/DuzWDkN7qZyCleMgj2oLAF/G1+KDtgLC2iUwn3fKhAE3/Lh8bTlB/QqOoT7+
A7YXUNdgisEgRKUTJhYnv87+gJKhQgDHH87zayiAdhEG1Xj8hTzIgPuMaXEb8Z71jPMCDsuLjHDD
IQA0kFGjndeyTnKMfivZjGf87573iv1yMn8g07ajLsngZLjb4ngekWA/9CXltH+IkZ1SRjTsZas9
FNqSecjerN2P6RyQQkORP4g0RBXbehWflhO8vd5NJVsB2b855WVrDNIVfodotbJDOFJh3Xu8rhOv
kcvSV3wIumdfiP8femM9AThFScJDSRP7YWnR8KEMs+NXJ9f7KzStTDI81hXxi+Ciu1ER4lld8ogf
cry88Dk3M/uxVsraha+HEZ+Wxjs/qIVMuyiYepjHFJYfDw47ktGDTMGsZwD2Z1RVC6BwLe8QFiXO
C6UH2j2fdMBBa5CG2WNqyyLfcjg3FvU1gWj0XLmAAx2iYtDmVZuUg2CRBIzNFPSwaA1EX2PJvkmq
geYZQVBmMEIEIJJas6sHLWlujWKZSz9QINaNQs4ikf15kIMztSTf69/oVrrtrru0bOi1X23gTmTY
tmANiUr6jt1T2VaEVRKWZ+cSmWl55+j24ZZfMkNMo7qOBcEISX9B9Jk/WAueDgCAhnbuPMkh9vnI
S9I+2cYyZR+eFj14N95wfWh50KZ+7VYOOP1xG2UFCWlRLeEY8qzjCsyQe+dcRmGlbgNb1wrKdDnH
VSIm78tnBT0VKckPH8+tqSoyCxL3TefLxxWqM6bMYjbiz+YUA2RXqdVPpLnYESELqOegRgMRh2Rd
n7xeKPP8UYkDUHcmP/QDj+4FxOUlwb/5SBOxKRK5lMZTXKxfGrKvY+owIew7dz2T5YZ6utjEKdNq
73ixZ5zUYmjW7pG9aCfx8k/zuFExBWiGeAL4Nv077QhZ70dfG615qlZmXwqW4V0hxAfvxLdpAuPv
nep4YICqUvGwlswvIl3varobfQg7iLJhtrUPund21VqB4zN+hCIYZ+Y/tKzpxeYz5/Kq2tNzPBVg
PR2hRWt8EgkZhMm3NEZq/TQMi0n+9ovWLPMTDXqzAqlR6zxTJDJNUfRBKYOnT/XLoJwGdAfvMVRd
sMFRRLufPpAfcgAVr+ssV5TH8Xl5lDRYPU5W5jKSVkmnoJZ6UVdIFkWtZ5KRjDDjeIPwPoP9BxF2
v77XNU75eqCg84xnpYMq1EVRjZQIRyHwZ4iMa221vtnE0tqDcHd8q5epL+H4ySLDIbMjEp3xnvJg
aCP73KtBna460wP1Q3nDUPYWWw792tHs5kLWLrb3BimopbXWnQFVHn2YHMZbIKBEBZKk2ra+GjpV
FwYn1Mup5cC2M0g9qiHOVtKq8G7NIThLQuKtqnzhODIaKb0YwwhvwrVALZtPArBAgB6bf0jg4YkM
41x3tFA76kYFopApS0se6KK1CyTmQa1GYuBh33dKLKGTEMgvvZg825jQY045tvWPNQjxu/NnD2bn
pnhBvagdKbrRXPH94SKYCCckVyCEGm1BSgg3n0OfR8xgOKNBmKpQV3I3IBtNWx89Uq6RJc1JPLVK
Pup6YTwqlhzZppVM3Mqu6n/PWYuT83wJx4/eoxSC10P+q6agtrWxionsFBQfLuhqIUZH8uqlZOYd
jfRg+hHJu66iXN3wwWeNY0rZGe98RnTLCEpej6vFyW2vUoFMZ9IeKjloCpUszW90/wWlm9VLY6Pt
9c9TlxaelM+YpJ+KoTqG6h7/+IOi/PkWlxoB3VbcfEQecKboRd1AZTdtriXgoXGnubaw7MIos8ia
XeSHggOA4NHR9fUEB5WQn2n7ck478huPMNvJwlrzUdBi+bh3XQMacCnmAqgMiW3hrdRNssh0ZhZ8
95B6UM/Zf3jyFStNDuRA5LZMcR6oMdb5edSfcOpy1VhjxDQN5ang2F7Yv5FbQbbLJhbgxBxJnr8x
ahdRv7T9QPcYbXohyordf0Dt2yvBi8gQe6rKfNUjljtIixsl1v/qg3xXlQyvlyQNiYMGdxYNyhA2
B+i/0kB/Pgifm0eIue2Bl+buxPJ7ExSc08t8e4Jha19W/LW8tSUj3DgJXH7o9zQZpKxQAr7tTN1Y
8f33W0Zeoup0bpYzY1ivzpJMMbwsAlyaEhH3daPKzQsdKkU6NABI3/i7llE2iw84kRqaHNU/AuhH
0mnKuP2jIld1uFmEKEzJ4tk4kONlFyiIhMvRZhMVz/ScZ/tzzVfxwM5TIOr0zVLxK/dhIPoRjZ6d
R1i9Db6c4GPjBV+RIifv5gfzPIig9LeWXvsofU8xo9QEot+I3O5XA+OIl3PaIdHnK6pb9LvhwXq8
wf/OLPJg+CC4Jpn/k0X7V2UM6gcVR3CXL/4nGVqdbeB7sxHm/uE4SbfxuHk20VMQYdTC+Hrl0bbB
UHejhCjT0zDrrxCpivMydS5ABxjjVrHrLR1R0McGe8aMP2fKCobccMVhyytx+TqFY4FiFJGOLtr6
3jxGxbaA138DDTWxK+Hhep+wImk283db1XUycNS+WgOa3icqrozpQZ6xjefBz7KlmcwKUXLzlb9k
TP885iw8VqeuVprhAqbEm8ToiuXLoc7UQ2lYFB5fUaTxcIl5vaDwp+VX7+GiUmgJQTXC+z2yrCZt
DjmT+jKpdSRLqNRy3CnqS6mgvJeUcqwa6AvXA1fASgBpzlPiYj73Ubi1MNvCLYeKsDTPDezE7bxA
Cqj4ExgXZUiSbI5XC/aLM99dVmyDU6On56yzqGdSXoGqpV6Q/Vih+qN6L7+A5Cf79UDmMInnnk3h
5aED5XhGqkvwY9yvA58v4p9aKhphq5fL9rfP6bBL+i5bxrV/uBy2Ts+eNThxAy9Gcib+zZw+7YEI
PY2IQjHFq96e+azuf1am3MjApkPS5m8w/ZkdAigRZ/yORCujMSwgoDzdsJAa++F5zvqBLyCPc0cN
5nxaWwWkdRCuvK+iihlQGST9APRmiKQ/u7BZ3Ocmp6plyCKT0Y6UqFXV4qFWv2udZ/pUeeWqLA4I
uqiPAD7uvk/z+Lfm4/zmRB6qhebJNh+8ak487p8/gOY6khqjyZRiR8kvqs1jIhGvao0LOC8GaW9p
G9dp0HVpVlhmr75p/WDdqPgqoRrSuajDYnHxQJqkHDAHwclqpAyDLYru5ZJLN+VU98fXtn5WT6cb
gcVfNFeTlnNgO0h9RzPbKMkOFPKg9imEJIGVe8dBjPsi6I4dg0vL/ti0j7YxQoNNZOCd/xw+8T2A
7UEVrKXz9cPyTd2tJH2he46XqcJ/aAG6Kczf4MjPwofwr5V2hTAWcSKm65crDT1rMo4b8BesE1D5
TYZUMxKLb2+nKvvdHboIDwKAk5v7ZpB233SO2EKVXE+Zzf3qx6R3XflKFjagrdkRv1qHlsPARABK
LPvHOzxUhPBNnPFXKSV3dwpKNFyLJASbCyZvlXXue4loaQ4pxka5Tz+E+qXeL/LYmo1zXCyC7evt
BVv7MbHKdqB2WySWuDjSMDy/lcGhKGDPVKnjAeOQalYz3+ZEZ7W6B1juR6Ll0DOqrOuQ+HYmVtUj
QoprKRC2Rst3os5EZ6cwWVkXk+f9dGB2N8Ee1njMDb3eqCcWfnP+JD6dF9jOreGGGw+WiiY9GQpr
dBr8myw86uUkrqT04HvXrDpbBTWVdc09Wt7W+iroVNfoYSZ8XiLtYvbSaOPGj9wuFWXrZgC1Mztr
9x03cANgCw/0sUbmfZDGtuxE3tK/m/nW9TSIZ6Bbl41M9r0UjwOfSlAI0mRDNGZ9tqKgzBZTaD3s
8V7+FtqnnEMIdsqGLFAYYM8En00CLy5ik47BXo+IEIbiOeO4inKmNQSiTEEpcLaCKdiFOrqs3Ej5
/Psu6pSoFKDQ4Epq3+arQyf+ePEtybU83ghcVTl3UvOhkSDSxnX6JmDaL33wrUAhChB1idIPK602
fi+4Y4EV4GnSQIEH1i6hprFi3MCDdhFPOnmzP7UGGOrzsCsDgcjVPYN3dbG82E1Tx+hKifXFRpGe
lMELFRxpXGOURWsZpYqkoLHaBzv1UMtU9jWbuKL6RlvfGgeMxSr3Qoj7KYm4vvSXNXTOAAeJMQN6
u8xmLjhMw9dbTtSnDadWqep3D+3NV/lxkN2RZEAfiHC/jiqV9zfU7bGk7gGLiPGI7JFMXvROjVYH
LmGUhCVm/rSPboe+c8SE+8aCOoV6fN41aJhZSPY10R+aEXG8DTrhP+xD10cdBTY/ZtUrU5ge32Yt
twuir9OmEP+CludByMTO+uyLTnoZE/lsDuv/o23KMpU+8FdJbzXZ8UYMCrU+StVZQZuICO6skhPN
CTiBPK65QtJBd4oR0EQ44+FWZ4Ezm/Np9G7N/EQq/Jrqp1lJ2q3StdeEjJEQnkZqXKx6XUEwEzxp
rOozIzfPiE2vulS5eA1s72I5tz4abwjra+HlFYKtcutzhZrp9T0Y8XYc+8hrzzPrRxHlYd9isp1g
dZaXTV+Kfwr/pk9QoB61dVz11seD8IvmdRkJjUs/JN2L5supXlBXWAuEmDYyfySBiHnj0sqI676B
xGq4qmFFruRx3Y6jjTvGEdSZWLlYQ8LARpfgmlcnxoQMEzrdgpF3i9tx4zAl6RPMM1Xzi7Y1LStc
CcqTBPuyeCPHwGp7WmPvjdgNcAdvHm5smwt9gAhkNE/RXYRzvWDQDi37PUKcg6cVBc5fbGZGAhvf
LgsQ+sM7Eu7iJAlFaZM/LDbneRnlSnYThcbF82OVfTUgROXh2DKaqsqw8fTiiw0AxTDJK6vtLmsM
3OgyWaUHO37t9BoORoNYFjK5Ty7fdazkRkraWG8dS7z58UHMJLqGjp+Fd9S87wwjQ8e5n69BfaTB
MPNTuDHB/K5X4XzWMO094S8qLiTa4hFAH+YJRJaw5XmffgqW6lHq6nFBrRq+BIymglEBVTrk+yyr
WxlqseAwNIyjaPJoqDumNvtqRCZRnoVmfeRnZhyK466npeDdCO1sEmZ2hdtSnPyiDWXc7BWAxO8L
5MofR2O+H8IQbotassPeSpb6PXUfvjfdhJw3THpQeBkrC+JG/wQI9huImFcxAGMuQoZyOCQB21De
w5KcShpmmHOazPbIZCn1JuDBbMG6aypbxn5XxRbPNoJSlob3WKFj6ldIE9UZSyOtN4Sajvblv3HN
dgwyY1J0Y8UrSGErsPDEmA1WpvjrBxsh6ST+2R9AmzJibqw4QfAMuL6e9lvToB76PuD70WE+EBH9
0Rfh2pcC5c+fSYktLLLOdlHaN5+lJjcCpCxlLzIRe8uSZ+J/UjDY9kJtwPnuy/R0RPujJyG+eWYY
dpj79sG6ykjXu19UdmPFchnZNLKD4gwhx5LidLkyl9/pegHqGFzWPvP9KF7sx14CWf2VvACy2oS7
B+OTfaH/36BskojIAy3kH4YNBZNuvKctlfqlVfH80kmVogNoXJ/vP15vocfJT3XyIbw1FgALShDT
ocHX5fFKNP6t5RJcWQvG2d6RAso07dNSdw4TqK5SD1rk2DsZFGvUe0eLGm6oqhOMKOkLm4i6T2Of
MX1I2qz338sxNjmPMEPXTlV4ChaNLIjr/m5UE5qxsovSJwqKp+gtpYE3mlSfktuElbDQyqoKbxae
20Tgpd4h/73J5XGOh6h6cITDynk1QsH7owQ3Qn6XtZLtK2kI9z+Rb+PjfpIRckOFwWPLRgpFPoo1
3RV+Nb5tchyixL78FlSFADYRWA4aoRTOQ92tGoSUCOe8ahB8iNK1BfTSigDg/BMPAN7TOL30llpS
FwU0NbvEJVY/jEh2DZtXptx16CuzKK19b7naS2CIVKxtJH/hryFB39kpAX5sISGYLxnait+CdDyy
785S3c6WKQu1oVMNsjSxuu48mVbT4lMj9iIdgKjl+0X3O81lquKNazULh2lWJeVea5eEEuEkWU34
9RDWTkZ5EsekSF8ikoHBQ6cNOCfJOTOaZQw6bvf5HSgfg/5z5g5Ycbqsbju/DbSCAPovBAJoAXRA
YAABlHfktOLF7sWZWVyi0LMEH+R7GzPoSdmKslZDkJgvFR5Ij3ewH+xItlY5My9MOOV6BIIpPAxe
yM0A9m93X5CGcxbTJEQ7XLObuzanukuQXzJ1aOmouoTYAVivXLJ4dCj9+DspPoTsS16Xj1aGBl99
hIJ1byUQ4CU78+43EaqS9dRi573+n2qxM5YShWUMBSd9Pk/e1IApcWXg2fN7CjrUNWGxRITP3s97
UGl+dhskphHEW/cOeajd+wDzsYmN8rSE2xJWwcP9KU3xkJfrPSXV8iWYB/rJbOHgH0c93Jqu87dV
nxqHFk+hnYiBIikT5VHFVRZDROZ+/naGNNrAjyzIDA1QWiCUVD228k8eOfso4z3hZNzT0dLIUIVw
yOkC3tHEZTOyj+F0/yf9I0s8e84xG5RUO0hSEpomXLjP91VPO40vo+EjgV2744Cy1E46Hhinkdxh
qok31AhH+h367vpUtnqGmjAxSu4UZI9Fd3KcMgvpy0KYfDXfPTVf+XX1/BQqNxvFE9ZszMzypYUf
Pc/wHoKok4ha9in8TiEtjtHItcE3PFrxsBzqGn01eBb8ATHx/4qqBltZ7TBImKJKUQcf5JEoAHj6
rvkrBVdMkT0a0mlGwpHJh8AsF0kuc9Tl5/r1/OOLdSMjEEqHozu31Cy/+O0Sf4a2hyzGZZTbQ5NC
wLwXR/F8X3xOLO/s4QEL+kLaTqhojOc/PDl2CKZPBMht1ez1rBTwrZFDbZJ+sFEOjfnCwawKLrfQ
L1CMgzwjDYi7V0c+2UrzAnLxu9Wxcl7iXazIxio2+UTFHzrOTsjfri6/+y/VM9qp92Q2lgggE+9A
CbtPqhOP2cGY+M2LNnJuI3rjAdddVfLgyfy1kbTB77khI2yzG7tYaDzAlPJzBySEurgrVGIiVHTH
sPdmsG7uS3X9txymcBBw4raOrk+W78TL0yvJh1DkwNoK/9KqM3zFXeUKFCBB1BrqTpyo2+K2P6ot
ZUqLdsAfVbAe6vZdMYHtac/Sbe8hMBCTSHn3fof73xtWixAT8stPuY42XyD7EsUiaAn0Km0G3WmI
S73qwOzxI3xvHqRTDMOgCuPw1ycpoK0Ob8wb1WPSQckb7uHNFymIRyJp+uMerJHBhSH/FerPdwud
v39rAkMAUcmzxd8+VPtKGnpWqz9Y4XgqaDi2HmXvpWAQSwavl1hGrDJg0soYV/FbZ/JM2PmO2KK4
/1G2wEajWucO6spxix6QGkDtWCcxw5crwxz4FW8hVcl7uxHvovR7MMWlPAzBSnBLzWHxRS0m3Sh7
a2NUt1/ps/1X9jo4mhp8bM3iaP5G6tSODUJQ24juQzxxo3un+hlTEydEg00XLw6wO9+6F9616eaw
/R8VAdSilnp8tllazPQmZogPi1iQaj2LnAVxKrJ0Z/lSpeNczpITG/yp+QPxuf8ylU8PYRZUlCRy
cUFRBQsQOrHdZMz7YxBYhA/MKxV+OENvrO2wGKdQBRMzx0v5WStWpEXQkiuD8vekWVoPnd/2kKqj
+B52uUt572HQlEnAtyZ/muO1tE8HccMDYVcMx8EhTV6GofGpfIZ+bnjCUfqAN63h/oADWHYMuPhv
LrbTq1gSuTB4dfgIBZrWGF8CiFV4mPaeq18iUkwVdKbFz0cYxg0lkTA4k70sJ+0cGeXNbDNx8NKt
6mTXJxM9lsZIatRVVM28YBEg5nSSO/89CLu+s2xpEqN90wuWw7w68is4bGDMrbCuv1l0hyuYHOlp
m4mktBImUlIgZlR/8uQkRZAEYhh2iZrxeotyaU2y78CCNqaeJIgDC/yGcbjwl8VzfphNYw5sdH06
VJO74/aySs5+8tOtEQJymohavTht4W8h7CDTmrI2tcgmmw3tmdoFHlWN6JjWHONXk34Xe6ROyEIx
B6MFyhQzbTr/HfBC3z5UZvAL4cX2VwDIJNy1D3PO/VMfmdX5sBOiNJadMaBTUiV1AsQF9cZXPlqX
EQQXyRwmPbmbpo7S9cXVaxEkW8bHdMYV6Ox6+bQi4o3bqFS10uxT2uUXdLIJ17ihQ7HWNghPAXeF
3wO1Rc275OgbzVgn72nT05H97bNX/LjHmz182l+cxxX+PMj3L3ocpb+My9Gg9lqrhoeliIFBg9Y2
Db3uYib+FJhZM/Q/O5evyvfVBzsMwGZLUsX0stHO/0HcqkieinolC3u8X7wtoYemauFqEqdtZpwu
tulT7YAo+osEGoGX0Qlei7jQQ9PVIHo3Q3Qs/Tz6GnZsa4x6a5lIwamFdeXwkDmMkcLHRQFs6qGp
t4CgdSi2eSeFs4PNLH9iXzSeiPzUTKfWhgLDDlIaedhu7N7JDhKv/G/AOjqh0S2sNkECNPCd7sOp
bFLUy7/fQWD0hcQjFqkbFbUemBB4SFvBljw3CkvPZkOFqAYSJX9P22K0JICYSAou2xKqsnhsZMgJ
BaxCRDBObyrHwnOz4V67i/7NYlh2RgReJoYqZ4G+IwsIKjmbCrXe6/c0HXj51J2YKwYaxjQc1T89
4Y7/XjB1gmoXhAiKpaFvZEMZ9rkktsmsjcNhMTrlkP6sw7A+iub9ldQwaunrL6WcrBQVj3v8MgMJ
a6ywoafDSFVRD610nBX95oYuXcxd103/pGcUFzKSz4PGeZP5vemkGFFv+VYymL3f3/a3KfiT4S01
a1os1HBVAt2IzA+YdKurQ363hDUSAWEa6XsECOcOPT69WJWaBJIKX9cOlWoSGG4l66JwENZX9ylE
q+S314V5WG/cSwmi082BNjCIWxH4hlpx7tlr0tFKoMufCObzVsNSpL/oAms46PWuyhuAHni+PeMz
FJVxLTJNg4tDrZ3mts5lyCRuKbXXI/dr8x+I/D+T6712nVFv7LU3w2QVybQnnMLzvnklHOd0fa5M
LOzCWAtX8Pv7ZTiJWSyvAI5JCfLYzJdsjiC68SXiP76G3C1m6xIMrYmwWiIcGTWRIObi90cDFXbj
8NVd+VcseIrIfbrA6ZhDIYJvmPa3m1EZXP5UsoOiGcbtVI/5WRrKsPQr6a07qpgWC5glM4pCH9eP
THGvMp/fHWp0qXbFzda/2Dae04mJy/SQCLxjv9rDMeLl9Jctqbhtx54dHbp+3ddHFSz0q6wPbqG8
aJyUXtOZ7/kt6gevD1zZw4f040XGGudNT4B/ubPDXigjShwWjfS2RiMagZTDEfhCRVqTEsWHmzJh
SEiAd6HfiJZPDOAGmSd8aD2sdShUkeYr8jNv7+o48BPI6HMJ1qE6fjk2NQuwKSiAj7PwIQo1q8vD
Rk+KmlyidyhNu5/6HH4okFd2N2LjPRLrEOReBqj6q46YfGq92PJhddXIYt6v2JzQNe5l60rcPiW9
hzDrFTJnQpsmZWDPv4ERSDs0AXjnx1w/mYU6tDvEGQ8zJrSXLeQr6xcI6/7PMSXHUxyc4Vc7q+Ob
Dl7aS+GaWmeNMLeZLCT5nNdVOXJO+JtdG51q8Akx25NzPeB1Mknjhn2r/wGZiorYvMpBA3CGpEQ1
ERgg1iv/p1tcmHdJGMSeXtChHEmKEwVcukfpCFSNDClj6yrW2d9H9UmflRWhvydXjDV9ALPEKTub
kUmEyz7BXkzdPrMCA6psXL3tvLEfAvQLWgx2+GBXsjZ2T4Cn4e8GAmogtIldusdK9nD6fpZo1noC
KlGmk7eypCtP80mrKVM/ludvhXFCsR33gTzNZP/2HhjBvZbJc0Xvi7LZLiQ+TJpxUIFW8fHh5IL6
3dSKI/zRvaSDvaWtIgOc2kLtCKD03FGtJyPi5jwmNM/bM6h5dEq8mSHqRoypbzfGsfNfDnScN0HF
fy6Ej5Ii3KFZg2v9l4kAWpuwXXvUiG9Lnw2N/x0FKGVhiR6muutj8du0qe5MBu4DKn/wVOCEYn2e
kspVm6If8Xjlr/kLJxF7stMD8Gyv5tN+AaUTckS8It+3E+QVK6PqDDi9b15Zkh1P9iJgAFv3LTiA
mo7kEFx+6XwZryJ4y8ia50jt/cvhgrUcGoUwyP4O9PQJi6H6oBBOgB9+6G3BFTIQfOCgXGKny2/X
IRtlF73M1WqiOVd4GuEhqtCNM6F3IIvy6KI6VUnmskCPXL73WlKobdbvX4Fud4VzOPXhdBj/5Z5q
IdUmgIOIkydzjFCK6LafiBAAViKkHJv7j275SQtgWpTs7He9TZWVxMsz/gIeKsxV05YvKgHniKl1
f9aGevr9S5LA/kPo0UZojsWR3ijmak064mpFKuCe965e/hJ5bnr33khak7Q5zoDiinHrk/V4QcSf
1qpuaqJmXT7yxVTfFoHy/e5gCYel9tQ0bPiCcE9nftkT4G8qTUNP0zWVPtMJdqT7bjuf1fZhBwwM
4ORqx/G/onABw0gIquyo3tbYzJNQqJP7445CzEkyqIOHLxiKTDXuqkKhuASeexH0KFPDu8S7wv8U
XE9Bn451Anyzi5FeUpAPwscX8z2+c3SCl1MPJYYm+AsoFsjB7K7BSVZGHMDUX8mrC3pLesNIhsDc
Gdv4crtS2kOyoU9DX7muMhK52tISLKOVFyYYmzf1Pm3SaTEC6sHnNW8AmjLEBmX2GKpbC+L2rPa7
19YKr48jTXov8q4mTXjwK441WbqFspTrZVOrMGEPFFT0bthzgiEYu0rOLHfok+Nq1BMT5GbyRLGd
ngT8m0KCxWZWieMwi/wozF8Wl47c+DM45shNMK6OsgvTCmjjMkxCZK1t4ISP/qbsJRfVJwb07TQg
JAZBME2plsTjc7d8NalpJF9iHi4V31CMw30mtXb+a/iNRnS8Yp/iokwsjb8esrpylB4DomP8YYSi
MOURnO2xNF63X1A9MsBZ8VnjLtUOCLv94bgNiQIqgQrhXiMVKyPFa0AWqr5nQLpQDaDELPAyp6LU
iiIhtW+lwYauvPKALkmgl1ISaHEiixT/aMuocjmLD52qJ/DscjaiE7mnXwOxDO2mO3+8HlYB2TJ2
pyyD9QxKRxf/bDQJxaFiHkFb/pcXna450MCy7enRIlbbAHhe49lHnM5IHsYL81ypykRJk8GF3h8O
yMHHyljiZGBHqH0aZx1w9AUHlww7i9TK7Tz+5OOQOLOU2sfVAivYH3MW1t3CdOGU4js/lRaARlHo
Hf0bbZYcM3zDyjRmsh4r74+v64Zf1ybO47OuMI36V08GNj14diwQ81gihJkSZopAHfgFyEIDjTFX
FruP3wrTsPqSp3+TVbqVz4OcVfN9p1UNEpUQAKdSqPbanfljcGfZwsSxVmlt/r6tKZPwhYoBhxWH
1I2tU27kRV7DznueKCXWRNogAp2CwmtH752G9FNXJ1sRlL7XaerF/BblleaCkl+tx6gEtA7RIjS2
UEUdJFI35JoHv1oDAO3BsNuP1umHDo+t5+EVWnqOEvHQ6nmazGx3JAXnRQBtqILbDgo2VAjRUv50
xL8gPZOd7Nx5HPgwVy/0h8HlGbh5zcdZOA+9CXgzzKwe/QKy5FkG3XTDMY8EIHqdYyDCjp/wENTH
tOMuwS0TAv98rPGo16SsRCZv0RmZ8foNGI76iHEHxmNNfYZw+S9NcOdY9U0xNeQqD2GD+D1YXppP
qfL9MTOBB1S26HKAKLQLCGqDLRl8lpGjT9CWz7z4MTfo08Qj+V3wNcAoQjZffsmk30fYYLYDWwO5
ang0iRbZaD/h9XgSbycGxqgwEwA6leVJYtWC8S/ydjU7XPG/cMshcy5VRd2jCDh1HEc7223TP0Vu
XAcCi4zSpjoQArOxvNcZkU50JGSFMftjWl2Rotil804eIb0Yhkf2TAM9qcPA5t7/iUfAHcsG9adL
t03VmLMXlDTg1tDeXLABSConKs5MI3f5ndChz8o6Tpyke/6QI8xlyLUeB5lS1o1uVdQc2w6O/p4g
68uEg3/KI0DsADodq5cW7OmwnkvKLvRW/N0Wbd/Sd0oHDnI8ko2LNmqKK/32X9fkUK5kVbKsv3V/
Fp9k5/LCKovGIDNPyO9l9BlimLl+Gvz5D+xxrBq7pGQXbY8qi0S9aYpA25Uk56nob9hCun0CdNfi
XPxIrNvRkeV8FqmagatwNpj6kW3VjPetSMlFLtIEqCwh87F7Yi8KO/aVo0eM9SGFKG4eD/5SNd6M
qj6b529tsac+0AZGezBn7kJvJq5G5Of48aFgj5/DgbP5gpNU5lncwk6q0X0jdBEHrR+XBIrKQET6
moGm8Oo5Hd3KgnKTGTFtTRGFXVTAljWXM1+s0ikfDZ98pbx7ATauA2YVFRotEg3xwsHNBl/7oKdu
zB41PVa45CwtytoWveWcpj5DubElbfn8hEP8Lkmj2dBD58v7csm5uyurwd0/QSzp0hp7jE15YfnL
i646zz1aOviPabpOx03TfBrBHCTugGbsL9nC/dxf+g5yY7KxTW36kW5xNus9FmcwhlKdGVZXb6Nt
/sZ3cshqjIf7Y02W33ZEAP21MVM4dH3Xhz5GTtbU2P6NpyCYuBWJyl6ElfWWEPDgwzH0m5m9Vf9H
G2V7T2ZsUZNyjLDpy4h+pYsy+n/DLCLkmLTcJYGkhJNZX111nbtkF9vj3UXbBjZ1JpsNePlYVluS
8uMcdx5gqMnI3PZ7keRozWTV2Eue8l8wwfz/HiEcP8+P6LfANW/w8oe0DOh9DM4J04yUe82Jj/7F
DeSPfp+c2k7UH4gtF3xqAC4MHwPjgqGLaXkIG9Cty1pqOhQxKETuZcoLTDeGEjnCIIdcCuSwixp+
jHD0tj8Oibb/rCIJgkIZXpT7OoXtOjPKR8OIzd1GwWW/Y5dxYAw4HFjCB6QHtQMYgVggye/DWcqq
aSN1qo9xFyuOpbWoBlvbm34b787vJ8EIh3aPVJYhXTzrHKS8J+V0y9cF2n7/BI7/f5cki82bMUMv
3WgT7q9MazgXVIiZQSQjCvjF0lriy2NIJ3UBmT7eyTr+rTXc6VqaEWVCDGGDrD27wq587dOLKGnR
5SZTmBMI/HiQfdf2s1rMg3Q8Z917nQCm8hpQsfM7aBxiuCnV7XluhEU9ZeZGY0SWancSokmHNz5M
2P6gTDxbgdWTGZbZvTAAkG3EU6hJ0MIoYkcTpYzVoZhMCLBL3tCBZKfIPL0iq+o0Tokz+bdyWMFk
VlsP+X8DvulFTH5eznDOelrzsdB5x2bXki5tuZhqE7HDZEp59R/6BjnV7XrAOGELzhENCAW8aP+I
ZcAVfwDnziQXXZMC3nFjJDmPPdHuDpEyX+mxSlPaLDhVNnEEhAHwHB3nWOhF0BiOeF2OCWFlajzh
/7sGqar1h7RyBs1PsnP9Q1iflWkDqjR6Bc7Tgz1BVYb7KUAStc2UdngU6fNQ0N94dK0B0pZ+lt0V
r5NsgXANuvDWXvdoqStQJItTSbCqb/FohSaWbYvUolpPy/QIlHpRESWbwHYzGYpKuJIul9p/Sf2z
rKKSVBmlidpLoD3KcX+1XZnf3om/VHg973ikyGeGhv7XKQWZoEUmy/3MWLrC732DqqGG9Vmdf4lY
NiwveQmCwjoAwbNaUy/EDQ6jGUQcFn0O/XjbjbZqb1JFrov0DCn7gV9M0b/rBfPI/deTTHaneKGL
/nZRyfL8lMSGt/dPeBr2gjgrDw/+MgaY2bNaxxxZ/Q5cWr5WhSHXf4yol00W/yBzH3yQCT7Ix6jA
8zDaL4a2YCmQBvU7QFlYhcGBUhEefelJPGxwQ+VTxYLvJtnmYFL+bGuM0qHSiGPMyto7TEXbnGaE
jNelF7pZT/Bn0E8IvACUfTw/cLvByXFaXeYyu/8O1HMWJg5vzxXYA4Bk5iCPJfWOG/XRPLE5oIHk
FNDyQs6p53q+oImLAncZNzsRACQMlVkqx4xK6019pQIzKEo987XzPrMstunODW5nSYGQV+imN1TM
2wdeK9v7ntO7zB7uM/zr4W+2gRYjzh9oXWXmwHLViEt/hMIrCvW3XIQuwZkq/xcEr+OCt7TE6sPx
gLHDREOmqWgOdfWyNOwShDu77wDLWmDfoo2sulLL/Nnn2V5BzvhZGS3DSsJGT/Wb3EPbT15ppFyb
tOBGAvmEIcB6fyxASfRDoufVXzls8utcagdW8YBriCOM1YrhA2BeKH6NjA0FWk2xyNeiLo43x5Hp
wKXDQQ+rbawueW33bveUXQQO/qj7zOmnIQVmePT838hxIlxzOVgrOkN64RW+8JPZeT8nLGFo5EBt
76urqm+DIYJ5SeS6ug7GpCdFaZRoMjHE8YeidqtzUeGtj7oFl0G2K0W2BrzcETZJZOdkPknx8uit
ImYdMhnJk6IwGzjuc30dnYMMDZ7jena3ZMjcfVSspm7ZigPmdOjikVZ5etWHOz0vchzfdaNe05AR
x5XISHrRdROVbxbhs23ytrB9bNKi/wbl781Nj+D1JJSuDBHxE3C7ICZ2wWojgJ5C+HjW0ROmKKbp
MXb4F/WGqMASGaq4xahO13AlTW0aiIKr9t5B9S4zb1DEZ6/fWDYB+5zAbNGECh1diUV6NGdlNppp
Ip7EyrzDdjf0JtHyvlcyzCmbJovC1y+ZWZiEnSHqzGZmuj5VtWl02GT3N4obNkWSlx6tS0eTkfqH
1bAJLobOAMgSsk2BFanRT9ZyOw3PRZ2R4jYFURt6WO/S4anu4muDTo4BQ01XzdtC+/5IszIJfAjU
dYT6DhuKez2a11S+sYaZYiEgwzR9RIIaaFtiEhRo9kuUyRmMCjx28kifvKS8HTl0R4dKm6DzWDBq
V9Iq0GtMwFecaB1tDCDYhsWJbXqjUk6rcPCSIg+K3DX2FPuScWIk4zdROOMODlLGxMgsV0Ibu6Fv
0fLZpLkV0lRvmGy6IEw+xsTwiZhkGYW8ng5Otu7RRpcwi0JsRvvLfBNA38fiZF4AEth5ji0PyRT4
Xsb9loy+5iLO07UWqYL4Pg2mU+/Q2GLy7jmBCiwqjdpGA9KdKAIwDNrJicOgnAT8PIpVqmvj5JUI
vmWlTrX5L7j8U+e1+CsDn5/icHleZ7k0RX5sbhjjzh8bycgA0HOujDsmwOJ3UlbIm/mSA6DU1eEF
Nsl27JQoBYPxYOekx5EFwxYHLTZQIBvxcvKl6q3z2IIkaff/Wn4Q/x9ypFzW2xBrqbRG7GocjTfy
3+ve0yMV0vN9yzM8YkHRbhgrYXdmXioWv0a4ZSVfVZblLWxPx/KwpClJQzvRHsPOwnf9A+v7gZoP
AH5KQxwr/14XvcIuOjdVWIYdvS1jVpGhtgTXMoaakzUpfdoZbI6RoOddhQ6x5tB+QQQYxsOah8cA
uqEVQzgZOotlcYPyf2h2t6RHYySQZI4m4rV8mG0wNoWOKQNNcXV972cIo010y8bfinK5zOp2g1No
R8jv2KLzBgQugO/+kjw1KDgzD+lfqG9aaY77UaDQxBmrFuY7ckDX+lzRV05j7i7VZGjornjfJa/g
GpCZrlQFocKq3rW8uOxv5neo3NmN98hVPnL0TG6w9JZmPP61Oghxe6WKJlJ41bgu+UMLuo++0ZVD
/1TxDN5wnztC7NW38a5fPCoGgsemhyMnGMBj61bTmeeXeVEWhtiNuye23hSVjTMyJbgFLOimLn1x
ZknTfaAtGkPg0smhAvC/FkHU8XMw+JJ+2p8b2P7rmzv0mvVbzgTZUwE+tyY2GEH5UP6N6lO2a2Rr
xk8MAGh3b/NMTusYOjRoI84cVZIintTqBUFJMytkGkcOzJnTZscnW+SrIy3Mevh7TenPV9GJPXk7
UeKTqT/6YJ8l3aFjz22ZczbVBK+lMcpyah7bglqO4ZMGDGAzfGEjadx7PIbchS4yCf1epUXX2wBr
zRg9VAgOv3FsATO6DzlDrBEXDOBysE2sZBCxhs7sa8NogZnEbtCpaJaMLH9zqoCSMl1fsSp81QnO
gAZj+5QuFAIa2wuNcI7CFNFc4JrUXW4FLUOUlvZr/rG/6NDZDYRmV0TTZz2kafeBPOj6QmXdXyna
He9VZaOQdUNeSKyK6KWOVibsFbzOafr1KDU9Cj4HgF7HR9nuQin+nGegPpO3PbtNgcXlWPX12Tr6
meFJ12rH6WSYLCnhEKpNAWF9d0C2W0/Q7NKOKMjXJzTxCoApFJj5zhHGvNDcTAwiufdDnX3tptRT
7j+20Xdvl9YACEs+OA247pMyMXvY6Z+Qeq9SG38Km3L6mTaejJ5CPySYVAJx1qcYNA6xFVNK3dwu
x6OI170D+DNh/peOWkyNy5EmEHGa5d8QO3DKh1RdPgrM9YJfysW6qY0goMNtycm/5F9AlBlN63QE
zEWh/wX5S3B+MXPwRaCjbw010fWpO5kJVJh+BwrHuy9eMGOsFxD3glFMbptThl0rCQJSqxGkf2xJ
H5keqWFbmpaZIG9DRE0+A3Y9sE/OK8syfXgp25uXuRB4cj4j2RPrL0NId7otvH26YzZ/4GDE31sl
XQjPD2XHJQ1mqs1dpWC6hAizgZkZC/tuckuS6LoCAGU3rlHLXgRz2Aw8ckITRWSfneaN1p4wrx1y
ECTp928IEaRwqcboZuRnVbX36m7wptL5GIl6dkBr0FAAx+L/6FrEOxJudXHWHTIxRfSqP+wYVUmr
KFKgp4n0y/ZAxeogAJJWbY1Foh0c4c8qB0ncJwoored35pss81VXfHXZ69BTTSTwMwGwvTVRWWZ8
TryxZcH4mm96d6kEZuvorY9GJC7rDebQo0/xsfCo/3fLUeGUcii92CkFg/pcBeiDejXuJVtsaQTs
U92L9lLZH8Cm5jC9hbIBTWqvQUvRjrjp8mxyiYL7We37ElNOCaE3eOe5t2DlrJzk7j2uJfBprmTP
GtwLH+YWuN07EvdVt5T8/pE8iaCVo/3UcWIDU1/qf8z/H9zWbQFjjAHxtjFBwBe/mWRas3aiPmZj
HYvWUQvvNgjDYwfZkbo89GH/9ZfQFJBT45GbGz6vvehpEurbp0l1M82BZCTC/X9uZnSIPDqHiI7a
G4zkLfZmK8pNMo3K463TTNHnbMnBxSeETuvVr2FsWuszcjSoJ3xs0/ZNtQTUEEUI+yh0Mt8NOivw
rRxkGafyXOzesgUGWNE73geDiswVMohhDdg4zDROYruAFcqeKSHliDL3cn3fTmRRoxcJVNJx3BiU
c79ySzbX8e6pqjI4V+nkdDyIZms7t50lqzZzE287i0LY4FdOgmgHMGSe1cuZ3bjySo+c6ujKbzB1
vEI/zK2mf1hvYk5/sE9B+J6uN/VjouvwJMlxrLQ4kBns2ZqT8PXFKhD/dfQeNwkS8GRhJUbm52ow
SG5msTUk1gtoF0Wgf6pFrRI4AqHispxB+HR7kqYGNNN4PsSwOibzNfAzjENQPEQbvMGzfnD5IejL
bSpoqCWGh7IPk7mslgBcp4JpGpeGWgXjupANUJDT5wPr5neDnAN+9LZPpWjvLoyCUfgHQZCPs8jW
OFpy5HsBzqU0eYa6/+Ps/+QkIkH4CEPXISPgrchJ7VRsUOSJnHUd1i/+Y4CQaQ5KpTr8SP1TkPFC
5+8l/36HfHNMXptHfaoWgiHaNgc4jjl2lzTcoMQ690jC2oPbpE0Ee3vy03qp+Qqso/+G5LUdIGOm
rR1pf79tpeuAt6V1LVEkOqvrReYnbJn7kZXKWAaUuSM9QLX5AG8cr8lWa1jrOEXdBlT086g3Nbn4
T0AlI8Tjqdp9GB2d+n3OVbNj7pYs+TcxsDqA6v52OD4QP9e89uTHsbZgqgO7E3RUHgLMrPF8dzcd
5R+yUgZ223afY9KELvJd/HQeCA/1Us16kS0jYOZEC3q8RFylpfwJVuq5KlA+fcGXQOA4KQrnkveM
Rgv05hknT5kA+7A+AZvKxLC8p2+ZiEmRkcAlUmpwxlKR6eNNom6w9d082d05IgOysmKTsFdoTMW/
6SBjPWAbHaDCZsVO8NVVaTo12Og+U58fWkDyYiU2aAyCIaRdXkLVG21Hd+vXCAfRRlDBM0wfsyuK
XvxZntcCU/w6MipCmT4CU6JzRwrv+U8EEwHfReHFxEI2kPMFnvEJ77qAdi++6WRteKb9Kc+YGblK
h9WEQTI7sKEeJtv3ixoHf8iNMDr5K0SM7VQeOXlgvwpUihlpVLeZ1NznBR4oNwx1Zq6xfKX2of10
1xW3EznmXtc1z1ukZHn2VTX8I4LRk0FAYZ/Uc7ITh/Fld5dJ0EBo4ePqp3r5DipuwD6cjrCP+3RW
c6EAsH3Q1go0WXJHOHuYrXWH3tQT3vR9R31TQ4GaU4FdQUbttUL4FyN3uycz0GIykoT+KUnuGvf4
kvZVXSjKGxRgh02b0POyphGl5eQnO/h0jgFmAlbBKkwR8sum1BV0Zt7cEZsKS4HEuF6MTOgVLD0S
vcC/Gl+h5Vwkk2DXIN5PSTMfQ81LV8GQTjaOIkfUSbUuMw4dACoKYqK7SCSE9gg/oOiOoH1Vs6U2
Z/WgwMG0x1/9550pGM5PuRiViW9eAPAjVgPE6c7UpqRW6jKjh3BRi+cZyP4bTknBArmKiMM8upuT
kr+8LXkn0QRCebvuHYPgpTvSttNXVZ/ic5RV/FD961kBT94iIT2iPH+yy/MT3+cbYYh++lziBrab
ExTUsJYmJcb1Rfgq+dXTvlxtRBnoy03+A/TzOGbT/W+68v852zDrR20jp9XJOgsN0AwSFUHoy8kb
Oik7uFiNaVC2hYthplNzsN3t/p5wMEFF561HlbrINQOk+Sw2HX/s0B+k+cneWJmMHQN9ISFAhccF
q9+i5A4Evxk/U2mPxNHHwQvqXIpPsmDb42S84OIHoLQB15mUuHnIQTpH78MM0uPo3hxGlmgATBof
CKXJ3SOj+Dut0sElL00/sxWVMGb29SrYeEx7w2wgAFrN4Lyzxgfq04V5wwtC3tnnHCqxf0UeA6Ra
6Kl2a0Zh0HYN2A5G88+fa3p3U7y2kWJxDrBMLFCIytdh+WDjmCBxBRRrhgqXEo5WomUkcv4B79RR
1h9S0jzY5a8341hqZEsjQb3r2YV67opUJwPyBiriLlyVk+Cg81X5lkBkgqd1kUrdhpWUKhRF5JwM
HE6SmEFTsW08GCoC+Oe+H63g+Lk85rJ6gtd1JNG07kMc664qfbTFmHJNULmpkd4H24SaIZzbUDFs
geK8G4KJgidh3X0rguPP2jkc8urBPvJx69AVAqV2Fb7Bq9Lot36KoPRhGmM1yf/PGBHpXLD2J7Cj
fDAYX43sV3zs9xjgWQNl4HlWACtPV8UFESwCYvhXGnEWoD3QGZzITUWINbsV1MNmfdOe2GU9OCTV
5JeJ4oxtvXI0VogboY2YvY0LBI49UAN9NEu6/0xswQBMLR22iRsPT7GLFf6VJsqoJE9vh6WtW9u+
sVeWU2ZUXqNbZ193FGrAj28KFL4z8heSlihh95PL2WquxOq/ZjRn8O7fN7+21ypaGR7a+bxNRKz5
1xxO2IitJIr3hMFBfRbdpsc1pxuZQZNXUX3hfIqxirgdcbJ+ujI0JWprv7MgYRDYABhtV8YCawKo
BwWCvc90oGDITMzB6lbE/OOFOnv9Jduslzu6KmDEo7xv7/d4JoXEiwamX1OTNZY5KVQo98OMVh8+
4p+Q6JTVYTVMYj8yV+pWootdY9b6yney7MXOhxR56EgdkLMRtP4s6RujQhp7l0rAzkzMDJqvbGMW
jq9q5nCmnmp/qBAZikk4sxC+GN3jyfCP2pqJ5L+OMQIRZsfd7SF4Mc4Trauh4uuziduQiHsComq/
V63cQprEeG4AEd0uIrhbm6/MaUhzOSleBMLHnQeJcYpCIxTekuMjeZ5kLwzEg/qPQ8SC5BGkUAZN
MYh5EqAqMNs1dzZPxy3QitmXOOC1u2XItaQhZs6nsb9vvFrD6lOfKDxuQyvPNCZJI5R9/geoTEG5
kkqC7YCOqJYmXwowLQGw90NUbDZONPfp4Qra8KZj/Du23PdDdiCsN/quVwQuKrrPJlfFaFOL84oM
6GpsvYwE9k+SGG532+iE/9QFGcA7XbLjXglr9uTp5ClHdtwlW4G7z/xOQ+Gmj6c7uIe1q70HhIaI
7Ujds9pJi2/BWqA/eaMvWcVQB/tdmMvy9kCk0+IzTpygZ6ulKn4TPEgLsGEAvWqxy4G7oF+eaeId
7lSemYcNESqRLxu4d5OLtf3XvVi2vwbWNRiPQNcb6zlcuQyWAG82549TjZT+OZYUAdjBxLKC/qwJ
oJhPWfLVUoMkL7zJxMS6MqH+U7+kRbL4xjHFQgpZgjPoBYnnxFWxcyMIeAuncHb46uqzX+GpGIwp
yYgit7U0i4AMP5zf7QwfetAD7lWbR6g5BjO7H29vdtJZ+ArhLGMoLAIa/yVCF/MWN2qnx1KE86X0
lHXIg4xd4yXj8GY5MreXTAmB21pexCPH16NsXN5LOHJennFgGKHLLQOFUiRRaPNa3b9Fs72q6ouj
FQn3oYux/d9l0fc26sydaB5ChkRHA1R5z72SdJiqfft8Sfb8q4P+zzSdfFOc/9gwkkmEJAj9RWJz
J43/i8WcWpy6AeSS9Zj4qhR7ukoH+JQ9o/wEk3Y/0V2yjg25qw/LNLm4siZskDWAjDS8tEVkom1X
78L0VGGrRFagkQXLc2eUGkOH6hnCTcSUlBP8BmUHWEt5GIVASMDRYW7Olnq0TMFpI24G2mmV61lx
SREX8vwGC6+zZOf4UziJQECuaadg+9fZy06JL65PgVFt+prEZi0T31hThWPr2DKc2+fjdi3k13z7
EarZElQ//1ika6EemyvE6xrUw75vc7+wVBBU1QruhMvNe1tuKLE7plNC8D0+S9LZq3llo1FhDxKV
+QlRIZSye9LzmcgZ6NMF2BTPM+2atd8yngh+z1JE7SWGeGUcZlrabPPhJcD4IlLl2mhOsKFm6zZz
kz0hnSjRHplnIAjPhj0A/HkpTMS6parBjHjmh3TUBYZTqDl8RZ/z+R5U3QSc4wC1JSJl/eummCSl
jaykljYP1yptA9LZTqi6q4eJlSJvXUwwh4/VOfINigC1xZbJHwPcZcdl8LQiEQBNOMH9RDN9a0fm
pZcP4GqF3ucQd6k9DhCnmAPcA8TgC1jyVJ+SAVo/NnwOynvdNDC2Iq28U+LtXza3l9jzV6xGgtDK
slmM+BAnTnxDF9p6n4II3NHl+/UIE0sgcxbl1lJ2vkXNzqFPconOhIVLLUS8kgcRaxaKrZG/vVGj
pSRPON789eO+RNHvQdEJe8g+bRNfbKqLQHu+aEpN1JBN/bMHcQwJ9AvWwdv65xDfmaTI8v6VO31F
e9FiOCYRpL1A3BJF3ZcOeZXjzG/QotIJFcUzzD5cVgHiODYFmq5hRe3ILPUptS9oJYnu9o0hPapv
Mui8L5KzgDM1CxEQ3gPIUKWJ+pnyO4WJfuA7cbkffqAtedpGCryWzG+2Oab5HTJkCm4EwJn4eoYx
9Iiv3rFWViB8247MpGOsAKX8o95OZHuKduXslcmo+e9Y5skoSud3twlMFFQyIhYQpWl32Tqr56i9
cJnxQ5zekyxhH837YW9sy4mN/p4cz/wVYTv60Bz4GkPHBU0kvSUd6XXvMWSObQhh2rcSyjKkMCGM
M85ULGqZQKgAsJNeGX/mLUMTSW8JUIp6TBkLkftm6zhpjT2CG4Tx8qBCH4xU+6uQVAD2gEU9zK7B
JSde0UZlJIlUnYorNRbhNnDppxPIY8NMCXws7FobBtus9dVK3huUJPPglfdJQcj7f7ux2GH2BaVA
MxpV/mCt6PK5CkPElV5/zjtGNy0iRp2FnWIXI/Tqj0v9aQxqMoHSsR8iuxy5usxi7RNB3dP/uvJy
tRYJD8r8FSRr+kry0QbpZ+PoAjwRYrurd6IfVEQ+gJaR/8yykDVVk/v0UeMF3GrXeZBftUVMofhv
AkGr8aPmQyqJn1PNuLVt6yZWaScbsIokkTt7HDntEGpr4L6LjEpoFWATASPhNm3pWt/yw59kfuo6
DZn0EUwji1B4Y51Z+lE2cq/aDtv36NNRj6hIeU2nB1OkIqjN1PBxbrUYx4efscHdewBrhYT0+cpJ
GAjt7Bx70iC043Gyivz0MshjhhXdYI6KUuD/bOYY3Gt8K94I6JdJUTnPUPmnFrcdLO2XD07nXzYM
iOnqeXBfoaY07mYcNTw7KSzt3JZrm11Yez9ezJja5wcipBwBZHzjE5XnR6aiLm+oB4woG+R2zls9
uUQR2l95Q3XUJS5mW5Hk73e/XeCLBaEwaTmj0bFnjDriiaS9H5+ipoCPwtdkCDLOmBkgOl91RD+o
0Yc5cmjpGU5KsD5Wv+EiX1DU1+tDQCvVvPT12B/DjDIlxz1ATNjiMut47m3yYtmwcEX8/zlubvoA
t3/UFrngvQT16vg8ket/AK3Kj1PtV2T1VZLrmdd35stnp0GCE+4p5SVZb/b9XO9iqhb36ySbna7m
1gbvAYeP5juG+o6t+o7wYo6oppEDXkpEBelCQJZXrPEnYOgkEUikWZnbkL61vJncTo/EAuUb+Nqb
OgJQqOYh4kPESw/3ud6sJBIBuVOKWrerZ7E7VI3sNYidg5BZXgoHnKkzw+oBq3avOWClrVKU475u
pkHtt09ixl741NSK7Z2zgGfYbaOwBSFpOcnUCPi2sPHHhv44gSzesTXppnYpPTdOAhO/BG0/1bHQ
7tPsz3FoomZi2DFY3367AFIxMmCOq+9zpf7gDxeQUGvC1Tb4eP09z3TUL45x0Jwadz8sLOBVXvx/
P+7aSwc8Od6IjpaPA1m6Bht6s5bC/46vkAi92Ckf6aW1zjxXWrLD3OvuMcEXOX+Y+LUyPjfzTrOl
AwoJYhwbf5Z90+RFHecWcZIjGGFhH7aU1LzaoOI2n988tXwZMvudLKsWXkm0L8NJsWutAWvorrAW
06S29nN1GH0upUKaFJDUfzu68zTHQ43iqmCIfiQ/WbIfje+fICQ1sYm+YCZjkZ1zXWZqs1VmGeeT
Gs45ynFBkrh8rsYdUhfZbyw2EyI/y51DpZqe59yhyBItybXp4BsOT/7y/1yiON4zPeSilvCvKwFw
a9foLAVQzpzMiEdIPo//OdvXm22bFoviu+gwMpUiJelPdrrk/p0Dn7AUzijpR08WEUZccVFjyVsJ
Beu8291pAEGYhOu/DhMA0yDVuu5q339l+nAHk1smZdc1hLlWWTFHE53sdmVyCiOUg2TqvSlhBizP
RsUSJ7vTpHz00w35r8DYVnuGrWJ/ZIIoBNqHbYnXpNtwAhzuWyeUzOhHG1k609sWfQ+TLYyxgsvF
fHF6/IuS2Y+YNVGxZEsnGB8VjSBv3DqzP3Ji4ZyqbvAyem/aea5RsEA4++znALDFWK3wC268eIf1
Jc3dq2ssrHJvsxX5pHWzT+aDWVrsqJEpbC7xERfLHEn18SWyJ7wovO3cWRP3a8bAEeGOqwBBZDxE
M3J0+tYfk+Im5BSzXpp2bfYx2V4WOyakZIGRqZGoMe2OEEoyTufThpHQTV+0rjmx9cdaRQ9/1nYE
QTE1r/Z8zpllWzQFunB38QxndTZpDS1XlOooiQ3vLNujjg11mrYBm+na0fT/x3+udwOntkAcLr6h
plfF4RWaqWkS3P7GYA2A4S3P9Z6yOPUwt/aoARpQa1y6uU4WLwRKKJfxp2GRcHVNezAsztSK3Qb2
W5sWOto2Z5taiXXW8WyMsI9pVPBOuyuicsZE5tgkYq33zT+z0ZwIOMYywtchvNXBCI1p3m/mRuJK
o3UZne0oOysmWceTkP/HRGz8F5mMGUxJRojqk4sZmOTfesnQ7VPcUmoua29IeSY5ud22h+cce607
r/q35tXb0GKQRM6gN8t1yCn8ANY2HwAw56dZKgyaBmazNs8RGXIY3CgwMaJ9z0mI7rXnhXqB5nAE
ReC966mNnIDGSucVQIHn/uPOdDAIvIDv9Kq80qDwfuD/lh6UW2wLJnTfL3p/XPrMYFGt9219xjRH
ILpex+LwX30ZR1I4izRzygK0Mvf+VT5U9v97/+gPFRELVpuahqpbGeCoN/7HIH7lTLmWpsssAeFw
dHG392R/3v8U8BaNeqdHcKXprT/FqAVsT67bLhZDPrliLV3g/RlRIWZIdHsV1K8hhUclIBOKZmqU
d3q1Eab01y3ZoKQ1KMPrlvfKhsA8ITYdc3iQ+ybr+d2w1zrSZY36+gCog3GddZXgkrXwUwSvO4u0
JKpmCiWavHNk8tjOpnwd+CQZZxShCjih7DGePjJnCyD3TfASAwCXtNuGeoxXkeitI7HSMf8shDyZ
Pb1YJzqGjKQlQaVv+nXfx6r1qjEyog9smSdw52N+IP545kJ4Rvmz59HW9+WW5gOICzYvUbBXwZgq
jVsvvWVKXMj1A6BuW2ttaR5F8iJ3g9zoBekOenOKW59xllSVzYvsYIPKaa4HJQK5feAvvVOW8uhS
fwpSFl2RKd0XuZMPf01cxvH1iNKw81urGC8DsW/6O9YJ3yEPy/OJCWOR5Xe6g0GDgAC4YSYnaj9W
kXoqSHU7r2v59HQrYvj1PmL/bEceKvIS0ZM3HY2j1tIkDyC8hED9F79+mqcFou30XK+yBoHVsyiB
50BDzSH+frYknqERI79S5nFH2hBIFwkjunxtN6wUYS3fU9bgTBwQtbhJMaZv95hpUAGsZ3nzsLsH
y6I7GDVT7YlRVl+X+LROoiFpckUhUQV2D2gFA132WXRt/3gZNH+4viefLstGHE0+MYwj74IjfKkg
Z/AlAorY+1t7mweVTMkOrdfT6tI+j98zqIjcLp/rN3358LqR3YEBZBYklySaHkRcn/w9pYAbayUM
HTKU/tAAbjckl4EMNrxSuj/86mu2iDKuz8HzE3JLws+Ns0jgUf6Ow1XvetV6pUVOdO4tGTAkT01v
A55YaKa9n9Wlkiwjl2fqsVqhNR0bhE2yA5KEVXxGQr8tI57oUeKHrwYmV5B/QsrZIhim74ApxjIC
QefDYQ4qHCa9T3eAgHszIPoFu/4dZ44hxvpWdHkcFkG17J5hI0O6BTs6nKWONhi+qyBPCHXPbDoj
G2cBkQ/E6msgFlbeKlN/f3yxhaRcWaLK1IjT2nXLuawZsNE6rD/zf6mQmWqa5ZJ1jrw4G9DNC8U1
fjnvbEOghOis4O71kJAqxaDCmEEwnh4Sxxhe2czWAZKsqZqWFObV0E5DqOs49jqKeej51e1rVLhZ
yH6PiZsI+spjE7SHDTgM9CZ+lJqwHJS5ZEQ3jMhqTvatLuEcvqUJwz7cKO3FwcEB6/fk5hOK+kGj
2QxftdRZHqLZPCf0vgs2XnibKcqVtDPtvem9B5hK2huFyNhzx9pf6bNBoenOE8rg2QA9b7yIGdz9
xqmIsv4hABZUYIhGVHtMOa0jSvEDN14VstkaD56Q67QeO5FtUkMvdFRUNJM0gqe5aYrTsuNa+G9s
BebUmnWSmqAPkKe7Dr+tqRXH1HK6JUv05rQ1FQLmuzAZfrPPF2IVkWLFPIUdpHKanN6fdpiKNSqk
6E0tsLw5XAI9wTLVvg94vZL07UMYHgO5AJvpsDoSLVZYQGT0VeD40mTVbMuHwhb0jRFDWWWrrFhb
BI+n8DfuuRnTu1joNbWJiSA3klIbO8DONSaOitrPQ9W6mfFjWOgPNdEW0kpb0U1BfFYnzlw8rHpD
IcuGjy0/lM3yVAX5joUVC2bHtL4Xb2yCxhHDwg1XgmwxGc1w21Hu299mzOWMy2BTrRBzbw6tv8BJ
znlcxn3r78j4ZW+VeGFXEY0wOavpYsl247PF7zHSBcJwfirmNXKrrJaFHtuZ9O2rx57Dkag/onok
nsJypOb8xtvEDN1r2PAmjFgxlp8d242P2nsOhGpNPxlnS08KfhzPJXHZPSkYbNH3/BYuqQdZod8d
1e0Cu18aUdwHPCVawp4rWrV6lgo7Lm2zBFp7D7OUHIe2bc+tubItWMk4fJAi1c8ch38O+q+o4v8z
DYRyqmNqQZBRdf0CqEEk+CqCM3XIEgA5Z1ifOdcJqSr88ttvWTsm+8yLrpYQPV+6BcjhcUkDLJh+
7W5P5iXjyU1itlm7Pp+tMVgwJmtOIh+EfxAIXu9l9oDWG5NGvf2722SLjulStTgiOaquhCey2oei
UccuFKAZGD/GrF+TXKd26k7Fx/yZ567/ci+680EPx1KQNKu2HENpyZbL1vZOIryh/+oULemRzGuH
JwaJUQHqkqGZP9hmz+BILuQXg6h48E6pkvOo621m8Nc5eVcE1ObRlMaQxlSMu7VCOH1A8Opcz8Zj
+H/geRFoNfu6ohC9gnInuQ0Turx+s1Jd3W9poqockY0JI3QVcc/HVwTA+8GVceGp+QlUM2x8f08d
UDOwvjKvi3FSgAZRB6esaK+4Hl+O8ToMFo3mk9NQfYKO3zmOnUVXBCQYQ2rOywgNS+ODiE3dIsxk
/r+m/Ex+GdABTe2MO3hXXjktFhgzfE0sW+GDmFoWZaQrZr88ucf4KHqO2EGBpoQN+5qHF+DUqjay
XRktLzy954OU178bOeYXqUBlh1Me4Ni0olIxhcONsdChX+0XY7K9IgHbjnljywk9l0ox7KN0EkNM
BXWfI1hRjErEpC9OIJVCFSNxJJB9g25sEyIkptR8TF8qFydU9OeLyUquJuKdlSOcpJkatQ31Z7Qb
tQ9LrmfW7mPhkUXWEPWKpa6JHYn/HIrIdpC1f43cec0iQiJroVCqv4mZIyXX4is6WRpYyngxFNsw
LIen9ARPIPq/WgvPMDOx2WWvZTQl/HOs7f7Kk3JPhE69+STOyNBQ+Z5UutECM1Fo3fs/R95lq/Or
jTs3ue3trLXRTVu0XG4OwUpoC2d4c5H1wO25XV9AjIUn3t58PdTtvUdSolGpo8EZg1y3mHnnFIDD
HNZj5/0jVw5lOYC8RwD/NajXSOyRF1lgxvAxcB75cm2HEfdIHMtZIdyQQfsvLTmvSuwsiHKz6FlE
ROp+yyvTsbqsu1NmJFYAPTdsvIJkAY0Hnhv1NzJEtbgZ/+nseNt+XxJPHlIL6Cf3uGfao6LjdZkh
EcyPi0M56PyuDwaj1zk6DL3z4DSQuZ/yi61GFH9hXPTHZfwCxnps+Ag2LAaAoRziFuG8lTJD8d9D
tC+Nb1Rh8xX5E6c744KCDffFaKLjrc5iZkNjrgEtmbnCerYcq8K9DcqntyoWpoE/dTFJn9ZKKtHc
SlAJ3tnXbkwTQv4wpSMK/H2Gl+7jpdfwoNgFhckzv/Tm5D7UwaYgsalca3z4fqfhxuLCUy/OszzP
/uIM8dZEKR5ZEafTAIfhAng4HoJy8FscRioOdR8qwOlGEYVd5Wpy+8MV2hnQfaFDfYlZYKI39zPN
8h2H5Qpa6U5gpzrxl9CoD8tdAK0HxhMTSe4+1A/TkQqZ6EKQSvAMMNJUYuZn8g0T978YE59lWaq7
0PpfMCfXr4uAKSojKskadxOKyrGrkm2jZ2GtEq5FOYKsZd0YwSt/GmNsODMENCRoeFeZBrK05a/v
E9rINcD0s/S85b+DBdxN4ZuvjKF5ajBV5Z14WHpU1f4GztqJQhJLdj4Y011VJ1f7TC4BFljTAotn
MKv9Tbg5tUwka0nGP82KhAsgLN0QqBhpkT208RGUu5eiatP3y/2gzjNM2no3uLNN4786JFz6g8i4
QJvn7pFSTwAdJCCRltZl4NftUIuXUADyXAW2hXfYzpGBe3SNUUATiMeDSluWSr/9gC9sRW/xFRta
JTIWoY9QjugLmimwM2kTIXZ47tFbdEYPJQVOgYwwmjylODl0ICHD2pYBkNjVHzStZ3RoKRyOs44J
eGscRJPX9X0rAO/GtOhxWqY+l/aXzUA+f3jGAmL/TG8g8kC38vpvgLKXI6UgQcO+P/Di4FnbNHQr
pr/VIxUd/i6mx5eBwCowaQjgMl72NlooZrCrhK6bJ18efX32wW5YY2lcMzDCvGfoybvVdS8zonZj
SkN8yHUcAbxscUeqHnJVQo0qn93NwCyK3WnyTTQMy3po6pkvlznl4GbxCtzNl5RHFW4kFDUCuaqU
HUK5dkCUl08KWV15sZKpq9XlDjD6MGB3kfgppCa+b12AF3WBns9oWEtEsGfzwJS+WVEygddQHaiW
TkgBmKPy3SLJhcBTuFfPr0eIxWT4LU4u9U3FIE1qK0unkHC0pYPSFwqiL17MS75kzply+s9KyV03
YE+H6ii5xOzipwXbyXLkZs+U8bKRTNAKZQT78Yh/d8DhvEHYP8m/o/YUJsqa7D5p0S8cV97aZ7Sz
7/w7/8DN3AzZd+9mPklDN8vn98wq8SEgDpnOK3pkNmyLzxLaBvYb+3gRS6+eFucx4jiBvgiYod4U
UtbvaOILxEneZbdp8TRRS4YjIjPWoMUfCIGUezygLnM0Z4N21SVF3oaL2DBsohiYR7u11o6vDvj6
sVBWeysDf+yNQjx7jVSM28mhFAhNJyR+jvmcrwSgVRotM+BDoMwAHqGLgkLX5RQYD0Zmiag7vBef
pU2FbJ4SOPiXwWq8wWKMS8biTr03JnOYkdfqlmvgOIh2u8KVAB/61LbTjIsJfNKuXstIsbxZTnEu
X6q96AsEHR+rphc1VJJidEgRNJotK/oWj/7iAHOSJmuzt3QRPSMTqcD/N+DUvbPAo4TqVk1duCVQ
KIA2AN4gOoq+MaZ54SuJ0Xb0y80G1ukpOu/urp2WZiA2146oGXJTH4GjfSYRvMbEik1zsrWpAniT
MpZ1bSEsAlUags7CaPQZl6TDR/dvXWO9Ljsfky7LqBBwKWoY217uWO7OZMm93FXCz5N3Sg3cx0LY
y/1Uqo8W2AYaYPZEM85TXf+z11YVyC5CoQf88KcUY3I0sUzSwAVOkJBEd3nx0qf4m3VTJkebIM0z
QTPq7Ci05FLxvdWjIu+xzTrdQV80Lx903JjGMhI4gJ2nJDmYSmsx6GqnrMh32tM2Ej20MWWZMtS2
GQbWV+ltTa7Vld7GNtqIqFzDuBXwNub/FCLrecYlf61oADrhhLpb/q0tWVTGt/8wTQiQb2O5eZrd
Sa5HOC59C1muo/9YmzthaTUwhQWlW2NbjeCW1HFLipeoBpolb/gYlQLFkomgKrfOv1MPevLijBu/
jkmFl/hbSEDXt5GFS4egdAymz5xHfhRYUS7mo/YifZ9eGYmD/O2lQcsxThjROu9FR72CW6w1AIMo
ebXu//c+s1IgGd/je7D1OTBidQFoQ2HC5EUjZTG+fxo2ls7EfYRTyKMaa6ovmAGuqyk807+bF+Bi
1qhWRMwFxahsDtEU3eGgyXUCWc+0RCfSVYvHA1IXLzkapjjA7VSzff72b2FeQWdBHgEQwLQrXp4U
xj72RQGo6EEi2wpG1CtByMyRuzTKv4vJihP/QO4ac1Reb+fbRRa9n1KU9fGr6ixmvhaB7UE0mX2f
CK+K1m+ORb5+mQR3IMdj5My5jmnkHDx7T4wvrqi3x1iSRrCMep5vM0nSJHyZ0ykz1/87yL6+JCuB
GYU4XmvpmwlmjQL5t6Z2e+fP6yC49bIgCI5/CSl8mUqAZ9ou4yrAp6IGyGQluSX8Rj+2zRkGhH+L
QF7V+nZctuJ6f2BoSPH0TGGMwe8J6khL1i59gyRFYQBjMZPgooldLNrkW9Vu8hG+qOd9SH7cd3Di
3HuewzgYo9O+wiUmDwXEFJayd+TCzn2FC9HCLDjsNyJBeFeFTYPA+rIYjAg5KV4MbP7FKEbGc9XU
IMaCrxLGQr8Ep8M1qZLXRiGfLVymba2F1xyYvp6VlTRtFp+5gXoUaK1/gB9Q8jT8BJb8/4D7EsB+
WVtA7lBHKUxB9JeP2CBgo0LGfblKu8Es4U6Rjom36qb57YgMnyNKGlwXuB4zFBvhhhyzb66xNxlE
+xElQ26+DZ8FvxLqd6wxqnyG8FqO2fzachkXiD3la0TbxnSyYlmDyemuuwuJRFS+CzJ5rCFMN1cS
3Jxq/4lZVu2vZWCF/yENxvvJpxRK3v8hYPlF+aWWYc5Rp/2QS99cbe0Yhj5iefRzVnZr7xNilJP2
3SIaVVaUOs2yMHODmhjzCAbnLJuxh1XL792wjPQyDq4YoxMm3gVharZKKXC96TKBYnGPcMjEV+sC
1MvXtI6gy54S26be07nZTJz+Dpckr7Sshv1i4NS/jjT2fe+0yOwXum5eQOSRMaN4+pfXBdI6eTMR
JEtE5Z78WydpH41QDqMcZ6GyAXYFiSQS5UMN9/nOGOjyB5cBbsd4R/EwWxr19lNgapAduNOH4/0a
rgBUfKVzAfccJ49zZwaqEamJ8NLVKVjoDR7nGdl1+fVyi699mvqSouQBSSuqhUc7mm93GKqveBRE
fNe10B53xYLrf8Is9y02p1l9rsazvt4BrFZ1Vmkd1EvGgTD9Q23uPDeZZBghjB4kqkt60Rce79S2
vRDRMMzwDIfRhHzxu/KUUd1ena2zXDW+/c8Tr1Ba7iomRqBxjsH2vqGleRD2tZMsZ9IBcfajNB4w
x90qVhvEOFOMf9zJEeVFPX12oJyBZjn9T3NRWjS8uDAFL30J61Am/nuEGa+PwIvSg/dlX0C5Dxj8
6FJ+h4y1Ih9nVNe4YQ3uIb6WQcZurN0A2cwwmch7MXTmJLkn9KQHZy6wsaMeqUH+SYuzVO2IreRV
2kTaUxVmkPBLqIHKdWaj+Q3/0cWlAeJ8ztqsHfXgR84myy2YP4EoLIDC4H2ZsrwxecRn4zuohDbU
+6DbB2bXmlSl8lizVR8IPfBC574QmWT3yGsNEBT6c0gV1sEgySkG7wxdc/INvBUW3+qxBuXj7KVr
DV9IxU4j00OfbUEILSfmPT+LKKHY2/OoGQ4foKLwrlYZOb57nDG90B5SCraUj+3rkmAfLkmjnAcN
6mGC64/j/ut/ltddejQfrG8y17Cp86WIwndDLzEKOGzVPciXoOO+txuRqacxWdpcSgsj/+9nPAwd
6rbOkr4uwP2g6xf3Ua5+wuB7An5OLTVTAp7rRSsdGQvxZPP3EAllsZmNmB+GRIoLGQQnJf3jJgdy
WClCBipGhwawo19TCfRDdwgfmkX/W/Dg2Fvb4/yjuRsYbz7vShYPGQH7deXTtXy5j1Qnb14EYLVS
AbSxRwDvYskZLpEErgLfMlXjpLmDyRnPFyscw3A4P/wXe1G39RVKwMbBdnbhDw4qudYmT3sZoLZ3
/ijcZl8dY3Q73bK3syYZIj4K3w9c9adC4P+8q/FwPZ/UTTIhL1Q2TMvdWG+gJG1ldBfBTb+ANSgR
Ok3YcVwl8GA7V5R8a0qy7tA2vMWbGLpn84gBVx0DLF2/Z8yHmJYsG6sBmIrk2WdtDs0hWOCLpb+4
s/RO40ky9WJl14GbVuKIo+i4QCwYajIhJ9+4ERs24XB3VL8jYhf1SbGuI4DxgvvW0RK0db1TP2La
BnFq6QgAbfOBYbRvAfjxIlLycbALAlHAgEp+Hn6tYFZPMFxfaWS6VgSPu3pRvmjgtEd2TCJGwSaU
TVMtbmiZOlI7YVW5JD3sfeogEmwi3CMJvtg2S76BZ2MKtgOk0p21mDd9QY5hLmUSGXKaFHBLZx+C
m5xXgbpirF1G1cgCz5St6psu7O8VjMYJJ+ZqoRUqFLuncngdeFNigQwv+CtcJc+Ie41tDF7dJeks
2c6x3YwEH/sTF0+YDQ/Yr2fkzzt8UvVIFjKNIlH2n8Swr9qSsdX8MoqD1GVmVrf5SuOOq05irKzf
VG195tK8zVE1rNtDtfiF8lBTMWXTttdlSKNc81cPnFGT/ZLo6qYW9fw/scnShBzjVBkch2ab91xz
6yKpwTDADLeu5PEnrT1LMh/trtfHFBHIscUd0bj8JAfCa3jePUUVLk8s83r7AnJoYbkH5rxd5IxE
xMeWoe8o0kUhPDOGABkRCapJMc9tsVIoTiXcV5LnDcavruFYd42q3VGNPxLHTYkd2fblTwlPNmmg
hAL1OdAwYJmAxzUVU040Q1u+SqNV9W81Uz9Hqw0erFFFzHi+uowjd9HRhEoixdlb5UYcL7pI9rWG
DPT7MEc/OVjVqXFbKQliQ+lb2bxNswi2dQbvjHKmHaOAhpgKLvJC/wPcCr2u/OmTJ3ysjFQcZsMT
eF3ts1uNng3c3NepcrliskM5BJDPxRVdgOXmgLwApwkT8eimQ7SUrvGheiBIYIyHdlZc+NP0JniK
hxB4VlbM2jfNwF7/0IlLriUtF/Z7A3DO3yrGT3H+kz9Lv2s1zcYNZuGWPORoW3yrJ38EDsFZx5sM
hwP1TbzRAH1Lm7k1mBVt0qrB08ezcmBBCo+XMgsneEedB25CIHaClJt3lWekkfHoeJho/bh9fehb
f851Ld9oZ2c7OWx1LuR5ElRSqTaNydC4TiWp+/SIVDSexDI2Wr5xBNAuu/zP96o33ZgWbkYM9+AQ
wcnbAEyjH6KUihODtx68K/uUZcZCMj/eTFrF5mWw1+VgVztiE8j0P2I8vcC0gfhZS1YuaRfRdIp6
U4ihl2zuyLs2C1yd89v4GtzI2tRqj6sSr/nEWDdV+Rt4aFm5YKLqwF1Vdt7mGn76P3Gd6t7ha1I7
yAmUe4iSELe3nf5KPT7ONyGRhmiDk1inoKOT+ZXIvzks9rNUcBngOj/cR1jAzvFkA6FgM/bZ8p5v
yBqxBZLgJAxRVVi1qhboON4hQzk7lPzc4KeWVlYFVEcl6JxDBt+2YRjIQmQDZ8IleqMAkbO3XTRj
uCw2qU2oMP1zYn9kBcRaXJfUGSRHd4FqM+OOn1pK2G76ferpYjB4B5b6KSQ9cePvg8XTmW1F4geM
I2+USyPbam3cWEePhI0l2jRrJoTyA0WXxg4UqgczXqotuNXt+0vhhQ/UurCKgEv/rSeHgdLjwrwV
JDP1VVSwUcs0c/OSHDmamIllPWs7GZVbw3lX0dkmO5lJIsZh76j4te+WHVsbNRVMXIrFb/JAVWO4
XyqGfyDMFpIMnpjuAIzQCfRyN/FpW71B6mDIGC2FSaM250nvHFw2UE12RjI9jwUHAgoJfmL9k2NE
fd8ckgR4hfQ73WdvF3Z8kcs82ORN6A6Lbi8fPM6NaxDhRXYjZTdxoiD6vSxDHGOwS/UOkJK2rs8j
HhnitrigcqPTRBrp6w+qtG5mmoTHVhALtO3syyQPds9GH9+5O/Ebv3ZkoX6liq18udQIAWqNa2Fb
9sKKeuk3uggSen86hB6MXYEj8euSZuuzGguHXCt5A835SUwJ2M75NdUmpT8btq2UJ0kOn+vHq+gb
fUkTv+zkskGKYU1byUDbh8WWC2Fv+BUsg036f18byK4D1MzLPQsdCahmbKPWj/AZPxDPLuFODTOO
XrX0FMITDSVcTdehF/HEIbDx7oKydo3omKqDDUUTHsGdUb2zXWrAeNCITTeCntBeB1Sziz++S2qF
/kqs7p4XiTYot3B06Emmx5iYft9vEeZk8ahFqYr2pBSs0Uj6WeK4CRKpcxGen67nXstiS7OLYHPi
pPU4m56Vrkc0qQM2rvbFessycsof/Fqpg5G3KFcRXYPkniufse+g8AB5BgTPmI7QV1fhw6vLCrzP
YRzxmnRBjTUL6kadZJbKOjyhgjes1ORrrUhXqK2ZpV++TZgN9CmwC4rHBbYAvH+RSKHrfVK7SaT9
I1gaLnGCB353mTAbfgNJpWuoit4m4Fex+oCKn+N2a1lNRaSd09R+PsKzBdMhAfnKS/gh8iZWlpIE
PF++LZ6nPSHWarkHkNghiU3NTBFiaCRTlF8rPrWEGiAl7LSzSpYj+96PozXelnjrTD3wMlAstYbm
k/eMHc2brYWZTaDNZVaNAFbv/mkgeaKSh2UpBQUpQcSpsBD014HXRD2n4z3QMIHDg50pvcDcpvss
CFTs7e3Yr/rVAlOCQ6lQRRXOFPWmrvn325YBB5Wh3S06einCpU2wQrjAXK4DA9wiBEcyA85PUehB
phekBJdxugpzRkisnK46CyMv2mbnutDb5I2dl8HhMDzoexFSjy7p16SZvjL+HYFGq8UQ9icwQfYQ
yDRoAbRpZZCFZ7cKP03WJf+nRYxtlXu2/ulA9sMBm3mYXAPtSXuXkjzsxb/3AqFmvq0D2SHpJBsn
TrjIuUgHBer1dSFmqeLJHz8VvjCJON8JPdt4Ukg1VcaRuwDO9upOCy2B0nSk/9tTTwLixUWH49ch
FAWntrHkUVnz7RKQ2Lu5hXWt8Gf3lgWsig64C+RabXZXrRGDx47NZ0RlTRMZlMViqX0JzccoBSAD
glHFP/fhQDI1/sex2pLWLLfe5iRpb/qEkTD4Z0FPuoc0pGu8vzhXhhjP+bVuTF4YYfoeZedNKZpf
epWFXODcKtfZRdcp5ZSQfrv4rY4/swNXYoFwCNimg7HmkVzC1T01rPKKTvMQnP2Ttxx/wCrqicED
4VN+bfeuFGmd5R+MY+hnC1Qkm8zTzVgKxQL3zvz03ji4U+JVkXt8rO2cqbvBLVRCgg/uHpUCFspp
GUCsnGop5vnPivIDSswmD48W5l+uu8rahVUofkRzx2MaVoZkRhY518pAQon3s4XPwsqevLsj++3i
vdFrW6cfXtiMui6u4GYpqe+YwyoKl1f5IP81mCy8nlXOZZW1S/H3MSJ1iftHhH18QV6SZ7OAHl3J
/WZ3+7kHyIDJW5bTZSsKObt9niFHx8R+CQO78OexU7J0f/1OaO8pIYtlhPVRAq0blu+u0o6j5gJX
JTHIkaWJT0vPa0BUC3XlYtg1WjMuQ3DOMrGbAVD5KkMaTX7UizyZylk1sJgdK99h38GmoBSvS+9P
1V+d07hSA8NUC0XZxcqwC7RdS6uR9eaANyBh1q0ylRhG07AW1bBgHmzuNw1rs3W7/GsohUstuJUQ
s9M4fLlzRAfrL6pPV1rtn6KtM+zQPu2m3WU1l05WUv1ObJMmsdTTPhpDwhj1/zy1fZ7HvS9OuWCr
btrT0KEZuHZS2Rt/xelUjwMEokDx0DKuGVb7lgQ5Hzm/AWDv12+f7gC+IV4zrQfXXfK7oSJGTpW/
vtaSvO+IXZqJtMMHfL+ZDi1R0WDTIi/pBbeff2JbJiIGHVq1A2wjn93Fku2KeTSJ50ct/gBDaF9G
fPesIzVhdkovHiLuIgtR5cu1aORVz+9tjbmYeeQuruIEYoaHHDjBHkU2H4axn2C97OT3DwQga/zs
zH+pcWItgBtD5SHNxBvI1/pBgZcaMQMa5veCcqFycsoXjNzGRnbSHo/kYdu7wVPS3Tdkr5PeWjwl
q54R+xl356YyQPPXlzmQ/PQ3OJYDhhHnt9mKxoGhZ0Z9KRbS52k7hxvhnH2I6b91ZDkvhfVCxEt0
AWKDWwOiLAz3HuoYM21NKjGD/WLa3LM12Lf4pHJgnBCceJj55YjdVNwYR3vIbwR3Q4HYZbodqU78
zou+ya1dH0xPrf8Pv3mGT0gu1ZD/Ns3TuzobgdSDOnggQctlSzxxFJPHJECHMtUQ7ploDSGX5bDh
1zx0zWr0i+uNT8JmmGsZ+DgpbOaaFQx14iglzvXj1NO1zBafpNlZdLtzZUhO/cjcEO3xX98lyriI
JJx+fNmBS0g3OXqDXUqULx8DBbmg0Ivb9ajSrbiiMBuXwV3fRx+BhPQSpNTfx9fFrqH0T05zgzCQ
m3By0yRrb5hJCzz/b6NwYNyBUd+0410UgsfMJr/rd3qi6jUnLUK4BOR+fev0KOUO79Hjk8ImUlXG
d57OjCPdBS/Pw/MmerKbNcv8v0317udiuRJreqj+ecZviFjenUQa7H16s82AUMbTEKY6qwkMtfyc
nStkLvqgEjjaTJBNbFGhTW7RiBkpV+DCzqw3zldjVxJzAEpe5RlbbnIRdagXDHKkaWePfpdBFQva
wicZrw43zH2CpWnx5EB/RRYfyvzQ/kng1WD6jhlbjDeXblfJtLhD7ri+DpmTlUv0uj4peOTKT+Jk
eMwe6rwzUm/I8/KH86UOB9bjFUE/iYPaOAFG/z9lBA/VOgqB6CGfB4vo8Dwh5yFCvgu/TMJsqb0T
wC0ZDlEmU2+o7BsIABRvx1feBLGAnB1rdqXpqRnOiBnskLzujwdR9hGOyezwNK9OGBhmHOweZyqr
IaWkzsBtN5b7V8oX7paboJ9gydQCUwKYsjA5JmbHYX0WC9kMn5xcetLeIcYF0FSMbsWLHKna5oDI
82+ZoF8gvC3Y0Wyq4fT8fbFyboWJvAfvGUucaLBOqIPX4flKPS4+FNTFQE/Zns1uBpVg3uO2JrGZ
YxZ3d5oMxB3I5hcCGOOXzThvf/+IE6NKuHLwUDseYPjrsyQzisBdhkBp5eUJi/uROiUeq6c85PMi
gsjWdbsvRItj99pPd9ahBWYUzgsj1MfYv9u8guGwEa1wfKY3WsPcZj0DNcQ8L1J4NnyOpbagRNNf
HfXGL+ienxQRxJJ693X/3DPI43OZLa5NUL1N6SC9zt6VWJmG0Mh9RaQxUcQZ0LVHUefEIUudqpBl
QXVMc/DtBeFYh86yZNrVAvk5o8oF03OE5aAC60wqCIGrcY3fW2H2gBg3aGnC7qMEXv55glEUs3DS
HNQoQexvz4l5jKmmlAwNeXXi/uZhkHI3B06K0Z2+Izun7UvXhIXbvXMq5lld9Qd/TpZh1O2qbHTk
WSoNqer99f/GUqnT6m1YPFj8dXTd7vZdEpDDSL9nefSNSl90LRlmQJvZ4U4s86l3QG87oi2pRfZO
ZUsvlZEK1vzJbFAz/VFxfTecdjF0S/Mtq9IvGlOcE0vsW1zEiSCRDupLEyeIYOP2Ga6EI/kQHGWN
chGaaNXowDCeNq1liC0qZvLeB/h7tetP56fToEdHzJWTlKeC79f1r6IxlagkENW7YPBMs35HEORi
4nNYIP9wROJUrSdqcen1fl+wecuNizSqnN0uQPpggQCWZojHxbiLHF/gNxyUni4AqBOH+kIm1Eak
vlAoz7+6xMdCR78eDYnRs5tDeDh64W77Bjtk0344FRrFYo1ECJlJcAhz1FpvfsdOQADl94y4Dkxg
3OX+inmbZEMyG63Ew3ncTtQD4Df0SDZsc1YoNoCQb3BTd209Fg8mTt9aPJXlyfUkZm4hKLWWjugC
5/+Q3VrGufVAeLVJKZS5sYQb5k1Q3Dr5VyWmP4TlwEBXiEKDX9a8OkwWgZLPNavYnHj6vr6EMYYF
ZbMZFVTVUEtq36qkCplC3nuwJSHE9S1CgMLpIrF42CggszmQTQPqyF5lXkD5/0bRBF1TTBAp786r
dy+BD+arKLMBxlh4Y8QEkZxJm9hu0R3bVsqBsXysRNARUhzzDZ06QP2QsVryhecwfbVbLiwRFH37
ihwGvynTR6vtC96MyO3JQM3pxWFODZa9bABB1wHDyymZFdir6wTAuftjI7GLv4yR/Ipst7tl5wjq
Cru9iBW7eoeLwAROxcFy1hpECQ0NGLE1ALyjxNa1H9QFgbMIbNHsJHAXfdqT5aIL2Ubpdfg7tykw
QUNHBzVrZjpPCP5PCQtsAQxhWoNv/ZutDP0S63d8wPmxTbflwNFmH58Ct8jt2yFq83LBDYO28CX0
shYrypYoSWK5Uiue+4stliiR0cJ/OWX0gKbAMSHNc/57LsU2oYD3C1Ahe+nVIQeW4WAeYGpoSnUz
rp3X86FVT/0b1dymZSLkU4lhJYN5DHkAnKaHsjb6wrt0HM6B3pqalVzq0y+i2J0IRLXZz9krLcij
r95HqeKxSoQJ12/8pueP5HkJkwHer8oh5He3KDDI0BuHyjzzxY0BZTOH9//Pt0YTWrtTL5guFzjy
NbxPx/nB+D+ELQLXHPgrhbqPabhTpLAT6soTE9ggXLWAXo0xHnR/vnWcd5rdjhypwZ2wQmpgmR4H
4MhTMWqCshxpQpZrqvhYjRRyenLim9ss6x7U33CqELXh2zlSEeAz3JEStlduozVM2uCJgED1rl0M
HHMhl5ZIqjHgxMj7qXyqFgAwdIoPfOQKhW4ynAVF8c/sd3ymP6TVcuKk/lZL1ySKkbgHJj/U+Fzn
mweAAdA3MdalnnngWsIapVxJ0gGUTZaWe9ozA8hZ09oXRatAYEn8J/bpyWfRfHN6qgV3z5Ie6JJA
ecQsqy7pBDdIXV+HSvtoWTnahDwPAfZg97ugvxEoKK/ek6nmyVVGOCgns/cqGwAYG3xsZKQb7/iL
3XsJ+3Biu+LbKdVNKl2MQq6mqrRK5DKo0xTdhQnt1V3t26ff4BVwW0V2weflBYHOgB+tH83dM4N/
BDo2ccHCBo6cYReVJ74KVdT/hbpUDktQvLsShBMt5W1qMVO3OUFro+mTR9zFAMScMftt2WG9y1q1
XQ9RwVAd0YHZUTbeH6IAqjjvkZYwgGebQZjuQ+iuv40x2a1ZDj5DaLPh+kC5m9yzHQoc8OsHT3w1
0fDO39c76qgBbNnL1suTWpnyGZdy/WDkqkZf5KA96+oaQj0KFYAe9MtfQfjjljUrXsC7mdbdKSDP
oIZH34HFVJrPJiEjGFRNz+phZTmmzeAO+/gIiZhcS8Xu5IKOMjT9ayXqjfY+sVVPdnagPbkmivd+
g2hUPSSLu3NeUPgJiYGJfdVZFuI1YgJIfHd9MbjucYjRLPpuf4Cp6OoilNoa4F+v1fsmDm5102Gp
/yeHCbfMqqdUwab/A75w1KPyaLqoPHkbz8MRolEI7L6CadCulHCiu/y8+EmtBe5Lh0KTeUP7PWbP
q5qhHH8UPZ5Ih15/8bEdUFpoice3cKJ0frDSaB+4aXNok5/ZiyI+kSiBtRFj2YMiYg2OCCvcuKLN
k80TTn0H7k8REC8tAgxETeZP8dudC+Fc2hESCsVm/kk/k8bQS25GBXoEAn3Zc7qU7HhUk8lIcsuo
bCNixHWs/4SGZh7Zwu5VYIeTrQj7Ni9+C2NNDALqW7Q9XwX5ugkox3VSz8E3SjRMwu8h+K841ROS
5Kit9c0hadyvRfPryyz2zoJZTjdYuLuM50Q1Y6aHWm0FcTtRvqqYksGCZhjnFwKL8LSg3BAjdrIt
mJJBAhtwIHUG2HxPN+x9IY0xS7S8uDNLmUgGPhk5sAl9osD59Q4kxF52MFHn9Q64cac6AyNEeLmL
Lv4YVIYhHNLHujLwsHJ3aYH2of9THbxnnTud2yRamEx0IoQtSOXtvc+oyXOZXc5jK2EtC/T1qN4a
QGrycJIF3zxSsaraftaDK854KYf7x1PL5IF2HelJKxey+jcyHCYrR4YIQ6A5RQZpXOs6eFE1lR1P
OSYg0clju1+ykOsV86/ySjNcdJrGlPHGgSpWZ1+yLtAq7taTD/cGfLhukv6Ugo8IjwxkuBZNSTYX
MQPxeH1oVnVBFFFE7nnFZ3UUrGSTT/Ab5cKAY1WcO4qqxSUOVUDstElOcqX3VWL1ZHZl/+MCOL4q
B5uL49/Bm32+6HW5Le9Y3D9lhYu/wDR0oZWSjOVv0xZdRdIjzVo/j8v/s+o+09e0LgcpODKgkfV4
PppFpfmUDZBc7lFo53mAXX2EEiPubP3MYvt/7d51Lfj6m4KdFFRmqGczaUsDfrT0S6C0DEJJLprs
NNx4nXFY/Hr+x5vXRogUpu6U/i8XNm35+TQNiG3u6Ew4/of/w5D8gUeY5RFmPRP9ldQW06nR374Z
Qy1O9GBrH85M+XJ7+iF4ZSUl6kjfBUVlECLMbCUWlglEkb0z2CCmmTe7dHwXFicCUu4P8ym7lKzn
jsdnfjzJL+WJ2UERbj54FOvAt/oWu1qeVIUVyq+lVi1BfAQmrp1+K0K6hM800DkMnnDP/A18FWot
gtXeLJjlln2iSP83a11tMFz3wkbSgIByv8rjkEiDX5+8mp8G7erRf7Zw5ux14QC9xBV0Jr0clzKj
yigNUAQ0AnngBKqPh7Tshnj0Lm9Jrlh6zKyJh7TXOUYu/VafRed/xf3BfQ7Fh2Q14lMUo7rT8bYk
OgmAt6AHbTFblHe/JG65nJ6U2VB2lPf0vFDDaLxQHCFeKuAontyNQkR8J+8tBQfktqSsfNob3ujY
xoDthNinM71gpj1Dj3Nv6oT4+6A2LNETzggslP+TOK6UP8Xuwn+tNMMEl/fJEeNpccdHVFT95p/B
grhcliwWC4FPzghM8mh261EosTJuyD35/a2QsoeqWum9eA4bDfmxFMYJt6Dd30tqoakBl7gcdAl3
O65oygAX68qICaAbp4ezX3BFqIve6kf07lkg/Jg5/8EhwMRRPP3ezZ004oKGN++yi7SK1Q8ftQWP
c5yKvVIcccHZQn/akRrG4W4Eb5SS0uirsDQnVZELTGSHaLjgJl+wPAiyR4wiDc+DRMA2jcDPxUoN
y/7YqIG6jEBFYbQIrjAdG9sE4Dj0RFngOK1BpvHyXp5XNmbQzu90ZLeaiijv8RPY+yoqd5Glr763
dw21yCgjkqyuF4Zk2wcNRk23QW5EF3PSrJHb2nbr4lnuuQUm73GgL4OzyPiZy9lgHZrkCCI5JDEW
9dD3kB2PesrIfod2y+lrvjB+pAdUZFxnaixz9PC5SLrn6B5K3VGoVybx9b+iuCcfINxvab0S6/0W
ZDFZ7gZI2i52gWE+oh/4RWPcbCLPZ6FhYq8vuoGVffyUFjGxCvXoZWmdLJ95DiO6IcSC4MvyNXVx
ASzVG5JSXVmbaqQtbEdMpKm7sAGWHil2W8pX6MdFDs8U+9UWdu92wcgpo0UN2ho1ozxPp+NKzFtC
cTziyf+NhN7saCwQ62sA1sFbsjAm8cKgclKpj8RFsdVPReJPtgCxGnhrKNWzc3xOvIxPfbZYni5K
88mFEmbCxbdWOLDU+4pidmVWjep/feY9kyjjzC7Nl4IUWk7VLLrn44TRHrX1e7NWMFG1c7R+Q9Cx
Mzw4rh2l4Cm6RH7KpAAGDUoMVIfeD32hZcpI5lU1I/gxQ3Dh4T6ye9Jh4xdKP5+nFqFxMacTSrvR
YuFZCAAtUMH5wtN2ebY3a3Wdimm0CCm8E9KhP/76H2S2/UMPPqL+mEIKq+ap2S0t4pvHwNgp+Q+q
5bbNCl2e6PN2x7BdAwL69rFdqsMbnojamZjMuKpsI7qmo5OtPliKcaPRfcJp2sfUQl0GsQMEZ6nF
QrqXtVvGEAWdgGV7cNY1hvUtDyfqWIQUtdjqUGcTD5BfISRW/ssoS8CAYME2bzU4B2lYM11NRNu1
QkUYpMiijgR0rlD3jLHqkbWbfVjrFf11HAVbYB/8rsd6sQanG+RP9H8IpaRrGdyd4mzJ37qoaA5s
Oef3XwvRMcPTo6G4nyn8lVE71xGLTJRbIZh0gq+neGHT5zSiDNfoyWbiU2+gNDMQzg34Kdbfs98j
vVErpup5YZebUhlMEHFzk5K5Uk9T5H4pKa32U+Z3hj4B4HGGJg43HuHEcujzQg8J/KYcoQM0uoPh
O3rkJAL7ZG3l/Epy+2TeK0fmR55bofmryOyfjUYwEp4q+2j4Fe2jRedc58qh4u+PF4+nvCmhw1Lc
t3FRYEPgxp6A5OT/n4iLe9jApNBpY/cRslZnw6HNmKmN5LvGyriz9hHEAKDQPsQ8AYKkXPbPzi4H
dogr28FckgHOAdHDdHd5gACETvUBVIgGXj6whqswttyGXeHsMFVmB2gFy148DrIf2yeM9pXatsjH
Msu78EQDzKHTbAlhNGQgPwt8FwhRi7kVLd6N0AENW/mEXsm2KW1VM002SOZ5H5c9BZ12cZENYrAf
5McNKdtr/JoPKbv1JWjDJJNnOWoSqe6sof+sJaZQNMcvpVKDTuO9qhIxcPhsk+kCmv2jiVk6wlbM
883pNLw8yGNCS1fjNEfPXWmY0GaAiBiDHNXYHry0ej+Bk30BjPY7bHeFD/rXqjXbYpD6GtmNo81x
pRALAeo77bEFpmzZhL+NxIMiWvIVNnJTl5JfiYYBZg3T3oszUoZkugoEcv6yBFK35FXeIvFc2eDB
0giOcywcw+w2KZ33tDdFXLY7Z3axEcuMr3za4mdImHrVt5S5GRAraCZyLsKIuJur8LhtnhNsCbhG
VR9C0NLole2PcG/ICu2xMnVVrxZlt24jYuLFoGxRpTtFcJ27BWIKIgga05hsRkiEX4LkZYOE9586
in98o1LzGex5+k5LNkWwJDa66obaPqkkVpZA5nJyR2e0ZUkxjiH2oqBeXeR15xkXHFjoGtX/KFoL
klFRLtVq2zjc5UYO00pDdZatvyMmbTX2wXQN+G/54Bc485XsVuUKsEw65oJL6gmDpCpfzR4C2uiC
e3l7IPzZ1Llkb8Fzx6pl5XlkXQ0UrHU2cPz972KhEoR2pH802xq53+HA8pe0EwM6iAYtRmZrhfyT
24M1TiX0vkCb/caeYmpK8Brzv+dSZrp0kjqhcUvVL5WCQ63ypN6+3e/NN6/cnXuFr/vFr8CnTv4y
paMy1+8emRdLnCj+3T1OyUB7RQaAlkuyleDNGxICNNfFGpv6ytsujSbojqW6asU8PDSG8JrCa7gc
Y8Mtq9Ya+i4eaqJ9NYMcqeIRLQvXrOWSVNAFHxZhzSXUaDqaefrJQKZiCSWrlN8m84NRR9NR0v6b
HVI9UMPnAhmVu2Iw90ejU7Dh5euEYnjdBxxCivZEbBF0wpcynhvylf79pgpNa7czNOHQQFEYdLYj
yVzAk/Kbj0nnsKKOrTyhxAgr5e4agcaFdG03vWb0w1zmpFpaiowpJQ27mbpUiZU2dqw4BgwT8sYJ
SO4EAvQWswzKmqswK/RZkUN47pt2oBzNFQRKyxSmk7+g2ghPXub6xicaFmYlOxTBqkJeqdWWdYhC
VzO5gdR8milU5NMR/P+azBjz6MCuOnPpTTZlAZmNZvBhmzakdmvQKndsXsluVgN6pA7i9U/lqIA3
ti/bJ5UJcrTflULmG7xOYVBCgXo9maGNaF2VpybpRtKndNebWd9yL4zxTQ+OFxt17Yl64HT+z6Xi
inAPs0qKMw+Mt6Zqtuz3nBj5mb4wgbILvjITUcW0JjbVUyutPc8zVAvd9Wgd8o/9FgJYas+ixxH1
uBABaPskhBsvZnPh4mzkVURJcv/zD4IdJo8GwqWTNEpyhTdPyu5Xqb55SBKc0pTaAPDMpDcAcLRb
DhWkByHJZ3czKuhKM30TDaDS2M+tnTDd3CSjz7r+7B13gEYntInlDzO0cbq/H+11raJdNJslmo8K
MWLeocNYJo7pRNInVmsKsx7jnz3wewMw9IS4ppW7spMqBOHMMB0jgJV4Djn1L8Af1CfMIzk7bBn4
ecEFknusxwqFmTd+5Nvhz0MtDL6QJn1XmYdUENcUy2M6H0JA7oQx8NR1jDz0iaxu84kifB9NqSxZ
DZVhS0dYtUcEr6pHrlZmi0p0Qh4/ZMMfuuDiddcZDrw6xZNENaMq9heX2Imn3HXPbqcbvatceMuJ
yhBnV3B1QqGGeF7aoAT84JuPGqDOUc65lGc7yM93331qvW900Lyk5QPpw5++oMOtdSavGCM1DwNt
F6dqKCXqbgyIhYR5aILfliA47I+BS4Pc5NabV2AXV3ZUfUwd72yaB0nCA44fcWaZwvgKnz1m/W4m
bw4avk3mGK9Ju6XwjsxSKwlxNkvs1sjmtgh5QLeJOeBwxii8fiCHrZoUK3HHYERwLFmRg5WXoeIs
KOxjXp64ljnkx1cOfJL0moYQpMruH4cvoyNoajP2OqKgEYlKq5G3B2xzXVW+TsnJmkMWTBWBAT0+
cy+jtiHy/oD6Mg6fWFDdAk8cwVf9awwp/XP3GVTuIq0avqHGfJOmiWMPfI1X3qHKnSUJYTUrtqiZ
ThBoIBX6s73cr/qmh5VqFdfuxXSSgk5Ujcpt04UkR2XUSad9WS5qO+L0bpIqY9F8/gX9MMMsGFOm
Zk+Kp1qT3w7NmgE3s1gGOk0Kesgm5r5LOApArhedmdTqWDYY77SfoKeG+Gq6xe2pl2E+YdsgMvRb
nmqPoNS+J0p3CyWmcMrH6D5EUn0RXjMyOJLvbjglSnt775nmq2tswIfCDt/eswgwoP6AbEb4XEPW
dGPusLyl6kGp9/xRoFECMDLsxCwOoWeLXEtJY9Lr9/+a3HR3enG6EOE3eXJS7SbWAwzCT/hLOt5/
wgQs/X8bRJDZGaDYHpSHFx3Vq9EZYMZApQMtJRccu7FzdjVIA4E9f70mvVIsRj3jTqQIDUVTx3qK
5d5gqug/8w5mMB7u+lHhwGQ033jNwCgtFUD9kkRvX/OoMMyGgYQ67Q8xwtVHMD8x5Zld4myuirko
HfYHihzS9X3JDEsiD8Twox75G17JnI/C1HT0CCz1lsm+OneyQMpSDJw95jldM2ExLmjUWx6BjZk9
fiv4KHBS/Gw5VWJv4n+uJ/owyVLOqa8U8Sgkj58HBy2l6JohHmycBwOa0VSJc+yh+ew39dMGqvjb
6hXY38LojC9fXCr1Uyuc/wRmJoYMgUr4TmznKESHSK7Zx91xOF/dLyNNlXsaQlJz1hVRHYsnBRQS
BRA+lf5rWWwAQORzHv5VAk5c7zDFw0hw3ok+Rl7txHXi0LmKSdXj09ERE64CX6djuGoWqSkiCv5q
n+jUb0xyHV7CPQObJcWO/hpHui83KTZIXoRjLmJc0/7nqm22vJuSSWYD1llgmhnxKQOzFXT/VoSI
fTe/cFFtEm8RETOUpiq35sAyieMNjGyIiVj6VIvNoQgvw6QFZTiye+N6C52SXOZ30bAHAeYszeUj
1/BsIDinK5R6cpYT53Z6GUQRwhaYZYfuLmqKFk7cuWCW0ZgQ/vRcHK5WJ8Q8Ze7X5oleHCfQLuRv
vhXNs8irVr+2wV5njJ3pPM3GEMXPtW3U6gvv2L0KWiIqQ5s//h/KKN3l3BqWJ9iNnnjgKJuNQ2wZ
UgcauydSwNzDSGtFoUGxhxe9X1JeHTJ9VeRGGs8TYJjAl5acyYBlrJZRLW5vgNEqBqH6IFE2m1CL
IqfwGkKt4FAegq4sZejZvGTIXCSwEcs9bSMkf3f7XKT9JUuOS2WjmknQVyG4lesARLSMRqVsmAgW
NHqDtqRr4/fxO80Bx0EXijQDrtq1q+VCTS7ucuq37/AN4CfdT4c5RP1cd4mtytWsqFCsF8GEgXwN
l6GXIX1hQ481k9jpHpnLDkeAJleAJgqwTR3+HJpaf0QSHpDualmHxlM3wj/VjlkiNCPLeIUB049K
7V4wM4yb0g3vNh9DWTe7H+OPvtpDf0QleLrfWqhm6VZLwmngESC9BbHdlnLNQzw1F9sPAk+sCLUL
n3XmpmrDWyEMlv8aB8qYvXxTdTCicI4NORYtM/bvSIyvhsoJIffOemkp7qvAMb6ycg6S4x1n3mvh
IMzB+zKwGfT55WcgvNfE/8WdfFRWaLf60YnsetzUwuXE8rt1NxhsFxx/Gq/juXsddlDdX3TmZyx1
3av5Tb5W1XRTTStC+Kb/UJiwdv+BHVyWv8bCgdiUreBf29cXxhO1qZy9MtSOBHAe1KMSaewejLAc
gY+doZeNxUul0q4kmxa8Jee60KlUaGaStdfEWowtSW/Vpx82G+BXWu5vib5NO/6wMyOUCVtSU6ye
9i/Jkm/eBan36ch5zm+OqaN7Bm9yd89hej0Q/jQi4gnuzW4HtRo3k4NWDXx5odTKWVt+ppgdlHq+
I6Zr4poY7CX3PSbeOAMHFBOWuhYvwzXS1WROeYhksSoUnsu/r31uyboeFaWgMMY+Sbvlis8jk34H
wKZcnk+h3uGtXP83Qt/Qi8f8fAmXy0RpVsCUaiGeDFGRRFh71lTUxmEtMNIIfgjeRPp4LNsBKhHX
Q9ku426YXzY9TYb+YQouUJIFYmtgXt1+B7SbMnhugz0vvQotSn3amxv9iuaEewyP6OsPKYlrZ4vM
fNrFH7SWi77m9fHYuPIVEysS6oMmSAUb03IiddD+mAlMTesrsp/vTLwUZwE40WXex/mdRXIC0kHV
ipIbtsK6jtpqrMVmIu/uWZPqEn8OY/CL/hBogZ6Z/0KDRNFYMkAn85sUP1abPGGRettLj9HFcuqV
Zje8NCyjwGX8dhuKoTHWWO0zRXLn0fixuhIEdsGHJOhAzGpV27pCfQn4rSiGWIc+aJewvPBIh6BU
yn0Qm880eOpJzktpbDQBLIOrJh4A2ETe1hQH1xKiHFQ9ZayjcCEa7WFhqXGvs2eIYH/vwqjxeKgK
+bxGTVCnfprnPvKeCYzijQGKrZB+A6jUeDeJbGP6IEY6W7zSpdAf92SEoU/bagwG/LLm3O4jqZZx
TV1hjqSBKVEmjTNU11RuGXZdU0p6w8W4UIkUEqJDNY6mio6p2076PmkqYCYR6R8oAdo3/lC7XqV5
f4OiG92No2h2k3xYLn0AWmYXnsl89MkxNSIOelASgt+AHfle0Y/KxvEOMVq5C5UY1iiZ+Z6IhBA7
GfswyXNX71Ie/i+8KDIQN/X7Bx7YCZ1TIpw0NuL0V5Iw/BebDTjDM7xeLG5zl++y5a0CGvFQA2hs
M8WrcrYHdnxMl6Il+3nEVB9O2peD6YlbTsiqXPC8D5J2XOJzEanIJz0+574dvo4RP4ybB4hJpu+k
DwjE5qmwG5UkqD7wjCDD7/g3Jv5erjd9YAeMVuqe1hgfkbLsc/YAQ160EX2dxVZj1776eu2KEXxk
KVnvYpNaYIOvcoXphf0tkOCPjvz61HrMSzL4FSui/zlFpnhXltcM26UVHFDgzQL66mKvFJPaYCYl
RKtjb7xwU2ptPiUC9/5Ce3FQhdwyxVdKFUjwAQdsjoHOzXOFfgScUsfoxbxqaRmqiLsCMiDhKBbB
olviZxql1MoEGnvq8d8Zz7EaQJAxopHh5wPKiHEDvuZYsyrIGY+Mzvd1ZEq9Cmz7lGYhJohXxWpi
a3zYNMa6VpfGRLVqwVE4W2u3isf98vW32RZeWD1g5TvEGKiz8qh67hUxSC61NFa/KWOwnR3adtP3
KOczMNWEUnPaQ3fo3XrsuoD2y6++L0Kli/U5ZV3JHO0IJC5v7gpavz3xa/ITvQAGNTtQU40OAdRd
nzvkrvN2EP+L5YHx5jVuqfXAxWPciNZeYCVoNkQEmtkLYeltSLTwz2CXAZEUXxV2jIUGtP9waEty
acFWArJsImhsCDgI86cOA5kn1De5oDdkRNZLM+DxLoGruJk/Z/sedz+0YqkiflZJ6Y9QXFwsKcfT
sqjDfph3ISSNp2HG3GT7IjQzQ29V7X5zEWgxhh0kxd0x4YXyOpmsd4trXd5rXwFxemNqF9ihkPkr
spdFYZLNDDHUx+wDcPlgwItZj/z5ZcyfVGjnTCVpixnabXfqIF+C1U1xS94l0/6qLwkOwKol7jfc
BIHdQEzY/hE9Dmj6bA4XSJU2au1wwfma8LZzOB8ofHXF4c0D1NZBHxxqFGkHGLvVLKoLc2qctyCS
VkGadZ+pd8pMm8vjDYBOnjkrrQtoUpysmaCDID+G2s6aecW1HfFSLxXVmuj/q9m260/VuM0zJFNf
yvYqkynNwsxPhYZS6TxigGCNrgkLI2Y7joTvGJCnE9G+ZCG1wfUGUgbANMt5RPRmOt1Ai1stmTow
lfKrBUDlLvXMXFWL4eEwVARyMPRF73vqFunC2az0Naderh9fnOgvr83MfzCqz5U9qs16vWaB8lwg
AXq1n+/Ks7c/T63h+PFZ4AkkNCua3OjrJg6Udkn/cXsMLVmJSBdyB+UhWxB+vFe9M2D/nqJr/V4W
auj2PwMr6T0kRVqJp7mOVAHFgKXPp//mbj+6dZPmO9K9l5728mIEtvNtYScH5jKSvP/tE2N61MgG
EDaM7XEKEQva+Hcy8nMZtJMBGIqZVTUJPoGvF0sLl2K4ZKTTbA4ZjW1YQ+lAKRc93B1HxjoUGSV6
VVTsGy6VGbeVZB6WIcnT1Ny1XZzznKXB0mrMknKP5YQaO8PIHk+WuUG3/pdtM37yEkhrQw7KUbv+
QdFF9FxUw9FrUY/82UOQGymV85muHQ1Kb82fdUMxFwpTjXcBGCWkQA7PKmDj3j3AANDuELUGlaXi
yhuiEVEHq6m46LzvxUDReVvu7+ju5Am9sRjS7FS1p5bsrZo1Y7geQ4JabXTj+XOnlDJDqimqk9E3
I7gtL5t+bWO4mce7suRnJbzKCjl+2TBbXg2WxChlb5V+gBYBvOUhFi/jXe7jSQLUQ1Qdcej5KE+y
EJxmSRTCJ1+BZLA0VhUtQNp25muBFYuSzpWJ0OLm4R9CE1UlSX7Va9p+21i688ECnTjAPheVrvTD
Xqi5J3pdoFFIcEriXcQqEuUjM+aPWOl8mb90CKQ9o0asjTL2IHdVX9vdkyZEvDgIKc7z8s0F5Dfh
DfLpO8HgmCImPN+5za4sbYqRK2v6j5i+C7CqKJga/+DeJ09971OZvz8exOyaSvbQfivEkDBLytxY
Hq6UHcfnJ50NjPeeVnsEbUmUVH/0MXpRLhqVhQyTtKZYqnI3Bs46hSMXm3JcFORT0Ku8tkczv/tU
CAhCUUhlO70DiTyKVtt7oa9eldKlhRRuB2fWtGVx/R/q39Le+hFQeELA0hsMhtRwRtoKrn3tS55y
ccaC/ZpbyhMcXzMbAUXAlCsN1FDm2EPW0FWPVXd8i+6AUUa+ovqAZLArVB0N7cw6Iz0Z61RHGIRk
aKVf0C0+7vwAxjuMECATSGtR41C3Leu3DBuUfGiuc+mZmLjo1I3zesTdT71yoQ85v/5FeTXJsuf4
DyGN+57h5Pc7K5qh7HlLpqdR82rWRiXvAOUrUOEHUWkfGP5ICPQPGSuQDDH+kISeZXCxpeRoS0Ov
ck1BaghVUm/h6mS7Ik2KEH4J9EeT17v2zDKfjcM/tr4EkiEKJ0COE9aIXYHyrHwgxQ642GleRsjw
MnfD1hiJYSeMPOSn99eiXkmPMy5mpekdSk5h3i0oYX7YcMyJFroVE3c1u0wD+cGitgqWwnnzFGEN
J1UATE8yLh1ChZikC27OE+RTQvyPkq+zJWsJfCBsvbP17jw44qOe/oIYKoWtZKgD3Ak8CSIFI6E0
V1K38/2XP0HmtcD6/Qwr30A5kUEq+JPBhi29lgxHiUVqykLwKjN6K70iXcV+iAldzoLLqMmcqcm2
rPCSLnetWl1RKVnyRuePdEKXJIO5TZeZ8F6Lm9CfLSdE4NNHzyhZc+cHQofppLi55KUBoYvqV3y7
yQaf/FBmMmQIZgNMGTDHKFI1Vd8I8skiDszkYB8kry+nnnvdbbQQ8P0dJc5QNwhGbqTh9P60ejfi
4DO8ZpRMlIIPzLjNk7wZvZhWlSBc1Tm7jS/vu7/WA2fUYVu4AhraqcNHYkLix80dYZTpuw==
`pragma protect end_protected
