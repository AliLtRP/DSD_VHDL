// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
B1eJv/sQaVGqLbztgnC/zSZiOnxQqT8X5te4Egw9Ch9bXgJF5Y2Vr9US5PjHEZLrNTmiMBQ06POI
Wf5VsB9Lz8elpgm1/2qnYzbKniC4clEi2J9XGW3O8hXOOyiXj4VpzWrPviZtMJBw9DoUahmqyTdQ
EzEmbEAq+d3OdnuVI81gzbf+CMuYXq4bQWEe+QnxspyTsnVTCWNUyX9OKZX6IgePdpcOZW3tipvS
LdWznuxqshTk6V9PIsAOK3tzpsFJsu3paJBkz1ErALXv1xh9NxpmX4kAe0y7tNZ1chf5UgUz4hff
V3sLUmUubF+8alzst5+LDvoH4dVVApeGeLuUlQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
DaN5dKWK+Y2+hyDld6MSFg2N9ou+ACKI3yHaGWwLrOWdbxTjvaNiXV9TszHdWgwfAltj7DGv8nsu
D0owEhBQRv1m5+yphnAbWKWUOb4YRxqFMWyTq61fh0u/6dQV9XSMRc83241oodC+dxdc8Jksn4rC
jpdbo7pr8b2Rp9me7+ZYTCwFqrrw1562QaqaoU9zjf/YiTtYBf79xQu7/F8aY6xg9qMsKCEb5dui
KlJwD8CWtFRkGhHkY9mtzXA3Hi+l1gTDOJtc1xTq6yoW03+ytlOYxwQMW5NL89tMk68tbLxw0VD+
pFue/Ry3gUWyhqXIBTIn1xtKIj3tzNd3JDyKqcG8SSxeTQ7h48/JJU+uEC6ogBXv1/8MKZ9T7e7F
CFC/q41p9/Wo4/eJZfhDTX5ciinxX5s+B1oHXUINyKJcA0qA0L3OA29MERushlcxbunRsuhS8JLP
711v68h1DM4oms338NfX4DLmAeXV7Y+AJtaYrCbIMjbTh3hEbzz7EMHAVufXO9AJetA0by2jcdUU
Epwtc8xW6OF9s6w6E19DPTL28wDaSyGJA/QbEp2iTl6yo4fp4jcMbfCClFvuEtljCwuvXoiFodSE
se6X6BR0a5ifrz1E9CA6RmHYykYqq8SsLsU8tTwJYkwa/ddnrg+Wh/B2KATUmJVvZB9JIe5PpZJK
p0mByIno1YFsLtvgmC8EJ/nYWPaOvmjF0yniUDU6eBVfu/3Rfsb5nRdcvuTx6MGCwdhTfU8idEU0
8kRx16u0tePi9sBeFY+ozu7SkgikMI4VNuAznooMNKVBqQs56zUlU6hWsm2oLOHzJnECCSOTmR6J
yxXXtEYPVgVj8IcvX94MTjyFEmfG6QwDG2xguLkHC44ps9RkwbUQu+hHygwb+y0lcZUGU2wDsOBQ
rTUd99gXSz5FvocPzhYs2EMShpWeagF5YYKapynT8VdtwOGmboLfeV0lzz94gjdipXSCS7vLfaxK
jI7PPfDsr+B8210nBz/ZQdQY8QW/Br40aVHEm/pacRpcPKTIaY0kTK0MDfnWseLUFIvmHVj5MgGP
gPVdbpt7sd6JIWHbVOUBzuZhOjvyvVTELqdnihJQ2v8RK8++a8PyAMi88sZLURNrCIC2FC87If9g
D4fQJ7BkIt/qAMtYeBXp3eqzAb/O/Jp62nyHjcLzsQwZ9Pvsp9OXYhMdHozx9aw4LQ9IlMvTT6Gt
ZQzrVsJiSpsTp5sSofH9elxKCcFOWoua/0DPdYxk/C8O1vaFpoHZJoVNnSasfypDWMUYAL9L68R7
TBXfpa8fV7pggjcxSf0enMIwbo22rbp5yWd/J/qeVQJ05S0HFS4a1ZSsRyKBSt59lNYHn2wrtI9H
yFXwBsWvBsnsXG2tRq5GR4jNVy6BEsEGW5eKmuRfqSSD+Pxd0ZuSicLqvi8tyrWKEIwUvJUHD2RY
3VSKWAEF8wI2+tATA/O6qHUH1lNH8emdJs/w5cGaj2PBKVyzwc97dQJJMhf8eTVrfeCcGyc9ned4
MSGdklHeVxizPwmRCbRsMn172DrN02Y2MixE+Up9iara/jQLFapHCAZRABMuMFVt5J5f4E0xS16G
Py4j4D/EKe7nELJgeIm1G2v+Q4JHETxfUewRqE+iuW85bjTMSiR3M7HRXcs2DCGEysYAJf8JymMn
fK0cQbXzCgEewloNmGqryrfF9lhxRZzt0f4wEJziNtd/TB9twWoPocLK6DefLVhi/kf21FwaAeCN
TVwsbqVuMJ/ajifenntKNeEzMth1Wgqk+WpRqxd6qhW1WgtRnML7f4AASvS/ogObAwSuEEf2AFic
rDCPe4pU0rY9E0i4lQDhEMg6y3HE5QQ99dh1CQJqGVt2PjNVoOVd7ncQyL7FZ95mnoiFYch2oxcE
1m3HSsrc4rcstzLNsWXtEMwBmy2xCaQQZxyTG9e/R0IrK0PY+gumL7szA/5tBVgrpsLBonJgdIW5
O12rIbgkSrRgwo7+6Guzym5ANiJnzFPOWZivtjQkYGLMAQISVzm9HQzueeOvc1b9DesDXT85VH4p
bsLejTjzlMC7wGIugGC+srtrH67ONSQszzHoMMyMsT9Jtj9sbi1CnVbPjRf/GfzOlhy5L6/xNHX/
U6INDW2FrCCmeiOrDVHd2xYiGUgSFXgP6JCCQa9BuNMLWKRhg/2naMzk5NJnSnp/xWsbKwGB/hZO
5bvfOGOoOa4csfKgNjuipNanD1XZqnXDHmZCTFAS/9qy9nbYKkg7iw6MUBiPBMmQPV5Zi4lbYNES
zU8gLAemL1/v/yhHOMR/bqqSuxrI5sd6tYNppTsn5Ag15e0ExCWjpqUaAhcSHHJT9m3MQ0j3pALf
gpjAKiVyOuWcTN4IYJwJ5WV/Ax3oxcYSoUfMM1YIHxtwZPl4/8TMXVLsSowvgxANiv/ZAQPE3fAn
OChFeWpDNOrqMaX5H1pOlkjXV3kHgopH3xpI7dlpMNvOCsMjfVZZaWqWPHfxPqnEwczPu9owj2KG
De9QEz8G4H8bflZM3ouIz5JOzvFGZ7i3IISrtfpICvUH+eR9ilGXfJhm/IH+dSbX8PrR+s9xub00
GMsIw42a0GhHNrZHBv1oCpux5IAh/EzyqaMwa1Q7+9++xafK+DC4vl2D9ML+1Sr8R54lnc7kEdvi
W9KW5ucyMwujwU7dJuJPcUgNvWltQ2+YVrqrvlKAXP0o5LigBsaChBF7GdeaYBjpincDFgF55ck4
3avbARVWSV2KN+4cZSVOkgnKfANDZ5mQAOShZMtw21XrTUOaT5q5aeKoUGrSInjepJuTncGCV2g9
SXIr9rXJmtRiGiYgx1DrlVJYJymalDAaGYFePkTOqZiK1TbVixtE87pocaD3iM/y1Lv2R1ZWKd+v
t/acpreMvgJ7PwlgIuciyowz6U3lUgfJ97Y/dYzAhunPJ9Rd5rt3ao0bxKbo8oulSt+LV8t0FeEO
DN7TZXyv7TMcRN4IEmMrK5wQ45AQax6H31ZmBNJWhqvLe3R4WyJozfpgWjvt5Ed7ypHGQpUKCCmL
biUyARgj9sRqblJvgz3oniueSt4CpQNmu06lOZlxyHPhHya0XjD5Iymlndb/5MJ3VnMmBXoo3cni
WmGa5GOgkot2bxsEgk0SPWUibPx3o2bQD4GV9vqAog2NAmadv5UWRf4jJqTmEzvCioOfNVl0KPXZ
i60Hu1qypje6ANQQUzQYRLBG5M0HY0Il0EDihVNZWkiEv9DN2lPeO/p7CjGGhCzKhfJ4n8j0L9u8
XzqCDGzmOyg/9adTXwrd/MbVsoOrRq6WXdCpIMhG9UwZaNMhJ8Xz5gYgY1GYfIvrZXHKUB40yDVs
Aa/LPO4gR1IMaMVfn85J41dxiNhjkXBa/Pc4BF7Xbx3Hcclvc8OYldlgPyG7cy76V8G1+buqMWC2
SKA7Z8IlGUK51d1XhnCoMdS/FyDoouJFjKF24FAxeE92oJu4LU8k6onEuNr4ZRncosvlLHAlUXur
kuwa+DvbcZSDl6VpJVJjhNdF+2x+cjrn6zjZPgOyqio5criS1xvbyTztoHjDXUPlfebDJaEdUNEC
S7lGW41peKWLSuajsBT5vHVtwlo8BZNepWmhyt/zdiAcBO2uPiBgidsKFuBdV+6CgNwEDaunk/H3
vVOxnK6bS5yYz7mEilWd/APYiKt3p3cEC9KtH5r0DyNZuS/f50RTVR8QsEdqAFGYNsXXHC57JpoO
zIlAJnGYn5f4tldWrET9bKyWnJcPq7iRfV23QdexySHW93bnOxvgaHf0UBdJySDZbfg3KsgnQTSw
aE74FIiP7StdyupEcwTLlKzWQQaCi3cMPUSGfM53m2eulP1qvUIcBYQX/2HLpOPKw5sJcidng43g
/wuVLjiOUQqTdrb0J9E6zgo3jOvSiJKoe/6ZvKUMLY5alMAHCQNKGIsfbFj2jcfdQPMXz72EkhI7
LP3cP11iC5OKUwU8vjXqzun2Yp3r9oHj+0mdIDQ+M5w5UEWICm5/mUWBtS2YVcAeHSdnoxT+/JGS
jR12c4v/+em6ruOrMQULcp/u1b/i3dSzktonr5iI8BeXOnqFpir/xLjbtMIRtEAP7YIVBDT7v2vB
ZVnbVkTXQ2ASwONO8FwwVI1yfTGHzHnER47bCvX1+J+vhwR04zz/FaNeF+Bl42HxTe0Vy1xVWtcr
L3LVXjcUTu6+/Jp3y9fo0XRbaMxngdDTmAl4ksn7Ygm7Mvbi5Lhl3aRAZu+5u++xQbapd/+qDHOc
N9jGCV6eatDRscV3MuXHLrtj76sTbAWKFmAgP+nXhQDdd4ZQsr6hmyvpFlrIiJmceWALjLhP1Qzu
Icn+mDIY/GE7GLshnAUa/tjhVrOMjKIIXSYA2wvG0HsezdFFYbYn9ddFcMxrHHtTHZa+CXg9CIZz
3KKR606DnBqzVrq+PsHFcYkX5QEngnjAoJiPqLrva7AwGxhfulYjnySuzmTGw5g2lBGZ7Li2wQlo
mo93g6SCeTflGAYiHY18uL4lQz5yCYtztYgb5B+Dz7k4GAYDbUBnMbyhhQXVB8CBPojClspwrp+F
qx9H0nW4+hv337u7yPpSzvjojX0ggh097qNvhuQvx0UP+lAaz48CbbKWhD7YfwX9Qbs05LpomLrC
vv7xjiZ/EQg6s56PGPG1BdX5SP1K9gq4/sOcoEgouRtqKl25pabsSmELKRGfVvMRgr5nua+a4dNM
dnPUVU540LWJ9fVJ5gSOe5NJPNLuesTZ4A/BvsJqqiQEGY9Q7m1CqbPymNjcRlIqVrPzlPtzGkZt
JfVAqbBamDM3k8Sc6Wlhke30QWyQOykvQQkw9ZEorJqDrkKcdwaPI8dns7HOipffxvpuWxkyRE+v
mEBJ/ldJlIRUNrJ9AF1OUcMrm4ec0JevrAT4/3q7o4t+vts7xzvRNML0fOGXDzbr3st3Jk/R1jnm
0W8a6+6LsHMhZdBv/0cdr8RoSRSOdVuYmE9m4wERI1e7/LzEr/wqzGiKcNu1f44bUgJ+ceBYkfUg
oZXQGgMdLLFLQLuuH2fZ6pfzDc/NnTMMwypDsjjxs3C2Np9dJuv+4OMXArGxVzbY6FAKZqGC4W/F
Eqwc+dS0bOYdL/h0UUCDP/o3o4+vqHvoHOWbG3M28nXnmAmbtSkJI8+6/1pSu/0pq1PMSnvJqAyf
0uVxZB3pzFjd0505K96fpUmDGDnBEOoWgLYG3ujJ6ahE/ykJSCmOc+Nkq/YgSagUFnqWjtn09/nW
5uHN2Xj1u5vjkytT16L8wLdzpWmjXugEIGNI0COiVTRlotvMW0XW+Bc7QXHnpHjPXuMQaG/LW7p4
5DqPRtt0p/rCiDYk40wV78PqR/QfcZjTLzyRs7qk7wHsZMg1Cp3ofn7GSaEuEuF96t6sgJfmn9U7
vIPZOy16idVPjKLj+mCikJxWSdMON4506Fjq+eUxWFjWVlAkAJzz9B/dJ/ZF6kMs3fRD10PXxTQ+
ugAf8UfRvjOcplwW2gCIWBcEfVaIN9jJwxldZ7KpZx75b2VveV0tI8Jh4EVoX6mcJtC5JDvOuIl7
hrmSPfVy1DxQjh8Jg0qZlgLs4jjceBj72AIl7Fe5Xno9xTzq3ttSVFZe3B6sOL16sdKJO0J7onLT
EatGebbCk6+9kd4cujUybydS/ckOAC6vjRSnEEfqh5Nh8TarO/q47Om3I5yQ970eQUtiXbxNQTP5
9NQ0ksvhOjTTfDp6CVC2KhijI4PSFajX7Ll452DQdySRCOLCnNdkUU2Xe9NPWR75xHZM2HJAg9uN
8CFrJi3Fena1f15mnWbjVsH93J/2R/9G9HoKXpd7fGrX7R0qOOXqfDVzvmZ0ylpjFkNhpVnGmq2i
gmZZyag2AKTzz+BWpPdvnADEtq1taF3J2sqIxQp1iGjUT3Ba+/cLDZa1uLAsYGqkT1B6u4cnFXSY
1fJggkj39OdtVdrcFWs4lcBC6pOn13aZaHWQJz6XzVgXJPrc7x/hCaSZh6uICmW0nfvMT0TyywHs
RmDSeVdc+W/iWNOYos8LQk9rhXe4G3L0PBoYpalIDYnjayE6axvK6GT6XFV4fPNeHKyu0FG5I1+r
6M9B208uAfTKukdLzyMNCpByeQ5HnB1bhVsFilZMLFc54FcSEiME526hEaF6ujBd7NCgzXgOfLiR
LDzqvLwthIhUWeP8kjhMSaJpRjMHv2pZc2EjYNw2DyH4jNsC7pN4PEO1DyePScdOzWncb31Syn7w
rG9UUSOwYmphBaq6pPqLHR5uQvX9ZbBn/DThWHglHHkcYdQl2wUmGE3S31Vc1Z3rUS9Rb3z5Pd7S
eWfgbR8JtpJ07HHatwgBvZAcnWmwl7ui8TzIR7RvAYoqyDNeqMd+t0PBHD+RokemM17MzzhfEzpy
1SEcN4tz3SnZmBcIZVShZZnSsljoRY3KhIM0L3iEb5VH40skzYNmcF38oAIHGQt8sK7s1MKO4uwk
AuyejilBkzV5dqRIRkuaTfRgh902B2QxHN8NS4JGjRQYG6OAXZ0KSwKe3AoG6g4rKGrwRA2/qRQ+
q+kiNYLnzC59cr8PobcPwSUPVF1hToFWRLbCHvoHZDfk0gde2+f604ZBc9xg5WMsVVgPSotRnZsY
X3wPWlibXHB4VmlR3yO7TedMplQQRvZ6FNo6moaTd07ECUZLtGOlNpXyphBX7V3/nsm1aEUZrrPJ
WqxeHf6RqtJvxxEeJq8GNKGiWMRKJp/B2DXgwHTlMm14o4GuThhoe9hEEXBcMkIawrNAlMt3qaHB
D2uyVqA0EO7YsAM3tPNEhjQWCyaSZrJtepDX44PWtN2X4K/PkpNqt9CxvPq1JTFz/upTOUUpFjhH
8tfBL1M9xCkCCv9el00Be55lOlCfRRJKFUy8i+e6yUX884tnR91MDUkMnTNVij0MFguX/Z4UcRUl
ouLZqgOecEaBWnIbLwU4HErcnV3AEewuvFHvkW6ZpDLaAYWMGCswM+KMxndvLpzDbTuxs2GioeUZ
QmqFn7/QI2KtH0VURAbgARNi0Q9EMHKz61bLEv9jip5v1D9Y3F85WvG48EOGbTYqFurQEgXFYuB8
UUbeSS9vAVeAYVs+EyPlZhnKwd7OwhtJyJqvyE9QnySgfv8V899/L9F/dD7T/9vENns5ZVGZeyZw
/wqMqRFhhZtXgAalcXwmrXogcnw5SNEEtophgBR6HNkSew0FGjcjf4HYx3pvkPW7H28LLb4idlBc
IADvIlihEICyQrhebNKdxmHp+z2cGd+K/D4EePeXng6Gr0bKIGH0ZtSqa3G0HqJio719mvQ6Xg/C
NV4RIf+fVxRyRwuYDJSUH5oJD721amXR+UEIZi4gN+V5SIMZbRz5UxfarQKHsE7u5uJo1vM+TCwC
nfN4kXiotwQ/erm1QfQ1SFWgLh3Vm5q+/6Xdt30WT7ZeAn4eewdUqF6rTDCTdz7Vh19k8T9Ob1A0
ttaaHNMwxfmouphbbzwT7YUrQjQQZoL/MWmlrGwYt2rudlQVoY6tJEACEqqIjDyGgV8jhEz4Wntz
kHXC0ecJo0mKkBeqwDWlrLCHeXta9N2cmYBwj/qoOvtxigRuj2v3+ZC4OKRJf/ALJxZe9kPqo6tU
ZN/GI9ciBqus4HmdMDw4IxIc8Z2xVrujRDAK8ovgFJ+lJSTQdq247tbhf9JYqfGesKyNOCsGHQ6G
sFB+TaQ82PXRsgCnQkUeRSoOkHr0NvhNmupRCterGr0QJBrSnBZ//3/WUOnR2DQXTRLzr3krl5F3
yXJmtj/G3aGqKuJswN0AW3qbgU2rX/6jeb6cD68VhGQFvNqqANXiVSM6HlIHSVVC56eOw6ov56OE
pqkxFQXOaDg/Jih/m9TwIW1bg0nA99ohe8Hy1Ei6Zf46AkqTqJGHmJN2f75MF1iDNItZzwbqoMe1
lFKRdZ1HHFy8DqxoCGRywyYrN2Mwuwk2D81GHClBuZx0itg+t3og9ytFjkbPNsDIqZ8RqbldDx7X
g+unZB+uccDzyrPcUbp3abUdmXQYFw61yqyUzgYe9GIuVKMo7qxPGANwCTWPz0JtCTGN3kXlCKKb
ApH6cs/iRPXQO6C/AHS/46F51oaXNToX6DBHQccOQBVvXY0ed5zQSjeyC8jmwqH7NmSC6dIaRSp+
fU0u7H7+iW+N6hNEosXTy2v993F0G8Ml4zJRPqAX/YtHlNsHY35sLdpnBHj5trnuXniDxbNgnPmA
bx+UGVTj0pJUyQFoeqs0XHEOQhpsXMoARYWoE9wApOY1KCf2h4g3QN62crX4Y2GUW+IXLkFCnjVh
AkFjsSPeSbqkCu8HM2MPYh7f473PjadrwlTYA2NlNOdJatcypHATF6QqJXD7Jg6buEk4oJWREs8K
wbwCuw+Z+XsZkKNvxIcXi0Y6tFFDsJVrVZsyhHOv2QF+R017a+djm6Cm3HG81ZPgKPVqPTZnUwv/
lBiPt6WVYdh2pmdujNV4VXQX+59sZ5r6umWowI8G5P0pL0v7uTr+Ope4MT8/9ndI2FQGIxISiG4z
K+xlOUAcUZwdCnpsL9Ynf35nWYKeuM+kFromk4xzQ1Gq8WCEM/RXA+ePhwXxyXaBnWGV3Q9L4Snm
s6wTHiYknNpeg1l6W5r7Y9QCEw80imIS4vvhyGBpMuVFYWobNT3WrJBDec/DRXNTEBK214zTB0Fw
SmOblxgTLp+afN8kHf593nb20JfwJnsRYeTW9h+gDDHIbIqPllXg7yOq/zc/W4IeXIEFJMNL+of3
p/ai6rBP6bMnrcJfTB8VbkiHF+EE3XoKfQBT9idMTWlXitBbP5f6hBFnvlW2g9/bxzkKDc6WQSCc
ciqTVNGijIMnHnS2dYjMeR/F2qQtvRAx2v0T3SLVQd+Ntb80Vz4M1Tw9iKQc9PlLNdhOYkKHDzcR
93HMsGUBmVyiXEK9YQBmjONYvq6UZdcFWGqxIf9fLCANfPz7ojjZR24jvpKxSeiDN3Ba5BUFAMEX
NDhJPBq42MlGMyj5vtu3desxPWBb72VyFAe6DfJ5qIbImEXvuq1cQFj1wVj9k5ZZIvRaQb2kXM5N
hgvXgCJeYMt2x44K+GaUci1pwvufddYU7E0U2LAXHu3RnDsrng7WigpuO8CXVwZs9aFS1rt5w8M5
USbzoqXyIwf4otVwwrGVPqySm/sXaMovBRsyJmw2UvMfNUspHbGdCEksjWMqyS3rT9iWLNX6StYl
YMTQsR5+KXKRTNGDpBSH/YNinaiTwCiBgeIoH9YmO2Y+wez5q0BSeiWJ4dthtqDpeMCTCuLTd7X5
bPTdIsMvbNOaZWrG3kjdMRleDq71UT4iKaTb37IDGLLNvfXK3jhRWoJtwl6Aga23ZC628AzkQeed
uf4TXXCYsOgRdx8A+cYJUxT1zKa8eVaDC6tjP+R7EgoCk25vY0OyuScqh5JU0xWj51VatFlOOxgW
voNN8s4Ti0YKzk8nVCpa6vgJX4K7Z9IcXqJF9NYF9MzYe3U0
`pragma protect end_protected
