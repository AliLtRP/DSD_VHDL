// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// demo_control.v

// Generated using ACDS version 13.1 154 at 2013.09.06.11:05:38

`timescale 1 ps / 1 ps
module demo_control #(
		parameter           lanes = 2
 )
(
		output wire         lcd_RS,                                       //                       lcd.RS
		output wire         lcd_RW,                                       //                          .RW
		inout  wire [7:0]   lcd_data,                                     //                          .data
		output wire         lcd_E,                                        //                          .E
		output wire [(lanes*140)-1:0] source_reconfig_to_xcvr_reconfig_to_xcvr,     //   source_reconfig_to_xcvr.reconfig_to_xcvr
                input  wire [(lanes*92)-1:0]  source_reconfig_from_xcvr_reconfig_from_xcvr, // source_reconfig_from_xcvr.reconfig_from_xcvr
		output wire         source_reconfig_busy_reconfig_busy,           //      source_reconfig_busy.reconfig_busy
		output wire         sink_reconfig_busy_reconfig_busy,             //        sink_reconfig_busy.reconfig_busy
		output wire [(lanes*70)-1:0]  sink_reconfig_to_xcvr_reconfig_to_xcvr,       //     sink_reconfig_to_xcvr.reconfig_to_xcvr
		input  wire [(lanes*46)-1:0]  sink_reconfig_from_xcvr_reconfig_from_xcvr,   //   sink_reconfig_from_xcvr.reconfig_from_xcvr
		output wire [8:0]   source_mgmt_address,                          //               source_mgmt.address
		output wire         source_mgmt_read,                             //                          .read
		input  wire         source_mgmt_waitrequest,                      //                          .waitrequest
		input  wire [31:0]  source_mgmt_readdata,                         //                          .readdata
		output wire         source_mgmt_write,                            //                          .write
		output wire [31:0]  source_mgmt_writedata,                        //                          .writedata
		output wire [8:0]   sink_mgmt_address,                            //                 sink_mgmt.address
		output wire         sink_mgmt_read,                               //                          .read
		input  wire         sink_mgmt_waitrequest,                        //                          .waitrequest
		input  wire [31:0]  sink_mgmt_readdata,                           //                          .readdata
		output wire         sink_mgmt_write,                              //                          .write
		output wire [31:0]  sink_mgmt_writedata,                          //                          .writedata
		output wire [8:0]   demo_mgmt_address,                            //                 demo_mgmt.address
		output wire         demo_mgmt_read,                               //                          .read
		input  wire         demo_mgmt_waitrequest,                        //                          .waitrequest
		input  wire [31:0]  demo_mgmt_readdata,                           //                          .readdata
		output wire         demo_mgmt_write,                              //                          .write
		output wire [31:0]  demo_mgmt_writedata,                          //                          .writedata
		input  wire         reset_reset_n,                                //                     reset.reset_n
		input  wire         clk_clk,                                      //                       clk.clk
		output wire         sync_reset_reset                              //                sync_reset.reset
	);

	wire         mm_interconnect_0_sink_reconfig_reconfig_mgmt_waitrequest;    // sink_reconfig:reconfig_mgmt_waitrequest -> mm_interconnect_0:sink_reconfig_reconfig_mgmt_waitrequest
	wire  [31:0] mm_interconnect_0_sink_reconfig_reconfig_mgmt_writedata;      // mm_interconnect_0:sink_reconfig_reconfig_mgmt_writedata -> sink_reconfig:reconfig_mgmt_writedata
	wire   [6:0] mm_interconnect_0_sink_reconfig_reconfig_mgmt_address;        // mm_interconnect_0:sink_reconfig_reconfig_mgmt_address -> sink_reconfig:reconfig_mgmt_address
	wire         mm_interconnect_0_sink_reconfig_reconfig_mgmt_write;          // mm_interconnect_0:sink_reconfig_reconfig_mgmt_write -> sink_reconfig:reconfig_mgmt_write
	wire         mm_interconnect_0_sink_reconfig_reconfig_mgmt_read;           // mm_interconnect_0:sink_reconfig_reconfig_mgmt_read -> sink_reconfig:reconfig_mgmt_read
	wire  [31:0] mm_interconnect_0_sink_reconfig_reconfig_mgmt_readdata;       // sink_reconfig:reconfig_mgmt_readdata -> mm_interconnect_0:sink_reconfig_reconfig_mgmt_readdata
	wire   [7:0] mm_interconnect_0_lcd_control_slave_writedata;                // mm_interconnect_0:lcd_control_slave_writedata -> lcd:writedata
	wire   [1:0] mm_interconnect_0_lcd_control_slave_address;                  // mm_interconnect_0:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_0_lcd_control_slave_write;                    // mm_interconnect_0:lcd_control_slave_write -> lcd:write
	wire         mm_interconnect_0_lcd_control_slave_read;                     // mm_interconnect_0:lcd_control_slave_read -> lcd:read
	wire   [7:0] mm_interconnect_0_lcd_control_slave_readdata;                 // lcd:readdata -> mm_interconnect_0:lcd_control_slave_readdata
	wire         mm_interconnect_0_lcd_control_slave_begintransfer;            // mm_interconnect_0:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [18:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                       // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                         // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                      // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                           // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                        // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire         mm_interconnect_0_source_mgmt_slave_waitrequest;              // source_mgmt:avs_waitrequest -> mm_interconnect_0:source_mgmt_slave_waitrequest
	wire  [31:0] mm_interconnect_0_source_mgmt_slave_writedata;                // mm_interconnect_0:source_mgmt_slave_writedata -> source_mgmt:avs_writedata
	wire   [8:0] mm_interconnect_0_source_mgmt_slave_address;                  // mm_interconnect_0:source_mgmt_slave_address -> source_mgmt:avs_address
	wire         mm_interconnect_0_source_mgmt_slave_write;                    // mm_interconnect_0:source_mgmt_slave_write -> source_mgmt:avs_write
	wire         mm_interconnect_0_source_mgmt_slave_read;                     // mm_interconnect_0:source_mgmt_slave_read -> source_mgmt:avs_read
	wire  [31:0] mm_interconnect_0_source_mgmt_slave_readdata;                 // source_mgmt:avs_readdata -> mm_interconnect_0:source_mgmt_slave_readdata
	wire         mm_interconnect_0_source_reconfig_reconfig_mgmt_waitrequest;  // source_reconfig:reconfig_mgmt_waitrequest -> mm_interconnect_0:source_reconfig_reconfig_mgmt_waitrequest
	wire  [31:0] mm_interconnect_0_source_reconfig_reconfig_mgmt_writedata;    // mm_interconnect_0:source_reconfig_reconfig_mgmt_writedata -> source_reconfig:reconfig_mgmt_writedata
	wire   [6:0] mm_interconnect_0_source_reconfig_reconfig_mgmt_address;      // mm_interconnect_0:source_reconfig_reconfig_mgmt_address -> source_reconfig:reconfig_mgmt_address
	wire         mm_interconnect_0_source_reconfig_reconfig_mgmt_write;        // mm_interconnect_0:source_reconfig_reconfig_mgmt_write -> source_reconfig:reconfig_mgmt_write
	wire         mm_interconnect_0_source_reconfig_reconfig_mgmt_read;         // mm_interconnect_0:source_reconfig_reconfig_mgmt_read -> source_reconfig:reconfig_mgmt_read
	wire  [31:0] mm_interconnect_0_source_reconfig_reconfig_mgmt_readdata;     // source_reconfig:reconfig_mgmt_readdata -> mm_interconnect_0:source_reconfig_reconfig_mgmt_readdata
	wire         mm_interconnect_0_sink_mgmt_slave_waitrequest;                // sink_mgmt:avs_waitrequest -> mm_interconnect_0:sink_mgmt_slave_waitrequest
	wire  [31:0] mm_interconnect_0_sink_mgmt_slave_writedata;                  // mm_interconnect_0:sink_mgmt_slave_writedata -> sink_mgmt:avs_writedata
	wire   [8:0] mm_interconnect_0_sink_mgmt_slave_address;                    // mm_interconnect_0:sink_mgmt_slave_address -> sink_mgmt:avs_address
	wire         mm_interconnect_0_sink_mgmt_slave_write;                      // mm_interconnect_0:sink_mgmt_slave_write -> sink_mgmt:avs_write
	wire         mm_interconnect_0_sink_mgmt_slave_read;                       // mm_interconnect_0:sink_mgmt_slave_read -> sink_mgmt:avs_read
	wire  [31:0] mm_interconnect_0_sink_mgmt_slave_readdata;                   // sink_mgmt:avs_readdata -> mm_interconnect_0:sink_mgmt_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_code_data_memory_s1_writedata;              // mm_interconnect_0:code_data_memory_s1_writedata -> code_data_memory:writedata
	wire  [14:0] mm_interconnect_0_code_data_memory_s1_address;                // mm_interconnect_0:code_data_memory_s1_address -> code_data_memory:address
	wire         mm_interconnect_0_code_data_memory_s1_chipselect;             // mm_interconnect_0:code_data_memory_s1_chipselect -> code_data_memory:chipselect
	wire         mm_interconnect_0_code_data_memory_s1_clken;                  // mm_interconnect_0:code_data_memory_s1_clken -> code_data_memory:clken
	wire         mm_interconnect_0_code_data_memory_s1_write;                  // mm_interconnect_0:code_data_memory_s1_write -> code_data_memory:write
	wire  [31:0] mm_interconnect_0_code_data_memory_s1_readdata;               // code_data_memory:readdata -> mm_interconnect_0:code_data_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_code_data_memory_s1_byteenable;             // mm_interconnect_0:code_data_memory_s1_byteenable -> code_data_memory:byteenable
	wire         mm_interconnect_0_demo_mgmt_slave_waitrequest;                // demo_mgmt:avs_waitrequest -> mm_interconnect_0:demo_mgmt_slave_waitrequest
	wire  [31:0] mm_interconnect_0_demo_mgmt_slave_writedata;                  // mm_interconnect_0:demo_mgmt_slave_writedata -> demo_mgmt:avs_writedata
	wire   [8:0] mm_interconnect_0_demo_mgmt_slave_address;                    // mm_interconnect_0:demo_mgmt_slave_address -> demo_mgmt:avs_address
	wire         mm_interconnect_0_demo_mgmt_slave_write;                      // mm_interconnect_0:demo_mgmt_slave_write -> demo_mgmt:avs_write
	wire         mm_interconnect_0_demo_mgmt_slave_read;                       // mm_interconnect_0:demo_mgmt_slave_read -> demo_mgmt:avs_read
	wire  [31:0] mm_interconnect_0_demo_mgmt_slave_readdata;                   // demo_mgmt:avs_readdata -> mm_interconnect_0:demo_mgmt_slave_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [18:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [code_data_memory:reset_req, nios2_qsys_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in0

	demo_control_code_data_memory code_data_memory (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_code_data_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_code_data_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_code_data_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_code_data_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_code_data_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_code_data_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_code_data_memory_s1_byteenable), //       .byteenable
		.reset      (sync_reset_reset),                                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	demo_control_lcd lcd (
		.reset_n       (~sync_reset_reset),                                 //         reset.reset_n
		.clk           (clk_clk),                                           //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_control_slave_address),       //              .address
		.LCD_RS        (lcd_RS),                                            //      external.export
		.LCD_RW        (lcd_RW),                                            //              .export
		.LCD_data      (lcd_data),                                          //              .export
		.LCD_E         (lcd_E)                                              //              .export
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (lanes*2),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (1),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (1),
		.enable_pll                    (1)
	) source_reconfig (
		.reconfig_busy             (source_reconfig_busy_reconfig_busy),                          //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_clk),                                                     //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (sync_reset_reset),                                            //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (mm_interconnect_0_source_reconfig_reconfig_mgmt_address),     //      reconfig_mgmt.address
		.reconfig_mgmt_read        (mm_interconnect_0_source_reconfig_reconfig_mgmt_read),        //                   .read
		.reconfig_mgmt_readdata    (mm_interconnect_0_source_reconfig_reconfig_mgmt_readdata),    //                   .readdata
		.reconfig_mgmt_waitrequest (mm_interconnect_0_source_reconfig_reconfig_mgmt_waitrequest), //                   .waitrequest
		.reconfig_mgmt_write       (mm_interconnect_0_source_reconfig_reconfig_mgmt_write),       //                   .write
		.reconfig_mgmt_writedata   (mm_interconnect_0_source_reconfig_reconfig_mgmt_writedata),   //                   .writedata
		.reconfig_mif_address      (),                                                            //       reconfig_mif.address
		.reconfig_mif_read         (),                                                            //                   .read
		.reconfig_mif_readdata     (),                                                            //                   .readdata
		.reconfig_mif_waitrequest  (),                                                            //                   .waitrequest
		.reconfig_to_xcvr          (source_reconfig_to_xcvr_reconfig_to_xcvr),                    //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (source_reconfig_from_xcvr_reconfig_from_xcvr),                // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                            //        (terminated)
		.rx_cal_busy               (),                                                            //        (terminated)
		.cal_busy_in               (1'b0)                                                         //        (terminated)
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (lanes),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) sink_reconfig (
		.reconfig_busy             (sink_reconfig_busy_reconfig_busy),                          //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_clk),                                                   //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (sync_reset_reset),                                          //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (mm_interconnect_0_sink_reconfig_reconfig_mgmt_address),     //      reconfig_mgmt.address
		.reconfig_mgmt_read        (mm_interconnect_0_sink_reconfig_reconfig_mgmt_read),        //                   .read
		.reconfig_mgmt_readdata    (mm_interconnect_0_sink_reconfig_reconfig_mgmt_readdata),    //                   .readdata
		.reconfig_mgmt_waitrequest (mm_interconnect_0_sink_reconfig_reconfig_mgmt_waitrequest), //                   .waitrequest
		.reconfig_mgmt_write       (mm_interconnect_0_sink_reconfig_reconfig_mgmt_write),       //                   .write
		.reconfig_mgmt_writedata   (mm_interconnect_0_sink_reconfig_reconfig_mgmt_writedata),   //                   .writedata
		.reconfig_to_xcvr          (sink_reconfig_to_xcvr_reconfig_to_xcvr),                    //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (sink_reconfig_from_xcvr_reconfig_from_xcvr),                // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                          //        (terminated)
		.rx_cal_busy               (),                                                          //        (terminated)
		.cal_busy_in               (1'b0),                                                      //        (terminated)
		.reconfig_mif_address      (),                                                          //        (terminated)
		.reconfig_mif_read         (),                                                          //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                      //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                       //        (terminated)
	);

	demo_control_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~sync_reset_reset),                                            //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	demo_control_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~sync_reset_reset),                                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	master_export source_mgmt (
		.clk             (clk_clk),                                         //  clock.clk
		.reset           (sync_reset_reset),                                //  reset.reset
		.avm_address     (source_mgmt_address),                             // master.address
		.avm_read        (source_mgmt_read),                                //       .read
		.avm_waitrequest (source_mgmt_waitrequest),                         //       .waitrequest
		.avm_readdata    (source_mgmt_readdata),                            //       .readdata
		.avm_write       (source_mgmt_write),                               //       .write
		.avm_writedata   (source_mgmt_writedata),                           //       .writedata
		.avs_address     (mm_interconnect_0_source_mgmt_slave_address),     //  slave.address
		.avs_read        (mm_interconnect_0_source_mgmt_slave_read),        //       .read
		.avs_readdata    (mm_interconnect_0_source_mgmt_slave_readdata),    //       .readdata
		.avs_write       (mm_interconnect_0_source_mgmt_slave_write),       //       .write
		.avs_waitrequest (mm_interconnect_0_source_mgmt_slave_waitrequest), //       .waitrequest
		.avs_writedata   (mm_interconnect_0_source_mgmt_slave_writedata)    //       .writedata
	);

	master_export sink_mgmt (
		.clk             (clk_clk),                                       //  clock.clk
		.reset           (sync_reset_reset),                              //  reset.reset
		.avm_address     (sink_mgmt_address),                             // master.address
		.avm_read        (sink_mgmt_read),                                //       .read
		.avm_waitrequest (sink_mgmt_waitrequest),                         //       .waitrequest
		.avm_readdata    (sink_mgmt_readdata),                            //       .readdata
		.avm_write       (sink_mgmt_write),                               //       .write
		.avm_writedata   (sink_mgmt_writedata),                           //       .writedata
		.avs_address     (mm_interconnect_0_sink_mgmt_slave_address),     //  slave.address
		.avs_read        (mm_interconnect_0_sink_mgmt_slave_read),        //       .read
		.avs_readdata    (mm_interconnect_0_sink_mgmt_slave_readdata),    //       .readdata
		.avs_write       (mm_interconnect_0_sink_mgmt_slave_write),       //       .write
		.avs_waitrequest (mm_interconnect_0_sink_mgmt_slave_waitrequest), //       .waitrequest
		.avs_writedata   (mm_interconnect_0_sink_mgmt_slave_writedata)    //       .writedata
	);

	master_export demo_mgmt (
		.clk             (clk_clk),                                       //  clock.clk
		.reset           (sync_reset_reset),                              //  reset.reset
		.avm_address     (demo_mgmt_address),                             // master.address
		.avm_read        (demo_mgmt_read),                                //       .read
		.avm_waitrequest (demo_mgmt_waitrequest),                         //       .waitrequest
		.avm_readdata    (demo_mgmt_readdata),                            //       .readdata
		.avm_write       (demo_mgmt_write),                               //       .write
		.avm_writedata   (demo_mgmt_writedata),                           //       .writedata
		.avs_address     (mm_interconnect_0_demo_mgmt_slave_address),     //  slave.address
		.avs_read        (mm_interconnect_0_demo_mgmt_slave_read),        //       .read
		.avs_readdata    (mm_interconnect_0_demo_mgmt_slave_readdata),    //       .readdata
		.avs_write       (mm_interconnect_0_demo_mgmt_slave_write),       //       .write
		.avs_waitrequest (mm_interconnect_0_demo_mgmt_slave_waitrequest), //       .waitrequest
		.avs_writedata   (mm_interconnect_0_demo_mgmt_slave_writedata)    //       .writedata
	);

	demo_control_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~sync_reset_reset),                       // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	demo_control_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                      (clk_clk),                                                      //                                    clk_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (sync_reset_reset),                                             // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.code_data_memory_s1_address                      (mm_interconnect_0_code_data_memory_s1_address),                //                        code_data_memory_s1.address
		.code_data_memory_s1_write                        (mm_interconnect_0_code_data_memory_s1_write),                  //                                           .write
		.code_data_memory_s1_readdata                     (mm_interconnect_0_code_data_memory_s1_readdata),               //                                           .readdata
		.code_data_memory_s1_writedata                    (mm_interconnect_0_code_data_memory_s1_writedata),              //                                           .writedata
		.code_data_memory_s1_byteenable                   (mm_interconnect_0_code_data_memory_s1_byteenable),             //                                           .byteenable
		.code_data_memory_s1_chipselect                   (mm_interconnect_0_code_data_memory_s1_chipselect),             //                                           .chipselect
		.code_data_memory_s1_clken                        (mm_interconnect_0_code_data_memory_s1_clken),                  //                                           .clken
		.demo_mgmt_slave_address                          (mm_interconnect_0_demo_mgmt_slave_address),                    //                            demo_mgmt_slave.address
		.demo_mgmt_slave_write                            (mm_interconnect_0_demo_mgmt_slave_write),                      //                                           .write
		.demo_mgmt_slave_read                             (mm_interconnect_0_demo_mgmt_slave_read),                       //                                           .read
		.demo_mgmt_slave_readdata                         (mm_interconnect_0_demo_mgmt_slave_readdata),                   //                                           .readdata
		.demo_mgmt_slave_writedata                        (mm_interconnect_0_demo_mgmt_slave_writedata),                  //                                           .writedata
		.demo_mgmt_slave_waitrequest                      (mm_interconnect_0_demo_mgmt_slave_waitrequest),                //                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_address              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                           .write
		.jtag_uart_avalon_jtag_slave_read                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                           .read
		.jtag_uart_avalon_jtag_slave_readdata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                           .chipselect
		.lcd_control_slave_address                        (mm_interconnect_0_lcd_control_slave_address),                  //                          lcd_control_slave.address
		.lcd_control_slave_write                          (mm_interconnect_0_lcd_control_slave_write),                    //                                           .write
		.lcd_control_slave_read                           (mm_interconnect_0_lcd_control_slave_read),                     //                                           .read
		.lcd_control_slave_readdata                       (mm_interconnect_0_lcd_control_slave_readdata),                 //                                           .readdata
		.lcd_control_slave_writedata                      (mm_interconnect_0_lcd_control_slave_writedata),                //                                           .writedata
		.lcd_control_slave_begintransfer                  (mm_interconnect_0_lcd_control_slave_begintransfer),            //                                           .begintransfer
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.sink_mgmt_slave_address                          (mm_interconnect_0_sink_mgmt_slave_address),                    //                            sink_mgmt_slave.address
		.sink_mgmt_slave_write                            (mm_interconnect_0_sink_mgmt_slave_write),                      //                                           .write
		.sink_mgmt_slave_read                             (mm_interconnect_0_sink_mgmt_slave_read),                       //                                           .read
		.sink_mgmt_slave_readdata                         (mm_interconnect_0_sink_mgmt_slave_readdata),                   //                                           .readdata
		.sink_mgmt_slave_writedata                        (mm_interconnect_0_sink_mgmt_slave_writedata),                  //                                           .writedata
		.sink_mgmt_slave_waitrequest                      (mm_interconnect_0_sink_mgmt_slave_waitrequest),                //                                           .waitrequest
		.sink_reconfig_reconfig_mgmt_address              (mm_interconnect_0_sink_reconfig_reconfig_mgmt_address),        //                sink_reconfig_reconfig_mgmt.address
		.sink_reconfig_reconfig_mgmt_write                (mm_interconnect_0_sink_reconfig_reconfig_mgmt_write),          //                                           .write
		.sink_reconfig_reconfig_mgmt_read                 (mm_interconnect_0_sink_reconfig_reconfig_mgmt_read),           //                                           .read
		.sink_reconfig_reconfig_mgmt_readdata             (mm_interconnect_0_sink_reconfig_reconfig_mgmt_readdata),       //                                           .readdata
		.sink_reconfig_reconfig_mgmt_writedata            (mm_interconnect_0_sink_reconfig_reconfig_mgmt_writedata),      //                                           .writedata
		.sink_reconfig_reconfig_mgmt_waitrequest          (mm_interconnect_0_sink_reconfig_reconfig_mgmt_waitrequest),    //                                           .waitrequest
		.source_mgmt_slave_address                        (mm_interconnect_0_source_mgmt_slave_address),                  //                          source_mgmt_slave.address
		.source_mgmt_slave_write                          (mm_interconnect_0_source_mgmt_slave_write),                    //                                           .write
		.source_mgmt_slave_read                           (mm_interconnect_0_source_mgmt_slave_read),                     //                                           .read
		.source_mgmt_slave_readdata                       (mm_interconnect_0_source_mgmt_slave_readdata),                 //                                           .readdata
		.source_mgmt_slave_writedata                      (mm_interconnect_0_source_mgmt_slave_writedata),                //                                           .writedata
		.source_mgmt_slave_waitrequest                    (mm_interconnect_0_source_mgmt_slave_waitrequest),              //                                           .waitrequest
		.source_reconfig_reconfig_mgmt_address            (mm_interconnect_0_source_reconfig_reconfig_mgmt_address),      //              source_reconfig_reconfig_mgmt.address
		.source_reconfig_reconfig_mgmt_write              (mm_interconnect_0_source_reconfig_reconfig_mgmt_write),        //                                           .write
		.source_reconfig_reconfig_mgmt_read               (mm_interconnect_0_source_reconfig_reconfig_mgmt_read),         //                                           .read
		.source_reconfig_reconfig_mgmt_readdata           (mm_interconnect_0_source_reconfig_reconfig_mgmt_readdata),     //                                           .readdata
		.source_reconfig_reconfig_mgmt_writedata          (mm_interconnect_0_source_reconfig_reconfig_mgmt_writedata),    //                                           .writedata
		.source_reconfig_reconfig_mgmt_waitrequest        (mm_interconnect_0_source_reconfig_reconfig_mgmt_waitrequest),  //                                           .waitrequest
		.timer_0_s1_address                               (mm_interconnect_0_timer_0_s1_address),                         //                                 timer_0_s1.address
		.timer_0_s1_write                                 (mm_interconnect_0_timer_0_s1_write),                           //                                           .write
		.timer_0_s1_readdata                              (mm_interconnect_0_timer_0_s1_readdata),                        //                                           .readdata
		.timer_0_s1_writedata                             (mm_interconnect_0_timer_0_s1_writedata),                       //                                           .writedata
		.timer_0_s1_chipselect                            (mm_interconnect_0_timer_0_s1_chipselect)                       //                                           .chipselect
	);

	demo_control_irq_mapper irq_mapper (
		.clk           (clk_clk),                  //       clk.clk
		.reset         (sync_reset_reset),         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (~reset_reset_n),                             // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (sync_reset_reset),                           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
