// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
cNpWyCZ0BmZsu6Pw6Ptl8JWKKA8Pual3ZcREyT2tvlVWYawBvALqzqBpRzPD3lGHRVDVieP4tfT5
pT2jIkibYfJIp5zQjlu69BpzHvYC3gw4FA5IojmCpVGrZiQeqVvz5frXxFXBr7d1owyuOJTywnu6
BY3gxX8I7kOi+e37A7zHRuCV5rVr+GMH8SOgjSJjzfdTFsK7FJzhK5IAkrdOIrh4bFDDoYHVhg47
bBK7XMxfjVxrGChgOsTVC5v8WbycdWYB+vr2d1cAsoI5iEanMzLwf3XpfW3gVjx2LwUnAMoXMiYP
wNcoJzVSEg4QwfD1jruMRUH5N46PCgvk+X3v0g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
3bIt6wGwdpl4GcUk5apu6itcuzeCSPD3F8CD0Ia7VPU0C2RoZEcfQ/bgZcOjZPG5c7PBKQmGm2rz
2+vG337MuQup25zbbvTrpLkOAtEFK73Glwp/WOMTMDU8nbDBQuJ8zd36b3blbYUohy86VNeqMcGL
rhg44R/dldB07Ou9k+/xpAc/lq2f94qgXNXtXqTQeBquulhBGQKuitE9Xb7bLVnUg9LZXSEjlnWm
HIIVTPDiCHGYm4N/Rli4Y9CiBCQR3WalNGRkpTuZgxBrM1lrQqfRkEXyJzgk+3B3ReAt2RI4WsB6
bxzMlDjDtU5F04xN8+MjxSJTAM4+QgxuczdxUO3BxkTsijdjddo18OoDsT7OcHpwztq8m8gXdOlT
Bab7mG9Vej1xUlrg9bXap07tDBZkndsG0RUpQXMiLhpAkMhkb+/MHDjFNK5Z2MofFH2Jo8/TuE1c
0F5CTX/zFoYGBX1xZ7QaWmM3GVSAh5x1gMk7/VnfFDu9k8R7GySF2sbkvsIwjWGrECOTBtE945eq
HJ85qrk3v4Iqv01cgzteYdHOXlAaLYSFpwi/hU5Dd/7iSSOxBOT108d7avPT7qDE5DRmXQsIV4Ud
kPVxAKGWjPnQ2brMfouBAjYJiY+qaH4hwa+nyKmoKNoX9bSHVGpe80A5MthSe6rv1smYsFc3qmWg
r2CB/5wy8QLaGuvM6B/3x4S9ZKg6TAEjB5XWIQH9E5Hzs7dKFiS3nUflhf4Yfa8B+TV5z3Vn9nXZ
qPyr69mqlbxc9LBo0cm8h+itqhWyWnOdG9qRPwzJ7frpDRLgCBBYCQtqsRtVppswefAh9rv13iWi
oOT4vhRM/R9wxoROCEiU5crFxgoiCXscS/Rs3IX7lQvwte9LbN9Cn5QbWAR4mwO7zcAgJUxxMgkv
QTb4XARD7P5JxBpetDTiN7ObTLa861GCxGQKnt358D9bdFimPND7x6cM2eOgzNv/I9JeYpA9PxFC
qNvVGljQw6QChSk+zETpb83Z8ba/EyvPuu/EEiGzZs1/GSaR6x3ZjUK3kvh1oA4SG4K17guUHsjM
OlR28kMblOsgrVDjGbZx93O9/haZq/Qt40S40/QMqlJlQ7nS2WCcxIw+yBJpALLW+McpQZm6e2oB
q9TgBhpHTmiqI3DK1N/vqBUS9ZUytTZ8p6iZobtVnuOrI6Q2jLITc8gQtGnZ693bG5E4cUE8keGr
oGJUD/hBq//cBl+zFNr1AoyZJdvZ+V+ouThMVeQgvIiZHjd/+RGCPNtRK6c7g0KL3lqu8HSWqart
2fWsEztJnp5zdJWZpWwPcMXK3SUpaWVlOOdyQicEGLYTer7uF8NYZSPX2m6TBjfnjN076FphHWBb
JgxTVi1K8fp+IOX67229n79B7WMsCn1QQE8omWm6fLidaXeobiC7jRRB0rOp18X8/9j1QJwKc1oD
KQO8gV/TJlK4YLLcHo+yAHLEzsdNuGF9EGIdA0yxBBTaAWv4/fam+gNxqkiqGElQDx8F+ljtwE/k
FcyT7TD2d6jpyvXm5qqf7HCJozyYHVI5jm34z+cicAPaIkHWM8wZABikHGY7DTOrnPgT3jGynMiU
GSM9c9a+nKnr0wrsbeH/sChQHhr3XoA7QKMmGtLy6JuSvho+DYeftm2MaCO34+7XEC6MJcLiLz9f
EJ2aWrAVYp9f55CLbLdbjWLhngF+CqFbLahWDfizD3Uzn6zLViOVIR/vTVQmA641iufu3rnS/1x3
b9/aOOmu7F4SA2zd6Nv7EwzQanPJ8SuR+qn+3V28eAWQF/wCM31ZV2w8ssUXS7sJhIF5r7qn/ZAS
8wII7a1MT16QNXBM+3Wg9lBRnXMJd/Trm6GtdPPT8WyC6+XpADX7RoGZaVU9ZRTbq1SykhG5FEDS
ccmj2HxaKyRgX83tfTerAMJsDyN025HJBdjEKnfn5UXvI5jlI2PjtJb/P+SswgabxjBlcF4QReWh
6aTs9vqJHzRUc4S/jmFKToY2Av4s0AU9WLNaLHnMPtkbvzX7OM9zQsJmewKmlzI7JsBQ/p2SfiRq
joeF0d8S5lYbMcyZOgBbhByW4Cp5kJgohXxaK0y/mH+eQiFg/o83ucR3Lk0Lhl1uXSac1sorjCAH
/o4kW77kNGYaslmXFXa9563EakJd1mXuyeEcrLLs+ZQuHwXj6Kx1e3zNrB1EWxz6z7cTHEEF2Gla
cehTrm7KRd7wCmqvAkwYlBrtk4CdEayRFOfSXqSa3muIfFsVfFstwSlFG81DRwwNONqXE0/0Idsi
lcdm6arPkEkVO1B1urmRCqHqvbgrdXXKXqgr3IKUR16EhZ90PSwM2NhOBmfqc76VxggnRoLV5bVR
YmM6RF8Vhm6Tvnwv7un+Y0MY2f9BP7MQkxK1IxDdN6nsoLF1ICsmxj2SNQgtP/71O9ySBC+xKbjt
4NMgvwPDdnld/qSONIUAarcKKHpcPDMVXD0BPirQJBsRwsJKxsdjTMDJFpVyX98XI3fkNiONTq6r
iqxeuR2RD4mcoxFw6NA/iqnqMQPjMVpubperArhKOb6oNukse28YiQo/d4JFAmsO6M1WRRDEHR2b
WPGbJuZvbKNLFA9v6tIb4o1xh3cFgCIk9yL47h/pVwjQl0kdvIj5tb3r7VvuZvOuiXUG49P+vjd2
imPAMj2o/lLwB/6JlAeumBsXskfKtJ5f3Ie0VcApyx0MgNMDRP/IXvIqwhdIS3Y4zDiQINZXA9LW
WzlKADZN/sJxhzXWp6oOl51ZOdNS1bzSlnZYgTd+7Mj8xRQZD8yuLt9bku7YzSdAf1MrrKNSrDa9
piSbXZ1NqIqGdCgwuGhEWPfZxw/GGPVSWmSfq5kzoBSJprYCostcqQ+Z5oYizbA2xo0O4jW5cOBX
7Xb36ome61K0eLdWtC5myYGHp4kLOROvRu0KZY7Dn7WXg/wORsg5WQZPk8UD0JGpr7DrDMnYjMKj
+RdJLkeX1r4kLQWqJU7KgPDAmWLDo5yvdEX285l1bzCQxt0cD3BKanE8JjVmaBOl6/rKAqhKYBS6
YlQBakI1b2yqx9zDIbbLS450/TQVbVTVgGo0xH29v+OJFFGDyCMoIQkNjhVG75gWKnYbJKDd+5YJ
XThE6mio82M+b2me1qlrSPHV5IwgtuuwT+sRxXh7ZMhEB72mxy6s/rI1fG0eG1aQ1CEi3NUrt4dh
Hl3wIbnezeVCwKyhdX4jL/mzT7TjVc8FsXs+NODYTuRpNQJJjJJyUrjOttfzr/pduVoa2DkHbdgu
oSPQ+ePfwd7DU7BT3SUiJLQn9HJ70MUltVcR0gc1WWXetWD2YB/3qfNS8c2LGWe0ild0BMr2c4vH
cGSaRK7RRLp8bwOqatbdAYxdKpfjcsVNE/7yichTBUE/9x5KvBROFsXmIE0eIJg4ea87y5MrEQwl
wr97mRbKH4hvflylFKaOzun2AfJWRiJzttIrLnhWvqyM6Dtk7rvZ3/FZ2s7yDv6MzPcFlHapO6wR
lAwthqQHnZu6zHO6G0hSKkiUByiBIWBPwDAMpl/XbhuDHurfV5XTeg7sdgoThguFm3PfOUjL0TE5
1Spqqx70NsXD2Yyl9HsLKhLPbPoT2QS7WmPSNjZzArKqVhWau+eGHf+gXrSnY7UpzijAFKpySihV
jkutuHbGt+9DbkF39zq/T2MDRMXHu6dPAH048pk67HBmdcLLVZA38gsRxWcTdzeysNpt181gRLoC
8JG59wMewTvUZr5n3gTw4Az7qH3PQjEPiu6W8GeKPIppp2bbfK1A3Nrv0JPcepKQ5FexClP8UuWM
u6awu55hA07AkH7XzHcIYmC6Cq0GVRMbJII5biQz1LlYPSCZ00OyAUGJal38GehL1JPm4F1q5SnO
mQxtQJUCTs2QbcN1Yjtrc61p8+sva+LmbnvrUDvOSsGr5GqLXV0QgyFxslAnUyFuRXsPvS0mSzdK
4XSQ5nErOSgw8917IAZaibWY7ODspSujh4IFIvNOdKNabgE+yVhL6FRYW/L87xLDRv7T8lm2smag
JuF1+omf4ZsvbDV+2zqcghKAc/4+qBSHNXN2HofJG+jo5gz14PYRbrpHmGvBeeMi/XSzKKl98Uaw
Fj4rmfya4eKp9iK6QDuANYlT7zigNSEKn6vGCcD7Nbagw6CzRezMVd/0s7AHgQIAMOb3Ko1ux9jD
6lApCz+PfRY0Ts3vh0LLnJCMav86Tml1FtnxUlxSYreq30nF/Lq0ZJ4CapNL9SjcYCODpgZGuLa8
N4bXDSLW4+c4DlZmY9yE/hPNjZFBeQG9XiVJqe7LaNjlPCNV138fiYePAKnnyzHZZXXeivJNs6uE
P9SwjKd347jXCdqzFwfWhD8Gx2TEepeI8y3NdeO4MHHrwRTqyqlciDnNZqMuxLIlBqxUGBehILgU
wi8yRqe2zUDijZTpSG4a6InSoNQgjzqYPu/2ZmF51ZIDtzmEmiqhUQNAHXeH+8HsqkVUNg9a3paB
eMNQEFTN8uhFw8Sm/SeLDBWJ3ykAZ4kZmnZkCp1S+0appBM+UvGoJYdtA0tMoUGrghHHII9KAgKN
GDsf6cVB1kvgYQhO1aSgJ/h8POx7Vk9clY7sYgkcTVYLJAIyM2sV3fmZEfBpxsx2qjrvVZb3KZeH
1bXzDzPvD/PSc3VTb+EyUC2nmMhkdM0hhEnvwHKJqe5DA8SBWJfYH/2XgNFVAhLjIvul09fvEv/3
ObzklCo62LLva+UB+mAsPwZ/gyiPcA22eime7gb9jI0E0z8UZgi7NsYFPM3sbt0hqg8/Rgq/qcT/
1m6zpHZSLwkkvzCco+U0m21BbKbDC56MGfXkbhnKI6aYSHohEuEhT9FgPGOw+4oG4Cnp8tFFscEZ
JlfV0acbVwkLOcFC09vyX7lvMZQmS8v1hQIehTwbWoK86WugsYNal6cusFFCmSUfeX91ckMCZxB2
7S1KhEC+UR+XZbv1fWoCkczRjqdj6qvbKZc9TkrjRAdrqRDEkC8GFvFXA1koldolHbahjzIfbLC/
PEjplz+MXB+4JZ6Sv0uQtbQxV/5M9aklviIFnHTcAZVmANB9b8/oPWKU36R3z4fKgbD9IVQMLuSp
E2EuDtn035r83R4dBrItj19p/eufOWXuxAsPP2stEuFBhIWND1ICItiIPIUBvxKalCjnqR3IREu+
YakWWo/M0comYEFO4HdgcXCXlZc7OLoVYwc4xusX/pbzXvKF29NBnDZrC5kcx8/Uc178gFSt5WXj
+6XCxtFOesmqKDafPq1AmoZj1kwHWXh4z/zXyfB+1ph09I63YMAkJBr9gRQcN/QCnVg6XdGGX70p
6tiA0iQE2y53iZZEBjwlSdhO+gjwbbFcIzrQLJDHT2iAaqGl7o32o1yoP9stfWQ/ZluTli4p0zfa
qwbibMYR3zd7Y8YzyytUEXD2J/56461MsqubFZaVUEg+Ejuxa0Jxpr+rAoM2WHLTEcIESoZan+Ta
SYO7znJR4GWXivpzr7NsfBrJ7SFO66HG2DLa0U9IkZOE5OCK7tQFbznPqAz/LiRiINjmYxtcmBZh
NivyahBwfgW46m+ZodvnQ4HRpVpSaE2Q4oiAnxHuIcESUOkuERRBzkZCsy6mjjVmPbM724tVVYpo
oQzmE8pWKBr/tY40UEvs/ptNfLzF1LsaYvlE/BXHz/4lkZ8GYmAp2XyWmeq50jCMH0rAYZuFxJl0
SR/qdY/YRLLVpdHn52CnYM1og+9F9p3sJN/6B7DXWbud8zW346onVUK6Y9Rc6aODiKY6ujq0O8Xk
E2r6deDT3KaVmGMTvnBBRPqHZX+duklVO+2/gu+Xtbdui0Qj3eD9Y7DSly/5rkgc9o5tqbw/ONuo
nTiHNA0usWjjCM6BBwxdHJhRqd4O5WUPizh40iD47OrTQ8BGnJuqmfWsauY42DS5wD2UtylCaQpM
hw/eKWUGdOG2p6tA/074MGhb7IOcYdpuQkBLybjzg5SEU2qDG3uYThoKpqKxeWMkOwcADSjT1FdD
szu0lmo3iZK+4lxZUccx9o6VrWOszMW96tSNpn56fYZIURB71ih1KMRTof62rKU+6fAGtbI69Fwi
0is76FZqSMPRLPFOZnLKHyRDdvG8Xp1MxM6ptB8jcmbArRxJIy3PBGGpjmt/ZkFvWjt9qtXZY8mE
y7qXa6z5Po39ys0zk5R/a1raKZB7B4ClALOPWu2NNH7C/5krwlp876vtMkabtq/f/RkQUU92IuL3
hkYQjcl/d45/c0I/59HY7o1EEGvq67KVXaRJzHuX2/Bh+fKe67LGDtwfz9qDH22oivPo5qhjQWPv
9RCE3cKS+Wa7WZimw/kbAgfg9X5LvMXLffNOpHN1fqeg1O8FVmEb/vQAjxrtfudGQlgP1K4gORMk
ZZpjCk8keoWs1GhsgFXC3EmiRDb3VyNNCm6iLFnmirH2lkmzGPwMgQSoUSocFDErXDUWIvqDh5iR
Y5kv4yOTow/dbgZu40yw+QkjO4kRnyjMCx1jO/9Pct9Vy6jCLvqtajMo9GI5bIwV9+fVst32W2sq
LdLT84FS7xqnLVKDHT79q8VrLAxO1urpiwSYWbnzyRxwE3kZIJbbcYJ16Yv+FGP8eGmCw6gwAkvf
TeFgrPiNu3NUL01mfM7wLAHHo+JPvzZX1oHnQvc1jEbFfvkV3FQ2ZzQGiOUJCqQ3wuPzxrN+Y6/o
gkkxjBxxiP103bR5H7qJZPxF6WyqKvMQS6X4kaIV88eNxDVYR0AWCWT78mJgBtFcxz8fd9SL+iJm
U7vxgEmJRWYerhmSFij87pqT8mHmTlfRtAgXyMxePwOhsafOFc8IfLvM22VjLS3UoHvsoQZLyCza
4C7075I1NxVB3iJqISY3ylsLksua/cVuRK7Th77D5bMcI9wI8sTdMDRcxsYJyVDq0BI5hIqXsmTd
hDNW8rm5xknqfB7JRMpEotdktbBjKc+s2yCvspyH6BHAlOIchJp1PGjvWPOAydmzPd+UaZmQXgIT
4G0G6J9iMy+F0EUT4hoUYGVcc1VRIe3kjcXWQRbV0xLrwh6N+OBbqT+wNlMDbnZN66n+1d50bIxR
my40vFx6qAexf24Pnc+tR3CfTvK8Qiep7wTRNrpEmv4VEYpCAxY2toJshwDnKLjuqEL/EJ15lmDt
2sGd5qbjdvPSIxM4MUlEqppwEs+kkJT4WF/FgJKD4gnMXtYF7AzTvyM3QF61OBHIE4RUyT1SAb/i
ZI14kl5IMdPq192IzZTrqzhaWuCJLGAKr9bRWXCUVTdbc1lXFP2VoKIITNgr7092kLzjwAGFNq49
bdYiZ7jfa/KuV7H9cpgQ+dM0neRmq5OPMM3mx7y8AKHIqWi8nl2z9V8MIqHJfzH6MsCp5YnkReGM
uLNJMfMb6o1FX8e1qPBikNJCODIppNBadJHSIJuYvgwE686j5IXSqI/HGZhS95rWSQxhQv5stzx6
jHgSpjv/gWhmU0depBJolnAmM76lPKn6hgKn/87Q91ucao9qISeNESjp3fdZ+8MWgzETMQi2azfp
0eTGJE2azu8OiWNJvbbWR/gpRk20/z+4oPKPOj7HEugkShy8NPVIb0zyuX6HWWmyPnZ+bsHUnTKe
El6yzJqmwDKfImfjZPuKX6OI9e0kJrSHdXl3NUqsm3OkGsH2PIqB6qxxNorGfRrSbDUM0hzDOGyD
CXUGIZq9qOMrzE3xlbp/RLpWfNn1yygfkBnOezd9RgwpdA9nuSIpJ69a13yuQAyFTEgzOz2TJ7NY
YOBk3ik1RzlYATrCE1DqJiCPCKTSEuhoBe/ZBmClggscfBZuKVk4H3Gyj0kxylrmMKuvq1kk8191
UoetcmBB6RzMeFcRe8gc3H3xiqnwSOOTBr6knZvzQnWXK5qOQLG2rV4oxK1myGZUBMY8iFKA1aN0
frk+t34QWEmGpBaIqNImzZXHOBXDFzR+T1qp6/HzIW7zaNf3n7qVa0bR+2VV/eMAfTzVpNXBGJIL
lWN2pq5CK7g5UYENI9FM1+PLxT271tqcvMohk1OeYP27VvKe/o1vSg5xCUbO4LihBwGeuFhhjU1n
SdhORg1B/gnkseCG6xGeS5t8/CJODUpaMSJ8OaJWJccjxGM2faZVC5p1XWnr+dL0c15KsG/OTcJP
oMGjS6cBXrPfWbx9MMgFxWasbHWcj+hlYHqsQO63FxW+t11lgAKQqC4f0uMKdA06YYrpf7W5ae2T
bLAnMlKlRsqrBL1FawR/uDHPbWP2A9Lt6SbOQHTQudgIssf+hy1weXrlreQvQ9g7Mdq9JBpSBTrr
xaP0jTUCnqvAKlNDs9pIk9i8LeAuljKD3l1v/n7t1jzecNEhUWoL8KxOORDV00cjz4BEPI8mwmnP
ev2Xi8DvmzKZZPUgIuHxCtRk2LBBByBUXo3iYkpgk8XdA517o+/hwjJuoRhi++sm3bt1g/WPKzV1
PwbqrMVPp4wnaigZue65dwDgHORUqvYEDYPP9OpgpT0nFAK2ROqfRUebafZ6SqEve7N0tCIV0EoO
3URVcweglYBr1MzUgbEPwS3Pbqi7C6kYakmtAu9bQtaXbU88LByaUCXkGiwu4RiFsmA4GI5n9Jh8
2M02cKDaBYu4c6cbGXVxPt3P6IOI63an6jT8ZG59C9Slov5K4Evl6iRdemy9hZvij/lZIpgwEwD6
oJBcxyc3FMcxSoXq25T0z5SFzMGmVwCem3ZDM4R2hyeohSHLTXioA4PV45EW/pS0ii1VIK2Hw9oJ
z64eIrepqCOufsjIOOFVbP6ml7Dz2CplKqS61WqLbFYEoWdJxy77SquCwcrSzpImeNTZ3+k0RfTK
CZmL3W17iU6+VBZ7q0K9Rog132soSm+jW45C1OWxgkxYbBfz/pR3eMfBV39dx26gcwy2uRYlw3ed
KLicyBZQ5c54iJcCMaubCx7RFL0H4amB4Y0bWvNKQeEruuWnqM7hpHyTsENREnekTAqx5LuqU+VU
EbARVlhIRLeV873SBe2rY7ybHYp08nSajrUnBmpuELvnBXqLqcaJXrGo3Sm7mY3Dpxiav2r5JLXg
kqRx/cWmWnOwZ0UGNpky+z9b6VrRCWJvoiylL7dIA7BFXS2OHJZQg0v4tjxrsZJwxPw5surgoo/s
iahW/oyWkHOc1A/xUCrk9uWQd+Ks2eH7TszqEgkBWPDe2TQlQv+8gzBLQM2FW/fXjvVnnMx0IPzn
4LIunMEZOYnnDKji8+5GUDTZT1VCmZQHDz+3Zh7X1myLQIxJk6BhPL/shlsOXHmRGv6yTwpDREOn
JNg5Mhe8pX8LaGd8mWzrwUOIsSky/L76Q5dWlrL4avoaQ2GBeULZTLH2SpYNlJECxDyDLODfk0Yv
KFMiuPrMJTtYNkXNzDFr095YzZTYBM9PwpZ1rdKZmusOylI30WMer/pp45wjoREfHGnY8zcuUpEh
som4SOtT7Fwe+BtnB7yovBDI4jJlHmgteJfFQZgjjBaRyh81auBG1kGsNfp4PBg0ILV0Lbgp9R1+
kjHEWBw7Yq69DE8Pc0OXeYdQ4yWNnZCIEtOlI1AvmqCrXAr1kZOUl8fT9tQJ0O0yTNRbia3gSP29
4N3UWAMd4+CYY/s/8FniYJdoFxms138xKRWtL1MmYUKPxgRIW9vndus2Lw/nA1yUWTdtuIvZ6l3g
uQxqPwXyKqA4nuwAaK0JUeo9dGZ0eCsgq0CeZPYTDrdu1YqBkm5Nh/JeFxhyNdycBrwNoVQy4cKl
5Jd1hJBjr1gZJOjIoHy3S6pHvszI69nROC8h0cvkoFcDYSAo5MfLW6jHMU8Wn5QDr7evfhizNXTf
RsKUEDTmjP5oALi6eLMC47tyMB/JMySxgXWRHXerlwOUhHoSV2br6ieqMT8j84xnytuZDSpUPYSU
haMsZvGRAAYCjwHrNixxTNJlzuD2/GB22o5oZwPBeZFW8brmoMPzeazz+VJdbBonfIAWyC7n4wxK
8JToRCF+JV/0d1h6UFyjz6PwfKlL1sC9sIMwb47Lu0gWRAzluh7ZqJ2NCMW8midMsAprMnnDdxBr
SchF9oi2eX2Cwd5Y2QBKLpBqnEjqky4wxgg7KZ/0FjdfqDCSsqv0+BDVuAaO1LZoCdRjNqT6Hlsr
VqCejp8KXGlMSHm2BD4fLncIqrkE7KjQgI9HkYgTw5Ob8YK8LXf++ZtpBNqqjsZS/IaLKB+wY0MJ
aco/gC/G9ACB6zDBBIXBDPC72YPv7WVTxeKjBUXXMOg0hcbKkYmQuWm886iF3H/O2oNE01mu9hh2
jwFTDr5juu1wcuPDpEsHqiETLlCEndyNWY0b/K6HUJxzTaa3T+4fYyum6yzVGmlprZH5ISpz64tY
x04tINjRkb0/+IQHyjlPosca3Us+zZ0eK2UGQNzKHBaBUwRjGLUYy1k54mfie01w4Zi+qD1xqi0H
ndF3NPYBob5GM6q3aDoOSlFDNumdsO/iqR4mYxiGBYR3HM/jUlb3bvCk6auEGqX/2XvcwQGwxN9v
wp4lLMEomUJcOQgKVo46rRGgPEyZuJBWGmubrNKbVLKN5E6q3eb67o8kZ5/iDgiDukZ+xAeLEIIk
CYmC6Nfmlq44AnTc8ciOkwH2Lsqr4uwQVBgTcdLX6SwMfGGVVv2eq+9t793mLIjbDG0j1CylRumW
GCgSXMwsqUG3fkOQri1dxzPvorVBmEAB/zaQrCihPx9m0FDOz7CFL/DqFF5eXIBLlRtgiQwooWRE
TmVfZQgQI4A+P8tUvxNV8KyEMYqlQF69F8TUEh9s5p1aDqMW+GtaN+ur7f3vrC2Okz2RGD4M7jW4
psW/qKaxgBhux1Zor4zyU8ERxmVhSaruJZdPpudUzD9Z1xxE+UwUsL1qjYp2nNLbnqqKNxaKc6tE
2AR1gOj4bSyfBgxzxa14PAAS44jBPLjvzize1JKtWToPgMdwe5M+pUAFTWtWoaZukGdRLjnPAei4
PrfAgLJc9uGC3qJmY6xw4BwEcwmQKf2OCr943hJfDkhsPiW0y+EUJ/V8GE911zvQqJ+1rac8tiEU
5XsJEHBIsGaF7w1X9mUtFe/F828SOu779oAhCfQyme/s4022v2q5L1KoaMRIGxmpqx8Qer+WCBvx
8+TgwNxMaynmuzRvUBEoJwLxre1lQybwPnhCxN4ep8H+JfuAbWrH8NYKaJORsDA0DBm54aRD06Ek
anitIfgb3StJrhm1c/Qk3TB0tivn0jTHAdvmGgyYZRYrX5r2oOU0E+cccrP1JCAHxsXQ1V0y7ILC
mWn7PDqvXZeheN17HVuyqhaAUSgKDQoz2iKM6fa21rVEmU5HFBuhop090+ik+lZqNmraVEa4Q6fz
+4NIdVRTFtni19VoU6c/vlh8ntXt16o5DeNce9qd6k+IyVPGJGNaQ1v9k7EAYNC/NoPkFZSe+bTX
8cGFOlFmusgW7+D7c7D2OHyM8eEr2xXV31UuJ49m1F5tdKVItBr0NDuWvRtqmrJqlcq7bnVlsdQH
xYoxEcIanj9EEGw5sSgR1IE2ZVd2QFn5vfSLlO8Lr0FMYpjfjpD8Jw+6vmC2euHSa8rcYKILT4IC
yGJ2oyVznW7ikU9kT8LinmQJOaFBtCZjx7MtI/Qt8EjedseOB7cXbrYapsKK8y6JcEVRQnfo+ty2
iNUzVspUTo4Rc3G5qous24rHGGrR09jC6bcg+x9c7Vmj2zW3h1MxhHz8Lizyq2kMqAy4HhtWVjvQ
jViMLEoFKCkUhExLujwAXUMF3mFQr5tWc2NVn9Frl83gdwEu1dsO0efyp5YgThoItSPecRQZxaWs
hWmpZk/rr4zhEAedNfxphy6ueZWsLLHnqIETRtX6cdfdLPhFvz0MX5NC9ALvF44tkGBUAWrpXrJp
Qv/0VsEY6HMUbyh59NlqJhgco1DfDo10wYAgHTheJic1z6IZZP0XJpWuCoNSkwU30QCibCw6KO/r
XliCQbT8deohw/mQsMT6gk3K30bSioAaUMao2z7wgF0X0OxS/5r9B/ckyPbrrdaYi81ryA/Rv4My
FXfxBSs2/3x0bAmLAvEV/0+2PlDJi2WeSgSvt1CpujW+/la9hqqoJP7R63Wtvm/e7JfRLLd7CEIj
jNa+krmZ9O5R+3SL7jQNvhWwKup/f0fKvosUMDnNEBs7B3Npk4rfacRzNUw5zbd5ls45Ix9/0nSP
EmileHnbLgB8RT1FqHXrkYRQQvONRuFBtI9S72AyQ88LEOB+WVuzQVEjBY/WM0lgEu1pgNyl0NF0
FbyPgH3IVeEJt7/dDjoZ38benEEApA7UaTaaAjCzb5a+d77fEBQ2Hkm/m5u4mCL/jYNbdqBEkyEj
KOxt4ygb/Sup2Nw1G5kTCjlFo2tXCGtAdzXnyz/XcD2wc87IGQsChIJhATEZmHrjw8t5ofzL4g+U
MlbY/vH2mcmRFLJF7kIKKzHqBf0n2IkvF/Tm2yqcP/eLnvyS2uD9rE2leuT+Dk2/X83TvQFU9YAc
JfcBbC54VEXLQdbpDxeFCTj8g3NVEC+7FL0VfpJHOxEV400Yvom+jLNz7UaANNLOhov73SzzFg8d
6tsfATfoG1bvvxdI+bzDKIJPDRgC93b19R1gsjcHG9vVmcGc268T0Nn1SNeTSWprhSApL2MPWE1D
sN0xRplW3nH/Do9JCR69NxVH/ya4nj7XR3YCtPBMUm5jqgrsgpIeTZj8ibTNcheh1TLQEY3vflHb
0Qa+wQhr0U0CNZTb7BhbwQl4KTYAap+TsE3GVeY24pSAMiG/EXVIrH/3rl/+hao4EmIt31Yls1Nd
9gzNllR9a3PDggZat/3pAttsidElUoTTqPCypSZHwdZpEDsk/RbQpI0EWbDsKTFojgENdMBmZNzC
1t7RqK2YYX4+AH8juXHlC30VZPNv4T+iuh2nOMuAQ6yagE++G1gJdsOVWqx9L21O47zFbmmR+hYp
2o86tYxqIs8eqR8yvnG0HVidpq4dlaiXNShD3mUScEKzJTgp5X1yG3F0erVnQfjI5NdNtjauw6Ei
z3I/x0CyWfMLfEZIgoKAicIr0zUM0E6mBeoVyEabXsBO8CsrBqOgynLjFQKFEgeIDfJ+hXQZOM7X
4+zq/wjeYyl0GoCmJYlnutyAA1r+mUWYcQMYvq2MxqSVIFJDwutfHEMbR7wSafLqgBpFIsGNDMQQ
65pQvl+MVF6h/UDVJn/lHq0v++H27ih+vofoJ2AK59n/Cwe+26BLfzgg5DOAdM0n48A/lNyj8qC2
MKgh9Wf0XHkZbArvoyGl86AAIC5vxtwJi/L1Bwj9KdEuyRcRJjZnNzzuKaYM0k0lwMgFOwfKi5Qs
qt6qWPDGXBkl0vs+k9N3eCx2gxeIxfximv9VbnKU6JZimnjInc4GtRAe/UYEm4JvPLxUcseNt0Fi
Vm97wx2T7uZCIDK0RLdi+4LIRljzOzDOrHKwURBHM+LWQjelI52qhvclvwzskfk/xHA3HYgkmCpE
3nvlNQjnosD6DmDzfxyOKGZvVzscY/sszma9+PMY93wQZ9aP7PQTV4EmeZJpVMDvONE2Qh/OpASF
RTFkNjW90a1U+CBTTQiXNPwvUXtNuuwLKafAL/jNIb4a0BOGopYwHE9uNST7Gzi0VXqBX4XADtrC
GgrVIDATRebih2Kqy3sLWYJCuiXHNjBK4Ixj7eRQvMw8PnH+ltpLF4AWCA7V1p4KSi5i1UU8/XLZ
g3ghYo3HN4PfFkq2HYWUzwTzJAUSikCO2rPruKniSSAUK7l3oIXhf3fs3yQ6Xz9FBuGfw0jg0syx
Mw7HBW55BrlNUtGoCu2u0DsRLSoV2FDpXgv9tXRx9QSk2RYimziXKBZqA4cgBKtKscZGqq7Sb4+w
lJq3AIoVkwqgw6ia/EeUoNtBE3Mwhls4XDPPWnapHLV9mxnnrLtlvSN7Q+c8/avzROjtSbTPT0Ks
4Hc3EeL6Wxl4RYDOhK4H4fEzl+MViZTQ1zwHoqn09sriRy12+k9wZks51Zag6j+VvaFnMgjY9NLw
ei0+zmNAkLHaXTGkhbm+8gRA7nql/fk1ChhehPtF63QK2oXV+28Dy0cA5dOWbruEjtJLdp2vFzYc
JR1suYOIquDsUbtuFpkSxP6DFy/JeMbUJimP3fz1Prc8fBE6IGoDvj3ZQQL8IQAMDEJg57RvtyRZ
IxzInaPibZM5VcrU8zCDTpgZQN1HbDp9sdC3sUU47ov3mgsIDR8pzN+e9L5w8a03frNBQ64Z2UrN
jwSSiaulXM0+q7TxsJgBdgk3/KCXMiUGTSfzI/YhRhKoWYfYybv7xJRPnXUvWgXeJgTui9hBSpJd
RxHuiaTX6Gug8nh0Sc4Re8PbRhgLPJqzMnrq+0GKxU6GBuI87/Mz5LHOjD3qGmWeXqTxwUf97z0D
Icc16nUVskQEXkMenjcfZGhf5Np7PqgT9nOXuyJEDk21Bm59ETN8mXe0YNgth69+WTEkm8viZOgY
prt5jdb2Jfa7q1+fD3SJctCkO+ZDocK4JgLshXOCvLzWzIU1RNJj5HCSHwfr5iaxSFUChCx4yelx
qfmObnFblbMU/7deC826H0wF3pU/ErlQgxkgYXwyK4nASrmeN1pvJVh03xnaZtVpRXSQ1L8aY2+r
gsmfTQTox2MB5UyZ6p8LauvNQpH07FS/QMC35IUZgzMOumHX3sLJOtFfr/J+0TrMVanw/A4toQQu
A981pEYjnlAEUt3uDNoFxwU5yVTjXQmnsfihpygS0D4O4vFHmJ9iBP+BJ9iZKqGQe6RA6689SEea
pKls6vNVsmVJxg1LrU65cd6JlZCP5P858PbfO8J6urNDI+xuac3Fh7Q+tWtdwmFhDg088c2ZSHnS
Up7E/LQzTBnyn/9B5kX1YN0jgPfRaOSXPGCNCBKfZ19UaKvPIGt8W9l8W3ZIrGkfwvFWsUqQiwrM
VXy/exqc8+mmv6clXQCI1A2USMS+7M0nL4eESjfGwRC2v1tNE2m6PpjATD5m201+z1ehuG5/mOKs
E9CtSiZQQFKKKKKlTrasyeBp7bt1bhgzjY9fEIvsno1UrAcQIJry6nSsJanVk+plmFiNfj27A9T8
VKFAAwpcu3rWy+wx8n6VNWqQDDjUrrUGi+/FgJ0cayILbDANNNWKtz0ykStSxXBE6TP8ND+h+G9a
ME2c8XMKGD8x1qnp9HcEVQwUyzQGtWL+jwy7vuXKUPetonzfaHotwhxGe1vfq0V1PKQqFN7nmrAO
aA7b/h1JwjWnlW+LnFxIHF92+YEaFPjDu3jpKVOxg+akad23MNA7+erP89kHvlvVRyIw+pwPHP43
del3LMxVc+uGyBJjcz/D28R2OHXKfPig3jZUoqEnC2oGy/ES7ER0mj1Zls7OrgGXql7l/5PytRRk
ZIOH0UXEnYQA5BySDfKx6QJ1icZ9VbLO3L74RCABo4GGStZ/62rlbSInHtcA8sMNlAtOjdPhkoNr
HITjIgCzWlS8napJeZdWQ6uy+F8p5jFXvZD5l3M60ORL9m9URS2XxJCXnzS2+1us8VTUVRsIVZ8V
GfPdz9Pe+tII3xXDIcAGI5dzHDVT/i1t3Gq7DHrM1uRmrKcilhmAl0fWdZXl6Q+V6YaQ8NVYMaR4
2CSz8DUiCskk+5CLc85abNXNXSkmod1HH94KDq9eTs1kglSbDPV1IovV52zcuCrQMVsTTi1FKLUE
QZVZQ/06Ja2Ld2QCK2VlKVTdB0lkdEQHBnT6R10BcC1Qs857jyHO8MWRtRioshRxRMboyusrhNyq
bLgXWEUWyl8rGP7P3CAZmhXgR+G/WLY5hXGW1wzeHgkpwyomeulW1N86ZM3Rj3F057yIyJxexEwA
g+DFpp6suUeaGqN09AYRuFrW2saMDqm+9z24XyLjjBlWS5XpaKA/bxIjjNaygtf+jGGj6fdFdbmg
3uNhe65oRoo+4o2rHYrfBLt1bBhhIUeypLrs5mPQKnCZU+6nxX0pDNK31/2kLau5GFSL1CG8bzmG
qOKQi9d6A2sIXaBmdl5a+2YEpL9UDWmjv/nKmUJOOlioyyz8p002vNszwR/O4ws6l2UA7dZp7Mxc
cLNp+LjXlPF3vfdxZ8HJyaIC/XWlHL2MwvXlmLTwwsYiDG2Wl0s/IsBMGoinHGOLBnUX2o8is8rM
fXem1PtjnxcWdvUs8eKBGxONmK7tRf/Iyxdg5mL5TUzr4yCSemCEHBb8EiPC3OHTyHvASoR1DixV
yHWJUex1640OLDmPCqgzvpgR0K2EZhlcQvxbwtyNJeBGiBryzf4JqbL2T+nofaIukQRU/VfyZ7bj
EjgsxPJKH21zn7+1UE3ECw9qZNN7D2a/mowBTqKeBwTbUVS04+TSdkrJCzkfFq92RmeWTzy2F8Gs
eodVnIbA0UlgyFow+3ArlIRK5kwCQfm2TdcTSefsztGWEtwh1dNRrzUvjHxAmV1XW14ywxNOTEzt
I2HbSW7ryOLp9lYGEiedwv5HzhdXGRCw/hkn2oQx/LAYvVB3SIX4+NCIOyi/OLUlIMXn2ZZNvfLc
xK0nXngTWdChebD5UUnXVLT92E2hHW4PNcCnB8bC1HrG/7w3yah70ypIMJKC6gagYBdGj3aBJMFk
XwO7+L/CfxsBtTGMSojsxnpyyjzC8S12/9h+q7AN1DvKe2sRcwFFkeb9dnF67ZkdwwzVxRQhUdia
YtU2yI0I05QBaEOEYOooE9ryAoUX50rijupi65A2U96hFGr9NFnXOldVhsTOjpxCwTe4FwDM7OJr
THFs91TIx/g13xzxBNzbGtbLj3eIhyQpk+LTYJmUMFH45tP+H5AAFSoocXcTzca4o8pMD4+dunq8
nJoPgfO/FmQgkaLmAlx37/C1PBm3khvN4b6AmnO430XHHUdefUozAEXqf90AZkSVssTuiHHvB0/U
Nnd75UzBVJTj/97uEFravOBu60/rB3gvQvV4xg1XKI6IMeyzyKTmreIkIQpFzWnIP7+rkgJCbfuV
jxzrM/QbBhbJlP0wyAYiD1VpO2X51bqEhf+SecmTkzWovBEVCE2YEKLswnftuuAefekI30iLrJ0K
ZRSaJT/oam2rBuCndQC1OVuAosI/KjKo2S68rwZhvHeyYHXQyersqfy43OjadUFtL6w1bVy8AHBu
e1ETe7eVnkSzXmNg7RjRUm3FLe24gtc+RHLg5pc3cq1Xrhqa3qDIb+UbFuznkzHt8VjOwFUrM773
79/KbsPmhm0q6IRn7GCgJ1AcH7M06z7OQu2MAwbfLm3cW2seCND4K2uJj6cDOXoL+xwAr9nm74ui
vueJSAIrwWeGaq+fIlGUt3TAd+XUImMR+HUBJTORHTghPw1lUgSvCYTYGaxS4VCRpUlk1Kb7bVEX
HAklbYtPC8A2eQBCnSGD6YUo7STXd4mf0lcHppI60TMF4AinBt9enAkOGsG/e4k+ldnqTTEg2m/I
8tpnN9TUd+E5NLXH6J5UlYUnpLbBZ0y4QN1eNvDC4YL5MN0D8hF8jl2NNHjyWor5vlYy827vOStm
oaYcl+yxO7zSw1HrSHEzW3LoCKCtD/PTIZtTbTvVXl/vZVwq+shwj8LDCiCloYueUJShlMACbunk
92P5b/hzDBFyJTTTNeJYptbNbWQj/zoT6dGQEAUbjfVjx8b6i49BtisrciuULDbE4w3BDztV7KLI
dAgiTZf0fxATljYuht9l6RTeE6/36BytnWO2MJcGEmt5/SdKsuTNdz/BzU3Lq1ZrboirXvE4gkwq
SompPaAKvEIYN1YxZb7UHBvh86Jww+5yfh9vqj/NQNXlRhv8k0gwzJj60Py2BGY2qq36PUtNWA8H
NPyX/CNi6Bi89C+x8V/v6Qy8xAXRMwrfJ0ZKlBdOHsdUTipf90iYzeMUYCCKb844u7clUQ0KMz2O
b/lorwMV70ZqftsT0o3wSBwAtSZ/077szh0X8oalH9u40hTJ//sU0Swyz+SH0xtlR71eKsig04ev
pduNI+NUS9+vOTKvPl2NJSsChCNDM3rvwCEMC/B5aGwVlrEqJ73bdfnMOq70OOFsj9NrQgj/epYj
HmCku3GQPF2ywAR7poa2fNZiMX2eM2XckUVR4qjEavz0JdG4w/vy26vfWoTN+1CcdD7a017PFsjU
fcwlWkXHyYov+/VQp8oaQXfSPLtt6Mr1209SBRDD96uOmIHwQfTsv0Wi4DustCoOjC+KiUOvkX+o
Gps8uXnu6aqRZeNPFI4LSkZbxM8gj95nmhxLkSzTIJ4rgf3mV8jsokL9MAGhlMrvW2eY9/edOp1P
zHP3dOrkkZx48Ja/krzdg2Qrsw9ZbkoihLJO3/Pnxjmw3BumKg5Au0vAnVGUnAKuOn+9uLkSpmrl
WzsshENJD1/fmK03fXVXvwa0dhqYfmjFpo5d4x5+FKluYajY6idLcJE2o1JgQzGINJpytM+RNHUY
dKt5qesA9/NZZPEb/6O56cKsJZNHrvz0qMSEpqsgqBkr8khPrKbtb2uQ+wxIyOOcCihmAB3dmZkz
FBForfCIjZGft+7FsXGE9ROVGchJjk6snbLU06cVTjToNII/XmHoVltCXk8dzCWcTTvBOC0DKwTO
pZv3i3+csaXxHu2F1S8wtswyqd7kt18rFiuhgxsDcNrs3tQZ/xmtydvd+lrvDuG4gNRZo83OpMx3
L3W5U2weQXTmSKkslB2V0NH4zfT1c51YQmpUoyjaHdxCMw0Vg5DTIDafSiGtkMzjQ+xjqkorCspO
dZzGWDYEznoFW6ARyv+JET0OUWzXr8uf9a99oDcUU5pRN30QSK4FptALDd7tRbeAqQs8uvBx8Fko
fLePQsIE1c5gm7TzHoz04+BByA+yJQ0osUL7zaXHkdvYubNRIQoM8rWu67k9k+ZelI8Si/9zPLEP
CNlsD4Bb5c/rzT9l3Jq6zkTTpvxiAEL8e3f/hTzuIVPGORC01+QnLXCY0gKsgK9neuj3Ad4ow5G8
xm6cUnh8JrBmUcJvAyCeKiBTQRo0joFdiAqoU/IWfpQO1uJHGqpHU+jvZHbc0swf5DpjdihmCElr
r92mdrGe9+sxHP9mjgJDTjjXDtB9DqttdGLaJ434ryNZroVuNsPK3YCMZGPwLGgpXDoo0FnkjeNU
lUO4r5inPUhRdPKROJlTXQXaXOUIcQiZDKmGbkkkUC4eKHiv7Q0Uky7U+18FMgWG2f4hKLlzieRr
/GY13Pul/xfzKbPdq2eB3C9YLAMhmDowslxIbskkAhhBIGMGUU2vqxDFYQwyb0vR6jnhXVQ7d9YU
j+wUv0I3WqYUc0OXNAQNFSRRfd3LcElAnCY1hj+qYEU+VuMNNKvn1Izx2ZZ1H+EDtwfw3M8hyhze
71wv8gbb/NxUsY0YBUtXSctTW3laBhf4TjNw4ZhUBebB6xaR2mh6Xk14THA9QZO41ZU8PNHzA571
YvmIHxylnow9FfpGh54Ci/kA5sGzNcEUYJDR2D1mNvoqLX/1kGmDMZHttVxio80sXbZP5aEXpX5V
EvhJ+QxgcxVSfoUA44ABv2SULS4IXhsA7lmNGbQhhyqlj5Ckm+weEJvuoEHEpvuRrze4HwXf+PQK
7oRSsjIH0qdTRDnvblkESwGf1fnuSreBXKol4uJT1OWI1t90RmgVA6qhCTrgybJpSiB1jwK0cGVr
+A0j7kMH6HWE0Eq+/pOpBKuqV6bYGgfk3UQhhfewjECFt8A2A06bQU2BdIzPJfc7PNeYO9d+7jbb
8XGhB1it4OXdBn0aEkl6wCssU0kGaKOVAtqDLpmZWzBuwaDhAU53By6yJv0xCLbOPk3bJy5wcXww
90VT7zjY5z1ek92A/7B1+bsI+ZixI7e2dCtvRM7i5/qY5+ot4zz3IsXPl5c2eaETEpo4K68lzb5r
MvhXEBBwfaSkhv5tT7Gj1N6+3nBXtFYYbkpEM/Fct+GzJrYmZSlhjkp+N7TWA9VH0tx/PwFrYU2b
N9fiexsWNv/U3f8DIqRipnRR6UGPN9mbQN621+sRMCFzaSv20osj76ts6rn3sXD7qY/pnqoXOjzG
t9PStbEJ8HkKVDuP5giWn+MgGRSm1r6cGoQAZwl6LZjbJRtvUr7daBnNh6stCoye9KicB9xkZ6U+
JpmnMxF2s4kzyXBltWjhkCexTH1+XL9Lk9iPaBXrW7Re/Bbn3FEH7yk9ksFUFdAh1MefshLNHInz
aBsApRobzRzRi59i9dPQw7JwiOIn+cXAHd8wcUdv05Xi70eaQYiK5NGEjThB8oTldfr3lr2fYYNL
FnLlG5RyDNRTWcBnHipAqKJPwIptg1Q4Wk9A6JxwzdlvEK5d/dTVgIu+KEO9wWgSd+jTEC/vS3F5
dhe4MpctJBEJfUYnn9OC/mA11zJ/nZLn5NQP+d88g1SYERTfqveNTf8d3OLu/iMgDq85fO0XOSXq
KE6tKcPwK7Olppt0bvHEpVeA91tSWFuRkFlQQBH43foGF1gA9uFLXloZTQEYBg/M2NPWcsqOfb0T
jTe+80lcUcSdub7degCrTT8PQ3bZ5geB7WiAq3kvKYX69o9GL4RcRCX0QL5vji45cFU53RWkeDtB
KcBi7Zl0oOgXF8iSplxcNi7+PKfl2mkz39dq+DxD8yt/6pJrUUwdQ2W8t6s6O4vjjtVaoTIOVdj1
GiUHyZ3OW8fpJOvNkvHh9faOpfph289/89ih8v5z2TrSkkLYHO6kxBWAZF7xeLgTr5D+5XknUHtr
UC/TRyaXLsuD/1RYk5byPiTTWMpb12DPNmCPcveOC+J1t2juZY34FFtULMJm3Lf+cFR6B1Lo8E73
Y1gr/c6hEp+7dc0SvmDYfyhaIRROUmyfNvDG9IgbD6pldHArqMhL3mlILXOcYPB/MdFBIJMV9XC6
tsR4oNvakp5g06H/rXZxUXKzCgy5dcsNwKHzI8Cz44ltfqmZ7d0IDTcqAgtUn225hqMspAwTeIst
ddqQofs5qRwT81op+KQChIbLPpBnRDYnD5ZGvtq2e3wXH6BrEFKex6gjT1aWRgwAc+a+UaaZMExV
/rI1XZSdYvl050ja1g0R+7WV8yPlKM4H4Bg71Z+hYRn8Nz5A2DPioFGizF7hgsJSSYJKNQDv2/KH
17FVrmx1UND0FPs+aASFFIGO5aKov57NXSINc+i4tTdxdYs5Ugu0vpucmJU60hBDxpQ4tlzwKBZR
Hgq7JHtpfXqLlBzFnKc+bvz/cpsjS3tOA9nHH/rpkzTlrJkISljTeZ79e4Wvt1G2MNLSkDxaRFq2
xRQO2mrcsO3RlxMD43U2Y66FlXSVBtGkHQuQm8Ef05xcAnfBYIW2G7ovsN5W8t9s3rkVnXyEok9S
uL9qOzYvIu9Ml0YkjFsdNYqLSNNElLIrUmCH9YcP2+ceUczwA3Q8a8p7Nm+GznjRwDFEuC/7dDMu
/0G7EgMKn5l6nU+5SpZvvBVM+qx9XKDnbD5F4wDCYoWdGjdOUGlRykIGqg6CRCWAgVpEyW+2kX3o
deapWehevjpzclq+FeA3SrybMvqbSHJgOk4m/9AsQr10U+dTT8rbWqVmpfX3Axnekd4D/rGLetDr
2T5IiDoVP7CjrjfpPgaEKgRGlu+hHdeyjSmPsE1KJTZ+AvhTisnel1yBUHm3rmu7IG4kgn897dHH
+3ikGyvHaGCpIneyB6Ov4+lQW0ETS8XAQJc3Qbe4rlHH66BdM1FMZw2mRM843rA1NG8JTvc7lEaQ
frRYkzSksHdK1xuZIi9+JOzvFN71cCpsiN86sg7XRcXp3RQRP/1aRbRrTg==
`pragma protect end_protected
