// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NwPCR/lwVC3WhDYa/dtuhOof6SZDBNTxAPw9i8rUayTvqxPSe4gP3a+vVKQmjacG
a6zb/zTdntZ9frRUuhVd31v1Pz3+MObZ1XmC7kb7rsAFY4JnVdRs1JlBFenJXtdm
blS6zGm2MN91aDmSdeEJAwCnzfhmBcVkzogInRNnK/g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9728)
tLP72XLEzmUV4J/40/4OUn+Lxor+Z0eoALsIdOVUss5SDyz6i6KoOe7W0+4jStmO
oznUOCPkz3V/IxU2GBUekTaKb9YHZeiheL5Aq+fr4BmCRO/xl3wCe1wbEiPlz41+
O98QBzdfRt1W0jSk+5xjaRr0F8ZcN4zs63ILnH2XeIsQHRSMml3uG4I3DsBqdeBM
e7ikPONr6uzxS5iJzzgbxG8bzQL9mvZPqisdJmG5O817KWiepK+l+Nis4A2Rvu54
8Rv4Uvb34BMCzsOANtpGCQHy5SHmJKnfVJBrwvW3j7lFEp/r3KKgrATQL6Hzeob3
+HmYZePyPMS8Z2yFrzyMNPTp2KrPHoZEk1pX3kXEIsSfLh0G2tDxThyEv+Dfk/QC
0qx7GBjYOMnro4yech2eMnfxnW076W6K34Av9xfSGEzF+nnGzSsmQft1nvvLmiZe
8q30MiARvx3aKCOW7RjCFoBMDGww8yLiV0YJWm7zWHkzd4uiz5j+Z9rK1DPRwSUU
mQvhPUadXDs4Azo7+//Ac8CqI4sLL83/HM6ubSOHSbiNqS6hy6vn7GgLamb3/Fpc
WSzp5C3QTLZ80wk7hC+SuGG2a+QSo+kmFwwD7N8x9vjeuc31XosVupUN3+obBXcY
IL6uo24vV6+NQK33vX4yCyjRQXvJr2LNg+341fUEVEC95JT+nEZs0fmRZxTLdiCO
1ula9Q4rEzmkKhrxUM2/T4KEQSPD3iNsPxKOTTV6AiGayobybZHt7GhvWPEALrIz
AQw+IIO7BmwElnpmnxVZfdPoqEUGL54j+q/Yjo0DHV4OfRkoS3q8ib2Dc7+kVeeG
d/Ec+/cpvWYUGoasJMcvhKjuNhKK4o4Tw9v8qRk6XkQluTlyNX09V+7SRrTjCg3V
yL0vh53wgRkm7MsRb9Xxl4bA0U9UzpjQs22CNAdBDjaaK71wpy37EiwaoenLnEia
3vK+SgavEfl+Pq7wnLBEck8lEnUmi2MUWf7gO7czuPNKE/yG4/iE3F3ci6KZtC/S
uwTpKMl+ZD7sg5FVug0wLD1hXONQ3quZFRuWZp4looqCC4ALQlOA5rTpoqEM3e1q
P1X+ZHtsSVif0Ww5wFhWh9ggvPnqbB+j7nB2nJB3fSicGbiKSpf9cvFgxUCftMnE
Vke1YEizHFAj94VOZLyakqEj6NFwVvYOJEIEwt4pcg2/ohgJJH+411rKZZP8g/V9
Eyxkh6AWm8kWZhBMNtx2jZo7BBzoXO3FiunkiqquV9XZClUD6xE14PRy7rZdKEWT
IzSm42v1txAgebT8tPeiN7JC1HafmYXkG+k+aZ+0u9tnGQRiKhzrGISrjGiEU6K3
TIZ0EmEVLiZzhXTq+Mgrm+TMvPyK+IRJ0jUiEjKQla2FCuR0Z4PVE0MXaIhG/sAc
fxAXKVuXGTCVSXSkJh8/UiuZaDkMEpwTZgrdKtJ+px8WZdeM+65IyGm4Kc/ZX7CU
vr1wFi26zOm5ukevCwjgJeOU9xUxyfJ7/6EUu2kClt0jyXP9+ITBrqmDV2/bQBv6
EeJpt0XcuWJ/2SOsgHAEIMMVV4FO5Mb913VldKaTWmL7LDeQ7pQ0Yrm+6D4TjL3y
hhGqq/7TLbqQjDWPWojBz3S17Wts0+RVGcy0OZgCTx8KD7FIO6Oey2CctkOa16Nq
FPG4hIK0RtJ6ci+4a4xl4DGDoLnotKtwHrjBLT38r/u1JeJLTG4nVi1j9e/Wg27E
jFKO8v/bbka9tnSWHej9V+j0H36a9dpFK7vzatKkzDAHY+ycyUa6lfP0zIN7D6N/
PiPUb91UsjPWseLzoh6wlsWeU7LnEymjMvbOMJ8+DRsyqhZVhbcTUQGr1/XxHvsC
QbZWMr/Y/pVClxcMThMfa8Ofpk/g5HG+Y/aCY6n4S3JFYPFn8/2UrKHCTqeKqsm/
evacGaZfJo5HL6EQMszUDe3wSioYIufg99RAeUnTpK+AT8z46dM9LWbEkq56wjJH
XM6VkIUOaILfUCWmD09+Yuy5IffEtObdOncjQkKX+WUzpJ4FT/hm41v8hSHlKU/Z
7paMGFHR0RKqkKPZaj2W+u+9gPXE491HYRr3kbN1t1uB1e/wYkoTI4VXott+0zTf
Si86MiEpsXOOVVuNpacMlVktWQXjb7UdA0l8fegNd73u13MoFm3Gd0rruEu4WFZz
6FoIeLt1s0Us8p/nx5w24p36n4dfuawKmJxm2pnUcQWqvMrNtWbZqHDDwKmsFDn3
j3WN3nI/E+CJZXnzz210lt8WkhHfXYFok7b0LHuWZC9bgokK62i0dcYVKXFa7PqJ
ejF/qIO/U8M8w6LNbTDl4ScaR8qgP2Eqy6RchnQNekeHTZoWFyLusQqskHfl/PgJ
yD/xpkbYYA+AWHdYEUFsIVBZ7VQOu62hUSbnkNF+LEg6qV0x61srmAHrvhWLnsrt
8twk7a2K8fHs2I2EQIje3Gm+KcOz/ljfvMnUuZyCFfJuWiBZYJqdRu8/Sm8sdoJ8
+YGBbTobOD4auBVl0IOuIgbDC0ZNxcHkm0wDFw7WGZQ/JRP+mRqKi9Mc6pUaR7cI
Ai2BwUcYMOS/5FcuSacgrzHUbsm9L5OXpXtt/b4A0wyafKKrQj5Vb7vNQudrmisy
xpcN9a9TNWdEPJMZ02sLJ2+4GYMqVtLqjhlvEJV3zdgs7+9AO3X1nM9+qkAyx8mU
0DYqvWNGAdqmpEp2e/JyBHBptArI11yc2cZPHFG/c4ChIZkxjy54motZLYmXYp5w
SPypJahvuzG2ifm9Twv5JFqoImuDyOp9rOGZDIllJuwmp5gr+MCWR91Xp/wIzCFJ
X52eHqulqZY98rnHCsRQJ4jNd8+GJ021eshqo5eV8jQHcPW1kLw8xOyY8irmP4ft
Ia4cbcH8hWQq54XuoacowMDBGsJnxvHp0ieGUtOEfmv1VI6ZuTsyIQ+D2CTUPmSw
u7Da4/+6mDckxwdKve1JXHYYgS+/PeByBIg2Z0gu+LprYNZ4LxPCPwlx1JrAHzkP
wD2+1oEmLX6t5BJL5qKoPR1hX40XeZ3NbhFD7EjxhIDB2oFnbm8HGGJW3gL20lel
cdWd1FEPr4oEILZoeALMJuCwWV00jc03A+haTXgJPb9yw/AQHS1edGXeu35NACXO
mlv8ZiUVrmCbSrbEUxjS17NfJmwRswgt7zG0IUkRbYdy7YxEEG0kAqC0NRVgWDcc
eCJjRSmG2Jie0e0MZSJ3P/DMGSNtLsJfgagfXou1j27vjOhJhxGCmzZXyGxXRpP/
lsGw7CuhlDuiZWqup7kdQ+Jw40R7OMhOg5rJ47hkQpLoD+YO0PMQmvNMhQtGT3Uz
4FECMyN964mZnD3oKorpM7d7CrESToUZBKWqkY2AjJzdlLH38NkW9rGQ5X8Oe5WR
DTf5Jt9my1Ql4MTnffqyLyYbJm3HrAv3VKzQEcbib5vhpQHuGK/LMb+NjzqAGnEJ
48A2lPq8G/eE09bbT8YDBtO8aYB8k5n0jsTjmKvA3cBnmkf2YcGRNOzKAgrXa98Y
4mIN4vfVSyCb819IUUa01pWSFMB0WR4Bb59rysxLB2vAIj/Eo/oh6tZFL1FnhoxS
5WKkKy5uQk7PHglMMo5WhjF4B0JIQlHZ3+oo7GVsxoqvUNi64qaBTYTya5iKkL4M
DJVIHx2vRb7XjzlzlriR17Gv3r+cLhuUssIgw5TpYrHBTXLilRfmnHXFtWXKN0un
ZuHkOqCo2I8mhFd1ZUKc5qYIs343jKvQhsG4ls0QhvavsX7A+NCGztEkmgzsO09f
XfH94eCD3fqntiHUb7Zpm7edLIsd3bYa+3yKnH+NeILY/Nfo/n2AJjC1Qv2uFm72
SG+ZNADERZ33op+kkvvY949FH9VIHn0EeFzYwP4lakj2Fy6R8gp10fjAg/4PyVs6
QlmY8PHW0nk/v2jyaOzpWW0q2cr1jwQ6Y3RqDvlgVOio6gO2AWXcQCcc4OpJOQSR
KIFhKZm3Fv8FPZaYp+FJQdNKeV5Q/hEVO+DvzK0eZ7CmBOHYewb001HLCGbXeK+r
j4wdCLLuziqQzAeK6rWGdJWwnX60XUucvEUQQxxlEH1lkhdrC4G9Z/ma3gP5Dx4l
jVW5VTeuTLbw5maRaa//Rd8W8d78s0iPgP4RED2bpgSkmh2oi2Z9N4a5/ZeHGFfa
i5UadzljqC1LKAhthiuAWpdPmkn3l375llhyxxJL/gRWM3y2YG6C84yh/PZG9WBr
sDCYpI2x/dj5ovQ1QeOf2IrTkEk7dRjBBI0ZE2QNSF8ZTHBrGd8Q4L/eevKyQGFw
WdbO+pISJk1VDjuSh/eH06TrWjRSmliv0ZY86W91x3KlGp1UlzU+ln4usX6XrzNZ
Tuy+Mv4Iy6z/npui9DWiJdsflvSA6FQz1I+f/LJFG91LPzUQtCtwU2mv3pDN/FEb
xzQonh2Nhdhcx6gBb16Um5IQTEwEwr9fxrpkFqNBDJwKjbOyJyPlOSKxYue+pVb1
/X7owbq4L3ptuYqmT9CwOeLdxrF73Z8b32yYwaAB4OyC74q4UB7AbR0MrYIJSR4b
E+H+GrhMmtN/upig9Pg9anYGsA02nNRWtwJSFhWnaAcNJPerWB1LAuNKgIWO8rgm
TIvr7ud76YAsZwDP+YC7ISRa5WjidY85nipYqN2wGroBizQUUXbjIdxEXsH+mokI
qtSqO1jCFHqhYkzgXBMImnIzB6q+1KbI4zlkEuT8u8/aCBq2s5IUkAuM6utMVw9s
tc2q/wRltS6GLywufBqe5iF8dEu91S6fsrlIZ9cwo7ZPaTH/WU608Yd1H4WpmD87
eFnP/VSG/OOGo6yKL36QpuR5g6QJ7TJSRmZEvJXMjyQRRi3RpZkMbd8+OEPLlBMU
f5U+HS88qd4YVY1vlPU5X9BrFvpiQkVis+SW7PlnYwa/lTdCrhtgGItkZa1evD6j
wSspsk1+ppHVYpJq6K0Hzk6Djx9Pa6fkN8yI/prT/tDwo4CpbuOcyvgB2LaSfXPQ
vW5XWk5xJj+fxpz3ph8FOWKqF0uViX9VDMTu0s03o9qF0UsOAzQBkiWR5huy70e6
DwGCRhcutAEcxcrD6QqJoih4yueX5s7GO9hZmw7THG2q+7BBjCLqC8K5AcHX+TwB
U4mRfWcJJnZa29qpVq8SBsYUQ3UTQupkAwlrkGjiT1xKUkvsHsRm+aEErtf3G5LK
yTQo64obt1UZFvMuDyrykfLCyPQEjVXHuxwfA2fuz7kP4asVOrqh4N/UFlyzmXIb
ja9cF+P+J33OInwMOhR9qTcNEmTJkS2Y/YQBoPiBSsByCuM0djvgnHhij6Nv0uEb
L/Xqj26A8RXeuAqSoUzcrEu88Qrk/6FWgcNpCJRe0Hu9FKcB4UEzt6k/7CY6c+Lq
hSmJ3YFZg46v/L8uVVA14US3juQrdlr8BDU3MKJJJnyaoO4GSt7UChXDIdLgfaiN
4mwlLrSMKgYvUnPee7/15mhj7p9QqBXR2Qjysd6xPr04pBvav0NJ7y/bx1IYdIbS
eAhZojARouIIuQ7fNOFDeXf9kn1/1dPv9dQuca5cT5D7VX3r9NDSDzuhYcVhZT/N
0yFEUm8VKZOQgOcdr7ds0bPH1zLBBcFQ+EWw1uP5V+fKsPpYFLMet69CI5Wi7apm
V3+hk2OgZMa/HUC7QRKYOcGz22u9V43oL7e0u+DbK5QPjfxER9hx4Zo6tq+q6dCA
RgyKLIfXG+utt62K8Rv4UA9HyMPZjkrR2yXXdT7ZuEJG9ZOrZ7YMHba8GwIoJHtk
zL0sbYshLoGf9nipU/jaJ7K3VMiwxsesNGytOsvsqsx1r8kKED5A3+cLmRO/qhvx
5/cko5lVN3+8puRAX+Yzzh+yUi4Y3fvcNWw2biXsUMfT4cEwAcjMpqb/fao7rqEh
xKvx+UX2xqujqBSsawLTP/GhHffpeKc8YK9jcfZ0Dqmc32xmwKRFy9cleZLtSFbD
TF2HtBoUS6hYzMWJ608fwn+Uw5VO3/0+5J5JzcfvK3Lt4u9t2VwZsdRaageog4/w
BxE+ubpCfKVPlAi/LUJP4Jemin6OUVrxsXmO9SeUPNnlrNUTacgMSdtIh2qoBouy
Khv1N/PQYY0Ii4GfMKUYgHXpTXonh+8VEzqyYPR+0XsPnTu35/K0gSHMpw8QZr4f
YsDyYl/cuBSHp37DSAMDfQ2s9TTwndi4N4TSgPI8hL5rz66lcfcBVdDdZVYa9Kfe
xAX9jXZjHQBqAQtDT8N8k+wu/+GmX9lIo/m5hMB/BYfUuBHWsTCioYlbwGhPhlrz
9ZN+zIL+L1yJtDqRccQhaEH86X8WacmjWyQVFHh5xywfKcXpK+g2y2s9mQ8MmAME
51XbKkwwL168kjueoEbTFcVwx4clOgmN4upuODX3AikM6VbsjDuo+EQAGH6k1/cP
jy6SMO/EYdcW27/8Rc/vX1UH4ulquZHrwI+FyhpykZC+8ZXP2rhIc0GPYYfgaNDr
KUX1+rRPZOC70PyhE0gFPbi7SgmYBT8JZ/ieqd1MO01k/E01gcOlEInKqj3wuqZv
Ub+js/47fiYNRl8ZQXkVeoRGjyf8tRPYqGpCkdbXDStaPaNS0Mop1umkavPSEwbJ
25+DIywRUOaewzPeDgQyNfIYsHZBlAs0uPFI5iAPSHgHsHChJYgulB5Hhib4DqMB
rgv9y+hFIP03wCJo/7cnT7c6/nuF0ku39eylfVE1Glg9zVULgwryN3K9xCwyt91G
thRa23njVrezAIejLkOSEDW7dsYdQuC7kmTdPvdzI5rit8E0r0NAHbImW60TPrz8
6hoPpqsRWPOuiz4cz06wQHjmP47AQ99Je2dor19Wadm210N9AvMht5tfyyEroGh9
vsTPlohdE25zviIkIdexdmxf/6BB7RCDS8oT7yJ4nv+sc53wQTgrFYRGmKKq41el
iiSmEJe1RYLW9d3jVrqZZwZEv0FdYKiRly76KNr8ZPV0JtCtfTInAZeCZuyNqTc0
Ac2Ii5JzA106KyPptJN1TZDTtOHp+/n/igtLcf55mK2KYNE4lqvc55atCRVMYheH
nNPlg1IXYfJM6AWbhpNLWjHs/hB44IfVzEpxMz9lkiW9S2SYBRi24xiFPPSESUHF
QyPm3GScOPWuiWOY2Baa8aJshnCo2IiKPmb2Nmncs2JyA8IabrCXyT7X+ZZvNSvW
4RnN9wNsGoaB10ZpN/LvBGKEd09AG4rlEpcUcZfLGmMEkBQkhExLePqU/O+78DK6
DUyRm7HlZcI9KR8tJZ2DFac5puSWtgMd58mOfqi9eJ0lOFaXmAuTU6wFECjUx0X4
bI8/QpsLCSM4/m4EBnRHCXWd2eMw5qpPwPXluZftZjpHahZl9GbhVhLbmks/1luA
YE/xo7lKFqMtnlxR/BO+V9ZMwGrUrGxUkVXkMZMGtc7fbacEp0fjk6DhJtH3skGP
ZtRuQj1OOc7X3anKV3BKOLk4AGnm5vr4E84YPBDj3aJqkzqQJZoEoJL46EgqtZ+J
Gl1WBoNLdr2nTDsrYxbbe6wVIDiQh2fC4QJ+5lWdjdA2qdm8DdRgZlL/CDIcOLN0
CloY1JdT0pitcfuVxoic85qWojCsYKaJUdJkVkdikPJCmrt3RQwvv9t756uhcYHA
skfoPLt3xs10Pq3AFtiQ4ePkibZXmg16gRR93Rj+t5p/azi1q2ag086XONZLqIjo
BR/eR1l5zVpW3Wya9IjG1Bke5xoYbwvHlOvPILTh3UIiDHvvPhUhCvLmJLiDDqkP
HfRv2VX8GaFctVsEr/5Q/wMVIdEps1xSGurvvdwzsu2d4D6zbqGvHAzCFnltRhQq
/KkW8UcpmIIMwLH3LWkOb+XRpDepTmrkzB5/BadX3hMtKs+1vq7nAifD/3a+wEcK
VGjoGkyC9BvEpu10hMjWYl23ZVjrVVFbo9O6SmsDN+xC+QFZt463DeRuRzev+XjJ
WVNsveYWj968GVj4AR4p+DN5WozHbn4B5Ru0D86E29Mvoi3sdpKPnil3+VJVw8gE
1p7Je0IjFTEcZ/K+Y/Q7OBKVb0Wmx6uZuNJ8xV+dPbhusTR2vakGYjLH+OIzQEo8
PdekSvGMLlW4tGfRA5cAL8jlzwBvMa6jXinwovPboP4cLoJOKNBg5Q9iu1qkaIL3
nOO6xgMdAe5w4xNCZvypQ7SO/vgaQ6dlAQnA0OAiUoDFf5GDEKl/YBjZh10R5ljY
wdLua14pLl27aYEz0MIlTcJGboAqmvkfElWEM9ipTptBLIdS8DmTOLj78VDBCT/P
7gW3+t34oqBczm8T+rjdPqlvxSsReh73KU9pICsWGLKJm0clo4NOHI6KnveN0Mtp
/Wsei3DKUbRn/FYDHCJR9bwyusFWRgarCqdokBQuTXTTKz6WT4yhex25GYZItQxQ
Z1mzZfb/naPyVL/ex4KQiIQp3qUeiHWEMhLJHWP/qo90PSdGDUJiaFz4qOxlvsUO
RW8CALlUffTY3NvLRhtRkitgxSWPuS5ztZIO20Gn1yuXzLnKR/BgfOPNg7+OaW1g
v5nJxHEtGGSsLpwNkdQn15l+t5ZbpA7ag6atndSXB5Ieq5davIVYpsKODMGk4sQZ
JNjXRti5960BcNfzOJvAYCZInEb8B9vC2IWbt7TTLGA3bFouoBJ1/SYVQx1AewQ2
bwBVUpa2+ExYGr53hFfPNNW5mIufgTLNp5BTI0uEeSgYYJPi7Kf7HyfGfGjYdk0n
Vo4ZKU1slgy4/oP8kMPLM9veU4npUP1dPwwYT2nsYL4FZnuwfLlGQORW4qbh+z++
ARaJLhgFT0j673cXODErJTvmRf/AZ4YLsDM9I0NdzD5Pz0W+lX6DRoYrVF2czNkT
KyKKIh2VlbXs5yMnDm8LE2NADRZSd6ix4jCH1WaCJ5nWd/lFV6g+Q+jbeVfMmVhK
STivesczaWtkZ1iI/CDOOONjq8UMWzc+SA8d00vJeLNruI0fvPb1+mOjbeijnTIH
dBfHg7gZYRsHWgDTd8hvpqP+0OZll2dpnB7wo+Kv50Y1nVKvbqIjiRU6FEPTfT/M
K+lVqwkMdqs6Oe7Hpn4whhcEKeS2StF82SvElbs5KUowUqzO9fxXbG4GEKdRmxez
RLDM4RHRkoOAw96xVRB6ZzzZB0jNM1A0qgJQGqm15TAzF/TJTM+P8kAAw3AjXP/M
56N+lnzSwQfa10uAe2XtKVq1gWI+xmPLdoI/X/EnMsok222ryoGp2V/hN6wuxwJ5
jQQVxKTZwMGqem+J0Qk0/2EO41yqWMThCODcKHV1joviRuUZdR+ffH2r5SK72qHP
bas4pg/PIJfq38cZvpVjMokaKcpx4Eo5oYzJRWyVOzqMIrThIozayVg2yfrbPHsi
St6CPEesAwv2jvtbtT0l8RQRRhkwXUInalIqLlj9xjopTybHqDgCTRkBCu8ECmVQ
djXU3hWUANFmzfOOi8kAmeyTERQnE4Eof94aCJJZJ780bAuIWQIDts6sqdhXHLVJ
1/byb9a7FRh2z1qPBy07iCwn3PITw/sOD1qv1P6QOvcoNFB1boNDu8Y80umYethz
aQo/rSvBZ00xNvvnr/JxVpJHTE0j02jV8r16oZ5CycjtftGXvy2swJcKCzO1cL87
rfVufrBszxT1NzmpR1wR+/OSnR4yUMRynC7S/YMSaZN/dUrEexMEjWVkRmPfhRWE
hTH97Qc//HhUbTTcgsH+ighJyR+0N2K69OEhjjKV6hUp4rULOIVuTqwQwcOBBITb
i9SEuRMoJPum6iP/Emx9dh83TxGD7g2IJwmDa4nT1SA4Zj+FcwO6b0PgLC0CnS6L
NDgcSQttw6fn+RDBcQ+ppHGlu9/Ye6gECWgUqVOui2cf8JiAuB3LmWZGZN3vsdRT
uK/ZwEMG7Q7LeBAIYk3nwS5UVSUuK5aK8LeVpzErgQbPferLmwC7OegyCSa+KUep
EoKXgWg5wxCz5mNXLlYj2SFyCRLAG4Nf20eQTl2/xMLeQwafKwiWwp/57W4r44xZ
konld8O4N71sPl6bgLViqJBSgupW59Md8ezLIQ8scx6B4mPNBHFq13vn3vxv8C+/
WPmCnmhxvzJag/ZoCXGZCuG/cnjHnh7TYNRX9xGipuDq31DcIoJZ0BdHm/o/L3Kx
oazPu42UNAjxUojuySR02tNf6lMmBgKtAwBHxsmaBONwiLoys282WaX66u1j54EP
rIxBf6eyEkd2f6saSazUrF08CVMS5jlM3f88wIx62I8YkzoVYEtHQzl9ihmuGBkj
wdv8dPtEdfSK9QXYrg1lk2U/fYl39bEktsoDkuJf8R7NR669T6KhqQq1SuIaXtIv
vtxXSakseCuBQrjaMWKv7uFTHd6c31QixwBKIqHGjBgDo4E5Qu6n1gKHjvJxw1b2
YmAGM7pfSAfzOCmzasoeWVGNzsjw4HDl9APxoDz5gtx26JgGUQ45Wm3uaP9/p2Rb
EkSJoEr/LdWPlKMiwiKWWap/ulqiL+kt38xav6xGncoBDSsW1VHm9FOMO97uL3/V
lhLNpu4POzCmHCbMHBRLnJiOKEEv+ssxaJtMxZz57DCRNeSV4tNSRv4QfmWLgMnR
CtkS19ca4bcd9NW3UxCVqPSBt/62XCyVmyBdt8hWO6wkA1H1VGHtf4sRT0MForjf
g1Uv6V0xgYV3Fbf62i0TM6vT1OBJloKUYYKMuWY/ewCtC/iHwXweahxigZzOqGQk
KIYkA638DyVIgofe0U2vaB0OpH57lZ4knSYbTVRKsqe1l/XwkI1u2bBNaZYCE6Wd
rz9HhAZ680bb25NJ3+iz3glXNkjN0T2OeTf0OLDYhfhZDCbHdUEUnqWCZ6L26OQR
XJ9ge3aaGGitH17HuYC+7JZsOPEQIXoBRK7nQjDKGZfRCQrKegHqcrxzfyjNLfHl
DXEHTw2AJ6BDJWkXQOxbRpzI2v/nnYh1YNujGS5ZSGu8mDkLSleIYiA2Bi+wCPei
IHLMM40vMQIasSZpShZH+6BBV0V+OSBZuySjUqPACuEnv2D2bezczTBYBvNOd+eR
y1AVVEZs4juME8VNkKLQEmJngAfdwlD70e0K7H0R05IJyq/51cG5EyRn9KXl2v2M
QPE4vKsBRtbndE2P7CZ+0KZ9gApNwRRWCRkU9vrZvbHBQE3Q9d9EWXekOw4N458S
Y8MMwSzr4jKObu5QoiOjrI+EqCJ2LygJ9V4PNxO1kkdaJzQtfccr/eOBvlAyYB4H
RVKlbMHhufhELkIdLvIMevIp7Ml97ptuiB2Vh3jUcSGpO4ILOkKnpj51xQ9RxgbB
wTXqocSe5aIxf+wTLBb8SoW9x5bzVEkF7i9ygNU8K3n/H8hweV9le0rQpRBOzP9P
76W7DH5a7lSEv1uD8gFrG9X9nYRUaKMMXBhWiek664WKkAliWIS/t44fBG5GxWwR
uyHTbJS3KxitWPVpB9rSLO7jzZa6M3G/xdGm2G+zrobhipfznNI6Fz0mJkmJpFK+
HIdBeznqemDvU7zoYfH20riPhwKhuIQpHjbFB1Eta3V/PAJfqnCA+6sfXPVzsPMA
7kBKYQe8eL/gFzvvRdxzNmhA5EXgU7zDM+OLkpQ25FfNF45DInfJ7aMOQloFV3UK
7rAsJ6BaznNogRciX1t0zsfbMhLH76DUZ32lfVcrb3QSHv1ucI71EmgBWf9RV8A8
JwtOjjAORigopre0/BJ9jztvph01KLG0FxFgeBvBmTjPtIXWuEtLP4d0iLpBS9rt
5p21SOsuJ4Kljtlct44ZTkgD1xsmIUyWMk8Uqb1MQHs1w/YfgaMxz4a7b7wk+r1S
O0ZQWoEuoCgc+Mu7z734ReOLRnStyPDDnhWfGMbucl/4WytUN8YOpYHySjtKR8/w
g4ikL61sM3tqO7rw0i359YFCpyZSFlJ3Tq0o5MmcBu6RXSPJMp3qx3aP164YFVRd
OfBar9VFDt0jr+x+TdJ8T5SpXN9h3j8VklqYP/D0tUbTs8AK3QMjkcIR8Qp98BCH
tnXf2qVdi7Pl3WBtGqu/y32dSYbJOXJHrQRQ4+6U/lvjqoU3bpIGH07k96+m2gyc
0b1xb9zFPaTPq0JYzWlkXWbwemzewR7Q83U5sUkJVzuiriXaclYbpV5BHb8o/Ooa
Gw249ytGRtic8kdw4azHnWQ7dZSaZLw+jtY//yeSGlc0s5MFny0TY5n0QpPIWqfY
hjeU1DrXQePLroTcUmYvSzknyHmL9+nWszjNFsBSh5PDIW09B8KC70iRBYlsxnun
e+HkgLFCgaBqH4ePOzOL6a2VoRaAbY7CfyPVfMyKJQhISFp1Ju8VjnvBUCRlN7nI
Od839JGcslZmd3rYZW7I62PClskZDC4jTwZfcp0pH75D8YGwAAdOSFbjQoCPoOsG
qQUPrXaKzPkSRCmk9FWgLcO3oqFVdZRKC3hTQCdRVH/kLO/6dsgHK4B3jYHrUWm9
436PQjDgJ3KCLkg/luIBKxLfByc5mxCWrMz0utdwefusFFkcPTdYLVAFIjcAYnml
CiUzS5z8Eh4RKkFz6ZLQu2ayo+ymJiLAHI7HbUwkmKt23GiExB7lPX+GC2jn+nEs
7wu470suh2QJzg9sZ/x7sYrTuT/a2N0lIVDTTSStNIEtOC1GsYTWjo1jc0f2m5m3
fl3SR4b54hoQfJCUgO3RBVK2arfZ2jGp3mukBHMVROX4PrWvBVqMb+Uvv4OQKld9
Gro7PJuelReZ/zAJ8b3QGuZ6Mhdv+1dkbtwKG5byox/UIIHCOAkRjt3BrvLjyMxx
YaflSLpdkDsKRnT4AvlfSHBWup5daBh+B78LR3SjaoTqt2P4cgEJAr7QCyCt6arR
RGW3/nw6LywTJQoQLn0L46RwnySi7MjbdkomIci1DPrmHrVZ2PkutjZFVpY0klkh
KCUS2iqcuz4IrJW/TKYPEloawnJH74MuJHaRwzTJVuLJwG9Ttf58yjgVX+7d91Ov
ZjAsrYpl6OSaD1zzsDYa9jWfWuHz/WJEqnHL1XjO+UE=
`pragma protect end_protected
