// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SnR07ZpMTJq/Ssj1HBvLemCpn37ewGd5o4iHdn/VZlLJVF/DKZ+WbDkeFjy/ioat
nv/2Ytc7JCx183ZLEy0Q1DZUwuEJ3xWGOEartKEu6Kn6o7kTM0nNpQnTDvAN40cw
ffApFlExQw1Lm56lXAJs8pqEuH4HbnOmaHBrBQ0iZ24=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16256)
P8SMjeTCh9RzT6NXjI+rpIH/2RLKZtNnCg11ukgSDPj884j9iusQKsVyBIEUOh41
NY1SxU2TMB6/+RtRAwFsx+mubJfLPDUZVuQxggk7/g2Xr6w0eUVBBmMfr5U51jSR
1xFs+ycGU1KKbSba2sifTGyRcJSeSfo//GgcA8rEV1av+rweuA3FYkOZfvPXnBsm
JAmkWGlZssOSjpyOA7VrlNPhO6my4a32znBp4xXs6ULq+oqGrPyjIuWBnCxA/Hpi
sIaGc3KT5IkXIwNr4uMsFYa6ukQBpeAckKDqEC5Y3jT22n5FtM2gvaK4fGGobGrb
Nnnv3rsrOq1N7kSXgQmmOL7SFbnJ4IEo+KU42Z16i6qAIU9cIsWppsbqXFhZExHw
eF2rWlJDtnhq3gfy4xhaqWkz2TEa/NQcLFi7HR5KaA75TE47leYDETsAQgOqGkMs
Hoa5jKnu2njYDtC3Cqz8sh382JV3aUelPmCo1WrT0gTB01sOk7bAtv3y2+nZFH7/
80/vXQ07wgH2xbTzstMFmh3mR/gDMvxC3IYD2epWISdm4KrOWX/+LveOv3vSvobc
80TrK3tIYj3US2fq7VS94bf7d3KjbTbirF8xMpIQQc4FgG11KcoDp6sknLegpZbi
XgGFAslUdYsyl/kNtq+PK956XaB1fEgvcXAS2rTDT9i0eymga49NVo7Sy0h82vus
7814os5ncLcsHw/WXeODQpu5HOUEL/FoYdb1EW3UVb35v/WMJA1053GCthkJHGlX
GiPhIS6145PXxm/xnJ2OdYXdYd4fSBn4Z15JWGoGWUUIQWrSIaRvR1llgCCjU/GS
2PgiP29vmdDIVScNZpRDz2XCXw1n5Ek/ukRRDBj6v1WCsxsXxFsg/leK5X5oyWwS
cMUnV+dDKZuJpp7/bAFY+zXx/SEUXmsIXt3vJ3N741sJgfwVQiZ8WOZ99eQhHriK
wlrLB4GKsIZI+BYOtYK8Qe07BWYALZAFMGxD1x0kak1j8rGEvbdgokcPzvMxmYMg
NfKnrIjP3AtUi6DOdDb64ChHuD67VnNYQho/9sYjnZC8EYq2RVMZjb+xFeVNSrIK
8MKWLacEkw5XzGo98RTD1yioqMo20AhgQIFTraDANZMaaDZJy1pBAza33mq8Kuqw
evPDq+/hLQ2Z8Uqa3wYCdyiq3YuOv1n4uG8xA3nlALMlYvYQcVv+vljHjqNms6cw
zJ8aG1kH2+QLYLQtfnDeQ8GjdaAc481jocIKxq/oXP3UVuLaX1w3cz4o221X0Mmh
27sPLhFYzJxUc8pXWF0FxZGt3N9wCj+cFsQrqNBpfh4vfM/qprE2svpo53U6FQc/
yV/sNvScFHODeI9QdL+IsRkTctbWMzkslEwdXu3Ai0ftcnldW144ishuAX+hoOK5
w4ICRyU6el8t1FSErDCdbP7pXpgM3+UfuW0xEEXiPD128ilAsWQCl8TwbQ9wGj9w
9y/8qN9t6w9g7HSWgZepN97sPGznMHM7xbkwTwbCF6egvLsCkzjdjEw/qfv5qLLg
/coK8eNY7rHGHCfKi8ERNiWZVyBCBFzMsAxC4bs3nwgrvtI87YQ5bSiqffouomgT
2eDvaIfukKSxSQz3apCF6EZnTPMEiiFMMrZk+ISNV97jIoHJqBrR7KnK8Vcp7CNq
DvJzZFJG+e4QIOcbMunSsKSChqwqpEmIZM+hQOO8Cwj1OQo2cE0yfR0++Hs8Q7N3
pUxhfqhBiAsRWD04CIlobHvaZ2YVWw4w92wK26EVbgewxl/FpIgiP1igm0DjzPYN
6R6l6Ie1Sq+KGgn0koB0NejV6rARU+qwwsk9LI1vcAcQgT2otN/mhLUcSjdg4Yrq
dPC/cA0vjOe1CoooYHbpQ0HPbdBjSdIz+SCiQt7LnepUh8wq+G9opsGBfW+lzXwr
iPFiZcK6+lnmSn4hOq3fF4mNxKV08pzKIcL7b6EZEHX88wtq5VoQYFCRuujV/5xG
BIjkFSgRxOj7Ja/mFBHErAeZUIL6O/TNDZnTMgmJ8EqUQOskbpRKiOEk1jCnVrdM
YifCQgNW/wlNS6qq6+LJMJo2JdIhWZUcdkKi6+8yUjw7lKdHsjcI17AP6UaWUGZt
g/ZT4W9tH5C3TNoh1M95jOUiLQonMtlZVbJj7QVPDAZins9grolZoxFx/btLaMUg
coVZQj04sV7imPyl9G8WM+X4FxT4IH4zKqsiNp4KLqbycK/rlB+REo+z7V8C7Sp0
WsaKBQgA8tHGIqQXJesfUrelDOCA+DyNAQgMKIvVN3f08DzoED+QBigcDoMN7Af7
2btYLbUlldUpGWNGptJJGfyhxQe/VsqSHYXYoOpCcXlHhS7FoXD9Pah+YKWqIYJj
gBPPRn5wFAuZDpGYQ9k3SWbJ2NFURGSQge05Ym3WlgLWHI2k3KrHwRMR3EXhc4M4
hcsPS7rNxZbIl5oyt5p6d7CkrJi+RFS3WeDvL2GXcJ/ts+0xi0tSEcOwyA7n8gjP
2YsBBYY+M6Nw7IOq10FmiCsU+K8NW6WAp1nGLQHVRF3u5xUbI2KvIH4dSXu2ca+6
comqLehBPC41IdhM8qdRZjmDzRtui5Z0A+hMN/TByykXsO0g5YlvKcbmzjlck98k
IbHQiiVcHrWnCVsGBLe/hBOthTvrPz96JyHzyT30qqHa4uacLPveCW68OoHmuvQy
5pTL0FgWRgxHIX9zjKFa10Wvuoc9hJFsaJaUp33JlPuFpQwisMmutDbbpeVW+ixo
DlL2SyG1BBPYZs151wmIQ2obJp0d1FZT5PQ9ZkGRqCjMFauTQF9YywtzfvMUwhnR
3pDf5s7iTHm3PznHkV2ksAszO/ZADNArwenj8Cxc5cebDMa5K5X/WYQ8bQSi3IKg
KFLwP2H6eJvDzvXDL+ajdfUvorexcGWfeJW/qfGicv7fJOrpo6omrT1pPpr8hU3K
qqifJo56mcRMVlkppEBeij0omj69/q764qTdAjDFEqbpZLqAuAJVfZgQg3ui8FcL
VqxagWLEi/YK1J9+DcM+bhNuR1PA8GAz0neL9cKK6OBNoZLmxjBQRi9dL9cqPaVa
w0TVTU1NR4/CR19cfrukkbkvBVmk/KMetbaL1GYP/xz2wk74E3JbM5ZNxm9EsPLF
fBHicNZBuZ/SNIsK9iBKQj1bpCOr1aA0VJikScWpXOw7kY7XLanIwbBFBETPKN9Q
7BD+2PkdBsKkbqxawgRwKirwMSB6xQlWqvOCwDn9yEYEDGEXQfh2n1iQOAOPgvVN
y3v7OoPsRQxANVmUxlfMjD5qjCL+G7qEpw2/hvgZTB7HkwoYhd7hrOw8LypwXieo
3sw4TAdj5i0PBpOPztzs/KhmsTzOE3RL6L4vhatShEd1fhGXOuEcwmvn/VxtBqBf
RHxoeQSp45n4its8/4jDaN6o0Ua+fkhsYOsu8Q0qBU6z+1cE/Lc3QCIa7d8GQzRB
SY0j2mGoxH6ShOjwSswhBIuEs1BUc9mDfrh8QTS1e7/x1h8610kPWIgn1BLVN49T
q2ZLEpr4iFkoz8l3UVnmyeD1QYy2ZsrxSfagh4+VaKp9DuqimNqHBTEehrNX1RUG
SA4MChqTNQ92eqIa22Z4IYSy9TIHaN857jcm7SmReR+4LjhLw5u//FmHyBZ2x1Da
L82u7qENDQR5TOxgfm2j3B1O25P3cHenfj78rSWBhYhU+WQBIuAHU0DPap+AMyBV
e7NWdk/g1QVOfEKl1AtEMCpQEU6x+qMl6hOQSpO6NsZOQ8ZiUh/tHKKYi3jBzLYn
4BrCWGQKtFGIrl0YLX7P639mSMWFGCAFW9ktLOIvkhUxKrVX3IogVG+rATdUSIjM
BA6qexgj58ABzUpKNWoFAWkgjwiD7WbeHJfbZSBxdL7tnU6br/Ju9jfzmtM3u7cJ
qHUWOz3Zkqsuy3HOibG26Z/rBY6Ux2eMGMFNLpOq8H+RUi+BG33hIZnxjXX1a6Qy
Ff+Xygk23oxlb11gJUevOjAgeIwzBb/avkJWZQx+DhP6jPwCJWT7ygSpVeFQ4njd
rqnqtwTy4lLOdL/QGtLr4e6TupaxB5gecYf1X2xXSTX1TXfp3rQlW7Pawq/fc8/5
sCpgRRqpzZxeIf1pKWX+iX7SpGEWb5/XFNimQ4cM1KA9W6f/WMwe+dCEwrtB4NU9
QQkFiqCGenr7eHYa27J75Cqg2bsxpjjArdOKGWWK9HqDkvrrZegP5ffkBTFQFaj+
bnJFlkp9JsLvEU7BpQFwfbZ/wqJpPO2gQUS+4TzUtdx0rcx6eMf1ITm+bxzBMUNd
DOZ4/7RTgEutFDF9GbLzQGOOwLFH5T2EoG+eyNlR7I4Kx1kjAva2s2JGrdpRj89Q
wvU26jppkijl9VB3BucxzhJVgz5otO38x9aPmVjLJ0KOzDdZMhALY84Ctl23eYut
OD1LpRpnO9s1X/4PddBmJCJY4EDJeKXzl70dO3cmJi/A6S4w0bHdvoDzHxP72irJ
l/pyHFg/qnEL4m4Odw0zsfuCkzpYQq9u+ANEB3tfM2ybF/rJakBI7QNjxkM8y8X2
i8VsX+1Q2s5jKD+5Ss/MmLfrHxt2j6oyeF3705EMnstDDZE8GNaC5MXC2R9ApEoc
zAb5hFoABCOglQc14R7tKv0Bn9Rqi7qnVF7P1JIoI68jZmiOc+jrHbfnf/tAhKMC
MdxDU+kaF1XIyukknWCU2nAzxHVckQBzryTQXUdnshYI4gxV1vZts6AMIp9cOmUM
B4o4hH8ZygF3l7CTVSQ2BT+3HHNgkuwYhjRg5VkiqJNffs5zikpHLZuZiSr5LarR
RFGbWK8o0iaX74KmzNSqLA2mmlG7jvPn0zL92zcACZennp6AeTsv7gHJCPFcIxUB
F4tI3O8AEn+ev5dgJBAuMZrL6GJEnGi+5ycxP7b3bthhu5Bn0kGMHhYlf2uszmI6
qI5J/hjguvwgsSv8C6RAGyxhdbnGT3dP1LPoT0DgsFhRCdnEn2gNLjReaNpGzern
ekM2y5Q81XTxwQ4LDIdmbQ4KTfHP9R1naRnykmeNytVkkWQxKT8Jvgt2ay2OzAr4
YMlgSwC7g2o5XflPS1EvIsBnFByx8528b+iEqEaulJQjH+BiNPOStJaX7A5LiD4U
9zuPxDYoMTxqGqCDD5OWKYWHV3Vln9//J5jQAJZQbutwkpqQmDoubP+/KOslFHYE
GNv0RxEbmnOc0Bnw7A+7hVsFIoGt8iWEfcnnVWp4NkZdHdQZobrTQYYxhJZKrc3f
YXAzcw7YGfJ6NR42KtqvhXbtWVcqIgizgs52V/zwqCEOLJrhY17YfkgY534tgHNB
MyQrdPpXIesXnotgYRHmHyeN/Wkba7tRHiTuj3q9o8xz0qKIVYkexFeGycGfr3U/
QRgAkFb1rUrI74hAc3mIW8kqAW+mjlwUonqNl86lPqZ8GE7z5zClNFu2Hw3rLKs/
Qjyg3MeLdQB9TWo6SNe/ws4vKycfi1lECdjFgvnHnU+SZqTw5ytM+YZa/gZ6EanR
/3U+Y+O8GgKKVYH3kne25M/BAtdTUutUl6e7flO5SOkk60PrtFTzyzyg0bw0fRUO
D5DO7Uzm7qxUjbdMfxP/cKXZhNiiBGXkqeXf9Ub7Frpxf9nyQFxmvcgIotXS2zzr
+JjV8W8CDG3Ye2XGe3UrAtDOwbEp86zm44LDpe2L0UEIB+aC7jLV3lJz9z7E3WSa
/SylDd/6hwXMe/9VR9MY9dKqeAg4zLAnfsJd+YC+66Ecr9myMPxQdqFfvV366z8c
jyXe+qcaChddXudpOY05axspD6EYQ25S7hLg85skd0aEm0BhJhqIgdcAs3FTMddf
Agqb7ehEac31y3yPRvMFtH3Jy6Ee9FnZaJyGNNx7aBwUgd2DzY6TIUaVRkdtNtwO
1hFB+sTqfih9mYLSBf5ID0L2WKf4cYedtTN+b99P2yw4QSQY8YCJ0Rweu/JrKV8L
TFZPX0JeRJiz/7dScjCVwj7eZHKQayEhQ8LsgLHLL5VH289hnG+Z4+B+cK2LXztZ
c+yk3W3XW+oYBEXWUnSQVI+5JJ+tlRZqFsHlIlSHbQmr1Yg7lGIZq+xpugPVqDqQ
LhRXNM4+hO4ZLGCu9Qz9ZHMj3+8NM/rA9kAB4Y7sKWo67P+lW8Mx3Ic+DejkBDGf
k6jLBjxQ4iflDz9u5Ff+fOo8LZf/pe233lj6igJzUiosSH0h2bz76AKN6sYL6+4A
KJ6FUlGJOuM2BaBg56Gx66Zk7ZWSjatP7WzpN3dmfVD09ywIqSebCZLv9ai4GMmg
2L0Gmnexvf58SJEdQQYOx/41biyDI0eDIN2lep7LyeWj7sJQbeuXDSw22rOf0Q3B
Kh2DaISgTqX2Ha/rVAq9OtUQ5ubYOt9gp1Je0hSb57t25g/tjbFt6Xhh0+Ivnjma
F4VkTQlxoU4j908QxA7eMMknEsYoYRsYrc5ahvs4qL5EbNv5GDn4eUJCKWR/khVs
Q0+oLh/1dYm0BtHQFH7HVB8xBzmnGaPR3CIlRnYBePPIO83rVAVmE98ch/2tyh6z
aApsSwUFJnjBSKDxTGokuJb+sNtbn/reAjYLLTdFLHYb160LcuN7Soc6lcpGD9LU
tEHBJq1CYvZCiBwZNoXhDQBMrZCO6IpXqt0hcnlmuHZNGl0/VfysFNMUr+8wQIuq
uXke1q3ahGttnkH2I4TDloJWN8IsRJwldN980fYWo8pplqIKqCiaPthGKwJsyyly
LZNdmRPmUe434i3kxx4Ymf2DeiQTc5IcE/ZWJeD8E/4oGB8PC36YEHrYpKsidKJ6
J+JhQh8x6hdBFXGm/E0DO3ByD2MAUXyVjDR35CxKvahqbLbR2iB+IGtv7xUp7lnH
jREDPT+dIQctB43YPGS0oijG1owZpLqDilSNLd3WOrmn4Uxbf1ZDtlYkk+JNWvFv
j9Z8I6NCm8oDY3wZq6Yc4KsnCSf6ZavBCQpnedQrsNZEXuSYvi8LKsJM9py/7Q7A
NlPj7uEW9Jfdqy+T4/V4ivjwL8qHgcDv7JRu6DskYNi/eCzhVlqyvfUP7g46NUJ6
I9MN1sqr1ZpBnlBwLq3XiC8zR7H2narlc7wNLPKw0Ys18B6Olw4sYvIaPI6msDH3
e75blZJj+96xFvgOZnVlapvbJThmU4a6ERYui+bUsK61iAKYkAbunMuJUkqcZOGc
qCq2c74geZzZ8Ot9T/6klqNwI/QlgEhy1Po4ZEbPr/7EINl6AOSEwk1rJJFvO+Ss
3a1Pz6uBhwOX09E/Ll1Y23nvIQttqtHKfzMf0w9C3EaYgRopwcIxIyn87NRcZDCJ
NkXR6cDHTHRtZF0+DIiD47TO+hAkxpwj6dRh2B0SImTbEGihwojOMxS5K+zSUNm8
C2z/wBTvKqonENciQ/IIqjqESImjckm2eXUy95tZVzWGCYQXR2mTQCUvXKBmDMgs
5KOi4V+mgxdD81dGnHJkRSxUGM1/OwUvgNMiRSH78Z8pp2CQz6WzC6JOAL14s2Gt
UJ5R57hOjIWb3InJ8CHzmaltsrVfeQUVLlEKpnaGVF24OFjWvQ7o263rHuhpn8xh
svewM+koh1kNxjx7ZYfQH96i3oVFsMTYkDLoO9ApYMXbJfOpaaq3ti+CpWENh+5A
veUlz7CKRmuZp4GjTunnmqTG6RySneWVB/VOKawelQaoUYZJApCHKcPrvwqvwqJ7
ZAyq7xv45hsaLrwKjwO+PXkCTb/6v2Z1y+5XwK9yPrsr96JbX1BkCW5tTtCA+9bj
oA1WNQGxiYycvnzZRh6Pg/MhyooDPjIgIsUxQJuKTKPfdEj3n2FqmSDvyNAyr17M
q+EAdHg6V6YzDugOOHk7YwRs7feGZKpF0k1Re3dlLg3ixl3kbFjMghQm//cQlQuQ
76eD4SYplt3E+7Hr/SX+NBiGKum6w0N9qLeU2dgNUe5DM+ByARpxBtCApVw77fyd
p2sqDrw9L7JgCzz9R+TeHYS+H+xZzU0i9UXgTwzM/Nmb0puBnzWRhQp5g9l8Y5id
bEqM3c1w9y6nwhJYUIWSLHw5FBHh56wBeLzeGhiheIagiwiKds7vvSFxlc5v2d+X
lVEckM8H6fv0m1+yj4lie06pioFRjN+6/4s2fsIV7Bmt/M3nKuPRulSlcY+ha4hn
QUukkViKit1Gwl9cVk2+A+FjjK2VnemfIMHXA/b+LGYkY2EL4qOs6h+zmk/qTva+
rj0V546zVXEInF697ewQ6/cvZwZEwJv8UMZvV+lzmbd47EKfFA6CJPPHhshSych7
TFpJEDsh4P9yu4mZQiImEDSD4rzfSpZJvkcW5Hgzo4HyEH8HCuOOFMnOMy4B9Msw
shAJzr69KvKuRqfR8kez7GLOoqFgnVw/94vYKuIyzEoKMrDCcZs5ayzKcrX3zM4j
g1kcxXL3oYfZScq7lY+WHZ3Fz5uj/F2xwbTtjGOY4l7x70/lg2t0zz7TPegnFhkV
90ZBR+jLgpDYwIVJhJaq5Kar4xVIoez2y3WPiG2GyTVG4bO4HrGNNb4ol69UME5p
Sl0a2SrRpRmayVmt1xRmY4E86Z28CcfyJyZn7rCIRKjAjJLhWGvniWcjebU6iABb
XC7WcRKEaE1E4EwTC/M7NChbo9ipkqSZ/x7qvEnb923pKovZVP+r3Bz4FYh3ayTw
HQr0atCEUTUJv3VUjbRhjxsYDB7/Xo9ddV7MZwehjZSG7E06jfG34OCuszSCzjCA
OP90Mbg4A1zy8M+os6et3DTyhLLBM+ZQJqO2DqrABqwSgXVRY/BqTgt/iJusGZaK
STooydwA0/B9EdjrbA+LKaWnImZqCXfyJxSvEKln2/trWP2jtQlwG8uLyXC3+sfn
jMLhWSpnYCcI2NMqoRqRRsy9NaEwyMB7K48Z+PHjuRkdLFD2suagXNCd6vUK9PKM
cXiPE93dBmYNBH42qJ65CCixcPUMj/hww6QYzG4mm5D6Ku32t9kjeSx1RP2clBE7
2ACXBLWJ72nu+/5hA9EVLGQrQ5obi3ciKUciGKFs+6mcGvifIR2fstzUWnZen6kv
UUmDbL0SByvCznKc70XtGzhEEaf6R/LKp8lJRW1jFXpJB4O++0A3dd3rHyZcpEr9
NCiZYqEzyPnLczd7MrZJlBSX3J5d4EGUsFLV30wAGKcrXqKZPKA//d6nDK4Hm5kU
qKTLlMamGj0B/X7nJqkdnWepCwif8chlexOeoHjedUhapgjDBzJp04SWKCC9lckd
s6HMekCI/JW/fmHZl623H2MMTtNZGfpJ/AD+zYB3oZiLZ9kTAwmeOYh/zNBBX9i8
YeTmAx17C7w5Fmijq3g8TNnQprOxCdPFKHI3o15/860R+fsVAomsVUBTxuT9TH/F
+mRUAaBg+oR0LdjA9d8NUCJ4b1W0AyxMkoEWsQdaVMDRrmfC9o+xX+g0rJoXY6hv
l6k6MzoDVRE/0YDTzUMy01lgw+CycxUQvfosravW8WjH3NkAdyNXo/POnYsevjOD
aszXwajWqgUtm+FQ0XRRfKyFBcJgXbitZK1MWCNXuMXLWdB7TLb1cb93sIcT+QWH
h2ciag4oS+Ip8dZWUrkylITzTL0FrvinAiBuLBfRw7ClKct9sTCFieoYSuTQnX8F
YzEv0LQN1bv52uO3EA5thTJK6sBlTmE2BbCsf964Y3F3L1iOeH74mnAv4LvfHU1Q
RLfsYEB3pyLvvyUoFoOyjsn8Z01UDnhFKPONbdoVmjc0Pd7Q9FM8iB9V6Zuxf8pr
h1oW29Nd0nMELU2iNAKuGS4dmVEJXd6QyZJyAbLy6xY8U4USUdSBNxblaFflBcv8
3P39dv72HEfJLDH9A4SQO9TkQQMaoqaIdgVYXNlM+DY63Yst5EDSRtEfpQkufGsx
eOJWpSrveYvbSKMQOgx5/ycHQvOF6zKQ5AgvksurnLX51YOwveqkBdfRvR9C0wrx
o9DL/fCKMsLDx+cuD2biOrQ3tM6o8xmMowOpdcy5PLwJsdvb+naSAGQDzVZKtISK
jpkwIwXiuxMLVlsPqTXnOlLMCZ+irCsQLIy+Ab6XpvSO+ZZXo6BojTQn1IaGESx4
LkU9ZEIvyhrso9hiNCTjCmAY+wYvyr6ZeapdmggFISY/6zHWur0PvkCKJ9mTfzGJ
1AB31yKUFrXz8rFxwmkW9pzotNYxXa8RpT1bQqb2Fxz2ByXXYbfjETMy0f26kJzk
PwnKjbTzX4umosTlRdxt+2cSOAaOXGbQtEqshuvio/KgSpvICSag1Z3deid3Pp1W
R4sRpVsSnbtk6D4pRc10RH+5ipFoj5zQO1hc1Uh1L0PhBup2o2sCS0xnNP/B2JCL
K2iZLLglRNeY6ypv478IJbAJGMf1D+ql2RItxX/6xbl/f6lRCRn/zmcaAJ1vkZ4t
w5jvALI4Py75UbPaVlt3nPt13O6ym2uV9WRC0jDwNiPjY8JQR0CBS6vozndG+O1/
mF150TOqOiYB7ZybPBOHyTgRiMN+9eU52UVfaPQTCfkMnHMsvlHdpx3UW9agHJQB
JRcuPiPwx5ZqyJ2OEFmzmSgKof4S6UHB8Z4HqM1ZznsSCvyfQ9cPY+afS5YMctvE
8jiBz1nfA4hjMhgztrVbBsycBxt64l4J6deNuV4kwkHKO+e0rS0tmryrMeb/p8QJ
OvNDewED13TLq1odj1kb8X+gQMVEEHUVHsGX7/qPZD/+OnkAnhInZ5dAo3gglAMZ
wIhlSZtVFo9SsdGhMrg3BeNA7JRL/yFntaw2j/hjPNkzHCOOaqKfMg5lJZDQdfFE
IpSJbwZG+RhUxhtZxFbZg4cH9YUB9Wj5duwO2JBqWWcEph1rsIKKe5AcyBRQI/wb
W35HGfrefSOPs8aP8sjWbE8vP5dx2VybYanGBFZCsFuGKzsZhPj1u3xvxZF1cxuM
IirL5IdwTs+Aad5nxoD/gGNESFlBkDPOgeIYBTR4hTXRpMfE/Kid8vahPZHZ/LTH
zzpvK0pF8IrPiFSBgSSvjJBXjj3Y7QwLTOr6JgU6ZgzP7G9Hgbb39Fn+D9VtXY+w
8GTVaZWe4v45UMx0EJ4NDX9MhDBl6CUlGox6luxFH4CfWzkKLraPLodS2VEBd5pG
GL4dDpSAzvUxZx63rrESvcZJLSJXLcphuB+4n/Y5UHrk76rfHi8nxTkURBbR0LZF
Guw7zfASX567+0rv5Nf/N46DRn1teE9uJY3Lf8PH4fk62wB5BIuVaNpYiE+s3vAX
45kuq/H6WZUZWB+R0tugv889RKprALxQmjo5MyZaUWiAEPbJEkTCKCrhiywN5jJL
8r/Y+Z0d/4H87M5GbSVQcjoVnKi3E6Or4Dotr34DczwvMUuVc0svx9Lj3dv83x8R
mFjz/rIkI3kI7mDYmG2ScvaW0H2/Wq9aLptEZwzl6hlwfrFZbVIjQ7sEdFDg/5H3
telFi03Eqwy8jtzuUDstMHCruK7ZfgOQcko5F2smQqKP7zpiPGK4vnjXMQmLKMH/
ITnqHruQU/P25+80UP8zdHuxqMWK+uQYw2f3fMMenVeRxiswjhxq9BeufJ6iPjTi
+izVJrMYwGhoFDR76osmF4zqBD8qFrj6RUKIqetSesXvTEtZGIMbGlaNgonnv26Z
nSg08TuCYOk2fTduL4J4rKpJe+AQfDGB/jKC5KYF0KuMpWjXg0t15IENat7EMlVd
oQzo6RHot4ixV6miTdVR8Fryv2Xiz+ZWXDUd5af1ftbHTYMS6nwf+PZ6ohbOhorv
NIZm+WKvJ5CtWyJajPlk+M78nUGEn2yRMq1YJjn8ykLt+Gp6e3mFfJQgbYorzHeZ
0fgl3klN1xhP4FPs1DSr0vXIbPheofzSHLePMzL+2eA7LylYR6MSTe/aUJWLphGY
5kEliqmG5OhGsyKmPF0VCSRdm+k6wcNKFbcSypHmNaHf47QU73VUGd36UnHcPsLg
Z90PcvveKy84QHTHSDhb4N2pkwIm06cl8N7KUdKki4gQM2BmwLlpnrQHE9uxjaPR
TbZPUz9sIb8YXaaTmSzJcM/Oc7Qlo2isdfcYgPbs4czixR1/s3FlEOxlaPW0Nzba
m6aZ7UvTgxIuFlHHgYyBbseeaifsNE8xNwEFQJydcvOwV/T4bIHn6IDht/dCIhCq
kbTx4tXhV3b3nfHWyLeX3UV3MH6nI1ARMkzfnDZKXm2MWZ4Vprx7Z+rOVClRhJId
Os23WLnU1/FSHu1BWJ7A8+V7W/bv2kj+I1PFEy9qJukxv4/ilJIMbn19jtqHnNHC
sQlTHtBG515VX8FheDePEWVe1W6wsJgOUiwgIkUcSwogri6LtLN2Z876P5g+D0b3
va3v+/+96Jv5nwo2/b4c5MFbzeaH+x5s1vHrsfqLzxneRnzX9gjCk2nv4tdyIiYg
UVFPST0NFjjdtnDK0KqCdzehJSKm2UzESSGJyLEOEFRbfJhH+eSCF+1VKTtuDyR/
e9CfMcPBACMFH/47mWJwgTbXIO7vyFscQiMe+ur8J7Yb7UvplKFRF1O5rsVY9Gz5
egERzpHls6Mv5VrDFBL9FtIYwWMjXwwqKpzVpjo0Mbs/n1PB2GU/IpNdePU/85Bk
hWTKnlCCahdXn+RN+yTMXX75W7RJRLwLg4mgYZFTTmcb1tsvSI7vGgvxvBGOYcp5
eTyd/c84rNggpNEeUZ3pT0DXD8nShQRhFpWI+HgAJt6CtBMWOWKhIstnsw7oq7we
KGB+AvfzDSsAIwenAoA8OevQvvOxsrHhdoDZ1cEvJqVtEuwz02su/LlJ6ZwNWh9r
mzYNWrG/skrgPCS/UqWzILhQ/STV9XkctxSJXhr28AlhcIkmh6vD7UvzRo2o1IeN
zeTynlUw2QJ+i2LOX8/QeaSop0MFosy+uYap8fJM0a79eFxVSY3nTWu2QajymxOW
957tTDH0ZSSC3faBL+OQutbAS+RzSqBwqF1e+xjEnw/dzmx3ExUnKNgp+/6LCKlC
9+9w72oznbhx6Wzcp1nDuU1nmRAXxXyRZ2zaXo4ng1L9W8TOY1pVmRQP4qDZKFxA
G1gdVH3Zrk3sQflYPxpvusb/oPQ9k6vjE1gO5anNn4Ky8iwXCM9XMkYyz31KMCsn
rbaD+TpqkDoPeCXiXSyjkGhFeCLGzDkIaaG9DKnvaTv0koG3LTQdL5OQedy4LHbB
+XBsV43XocUJw+Pi5OsmzrJy8lKBJuzPDN1LLD3N+ov+S5VpwvmNe8VxDOK8yWLO
SlE9C6Dvtt+LB8Nkywf2DNbuLsyAnCswgMcQ8eGAR6PeBVWhXQnS/gLcd0maKBvv
apV0ExSGhnY8zSut8HLrTsCZVq3J9SsZXSN7BzJvs2oEncI7bkdBIeSy0UTe/0Wt
0F+KIDVMdVIIp9KwuNaZg4romq5BxGGsUOJxE03ULP0UOnVkg7K9P4Q9S610LTGq
QEuDOfmON2tJ1laLndWEHepeYF93PTd4YN7+EYiz/Tdz60yIINdMPs2OCTCS7be9
qOjkWRsBbe8Z2ipgi2vSaFmOAyYY6zOi4lwV8xkJpg2YmwtLjQ5B34uZ42uTLcks
bF5kAtjv9YpL5Y1nndQQR82vGJGEpPYEVZAHLneQ4NTUYUrU6qMJgkr1+UFqlp9j
Ktm5JSGtuc1omQVhQIWlP4p9ODs2q08v1ZVZSx4mEfBd2C+P/0cU00mxpwYuvq1B
snvYMWMmjg1CE7B5byRgVClBQqIex1M3txdv4eVWK+OkS/KmcCaAYKb+Zc8Jg9BL
ew5KjoI6kb643uwxiboDeQVRyKilqaLo5EhdmVRwoEDUsAsGSi1g5AT4ucSA6NAi
MRbcWJ2FD6hVhCGh6v9RHu+LSowpN3pWT37rP9rJyeJX4tgvd/GIgw32kYO6RbVA
6gUkOsYgDECTdC4HiN9DMhvbxMjPahQyfwYnH8FN7cLkc1aFGW8pkDLWNmZ4F5AO
HSgPwGLE9EOuWTUjeyCvAEjTfhY0kUaRtI7zQDTK5GuU5mablFYLEivkRZDyRpaj
czU78vYzKs2dAv5iOyOYnBEnNsZWbcQrDEVP2yC+UwVWIMgbOmD201/weKJCNMuR
xS0zliOp+zgLORxiGwj4J3ZP6x+5+nwDHAnpIWMq/D/4uGyRApWFaWuk1POkA3Pi
U4UzO+mNl0nso4MUp3kn7v3pr9DrvQk8rc9fFGoLxE+6pBfcxmVqBSnV8x2TVnLj
qrHUKBmj6qpPmfuPAzE1YE9M3lDWtYxtbDWE/TfEwKeDq0qPqkRfieyhnRD6FWID
KINRV0uFEdcpFEeXoD7xIiWn199ATjiQGaSjBkC0HUMUPUv5ilneC5InrbY0SE8n
Z7VZtsei+ABcJViLGS2vrS9P/VsIeMBTGqghZfqzcW+fZpYLSuZVOR6zmT1oVGLt
sOPaJwTN5LfqslvFhDONNxjMSCj2k4viIEYpp2WJgrLNTxQfmqPOV6OLRGFEcUyc
Rg5x+4PkzNLOUau/LecpS3Mstp67UY7pRwMAz694jbvIQcSgJbL6A+TrFkUkgXOn
dBUh9fm2QLQy7c3oRKd/t0jcPTUC08jwfBxjp/ODLqQmuEZP3kTkzCIXR8rFKfUX
ldR9f4Ojl3NxSmoVuy8RV+0qUULfdfqjlfFVM6c6+aOqgkYyadADB1ZLyPExapEh
8T1xUlhkMAkiqbWzBHK8xFfOmD5s7atbC9XG7R/XMAYQupIHObH/bayDwQfQoGhC
st5Rh60VwvbDtRn8+dUesPBIdM4w1FwFW1WTL+82a8Jwt/WFJysc/ZKk+TNUoRPL
0QRzswdcfyf/30tNT/M3E2CEZxpuHfxMP+XEdLz7cCsCE8oqIcBrF08bUBN4lwD4
Wfeapc4MzzHyXmpVWaZ8uTiEZiMWNm7GSjc6QXEM1vRyUGEexxLaqVPsU/DpFPSR
lxATKq9NAqbXk3YdJQbqzXAiLmMGAwhlKf0u291dEJUr/n8ypWZ0sqVyWgjz1JRH
mwVF2PnYP5M3rXvinZARnGrlGG0gyNOpcqGXz4puPfVy+eG/G8N1OB/HgO6i9wrW
3+fgU8XArZUOWQckYaqcZHwk72p2GowfcOjVk/kA2pAoQ7g1clUmzek2ejTo+MRQ
jE1aPcK3OVZouoGmOXDFF5WC+ighvIqRE/X0LytS5Z7N8ruSLACIcBrf8ybEpCLR
DeHf6IUlI7MW1YG0TYl6KGdurdz1NoM738TV4u0shfvKDDjBZ5ISgV2xL1NL0/Dl
bZ2qO19NiOIega0gfIUjpi1g6t8uosG4a6zJSLvqpJec6u32iRn0pTil2DryvO1j
HXfbN3FMjnhHYVlvfhStdWSGjozzddi/sThj5Wld1mtMoILvLA6fQbzjCTKeoARw
+Vhzt2qKf8TPtHrS6DBLh/dz/5I3bHPpyMdbEB+EeZ/Nm7VIjRuFnxk3tZOkdtdg
/NTl2MGT7Z8vGWGEwl1fsofct0P1F870uv8xb0nEsmeUi//TgBgoynKXYnhbI7xT
EW8KcpUwLihKu4tTnsmVSH4XPzfxk1dnzPvbr/xhCxil8i0QG3hQ8nz3x/5VwFf2
b3MtROUZQf4YHjbypy/5CW4hUo8/7WWIdy2BhBKS6oA/L4KU8ov6MqqPaFSoxDnP
LVfRVx86biHnXj8XTdgpzhxAY38CJseOH4Gst/kGNtEYCpUXR93cVhAZLLys/LeB
V9Wvcd4s3KRr1raSOmdsKW9RMEXOmssZEgd0COXtlDkX7YGAzIqk7wax/873GVdS
dcNYbzWBGsrNUgBkUrfT9S3cM+b122gAfSXaNPqUnc9rRQ9O2/nQ1xZDLdBI/HTo
wY/nTZmf+I4XrIsyFlaikC3StJBrWHuk/XYYtCcS1k3lOq3fZ0VL/SJS4Lj7jMKi
qZfE2/qkA3jzGn+3Bvi7geuK2ahuXR5dR+1wkeQHE3s4smpltCD8OQ6jMfWxxbKU
UxU+KnbhiZO3xmEkceDKsH2HfuQnJQfM3muEJQ+PnOrw3PZQGXvhG4IqHYvePYc1
Ob3C+zM5RytmfLfOUMEl7WLwMbOZMjwfAHKYqSFp7HsHTBqWTg68MxV2vYDuvZ1k
ftrmETwxE1z1aKoTDWEfYsEQJDTJAOHI8q+1BBW1yjUZzIDPqBf3jOlLyDT/HyhD
Z3/Wqjf3p5FW1I/K8ygv/C/byvAETDZ6NdjRdsM6bzfrtLNp469/9Lsv6twKsHln
DHfGANQvn4iKRyKZl1AYZGkYP0b52CFeimbAO9skk0/vCpVMPjnsDRnw/MdK98Ck
0poF8FuQstrVvqEM4A3vjPd3ryQ0l5npDp2tZ7sSxCc8YtuS0xlHK5kUEVuGV/JF
PR+Lp+CW0ycBySh+ffbgqPmt7kqpsoPpXW5aBnZvisbay6MKsp8J+tZFbYUrDW43
vrZ9SD6I0s/zrg2V/FmF2ST/uWzj1JomOUjwGuxnYUzO3z675d2SYjIZFA+Oi2vC
gIf68OS0jyy87mFXICvP6dweVPTESJon6wpJ/AoW/KgLq4vSi+IkvKUM2iu9zgV0
WSnm0CzxW2DJlPvbZQ+p8PSk2Dw85h8R+HecHU8sI1rN4zzzVE7wJzYXPUSEeAEd
ObNR/jK3ibtiMftBMt7L6gbJ16mlzJaerjdyuAgyEXlgOzWeYWpw30US2YcGNNe6
M5C5/zhl+BQyqnNIlKBvt2XrEJ+vxSnKJ+YoTIxOcM9NlsGYUAaKP+/DHQBsas6N
+Ivi8WVwRftHElAnnh9ebdxm/4iIY6MxbMsbxoHOfgSt/Z4K/6YC5+ujug+0p/wV
mATQhsyHivJDkfR/YsK0c5oe9LfzV4cMuCqHupk6GVl/hhXxh8oTgNiDhmO59DLr
CYZe+2ylYagMGJV5e0vm3bqiuAkNvhzpnVNHXIyOiSopR6TEAX1PKRVO+/rzwzkF
jJQ0BfbD8C0EiTGP7s+LBFks/MA2GooN8PsbJvYNW+B8DcOMJlDgTu9i/JOlEvq7
Z2jyZ8/2aMwgYTiEc+0IvQbtfFIvflssJRlgaU12O0tHm5x8ZcBEOVG8ANuYhwUz
pNykHro6T+JBgf+Y1QHxLLafAXUynX1tfi9W6jPM0MsdnCXfGUU/H56fmkFjgXo3
ZTn1LfYkIfLW09/4OM1zjIWpQQdEy1L911Ak//5ir4cJ2qwLL/xlmJu2/Cs5dWVh
YD4J2iap4MLRoQtyyVSZ9wtfeUT5vGt+gIIxJMzPGe7pw9ymsqN0CwVDu16uaBuG
MAaZM4dFKMOWgOIQCVljqFyH30tQGzLQDsvsN5/06PZ87kkcP5aZTm8Pl1UOLCeL
xS6AyA8EfPs+yOm++J6wL8YF/sVS+B+Ub8canSHNeTIbbNGglRP5/SKfVo2CfZ9Q
drMLxMOyE7sHEU26Y13l5BRPw7EztHsCNLXC7WGEaRJ7Zl1C5AgD3bZEtlFY9emO
j4Asoh2SeNpX+B7R2mDjeyGajntOumZCzzmUWS80ozvOe3WHIJ3Ai6/uaBkTjrst
dpBpdNZG4jflnF/WU0xjil3Ng6kAMhwXGNQ2u8oHI2JchQ1IriSg3jMImDLA2JHZ
gWvf6A1f3lnXBdCzP6mw14fJPUu3+DyM+C81Px0LoBh2MjYxc9EHzjqC65pVZtKR
2pnlhI3O0BMWsAEiFtuQrdnVU3BszzIWTFRjGYs6jdV5Yy1fP4ATehfJPQRuEslo
3gwxzdlSdZIt96fNlRFfF30MCq6JtuU8SXJYGY/z2WMbzji9H0mtr+E5aq4rggiK
NVv6tYqXeBpP5QD8wDeI7z9v3q6BfQmmrc+QERmOhvymEBu0kUM8XDt0bxQ0SXtl
O36hadb8jFe01a95HnumQzwaYJdqY/OSLES5Ti+aPlLouhdj7GR5aMaBsISxH8Us
ftB5CEwWWgT4enslFOk5f+BrBdX5OZ5xFc/NTiySZQoL/5Q6qWy2PxUv2KKT3eHg
RdSojurEeG2Z1dz5un5mgXtwB9q/s00TH3C42+Rs75Uf40nUjTbL70MMKrvEhmum
w0/9tRXjRgoVwOEttTC4H3lZcJnQ1d2UYVAew0B1rgzWGmg5/JJerxEla49SG4Rg
z1v+YYvD9UfyDQMyK+zhmYsSytchzaUWvxyxHHd/Nz3AdnMI4oXyvVdBKSjDq8DW
9QubkPg466ynjWqHytkPCbpNiqHaZZsHJsPNXyAiWdVQ543f1TB6ANynuud6AwkH
PYWSyZ4kABW44TokXx6PY7oLp5BYwqmlrbnP16YlLL5XcV1185O3fft99kK8Cdsa
u3254Y9FI11DDULvUhZRS/Kgn1bkDWEmhPCc5T1vxQBE8O+j3SQu1or1Q+VGbJMZ
Tw02k2h6o41CSZ8DV0BU/lEPv6G4j4EYYovZFP36H6qB3n7gzeOaowT/MGX1NH1C
9rsmUyOxOGG6Kky0bOCs3uofA9kAmWX41+U39NNOFmnWCSPhbrcyXXAGqJfW4sGV
uLAq1AlPC2KUqVvayo45xIOlUDW+XkHXGYNj/15NunTv8NJPY0ta4d/biB+bsv0x
4Z71SyAV5NwbaAxQF40ftIfUY60DI5DXxZ1V3raE/r13yktVkej97CTQrM5ARByE
wf6YQa7+nIhRTOXxMKsVZ4De4y28mWExwGSlfzFBiENWYDBY/yjQWa3jMIdkIg8U
YEPFp3qL/X4MOLwTQIePXonATrel3yrf8c7kEC+QwvtPp8dUuLz/cD4j0kzLGdF0
0dDEunLtPlMjDYuiGq4T+XoyAI07tzThp2bnB6p2dQairLKSmsFgyxUPnZS5vEJ9
LnFAdxnAikoDlhVI+SyIjhzP93hal6ep1znpjtPTiL8L1jSajWkqqCjB0BAV4yMJ
vXBf63/jp+Mh9i0hgnuVcp0mQVnmNYCyS9HHV96Ryt5gv/SM2Px7gEuKv9uOQ9bE
Pr1+VclFSJJGpdaq5d7y7j2oXYOTct9rdzhKxtc926pxWbhuSrwPbpgN2RE2HTmw
MTBcowZOmu6SYKfGH9UPN6N0awtWq8JSN1QIACJaNMxf7lQSUQ8RX5/qcsQvOnIu
cWwXV4YdjgeFy6AEdUAXVZr2PHLjB9oAbdXbiElmSYYmDxF/Z0sJbm8z0o0EZ6Ni
49JqFzcArMVQxg48uYIGalen2A1JHMMsBiEeP12E2aqqSXPSkvfxqW3xBLgMrZXh
GdDE9YHo2IROSGnRBdwZAbSJVVRCvImK0YBf59BfJBFmWPCioLv8YzjSdSrnKm1+
lOrvG+ht3OKBP0obmqpN4E5/gTopCRZpBXd3DttoSHtFrM6HUP6yanqCG7k0yisr
gFKoPbHULwX7naF8moMgUBZV/zZ4gwsJcJyg7xIK3fXXHza5orFQ0SAFNJOwWgfB
rpZ79JFMSz9INg085gayppzCK1qLZXdrXQ/c4YIhCsqKdGIXCGcwDxYVU7Jz+vCK
qOnCwYHWfJhw/tQa+jcE+e2qEt6bqxQhuXkOGvnmGvQ/vJIoIlFYlbc5yT8vdz1n
L35DBf5IP5UdKB+baGq+wcnkqzxGxGsTR7Zkfscq8pBauJRnKf3VVjYDAeZn12rO
HvzS+niyowUXH/AR9dq2vn+s4ncuAxFb5qZKyYfxN5tIspXR28Sko0G6G9OFjtOd
wcrLMEdmslHKKZNNh7CoGvES7ecbvCPxiQR+QKcFIEch3FuB7WHF10t1cCnzQqbP
EPSXqWyLJbv+P3ynH/qGBZR/j3HruP0pYW6R3s2Z+WVBk9oHvPWGND3vbXixvDMb
PqIaS8lroZpNKR5QHBHllHrzpdexdiHAx1Qm/V+yTqFeJYPAEPXfladnyMcHKzQw
XjSGcsuWmxOYBO2ahdVyptArjRTCl65iuB4hKZCa4GBGLT/QGkQTFaUImW/uEtUh
TBsOA7dpVUUfohbdgxtCkask1YD/VxS+WAbiCZy0Zt54iVWEglQog2n+gZm9TD1A
BmvBxk7/Sj5rf+JV///Ds59HzwXP9OEIotK20gbsjzYzsXbX2e5REdhS90Q3s9zj
ms5RExUdK6q0Ax3Q1l2/GUqw8ZfYLNg5wrOieIizDrygFcmu/K29d8RTBQZDDVl5
N+7GIkO8q7eYhtA73FGs+1JpBSjoxF3WylKgvkXtEHscHqiaS29/sOLp4+6Bv/aM
+abCIxL6eFMSRyqVz5fc4gJwH3dVC9LNl7dwIGqz+scOzkbyyPFnO+q5KOWTGhfJ
pJ4M/jbReAuFCZESnapD10Br9wYEOGI6985Av0g+gI52wVKCnQvoA69IAMhmeujL
QtfyDH6TBWpam44aVua1kOSWZ5bOFLl8DCi6csmmATvozsZ2Y2shV0RxYW+lT7Ws
Koh28nlDYYMEHXWKqB9yGmoEJ4WxNQozFPRUWocG6NTouKWxpVEuJ8O6xj6bi+JI
+ULiI1Ac9qPNAaMN6nksxbxb6UZFbohau3PLABZItiPZlPs5Iz9sbfZdVvgJB3NJ
hRobnRs1i6Kax+b/AosUtw4+UGra6Xpi0RpbOzSC+fw95DNenHA36BRNzM9Or7/s
t3iADS7zKWk709DzqLsdnY06pRYXgut5XJTYlsSH0C/itYdiYKoB62HFoAqss7V2
3rPqR6LIRpxHCFYXOMOPK38f8FnsRkZff7gYvowrSXumJLipVLrtWJeK3KORWL8b
NlQGY1Z3i/n1g4VTVTIH2pNxt8Pzo9fNWI1MMb+EtE/fZpJOBKY8HYGcC78yhPiq
zn+eRuLOZquhVp+pPR3GI4AnAFg+uZ4chUGeHIz6u7GRhW24p77WtXV23HK9Irhj
rc8lwPLmT/Sw+KPBjctjFYTdqyEZM36APNwccNp13QssdREBRUmT9e4jhZmf0ErM
le2sIBTyJt8Bm70PCGfoUgiuBoSIy3SV+o/G64qMaAAPLzfmJ/pr0fc2U+Uxd/vp
S7ynlEwurgozoAk1YTaiIPSf512l92GO2r1WFDk0nVVJyHZqEhWfRe1wvMjraW/O
yhFcU+HQ1sNHppuhtJB9OORC4sM2b7gFp8wlASE1viu1Fqsm7xg9If8zRODNiHVx
r6xsb2EWA8Miumpmnbl7oY+akIzNBZ9LmTuFuMQzcQ3kNuiATn9Bf5nS2/cFS1fQ
L7SUz60kcaLGbFpiu9CY+zd7VN+04Y/jdKexrsUMp5NMiO9Rgc9vHQTzgnyxF3Bh
cXf1F4tu1a90KoZMcdbEJxVzhu4PryZs8FMwBrlY4QWIOHot0Z4oqHrCSZRcDq0s
nBjV6Sd6cNA8ZFFq1noQenUL7HHwCE16a8Fon9MzavM4VsJrEsHKFF0FBZGO459n
zuMERhH2chM8/l2dgunaMNV8oov9+EoL2yG6Zk1Re6RCqeL7hYXwzkXl2qYtHXv7
d0IqFZpE360ELnf5ZwWkFZ5mXSzb0ASJ3RS6ShkBadIWaXBU6g/nMO3i7Cr/wIpZ
w9KNZC9J9WIpa5VccdfVTd3f12erlNPG21VU/3v8niQz3cFM9OwsBSpNLYENcHEX
7/HxEIvEBAYvlzimNnKtq0LxPBeUcyWrV3GBO9nvxJP0Up/2ZOHZnGuB1u++vkPp
I0wQr9dd+jH1xYzEi86LzDTybEHWlCJeLEOYH9yy8IX2ojbtuhayPLPUqacWMat4
FfMyyiNfxMptsMohMpCn7gWTSBqnMA5HBG/IaveyTrGhoNu3y9ikrra/bzRBzuxV
54yXm7kMQJhM0YRyduCetDLzKe1CZjde09ajJ9DO9KFA61WoMANV4AbtnXyp2oT4
IlTGNI4xwmjvuspI5Em3wjZRFHLbwK1oVj+qNrDttm8=
`pragma protect end_protected
