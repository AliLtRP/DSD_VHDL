// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
newZGTtCgxB3BiXggVJySdMvUfDUHdNyNwvXQvVuAlWVVTOCNlMFCsw4BQsijkxN
QWIw80yDak9RF1bbKKY8NCZbltsBxC6emBKMacCEfzWda0mDtrX1Vt5HH2lYgPh6
0BdjJd5SofN0/ZJj7Z1FuPpzWTnDLqAUGP2RVk8p2ZE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9168)
xB1qTIynsEY7jBUF3iETaAFJ4AlvCFX9IzUJUmszlJlUvzwG01RY05oKDbNbkrcY
YfP3rBwovyebXOHQulmc1DpN6GHFbJORtPHFDC9UiRkmNbpsTGWoPg5yYVc4rW4d
mBpL/vS2A4JOuMFV1/PVuQVgLoXHFx7PD7roG3zp/RVRltar969ISHG7IcchygQC
icsSFOkKjYoklq/K3SVwG1NeCYdVXl2l3cfqQod4o/kUce45S56hMzs04a+bzhmx
1xBPQC9UZkxhjvqqziGMUnkkqkDLXUDRde4Sf0D8i4X86jDAaGkNbxFwx1+tXRA5
IGw7BFwOilZhLJi/rdwgSyilyWTJwHtrbqOdbhrEvpATVPx+G7csvB7OemXQBQeU
uDqEx6R88VtVYd5kPkDIsjdaxlUU14RPo4CagjQH1B36eqIomk4ZeniS+CEI6vUR
fv5YWB3cVdLxHoZ8oD+EwI9x7+ACMzbCoaOooAGRP/oMZXE1Ry5SyPI1u40+R6+C
DyR/uXesEljIWa4A2Yhmh/TRq3/TLVHXxKilR6thCGQUI2CGVYMRMb1WczITPO32
RxYTxXH52Bz3YRr+7upISfLhha21xT5YlPFNm3+mIslgBM3qE9YY0MqcwL6SVBSZ
ytBAyClT0meq3flqZ/5ozk1wGrrkX5LlOnAj5n5vTPxXYFZYlslkLjHv5blEGJWW
JyYfDmFxjeRw/8aXZYgYfh4L0g9cX46bVU3ddwlLhDr97Z/HmCpeTvB3QpSC0zYK
Scvc5H7OlKBB2pSqplRzz0vjTDboxXeiMvOsfWmqKvHTkOuxXp/tpcq1Z1Vpkafq
d+TCkNieE7r/xbCi3B0lOvkHpE7j7IFPaJQv2/eCLHsLbq7qJBszjU7NHZlAjBea
SImnG14Zz+2rtXeh7gNzeLLlaTyVVIAi0GZEt7XeExP3UxAPbJUAIR5uhdS1WmWF
RlJzPSWjb1J53W7+J9g1EWTusVfgMVL1epVZB7l6EwH0zkPjuGpilChcO+/I7ucL
MZ25BFqjsCwkoCNWmDjMNmav2Wfa+dMAStIGCwaLM9Q1emupaIeaRq7cCyCtRDgc
Kj1EmwCWP7BBWfxFWDbezEeYeXBIDW0fRMPjJ/FDb3Y6fJGbM9AyLcRWlo5elQ0s
QQvyeSAl+HmXNo7qn6umoNUgwj5sNggx/SLgY/+iJYtc1wRpugwZ7ECAtTS23w+a
y/AmIof36N0wqKwAH+Cg+7+9sYCCuye3rsf5VnE9L3H11hFThITkr4bfCPCAQkAz
zkRNBxSiVmUNKfuxGbsskMtZWvX89mnY680Q0JxdaTyAZI2BKSsv2/dGk8gN5TxB
wFoCzJMmGvbnJzGehxR02mv7LLnWDwIfOo28I6l9eTTUtmvaY9dYMFHUf35QleMF
3cP9qiDATuvXykYEzffz25jXVZR9DKALciFPRaSjOJXRNcU6Fa6MRhaq6nRDCiMx
TlgJqkmY7Rf8tc4UdmY2gixWzUPt9J4mVrWklxG2w5v2CeksoL55CNIUJZKhBdwH
KpD4cjh6V1CojkZxL6EOlznGQRTFjWHB3dXaXaArwCtgaXj+Ug+7n4y7ebRtjZUh
zhTYQEJCjVoGWqC7GmJhta0J84bCYuARaOLDaWp3IEVpLWVJ4k+fpXgOrJ2v+29D
9UAMeBNsxAiY4r2J7vKKvDfknm0wPUNmoX0KE2WWd94Jn5xryyM8uzxTJA3sxd/E
BbO6AUJ4eumMDbCaF9NWcCGa6gcMQJ7mgmE4ukAFo8ctPkT67RPnUx6cYif715zH
Ic8OvXeCdxrO9FvVJsHybEYooh6JgPa0O+C4WhMr999adW38+gmrOdItwFLSU9ws
zX9ZvnfkP2Rvl7VIecJQPQc98k4pLtx6VHJOrFGZLjitRfdTGiTr1JJV0o+2l/WV
9TVvAdRaSje1vTRixuUNlZwOVcmH5RG6mPIiueWlOo7fSo7ZFx2zB/438q5QFy0J
MM1KwkZ+4Gy0+ghUILAjjjbRetENSn60yvk4EUW730+NcDad8OerqL08AxgAZAXh
FnnWG9ewyaEjDLElwJyjr/Q7B4brmM6g+pgmT7Q0rcHZNYsM3UG3MQFIuPh2GC6V
F1JcsNJ1EIWCH71Y2P2ATsznNZK45hK0Qo1dmzHLTRtS7PSnp/bzLssn0WjZ9IA+
2pZ+5VBkV3FRxGmfYwPSn58ndhq0LyQNjUuHJO7eHYwjLxyqcUUDOP0IFHQlj5JD
xsePJL+UX6HlcvqlNoVrJNf4nzPqCCBUCj24cFCyaXTFPQA/rJ1a8AfCHRGPjPyz
TPUXqAP3+Xm+TFLF65s/wsxukM6E1Nx3knz+QrsAjOpbmKqfKbO/+PTHxd5xcZIV
lvZaAiLtgSEpzfHp7aMXb0x9L4eiCkBgEAIeTImgmOrA+ehwsKoDjrQEdqEId0DY
RX2E3Vz0ZiAj6BYgHqtQSML0tJKfbE+obax6KdofgGipWGAaGPOzvVuKw72ojhH1
uw/XSEwAS8oWNklnSePbg5j27PEEVDNrxYG+yhzd4EyVSbePUgpQpVPv0PyUgIHv
7Ka8wAJh4FSLuV8yyhQKFg9qE8llqdVzqgps4nXN2Iy/1XnVADmepPJRHTO3sqlb
rRCqsYjVqPzXqYbnca4gf+NSUj4b7i6rAmeAVkV9kU/rlxVZwiUduZ8IHdbMnmQw
Y4GuAk/FeZb6ZpKvRTeYU7f5NWlFJIZLTg08wG5d1HVIY9smm57HsJAnE/EroeP4
q+iBN3g4GA90pHC9fdgCL7czZU1bxBm8yKhXZenUrDWlUzwo1MT7auL6fmIGMEuy
NJr4KHRCujN8f9Gz1D5VQZqbvrYkWuWcMzSGxzPAC4j9CJ5YPcB+CLpM7wEdx657
3tkPNA5vbMyn034tlkHM/eiqpmZlncvNJ+lEITBl0gl7t1m+DYH+TgwYsCCy2BrV
ozYc2a+WMBspcEbiFkLrXV/hPbj8dwLLxvG2b4o4g0Rk7c7Eo/yxMWY2mS8l/a9V
njAvL/VsMdahk2pCMtvjyEAiWszFBjLh4jSLgq8qgWlVTaEUBLtLGBiNgjqXMcJD
XyGnKc9sA4/hfHv0uJtweoWvC6GYmJ5WS7ut+KCtSqch2W0wTq5ruAPBl2h+/4oQ
bDldQfhsjectlwP9A5mgRR1a9Qg6Uh0oI9zjM2ARxb27BH5Apki9dzTbQia6R9tP
FHLZkbtFGf1rpu+1eTL9+Y4oho0ckYXgkt2nEFpbevCW4eRPHSPbE2bRZ3D1s2ZD
qTPNIxUTsQjfzlkHnaSg1+d4K3dRETwmn/rk8fWhQICJTyfNuzABNbP6m7ICXPUI
AF2WbRY+5LaSADV0Zdl8R5b+DF2SvMO2nQKDrph3n32JCoIuEqswl809agsjtf4A
QgtQELW/w8ebkvdDpjQzE2krR7kJ4BmwYL1pIahG1tYMPzuGoQedzfpPrXS4D6jY
Tf94zVw9/pEB+E6hF4vEd1lWmLwDt1xZ/hrpYycRao7ZSQWw9QSXef0j4g8Ux6Ow
tMkddUfLLSVsJ+Ky8a8cwCqbiboJeQ6l+pn1zgArUqLK7jxge1tYLHoy8zQWr+DF
xdIMl7pfFJxFyJjgZ+NoNxG1nCE2bnMqDgcrh9exlq0rujusQjyfk1hNi4NsqmXz
qa5Ji7lrAk7dyAotth8JAUwsBNpqrF8Dc6TnF9+g4GTYXsEL0ICzu5nK9xO26KjA
66H3KSctPqUhCpem4kuhW2PT81fho+DiT9ImdtE77wNyhKU0alj/YDveJKQZgCe9
hr9jPSeNGevBDz7JdgqBmfnSXN8W6owS4G3f9HZRsAT+wXOJXhQVgnS9G8x3erJ0
bQcuzCr9uxN03q26tvpUdLY61shU9rva0g/OrRLYS7KYShK/WfdT1r5nfgF7X8us
YYMsmt5tEmIKnxmDy+7YyQVwOcm2I+XRKjZYt0yblc9xXpcvXtTnt0vUk+bqnMN0
2xYkruDvxeFRlypwAUai2lAzcVq3XwGUjGhVnkClxrUxMSDZZvDrAKlxWIoDctSF
fI9BDPbchXezkV8yzhNSsLHlnPjy+Bym/6JvDY7VO4kK54WlOGHbuLKPomi6xplo
2VMxjTrHMnWZS65wXabcCwPnGxGqWpei64JQpqwFE87sv4CBwx2jw3XcL0Anr5uc
MZ/cv8xVHgWbA3HPFPolc+N8VCBBdQX2cC69bRWuQWzrYuE7J4geeR3Ky9mSRAmJ
K4BbGfAR1f9+6sPpgoa7ZcNibCTQxLr70rDYil/IzWS7GefsDvW0p7W0wHSObwY0
E9FQygxvqrTfHwmf7nOtlDDxSlthIFroABOhHIsqwBOgESzoJ7OKi//1jPe+MGfc
33r+NBndQypOlzZ5GfKvHLwm6m8JhDdNmfAP7l8GmY4ajj8STwWd0ka2euGTnnSP
tjHxwNjb8S6aPD5qgv5p+/RKf837zK2hiABC0y8h339vzaPYlMG2fnfCZFCK0Ofi
IubfB0ZQXZh/4DK3Yohi9794sCbusBfzxsyIB518rEc8uQ+moyv2TSYXHDFZY4+W
gNMB8fJwnmiF7BX2AsbiRANvcSK2q31re66XXJjvCeXxvO7pOQkAlychTnxUbIkl
UwDLpmbGFYTxxSZZasWF8T1dNAIyhagqK+Op3sRXBz2xCzJj+B+I+pkzhab5W9ik
ZoAgGTzfzGpiCqY6dsS9tLR9d+E7mosqVuDehRT/67vP2CG+jQtox3OHBFwfZzWW
wdVSWAvjd3zPdFzoj0Sg190Mshi8xT4B9d0PBF3YjSlu7zcLVUWH5opDyeqYbC0H
fWxurFloYYDkAmlxEua52zMi5tL4uK8MJAaJb7NxPZxAq1+dU72qsRQ4o/O1MXDD
xUmSi5MS8bpSmMRi10opgqBUi1gzV+c6zx8hO9ycwLfWw2vKzZU8gcJa9FpyX7cc
/hIWnTr+S877LOBQm8409kDvmu+RDf8wqgJ7Be4I1JhXSlidbe4FSmEbcb1FKsq6
x0882a5oFhQ9c8E8smM4cOeyIYTt9BWphZxiOAuKDVBzPZR6GqJxbos3ZAsm7lCM
KrNlK2sB7Vbw1KDsX253SjoviJK3B4QlIunr5zi8puSsmCFMpjGSOVwl8POBFOdG
mo1BJ4C0vot6B63XE+Aeaa74I6YF/ter6O1BN4M2yF4Af9U2nGYoP94D5ZxyVsYH
Xhg1ABoA/WHEwjn7tdpD2kWUPcn2escR3oICxp/z/FnyTn4Y5mR/wO+mqYRh9U/c
I7CmwyYQeULLBnHm94mAXCzRcYTlF+Kowm24x1YnRQgoPoWTM3fWpH8pv3Sqnlk7
Ll43TDDNaMbzYaFB1gieOP4FAzQLi9UsZkyiqBwuQ9xYXaacDWVEfKy5tjQxAKQs
zAuyQREg90lCKjBDOvH/JeUIbIPkzAc4lPGFFEcsnmb05uLrxDqSsGoRf6tzppGA
rCgGKxFpCReBp5GyGNhmBRfbxg5XQ/2satDR7N3qChfK8HUsw/uwrXVNRGTWC2Tc
+/Rd7mwRAJLAAH2adTnJ/cYfMRacicgYOGQn0OTQU2I6bnC0fu2H5egUYrPDPbSl
Mz/VbGZhtd82XcPoNjfghOPTx2L3o/Qx4f9Jkn0PxSqEP0+mhV9qhRBib9HnghmG
t2Yqfm2GB2xmaTXpuztBvdbKqKH7KGcrvEXn4x3w8VKb0WLmpx6z6FItRub+cWmF
getVAe9kSkrgbwHtx2eJl4CxDzGLnL/Ies1YyoZrbbZzIROas/4QhBCHeoBHEQut
SFW2IrnzrdjLKppNiGMTOwigFZ8hShsjzEUhY3wDKbJqasF4PO2sEVPb4u8cxGse
63UGAOxZHhpT9Wh7eBA5yG3m1+zbCNHq8qenT8zaSEYA4n/vA8eI1PO8lhl1s06c
M0jxUjqYtqWqQkRVF9Qb5chlY7F3UK6dPy6MqBr3ujkXSoTYDCREH2s6ZCi7Cvud
nAL6OZ7q2CeQW/qTUAm5/gSR185kVeR8QNKSL5e5A7Lcw3AiEFeaE1gbOk7h3ZtR
Lafh6dMhv8ABz/rKXpCUfb+Hmd+yHnERav2kTUELHhZ9YEEZ3lFGZZcNNwGKM7hL
5CUqS5ilnANxq+/DZOweKF1HWtyw6GWcFx3AvVgEle8XuOuOYQX9eaAb2/0riGoy
1zcVncZYeAsTi6SU3JohFrk6viUk3OtkFjdAMOom6M//UVgG2lCWorVtvtn59wWD
CX0Gv6sXJcOPY4x2xkBQOh7RDjPs/ffsf2glsxHyYHKzRhZLnbZqH0H5UT5W75px
bE4yJv7Syz12mynA01Etot0Qm9CM+SuKRjHKs7DiCxnP4jCXmjJkkjPGAHLO6I8V
EttBtW42w9kFvW8zx80+WSqkLYDbwS8MndmlJ8Bpdo4sBP0t7ayrKq1Bfyuek/8S
4oZllo5mF2J4CjwGyWFS7+BSnmv8bRoshJl3CFrAbUu9x0smjOrbnJkSr9e/QWh9
fRnfS7qjfnrDDsEIYfc0z5/hc7bQyeRnB86EFydaNh8ad2U+k85VseDCri+bA+sO
nop1SQu1Fj+jwL88rX9/+7jc1Dy47ykWGEm5nP/MECMYKkiYtVutCNMcoFXsPqt9
yR/RQaNn/1p5Gg9YeRiJ89tv9L+NBRsi4pKkvsJHs66ctWAAbHAw9UB2pZMVQBCu
2XrVh0ml0hwE/uKroe1ZOXlUrYGtiC/CsNyEs7ej05WMar7uDLjus0yZ3D53jS2S
SDmBroWP47um+Pk/d5KDqU1Vo9IA0HKCtLYlgeZOY81rE9hX+M41QHWukav2kJ7w
VbrrtpY5FxuBhjXqjC4yidPWWMxW6217F2etkJ+DtFCAO/aoa0caofLLyUJNP978
VUUdVt1JVqd+1JAqc6LM4FyyI/bPx2Mq436oQoQi5Mv52mCd2vrJk4UqjaVISPlW
dr5vl1rLI1IhxgEHeSo0x2B0iDqxFKhS0p42bBwLehL4a7K6j6NnN0QCIlr2EG0d
Muvd0kWSHqG0zgPPkuKX9K/cK1sP7wufvWbUgLo+x2/9fhltFn7TkEHG6b03sbP+
GZ1hKT1RFn4zciES/ORPnuDmDQbz0WRlfvvAzaEqezrN6motxHhQE33JWKQnIsIn
81PMYjT0Y5yHK5k4gqhnsjREZc2Wu/jv3q/RGzxy12dTMO5f2Bc3GndLSPWgSFhh
QGXOTCj3YDZEXNGeFwF6OzLYndpdaIQdFS71UK2m6DJ0JZq39OkepqudoHokpVu8
aJ4ZuoeX/9LMqZRqyhgggBQ8tv5rtzwVEmEUTI8EXOYlQJV+Z8ymh8h3jFqSjTzU
caoI8i4rwplJxDFhr/4Tn+CTE+JS/2UR68opiUDXsfpXso/qh1iII4F4VZsAuau9
1RWKBfPkSny65s4DP/t4uTpY/6Qj9XxBFshOuwlkeAXTm2PONE4AiydNPqBQz24A
+kOG5rE6yE580qdIhvK22ju5Yt+u4CnI9IuJy7tJ+SiboW1JUnIuUhaaK7skVJ7v
J5VhFFo+uUZ2sJ2rLibXHyDistiMGxSUjsGD/ZztfBDI3SraVQ/KXloJddr0m55R
hECF7N1rjDxZidHEy33CtG2e6A3PDVqBxnE/uFABSJE8F8pjI2a0W+iD7CSo7YQE
HEfNJtUkdqltiZAchtiNyrDUfAn6lfwU9DPoNEwrP6twi47UIy1LL73Ft3/uU6Fk
CNSvrFOWOwWSoY6deOAMa86jSy6zmY1Qd1OnKIvgVlGv0sz1Tb5RuNTfsLZPWN6q
jwAD7iXFS6bqp5CM/wdRGzvj698wtha2zvRWfPSfwKVubjuottsCth6HSRjJNwpm
O+hyFCcbquClmauf0LujK6WcvEOOQmQj5hF5iyxWz/44Uc2WMf3qaHFAkDJdEcbn
EC3NBkUP49Qzk0RADOGQFGZLiePqtcQfqzOVLhFoSjRyyKfGQ7tEaAug8JeD5LMX
4DsONYe82ze+zkiLrjmYfhqj9iiTXKmoo9c5K/H7R84wnBpbPQZsgm3yI7pH2OMZ
F73h21Y85WgBWpG4gBlFEqFRx84GEcPkxlRe6SYRx+bCwuU9n2gxRadBEHjJ5p2D
Cf/9+jUqKRzssZqS3eveCWFN8ah87KmVEcun482Es/LWqiaK2BCA8IRk9HJuzKyr
XpjM25D3OsRZHg3UcNy5xjqo6yD+iTAhNce4ctn+MCNlmZjQKglitN/kx2oCdRwY
6kZ0xEHdSjXJ91vpNjb6zrhPCDtW+wDqYzgDnWIAEidhM11cay5rBI6R0J+66Kq8
Mz+Pjuglu2jEUY6V31NBwqRaiTF1OqSjwUD+ad1PPtH9JpeyfuvxSjPJGZBDElJW
c6AC/7W7ZBelPLnyj5y+H0E/gnl3pYzI3grmDb99pK7AoTx9JN1lW11ipEiZJtt/
UhQBv/MKvES5hioIFb3muqAXF6gsp0yweHclKW8zCRcsH2yWvc+CM5+LqRD1LGtq
j8suRbksOtyMxMQ6Ha0+ZTJzh21YY3Ps8b7LEO+4U3SIPsNw8UOyJ+RWV/kcm82X
v6FuTb5H6BapIUnpgiRt2UQEAtMkiD8cDnwW2XnzKqoLumILbchCOIpCOGnj9IZJ
atzBrUExsEg20a4HaMefAdZTDs0/rsQwtucdTRIRDRYutbP0c/kUEvWULnVo/uSG
tRHjk+axhXYA9UDR3xLiSS+1JfKxQn5y/hFpc19QvXDja9YvSlCzuLOxdz8YUeYw
GAUyxkMZZ1ENrwGTIwCRRhZOOgZCxlVMWOAGgW62WFsV1ik5wehZoo8WfgflGRbe
eRwYb+qL446vANkG58c7jluPvNYCdooua3R2FN1htU+Ks84D5kIgBo8hYGKgfWR7
+r21v8WsX/QvoDUvCIGEWgv3ym7i1N8YhVCXLjTocaWolAAZsnaSrHJ3avQF+Tx+
96b5bodBjHozyavmieHFVWtk95xC8THSWlwZeoVWDYIjkee8JH0meEPdYC0z/uFV
3Pm5tZrDWSZ5N9kMuwPhMrLLbrH4P5MoVwHe19SoauDaL7TYT8Dc6cLYtDJjieJs
YCQgJW1lDbFnb1Xpyfr0zbfLt8cfx83DKu6QZSOHmq/kns33H9Dc0vt8pafXzP7v
rYE27KMnNPloKaWB7EKyQIJ1bNR1UFtKOrboiwXxBskrJ73MusX2fV8OQNfy9FyT
xdOz58FxWluFzB9tj4M/9XpG+zT2e4cKOJnlIA1gpA4VHxAp39RIz6rYbuz0q63W
PIPDpS0iRzxDv0+kqIOEsPZqnFBrvLOJCqgqW36+7DTvh+6sUht5FoRN6Sg+k0iB
TLNxlanNM1Fq94GZtfsAZJ6pi6socHSpaW0jbEaKHuJLgSn6qeYxW5dhN4qXkFmt
PRR6Y/pqheeWfR/eih2JE0gmfuNZj6SSbud2bfoHJiOpvuGCay23dfonLgZjnn4y
LTJJdORd6ZO6/qzi43gXda8sVYiOc41lqWuW4YCdsXk4XW5gRpr51UlLXzyfPQbU
0lZCbrzZpvTsWIlzGr6onH5ml9BjrNJCHv3wtxvWI4M7QmvrvWO0ub1gOg1vZ1Yz
1fWunWO0j46qfsKLPFDYhJvXkgOph8TGSvJHyT9q/MqK3Xa2OFyh5leKGVueAUSA
gARwX2ZbYzxOnCeCYspjru69LTcYz8sAryt2KZnsaMy1IDFt1oj3a29G+njgRYT4
2mEn01b1ltaIVcI6dDwCwLhXZcH7GwnfVLoQ1thzGc18mfO3qpSrpGvqQ2kbbNDd
OURVfewDP7f2mbwtxxndUSEBwI5mFsNNnpVUD/xXfwTR6pxPKGiCwoHQt6Ya/nyz
geCTLDDJwQikn2cV/rXL0pkdy+7CFqSGvV0OE8xziys7JI+ne4AdFOu5w6RdwJkK
fSpKpiZ3CMSPrBAssIudAZSPHB8+GDBgwy+2Y0DGhIsfsmefGijPjyUtOFNM09Ox
fSC0ZYCzao2ncOkCIFiXLG89dA6AAc+ETkVXkDhs/yp3RFoga8NJCqjnI7TgC/Tq
HS7/M8G6radBAvI5i7IqV1bNVw/p80mmi3upyeVL/yQb+W2tFi1caWrjoZNKdb8t
1zMRhUkKx1pka/ORdWiExlcOy2udPASb7FHiwtw1rgx6lf0uiRsBdvKFt2mwJ9Y/
7UB1hRM266VAwRImKRggfF3zifR7YabKUUtgaF0YlnX7Usptq3aCsty2GAGbUKnW
ByrBGREFdgjAAZfwgYsQtgThsaA/VomRx0/kkG5dkY1hLqLLHN4Rs8SL9YF1nAFX
6XgVbviol3nHjVaq2MzhYuHk5FMlA5k3dXHLPR36KQwSB7wUYi2TXLaBEOu1noPF
p7jebtxO2ThsdvYzBTtDkuXHCWUff2G1qaaKxbo6Y23LM4+A1FBtjheMjkDi3Njx
YLXv+IBOQiE+sCD46LBrPLO6szY8kWum8zbukI3KuFEl9pAfGTSWQzBUPUeJ7rce
XKKCtNKqPq4eU0hj84bHQ1Z6qY6O8iCRKtO5rI/yVJDfmyTQgafc633efYVFJVTx
ttO9yEdc2k80Ot5WV2Gm+3RAOgqev53sT3HD4ADuoae5X9ciOAUP8QUmuzppje2U
NrpSXG+Yik9lst7V05/MC5z/NFZThQQSwmVunikU69Fvj/TJGrUnGrGIY3OJaYDz
jJrqxKqc2VVGveXZZlRNE7hcXvg5mI8gCaMpkbYOLRBtfQPhZ5ufgSNp4MlxIUD+
7ZF/3yqb1QtYLf+3DqbtOG9FdbQPutan2axFZqAN2GSAszcgCnbG4JaVgh7Bqe1C
+A4On1jyako8HvnuS6lQWEoR6rmOyg7ODTBifDM//I1Ds/jlcjELJlA3NwcsFuVI
/bdCuYcfPTkuh47gqoBjA9o6Hd4oG9cPLQ/8z64nQghE9ZmsanDYLr5yiwNoPyCE
fPLhCKwu/n2Yf1b1YrvGQpIxaorzR+EwaR66KHc5ks7JZH3MTQp4uTzQfaqBJOm1
rM7ThsCAniNYzxjM6wr2bKr8r5pLeSD8hcHt2mIXztC6Zm/6ZH32YSwY+jLnupWM
N0Tdf0iP4z+NeoTiIUCXnpekr36kwgOEoZ4Kc71ogyeqxCRoxFsR7XYvBTvjJ9w3
ITsrGuI+wGM0TH782EbmWh/tYX/+sNJ9IOmzL6+6UkZjRUVlO+W0sVDroAll2vRX
bfMsn6zB5BV9i7v1xsCwsAipNvzO927AOAX0CeVwsgQmqClA9TbSiUo/nGK41KMS
vFRxLPOINjqhqzkZapx92KRc1r/FwbX8/c/j+W2iBYO7rooMPDTFIi4kgW74kxke
FOg8bS5vSraRKnLOlGAM3R1UXU2H/iJxOG2SkcgOBw8EAOT6uyPhlGx6rnrPHLnQ
oNTxs4kZ+YKlXiq2O+wL6Zn87gqkuKMDDyulLBBqmhS/7SBstmm4x+srKEH2ivfs
e7ECN3IDtepoasD4S/AKUKBQOgTwza0CCsJRrmRmBr3T5BWmRv8Uf7qwEsxN/H1L
hfifJqvW7wI6UXoNxBW08eCCsuaLz+omnsFsCJkYemxTdqnEVGAnjrIaQgjrS58g
z+iQ+uZBioOicrLmkbBKht+8hX10n6rEbF+VcEyohop6ZwLRIWwGB2k0RlOEtciA
zQExtKBYQQSAmtTdi4/jVJbWofdmd5bKte3km7MbTIPAbLEuX9BRYG6IQVfLCLNV
x/E4d3nX+iTII7wSUpwTonGWChdWNdHhESQAMthSDHr0V+OiePssdEwsgwckAlQC
Yrvvkwkc/MuHZBu9UPvlW8mNImUPhtI6LgyAOGIr+9UpOWCutvxVjdk2BlPZqlhh
iZgpwtfhzS1NMPXgpUxwIahmLeaTgVc0YCBBbdi7R2am4ZAKqFhVAOlWDVfkUKMM
K17oUxBF16ND6/NWxfzs08t/LZSv/uMFKfB+37/7VPP7DNp032Zw2snmtqzEoB4M
BeqtAGZ2KDpO6v4OY2RGb4U9a0hr33/Hi3QUmdIk/NF8Lo4UyfRki9xkOjQvoD/m
/bDeMNO4T095wUJT5P7QHSGiO2iEGN+LWPnS1qzZsF5xg+n3cJJuIzg3Q4YLTO/w
CnwM3+RlBtq38iFY32MtoAfv0d1CAyLx91GmXIypcI7M20r6S+wwAfxMfTClP/Vp
/LQYj3sfkUF9UbRLnExalfrxQyyr6vk0EUGNWu53a6sH+rPI30jxuB77hFRVxHjk
HvO2s3wDW8/5yWxsYAesbUfN3EEii7emDZ0EfRiTWvlgSYhu8yIkUia3xM2GIk1H
`pragma protect end_protected
