// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X1vR5r0VIydrIOyCoBCYqBWH9NMHWQ73q62FjiJ4AHMek5WMOXx9L3bB2YyKU/Cy
Mq90eFUSDuLxwIUiJ4N/TDSz/Qa0v/swFbwVDes03ib6VrCGsU0glaog6PJw/Hu8
qVAqB+6RuDkWwefpZ6VJDM6rZloodsRxIifDYPk6jr0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7136)
M463d0cMX3qfB+BEIOWMR1944fVRt8VUu75+f3gXKOTOsD/aXnssjpLmrreU9dfV
yWZpo0lZ7O+o/7EgBvcRxhOvcMBftnNZcCtS5fXkVs0e/seuU3nRsIkek7CN0NmB
jJvsfCxWlGx5j9cAk6VKLaxynAhOTyWs3KiEcx8CfCNJij/R7oEUdCcRZdveo87s
T7zLwPjdDc80Xie2AITCXXQiTek6V7Pwrexhc/sU2HdeOH4aJ7pzpP2C6yDnsiH9
cXQOEit4U8CNkNfFYH4dTZX11wN4D0NBbl+SUya4Zv3rKc6ozSFsbVMzqlgsQTu9
Ui7gJ3FH33RDtqwtaePL1M/RfVo8aochSHSKtLsR7qaJr6UNBjUofwGKwyO7Sf70
5HanXPgCiBLJWL3nYf1DPG9NFkeFK1Yr1BwtdYTkBscmqAe/Vbm13RlPK8cIX1Bd
lIQSYlVNLQJA9RTIY6ATUrr+5swh6XQOI8p4g1UTj/dLt4nl4s8E4mpECSQ4FsGg
wpKmyfp/oMgASG1akWAitprZPwfSHTA1aidC+FYRf8+yQ7uQGxc/OYLpPrW5Vd78
HoZXSVnBEPKg7c70vekS8V6d31+KQATEPVn9Vg5UMsrM77Qjw6PIxxdj5Sy8pO4P
yuKp2DUEs/KvkjVHrQl8JcVARFOd7XKApJEjFIL+xd3NYKEumdJeaHmGTCpnjGW+
vQoszGTeJW5nNJuTq7DnedckyHRGXyouYLJVgWm43YtD/JSw1cS83+rzogeqKwmU
hlQbDqUOryB3YFv6tbiNKupQ1aIYpZPDyGX/2wPsrk1CnWi90ceTDwkw9Hggw1OL
77ZkRf5LP1YKFL6XVqizqTFtcCf8AfdZjZa1zoXXPa23AWmcPV+beCiKaIXBsaED
WMSQJwLpwTp8u96awWlkXCLIbd7ee5VsI8vDSlBRD4QBjOLV1IZ+PpLZDYHi+HL3
+6pC3JsRxsd1tlGqpGmm/OFlMtkvHmksos/J/9BPMTSyMJfaR8X4OIlFlwGgg/0h
YUoZAwJ3486rfw/8r6V96CTLi7VX2btAy/bEmj5e7AUkyiGRIcmGNChcFlBD3uZ1
cmHiIWzTLMBqBAxhEBmJ+93OqC2MHUGQTiCVXroH4X9OLoI1u470D0u4VwDoek+3
yFqMrwhQGNGpvhoPVQFZGv8eqtbCyyU0x3fghcVRQ2vH+4Bd0VOOuNrCqgQ/pAQs
xwqMEwkoTueXpogn/PjFDxZC5KsG9JRiSmzfJ0yLHYXEOCAc0UbBN+lCkvFdQeW6
PY9veILo0YTFFcebBl1HgrcgOuufjnOtHi/7lKZ/sRiRVClBgXcOa4QF8OaVsAwh
YRaKYy7zAkDj+30sKRANIbo0Kap+qHgzwvclm1FsdK1BkuD1Utp9ShklHBnfc5gj
sc4ujR6I0AhCDLDSWhGZhk1QEYEqRpg2ji8o/HOlQoNt6R2fQmQxbauIjAxwq7eu
nxQ1RPh8HzDD+Lyd/Gf+PxMuTdgwss+qSMhd7x7SbvYp7sAYfb3GYYvBFrcELJ8g
Qi30yePW6naxeKfGoDo1A2bdfEXAtrRCMOKY5VBDG/gJSwxBNdKbvOK/moKbOVOd
JtpMciTfXZL3BmP/QzaIuBRJenNTGSRWJyI6m6fw1ez9+f7TwD+sW8/bBNV3HJCl
YXN6bFHPCSwNt47SmVolYXygGYnk+QFHC4HMsbPeEbBdaj9gC0c6FfM2xkMvYV44
IYPAqY5xvCOaeRyONsqjqHxyFEbIdsp/nt/Ac4fcRfoMQtGw+/WPgkI37EU7+C7Z
1LhQdX/JTl/txSdJqx3NNHF2Xll44j2WBB8gCQxbP7ifnb/nJJJhwtTB9N4qjAUh
gcPbT42ZoZr510IZBWLhhgTofnQLP4H6ZuwYfYl3vSnNTV69Ilni+tRTgPzk8AYY
ClF3k1Pli/Xxr35pO2mUTPEOMoENu0tc6JIffJMKDKKONXYqArCWMgilZHhrQxmc
kyq27QPLDU60sAJ/qkiXcfXvPDLLj1mOgTgLch0NeI2d8wWLcQNSLY/nKlqe6bbp
mJzHY1f6j24JbciNQFzsNcjoCaupeq7le89hHQZDML1b9nJuCbKFmuH2JroLw0yq
kcUfc4rYjjyPUs5CLfC2BOQrqxHcpha6lQYSIbPfuvVlHV0LOLTRpsJR7UliC8p8
DGkypLgFpfPX1RtOBsjd3FktA6FqX5PM+L4+yFfFcvr7MQgxmUYwjx6Kd3UGNDMA
+YjHQEz5H+rhqd14pyAcTk7dPkZ7sKADfQG1uVFJpb/ZT1wM2CiIabIarmJcR7HV
Ou9DKx3LAlQ4gIVGHH3a56t3wsLq8wwRlbm/n1HdKoKk5aDcmgYYSiUjiSLyYdr7
ufCDP+coCEZfk5eolfxuXZADtlSctCqNcJBK7IApsQrts5x9+d3yw2+PlekMmHlv
m7J1pkjoBBrLqy/IKHyu/pXO50nEEinHrxss/y1MHcY4TndxCnEgfc0/G4wlWCcZ
8plguPbaHDa+qYm2pEptmpL9MfELC+b6LI4EmqqttE2MKyYDAJ9jj7YWrzdsQzOP
VsALm9lREIk13yDtNidhH2N5/SV6VEsYQ3B0m+9qeEHVUdr2dDChUEdtvvqjKZ+V
FcnBtPWz9/HFjzZV7XZhG+4Yta3VQH2vHP2UVq0/yX+rGZc6CxMwBEM2g6BtYw+i
QCLP9LzaC39jnGrN1kRclrruWsuhNUcYuwCno/RyTQoCbkw7cx2NeMpSK9mLGK/G
BCjKvbA31rTBY3iQoLzDUYqCg/Y6/LZ+FWgm4neqSGKnkAy2niaLZ3TK9de+mxXX
aw5lEQk65EbttZu4yoohke+kLp0AdpONjtfhkau0AO6O0e58h0zK5odN6JHjEICh
Iyut1ttzNQQ/6ePW8lneH9E0XtzjiBd4Pul59cHhWnc1i2AGyhFG7Bptf/cuNy2X
H5e0MZ4lpSXaPbW703oUQkfIeanzK/MADQWqYMCnFa1h52y+F9O0KS8XSyTQBZhI
8dHqwvfcS4vN6jTktamYoT4NA1dZNNOPd9kbMLVtA7m5AVBBEYjfzbvK1HTsdTul
Ij/S9BY0Clljsjc3ZJayTPpHUV9665of3B0Cqt/fPY0Jvp0MjMX2dw9HUUf000Qp
mOW9Ue5eZXAzM05/ngNmUuwiQNiOvgnXbuje/J5Kz2rz25yFU9lM0oqaT3491yPW
nBuzx0GkSla2JbmU1qEA0vLVwb9qid5kLlTAVf0o+3uS2rTg72CEHVxE8Adlx6mW
h90Oxj40hxgS1/wKqnrLmJrCkoawzqTU42sZNmbZnayaN4RdGAr6KFqCycFtvVVj
bFdIz2YpxagxOV77Cq6rIbupDBlfMO/JHzJhYLPhY8W6uUGc12hJUTN3qZfNq1pk
TWyckyInnZyH1MniCJUdgCx/dA93lVxCFt6XqnYnk/jsXigj7wSQ7XyZIH3tOFAY
bK0hwa4TbLvf8kLiZf/b7quRiobCoEbfUA1ofL0zfQVIwYa30yF+XtunN4nScj26
VESrdU+jJzeK85rJmL6eVXfG0X23DOrvh6Gfjsm1newfHLM0RUzOoOGnw/XKf1fk
oiHUu/+eay3R8xEC2v/wIzO+EQK2DsgYPwbdOjOySVqMcVmSXo3BnFCd8BMn9huL
65/HdUMs74uR77eOTtI9QoP+l1YX6AJCeIZ6SAF5vAefUa0zahC1JN7SfcZZ+DrJ
/LOi4OVVliNJmROzgk5fQkGm2mQKYssS8lk/J6U2hVvLtiASykPTPtAc0Fj28LVz
SNBbB1JfGoEjOY4+VUtV1FraR71TbQGQhhSqheeb9AkARiuEci2Uiu5r0/xazV0y
XcJxpYAX6+0Gtxj72bMvTgO94eGmFQkcYUoOek5kTvvMoMqFrJ4XHxGpCzk8ahfT
tWau5dngDjWR2nMBZbKoAGRaEhKy8jm1oAIJrLs4GCGcD37K8tWjQ/J+IxltKffl
pw9/uL1Ll3lpscJZYEz1wceOQm5LgwfxNWp4/Tea0yQjHMINUrwAvVs7ZhqVH/PK
H4V0Mrdp2At6NV6NSRYK8EgjAlc22qsLyYq/lR3FlxPkrJJlOu2WOJ6OIBBO1ZKW
H8J9CGML6l/n7fr3ZnQY4JDNn3Ba7CJu3dxQcut8+YV8EBj+sgJVtUfHYQ7YTbfj
b/iYlsmNliZ196pPGCLojssjO1EX3fjnxNOKSLKDSHHhRAjQktd1KssZfeZAM9YA
AuqnPbjKXp8hWmA2nFuxJaYXLeM5wfODknfvrv2K0zsnF+taYOT97ZK43362M3r+
A1nub0jmkAix6SgWBCq8NibKeTeVn9Rt/Yb0sfhplHTjyg/a2D56DSPfABq+DMHc
5buWfExDCLr0ATqKVI1OcJ1n2gY4W+i7N205aaJiJyXUnVsA29jRis4WlqkqWVQD
iW2P7H6XN21tz/gw48jVNvgruvjtwlzHdeisZd3noNGP61di3tt8EijEZcRwx2Zv
xityXOmBVHwYbuFk3VLjHti4rb1GhIFuEWrhU6OVS6A3gvpBPXI1QU3z39cqHmlj
XneOhorSQN0s+nLmkIkpwYu27Rtamsfn1SwdRgFhiwrmQ2lREI4x7Jg8Ld66seop
q2u+BdE2jqPS3LQvFzcTYQkc5664hZtFfJUsOzdiCWExeylXVAn4fLldHEERLhLx
TMuu7RWCtuM4Q+P5tAZxlLpsEjVxxRgzuTP/w+voWsfG9vH4pIDN1aUzkf8E+PCH
I09wVCNGMPQe/YgRPMmAn9P4vr0ywpnJKRmrvNYtupGQbTQXOy2OJb/Od0lVN18/
f+Ho1ra6DWmyfzhsScYUfjXjoALDzkYUUGK+cJoAWeSsdCH17Uew0Cc9fsfvSwOI
jSzb2vmHrnSqsvFOT0W9gXAl/3/eL2SM1eH4NyeNgmCOYjO/I7xcv6X5kmu+dbTg
dPGeKOdzXA8nmJJmKzGwRop32aeFVxSD9kLg7m8BFOX/nCjxXY3xEX6xx7NdTJWq
95bDzs0O+CKEq1jmvWCduo7wHfZmkz+F/akB3K+dvU4bTvFQq7F/+I/r7x2Jqtj+
EWcKWwCmjiio3WWFqCcyuUgjSu6y10p4+qMlHkMVulr09dgo8tfx6mL3O5hW3LkB
g4E0guSzvwbQczmHx6YTIh9eVMylcdCnM2g9xNLcR+mp1URO02sPN08I5FLvHrdJ
xDPJJ548TcdcvU4c6W+QhN7mrLh/AEXdIpqgp7LU55bBcmJzQ+qjcvnWDY1c0drz
KXxsGDSqKRAFIrgekm2fpydXRkVJoJ1Ziz52WTO6SSpi/j/ZOUTlUh+Q+kHSmj0y
J+/NvZiuqmKvoy+qCoCV9HitluNKNPBJ9KVr7El2a85jgWMBq1TGepdvTZup+YTT
vC9n8s1iLLrAjZa5ppQxLO0QZQZ8K2DoJww48K42rygx+kSxSObZ4BvOURx4INJ/
qAkoIU/h7AUFcU1c+sABWbad01S3haKVBxzB2m40yu3pWub/LJwnQtBGmKeDBXhM
z0zdMJXXv434WScredxq+TgeCEl588z7kug5c/5uoW+D2qPNaWg9/tq/W4DmBzZS
tyRX5BHSDU9CkKlMKtADzEEnIe67YbxjF8A4oYN2HNEdLsX9ZUs0f8nIulTm8gQQ
3TxeqWrM1XipnnnkHOmjJ+VriF8VER3gpXfIl6sbiP5fOGqAzhFAYbT19lQZE7Mw
zdsXG/wGlJmNoMpwssNXEtObvsvWZx/5V4YmsX/zZVBQ3iBLGWWMQtq9bLG+ib5u
zuj1DtaD8Xx9a15ZdyYLchmw5T1t2LAbUFcu9Jwwakln0hykpohghuk4w+tYsIaj
LG1qwhylAPXlTc1yeiJFUnpEGcvVbiD2fr9SzMhvQJTShQ3C5KB7FZ4CyxEnMHhg
D3pwMCerRqp4ZVP14a1pp1qWNerRyh9kNYIpXsBCo9hlzMIiNcqNQ+9FWnzShS8H
+dGUE2knllxkG7HkogN+dooZxZqhFxIfTI67M+WTfYHdk4L65qxTZ02sjkyDLPpm
cmEQeGTk8bfsPU79Zyyn91CQbR9ElRsq2FUxnm8S+pUOt67/H/sZqkeccAmZ6HBZ
OCj6nBO5S+sitlSV7pfVE2dcrqKM1WySZj7tJ6ds20wIyRtu7uBoNI3K4k19faAK
09AWb9rzIwx/gU8LuyiEdLSBaTK+JuY2cHmonecXi55F8GpC/5tFmNKVvVfe9BjZ
q6qRwHgMjwoAArhBzErVdHgNAxZeZMagGd52o4JF4estJg9+4mMoqdmbGQwgUrYk
9iV+3E/CCA6zctiM0OEsGP0LnO/reBt3EfrQkfac8SSgKMekWvgjIwfgu0LDP4Nw
JIIq/Lk+hk5LNW5vB8rOHUJ21bDUsTypQoCcsH5ju0j0mV3tP1pt7ntioGWA0tGK
qNadNF4lxOKtJ9bWAhFk5qZ4egz99r0iWr+HsAxmiQTv/ed5gyPAInbzGkH3jqrm
M7vR17yqcH6fhyPfN1qxSTc2gQkKfctazRh6sNZozU2LLbxcWx19RH1FlzbdUwDw
mfsi6A6E57PKBbCIURp7epIeSUGvOnDNk2dZabE5fczHn9D69QjAf6+H3kWnO2Hi
JEAudDn3zFPiyq+UZMKWzsGlKzhp9XUC/4lCSkqvWFzoEU50jrZ7BGu33KRQZYWK
5T0yMta86buDBlWosuesCOQUlWUmiTwPZRtgYh3yEiUwqXe4DF7UhP36s2V973UN
VPfHHuA8yw1jeC8h47zku1PLl2xuerbBr2giN1TLe7Zxjj/quXnv8LAWCR6fciMi
9B26e8KO2q8/kiyRdED/O7l0HTg3FF11iO5ephY2U1fFut336cqJxyBog9/qy/wl
WaaNls7Ip0tpvCD4TD6NGKtIlPJdtHem/oYysBUOTwA4NBs7Kon38vRV8Q9Zg0t3
mTSwCNOPq3/8Rshvpst3dSETBxn6abQBUmP5O4AA5vPrluQzEWVDtTqS8NzQ818K
Ags24ZvBG+jj/6a6l+J+3qRM8LB/yJ8fl8RYOk/XptHEgdsCf/ILdwxtu1CS/e29
5a+vXW4fBUPctAmzBGIJIcf+sci3/j794yH60kXzAZ5aysM55pu8hsWKJo7dCzw4
RsVpBz0WJhA4OgHzZ/SHh98vBveDY3W3tMxGhnGG3SWHQc/WkmoFT3wkux3LWCrN
rf8GK3UmGJfSXTROoNGKnJrRbUO4RcB8MEm8AFKYprDxCWEtfMPpHsEk3ANo99GC
E5NJrN/hcjUvD2XEydUHn7ODgu+T55EP/VZn4vCUGmPdVpGpnq6Uju/JC6SEfv+I
0ppJjnSmqkVk2YMHKfeMm+CLZHaheYdVzkuVujq+Wq66aZ+AB5348rD7tlTMG6v1
HJL2ORJncuv9MyZkmEyzL9mH5YVxS71QyAOSBeDUWQ1knLUfJISKsnHOMARvflE9
GiPuE0Qo/RGcvyWYUCxnrFVQqyKPxiBOYggqD6hAMHOZaZqIQDjLbt8jhSPJ4eP6
IwhMOtw1AX0F3xOheSMmncFHxLDQN7dzSnrSN7thikiqVW9qX2CkntmsDVWqELNO
9UDhaCAQWG/vWkRxpVQ/vl9Ou72X46Ic2m9soiY+kUHEU3vblbzACXi4FrwXzGUW
qtXV7BYhLUy20h+PX8AwhK89GuUxu46N0/nhPsZsey6h/ZH0MRpqLFsogIUWxKiB
GQ372luBtqC+5Q1U5We6ZGRVvtdb42a4M+JWMPHRKl9bhJ+EPe1dhSke0LIEACpx
H9r7Raaviw2DgtXobKpm9HI4sncf/nbXedPSKYu+mKUEVCJVFnMERLVbUelvWySg
FTEgOwZka0/Jt1Wgh+NflmmC2QAfI6WoabPS6U6HzzoDK785BKRwTfPY7jc/pFfv
uW1tSiR9462nq/NXYY0qgNY35arPFMPSLNw4kxJVsvnrvIkJ8xlfngk9B9hYR1oV
IANyJ5TnvSn6mWYgc6fwM7Oie3bdWYAX6XjRW64/9h8MwUk3+B0B4fD68447EJGK
SGkBu+rrasSN2wVWMl4ne2FxvG5I27krfpC179ZVRUvJg0tR3A7vPkks2uNx+oXP
q4NRrrej+0KhvfT8XnF68S30orZGLSApGp1CRrZvC8li1c7o4mywe4KlM+JPZaHv
u9fejKOEvzLSlzPEGKn8A27ZbeuNHhQTIAW4TMiAN+piCDRwd/Z4hN+3xr1xa7x2
JCC5eDGKn8+b1fyBGUR+V8MZtnYGAzcVUG2ZXIM6SQcPuApC/n9XkK6B9W7WtYJw
AIN5eI/fG2RROO85FPNATCAgNNgNEOlYokBnlfgEBhSxMtXdQYFuFnXuXduZEfkl
y4ZxGHjJdU+6haFfl8GmPYtQM/VY7MAB15HQkafhkgHfl+NT0xxlVy93bB7379l6
AkB+BIKtNaNJigfzH8W/+ma1UkM23zf/BvuO3a/j/PUd02TLSEalgJ2XfsrBAEyU
ouqpbYw6PABwYrsMrBELnNnbaaCB/I57J7wx9ovoPPU3u2A/EBkduecw1QVvyrHI
4oxgQIv1CdpUOXNA174T/JcomWV9ceI2jSWB6ZX6azCHCfdbOPjkt4PkZ/CVhgdE
77LMiTDO6NVb6lcOTWTtskvnZIsCduUaWqP9XWqt7kF/vpfjPrcQQHDrfBpuMQLz
/k0ifalb9hPwEIhXjmBwwNoWszg7xHragPsAwqJkPnnYfWuuTs8d0DwRT1y1zE1t
SGW87qc6JVOQDQmyEktJ/G1A4Wgr1wEgveFUmwtGOYZbPZl/qLoqdIBSHmL6e9Nu
o4BBBady6HfpGvrXPZutdTwMELn3Y0OHKLpRvCGpPRQVkqJDv+j9ppfkX4mZ6+VD
q36x1+PKL4Lz6oMnm2ahd9nYjdhzU63OkxZgmMMuotqnhMxXUUBFV9/SnJ2d1+zb
0KjFUIwAJNrELDgUJrZqW0uDkIHrnALiRlh2JUXTS63mpyJZ1+YUxakfgOpjXmYi
A0XQvD/KCyztr6Be75hqzAp1rQZKgevbrjtLL+3eU7o2LU1Xd3ZLClcu4VzmMRKC
kfyAwqzpXwE3R7CKyOziXmprhgqpIaWLtPemLBg2GO9sfA8T+DwLndRPpq6nJtyD
iIzRsGWbh89lAriKezFiQqxe0SjtLcSIR41Eod183pdj5sfRf6mHiREdu2CiJxtr
VB8LIBSlCGeRSP1OWgVT5knbqYGXlkvEPoKRUia+zwhKVgot5CbHAcq8qnN+bcW6
HAURJGtwnwnGLUW4TASniKYkakTTJ+/h17V0E4pJlBtovox3q3pQSiXKa5zUq+of
WWIEqSOoZz1ojGad+ApVG/oKMMmaxx5I6YzGZ3VrpEsOeZApvRNT9CnLBbJFDhAY
lJXlZQuB6K5LVym5m5ph/08ZG17iEPCQ9MrbJyvsLPNcCztMVisXTtxVI/tXfRrm
hpZaCVe4CxPhnFciQTbhxyuFI2htnH1I4QZz6PMcuNQ6xGDr2lKgTQ8cYgWc7nDV
BTFCjSXb1msMFB/HYVKBb7lquPmGEhcvEg19qGOQXTU=
`pragma protect end_protected
