// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SfZ4/UJTHUhAnhGdGgQcvhhVd5BLhCqSNuBFC4f1Ox+F/wrWAA/UHwzlHNew3rj6
Z7P28Nmntd5UWUPZR2qJclKdskKSewFilAlklAHlo8bDxp3SLBH/807rPl7YBC0Z
kepfiXZ1bFTlNgcRFdPl1FjRWLraAQbdjVBpXLOE8pA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43264)
EPaeY651vnIFBMkcQssMXTzm6UIg9ErgRh5W8cJ/hop1B7FyUFWSzm4YSUrrXGKO
TDxznZBdEcpPf1BwPALIuiS0SqQIXpzzHb9dYyGjHolXJ7lZ/GNw5zFIbanmIoDr
5lGMQHep6LY8pkYgNdYsDBXjX+Nx+WYaziVGxqa70DfwYOrW3DI3UUhYOO6px7zl
cQ1wQ8XGVi5E92uMlHdkE41vs/4rwc73SFyXTLWT7EFlTstSClVWrkgmwSCkO/fH
Q0CfrQ1UMifrP4XPbESB93bTNXoZzG1ULt8bXa5ZJOIBVkr6NBuM0dc9t3HAyZ8R
k8rBnJ7Xn7T10JpQJY+vxYHpKDHMnWt5iI2HzZQY8CdshaIfZaeX8m6FBbqtYSep
SioATAatR4+4iPArBBy1pvut0GtGXssqKLss9OJQOcDnin4m/A+py/oNnMv+heKt
iZ40zDBvsQud5yvSIRIYejj1AOdhY4L4veh/crDky1x2cF27Zw/qyAQ2j+6wVh+j
5PUU1roYsF6FowubwHHUMaW838oOIhVg/6QPcpDpu+ceyGxZPLZ9VhEhOeaVM6Gs
JtMirXI7GBEla5bs4v+CYCjynrjJnus4WqpYdq1y3Ni8NtkWZNHB0UVAG5tYYHB9
V4jMAqbuJ3U9z5t736EwNXMIdL8siutgmN70CRMUWD1iKyl96v25BExyAgpDrU/h
VoF7qhw/6VRJ+opnYABlww6V6Uw66MNG3N2v+PSwpgcOk7g5kRP0xuKAqM1O3Qci
AQeISoZOHsyceN+ryJnZbrlvmNDqEGOcJ28nsOVkSZoWG7ZfQoe+7VSzsDnfZYER
QP0yKOllcuv9NNGXHovDRhUBMPn3VvUrDnlXvra8TZ7SqtA5Df8IIKACGvzL5QH9
anz68p45ecwZH3nLNQct/s2CsxKNxg2sbO+nriUfBn4m6rLegk6h3/cmUG5ZR+Qz
8qZy9gXd+cntmsxZaSZgAH0gWyfLUSEt+8r9XKHF8AuCEAo9QXXgn5N5Jda3NjpT
grVohrZGxzRtyrWDpce0I6WDD37egYk//iymtZRB0ELTVIeoVyrHdiId+tcJBmkY
NM2pPAR0omTLzp0LQ1HD2if7MpYlpad6GQBJR+mrImFuzc7kDfj7H1F8EXj+966N
RS+R2jEHoHivCfedccTUBExy0UetP3jMXUqjRSa0kZxwXOTGyUbbzvLA2m4rHeFU
8GljLNwESYKixRMNINhY9tspQFRCyNIeGNbkjkinA7OCzzSakLd4VaWfH/b8O2+K
/xtCFd8RwMfDQlCBOXtV1WNhkg83g/dMglOTXxVK8F8zi1HSBgb2klXL05xfLJ1Z
Ga34CmqxHiV0OQM1aHxeO++CyS+2gX1Nm4eTg6BwGnkbYkNwb1BlXKJi9sk5Yl+J
Il4OZxF0yWFYhvGHSElMN2UrDm+bOhncPbRdgddLDSCbvp+U2hgmBOwhYl25Stfo
IvqxVpW7puXxXhNU2kaSPOe+U7ZWG/lvZCGeXVsvVF8Lwe73rt+To55ruFan/TrZ
mhX0f/p7EkC/jTnJoiExoXktl5iVXO0ILIUJMj+DF2qjKTsWbiS4qFRvvuO5SlYt
pTwf0iuYR/QX5FYRrVtN05Yx73bNhULMlhSLC23oGRA92bkWL+7vT6YVKU8cviVG
7bKy0psXfDBKMkzmN0jE75pvhRtZ/y30i/A02znB8UrOT6cEjI1nl5xrupyO/EQr
eA2RB8MWlhvF2liIx00NsfeMYjzK3pOQTVcxqW7JhdQOcjxzhaR2Lk3Mq2GhD7Pa
7AhQKSPs64GKvFYVNziw3FC2BpbIczIIebgimJPgptgeCfJ93M3mX9coBbhqkOnt
TgZGUIq5YrCG324qNLra4nocDbIK++IdZaNJsQHGXMWLG3vFTAptNz0dVKPFmudl
eCAk9gIwC62cJBZDzMFMTm0nfMbBBhw1PJQZFNZC3ybdF+woZwePrSfWE5dc7SeH
QxSk9dQ2Qb9P0jTAvcJ3oR95prjFldH4iShGBKgSQ/Svs7A+w8YPXnfXaXTFtWHd
Xad454qsqkFyDZaT9jwjo82cSQUnSG/fgLnEm8C1Kag2bBw2Y+t3OgO1XdTewvra
+o0Msl6DOxoHMD9yRirqaRvSoyeZPOnN/G5YMvS8eW2jL7l94YMvQ2FmNz78kAOI
Ia//fgIy/TWu+Dkbedk3UyXxSXFp0nQnSO6uVHWM2p4rV3C3YF3Ktpepa52f/feG
BVEfwVddK+Y9rRpFXNfZhxQmIxtVjqo6X/AKzcKadbyzwbgEwOrVjb9JUO8xLxAT
VpPS2rKRJwUNSaNg13rR2/GwjHztdmDFtwbRetiWbDYFOFVS0HQEdcFktzNLaoCW
FEy6W/dF6E8gy1Tv6arzrkw8DxelOP2K4/VuKZgsesKPsoBW51VCmp6NH5X2JzEo
dwXKEEK+V1cKK3xvChb8oi8/HNAnFdEjZ3qdfEZZfXBGFeJFZMkq3c1KVLvfwB7h
JZ/cAwFZSiS5ARmw3e4kXSwUVPL2rQ+JuX2Wk+ooGA4HloFPwDm9ojUjNIk2ePBn
d7CNhzQqv/t5PN0VsVbBxKvIBbjRSPUMCMKyV3EnkdvYA0O/Mbg1SokLLk0tjAQB
38XVxDhPkTMocKxqe4QFroLVYW7acqUZCDSVq+UF5R82mvoArY01wp6QuTdbF2nz
B6NENrXmFGX8FEjWkUNiULo/Sr2H1VB76ds1UOTqOq76/CHOJZlUZnpRPg05g9ms
IEkNIBijzR/aFR+yJCGXL41SPFX13v151t35YjlPiWJPhTK1gIn1ihhgTwqUwzG1
FYFT6x5rZg4yFZKo2N05v2k+2pagHfXWKB9fX40xKoC7RphdXXxRRPCyDkH3WYAH
Ip7DjV3zu6navKD9gnnyKJQMQ7KGo1tz6ksyDKrkEKe6q4wGHvV+YJdFA/PvTSHP
eElCSPgj3m4wvrWK1uWM4Wu4LAJSUhUwP+324yaFvWGmcWgj+m5Nk5xFDGsK4T59
Rb4LFzYl8yOj3eV1FbFvjgMRvasVRB0msgMAcEr2S9X4gKi+7Pp/hcg/Og1Bn6ET
wwoONSxRN59gN4D/BZAz9evlhfvR4ZxeuLEQXD8Lw8hfJLZJu/kpmemt6o9CLOrd
PAVgs7Hped8AowZ6MdjQH4ZrnXB8VGCHmFiQetsFHOlkLteL8HYHrFsWyWA3Aieg
yms0fSRM1VSb7FsFmyrvU2NJokFaINnJBZ8HEzTNZ1jmfWlwYl0ahzzZfuksnUTM
IGKYvhMfdmILvrb4jNTM8rH+640xRsog6FByQqSb+uliQQeGZhiUJt60msn3mQs3
y2tkQaZEb1dmmKqbHSOgr95YodPSdCqLKYXOfRNwyQ3238x1H+vR7Dq0iX5eSvPC
wXcwCqu9atbjMhc2EdFCabj5QuB3QgV4ewKCC2FCEZnXttxeR4SC2HdLXeOyW063
IzVZyhn+4H16/KvHI/qJgE41l75QFnPWm+cGVB9Knlp/Ylme1qs2ka52aSSJIiQy
Xi5FY/Tc2QdKeOvhNTk6sCvFRupDqzJ6R8cPK+aF1MfjWya0Yue7BypNW/qn/9O+
oGuaVJLgnuSL3OiAozEpYAGspra2AV/5cW0adgHp7RpHeUP9tMBvBNXfAug4EhCm
wjyIL+VexIPHa/z4E0DLhWbTB+ReHKeh0B+5cdF3nVTPXpGIQRYQhn5flixeC6WG
4zDa2KvfUJuCDYgNIRE1Bmifv85jqAExOeBNsDN8xTyTGOVtdk2rms8zaHUodOxf
lpRUwSf3025v0pPbNLfvWJ6Oqq/+GX9AdtYK+N+JMahRoGU+NPRkXwAdN6rdK5ls
mmSaO2L80R11+/zSSpU6+OWN4ophaMWLT5BzIf2qUP0LTcxxYPiHamYCKmyan5IO
xHtq6iaNwYyrRQaouJQiPdoT5eN8ab+WGzrxL55qmFVWDtwKjeTS/f8TZtQzGF2v
EW+N6WIB9Hpw5cw8UVc2eTEphh73qkzQKJTLQQyM3MZjkHgCieM2LyoUBl8+o/X6
OLA/eAtGyuyehS6m7FTLLFVCGTcewWWLrysXixJtVqiIFa3NEWwFwWUYJP9OxVTX
EZVbqI0J3c/eKNXZG5C1PgQ5V2T/UI6BtCVI3FsRaGK5jB8ppuyOK4gBhgtXGCGd
xxbQ3YLHF/cjqPQgfpchrvS8L+l6iIZ23b8R+hxjTTgr+yc6wMTPrU57a44QUJXl
vik1l3AP9wpqrQ+SyuRAhRZzjqUBbTPuuenJt1UV60qOyLmce5SyBANr0HI0nQ+S
fqB1blKwAW3uWC+ZiZqAppHSQ4Tg2edqjvTTL8Hv83+4KE+AN4L6osqiMg2Bi8IT
4cHIRq7nKXzExb+gMz0B8px6xvbxfMDhEzpuXofq/x+W8P2KUSLQFEUARBm7T5Dw
E0ol+tqzkv8q7NYomAtGDYuPC0jzHDuVl5vBKJ0t3BON98Y7TZvIkaL9EjwzIScr
f91QdI4vxe8dUEpc/twqV0KHqocVpsWbbdAWKGkk3tb657pkfgVSG3v409M06bsv
0bMk4thXC999cm6zPbp1+zZkzYQf+DHRGPHj2nXInmi0M1qTKfOpAc4X+TfXVC95
GzKu/BDQr1i8VcPLdfe9XUSql45j01ppIKavxCJPmRQWNpiDx2g8N4OubwF8neHP
aOjoGTEqTaGsBIsrvujI/kXIFw2K852KtlfNsTHtY9jUhfsQvMIr/lHq3vYMDzoG
i3JG8L6m/EP0N8SFpwLeX4O9VZO+cc15HbE4qq91wxNIgT8rNsEXcW0VK+5H/i1p
KVJ30Bkh14vNS1JLu7A7K4tS36ZCJRA9nAkKoevHLvclfwN256a13x9c9p85nLdH
aMzf7nFkaaE68g1FhK2YSG+nmlPUP9ZXE8izBA9PsraWTtFJ69ieZhSKKnskFAqx
oveJuTPoOn4tWAniDyr9+9uPxIdQMtuzw9HAa7yr86UrbNZqznZiXyyYcFJM7dQ7
Vv6sYjbkW19Tq7izkjB4ZwsOGN0Xno2NLqquHZxSvBftosynd1aWBUguANKNN5Zl
AMmcDdAuP931pkyfyYCuPUTZtcwHJjyxTl36EYFS20ARlEufW+mTJ7+1H76g6JiN
+07zptuNmkFsQ5GQjml/AyP9vCwqlZPq5kKrW8yqE8lbKtHUnrkRpqkKFK3XJGnY
3RvHE4+1EauPLOZ5Y0f4chfxdQXyh2dIHPkJPcEtALqCD7NcG9E+Ef3RhUkySrzX
beLz5dA5nYofByc/2c318B86sEF/6GbFxd832JaqJn6KbuKUen0Qq3bSRajwy+Zi
I+APgHEpw2yUZSss8EWxvOBc3dqrwDVQ5TNwprn3cYG1jpBUHTTFU3W/JHXUls+F
q8SjKAodS9D/ra50no6ObSttZbjf+uklqbTHKHrzxmRibIq6wLsg95MxOgbiwxCr
EMj9/3JsnnTMMRpuv6zsYbVIQ//9HB1R7Wo/XJoLCiVY4D4vpn+1pFJZgH+VqG8T
mDK6l4CVzHaHfm+vT31e4rirrAwRhfv57zJpn/ESmVR57cscadR0QvyP5fr12y6Q
tefhwR3zF3V/Ntg6wSBX9sP3mP4dw3gsrFyxYEGpT7Sp1OkD6UsWDFxXF1cCfxtJ
775LnB34hSyQplCTdA4TiPlZw3GBFKUB1FV+gGDNhvwkaQyu6jAGm/OEiXruevCH
MuZOk3+VCq9Lm6LRgOfoyQPDHdGtBxM9Rxd19tYRxuJ3GVB+oylehJQ9vC0R/Ivl
c3oqpjrMgKAk40mA3YYW4thApZ/UjvZ1OdKHAbIzP5PVXERrw9iRm3zubqTxYQnb
aypn1V6QuceUW/FnnVefZ8cCjmEkknAjeU/SA26yiQS23UTjkde2FkPW2OgQ7TCK
phZ3S0rpA8j6O5Qm5A65Kx1VC2GfWkPtkQCEYyUmerO4GgBCyewAndTyh/Rt8wMk
bnHVILYjgdB8iMxsu/ajzqKFnLM34ubhXot9NaXI+zQZt5Ucllf50mpUHgMMJgqs
ehz34RBEb511cvI14rR36TbQV4tIonRCblm/6b+do13csRHF4mz12pdDWW6pO/nf
idG7eoZqY8z0wrOcL/Xa8sEPIlJT9K+tVLc70S3DkZgugGoHOIPXJRmZlc2bJLC3
VaMM1w19upm6vhQiUuLofjzFP2Yb19r5PcjGfGivGgiFhQuBTAHG3O2Jl3bgkfcr
MPbsJsDczu2AZxseYlWQ09yaMfKMdP76hEuDmNPWPQihW/Z5d3wBWRwQL/p070n3
uZPwhqnfn1ddpUJYB+wkip0Yc9gqRodu/zH5F7MImbkRc4yr1hfIDU+iuEg35n18
nOtk5Wt3wbAlzCMfvggrzTiaUzV8FVJrirYRjI37nT0Ogs5J5x9P20k7QTwWCt69
EmRPf5IATs0w95v3uYB1Bqwml7tNDm+4r5XAoMRcADBN1mctuot0Arknnzw2OHOF
PgVVQcw9JwhA+HhX5BVyYCz6Z8fbHjKP+DwVmTW0uN4uhPYHBKYeQ9Dd+RUmXwfx
SYDBYOxW3cIam9dcESo5ER/4lXXasQsZR30hClXVR2G4T78GMulstdo768oEJ83+
M8bDsHvn2REGXE7dEdfRQnj+r7SGA2AGpzjbnX6bJktMYaHEroLxrSb+k+UR8ORY
ZTBNcflGmn3RwHm1Khb1bVhLiUmFIcdPFZoqPQI7sq33+jl2/4zr1vczc87ATOz8
GHN3Thimww9DoxL5+8S5DXqmwCmhSIhIOWamX5RzssZGg6tvvdbem0Dk9y/UPqJG
qLtrByvPk487A7sfh9Rcc1tDHDKf1htp9wNbcxlfUyKuDAU7xJ3HehInaddfTt9D
9bGftPk/1wpPfTdzn7vybwOpAYUJ7elGRj/kh+YUlJG8/BTjoA9YJSE75N44E0/F
tJDx3R6aWBKE9s61dY5WB+MQR/ZRv5PodjTg382c4tydB7cO6HgMDC5N+zuRJEZl
KCGwKGvDix5e/l+q8BU7cK2m/alTBwoDmepgRKwas6U6QFvIs1yvzJTbCV827u9h
yKVVkcUKKZJOrKIlLtTShMWcO8kO910hpqXXHKoXCUb0uOuJwfX82KBGsQSPMH5k
rqxbKe1Kmhmac9K/c/0Hid6wJzwReIRqfYYB3U1TUvlJtUrxGZAwmZDBwMBJtbBT
odeb1cKNjvtI4Tp3uOyOv5xSJ/nFNEviQkmhwuD8oU6bsYGb9aHYnUpFCAZNj3vv
mpVuorY6GBA6DRz5yawLM2OOFyRHtYzQFbE72a59UZZkqB4LlonVtrdvEjO2cAHa
RoCAnok3PivimaArA1wnPpT0i0cgYXCRyrAaRa542YQNYshKvBcPzVnxDqQRcwO6
TX1kA7Huyllbt3RYJjdTNlPeabUEfIaSVrx5MtkEc5Ch0tAmlEn1EFlqG7q8drHU
j+OJ0Vz+pjwY6hIYcW2psKlrGPRYs2ZA3g4oZOJ+DbYPmYHfkSoS4wT9boY7aMtp
KASrRzw8KopsvCsjuQ3cAsHkGrTRcUZieq2ZbdXtHLIRzbZyV6gkbu095bH0onm0
5rlR5XRqfhFdOVeAKVKfaK6xyea1wJkjURHRVLHSXaP4xFyNWwRHzlNiSxIQ4cX8
LKkMpiJu2vsVM/N2rVhuNxgo5R2Awhckm1ceUX6+c/tOl6/ODMcuwBCimgADhg/N
WP4QzDpgZtuc0Vu1tHtofswiw0OpViu2KDiUzm3mLhOG3xDd9G0yslfCjSlgYHVK
DiAq556Jsu7sr340HHe0zT6icJbytXRVU1pVJvYYxhWSnN82D/XEQixPqpSRch/0
Dfpfky9bCb383VZf4Lf0v8rkeaGjp3dUOpQc8TE6ojlrPr+kV33LfRJMbdmlhO2T
kHGAKAleuECN40hb8eNh4ALHN80GUjmc3SUnrZzpqkRiJfFnfc6YG3Z65po7DUa+
Uvj3sPE11bE9eeUHAF+3hOU16z8LhxFiw6ql7SO+dijcmBOs2+OzL/6Y3UCCALIC
qWJECrJ6TcD7+Ga4SHEOMXojnNiK5CmJhNkmWsfzL0CtYQANiVxziEFuZWJhLooC
8frYeKou2Q4JJcsm6zbcCS3ohdbHzaa/+NC2QsaDzwfX7Hycpk7srC7nQYVesTDH
KlLSVLPHg0V4ox0KUEYRpJzuMxaA9zN4M7cqFCbpRg68cN2pXAdoF3NT2MEo2Xv+
bTFItOKp/SYoqPolmUjeigLR91gi0NvcLoJdWJN4xEkUHs68eDHemClzriCB0CtR
2ncw/kOZVcSk0r29cE+Vo38GAyZ+GApb+1RVKEjmLxNVddl6ldL7SmdeE70YC5jZ
sTD4EX3CpLS7Hacid2DD+CWWuGKvDXr5GE8q0UBqVLG3Y4PSWz6K7eQJOgnvglO3
8dJF+PY3HAlM+4Sk6fM5E6Xw/tL/z05emWDbJ1b0W0AasoREm5Hz00MkdhwDieoV
B/tJ46Y3FfCnVIPek7IPOf3SLcVcymHEBgCEBnbznPDiJ4M0WLWxHE/9EAqfAm0k
XsgCGuKS0OxyC36M6rJdgZr3k8y3BUyNbDvBy7lbffquSQQDdKmmcGAIbB44NVlE
KJHr0aS4hGdgr/vCSiEuMJI6rP/fhPC9iXWKKEtg/SYZOJm+u9tFzRRmLuraoXSp
n7P3Qcu9AC6lOQILRWCIsL52JKyvsD+rW4jgPhdXoGNyPjV5o63hdSt3cqy4WH2U
36HB0Yn/B8Mc2Sj/9kEsQpAcU23BVJtD8i4XuJUyIEESDPGWkP+J8UsF0xS0k+lV
4YEgjy6RQo/rE0KR2WgYFoBEm3Lg5LGjHvz+ytQlGsB+/CIL46Og8QapJp5brOfh
IyrI1cG9yhcPaGuKouRI8vgNT/EHdBMcKcOYfhczsZnTugD0yTPqrMzURxFyIfcc
xyHZNz4wvuWsqcdvYhqvCydUEIRsGJrYso1XdHlxZ9/hzghk+O8gHhXuZpBuFdiK
zAfHJ/oqMa2RNbNnQkM1ttIQGdhIc7Ub10nmC1cbiwYvFimJ7vQ3ntnFIsPy3OyH
GpzEOarsTwRZyFYq14oDOI0TIO+/bCf6lPQEoTD4ktuuFGOGQp0wBwjUig+XM1lF
4nPXLWjC9ytEmKnFuaPLrIa0jYam6ud+CvWaePELwC1zpAUs/6CURMsEO1SGqTon
oiOTUyk2ePGlFxemOdQhMmg/XWrUoynfo3QQW93dsWVIF+z+MMyE7PUqHChtf202
6/WhX4rimLwbEiZhfGMgI7xEPWeM1hj+B/46G8LGiyFC8aVXhCsnN34LEbCz5iyA
SF6OPQGSokUaoyO5+q4G4El0Nee3xP2LW2GvcH7HpZ/3hcSSd49TPxsTqr0fj3JF
0LjGUTv8hJ6rh5zDGVAheOLOsLaMaRio3rCmoY9o2frR/R3KGwRoHRohgMgSM62Q
gQKKmxZavhqDu2CW90JZREcGI0f+/MEJ2VTCBdnYyVFwu+ez5f38Jx0/T3uG4eti
GiR1ds3o3+EiGrFy7idRIpXdXDispkE0+p4mPD+8CEnGTYtAWox2uStfzuFkBizK
GYOmL5qXmXqyJ5WywlpzvJ8sKDrzMoCMTupMlkBEsH5wzgAuJoyabhrhwCnKAYfV
Z/cc/6bqF2Idm8XbBr8XtaeX9YPytHi1zQlS6FwDH/ShlZ/9Ar289LBLwGPDnthM
KACg5T82UH39lG7XhIsHlW4JIQpLsn6Zp2DWsT+B4iIXBClkb3i49FTLvgcDgxRz
2PblqwliUY5J1+Fkp/LMVj61bOo2dwKV2AOiqczj/s59IQyW2yN5tnltADgYz96Q
jiPidOkBGh3E7M0Z1OBkt5n8CmSc3XJIBLjawODxeO+rxMTg/c2uB6OUB6PUK1b7
Il/7lfELG5Xru+hnLDGal54Pi1mj9uROmZJahzYRvIeUWOcCvy1sEX5u2TXj3Mqf
pH2X6sFik3zrtXuWl/uVtQPfefmYWymC05gMiQnFTmXktQaxE8dNUM/toMbZX0B4
dwkPSP87ESanXsBftasg9Y1/YOYW3RrkC4Ecw/IkEZQo7ssR15JUbk05veA73wpZ
1Ix1xvvr5Y0lbw2AIVEE3ZEn9wOTZwpiFWvvNR5BMXd8yapInegmFeqHFilXEk3r
RySgTfmyIiuGcl1L2EKlq01WFMiXBPo4ujmhlHdvFyDM/RkgHGRTUcQHqTwREAVH
T7hpcdZ7rs75iBcqbSbopZAQ5XVDaJPtX/oxnoAZuNGrFNNe43SsdD8h/72V0vhl
aFatsvsp0P4l3t8yxbnzcFGJMYcfURFVoFCruj5AwzWTLnodghdN0dMturpaNvbi
rEjwaL4u/ZN8OW0UwygGFHmxB1ZQAmtZuG2nIuflICob8bqNZ1DkGuSZ5I4o4ZrW
0LQXaPE5+Q1yQFAoC84+LbbUZ716NBJ5bqH7X2z2byavs+CL8+tFi42bInt1bHQw
Nuz1p8NpbbhMCK0nA8aX6JG8nUaubJMtbom6/U5U5R2+HRFXYQrU4YQ6gBWBxKZf
rwOw/VnowLq01fmnL2j+3IjgHoYyzJCY7f07KeXnPZHBKaLgK40FynaJbh0fGtiv
0/Yyhv3g5HRtmNFx4U+Ilg+wsr5P+pxhjii/UrlEuSk3vYexouvRk3ouyKwkuUN9
vnKYwABc27qXjB0jaeYKidzBunDlHVBaDBJYFz2tWTj5BD3iO0IhtpqdKVI3QDG7
LL3bpW0NlpZdp9jXIT3lqSQJYGSb52xKKOSulTSEJyEm3NDmV8whNGumYW9kk/tJ
gNYBuqv/W/EQ87tddSLmcdhZ5H0NRRsMn0BRvxRHp0UOK+bqh+IYoclAw6oYfawu
HNePBuljRJN30TK35oBHRQ9AiXpBGYyJRC41x1wGcuvIe8zJYuj2xg5POeSIxIYA
IE6hIjVEnCO+DIkDZHvHyUaaTnWFhfAlV/J1OKAp0jpaOAv8lRJFE4QKSlDUUc29
pFVX/+qINQKd/fFCe7Xf7FDgC1ok+VS9WDmSdomcuwqkeW2lwt8I8APfEgN0h2KP
wgia8vaBYgY9YcAAZ1T0ttzO8eFjGTvy5BSJoE1MTau0SPNHuaYj+9CIZJETLVyl
6hYmp+5hGCunL8xDpBaLxtOOGJtnjcBlhsofNjA9xp0X60XmbX8b+zH9nFw+vAty
9OE9v09ZN/lJl7ImvPw0P3uy3FFBO6EC7Jee5vOiy/901H6pEgkWSwPJpliBnUxP
UJRehAhIgbtlldO3aQZsHvqYK+LRazw0kXAczFiKgR8VpQ7os3jvvD4YazzIY1wH
bT9owLVzypJEtKyVyeOG5gLNeSp4PgXqCm9thUczg6RNYHhwoAFY3vqe+wBoX8Iz
cZ7NhqidB52WB/UkgJbEEzMVaH3I4nZxx+bTPEzwcI7vm9f8mU1qgJw1al9xwSmT
vUSmMkI9qxpoXO8PxQS2ob8sppkZ0/D65x2YuRmoiFRury8Vm/1EptQa6/NxyudH
IlXhFlv+d4QtiEkvjUa+E/mkS0Noo4DWDFr6mn8GLCDZpw8gHd0i4N9Wn/NGU3QS
aEDBQHoPzNkPbKF1u/8rvGuZn0YwAKIeGv+Ro76zTlKaF6lLWawTCZZKFv8u77XK
nTCy5JaZkOCVLhuajEJ4WcTuqfW+VhI4zMPnvUIenlKgoG7KLnZRs6/m/LD3G8IU
+7jnuIfRMVZXJy3GCLzLBFtz+k7XDKNOFOmx626ACp46+Z24EVPZouzWo6qHxQAO
+gYCSskIrigLIwAIG1UhT9zQvYzIsIe2dGc3ASdKxUt6+LzneeQzE50jsPrkK/G0
F/7vnXzCWHLphwx00EBzMAPBpdg8sOGc5evbjktZETZe5j7iGRV5/521SeA2GGGV
OtWoZAGu9NYUcy402LYz/JqejqVy0ndgWM3PylXfclNnTiC+mSW0KR4xD4Ua/uUH
/jn5acd80CwyLK1W+WrSOELwVg2jd6SNseIlLeScyo0nW3pQYPcjh1WpAdFGP86l
7OaW/4gNtuTB4FQDuS4GDhJILrLzQbWfUjM7a/KHHqjK75D+SufHkdwEIvrnYr2S
sVx43AlIKxE0lcDB1wZqcC71stvSm/QAK9MF0k03Ca17R46KFGLKfjZavdwcEMkp
DFQkqjSgYnE+VT4ahacNJgpeVm4FGa7hGXYekwHjY18NNlbqXf8J6kB4VbEqBSq4
qQ3jwXqCOhbvaqsolRauwjZYD5TaLeiNKEkE7DKhwpRDa9z7gAj/sly88R+9xeyW
3vkQ4utRc2G7CTF05zkFwbqzJRfVXc5dlFIZrTou4+JXNH0hfulGy7uAphRSchhl
XMCadh2Ti4Zc8VA8DOgvyOeBhNZazQX2HV7qRX5Nclp6GsylnP3PTP1jzctyahlY
9AozLFWs/Px8vYi48qjIZVVf/J5uBT1w80kbd8MkTRUOnkmk6Be7w2d/EEGU+4PY
Tn5HupwrJ6mCom5zwcB+thLTaP0p3VgOGvDHD3XbtXizVT9/T40GpY85ncCtBZQg
qmdxmQwnLzb9mvsfz115VaEPrYjIl0SshRHYse5ie5aPTLIHzj+xTLyor3KvEGHf
LjeQ/p25BOBZwOW4WjDUZoMi61DXYM4s4AKJni9rFQMPVX9OFxIzcl3BTxN2d5x7
VDYOtrBS40UsvCvw270e1N4k8iSdXWRp0R4oGYuar+/j435bRgqTk2KLW1iVDb41
yHn8YiBJc9ZY4Hd8Q6WaJ3pqRqHP0MAHEzPjFMrbEbmEPLnTQLiMNWhGLcGq38td
7wIUK6192WDSYad2BO7dQFjWkYO9GWYt7bTNJo4k0f0oTSoTHoEzhOrWYqJfKW8d
Uj6T9kilmj8/BFTrXSu3szJzq47bgxRr/3REergdQPcy3Dj54xcmlB0EUHVht7ox
KqgEM9t5cLV4+GPrqi2xU3A5Tgm1kxXUR3C2wYWUzesNkyfZOXd1ZCJ297HmjR/Z
+nO26P1T2J+Z4qhk+NCkIKkUsb/H2GQ8j/r1+y0nqgPX2nJUNFodpIo3RHzMsDLA
jRPygCOhO6vxfbGCeTeiNkn3CWRDiJFGFss/oXcj8k+kzbbTeUNVTtvukdLDm4RR
mpKI1JEIulsEAjgbvW/vbCH/Uc2qtvY5YP3aofBhWtqBYt2hnAHgvH2tN/go/B/j
AIhCMaMucK5RcRlngPv17rZzpHYFn/EH4ntMkYd7v861gqTjaU3+LrLk9/FijIg0
N3dhBYPFScLFesFHvh5YFqJoEUAA1wIiT4506zvIH5XAvUGm0hTqTqUMJUMRaIW8
fYkB9qLekGx7lfYXyD8cuL9e+BNN2vzMFkYr5bEVVrzpfgziOQHhSoBw7wKc6V2Q
Gl7BNRfTTp+U7/cP8X7V+S8CZnjiweHZ4m5xvz2GfCXtsePKhyHT35UxhwVAD2HH
2f2v65SexhYtKq5F23MibWNEP7HQZP0iQBpY7x48s9ybD00M/+VBVfdcRT1/k6OD
pG5Yys9wF7cQQFiJON/1uAM++cK7Jy4d3dMSvdCH2MC++cNMmKvpPtnuxr+ZRnhu
i3nU0uLyckG3fiCtyA5M8Rax92NDYLJJQwS1uUWLuz/OHrq8Xzrufcqkrlg4ce6h
o9zxYf5hfH1s0TOpT5+1shxp29q0461j88fBuspiyfC344A2YCd62Hz2UWnjVUpO
WV0SyvZ3u6mDm5yQiM3jxHlo2+3D3Yj5xxQGFA2qVcvqCobtD+yK6kCIe/qdTpA+
sQTwUU2huSndhQYFghK4jr9W6F3Rtpu1G8ffplZpwMlLhUo6HBqLU0QeopDbzqgJ
kOPN8g/bac+swkHNAFGF5zHm97OVTyPoqQIY69+wkVQcSdXvWxVOu96hCnAzhrpk
GKYCROkrHuQR/w0hLyq+eQx8NGjDx87ewdTl1lSi+P3dDWB4Tise6GJFQ6wNq/dq
WqfKvtTHQcRiVbl2eztwHBUSlK0dSjMszPfk6el5lIjQxH4rT+Sne+cXK1mr+SAx
qEF/Nlef7Yd0AXaYYfjlJBtCxFmtyEHO2LqUSgKt/uCQcuF74J1DXQ+J21LMT1nm
qoUvZY9DMqwdCPAvyfT5i1uTxzppzxr1nwg/wWZF5+DJTiw6x1Cg4oPEoEondkIN
xmAleF/1sB3dupvr4qJ8B+nQ1c7wHikH65tMGAynGaDQlmNl9rQknLUqBY9N1Q4a
cCby9BZ+2yLGodPdONcXlxpBhore4C3tRZ1h/ophoIQg6rNxRUCLlUWsvRvg9gdM
JI+dQ+l0H+iMkG/Zl3mUiPzOT2D8LeFdIsvPGEuUiPIZaXjvDuRLHbQlR4OdC0hl
wJwmSK3X6ceWvNRXar52MSTTSl7f7HrK1uld32I31x3mRRgPyMtwpB8mEMQLk27L
2KG8+6QOfTEiJ77NN6CuYYCpUj3V3g0ZdEDzM+K03QtM/JxfxZw4QHyOEhQa5C+5
0zOHDCGix8dfWj1ql0XSUUiuaT/PP4l8lupitO6gpfIbBHFc0Jy/td0QIKbScfn4
regHW0ZtgFoSswIew9racso2OR+fywA7zQo0EkMo7enmaUvlZYyV2osNxPYVie68
klxLEDojyTNcEB1ScXUAeTgvhOGxbFbShgxCiPK2D5rTgPYWAUM8OynP/NrllI+b
EX8wFr2uRHOKYUiIScmqZsuD0k7bhEfvCDFYkARWo8oRF5v9ilJ/K6ySAbtWERh3
HWLUnmltezWeUz6HzF3/ZvgUR/n7iXIgL0c66NyhBe6Zkyq/YI5I3k9uoDiQGLZV
LNh9h4SoKuvn/saYTe9nnn8PxzbPwn5STSOBW4v9I9IGksp+SfkqJYmoZHWXkCHc
DFk7E34WPAoSP3AhraIMANWIjwvsb6iUi3hTzAfMXMwXwxIAq0xqKhYBz5xHcAhS
Ud4PV73H/7jB8elQ7Pu7d3hojGgsN+53kX2byXGkMqrJFbFX67SrFF0zXtf8cYKu
vA/O6hS2l9TpIdOvqNNbVQmPO0LA/Ue5yNV/7RQGPIV+d6YdWw6mfprmJDPBmxvO
USd9QeW+u7uE++RBIs86ixEwdzHAuY5vITBaHHkWY5xHsAWneRCTH7UKJXqu8prI
3nM4vlJSZRhSEg2HWzFUTKBW2etzESrofZD1NybezsxytqXLcUFjG7RADKRl50zN
aH0BG0MN6RQB5cBxKCrQ+CiGFjBuJdmW8I3bHXkFuSmbvEuMi73HqkeBj1SF5tFw
BqGnKjNOGOM6U9nJ6hORxQjv9LyVHB2laiWBFD1yE81Eg11pCVL6qrpke+Pg+qOX
L/ePavgVaE5wcFYthYKAH8mIWajOoptEwTpdWU5VvKszXHoTShJaU3QpO1EYqNf9
uUFBERkFgNLySCpgDF9h0utthREo+JTiIwJw2Q7CG1Ik7mT+ISedUwl8uoh286jx
W3pAFTUqWMZNDQUxjn5Mcj0eGSw6ZDqAlaXs9VerwnX3xxqDkaJ70qqJjowz/aDJ
FC9EVU1E1HT2SNbj/KKfmTgeK07AhK8OyQE9WEXcT3NmdHthmNztgXCRtflX49MN
+qfkG5Ea/owl3MQWujCt7+JW1gsw6JuhHGK6TgD5SHVzNViSFTFnmj1iBybAHK0Q
X1Ufi+7a+VvZrMdLHKodsjSFnBwWNtaUTMW1OEVQTLRBUNN12QZC1f3a1fvz2zCw
V/tRfTanH5lO0Lbdx1SFfXExSbBQ2uoJvGURh6lpBAZEzxZiEYytiTSFRTdeHfbY
BWdfJ9ZNFoNwvGD7Wh1eC1oqz4ZVvPIpmW8pbmDhnT+q+hHHfS2Jl9y/u/zXVuyz
+ltt6WNlqf2XxTASolsv6CudKTI/x5rYhIie7mFKfmWOOmElozi5tCk2RIUpZsO0
K/uAbYZtzUYkWL5RK+uWRnDQBqPBGd+/KNrQjTmudKUbj+DsEFUorac5uCjLzJg3
4fNsV3FO6HLlmYj53FmeeT/KhNCRHyHmiqcUrkD3L9Jb9a0Ky/EzJ7X2sd2GHufV
KHl5pigq6huebp1LBNI+h4CGn5BXPhZxVIIivc1aVctveIv9FO0XVHX8EYif9t2U
8zDfaRjIFaeSfUr/qGYRnBGOffT9dgmDpg+Ej8kcdlS/Zv8m0Tgq90Fxgbr2AMtn
aFBbqKhQR7QRGaOEioy9iJzqtPppi4EN+FQY8tDyG3ZfOvz+Lk7I3kaGaZ3wLyM4
WtdM44eRGOavcwjC7h0Xds3ZLWUsVByPlIkTa3ggj2RvqqHluJZdMIMorcbZdcOP
jLXEBiT5NwYdEVy9rEegqmIHJyLfxVgsGr6kUz0K21qleQNJJApT1/HAWgFinkPQ
pdF9urfFP0LRr1JOTiTNcHLfQQNGV5ILvklt9jXVZ+TLc7S3Zvm1cHZDugk4y+Tb
B3wYSLPjo3nFd9J+Vzm/0UP4y5n/uJCS2ZaC8xp/Yz4pYI8CeKxbk33X+EkT/HXj
4TNc5eYzewYm1bBHcg1IZdKPiDroirfuST5JbREKsVP3CEMEcwqGHBec3r7STIke
JF+Fk3aRgzcoFPCMaHZp2uqIVH0lt+qjdaVRy8wTEtJFcwbJkJJ5p6Mb++3np/hX
uiV5SVfdBBqW/6GJy5mnygVmmA0lwfJ8f+4E+VMh/WkPSIVAxj3XCBYnazvFLtrZ
Y/ouXMQ6Y/qi+nJD/mtEn5H0C5fyE1DzvVysQDkBl2Mq16KZNBex8z8Yx0QQkn3c
/9Z7pjT7K9wMBlzreDvK627cYvqSGPFzSZUsJ2ICUg0f/03FLWisa9iK0vi2746b
ET2sbjhcong54VwMdGjOzQDePG1XeyZKFwSpCFOM9ySDsEf5droqt6AOGF3yUrzk
ZKG9oK2oEzmprx0dTiU1+KpMeAUPqUqKkgylegWZKiRwxLCyrm9jvQEdjEExodnH
elonojpGRSEKWbnforHAmTeAkpXMWEHZFXdfnNcaOMwEQGp6xfo+awD+62cWcDwv
fUQjEzPO19ahhJslEe3cCnAjIXDs1nWeGGToPlh2tF5h508iSouhkjBRoqTtJ+Mk
DZQ+bJMFIRxFdwljGEvCct02/JV7KT15x+OJYW84fzD7XQrCAQTIUsrjEW9BwQ6d
4SlM5cDioezJHqY0Jpn9e4XbWXboVmnnyF4fWPKVMtqP4huDfIRvhbWpIT0CzrIZ
XCoXHThbTr5L5jKWPACR8KVWRHObpGWpb4WyuOb0viRbeg7nHT/iSbys3VL1J7+Z
/texyxIfS1NsJ/aP7pn7n5Xr/tXyeOaaeAzFNPz225ZbShTqQo4hoNZlmHG1moHQ
cLsWATrnH4VCUvhcul+nAaJcVRm2AyZe7Q/BNVYujvf8V8H60jSNGAw6QbqYdbHQ
Rz7vTVSALtUv/c3XH2+rCJ1wyTyc8PgR9SQvi9LrbK+Bk57+Xj7avL9gcLPxEF6l
xLBAQpE7n8nDzIsCCA9GfmfK82JlBRXQTGPgrJ10EihAx53ngxrB03jAJZF1RcMc
dxbv3sGdteL3EeHAMOZopB4Pb3Jhs6TmAtVfzySIL/5VnKZxx3x/zyjWRrF3lWwM
UcmONjDIKtbNJqALyXWErBFhRPhBW8nhUqQYYRfah+F2bcc4163zmmLInRcCd7e8
dTUvy3qRUXN1aovCSAxQfO2gcpvGkLKhev9T/GM6jy2+6upuqD+xzwoPcBClbixJ
ioq0pTR4sNdDZPmOMzuwwzQCUUbKZ79oFkpsFklSbh34xXm6WgfjmE4Hlr81FjLS
B1WCdC2TtMeMvSlURz+SkAj3J8Wwd+B30FXJaXYfczs7iIEsasBuIDJoFiFv3XOS
Co3lZpWqNcp61KtcMgJWCveXYHax8w2LmIy1sEV9zUBASrpLbQl/yVW/b7fA/xda
VUWQ4GLhPYzixzsbdREunAIBHTjkLM+KxSN4y+EoQhUuzWCVgND5zskad1oWbq8s
p3yZE6NkSiYVH9NQvE4eYR1jtHkF3hiNl2ZVGjnge8l5jhXx/+A2+BG9WLzs6XH+
3elIeY5r8wHLQi01HQABZa2F/MGntHAyY7DZrUxACMs1HCn8O796LmPQ3iuGif8t
LQF+JUmfUqbrJ45HTWloviGaYEN+62RFmbknPLouewZHUUFiytNqxLTL9uG06+pr
irpsukxRmhQUtJy9GV/HcjHbNA6zhJjPuWW5PaF0aJGHgSG52vdWKDYeG83tp/JY
uWo2cEh0/iGDzR1YSQFmb29TJkxKccdWzXN65P5xhcrPIvjDAJluHq5cDgQs/Zim
GkWWk1VAK9vcYEag3uDFoE472qaRSEjvZT0UtxlcPVZPW1N3qQB8E7ac5ChJCd4e
XwnRfeGvOMYcOBq7+8GXwvGSucnjeZyRDG8M5PCtHHP9oJfPnbaXV/HFbn11nlh2
hB/KD/ippUqPd6Qa5MUQIOcOuamIvPDu4abDYj5Z1KqZNqdxREeYqPOfDq6woXWe
ejurv+eWsV8GnYK/vc/hzV4N/PjhYY9DX2NcxrbaYG1b4Sqe2yyaIgA9CoDmFLiN
ShiaAkYAwNYyS5AqFXg4K6xJ59TYX6oUp6fWoBWkfejQykJ+1jmi0bejJVe45sds
Q5wTM0DVQPWAXjujljgUEOOMXXMZlEJbJTkqGC1owdCT+0ZUHkwsIbiovf08HpIn
pcf/4fWa+nXlsze96G0F/6pDfkIoWlcn1GTz3UBsfk1XVt53etoYM3NprSORPmXc
yYeo3IFluiedeH5c4pa2i/Adf2mKH2EhgNownxHRJ5XlKP0FMrqpUc/r5TI2U7xI
2jQpzce4Vv8zzEPUph63H/x4NNV6KU4pdi61mo8BT/51J8f4pLXePOz9Yzo7uL/1
as7pQ4iGc9GpBLvv9Fmb5U1fPWB4miWcKdyf6ugQdLxaTQU+OW1VWFkd8urolqM5
WZQ+z6hkmsJKY2KcVgYr9uDGY5xEHrXISFOmJ1XhcNmZSXjwFReEoaYK/uMctbzE
sK58uYKs4/GHDQz95Wrr6kh46DYLV60C8ixvJx7627CXyTiiO2pSMlzBxSJ/P43y
AhdyP905kB54bIlVS9sc7h07ixTyTmvNI3KNKmU71155WZDVZEz9FYawR28n/KFD
v0ziDG8RiKtKzxwlwpsFbHS2Pt0KCmWVvqA9LeQLTYcImawSX/5Ko4mQUVpL6re8
1xVHyE47+BBJEcz4NjhwTDD+kXdPlk1d+kHtX0CSzx48zBPWGRylv2fqDqtadhLt
nDCEqMFI1EtfICWbb/OrE43yFaWFNl8hXYOdUkHGwdp+YMhsIqT/0ua3FDS5ETQk
gGYmfIul0galkzJ5doPBmrlfubiSv3Y1v0x+fu0tkkNhvnCeY1T/O1mFR6kufFGv
pd+g3kt1+UdwYExEpdDjOD9Ajyi7Z4qDYXZ9aNVEZmCPDkdLaVS3kRpuaefX4gdR
9eFdxnionujtkKGMbRnU4uTRop8tz3J5ZIHHxuBhbzrgRN2g0fp/WesmOE9R5ZSs
uYIlKQj7BLGmcRg+Mh8xt0ky3yuEXY0cbkW1WyooOIXXb7NGOv/hotyahqk4JfqO
JkUs/6/uioe2RKrjAjc2RdevN3O6WbD21Hd8lovYbe1YKCIMK6xjbdwRC3Y47fWd
uyuI5UVINs7csQn7wHb1VnEHAm1Ruy7egc7rc8Uh/r979lWhylupS4JCA5q7i2IE
jNa9qUjxpZwApzZ2/hqyAGwkQM57UJijPOMYVo/qeqqMwTqX109yZnldb6r1Dvxv
ieKC/ewkyYFYEkfn/4rRjLJv7gbCIFWcGwpEzU1cNsshKXVGZGsLjlkOGXAJ9pLB
0PoZ3cn2WOJ6z/gA7NwLi3oYLODbo1O4v7riZvb4Yl1MSThaICaf7Bee3yml7PAZ
KKfHuGF3NK54ezr2jLSG7SoPLAzXykx6Jb5Azk5dDY8P2vV31L9cPMKlDvb7ZoMZ
PO4h5ym1R1A/X3la62H3ZnwzHqyJoBCdjbi7BeVfRiYKNMPjRSHP/v0KGpHiT3mv
EzTmhI2nWj7JKkXpF0wXzqkHtOKdB9WDqEHJapfzKco06NKyEftg2I7L3SBY1ly7
oGR1qdOEfJ5Ni8gXahAN/sHW/CdZ3XZDD8jXMpZmz2sLhaUnGzKnAXG1tQe9X+Db
gilZ4CstIsnU2sZXztKtUJrt+nKPJLHOU8donzeyJjd/bmaApOIR8G1Xj0E1S6O/
lbYuT4P9jPDi3L8aO5xR0zKKApodVvJoaVSsSjE1fGBrzetWXaZCc0m9q1XVLshc
7keiL+NHJPruRlS1eOdRw6z9NJMMILl8v/BqNdMOcsR2LwtXVSQFvLy0ohg9udrR
u0WMqB10xTwrFh1z8EGRqg4miFOz4IvSz00BCNUCO8A+ccvhpL30vaealZtiPAZP
lQzD58hRppjN18gf5liFueAGbSHP0QY1yazaWcNMzga6teTWZ6NK7DqxvBD1OnG8
R90dSWq1mxS6GJus74g2UD2X4ER99JB7lMO/CDeGZvv6Gmux/M3xLdmh9dbI3roK
kJrmg5PoeGzQUBOTWzdOQEQK5kwbHPWOIs906XoUmguztpbjgw0VLLAlqGdbMddP
4tw9tVivLtIY3LdfvmEnC9le1aXj1zMnVt3Gn5EnLtlsBHsto38EwvwijWg++HQi
ywuk/jbtZoWYB0oPiR6ibIIPqDm/qFsis+1JYEK6fh6Iq0gS7O8lwqyleGHEGZnm
8F8YvImO6ENRR0kXk1BHoAA39sU6McM0WIhcAWlihr2uGGFtHE7+6Zlp0le6FVLs
CGJwPZQcICXFriccjLJHBmu3DDLpcQBXZs5rAqAdfCl8SPqyukxo0fbtR0ds4XMi
Av+MVNE1R3SZFI001pLFRQkPXZS5ICnUGxIlKvYy1KKvtlHSU6SxDU/3rjsJ7M+t
wrdH93kK1iO8UYsI6OTIEUwZgheIutbzkG8p/zyIDxzbiCuecpyaux7HQ4aGAYVv
I53gfV0DY3mA7BNqvIMKFHp12oTwNZAYwEqkA9JvT/IVMy9m/ThU/ync2AQ3VLti
tvKXaSBL7h65x/XZNV3rTmH2ql02/LklI7wI/plZeAMtLs0qBmt9F57pef7IbRC2
9dvO1cS4dknchUN3nw8yYVVAdeTtPOh29IoJSBiAg9DHlhoXTJHz7mMvZs18pm8K
0Xl0n+nwym8MV8bGpPDIR9gah2gCu+NmawNYb/Ro+nKL0HPIQeujoQHfkxbzc9Ig
OlHoqjmsPPuNxlVmHHiiEwcYXNu1Amk56Z1tHte53H3euyuJKDT39D1igVf5lpEO
10CruP9RrNvI2C3ZBtQtkC6GUorW0mUPKuS+NIodEnr6wINCnnfr5X/bf6qHbss/
nQ1wuYSCMrJPpSkn1B2LnXKxDsYlZeNWIiEoDtg6MrcLQs/9Y9IBjui8eeH+JymI
9/4K25wvJF2G/jBVr3kW1G08ap0pKaPzRSmziYrPP9dE8YMkixnDULUOENpO5gUv
+3tziHiOYjlqZ/4fcROGhmjZ3/IPIGoZvPn+ZZDzCsLqFq0ifvoUnuozOffPtOAT
KaudgLr2HoxAm7WdWpSw+HgUlZy3gRyPpLFqI//xfe9r1y9xP+vwlPbtTaMZPWpg
G19JA2DKbYqGvv352Hhvjnck2sukRf+jPNBZGCjWGl0nrR6d1MQuOer55IHrDNeW
3goXfK99J121ncaFdtXRcyiBy9Pozx3JBf2fDeu/Ehnqf1Toq3zNLVHn4kEWNp6R
K08I0aaG16/fIRL8oqa+bEfsUhQkGXkR8GwrnXNB7Xl9/e1jJKJ8LSvEivjf6RbC
nNVXEFUWo+wqhuw5q/ISDQGOT6VZYRKyGuKHFdyt0VfUgEOk9Jx4fLSEYSkmW1f8
t1+iOpQq0nsSYfCM7dB/yjdyoj+Ngd5f+Bvovd9QoK0aMxns4rgxKSMLIse4N/aZ
/97OKtfGGZbe2nCuSt+pXnBuF3yg5s/9W6Sdly7sHaLtMUmXu8LJ4sKxAifjNBoo
86AJrOyAihRx+tllefg8Iu6j1qPakvW7KHfZdnwrZd7CanQfqaGQn/cd2MiJJmRw
arFJaDFWYfx3DUPrY22riZqrymtiDTwMgr9Y2z37t66Uoo6jQObfmBwv4A4N82ht
QLk6fEjXmhyhWJ0yvO/J2X5zRYULazI3PEq2u08ARmRaGwd1x8Z1UBlmUPbGHNB5
WD+47qPPUOfxLJGHyWrxTIWmh5bo6P3FYalmc+5EXZOJQHFUJdAe9FmoPfjhi5qK
+wr5C1KLowTc31mTJtbO7EzyrKyFBjSz4ieFfIkFDCI7gyTh+raFd9TffDeiquZc
wMbRx0U9lAohRmce2AYQfjU86CQ/2mhozim9s/zi1ONZsU9j7W2GEaSmBGw+Ylf/
KbmUs2WSLd9XL7lBkIammaJWEIU7DPBuDayJDParc1p0x7vpT1TLVx2F6fUwD8MP
lvaloZdGtm44M6FWCqJyAV14QL+ZFGc0vRhSiwJ1Rp7e+/LQxt3yaJqmQnjy30ws
F683MMzDoUuOWEuMFAdIoINBsz7QTonreKSyCfxkfeKwxvL8CNAsA6V9n0/nAEKk
TrVg8ZH/tqnE8gxWLY3BiHmyqo/duV/VRx7Pm5J3hhzjo+k1C07RYhtFTDefDyoV
KbGeEhNgu8BL0iTc+K86PIDhbihoEHhUYLDAXytofQ552Q0/uM/JYV49skkoseqy
qmYsBwtO/smjQchMwnoZk/CropmDgNA9W0HKmhmmC7A5cinI1ITRclugXArT4A1G
5Mw9kRTFDsoan4jWaAho6TWYsw7mbSIqGd87Zp8GByJNcnfDPj33EF3mHB1kh3E1
2HIjnYRsbHNfO9vvFlC/DweZZ+BCW1NYJZ7I1YruLD999kqw1sUTyPSNUscB94pm
pPGu1bFcrDPqKIbKUph2DODcWEXge60B4bOvZrpUTMg+Hs5/E2bSQbEdHiARZE3Q
TapcKIvQBm7yaomvvD1cr8f6DhuSE/0huf4/LW51FY6yB6oI/2tWP0d5OLSgSX3E
DhoKCJIuEyGcZ7U2Q6o5W+YNhSdu2ihRVqjofq3lg49vvwCcl33VlasBtt+XPeEw
KVAB05s0tYi2W8INZ5SL5H5YWaG+6+5IvQvv+1mB+p+8y9eNdJbl6IkgEKi5MgjC
/NVmSsszTWFf+wBCaNX/eeykCWO1/P28JNdigJo0fXjlpBudRbh6y5CrPsqutJk9
9Q3ZMCEyAatL+2IGGafDohSOX7vyFQF7geb5S600WbUbp4kPDVUuHQQj/BwriKQ1
Ys1PQlBJ1st16l+WhLv+Ex/YV2yzfE3t42ZrOGCw4QaL/JgIQIU8aAcJM78/vPh6
Xux0bTRCQ/Y4BJRTSOxPWGhZnyOWSbIB1GqRLzJlmGzAIwVutKyB2C6ttYhSIveB
0t6tOjs/diYR1RApWkHZmULTqY/i7yeRFosVhc32UFk/2zRc7XKq9iwVTM6Xw3Ej
fS0C3k1El0KjV8tRIjJeM7PN2Mk32moGZqzI+lOBP1y3g9zotXB/tyZCKG5SwrOU
o0J/X2wPAVqagIA+4dorY4Fp59pd+X/ioxVnAY/bNWY8/I4PfzZ0MRhnYDhdZaWi
EPdk5pytq7ltDjHbo2WUJx6wbNoVJHJYiCjIux9ve+DchCsdMY9yfnHfjmm/9YqU
+4Di71KR6JG+7yOjTRuQ9p0fTh/pBakP6zj6sGR9STwmBChx93x/40Re9w7Xkbg1
t9iYrraWRbeA9RA4/VKPVvrIHT4lcgkNvmntHkv9rnTCDoRe0Yy7CidZBDGlylOO
CyEi7suk5EoUzZFqOiRUq5k36mGblA0TgxkBC/VCNVTaLOL4OSHBtL8hZ+uKFjYy
4fVvgGsLSZjpGBJGOj6CGjb7vc1KduYAs/wIsOogo3eqtfJPYDpdEGKwy7ZzM9Is
N+R1GvFMWRF3rouCLHYewzA83th7ZU5lQsPtYjQiadOgPgkO7dQjana5s4lvrIDC
Z93z76JeY1gJKzgc9EaVyAIrPGAUE6bJBsr4Ey/WRfjWxP+AUn5UvFQ/qy2xkU2o
QfOzrAORDHZM9wPDPROoMS7jbrvU0KlAf00LK/IhfC2bPaUC60uxKUsrsTKHB/zP
dn7UnUeaOsm1pUJmvyxYoXyqVyNk1x+4ZQ8pYFXWJMYUbl12J1g9vOsKRDb121QI
cJHY6xCVSI4VClbXlTJDG8AEW4deOlhY1ghxu+KJ2ba+8avKfeZTDtAPfQLpT1Z+
wTJiS1oFpLydlAk+8Vc9aXlBysxkGyGgEXsBJ3XcqcbYImDrr1o23ENA9FuMnLPq
fe0HwtyWNw/8Kzi/QjNZfilWnhvBEnU9Cu3MzBv5USSYFmgb/fv/v7UGinTtySvQ
COwSl9K3yPkJgSAO0p7A1fT+CYXKUlQ+wiHQerCSIUAaiZlfJXuJb1mYT/+ZvnEP
6gyK2r602t18K/CwrriIgJaiQYW703UWh0rIj8yOIP7DG/H0H6L03ll8tp5+aprg
USXMvoqvxJLKuFJUDuv60rOEaOnmUz9DNi8O4q0kgApvC6cvpIF1RRdoIeYTTgI9
vMbQkz0b+093+2wjJWW6ylGAH/fXltGTeTE4AuprsHuzJSfHjJkR0UIOvshJBHxN
NcYxefgiWxCvfjCUEvEBTSd3QxjOdq6PxwxExXE3ZjxM2oaKmiOe+KJeIGoLwyM/
ZkTZ7p6oi8VnSW9tZP2nkZmjsF4D9AP45cUJPSYvmtCBqBTctD5j7Ewazbm0GDNd
eUGw/kgXzgR+tZUtEOoGfD302DTLFf74S1li2nEycAnHLprt1sZHeCSLc3xh/Q49
dHBVDQFdwiDM32kmxEZa7apWfY31Rdpdd9XkYLLxmHw0sKLHSllr5Uwptxkbca5a
p5MNWbAfzw5y1U/EHPQBa5qT5fAefwF5VBjh2c7Ov9i3J5wpCxeAXdiAiy6xUo9J
yaH4xmeglM4R4n+Szm71COF2whdAACnYg7BpcDsKImZmpeuWq1Tn3ZYozWRuPYqf
VisE11dm1eUM3zGY8/kujWOsBY1S0n466HbBqrVhuaPvqP/hYy6nF88I+yrzBAaF
zl5CJ0djET1iEVUqrAvuwb0O8RHuT+8mN0tyNoCfyjzfyvR06/WLqPB+pEWUl+wb
hetJK7z6gfvlisOhYuwY3aNGAwot0IygvrVNr7YA5HYUQ854TMX/V1yxswFc3wam
ROmv6nhr2fFoSliKSSkIrmMibChE72eNhIJ923ae6BWt42WXQrolcFWl4lfJB+/d
UVdX9lyC9bmW/bNeO61JNpAsXeCEGoHaI2Ru+LrF1cqUyRODBp0NSCzwnmolX8TC
CxKl5+0VWzc0ty78fekziWAgbbODUZZy17zCdlZiwqfluTq0A/NyXI+jdv6g1gii
B6HbG8MPaEOckxwGEUavNi1AiYV2xoQgNVnjt10+32AYRmE0hHDe6Qy4WkkY/K0a
aS8+ZbdQJSfyTIF3xwCAnoIWGfIHCtZRTzIdyeLlBWLS9EowngSJAAaxsPGlAY1P
aKd+aZmAu1swDCF2p2bGlMhpo+iBYYjMAvaGoA9Y5MiSljsE+sskqeyo5a5f29t5
TakZQprDDkfcWHj5Zlin6e+EQbbQovj5F7bkOye0kEVsDGCTYWcOsc81bJdEk9VT
lZgt/x7KP+v09FnpZrDa0Ozl9ZWd10KQq6lAQqxTshXcmqx+UbHXtcqkP8OPsnPb
BvWMKEBS1+04zXsmgD4J5QwhTkZa6OkiDlxUiyVf01KQ8mZWLlW1IOD5jyZeuCpg
Z9ivvZkKwRITt4Gy7GXTQjS6bYUGq2DlD3/FgAfLm8tN3whvFGax0JJB6MgUs3GR
6+1k8UP1xgCqNTQgklQe8zp/stUL0/rsoNxPxiheGmvgrT4bKb95vDKPGYqe/tPm
CsJFP+eCYI9eDpya3vKmbeySy4FGmKK0AvWbtz1odOQ5mpJL3GAfYnC9W7m+aKF1
hB3ocgLc2Y92JB5ai5LJpF+pEI9/Rzkh7S5mxzib5NUtZ5M43gUd+6SfDYVKJ3NC
EXv+qdNXGt1HfL5bhQ7V2U8dmtpvCxTp6mlJSCd03qv5QaBCzrBxG+I8zlMBptU4
SS31n/hv2vJuP8PCCZaeI0cBid4Ey2aAel72FkWUkzf4JmyjubIprcfFqKsoL9jS
u+3No+EAuFlQLraT2iJpSdEwROwnBlJWNjqfv8l9jybAlYios8behJFGtljTg9NF
LmTgNlQGRALDEbUHEZRoj25LAjSMfey7FH2e3eyztpUqW/NAYS+U3uEE+B2v1o8g
uvKVbzVhqwQyNnGqRCjFMaBYuQfjm9Yy0SVoyKWO8H+Ma8dNYgASIeHkIl9PxXAH
NvK/Mj1E1X/T32dQXDc6NcyOKtG1onuadfQL7QF25nhLDFzxHXoIb02xA/R2HsTi
rcLB155J2QvnbvPem/fcxO4aUYTFK1he95XDcB/TiLcaIzYAexb2d5KVShSO6OwU
xrp/lrxziqZ8GHwKwQwN/zorK5n39fWrsGTXRh9jbavkX3iPBeHJomak7ANUd01M
HOx9FZpIuxVhjaV720D52Cw6xX6H164P6WLEkfJxbJta5FoOl/SIZoW64GRMtJiq
aTNWN2h5Qk8jnPJ2XO/6lTaDU3GaomqjuOoqvgSKZqby2pT7pThGrFpMYtAHngKw
fCj9ZAXC4IFceTEgp7hhqYBPS5A+ThbBrdV35g2FiM3JrMKyW6lR2Dj3hAPdRCpY
TelA8ReOviMt5tHJc19h4bwNMUEAqxXgWb9X49yTzh/ocBv3RemcBGrAH66g6pm2
KeyJH8HRaaHqifS5/NxWNXMGg/dKZLtoqKSDlbV++UR/w0KBpRnO7zSE7HmIQ/59
MAN9bMJ6VPfSUnNjD688u3IcwGjSQMLZucv1AG183D+DxKZn9X6LfP4nyrhoodkz
4uo01qoMxn3xfG3uwcx5dZDsmfSycMP0xBusAJ9nPA3QwrSdTWQBTOUdRwKPU9QC
2G6oqDFiTnd7Q7lozJrZlaIBDvvCziqL9aIb7ljdhuaVGel1BOpdij5JFxJIj8uj
nMXqPAWBIsNEhti+hAiMkgtMPWWlIzN2A5uIhxcG6dRUm49BvSesb4dKfMFfNIYM
mMz7ScuQkfY1NJBvEscvGZsB29e3S2LVBeL7PT/HGkKhYFsNfyAl29tmcvPPJvIn
FYEzbCIur6hXVQ0evBTW5SzrH+ChNL68ue+oiJ/L/+pgt8qpMbgRymdZxYubmQtX
ImzjkZyyn1wEh3wU509hccIs+DkVF/Zuwgq35L0U8P/HgwmeAy8b0j7tNW73FIS2
hWy42EPfZWWHFDE/Og9d4srSFfKg6mN+zoW2ACey0tAtvvJWFPlo2y+kDrbwESpw
ZuA9IV+pNtxm7rT6pKLmu0oGTFnbYAdExEEH4GOuvIyfEpYIu7tzE1uAoysQCszD
O4WjS7PThQuYaOfe6hGuFBsOJd7nCdIy0BVYR4akFDdewooQCVtzAdfAhhkRIcvx
I2up8F425tK3fKU/cyprQNzoaK9fkq5LCXlry5n8+Ebdbx3ZafXz9PWbKjjrnig+
o4bdMmjWPUKknR+vG+hnXSWOz14Kd+2B+qTgP9TC3mtzxOy/Kgo6P6409xJLkHSK
KJc2JgskAbTPBYLKwN7pluYEs5I6m89q3KvyCfscwzm36KmxAXEfQdAo16lmG07T
99n5E12tkK0NOnE3AsldHCQX5WGiNCgYCBSJopy7chpknvEjSs2JGd23w5Gww8J0
cIbG/3FEOoQxozXaG6JViv2mIWBseUZTOn683iIFChrYlkw2ZQ7qajJkt286nNeA
ro3MhFQ1neX6FoZmzJlKRf1DIcsc1gA7JOmdZBSRHeNxhw6tyRTadY90ORZWDrJD
+PipFbnyquqGSleHdc5lSQ/moD32z1ZQO+rXzF1uVzEXoR3OXt7YbiNXvQ6dlVNd
xxVg4LauOq1kwB1wdq4GM5mzZgKCbHa+fnEAc3FetXkzRkY6W0947DfIAQDE2M4g
Lpg3zFkOgB+YT7fXnKOtK0Pdw+Q9SflGHlZmlZ2WnyWqmCJU+pBqnh/54nlMyNsA
ie1x8NqU8EnlQzDAnl/vv2cx8s2GS6u7TXkbLSGJ1+YYfyfKVoiDXPhEAUsqZ5Um
V+90tjk/dKKKip1mVfaZ1pHFdlUu5zlvvGy+XZqRPefkH1FCq5pRM12CBDzjvAKN
E0qcHCChrHRyFVIOKSpiCpSGobIntREnHxus3ENvyt+PqqlIL7b4Z8wqBAAGzXKb
OZnEkLKz5sDjpWkoCEQoiXvb22KFAm/yo88/IEWzXXbe9FO3x0r74YJt6K1p4ial
mSYHsWiZZ2dNT6s4hxIwU/ymsvzrasLf9QUdYxEOgToM1YX7tgs3tAhonLOuEh2s
EBLVtM02axNqdDvEc9v4vCZzf84+13y+S0MNT7IuLynV7+vw7HSTGHIBi99mZZBi
EkfSofyfTqvaxMjDwZ8QvUz3m2G/GalO8w8WFZvOOwXwGI1HTL6X73L94KFHLFtb
vy2pIHusvkJ23VRyFVn4ujB7Yl2IvKKv1hwfPBt5ET55+I985FNlfFFWPnqWAaHm
zcYIX9KakdMkXWkgZCColt4UTziDe80Lt0GuxiYWjHDZ5aGq9k1yb3X+T7blqPtd
wwzfFkB1mMMkLyduvb6ay2rtk2TnuuKrdttf0M4u0BDbZPD5Sv/ZdH5g2BgELPsx
BZhDbGUEpeZwubH18DG9fdQpyV3t9lihc1gufTeHYYXurEUB0MwWpmS/qJVCsYqb
2uz0mv6U/pMla3qUOwb0HVn0DFBGFQJew8rfHg0xsiAtP1Rez+XJUtdunzNoK7CV
acAaDmV/xUiHA5apn/37eEbGvLpiHbWLSGVxqkiwMB6CP6fbMi06M0fUQXasLdx1
m1ffDlVIMkGUwwIUSSFLaaNLSJdMKtR1bQxOAFSMcdOAYaBw6WVg50Klx+KWGPgM
jwXtm9OwbCl7K1ne5F/mGr44DHH9er91Jm/EGt0dcbcMFNFS19IVM4BYz2j7EzCm
p6gjRKda4+db7FeMAlgtxqwAr0kj2Mv+DWvTuRUQcYFxosrNKZaarv6suAMQh3bG
xnfozXhkLaKy79MXsjqX/OT7H5jLm1W1q5Ca8PIw3VS5StBb+cfqIc0YCHXTMRxV
N1iMnRFtbjyziOHC3GHkKHK5KlN4c9sLwuFu5N76AYOKWogEQqfdGBOYaWPxdewE
zdP7+7Ka7VNeXPAvSxi0p77CK0P+tPGI4XiJ2hhwlGmEvTF5UDScE8XBhGs+d7S2
n8aHTrrsr8yeTqdhAWOyn8DjMA8sxDoTUKipdk5d9s4mrTv4TySgXCVtQxXDgFDA
YzVXWxuaSjXwTcM7+n+w5lvkUInBfHcMFOEg+JsSqeOydDKZ8Y+Ikq0DDFcqvxnM
YSYCQOaEK7UeTRRKO3QYbG2ioed+VDN3b0KTd47gz4Q2cjLDQWssVNoWr5QD9OUI
20+t0MUgqlMaelADpXxJ60s53XrQ2mQZmBLN0eZpXPXzCuD+iKt1i6JXCNgENMvZ
cu0cGHSg/5pAGmmMBNE0/pzFqQqBu1aUwBzXc5usa2bAFifyzp6O8TzsObQBj4LN
OCnY9625YmNiKlH7TjICkAS9c/5jsVYhmdYR5NikSO+o3JoIWwF3leO6vbICNSqd
5zLCDX9/2py0FI7RY8/M1rF5AgNO3233hDuXG6DHrxzbjWfLzQdMMZoUSjPI1Tki
1h+B11xLCJWv91OAvLw/q/Rz+iQs1soCzJiylxxKuTi5Kgyb4di9yloh3Zvmqxgo
uC4UPlMGXKhwE3i1BnyfkAdOpza9Eq3MMN1sK16DEE/pxBeiGxx8P8UePSDVejQO
oQvJ9j+BekeW/QdKAFUAIaHSofnnGUCfs22q9YLKqHy4PzFgzKWVb6sRkfaJ1wfg
F2MyaTA2QR4b8B9zcz5CTrBROUBtb8zrj9GdH6ssLXFTkeCaCTb1J8eNiLjk+5WQ
QkL9HW5uJXdsnK/WPSBGD80GkPYqzt72CKykckvAEyA080RhlsN52RfqqnTBOb5f
GCKaGr2UCH3IEnWm+aSM3ZqI/HaMo9OJsA6iTw3l4MsF0rDEOlyt4kXpo7XK+ML/
oh5IUPLAgo0ktqjJKKrnpGDO4B/UxFK35kXxpwGvKgqmalLm+hs+tum0LdNZXYtO
e+cZylE3JA+s6/Nqm1+bYMgkdWFDtcjSJadXTF6Vn7VrFhqQDacDBnspSmOgZo+U
IKVhE56sRkC3lMAIUJHTj+E11pzXbcHw9CDxLlIalBwZTxYFIjFvCibeWbZTaSe+
SeGHkdkCvc2L2Xds0UaGXjKCcRzh2axd5qPlp4kXxttpTCFG9BuhZ2ocN9oq2SqO
FNBT6gUWGpnnAXbi/8pVqSB8eZ+LqkxzUXw/QoWu3JIXy7K5U7iNM6r5Cmk0847U
JubQ0ZOifjuUPxZnV2iUhpYs/qfkAkjV4U171MPKEUtNIWCW7qVoO7xNIdvzfrqY
d3njECP+b/be/ZU1uzmczjWXzmKk0pdPMovnFjvDcGg+47S07KMURqNktQjsvWwR
LsiATVi126qdJq2mRxcATopvoEcEFEHVvZTNC8+1q7jJNEdZkDbn5dI6lyyKY4Nn
rTVyD67i8UWS/TUEDHfcoomle96EV2+4VSefweKaHIlXiRiWFbm+6wgNWMtxKjEf
d1sdCg9bncSnsYQZBfTd5PQnH49p0BoIvruM5Ui/4rqpYktZQHfmS/wjSbJH254g
gzrLx5B8xd5mnD0aWWqN2q0vtbhDhuJCqDdLeZCNmDstDpVxnieaBMzcSeQ4G+ac
j2zkRzvzdOEJEZo5L1tHupfQcAW3B4oDDWv0zv5AmtgI4EjrHABCfkwOdHUFBhNB
4qfVDtOVM8nvguiWGTEc8dwjCcsk0k5utYB6/dKTnLuGdH1arTfnD1En/CphE8jm
6o4VJW8dtAKDs5yMC2ed0r+JcJsADx4HZQkCvQ3SdNWEr0UVZHUgr+J+xPXKnfVG
D5VfNx9Pnboa3jOey6hFVBpYl28ErEEOcGi+QFKSy8L4emOknW7hJCgArB8mJNj6
Hwej4IARnX76/s/qf62ULOMvqUSj9Ce72eq3ppJ5kZqeRKfr0mz+AGin7CYDeVHD
uu9a6wJEgumw0nHjLM1FafJ/P9Ellp8aOdk3xpWOKxKBllpf9dx1lMthw0yDbYmu
A3TdYfGlCf+XxIk1Vm+H0l1r64dq6Ek0ApN3BbYUKGbQnnwwKJkGPmIXSjR/Xie4
tHzaPRp8UO3y8KZDSupX5Rwm+6VSWD7ovbB49o+UX0sYFAyHvkwHZteqh7hpytJg
8AMyhpguoLFhxL633fn9jeiWl5HwdJxInbVF2u1+xyQqNZGiApO2sjA+b3+PLEj8
qyS7Kpk6RnZn6LbY2tpSl+KDh4bMKy4+hJi0Xj42hv8sLbwZMcThX37MmZ03yCUD
Z9nK2IkTriat4bN8WBCe59GxMHSlcHf4/aEO5mME24EnfYVwoYGsTmgt6RaPDW6+
uUb2zrpqZMP/i8CIfPe4OL2DE1mH2mdy6SQPJ1RQXFmOsQm9TNpnht/f/pPYur9C
hoUi/StSLSt8iIxQAl6+mEJNFjeJm72T5Iw3tTDk7/9xpZ5U+cXyznSxDX2+Hgv2
I8/OzufJriB8ymXiB1yuVkHRCzBj4ZrbUW3vpERJ3ZPo4Km7OSNoJstjxOdNqBd5
B4CsjTu29ewowWEYZM8BuvEjoW79CZI7T7yFLSaRaZLYf3ghXNNE/B7v6+5iOES3
WWDdJZ9yxOy8EcFzUoTvnwugHPyUckm2VdLakMdWvmxHzDQOweyGgo4wROMBZnMQ
Ft3S1JetIeE462TYTsJ8bhhHY7KI4vWh+yehNGayMD9MMeI06hOYYuaJzcq4Xsvo
h/0KVe0yiKvxWStV1HSG+jTRMigNN98h0HMT4PGUkBCMNdjdXjhrQdftm2edxWrH
2NzT5DCkoS4dxFFFvUOCTuGveXESRCmmgDTOR2q+lGQntjJn0Y7hwsb75vvaCeny
gIXmj7TVm14xcQVMXwI/LkuXJwk0FNyjV+HukizqQED0Z9tSnp4rXdsMkjgzB+6I
Z7avYCybvK2DZnOoupEq9L9GmGegVa2DW2AmxU0WT2QXEFy0lMHQs3Zc64+egRGF
IdXKC+bLjKmXLtcWYGy1QT877FqCEt4Ufa1QzNtBt0jfDry3NDn/kh2ZbA9eBbEy
oLSjQjHIPbHuU9uO2Nq0f0WuWzt7FGCuiARZi/BOGrh/TQeuXauxIwU+W9TvqZbm
ialyUfwUYG61y1/8oSuUNZAHjvEt64TkMvmI33KpXWJ/ohTDsLPuus1EcdNw9CzF
rBdwfJV5PqodX1cMR1l67BSieuI6P7IohyHmVBW2ZRO+plofaSRB82p+B6sZLowy
+kyROEf+IiNjZjK0TAPa2kvgpa+Hq/MsQ5yVmRouhdFxM7v/R8pQfcSE2AOWaGqN
GOcqgabvipulqP4TwpFEzd7mL2J+0fR8tRRBgav2L83EvUdPaywCtp93pe2KujVc
qkGGYE+sd7yIQ/oYLC7lrz11RNMoaa6XMfFhgPjJKcxvY00N+4R1g6ilYUmtAubO
WdLzqx+VQerIPL8ERSPWrp6HmwJ3NyVLQd2d6FVm6iqCysQTx6TjanQgHhSKy8PT
pGP384rDRJbbV4Go7ii7Jeuy7sVlsL7Hd5Tw/JM5tNx2z8aL0SpApSrmKqFYpUWj
6kfSkEfKpHRyFa2XG/kiILtPDiguj6XzTSVt2fSpPpNYWCk040qbXMMTajTq8glm
Wsf0r6GoLBriiCBVBSRdOY8W3Qb1OpislvGluT4lfOOK75EgV6429OKwhvaCS+jI
jSIAv+veGjWGz1Fzx0KGmYGNF6zFzS4osM6LMcQ5tjJUy2zAzmJLcitAwFygULhp
tVNtRODxLw4kumKUFQWGJ0O32xpxqPGi4uqNezlSaLNIbxdgtuBYXbhbJ1nOc6tK
WZHoFTCxzHbupTuT0HsVAK5o2wtbWg/0kZMEWsHGoQDLR4ulpsC5W+OZ38Evfxie
2iLzHVN29qn5RXIl9Y+DLhjImW0GR7tG+/TLJyxq0rMabqoOf2UHKgiYbIBT4W+3
vDlgG3Ky5K1Yl+yeWTujXvwuV+YKvdqwt3KpDM7at6LF1My/icjdqm68hEuo+Wzu
/m476qTz1GDiC+reqKQjN0NRfjdZFg8+/l7yHq7eLpw9oUIgefJ6Xu7ciikh4fY3
He++yN62FUkPGSlp0d1zntUKN87jijI50SqX4IztR92TQKiJXxQCvUITBJq9IzEr
xNMR38vqH01rrOyyljNhbJhowjGm4KOnWBfOmHc0wVnUsQqiImEYyZi2o7cfnlg9
jXX1m7Hs6k9i2LvAf+nQEiaOeUijVBh9GtEsybRrKwFKjoI3usORWdKfUaZ3nBrL
KDqPey3hvTsyjz1S+5iXnPzp2AeoPdcsNaPZZyKWM6qFG3d6QfydomjwC9glpPha
EpMvT5oR1RNZ/CfIdPXrPLEq/0Osipc3BQl/DrWe9xSBJsmQ+OIo+0xiOdKFSTmt
GU4XuqEJbZIwWy15So+5H1oZZ9FSC3xlf4a8HzbhSHyrP0/V/6UPGjoVrpV+5S3K
l8JL+frr0ls6FDjEVMfbTr9/JzKrelAZUpZ0V8qAVit/Vs99oIXz8uzJ6d9cd24E
if5I8lGI4H3RxgtLfnTc+jj2w9lE9UGAUHkMxonSwtwry3Vb5MZawfEONqIWq6wY
UkRURt03TUYazrrriJwun1dEBpLEMRFqlwzmnUCDzmAK/VTQQDWmX4aWVCUEUcGg
EsMuMdRwFVRK7lsjKURcU/rsuHcdWylpSCMFtvpLzDSN9oYhnBA35hjALFFwJL4a
nZZzNJH4RqPj7lV9NtDJA86Q+nijHzXj0UeuxfgByamRjI16SAwyk+KV0V7ZocT+
OnY9DILBGSQFPDocRyin3jAGSgsTO5LN+8Peo7TLbbO61oiPm7rAxVJd3jwjNIJ+
sW26qOo1XawfZ63KHrseJKuW4YEt9PrY3JDz97DLFRRijHARwLVRHIDz0lbxc+Oy
mQhfueitThaBAvzm955ZVNPYwfxf2aCwVf1rnzxE6tew6hjJnG2MnAzwWKwrJ2Og
/LSmuXcxeLiHTmQv55KkPDMdZdSAmTyvRRQ+hY0s4WpmfxnHpYfRx5Waidv5FYwu
Rm7f7J2M/6S/iTXLsrh7nH0NKcDWv11T6MkFfKxlEa6MWBwssZfHqY3xyN9wFh8V
M061m9K1mQbjELxU/1dPVMRwAHmlVOddnX7hpzGbkxk2zo6aBATJchPk8odIqmcQ
ccn0uM1B4eptI+QAnrdV58M0TY7ySG2+M+bruA9TRTGAtR5CqTnWuxbUDYVRb3O8
CG0dRvIGWHs5F7jNX2V7CxA/2M2QOgKjQ64xsZxuWbo62HJQpg5LeNLknw8B4mIN
SeAS9Dv53QLLXtioqNtAO3rdP2s6vcPuwNRML7n2n1k/5M3xPHH/PLyHjcSG6rsR
IOh7Qxi19sFXPsIVfMzVV5oPm5I+W/AxYkA1sJnOkrYLpfrFn9saY8uZ4XzWOupf
A47YrdI/kVCUWenzCYSRRE3EnDY7JlQGnsW7gFYeb8iEfgie/1gMu1pSk8dGSwVp
9X20hMS9mmr+mk27V+GSUweQsyri/jL0vQLju831C4EtcZWHP2vD7R3v4TZoG1dE
DvQpSoYx7zDHF5yuq1JxKJRPHP9IsuRarwSweysnOi+TMwHnb2etzDR4X/kcI9ZE
Qn/ujdpT8ddbKJb/qODZ4ZRvOLYnygR9APJh5G0+bxGxQa+Cxim2VXEIy9GoQBzL
NXiMNlEsJ4XfDP5A0Q59/pyMKI8B6Bh00ILV/D0g4sZDzeRzctoQHVRdRpLbbfYt
PhiwRIkZ0b2oElRY5g6CoM1492XhH9RYzdZN8N7MdXmuEhQBPg6kDDQhcRCbbtJh
/EL1fGHvyuTStWgfONpATT2tG+iZKZ6ImN6vJl//WME8iugRtSNfAzFPFnMrn2uq
Csgc7Ga1tskkJiHECYrxtFbpmFUJhtGCtLpRtJQeh4WhQXaFLZ2IAdF0bdEhN4u2
yt7FjQt3KlX5VjNUJlpNPtET2yqJCuWj0CvSdRPyy5Z44MeSikUG8EOuWyHAu14K
HICSULEH8HKX4wG/r12kU+33n5fQqc0Pr9JYRReu69Oq9fLT9cSlkIAR2y4aabLP
Vs8l69jc17W4s/IBN51tWgfypiJ/hZpqdz4S2kVCl02WZXBQf6pf/lGPX1NpP2a7
hE82x2QlVZPVZxB/YgqftTqhE94wwLuQHpIzYfSTDGjwJEgOifrYrt1K6EA3b9ET
ko3fYoIgSvlO26hjjTQ055l3f7csk8Fd15e31nA800R9+N40+NG9xsS/bORvglKQ
4imffI64sfGw2+yRgw+zQUkCky3EYaYlGo+QL7yYNvo/5vdeeqrrU32UNUsp0o0j
2SXE0B+jhmRNiHI9Moo7qd5fW8GfeB/QzoESrCJZT3tCuNWHIQXBUHUEwwZyrlgB
QUfCqr9LinJ5UPfq1EhkGVsIkF7QS6hj49Xf/K/U9q1FZAtt/7l36w0DJabtgh3x
hctNvEB2QpT8ULVZ/JZncOqYHbZ60NvLf7YAmytgxHaOjlzeqwycf+ycG60s766k
AwnLh2HGERUhEiOHKhzfCT9Bzam6LTubGx3nMi34uFFiQsLCQ0e/t3eEnvs0dxj0
jmLjjYbRm06ay7Gz6T1X0AIsTIdgk0yj8Q3PQm5YEkdYTOrIQRNKQRkdP063a9yD
+T5Ski6Zgnye1POK63c00w6XAgN9MEvIlfIn80DcALQvdd021H2oWRmpfDK7f1WY
n6WHaSWBLuoNEjdR9SHmdlCZYjHwLc+9DhI9Q95PmfNp9xKWndqYp5oS9KnaS/dX
+H4VR8fvkWB3tJy4dzLprhuYzGmM2UqPt/S8UbxZcitAtbcxpYLUjXgG0vV+MhHA
1RbCHrbcEPS+WR4W+yOLnNkmLPKmsyPhCVb7Q1amcNMDgNDNAdmxMO06gQMFw5sC
DGSnn2TJPuCxlKtRa1KRBkqffZGJw0C9p8+SpE/Yj6Vevo9uxGU+R4i2DxyAPpCL
UF3WI7WWx8Pn95aMxexgGWxr7YhLWyVnatFmZjyNgfzVTEbB6vuno/JroPrvBQov
KcTMLU9GxeLCSfJJ+sz+mM0ZweRWpR4UoXnAYEHDpVkAuYHGxxtzlZLqeJlegxih
dYhDopfcozj3ZxuI2VNMJavzVS+E57eCAUcpT5L27O4fqEOfc98Eb1CJ5Hf6a25h
TigT/TICXJlORpof+lJqVdw6u6fX9LJDuy2UM3DL5Ah7r92IPNG1xhezDBvwTDEp
2t7bU/+BF5lKOz8pK9kVBZdFLqG301PtUJktO8iM+oTyTJcrPx5cgShw8cHv9qxX
lmP9RUV/RsjI3MD8lnuWnHncOt+YPSa8MaKHjkL2J9Pvmsqv/P1OczeQyGo/TgkM
2edtcIAG3JfqCJrQ0w3SXFjefPOwAEeAAGcyxQTWSI6FgWwpI3Rs6QTGQ7lzSPoN
ccoXGkKt+rdY1DeGYetmrd+PbD3oMOwmp24bePRb/xktE3uRvzSXUxWnjw6390cu
wf9mYFxDOikzvvRAR5uKH4BGAsM3Myj5zR8Ks2RupZZy/IqHJd8Ks6ZICWxomNEC
gWJFDmiLsiVZ6pznjDGhqgayqgVhbco8zp/FRFm4pmzGkRYtGLajAj0XQsw4OAJE
o2UzRXKWAvstWhbGrsC0hpstBk8kZHOZJOfuWmI4+awdOXZWfqtFObiwtliSJkmv
dOSuJor/qr+KOpGTFiSUeqN0vbhsTq3ElEROyYGdIzOPypfP4O/GRLjJaPSJQmx2
mUX29mFCCK3HVyaZr2EtAz+0zJAcL4eGIrW/7Keg8rft0zoY8Wo9UMOi9wbLCDoS
so8TKpLcBEWAGeRj3xj1AFqJwDDgNZfAelI1dc9cpat1nYmEqCOfglCtL9xsMnZp
kv6aopgVrKhmsNopj8xrCqGr8nUaRpXfEno3INJaqub/c38cO2k4+eJQphmtsxVk
mWgO25fBvXW1UONO0ViMbIQVWK0CltsPpi9V2QLiXqYczIpfhFY2nl8CsxYNptrt
Q4GY2ok9AGzMbKp14vr3WCdnN1EZm2O9mBsS0ePyN/J1Ho9qYjb8nUQdQ4RFewn8
wN3SWDwcxszdauUFMt2sLMwaC4Th0oDzOuF4IsNha/Ne0mnauSPP/Syh9uM2ax/x
/hZtQygnA5jbe/wfVyypHeoaNkCfibWYuiZFJS1liTd+rl2Gg6hUqipq2w5w7hN/
xBQ+/OQunj4xwOSIL7YcUpdG+Vm6xxJ2BEAJv5ilVTeUpx/cqJmDgVuAFAK/LHRt
dlgKvZ1EqBV3fCIXi15/HBuWZAdq/xP48Gc6RmzblcOPbhdUoPkKwt5FW15w5Knh
p3titYA/nCnRdlrsvvsBjulCcfZRdIojcCm+Rjb/yNDL3C5MaOhlxNwMfGXIHaQz
8UECiFEt4n7AafYVcBWEJ1DXRbqrOdm+GlC/qsU5fWAePi4pduqyFsOt5Wp/fN/s
0Hc7gTY77WWVcj6uUP88ba7jU/p2KIL7R+SDBAxWXpCTxnuzyO56le5LBTfyBM2Z
J2HkjvoNpktPOZEM9M99ZzTugIGV4dvpzeqCYR6FWJKFOJ3tsmRJcbVkZ/blaqT+
/NRHKoHqPUB1ZptpVmqsoPDODlVmWR8mOJZj07pPXFu6cbLWvrNVvenwirx3eyEM
TMiJmTKli38Und3Nkjpmzen9Ia5Ylv2Uvgxct4IqXCaCZHaLgLBPI/2vbuEwtttE
zwdGrdTERVTNncq/3HWpCqSr21+zLGSxg960DkCYysvzg9s/zhPy5e7qZDIPDF10
Yb/Gl9ismRMUnOmMxrMC3aPx6ZXE96trKcwMilatp5r+SFc4kj1wMevjaIB2duDj
n+LcZAGXC4Lj1BYw2f3+yF7wFSOlPEaJZ8u9A6duyhcVWef02JydVJaHc7V59PoK
y8kuo4quMRyc1hRLznHcU2ARo8cJSecYvGWADmPCxyP7s7208X+P4WB2CGEY98e3
KwJvHkZyhDeIgYhsqxsghqRRHH7MJxORkdXe4bdWTdfWvcKsKCNfKkISPDA11/oh
VMt+ormozdw5R8FNaD9wsTkLBduv7OnY0neob2wc6Z/4JHLnZO6f6cYBU71QExI5
XLUiHIkX7Px3bvhqtaPBau5w4GYNUC7IM5ZWQxFtzPb0bG3YzRgiTkNi6tyFojC0
miGjNqQ4mxh6QKCkc32lc+b9eJf8cLiGDVNDwYHuFsZ9K4VsWJyZxYT6FTy8lcwI
Neou8FjSNhuhanlOYDfEbxXQ87GsMVeBaKs47eUBqbIb3xDeo5YmtvHg1tidqc6x
z4HUaT74Zx+317RHhPQ1Zm0fGSoYfQqc4sFZxS+UvpW8SzpA3PCo8oNPaj/pSJms
JKY3frEGKp2s0lnjnjSQxR06Z2LLOBR88/+4sh1qPBOaMMTEJtBD6bd/sC2HxE7E
m7GgmjmXEjpGpuBBKliIY9WVyOTU5ThMVRzLtBNNQe1BL70WxL/RrAXq9hNRcjA5
U0K7ZuQZN5OKtW1RsgRlLdC0rUfS18ZErJu0i2FfhR1fq1PkYOWDXRzFtwKNWg59
c4ZenUtHV2PV+8MnIdY37oKlacZpi0nRi8XSLZqjD8Ro12eZk45Mv05Is3YKAXZH
YcM3W7GUN512eyd0onxli2YRz7WJt8xzOBh4rQp7xixJom8Mn9iTVCNduAaCsRty
wKdt5s7Uz3cxawFpeIaKqC4YLyf8lpqO3irEKBTEgfRTWiOKt3ZRqdLGuxGtRuIf
wjsPKeu2VzeSLevqmehqSFMW8bHbU9dZgA6mHFIkz7oAs1IsphLwwqZ2oJzaRCnL
C5ynDQq4ssCZ+jtOHF6U4B6YZsiucCnuu80j7oX8GMGHRSzlBGQbOyxxcOmmO6Up
FD0iwtrVQleiW4nig4+Yigcj6e5UgpLcmcL4c14o7/u2p0xVHg4aaX/hqANjWcR5
bxaDVhaCJS+V7bktys8u5rAMpC7bob1h1zdI/jfhcamTZhfAcuKrjDuz4rEyx4IJ
lwDkyKLS2vcyq2A4m/k8GNOvJ7AKhqjXFUVm1zCAoRK30iTdNtsbaHhwJa1uM7No
dPKdfhMzz8QQfuut4Ygfck41HzWh4tNRJpgCJ+af2TzZxQhiyMBxwoJHq9PLZh8g
1xas5VidmndniFQLhdjAK52sQXUqazvBstWJOu2z/xjjyXqNx9a02aQ32PbP2kpN
ocxyhX9Rimb4FT0BJkfQR4RVl5hoXKViunwFpSu0U+pStP1NURIlAGdV7hfHq8O4
WkgF9+vhf8VUqeNER4dqXnDS6tFAb9X3gCSIyswpN8mZroLKfiTA2MV3I8N1DSrj
ZC2vQu1qbH0iSIUwl1IMhRBHmr5Hc86JkvTC3H3IZT2+M9xRQCSzEVeaUCIkhcq6
7k7dfCn9I2YgPVu8X+goaY/DMu1osc2o//UygG4sGe7MCFV5AupxB1vpwkTRzr5O
iCbJpTzIyzqDbHkHCwiVmTt+vDUVuSap3KmcV04sgz7egKbUgijJlc8uCIy4gIgg
jcbDUMcAzhzx+FKVHdJM7YQTrUnRYhJqf4q3AMvxty17cSvcYxIcXLH77OkV8JWV
KkKxxygkKjUZfiqe8HMrAnUE9SBRhHlKOqBJsB7ej1apioBUQkblxzkTYsslQ8ep
KF8XPU8U3UMJa2nsQ2tU38Ve8uuOI3ezgN1QznPhe5qu6so9V2WnaxJrWpnqVtwR
zvZAjESoB3LftsUnlYsVsyy34UmEOGke9c6TUGTvN9zgYN49WY8lbZvt+4GtZoII
3Fv1oNoM7brP/diQ1PyWwtZ5SaHZEwq9SygZJS9h7IW4fD3JOb5bA8G6rkjM+t0d
2fd/Cor77NmlhDq/+YoWUyrSFHuqiPsb5DmSIhgIyN6JD1ru50fd8SMN3eoF49jZ
Tg6SNw7eUtCztW8h4gEbT4sU3yki4Xr5KnKBd+C3YQEsbStJyNbZeEzPUfinRNvL
KZrHV3ieEWSGSyCLRikFjAe6ccVJd8CNlR8Bf0S+kHeyGfOHstscik4miQSwU+GS
rgg7pAOg9l2je1aCbCzV3+fcRflBu69UnZoaWWOcM7qgqZE/SEjgL9KJn6wNuzoi
ZkE18xzib2GIbRsMbY6P/YBYaBt1kGpsqMPHTyeWpdRmkK+pgB5u0A75AP8hVrKK
umGztjna45dNWda6v6VmSxL1untgAZBGUPNdyOERz2MCcfArpR4EhWsRnYSDJ4gP
n3+JVgUZPVb9YlFGd8cwgxDqpsZD4vPC61CHgObTH1cXSXx9L8/frmi+mpubX2Zz
tPgV9AIevgg8JAU6e2+oivT4zGv84k2Dbfs8RJ2VHYmU28hb2uOJGKlmwq1jNSCB
fT5M9p16r0La33TqGl72m4wIOoYySulcui0QW7UiuOC6t1J6ojqCw/pwIfAe5SJX
4/CEeaBZn4Ie9Jp81AY/CVNWJcrnWbSjeDvHwBkLxpZ7F9amIOU+il4fY6aTVKV7
Djgy0evI5koGpjuo2ZAG2P8bTwOnmoEvZlMeMwilYMIm92q1GC+t+TtXwYixete6
vS5zMtqb5KgGmyh+TEjdbhktWrWEkmKegikdChdt/Hf2Ss8JY8T5jIy/R4MwmZyc
3SzrKtYhsrWx5gU931SVf838EWWKhJONm/HN6yLPgZ533CRSHEo1hSyBB99f/Y9v
aXI/IlmjdbNJJPaix1a+RpxPJwMOuGXXoa/nIKsRc8sypD4lKLLCzjKiJO+gXwWI
JrrqctAhX41EnqWb5arESuMHlRXmXCLb2cWFz2LjYkvOwjhm6x1MDAkMnGfVSiLK
Y1hSfppO9g2jG5V1xdaxtqi5FviqTFthJ+UGxSj4FJ0mB1RbnXjlCKBxQ8MCwYTu
6JpAZYUErY1zwmLrFLmZtgs3BCPoxOr+QcUH93trRIwFQvKyULfzxNvTV9ZX4th3
AojAQLldoQIjXK9eZHqYrWyomwrdl8GGG3IUdfHK2C2zd93JpHG6x5r57NghtZ6j
2iZzdTQeMpfJl9UZDbuaYMKHoT9JxgboJnjd/J7z4W8Q81sfWbIeH6Ir/0129lMX
4aDTpoCnPaCEPMNCHzRp+f18DlY1uimAYAZh/xgUgBH2g/6ru3PmFfTC1cJEGKKP
ZmpZwi4VAOT5oYcXRSWI46U3GHY2Hfshc+2YPNvqFPjIoW2G5TImNkBHlvc2aEru
24mR7mBl/5oV2K1fe3vB0Mjw0ZiO9Rjd3f6bKjXOpxnopAteVj8eThEeHujOQfXb
rQPMelxPTjg03IwMS3x3MM/l38AZ7WZNmA4ave0Sd5+/GxTNUqXYZ7CLraDjDTRf
QA8QAjXfJAtjLwzAtyhTIieK1AnkGreFDSQDb9PEu/aNElAnuTci4hES6SWOgZxv
Yu/C3R99fMNxIYxk7EGqXIXv7ATixW4uYLjhD/O2ZG3TabYnsClwTQRxyArnSqIL
lyS1VpZfjTw/VeTwI7uOJDPzu3EeyrYRlVoI/VZchNV4QMgnfrWHITCBwmPo4XwA
MHUItJdRGZbLhNKJNvlzQKW8Fsf0aAv2idFtZHB7JqwL6giqbzZWkmPs96brITkZ
DvSLvtNpIonyGn4D+UhVg6367E9PXncMxUogXUVYxOUKLgNfqrG2H17zajQf2evO
t+Eo5T/f2BTmYp70ItpfSqa+JISGUv08ztxndnJR+Zlyg76woT/cuE7JfnSpLguX
CJv34fOq8BAvZXdrOmypG0I+OxPuvCiMy8fM8hbbOQOL1XtcAhZ1iRxbZtwsEKUh
6nHMCPVGZhfndpwadikXEmH1RrC3d2YMWrrZ95zW2Tc+1rszYAF24eA72WRy23n6
KFAtxCH/OKm5hXzi+YskxkKGSBvUOcbDq/QCdk6Fj33lPJ9k+SAxh9NEyR+gW+w2
6css45ElG9UmG37OnWt1MBb8SFDNYPMCVvnPYYhF9O/mYbpo//cDz8PldzVahJZT
R8+GNk4h3TIIzECg0vup51RpHZ/Fun4LwtlIOD0oT4cc17pxxUNIF8Eo114RmDin
OtVr7Pdpu9WPRkkD9mJnWutHBz93FxsVRBs3EoQoFtNbDttVs+HStiBV0zfp/+rn
MuaYGZHi2dk4XcO1opfKpjoliBYy7MWFfKwXhSJlFzcptqfv9IEU9sTLqsYhyPax
noDALY9AIQ6yg06K6Z/8BN2WdF0hv2sKb6dTag1b2Wj3sb0rrJOescMD4ITqnvOA
izXvaKmoZH4acwOCgpor713xfuDC3kUyCSm/gwPYXFalH0cLF9Nt4k58Z2JeHWm+
H9/xdTY2viLV+KXuIImXEegxMk44nx59MXNHk9Q2qStyOJuHXjywuBHILvAJNp6Y
6UFQ79MkMr0Tkc8XmBxYMbMV8lJtgul6HuP4bKURFpOGP8EUv5TZYlRgWSbEtCa+
dWJAUNCkaZZM+afk5bzMCfUb70DRcnK4Y+dZekVHS7nWAcxXNjI7kfoZGaExLn8L
s2LnEM22e4izpNUPSb2zDOJtIDKp8jXvmshvzDWTyPerX7kZRVGWbf9sV2SpNMy1
qnTfQVhzF5EHEEqft+y9OaD7akK4QXDAsZsWKH/ZBiBf20T4mFKJxVq5Wcvg9NI2
duSrKC9EnEXhQVubthjL5XHUF7ca/JWnEvzI/Tb5VHDVi5WSX8R/NikXAAneg/x4
YoCe1VKmJGWAmg6Z69zkiTGTy1B+KdwX2gRU0Wb0jO/IjMZo+oAhHdBhrGaYv8ie
fnrBVcLYSwHKPKYv/XVcyQkZC/Qukm4ukjyo0g1iOxjai/EyXOjWiBgTJOMvDYrO
W8TShZzCfhe8MjUYobH54dzPMEmsxMDlqSxSiRYv95OTIRMWfFbMPv6JztiX5VbR
BGE6JzLRgIXuCvAqOogMAgwQJ8NQBdRrelj7341EryqnKMBG4SNPxNQjNUoc2rVq
fqBlL32LQbWGkG/fB2bF0Bs4zTyKC/8qZTdNdYY+UXcTaZwHlqcMm/iPPvMCw8wa
iRLjZGNYLlv1UGfz+NNhnjK4K6irTy3VTmHZ+J+r5DOG9g4lWLUfPAv4091SpFjw
qBTBFfWePeKZlWzFCIMQvaD01caZDnCg2h7FqHoCRAYfapflsqPcWWcKDad2pSIn
7WyGB3HJbE6csA9aTmIiXa3D2s8h99i7hw3S2f0k53+/J4Zwk+6E61KX53AU/Jt8
6QhlGFzNab+0zqIAZ+ztVGB6DOdmxzwTwmNYg4EfwfgO+MwjNkr596ulLEGR+Sr7
57+BY2+yTHQTHS2ZOwfL6pKNOR9Pxk2j41E38ZVnGSyFMmgmuv0ZZUL/it79VQ7D
/cBDOHtpI3FoD1WvhYkKuDHMd4U5PMkbgJw7OAFsBubqJPF6gVfcA57zKNzayXkL
FG/t1n6sVdp93UPtMkmQdLT0YEk5FQ0F8UjuE/ffAyFvnhVc093DVD0cIf5PfSc3
8tLRll4YSGcih8gf+Zbfpkqui96sPjkMbOefNdCr8JM1enHe/ar1/y4xEQ0OOy1V
c6DUUhaCbfcQlGUrGARyFTiitNJsnHMpxJE3xN7vjvDFg+W8I7YpIHGOV4J2UZOo
xcB+NyiLVaSxcaK+yLtFNv0c5CdJOHbsmutyJqbEi53zxD+9VEWJjrWRBWMSv1OG
jCElXXj/gtz4Zh27st0EajyHQ8YsoKsDDtehAUKH6ZNJwv/MKZTK8/HZ/zvHOunX
nwQHAVZ9U9EyxyfLSFtJ6n/uVAV11TAP8SA9G4PawjMD4IM2KudOcCPKI1kbusdA
Q5APENLe+jEaHtFL94NKYXHXWdSZ1TDkaezkACv6N/u2GXwJr8ckDmyYIqkIHKrT
//wUFyIYVjkMPVySlaVVA1LTYHVdbQMIqeUi2+1iJM04xZmkabx50Es6AViQPcYA
5dyA/KhDF5OrcCaPdDEKZqZT1nIgkIXA70AJ+F8EnaJN8jbQo3ckuzNcOQz7RuTs
tOrmwm6HFIiSjE8hXVxI3KH0CjulkYyqwFIEtPBKM4WXlDcU233S1B7Ldk1DFuqb
SPw27G8g8ebhKupks2wHmONCYPplMq120hswlXgttaQJn7By6nAUJmg24o+mXQ/C
MOr2GhjhotIWaeRXXuOrA34zr5tRdnvHXYQOevJrdRpIpTTenLSEb6jG2ju8/9Ss
UtH7yb4g4Smqc2eL2wGRXZGTZnYACykb0ZHS2vMtxUbVEkwQwZw6d+oHbcScb1br
lB6zdSHIgTyuzc0sEzPjxt6+wOActUZm1IHVk3yokA4s+ddVgwloaMazf1aPaOhQ
7SasnKhPZSPvunczuwPT0cmVqLOZW6MRdfM3lSj+UrdVVtWCs5CdWDMbyZ2HfPT7
CVT7K1Pqqd46YbvDvjitfAizll0x15PlTNa6go9FEKkBa64bjZ3eo9PiR8DNuY/u
SbHDujL8DzXRc3o5tBFyMap8CZy/6Rwz4XQII1j7obGaRXGOSgBvYIpD9jamoev7
H9MT371BuaKNrCRN9MdMSbYfpUmhbIQvktdFZrHQyf5pbm+9/NV0q1iT0xyjtlcZ
Lg1pvmmjVuaarPW/SvGVY2Kelo4oy2JnnsjqP1BJw5yupTKO5pjd3khB8xtKpl1Q
HI8u88v7ZSxmAYN8TW071dM8V5Qal41wz5sD3+lB/I5VPSlTUWM6nwnybMmy+eLC
qbEnIFh+QkWuz0+HO70VRDieIs+ch12L4ylnrY7P2ySY/zJG6rvLGqqKrEfEF9/m
H/IW4U5eVsoPRZ1wwxPDPkU2Ifm7ftC/ceeheukTJDblmqTXFEQuq2DLyhNSuyZc
y4EDXYhvVJWY4+lDrr/cMCRBgCEDLBDPbHzBIJrghHC7h69b7Akb9iG9bAU8ao1B
tpaeRf+LhsasUhDZbKOmqN5fPkgN27wHpE+t13C6pqCPYgfwRTtAX5UmXYBK7lH1
U7AzEQCyXv1lR/jiLo+/DTJ2jGRjPeFGJhcR4fvsvY3Tn++7kJ8qGj+2wkEKVjRl
M2ilDVSL8awUZatFqzuksVYREZD9G9TDFcVdqGi6HSo0451/6yq/eBi5kMet9CNQ
gcel8uonapzENjH/9K342rC/3kaCgDrEUGQXZb23/AjvlgLicPw395lMAUkdcwzx
oBzVgsw4BRYoAnBO2liV7UyL4nsZuyrSCcN7iv/DaxP8ZoKvVpSlbdU93BWq/X+f
HBtb6z8eZ91IbDVRz9s0/GjgVslgExckaLJjQdP6y7Cqxm5LMhMhzpqChX/9jVXW
Z7s26LvgQoE23XbYL1EyJwupUJOwh4aFTpGFGY79Zn01SpWD+4dp9CN4B4OonDh0
Xl6VL3O2Y17qhouP8whZH5hIu8JnF6k3XTrwwcIMgDOJI7x98qvCNE62TkQSfspD
tnmE/XDC7DpDhW5IA37tLBYbNlgcT3FvwusIv4L7IHFowD8Qkq7HN5kO1V1jsWZO
sf48acVxFP/1UXOZw5mUqgMnXjs+gcBX5Vgxi75Hk6plajcaDcNp+QwUkDhpnzJo
axgnQ56QedD44l9QmQ22dP+GQone7tht3xKKy4eGyO1pFf1NdBRXTmDRfO/7RreV
U3x2PyXwHKXjXd8ak9Ev6Ofv/ru+BXluFR4BVZ2nZMmvJhkGjlB+UxVIUcRVxIJT
VsBuXyjI+pSI3U1yN5Uk7i5Ih3nW76vTJ0dAma7GIUVfe0DLOV4ldBL/dD68sQs2
HEcjd7QPBRGkv11ZXN1Qzsh4EKiKYJtDBc63eBWko3zEV3o/gH7dOck2CPjg+r4p
793X2zkA5gFb+jPNVXPj4zntl8VXA7ssg8hWOdDlanWg/EbX3SECLSC84f8Oi1k+
J9qaa04PgBHIZ793YURf6uMaON/7EO1yaUYNPy0ZNd2H4dSrjsQdhaIp7mMYR98x
7mm6DJ9r6CrTUgWiHTNlk6uVExK4B3mmXHIz5AMWjYmBCk9ZWv6A096JgsTHeljM
MRyUk0U2M2ygVy4c14vEsz9IxjGPPzTMOjNPmCDOqJgZW1TCYVrfeQRG1gQi9NH9
Cea890rypMgPkzgsqlgg2114tCxMaYGZex2wo4i/fdtm9KQOOc8ePl5bRsd5/mx3
VQk75weTk5pI/hATeT3Oo795SiQgdMZ8875/E0Qre9MWXjlZYNCcYhvOaw8ATj3r
nOJ476LUpG8ANvSFygNleLEGRes1rTltZUBaLBFIZQ1dD1g3UXEi7OIX4dtbyMSV
EavAP3u3RMMdXvu8jaeSbiyGL+gQaKie/20y+0jeQw8gxp/M8A1XhiezaamdirOs
7LDC52N71Y8LS3gjKMJlEg+2ET5RMsf2bO6Jg0VqWiw2m+OvFgwWzFh/NGZVDTme
16CNRAbRCgcLwuCbiUXfGEswGFqST3YapCg4IfE128ucM2myfSuR+xnb7R7mgA9M
7gp4D8m8DvTLhy23S+RseUpuqt6B9kmXsgyjiDRDXfVOpI0TcWvYx3j2aa9KyJP1
phbVxi0Xpt+UlaI17AEWqhzjb8873SxV9l9kTOBlBeEF2EMQV7aWPzvleM7h81cN
dzxgdexYekIfSxBnFUhySg/jma11l3vx43imQP2bEgJiDLx5X88IQqeYaNAuid/i
aA5wt+LMzqb1zTzEav3H1ZQYy2OjPHnw9BDu++S8g9b9nUTduE338mNnIlnQVHVU
7dIEMy3ZuPn/KZoQhQwZqknss4qE/Izlkiz9pkE+PN1sh/EuIemwUmnrFTY2uM1O
FjJBl9HPEcCkjK667gK9mekPTo2fu10Q6/uH3DQloFiv8AxzdsmH1Dpr7PZ+DREN
IgMBp8twTmvvKvktjuKDrI0t2Y0ultmMnQrBcnymWB0WISrVZNZ6kVcpStPYPbZt
EtT9vUnW3og97GooWkgUTfhmcRVB4M6TQe0sHHlTO4dQJ/19NhqZgFYj0JdoZvU5
OJ0fAhMs8nICvQSlkBNgmKfjFL6Q4aEnE4hnuMRHOjYQFVAgDxl5gHlqqlYEXuNi
AfF9LTcqGjzeh2TsQ/vvORD8hBM9mnw+VI4+R4KWR/g9kUZ5OR+Sp0h2vgdRm9cu
XyZ9YJr4+sP+91TENG3cFRLPdI4L97Dj2Ran3W6Fh2Dv6A41/6w9ERGf3107KKq0
qvl0uoHQoMqAfC9jweZ7uoZgIXKZFh4JHrc4Ms96O3QtxTpapcZWI2mGe4lMMfe4
oepLSylv7eyElNYTzGTLiysR51SGL65Co73gbFOzYbOciHgsnwhW+N3iWYfflJld
ugTLTW3XGSYkAqCikC2tur0HaJrwDe1ROfzHDsUwLfk4PBG0g2OAN6PZR4io2tvy
x5JNqB0OGUs+hHbMTiT0hHMKoJ+nFdkoBxfHSVrmAZ8zo9wx5erlJWYv6CwUf7eh
ih6TGVsc3evfYzvxE03oiMflTs7MbdfpgUWF4NDBsSVgvUx2aPJVDRUB71LZjtNj
RHyYsbTICMnRLGLNGxN717iesS58Ulx/Qauht/fA/ARofQu9dpBTDJiLp9jQ8KM0
Uu5QS9YSUZS370IOKu9vCsOCzWIqFLv/5vPQARe4v4zslfYM0puDg2zIcikzm3Ht
Z+ijgiRohQxRHHz+cCBuUIYTCWh+KU5Zmelcgkde1dv3ser+q8S+KBEY4nRMKLsv
sWd1tGBspf5MhlA8JBQy/b3w6eamPtbwjbuZrqyzuGmUQTCrepbKPL7OJMgNDdXs
nsOzgsdLVAI4p87eY+6DxEygdxtALSDj9dhYLRZwT19pMe4puL3WetVwbHKly7jY
zNjxOr5idF1kV4zIMI66PEtaRtYuGFOva922zadFKKz2xOGxXLJvPFoHRlker9Oh
+nElDeOvAYah0crLLPVnWyGMPVd+jOyZF28na6ACyXESQgYtYWccWro/GIY/J6S2
gSlPXBd+tEgu/pOQeb1Xs8+nh8lCrRW1BW1SYPFtRsH5iJBs+8xtZiTTWJ8Lo/wb
MQ+ZPx7XbFdd/rK8a6SOCGraRO+UdlVDYe8ER5dwNn+AreO0ICCSKxVY1gY3ZVMk
44XzpULmZaWLP+ZDnImMMt5c2C6XieqdmAUyti3irt5zU4YgViqa68woS80FJeC2
NlY8yudm2MkwltaHIflfbPLDEJKQdzxmqUvdtuHNZQwLzHpcPkVvXjnpnQdzKKDs
uyYju0Gyj5JwElwHCtXOUvbbhvKBQKPCYDHf0F634TmbfuSc4CNCSQ5rduZZ7/2y
afj54+sI256S0dLliV8q1AGMpeetUIhsItnEVn0ulRy3Tld5+iOIZlEiDsIxQWRs
WgQ0eqggS6A0YapcrsIx3DVIDsSHF+QZcvGLkUn6Y0vYQpROl+kkDQuleFZVaTkd
kEkW61MEHOSBnoxNDR6ZrI1Asen0Tr02+C3kkwiMLqDWZm0HDp2FaE7n7PxWrj/o
RpzjIgdJWXtuBn2/bti4+BBI8lmEhhtKW1YOcP/rTdrE0ub5bRRzVYLWKQQhgP1t
GFvQwBv5op4xVes4dmph9vPKyT25BIN4qQ23CnrEyLFBSzBUlYr3aYZ+h5IZrVbK
B5SYCeOhcm1Dvy1XqatCzo8DY+ipOmjWAqoABZt+WqtpRHKM12v62DHhVnqncMpx
CyXZpJrk+6kMEdoCeOjkI7tjjwEQtA8lhJl36RIL1G5KJMjV02QkzACDn47f6/7w
iUg8dGbwuPPhuvQuVsl7QiopqCevNEVZYVetQcgtii8qSQqW9K8Y8KH5yeZ687zh
yLIPRxP/9lSN1vYw6iRVk/zVh4XSggQQEMLbZ+52wdODoHDixo6Vx7JCH8gDXLoQ
are/QO8/4dG4rT0KVEVRsxBa/LEIma/x/c+rnYSlXtdYx+V8zzXX9xwCbbWoOErI
R0mUSP4ww+nLQu9hPCeCzuhIi7kP4aKN3RpIqGOwPhvTIOml5LzJSGe2rbRHsvYf
BQb9vN0m5/mWiufjb6ypPjY7A59AyvqaYcjwrM+KX/rTyQg8MlgZJwkApgvfMS69
xWicOFmxAOZ1cdz7lGOAFZiamqJoowiUGDKrsJMr4XeQ4oYtOQljh9LTT5g231JI
4C1+vFKDWGWDMxgmkHWDY+VtkDggF3ZTIdX4ROgAebx8E8iC1YF9dimAf2vlzKkD
ENajkZMo/WabaDl6GOYmfeyI2P8+D6v9woJ5RNfdApaKNkS6Vg2H74SZqz2Etqdo
XOgfr2+kul5zVL+DN9b+AQ/28iJTfDf/KZ5NoSs+XeB7LI5MrjaZgCcIGSoa0QFE
mipIgmzsm7/H/7rbcv0+A0vMMK3yKT32gtWeCTOjxV1sMPxPdeQFP2Bu2YqI3s72
A0G47n6hQ85U1M1lSfliXwsTFM6YFpJReW4omRjOG+UKWBjWFEf23rxzFkXqtH/A
a+LktneihXGoWgBUdcrwEjQqp6lc7biTr7lvt07BR2vXfB4dJkWLT+1y+RGgk1Vh
MCsprpjwfb1KY0JnSX9FHEdRumHY+sqfkfP3dCh8rlvown00yrqh/+90BmHqI6fp
AtqHSeDjXGYaTJEkZNGkFwKEwSDYFY+0e+zxUTgsR9eD1oTJuAKmkxSrigk/Rfn6
7J61c77RdIuuMci4SrvkJcjybwduJV36gDYzqkww+dXr+wTksREOxBaXBMfFGlnz
KQ3a6YGdKzeJP0cSnuSARE5TrVffQ23Qhr/dBBUFcYo8Lu5VY6WOJK1BxnWs9hV+
TnVy4j/slntzp6TT8gGYozSQBAFvDYSlVKo+Hj+YPdgzp1WWRrpYA5Ep2H6no53H
kqobQJQURx0VzSZpUOTrGGcLG4PNU3Ku5S5iiSpTr2otyT5p/Zs1MdgzNIa937xQ
gKp+frwrHwzY7S01sxgFPlD/jDy3F8OoawGSY8yfIEVIT/48zIT+1EXu9bNIPFVO
B9ktE2huxpur5T4yJ37BX53/TTmDYqDyW/BPFss/+ysJYhBEbfqZEbkx/ZiePcb9
Whnj9cqQdo5C4YyLg27Z8CiGCYfzTZBvkxkKFSmjmpfkJo6/cegb4bOJYI8lBUVy
qZWEkCc1X+gtG6FsZvPUloWuqCWcR2dUTUb7bLWZjvUusf+P3FBngF1Le6QmT4jU
64abQTD9ciM8DZmzQmpiqh/YwiSK+jEslnAUeApntHdU0FyUIiCGaswyjSGDhErS
vgaMO4lHKOJumdktk6DkO1O290iefnQQP971c3xaCJhvsn58NkCprpVcSTEyzuX/
81vu0dZ6WL6Ey6vlPE3D9SsAUho5rMVZ8+TQFJve5+baKkQo5ZhyCN46KyS2yXY5
W8V5h0sgi49G0EKSQyZBeIbSjdSiiCAZHBN6FnBbIiq6o+rhgES4Jt1IV2fMoiZV
OCgmxXgp+uedVDPXU9S5NOJ4Jm2V4kcPle/wsUOXYnAH0LxRTwL9TIv+yd6R4BNt
WNYPecqMgzJ3zhOqwxjs83fIHO8l4A5kkmwDd0E+F2Ixr7BiSFuf+jLnxaADiMDS
zlhopJMIlVbtb0DTkoQAVWBOALloOg05d3VaEbEL015ji/BqSSzeZRWIaRR3xABe
Mh5DFv5qaZt6xdUpsPUTySIhoYdmgu+Jh4SQXx3g/35M/ehTbeTNpcGHmRzi/+hg
smWPCrFTF9B8+DJY2pgct9g8HL3Den9L8BJUXBtQkFePoP8s6CKXONTod6zfgh4o
RzdDWfd6jyyYDuf+pze6pUiknS/CQIJPu3cTY1XD/mkVT6OlDENSSK9Rk7GEeUPT
9L3WQU2sLy4am7QRtdueW7R2cfQSHMJE5uAycJXtEMNhv/NeCblZxdpL1GjLYing
daIYAiLlhAll4g1aW/GMRNDQ5J97LuSog+WzDmZwpdtBBrEBLrZfoxk7tdEwE2Ut
jGGs/aqWc1pZz3L4wpZpW9odI1gmXX6wc7kiAV/mdGFDFtvxh8BlYUMohUGbC8ve
wp6iXOwDp6xPp4SnHLughH0aG1VgVpqoxuXss9vWMu5bS+J8Q1eCx+oaPbAsR48l
SFJDrMeRJw92xV9ilzlHq0OkWE7C+lrwhA9tywFjxCZqlMShsnLA7PqfduVt6Rti
c3/8JFhy8nykrODIIoZ9V1/7AhEesV0su0IbKM5vooSgN8ORldIWYjg/AHQD3H8X
1cVOXzVLc6+I5D8HTYrXff8lXkuOcv/kX4Tu6F/WrK1QwliA5fAU9T7DN0jx4GQf
hnq5UkILmhPd84XqxgpImjbNvfSBSn5OmndiwDltONkefZLbWj0dWMkwK0BCtuLr
Cwe+2ndbVg+p20tQWaP99miCdLMfeh3OfZfxWtrcMG459f35MoDJeBo5sZC6EbE9
HWTUIbMcxphVVge31s5c6nCNDsj+XiLdMUgI9mR1vvP7XdtYIPW9Bh+z7EVPV61s
kaYSnt4uk5joV34EFhJl7fOfao9z+1EDQ3J+VLZtXhok0DjJ4eihJ8eQG+u1h9gL
w5YRcytXeSWXm0pk5VK9tzlqvoBK0Z6hDlG0pF/sQ+BjwsIJyz5V8ZaYejz9vxMY
Ak3HDT/U32rDpoJVrPTX0fu7tLQ88qsvjSwPKRT4fGSxEVrTEw+N4RH4ZQHb9o1e
n7A/nNu51vN7obJUGxtb7WFlfHhaltVEm/OJLCnAmb31nAU27mfwOBSCpkxKmir1
gGI3NjEeTkL2ZjPffR0lrKtv4hnJjMw4Y36DoiHAQs1+v1xUJwI1FHzcKNY6Fgtx
CM9dOUzGYGabE6JmsKpCEVvJ1DwnSbfPADd2mifYItiS1nllnGqU7GFi8WtjOJ11
0ztQ2/avV0cmDf73jj+OHRv9Fd61LJ197+Q9BDmKvtvTRqbqBaKgTO6B4LRgeUYO
dhWYchdGbfXth7iGUq7gJM8Omf7/Oq6YShKPfmQpJzjNajDGhsViKIUUJQce2Ufl
qXtdZzrbO0Nc2K+/8G25ECmdnCCBJkTlS8mNu/keo8Is3KSDlFbwiVC7SjQiti7k
2Qci9d8ijLgReL6olknx2jVF2/kMdqLIalaje8sL/weH3iz40ZuD3Rcaa0MRAaP8
4YX0QUfQpqnnTBMQWxGtvMu6zNRKrK6JkYP6CbrwTSqH7s2OeTzTwBh0JMsCN1jX
uAXyLzhBvrleQE2MnJJUa9cR0tW26u7QWWOaTQxJCNJ9KycVNCftaQ19tp+sh9g/
PeQoJB0xI7CtnFn/J+L7b/aDtBSZmrSLEue57l65dtcactc8xwu3GYtlEE8hbTsH
kNtLH492JMGSTq7Yp+ZKWnd2Zo+bRamtAkeKuvvdYIQ2Nk++MhXYGbSs941XvhNY
Dsp0pC0ZGCujkRAzKqas5e5nC3cSAhTw7uD8GSgxwnTlbNzxqQrVGOMd0i1GBeDT
a6j1irsBjt/gticMllzk73rEFjWkKU4KZxR1rwDnDzvSNY6C7faF+yXJubieCFtD
2k8A3mP3wMXhSTd/hY/HkDg2afdxQo0vrQTPGHYTxldv8NdBj6sACcp58Mkx6Dei
hXzXY87GFYYC8V5En5Z8H7pMaKYOB+4VBAsEdCj0qDqV9R+X2u7wvHoYcjHxbxG2
rpHlEOyA6+02bdxbdIqa8WDiC8pX4FAaSsNfQ0A7DwPHwCkfoid9/zd+FuCC1mPI
ItAuVOr3vS8B+DkMEgoN5RLr+9yutV6p35qq2ySXlLWRDuCH5G72AyNp/u7k4cmq
dAyaXP3q6N0kCtOlDh7B5E39qsrRxbBVo1JDHwIgQRY/3g9qVhXOs0+75UtU54og
Ct4InaiNp6KvkFCb4nSLg3yylsasdZihm3mAUekRkBVlKNSVsn+Sj/y+5DBJrU2X
wg9aDwR1JA+Z6Q2DBMmeuPRqoDQx5dO4i6dYXoK7VxKtUI8s/t0PHO/rEnfhwV0R
JF2dQyYNGT7k+X7tgg0Bj7yzRaFh1oz0eIvRlKh08/CxMAv2f/mEvui/IeiTX3S5
6AQUB3BqKuZ9r3/PCLb2w13sgCJ4asupuBUfNomdAU74hIeIzmiROps9bLj1ng9u
656oFYcdcQfgJy62/+/6GaWADXU7r4n96iNzMAb1PKw3DdriSPSb3PF4907vIK43
h4PEajjp++7X7Goq3ZgaYH94R2MIbrtT6MtI7Nrl7rBtr4WSNsKMnacEoXGgkmwQ
Z2YlpSsE2wIvwr5yDCvMCpdI2bXeQR7NHvR0l0xLMGuSV9S2YJUr0ilWhBzs4Giu
0GrJEMpEhZmEnAGRmS8T2McYC4pDjeDAdIPzoBlCWX4S0UC0EyFo4tixuPPMOzNG
TRCzPchHM+fux9yuRst/0gENATfAHTzKDAAMcm0IKuVJ78OUuWGgLLPw8gDQY5zu
zVz2zscoSrn9oLGnWcmEjAOPw4TZSTPzSbT5/61XrBWQIV3745sojEwpzpOj1Uml
O/jnc2v0VeTpRbIFlsVEcgG9KcTAiq6jOh2kpYtHHy7AaqnGQwlfSH01bPMBHHGa
7risXWg6VgOUr5+P6PGLipKpK6SE0WDlPN9xof19EuVFtknFRSaAoR6dQfd9Y+dK
PH21FkSLjrcniqRWyJ64vnzv7XITjm0Tj9sm6zd9hh25NFE4xiHpyPUCUfbG9mWo
BFg97lc5sNLQAFNZisW/CZ5xDfF8DHZP0cyh/bYygWUjVqx7ppXGcTdhaVKLx+h4
2Hqwf1+BwKD7A5hvWXjLzaZhCt8FyRjcjA/pFlW9wmzylNrXC03e5rXG+VuDf7U/
IGu5cXVxVXaK7YpV2Ri+bcGFDNtvz+WbdAui5DExQiiDF2oTM2NUVRVmPC281UXd
beZhDlAUul6mMuSJKIum9G29zg0UMjdrdyWbtFGvdwv6MMGWQK7SKqh7Yj9n0ip1
K5qEoyMOezLadheTtNJZcIq0DhZMQwNi9uFpk3+5q4jyiz1xjwr5RLLHGoiJ0svU
uEPWQD9PvLrxKqAM/qXY5h9yjqYtWAZ9vzsjXUn36FceqKGuzbAW7gbpcNq2oTDJ
2RsLusrSO3G1id4rC/psMyrDT0ocJGwSscl7pSvXSLS3nlh1QQWu1b3nzC7YHLnc
TA7QKoTWwH1OjOe4xtNi6V8leTdImUIldMjFDp5fmhzshQA67BtWUoXDuS4TM8WW
VqvN5QbyuvNX/kFLZn8IFonW8zPRP3l92UiL/xSuzk/3Sp07/PNlPM1bADCS2wfS
6DAYG+7gXumDaijQYTfAqrhlItOG2IGbQBzbYaNr7LMMpPZT2sS7VC8if6uLMm10
YPl7FrzgRPVzgz3FMiCz6loFqKdrzrY4XwXuifHQQGpGsEA02RxMxLdqaJMadl3k
NPCWZXXQeTnLNf2TTbkGF5KVYr5Ty8oP9inJMyfdjHMALWCkng9wpRnNdAgscZvQ
76fYLOcKsTIXDYT3KyY4z/tIjEgAmdhhcFBtSfIlTt0OOWr4KBIZlNqdYRVoG2V9
5wBpjnNRy7RVj3KQDihf/8it5vbeRNbvmhqO8VJupg4Je3VPTUFrsrdU8J6IpPF4
YbPb8F4Iz4tO1FYbKU7Iq+KSLGlVLXHnNbJwp3Ld35mg3PRGyVN1tHLkhP99QJZ0
HlCIKIWPcuM8XvO3qYY591IsMiwptezAAWKbI6V1OgGFUGGLcKkNgKAbkaATcbaK
X4AWl3PhPssEBa/kKYTYyRX/abF47AeQ6C/h2PSYryknNavbmvmeWuOY8J6eRxHJ
HiRr3S3IGYqVF3eR++hviTb2F8ArfHmI1f0JUsT/AU6A8XSjYpiFUepB82ZPuEc5
5iIyUm9sH4Gszep0LAVnSSmnAUanKQPFJGvrWyBJvVwsXgyZPL8m4GPuAwKAKBvJ
S2zgH8qc+CPppHCsVmlnqubvldnYVFyaoVZOJo273tb42IuXSsKuRoETTpcIGawd
4a8oBAcSsskHEppYOwsfyMQMs1P7E8EAjTgPS8P8gcy8hy8BkYN/D+/7ysQUNfPD
MYDgrE5bkWdHQoE7TnpcmJk1D8iPqYwR0OHlTHXq17vcMCGJ7Sud8aWNnTtzagmV
Gsa3QglH9iXD25Rad9+bD9DxkPPJW0Cc24SGdkcvlYlH/KIBirLyInGcKWENjru8
Wr9AXs90ApFLhvdzU4ADzkmwhLQG5mcrug7UeKoZzNfYWHKQG5yykqBr61rkTlst
YIubXG6QDtfHgokYblznrHJGX4jrAAsnWnxOYAscxjHhyezgXPlwF5/kwXhmwwRU
OjWw/YMF5fLlcaXBHmeNyBeV2/+MbinZ9oouvE7JVyv6XMCTN3RpeuEu9IlU6FU7
bjO+kSA8CYVLZd/oh9KBWgngqmXkwAUidAo0GQwSLFZ3pPTxiZd4SfjNCuyxLQbf
S7CtHWWt7DfazR98Sn14P7lME44XgkC8cjSk/jd9amV3Uo2EsGQDUhEttyY35fDi
+wpszF78vueI/M45l7Mjolf9dLIF991iPxFgNe1kmCu33cQECYcu2W/PWBDrun6G
mDi/oAOO4X80goJ8/S4oWT/fRy7RN4q+sDGWA6hedZq8LEU3Xbv3moxc4j6CUXIr
aL885iFrsYK9skuctPQHoUVAN4pPY7evBPLOam+R4znLbstSaBR8X+8nvduK4UKe
4XtmGT3ZSO0JAFxKQ5+M2kNVzd1fEhyoIrVoBjlUQO7UqZtcaxCBra/cIp29NByh
DqJk/3Qo27cNx4Dlcotqiw5w1gzAAqqGO8MimcGPffGR6VI8C4zxLmtV+HU7MmK5
y/TB496bJ+S9tahbuIjFD9ki3VxDAjavpQvDG6pBTsTfoezkcREtmGMxXddM38IK
jIw4S/VAPzENEtphIwGT4CaR16EGRqs11XAOOyZENM8l34C7PZHK1Mx116jVh40z
O7HdipwOjy9sauPXogRabFcr20FFGRfPGSY0kGjUhxhURyAp3gEIrylo7RvnZa27
yr7Zh7rVb21KAK6xT8YoKQ+6S6/RBVxYamQ3uD7mIhYgaYNtrbUz3OJKYS/A2KV6
odo8hczWulU1ecuZ/O9SR6OGvDdBZREiZ4rUIXYOoIA6IimBuudl0UgszITnqp1d
Yzp1j9VX+xRH6CrtdH6gmSe7sdyX02m88fM/95nleG94eB+01jfYDd1LGfBBkmIg
v6rtHbSMcMwUOCHE4NphGxoaWi20Oc6m16Emje06tMKKuXcQzA2Mfb8ON8+O2CXG
tolHbPQgW+513pOcwDIVu2g0wjN9q6SIB5dAAFzUbQCZXDzrNBVVW1M74YSO9v8/
c9KFS989lWnMqFL7GpEyQSsRILgYgi808d32ue/QXPWAYTFfEXAx1AXB9/yYZmcP
Rl3+p7Z1YQXxFlwJaTI4eGBfE8++F3NSihjQCQutuGmmmgsFlNlbXHnDigYiKPM/
H1VtvugRW/L/nM22AhDuZ5LYoAEtRF93gNtY+cQj/YcesZRSPvlh3rFKcAS41dA/
0BsGNCxfbskIx26SG6zedQ6azuBp11ZVkk3A/7pLf7tjOZmRcdhud+YqLSZ2O5DS
pg5LHwA1LYtlAblRgoN/J0SIdd9scLZsHPBAxrH+qi1Tl7KKTMI93k969mYfn2A0
3fl2wPuHGJyqxb3B5wqDwm/A3JxHMHf4ods4i0IjFrPDhLfDcFG+G0+ubpFQi/6w
T9zFfp/PTld406ETF8jQ2+MWp7nzdEPx94ucBao4uozRTkLO6sNdJEtHglw2yqbP
sZG8OL2yHZr2VTQJchfb526Mpy1Er4wd2YqenSoRbFoyzkk3Svr7PoDY9tivmB6h
81Zth5UFFD69hP6LSJead7L2fDirYJ2fk9MOCxEq8e2EhA6lL2tDG9oE4IQLrg6A
ZkYZ7poxT6AbzMQ7MG8hGwSjGUwAmtKprFcZgBr2IV2VtIYIcsVIgfele8Om/8We
FzzGJq7loZVo1hRiGMrrQ11peugi2PftCAxGcUCM136htc8Iri3dP65Z/mUgh9+/
G0pGR4tSzQa+fh1LLhqBjikZOrzlIHh7EFUT+gi+bwzrzfZ5b5MEsQBO9KWlnjy9
YZVXpscGbJVz9FxPmHuUPLz3kTb3eLqT2WJISkDJUg7JLYfMCnVHfNSV4bU6AppJ
hLEtowK1XnAhJJB7QcJlqo4JNsth9NYC2/dE6Oejt6HSJ5DViY5FyCEmPuxbbP2B
r2edznov557mEhmfk5wUro2GU16xvmXwHFdneXXuGu28v687DIsmBwvu73GmiHpT
G88zmGPEdRHBObVxFd+gfc/xj2uGiWMir3tVoAIL/lHsBj7KSfIgrKPVgVhZ+Jh2
5PQ/q+CofbSHLBN+pMA+DmEiMGULBslaueRhX4fqTdNptzFm1uDlr/uTomi2pmPU
MOUGciGZdUHrRNfE/mVT2zA5WeLqPnbmnlBgOcJ+QOR5mKDbzusA4+500qAuBLyF
aHFD+K9riRvY2CZnaW/9AV0y4HhreN4AaOKNhPqGditf2E9dEfpt/ewFUC8K8TuB
BCK6ZUe9DVqESK5ZYXUwgOUEay0c6HqDz+6T5lGIpQKcd90Xw4Pz3p9NgDo8X9+m
+o7Ucjl7FkBUZvxVv51xXFfEGnJZ/cCQxmXB2+or8MgfxoB6RFmRFy9gefivhCnG
Mqml6lqjOZKB9p/WHt5cr9xjvdauHt/niYuiCwDK/T23tJN/R57FIuHG2qq+dR4t
vKSfmgfRnGvw3fwoCVFPAflsypmu5HsFbXcfXNnPNPzSRO9OftBj9i1mUn/ft3px
bTSqdj+JdVr83yxlj2Dpgnw4L7rvtnDJSOr8nbUpBcQ4cUc6vxrAjeW8FXXdJV0b
mQ2R65I8cInIbAnDi5W2eg==
`pragma protect end_protected
