// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Rxy8DOvNqmsGWc+o7oMYb7Z1JxmtSMcUtFDPhgd0fqCYR37TfRXZyQUyymCbXpxod/7XFuVdOtuB
rMCqILlf9QkIPAUVZODpX+FELzL3ZMkdQpuYQLR33cJCH3A/pvdCO+CbIA/zD/qyJzZMXHAh0zzT
rRE8K0zu1ZWbJgCaeHjZrs05BiNxiAKsV0AkVTAZpkbdlpQMQS0kI6UcthpawRgp6Zj98ykc/KC7
CBf5GY1XcxtdU0pb+jMZ1tidUKA2y3hI1XRLiMiTTXTKOtM9MChTrNSSuFdlFEm2EGhxOCAMCObe
gWJ5QjDZE5lGWTXqgDiqdZLDBGgEjeopvsYS5Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
YDAvTeixWkMUx4Y3tjjtzHZpVIyu7D/m3rF7Y0jDUlNKWmR1OSbJufQLmokkUXXugxIReP5rj7w7
o8ZwHqbOQbEsSu5+uZiCQ0078sWCQJibgQsRHONDLE9KuyAfWPaA7L2wXhSzWHTqEczWctm3bgZE
cGciuAHXaJ+2Hzgc0fk5YrmyoP2oK1nh050bTvjy3114VH6PgeRQZ4SFIQfNY+AGlLXLSSt5WcD5
GdN9PzRqxQVXUPfM+UIsDEtzodmS3aAtDnWw9iONqPcBh1abn8z7K/5e/0UEoTCbVMBTf8HHLzvl
hJKKYvTA7fOFS7f+rL+gNMrU/EPVOZuDFBvs1Ov/zbonJWTyi49zDr4rnPuo8PhgYW7dQiw0VwWb
0zA0LhkQ47cMZS5i8MvBmNF9D19r1ml5o5wd0mU9P+N5L0csjHaugiI6SPmi90Mw0cHEIZpcG3/l
xYQsHKA1miUj4w/xPGo+37N7CWYOgHLVuFkuQ008vOmocZ41Ks3d7ZYZZA2BYyCXqYJ1GeZsIvv3
BxbiHtWV7O0suawnzBiynr6c9mLRk77bAva04CD3AA7t3XRPJ4kaNVsczyvtSppyjva0hPVZKato
KjuxpbbVwnbKtZiLQqw9/EO8FqRe3YKkdgXriSmFuE12OXSJrWGLgSeNeBDA8BexDqJ4zCph4vKY
Y3Kl8zsbHHxkd5FGg4WO5qhUDqs/Fb6NmbY2FUBdmCJzm5qM4hgcCj6e8I8j9TXfxNzx5LLTr1rW
/UVjF3BF9uYe5Hozm2lU6BllZY1s1pRTOcfra3TPr7R/Ddinb3V32t/ZTJRIQ9K5UMuio8vGtwDy
Bol8THM5oUmnjtblb0U0YfJaKV/u0HWEdfpy+cOIzGUIVMZC51gZpNrJA71J9OXt2sJ5Lsc7dcqZ
JwiIlClSEN2Ptj5GKWchMBWsufkRBfGkQjDYdCfq1bjxZfa4/tCvUSkOU03nzAOSOvTr4i6YMbVc
t8Hf1WYILDoIHgxR/1bcIFMIKtE7HLB1eSLjgHeKyjNqcosFj3DLt2DqgpIh7cmxO5ISZS/NknWh
EXaBEux8Lf1xh3dv1JeAh+rwh/6/NuwO6DDfkQyP8DrRqhX7dlFG9R+NQxGT10w9bc9UqVWHyf+n
eK1C27PuAS31wak/T1TDThlEfAA0wcTf7GaQviqkhzze7Tp8YHHxQiNhSSGRO6hJ9rpI1kQ0Sad0
WEv5+B6yBX3sDkiPiCvFcKyhLptAyMevaajiYCIpDFaX+w2LG/zTbp3NaCCxS51gSLHkt2aZtIVE
3o/LwZ8ROaJMMOBDgJKeQGg4pbBJ04vPWKx3+hMtUNOfuRcnqn8dwWXvwKAs+dW0NdLidVatypfQ
BYUwLI7ZgIY8uUGDMHGMj2ZL9Ovy5cAP1CxOwtmQltuiCZno3OPVgwvRuuYX+uWkU09VizEVv+QW
cfH8MsaChQM+e2kK8RXUbX5e89PDyajrmGvfOsZyQ3CzbVrSHHKmjT3Mc3e5KCQhkCEzFOvgV1n+
her6Dj7w6rHS2I78hUD+n/WlnL09yuB+5BHgMoIrgMcm/NHbVXzvVUE2GtbJuCGccf8wksefwHRS
7IFUMJQtkYBa6X8sW3YT4H5nsNURwEWpoltt/xvOTy7g/DUAWUz6HzhRzY5IMSSfDjZipuhFE7Py
CoeLYtGaFBTMX9wRiCCOTHNPrYj1saeMGj1GaUNeDsL3owxtaaiuXlmLJr/NE8fNcMGROdqB67X0
l/6L7T+uWI7Jk4mtYkgWUBT4UG8yGBQZ+h/AlBR0/pCvrC6VIU0HoyxUeLkvAy06CdrH9RSESVwC
WwzJYV5DcO9tKDIVJ6sW3vDpH+xJ7OIK/Q37ZlMhn4m9+jHj3MDfMEqVEHhd5lC/Yv6asF0Fadg6
sP6V0Yelbam63B7kl8QipS0b3EF5jXAa/VUtPumZqMlkXBVYW8CpnQW+hrTMmE25R3/bvEqeIUmG
Ojrlwvvl9xgA8p3Mf2b7DDq9MxN1LayaxF0uDLR4cwowrknVzYv+dCWBcSM0Y8hmHNhv9tpHD5Hi
6NHMKjSPvVV2RJnJ+ThcpamY7l/3DFLRsUw5ZC5rzJgCInmzWQXmXRNrMv0TTeD3pSogoKTmh8oF
4MY/UV0mNBD4eIqySB0JB7w4rsd2xw/43OUmLkgFg75y+/t3wOmJKtGMSSUUUQ+tL/DaHMAQTQoD
TmW4zaBOQMTh8cGopIIwNn+F/NEMNrqVf8mVnpvQy9wjon7abM58E0UAKz6hL3d67JwW/7RiDREW
3KEHeRUho1T5q4w0tIFYo5F5MNQVMK0CcE5W48YOolxkZXk471C6CApaWYc7oLV7gTaS0KnVOKBY
eNaCYxnNwf5aSwp+eEniLAlpt0UPJXUm3KEMyz9W7L6YMSEOfas5Yh4fTyqBDy7Z9KhsvYgS799/
Wvk64e5TqacnTqfxPb/UxhoPYzdie9FzITTkJ/4Na9JCpB2Kuo00GyC7ltd3sx6OjXAiG0AduFQW
AwA5BzIdxFNqUTVbqsi05Y6u6VWNjgOLE0mI0M4t9TkH7aEmtLIemwkuJt71T133bO2+K0613Enr
9Y3yg6sos6xPSMW5QIIzL+x7CvmQ62EP0m0RVdmIAiJka+B2UEQxsPsBBvCvKqGlXTCH4yAgplrK
ViDDmBu2IWPHU3j1/d8ztaKerSP4jv1GrwR+w/meoy/Y9DWEaZ7s7PoOjoMb3bjtvnMJ2hj/jM7D
BX0+m3Ce2LdAF+VOqeKCgSRKF7d1brHVob96BRxkS9IaUOG6o2zhrkBe76BO0PP3qheWcOIpbe4E
ACNS6v0I6IMkiTcbHHXlSrVGMGzujjAjWTOK6UDOuynNxllk2Bkf1Tr2JyTZkLPJGKdMgCanw29W
xxQQ7oYhIfU35aIIdCL4ICJoDQkGrlcf1OCS7eYe+JtHeAzyc3BhtJm0trS1lg3zsX+2/2TFuJzk
yjp3nS5mHWwoTtfSIrl2h8+MDw64i4K157rROBV19CrvXl4BmJCW+I3RBFv+SYn2d+w0BHVrr53J
YwIDFqQxN58JYLUeOwPCLMrgDCiPlvDmbX846v1VNohDvok7TcQB2SwvSV4sdB5pXK1Hmipzz67J
ggf3AbRFQPif1bZmkVIo/d5SPLNneoFSpDe9937OA89GrMP3RHh1bk1nT3QfRMOnfE+25b8kXhmJ
dhbZuLfTIEMlKttBQK3lBaGkPbrc9t+4+AlzfJ01wEU4v2NcolGQE5Us0cajdWsEgh6xaQJzKlmf
M5m29Bl0s90eXbo6n18v04ZJ90qGRf96Oh5W06ioMNWEuFUmWjXuL4YW7MYHJrRTLpN4ZNd77Jxn
LhqKtsLl42n+Jfw+g+ncq34V8aWd1YNsQ4La4KG/AL8RgfEysf92jEir7Sez/DJ6Wndw8nd07Mun
z+dd7qFIN100z2uxDG7h/QXxX+YPXA7S40fkD7xZiHFdSRyOSgiPb990LC555Ym912+utDsGQnSC
VCnvcgK0akihMFunxv4kwAn+5PpXpOBjKcNsI1wdcxVBxbqzjyWPrjIcsqXF4CegMtVRpZBWlRw1
rU+zXbMUuLXte/JD4nYl7xm0+SCa4mNlnbAeDg9D6lP/a62PwX0gMT33kjKax//83I0DXrGarjKx
OqoBZhHDEeU7ToYAA2eimtEsH6dg5ir/8cevN6Qp51N4V+4pp02VKukSBESVnAMLKouCwtT2Xul4
SYOaJd5HRIR8EbmiQnO8fanxIRLrqIRtjfziNf3RjkjWtzELDIJ44QAbfUCACDwCh03tctejNwaX
9U+aZBLXZXXAqYHJ7EqqFzsYshl0hXGjwN4aYLPHNnwfMgSIyMS0cw77IFshUFVesovinwOdPf/y
GobihlH7NYlzE9JTgj7dW6sIUEW+lckFW6nZz8cZD6sjKEoeInODId9AQD+Tcpr3zfC315DJ39d0
anHZd4k1zA+uy6VNaiJVw398sLWoJ/kAc+g3nxhv1jRxKQnFlRv67M496Ulq5KbuGZcFJyE7HJs/
B6M/841OAgvmRZr2aI3iayIUSON8vL4HJgTQka62AxaEVVkEMOKW4gcCDBB2J8LKecHGcEJXXLF7
EaSvFQNyna5skbnXFqoZ17UcfCQrQBxtVKGkOoOAF8ZVRFKjkSsPJOrdgFtot+bRH3Dj12m0qdx+
F4LI/NwMhHM7lPyrfQ3Mgg4ZWtjmh/NZC7KVOeMYjdE78lDtIC5un5JRylF6aw1wvXvjOVN4TVQd
u2BMCa5CiceZ2o1X8BEsEss68B2ik26fw59P8n/Ng0gy/yE3sFKkWx5nnrrj7ibtFplUN2cFR6pq
0clULYRmVKYV1w7ghHOccavbVqqlbvEwRMlecAgeWnzTReNpEPingMZXHCo1r3q+q+fkWah5OLpG
EatkrR/Lyn2H0W9MUmmiu4rlZ2XdRXnJjfkuLzz65qmPOlZ6N6lk9qzUtWL7m/T3VaX3rp4v+EFR
cwEUX9ueLFn/7QFipa4PMpeBOYYuIBqDmQi477iqhm/OHlu6y/hGggfKz5QhC/8Qgd3makfC07vz
6DnM6Gw/6cu20QNfODiv6bD1dI5Kw7hhZ7JOTJsfY7GHp5IiURS2J6awTlcWmlFKyh6JTBgSRPrQ
UiufRlYq63gX47nuOenXE2PtLDVBF8LBLpEsN1ODemp0BUdLAd1v21MDrWh8e0DwmP3AeDdlVPNP
E7MBSdqUP6DhvCibmJL58XyMeyWzlp0iTFDTazmCZEwVJz6wB4HtTla4MN8THCgLVTlmLz16Gn6N
fEztxzmZEI30xnpByWDezqwzoOGovD5EGJ92LSrqdiZfNxZ+klALyFkwSYUbej4dWqtXZ7+IIc6K
Qtzzyiz0A9Om0d+VwLdOgR+uHxtkRa3erxwuzSXsbFZ5uME7PZZequIiVz5FMXgIfAiSw1bhL5Ad
X6mIfaIIyGnYWoz/WT9JBaHA1fd0OwudcrEKQFlYTvblzXfsb87r+fyUsCNOFJDSaHTDSho9q4qX
ZBzyhhw3TdQOUgHHPyJ5Ak5Et+CSxyWxlUm9Usmd/ebOOFeTWZz4W4N09jztiL//IE3Qm1FyaWlF
okhxibpDuW9vzh1GcFOVgLH3y5zTfjflWf4EsDwEt4jLYbj5jIkgMnxmHhG3souOm66TssJF+oEA
aZormXVYLBSc5d12PrQ5EoTW0F+/Kpj24qHskQ5mBEupN6IF/fQh5xTfF2/OK36/FCUa1qCz2xj+
P7am+8z4a4H8qv5Vt2HqyrT8382dP/y5ok5s7NM4fNdkOo1c8CaFPZ/D7kPRyaJUzBtKL5kCiwds
d1SwcItmpwsQAO6llXGGb1u+yoUlBf9bmB0gGBaiDDgZjpZSr0b4hO1r/1VNmWi6484V10OqSQBP
CTSTbM3nQK63zzky6pXZeNPeudgvxnnyiW+Nc21RDdtimIXkVORU6BKAUOspe8UnG/pbM1f7mCZH
5ajgj8LbiQ6jzp0BMcIzgzxidJdoiRTXYsccvdyXa0AjIN+e5O1N48TM1z/ZYxGWIp55Zk3OLMTc
4bjvuLruWzgg9B8KP0Z1QuqJhnujG1J3/+lil3JoYEq2mgihtmqJeK2nMxAInU5SaD8ZWMy/bk9t
nWB9XF1hsviwF9jru2uvxHBOfO0E0adUvfYcLro8QoojHeldfwF0oMfll67mmdr/YkRngT6CA0a4
fqjr8bX7qk8G7Fq2f/NG/yBSBncBAPQ+Ezc7mAX/4PuX9kS5Bhc+TYY9D5aHpVp4NBHbkcPS/0D9
aGqAhwHMvQ5s/ERHnmhzREI5tTi/0SumlQfZg68Rws4hVoqWkaK8iRH7dJIwKKodSJFXyIJAEdPq
lwaUzuJ1Af9k8iYnkTH6LuWUI1ShMgzhkbmju2g+N6l1iCUfDc5oUMWUUuhowOamlE75vJncjA9T
FM15ddLlybx/EjfebMJNuNIll4zYcC5+q6Z2gYkf95rpZzckchPhR+9ENPurmU+KUA4ceU/++96A
GsKYnVWnPO67dkzmU7NZ8Rb6R+E1/z7vR1Y6LAxSs0NMKkjl8jciJoRX2G4q09VoxutdZs86u2A1
PrkMDbNT4EfmX26WAUgVKp6v/wLPWzPzlE0EaMBDBfJwL4YVLINZOMV3mkqvdrL1Qa8uGsYdxpqF
HuzMdS7ZdbNJN8wNmgy47X5b0amCBp3WRFts2SI+oK8FOP2TaUeRw9x6fhdCb65LfGhrTdDonxmA
4YrO2iTLMbh7gry9L66CQ7ohuV1dXb9Tzt3eYOARwEnmOZAmgTogLUknTIM+yprfXVT4zlMYM6DO
Jq+yozo0aj9UcDhNTvQ3v0OdxrVCbsyX9JruTrQHAVIb/NHVLlHpq1sT8snMvxssSyRu4k6FrlD/
E4HyAbatNswIvGI1XtIxsrUQ6DZA9fxxcCUgpSMbwXWTvUfFj+JRnoFzwLIymFfmcQCMqT/taJnF
wFVVlNjfSOHn0JIr4vzBNmILh+xJvLTSke/szY0Xpr+7iECryt7PrrF24k950CSPKlCBMLzCF0Y1
SNsPIIIncsVuD8EhHoRFbNVcJkgurGqzSuPgy087o5ZhBf2ChBY5KexvUkFZdZj007pkez20WZ3R
RavVMe8wxNKdxHoFNaOwpQItKkdksSvOIE0eM4gZ2oEsTvHzEiwbBopCj/WzB0GJO3UWSjvjnJej
TgW+HUM5uB6tdwg2FShPkgRwHM86Gb/RoONspcQNcaMFefnYPUBecZEYzBlR8BpDF+xLVVGtXp9D
dy3DMRtMRedO1V/7YfKBlgVpMBU2VAvjwEyU8WamQHv5nI4Vnyins2HzhDsQJTfnYvxSZHcqDT13
Mfvt1IA+P87A3HrB3qwgAbCP2VAvnjGsl28bxJkfmKGU+TaQNE1QHLMUjAvRlL8tQWbyhNtxQj96
uMVukQtO6H9xa73Xxkd9uxaYULrxxeF2XGip78Cp2OBNBEemLgplXtLtD4ZQrGDG4vZfG6i8asAj
p02ksfM7MTZrCl1QcCaRhfSV1XbaMDKslDgaZG7mMXBLWTCBKGcQrSX/MDYF63SDMG0xntAoCyo5
ytj31V0llCjx9JXlWvZnn1NG4oPCSsP+u/uW1As/LQcBSQF0G+wnZdPeEP4m+XEz/Ovg5syNVdMW
9dyWuruE1d8VU/+Rm1nqJTat1iIN+GETFZgD/ffwLiHZwjudJFyz6OKRH9e1tIuRvSjIT6SBf6hC
aRhiAcodkFN1HDyT+85eb0jIXiQuzvhUck+a+XJCnhWwPHbLlWzNwmcJYVUno7F8fD5VC1lxvlbK
2Ep6G6GBzAEsEiJBZYYjXsLySrSt8pC/dz0KWHqSNvpua1MYfPslItIPr7FV0s0sv2j8Y5AX1Guu
gEiG0ezLcbp/S6bm8Pt0U+g9etChyrPlWY6zf6PFk7WXPd+2kX5cYtee2SSSU9IXv6Tsg/2/Cd7A
ZNclBXATLVr6IeUBiabK/zpox/GLXBQjptqUfKqKYQVKvN8HjX4tEuGDTy7fxUw+X7AhEaPgSMZL
o1098C6dCqjGK8S9gRziTDd3OzBE9MJsZBJ6kM8YzUtV6txbF8QO0oYN70PcZfSFnf5fSTU93Ali
67rNw9dnK3utullbutFAqP+PZYnV/fiZRbch4COpuqyJtGgfYlLLkYhpajrzbQ8/sFxb1TQ2ccku
cCk7io/71L+9Ovujp7kyOHuuIjBL9SGn9hBTNv984qURXO1k/2duKjK5B4siWb/p8AIRYWQIIPAW
Yhu4eE/M4sV1Cq/fVRUkYOX/ILCBughsNBr7EethXwTsdvKIoOLqioHEYRqfGIDK6b0W7yA0ywGA
25zmvX4NaMHOa4W43ivgQwbSbMsPcfnEnti6pwLUZYnb6/JX1LJZB0ULbQ48RRKKyZylCxZztlMc
1A6U++y5eMPc8gs9Kffn2ob3qXzWs4xwh6XIunCg2eQSQvx6I48oszNeLJMs8gIepwiNzNF2IEZd
PwTyFQ1SO1IYQDde6MTMpTjRqqtgirgovm97qT6y1dg+b/VYRv7sAZmFkCiYl+LxpZR1IlGPNpuy
FSAQtI02xc60udRjXZowpwsk1ZNrQ8eta6+JAYpSwIEp2nrbJuBg1F5KlNdGTHojNd4XCZlH
`pragma protect end_protected
