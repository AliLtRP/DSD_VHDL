// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OwcBA6a3a7qSitWMp5NxGnP/wTShkUP8zXv+L/zPvbutDIi8ipftfCjHybaY6d9V
E+l8hbAj9/dfhTRSEsoNZ3sssmWvMucLcsKYLsKsBcZa4FRuoDKNEp91ezMmQFM9
7yHqhqsP3qPYqVuPTcWCfFSvl2TaFYdlg7y8LL8iaW0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11296)
SuPrIkYfuEEaxnXQJ1nEPTbX1wt2qauTK4krBwFo+1oqN4y/cd2aRiPKCbzHvJ1i
QJj8qJqpgn/cItzbJvif45Wd3DzX2OLLREWGEcgHsMMHvNubuyrtiG4J3j+aOYYi
cJdVnWuDGVNUjJpLNYJw628pYEIutMh4OsujrsUfB+n2ZUratvWoPrszuIw2bztd
kQVn0/R7q8guQtm+gQQrMYucoIZ6kMtkaC9A17TAL8REQe6U7pRYx88QW+KTH6ZG
vD53QMD/0BQdE1t9gwIVMO/5qt4em03vPbb8HEitggZAAh+/ZqNmvNnTc/gih0tz
jk+6Nnilo6IgQ3fAyS8Uyyha4PdgcufteEeea4a3NNc8CSQWjFdbHyf1Ic8lnaPA
Ep3sIjsLu2qtPlYzOkd2ye+D0n5dvzCJotkYmx7GyglE5kchQAU2ooXlGsWQ6lLM
bult2JUNJQyu8UQ2JrdBtXW7x25dHWz9wDvvQT5JATDpnwZQZxZgekkfbcn/z/gt
a8iec2p3gnIn5jlE8YydeKrJwtoJmOmLhYObbkLpNbEdQASTYhLByb9N8LeeLJhF
bz87hfVmIh4zGv+Pyv7PzZGsFi8U62p+/jQutC7TSxuw1CUFYbm/flCfxIOAdIf6
QnaUXBXVu7YvW1cj6mkgOV5xvH/b9qwhuLp04onKIRoPARJr6Mi+ZVsPFHDE3Fbb
U3zXWOz0uLP2UthPj7NbI3EZTXR+SgpoUDrATZzgRf234PixsTITXWC4XOdh90V1
8mBXIw8KmWeAmL9+lVhyVY1JgkCD3DvUCN/p4FZGcnhiOLHNbLjMjSpBuheJhzvc
GxAQi883FB0paw5uGBLKOFlZ/0TFbW1KVpyU+WHEkaWaGW0vPk0tGY5hARApijk5
bO4kZfhJAM9Xcwn3A2zkz6w84gR/nhUA9ESGJZcPu6PAuAzgAmb0Rntohzrp+S79
zUiqL1/EuN9vWULWXU6b7r+e7x33bwJbamwM0w145TwNnVzukjQWKiZYJdAqAzTF
c9yyNP9oC6A9LRKu+nj8HfCh+/ULs21+ZWxSjgV2ZIMKoVSuYCuzvCOvL/wJpYar
IB+LqsrXzFX13pQkz1H97PONQUsv8lQ94ACknEDcZn/bfmXtzjT5FZYNgWQqq1vp
3bsZUKHfxwGQ5nYwM3S1KMJ++t33Mu58o4uz0mF8Y6CgQ8vrtswLzAJb4LD2Gx3Y
g8o2ZidOQMganu9BNEjC2nGvJoa/cet/jE7K4iRJKndRq1lVObrzr/hNLsbfex7P
Y+fcYz6kwGWEssLzTP+ukI2kCeCsgb5jZscGJeWZijf0+Mf3xxsaWZvGLVGe2qgB
6aHNdvEPx1gUWSPchNyKP4j1DoE26E6y750hXJ2ElxQnx++gLqZr3BUHyexMWPZT
7vX2lJogs8f/19j+hlxhFuTu9VhNeCsDc31nC/whquvgW4WCy0tcvdTM3TQqAkbM
4ILiZyz2VBs0lantgR6/WiF3zMcSpAoVxI3mBcseboNWvLDo0J5hsLyCyh5hN9Js
ZMy82Hc2JKKOh0TZdKQZeRbkM8N0dqFJXfa1PprfWVb6jJGrjatZS/aoyBVYH0rE
HVIhIrGdPdcmr1Nh6YOuClrlb884ikIBJDbhV2hbW61cS0bNwAg9OD3Z3/DvDz+Z
V8A2aJiVoWXZ6ywsoluZVRb4lBUY/HvVpzHwZKnizQBGrEW1cwAoHDr8ND77+vkk
9xBtaFXWxbjCTh6OEDQfpBtwoJnYHd3qu+JM/tfhoP09ZK+4EQt3crAbPINPbgyT
KmLKelkVnLJeUXU7lht1yebAsOb4Re0nmuHKuYX7BY/M6sNQc0JsyLgkk131tv5Q
EI8U7cEtFeBnej/SAXrv+IjOuYi65cGaPAvfmMk0OCpLDvdqww58iGnr+uDGX9RW
hi4PrZ3F/Gw8dXavvBQS+TgHKa+Lfu9gqW20Cil+LiRioqnvoFS6dzJo/WCvpEWN
dRLEz3oCEKnqPhEU3GhFV7mPubnVaBA/DN6WUF5GcQfxOqLPgtVJbj6RrboCgWeE
tw6vSAKjSs6Y9vnZsLQnPjkoRCRurF+0W33fUwrsB7wtiC34GCnFTjfz70pDBE6F
Bs0BV1fJto2MlykugaHoFgjuPhKRJ/RQZkfoV9xJ7fSEZAfKcyM0DcfzFt50t90P
QvIy9YwycaA63SVyKEhY17zmf/tSRK0bs/PWo646h6csTROrSPoWugRMK3TNRdqW
iFS4htiZ9Aan2yTyupwnpnq/bZ/Myq5ygUMcvTmvCyvuuoOLOY5xu+JVg1M6Kjjg
aj78dkBXK1kXG4NC2DEiCt2JezxtzzbOKa8L5eEbOGZmHuaNGIFqVFZK5n1EXEQ4
H14CVcuCl4qSOuOSq8AOx1MXzqNFw52PWYxKymSr+uh0swbYMMy5O7NBu+Zdi0n5
911LMyLtt2MWjvPSHuZarZUBaPuditsxppdmkFaiZEf3BUsqlmglNU88IFgm1XHK
XL7hx9HfHb2x4AqXJWjz/xiKxehi/w382OCRG/lJXrsax2OL4YRcULazsOIGBDIV
Uxy3h0nrWZAarlWzXw1GIh55bQ2Iol0+wrz6IX2XEBRHGZmLA58hqY3jHXKk0rQn
VK2YQgCIqPG+zX27V/+AXknqnLSPVmTLvOhlO1FF5FOZGgICHeRn9ix4lQwewrhk
X+4noY0DRlTwNjDp1y7wqc5OWRqQRvTX6D+BbFrAKHUcfb7RjN7VpdB5LMQrJ1cg
M7Rjz/LjjZyf867I+OrCdXuBZMJXRxYB7im2Y4InQ9YEtPN6uVZiud7laUq3nagX
dxnyp1+7mnsmyzK5xgxJyNOb66C7NcZLst2Sya9KNPlRLzPRelUd3vKQIpla3529
63wOEBAGMb8c7ZTgtH/RUc5Rs0ye2T3cZ9arycflS703+/Pas2QInyVuig/zlFxU
buyfbI8orvLjm44YG60kpBiWd2EqjYBPlsdRHXh0hdTGKj9mB1KAX0XsiZOqKwil
6iZvOQwjbc0tE3Dp++dxQ3DQuEwj8SSYhLiPn6PZYEKwW98wWbjA0paVo0oSRwnK
FjVSEUAsqyE/OTCeErRNOd6o25GLMmRcmE0+5mnNhbI5oQxHzpx6Qo2hmZEPgoyA
wLeS1tJKGLYeG4s9EK+ZYsL2Uss+0Y7QipQP0olvNRGOxnUZo4S70Dng7mZQjnAl
c9lsEtkTaHBT/wGVrRBKD5lB2qaTxKQ8ivlnY/UL87OkPKNr50B8Ij+R+ndpF3OT
1/m9h7b5qqF3X4Z83BjlVM4T2qzyUX3h0WvoG7Vdgf4klCQ9iPiJ+mpYZmO73Bjx
LABKE4ywo9YR3apmuuX+UQoOrxP4umkAvuN5hfX9hxfIUEMx0sqQ31Ds1tibYe2j
c76b4h3efyyXXS1fepKy/5hOoyaC0ZNFVyKU5Wv9fmlStY31ZWGzUxTHZ0B/Ui3K
jvBDw8x8GlJUjrUBXIJYvnDEZMgfbmhcXFtRCNCVjVnQGKmll4tLQiVrCPBDKoYh
yAOJrlxgwczzV+c0O5U4TuKQ6FIwPaljAo2MFQgZQbVCDIA++VOQ91PisTs4e3kE
4ZKe9QkUqKB+0DuUFDL7VzNs/qFBHlGuh0kbPDTCCRG0ldFzmz8+JL7MC/C7rPG/
Zq0ixuH5F4S9vf6CECHwp0oejoBbYiV9GVpNiFWpvugSCKWphpcdbkYqE1vXRj5l
rzL0JWp12H41q23toTozUrtq/gmYNUTcFJ162Jww4Rm6XwZGRgw1ErnRlwovbqct
o9ZT5I5MsLkfEq7ed0F3YGiRj8jdGoKJm3DxtG2LLcvYTEHWJ2W7xRr15lWNycir
uR7oRKNZ9zxi0OgNzGql3LRiBXYYr4boyQjkM4CLfTPprSO56H3q0a1bKmuZUkG+
VAW5lDwOvJECWQl4CQyGB8Dpp4D0N9F+NUCizm/hu/L7TZtOt5odnSy8Jd5f42Ib
D05C0j1DwaZgQ87iwiuaYVLX70Rojoky3ZEgN6BgCTgAekJA/78VY6XerMQf7G7N
Yrec55RRglbjqLw7oVVoUoOnJWe0LhUMUmXAcaPQhLabyUgkrCvk36BMYTS6TSGf
r7gTnDW2jq6Eu89y0qXHswnT52VX49V+lMfTllwCc3v1DpTWfjZMd2v/n7BXKQCm
6h2GXO11WcCWRCgqmqRf8eMJulBTQ5nJXkG/Ynjqu5Oeny3VuEcbTFcLEy5qf/1Z
6U6enNCIgUCEwgrca+o4rN/2xprePn5SoMxLqfB4xANPSDtUbI9gzgdIacrquyh/
Dv//7HwiZyPA5sAnSYwNcZYpdm9jESrCxq9JjM3/+jFfwrKZiIPNMXJRRVBB6o5X
KAY596ZD5ItTOdT56Nl4UcxdQQI2TSE38RG9ITIhQdkJ+PpJbfw1C/NOALSnCw6s
k/EfAr3+lwaRXz/RE0OEeE6RiL00mPykitAFCRh2fuU9hCbOBfCqdoFY5EbMqJXK
NzQuGqHX0vcml8zDL3XQJZX1NB61XnzYp4rNiUqztvG22a6rSbCikDHu3dVqM86H
KRyMSlyAyyMdyOmT3OgqYc6nTDHOvihRdwo/42HI2Fcz5nyHZjP+7uObxg/wKgmm
S9CD7tAz7F93E2iimpq1XZAWNWC6QVoe8WCTc8XhN/rurhOaiIPBM8YEAY2E3UIS
qBUsp0LOwDAqIRTNuaw5SPhvCOvNwJOZfPBmrhOMwcX3RukixepsF6VBRoAsLZWr
AjcazI3Bxh+7ik5pZgQ4dB9qVue0D6CYgXn/2hYVxcImtF2vtB6YGU1zcvw/wXi8
gz9CdeM4SgER8j41+uDV3tr+X8Todub6lVFwXL//wcm5vPBN7YTpS0P2ywlyeQ7d
kMTnDwzH0f8Qt64FFxSbSoud9LZ3tkwR24TePaAQcrv6uxxUS2CIgVQ80bPt3N3N
RQ1EXo8fEAoh/V8CDbk0WZ8fmkzBWuvp1PHwV/76PYyYyUXm64ak6Cancp4Wug+o
2352AqoqQagxjUTJfAs8Dnz95XGxF/f3I1eqsF1phlmvKVPp1MiRZd/l92LPAxMJ
ihSPSznH9ypVHLgCbLtHBC/ndjeynR5rIAHacrFCq/XbPNPCVxmEDnArvB2bYTvy
vQpU6EhogTzhfW4r7xmQaoNeMl+IFvX2HqUrV53O8CbEyFFU1gzJz3E4925bM99k
DzHESKJ7QroGhhCo5+8JXY7/znqeeJlYiwXb4h1J96KxQIcNi173RwM+v5Oryk/W
2gWnXIceOgc3SsO0uACsJ3y9Er5x27ZWmnzI0EyKGgKjaV+dmySN2FYkHKr9oPAF
UDmf4iJHQ0/J5i/QA6Z/gB/la/LsaJga8DjBLgGWxbXdOLVT76EU6AF5UaixP1sw
XzX2/iXgq6dy6Y7KBX8FmtFoTtYI9ACXaeehpFZo/2s7RmwstR9rvuKzBI7PxfQk
voA5sBzXoLCHBaw7OBYESw8RJqyjWhSjLCxOnRF4JMxhU1p97HLKsOSxnspj5tne
1Ec4enVy/XGoFiQU3O616jXVzOH6yT/Y4C9sfupby3qYBB/xEQeMW8iTTks3VN41
NZP14SiDDW5G075gTmty/Q1Zpshc5dn0zGRY8ADBqyvXd351yU+3JcIOyX22xHqm
5su5xY+S7cEuw/xP3gm4JdqFzlO6XhVF3aN32eNRFcoTMaZLROqS3Ru8ImhWuhN6
BOyuDaIt/XFw4+yCkbUX919i7Z+TPd/epW+TIm4QLCgK2y0j88pRANybrNaeVAad
KMD0pK/26YnI2/EMkpM5XJYczehjrUQSazFNNDMK+2xV6qMkKmn7s5oJ6ygtB2yl
8GUxBpVtjsWOXrwf/okoalGExfmSCNoYJDGDheX0UiYx23fuft1jIzCopElokITB
IwsoPdOcADlt4rjjlEB2B2pLoeyrjSaqz9X45b3NzY+2NBRFn6l9KKg5StbgoHn3
CeczgTglJVkhO6yT8ocUn07ZQIPy5J1X2Qy9yKUfDrsBv7SA/eYKOFC1J6b7sxMv
nXz8MxV2nQfgCyHdU5kzz50bFBaXm06PKB63ezkLqJivmAvLWoRnvhtEr+na5pw6
H+hjQUR+tmTD3Di0MsTA1sWyGlZ4twj6XREHx3ews+PsZPXhST/hyiwc13Fn4CAv
EJ8C51k7z5Y8ski9XVuWUpSiE1k46aVyE8uvnUxhIbwnXoO4D75KHbpmCtUrPS3s
iTWWXfmqpgSOMySotG42astJ+8m4H2NiCyxa/USM5pHYloSOtUTlS2hxcJ+CTSq5
SOcWQRwuTexl/BcneDnEGkoJgRwTW2+ps/cnzhZC1WdjrI3BKcP3UL+/3E3h/8Ng
7XAxh25XVlVmlW08Eh86TeVEvPfx+J4bJwA3gDuDnoSI07HHbEnZaLCfkuZcl8DZ
sKrf5Hsk17mOmSPm8lgYp0Oblh8vo9K9F2YbEJQN+RIdmkOE88HkayKlSt5a5Qwx
xekUL40+W65jK39FBogHuYm8uuQ/eICPb7lJjLahrKU11rQGsOgi6if5x0HFFYbL
eKsl3sJjKays1zD2GigJ22nRrmZMjOvcnsteTnXA7SGkk8LCdPuPncnLYWf+6w/D
H92fiP3/J/Xof39jI9KmYdB7XxIVPwRoTNZbhSy0ZSVR3iwA7d9ArT5n2Em0fc/n
2xVbOcvNrVk2YZmxudEp6RCbdFrlB23h0xtHd2Krx+UiZMM4SyDwUVtgQdlz5KXJ
xlkbclstuWj25zeFMMgH7tTynBrMtkbDxql+xLJ4rjnslOj8mc4IBxfepFUNjlCE
Dn/26xcFqtW1IEdjiLhOvMj8sumAM6GBk+Mdzsz9J106pnqIlhhTE3i+Uh1CD7TP
UUcJbzayjqcBknZ9/a5N8OmkERPJ+k6mv1wmRLwDKgORo2I3obFUoGeUe87aTuLy
W3PcBXSa9Yrwsuzj67uswGJdMRTPPYYpa5pWGGEEUfpP4mdxj0kCivsaFU50Rymn
3N2hP88QHiZrXROIy6EoEEzNVhACS0PsGVl/tfaCkElb15z3ggQavIkkKYAcy9/V
11h3h/TMweKhd+zaVkP1cg05KAwYQCJHuCe/4GEwDJOPGQvyPG+kR418UR5/gQto
lj9KU79+XSvBFvKMG9rPeo+NVp2yMAIW2Q+Xcn8DnjMxgFqttbUfl6EiMupUFtjg
3/VUZdtIEi01tKcJpnswo7ElvQgkDoNstYAlKo2cP2mQ+VSHsgz5O0slOktTx4uP
xsfeiPGP/0DFA3I8xNxjDIHyud1idgtnDihiCArSREC5MbjWBs3klzgKjhgl1mB9
xTSAxTAlLIJkiydCBWGozdZpaJgxtZHYxhYKiV9beIjPQ0+Z8KU5bOqK8Ax+zeFQ
t8JC00BK+kIhExO94tS2B7OWPmLXexvb0OqNf/bAMsE4Os50FaHe+nLuwnDlTWeT
GQ2ahKsBP6rdc47hN0RR+C9UhLderebLK1Ersa7xdlUaskOuZS4Ci6Ymg0qQMSgT
CYqL/f55qvjabX+M8PC4oXb5SO/tP16KuGYcdANEEqt7HnLuT9Zxhfe0nGmCZeci
mgy2vhGZppBnwkDtWcgrQC0xrwy8XBCuQLTNDjz0dJk6SAj9kvKeW3GjUDPMC/Dn
IBwoCjZ7IdIrxRFz9QrJXPWSNAdGei5Tf3ofuwKjVmSGXva8v9VVn1R73lkNpZAP
0ldGwvw1AwWh16ij3be+i3dGcA0zQwWOUKLFx/4Tlu4fVV4HyDgrKmzdV36dJ6Xk
0mKj1QZqEoMxeakBvTLCEKuRKT9zsHSH5UbsGMnwiBujwKRPJmdiXj4+62tCdGgL
f1O5qUsIDzPi7u/6+68+9LjbMIGu+FQsoEJ4q2YtwUUR03HlOBtiiT1f2MLYk/Ew
81q8WItPvK3ESkgY9+PowbUmtVIoZ7VwARurkN2Ti0RFkrWk5AIWdaIk9kEeDHR4
Ok+1P+yb+j64Q9JZkJJFuzHxlZ0Y+sdhwQn6L6xDKPcv+Yi1BapI3+Z9BVjsAki2
X1+mVGT1Mmz0tk2HCK31BfkrFyTNAFpZ2NIzZ78n/rvx4JqS25q5DRbPJN6xdmVj
XYE+/szPYOayMVMOG54yKwjBN+fByKOpiEFKGkTE8HS7S9JwnnBavkrGMtkuarRv
87MZbPvyUzV43lxWOBNtMXcAXvpmbpkFAHC4TLwC2ah70EX0L8QrG27StaBu6krU
ImLYDFKaRQki+ihNzkdqToMVBCE9BF0M5MqyFjdL94IVWuewZ+s3NIYlvAcA3HGf
Au2riOd8W/Kth0wQRjpHspdxTKVYqC19xpqrxJuy0T2oAOMZU37nZxtFzDUD9qpF
DaXeR75fAqBSzJDY9rBDmLXbPeh+fr2wgszwzq0fc1I7fl69i6iQMxlKJCfwDqHS
etURInKtduOlrzz3NYpxTbWrMz9YCt2GoEFxSGCXWpb/mQj+uiS6wDO1+M11QmA+
KgVwIophBa6O0CLp8mACAu03IeAzIalT5ZuyYRRuSA7CEcCt0wEMkWu6/8BJOF04
SFvnm8SvD+ssnIJus0X9J0C+NLxXFNy9AoIJbHmsqBDLzOMcaVnAOXyWt3ik1B+N
Z7Vul5Nz3L4OoZ75zwUuheI2NX6F+wT/Hwnkef1n55VKdRXLdv6+Uhm8iy7BNPB5
xvsyVLTUwIX2n28NrpTcWgoocFO25sthcnlsjJvsOElo/VVC14r2IKx9o0pUV6Yn
DEyhwkXARfsa/au2x9HLIkOpqtH7sX+8j1N+kibi8UqPGVNhAdsBv7W1/4ZKDTGf
RJziCokIlkjxK14fWPgX/6JoLEKtKfCpe2vZ87d0ujTi8bC/2Wb98aSU49K6QJRS
lrAoFVI+HhUhKYyxriMilll/0hlKQihMzUc8oISjMCUExj1/UXEQT2jjDg8JsUKe
FG9971bCkqxWe7wd95YzXu7RQvgEShV6nphqXDP63o6CdoGW8ObKS7fO7/KfSqSZ
u4Lu5J9ut+aFjTgFUVF+odCVw3B+4pareGjxDRvE+KGud2p0rykCb3urxBoMr4jM
o1MGF+cEaLETOJALKK6Hnq1LJy0ZJk42i32YI1sdtCveub9vZJ9SuNCJtkNJs8JQ
qb3+1EwcO6MiCFEO95vguiIx2alpGSrcOTOnBSFuBCryx+U9Dv/gk3mJ4dxS0ZzN
OLCEqiarmAun9b87jM1jE3k0MMAIgWYgNZKkUmfoomkbIXShtOvpFYYTGGoaZZKO
0pwEpPn/ZTJhes1GB1O+sqgNmCiL81wt5ahD0aOvw8UGe2xP/nESc1wJbYgp8lWt
yUgS/zOE4mQFpReF1zXOolinXP/fUNHPWYZ3rEiVPKgr6Ytdu3FxIDmRnbJQCzBt
ftvDHjNrqR5f0YTQiqNGTeL0lezitAo3OkexNhvRHsXGcLRiP4ZYHuNnmR0iEyKd
bgV14sCVjWg57spQ++fplWvFU3AEe34/Sv0QbraZsyNaZJ29uk1hR1EK+br1s335
y6XFjBt73VrjXBXrCe/oQifPy/GosuVE3YdBa8sZ/ztepUnW5/gn2qMhWsLwaoCV
qZcfUsIND8phFbd6ssSkvpFpnEPLSPSZQ5B2538Ic5ZMtuqZZFtq0uO69PTczjrY
Lh2cUc/9E4HdtPM491I0KxGYLdV0BNlSdCuvKBa2YOH0i14xFbzT4/AGL+pIwMu6
8HQgbku50ZKarajBWBaaZt8r7NCxcXzcpBpqgeiaNZ6E3ho7U1N9dssGWjKgFkkl
BP+IFrcQZoImCUF6syhqkMucjZUyZAkq0hoWTVCtIvofehjEyj+GeNLqyS7mLLUl
mpKoe7wMgkwFFvhxMbWt72Z3mmefGGC1J4c9lL7GCpQ7kgpXcqaE5RAFWu1ImuoD
C0Z9Szs70dtvVUMSCLoQcQdKEHGWxiWPwQbTpg97J7Q/brem978mAReV43HrIyul
N4yHMm+vOu6tTc9SMexRCzeOjiSRGnaXdV3lt/j78B4MVBlw4dr/TUBIUCfYpkqD
4E6N7XG+ti2aWRcA1gWr5qaao5nUtHpFGGuwOyCz7DNS9pLDpBwJPBVJdLGa94yA
l6YMeQt6x0CkJUAvgNXCacUd4NyMrNHqm67rvoca8xeOSmz+EKre0R0cBEd0eh1d
BZKRRuNPV/T8Vowt5B1N3b22iA8z5OnN4I3uiF+FP/1Wz051NLLyuPgHfD5vdK1J
wFy1wzL73kTY9a+XJdniQK0tq1wsE3/4Py13CYEept6G+hBzxFw2vOijhqHGOJNg
loh0Q9X5s0P5nsKNhO2/p4TPEK4C9JCW2/00zthOGaUlyu8xRv8yX4mu2hIF1AHC
/n1TTImOKu6qXvXOqjEC6puYGFzkYDyYeAzqGcAkxrmlcLe4gAVJ7tATFZi0icSt
N1hhEkDlp5D1t3CerTskq0tivfrufjL854YrXMbhYYxVn/BNiB9gIaZQ7Urcjs1K
XK5c4YSlcELOy5MozHGYSwBw6xMOqkunl5KvDllcRfsXemhqVJUWphlVzAujZ7FL
epA8UJ4t5fOyIWj+bJDkmTeg5AVX6rl2Yq4wxqv/taiKtHKiCwxXqV3TGvLiNsm/
AQu4/M5tygm25XmMKdf/+HqLMcT/735sqevsfRC9fpSGqNeU+xa3+JiX2i1Jh6ox
hFqV4GM2rRmk+oKnHeqy2Acs8UQfETOR7GP4SItV7+HyLNW79BjvbS9rXw22jxgU
sypxNxH5gNRi5+9IUVA3cKmd865jt6y9Vj8L/lCv9H824e38R/BoUIadiJwVQE0B
L+s0LCraiFClSacqzK4Qq2ciaXOJ0p0qRahx+i4k0soE1YxaNRa+XTZ6l6LB3YiA
Oxr9b+U2pZ4LIwxGIjw9lGpeXS1cS6qD6zRf5jGzfU/59O9w83TG2ph/ruTy6s7X
mVc9xajx8qAKBzTELT9iP44rHVZTXnPWgCUEYGNrI0LEK+rrxyaTf2ubx3uBzvIU
uYEzM+hDAQikdaOQSs8gJ2Vcwob+7sPSysYRG5qZemzQgfoSgkP2JqBMZp+5ejsF
GF20UUexbGqvQCarBHMVY0NbYMKVO5M/FSNd9nYQLpd/GhYkXgTiaD/NhD4Y1q0w
ilv+cYaDQCrsFaTC2rmKf3JbH9bfONMA9bCLBVBuUb3C/qKuzsyrurp6SSlAsbN8
Lu42pt/vzoXYvdQ3nSDNqJWwWfyAPgTVRCmlLeRxxE2hgk6321kUd15+30h+Ajbn
GnxVUEduGnNP5HD5SWXgLHrM9fO9jiDK0O52sTh1vv/U9M1R05N67eGIxtAQYQ40
zqdAfvZcZ7h7ZtZ6KHA1297EJuSlAiXhxy8bCH+4fy684W73hY8Ec4BUTzT4wc+8
hYFY+UZ9bKtob6WpwVjL6e4D+VnwnRgWyjuNQtIA+u5yHezPspyx/AepHJC5u5KW
sI+t5Z2m76+U1XzMdVxXgRmnKpJZXmbvoQkDshflIoNXS2jdKQWrhsnB3kjcLJVP
D8ajjJntiUTLAR3tQvzqihazHSJYg7LZqI8u/B/XiYuKFGpqOWaikWXBJl9qsh+5
zkUZOTKRLjwMUo6EZWTLq+UxLHoSATm+DIV+gMAV9wWl8rrsVD24bGMje+XisXb7
oes7SO+78G6ybqn7jlvZlpDqjCE8neV5wtWJARD2mQrLyvQOv5I34/yLZwAAcSj1
xFNZo433+WCckwHZaiTsFfjsvdBBAPWDGlF3UXGsYcobLtOOjhh+DmVph5ffF/oj
gYEyyEv73qknT8rirl49EdwVXrt/T9tG0TpaupXZ79Ks3mvUSoOLQE/upZthTpzz
3j+Ll8rJENOfZQrTx+R/TSavSagIHH9+VVou1Rasr6ABiH9yovZzavA0mwHIRdAX
69q8GcvFKnW73kwbo/BdMIjhR7TVGnWz+MwV1AdhU1MOTzVGWcM1zQQjITk2clca
RHDXP/+DnSDtVeMIY3+6pMP5vgDmaCGlyhEMa6e/eKJBrXyAak1X4Afi1AoELZml
GRoO2uVcVsKx468w+P2ch7ItrDyW4Ennm2TXyBj2cIkZHTWQ2N8UeWYyoXLWVkpS
t/dEne6/sSm8nEYn089oBzxMtiByZ9y//5Ce2rfqdLLTRMB99QiVIMG6ZCK3D9SU
hQAmT7JX/mAmq1xcVI1HPUYQy3pnpZswMkRtiAdZOO+HW+eS/kWqg04plzDg8L1X
iVWAyrudj5p4Uz+hrsjs+hPlrDhTdnA7zgcVNRgLUUYcoENrprMLyPx4ZpPFAveK
lgKQf2R+/t/gP7jspaRgO12M2gs7Bcv2+XtMabE+Qr/rHeuZ4/LC7YH/nXIR8ZGX
zqy5npK6NIuuEoOgPV9IQ6d9j9bVl0Ua0U/hM7FyIVi8CRaG6KdjJOjfFCEuG+FG
qVFBjxUH9kgaaXnB2Pvdt7HGBukYtgbkSGwUkHxjNecvNSU3C0idXZ04uihEdjSG
4gQOpgbaCOUyYy8ExLFZT7H7mqrHaYlegNUl7Ms/G0jWcgEnnxjPawbustOJrJY5
MnfYEjORBmIk6USvfeeD5v8hlZKxnxdGnvtwLmoDvu6I7b3AZfQhvPGCdeuKv2/h
eCnacGrh0nBzOoxEVCEckqFTXOktlk4IeDlo+XRuh95HrynZzopKkTIqkJu7hJRw
ggAmDKz+r5Q6c4FHivr2jk7hW5qpAUdkxYbLerEFs7blFQXKPuvtCCvwjiZpAd+g
RuWSwY/u/nM/VOrD6wUf8Nl48d5HvNAgkA7EzxADWqSwqOtYFBMrHSib8/gnhNqm
OinBbr+SgW/lVEpP0xzR60E4fJ739wRRI+4WHAaf9wi+7BSS6nVl18ExUUqB0yXQ
5vzFXJhWEu6OP8LN7tXzAKLRGxKYfFTx676ZCkL0/ImvAdBDkCCH4csKVngL9bpJ
At6W9aMLr+VyoUQy/1DdyrDeWcJzGGA1G6iTX3W8dCWrGFVBf/DjukXtX1lYR2qA
AyuAnIyxM39uZPaU8PvI61g5k6kYzj5yM9g4rW1bxtt+AHBjCufGNiVmAK4F56V8
WBiglYvcdmaqvw/kGKPdFIv7Nngho69COHRRd1bol1dWpR0+QB/s0uCRdXkFSh3v
ZlmAYVAhEcLWb0A7EteYIX1vsqW6NqE5DNw03FtXNNT9zRkcVfLh711YRo846hmG
BRX6PueoNECvnAh+bxxX9OJahVAwjMBj0DTymwmZAYTykij71beAvNBsVbFwmx1h
Er9Ub9k1y323f/yvB2aPWj3QqCZLNVZXte2SvUwG2pJ885rm9AFBt9oLGszAGroB
L5+TVFfl+6+YLsTxZDo4poYgGDnqMwXD27QQhvt4o2TOcx+EaJhmH9WQxf7+Iq8n
rUV/YTN/ys68yhPLD2GmkDwid5cxSUdbuckZT7OwvRpGr6A2DSrOvEpsuo6BxTxk
FPDI/Olkj2gPKn6pB5BI8Ft6zpoEYANkN3omuW6ijC8mJkwCQUK5oGUc0TvyYEoq
C4IJv9eGdelqfv2KXt3UC850DWSe/oyLwH2d6znEEXcLgmwqgYJ/m4rCbrSxS3+F
EStHKEedlG2bc3FQOgGhCdh83jE+YsH6XmRQj9ipIc1EE1+stsamXDAdfdPYXrLn
mFdDFOnTbSeDznguFemicRwa9PVN04ZDrbSKSwrPgjDHC1sIObb8dmhJsgJq014P
4cFrWz5WXsjr43C3KA8FlnUf2aNOTZCqvmxbj2qwFsBSVG4SEd0dqNquoNJYxIFR
BY+A5e/Iq7UFqAA1mXjsUBdg2gyLsPjvGZ2pgpSfFJYaUr27uXN4BzPbfuW6DbAJ
w32OP0Vpb6Z0UXjrbEdj4ZMr7nzVLxYrrEgwl7x3KqG2DMM3wJ2B+m/jDF/Ni6+q
Ld+hHuz3xtXCiBDhVddKuiPNZorSvzgsEDasuyOB5YumD2rpHE+y6U8BW0KJD3R1
o6UBVUuNHgdBafUdU7sqnSS48uN3FDJa0kvfM/Tg6JBjOf7FXTkQonUfP6MXzNwU
hHgHdaNZOZIKzduAgHjlKAtfWPzPjYQRdUtwLFQEZNSjKEpg8S+hfBFWoeO9GNr+
jW1xCGimDsgEWP2GqeYTJHxWJw3q5iaeLVGk8cskS84t0ViRzT7q0TmCmQRad5qs
imNjgTlJxJjYr767DdzgPt3suAuTQO99EdXrnuuuMwrlOREPQ5CZS/0fE6Z3Ohkn
AJW3g9x35y+xLQeBCOfxagjU3HBFCTOTSGZV6Ezn89qsAN+/N1bGB7Dp1KZ8GOsJ
KiXpNvNQEhLt2K5QmONTYiKUspWpV33Obq7n0iH4HdhqutBFNDUdWOGMdIeubLD0
vObMtCPzusRQ4uXMOKTnPBdCS4PDJobj4Ex71vojw7Dgn8n67X7wl0+iX5hlLOBh
QoQGHfqOFAwoBGTfExCUJYFKMzjTjLob4fNc+scoBdmLhaMaNc2Th43Fl3MTdajk
AKR78NS+dUkdGNh74s7YDXj51E0FDlr9IkP4Sne3/cdQSMe84Wdq6MnSpVUdiS5w
f+6VCxcDOHidH5zzZTW7cGHW6rxhrjWXsv5p1nB7EL2C43/VBl3PKhOtS4nHRy/J
XzbPBOXHGMAohkH+kbRbIIJbbbw6uFlWDQg+jjoSd04kzRqLXtL3cHFA2Im6t/eF
BEV4MhpptXurAiQwXwRgt8MjIoA55Wts5mmh5TXD67o/C6F9ub8B2X9DhfG8oGeY
qvQGNOOCDYYqagm3wkuRxWvTF3x3dryNskNObRQYy14+lMOJejd/UPpnEOPfXtCr
GSeyHLbef6rtuhxt7dlLOeUVOLc/8z+WM1+lJX9fr9GmOroiyI81b29k2xLeFyLn
r6iBFyrnso9W/wM3SjDscLGUMxZu7x6J3e+qqb9xzvDYeqSTutDYZYLj4+aFu3vM
qVwlo8VMthhoYXID33HQwntwi8q1N2LP563Yjf+vny8NfskqoF59yE/0HDdlVNRI
655kU1AZ/sHFdXMMFcs+GjPBcGdOyvBg7pF2PtgIrjiB7kykVEk2ypc12mxjDVCn
9k1ksIER3HIsugAtmp6pUd3tfwu85HmsDq3k+3iPaywMpgS1uEKrC+j34cKZhe1z
kjdS7oaOrd7klp7tEwW6ag==
`pragma protect end_protected
