// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PUqYSVFkszVowrfzlWnlRsg5D3r3s3UgEkC0EXGOt2t/xbnEn4q2y2LDa3arBPWM
+XbBTeZBL11djnuHy9XEzXw5yF/6jY4VPeMfFOJd90rVIrOsHGXZgBBptTCAnQw7
g5bO+uirEfn4L4fHhCJxTmzD1XZwcIvLzCVUDbPTVIQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
029T7E3mG1nfbTE7M8UCJ1T5M7OJGCknEj21KSqd1NU/T2hC71sbmspWfM//o/Tv
bxVsozMc2eQqU1hQ3vfwSe65QbrolKk0gnBcXMhy2uB+IBQMQICm7GrRgvuZavBh
v1plb4jJwLe8q2DfjEWIhlWFAdbTWBN2szh5tXZoq6LrjVtplYFKBhcYJSD6ePcI
f+XA3Ba5sWInLs58FrMfCjNDtLkhXi7RWpPlPMzP8eBBW3MMVyjUPOq5tpHjcQMv
YOnBSnAETriJ+p7EaN3Ln6vBvGROmQ3F3yGFLmr8+DZCcPiGivB+Wwj+uXSH86TV
kYSOnOCbVsnTWKRUKaBLuqcmSXiZXgLvGrQvUyJ/qsumGdjpTIRlzpVENBZTZYbz
JUua3XFF7zu3xKpBO7RBdaj9fZEQfpyDuQaf1/YVg5TAivXxfbXypThE4cKYId4r
D+bPkvAh4YnWUASKiuvJgoZ6fDnz2RqEeaFQtKTmEWV2unxELNe6cq5eTR7XX/mD
IYqUiQiWINGSsqFucOpxerxJ/pXqy9Jczm99Eu5VHRAbokkgLfnUWCIoC/okh+Sm
Le2BrulKHlh7QlrLvZauByTOpReL91I1dr3mXF90qZcsxDKNDDgnKpEGrNoEfBaa
DS0xyo+n0fRksjicnv7tIIVvdw27g4ueTsbSwPgNAFc1sMRwVGMVYqCPPPv0WB80
xRgf/iQHN3W+KyO0yCxzXZ22hF4VtApCNarxrvYDI9tRQfukYUrl/VTdJgik89FV
yM3S2W5ubPUK3QpyZhwg6C5YZQoC2g0wkC60rVeoFOAVRcefX1p3QcQAMO2IuTsk
XCQEiNeha/tYew90e1hfCaZXXGIO/ZcJCu+HiGva8V2oGVbJIWr0A9A1ThRBbVGP
GOEe5Rv3pykWAp+mXSmX4VCw6yB4lDu5tCXVDsPhQ5Yv+xq4/Fq3UNN1iQmZFnT6
7h7HAORP//tHnTL2cFLbpkcAMz/QQpVAjprU/INx40FpzuLXw55jwxg77kOlXQ0k
87usfd0pJmbOGtJZtCXiBS0quxS1LB9IeUHRJ8xfKGucie0gEZY901Glf+gmUpEe
3kOCwPJeo6qilfdgHo0K0J8FJZUwcScD1zk/3Cclzi11YJ8tePiVDMVP6e9gPP1d
K6gDV/uzi6cOuv/FNa7XrqeOE+x8VMwtD0bmEOjd6ppriDqZi7q5l/cHQEqSFTgE
JLZPSDoWkUH7Q3Od9t6DZjRQxSrZsgcxcH0zSguREKjIH86kPXQvgK0+45a5Iyds
bXuD4kKuN2KnVeq7P387Wm/S4+L7XqzxXhTCLb2/TW/ExNz9yWM5EKyzgFl7t/zd
HHPgO9GToSnfZC/BU832YlalLHtsdT32xnNugWEJvvr+7+gOp8SL7mPI03wFys1X
pJ4NkXcfMD382PuAKS7XJztegUe+OaLadjRAc2WjqgHLL0/axpFbW5tQA8SZXMBz
y+kbzw+wHY1076l3txxYG/ocHV4qafW/H9o95Gxu0bZqK6IvvLCU347cLpAxkfrB
cwYLCkYtSXuCkV7GxPbX2AmPU1dkmI+P0dHcPi+6GgnvUz3CG9GEOr/POFKQppDS
DHJBjdG95Q4/peaKSU9yR2X72UOTawxHOWg4wdwt5oZ38MTsp3/N6zQNSHadagX1
W6GXKZEyFPrcIZ2H21dfIpS4H92pwrjjRJCNkeSB6pNcV2xEyssMzVmdgM3r7+bN
RJvjk1XZV67tPqlAc3/PdsZRJ9xZPJEfVSherG5FMHq/ssxLbP/5BN6JtfOs4ZNO
yao9b9kMiApLsIZH6839UVADd+3BD0xErSjD5EewQjhgpP67IOJdvlUaGZu3gf0K
pK9k+U7Xoe4djL6rAWkW/gEkzd/g6YXtHUZugdmJtfLY5Qpr47kdJ73Gvf+lpZzp
Zil0RJW0O5hC91NxKaHYy9gOe0Z4NBq8/3ty3df0nYzVEyDVxRvgaQgAVh5nvfA0
cl+lZqfSXLSLCmRrq55FD2ksZq1XGs+2ibmalJAhQKrPMv2IC+z6wprb9g+vcZnG
iC1QxhU1OdTul1QIdwDo7msOOam7PwqIMVwbWWeNebviDLf8tjPom6jLS8LaSIeW
OW1EVhsowzxfzzWsVOuWy1sEe1pkIvqDlGkFag75DfMXhTftzUP8LYCfcu4EytGQ
yLbt7vOiM9OjnKxfkvMrcHF5NANN/pwRoryfMpP3X54fatk0PL7Tot4KLI4FclHl
rrdp1Ko0phJbNkA3XDNzUKbrk02CnFRjgY4G2JmPN3yJFYQY7854BCNDvyRARAHh
Olv4SCPu4/UgYbIqHQ0wfBnCwCqC7dzBBb77xHhaI/99zTKdC1JCO+sp0qNDnXBs
mrSgelrEu8LNtu4nw52Ita2HkQMKOejcGE9s/uj+fzpx3KZlvgxbwAVezJGPmwGh
USA+qbP2D0vL1YGI9E1X+5HRElYF6a3CdWfR3+iA5mfcH8ikCj3Q+RXDyPhCKrqa
Ty/bdH5hlVrBav5uGvgesDw8frRc/rKMgtDXi1Nkfst4QG9RTGQr1VCv2S9psNEV
jsvFESJTfWN5LengNWmwqG8+eKbTHpltG3HiGcNLY5Xq0x0kchUQfOKrdURdun75
0vY9zVFntwQAjU4ok9BmlKkC9i13owJYmCFAhpXN7VoXMNvs8ZxkzqDbIRzV1dKM
VOnWL9vjiS3gJ19x6ES5GEg4AxvZTed869pRRlxw608uoIA18GfIFRgA1tLjYAP2
aoaijZxfTJOSyCS/wiyM33hELPnW2LWN3SQBzwMAOrWpPT8StmiTuZ1811zzPyN6
DYI8xQd/UsTde8Lq2Ir5ckc1kjuxVB0AXV9iK+lG2PFCr/cBikLn2K6/PpT03okm
WbvODvtl05JTu7pB1FscB6LDemC/6jossNUzMZrYNGvi8Xi/LXrKTmN5UEXRpMGt
DzcbmNa+Mtg6DDI94VB37+BfQwevrgLHOByB0nDlIe33j+pAQxK4IiAKldZxB2IG
meUkzaZG4vt+kL2kwctYj5HDo9n/oWqcGdvdMaDY8og7KCE/EDuyFP5MvYrvVwsI
2bNA4JZ3pvQ9N86cZwEjv04YYUWcGdMso2t8Fby7fRWJ2AouJGfLJpStZtXRZTwb
6Tb+I6SPxE3FU33vsLJqFaV2n+eQ/wHNDS7OZBOEAccCfOQcHRbBfnVL/InVf3IU
10pNjhyriWPTeldIynEcuaLXP81qDDpls4SsO5RoXKF1Y20ELP7JunujPgDuDVbd
UlD2N89NmHEnAMHE/+hJXAZbiBO//8mxmrRjsBw+GXBaGLIjH2sMC6fIXHXSlzYl
3WloUCvAxT0ZOcvY0fc6GlGzhNC7cI3fadyDipmznRndmMsJLm1I4DeowCWUXb80
aVsPuHtS0r+Vi6oJi4QmA7i5fP2DywNf5CQqdmiNHayJg5c2z97MGNMX/E+m/fFu
h7UDnbatJEA8BGY8/gpbgxKGBhrRF4Metw2qdbDZeTrejH0jOaA8iYX20O8pgiDd
3cO83HYvdyp1TayybHKK3k98xhuB8vMXkHiwJPcJtOIs3ctKBM6vNUrj6fGtQ7Pw
PJQuuD64yBRD9Y1Yq8QuQj7kpZ5f4LIXduB+e94tWqRjSYRYKU7SoZwwPXmvR4If
eZncETr3z7emMdwq5fWuAN4YJGEwY3lb9Vqt1dw6d5Hdxk3BghonY7BV/ltOGcpk
yIeReZ/y6NX1vbQsIU9uqg4GpHixEc1/q8jlQD3qgNxlFmTrWeO4i4tTrhoZ6nNh
fJhBTHDeq2O+u8G7lYa/rBgvOIkxt/1vVK0PsMvxbaMEvle1+bWj3Ov7SqpvKBtE
AWf+EdmysoK7MbAED6mJmncwHJPvGeW/RADUjH8L2lGyeeWcQXt/Cp5+baIWKFqC
z8sx7lXWqMtVCgew/thJEuURMCxRKEeEhgEz0lklRw9mfwnlbNZGt9V76bgqw9xF
tXsZcY2SOD90IAwjk274Pf7EHOgTxZpOl/V69Fmrrcavz7H5dDOJbLUT4rsVXoNC
9fo7tB0GDngjdUVyEjE/zzWOknvwOEy/BAO1MKbG0d5/94rTuzDoKysP7/4lsSKA
57ERBZcpZuKnWxgiWN2Tx1IIEQC9O6HL98NmquSgC6Mvf+ZccRbTlUOs8dNYRNnC
35rqrp9yhgyYTVc1GV/72IzJNo12cpUVdV4krUac3kH1GDP6rIqQA9OnVUvpSZya
uTXcGjQJ6l2FthyItZz3xwGaD5lDDienJr6FQ3d7rjflJ/8v9gG6C+edWBqlD5fV
CNiCiPvY9Xt4lfdFKrtpzbAtBKmej+k22GbtTzkS5p+RBiKl1lVf+jaJVX21/o1u
YsaxmPQxNLn5k/wajv1MdFD3eCBdKbFaQvgHqssFDB2ibTQEpC8nQcw+98qMcR3U
UT8AB8jr7f+glCquR/3/ivJe/61cdSL9RJiixnzhkXOrtJIn5IJRJrpULQ4jPhQ2
cRQ6B8z/YmcfrKpQJcxMKFQRGId+VKuzj6KNXGfbVjkgHM/69CFyN2HhhUa/YA0k
tqEQ+noeHzdkjatsDQIGf0A4Gh6zaHaAEhKWr6y5oC03Jx6BpOxbQLJpGugNWCst
Nx1oy0SamEyaWCOz3b7T89ZPbVEV1zSl6gP2CoPSaVPQOFaTKJgh45RZ0HAgtkBM
3589HMglaBPZEg0+rQP7sUBJDYSlpXAV5F5YWaYOfXzDz+tajW0PWQ2cNNk1B8R7
hxiJQyA30Hq+iOUobJKKuP1gtiLtgpLEkTGCDiw6idcRyug2Kju3ig16e4mhkKlI
HcMOEh5ouopBySbMkicmF/V5mNMNqxr+LZJDJAu3PNbJ7eBeONkQVPvHnMux7cZt
y1aL8HqDbpdl8FVT74aVLbK3hHX2TgOamG2hEGN4UOzCkdNSs6bQBanFqYTyF+7Z
8VMqOoBiDczn1OVDHZlNBkyovPgt7N+7HKhr8hsAChUuT9j+P2LpGqnCPR2Dgb7n
uwwFLbJbVrCdA6SccRG0vevaPRSEeiQiGZWBASWOxgDASiaj2Hc4BDBNIEei7rn0
xs/pya6Z3+4HsLfHnj0W0VxGujGrF+7X575u13+F6co9YBMtUM9AVDjaOYMThdmP
PPie6pcYvlSR72slEQKGvcUduF74CI2CQMIIuQtIpsQ11pagh2U8cO4I//xsWqNj
zM30PFVbgCdtoH7QSQooqmy1a6rnBDuCSnSVy9dWzBaJtSdBvvKQvozmoUzjI+HU
21SpGdvDVCGGy5WZyRVNiS+uxSYRWqO0XXKGetI0IQYyp7z50wjXS79x+wKEq1nR
ECZsefxWY2yhLlqXMh7s0U7bN+5d+lwhlUE8KDathF1uU2iYGEy1SQUotVYwaOJx
TOgXDiPub2HP4O38xRFwBmMMCFHYDQY3Ouw3TSjcxyM3vyVZysxvGuJwjH4tMcyG
9MZ/1PEceQasjBdDH5q9u9FPkSX0ESvoUX0eyvDzvKzHsxYMne/tIjaQnJrAA1d2
/zc1nvM0ecbUDvEq5XgHajACQZZhSqkW33XjGnUmuX/Zp3VXXwguRbhUvpjKEvqG
/5/93hlAa6Vpy2Pff8VmKdkCQpw+uUr8pCqPEysjXGksrBolnNlCzuYWInCgVbzh
cuTiyopw4JG6cc8X1YrmDqE6RbMzW/sP/+wFumyOpB+d9mcI3sd2TDh22XRh9a8K
LvJ04L5gP1BchP7CfMpdN9v4L3Mn2aOi17K0jzuZk/QGCCk8f1m2/aO71GzixZbq
qqvkfz9ZF8kmHZRGyDoogyfvhNIfwRH/2UtKBN5eYqw9BAgQ/paE6MF/f3hGV+Up
GvKZTUfTY+Pr2h7F1RLMdqeU+0KDFVmykmjILCDp8TD31Iyd/AAMacJV9eIX/fVK
a5yWwA7ZKEiFNY91YPNQCxPEqVqFWip61fLToAz6338X0YRA3AqDDZ0FADLm7BGN
38tDdumoYDobne8DBwOaUd6UVlDT2pah+H0jELE9VzeJNNaQ6wgGGjcF4/Sku6+i
IMmuLbDB1EP2ed+NN/UJ3F6GCD8X3vS1z9ETD8e99HOSHgtnaKlrDjU2aub4IOV4
M6NNypbVuUH73awa+BJvKe7PkA1KrG/mXKnOr46D1bhSDcqOTYJMquFowHFGny0g
hlLYYC8RH3n/BVJ+MDv8UjilT/Q9Uq/PY4go9EKGXaIJCeLHSKW3G9mIjh18J0s7
ZGMmeZnZBM4OkCjzKA7wQglhSFFgw+BRrTAb1+1IjnzS87G+p6bQGYHDSIFIznlX
a6WI6V0YNhKwzwxplROOKxPElEMPm5DlhyKcDlI23axrK2z+ok7TX2sZY6jGWcI+
62aTKPHPvBeH7+UnI/G5ovxridVi0GDpOc/rIhZ1E6BUhApooxNgpaHUnZNsYOB3
T+xCumXaHmPlh01vm8Xm5sIz7P8O6/iXYqURcx6TQKfKruu5wyg9DVhWwMzC0C12
/fbyeqnjVuolWBGOWB/PLVZYqiHvJw3MSP4/sDwYa96nxN1ImEkXa8PyGsUaJfCz
bsG33ua2t2cBZq1BJb1t/YhHZKzSUa7vIhexhNfuMb5FxYM2dFsaLUPDIT8gy37a
Owr7pTxZqqrBpdDl1lffRdUUTQNhecjmssno1XoQqlqwqXgwU4fEG7tETcao5D+n
/ROLsVVPKRE2WTQ4V7tJhS5Z80iDAFPD6+fL8qUSBi+CCu86hN6C4sZ6Qhz+K263
NVMcIWkXOMRJj1en+l43yweKb+YLjrRmWDw4qy+i11gQixs1mxPfDrQrl2viFx/H
ZzPWZ06ndwu0ZsvUis0ochV70FGu/kO7aqyHaWRGLWOTSWcyyY+jC/HWuNPv6KAS
xshaHSoD6O+s6zRprVrKJyZhT84hLtJqDcDQXMlHUWFhail93++pADixIi0K9CQl
qrLgHPOiMYw6J6dCo3RP5Og7N9j+uQTCaiBh46RRemWxRofKflC0O2f+Mzd5nrI7
HbLWiO+l/nDLy1gpg/iqQ5miT0ze++36ybY5qO+UQqBGmX1TNeDJbrR8UjDKEFw5
cXlMgw+GCf1DvXbgSiZv7wtc6P8MA+3WgK5HfKvzEflvLCX4JDd3MCGFS/Q2ZwBF
MImFJKcCd6oxD2BhwAl7xzyYOKETpU9CjVzG9PbQfMUO+Ir6v3AkHUz/FupHEuVI
Y3RQ/Ie2WDE+N8QHtsKqlPNnKmbyof/K0j7Tb9uoQojMB0vExNiirwq2K0XQDvO1
Uy1mlAdOGbdyj4zpxyHoxzRm8JuQKMyjPHH1zuY2d0D4u2/QOGIkI8tl1gezUVZ3
NfRJq5b+QM4INjPiw286lFyOP8BDqTb2fFtBTzkvIGZthGV2jDbb3/EJEqKiS6Ec
bi5+5e/gnQ6WcUQ1Id/Fr3s7HKRPw2AP8E3e5UWxeb+5wJd3ykoVnSelyKkGgAmI
BWGxLiWGNUXldOUT1KSnXVEZ6Ed7daXc4gVgF8Il+WJF5F3Rn5uKiOqnuw8u7T8J
6IXEYnsWPhYl2dIx/n7r8V7cXHNcGGTjBbGM7oRSVwdr5UfaFlTNcV5prEoU+d0J
I2LMlMcnyDBtEY+IvGaMG4lMFxIydh+aQT7+WopN9pigRgrMhzbfLN1BEuqfSrTV
4plYJ75VqdW5qwphBjI4c4OoZPNvm7gelSd6tfKhA619rw3lkCvQVA8ZWgAlc19R
KMZrmZv9gr245D80Z+0WNyX1gAplWERE1DTRgx9RlooOuP7WguI7wXNOIAHG3XdT
iUvh7GM/dD6beJFEWTrUvbuIfMM+U1eLRQQscMy6BFfc41tyA7jkst+ZbUQO+qzc
JZbhXDUF7eiBVA8sry/PtpEnRmkh9J9q06tr6UilED9ASRCRN9gDOEYdoJGDbWJx
s7mgsfZ13Du27SKH8aEaXbksCEWhmRvxXFSZJZLydIwZYgSdWSc666Xf+iBuas9e
W3ZVNjRhoXRvH/gYX3LS0FOZywnxUiRUZ7+z0oJAViVTl8jOP07YkJ55nAGmWteU
ZwYFoDqIZhUrxsBuDhNjUIsjgRjiFTRJh6ZSYs4f8NKv31Kyh1XV92d3n7ybBxqx
qhzJtyVhgv8LIRP8UqjbCt6hz9m3/GbkYf0R5K7DWoDKnQzZDLz4NdwRmh6JvGNB
ThYGyPpfvcpBVNR1ETQAHYJULgJrUxBPfkYdwMLDekSHl3MtFnSxH6e/4s3zSJXk
aYAtekBobdSQlXB+HjX9cd1AKbVZIjEB9A6e093c64hQZj2gUJUE89HB36sTt99c
b/0BPZRTZsPeRIF4fZumeDkdWBCfNSuoCVXIOubzw44vUBiNTjUgnVuePW7cfi/v
AbiJ3M9rsjq17CLxYIspnmYQ4T/tNd3vU7YQAUXRJhhIY/cZcsTrqJgySXFBE2z0
tkjY87Mhwq9k16tHpr+UgDDk7/d1ffGot1j/YICtwNBFZNipDF6uXBvfx0uguiSc
OJ6aYlv9rgWJ2HY2vyqV474puSezg/t0g5K3UltSv1lRnHz/1Ayn9POpcEeZZ0PM
uoAelRT+oPZH3FvMbLx9KezkcT+fQ9mDr64Jq5stEBCsbtMWRx51I8L7AGe8JQg6
L3U+VhO7lcAiz7Bqzp288pgrzwE7R+J50qqLVjc6N/+f3mh6wjEVMRWi1LXjNj2s
J1xp5lTP5Zt5HGpGR9RKDomBXUSHlkxcjbpVQne9MQ2xZiLyjKGumzf8p8Fr8sei
qUnhcoW0MgrcVD8icYjuKoyAEchlAL+bScVOzFi1V/liHMRLLnCZQUdeQOnnihAQ
5yWn+KacwRrm8W36HFS+9GIxSeTmh0TD7WoTjcm0hgVq6WI0tZDeL5l7h96jMUPG
AuzTX4sZDwx2NTkcuvVbR+zEkHep1xgfqmb2Vfo4jU2ExS6KVeq7zpnq4WCDbHad
DzN2RRoCUjqVSfIn6LsLUzl1fa1HMahZyzd+t1QfxVNQ+inDTHyImzofFj05y6Ce
GsxJXN3etLoQYnqKI5s/FDEsvjJvo9Es0hWBLad3IOOX95NLFCCkZVWM2ufXn907
AIsCyV3kmDrB3Nha6KUdvWPmz9AXID5AMPt5nG9uOp2gtO9Sj/uB3Ws9bZlZ1Tyn
i3nfbg2lPraqAIJ6td47hRKdmkO18/EJHq2rtcHJvnmQbmWAwgL6CjCvNC33Aqi7
+x4StBmGvJX85DGfO+NHObp7zYI4PNBTsCtsLFdgCFm5yh06dqRIObXofdHKeWxx
GVPJ01C1fUFVH+p+96Sx5eP0QdryI7a8i2wZuJfn4SjmbwqFiveVPUU3HtefdkPH
Mu+fnY/Yutpbjd2g7DRmUiWzdZC4LA+lN/KRsTUiN/s/T9PNyCcjGDoXkdq2znPJ
pzwc5OCVMm8sGne6F2N1iJaWZj/Zns+ui3z40WcNuit5qeZhVCoZI7BI9kUfCbgk
aBcOIhHjW0m6006yjr5IaKJH1gEyCPgabBeYVA56NJtbmNYGEUh3eBtlrHaj7GX8
ngwlV+wCfUqFSxO/F1v/c3rEskuoXqLVS9twHddbZbLnv79enQla7CuFIz4xHWIp
mYxbFxU97pZ1jRQXv3iFIhpBFDfb+3XSXemXz8gNBxC29+JMfxlWdx0TNh+Yozlq
1oP8d56oRXa7PDgh/8Mg15aZUifHcVF23uSj+q7oKOoqU7Efc+pvau9YcVLc/coM
b4zvs+YcAf3jzwcxNJHd2ojZI4j0EJRv/43zChfh23nuglanIKP+fvs8Lvui1U8s
e5qjFGXFhFHyHhXDgmTmqK3LV1+8ALIosxyNJit3dRZldd7SVd7hjJ3Amx9OWnD1
6rKBfTBQVXYH4Y+oaNNiBU7AaiF70PvGjCinoGcpQiibobTbv2tD8uSYPWhb9/D4
wtUXQEut+jiVIio0yUd3GjlCqLoZEvQsW90u9I9/YSBw0+VCd1X796gaFx7PmMyu
hFBoGSEiTItf8dZioqZrgbksV73MGPNl5G9jnlrnFUMJLEgZfkFfiiBJcHTE9Dct
lHG4JiRI7YHl9jXtjdbFdXWRutGB68HRVKA+1l2DbBsY+bvcQroscFtxhd9OSmu2
Df1WqX4BCnkKhmDkS56uBjzppnQFRWynreXxoBmxNwO+3QnlOrq4ammxlW2QjZn7
/0BB6k2b/+HT34z8fjCDBPmEKvgjQr+Uv1y9X49kLN1orvNFdArSiM7bB4pSfAlt
e9Pao9YPwqNBXK/1YOOm6Lv+m3/z6a/kcJyh1hvLgP3hX1ynGcINU0tUESeFzQub
Yvd1wNwe6ovi+ahL/ORazzjO2IVhvjxVt32CHQRyoXhb8Ey42gss8YBt0oTqoNaO
ulatm7IcnFYDToCMzvJOb3LIuVO3+20E/y+MgwBqHphD1QhhntipqHGEF9+ebIZL
quEeK0wwsV+CuBZGdp1ofPA46o/1PxEZM6qQonbX22rJU02mCPXAMyqun0ZrfJdc
fLiSJo84w7usqlJ2jwTXzwOKbpy9pSfhMGP1AUPOHuO2k6CQVFXxgQXkeFHR/IG7
cokjia7UXGRmSsZmbDGOKwIkDpXfbYXgexofNZBrboyvcPIDdURmm6rnm+duOnmO
qiX/bnbjrYf3Xh8aUw6VkWq5n6p65BsFj7fh2zwlbLQQ25i89fEdHUJEdC4ehlkO
RQ3sVwOtC+QKDmY7+niLxas2NXMP9suCB2LKgGBDECOasYsuv+C39XRNrfxEmwzj
wANBjuDaCQVh75qGh1ep5aoEv+JhbNkzXsi0PcDrb0zbvD8PsonEJHbcfXrPS6f0
EvSnAzORTx0tHpq90OBHfCbX4jK3ZGNpDu88aEDaPD4EXLEvhmfvRJRDzSYIKUPP
RCk1TGRD/4pFSy6ia+pk1AO/embRrXmIRnLxnv3hEUQScTpeHxXuJwdIRKFwrhI0
kMavnhUL9tUFEJ62FgBWpoc7HaMjKWXEBdqbE01q+a3bPTxwJe7o3UepNisOss8/
CSIanpXSp6ObDzfSvuFxZrr/f6BwQ/hEohK9IHjooYF960VOMIBky0XfvzUGGnOw
YtDCzPwmI73aNE8SXm1V/ZrgwW/OI7qvI4bvYwELOBNZM4LSOsE6wHYKef/zszNu
EurfZhwtNHrLUDZWF+RCFFB9Mnz2ODA4zvAuo+l/IjlTcITl/B8h/AjFY7erzQ7f
efYGR5aXtjJicJiexmYwBVFZ0JRusGwR4iDvVyPBf9EWard0Dja+OE/okH+sTQFX
uIowhxhsVcsw40Dilom0xOG3FsXrkUI3s6ycYN7rfJ1nQFZnjUGsajFLk3kdboil
yLHvhdzizfyFwmZHECPgr9hPsC6vES1+YlCwLo+3SastJwSxdvHegkS5OMtz/5Xt
AD5W+2V8aI9ONAiug7nhqT0GJxbUGtdM1zjuGvqms/Inm1k3Zy9FkoaW01xct1DP
8ZqoSASvtQWrp/ruERS2C6Sjk7dCiy1HgrS+dWU9G2MxwMLZMvF6DHaJkU2OcD47
snG5j93jIBcGQRdhI9W8CzgoL2PuT13nIq6gN2PCWmkJoFkHsWOluueRv3AVpwcW
ER1rd1Ue2WVwKjTzsoUMUkvqIDF9kHbH7QGv0163bCro+2APeBOwUxg2WVuFfC6A
PaAdUcrDUWGCRWonde+PloUN/CRP9P6rEk9xtklPPu02Sbw5rM64F77FiBSBYv5o
7Pxij0pTodqM1Y11uWrPcr9jSWPP4mZCu/R3bMKNo7cXqM6nj7s0Gr1+lBLGlveJ
W2hNIKYZwGrg1FlKNVFVW8A3O3VWCiX21vpFSPXp8y86GrZ7LVFNq3x3v/ML+tbv
hVHNhIHMmwUXVdKxrB07SV/rHXweDeGju7PEhCE4gH9h8bOZW4jVN2wHU+mi6cvW
hO5e5yGsJxE0yvGieaAJhtbyUm2t4X8/V0VMePvE/lQXPcZVQBJ+mCa3ULcBL3bG
Z57p1Oan/uusIFhj4brlYbMwl4Zo4NgLj2Sq2Ihg9+1P7YiWltwBoR5tx2nLXw4x
SCuCLbMQ9opHdTbUyBqXOOcHpzdgB+Q33x/4dUb7hHWdIt79x/VdeSz027GnOgYJ
K9OKD9Ubnd00r7/zmS/BkuVU608uACeY8toy4U1R+s1kPHtw48/UJI9YzxOj5WlO
seA9PpEgezkgMLkHRoOW3EpMtCv/5eJ95CypEhJDV1WgglIPGyJZoPIvMpTR0wWZ
BknY7OiddGkDvpnv0kJw3jFP9L26iZGKSRHIRAN4kESNxoqONBQk1lwCQW61exR9
ws5C9mOxc0GSyZViD4kMiq3d4/AWd0wHLfoBGUctWaAGhQk38Xriq+tNLjt3/ljI
WuOYM5OiHb78oaTtB4eXBCM5MEzUb00jBlh9DVPmd6psrbX5vNNt0lrdOOnukbkH
BoOrd1V1C4+3tV2GTmDSoRFNZswgYiUXDLx1ns80um6CqwV+7iLqA1yzb/lt4aLl
COGEWZ4CA4IxJQ+RaoEH2WEpCuDTQx1B0kEa10v4PRcg67fngw+jg85DVLhtsTVE
P4emPLhPe/1oTG2XgNr6KhYMoELxZ6BL5ksbZnolF2gFXgFKry3qhA0rQMX4X0tQ
RdSQ8emS/A6YI6bqFcdYqtjB7fQP6BExuydfRjZ3YIkNUZ7+xyVR2r4qsQWmkHvZ
336KxmIAmAALo9CTEkxy6VjyCW0OrtfmHBLbfXe0cP1IHCTxUPNReFYqfEHEx/wG
+8Xna2PXpygoOaTUV40IhT7NirZu7npYOjg9K9LzpdXYdfBJkDw1rZSxTU6XsZUj
udm5NrRpjzDQnqnLYTcVXnH15Q2gTyAzvkT0a1SU5utcabXFX2S2+2o/pz/swJ4O
PQRvVVSXNqkrq+hgswuMvQlgsZhRBJYt/wtBDXtR4nPiEJMRf+Rtu8rX8snZx0Tq
OHGQQe+db8yevDBRcHhkR8/1VwpZzF/rJu1mu3INgtdFh88jxll8tlOH0XF/hpwL
k9hAoMYCC1mF1/vOUwh8p3zed4eyelFI77jTkP20EDumKhFCH1MzJqkPZuanCcNk
KFJOgaD/XQqKg/x5c+UZCuGHkn9pwm6VgQ86w2HGRq4B3V58qiGtp3YCkFAbhAVm
kcV1ahLq8dQHN0+6rwjVlAY+I5HO8JUQcbI7oRpZxf5fsKRqVWntQQIr/jT21/Ik
A/58Tq7SQgKDJkIRJkwKLkbt6zW3fVc4Y5a8sCscHGhhS0V4GNkDyZktU+P1XuOp
dA7nEE0NuqvfD5N4ZWYRPPW9mOsCSZyGFLPNSbp43mPMvEUn6bDUbOX4xm0Pe9u+
XFDADyp5/viN+VkyAMk/AylzSyhHXDFe7m2+dIYRkaDMolNXp6ngud+0DMzG/a0l
IlADB1Fncgw8PpCLeUq5NzDoGlDYlOnB0dS5E3H7sm0UPHjl/0mNLFHrZIRrzEAq
W4btXExfS6M6ytxq/N3c0RVSKzACgWNyOVBEW5g2l2Egm1sKQV7d+0u+ZauldBYs
U+NdqLwBAoIz/iId3G2bXjiKvCfiqM4bLdrtC7neWHn5YUbNymWHQVLc57TUtEkl
t5ZxJ9eueEwsw7xI09rsiSnfzFdPA4BnAAP7QnQtBySVI79ge7IK4NAW/jSEUVSk
8uaK0j0ZZvk0kohZ3OGp7EaUS/xy1ThYD/C+TKzJmw0npY6wNVsjsgKajYIKZpKY
JBDMgA/Pb2D474nT+yGyGqmLebdM9Quz4HgzUyMNXx1qLP0377qcGQfVeKiXu4Pt
3tOHyqm0UmRbrjcC+v/stzA7Zkr+SzGQyuF6gjWjNlRWoBPdpn//z/4ocP7GYLlI
pkTcPKgGsSjNhQ5ZzSGXqz+mMvKw9Ty/bWo3Q4/m2zFTpPDvts95DuC4krhW2ulb
MdXYIIfW9FvDEWUInf0bU2ueMSCfoLQiANuIrU3VtDnhxkSZLlIcuBur/zY0qA8X
7Q491a12lUXz8/v5GuxC2uMLjVdV6eB4bfIBx6pbHd4ruhb3sFjSBYro3mTNu2TW
qYHQb0ozMlq1vUPItWnoW4NhnnhvUBApPD4SAAr2UI8fVzpd59kXoaSQgcH0b7ZY
jK09tgWbblR5rDuCV6EQtCIt7vuoFkwJ/cEIlkLEzdjAdGaiyREfNOFlm2Yoo+NI
sqMVhTNzrCFBWaKHBpj20MxyOXVZm0ZHMq6UdFoem4KLiuaLLNsvfWhIoXATAOzR
J8hvoJl2fDYxPvbDgJrbspgBYeFHXxazZW47Smn0pmYg9QN0+pLXa6kVdSBa8Uyt
k8c57KauK+Zy6CBoqQSYScAQz1hJjO8tSHKhkU7jYI3ai2md+GSS6feSFlpbYn4+
FR4ruxXjUmfDxzh4W6sonTyVf7FQP5CAXz5s3Wp4G38eNEkNux/q9Q2e84p9qOUe
CKU/T7ODVQ8K4RRghuDsAnIMxX6NzUp3g78Ec59c9F+Vc72Eqicg2tdvbT2ZGVon
t6fw3QlAacBtmzxZh3R2XOwYjJo7HKqPyxdbzHZSdUoal8e8mlHscpdKiUAulkML
rBtOwGVX4UxT9cAClwsCxHSr8wbG2yIS1aHnvzvxiAzrp3R0kqKnW8827ZT2mxCk
2ay1pmRsqYxoZ0ApeiBKH6H1My9e64gIqtseKAkwg9V4DrGH6apNnr4i6kPpgpm0
J5hyFF4slz/Tmn0zrNdxhxPJuLgxtW5Eo8TUmj/qiVqF+LXQ7KBIVw2XLbEogmx+
8axCmUMte8/ljlAtUzqS9Fdm7xCS7LSM0YzdAbXPjtio+qoyuf7o1Qnsa8GxBIGn
4dm1lK11TRjUEtgg/29JNU54ACHTmadB/XADeoo7iWudyr5Q9dCKdaYSTQM1kR78
+ZHfHoMJ8m9hKq/w/HACpqEgk3k83dr5Pn5BYQqi8rM+BHU557xTQaDDrVO8jKu3
HRZJMrovYFy1RSuQ7TORWcTwHpuJpnPp8rMiIoXf74AHyZ/yguIf7vILkhJU5T6W
N0pqlOoKIrPbO0AuvtBQusOGIuHweJyGEVXO2GmL9doJxNBr8EBFlB1eekRFsd07
q6294bkMhzyWvsJc98Jc7cT8MwUdrS7yO8KPcMYyQrBdt1wYagDIlMYTuJYINnzQ
tslLHtOlDKq8GtcyAwmpRp1iBsz4TGUrsQpCUHBKkZg9gV9siGc2/7n/WVfPjiIq
4a1KH0Xsbt78G4a/F/fxPwjYM8gOXM2mGN+7K7reJY7bEzxAmkZM3IrAKVhmN3lZ
GT2YaGl4KCui/CbbRglE6RHmpbuB8Xe2PCPck+HAxn0yqVOUTWzM8bgQEtZzBK23
JFDWpaKv7LMLwO/h8CyQ8QFl3fx7xRAMqJci7qFFOqJhwwvZkPmQvxmcE6+Ooy4i
E4l6K28vtw+Li0Z+HsiFM7yEe0no2coOfIrZQQ4iH9xdoFJk/z13Nmh2PMug9ZsV
V2p8xGmUkBMqqdI7KrgeK8KUnKnx50XL8jSvCuDEWHHDbU6S+8KURbNdAG40AA/x
jUhlYP8+RxKqI9VF8RwJ8FWur+6hCtL35SEriMt1CAxQcTF8zhLzAgA9QX1gAVry
XkrEaF3iKVQ8cd1Qa8A5OkMWhBf/grNlFLnE9d+VKVc+IWV4zXQKzPEYlVtoVulX
WamTI32wn5f6qOPCvDs1msCW3l66rdGajxIUkj8BVRwhmaWXkiqMVX/mAGKV78Q/
6SqAi+PVtzyNNNaq56pw6z9wDbmFpujiBJXkdLueeN8GM+Xb2IBrwoG11MQ7WppY
b5GL6hlf4LD9mmBwApIkE/cyfvXEmNHSu6t/af6b+hEjFOcLO5K/SVY7UihTHsFB
HJgQy+FRi7EhHktDlqs1A5Au5RebcpNpu0WqkhrMf9Z7T8j313ozjWtV0f+5aACb
2nqzL6Tw+zgzEHf17OmfVRyD7ZmgOSa0tg3NYtXCFn1uFoGdHem4QMkRKzT4MTpG
2UH5wI/jCcKNitgYhxf8fAwQDbYQLxi/oZd4gbJLejJmLCHBP/Y/yU2JJUShCeQc
rpa/o3UyaYsTLDLZOH83KDDvLJVpaBlV5IfsBDburWJgU65oOoEQ46IzWkHzqNEh
ny75ieovMziIK8VQVRtngFAx6b+G7xQjDuO2V8GJTJDmviMLZkF+Vp4/yZBTAT6Q
eRpBJa23ZSbvtnpG9BDbQYlHfKpbBEzWwThk0AYsdQFh8bi7uuSFTIQIKR2OLdGL
AXHpipMDS2baGSmNmSGT/Tph1Fir4UTijjkw7V91p6zipaKKTyq0v4agymWiHiWp
lnebAUxsYDRg6s5vQTYP2ZXUYheH8tN3hCYYvbpCg8cN1GZJlr9znQWMe56rNbd3
ZZlzwVr6FDfuZ2HS5fftIt23+Jmc9rGGuEUSJVSOt2WO0/Hwh80q15pVVJr6TzBc
iR5kU7Ef4F/0O/pXP5VWBOY/BPBvErH2V1KbrUXAm2hmNXRXRMyVwEEIFs1m4VRE
HpWL3EezfoC82ebqbIzt0IYrvhe3lW1c8SjGoGj8YHK3A/0gf5rgf+VI5HZ8TA1c
mYbC5OvjRKXZWA4npgE4x0am7szuHiVJhHBzW2tQDDHM8gzy2M8iJM1wqAtON5p1
1FCNKDRlftEmIxO+kLSs0+JDgG/FBlnKdEcDXrPPW5SP7IfUuG31+I50gX/PHSzk
XxXpJROs+vGTafrbz0sO5H6R70zz/wznaH2oq3JKcpBBec+j3chR5W+uba+RsoP4
XEFpyQuxLQfWM4rIaK6dHsS6dE5ZZ8XwYPCjWgNwQTWaoeSfbzRmeQsT8ChIyYUl
2teOqiWObj5GFiJ6PhpDR/TZ16wXg3KoD+4NKUSu5/kktKqg6p1hp5UR+Q2peroJ
hLQKjt62yyQIWI9bB3XoGTbWOiyJTe25FFg1oDWW0JcAQajoXas9eju2a56MasdP
haMe1znA/t6gfB/wtOsEYrilThOPfL8TCEu74G1a59JzfXBCAQuOcW42fMKer+q9
6QcbabSMCeQd/P2zt9N7R1ceu2XPMWIf8j6A2mppMJIUO5xJhL4CNM9huBBufeXb
QKS78xIJ7DOv2riv9Q3a8V4pQOBdBgI22xHsya/c3qg4ysLTtBETJJ3Vi56Dcpww
uifKcW7MVrIdeT/hiLyFfKIIvGyJ9R2LtLKehjwWkN1Wp/KnbVImRtFTq2M2fCpR
tMuzniLGfWReAxpr/YUGpsaHB/MTzCoPC87BiiGXJJmlmYZMNI6kJ3A54BzXUoVd
jmB3DvYjUJknbYUBl8er4pMaIyDKTv1oEl1Lde1XpO0/SqstJgo+UEJUyke7O6X2
5PXZ5QV5AnS8NIp5Xz+Gtsh3r4yqzOZ8oqsoWV4Pc8d4kgSI5bhSFpUJ4KEQWB+1
CZrrDq+86aNZwff4hldxOopU2gkTXsT1fRd4tqXC9NfuiyEAGCaxCRBildGIkJtB
UWv/KpyhsZHioqiY1OEWuU3ewpe7uBrvU1Z8fV73qydak9MSGQlCPry6HqOtkfFX
k3LRxLIGViFw+LViI0c3R9VnV81JEAh81c5A9JsVcP3YCprm8lyUFapzVS0Q6oJb
27HPcWosxBCVE8pD/+03EKNu2imbSEMP68T4H6vaKrUsBVtk0l4w04yAmyv+nVuV
qbjNEZZOINoAgjASPyweSFKqzsrvl7cOTE+3tTuSBoZFY2LjwMhRJMGt8+DGatG2
fAHIo1CfRrIgUTS6tpBAQw7pSsJUHMrlf0ID6Kxu7XLTZEL67tRDANAYlreZILvv
tv37cYtpNu+c2VqZbwNIHhmH7MkKiypq8Y85XKZbIrr2t3oX92szirD8QS2AL4AE
raC5gMMRJBnobDe1g1Ciy/vxq/Zasc6zckHz5fA4xXhIKETOF4x3PJ0B3EV0D76j
GRarhLeC3MsDY1wdqFOGzP7Y9bPKtprBYzLXxt25mAGDaFJJnvxvyDJmh3ZcrQCA
ehxvo1njMylkMxmKtPzMVE1pEmOJ+0tNEt5sLFBSqEbGWF4nDXmGkTZfkFQ13S+T
JelaBV0J+f1gh5f9DoyP3U+0XHLhk3mFwGiz/bhg2h0K8o5ggg/RpxYpibM8McxX
cUcIf2atIGRTPCWw8w2xExlXw663Xc/KwBpgbSnU3P1rAXHX+SBpbleYwfjqFiKv
Aclc3UPqnoDkq5FXBF8YeXdHUNrSBVkF4MEWRhX3DQhwP2zlVbxf4C5mHEY1bHct
847TpiRWnnaPWHXe5umqgRiTg8R4ebaC/Q/Sqm1ooLVsCgEfl0HLI79hWTzTwoWL
pprTXGO3GhtqkBxYm3RGLeYy2z2/SvDosQbp8xycWTd1qo/hz4yPTnwHzpn27Ybv
iVbZUxJ8ZovsbCxn0n3byhNZ6LX96lRY4GDM5TFmfL/NYMXMvDZsx3ICqqjgvB20
RtoC3vL8SwnK5oJrOBbkD66RxEn2G+i4FHT2NoFMbuthBd9I+o2DNJmWQ92cVETV
Uk8qxT7c5/EXnEajbifouDXqSnJjTwcesqnfa+DzzH4a3pvh7c3uZJB56dB9scgi
Ri0ARcSbf6+DKoEqglnUQheWTuo3HUNhh7e2gxpFiZWXuFhMkXieQEvObSQXpXJv
l3avDHU6mDdP+/Se8w9LVa6lvMxgPwNZXARS2W+zUPyqgTKwpMBDmRSq0ZvDu5Ie
lmbUhKWzUOTMILCYF46E78DadRIirRt7enuKcP/sEzHba8XXsZJikqXjcbOcj4du
F7JFc/GRhv0LMgXYKGLq5EJRxEr5PL5HDFH96DZmsMoPDC7/YEjxuQuALMzoI2DY
Trg1RZJGTOpnmP8dtEXIN8hdn+oyqH5jaR1Uek6LNN78OToILtEiG5xpXNYOJ2lc
eoxZwZkr1jhQMmczb7xS+cSs780PmZx61ZShTEuhaFsUm/pvtscc32Tq9GEjDOR5
YA2ft1XB01tl58cGZZXabU1lwgzi+F3eCxBvKFONI4Xm2bpV+vbmFpxVE7gvEOBS
B9CvTjr+/PloX36j4i1hXLattB5tPc/Avvu7bJIiBJCuyWS/a/Iyullnve7pdnKt
TzFXVDPq907glVywwxEn+DwnDIuSMj3rVz3z1xowp39KsoAk/oEvbdTuCySf77HB
joZj1w5fiOgKZz1ePL2EQ6i5O7L+qByQbc+bKYcD+38bsr2nvGt47qDVg/V5uwHE
DqKhKhKk8GgGD9iPHKnxDnsDt1WCf+us76hDH3LznLap/aHebS2+CLzmPdoEwMCT
LWGh1pJyo1mtEFzERjWF2ZRBNlCSshZeDttAJAEnmnFTgGeufE0USleCRdpuySzT
8iZ+7P6y7bwUhK6os7ZV5i/aLx+ds9izTdv5HqznpMO65XfqHmK9P02ulsqeSGKh
EJsv56CdM+eHYa0xW3mnTcpnssoGkenQkJwA4S2dAMhRhms/wB3pkbPTjH24Xynx
vang+QGP3FG/D2jHhgXL5I7A87xUhXsRMaW0PwOFuwfgmRT+0YohM7JwzZ6P6PkZ
u2bUBuZdMaM+x+t/YhLfW4FuixFRq2GjhQYkzqZ+fH19xnH2os24qPV65JGvOZFX
8uLvxqC61PSgVlXlJHesxQI4rOWyjXZCK5tK264rDTeGr38BX951i1iIkHThZjZX
LVeJH2p5/tx4CZV6D4QQCZDAMy/wcgVSAjLj5nMsz6iIII77x96H5RaB1s6mGJZh
AkZvo/7RU1NLEhjvD8dHnAz08lzAnTOAJ9FnHcp3eGhb6srpxgpwumrHb06Uw/vw
ki8XcWN4dZvZaYxfIMsRacnb1hKWAizSZjZhmzWTO94ahmmJHCDPoIsG/D04LlOg
yH5lU6NfxjcNOCtNaGz1x2cqi4xj3FCi+PAawzyTlZ57kyYBC4piRO4H0PhkjDNd
4HT7VotSVEkMARCr3QT+xvYQYF4A4NrqH2+5Ad0CxxknUOOW+qYe6N6RJV7iCvdm
XoJjUKHpDrolKzsdrZdDkDeRu++79hWzxNcZgvgMZDyWEFrDyIaC3Kalnn5C0+IJ
lxzpjnNi5S51lCtf08vj4J6h5kK7sHkoE6ypn+UG7+11R6VlhZUJWiEmVi0bA0Al
cwS/8KY8dSJl5gAeW3jkFPc3Dw2Jg35WLIT1Ucl67GBzkgXFhJIJlikzNPqjhqRx
4a9mXGP6NZcobWRVm+85pF4xhAwXW149IxVKDA7gg5OrFKU3/a0HJ6gv+Oi25XUD
BKqWmvk2mRPmQ+kVzIzQeJI9SLiIYz9v/IOxKhhPtSROl5QCXAfjn0mSnYmxU6WA
reM9SmAfVCcM9FxNtm2SgP9yJAyyUCD8URYTyQCRCMfp6SSyIRBLtbFAitTmtXDs
2VEUwA9QrsNRubMt+feYQNZXnJDy494ILOTaB+n4ZhM9wcFWRXGe/58qOoc1al1i
96RwwhgFKGuBvNk3BSy0GqELXFQF2L747tz1EKdELkEwPzr+rdQvnETJqndKWZWJ
X0EkKzM3qn9W8/taVKp5OebQ+7vRsxL4TuO/oy41Ib4t69YOJDw+Pb38JNvSfhoZ
mE8ICqshKnY5mGQkI7w33bwUjbsegeYOd61TYjIV64oUHtZHHxaL5vZdBektPDS0
9h7jjQNruakgvdz049Q2Tdp6hgqc9YC9u7CMBZVld+x+/Z6ZM1/hs5jdEtdehNNj
8jpycOy4EZO+eynw/ZzsehyK6xe830GRYiJWpIqqhIlfVGJrdunbGCVFkKNMHWcP
gKmXnp2S+kb7HT6vNftYzIBfCFnof1bJB3PpchH8gcRVD9YIXRyte/yrrj8Jq7DY
ZcxAG/g6RcA5bTHo9uQok6oF/myXOWrbq25FqQRUe4Edk6BT8+MBw0uifursku/L
cUvy9r/nSIUzu2wVq4gHReTpyGm7qkV1G6Fnp5Fo+9Tx6qKdenQBGnGN4B2awxxs
ap5ipPvU31vtDX8z0aIptBbJpkKw4j23LzQAZbd0HE1OT1Cy7xc1+BM9LwUIauUR
tyb58275246TZrhYkXqP63RAUPryWT7pjVE62KYOjLxUCtV8+cCZoFjj5bq+1AHe
95IEzffS9FfmR09LVlBXi/9UliB80lqG8kjPG6mBUPo8JpCqQ+Rsli8J4w777WVC
NJoslTDuG/rgKguwrbTGPNFzwE6KB52YDi42nRH3tBkj6KRnCVwGz/cyvgRwCSwl
FZ1yWdzEPzrFRMqswQkScmUk1ECJtT2me/zJJVBUM2WHrHcF4nwqCS9VjowRZ5Y5
sQMWS7lujknt7fctizetXOLte43N1v6A+RfYwMbvw+Ao5w9gkkYNII/5ULoA/XdP
3wta7wf7xGrfq2KPcZe1wZ/L2tuAE3DlWRYRNOhDno4TF6D39rm7X6OYqh5o2e82
Bu5yk02T4bi7qSwLofBxHS1nhCI5KZGclNbzkPoFTh/JZEz7vE7p8QVMd7o33TDN
7WYECnR+x8aIAAcUPGTkPg+n93FZo6ATYU90YquE1+h0AbnV3jb5iHDW2oAa6PwE
0Fu0x1OEwQ/cGhNSbEXez54Qc3gyf4yW10n8KazOubyurKrFRAgRQ+zXrsueFhIo
OGex3ZUo4SA67vi15FasHr7e7ir8fcNeO42k3m/RTVWJ3O9OJ5TU/YhCVsTppYVh
1mq21yj2b7556R9mrrUazcWothqX/zURAcsQKeCPqJIdt0nvfl6qoB0peu4blqJa
Z/x19LGFn0P6yeJ467y8Kb6wM2Tre2ACOZ4DowBf+t8gwH1Y0s00G18c1FTZwoHK
kZNRr4pmbtJnopHp/TMAgK9Q/+iA8lrRXwuc7XD1OCDoAYftoxOxmfqkAvSMb0dO
9FjMHutqyHum9/xasOjc9kzXmEBKbdPJHR7l+NVUzevMpI0OVnzU2wl1i0xpdwNT
+5/KyAItSgMOWxOWVHVPwNcUTEDSvPjKE+fS/dZMOdb+O5NEhv3VvHSuWFe5rVK+
CDyF78YB63Gfy7EpJNFV3cUG+KEOHQh19UlKHXAAyF4otWtPTO+PJGFWnvDRd1Oa
78KLgVy2l8fHhP4t5jZjVHGRTVk8td2GSHq1MNDekeZglDBhs1A1Fajj0wM2KE+f
8ZIpNFqrS5DmRHlkU9RBMIgbApfwzTjV4Mm/1LbqjUvdOcfQ5YFf3Pcrd3cyYzBJ
mIpRVwPG2Vw1UHvQAVX3K+SlJcnayr4mDYpG1AQ8iiD1n68jeLiSkdBGzqT1vkXE
GmEGG+dnaZWYqym5va3AyxVM/jmkPClndWqtrmVi1WGcoiuPpAfndoDkeuKOTSMu
j9AjAdTIiyGNzfFwAbZV2IRUQYMyB3RGHs0YsqEnzyYaFZLoCcMuau0eh2p+oFUu
8PQpYhR02nBelMm8dE+wY46n0rwztM7fykt4U1AoWxfYkvOAxcUs4PRlMHKaV6/N
zpYPdyXvLXBDWKUZq2d5dPL4jPjJ5WsGbkqDsSEXJCSqvDJRU+zqqiJ2qwEjEkP7
LH03wdeLxT8kmdShlnLHOqIDQsYBAyo+eUXydodD5xspa0hVZiEjGiDBAyrZ1wZm
YGXq6/4nC6LGrX3wJStmCWeIVa6QTn9BlnoZKehblJkVfLOF2Y+oZUta6I71rQU+
NT/BQkz7djg/EQ4x8UrrZV+OFE6zMM8Lv0WNbnKl7Iz5pfiy3mUhgpvAdRKecm5q
2KSxbR1QXcPrqZ1QEXi5j6xmMLo4YD8pAYqvV5bj5Wj+aPFSlWJ+OfUQjsAhPr7W
Cs6GcqFyZKGPWXxmOBF/Rp/1OzEhvsdM5nQEnX3Z/kJ+y/u7awP0OL3pQtXEHY6f
3CxceDOaHzMQaAjFO83CUTtuUgxKkrkaCJYj7GLBmrCY5lIR6AudjuzmGRJ6Jngf
PsXGUl/3eIuLv8HGWzVur3JL+xPoOvTx4BN24//J+qAS2dqDl4N8GUjFlktYF51x
A7pDu7CjAdjn9Ytzq3JTd5HaQjdGMVsMCPgGzakWWmdFWdrfxXg3Rr+AVvsATNU0
wAzts2XXTh42ZH7QA7ZIm+TEdSGmRwpmyxH6fU6C1+Ic5k1HyebS1tA3qGZIA6vL
5JswZu8RFWd2lEMfl0KAoqQ+n1dxTusm2cRNGo+7L31urQXeHJvja1H+sDCgp+FQ
LsiIl7T3SHjyH8r9mSmz+u/N0ge5RTwRo6ObV5hGRlFeVO7W/fmO+0VWG9o4Wi6j
8VA4jeqHa0Iuy0FvXJst8eIP9nsPz+V9cGntZ4kpy4lweRtqXzwJwF9RnDVH+kmq
YXFaN4g1xzxAdwFsC5P6x5L+2N5yUIFKk3neZFfkL3tDM5cmajzI73WSpc52xaL7
rNfRygMMAIsaR/46vBWy8VTdNjMsZUk2/u5UN5rRf2QqcJgvJn3kDqXVEw3t7Nkj
RNYBpJxoZgajMemZUWHMrnCdBZtlTJ5TP/ylal174M4e4jCyhSGlztFPXIcZiBCa
AZ644dDoaHVV2hUkKW6gDicJIgkd4wAhqLIjRDOfv/npXUmJf4VvodLtFiU14v4E
c7x6fdxr9tJsEIB9ZH56XQdl2bgnUUPWc1ZdLCGvgELhHE9sxcrYDfp3wwoc2Mv4
JBjdWswyVpnnBVEgSFeH7lapcLOpSipLKlqo6Gv6A3cUkZ48y8Hd6giIdhSsYHJ7
wHnNUu2/ynHzZi83H8tmgT+aoA2uhXBhx6IDM+6PW9bCu8nlCfmvEgsNHOxskTAs
GKRvsSelHDn0NVdulJRsz1E1xSDrQwVCTAMn9uhJvemT9jd7ArEZvTAS/91j3ejB
ImHYrEkQgm5GqV2eUAyLK42Pjxk3VjS1YhkkskeBTkRGyWU3S66nNFjeregXJrHE
E65I9ldakL9PWL/UtORzbG/U4esv9Zx2fSN2ZgGXD5T3eTKScmQ7JIpI1XzJcd/I
Y/+d2+yv1TovBEG9+sfl4FIhegUqxjiQJ9WPGkKygz+lUD3rJbXuulZ8oqy5KRLR
Dwxk7uRYBHq5cI/0zEiudgzVyWeCO6hO5BgAAA4WkoruQw6LClUmokY9dCJE1P5l
j4kdfhoNIdMLvSiC+0lysU6d/HHF2ld4az4VicPQXWUTNHUmxfssLvfmXfWN4meD
80TGL/NS9rIHKvfcnKhoqZ7IaQ1TSwKH64G4t3+1QGHpOLj9SItL85z2IfziUJZE
Xm2xY17MutkJYRCxQFjUQWIIwMeASxp3vJom/H/0Oz/QLd/pp8FKbL5zpirTlG+t
/pXNb6dDZ2Yvp6X7v1woSrhERotibayHhMZ7r9M99sBeFJVxB7Z/s1wcMxO0PFaQ
wQyh28q1tnWEmc3foboYmlDsvd3019uhJzwqBhKlX3ws5F5nQt8Ph8PJdQ9sSNMd
3r6fwLWJ5fWDDtiuWvup1xuXjYowtXxVc9Euom81Ttq+6q9SFoxZsyC+oRZ47Kma
BqrLQMVszLVfJx0SJ7MSNYVg6E9AH54Ipi7EFwRh+g6cPvQBhoKHqF0eaX2KWYRq
HY8q7Grdl1NmA9z9fw7dZ3J78/Ph2G7N3uHrkmYCWnbM4imSYQDNNtUDQM2oPSa/
v/Qbu1E4Hlts6J4m0VFSz07ghxd7R+/NouVxkX5y26w4ffjcx8gYZY1jzdSVkp0h
bXWTIKSTE/1MVqNcjWHzTO36eLF2ek711UBvy7qvdW4FZ2N/cWPHlpRIWErHHFOl
qUwwi2FOYYhZc143VJDU+zrrJUazhzBQg0U0xjV9woGDz/7DgSrh1fNi6I2h8LCL
kRAE/QY9BRtLCa2RTO3tfvTRbMftj6yJTLDhGI1M79BiO6UkdIgt4Nj1QuoHtXzi
DOAagvceUPKTdkhKyzjk+/wYScQfvB0KPGVHVMP9GOrwjI8Vp8dIchE4d2mb1w+i
zgWT5GbxtzV+JGyHR63FgVq4xgexw9kGkJQq4Rfrcyzgj79CJQZEUyEJJzPWyQD5
bjMltM87a+X5bmj3dtOfJkz2+VOXvShHTuiZLDLnHNn+clRvOX+/ZJaflNFYWBYP
qfATA/Z6SIZy+VsN+XjsHyEmphpqM46+Ydy/cd6rBadUbcl7tKT+cAz/GJx/wyST
rSM/wnvvGgb7aeDk8FwAibJ8s92EILuOUJWKHd2cXg3MahbOqbbGpTbr4RjMi0Xd
d11Ow3BAYosqOW16PcKEVV8ioaX4Ibginri0yg9nqd2/2vvRgX2sd4x4fh82GCsy
yuQXK8BBhtRnCTo15eUiwJkBwjxhHBV5YOUuincU1OWyAU5l6v+dHwJxFlV09SP5
0r9ewZ+Jgl/4tKTfEQEdetrpY9qR1F3nMRpO8RCHvCrwo4ZT6T7lEi3b8oHIXYD7
eN92pTXiDpzj5QRPLs5zX/FXfSn0YClEbdAvDdeE2Gtx3Iji7z2Ir67uy4FOTwEJ
TCLHMNeMczU63Ig/12bNWMhMmAim5nAhHlEZzNBgFwyntry+J3pu0gVC9lTjdddu
csYA5vMsUJWk0cw6c9BTPYb7O4i79dhVEHi+rsETQlDJ2DfcXN/fMgvJV+9KMBTo
ICmmjgNC3qRCEpQgR4BbLT4lc6SCvyrpse5EmRQjU0EfOFbEFYX1+3O5ka+KoeYO
KRTo/w9ErFSyAFpesxV2jF94XS1y0SvdHSFjmsmw/LYIaaUYdAJ0nEoRxIgTvF0C
C15lB79QatGommGG9yFm3b1Dah4yQTN1Uoy0QX9+X7gyNIwe5RmVEBeSHYqmoiMo
yc6NY2WHRFGjADPlDHPOtT36BJnHj43Ad5CvX56F6iFd/mrUvmtKamUxi/QyExQz
BGZgutSd26kizCLMHdFJaNW2a9ixSaEMGP/tR17CVYtWB+piM1W0zoYnZ7coWghn
ojIx9mRcESxcc1efFWOoZ+1FXZlKjmGzpoi+7eJUjIC7N1I8RYoFhdQDY/8k5jIZ
N8V4plvV7EXp9woGzxqBWDYU7Vz+4mepLMNvuZrn9SqhBPdAQKcBAz5kD9P/LKTX
pg/FmdsbXqERKd3CHIHOuGGqRMKPWzsNlWMcSa/cdv51mlDf9yeZTZgfSOhia4Lu
3E8wKIwWkCPQEKTdGJq9I5agrPukSe0MDyy+Zmjf2nBaWypqv/ewXC9LU5rCEvM5
D45CYkX7NYt0eFG3o7HAg+Xq9FKxIV2oMXao9oSLVD7oK7AQQPHKHLJSlyEgD9O9
hrMQ2SGxRDI4yhHqcu9ViFMiD/sZLEXQsMZOEbNjVww+4GMuOClCfYnz/+fYStqQ
IPOQmHtJPov1FGZ59hSlazOTwwLsu/GQjE+aEpjvCLQrX/UtiowtDbPPM2k3l44+
jHJNV4iARM79aLMZLj6ATOlWINIudbQRAXO/AZqUXAyTAz/BEEn8yqnL6M1rFw4F
hDsDnV9TDQmmWULzQTaE4tMvwzgO9g2m0yvBNVpwBe9rjQ4TDxypdB4d94BBF/Rx
H+KhUq79WlxClJ209VOlhu+EGZjD6d3U3KO/fASujZL7LHov2Bt0GSzVl4BJaP5k
9dbw4dvobKb3VWgBW7Kr9H+03m/suft1yK12J56Izfz+wrmqSmbEvCghgHXuk3SI
AHz3Vwc+06LEn2bwfZEv/ca3CayVkkxXkMUqNYM4b5Q3G15i3kgPbuE2I3GRJt6j
CzpPL1emd7vdVbsttMCe8OlfaTF+W2Mj6n7Os7/ggTFjU9aBWJzKwPgdSd4W20KR
UCBZnawB6Yq5txxJAGZ3Btfhhn5jotPhApMpYaX049q/GOO9eKqIEEjyVXoqyNNr
Zvz9nTGdlOJdcuzUccRANz6qINz0UxEmsxbBD4Jdfwl2Z4QjDGddQYLFku6TWjei
k0b5Vgn+IHhGKzWnXXoD4JKrGByg29iQ4DwgGYgcjKgLDa7qyx0kLr61hpJgXMqY
lcfbaqPbWmGwLW5rASZAep9l+JqjR8Ufp8e1tfyHElYu0C61AVtuSvCIswu4+5Wa
yC0T8ie0yf8ufBJ17N/JBvMFk1aeoAnTVKFQkpk9FQRf6UZblVLqAhxdgmUV8vsm
HYToOqOrtA1Vt20eQLK75k/PS9/i0zJsFoF3x5Rm54m/JQDgnpAiMKKW3wMkD+OZ
hxx9o053xkg/zFxy5vQajaIs4LObg4OtKe65YISCB9SFH9ed13V8b6OjkoanONC/
8lpunuztZBQbanMpFbJVWu7IjYXmpySV1vQcFxyxAlfnLcvR1hZqb2HcDxSnlcZO
5H4SiyUVEjwDnQspt0yZXUvyWO/3x6fKGNUwpMugzmvaFwJPcziLNWik2MjipyUR
MNaWMtWjuYJeHR4UDSysF0aBQPCuaQ9aEkUKfv5r29gP3wHadYLoNaASkITS0N+u
0syAM/wS97krOaJpxpzHp8S6lHWFHQ8u7iuD1nQNf+66dtsakV707vJ5lsxBmM9X
3tI7sp7P1jWBw9eIL0JcPbnnD5+1n3a7Z8yzMlzDh0E6Zm+4O+X9UHVbhmTFlpnJ
li9sVnr9D8+yRaTbaAkQYxl9g2kHkr2qNwgBD3v4Iivg+46akYn/GoYiByVHXnWZ
4YfEzaAZ4B/I9/VZI5QWA1p31SjS5VCMGJ2dIogUfOimKPWBIMudc85MgPy2/9IU
Csi/GZ4BG4FKR3S8dF2uGMKGMjW+9TaGomoX2tsE1ujFsRkOzApZtftOXLVPmlqa
u+n8HRqdods3THHcODc9p2Gxsfzau75j+q4DicLLruKwRyRNvmqA8QsjXdBHexja
1iZK/dnO6HA3G1xKY+SbmtzYdhIlSdOisNz3Sbt0EPYuFvS4C8nPad3wW4LFzYhL
+HXKpJXm8SwwO+bh9xVqStzGKPdaM7/oWAaPxHOp+C0iMM6qprNTwdBXqH5+9Rzr
oO21sTo/G45J4boB5OfTMSdJaCFCqKD93h6QnOF5IXowopFE4Agq7xT8x91k9qC6
ouaL+39jfv2RoX/NTXxY4HI6ySnCPDh6Kvqxd3xmoFUkJjjK8UwdZY6akd13O3Ui
91f0hMcryuvFN3zbCRUR9GjQyZ5GmvajtRXoB9Xurbw2/tVgxD924m3gQSp63CKv
KQjZQoNqXbRB3EyBFQ4A7YbLGqkDAL9YEnw40t371F0apbH9mXkl9BYorCCP19V0
5C66sSkDsXW27orCdeKKliLlNdpqvKBufB+Mhq/8nSMzvl5bvgoxGi4XhWKBAcz3
uS6zkQe3MwsqimNmIWAQV5ilNPoZKi1JNk6W7XrnX04NHjc6Dx2NReJ21XvOpa09
nRBBrpKMNZB9Thdb8MIO6H39YM9YB1W3Awagyc81cId7jI+u94kQJ8UqRTHRak/F
R+uqcRVXedgRPuFQnVLK6o5wyz6iDUO5RXqr996JxFPBA8DYoFkumCqwytxKvlXy
mvsoQwS9R+MXisv+jCNc+R5JofMi0OP/UsB7zeyoTCtvWtBAJQi6La+ld4B08QhD
G3vrC5l7aDRCgieoK/FfKqrCveY+KBt9Rv3XbK3835etkJ1G2iLZeCnJqrQcgsTS
HyolccFmnej2BScZLGHPuEmViGISiCsfMu5UsJ5maQdBlJDqbwXZBCCSaMXJ1FgB
9JnWXfV1YgtyUpx6Insqrfn2R4AIs03xIBeYGNtx3GBosNgrlg5HgMvaYNxS5+wd
K2jfmMh6Nv6Ae6GboC+8abNwKA9zV9Ax1w4TMOdaEYyUXUNDrxhf68wxKk1Sl04h
NbNkRPqCMdtQg4i4Xutzd8RZuaN5N/ZBY80rK8KTH1U9l8or1IlFENJzYmmXa6oo
z1M038Eck1l3ildllqexm0AoWmwiuhctlwG0xl11b26WhRIFeub1VeZ2HqtoIC6U
AU39pahWnYnPtN14EKpTQzifg9yV7fdrzmYHaDnCSwU+OhOsnCKp9B1XN5HIFlVQ
Y6E24rmmCJCaTZcENMct95ILe4T2hBfC0+QH0Mv47pYPvkfO1nkxy8aV7hEVRln3
nTdmjACIzlWSvHdYvQTPyRHa2/1vgzbckhIuJ56b8gCoMypHHBhuDwLpNH4EAvFk
LAYZW0YxLRaTN4iByjEESQRdCDId+CBnathasveP4Y9K44Pd7IXyW0qf2ycFObRt
cqvFxyfmKvBHzVuQP7jZRbFwG02fjAVXGtKM+7HYRTTG7TkDf2yb6wFp9FKdtjEA
Uhz47jB+81uqHfT64TETQXj/H+7xEKugd3bycNbIleE9PyyLlwtm+tp42axPFXFN
ayp6mDbwDJtfCJpyWGbAATRe9tNENLb2j6Do+t834vXM0MkGdqpt1CCfEPscWPrA
jQw3APXEs/akYaw/jR0a+KblozQOLedfD76nMbgDRazI0I08GwQSAAF58h+7f+Be
eYeqy3/LEs9USdClesO6mri/dZxlqjYLBCE1FI2g5jy9qd9N+6ykEZ4SVXZE9kFa
7v6xdXuASITABIJ9biaNZ4AN0kEzJ4oN1c064ST6PuL2+JSNQyf/wLseGVINN3JQ
C31yUWUg4G8Hy3OcI9ZhyDJ4UVH4cRXC7W5zJhRqc7voXTJp2+Ga64TNM0IzT+Iq
G85GXzs1qR6NNMLrvIV3FslEzTvQfJmfXTQycY9Zyo/R3SP4RqjalOx9gT+gUDA+
1ql/rsRyQycs/gCUr5EV0Tf7S9k9XmSe6/7SKA/AXYR5yQu+up5WYIsL8HUSe9NK
JMado5ZKjnj7Wl8wZYeFaOKCR0oOhjqO2Hk/txcrf/wUK2+8EkklHiySkIjk7Hjm
MafWL333B9PyCpSv2q54EPmCD9USVRUqEa6su6xSK4CWliwyTnTAr8b3SFR+ENrz
fJNcljGJbEuAUrGb0/N3q0QhQgDSiBSopOU8eItGk5h48uDjbCp0QA3Rnt6yp6zA
n5YUDkmsSHu3+Vjz8liLgJrbZXmVoZIZt7HhWaTzjMWGytrU6yrj0p+cWueOBzDR
+/MmOE6+FWrYxEa/hZRs/iWGbWAHJ2lpsmD/kM7qG7naonZWZBxlKG/M834ZeDZF
UoHxXXZnZrPdw3u9rRgIkNnwOIySs0n1Su60zBNXwB2OSPxgxWDDmBojYitHwaCc
YxjUPTTXaR+066hEH5Rc2t8uL9NH/rU9BMnVwNl52yPmL/ZzM/KgchkEcqaM75cL
RmzOV+4Z1rd0QwZy7Z9NZQbPHG8+i6r2Tk2iCXQ68kLGZAtpgYteJJB0ARrJoXgs
nIA7IHDatfM/iuvDdnATX1XrFMmfxYoV+6iVeWYwkeyCM0cmBEWV12W6lK4fTjIg
AxVhGYsh2UM9d+hkLswIEqJTEYR9qrufqLZfu+YV1D9R+xEZMGUd9GcRjLGZ2BUW
MUNSkFBXrLe97/+9PLnOkoe2DCb3u2RzMuBN/eDtgT7RzCm4HdJPpPqyl+/W3yL7
k2w/V2Ipn8L5T9d7MC5KT3c2vLQPA348kgljm9YgHuob8nPIwQqkpgPlNBhaKoYP
thP8yGTJvZOUqj6k+w+5oPp7M+vf5bryoMOvJbV62EGhoy/WY62LM3DpjM7mDYkV
uM6r6VNEFvYHU/5Y0GjbvmB5b8XeuHM6+t13AsmxfOdr5ELUzY+kM3ntrsJRNSDx
lakHCJvYkMiC8cabpoxOf1Iar717KpqOFNMzBXy1wBN49WnJgJCa/LDMuh3kBwDU
wnTzSept0QQevWomQj54rGWf2Kg3xuOxVsUYm95XM+2UGznJsQq/8ZstjMLqAXbZ
/DK52xLAyqbsC/00vvmt9zIljGn/et6E8EPh701Y3QdYYTAk7nTHN980ZKVLB/xc
PIT4RKH5CZ6TvXjI2xswrw2naTCHGX3tZ+KDL3CV3MMT+0Q34qd6vX1XMiGD+ZE/
TfeZ6pz4kXmGqA7SlWQinqabqQz2YZo5RFddepctgoI3WmqEj2cuG896vUo9SHRI
96XQbLDH3Ms71OM4kOBdN75V2637uHZ3ybExO7bH4tpY7mqBE5O6N47d0oWYCrYZ
2ksv4VlYpYeguBfRo4v6Wv2/1LhqdZhpGDNwekdfcFAGRkBGVLgiOTeZrTwtRiUl
FUBB4ghxVnuFLdi/sYvMFVIVmHtlhchFnwwDLP1ib2AIWQlZlzLTwI/53x2K+5SW
Zok5GBdP0cboti7jQugQfqj8EdKfIGKQJs7b3pGUBmuePs0xD+QFmc3TPLhSzhx4
/297FsNycN13paWCSOKzr2gF4JOey18hznzn3IcLA4nW4258+dYhpx5BSOxHAHrV
KjqsujASoGivdpzVf0RV40jGemizWn3VHmrdEb701HDpNuf0YpEfiWMfwDVKI7xp
PECDVdEO8z9C38Hf/vZ0BIWJkzGLQZoPq6fErj/v2zqAliaeD9HwxAmJntdZc3Vh
VnizyQ0e0AFPMK1z+Y+JDoihTbhAOb43ixa077bWJSZzzB/et5XF2PHufbfIlv+k
cOfCFggAJVlQhEp3NFN2YQ5ViJSv9NnG7OO+bd6bOKQzLlI1vJ2fLPFpdxaF1p7D
3F9pxbby78izivwE5yGmBx9I4/jv4tOZ07hoS30HfPNRtgEdcaZ+OuhDXU7Z308j
vV7cm9kvXROpBGFgdOxo24OxsMqIiBNpwAzxO7jPjHc3gruLPn2AAzbfDUD306IR
t5PvHC7WfsCN34jfodnl5whLFO1OKUBIjQZbLzKoHmXN8KneCKstUnD/yGB+lIrl
1ped2tPrahYbYIwMLqIFpsvCvNQrOM/f0Vv5fFLUADj4lBEm0epaDiYkIu5j0OJq
OJiJz9f4AEO2mAtSrD47FpX7HrViYwUPDOh6rDmarZw7MMTtJji/EJjJzww5ZZbR
h/s7D4DTSWtf8ijcoc0JfvemEM6cNzHG4EotAGkV7LkqlekDx0Clwj3/UFvEM0Md
G2I0LsMHoJ63nMKvl5WWFVeNmHh/MBZURHXkDICx58L+gIsC0Eh9Ds2NfZZBK/0e
sgmFCw5p9lhSIBS8T3yRdPEsXZ6nxGh5MNYbhqo9foz2yYTgjof5AxA5P+G2O7Iy
a8b1qiesYQJFaL3zwUXmH3MkRst9dfnRNFdUyAnhMbmTAcaRNDfx4zuUhFjl5dkU
F8I2t2JYW3fEUWWFP53N7Am4OmQlE8nmQnkSVrouhQhmi7z7vcrpOev5HyMMUzOb
7hHWdTvfgts0RltzqjfpKUIDvmVoNBt38Y9d7sJPOHgM9HU/iu4NsMysF566MARQ
qw7U2RRKmaraent33DRlMhwHPQ+xzmHV+rJyHF5XV9mtDOJtfhc/E+huXxb/Z76I
kZvRjFHpd2C9IOyPTXKDlPrvzErGA1mxufLQac41QnDBhPBbEp0PoYemiR5Bdhev
QXlAAoA31OuF3jntQt84pR6Vd9BorYlNAdUzo/6csLiT4u5S6JUmDvCNEUeHB1V8
DtaFRFJ6hAKJ1c7a/1xcEmw3in6zDSvSpD2sxZadainkErIrQoXpsxyVobV7dg0J
TqHYyW9FL+YUrkmGw3ntavMlmG2UmpwZJoVwcBQTEfqhPDIV/gopgCXe+M6eAj7j
H1BDxGYK4q5XRzO8E6CvWTFm3RZAdWD3bxqnm89xhng00UL+/88msblnKA7gm2wa
4gjwfqWOp6RgvQ9aqvGBzpxKIgBId7reDr2MgFwRZKBvdF8kukZsX5bt2FQ/eDsg
JPv1995zcMCTGuudnvcP1rOl1fdZA++dDrR3jkNLEtoqtrd07b9N1XM1W36Jkxb+
9CPRgzootwbBzPUGqBUKf/jmNSaD0shVjmT0WW2E+Bc/prhQuv66xfbyZ0PyGtty
gmN4ZUpdSG/qTxpTj6pK18IqenPgIbXnLmrtmEU0u+kzKGkxR1BSQyuUFZEHsvA+
bV2mBI+5zqDJgKbyVbgnpYWOfjQFDkAqBroOEFOTRd7LjtAZWmuOniHVEVN0ANos
KcgnBebrhngEARwb6Ui+uSofmB/j7m7MeoCkzalH/xxkjt2GkiFunTLPx4Lw2WG1
IK4SKMnvKhZmH9NM+DlOvPHTQd6H4HTn9R4y61MhudRjLnC21pt3P6YDdeDOjCVB
WKUGYDXemQ15VvHzPTvkAjiIfkJuEuemU2PODyUGJR4TO9qo2w743/x8AGdV4GcN
pzJruQrDYM+IaOHNYp+c/GgK4+lKFTZP42NWDBLAuhAOSKWo8o6bIBNGXV5OVe7y
BIFmdIXyy9ExWbwFFDpgc0pjS253h321ZYTbCVnP88OEGXTn2rOPe7VifsnKpzrA
S6xV4tqzv5gnNAkB1x5apmIthAhRJRAQPSBspMv6XINQVVA8cuf3+GKtwTYVsbPf
Kt/Ahlhzt6QxJEE9HjEqpVmd3T0zGOME7wWLq4XunvhqjfrlRfiKUNVQ8kBCQAN4
Bfb10qNVmEjrWGjuK3Es66kHekkiWuIP2DR2h2xogXMm19eH0sBd7UkJWqfYAVgR
9VoM/O7b4S/w2tcGZMx8dusGm54cDUpCXM5DKa6Uc95Zjy8N9Dne0kP1DnkBMwOs
a9cEW8erDkb+mik1Ml/nJ0OwnMYur8DcW8fxgSR/wCdwksjr3Y2A4zkHSnVQgIop
4zkqgfehZKim+OREMYDJfp6LGymCp1pldkzkKL8OQJA36cdPFVSvJ4MFpNtJhwj/
ndszPlCVrvrWrEdjvtYO7iDX2jgbrUAEdDHsJGn61RYYmflTdRcMH4FNtConkxCv
xqcEjI/LiQkEB6hCmiOET/4Jw9Jhl3pUsqWb9xp5vl5PuCXoXveCvuaPpJxzJCIw
v35W2d8D9Co3+JkGYq1e1h2y3ZDo09wBtbSVKkgKfG1pPI4EeUurTN/ZUPhQe05+
KM56elYl+nDcM3FcCalvxraZpx9fMM+eh9FJ+im+OU0wJs1gQ2I9z0nrzr7AmoY+
K6EA1YkgLF9rcz1uxh/+990/4E8aqxLByKt0dOip7lPrU0VqYvBnxeMq8NRieU7T
7EIwFnE2qN2Y2PhYGH1+YslC9WEwqkvdiFz764wzpLZzd8AlUCeQI/lsRZCIjYTx
Q+LJxlSUL2dXeNs8LuZz/p7ulM8RlAIEx0V25LUsDzvgIuKWvbQu5wK8hxyur/rs
OcFI4GcF5E/h3kacNep+NAlHD4BTqVbozX4oPJk+3PGbkeUVVolNrNzFB4gLhhWQ
nxfGGYZyDX9G/oL0Ig0HpQij94RozegvwIAIXFrfesMyBP+SzRqhmhdhcisHdTcJ
aa2B0DkKugdsaawddOg6g0UMlF2WYMTPVGibnpjIje3SOzK3JJ77EQKUCcqyjR+J
HQgYJWo11SU/OwI1dzcSoOmUtB/mzWq/htN6knVkF0WKDMgbK5FF8s61AoKd87XQ
ZKqJtFwzH8sZvbSLmw3v3yt/WOmxxnSZ1aVdFt+R0R1lOFdI9nGOT7TsA/sJMX0O
WOMDouhvLXwd2UkdOBp/eHls6PrbAkZHrXVHQt33duMhO1zSrZ1F/LEvujGW0DTa
90baCvkzGH61dbB78kQpA9V4GG5v964n+47yT+b1joWG39ZeHXNEXfRO2VUrGGki
ZqNNzpzQOejIq6sWsVMPnRZ6aSB0T3KTp6S7wg4VDo7NM7oXIsOskIYrig4i6+WI
S/4zm+k0A6a+vt2wT8jMGcFXHENBJUBji0ycLneuFSHz38WdONaN1nIOeuChaBnr
qcVM1THjyWuzin3dO+OoLk/MOTRAwPcyy3NJQQJtRlkXtsi0TJCvPJ5lQHHzcSBg
OTrk7nsSybCKJlDHHZ3vLR3COA/jHwxcK3zk/PEmeNIUl87VFJ4fXPZRQYzF9Nl5
MKaOf9sYC2NPmKkQZliU4avH2kwcM3M+wGWD0yonaOgCPlnOQcT08oX5onrKVvPc
JX/aH7RdvolUjn0rtSRCf+HqInlfZXIvVcnvN8hFEqi0DyyMQQy8+sS1KsKewDAC
U56KcOIyQb5LLPvfC8oJWrVnkwbg3+0b/Fop4428ne2o2Ajqm3iTC7fB5yncxYXv
+NC5YWuXwPNS58S1Bp3z2zDUfLPDeb/lTkjVHV/378e76g0l286aIGw6dMZfKEE+
i0ViRdpqKXMMmS5P2WGN3H5zpq+kFQuwutLt0bj4jnIPaf3kfNhmatROSlZzDPsA
2X+oZJ3V4KgEHCBNfENmWgGdmWF4uSZJ3BiXZ05ho7gFFc39p+o8jLF5rboK/GAe
fTOTk+zhtpM021KqxyYqAfqsM49VYvsuQPuYE4zWOK3IoIMQX7e0Go9isNFrl5pf
nHfkxWgIwmJMtA9Mb5rWXLzu6Xc0TknW+swGw+zwBBavgVmQ8yan2nJQXVpsR0xU
awNkXnCeOkfqxoWKt2R6eLR7FUxq367KF/l7ah5wysOB8G44w71OWw5FzI5VTT1u
iAw4lFrsqKR5qs+mYN54X+HDbF58+q9s+JcvIVyCyQFofpdLJoh6hOzm0K6ZwtiL
8an3dAllbgCMEyuWdHOrU7x0iub1IDI8ud6FpmEemgB/Ft0FRWFUuw3cHHvRmWke
x51dlw24U9FW4yW8mOBnoN+85YYSOfHYyT/qn1zmDyy+4PllEl4wpeW6+GraT/BL
HolnZGL5NdMMpHUG/kkhFZXVfyRyOa7bDDcvVt0B2iqensFua9jIsxxXRTZJxpH8
Lz1jlpomF8YShFHBnwGb7nAQ6gyvRLpeszNmlcj+E2zPEw0qkTZLmnW5tuMYmbmw
GIyZ3PBdYsAMI7FWQqIG54d4ZlOtUx0nXtyTwinMVW2hBDUkFWbOZLPZIhwXNHLT
9mE/g3SwmSCgVUSbTIPAbY9y+L8HNMYKpnRzVfQkKcrkK/pjnTNmcoSBU4vIFb8k
hTF2I8hUfr3D5oOTJQKuq5ODUBZ7F3C9rHKDjmipnF1+AmWtBnLugCSTKU4qsQml
Gg+Ho+QM+K6voSb2Ka6tZqarMqs5KnHO5zLQ05zMuW/f6IqRAmMKxckbjCpCpeV3
yeIy2nEfQTtJUZ6KTZl72aPKgyZ7XWMWqZkMg9XgVFZifjj/7oqxHDN4onog5DC0
MxhXbOWQId1vDmLyR7AJ271c2GAbgDkovW7zoxM3oxzj06nJkrO822MCI4xOtXIP
1sMJQjArN5ZQ4K5J6v9wLH6mu7S2qeBWJyy60QRA7L6hZgPulK4FWXQs4OceYxfm
m9wNdgtcDnLPeLqzEdoZx7FKcXxmT9Sf+zKpPMuVATfBAd9t/6/rBMJh6AjZg94g
i+6Q3iibRm+4SlOb7sQcZ+CMzeQDkiztiORMELRtkpEgP7aE/lIV/EsUX6RaHFPE
nTWySp2CLwp4h/2ponyOveWASGMVgm5RwP3h6Whmb6myKO++TssTKntRkfR8nU0B
5S3uE2PPPvOW7g9gbQAE9Av6dkqKjAlbgsdZoamF5ZiwS+vMj7FyT+IGyLwaMtSR
21tVNzuCgW4oRkWkweTP/QaSOOGiO+zz7I/vCzsT8PbP5UQeS2eNJK8wYvT1XM0K
bdS51U7gvkKxQbSptdcP4RTNI9RNnwtUAyEArsFq/Dwa77Ybpkqu6xxVm6DCIwHJ
e9K5fuifxu84Nss3fvOoM5FdBdQrnV70x6oTmwgjdycNjF7wRotHePiG7Ikxo/28
gskRLIxQr6Qa7OP2OVO9bLcBeXXB7nIGpNEwgGNKpmKJ79NOQFYNS/o6vIXfhTfl
xId2DvDCTYodaIXGK9SynuYS5FTBzUOEdYk5mWyz2sK1hj0ljTc8mBgJE/HprBms
n4N2aHmedTzzxevEziwXFjFUlbbhW9GF2O/VEaFo58QG9JJ+uWOZsGa6QKVkCi3+
45KWnjzdoXDFmCyM0U7VudwfsG8a6RrmOoHfjxf3Qfo/At7Ui+xOk7zfwBIs4caf
c/oLmLlVBc1G5ErdCZkVOam+dk52lhr+pUbCyiJeAddShaPX5DOna/auwf9FlKly
FBHy+bFLIaO3I3qhEgI+r4kQBopl595zgEmImRCEmCjXS5y+gCHa5tGpUWkaA8Zx
PtuyT/Wn7aaXkbbVxykaJc2pgBG8LrzEMHUOTUH9WqGXHnGbo5elmnr9bHD9NbZP
6CA9CLMW96JLxbTh9xw6e+2KwL6XB9QLOkqXeyHwWLJ9QWAIgAnFdMXmPaNSiqeu
LV3gH9hW524FRbjHtnwhCaxPEO79OTDyAeyugKfLY61AFHNhbsM8cg1rK4cdWxfo
dO+9rC5G8w9anp0UF2k+UvgcYsXyKVHu/j/2Ag6MaM7In54OU1/fDgHdfAveZKi/
3qjTzqGn0IHRxGZjF30WgG/u3Cor2ITfXxXSSw+bKt6toEIuuikg4dimNAXOeRJw
9AOzJ/6A6Zynfm9obEN+NLcnnJENqnGEnXO7QhsE/uiIiQ4i20B1x9+VAW9AH4RF
v59yyww/2MF3hm6+iU7SMCjhHiE+FC4ltItcVldtrPs8XQMY5fhhkb4jyMi5Pvqn
1XSHiBQBOJ1BuLQeXFwmuslxmaFer2eBoyLbIe2ak/lmlDuJwHNIfMj0qSA+lPZ+
Vkow1x2hQGnj9vZvcVq/72w3+rgDAZW5Fb/7INX+WcguWOFtJ7m18VLor8pu1zxh
9XQnqhXzvwPTXS84jps8fbhaE9jZoX0L11ZCz/WfVkjVLaPHFzRdw3OsxTP0Ehju
9578GGmNyKv/OoMJEEnvvQprVuPqW5LpD44qeAFF06/ItvVL4EO/ZzX+V3QIrvF8
XY8fv+E3CwykkggAxlfBXeV9vMsVXCrBiPwtkmVO5HfA+WeiarhoDolB8bHg0nii
xf+UZofluBrv1RDyLQQSGydAaOKNL8JKfBoqXzRpkxs0UKj7DuD6e8gSe2X/an3h
ValmUUxU2VpSfZmbvAguwslr6dIADREKRhFHEFy3NuNLOSBHUssfhRdecq4ltACT
/6WHdt8qO2aK4ZVtqgwjfpSZLJwHIrEXyQPeynFGZ+a2xJXps2/kupDBFhsAqodr
1lXz8EWUiKTmCuAKnTAKfBofcmw9bm/ppliXdnAcuHFGvVsuAD24K0RUCBYcIAmu
d/tf/l5nd3DxCqbn7c3HFcsYxmGsZabHWbSvuv1Ld8274zty0VoLZ4anUo5p+9tI
Dxf578kML/S+IKx65PVSomRcIc0fRVaE+QliGrpvypCKulhvIeZ5ODwpSRPWqfr5
R73K8l/WhFD+Rww/bpHATQ+8bErLH4iMliaf/im0bhVcHtXnxa4QSVegIUl3bucv
MSzNHAFvK93daGQo3vMMuHFXcuzPiuUYVhD67cpPi9UpgZfOO35J0qBhFa7k755B
r//gWdEvEe/oDe87Ft7xGVOtzDaP2j66dddtAZRnIhgglytGAu9O+bZz1QECV4r5
1MKyB7Hd0xRm/rSh19moVkLosSFsGNadLYQIEshO9OuGoDLc0sh4TCDmBC/OEvyP
yggI5mBGxhzrszqCqt+FbjB6OPtDl4hqgOJgKibzLHsdTangM4GnbzPzdFTrX0hA
eGH/GuRUZmwn0rQb7ebXKz+jUD16xlnWldg49OxJazozhNtnzJ1f79tWIEtVWL2p
x9It26lYmILHR1U3LrcMHAwnG9jCmedaeBiiWUZALi+CSfEAtr43rENKlWnfEaXW
rPHj2o5wEcfnlK3EP+VxdITeJim7TlJtJmm/Ip+EkMDFSCmpLmrE0pI6ZzJDXbXN
0US75+gfwMl84J1OCZeJOxCDLGZEN+Kd6FGSEBG2U0zduHrJgMs4zPzal8CacCmZ
or7e8dmDtqvjllAp9l4PfdLZfbc34DPPDqO8lfafXlG0Ow6orFdWdZ1STXEvpTxM
THUlxYS4qx//yyfvo91+LkRP4lrZRYn6vQYc82OnJ9jrtxqAMJb/YRDNlq+do6Mj
FPo7URvj52tcYqRePK3pm/DxKQYV+Jp7JJmuqQl+cFxdXUdqV7sSsOoQEPXuK2WG
dpH4GmTzZ/H5pvXEUMT2oMkQEEUNxDQnEAWqK54ZoLzDGJqcfLe7c90KNUta9F3w
NCpAaHb+SdC/8+wE196mPfBYVgmJ/BpuIkOJ7Ze8TB1QM11N8t47RyN2baO0O81m
`pragma protect end_protected
