// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HVSRedxzrwHbrfs04/cA8kJm7jp5M1wLChmErB18BSlnIp890L9Sq4v68CPfxe4/
FbWAdmrugMAVJz9K1TT2BqOz/yij0g1Wiymtydorh+MceaNVkypa841/g49TsWRb
zo2+PcASCVYXnmYA+O4k/RIeF6EXCZfwi4VfrBMZKWM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62576)
aQqbcoNOfWu7WG3EV90+xl8SfAb9PhTLVAUcEJn2BbVriEstmBmVWn6Rc1J9gEwe
xjbMa7+kNwyaO/lMVnmQ1k04yrarIftR4AmVKK9qjA7AwWzG+7oyMmr8tSD9Qfhi
qL3LUXgtLcodQYJi5sTpzBsrWmv4S8ndtqMUBNP89/hbbZs9tUvV3aFmaZByMbOi
v4FQwuZovkK9t/6Le3FGaWRVdMDJE8+H9s7NzFDM58RVvfpEOaAeQF6Pre5kEjFK
0VGt/U5e+8EJOujg3rJYvzziSxzT3m3sCK9xQUv22VEsR08S3E6AFagAIWU8/ITu
ah0quSdr1kes9glPrpcZfx85I5FDKPDJ2dPRBPZNA4NSkWY6OTbjKnF/X6kaiMnN
XsSLOk+jp1XmSO2Zss9k3Ov1PaNrDMz9+iFkh2JV6224fxswOHhcjVOiJu+dItoh
Ctm8mVYDr8ERV02Ym2Htfd7Sc5KPiduXs0jpwjpGMJJJjTkUq3se8iNHCrcsvCkL
td3nDlqWx0dNBHf7gPwMgBex1Mczwuqz/GcX5CiFFqz1T1Iom3gwHnmBYpaxmwtn
oyH3feN3A0O7zsFqgqI0X9yUysPkH7T802oqyx3hpLFfCcWjUit6KGZ95IG7t6Zf
HJsJAdr4yN2tzCXpZ97Kp7Ywor6bUV4eQWVPopwIU1tV2NIrsNwGR7Ay8UoDX0zD
fJU/TXyzwEwWUU2c/8CQH5Aii+BIGOnahkUoi8Jc416ZMPqbQAK5xGeVosH3XCsr
d3jjdTJTIOP/q6K6m6DKna8VvtxRfj5RGUf5QmhBWN6HGsnefQXgM30MhfmgZ+Vm
cvpxkfXitrqhN+f0rV7wpDs5q+vCsqIglyU0RB3Uf/4dqxbFjK9aju9xOMOEzNsG
5f2mhfiv19CSrVy8/ATK8Qond9Mw3UZTb5PW/6V90vxNWHz44yMVWrkKSYgwBxg1
S4HyuJh3njH0dXQd2NPch8x9sSm4m9qgzRt1Ku16dfrAIr+PMMzKttBEqo4egO08
8nz5Ev3C7hs/l/+VVLX0GOLxLKnzhoLAOPBZzDW15TKJnX7vc7m84V0ndOQ+jpWV
WbBPM/xkBEuOMVSM7Ccqb7nJX9u3GU6+gcZ4PAyTsKV5WMR7sIbjGngNMOZV/ooi
2AJtHu3UWhQ/dCQzi4kwljk2GqLQWJprq0ilSmcn325l/NRlmKp0q91HZoAkW1ID
4+jbLqT0otUgfpdzdodF7zraKMTzuQZp9BEp5hMtL1mz1QAQjT+QDiFZD1Ak3q9o
V8Y3qvTjAB97c105CN7/oQ6fWTEPdmQ+QksThUhCFSD4jWj93uPYmqwXXHOmDtEB
+zhwaf6l3SkxSNV3HLJ8vXO2+8J10UvL1zHENBXfyqX7hdck/UycTq3uKr8gN7Ta
kyUgADDRDMY3vBBs6TA5Np2smvG1gh2Y3Ux4gh4WskwagdK5VYM/NKilHJmkYwyd
sM70ofvf+5/9SMq64C1mviTgvSVw5O7LYP1mVc766eK9bjSKqH4AYteTn3nCYn7z
BqRzMX/9bXyrd4DOfgNLDiP8dpJ5cVlQeIPWrFgA/oDKLsoztF12HaYsS0uenMh5
YYbD1NxMrMj+0+bN+g+f2X3iIX8pVDdObaTVDpKgP3xBsZBYjrK9+1Iu8NAYmPHF
b2R864CMF8P2oYiHg7vwEDxStw5iDnSh/OD7cLN1CiLogt6hhR8jxUbLn8s+Lk74
AaJ8gMyizGgR8gENntuWr/WNe0xNV7OccFCgD8Jfs8y2GQcnuPofkUN73d+a3xEP
BETrI/hsF7r8DyCTCJ7u8hnwwf5tncPPIDazBNn1sE+mfjwC0bgDnMeuv106ywzI
7EAga7Y+RGccBPtxuFzLFKV4z0Qb9AG54Q3tMoY7kM1U2tP21T1cTu6nQsSiFWPF
EVbt/f9XW2HLsV2x7sFqbdpdxQaq64g/3TsSjbUQEOInEPXnfgZLlixk11lcNxZf
UVbZaTPKRht89b+UdJaiRltpN+eVoEtUjWu6xs/JsM2Hn2Eza6mfl279QVrPNEcs
wKt6HcB0UgCxjuJ96bKSK5o++NexLKmMqcxlQAl6yDWA/KZQjrsXhvUYpEbx5E2P
GFkjOUByQLGYa1abBzWqHIM8smu6EuNmO3oCKoO45OQsG8WZBh4QJ584b0RApXEy
D3OGqBEVm/oVR4AF1UIuwpbxp6kbkosS7HwUrwOCeqn5bl/NU0ylGKZHwKHMliMd
VQ5dPMTLUZk2BOTBas0/kh1y4juqoCx2YKhDJbi6tGCQzZqRsGCMjLGaj0rva5bh
5uh1kMH7os3MMivzm1ESS9eL8tMuerfP/0dNvn+nmwKmMRbXSH0B1/lCwpDyAMFt
p7Cw0/3aaRlrSmaoXKdUhB0wnPLuMRCCgqD21GFgSfkWoSHcseMsCBwBf+xZfWN8
sObltlEkIYgaGgChFahSOw8g44UtbnV+6bXgTEkWFTGOTXQXl7cankn+eOqgfhlZ
8q+pVI+0cIvQxT2wlUKmFWbYmxgud8kcXQyaCLZdRVzSUcXp24SDhwfAz97NEm3o
OV18lea67sdFsgxyljmWacHI9j50Vq9TFEkmWkRPQ/YhzNWlKtnOqvM+qL+gdh0B
tv5FFG93xsJJlUllS1hkPzlFuOMaroAScuQciBWbnWevTl45ZdkqjKOkl4BaQBZV
pTFaa/vBBD+WWU6/It9mT/am9LuCxQlbRxGRwcx7D5KXoCilyrcvGwoy3lYdmSoj
tCNlYsJaJwYh3q/g/trBrmlc5xElnJCAlkVxj7S9Tdw3j8xDU9BRlgf1xiEctsE+
vaROOPWNrcekoye2dY9bzP8lXbVmlOBwFxMN7nBKLFT30gEgJHmY06B1ExbVQw4F
VuAmnOkKi89ffXp4nc0cQx3PpF3JuOUwYS5oUMrpCiFXN4rODpfxQ5Ue/wUtokCQ
pyYYgq9LoJHc9mEsgqevnKjMvnq1TPFTcZ/Yp57qN3cMufsQ/IIu8palqcITiyqT
MjKwvPUazwoyYQ/BSXmBCFmkuik9Ay20Lcbr4CfsUDxX08TTidauvo6edU5HnieF
ki9kAdtnfFbesuYclurmDge3X1fWmNAQk4JcP9cjaOzgaJJDMZD3n5Ypw3NSZCfu
Y6NwgVqKywtEWkibC+ULNPJQjOlBVgDDwKw4lswFgUZR43pIPdj/oTWozxe9KzlW
l1ji+GApua/BB35gr2Lq/AhgoGIQRmK7o94rPgoPcBS4+PgH2JhDkvLL5DuwKIFz
YluqdnBepnbHSpzYnTkUPa9eRQbABUQxAKdsxSdTUDb1BmFz9f8YJvDu+1OabQTz
8SM5w7MtoI9B4BePwXaV93FKin5Uh10hrlobTy2FOK0vJoBCM7z259nrp76vvjjO
a3DbEioE8TpD9PRKDtg8fDQXyPAzOhHN06gB7JMzPmVm63TGgQUij/fmwnEzupZR
6Ia5qfASsnHSImaAKuT1CQmSMQYarxT+hoOd0NO3QiSyynGu0iUp+neOtbVkMpDP
8FAlp3t2esmdV0KMs9gGd97PdsUe1AVRR4sXpdr87Lt9jfVLLDRrzSDwHmL7IIHn
BMaMexkt1h1LXXsObzEE4Ndeac0W/xLtHStAQkiNR3wcxQe7ZFrXd2mNOEg22Y2o
jkxhljFeja0x8EL9cFKsHYXhzKAIP5MviJESI7gDT+gSTbJvJAfyChvi8rhXlUCb
Do7l3453doto61YoHlrM9y3/XYN8jcl3LsJz+oN+6Z9JRYL3Dbn7qGQb0JW5fmI/
Z7QeIpdJwn+m5WHD7ffxToy01IVq+0afGWnzf4wrBbefWvhYeD75XuRpsrlEn+ph
etC9J4cF48U9keimKFP5Aiz7Cykv5pkaN9nbybBg9eJiinzqusSzpZnalCVcFY23
7y24kBekFfQaB1BfHZ7fGiFXdNKSQ76vEoUa28anXnqrBRZE6UhYRkyy1acHW393
hDaZZIktCPLNqIfrIq09e6BAnT3mB7Ik8Q2k2lPMvcfzcdsvnKeHF3souFH3tBbi
nCDA3KUMlePcmLzDqaVGNCeWNNXY8c+qtCcE6Beuh9xrzzEzLgNcFTgadbTJhjSf
vWrdZbjiEGukZzFatp0lxDzzYRduOXoVrFTBp9Jdt/gZSp4e6LcUKIIHayea9dvV
T0RcGkWX4aS6kBeUh24fKvUNcKx+lRflO7rVHE/PyQjBOxaNGeXJsQ3/Sz1+1bu6
uTw7SSFW0SHWDOzLz7Puw/orY//g7ErldntghmtbXsMot/HVDvrBhTLz8K6e8USr
b2eO+aQAytDmgqh5sF7bFjKYthuX0Hl05kgEzu8TmSISLRpsu4uYylGAkZ/ihz4t
0lhCInS7EkD4RFHXG8mTreLL9G04/11faEw26zAdC+L2Z4WB8jnWzySTFFY3+18l
1QEC0jAqy156G3bu6uji19p6MXyqme6qXj5mmePHgu5Zav369CtJw1MTsW/btiAZ
3cx/he0BxoTtoGbouQSI/qZhD0cPvkMKA1AfTyT4ESlL0LV3AxNG0Pe8TNQNqy9x
otesVA6EuBk6Rgd29VGw9vsnjwilitsSrfFkY/JAhaLVim5ve1zyBJfcbAJa3Wv8
EQ9G3QxK+vDK27stuNeFqE+YAQy9IcTGCE+hD6ejC/JJ/Hf2KgwEAfLJ/7psM7LI
RxUazaN/Wf0NirGl8Z4KQZIKZRKQ20EF54j4bHfPiuZFfp1Qb5p/+VpgUumsr6TO
a78JJ/7NKj5YZ9zYAMrGQd6d73AWSDW2GXE6Apvv3IE6rSAA+ep/s8MBNwKHN5+k
W2tdQO+4nY+gRjrIjFq0zPxzB0RpIoXP50hQjotGITAkvjHVXDcgy7sV5ETZxLWR
LDq1/hhwFWPaUGQJJF3QwZwIq6Zt/GI4iIe2nXUC/ZmUujRdg60wH8/QjkqtpRrV
XIxv3LICCOEePVlHHRNq5Z+PfAnAVyP9zVDuE+3UC6JX6MS/uXfrcUjNq9Y6DQnF
h5XqMxZ0eduXhMB+i6eubLvd6wLaiFBs4M/LnnbhvFyvQxGNtiYtsSdE6ArDkoCJ
4a6tYASSyGkolNBHUC/F3xBWgtXpFqLdT2zhzRWT1C2fACleAE5C7Fs1XehIWAHi
ZhcnO+sbdjjIWiFkpLUIAXX4ob6943bbOma7W8Q2ZYvohBe1VogM4qcdgFD024Ex
y1HEwyR9fUKiN5lOv+o9Czwt/DEwBqtUU5xs5Au08b7VtjRnKQn7iuffrV5nRlsP
JaGq1YP6fx38qv3VqgHVeIuW9I8E7cIoE6nzoY0w02o8L8xzdrhDHHVYGQmJeMtV
JWAs5y/IKJriA8zNS0U4qPRaFVmtXk02wbge0bblx3k+rxXXHlCZMzwJfVJOhAAJ
QdkSexFWxCP640+1H2t9CQlzQbDuQeiWRKg0QtR/QvB++0goOWvsBvpVLx3AwwhN
kAB28bLQ49nVrh5cX2lpg9u95FW0d7kwuFvZVog8VzSfZTcvrQ+D2lBMdjEkwBaA
eOqVhiaP32PxuIIYiPGwrOwncMtUK6+4cil41YAtAYolBX+APssHkct2TbEjKFK0
kK2fo+39qaNpHgkvas5fmQlqlZUGb9Xa49z66GNkZ0rosMRiMLPViNszTnk3sS1O
B/DcRhWZDKs124a6osonTM/oAoOxudcX87BZnqNVq9/P6DvEOXNf2HUNtQQUV/s7
CeS3foOTv63wcN6vCkM14CApx3VAfC4uYi39jykQGDxSKDuNeEcWW4Z8hDOEdOvh
cfij7/RqnbPaEKgPMN38ecWZn41xBoIavUPyd5WygfkH5rQv3YKIjoEnQYsxRO3D
AGpkg38uoRFgC2RxmOUXlN0c5j7tnfjfM+8/q/YJ8x2ZEzJ3MYNwayORRUrk77Z8
MVOkTt7LJjQl1qzFNrmEX1eFyqEx6wIP9AqbnrwTGBXCx5YhrfWpbB+2qXROlwBK
PBwsR+YqPXU6UMhDoh573GcQY6FFhoJMnssclBgoMIumUtyO8yWjaeeWykYhfIEB
9ED3+wzZ38xE8ETv+7YjSF7UweFb3sx0XlhCOoZzfhVeQENZ2cB81aukEkXSrDSl
I64gOiHPPsWg3iHNxBMv9zI/PF5A+L68R4DrEbBHdJOgBlR6U22q7rnDz9oSxrPp
f4KylBXpDWHkuROOAcIhRDdFMmUJYxzlNXoUR4mWWZXoTbPpWWeHjE4xaFJOonks
k76UNeccpKChlrSY/bbDKtluvjoWmNl3Y3l4oP+wDy6Ce3TT0ZWIaj+5eSo8+oIx
CS3tHc/Lj8zNvGng0X7s3YfkuFNFJgmEHj7ORS8N96WLkgorddog/oAk3JLDf8NT
1u0LvLxo/DL3BKU1zpEHDG5L0T/+cYwN+rk5i9ii6EsF1pQd4wbfF4eKpe3yfQNy
dRqGnr9Qn4H0XA9I0f3FLpK4sr5jz/gI+y9AFNnpr8CyXyOfWBBKm6jZC89GDUt3
eJwU+RluerQUE8cmMBJt6tCCli0cS2CvNvdrxvgNsO3uBt+CVY1fu38RWXbPhSGG
zR2TCiSDCNxyIqC/SHqfAHIzKAN23XBVLMByirLn0olNMZDEW/3hbUH+n0V5EK8w
TcMbSo5PK4VlD2ECIwQGDhbH1NPjtU6mvxYiIZf7kFB/0p+Co3y4fFxQ5r5DVHEZ
sw4PwWZIyhe5pZRviBhv6neqdyS73x1mtHX7+df3TOG/AgnsRUc7R6DLu6F6AHyI
FcEMqO+5A13jjCZ0c5F3windxPH/qUwgTU3Li4I4bZgEHOjE/dK17DDArZRJ2Qi4
lv3f/FpoLCr8ZNxHWWIgRtX+AQiL910J3twbxurSuHkOuUyzeoY1seeHXL9RcnJI
rI8RDXeei/YqpWPqbjittSQ0ycmAwejADNzckJvWU09yAb8eQvzI2RN33Au4u4k9
uh+PJ+TffyQcOxak8/LMVNJl1Ga9yBrY9rlq+gtvOepMN6Xj6cS7vVawv6RQQsYO
naY8vkMiT/rKc21B0VZA1NM0vzHWEsrOizTpx1orNnJxbrMUCHJsmhSYQ9O0wqok
XIDB1GHhQMLneFJr4LwEy4av83FMgyJAoCtpN4bM+A8DlfNUFw9OD1ZMcs968CX2
ZGlCwC4pc2dj1h2LcdRbICK/lHX4eYSLK36TuKhlIzCAeAV+RNlD33auzi7/iiw2
4icXv4/BKpJwhu3u1trlOrlRnTWvo7If085jOASfFVYTLj2JVUrKczww+7kE0TJ5
/eCuUIvoCSpyBjF/mpgj1derc3a9uXiF4iSJc+MI8ZqAo+9HttPygnzZB7mxftwT
rOfCpxWt2NcJJg1sujvhX4zFnkyAxgkwR/Q1ENWoHEwChAnk+9i0P926kEiY8CBC
OrnxcCnrz6DNInTmme/lZG2Ms1g7HXTTxcApm+EpdM8qito2TT5Nn/VoXyoc9eGf
XpPpmSgMGbfPHj9Jn+hh9u//sScELTojdevpo6RvF9u4a2xnbjA2wyya43FxXG81
PtHbmZUl6pojQPl8IeUCWjxkm5lDpsThA34QEzD/vDu8EhMi8EPbTxh7WZjynUNl
MjnM/Bb+axaZ8mSct2j/mjhe45ajwiUkSY5ZrIVBU/HX2CIKUwhNx8mH+Pk1cDNy
WwC3/MmS0GXShivOIY+Hlp+3Wzq3erPJw1UvDEL2GNFhDS+2PNQN+IutM5/l/ERN
OTHiBn7c23kFbchDUud6o2f/aaus73tDEiQqBpIMf8raXLmv1YQTBo2xgR0ubDcI
HEOcim9SwTFfxCCQuXHPiM5eOXc09FlFyYMfyOseENutEUV1SZjApIceV3SYk/xM
SP1dDk2+CgsAAs7FHdA/uVr0Oxx1ZAE7GCsP0rpcJsFHLW3S/Q7gCp844bCnQgtx
7HdLAzzP98NF047Ugbe9bTPyveJyRIvYOOgEEokzVW/KO1QIh/4F0qRHRY0e/u/5
3Lo+cC3UzSxUMvB3/OHbhsOY1Um2/CMFIBKamevR5L4VtjU3vFbFY6DXC9KFRulw
NuNcufh6fuMI1Gw6t4KFtqXDN2Mx9l1NRDHlFPMArV1D/SOcQBqLVHUPPuy5obvG
KpGgRXaZVtEiL52JIvbZAbpmAFBv9+72jh88l75vUTjHwRVZgpMJ4mikPktQqCX5
g3Hnx3lStLByukCeZlPDlIqfMNlMLLgebQerYBAKfSsI4dcjyi6RC/pHNHnhJTX9
VWPNT4+kvswPrRKhNLA19FxfWKrnMhHPb/Wjp5TjnF8S0spX6U5ZMRUu/DId2HUu
p/kgF5IVjE0D3ZKZ7On7mXTR7icLF+V/eSL6CN+FkepAyySZTlAqDa2R1a14jWX6
jaA7RyKl7KXKkBRJSSvzm1O/6/f31ayz6YiA0KX/rFpCAz6gLYPfaf6wMod3IO5q
HBgWyIfIv3Ss/z21H8UhMk6afFzWh3xdQvD+hxF9ylt8iVIV/g1DglPqjnMsnAHw
NiVOaPCKdXq87fnnrcR8FsYXXLMi+gOFmWoB0VUX3MpKPqOuZSuyAflP7mT9eW3D
n3GIPwEn53be/UzDYHOS23Go7uGwiUffFoOTdCaPNc3aEm/UWCPhXV2835ScBuov
1QaMwZxUuOcxMh3weA5fwqKHfJZmsxiHdSipLu6ltmVHgjf/iQCImxtGsqfTaUsG
P1Wk7L5VZIBOWxIk4MtvDvKeA5eT6giSqed5Z+l8ogOG/zV3UBjiAfnMQEC/cG69
s28elqsWjPDVAeNOxmTTb7xORLmnVyF0oziuV9klEo0lfnEpjhpeCsYu7R91BA7c
KANxF46/qEl99I3V+Dxe656V7SyJnjw44LyS15twdcOIEPv85rmI9HTJWbOa2XXa
hcWPuEbFSjPxu+FenlZuC7psODrreDaIe15W+u63DR/e78Yi0nHBnUDnWxVu3MzM
CyeRlAeTI3s/eIIlw8lAUsdOwe6nNT5tG8HzwA+o1kXTDD+KZ4yADa+AKoUkPKjV
2riOiUdl/TCAkLD/gUKjKhN0KwplMtJO6dppQxIIW6sjasQTwBL05fyFb2Shswdj
QWq5DMBOocZGfDxQ2fc0r83jb8nsLAZQvfkmn0RgtggUd5GKi6MJ3CWAbhddv+lv
iyi8QOEmkS+nZ9uRS/fx7waS8qGG87FR/ZRw/uZps89Vmwa4OFR7tx5D1qpwdxGo
psnVIJYoo7euJq5pkSj1XzYGq0izZGoJIslvTp7an2syTPs6Wsl0EVfEnauLXjN5
9TB3Yj2eDftNqtGJaDiu8HKENJH6R3FwrtxYW3w6Prju5s+FDhwMEn8kXoZWfE2t
yr4LkoyfpEu9MWI0Uq9iB+ucTjkrBtmBjJEup2xilkZGgI6ro+qCVa0GddBH/kHp
u/Dcc28p7yWx4PPWBpS6Af9qmNRAAOe1IvbIQOMGR8vfDUmbB8gM0diCLaRsTx1d
WddD0p9tpC90BLNEaMujyOZ/PlrVtC7AR/fdxJYu8IURyNE9/UQkiOjj7BOIfxAn
p/xmH02VTq3t6HgBvkWOpFiRT2pV1qpzD+9Lw0E+A2n1HAXZWNLn66hKJw1ykA15
LyGpn/YJ9RaGDhLaxpVgKv5HGktf9Jekz1SQ/TCazfsWPqp9sdc2WYBfeG4+S5Zw
kw1tQGuUNaTnmd/Q6ZAL1WXam8g0OgUwgO9LZ9UjNEplIjxZACphVY3klJG1ROmF
Hl3vq7VlWLIKp8Q7VW1mpxPPFYNvtVMN83a7XwBzHgp1Syrk/2qvLlH/M7Z6UGV3
1adBzk/CYUrW1GBPDSyWRUgOCKVXgjpBmX33ZOTcPtPu/aGpzLefAXG+FMemjIzT
FuDDfPy2yoiZ/cu/hln6CpOEZ9dfSEoRSei0WkMYj0XRcwJ3nsGu7ax0p0q+IIwM
G0tAdSyO1QWEdAkIH/zZErCgK0asP5OLJ/CQFUzd5m+mOA6RN8xXLU57IjCnDLia
qkCjd+8RY4HTGtcT33PomTgnrztW33iX0oqNw9g1dNEaYtS6MUPYXNo8Pojkffky
2OPpmN9rkBuYEuWU8HWpOwD3M3X/z4h2NPnEQ00prcVS8H8fL8uTYDvYHPXbB1AH
KGE22rG/APhlJyWMBNnFNcw5m9tt5UL2704L+nw68tZN3simaTSCqjDcAZhS1qwi
45r6kMjhw8AXygUKrLLELtNROM8xauHyBGeutqT3ZZZdEmJXqITRD5o4U+GHGrDz
2HGkS8TRaBZaWCLVJk/LHwsSR1AhIbd+bN8AkGHlANPrHz6uQtrJEjKJUD5QFjLw
gqWADzz2pwgvN6tjrgQtGM+aThKHHe9yNWXgJRPwpTBX3V/6PTjM3seCp7VHUDDC
edgzvXUvJ5IHmRj4BZ3QAin1QrdJHsHL4xfK/8gWYeyVy5/AJL16YP01mRv1Gpxn
yzHwejqG0vRx+iOcMg3UsCYwPaf0LWDK0NQn8sBN9/fulrrFjn0ATTCttIsXEmw6
EYcHwI2uXY66yf9qOvF6ZIa4uwhydAuX3As8FfxdJALGNFBBFcJVdJfQYBZeSQeK
OepS7bqSEJ2i7d1VmkdUE8H8yVc4Ujovxp4NCp9Y9nP5+mvn9umo1qe5NntR4bcZ
gKIFdoxDRJ3kItmmmPze56tnSNZsp3pw+vRcUPi/CyROMQWvQUfSmFlAWshy/VDE
1TsuBDCGTmJlzvtXpwS5BpEkc7WU7SSU6XXKSXB+vrP6n2amt/haqxSLe8B5cHGf
AsJZvEgg3KOxtLDB9rFDWL8fX+9KHOymaE4lNrqrly2T/bFV/IUiMflLqO/+Coao
WNN6FOSUPwBMG8TH4+ImKpVgoL/6NFZQUsdlBeR9ocikam7gK2txiWViY3zNOgQS
VKfgKpuMzRYdSVVfY6v0udJyyCgA/t2OSDrjJx4DmqCjrS9iHz7zV7Tar7e5eFFf
vZGbDobeh1LYl5c+3NoD9La8xfCHtZcTDM4I5OYh2Kq9BO8qUOBHAvQ6kZz2BqZu
gBXg+zGvOGFA7MG7aTwQGYR659S+aFNIoeuNJiYM1UiIiqwVCB4BFIVhfdD3oxuO
kXcGngr/gbNYwxYnO9s6qwvYMhaAy10f9EJZYdwMlOGg36ZeFIB5q8V4d9XakQW0
PVVq1uQ5iYmh2Wo1YvQ2syxE0Hdv0mEU4owLuqmxT6isut4PW6DUbOPp+bXdYO/J
Gq7TH1kZSSjQa5X589XFOZml/DBRs4v0xNEpVRt+7PQD30S6wVv135GGnDsLzkHD
lxqoZZttHDunqiJBoxUEYbW9ysbNyBZU95RXg4erBrtCCoMsUsegljp8S0wD2YIQ
tHMFqrikw1nFLzNEOGLlfk9wPty779kCHaDpQyHNR7rwn6FdgKn/zN5+sVg8vZpi
YrnDUXjm6QL9UiFE4NI4T50uVgR1Yfb/oBKzp/N3ev2zdWnbTy+OQIP5SE8/csjT
MmZfGicYEaiNzF5V8oHVQ5cVa9Sdc5+1zpdTBlKVU735Dyr+NWyTcTIPUjxpuhHn
/e137WMqIpyovzxdBbGUYQeSeUs7JFlq9EDjFZwVP0ln0f4a5cUI9v/GX2rOj/XU
1er/rXib/UhJiHWQVgyRpAjKAToAXVNa9IqH8tXsvAH5x4R2qz+hjTaJh/C+CjxE
8/kcGfev2HOEf3zjmnZAiAlz1tsHD5bDmCwcYuYldITHU7HpsUq0WCw/wk6ozAbV
RYWYr3on4qdWGRTUcawO/CGmHswVNyjDQE0o1DbcnHPsF6ze4PsAig5TyALXCkTO
RpTOMbGA/8L1z1y0OOmxx/lPFEZnycuYDZPB2oUOk2MS9F7qviyzfRXvNvyoNo0C
EgOEtARsSyfw1/Hysi1FL02knvZ+2VMEVDjdCWJXLDDq35LuY6aLiQZI8e6qRfgY
d48eiEDXI9BBLDSD6XwgrsYZ+mWta71JkiwemRpLxN3crtV/RST9ULMlzwkECg1w
CiDvedbaFkq4y1UEgriHkP04f2z3lWiHoRGbzdLe3h31qSFcV/7mCKwHmMqhOdBB
Z5MKjtA0XmIzuoO3Xo7ihHL/tfHDJuCV9GYxHlpKJdbZb8u58lV1P8OijLzH52bR
9fRBSndW06kVc1b/4A+JvygIR+er3sSeuUuQvA/S078atZxLJOfghycX50Ew2t4n
QzSJp4blM96dhifFGb1qvp1L1RTJ0IqrrfcZRgQ2uAOL7laNq+fkOPYdFKnmq870
juQt94zMxglJV5aLAGSQmNai1+H4IaNToPfIxWARV5lcxf86rDfpXzgHmeGSAIDt
0J7N4rqdkTLatPUe7pCZWT4N2KZAakNNNu+YM5kifWvz3CEDNw3CnlmL8SWrLTK7
4VYCdd57LdRorLOh1wJRaQrvQPQDiEUO40h+awa4Gi/VkH8zxyZ3TxB/UR3tMJDy
E3OJNkJr11gNp5HE78i5BW3zgdinx7wOlT8OsWGeLCaigQhDpalmxoiZI7Ca5pgi
VlzDjBt/RrnIRX0YHLf27SjQgN7lrH7XLHdyzbNnqDJF+pfTLWcWhjfwzTGz99Br
cBuuz75WnkuqkdpK2XoDAfoaAVaYE25Q6yCRnQb30mVisk2Ep1SnrxygerN3KKQJ
vV7TBv67c11giv52GBAR8j2fn7ye9Lk4D/tF28LKuLzDovkhkvA06pQMtom3goYS
Zheq7BgXUTAmrlwEkuZpoNAS1Vo0QfmF8RB0NWRlGTAG9YQeBD0YTGfby64b+6go
uu83hnZF7PGxMvTibK5kI+6IN5vMSTV05m/i3j0kxn91ZSvAQxw0fXWFJeO3U317
wnd0MCiMIdE+GagAtBQlL8g6jVJH16AY/sP8bz35DzqoVahKO99siEJTmYeFuEjp
P5NdFbm6VBZpJz5p/Vp1CukyO21PUayC5tb9cUwAyEwdHL9ee+jhFFXaVUUeKRD7
cLqIK0QeNzRnuhKonNxuwCfO6E0DjJZwP3MQi5wIv2ULHAPFM5k6lyy/tGNlC6VM
6qFk0aPSTeAbS7rR0OeL0YnsVefknEQ3ozxXEwAz1sNVEqit1dSfF0ukYluy3DvV
Rjt5TEzhySBSGG2dU+Ovukqf+hBmK9egbzc446llC1UliMXGZPnYmxmi+PFKP5kI
f2S/eQxXXAVs0hNM4tq2m6o5uGOWA6gLRQhRZTmukx/kyf93brciRp9IMGOpD4ls
tfqL+39msFHLCMjz4VqRCQFlZ5eZoU6klTPrgf8X1EN0hG7T4zztygJd0aTJo/qf
CLyYehqgxFVfgrhraxrl7skwPDUTJGqszgaNMr9tj58odX0tWvaJy6v93FuzEYpc
ebdy6Wcy7xjVam/mnoxqsU1WuvylbKrKFkEbO6g0/1hgCvDqxKCUZcdN3M4Vbymj
nTNDm1ErARROT34aFX6PBZnrsIeenUqCecVJmgqHwswoqsTBb+7G8Cqq+woEh6Zg
rrusp4l6dngRnL+OxGfI69lHKvNlHlYz31f11w2BPJtzVCUabk1VU8cUH4fvfp4I
DQjZqlbtfQel20aryFBdwsO8acoHh6MfMpg+8Q4ZooVCK+1ns05u1n/C6G/1orX6
ZmqNP2uGpPs87fBJ6iPWDyDsOzAktTFIEMuv9sVQejiCxdcFJYCqATG0JX3KYrsm
zpoLSUMmAaWe2J4Pr9nYrVB37KWsKpg8R7J0yHod6tOmLXG8PaQWNeqIw35WaDAQ
y2Nyd+85ZUBKeEfTU/w+rDUdUc+9B2AtT9WKmNuM0mS89E7p9f5mViCxk7+dTHB5
X+HpNxUXKTnH7aU95JUGK0vRyx0TS9EJf7FLUz8c93qD60pU3ZlgCdCHmuMx0oIl
iAPcDLZBYZwAdt01wiHlUF6m3ngIFxQJ1r7743x2NVQ/YrV6wj9yL26AqlJW/7V5
k/+6wNYAfnEQzEsRIh7aHfxXc8bei9UBjrCixEtSaFt2fQWjqZwnTMStYepKuETS
nOSGmNYhDbOrXY0wB15tCwrWjY79iCafAt5nmjeA0bmXaECLyN7de7CjDrbVQkK4
hV8odQ4hJgWMsz6myDRk+Dv81w0eRCS8en3HNPxyvwcNJiFWRFUU/GYlQtOXYIfu
TAsVC/JTKLV1yBsf+gje1R3MI2LLb964I6F8PnAM4/FS/bI26djTezTHSAf9APEK
M/hYIoLzQ3fBzIcprvuyPQGuCJNw1cDIn7+J6ploN/AaUoGN0OUbNHz6bLrsXlrS
iyamGYPpGgm4hD7JVa2El7LkM1oppkoo4jyAqriN7IS78huA/j8CAl8oTCkAy5l4
qizNMSwuaDzBW2KjrHfYP4hOKjabho/BgQ7o/6RkBWXHSiVCbuzYgrimseSrZIVC
yKQdFYh2t5gtucRt8rkT9AZFjIz+ed3YIbaFT1J80rGKd0ZH4FXb5/Xe9PsfH8sb
FP5ygvRIZV2PIhgY4pNPLVr1v2W7FnlqQcKFtQRt3ls1zD4qa0zTy3s7J2BYhDuw
R9BF86agIZsOLy0ax088YjHFJGo7ehr2lXfki6niis/3d7Vk/UO2ZampgPLqLuW9
D7E3JlB34LDBxnP4hU18MwGN+1IpJ0nQMgG9+7klQAXab1aHJZqmmDddcHE1jooT
xTxADZy/vwTO9JKhaFPuPv3aI0efupAhHQr+8jSJ7eGhH9ZJEpxntbsvaZ0PI/Gf
713Zu0M6uvsrRW23TvQ/XflrBMiWP7srjKn3zFTzroKxaWLCu81b3gV9hTslj4Kh
Ox8ncjC1i64tU6QTM8xfJZF3aJik9qanf3nvWLdprbkspZB2Yx/5sMzAZuFOUYPo
RjKtbCIu7qkRIegbkvIjpx1bbE0JqJCem6K5xnnx9BFTJLOd+Vdh9gzRUsyFqD19
ruAtZ5m0EIBbKa4famQgduGG+wDS7adfeYu+4//cWk+F3q95P/u+7K5ULwtxliuC
M4UJTrUfZSkQrYfIm28iUDpiR1XpE58203PXY/6owDN6QIgVq4Mm5NPXKts6URDk
IAHpIK7gyug8f12vaXEDSGBwSYLM/VWCMSsFQbk8yVTEw07039zQaCthqFe2z2r0
DlJUmQhRtM4/FGX75s6RIG8ZWyq8IiITlzae5QiuVyzYDUNcJgI9lZoe3O9lNtIL
3VqdXCl0/Bahh+/NrrF175wrAFkuIBdrbrtvbT1l+rR5W3QiOeSKc+v62CEP0V2J
t3jTpMbFWZMAIiYUEDmCzhVpepG6QZH+Au7VD7u0DYYaBdaCw/3evUbBZneJGgwq
rcUcqmr43NyUfwZ37EVFqXb5AvUqJ8ftj1oMNB7NyjBLUowz9j15XPyhniN8LHk1
GcKEAkXtF8YLJq0PaTGbS0OIuKBIE73Kg7xuo5ywcHX5qdxLrSgFfp+wkWrEj8s+
J+sqMod6o/4oZXB2JaLkUcEU3PfG1mM/mabt/910Xsa1/9ytfePIzWptAunISJ54
SIVYapKX6BkhiKcO5PSs5ZRxB8VHPZnXuRIj2JKjTc+hHagbcWIkj1PIb1NkRuO/
y30tjLXfbHW8+NWZFFzRc/GDvuq3BIx8fygtyrbepnm0dnL4+Yc4+e3NOlF4GJJ7
H1jOGWMXSW0+jsPFRE7IS2/xwfJXDddF3SD9+uqlUrdghI+Jh9jxcxbS5PV5/FVu
hW8P8T20BthZB/ei5zRmXgU8R+ZTMXFTMzqPFhIjDFo6EAoADq0MR7p0X+uEp2O8
H9HiUL5sE1Qy3sjkZi2+sE3vpwbRodAetbmR0nTuFvBV0gWMXelQ9SA9Rf4vuGwU
OkrjrTzGr2OtSOzlr4tccKghCn72w3e+qGUHYiRh6+IqZsJVURa8dWUtAAuVFig1
n6KT6NxngOn82PQZotyljeKPvCUSlp8WyD3+7+Biqpd/dHwjrn0bXxVNw13IaYkj
kkD+wJ8b+fxdfUkFw5SeUsMQWCPPQiljbqX073rjfgv9cmf7YhzJ9pWwxTrhEe53
sc0MQFpp8/MjUqKL7C1k2dDSI2yyOEXJHKvFSCd/A7crUQERi4zItUDaPb9O4shI
bfmTvM5zRC5it6xj6E1AGTIpY6J3qZ4gzHefzYvEYlqkRJWtA/HvzkwK3pD2Uwn1
O3lGJzQtau0rQtBaj+T8kVI++C37NkpZ4eSvpQaUafkD478SvPJ/A9CDj86fynW2
SRTvtPqVoW5B1Z5SMkSUVK3o5/vAx9omDP0xv2PtEpH19GTdYS25Jm2DExVCL5gA
GF4ZeEpHYE2ib3+s5wkUFaQYlauXuB8C6EIJZaJKc5i4vfLUPvH7jhS3So436zOK
4uCMiSi7invXSPigaPoPFyXS1JzMFUdRy65ekbQIgy2E0e9jQo1hahaGs3GUPcYg
VRPoSDd5w8PY4Mbo7AjRnXzKg63dB01ftZsmWrX2LbAPyjIZZZvnxMSCPzJ9ZiXP
MM1lupn7mquq8QW11xuNh/n/aCy5bfai5lIhRv708vKIPvVQkwcGHsvHyY2mEOV6
VVIGvFniB3Yh24rxoggTHkXqA1EzD8fz5JlDqGlQrJzvPtcapWhpYfYMmhFeXw8U
2udrQxF5q0H5MP2lgLiGgJmvYPbvAbLC4Tgunc8cWwAjKxdAEsqbCc3DxQKUBBiS
qkoVs/TBrV2qS2GAQErHGuZ/r8PLSdDNPATZpauaYwApdp78YM9jTTVjNZfyhwWu
+Mkok8GGS1GiPWmIBP/AR5XXOxnbYhJu8zrs14ik71uC49VbfhQBDEXkjy19gkWR
CUOyfYJQyKadzDyiN0Gs4cTRiI9vLLYnuyU8DkOuqsmGZvP6R5XB3PexHdiyVSgZ
zY35ePsYwtPzd2X1010UJTOVBtHZtMTS3w1qNyQdfmeoD9xbiB5c5FKpcFLZ9xO0
e8adUoQSNC8LscoOFAWnO/N5VqSHxGxWh+QodWPC67/m330gEGOv/2qtKA41E70J
d/Z6cOdflUIM55OwvIIr6ssFCmb1K0fBDGreO6Iv1HdIElsQLxLfMbKaSqNhodZK
NjEoM9wJOvMZnD0/0nf1sLlcwAp/dujivRZcweMpEwbSMPwQFJHaajKuyPeW8tWo
TDXOFTDDy7QSce8FGe3fP7NIhRv+faAHcLlI5lglOc5wtlCoMVFkQ03uDTF7fr3Q
yx0WUE0voJfkjOD6eaGrnMHbqMCbhM36zkezbkV1HB54YN11KF+Wh06Kq8CPUoiB
Fvrq3aMGhW3I8A5rOdaCA1eV4AunupBg3Lb19r4dmtH4dTrwFBeXXw7yC6ZVD5Rq
dlGC32dZUiorVh7q/UGD26fDBVadBLwTSjznJziEt7WQKM/IB6seH84TueF80p6w
xl/baCRGG5EzK/6+PqkEybfQ/fGeDZymLbGdwauiQvbaVjalJYabhdhZcm5EJYt8
6GS2cq0L1JUNSB8BMiEgkxUQwBOFELrVn90cF9xLV7aANzcg1Pr+pPJAsXKFCQyj
Anp1i00fagwYTvP1gPAbHNCqnoEM/tK8BoTm5ndCF1/prY3NHxWzUv12hcV+4uTA
aJowkeC7CXVjbvkZpASWzENpkTvC97+jRJomhPrFlvfPiPofVr+s+ZS/SgPnPe8v
EGjNkxOMnPybtoBCxLjp11hrwXsjC7jJhAsenrRTlUpj43D24Ri6rqwaq60uPkob
ZMZWkhC4vSQQ09BEF52/s49v249Fo+viMfOl2RDKnBhuDB3OQfyicYrlqelbqugd
ZNC0KafnEtxmJKHy8Qbi4eS9xRms0yoBYwdwrCx5O/pIlUH8HNHUk/6T0tJ7Zupv
zQegaukwA9apcWE3oqPyDrzx1fxq/AqHxl0vvIM3Q054C8F6CVaQ84sDrW9Fhmgo
/zRULJtvhIM7flgCK07EjmOGHrO8mgAvt0bAAnkv8avHBgw2RVySk9LQgZM0pREs
J7mR7Ir/KcnJTOVeAtSysCw1LS2wxXdQB7tS71VLJSNcpNjzPQN6UXfe2r7Yj7Q5
KtKW/FqSK/0oiHuhIBPu5+S/TYvplbvhOpnP2KlI8uljFj90pq4/3bomWRN0DhLK
UdOWSp1RhAEmKxKIGVc/tU2gr5pVDt+lPtqKk/crjaquT8Qi+AEHP7+ZgI717lPC
VaNSkMt5siZdqWwFkIosHJGn2wVUd2YQTxI3aCaJHXClvADMM0ie7EJW54vm9sFT
pOiZcfpI6XXhrPe3eKPuUFnGLOlDvG0I5Mk2Z7YCRbZHrXZwRLg7yn6VDEgt56PC
t6bHsyJ/OpDZueaSMXL29fTp05IF57TkxTQ3vNRvPZPPtRxpuAOSo33JYQhHSaID
Lx2aLt0ribg6KzrOVdoeKig9Vn6YbtkW17gc99ohf5EWiyoVseI4FcpvDDcatvIa
O0tRY5pQsUP85pJpmpR1yQ63Vx9ti2OtWaPFya/mITh2wxR8QJzlEO59iYxq/iOn
+JFuknTpxiOze49bpRrlqZyT5Ah2wVLoDYlbHuCCxbQaKR/Gg8Fq8q299EikHau+
pBtLkHi5GW8jGjs/7Yzt5RMvqAcPFtYoT2yQc+KFQmFiRoS6dTQTEnt0xsgGsbw2
BShtgGu/Jq7P202nxgxe59wzsrqDiKW8rvLoD1ztDkVxlPt5wOpH1OVWLp5M0sjf
lOfBOwRIjdf3xX05VpNi7GRD9n1wUeNrwG7qDpAColxNFYIBvR1+oeWS7SuFgp11
IjA9Ew6R//tEd7KULdxKc+OUJMT6VbwFsHp2V7Hos78IaTmAuGi/GEcVtgyMLqRs
7gPx5/ztUFhsgL/2aHFoel44s1sBrNGXugcgfhqIIvowKv5LPPWCobeo0jWm1IBj
NJU2M7/56HLd13MSgsMIx4X/ro9s1X1eRplWmG1+Fec+pY+Y90ZGWNNboD0d2dZ1
6HWawD1HBdgqj1wVlPM+ubB9yl3qt4qIDn/AminImQ777ssbk54Emz6konrAsFEN
A0KIsb1rxsfxxta+M8N0JJd+XNVWBy3SpPjD0GsSiuR0/2fj52UZ5i5cODh5+dqR
50aypmh2GLyznQo6+3EgLXstD/3RY8vanFd78jpsMFh4VcP4AmjZOftWcjRinPbm
MzSZJo7fjVueh8Mz775/pTmfK3K7eG60ZTOv/jy7inXCVD4WWXUan3dLs4Fevx2/
Jy5KH17DPyK+4R21ut+Ke3MtbzXls4nx5OYApp28USF0KVvCpSvhJHwkkyYiriuE
JwQoOSQe/oNx6/xSGgEg5RLhrp0IRSbi1fzmHSjcSTuBTqcyCW6Y4SKycnMR56mq
OGmB3RVIEEf/uJqzUPrhrYJq6WBLugRG/eQ+0BrDLaMkWn/2Tbuj7HrwfOzz8Iwn
UAnqgvpNrW0ghi02TRt+QH9gM0s5SJwB4EXqVEtw1yfXw9/fgDrgTM4bFUXNRG79
WLpHgNdn+2nd3vB8hD62xRHmxU4WpPHSwRCmhL4fsgt7b/EBLM/VjANsG+8W0cRS
4chyh50HG5xZ4mu3VlAyOjGwjJdq8j50kIs6g9TRgq+2uoa0d/rvZm6L4i42Z4pW
0+9rLal0z9GlPXP5z50mcIsHw3BTvxbt0MA9iqRFqKctLOjQYCNL42i2cFM9+iqu
vFlXNKlkz08itm3QvNxuAjx+rhdukdjPsK6/u6NE+JsQLphJs9Qe/1HxKSI+ZBZc
95EiqjD4UD1VjZ1DTQt1+TnkOrLGDuZ0jV4ynq+kmfRKsyURYn6MUiFczwICy4G9
rEkLRNHH1q3djrgJ5TUA0Aa9YIqrWccNVr+Noba96Sl0Dr8lmq413u4qYhcfo28R
JH+CUldAW0SdF1cmnNUUm2fzSyooRVjW66OlL/ySGUcw4U3+raobVrZArhAU7rF9
9xrnBwGGfsdDXLTmAebOU8VRpO4j1EcpFLHqPq6AohTq8FygnQZdZQpqOhe08Nzk
jx4O/gbO14M0kyma9jAylJjGmcIrean2iTiXgEU3c0DClO072ZZeIx/RrEKnLdsR
9wW2aKOQDb9plGBdmdVwHTzNICeH6HSBABHetu/olAqHc3hg9ItvMwP0LRY/ITUN
0rZSZzzCVD15J6B3yrCd2wJj7RukBLJP+MWxJypzjub6VUPJ45TQeSrVANvdFrfl
LUjNUoqlPMdOwrZnZxF40jxH35oOnee3FDg8IqFaX+3S+L5GgFXRJAn2zPlzF1b2
omvZXXybVpXBAlxzEq3/fXCQkH4qXt4EaGLN61yZvssG3GItv4x3m4GRKXyD+kJx
9tIkxrU/fG8VxBvCV5FZIrFxhNNCf4m6G3LjHz6ME5f6M6YzzG0YhgMiOvVQAb86
E9DkUX2nWQjhlziJNrcSkdlBOB90kvYGoef9Z4SpYdzQ9nvhzWuLnoqqTF37nqcx
fJW3wHO/zIjfozhp8EXrvDLs21Sohz4xjJtgO+EC2dioIWvXNccpZZNayIrQCSuC
Rs/xTw3jnGLbS3H0KpYdG24jIsNy/RXAIgkhq3NIM31vRcx6eYbeAWGvU+ST+yKq
FDPoCdkBzW1GhASVJKFj1sxX5jLb3e9gio7XhniQbsPhd1G+reRV5iXX0e4x7A5W
R2CZr+l63hDEUorP9awmTGkxiwMJc9SZRp0OjHAhe/TA0Nx7spkrt3g15URFjLTa
sh5mwGLycHDUbkmFG+Dnb0AEdnVht0jWSu2cG/MCetCmkuQJ9UyKZ881GYBPNfPz
p7t55UAcXs8SQSIZWINaEPcIVUdEQ5PAJZCw20207SijRMxYMW+Klu0xEVin5Suy
1Ok161PL2dtcALVqVewG+M3A7Kp8gWd62UQrnAds6UGaU7Ibdx7UD47O/sJSil/d
W9OOP0Mf3RFX//StrmRbxRPvnm5zqhfY+3JTrKsJx2AbYEJBPiXIiI6UyHyFlbU8
rjwqt/kPreWxLlSM67ToSNXGxYCJBZnnOio/dstWYc7NM4rUl9oPle9KG8ByXozw
lFYUJ8TJGrImf12xZPhd7h/lGmqc5gnoKIZIiMPymSee/OHEwqq+tsgqlKkoPjIX
8bTrYqjFxoyo5EbnVkz5bj6U0Ai1aq/LBXCK4Cv2+PyqFe77Q0COi+cTuGEsAtUD
KcDRiR0Nk8Gg7ISQ1fQwzguYgCDdu5ZZ2pvRTRa190AAeyMgVE5jzFK1ZIsF65bT
/K4biG0+lKfaeIx3SMRBwuyWSZFSIcsUWiWYyiU5e7dkahpHUMjbEfSj0TF9PAl9
R3zOJU6Y+B7/sSRQ/z9bNbqQ4X83/DxcIrQKSh3lQaHlix9BdghzI7DNboCeUsri
O1mIx0X23C1kyQEQ9XVVyPBQuLzYRzEfkRlL2LsXhfNyTbsQT6H482PkzhoiHy1w
ZUX0y+Fp8jkOb7NKhQZsw4KveraenpMp5NQHtEyOycHi/yqgUNUN1YtfzFfX6U0l
I+HoEa1jh+fFQ07E1P2Z8xVP2bGjRe2zISFhBj63q9WRIQRQSgo2+3Z82FESeq4w
1xYE8O5Eq5wDHP+4p8eGGRL+yjrvn9g++j8taELFFvID5qEF+eiIx0w8WXiXpIYK
pvHIzFYeU7ZwAGmw51sHWOOpEFzYkB/jJZcRD5TVqvqBBdrScKSop6du7q+6rbhn
sX9qGJRiXRJcSsKcfhIh9ax6yHUvFF8xR7+9ixK0sje7Q/EEKB7QBeAOMKXD8x+8
HFubKgJJV99I0EwWL1sk3uEnU9q5pq+lH8LAdKcvAwaTaTM2OkzBkw9OFF12jrc5
QyZKBUybuTT/s/MEH4d7XGkFmUZt8jUavkaCf6HopNHO6NGcjkZJugMXkDMHZBny
ojuhmBdh24LN6/rR+1xKO+kdJo7mXfZ81i3wGpPd5Hhl3847DVL9GcbUC07oUMWl
Mn4fFJM4S4QRpwm4E3J9jliCp4j9l+O1mld1/PWCu175ty7ohjIsdPjNVtaD81S2
FWaFdczdvB/XyuGaMLucpN6Nzl2fYyt1hxmmUyVmHk8v79t8iX4g7TbIH5UDt0GY
Sh7noiF25O+CTbr4PCiiK+vGBrrgKhMcHWk9YyfCUzKVmG/Eia9oglEJNFPldKdG
yOBRDmI8U3PnijCM2lG9tV3NXjsrdWimZ6J0ReRyJ+TrvM2QOwJ6/cLiPGTAhZX0
+XnsLPij4moUBcVjjDuucQmeq5iVg0dzvcXcOG4P5APXmucwUaZkt9MGCxECjZv7
R68/ecI3ZsuHObaTR+mEE5UswQqMuIkR6lk79b7rK8fXulDJEjVZ/O4CPwwnRRKP
L2Nkt2M5BTLemUC7lnmT+T/mVzz+xXlVINCXI+2LkYiAWK+NdzI6XULA57sZvDL+
jybgDXIY4brW78RAUmEzYC+CqfWurC5eebKmF6QEuSJvpoCf/469K+c6svTrR+Fj
//42SdtANjtm2h+nRN71OFw+vPKrkz+SuavvqD4jUsVt3cXTn8+Xxoz4NdPqB9If
yz788uuvfpF7c26Gu/GMnCZK3AIWHvzLaVj55z1Lfa9SYBYDyZT2IJZZipBJBhcF
rskqBCJ/6Ey/S9M3QEB83lfhiHWeD9V3S3rvRasCutmDJgliFP9tWe1bu8qVGSzP
+uVN7ZE37ZO9A94lGii+Uo8cXWF1ycHJEj657QjvJPmhedeO5WXDvesg16D8jkk6
XsHbINlO6vpYufAteyJET3vB2ZjYhA4LU2ULOfoy+hwzXGinqVsFA1WH6Y49R9dm
QS6ZVNJveRBwRxO4imstbHTwYKWixzMNCGb72Xh3GPVEihZddgLnfWi55WlmFb9b
1FxBWBTh28QH0TGPDAGVDKJzF9N2i5mHLFKr6JwZB91KcTi8QyRCHOKVDKwJEtCV
Upz1pMZhjkAK04NO11D8PBRq1xVDkq4k51iXgKvHD1Z21AUX2b3p65h7Z5AUnKIZ
sEjH01BGYiLweSqZsuNIUPc0SZsUVAlxylvo0cTZbW+SOO/JYD+7oEcgsPk4SKoA
7XS5XQEr4rY3N0W37IHgKR8C6XwSSooHAIAlSjHxwIXOY1EsknAnyAUaxhuqKrBH
L15qguiS82EO7ugQuKh2lzAShe4VJbf/MamdLEitDNeIgpFW7UXFKHOge1+/p33O
0bYhoos5V72yynRCm1yTSGZaXhTy9XCdrgkmYpIrj28yaTaSKXRzlru9AmYjfoD9
5estrPxs26AEVukqiubqOi+VjAHWPAYue9bmuE+BNImiXjM/nFpjEBRPCslV64eD
f+8weDN0s8uUHNFDDVLCxv1lAOYSjRcgRRA6gXqcs9zDIUf2NLbHQLyJ++kRJuOs
n6/DGFxyroAaPHcWv55benx1WWKdHzy+3cLndgWgchumNojsqq39oC+PK3mk5nGr
OezSjuuvxC1EK4aF5xnP6WX9mJGBfnOdG/bijjZfSpVFdho7+MSDrXjppiPrUrQc
ib5iJAXZJyNtw3TlqKkgF/klmj+WTX0joX3Odmcax7U4F2WDR8lt6lMl+M7gXPU6
uCViUClzHaO6dxlAMTh8CjidSR6QW92Dx8JZJIsMJA5mRoQJtgIHrwqSzqytMU+u
oXCqjvwav46W5fZpGj54GXa7hd+YnL+u6eCIqTFRVGdmDPopxGO5BClrfLEY8GVs
oG3+9172p1vvA8UmCeFXcaMu5NJK/oix1fEjDAggwy9XfeJ2b8WfaV+y4iho6qdi
o5u9snkQ3vkh3dsjw7mHRrizbZYb55Tsk9kod35HPjwXUlIgPOdqULpuUyHhEB//
wp9Hp4kYJRlKw37G9Ep//uhqLtX91k90wrl8KeUVR/Sjr/iyG6Pcv2EBXk9YgZs6
GyZ0OlQvpBcnLBIbx+ehMJ/d32bhv4Ud1ZI9NULePX5Nc7XywwR/v7bpRCXt072u
6omj2zoE8zomKmlK4DlXMYDAjAS0T6M/zy7BMLgW/xtjv9IpU7WugIaIs9Dvyli+
3Gnu065JRmvkF1hp8ekyVU/u4WHSPhuKIEq/DjUKmNtr4VeghxkVvQw0v6Nyzu/S
zNwK/r5WTHtpSBfCr/7OtVHixSez+A9hSUh7bmIH3WY3qCTbzvIYdNuQ3vM8fBXU
EVZyiq4WBilhqB+5K2BQAGvsmqTfsIGoO1RGntawLtVVN9j5wlJkSQ04hggk7hyz
gZAJ/cbzj4WLaMCGrSnsr/VAZ/XkybMg5U0D8T4wRsoFjtxhOAqBWE+WOfIXRStq
lI6kcghOA5ne/Zg+pUCO0UCZxnizfCW563xdZtWH9RlPNOhaiEvEyy4OCcIzTXiJ
bchvXglhIFNa5rFAHH8pJrVwLKrtUPCDL2QkSCI8TcARvGLCH8jbNnSMK/iC7NOB
tNGd8JusDqQLlif2aC3N9OWU13HoOW0WHsMDWIfkokZpkPn9XZ5jgSOcjfAdUgKU
f9Tim1aU1WZQvCVaTZIn7qvj17ZTnBX+9TsD6p2Pap9KkXhIgq6W95DRQ9ebpEHs
WfbrqoFXojoCpLroOz0ZYETumRC9XOtRpJl9lzmiWM7L4wJ/iZeVuJ/6H+raxnvC
s1Ia+olAnpZoPY808gbE8l/ol2LnsTpt1iUw0obGx10TsxbcocsdjH6eTZeCUbXx
w91WDnqBKiMwU2afPlpHZJTQMPABIe+hkHv0BFC0/Va9XO/hlQO7hXomnclpI3Vm
8HXtEAxTsZoiPbPNjk9FuxHcHyUAb+/gcC8DFOjMTWYzd0V//zj8T1pDpGpcfwUL
aVJwabZUnCUlw/FuYLe7Xp5bY2KxcE3tOQSJ9U83R2WehkarOR6TNk05jKkXTRuB
teAu7YqVG6FosEiXdw0CpJDSMvDNCKjuB3sOPPoCzEBaaYxAyjDbgidetItOVKrY
5n8eqq9h39c0aZJ003YDXzDM64ZcHSoaF+9FW9uNsCQRv0qTw+Xa0IFy2YyiBX4p
uKoM+PPdwhfaoSJWhj9teBHz+EvPH/Gf+IU6ofg6Y3LpOt2LRoJXnx/O6ZqobIAQ
gLfttpkc2RzDUZr/uEMzd9xhPWtrUCeDuM8xIsOkojnOFodXg/1FyYt/9uU/TZul
OuvdQMwBlT/nlFdQDM2G8I+/U64BqQtESbSQUjVOgf3eJrLJxfB3whHBbNSFHX6/
BphGJVnMlwbkZVKLTtyCgoRvIYddTvrCXD53+U3bDhx5HAIUvRVytuQ9z1OxROod
WUj0DdUBBAZRSn7elcWTyjlQWv6eMIVO+uN/y0gYl2b/+mhGEdpMLOuA0xbtnRhL
95GoFKOs/AXLTHDZmOlJEt0udhKQDlnU4bz2YJHTa+bLa9HzXFNyoig2vMA/85iO
oGwOpG5SufwWHh7wpQQOvc5Prz9Z8IavB4/wnAP4/XNuQp6UB3mra3nCS94MVquO
tO2nTLoyU4OpRHblvly4Yw1qjb8jmsgtuUfFnDJAf/o7O6DGQhBA02evnaDLPdyq
/5WfC39zdQV1Xjj37IRGzpifqWWcyeifR4TWn+QgH2lyLZeh4j4KcsLhV8iibvV3
UuzeiRWSgBvDvNq9q+gfBKlkk6CRqwfJq3r4QbfUux8RgmVGIkogAhCFI52etJ80
+qUUdc+9G7qa/PRkV5PpzsBDH+O32zIzPmNdfcLgNVBg8IMuaCOtqeuK/m50umlR
kNXW1vUnwR3HtOiXF5oSmSH/JxKLanmvfry4uIbzChJjYPKyYr5t3Fw0h7ndJLFA
DWjPrwAVKXZ6NkGPI5dHRkHqyEGWBoYnrnNWafd84uFuhTuGsit5ldDmZlayU5Ta
vHOosArW71UxPPPa4w4EbVUPJmOHTOmWE3KCz8RGC0vKALcqvM6LUxhPvQzSMhCk
mT3JOBLkCiLk66Skm2L/kkMGLB8V0nYWFFyNRMSdF4RzQOMmNs35vzIVDo+TlaaX
VI948JZTy6erpnxgSK8jfa2pOvi8zTaCmY8KuBBsa8aKaHvKeDw0GcMtrKtJnB7a
yxHH+zRD5N74QMxZSvMVmEGibxHomGsNqelGKumggm7SaAfZed9TTol1VjdUtmb6
0E5SHNPe3FrKeOeE+N9uUZkI7UTCojrCHiB3ASVXPlIHAOcjJDsi1P8C0zGC3aQS
lFC6nAXcflOYrLf830qISaM8WohymjPcZ1ruIq1H+PjJcQhjXZLs4rVlDpdXxNTO
MCA0dm57eDKxYo8dXUNQZrYTeyWUDxVM89opyq5NxljqNBZH4dqGvEgCTIKae/r5
XpJWVOaQoRKTnubHYkyUfsG/4jqZbsMroIZdSTHmqJAg5EUEP8o+B6jHcIZRfp28
H97zt7lUJckgu/RifEaH1QRXb6peeHELo+Ph9PYUTbXQ5kLwdkPLxeYM97bHrRCj
RUIaFzy1GLTRkKZRw+MHPAT+LEGvqJKEXcSp1U9YkdgUUQ7GkuToFYCUSh68rDMi
L3ojOxD4FM66QRXETaxpGyj8WrlQ4ZR1aKMBf7RlVGC/WubSOHKx2gR41K0wRBJP
XjTYj2OnMIlYJajW7pdkME+S4ioLpHOMMq1OTAm8/+sTf+Al2KfYtEaIHnsCf1H5
TFH68GClSiBsJWcV9xXTttx3Ygjdy7CsJqTkd/AM9aeCwdXDekd1aYTw7XCApB0h
kghUUl3nPV2+L/9x/5QY/iQEP1ohfm9q9F3C171V8+A2PGgfm0Kk3exVVub4iFRu
AuwieUCvuRFs1e2g3j8PYqYE5cEwZi90bhE/q3+vrZ6h6y57oryE8JMPQlCk/7vX
WlfS6YHA5IHqsoX40PVI2QYH2xLp7YP9zEPPaB14SGDu46ovQhaD7RPDzf/9jsDR
355OBVji7FuMOWJ429WlYGAtUg61cQJcF50EFOiJLA+nVmAKYNPSOw8rakpo5Dx9
frbQHD8US24jU06H1NsTPDcxZ6j1ocg5wtHuxX0F7yRrq8iRAn9Nwf0gg2Wy0zE+
d2r74L09glhU/xCjV+RTPCTuK0n8gO8CKgeemfCwjQVDCPiCM4lCnlCeZi7lmwsq
tKW488o/HNtzlbVnE6ZSAHls1gFzZwWSb2BYOOhEPd7P+d82+dZkDys0WwpO2gew
t+IxLKXPTULpmpM9FMtcgUQ1FD41fqIGp6R4+12Db/8FHZNhVWkVu1rilARgVg7Q
YTUVQ9DwqCijwuF7PdhVmYhK6+z1pOW0OBTLkyDdXdTFDZr46B2D312te6Q+6lwr
ko2yZ0RCJfBbCSO55RVuu5d+7EUUlpREoq6BkUbv0gztKWOxfmYlNir3ryS6gnVt
DEekQG+lyT2HrqkadZfJr4OA2t8ZKHtM6NDdxyDEBSbTSluYOe6LUyIcFhtzhCgT
ZV0NUctEAcSpjwMpIXqzlX3KpZvCy4eXISpoAr9iIPKMIBVADm4wpcEsppayBal5
CxqLoLuO7hJI1ANEW1AlrdWTSFf0qeQVGwmC9hw+XVBGUs6yLEjrpcm2Qo3Q5GAs
q5sq0glYhRDhSnyz1ALmth5Oo2hDzwEymXkAx0iLX2A8pGtCzWR3D8QZhTBnALM7
06EbNjy4+IBb77OQKj/IyDBuH2MtpBTkTxJXc+J6xDNUnUK4Wnzc98yh9q7HC3Yf
p+Pbl8rF6ECAOwYtwrBqPal+vei3c7DN+IFimhbBVKVWhpcxF8+slWcy7MCDGPPD
SBiSuJ39BgJEu+lcJdXJqZ1JAu1dpM/2oXFlI0O1XTvvs11HWWU8wueVBgpEpTzL
GSZ0X23QdxQap1VzjauZde20Y4x6tm2mgEIDRm4cqKZTUt7Cn+ml5piFA6atqlmB
edy6IC0rxFTG2aLh1kgJCcFDSn0FtC5Y/F1DW9J9u51Y+mUcgmVNcAZ/aVL7BEs+
XoRul8ptwFU733VDlUEfZNextB1khvAd930/kyOq23sUJ7MGSI6Hrszfp7dE21Ns
aoJuPbDnTairhtBAAv4W9hsqzNFVUy7K8bKC6/4glKKWWxR/WgAfBNWMlUaYEteQ
AOuXTgGVxqw+UVfpxEsSPRcaF3BHb+hR/2Fn4bfHELtSqgfzLqpROytkCBukni3A
FySap+ZDYoXUQ1eQjxgSk/wkIFGSufusdy1srxyiGXWvzH4X1lrCBSoKteTIhuQk
+Gxz/e18d/t3F2EqYcwubUsyL2Ua3qhNf6zulEUjmJz7PLICmk5hLyJ3gfWNdna6
B0aiHPsjceV/eUc4xrvEr4bTeK8EYRHcgFx+WyUsIfvOgoQttaBPnuFQXsDmjP+I
u4fcvVPUz1w/01LYicIca9V/Qz4wIuhFbplPBGwtkq3sqtEc3FzgbVq6JusQnZkW
Ivty2+7sHRdZCIJVFpPEqyOMynU6uFaU0vvZepNiHBtgLVvK4uCMk2dYNbmG13ld
2LWvyI4e7FeBFzNaN3ZfEdJnoQwgOQlmGM1bDZ8Sp3w2al1DD7BytgyV9GASVMcl
ruwUg/r9DUKVbj+LpfIEflAt8Gu79HjWPA4ObaUetDailFm9kkDH0OSyuPz97lkU
Xwh/koc+6L6Od70uDLaNBGX1JsHz5NzyknalP2Z9e4/Uq6uq6U5gF6mTxDYza2j8
cVBhc8gHP0M17gU12uC+CIw7SQwoec8rH0CWKNPU6XzgOBKhFQXWaYwKvu0TVC0e
IVI1SmtGwp+/tzmdSyVpszul2kFQ8NY6vm8BLBZqWv5etNjUjd/Vnk1EfjoufY6i
x+SmWj97tEH6xJkHaw99e0OcTMPtJ6pbjuqCB4LZMtpOEq8bJxAKd4Se/p8TXz7W
4y7C/AW2xrvoY2aNnDlMb5slI7wxkJn8e0SgcaOzCFQilOJB7cr1jMvuXv3WIkaI
AyAIDiHQZVUIwyLEVS7NVf0+ML1Iamw8ISNwEXlowYAXtlcfBCkWVjxiCnxj2O6c
B+2KMuhQb11i2euDTdg7PFJItOWiPVNuTIVkLi22lVHXzOOzfBoX/l7X1jmyPLOv
c+yWEXotgyVwokXGmtTEO+SE9ePk86ZubuERBYtoCpISmIIWjOWB/CpINU+lDxH/
jLTxAJ0nnq97R9hujnBYx+glzvME8AjrPLPqwUF3heshSMHTkEi1evkmjYdP+Fae
jIbB9dTxK4jm6mfuCj0O8JA3bcX3OwjJ68dLsXpwCLGEyGBrV8Tgn4ib1oFsZMbP
Gwvs0Lbe0DRPcl59TYYTOX6C5kJMZxWjLbVfhhev4bqszfuGsTllT1AysGGni2xV
xI0MRSFaoJIOGnXuhjPFFQlMTSz+14LKLOme00MBFu8ePmCeLA689qbftf3Xf9PK
m6wUbfp5YA2CB8OtmdPCwnSKFMvOmVYXz6gbVR3+nXjfnslw9PICk4yq0FyVvvj3
7lDjcW119WN9exMoo8nO1XhOgyd+S5NFkSOF+MxnyWnOWs/ZfCjh8+plK2TW8ytR
/1LBeFi1q77cV6X7E60p3ghU7dZAssxn8Tdeg4YtDYI3b8KUkxeNKAhfw0VLc+Pu
8oidr9+15ifpxDoSyQaD5e9y+t0bckVovsttMkpfjwdiJNcZVg2Mnm+9+NkDRKaK
meUFnK6140bK5O3vifL8sU5GIBdgpTaffIdmpLQVMuOC09fzprhu3SaJxfOnxFZS
GTijNPEOSLNpOjwgHzmL54/AVw5X0QHSiQ6n8HLhGm53f7u3PSpm14DICZWDTe0+
AFJ9Js8LXoCMEjwjKGsxUMnbhsSx0GvwA7iQ+/qvDkAKTLz/3eBNB14rHMN7byRM
Wx1Nu7H+Uwul+8ak3d4bVedgKnfHaWXie0csAUVY0oFthvyQzUTZuAPEGRjjb7+9
92MByXTGZgpbmErd+IudLrE+4EkqevLn33uV1tO+lAXJroUqBzIUxnMdcC/uwumL
qkK0OUyXbJWhSUm+TsPtXjk8MMsOwe/lesJ7SJHoTV4eDWAFJTuEqpwlItFLnWYU
ddGyBNWM/2XcDSQ28FzH307dR8Xr0bpLIHv1fZx9aVATNP/HtVtITVsd3q2jEYfO
FfEdTxiFwLv21TDfGe7Cbubz1P8dJv2RAC0BdhUz13KVlT7/HIJ6nBshA6GMOqR+
QbvwsXm52VD7cxMwCtREKsakxyxvbYtWrXkDrCpf3dHm3zYnkcU4/32xmjWyivll
SV8YQcn/+8aM5oOEf0CJPjwa+Lnta24O5a3Iyx/+qyst2hHM5BeLWCwZlnkz1Pvk
bs/HgWXeUvTmgJxMlQ5tBff/4oYXuhQ9+ZGK5WTeOpt7iC1hyLAY55is60IFHidX
EUx6ViS6dp/51noZiBud/K7tCKQs7XmYs7Ok42nGhJ/khSfWinHIe8YE+pdzQNsi
YFsZkbYxoiaKO7hoHtOAbLra19nk8VkVH/d4pCxJuIc0ngkkNhr+DKrpMq+Z0Cux
qDbppPOo9Si28AZU49UWAy3tAredcaHZXHNidDvliM4AHdr9mPC+Ag++cinXaHhf
EWNFWUGHoOix9QI4XJwqT0lhcLSlqcDIi+ybDj44eYgI7EvQcjVm0drTKDxWm76l
HLJiWvZQpiP1/7PdfS523iz/zcgQ7tSFXGXK6MEQYpGS4QqUfaCEeQ57omnjVqmK
0oCOph0z7tnvC4Jho+c3T/pKr0Xdc9GeCxd28hcRedR0rihNGat+G40//rTWNsnB
osTavZwXmWk2PJTty5GDZB+taVsKzSufTMLNbpeLoX9RqxqQ7+adQp6yQ1sr596p
xJ1yq5Pv52tqpw5FWBJAkt708jGlkWDLgm+vr6vFb/ULM0/r+ts/J7s24NIWGXty
vwZ0mqfMY5UqDRu0xEHJ80Pyi28oQHBMfN0xSgiPY5/NZZdTn+5mw0TZBL0s9kNz
ujsC234iW4sCUr2t1DBc9Md3g25hFrVCqozWgn+JBkRq1CQl24+d4XctINJBBAgY
7jR3/0EhIARouA+U+RE41Z2dSx5r0te9aHqc2oEyDl4Wo7XZgEL99r5pUjwbgX/m
QYLAtCXGeHTJrex97GFRzf34H5GYVYbqipWYY+QFBkLeMDSjbsVjTz7FUgZIRW1n
9oC/LIYJKFL+EixbH1wjmmxeY2A804zI0uN/gvY5WscVbw0Tx7hpWB4QfGvO1Zz7
fMNX0xusuQBdx4Sc1spc0+qI2TdrwfNv1b/6ktamJ5NxTSge1HQNhMaFhrUnzi8J
MT1Glr9zaq/r/IhrKLmckyXLDRvWbwF1T+7MB3zjtGWt3Xf6EGLD5Xis2qUovPK6
t/bDpKUDfer6hSCG5IcpIRXiPyFfAKJGVqdnxMXpYQxV/ZHqtVo73AG8l50Kj9V4
7u31wakmVOKB3EiXa/+27nNRuqHZ4PGxfqMaGTdOnBCZ9tNiwtfFIIU8RMc5tJj2
UyKigFiP2B1R4Sxlr4kpJkC1fl9RlHaclsWhYhATZg9GTnAMVi+Y2Xnq3G1erQA0
yRnshZUkEmJX0aE1cdXzPVSAl4QXXu2fOtNK8+sCA2cnbkTROMOeBlE47GcbwDxs
gZnSY4dFWPPrZH4hETvcZpXmoj/7jYWWhRJVP7dAA+V75LEMT5sn5HNP/yauNzbn
enKj8pVfYARTxL1H6ZRCNZz83hZkhh4Ymb27dQbLJVCu2gsvJ+t0LCrGrlddaXFu
6+rjXNem2aTyMTm81uT9snQJ0ZiuO89E9pDWr+ILz7xZyk7cJ3VIg/SnKiF9Qz5K
0992lRg5MDlvOBQcivFmfZyOHE1o+GY8ODb6cSlvnRvIvyujLoi1N8ddVa+qx9Hc
YSsyKLyAlXMrQ1zj4WA8A5E/gLzBeXhAVO4FG7eLTgBF+K6XuLErCe/frDhrDTDL
bYsvt+8TyZnyrgGN7oLMndH7nePs06Z5UL8yZyDNRGK6vNypDJKDnHdw5enjAOgi
0j5DnVkWDuxsk1+7mgB3tgOa2t74yVrWSnuiFIo3XR5XllQ255izzWRADpIpJY0w
yicLDFP2Ve6GTu2LHRppr47eQwMcc0Qt2FT37afB6Du0LZJ964dOZF35Y8SOxMG9
Jgvz8Jo7nhX34hso3V1itA6u6+hvlL4fprkWeSXrLQO5J975IQZcNj5fzNJlGvf4
5NaJwxX4ZWtmCG+zL5qduKstS0LVH4RcvMNNutDPjfdOHidynTgO7SkL6xHQG903
0UzOY1AaNha4fj2iuvyUXWi0YArxl3OoQYzH9hWcfuY8YOM8yVDQFS4qAveYoYGS
NltBNgUJuKD//7ZY2kkAmX10Q6piZpKWngl8o6tkuIeuIHC/wCvrauKnWDQL61S+
KQKefISO1Hpewqfanfl7qJomSIuvmib8v3nduI8AU4gmuadVTPWizUPCti3x4G0e
Im7Bx+so2TJacIpfU4PhIb3xGZgddsw8lagfGDLFXdz0Qo24Yi1m7axKIBPQ3Q8D
MxuR5MOqeYaHvgeCYaQ7I/knXjRqXwWmzHXGqrRJzs1qTi07qVnqGZOqxIJSCWXP
MwniHIIr2N0vOmv9U0lvP/5XfBSkYks01A+ehuc1UgQ0DxdZHNkUcXmtO9hYfuPp
Pggs1WF9eAMz8JZB5uG05jqiQKiGWBQW+TQ5cAjyTEBN0R+eUS6eHf39hw8hBxVq
kWE3LbXwRbWfej+KGvLVAwnVzAWLPesZpGeYJHcL0AbFirh+X49T6cv62dMNrVSq
iAhjtN68L/tHK9vpuKtW/83G5nbSp7b99XQbI3tGmrC914TiTAl1WV2e0Mz04jFu
SKInH8Jb3tyVtpmzbY1N21m/vSdapfKQPCCWN8+NTSAWFhOtGCWlx/S97XGk6Rr/
kywsfvyoQ9ZywT4p0q1v/p9tzmAGlMr5z49uxyiqwVr1q8LOrurKP92rMlaQTz2q
bmNpNbAKXBHuC/n4ToQrQortZwK1rYnYhuzORD2EjVZ8uWQA8qRjJiPaKQ20D7EZ
ojHOI061gAaeRFy4ivuIAncEkGmxNqS+/y3T6JL5vd5g9eXnSJZkMOQ/NUjDU5aC
24O9lrTaKy7/NyaYyTAUtjNrC924dWsfcH0B25Ms5rZxvRVJJJRuEHEfFxUni77q
BkiVqdKhbXwLs23cNS+lzPUNMpq3ithHGX9ERHyXvpVMrPIuc5JJT2MDBn9Aeciv
4gIj7Xk9na0Eg8FDyRsXzJIIh5rg17m5iZrTrHyBUzx92YgQHlx+56w9AazIhmnw
PZ3LNfAO1rBoGeFzls84SjYhIy819rAlGwsDY2SARYHYwr4Lkfyhuoxh3WTdpW7g
Gjmes0P60kMAzTYT17UzoptgifO7rzEZxbPuDEdvcZ0qkRzmtzHSgVF9VtPTAUzn
65UFhdkhZHd9h/g/MA1sVKVBD5R8W3az7XR8HAttHQaGkelvGpHAC5C7agriLlRR
8I1iYJW9ghae2gG7WtfbVHZ+Fnblci9G80G/YTWYD/+EoauvxlW4NEzDqHumEkOJ
eskd0TZIj8g5/ShSFoPbBpf9frgwXA4qYwuByx2Dp3WHFRq4wmj18k7tLqSohLyP
cq4J1qIwM5w4i/efzBitpEiXzy+yCeKD86YRIRNcgkgNpwvamWu2ARJtiGLWr8QF
eCEPB5qt2i8ZVJ2ciQbYtNq3CZK8GGk2ZRVg0RhWjYZa+qOoH1XeBVRv5fDYgKE8
EZFJtGpWcNIal1f/64zAbQudEIxH5OEPktdmQxL6cyg+0j3rafE2PFkVHBidEn56
Gb85uZCFXxRNnth6cyO/w3eAvZ750nBh/v3aAFxGjJHCHoQiKVqUZUpgf90iKbMO
mRQfE2YeF+NkyKN9zsOylR/GTqu3Nt6dTGcyT1GlRSSA098sYXhpkc6y3glOX0TA
ZUE2so4dZFBL+GWgJJKOB6NuSrqIPk3m9aEQt0u1gFzKv/w1GIxTdBc9uYkDMSA4
SvkWoYv4ZSby5A50lXRbIhY3UZx2w67yqLchVdXqEoViZq2pDp+S7wjSihKlmg3X
wtCbH4aAy0vZCIzax/ht2vmqMRBJN9En2U13YIbAZgWAAI4VRY3LRwtdw7YM5LKX
VvEyOzRvMcJvdNpfTfuZBI4ImT6aI2l5kHjf2+YJrkz+uOvnLa/gkop+gvk+BRGY
qeplU5ZfmcTGJ9+QTIk6itDr7+uBN1hmq0dBA4Bo+za1nUMdZwspPohSH2+kNjIj
cCIZW3VcfYb3E6G/qH+XYfZFL65gmObjeJe799W9uNyWv0DgQ6vrxrOpwCKInf5s
jcqBIFe7cfzzshO7En0qM6O+MzPgPNgZWRq1RxnVivxh0r1YkqtKOSWc3icIbCHn
goCTj1LFhQw59FawOYbWQ9JnOXA9jfwFifzZENyMdSBkzbO3YZm6qWxELmcMyA1K
gdXVCqcEh49LQD/pmpUp/HLrqgI8Zx4IBqgyR2VsR3UnYB0/APjtDglbu7YkOkgb
3fh8uhogliyFUDUMbpnkvQYcYBEvl+R27dPyiXEfsHf+mmf6UHL8RMLBJHEM2L4V
a0+V+AlN/ncbYUlmKnIroRJnzf/LED/3pSx0dy6buCyubzWN6+j1Xj3lORNeWk3d
RRJt6ZyR9vrPaYNQAtHDX878GYjErOv56sEPOL6d/enZ8R+ykR247zs4pPfk4AJl
RYWOG2cmx6lOtntyNvDd6Vs6ZWobGmaJTScH2jRqksCVcpWt3Gv/lpiiDTkJmPuk
zpxHlVd3mTxBl70qI7JUK8E2ROcnilj1XcJYkzTXvPt8ssYVOfdqCYjnlb2zvxRT
ID71MR4o0ZGHiP7uKr9kPHH8peHvfIVrjSDRX0FsF7tuTdUzl3pxUy1WUJImO8gV
8uHhklEddrmJxdK2RnI3UIeZYBNxXjDZg5nmo0MqD/RP/yjDPHp7p9KeyKlAvstK
tibEsuRawHO1HNSzEI+HGpcBtz1J6PXXLlnvAst4xdXCM/jN7C62eJhUzJj/tpO4
Y0tHPj5ODj7htiRzMZOkGjnTDu4Yim2PO47Y6Vj4Zh6AddKXAUvQULlDLJEnsTJc
COmUKYgsT+Oq9X09rbjumb6F2x58v7tGDteA8Duq4jLIB2oWqDWXFzqykDRhEeXF
2oLEcsJEukGiqkfbOOquusNIAVPGb8sdzqero/IhnGqCBUoZ7lirNCMcz7bzONcy
VzX3fSz8d2uBT5UYLRbFOlKlCR0gRaBrkgQdAfDUdXHmwlIrrL2gvqNOzIT/Cm1q
hYYheWVgbZ2qBxggN70d85YbCCbCtA4OBpvU8eRzCT2mkG+n23KoTIM7Yf1ehN9p
1CwQ99yXIAQC70JSIsciXHYdQxW5on//T2it1yVps5U4oZwK3OW96Mzw2ucxTkYN
DcI284slwaskW+kkdHF1GKPKP8NYbJ0wmNiWV4eFZ4YJW7cGjqrFTZya3s+L07yg
HScMQ0BX71En021y7saNHF+gUKZYhCh0nI1hy/5l6HBLe9vCa2erN6/VOXopxHa1
i8OsCvnky3d2nRyomJnZyr9XH4bw8E3Yxz/Bk1Adxt1Li37Q/BEUBCCAOwRkeFVd
I5cCtzBj45JOxaWOIw70J6CuTPofxnSQaz3X/cg9+80wcFf8xN9fKAyLtl0vTTKn
pWwROgX0+fmwuVNogcSII3sjKUh4BZsAi02xoLjDz+sSwZqHlaiSttqoy4Ea3pkG
vGwcfgof9q2Ejz8e1oKGy+UFXpF384G+lVlQK3HQTfkOKjDudwqnsbx0I9zJTt68
/cXDzcRrgM/airIjvPnWHnt4lk4bglvxOX3feS2qjMh2luiFkgZw3kzJ3tWrP6S7
q9jzuXNSe/0quJ9D5XHPYaP+mOWhCD2ZwmRwXSL2FTN529cd+o1e/gMuUmVKI/5T
mTrJzEG++gWLAjmhJyW9YdlIh5E+yqA6UzwvT04Qco1ESSRBlRIVBTcTd3SNDZra
DPQE8P62b4gdW4jaiS4odVn1Zp+yEq4VKE0HPh+khd8GrDeylBZulqQ1iWQkB2yz
2HLTS99uhhAW7na43bbSAFN82CA6iWV3xajLJAA7thyIg/F6vbiMv7wxVGcZP7zC
y620PrOk3SwX9dB4BoaSdHbGOt88ngPpywPrW61Mn8uTX8cwYrI0vGiVEIfzO9Pb
6L2aEO/NYNABSvpeScp++fJbTfjbSDtoqendMV3AU2nPACa240WmK3DUzRhj6NNH
yQMdubkVfsxoDetPBH8EsDtV+HHCMG2ID/vIrkFpQFVqR3kc8O43snXwBW37gapW
UXhEPKJpdXT++dIC6RRU9oGfPkfa2u+GyJM9Yi/8LZIxjv7bniylb4YkkXiqwg5q
AjYEnHA2K+peOxcO1lMJl5D2AuyId9ObubHcOCobbzssmpYnhNVexE4Rj6JESU9z
64rdjqOueF2+Xo0ITpKo3FvnuLBmNVhea4hDCOD/J6kjFYf3DTMwn3H17sHxpgQ8
nis1Ya+HJJcH+c61JFgAnWKPHRUbHVqDYduAAt7JOCzsc3IsZeb+3nbs0fQm5f8F
4UNCjwAonjJMRWLcUk7LWdqZt6S4BW0M/Vqxh+r4lBQzTaZCUvROs3nkW4r6hU+R
LwVj68Wz/Zr6YcPS2rTR4a/fEOJRnTvsYr+O6QLZF0hh/KdvJ7LLSeYFUH1Hg7pL
QRfwqk1xUXxVreAFXSi+OWSkWQqHSwskLPBaYHVDxm6+CoY1HeibGvIRZgQPuWCZ
8rPZxVQy+xq2lWv9HMoZPXMT++hXX99g4UmINxyddgzlg1ZvSapWT4gqrdSpFJoe
fKeV2Md/4kwqX92bDKqhLzxq1gofMRVNCv+D8H8ZpL2+TGmHqPPRKK9fRaQRK+w+
OeQLfl8yUSuSYuwE8I/KZPY2IuqjqA8kYsaoGd+hfl4wq4rOyDJtdE51xZ9WPYTf
YdVtD4sHU/cjhKBJENRmkKsW3d1i1ZuxTL1Cz44PjRpfIdYJOlwt9IppzOUvWS7T
3k5ro2KQUr6vigteW9L6DI2HjWpr6getmSI6RdTID4qvC4DL/PgzkdnaCqiSN0Hp
OZdWUdVC7a+t+u2HJBI5GwfMV0Nmk7DfnNkZJb40hbRFrOlzGNaKN6i/kJCzNaEx
D8zXaW4/sdOov+bGmG2J0TVFqmFTspotErsbeObzIgnhlxQ83lMbBW0damlhremo
Nv4cR5dBWOAg7jrsaeVs0nqNn9xSkd88RSc1SbZrPquRHyriTBno46xZ/B+94igJ
DdRVZJLDvufSi3f7q20/Wn6TsJpTuwdtpLI2IDrzOJI0tdtXk3aARZgsczEccL+q
JPY7SBL0lb5T2+67KEFL4ccbna/W3VkPIxFQpshTtv6FoKaM9ADC9wsY4bkhXuqi
pLtTgnnnxghvKfa6y6We+voKKoWBeq0bKRT0QoRGD9GdVVz25jvuqdEdYeuBuGvo
abxrMFLGXLcnPxkLtG/RReJxdZGTM9QCCOVYDHO5AfYn3ww+dBm0SNBR4ITHGI37
LTxGTg6NQP8weBKkAJuWDTpBwXLY8epqwy2HwoPV5f2rpV5XSTSyOte4mZnYZYZ6
4GJaIVoQRsq4ORVBwCtYCikUj79KRQlUUreNbPgwxk2to9xM6M2c7UYelpvLdA3O
/VrBSdiTFZCj73wef7DJLGwKD8uJHh8q0u6LDf6Is8qkQ/m46nkDnPA4Nd1Z2I3w
qvjfUWpcB2vxWOFJhUdMra/z2ldFNmRCFk5lk6Po/Qq/zSH/SHSbaCK4AgA5oYaX
ti4xHsq5Biw0ODXBy4HlZhK5/bIt3FVdEDw6ZGNfnQuCvRzkvlCBCLD9QtKDWf6w
epo6AgIBgvpPRgIz4lZdWeWf9Lu5Ft5UcXqWSQvq7JvmW7gWyXKKIcSer+HyA7KD
eWr+EtRr0xnpVjnrynEkULf4DfCqeuWIiBiLXKJt1Xhxm3jq2aR1fZjHU4uqFlfT
wklOxz3XC6FXBq16vsrhyakmZLIZhGAlDTpgHq8zKQMHd+ySHkaQdk0g4QLTdkiG
Egzk+ovd9QxyoDUtrydgt4RT8XD+pvEoiLkpna7vgOnXI55EwjpfBhMXAcW9ZlDP
t7qcTZ/LgQYWj0k9dL8imJZ8d1UlouUHNOpAgjUj9RP0KMDWtEs3WMVs9rF+AmEL
nxiFBpzW7e4q9hCGBUBzD5av6KLwMhV+LdgPxEYt1P4veulVqmDSdE/JQmRG3rs8
+zf5g6evdSfGkgNK9A8F5cui5KGlUBW25SyqxrSBgz8zFX+3XNKuj45LfKJKRe7i
ulZ81M6+sWblCMxAFFkgNjCmI0UcQkDe6+3vHJMxE1FPYINScIoTBHczd/vS4pRT
weauur9PDJrjkfaRgLwPyksYNWTY/ygnO2gxOQbjrPw04GDrNClcxy6O/cWP+25T
E+7fbkcVrlDCLoyLgOqTQyyRCNuG89BdZoUWW7GVIZGj+3vBk+dO3ZKJQS7IqafI
I9Td+FsRaJhE7fpr9KZ7Xn0t6q2uS5ZLEo4ByW48mcq4Wh/7qcFKU+M9WYFeNqCV
PWjSanbGk+GqXfBD86344tpk1+OJVjDgj4toTAsEHsgSs45UJNoP3nA0ZgNU4ezQ
FKiarsXfWUy9EEYvtvvwSD+Pu5++PFSvNE827PilMWkiuG02dk2nIWb4LDanK9Bt
wieYajPkVt5Zm4hD9w+XCyLU6WoVSzxpw4qBAOjopjYX4tEDAbzIo52HchxAzUM2
BhqZHKOZ19EtiJxKj72XzIrTlttaO8zyGPhpQClKCfyukxY1MhBbhObKYUPJvnS6
BYkB0AJ39HDGFG/8SCjMCIZ0WgXhCdKjUInM919ceeM/hYnUhW37S1ozeFSj7GtG
nRBTLR9DsaSZfmRMDl6QImnEU80UNvGETjgGJcVpLW/1EmABWmFVT1fH7ctE7dSJ
szhAHgmI2lWJjzl3et/0QKP6PcSIP9KVAvKJ3pagmpPgh21p9M/sIoWQfDDcgEov
LHMu1izss2lzAAgatIToUzeHR3RKmNkfn+mbaXWi+X5WvDdECYbZnZ73QkVQ2hBa
wIurPCcvqTcY2Fgxo3KUA95zlhwJMl1ulj7lPpOTl///09w1WuFiT7Dl4/1cSivO
DSji4XUaAbIkVnbzsAC7c/91FOHyitqlKQexqzitT/YLKNVuQjUaxW6NVWCmwP/f
gj/vWG4CN/1h+8OK38k6AvCgbpGx5bzylTvA5pgEJpFi19eyr7NA3OHGM/wbw7SO
BALWqwbjqlK/iXVISrh+9ssy5yVRY2HgmhTnoBxJXab+0B62N0oILE+bqgozlaj5
nOoyaZb4EOXaw7qDObTIuSAX3F9kg84ck/f9vGEFtuFQgWb7FfcN6KMuVXyXElc1
0/XFnAVjywOd0iT5UYFAlHX6j3b0Iv9ByYsQ+3oMscJp+7AVUm2hr22yqCabhKCt
xRJrUVvtDalGeIuImO5zCx+28+NgmXkLxqth/kwmhbU8uDojLjQpBE86tE4HtdKz
+mAb1bJbOZONmoliL1oMYnuYTil5RWpSc740ey29IuJugZFJZuQ6LHWfe8JQkgUj
HjjPkeZ+ScLCHn+S/ehDyAigi8xpdty53oYjynSpdc5fZjynPi4aHeNAVewNDHoB
T5KCU3wGL1KbdC+WdDXWt4I0CvwC5q3wDGhZrkMqLbMu1uBSpLbyrcaz7dznYUXr
/2nI3sli2AxSxb3dmqh2X2r3KoDBBuNjB97MfrgGpf3biXcV3pdODugEoLMuElFR
zytWDzw+a2kAXgCtZvzP4+wBnQ899Fr8LPi7WJvvokNSyF01whuRv3alyoL/YLbU
BJW6bzQmPCDsaYmgxA2/oLstNJR0RAkJ2nLZDBsdRKJZwfNE/ciWIXZOdKGIRklI
ljM8nmkGc5aw0Ybl/hfXCnJOK/LNSIA7vgJpX6y2u/LgNfGEJuBRepPbEV+2qNuf
bsYgJL11chJHeLQ5OH0TD+KHJU+l3JmIMg94cwvfpWrR+6533tgEHmmf3rk2J3T+
CYnq2wv5Ob1RQwr3EdjPPkwGuOQGHp7BtXp8zVlc0saMA+Q8gvt1sPdN8AH3I/bZ
SMUkVeAjeRmAPvd4V7lb+V/QHv7I+1eGg7hP+VbMzrCyO8JUE0A2A/A888nyya3F
civL0mXpEwdSP6CyF57q2uCTZjsn0gDnsdh+bwdPeXkRPMtsZGkf3l8HOc1IlkL3
YpJmtBTSysyupd24r7Br8IwhOqlT/kbcZZ7+LnQ/xekNQjafSijqHEcaoVQzHIqJ
We3Ap6SU1moQWlJSfjD/TLCcCmIkHFqUmBkTCFx4oD9g86HsW+01pYX0UNKa3eCW
TCUQVlgh76w6+qmQz1OHPAsmpkd5jydmmP6kEaOljW/gTtPikBkY1ToAIy8YyO/7
O/yFn+1js7P9vUhYWPNUq3mUcBLTBmR+ldgv2X8EjeKFO8ansme2Tbaw3Z9o0/Ns
9qZSNIJFWn3ayZveQlljzAzEYr1liXOwiK3SmVRMbgblwhASYipAZPfYS87XwVEM
O99vU7Z6Ijnw0sSkj03M6sS1N6fP8QoiHZ0Ow19j9sxVG5jFp9ZwnK3kK+e0qVlT
MXC2+zef18oYeoP3x6RnrwGkHpJeSlmeg9EWIVvwrmIYiPGXpLqLRnwHu/M9oLDn
H6hsRa/9IKcCHINMEsss3mH8FMfG4tlsZW+jzYoMBLTk0sPPpYzgmgjC210I7Umx
Ar7AwF+yJWz/SAoQGvXOCSApdUbncXaOjwW6K7z8hKH9RFciWrrkvyaF3V8sTZeE
R8eC/KbxTKqCr7O+R1t7QUs45XWVjjWiCAe3SXcgon0JDABibWj/sdYA2bUXh4+L
WmnbghK0OaqY57VRNzVDmQJ6oC+nHyDQj1uVP7G80qNq9LRLajkfXCC44tMQz5aw
o/JRRACyVuDnGY7p2lV4gufuRRNSHiiEKIocBXKQxxN+XCjG2mRce3iEAS17GOf5
GRAVLemMjoqKmiTYq88wRDybLvsQBAAExBHGMc9tvdBWsncxTOR4L4jUVf+XjTxg
RSQFC4UQ0pqseMp12OOEFXNtMPBNJE9E4u7gVVMGiqZLZ08WBuLC8yofmF6issW3
bn6MjoWTi3N1DXFule3pn+CGZwYgjyFi9iNpQQAh0l+yMsXWD+j4E3B8w98GJIZP
BfCsPcXtUuQn48HRjvGo6/FVYCb5vG7ruYu93KIT60GDBlPZAkG7DQzr6juqBQiB
qw61t1nuxdT9375keudqkNNFAwLPOlwJnFVrXGgpakyRh2npj6LI2YiIvV6eO7a4
+8loA9tSqZ6Vy+9xRsAIH1/RrQvtzPkZxFlLnmM41Pfs0b9u5Z3eexjT49sriPpl
xjmh09TdRFPBXepTxUCZ88hY1v0WX02azEckNoVw16WO/RCcX3CZlLVGVqLDDfSO
Vu7sudfrHeuAMQbUQVFvCTSLVjR90GJ/x1enKypGriAl36MXFCPlKYiffFYKbXgP
Rs95I+FrLoWgyvs9zM8ZkTCpQ1Zzj3PvCQL1x3asCqbwSyifTOZZfRBQ2w5CdtOr
HOrFOGSFeCnENWeFg2hrBf+YlPTo2cZHFHz48WogFr8OTG0+m/8xrhoe9ojxlVJk
0CNN8cV7t5+xNzPiB/vsDDUm+S35/dyyr556u5T6Ec7B+q+7Y/0oMHOCHlAwsqVu
y7DEsYKr1OBhFHwxxAm2HRvwmH8QtIRwWabG3oeGky3gXsErfVCOyLwd1qT2ED6b
1Uo9ujxclUi8Qg+CsU6jda1GmYcmP0Btqmib4sCTTjGQVLFoa7ZGS7z8mhe/JJVp
ddOvLvJk6/yLadrt73hubN6V2l8abJuiSpjsuxrPdYZ0yQjQFbMR4XyCaCsryXuF
T1cER1ugrD26ivuCDa9/ijAapftMEQKFIALZPnX3drTRIb6QhCm85ZD+2GvKbOXs
+d4TlYE+wBZmBcQaBmAoc1w9NRoTFMmacvL8GuYH7BfuCylYCv7SyXEvY0pAdfAK
vVk9g8XX+h0HHD10aKW1rZALkl778KPr/qRQJUr/atrGb+KltM5AcSWwirM7NyTy
MsFgj9ZyrOrTccr9o4zFi6c82y41VHb/56J1vC5Ladv8h0mWnpNjTLiDQyJtolCV
fIXXv45fC+1drbqBSHVisA04/NZ65kP01hzkjVxSmxOEWt/4uYxSFP4j0Cdgem1w
i5+tHGCm0t7hQ3dpeFnBnZU3u2o66y9pakN0zb9E33QfWggYRyusdLPXxQ4khVFx
FmW6X/+nQF0oakTgv48TCuJczNygZMdq2PVeCvZRCZD6tnNxf6qBk6mMJfjvvZIX
x3DeJ7IG3UZoDqERQME843BRETeMh003YIs57PAnyC8t5B/03UipdsURzTvAXBHf
Prd8SnLaxlYoMAWxo9w3P8ZlKomawwF2g3cDeh1QB4JMbDVKwodRcyAhFl/8Z/Gs
viB3MW1zi2HYE5txULBiHvDyQxYdLEOsLrILiQm4SA/RYMLhJp+CKUEznW8gLcuI
Ehfsjn++h2466nEnsfq8dOQ7S9mpACqybDVj3iDfsi5fEAsRcq1tHxd5th9wgCdb
sdJBSPkO80WSmq0+9zxkKn3Ce8E+7j07JzARKU4TyjuER4EmjbEKJd2GR4vmv4ci
I6U4XN+ZkpQMR8IpltUFD4yfthKWQV6trwt1R2Sggf78XKCVnKjCCc2rWCM3mM+D
bv26hv4vh5/7qmDJOOwYnNa06YvKT43Oh2LWVSPMxd76vc65vuUj+oa3r1KnkVdX
oRIih/p2GexGZmJZ34YB6fg4+H1PYWhafWlRHkv1YCSY31tnP2tq0UAVJxq3UlhY
WQQ0xojAxfuHAxuTPXNxIQrSsJYZW7Pagku/jHQI7R+nZAcBB/MWWLZ3UGMcVri7
3ZyG6nwilN4KPUG0iWSNLJ5gj4C8iObJEQmWQEvu2q3K6acMFdlLFLvO77rjdwlW
4yKVmvfPLFDs4ut3y9qa0AAd9OrdskVLne89awRj+udTzd9/BGa1Wqt6mjZS51/+
5PDXouPMePD0z0so8k4cDilKIMT6BLC7pISU5ldd7aDwQspk30t7TdV+fU5iBI4R
pvbuKDbE0/c9VbJNrbaa6o8CSRMxmXuOTk52AcOF7HGhxWdqidZKGBMQJORKoO6Q
7oI2DbmAjKTdNhuwwOpLedX02cKDNlfW9eUqWfnB6cmVmc/iYThikW7YxpENbXs+
Q06jUh3gSG+leyk1C/BL42N84ShCJHP9GaC3BEss5CKfO6tBz1DBO2U/cHwAU8Jo
TSigSugN4dpKlz9gBTonfpVAesqVg2cYdth2tphCmxxi9z5YTMsgommuzSZIMg00
hwsq45UdqeRPEPi490/WKrjHWGLFQfd55ya+l6jcmk2Urt2RMawiskI4OVdbcBsW
ifualOeEyhxDFihZtqEP822MNFLXyYcpNlqCSye/avGKCXl0NfnHcj0DLKU7uFAO
C3cQ1sGGg5czsKxqqt/pk1Ey64ZHEVKF+j429oM6z8+5lbB8F2kEVr6mG6Pv/y8P
Fi/Jrbm8nWqD530FltlDFMANUtGSHcSZYt1cgnJE2XXHHahCaOvnnFbwN9UY0kU+
/a1TXzW14i1JxwfmhoaM++7Spi3eRhjh4+k/JPPxVRDqb6r2pZ8Rf4MZnXW3Fkx5
4eiav1lOPG2Q1TtxI4nX0BHmP81o7QTCzD+uvlSYW2J6cjOWhLSiudmu9P6h62Gy
BXenGYdrdtRHqn89+S6qSk8cZ9/dKWAre7NsYmZmDMr0/gz36UlWNytj/D26VVow
QIFxhGvaJcQyS+QvHfs9mIT2nNENZ52PDKafM5zTlqCetPpTsfvgnsBscXfA3V8C
L5iqh8mr63uhL4MPBvBnxfzIy8betxDvDurqu/2p8+woGE+4JZ/588Ri2GIYACdC
dA06cbKeAYn1WIg5v1YiYWhkUd8AYE2Er4rCgwTInmGT3fIwYAu7S9QXXzJNrovA
U+HOJkw/fhoFCESOZxYpW6JLoVkAGJbMBmu/NFOG2q5G4LM8QtoG8QSehGjPSQnL
o9NYwk0676BpMc31BJ729FaBiS3kS0F7AyU6Icnu5zjwGrthrbumktueMcI/TV+u
JX7C/KZJTXBeLeNGWrkeZ6zG8GxyGSrQ1a1VaJT55GPORRXTh2dNAa3HKZGxwEZl
GAUJoZDDLHKBsHUNa+/QRt1O5p9QQeuppx1fVjq7/khI4EF5801ibYnyASpIvR0H
Ek39A2nuRZsC1EaIarX50/l5adtlbc+6J4KiPl1VfBgKDqd+biyEQZ+gV0qSfggt
ynnyBDlCqPb2EzJ39UKm1DCWcaA+y7Pbp6TzdjM4J4IJsNVh5kU6o6dZ35R1oUu+
CThry2xOIs9BLX9O/Wi3cl3HkeuQIT1bovuYq6g4Q5bLyy9U/hJEo3XzIPekPzpA
xs3AvgoNAgbZjUwDtT4uN1DRLQ8VmL+RTjmpXsfoSVWJbBTT91JuA67hTp7wWC6+
1RHaY9acDQyYm5Dn6I/F+EL5MfYKxEzrvLliHZ3hD1/zWbfd25OV4DPdXUfeLSmI
l6NIY+ptu/a6jbrv1RY+8EPZgrA/EaTMN8GVNJrIVsfOVFAaTtn/Dqvm6WXzjRRf
fdyOQMMaa+osO6JX97D4NM7RlufFwRhDEFrFZFcXo+V7BWCWgy3c0fDoLxaPrjEi
1TrtwZhZt6w8/Jm9sPCk4ztdaqX/+f98qY7V/akvG+h8HlF7FbMNuG8Irgvg1X8+
L7aSTX4kKPFDycPV1/ZTAprR1g31fXXlP6KzLi8E4F41YqAPrxofFDJxaXzNhVz1
ttoiYahobo2RcG38PFVudYusraxAPeokHb6BGjazH+Y7PaOl+IxXTJrv/H24CpL/
NFrjKU1yPtzqVDRfE5UvyDzxnp2pgkOqBWTk2Hemx4drQtdIu+qfOoIEx5xL/uE+
grZGSN16q8oQrTnqHzHLzhoYflt7Sc5II4Dly5HoTLKvcPMSufpCCYjj3WjW4leK
acdIjDLRuLi5S1YysNnXBzuR1fI5sE4FU7AvCmMgxCP4bFuNOZr0pKs9hwGzx28Z
DtVwZHwnWzug8I4LUJyVcizp7zxzD1be6P/OST4vp91GdyGeLRC2bhw1AO7yqE4m
LopCZItlOr+bCzXAMlfGyoajBF/ysTsttjX3BBm3wD4mIFjs14kv3uRBQ1yl6gLn
RkZjBzw4VKJCMuyobJUuWCKbeKqBW7s0MZxivnpLWKACR4eNbPnjy0gDl5oFAjWi
NtylK/Tid61dU8N6ziddI9K8UVC4eJRFzc5klSIXv73fbscPNrIyaFg1c26bteij
if6Onvp9WD6uqjD9SD1lq3V2JOkyaBWGObtLfXHVO8hV+Jj/JrBshJu1CzyvVINE
FivMfH8ncPY3pC1EpkdqSnFVoWYaHJbXgNlKLYMiVvaXfGstuYkQDFoq2I0p8oWd
UVKLawm/IwU7FkICJFbvRitIAG+V7FxeA4IDi24tZzSnsDGeAKKxPjey7i47AZxa
U+y0xtVgCq1GG5WKkAarVI01Eia8OhJcivp2CtVpUZzi0+/cN90Ps13KxFMI6/1N
hcs63VZCj6f519wepPHT3Ec1oSmMoaI5HfvEWcemBaHNJyc9NEzShtXHD45Fhc3w
qvnhUNmFd662zoJDSy2DT2JA1pxWwpkixaziLmYGtToyi5BWBs0Yh2AD3XWm70qL
Nfr94NOZD2aAyb+9n4QdtnDVSz55HiwDYtap5ulDsGC3tLQa0186pD7n770PffDY
tO8ggTiMbOc0+AfgpwJRsaiCuMzZ+eUJSZkG/8XIO9k1Bftc1X0ut6foBVizefOZ
4Nnr1woIlGsHBAWM3b77KRNH+bL4N4h+NCYTisyi5OuElrddnxxS6/UEeSIlASnf
BJ4OHx9fB/b7pTq6Y/RRV7kRm3lCjb7pWf09s+XWRQy/u/cX8WT1h6UDErf4cgey
5RoqCk6q+1m686ZsVdvwfi3FPV8M14kwPECY2iB9Jn1CQPl1mnWqQGlhR5+sP18R
1vTNGkTfQGnZuj9KywCBpJpP/2eN8cw1aQjD8ioT499MfpALLvAZnmUxXoBMgHYV
udM2L6oVnZioyCe04315qsE4fXps4r7bPkQjA1WcIpegcjdo5p30NXimlzYwj2bv
TCJGfc9eS7XKhePOjAtRENSV7Yheqa3b1Jq+9XLeffv2g9o15bVl44D290yQQfPo
p6MB32cAc/F58iLnC4BhnpunNi/Hbgn/I4ABqcqOdKxEqUM12shfBqR6DC/HZBOw
PK4F23wkPv8pdP+lpvVE2xDW133rs/3iBfn9rxaqWICvAnN9hFQgkUgqRfSvRnMi
jZll0y1xjXkmvjaAxMX9rJmfZf0Woo5LAg5VBzlUhMpCKJf4+ntS148gfLPVOXbJ
MWONTgAfXHjEqFFjCvOHCwLrHAHNjhrKSxsh1vFI176Sj2mzkJY2lsk6s/k4FLxy
6Oe5+NKKAKPN/hI6x9U7Aqh8/xQm3XlYdj/dfBudcqHZ0WdPev2TmBqudyRW9+DB
ykbvpDc4rJSxuKVfSTycK/5/ZjGPBX2hhLIuphSXLF35loZnO84sgiHpR287nNtE
Tpj+U+QPRS8LkwaRrTYNAkxKrttKllkEKjuyVfkkU4HWeAgjRbtw77x9I2itJRlG
IHIO1JnvHpxf+Sdshl0R4RD0YPeRqrI2tmxsyAqc5svmhSfPsKsUVJi/8ofabeZH
TH2kRQvhiqFapDSFPdv5LMWBL4ctB0aPvGmzyXEfecjmTq1oh1IyV4nYuLlXnWtr
Cv6wMumgfmYoWEKnigtquj5lbBid7yybqYLusilK4oyzsNSHwsXtZBeY2CEw+GWr
Z+yguNSz05n2g0Qse+opruuUtn7swi1Mg6Hgt3Od7HceJsGmrKIpg15XHiOfYq2U
b8WSQzZr6BXUbiHKatxVCL8ShpN4srwSHm6iY9XD0PDZDzb1Xps0xYz20EWEcXQX
V0OJXgC6Vm+X+ccl/rjz+v+G5V9pUSRY2KJ/JNE1yY4tlcB4Z1SO+J9cwMw26HDY
1RXYixgTAE2B+SaBl9kXM4207OYUnsJ0x9OAqSB5P2vPXBQt3GT1cBm3Cxt2jMBB
DnhtMQ9N06X4wKsZGHSdQnjKjFV/kHbq+SqDwE5uGuui8YgWd0qtddnaZrplHCuV
5f0dfVv+1MpjGZfOAcMuE+5O3XcZnOK+Aq2UM83oOihvkg1JjCUqQk8isO7Gg4/5
PW1Iqa2ePXh2GJow9nO/m2zvApkNfVxKuwQnSefQLgQWvvUJc12Eq0u1DvYPBXsy
+fTZErTYw/hylQ4LnaEz8/mIUNZ8Zen+mMgmmp3ZWqmOqdEj8O7kQnpHGuageQZs
Cdx0hfNtyTb13SYkdWohRlhxdVwkAa5cSD/uohhMR4Pz6iJSsPo32IT9TJ7ba5XQ
9khvZdFHhgYJQFu98Al5O5s0Oykd/3WBMY6PKpQvZNgKbSZ+qbY4mXCNfDASUrkT
av4KOBdgRRE7s1LQweJ4rCCRDEKs89wZ0yB6Ex9/6bLK0aFjbDkFpY+mKHKH7KF3
9p2730DoV/FAEinlyEd9OoLpRDPXi6dBKnmaBHEC7nip3lDMltNsFHyvFQ/J4t1e
/yolXOeYy46Btojc2xavV8vo1Rbs4c2B4J9ctqwkqig4jRA81S1aJc08GdiEY0Fu
BZzKDwcT4UGkLg/5cBViRP7xX0de7Yz61ozGEdqMLG6rIqitEhSeBb8ZUmn6hbBC
VMHXGov1K61dzjP4YT0zeT2cr9DpChyJMWQOL+ba0mJiXzUlzxWpVflof9jGMfSd
chdshnnymJu+aYPtL+BVchIXYRlpKDGzsDN9PWLkr1JBo6Qwxn4kwg5+WA5THjTJ
54Ip4Lop933xSVIJwTkI4Ui20kDLdqwHv4PSU/Lr5XuC39vVyiQ5Pt/O3lYiC5DY
9cIVtmGYVL8jEh+04wOSGu0ZhNWJ0lUdzi0a0xeo2JfkkQuRv85egw6QaPW7kMLP
EluRnUyyWLR5oGQchoFtKfChRgVzelvCU6z+gtavAO2h1o6x6jFu5RWiR9ADf4gY
DbFn25UgWmzDbR5UZwFg3BgJ0u3w8IUn8XXU2vnm9zyAXMB25+0a9HyRaRwtn1HV
j09Bi4zSKd8YUNatoLjkQquS1BHHYVUs1HoAltWkMNGWXigjFUo5WMeGOsljMuu7
BPfJ7hWHw70RngxJgnVu9sG54Q/RphEfj4NXQEu25K/rB/yA/ykfYrsqcvssVck+
5Jzr236+mMgrvh5DDlY7jsHlpfZ3RHy1b8b4OYlWxUht6KS+XxsukigKTUclyqgu
ybj3qs0/mK+wdFXzJxKqni7klXONEr6uKv7hmkFqVzNAxeMqhUcryuHL80CQivsv
PeCnxMgOlyVYPfmMf6QWxYBxd944oj/ttUL0Dj+lDynMrs1aZqeNn7gX6k/qdXRd
ZAH7xKNHkELzFe32LhNak330ZEStQNShHfUKFY6OUPhBsU619y+hLetuoIqBSV3z
dVGpXU2tU6fs2kp5RA1+rV8+YnVifrcj7D2iU2AoDrCZ0lMVD5XvYBc4011Xs3Ge
W05NZg+kRILijpT8B/s1XmesTt4sJs0PSpJEXCJOrd1P6VZaRdM+84OK9Drwio1M
oXEFgabXsxIobmuHkZCGfVR55KQlG/Gny8Jkzp3x8u0jq6hEsmk5lq4E8C2wv9Gs
uZQ9gZ4IjJvv+v/R7BxIQM0lJgOBA2SEQr7G5alQjwWR7tyHRoT8yIxvDJs2muiF
IXJetnejyCvLRnzSpSb7go4pXOKlp7Qn7bz3EfZgoaZleiqh0du2sHFSs67HaxgM
bRDbCf5WJrN7wd+QcFDgWyvc4xw53u/2jmjp1S4TCjg8EPezFI1tlrDbEklRU854
qzeHMeLCvpTKPUORDw4DR7VLgdJtIYsmOSSn5Jyhj4KP3eE1DbrH1ef53e8wk0qE
Dyt0RZ/zV6NHcInxEEzJ4DNtkXG/sbCKA7Knlj2z888M2fxB5wenR99dwykTeX1o
tnURUWogmQoHCzDXKX26XCvhRKNbwGb4NwtRKCYSBN0gC5qRrpq/Pr9656wx0eH4
9dj5TD+F7+thfcx8Awnc3QEfXx9rJpnaysVD1yVqQJsUQ2svSJTkJm/ji21GxHJO
tkjqizpTFK4HXicwlCDmwh/iCAb/4E/pVYcTQEAnYvgU2+i8GGeVCKTrqjms0Qky
x8GSsbDDfNV/aeqjsKwPn6SObUHTnXGS/IOrcK46P5TxQMQzQ/CDDAeQahEFIBQr
GVKH/GnpPKwFwQw3G8YxdUSBPriZjd//JUTUqaNoAYhCUMG1a2qUvlW5o4ucgbuh
vaxzipRJdNMcRkYFdh1PQKgTon2MEL2y+RdBt4Vt3hylwDS0UVK5EOUoWg9cb6/K
KYr9XpR+HPFqTXqeTezERPCrVnNPATIqM3EoFcNd/PcvzUN7sgug9wuO7syFOV6R
2ej2uyaiQr89N0StOGQmByU6xS7flV9GhQLaqYNYt0gQpClt6ykloWuP9VS6J+Dx
iA/7PKvquuMb+X266tPEm5Wuxdr+FY+TC7En5Mdwxj767DGwsoyE3GqKWeMFqmBo
sRAOwXyDnC2wm9Kh4hI65ORMc4nN83E2XaOdDZuEFZCL9a1DmHZAJiULWodDw/LD
d9TKaIS9hO9s+TAiZ2fquQA0a1U3ce1Cxi1FkFJyEMpusN5fcmet7E06blvZ3c9L
TRBlY/9ntpLb6wOqtNoaCOve1MLTWd6fRIGfMOrJ2jFRUAQMZNJLzFN2zojS1xTo
1dyPLALHI4q+miYg5Idgr52+wCz7hD+7zIp+dKkyv9nh8YQiudVCn5/fje6kQI/s
D+0Q+ayeJARuQrkyBQbMPVHxUs7PPrlcerj411KwnxUgCJshC3owmQvVx9Qoc5oA
jEHvBkRtfBZbOKYuMx/9zSxYmoqiJtw4Vhf0bf3YqTZl9HW9TN5521Asxfit1TeZ
Dq2lKGuFN2iMIf+srJw5Hpw0qaXQSAOx/fSpDCFogHc5ifB2NlfZWLb1RV9Kd3FG
EyrWptTXCcsqWVQe4cS0mUeFc3JuDxZ7Cw0hmE9i9WaZdJe4Oz+gihqYxMOb46RY
9lej8bexOe9F1+TVrMoYeNA8CnVRg0DFDxmllje8kxSnlp7XDtZU2XXgbMSSizTN
+v850Gc4Irdl5Ij8NN+1UYdfr3OQb0alksvao1lpVldDio2kf1mpAZDRqQFhcSDD
hWchx6dS50uzkwQl3d4BJjkLM2mH6QUQUQgrgZQM9nXfhg/jPrO5xf/x26W1tlYf
hhaALZuD2s2yxs9fZh7hgT/GDFdFD5d5j7YP7qAzmpgx7jxPyOeVd/uPD9eXZfR1
1zZU7x+S0cqoA2bVI6J0Ff52kibELjAwfUOxDnVFS6eY+nI4jsc+fxvno6jTjAB8
2C4Y6IaQuNBkA6dEIz6G1wb8+7iv34UK3o4dlGrAhd2tFXG8d2x47BBOZfrUTeoK
c6PIbxOnzVFY+AZ5C4husKG6QuEWuxwAV/3oylpKUR8+57u5Y6DMC+FWSBYQVA1x
hb869tITiE9soH+S4Gclx1RNUXbCqJfF4j1468rkZ1vxkWpsfhSX9aAJ8/3WqS2Y
4pd2kUMXbjQ/PZHEntMCee//bm3PH9gD4U4EbFG4rxbaXCHzYdnN40p7yETn9huQ
BtbOw7q78LzfTmmLVszpd6Yn1kCqrklrajCJx+Yk9wJ+gAZQ7hEdWAOi0/RcIKLm
yP9NcYTV8yMPWxa6ffSYwSMkgr17p2Mwy38KmcFp2yUHrxALxeHw+xTpV/1JsRw4
W5uHqlgCzQPqyz8qn5YzFBXuBP3zsxV+oaLUx6ncrnE7ZAhJDaX8caBZfGdF9x1P
wag01oi0R8q75PYsdOv3cEv/bagjUM7z2vrKr//E40/rdULYptxbXGMLfJf6nERq
BWrDYUJje/cpeh8MDYACUafbLbvggA68lOLAhGWI9Z1A2uMhXeRsgd6W8BP1uasU
snmf2/UKPSLms7K/6fooni65TThk2oF2sO6PT6MUOF0ZSXS/JZFgGVHKMrX+lkh7
VTICa9WT9IRku5VAGbhO/ewlEj43vjxuO8X0pxH8i2ciAvcS51cKOjXD3m+SjlfM
9rTUSHs4RusOzFcrbpBH8arUYpZFFhmlE6jGnLzHUCFgee55gn1uDEtPqTJtybXR
DzVZ5uu2TTwRRKncxchvaBx0fA20hfWC0+MMj8seMUD1AipDgxaQg+X89s4hSTdS
sHp/xhNbKBcWy3A4wp8k5TTw2aTmDQwPZfDK0huNyvLU6H5D5wqRQdDEDtwgX1fv
ZmDoGlMFlGLIBgwcERMQ9lgwIxORsFxTccQGweCzzHs4vr2bAA6Yq4c2XHC3iFeH
frM2WctErbYBO8FijnIrZBq08/U9CZSRy2lSQ6aFhvP0OGYBk0P/EHav1d4aylo6
QoBq7tpNMLxL9Y7BcaXTACKvokU6lTwc6MqAx59zwOuUjqgFOQK0WQZehWmDUyRu
y0PtREcq6SflbC7dEGPTTrlBSh6A5eOGvcEp6TzN3LTL3e7552mGd3+ZdpHVNJBT
ordXMfJqwfRGE+KPXGn0xtcWErcF5qMI7FiAQgx7iZiRaeH/Lm8BI3eBQDwnk8NG
TY6/gxdL5TT1pVBwcN5SDLWB5vhRO7JTPGsaGdI9KxhY8d+Izn+6JQB14w41sylS
HARaBxdDxphpjqWnI0r13czco7fyqezZScTwZl25evWrM/C5fuw1vKP8xfejUwOU
l6fCTIfyXHEoflw+cNsod76EJovrVMVWAGBx9B0qvDjt3tTq/CR46rzOwOWuCShq
idQu6BwUbKhTO0aJPE2DRG+6ZbwvebmCxlgdSOQMpkC3mX+ljoiwWNuiHNuG/V2E
4F95/SasBGZlhKUfHINITaNt/o4HbdqHhb1tVTr1tYLyTVJF6SzyMEvDecOtBj+f
jCk7URoMPPw6JPv+TcMCkTPiI7RG+yYhFPeGNvj5xkB/hOk7aanS9I0XlVwEcHC2
h8gu1HjJQh4uj6H6H159QCWtEuw/bBEHK6dd7lTpfm3dXYAdjoyAYjxSd+nJgw4s
CUMSsJU221u84PHtTh6QhcbLUgPcLjwou/jb01iR3JB75krLQQub8HqXJ/jQNtD/
Ewhl/i00TosDJXLdfDrymV00S0FttasssIp5d06FHcF6OPVtDNd1CKlj1rL1HcJ5
BnVwIQVZxKtYiBiKir6+QU4ZF9ukjYjHT99KAmj5rQFogWBUds2bJ162duqNxIxi
FgJzucofjI3iLqXiXaPAnD6Q8Ch3jqHlH91XXS38bgRXBbaHnrXaQPGA4RJ4I2gz
gfqHfZB9Z8VNYwU+eb/AxfspxCaV+lErK8wqfE5tYVtWxHCSunwF7h2Js+GpcRWa
t2XQ5tD/Fi+E5VpRhI9zw/wYLnDVQWYRCNxeHYFPRAJq++lkJ9iI1ZEsVL0qZQ6N
kZoxpj/uVatbQrBePB8Dk/PN7kP+En09DHopjyHFHhDsol+k0tCTjje9t2mF1clH
Tyi6wEMtncTXx3EdSWix0n/7x+hzuFYFDBwA3yIn3E9urc41IPmmvpE9NQCxI3NV
mizXLUJ6wMaXwVs4eKwAjdQjGe8qOQAmq3wVBzaYQ8LJiW5n01ZneP+5Ou8uHLGX
sge7GIWQ4hT/b2MF7+8NTbGP3PfsI3h2f94mlGE9GLxOM/BkkOgd14L5qWpcCX5M
yRGoMfbiJ5x+zcfcUbIbTXoCEEJX5ZMFIcUrx+hRk6U0QEwNZbmOZwOVTd0yySR5
QfCzvuzMI5YUZmpV2YWaFB7SMUKF0edCun2lAzCyEbixHuRA7TvbWaT1CK2RybjX
VabMy1nrlXwrgvIojHi8Zl94BJdcmJmkPLniIs06nTbNxi/S8LkZui6rZD3e0BNo
mWMv5PWYQHUTtOr9UkXpVZWxRM7A7+NQpgUpU7uCx7ABt7QvkI2CvZSCvgBrhmzv
st3OsVl2NVpyDfpapwis4lmLuM5ReIIsY9lxZfMdp2E9D3HgTh0JogrQc2sWdmQ4
mN1SJMFxMGgSfGktI5gdZh8b5/WweEJ+cyC2biw9Lw6XIoSobXWBtn2jgOMC7LNB
ze+NZtsglmCB7Y542BwRT6Y3w+DfZWi1vf3LF+YlvF4L7fQlUV/Tp/uQbhYst+cv
NaAg1qjq+XUIuzl+3SLcNZspbkttBaGKYwQ40ZpxKlkFNfEMLNqZAcvV4Ot2m6Bt
Scno48nn6fVsXsp48iG98tOogOgdphcuwUJ9iZSssnPzvVrOtX8Xpwb62dgCZxh8
LoQW42iUJPHba3pi8DAJtUNY2JABCCqWTTk0a4zMmB/FvDZh3BvhaAXMcx12+W/f
umwcoR2w0YOLvs3TbjcvGZAj3veOuLGAy1C4OXGsgf+8aWhY4dmERlnik9f0fTD1
kjQHogNuZCwx9ROUxhPDFa2eHNom0P++XL994c//Upx5KXYkoOvU7CtjT59lxO1R
aH2yX3eMTT5YtDFTIPXoAB8wyMlLa9weTAFCWACDaymsG6n1tjodfwxczqAtl0Cl
ND5Q4HbvGwAoWb3CYStsrC5lkUGJ0KV1d2Nx2Yf+mPd2itdazpzr1kMzcFx1xJQr
r6NpIvvDVKEMYgys0iA7f/xhIettrrCZwNIBy8IlT9BHBBlWFJ5o+LL29UvY6uqX
+S9TSrh5rwRzKMWKxR0mnN0Gkp74MvNeBX/F2nvgxscCcrxev6izaEh2g/pomuiU
uxVESyLro4bh89+wQqmOZSMGc2Acm7cXS8DDGUy6gLM6DXPEUOpY6DOlO60rthvk
9tVllwGybWc/BxcmKCcKvHGDMClS/jL9H6Oa7Bxf6JeZwFB9UbUblHfXSmX5iJWl
NwGRfjs0EEAMjfSVkF7WTBI51MGmsUqtvFbBbadnBWSfkigYb8mTCIGvhKdisCu7
evnU5O1cgD9jo/Mrrt2nM6TuI+kDZFH79NDqu3thHa35IdmcMa2jBLGKq49Tk/O/
AkhxbxyCbzoSyeJeaDs/pCowCbWiH+rdKLXayAC7w7zmm+wRTZ93fj2Nn1OWmxu6
+XNsnm5ruNxCfT/ozmn5SyVZKIYr1/65No2v6XQFZPttKHjRub8sK/un8BSao2mt
qDriS5XkhvgojOBuyyM3z7V32OQ4LUUKQ5TbZRaXHSu/eFjShNDBetsu/7mv5g88
TxeNFff7aGQzcF7KPbwsZPk9bOn7pHm3veV8leP82oh8n2l7PlZ5v47gADpSHuW/
ezljQdkriVppN0iGleaqg+Z+xQdjpH1VpBcAt6ouSO8Gi3aq/bXANTOEIMLsBdH0
kcl6wOuVP4toE8uNusVGYH04XK1NXt7okzKEbCIjQv3JULqO6gClcPpWl3m8D5eK
ciElNRIT4LbjpxW3y5QVMk3roBr+YZY4XoUWlggBV3rrimJRNsCt0hEh7AnL3adM
3o1vkwODfAJ+fO1QFq83/QhjS9WvOaOQp9SpO8il7vMS9nikXvXx6s/aU5Ac6ggz
5gk7RpZ5SLyp1c2qvIfSG1ePiOmHrLZRplY99x8UmuAeUlxvSrw9GGTd0VEvG1E0
ehEgWWUwtwpSd5HMazuypR4nyE1u82oJ1MmMu3er3gtHrDCPZOqFCrFbbsG0g0hk
7WxEbyGiZSkLKkw0pqfHyTNJ4hXweUrNrQDIlSouANquQdX9KU9sW/DdYJqWDWua
VgDqNlCZxU2H8OxKmyLY3dIeajwdcxGAFjbWHlWSoQh3y9uTwRuW4R1yxfRAj/Xe
SqwSKa1UJK2dvlTCxTJUtZPXfPLesJ+1MO6rFJIrPVJiL4cD1jIBKK0Hrs4emw+w
dGMDzdlk7QstgSgpB4mfm9ZnatoLFoC2XyyoXT+wXGG4/5fJiavmcS1E3TQVwUqr
8vSznjl7744xUUDToNd70nMNw3v6DjaZ/8o2a7jD5esRYxh1jk9vbVUrnQWCt58W
npGsfU15gSw0tSPBF1XUOiUNmvooVWSzugkixSns1BAx0jzY6Bspr5MtDnTxV3Gl
eKSMT5RsG7932SmG2CEgax8Em5jmOJP76mnpfiuE42sJbEdq3KiIR4HfcZhKoojb
9antK4SoNrU32SXpuBAIfVvvy06G6X+TT9Zr0BO3lK73J643pfRShxZTV4tVccR7
qhrboqL+4J2qH5sD6hgSAfEEdaKl3lHjO3dv9R52lRgk5Df1MVACM/U6Mdu2r5Lb
N7Np6zeaPbQtG2Zgp4zrgDA5S4woMlrtqNbtwpq8put3/kJbFHiz5yCsPVRTW7KW
EQj5Ds93LlC8dFcQgMfZ5kBmWZ38GCja+9pMHIahXvRjsjtddD54XLVxnFR0g1HA
TB/eY0tUVxbmuLSg4fYH9wT3l5Wk7dZCXIB0kfty8+NVJ+MbiIjcmsvc/er0Tnp1
5Jp1qrSVXUAD4liHlMEWTJAIOpEI5mLN8rMOCWkONYygpQuAChx3J0yYLfvBpZje
yw6iT3k3MaLn/XI49QX684hQognl7p0B9mWazmcYfEXwZjwJQiD2KUFJWnzBTBqM
HwOcorepVBZnBHiz+m7N6Mbe3UvHtdtnk+/gSWbiXZX9AN2k2xgxVkqq2ojV0BMD
A2zao0fV2dGDxy9PZDKxAyLnmBjU4QgmcwkibyM8KMc3M5BPnpJRLdXZHmq3DWSa
KEgNEZfT2NbtPzeGVbF5za7hyi0mqjA/om2ZmWrIcclTgndrl4yrsluv/cfpAkAX
Sg8OFWIW3cKi6DSX4SyfqI2D4LHP22LNbDUzOOw8UHEBoCwOsjjF5zBhzV3VGNdn
66ROSETtv91kR0ClC4mBbHJW91yg1PxkZxRZYDV0WLrG4Ph9TEcedNMvg3goo7Fw
CWKGJUHs30Ps6PRf0ShpyWn7BRuJfnSnnotTojz7vOHr4sIJm0vnBz9/u+bX1pYO
MH/CzINSlAQdKaQEiVXTG2UhUdSGkJAm5SmUHC0POU5XPo3EoGMf40ITDeyD9Uu+
SYilPRBJ3ScoqoYRwe/vHNm1wJveFiGCPFvlDf0LE5AfYo1ohalQVxOljsR+ENP0
M8OyDBmZE+Mst1xwN/ozh9ghYWzvzfB4u3zPWqTQPg50mlacM1oiVliL9JE0tCCq
SlAPLLJdnUhXRXkdZkd7elZQnWxg/MPmp0ybKJngHwhLGAF6Uo3cSYqg9Cs5KOEQ
gL0PTEZ9GjssKVKSvxJTnJDZz+83z+jOGrN3qPBL5SqVQ6/E6LRm7a0rtAr4xBV0
r77VIG/lk9xRxyNSHAaXOrUP70PgEmNPei+S0x31ChsLpWciKhhAD5SsEMnoAR7l
UkN4dwgMYfeyIbUcdGLulqOAsIvH97bx/VsbNNCu0MM13/YKUH/+Z0JiAOf7HTdm
96gpjOsC+rqKekWhCQd7Qp4Pbn57ayJhM1bH8ANaXBHnoQMw8pF1STsxTNMuIePw
+nghMAF1QI9zEXhT1LqkNhmUqWhhShriZOGACc5n5ngBedtruzKM8Y8JeGGIBki+
UtZUNiT65GH0LvJN923xz4t/FT1PqmFOLxFtYgKtXVAWYUJINboDzkNQ3rAlE5kO
Y40T48ujkz/oa36lOW94hApALvEUOmu2Mo3sOWFfbt/2innhTDN5D6Den8LDicYp
C/Y4qoYxmKioA1nbOHuUbtTfuvTsolKwcp7+4vJyAqz+CsFSPTxmLO8M/a+WUfvG
3RSu7zjz6ckWnc3SO8I7EQ3xsvF+9EeZfq7tAMXbQJFJypMLTayII+DIVt14ylaI
7T00kY/KQGLEZB/c0uHA4Xgf7svjiA+cYGkPI/cTw9plMxIIbs5Ss2Net916Ssb3
0lOcLtWfwyjHyCN0jq7AFPZIJRAuzQbZYS/N2wubKRmdTvn+TAIvDtkGpn83j+J9
TKK0ZID0goVYddC+MP/ByvFWlxiwXBVrPRc4BOlEGxq0pUw8YzlZ1oEGCbTaukkc
3XI5hvegcbwKBAfaf5M7HCf2IjUvbO2dInVppqwI9+ryPyNTSNd2Hf9OTwOMf8MB
Z3laLEBeshnsIDdUVgAXUxjRfplR8P7vgjY3R/VoNdCO36brI35PdKxk/EmQzWGD
CUca53pcvvRmncwuglcK/UogfI6aR1Q2XhpZuy+0/W2yjM6pwQoipZD7xw+1l60D
QoE/0sTXSu8mnwQAuxSErcLq0r2o8A0TvFxwGzspOGBh5v0gOo8kDVlJJ0OZbqgV
EBvEvE+xqcvzypPiz99YDw7avPraSKT6gTP5wUojSejy078KZnD26obxTCk8o7zI
BvnRTDKd+q9Rk4hx2pM0lj+a5L3kxIwk7p4BBpPyw+HQCSIfoE72ouhk+uuD5RrG
WWhLMMgr5qLOZnWMsJ9kmniMtpk+qHCKVHvrDTXnNf3A+3BuE7vTjpMySfpzZXrz
XXNqkX/KahuJBoOiUAYmOxh1ziutA1XbsWWg5TN32IREh9hURlYuaKf/z4OAOpRH
EzGJPl/WcjjkJHqFczZizX9Mi96fge7Hmah5LpH0ole7dJ9+AfKc9YKj5LTgx/Gq
/sVzDkBT+XhcI+d2splcA8yxSPC+7lZqDjKMgEi7y6akBtCAlPwuqBhogIT/aWDJ
riio50cocjOf+V6MDZbyfCwKWlwEMhoSpknwl0FplsVKhxaCrhyO+ZzYmPYxfSiy
kXiPxyWkgOBZKMj523knjLKYDYyMAOBs1wBwfrThEzojnv9yN7siy1GH5J3uYdIl
9/yWfzdDQAG6YIXb5+Zji9odCEU89NeI1ZGkljzXJZn7XJ6j57KpFSRkiJL9d+kf
R5IUBmiSYdaksrTuTq7E0UUIC8jW4a7cBJVGrkNJtS30Tpgal22vscE9IFPtFbqL
/0PoBSwrn92EGA5ik9gBRp5nZ9HBdC0Xzp0eqiSNeC9LyjQYu87zPBGvsmt2yHpM
U4LQsVDBpCmnBkKnuSiDFcK2MlysDw2+f4/iyjcZLAKuam6mg72MT5Z/Xmo/K9zb
C7pBvAChH67HDtGCQnGhyBrDFs0FMTqJvAeWMr/PzEGCp43Nmrk6XqESHi2dQVX0
AIOT75K8jcAn3mogCqL5PfOtCAQGh9Gdhq9bw2/AJiOv/m+Q0E8a8xQzMm57s8ZH
X6PMZbPbR1xzwRiB47N7aTSjjCOBOCOx9fa0kVvh5MfCgFqZBzT1yFB9Kic3oEph
LeVgw2dCDSLFnoE6hiotQaBuQzmyCqbZuy82RWwcY7x/VQEWOfuJc5NnZKuRz7NY
NRP4L8E44ttiXsGLw7j0Z8JkZmABTWsoaDlvoNEonhA4iM3qBP7DNr5G3DBmA5n2
Vdb8xcEh8hrDfaxxmjKN1tnGrpEhuGeEIyW/MWN/DSXMxgujFgFitR6ytd1Qae0l
oVhFRPvIsroyHqzrMozcXxXbWyixGMW8W/3BfdTJvo6/ayP0ItHzX62TioLd6T8J
blDSHR8qDGIKzfnU64tkPdjhLcYOvs2+3cl1ph4U/PDUZF/zGm9ha4aoxalWubkj
vdMsBn5wq/lblxgXd9lpTbC6toodzeLGVkOANhj8dHdaZyQh209MRB/b5NwmDYYd
QpcBpMDhnWsLFrPgFsauzAzgcMHkf+hRnfwIlhlHB2Efmmg+Qs1/HHMjGGm4qA3s
NLtiofMyuuBM/wXNs90gRhg0/b+ReI4460EwQrTmsSozkffMeo5L/paVoE3WcpxS
Ft004ENtynftOsEZ/zVPgYGBdOE/i9hvXAjBZ1aov7jqnb+UCfVXblMzdWZTPPpm
yXbPia06t6EVvIGhtZBBZ0YKA65cDGCrdYidLy9iGrp+p799H/417e6SU8JFJWSn
z17ZBSujzUhN2wqIZs2THmUUf90pZ54z+Vpag3Zutu50Tkj7euuKZwA+I63NKHT+
PZyU1aTKAI/p9Jpw6Z2ri9aN4kBeux7NP0ReGfEYQl9u7FdGSYEY9PV0IvLA9ZqF
9FgARejDaFnPx4RpEWBUEovMbwy0omAuEyTawEvv5eXou9nTafZPkkl9KXXoE6Gy
Laq6WHJQk5jX5M83/EZDULN0mhhvOn4oTOTtMzN9RIR/Dx/JCVXeZaAfSyq4pESJ
1g4rqUmSjezaw7sCAYdvboRk/MlEpwNNmZOFHYNaSYmpnia5GANYw9v4nKpMl0fS
LX7FCHdMDRjkBBif4oo845KFD8W3jdj/dH7XUXv6mITk57fS5mKKOzHUnbgtVR/y
il34SVW0fZI+7Ql/EKdFvmxCHA5Y4Usi+2t8tGbEja5yUuIplikf7UwX3azhxztf
NV8QJOEg5VInVtX/uNGB7oIOT+/VOqqN6G1FP1WUaqDwpyqmneJuJO8tAadrMek8
1xwQBDPKPR8DDI8vmZTkuGqP7SLpUTW30aazZUXvjKsEAWhfyKGvO4ig0e2MHQOu
Raxk4gQEncopK0xn8Vb3kiUuiM46YkTxa/NTsaJ/etcajKq081vfhBfWCSRbD/Af
YcjO1aRu2OLLEM9Hoz++L08xyZjcoKty+uKz1JOUpx3+cReM06FNqbbDLvBeliAW
0O2ZJ2P1q4bBLqI2dLbD/9N3u3TU+iuARFxcoIGiwsipA2dbng3N/OGBhDERFjW1
9cK4G+m3IbQJid/+t3y3vIDU/9FxweIIYgD367R5qRNsvj8IkLguAglMKSCw78mS
DRTf/hOsBrL4yax9BoKW7JSh0ZrUZw0zvsm8o/k9Cx5wAnZAP83WtvhOCfPLY5J1
8sNgnX+4nNmCNrXAOP6CpVfqw4tUCHG6r/mashyNIh9CiNfBTZGoejKT8kCA+xn+
HaHizMVkL+lIzAKgBjdSLc678WWwLs8ZaFsQT+4XX1iP/inpRUIdtlUOdOBLB3JM
ZZoyYEjDYWCPQFafZVRUwL5/VFfHfMYqw910W8RYFQR9WJZtYPwnToreZePJtVl9
JzraQIzDGMu3pS7YB6DA2LRDC9fs+43RrOZb2oZLjpuF7OiqMVSOTQBto7WuVZ0k
cOAvZiFqUG7M7KcgHgMjosudZkrQHh9qHVM+mkZ19vkhUaWOv8CDdQWlGk9ER226
fGH1ub2oaQQtO/xJYTu5UStYLeqN9X5Js4IHPMptUGRNeVESAEElb+cNa+cYrJbU
NecptcznOjj12JMEnvRCK8ml7lZNGUbqmmfLBL9kxsu28qHm/0CGQ0Y/t317XmbS
MSt9zOpuD7Txv5kSC+lPkiJHJO1FG5OfA2c4uemxjTNcfrqkYU0Ik6GjsEUf1nOJ
lkpFDNDyhd5Lr3RPFwOsuC7n1ruTO80IKd2JbZ9/GAsFpmtrCvBXiG7fQT6TAfT4
kSs198nHNnVRmdVGIiejMvzyHE/1bfr+4ycTcGNNZnbeVyvY08WT0PzR4jtlila+
Eh0kR81YqTvjXc6/DbrmfevrC8mLE+/EtQx3BHQqek0R2rk7p3WT3KHdvYrHEwLO
x+Ii/aKPJsnZxiXJUKwovooc3FvOOkQ2WzTYWHBK9R/Y+1Hg7cY4k1NNf+xozCBk
ychFd/eOB7kYYHB1B15bwCCq1H+5lULHlYY9jPNgoOt/VHom7px7eb9PRJakiypR
CeaAgg7CxEt1NbBJt55Aqc9BP3x0kXnH/rLN5dxLzXBL0HVgtuiiwCyIJ7U8KIVr
8twqTUHKvrHL0ODJvjV81gSOrxLvS83w5jWscyq76jPauHoc3mJ/nFz6CqNFP3BJ
CbPgoEklWjEPk4U0blUDO3Gy6gGX4UwMd1itpjS70y2z/cVWPpl/C2VdgQvU+nkC
o/MmmfxchcVpImVxBi1jj6m9sw9jShjhFQOnhj0wwQbyiFbpW818BPR0irEwwn7S
ZUINZuQSRjpOyX+Ss3ZDSEBiom6bjhs7V3jnD45hd5KC/GtkE64Dr76Hwvm8FfSp
8fJWni1HYpVXGqtgCbkhIn8/qmuChqxYZzOv4gXPDDS64LucOI0xZ/xcsXwvCflv
gLoXjd0D7f6H8UGkKPQ8WmJcJTHP/OzfAAahLkprNGa5kTr39wCtCrrH5kzMS8Zy
AREAtZZDLyg7heQokYCcJETgAmtEbuwAWIpoCtLsn6suJtEPU4l4IhZCFNVyqmBC
tVSqJAa9EXOoIxw4lN1uDhkr7a+2UZeibU8C6fffWTqsJiBxzAJDHwRvd4CHRslP
4gp4pWEPd7Xz4xr5CTIbN6iJzNIUjS5OZc+M472R48cHQaE4zX4GV/jixG+tGm8t
GkeeS0k2MstgGlBbt1GI3Ko8ZdGLnHCdE99lVbZzzsetmjDbQYY2NoRoPepeyWCS
qT4xq+7m2l5XswK/h4/HB7gzIAYbESQ4kCRk5FFMPAuDxh7UPaJ5sP5JI8MsATU6
zSUvXwsIabjpiYN6j1UTH+YqQjYgB2YQxbzeae6xr120rZ+vogDAY6qsP7+olPkq
EtvjLxWZV2MQnJFPjs+qNsOG79iiPiS2A4hT+4zL3vEbM5G6Gviw/DTZIOx71NXz
h5fOgdSEgXcRxWmln0TKLJAffPrv/IEkR9jx/7t7lXWW2fcz/UOLq+VnG8hHsvxH
Fxc0JgUKnOALV+XDi1vfuBQyY083IxzQZX5cyCrszyLv2PAnXCnKnTC2srtAn3+b
AZyKF+fHsU/WEhHq+WNPDaJqZBozv2FUac/1k9xP1qOPv4OsbxQhn8f90kMY9cXm
vR1xh8IL8AMzPouvSp3lRAHbuVfhoOuFaxGasGEJvij2wGdWgBJ1G7jLv3PqUv9D
BID1d9aP2vkmAG82uOMGTwYtUJNNhyJwypna5CopA2IXhCrzw78ROJmfobOk5x+Q
8YU+HEPs29mBSU/KtkCShbiXVfxjD2PNrsLpo9XlSu3cUqRlj8ZujjPielPt1YDA
fgmTeShOVokBg+bbfeUAHN5fEbkgJh+IWYGvxfceB6ev4+qGWkCIXjF7YRKiiWNP
XjfSPyH+58PQsEhx4Jo+S0NcCpMUYUclRFnzlIuoCylKMW0f7bDNA9JzXMN3V8BY
9YnDWxAZS055NU4IM+yDcKrNTq3f/k0TjMH6LYu8Fh6MwgzNR5f3tvdD4FPtwzTk
j8vF9bfsQIbbv0C7SN2ENQ42ma2T5xJTMajxc/ngzQ0ODa/uHMUqlQyXLgIxFsul
mm8+1b9+hTlJSXQOjYK9atej7pcdZPcdzGF/CtVtsFLopRVXoBScQHfGQhIEZFwd
eoP1xryzWRyn0jyZX6FYGTXoFyOHAXfbBntA0E0EaVoraeX5WRhY6oH/qKe6rKvm
kZx7acfd9g7NGFfKdVmD6lKmktOT9lMF/TJen0CRYuyliWyJIM79DGILj4v4x7mw
x91RIhxDVyoOp+n+1d4Aaax7mrqLxaT0lf1wAhfKCtdkiox/pLebYbnHXDp01ZGP
Zh/Vrj6fW0csgoFB1Z6pIh2x9jglJmj64S4r9cbpt506fxM5CG+EKLOQtl2ZUgCz
tYf5PcR9hlExTy5JvT4ia0GNnz1F1U3N1+8Pp1llFnxnlsGm2PGnOubDwmCJhhUM
+GgN4s2iYePg63eDzatk3QWQC3UylYZkzYz/eacIe1SBCw5I0Tc8h5VGVpFtYbJP
OHRBSX/xZJz2O1qJK4AZlEjSmNKMIdC+SqS4ZGN8dC+s5MGUi/wd2EM1aL1a0EJo
LI+arbBuOjseUj0Hjxs+MW9mpwdkMxDkoat5WHeom/hbamjePCc+7lrY15K+3AVC
N64HZCpUbXrtnF8tgOunRG8taDNrj98Zk7jQ6jXMJiDCU7C/a6Kqn8zXutr0/kqJ
TJ6X4c4kPeLqNGJfrsvOMygRvILvSO3t4nSsFyOHg3ywiemLLkRbaw/eUl2AAKIl
6ZWM8MkHsifj1rARLN7Yk8++TnRlragf7FBQyT9XGLELW3Uh8xIi18yi5Cs5zENd
gfN8FtJ6rKQfOeiRilyDCRqFUGw5zCUq2RjRpG8qxeztFGimE3YouVq2RU2mjwWf
6vYcYSTndyPu/FLpNTHLlPlyiN9ETmCK0SbMjcdYOhcC9n5DXTCH8uhJqe2qaAkT
OAAMduxYksM1jm18fO8NZsnKhPlDHs8kLjHeIjPqp7s5k4bEDfjBTQ6ioN3NxbN3
hrA2ZAJAS+zaRjsieLnDIL2+ayR5vU/l2xjZlNR5jtcyKrdYbB/Qw+bCQxX49bZo
d/awlg6LfkX06LEQHo+rYGIiuVjLBBiromaCL5X3P77VWjzd+HMc24ALZ1NuG0Xl
TeDximsnx3E/YhqtChRQykqE4T95QQyJJgUdr4QCiqqpcFVFz+z4/Wxzx2acV9d5
VEB+al7gl9nfcXqqA5gzW7jW9ZKuxKQUTumEsuMMhgNK8X9mOQbNntCLrkxDFEls
rSuEujUA+gBlv1kEVz8S2l4IVg4mpTzCLlMdzQwOWceef7Dxm7sXeHqqewVzXvAG
DUpMsO74QL5TD/dO/Z2k9YgcNHlpjc5agz98ueYHK+2OvqEV5zzpYP7yF25iB/Gr
Ago8q2Yx3L6P6lksVDlLNC/n4Nvgnz1AF5qmloHSSD+swYLy8jF+3APC5rnF50rk
cYPQca1y309FbP/J2c2DNmiMyzCgFfnvm1KVqH39c8Bz1PdCBA5mEpRZTS/OL3VX
RdiaMYBh2V93kYtUyRNpvQxcoS3SHhfJNfoz938Q7yRWdPnhpzH7fMN49J4pQY7O
c652GjokfxqH7QUtOpzfzeNB5cyjqCUXy2MeIHEaqcFjEpRcrdOQ4gSQSYwEv2jP
mlA57w2bVpK0reLoMP+KNbBXs83HD7x4zKtPOaKnCgYjbLpHJ0j6MaxvbJ220u0K
x9j1tvoqYGqlvALnl+8ni3gmIOARc5yw0jDI70jcka8A2YZcu2GWPLXEvGbqXpIm
PElXRyMPNnnQ7FjoHUgbBjfRMIy14xalt8daTYz9/rdJdjsL652FoK4q14Q/AR9j
UlVtTLDjOuTb/uAmThOuPV8MkUjVzu8fPL2K2Edx8/EkL3njotIBYn1NGzcbxrfF
x/7t6IjvijP4kO1hBw33gJlb0qnFb2LWKlG+qi4LcjiF9oc91YA97moanGZu32nY
hTW1cotYh8a1UEDHnfqTDjLC3+0bvXDaADeuPXZORxyOx0V9cdvuvc4yb7sHhspE
+7vuH5u95jwBlgbyhGdm0jVXkirkaXUoI5by6LVJcIXFmKRcGtVHt3kC8CvQ+wwg
SYHcRukvS8WgW3Yy3ib6O4dUwdEQgz6zWJ9FYsiCvkyZMEy+FJTpXCxZFrcuf7l7
VSKkoycK7BKoN2wFXKAM2aUspk5cCatAotNYLSzKXbvq89cF9mffjW0lpFUC1tOj
ojzFFK1q3xGm+KzvdmGdXODfcB5fV/dL+eANRdMII3gxY0A/m/x/MCDIR6epPI8F
3JhOkSdR/H+RHsuM4lsORGDH9aaLEO6vzwUOe7BpOuQWK/Emb1B7P3AixxXQOmc0
xVvilhb7QL96Y3cVODzE+MQyy5PgY+irJyv6CN2ltfMVyhPBVTdjV6mt/vhcFuoY
d7yRqOZKiwY59hfho+OtqS4Zm+HfuW1FMgEfPzh1xS13SB5D3V1HTL/+0WF6A8cF
mOd6BY+v4rUiw8gY0oY45BuH+4k+SsC54tpWnhNLDauoH9qAW7Xjekdf+rxMVdgi
IxctK9EO+U+rzBBN0AyPzyr07c8i3qW3YABotX4HqRMb/XtyplCX97ioKXitD4Hh
7rBRbGCy1G5fYLgWlel1hkhlGbcz4HMJPBmsCxH9eRkAAEgOxvvAN2wK+sCXglA8
7XulD7HAOMZoZmDbI56joRMST2ArXHFi3JnOWORL0H3ZUtkW+AHEai7UE8ca70FN
YS6jAuL8ikySnGEN8rjWZyBO76geVwo8fuW6wbsrQdHZvAILx0diuZhO81JzKKdx
K50W+JYgKzx3Qa/pkQV/cg8tEPP+szYklmTxEF60uUQkeSfD5xbhddOQL8aKkA2J
vcWbmeyRt0dWPM5qpOisGPcgepNmq8MmTGD7z9NZ1zDz5Vg1sR+Ww/qRIRlFJvBQ
AegbMhBfjGgRPcjlwrqzZp2RvN3lBOoDwn0lUNrwvOTysUqVBbmAVhy8b4P6LIgY
Ov1wL3mNY1jtZpBtZMtnpLMNCxE9vVipD3il2jt/HcimwzrC6wyDfquASdl3Geq4
SIGwXBybkHOz2hEfq/BWXQsrO7e5ZG3IklUrDYyHHk91naQIQlAIimHc2GSLE6XS
sjFKFdlih0XEsA3TDAR7Fp0Hu7oweEAU0Pe75lOBPl7IF5yzKuxzdhCBQBwZIPxy
CyXCOgXH5AwSZ5v5uTf2YGYe5OwgQttvkjQLdOLvbEZOLpoQkxbCFszOlCW9Ws5n
Qs5ZW3UJdcPVDchTp+qtZBNymVNHMLki0TlreoI69cnjyIDlRq+1cpfd0tzceKTs
UO998tndq0Mdxf5BxlK7dCO7yLUHnySMCC6DmoCHryB4psZG1Xl9fuGfoEg5zp1G
X7jOk/bx2O2+x1QZggt/a7taiYPLfoPu8QH2Ul7xDQBWXScvqXMKol+JF4OzlgKV
FYlLocFl0I2iPBBBMn+e50YxFuA+zH7VdJsYzDAC5bmPlSd9b+0TsYjtRsZpMxzM
WTOISciln92CFtM4ien/Jp/j/FDhl+4OOkaqNayvYl6/zJjuKS/kUBUgzdzw5GrT
r3D3Ppdffz9u/An5nxxUFl3eJ9qCqPST8SjQZn+trz9egnf1IeXptXgi9/xmt8qn
gsevd8tQWRvo45u+eMyL6YZ3s8NCtrY6a6yfLa1+SVEmPyz/urgbp153a0W+ngbM
RQOtsByYPgIgisC/xfTOfvQM//Xi2a3jTYqiYrJ75lb0f7YGRm1Zsdi2d1dHao0f
PAanrarLNZn8cUryjpDq9Al5cvJaJIigK1irKNPvezMTkeayiF6eIgRkKkwDy94O
kn4WwAbKr3Th2Ie+gC//5D8lDTK8klNoi1xMWYKlhm0kj0/7SlLUNe3XTV1x/iM0
3hDzPJKUcNw7trrjZLEowgXwpuQbOYbDr2GeUOFMWhvSTp1cQkqXKACawsFuymnl
VhHHhgPEVhHBZ8podEU8elfNT4qPmXGZ6NFTz+unHkIoleifpyq4/hR7L9EjJvMo
xggXXtTcw4/myXy2VYmGT1Ypo+FyfGON2meSvKB9hvaUoBpPmVAr9w/F6vjVhblo
HzWa1BT1iX+yuOuNHWmB1fLIPrTGBbIpgm7bpcDJBXOI1GfbwzmTKy3jN3zRecj0
DJfk/Udct841zF3lHZHqXY17UY4EypTPdXYGV6eSflONNZeCe2CEmjCMU6wAXOe5
JwkwFAB9fthIy4thQ+VTZHlIf5SoapXtU8V6/FZ16pVmMOA/zC/T/BH74ApuVoWM
0Yh2TTpjxLXhK8dSwDBXoPGFdQZJpJ+B4BrkNpq2B5OaD2YmRI800UICYuc4uvfb
WDtkWLTwBfk8cwmSRG6fgZXGZi6L6BVpCtsXeXdGWR6IESnt+LX6Bw5LslasKCs7
miw4kpm1HY2ZHSVLWDqQ9lhzF1eeXni+dIXgl8uUDPAmql9nvtSQ3BeOeg8jzpU1
wb8HHP2SQP+s0UuhNJvQCW8ZE/lzmE3lAODGqf9CPSnfHvYt5kh7MC34RzWfwehm
teCd0XGDzHfHOBZbeu3wUmTT5t3E0Aq3dcqDm6A4jz81Xr/FLEMwWhZgiBcOMNKg
N7H6Xp0IBqUCf6J8odEhtJbbVE36b6AsBtYPUcX6GnFnh83PFk8wGDplwgmaaA5B
U9Pntcosfop13ekO8XN5nbBFtdrFojV9+XWdlps1lMjMTzwtOqLuFOqpOJyL4SFP
0ABxou706kwTWaOinB2t7Py/Uhmq1OPesS64FmEznojz+wC7tjfbRglKurEPntsp
TTICcc/gzdbeAci2ZnweMHR7RexsK07wqxX9/CTwj/2B07BuztaURPkdK1Bov49i
fSf/bttqw8m4WWngZ6DI7Y9wkkOaQWL60+fPxUz5yiNqb2icwT/Y9TkWn9axQ9SD
/XklUEPCCkBbFeIAerFeB/B+GKJmrwjWawA3F5kNxTCn5onFZxWjqQmfDH4rBiYU
BunXpNTLE0xksoidYftFicEqIYiUXwjO9tiip+2yqytzzUfR+D24BSSeL0wiYYuh
eNmKQlnP2OLugXKP0Dm5SYTWQhop8xO53VLxST2SUOillpSmFgXxbYowBasIyXG8
/Dzeasu6TiRjBJJ3GG5QSmfMsJkEscJXwtJQ+Q8nhiXz06zvNJXVTf6svtp8G5Wj
OCufOAY2r0FeS3W/9Nixct/AJn4lzc+U6wDc9bcQSpZVzZ7XfX6u1MjG+o5kXAcO
YTYYdE9blFTbM6yYSbBo66gA5ZKUxF8ZD1I8+UaUxVkyXfWQvhkXVyKsm/QeN28M
QX37MLhpCkZLCg+GFkreaFg3RA/Dk1nb0tB8pfjijHaGQHu0xI6HLBjiAg8nRq3O
X7xLuxgws7QNfy33Xkwq9gI3QmLehWcg0noqc+8P3MkxmnG86bYI3jPNp6j/bhor
HH5zkePhteamQs61UHFXFzMLsOHctWqRPdmsUrACHNHWjTwVdR3a3fGpwmEtOitg
Ak+5oFHLlFlRKuMjVCxIgOZqKQ9n4/GZWomRSf9Saf5DtbSEaLdtjOaNmjW3dg+s
NDuXwM+5PpuNmTlmuH/HSsXYv7OZqcbqwn+I1TJad83tECGJWwaqkPlM/79UzApW
BkLpaxjsoSyVgNUz6Gj8O0DOyxnHmyav6MUNStSKy3DJM+s+oYXSCn2IZibc7UG+
k0odhYx9cJAORGqDbp//WzUzPW/38OketxvTDUo5ZScc9lbBQ1Yj8UH2XcmvAYx0
Xik1sRJeGiTVfQBzffg+p4lNpia161j8Z4wGNRkTMFwOwydVKyZwv/TH87QuyK8L
tpFL6221P9842Tg3ZYJs35K/20HpeW9NnGJvWIZ6NiWcupr3O8XcuVSPHPLQTPbq
HOZ6dEcmUoLCvcsYvB4EmbXeknkRMSTXYGMPs4logwxwG5rnKfZkNappinmcI2tP
sZU/EdZQIRNqreob15wLrECyRt3EGA5Zfn9jGnGgpdvFXvxyWHCTgKzB4JSvsvHO
1x3EOCtQ+uC3F4awI84K6jdtuxzP30L+p89LvfP9A1i5i7pmQbxT4phhx+9DfIUY
69zMISMMga6MdPmGH/TBYgIaKtcQN0BVpXTdtq9KzC8x8lIoLUYJLkS9884kvWm+
zpzDOXfsxtIA6ujtwPIAcNh3HTj5sqmHlHI0t54LSOnc8jDQ8GnR85YBQVGfVnWC
7k9GBDoadIvD+XUu0XmvqAQMYCUf1LlVLe86ojcXf09T9B75v0qUo9neni+pB4TC
r/kH6JExa5dk5SvqLDKw62Vp/LDuRPSl3U4oIIaZzVZXu1mH4X5vfTLnm5SqCLl8
Vw2DjDkdZXuNg/mtIheVi7pOzYlMAdWAS3azunR77i3rzUsKiFwE85IiWI56Gggi
oC9DRT6uSnfMXv+viEtUCvzC4r6RdhagxpwNfbcXYLcnOj0xObtLvlLHkrDw+ZU6
pHUE+mqsGQGydhnH1fIeMcf7GEPOutG3W+mswyQFyeiN4hLJTIVoFVEECko2L8qt
zHpGo5olbxtclCUOfKFOcwy7xTWuNjlF+yAdzpto8/yL1wyMBFBC7Sb+Q7GTEPWM
azUI/6LPm0sh5SlVU1DgEvuj1RXNQtswOlALMIOAnY6YhgDdez9kKn/WCAxJa27q
9SShT4anpZFmJXrHmVukuVeXBwpDPyURDlNmJf5kjiqbwrlfGdfN1ZOJo34hCFvz
+/r8Vd3q/hL9Sxo0riiPfbkuJxIDDdQ34kbexpGm4I8m+kxg2evS6380BrhXqTUD
0oVgNIpe2UeFtjSxANXFeDrI2wQWX2Zi0RZ9qVXjfPj5NNd0PNihV20LmqERsLAY
HwMCOWRbY0MiPCIncmeDV+H41zfSQB9AuxoIozlI1G7aEMVrxaASSgjcfsH3A11F
bdJAYv3sdrRKzn0VYMEjS7aMkeEW+W7IWGrjFD5GC3UwyAjzUgTkgYHJtfNLd1Zz
ym0C9xzZdlbbbdiXD4619ws2HVQb2Gn7xlnolN+5I02PvXqCvbePlHDdgez9QAsD
EYb0ncD2XAxFRDiIVEuaQlMrHHdRE6NvjYq6jvoyO8VVdfm3mAHnL2No79haVgip
KFHDnNK2XGlSGae2D2tefTRPHwhFREv2MKlkIPr1MyyZ8//t6ENE9dLxD4atTCTE
bNZF62Z9Tdsvi9vbfWgFF3dWP3BtsaUQWL7hLSmtUaBDQRSbl9dbr4e0TkbpTqHZ
XREFwbvkN55oFHrKuAVBR4CUsMU2vX3c5kpLb3RZB5TIzu+XtGAEErkijj/uXv0M
tMgR8JdXQtNF1dkZfQnr6PcXdVpxe5JihRKkArDoME8Qv02Zq41M+6Ujaej1f7HW
3pSGozC4nCC337dj4SM9iPPhmA0sn9rxhMK++eSpEsepHLK4lGlKxRboIGylFKeV
ExG0WqQi/6SIydrnYqnzlngdk5toHnWE9ZZNyEcTwfUMB6MvbpxV9V59/HMkjMGd
ABh3TE4v600CzcVm7Opv1LSDiPIdpaJh2jAqT6Zb+UI9cQa8fBqnbFCHQTZdO6z5
lIJb4mpuIN1tRu79woZcXPEHnFJwHVJOcgNYbTEC+U8eh+YolG/E4NzkxGLhznUE
0aAyQid5ct9pbP7zLmishpIMAle5dhQQ+bB9VufdkZJJqGOaMM3xwFjWTYEe1IyP
Rl5y7Qs0fcTgJtspWwd5IqBldWfoJiBNwdrJ4I14DkRoUucTKfi67ZewAV2AjacK
wdnYzFDBZbenZaaq6AVTAdnZ+fP4qDHSJ+siqDlms5owwR1HZXVGlKzdRp1DfhFM
08kloGCkbKQMUo4c7ruzwCO6EnkffXesq5cfgFgd9xvuuP+qdtr1+DqPWbkrPWVn
SWOYrLmzM6eQjIg2LJiK538st0kRpoKeP0ipk+2qxc2Gv0wg3vXf9rKZ3R+zpRNb
uUhqqRsOolgikwTiue3oVEl4HvLhc8g2/a9f4gpNAQW61J0GkxQE4agEZTGTLBP7
/n0hcUBK39AifVPA2O0UCGIsITiKUfoI2GCaNZCThP8Ra/Aib2sqA0K13rPfjp+u
dGwoiiZhiY6J7Gj8KPzCmQqgfEbw7KFnjKQGdJRE1JyZ6HA/4rCpuxE+l9IRfSrG
1O9RHVaBjT1VZBG2x/P2xjIhc5xFDfz+B/+a7865SQSbJSAmdd5xpC0o3VR078K9
3O1FCt5L9tFE0b9rTGg0nrK4yKg8MWrroy3AA/bWWZln21h5QWkdgJQJiA6jmKCl
Ezr81Qkl+eGioppOmzq8MEknOfnIDFMEkX0Z5J0gKJC1nGOfHtEgq35BR3VIAgpm
xpiHyIXgycWfyZ7M50yZVtWm8+cb3KEPW9uPi94DfKEAIwzX+TunHvdDjfvDJM7c
ZIX/5BIGWJjS+r+lBTgmtMN34nSYstuVOEvqdAyRC55xjtZdHmVy4sjA+LaJ7DKZ
hmTYr/TYooBVFFJekFpoESsbC2h0QqufssFwG4V8FIuVbWgqRcs97VcNfAd23I6q
UQaYsxtvbTbTTtX71/buzgY4Q1GpvxHWN0PzZKv3oHHvzjMj+1wGdjRuMcrKghy4
mKJ/R/B08S51K4OC2JP4TfWeH/k2HkLGq/smZcn6rjnN1JaP8tq/iVohKooV41VT
LNC4Z2FoopA/uHeU0UWGAl2SDY0EjHQRoFeU1OzjhHXGLYKCLubhlbGUKH5muj3d
hLyttUOZMMlshwhzqymZQjLGB+FiWmVOmAIBxMFSn3EPwNTXJeL9lCU3fmKe8l52
/ddxuEbhkGLItfbdDEmVZ9kKDkUcaeu4tZRxEDxwp3vkEqZwbixLGt7gdHhsFlMC
4Ccg8LXN6Xl8IUNDpuO4G7HHFQjyk1AUvIhUPA1X0oQuEAyXqE1Ml3vpFCEzmyLW
ba5p+X2/9quXOXQPntooqksucRivSFIzCBB+gDeEQwzHMVsmbiNpMS4TLx+qoV9e
6SmIgVIRB67IQpSFY8ccG1CNyNd240zqAZt6gz43yc1SJrJx5QvZOj0c0aqHJJxZ
Ip9knnj4DhG/I7c/7AtvBPV5lcb7UlHiw5ycBAM4j497559+z8Xm2K57Hpx7DvVT
6z4I6FqowhRxU8Z+Qt8FRdo7cgN/3I6Yamh+bsW5UjeBPIQuXMABI8SEA4byltxf
u4EXQXhltqce0GONQxe4EXuGSnIYa0yQ7PmiAmf/SpVoGJ10AOvS8/bUKP89kHbt
Vg7gj6EsrAOuw+TqMPDzHQmwoh7bn7Ae64oIgFeSB3OkLxKDMB/Dugf2PxdHS5vE
wEr7SsxCxD8FM+7IbrtxDgtb+Eykpq9dbnfjXVs8A8DGSH1VE2TL0ist9uwxLHFy
impM77Rdc33MX3EiDQxpAAumGngAOnAPbGHPC14gqGiqeBgIsal3Y176A9TY1MQs
2DnhCH/mUrm0qoqfpWEp4YTK2Vm2jHu3r35NPuWVHAzQGWfTvTborv5phNxsX+zW
mp1AjOiJvC8wQkt5tjFH3VD6v01tbhWEHm+e7eAAviXJjtQpYTW4unCIgfj/53nQ
njU/outu4Ngc/D7y1F8KHY4NNcVKuX6OiKRxmGBYesTEnsl+54UAPm41YdG8weLD
D+cQc6YXxKQSCzni6c85XTFi7gPS0BMvroQVMkp6gfK2hBah6nKXkh1WPVWW+xgQ
tITwLQ9UOxra69hcPSEoOZVE+HxjufAgcRCfFkB2Yzdpetyt2K05gRgcn8tOYC9T
P9La58pdZDREgv9aET5i2+LIodcDH3Ts7CBs+By0mP7JS1tOz2+XbrzOCof6oUfp
WqWZ4iGddnPV7fEz3cVnOm5HBt/90gQc9aMcUMsIVLoko1lcWbrsYLJgRgRVzoAD
jIsAUOF2+XxUCJwaNwZbg3zkdysGNv7QZtcMyFHwBgQsdDJmujLeWrhD4PGbQusD
+X1WN5ls1sEoLiHbky1OPO4cTHjTSyU061rt+K5om/rSn7fMGw/oIRvVCiguukdu
hX4+kfM5aEUVdo2T73f2BVe2enBtXfUZtxsJizadCLnLGhh1IH4LSFOTd5O6TeTo
bOvDOGiErPbGhM5G9RSUmmPXQPpEm460Qa0Ov6n8gtM0PsSRS6nYLCopOmoZF+2O
ktx9CL5HKAeVeutRypc7LsUX3XYFBStaNGxWePVGn8vtB9mO+ZGs9Jy0Hmy1TPWo
RGIBMDN2J0+mFl+gfM5xDwvUAI9f3hiXHtfR0tZ+2zOlo/OmUgjWlOUr/SR48sRi
CeX2r5od0Tuk6U0oobotCeQzEifeCVXcvj1mQ8fRm9GysP8McW60acDqGAkakFBl
EtxbKB14/UzYL2sVexnH8MNi8l+8PemKYGxSugb94u5krzkHgevIw3T6KRKq1SQd
OXHEv4AVsYzuG/qXlM+Iyh2cRlqgXhIX31Fbag2PR/YOsRsZhvXw4huXByMhumee
SQEmIOig1TPYKimvrbuPTFOSt/YlVuPbkITiL0Wfa+yYO82703CtTp9l4CgKkyJT
k5Mi6KuqXBzBPrIN4FtCryYXutd5SBwZadMBtkj5m4J/mrGQBG42oyqULjNiahHt
K+j6lJ/PN2OtYcSb/7gPMGnpAbG7NJ+peVTHPKP0PedLhFi7ZtphZQqNKUDbMFtP
Afa1U3RAfSO8Gu6GEp9KHE0SrQh1ZMVxYFUN1jimt1dlX8hsXB/LMhtVj2fge8Js
+8OmvZ+re5UeMkbpNJISvlCgBCvNEWnULBkHYZpXhv+yLPnf29Dis+FK5hr+ZBLb
FoDQEb58WQpPREzHVBHiIH1nInkoMz9SczSvwA3I3PzTJAXLBwriJwz3jGNIWp55
jsUwSSG6zDtwWn+StQxhfaZT+/UkJj86WOnDxHyT0trGxavTtit/SrjrtvdCX+Mx
Kx8gk7Mu6qbDVh03J4+p9Yu/4Uc3mgFhIuYR/3slPi8bBEcgSovHBOxWuy4R5GPd
ROQEQ5LMZWq3ljqEd7a1LpCbV5WuUDss1lMGi3rLDXbAgfmyfz74ohD/oZwCiiNf
jor4kiEJl1vXGlvLuY7JFBfP3lecU4KsFk0PagMfxJbVWH0nsWrWtZOBmvNEcMeW
nDeUkuGpWWEwj5aOCsBOYmST8PPKp3CHyhp8feid7o1/kZKyyeGeVQUGekyWGsXS
dbeg9Qto+eh63ZFjfSvm0HbtID9kIrs+CGblpZJiEurajoHGN1wgo8zygm8FreQa
PWClSxR2uMCnvOvPmOnb+aeiLho4utQzVQUsAtsSU5XMurnfWiD4LudkXspk/FBr
Nb3w8JV76SBUEyq/kjxyolonGAbRpr/BknZwrbmu7jyMyGrwihSvO2MBv5+F0lUO
tLM791Q5oeahUu9TlP4Jt9WxWBu2PtfoypkerqGqbMM5gTayyif2VgLb9Z33L9ny
Mq4MqxqiKSkXwNGCTtKfaC3lEb4xoHaxWLIIzUgX8nFB9Dt+DaBqns488yblMCeW
p4tg7ixgXc0LmV/ONlxyZ5L9wENHxR4HUvxAYQC9qBLiY6f6oXI7tplVaei6E3Xj
o/EqRkElhFEQ/fAAwdPq/zvF0amt8L36yeCjt5skVLWYZ8P7mYF5zp/cmMHnLYur
zAGWJ601ntCX0xgm0ds9elRnr4LSsU05Zf4Ris/iYJH3HiHrx0hTr8zyiwX7blV2
Ksu9qwECJvBTzQqqUGjSSGYdjqyBcrDYRjdOMdvDK/B9hOjMu+RyAIkT1yIO1aFJ
kTR1m1Gp/mCIqrTIiOX0FG45AwQZEhBqDBjZgn7OAqKDYjPYBcb705bV0YAggGOy
f3Pe59/Eg8NnW7iUtvMBK1cCE0udgEv6eZ9onRytPhyMNlG+JJICTx5P4R6iGxcL
gDwNjJaC1eLTn0ae5/s2+i+N1qhl+lXABKKWIGtsvsU9Y2q99BwSpGL3HZaUiN2Q
HyG4S8ODFp7aB2tNPSq+EdHzTbqHnkjfftVSTCMzg72+LOSkF86rUrKzU6VNsDJU
nmTDclUT/QkK3G4DplS5RnkBposIaUA5bsz0HzJqn+7ssOitb1zLHc1pIigMxL2U
3l7p/RVFVNftBkl7iu4pbBQd9w3O5JV7Ut+Qcqh/qjTLGyhbp6nZZv3wu3V2RSDQ
TwnkBXfRkCSvbj5PXDvB4ft3Ge3ykxXlummVp+G6s7Sb0cZmlhPkuNUxXz2oUpwH
Zs36EGBx0+i0P9LI4EkGrS4bwtAkWUqKbzjeTS+mDMIliO2fVJXgRZimKoLZpe+w
YwUOp61M69tOsa1His97FZXkH5FehQzz499vetWcxcsI6P0a2LZHTzSQx+5XRswj
9Yd2f/8bEI7WsG7WYB65IakgVHOY0G68+8uXxW5wrmYRPpLi9D4QPQqkGVLED4d5
FAODbqlG6NaFGDa9LX9pxZyVCe0CIBp+0oRz1wXJeWVFI7WMCctT5u2gKp1d8kZH
VG+rJ5HW8z2ngzN3Xq2Aa7YzKm+JtLyVLR3z+i0e/9G2Tc84sqib3A82zARRWrq7
A/5B4t2ZTuVSaLZQTgkxCa2bjKIyr+0LK1fNqSA4i0gd8FPX4eRiQB19C+FlEfNE
Fcd8kQn9CpMHgF8xZzsr60FcJa4Ct3eNeRHkkIffkjg9Y1CXM3CmeSprmci5DABW
0XT64iMebExCEUo12Mxzfg1u2JGAc1BkwjERGFqcszP8FqihkLXMOoVfPai42/Fg
neScgfCeB2PJ0yhfFtSiRVnFWas90JJYvIALaCS+DMwD61gmkDTOv6aymGFUBb0Y
6NVWyLfLvRBGpyTIK0gYzlMe7bzTapue3U7vIrCXgfaS4K8fPHT9w14ktdCs3GWO
FTu3itLUF+nnfBumD9/3GWwgAykNgBI/glvTC3DxhjJj1/2lThhHGrppEm/JsB5U
jufnH2TS8WSp9TkM8GGdjBOsfJC23a3ePCkcRjRoRDqH46eDVEvrQGNAGtXBMLQk
6a3ggoXSR5Qvuz3ctO5q47zp7mAXcu5cQEsuWdiZh6ZOrp7vTlEOQ2S5SXhtw7T3
Ha9XsyTJUpZstaKEvJ/fD0K83GNIDvnf1Ntlgbv2ycZLKMn9sX4MUBwW9nzmazvU
FAV9UvB2QXgOR00S2lN0EnG/6E7UtBjJ7nWRIwoQn/89NEeucrI+ZlWTvfh9bPS1
IfFz4WmS/m5v2HAZ7kxEXvOGlKFlM/6zIaO/aX4XXFKoxxmFYEONnt2G7eZj3Y87
fZUjsljy/XKV0YkpCvN88/x8oLI3a0KhNMEsjxowAqq4XDI7u2aCi4XdHi22xc7z
FWz8FWX53LbXVtCLSsMFV+UO2e8zVGx5UpXA6Qj8xaU+8NHEgGIhjwMpGwsET/4C
ZUoX66R9AkhMxv4Yww7N734qIU3Fp0IrJC/23hru1wgkdVn3B7LuSoTJJBhBd2f8
kEjfk/orMkoDt/wGkndkEN3LGRCFTwmLst8IefJBYRwrBDXaHQc2Tn051J5xCE6x
dx/WJxOWgEBwScBUXPeocDxrQ4BdgYGwyEXGpL3Hf8/J7bCr3Czj8vbkW9Dd6Km8
jLIV69sIYhJbEdoYNqrmTWZKMD5uJngELFYEdqGsxtLHeYfgLFiv/HIM0Qqg7Jui
ptq6LmFwJEXAwVkUcbj0d+nKM2UvRTTv/Da01psUElbKeyLIRIwP7iht1erjGAoC
nhBMLQwtujjVgYqM6clck99Gz7KBH/bdt4dDY8Wb2bsL/GIC8PkZQQE2LaCgoLhK
3w4ualfygby1AAJJ7qgO3AAhZWEDer7IAfG1rflI3x2ahfvKr0UOcq113iurKNvu
LQgsWUbpYa5FTNY7vaei63PaJDbVwK5EhfqmUmQPgL9Q7jKVjd//PJxP+xagGF7x
2uNXNR4SfMXL9ky3Nd8eUeU6dXC5x2gN5/fbbqKxqcgwFrgIa5F3EW8zUR9ve9ZW
08r7XOpO8l916o3gsRYAOIY9PHZX4356KHTA6XwHQr+fhbFz+c7FZJowUuZJ4kOu
GxiTQd0hf8Le0epaTL062/qEMGgrIWNLgIOmj7LvBwCrzz2/cXMojatqL3oIj/WP
lL0Q6ZC6VIofbkwuF4N0nV0ooHjlR3SXyvT3fbJDlN70n7PkQprMmkSh7fAyoIbK
eknEYEVlZfct84OtA12YyyaOdfGuU8sWWPSKSiKbHXIRplMgGcrEBwsIQX8ahWZC
f3D35NimRrUs2xBzHS6lKpPmckjVfbzl4e7ur5/s5W2T3IZb2XLP1v9zBgCcj7tU
gJ87mp1aaHeGZEYxvRLmszLwvyp+nOCZYGMtBibc+rR8eOmXjgCa8Hp+N2tc4rqv
1IDnf5cxgfAebSMT0XDuoG0X99eomxyBXI/x6mlBw2fUki+2lpHOjS68VcDJmg7n
XqYNIIJR+21+T1vTkNp4flhetyhDPGHJ53whxEyOODMol6vTx7KA2/8ag9N0IguW
ZAJwQbcjsvKCa/zOQBu/Nh0whsF7Sx13vENzNzEtsrUedS2wj7bwb7K5Jesx7eLl
BWDcggI/7eo7PIkaa+ejV/q/0gT++ibgMseCiSHgjQOUMsEalK8TNV6TG90R/cO/
uQrYSyeASsTsc+3buV2NKejc/JBr3X9FJIul8BIb9la4/HidG2g5qXQKB5TaM8Av
Bf7WxmeNreRL9JtSPkkh0GKa17/SI6GixZwbgFnMi4lrmO1CQMalLpmyX+Y6D7oQ
+90itSISmsyHaEsJI7spEK8gL/Jnnhf7fi3sMvobkSi1T6zf0qGRTm4QZAZYC33q
2RyzgxSHmo6uhSFRIFhxGIxaoy1D/3UMx9L6MZKktTba1ICrd++SP0i48EerCleE
z/WeILsUj3Z/qxgw62/IphRnovGJguxv+2dO+vINdCsXMgunPmUS5/51QbbcsxBZ
BM2CE7b5Bka1/cUj2u+zlWGN6s58KNw1U2o4IKZYDcMzzV72cWgUxjA/w4VjlUGr
oruelZnwolN02atDuJE6717GzeJ5VTvrUMoF0Q9js+2WxO30VcsnCehZ5VXnWyEm
0OwRPHT+YUrnmIBQ+ORt11sceDbsdo8yNN4Q8STiaPgFsLirW7nCfp3ZQjvLNUqV
IdOaQSjLEsmfIo4MU/CsN+Ohpg7EBd5Q/y+jwtk4gJsB0YX0WJmoI14AAyGapIib
w4VbNsiNsXw6bkNwjVfZMXgq5V5ufMS5x7y2v8kHvJL1RBvzSi0Pgg0uNBOEaqLY
jkIfVh2nrTiZszL0aEOj1t/R3cHiCV9Q7L3QrkaE6HLngzA1QOZLLbu5ULkz0j5Y
S1lk/xV2hcAfc9OnyuKXY+a0KL3F540uUhONvK17mPf41BlJRxsFkSVrPljZF0P8
3JU0m19ssJNbLzRDBuxrVH6n2fRZjhG8KYTSx3+1itPO9i/teWQ7scN5CtKzlfQx
dODYtFddZD/1xvv4PB1+z/IGkvDsOLx6OMHxwG7pzdbPOLQFFNuxyUiaJGz5C8PE
hbvLn6MGyrjqCenaq5Xcq5tSnjRQHNiK30xmqKn9LqXXczhgLeeUK2xWiWASAKz/
G78d535AuGLIOcQi2eUhvR8uQIzw5nbPJljjBZekngWEKhJfLHxhtoCopYCfgsbj
ziWbAcffvdVelrLKhL4fBPJoDVNzOtUSZHRg3xLBHJTXo5yZU2taXIbeQvnL655K
CcD0xzo4BzOR68QE9MYql/n2MxHH+qk9ZNtSwTGdaOd1xRKUO8UyjjW3u9uyHbH3
jkveqznvlzGG2sysr2POP4nMY7mvvy2XyajbhQUgRUQuJKq4VPvqeJtClo9n4FAS
z2qX+fAVsSuy+Ug6uxiMcXoKXRkzyye4hg3f6DKGjqzZGQrDYoeGRL3SMB1GwvtP
OTwmsAtFWsomIITAwXVyYV4vnuV1Et2+m5Q2Wh1C7bz1+qPPXVZMUYYKvmuHycdW
ecQylOZPpcE2DOTlf91qdcybqyvSGOgYk1Wv+IEr8/6umhlpXzDU9bAe06kLfcOx
70yAnIEFS5NS8M5cwQ1KSIeDPAkiyTD++FNFkclUPM5i5+vYb0OC7xTuX4OqoOIV
j9Dugi/liJTmvoUe1FLWpVCIpNoo8gz+5KYv5qmrNpb3A01iPEnbhLQm+p9Pq3uY
3dHhoXb3XJ43N55RRVSmhYI21SuppLYtwPHNOyIrF9aUiyFM5vhaU9Y6aG3CDmS0
hYHTCJ1g7v+RcLQowDWe2T9pZ1Xs4bACC1JP1DIKxCyephcWAKWJyDGmesSYrtpK
XfV+SpnlBnAveHadIV9fuRAAG99Zb+Ne7dudl28Pgxd7s9AkdHx7BzvEj888hAJs
c/w8jvzF4nfmA9ydz06Pe5HIJ2ByclQSVlQxC16oCEpYFALSlneMg3I8soU+bBqJ
AFtHz7VZyOgmlpGs6wOX5W4n49GLFcpjBAeM6Hs/3KUKS0IXAtfGY5nA2DmX12c6
0i3xiJmMK6YmFPjJLavkC9U06w3duYR6DTXpHBAVxSriVIqyvsEpqVKH0jwLDr5s
D+DV9gIazs56+i1KeKal0ifAtrQqKWgjP4xL9jfXXJyZ4jYnR9qDXiJKJLEFnttw
oeF+ZpZVaJWZP1hm3stvL3GR66KPr1bqITBotq9IkUFQtQrS0fXLxGK4BY497oXh
5DTl0WV9kYkP00NYdhFXS0fwuwy/NrfdEYCSXBvOkrCR2FZxMSeFJ1f5VAUq/VT0
MNw9ToD35p9DS+QDfDVbgkBGjv9E702+guUvS0KzbjSmrUA2ZnzYPNDi6fRTHLfo
VmBA0a5A2bf0CYw0pzjMyKF038+0Ei118z9N65V+tHUFw9nSKxgD/y9u3YLzZtEy
1hF5VxKQ67XLXn9/tXhiUJR0298yHWXiwfPaKoFo2nScZPaQKJx/8moQpBb5RP5A
MZRNMxRWfNWy08v3bjdGV13s5y3eDsmkJmf79aHsANj/li2gsjA2a3pw3A6hINv1
wQVM4BQIgw9e+HrtG3W1ClCrG6d7vg48UFhsrmtxuxkXlWU3NrLAg4l0pQNSiJhg
hZLQrZmdwwNXf/ZWIvOFdfE5KTsdZAbmbCx4cA4xO8LdunWGYR1+zkjsR2c7aoYh
WX+ztf8Yd1lXURG+6+sfi7KSCq29LPFFfaafC0XaQ8ujr8mO3DDCeFbC8a98fNWF
aJoJ+OcmhZJZh9c67sEA7T92kk+3mWbxW9SLeogp8fKQ8ty7lnjRcqQAZxxEDGiN
NKYNoNN0Se8Kk5+pgn/sHEhrldntr5b3uzsPVEWlB6DduMOZUveOD7JYq6MUN0pP
zAwUbqiM4ixp4vvlWMF+s1NwWUfD4XJSJBavFk5EQYgjF2coBkvAHaZ0+UYTYHHT
4gVfflbtU8IT+Iosw3eeN0lJPOFUyB7vUFVRkqwvj8x6Weq8vDCOCG884D6BdGyI
v8TBo4QjTI1mQWqVKUhUMybnZTfd2ZSvmvB3jd9aqVJbda+3+tKvAK+bamz8lbBe
mVBVkachOmnXlYuzHakdVUU4hPe1kP5qR14MNGeGsMpDwbr+tBtOuJ/ii6g2TUv4
Ug5wJtu5i2FhfykAUqwRiosV7KhOaxOtxfGVFc9lvBrERF1BI3/fkZ3boY5LSyPy
glFpSqTnZh0EWj7hawHXQkqzPtXJj0Nx4YOJERH3RgsiZwaPdu1JWmQwCUtpeXLF
p+UE6iOgu14nkc4q0OdkmMyXsJE29VTmhai78rRoVOC08CqM1yd6GBhaD8DIUGcD
d/NorAl19XMZsPxNUk8+7TZuJUE08H/ebIKvuc5vto+FVXACw+/7ru0HLLHQ6VLn
BbDlWlDJkTZzq9Yha3SlgZ5wez5M1ZxJ19GwK9cRkRRTKd1wer445KW8+emrXKK1
S3I0GeqcZbpYN/AyrSWhm+5/KGMQ3CEll9bC/SDQ+SII7jvRCT2lL4EogLdUSisN
clWDAhg/LpRc/IPwUpZWoNA19UAGXwqhN8RJDs/PBHIZKHt7ImT1mIBYRefnPCxz
PtvxZyzavTUPkuQ/GBRfbpZSpVFGbAvCTluJuS+g1LIuQT+MptdIojZgOsgrZTTV
pcRWRYK9lWN16nOxhaTtYjJfN+5A6zbsdzHQanGRa/PZysMWS6T9E55Q4W2huJ9n
tVRWQjxbUtb+M1MmhXbrp26bbW6y9+iolzp2O6NkP+Pg2WZ7viW4M5eW2sic/QRU
9nH+fKv8wO9zIT5Qc+i1QM1d0tl0LWNH9IIOnEI3RkXReCmXflTCDFPzTbJKf7qV
9ZWWCLCyOBhFV5nWEogu1xxrszzAXpA1LVTbzPdSolNqVMj1QFnbrQwKj6BpuPXB
W0ywObZmIwBSMA0FWdZdD2zKgEeuXfNptfDZvG/BOLQI1j954T121sg1E5F9K/04
obRhUIISF60jGsplbThY9VDjC242poMxTSzfEIbEUz6X8UrhC2QgLXwKzNV0Gn+J
WRl3V2CqLeH977XHxNPFmxe5uV6BK4EqwcyAv9XxgnU96XE3/5CEyyuRvlby+Gi0
jOOlNmPtXgECuNa4xDyLtfaJwLtiNhqxTOfwXM/EINRGrGqZ6O/DG76tO/55qgHg
gfWAJWpBEAFtLY/k9rTmBdo1pr2aeAQzuvWns4IdRtrvuVHQT2fsBqW/iwiKNJnt
rqMgRrLi/lPdREYFM0wGf7OxwN7esGanf7k9+zaSnCvu26ydCH9F41uoF3UeXOXB
a0dkuhi8GBM7reGSVeIOpGWN3rLG0LneY46lKaC1VmrB6EwYTYE02D9KawWcHBFm
JFbAwUV31Qmwj5naxoPXvKvUhyEBQys1IZkMME22ImQ6HybPRT+VZKDuZf9EYVlW
SQSU8LVSqTWoo9lH2JeOyEgVL+nEEKOMxQihfniKnT/RnBDB3yxfF5YelQhY+UyC
PzXRHK4PcfAOwv8jAAv2nWzTC+TA69rqG8BcZ4P9v3CF+ksWPXVcC5p9iLLbQhk5
MbmHlSLnUSlruvC244J/X7aSgqJ6AKCkFbUbgZgeOplpprBNDB62wvwA/urd5moa
FM2wpK4CwuBUGSAC+aOoE0hhVUYDjZhCLkFxjApNDCbrPZyESukFnBuleO2FpUVS
L6Qxt/7ef6S+fk9KSuF8qMeNCqcclqTcBeK/9i9xm6LeFL6N8RRlb3LzWtW3NU1t
fsQ0H4ULkxBtxl55cr2GnpwkR74Gr15OLtvNMMDWsODaNGbdYz5niN6XmOX+VepU
tLvD4c60I/tWWpCVMIhQfGoYRoVC25k62vipCa2Kjrw0fCuZ8zq057JxGn1PU4l3
o6i4UpV3O+wQCtTKy0w5E0VTjHeEpHcuPgAML16DolGSj/RzVKdiWYmnG4Fo7dqY
52PW8umVC/yGoCVCiKBH/KdpEwZvawOr6vxsHKBv0pxMBoQ+Q7dzpx/i6nH0THAF
QMzq6dS1pgSkbb2EfCg4tLNnd+rTVXgYsxcgX2NeyP9FpgmKdqVyOAytJN+UVs2+
GlV7YHzI0YtQOxYQxVT0k7InEss9aWIZ8FnQBGBNIhqDtBhqI6Csq4sfzVPv9Wm0
icIfdA/qLXQls4xvzHgaNANdjrU6bTyDBEMycXYqyLPr5+JBIoBBXJyoHfdNkbCA
sBG9h5IJ5W5kya8rO/Ni9xlFleJ8A4YKnB28Mb+NXX9/hh2KbsFPYW/ECtpv9Lj4
767aeP7fUmIHjVSjP+DbvkUKTSkgzKoEUQLtJtYPiZtpOs0cMeULhD5P2UeiJBSE
yiE1LHilVE+LS/+sz4hoieADONJ5JMT5NC7srJswS0f7sXuqd/5aLXzg82zzQSvS
RABW64Ug3Ho7EVQ8jPTDwSxFZ+fD28nNZJufwZCf4OAeNk0wndqqgemMZ4o3+LlP
QeN+GrPDBNIC7AhoNfx6dKg12s9UgVuIaLZYlQLp2KJ1sx3MtLkbZbmAYWG3muYy
soURmUrCj9qZglAYAT6LPCpe3nIOAUsy4b1yfKyMva3PSEli3cSuSndPtoQYxlpr
5vLkqWqh2rM0clIeknwf8NDekMdOj3TlooYXtfVXKLZusUtOmeckpeuJR8t43zPs
P8dOr36PKbW/T5bfe8s8Jw94N2BF2Qqe8r+cfaeqHtXjUBvKLj/6kwEFksZGMX3t
UJNT6DW3U/Eg01oI09HiPdNT3YEGdhbTlg6GoFwC/S+g/HVB+L0lmjYQAR1bVTjh
eXFJRB2yJhLKuTmduqILdIee121ePbXHk2sD2uplRWqB0bXJijMz5qlB/NuNB18/
elyUSX6bIhgwHgCLXw6TmoocAko16ZNgB6HaCdjlL8NfJD2kCONlC4dryhNtYzib
52F0nmsRS/PFfgcTtghJ8p3He83Izit4RqDOZXis4x1Dv86SC0np2/m+7NTMBpGK
8dXHqhRVsdX7AtsROZVh6NsB7P291aZBRXHDawaXbdtc6QvLolZ+VXBH51SjIdtH
GpbkvVH/BNb5LpQ0CuqZT7XBuBJrefAV4T2ClDTRwukhJ0VHyvk+uUURpXFOZ4P8
qk7LDV0y3wo5V+eVxX3HFl+kj77uxou0n3suAgSoEqkCw+e2PFVUTOsrreLVZ+kf
SjGphcEDjG/26zoucq/i9nfJwbRU8irVPB1sZPoljD+Mb/2Bm2kmjm9UKw222W61
B5VPQj4GFa3xOdlOJqp6J+qxZ/W61s9hSHkhz7sQudg8AN/cJvGWi0uhQFgjTnRn
LdPdT2uor+58EL2xiOiJnTnF+fPYtnpaehNw8gK8Mi0Il43NQJmlHjMq5xLvHySN
FWAIf82O/G9CmRP9Lj2P2CatpXh9e8sVcCQUWAFYtDavccv3ycUVOjVN38Gk+gQT
qjP5kSJky9FTHt1MoWACD2VnxhzJHpDT28GHeTmg+PCIfDJNEaGPDTfHlRDHG2hH
BcR9LUU+nQDozaZLmvLGXRb+h1lhCW5nMF1GHg/Wsfozb2jNZJdw3ChQDdAEB2sq
uZWUA80wPz6UEPsgmlAs7bzIAwCig84ZXCpNEqtNlzQfafq6M4AAeJDZH5SBWKli
l1xROTap9XonNMTPpNooJOcBKfEFPDJpcF0c4fZkQjqqQ6VmayiN81MeFbGQbTx5
VucDL/fTt6scGSRugT2gTuYiKXoVTQL8Cgrz5blWNCWQeZDKodaI5Nzl7s8smxQH
TCM10Dc6Bv61FO9o4xCvT5cOFV1KkbrMqZxubm+WDRocWM6blyJ0kg7JLlkoMr15
rjBnEHVk/y6FNMTayzoaueTHw9papPyqHOY5S2JIYzBpTQHXnqExj5kwCJPXO+MZ
Mx3mi6Oe6s00ZkT82HDIbW+VFWPYSsFGUJh9erJFDTF2sEIqrVlXUhDHeK/3tQQj
TePISgvVeVcoNeBU/4VYJngnyVNrH2NeJseB7vtz4F4R2qsrfYTLCVaVoUupYCuP
qKYVGJQUWwV4IU2v+NymIT2vzGLk+TOSUidMwv/uEPwMUSAlHnpMBtLkVz/lQxXc
ZR1RlUG5kpYx04rlne3mfKXLqYdTyqm2om+UNHDzdflKnQ2kJdQuYu1ztBU0pXqd
8lLUKmLM81fmEMfovR2Qo9IOcWURGwSZXFxBVSeygPqx9Le1ODHqrHUoU2e1dZVs
X1oBd3RiEuiUQLewlCOod21t4V0WzqIlEIv2Db2H2hEX1sgbTVIL6fdDmY9uG1z0
kBDWXPES2nfVbVg3NUu53sFTxoTPB3ma/QiokFVXqxNBmYL39CF6BAgc/Bg6vWY2
vThBOBWV0tKt7jnpKsS92H7cqa+3vHhvyDgvY9ySOYxMy3SHsPlFpJmCF4nZ2h8k
Z+2q7gY3AubueXs9x+krsLs5wEQysilYFdcl193dF9M7SFiLpZEzN4+rvP6+grUB
6WHe+HU/Fm7ZJGuwWhjJGKguNqQgfocGpDCMLskELxbaoX98AD3qiqh0z1ntq00Y
Bpq1ulcEyyuPwUWGRzMLRJcrrdB9+f5MJdTdrkLr8ps=
`pragma protect end_protected
