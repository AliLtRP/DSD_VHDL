// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A4y8aDFR2k2v+few2qTwPVxBrhxlxsdBrOccfEScGzOj0snqdLPk1llES/F0xQYR
k8syNx2daZI+4ppf+cJS0nlK6R8F8n3sxJLO36RyuYwQm5yVORHoH5TZ6ygF62uL
EHEQD+Xb1I4lMbkWj6JFVV/sldd1d/0Bs001+l8V5zk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6416)
tn9Cjl/t/JeuaK8dAd2kCOnOREGBOE9nE//pvnzCr+s5aXDkslBSDQq5tflVBTw6
OqEqe2b713jW21iCN4tCh6cXZ0shHBZzLYVbxKK7jvbZTbYe3clfgJyq5mi5w4rq
6ZqLSEjqXG55ntsiJ1zDGY+zfKji2WGx0MsFP4+CHZbcOalfyUNUa6g1qbm7Ec89
4jT9Ad07ZbECD2IOB2bx5o0qYfNbW0mydCrp8Nj7aqeeJhJPZFDF38xNtKGlyeJ7
Hofj7XnEqiq1jg7xNXA6234auPDfBV0g8iKMQMHQD+Jr55LnQotYxAWq6RmCHHbR
QlbXktykThMx8ehKkFuYAMPp5tsUlqdpIhF7jvAwdlaRjSRWGxgPU3whI9h9k0Bv
D6FDJWeZZk5QUH1io0wetEwCbccr+kAwigenrAoWNE7LRCVZ+iQoMBhDEEml4HOd
MuvexiqH9dYvnu5NBX/6t7lKVGSgMOrNAJYqXCr2JKAFwZ3rapV0+ChzJyTmntea
Guo1t6ytg5ZhrwSfTcV+GdBtw1Xs8EAmOA42Zhf4OVzBp9Q2yrKohHYU7IgDBYXx
MJDdhOkemkpVNcrcDcwlNUHSIJPZ3PqI87bT0LYVKrlIYdv4HVMuT2UUX3sG9GMY
oR7iWwtRlW9yRO9thbUSCkS2/dJQgXqI9aNX1ChJ87A+YXUaVp1swe53XNeaF2lG
e1cX32mWtepZwIWxdkszSNU7OimIsrV2mCZBRKaxDptu2OjDQuAlcCA9Qf+4UY+O
kl/A+8+0wyIfcNjubGLdQHYiw5YR1rIxhevy3wuUZlI1rCbiaJ5bvDfe+JtJ8o8g
nte8D/3pmzBZMDVmIyMDpr+hA0v+k4gvHBSJKkE7xh64PMtM+a/vUt2QEpyW5AsC
uMUWocVyUWpwUhUFmD0Zhgur2HxfOMb6XRhM3nWGFd6o4Oobg7XtXR01Ai/tmzFo
dlGSgAgVO6eis01KIFaUOB94Odz9pTyuw3rCpIjmZn4ejT+Cr1On2GHB6dKgZGuv
dpoL6FpurD0utI6IbEY8rjMouvETTdICEy+iLKPQCVJW/dr+SkWv8raJbPuRL2Hc
vzmB4q2KFOd1eK1WkDPNQ8GddIOqSIM9E3ZH9PMGQE4TF461M5Vxs/KkLsRm20ho
M6LkrPA5jWMXdHcJT7NESNlApatu6DbLFhX9HYHOlLtLBns5lEU4mY6uIvHlkH2X
hFtuebt5cKRKGs/UoU5en3yWfFqh4S7FhQyoG+wqSsBVKj5rvSOWxXAU6V33Gqlg
dNi/sdiTkU9G9aHlVsmwIYxZjsz9x0qydZmzk62UEW4WT1PiKdfdcU/RkzDPJvLw
mW94LE53tGkT0cwyGmxbJm1xzRakbmU44pgtMM6yvZ/ooOYtE0M8y9YsnLti9a/7
QDgDExgBsMNj5xq6fyhuobqVKp+X8tvGq9WxjyLUzg3xKI3LnvT5eN7e86/L2lfe
BcdYgkGPp+qIlAaRyJdrihSF9ToXI3UOsl2GgXyT1qNlX9jlOpHY2lmf26kpAkuJ
yO+TT7btaz3KPcobJPEy1blAijUwPv0MasZXK+hj36fruwl2whYalBQVoLzNgpnP
3e2Fqjw0odzfSalWS2UcJbIar6cnT8hwbp5E0/BXEkTr3Jc3q/2hewJQQS54M2AV
LO47RbUSynrtVQRJaLxnUBxF71ow9brGJ1b0MKU/wHyK3vlkGRq+ANQEvb0TeE8G
C1+Irjioi/RpRPNSwVTmwkv+HQubyREKeMjvG+A7ubk4qeCGOpAigU3O/bJhAfoL
rPHgxTc2lB/26POjj+vlEwPMYETLSYe7o9A91HenSIwq71DwxiLKPsTitIGaRnIE
u8/kjxxiOdQ4THiUE7L4qBwUbDA5igEByA3Xfz25foPlxokILmYFjKuD6HUwATlf
YMLoOqLrxJSob8AVDggfdwg6n4fJGDx3UcpjDZEB1o3ZdQcZuVih98I/a5DbBfIZ
raTYdMqZlc4N31BkvqccesO0NbBvEBYYh/nOLMo4L9n7WIwEFLoz3e/+p3Aw4yOb
FO5a4QYpR38L2MGCJkgj71CjwOzMBvQsziKtXk87VaaTUZu8L6iDp1CAs/u3oqmt
1mNRPTtSob5mmk6jWaksnzXw+jXfinttds9nxXrLZUMA/ExvA5lcQiAXUZ0J6Pyy
Iy2LQd6AqdnTPNa2J4d4lfY7/P5myLtaL7diwaT/q1SsFrE8DKmCYok+7q/WCO15
NzInbz9UMSaLcj8tAXcJnLv//Kjjnuje8rQsk/v1Nyvg8Sa8fpPkWmqZw/l/S8TZ
mQf8r86+ht9ScaU/AwmxhQvArZbnVNFYufONYJ1sfq9pzEW4dPophKcb0/vbc6Jh
i0tFda00RdaOwREb3o8s3AeeauatOY318opLS/vwwgqNi9k3j0eBrxtpThw2WSLl
+34psRW4clyEdKdgNZyEvfyKF/WA6oEQEH6xZUDkHkKTZhqzrEC5KIMCQWO8bxuu
3ErlJIF9lrVNa5NBAovu32inuYy/HMyyNRgAVHVHITOWR0B7VWJq0K1W0tfYur++
kQLy4YJuFzMu+Trgtdd0/kLkLJflA+2d6He78Pb/iEMzu4VSaBJZY8jLKj3AxBy4
3XGJADhiXgqQiIj/ork4hGFn6u5hbqb7dgyKun7daGgYcQCvb4E7TFpa2z6khkRv
xZlolQ6Y42/hMOOk66xt4wRldavrrA2QQjxGrvD1RuZepT+t14qHvwZ2vhTs42EQ
2ZOw9O+Ogu1D65XLrweCTyymNkti0E/wN99REenQum0p7+OPzeHEYa1s+fq+Gyjl
EyBnlcbJh1fviDYTdAJJ+cFQP6mFhIZUmHSt85NTBnE1b0CB3kDC0OniClRrnG0F
MD5a1iSJOydHAVKmgriLxNiu5/UABC7w2fy7qyZZKK/SV9XLOiOzrwbO+9ymJcQp
nmSGvIKymkoV9QaD4WxOtgrn0LwJZuUNCL+2oHRKk5I/oKyqQTpijDZh95JKiMkG
mgOfpVsmozY7HpXRNmKZ3Sl84LaQCIivewIUf3YGtWuGHwWsGFTkzCVrdbmMQRZc
HZL9tWzQ+kmMSJGm1k+izaq8HWk8hjOmzJWgQQAbUsPt9bJDDDJ60FlXaRTqSeIP
nti3I++EaeWQ38yXC26a6PvIZy+dMilxk2DGSxiT0oKhz0J4NcC/uBcktnW4Ojlm
wMlxk0vA6Le7iGsSqBvQUbNx+FB3ZdLKUBnyCaABXvVtvH3TLeW5Fnb4hTyfCoPK
nT3+k5VNYkj9wYFAAQNhqRtnqe47tcvX8avuaMoB+is/DqD5c4VbR3sDctd8lKhE
TOYrbdSYnpFZv9LgC2WSxO73B+5BhVvq2IJq9NpDqlFdIlAkx8KRtX1TrPN+COxL
x2ToK2HHKeNGNqkx6MWNdthFk+yWUPBbjeZBSp52uTEXZVz3f8MeGz5J3jAJc3oW
d2robnupMOG0p/MWu8Pupkk+csVe3BdCD8GTerKMKyJIHK56TorV4rJh92WvdCxo
+dfaoP7PfY+LtNV+iv1WelhS/PI0xdKCKMLNVC1F1T5S06Ea5Wqf43yCkuSkFoQi
7uo6ZZBvYkCYY6aIV2LqQwg2ckSZTf6VE7H6PeJ70vAwugk4ewzGN8yPKGNvQbOc
lZB/wzSvrwM3Zt+h5UwfTa6dH2e6+qaYZtu3rw53f9IzEgp29Dhx50nueRPxBgRQ
n4JFy1EfkDIaFsyNENcqQVk3hTK+MO1thyLdvoRmglnH4J/YKG4pk58HC6X5N7Sp
0JVGvwokXpoKULYF0/F2sh5FLdP9tU+5ewWI/Sbin7S1IpcCcsonGWJuDzkujVM7
soPEQOzei+SlDHtKwTui80udm7GoVvZ28OhJXmDM206UKimlr+wpsh/DRTHHMIwq
PudNo9xOVSSh/qeNG8hcaG2HVNFr5vPXMwGz0S+HjcLihHf0JlbZq+60uq3tnZzu
12rs7zudwC857+r7Z2YYha9IN2YYmM5szntALXbBJGfeVV5w1zmG/2wCwYJzpms5
nxSXNhMEESkSjjs1INO8/W0Uc3cRZMCV+vMiBwOMMa++wYR/qzwI1eBtz2PvOafC
K5KBlAeJKMtOIeEyyIvcTjO8ZADt6AJro40setwBPJzArizkHeJhLOTNyOoI5jCM
bTN9UYB0ShEgeL9M9GJgVva14Fy2QWZH5xaFLdLLXqHh6EScG2D0+E53WXCn9yWY
6hZS/PUtW2/3yTDbQlKbs8uvdbYdAs53IlYTDpEz1LGfnEb4k9JUjNH4Fy22gkBM
+Ct3iV6X3XdWyuLPhTaI7pB6YPwk9qzmu9vf9jyVYoN+laMdIdRLbwf+Be8cTk6Z
fen8fa5lG6oPNqf0K3TZ1WNV0rHHUuqLxTrkl7vsqqW5Dn7fYJ6aKTFIarjPym29
dHk0fdfQROq2rs9CoZw8P+p81eahsEDjZpcrGGvd2tIDSN8IkxbjjPJ/LGaS6mpN
wMr9r56zFPaLC5bEadw2NKQb0Xie5sQUhoXOqWqoAPNmBHEXJvkqlxQulrN5mjNc
1jfeukVAQyPdgFoAXyQrytNr4vMv7pKrtIf5JuPcjv8MvELobp5i4vInVEOHemsU
cmiIN/hXQqMCujM4tTDtf3KNL0dyl3pgEQ+UMirQ71SEUfVSlryxwyRM4u4Eg6Wp
xrW1iOF0yZORF2j9VyTvR2oZNJx+wlSitu7UXNA4Lf0zZiL9PwJ9+PcohWp4oJlA
UllOtB19frC4qgR/iVwtSP2ILMUH1cDHUkCx94v4qB/sX/NBtXgSLZ9vOKasTymL
j56hwibzhA+NY+fI/9H1MyzuEpAXgD+5h+EAxmRcKxUk0p21KyLY2DufKN8/UFS5
NJT8pw/8to7KAPAc6B33DrbiXCLFSEWxNpWZTWBZWlAnORNAgR0BIAaRljVryTDb
FRBQShH7By/OFn8Ddw6HSVVc5CMCN2AP85S0LigaIzF+5cxhEaTS4TAkc+o/dUP+
aQQLuKoKXejLkLWDC/kEHBf/NX5F61njO1NYMSoUyFkLfJhRv8z3fTcavKVPl6ch
tpmyTUnpupOs9KAeNA1d4naC93aYfTpqx/bld+hsdZOwtbt2vkYBI298MzXDct//
ZEaoTa36Q2D9A+eM8lEkBkYv4Ee/fqZG5j/tlJfORtEeN8rl/wbkboXX0tPDj/83
qOqqcXZ4jlVwj9jVWElNZelQGCZzSLMhsOtjYr9DTkAMytTTpjN8359zLUQHbD+v
k1ZrmPFmBYbmLjCycgVsLBwq4KjdP0AF1f9vAuReOx43EEOkhdS7d1Drv+JWl52J
xxeay+69w13SdTnO05MRHTHZ+SQm76clyTewFxrhaIyZtAS8jvysZJPqlWqJ+kt4
wt8fmzXAr3YmH+y5hlQ+VaQdGCYg0UTJE0Be3DR192hv9lxHdkp+W+XaPQNqbQtJ
oxPz1IJl3WX75hNTB+szklRepT89V8uUS0unmNJrNC+Lzkb6MpJROWc8yhEOad+l
/5zfWaqcaC/Dr7jjvdDcKS2kPlKHQyltoHwUrGJTpjL+pWd5718l6vjLkoYrSdme
UUZK7NnFw5ndNMGycBaICkabrAT5y5zW3l6HK1mqPxLg3YC5AnmlBIWbEv19rquZ
FKcdd1cS7EBV83lGgmDAQ7mYJw2qWLCbFjaefcPzZEPrRsx49GcY8YHA/DeXygrQ
2uivhUrz6JqXnhUx5O+Zqk4rlMbP3vBkGsL3s5GT2ZmGB7p8q/t6gKHtOZRBXOyM
Eth/2qeEaNBcxXFHeIvq6UtE3AD3XkJZKV0JUBU46LQWZ1Y5vy22MCOFh7hxSbX2
Y+8Vm9NJAM+6D0/PEnSAAXamcuPV8RwN/u73SGypG9iMWZ7Al2ShdhOOnSS9jjZg
ZMHT37jJ+cgQatOPbPSAEY2dL4B6nPEydUcQthKzS5M5lhqsWg3Nrv51CucG0VWu
3K2XRV3H63goFLiXSugc0/cuHiLAC6wLrAzemXCv9g4uXR5HneoXNfhPdC27Xikr
Uj6J+Mzb86LBRe8Awi2gUMPGWQPLHbrS/egve+RK2bq43SLFGxFBq0lxQ9JCuoyP
vx4AqTPPmpFCEkgbY3g93OunqfNbl6KdxcudbpNDtZEXw9jPZOx+ou0CTiOLa6DC
1+20NJPs7vaylnUsl1nMD1wWZi7GI/zCE7l8S3NXgiBJiawKqtKdeXF+6YPsfw8k
oWXLkUdgNm4VQB5YEYx/mm6ja1sUaz5ovp3Pb0J1+6/24F6q0jBnV/enMAYyT3nu
Xi55UTezUhz8qK/lNLCEhykBvwA79MBr1jpGM3Azba0YifLPCuaIl7zKhbWcEzDY
Mz4e1qB/F9LmjO5yO4E+oGYQ/4tXpBBnvyxfvbL3XkkD6yPpvZhhIvoBkEPUEo/+
tu4Ss5PbA/5Slej5DhiXz6gRMko7Zy598lBVWgPfQINtWFVlkaUv+0/To79hHPSC
mt8ogZcmM/h8b19yAGETH+ZMqHz0OhCQuEBoZpAZyQbNSUHB4NE1ZiBiDQvRC8V1
7Z7zCHkAggqT9IXjl8hCuIEdwFQzbpUdjfyCXRD/e+MAGGBBHYmCFc2cHNt/uIHl
/j9ugl0w6vPVpIbenyGBbbKEkNWv80G8Fc5lJOS1/42gJl/zq67r/KyFmDQ+aWD2
WRdUliFjGkKtjJUJ7wKvVteU9IyOasJekjAhQaUd3LBg/L2NE0M+Gj1X0mhJW0GZ
fm+zq6t04abth+0OaNXu2VHVNMOHC/UNObrQQoYImFYpClFRfhS1eWaPH497zcHO
XU037w5wYf84CGD2wKIp7UbedvtlDuhX7F2u3XFsrs1V/CPJw6SmE40fEqjxmxGv
Wdg6PaE1dSinYc2JK6DEHYIUxoEA34kT0+Ej40z58sq2M3vfjNVJpFMaUSVjue4a
FhXqDHTlxIKy+3984DO0R6NWddiUGGuDwjPxUdk16EXBhCa1xAMSsjFiPxAJNnXn
Oj86vyt3/y9BPaeH/Fm1X0goR0gkQ45fietCpeyG4a39j2FicOMYzDGAZTJPWTRx
ybSLdebqlcP66JcNuizk5y15EUh5gu6xvXxBO/IElUK9gS5ZjIfa/BQYdrQJ0J22
9FXR+XJW/mUfTAyG6Nhd1F0PL6ER8ebJljztu+7Jf/vdaZpb9knAFJGmk6cUTrnw
bUuxGC8Hv/vjOuX4FEBeyyP1CSoVfVQjWaTSnUwnqtszMATqVKl2obdNQAezAdyK
WXjJU9PfmPB7d7I2YuUkopuFuLwOXrTZZ2y47nZyTReP/ca3EXbRhWxui/hD9BbR
CMUqri6nBPeHaKe10QbsQn/hxmB/Q5dyoEdpW1qu3KbNZHrs6+28JQ4zcGDrIVVM
1vOUben3J1+l5tQlh4F7UJeci3fieCa5mBRrp/fHY4xKJHki8CojU5yr0cUug6ev
KGOcKgCECGJVUi2nK/4uvOk7kHx+2YCEg/3o/YzAZqdqDglCCcHpkvJC1OUBrhRK
eliGU8HinX/F77ZsBm4Mdcgv8ueGjhjh+q040f6PRtDcujByr4SPXFdPIe7ChYsj
efFdjPn+8IGFBqfGynP9/h0JFgLerGuKCT0FxR2iP+IFuUD5/MmGsBJPUzuIQUcr
3XrN3mUMGFaCJM6LUiw85L3CfdCFQKTW13IJ5SKjgvzsKvsNmcxN9m994TDDsWZT
sIrwWPco2laV9HLW2Ewue/UI45yXrOg6kNBIQTNOQJa9nyXu2m940VbMS6wWNYUn
K0Mn5DXE1UPewB+NiPPBK7LPbHBfdFOwDk+wb8pKDgjdy4sC4ksliYdE93Du3yQO
zrVFo8FIfYLSW6sYsjDoOT2tq1jpdObrU4Qz/pHlNwIF0yVEmaHxqBo7UUP8mPie
VxQpZmKdROs24sVwoM/LXjoIBC2aCkzskOq33FIpyBRcjGxTcyJg6JXDnpo97gFt
IoiWoXn1nsp7ttMPgOhP0K8e0nudS4x5jOX4ySkQbenOqaEBtgWCfacwBEDvIEKd
Uqxav+OvPdV4a5JuPbWFSkRRwdz6ldR1EXAsdPxy/CYqSFKP7HbL4tzBHtKFKjMj
OPLUHtMCUtrZdZBsUuPJhRSOyz53EbE1MSmSr9hvGxqBhKSA1oPI2E0FBHa1jcds
Z+p9me9T8JDkWiwpRY6F4cZcJm7ioW3UBNp2PpFoTAIpZFq/hPm5pzTtCFTmo/H1
bLN4hUmkV/WTxoh0rFEGgheCQZWJtkJ5AKb/NxcDLukVgozNOV7aznFAuwDllx4P
GDjNBU0ivRkeIWx8FLlHc1GpTXCHaSwuCIBu3TmGvvZGiU9+XmN5Uahv1miXwJ35
OEVWcrSOOE7ynDFmIR1BYC/mux/vHE1ZIGEZFr1JRz+N0CrE7uJrtB0U0CRmxMt3
Gx31rBm1bvnYJ7ck32fY1QdL5FAN0atRICuqNlljvq0Hxjq1LfFWBLU8uIzp5D3t
BrLV+FpaWDGofS97xcEcYI7WUIh0fnP8KPQQJwPm9tOtTq0H+F7F/NtQ0lQqhYa6
KnT4uVOWCRycWXMoOFqelR3E9bntW2CvonRM2qWfb9A=
`pragma protect end_protected
