// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SJY+p7Z4QqYd6TSaHSo89yAJtLo3ia1UpPvJtLpz2obw7Fko0jcgnTKM6NdcvNbf
IsxKLr4QydvYKkuVC5MJj2IhNuys6yI+mnHyiLZWapgiT5bHR+/6roLOXt9DcHjr
GVV2YUFSkMcAtDRzHdA/M1v7Mnf2bwJ/8VSAwgTr6ag=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
27OmaKLfxXaU1ps4f4gXdQ8FZSFhUk4ltMvXuesasTJeswuDBUx6U4z/ApnTuI+6
zGpxlryB3H3vcpOfbP+EE0xqGf/zvu3EbN3vFgYjLgo//VfCACmwFPA2GUkZFOsv
v+hYm0xDM5AOIwdbQS/0mNLp3Bo8wJIHQjfRHa21Cin2dx4bNUoWySjWefVbLBp2
FBIsodVNexsabnpvsqZFGrB0cqkdWimndZ3tpEq019U4UGQE3Gv+PHw9isKv6EHs
8D6zosv89ucnmOUWDuMKIQ/905C/NSznZ5l7n/3WiK6PjnWvtY98VmxG4zqgC/5I
4Xbc367p+uIP8rjGDzWsPf4x9i7x5pSmuV5DDj5C8VnZDmiiHq8xk6XRfuY5nEV3
U34mMh8gPFONHqVhQZECAyz1ghnf/V0JcVraCUEkuR/h7lbK4+XEkMUnEiPK29nt
ZPazug58NZIUmlBxAB8zC+GvD9fHFbgaUtaCUuyLFmaIb0iC+h2zyAGH5gLrbLWk
DKdUUWb0xAOm4c8H8wyj65WplPYrbVNclEQNfeGMNqVV6LOQaGACSGVU/By7p/jD
4oHEjT6SKCWZ0d592H9qE0yDV98mmeQU6vvg3y35bDeD7FtnvHIjVCK1zBkiq50G
+LERwmXbmx8++UXPtGYv6cb/2fLdM5OW60yxE6kGBHsQzGe8BNPXN2Nws6f+WhFF
dbqlNlQOcH8osoJSzz2D+0bbXWKD5gQ4QIUJvUyO4dgwd05Dc2N+47M/iLsLzL1A
donPEebRf7RFSfCxwQCgqNEC6ebLRjLalsZNZlgb5rZ47LbPi8cR25Nvd7AvpxDr
hNVO/K8BlQWtXIJZtRgIPBE7emmwAxGCINwbCXtJ68G3Jq8VHM5+cLXk/O8Zm2WU
/cKct1m+ZSL6rLfLgauk8vAAyLusG0P9J2/grK6n49ZdNkr9bfWO8ijTnwGzbOp8
6PsMR2/yfY74NpK0gCnhtZdGqErERwieFkn6qZVPd3pCw2kY9kFQhk/sxaDrE7zZ
ZuIUdEi3PJ8nEK8Pz6V8FFTYMykQEujysNaERDFjMbXp/aEyAOXICgC5zcnM0QMj
jJZFlhOqy3m39tjUCz+PnC3Y9VKjqXNZuzlbdmwnsjxnvA09jScWGG6cIywK5OJb
QplvxzpUESNlmm30IDpjoi6ffSQuSXaCsE631oOsBOoKXw7jORX6R3TIrnk383Qw
0cz7Ycp97M1/lOyoQWcHnVzIcsz25Vmo4tG5kIsL8lktnR2+VQIWIIlmE+bsk+a5
Ff4C7OxC2GlmyD7AEm+iGMWeAlwWtRtqfknHjaWVmVktpSl37nPSnBAYzILgea2d
m0uX/UURRd8M8/emwcu9lEmj+lZj+79xqz2L+ERFdrKO4nYnWC+iF7D3g9Xb60WN
nq041wFFqKV1bucH3s0daGXQZOSujG1dEGs6EhFNDVzb0ptOI5g3yG6s5MtWanX/
pmXh1i0Ic6XuUQne8KQTMW9Ai6knG7v/2ArQ7bp+dmzhXjWdHRjBC4yP9q+LHleo
08O30TUh6NpILk2TLjDoboqR3D8wQ0zWBxMTGhK09ltfM6pZKj7In9S4p6xyD2Me
uyuaTKC71hmddJhA7zxYnnONlYoXLfnuimPESJ1QEINyu6KKEcIMJHlFXQO1Nu2C
XiZXW7YotNlbohwtplOB5MqUXG4Tw2rvbEhyCRtbJoRRKeyl/LLMbt7GQRjZmYH+
hSsFiCU9+eIoBMVp7fWe2cG220OtE+Jyv5SixvEMppxixAT92yiGyLhjk4KQT3by
uUAdeozBFrIl2lva4ViKUXg8FMVEzsJLdrlr+mrQflyMr+ZrC1hQE/NVC8AHsHwT
iukrrI8YIMBgpTlGV3lX1dBoDeM1tqYim0RQVG5DD6UN4GJwRYdIHSz7ZnQQLe3r
hCQV9oE1BU384zgSRE6ldnJxYnBTreHHtqd6frK6y2iAqgHgebB1+Z44r+jcbLdL
Z3J3GVqkao/3pMb4ov84A1+mR1LcRlLLk/DqTcFh+i5Bbpv1hJ4OWDjnWM5XoCI1
MT4BXgcLrozPmLfM+QpSYPN9mWPf4C5Ab3alpE+mB8PvXgVoTywmWGdKzz7xul2v
zjhg2b0pzD8vtJesnqz8ybC8J+5F6gDXQe+cAdbggBl5QLoaDmoeJakHvNHfCIDc
3cKhFN88ByftAV7kvkGcFxINdnAvOjQAIpHrCZctskGEqoun46FjJSY+PxwFq8qE
OYf3XhvaCF0sjv2ezbGgSTomKGJ2a2RuOOicGgRiihLRvx1KW3JjxHFsQk0DKpcP
jJ2lDPo+g7y8Yh84M9YusU36xQOF7vDOQkgyqp8AnSupnx1jfUw67jUFUTcAL9Sb
COTfslETVpAFyPDZ+ANc59VB6S+so7P1g39jfNRqT3zAr2nGXMRBSKMaUzrFmnN8
W9Ty5XnAtPw9ewddlyi8zXGkDnmwha8FT8lyVE0muWZP9fWz+uecMfeCIF17YGx1
FMXtjyVSwIN+LbNyRmzoX7o8kwWg/NwaFpqIhHlc5eQFLrr44l+yO1LwXKI1tns7
j+sCfN8orAXVaQ48Ps/c/CsNGtva5eRcpWIavkTvh9T3eEzln+mz3PIaGBWmRX0Q
TEyD6a9+vu0e8R/m10VKIxkXC7vUHFyo5wiEqA9Zr63KNA8AbTeG6gryecyAxD13
i6p0NB473wtc65+awKK/9EwSgjUsM70MdxgtXnnYjgijXUBgxma8SOpdSeOjx4mD
pMNFX8AHXrBQxoDj7esUohjSga/rSx0ICOY2D5h/XN0i1M4M1ldT4bb7sXIPrCyt
RKpvg2z5xIM4GbapncBb32QiJjweTp8CnoIXj0qnHZJj+1FPn0rE9PLpcXgWHQpB
o9Zq7pByV1U8GUKSP0Oj/cTfz611ibz++jnAA+lU2dg4doPC/WqRC/0JQpYZnHeh
Fr6pHXgZlTIcPK0Y0pOUYjjEsGvOKrFWmXm7v6ZDyPIMxMitF52adYS1nl5X7pW6
EG9lWSr1zP0E2wzmGPECaLCgXsHcBoDRFjq+XSiwh7kTsIMeUc8O32XytaxeaxNG
lXsTZ4XxIHAxLwFN+ohztQlw5z9kEnGY2B4SBdW+nIT087lje/kH4gYYWBeko1br
aiDlo4BUnezBQBXwRIIbGni2rnnOZau8OjwGx3BxZeQXsAGcN/w+yMRlAEUU+yam
bvYJyGOrxQgWYbJ7wW7KD0uNY/GfCB6aSLp6Gn6mNHtv/D7jsxX3sV92e3DY84OH
ctx8teLp47cWSP3j1TEyLA8eO1tjJ2lpYZxv7QlcQZITtXgZHfmdW84VPa3DNGh0
6PXzn4YguU/A/b+sZ8J63GETTzrUs1Y9kEKacafFx/K5OTw81alLMDIQHyBJIwUE
tj9vKfnv4TkcHPse2Krcao4UEtJlj2jMn4SGBVNXki71ZsKNdeWKIZb1GVn5bORJ
jcvFdklmMn9YS2/HO05NbHftFkt3HrkQ+geSw+Yz4gGd4KwsralqGed/8xPLt1/f
XEPGvzZL1zusWkJytOuChb4karX5d3bAmhXKa7Pwr32ANqEY+W47PxEVefl2VSU6
PgARQgn6ClMrOxt2NibbX7oHjSweLvNjIAHtNXj/dYKMHqFSyQhXuicat/qvBG1f
dimB3/p0gXlH0Jp+QqKRguYOGlBVCnSrTnkWpqloY+hAMjIzbdsIiQhYo2ySpuCd
Rx7CANxiZSTpT/9rFlrsbY1tah8QVz3QRs8U+DH6tw9p3mfNXYQs5jyWAfJjuDMy
jVyRylut3YNJDqwIUQNNFfMFIeKurnRWpAjf1NAUdWii3JrzB8e6p+8H/PDvkf95
x4EnJpeX+RQ2eosqWQXQVmvqKHQVblTfnFhU6vHR0pKqFqefbtGaxlVLdizUBzP+
akZqtSZbbj62bdLyw/wfKJe/Zq1JyntYPAzzwoKQXLwwyYDZ3ujONpp+AvuaAGDS
5GNXkz6Ar6rgMPBVcBSlPnt3joVcAuomtqXkFxBqFF8lX3LICrMb3KMtBInFA38Z
SaiPk7H3743a0+GVGHRBJL8qbeXsTWzB7F0gF+3q3F44Lg7YIsx3YRJcDv4Pp+MG
raDYkpaEtIDUFXucwPGvnIXej3fM58jCuPl7fGBw5aMTFoaYy3+Q0LAa3LRTLIEC
LksTclEq8+WGlb4zBvfLqB1jnUX2z0dmmwlzuA1CjxfKyCArzPcvdHeDtPxh+vsI
7vP0tj6dHMhCNAfA2XGn/v7crwJakwLdgt+Y5G1P/4BfmZ+Jxt0j2YRjjRtH1S2D
ETL6Bbz/GMDo//WvyxH2HMuR9apYPn1j/yWou/Ug+GZFe11KvgycpQeYHq2RjW9j
lzwyCJrqMJkkKh3iHlS1KgYaIAD/bGgZv5g57IP5hobWA2Nx34SYdlk9lCSPExzn
Qye4iwMvo51xkFmcQ5TRiT3dfoJO/jUpeRZ6Eywo1BsCUaqRnQbk1zA58zk5xDU5
5qsqAPNb9pRxe7Cpa8yQOk9tuXyCC3cYIe0h05aLoaGSmDIyX2fI12er7E+1mVt2
KUXM/bWmG+i7QVM2C0cfa7o/kUOu3t0cf4N2rTGNzRPWwXnYfnvW2VZE+4DS5S2n
0aTQKocw7PWU2yUCUUgVQb1ixh+EbbxR4aPl6lCG7Iw2Hg/qgqwZaHc4JfKTanea
LvavdNEciijQG2B+WN5X5GOqzR4pIYkJfx4NBlu71cXdJgTq0Ywc1/dfDc/WFMt0
xAFMt2rnODQzZp0WnJYP/Wj/9v+m0U4BRNTfrq7GtwYZtKTAG2dfIi8WZ1DMJA/C
aupmgantUYFRp8LRRdEV0p0r7ZPMJa5X0ykxfKjE/XeJ+9CqPpCq/8XWRP4HY/Nk
Ut62+ZHp5PNCXw2eDBGma7SEgHmJmxx8DhQnwZs6fWVzRI80S8OL2eDbWwLfYpD6
icRrpgRzLp1B7DUx4Bim5iUAWlcoDdMCp6cPUXPl80P3DLp/814xd3tlDHFUYMF+
Wua9OeWT8FBEqnpqW5PK0QWfwfkAWCvgGrpPLGya5KFsjcFU+TgCk0OFnOLZHpQn
SXBED1DfBASr7onvub5CLyFb6XJ1dP5eXKDX4O5zA36K5FxazxmAVQsuycN2xmhw
5Y/pGvxwd7+OB27M1qEMHFQJ5D7GnjlPNkaIYYrlLi/BeSkX4m06CJmLtDDL2wJz
j5y65KXCcdU39G4A+HuWIg9D+zdSmh38lfeAHccuEQhw/15xktGPclMEnW4Zbm6b
Fnx7gvV0XWeTZ82YfLP+NGpuvQEHNpi3iAqhQQ8rWL4brG0ABa6CFSYKSsSa21KX
dBXrv65xFKNKUlMefvK+8GCOrxJiAUoBIJ0PDBX37RmWkKMlRhvtSs7wCmucLgWu
1ijqdZ/rHZvZ/kPL7nFB7sKWEFdBN+PQD35jZXehK0Y39XRhLleVZkqRhZKC08BZ
jnv95+ny9jAWwT7u97eTnlrE0t9rkfG78ng1bdjn6xOKuLHHlVY9650sGWpzLvA2
jVAZ51MW1mbhwXb0e0LQxc3ir+cKimwFt+XAy+y29FWRWmU71KidCsVnH0wjnKuL
ZiY8uapXeZscWnMFqa/7Hj++qH1v5OCX/scJ5wffJBU5kpPT5+xzl+Agd+bH5TnI
tMIWwqMPlh0H061pas6xMoe+jiKryDpfDCqWuzYR0j+UxFLTrBAjkL3/Y+S/Senu
qtbQL2JNQSLv5UCgrSarKMeFMW8N/PLP0lCYtvMn9o6uwFwLSksNNyO+gu36EoKi
WDPtBC4jDVwvbxB5vgId7En5vL0ICCu4nHJendAcrzHtt4NtzUHAWV1Tta7lICzf
/5GYpRljlmHkT+WyCzFPjAqnoExaZQyT5LdsQ+CQnwzyagbUDelkX1ZZDcFPblWI
2C+P6qOrQ76Qy5bl+NdbtHLVQZtyABl9ovcUbGPWLEQ0z4Wd1CVyEIz19ankLXmm
w+WwrSZ8WKQjwuUKOMhqs46hAI3aFMZ6OvDAfpoGHeF6RkufUeMqs/973iIxdl8s
VIfnQxhloO1/7YQgCyMvJDMu2xsBVYfRKtIU47HTcDp3p2co6eV9UtUrOgTjPJ8S
vqmC3Le9iQABC9iO0AYlqjWspwBTRiRihmuoDbbe6UIdj++G/W4vbvCVhq5M6m/L
ZgmDf6EYAgbXC6ZdU5/WhFQQQ4oqtLDqyF22ju+6kmHskJQ5mo/+NEL0JCpaWAj0
e9+DRwmvUdC5j5nhJ9DZwY6ksCIWyfwUfIyjiB9+ShCNUyCulC3GwDwuQnKbDuaU
8ZMROUbQotaALtlbGFZ3L+JhKXu5thCdW5I8+1dGqsfneCdo3H9F6AqHZ4Cy0GSD
e/046C8lYIaKB3N832aDjoJ4yfrjwqFXkcm8BJMm9twwRyy3ty3pnZm1f3TG6px/
8z0KJECSVGWuTlxJbEjkJTg4O8euvcKV0Upuw5VinpZrhn1dfZGA3V7ZPWHgMnCZ
CVvudBHnTy5ukUs3d7Aq6lWnPphlSOHLIjj2vjeqRZbDJQg4w8782GzAK2yAznoX
LlEjvHnQCDJ75b+5Cw8W9dR0WNzsiIKBgPWI8lVd4dNO1w3Yx2PsHOnLYycnl6sN
pL60iT8lxBfzPHxOaW0E/wT5WUrckNQuEJn2g/1Gs6kjguA7yc1/IMQisI8AcKxn
Sv352bhYonPzLWxkHpQODws9dUzLdiNGzBrDgR2UjLFRUIiNV0JiP9P8BG2H3YOH
VWPIrGFoU2hrZF6Umh0xEwmqe03C1j8PSsYu3CPxNwieAekgyDnFoqyuNqNmFfQx
dQnq3sOgpzN4Y7/7r5gslxUQ2ALzZCChnXrBvAMAAcIiQdUD2iSs4faw+uTXJWh1
/Xds1/qddAEdwPx8d6AAg7IWO9G3wbRPvA/2NEIrmgIyAWwIekkUCs9PolZuUc37
2/Lu4MGhCf20hB1kaE9td0MxIOInuqrlaIysTIAyWRCbdpVwK8tm3vY9+fXGcFgs
Wqh6YfPfqRt3nGR7c2Iw4J7Z8h5M7GgT38pdJsAupB5CVlg/K4FhLeXzYBcCIWQz
051xKwfkNuqXHPxNSoLb3+lClW9M2vXmADDUqSOZTPxC1enEeY/hCQ8qUUokMZ23
EWXnHU8u33H+1hZTcYyzaLYvLw5P4HGG3YUNecoZ3vpI86iTQGqXpZ98Q8p/GklB
kmuTZOKua1LgPxJqKoM/QMz9DG7WE4FzIphf8QasDXoBWUw87TV06dCXyL+UsnrK
kcEnXPrSw03Y4oRXl4fpxI/RIwDZmaACMZFbzcTWXcMo6CKwpLCivAMnKsF1rwNn
pyox5c76tEXuNOqtVIKBwRfLGMA+L/rsjtUepl08SFFnYWUI0K9XmjaDS0h55y6n
3oc+lG8MNJSUmmYt0x/MKa0Bm/njTtIe0M+3utCdPT9Zl3yWid5MCIQsS11w8pBB
i12yrkZM9wIOoqgXqhCnZiTI7esspSG4uFyLtz5mlsdPEE1J+f76tvpAuxXZHeMS
i8vWFNfEW4eE14U0MJlJr3TxyVZYykvCV1pqBvBBTUFykHpa0prp5WiPLF9jvW2B
m69KzpZlgRy6FA0EMScvleqVeTZpKCAYIWINvt8NxIZbcdcPD7PkJUW6gMqnbDLe
bjZdgqAkSLBdsWjPPhxnI5L6icE5nQUbTu/SeXjydhoi27xS86jP8gq7NpJ5+nCu
OMXfOdChNv3JDGEJDURc7FWSfjkJdv+2ysi8SS/SjzVNd1Kz7n9r+UeFmBB1ToFl
FdHrHwQPn0+UJDxuskK4D0aBnzNZU3xk35q4aPDOhBEluLkXaGZlXcnY+p+ypURs
2ET3IXKl+Q5SYfFaN8gSMHm3O5D0DIZ0c4YvSD8UuAkmaZuQXiZ0FuKWY6SGE0z7
yvTRr1ZWmLQayJMm6gq8Bif2kMB7dQlIczCPxnfopzYOPv7UV2GaCXA1JJrHm10S
QZFetCOitU2GoYJR5eXGyUU22fA9tIoVchcHsmductzzbWxezykrKyyL1n4+4XtZ
jF8oZohtYSRF2/FgsQZVlvC8sVtME3kJ0y4AiDUsJ0lzD+cPs0pXE0hFPOXyPPJA
W7j/Obk6hh9380tIKe9X/Kcsl+mWReblWDvOqnWsWKw32fpxOMuSFajyunPpGd4f
Ia0Czx2z/sVyZ4VsamWyyLVxMbQReIHla8A67dAkzFYmE4yIiNkCe/sy/6CxlYO7
mQD0EcB9SqC0OVnchjJ5UHQaZSHQnPTzn77fTLmaz0F55GTi7O4rLUq7EKUYXCyq
EJjRFb8eeo3yd7N0RHRNZfxq33eimigJC1LXpgkVTlA/cOZ/SJLlarmD0YR5yUPz
7toccylaamzxj1xWAU0j2RDuUYLSTpvmfu1DHjMkBPuwL6jzubt9ZPbvmO+hAz0o
aL3urSky7SekzeBEDR3wtrJBMprlYNgCWmWkcDrG7+mkFHL0etuRtMuaAlxWMcP2
XoWqCtXshv2Wu/wSlz2MfjxwdyfJ+efjmR1VWGhNh46YOXV57x9R6swLy52TnPVm
JbuZ60MXCQ3XvBePbsK2jnDzPoa7gIPgHBUp74aM7mJjHsJusMzKOQQtQ4hoOPme
/o3CnUGBsu+30Emn36t81yasVKoDt0a8Kdj0CdvBCSiYYOfbC2va8O67g2uoSEFj
XrDr02pELA25A7j9g5JF9SHnwn8eUvApDY2oj9Y1c2DvuX0pVZZyXBtatPXIw1EJ
ivKd8wmdJhtwMt49Ftx2oP+7nNIHM1uyZLPkBwaTzG6SKjBCJMBLqniyvyo/bIbm
wHRGBfml9B3uZp6G21uzjI9uI5KWA7cDZQRbvIGOW17GkWqbOCCguh47LxN5dL21
IyL9prklrGFj27ydYO/2WPuthVdv4JXdXyVep8kgS/7Pcnhe664uyIJY9jXY7IZ9
B6PlMCuzywT87iUp8t5EUe93U46omuUabk1tKZ7t6VwOiUUWKUuphF0uA7JMCk+L
Pgvl41B5ppYlbtxOuJfm5eydjlreNCImJAYaFyd1vUYbxm9z64Un1uddcX36qp9T
DNfzKnpRrKXqr0XaOseeFNTepDbn6csJmLgjROLMS/UkX6h4FjGMABEe5gK1hyMl
x18QThSbjYOsjlE3xjcvadSuvQnBkBdGjTj5PQakgkOszDy879cdafEXezRoKfAR
icNXfXfgEHi3M4P1NPGz+4elODrsfPdVERtXzxZStuPQDwY2S3VN63VW1Z4ww5py
PCCfm1HKDI/n7gfmDwnv6qfeIHuEo+prEs8dN4M/7zg0u048lw7n9Dv9EoKRVPIr
joFNZfI6vwehEAry02hllHtJcE5aVtweVwT4RX7g7TAq2m19MDyfKiHk8KZjRlpI
O9Xk1Yf23ZhVlwOwu/451EKiNddkxMSF66LQsQGC8ZEBZTlwlPTZkekFtPBB9u55
3VdBrv2YuSGSC/VpezZdYH5tY2D7gpN/jOdOTflJMbpWViWNOeANM7cyinhzaNC7
HMsqHmTi+xST2q5dkhLPNgeCN3Mq7r1j9INhBhgPYzqfR7Sh3f/pom1IZeuCcwQR
ZpFJpngTjDZQCnIOTBimX/fkHqz/8mknJJsg99tWQh7htKrltgipIqUJA0PJLF8z
MxKZl63QFz1o3snRQLY874RBIcbnghDjVgqCBVDKTKfY13qXePIHdDTbU2c4kiph
Iq1us79dTKqd1qxRhGlVWRvWq1PXmS+vGLaR3f+Fh1xnH9qZ+70WL5qiDeR+aC/Q
xU0aghuAOXu26WwsHu5qHPljPBwThbikXDiWSrwHBCCxfKXJ4yHJfbb0Je6cDrnQ
ytcZynlnik9maGyxHgVE5DFcu+jeE4SFyADxg/SV0vOnGiMjILNLgSiO5cVqb6m1
NWVxILrh65UvpPDAkFY7vlMYdkB0gtCwVdk/J88LD3E2k7a4LnLDxXilyCWHZ+os
zX7l4ama1UUi8lwb+J1K7T8/e7unpJWRmHINkx3ifPSeVxLd3nyEavFFtm7L96EG
++pAzZYVg1srkt7190xOIGpBbC7O8+tU1jOlhkArpVZ5MfCHj6eDEtvAS3rhVl3E
NfKV/n6wjCOurkI9+ogglunLO6HOf2qIlnOyjPDUeAMKTgTVmIbUb7sAXtVGWmri
/w+L0YLckxV30bV4smV31pUb7A1PwgUVMqqduuMHNMlLSyz9VU/Tet44EzM5jzop
SqCZ2pQf49Z5x39hQtwYFSy7+xf/GfnKv1MlSFBpKVduTlN+spnydi0Et8SsoITG
l6OVO8/I4SrcAeS7wAbdR+M8aOqaUc4PxCzcUrPKB++RHeEitubAwzh7kGiNJLrs
sTHrhPG+uV8sOMhclsoE+V0Fw4ahEWHguH2QknaaL/wUTtW2wWeSmnuLw/2bbjY0
udy4Q617W0mIwypXRiY5vvGLXYrQ2rKWaPBEXHAhngkauqqcKlEUYOT4lC7v1rkZ
4V7vS0uOIx2ZX6Qm2CxzNlxI1Mc95tN5S0yAvyn5VgGNl53xKwptnmQammKeIQQh
13jg1fTxbrDKXEuQe4JsQxZwtFQOMokRKVehmWd/TaqCS4zNAFkKGJBpkO2JOG5O
cCb4ZWFmbdwtqq0jtqNa8+lHL4mHnPcnBhxcC0t5TqVS4+0afhS5BiO7IQZZB09w
yWgAW6RLPw2Et3zCGuKXpQoWmBz8bKAhqRo+edhw1CrzfKQqCVahVzPl+/FV5/oY
bD/C1cDIa/5MFnRjnLuM6ImP0GqjD3mU1hqslIUB7Ntgf/u1S8oLg7Rjglqv9Z1D
5fhzexjKKsZyniKqR0LOkmzUSDKLGkYduR8VegzBfvzrC6TJWF8GXXKbXmtfENEJ
/ROCUigzyAxUKwAwL0ZIiXoidf5RpvBw+nRfkzeS/6FgFvvFmYppIgvsEsTo5u1V
myy07kWHp8XV1jJQRd1eLYfDoF31rqkxYkuhvOtSBxXQuTZexOnyBplqOAiA/dhA
Wffxfz5Hre/1ljOj+LZi/nEwWrebfrtL+c8/fRmRrOfkySsvcZOJEZyzptYu+PwK
HvpUlX3P27u3JnAORKNx2wR1689nG17sHRyQ+dBJPp+yORjW7kYUuqI2/HqhkGUv
yNseFx+kFq8VkaGmTbJzBXPHlIOomLn+D7bMBQFvc3mVhP40gXN5eWpj47iw09v5
oCJ2LPuEjHp66b2aGFniDInJbn9QY9TnCSViD4qUlvhPCwqF+kRwS5DeyB46+JZe
cD53AhV7xoFas1i5uQpPIwsgDfAzm5vm5YrseaCTuI5KxS9nTnE/HN0ECFW7t3Su
g1pHVFvKAv9Yh9ncb3xS/+Cu1iR8wtg5gNd1byMPiS3TuTq/TdHSCT1/+qMwjxji
7Hj5g+FdM4/QFSucwIyWQtmGGG35szvKM/UKppD2fQCutmlWwLMPv1nGPnXRb731
JEz5I/Iaqm7896Ex0dKVyr68h5D9mzDgOKvyiJvIFEIvydSyXDxzo1fymp4KhsmD
eZhisfyjPbPyfXcDV3EMkMtDarLQVufA11zKsmzTZN/hIhgXdQGCYVbTQcs7ZJb+
TtsHjV9vDrUBJXmYxx+CNYlvEARWePleEyKJ1dOC2EsWWrVylxkNGBLTP9IERzW/
PghSNHZikyxnRbnYYm6Vvq1NbKAhmSDCihcPQOEtoGGE7zocS/nP1oYcjD0XjQ1s
rvnm4ckBx4jhOBFpBGJRfQ9TiJICjLMmCe/R7dLjdmLsBopTUfbwij+OUv0DoQCv
k27fne2b1ruP+0w6L2dDbb6/BpgWz+iEwJre2O8tQV2XrLBD8/M0xN5URdZ1CNKS
xtBkeMHzMAFcqtkh829hj1aNrkp4oxGQGh8YQj5kF08b+D5rDcJ/vNa2Ys3DbRNe
xgH6wYhbEDPSSPY18aUqPWslPV5QI0OQyXERZvMQT5/Kt5E8w5ORZzVY6R7ksmN2
FRIB5K7vypNR5ZExQF6sCcjP+GkoPyuVk5nd0Z8v/jZTBlxJJBlALqW6FbN3RMUk
Usuy4ScDN0jDHCNN4XoEwyl39MuxQDThxlz8FMfH7/7cDOmoZ89Vx+tMkSlgoK2s
CIXquNZvK6XVgCu7SVHjdSkiO0hYPOBe+NbSNJGjyzeqQdhZ72xCoAqPMXKsKC+l
9BWhBz5ZFHBjHz6AJSnaCwNutVWkcJCFwETKqUCeEIxBTluKlEmyjII6dEaa2Lsb
E51iU8P9Tw6a9SU5gVty3QiMXmf+6hahF1pPQ9GHiKr5d8LhYzcNVn+vEUExb38B
Fwt20rPABsIXGokOXQIu75nKEcBH2ht1WCDBkZA0O/4VMuYncdD9m7tvGD7p9P36
b2ODngqQtPg72Zlh4VP7vitCxPGiEOwuvQ/DXK9IW+s8Bqlg+/GLQ3bfu1bsgSxu
G9liSle14NmwYkFvUb+q/9e+d/zENXc87N0RAAf41x+uH2+ait//J2ZYQqYSSJZs
erukCB5pyhKigeekoZAoY9zkgO3NvXm+2hLa/YHI2fvT6Gowgy0HFvPOsAFBmZO6
DmXTjVrGHfydxNwnZWO5euOMqqqddiFrnq2hXrd4su37UcIPzDRkPz2tQxcKkCFH
tC9WwIrxtpgncB0977PEyAIQPPmfUV5aka2IgBadwPAt4O6DdLyzEP16ZAlvP6nj
al7+virXr369+i2MflwuDoG0pFOXDZ0ON4NFh79PuekbGYamCN2FelHlyy6MMtQs
MroH7nPTR5cej6SE5sgpr992pL+4E2GLQtL4g7QxZvOQ0yKuroUenVKfr5rMiZP4
BZSboHzUSEmUtJIsPEvMx7EUGRqzS/bTt97RXe42nxil2QJwnx8DAqe2y03ZUkXO
kCW2plMWn4EGZvoS0alS82E/f7M8/rHwoQWNzEffdJzcSP8N2lBik97de4jishnU
P0kYnttfcUMC+hbQ2DMiHnwEPVREukEOmxaP7kp78WakaZCODe4HfZvKZIQ/Yig2
P1Nq+10AR+VFmiWYcAcK92oyXeh/jtBgwiis9NgC0jWE3/W7Qxlue9M8snS3NAIU
idyizCzsbxA0VXRYW4OHAG0kLagNBfJKRFDf2dD6nsB7Z+SWXfwabxn1UgEr3nhz
oRkPhu5BE+Pz8wtbBM6vSefnEysGLmDAeR3wXku96fy9CWEA7J/VrBooaNCr+ARI
EmR/j3aCRcM44gt7sNBKjN5BHKb3hFar7BafKdiEA06YcFINp+bP465oocbj0a1J
A9tVkQ69WFRFCuSYX0HXD54o0ARLHkmFrYVSGEnHcagsrDcMEDvCLLwtvSSCz6pX
V1gHRGhiyczWL5LnSqbeGIz9oRGT8msidBIFSTQcOlrjiuBKrq1C3gmP+mQHyCwN
+h9nbONH2OFMU2B/yINcP/MLPS/DUh+LomiXzN838WhU5nS9zE8gMIP2rHpMncni
LnY3GUF10+DYEHJpei/t9aWiTuL1LrHGNUodngedqmbsWB2fWhcWDwZygIwNTTgd
GYk2IR0Mf6vGgC8fotedm9zzNT/AplIfP33kdyLHhgCyDNJjpddVCRqZQO0n5yX7
SNZj42oOjb2Or0yNgZZUTekvdiMn5G1dHSyQjuEaqt+GhlJQuWsPV1FjXmsoVoPn
3zS2yTSoOky+4l/NF6fWTw/PYRVNrZZEYPOOQ9RjJnG3vZLUBqcUXXBE+QUZd2Hr
C4YEAmPTyW1fgRJ7h5q5CtLgpktYC3ZWEvhr787xQengH1J1HZjtUxlCSoBiOR7m
oNnThEAlIYH1K02rYuiuYuPaeE/2+XivY/6iiQ0melJu2UJFyjhcOkrilKNDbyAs
awM4ED30fwfZGla8MJfe5nT6V1ylhzeJawJOUZFTFWxUHD1oQDZx5nbsI9dh57NG
W8XbpgYdEUuSUAFBGl/F0PHZ6utuvCb1CCRkJehJ1nKN3GhB0YXyuTs6NDigHTpq
HSX+YQqKFc3FBUfHjEj8b6hAXK/qdNXxKVvDniNAlvdq7nO6QCcZrXu5yTGNooEf
aUuEOV+YQ8kdJucbiHow0j79bJjYDg4K5u1Ic7eOUv4fONmTo+jrFibEnu+gocXj
ziCGH5JM1gPFOxd1nwgDLM+R3wtlO8xt173MUjg3oBKokhiIdxKsmy+9xfzFIxeM
o6hwiXgR0pH8wpOtU/6rx90iR8zn7tpshxd4zGO5JGNu/HTIWuDo0lEoN23ZH8Js
USmpdwRfgCSqUzGZEjsUZZg5qdCWMBZLQ7fh/pH1iWTiC6t+JKSup+1PF2dYDf5j
IObLjd3m0WsqCLCI/CCg508dA6pgJWjgybT2b/cioiIwNmk7bBqnstsSZLH/GzGk
ulhc1Dv+8J7a4yXG9nFCzuN489X5aok/qwf6d/PAP4iK1+cE7K30pAIcoxo00pqu
Iit0SQeN1GLvoTfM0Wlt8+JCGpkSqiHDu3ZTiHBjTxehEDIKM3nao/H69vve26i4
4gi+8b153TjKrGY+85uUHehRUeeIZILoRbH6BvVxf2b+S7Xc9o2iFu8gzjAcDvCk
KVxh0/bgo57tQWwwRE8qrgr7XS5wFiJtNJLUi4UPXXbnn9rgWMQouj88nra6YngZ
+KQo3LdR0KQxD5PP0QZPIIO3W6kw0H9n8vZ6VYveSK+hwN8GSyMpeeBuKK9PF6W2
Lcw64xAv1hjwd8+xqgazG3Vlid69ftJ7fgcmgNaTudCx00pbIvAW7AFL5VjjgxXv
ia5rdUx68XThKtfoJQOvMqS3KfPf1+mNLrzqSuDqo8b8RYQkhDKKv82tDFDMgBjJ
KKv/OC/EbnptfoGSGQzm8QJ1+n3aND8n9eH4As3kfX5W2g3pVuPEygYlc7NI0AkC
5WvH8WbjsXhHDRpsLlnupRMFpXK5EUWfgsyIIU9EUO9cJdHVWJBdsjhPzr9ajqlD
PVyiVZJrQc2Rv6nps+i5U1yjo84qzkh9dfva6/uIOkx6jQ6atb2X2rgVadfaxeuF
zAm61/b1uJEVPhH4zTVL5NH4lhYzV6BU13pSzRz+3x+h+3Zi7QWgmwVehwSS/5OV
jVzeunOuUTTC0IQd6OjS0qQkLy0s0mk7sMNI1RnyFnCBal4DwEQwJKb+IqUFHoVD
L7erMYijdDvkXwd228FEDlDf2tb2s2s7UgAx08itsEEbI0QXwtLfYNNNosb4RZKl
BGRXqrx4ppOZQCx/WOuCg/+o7Goiwj7m1py/EUcF7/P8dK9gjUmBiJ5SJbqhWtTe
xb7SX71lej6KPE4oQ7QmpOlU8xUAu4cUEsmsOPuJExxpiiWbBXmnwAd28GCekicx
/lk4iADhvn19ehGvznBlWBDA+ni90XFUuV64iwtbgHgbjBq5IXke6/IWzxhD3inQ
ooZKQQ0xtCaTqMEftv0aNkR0pRrNnEz+PxO3bYPlZdu2HZTCrZfWrmQIJz5wk0FP
kt8T2u+qWm1yZPTOE+AnaHc2aQSCmJNS5S8sJnsfoe+axDSJ5doU1pewblbpKi+B
prHbTqKznUvIA++Vxt5eq0XYRYkpAbOiW3ybF75PEWcGXe3gyzpF3uTQ+cA0j0PU
UpQTa8MubJF4WUBZn7lo2Xm92VOUgCIM5P5zMnKya1LTwKsiPwY5er/HgP4CXJtR
CfR3ImjW1nX2LMIRO/iol0jjHMR0t9uYQedFCeMLUr6YHQRBtt0xFS36VqLkDsde
TJcRIWVRUhwv80TIc82FEavkiueISpT6xpi9VZ9g2QPtRwUDtUbrzibnCRtqeOvi
35jxmOs70N6y+9PdOq+iJ1sQ8JWPKMbrR9LL2y9j+x9ZPZ0PTb7ZcPtQm5gjt0q3
zGaJRBQY2jqhlR6xDyndiHn1KXrwREgV88dNI+0z+jy1GPfHuZ1FQSbYRiL9+Je4
M4zXGI73uhcKmlpG7H0DrxtBk9vOxWWUERqF185MTIKK/jY73BCqomJeGy+VPw4o
K7gmulKDsv5kksdhqzszs4eYW4FlzKNw6GxaJKiSDMzU5gGwJlILQyIgPELgHytX
+CFbH/koycRMSr6iljrk1g8maVZfOP3u1gSE88czD7jddqLRO1gYwKZwoj6cZqL5
/bx5sxY3YJ5t9i8kgktvY+YKCPLzrzhIYYta4NXzZ0JPTKYKWv3BdzoSrmtrtuO3
qHwt3JzkFgs5xJ6ABbngc35BNQD3V+BSS6/En8EJXS4jcAIIC6u0eamA1CzC9Xog
+uKsRPxB3xcovf5zxH5Xc3zAoScsOAhy3eVe7k0RUXcZZRzXcKilarnNrQI1mAf3
PPJY1wvijfKPg8GtT+88s4DUv1YJsmSND3aDRUFhPWWi0LuaMCihxARNGwpktJ7f
xA3yCvxgmEmUeot663Lo7CSQNRqmuS/kmRErzDs1nwPWBTK/hiefB6k/DXa/tIBG
Qio0CInsoLf5p1O90wwK8vEJJ26kLZvEUmNrAa12tyD/UHYeD88ICBbRgfxeIV5B
/mPf6xei62gIsWWplesqDq9z1P5Ez9kJnCQQgtUeWC+e+6ClyoBJcp2ICOHtYvGq
kDUAvUjxpqegqgYJOzF2C5yM2EpN+5DHSu2y4MvTVYlhRRaXfCrRyhaUx++uMyyE
aH+n1p4MyNApSbaIIEGCMFz8Apg0nNMgMsP19RO9AwIFBsycKQOPrPBPf9DtfNd9
P8+kP2Tj6tzo9+lx4tOCQFJBArXYBPoiYnBmGExLqvPki5qydd2yiPAk3eBuiT7K
G0n7sNyUZdP+L2fbSs1SGzG6+we9ZffOF4xm7C6z0va22JLtHFCOUnVs6gmp6wfg
cG2srsPK75quBLJC5+GptaTpFlfWNY1BZiAwBHgUxQWP6hFDuQI4GbhsGNQESats
wlzHsVWs2/L7y2b2m4TzZNufz4ERCzE+HzXePqGS3VyT8wujdzabqqlvuBeTFEGk
cLakw6V8ezyUie2UEgz4vuZjIoZcqBiGx1iEEOD3araMRSOrTMAumDQuwzxq7T5z
nEtnv9lfuaROO9IpoJYdgxmsSPk9iUyTss7rdWOqQSsFbITCmmlEvL4WxSG6xX6U
xRnVrFjFZUySHS4GD9jufrBkmqjpeKM/SMMI1PLz1ski5nnXXFd/2SKewTLV6FIW
YJrKUK5B/SOwfT/pPL+koYHOw8LPldRoEMMJ4McNZq+a3Lrn10h7X52jC9M71+ue
5gM6cD5WCw4zRlymOB3yhn8SzzpKxWYPgZk4tuNfciPTS3ewYbcbcBt2wpPoXTl7
jzbgQA9cRyRAmlCZiQD5m1HUfvsm+RN/0REJqb1AsRxa8ArlKb0yFF/nkcUVE41b
3VDFQbQlVellYTWJhnZlxk2SGTI15q1IyZymuFxYSANOWcu1D/j2h764xq7BewZ8
bqb/7UJ5BuszJdLHVbyKZ9Llqe++3jpQI3bHGyxP0DEFuNjPb6L189HxIylw8kNC
6fuDtnLg6G+ywPDGEmwfOLhHAwMjRuRgaNJ9kXoXZmo9y+AUdlrOiIYZvPqP0fkB
R4IFh73Hw6a5HJiJ4FErulbwFSX8+VArFWb3II4NMjzLg4yMp6WtJ3mppQYmuD9k
426HNGX3UOAti4dwfNSDkuONsa7+qN4oe6zATkO8JKQqwelXNsJZE9iqRyfEOJAI
EYjBnpEo/iSeHofVR2OG3aiebj6+KUI5tVGfBosI2YGv+iOXqPpaJD9fdKU9he6a
6Wt/eBkz7ie4wIg2d7Csk/t4k/2VFK3SOTCt6yDstESHYZxBhSFpJEDh5DPE3DX1
4DzpLy5WFlqOiy+8GexuGVNb9VCXyuEMF2oKueUyw3ZzgNzfUTRFIeEB5OJNKv2z
HuKQpHXnjJWcWWyv4cW8QqTPRW7VX+821qLXmUNwwZYH+zulozUqWYuCiJgz33FF
I+XCI3S2ht+cEXdG4KdPSuycLun1vDcljHxQT3StTR8ezZXZvUX59MIYAH1q8ElG
iqlcCaeNoLAL8+qdxsHvMOhp1Fgw7IgzKZ0kaXEzuysvcUpdPuV41A2vk/23kKT5
hVUfYUIKoCvTWjwi7b+nACZF+ztwB+TzJHmUIKsEf7MSolJWXtS+EKPRar4KTFjn
ylBtGIxMsOeRaO9Hz83Kaz/Orsm7ZzTFaKrhR+7ZucIRE6J2pJX3xJZBpW97K2u6
7TTwZoe8WGjyTRn1RKSU9TSwu7iQcXxhFkhWUkHO20CyenROXWYOiFNb7c9Ahy4t
/Mbu+6CzjiSeRtT9OvnvzwknvY0FfGwoGPAoGx0lGkDcFqDItF3cixszmCjl56uT
Vhiy2QKP2wXIo3EKGt2TVDSPMVr+oq/9SfTr4291ukKtl2iAl5dzAi0k0vDbbuEV
+fnlcjWU32tAMMhTx/SoDAtOlzpmkNa9Tju4qIq6XSdLs2ZelYbVCDchr2uhdoZb
/k7F673sjcVg+UqGGUKmQU85KhSYH9Y7RYav6wnhdogdkiQovkntWAJ5x/pbP1zX
ZpqLLpKDWjHCMdNSQ57f/PbLeUSY3a8pjlrsGl+b3QEpCVQCz3B/Q3RPTz8jK48W
5C+SloDz76eL9s43KiBzH7czYZm+KNdeE4C7snMEOEeJBuZDG7tnh3lFxfvZPZWs
LDKuw0796tEDlcQubX6VrF4sxTYzLfEN0ACIjKA++4yIyhuIOJzoj+JTUeDbVZ3d
i2bF16EeccvwtcqGWHWtzs1lzIcNHr46xJNCGt0nf6NyL2qLDRRQenyqknxvp4Ax
iVQWvuaYbGeaY8h0c9rAWpdhXHSePGpLGaKhlhyHdR3oFHv9KoW2JXzAxiW/659Q
uBj+IyTWg8VMetIwHZAfVib0WpwLotHWPK53axRQZdB+5zIqo2Ko1tELA9FxRC4N
jgBSFvpuAE9vRC+vKUascuMX/xRW8rPXo2PZjCs/LWNtIg2kxdfqEwVegk4UDjfu
dZARKMp3CdkTZc75ihiKOp4uFbEHqOoqLNVn6Zp3y53g7AIdnSFYRznv6gjoNOHV
LYvnHoP6pXEru2k4ZI/TGjUEsjXoLWBJ5RgBNfVrh/2hnBUb8ZiscMRT6EE2gJfe
WQcVS0AyC40aw6NT4Vjs9dC+C4c1uwdCkC+xhvnehMb5Uob+MeEnEYqEnGXJZUWU
p5ukaF13j5ufV6HStGb2WwHjY9G5hsQOT1IIDoLu5PXnlW3RyoXYNIF+w0fbcHLL
Kq4RrfhBSJayr/SUUMr5DkPvpZAtIUgfGIWbeht0VXtVkT/1v+9kH+4O/nZIv/07
BNTTnW7ITFe/IvqGgvuPgwSZEiEQOVjlhXoFD7T1K21/BO/NC8Qv59V8pzisZk8X
yG7oVNDjDp9tkyYO+GdXqb0AOEXXy/bSO/YHYlM40BhwmNwTDfLFaj8cA9nolLCl
ZUP2kTzYPNIHuvoOnKaghrQycmNlFoXLwSKOyepgSNwFeOleJp3ERgmL8we+TGIt
DP4xXaUm+PKQlijEJKPKl4XUmNkqTadZ1RuqjgZJc5B5dXUzOn3L4VAEN3R9FZEd
+3j8UT6G3Qku4FLqYXgQp7fA+uQO0IwNNx/BT7Wh2pGMMMZrRoh/hewrD4NSCC/0
bnqWBB92tSGUZxWMiQhHo4F2BT0oYQLtu0HEd0akAHHE8zVgpaD/0MbcI6xE95Eq
NyHECxMRIyPyrRNz0wouyWc5etaYGQs3dksPyvymul+C39pArq7PvQTpeYyzLvkT
FfuhhEqkZdzFIOLx185tMvq8VgQjZzUITWu1KVj290VmZC6333hiWwhBSRFHlBJf
fOZK+cGAlNX4VMxXO4BsLWN56hRru+QbrCbYPMggsm7iNI17bWoi7/OEyh/bwky2
HOidKocgu9PgXE5lOj4L66Sh+A2qPBIVf38cacNCnHRPTx7W5nNoiwD9M9G3uUWk
qRPeMfnr7d/pGVVivw1v11XXylMJ/+EhSS8ZyiMUcVAijk1PtPAg2qjcyVjt0cTx
qAyce/oN9s5rL5QcfZWM6N9LjeAwVpBx1a1p8v/Mv+LBdlUD9RkTWAMz1UuUr4xh
DC7TQ42RdupQJqy8Jg4Z4YkZOrDXDn2X12T0j17H+NDdo663botLihoBpVSnZK8R
LkNpNp0JKqfBY+74jgimC+HYmGr2ZM0c02Vkrpk74mdRX6uw3q/lF9/WjCr5l/in
GMpIc9lUS5FODINTJRNfklcZVRRLy+u/Wgq0Cqc4CbY7xgZ+DGkpgvT+t/IYAlmE
cajfI1sA77kd/ZOM1jtfngfFS4ag58Kdkiu71DJUbjL84cwV0pZaIxl3AY26JtZW
KHHs55i6gcoDo+XuI1lgFrFCrO40d/hLKM2E5UU69ys6E6KSWePtDfo0EIBixQyU
5/mhLtuDMber+nR1XtIhr26l4jyjJp2ddE5l2d+ndhc1EKmcgyAoiRLPu22jzaW7
l0EPffslhuL3e3/PU33s7yDPD3ykh6heB6wpqCW8jddVrp8mhv/nKgktQ6nanM89
ZOrA5EZ389UX4KwTAb82FAWVkGp56lhr+tsOOLuZ6lWWSaLPLvH/lkcVtOVrfTFx
LgbgAtVgN3uW1K+93qsJwgWfnpnSUzq8DeV10lDDpNeYbVoJCiOAnZzs7Gs2JDez
fezqtfufXBuKriuAbitDHEVAp9xO56WZXXSMHlvTsD/m0XqXngbaDauRaUEa8jys
y/xPYP6+9ayfC8YUOvhmNjBJnMqtgkgtKrE6tAC+X3FnAHvSoVzcjCmYQNQKXQiJ
MeCdrc4ZeU6zjey1O5xP9ZwT7oTuOSaRlENuIcEBxjTM002A46oRTs3Eku4y2dQQ
+XLI58mpiq7eidQjgzk7bJN1Mz33lvf6MQO2mHqjF+7H8evZJ+Rcc0sk6VJpN/E1
D5TjgNxR0eVjIB2K+hGGVZ7pRU9FAVp8FPb+cmNj89uvzHz79rsbRgPjiaJH/vpd
QTbmT5RzEU4Fi6WIziw6NipnOFg57iLlfrmALdxZ4dVJeONkMj7e6Yuaeb2SxOP2
hrgAdC/aMfMB4CzwEOj4wcAF0CCUUqzqWh33GiDv6nUu2cwbfz1VRZEkysxii/d2
eRp2nssIUZrsVk8Pa7jVumalRRZu3E0EZ7X1f5rx26xUdqebT9Bjh7qKKyrZSIDp
1doIl3emhVRsJA90mCDDoBUNsmgJusqly/Xjq+qkzrGi6q00Z3DwaIrGsbBM8d25
Fvm9i3yr6x5RpRvnCk+u6Zl7Urxcc6iX50vTtfGKk+DhCnQridUEFnCY0g672BNv
uykCNLRRFPfiygA0eEFLdbn5tNBfAwt/zUA43h8pC4rYfiy+G3spLR4zlDFgyI9V
Qp81OXNl5ZOkj4cwVfBBuBTYIopljb2wEr/+JtQHIDfT143R9wCePlrstZ2ilHWN
C0OMNcJgzLtG0UF2WeRj7soP3A9a8Sfdy/7YLpTD592PNO4KHPGeVcokIQNTSKaz
hXqHwXylJcUjH6BSCGDG3ObNNC8Y01tINmmLK+RerR5c9c22oYmKi8qWUj9X8fil
j4AXLVkMyOpJj2XCLs7qrvkY4mnaMwFNxHdMIbo60AHkJJ9KNNz+kFLmfXlft4Jn
fbv85PbBLqAYl9XDB4dX/Xvp4G2WLc6DIcsJZ1TYkIRAW98DS3BdDAKn8YHcwqr5
CpXJ2BhFqO9VgBmTRVkKtg/0syLq1QhrA2Ek+HdzUs+xu5fmAa5toOC5/mdRpVkL
8Tz2yhwANYmm7ZuLi4OXyGmUOBzubmi0d7gaSM9ST/ovpHOiHerF0BbfWzAKO76D
jHXy9qSoX56VE10Ya8+qKHjfDKveQ2+HBaXUsi7BHUa+m9QUV2+4SU+calMhEqXU
0jwFLWdO/fwSF9gES2+lZc1BZDqi7c6G/WQI1j3CCbRqx2EoqMBrYdfw/ex6s3M1
9eT3SrdNZAzH1KgOaMYtcpUDnGGQcl5fTW4biHTnmfpyvCqv16HV2bEBPxRC9qtD
cVESR6wKWKPQJKwmy0jk2EHnBQ4IJLJa2/8NfuTPa+zLyj5K/Rv1V9Q209mpjiJY
8d4f2PfvTXoXNQzHLydJNgr3Xie+c4lCOIKecMVO35UHlm8x1lVKy4yPW39ryNnH
LG+RJT3Q1/Wn5fDuzTX9RanMf+/HIEX8uPXmYUpJqWMyZ05qhmqbc0+4gTrEe3Oy
bJBpZGIRMAoidOxBsjVwrY45mkmCkTp/ASRxhucli3IYt9CzkdMbvs1uq7dx8Hrq
1AOgNttn6jL58sdlEnnZ8/nZ0TyBULFSDPUjuPlxbwlZNIrZYXzcXBJcb+VeB86E
LBlq8q1f/yTm8YjtKBkVU4GJyemHjD13N9zOExmQOyjC8D6+Ou0HbCKrdgWkVvgG
0MI/zP11cgHiUysrAiu6EkKKHkkE2Y5pg3eAb3VmbNy6vtiVvZz5DWrtgLzR+hD9
6AkQcfljTml3scMhD6Fp0WoXajwX4FlLs/VqPkYptJdiSS30feM7BA7ikELvz/Cf
4j7kyEGVpxc75i7UEB+kPxv+HwKZN4katK4/hSQP64fs5E2AJBYhODJ0QyadDIzZ
rq63lU3uk9VPFMkiuOrX0WE5geh+W6fJ+uOid89dHTO8s1/3TtVnQ5/jgDiBMT1G
2KecxzrJTiFMgJ/tKI6I00gG0ALoSjnZ1xlLLdzwgfqcAGANkHV78U0EIvBqX6Tk
66NyF6GlF3t7wATWoeYLmCeSpTEpoqLL/+BetcDBPSXjvn1S7h0oytOclSolAN+z
jXJCL2FaxN+iMGnz36Dou5SN5IZuxHK+N5ofax7Vvrgvjg/bEEi+U+/2tT3wyIGJ
B5dvb9QYVtgbxBv24g4OO3fPZx1rGf0PHALjDDl3dHPr43s5ZlGpJsIHedN3Hk4F
NIzDhVPH2n5GjqdM5ZoxoeZCzePBNEnKPmwffn1yj0qKs3IOFRrdkLdR00DPnPmq
374SgjyRf/JajFQHNPJs4LV8q/nbwdkecXXuiA7GPgVj6mojC4xkMnDoJMwsf4v4
j5AILSw2dWOwlOQz0+lZD3FYgqKyjbLGVcs73OsvK6a/IcW/bvvAF742BTfm2fQ+
34GqdM151AHrDGpZSTMnp0WesafhfntALEkYNz93HCnCeC6r+BDnpb8ZaWFM0Fzb
PsWdaweJSvuZ/pY1iMDPn9Xu+sAs/Y3iUu0DN2XYJ/2A+7zTHSMzpGf/0IukpKml
XPenE/BkGriov0+SUJMJBmBnP+Jqeg7ftx609KcAYS6+vYNA82xTy4e/h7nGEsQZ
6kdHlg0JvpQWin8XX14ttwBb/NW/oBCONwOq0hJFKh690vv+msRjwu1EFCz5rHxO
1Jcia+nkSBtcl2hYdpGeDIINTGI8gVlKJ2097dWMIAtW6qAFTmWWCreMajuv/j1/
Nt0OGOXDTZdHQJWtvqb7srPLl2W+mJ9rOrrIDSD4+c7nLRBFS4O6tAY6lHOYo6z3
g6OAUW0kajA8S7pUja3GJJz2xBiJ2mNh/Gi0ryW/FuwUfCu26NDuCUbjypzxJFBc
k339lfzfBB5s6ImdqN52F3TTDRjF1ONPf1d5ul4ccEYBtMgoDUdytmzIiZEw/hIQ
CqSx/3qErRmiN6jSd6VTxKch7a3QZXIh04yvKowTPCwCw48JxHTvtLJM7a3QCo6N
JsyIPe4xpnzgWHO/xG0QZi59WOlN1BnPMoXPQI0QgQT+4gELV/Pv8N3PlkiNEkh8
HCrqykC92rXXCeW6IM39QhbR5BRQEehehIYwmvaUcBySG/iGAdrMx5kqf8wnV3oZ
pXqoQlLrK5scn8moufmI+ucIKgH9p0jVTx8tjIrCi5TlvfWVrY7b7ENir+ghNevE
rCDxaNY49ayHOMcJavGaZoq9Wdk6NGXfFHCjIuGepBgmIakyrtFOtLOYrdbuA+qR
d348+yEgZS52VAFG9aA91KO4GYrXUW6kStBpLFf38h6xGiRCwD/49wWCdVS3Tvh1
eX5HK4TocyFfjZkfVsOYDfbmpRNIojqCprOI8Rk45N0J6Lw45rzb7aTUF293gUMr
oTtwfAI+ceXcxlmK4tqWvcG2d5zQZfatsoWARZmYyr5Ww5WrH3N+NNe+VIFb60Wn
fBUi0ryUnjypajn+iisQarBu+TBZAkYQ7WqwexqiDeP+pVCF6JcPliTAZCAm8kc9
a5MbKhDc/tMDC72PUyqCUN9xoXbM9tz0zIRPrtIjUXRWZ9BoEQMxdL2GxPnyfDdw
2N9ZnT53fjLnqDHUnmp5MHfh/cCCb56jiZ9TT+oML9wVmafRlkNXp26/OA+fEF5b
apWj2yhPesspuDBlS9Z21N2Ottj64wq2DBNVkzUJWGYwmV4acn5XnZJ9w2ttU1eh
a6TockP0u9LMPBPbDUDMg23geLCljr6UtnAyqAgrNGgcNct3OYg2Y4QiirMW8Su9
jryDjYXQs355s59hyWqqmuaFZxbFv5x60ugNbOS2UcrnnGPU4fWOMk4s8o0kzpfA
lrHuRcVPlM2dL1WqydJJVh7nyP4e5H+TLhDrH0qP/xBCzbwmzmtqhbMwtMVOXlKL
Kz1guIH9CV2IwM9JDXHEndc7qAYC9JX5lQYB2+NdjIEqsfS3RZKKZbExJZPUQDVt
Axnk11RH270tszX9IN93SR/a7oFVgwWS3/A6O2eWdoATrwXnsFDYi4a7iguRMWeg
ynAGNErQlcg5/afmbcukJpJZybPpOfRtFFNw1jl+l7D2tW8Tu70yyoj2xrmz2JQw
+J+jJa8MGP6MuUeCyuPuIqDzeq3GaiP8epQhOXggTu4wSLEsDn8a1Xz/z/EL6Fps
p8O4ch/UvGRti/5LLt6kOGx1O6erv+/+IfEyhBSD0VYUVvYfSHxFe6LFemWfiZ8t
rPD7mZ7MC4ZysgjcwgywbX49ZdxjCPfmVA6t4jOphu2xsFTufi2vcQfW8mjvh1PA
G3nE00XYb1hWaD+m0RJBNa49hRzD5MCK6XXD+PqPiQyqRnTl08JUwz0estp+HCKW
KpVTYCPYyo9B99lJxrUHZj/Gb9m6dcBZIidxLRuvhDVHV9m3quMWI3eQzZLWn0tz
RjEu18qMtmFyJuZLTCk4RaJPf4jJ4I9CVVpFNMXAVwMeEhVFryWbvVD7KPHdDn9W
Vgc4BO6Oil/A/IP0EDKVo4r1/SB9LZQBOtnKHf14Q3zAPC4O4kJjXrysg6yo10Zu
JZ7pQbz1mZ7CvUs+zwNKeM6xlEJd95Jx7L1aJzbTFoLMdpAAVyoQf+rRowabXUoi
9tvisZYsY+sjebeiye2bn/G4X38wGgvSCE2JM9rZRGsFQ6HqsliGb5L6ecBLD222
hYuMBBZj41YSuD4u2LoR6cXrgbdsczpvri+8CHmz/7uBSELTTDxQUt0KfVvWe+aV
P4vh7h5MEeRxa5nqoQ3HWBRSAf3x4Pf9F8eV3FdWYBvl4VzEY/5EOSD5IordyseX
nICH7VR9oOG1X5rYVS/m9sqn5aZEmH+6zwh502KTQljyFVKrKBbnUHRT6iPWoBHG
QG7n5yRloBtoz0D2RW7+rmuuGwdTBC7KGFaJCiOgQAUqq0CCky8mpb9Yau6c5BOp
IWAQOjgh2v6noR++Xk7RPsIUVms5eogMtpZyIKAx8TJSNfx/HwaC1DSB5tUlue8u
/JLoLuDrdywIm1Gr2o6VFge1DQtJyh6JTNvMPTVzPLpgZpMN3b86BKQyDBn2EmMj
oA6SsWpJW3fcwfz5OBfPgebvnXZdpMbRI3j2i4SsXtOE7WA1sgJzI6NCXqrDtmtT
EPslCsVtrKV2JmpIizSZJrgTNfT8gB1ibwCYqenRqiakQ2qr1+1IT025hVEjsnph
KFJjzjX/fVVEY2GnGSQiqquKvBNh1hCUCrhVaC5Bg5HeFYztLh2xT83E13vfGH/d
efaBAI3urLY5YN91N1qREav67cUKFVxvrzBIJD9BicIWlSuZGfOFZr+ioa1L5Qwk
FAiu0BQphZqbFK7S403SZw/nuufBQ4JKpEpmoxQGB6zsiTIiOPi3bJ9JHX+SnygS
P1FZFY+7/S27OGRe/2epDoo7RPnJ0x9kIDY1zND3QC5NFSnxpjJqX0CiW4nKQOOv
/4rCtu4d/bs2tPNL63R6zcnuPm8miwQ30PH2E0qmx2fB5udjAhN5mz6GNhQK9ZRx
QWbVkTC/runUzeBq7G3Zbm9BdEZO/k9mzwci9maJmw5h3AEH9Hl92eE9e/0bt8La
vwNrYh89QPvxaGi8cXzWNjwd5OI6UDeFwy9FTxzspj7SdaWCsIGTC+RV0zBXIXpR
9bC8yAQixYJOgzQUz4mOMA5Z+Gpp6J7ON9/+C6hFNcBNxD/lr6MuAhQPk3jUtA2n
guSA9dwH0VUxU/yI001D3GXRyFMxu8bmptBK9q7hvbzWP2fuKRztmnTnLqxSokBF
ytnTeXf1SP1kvGcKuQETu39J9PCioS+Ekj+TidN5uOTicadwFWGXaQ7PjiOP7odh
BedPjvIYAQ4I9nGSExbVbDyPIh5/reyw/SA8jQ0rNH6inQwsGf9zWNN2li28oy+X
O0Xczoq3ntZKbx55I9epIbfKfUDJGf/X6xDfxIHdJMw56/NSyh3+N0qz4MozKOOm
XkHrahEcnkCkzjYrkSW3Wwk8mlvdYafd91n5Pm7ShFUHi8pDopTfIgsPq5273DJG
N6e6ITVkFg5oPpPyQFMtlfxwABOAcHxndpX4KdlCtREuMXsJ16FfWMgBMT144znI
0kjRT2ZrA7E8K70KSy/XMxn1GrK2fNUPJfFXoZEEoRrj3mG5EJ3+XxvvI/3EupfB
x34tNQnbp6XyDHvxPdrz+EyuiZ/o9h5hyyN63yw3yQr8QMvJgg7hJ2Zoxec1k0Dc
Ck27uav+T8k/qGAUSKjFMhtG6lWcGZCIzXezyVZyFTFTUAhHYa0voxyUgEV4jLlt
YYX0BBrmki6HDTqVfs4MhNWB93Wv6J+nchwqsNsHfjvyj+7EM8rSJoyiy06epePB
TaTBe3cQ2I2NADgYlEzFslkyJ7N1hrhaGJneWGUMAXR+lRKztLv0CG2wml3W9gv8
VDmXbaM4lFT3zSfP1IX8LXqxKje7WJlNiiKEMI5KmFU468mCK6/hjz+5rGXoKP1I
JfCySPvgiaAszX12XkzoJGqNHCBxCwx58y+kUkIgBTCdWnq1absn9/3mE6i9+S9o
yPUSdpuTa0/0xxmmXvoG/ZBb4fY0XjcB6koC/EVFeGPJpjru0XJF4clvA1TmRSoo
8NckW3R90dfIgUhUbdU1NhVHCPoZPjjDamsBeCxMrGKZ8SpsCSi3FVFroCEoy0VB
VcD4lst/WL/kZP1Kin1AlpXA+5AaS23PH6P9UKceFmITO7H2GxodUYBC9os5rlJM
tJNxJQMfrZgLm8o900fgRGZIVY8Vmqh2dIcEK26z4QyqRYtxjjRbdANmcEsepxV1
EMFMU1dqXZG3y9Hs0gx2DEXCYG8nUOB84LKocG9zUELkn2seYdxb2CylwdfnfGLH
acV/f++oM9fthm+mKBqjV3mjTKfNVaU7LJocylfSYDBpYX7a8XEbUgL4208Ydx6Z
D8kYdqadqi2AvIHBl1Annf+e7JhlRkTEcB96LUdGiVKw9mx5tMIqyS05hoivVWGC
HI7PGkNgZ4ZD3HtgxznWL2FIDVf6iiz6PHlxmGxVkAcBX8ngnHWMKaVUaBzEcycR
sNUdGloReRDmG9/FEbzbqm+BsTILoYIiezgeSKc5DLixllJn3k3SAV9thLV+XuVR
p/ky4wzvbakJwYcqx4S/OBD9e6EoL8KUXpBSzevhjg6fj3kTUuohmcN1F6Rqe7MT
NXLnTj787XUEVns8L2cfoYTriucB4wjMQKyEzfZAx0tEe95DRlYc/SfmtsFOIOfd
KmNiwuuw81HxnBYqmwYPjukgLcbAPugcq45/pScOcpnwBlnxBEUHgJEt9H6Gmo0/
mMH/q+RdfZcWFpEfKq4V7YW5NFax8uUr1LXbb8Qa20ti1UXixoEXQb5maxmuhH32
c10pY2fsfoXTgVIWaohxNS60cnhF0wsUHMHyIifDphOG2NSxFWKHIhZLWkOp/s5/
NgPm3xMcuXCfLCO+Kta1G/CYW/kugE+JsP0p35OCS2oHb5u4tJPjsFOwh5JqNxhE
ltNELrowWS9v7mHjs32jOz3g4ajMJ6gsKKtin4kHb4HSWDTGKfHm8duTIaXg+C+U
+Vb4LaTO7ZMeFb/SJMAycsuA5Vop1a7ijfXrZXZrBMhVkN2eILmT1Rp3GGQl5FuZ
XlIFJ+9DEVV6FCyXDOqJD7OBiGymsrdRfXFfUPKCLZ6vkFKqg4vtCjbaPly2CsxJ
cpvuz7jR43RDTNTom8bvqjc7wSfLEtlVhyhyACrCxNv4k/x6wh1sk69HbWfM8nZ9
edemDtLU+aJCZoHg20Uopn4zrEFWZaO+w1u8XQQYJxVwcEgu44rLk+jVepbLaeXo
uzId0U+PTfQNaHiv1QGbp1x0kKRlh5OCDxm2cDGKwgoZxexaiUCcXnhzkifc1nYS
qlrHNex7Is58ImljtVd6Ncj2xwsFhNECMIO1TiI7kHe5uQpp57psSiXX62PT6fsZ
h+bkZ3kLJ5vdS4C10u7tbKFJndaP2ryPRoVsmViEpy4S9e8zvor4TgpfQXpQ68l/
zOhLeQQ20j7n2SmHr1+iLIzLlMHmxNwrf2YZ2aAbT09nelSdnilXabQPRK2jgDFw
iTvoQM/x6hemXPoXuWKnwZFa+pQRrhxWm0tFgOpFOftLDefN+xXd9yNjuh7AxhRa
G/Q1NgSJhCCxXLGtiB7pN5nxg2AVEGdi/2Nr6847StEhG7UH0cuwL96frht9Lof+
6QJCK0NL8w+1y6YeVPKjqn+uFYh7Xlt+0oC3LXt9rskYZVuTb3Y61Dl/kC2egEAa
YubRedxoHBt6Okbmo5yJWAVym5WPvvuAUSNKsqY+QQSbQwskNiyjQEnsBmh3soDQ
Qh5IfpeUH6uXppsTNb35/V139FQwLccp6Ttl4UbDVPNRL12NB5M41vBDjjhe0oog
ZpbhpOr1GFetPQcVT9lqgwfD+aoTJzCYSi5i5pvZ91SNaDHtFuKMcITIYhRkJgt0
NnsRRgDVqcSW279PA+ZNSobqd+oA85OFSxQblHeVXJdcnqc4AqpMekxhIsgBG5B6
NBpx7Kn1cJV0eocp+8EjpDGOT/vAGToomfMhKmLnGkDjNtnm4gChmUtgP/UOsppz
Q6dSzbUH7KWqwIsHP8oHa5xGC5braiu7nQLgi9oLb/QsEyZ0HoGNdnvJ6PTsNPyC
zdirwgNDDJZibQ7QRyBgjn9TTnp2yjWtXkXCQhcXDa2d9d5dhJ7VZ1iqZAwdUiPi
HpA37NaRdHoWIDv4RV0GepNDGkWSjC9PKUsoJZIOM5XGdrcWiLyEoh9Jb50LKvU9
L/HwLOsAB/KcQ17B9uOwOq3ZWOCgsp40XT5dVjDPQ7PRpijkwWswKage4dbgleH/
51y5EZggv2+A5b1nZ22P8XhuSDyQ1rJmSoaabcwQu0USr7BFR6dJc69912QLgtyk
ud+0PQDI5YhaI7SGA6XlsGgWnLUYiDLHYOk1Z1ggq+SeTji+N+thN6NjIePXu6w6
sQcv7IRgXxvqrjQN4qAGmRxTxQL9T6YFKYFXIg7RTAcnPOem7PYGilkBzTL73eMr
2qfm/xm2Q9i1xP6d1GxwwToaJwDKK7kH1Jj3NkkWUrgjn2/tnchsMQlMT283eQRx
YU+s1TzvH2WOrDGTajo5IBbKwK3egYAn2f9wRqQoqbKS0xDA5P/sz9NoWZyKrEwn
RzIa1zg/xZP4sB3kdGknm+ZmMmyt6C5YcZo9NtzeffTvxkqFyfWPCvDkRCswaZqq
oFt4vCeejgGNswOGAiyzdfOSxV3pezoWkqmkpRzNZo0Ua7EQZZcxw5kkAtsjYVWk
RiSiurtdEtKRJP44ZDNgUf2BpicMHPWvDwuFd0hzJG/++IZFs/EpddBB/DEv+EtO
H52VgP38L+rHvdPmrtH3ErOEHB1bqkJ33rxZ/uM+fwhZlrYPGwBKsZgvQ0v48FHw
84x+5OC35jiJwcNJh8dOzqmD1BCajhE1YvXTKefXP839MJIt5QO9oJRFNuHnST1c
28Wi+ROPPc+KTojqzKU3dObkp8PJ4ZJ4d/LH7PpzawR+YRwzy07gsEnaBNT7GOV6
QrMBrXwTiJAzNKvPDfn8KFMCQzgG6aQm9O1bRfSTTTxoJmfcCCjLSA2GXOCMb4ui
zf/Zvq3AT8GsvCsGGPJw+8HYqc66iY3afpCNpKrU+OqIDVcEH5UE+vR0sEQAubDu
Qn8rL0ibBe0ds92xbOzzk4yVGd5bDkx3x1zYVvqwjYLmGUYo8OQc0grw1Z33astl
0IQkdVtXZtm2wD09nkZ3zUDb152cAzE/oiZjaMXk2UYOdQ/VrC+/EHrn2P1XGLeW
vn9LYh0OnWLlNbx4/WRsiYsYXmm/8Ync4cjHKxVnbeB5f0q02RmUTwT/GoRpsxlb
FimTuur1BMlKrn/r6PPsbIlCfitc1RFWFNVXcln1MJVMUqZa5CjQuOto684I8c2e
j78jnVLla03+mfnfDgbaYcNOXtL6weXJf5MwbaImaz290nZn9mJLMxUmHfQmAyg1
ExFHBDvvWkkipCxMokRRH87hidQ8jXSmEKyCkf8KPVcrnSImGIxAbAuyfpx2MT+2
yh5OgOFsndpLgP5RQAknyOApsiMvelmLsbtsdd1n5P5UU+zyjablT6k9Sv47TzAt
pwp8Cp2AuhxdhQs8nHARsbyODbcmSB/kLfFSNMP7RbT7D8J82tG4U2PP03CLpILz
pCriaTJQj5meHs+Tv+kSkK9Iansw4VLij7K7qTK5uh0zub/9lDpyN84bdWtBMLAw
w6jzhUA4ma4E/b8ZEzF+Fne0QLOqj3qeJPkaY/8RfbEhBOpsjpQKUvRoSQKl6TjX
RYKESaA9uka31WIBGq5ejYXpIkZmZnb8t9pxdbjripTCq7mVRUXYwJdzBGzdtl3p
/KTQO6C2MpWMd7ua2CD88Zd2PmFJw1f7Cy2H8H3Jxq9yggeAH38gS17ej6CuktFT
vwAeE/07+doN4o8P55baAOYfaU6bLAq+qMEFF8hA8dixGAPj9wVs4GhVglqQH/py
IaCS7SgKpb5hDUrXuNJkMWw8evYhgj4rbC//t5hcLPjokc5pNdglqy4tu6bkAK63
L9dI7+sb9TjlP5iySFDygP+qz2TYEJb3LwSGqTMeSjEwg2UMJ+W/PKrydKUWRD/s
N9qQIzhUTBwafYFSAjKNvwEhGklzyR6M5SMO2mPE+mrGQ7uPc79ZFx3cSqXR+tou
UzREvnbuwwsGlI1TKzXZEFyyxTEjej0gK4Mtgt7V/yuDoGH+KPDRbEnL3HXvxN5b
LgbskXiCRLT3Gkkn1gz97NoaoG/rhx7emb2Bb/5EdInC3LT54IXDwSNc3o+6oVNc
09WGeSwnT99lKlT/8kw/LJRq6LdQsbzdLubY1FTl3YUHLMQHrw25WW7drmYXa2GH
ko6FLcTOnOV/GRJ5/rS+5iaWQ50IuFTeiFHmigh7GZFmfRpW50RV5HFVTGf65BFW
zNaKjSOpg+pKwRtO7IYHC30UD8OJ4PeibexlbUS+jGdZhAIcsVSfu7PLvsjPdEE5
lahkzxnbxupYrz8OrUYnqNV5tSE7MCFN6W6Ba3qAXqEjU4KU3my1z43EmgPokQez
9Gwm6ZmFrBxH2MowbH6gEow0u28gBnXieJkkrJuHr9xv7jQmiCw5oAzBWfnYaqiT
0lLoTXTEf6lesxyZ1pLrE/W0t8VftAXjq1LPwrZedFxtC+dHomoz1vZHUd1ab0oi
4kR+bTEhgHsW9wdfnAauUK40392q/dV4v7sDPsfHQPHcBsyoffS4xcpTn0AHA0K6
dW8NZew0sTlUR/pX2aMWlA+zyL9Nr93dSnhJ248XtmfE3rHrNpyV3eJ4tNfe4H1c
U0XwC85wtAJZMjScO9F6JXpU55zxu0kGiEB2uJQq+0f9iVg3ad+uz9NhjhIHHJC6
vOVFxoCis5zSy8WwBGOCBPsqNrdE0Q2iyN6YJbjq8VJDqA+wNiQJjycd9RqT9AZH
yvtmYBYB3MwUTJCrfs6lJDK7UJEFPdUmPA7YyLy6f/BB0abcbo/x3qchmgSpLtu5
4/TmkIP0+ng76uwNBZMYC2f8xiQfN+QB55/s7Q8D8nfprbMrA3/tA2rm8CUA6jxD
Jkabg82IuceSQoE3CTRq36Tz79BPOQREujyIAhRGzkt2Arnc/WaqxK0ryVkhMZja
ySZDtz7m25p7A2k/lhD77J5UlSNwyrHoCUYjWYAKrAoJLqKe92TGr3VavwzpOJtJ
LXQxStoorUi4p7YoK2T+aaOQBVNsoykxeQQv+wuGREJDG1lNgYVVrAKl2ETo3t2K
yfd7oDUMdOObUL+tJcYkMJcwO9xJG9eE9YJlrVcSB8Gv3i3ZH51iMYdy98vF+fk5
faDlz/gNlFCSlQG9xNdJrJ3AnSYKKEvX3E4rb/9OeVSi9WZrZGkVssnweehVZWkJ
BhkxeBz4+y9tPDa8CC6BRHehVJ0uBZ2UEFQ1foBRamg25dwIOVwYKmbtwVk4lqhS
Fksmy7e2ZSJBIjNFAtVnFO3gYVnYc7Hlv0ZWEw7N6zyYwnptjRxi1BZGOvDs50I8
5jsF+w0yukTpDClER4IRs0W1SQs3KUrvB58vVXyQU7rLWs+AM1w68b6vQOJ47oV9
DD7JarADw/Frq3aadPc9MykFrkfdSZ6nBak0qO4xxecpblXkq1YI4/dHMfXOHyoS
+Hmu1qDZsY4VLqtDfSl7qDMV8prMjFt8IC225bVhBU79vetoRLjRaCHJB1o+x34k
QrboWhWpVFGzMxkd0XaNwcQy4eecUxuCcQQxLpWeAQuTQv/dicgPJIyRJfdu/bBn
QEXXGji805gnkLOWFmGBxxPFde+z2iSXbpX60ncnnYv3U+GiQK++H11i/Cflcjge
hWVtYs9Wmw2ZL85O+8uucEjwGdiqVrWlmrtk+NQy7QoTv6Dz5Xm+sKU7FRcwPKUX
g/rJ3wDDS+lUrTBf9BwIFyD4aOTEDUdv0uSBdQ+wjCE531ivff2lFclyuA6b8S34
bu4Bi7rn0HsWzLK4D/BCouSvyqn2kIdc/eYyrfZJQsNIPkO5LFGniVMzjSoL+fvi
IlFlwCmHCwtrXnyUGJsmYswqDpuTa423+o4siDcuWW890TgOIFHke6ddb3WICun5
kUmfmYzQoxTxuBZ9b9/fYliCHaOLMjRHrpq83fHE00k8fRb9/pwLV/YD4gvAKsO4
pPhRyjKOwUcbAAF7l+V/S9/oYwOzpMcI28G97q5OlsHaLf/fckpXvT87dWFmaTTf
zszH2FKhBPE9oip0/LV3ZXF5aT8bsZE2qZQUqaS8walrLu+BoUlh/uyvjmp9gncl
ozmAvz2D3qO/dWSd375FpLbnj/5z1OGfF4Lip4euxFhjGfSlq5GCkmrMBr8sGqY5
wFD3jVu2SHTxilwZTJ67u+9O7v/R4Bi2Adesdz6MFHhpx0Fj4kj/Wv8iKdW7BEYN
0tt1hK+mynw/Ulsi/WoWU7KbCnj8oQNkhnsdCIxSh7G7VG1zSt6FN+X7DriZ6RGu
YTpL7GKz5mKAQyvPnBiOqVeL9L3Py+XZn4lUpMPbIkNbJ7mPCn5v1werZJuf5L3I
gMtzEDujiFSg/AX81SlJboUit3RX06/mqIViQW45jhr9X5mPpgVJYuSnI0TZnfKX
PiQEoF1cp3J9V1Q9GIooAeaGGdtkwIibmv9gLx7KuCGpzgasIR1gDY8EuhFFjzjC
4/G+HdzLSWCC11CrQvYCKPizUx3a73Nor/3b4+Ea/USwjfVOyH7/IvyDI0FY7Zz0
KS/fOqjHqPhp0/lh/q1CbGuJ+cyMPDxAUKD0ZnrWqoqA+zAxx+cXx0A/DIryTc0e
hVDrv5cdvemc7vaXVHHptUfpNc1a8n0FYfSywuiGDbSkNttOlyw7qV7fD6NSrPLY
juPiP2aTpybskTyY11RsFgI4Z9FCAbMU6nnejLBXcZOAJmBNF878tjG5DZ+3zKFY
wTiUhVt/pw17MRivH4vOJDD0ZaS6ZK6nIpuN+ckM6DNXuUL4cMEQit1bUHom2SKW
TecJVCU4Wr2zcmXNZ+cemcFD9LkzwAMVCZ12qmhxDdJqoHa14zeqh5fA7Ztj7Lga
NDkN/eCaP5AJQRHNVqsXbIafiZOSZj6ZSqHqLBYjrdbwfTMFLp5NFgFxZSXEjnI9
Frz0S4nxIVlNRU1YKvrM80v1gZmRgEPtu5X1VEkrwARGFnIyMHlg1Pn+0ZWTHuJb
vhLGP6WoVpmlNYJvHUcrxO9txbgoilRaSoyFNsBNjjqeeJJF5lixPjEwMKjL6K13
U85vEdUA/6SpbnmZi0whUU1k5kLSPXUIbgQfZHCzGiEuMDk/j4TAg4Qz9kiKU8IC
XKejchS/HFtRo5688UufFmwyCjXYEg1+edtmJwEHnaxYGGZ2oBho9sUr+veSmlsK
ws1ept/rSK6G0gqaYmWFmgZsDe1TFLhmkpbolRx7WBc6yFqrRUS+N0qC8+t6HRoQ
i2gArwTWAyxIcF/UAfKtvOTreh5XW3lTzOsQYIcLPYNncNM7n7qKfztaoZ2Lv58P
8+WjdsIP6JhfJsbpLogkYVjTr2o/eqLQNVjqV5qtuOJMXvDDYKrt++j9TdX2rgv5
a5ztpB1WVmdkH/3QqYmP4QF5qKpYFpM+8Z7lZBNbBaiCq/+F4X9QxLCUG7eqcOFB
TnY/02hk5EsShxnIOsJNbqtEgO+zn4A5i1Bp7Al/9D60KXTFS68Bp1o+WPs1V6D5
Rooh+7wYyIRq6pK88ZIAfO39pNYOF+3ow0mYKCvMhFTi38nlGeJIJSC0sW04ayAX
9AFaPLokd95aiSDHLnEvT3wdUjTChNeZ+z7XLnlmNufUJcox75a8daaTHbB0XsHB
HN3B1lAlR5acmC7bmANmf4KmA4d73j0D8zqPx8mYGFfk/svy2WeJs5hotVxLWvfa
9CMa+Ii+Ij7EksvrsMhHGf0OuAyDfErhRp5CHpcWWmt1jEbguZhcSKhEE0R5sgdE
32TOnQ947wPxK2xybpxE6fvKwy5hQvouTiYcWPc1Xw5PdqFdqfrtcX3Ksovw2YKJ
/2Smv2FmuJHnfMMCJZ3x/ETxqiPGKChpzgVDIBRDEXSOOCxE/Vm4fwNWMMkSmDZt
gXlEhWzlq8rrRNsslyO8SqoEtmKKu5qYnkyGQoK7goWw2yHOTKZqyKuePlpqxYIg
CNoz+Z7fn4y1gFSvdqlsOA+NF2XGSbMeY0CjGqDuRMjRNzFtOjSBcVf0DHioyiGh
A7Z6lTU0eI2d36uIkDAtonhUaPYTCz89CEsz8jbGHN0bD/zvb4/N8LQ7Uectmn6B
OXZe2MdKhxrvyxEt2OTnSxqgb1Tt7rZQK1ijqbhjAPAeWOEQYyul8mslCec2/KRm
+rKiBdBdgBHL1ANsyhSqU7mogEuKS9sqog7YcCNBBU71Z9ycOtaa5FEd1T2A+Opb
0vF8bFy8wW8efuisMGx+2XNSTkyCuZRJ6s0DVwrPFT54cfbYJGd1D2Fg9EhzIEML
RGBt5DPy2pEohX2t9RCWiLIscdgz2Pb6iKMe6tHvdO0JKmDHl3QElqI4vk06BWwH
AK7ZuovngdNzZUz7kPH59FHr9cJgdCXd9fyMLtEk2NpI84N7uwv3mOQhwgTL1yDh
6HJFXbgPLxz4ggw8QOL8G+M6KyK+CDqUV2FTmPzDGf5u5736XFfoPcSYAmlCbCLq
+cU92B12Fzb570IsirwqdfCGAs9HvFEEsnyuAhIuBbd2SkEl97iqMvROANk80D+G
/icQ1ARvX9n9wcpLe1vvOrdhAPcdSzvBhBZVpsVDvpaX+pDErnyB3Y7dfGlyUHw9
cBgRblYXHZOZGVM8mEqLfWfBKeVXBMM6mUgHsw34x0uOHyD1AYpej8BHHmQHOjk9
TVpeH3zqh6u/UVpIL/QWsYw08KFHeG5cr5jfrpS+82musRH0Y9iZsvC8qYJ1M+3d
BGu+x+JE6iIYLYg8zAKaWnXBTUa8xuB+hWtBd+rsxjWIzPv2s1ABi3r6+IuGys48
Rd6t+B6nnqMLh+6kbIRkpKkmDsIP3fSDcq68Be3gID1qAxsVoN6u5RpW+hlvT1rO
ykDHc8QfVtDg3Ay09AqPwcpFhkd879GXDGEHLoRDMR3kFSwHDMLaMIVxmss1fhos
xV3Lf2kwagfD28+jsum7DcBawCudfMht/UpiB7l7DYud0fjjmThFILH0kTwpiGum
b1W+lj+qMfzKEHrcXn2Xe+KyaqFj7lmfyib4q4R/8uFFalaDBCp20WXoLq5gKL3+
Ewjk3K0OX//QzlzY//TP0eY3a4Q4EB/hYb7bFG4Mzx12kHfpectfjoBxL56o29lI
VS82v55XWvCQNSH6NAs3on5Mqnzg95YRe1V/Od5ShPSlztxB5L4ndxz7YwJM7C94
suK89lyrAF4bLMUJXk3fsqk/sW62DuDToGlkRN4yxbNTMOd8FK+XbqDtQ1MlzSxw
ZS059xQecPcfSLQX9NoXg9sEJMak3yJMM7gjQFwNDRe3FmcAB7txYxzd+XDcTwL0
T3ZnQ92gQWpUGsDn5xzKsJDLrNl4EsasqmQyQXV7qPQFV3a0gAhdOSKqFXohNPy8
c1F7/MUiZO2+t4YEXHVCkgKK070z3p3si8VKPwa189wEbhJ58Dk5TxSb0+Fr+Z88
f+PJWkZIZzj1nMsVNdO7pWTAKqYL6yMmkX4UWFN72L6g3qR8cVWO82ESREUNl6AY
S3YPh17GGMWWzxIFtLYTVjLJjTrWh1OVIDwKUwYyJ6HqyVHINwF1S9ZujHqIJcyQ
T5YFyJXRXdVFIm7L8FnFk9aTPIKR/9nTQhpE4stmOvzT4Q0SMb9kbe9UYtt6mdA5
mui5KlqxEHQAb4ztJQpECnK+x6iUM4mnEiHOFAwB6f198NiyepZvpm/y8FoNuYSB
t8avaTxUMXsTpqFLfTEpvzSh7fkxyOcu/H0CDXTJACru0bicITeixnzZTvTdPo1N
K5Mwx6ZPR4JYud4T/hyt1AocfAFDfYJ71ZIEuTY6+/lEoQZzZvNX1rfPV0zJA+4f
y1jgDv3uMBcHMH9TUOC5g27mKoBzgz/tzpOARCLR9wWz2gVHcgXippqB/7EA6Gdd
oAt+YzUDZ7taH30+gv2Gm/BxOZZ68TDSWyBo7gNkilmLO2XAFiiVF71nBHCzvLiU
/OYpyC0EbHW5UBEOjQai6U8YR4oh06xGO6RiaRnuDASE0jCN7d+gu2fTtNtND2ty
2fD5P7uXi99Cvkr85s6nxcMtUgAZVNuTk74GROwXmdpW0JmwYLYlejVS41WHhP8N
0zipWCzU6ihSXQkX4TZJ1OXPqBizqd0Sie4dFUODVoeaCax8r/vTLqRR+R6g03R+
3tH+B/VdPnHF8m59fTZfLYKL+xfBQTMXlJqlLk0IbX8=
`pragma protect end_protected
