// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ha/Nk6lZxm34dp4BxjWjXQJPqQ6tMkZ9urpjjgp86syNewb/Spf7stcLa3+O5Xl7
rF72M0EQnlB5OzX/8jaB5H+R7LDYS2/MT3tMWw6j8Z7AHVk2aW0bPXRJw96R5Rsh
y1Q3rANttLNas1qNYE3VBjLtWHpWx/HR6fY1iL4F5+Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10320)
XK998GLR9aEgkPwB37M2QCEVVDo7IqJ8axLd5bwHnFP0VMSJe5tP9wrCRna2ZAFK
GORGiRTjgVtM80qgOveOQRQjpzAlPpLjn9m6wxkv7qy4ENJGr3yJMoRflX5s7Paz
oTZGfSIIFYUSOVqa7D3K/NTiqWQsyds4A8wfZGxu8+26jJYK9Jhx5gZt21mnXJaz
J0wBZ1cIESVuidGji6fCYjEvO8YuvglF1j5vqxKQ6F+JRBBG+XqMydsH/DnvtGCi
gvdDvJhcGwwv5bEM8KqgyFQl06d++UvcAJozaN4F1owXFPD5ZKFBQLMcbBg1yTjT
zza7zXPnAUTl8HDFQlZgXW5/eWqiprlcgyZAhwmGiKkn6e3ltPAvwdHNBR4jZDTf
NCuDsf8OpE5QhSP2LEt8LXrJXxZWcxyGxAVXkQdzI4JEfE9iAypIcuvae0sZ5dZN
8xgn4rm3iDL/1ONoQAvinPg2goZzePJLi9xIOI5cMv80rpPYgXpnA6t0OZf2OVta
b8a/S7ASVfyHDsjXdDhlSMAuszO58MzYimFtulli6hMiyrM/jne3+aw0QwuZAW/C
vx9zOv5Mec3AvdjMsaogr6vxsdPINemsGiVFQudmPDA7/whfNadhDofXswCKSicw
cLwWF1kulCeWywDBDLucxgG7Coe7cCTDkVGil8FTS75HI81kNLUo08mT0LxF1Odx
TLZ70oqPQsIp4jUHABcF71zPWOfh9hyJT21tMy98J2ALiqLJGFPHr6a++uWqWOuq
aze09jCAuhNehxVlcFxDcTIIJGzQHfW/KG53OtZ1gRdyn7r53h6rQ0k7MBepEekG
srGp/hLsYmJy8tco1arrEP9Kf0Eo1SnNIQrZilAN1MrGx1jTL5j+pBCufKDzv+MK
CIN0rIw7PHv2BPm/kPHiu2ipRF7FTxv8OnoAS8eVmwQwcEZ5qEIDOZC7qyl+86GJ
5YBjK+vQJSD8tjFZXPToQ2YJ0N7pEEP6T1gxutZf5+fDnSN7Zc2OQ7WE8sBBdmdr
GhyAJYHaRizzPnoV0yno98tjWtIfzxuy5nDwbS1mA7Vn28fge2PMscfw6waaq2HC
ISJC2Kr3hEKCsRGMFsSDOWwKVL14uH5F8CYtsxT9PhIaHkwbCUuofXPVSEIsYQnQ
z8BrTNtWfUnh6W+IaBCa6S3+x/zlOKM+8qCsPT9m/UknqDGAa63G8QFjAKiygIs6
mN/3//l2a6id5jDHhAHFWKJLatC2Iuzdwcc1rjh9R4qf3Tp3sP2WS9TZW/oZlL7H
i/mFmqTsdzUZVsFUfkpVGRFDUrKzFja3hbmytPApU3fELygzK3l83Uf5b7X8cKdJ
YIoSKBe9WSfLX99isUC/CYmnXIh/VgUxoh50SXhfilcG8iW3dE1TSTP6pEeYgfZG
4TKIsjsX9HzTInEfFOlQ9iyDkk3XH9HSvxw6DuWBBn1nJnsctvjF8mhglspDOA1G
wiu6qadD8XSekSGqw+DGsW6aGj9Jzw0RYsqFS7ToCKE+QaObitmCLrwCRRHU6Xvk
+ufmdSexIbYNXH+aZszEh3Q8JTgfWv3BwBbw3c5wG7L17zHPXUXVk4KSNmlTTnvB
2okKzpUwpMqWSFUls9uA8ANrAvyRm/IP6CocPc6Ut1nq61IyOrwngWNv6awZ3FX8
VrePmwkqIAY6NIrW9eTGAz+iqH265J43QVlqRzczaNb4MZD4/r34RJpCBGLpH+0P
jCfMAGbHpmRlp7c1vlte4qaeNx1B3B+izQVXzAmxKzmMPnrP2QM6iaDz5q4m5vgr
dUEq9FshgGNYkXvvPXCkDExSn/eP+wurG+zl/QV7DnfNZSf8y3ysMbv80CmrsuBM
8HAS/tpRXAAXFIeRe6fe32jPx6Qz806BdrTJHvBL6lKQhhXFrr4cDF2BCwXwXfzv
+vt398zDHWRAVuYBx1o8xmTCW0b2UwapmC1iH0gFT7kCzYnoVbxI0odgylB6eYPV
NVUp3FnhZH75F6y6CT0sSZZL533tZ4ABhB1ZOveYp1FKEDvpZVa7m+6ZeWNpBlOK
FlI7Srp5GPCP6e0H6b+m9pY/Kr43GgaU0K4Jb3FwGytbrLdS13B0IhfGzykNJWCz
HLeOF6RSMslfV2PW6pY+y1hebJha2Kld1hjbA5KgLTki1PVWQfWJ3Rt+hQIsEM+B
l0whtNxBhEfjOrWoRvD0nC27caWGOPUZgUzoE6OzZ2mnyKQe6rjA6vkXc+B9Cy1h
VZTc+9gXpuEFX4uuGb3XbeW1GcKdgnIsYoL04fNEaPgn5QrYoYm0UJ/97yMPFCDm
Qkc2PbX4AuBtmdSv3/Nb3a7tuItNmuBUBmQ7gTNLwTIK8GI0rsTxVtap7VqAkaAC
e893o/9HrgMxkyfITSLOYH5o2zx8NGaW8goTDQFEU+TtBu4KiCI7YcAcL06xYeJL
JAPTPeLD/AXA/nfFRGWXT14qaMe2VgX+FOEuIGGZi7hiC4TrxovmuszWy8bD7m58
Tt2HSIEuUYp+WotM0hC8sh/U+IUfUCKYXxjxWtde/lzq7bGYQHCEpsLOzLJ0+diz
nqbO8Y2TC37l4RALuq7V+O0gKv8EiWy0hAZDsNgXXEgvMOX+K9wl92SjBQ052tyi
oCCMrpa/l7VlP9JnkvRgOdenXDYfun/upza1IkrThRu+LfrqR3d5xGijmQbOlZAK
X6F0Tl7nDy7+ndg57751LpGbCxcHnfha7r/91coKTK5SdsgspDQOAfOjFQW0FIlY
6QVAjBEMeKQn/hXIy7SGdJtkMuB1EgePUg/f+t2CbEoao4JJTyJ+VC7jOtlcGZoN
JRyUD/RNbhWyK6n8+fUCMFtzg+2jrPVwkjaXzVM+UitowvqdWTDd+Qcf7gslbMq7
IBSvcX8N64KwbM+dYCzP0KdYa9Fgn/xYZw307qQOIc0voz8K6lslLmP+xLMl+8ow
9hPLvLX1I4kNuzZwtYOkCLe02ZKRC0P4JUEwogQk7kK2DAiDwayapbXSMPsBSreZ
aaTVoCiC4SHSzjBlzwuR9QK2qsg5CpomQVYDrh2cC9ccLbi+yvSTo738z+agpbbY
tglep921O36zX1Wcbwq87y2f2NHUHqbzxn13BqO/WsDzfRRnoFvbXWI3jZ/nlLUa
mn1/Jo2T5uWjtZtLmmhp0FiYa/9BO6ipfntzaEZ8ClsFrGdrH+V9ghjDhzWvDG9m
YdnM0/HbR59XdVXjdYJW2fksTfsNkplVdFYWH64fno3KhZ9u5MdlfYCVyJTTPUzz
kqTsfgSWFfa1OZxdAIWb1jLhXDHOHkw9VFDjoE+X716CzPWDo+3ETotOSyteD12q
s0Lhnme8niR61GdhUbaamKb4KXReXMBFq2UGhg11o2PPvwqjon6AeER9M56EwzTz
EW0vM4amkIqOIZggTcRUBlopC0mqwRR4Eb3O4ifw+hrKxNmp4XK1/xl6zU0eMRD2
S8tXrNpDoWF83L14Sf/CtZgDAceuxY6eE+wpWpPYW9SdIuH8Ilco0ow2cU9JsC8x
kLioMuU0KuTVcvoJhBiWORJdRg6kZMyNp0o4tf5qhOvWqy/uzhr5fEu79RojsUF1
BfdBLwWDDAUPu/D08XaEDlUeLYXwt0ZP1JRbcQhzqHmaSVkBqZ9w9tuusl+ah08X
A0CVrTV3MbmGUgyX1yZ8D90jddsalPuZicIiWKKW0fJBAR5Uz+80spXn+vgJovW5
krrh2fFV9Du74tHVJttVVv2N5hR+jhgIKhmQzeyTqrV+p4Ft+hbHJE2XAJLueWYR
7MUS+H2d6rKmmEbVf5/bhaeZw1lUVBRtNV+TfMC9lH9zqi7Ye/zSN1z6Ch6WEgBO
WwYahGFg9fmoOC6UBKgX8/IN2poNObiQYIq8Rc56dRhxzjKVVlQDsOqz5+gQ6hFQ
59vRY/jD2aGffOE2QW1mUcL/ZKJdJGWuKULP2cU3PDfDPZe+7a3G64BzUvU/KPaC
GY81le1SPHl8YgPrXh4dgZZuahnXiXPm2pVUrwAxD+0yTOpKgPNLdV6SIG9C6Q70
zXYR6q2FAc9XDKGeYioB2BTOyDh40GUkaDTv4Za5r8nMyQehHb6ZcOegib4adA3Q
zljHc4bB4I/KWGZPVaNKq2fcDQjjLbcYTsydV0woC2Ib5CWbYnaaANGaq+wzsG34
4jBoRsjwEcKquu/1MeHD0p6jqXbgkkrJameJNvMN2o+Ax3sIUpoIetURUq1HAncK
1hEPW/WIfkt/Uw07Qd+DejQ0BlI633lqo/wZZQB7nJ2JY0ga2z/zCMzVzeTsZa0F
/erSyj5BzU+ABwHB8ZlmwWrjy36DTRREESPrYQQTlG9i90jFxjJtg64e6xQOcZoV
Du1+YEMOjnuqv8iklvf29hQWF/UCYhL/316Flw1Qkm+0hoegEy+lELqqoPQn1jM+
Chglfkddkem+GS3wuHht6s+hDiQU5sfARwk5Bs328it5IO4WSuDQjKLm0XeI8J+O
VmPNr4LhwtSwFt7iiW4TV4+6ONIxVOfJslfGv2KUW5c+BY/hf/x2+QpPtRa048B5
D35g+Q/CW3V1D1Wj31g06ov3pLBCkBfmTX1nZk0YgStlsJToapK5QN+NN7XmBfFy
SWec5pBHMNU4TRxmgwP7abkmaMMv4NXM5JTVmbyhI0HHyw86whi2J+gc0olQ11Yz
fhn50+ifZtKrtHLMnq/Fg43uVNoRQXjWNQMi0ztAKfF5ma82fPLBkhr+dSuuhRAn
tfqBug7HRaqfH2/7sHJdq2b/Ud1JXMlAMZjVV2wLM+th9F16QshQXxCBNhNdVW3W
AmexYNYJWHYwUX76pDE7uyxBVRoOBMtaFyHn/WpzYHnXUqsI5ID3xy8Pha1bMJLd
7i3mr9se4CJ/kjvu87pmoD3LDX5x8O4L0yxQFoI5p3B3XryqqJKTI/ENHkuwzY/K
BOcyvAkubIaXuyt7DpDA4MHHGu6V75ZKmIjTAsJhcTXzBDB2yZvA8rq1iwH2unLM
0pIz0tqcf99mA/DbE7XcgXtCZFurF8fCmxDncj+k2+b8GB6nC4sNHXDzIv2yKblY
rWIK7BEJ+V0KnIaIg5oLPlFDnjuhwXMJeaBK3aMPOYRh31T3+j8eBCXK5PqJ534d
3wC8rIFbBRxap3FVrGt+bcoNyYlj5+ItHQFSrqKri8jCpquCHWtqz8LWnD4PQ9Jg
ceNp627SV6iaNgzR7wMMWG+eHfHnCR0lxf9H0YK3fNRt6RHv9OylK8A9k5VQWn2B
bMbplHJerGS1Ci09UMrRHGlfS/dbzHqyyww+KmSoatm11Mp+CZ67nTRBqcmS77KD
4699ijJlJva4EUX4MtwnVip4GmU/XQEoykWx0bXu0LkpLTc1hAsPEkw77X7G/uSW
VRzkxgwNji44+OMNUFLBICv9osRgm12g83CCpajGzPNhkn6jmweycydn6XHHoCZw
27roH+vEhdwdtp3Bv5ipZc7GskiLGtN6OpHB6ThpOIpRaS6/Z0DOg/UbXZj8kMqa
aBBSFXrtum6HbTPIKHmheJK0NtyeB/+IjCIZD2mGMnGhKVJOGTyJNaY3chtjHjGq
LhmTSqfqfNQ7ookpB/5p1TkGaOA7JMqWK+kr+MlvYEWk6xDVTWIGZE+r4feTFBvp
T2mPde0Flx7IMUoexrSzgxosPrp1stFZvG3vU0c8Pt+covGEoRWIg6ojvOw7Pb1H
o8/2h+jL0FGyN7rGbsXYSF05Px0sBOgS/xaoiE3etdnOMvek0PDJ0oBWHJdOsgcm
IbgE4yindqEOhqjPV0wyMPFGnmo77uY9nfzJ9tUM7TpAos7YCBz0oYz4LRXAGhc6
1XZs+eYy/o1FeXrZt5Zi1MYHCQxI/qQtRrXFSt4znxp3wbANbxjbZFAbu6mSSpAE
RqX6Y/sx50jCVkJv+7EJuogVcWDhV2Rzurmf0ka7SR+AW6d2FnAx/QVxSfgOoGYv
jtsRQ6au4IJfRsExuYpc04D29QLBTk/uPA6xoiDTutc/DNEp7rj4o/CekoaOYSdD
3wSqOnD6rdYJYX4ezS/8Sd1LSqE2xcrNpknwAwxRdX+oylqqyLKxhKnRzHQSdxRT
soA0p/3Uk8runN8k2xizMxzQJkzrZGa7GjCNNk0qiymqnGtjxao5b+oMbh3RUkGv
PZHqaJWVm8DdrT+1RtQXcKdWSLtkiWW5c4KrR57meYf/Cgs+Ms96f0f63jK8roPl
BtK+2FqvJrIUdI0CR2U9chgOOOEpq7L93PcPK4RuAy3BkchIcPeZegqR7jFtVrjH
YLTNVez5SMCXUJ2gcqrzizujL+8WrOgzq05kpcvlzIxP8HYG9TWwpi3AjuC5z/Nj
RV7Rc4YDaEBVeQp7+4WqyVryjNR1M6X38dKzYh7rcWh2rQjwtalBBKVuj2uHmVPx
9ti3mPvOECvghKbznTngeQ2wlD8Ez+vLCaWeBV/bb6+mmpJh/NpcbuNf+oxnV2Qy
6m+iycLXUX9Azvm7C3ooP++D7QIoOKAKeHbg70EJE5k5fUf1WpyzZrarfxwqy4Sq
OqihxNCO+FNq+OqEPYl2++LZTH7omQuJI/jro0pbWOY8SdjPTTe3jqmhZ+UN4AUW
UUvxMZMISi2Bm+S7wZrqL/pMkKLWI2LL/8TyLWj89oQPoRLM8M/kfiztSwJsEwGb
ZhVxHw6pzcaLw8CPVsC6psKll1lMB01hSsMgoEK8CQhJ1T17QDx9vE9t1nVEuefX
gXMta1CppKXjIhPhr5RAecav3euRD8KjMVDyI/n742TscZeb1effkcqF9cNY6u3t
e4jdP347bj4XjDa/T/eLUyujZofhchMf8i3/pOBZleY6YxcbpTNPLtqQ1EubxHsG
xLLWTfLW1gXIXM4w9VlfmMfuJwrmKFIIxEC6cv8TBu42+5qMfwmlo3ykybCWY4pA
7+W7XjVXHxf1ImXrRnMGwVQv1CnRjCIdAxSKujTb/slEAeFoJsPZDYNxO8X/J39V
bGwemsIhcy2mJIfYhKPF5WKoEMlYzyt5wJwdYO4W2xd9iSdE+BN2DtrZpf6YYc80
hlEYulL2cS4xq+AJqlVfw5VWjxayIgMgp/FMQP9cmechpCYjc+ZrW8855GokBeU7
7rgILsKpJHJ3Do/4chcZWGinuSrGYLCmqacrA+HfpPvfsHChkvH25oWTJfOWaXWT
gwI6dgHbCqBozrQEbT77nPipiN6ObZvUpBESHhXMcDsmvRaiORE2VOwjum+EbpRH
t4yR1JxZrsldWM7L4CnlvHpjD2pinvTzg+d+7Uhc4s4FhC40N7dssMblMQuntuOh
yoU38XUFcFx7SaQhGtDBEoWtdjZj5+Jn8kDiql+subuJXOkmfdxF4CXfe9UoEtoB
/jQ/hPls/Rqx/aDIyahBFJpA+rCeA68mjEPex8HrYDCky00nTVRyuPMV6Qhzhi/t
cNbe3UTqlJ38Vh1ZaVPuBQQpZycfIb8KuubwMSgF0kEYHWgNqF4O1ze17XOQxGG4
i7nuzLM5VsqlZtXNg7XKQY5f8/gjLoCzrUrZ05eOfvtKgS2DeYE3olY49GVwJa5k
8tKfq6oJzed4z3eJMB7ZgpVAyEGMPzrxeSCYPT1kMoZFsPSaGCqY8VxZ3Pkh029+
JASg7XuOirRZnjq3KOqG49WVHANo8de8VCbLeqPRwRpmJKxz6q8g9VMIr70uCF7n
pBBHTyd5STc/Kyv0K30HciwIyrdmPIHx7i6k2AfDfmALW5YCtCrbTN0Kk5myNWFh
MqsCHcz4q/WiDevheapl9UMq8FO8kvI2px2fu2CYEFK7rQXjKdn2BkxWA2TFnaZh
xST/f9stI3oXzY2HsMcmO8fynoegbLA/KORGEXcYenlMpYYzjmHsqZJV5w7J7hWa
rS0YoIVgu3OKEua1SiBXECCMBML7Jo5hnbtaCkCNaeztC8jXflrWABi8TxS5wlrN
UNJljfduHCIQnrJTQSnAuCbNXVQ/KwAJK0b1qmYdoxegXqQichiBFz6FEa/93h5l
UsAh/FSAPGWyypulh5T5AkW+1PKl3VXPUVOr6fLMQSRT8qMTP3lBQfT134cPHIAg
Mso6E7tFvB3haFkKJdTOXuJHtLXM6LNI/k7x4W1TCKo0n3uv3beDCI62rnTtNywN
cJVU6CULDS4sbsjAFR3+P0SMgj/BzT4V7ZuAK0TIVSg9pZ8eUM3V2Z8k4Iv36n/6
4uitDrlF2GCitPvplt8pSQbUR9O3rFlWF/4UlBhleUGZgUqiIQAwYv4Svt19HXW4
ZVgn9dhc82G14mhxexbjJU7MhNXOvDIvANoLIY6ikEqd5QrUHF3f9RWnZlX47iQb
WV0BoTRA5zLWS63no6W8ahQmx/VdM5CzRj2gYp4n+TLjLqlK2fPVoCQhiFqKoxPe
pJ43NwQ4j56FQPgCAeIFwsIIt5DBpvOoHG5f//60K7mIw/4i5UCeZ6Oszompz+xX
dHscpaQ+GfpvPwdhKpetyMJmtF//EsCYKUc83UtABAUdG5+uxqQf4p2PxBX1e9Ee
MS18livivt8azIhaJ8zPWDYlkOMbqu7aH+UNuaVPqLthtKeO7XUfHxhf7xZWM8Jc
9GCHkdF/84rU75BqfREQA/7p6GNzdmkUILI5e7ajGVmVNQNtPzTXcNmXfZBdIF+e
leT/jDAtrB9Y1c2fhZXBaWRmW4HGI0SzVow6dEFJU88DoBX9RmECmXId755nJ87j
tySW6pk+wdfTHmn2gvpyYkEubmK+ZHq76NilEoG8d1gcIYXu7tTEhxB3O6btPVGe
3LoUjSslnBshB3d5Mno17UhaD3iThnRrIHluwmUL5UjzPlJPystWSVGM7DzekajL
y2xsMoR8QLEPsZBe2k9wZo9/R8YvWYhGePuTib5iHaemFt82jp7Asimo4ql7Wlb8
0/pqQDtJhcu6Hf30gqnahPBGYXLxJQztJS7RujEg2Atu6qcj/phjo9kJXHlaWloj
iYVUySingswbabRMFZwDLy3Tiw5fn4hvt+wmXFyF1jIkwxak63sVbKjK57W8IoDO
H+AwLEe/4we78a/nMvDPjCyRuYyOws4IZgs/c9g7lDijrzUClMz2YqDuT2/9e70K
GQkG68txKLmOUBWvXZZcUCrd3xKEgPwTAuB9oTZ7UtpK6Kz7EUm/80HQpH9Ri4ij
ipNV9HMGfAgiR+kRgUWV/3wyyJrpOdE2gaAFyhCZOf35P4YTJpkuj23LPSgoXD3v
c9CSn1jQLbbIkPlUnn0V4NY9Am7LEPis1Psl7jyF0eDLjyOwMQHVB1i/9sXdXOyu
XQN39Sd567VD2ykUXRy1c3RpUBEq/MMtiOmzURgO7RNaVb8KueeEutnpHMstQpwR
ZoGPsjnudmo9W1QHy++n/nku9jUE9YRzR96xxSyuxfbd/2ve7lHQx7Ks2U1y1emj
VzfnISJShGOH7BirnssVPac4nRvs1pzS0oS5kr0vgdq1j19IlLXcwVuQtzDm2EQx
LmkOX4MIsS2OrpxsIMTJAlp4FF6vu+MV43ieGwnIGgcC3UYJjNKB0mAvottTaNh3
Cdt4v7a8VGCgog992rZaL6vK2s3KrjiX6Kf3RVQyawuIUHRhQqpEnMlrngwp2n3x
tWHr7X6QBlMR6slFeRj5hjRi2AeF6Phz2Oo72Afv5xb34sn2jCA9Lakrb91Deo8k
DXOwwVCPTaAj9GzK2zY84ic7q00YO/1y+A81cJkntRbKYOGxmgvI2/10vQBu/n21
IOrUtTtDnuVjaQ+KFlTd/tmfx2gkCw2/gLbudJTEfoAHFp+FyZPdF2zdW9ajwKZ0
KDf4noodsFisr4wsHtJAfMWeTrZ6Vyi4l14xp5BNZPuRdnZrsgbvdQTsy18oF9xa
BFci9UJi6EnPe9s+iAZiJb/OwZG0Uy26A6ydFfUHI8PJp3s8Fs1la2ok862WhwVj
yARLYWDOWkoR3H/6zEUgMKsv44Gf9lVGkBlIaoXqWY/1AwauYE2jeMfDqOY1uYLF
lswuowRKwMa9KC5xLbr5RF1yG8q1JCARJvc4KtwkkIWMHijD6etcsiq74IqPiXGr
Q6aFzZZaGkdIpryx7VLgiVoWxR+f3U2A4ul6TkVjkdsy0LvPT/FqScLkO1TSUtNj
mjClD/SsySFtVy7KJFwjE/xtQQEhFR29q/RAQcWtbrp68Ggh/8PsByBpD/nc8uKY
pTiWqKrJkqf5aoZoYZPgia0I0ZVcw15qfbY+hvK4BBaQMHquuh5YOiyQNPXJUD1l
xZCf27ff2WmOES1H+8gWB6r0+poPsVFe6JtBEDqjEzSBon3c9AfSu+D0DU7qWbTA
/Covh+uea4F208SpSNRSYTcNl5o0c0e1ugjzG5OSK0mU3H3IrZckjka5shDV/jsl
LO5u7G4aCoXrFaFWEzTP3YwkUJgP+WGeAMmqsTbCszGxKxBgRm7yN112X6aUdNmi
cnIR6tH3SX0EeT3BKu4tTo+54xYLl3htq3TWK2OaSNJMgnLNSXyFuXNf5szbUIt7
Sau1q8LKZvf4513tI0fIHtX/942FbbqjbuA3PhMVlPexHw9NjxIgpSOLJWiZaDgO
3FZRNBbzePixSH1NJN7HysLSEC1m2JqQFGzDqSSWr5QLqnlcP0+UpMfwgiFQHkgx
nHnrRA0sNL9r/HE32omN3QaxRpikLaurMcDPOHzAWECSEAvRBwtPIngAObGKEFLd
VCmbn2I89x1QiN87silnoCxsCaeEztwmjIyeOuDm3WPTlfcMI9zna2Fh4CXiyYmT
iMU5qTyBNoewq/okJHdGef5RDe/njtA171sAE0ceaEBFwMGTL7XSB1t2AN5JJRPq
gWHeKdfY2MLME/2wyM12EryWzry4m+O4Kjo1jRmyQbOWyFFTBXmug8Nx2XCU4aQY
Q+I5sQ8Vaa2/CkHfCrLUSBIu7U9BXe87ephWlLzG5u5M9o8rFwKea9LnvAE/fKjC
yh+BrYppbrNEVp32glszv6NtcNE5s+5W/dFq9AgB08zsrDcccMo59SrKW8xkFsUF
cEOnSRrZz75HZHCHyYVFxstSadTdc11OemmNw4lrjZrYXUdYgVoJ2OES1yyYqGZ4
h6WsI+zff1BTCoGTvgK2fO+13DFvosAK+OO1Xd3RNeNmNOxdX81ernYQsNgfeJCv
sSssPHRXbg3wP2OlTQMsjwTvoCZKBTBP/fxI+FIlBAOwD2q7aLDjKcLQLBPfj5y0
kXVQNH44R54picID8IBH2Cy6L5nEVQze5Cc8lQ/4OOUFV0Op8j/wIfk8vWrIaC2G
3GWUbiuUor5gjyMFUrAFbgmlem+YKuIKEUAN1GLItxxK1U3TnsYDif9pDtk6wDX5
PX3CdwuKGld9qnBpko8oGFizyx/dM6s5zCJf9ZMQU8tDTbYPGNVkt46YjMhhufCZ
/eKIQoLrdMBge+jfJiesYdzs8FyAqAhcffdP/2DgVLDcYw1piHMJUyFTVuf9ru4N
ZA8fMtTmcjBQSrRZPH5hSxmebIdfMRZ6Xl1eH4GYehWV3RMFJInk7jArUIPdNlS4
0wCbhB5QrKbptkr8iXynTGehEHuGmuF1Z+LAYhT4HcRQaB3Se1LZsgeFL8etoK8f
NEfIa9XIRFIUO1otwVo72dlS+BXSopp/nmpm6/GD+w4Aq4Pw1iJcB7iNPnrDTCv6
u/SDjmHFTEj7XMLPafS8GrOfBnuiWCCW2yfU0b6B0cVVhtVlAdPrsCd0hpCrPQgS
IzPvDqBu4iOJiVyJ5muijQBsHHil4at1S9TdtCelyEEaXFjeGhYNaWlGhC7oYh8q
+sLO5VxR6dOpBptBuPKTJAo3yo8UEBMs3USLhH/5c4kTAS9C3rZ6S2H6hzFl2ifW
3AOAvN6jHUhpuBHl2DOZXPI3rzBHRggjJPxZGqVWLRtI6lVkZQpsuAP+wumJGGlz
HRSVXewP5DCQ6F75XJ5kdZ1XOzETvjMphoxJscy4+qHtUxsIH9vJDvpz7PM9tY59
7r///LjQPkme2PSM2AIfLu0PPZqp8bMq1KmwAOledMZuVGG/+8XGq5LBehB/pFqP
uaW0jZTIzdFnFtJXo68+moDg0Hm3h8Qe4vkAtdY53E71JezTui6ByLDTj/8ZmOeY
RfVpZbHqMEAqXYxX/prh79/tqE6ir5CUYCc2ehoE/MqFD3RD4lTJidFGH4ehtIal
1VyS7mD4c9KwXQS6D75bAZJ1LArKfPRn3GuAMT3LD/jgrySgVAu75d0e5LjbMYrh
mrspYrAhl1Hh3Q1XxRMYYJM5J5AmcF4nR/JLb8Qpdn0sIlEYxvQ8w/g5JkxKLLKq
EryHX9dhKANVPJuvFPEmf0SjCNYusGwyYgn33Myq41bk1D4AYkab750bV4EHTwKW
9KOvjkPThitZ0OrJUjBoyPmhCBvaDBd8gdefM01+816PoDGXCtw10oAMx4iJMW8b
odXIBzproIldOGBrbwtOSASoS+Wr+xWhakG21tKhtMNqCfyM4Tbs9+Q3glY6Hiw3
Q+yNiq61n/vw1I1v3DE43DHKfHChGpKoseBOeyZGNiP8U/9V1O8023I1Tp/iou+k
bGBPa+jK69EbidVHLPL3BJMCwbS6hU+D9hYK7gRCgl23Oox2SZlGoVfZg7M9EVBA
BgwqUn253x1VnG3GdfrKSvuUOje63Bzph4gQdxGj+S/lebkZski1lC6qFAbBuCjQ
bH2pA9Y3yxglVw5z+ZSWyFe6kUmpnXxM7gUzn/5qSvdhgqecoJT6EVl9HjQ4TtYN
jCqh2wWD4f3hI9C8WWabrA4aD8AY/oMXQGIWxJgg1JLz0PxyypoMIgkh125cHRlY
bDdbmsSE3INitqiNrdc9KjpjMLcRknTU0iy79TmS3okL5qwm8BhkOwJFtA11dS8L
iXbfWmYVqmqxOK4G3d1Mae8hbiXWeDNqwABvmzsO9DAwbc7RIxJIKTTPFtnw6OlM
vp/s0nuqpoa5buN26xdk+kRha17YPKD1xF3m1Ce8uK1mVtwZDmTJ9CscqZUabsjW
VXpVugeWl1IarwBIY0iQoT9W0hDFpJMEtY0uRU5eWFo59fUkhMB3pvsM9yPbPlDw
s7TQGL20534xsf1q04Qdsy3NjhYam1xQJoemtWxpOlhYxp5ow7x10XCe1urvaYqU
cM8/y8MHgIqiVwJCO5IVMAsa0C5LBAD4D/3D8Ja8+HFkn23OdPXGFJoRTHJaz8OO
w1byONaYw5iqf7gHIZtV0uNQFS5O/CyRD4CbcJKs4xtSY1L/55g24s9MTqDCPGVZ
1gWJOXWTVWXUKmpBu6NwBCkBBwrfS0gWG358Lcxv06QLwaB4ip4tzsioBIeJcsMk
zM1L8szv1ko87/Pnq/h7JP/kP5/XRwtMt2z+QxmakVJ8kgWhkrC1jOeWYmnsOMp4
YJYcNGbLCeeu41WvF9qpSFg0AReoIf/zMvGzfiptM/8bINQRdcBHX8qANYdGdWur
hcoNHPf0loIeIkutPb9BR69xvEm+2fatLQiVIunjE57A1nk9ljaLZ59bYNhdjMBk
s25fwk/aSFuCoUnDetutsTuONveBk0RjahbOA5NpLzJoJWC6ZGtT/hODvINo/hjW
6C8oln57rL1C34ciRzUy1huUycGVrx7281r6ky2teXdprzknfnDgw66x7npfwQgL
VrEFlfRTtZH1WaimPAD/nN1WvUf1FxmLi1c5mcLqGX6nv5mMiUzyKpbFamcqVKvh
EPtPqtdiN6mp7YLt6DAZkg3fAUXKcYKo+fjTjnM1Kt1cExg8VglI9Rf2Hr5Xq1hE
`pragma protect end_protected
