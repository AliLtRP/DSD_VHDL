// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Mnf+zXfVKLbv0+Iy22maW9FPvOCMQA63+Sq9kJGMM9+hntPukFlfCfqqxJEpCpuSdnh9jC/N56Uk
sX19Z6ovtUeBZIJM6SCijKP/GaDW1IPLatXTI0iFOuMgKAGKlXidR43jpMkTi5VGhsnYJ5rvF7Fh
iWCXXLsTkzphCiyy35L540pQQre1bZCRYc0dwK2j6Q199KogohpaYscfDp3xHtvBGqxamHkI34Ok
mXcvl7Qtuh0DYT102zRXgblX8tteDqtK3XNOjtb/2849n0InrDOcoE+748gFGVDJcilbI/SwoGaM
lKiNHaAUDXOdBxSPsWuUZBXb6IJyJE1zpqgf+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
rNikh8nbeRyF4LwS+3RewtvqauqkukiC2L4fdMV89jfRk3OPLII8nWDZEwYIRO6cjss0imeQRWNd
HRF0J8bibOj0JS09ZnHnwEltHojvmTeCmX7OlJgfLNylFqfZZkbiJnGpmD9NHipRzTnG51PKijpc
8AsMNmA32E8GGl1cnD5eUHtd71Ja+VFzysgauCVmw17WgKLXvO/p8mt89opd96qf6ElBKtggHCzT
+LOlw/PeEvG4ZVeexSIQ74UPLVksSpHg7yVyBT97CT931BGuBiUlGBtiz5GTIq3MBKvVXRCkpoWB
Ze4gcQKIvAQ99FVqvYl+MCYQ6I7eUvQH7cKAWakx8sFw/EUiffvtbHdSpZbibvIoL4n5eFfEnRg9
C4Jw1ssiNx3ZXRkJ1EnNNEzDMP9S+cby5g7+y5EApDeWQUY/Raw57Bbot7JKEuVFqX+jE1E2MA4K
ExV4/c7nm7fwTSpodx9VYnP0KnJbx3pH8RvuzGL/QbvivGWGcPFypPjseXnwjuwwvVlFFp5DozFF
cPwwSI1iJSgMmecg0jFGe5lCJq6Ah03S5QXCcOmjI7fuYipsIV7euCa/xaxBqA6AIVIgxHWCPIX5
48Y0c3TG7R1fv9z71zk2ncxPYHgMB6ccFqZe9fGMYh6xKeaGl9K155IMcWQxO7LsaVIqvOEwhf8Y
+61nHASgtRGZFCV2mo8HC03UpJbzJqVE/VHdA+dp8K+rC7vm4+qjbk69LRKwQWTYUQDzeWHwmCmR
0cchkVgeCAHW+JYN6TY6ULa4VQFAGfZaMkN+wZvoqenGtrefp4rD8lHKHFoG6c/xV2RiXJUoypRd
4W7iSJwAYDjZ3ndsD+NanJ6psdsxgPkcWcdr849ckY2CDpLd4UktKPMhvqgePrEv3ELcNXWvx4vL
VUOnjGjqUJE8F7CRstT5u5765xyXcrfkt1FcrNHcVzLsNC+Ind5RIOjBCPAfxVkz7q+NOdEtDKKW
SXx/ivEr1fppVjYHvv4O6a98ib0AvWZ7TFeH3+UMLHmTW+Z9aedy3PmILxRvaPLgiC05dvgCu4Di
vK7enWYY2mEAUi8mkq9AL1hgdgDDKNasst+l2izyKaxYmESGOZVJM1jX6/BCdjqp08hNHLrlGaaG
9Vsgkahka4uUIZfR7mM08O9QhoN3DjkSleG6E214CQQW17aoYNP/wtYBaZdIBU7xVkxslR7hoVSs
rkylP599thIh77/qDWIZ1gEeux9SrM4TPl9geurTUrQIQcyz2GtN/NBhRvJZDHlYTzq70uJQcH7v
cBlNdrwm8VFY7/46r9OpAiUXOFo1G0SgWiDJYqjuEeiYH0+2T4b5Iu5HvGwctfyvrr0a5kPDBATT
LvgA6gNAOokXvZq0JGRX5Uxw7rJcaRlcfwWcuk2+uhWCSbEj/e5Hs9C0BeWSLrrVBJfFFk8V0fqc
ird72PVBzwEcxRptcAZBDZMozt8X1XbO20gs/kyRVFOAAUa6jMCFogrcLjW3iYFp1xuA3aVr8/NH
MECRqZFqPQyungg42X5rEOpSEL0BIl4vxtN0lT+clBXWzGnoTs07cXzBSrUEY5rYzHGva68Ykwia
fDT9/SVff7fJTqDBYLezl7NjyOuKFj6gJHpsn8G38/ETloNkPZbFsw6isLqpWf0zZ3zswToFJohF
Yj76aGVGn+f1AB6nFUujVuB4+PGozPE3a+wpm/q2qo7HHc9TaarbA10UNyuxTyO2aV5tR+k3oVMH
rQs05tbvGJA44Cf8YT4OxZa7O9Z72r+RVBFPLJXaJrSoH+jnuafBDWDEvgDnTjv+QTiEzIAgKD8D
ecvvWukP+kR+YIek/bhDhZNfbUHo2/xWKDB5q2EsX3OUN3Ql4Sah95k3inLsIMr5SYYhzE6CroYY
gk/kk7tXl/rUOXpV0a6rnDWOro49mkLMfHEzSMNj90zSJMmsx843Fou/gBHqQ30Au878Egdlq8Gw
KUslBoLoCI6pfL5yS4a0UQpqcgpsqETt+ZxJWx5UAqRA6BVYTUpE93B22P7OXvPMsJSInXAigyUF
NPFwZDEuT48IRXD0B2t2t7f1kYwrJVKcD+TZdCtjDykhq9GRjgpu8/OF4xNBmIGrTfqi8DRy3V3B
QJOHgDTFiW0sTgRMWuvEjuZ5s56uexwbvakgcNds+MGYI8yuaEpc4OTULuKGzbmBKtMCgypu2JAT
O/riIxp65tBMzfz7njIlF6EzvT+0EoIwIR2dHirSL03p5KG8PgtbDr45OlAaCoSQrIfwReYPczWE
uSt4pv5Pb6t3FUv7NB0eCXC1Ao+lo3Q5kkrdP8SDnZg4iY/hTrwpqDIzsQz05hZApU+BHhK9cKQp
K+hrCOxFfwNPx8wcAB4V0zzW5clD7U7oYtiLa/fCI2kD6TqdR7iwNg7U7oJCu+lEbWASJDKKeHj0
y8iJ9Vlqo2BKcVI7HUGPMsbpr9TImBbyVxlplCPXbIa8UsFqaaELEDMFrbZ0Oyb14vy3Bn5nXtfU
MGfmURs1IPQm7aHBgjZek8Q6U1BLx55yWj1KkDR6VJuEK4bSZj9IvbKO1VUondRLzTcVXqD2ZNen
ram6QTJIFgB3zOMEx5zHghDg3zFImyNA2maozD7uJlZX7FOP1gaM/LcUjs20Fn6i7jpxvKfIWr13
N6Fj6B8U7Z3GZnryerB1iKbhcADGF/1/IhP9fiqULOlg1YTaYhNC1llhdCv9cVLDthf9hznG4Ayv
bard5nF9zs3EcQV/JtgRMO9kyXiz/TaYsdexVMvfAyy/jLuVxIFDjpAGGSw4S8sWFlKmAK1KXWgj
A3Tn2RbS/3lniYe0M3VDwp8Yv4Qll2Q90UZ9RlLjjDcTA5iLQ7iEJUTu8jNAquP1tZL/It59YMYr
sXODz3/ivU74Um8qPO2P9NkznbOcOFkj5fX1XRPcCeWTP2Tl7rFBQ5e43p/3LtbjcV1r+iQ9Qr44
e4IsGd9LFL5FvsoMMh8t0Lg/zO7piPoahLQ24uRbjOdgLgvp85Y79l5cvSrEBs5E3fEBMtIjDw/5
KvSXIkdIPwYLZRt9NikwcvyuKvtdkvqV8+4csYv9egM/w+NWRmx7lVDgbOgCfdmKBMkVig97xQNE
OMI0il1zzPDYlRmL4cGR0ICCrlb7PqkWOs/5f1ch/HTXFNUxjvwySi7p9m098Bx86S6zJpV8LbhI
hNzScXJvmfomd8dHxLO847nybFOrkHFuAdnbsASWEXxip53Ns1GpGVntXeMbHYfv3tcWwmbXRpwc
qHg7y4OPI1iA4TU9kZn11CnfMFVp6e9DPrFVcJ/qHeFmqvwmHv0r1OaZNd6eJfmX7MUkPXJV3xZR
lb7oKE/aK8YsxTT3WL2RQcOeDKblYiG1TQIOhkUYy/EaNDJWHZGeN1p6aTJATOxbU5yxHBXi+jmy
Yev8ZItMqM4EY1ZYWe9GvvTyF2ehMJ264sB1eLetBtz1qJpAIWJ8uncChw06mnrHjJRU7h6cMiKY
PZFz933sdnbekXrtCMvcupeLfrghHW8vOq3FO/cWDlzDwF5kMzrYwzODUuWKkDtg5gT8U0GzmEi/
DqqRe8rxlwaLWuTsGUw4bxGSG4FXUDzlBJ7nuk1w586S4kBbNNWSUm8QqKvWTBKrB2R4SJWoB+6Z
2T/Lx3b5hdECkIo+BkIwCgeodeQvmzX7mD/AiKu2Hm7bPoa/1HkTvZ8a2iOg2tITMV6htgOekIJV
aTy49mHP1QldKHt2AiIR4V60z8KPvpAQRw73U/FYebTUF/qQzuMUKt/M9/5btFfE7Giblaj6zyPs
EgO5yct1r2YkBuwp805TxqrLzzbFxWgoKnfj31Ju89t4wrCezQzliqoMow2yT8ojRDqKQ8c9jJTi
dujtzFz7GyofWUVKrlngsqWqC3o45FfzdTXrpOmnJTXvqHb2kqk0RtM9o0yC7J5aVO502wmV46tm
+QlWiPZ0eeDno8nRZnp+aOSIBYelY3dr2FfiMnoOv44K7SE7YXXSvLzvDPI1Xo5lS6TOjbpZMUbr
I6TUiwCSMHHrgN7ybNob62NRLR9yJ6+ntyeTGsejq4gIytTGFvWsxvj5yk8hFDfWf/ZzHn/g/RZb
6qwmXCN6sDWld4Ilp5CG3iKoXmw7/d6uyA+sYIVGURaf3a1iU2rkQkkI8zYUJb6RoiUIIcAAGvvc
MiYKVf7LNPWPfE6dc8/UDWUeVXLcTuADBHdVxN+BUeTDh4cEZJJwPAssbB1oiwnjdmH/6S1o7bdj
uyf+NIRd1SZCmrUPyKQTzogrGxhOwKgqkstnxasCArbxLdjPgpKF9T5oPHB2kTZKgriXHtglXQ08
UBudCABqRqS4G3N1gMfCujDUtMg7hYtrCc5ZQHG7GDJYLJeh7wDbGwlz9zcl0VXcupRvpcGIta6V
BuSaT+iZQrsxj61CXUCYp/1Uvz8vcZPuJA7oigZF9LD+eQCu0bheLIW6V5YEiboTURLbw35qVEBB
QMo7zff93DcXEvU9eEg3RLIF5LksiQ/8vZc2IKqAuZX7fhY7vpUHjsOUmEA0LdPV+NhQWKFRFCZc
+PNkv4sq2IoSzu/ivc/WQycGZ3t9WZ2yufQ6OepIM3cCmwMQwvrWEtqy+agr3Kbm3Z0oEdJRuSvp
yJVUMbK1f0iXUMWN0rvBS6WRSQLSf91w86yb0j8Emooq5CyrvaS+prM/3YsKpZd+yTfjUK4iagw3
N3M+r2c5xWtjgJudxDPMCoSC77ZUviUFkOs9xnAIPv2dxzyoooZm6ya3Koy1/4gk0zye9jFNAWhM
R3Lan3OFMeQDKdhK2pr72zI1Y4iDWKgneIIcpz/WN3ukoXKz2LtimmFGSQJOEn/Pa97gjfCURTR3
z8c4FrmzEJffkKkFxvC3gU609HyKdl8APKZpldHRB26k1adAwzFGK9nzxG6cw/oxiztT60V5yO/t
nei5koO7ex2qpJVKTlHDTptBMpvWazz4ihptuDYxeKTzl1wlmYBXACxgYY0+CHpB0x9XtVLV5OFi
Z7GGLcsbG1IOH4OrnrHjVr1Xz/n7ShUZBaPZJR+tmJGScxJxM7WdW9rdW4BlBOCyTkrOGIag9q3F
bXP9wgCSLwGg7Wh5U39nYPXNxc+Rk3bRAEpt6T/9g0Ivi7h27I86hzneYHH75n/GitZLQFYx/dAh
QXSVNDtLnS+8YHWuJneSEQ4R42cAgbPHXCF08kFf0Z7hdSVlJTNAtvecrz/Wzba0B5JmaqOWZEWX
1sWrkZ8sPPfJmkce1CAA51eagyrCKWoHkerRt1Vj6XAInJWeoCK8OPRSfBhyKH242cekesYaerGN
Ihcm9kTGIEAqBzZtDPaWCivKTnX79Bawe3iczfGKKDDrN4B0rdMKWhuB5MMuVEaW0YpQg2IWwTkM
nF5miGlw7nsrHysJko5NErQ/EYIhICiDjX5VtNrzJ/xLKWQRqmFmGqBbW2R9agIVDR3U+CiR3nKq
W7TUclA5++qv1UAYQbBCpWkn97kPomKVqfZ+vm93n50yUl7Ces3n5QvvBmRmL8ObWLmGqCDq0o6c
2tt0ayaTLsPYOywrc7MF1FzRQb7zEzxirfYE4KzM3Jua+h2p8zVS6Fu/jjdcdjD+dvttVNtDCe1h
dTQDzm/t38vF7R/uD++TJ06UJ3SI06nNSllchF7Xd5LfK+CREAv5bbs6l1rBmZ74aR9idu2v8gOO
5WNqfRmf4KaSWCZ7owI88+7h83OMXq+3E+51bluBQHWqviz+TGXsvtVAVTJz7QhYPRO+hf16V/Xt
PZMjj37rmaZm7c4Kfv4dO+gKUCv7G/h2vQ50LWTg5GC0L7KehjxC2UW73JV+PKYPjxOp5W+jGK3v
zq0HoAOBuLFcZJOxg+6JVTNIhp3eYOWLGot7bzBlLhHyMrz53i1WCb8eQy3WYxDZ/siNcoAOoMdo
wtczEOYt0ObBO4Ra5HwYtL3Mv7lftHUChqHEed6MzpEQKBuhVJSq79COr8pQ2QgXvbWUD8/Rst7k
RsKvgQJ5YE7X6aHfhcGclDl/6iAOystk88JO6t27Ld5fOuOlzoYfGVpP05Io28ROIdRYdBJ+gcuD
SYUwimeFZ3xXljHHtjo0a2VA1P6kvxR+WUovQYKH2VLU+Q3dbHttaWMs1M9NOJnZdXkiovR/110E
sp223rds375xnfOVtajgCzKP+zlaM0uJIz6AsKMAx5DSBgJ7XnV0q7UCsXSzy4haXZpf6HUcwlU+
fhed0TCI88UNH8jodKptMLvDFIMoEMX5a0CHjGUYhsd10ZekfUPhHnUPyhsuNaUCkBAw5xwUodHy
JPAqMQ20XX3kt6+TmGqLlWTtZLkQDiJsHPAtTawqlWXvoamU5uB+Vol9ZrZJRmuaM2DdRXkgAe+J
FxpaEQOVeEdEsQW/xjH1JtSizFvmVHqLwDLZuZXSnoXFLs7a0f2+2r6gLtiMYsO2+Z7mkxjIk8xU
Hc/VJnaoWKavg2w+i5qScoXRpZ1Lx1yosovfQghOhjFpKhJ/j2qoBtw5tHsuIlZwFtHvpYwxYk17
0VOXKbuQnvkohhQDoJpAnaCiGTHwQulkQbHYXACpZ1HnT42v4UglvOP9zyzmFi/FB5Ne9Kbig6m+
INCcWe/05RnE5bqt+7kS2KnaAcYmJp8c08l8djFNl11q/u9DGBZkI9xtUwh+Obu7IwK+UgzsZ8ke
8gFH2rONSMOcrlV88KiHGRnLxmv/Y6Wm2FchOyoa4/aAMnsEdBc+7ODRY+oHsds4T/CQ2uQ0PlWa
ZTqSBQtkkIYUpSFly4Sj4BsqQqYs23jV2aOi+CYWWr7X2PeJXlKhfFrh+jFQ0lwtUvPMSzAcPwJc
O3oqk72Qv7nRSQOivdwTiw3MEdyqQkyErdLRZXLMEztyhuQKkCfi+0nISciD4e0yOZMWIy0D1O9+
Qs//8OgVMSr13eyu6OtLyosh+KmxHhF66RwrA4+aG3JQe33cNNzEwmQuBzw0TrJhR2SDqePEucpW
8OvMex8dJgKgVUnd/8fcEUm8hxZ3w1k2QgGD/WInzTpRM36M5EdgL4bxgAelqsFsvyqnK0kH1ehn
grPFqCq9TP2OVQHZVjrLBQ0mgAHhoNgyp8rkgLAAi6K0t1Eh7QQZtAJw+fSThtxL7/2VDwRCwOY1
bDNSvAVpPW2brJy0DCkGr6+RW/ucOod/jNTsU6Gsrhn3Qs/dllJaqmWS2Cd2poC07kMAaeDta9dU
TRAngBPUOHJqDiIZ0dmPX2xV4YAxLrvu0jl8oimfd2s5mss8H6NsuEy4y9Iv5dp84dqZ+BXPwjKv
/yYuP7QfWHfj3HJZmweYmfJmBEwK5DQvxUZctfMvn/SlN8LrjwafrcmTRMziGgS37j+vg1a4sczA
IpD26JqGfMUG/E5l9PyuR8uC+oh9otSpWBBeuNbjUm4izB70VJ8O+DeRcPyOC5gDDqjbkuXsjQls
yA7CEQ7bEbokOu480PblsveoY7QWFgqleNMhS5CG8V7QH4Xo7XaIMa8OKvh+ufToMtx4mrwHmyVI
QFduXQX3V2ntrQWE3mbc5XZwWzRd9vHnljo67iiacUU/R8YAChe2atp1LuO4axmSpoAhxMkx7wct
f4aDht1WuhoWHuMcTxJn/UueYoY+dEikvgqykczob9NZo4My+bJCw+nqvrReiSSs5B6uHvLJC3g9
OjIin6DJEg4yTA3NYY7yj9/ifUnOxLlqtkAE+YODD8IjYtIlCS1ws4zf9NrCoUWwqjjePXcXNNN0
2GlC4q0cmZlOf7qzqPAVyTUjuKuhIb+bx0xvI7+Tpb3E3WgGtd70FD/ncdj6yssZAmiukNlxyy1i
KOTeWcImP49ccMZ+y8/h7Ud86vui8iZ2T7Ub3uaPhhDorzMZrIgT8zUEQFOr3kCKoDmhtYxSkVKo
1mrTHk07RJGveRlLKSUfs5u2TzasVv/v70apZbAZ1COLLvCTjSBttsXSd9Vrw+Xb3Y9NoBaeIIaW
5rxSnUi+nkFJbzfE//8Koa7lAgJAyudzzaDTxQ252wuz5dI5VWXzQY2BUgsK3Yul4EYB7Ym4cfpt
GHGw6vFj5NcO0baXeoWLvHptRNWFCLjl4kC6E8IOaAbyVSAAmz2xFORwxugaUnn9bac64Q3d6npS
hz5KffyjwXwLhU/zKU1JpyE+zvmIOV6WPn0FOrQXf/UQEwtMqrbs+i+Cs53IDqEHVLNnYOvLfBrI
2tOfU6g/f5h5Cfu4SM5dl0jcPmkQ/2ZMSxH9gW0orhRnBGXsgpyzyVIDjm6HiAAg7ZeuWDau4Hwl
jwj6Mgfwesmqibcn+t1uNvQgB0DE7vajFRr9mrY5DpIb7UmRmLqjRrBT5MnboErssmmKcfn7d8A+
7Dwn3Lj56IBgy7eflqKAndc+2lwI7oG/sFRn1RbKhbriW0kdZDOOcAnk8xK7hgEPBKqKxnbdK4r4
Xd8MNCjTThALeFJ4sedmj7OyZJQqWBowld+4YG4CxQ6nWPS0Cdgmwe7NFBnnSxgqnhe7JO+40Jtj
QY+kDyPja3JPqvZAqibxCEb0eD7fWmpO4zIhIOvVw9Nr6xBMHlXuTQpUBosIGy67WCLnSm43Gw0M
88RumgXuV7v62ho+kBmrAuL4ycE3dfFK64sXURwsxn+PHv3r/7yXH6YlS8Z4oxYz0YupaGvt8sUk
dVUYmbnXqN9i1RJR0NyiUp4hk4tWbbsJ8v1y9PL+pgawn6nJwfvD2ZkSu4BopAD6d/ksw9Pu3vtd
Cz/1UK5/Vp+DrpXxqFGZ3xSCq+QYk9ctFcmmc2VRMBjYfq742LGj3gk7IWl5JyKRxxEu5i53gpEP
oTC44qjoNbcOlM9Qi0VyF9YT9til8ECmBkylltSDbsMHLprIzXyVjK9KfERyQdTaEFb4hn2yp9KF
9GeDX2/4dHjjqKtvRNTusdSQ4gzvwrs75UFxenwoYw9JzzlwdwedEfCjkWrN3N+0CpkfVS7whOdC
yHP5PQrFrMP5rljaq4rnEfmjlkKwnpyg4nZ40H01gwsPZbf9zWCRrhgd4MvtTc7GEeY3MXbhkRFl
m9fd4n4FP41LqjT7DLKjy3Oi3dmBOs/i47n123A/JTiE4g8dJMCjtnAY1gFKHroLGvR3CpwHdjlu
2hzl8S7SEDe7WieZQ75Q0p4KODSVMhQzcRwmH9t3DFzrX7GK3QNVgz7AI6I4PXh6Noe6V2z3KyCd
3mG/eK+N18DUt41qjcryuSXmQPAb8LLOWOidccY3VSevXg+NiLopvRf+FKluI9EDJ8NnBIoGn2SB
PBIGDiqUzdlFTYd1MM6Ux9ffdku8vUE7VrJ7IDk5acWxGcY65wbjKEpBxIash8SvBOfzBy3myHqA
OXRjo1qd/a6xX2jvYAsE8x89JMAkDRB+WUHqpV9XII7yOF4H0ItZPCg3I3u078738lXoa7pqqBrH
KSpnIEK9KZ9HbKb/HjBTZGCOX/QNZO03TmNB6W+9t2+ue1nFbx88il8o57IzAas0IOuDd7+AF+LI
cjzVpcPyS/ECEO86+Be1tPYgQl7dlwdxPJHgEVp1CuEcYp3NbJ1SRjyDBwVpV+pGlJ2CIjT5Tk7M
3pOSBPh8mf6aBu6hGNuOqnd6eDd3ddYrtZKOfdTj5ebwYbfaWQJy7huNTrxdtMdwUoWXOIV4P5dO
rNND4e24LHMgPl6awci6K87cVDAKfskoQj0UguWFLyPlWRqIeP3z3uHTOTjpTejZDLY6NG7yYeY+
d+/85ZmRJ0dsdlSWeFe7cVAthTVadpfX4XMKqeTu6ZpSaD+lNDAuZeC7qcylXVMKRdQ/kVI2m818
ZUWgLSiQXSuziWhVUpdM/5iBKA4j9gwxlyqgHdso0XHrwZy5TB+rSTIb69SdJDT2iDjMLRwq3dKT
Ye3CM7yhiKv2HW8htSgG2jarL1J6/Ib5tpKKwiP9tEpfkOCW6RHqQAv72/IM3IWmGgfMiB45FWi5
PLd3phDCSbMKqNTLXXtA/qEOk5VUp4PSBjm9qGaOqZ+NSwnPU0DNNklEv5v0lO5SNvjC0I91ZPaT
1oZxQ9Ww9eLZHIXKDxhN7fjAG2XILOoq4HnLrzOxno62SA0D0th9oYw8OAvfQnBn/1atLDChkt15
ICmMNKnOLZXD3MnDV0bzsAvqfJ8ZBC9noCOL1/GaRhlz48fHRKEc+qisrXpdhUIyzXZRUy0vA9+f
CLjJsIhg4g8N5oQDA1Cv8aSbcWIL4lJaVJgB+HAAb5bDHz4WdlZXxRNuS2nlauA0Q6mi1eqIDlOB
z/50WbbOySiKmHmBX0Z4ce2VNKENKMl48rNYvlzBwMSTy8GxThW92gxYmWn9RRIsEAwIoOO4EnCZ
TE2DgJEOagcZ/S2UGAmuclPf9r2muBUTber+hORvTSE7bjfxD7pt3peUGl3NXnVl1YPeiMexvFxU
vsi8YmQg1duSKhWa9hwxCf7gGCAtnqwzgAfehQmjgz9FK+LW1E8UU+y/ZGyi55cngLIXqFYoE58W
XTkJbs7XQ0xI3+Y6VWMf0vXsgXHVhsX6kY7lQ8gCgS01K4LTN+/JmpwS0OzpcmNXzrne8F+WZxP8
Lci0/gI3jFuZO86rgeb+SvzZNF2Cn1UOYOCd1GrYbo8VieMlkT1wQJH+nTaw2z4cxbrw8f/rX9fD
3G5LwSzaYeJpngpQSaQc20fB35W05Yp6kNZ/EKdaeqHk7qbzkqlbzIEk3jz3yy6AjtWVf6D3b3dd
B7YshFe37t0fVCWhRUgK5Yehf7YjjMdgUiV0SfXVNhSB6CrZZx+U/nf+CueYY5cqpueN7nPHCsuG
fcWXECGLSfgr7qZJCY0xLhLiws5QpvZd/Ju6ELnIkACf8Srjs56vLgfq1+RA9P6N/NcU/fvFIbWV
3XXnCYOC5HQPlcW1pTNEmt77/G25/CdsnHLNlb3yN9hoKp2ax2RWVOW5Tgk1tu+jacWvJgkya2Sv
H/z0q2QyQTKaE51F9lWm0hHk/TegtqHVnGsW14P73FOQbjeT2hPT1lJkjBElZgAZr4FPBT8mr/3r
6OaJY+Gn6aW8d8zE/NkWCU1LkA1nBA1zgcI4En/6XuM2sciQNXnuDPNnzlH4mFDpo/TvboKri6Xb
Ze8PfFSLG4OdxTICAGEMgYpeuyQxruDk+FSQVjSRixBgxtfqY4ZkPJarV44wXy/9akRrhveyuZEt
JAgtcldr7qiM3snhY1R4YISreAetRgXbc/fKobhyYKdreY+m5NpCS64MlqKTuNJtVz/KWw8w2zIz
FxDdMAC68lfHEiQkGVqpMnXAUYZpCdkuwEI+04F1tNqCwtx4oLfTGTLdWlHCJBzdBqz/FCEAWSBr
M4XY0ANVg3M1Yl1rJShvHz/+/IxZb1HoekGmGhdvnC5sl69MKxejSMvqnIMtrQlGkbQUOLnLkmsU
KZTErPcPcrBDmuxBYmIxQ2hfB9CrwA3dxlRRKunEoqq6QQf0d+K3DIgEiL5U66uPXXlo/F6r8iI/
tWm6xGxK2UOsyjCabjqPTTdu1DnZk9UOzJaMC4xHM58WrwRtCm++olBngEMZpUtLH3neStp5QPHz
Gwk2ntZSFR9rUq1v0nNwr0xa6hvZnTfLQgjum6yPIxUzWq+yc1/pUn3GvyqsA0EZHd2n3lnkq8uD
rl4rSkyQd66YAbGT8nxtWXds/6jQboxiQiHh9VoK9YqttJp88atWAGtBRqc8EX35AcHf6D+J6U04
MnNYc2XEnGzy5B4SmmWSk6wiu9aZWYjIhw7FfBRc0T+2o0Ya31/QjqYuQr8BIdZLrWbr41dnR3Km
im9i+utQQIr0N3zR4OoP8zioLBNhR6ndq3aOx6QhMs8MY8B4OFifSRUrtS2NWklMqwU6OFJ98zb4
h0SvON+Kngx0WUO72bZhj2+P4AXk2UW0FecwV5Yd0oFW5e5Mb6iQo7/3NaEMvTY6jl64b45jTwgx
WZwCoc3ywaNLnh3DgWEkQvBe7OxtjhMAnRRuvWzf4IYcRX+d0CrbeH5ZtqGqmnjggt62B05HJnuv
8o7djshbyuPgNIq5Y0DGx5Zy0RF5SIJ/OO8MPRy38cqjwHLdUTHrMaLdMj6X9XkqXWv2pXuOx/CS
b0TyLJfCiY8xIL/1qFGK89FDcGl3BbLFL4n6/C1qIlqWvaT/XKfmenWIhnEvxkXm7lM7vqh7IV0S
pLVnIt8w7L/agKX7YWj4s7u855MaBbj2l9I7Km7+FGkIYoNVAFCEc23AAjdjtgVtIlf9agN28Dh4
k39eltVrmOBqUaJt8WOhqFZox18bRR3OV2z8qT/oqiWwVYAFgfK5lEY6ZVFPsEjckDCga/wajBE4
vMnEyYK2dXoKtGGH+ThLViFGEvGOMhFJInxvkP4Tp+NBboMqnw7vcpRYq5XFCgwRh1/Bsjs7yDdx
ihpleUSUA1jRKQDyMXHVLVC61+MEeD+Du36UIygEVwMN3EvJ8pjpxHyxIbgDzwcTVFCW1flKcZkf
+rL4MhIV3/ntaDKJuZGfES3A6CqM/i9sKac7umThdMO28lW4CvcQyeavf861nNZzKCc7CEoGzUNS
TiMpVuKhDyfVlYz+ne5YCrV5bocKuyjB8ZVflKgf0Lf7vojhZ8e6EjgqbR4jtAxrAMsP2pRTgoJB
hIjIPFIHmfpEbxkr7EDUNdE1pZXthQNDtlRhnvtckfTAmPBcJ2fX8EQhDXCTP9Pcw6mUxNUKnpjO
Mp4wqC3fs4LcGo/B1znrNwSCyGkBgXFZxaw7lI/9T+W/gUNRrWyQypJt62LyUETEAiZEis6t44GZ
rtYzj+thNF4YvPWfRTQkXHnH3NKWSHjBgVybzhWZfPkvPmb9qoph5HcJ5/E1QepxOUsEiYpDcERs
SbN8hi3L6d69dZJOhBYgwkMQgOKVq6w0NQNMt1zb9qtgIn3+Zj0+faPdgKGobmYZDbWu5RPbFm/k
9hRHQmrc56LO3dYGanKLYuy5vcjIlaBsMR6js7w6CVowuLA4rNJwKTlkRGxJivMTihZsZjorDqRH
Sg/2AH3ynignWsC1XWW8byTJPjXur4ziKx7LLNGe7D/oPuzf9Dc+giY6SsCqOumu2JR1oxdo3Psh
gtp5lGmbBezLx15vMPb6mkOWKaeA6FJTRAg3sjwAqXxXY0eFojwpm33ZT323NKEM+1ld/V9a8dtG
W2ClcSPMN7ycGofKmMeor/g7Vxy5A5GK64/Di43insz7a2E4kuRo6Pb+Pt6T5VMGLKha6te5huzn
Q9ZELdXoQ5MV9fhfGUI6HvyGQdiA1Zanu5cSrnjneiAR90S/07dG05LeqgGJzJAR0I1dX77GqM6K
zjinRPGSfK9ScbvAyJsC6hSUwjW+ttA+FdU9Tk3eQBQxsUrwPzeIKUsDvZ3tZm6O78FYO/6dfuaS
Gjj0iWlYR+Obzrz2seLthJ6FxhH6kubMPGlrD1qOwfXHXtqxlZCkyEmWtd0+D2UE+GcgZv8MWEGj
ubcq0QPMwvyHHY6iITf9aGiDHEbr+WYymUeoDhNhVXGURZFaHTLNJ8oQUCJ4mBgFNtlqWcSwSDtQ
WY+n4o2pMTnYFwM1bR5aSpZe79JfvA82uVNWm+vm3OQiqYW1/hLX0lmV5YFI4KEdFZkmBzlMahHR
ZvlX4dhhLJ9sqSiNSKdNz4D0xim6XuxU1P93m/xyHQfW1Rh8gEgx0koG7Fo87NAQ9qzucSSdpDOj
AceE95tMc4QONQohSIN31ic7dUrGbdzVmtNH46O/Qv5/RwggSzanlZmV7J/+4ev123HBGSiL4Lts
Z8meq2u4Y/axvjZArdhb5XSJRV8DbVZI90BiSrzgV2eDq7wmyT5R6BQ+3V4Tr7qZlcHZYV1+uEeD
SPImfnYFsfroCh14lnK6AyNFCtQ5/kXxS42YI90PonCKEhlHVO5RcGUUQ9UY0i8BWTD6nN6WT5eu
ylS44Zy9SUacMi5CueFx2aDSSHB4+lg80Jn+XeDjxZ8Wt3vEVHd6Zu6O8joJJ1yzQaNiUHdq5fU+
n4h+MOXJthmzEArtQsuB+D3OVrSf96SmMPQrX3OmnGGeM1WnUanLfDttNXrrW4RPY1m8CdDBm0e3
DldsEbFj2IY/DaH+/MzvdWUP0bFHPFr5uYqbjcjBu1VaUFDOHeOFulKXJlfPrbFRMWPF7yl9Nq32
QVmWpWIyY4It9kEiaE/Xb5+mztAWuQfmEoJfsfuiIkOHiZjxoaCWS2ANOiH5i0VrMf3ufJER9fuD
x1X3Rz+IooBazoQayszCXq+LZTYXKrJqtab98A5B8scr0DbEWkynYs8fym1/TNIfeVuhu64Ecq8K
O2JdFWKjIZxx49sUYVYi/Vsgftv3wHWUviLYmmOuP+xNjiIOTDdqmZyEHGw9gzwBEfGhN1bLwQRG
m6ozvfAgZanA8te9RfCNuuZU9bp6Gobjb29oAiXoCoBpyYCHsPJA3VuzICEpSUlS8KbWNedwN4s6
sCa5z9sBqGTm3juJR63JrJqzi90ure+YjVjWn0eiKc1a+9LEuKXIJWMnMXY62nsoCBnQAPe4fAAE
wmUTYGrqr8JChnRgFpGFs/oaZL9vQAki6sT82HV36zGBSjP65Hrq+R4129vDzHlujdRPNoFzSXNt
fQ1SrDwlKEJB2Vl0gQ/pZtvjUaY6tYhXOsdmc84xonBMyMb7TJany+Nr5xP/P8crwq06WUDtXVkq
Dpd4UV00iop6+mLPpMRBBD4fzYxdH99FKiuMKM2Une4kI6qYiBRCmqG1MM2p0a/FCxIhoqss2TSD
8QD1dMZIuZzUXHcVC+rJ1gJyqVkLLvI49OomP8JAibrLRb7RNrUj4HE6eSmydCXCsSX3Uzu98QTR
oPAiRWRq8JnlL91ZLnj0orYz9U4njsHaWrO98RiDYfWJu4CDNyaH79EYX29X7KPGChLX/hW0mynM
gGRHkKgnTR3YRZa5gnAD+rAdx83W4gtmGoyjuiSH27kYbwwoiXLIcKZsGXQiMkYdn0mhmTgPGM+i
EwkffFjo/xN853XnBkL+k4kc/pX1c9IbsVKwo5lpF4FmxQL6Co9rn1u1+/orucMS9ni09C8aJV6y
IOmuzWN+mxNXHohig91uSDv7/qU/RyQhzFFsTc4Ol17zjWxfwtIpMkCKIf+KUQkkqmF1ESmUghQY
m/Oi5V6dkkY29u5R57sKWaXFq4Pztp3Lao4IXRLJUBM7ZeldcKlnzawZIMIYgPqPsxuyGOhp0CJb
iyAetXUTRJEEUTvPzY7OR3ItE2lQ67pg50zeYNcKAsqCzFmBEBEl9LXBywAjmTisV2jKT+pqqW3C
8w5Av5DAOvlv6Glum9egH82f0VYhDwKl1RSSL6rWYdkXCKby7NkurB3tAR/1B4TlV8Tpxa96G4bS
0abl0mVtm+45p8LBAg8wfhGarvIuM0oi8U060xLdaQmHDIRHwvpHRIPcwPn739rJlUJAWNjJ+YDz
99GgR1O1zHNSL2BDEffPp7PK7XF+nt9Zhpn8Ba+5u4TVfEn60ItEWaSBwFtoYII10UFvqBi4qZf7
csXsISXh7qWh3cxKsEl2kaf/VKSqrkkdV8p6zsS+YJXe0vVBH1rRkVOfBJrO8ZHdjC7ruGDZxx5/
4mqRQ3gWvtO0CQLXghOnkNXzgHSThGjkPTWJCrIhhRNeRQMLYzIByU5ir3lDzUC2Fznd9Lvul7UL
B/0u29PAxemVqBPIOtE8HnhW6GqRL01yg6NHeHrf5bsYJbb6ErkRxsWsPpFDQadGrVkDfSjmaEsM
FI9Io6jx3XS3vgR/XBKAP4wirm/6CnkLQE77UWilCx791Lf2hx8sctxjSdePShgTaUFGoZH0tMl/
Bd+4quRUuEWkmJaDI43aHiWYenyT0abDoK3tw5ASB8fKIV6c90RJPHEy/5Ad5ekZaC2iMU87nCVo
gDv1ewiRN/E7dyxcwPUiVo4t/pVuPQcQP7wIq49KFshU01UFaEMxEA5rrqxr7DOHS+t3j67G0pKG
iVurWPtPIvOks+xVHTevFu9lwPuv/G33nZ/OvdZBicvVKWCu6EeT+5OUxG5EtMPibvfmkkpa+2xC
39UbZy4mPF1qB6qXQeG5pcpTGKKI3P7k/TDa+mB7J++FUcwH87YEx/RLFuLW+nXQWsy2YGTkVWkq
BCHgQ7cS6oZqnnpRFGp6R96gmaZDZUm16FMu1wTnJiZViJxXEztS3P30gG+DZQMELJqaLMdbkoVz
slcADxi0KiX0fLxqqyGVBeR+CzDdQhFoLxam1nhPFZUIJ9PvZIhWnzWQb2DkHoHsK6FC0h/wCmv5
OeKVufwjvOe6ETf4mh/ifNQ6vBuznGLoakyKVXr5sP92pjjknTPudPZJqoeCkVBjnAf5rkip0STJ
61fUa/TBLqXdSGNA7zNLDo1zqEhBHfW5Vyow8DxIW3P0U+ghg1a5+YFMtU10Lyq3AzyEZQmGLeG/
MwQ2yO8b6HlTAcki9bJYJKz1Xd57gsVaN2eDCzSRaCJZraxMWUcDd2DSBMYTJZ8IIB+iE7whQM/i
y1lwAFN+Ea3YWsrK1wSzXc1JLSymqXeRpjjaTHz1szNPWx/9vNDG4aX44M+jRmfL3T+vVsMdpy6p
C9/VQGf7Os3XFeWg7YygN4Ac20sIUl3r5aXFCGedsMYfLVh/XIUyqYhQG0xI6G87pYMPahd3oe7e
SPaZi7lch2g54pL7ftVNTpHBoCimoY3/T+0cAjHlAXqodMMwMhWJyn70vHH3dJy7NP40RWM+7HlJ
8GSK6vNWDclf0PEB+Gfhr9VOVXwj8AUGErRIQwrwICw5O1UI5UfwUZGgj04oOkcoLZuSdlaXnshC
Kdi1B0+mfUppWzp/5ZR+f5h43+8s4LiMtme7IXO4XkAb753CUPrdYD+3OWE2yBbeJdDz4wTemZpS
Qr5mDmjpCpcjl3UQdGynp4N83XIUkzOPyqXBYkGHLTdUHfv0zRxDJJZYcBkJFc8jm8dp5H/R3SlP
Roa4luQdqyl43wMP2YX/AuaJww5BOTK2sIUBZRU6qHzAeja8aUxy2xnzymr0ecXLho0U/MHchlhQ
of+VXiZvJPiVzl+rzUyoWliCUa/iN300oGHUGDkJlQ5Si4nS0QcMUTZRcjr96yo+mgIdQCoipeXk
wxlA3VvwOZE44h86nR8OwBMMYUbRKt6ovKE5jnXBLBpEHQjrw5X5QuTXhHUAx0Q9YacHpcS/1E2u
FkIJlZ4fJpBhHQW4ce9PY0S+e2ELP4GtcG8sSaGh87lr0FJF9FIt2D+KlodpCGpym/9v+C/J22da
6Xj57p1ZuOHPTRH9nc6LjCTLiiiKZ6VpFjQpH5+e7PuTWGU1F+YmdyKrt3bnCRsc9kF0LtL1np0t
UXd69orqe/+TluEaVEBocZbtKv1PfQ5CBb0z5DRF/qmNLT6cOqbhupn7PycqzLPL2kjK6CbKM3HA
rxT4U+JvG0pYd+U1ggLvZzIlIOkVRKlnCx+MKwGdLO+pd5W4yeRit4OdnpnMQnmTkgoloncBH8hP
ky0IcH3KH39qp2CfnyNSLPMk4WhT6nlawaNk1j8aovTrzRpHG8+YyK1tTkB9TyK3N73IM//21yqu
iUhQuM+hTNsqLZj6/Opl2Q1Uy/qIoS/sleAlOshUG2KM3VKNHf4KPQQL8IK3qGa4pNOpdx/iBUMJ
ErCXQLjsrQXuGdt4ba+DTufha5tSnU8wCgGE4O/04qc089Dsse2AK1JjjV/vNLDV2RV+KJ594V9E
SyDwBn/RSzZMg7zr9PMPoSgNIhVFj6rxH8HGO08hbLmhx2vsXyqlnYct0TC61hUIqoVXO36TOmD4
zCzDFHlbimXkO8sJ1Fai1PjhNCFgJdsCYnonKLIWOXyesNA/f12Yy6rpiIuB8ooroE6zx4pA3xaP
MecsG5UYNPDu9mTr2mhbV9DraIN8inq5GNPE+dYAnjHx4qZbMtDTQrmyE7nHUdeBuLuZTa8hxpug
TOy+aVNn0VjokDqNHbfDra0l5bP8G21k/troTGkq2QWuNxduMmxNV/k8xyp4CGhN9r/YRjlNMGH2
jXn6Ll3hkWkq8BezRYvcSv2SfAhJGxburgkFn5/nAdwCZmv5nJcuwqoGsZTp+8ZthhxAOY1qGqwa
Mwl0ep/MyZF/MHsDkI97HLZ5yM8ASABkWvtr1kFlhmPAFEwFCrnxmwnBym18Mm3qfcEeIadWnkFt
0b+LcO3U6/PZ42G4POtOXwFAN6qCYw1v3QJBsffeaqUbxSBBNGOiG2xN1pC9BvT04zU6tUeotoYg
aNw1d7p6FGnErBLWbW7cvZxo91duRxr7umi4F6DZNMIGo7/16rkC6P2dbhNZj+eoEA/3hPb22Z+6
wc2oRuN4C8FqHkmoQVHZT8hJQ3qZ/UISEmOG51dil3YUMaXgnKaMWY3Gbrh/I5ZF4PRpZ6sXg9bS
buAPzB3s0WN/V4B5YUw6xhFGu59jIO8VJYcKWbQLFTDn5B54KY5QOjPs2HNyMEIGcNabt2g+jUpq
cGtpc+9CmBpRcz+V9UTRvqz/eof8gYwh+yliuNX98Gs/Zd6jkdkPJIomtZ1+bsEcFykbV8MaNGvs
mTE5g1SjWXfhrtVb8lyScAu39FV5Y22840FCZge21znJ1j6ts0pJJ+Sf3l36JdeC34QglY7MWNhm
E9XQSkJmSXT43SIo1G98Y1Vw8LPGzFi4JIvooFWA0DDhSZYNXxwVQqkJYHNJVHtHxvX5toMShRR3
WxGvbLmVhctIiUPlBjUJP0HlzCRb1E7D7yecm0DB3uH8u2W3hF5XhXW9yggjESGR5kOewJzB42G1
uBp1yvr4zAscRSV5fd3ZtEIEZzYGQRw9SPUhG8/aoitHaEdwOFPDWnAUa4och1EBVD8M4zHbn2R7
c4QvJ+MOes7tMMPKTtQj1HYtAEAubrxUnrl7FAreXOllXqr2ZO6LVQkIYp77kiBHP9zIwfw3siSU
h0oeq3atmJDx90LLGTseO7Q8D4gR5iGJQn3IsORx5jTrNTeC+/SIS6lL/vOqatPb3wxfi/gQXbN7
VIoL3LD3zXcoPOwYqTT/fb7eFpG68I4i1zQGQRs47TdR5wtSSVKHLIxT6qXOyER07l2dR6dmfxL+
33qHOHe6duTTRE5OUhRRQNJiqhkcvCGxWIWvAWBygPM8iT32XD+PTb2OwyH3Yn7EgKSfgO8MI1vt
JHzC/jaCkb9QEF5DShE4VaplEBG60WMvdwCbjC13oxHXBmtSe75UeATkNlT9qh7AM46nfmH7x67S
WlGyvbEwXcg3HslB41M/KSMqQD6Ot7bAElwKPIgBnqD2YYGJ80s0jAAb3Mya2yF88zpAJxcDKT2/
LFZMc/aCJBlwhEO+vKf9CaXnf1sHjoJtZrAyV1Y4Vr3Fh8tE04KoboabVDY5c2IeLhFjP5GMNceu
SioLDsIoWt5zaXoSt4r7ncidBRTHJHcJaZkcwOR33vevZZee9KLUiwtPEJBCZILl6cFoFuSPejj7
ttRQaEW8+v5/q1B/HG2eyseeYyYbvej2T0dAq4M6ujoWg8SQ9sxiStCQr0GI5KtLcCr8BTsIL4u0
NCdhDxzPPqne9cuUIm3Cv++rYwHRFOkaAVeMnvGtNLQUKeFBF36fO8SI/qkySGe+Nen2Po3eHPEE
8184szNva1e2PJgdsMi4n1BEvI6dfo32d/DSTYsgvNAVQqlyQqAt+rDJXc1l3no8PvNE0z/ac4Bb
CzccrAaJKQJ6pu4GBvFYpmoZR5TTIABot+jRCvwDfEoUyapFRIR5vObgJBfjV8Ysi1i1/0BypQ2c
/sgKOLZcjlhNxf8AMG9diiLfOersfm+/QQNH8z9+2lzIJuo6s0ULe9EV78Ho73QlTQgX4SN7ihTV
/keczKwX6ooLhRqVFZ44TR3x+84ESy0A/KYmEiUxv5IDfT7fVYq9hOlC3ZUxNX1LBY3xqk8qBTwu
7xaYZ5sQfWKT6LXgY1PlAguHJpYRvrX+SdIpvE4pJtPw9Gpw6y4ZKMhwWBF1TPf8IL77KVpeeEEz
8l4ukm+jNk9fH8llhlhQsVj5CfqjpZWPEeQPQ19AwHUt6aXj0zrJeUaQXDDqcvlcDFd46eJZW5vC
znC99E2hDUcpowzy+DY4i88IfUj4CGvzZnrjl9VuFC56VTisBIZy4UGCR/7qH26P6TY12DYDzeRC
EkGe0TkCE4MwbFzshMAddkNtqI/HDfI91z02BA9C8rkFvMFadt3Z6jrvEjPVOlL10x0cRySkGrzB
x4SI+WSim5kaIM5pjqoNM/IHKSOZjNKuwQ3Ir0x2+UakOV5VVNtRBTYpJX2htEfJBhYveS5JOtQ/
p1FMk4q4rRJWPgBN9oYpjvxIYE4k76CGDJFy0mjhQbecJsdwj5WIeTaV9lUYAtc4xRvAKO6dkKlq
9tiVvPkv7ILudcXU0NarjvjeNOBsSLCzGVIxVMF0QX+G8MuhQ8o49vG41PpXzvbDavRF6ALEdMO+
WI60g2giGj7kuUHph2jFX2+X+EY+BldVX6qt+id/0Cw/ZjIRQ1RSe23xgvcsXKNqBxj3or+tLR60
DMuAW5tmNKX8zcBHjhgtn5fgRkPUfAx+j9/xaQxAUuyzr7C1tWuGmCTLJJs1r0QpQcOMCiMur3ud
rVjHhKAMXHmpgg5pKi6HoZ6QZWowc2rJ2Aswcvsyxqowg0sDl8Z+ljT63jHn2vqES4O21VPmAr6k
m+dfy03PJAqi3jpoWulUL1bw2PxQvuW8pOx9V/j8i6zxjZecKqCZsfy9wV5z+h6e37zi3yjhLiZa
WCgEKCnVKqGV+5kBcLqa767iK5POKBQHRTSjUdfbW/2KptFKgrA1f9YjyMcsruyWXjIVnSOohR4j
CmYlRJQPX74/XHf4wKgZ9CXczDDHnXAQCEnzGBh/N7FLvzhtafEKZNxHlXdBX7xq8Cvxf1OjH9Ig
XImt7vFSEfggEXR3mnonpo/u/RvXZ3laC84ett5s7hM1vt+IlT7Hp9UViP1PzcBTfH7XINazhZiM
p31G5f8g2eld6AiVD0JGCj1VM5NZeDVnjzRiiVnehD5QGslPjr34UCS2nkLUNXdtrPTCokTNOIJ4
PZ6sfv94l2sv1IH3xex6+DN7rsmnT/Yhn7RU4xZTagxcdc02+9tLRlkbtX2XxOnuL54X+ujd1nuW
WS6EQO+MOb9RgMOEvg+ZxTlMeVvmlmBafYvo4l3qLllDxlPMX60dkz/m6oISrXfubgBBQDn7WN8s
pk9emivKNJSWESH433/pRoDtDP+nTXrUx2EWxsigBZahWQDdi1ouraFPCB0aHCd9LRyvgxOpLdk1
ZdmoQV0AicBH1/5uHlF39OWyrcOuXgr3DyLW5JmAxCroP+3xdNfP16l9eS0pn/COHsRa/7fkDMQJ
GZbcOPrhN2dpbPn872nBR7TPncwa/cIv0XyKLrJjKGv9sCzRLBMzIRT1FL08UsHpq8XM+WsA0RsQ
nmx0ay6e0HDwa0mDnzHNw1h46Ez2Fk+calJimLKnQQ/K+UogpK3q9Vw6RqXTqjDeQuHWZUOxM8Kd
7rMrtJjeDpoupd9KgKOWr0Vr6uOtdvAlDX97gzA48dbL+FpX1+K5gOYvaW1dtqgIWKmu2m1iVut0
/vWi0dOz+UDHiZ2j/OHx1N5BGf/q204f4kmznP2t43bMOBDrBOvF2cerry4aqfEiKCZfTcuCL+db
BhBG3txIPuRkRXn6F/etjhIF4zCA+f/gaScSFzbG3Z1H3W9kkjIEhf83V1m8x10tXfN4FBhDw5Yi
VyTsllYwUreVs7BcGPwHArNEjriLd761aYhyFgiD7Av5anctIQEsSPxJKSuFGpCTi8O27px5bTSK
6MbBlULpHiQYrXi+xstarKQbYNRaujg1PuiLpP79vTr0fjz5VhETQnhM4xlPRHRx/MzpBc0s41dm
zvvFY7lgjhTE3HBk31jtUaoXFvzcZ/tHbESgdH5HEKEGEKMZJJ1tzNgJcPV9QTT9yRQOoO9DJgrg
qtPtVcDs+wBYFGQQwNpoQBOjxvByG+xCY4u1XehNZa5cN4/3GhP+BDw0IuCYtOatpbdBhVCuuxgR
nPpPNqlOGm4nTUaATf9OJbyq/HxdNg3sLEPyTmnA4aE9v98b1BvmuzT4AanxQe11YkfTjmJDrplO
QR8/08l1N2SY4jXmUFrOscXC3bp571xE03mk1bMFvr1ZiClM/mCuHO3JroOw6jEW/jHPiY75relh
b7Z/quWkGSfGzeUtJLCKphEbSw5O9KAOoTI3ew4L3beLCONuc6GeKj4ZCY0/06/Ez9+4r6uIVNjX
r2OewbiRRO5RCAzLbpfyO0QA51VenWpY8fn5iTSc1kUXAoB+ewrA1XDJqj++7l5lVt7UU9oe5nV8
itkf0qTHs9SSF3Evtx7dEpa4Pkh9PsNK0v64OkzIlG21kMPOEHNY+7YSHyvyTdA8PqB36/9ujZAT
8q9O/99Igqrlj3x2X14mpu9YB6Ewv8aMlds7VAKDyVMShECWXNbFB/dRLJKie1k7c4pLMN59OCfg
KBYph9wb49KOcUWzC0Xr2vfvfKzdj9GAtRgYtXUexC/uOrNnlk/7VHFXuSVVI/cH/mFqkNJ8IcSa
VkO06UjxxOZwEW+jLL7bxx+BGGpPgV1I0F5VJyLbyUyXCcMdKznSfwY4HXSY7duMyraFlZoM3MbO
4Y5teR585gSChQiwkqcJwmW+z0Xv9MDZ0cmCw/oABL4WWC0tCcgqEuhdOUdkA7WgcteffxV3GlEZ
50R1kkREnckzf4IytOc7C0nnBfACnPS8Ddx24z55hIA4m4md6bnSj3yT1qosTl7DmhBlkkT7sybt
OzpV83hqdXmtaK1BwexeeghqBxMs90X1ENvUcfSd7+yJvJp56LWXTHNiqH/NIx8/NeH8tgKkFk3V
nanvPH84ofzJHIGvcRsWaFuvu2dhzIjJ3PvGqairNrNLpBs4tGuFnSsdmWQ8McTLhiM2Q4ZuQ/kT
DxGTb7idYS2Pj2kVsBaZDiISJBHhK+pb8IAIf70R3ncoddKgPlArDkIp9oCPMJWNGBe7uyN28uS6
qlB3TY7eAgnnit1aCcUoKEnI/6TDbw7Kv2Q4Z4pGfguuMMVFRB1Qo7XX9isVYaEvRAfF5p6f0ImT
0M7/SLvC14NmD/kFRQr9IoMx1APHEMYk2f2BvHXj2xywMYwcSrflBRLg4dGBZv/o21nRA9NQFYH2
g7L2ECIQS3jNBGnkTj1cfrECaXBeyQMWMXC8m2WkcAuNT1B1Ij7YlE6Gs7+BwCbJ6iau+VDYKFo/
pNesjo1Ki4be/T3zSDc3a371OuJJnfBbBYe+vHeK3vfR7MhWmTC4WF3x+R8SuD4h/ptaG/3QSuHH
F7ODnPMIlaijNWwiI8FmQH40nO0PqLn5/ntXxGHugzlBKHjdyuZ1229F9jZRz4NG0g2YmfSC/8os
AEN6lFWxwByxyYsJorxiY//dXYbeQUL/573y5GAAyyjDMLc5hr6LwuP9NVRAXHStrAia/gn3q4aN
735dtHn7gVkDM083g1C9D1gtc72zijk4Q2Zr1SAuRF1wB8e37+giWQDtSQdHKiTZzpr+8HX0m+gN
vLB6ui5ipJf93woej1S4rY9F9etux1sUWqI0WJ8TjUuuPxAofxV/lCNocYTXCOU0jUeCrFDdemoa
4FWDCKwG4GHG+ypGhPMSQbNquEkF1ycLVBzzD/2+FDVAq+lBX6dMhAGZkTPsTZkXeXLhwT3hZU6O
P9oklfdNcbBompcfxepXyMrXr42IhVtNfcEgoezSPuwNd9lhphOswCFz8/TCxQYEVE3rSwXZO4I1
C3+0syk7x4UEoLEIiFP7BHfidyLs5t77mvVNHS/9XDBqAlwzYY4cN+7H1T3OVbuytxAOGkdPAu1M
Ew4u6ZQYF8ygPcCIK1/NWG9bOHvbXfKobMk9w02NrCYd3bK+tovLKXEzxkOYTuQ0DmvkkKxN+vwq
TROhOngzTiMqKCEosLmbTI2KUAiTBHHj8xtL7vVz0klWdaDFmBuE64K61+EUH+XfDTu4/8GyX9Ao
HTRMJRQx+BrO6wt8bkolgDCnovSonmMPJp5YVjbnnbvEGaNNK8B/5Vo2YgB1frOQFnsq8vBj7B+E
eK2QgDa86XIYQTMI/nouWrTqD1lWLINRvkjbRb6/feZB3aYG9Q5fRIxHZer5rRGxz+61feALkr7I
csnk+lQEKGbDwy/HTj3d9NyRWGZBaljE5gqKirUnN0lpLl0tNUuR2M7tOQNXyn9TyZWtNaI+9dno
KiRYgZ15O7+ca/YKerP2/J4L7Wqa+PF7hGYOIFAElx8Wicybv2/d9lwh1+YcXGN3xg0zQJql8JFu
FtMO0ExodG2ghiPceqqrks+PDlS4ejuPTNnWGyiD3JAz8Qy5aMczJjDmBFrr8kuslmZPu2O0LE16
Gu1+ELo3ka2RSJUFqIVoF/OPrraqr7D7b3oXgc+k50fZxvVpBSeAYF4hm+05IuCv53Ff+EKPFlYa
AzXtyWRPWwk3vqbU3h/7zl3OyJVvHIEy6mLFtHyYZuNTHjzf5zu/rxu/nL4Z0197Rt+LNRbaIgCM
QvYPosVBQhJnnZLRHRggA7mT2iYyT0Ni4F8c7vP08X1b2q6XltZ+eu8O3Oo5jdGl0BVvFwQHysF9
dvGS5gVFz2AySADT68oCmdORuR7sJP1l3Yx9J7rcJH1S99l+yzTCGVlGjTjxcSPhCg3XCdH9B8RC
RNM8qAUVCc2gxkwMOXiHxMNf9d+DNfa7ADiCkqiqXuy1GhMqyzdsiuFu52OyqGdujLsxzEn+JCGO
gVdlAsVp5M8+mFBZQBXcm9rfJsDl/FUiEufeoVhW9+cEmzlin4kRc62fRImjUvRQ7q41TKiKAgeO
mP3aGePtjMTFnTK2quDX3hKQawXp8o/XI1OqgASlbJmAx22v9qiTyeduyjvbP+TCXhwJu4PVDEeN
amnscLJBUaYzeSgY3iwrTIBPskrnUxN0glDusu/QFd1hsDgAMSVfIAgT51T/63Ecc6okcWgrKLjy
4DgYvztM0S2Gh2FAFXLA/Yy3dvu6I9FbwJXrB5YH0hviWPjcRnotWDvSkyV/Sdrf8vhg2ZmkzRP+
My6a4UhNdHwXU1H5XdfR8nRkSKOKfWSAuv7XlOnviYm+F7AeCATmnCeYlP8OW8yrfKDxrhDaSAAi
CMNr35QlO7ospUT//vW4g7vNWCDADOy6wbBOn4nIKHDLwRBHaJsCzVwhi6XTVPD1FsVfkUN77SIF
682Kawf9OVhjlNUV3ONUNW52Q9EUBxIiN6vCGImewarsWcFLYeg+xKnCZ3aq2ij6GClxokslk+3Z
aCUzEy4uiLNqpcCYnk1pomrofTrU5h4gEZpo+Ey7hRt/uBgs2KueKIPivhQoF6K0anjzQsmsoc58
70xSKa2p3Ufkwjx1u8waGaMdolTpaRW5a3GPe+Qpoa9E1lK3GGahyP56sXtukcdjLeOnFcjY1FJq
STvg/i2fOyIagT4/9KVBgHvcrf4a52mAX/VK6z+K7HDN/Uf7U/W/gQeYHZA13aZC4W9X0VvXzcYT
uT1EN1Qx7Ce6jXUBRKNbnJ8EtDWBDMhTEzsw7mFYAOMqBg1Vnlpx3/fQHUQ6rmNY0yklzc5X4x2Y
dGdXobkHHkCpKRuG0EjnnN1l0qeah5S7EQCPly0RA9OBQ4KND4cv771AEFbvVoo/gvvA57huj4wL
c9/7QAfZ1AzHVxZOE8rypxorOoYFMmeG/h2124E9Ipd2mQ9epnB/1mczksBt8XhKG6AXqByNhmj0
xN8Wj2juOHYVOQLmqT0Hi7wTwXPg/yakFWKLSWKvVtlxvEzPk9qVxNOdXlivtfTm56+ML9tL7Lxa
w0q/bPV1B+6i63pulNOH84QqRdNe7iyWk0Xid1i9QhCEc9iipm4RWpfIImJA6xqAAAxMs/wNbHlr
7Ggmi6v3sbHqOlgkmjeki8CJDa9Hi8HP+MW+M4BONjI50XT2jBJs81XaoaM2WCdiexQ7zTMNJHpP
EBjWF5D/Xib9voNgTgYr6s4DfQ1NcuZ9cnce1hprPUFJw6gluUW1+PK4JRgT/SPZFhIHXXNhRM6r
GN3QFmfw49rklihiC9DxFnDldWpYJauyyE6ECxS2emG06Rxax8PAsHt8PdWx4AwwOIImgn8FmEtG
WkKZHgxg0QTqagtpvRWqVaFF9+xBinftEpEufsXfW5yVdShMen9eqgHllvKS2gAdjxtWHcjUlmJL
yrF8EUeJ9JcxoFxyKFlxiFI4ht48Nj3oykx8ELgxlBxaws66C2pmvYn1KA0e+YNmvmTsWlZo29uY
8evmubZppbCfkYdDLNF7U0Tj9Iy49Ia3sW8vfFWXHsChlZRTaH5VcDn02sAyc/7BqAA00J/i9Pcv
HSAXQ5Q6gaJRzVQriTt+Suy2LxjDGLUjPalk2wwoxlNVh0bmzbZQcuenjeqijmFn1F5pRuHfActz
9dlyG2QkwR3ACU04V0s5IjpasilOnIatUIEjEaxkUxxwRKLTvyYLbaTW4WzL4rokeVOhFzoKQjdU
mFcfjgdRfCyVDPhYMnpfw7EIBu6wwndgRHxwO90JhwhtFVS+BPUT+aeyNtU0kkV9/THGHnnVwYcG
h84Pdz9Nu8b3r/1uC+HWjbzrW5288gSZmoXVQzI309VAfUvpWv/6L+H4152Pw+C9GKFqH/EvRvJA
r+BDz6ohwfGLr/U9K6DyWZn6OrMdK2VpjHc6XONqjWoRab1ldkY+HvIOffZ4sD1vhRjWuk4ZzRPE
kktC3HrfZI9rG8olmh01tbcFhBetNFx0R9PwiolUY9NanuulJjfV5uvanyAkX9ufBAGkETBzUzob
br8ZYJ7NHEoSefeX4KK4KrHxgZ1C5Ms4Gu0xWZONzg7qixSYTXtnblAMxzlAlXCf2GVlAdjQ3Ibc
26M2b9PtJijsT0w+3Suu2f3w4pXsmvctuY3qtxRoyO6lZArnpu2r5f+ZMllljSd0LaBAUN+ILRw/
LsOpQUmCAyYwd5fbz6xjtcqjZwfDcX0du4bU3lFuRbSmxdIW13esnU7mswoLLUi8wUsJtyHTnTE1
PfFyGZvbjP+JwrwdBCZUqEX/KWazk0UlUivXLaYOhCaQ+o2IRDupTl0oexOi2MYKb4WSm636ZwFd
HttEiAS0ceAclEvWqKWErfqIJWGz29l9fQVYBYYYmqN+ajK1z2FnztHkSVoDsPWJ8Unfj03IMP/j
Sr9L+GSTpT1LixB7jsIcrCulCUpzUbfdF69ILCcvopa1yxYrBT59BHUehgLaB3hZ9QEPl1C9VTr5
BFL+Ij+nB0/fpO7JYkP7ky2pF/smJ1diN0+NEV7gwBAe+/027mG60WHp9Gm6F25syAeCh4mGPJJG
OeZ6xVO/iNTDnrMhSHNt/wZHO3usllawe68u8SKGaktMvV2SvJ7G9RxPlSZTpBkMy4SlNel661VP
RzjCPVeubbzyajP1U6O17raOz1tE0QjLqwBJ9uqu7UA6KR/8RY7OArTNzuZugEjlIMdlLsFV1yOc
datIY4zqmTdlYdsdP2p0OzBhUqjKx6nswfQSGOZGfDVi2LkpTGE0Ct6joeQ+GJR8Gcqqcl/sJ6eF
JqFBAmyzKCx6ZB6EpQzJOGTG7QiDe54PgqkTUN41jfFigPLP0NxwokVXGmEH6Luv/M0NZO7Rurex
dTexnEv6R4iZVJlXA+N/C9fGZuoBl6FgeK+q+ZF+F8iFVU2bCbgGXkTEM+TBZtjUDMQ41gM+yaq3
M8BeGAcaWwGhXzmB4asySqtUYUObYsrFdpMfoMiInKZnEHui23/53GagfOe52KegmrzDplwdR6e1
yExyzFpw4fMgJQIBn/hF2sIAt5Cpfak8f6ouOYuxTZSzJp0JOYYwQiRuASIX7BdgnmYk7MpSzhh3
FU1YV0CLqrv8GmFTmdlhbWM2c1rcb62+8lOhPXRFZAjGzvSNcKpirtGg7scWDu3RkGhFv1PPvKCE
HLQgdizAUSnGjTFUbeug0RyyKq/i6UdUz1pVQrXBjozYWFg73IH/uiJl955fRufeI+vloHuPMT1S
eBvEAWwBW4pGmTA5ijxcuLHVsnruWwtOwQrb+VAFbAILij4rt8yplRi+SwKl6aZv1EbbNGxwun6w
ReoOiIsYeZyHKOLCPDgnrQ9jAIXTmTp5dcCijLhRCPeypdIqSDQbiCw0SV4DpFwZc4xYCHsTrjVn
OE0Eg355kR64F0E85b1ur5vDckiwOIHtMFi/OwLMwnje07xmx3Mo4ack2vHD6Sh4Rt2kQPbB4A9v
rIKtevlaVDse2y/h0L9ZrpJY9AYL0GtnBh51LYyz2JqT0DaTvEHXc+HY9FRKml5Hhla7pW7Wy9sn
I/QRQVGo/vVf9yti3QfCcEVFsKOvr65FNirDkI8YxmE02B265FXej5BIinnN18cHbQ7pcLt9wpMZ
vDdqNzKlINsjQMf3VS1jUegIwbYoCX451dsC5/e0ORCrmth26SBCBK/Jn9Tgoo2LADP54+kf8mQE
XRGwAc9ntX88kxK9s3m4CbcGvbtY0gv8bzy/x9dUknKvJNhjZobhXbl+0DUytYlDKKfBEA/mrxtH
ymvnpUxoH3fViF0wrknwnfZROdb8EPfAAC9K7C9+AsYtS78A7MHL9otceg1WKODiwSZHQbWcB/ws
Ld+asrCbPBg6Fw02aDbHY35v4EgWDHCD8EBVUVuMgex1blpMRB7hBQt5BD7MaIPDAQ9ZUI6GDAqg
iVj7XA4FH8plJ9TRiEX+sF7CrfipJrau92xPjmxi3u6mmXm8O4ZSni9mqgFTK9BQ5wtzhc6Ndy8h
rFP1kSGyZNv/Dr/Hd46Y5wrnD2xLkjr3iogCbBvDKwXNLGC8q9NJ9cr9DcYfXbCO2DeQxVObTl3b
nkKB5fytuo4haTRZtRcj/NTWxlwtlHTGzevq+wBkosAp3pR9FiEWGX4ois3gwWK2YFAVCMaCFgWm
0MF2XxB8Sjl+8SDgGzwhMfR/mCWKLL++Yh89Zs6RW6Nx0qG0fZm2Utjs9FhD1tZERVFK/5P33MWK
75CzXq/qjPT7sJx19SWUcr4CGZdML5p6PH+awf0VXGDWztdqqjzh3QB6rLtGHkn9+xmz0XYF288I
y348LO2DekmEOmi9KJjxkg3ukRwExnnjsvNOC7aRgFYLApziKMMLu9groy9fR7r5ycLRpbTYmsDw
2PvYwCb3UQhXvw97k+okccAKEPManf2rcTkFcusGseEgb+n5RwqALZ+jLN0/iqRSFyS5Zm7+IxW+
dPiMVFBHa2tblvc5OfHgeh30SwioniiwTJ3EzTJ4afhT1kXguN75mVkIFOMDrJHUEo/8vWPppvCN
bUgaILxvXk6vngf4O00lwgVGtAHXfwsH7k4n/74eUIUQGw5TXRF88ftppgXOxeaKuJmRPJmgEV9Y
WpJLDexaP4f7mVdxPydHAyWM9kAcl8VnMvushuw+Vp3NL9790L0qWiCn2TDJAc2FE3Z8jhZq01eN
G/WGB4AqnbxLQ6MgFk9qlUT1jQG2qVBnYCPv3OuDsKPPk7EDP4XA+yaJ2eut1W0qR2ArcPd/yQ+d
LFJl6QkpBkWTbljyixhLJNHmuHsei0e4jVJRPRp7Bvykit6PBgGDnXOT2GUWA+6xc29Pu7dP1Rf7
e0xti62P+b2bUYCA7eKf3FHpUoO0yLHjZzOt4nJj4IbMIJzXbyXt9vkWJNvA+FNEtC1GWUGdLTq/
9gmudd7Tz8vy3uDZKHh/7g2i7dcbep9gDo8rhJKRLCupwYel/n7RpUDCmCk0BjJjP4fP7myDypU9
HLX1sYuxoohC1AD+fab6TB2FveC4rK0grSSxz4LkrLocwVge0XPgKDyFaZMm5Az1rCtDd+9ui6S/
FBK4Kp6Q7P4sZ+Lh5ncIPcl8wmqXUq0jsHaFxYKA9Yh0SBkgHq/EAN1LVuCcBDWMcFMbW0ulVudq
vKNtZDA1HGwFMJ8UuZ/NjKltUYuWoleaUcie025Xp2VirRzjHufB4qY48LQF/I0/jv7IoCwUu0kk
SrtG3mv69yd0Mv5LiT2SmhJvt5eJn/aAaP32IKgXzsfuOg03767aqtBAPWREhpFGh9IDK8w9U+vR
Kz9sFZxwDMkwGUyJWtd1Ly6Q807WCI0CHzCEr4Xkdx9aSMzror/IDR7Nnq7myZN41Hq2r96WoKGk
obI1HT16Od4w1F0p/6eIHWaW39R8sz22AMWDsl6dh4lN3rU1Q1QmFFQnUnGe151UO6vHc6ov2bQ8
GunAB7p7az7cKLlDZdmyYMtr8whI6R857hVFgJopilO6zSxYySo/E8U1FbPAZ9qphBvE8NgzoWUi
gKVJBUc7BwGvKZHMgUMZPoFUTfsFMfJdF9opivz6OaeHxa0EgaIFPUcxPUllHzeRUQTG/OC0wAoL
XFYT9GLaN/niqWmElljbE1bUZe65ytkvGxpdaZ2VMHU1TXs2xwTFcb+uBTOBAdqcMdfASz7fPkFC
u1nxvHX8lrVunuEBAVB94RIGyZ9s5YaAfsFv6g0SBngLz+JvMA7QJhnDiI6n//10g8CX2GO2Pzwv
N81Rgibgi8IAt4ZjsAoc4WF6TF2WEeZ14CfLH2uCkgmsyg9UANMSTAdRnUg7fWRflhv/S/6uTCme
9cfqwe/nu4DEWQWI0hIhhwuF5MDIUdDo9Pcs8gSce/+bBFVs3L0fO01LZz2sNbEX9JnH7HY00Zf4
Ewj1GU1/KRY1CivKWnXRioyJKq3U+y+GGQWygE5+tdZ1V7EdiD/o4MIYip/S5inC+Zqzxxm8fCde
gho/mR9sppbKQDWaW6VA5Js+O8pdCFbnrZWTnm9NIdDXs+m2BTusmhrbrBOJjLMC0rGTxEIgz2iq
6UStOJzpq7eZkuzD0Krwq6bJfkNWdVxb8kIBE+4HqyZH9zvdNlEYg7iymZqNYJo3//Zzr5/S+CB8
obRcNUmXpUFrQQLlgP2GR1S1B7rEdUE3HULa6EWV92VOtK1lXotrJXWk9Qkfc0lXBsmioFQfDYJm
MrrClo8GPbYwwQE2mGft4rRj8jR2XU9s7yBC6joTJ92lN07kDwcUpApTHEYycET5ZoT+/Fiykb6e
bcD/wquTLcSQHNPwrmqIOiGH4SJjMmWn3pLPrAyqgWS+3fqczZatoqBOx9X4sGLwc1quxZnarOlT
8wPkKmOc5a0MCgDewbrmJueDgs/x/X57PTIQboqc121LT3jyV6zosP5+PDYDgdbyI0snIgCOMqeg
jGfFs5LkLF6fUHF6FobWqkZmNwcJC7/70aJ9fCGJ5ZUZIboV76YewVZ528X7hCcnnyjgWnhqq4r1
RsHa8W/Or8drjxoGFL4svj+hcPDfPFKRLvq1vC36pg+dWwLCGOA07gtELieRbUcYdrzgLh2w6q6/
NiEsGAWr0FNSfWtfiZD+4qu7Z/lL/XDi09IirWRxLulv62miiwmM9DMRXoVd0QujxAUlhmdiEl8I
UVfTemwZ6YoZE8CNOg72muz21+x6BvhSD+MsjOiVBwvEJnis/O6A8aYXzx137WUG6Fv4uKUNYtVY
xE8gomxYIqZHkHwP8LYjT7GnATf0wk4lkNQQ60EJnVqBj45riqq7NBZ+b7Sn0wPh9/zxleRDdz0G
yOzj0qhjmozJbAtR6px3WyFcAa8f3dAs8WdGX+a8GyHjdd69wIVZSbuSpTt7VQWuNVR1lL2SJtK5
Y+6rJ1R/9fcVQvfR6zq0niwEM5XflR4ROhPeS+56xz92Vf/XIQymuyJ1pqXRR21vNsS9bjXFyYj7
vV5g0ujrQ9KNQ6hDp/MhH8hlsUlHmhG7SEqpVWM4JuhvYpSh1I+zqYf37Nq33wH7xdN6eTiPgRul
bWYTILwifenrhrYdEvhrUZqydfEv61iq1vae3fb7ptd1ODbCedIk71UbRQX56ZfgDYXPDqvaLh9g
+tz7vbw2z+ADG3SDbNhhII/I6wt62+fsjU4LKs0TPLf7H/ox9gx5wTU+6bD10UBfHMJJdp5PeW/h
1aiFyHN9uJa4Gby1l4u/yu3jhrZNOBpdPz0lQ9UoRuStIoorzpZb8XanaeY1pA/ojckPvBvCBM4X
HwikCE9iQ64g+yfdOGmnECuyDFN2oQ6sfvcqH0Fz6zL/TLiDAYEl/fHhNX5zslNGGfldNfmIQjJT
snrsuTZaxrAO3tRPii3mSYKrwYA/H9aZ11I5j3cAaoMHn8qif0Jjk4DpS+7uygYRCN9fvYXinfur
Z/bFdjDCpAtDsZmve78o8p3fDUrnpSxOL1KtM9uqf+GYUCDHoRYj8Sm3HyrETJ0wlRJlBBmVt9vn
rUxhZAAs5ap+/UDXK/qWlHT+7hfqiC7wcwafp1RpMEB6cOCjxw9rjZelLZyw+HgnjjMl7xP0c6L0
lTqcES3m4aiy8goiAP4F3sg1csDc5p7tT5WSeVn30JBN4EHG7eFIl0utS2mufFX4TiJwrN5fMmPe
9v1RUSj1sfVxQmc77EOEetgA0D2HvliodsW5tV3nvgOKk/tiT4UMmxtfraD6dtsMdeIJKQMmsl5+
/fT71///n1USuwQyah+Jc6fkCP6lye7WVZA+8vM/NN7DaTCslGkA7goJvDInea08bIzRQdeR+kSj
EuJ0zl7WfrEug+jj4VDtgO9t6/9JOcsemWbMAshS6Rwk1nP1xy+gNdb5NnRz/OL6kEFH+4f6E3YN
s7At4kzVZPeiJHqyBD13AnQQaa2kkcQACFIl5xZfZRxf+RyZPZWF6AV1Up4b4ueMrd7QthcSpzXX
foO5zlLsLVKihOaQlI55lQVQAB89hLDvz3wb0Y3MB9l6FlACbd2DQNb0rC7pn0NoAonAzDLav7pD
T5/cw1UAg2K73YwiLxL94lKKBPQ0cVFWWjGCrH7etUU4JaCXqpIsR37ARSzmFZ+07L/LSinEmGuS
GsRQdyDQcPAa8ubjL6bTV5LVWfOKapowwJE70ztrxOveY1gDZMgiTKuZQSUdWdWG9z1DktmiuIoW
JLzZPXTiVr01haJs+7xwZc7OXl4LK4HGr8X6wyzDzVmXklJf0i24iI6dCvBekf+kjnnwLsqGlScB
PQc9/s15B8KbMEtRmOV/lc2hPr000zxoR6HoYNuCJUjOmLJAbDeQJ6M+6Ku4aiiVXkMYP0vlLoLJ
+mKxkEjv9xrBt1T2YwSyI9qbMf8e8/Uimv8766F2mL3j1HwlZZSbdZYpoHqIfbppwvq0p4K1N/1T
1Vo8T6ZbblK5wzL06FJ+ZJvD3Nc097ZvSb/N+iUQRmt9TPASIuOwRUso1Q8ZdXcmIu94HjoHH8HY
7T3S3BQ6jjxwqrDpXeNefl2ZAUff29tMwMs6TZtg7eY/YtwGsO23SjGShVV8G9CCgtyS0oubvRM0
Bp9oWtHZfmrnOAjv6oIly6T/YRG7Ms18SCArTcW6X7Ljl+NM+tvATwOznTB23de9b7xHZ6xCbInn
A9Isdl0V12nL19PbOB7Vv/F37xtsu+XBxc8z5bW0MhpKpcYMP+/u6WBqkcQOnHyFsgKvWUXkSaIr
8GzmR/ykEE1ffMWn6p3gtlCYEAV4STJNMUcm+bpP8Owtb0BaWiCtn9C1O1myJrL9or7M65cBAB5s
I0r6aMgH0oAL7+f7FodjiekAgf9feAGjWTIalAPh7O8g+USbT82EiQV5Dows1Rr/nRlJm+QtT/q8
aUISihQppLSe3klPXUHq8nbzadWIyeCxzqy32EAvdAvyikgRy8pyF4M9lCFx/XnmlzcmKfQ4s8f9
9/llwZRv8uT3mA0TZeIg0HX2bT60Pa5HaBzsqWGVj9Jzz/tFePl1bR1tFN2HwPP0tffu6LacGgDM
CrvuFTBEO1L4sQPxNv4POZ+831fA0yjXOvcvY+07hcNEZanS9HG7+WMTSYLsnqUwNhpT+W5FY7BU
j3ng4cs+3iRLNFwzQpY4mMX5qTK5dssUwW6zp79/SJCabgysTecip2cF/x5YmjDs8gO/+X70b3MU
d2+qtnf95TPOknoNyxo+TIB4g4cssHoyZxx7NFmdV9N2tgirYBkxSvNTfeQ0SfWklbtForxmVu69
+tTeyo8F3SOw4DMKUBvgEAFfhewr6h0a4yzuAToKZLazd7lUsEr2HB2UjRmWAEYcKABh+b3FCl9f
1M9hoyA8ytPDlCMd68bcuLGKMk9oVmVOJUrF61qnsEJKyy/bwrNRoqr3gTHN4St1kDC+dx24g7N8
8QhmQeZNcdLLYJQ2XxAgzHIf2DUWHGX+rCb/BmHymQG537XcgYOTXF5wNLR9/iabt90DogX72nFG
iKP5T2V+Ht2E82ahkDxJIiBAEODQTAtDsde+tigrhgwmocLC4z8rgoWAWKJg2drCE0Rc26ny/7hq
m3Vl3HM7hnVh+MsTmTCR/CNekTIsiPHUJmiFMBNn5XY2jDDzzipm1wQ85uw4dQuHivyj/fywSTKd
+onGPrC4rxvEpszS6UnzrkdNgIoKPJuNh0/6u7LYXUzN5PdQAd4hVtntRFAmnaG3a+GLmlY9aITz
epi11ULbmP+PpIQqdtPbgA4CAIe7ZMq44L/NrK+bT5IETndLxF5VmNV1pVIcPovQ3c8mGB/6ovkK
2XVYMoe7WZzlg2xljOWGujpq15s/OAv9NQOSaCX1R7G/SRYQjAJ2ZAQW1mJMW8A6gxt24jvIifu5
GhH5PaKPKeRrmgv0h0jShp/gsLv9jY3cUtJwFKeYbS9y9EY49q9sAkP1fDdpp6BVxVaQPaj/1nVN
L1bS3E3HGTfvU9mL/DgsH9G1iykDMM7m95OeeWRP5aHdDYeePZoL5X6QjIeFMfjWqgwHRD4H/Kj2
aEwpMVt8Qns5Y63b8GDK4pmNmcEkO/P2R1n/WCHYCBaPSn7nClNsqvVD6pJ67C1QD6KyvFQ3hqyh
R/5TglUzPHcNtP2EJ8YQwHpCeF1Z3INr8Su4a4i2VYHunlM/p2MKocgZRlEGjQI0jvWy/Nzd0Jkz
6/wJhrYSDJ1OnKIyu+O1G9wcuNTyIvAlLnYGWjWJx0XkUZkB0F7Pm3ViaflkJvSZm0XgXutDGRui
JJ65TUEkaxPbAh5qfHlUdQPDITuuYCa+MCJGQkU7/L5avWsx11R2W/TkV+Jve3CDZXn8ABIShW5/
ylloRZDeSUySRqEw3kdr0urRU0xU1LQtL6fQGqGuHKd1B/yqFEN/KRduSlNtJjS7k/dG+fn6GQKm
SYFc1f8MiVJO/li1cPI+GnGwAD7EtWsHv08U/CN9yTUqSDS7/R7hAawCprhgpexoj4/H8d+gBHvZ
lLwa1Q/TfMvIUPuAA6+kkxf6m0lIBPHtPOCj/0h46xJi0BPV3WuhJXqHCzan3QTqmZPv2BpaMhDz
4nN3RjSFiryzrwSjJYhXj1X+/K96FTQxwrOZEAIthi068SYiZ0czaM9k9o8S/JemIcXiXnSKOsxC
rW4kg+0wrGijcgvrl+5vRbQ11R6vo0IBeZ6SQpenuzLL3liY5BqWOvK+jQaU7dDF53VMZ9A4U8Wd
B01BUz+5xQJoHCDtLvkruaa16E8o8iAl50xghqVHnd2L3qpLizdQUSS9dztodYWJdSMT3WSv0vvt
RQLfcBePQUgSURsllC5dkW2kIAeiSkl8G6xLQfDouLzdt2kk7N4DPJpTgjql2Pe5K9jdbpVhn+4S
ebwiiX06sGhBpo7Reyncrck0jKlGt9IAxoVTtjkcRFxZmZ/NUcpZhkQvm2bDwdGtjdjDiozyTN1A
jtvB5ziuzcArZUp2okPoOsTA2fJyVJNrsn6/2qFJI5vo7ieZbfsbHB9wfHCv2XoCYW/benw4RjS3
/sEfge9facMvZ+7CLLVw1+Fb8rgLdT8SWIbztE+34bMRiYwrHcJAOs+i/xecpILVUGiyoRNi4936
RDfQV5dTCgFZtRfhuGTXrLWTNdRWkZWNB99NgR54v1hTFwe90NsAe0IUZ61YUMw05XRXOe9B48sN
DcaouD2OvfG/jHoTZC6THbEL+ACm3uVwE8OLjJAXS1GdTGu37IT+DJOWOfqAZQGAK8hDPiFFcKGg
qna1EvdguKGOhbFJR2Rwog+uNzeUeFqruBw5Zepn9EnveE8PF1p/HybENzOcF3xbZPQNBL1cZtx9
mcx0NIvRHFsKjESw3y8/OVIZ2um9JsgS7dy457NLYJMO+hEvYIAYt22r9QcHnaCINWPM/P37X6mE
tq+1YipaW8ya8diN0iAz/TSj8wrk1tQE2JWgfQ9ptg3V7zbKQ1De4VBryBWn9Pau0QWZIeAEdNJa
dnzuREG2vw2Q7M0rJX9867o1dqJ+m3ELSisgr4ExuIWW8Fprzq2/aYoE/tAPwrtqdYfebxHdkEX7
i570E9AvH4gfYSyy316RCCwlKQMX3K7Z+IVGoCb1FsDpt2Ty/EF5VYtAj6fxNrreRva0whU1KrsR
DH7DOgCLqJFlDBXoqGJgA9E59J1m+wt61lYvZPCoKN2Qn9qPE2sCF8LLRvLqc9HxaIs4ZVo4Tl4D
oUYMlNdoW7b4DyiZaaVSQUMwnx+XCPXvVmv3FDWJpZYRS3g+yo7etDZiR9NWUVyVXQbW5kJInafn
rAtiVUcjwVF5ETIhwZDI5f+ctDtrYd0hXaW+rwI8x6WWFO9+Q7oLmiULpmSKwMJzFcTom4hRGP5Z
qHoQ1f6xzvV8FPOmD6xx9JovYGsAsltF1wt2XJpfPgvt+o74v9DMy4DgmsjWSUl8WoCFCHaUzEgX
Sus33h7eH0b50oy88El4TntUVW/JQyboWyzvyCC7vFgnJ5naQOPZAvM99nxnhMjl3GalBiFImgSf
r65vgBrju+aCtGWi4CXNj3YAnltJgxWQEQAvnJueRs1ul9p7lNrL5B61TcDfhqVqHAdOSg1/6zVU
9tPtTYMWZ4wOpYvEhhyxkdnc/ExeAz79etuwpznC8DZeMjbbugNVLO5xv4Cz/orSttUdBU8kY8/d
Vw4qQKYWjTbq/0eswd5WfCgh3fbyIaoUFttUEGr9OxGfKLAp7Urq4PyQqNub45/lH4rU6z3/oejI
CpUV+MMXXnFFnXBZROkZCoyOPMhyvX7kD3a1lzrRXHR/VtyxgRfTLs23vk54PKEn9gVTzbS9D1xH
vd2/uiVbq688hZWE01Jm3xyQF2otdZaxfB770M/RGdVX0oG/L9f4mVhHEknWxdKH3z4XM2FW6a4Z
QvTs8ibYbjct6qy76hPuuOT3gppelVQGOil0hyNkcTfuhB5dFgsfwhavR8DkPpSe3FEHDGkHy0BR
7MGBOMO50OTqPmTVnq9TEfu+WcAsIodTKVdZxYzwCvpPrxriNBvGQ0s9U1n34LN4z+OWXxD3Cf8Y
tdc2XAJyd92Q6QLYcJPbvGic6ExezjBef0SYnRmaO7P/AMDqi6XaUnswhL+glwSLAfkL53yzsHCV
RHWc5b1eGDBEAEq46M5pC3cqfp14AnqFH0R6QIrGvC86JqQRwQ2OVVgTlS9R4Ch3GM9tRuunp4vz
vIyi/Z6UCcEBp0d14BHiQWF+8/1pMJf15XaNOPuyr2yTxBxUyJluo1Dha+rfqYUP+KPTaQKnFJHH
MO3MsvDqxibhJAp14XnNi7AEwjgcKzyph7VFQsJFLHp+zi3NtAPCMubaA5X1Pi9PvqYsA6V93MxS
BjimnByAvUECVQkLdnfWcYTM94qDL9Esq/Fq+fWUNMqDiINvc0bCXemZx5BtBTgJuixn+2nwZRbT
JGsIzHaJaZ4D7buNoiWWezcM/UehrthbRzy0qIFj78/OxarBb9a0aJh3GBUFnOFzsfKqkcZc3UgC
4ScsvkSxZmTX0AOp7mOB5FUw+ac3GXXz7cAEw2g/UH/v68JPUEB0Y59AcopTh0e42/pEo79VeLTl
3jTzzXUosYQ+a1zE3ydyZJaxnikYZkIXALXn0BiBST72JXj1gDpwyVKsfI0fvg6KVGKsW5+0xep8
gNXCQRwa7y6RncrpjC0RfjhNoYwHTW1xxS9gStftSV2GI4c9MxxX/Twt5ZQPjLLE2wCPA5bUUMXn
r/mlpSGD/otA7Go6u4RKyXDy5sFnD7fACs2+LK6QUMmM+mUFWZqI9FNfAkwzjtA7Nv+ACXC1rgFW
4SGi0Uwi/H+9Mx+XxOjRIRBW5NbyHlfjjcFnZbB1WO+0wO6KSVD2kw+BP4hN4I7IbuLQjJww0TbC
mBJv4Ccj5a2mFgZvVRJs4lBYLusVfPrCahXuA+pNa0ZzE2glA/l+q6TxkQYTmnB77A0cgA8hQQPK
00KY9jfc8WfSwY4UW3yZY0i8qq48D6eVJkBZeRk+ktLkgz2QOvs3IZHPSzhmAKjHzd9M07zpIwYP
tgDXYz/Nc860Iy49C3Q4fWHkJZxotafclH/bI1GnMJfls7bF+R7dqq4TmA+yoMnr6sddt0OGRFT5
LJzrYqijeLX65THJbZiDVUQITOmUiBlc7kqYc5ERKwYUrsnQJL7mgSjfUL6629QKB+YA9DckwN1E
cDPZAZXufMA0Ft3yKoDPzHeJCBZB08/OC+sb1mWIwZaKtR7MW2R3EWiQfmJtrIcws6R0mEONS8nj
fS31G7yGEUOZUm7Q02A7GbZIBzHLtEniOHnQ9AAewK9Xp5oQBLA1olB74+or5L7XfmqBqqMEtN7B
eJ2t7HxWrR9OsR9F9+uYjo4nS0q0h0Ta81z2Vr5lrNt7ccbGQ4j+4o+wQSponKRW70tm1BVzCxij
qHZPZhBNPf1ehs9zeocxS6dlbSkbi7zCE7mg7w9CTTELoY5maA5TM0rEqptmsNodav8cHhRzRRlf
+vULDHD4M8YYIrJgg900xT5SHK1TZP5DOvZgfkWa+IjGWcMzU2uLIUZDS2nfroGqKVr9llhqKt+a
7vug3tarMcsIysSUeDXrImaRMu8lxEMp3b/+zPz2nZ6P4SB8YEw4cSg1es942aSrqfNEmTzvmfB4
+S/sqD5HK6Zb45cJTRI4lPGCxgTrmT5ypXwaQZ/PM0AfNP9UMezdKEju7hbtm/bPoSEgITgHEQCw
9O4jN+XwKoeeTy15ZwrfJT67TwPb33H2LQxseJXvputzK8b7bkxWp1Qlc7Wuks7EQRqVGjGjWNgJ
za+E9WzEg4MwAXipXYDYIjpsXXIQBrEhS4OyW9nJVL7hTeEOK2e/NbWGq077L6U1EkaA9NUBf8tt
uDj4eQEj6qu9mfLH2aE1egxttqnh2EmIbv3uGEuHdtIMjnIlTq1fmEydqcVmRMOo64ulZyIX71EZ
QV6tgLuteKEbSUUpwSV22IBq5ZnDvh0L33b6/KA9Ae7AtzT6jsuwA8FbzZ9dWfpaESMwutnGtxlO
Ke2dtDDjow1iuHLQoprPAJbZhGFwaCni6AENOx43YlZz6+KWtpSTL+s9E0nuS/EE6DFk5u4FqIv0
2XhZIJIbT8u3OrRQgoApBp/JV5YjwY5amSs/lNNhfuMH5TXJqGPczrVYNutwo2j1ay9o/TEBm7jW
G2h3yovHng2rkBVLEhX4ETihYX6v921bxuDY9to03M2n7fpTAQBmisrXNgwfMqg8kF3QuuoWOijb
kShxRPzInKjZM7Ifvpkfr7bJ8UO0HCYlSboYhxr8k8AIgbZmH6UdSlTuPZPmmnaU5ukWDkqGwgFF
JB6rQFH5CIlX8ajYNfPh49FBF+bK6j+JNxOvhUuKkMH6nggsxZsxv8VD8EVeq4PNsNYeduCMjfm/
ny3M/vBLgyE/uCiHKEz3u55QqSI4tCIuSpKLfMIjpyyvhU8B1QkzjMz1duowZRV6pGuJknDtAHVg
kDuTlJEuFSQBi7w0brhG8vwVMzTQRt6ekzo952ungXt8Ajb6A0c+i80fGhnJFZJR3Cn9CMrmxQ1n
ZYyZEzGf+7AjXgRKepQDOdYmExdllvUjGC4P0a0OLK0mKxIsOvzBGKrPYlHkIAcOMBIHFlcTM0A/
uk5ckeCHukA0yJsuSEMtyYh/8fnLhxSkEb0SBtULmabzhhCSVSbjsuc5x3heLOUVed3U6fdHPaBK
Jr2zjkdf/4UEJAF7BxWndp9mRLvKpx1euMI8oLc9Vj82/xCTbZ4qYfGSFwx89cntZOwYifpT8UTV
Ni6G9mWkFnLbVgaKh1mK0DlMXSFar2yJ32u2WGq/Bj6kGpPN9E75AzXO8zG7j8jELbkkweO+opL4
pQGyic9mkZ0ZUD9pF4p1Za2rCRPV8W78pPa8FqbKeHS/u/fiG6vkQjEJeo3hl/fUzs+a7UFDoCt/
0f2Nod3rn7nzIP268Dv3BsrVgq2SW+e6EjU/YGS5PftXa7NT5Rcw8tM2QCvRkRAiLyT0mxp1zfes
q6KO0AafNsrvi5ZB1rtiE9/uP37jp6woWczhccikS94GWM6OmJ8ZGyNk8GtGD6DLp1aB0gRqwPUr
BQrJefzoJDCkoQ4xMuE+J3Kh/8suy64JnLMx7ESHFFy4d23u6wdR0rXtJUpeS0LWRQvhn5axRsPc
5DHUhDko7EmHC6ptk3Z7nvM8BZXS8vnGvQfT4O8pnBOHM1crqz611ZKfoggw+v6UQEEsYjCeIFj2
Mm1KHAraTS4/1VKziTsZ21XbCmSJio79z1p2HX/mlbvO16nR47DwLjgJsb5KLU+SLWxgW0lvkqZF
JGH+Bj7ak3BKmfPIWwwykGvfDq3+rDfJVYrfqaAc6L6eXK/e2pPOIUo6F0x/vekex1NBDa1yeZe3
FCwX+nlWGnNKhM/Iuoa+u5tbqXF3S6Dni9hcQkg4uvqEOldPgFVhWid0xtMWjHJTnZe78n7Zrupk
Snd7qEshCrr+Hz8PeblTp8rKBGJgRAagffn7bnimhpPx9vJS6VIcgs79fZihwNpK8oQ31/4YONd4
NkA9B/kL1I8RrHkIduuyQULyJhNGw2k6fAtBo8Ojx4z/Pj0OGfFQE8vayKMTCZkGEilcw8UdHOwA
OfyaWQVf95dPzkQq46ib13f9BEWGTTT7hTapJCd8KZEJWKFzgA8IK11YxPD9gMfDOIdRTJ5LK7jM
EciQ7gFXyPdpnSbpMmWM1XKVDcSXiYGHk19TLzOCq9z1gORAyOng/MosWIeBYkmKMktCeiArWWXs
gKG498h97cqx2rd+8KIrCYci2AW8UQky+N68HKzI7ySNp5qMXljcz2rJ6x4aATg4KfRkdwew7CRH
93Kae9BtKm0rWNP8LW1a9m+lo/BYCZO+ksWJL/6TQ7hBeGSxJTDxZFG1V4Fc9y4iEoIfceIgDBAE
WGMHjGttGozuo0l+lx8UTGrXFYTbXhs0a/Ew4D7BBXSCADyR9tZ0qvLyTsarpoL+1hgoU0niNes7
TafDdZP5rSBem3jxYBKvbh7HVT9ufv1FKH0OetnjZ2ehy9mNw5ZkLtbkmRMTcaZw0LciyWt7xza+
/8hMzsWzQwQoUzgSWthRkRdewAuOpOy1B6xuezBiIDPUzr8A9839bSXXBTxCUZmMd+aF4S3xPoIa
4cqOEtOvM5/WpLZjZ2zymercxNjhV1TRb8CzNZOCuwFsnnIr/BDSo2RC+0eH5B+ryqw8fyTtJUHQ
4qg2a504EqwGKrK6yrexcBGbXqhxlhMstIPMr7J2/s36TN9dqi9soGwj5JRqkBR2y1zzJg2FItll
o9d5j8MEs15Wixi8FyMk1M0hh/PN3ESz89fkXWvSKhA8neqg27JTSZn+J9+GeSzX2NM/utUHPV0q
OAGE3S69HEptuXsf+OTtv/MVh2BqBYTH17gKQrmGiX9XVP81XvtCIicBTxAGP2Ho0RS8PqUEs/tn
nqEopHY52qAjGwMHqRjUR7aBjJjE1zRAoiW69WNhuhOq/Hiu+bpz7WACCKaMxaz4WWYV8/MsGnm2
cDq2FgebRHCVICezKHxmEWdD84vX8W2XzP2nDCZQjOU7/HBeerJMeWEFqiPzOAkgnBvjyXvvGl0g
hIezKyFbBAizYVu4p59zTbwpd4iyuTIGGF9JCMQtjJTb05x8XKa3+tmKXMaBIH2LAWnZM/vKUZ3a
hBYz/qTyWXVr7iKsJHp4tGXTN56oXzetBTWADn6SKBjqLR2z0bxiojX3e8LKRawtw7y+ZXqpaO+J
MZo8oX4txeVkUaJ9yH7uotTcTWrnDLVmLfQGYnzP5868f3xt5Nc0O4Bj0/wYy1BqGRL8IZ0dObtf
LMQuHLf3SRy4pC9AsKls0wF1pkwCGEGusxAQzOdQKvwUH+53vytfg/ZeDDlCRngvGPGpxM4eQeKK
Ck4jWW53fBe6KWqYKDB6PRGesD5HZ0Svw/UsCCG7rvUoQY8ft/g983ZKV1l1O4hiimCvgZc3mpTu
zhaOwp3NipaRIZlqqFnP4dzoGb4UFbI26DXobnr9k6CzBYbMhKM6tZCvbIansBIC6v9YNwWbckHK
5EfjIvPu5q28nuIjF54Vcl4jCH8ZrZHOaFkdsZpCZhTLJfF3RoXvIjsXR0bZtNV8902WIYHr14yd
NbAHvKvJLMYIERyl1HytYm+7YxGpRd+qqE/5C8fR723U1zoCIDi5jMjpvougLnO8YYihllgaZjn8
BvtYgEgRvzFf+xPkd/FlBiZDvk1HmqT85Z5AIfjo3gd6wzP8dpa/H5f1ceYi77YAGFrmkJVhqBbz
HJ/W6q3Xf7hszYcRUZu25sUyqsQGRb/CZQR0U2hQYvGOic6ncV2kkcNDGc/RJr4PpuXd0ilaSbeR
MQk50McquMwNlWVZxTlIZSCG9G5tWyQmc+yYzVXkX7oYp0N1AwDblzx7cy641DEgtarXPGDWkyVQ
cdfkV4It5uZbo9MUsmo1lZrkx9/r6/vs12LPBRZyke9mrGA4AQHvsyWnx8q4zJKcW6x3RUvycokP
RToHz/72KBZeczzgnHL4x5oXmcyLMFm5JA5XahGI5BRDX/naFep+auTGtbs70yctbAB5IZor3Whh
RpGsikTjmun+YsHeqoLyJ9MG6nkQiMNrS5y4SzCGp6G5bCMjyDzMTIazg/TIy/wR+zhyqhfF/FZ+
T6DVsEllLyo+BTgAwRKcdzenqK+zhKdS2PUy30rpvb9q6dG3AbpE0rsXKdvBKRbDw8ITVAjl62ZL
sXG2EWVV9uoZ9u6PHLwjrwO7F9EFCMt/5Zv5pQmouEa+9eeAnavnuiuvzCil8jPov/pTNWuAlE9T
EFrk05LDnrhO6ueG8/LDtBsnqgtbMOeP4qgakXTCjJXOnbhuwUwXOx+Ugfu5T+QuLC74VwLFiSsD
5eXcAkvx8rrkQZpBf/ll2+geiV4AIzsAadeTnvbWChUY0AQNtIguvT3MWO97jyyHBdWtATFFSiYI
zT8OG5fPVLvWTP5tH6Gz7I9/lc0/9D7KwI6NEmyOYiSpDXEAONLGegicPqN1Jrektq8qoPwxztgK
XErz9YTZwowE6Id0v0gLqguNTTbF4OKicVWf+saUUZfnVseBfBKxkdocH8BWYwZcswJ+sd/Eyq0s
EYRcekR6XUyYtxqcQtzVtow5D+ltEg+AMEPA+Lrw5cXvE3YYTJpjn1k6RGC7UpW4zoLWNIP1q8tu
No79EplsmgiRWlOHrjQ4AcS+AsPdWm2Ot+7a3CKp76n5jMXnwJntoKun5CycjjoLB/a6jrkdpg1D
oZNP9oPw6Be+DmXR9mpH9E5YQuSxJqLBqaOtlWOxijrbRA1/CdgOzkMGBIn3QuSEcaBaL4crjE9X
q1zNQVeG2zbw4Rnt6RGcXuR+8CD4ezOiflwki3cogI057lLOM9TF5aUxDTUAZNQ5aBq5AipwqlGm
/JDCJ691k3Ddv+1dALk5ZR+2D6YYrarxRHSWzFZFHB6ykk6F2Eax9B4L+MZXmVXRpkDE50YOw/ZX
1Al7fOSSj0G9WkPVrt36bqAAhZ1JsWOpCm0LYxb/z720qeLUWWuK/rBO4Gi4b922TRay1QbNYYio
U8PVgPeFqe0gTioiGf0xiYvEtcohA0WBeY5M1DQYchLhVpkMF5/YYHSVjoNdSgRKuYr3rrExN0GS
ZPggo8GzypNncnyk9BLj8GH8oDuGs3LSlWt3tSEcItT19UL+CGg1r6LYHVIPwF1OXkUQvSBDJqkQ
rstidKG4x2rS/3zuZoO3BepHMLK0lmdyb55JXaeuQF5dh0KLpODyX8F2S+3ALyHiFE25HnsvedNB
P3U5Q9ibfQ1O71UXNh/vXwQDSHDb9shNFCrsN/hzf9y2RKJBwFvVGLu2TXT5T+gHJKLNPx03Eurh
ZiKeD7PU4J3HK4RVXY08Z9fEqTo3nGj4sLhjegI6m9zLZRlQ3kxTLizZgukPSzaMCJ2544UTepik
n5y7LeUbfwnEDSOOtwOrA8db7U/H3MXJ2uTltEnNzQQDGiopR/DzySIwTVGOYUUFM/NBxj21Hnye
Ub6vcDMXkPl7RBc1KYHf4lW0StkHvltMNlWHpNZeMQO9IaT/WEHYj5u562CvmPnLyOIk3CnhvTa3
TJcYp0lEm7VIzWEbB05pEekfEKz35l8jXtzZSBvHxAt6tlpFIC2C/tAWOAxOjzNoTBbBl35sGqIj
Zo7HkYL0oz9ahwBlLywO0hHdwtfd4HKa3fvILZl/snwp8CfZbB/xQAkDT3tIu1zc+fqKuIstXFcv
IMxQB48cSU2l6NrY3RwchhhAgeQmlqqqWVYYN2a/lZTkP3CJkDMDgC1dffHbTRnvRPVTRMRvUr2C
/r49IkOZM3JK1MfGOErcEZ7YGZkZxfnTeSZlzsaUlvrjM3jyLAgUZeoSHGLOvUYtSL5skQq9Isvy
KLB2JGl035mghKGwtsCm9GlEQy72jpCRvZTcsz7ZvRlVImZPtzW5U/pnUb2KfhFqjwIbCKky9t2G
ue+eHg12inB2LHxQu+zuem366/T1kv4bJ0Ci3OAQPcXf+K3eq1+AzWuIiH8+DBjeAes1bDjSloVs
VHgDcU71I0qp+RxNL5xlf5TdTD7GqT3emTAZkIOAlAWzqMY/o9z7WQZKdyO5h7B9lMtzIE9jHidx
iasbpniBLnbUutWML37hVdgUAkNbv7A54VUmiBGrzS1GdqnuRvNX+1ZWGDR/dHhaGMzYMy2qg3su
Wv0pWkT/7K950zyAPDx49ZbElQc4VefkMn5K6F9Wcnlo8bL7iclxsJMuiVxHw2fZIt86OYKZdhMI
YfiDL4iDYAKb0uilbBYmpJD7WITieJd9ipFU64spQgo/hpYgUg11RKnJvNqMvuFjNsxP9EVr9vKc
mFi5haByU4Gqa/RQAvl7AmihneuOX37AXVMQXvogO/Hit5dAMdoUnlR4RRA6A6eLKZvkRR+9BD5m
+Uzfb/IDDAa7AJ5IK80sbvxCb53RYIPG8UP7LC9JfxMNSHglaixS3R5BfU5QpZ4K99IB+YuI4N33
tq95up5rLWNtC5ykYLzysR6SxO3f3Iyask003qxEfY2HXfM56bGNSmIfNGvlYCRHsHQM3QHDmOxT
PwYKx4aA7g8+Pn6NnMxFehbosRObRnPZpn21pHbyS8Y0G5mjLFlaiaDiEztC0XdYhOecpkuQjB5Q
9L4ZOVQqEdFcazPDzk4om5L+yiH5UB64y1YaYGL16gDZAD2KOJC7qkz1flXQROw4DV91BThuvD4d
AgZy/3RLHddu/XLegAapKMs4vSU2kzssZiepIY9DTsxYuZglunLV+LljdmwtG61pDdpkw64tB3ju
JOCmdezi66YPbaduhHuIKULG2c9/24b9C5oFuKpwobc2ZAGDH1YlRzS794NkdhFcx9RaOLHauaQt
sOnxhtncD5V6cyVRjWTjqsZCbwZSIUboTjF+Frn5+0HewAumxtozkm7IUHUzgzSR2UsyzC9mxCks
+PwjRtVpYj9PHYIGRBgv6zRnpPg+7aMx81EGaIVyu9Xy5ZfZDkbPBH6XIOacQuHTV84DDDOaTkAs
evb0C7Bg67JTCPuRzDTyCLF5ko8+ZdtnFWKtgnTgKfV2qTnCTgkktgxzfjyhU6vYorMfcrJXyQFI
AvP0uPxv8S1kIlXKgJeyRysNitgb5y7NZG0Mi3X4Av4rq+12edrpvnV7jE2N3rh4OHCv38DSJGyz
dPGWlCzkO0ypR0hQh5NZlFVzj9cI1d7U42E+G+HeITSmD5OtQrTZIwQrjvXA8w8bwkueV/WrEwdu
1uTlI4R3tBlEJm1QWCaDTolE0Fh0w0CnJULFlQ3VsxtfH4I7r5BFoh++WtzAqlje6RhwmOGVHNux
XDf2U5Qk114uW5rN3ZbwymLQG/RTPaOvwoUdX4cW2r/WbpMUkYYSuedGBF4pSWtN7gKYZGA/FMoo
NPCK6dgXqRXXbxz8T+6tCivdJE1wsLxJXqmn4Qx20VhOoOojT8cFWgOEE33zUttbmK10u1NAqlpf
XhFw10x1NCvHK7TgFH8F31Oh0TI19+9/Mpsqg8vFMepMF/fIwvVTGIaF8CsGJctZ9IJPY6XgZN6o
Uk9fWbTrNrbEvVSEBR+rRDPG1jNOVxMkFYIsP3FeKkm//C5u/kvVEZAXFsigQK8fl2N6eQsnn1sN
PTo5SeQ838bNwNasl60NjzdGvmxq3gYBMx9Swj38YTK2FP8ei/32by9vWogCgsJaAoTguKNl8eZO
HDXzUzHca6ut0Wqj2IkF0ru16cW4xuQawYdOFGbVkOrnbft0m7usutMR4DnJh4OhQnSZYEysl54F
f87FMD5Nn79YKS3hNXgo664r0gNg3d3dEyRg3QL/fOJHklC4/sX9IIh0QS3jsRiHi8C9Oqv212TZ
801pbYIrnwzkxgD8rkJRDTWBnREBeQrckyEgMyIADlv46qO6dpC7EJ4tvcC6aVLipPlNTzPW/8R1
PPYtW+8wo0wHZYVSRaI3YWTKyBsJG+ZkNmiw+AdpTz2+X9uF5PEtzcekWj9P1r4nOJW8zgLZ6cB5
BRXoULnnMXcIs1j9Pd+ETqh1aCAyKfXpVAPGdsXrzi9taxjibM0frV3yYEwLFKHc8x8d3Ps2tdKG
2SkYx8pACb16F3sOvxPR+PKUX6ge2pkMoRodGBKjHvS0BGeV77qekbLvxSCDzGiDmUSECiuNb850
lrXoocZsdKLh0CvIb8t30+/+EhYvkcwIBHR594v1ushuCSJQBfI9XDTlVfR+v2ha+n2Lg5n7kPka
4nonL2sc70nF/vAIhyhAikxDa9m4mp93uUdSJ/Zoxqy2og2M/qdS+kQmxJR5umLuHoGwHYhjurHJ
mz5Ey7vfRrdCT/tCvmIOAaRMoZBU8p30zzSn9F8VNAenq93hQwpLOCJ9kWdZXJJMJDTdRG0FmVDe
6DVT7UZnmNU4TltPmYAOnzXC1R0KWfL55zALjr7I0vRRgPRbY43AeWPnQuLKIA8QX0HLG05mL3G5
gPyxy7sl+4cpJaGD0/cbLrEA6mR5Za6natdzP5rfd4S6IkXYL1maPxgGpKBThIObZlIlH9HXf91Z
WYjnrIIuKGYmkuwrKE1p/b9sL9w+Ci26qYkMAu4LbaJprkJs4j6vbAxUrI6f4rbTC3UupY6EUT6u
u7JfC55zkk3up7sZPb2lzqaaigNThDW2hUpIxWsrdanHsAfWaBuljzopBS5P1Uy/sFo10T8SAsiF
oCIB8obq8AMcFB03/msDM6Wz50nMzNzDHV/4y+WM0mF21bSYV1ZodW7ak/sZxdb3CohLB8Wm7Gpv
oFb6mClNI7zxzSt+BLvXaQM1Eqa62eFo1h9zae6OOJ+IemtmJUuW039od0D2YdxPey3v+lM6IV08
L8uq9suqmgYkJCWh1H/GStSG3pP7/szri6R9C5PXcEMUH8Qz+K5skq9QXZTq/onHf75/fj+oYkps
gL6eYZsyCLroFI6u67S1ZlMHbMMaWWhahoerA/R9jd+z7Sbb+YJ6L1jSYNpkwBSPR/XnMZD6GVxr
tniy00fiP6cJoMB/Fj+UCMy8wgZT2AQbL8bFtUYlQHuECj+yOBuZmkvZ5H+Yi2POWM5HIhDT6Wmw
GlGrOkS/mIW61C/xHDhQZBqoQjU46AzwHFKlsneAp+uhN2vGeOi5RWDVwa46hijLUABXWT+y03ck
IL81nJ7i2JL7Knq5yj95JWAqF9ti2e5ml6cG684Fgp1/TOqiq44FtAx8+h7FJwbUfm+cijWCvDIn
NU1PysKbAeYmlc8zkd+viq2GkIPbsMvjrOh47BWt5iGPOp9n2kiE3mC6AK8No5K1P6RObMunDLXA
OAmTqLQedKKfUjfH/8y4uEOTwiFgrEfBrfa0Rtg91hI7lzU8QCWpcwJLfmIG/xK/etWl45Zlv7kK
HcNW3b28jyjmqx/z/sgBVnQHxMs96gLAyZR2STJiQqbiU0c3d3NObTFrr5qqjh/y9nY5KThINUEz
h8EbsIWHLHWpaMAuQcsw3gQTAWlOwHuWPZdqQ6ada3lWzKSbAIHozJBjlqCS4mWtQ4QYay/h5q4A
J0tkvuGJ465ipCowCrFMHGs0Ub9n8okYIGEugRstLd53sGTJJ6Q4wwaN/5O//d9eyQZMGnZsk39N
BpBUFb+hAHx6Cvqj2es071PPlKWQ4ILUKjgRINppmLMqLnj4CBf0/55PxMka6rDs/w/OlvkavNki
ptmXDqN90nlQdUXcFghY05IG6ZXt6R/BcBRZsTIQ253Ryybzdzx4sIqIvdknAwrXujGCNIJjiVcK
XMAF++dIrFz7hl/aQYXV71z7CG6s0sEHQgdaOxfthUA6TZ+COBTqxZBGch84oY/FxSx/m/hO7xbb
lWTnSOYVYISD9XtUtp+0gM5RcfXkPG802rUJOj8aIrxt15UOVrvqjCrgJkxa8BuNsdYExMwYdMua
YruBQlLi2PTm2O7d9ZPBT/1hlGHF5oozhxn72wI2+tJFn9fEzhYin4NFlmsvK27GhZRX+5uumBb0
ElpfymwHbLa5LNr+I4zJ+JqoblBwvwFGp5KUoigucM2X5FgMKHJ+sPtDI8lmEEfsx5xxeYZCgrWX
IrBLdrQE9Cj2YLnsk9HWflMbAlh/V/TrgvOoFUpLKhG+ovNB1u+pKX3hObr031V5S9Gb6UT9R5uT
KVLjy+f2LcK3BTbTLLPAFhizxkg75azkInbVxo3T2RMnk7AcxcLCbo5/q0ofl/ji6TT83p+P1LHb
saX108W516fD6WT0M58sRThkt1MlaDuMoILuMuttB1LNNNK6EZtEsK1KMWEhuZbBWyhIYdWe7HRS
gc5Ct5DZrCDMtOuD/jvKywtNZjIcKyXbFyS7s6AcTCHcFXjNtXDcLYI1CjjnuNUAImGNsrbFZmCx
Z0mYS4e23qSNSwBqVZbOCqwLdHhOCSiF4OOIIF+qPrx/K+VEI2jMcWlSMob0Sx/IjdNXlkfWSsOP
hAfbgI1wKx/EZxvdC/ZLLC1CQU5Qs64/t1EL0IEBFcMMMBdVthGwlBQ7XAeBla30jIytj7cJt2pu
jPKN5OBbIqBKdWNI7s+XjMZaYx4pmBcUiBPctuJAO6LlevvbANFjC0iRdr/7Fa961qWPKcqtP8q5
j7oZk/FMqSccg1DwdwpyCYzZ8s8DhrlGzwQr0SkeJQUbvn8FXGsE+j5HHZdoB5OO0oynTY3COb9L
FJnGKINowPFC39UJHOv6H08GlMqkUeXR3xpQWuTRv21hhsX75Zyxh+TlFaWIJI+aGWunQ8YlKkYe
sKZql4HoeozWs6v4M2ti0iNA3AoBL6e4iBSQETjqVxmSzJ2leKqm1z1sU8PHWl0FqFVamroeax7Q
WdS1o5AkNDtzh5ElA433SXKg2Bxvf0qH8QELk669r2oBLErmwl6BTzEM2I6SAVZ9q/wgxgOvwD+d
/yoEVH0lPZUQzjqy28oXjFOPL/sz+1w1s55E5X6NvkbxvwUhDVP7cU7yn2D22lWt7obzHZFKLcjl
MQpxNvrbxeaT/95mtXVhpSfDoINS8g5FA1LcWxRHzv1rNHEJXYXl24KVp035r6jZZatU9hbYqHaP
UBZ3wzlrS5RT5pXDShm5cJdIWi42i9ZXn5K6KpVrrT/h4wCjXf9BHO+fibQvAXezaK/ykN657brE
Mf+2N4VK/r7tHcztYdAysjDxV3HvQcEjXAkWS4tUX4UABlkFQZO8FaB9RlWsUjVoV57S3XX9BlIl
e2f8C6HhcSgVZVlBg76z4YjXwsKdM2OwGM5ZXTe/ii8Pd19zfztbsEfKF57yjt1dncMN8wKYl06H
AxrwZYuerAOIrbVrw6LaJFiru4gBB6DuiUBRcyzYgrBxn/cOSu+Y6N+H9RWCtzwSfPTYrza6y/wD
cx3xDrDzylGQcMCf6R+ceSTC4njVXXxzzClvowfMFmQfVITIHzLlqSyloScIeP3fqtBNbcuQE8ma
KPt30WQVZYnG7Y9DB/OstizRFgJJlNKK1ID+V7ZsSOpcWCx8H/p/UV5Aa7MQueGaGXUBrtHHYEgC
OpDA/fppYH31mID+RDL3KrxKZYiEh2ZWDIC7b0hUZMrNkYjAXLII8CJxgthTG2wQWuJsIjnvzOf6
BfldYRPGgP6zaKz1YrDgqVMRlF5Utocx2yFQk2Z6xq2HxBXPEZj6KZ7Hy3yuqfEyktMOawqTMWiA
F0VsUH2LGTnwKMlQK7eZqOcTVANeaoJHfg3ZsnayQ9+6NbZUO0HHvpYHhrHHtiBSQQh5INGTddo5
3u7FsGi1gQYZzPuivKDe+WiQzHdnqRjDVh5tIDwvetBwPdn849D1TwKyDEIZX5TeQEfeVVH9X/ym
zD1p1y8qtWnBPaglE/Lrwr60YNFTJ0wQdRMhri6ryBqSe0xyfvuZ2hb6Q1wVeCxeczyuudUeTOcP
iO9Cr/PXchlXGrLw4wUmXK7t80WV8P5fnZ26HmPY7o4iTrvfmaOQ7dGMz/vdvTAagQYZgnDM7qBg
tccy0B7HhN+x8T2Cj1VC/2JP2+EIcDf18KHhBpGAnqTaG8DXnD+yobPPnhyPa2zPtyRxpI49l9Zg
lyprOgGuoj9hmBWGPkWaZD9nmIHJXQfPPdeH0xOPkw44jRSz/+LeiJDPKEfxW66sN3Jp2hQO0UCO
qODUBXvbtIpJzIngPdk9qEfj5zhsnZiuuUnrEs4dNnGuKLRqBTkw5+o8dNgZRzx5d6jPUPIHUtUn
AQnNgTH+UInGf3sZl7dyaVYqh49QO3iuYqA7W3CMqjhm8nHgblkR5S8LnK1SzbzqupknXEFXdMmx
zg0O9gdcZcP50XjlujrpJel/88hJ2jPwglYiZ5TJfdkm2LskjuFryR8+zE+KHR0KQ5QVSsFwiNcL
ysIsKCI04Q9az0s6xDV3X0jyeOTdJRWSPVIHnLluDTx9uelbwfYr41Sp4aRZWbfzFfVe13nyFQ8a
jjTWnAZ6CkIoFuYLWEY92h4QC2mu69aQWWG0jBAPXlQO/nu2LRAYCKA2BxmxreuDl5HZHXYhO6Cq
3OVdOjiPIjKwK0VyQ7DKQKJA/4+59e4uQDEABMTNRR1/PQjbYBon5GOMQ5SKr73LVcwNoEwTRUCn
UofwKy3kuAMHBqQf5balf37wYlWKXmJwZmzKT0eZ+yVp5SfSqYtGWfs1Qs5vx7CBi4zodtcNUHTu
x1lLeBREyckhL/IUEM0krTsoiWoMq9hAEeRSMnQuVYxQTgRnzJOK2W/Cu9MVPRyjmtrtEiovGmTm
jXZuxCQhTfKbUbRvvhs8PfbfO4opYO5wCBXFaNvmj/9MYAsPORHwAtxj934KxCMT6xngdOMeP7ga
ZEqDC6OAWFmYClAXWSk95E5fPaO/tCbEaflwzQpYZkh3qp+fVvnH+QoHRDR2N7/LtCC3G43XudLX
kv/X1Z283/5ySP0rNnZw//t7Cgs7f/P0pX+1wVLOwDhw2qtr5l+zL8pAGan+HAXu+KpMpY2HKSDs
SYVtTmfY746DM84vxlFlOsscDseTQ9ZvSTIKjZIqjX0ZksOE3GSqRp8j9lRctqRs0fFYY/VkHP8Z
HvKBqMfz9Q1dGTdFU/WvIYvchLT0g8NX6lbD71Lz5r4iiPDFZMQm//AiESHD4TarhllQmlnOh9Ca
SXGC21pZXsRa8ev7a8FAAc7TAA9vh8FaTaJEsWdgJXXlfBX3wvJYcErnV2K3kiK/fyB5b+lofx10
3WvqNTtILSJy+eJ2MdAMXJq76Ojv8ZQONG5aUMoP4EWvMUUb71AGF7EtZUEoFfYY30BnSC56iWk8
eZHg0+j9BJW9xGY+l8JJIvJT65aTHV+U5JEMicXVIXpp/Tef5xsMnsN8RELkxZzzUDnDI0ctnHMv
irP/tg4zcIG1D/onOSb1bQWgn6fX8ZUZypRreFY4Ya4FGDul55fbB0xkaafNA+BXTYAe3A9S5nd5
Xz2myRCdnZF2unySc0JWdRfng8le9J0apEmnde1S9Vt+zM0XS2T2goUS1TKvqki04Yle4otV+LDm
jRq7KTnvOzAPENGJObof4CVLdK2NwwC9Ez2fjlMisSRkjtPdA+CJC6zuFRjM02B7qQdSt653fKpp
g/yiStQF/26RYovPMwXfaJdEmqKENybGD1PmYmQWJMKPBOwjL+vQSwmlykd8uGnYNbtwf326FP30
rlyL9f2W0Ci/0QrxYccEwcy3doWO/G6jNRhXiigy+/gt3DA8JFcfPlGYyl+p6UlxISA/wb4xwP6s
yp/3/d5kRZaeIgO1ejTQm6dbN+LhGIYerKDKzCgGL6II8a0eauiINBA+ig2P2AJKta3z9H2b7bbB
/HaXTS/JFwdnbRwX6kBnSN5VA1TpzmxEoGSJd4HNnPpNGQ68TNjzBNnFSAGlGExXQll0Dg8AnxKL
VaRW/0LbHGTWZavMutHr35KUMakoxnKYK47KYLnwieB4tLHSJxw2l6Itikw7hoU8kL2HaqAEdsP5
qRYsng61GYXF16fCK665uaz5y3h1k5zE8gg39SwckrYM99/COSrk8f0dFOfXrko+Qyc3MVqjl445
5pTRd10Y1okI2YgsZAH9PPpt/BVMbXxG1cLLYpSDsulp3fV/gnwgijXE2PAkCT00Rmm0oGz9CMMH
hOLvBDQ9eWClNnBpTL9qBTuJ+mwYkFn25m1CyWFEPYeZ5eL+8tsFaxXt6JdtMQ+48GrDaBQxx8iI
8Un5v172c4WWBLTCvIfo+l3kWEEireR5UmdApmuQzKvDJKEH+P2wH9dwTOgldbEbrwI7gt1G/S18
z1OKvBqWz8kioAMwqKtxIGT6WqX7WOpyE42AoUYW1KVTclvis9FqA9Vo97t7nykxWDyTJI6O2ohI
TYSweGg453pwIBU0OSQ8pK6LvhP24CHf1EdB4IYKCgq7NZC1ZyQe0xmSmQEQGfbgimQIMlMDGZ3g
Qt8tbyRFo0CK6Lq57Rv11122Tcy3a6cmMS2vqS82hx9EIxMm3rKPEkOYWRUkwgjObeS/UzTt9djr
dZOOe6C2IPUhvHJCTZyKqWZapLLzDDRP/zq/DkJpAsCD/SaFHvZDuAP8P5qofRw6chZBQsY1mIYA
J2CGvLKdHnU+mZAQ9GV62sqf+waC6T7Z+0+KHohiXdqRYepn5/+a9IJW+feNqSZ3nTnigBNnCE2W
F0Nt/gWQ7riPdIDx8v38hX7QAjCLBqVMocDcHXuhkW/c1/iJmQHn4fnGtmVEXx1Ptb6eEyOE6GmO
gJ6zuyVIrfYhQgK1vMFNlf10vC6RqfKHBsUKKUjc1664OahM8S07OPk42ur4vOwPLorSK3H7k408
SOYiZuQYSJFqSKZhtc1rxoSIfBItIKpqw++jFm6ha8Tp5ZCFUFVQSZhyQffIylIWuiOlr7binqLa
mwR5yFETX9dvnG4o+Gh5de02V2XFfUN1ur0Im8i3KdAzz5UV7YjjtugK4aKkYGTPGZ199j889cuw
1WxhSRId34hNucHD0lt31p0nNX8ZgeFF3aUDX5yccLk+SguzPkJ+s/KgytZ0AFmLtVQwWLc3ABx/
b7a2fVkkveKqaHi7L2jmN5vnAAZhGJPlQRGd6VYVPsRrDi5FAWJMEORnwYfSbLG9Q7u2uev4H5vX
Vdjgo2TeWlDaQT8IowS4LwoW7vmWca2ZVwo7p/8x3E53cK40J/1cXHnkiHptJUXax9ouCPlGA2nN
OCgXmwtC5iGILU6K85MTBL02sjDFKjbcosBG9JLpvqdzUmqriMSgS71h+sswzz5+QCY7pghmbH+q
/mWF3dGTc1tGuPYhA/XSDu0C3OsvyH0huf2rib3R4+CU6pm1qyoZgIY7LVIv4qsLjY96URVwBFGU
zEQEBJKVmLIb4WfgiKJ2ogX9YKNMBwja34b1FdZO++RnP0krepDjM/pQ/fOqPX5TVsz0hknJyxQF
9FlmB2X7k4QIkhEHCGhGgRTJRLukA2koK09GjafrbMMM6d6TWSpcOMSlcEV/uq5huupPz00cuzR/
E/6GmweqOeiZ18dikWhRo/pvBi1TvmEvdDYeI6pk3jh33OVSoS+Csh6hwuQhNcE+u9B1HbxUE6hE
1Tyk8PRqvsD6tjpMBbTRexKd0HhNmHYS+QoU14puns6xmlanhmPoAr6XeydVw5jgSs1bWYaQa4hZ
Ku57JALZpILsN6OYjVMT3k0QAmXyaDzyBebyGMGoNJNL0NcqV4tAnUw8UgouKqLgy62nymMiKMDu
2D00QqaU95KOPSKPYr1ZM5GuaHwlkvTLmKlyJDPCVBbYjhlwEtr5XSWUvVXbRVD0tnFHOVc4QJ+5
37/0hz5oej2Js0oi1ae3PWp+/5fC0oETZNHRh9kNmNoxLXR1Im669gvGq3QiLnc8mmDXO3+8yZyq
izN+D1OrGWCIp0M69bfIMnY4mmQVNd+yMA45/8vdEaRBcAtm97/bikitFfKvb4Fb+iXJPKfemMPu
aGvCPwsm5UBLxB+h4Xz8o/oldiYEuKEcfG/RNtrvmF3TbTC044JVVDAhA6zUfgGHgfPvMuyvSv+X
2HJqFCA+OwWfqDPobZPij2pQDODGk/YHQlVKXVONCz0+fehG9NkzoudqIDDdpVFO4Q7GkUvV84Rm
Xomo/jcbOzHcL9fnezjf2yUcInPI9fUGcQU+R6tVZY3TsfBr0qp0QJStwqQVpxJCbfViacRCPvvF
u6y161xCQfmah5I7CpVJDrhI89aosVROgHE4/6H1pZmKO+KqBzNroyU9M8Y85X7g9IeDbO303wzH
u2F1jkV0eN282xCUK0HuQZa7MvzQfDfJIFujjWBfSfaB98y3V+cjfSWZNdVrw24xMo0pt5P92JSV
733fTcuh/wwljDYwsxlWcosS0vHC7Kjhv7t753tkW/R79E9tLLgUAFHeJ5HFc9ewvCWp7vdr528C
z3eA5PV6Rfi3vVaj6Jl8mpPM0yZWzcOU23f5+cEuprUqb0AoYGJL7OrcK1ODMU8pCP1Tp1zXpbjs
Ah5qdxHGAQZOM919h1oz3rPgwmZVeoTCE2sTpB67EBf4lsCMBMZUhpVfu/ncIGvNLdoGjH+jrJlh
hF/fc8f/VP3+gmjrD7b8bZi1fNapUYK6r9YN2Vap2dbAVWm4ytL65CgyjaUISbhk4HT082mLCqMl
/3NPdQ+NJ0dRyydRrjpInlWAtPszLGxbpMo62UX9oX5nnMsC2e4Y3bN9VvWv34EfTOK03eyodE9o
K8u0Cm0d4RazsGXvTrNzs340fH+esK57NmDr7wii94xCZJJHVVW/LvjFpxArpwv3BJhh2PRJf1VJ
bJILV0Jbmn6aVbsmxpzwXLlx7y/Q2sSEatLMos31iy0Ol9ZxeIGk3aHbgjprK2Va8Gs5TaSmnWmQ
D1qeNui5toCpZjjpzH19TrxkirpwqRMTy9J2G4zXoTS8QjXSTmHwqhQxrhVHPnxOji94EznRsEPB
gTiAfMx8ey7tn/LXUE4/dWr8OrFRnSZXpG+mpT+zQOIGt61UpRiJBedQoOY/GV67k0zR1wSZMU78
B0vSQekG3qSrWv8GxknD1QDD8nyUSS5zakM0UsZIrhwbhnrzYlQmh45lfiWNOMGfLLeTaWEB1HYi
AAOW/I/r3IyAx+zY1dj9c12bnHRPgU2JfqQ2q99ozDB2zo9UHY+z0eidQV9i9OQ27eiZz/Cc74td
rHMZZWkuR1hVRmZ8BOo20RyUwgNuBCSAn4HvpEjGw7JOPzDy3wQow5iKo3FlnI9AVBR7VBIaWBGW
tpualpGDAKOaaBI2edBlEItwtM1BOnfTl6JpmDUJOOOHsGpGLOtvzmCSiroljhjkR9yhKf/SEhQD
+P2Tthz4zYFO98nYvRGa5z3X8SaEr13RgirXYcpSxJd3VU2Gkd+O4djjkEHf4wZlsHerw073BKQe
tX49WoHfGYPnTCrZTd31dwdlVIk8e8w6jmlHbxifY48Zo89v9Re8NYnJLkzrkmp6hGZPHj0s40H+
F2NeIza627oOis0YyT3fTRK2NGJVjsn8ORRkrBGJxEZ56eVJXEdKZM1FiDooqUoqI4C72abIo6gR
g5GC63gDnVz2HiRu/F+eh8YeAU2nlsGd1RDkXKkTyH8EVjw14hiX5lxGfrBiKqcMPwTmoLXBetIn
ubNUt1HjwWWcxq5jkQJucEPsf5k9udiku6tLeASTCECcLFLxe/1a0EAW7BCjokvnZw2/Ih1DXo7l
oMF6c2cWTcol95yoVqEncD4lGfYqGD9SMEhE1AqKiQ50TfU5jyWPCmt5/i07eEIiAdxMPtC0M+oV
dvqXVxCBwSxaduM9S0MQoNC+liscrI9jERbClr0xozM68nFd5UU/CGoeJd04V2g+Mt7+0Jq3zq6B
e5M1xbuTvu9kSGlvoq5lkyIqkuS8ZrgfiFWjHw70KNYIT5lXX56k51XgmGjkF/RKT1g7jt7aZGmG
3nYCn9PUW6vo1YVQXLpOIeAXQD8LKFQU7MZIEyf7DR4qzxMAC0f/PwtWdPv8uBh7fg5/mL9ZSCkW
ja249eDxxfo+KMZ8vtGuA8U6lFRe+4E9Xqj9fg6dRCV5fYPKY+R58QO2HSdYNJQgCwsmvqkp2ZOQ
EBRhj81AackHX5NI+cWj7VoHs4pmCcGZrTMBR8it8JCgiB7rMnT3jhlO7NOJIgAGPc8+vAoiKXp4
TUg69HSMU+BTbA8HUsh3OuSoiTrQ4EiFrFNUq7PCHIRRskgMrC5KEfJmi8sL+gLjdlBWucUaAzUB
JJP0dcC7EZKzZcc2yCr//DdqGl/JKdvnJ0FvQMDIGstCqDHmAlECw/k2htkZ3dpTjYnMAzgLfTTO
GoHk7E9E6m5SfES+Z4cGomX8jaMrK73dRHUYuA3q6wRSF3KHG6sxYuoRE9ZYwSadjhWUhQvNJoPh
xwhxgzYEhGIO0QKoX3n+VL6vb7xwm9T127Jub+1eq7av25FqAMiQpWae/R/IOp1oy73Jchl6Y+Dl
EwRemWIN7yEGP9lpq/x51SIFiBoqEGgq66Ww3kWKxJluWu5nkEJELnMdPxZUMm1R/znUjNP4IMYd
lI9f+aejqxSh6xVGaqipXYzBTNaI8RiJQRdUnneG8Pl12W1TIRnvGuXePosx8+BfWpjTtVHpOSEg
sRW+tL/L3ioaYbS50H8E6iMGLZXvPXiQyMQHDR9tTdTARUHvaDtfVKlDpGjvWUVmJEaQWAAf7enW
y0IU0Y6C1Qj/EDz+W0t5Fy7eFoyUoq+uzLLMmZP2L1vDDDapbYBQosbQnVxHOt9UbcanXECYALWm
oocx7/3SmFZUfAMUlsl3RaVpFJou3FcnhHYdDDhY+t5AmpKKXMpMMYkFu+q4atr3ZUhE4nzBnWf2
aMVAi+v/u+D8tIK/cXQNeVoMnB4M517Iwjus8GJSwR5JUUqUuQo/iqdw9wTbRR3ZYvucvK6/C6Qz
Wz0Tc+NouJlWYbo9QQT7y4e/hhZRb/w7qRf30gwYq3xxTunR6smNOKkVESAhqiFq4uh3woIQJgoU
8Pn5U3QdJpPgjT7wISndyomh/P69Pmy93KyDJhXEedKTxI6uG/WtC8kMBReD0j/2fMmaa2cllY6Y
ZTfZrmL/9uZX7WnDCPj2h/CAKssqm/1oLVYM2QPEkXwvj5HqD5ZyW67Y2VT9iAJ4cpMOHoTj/YfW
4I3nPDk8EuUg2YGIRaoEmEw/oE1uqI7CS2p+t7wCz4bcLjxW64ZEXxC61KNnQ0UuIXaZj2qLG0T1
YXkJWojfPmdHV5D86l55C2bJY9y97Ha0iakWxndFK2JuEily4UttOvvnLT+J8GexNGt4ZE0Vr+W2
2RrWjSfJEE7vKA7OGo0SA90z3Kw/dMP9jgOg+CJQF0CN43AxfrpH1ML6mAkguu1Rr2A4bpzowWgc
R/JbEP4ndhZDY35McOibQ4Qw6dZEyBTUfeU2I9WfiQdKQpsh0QNp3Nk1JhnegDo5JHxFtEN8lER1
8ZkAHE2EkOISihm8ma1CucOU9J5LClrE46eKkuHKycn98VXHzs2Y5Ehf20piJlk8yVK2qlzUArxb
NoUz+w+w7YFyyMh3B7yVDQVSCWWhFZUOTsCdoqjCB2IqNg3QetXvW0joKeOfSsV3PFg6JOAhcegl
sgO0NOLeVEClNJO84hDAPJJZwujrOSURzFAoSuTpp043TOFWAzqx1SLiFELb2iHU1H9cbxnu59pK
0AEP8C2/Bd78HeQJElUtssujn82wQoonYHkV0mWsCGrCACe+55NlKArdpcZH2QVItN910/3Fxn+3
uHTsVqVpUzwJNCm6BzG9QttKc6PIFApxWbYYY41Kex74V/5q+AYEjOdjbtWRA2deHYRmyXMmyEe0
ldN4C8e24jrqOGJqWhxk3qXqyaDfHXW5lM9pRmlJgJ1beUyFLzII+7mCiWuIJEiNkxuW1k1K5lk/
JJ3h4yvlLWUPzlSO5LnaZtXS/t+cuwaknVn1ynGOd0ggqjWcmLOpQYh3lEjYzLUlaPUFaD5BljqY
67WVUs7/Q6bef+jO9K+4u5LFSupD/g/ify8WF/A7sJcr7vk0MlX3KEkS0SJk7FB2dmlFbRFcNDwf
U3iSOU4AmV0O6YQK+iNn86ctzwW4goKtm+8ezS8d86PLxifMS7liMvgwb3AYNdBdXwiX5JWkuOJf
+IAwPKiWTDEYYYSGPoYj1kr2kWH1KtXJ/mZrWtt9yxoUrxAb6kuZXwWiZOkuz6/vUHLSGUx7J8lJ
Trh9zMGSKA/0Rek1TjPWhf5M7fFSePCTk9RyqNwhLUOEx0yWP6bL7x42jzamzuzSUdrOTtKtYs2B
itnk6HLTtsVtZgIGSo7XbT9dY73IYNYmPckHcfJloEI7i3rZIRyHt/r/HSVn5f23bTk0JHT+4trT
YoFCe89Ik+Pc05oPlH+Xgzfnqn99IZ33JQ5+xrRtu8dqJKOfIpYnpheNDc4/UIMY5JjUQ39fWmb4
0ESb91Vnsr37IQdI4uYJ5FwkcV/61Ctfk7+n+ZRIooKRHB167BAcVw/bfKizDqdL8xsqBd4BWSp3
hL7Uh4fL0/NB2bixNq4brNQcnNWSk89nTfnC0EZ2ZQCB4Sk9TynhhcCy3HTWO8NYonZVSpTS35ZM
sQY0UnD6frbqTBu1iMvZYRGFpN2Z1i80KP462YL0rrULpkBvBNRH9uhJwOKAjNLcmocgnhk7aFlo
e2CEKYuBuEg1GldU503T5Ao2z/srX1YNrT7WtiBHUzWkt8m1M7NZ4qAgZnwM3sS5g/PnePvI4kPd
Aqri+2iB2U91CI9U1IoRq19ihGDnOdyOwkeyKAQTKI9lYOLbrG/VQfzeGFiMsWtPUlhaVnaWALBj
2AU0DRBs4ZiE+M8W3GtYh9QE6abZHsum8XN0rE9kGhuqR6QdIbdYrOMmipQcSH+f9Lm6IbbG/K6g
S3JGUk2JigQqfGH+hAP8IRlvvfTJszFU5nGfuUpf/hjnzwdxx4oBGAhHQK75r1fBZWPudejaXPPH
/7zhgy9XwKynyb3TUDdeiciMBzOwg+25SBpGks9JYNpmLsTApVhT2xVcK2vTeF/P+Mv+AWWLoqB2
13GMBNUZfAiil22Cxm57kPF3XO7DSnkr0UcHzn0dUhimbg8R6Q9omuqKWzSK5wN8zdFOR3fteFt9
+oQCt66AaSFpzdJ+vpUo8q6wmxKSRkkFw745SbepQDfU1DXYFzgqAs6dmcI/QFReRKMSBCps27X+
xvly452M+/Ygn8ABHCB33xp5rg2LgyJZE5MBncbc5CMJSTUMYHCNM93pSret65AW49Qu8v6R+NGR
rbqRo03wmjRhHAVFdCCXT1VY16/YCofq/T3eM091MzXb4Jx2WSGy+DWrv3Qeyl0Vztma2v1DFc90
8FUVFARK41a0yTQv4CXx6SrG1x9tPwumFrSOid8txm5chEo+P7VcBaWSU0BKYr33qFxhAtWhhCFO
ZAOhmX+Z/SKx4QlCTu/yfb1l/G2zFOA4DsK4fDgr6bSX1OXVnmxBNFWJHUZJhVpSMQtcWLNJBODv
5g8LuDjNapHK8IJCqQLmXGTe9fasLL73obfVezC9NFld0VGiwk//dN/aDneYnXCCT0QUh7T5M7Y6
5+f+Vwi6hD7ZD4l5ivS0qNMIMh0KLuDtsWGJsDLWarJXT9f6rElaprg3xX7tx7Lhg1B52+tz50BX
VUi3mjthcjM9n+QvubuJ/A5CnWLQRH0Z+Yj8/zZEhVTQecz+eK2U2m4VmlZQMTR/o3NBVxprDAl0
cwax2kV0hyRk7vT9Z0Xfn6VCY9Ql2J0llGb4qUVg0BN1dWqCTp2snA5M5FLps5IC+PJsOby3EInB
XvmSE283fYUAWHO8b4CbeQC6D9HB7YEZvLfuaTj2N4lJ0jgm0BY6DbD5SXcM8/NMft+Uc0Ni/pKg
CwEDYvQ11MTyAbTyWBIld3b2xNz5O9Ax4/RhQE9cPtWxagTL3cA2OsyHC3XZ6Pnjx6ioQRXWDgZG
oLBEP+Tlr8SrVITFd40EllxT07LydD4rmLj783WyPD8HaaZvvUAhaKbO6LWalandZUl17Zdhtgd4
Wp2lirnYrAa79GF30g+IqgAi7Uol57UvmfT/uIDG6NlBrpxqP3sigJBW+pmrNe+FutJX20bcTc69
78BgnvlGEQzyCz38Z6+UaB5b5scoOD1oGuM1t4nfH6nzMHhexse3UQzklHhL3MiAPgc9siRhbOYv
F1B8mISAVxoO9vWBCXzG1fsNOk2AwA4kbikibhhxONZVXYUjPePXk96LX28mjFUK4iWxepiS6LGv
64kUGdIYqgrctuxDRYC1S7YE9USuh0mw6SV70yqXyUdMNaMiTXy/ok0SEpiKk7PZXA5ERirdvTIB
p8furv1p8RjFX3N6ldYgTp+qkFwUjdm0NGKizodWgTmulrVyUwqrFnjTzqyDXbP8MJCmA8j64R4g
YRsq18I14eElqx2yGjnv1XmKsucUTkkrnXY+Pk4bDMyHEY+3szxfZrIiUQ5kVPlMKJUxwvXQ82H3
iAQNe6mWtTG086Q2hwnHQJd9GMJNfJwa+jtWTRBxoj1nJma6EO7Kz48GoqKDyu+mvBSqAYlmpavS
r0ishCucgeQP2F+MuiU/HrmydY3hOKSNgiJo2y3PXqk4dXNsR2cpfVwnzE821D/WoLSuCHBAZURQ
716Z12s+1BJJSjjwO87tFwMD6dxIaIajBgnrzzSpqtWanlChkaIXocZznHVq9tkyHjc75B362qSu
I0cSuS/Wt6UuvwsTndR6+xoExrmrzbLknwpBEGkDM4ox1AjUpgoa0z7gkyXT+NMEYsQd7ay8S4c2
ZkE6evb7gO6+Mdejos+1W+9sELUx8A47pw8ZTj9Jn8J0Iw4NKX6NNdp/yoATdm6/Sn/oaaz+yiIQ
tT5fW2HbhXkSvYFYSQwFuCiJIs5no5UV8TBC8gpdUPZGPaw6fhsnc+svj5EoRR634hxNKbyCW4Hh
paQ6m90p6dRsuAdNQlozKsElTZsiJUE+/WqUvd4KSg0ZMLJMgsqOUYwo/iKOZ/I3P5BHPVweeedV
zdGdg9zy9C7d26ugPm0PnafkWUN4Nm9VQHwanQCAl+ZKYEuozxcLpzaDLZ8jh84IUG2CIdEKYP7c
hdkf9ZZN1iBUhb8gIYoS8D/ttktUSvvyYvEDa9OC2rQAAwaB9vctU9Btl229xHs3nL3IXNWGlI/3
EMtRYvebuM+R4pLaxpd6Q2Ju0se/ZWfkgSwmb2nRwZz54RTBJyCoMM1WOXzXKtwfURGfgYaIW/jD
+GW8ojIyYEXrnbxB+ckOxDZirOuMqLmuFOSBVFJNOLYfN6cS6JS7rIg4HBnsdKICma/jRc3e+Ow7
UTE4+j/8wy157pw4vgUWfObVxX45qN2U0dqYxIAcfKnvXtIhS2s+XRkB1IMCyWCQJK8tn5jM9fS/
QOGnJ+RX9dr5yaKJrPbsp/7agwm0+gMRF2vv/Pkxj0ZP4rAKDA/SCYaVl/fZWjc+d7/H2SDs9Dwl
lQady/eB4qlshfCW+mb9viJ5VsMwDHYK1lsbesknypxMavw6/eC32NInfm0WGUHNYmDZz+Y2sFfH
tezvbNszkzKgUYAAJwyV+MniieukJqkRdzxqwOdxCnf1jo0RWz/sH/Lj8NzhsMgkg4kGRrmBsEKQ
YE2YVbicGUh2Cdst4+JxYLCmfmcF31dj4kdlmyBu1kbRWPr5UbjQDZmphn6AjYrWazwTrM+eCbXl
agHWEmOpZOaQtvi105Liva/1QJE0V5dugNdPQ4Y7eHixU1U1AyH1pnMRdH2rmc+Ey7ySFGmUpiuJ
n/ldCQlV8eGIw690ipSFGzko8tlM9q6wwC8jn8aC1cWlhvRAOP5eNe0S5Ot0LPywFoM081zaHthf
SaQ6ICUMckaWHpoHu6Mubo1Pak7K6tDWEjlg5GAbWNBrHjAHPzn4dfVSwHhtS+ie3Y+33dvIlfbz
pQFppzYQt++ntTWmyJ3RyadkOppWw2n1gAYTcLjr7hUXLLtLkxAzGJCH2Urf7dQ/hlHeY7Pm3/5M
Q5lV0BlRWwTvaPIb4ZFviBTyNYlRGK/pjphAVvphIV68TWL5Qv+0aFH8hops4XFRoq+U8ak4cHdw
pdeuoQQts9+MmhsjvkqMhEnjHnTS48LAwMG2XHDPpbZZcIGtZFvE5NWrIzy2lxEbVof7TDKNNXMW
gkRaLbu1qG0j5oe4E0O7DydYn/vY3J19hSzwPmtw8X0hNN8v8nARHwMZGLzPlQ4nd6kz3dCDpag7
cfhJ3jYwJWltkWj2pNlP1dYN08MNwWPIaJUIihNz9LRJUL7c6OKnL0MA2nS9LAyVQ30T3Y8cPASj
kyRJILgUlTiEWURXDs5bBQtGH3gSSnb8RvTST/O6QsXRnrp9jJCcwde+08uNMDechqE07B+Zbjny
TgRFdFe5TvL/yLj2FSgiaJ6vbWrOi3ReR/Q//nS12CvNC0exwwiUXAUMTZwdJqE8mHRT19S31A2v
FcO/TtPL+6xDAResR/HvI8zYjT072AsVaoIOirNblPyCYPMlQcKMTRQDL5K60tbbpd5Ma/HFySsf
IBQE/tpVksdqYNXsEif6FOkE6YiUpc+KwhydcnqnGmqhjw34KouUg3TQp5HMS6cPGnOmSRLLdqPm
m/MFyVZqXNgMqTlRXBmqLJs+KlHpHtbCm/56iT+/KzOJqbFDZZx9pW4la86wb23mvGFn7al/Ncow
w/SoSSt1+qAdOEUREbv73FvzUu9gj2XWyBQv4jrVKc1xPfiri34oZZkGbs5clMRt5MHasmEY2ImT
UUKnMYlMlzs2qjfXkD/y9AiUAeIUqWqLmc94DEFFaE2+521HK43FnfAIBGWsePDRuvfYJSdSFoxN
1Pba8OTya58kCquohUCeaAQkqD4h9u//m0++V9WY1f64NpThTZmx0xB4LWOWDEwln7XIzYob1lQe
ofVqCpaR2D6rEID3Sv6L4fpzPB9+q2ubX4mFnQCLasIQxQwGutUHfrCRbneN7e4/+WsSNHM4fD2I
QTd6i4bRbBEnLYhDnPDzzXssNXmYduxl6xCzpWwkdMbeHSksS7vsnlTfGxE+VPhqSicTAU/f479m
vvn1JAo4Vo7qvnlgs7T/+ZzM7g1e1hVsoLM0Hn7U3bff7pvy/UDYwztxFj8l9H40wtrDntKKt2js
3a4dOGkXDFwD/UDAI3maPA/evCxnq0Eget20DPo8OibXauzyaebTjD0oUAEDWM29qRFJyjtoQCHb
Do5YRV000ylzQG+I9GDRJRok6lDuqDwcwFsL2+NBr/OLDjCX6kGU7CsXGhs/4w9XhAgQ6YQBvkE8
PXcIRxRbEy5u6KZoy0NJQXaWMQ4f3Ret+zgj/cC2riflIEJDWobK0jVWysb3QHcu5OxH1fW02hrE
0XH4/kXa1iEt0npiQ5zT9XzrprDVBQPt1tk3OHx7tmvgRVhU/2V2RChAltjdzoPWujuZmH5QAxcC
43AV6VrmUKH7zy8WTO2L+tW3DXSAbrGy9BQf3ZNa8NVDThLfn2XQLmeHCeYA0srY/zRLiECrCKJw
N3irFUSb8fQk/Cn/hVSKoVAWwZuBfKnHs+T66Fl903bLF6ceHkiZR4CQHUsEw4AmUacMLEfsMCOL
rliYoOsbffljJzz8Sp9msPRSMU+PMUHRvq/r44sibOWho4Dutkb7IbkwbhhCwJgsJWWJU/tLI/nl
BbCTSsWpyJxOVoDH/myRGX5LFQofpCFESIoHuGUJSP83/6wEcxw91wY2lNovPaWUNgE9g5xzk2WA
7io7rVLlq0vIbbp7qS6MWo7TqnIHYU0lfJY0tjKUOaJviBOM1lc0CpkZQSv/cpHx+bERIrViChaL
Wds6vtLJjh4LQ6npk+hrMyzIzgKnES3KR9Y4aaLo/ejTWxmuwimivL5nJtbkXciOFcp6i0HU5Dvl
W9XSPcUkjwaWnDLz+a1SO4LeZAq7S1AhZgw+Uw8+0K9MPPymp6B4EIh7q7CL3UIiMJSFZ2JJI2Oo
GgiMXBgZlt3Mf/wWoXhGzLuBFNBV9t7P7Be8netEivhmaiFmC3UqAR6rueEq7Ipr6G+Jk4t8CeTB
5UekHpCacburprtbPse5MhegwUZ20ITBEwvtzvlBUE5fFePE7qENZB+8bBSNCtZD65ej8/0xWLfU
xoH49bwGV+aQBANAodW5o7dEEi7ZUcWYxHIl531og6v1/EWZpuyNr9tsCiorBYvKpL5y337WtUFk
JpTmbBbF9ohbceGeZNe5lx4TeU6HogV3QWkWVhqxvyyA6j9bxMcDjtw8h5pw5hLG4wFeQ/bZZzqk
3DgO1VbmWrJGyoOIrjAs+QbBgiUUOzLI8YOV0WrNfh5dAhcOM8otVqXnrO5/+vtyzEI4vkXPccqa
RdPuYTlvqiyPZg2p/NhsFuKokWIqMZ/T56XhA/AiLv3Zad3KEbXJ0ofzfbv8JyANbCfOhBRpk5YJ
vLDnuivH/2HcBXKRp/i2ytWcx5+0I9lf7gVeznn3VvYX+iHhP9vMsbMaDnjDGON6+fzFy4h7wAo+
QssBJjywFvcV29xBlLT6KcJEiXd+drFEOSsc0VuSUjPpU+rr+dw5ryHRDm6RZqDzxPpqHzfC4Iox
sSp9Kzh9C2TNXMp7m5nVNrKZRnL6CNm+260L+Kxb9s4wD/ogYILu91GC9Fyt9kmnPeAmoLBoyeUO
UG0D2nx6DUvWCgevEVzsiI/4i9up7o4F3Lvn99Q5QvQDmf5dWZRo3kKFS4bD+5BrbEYDVhzHGFfc
Jr+Nx3RAZ5XSn33eD+vDWJ02f+7eYsyrflRvydjvTXPFlJfym2WxtmLGY3UOyrbkP+OoehGB104W
4Ngs+uD55jT893atyULlPWTCDo2Kq+DtLEzW12XUalWYbSHY6TNRR7AeKu0lGP+JPEKhpuAubYpK
igKTtvq5kyHFojdpzINVGGwKd7z6lhEnEKXLpVscLZsFmWpAqaHJxMz/8b2lPOqU/zup03D+VetM
TaZfl8nBgsBsXmsNoeGuDA17PmosLCpih9UeiRWUFn4kf/ICDbN368gkLWkbER/bl6CrnpdG6XjY
P2o3pwltU8oAArltNwx0ifCdFClQOO03O4qxrxpEzNNG0uBVJzudlKKDDZzzzb2Tur7+3QC6g40D
XfjCQYcvex/S3XN0nFe1J4qmrt7fEhYy3f3Q3KP7WXiW5+uG+9TONN8HhxHVhsFwkWIJkhFQmJ8U
5XZYoEYfviLPw+KzEZg8qJ3wuPCgN9FrR0Ux0Y68ysh55IJkujpK7LdVtYOQQwNJ0uMCF9yww5Ft
fA0ZS35EDuyNEGpsxlRz8iSBqmjZcDAgJeHUJiAn0z+iLxF75FiNodnoQPf7+bhwa1lg5OqD+3Z8
RWvWCRiPue+r626/kNb9y4pRna1zDlw27SZbGPqqXidEjCLsPycdHleYFeOpNOj3ulPLFz6abj0i
bQHT2cbTNs9YZ38EcZP5o957T01s1Gb21Xi6NbUP1cjbpVVkz2RO6NrqI23yJhfzvqKX7MkZ3lH8
bw24JZsE1B1xFSdMTi8C5qcbGnGDoZM6CYgrHVFEIRaIMh/AHSacIqveL21i05cABm9AlyW4sXvq
0e0V8vUFLQi8t30lEt1fiYteOp693g5rHmdWp2ozl8Oebyqvl2sANTTc9FJEqeaRgbOrQp3ag8bG
JzRb4r/1+fxRgnpM/j56An1peVKA95e21wA6HIxH102HCl4B0K8IPLQcjtXw83sVlRujY3TcV2Hy
OkWyGVzw5YSbAzKvcYdSn6g4i0FwnO7JTrF+8B+SxyIL/RXxnToYljppT8AuYRzgCaImSXhcxcd0
w36DOP7v152miekASvt7yA3ESHltRTSa8SZ5/R0Ebn8RbOju7hfTht9tTl8YzMAMhDjVeru3F58/
GK5qvwehbkdT/fnLAwbiXik8E3up0RIrAj0sgymqghLZrf2/M+PSoNv2lxVtgee/lROXl/HU52vD
b2DGXmfne+AajJUjctO5xHcBcT+WZFZg1uejnnjrVzlIjaJFVjphTQH+CwKldaT6i0JyG7QXkqpG
dRqdYbDvjlu8gMZxHFIq3/VPDNqi/sUwclSm2j+/VUhsBT8FVQ3CDPepQ/iJp2Dstgf5Yw3K5K11
D4N9HqPsu9UKDxGWPPy/eteP5CYMgv+r5FqO5mbYGEnrbBiamgNXgd5g04+si8Wc1wJrXogKuHDl
sU1hZCzXgOkiIJ/bR0Q6ySVY7N+zyXRBveixPfZC8eZaX+tF1N7PepDewXZQ7uxHOD0Qh2Q8MsxW
KlJEMtmO9EEiUl4745kiuEmVAJ2vjMrysPO/LWLXNdHLoJYXbSEu5HRL/uaiIVIB4O1WWAkldjlT
mjONiQgsRSsjA/Itf2Uwf/VZDhA6pB7RJdUVqfL64V79A/QCbnGm8inJULx9KiB/vEvUM5MuZcgj
GtoGhHe2JaFx628ie3rhQ+X5EUZPycscBPYRliW+TCeu9zmapyAy7WquUndDMHIUA+warFfHgHTC
4L6COj6fVb2U+Ul5IUJf1cyLTfcv6/Ue8JlrXkr9ti34FohCR8rw52i022E7H5C3aYG3h0GNxbml
qOo7yAhiW+WLN2IkB6zCd6+Feqbs7IgVL4X3QBBzEpn6WZxFLL0lVVgNerDZuf1MLWuaPL6I1CaF
nMhntJKTEfh0yGNXwVDiz75osNr7/HNC7Q19P8WuZQ7Ow68mSPyA1nc4Rzh9LRQmt9du74hRt7AE
GLF6r3wTPXMnqCpZfxNUCn97GGciMfLtglc1OpvQp0PZrdvsemf5As8wwbhLFEgkb8SnKcbEXuns
wKIfk07GaFibDtza366FIlU+OqoqhNPt2EqIBsSBXsq34uKgZSJObgDV8+kCzxCOCqfaowwdClXj
qoyZ0V7dO6PCOy+iK3b9BDEoPiCh7SiwXq6bF5/CyxAPCSHg3u6ulOOB2LMoBtFhxP+zE3jNb3Dc
OMEnwc1L4XsfYWXZDL0WkJcc9t8JNHQi4RcVcHoBTrr2vG0cHlypioR4P9ebJaHOznCsZyi3949k
4XXUalQzsbct1U6ugwS5Ls4ZY23CGktuOARIqNOiLhlPcJyRCURKVbfcC2Gt4392hBm7l5ckuwHD
38AorUYVFhwKOLIKOaTEdbXeSwT1DoLmwh5Dh3XHdgBcn+ppIbv9zPPWDYjN00Izsbt8z/ji2hks
a0Va8V+b6dycY7KJRsgD95erS2UnPw+BCHU0FupFCuLCnZXViTu76LHFuZh+LN0CamfjKg8H1E0V
50aUV7VZXueeGiNtUjrvoohIhBZRtiQzlNuyw7tkKFjS/ooqWNk7sT1PQkYjMe5bNJ+KhfISUaND
cosMg567Ia1i4TtnIJ2y8qUi2nfp0oYdeiNNp8YMGJeKwvwpQ4s2Qprp4ijnKMm3uKkWIXxcEtN+
8MB+g9wGAh7iN8b6XST5j00UQA5yLtiZRU4+qLcgP7V4rem6UVCmPwUlE2Kycs67qW7ZPPobov+M
sV1FtFzZpoC2pn308AFrc6mVX7bN+0gL0ejYIECfP/EO7mGhFV9647sSXOQHChFmtUd64eTOaRGT
NLMa0nBsvUB02JaIq86L2172+MJ5pfrPZkaD3c5TuEjrdUTEr+ttNYJ7P6m7d2a1KbW8LWX9hiXo
/MzfKa2CcCFaHeJE+zi2aAm0+sBZq+cp/6S4npO7jSv+TjuDu1nVCAyKdACY/vjsOATtNNpdCxa7
qgRnMp3quxGdoQEqVkLoGO8sVcw5pDIGH1e/i2e6fQoi2fR4205irbe9jphDKQUmxYmS4Md8xhpq
mwDEI1CbrLnO9DN8OUDGhb3s5DwOiUC5UBe5Hp6UoTJrHTDVh57ZyVTQn/3qLbI3PjUBgIS+zC1L
9/o4fT7ROajcyVbdJOa/CAPHI5mbrEAOgR9OswICJczYdK4t2tYglAihtPbTjMCK77uPsYg9H4AZ
/XUENukTRdaV0WyVZMHvCfO8xV0cyqQwnQppL/F7NxXaz9kgjtl6JoN/eh/Wo55jRKaCKldVbfb/
rMPtohCILSn1dViQfDITNnPH9qWhyj/0sA2Rn7q8bWNcFweTpTWmKyM7k1n44Uwpphtp2XjZ5kI+
h4xBXG7yaaB6IInr/Y7eSLZQuRSr7vIl7bSj2gI4ayCJma9FYrluQghQyksjF2MDMVy2Q5foq4Tm
yMFDP+65WEyikKj2SOc0ZXbOd/kktkTBOLzJTqUhnUXLyjLnBwo55N4lHSbYkO0n9siS+m5Ld2dR
hpLjxqlH9PYf850OcCi/Sp+9jnIyMLRmmZNPkq2FnC6Y126QDatFFjjIYjEkKao3CuMNnJK5xe7s
mlHw7a3ciBtKpiN8E/T+B94l3f1HGSuT9wZKVWkpoSr5rJUaEIFh3uvi0AWndGoI46Pv7ZtIbXQT
wE69lFG1rZ2VQbGOouacw1/RIk1PXFsi8pXetw6VvGZMoZ72o9nI6MHy5E348oqaeLgGqF04hFPR
0jJT5Kgrd9JnsvkpLCQo4sIARY/qRl8DJfN5bo9ADsozDLdx8DPlw8Edngqe8zuqPsU6rshwKFW1
6P21oGAfki6MF2lER3lJj+OEzntaqGJrci555gZLlNvccEiV82tDHFxupdjq01tugD4Zlzr+6Sff
EVSrgH9ObCZOpqkNk+KaT+UiANoL7/ZJuPZY5TX5CqtGPbJNHP98q7ScU8222YV94nudjIoziJmP
7Vq1FA0JTx85Bd+GuET3yjtKZCGQZk8oGYNgw6Do7BId+Sers70UvaOBmV7DpT+lWRA1zVJesSQC
1uTnGSjH37vI2nj+IiE9sWeBTFUJAPq21SoaixCb3aNC4pIhchZeDlZG8ObX9VLExiX73Zi+/vnw
PIjbGUC4YgOXrJIEaRWfGBr2MAHurFpqyZYlOaNqRp5AM8oD3UqrSLJY6iB/8NAZ99Ty4mypmXMi
DMtdakRDHAhejqnvNbEnbOAUjGnCugee31TwNYOavN0YW0CgT2ohVldX58BP7He0jqyHARopmMO9
2K2TF6zN8EysEeVdkW2UcF++IkkVbxrT8RtlCVLwlXk2YjAvkI+wxvS4gNaXbec8RRa3RJaRRaxr
98QMPGJAcGXe8ZvUtkia8eKdp4SUX1LmNlsDsu1lqI7b3UtODC/90hIqCKmTZpIx6mkG754YBMpE
Cbp3KdFG8ZEjdfkUIIfyeWB3kAdDCH7T9/HxwO3uyxuO44FXLYkKpb4Z/vmaCGGagw+3dXcXx5cE
k950XrebidKNCUU00ExDNv+OEM8ezg9rBc3Qxi+ISd5KoWDDKMBnNGGLSofNx19fxXZLVBIIfUgf
PNiR5ojY6d6XBSPBhRM9BSvk6sBRhsGQaSrclmr17TTeN6JvrMVkBe1Nwk6w4kC2F1fDf4pyNEmK
qUnYtAybKkEVqD+UR3DB7nP6NoNa1ZL5OsXcJXDcYOCqiitiAXLBKp2dCGQILMY0mRAOTqI9d45n
BShVVaiNyt5RZSR0UBtM9ThmanNbLjHn/zlorTxYlkp8jF5EOCA++t2YSHZctXE4aPa0zpUt/3dM
RKeQVoRTihy35VJExNyME4BnnSbui0HZHqzC1EJLgIEZnQMo766W33AuLbdAKZoq9B7wFvJgV4Cl
59ZPwnl6B22P/5nJkiEr4D5PBNLlv1oJbMBftDxuPnCXg/hwov+lh74jbZ9DZ/Uwdp39zm2jdNQb
3XAHGrugxMpo/MYzlamukbEX4wCve3kEo23hIe/41ED61oE+gawTu1EYjGPr5c+//7JtTa72VjiA
JWXm588WPiS8Www8/YQT98LVsUTuZe+nPYSi/OpJQ7F0fe3Ip+G75T2ijToLR7OFfe5OduIULo55
etFmOKv3Xvqk8FmpS8bfqp8YlJwdrUVu+MurHMa1N5PQP5H7Qze7Fsf/8d0lg+M7tLwMvitOupeP
lCkWldsVeQwatu+SvLVagUlLOWfG1WKYv+eEzTKo/msOxi2rrE/JFb3lXOC8ClFF8/v/59uHHHjs
4D3H6msQBA8T9ZgR8+I+ipQrGrcFdlbCS0ar6kgisOcqxXN3FyV4jj/IHpqeNWVEdX263g/025Gi
l2fXglrP88YFk7Jfws100xgXODgDP0xotu6sp5YGAe1GM96iqk3v+4DkVk+rDD/cvZ8JLFXq2d0G
CKJJx8IzGjvjZSM4aWAjBiqZ1CbFfYm26YdJMM6VdrjBZXkx+1QRxIDKLQRbLPoMcUJtrWHaG0+L
d5NBrp7erLOzrRlA7GkKMLjdLg/rKFBo3V6sVahBIBzckuYXbak26gBwYZBD3lbipWilW1fn6Scy
3/YabkCriCXke0iTORWjHJzARBHU8qsAPosyC6AwZ64UHXR9rgK87bui0ZKWP9mhtqNz8p+jBrld
Ui1HAkSdGA2RitWRVFym4kSchPzsIY0FDEArDZfcWuBuTiOiUoX6pyvKE5f3SpK4gbFX1cKpYH6A
57YX4lTZ75pH/wvLEjKQ2zCp7I1AGLdIPie/8xm2iPMs8wg6j1A4W5ArZgzweHu3MBUIFUeE5grb
nlS4y10+EYCs5uSj3B6qpNEdICEawFk2hct9Rn1GdToYNnai6at1pi7qXCuD+Ub+9wONbsshBfyo
EWcDGgJw518WtZXmAqjTmfBw1jLfBXIC2lnn/yx7uf+G1D90ZcO1Y0s3D8oSLuDf7VsL+woxNOIo
E1FBuAqbzRCSGopDzp4oIPjxPMgHzme7yl7Du2uQMq7T7v6aLgxEjMJvEb0/ViBElsJ3UovDF3wz
r1shzus16LkfGd69HFTcGgRzxC64DJ6ruTp3a1HJBTjDK/AGXAxKARiCEePdcBBB/J8AUU4WFT6E
ade1OW8+jpkhxMoiTw9DB1GKGW9Ad1OS9WrlJWhR84et7CQtZkUH/IvZjPLZgNtmt9chy7RSGfb7
d0UW6sD6GmzTFx+1JFm3QGWRGSoh8aKN0K1pBKMPtTnhMJEQP/F++SnTpHLlZCGW1fulepOPsVw8
Tl2NNMBzaITId+v4p4SmWbjn1mJgM2Ivi3yEQvXO3pIv4xeWGDLAbs0oWAzfqknZ5nJyQGPKXien
MQY0VaJi5746QcwM/YV4D2JvaJxfO3erCVKqndf4PEtuHXLcDfbxqX6D+ybaK5+MjaSstYXwPdoO
tOSHBDbhiejDuIKxkGsblp2KksYh6MI+uJe/B1RVPVL3SjiWyxuIVQ+Wx2ym8SYHkAKW/Jb9GLDh
nvR7Y2NKID0JKU/2sP2af3gr3iKp/vW0tMBbAzpSEaPV0oXcZhlPelR7EPyEZMylOYaNbbsgq5P6
pAoS5rjNd+vSvTtCVtlUJf2hblXSzCiN0ndNUfI7mR0bIQBeghWkCbZk/dP2q04Rb+mAnCqLTRON
UCAUarzI7RrEN8oIBeay0pXnryB8wkVuXPvGnQZnZ7idNgSv39gWHHEu6Pd2xXREWrtvYauQOOMR
zpTFdA3Z51zZQODKTNIBnaliEswh7d47QcANueYuRyFhSeM3o5n4knkSdztLdF87/SxLtLSBUGBG
vnVfN3VvMkrj53wKT0eq6P5QkK6zFMNUlxfjdTm8mvjvrp3rJ0r1vV55lzmhhJYU4ZsZfHmLEC27
vk9dtNiQwFFiA789XCkrDshi2HLngCA2IieizoLqT3pN/JhkoyWaauY+QlML9OO6xyJaOIW2UV3t
Lf7Qr5HVKI1Sklh53YKKC+tzxsUm5xI6DVP9oDyxs5NIheh/ePJMsSUN5Q62oQKMG7C+4tNxr2Ga
xm3wDovvJnrUI6oJZZxWCAEh26RNpVnzsuqBFQ2r5cyY/8E40xdGgT32OHbJWcs7IIRFf+z+Na5a
1Jc+etkfBI4eLvTky2FwykJNaL39x82IdjBo++BNBluWe3NjRtR8CFyMOU5wfaXKusyCovl5gYaN
rkbOBzjyB3FT6QeK5l4s8a/d6ce7+dR66ukutwf+rFUtm3ZOPVG3j8NwMMbU3HjHTMmppfXYpTAO
IKkYMOrIyJKiuYhzsiFLod92TXsW0B3IQtm1biEInw3ZeZxirutCMsfcfPohB33di66C/XovovTU
EdYDiljkpuQUOFpSBm9z2r71JVwX+N/s+gY2sQpIGhY6VvvvnpWA/3Aj/sW8jnfZ2/lSTZUq542t
L2+3yHiZk/V7wZOLIJ4eA/J1cIGVOSPuSda9Xq5e9gK0SWgezgs7TXv4Ppc0oqQBoLOlph59ztTp
AwokTSTxphOFqZG4UK+HEYflMqv1rISFX3zp6QEaTgEVKET8zmuim0hPMjYNv/Zi6EkBppFO4sRA
k6Nolsrpj2iMsZ2ij/LrI+RgYM/oXp0rZV0eF2Djay76X8hCj12PXf3j0NyMF+axqmaejW+9li8H
0ex0Tc42MFrNzHEZ0Ip/FEJa+SjioreWVMGtyTJjPljrFdXjDbPJk79f2bH9FPRXTjmupG/ZA6PF
088QpSFPUMgzdi9CA8OYObtb5b8+LXUs0c11GNpyo72Rm5ZKchiEKti/Srpr7uWZh3aqscPAmF4o
ilounZBwpy4qadqKIWtUd1OHnMdHfPEFhYnMTHwBoPquhVteadmXQvJiFxBYzd6BFJLE93SE7vgg
TGaLuurprx/E1mplBt95bqLBHU+6E081lEt3y5g7djCO922QRkm9IMY+js49yHVbIl5FWpZ260H9
bjgVfXshO1zDKgjJ3xkRXnLVl/UsPSxh4oZGrh6OaIExvZbQ6xIjjvD7BwRTH6L9UmTZviv7oTaJ
mhffkNOyA99wROjyBlnLAmurwNWc90RI2d6enzmi4hgxHUd+0+FY9NqdzXTO4tCPPMUqUEFygIf4
89DepqlCxbdTtAg2MkgeySPkpqw01NMtE3UPAiL2uWMqHSu6OQWbkeBY5bpzBn2p5Ol1KVjb2jqM
+sPDRP0BQhZR7hN/grRV18FtiQMmsozxbsbQxWXbyEriFBfkZ7JN3mXHRbOa/0M87eDcAp7Oz0Nx
o39BoKC1HRojkwbuF8hTy+YJJSAnQ7gvZPzHPAlOd5U9qn1FIWipU1wG8gaLei8nOoW3LkxsV+Tc
vZQO/pvVnlxYpjEdVp8LYqdVZCYK/KYnwQ1o1GxHq0bK0x5xYXbqcz/2AsQQmRsqUGYnuRGqkczg
3bezv6/t3kLOMJxwl4OG5jrsTbfzGGummytjhbVkVhRngaoDyrO6BquNc3DSJLkq8GKKMUxdnxBo
yvdfh+9MxD7mU5f+HP1pMJ2ZsgqA4ccFarW5VZ3alGCIDW+RlfJpeJ/UtCM3khx/ZmzfslA9JSsh
EytlMKQ9xBpM/Ez6ZqKdpbB0N1bliL50edX/o1xffl8KRgX4XnErzPDcS27EhZ+x0TZVrqTT64RK
IGbbeBil48Ta8RCCf6Z/MERRgT4byVRJnz37BvWG7wQUVxXYOZD92l4tk83Obq8rjSVq/JlLDNLy
55ZFvMBTUYErc8XOZh0/ySiq5OldvXcK2CdRcobqZhwkCAblYLqW7lpc2pUPGNEkJp7ILVwJilMX
wmebhBbWuyXu354Hb/LhpgH3ZCm2DPVSQ/g0hEKEfhRO7GhA8W36n8gBF46NjQJT+gu4zi1q7jCc
6B3NFW8d4LHfsS32lFSfpCu/kmrPs1TZJ23aReCWlq7QVglcuCalkxUEzBlRBJZEOHgGiblx9ri2
bFZt8KD2/ZgGih9u+PA4fOlE5kOT5Np5uOB/6mPwTKs8JrdaTAiAHdKHTj2yAHblyOONWQMhYFJz
fRZ1AKcLw6MHNblTip2+lEC5zPf8RvkMlbEEAdqZRvKaRpqiF0GAhlMMWhvqVzHDyDZyhJ33B+/E
v4j/DbSCN4P8CVievhACQrPuB0eKVhnquzk0tsfnhELaMdJ7l7MNlSyncAH0rQb8zFkBLoINbRzU
WNAGYW6noz/6YVgMfb4gZ6GJ6rMS693W7IznGtdhXWwFyiOemtSWe+CbSgHEkp/YXf+EZJnaMSKb
4Mu6VOVU0l4IWxbpzz3M2ryxZwUg7NJk4P+oIxP1UOu8SckIRdklw4x75f6iLlhQDLcSkGldVsEN
boJ8ChfKdb3OwV1cTY4UilI+TUtiudXz3MVRnfTieHVT//UhYryo3LPWB70Dwm/k1jotZohu9Q8m
tD8zv8dVRwh4bHL1blK0MOGtpi2L5O2SEYGs+ezGL85jxK+CjoUY/Q9rPSIPcLLPOO2ERRoycM/1
n+EwIzsvbC3P9nD/6ryjsMFik8wK5lysFykakqpCqyQyBkw11ug1Pqt7RSYexBzlIjv82bWEY1bZ
Dr+aZfeM+TImge6/Whca6C3uP3g/sAhCm2Ovdi1d1QnHT+BAax7RRXDB/VWIJiFDY34RcDS1KXvf
s/6DDILzOvbEvyA1lS2EM3HbPcMafw/jzKIFT/i2wXUzRrjuzIY/MpBiIFJ4CpoS1WOoAuo7ygTP
u9oU8fso/aV0pwAiFyAzGO4h4kIbenyjjE4G933y7q5wiaWlXQf4nukK9zsxb24J2ULd7gPvxT38
KkbnsEJI5nt4nPYMUtrA6/TRRmonSy0tqs5YXvEc6AJb+Dtgm+/ka01R3apOmp/xOIVhF5dBpbke
oOLm56I6jNoI2wn0LbKFioFo6qjtZQiDoRvCYKekjP4nO63JknJTiAtlb3Fjgsib95Fn1uZWgh/P
2ZQVgDkBm9yiCxDyDH2K/2hYoQ8rcOp7N1pHfQHvo/NtjQ0yLxu2qpGJVumEFCpZ3F6QHpQpY+/t
hxVlOTI3Fob2ZYxVB9qo+1b2dWAYWbjPbt2MNPhmBAvUurESTsquc0hu1TgL0DWTC5uUItanFKzc
9tCBkFucyVflNE0cDNiPYStRKEddfc+S6tB60Gp+anYvtIOVVukUad7WhluS97z2dwhLblhFicP2
dBvnPKg2gwY2Q7TQfVN3RAizj3wSOsAWzhFYgapzEnMriIx3Yg0f1fdTtXfXXS2YcC3E3I+8ZYj2
FOWXew+qXYmKkxgQRlRULo5UX2tsjFZa8Dt74xeNu6I1ivF+dqdAPXFPKGb8MrXm6Lr5FTK2P8Ai
P/NpFMjnzskL0+pYTDeEZqGNyXmOJ3LsvT0JLpNdfZWvp+X7wauaTJpICWk1+XTuLI76Pe63cDBI
kikNEcfCrulIAwBFFXVP9AAdh1iq1Ikiu6t4on2nkyfFBPKUWZjUIVf8IN/wclvozg99r7foYSWy
5W0FWzfxgffiD5ULFzYG9jqkM4jiXWDmMnfsGCJ04Pf/zzlqorcXwM5Td0KmrSW+1vv/BoQHcjAY
kEUv7TZ0DfOYoeSDlhKxFcWDBEC8K6i6QCAWeRV1SXSs+v6a1uqTlvW8T7IRraTwz0IaVBWMA2r7
scyQUTbcm0t155AxvwlOe8WgmeUeMNBf2FUwnPh+Q2AOqVCnaAtMnaOSgSa1r98vS3tc6NmH9JzU
/Il551a1LzAuOUfDM0v9CyjHP2yeR9hcCojVu0vSQthfZeJG2ou01azdDWqeJc7Gtq+WPS3251JG
S0vYnggwfVakEH2Q++g0bhI5jyoSGzYnMX6fNtSNITswXjqY188IepUClij+mkn3mFFTzYCtO/Ku
KAEizUCOKwBu2zjTFGhYZq1Von9RwXBaQPrg6wkhtUg5PZlpYFd/hdpvau84S7O75uE3aI/xR3F1
xO6rS5+IrKerUHmyW0faEXukpQLOIkGK64GtxyZ1bUki9NJXX2/m1YU30Ud1is4vArAORmlpW1dg
wV8lAhT+411Y8dIQD/jgThCHsiVPJVXtMYohfOFN5cINhvFRoy/yxbVpalsbduNyzSlXE7ZRkk/y
bIcn5bfetJ6ExsbNnEfJT9ySbhT1cMb60RhoB7/sMWyUQ8RlAc9utnSdwLonFldWf8Hez/n0hx/q
G8NkASNYM9kj38MIXeUBMwMk98r7i0yVTc8VMZi9xCPEHoMM2UAUYgK4u1iFFcxlrARY1BDHZ6nJ
OCxAwbrvN7VUgMUabf9xX+ykt4HvJIUelhwhqi+tI6Yy0OKNnRtzpqHgB1G4pgBjkLdfIPvZcj3C
YkUMvaUV6pSTQaeKTNcBMlGBnsiCWH7sCoOuvS5jdIWaWomS9hvK8d9ubfFZ9jQPKqfAy8iZufcL
dJQJ90NUKAtiTKPR9gikM43zw0ul4IngaAEa5oHak+Azu8js6g60f91xxOcdCCJK5JcHz3/wAUHU
im97cf9XEMbCU+AeedIDMK6Leg6qZ1YiWEFMOYJC12JDQzxCVaEN7vN9C3oRPTBaPgjLidQidCl6
Wn7UtNCwcrzpz3N7Xs3mB/KQjTsXsGn9IDh2u20X+1jMrx1RNr9w/8CXQz//QNJyX5TNPeTp3ABe
YSpjn1Btw/sXz2LJmylwbJ+7xGNLcr5Eq7C+xUhpliSL8OLqwA29NwmxD+vpMwnNfBJqRo976d2w
Lt2fIOFxQp19Ik7YrauoT7S4QjmFf72Gfz66sUtmwxVd3X3JBCCDhzv+iW8wx02ykdcK/czuQzxA
GnmvQAIyowpAqjpQuQd+B3ZwvEpw/E1tHYDk5GpXFqF41BbNZBwU4mLnGFzTyvCy97Ka5mysDHxH
IXp5n8z64lFobi/Wk0K4pRfPYrs1HIPx/D4RpP4wN51pqYP/ffoWoOl4PwEtKFIhqMqnay/R0Llh
rQdA18u+eR6LLCEfHnaXx7e9x+UrhHjH3IIpAC1/6ViixWnOwzjqIR/B4s2XJr0h3NWoRXOpH1wf
WVGP2lBtbnSt/88LnTDm+0mpA0MBTZKbMFPawQf0ihcr8diKsFfOAV3XJ/luKNy3ZCY/TVOAlE29
qfZaf6r3LAQqgK3SBAVYXWfztK2PpoG6tLkeu7eR9IeSn66Vk8RgT5lZeMDXa9zrKQlzUFT/C6xT
Cl+FvjBnW+LGOrJRKc5cpjRedhTgSm3qjxVCBeJDoBp2/nr2B+SceVALvdXoefHiJcSKfN2Nrjrk
BIlRIisVdhSJi6QyZJ3QTetCTLe/STeqR0l1cAqgdmlYzulnnEJS6IJrA4DqFvuqekDM6ieVXv3Z
pi/69K1kj6UIyEYLVaN3iDVJDVbip3NKDza095sHK4GzyGSIlPyCKJeuxyblPP1Bve1dcAHVFnBy
W5noskHtLdK2VbaKONl7Mw3suIaLE3+TKgG0yqLWS5v2xzDfQhzzt1x1UJvhUwtIz4r6QenxgZYO
7/FUH9mSiLI9CLhvI6MqTcpxG4dMwIIfbqf/8cQTWCY0z69c8KQcniAJaywLGZGhE0Bfnsh37LXn
VvQOifoMwc/RG4WsWV+RTcTFhgroORO2P/NuccTko+jGJYe264J59qMoUhDxizvm5UC/s+UczI/L
NMXMp0vNjyGUHRIu0bVaSOAadGG+NZEPwYfTynHmfhqj3WKWVpJe6bSYbl/Sh6vJwjuo9w80/XSL
rX1bt/VPLRPM3/x+qliWABuLa6BLcKCGG7GLqxMrBHDr6KFYysy62WeeI7Fitx8tMMfZRfvAMEpv
A+aDMJhARIxUxi/FzIL7+r9dhEZ2gmVdOolrWw2Wwd0OqFl7lNmOndRnK1Y0Yi+UMwNX0TLQfI5+
bbGUzdq9mtf5qQ5wbHtA5NcOTlEOoag1nTjPqnpJpc7GIz0ePhyYgDR0+jAtHXlqb+7/A6j7EGUB
V9PA/kPy48OZlCHLwiQL/rnNZCib3ZpAA4xJFdFV1WRAWsfwRf/8+uQtCi4ew2AInUjZR04BMNjU
BS40luSQB3qZIAQB0QSVtY45sI7jALhjLXcBpkajyvW2ju6p/LvCp+LeRs6S9z+iViyWd5wAuVAZ
xTXiHfV9XMrqr7FH0ld6bg0tGAvvZs4XQKu9g/4qqesAKBW+1LyACepfsiVsB83me2Qdp854i2LB
1BQmM1pcnI1/kPwCQ5W252cy8auk+GmYxy9tqPhxbUR99xUIYxNewaLg4EqivhjiWXUSgDJIb1L7
8xA0K/tA0KckOp5an3Q3jEHpB1SIScg9vG4Mx+JYBgNeln4tjmOHJizQ81YspUBZPyUv7PGzjDcP
v5qmn4xkNTE6raHqWLg6bgLXfJsQoi85BoabIasKLJpfXgWaATHtBi/CQP5TuCwGpxv4KhvQjvM3
hob5ZaeyAI3HZdzwbf77DaztqtKuIpCZNhabBcJ73iP161nGy9JFkx0F19d9ozkdTtw6vZxM2w9/
Mzv/udhteOzHQmN3y1B8SCm1UdqcQ2rEav14OqK9vBSi7Tvm+trFQ5ARRXf1UsnigPGyctpIlNLE
n6LYcxCXEjyMeC7nx2/RJB9KCBvtiPnWq00EAYBxX/QmEOyWhzHYMbi5MCaA5CzKyKygJYGt0owa
3p4zFBGNf8g0o25/mdtLtpAutGIFIWgMda1mDvCrxKhWpTJFqtsqUtplXLDaJX5jidpyFlU+M2qG
G78aUA9Gnwk57I++LycztEN6RjKAd6R8vi10LedZQf9fIXEJbRHD5ROlu27wj12/KF8k22iiEqRA
0B26PPOduFCJWENLiMA7zJ2QCPF13vuMAduFQ8tRincECzboC9Oqv3+7+KPZXlGvtWhf0kVCvmjG
GC08sAhQajuV8q9lv7GST2yr+kuRG/mhDayZlCjBGJ5Oe+1JQzftpR34O/3F/1DbnfU6vtRARSIN
pBWHXkYPp5tLF4h0+4M08jmWuXcY//6rVaXvTB73tNfhv2PcUS4PPr5gssNfv2xn06genB5DH8O0
RlPCUA4gMowdJwiYG/Nk5zJ+WnfMT2uX7U6f2haoMLAEorTDhAhyEP1mSw48zjvlsowfSfib4Oy0
ek/DerQwDe35H/b9ZBJe6souTQBBH7tQdirItnZzGNd/TkgPhCjY1nesND6J9AWwZ4HOf+EubAqD
+mX6pHMjCXaUzmWxlErHo8vUapqhV+0m4nb132LgzbK/7gsECSQHIvMaZfdfeQHdxh0owAygNELv
pSw99jyjt7/3Ip1R4Xr0CmHJ0f7hbLVMVEytK9/xOSjP0b5yLw+htFbuYvg5yy+wixwzITq2K5U6
BuubvGoE33idWztMnJ8p/1DZCtn3NrK+muLnmCpZ3PfeF7nWSO3/Om/dT7IXQa0oTj/VyBPuBuYE
HSqn9g1kaAmNPZttZEpavWL9fvp7PnyYKPXQ6Mu+lnIR02koopnV+BslzuXE/Oj3hdL7F0uR2URS
hqYfmGx5dJoIr7n836/yzlDLkjOU3fT0fb0LkKRlprcQCI0PvzTPzzwVJH5ZRIbvRx3Yntnx7vri
00GLHD9KXnp8wsntgyz8ehGEU7sh01nxy2ULBYqfKPYA9MXM97diY/O9VoS7gc40W4eONGBRpvKQ
tgNbgSabREFsWvGwm9YMgOro/79+UAinCsPzNV1uuzJIzvP95H07TWthDhuQLSMYY/d+pzr2A4C9
f5v8KKrQBG9O6SLLjNDTUn5ZM9dwIq66FOslms680f0NQnKjucIx94tXma1pVBRro/QjT4yImwCv
DoZXSm+ULnKNpbOzsjU7E9uCRRj26j3eYxfawIfYe7ubtA2Ml8KaTgAV7bdwDu0+ZSCwaJBj9gJJ
mRrBrxciuXg0+D9UR/ky3Ckd5v45XtlDx2TeOPlwogNqk2qe0OZ849DwqUGMsrJkhH0Yr9hUJhD0
hCgkARXobLShUSJkB3tjB8rYCaQtWVey4I/TsGdF7joUI0WRegETDcBIYHQxTuB8XAuIPMRXCN5e
Z38dQ35wrn+tt5lhypdLqirl28IIwyTmSX7e3EhECi9XYNVoCmV6+N6sYUDtIlGkyJsBcDzm7a2H
RAeoEr/YdhlJ+NvBBF3taP4e0Hei9HzFXHKQkU3oceKkwTmUDwFjdCFPKQs1lRUOAW6jaIl4FrmI
38rmnzJDnZ4IcgIXKdUHMBFCSn5CJN6Hi7ybRsnkfoL/rn4rpW99YyCnBrlEZSg+V3wFSNkXTwLh
etEqvVC01WydyP+UQURtXACZKSwGmpicB/VxNs7SNab0Z1BGeT2/i6YmUzNNgFKtFlhS8WiAUSLY
ECpo/xB2phM+2+fCidrNTGxenCo//JkS2Jc/wsPwFzeeuURu8wZzvFpY/ySYUv9fLsn6RwIhax3G
IkfI2EEcCowaJvXwvYkT4L4wOzCeYt5yg/nXsl++QKcfdXNL8pM+x+pmHQ6qhjlLKf8d7Wr/O862
qvU21NAT/NhSc1Pcp5JY42kzRzMK/9jJmqgqcdo//3t9k9S8JJREzOzyJaw54wClFQ9bYbGEettd
HrMlOfIOWUsdje3nq/pQBIc1+InFr0H/7Jd+sutTVaSriwjJ00qCF/SWlFLzYQ7ers6pyEcY/K32
AY/JN/KXVjWm+CZH1nseyvNP37NIS4IkcOLdGAxpQo0oo33m3LpS4kiLLo6SsYCEO8ZV/xqvxK7t
odWgXkN7vOX18s/ictdqa+Yp4QemmeKddwwBCHIAJ+cTrfEt+QUUIDm84ktC3R8QZINozlZPEx9b
Hl6y9gn5Xzhv32y8yYpUAXFS5dXf2uMAE0ngp0ukBNY/Um3WWynpU/J/bW9sjtwAA0DreqBJu9+f
9fDvk94YG3j7vC3QHmLVYQD6vG2FwPI14FfqF7aoxmnVlTpLzWhiznuwcgtYDzZ+XOxnzhahH+oV
mr3flHvSe4USXSPgQHwi933LtqSm1GKgQeuxam5QpDaOHo7G2Sp3foYBal7k2DzLn3zCj3vL7F24
pStqNWvIqPLA+SPx1ffENBLsIB/YJH4H3fQ6slOs7F4FbJ6yVySG0NXFrrh4sekzkq91N0NKFrC6
iDnFfAz2jQUd4yIA+795OqArDy2lHM2SwL5VutXVgesWhuZOef0B6zgNJ710ko6fZ/XRnKxgcCGI
TPrjp72iGXkaD/8fuCSW1uXA38k1t4qAJontPp91jdejqyxlDV7itFm8fPQ+9HvUuinLOCiUIoDW
2rZyiBr9jqFE7fYE7d/RnX+qUvZygfqAAGhwbfTZDjEzft8Dy7TAufi0B8BtZ0bKBuJWUixxeGFw
Uu4n11KG7ogmAu2yDJgwGfDmx8nXfRsSY9j84TGN3eqzPdMM7qovMvXPV/caApnqQhVL68bVJGW/
G+RdzcAKcp5+HzeD7s2CSXUGg3s0fvoXW0LVvHPlMze/2ABw6Ae8EcCRglQ3Z5CvmXpptqEz5j/V
PZQF/iaY+XMr2RcvmtnAr3whrdeLDHUlka2CyvLhKrfz95oKBFs9H3/QIkWoM67OZeeAhBIEbOU/
YbxrciTbIG1cgzgWTEoisivYVvgfXIxs3QCPnPsfMmhAkbdI2o1zBA64CXFP+N4KMxncmhVm14KG
wexMp4FkAE6I24ec9KA7Zi8NTfyEIXKplYWhmvdzu/YelmvzRu64b56RGE5XCB5aMnfx1OjN4MV2
miqK9eDnXjlgYEG7gppyHVVbZYMZurX8Csq5UdVdpHXVVa4FxgYh/jxRfqE7lLv/WTNuLyLOy9G+
hGYj+XHvf3kRtI9by4ML5iFNb1P1knVJjgNhqArbze7iYevendPXy0AxP0ZQogu62w3s4o+FOVpg
SmMjxXVXoFhkQMqAMsBX/nJGRJ298yHuQbcXQiPa9PnRXbnPXvDk84E9NfPiFw47QvgPsOIjzyYs
1mTgnF6WXHdWsUWis60DHyvpB95c/zKsvuNe/Mzv0Rx6XcaXV6qr1pwVskAq/pSPNpgebjgHaZLM
bSVS9R4NsPQedkDH2XNAVX6jV7zbLBu0quE2rlswm6LgP9o+6BVXS1P31pdyBYo0TLrOu3XjTVxX
7nYcIT7mSw6pqCly66uMqg9Q13DDLvjutErUKOVPVpDfnv559dHUgJkuCiwQWC46em8NvADI7vAq
W3WN6zP7O/qLcg0/nfHVsapwmEqDob7QlOqxH1Wl6Zg1J8LT2lnb0rsYkZY9N6GGRjFXgRlOUkhU
Xqv8fwcqX/Nx4eNSjeWi0siWL/HtcRrollOd7iv5w5d4tGOX7zxRxo2Fmq5n+v6u95WQy3SkNjZ+
jbOLmm0zADcO/pG2drXwR16A3UtZguwNI65oFQSpEKPD3sRujKtP5eKIHIOYTcTJBr6Qfq9OdoYB
rOwWaJ+g/UdZNEuc3VpC+AwB5dgozqMdVx54ZA5NwehRiDWj5DWobv8t5eMyP6VEPlfTf6ZMMRBb
YUq87ELDBjNueUH4o/iwyXgjXqqj8elwt92lYyDT/+cqqWLze3bDAMJ325VL2qOW7xXyDUCXuLwd
vEveboyOc+8jrbUQplet8YgZjULaKngBHPjhkAIvtSLOlbKsB3tk8diyYhJGaPZuBZuCd4S06oac
DgfKghSImayfKFgmC5En4T3yz6Jziey8E88RB+EyXwuGqPfD3mY5Od3QfBK6YL7b3usL6N5HPSPv
5D1vYrVOpvYj6iBTP9KKof9XxDsHxePoiCBOSnoMEj3QDZ8QCu2DwmAFlJ1Y2Ik9miwPkH9Lk6iI
/gZI9Bqgo8KYcgImI5xqb1RPYvhLZSOaNrK9bFY0tUyCY11Iw+R+NtBfCjekEhKW4kXsyHVhkJOB
0rXwoyvnhdYqq2tyxBK0arFOtWEP/UgCoCvLG2eZKAhp8uT+3GMuVl+A+jBEMg6dAp0OjWhUm0XH
5fIBaAscEsIcJa7phS3Q6qacfYCywD5wGfxDPJcybtVfRzd7vdKgg6j7+xMrKciyWbeuHxsVNeF6
xKNghmr7O9TNVlgrgWbQ+iG+Z8tZYUP0iOc/IzJ6E1idxaDiKEAwexX4/tIE5Zs6VfIeDzRBof81
hvAkebiqz+IWC31lk2OPb95uqIZJ75v9El71eU083oGAkRGz+Rswj1Pf47ZXY8S4D2Qaq2QI5S1v
g+6BzOLjL5fcomb51I2ngjEdHNvKeKgqvboECo3FF/h5DiQJ5XpFDav7Q+OLGp1hTHTV3aCREtCq
vmZFGTJX7eAhyOoQ0JUC//g5m8K9YODb34yiStoyNX3nhOmQzth9NnjpRs0XlQJvjCbUx3Px+IaA
OnbIzUSIZoFCVdFdhVKz15Q/1o09dDtwFaUhcNmNjFzhFc1ZF0l0QeqEVLf7z/lHDZFcKDlKEctI
ssbqWkdikuawYXYHw6Ki50kTY+SxwsweElSkWghCvQpYg8mIy8RjHnPaOlVKiWMigEkiVWa6J/Ye
sdhWbmjiG9+EnNTcYAamtRPLgurdCAgLx+MIrK6xWQZ5N6k3dRbMc6PA4O4AZpytLxPuS9LmaxWZ
J+nBMr5thbHakz2o23QY5GuGQq4/UJYmGc9FqsaBWGsSBXCrGY/ZZzRaVbVM6R04VpEbKrusPaVy
ESBl1RhAfYsJKBJK8E048axlZY4v8M9FSgCkbN/UFMbUZYJJVh55ygRAr1yVHSljqvzgoc+Clxkn
ZqNiC7aYoQVVY01aXffS4U180tHFw7xx0XDQKFiO0NHVFll0HKQjZJ3XQpyUi4+suM5meZ0ebtrx
18ZRQYqImw5UyxgD8i9wKS/9l/Y71hJoQmheKjh86/n3/O7A6sj99QqyY0+PDu0J4dlQp5MEzHnk
YIt7xgjh1n2d9fcV4vnvDLQmgAyj1x1F4oePczLNDhjVgiSZ9Ll6wwSyB8MeW0tv7kGRBVPk+Rne
oUVHskPrQlyFyDSgP5bcZx85FIQsncFZPFkh1sO4bio2ry6nHuXcJ2QdMb2wNykJVt5kd56In/cu
Drnb6XFV4aPw17EeFVNuxbHrqDKNzD23YPXGy1Elifqqc7HykCi5IBqTNmSXIfVy8YPPSksrNpIT
8HvVnCLyQqmYxDfQyR18rz+PysWq2bWFJ4yc0GOYWc/IHvPjlAW0bvQQ8cc5ACm9QvsTAa//5dZU
VzeDAdr1qbXGQ7aD6BsTvFZ++T83a62ntFv/VgHZW/y1OCLWb0CKaAjZgvTdQjTZTiwEARR13ixm
JZ4rewiN5OG8JoqUStAVn3xCbw7jhEfJ2uTJbCmKoXC5JIF3RI5yL5M3SDg93G+6UJMrlD52Y5TQ
LNyHL0nYjLjJzOw1hd6+5r9ZCg4dMwaNav+KP+Ax+gdRVXQwOsM3zTs7uoHpJ90+QE9yUHVyzNZh
Xk/NgjZp5gvaYNjhlePgYY5aZzHF/m2nGqMQfUT66xelPr7l/H2Yhx1m8scEVukOaKD6CQ/U1dHN
SGQEBV3xXl2kOAKLx4XJckYTuClPjHb3FmbFLonu3ThniQBu82wP1clcXSicbW516qkIoGrQu6vF
/QILlz5wRz1B9YNH7xN6wF2Sg9UuHuFxyNYYm+nPRXXVQQgCffNMZK8UJ/lS+xBanZ3+k+x5KJSU
hezIXcLq3rlZs3Ml+ScEhHO8nuecJojjZar0n8D4f8wRp1jORgpQjOHUkWdfp3WT1Tgpam87fseZ
hkGOUo4e4fbrGYcX45V3f4eu8nkFqPnNiOOy8VUj5uOmJOu2hjl+E5b0/h9oFdv31ySUkhklMwTj
1JBCOHjV2UqhkLLLm8pQn6pf69KU/a3VPdudoHpPtmGD9jkpEN1NK1Lk7Vp+Gpf2ZF3tEHQHUu8N
vg5rn3B2o442vJQaOxjq4ymPdZmdIORDtWxSYoa6Gm16p098I+orMHoU1NYvVyrrd503LY1+tbn1
Ob8LoXdUSPLboKMQ2YmgMPDpVP8VCC+AHEm2ooeZZZ24az6n2mCXJfyYwBZ4ajzxgb7XYo1K6sU6
ZzYJ3CZnwqwfO/Yl6fO1FT3+NjwIRh3mZDRdy9M4u/ne45lUvM4ThMaeno5/PxTxIxDgBU6wHjjD
vZz9QO/yiYc6FInuugvC2ZxSdVYBYHHx5M75wuWiYF+pKo7XxsvEoc7gLLx90eLlJ1izi0yHlnPz
F6ss3KOHz4zZHWhlJIojh978jY/COZwbIUdxaMSO2LgfSCJ58jGt5YVn13LKUh3fh9BAWj9OxOJG
pwCTc2RVv5xEaampdx3F6ZQ9XVNgfZZ7wpWT4Y2RMoiV3RPLN1EuCl2UB8yTDmFqLe0ksppbNZ/Z
oCwMBwzJaugKeVJd9oVneH1AlWyeYUMUNPEOzXs+hmXO0/Ax/VrwhFmjdXq356QGymmaezmHLejy
mdKh0IfgKjKEzEYMN0yuLn0dmctzwm5vVSrdySsC1vR26XiBC6tQpkv0ppeq4OZjBhJibQmuGO62
8V3iKX1Hn4vXvMwGRcnxQYdSwlT8dYKU5nfiLwuQb6FRovktjW+EpdBqG0/R/Xa1I156yHq3kUEr
oX/XtRpjWotaAWBk0ZwTg5WuKCd6hA6C2zHro1JR91mdbxUKJPMaEDEkc55jqy2CDovo9NHpbhHN
wvoS3nIGIOr32Ep7yKoT370SEOmMvsga+F9+QSnwZ3C7WspU8ZmRqAcSgDWO2pUb57R1GaDT602F
X0OODeu8iLs6nsAywUCqZFCLXw1e9JnXsTdgJmA91Pqno5PXzvLp0B6v15a04Q4qXvTLe5NbjU2U
HnYe6/xbMwOFF4lQhaT+izy29lB5t729GYklL5B55oULBU8fG/R0nE9xZA6WAQS/3e0qa8INsH9H
4+g/rpYnylfseOe/2SaCiPtHgBtQqI7/+kJvTF+Eg5wxvMl0Kd7SQbQsLHYGlyJ4UOBEHBPS/ghs
vAIv3sGcMd7IviVUQkMBGvcrYrGO2CXoRwUE4VXRlAtaYyXZI1TNondzIgcJVMWTW6+qt9eb/oEF
cyLLBsc7fEANyKTPj3DMXNhyxn+rbnKlqJUmHpur7xBZcMrBFelU4YMlhCispyrfK3jsD6JP6GUI
WVqryibjbe88+JbUJ5IGzdmSsY95fWCLRBvyblSnT64Tj8dZJ5pZVZsEA9LU8de94zrtvToRRoO8
Qt5lIEODjCXQSVqcoyuXGGinRg/HAfuZxdJaN4fnboYwrUCONcDqYpUGuEStbWtWRFxiN3u31OD6
6Gur7DtY8oxjRUrO/wCAfeE1aMci9id+mf1u6GHvPZgL6uhDjSDlCoWagrFz3fyNPdrxbSiXKY8v
f3hj9lgA3q1OXHgQ/scJ5XAxyhCWPC2lhadNRTZgq/2V0r7kwdTZXRctGnVJmbCl2Is/XZ4HKczF
pA6VrH9N2Jt3yTWu8/eHU3vFvM1SalGdpVoLeEb6xXAuKwa0wWpHDuXmBr6qDrsMEYMzthMz0Kkh
+M13E7EQ0AZhj/QVbdQElhDPSsAUj+XPgDHv/f6mYz6VymCVFtWlMYERDCXoLMAfzldtYkqbNe5V
1qK7AloG12iX4+AnQuS0ty3zxTLwKPU3rvGDAFE/RNQDa5KwoeYu1fI9Yw1ZU8aGIFG1vqqlVWdR
7sgNVLnXLFCeSddgG6KnrVJ3Jxq2yG0y8kUdl943YEeNAUf0G6j5ZTh66RbV3fsIF+WHSPZK7sq7
ICzooSb5Hgh8tanCXd3+fNS9ZzDTPMczAUmUmQPglT6f1gmsb3TR+XcN5+gLVHE1HdRiwL6CacP/
yCznk5XHhpWpFpnczTQPN5q7vGQpcCnmbFydUKXNt34N5RGCk0w9JSkBHersrAiiW1nNnpVvKvc+
3Kf0hn23EKzwJ0sQGX/Esx3+O99MWUq3XRrCpwP6l72nkJ0MPPhjcyHO7efnR7AGSI/dkjswKTrq
Tfyi7iUWce00QkUan7Of/q7iFfi1KfexRFdR9aRxXxL+QHct65o6EI6WlKjGpmLuyt1TpIOFRvHw
c1EN0/r5+s3pSrmbuec/YMnnlZSDJavDc+BHdE0pUgI8suDt5E9HwYXjBnxbCyMUHQVt+EKH2pI1
R7sIEumCb80OpFFkpk58Lq1oOX9bklGUdBQpAPpSp8TPttZtwedFE6acZ8+v04pUNxzSemZX/CtY
AXc+bnNyVn6H4QnCyzvW8nYMdClW4SAX6xEU/17luJv+xBRDBetlVz2b1YXO51KVQmwT7AjooYqH
xAFH8t2imCLfVtFbZ7hcwdvw5MdYyowjEXG/3U1vPjb5bI3a709NVB/WkjlFFJeBr5UuMxo7TvPg
/dAyloofuQl+6/ZQISjj7d86HihgoGTgW/dmaO1xY2DVPzoArtHcyu+bDgdIoT6TTJnO+H3ql1a3
FFkeOcTnRaKotzCd4PIszwioI0cozshJ2P8mKDagtEAV1ra/Qz3TujQLOn8osYE56sz04tEIH5Vl
02g4RPRxRjoCFuLmuvSn49p5SnS89VugYjOupsdBwbEUy/M4UmFX7X7SgQmbq743zA11bNYrmTK7
xgi5OKPE51/jDb5z8MAPnCxxBVLlpOF0b0n12SpC92sTHKV7ys3rBdJgwgLH+yhhAhv3YWN1Ss4X
wOHh8xk9Kf5CF5lzskzm19yf8U9JchQmKJvbefH1pCqWIbQRPDiLr/cqTVcR4aWY9kaQqNfyzPba
k4KKrABlURtEPy8UGOeWcrwtQMWL3GQgeibgsMVBYenV+KUgN2fmtF1NocrXg9meHwmxpEdvNnWe
cJyEstrqliFET9PFXLm1Rimmje7FV3pX6nlVqA8P7AsMU+AJlGKkCdkio3vusDjKhe108UXMZNv1
CApnIsUFp+EfItDNZlcBv1MOYNjOKN1kzKzEsN3I65DpWCZEJr3CT6MIG4sgXPMm6V4MgVFd5w9Z
wmhAZBjtuRzGt0uC/YiPBFgUg2YlZtq0N8QERi2nimqjj8S0p7jphhgBBjnjRW3clzvab6QCz8zD
hm4/Jfu03UMOQF16Wur7xd4SvE2j2a0kSSPsI1BiDZU+q4ZeYPjiZ8mRBjF9oeRmbGRzXc3Kt8Da
gI5w7BbsCEmv1TdBJRvh2JWQKj+MoMWv6OHjLGw11C0E43/HGCNFU7jR8XiAGAaFYj4DTrPrsfed
+bGpIoFmD/wGtfHUvcON/XbRY3rYW3PaN8k2mblY2JHeiv8JbX70HeSWUBvJHBbRRzSA/Ka2PLnT
jJUN61pKfwQbtLCLNmAsOTzkqebwKD75YqCJcSlzHszCrznun5uivSL7TKW3UvVqPDCP4yxh6m63
P8mTWP9jltSy7JwTmHZ3VVl24xkM4H0EZnnjqbIebUpO3H3xNs55wOazQgtxDdPM9/MpjXGnHhwk
Ak/q4AgWRMMa+/gn4LoVc2SPJU8t3jpFfAdKUEAyALmIIwgd4RKujYUNnw9EZ8jc/7xRDlxhUo66
7H4tmXsMBoRw48TgfHmM7CFWBkHdjBzU/6dXLH1YhTEjTmXH7Xq+L/xnZuYlKfOwdMNfGq9ijlMq
1ZWz7BvjWfRrHlDp6J9RoRhPjRiBYj54CIGpbzCxkfuCsibjHY4tUEXMtsQ5EzUE5sYmUyl/N1UR
iRMSsLeZnm4jG95Lqgb4aGaE3ddfVmNgo3/PZXS4fPosH0g4M5ZRl1oKMQ78sntxpvwERhMITOKZ
t5K+MCjF8aYNtLYjnfsOoEfK3QVN2fenV+j8p/NPzoLpoFIdQb4USYoIizVWOzeaXmhXWMAkILuH
8lED935dZmOMJE2g5IiZNiw2tk623qYdHuaQIEQCt0wZcW6hDvS0vL9Vu2UI6k9Ty29TyL2LrdJ2
JC090I9XZUqSB4CTrfQOtS1iikd/6r9p5yN+FOWZmxl0QJucxx2khYHnOw+JLFtysKWBLXLDsq/A
azAZgWKJTWuRWk/ekH0CkSuH9j42inqrkEIiP0tp4Ayia8ni36w1cSCBpKqR1GILNVI4UX4N41Uh
vh1lml0VdisBrSvDT+W3KZUiIHAoSgikDUP6HSv4oTUwhLT/X1WLFY0ZX5XEnCGluLfz0JxcQgHn
utRz8F3xaj5clbm5xjfxiYX9RPjf+YyHqNuPWfj5tC4gS5dzFg5naVTczHqsMkmqRAhRFxFpnxZ6
FiM6HiG5/OhhLOXwA5dggTnBuqLovxxWuw01Mxa/TC7bpjrJ5m/SyLkr9lC5vhQ3T6i8f8FR58Rz
wjLXs3IQBpoJ+zaEC5xzBOZ7y7SDzqVj9Co92RUB7omI6iv+MV2GIG/JJJN1hkc7FQQO9g2p/FXS
aWJw8wOqWlA2e+3pNk/EUR3ljmVbdsOVPb8I+3vs1BhFpow/rjFo36nqhgmDUat/zlODxZhgsPiA
6g0G0oG72Wvck71rrvhV6oD0Pa0FX9AOSJwKh3fNo1edGTRKTwmQE97Zj1twrnbRfWxcUl5r1sfZ
W3OqEPwq180deWGYUd2UcW9Y/fDQ0leXZEV9Eo5VC9DsE275UP4BMx56Hls/3lrTtvruNBVT6jW6
gu8CnWggy2lCgOriFHz8ToD2Jj4YuRLiFwkWPMqV/+fjIqEpZBzNHnDUMjwL9+XWg439qCEkGlpA
ISGVTGVQERZ7ytdUNBshF+OJwGptmsqXicJdzP/f8C/bVLIMG7k/wTpeSj9SdbyggXdeR3YveeTM
NbGjPPp0N1jzUY6PR75LsBYnOeRbPEyEPOs1oE5NDpEoTqa8+Jn/6sm1G4BsAa5D0cMvcST8BCIA
f/+pQupHCPmGgrmgKVMW9dDkz1PdFdroduFEO1kU4eWuzRocSQWojzYxM57/vnVI6esl9KTjpl/u
XAebNYDyE7xifK2T4PttHNAIGxHo6W+IInK9YmtP37pQ3YstD2GU13S/v2f4VcK0ae2UWJGcRSob
2V9Yp9bLb9FStGVZYY6OFlvpFZKaUditdOXLow/X9UECNMAadPDE6bCjuAHJaS1PDtNllqKzOiyH
NlmWCwaJGQEjN4SejABwIKIr4/tv5Mx3b26azpl1AZQ+fCWf6WOfy9BILuMSKw+OVBUvsg8oXFux
KIch2nhiLj21VY4gOnt9cx89lyixglQl9b09+Lo49KXAJ92XzZGN3yl99APo1vrlyyThpIKNWaNg
2UoYC7SiVKFz1+K+mOw5Pj7lTGPzaLSh1RN3YICasa+Cn9CbtvW104HNFRP1jqD1Yo0Qwl1os2mh
SrdUX5OJjc3bVDUPQbqUegybadLKxpGq+edX8cdwj+Xxf8vQIPInPunKvTaHKfyrG9Vak94hrKP5
V/0IlsewdJci5OpSpkZq8fzPuJDQ45ovL3+JOqqb/CjayomepZq15FU2LiDeI1s5pMgu2+1cVaKu
SRIjMC7XMPSmDaVsAIVwaOTWBqit/TIKGbf6A/TilE86VJB36BJDx57jp+7LzsDuwo8uZBZUoaMe
/Fmo3M5RxQsdkzJnpMBFKEHF419U7Hfw6kwUN2mN3A0htJFjU1wnHGBHbN3vrPiDfyFLm7ke4Ibt
Q1ClsnnSP4Wi2gbACP64r6prfcWmL3c9FVYb36JbAzXjFfJ5maW0cx6Tvg9nqOmq7ts90MBeixga
8JYoJAbRo+QehCnF0oZSyUjnwoGcGvgZqmLnWQNrL10jAsP9gy7HKCxNmWWFC8UFPEbF3KmJbZFk
Usj0Jh4iPelvLmYnqnbmonsMq1oYrVmsCdPSoSBJh5vtYqhGHiFAef/v18eUCaqncmubdCBWbLoV
RmqPvBbPEcEs+vzPOg0tVpa+3fKdCwqKyxHPzZ7zA9Eer5tw2+cVaWGzn8c/daofS9bEQEBMXgRQ
ByU2M+BGuWudnI4VivWUfOQlAoCgZcqbMkpnd2ZetCfkOGZ5Gu4W17Slt7CW4U9cJ9MN93z4EG+w
ErFBI8FPYcgwy83C0YODrZ2czr5qfHLixOEx7H2cP08sfMTyvhbzz9eVEYfQJrRom7kPOhrYBiGC
SEOyLWXRMRBXEvC/AZJdlT96yF/9bYMX5pA6SRAduXXQ8H5t0kBo+UvGVuoprIXEqVqTkVDJwSZ9
nP9+mH4ZeQWjNzEr4okJwFrlKGwCLXBoCelb4f4Sbv5H2zP7CGB1TfJ80zlRBwAa8GQB5aMy2aVl
ywvCiYMwauP47ssZTca+BYEY+Ec2YPna0Ef7agNtesBTL5eeeEgicIomhvClO687twO582pciV9m
Bgp6KBg8JR1RcWaas8L6Gzd+5kSKthMSUAVhUj9vcVnzn6IIR++MfB1k/6TmaJMicfemh03vnPb7
5Q3FnrHhZpA8LtimTIgqi/khNVKJaITB2UAWh2JmxzvysWTmbtHV9u/c9oAyHuKCZnyNJUvOFw7v
HGpz4ZorlNMEw7OoGLhg83QeNsLV3LojHwm+9AhMemI7UJYhwQbv5ArFbYpWpsEwMUMU5850akW0
nWDwQkK2XDNO1AL9aG7kL/3uq0vZZS8psHNSv4/bqHgJW9OyGueaBfgyCnj2Xio2rMM3gQ4xn6TI
ZgOSJkq+Rq4w+l5GLIPwDoU0VzPMdJb3Q93yd3GLMvOMD6jbWolQKS0ZTsGtuYUy+ADUzqk98WzS
nbHYIxhatu6OVmuZ26ZOwJ9L9943k9RTfGnKFZbAvAZ5LxhbRQzJYymoD7va9gS59kfdY1dZpEo4
lMbSEHmpnW6a/dk3UHs3CVCt4uSRN1VmLGEMXf2YWGMmHPCWwybXESEZf1/HMsdMtnMBwOeSjgVT
EYV+wCa0bYwz752scXKc5luGk45qs9z2gqd6qaTMwKM5yWwfY6IkmWeWD/GS/6cp8DXcdi4t3Xeu
Gbc/pT2EbvW5wGEVQLrHjjhsM6ZIhEA8UDahccNLMOAi2NWhNTc26A5w4i1TqyZtkR28zVXzwzF0
4N95IP+ivVu4WB0cLHAp1a5WJKbpbyTGMDFY8o3wWNWrz0rfLKwFPDn9d5aHtWhy5MXiuhVh91k2
CBEHPVUemYA8LLCPqdAhJwS41OqfPlLEtp5zlZVLhQZs2g6paGO+N+cMi4luPeFjA2/seZMRp6DY
sD62k/FBILm2BBTuY63vZ+Q6DOhgIKieeEfW58wOyua8+6vy3OJTmuMGhlCcnnkc9s8u9Lb7v+WH
8hO62VCGQ6FhijryPESkF941rasRrmdRBxGQJ700+NHeAhonWAy4z735NW/Eh/cXrdkQ7QmnZ/6p
9x4L/ufCHO13UFosq4W7zy0mSxkq22savHW8/X/tK//8nXl74heCF4atrBg8i/XJdt4ieSdfjLR2
cfQQOq+xF3DI7nnS6/2NqFkABhwR+BZQLgCvM5hKGOVfIVcMRA+Beb3MRLSdVq9JYb+wW3fykIZe
xmAF+6iPNY2q17OUSwhia3JXN6MTovnhC2T74Yl/oqWXnkEaqWL5wAMznrCdwlWn6+6xpQu8yEWq
WZG0BqHTwXmJToYupB5feV0Q+HecsNysyUQ0RFpdE6jIJnxQvKQItds5BmHm5a3vLvlwv6PmC+qj
ksWjiF6Iy0Vl0dcYkhbRAyfMz3O9MXKyleKZ9+BxEn6GT7vmWXFyMOIbPZc5umIRbJMhomO5XiTu
vonL5O5p7KYCLOAsD1bsiclku2rIFkz7if5TqfqMm2RE+qx/f4V+ckNxgBiqsJLtCNs16YhLhVu+
yWqTO0PmJiTa6gXmIeqRIoVwBOQjgnrkQkHiPFZekQiY8UbXd31Yvo9dBCaGn4uJdA99MAWG6Yih
0UejLhL5kn9dIzkIGHsAZe16jApukQ/7+NQUdwqC4AgD4Oz5xr/Mk2d9K4Qumr2Ujqv5/SYQ43Mm
z6da4jHwvpDXdm63d8gkVVtWeEnVdu3ojzzJxnTnDAsP0wN08pxB2YIw3A6zGCgJTRow17L0tof7
moZx6j/BvwmHFGhvYfU0oZ9nLyyU5QGob3f2dEUTZUCz6PieC/IA+oO1FFqSlhUrgqOCVhn5PB6V
BCNNSk8Ejiw62gRVMGViJiPihXarUKHawO9pHMKddALAOhXPYZkVx01FutRO0Zmo3w+lN5xlYSz+
r1lj1XyRepv+vv45z2Rn8q11tgvht44ZYi6cavTnlJkhbjl2p/Z0vVTLFk3Ch7MiyPmi7jeFQC22
OjaZEPhnmz/eKc6Q1dbIugjSBfyBdA/r/1QU3dT+0e8ahPhLjATnATDTSYx0WeRpLgRLEr1xPmNY
2xRTFwAqyb4rIgT0HCsS0f+K4VVSHexCieafpe78O5rrU1hxl5f4P8tpbMiokVfUVbGzzfrvXVDu
nPqy35FhkTtWO73/eFSxBXZTvQMcFb2ol0tOjSgWLsLwCqr4lvQL9k8qaCh8jEWFpOwPKuMVFc6H
lXnr2OEoTgJTX1qQZVRbBzgoZVAOrxBTf4/oNzsCVjf55pc+S55I/7WN8s28mecXnCStVAbsjsjN
ZTTAoHW/YdQT9VezE8bNo2o/Dgh6AQMJOIIXPBcI6Ijob1lZsJCkJHwHh1K6+tfymbjGXjcD/xJd
iIOfM9rkdiJNjqaWxhYMJYuPu7W11nwYCh4VQFBnbiYYsnpB5Ve6pd3VgHWdM031/muVG/OVJFlv
Ljxq1lBriTnHWEF7doaCHdbuW0wQx2edq1Lo2mQCwBybq3ITUfrjBBZlrRWnI13xuAQmZk4J7gQd
L3L6ul2bC8G2FP7F/T+B/VO20H48cU10oFQp9Le5r7E1QovPSLHzvO3a2k0oH3D8pAMSSJCYyWix
MZwWc7r8TTqjC9J4tAiQurWfIHvKP7VZgTvrWJDdarGmBhrYZUTP0RWnWJQcR4iPJ6cnza81YcPo
yPcZuhTB3iPxvlFgNjDbmnZNOWh8LmiyjKtqnXKNqKx2L3BiG8KXTTtCqjraW67gCxTn6uk+Sk90
lgFf8/+cvSIWt1o80BYSQKpboFAh0evAED+un8XH9L90BjP4mbLnZuyuxyhKdrUPeZhTtErySbdF
lHjibherq0olCHfjdJTl/oeJjw74fcYGxhDY+Z6NEOIszxEe1y7QDbVpalUUgFQSImCvtIoeuH/b
utxJa0PJhv/IhTe+6lALXm5fwz7hPvi8jqF7lZju+WAeGF9zBbSejSA1AN1kqjWDaLd1NNuxfQEE
2R0qVVogDi0ifqeUtcD0H+HQxkM15GWI66SNkgKJGYhqZxOvH7RxgZVgyEZcMrpnyo6G3NIctRM7
zvu7m3ZilLjKOJq3fdEtudjvCk872AP2UO9sPm4NaBtL/UXIdIQK3i4ls/20vI/1N4BFaLdL1IHU
d8RP54dBnVHyVUoSnXfMadvyztLlGYxyDHt3S5lUmP1ZxVrXpRetImQ3fZ9zc6AG7yvpNRs2NSdQ
uVMyUCk4nuNgDwlFeLnfzUKSEFaK1vuqBs8J1Cg7iLb+jUwdgrBAwLsUH1S2FGy6VsVDZvpRFtYV
jBxoT6TuEMGIwWanlnsNBeClWeXHnSgQvJyOCZKssWsYbinnP1XiKMJ0C7BjxtMO56xB9TNaYEFJ
bME0e0s8D5yR/CpawM3KQxvmwstE64x5385aNyXDHqbWOJZmmT3XvXpX1Vnpn97eAjDdVUsTwkAO
nAcWJx5v/oR7EIQtdXAAXuHD80Rw3yYfjuQjGIfmg7QuBWe0OQOrc+WtLBaZLYBsOpayAMaHvo/W
UueyS9EHN8OlYvOpQVst+WDVlQYKKgkEP9sgR52ZIJHQW+9owvNWvv1h7eV8yWcQfRWHsHUPl5Pc
UWU7eqaii6DyTP+5CazbofP33A9mKWQYdvJ2cTKjefV6Ak4smogYrAb/WabzfoaR4ggvMhTcQV9s
PvcZPpL/gokjK0WKOj9S9JEiX66hmFXZvBxmuAB6RYyxezvO5W++XpyWnT89QjwEKR5Q24qB4hq6
V868EJyh50ZUcfRQufZavWW2UOvpLtYJL8C0MSf9t7vEL86ldlUc9p95dQDQ7/iIyLeItL6iW2/F
tW3P4phbWuocnxhKg9IrgTNX97+mUaEDN34nhM/xTU1aJnXoYJiSneuPxic0uHIt6j6XuYqOLWtt
Vvv85qZIWpudlZWBd+AGy5zPxK/4d3s2JIOdZk4qBA0lPr8DKdCzh8i0LCHhjEAUUWtlbLm/t6Tt
Afi+Htevbqfgf7uvLyuiaFkSu/5zvrEFN1XUtlMccwf0pUshwu3oPBRTGkmOfpe8mdnkmrzlHfYD
nEqKRh2EWEwXzw6UXRYosVbP7XdSIreSxDl85wbGx6OB1w8sz1bIi6pCeYcN0hv4eFsXDN46bN1l
lCaIkfBhyMLGM4+Xg96XuA+3e1C9CeEj0066Ty4sLB35ubuzBctNn1DWJKOskXyf+22ELk3+VSdq
hcdSxWcKbrWYYra2TNiQrtcYtWn82xlt5g0AlMxFkvsVqfMvfVjtnmTstgt+oxAgjDd5gau31kwF
rFGZq3I6G8jvnWx5DiXYJQMAtuoIJ350krkmWOkcv+1/foJPTVXZE7QrJkJKgMz98aRs0C4Uuf9/
FrKKMLuBbI4etdk5DEImrgDXod1NwqCw4bonLKLfckWXKi8CFgX1eCPTmRdofYAoVn8MddWM92Q3
ZJ9FK291NURbUIgato7ZgYNDdb3sxHAJfrqvoCoRl5oBH0ZAbPQuvKJ0qXgYN/Mm0Uk5rIW+QJMM
BgPDvz7jCTH3TJgb1DZokklFDCoeNbdH3RqLKfua2h5uJkqTsRLMqD/jr2ZXssBDy3m3qdaLajOd
5JRiXqHyikz88a7sU1rXvR+QQEnRB58rB+yQlBa7QElUuZt7grkQm+mJVgP4LOmGokJ5JZ+T/WyL
`pragma protect end_protected
