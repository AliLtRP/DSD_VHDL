// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ROd6ssYCOIj2b4st110cMCyZlM4gjBI7adpeB7cefx5go/BjTmipjzHCaPfpREEt
WDWhIBCaJlpHjWtnpwcDS+4MKR9gUhh4xZr1YKlDoqpRz0kW6mkK+6hGGhm5KAoG
waJ2qvYXEkhP04sZOardl6Ya8dIHtnMMi8FMo6hRNqE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
aDDxPScOkAWiRapN5QxabpY6746fFvCZyJ64Wag+SxB8u9VUfVeNZb/7PPRp4iwB
TIcEyQA6LsWLazb6d++U7/WFJYHa0dkM5fBnKzC1jGTmGLws6ArGU+6SMxynkWJ3
F+JiuFXHAOecJEpNKjwOBVLpmDyFM381HMrh34nwzq2meI5I1ypUcRYpAtsEe/kO
v/l4DiYbkWQqW7sBvDf8R1Zmy6xvYmvhTgY0ZMzGyx3KGt45xEPydapqAwYvchGQ
0x9q5wboYolzaqNkfVn5ncllTzOkchNct4ZWKlhl8rJtBt4S9QGiQXXK2pg5Mk6T
GAmFYHKfZwt6JaD3sPIDco29Wq7Pj6jSA7u2QL6luCUnK/vXHry5uaKa5DzQJdF1
dUgX/JijqLtwOhw8DYDQVG5Qrt5kPoDLCFg1hLcVJBVIvBEg1vbaoMYzM6P1tbTh
FcvCa81PRHOTAYKaoNHw+SmFfxErQAblSKECD5u6INUXPj+fD5ROD5X3olcPU49/
QTn5QyfJK5kQKIMRTVdxfNoJIbKlNnSqiMLFjtcCT6bmdu46jdeLY/0Hepb5Nw41
z/G4VAOzf00lWHp0/sM+0lNKSLilSu/jm4TFPglg6B0aSJOoZGxqan+MGxe5PGfB
ia6+VqjrIxJN7T1WCa4jmc9oMO8Fm5tzFnZzc4jvtCwzUq/EkqSi0GqdEdIqC+GT
o46mJJ02V4c02lRxE55mIhk8gx+mxdiXSLm1E8HS65hx88VQiHm5+A6FuuRN9NDw
NbhZNT+17qI2g6Z9Ydac0xZLqjwqYoW27h0M3surheVPG6y4hdDdP51OL/2n2XRQ
M97iQDZYRnaZmavVtKxBFrAQIczCQ2EDQX+GzYxbccTiB/amxmfyPOuX5p/lBX54
9SwhtUutHdmlWilw/SNDQnATBlVlt+pmW+TrbPK0EZTDXTL2DEUKgB6vhWL4J+/2
npodY8Bnb6niWFWXvADOVWd8TL5DpBgToLrdrCYUc2nJZ2RLfWARRxxPFKBk0nn0
4s9N06Z+eOHAFfP6GiqqKG06a3Oq1Sm/deqcPrk1DU6nigjgzU4gIcKxky4Lop/e
lZ7YENpj+Umxr5sxCxRQJKovQTsPk9mgyRSYBDQZMnc78vN4f10KvOAIOHh2hvxs
Ia0d/pVuxZJiTtgsJX399SQ0kbREcc362xpQ/ehvHiRndJ3D00rYLs96nEsVNNzQ
i8jq5bTVB0dsLvffwuJ0nL35dyXUuIlbtDjJDJ/19pVJg9USa8jCkY3eGvi5m4AS
cJnMzNT+dHTYCldBfBymZdJ1y+tDvgmRmn62VApmHjLyIqovIqSdqD+gw9p9+kMf
KtO43S3qv4St8/Dqa7ri6Lpg5XDWIsLi2YP958Ox45wyKCfbStD+azbSa2KnOWHt
Jsq2T/tZ5xX5N1jp2hkwgz6PHJHjwTMvMN5RYagJhsX2r7zMDo8sT0WOy/F9TWj+
5fPp0IjFbFsCiJJqLx9sLU7otE+lpllPAJGYOiRdqxonFEHN+ExqRRoevHsC8Lhi
n6QnxhVVwMyrYZ4d8mB1Et3OufGbDIrlVD+qWR2ci/Yl4tQ/psvPdnEtyKYoi6Tj
ZtQBtOT5eXsOCtqZyWtrAu0pQ2paVK/RqsutyfkbXzKP5Dn76mG+nLvCpO1Zhol1
4HSeGT+Zia2hCaw0NR7ClCB3xxBtHO8EYZmDK4bVKK1Pgso8FbWnbONBmJFrJU37
adFwA3M9/006d1ZZxRPYuBCof9UUExl78CDt9sW7c4qzmxNAHs6m75Y4OuA1HG2H
5Ohh7g4wP5ZLXtDYUVuoth8JD9QREecuLYbJm+l/nWKYOeUW0Xa3d69OQM1UInUL
7Kg99e/cSpUAJUdouS0oih+VzJaQQXlg0U+FubW3aSRmdGWJqK5jsDGz4ohZaclN
I5JyEpli7lKhjx0XjxAFeHJQC9Q5ELJSzGYSGUzpMNpKsUuTZbvVZ7vqcD+jXfoR
lDb/ZWEN4BekVYYTKbQPuPRGOew0tSxBK0R0HxlelccUX+i8xUBazjuAqNYIdT9j
HopcsWnN9wL84aGzf5CfzU6uvfLo1JPP4C2yG4oz8RAwj2TTsvkfUScEy8CiPYBW
85EYqcQMcPic5oOjUjl80Afadx6hBWiRMsXRdBshgKOaoz2h8LF6TKgq9FVY647M
u2Fr1vsWvn76AA2blhpXTxLOmBaHW4+XHK5axvrF4yZy6qhpNfKl5m90cPDXZB/P
VR+hCpJ3jsHtgUhdxq9hwc2bXjJYYC9E8yoLvJoTo5dzQqs3qwqyxBRaQHS808Lp
1V9jcNSjKwRYarx7OPJ4o9W/TIyeyPboYjAjhQYZ3YKxD3d4lSoqCzF6EZpe7Hi+
AW6qsvLFEtYFrT30u4V5yHk59DYHBaNdKmMdUWsfXoEonwDALxvnir47HThjv+yl
q6Tw+kZcq2PiY5lt1IFhKcu01JeeT7d49OcN5NqgDMT3aR/xg5JRtedZszCCxiOG
3vVgbvCB9ZKpJkUQQ9h9SGIQx60kFN0WG9T/ixIfzSVm5t+NecBsv+fQtKTNksRi
rAdXmhf/nWoL5iCQ4qwIF3c1q+1tDCJz3UmjYO6cflyju9fOz6uPKF4jOnNt/KF/
SkI6itTrwXgmr9wXeso46/NEBd0gSmqaetq76RDU8OHfYqdwADrvl8vbGI0kEoLH
R7V1SwO4DjGv5+4rYs3mi4chyZjRJ+kUdG1EbD8oAXzhuEAls+6IUqhWgxuBCNqL
ke4shWkwYITwAxjA135fTQW8LXvrh1yZ2aHpVD6y9VPPDEk6EUdEdeqQRUfeNB8b
AJBjGAlku0ARyLBILEyIR/0m9btRS8aj3/oFEXuJtATKxBwM+ltMC3IB6Jv3O5Dj
nu67PFVRk0Rmsyy5jXsxDMFeMOPMRN8L/Zqlq6h31Gv8mV3Da7gPXZyo1/ibfJls
Ba2zVJi8+M3lrEtVAenUVBmH0i8StNZz7Yu654eqK2Cz2rbT0ithx46o8ThiVEba
/cJdUeyLm1V4GVM+xJlUkF/guyo0qJ7dXcZ82j0W1SnN4LkVPqr8i8jxyVRRMHQB
8R1ytFdEBa0tZ3mdqRzAh5NHtVRNoFlnFbykH+j2k7gMHPlHV1+uwU6DERCcoV9d
TrbeuwSn67tlb4dIYOYjwPLyjWJuEA+PIrvZDcyVmNuOKwPeFXIimxh37zWF8yS9
PJlZ2v0Fds/oL/QD+rpVJYrscWGy/ext17oiOxRQxyRzyqIOkpkk1Z0vxRO5oxhX
1qGbLo181ThfPfDt+fl4SvRPlmZgkCEPMCI8TlREOg32UJyQaHVtBGGxCP5T8Odd
dbu4du2H3rOYc264Pc39fUUo4WCeCruKJYkGYyXnelIi/T7o/Km2fPL/ca/XQkHG
IFmfWa2SWMNazCXPgDDHlXH7b88CNAxUI9Mb7VAD1XtgC2ou6ahrJaOLEy2NeUrk
wH06v+chlWr9ygw5fZXPhHZ6hgyDyuSfbM+voZZ1/bjM2DdpYXyiSVoArsMq1ozw
qL1aJ6VOEiAdi8yKtPfJkxoOvs8rQbKXF/bkEM/YW9rfYQYYIyO2yMMO484H/Dx5
4ofenl40MaDF3Aaax0I5AnFOTfjJ3oGR4GtW2Xcxinsujuks++rAPlJTvm5r6FXm
2GkKK/NAbsLA2Ci2PL7xzeS9kkrMiIoK0Iw0C81mED5r7OPbtaln3irGHLl+Ma0b
Sv6z97ggSIzIZotgZn337EE6Jy88si8tYnGdHfYvv4fRZm3tIuwbG93LkhAc7Kui
9IqCD+RpXAsXiYnizzL+A9NpDuvyw2dSu2+4DjIdie1YEzMtL1M2tyCgC13x00o8
ie+4TT8WRkvCIeYfNDA9yfLfIffsiPvvXpE7et44joH6xajBB1BW+5zIuEfEqMbz
kI6Cy0ictodTleopJbsPH7MAsckTGEuE9y0EM5nqCdXkfwO8XxfmuUjJ0EU39b9I
ZfWmNy+H3dAdOPPsjtTTss7CRs4rW+cmSIbJHjH+N+Pr3FeMjJq5wj+LRjNzdcFJ
wEO3ycB3lre5YKvWsV7BXKMvMKe8hIi97I7vBcOWu8ISgO8t2maj4WyyvHv8adk1
NgpkN5HjyeJ5o5wEBK+/Z/h4EjRJAwiuFeKUlsrdPtwm/S+2GUp9xEluw5iF1/NQ
IIHwzfsaVpuDv+SpBRMUT5JuykOCdU9ioU5kxJB3+iBkxRkjFOu51UUs5WpXKoLT
0yy0o6v2+REEmVBleyCvERzVzgtJ3GLz3O1N/gEaYYS3SUEobsnfRrMUiIETajTi
3HhAFqaMUmiKtMRElM7EhJnddRJ8+Cee7HogtFg63IWq7WgpTlU/nZxrL/e6CxpQ
Ng8glPWS4sS3302NlMzPfjiyS+//KAAYabM6TWaGcyBCHP969yH0P2d1lpr2ymFq
Me6ZHiIppctd0yWRBdKvfQLYUoKQnD+e8svNeL8Tq5Q+vKf8Y8SHnaIabKuGyPsw
oLVs/qs+FpYk5IHvq8g1FIm0G/a3CyaE3vu88LIlTwuQ7TlHh9gOCauquS1m2wba
jylolE00EC/Il9rF4dSYqb+Eay6+s2cfbISAxX/YBaDn6pgh448K3SfbnSLarRtP
nDkyRUolilxNUrGBDfHaxrmS6OS6aBogiBXvi+LYK+vhUDr5ceCAr+er5A+PuU3G
Yy66jKzYdBA9UDYagUH2rx0+/1RwGkp4cfGan9bK+8JbuSoRckzc+jUJ8wVuh+Hr
RoZr9Ms8gGgCM7/ZPGLKKkzi3/DOaFHFltrMn4BxBHhgnblzuJvSUac3jqTjFNZU
1Epu4C1PB79pIeCJxalE6HVMVBPli8kro0RyDOj/4HlXN8AuRBrDzh7AWut2BOmw
FNgaWt182DNNCWiSHXG3h0u5L4HpBY1xFoQLL7Zfb3aQh+x8WTDpP28ngGcNMmgf
zw5UlVdtv1SovEITgUuwvIC3PoyqmIb4zKKHspi2rB6i1KNyIXeZrDDUWZ8s7DMu
q+Ty0kNHzGT165ZVa5cHn7KjoXjk/3UKYFxMv10KHupYsNJyFPOioWgsYupSlujo
jslkAb9SzxmI3uvNZPyILfb0WrCZEsl+HgydQOTCFrXpZF9dwt9SJ8CxKF2SMlOB
aYjz0CmMpnT04ZsLRuhZJjy6cyhrcb2LWJxs/pMXeuxtanc1bILpgOQjeSuxWqMU
WZXIlbAMo0EQXx2KIMocX54NDoAGpFAnffaJNgtanevdt69ZmM4d11acBWzKpGQQ
oWgMqJXxW/s8hqpnJGlQxdSE+iljbUD+qxK7SqiBK6cXVXmFgNs6xYclntpDzmcz
/6Dxv0YdtZ7u3wgW7Xmz0M8bZ378z62Kxzq7/xGHtxMFI8xKKRxmRk5hm16ljI9l
Q3xRSw5ACFRJmCFoOPhyT8FuKYP05MRbv2gY36OG94ookAvS+wi13lblmDvbffwR
kLQBnEqUMOHrXzt7bhPPsuvUDSFV12zySTyrOLlikTTIH8py+mU4FEh959DFnlbL
LX8soThqfYPDJZZ1bF6XxK2pTVlkrZeZ7RadpdAHjjD4c9gYpOGr5e3vuS+hfha3
RcNGjFElvQ8ArAVaG9nAdYkmKNcKPVHAbIR8jIF0XPDCQHcsdVpSJc4KpfqVhE8G
cxGpoIIXysBwzBmNtYuWUu0ntolQ4E2Mlc0k7Atj4EYBHRFT5xd/Jp/thPOJMBM1
90v4s69dfF/ECNLGTXLp6iXuTgUyhfoErFWNzaAt+iCukUJ84uougram9rotlayP
5kwOi68t+wzCf+axm51pQfkNKArIVBt1oEjMLFKK33xyJUdJD04d+TYqTpahGGHA
0wvga+ZhaEfYhJIFtUqGD/TuWjms6+4MqC5Y0FmOFkmDZwDdPnKMnfJ7sOg7TLnA
eYEtlNbIwyKTp86+anlrrmzdrcVT4wel/i4P0hmkp+w1CCseCZshzYZVDjwl+/C0
X/ucb5SZVWuOZtmgYLs7Ap7SY/QlXciZwdpcK4CWuMknyVaoQg20rEMaXI8cfKde
fc/+7x8qiJZ74vsr7Is44WNbnYf+w3sOnMnlOpQHukXM0BAR7G3cAkYCZcEhGJh6
C5UUw6VmvTzYB7WyuH0X4g9wyYxH1MlYfPVVyIbKx2ZVtj67tg5/o2n2AFLXxMPG
JmaOrt6iIs7T3xNeKUfJvrfjGyU4GSiil32Z1S7SPo5EuPpJPkmUOyE1lynZOItA
rBNeUr6kq+mzrhnELOnb0Mf2N7O7slbR1iLfc1YywuHKkC5LjvG4zxmncRymbYxZ
OhH+vR2duOjO9C//Ni0BRfKhvgVoUfLU6KckUaGa/KYz+QVK2Acy6cCdk5heWyso
+s5xrH3SCWAHRfv5P1E1xHjTHbIKneGzBWn+xzRt0HhnFyouzfAI+roP8Xf5XbXH
3bo0gGij1MwiXmuGCV72N4boiUUF+Y2xCbUAf57/0DKbc7jRNSB1/YdGHNkNbZME
C1jRmGFLpTnEsOVXptQEa/PbEb4mL5VKF2Q6ic+Jr27OqA2le0+XK5vqf/q6klYt
vDTtxOaQjcBNxp73Fb9783jR2PVWUVLvGOvRN0+NMf9gpvNPJkOhzb06Q3WxIDTo
slVuXOK1psgVC/fjuqKA4ktm6NSwLyLbRqJiMcO7EP35icMMUpHmx39JstQ/3EMQ
NDWdob+yOk431hzLgsVD3OAu2gmy0oyEzaz9ncmMfIUcEMMy83v4BhZmKi1lmcTO
0Jf4gOz0UkEtxIeXBlrF03B1TIFs9ycpzqxg64RllvOHVYdpCnH/PShzCze2pHtF
zLvWGhw8C28SYG8Kp38d1DmTQUNS3dJH/HdENg0X1DsE1OtxxPqh5NaOhfMqBJkp
hQBVSr81wn5CKvCX6N7mUI7vlaVZewQpw9JtVK+EjXGFVap8Fu/f0agwwsJBGxNx
1QKnNg7P7r7f7O0Q0OHZHx6mv7//bJbuECkMvDSzyofcbZhz7IMDEF8OV+bbEWds
mkJ6yAKSgZBVgUKGprXvx+Kt5sySyZsv0eCuvjS2g9TwF0tTriAtAO0Lmt/N1EtG
rKvD+ikgNGrHu/W9xkJDniucEThVFiSpoB3lleihUXgZXmZW1rieGVFj/KHqMc1A
lsjszzHr4CjX81nqOl16AU4Hf9Ow1w/x0mkAnX+t+pzNyAm7fEwhYR/iPXReAst9
0tAoipuX3VRSIDIa4cCPgTRGQ6qT++/F1Trys4ExgzJ0atMOZ2LP+FMisK/8U8f8
nYJJEY9HqjVvIblg47FXYOncW0EOAnIoSM3S94oX4IEXX2zbzFknS/KAk/sbJoUZ
owzAOjWUH7iENS6cIMUmLzsKrcpc+fo/3P5ONSjT84RkNnwispVYSmBWmto7LYqF
0nY5sBMTokxbBEqSkjWbA93ydIvTIF3GmYm2jIWb9ENU3p1qTqn6Q7Cjp8G88oT4
DELG0V1YIprBCiTaVIdT4cUdSD3B2sd4Hk5BTkaA7jk8sBRsn2C03ziL47NukWRQ
+dqiBv8o79NwiOefiplBePNSppCD85EBGTVCLtxa5eIs0QfFY5fV3z+TaFbb7cEF
3gYxOqMdUNrIoh+45xLvMJGokhcHqnMysM353JumTYU=
`pragma protect end_protected
