// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W9VjF8BoTsFqRr8B87U4Pzsak46rYaMgjOEI3RDk+kU0ZV9/6MVq0GORojJKywtb
G/DtXNvoeziai8s+wPPigYf8f2ZbhG3sBNVoAqRyWk68S7SunRYX3YZsY2kOu1pf
nBSlYfnG3O+4PQPJ3lCzulWl/2+jvvt5i5nlcgEwV7Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9424)
NGEvqdgs7FOyHnEPuR5eKAe9T9e88AER4Ii3ETk3BBaZJmhN2beUCY9MRciJoOjB
DqE41yEh/eteUS8YEq4iBZxe6FWCi5sO48lH7Jf4cE9bmOzVSML12wKXLcVuRSxA
PL8163hkwLGsbmFXycd05dMkfZWKihMll+XpvFHzgUmGrznRQdSX5o5ZAPQUV54t
IAJCweX3zonJk4tEUvwLBN4c0kq353pgm5enarg2dHpcS0KflRj10hm++zRtvIuy
vHp+td7mlYnMWPahE9JZ60/ekjQY+8yUdtJROj7yh11E/M7UowYX7oK2KX3Rb/NH
si2WAfG0+P+GBn4AdHj5GNc1hc9D9t1DRhy5sr7sMxQljbzA6HdXN03Icf4qPBaA
rRakJYR10qttraybRugy9ZvIRw0cT7uIcfZn/7z3EdKcGDjXB8BrGw88FLc4PBcl
LxSNl6ratnHyPYz7/vVMnWeXC20wzVb2GqGhuQBnEt8yI2Yx3Xb/InBZofC0VLdS
NN+tPfxVtsMPBBDKS9z9oBK5s+dYRgwAdkJsJJlm5J28ZjuIl9fX7WdhRJbR4yp0
TeP+LW7PRhazMKeIxXWfuhTMk/gXhpCByF6Riz3jyNZOPRhIls+EfCqv5P4p4Gyw
JADyXDZa5i2DXeZ31d1FcV1nsiAuEBtrqQa7voUTHYJuw/1Awefy2XzyvypOSuBv
DeiyxsjNqNieazu4Ipo89FmvNfMFwH5eEPsjq1k8L4iW0cMeMBdZuBlwFANCngOb
bWBN/3bNXb6jkb0rJWxYNi4JjKUQVnPCIIgc8pcERYp7AeOwNQoqFqzHX6ccxet1
fx2Wm7KxDmKBmhFYrAcFT26/lFWqZki87wsprX9WzETSBfgXjxkbyCnyWVEbzcs9
k9p0LY5I0Rl5YgiKhJXDQR57GoC7tP7ftFLSvSk8Tp+SpIQcXapjdfKyfRZgL6uS
Qj4rExCocB4Xdg4pufeJF1o9TwvJwl5IT32WK5AVqYRSMTkdzX1jIxKBAtzLtt3O
GSQGNV7QI+BHQHAqLHBJsx0DLYtCUpe1ARAVXzwzMCaNmkopu5kAkwlgXbKlBqNa
XdJZcJ/qm+6YhPZQZDZYgCe7bgE0T0cXkiC3YBIYZAE+DWshqlugoIoQVfv08Qzw
t4H1Wrt5eCWtal1BOmTVtwRB5IxkQX0kHFbKPYQL3V7thuJpJoMiCrUK2AFrkc/7
HgmjDK4rrU5UJkakcZMjU9Q8+98iwogMbC+d28qnor9mIkQq5GmNIT4gXd3eG7dp
lYKZPlCm8cG3THxQzJnnPFYpi3sVbaGVCM38/rzPRVDdKI7kONgcNRLBDicH47In
wStLa/RCcM97vrBSo/sI4TyzLdGGDO0lXDG5s5Bt/bOLHbnMXGthCQhfIZC3bl+u
9QztByep6d3eKO0cFWCzaOOEVvCLjhmFpR5zq2ozl1KkENLAgj9LnXyB53v7YfTk
e4ANB6BxJ+P8rQTWUq/+I+7kPgcipD5m3XFBoydY53WfKR98qnsjbvTjuGquJ94e
jE8+6Xu20nSasjmiUwgPu1bodlA5nug71200Fj3m0tJ3f11+RWfN7Xd1iw4pmzgl
jbBKaKui6E9LWZBjDecvg4WJFdq376Mmeyihl/rmTCKkd++XZ0dWlDZwg9haKY2S
czpOswo/6DIzhaOvXNHinEaOwOcbCufdJGQQQLMB0m/7aa2XRSh42mVqd5BG67cD
yAehSi2U2p1HSi59Ajt3xsyjAfuRh/TQwGiHoGP6P0HFN7Q9op9S02iNNyVhkdZT
kjLJPNzKBlhcg/tvZkPOLIIDZMd5zJfnhmF4dDnLz3K31r/rvwbf0phXyxxYZvkc
aF4UxqUm0+AxAXrOi37fyBsuNkJULKcTHcaf0sDdW6xVAKKZA8ZrR2VrMvMAyvyN
PksEvKk6OxhnLOBy98j7Rkx4loe/I2Y9y1e5rLFJblLJQoQCHPSL7OrNHGA+oB/G
OyiSehQiHaEHKNdmBKteAK4WClfI6I8Jpr2zBU0zv4oaIYpzp5Tr52fb/SR0co2v
O20eO1G5Z4bGtWbP5k/piFrkPLfb92mEsQBRIejbMiXNx/btphXtIlHbHLKN2yaY
lpzhLiBpD8c+GloxerQHcaOHuNefOaVChNpon2XBPOFEWVElpQd7Vpv4lCLf6Ins
SG4Loi4z/87/JSB8jxrsZP3/A2gzXWoHfiUA2+uN7MyLV4ww34Owy0VAIs9jyy5j
phohipNvaYceR56S8YE/6h+4A9B4OzXfQOACMAbUI60FWSOMq5+yxLeJmyVSgIYZ
T//eL5NrHai60Z9db6KePp9oi1Sjon60RrhI0TmZzN8CmLEc/cqLBknhs02/uxmt
cMrFZYbNgKMhMikO0/S5YlQB4rrH3Y5ZmrD6MaKXHnUfLnGZZf+pMcwXLKpcxdUr
sishm68++TNLuwTziWzi3/TP//hBJlg1ipk/kWQFOu9/ksALiKqnaM5bloWL1297
S9i9OCN01KOYx9nN8XTiB72Akmu55kTDLFurh7Gk/Eq1awzaWiiY7+uKKi1w7fCp
P8zc9cbSrEUtdckjTDvxfa88jsByB0JrRK7LW+pDsi+S5p4KWByxIEeiXNCDiJ/4
PeXV13y2lYBVfYt+7tKLGcQjWAXwX5vu1gbsBQSEkx5Vj0y4AAQkqhzVkGaVqpFw
GYSMFXvAliUwjLkv5596TySEG1/Na5SuS6uPfn6T4cTxrnu3+Z6O//+Ya71CkGOs
UCPL82b0XWG4yUF2b+8+TGShqYzU/9OQpECliNlNncCUHGO0Q50A4zVkGSaEAfiF
iUqxNAn7huBn4ATBLmpRPlrgri817K8hbswHXx8ePWxyqnTURaI6JUJFcNgrgFQH
GINhGTsXlVz3dbKFMrScg8UMFmLmdeu8UxglUYuPP8dSoiBo6lvH7TfZNbjBmNx0
xemPDKYYmmma4r70S5NJR3Sdk0OeNRxUly/9H0Chmbx7MPQ8Z2d3CAFYMprppFdk
N8KIZeYJ12QjkSiPgMpzDSrdH1ZBWHg2p9yW27MW4QwByrD84UP9Y2w7sqeqhqUf
3z/UAnJRjzdcMRYIMT7LEbMDZounuKEcY0ga6/PcmM7XncTylstlhjjQOjpTW1Ni
QTVwjMMhpLUwsfU+XEHmiBk12UVnPYAvt4UZmN11EjkGRV9KpbRZhCEuAHiLAab1
jCjrK7TloK+V6pReAT4A5dVVwLCziHhE3bD/yeiJQTv+HCD3TEjd+3o2BJuGJNZd
DvJO9FduhxFCP2VxXWVNGLmnAODsNeQCH3RjuTas0o0ahqCoqKBiVuiMaGYK8Zaw
FhvODVLh9r7lgRNXjLxIpcvVpCQRqKecZjczGE+sWgQt3btgahIOoOcedPEl3XwZ
lQWabreLaql6wQMz62VJncYDV3oaGwgJ2fMMKNn4y7eQIQK1urBYlEkhxY15aL+o
TgzFDVI4ksA9BMf1hrixkGeujpSlE1ZLPrOjpbAsPokHoy3jpp/yXsgjII7j6Q5P
a7cWpVWAb5cvaDSOCYSJ7SP1XHgCV+qmQYSwbyvWePN3iy6ImuSoCFCh6URShP0c
eeJ1LV23gAAG6CiAFgh4hcb2IQJFTqkLjKWXQGAh635OP/wi7thzynG0v7zf020J
J/RS29P0oZ9D2SRqm/U1TquvHtFpZa7wJq0XjVgYx/XVDXBHinryIvx0wi28RE4e
wXlBJEPUpSFHpdksVaU9DmVYvJUOkpYrC/tEuum4pnPj5RIeByp7HjLo/uNeYPfA
tuTaga54kRjnXanyTbTXl+FbJODysw++jkZTRKVo5gj1oarpw9Pz1dHXrE/SJKlW
w+/xg+rKDGqWhCgWSE+UXLl+sq/iM3cQUHlqHOl2tGE9Q5d4u97R3tUmEr4qDK+l
de9+QGlCXYjooHh/1Jx44U+Ym2CXi+sPOu9VfL/zCog+Y9ER7rgVzOx5smBj8C2P
zVeNRnCxCWlauIQmQYkeLf9cRIz0FmRfMu17SGuSJN8KdTnBQWNlgxKRPZhy+rC4
XyfABc7bC7MdD0j45ZqnBuzj+oLoNJoRAFmK6DNZ2mTIEZngVORDXPCc+DyJf9GI
iVmtpURyS4N9rAZD+0eEUtSFLq/YPLNXbwkZTb99MjlIH+dAJUWdwkpb2CeV0NQa
5k+hPhTUGEPN3gPXPzyDutl7mud9LH/KcoZZGeQy7a15KA6zO7poR+9bXqAg9IRv
E3BxUHyAsBRd80JqljieW5ESnJ929Ek9iKgXt7uR8rT9n/i3kxoxuc3mVkleVpDG
eyZSZnXRSQWgVEQ7i9SrRyg4Sl2XhVj23Ye7xy45qKmdbzvLX7ld5iSa3HtJFdSa
/vEEqgsEQBkf5pLfBA1nBGlBiB7uOmab9Yz49+41SZhIP6RoK+CpHB5sCLWs6YYU
OALRCb7/U6HSgArYCeeEplfDHPsXIdCio2S+gjOMS1zIY40gUIET7IvEMntQC4/F
15Xab/t7O4SCv3fdbnZ/yrrD4+nYw/n4yiNm5g/r10jfUBzElNrC+EXBWVOBhBqn
Ak0fwl9H1KNVUdaoEdZ/YaLfEmmJNXd5R9e0EvlRJ/tb/uyACZKUIsftj7FdmR7+
Fi3LkkIe8Scos0Xwy2vN1D0Kl/08e6kIQkOx4GyZ7uBWJK+cwO5geZ0xe7epjc7j
WPk3avfyQMAO9bhNgcViCnt4nKLcj1VM3aXK82vwdLkVGcPg62CuoXV9VzPgGzFx
tmywczPBSHaZnmNdFpzGQtHtg8ctpJZaH6ag7XbMTzi+LDgipNMw/SoyrGPBQHlG
SIRa7vBvszyBCCnEqf4w4VRMqUmNU/zDkchil3t9Jq2pC6wYqc+FQ3aXLXoQOSaV
iNxlXUoZ4S8T7DCnJCrw2EKt9fikFVyHHJY7HJQeKuPGxJ3yehIJVIngldUmeLXe
TMV7pJ13ZXq5AqTqGYxetw86+5D1+lwO+4W3CMeM8eXpKtCJRcFOPxuNCg5QUOkM
W2OSBwkt9eoDiFoLRwrlQ7YFTYZublQ0qmffuNNp1mbS8sUHDnsoFK/WYSf7ghRF
tMkzKVlbbvoVrT2qyEKT7EJGycnFWv94NhaJAifOY521nscCetF3keGE67rKWNpC
3ahDh3cRPpdN0oeAwxdykd5ovzq958yEzMi+mLkkSDbbzEW7MrdjMqCXesP0o4v+
F78n5R8a3kvjGZnVpXuaNpOftLsBbabL23f9XsVsCIJbx8pLo/hUbLW2eH2XnzSI
TDT9+idjWU3KLB3mlMgEq+8E2C3E8REV1b0jvuAmKeANlEBVrtQTn7QwhYOWA/Vh
2y1XEUMleYbgPdpvM5KKmWjH/2YYWGhHRHUZ0tTTMfpDu7CGY6JiP+ZzJ1GAKM0X
fjZO9dP/JCRMNhrY5YNS5yUfi+cmy7ZMhWQjou5aa1lNUP7ZF5SR9czCpfOTZkI+
ECrnE4KZlwxjb9VOFThUMLHJwvnl3QBOzhRlTWP0QdYGSHg2aE38KstU2TRr0FpP
qzkpH+QF3KZcfgeJm5jj+QTih6FXbGdZ1fPR2t8Nasyr64VzQm+c0qhLpmZyP431
atqdOjXlpmk5AAM7vn8F0FEKTKgjEe6klXpt+i/e5UGbmB/gIk0MHOfIOZnpF0te
MZdBkR13QOYGkP/6KPyTHfI+2SWtNyNE5yGriQXkzXiikjD2YPHoURCTTRSLzxQM
ubwOj0rqMl3Ut6LbeheQJi7yqnvElkalPAQz2+lJQApRWmbChD8PpqC249viLQpr
oxn0GFwnP59Ou1r1PPRrKu5anV7tORKuYoOABru6QBp6f3qOGs8Qb9sGMDMQTvuC
GbAIh1pTMw4pyGkZg0vIhokyT5mwgvJ/yLpo5jocQ0X2WF9GhRxhb/I9G3Q4p/tr
4iBoXnWhj6NbnNjk17F5VdyU8DuMPAFlhEEAtfUVvAunv1QXYYeJaLiPIQv4I4De
hWmjQoBxd8nqXOvVAnjgiOzt9HyUv1QoXoL6LR1+MUwSBwEahZoU7AQX3Q5F5HYw
oRoqxkXE/IrPanz7TjTSTwba0ugzWo4moGIMuHZ86XZyCL9xJV4YAdvUjAkhqVEV
7ZtNpDc7b61pG9AHBJR9u0YATR9uUBqux/Sl5unazHLHSrXuFi69ScbOLqCmnb/m
p0TMJi8TM0+3qqQ5rH2y91nc0X56nSVjgsV2/XAIkEXHeUr3CHtc7SNJRoV9lDgf
FaR08QGKIrG6f5Z4k3K8y9rUNSLwo7DC1TZDLdFfdxxnCLrv8mUyPfN1Dek6s+aJ
dTSY8YF5OD2hZz6WvJS2MRgOQNYn5maH3O3R3sRRjuipbQ2J9QFY/dVmfj95txmj
O/DjsgO8LI6HIaHPPdlq/yRh9PGSn6ZRe0QL/0oB6IS0fXHkaBX9SsyjtO6V9awn
IRkOXzjLysdJFGiRfPROdgn84Jf0Ff01l0q9J3+/jEshw0mQoflBHw1ofGtHUGl9
INxPtqz9WC/FUjvfj6cc79tVQNNd900U3OBM/C2Ar9LVuv8GGYStZWXlDSlpwHdp
rstk897jdVDowIHE+INnS0ca6DLE5FOEjhlSixmOHrbKHCWfp0SqkCUMNS53SXoj
CBBpHeCa7oM0ujrXXWW1j/8Sxz4HNxExsfvC8M1pHMwWKlw6y2wG7AvB8C6y+c0c
SQZOeD9kUgPT24Oy/zHnmJaPcqyewwIl9Eb/SYaejMsMTXe+aokipeF8l6sJqQxH
6nfLSsFhe5j9b902vXvMEBZeXMCwqkg1138tXXtUSyY1sth80UJhPLQ03nYunNw1
YbVf3f5SuYxnF9IS7Osku0sdNfhvtW2OrVAGwtCyG9QIPP5Qd1KzS9Oa3YXBB/+o
6Y+GubIgEwIYQ/ZBcp0YhGCDtOZffkmjee7fvEQIJ2KClW0AqvEXl8C3+HTMml/x
kePs1VsYmgVaTBf85k+bRBWPgDIaBqjX0QmPKSLWO8KYkFdMEMpaE3bCIGQnlgOF
M8S3eXEejGnILb9yd2w31SHQEry8tTEnc/GX8AAbtnC3gxpqvktj3IiBa1ZUNcsc
z8iJLK/Vi5air8fEEYgc+VSiqpdDmuwhAIsNdIuoKhhj8jiZ/fkM8xxFoG70qq/9
P2/y96i7udDwlRjRLAW4bHQSXpsGPgrinr+zRgU4+BU26rgBDVD1CPkV3I02amPT
sF6aZnyyrIgZLwlMQ0CKZp1q6xp/Bri/JY9ZHlDidhg3UIdcGZL1j/+0jffB/Sau
LBXSo6E5NsYs7pGzEPbR5GrwZlwzguXp1geirILdF/eV1OhfM9azDsng53dcrhK8
irzxn+8jKAQGywbcNdG7h5OVpSfTqj0i5KhAZsFAKNhdhF4FEzr8Qw70xw7hq8c8
79pQK+lcwKENx6TW12nWUgEQwB3gcIVUvd5TB0gcfkMuLJnNsn7bkOWvKm60ltz2
KtOUUFjHjPehajJv1/2W9q8yXQLra3EZBJf7H/X3EV5fAbIO8pusPJdesWEH04lL
7WnuvBp+nmbsNYFOOi5iwQhcUwA67EschOBCe6UUavdorZ7VfLQA5FXs7VnMZsbV
IcpgY7UDZhS4HLK7gpdr1ZY7cI+nvg1fDN6VJVp3BwTfQQMPlig+ZPESkEm+LYPH
lt28ZfbPMIM+MrHYYwVBqmcADl8R01FaOJGqrVF5QIfYOuVQSTNrXEhljNt1pxj2
hR1DFB6bBTO5On84ZUscKpejLfThGXi1pBvYeFCHyCfNCqgYFRI5+gveVmn5BimK
vqA+7seuDv82JZG8z+jzGyZGTnfaY+mBKAc8BeYVMF/Nl7Km/YSKOEv4jka4N9Uk
ODKam3oSv+hM2Dt7X0LmYd8aWLw7GmXvPLdAmXRZI81iJpiVt+O9PjXXn7JFNTtx
44LrN1P0ZTJaK3dcRR4qbRh62JQbNxx7n8SPselSAluj5+H/iHapWwkPKSY2NVd9
802BHntof3x5ZcAWkO90XAzesvzapMZF3thHIQYB2O+s/8vtiDi1YbmRJF3UaM8N
xJY1JbDH2fU/Rg+PherXAocGPULLF4ZdZkgOPfjwgFW8RiQW9NF0Srm1fdtxkLtF
rrh4viYHRhwKlIy1CAt5b6V4ofeNiWfFEYWgeXR2EbhZBgwST5MQl2x4/t9sbYud
bwbIIFe7ktCxRDaGLmdrWFqTsKlacoBrYhl2cKNRq+ACafURcksMeYmnm1JTEAj+
2CExBYAKRLWE3C179SVyHok6eFeLtZDf9xcc+xPVWL+kZLMtziThnLJdSzQ3gQR0
L7QMiakYpS5EvMxfTrG2DqL0gu2nSiCtzj4s9gS3sfuOjMybg8orxVZVfpBoIXwm
3gsMu0KgnD/Rbjkca8Q5X7ZoXzpE1xuBbmCWYOA8UjdJSu40hYGqq4pBqTI6JG37
30dxDv1EiJCrlsvFmjMqE7sSrlnQAYbHaeeuX01q4N29tEmFg9q58Nfw1YFHRTXC
fJXjIerYa80mc2bxy3TBA47Fayur+93vGfhxRccehOkMQszSuwwhxOnPUp+fv/Qq
lg/96fGJ8Nm7pc9+HEDYT17reM5kOk0bv1QjaPHL9JGQKtelkk1xaFRtyMiiCYgf
hSM7QryT2Psu7wZ5GtTIPprItN5crRCM8GsFRtRbDr23kCzZPc3FByg0FI/zkiH1
kCZtvE9WZqUdvZRlcGV6+Ialwcnjzn9d1AaanBWvQxnuJWhXPfjWUHC6FyOn/Opz
qTR3YOshlpiyYpr1hJzDBa6pOE1Fez5z1CzpNOMmlO/HITlaSQzBx/nYOGGUYkmt
HxFUiEzk642MnpG1hDCK628O+zO8TKw9pnfamDpxys/GhRROIUtQBkUOltAEgNXp
n2vkuwxZp9puPoYqcecnXM2rbguA1RtfFPFXOPpAJcqluHRdox2WBoC6EqKyUVpq
L0jtkxmiuYwJAtkqNxKmRGdXNeM4EQUVRTZY+DvGloxoeqxJgbRCPebu0a0c/Bbb
fx1luifj92OIDGOen4WymEQwVcy6FBNBJjwywJq9shw7rLIIIeYL1c3KBMEQY8/h
XeyQ372wIAcXidz+kAzvfdxJr8VzLavbVaefe08/Vxq7dbFGVNENtgdezuJRpfwU
2s6J/hgZY566RPftXVQewqMFU6OZuxekH7vIJrPhO/wrAgNGkt3Z3o5Qgp+/NhVL
j0lrgSUdgwe/4+kLbu+XLwFqTGqtKLIRozoEPpNHFjWXJ9oASmjmxEoPPWAR6S5F
dyNHwjSxj7HemiwsIT3lX7xkvuj/pHrisPBGuvlv9PxebHe2aNB1lbcyzYw1ZyHr
sk6IHI1kFS8k0jJL9L8PQJX4vg4wkAZQHjgmj9oLwl50bn0xybP76Vp2bZe4YRvW
DiW9Rk67R4ZRijoHo2UfZVhw9SyhxROTGwVnvdMQ7V5KHmXTHtWzJKfKWu5UkbtS
lOqTs9pNW1vkKRgOlHjQNL8hjgIyd1tTa9O9oaYnlPE9CO98wyM9i3MKarQInygu
slJf+8LK3kVpmK6Tdhv3Dl0PRoxzIFmgTcjruKbwtX1cKrCkXL+3RutiGuhRlxOw
xWpwCoR7xXuhCrFAuiLKKgGNaVwbCKbMse8LgFtU0B3uvpxBmno+DFEPMkMpgh70
fx7xDN5x/iyuCvhYlxaOAxOZqcmp8Wagl6d9j1Q+riGd9ynIetuh1GNf6AgXNnE7
5wKvyER9MhDep1d1VbEC2NFtl00HGlRv60cDXFPjP6v+O6nU/QK5BGCvqEB0Crgc
qhjmYE+2dGN7xWlR6MAqrHXQ2gFqociuquD+5khmv5cqJlfrEmFuwVw/JzkFvYae
EZ5NNH2xKeZsUmLEBBYLnV3basBMgdBxQD6MYuZV/sFqMVL4vR9nuTNBA5yz3nqO
+9jwZ9J0YKHVF+8JbAySDuf7LXiNNQGXiGdlRq+Kv7b8qurRWyl+btMah/0BqAFd
BliQIb2ZvWwgGPFnzjjre5HlGFUWHo2pQLhFIg+BNY/kkSSTBbYSwF4FwnSH5dR8
u23/Y95JtkJSBMT9Pf/vmg6kBv26n0sm9l1TQb6NYtPOHmVgNo1FUi29Og3ArndZ
dQJvouRNBqe2ksh3HjBBqBkvuiAS+h7NftDI6nD/Vk0nIs81kMGxd7SIbdkSCSyl
MaqZ6vlqifjQImZWJOFv2Vz23NQH0HvhY0CGhDbQyqJHNfC7PcL/DdfCavxZZnE8
xgnPvQ953+qfZ+JxtEoRTogsZp7iryn0G8G3UQEel7pl7AQ0QIebuS5ccoXzR/Zx
57l2MpJBONW8tnmarWnf7WlbmCfadc8KjJG33DqtlfACKapBuB4BfUj/5i0zYuAW
LrRMT2oNn/H/rIXOjY9TmN9zlinCACfs/bGp7kYV3V1m7rv0lHTk+wVZ/y7NtSGb
tApTOH9lHxSauxmIHsiDEg/lyq+fOUnmGQaaOkoPKzwd55dY81z6yaVbrnlWUFBU
ShfqnxDVzUh97svCZtVfa7kW+JDvVpVJKLNw0IRJw2SoQKyiOEtcDivM/VcLr4Oj
vNtaxLCbVrxUfT9uvIO8yUE0hrMx73qoXBlF60UXgN55V6Nf0nVKC3FSAxDoz1u9
oc8M7fnfBXBM8R2uYJDwgLRs/LDwimkVTDgWHD8LjiWMXgJTRfFgbCaVqu9tHYqu
haVUYA6Cp9uLXDwtwnCO+1zTm4J3DE+gCyGeJKKNceSiEuFvlx/j0jySq1ibJj/L
33QS6/y2GJwb9la8lfGczCMyMhWTb5RIR1DfcP8pF9xSWIwHeOdX0GRzQAjaGH44
8Fgt9BAfwrmdaGVqvHiaAoRMk51SOJqGTj6C9QV8HopPjQAQL+lMYc1MFfvU0OYx
j6H4fqH5aTmx9QRWqOrHAObOqH0+iCqf/4p0t3BLQkLAySkiNy5v2+uubk2fG3NX
kJustMXnIEYn/g9Rs8NJdKHVU7L6CzhTtYbc59sXc1sOJbA/3PhA9EoSRZWxfbLk
PpJ6kpyhxA+OwPNXORv7p+nvtqwZK7xrusAlE3ft1ECD6S1CCFpJwNh/J8GnNSaT
4U8o3eeRCDsQaet4f6zKm1MkQupCbYF6/NzjwD1UrtOuxQaORByjjdBq7BTYPCt9
G0+07oiBCsl04Jeaj+oz6gXXAg1QBM8HO6ScBYT0eC+3/YIMltzWaH3drkYq9+kc
IfXUmqSMwLrAIyObT9RvySz+h+3XrPyfxMQkUSCtHLKKOado6kuIEi6l7YiTdZhq
slqFi0RtrRYhnX9aAR+01DfqQt9HvvczyCK1QWnWarfbB6l/PAsKCNZjYyiHwvAG
7wGXkTB3P4xAnZ0lKmpUad5x/nlfIm2Fam62wNMmrjeGSTz2oaG96ZbsLviH4wG2
bPlMfun2xOhXBR+9uwNt0oWT3I13PpGQXE3ucGRXGsQSHjlf9equkRDyj9Fmj33A
9SVTyBKoWRiavvgccVatVHEzCmhUBhMPQqTot/2Y/MPCIMTgvaCSem5C6WwuUJXD
QnOwGV4hLHM98ff6pSOIicUxzIZp9BtO90VrNnHCMylwBm++5Nqktcqkf34EnfQI
8BvO+A0HG8OkS6dzd9ksktW03Ef9X3cIOTS4Q98/cJhB2HPggtDXYXAN9cRZLiD3
sxI9Ki/EB6DtZnhCjRqfGrmHaK8LGbYXteoBeR2IMgnZRt1JKyvGiwVsQYSxk7Kd
eepUWPtjSKJby6/Uhwn+5IqEfK8FG+t+UOXgIsENva436nxKAEBQK735xLXuzGwV
xOfUpnQeJ02wIEXAPqqO8kX/8PMrv7YfoHbFssdb5p8vgDvkWCJFldXU432A1krW
nRz4S3izGKRpg/BxNP5U2T31pC75Jn1QBjJrzTXRvP87Fjc4gP7OQZuGbeSlXcxY
2V904tRQgkoyyi+6rrifim28YoJd+CRWlyksDXg6oOBaxmLxi0ioYArp0nNEdyEk
q66SN1w8xSpsjhMosJ93dGnRpUmW5VnbV0MZ6M6g7jGVsdIAP/SdgpadzBDH/51x
F4bpkJHLBmdQYBrCQ0eXIQHk+7JsKYhku7XXjgw3aj0DRmgD9Cz0QICQs+02kp9+
v2BfHFzjVKc15AJo2xJNdKrgOlXRd72GJlYSxnR1bdYSHmynfX32ygNnH92FDzmn
PfwvYDIgLaIzaeK+aVOHZh2pNBMPNOhgr/Y3HT7x5BhA/n8lQouoUE/u8CS2OpY1
2ZlqBkyMPiSRs+XldkjZZpztZbeAzlwtVjUTRuou37tlrjHpaz7VBjkIkzD4BCBT
hxZ0fnpIyh5axk6xMV1xDSN5F5EphOy7UwzRSQDJD3+iVgDDtC1Dm+RhKQ3BZDUd
MSd1W3LA1sFV3qmt0B2wVyWbHM4XiuDGtFINNBWSbztrzj/3kKBfVVsrE/eyEKGX
P7g2nfJQsGDL8Y+fUE80ZHSaJSwmysCSc10TGyWM8ZnsNcOaNhrRg52/W2z5d5eq
NLtKvxlrE84RETIl+AuyZ3SjYBXHW2qwptYg46Mohyz3v0w6WOsul4490rPZjNwN
6D6AJw63agbplCoDEQTLqVObQ+p4PXNl9Iz7XZFKx77Ikp15u3a0W/h2WIIP4Nr9
Mh05pOjV3ggkKyRQB+rBAg==
`pragma protect end_protected
