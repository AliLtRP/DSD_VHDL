// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hApcjeFvW7jualcUmSMXGjfHWghNVDFApO++yNc1zaEHG0u+DCAIXfn8sRv2QNXC
1ZS86Wjj5WJmgkZjF0g+eE74pEijIyA0pZNf/OGjOCSszjgdgpZeNsJPtKeJvZG7
hG348DsJQJInpiH33LcijH4zOc+BQi+S9RkvZla33Hg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11408)
l74f94KM4NGIIPze3JmENEN4Vs5+rjBPR81wcxcPby7h4JaHL0VL0PeR/92UvZ81
Y+OW5Mj6MuiJwRozHEp5rVx7ZcMI8NvbqPvujsDSSnQVikQUuRtcelmwLpE9ro1H
Z3BthM0J2WG8V7SOKQXjel4BEvLJIWzfsUKm2fm+gw7LHzOrZ8uS6e1e2kTXxwp7
vlWp3eN/shjGO36qMS5hX/Q3kde2THnafSB2/r7VTY5YOIT1TAMaIjbtMIKieHD4
I63Iwzg3QdXc2oge25+t8p4MFdX0UwKj9gPpjYSNYmjo7EZpyu11sG3ZZUxXHvfj
9x0QFNVbyNp7hc7rPEP8Dinm8LTQ4iB6hbprqW9mrRxe1q3TTVVKTHyBlhg1T3GC
q9fZ4iSNmQF54r/mUxrILMVlG9WNVjkohfa59fLhlJssiuon4ht7tdLoRfHZ/ssX
hdPbmtCYGOGLj3pJKVKH+u9dvAgPd19Fv6xmEU2ca1lvq4K5WsRvQxmRQdg/eXqA
cBOTMhGejbcVCwE0IeykSuJK8oSf/Rrch50r684HX8Cd6Urj9yN0TeX05TijdRa5
6S1nC57uzzBaJQnm0bueehYdxOfG3+1oGKBITEgxNhwS7OSKdrdJIKKip5xi7jeK
4zo+o/m1UAaTQW9VhdjuxWsHVW/iDC5mEcmaGHgAaferH/hNXI5kRfFes4meU3O4
uY48DwfGm1aiOGFWTNQihuUMqtgxL6r9pPfmfGaG2x6LaUKdkKalCwIfd4f1PzLs
lPu79HeHQ7XU0C1wbYce4bGRypSJ5Ic7zjIITn2df4zCn9hTacpvI4+4QP2ut0KW
XD7+nXNJJK0WY55dSAiQFPi8gm1mkBr14c79ppOkDXhzjnzH0bDJvaOdWdoh7u4l
bp4sWJIqLg+2nfu01oAYZV4g8cmdogmMc++dLwjK5kxkPM2tmj12UQte1xTwPJi6
4rIGGyOxgpr6kgV5K/ERv3vUYvhG1duQgNtuK2PjlEb9z+G7uBCWG/Y4v2Y8Evdd
G5QYCzVrKzlnqhkpAqbBHssOLSfJqAt67BXLiIA4mFYhJL5f3oD0Jpv7TzZWJtjj
ZIVJpla83tkd85a9TPsKOVgCZeSAGA08Sph9wCAl1jR9KQNW0ev5TwJ9ltalw64b
gmPIb7kS35d2WNOAgagyhfoTz8b4O6UsAWm/t3qcMxxZE8/o9gvv31585wFELnHX
8q+itQYYXQD5ycWgp0gnTZnTThG0Dr+QHhZfbNHSh+uLTsA9fJcqLFovkjU5nBOF
lk945CFW1QiI+U3asTzq/3P6S0ef74QQO7qxMjHmxt4XJ1k86V6o7k8gq8nBU+EO
nNsKa9zD9pLPX2uvbSnscs2OsmxIvrVsPm8GGxSw7IBmwxsqKTFEkbfq8dUQRToc
c8hmyDwP8M6Vyn/vFObIW8JU8H6wqlc2O58PxRVjYssMCyWbPHJmJboLmCvYhPjS
nvyhu8dwbrQifKh6tKNPzwj96WS4qkd4D6FsBYP2b3liWk3pq+HIqaUbsV3t/po+
RVmvlNJpP/WXms2xtcJKo9EprARghDqMl49Bd4VHgaj067mff1xjSXK52oQ6zHq9
XI6b9Le0KshA+pbjacx2r2rPn/8DFpqtuyVbJJvlRnxAIV+iS078JVgctRXGzL8W
uFndN+5x7XCrdacWdDQXA7CrZyvYinqwXKHSe3Z4hGboS+bXSFgu81XTmlVYBdlb
tmo3mFfD8hxPpnTqaClxgWXcPDluHH52uksXFyZAYUhB2bvWv1AyX+j4jdjJ/03B
l9qgPsyL1Hmx0+y8AYOYKvGkkTF65cL/qPQ7niAtTtcp5rEoYqz9LYUojyhGjXf1
P+gIoqgbJtyStk4OjIJQAVMUOxlr5hnizU7IazTLGFtPdIXs5WvqQLH53wH8hrlC
da+536tzKFobXrhGNw9DHf4jjVxA+juAZnIb4akcyynCEzUIGrTEdVhQyJHVQVG1
jc8X+f409hxPPmE9MxItGac64Fzd58y+RGMLBQ02CRD4fs6q87PV+s1OIrAoLSwz
0rOQ6fwNYUJhtmtKsSzdtmfLFzyFghdTBbeRasIaSlrt9WoQwzyxJIgT9KNrM/vh
hwMJuzUVTRmoGbWAS5iA3MdssvmRJA33Jex6c6+4GbJsHvhXmMPxHoMEuEsnuFMo
/hyiOThnhZJEalh34MUecs6PIn+BeIuJNIsBwsXMSDsgycFZLwHywPEmb3GVStBb
ezPEJHBPqvLGxOY6Zrn9MZc+Ne8qOixZAbQ5OzA5gmtC5AZ+kMG37rEMSBahEsz1
EXJeRlGwRbIIY6sB6Pke09UONkqGCcUKT5n9MBH+LRXcWOm2yYyeY32dRd4pPC5c
PvbTkFzyFr7SREF/2B4UIKTpYWKLT7NXOAhn6CO6fv6kn/xHRPkOc8KcahroEdWf
bo9cBZCHg/8uURuAnXWks6twbFb5oqtkRHK0l6rcnFTxRoKm0gXoON51kQ1SvtUL
P/b1GV4sMYAT2zuK1kqW2nI0DTPWwq+rObbhme8i9hod5qx5AR/yAPgtBmvspl7F
hWu+V5OhluyhKlZfphkgIUmiEdtK6XAYOFcYfHxAPlaEhTxQDRLqYDhqUGdGBhMs
XfG0iUrj3FK6T3+koqkZdXwAAXbhmQr2I3u8Pe6cCyCqm5Nsm2JsJdX8fz+f30JW
P1nCyr/rAZosKAQLxj+C74rZkxN5Evj3jImP/YAQXjw2brcah/b9IJ/6hS0/l4pO
qMejm4k9I/Gf5uTp0qev3O8bvRtjstS6u8I38PvVO4YrdESmAgiPN6IwSUkzyzRR
+K50cHBd5TSo75nkScSh9bSvsc/sEeAE/teqvvXzeJBCTa+IfpUZv+8K/FR7xaTc
3kOSNpVM6EZzQ5VdSGfSjjq4bk3mcXFz6G7BqdsBAdaogJRsUdXde2DlIa8CYtRE
vhDT5/SF54YyQnqlzrChGTBpGjrAT6fYJD4GOrbsAtJnIKu2e/IUkcLbkWTbfmvO
beCMDVvu1jeClyOjhhyR7xsnHsEotfE8ZeGm9lbR96IyhgUFNifo+HnxNqPalOw2
rE6kfHag4m3JzQv3R4Zaaof3q25nQJLJo7UpUwLLL2Gw3+zSh9dPNeQFnRfY47Ly
CKz7mrC0+slgWBXcqmvvWLoXsvhjATSRhvYHAyNTe1DKmCRwTBTz+FPBNr8DREpv
ed+Uoc3M17cZc9xhD4mxfbQEKNX6lVvn/HlnbBtxelIEhm1RK8q8PCP/V7v/7Sol
L+s/3ThGzDysFLTJiWof75kYT8kNc4Jxu6SI5x0rQIWQvywM3MxFyh4E2CfkFZXu
fiXtNS2u+4OIet1biuZQNSOIZtarypC2FBw4hdhzQYP4qam3nML67OG3ZqaoHtKs
Q7pPP9ronebeFJc9FJ7soPv8sgiLMcwUUSgG4Aiv6ipBi0BrVhIeWv5WhYAtJn0m
aaZSxhDPB16PRuHOOwsMZ3SqFqLeup/TQdv6ittpYjxQtVfvoCRZVGwGufkFGMDO
bMYtHCMrKAUP4WOqrh3rNOUM2RHLwxHsO7H6FWpaRZ2zNEcNFO/ra4HUnO20iW5d
bhIvPNKVnK3rdp51LM2BQED8lk43D6fT8PmVArn+hdh1W5YERy2FxWxv+M937cvs
k/NPVP4JL4NlUMbqDiSIsX7vxSc40dGB6MfgGr9vHezbRWX5uyoxZE59helFsgDQ
uDydJ+L9UCVpssVxMiJY1dNmoqOwSKkwKsheUIY+TuJrfoOP+/bWIApT91w3ht3P
OVNK2vYPHnmoQcd8+u7qz6vmuOs3587Bjz06lsqt2U4AV156LZvNSBE+SpS4VE7F
bKONpPZM8vIr68d7spJ8lz11eXt6Uk6MiHdmo6a/L3VsXe4opy0xO0U7LKv3V2kP
jZmnZ427ZJ3P+huVB7j3Xy7F+SZ0nuXHimV8pJhGJxaHmLcrMjyMsSJCNp81lPpX
EqjC8OQavBfTARmhCcOdJZGz+A2X7UP8rmLfmLxGE/EZTmOcKKfBhyWQpJzwG/TR
lPbzd9/JtQ+I8PgtsviyHV7hCHhSpwedXSl++SWje9kbWj5mg1WEifsmKmVEe8lV
OJDYEqDHI9Se+FIItWpGHZ9GfqKgzN+KlEzID7c2ObUU997Jo22hYUYeukswjGKa
ps4o4kHGDhs7vhfYaSdUVPYMsPOFfnL87M/JHRxa/MYRnWuR+Aat0KwoRLwvqoA0
Uk+/bpd3ZiP5vEQZlrKReco/n/VtzxwTFEv/uIecmktXfQxPWO7k4HRYHlVfW/Ma
MBZZnzCg9hKt1WxaaFVBVIokoFRQTuPkLCV8loOWL1fB7c/Mn1/2LIPp0WxJvo6h
+6GnwufzVuNJsVOn1awt/a+fHPTikC7T/DUk5AJYvShp9La5U2vQ8bqWnMhzvlDN
w115yLmQvMje2tQvLTmZu2K0Nw0sSq9QOCxzw+rvJINJjFBDHm/Gu0sp7h8G1Ilr
uCQ6iGRIEWAc0YXcz6E3MWh0TGMs8PfIEkJyapQecPuUtLs7jE7Zj9pUc69F42qR
xQxsGVQ4IMp7xr+iVwj5l+YOt1TjacEvWBdSBx/1YZC5bC3Tom1RfB8tOmyR3908
wjLfepMyGNVxsug74vQgNU2yHpOSf9ZDaoyIBcvpsBW4r+dyXfGSOA8mR0J8S8CI
yucI9LGJwqVwMZoawepjiLsk5rWQVtLhZrdlTI2MGvmIYWJPm7VyNor521VYZE/p
mhTL8QoauGpR6e+8FhNWV4eRhRbOseOus6B0Ks3CDborafmPe6VPBGJOc+PofgPu
gYW5haoc8gWnkat7sZiyrcLGTN/OLBSuMet9uUYwgLGJgJCNmznYfZsv/VdwZUWS
gbhNopaew3zHUZMjXpSwZLpBJWxuwO1hmc2pCsOJfLRpr7KJ4wfXkBe8gm2erIEN
A7icLXrRtWe47xMTJXi1HKt59iOMiTJzFPt2FCjTxe0xrkSHdvkJ3W/MZw2xs3A9
r5oHw+Kg+n4VH70DOv1xrOmi2OUGDlu7M+2+XbdUr+6ZRUnFAF5N1+1tRchv832a
I+CfcbYppZJ44lG5BGboPdJu2i1kzgEmXAfeK0//V6jp7zdthJZqnWeNKlYVj8y2
MrrtVsWWkrXnMBsDlGiIi8z50jwxMoUz9XvIP5bSngYF/NUGY1gMyqXPy+RWNw8G
ncxFkZCnTKsH6Ngf1dekvuokrWQwZSodwQEVpYN95cGHfQ99h4NO61une9hE3WQR
5STw9USCNwuPF/Lf7yHG1ZxDr+xbiFdDnE1XS4ZMHy+iquV3X+ATkrILczlepngi
zeeXtUDUdZwz+tVLrzGgU+y/6BvD13j9uf4IItxy0yrh6yySsn1pQNjcyfEayddS
MQPrd/mLTqM8PpJIIJxyqbXzUMCNr9M+Ce6IRWUqY0srWUJ0ObLq7/hqvTbajOXG
eZamcpwA6NiLjricflTEk8aug3Xior1Eyfju4beZNt4DMThq0ZOIXkckHn82jWLP
ecKUBzk1gjwxjfYFEfF8kHOzTNWb2KNqLNGH4/aFQ3oj180CM+sjSiEftPaeFCIb
jfISunD2yM1cO2l9sJ9lyi3hVZuR71mtCxH9mfKTVEwytXz9il7YFw+alCpx6b90
8uY3aYMxRVmg2sT8nIN2xkrP6wOKI9NRapTMUXSDm6ADc/RZ+qo/gagNc+qH8FG3
E/5gWFj1Sp3boNhSobLRQiRsbm0pf1p/J0cv4+Sij3yEeyWx+w/T6ykRO4pdVeKD
A+w+JWs+EOhobBbpoAzEalRFSPfMtJQ6VCbw48q9t+0WyJtSofRQ2Q68ni4j/diP
yHIyLThZsT9/I43HRKXP7vLbzvGZdSsFDeZUFCsYn4gOWCbHrS4hDMJsVU5J6uwG
A/gIQ7pq9r+GOWYByzYqdGNyK6ZjZN0NBkGSfjcq30rNrSfwR/y+Lh4iRS0NcqPF
0WmZojQwWvvkGiST0YQCnaBMcW5WuD4aLpUWba4kor2v0jMvDVizcfNOMfI9+xuE
+ftBvHQiIYztFZRlbUuR+h7gofAEYgYz3nGlwaNy7KvoU6CwwXqxzFkDRUVceQNu
fL6bze/XiOPt483086c+0z6cX7EEeygh34AWmWEg2SXwf/1ojuKQJRlIkI+kBlUj
vFMs8snoQy6QPBSyoU+4WT2rFR/SkfDnyFOG7GtMO4zH+NgYIU/8iXrv7foo6NhL
THYOdnXtw1WKaD97kafjOj/dmwq5rFqdY/Q9KVrRpVWt3wbM9mlWw8eIDiVx/OXY
bFaTpVyfDq926oce2CVwEL/4DJEFgJbqFZEF3Hz7+IAYwodq4QyNx1Piy10gW6bd
ouvutOeG3LFsxCi09qfSJglj6KUBhx4Ozh5XserzWczzyjimmMX+T+1A1FvN1cSv
08758pbepGGSaOeQF3ELUTqqDtgMyAqgwevBP79CbBqljg/ne+qZrThuFaANUNux
9mPR9k0+GIx+3nqLiUi4RwIRxUq0O6KCqusmbZqQmSE4vUrZ7d3i89mktE4Jz1dc
ncscG7ICSu4fkrsdoGFhTTXWTXr1gN+1wRO7BiGc9Vu+0IZVw0lnEvuEyibH2bx4
lTck7aAdiI86z4D2rPjoufJLR/Y1it/swQL9bVLYFv9CiqohQK+Rujklvg9BP6nT
HBCGzclDNxcDABvhRI6vsDFW5oyZNxmsibPgUcTAj3okXGb1lZw/93aVPLDvOl07
IHzVmRdWlv7zVNVnC2KxKR0qUe/AqLbrj8e5HO08vtMf01l2p3UJsrLkiJErZUW8
Z7HtDGbK60e4iToinEnODLpw9yOICWjS2Sg9PeDq+i1DgjgawDkh6mSYAw0qD61L
KnHJZy9X/QY9CEy56jSKV2Ys4Jvs26UTyTfvEDY94YImy+7TaCsd+i2VRuSq26lS
B9WA4EJQ/LylbgwaLyCqipXF5upRb0HuS3MQDS4a7SDL11ycHwjHbZHLyc/RWq01
sVPMwUNWauJf7Q4TkdpsBjwbbmGZZpB0XnUt7Y69KylBcMgpK0+f6yEVa9SrhAkj
Fs26Bfh55CXhIWxYmL9KsN8ViHILnoNgyGvlDWT7rMqlcC3zaU7MbGZtalYdaMGL
uY+OZafQI5YRF2uUEvdJMlmiRr7v5PFCd5FME6cHUDZBBCn19+Wy9TU1XmFPYlUz
tbgQmPz1O+4dGTLYmzIOAOmVnVMGWvB6B4LZL3CR735yC+8Pbz5aw+iInpMjk0BP
hJT0OQma8PBjHCBp7RGwtIA+W71GLL/FY1khUYA5p404WbIcoxog3GbKIVd17l9d
rfGtPoQWvAY+j82o8oZISqVr37rbDbw2vxwZ+kdqcpQ23T2eG5oGWJwtxPMKZDaB
xugNjcej8JYgPDz1viNOZHkZl5N1ycSNHd/AtU6TOl+zRIBMFnYBwk74UJWT19qR
AmVJthd0dJk4f640Rsun5oCzTK175TJOStKh/VjVd7J19aI0gTXNNnOS/igsB/E2
d5jdfGIkjfa5Oe8JIcES5fjhP+WNtyqidaArf2cIAhqKE2b7btCQHREIFVCdbYPE
sXKgs9GvyM6XvI30MlTs64aTIs63aptIPgvAnHpHk/SF1w5waqDO323j5TYQGZFW
/XhxL05cclxSCZr4eE0CqOCpnjNrg2Ji9TNxIkhlVO5a4G4XBGgeJUvRMJe8Rbyp
L4wEyh0ZdKy7X++ZC6RQ3jP7Uj9OVFfz2RvmKWX67rUyatQdBgThHABlQOthOoRG
6onrZbGODmnFg8rB+Y8Vu9bdowhC9Rewn5zLixyZqscIIqdqb9E7koIcf5nj7AUI
j05eb4IAQlClmM+m80veZ4di26P/Tuzy/ZXBJKZulBFsvToOTb3AVe9X81togMju
/dL0Bg7SaulpjHIMNb+SLUr4+7oNvwbJAhSFIZ5joqhca9p2shw0s9gSd3pIXIoo
Axa8+3vpsn5Qk0mA8G8GbZOQecGLDaIy69WmccEzrRH4WM/GnBeV+/hy+NAquJ55
HJKbL3pKAleJ3ag/MnGtI2USIl7IgZ0YknkCiBEYgx02Y13g3acjwNkx/VFitgOC
FhdRpWu1KIwoJsWypXtQqHJgqkAVTQXKc8/AsHoxYqsKa1fxq4SPMkm5zBLEdha1
Ggv+jAD8UJBAvVb6gwmIny7GA/tS/otZnv8PNGRVNkLVnV2Y28++IgdeTf8LoNiW
Gz221GoZbUPIcI7dcTqjVuxpIAtHVcUaOLHuVfELV91GdQ8X3vuDZzhAuprpv9xU
ECFA1bI5nJ1dY1dHxydClwGnh44/WBcbTB0ufdg7a2va5m73ucRH+zZf4fcIKPj1
UiLH/A04AJ1kTn553oWsizFjPiv2jCMcYk4CXdZy2L4SasVLA0QaDWjHXx1bn0XX
PYxvHLR/GHKlVzcaWjNf9CPXjzBuF7hKk+iopBc0yNWLs0Rt8QhCUYCONctMSw2Q
FPDrbFuzcyWLKT/w/Yq2IfSpPd7BdbxXYNpIJbF/T6J4C6ZjpwFsCbc9sAus9FFB
2G146HiUo7YTo1b/MQ3rH9QOq+vGog4tpw1LpOQCs98s07P7sVYZK5bjJLHzHDkG
5tkKTIbHwTdmYMAXW1ZwWewpSPgnudhRzBEdP4pJyxhyKfUSceYZOtmsoAgafZpM
WiQ3lrc9ootZ0zxZBSSlJL4QLPvCyWu3J0mnGVTSKQaq5jekZbBEVUZypQN7tEje
i6BhDRG7YRhUDQjaKPT17WkQSLt+1g27NkDnLR+6AXNiM8mORn6Q9gbIHHi/H6Fm
F9epkznPoxfR5v3cED6f/dHJNIy7cCvXXggQ+GPF6LqK6tjiWoljYYwr4eS7ObaY
x8LchmA1FO4gu2nXyPo9T9IAMYbGWF7NVzRgbuPmCUgx6VbbBL5apX1vzQAGbenL
3zbcYCHGj7qIS+3NdKS7ROqBeTa8SkyuyvdKdIQmUxA7V/RCWIfvBKseDzQuG1nZ
jpT7vQxZJzF6Mz6pjznlqJV9HS73dhzXJG/V4dUCtRuMg97iGyGv7OEqkn7rTS7r
RF/M6N1IHH4TbrGwhtu1D352yqCqWSRVZ1yH0DWztwPlvUdKnCdR7DhAumfLe5O6
eLTEtnLIBmPinWMrLhipGd4K9ZUGGMtIeS1VCTyVWD6W0cA1u8JprzKUJrm9n0x8
5Gud2ITWWt3MFzH7ADX7KZsvqrkOt/PxnVNClUEz783LPzG+KvqIj4UiKBmJ6oiI
obO8FG4cWZ8qimlJ+Qi8FzqMIkwCIMCQTClKjneSZnSB6vNQwUqaGeAlX2cd6jRt
Zrmn1I5d64F+wdlD/hVnfJ5mb2LEQvKsgROmVOC224uoLE9Uh4LLqB/afg3tiSpH
/qOHmcKbudUqfmoMYk9uxQ29B2akKQiJDwAlpr+2R5KawAeP24ufmrR353a73srU
g+KBhWCvI/S6uL7QhB2sm11aiDwvZAywxRORax96cu3Bc5duC2JCgzgAlMYuf2mT
Cx9vx+lxMb0o0qjU5T1o451hB6c2WJJF18XKVH/cP0ihrq5Qv7gYZRju1WleyeEA
dDk6Xa6vbk63Yqs8vj/RiVwc+YjWbhcRIpkKnonJHGXMQsbUQROdY5HH4+6YjM8x
vdGXhZyjrebmBj6DF772mOTkMxjWGhiB3E1KpVWnFrPK+6REU1dT1HyCdscGFvSy
ooDcSl2bla+Gc3Ck62uMUF8tiyDFTFtmGj3ajgQgtJ/lYAStj+wGhw9aoeWJ9Y0D
14nK4aG51IDicreVEcyPwOl9bLFNNrm9i00V7tMNVNgWsRkQwyIYIh19wDTkgcHQ
ZVmpVh3QRVTas64e8jAbRojJibDFra55y0UhQPoqOIg6hA1ptXUq7pElegtPWihd
z4hPcWuUIDjlsKKmMrPEgdrl4a0sT8eTCQlFmpusCEd0IMTDW6Ng56yygOFLSMs4
o4Z+woNrYyeEawdOLxG1TUuxghHCkLy1zdvKqUhQtguF9ZB7Q7q1hL97RvUz6i70
LBNzRYuCFnesLeVWhiam2Sk+wcqq+dy8d+qkInsoho9JodRJlu5LM/h96HF3pYhi
5ZVRPxFtBK+XDWhFxn3/bk5oxABZducjdIwuuLCPV5h4AqPr2On7BPaCZKs371oe
otLC8udPbg8Fz6p5VbHt9cUP83Ryha3fB6jGQ1CxZ+MQSw/LlBqDHtia5vSb2Ifn
gon5FBncF4rHPDRopWQugi4QbJnaLwSOH/dDpV6nRfNUE20ojq/S1f8B1FUF5faF
LzAtLkdb7zK2TkJ2vairhv17jdm7PfhwxAIwTN7FyFDvT93djXbCXy5U0Bqx+OcX
yqsTBVzOotaQAJSVN2/+ymKM5nZuhw3je+0cV2UlKrnaSh2BhwdOLUJR5uU7TZsg
mn/ShvZkwpd7nRZtJ+nnyi1s2F8GbTYlqhCDjRaYVEFMTGnW4G6qY7GDloaPhqRM
I9INcL5w7PazlExmMwMk9P89zuGL7nvvOgwIIhwh2x8RhE/csMb5st93SWkEqF/h
4+HBod+w3KYhVBLu03aEGkwlNEGhoJfW7ub1dJKPdAaxhaFs4HRcQ1IcGhYSqhIf
vaSaT9eGU4qaY1xx2CN9f5aAd1EfNj/3wFnJDWZPKONyhDdoUVn6WEr+uEL7Go+s
TDV643zE1qC6Ix3zrBkthpiXgEaQKBfjL0jHaH8O1trVxUaCH5OjyvzvG3/rPJu2
jqOlMPXO7VwRPlemsMkQt4qhgyBc5VP/VuDPCr9Mdg68fGmWuQic8CLTpVHcNVIR
Lozy+kNJZYxvxPmV5EUnVnJrT2Tu6pkXh6K9fzdsCm+T4dWCxd0VXvlc11hxWP5A
c6eVP/ZiYKb77tHPYQC2YmC3CbU1+1rD2Aw6enWjiEztZBSURQfYSibDsH0pQno1
MZZrrwWwKi0XSeiidGPWKWYsut3DzbJD8QPz417fRiXKMer7IyyexOwhFpBPDZsn
k62Wg09A6MD0+1yZ1RxriMFwvviKvODS5f2Pl2niNPWmvu0DDnsWWaZgFb+LLoKQ
vQY5EOBGxO3PeltjzDv44vW/YhKSw9rEpVhqDMa53nGcUISlIFm5thDnnpD+GW3e
lMIeM1azOKkPiW2KsVbKWbPcYOy0VyfYGLgySULy2wmG6CpoE9xK/hR9I1Xl/Vx7
bbkz1moWJx1rhM+qZYIdgMfw1/AcUYwYxjgn3llcuhzKLn/H9drx+303D8I47pzi
i2edz+h43gkDx4OnrIuvH/mtwo2TNQtoemav+C6OH5qR5Gg/FXuCGE7JGL+KHhDb
bdBsooGujqyVjB+WkSBdiCol7um8QhV8daXNaMf42sWX7DQGj8cF4tuFesjJcvFG
9fUwx4kax61JuVXOBD4zSlNgvv356gqEeq9nTNZ01qzLE0yf+2NYDA5/onrrxvNb
fDT7ydW6zYO1wWFKY/Qw0lNEw5fmu9kdKT7gYaXNg61TJ3s3f1UGEcwsktkxqe0d
utWU6NHPkDkGtJnpAYw5iGEwYaioN3QfD55bH0U2yStxKya+JChiTKHZ86wJzMwF
xPTaw5UrBbqCD8ePR9jJAEBbuOOTuYsxVHjD1qdDaDh0YwKTfg4PqoBW9/lFES2X
Ln8NwKqTIb8+sSwdNYf4uX7dgSiqTAbEk1yglg3PYhRybD7OMlTqt+tP2aXU4vSV
v9EE/7UyDOD58svLGlyNZWai7yEealXgMpBTptanfznpCcHZxG4hCYKFE0xF6Ond
OKT9aKzqk/Shb9AZAXgRHeO1teg7TKAUQhMvOxZgvMYjcW/52ABeAXedT/a86j+Q
ruGYMItkhKfNQn0xrgJrmovV1PHUAFr1Sn+9B6y+KSMhmHmVuswhh1rtB149lR8P
X9G7z4qIIwOJoNjt24DU+/rb44Q4BLUgOELU1vsxgZsAUjM9AcIYzbJqlqKqLV9T
ubi8vDjkU4KBYXRY8xly6rdaV/w2VB922T0cxWlxdk71UYdU3zJXze2h23LDpuXW
y52VsHkgSjBhYSQGmyrTYLI8hE8L+s02n53y7Ts6lNo3CY9i/mEK1W9jluzTTPAj
sdxZooaRuRZ6XwrH7/TfWRChVXAiKSSksIN+SHFysW2XwyZhzqEP3UWU9spzV+ew
GwRXURGUK1fZWKBYtlbbqdoH4n+Ug8m8OcX73PjSXQriisx6IlT9vM5XYWWQNv9T
sWaOtemk/+oiBUAcSZ8owCYyF3yFtzM0MyJHDc3ngDLDs4b1ZSSImp/gePEzOePt
Y4lEACjjdPtCZ00D7sh4sOqThh5zk/7edKPsI8/+J2EwNMZhK6TanEUdw8by/NBA
4S5WSeE5VPcWdFgp3RzTOZHqo3la8kAmUcRRNOxY0a9Fk0v9s32N5H4jR7o94YPA
odlKWeBt1lhEqORfzxXOSK+QDGE6h/HH5rWDt2Ibuzud/CLim6hB1fPHmnakI42V
q6+wWU5bDRJDmrqIFanL+Va2J5ZAg7yFbZzoVO3oKK4Z8ncJzjegkNv3aKVfCEEe
TAdZQU2i2mnLEjgHXD/Vx1AUTu5exeRrqd5nTYd/WWwrc/mPMGU0Glu7EdGULvV/
48uU4m2Zun333MkhVOrcw8+fltXKyuhQmB2NATJYMH60e0TQSwY7TuqwHXeIQ3KG
oDpQ4RaZxZtsnyvapa9mLs+PKBeaOyKk20I+WfP5k36feCd/a606nMQOxi1dKsLA
7BPAcwkEvY4bA13rv3tXhFlCSPjymsLaGi3VyAzwmwDaFegSwe2UIPAKQwE4oWdy
t4MsG8a/16XAk4ua7cofA0oao3GwcyHPAakxd2RJa4kt/9ut6VzM873pg8aX4cBC
u37OfyHVjM4yK25dCW+Egwc4QCRuMeDnHpnbozD7IBkoClKAsWbqTRtiJdF3sU+T
TNJ/a4vdTUuM//FTFy3xAARViI8XIASLG3vjTOhgy+v86q3I/6rKvG06dGjRbvnr
fmjtPy8lwICpIFUkJNOGg8eTTOWUOlRLFgehQADNbY+8oNlEyUH+xbWdGVs7X9NV
xrOILcA6fPmGXSNT3ogt2C9vOPtf+YADXBG7O+s7J0rDd/xCoQkvBFa3t+iTT424
KuIyEWfHiVMiH1eCF6ZJ6FrkyngQZwkL+rEdv4aLxkaTYkoE/jAsk8DaqbaCW0KO
GDCnKg4wmR14nv03o3Y63O+kog5o4sG5RF5cbEIIkLe0azPtKfDX9dApac0uSjJK
ATnxv8/4iYppZjmLYG0hKVgddCrWEXGN7wMdCq+OfTRGebiVViWrb+yitEo2/MnL
psmKKVx1t5Q0eZtHVWEBUBiK8b1ISMslfb9GWtbPkMEwrD6Sw8hkVMnfb4Dttyej
welqNJynCQONeeUePVqoUEBrMsaDnwMuC0sPlXXHXScuzat3OpzQ74NIkbZt555+
xewB2/aIiXU69eLdw3b7nN6SMILH++b+42B+bImsJ9oA9Bg23f49GhDi04/3+9xz
0sZFn1k/xh+2UBZ9BsMygZNwUAirtcvXg7E27X/+WWkMRN/rRemYbh08umYfy2WN
ubmk9MTsz6VdEqjXMbUKwIKifs2EKi/p88ziTbmayANuofb9U3Ud4AAMPShJs7Ky
dRIBf9Hmz4Y94rK+dmtZjNjdgI0dldnz3/Ms0ynXhgzAc3MLUr2nO6J85NR3emUp
1yWTZS7z7KYs2qmhOD/aaDiH536/2KwlDdbWF7o6e2IVSlSNKlAhuF+iRe/7Io83
AZDX8LcDjw4iZIm69nvvmL8+2u3Cn5KUQqymEjM0s6XmhvNauCOROuUOhEo7V78g
wIsuWO72a/Dd6bTdXUma7LxJGS9qHbOELangzw4KCmBM3j1FBP9hdDdh19Kgglid
DIkbYOMMePA3xqn2C/axa3Fcp6NYJ/tqCLVgT+6ud8j6C2vN7p2DLrUs5yMLgevv
S6yXb5e8RpZzXcxto4X0/K+vtIpQMsvnwm/o0tmREzsHpaJwF+HegYO0KVqzbedH
/GbGo4kgxGf+TOY/s24PZEoSL0R+UV17fJFhw4gSJgFd/ZD8LvqMt8nrCMAW8F64
yPWsCKhCRaMgZT6QJKSso16JMsj/tn3fFM5PPMD7DvPEgRie8rLKzy/syC1YNX82
TPbIGj1D961UGg4EdXC8C6aQpjOyi1Snni7ULRxrUSGNrwFqfxOJ4dq77OVQMUgW
9rl+aT+Imvgl0ZRigKlRKWW1VK+y6un5r5r3mwFx3x39+btT2F3qIb4YL1B0yJoi
bLYLedOg5jPE3KgdXI7NSL1qXbc83f0oxJWm3YqoN3JOW45VIpD6lUv/SBSvuHtB
2M2ewuJWtM1btgL31HsSevbbBPlLBwzZovubfy0Q1Zgm6+t5XNdgD4Z9i71H68WO
r+aJ5w8NwgPyIWwrn+UMPYrCSMTw2iqz6CgFWLEj5VuQbRFg55yYqo/6a9R9aoX8
eJaDRMLh6l/YkJHaGn00tIQ/7UMMH7FkdOFRvyIcdTq1L2scEKiN5WAAOVsBhMJQ
qcoZHFrsGe0Tyjt3j293/W2T8hmwXcw2xALrmDT3xqLzXJsEqtk+IkvYX6/9oYlw
6FjHTWfqeTyP9+cxJVuYhXTpXOstCShEEeE0DE5iZUVdI8Cvzx4A9d9b5vj/I6aL
RnnmitYMPNgb4zkj4soK1xDH1YoqxLnwcsdXYfRPHU4pwpLIH4gA5+zmrKezLUlR
olr+XGvTLBAIkum1T9hQLdm+CcaiROZdgnkmw2oblFFrLZO4y9hZj5nGL/lZ5WhU
ziF276b0GKLwZuc/ksLKb91T8MtV09N7GkQJo+ACJ3eibRiO31xw2aZKsP3Cw1lY
ZSi23qZXTgJRdY+wM4JTkhwkVBscw8KbcZ1ujeDanwp5XJPipYids9HFYTS/qYI+
Q6ls4dHwi+5CSIRui1VMO8sbwnbcOGzH3VUv2cQkbIEkc1P0WUKgoZBUE1/ERE+p
y90S/H5Kat4BHLROBzi5bgKOVoIhxDroenz4wQdOwHKi5kjInwT8SgQvaeSyAumb
QJjTnuE2CdSLcHk8l4i8Z3p8n92eJ/HcsD3x3BSdfvD4BOh9fhJZUuW2XVYk3ZxN
1p/hRiAQkwunk1YbepYUWxNbmFXu/4Tw/Xj7ne00y/KCYamdk7+75c/0FrdBOKWg
C7iiyZaqtIPEzHSNzuYk5NnixA+UILjMF2H5qRbgLALMrecOqti4ht9bMNWg98Tn
mLfysKlA1oYyMJE8w2yhAvjF1Z94A7Bps3b6U/LMORQ=
`pragma protect end_protected
