// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BS+OFBHhaoBKr0hiWschngu6BVroUhjmULSZwZq0CuSKoilffDgaqopExvZTiBUy
6P69HQDH078OqVp+GNKQyIyV3fF6ZjwvME9aV7vFn0jwGaM67XZi9Jvh8g6LcdYd
DBYvvTgGpWOhEC4b+tfd+Ze5cfzhHoatJUvfiCvKKj8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6880)
B0dG5QhJwJxd3wTJOYDHxH7JAgr/hbmEUNJh6ZweBuVfRl/pAAbcL/PR5jG88dK3
RhBKFWq/osa6oM9LAv+s3NBQtuvUCnsLxq/nflW5wJpI7xXourMhFampZTGH1tHt
5iKIGqxWhN+DXgW7EaMYDojF5EinzjbiJhMza2DTEsUcWxCvexGffmATJGrLI6Ul
bkFiXgZRYq50yfGOccEEzrmrBNcnalWWprW0gNdX5qy0t7BYI0iGFNeSPsHZy0gI
NKF9hQ3C9JpK2PKjz+aOifnHzQbegMA4EV775fnetTmD2nr4JgmuaNx0w18bR4KX
uv3GMf7i1RE3Lqd/Z5QxPR0RfIDcvuhuOSEfupfls1OmDd7fLZJrm+tXe97wTZ5k
ewSEViBG4ZiOnXVEbuFe3wYQRdW4Sk0oq1+mObaiBR00QIUqnD92FHEeO2FY89iv
ej6V6Q/sctDU7SvAd2dpLAOHNF0Uy2vazmxiQthflkuLxUiuJuX13TLdfRiIr0MV
Df5Jhsu7NiqVMEnB0+4ImfqgDEaUJyqq5aLk2kjCk5x3EWddy95inkodXVdPLEYY
r49+dszytIrezYBez+6H6lpWKNxUNv4hY5QzeEKps4ewoKCoav9+QwX/u+friLrh
hIxV/2iUTB4PPIWSPOajgq32XfAeXUPLsH/HSq1QaTCHZbAE2K60A8nhp67xynYE
ofVcTL8jEgB6K6SfznR6rB+G8E4zMvHV6I+yNHU8iNkXroHaUVHC1GMigTYs9gWZ
X6A2J0WX/JfV3pJ3lV9ZxH76K0KauxrXA0yMp8KaCE/Z6MFpBZUYrUeAqYvVmSbG
nYNgBc7jT87WPurQqTNqAT5RFDSvacmYF3+QCLSP8d3uWf2INtBIhdhaqy9hOoXO
PePG2QOT/MVpesVWt6aNCNJpsPFgyqEVGdz/PFc7CyrJPPDHO+QVGnhea/Q/Uv8g
i13nrNqkv1Pdn/AByBmSU7S6p/PWtCs2pYKZrytSb+u/HdGOm5N3ZJLpDllyyj0p
TNHzpiqpIxwR8a5mGQOgQjEms9rR/2A/V+jGPxQrC5uyaR0vxRK//ITpOCwngDRd
ugns6PfT2apIzEmDvk++YXP2Dvqptj3uL8P21ZH0PyvXYoTGbL6tPAvJWVR2KfWR
R+mTYts2euMcnw6Jms5m+twyD2soLlaMKl8BfCksLgbxfWH/ofbTgWlT9RUIaYwC
+ctyNEmVF2SNGHtlPM8P/PAwvXqDHa9Zd/L6Rkxf9/pHJPbHF/EeVzBUfCwGbuW2
+4tblIhs99RUt/1Iw740qtDUuZoWcHfWmgxT9DZQFzIGu+lp+UltGd6/ZebjkvbF
nj5/hnuANMVjJ0nldkb4CeLrcgIWYn7G7NQMMYodlloRUNgDPxJwNSuJSAZtAH21
CZSA+rX5fn0QP23VwDlSH+eDQZx403jxiHEw2w7R/e/Nv8zTA5e8LzLv8IJ4XdsT
pGeGK4zjc09rtUsAIwGJnjynbHEM76ggR1lGRBK4/QqxiYbPkTJxzuXTMkddiJ7I
0t6Ez2Yyps7Xc+ryQMGHDxKZi1vcjohe86qVYlx/5ikxLx5xm/NqrwRxT0AoLdzN
VjzGX+C8/qjzSXDPmV82Whk4Otqf6Mn0J8d0Byc+8yDSPYP01rJcuF3AuVGqR8W+
tDXAaUeOS93vdtzMMQONs1s1f31i8hvJWjxRW3vdcv3ijuV43oZnGVUcZucv34C/
GVwNfj92rRrFNS4gZ2LrxOq/Ke6XANcpL1bXZSogyq6yl/DVYWNab8NeoP+WmTI0
IZISnY3q0wFKmS0agx5+TTnUW9N5XxBgj5a/VefDQLrTiplYSTbfT7WXUt3NsUNr
kcTRPtccVwh5rX2fZLsWMet5Tw7QZrIfDGTYvLsot4VgFlaVYtByX6PJazK9A8A6
iKIkuLKPKEnzYCK9wcPpTx8jmqJUyUSKNQ0+6569sapOf0jGjFv4V4AWxFt9/sr+
jo0uvw/FZlfOAyt3rrIs9ENlCH834u1uI7vnARvGkAu2lnWOl8IxIPipANKuvcPp
ZwIAL88ytVV9xiZjtiYjWShMSuSjLAvgNCVdZQUvEQZV9oJekjSAgNd/Wzb4h3oE
prXi0QBTRQd2XuD3uHBnb6UTBt5GGh+y5DDscC5/dHc+FDPdHL+v6NhGLuOy4Hz2
CKq9mJ3X5siScB3e2PWmeJWmprVKTMrIe4tFHTGHwrPH4u+470e/JOlaITV8r3ei
szUYRldTX0HTbl6FPECM0PMMLZC3kkjOGdpgXuj99khQrf3PeC+/5PVcHtrC4UKT
IFLoDpP6E2Eb6zDa4F0xmaE6Et9cXq6H6JPssMNdKA8P7b/UZpp+3LBoVp4Q/PWB
2XsxGvdji664DdwFENatRXDKdNTmndz3kC6nmGaWp0L2WNMuGUEfKUVsSS9j2fTy
aMtTMUnec2ZBWvWOqBuFtk/V/swZ9DSFuCZj7kTVqcHvSgBEuepq9oAIe6aCbRsc
8mz/a6VpKVcS8HY0i/zodo6IiEU3yaDf8ngupQoJqBAINkxWYrHXufE1K+wctBP9
V7b5PwqtEiySTk1UVSV1DCK0q/pUxkjXYDFANa+1m9uWpXbSojZQ8pwi28cSPXSQ
rJmAzvhCkXJ8fNOwtPqkMDJm7lmXVhet1vUgeFUsnBTFLBgPD8nwkFpMEezyb42q
kRY5ArxIwzilniYa6d/aKXjRzYpAAJrbyiw3P7w90chJ9EPEMd1eVT6PvsPnLkV6
TUoVfaAolJVNERm9M3hshMqyLx6oi3ltmLpfZG15j7rHRN0x0FYfdJMC0nDHVOuz
8IoUHQgQ/uj0ODGJ8W/8SmZBKWTsE70rZMKJTg5lqsCBlxCgC0m8d/YE86kotHLi
0yu/h6wBV8GEkvJdmU72rpcFRvPSZEXnP/UiGi6lr8Ceb+gIVyifL5lxXDGcP9JF
hck7p4pS6JWEOe1Y+v2t8XN7w3uqHaR2/Px3ZDITTerTM/mSGCv1Hnb0EKlh9kW3
cxCrDU4ZwuAyzHvRQm/ahMbsKOYTjgRnEsN630A5BxlO6UnSJvi747iGbjXKR0vO
vSiBTWDxMmsSfwnDmOZxCrQEiXrsI4hX0DP5PQexQg0A6QKQWM7qlJLlt8IqbUcu
5xnf5ORg4d4YKZPDbbBgpAbFIuxbfZwu64YnCNNSgFX2SiZWyilMVAosyrgxKoPL
NzNACvGZ98MVXNJFB0kS9+PMXOQh35QlJ1FMR8otAMjaTK3rTd66ekm2ZHJjayc4
RTJ0ToZnZrOmzDfeZJ1K6/oWqxBrj2Gs75dYXhWVYcZWtRyFPe/Bd8g+ScHydFvx
4RE9JPRfjqF443Kr4YJlbe9WGgV5/acDF6YcMEwPXzoIdm6f218q+i8x70gFtfqf
+fZxCPwSFJvZzx/f//hCu98cewJXar57xJJ1X9X9s1UILlLdpdDkZ6dMIsYssLLk
KmT3jhZ5ZopyvHE0SqEZgsjIodPlRavfbzW5A1YcPNGiM65n9LZdOqglZf2Hegj7
n3raRYqNr5s668FqLhYC1NOW8iLJC/7475U21mUKF95r5y49YDEeavukR6/kZ3hK
Gr4i+Px/LdIIfyH3PAR56QZ3gIECVgIwb/oR31vxwf8A49ole63Pu6S8gmXzThje
FYcjvwKesaprKGfLbWTpQ8PxwgCb8/tyuxKrD3BHkRml2r0IlliH7zdKlD2QPXKH
mjPPQbNYdRa3KwNFtrwLf61DMoKClNF8rx/rZ2uNf2f2wvhoMes6BHNabhWFUmAR
cdBufAiC2RlmHNyCofN3U37qX32mDNHNKeYYhzc7nxkGLK2/517k5KXLppxUBzYZ
7uCJNjLTSXF6heeJrWCS3D9YiCPRz5a3tF1VZRS0YcC60+7kESp/QALNpTQMye/z
477Hs3k9F2woWL8FF6kgoxmDywYZVkpeE+8n9MlH1fFjxvbSy0kGqgXv2TwXmnwG
EgilrALYdlNqtsG6+dNqeC12WUeAZP4mtTfNmBWoqrhHMTIDn/hgqhFZYp/cCq9V
DQzgfzEsPQkA0XBgnSYGnBEJm/OFXF10oN7gFpxrMbHPiY0awfIAvTY9nW60ACPj
1V0xBlJ1skbh3H+s1XHUhMnNtAr7UwquqZV5noWLRZCmm+NQxLmjNum59gyZJaBK
zpg5RpB4vHdAIijFcBLa5yKJM5EkdK84XsWzmRzyeztb83pz+7SmlNej60YK8GIN
NlAFcvKDQpTP0FG/WuIi6BX4zhlbtqfvs85MJZBG6rJs8nYkmY3RvMAnR2CrerJb
mMAkLVon4zenNm2pI257VPxlLij/C7C6hjwU25uyVP3i+5CawwBqbJGzF9e6uSjw
CduH2V+hWPN23VNwgnGA546R0F+dDl/BpxVRn8lYUYMQmtUW4pOwo8KEMqTg4M+3
L8wOrBIGKZth3F2hsqcCJktT5eEjZkFDoQUp0Po61c6Yi8XX95Rj0MI1sDFhUwm3
yW7nDDzhQoEQWpFkx3DKK/3LrHK5P3xx0LPaqm68+rOu4sWY/7j6GYeTHtNwGdG+
hGcZvy0f+nPkcekpjJx/Q0+Nq9WIk7iXbGnFilZXGqkM3K62dkvioJBaFpY9MFIk
FJ3T1UTOxaLDKRwbpNb05t986abt/vQpH4S4lkuBp2Ll/TGmj6kxGwayQEe1FPXa
ibTAbLBtr0FTS9wiTpwqcrqHfMtpxuIQ2M4kBYYx1lfKVjdt523eQS2Stpn/CMuS
diU12IUA0EdKpxJfPmE+fnu52M1yNZmWDOpsx1w7AXvxKSaECe6uM2MPk2dn8wNo
ClypCypn7CoCWkOUEehMeF21t3AmS9JjECzNtZkLXkAhltpjcn0uLXzpIvR5gYuG
fj4/PBB/LYXjSPagOzQmh6y9onluqUM2zPte0amf+cU/1g8cpUbJq5lCqEDAQffi
JSLE67Y0yEruX2HwBvvVmTP8qKtZPzEVsS/G861BvjHxcyM3ePmzNQGwAcr+Giaq
hGmEB0AvnpBQOYfKCyo4Pbaplaw0BAcAR20bx0+QLzvqJ4696iPgrgrthkL0Ocuh
FiNWYcPtfsR5bx+UYcTPdUxKp1AUsQbcz8VSidQqiYPpEyw6CAINv3O5VF3o6/ZA
E1G4SLZHamBui/s4rcpaOvAVCGF6NTmdgTiefa15HsSpUtAR2CrrrTGv9Yh6gm7q
vEP5fSSCeIG2mukCtU4nUvlM7sRT7vjgJiXd6rAlW/Hv0MoP06WLIY27v2hq+lG7
dxPBUYiVLzbUa6dOJDPKcYJ0ZXKii66OJfHMyE3u1HrYgI0dBx1oZF+GOwvrCRMH
hW7Ss9tnPR9ODkUcj/8IAxbMMwzWEfeT1TzSez1GNgdYdR/r9eDSBez7OyZAc9bW
VsMFXcCj6rwfk9qXpUsHYWaU/0LUPy6q76ycvcPuRl0VybMPy81hdy31wvPuNlzS
kLd7q4fwlRwrLMwBdjSz6HRyS9YRHT/qL+jpoU0Ktnvn1rovtvUYh2YXC7dfbiZh
PoUvk4gHdI400mcRdroCj8H6+fQKGDS+5mEaGGH5q/BPjWBBnG2lc9BolMUR9hu4
Oq02+KZGMattpaA5r8PysgpCWmctfhBaslcmiMpMSkb/QzdZaJuhf2Tf38XWmzQm
OeacWt0tlvLZgDAeyQkQUmkZ9+zOz+aV8Pl6EirJb6NhSThwtJpTDvB9mi8UfHRE
dzO31mNsX3jiHpx1wSMKx8Dza+eaSIiKh41ic3oljN0GURhAeEB6yGdu6OvQF5OM
YfjVe9Xnd72FSlKJIGwTGh+9jXYRqaWfEOBuzwEaInQD6bM7QkR2dMrWu0iNxs4r
ptp2PB6UNKBFdnVswjgCY74HEwNF50KjgexDd9pZLeGGcEaA8rsQvvY1L/1F4LhM
J9vtAWldK95xQ5mEjl64jDJiSNT2Jcc2vp2kVXsYcwHpMBrdZxCwwHNF1m4jD4f5
zE1HNo83gwGD6k6kNL9vcg3ycli4fKkaMAJWLrWMlkKuo7RMdXtaQKcIVpqBMbv6
mKx+n02P6/anltgK3FQrb1rxH9Oc2cPziensZmc74uYuLonCAk5uv83IcTvvyPsf
Nhfz53knbFvaLL+/HYtmkOyGnwvKNsa3agR34ncrztorfoId/8I8+CxY5q+3U+A7
VPJwPR8xHk8njjWGM+iBO3RKnU+WBLZmBUDvzG0DdwRxq7jgxelv6RF9bqYxqVnc
RLn64ZvfuXhw1XRFfSzlesMOmA8uybQOmW1Kfb2u95M9c93mvf+MEAV5vkl+rxIv
+o1c10TspDxdpcKz4bXbeDOJLlJwnRQLrnoWDCv6ftXO1KXI5oGjRAGRwPRBXJjd
Nn+QpM6ZhCcHcgrEdmhIorz7AK/lKDvRLOrxCZB4jVADIFWwrG2IUZHgoYSYAi6o
uyWVeepTc5796EX1kU0CsljUMXht2wYOoLgHVHxNzQ2dI9Fu5osI7kZywxqPe00Y
a9kKKZ6AdpavQDNb4kmVRcwPHL0+A6wzlrWoVOnKkutzxDXsBgCP9okiU+Swq5On
TFXIfPIqcbYCIxCSkqJjhuDoNxuVnybAMzgwJN7EW6CPKQerNeSwSDedCfKMZYDx
Nuf14tVS57Q79s1wiS8b99SpK5CBLwW73uY+FGyaL+VVTG5CG972luoKLV4+5AwI
hQYW98sHAgvNHTivPvzcMRXdWrePtCUp/PPz9OGkZB5b3VBFQTf9kIL2gzxQVj1i
lZPXJMtaZiyixhs1oVtrrxYF0zQXMxqMhyuX7F2cRs9HfL7zh4vzRM3U8tYWUBiV
C9+deRMBozQWmv4svUDKU6SjG0Ftt1w/gwmiWKjn3hupj84RsEyiwp4E7RW/ufeW
k9rBoVc9Ja9cghfB4rUOmCacyQIijcR8eYul/AykVfGYs7DAcDD7EbBEC5mWqez9
ND+KYYb8jdD/V4grvSRz7TftYVnBtYh3tcOX6C47VLBAZDsmgWy0hme8vVrjy5Ss
MfmgW6jjPwickv65HvBsuZXB00JnsPizDuWmCmbp50iz/hTylB8Alp+FnBNyGHWh
t/MpGZhnWDU/PHMbzxhP2QOL2JbCa2j6jkMGmWn8dmGIWtcGjMIVBw0ioDeNpxHT
ymFVz/o1IWmjVmDiIhcnwByiKkS/NP4q1NRjsRnf21PGm9IJSA09KV6HMWIc5uBm
yqDqPCFAmbOphz4lBLRK+ilvcbXmwNypE0d5GMOZ7VMHO9Ho+nzoU0YcGXYuowss
K6z1MsL0QQlJlsjmsveJzdj4B7qedn98rzBQcInWXOD113xb57Wrhm0SogKH1I8S
zOls5it0z9adIYvaHYSaqEqKFZ2CJMuPehBnRpCTLRHkBEzzJToJCMt05m6vuSIu
ddzoRKwvjvszOCWSTGwGVFdzPVAY0RhQbd7AJTYuxXdv6VQ2JYmXouMHKlBuUbIm
11ldPmTNcQRpHuIHLSPZn2yBn+AmZMu3kZZJlZhhs5Ly55+c9yYdz9Q9R0fl8VVm
MucXhzwijRY2reVisDvg+irvTzhohStCaDotI87DBq0dDLb4vosIFjbhnBE8iJcZ
fih1M0YHcTIrPzZ6HobqsbdBPhOptpULyCqWcYyCpdlfjPJSf7kHWLte5pNKNZpk
PaFmpRU7ixUuuf/DrsWPdJNI1BhrbfJPBi/6ewMNmGuATx6jxu3vKwlLTQihHnp0
YzjmDZEWr51nNG6fqtQJoUDLq7+7D1ioCyQxH8RAIzsA/Y6RngpCRx3ynqIqXrrg
iof89kAZ8fyXx7+ulSCbSzwkUN0/pVX9hkt3wm4YfC3vcu0YW6aCwjNYtFa38kCh
NZnE1w4hnKOMSoEmdS0yJ/RVLNYEuUzpyhilmxiDmnOPFLvUdYUbqY8cq7KTCnOB
aFN+3PwCkC4yjEGWoY3VyqhORXwFt77x0PZqPd6vtdNypaxXxR0UTHbh23CiQNhN
OPrcbMRu6MtOpi1ePKQ7daYhrR3oWeIG6gbP0CVXXuK+jKpR9nLV5noWlwS+S6Za
D7qfzu8Edag+EQY+/AA0povlqi5HZgW3udspll8jdswtJzn3RBqeYfyaE2wQKiLW
dPTiOT7Rgb8E7Ir6g2Cz0xsS8tgv8Rtnz17jRhSC74NbQ4Sy3gB0S5uEvtJiGnFx
ViFSTk77UQw4eybeaMvNOTt+Bq8rMSelAkJtLf3JXOIJxo4DAwjDZTTNkG/Zo1Sf
ACtLflgB7L1JsaRigrvMFHMTdg142Vsk41OPkfkGcOv2vN4gw8KQW3bLokuCNvHU
kxiQF8OttazVZZ16aWAVxWB5I1qOIE34H/iMHNUVvuhdZXH7diqePc5FLpvnhmSO
RoieMzOnrlOI45y/gIEakpCAcEt0as+7G4pUIiAg7kYBj6Hb9Myitg0FGSyjAzDR
zuNIxxkEGpTh4QgEqNhrq+ohQ2IpAzNeVmwXeV2qoq1xFjNZKtsudRxlotTprUWb
TRa1+EBVfhTNlVspVBGNJgyMNJ73IjD60M0UzAAcw4ggIVQvyonFUCkI1q8AqvYZ
v5/4Xau+oFbct6wVZ2O0TgFD3qwoaffM6od48TnJeXFIMVy6+3ICXIzL0NaUQYAd
HhldoRL+GCQejDx+GE5xvLfSkwbqxRM2QgJZjDw7p9B8eAGINwrAWVcBrziOCbBq
0vf8d7R8fTB3h2b5Udv4cKil+A6ZDWPQJjoWeV8AHwqXAKNhGTM0zFvPZUDcX2D9
ocVh09W2SK4IQFqSybRAXD60YOMHBpOx4zPKVO95fyYQbTnEh0l9huewBNiSjVbg
jnc6t7cs1tdYco5NzA5R9Y56hKjFPPt55xgXXNxJ5mLI6iUoLpUM28Bb7sweSlKZ
+A4hQlkBj9Oz0g34kxM3OZ8tc5AhymnNhBQFrMPluO/GTrfIrev1gwzXL/SZnMJb
d7Nh3kkdPgWyEESWQMsS+6haEp9dQ0apbMlwSPEnfPccEmjtVWDDk4xj+UHkSMi9
tMvKEc+Zk4H4ZOSGSoIbKLFi+nAqXHzMp0DFtW4Di/hMVywABIqUJGCm4vqDnv5h
Gg6lUtKUiQck4SdEgBjWyoK9nXyxbnzygXZpv6WVVuI2IlZzpMS51zB6UhDaAKwO
q2tT/6XjVebB+Ry7O3rpQATD5sw5S0zs6rocXvT0q+yZfZuiKzRPWsSycn1enrD0
byZzcKVOSKzAMLOVfCTUJw==
`pragma protect end_protected
