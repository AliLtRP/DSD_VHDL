// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AfUZX2ECh1RZvRUVn7GZGG4c9L9qDHYqueiBIO/qHYNSl2hZJw+t7fW82hpIJodp
/Oa7vGQGxZqU21heGT7AoEwaldkwnzzx7zAXzqEzeE600Vrx9Md3P4Ya/TWSnFQQ
oQnZqbt5Hh6e0YHiOhispsnYx8nJklXLO2Lx34bvWrc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
Q/gLe3OpLfudIyckFblsZiGePI6AhQ76fD69B0C4J9PuxMoBlrTPjyIF6yf/1T7x
TQ1OEc0KsTcZ4l1Osh1UtTaDFrvBjEU052ncnjTJNSL1iXPaME6KZHrbxEDDb9+G
1VD+N5lLf6ZOeyl8uVgpzsEGT4vwZR+xVnGATFmkm2gLTnOZg3T+myY51Ug5xB2w
tKx4cbnD334I9tsfcGT1BbzRdFfk3blT+o2x6RXQdVpYGAD2WSzx7Ig/opQRvDM+
EwgWNPx9A4QwAsiKMVfwYCINbJ3Sjwg2+LmcnjHD5lWD6d0Zpz5y7+Dckmq07Uh1
v/GEg61e0CWyMSSyLkW0oMTLX3WkyxSn0B+uEtoHoY3BXEHWcFoMiCWBmXoFEUzT
5WJewng7mJBesa7vX5nnbPi6gh8jgsbR0sKyyjlQER+cRvDPg4MBX8LAKlHujGNe
rennjhBZXaMIT9yjq9J4njmTAOmM+mKZtTkfiBYD0ErfWk25LPv6mI/8uHF0S3RQ
aSdA4dsiUNZkmLbda91BEDsjI+vwqKGkxLxAPBVAGxaFkB/gmAKX+2FTesrsLxYK
tgvwWL+PHOdQn0r6S1cYB7uWWIt4UvJwobQoiaUfzOaKRqnH/Cn3L6qtEgPKUKwd
fJE8yJcaf5DE/yCa4Afvhjj6nO+1+BCKEzZDsx2j/emfqdJAR1+xnFoW3ZX4nCcs
cczz2ZxpiVisy9TZpKeVh4ONsHSqMnLg5AaL3vVnke1RY8j7txXYadsXMwDH5Yzr
w/4ER+FNTp9+NeXZdSKMeAXEYXGywO0KFullm+8IAGGzNSOnT6xRF9S/QlFhaWnA
3wqahlwzANLiB4WTVxd8FtFwX7Lcf1kpKFXMvi+mydVstpXFdkLRJvVTWhSSRYr1
7QlnTDrXTIq0VI9171PC7plR8vbwUNWnRhqs+ogXJBVh3KY2ikT2RnuW5HmWULTX
TzrO5nE0R9LpCKzoE1/tRwamSyRPD3kILGDqb48Y9f+xdYHS40hJZ/GLU9yKcxgg
Hch9+ZP14ri28nKqJnunzVPVBeCBpsSmMfw04EI0Xjsfr0LJpgznXHhk6UgATboP
mqJCRp68aTs5ER5Gyh1IBNts7mYUkMqlLKjprdgCiqq+zxn83oGo0MgMNq0ocMiP
4FpOFz2MbAmZ+aVh0jApQO95MSgWGximPfCNKSA+lEVuwHAjAqYjSChgTWVT8nZO
1Bwe2EsUx4dhuT+kfKhlqZFeRfXzHGLCFQ7Ch6Rn/XO+vQs6dyPQGx5St2iqyCtV
7t73iMghI9CkiS+biAMHWCBAKKssSn/m34EpxuqCRpUsjkATkseW3UoVI58jBMH5
i2ita3W3NGzWuJPL2GZ3Gbn5/UnLT6aecA1tJgJp82bAPcYt8A1mvumV6pJGmKKH
o51DfoeVU+B3vABrKZeZeg9AL2fcpMU4I+XE9o4y8hohnfVEnO1uXHgYw6iDcB6a
NdgrYIG6Hfsl5ob5omgGeviPnLmWoFWULjqTq102wOphGemEcJsjUg3FZ3FxxJuF
lLipFzbON+V5p7W6fmz5xptcwiRbcsOsb0r94fKm2390RLewRWLUv8TZS1APlpN4
KtoNWhBdmHsd8OT1mAKmGH/F9IGx5nQLWk8z8zueXKVUc8V0RBnIYBYcnezZRImV
QF7Ikm0PwgEQRSTemlDMI7sfsvhMCqzkCW6bbkHwz63QG0bGCWdy4UqoPOnScaMV
WpstCot1eir7erfUC292pSAFxQ0PmzFeWqHMcoNPlt5IZjkVmC2sJQAtNOnozJM5
LR/FOVFvWPcK7VB3a+lsV2FzrwgGQrJmrGIj0CGpvu+q9k84ORBJ4mZmSlPATP0O
mEUqASURtuJar3HAAbCxb6A2xAbrdwMtD/4L+38ovGWemHMMmiOpHucr/s5Px3+j
3jMYcqFt3ud8Q/KLsic8+41maXKaemB/IIWa1Fko6qFo7KDMff2qc/+tk+GaU4Ac
BvWIGYhTg+Qw68kInNc8S2qw2+RwWaioho1vW5cBm9VhLXYfhIZ8eKKZ+46tTwEs
Fh4b8G7NtoaRtR3mHF3QDmez9Wbr+vUcMy2k5hDaQvZyh27cFpDs3Nc9Nxh5L6lo
HTQkd/VTvJKMRU40poPuK4hPFl0aZtG4c6NPEtB2xos5B/O5cWfOKpk3SQcKioWL
ZMGwKMP66gPvYc0zRQPq90ujljc3NQGSsT8nHKyOcS81kVxvzEL1osEKFom9sRRw
21w0pKAojjVDf6hewiybaCbTCd9tDwPkdH8Blgq4y1NKVh99lERy+VlR3k/95Zrc
Cy+aZykDVtO05a3dkfC1HW7GFk0dBTlvNGhgiqH5TmsLMdZ5kKIfmUtJyDt8C+ta
BjwICcGIQCgAGklyoYwo4Y/B/1gnyFjxTjKf1TUYYRbAjSe9fzeFYMc9Cu+P4MG1
le0qa35gPey2M17A6FCESUYww0ErjyDh39nGTcS5Uihi62VVnX8qCSvqiflNltsh
3P8lO3z0WU4wNVU54CkbEBlCxUluO0SzzChjaDYuMvul8U85wkE1vh6Lb715bMby
Gh260hgPmpnQEm1n/sVw2VjrdZgZGx0uQ9bR69E7QBn2KVXdlMiP/GEHHRa+mQV+
TtrlRDhJ6E6/DW06iALgJTgenjg87sf/YZZM5vvKQOER7AzJDmA+RMpm0qCFYs+/
QYmiZixvNR58UqD4UxGzY2+qxEG4Mh0GcZPlVD/Uv0XMCJJoFpUvRFHvFAz/Addt
KEAZpzXgVGWfVKGwaNSeoT9flKfimhVet8274PuUZl9SHTqNjwefBKp/eX83/0Kb
BvsxDqJuPV5sUNQPB8SJ/4JDMMAkBBmf0Gi6FN5bqd73UAS90RMzuYgybruNbNN9
trejGNikR3RjyAxeWOau+sTKwKfsr+u4of7f428dhFrHjvf3VL5p3MGHTpv2iM0p
3+tL5B1Ue0JK56FDEb384vOpPkpQL+HoaHg13XbFdaHUR8tXDnf44Bgt5Exbtstp
YVvQRJ5xqQwk1XbnTglFf+zoEPvjA1zD+dIQRgM5Lfdir8yGAyvcO4oXtx2aQNpg
RSneoQoO5FMD/t54oqYkWRKEZQqSbz7H3/DYpKse96/pBpiRnNHwJfhXGXXGpHS7
qu2Ie/olU31Wggab5Q5L7k92BOYqAUZE78YNsmBGJlSV+CszQhPNGlUBRCpgtaHc
sF6bMChZ87/9mIMhewNkB55L9enxiPUs5ENaR4OpInBa7NANJBx+qLRy+raz6OlM
KbDitqyUlAeRdoTZ7svEFR5CnJWrHGE4iDGLaRPjqzVmAY2b9rM03VjySb5gAtcG
ZRhsM2lMgOUx+TdrjsbJtkWAsxoY2mvSjJ3ui+HxCed+Z5N6UJE7VaKF3C77uGsq
6wOLH/304ZfHeqYpGyjr1TBxbkXx1Rkwbx7Tmr3OBEJc/FH+tMwptR3PjT0QrHFb
6rfOI79U+2vBxCeu+dy8zmMrLC4UwNuRwIOqRTm6oGTGbYUEKpWfzCsmqJXc/a9e
TiwK3nNLZ9DbUqa4cKg5xdWX6n1Uk8dOsAP8P9rejTC904BgQ+nWT5fRs/3JgT6L
jXXqzLD2Fh1EE7EkorW54V9MrU2pG1VtYSmLNImFhNJbNy4A7JVin8b3RnSYyOVa
MkyABenVC6tRmczL84EyYi/LceFynMp3BIVAoLlMT1wt7U0MmH87UvwmF+/7qlsx
77SUj7ocN+gJSHl6La5P7iey9jJnVnqIVFTBpg3zOsplJH6yOR7UvL5YmIvLQsGj
E6ktkFkxMvjbQQS1TDw6RP4c82uGhCmlEhxgXyw9yjrvGlPW0D70s+2pE4fL5O04
XuBy4glcnOzLYHyOrNYlkZXoFiF1d3DlDVvkvtr/frewCm1wJYFNuRX08xrnkXQi
QgpbquB6rSVLh5DQsZbtixDeYCydjLX/OYMXWwnaGXlSU33O1sjZEQPHzojUBPtJ
7qjIJJtKE6wHfXkILFzSR+Xu6BaaNbJbumKS9mkiLdhtGZzUbT2VE912lE1GxaW2
nJcxOZg1xm55LgktYA/d2DNjk8QjCA0t5Mhp7I/4L405qjjs5uJf250fZviUK+X8
4kmePxBHrT91iuV1TVgWvWEWCwcoT6cNoavS0mIXIu8JyWnPUZXfZSO3nol5V1Zq
39ktxWW2SzJqwxXIaGQP1RpY7jWDrF/H2j2a13LROKjApN9VjHO3ytX9nVvuFXSV
pOXS3Bent/X0cQVP962unMYZNgxeCnAi3o8bhrtQeCpvlq5DpwOaKOqO1+EQ5YEi
7YIuJSj6WdREFItq6/rjIJV3QRyvJR+q26GDGYsaaXxn0vNZq/AiF4kvsuvuNCEh
JikfhZDn0gloCyg4S7iDglLXujis+5GPklSLEI0javLdRtSIKAS1dAcfBIphMdpR
5V7YBWEPAwRIluifGJqZn0677uP+K2k9KSxK3VjknIVjjUo/trO8LwI3xi2u4L/T
IMbET8pFHrjPylnWPLybubgI/rATWQF+pJFla+l4FekshhgtC21hnJDbcL4vpK1z
P2VKvqaNJ0VTuOPsSbJ0z1BvzPSGQmCK5IzK9YwospSybAhejf2nIJ0YyNM5W9T7
WWHbJRuZK1YnROzwFQMvDX6O4cSQw7HO1F6h/L3VuWjDHwSe83MN8Xfh4+Hd22c8
A1xFip0SyCxsp1i0fcarRsLnqjicqO6YhqU/7G9yETnOQMwUWwVHigcrahMb5wVD
2s3/kqwI3tbpz1cFC5xjpaesWm4otZujlEXrkJ3p8LrArxV9ufTjZ9BkCsv28psf
rpq8d1NpFG2gFDjy/+dB9ek/GPZKe21BnKhjXvVdxQgcgv8FdflUCJTTR+6KfaJS
28ina+osF/yziYSChwI+xPL2a/qsRPFVBPmrr//JOfP6UCIIqr3XZaswNgH5AITd
neopnVX+zSbo66BO9YBTfP4BLnd6Wz4nLUWMwPxg6OtJOB8bj3+fxLDXuGB8RkV5
VPHb0ngwVIQih7HeqjBY7cecA40Dim/ZYj0E+S2+xG8ZEGRSLDVVDhmoPqbCIIF1
kwXMMhjUC4H5YQ9XqzPtt4s5sRM6HlGyimwx9KMT1PRy5CldlkWdL+ZvmO+vAemB
N/mncg+dmgPOCSfmKbq7qyLGDVBUSfQyPYbk54tzx+o6coOjGc0e8g8AFoyKQhTR
/3bqQbFyMr2rno2wlfa4yEaQDxPshR3v+je1UM5z5ogV/f4czK5lH6IoML9j/SwF
sEY/MeNm1LeBQ8xXdHX1c1617kYHJmD2Pe3BotK2tpH1wHV+Eg0TZ9YQskrn+uZp
EuHjEEkISYkgJ8ZRIlp8uQSkKbEakerNeG4qlSFr3yb4rs2g1+gEtfYs9J1bZ2bm
4HN3j2YTPmEsa7FS8Ln/lTjw3YgwQe9u02E+WsZP8kT5CMioyY2hLqZnjnqqoFtq
uyeUPCIa+/wI0VgH78O6tOSKlzQ+hie+uzEAUtO3OhBkJstWeJIbNac1EcVfYQBT
wPF9uhFMw+jup3rYDo4vRWYlQ9Pv0Dem3BOTIqtDVUpfL/ytBTDaUwRd+XiZs2RQ
SSHjPOBLdL2CZoRLWicfE6FgGUFSPF7JhtCcouzT2hP2aJMDPMjXzvv/ogSep0YH
B7JYrbqo4fPlhyz+VTo0W/vDe6ZTfdJntfQb4R7XV673CGmlFWiNbKxKB9cN78fC
dzs6JWLjeGRYOfccD3zdrTO/FoNLP4Egbfa7Ni+JGGZyU12A91k0eMhTxqd2+nqE
v9S9yY4FePK3cPOsDhlq0PwlZcJ/C62M3GB+qfX5auMa6pQ1i+AUfTzTYXRiv1lW
R4RjVeRUI44FdBpz/syooVIXqB0MzSDFIQ5INonKximsTa8lJuIygwrTp/4q0B7T
TdLqetlC8/uWVS1SgsAlWf+U6uEAVPaLnqHvdARZtQPIrLCiEWaYXQhN3CAjHA5T
fJHav7saJ+Av1RxOF0IMdFYXn2tY3Xr/R0GJlOUAzAPfbv/8hOQYEmDKRmzlNAf4
7iC6KvR4lNSL01B2aK0BBqkHBW9wk+mOycpnd/tj4sRgRHEnuiRYINEe7Kcd1ryA
uKgvEhiZY/IiIX/qPUvoC0zJ0QlQC+cSSKSzuHS83NnrqezACU/cyn+5/d8WobSR
yah5LMN8sxE2rJZs/fYjC79sJQkK3AF8ox5cnj8HOm64BMeFtBIDG/76RhEKPjZF
ZSJAqbf1S3z3hpf4mxv4umIhfKO09VZnNqbwUYxSttgUBCGuSSqPZ3dZvy0RsHh1
iDgCXEOg/ovqcGsQH5F1rkvy9R1Tk/EU4vU9LvTVUBI6/nvAemy2F4ubbBz/cGp1
/I7k2wRwp6PfwTkrM5t/9qK3HKx6kZVXpEMgtJ1qLCN5USuSzFhZ5XmK+R1/Gel4
Jg4ta2semDx1AFsSIg3KUL4L1MAUReiPDcpaTVcHEYI0CEppMY91B3cdmRP2NVNs
WOXg8jHecqb5VyGC+O/0sKPY3I6F6zMXhAo0RwAmDlIF3JBJWk6WvxHy+Iq7N7D5
VcwV03MOSacousXaR9XaQjfVDK10Fed7L/4Fgb5NkqRB/jRysSU0NT/h1LQfz7vg
1uP9Q6n2SzTbhcRlQ5ZYolFggM6B6W4TFZ3j0CCq09glrSQ7b0Rv3cGEpqzXREpU
QgYnn0pz+WnHpAyYZ7AJVy/RwkCfMZASNcT6G6+yneVfA3lbxLFQtfdyhcv4yrQX
xA+Pev62CwENvNe01Q2Lt+hG8OIOhd0VTrV/Rpa5OErZcJKZ3aNLt7XuUFIhfkb7
WCSM23OhtfGa5rRfxj71nRK5davfTY5W7hdx5+bu1vL83/OgRhrjgU/eKBvWNeIS
dT8SdlB7sHvBYeL/WJh9IdYv5Vvr0aadWMnFbaUWYAu/GztPKrTswCLmjkdM6vVz
vH6SgcAVQUoSVP6SdtewaqO3Lb5Ftc/njUdWgEwGnUQSRp/iBf80Ntii3gUZ4PCE
W+otHrVgvZQgY90y9SBR0WRB4624qaGDWJFYzO9++jRlqB7XOBpS8EVLt7+XNqNb
tAbyzF8Da0tHbhWb8XSWwk4gX/2DTcsCbhf4IIBkHutg1dJAKMr+xpWo/tEmmG/Y
mIJLMQg909M8fQOmxFKeEF07p5YvW3xjE2SDNhMzIHnjM3m0he8ecICGEE7YYbzi
dspfRzicN61ZJZgIUOMfuByoPk5U7qzpcRNT5NJznhhoaVUue55YusLj7cZeomkf
NCQWroiQKILXuBhtfSe/E/t5CsM1zZDgvDzWWXzBQmNo8VD/UvWoeP2izs0LphOo
q7Uok6+M08V0ztxYpcANh1gYwCewSVRACpjjgoOG+aaXnLvNSyuq/GiJrHGOimDr
rW1E2PDdjemOUJqEz5aZJQ2/MvMZgxfYy+k9mBF1GreRzNwbMrV9eiji2O/3Dhs5
bHnaPtZ0QZJvDWWViq8NLA==
`pragma protect end_protected
