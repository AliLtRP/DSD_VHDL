// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ManmcuQtzH+KoJtDJ2TrQ27lHrzBCh5tWvPNF5J8MOIeVXt/O/3nDt7hGCcogFBg
pxTBeFIcXtbVmZwvNXYyStcovsmy0z1FRLbZuHeuZpL4a0wGEsdsfD6CRXGzmFQz
oqfC9HphkaFHCLatY5bM8/8vCMr01HBWNuvb4CCFbAI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6384)
JeaVp5GXeEpXHboa4/76g30Y5Z2z1KqJZ6mrDbu0g57mvOz0zPUJyMNpFuj/BrHS
3SLOfsebeWYIIUDMZ2ystIruKKaOmjFKUP1rmclIN6vnEZdBUTKRVshoi7CLHA7w
ThFL4oAt89Iz3suX9E9ej0C4S7//iqM7WRB1UrWw4yS9Vw6i+AJH1kqoNUlRrCMS
5NqCS5bnSlGQKS3N+apD1SMRE7Hjb7pFwat7kk5w4Zwgv8oAtwCIIzl0E6KsGb19
PrqS1IbILO4GmDH2RWajVE6I2ln/cT7fn1E/gBcBy2O9S+7I0+7mnrp6o88e2lVK
bIbfcEYwnfBSrkfIB2fSKj5NuZwQtWSwczj9TYrvX/XDRbkgm9edUgIlub+YcBAg
VDWZHIYwNNMszHJrZdQxepcpSvO8VcolqJ9FLsXRr+I0BA9gQVcMdD9WML+qcRAB
D9icOCGLDo680QL5Cq5liFspiFqI0kA8NuQFtiBg71YWpaPTpNI4PwansAG9wEtG
zwyL9s8gEsLAG8hTsbmU5dKsxUg2c3Xpa57n3Egd339zVVHjdlgixrh5Z89xcSiB
hnteRACEyGjaScfVS2d7MUetbQoK4tI1KQ6yBvFu32lD/nuHC4nMh5t4ES+92Laz
8sTrOBRhXUDlu3XXahHosxGhvnrU4nEQor/NvUS/dPj8qva56wW7QL+TWvJ8Xw/t
G6prtjsaB6zK7XQZjKdHE5PqxqloJ4IrEN4Ebs8KEh+8dTbfQbv4OfkZefk/jMA0
W94uJE4ARmSWR0wR0e9V1iFCxMKk1Q2bq707gyHsk1usp221jOi8QAdePPb4hSWd
5HFrxcdlSPOKVjc/Ck+eq68GxLHQF01J4XygZDZWdhsC9QqPkW86xgc97YILXGUT
+eRBpysp15Vc5UM7a8s3YYtsw7PQvZa73mIllXNeZ5z5kcQlyjn3f06bcYmoAABW
VmVclDfmmfzyYH99wBldKOuxHVQauAsf7JVbKhHZArlNK5Hlzph3FMU/dBOax/ba
3mm/df1JZM3Qs+vxbrb3VpQ72f9XcR5FlwbFQxf/hWj6c4r+1RpUGYyCCiRiGMGa
OK+yEWJa+FMdEsz4dtJVObqMjBziOOS7k9N0FkhVF0pce2Si+We1OUdZlrNb2U17
YRzLwIbZ8BvhjXF6Bq26Yo+TNT3VTMWVae0AySCnZ4WU6ZpNqW5RmOEwBNoO91a1
ZYVfRtxOapZKvWb71SqrvdCkoW2+vfLX6Eu2zF8CpTlOlEzgd6iYgI5Qu23+dUI6
34wfzfmVsvEGdX21nrz+s5DSHev2nkRRljBX1Sk+XAg+02jzbf/0njmJkFqcAq82
JKnCR4K2g7JkdgRnAwO5U9KiPw2+3ZmY3e1soODoUAsl7c4GjyPG5DDganOLx31d
3mE3FM9730dyfQ6p99A4x7zRs4EPf/nzwkxKMVTQjyBbd/lVh4Y9hnNcBD/W7yfj
/9u98M5e/gzX3w4vFRoOCu3ulYdU6sZyR/MwsY8IroHGG4HoNsBoTlYqn7XyT5fJ
YiGp9U5Qs/c2Dslxzc4FubwRqijbgFyDCxb3aoeU4PFPnV1A2Fy1MtaE3s5wTTM+
ax9WGdMXJFW4zVKUKCxCbk6MsLaBGmMZtHeYwq2gunYd0uIHR5CsNW/64voQJD+j
0SaUpJG3TBrfw+mqq3KRMEtv/HU7XHT+Q110AcaWN+DrEf99iKwUNm6Yho9k+1+f
/pMuOWzxO8C6sq/FkOTo5I+JtuYq6MA9mb48KC/BbKUXnlOLO/CZMuhlvVgObIZw
Rqj8jljlyXWdB3n50f5jPRFkkgF/QmH0gpBl9/6RGAqfETzKmNtTxQcIvIrO4ntQ
cVz/0wCBNpY7KzNQHcLgHGjxczt/ttDDyU4vrlG663AJB64gNv9BHjH821OnsoN+
VXKyZ2J570SVucGrxsOn2lLRtvztrNIYvmkWjj/xqYdi7bKdGSabA5BRvrSdPZCs
FdVfYfn7gHJ4I5hp03/SjX9OYq8ODSt+Muq60V4xrsTDrfyPL6MfgPPrDlDh/mnc
jSW31hUzxHnM0t3+13DC4BYQqlrNN+qU36w6fK5ObpFmRAF1TmGay2IUQALtT3eu
dPeq635gFeTZqCIlSnb3r7kI6zZljXyetgED1dsr+kOHdY6jPNn7NQxfSjWM3T+V
JeokMuKwIm2uQNFCacTjDYawAToZJBY7xRsxa0rGFi0z0qQ1k2qEhRAi3j53ja5t
MizShe2KS59M75NEzNDMua6pIdAAXBcvM7Q150SD3xw6wknRIJxUnJ4OXWe2sP25
QtUUqgLid8dagcOljCqadkMdeOvh59HdA3wEJEjaxeWq21ReEcCt/KGutkiY7fgY
X9ysAkG0XLfvdZv7cEibZ6UwyBNxIo6wyAACOmHxvN1l/aCe91GF/0KifgJb849X
SVQAjcuL71CWO1Efw0YFCaBvWGwO3xqJb0WffzW2p31cCRXuvDm+6FDF0yLoAtfa
0ZlCCWZihLQuaOMZNLLSyk/bSRxmF45L27hGiFqgwBv7MHMJla4MUtN9av508/xB
aeFmnCuyFwdhJ5lS9UiXFKpO9T4qj9XIKYzsauFELTxS2nDyBUoSI6xpTcncgAI5
nAZhVGO1P7L8DijbbSAv5Iv5/ukMEWT6WRufRY8nzuAliCW084oYTV0FBZjHHbVx
0mSfS62M5BkJPAYQis2j5hz1jkScUyoz06EhjWKEFoaLMQHPnV1zyCj4p66FqHHT
Sqz6Th51kYRfiRXoPqfYEQUqYbiqyWoTxGzkvgrc2Nojwl9gFcF61LsJ6M1cfxE3
UFrTK5aGuixuzQktF295SIzPlARQ8bwPli+10hkfz1BR7mbjhAOkkfhVkDwf2S9/
pYLzqyV3ugyrUdQzq8J3ozT3Sak2JBXOVCr+XTcCs9jsJICAii2RY25pxqPoTtW5
8EpByKpU6aryNleLhsPM918kvEDa/o8Tczq2OQgFduIDHGPidxo6tEAKtEF3YrpM
UUyKyTuQMFhLTyM657irPV/6IPW1gPc+XY6V4qx7KlimS9u9H7msvgJohDDWmRVE
qFkvAEQYXAuRK4E/n/sLGwowcQNnn2F/AzZYZ10mZmD2FTGZE79/p1+nFqdMjSgg
xEtegs7EXig1rl++Vih9F0A5pahAJ4vC7NjBo/0HSl63HhgCyLeRPFvK76+XLF6g
d3y6PvIL4KQe3zEKzuBgFWk9Jg9d2kMPfQytitEqe1QXwlHIhKQIp5saSgsoi7/l
SfJuDl3QfxTciqC5gSu0YAV7gswpPyMRR7kZV5NQNGD2pjlrCplPXv/xHGvdYwTT
0QbbWw4JNErRp2Dn6+Tz2aasudW6P5D0Ar8LIR7heGXt9p5iq+rCRaL4eWXyh2SC
tQduxQdRDQKNj+kE1z8ukA2XU7uTkmAZtZ67++UGPGt+hDltVzUzhyhzLXgTaA80
p7F7VxWDYyOG53LAoaFh2CYbNuBywshJFY3y0jvDuJkHPfN21TVwFmZy+2Nc8BP7
W5VE7BvYXwB4QfpwexIOVK7GezbL3T7lDPowrcxMWyYfDhj3jXAqQs0ploVRaM2I
c42cvZN2pGPZd0RaLX9bxEr1m5uy/D/1OQEcljkRBMEYvWNEmNzBIYdY3NHqjq4q
J9z9OdmEEF8Aha9x6iVm78JXBrJr1EQs2UcX4fK1JP0UO9V/qNFMRIzsqKeoI60e
s1gDNKbGHdT3gHcyJhKENG37x5gBC+mYC73YaGtC85EBpckjABWK0XGVOYAzzsCd
6iwiCcpDCh/UAZqgZ0j+bZJzVhBx1AiSBvTBO1m0SdTcvBAZMrHeZ8wVr8NH3Uyy
yx3Qo5rJe70YQDMeWA4iIr9BBiNgzn5xq58U/3xUj/wOb4gx4L5TsNjfpmlqVzwx
SNGsPPBSuD3G3MbbQNf2k0Tj/BvZhne872adUGPXeL9CyLB1LBl4iNH8RWLkkkRs
NlhcKmxeo78y9DL+i5KELnOwRHNBFRPhyeoVslWH86NHChQq1ejsW3KBGY39VBAN
MQvmk31588Mj/aIH08/t737linxwlTlBRptWDr2O4AZxR3pY44TT5+0O+qeR1RcK
wwbK0AKsRl0DRyYPzraIvKZ/I4/iY3dglMMrOgYrWbf9L11n1VaZvS8SXQBeE08p
cbDzEV8I+LaJRoTWrXB7HUNm55t3e0q7fIz8Rk1onhvu1YrPncYTyE7WNdZZl8mr
QhdEBfGrEPh6IUesLoSLYldWl/Yzb/cNXVML1j2Cu0FEqg2aKFHJUg6N8i0aOdx6
xYvdSF4Rouoh5pDOP3NTcw3+sU+yE+7gxh6a1OA9XFKSTgNhK1BrQdMUBTG1jL5l
V8yactMZayUPU+YCQpRqYAaacE084+7ic4SUkHfcdJCVBHcILlI6F0laoSaKj4W8
zpI+VVHtPRCEthjtpeNsjAWg4Ok/wjbnrKJIXGapLNllkVlZ21BeY6gVC0afym5k
+iwklu2TpYiSP25uVmovUULGn+t4xfINtZC3ErNc/uKtXbGjnT8metjEH/+C48yR
ae7mbMwzbLu84q+Mkfj//liH4gK5JxOT3kF+YWNFh0vzhATk31n79vM6e+A0fMU5
zyXnKnyF/NRjH+vzGHXEdMU5wDnXOis9A5MGusdRHyI0VzKOK6KhyWDcKnp+cXLJ
2FVChe+fiWQtRGFUkolI4xYk6uLvsMoSFrX7ZK+9NnQWt5az1iCg5TsqH9R+95uh
5h5GWRJEe+k9zVdzW36C8vFngb2yEVARtgAw2/mHsPl0XWBOpkYT4V3Hdq2psWb3
d1UzvzuTBLRN9UJCBeIndxaoQsoQlqOM2t74c3uiQ/OOZR638uQyMyYB1mmHRcpI
ufXsXVyvW9Dzdfdph18WVw/HClfrDZY1zhwKHTlaZvxnNOa1LF++Fqnm6D5OPNpb
4Ty+VhPH6cgGs0uF/lJATSTSney7AorcLGICm+zue6folLaGCt2Xks5pvc0YE8Pb
1JA648isH8Z/wglP6pY7b+aQYF4O4VIHmgccIhUAUpoumloA743WByCW3zw+kWmq
S1rBP78BDNp071Uc4ac7Oemn+AS51Tuv2NRTHku7iSlt+DnKMVm1mp5x83YpzXge
kJ6ZRXg2T/QJ+Ont9K5ob6sz9Xn7AlYAA/qPIj3/ZDMw7yRVwjCKz4/25wum0v5w
brqwh1W9JXl0y1p3Iljbp1hvSUfZmHKiihHXlk7MC0PypXu+1EtDo1xyWPzb8hE/
MQqa1j1n/9q98HZM3iSQ4SYCI48qaVrjlrTfJPZkjXkPU0lktOxLZOK11hhJeZbZ
RqnEcY+ZRXjZ4rHI9Y7yDUXrV0ZYr9DKzer1Xmz5V2rs1pyNyV1TpQxie8XksT4W
WguVwpWELd1I/Uwlx+XqvEdpu9HbfEqjFgH2nLjq0c5lGrEyKxlPrCd2Zw/8W5FV
3Z1W+Q/huJ+90wVi9qmz7ALaeonEfXDohUEAiKjdCkXf2g7lwGserLx2PrzspRX9
hrY+nYVOcQ57MSuvni7d9ttHIzRoHKv5UkZ4O+ya75jQxxHaCE68RXYOpOz+Khf/
9KNMbAoLzXevHn1HtBeY3SeOtU4wL2ayaBEx01yPzFO//X3kGmY0BXlCMlJotPwA
lUOkO1ALYyS7zXKRIB3ZGBjBOXP5uB5GRvRQARiBX8f9/fjIzH4Ou2ZFlyOR9EGA
3DYNvFOt8/NjnG5sAc0d55p7OuKKNFToaqmCjx1PYhlqOHY48UkFjrd9ZE9reRDX
0WRBuoKJQ+WzJwbMPFHE67gGSnOKyjZ8lPLPxxlF5pCLRW7owetufY+fd0d/2F8y
c+cUl9ubDQuxSUtJm/nx4dZ7CRu9/6TulCTpqHS7bRvaSDdofVNx2uAxHp2QzUi0
G25/RbKVh4Rm96rhuPd9CkP/68fidbQFa9nw/HVLZKeAOxofKXPCbkPFi8jCO17f
CMxO2wAAKiTlvQFwC6TPEg5bZWT3eWM8KpQZGAV8j3Umms4IJw/qlHvMihPv+ORZ
mtDaHzTi6yxDCT3ibXfBlwcZoQM6YPIGJN20VLzQgjbOvApg+pCbh0ssnftKZmuu
kHS3yxHB9tFjon/5/cpxg9MxPCCIDk06o8F50KdnLrO4qpZDppplj2xbj8MvlUSr
cOd1T8cAHl6OE1VHQ+1ir6DMu/dt1nIuUhe8bBNkNrDCTTxJdXNFYrtm8cHHSAFO
6FnwU81217F+C5/xssr9uyIvZIbYY9EE1I+GYUdk+ZGJVF23j43wuxR8CDSnQNHP
0/GgvCtu/jR/uk+9DMQVL21UEQxrjMn4tO3Lv1JbhWw5dPp42m2o2efzJ/KrhnAi
mPIEYZS6FHAV/8ZSCkqmahhZKUAVonRuJt84UjvpaxQzxnNTw6ULNlZBkG79WBDe
fPjVoOL5zBberWkfC9TGwpurzt3oayqZmuUfixT5I87GvNdLg9904ua9yHoznDsa
U2IOEgc1dwGI63vjcM9IVyCRrs6GSlqAxBw5cL1iV9rZnER6gIvDE7ToXXCQETRE
MxOld0Y1JWRd+llFxKpr8DcqcFnWuAvsPo512A6ZBASZ7YPbZF6zyVW3lAZgomY5
+Iu8nmy2DtmYrhfwE6S9f6cbjyDIHgC4sfEDHdYQSrT0pffRhnOJ5ubZ3btuzOoV
oGE/XgOok1fLFL/hwamDkprNzTqb8942CaE+0ovk7YcosErICR32jD97cxr7+Bmr
SVZAxrHCNvjJVxYuaQk22cM/lhXk9nd2RRSmlrsmsU9L9iknhdRy5sMe1gBwdHdU
pgQs2HPTKt2jpKzTFvMQOdoQT1nJZaJuwsESp+35Ii3TOTsMWv1bXFB0T7I+Ojp9
Mg7u4fPUf8DxPMuJ8o9NoMXhu2+qH+zuByq8Sd3X0Vr3xI83GEK0tkmbAMr0VJ4O
vD/IeQV97ieAsDf1q8zw34OFOT6GH+88XQsQnVagJy9MhOjsLrlvWMzDgB9WDyIn
VrePx2iVNe8hm0TazzaEPoOKqR1ATmFsAgXKia1QgG666zYdwF4nQXd+ZP8ojInW
CwOTNJxYRnywrammiCULT84mMRZY/lCFym9/QXl6+Fo5/xwkdneNqL/Ko56Y1cq1
wCU1SdB+qxfEyMIQbBIf+AnLDOeiZkGfoLaqXY4PfgcMJh9ZITb/gZWPLbcmwXcP
KqagFC5MIct8Q27C1BJLB5+O+dSlzUvPh0jyURdzkd89fdaam8T/kf2LULunbYYi
Aril+oJwSOYpvMsDMnzSiPCCVXmWZPaUdDlppweILb8HT0UN+SP4KkryBS7oD0gw
iWfTyhrnAme3cx+TCXQ0304aqfgO9Bf3PchpmCp2LecF8laDxgdgmsM2flt1Baop
XSFIUjEf6mD49YtpMK2/bOHzZnuCF5Yckm8GaPSZf4Cf2Z7gIcMj8KHfTBi+ECxm
xfsnqtlo8osDey+cgKNKUVmvrgEkg5Zfso3wT0qFQfr5m84o0YmIa4hJ4Zf0OjIA
kYzhOmFCInMHgKLK7DATPZx2Am0G8HWF6JScqEgi/jIhxkICnlY7Uh1tmD0PhpLO
EREKow6H79bI0sGcPWMASUraEQtvV9cRjbvBWh77Qwyhjqxbvy03HObDjx4Nw4sa
bqQsdXZymGAsEO6AY4vioK3SYKaaowvYfvsP4upJ03IJjwbC19IclUwgR+TtyXbR
/OCU+FHNiR56o3cOL++NvX5W2mvAmTZqpkF+9NvL0gYHLswDvfx0xrbn2eyfF8W4
a7huSD7Y4r+os0HtuSEnZtBH0Nhcf4JDvd+b4n78jVwhhllpiq82gNoeDDnHwdIl
6a9hU5FCGEfaI/4+Kpj9a56BsGxFlViNCKzs24tMZWwoID8LUfa8FRDxW4BmStAu
mhjMYFeC4TNv9ptVKtxXglH2lg+JBlGJ1iJ7FAc+uYxr8bzNlREdFPOI7uFT5CVD
3P4OBV1hTVqw6oWQ522XQiUtvNEu93IyFd2+x4jW9NMEnkxNBkwb30oEw6XwiWYG
8nICzw+7xGGqgtHHKGY9qnZw2kInSw+EqMAc6s6WhUMPDUgvoOuaFOemL0S+4yce
HHevSkOyiCtpd8Jh7xWW9WUYKWXQO6TMnNAfO4M45yszNWCYL8uZB1iNpC3KEFys
xAH21dTb72j90XTnaIAlVTYS1wbi6mKdV3Gj2C2i+l3B44lVQl/R5Gnc8Z+aexmd
RpJEDmjgj+LEj/GXaNljLEbuA/n6R2ZFsw43sYOHR2dnoHyEK922vagnMM82vXtL
d6nEBiZRPgOQtSQjOYqic3ojVdi6gcyIXSCJEfdeVwTz+jgh5CHbM6BCsLbAiDcU
txEdfXuQf/oWmpT0u+1VpcKE03sR96YLyuPSjmW796pTsdaeOcXfrUeX2jFp7IS1
e4f6QVwQ7/SN1tgPMmQ+19qTYICcymphnuI09kKr53zQQMywIfAPHtBary5Fka/z
59qtnzZRfAXh47dXJGb/kb8ld5TVpZG8KvKPwhHscfDSHMzKkbTonO00n92qt2Gi
`pragma protect end_protected
