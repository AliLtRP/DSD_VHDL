// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NWVnlzL00mkHDA+Kmi3YWDzkJU9IMwouZBEosTl0VZ/NzC6twDY6yQt1KVGua73k
EQmWEQcTBGBoG6OElIjQc9dEyxSN2a8sBeJeCYnJCpW7bBd64q3i2LA4JUUYUbcX
zAUei8yErgd6WlTn4socO/qWNLAIZxN1ur0a3YE9a68=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4816)
F6iroMFEXZX+4QqPoWzyY6pHxwIA4A5RuIfKXa989smBzgi3v+UofWfHbMbuFd1E
GM+jrn3u88Sq+5wgZzfvVY6LEdInYZAOoImRnTJoGIaMxD0AyGsCWyZi2m5OQK1d
2dECnfS9kr27Bp/5/Do6sf+6FWT+nTyUF0zmyfy3G3zstpjcVi7uvOlWWqBnxcAx
cP75cGOEbYIWUGLDblvQYStU22d1qonyGyjnnw9htGAoxnGQbUceFkXT4gMQR+Da
NA7DdXX9iyttsb3LA3qJlAbf80dgczLEyP+cvH3sqZc+jTG/P9bTfPzasCF/KN0W
50Iy+M4MFH8tSLMs8CHru3dM2iBuwITK1Ujgkb/5Hhwn+hDyqyS13MgY4KbXug3x
wlkqXdsw3KWhrLtWX4WkcNiozsY1KRKDriD/uahPyJUAiiooVW/S6wopalhQ42Dx
2diDshxFno5hgrwKn230hxrWwDS+6YrtHSlVNkj3em2hfI0qKQx4qbnrkIOvwFZg
ct5P5ZGrTcxA63Y7KnCKjxalUs/bpPOS7rqc+EKNi2d1W50uYy+oc5zl/1mJ58FL
iaOua+yA4FfMe3Tqip/IqzPrlRPJDCgLJ42qzsk/eBdajocxHVh6vw3pdV0i/e5A
q2ORtmWYtyrJ5xdhiC9P6E/A4De/qSTNwbLPD2qMKYMU47ESGcbb82FUwumQA5oX
sXxhRHfUb37yagYnKIiDZQlfHigXJBBfc6Xe6Hx6NCWIy6+lqYmwd81sHU3qXV+S
exTq13tj/D2Auk4GO1ahb9gSIU5t4+wppwUZUHlY+AsJMMd9YXN5fyjjnAj308t9
LocInIR58vR8seKp6p5EdlbEN9D0PumS8Us5s3YJDZyi7hOGOTY2E0KFeb+V1x0Z
ISxVdUy10k0U/gEJWqAky8LaohVlM+8NDMxkijIoe/nTcCBiWpTWekJJ3m4GgxMX
nDSS/UFOc73KkgR0OEqGJM+8Cl1B3yfwOv8z+UcmQGahMBYke+NBUG3ahEhOBlq2
juUT7X4qKxQ2/E1NkxwNIFw+zlRpvlZI2yUe6eQSn5+OhfwHBl8kex/B1lk4IKeG
r+v3zmzVAxZZRy1Pcw5xvgJRk9W0Hn5QxZCrgVned47ihJFsuv0IRKhYldm/raZM
OutSUelsm1ay8Z8WjaW/8R71xZBtvFzpQZwMwakpE6wd0r9hUUy0OjYgEJHsLSXp
zW3xoRY9AYmi06xBeH6rpW+KVevbgBmzzSiYv3km4aFkzy5NXy6zV2W06PjWexO/
FXJji5piZyUNqRwbME9bEINhIoXwVoZy7hTbQ9Zlylt2Osnrj9joiOKH4R6VJoOy
f4fywC0vAWx8hrD728QHXw5VL0WQuxG2UoYPinBekGVHCuCgXDf2wJiHXddogSYy
wgUmoWHvH454KLqPgpMIeGbQEXAJX8m0jU0cBoY3VsnXTfF0RMBFsJxgp8yyKgi4
DvbP5RobJAOiiNh+pRgWCQI7c1H59ApeSCguQO1se+AuW1oLCDTZitPVjlihprLM
4kw9r1qKN39+/imbvQ6aZXnKb7+LW5SavoosLhbYRb9WuXU7LAXQX/qTyYPLeb4z
HiZnrXWRd0a8LMYgEKr82KK+Ai+CL8ZX3PR6FaYxsimkA7SHppaAmT6Sv6iovBi+
8d8Pk/jif+41SNo8PUqyXtgJ1YXBFOmCerMx8ViAxVdEz1MxDTisXR1taMHPNqLa
v1zlxNtLqHyf7fB0Nt2Dtz1ByZZiNGskqLygnMbcYso3URi0GIWMCk9Y5Ehto6Tp
oTzupPOJ2jI2+vj7CCot/p2NrrSYuHh3Gc2mz6ylAiG2DoWNo35c9F5xLz9zlnOb
sOQfGUwgXWWZkTLZfNy+GUL4mWWKtpSyi3T3hjtAtyt52a9wtHCEEtIWfLF091zz
/osZSRr84XrbduqgK6njDtjFyiQ7C7xp8N22GWYo/vOkl7VS053DhdOn5fL6MVhU
QSXLRacwr0y2einm/n8pniKIlaJDrHAZx4n5gnDM/7v6/BRm3HxnoTMWpJmZ7fTS
UqLXsQU+/um2Hhv3/2GPIp5+OSkj/kdbRXZL/sIpHu6EU69Gp1AAkmcFd/YDj3kb
GDj9pGAfi+p4DsawsFnyiuKhKEz/ciimicMXb4NovDSNY57Gj2hZyz8WHM/F0i9a
3eYaKWhR4wZ6lhR815XQziGnboU9CmvsPKUn/MBE6uj88zWGZawOhcVAbHjno0HJ
bwbm+LcrQs19Si2pyZkTw3VOkPLSGbbhF1WkBmkrU9salqDNXlwzZh5FnRKR7Wul
dtmALRY7+anm4HZVkrlVTyuLwrX1tb27lea6wMtZtNMsQbmwvvIh1oA60hUaFM3Y
mpjWyL0DEPt8EDc84S76EFo3wMF3AYstXfTcmJajmoekxD+JgSxbF6cxVypuZu+S
G2dVmxMbjfbwC0I9U20T2OyCP5Bh/mwByCpdHGqy7et5APbcv5FeqwdFy8L68a3e
ywgP+KokdQYH2VzGc4uhkA8FH3I0PmcWRH3irpit/Bbptr9RtHf+8BQh9Bba4KfM
mZ1+O9p0CY5iM2TDoMIUAF0OyBuZxquuiNfhG0gYORimIRpHmSA1gyqD8xrIJqkp
pwkfD+2vq27/6gydZ3pa3g6JS/ZJWNLRG0v4Xv0M0gFn00tbwmmamWJJjMeNzgip
k6fOdUEADG6TSu82+/MtkhuxFTtg7NyqmzB9unSp2jbb8ni31zeARWUoyYJirrAb
Fn1eoFO8rJthKupoMbRPt69TtPBoWuA9q6XiPN7CkhzbycYui9sLg6lIq1scUwKu
4XNQyfL7RBzIdyojAs0Vn1kC5t/04q5pXje+gEvLBw1DjeekCGbqxrARHWKtGaJk
MJrhS8foO9rN/iDEm1pAhzB5uef6Wi+h4ZeiRjer179KES8eBKlkb4kXPtPCj+QF
EMIGaUfv2YNJAlayuo4oPfCZa9cBGbmwQqhKiaEr06rZ+7XbG0Ii0YUNLCmnt4JQ
9y/0FtKMEl3wEjt6RCl1uoyr8Rw5Z/mIXKTetAZERiQnYUHl6u+bLI03f468BBJT
88Q1jDpKPu+mjqsubYwJcNVE2MsiOsCv4l/oO5g43r2DwxyDXAUVXvIdg3KW1SbU
uHNdEGd4ce5cgP740UvVh+QEtTQEfMjMEi+NSu5bKx92O8LNOapfe2LvMqdi5FkI
LsHgbLOeezELP8q5csYNMxuTKb/QhG6/lVLotw9W7cSkXNXQy0SU1tEo76jg8oWI
Le2cNQOlvn28BmcwwXhgRPgCTSpyiGeEav1Yf8xb96xvIY0dtgPUkRBnN2jaoxbS
QhA0w3WLJGKJ229dqtKl31n8/V4HSumHIwXsnRR9IKNAjFy6maWyqd7kdSnzixow
3i8LchwdeH135d8X9fgSBfYted7mRnnAW1T6//Osfdv0qRQMFSO7uhHDxbDELxh6
t89SNU0dpkSNzSqHRsigWVhWd47KZYeEmnemMp1gY7SknaoLoCo6Uoh/jDuFpEOk
yedOls3NrGSnoRyDr7Z4Nsm27q74OOUjD1rsZhaQ/BQL4YI2o0W6Ag5BmzV/HM/2
xmEoihGkXz8zu6zRdHiVlwkjpDjWX99Y/3+j6iF2BNo+6dLaQlgvmFaU4ZDWbcES
NwRpm1ut391BtLB1nTVonUiIQ0jNMZLwa4UVAXOxsGABnrQfDDU6kQVqdeXJfTU/
2HuTJ75khSAps1ibaKxrd9nbHnT6ySU5KA2faOnpssDQ5TIbcY2co9GRuf8i7lx5
STpW9crYMtPLJfpd7QLV3RgHIHInMJbEydUhkw6BJd9v/an94WirNFQ8JgUXiaZX
zrEQjxUtKmC3/U3nWLew/DaXeXXyq3apeGnAa6X+/sznQymZITrnSATOqqxyKRbE
2OhAoUhD1tuo+Kd2sdL2iHrdwTdCe8C6qe6FSUPkZLSSQHjSuaIORAs212Z2VFjj
t82lISOvLKqy1SNybtTI3DOFyt9t27Fdbmg8+b0hECxAyvkFSdigKI7Yu9yx+Keu
/TMOQ4DrI3eIIXeO0YyjCNSKNvPDJxtg2/Tv1lsYGe5YeNL4fdshYPjCS+iAjVkR
8XdthQoUiM+0/0N041zgJRMz6QJe8flsAIUKVcq5CT80sUos/9E59LnUsgIxgxvT
/6F9qGGBP/j3SCCWXs0+I6mCF9FStrTu/0MNFn33Sd0w6XCF5WqQUwLm49PRzWpi
Ke7w4Mi4eg1OKzS/cjG9MrLnkrVDnuYHeIdbXXyXj+AUtmJfvMlWwJ88P5r7JK0L
v0hRwZEtlPUUtBf2eTc0TtLpQpykXPDGcysRkUzJcOa9eQyMiMvU4bElzgVSOZv+
NRparpNeS9K8yBubFZPZfhKAbp2B5FYEyqs7HUDmNu/QQ4/ShrLuRizBwBblz9Zx
ev+bybmuy19cN/I5QrzB/IJLPC3LEvnmAFCrsbi/sPfxu6oGUFfo/Dermtp0brMY
wIliYyaZ5OPYr4YyXHcmIyZd14v9VCh8IKHoRyO5BvE8ODAMOsIUO7xwi6Clhlz0
us3JkauMqucL1buQMMFcZS4WLEth9oqVnd8L6AURvujKKFC/rc84iqvu1NfwkhF0
lq403xTQ1zpHLZLqqs3tQ0baiVaEzZ9RC0Nj6URhfjJrwodue75aJxx3DReipoff
1DJemeqapg4l1KBoqWdqVa15b8KsEHeBZokrViBtt7QkYyPgQ0J/Ax9AkWcPWwzY
kyuiV19h2W9ik+4ElLLBaRCAsQ5ngTMQnKHugdVjpREVi1n4TKmPwx6MYlSIQ27Z
ZV60aWtQDYMIfuVz4l9q/YcZmpBZhUsq5L3YcGtURqnP4yeFt1l9UXPKVT2fXDX7
U6rJpRULGy4lQye15jjqc4BKAQDoxfxX0QQGumjBZIzhOR7S8aqg1veZ8Fz2gcZq
KHEZZhkw+9iONKfdC3uJbLQlKG+ONlnFHzXvOCrz7QMkyTiR6w4twhp68nbEHLjM
WueHOtYa8toPWYjJfClhWr/IBHiUD56/puCkfsJwhksDQFS9cEMjMXRJNY4Xc9Oq
ZazKhW3ow/XzuLd1Yb0siUKcZ+1DG9qfX+U434Rq6JL8wuGrGxxrPWIOMbvmZzHg
LkILrKKfzR3+u/wpduO36k+txR2ShjpxCckjRbJrRucJtm+4Ogl1vaOBsRsrm38+
6TgiPnff+4nBlEO7KRBZ4fIWvXKs0/SyyMfh3cj/r9XUhUS9l+szia/BLZXnGH3e
7fTNZohHIh1w407g/Zel7/pL1Zr+iSf4YYoMMxSqcOjD7Bzv5FnpHeioXvmu+gkL
KFPVuyqeqTJTO+MdrTtrSQ6s52qrVk3GiGEpnV68diKu9kfJdkgdh7UyntErC+pE
eJ1VqMlerLgik8ol01S36WePSXaL1x2qIjrYOEYQxh1cOZMP27jnjfMaxDPPgkEj
w9tRjmBnwv3U5G+ifBGOCbf0alnpnVX890PEQI+508+SC0OVvRn+WekILpkeOduU
mBTyp2hStsUj4n1zA5JO1B/ZMCdUpGZy+0GPeEGw03s5Jt14rAUTWvOz5aRi1lzy
5C04jr4rtPlg0Orq4c8sosizLH5FF/rtmhAoE78B51hSXxlK9XLjQ/54qDX75Nwa
8MdPxKuIacvzSHVxFyOp0BDiHQ6J71ZRRGGPbQZLtwEoqy1+fXGHKhG9f/rurfnK
qPO9VJzv3ry2/vh1KKzRb3jy473FXrEy2DyRVFbrbFWOdHRv6Yidh2QMnQjB2aX4
O7Y6m5v36OlGnh3AschvrcPvwcnTvQ+vaTcyJC4uBOikTmalFcaopULVRF748DPh
nIvtRWPPYcHRpRoKmR2zg1XnjG//3/NL0lS5tiAx+nDwSLrU12G9KkvFb0FXCmbd
RHN2vdXMGQLdX4mGyMsaAfYNn7ghbUCOoE/e4zBZe00Kcq17UVAoWgTgjOBdf3lZ
+Q4ooFEF72VoTPis+Z/hU+xx8wDSmnkzptU/284PCEqNg2xNcrWR8rNZwjlIOaHm
Nbq6lKnIp1KjavKmUmNMQk2J0JZagyLR/uA/0NIp3is/XSb0hlaeeGXq6f+cEaXE
YzT+7A021tG/dpkoAUsHBqShImJeSsoVsk+vsaf3J/0Lgkq+/8q46WgVUaUV0nY8
gTHatoJurCmNzXTZzaqti606q2elns0bv0e7Z+JywYVGH4L9JCX2aBmBqRXpbntR
8I/wHCR0mEnlWPMHWnDLgwuXp4Jzs6cppyjLj0k8Gqbkyv0BYEZhbqp2oy6LOlZe
ZDKgkYMk7zr0e+iTeiQcQmDw+AVUMOCjHuFFzZTo+W2KkGUx4dRzCbSHrA/bRspe
hTjGlgV5BlDpS/gG1q6QyOMLNcO+Eg3I4jCm0nwuy0B480Q8i8FQ0q8i+FcJBG7M
RZIROFHUs2LEiVMlo/RQXw==
`pragma protect end_protected
