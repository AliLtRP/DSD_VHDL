// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fe9s0aE68j52ivDJz5BbL+vva0FeD1MiOXrwjrrNMXgC3x03pfLOr4F5gqHWdv5g
+ILoS3GjqrJ/20X3uXHBArLyvznjwEXYM2iFVp/sCnbSsDoj9nt6fVltLVd9C7TT
N4jLSK5uywmk+pYonMeby3KNhShpsPUaPD1ZXbw7edI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10432)
PEUWkhGN2YDBC2qfEn9B90BkYFPTsSU4F27ARsWKQaQvLkmIWrib8Cr7jEtyIFfQ
cJcaObCoEro0UDzRTZMeDELr+Cc4fF6TqN5IbO9DPr85jTl+QhquCtaGctLblOVp
na4Fp5lb/PVFStp8jHG8qNOf48yHaTxiUsbTBGNYpRPwiYtLwI1iFeVronOYa6DX
uxJ0eWf6QgLI4YtiCYUQ1kj8DQw6PCIpUWhGNA2e1dSgFxMZn0cOCq+gwHqNVsvk
xsH+9R139yEiIfPBSJ/Y/IYqkWkXK6/AbkQBnYsOePUltrG/Lr8oWJ1JyHIrdEP3
Mb4R+DgV99CoR4fFCthL77dWZArZacSIY+xXy1Qg+0zJBV0O+Lv5LZjNFWMIDufJ
u23P//EH0alhq99ioMO2+utcda6lBG+H3qX3hoWu0DmagtGsRFRCioEsMVj4/Iwr
KsU6VpDpvZtnDGGNxE7Lzt3Fh6EHqk3U7bWglVDPKIt2sn2290Nqj/uK7Cl8p63q
S3V4n5GjA8UeW9x0KF/kcGK4Co9Z/j6nTCH5L+DFc7X5LY1KDjpnYMVtMdiUySzT
SHchTQmL0eAkvcI0F+fyKJTotQXlScU3m4fX2gceaf6gbxXGfeogvJ5eB17nf8TS
kkltRmc3E2LSS6XdFnrem+UPQuILX4/kW0rhni0X2letF470lfZlh1hGn4cUnDXU
vUDQqfNWdz8cfvBQa18vvDzXawmYvOeG+6N1jfoOHvlb4EFJ8CHYYnw4kul6D1gz
LkyJNd6VHp5FyGSq6sKRnU1zoFVk8yOZCscNnt6kw8Ti8vlrWdMO2VIz22jALSyH
2eyvC1vaifhPJ303v1ZSOVBvmSgZFqHWZE8v99JZWodBtvVNK1PDI5Ik0MdKqJ9Y
q2iPd4O4/9wStLi/1GCHxIWU6WH8G7KthKh50+sNXeQZKSOcy2tkPUwk/eZzyqTX
w/L2zFXqzy+5J7J714mTCImLBpSgRjYqiG1smvyTjlLxIpiBZQtpI3IXxb0eLp8h
EdE2XAXFWLOb2RfU2PT6NhQ3U5AA9jXg2SbRzWUmfxkzisbM25GeRn23mHO5c6Na
9XjUNw7qhClyzOsMa5ZA3LMvhmEdDjfxW35Czffa2MaT3RAIILHMhzq2nf7QkmFP
OfXWGPSJiTHOuY/WR3h88I49G0SFy4pfwuI7+qYgVRRUw+lUUZsTpAuWKL0KEjAY
xY3kIAIUevsRfYdgEoLWM/MN6cVygHnDf5NJ0wNnOshCPlW02VU8/zXP8Z4LdCi5
h2IXFYq2pRkWmLepQJQNXezZAQZAVY8NDc1xdC+5U3E3en7WxSGBMitKk39+Eyvu
f1esfY+ORt2m5p82lUdMhQvbhcT7ZtXR58vlrYJIvEcU20lRkCxTQjteYgYZAe9R
ymBUfOG9gYJkLwVemZc01pBa0ND4Y+fjIsvZpvlE8dDS/BHiGCSM8Qsq4U/QgdzY
DIlX4wH2v7d1Mhg1XL0FK+nmO5TwPJhgoBTzA9Pt5lGFBgetC6KA97qi10dBmIxi
e6VBR1YUdmi0Y0LWff96ClByywiXDO6lLB1tApXEsdRr8+lf5yGnMgVMIiA+qtZg
EoIgA7GrHcX9ErpA9AVZ0wLfctaUFHIOt2CBKbaMBjRSZCaea8QnaZq5Lrqkb0Zy
JxZN6u6UszN6cHEjl63CsYMl4FQBE1lejz6A6C1wAGIQPODObsKJ1iNpg2wUkbFG
Vh/UII07s3+s/kJUwtvAz6sD2hXpwdYQ9b1ybg5hINbVMaPZ1DBySUqh6a4CwLLq
QQK53gyZ3N4tYvsN0KlIPmKsRNUhL/ZvMUa2jQuuxBIOeqS48S6XHm6x9sbJC9yS
zLDjfTF6UU3NWP8d7rui9kw2soZQR5Njov6KDt0CYbSY5NyDWIQWbeOq71lr117A
c5Ko1Tf8iIUL/gNA7i7nUs6NgjijCViXhLPKO9WRXAZC9pAmNYXYpRBsrOA101F3
EnjYfg3/c9ONCInsHMO/XNHX6Yl/8ZoOPHsTpqoomNr5Fg685C7Dqa8Ro0LvaXB/
IUvJT9MGRffsNu8DlzQlqhQNypqpiYZgfZnej9eU3ywR07ZevkM/BGrSYv+/NjIz
L6qxIN+P+CNTjy8leEVf5sveUYU1C0j7Z4bERY9JTESOwC6dsLPRsJjqaJOvnTcY
+7/6lvQWWhqUab8DDleoOMsVI76tVqc3j343XCscO+5M8F8nkgcj2VsuGrjpw2Dp
WeSsEn/I9cbCyYLB+0GY97ofmofv1g6MbhgA49UpUv7+SD5LCBhnucUCx3xD7KdC
poJU5zTsB71yjuuxFI5ECVut7ZUJ2UTy6gOdzoztuAJ/ynoYv7i1ai9bu5p2s50C
G4LrzeppcqCESD/sMxzks1QyEImRQbGJwepc2V7nbjkBsiCNPruZUEBaCVyPdzgJ
KyEukFqUI3dubWvJhWnSbD0aiVd7jWGDlVfPaBGVMMUXxWQfqinrMVMnTEa9M2AI
gu24nlIfPGqtt4Cvgmqf6N/XXoN1ydTiU6SplCjD/rZIL+z7BOz8WZpNhaA451WM
mNQ3zW/TCtUbJyU96YWFvpKIuAzxOCnFd9VGZxTKICxvZqCREOQjtv8H/04g4WsN
XNe86ahZ2LesPpW8SiSaAIkorV7+o/KvI/TL19hs+IQyL42Yc9axOZaPl1GjI/A6
D0TibRDCz8wbedaVxZmnmjKg1fWkkppQln45LfG67T4XMvmLSTUoZhZnG3Fu5LIf
WSYPYX7nBHqSrToK6/gR7swIWzxoGQBcx0x9AodOSf63gi20pYZtXMYfVrtLhqRS
qKxPZFFD2ZG6CfJ3qkHLINQgJ63A9MLdj2yrfkLQsfp4tlPwsHXSh1eO0+V1DwhM
AnGGgwbmVSb6TIGG+7gGPJOICJAbweomFoZ3qKMQOrm69xcUaVmsSU/ygllAagRT
UlJYEyIDu1Et2ZgGAy9ho0UNgW/tcGk3nlgoNJuKxeSWAtHocN5Zaxp55z23O3VD
mn8VcMs7CJCl7JUH75E0iQHm3cdMTaHgVq3nwzmcLvnvFMZaT1H5tpNyj/BJQE2l
UDuWuOphYJMz7yqWbu3TWMrrd27W1h5/aZg5dBzxHrA0B19gHev1CKlu8wWj3tDz
3le0dHY8m/j3myYCVEU4tQr+H0mBGELXWxlsR/mQEs0ePGn3nWqdQgwlUYvVYpeH
fR1xa9nz879Jc2TPH5jHrpW5rNrXshf9uY0udSACSnmfO9DBFUg8aK/03xw1WZuM
KjC6NQH+IU6VSEKkjpSMkF7jBTyKkEfjGbh7L1XTJGIRkr5y+dXiVo00LihFZSRV
aOnCiSDVuUJa4nylXWPUoZXAcKBxHEoeLzIQTjWdtidBWve6zEqNglqRAZZc/F5d
ax6BgZDnBD6JFmhY6FNiyjmNOnXepSMnVKlIdYc/PEu1XPJ8zEQvBB20Z2YiGJTX
rUdMYsmMgQXzCtJqIjRsIDllxm3zX8k1MpAqVA35OXY7i/LlBLiRpvIrvHUB3xwf
DnaQGtGolx8Fv1Sq8bYjV+71kAFYC7uZAboIQKf6hJ5bsaT7xetK9QhzpxaMv0aJ
eug+Qo2xl4L0BVECxJYgKj0Isc3N4cFUq4Bgm1/gX4OfpjVyOmrt3a3TlNCJiNWv
KXB6HhSlEJSZbribAkWUPKWINDVGB9bjfp87QDFnIXkq47eKnRSuv9h4q4kKNPin
6KJ4eUk2WyXqyCi7Kf1sXdiJq+qeewcXFpKq+huUVVXPr7TJqCcwh1CmRb9e64y+
5fwZMQcRHymjMb7pO9CmbKKVJ1PA3G5bmaVAM8PI9QGCbIPCRcuoptI3Lj4js2Kz
Rqd4VdJ41mcfM6IbTX944FU9oxPEiZlnWxOSUB+ConQDG9IHna8V+AQDCsnaG8OC
SJ9eBU+cpeCXaim4IQ1/sh7eA2jo0ekUL1JoRe3bvekMeQaHyMEt3dFG66mBDaKP
ic4zI8VXchOhsafptfxV6c30YB97udSkSMUN1SScMpNuAhSVpfWtAjwyV0aWT9sa
5o1/YzaXg4VvBFge89oo52kkBBUeM1GAuKRE7A7af24t7SuA1mWzd7E/s+vsomol
7rhuikHf43UHOwL6NxqJwwXm/zzqHCL/oSkr7GHTB/zCqCIHoWpTNPGbkyu322ju
dBqDTRfhQRDJVP1WzhH+lu5ZnfzJTI6CllJwQFRohkZDlX7/ISRAwfZy8C8S08eS
0bnOHjwyJuBCLwmxsL7+FDWTC+SU/dTwkPnt7E2opxRvvkylgQlWkWjQKSJ+kv4h
EJor2p56dN3aKEtKMbEzKYVlUfdQkfk8r019Nk4yR/+pLlFPoo2CnxOZZea8WEMH
SOYfvuZWMavy6qE7h3sr1zle1rw8szq3zTD4HzIcQRpxaOKq6p3NDIGvD6tRrk6p
OAC5k7aSKZqaTjHs25G/gtJwpEdiHiHapjWya0cZu2odQGFTVVsb4KSiUJ5UjF+Z
3ZpQxEIvHsLx7TYPKN3RvaZfM0N8i3lKlbgMD6DKS+iTHz39gv4hfYrAbs7YgCil
1Yvc8DmjmE5nuKs5ggp2c0p7SlqbOH9qJJZJD/u21WMSO4Y3AMRuUqcDRo8MRPZZ
bn9KOKZPnfLpBBykNOWnssLAIoU6xYCwkxPFXINGGxTXpUlL0+Hx0hcv7sXgxYQQ
oKCql8a6/3hG8q5AfMGFilU8XVkYxRXdKGxCIBkyEPfI4g3FzQVlVpxVhMgXIsVY
vthxBGZsxMMT1YHvBkbeTfGXqxs5nkjlCpPS5Oeir0qZrKUfTgVI8qU382XQ1lmQ
Vz5vuVgpzPbRJ57+L6qgkc4mThs/Sb0zDfWJeP+Ge6KsgPX4NAVsTA/sAdzCC5k/
7Kbm+K8Gosuz2VmxtvPE5wIFT2ow6hxMzhz1/MMMlsnPA2H1AzMi8n9dK1XKvhtP
3+ORaQ0GBulgPvCY4AMcRUqEnN9lwFDpOLgLw7D8N7l0Zx59n11mD+haIubLIBAS
6YjpRRNuNi7Wq6EiUMjuzWaFq+Q23HR20trkRI7KrCvPLbBHa1cPqAD9QQKEIfZJ
GJ7cwSyfy3hk0JGVoD5jYPDSM+qMwvJfFy22bHBkXrM26URMiAYbTCwroDzlt7pj
O/gxgJSpzN7eEZxYWuuIZllUM1CnZQ0DxiVECfR7YtS/P+cLhSVhxHMdoMKnTdkU
7fVOxW4b33FducZVYcVPqIwxpUxgRlEDCk2mCGCXPIit1B2APZ3EJqj3rIGw0ze6
2ANv9gsuULsIAfOFuH9ESw6mwzT388CSxmjodkYniFtBaKDyHYOpKowX+AfqmzWX
wg8amgclo/L8PSCJd0/4oh6Oxv3KE5bl24UQgUBnbNVNMeSRjFIjSK168gMwswQP
miWUpwPzGwtGh4WWZcHzM/MzJSmima+IJayziegN8f4Vi7MgtFSdmBc9qpw3Vqs9
7a9DyYGrZDLOwCIefgpyXxXjlKgvel3mBhfjDz2qsi4HHYbl6y6SJaPyXGX6NmKi
XUcYt8E52G68rrxmD6+Xpf9m2Ec1XIT0YYHhzargT8GnpRb5qDe1QLyYd8TwH9sS
DVyEmxIz7GTjianIzPjfQS4+I44zpdUbx30EC9ySnscPdhtuNpD+jTX1oiO2XF9K
37yWIllDzgqzkJlwEmBszFXGGkt7UHkB4rRIjiw4U0myTwpBrop4IVUTM8Aw7JQc
22j4L8Ox+qzlEZnuuRUWaRaYDlu+J77KraOd52Z0V1kUls/yymSfdGbgIpddzy1N
c65QTdtgz4Q1ESyuQl2+rwwvihzq6RvUOnS3rjsh+FvfP5OTixtCANlVxGg18BX0
yscOKwhwi5jQT8BwcceEhDgbe4thNitW++A34CHFsXs9om0cQFNEnXqm1zY3rNhA
1mznBH04UQCCgwOGvqbDgkBzHLJAW3Rc2yNN2WXIUleKQyeh6Xeu2af2BrfaTkTL
YbDoDcNo2U7mdO7Abfi8OpThiruXTR36N+zSYPA5UPlfdras24hI25nd7LGOKfMi
qPGCKp0veK0o+lBQJIOtoX6EXRbu+j6V73GJUiDgqxY9DA+SwpYDr1bKLByV9NKP
+1ghJKGEqt6tU7Au1dLWCcDw5y/XyVpQMEBtGGAdOqZF7P2KwDtUca/VZl37Gz9t
t9P4zoKon3cZVUWOBO9nPEgZkXGfNeUn8BCF49NmHofu8PXLvyhTN7lP4q1yTMZT
5qFULyodeJH/+bdLQ6B4W9gC4Jiz0VYQvWzAsonvdTd/DsJYaHWYbpcJPebtsFDY
8fGU9L7ZJfRD4wT1vyujD4cuKspGNSq49Z05vIychVxRRV/xSthNMF04OsSSjKeN
MHYumjQvxHZ6Bhxo/rFJZL141fZTuepmGJKnmEUteTHP5vH0g2P0jCJFOeA/xhsH
2UPWU38Ymk5NNa1F+dRMcJtYY8xzUBPNPK2UIuYQHFUnkAdOL3Dm9+4UvcUs6113
54itawgpsOYYkH9P4SXs1Xw9vbqnEWnIFHmlKgVoRi3yEEpNkP9mzRJYbB6iNBGL
kOnjEpceMulvNdbFvX9sg0cj1C4QDo9sZx8zlMV1MKoKH4kTKT1Gnqf7dr0FyX5/
7I4rA7fTJVQOHj5s9G1TrEyo8bFnRHwgDel4nrZlNJbirvzyM/ZYAdwafpXDHAoT
CjwJNbJ4FEf3icetMB4bH3Z0O4qiQ0YXHWRPXQWyPpGlJ78F20epgy/vO6vOYWaH
Q4e6EjayZxLGJ1xJMPsxfjmeWFJ35KAWBnpp5+tkhmT2zAMCM+HH60mPDF9CVkoT
gmIwwIey3igNFpHJqLvcjiyeuJRcQbYBGSAb4mADVyeTjUk2dwL1M/dbeywizYoY
WRr3/Mg++pBb5sDo+dSgkhgXDu7pEzmTRP2jKiEJBz7RGQvd3KDL4NU5e25/MwWu
oG/upuPJe0yToc3xmeARfdor0rI6VThhN7/FtDB1lz/VTbXyIoBfuwq4yVS7MjZE
AW3vDQWwcB9Jx3rAh9/64mS2ajUgWHc8biiCQwtaSgyxfauVBvGkTo1atsQp1u1T
Wwy6Rj+BTplUTEn5o7uHZ+/CWel7wH4qNyLq0CSFRDa5JWEP/4kaktuZWPM0l4a8
KAKzMn++Xg3NeJQSj4Vwqja5aw06bxNIpBSxkpW6joncbEC0QbR0uboqdxV+xPFD
hcN1pWLIIWTQpUt8EYaWCJIRDDo2BAI65kXDdUnQQ+wP18cdJJrQD1aziXk6o+u5
XymX3uJMMnj+x1vZXD0kf55DfXJxfdp7tS06GIvpYX1foN0mJQjLjaLGaGaMrGLY
fwKySnrVlP4wbNbX2ZtN3a+8Sl3uJlrkUz4bpa1zVbb9RzOKTWXfXzGFGOLZRbbl
swRlideYzNOYpYJDGXd/7uN3zROJxHXrG8qB8rAakvQLujH2F13SsvCPqGvZR0/S
QNvFWmgM1pNIkjpLj1PxZ7uhRCsa43UFtMs+dQNsg1zpjJkR7fHOnvlVkrT4wx6v
V9VXy6i1KF8nezU6ereylhYKhS2dPyT+mLgBIMqvHhdIihSNWC6+2ppXVwbMmqIz
8JMgcs+bMp5RDCDUrlM5shG5XREwVHxibi65l8ImN82gANiyjQzpYXnaENykRVg7
tLXTsy1qCzaJQrg4YfZQReeOJYifXiYMENGDVdmQDt2dqori+XPll7VSA5O1JeGj
mgcpTqF/2hFMyZaS7MvKDnZQDrWO1IX20CwysxwjvZdOKDkwTkACMi3B87rcYIEF
P3bc4k+MO05pRmMUrFZrSqR9aPGPT9GHu7g1u5ld8HmkA7nk1WuABBCW2LRqu1pS
m2YqWbQofVAXucYC4kN1ojFz4FVvvFadKrxQp8tW7NxedSFxFeZD8AwZ+pDsieDR
jMl3P/e1OWi1kUXcmu1vuaYzychyuxHYIvbDK7hgJXkD/bMcVgbLsWj3aoRae/d0
vcZa0FUBVdvA+z3jJOL/iGlEnOBs9XsnWxSNr2Y6OWkfc8ePE8lpQfA/wpbIbSjv
bczjJmzdC0+nlyuJ8pqPwlUjm6K9zRg6CenCVi+KKIgJx2r5/2FMwnUHDh/IXUIx
6Ek6NWrC5EhW816SeKkPH/T3T6BHFk0G2OvJN6we1uyQoae+NztTQGuMzfy5+YJc
8Kh+FYJVgdVu2jv2S+EeTbO0njqsqnC8BxgT3q2MidQytZLXnaaYqJ6l5t/lDto7
fiuDaewAiTNj7NpvwAXihvX7uLXTJBZdYWwUUzpXiYE5KSmZNCv7afSy0esdC2Gu
a4W69fxF6Td0ovtsTVFuaCJ69mru2g5Z8Ym9e+bBbYiByorvSZLxpxPwxLdsG2O5
7gBJD2pDrNpFTBOWZTK2HJMfGnJqKFMBPt3QM7AGxmKWhpPgz/KCTBKQMdBOryER
7qp2kqFM1/qo3QcalJ/tPfwfpQNdAXr2cuPIpaiJTeOjHL5vr++TUjKpIdlY+/LA
ZyghwYMVUjFfssufSwIeo9tmnxtSlv/9tpUnPkcFjCxfOU6Pqyg8GnXpR4Twk9G7
3WA+ABzLlZrVnmSltfsc1SwqqlD8l3pWd41UL7AkKGLFuCPmm6F/dZ63EtZexdcd
4zCSnx11E2PFa5hx5QDaCq6b75QPp9H+7m8+o734bJau7HvHphfoQG+V3rEeQgXe
JPbh13vhwsMkdKxMn96TqnyUDJ/F+U0z5R89+X4KiG+ryUCmZsWKImvsBSxzWnai
tfQJuPlzKsrIvZshjv0MbsX2PErc8AOJ1yOYqNS+6Q+OzrbthNzsb+0yzdPLxjpw
YJOQrc56FuZs3pO7O4aSi+fcpBhqQRdRfZ/HthJZjFo548uUIAhMZ0LeU/Ly3Lp6
sArJL+cdeKfFUIHaVLEwMO3QcV1NupVeOI7er2/GpQAMu2RNAEs26wOTuZDjbLsC
LbI1WT6JM1Spx06FX0qgoyuTJaUOcB5+D9BOeNE2btgcoporQqqz/sbPktvlOT47
hkU3csPb7j5AdBoidR/xGR4865b5vyqKpHfxHK1QaalkgnPPQtnCpit8Z032Z8TU
V2HyrlCL+et1ughuF0ICPkk51+i9HCePbS+4vOjROonJYGR6sI/xVqyzDxBY8Zon
naU65+3dXJQncGlwTM5nWEe1Qx7uMilb/+nG3nsM22xzqvuen6xgRovT1SK4Zewv
pgwxC3VItvFyJ1Hq/9AFb5JvuKEPRaeUar7LIWwvJkdMS/zffU4su0VLwHSgsmN2
A3Ey999Nqo6nvKRPbxPKhM3yyCv/6ObjuEJNkCEffYtShXdbCcvgWlajQt4Xfzrp
3q5aINekWsYCY5WoZIA3+bHNnry8HJ45yP2u71ChIdPgDSxliKs65F8YFlrGibIq
1SfCdg+tpq6/GMTBVzZF4s1II8DDOIxOfR3iGgsl73b4BUsjTh7pUy1yH9aJdWpl
CQl56gXiQINb1oZp1O9LJlVTxgQPwEpKCppoSNu+sBQx+wdtqZb7ix1rXGls2KCy
m155ZdWRwgmWSW92Ld/7llZ1WsI76hSgVIVgmtPwaxNHnl4YW/O3pWdOAY2V6xNr
+CoxQjAR7rSR7vK4l6ls2Y65bHYYJXrRETlQZFwNbvs1zTYWoSQBsLi89hN+EXtj
MRM1PaELIgwIS9sEhceW4HE3+t8Ouo+BNYQYkR6ceuGrHHwazSCRFE0lVzSn0Ui1
U02g2DJs/5mjI6XyBzzo/V3dRIAjQUgcBYjMvUtLgnuwDN/IUxjC1Lkgijv/5bak
8OmPDsNaVlnbGly/agoQ20gYwS9UUPC6nxgrTboNVeaz4umtWPUOThTFv8ZsJY7i
YlJgnii/DGGvvLV6KU8zn/G1v/qx7FGg4OZBMiiTObIYSP7weW02lvmuTeLlIiZd
MyKr61GUBJ2UbgYoC9TakbEjKHMBcUNTcd7YHtAIZ1aBZf59F+TLzG/IX2/2slSf
iFecB9O4UOiL4fwijv4t/saEXGNFXtA9TXNywjhSD1Ejot4CPeFfi0iOuw0vaoCN
WjOJuevdjF9GrPfZhiRnyTzPz9ToA+g8h9nnUSvQzrvuuVgcpqYHJdPrC753QEMw
ZhbqgVfoZIWZ3TVnt8FQL0TBhyXob+Lrb0bq8wQe44e5iZ1JiKnQTOirhJmaLpT4
Sprj6yOqUOOOPx6QWMDeyA9PVMhieCfOKHQtmR8zf/PTU3rMfzgVggpOoHMDkeKY
hjDfBcGgzMOas4bOzE6LxgMqHCLrlraQrRN3TCOKrAkjpRlAr7SaxlwqQLcrcb7o
GKn48wf5gVS4UJ9DWePLKIbo9+crXnkUyn7xnAZe7K9CbfHkkS02UWEWuSpZOmDU
2+2hMWAd3w6S2ntsZXrX2A/nUZnNsL4kXBe6nfW2PE86bonlLg5o1+YBfrTjaqQD
D17dDjlvN3ZbYysPRvRtP8wCBOyBlXg/WD0cyMno3LkWlRXpmdXndof4doUMxGup
/MbTEcftRlXOPAdZleiAzdSqcHi24tdI+2dnPaGB703uK9HGIWMjx71HekNSfH28
1g91Yx84s4180qUXusRlB61mPobNSoNWox+onhHFpQYNG8KBnycIn54wdbIyHqWU
+vfZLKYDrPPRx9pQhRLunnUZPOiItLzf7JhJahCPjvbq+MPVRFnXzj6n2Uri9KKS
6ZmHk1NBMkMoykRqSc1ImQKa6EVIMLXocKz/yZhpXdBsWg9+xbQF/q7qJ9ghyPG0
7XASSaKussOqsPHKUWKln6RsagHnlJqVfkFOBlFBx5un9PAVW8BX2Gpgy0pFnxz+
CTAIqTraZRq6MvL7fLN/Cru74flzV3rQHGsz7fcBkKxeSUMY+NuP0XqSegSPKVlx
j7cDVfUgMtIbSM7wXlVog7GdDem77tImXQ5X8/bFcoeTWPTPEJHg8FlVoUnaazVl
ZLd1URBAmBoAVhytQ2KWKGKfon9JLZnhkn24cdU53ibaiA7i86VqSUYGvdqnlu6l
Y/5wg3Q73ee3W8gwHzz4RHn0MrhyIC4Nn7WR5aH7hfc0HoEMOWBuofPyyiG6NkDe
PjKkJZ9UIl59GsMxavfrsFVdoL4s2cTYZ9SLk08EHLTFWjlw7OHVRbipZmh3ZyL3
7iFHpPWr5SiJFqWIwgObxUzGscPEgenMQRmUZGBbVOMLGTH2a2qnesEUSX2sU0p4
Wkix54t1iM0dLMn9x25tN/NdXkfhKl1nhO0gbHeVQdgSWfeFI0kpZfdhFg+PHZOQ
433vXRXQEG7I9iOn+6tLNcmX6ibppiiU3bNBiGnMnBpLljXRpfk/Dg4xvksKf30T
/CRFd5FCOUB9BaQk7aZnZMOpmUMstqBalbx/I11aAJzU/qGinbxLlfjHwdwple9R
2n/zO7tlZU2lUAR23UHcYVAu+uAp0Rt+btG/JJZyq+3OJyjWA/DR07zOBU+yc28q
3gEkrETzJdD67viwrGa+V0V6grPxlnZDKDIuBMO70bxv5ZCQ6YVHm1L1jMZZ+AZ+
puBwPiPVyAkJ4Pe4ex3phoJYHzsIg6cbaIhjhDm65Q75XBiYgsgU2xFozM4ESEl9
yDoO87LP2SEarzv4IFi2CO4I3v6OIr9o+TE/QGVWsIFeaPTyzvJbkdAlaj/4ftE9
VA79S7C29Y2UWoYe9hvWkA2MEz7WyrP3PnkX6UVbpOzEH7PJo4WaEM4gsk9Ulh28
ZhJYIUS/9Ic3PieQVJtOZRNJ1OYv6CTT094qAuwATFcrTzgfAVQIV05zA63LDpqC
k/MyxLBaOQ6LaQJUwH2xPQN6dkb3FQF2tH7cEjz45s9nQ3JQA6WpSDCs5HeVE1WF
4+5xE97xGJ2Sqwp4DOAyK0q7wHakItrRsSEjGTviCTYe4FwJNlX5uJe9S/nAa6Fo
FaBBYLcIfC6vDgan3YwfO7dMxGnEwe/dDo7F8/1Zchm78aOwpk3ZmdmKCCfHDqKb
BGAAQ3A6z/TXnznBpq9V9tc9aV8zpgx/a4Rx6umPuoRMj8MMbuUWNXv9RQw37uol
L9EV8g8a6Xaa44sMpNYChJmTp1vSyBmKxxzo502n7NP+lOBu7UpFXF4h8IGRfgys
9XITyT47RHDdZ6jqgNWWADd3XMQNaqZVid7tcz84dUcFU6YinygwLmqWUHVA+uaK
44zsHvtLmHmyIN10zr47OdU3WrKwbXvwkgmZyNXo+31PYTlS/Ejp7FfIRqHrACvP
3cX/JD/98UcbgU51/S66xt7VyGL6WGhe+0MMY7Pbmbr9j+K+p9qpCN+7N5s/2vdB
f6WDgpRlAKaQBX+zrgizhjPdm0s8YO+SR21PqRrgoWl4KDKTuiea3Yn4NwP8IcBm
ceNj26k7EM3UF2oPZ+2K8yLAVlkSal5ys33ATPxxr73vkJzjuJgMxISnH0SJFpkj
UG16su6QnD/csHPylktqzDy/TjONt/cXaEiiPvMGHvCcJ2fb0MMVT9//OSa1A7r3
dUZgg0Iax5w+uvVON1Ua1AsMQvAFy+P99IQmBFiGRADfc8GlU24yPWYwWsMYZhZP
+XeOuaPruHBASPJk6EMpxH8kQb0Ekh1h1mO1EG2imVQDm7RJ0ewGgyYq7cGfUM6z
XGxuZMyrR0ELso+KQjTGf78ws0CBvjcy0qDwVd8jr8ElKX65Ua/x9Xla05BRqB3+
kfqA4uL0TpUKQc4g9NgqSt1+FBAdiln30OMoYpGTxBDwk2o4lr/Gc37GVUoAt3oM
CQACf9tdacm9B4AOVSW4S200lHvfi5DauHQ9rahN10HQNFbQOpZ8fHO2LzP/mWZv
LEDywab95CSu6akPyPWLH6DA4yR9VaDn5fm3VBmVKbQhWVAfSCVMnJjUI1WPvoDK
mbf79HCupIjEly8v/dLYKik4X8Riup0ieQhw14+6WC6qy4Flo6U1k1NBjKHXUscy
Oe/6xFlklq/Ii9wPmH8DzymgEsaRV+kbaxrR1kLk64eE67kIo0hKQIlCuxt4eMEs
e34bobx7tb7n447rIBriZLiA4rdMvrH+ATAbvTJZH/q20THq/GQ0Z4UehGA5J/a2
hPQRUghrdKnf3Fstgp7d6JxFkopnlSIr4klcKD6YZ2JxfF7xvGWUaI9HIoHedTb+
BwyB9ulpru5okURprEsgE4lZxN1EdajZjMm2YDQyY2PqvhdrW3bJmn326Wb9poM2
rc0j6MsSLv2sNcLhIRgAkn1wYNDQrUXG4V2aySAz0RO8HgugiZ8KYZ3QQydUSWU4
8hrlfU/Nb+SMp2Tn+iHIGCp46fkJNm4GUl3Ie6ueArwJbRVrQOmJXPaumgbqRNxi
QhFUtfhooGCNa4srhoMCb7ZWAYHL7XNJVo9UWOYZh+rUeyA+eO33irBp9Vc1z6fj
QeNDWderkAoHKV3Zq4rP+NCMUaA27H00ePNa7cnYSx4cb8XeezRJUd353bP2JTEr
FML9+ASZqN99XQtwJcl/7+a9+q3Qcb6qEiT8oOZYeg96/alQIQvh9mN/d99KGtFW
rye6yaI3Zvp8rWeGnU9kCXcJcR/mA8AfbTRA5rg0l7IvS1ZBUnKdD6cxOzq/VjNo
KRb6yq8MzJ3YXMTkbMlcFX44BYi1P02M3/J4z5PQxgaBm9WouPF5YbWyCOGXDzbl
bfSWJwKG9yT6TCInhKWOed573T7llKYyGyOnbNNSqRZTpPHxp4RhzvIQkzK6DWAl
XlARt/BTorfc+wZfn1Fw6QYebJpmVRlTw5pAqtNG09SJGyktTfBk41sucHAI/75s
a/33yFgR1+v65MnCB/fKahxYaSoS8PCzslq1zRmrnyMRPzKi+7Q5452L1JlO4g2s
i0V4yFouaqP6y3gZDELdt8puyUlW2Dd7Ss7tGH+H5VK7/lF8/LuJKrHmnBGQsDZP
bBuuXvojJj+DUC7iFoRujU3Hhs64qXsU8b//5uP5TrK8CPJlzUCi96t+FirHowvp
KP/TL977SaErALk8/Os9xA==
`pragma protect end_protected
