// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MoGm5kLySUGxQymgVHxttINOWdMCya8zWpTZRfz1ZL8AojqeHErTyan3U7XUaffE
aI+EDWfFSLZMhgbVXntdFldNd4rDB0+/XP9EmjHQYxMsxazKbRVg1ilpK82fz3PA
PWaBRPTnXuXreFeAe+yupsAoZVGDHBdStMuD6qh3unQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4336)
MQrms6CEHmhObR9zoQx3UXist/xpjUbHBOZOut3/9pG6DxlMjxn/AANiRPqWgWKf
wu8KDP6DXw/7o/Ud05zXbl0FbO50ncTn9UQmNHDKE1VfnojlhYCcBwUxbUC4DafD
Dtqg5jYiPx567H7WDcFqMp4yKIcy9F8SCGnEU84P7RmuHyd3IPw/hlKSrAPB01EM
s+WNR1FPnuhaR6dnRlxfdqSWE++8xhXAg+r94590dAGlDHjH1tMpsjcqoEoAj1qz
H6QU7HZNUO//DDuzUm1KzrlR6wbowzzCOFENvWwN7W15smgNuRtmgr/UQpf3er2M
+ct5Qlzy0NGK/YzhqNdjf0Wit95gAz+TuPoAqTcc6W0usUcdGSR7nKgaW9DxKVKO
cuDdD4ZkGkln+akpovRe60vdLWhg0l9SRo1KCqlYNKsdayCtVLQxWmknomNDAiSD
IIFwFY1KeadtIuktkXJMOmvxNdVV6+1HMwdb5zaGOc9Sx/fPKoG67QeBsX2ICu6Z
0PHUOo/Fk7bikxeRi+k+c8SExWBDSqKfNV2QR8EGg0xXuRO0toO/lguK5qjuCMUr
Io/rGy+2iMBGcsuvJMCREjg1NFLPW7hYwAB2NLi5ip1zrReIir5qHjW5BsMuAjYD
67MFHwhUHHyNcuO5ze4PSxDejOpZkHgGRd82shc6q1nPZattxsMi2LTkOAmYt22e
Libk6+yEyh0UFfHW/05gUtH4Gpk4q4xjB2pD4mCXTYw7HeI1GzwpQw6pqDYAZJuI
yIlcgy2DDvUHQq4akSQd7jxb0slvn59O3udkdx5H5VnF1hZLfwDUTqOpOoKX8v/S
i7lWR+XDTq+Zm79hlJnWdtEqviNLHym8GdmlxrecpbtaZ+aQ3e/83V5j51dLYpV9
Id1mpq7R5p/gljYuHH2v97QL4Cu2zroRwTNZgV6OA5rEG5ws1LjsDHIReopxpU/1
mZstwTh2NRNBX1J+Vj+0AZDDSXWS6Nl8/hxl/hsDPrV1RD/5m0vtX1J9Gegd2GiL
aLgtfatB1h6e8mlBZEOMrAvGf9FL8CCPmDeLjMl2vvXEZ7XWgctpFpWEkzTni8lF
7pqlKTxatsguTdCS73Kzu6GhdOGyM8hZsZC+a0XIMmi6LHsRSphHMu02ppYqsxD/
YGuKmd567I+5zCcyV0dn1J0LH7ItewVoE/PMGC9q61wO+t2E8VSQ3+rPnm8nqhpz
uAnsW9CROIIblTFuaw2kXfqsEPMxlhNnQg9FkfipvUScZJYmfL9Hz3Ae3wUtJdWh
wRGrIMKIQBInQm5fFE/wPPJREsVou8CTzlEqaPY448uRDCOYIO0GbGyfNaLateMh
/oXc/siZYpbu1RlCv6eB1kDUEdsvjsnrjF93NgCwgA9OUSSzsZhvGXniUPLsyEBe
wNF+blpDnasFZDCulZQUIeX5JGvqOJdNXwrvHTw9vH0HuneeIAXE4d7oPt2kLaUO
9+o0ZOMIQLikIYa3rFLVrmogX2Ypr7EzX2F4T9VgKZ75h9CHLduJo6cVYgcfZcUw
DHsz7AD83c4+5aS6D1G6P8UQqiW9xKxl3N8w1RHmy+I2bhqigeAuEIltxiloc/o5
CU8UtDr1O2CJTtd8toIyFP0nvwwFRijxx8THLdNk/abky7oG089xIoJlQfWjEqio
3HE39NzJS5qgloVWaPpuL/kSVaut/5oQvAmOXLuPVaMPYoGeRfUP4HdnxDGuRdNX
imbqoFujF8R+uXe7VHRaLEJZdWzzSPUpqsLYqa6My7McA/62ggQZ5Tuz/Pw4b1wS
DtPzwA3uB6LSdeTozINvM7ZMsquHhprqz/zJfhiVqCWPlP08ZzuJ2bzsh8WqS4RR
7H6Il68xjLidqFi2R8YvcHoPeK5wN3UmV0MpQy+CXFUyLiUqH88GLmkAXrUZhsBV
wTTuhNkjlfO9mt9ATrmFmW3rjXXIE0B1/Xf4M0yQR8MNVM+2zXNBIuosfIpIP51I
76qgKPe/BtfS/sUQ00KkKt56WZC2UtypFjGGakBJKEiFG9w+QhYs4G3MNjSaYf30
wEC8Hv2CCYL3NPSRqNcq14GRlq79XkL5HsPxNRa+hrgh17T6HxRB86hYrJRl/grB
osnqciAe8A9Nj15mZb//nFqbJesNW7mjh/1YsGsWkVwY7zerkeKuiTYiE7SnDZbN
h2WFQmriPJ0ROE7nKUP5Z/hLq+txWk1LKXO3KSu+7WnyTyfAVBquBmifpEtmvDFF
MYoI4CghIKZ++qwt94YcCBLjyyxTb5+BuiK7B3/Rt0OofGfLPSOSGgoolq6EchYa
BrJyD9e66I/6p4XsmSfZMkDYh48VLqNkP7oCUOp4r+cea90VIGHW642VMAQ7Q9px
Af7wtlqQi2qkak7Dw5uy51GMWbG2vp/s0U6aRqX0SSneINCdrWg4OcvOmRkEj3Rt
zUXGNt43XHFAEeblhqCjA5xviufBipLgkSrWDYSQjMLTkVQyJQbwaUkj/M63WoJM
H9gmJdKJeMLXNX8gIfm3ChB1k73aNACH9XDrdqL5uzi71L8XLR/6lQlp3Glxj7zA
scc0ht+M0jZ5IGQNR+gxloIyzfxP3TvUhCYfq7cropSB2w5YJmgnpp6qi1P+g311
FLoGZAzvfvbjVPawzHfUuV1Xry5oH0obwkSHvdIfgL+1McSh7cTAY+URX5cvPKmY
DsB1QoYRXID6frsia3BboVqxuWdh7GpOH591zPqvT8R7yN2gRi8k5qWdfaPaudxZ
D+w3/VDnd6HYcQkuE7LeQCHBYnBEv3QXRwSbShPQDCnjxml7jr7lEfyRD0y9gTFu
hKDch+oyqDruF4kjq1si7KQGSNpsREuMxfTk6vPmXQmLgebfMHyADTRZN07g9I/M
gHt7RPOhQdJlxXlvWhoBkRhepxuzrk0H43+OFtfFrYFNMfuDUH0JOMWNRZiCanpu
yPLC6b0sMfI8g8wT8I9F67CqSVeXlluvsDMdIxa9F+WRBueTEny0MXlanwkbKENU
l2MmsReeY5YBe0Jht/GgRxpkdtgjOtT8blWMJHDUCZ3qHtV3D3NjE7kRi0C0Dthb
Qp85bafdloCxQ9eaaU6C/7F8FHuWl/58vohl465l3LwBleN/Byov0j0DVwaK9Fm/
AfOXzsRQOQTaCI58+Z9oxYQTPqPJtz0szwf4amuLtsNGTdXG3HLyENhrVYAw6Xgy
SDw40yTkvvYGVFz0TUp8687ijBRyHc+FJQviOPNtIF1WhuaJJqS56COH6XZ/OjtA
nVj64gqDZ44kvHKDhamTiz2I4gRrrAhCLo+WkxIAd6d9141eruSMBOKUnZqO8+OX
DVQiRwMoORdgFGNOWOGjPfCKsf9t2Y30dWPtSLUcI0/JQtLqVun9AYXNphtGL057
/Xzt1GAu4Hm164MQrOuKQFRjfb7nOFpNb61ZyEVniOIvl7PlfmUn4c6rlTQ/9BRv
AZDR9iIyycyPqfJaAWnX1XGIoqMBo7nskoRk7P8ufb22b+Wx8NCwLB2DYi9CCXgI
9ud/H4froa9/PNZVk20Rg36PZMB7Ds3Tz/bHail2wW0fcBwxglI9/GWyMXa3mzNk
JKa9GZPsmaac4N2S5YE+n6W6Wq2hPtiHMX9IWNsrlkUAmn0A6PeIFQh35PTBnv91
s745yyq5QkkJbs1KIezVLi9M/cl2/f2zv3lrgmpBRyC58Gv8TTRnNycqN2Lb69Sp
zXGlStT7VIMowx9Ibw9Dp4sd8oYhZ8l15V4Bu5zWOYbJWGY036iV51Lkxz26QHLn
gDJHAVXf9Cs/6dxhujhZd3tg+tX1LLMOfj6tTY7gC7s4oNdhDc9CyXqx2kZQjoaP
tQz4zp++oHFuXcaQ3NKfpbmKW9jV093M7JS7X4ejwQ6MvT0FRmaWZucdV+nHEy8P
k4E0WJycGrW21snmRjuhnogCnDmdi1CXBY2+BlSG2Bn7GrcBN7T8tWiyb6tnm8VB
YloiWj8kiRDph4zlLSccPrr7keKIYSsGgw2xLKYxJhSr3p2GUmCTD2rx/9oAcnUI
wUURgsppOqThdrv70TtndxqgZN5sHTTE0s0i2Le1QKwKGXC1lPW0nmqP9mCzsO3F
kRnq0woO+n+Vx/mK/SEGUnc4/4LjLPMO5aRXEKbHS7AjaLuvWAoOYLZChlYb1+WQ
HdPwFlGbpzOusRuv7XbOwO0M/8izKNZoQ5l5AfAO+mBhf2OtOkk3hIXwoV5UWnks
4I6l0TzLEmxqiEJXkS9jaMgVfDWxZfCj7lHgbWYr9+HlFqpGc0oTjHNjX/fhUIiC
0yqbNHgjrJHX97Ff3QXP92kdLJPbJwSthLU/EOCKSjmgJz5Q7NTfc+ESeH851W24
AaQytvuYWLOdckm29VqMdytm4z6F2gEtKJc40zzCCvFzc3v2G7338Zb0f5AOgYV7
cEYIKk+NqhUsPzJznIQLvavaGVGjxAJx1UT/azueybcAg3xPNDyOzeEcbMhdhAil
97XHxPHqUl/YpoNJ+wfv3Ne/EfZFDlMVcvthkFVksAwyGy/vAzj3MTABQ1p7ZHfz
+FjC2nAU+NnK0Z1iWcKNxdVwx/mn7kjskCeOBX//zSRlBbu1MlECospexGIjZy5K
Mk9IPZeUOZ1z8fVLD7XfKwDbeZyjFJV2vSjkmIy7B6COO/BF/Bc9KxlsRBk/W4a/
IqFrL6C8t9m205ZMNq54wm/pAjRNM3TiZcq0BnkIR9FO0oUa8kzY05kzWbDShT5C
51igmLu7ZorsD3rWB/4jjxA1YYIvgVCROfkdp2vI3SSd6GLxuApUvfmisXbnbp8f
8kMpjpD1kC8pJnzgucaqjsd8e/BAhq/Hz5rWbuVTAPNFqqKhB8QVFW13/ikdFCmS
v+/ZFxe39aDST1ZmFwpwPPeZxen5gpf24FKgWPkrKevyItKkz9SPrgLr9UNp8Gze
pokbcxF3RggPZ60gcoe7F78iyCt4gL5rlpLl3X7CN50Ws/t5w9cVFbNOobjuboVW
ny0WN+Ic+TeKB5aIXE/WBcxstzXUSbL2USD3HiF5bn7bG0xTa9afyzdr7WQqPwbN
nP2UufmorEGli4iNt77QcwjWUTrjXi8uETrkUyYjiWX1d7pfAPtr4NNIJULIDLX2
vb0npy9InppLvV2wcNGxSKIxXkxWMbKlHabVjzhrMUNfB9C3MSk5CuQdzO+530Ei
6109Ms7+HjC2NFSwRNaHIkxGspsEd8+lJ9FUcWwGz5CX0W592PQmHAid9HFO4NdY
ncKHhHBDxYofcBzOwvoWDiuNvA2qb/b9ucmeM6dSiUe9ifgTZ1HgOMY4ipvvba+C
mQ3Z/kZ2XqNeUcwzp2t9Iiqa3L4AKKc7p1Wo5BQOWFK7EndDrf9sSlezORTBJsKI
PY3iM/d2kjzTVos6oNrmNyk2MwosYwjKOJ0tp3VobSa2k7p6zyVD3FPNS+qXwt4f
V11vJBFYfe10PKxD9bt27ynYi18wIcDVbaF9YaTE5Ccv/nzgNQ2FXz6wMvZxOsUd
WwNEMy2GxV4bgQT9W5LOFfhAr6GAuD158HgHxM9aOSd6lRUPToR2oVKj/JEeu2h9
OsnTAKiX4l13WNkEy1YIM4Awqq8i5AVIbfjJdhVNiBEkNOVFMob+hEUoa8PwT1nJ
mAVVNvpnwgFJFitcdr7QfJRUc5ylvRBF5BzPU/GrmTT7cW/oiXDhsRj5SYCQSpep
lio5Dk5elkQx2u8HTIIlxVdOXvvSl0DEnKnPK5hM8RbL8Xni6Po1STq8Mliu5zql
nwh65xi8wNqUL+aqJQwdaQ==
`pragma protect end_protected
