// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
swDj6Q7u5kpNdoAkB1p7XEKcq5F970gQWB3IoRqZ8Fu/RTJZKrtIoqtJr6gBWqyv
i5B6allyKccdvzMcBEcKdJBUMimBw65kx/KlZOia1Ng0rdSahGJJtOYJBeB3ue37
bohjQrwaeKdRzFerIZPyQ9akPpVvs17FaKumnNOh7cM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7264)
LbI9YuxWa8+1njgU7Y4gPMb7faGvxiV4OmNid1e+zK8bLfXxX3ZUdM+W51e+/t5I
RYPk9JOvsXxHh5SOOmZbC/z37uBo4B0Em81hQmTCceP+nZ+tgrHF6NQ5i6p8+iUY
QoTsgjfILr41I3SI3NaxLxuDTschz+ZrhkhcO38JKSbutNq6aL/cE1VmbgT+M2Zb
CsclgtuYVzi/IAoo0ToO+JyzVZAe0vSC1MBbHIVVji1NghBvNCSw/ibyth4taTAW
tPgS0RPS/+9t8k9t4CtltieKaiiHIvXK+E73BcK9Jc0k4908d30301gXDk2ORpEz
Z+22lieMCjM4k9TZb3xzZDoU+86P0bToV59RZGVOlkz5YthShpLz0MmrM2gOriBs
9Yj0y0AQel+AuWWya1StNXApgU98N34w25Utv+YpqSRpnpsGR9NwQjXw5diwlqdw
XUCrtZXeyJl3gHcZUfBZ8JXcbJPFwJEsZYCMXlRTjmY5OsBWKobz96lK1O/TUaKx
jFWbfYirkfvRCufzz7PgImAq8+TR9y8v8B2m2jUlydaMpdaMy57n0eVLIV5EB6M+
GuK5S9kEX2O76cqyoc1d+H9v2yEotPb6hHvIdNlN9iemeAvDbwwaADC2QGTCKO6y
KL5W+ZeP9UZ6uj+guFYkGv3HZyAuMYW9CfAxcqXyMR5Zb+kWOt+oZfzux42HfzAk
KL62p4RbCLPrjZ63DQOtuUi440m0rvt7+4u7E9V+7JVP81Mlkcgp0FXx5JY5sWGP
bdNWNij9IjNswi+u3CoBpr1czbF9LHA/mF/+ke6KH//1fUmzpvDVElTNNIPyEWHO
Dsk/lSIiz2HL/QizCiusTVNsnw+RQCMRcKw9+pmVtzXox0rqRtvRHNdpZYw3Y0Xg
vgd06ZGZwxwbsPcC1RRoGvCaFrwL1SVEUOEV2yf1Hh559P0Z0cmW7McQRnwLd+1F
iDbVH8b1eMIDlt7lrYpIuwDS439MOI+51T0dZNyyzJx/RWaYQ53fl//ke1BbRRjG
/ow0BNM3SNE80xR16FECiLsNfE+CYzFtdbkLv0Mc5BzhgiTy24iWDLDaDOVNxHYh
v+YDFRugM7KRP56+7CBOUWNRZp5An/HKfhkSh8eII/rO6tA2SUzSWvDUlNItFAUO
V7UkupNyCOvmdO2Hpik5Of2ymDrqy2l1y0mlXabyKJYNUG9C28/LtXILqmqOwzz3
IMNQ1CvrVuCgyfJaq+URykbm7ypEDKrsdzR54/8khLBijRDXBqCpMulpsUFrFppu
DqhoCqgPdDAY1Kf34ogCXy4kMqIKSNNeWeibffLJ378n1QdVBIzycBDZOpoK1mdw
x3zFePSqeiMBK0H3UAywknVqzFEz9pJbuxQqLjaEyYVnPMJh8MZlS9oC3YKJkvo1
9PaVeb5uHWxT1xBtSYqGoPNlyxgo+r+KiwctzDK0hUwfJa3TX4TEonoj/jSVjTWg
T/4MNplrBxk1xwk/klhR4TZT1ITjegUF8g035ZCAt+y7lhACu2JLermauzDaCmYu
q7fC2ieqzURVzyxpi9OdNUSnvCINTeSB/on26UrESnT4/XTDsdKIpphlDnXZ3jwz
z5PxHutNm47BNI7Tm2kQs8oN7YV3D7A67kLnf6zwoZZjAUf3tfvihnN9eVEoY73G
lrlnaT/pHeyuo5RArbAyU4UuWwlJSwVsFEyAVxg2N9b5SLBVOCjvEa/RBnVLvbRS
xW4/UFV1n7eVRYXnJX3xMd7OulKfY4mY8MJZPT0PD6W7efW0/aneSLvdUC/QrVaj
LvJd6eXmnaZ0uXWCiiFYzxpr/y1wgLiY/McXiRVvt4Af4lOWbhSl+pwLCNk20Wqn
34J+C3+iB46a7Nd/0YcvtnG2hhzJRlZfoaIatzGpz1UL+XJHSjM5phq5vFdkAv3E
6TB/rSMzslYhw0a0jDOcEGLFV154L+BxAqYDWx+eB5eIOZ6v/U749SXYLibXgCCw
Qr866KZVuzG1CWFica3ZdDptcKaDCpBvQuCAMOOpIgL4Ughu95ciQuhxm74KE6V5
XVTr5BUWroGG3CVn6NAlPMDr+5HeZbc9L04+qnVPC4A/vmEKwueSmjFxptwy0RH1
WVUX/+uQ2611pWKMQCo2VctqD9m/3UIwPtD7sMLeMX4x85NlxDWwxdvz2zKVInvT
7e2e+vXBVdl5f11I/YdRWOolY1D5sHJ7bBFVg0qrOO2pBN32RNWqiAYzsqO90TEG
O3Q/jDnBtKV+MTc1uGfytP30i786h8uZJPynmQRkX5UpYFeGk/MTo49ez4XffghI
S1qyDs245LpYTLr/abKKGxt5hwxXEQ9/+KAutn0lZII5XtL4NKAGRUuLx4HOqxb+
3u4wVzjmPGdyueIgwprZfeYVCgIfho5A36HF6ogfvNk0pj3E6YyFP5z05t+Clsi7
2G+gpHi53/qUBGB96lrt6RFTLOnqhjF0jwnIBTBIdnwE6cl8v0ZXc34OhJUg36oD
ZgizFwDAzEBNQ9AAZLzuk8OSZJvoXwTq3fzDr7RX8YVty0hFlynJts5paQsl9v1c
fw4J3Tgp1MPYk0PeJmn31LVJ/YqH/DQTEvueqSGdFFGPxY+szvREv9jXNPB+yN0R
aaJEIIoAyrKQScgRsu7hE5af2GZkZUnX2rMxhdHvq+pipCeluzu1Q0HqQiN/g4K8
Rj2iDFxjDwQswr2XQg987sYfnlPo1NJ/OxZ5ac+m1AtPzD3wqHZQZ9vZe9K6PHn7
44kHHdQNvzS6dSULQYw+3FWKFB4qtMrep3jwgG46KkfBJ3NsvW5fXz7Pw67n/o8Y
cXYyLVL76KyO69XQoEIpzWfjxFwflar9jqHPP4aAjbDWz+xrDHg058TKHL+n8yaw
+KEdV3VSNHN/RxXwFGQkys/sT/xpcgfQHFYdxE2aaZVx+/TP21yueC5LpQYBoULe
SfnohGWtCZ5vR4dG1dj4pmvuazCsBZNm4GBBQW3jh6Fjwq3/CTR861D8wdJ47tHs
8m8gz+oeiQFa3ZhOwFew3F3RQIMu8NmuSlABOq7Nx+cxGpJKaksJ8Mg5fRuDz1gU
O5Spwso11knqky+E2VjwLkQgcB5cU35k7B9wqlo/JQGFKoBCXnCcGRnwBDik0NoI
ze1iINChTlzk9pg/sVQtSDJvR5YhxBQ1vai+1qukwJU0yU/9Poql3xw3kk59Dm+O
KcnDYLFK6uZKox0zmqF8NOd266iXSCTE+n2PIzafKJihplJ9m2zWb4tLu2DyM/Bb
NRlBhbKGampZstSck1ypDaotZBpZlcmi+yejHC3at98CT5pQj11A0Twk7MPCWu7M
cLXEwK/kqrpyKGJH79PG1vneznTz/u5EQhmvrBiAQ0kXWDdxVhxOpLQSeVUPb+Ab
0mc6VytwJxms9Fz70dU7Fm4sAe+lyswBtIyxgyeNgoSRPsgMoBzluaT5C5vx7HZu
IAXisHA4GJytZfu8wTs6UIzwn27+oPQfCFrDh8nXGOSzTKDKV1ObKnnXuuVxrR6e
ZMOyQTP272jlv5AinkuHHqjCzkbntIvGi2eXUST/grmsBX+UxGIxhUASrlqDoTsb
6PYrO6R1w+iPdHpE6EM0m2hh9ROX36hKqKG810fm3+rGVds+zW2UCwpnH7alIyb4
JGZbWXMF6OiHFxI9FlGnmANuxU82rGHylnrJQhJZHjjwcP6N3lxATftExv8eULz2
OHSlYb4+cqPeqr8Xev7v1PsBYxx0kZ256D1g1Fuax7pq3WCFVm5u3RxUYtTjp47x
FI85TDuJmQKcQRQbTCdThV2zdd3oRlg6esqJ/SSHw6inJrTSPRZy20g4rEVZUb9i
IdaGno5iFtEQTSjtlA5UjR6jncNdC0Kot4Xr1TOAM7gaQU7YWhEJrjchCEIGLDsG
HJ/wLPlx+UysnmCR3rMuCXIO3FoyQxprip56E9s+Jc/YJOKHtUwmnlOxpax4pjvg
d+LlfaBVk4qg/NvQTj88CS3PEwRPfP3rDuZI7c67o6jw8pP6MfIYoO5gpAkrkVsJ
Md7T3z7RUnsRY1QYc8XFQteJqBFJy704nu8DH8XHfCcTJLJH2LIODz6HEgPOiURM
jT7n14IwU/2azxug7hQ9zvuEB+2EBgO+dayfAkjzAnrGyWC0K40hmjtegvS7UvJz
beoH7pLfIBpqrBJrCFhITIa6H3N4QbwHh3VJcgWET4pJgLe/I3X3FrjX3HqjPkCv
Vc+QTdKwuWsUtwBEwacriAo5jZvUcuMWVFeiUVub4kYWtHyX2BhanJwGcbG8u9be
oP1M2nEwqKlfF7JL1YGD3AYxDHZULDpHeewhMr6cB9kmEB1akBgBmJdCLNr6a+mN
fcQvjfOFrl/0ueowm2LqMW+3iJabc/4B9CqNRnKX8ZON8kSJQnBMO+DbAujjex/T
EPdtT8RHJ0WK5qlnkGYKVKbMykfsQS1yWn5wbMM5tOIueJ4jqA2x1gtU+o8hMjBb
9zrRWo2IkI6B18xttR4oVLBwL3Oy/PBW7FWjpLbcQbi45LrMqyl8e6C/oltbneB3
Bip+3PgEx53Zs03DhcYfGkbn/Yt+QvmXw7KT823LdWjmi39QPx88gbwGHAAUd7uo
TCcJjyGCqU2l96/cXLAy6PxuhVneI/0Rlm3FaK6npX7o12DaDwEn157iJPpnnDOc
pWHaIVy6K9RmldOcDIWac51WjzIUDAgEceKJKWFI01Dj4dfYwKed3p7bD+jg+0sv
oV54v5Co3SGBeg82Q/rDRs68cOfSW08ZjclKQcajJ+L7zuK564h2o4NUJ0ePvPwt
/eWQarwYWwnwhpkvgb7BsNNbLSwutmS1KSJTbdviWhaFsGv5qlFedK3r3jblzFr0
Gcbym766+JMzMRpyYQp4dqNz7k759+oNxkJN6Ry2DCF2fMCQy/DOLxg+dwUFY3Ou
Z2Tqb9mCiDZdihQ4vRH73PyeLQGtrgoN6cnMwdkstG7C8AlZSoZG5XBTUdShUTa5
K60vKcBC5IG6bxYEUK7+hKiybYdjrclfGGfNU4CHqg4seRsq6CIjlPoUm37VscSM
+KJuJe7dT2BXbVCqOuQrnOW/ga/G+RcX4vHtEx7kg0QQzOUBmPeFtbC03aP9t/o6
bQRhFnKao7sEnspBQP2zVsW2l19ymZrEgxiVVIN0NiOLIl19DUPBbW5mzv4fNwwu
d2fhPC1iabk7J4v52igF3+07zNcYUbjcXLbhjDdU+gt8dbYZZKdnH7jr/xHOhg3I
oW0Dk4PAbVM506KM/XSflaOFvxjWWFHuerPf8Wtpin76Air1r+vQZBgYCeYqzJl1
SujCb83IxMJdGy15W1BcRvLFFUeVIMGp6DVNutHPBr2LlMSK7SatoZA0k6Khrd/4
z0rn7zHftahoRd/JVCyiD70UQtlomvFFMjUE0Hb7ds52AY9DJr5tTwWaVY5N1JEk
wOclmWWRF4HCJqH+7GH1CNBQr2lMTYc10EJH/bbnnqlPOB2JT1AQh472vyNQsK01
safNuX/VIXzAU7fA5JrmF2UpAvXrezP8kx8mkWwnreQZM/3Djp7Dbe5Gpc5umVjq
60Qi8yLNAnbvZhUHkG7z/AKSNgxv15dxqou6d/wdxvfFzPZa9QN1yKGkN84S0288
AG+6ff6IjeG3xaAd6EOjfbZezg+wK6M+7gPfjrIKdugkpTaq6Pzztuji1B2N6pjI
gPQDwzlNJX/l2/rk9HMxrRjD3zslCRaQ7mAHLKaLZRoxvBa83C0EF9lW7Slofy+u
Y2+K2K157/b2S17N9GCItaAwYctt0ZAKoykkvoTFmzZiPWOthGYb2s50JXpQCybC
os1wyUZA3hxFSQl4STru+OOZxv6vjkq4jRCcetYi/d4UjdGIPKCfb2KlcBi9TsK1
uJCsR83phq3SBF1ruMLnpbiUMnxVoNLc8/UHc6S6BIoHzXwk92k3w1gQ2LFSpZrd
lqDzuCyy+jpjGHvEwICLdGSMqlICHAxvanFPiHhYuipkjzCETl9CGVXKAhCkZy5J
LgUowLah/9Fygj0QFo992AZs//gSyP45KqcGQEoXSMuAgj0q/u0rNxfEXSXHRSIm
G6GgffzqWxXIMlhHRhbs8TpDZwTGUY1UjRIZ7VUdFkXqLZomhPe6bOEB9sxp8bLv
CSEfoJ/dzrbVvRqCwL9zGZ5gZw8SqG4r/a20sOnZCO9V2yuJ8qllA6r6W3b+nbO5
7yFfW8MuxkXdT4yHpwt7bKZGieKnhjNubKy0kHIGRvdRV4blVDoMujwb+mxJ33Og
+BL/zos0zkqvg9eP1RcwCHHMyfvFIj9DZPrxRWc/n6Sl6fQ8i3xus/apTzDOLP7P
dpYg+7Ru//GyECLb06t0c9vRWXKQbrhV++1aDYVt7wsxa5bVEJJ5WU6lS2uS3aeq
hwSbMJAB9u27cSLlM3CP/fi2lkgF3tYPolDsy/TgnwLmwiIecMvRGYy+5HkXpKoR
xbyCZS3pRzqIJUHaaaP0NzFs1wCb4qHcldmmMdKgz9YObtaSNADr5xbPyi1Eb5T6
eqH8nsRbusL7TJUWprwrViaHn6tTEiFVGHJasOJzR7R4CFqMdkW0xyPOFcbD0S/7
x3FEoHRXilyJMfOaQb1T9LvKrYtaFOtwgdvQFHW1cSaaXNtiN13GJscDyCeKWJKc
suCb/dfyXhIFdchFJgafQTv4Byl/u8BJt5zXhqKg3HdNIzvklRPna4W/VOSwGRW8
13Wd83RG7MoifPZioQAkZP/+yKSL76nfz5cmFvR9rTEo0FR2Y8vUx7EeD8FuM/00
CEcEoz3WQ7N80BfkXN0FOzqZ1HCOi4WHHwVjtf/3teYziCbR1NSYhqS4kg9m70Rt
bGxsoXBNz6vXlMFK0cc0OTC17OnaC3qsy2sYhUKle2bThUsDsEsy+y/ZY2sPB6zp
vfuwZTursNGNbPdWQvtht6OchZwXOlZyuyHmmzaQukjEeRZzc39NxFH2L/j9oqAi
p5+RSgevco7WUWiBd7p1brIjsAW+a6jrFgRHx4TrXuAwWR1N6sTomPGOcmsKQpq1
vy2KRb6uE2FIQ0fHoWMwkNB+dheuH7xdbPfxBagC+BaF+eSm1+V+vCt6qdvByy7Y
7j3xElFMC9OolkIEOdgKj0XRLl17uoogrOGJfKwEO999+t3hYSK7HLiUwY56Q9+p
/YOLdxnFfABdaqoU0u/+sD5Z1OwgFLeiwvuCK09jZ0TWIdqEEE/6n3FFD82naF7x
RJA5+J9HhsAVN+/7VKuBSWbYIOHo47yHJrtDpW/Uvzc7/5ZMWgl4Q3zzri+KpWTs
6U6IzrrJ7N+EWawOvcK2+cTt6Ton0UG50ZBf26dwnmdd3i9VU/jRGer3wy8LI+ww
UdTKNS8HlL/qPOvt4p0zaaCBx9FtIo+tAe8yInEkxwyc+Df1B2wc+pJ0uhAMym7U
NT3fbNZs7+Dv/a8ndofuVPBpQC3ulqcqT2YbOCN6lYkFpc5hXt3zHgRNtdLk9kWl
cmwovPB2cVtcKrYWQEf9EYaLKXGk0PXTxsACsapnn38yZhsofrGG3YDnMnv/Ex2A
ez5kVnPmkK5tDQ+8ES6s3qR5PjtrLZ3twatzE71b0XVSQ1NKuEJWMsXIOH5pJIrB
jLX1D/9z5oAcNBFbvEneZNuTcLs5CoUF84GNtvXyu69ahmAGCzzDVrRh9UnXaByj
Ga5lOc3YEZ+NWxNPDSsLPVELFcBDS0tRYqFw8HOaS35jbnY/Nw4iVh1LW/joV5pW
8r5myvEXKVMbn7nreyDRDgvctN1EvamtNtoxPzfPoS+eAybIuoStBOzn2TmS5LLD
ZZU+c4J+Sn4Uusc640WA9damcbPolPbQiNvecisBViBFJPmiZge6FpjsoMcMWKrA
HfCBVqyB9omR0kasBhOEoYez0aTk79tZzIIWTofOlvNjmPcJ584E1pXbW43YPG4Z
uxTRC+UVXYU2QALCGIeB7rqvt94fh9xT87lHHTfLf9amfkFUA1PWikKBpAHMsFVF
xSF69XReEsx4GYMSqhKxQYjSlnEMKLOTqYaUtNCYaDslPOJgSLb4brumoejUYNAW
fVflxTn3nr9pNrnGUH4y8CyWvtDP93ciy8pr1w7G9mXa8ajAg5q9PliSKLOtit7f
91KX8L+eGLHn4AM7k+ZLshxlme92m/qbA2dI7AtbxTBVesFUPxdgfFoqUotil1Sk
8mReP3XdiRZbmfYz1G3dVFMR+DZ0XP024mWMgAa65T8lWcmFNRoN0s1dFfHYlWik
z3dGgL2YCcWevmX/XXx/K1JsykPMkipd54E7KHZ42FmzPu4nVlm6D6IPQzykYtMq
Ul/CCFrFue6b1UHLksXQHL5GZCL1xwmRRSIaFrkYluK/MrWZjfXU5acVzKPAhejF
s04X56hu64+sI7uqmbg4WmEup8lY39P/1AXxcFtkGBvfzhI1IQ1N5QvDhg3oA07Q
/PV1mELjm6d0wPB8TuCuYT3lOvFZtOtLbazxqwbkmfO4jYRxkyUwqFfwo2Qx/qEK
qQyxifaXNyFMqHMUbLxTlDHLe70ZyZyXodvx07LT/aHLSZSoyUE6VQF/ePyjyWM3
pOtGvC/3SfzUd4J65Ya0rDmPdq00tRKDNfhGdJVrXUN7CjTWlucXEMxG1gj1Z8Xg
w+svpI+QTLw9YEAxTNbo2ra8tf/ybj4LxSNXUE5BDqPAfSUH844OgVnMWpeFNcPV
xhuTNI4CAz9IOVxN/pf17f8znGQXt2QPzo51YfXHjjt0v2J5ahkAb2f7oYGUj3qs
tlz16q8dkd7gakMX6F4WJVgHO7rPsffN3XZ03Ga3z60fQqnyvkwlEmjUKTy9nKks
LsbIwvzxkW2K/McXC4weg2yk8/g4U4KVmkE3XIGQbKEY+zIHOz7m8u8QGbAuXq63
BXXFbHGwS9lf7pdZvNU15DW/1IEJoK0TqBxPJq6pGkqjV31NHI4Oowj7RyhCGfBK
Bk/eGVQCNgIW5tvK+mZwu/e0+M1ENKRccZAxoZHp0CbgBHzUCKw//QtM5J/+CpMS
3OmgBp+krizIC0l7tu34m7MP/0r9Wp9YO4XdbjCFdyC2IvqYR4vQedSGG3NqeGz8
RuI0k7GzGUshC37pq/IEJ/gMXC7qLcgTSjdNQKcJCIZIGk7v7e30pT/4TI0txBbG
2ru79P5mmVqnEHKJPcfg1eMUzsy56EadZuFxkKK6EirnlSibeYFS7C2zkwUGpOsP
i6pT31oHgqvfj3XCoQ4Ts11C2xougjjWjEnCPLg0ErpvVKlAcAD6hYlYa0BYpzv9
bewpS3gQ1mPPJBKy2vS45cWvOxno/wKUQ5zjX9a6bwyYnpeigFCkb4Dg+roA4UGa
mEqqiHSrSD9/qAnMNA+q9x2XrVc/DrY0onVq30karFDoejXAjPCZZO5q0YWpE/9S
pULm4gRElEZOME6yTnhK0kXBYJdRT1dLRzEtvAh5qGrW3dUHrxdDV6lcH6GMPehU
nY7uQIXy9f4IqY3SwmFHVy+4H1+g4Sut5MxzvSsit4eDmvWwBvH7Z4ChVfNBP5H8
3/Knv1kthi3UGp7SCTW69tMMQNUp/sUGLmgzcyODrMljLIV75K1N0nTxiSEi13sc
ZHWlH8/xXsqwEGmEdTLyniVp4r1LN46BRwUrAqBmVEVwy/Q9NqKv33pprW1yczcz
odAnfpLtX0pP4xS3b0o++Q==
`pragma protect end_protected
