// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L9LZzyqbW32s5a/eDlBntN+QbkF/KdKyyy1AGoo+HGa+10HFB04JbVkHkcHZBbp1
MK3uGlj3a+qGFu71SfaxjDb5sspQmouL0syu1JYe62KlO48u5pD1pTm7+iWTS4np
6+1/1AH2n6paKWF4uzD5a37adKUkKe6zfOfFpthBXes=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15312)
ZAjnjN2YwpqwIqSjG8mgE5YvBILpUZC+SAPFupcxHqqlqgmSzxc3AmrP0Z16pkDq
8gJHfMhr4hQK7wsB+FTPXgRSqkd6z4QrethU+6CO/VCliAvN+gvTQ63me0m5VXgy
BXnK5C0E92HC9hnht4u/ELgrQ6iVlrMHkEijZsmMSpPHJG8aOagDH3l0WfNSWx5c
qljkT/iUA4WOlpfPQoHoSk05HrkdclQaSJAC3TbQUQYMfn7D6JxU8mxkXNJJKwSr
RAAm8sGvyeOuecFSAvDUPiGz8FffvxnEPHIQoE8Wffc24LWH0rclppdgHkD7+Wib
Z1cC3fgqRakUsT5/SZU4ijqcE3aOvtqFOEvKUYYhne+hiOcIH0UFgXNEfhnamF0r
QGNGc5DbX0u+7/J8WQ6nIUndwb36JcIazeMyh5GvjRSD7qTUmmAaEN3iFNNuX10I
WtPuSXMYXYnsg6ldEhVMtruySTrc15TydBAdyYtsLRqPjeDTotLLdYFI3mtm3jek
ShLSVTi4Ig/h3zU6yrJdP8PDpw6CsJuIwifpIjfrXQzo+DGIbJSzK1JV0ybeXF94
BSAf5U5671Ho/SIu46dGWTAmHM+VBSTZrps/CM36gSsVBn7zpvis+7+spUDQ6CNW
w2MDoNxsmtIUjZNPp12Yu1gfnIL7z45weBAP6gqaUp6O3gfv4uz7RDayUxMX3s2H
29ofrgHtviGiHWtyEMCR/C6Mwh7veVKZ0Wi+LZR+VWvxbDeugzmjGcXEUDdkf8N4
w28sQ9Cr8IA/OAjictt2OBL47QZi4wNHR2Mzm7dgbOQsN9go3p3+MQv5YEKq4ONa
T8a6NWKto80Um+M/nkXwInVCkOxd43yhQrxDs9zL7hTJ3L7YIC8qcTtC1zMeLrSY
Zug2zyFKy5cChXUGtiCoOneoFHOn1wiCy1JllILpSye/89LtJwriFcVOqhmEFSdV
vS++Fc4SJf5aiTdZ8mNSAOSCgc0BJ20PTTTji2lOLAaoSHKa40P7JR2lIO3CPS7w
ii0aCV4dxRp5nNMegZWd1WLgYVFLd1Y5HyQCfY5LpYVIbLR631Pkc6uPVZFC7iBS
swHW9VK27kaaE3nM4CyY3CLxybbF6vQ34tsd07uO6+OzOu3kP2jT7QMplC52ndWH
yobBU7MmD1w1qNCYeb1vMj8qPQ0PFB4TSEFS7XQD+T9Ym85WVmnUYZOdGXXA17af
WutJOWlgmJ/4S1M0w13Cu9cYQnUu6MFlCaBHOKpJc4CKUQsw9aje065X2UWh1aD7
kAA6d0nnN2xC9sED3PCpdRDkb6R1B/PP2gi7WU/4cg5u1Kw38JrkFDaRobYvFPy+
5BWmW+pYsIPLtMGif7R7y/uS1eIq1JLuJHsOdXL0XK+WH2nTBtBcBnmwTgY2fHUk
FAlKWwVxgz1/qEASPLrT1Cdjx6U3k5R60n3ewVc+6aGCR7TvOiZF8s48/nYYVNnP
6RLckKL5uBCHACwHE7SJiOHCHzD/YkUAriGNGJXtdCOhzRZ13+Ep1cEVsVannk4l
wOWEQhOyCKGhSD1DwJgZCCpH6bDC4HonxBuRujuSRYKDagUvhijBkKN6HUq5il5X
aMfyzyqDMXiTT6+UoMPQFOlC/92lGGBf7+ysymLXX/rAMud6zagACG4eTaX0bt2z
9KfGIpdg7wbbcY4FSbjWY1ecQ4dZEXZIkiB+OLKn/iyeFb7KBcsDYz8bcjGYeqVf
wKCWbe+6WaHQOew4APMbhwxkC0h9IerUW/C/jX1v/+7++SRHyC669h2Lpro6jRJ5
iY4kNJIJL78HTN3iqKNaStkswBd2oyznuYEmPoD8FH6ds740e2eoMl1P8ie6w9pg
mkL7HF2I1Fu7rCz1r7iQA4g6pSbHG3PS9PZb4RDSXKN9NIlGMwlAJTBedBodfNRt
3LmmEj0j8U+QGhdzJH4So1YrbdktkXZ8QM10LC1g5I3tluYi33FCKg/vdXf0ODAA
q4UsILlun4DPlII/ypcAJRz6QAGuwiH6V/0gHLwvDOWPE2fBNGlOy8MGE4MgiRgO
vqsK5Ky3q1DUL34sAoEmRG/Kv6Iyh2PwJIpjoDgvB+q6rVxEPCNI53r/BRXToiR7
SeEwKdWW+QYzS8Y/VXoTiibndcAJFBsbsVypvkF3b2uIenIxC442xDrwnRM3wHpL
UL6V5uNFyzbClUBHo9A/2lrT6e23NCPgypNEbcf01qr123RAlN5l//Awc4s2zvEw
H6g+kAtsRiTA+2fZSCbNH4pUf5kH8zIUFxXQ3WOhCuAdd8VbhIAurm85VSK6jq6d
5BYOEM+Y0FidxJ9aV0N4RG9pmy58aaDGkrEIxbeLXYIziODQVYEIGcRKTN0VxsjF
BEtk6udXFCYjs3SNzOD4n7aeELB/4723q6dzLJEYE+Hi51NsDlerzlSStsvwspN6
izLIa+wn4dNCjBvglRVHErQxDl5PxyKKC3tFziMULzsUq8cF4sNEQnnRrLA6l3mh
pOLqzH+nbXCkoi1Qyh6nVOcaxfAlspNyhVttuVwoeJMipNVPkTNXvd2Zim0h2eyg
E83wFWPd1pn5r2dUL6KAM/uN9XZteKHMPXjUItyNFz3BLAl70UZfiAe71X8MISmX
q/kdFA36YyE6IPeCxBw7R3op4US+1DlNG8vChiDIEvZSAlvnFVNAF59NZVyDevF9
ldCvLKlXvjhTYDUu1tfLtDc7Q3lSTHPuQWpgwxEc9fCYPtHXx3di3OhffttLPq4E
+riLn+W8Wz2+E3c30q6ulE9RExRcbUypAXJOP7fHww5SCOVqkS7GRNcivXAhHL//
v7DzZVxRDpQMz9C6VbUSb8OalEhd0JBvkUmaa6BBxgzbt6yOg+DOckrJ0KuNoAlW
tKOOEiiNu9T1UqbTvg8PLKnzCwUv5gw2ni2aP2zmMcWRGWHfhV+aSaz3JSLxdfzM
JJnleA+KSkr2HTJ/r5KhxPNjAchVjmwQynhMZeH0vpaewdq8jmZh00Jq/Bl0boS8
PGk0Y1HkCd7oE0SFUItMOpYKxQgYIVC2m+YEv/9fxFx1S8UJXhBK+zySA/AaDEI7
wnfzp2SgEoLFEy4njIrquiO4RaFHV1JTiT1xKtgQmSpb7+Wy5KtitKYoHtg1ts0T
gtTwETGUnzAIC49LqJB61ivPIEQpe6pvIDDFRaTtArC11ck+SfYA7eMntkm1HEjU
RQpktSRUf2SM07Lfe87ji57E8rKyO4nvKZiPaYf8L3YRhAohq2+FeagvWPdceeUO
HZghtltsqVKYLQ7kVwluus9Hn+ECzfo2AtZxdKB2MQHJuR7wI+bT5qt7mpOYvhtU
Pvquna1awszKEH/wfrpFK3Vv5qhzqEDsoEYax+k5z6rxgFAWZsHLDqmlYEseF3oH
3ovYLcvrmOAVFjxjpjtg7pTuT507YiMXIcMbzBZj0ScmvYpFaydcvYGoL/aVOwLc
ESo3HPP+C24IfkO73how1I6Q5Z01wR7ehURHXciYrk4yBubErcW642iTMYgyIRmp
bcxlLaU0VMRLspllJUuwuO9U2Odg2nABH3qG2dN7xMtN0gme+6u3ekvvk7liBkEe
quGAchi8DxQc0PXRs8eHoLy53/yjhJDl7pVlehtG+3o5k0ytfeJqGPaqfX3+MCuf
MlTkNctbcULOsBQ1nLcLrBZ328LaWDh9w+q8gvyeBGTUUbp59EBjygc6b8rFPmZF
qILcQ4mAAYimPj/wGWyLCnfxgF4dbQeG0Dp/zGT5Ll9zoVbBR6hbbXCvTf61K4aD
Y6d8S01sKGkOdn6xrZCyeiSRU+v/cn5OUh65w/1ZqBkC40YYTmcwQMUp5b5LeAN/
PI1Mxt9PDcjcrqd+eUdCjT6yrYzdrTmB4yK4PaeP6Fx8TF3I5M2t3TfZhK1bnG1k
/bIA3xygSbzgxw9nMTvBVq1iVSxH11IRo79dDMFxuYQZyi7YjMHSTPp5ozh5KcDr
C7QSoam7pwAWzhDgr+UryNwusDdf8YgSGlIQ69LRSIygM1Hrxc9VizTrlGZ9mj44
4BiRkEq5megmIhhsCGIOjx8rJqG0HvbXHKkbvomQAi5VVPd7C+80qtnBzsMzCMjU
eqkn7Wo6EI7v3Qz0/LXrUyVfqurgDk1q4/T9pa/5kzlZIryp4AJowPWHhMgHnNPV
LvoCQLyA+hzosCV+d3019AVVH99WgKgkzm6VWD4iwM/pDvhM7RlxUcrqiMXIEhzG
HPlMcDPPrYsaJ0SAe3jJEaafMPxs2bw5WsUoWQEudJQu03CM5Lw4R05YAt+pF3QP
tDnxm/NnyGvZeqJOyRLT1Lt7Le/eoOfpX8zL9Err1CgQdXPTT4W2V5UiC/whSQVY
qahN7g6e8HToFhibuxk3EJe68HbAFVB9KvP1U9Z6diCZzRae1JyyJPnkYrL93W4Z
hQSw67FqinikFcpcsgv+wYmuAhPGb8riKtxuSbIPmjS/Fiq3PukAnG9BKd2bQevR
FI8g73wpy9vRe41KQUjrcevTNXM+UlfjR6DtjVZLCJsSPiew6jWYE0H3q5FRQVlj
OamRMQAx/t70Ap5Walc7v/TNSL9C29Rj0OaLwQt6AD4bkVojGoZO7snqqaQZuYDQ
05GTZsZTbSc24nelhNxcdeS7465DxKPglO536lmxhHf7HBs3TnWUGwuV6OZ3gDq+
wICIJtkw60itk6dJf9clMkImI+M2EqlEUFTih3UC23SlrK1AjnGIEj4P6drDHwo0
Yjtkh1beAguktBqz61QwOUb1zwNW3au0cp6yKHjWyC+LEWCsSZ0XZHQ/GQBsY9sB
dBtWFukB10gEhwJ7UId2a7SffCLI3lGGTburhu4mXRZ8KwQ8+46XOLkgLfrhSPBJ
qTgRI+5Z3+Ji/heG80YT0l2P3XN7nJrDzSJGQmcIbpnjMRyx9HuK0P+vHPi9hIi6
ESakmBe8frCnx3uAqFtDZnHI0V1MfY7p8MEnBaZC/2iGkGxNE/j9DX7mf2pRaiXW
DGYV4lP1R8urNARvZjjXfqE/NuDlhmPgFHSDAIEu7EQGARdNzFo2TCQf+ivLbLfV
kc/e4bt2Txy56nvxx+KIva+gmbzAn246Czh04J2U9zRV/ZSS3ivRY7KKppPQQjwc
k4cSKwgLe1YneSMHGny1niho98cTjdpZtQ5C1YRez92e3MfanASdZ1KHoCW01zyu
iNqF1nwid1KQXLqiX/iJ8rZWQGYd+DFr3OgwJIT4mfzLFGPnCRYYhDsPlxgjFJwo
0HRJjHjYA/ZBGr0Plk5vJ4Y1q9Vi3jNkw7Lz18DuSz0JgpFVGOHFTDPpQ8q8EBLe
9Z54Pk8P9JUcN/Y81MFFyQGfbQwiuCA7hQC3jwJMGIAp7v8ZJn+WXMneoVfvLFfa
ECNgLY7ivUY+aqtWW4BM7alRm8F732Q+9DjpD4jRRXU4sitfARXmzU7PkhENodzC
mXDamZ9vaw7wzeGUf40nSGqmr/0r4+B1FunT53Q0AbplTd4bQqgnmrGMSm+W1dbg
Wd77SmjFwPhkMuLwlj1hWsHyUS8lwlhIBjZQ1QY64lYR8+ESv97bHAxxqe7eEt20
ycPapmFMH+IzoLC3+EfPhWdVXzmrfGFEgkpxtr6L/3v/rTdROvQZguV/nDIWWx3U
c+xSbF3EAt/mfGllKip6Azst8O2Xbz6Mi6xscuA/vJFamJ9EvsdaBS7ct7HRHJBa
vE7rAd7bwz48PnTreJQvCwbeETP549j1JWQG4DOJ09j5fklanWQa1yNBSIuRIhPS
icOIsorh8JBTBf3KMWsJ7QzDJ11+/h5kHYRwcvpNTVpqTTqJITO8f2QjjFhhIwbG
zxDcNYB72v5r6GzcSVP9ZLyfP2NqFXk6AMi8apfZOTiIWN9d7ls+mFXU77kEoHN6
80FTuqVGGjKWIOhxvaYIZhtFwDiRSAZQs+iEiI/AVpxuuOY7xiql6jjKv8OVeS2s
MLjm4BYzG1oEb5ifZ52be9sS2iQ/cBayKgMUUstGeLDdXjwON2gQQiNf/Rc2ODjH
t1Wy+v25Hgd2kBM7J6gBEoMsYyk2YZeBY+pDuz8epcKkShmuq6ErEWljO/N7DlwY
T2InCdL03gIWLzFGOKiSP4AXeqkonPvj42KKjQxqIosAhGIniC/Fsj1tKhs2VeZO
pitdm2xdSUSbGe2b+QECmMPp9KlN7Bd84vneyJUAv4x5wCWnNQyW+9dp6tWEUMt1
vkMQrIoR70k0V3DApys4mtDg85/FvT0xWtExjRfQI62VjmDM+L7zlSJkmAfOVrDq
+d9qH8OD9Ow1Qzwu1KPaBkd4s38KjqZylgZJxJ1W4gv08ZJVXL+Uj4r53seYu0AT
50SJRJ+2I2Uva6fPeamGHM9uTvRShLjCxiQ155cINNt4ScKHYDu4EBBr4cK+lTag
5SL9jZB2ZTKrAnRFocmmPxjIuZ9PItBw+WvfFh22huZzEvepMPCeP32N2NG116Mb
EpupX6DG3gvErxzWDCjrTlLa5KHMHp5u13PyjqVez6GzWLdbHjEeaRjlUJAL5V15
1aDpiS1ZQXgZ6ie/m29vpGJ3ZeyK12tyL/Px2Kp85xJeMnmKkngVvygsduEGydy7
ymXtSp5v7dyRy9DFY/YCkhWhAcVdBVfhEb6lQM4lT64RiwSn5w++qjnmkJnLVC4T
ziTKuuo3pz8YjQiR18ZBiJSlBuWkRjTEMh1PBDK9WG23d/zV5AD16o4l8Yz4WicK
72tBfo8EGKuqiYcxizPllKepLvvBOnV/ExTgtkYZTZpsatrQtO8OpCdlnGlpm4k3
7GYlf3bFP/+7J046eLs6Ex/sXWl32UCvKv+QhIM6NkoWNvm0vzOvuHvJZiNuoX3V
oFFdLQzs7UH6t9uvgOiq03QWDBHdAeaKJUmU32AoFhyqRiSn3gfuONnnXQrkbE4+
Sx9KpjF/eKyKPu2R3NEd5r++hW0rra0R6rlvnaerJTOKfUJKGF1AwF8+rIiiqv7q
u3mzYVIbEIjPiPk1shV+sZueVU9SbooKXVXiXw17y5DkRiN2FdBjrXGIqcA/vkno
EP2i6JS1LmZQb1mbX54t5XS3cjC9JdDfeHaqhp1D+voNdz+PYLiVFyEjVdiLnRGi
/aDaYvdKgyswEsV0oFdLOPdnG5M0cDMXH4xSxI/7swhyP5uM7ahGqz71Ba9H2Mub
976wsJxqs+3DZeC8ejQG4xoH/433Bf49v7+VydirYRJxb5Zq1L5yoiUwFUYHJgcY
fBK64g8z1xgF0//cqk9Uro11toPkhScjeUHXrms+yH507wfvjhRH74atSruoTsIc
RJLLFjxyoBT72yyaLDA7ouEY48S6BSRVu7W5UM9SS5ubDDnWm/0/YAxB2bcSO+Bt
hQ/MBtmO4B5x80DThHjeud84T0r3dmU04pEiYCsNOR7mUjmwHFkrtRs5avVE0EHk
kl4YHCz8bGCxBxE5QHlkFn7dvpKy8Yxezb/S6h/+F4m1kV1MTbZ3H2KrRC+8zMJz
uOYJW+cnF2OTeX7TWeACy7MJZVLxnU4n12h0H+1F3/rP3Oxp9+utmmg9/INksvun
yvM66KOPu1LqT7wN+hUdXWCiY1OR6EOr4dZB2OXBUecC3gTYt0clrqE0Tx1DOaqW
sH0uxrhp1UNcLjrzhGLVYqaHNiW5yhzftKq41tq+eyvxURdZthb0sc3k1RaIzCIq
XLU9vSNNpioFWMg64t1AuknnNoEP471EU9gmimL22N5qNgQKI0DuYgc5FZjRBqvO
61QubKZm5vfZ0+DVF4Hz7Hk39u+GoynqsCtRFd08N9DqnwGsiFSWJivpnO9hhL3g
Ct5A/olU2J3/VibxcdZSbZr4meN0pcah5LvoxzwIEusyR4SAN/bPtrhmwEjOw86R
c/EN9Nt0UmJPAxVZVNAR056bIMaSqf7lQN61RHJov/Z1Ngnjg95i0kg4iEFmOvMm
3Fc/mUvPhOD5djtS+Q0mCKPGYicpQ/jRPOAm5HW8WXWrca8jwIA4FhBvdNPSVhAE
BqxRK1mc+BpNCNk2MO/lPDcSz92AHVOPEQs1DAd9Btnwi08mfZ9dL5vlWPUQLHiT
xAjVvL2qV/da6jd0aFwHhuuj+XidsyfOfqOZkthu8Anneoj3+MTmg/rHV3mQckOk
tmH1v0BPIS/0Xz3i6CiFJYXcbVpZGNgWJpvcVjOvPfvaTovMZFB5dPtwxuNp+2gk
IYreob5TNv7+1kxeOUW9nsFc6woZ4aAhms3ws2JYNX1DAcX5G1ESaiz8eIqNEGQ8
6ByxAYbfU4ZhmJRTQYCcrF89aniHrsDyqOyCIpt2gSOxd1+3ISXd+9R0qxKS/BNG
VhknC7UUJEItLc7ewjRKidMy5XUNOXqSU0xxGvT+WbqzsRV73io5+rc2UQQ1cvBW
R2V2NgpiH2Ja7M9EpoHJtLcwaN7yJyHmj8gOAH851v1PXz5yyR3DDIF37YOx8IoM
ncdDwUj/RQ4efFqxrJeMcHbobkC3QRiwIhSiUiJ2Fn0u9FkOZq85qHFBlC6u4IhT
x8FGraZmNdVs/AnigpWk1xEjd6KQPsam0sI5FmqF9OqbLLOIEk+moPuR1p7zAp1z
0TgpGBMkZNp4qdpa8w6BvZVZdY8hMFoYkqMo+L7K/OoooeewYbZjJD1D8+S+Z1/O
bdyX3QkvoNpaXSD5s3xxATPDOIIHg01OQP4jGNCuPQlQE1AF11WQCK06Bz2yji7Q
O6BpAHMQCgnEGAGbyVyb+HJ0qZhVPbprQNJejejXNHc158Z/uSe4gv1iraw/rMr4
EqIRyked2Prma9mmOVMJ5Sebxyu4AkP+9usNEaQWGkEGiWIHoX8zBrCsjsfWz9O7
5KXJbD4QNvVEMOUR7rAxX9eUmnTpBkz8BEkPQg3I3HMDjYlF4+Ps5a3AvCgtxy7k
7XIGc5iFHepTzBEMqyvxiCDOh4Bmcw2jakmIffFKRP+5BCtgQriyez8CEDNaNwY8
zl7Jcl4amChO9i6bceQXtX1ChgrcS84LBKtksbKpOkRvl+H8qmni9qJNM9sFY9ko
rOp4JJQZUUOkF2MF0PsJ09q6lomVFHz1djNi5YIRzuSWLHhGzXCP5xYLCZqsCYzs
ZGI/77QJ9wHZKxvY9MLkrLKSK+T4EGMxuJGOgWlfog9dX6Ks20gmnoArywp80Vnn
1xMQTXbFLMFJn2UucrpQp+WE6Xq/+k6fLqnEmd+bd4f/e7JPF9dWBOa8M6Z0IF2C
EKeX1zhpFekMdM3cLPuMqXzSLHDBBqID3cJLcjthWNFyFL234PWS27109FTwYcg1
BzJgTJAROiuJeJFD0dnFQ3voKq6ZyS6ZUU0RPwpyvUsX8RdQKGGXDwDT9dI4s6mq
6Se+I3repxC5bn2m5ICuHr82Y4kfD6whJKMndHMlvSmJ7px7R/9WkMppT4Ij2wMT
E2p7ci0g/nd5xDkVCwX9ddIYhBouVwbn+3x96RIb0WiIIvYgnoFed5CfbFYCCr/O
/IGgvRfg7NEpGfwGkiXnJ4AwJNRLowyzXFPfMaTF+6vcRtHcIVVoRlTdhmWBKF5G
GXa0QpwFy69FDHTwdrnaM5ShI6r+73135GSerwAlv1aynj/9tPW4JVCHCfBkN64I
Jd9Dk8dNBI87+NfBzzLarWxQ5mSW3s47dZ+gCikGpE7Wp3sxMqcDv6mwGcUz6kqg
t/iocvdVdFpMWTswL/IVhiq/RkDj+CTNcbypor87xZp0yeFwB7pvxRA0ddHfdgKb
K3h35U9HlxtTJ5UkM95C7/nDlqmZPI9yW+PpIkurAMy9m/+v/9sL0cjHea46nD6M
xtU+g7V3E0oydkiLvy+0LET1spSWZY2A4qpfy0m6k9UR6xR7P05pOO3JB3+QVe6/
ifmbavtl8qX4YCzpZv1NZeX8Hj5eoskyUGBTJFGP9hoEsDu507favMdyUuHAgDf2
On4sHGYGPmZ41OiZUx/rT39ktlIix6JMgtKo8C4gJIlChReAIAgqg+ZgI4mJdJ1h
tdLaRrbrBP7vWuvuN5G0/6kn0RQZkYqstyX7Uie6Tlo+kQG59CEHUvWgQ2mDU952
XViCJZJa61ozW2VabL8CvlZq1KnHTP9gyMaHQjnqQGmqrrthKS3/qevNQ9KpR6+Z
PUv4AVQO7j+Qz3cGfFxaLoDsZUQ7C8rqmc83ay2OIUiasSKJyqtGHqlsQa5HBqfu
RkdMuFXnF7Eik2+ACtEdTHIu908me4HNVgNvszo77NbTiLMAY484pkn8RspZzK7l
inxF+mSVFdLoTDKtQXYce9GC8ARChqQDPZdUGUCz6noSZTMrPzxsJRwlKIfC9fAs
ylGgDVs0OGZkN1TBpFZ6IdifiISXfgxHjZa5vtlE4w3izWXy4lDziJ3Lz7c5OYJt
mmhWdeXvrt7Aqp9ag81vjDb9TV8YwbhFRRiOjfikL0D1GFYMoodm54/qWJ4nXZoY
qPbpFazRW2CG0qgW2b71Hti0KlOanVY256OGkIeanYVzP65qfSjqtKnmFLWkwmlm
+VzEaPbQv5YJB3VP2LPS9O9tAD6iApxbLscqWlj+eK+gmM3Bfu5dokZ+27PaSIR7
XwR7ZqLOLLVWlYaiY2Uzjx/V6U8K4r708cXHdQGote9N98oAkkKujZ/EDLB4OKed
cvVUhV/aWHVW3ggg74b9oQpsNsXqY8pYohi25kFzJ283waZivKj1Sp4vvyZqOR68
KeaAMo9SSIuvgp+mqVWDbDdghSndyI3S6qn+rPrXeXQKz5Bp/NK73YvvwoiAUbPM
Bv8nXDf5uum0mfZcuOO5ZqkuNd5TgtvfxHkExdLJEbDCx1/tq7M2qzY0n5FmXdxl
0fWdkLI/oIHtXy+jRa8v7oCAKG0NKzfvPZPZnELXF63q/6npaZpK8gZRazayuU3A
eJRmdqKF3X3Xjx8wx12B98iMLXq141p5VdlezfOwVOwy55+poSIKx8C+D7RffcRG
qASW4VjrBhcEgJ8CCTYEunrEQkTcKZzRjAGhKw8E5eTZQbj7sG3lZitAMmrj5xXz
KKUrhKH020a4uofC/fvu80zUUdLNN/CfqzVync3vbScHi/G9SOn4Q7zryXmkAcP/
bbVdlYgVH5z+cTsg3Dp3jdB3svi97jzWtv0YSWEPjBLVQ1JUi3MkJ8KK0GE+U4Un
XqOw+GxDB972aJ4qO4W0LZGI+6bjzU/GmBFZmQ4W+7mNrx7OqLGWnEoqhD19Ndnj
QntKrHK9jWnVNp5fRa7rxRlb3ANF3VdxZaDWjZ7/K35hhlfTdxN3ZMmojpYrp2J7
NNMid0NtTsu1hxhFAgCSG5tBOQvUk+p9nQm4LdA42kO6L/LTq95z/sfiici5TfmS
QRRXh8aQptVT5WmkKQSeQ6PkrQoqU+gc7p0uJTbiCjMyLcsZH321vB4PoEr98mR6
ftFTqfiXArm/ODc8lE20HhGl565HNvm1ud5krpdP/KDoAoEIkSjM01qCvmrQZlN9
z+NctEVU5a+YMQSYuTdJ0mgHD7E+bPMMY9LcOxZOSh+MQqSyLm/ssyQu6cjBv9sd
PZkEsolM8LIHBo+Rss+fWFgXqtAy6VynkJ0cPisWcys+GYuf/VG8+UZDf9ugXNLB
yDuSEaRi3mvDu5cyd1zQTDerxdWJ+Z0kNauIxFJzK/E0mEZ7tgPUHifkKeqgbbYD
6f+at+N36X1Lar8Jg/bnFvZXcYrAFq5WYDduzuVIGZjG3/a1K75aSsfLcM21EK2c
p46c0PuHz3KvkdsIT/YrZiWJAAfjgoki9LmP8y3Davq6YdLFpD6C31CfgreaNaXW
PKgiDhbNOGIBzkQ3GDKM53/gkj4FjoF0gp6HrrPizJMNEVk04JXAtMm0zz9Cxjve
dpoh35kgFkyJXajTCmYg8qYH7SiUI88lMliDB7mEjh4r+e5xUfF2OGxxhrMop4QD
+BrVRZwmFH6wtEo/iHwaBm/8EWk8Io1OUQuR3nM4QrereUzPkd3GOaqwMBfKwmdz
514KbMueO2j+PyVk8PVvqqsaNE4mKsEcy5Q07qze80ySvYjnkcryeRHIdpTBmpJI
UH+unYqY1NOJfQRR1egLlV/VnruTYa13exnZrRx+b4Nw/Nnm9YXWCpCkSeT4ZBPj
6u2r+sizIB307r+XZ5qqrZu+cg3rsuXE2piBD4H5FbgA21NEKGMTqvam9ssHwDW+
p3KQ37qDyyMXWm/IfTytNZMtWa+Aew+IhyUF5do3JbEjWwFvnSD5BrLKFnF/AHbu
rmhNAxba/T4SZoiYr4pUGl7TG9hVGVvmpGjcB0pJsgfoUrhxSz9/dVHztSGie/gU
xXB9PPCVijTyNc9VT+fdjC6KY26d4SJZjaNPO/J/pKL2tiD9HgU+jedYvsV/ZnFB
M9jZGCCD4K5PNII2L4qjQeuCQEfpnUv1fG0VtCtRHE3U8dkoGLQjdGbLSb9Or+C0
K2giJJeRVzmXQrjF3nGhrDsbcmW4qQfaT+O+w7U7IjsX3nmBzmoR2W4Qpf3zQidz
JU1zk9nEqRlPhXlHzn4C3k62c5CAU3BoVZj+K7wf3b24saXsPF/YvOjPEWE7kCwJ
D6aU2RF4o7p9UaClWpdKCm7qVaGBpjP/rc/e3yQG7J010b5ngpc617U7YSHwVm1A
Hv9dM7ulr2p4iGJFu75nKBxp7Lx5ZAtLx7mGzV0YMoP/5MTDbUQknaNiDBwmZ4Nc
et9m0AHvof2E4Ec7QmdZC/PkJl8gvI5R8JUOV6C7WabKBpdQvXNWq9mNuf3lpkq0
A2p7LxufNOviW/N2jtymB5yMo10khJqsRVqipSgdeuhQJswnytSXjvcO1rjpAvv6
rHtuW/1nPEPaNxueWh7j7ydsBeKNVQyFtGtjGgf4YfvS+LM/JW0Pd3NerMFIA+9G
HGPY6D5oAXc54rbsA2eiRLqR3AiYaYKR5cuAl52RqCMBCW1cTVNIozWzfoGJUIQP
b6zDBOskmr8aiSwfGuDpuNpQoner5cp1ZP/FMUrtvIOmIDQbCyNl8xWAqvUH+Bfe
1Tg7USLl6j0F8WXjmN4FauQGpVYYWNTr1R8syhbLhbxxOPf++DwwCbh1YdENybBF
3qKG13MUr++rBVOZOQg3I+Nq/vzm6NVBNbm5iG4RrPmY0ldtQRTAVPlDBaSEpxon
WzdfGrNBb+qZEneEeJ6mI0GhlCacGi1rfQgN3fnFBIBCr7Btp4Cxc+SPiFNOYdxF
coiqdVS0vsy6xlsjkiZqZWs6h8LyQMRbexOgBkl1yN0TKZCNwoQbAx7PpzyueyVs
9LgQ6TbFVqc1cKIBKX+JRyGDcjuw4M4ljIlthSaDAhaw8JEVP6UUYM8H3R+FvJqa
ZB6fX61bOOyq9iKnTnvGWwh2ZfqHgVSKW3LboWLa2bhQqdu8YmDvdygowi+ifRtC
FgaYFXkCTRa1nzt9cGlnyI6DnH49jiYPk0eMc2AHO1QLVGex68UBfWXuKHUAEM7B
aDEGyNgemDi8nZcI3Phd/rQJB2+8thpV6wkTErAN4gZlQZtc234sck5xyQPu6Qhz
RtultTG9ARYR7lM4pPUNaB/kZ72HBXxqJPv72D6rDiSU5Bfv3xoOsGKzTIvWvj40
JAjgAQIr/Fc7YAk7gzZ6DZykZKnZ56oQ74IOMX+391BPmHu1nQddkgeEsF2jsO0w
nm655s8AQZEn5bNPgbpXNFo6Xw0VGwyx1v48r0/zlgjXD+GfEmHH3YehcPhMkGYo
VKWwt+iLySG2FtLZ46fq52IUz7iFf3/yNWi2kHoFl92Tn6JNWnHpaDAbZUQde+RG
c0dPNRJiEvl5UhltioEIx4I/mOLzm+4oQwwlzV15AQc0yVYkgo74/0Cb3Hf+AKif
7IkHZ/WbjdJFXQ99gYjk+Dwyn6zyZD9TaYBpyfhuViob/8joxw4oTCoCJbFEf+ys
XYQzeLzPrWJ69V3HUOmh31qNr7lv8F3vO7+chohHHAdICeucTCS76GZbGz1MYiYE
39kKfM9UFiPwxwj1xT7Ri3OfY/yW7iIad45j5j9XszG/wYhY+pvVKUsqcQjLfwUl
okkXw7baR06H5LrGsuxe8P7gGbaJZj48okxbNt6/Pi+564k3t/cQ3AUIv/LkLlmS
oWjm+hz4DfSZuGzRS2xonmeGkpbnYh0krJOiDWoTgzqjdWwRdQiweivzWOq3ooQ1
S7rRLDMurc92Q+JccbjIeDBL/F/9+7j0Iz+qycmagXSeuk2JjAZCV/MIU4LhOxuk
vCtIo3LhQLh27SnG5OaGnZGjD/oKGWD4kcef529Chb3EskO0wvTeH0vo9cVIngpY
ZcDftlz9Djupm29UzUPjwfjqi+KNNgbZr+Box2JtRgSJogdO38W3nL4UuOP/VSBz
RfChjyDdzIZFjG53jf5ugmcU+RWfmW6hYMuHI0Pp3ODCvROZd6QA9r6w/kBGaHRh
wtKb4VxW9YvI1RDCK9ewh5Avbzaod4gh107D1YkwxCzGcY5rMWCheyzQdPeTpPuc
wRsXHMUtAvi5qrcc2grO1bG2IkUp5aKS3Ro9/fDCbRtE0qJ9a/Iljgs/4EiVMX37
cgVsro+j16n5Cu0DpuyZAIkWAD4Yrw3NgVO2X89b+9zgfsqpB8fQw+SSIE2WO3Ch
Ho0xtT9ZEfQa18VoIObgUZyP3LqY4mCMmWgQG/nMs8YrBlm6E433+5Jk+As+j5jv
Mu9IN7gDczulOUnYMr5LDDCeE+pN14tBIlv1vzVnPSuN1sEZDMu9wZ0LQIcL9IvP
5s7ZyZF0SkmLwXR7PgxHYtgEgF9NFb/EriO/B2fcRcSzdf6dlDDJNOR5T+GVdZHN
d3r0nCMdqhel37Hhmuqr3l0sRvWj5Tfv7gYRtAW6kf25tEvrzgva5NhzgV/ymXgY
uwFhETh+Fgvn0GN9R1KktGoXVr4ahqE8Ic+N4nxvyDAazskRYg6/Fst2w7NODxb/
ZAjLbhW1kC12mbTCb5X6BVBkFdI4Y0kTtr+Ga16NmX/AKUyLZBL7Giu/6+KLH8H9
8T/aqHS8xGuV6ELGHz1Z0QYQ5qZCnwNCa+usyxMiEa7nBSAkfVvqIkSRfXjdN/o3
lEMbuxZxOWXk2g3V4TZUxjVZ8pW85/yCj1nqK+SWSUwtClE0N0GDSX/+28mDfNii
dvOhkoo45eCe2hyWR8LoBZpUgRfonGQWkWADqrKTC3NcOg/vQ7B/wID0ebfVt/qJ
DbEorzGe6SFJIs47ktyrTYyOOtzboPcMcfYNxUe+PhLqAIBjWDbOsGBhNx7b87MF
fU6xf4roDuF78pUZ9/L0zy0kAfRHcbG43CKC7RCFH+SrPu8TEMgUCyv2goTyOhUg
LkpXLFkTN8I1dW9mcuOrlD96tf3WX01ExVJzTPY6b4MxVx34tLm5oDUBGYlEamyx
dsNvnNlgfjW/AfPKpte8b6pPc2rZdUL5uo3zaC+8VueqkudXr5ElxVbIs9cMBn0Q
h0DyBtEaS1ye0FpZGlx4ffblU0uEzQWdG9bggUJd4qNnw4bom9bT2nRoPGje1bat
p42UeIy6ABe/+rEKRKy+O7ahZa93g8ok4LB1kOXkb8kNWpaMbS2lay+GUx/wSfoV
9S6mUP9TCqjeHZt4yeacutpsP0Uhq4aAxmWty083EDfwyIU/XU+rGLzA09ok/I+q
sAfagVlY9X2skkCxYM/jabQ0hKVJanRi6rmVujnkJxCj2yepe5faHfIDxMmzWinU
q9SqqfJA9Al82dB3ak1biP1uxd54QAcMlPIqylcBWiBeft7QkP8ZpH2DWWs1C+K4
yfaa2v/aE7Q51bjDp70ZBWvOXlZMCU6a0VvR75PagA0OuYpI3WvoQEUVbjLoXQUx
EjVVeczzHdf+9QqqSAFRFUGzOQ7HTdvKZ9Ra912QVzxivYzm/UyeeKn7/CMLqvAT
uKGHsNLYdlQeimClPPiLD3DlTBj1H55akze+4U9TVLJAHEl0YKYoPG13tGGci2k6
s6/WzBhdJbZYU02fzrmW57MPX4JGThNwQ8X6JA1eBTXP9xhaTEMsH+pX1t7IN9kp
cY9YAl5qvRwGz1IsGsjb41GtYSI7EtVNFU6JHUgaRgyySkQn+vMzJTyORA2NTC+F
YQGmBMBCZWKpxwBL8bW2Nais5XbOuEZi6zip5Yo2GYhAPXJw8o5qKtkAzGpaV2r2
lM8kyRcC81m2P7C0dJ7y/NXsQnh58LKpuT+2hu71YojMH3UbvP85pU891+zKOidu
csLEni0G1JOprgxlxuorvq77Ljs2LSWzhsy2qNyqWKFyaPGuw5U/uTAsOI89aolx
aQuwmfL5DF59brIK/GCCEoZ6u7y98Jpgjemvne2G4Zf3XEwT2DwRDULmECENyslK
7T/uGX13PUoJfYzFUOMyq8u6faD0h4w7flpJZsta+h7npF9xLrRmnUhlsUCnsfJQ
LViUlwgAzDYnwg8drjqgKt3/6l71CWZFcEgOM/g1WeLrQON3ac24GUX4mP3PJe1/
Hq33Rh2mPTjgZUDlCXkroWNsd72Sz5/DKX3vceQeCa+aOV+LGizGrmRqF9xaPVrK
89WfGkKaR4Fs2jIpGVY/nXv9hRepF5IOjnjVBypMSY8V+34nMzvTDtoT8tHZZbkV
L6BDsCigA4y2n4IxGdTmCZc4oPhXlRUu6j9ah7pBNXT6ktVmoxTpnJ0ZCc1ilA85
kEKpPHGRLWJ0TpXEN1SP4YepL8NZTMSAyJ630YSda9P+8Gzuf82nda0k9YAt9x2q
A3GZdSbBUHp8lTJTn4cKMfOIZh0iPUFOecUW4toNt9HVSeivQ0pbgSt9G98m/kQL
aiJWGr7jECl8N6OnvdYhganOMwUsCUHWDS0kt2fa6neEg2meF4s5No6OovXNikDz
oaKG1Ykeq0SxxmklTXEVCO0DzM2XqR8+eJp+rIq7AVVuEi3vI69K+hM8s2SuUsmF
0zSB8A30FQcfgNl5D/Sm6/FY5ORIIS8lx6jbjWMSsr7DmTMSdPlsFP/8IFdhCWLv
ZTk2uCdhkJDKxv1qOB6KLWDCMzUFtP91aoy7Ubq0WIDahD3TNQhnNPT/pPAjU6m+
111Y7q35yk/GWQO8lE/gDcM/9/kCQ2gxqF0to17UYZARPU5BAEXORsI2ObO7MNHs
0ntkk7+pirsjXfMv3Q8ZSuuvj+Hz8/Xp6INHvvABq0u/kJGSTnx1H3iAPea6twen
V3rlzPZBvrc+cVtfiiF30B8oRh78IkJCE+eYMQ+TY5rm1LKidQnv110Gg7U3FFx9
4UD4SHNWx+Txv+zP9oKKaSk/rBeh34ktyhqTVSxzN1OanKxOTHASum8yBYLlYWwc
xma6NYYeU4KAEBDgJtoz2JSnjoCaaj3M3RRu/l9jQYTppePK7LDnBuXdN8oBCfgz
5LwbWfzZw9w00kWmtVpng57qw5ba6LnJCO5qnnMvY29NF0NOqelUTRGZE8TLHRnY
/+kf0hwvgctNP4ss5tmad8DuV4xt+LXnjletZmYhi/NkGB84dHteoA92LAKvvy+q
CP+ehOsqCx6beGcpB/vZz3o5SaHRn/CUIsHY6W+eC4/B4/DDabKRcLeBaQQW3LDl
AcSW7K12u9DSwIXVKIuwypDRkhUrwcyTgMYDwpYR5KTOGV0JzzpxuRnCn0SsrJYZ
/4OJMZaoSS/zDqzI5LvXMXwXK0Ijp8KeCy/9eGqiChPFngUnTHeKqjUMBX5u66t1
Dn80bm7gP+uaDne/Bw5LkFWaNcbCHjT3o4Z53i3N3V92Er9k4Cmm7PywZNHGSlLh
7l4aMVec3n0vx/iM1PqmPfgVAvAaO86P/AvYr5kdPrjvco7YrLjLPGMRoyBZ0R6+
mlgC7TpcV1dHmfy4x0v0W3MKJ0K9TDLyvDyzT3kAAKmJhbL+kRK190MXg3FOPXiD
Y7xGP5W7PBIeV495t/sY1fceZ/qZbhtSPlvRrzMQNCEoe2jpgZHPh6gNfKlE3lrg
Qxt1WupzmUoaUVd8GXMQGkK2UdSAKleiNfiCE21Yl4+AXa9oofNdxaHHZIS0tyfI
lx1Jc4jCunCKK1UDwxxojqXKeKx1kNkkQk++GM4mfZe2WpjsY7QUEZ8AP9Lr4SPP
ahy2+0Ko4pIE8xAKos5M0xji4/VJ/XI4yPOk2JoWfAS+8SGn34oAZrIRnadI3sFO
GEIO8tej1bFWB9eJPi5twk1k/1pKSpMJt+0GHMwwPeO75sGKEcvWmZKsZ68dJpRj
UfY+C/U+Oskj8ECV3xIpcpec3Bvrew+wPu5+mdi9HYI7UOL/wQqI5Q9n1piy9hNE
aE2sbId2jk/GEOByNaX2XHrD1mhAN6mL1qG0Gpwau/xKX3AxiLwvSeDZAr9ohx07
K2afVN3+P0vMPJ2qpKPIhnzGIjN0lQWoSJs9RpcdJWKglyiY9CHoVduZhLLVdrg/
EpM6i+SNwGIJ13qY1oy3maU6VCm2wdU6BFm9tg3pwyMfKfzlXHDJgZ5CCgdubpub
ND2xWFQGzQ7FAFwh35knIF6dPiC+O7E3c/6IDHb+uW1sv5s52QwFR88+l+mJbU6H
hQ+LzU1SHHhq/3iEgJ00HX4llYEfeWUN0bokb2hDRVyHFCVLnclREssqTt3MGg5P
deWG8vDHbNq/MVTC0Kdp7XA7gaxPi4CH0rKy7z+5/pQr6mnndWLhNNHBTvA8dckf
pHLIHsNo3ouyn/Clb7tqfrvmNKtkv/fsyNU8+Oo5bGxE0azI15emKs6rKl6/NesT
4NphLJ6IuoqH2M3T76ZemSLLueTf9o6q8giMpKgAydgyJC2BIZWQhn0kOlX8RzDN
u+kn5mD3tur8k2Uagg88BtwqUnZ8r8ztCxGy2vXSV1Yjmnr7NZMAh2qo5N5amIjA
qGD7sOSJ/gPkjyxuEuOVT7RticGGdwgpoPrC5/tTZc8h6GvSqBeyG6cPKu/SGL3t
YlCDiKqlq25Te1Af1iLsDXbl7GdNIn6/FzcW9a5HVazN5P2b0/7zl8BaNRzu3DVM
LsjNgBqfWe5v6Yglu0IZdaCuG6NjRVqummj9bReCj/JHbZAwA4uOrSojoIRV+bE+
sn2yZoohBvVrnq5WWXOfGW8kE6ju4xtvlDpJtBF805rGVNI6IAcOFkRKfIF7Im8V
BT16cva5OlB9/AislCDSduMECfeYGU0LdVHSBWnWCkSHyPpN4zAFzFyBRYsSExRS
hxAqjhLyb7RGs9kfE12ZXu5XYOCymS7qQl4yqEzKajMRfU3hnX0j3x0nKD8OczxK
FaBUTS5xstvCcLk/nb55Dvm6gIesZay3Rbq1kVstjzIEeGvpmujgvu56hyhsWtRu
Nd3G80V7HW/VAZVdeOIupFw4acTpST71X/P/fCVrhout1DcMfzISVs1KDNYpf4w4
nFktmirJXYVNY3Iv7CARphuYdBObvXS5ueOwUfnWFcZfnDDGcLCc31yW9QZRhQmm
0lRYg9v1SVCJ2rMzz9VNnyDYaKfF7MkzSH58j4Imp9RVR3g35B6EqC/ZN8XHORTV
OU2+2XTcO3J0ZMpKZDLn3AnP+NBA39qyGt6y2OpM/1iuc8BZ8fMI5d2CK9qxN1bU
4as+voNr02uMZT6/u3sCBS+ujvtZB9TxPxUNjHNFI1QTjSlM9ODaZVl+5ZgsRrWi
Krhjf62zy1l1hgYRa1zPAHiebPx7UPRdosARzXYfEnIVIlE7xH3o1WYLYnaJxcl5
2Kv1i+szBGXQnCm4ePwg3rkpOPBVkWQ/fwf1k8iw2X7hVQ/l0aGiU10wXzMPTPTV
/pjsOsa7tFSHJmA2H/RVp8wITjDhb6yfibztS7qMtVLT/Gwo8jqWripw+YdWKEAp
cZZKuGi20y/4CCkKKGM/coq95E1tgqckSjhDnDp/FglCpMIrZw2yHqib/ebdtaeU
lieUIcX/07TZSq7YZFR2S790DXYbrgILttmwLYUN+IaEFLwL9uLNojYn7M7ydH8X
knOgJvBs9Km1PEvxG6dUvyD6amdmQLzDgHftHaqdj3qBzlazX0zW9V68/lEsGupF
3vjpZK+U1ElqO7P5k3XduDmqkqzMjZs//HCx6MQAv1ydCo9qMLXYT12PJPvgB+xX
eo9uiKSQqQZeqCBV/EIWohMHx35IsoqYG3e1fa03511cdl50vvJ9PBzpGYrbF71j
8m/R3iMxFCAtjptli7sj1v4JOh6EszxvE9Ui/dYtCQp25wArdM6zzzn/XoIzFh/d
x1oXvrAAYcau3ijq/eWTYVzkJ0o1vf8rMhGumeKvn4a3pH/3oa/BkRL2BK6aAH3U
j/kcezk0zxhnzPz8OGyw77tg3jnxlavDrXYJLKimkzTitrHbr0Ouyq+gscKDXpd1
kSThomo9kPl/qUqPKGWmVyaT8A2rALgSNcG5jkk6pUsVs1RVk5K5bLCJWtPrTWGO
Maj+0/dn6hPCG8UB2wWwO6ZiJEkFyE2nkKju5ESafh9/5YIXSqH0MC0ml6nQKASG
`pragma protect end_protected
