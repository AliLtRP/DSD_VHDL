// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FTfWeNPoTcNcHkVxC5zrvbaO/X25tlQrXdePs+Umiy4lkSzOAc2TEZHDvXSNuzw7
FQs6iuSdezJwKisgh0aCTeKjT0GWO73foQ0q+xwPIGjJ5xa7gQPj3l5QSjuCjgCv
JGZ5/ShyWNAhr2TArYyjrf1cGlKZJGUxXCKJU0iwl40=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8720)
6lJFh7XPpYmd2sg7fclZRmTVHLf8qkbxU5Z14e7cVJzY44eJdscnuby3laM46/fy
hTvtE4U1XyXbrgDlDQ9iAv/rCf9g6GYc1jImci/CxH+iMq8FTHuiWvBQk6AcEtv7
zVO9sdRYuMupn6Vhe/KKMGNxE2L93meY8oOzLpwwUb5I/mzBuV07zeFilSRwR3CA
IMSBMe5hF1LFusbcOyvYwCX3OD2vZvtLYFnBZsdkhjjf7WDLLYSk1B412s0nlVEu
uQz1gRYTAPA/xzzeYPNSKcCrvfjb8sILqTxjFymy3B/oid4GmnM+00s5OYEfvxBs
9qtssbcAYq44oTHHOOEYzPAfO+Uh8dSao5m8JldgLXeUBZXf/LV96aKdlRKZUFQ4
Gte5KfvO+SuGNUJuehIv+UUkS7s1EjDf/gucf2fjipUrAgOhCMNvwbu9sJE5/chH
CAcH7HeeMqr5TryxpshC+5LXqKGzJ0h/fC31dBeEMokPEuDcATIk3VYj6/oFbcrT
jGjaKgGNfMOQSwUJ2R8/HgMPjk6XGtTx8PJ7ZFP5GChlWBUzruvk8cFyNPBo3t93
RKgajKdMsxItcIyAVzljIXNQDTzru49LWg7ayLedJ3uUzCi7LeXcDluRu8oXMcVr
479Tu+Hkr6xcuokmMdm0h8Y7eS3Am2w4v4zJkmc3biB+trdW9i5A26pBQx1ZThby
3F7z9UhFo2ePqreAXhGazWhC9s3h2XU3iRLJReBzfO60xJCbd1QzGJPSt1IMx0R4
hdPL9WqyG3qBEyGuDhlu/w8wWuLyQ1JHenLW5+T+yfCb1ENEg8EwR2ZRlULZqjLy
oZBaY5eafTuy+VFdGhPq9PbY2u1Ja09/jrqGI5P6HdKB0MqdR4Ei9EYu94jZZQcS
/1IZSRWC8dCuRj5a7KIThzVyw3Pg/NNJMG3Al/ws7ySmyMaVBzetiHHXM4JSJK0B
wRPIWJ8AeFEhrFYWppFmAFVXv7QQVokqT90it/S0tDPEImiUaw6VqQlBaZzGTndf
kRN7r8E/f302aDkECe/tugANuVi22VzD0gvaXQjA/lK+vfw98OQo9Ycqe9vWuECi
3ZPP/LcVHDzjWs6VpthNkBvRhQTeE4qOcHQPdYqZU+VUUgKvW3p0DGk9pwj/1AO+
ZKsNaCmigi2Q43yT+6uqxm0MJTFRYFfn/i8BNGEthAZpJiIyXQ59inn3oiUm77A5
GVJwLOvAQPYqisZ4onFUhmJjmWqUXAZNSGlFJplSNuL3Gn3+vyrXbQPmH1jCYaJz
SiIRL0jNcyJGmXUw39aWqvg+6r/Oux4QNFK7T7J4xWOwz9z5UNUGvYNT2M2/XiDo
isDablQofW49uZ4L7/m8hph7+BzmlXC746K8Q8VbHfQ2ecXpwpSbF1RV9rY5AklS
HcrSfrtFrZ/nJv/iO3WavYWmTKdYOcwoPkeCHqyd/7i9CO+yRMkTDBPgGuHvAom/
GQWDs9Ds6zK5Qo3XRbeXUqkgs/yCQKL16/fG/xffOZg+bWmSgnm+fOHuxaPkILmx
vOuWkN22gqZ/YKxZYo158gfh0uEjSdmuYO/j0TWBnnmEBOCDhqDJ/HxTJ3EVIJoL
C4Cb8RKtpyI3E/tk2vYj+gQ8Rn9v+E0x7jeH7hNuyjJjY4pGniGamvLk03dJMpzr
J56rJhugDtLXDU6P3ke4xQ4BguJ+8J3f6mehqcpHCfiki4901r3v/UHQEWeCfJct
AdHHpWY6833QZW1ZoNKlbyV7wja+Prs/slt2NpPbymQwATLj3nVaLHbfnTFcBsze
l9QHUtVbfP0WKbZKQTDOxQCe9Ae4b30kXwpZwiuppAsy+mouUGzugPVJ7vrli5Ca
lsJG1tl2+WhXme8zh1pEWUB5UhhCN4uFURv8zbz+E7q2Nik+CT8bv4dyvnxkqxh9
KrQlUSw5jsc3/sn4WzGODRo4v7R4m/d5EerrQCFv17L6YljxQHLjrxBWjkukhoJi
Isey/m8Bv8RsqwZ6qUcT9d/3Euuj8dTAT1TXXedfDssqXuMDVrDo8vR8Mo4RNBa9
XbbxOm0dchvBX1gcO7STbH0N9t8R9QhDt1+R8Qci9PQWec3lpeSbGLHuXSYZR+rV
ktSp4dIrz9gneR2zvGcAgaBjx474tdkArBkIyV+jUnws46nCwjtLQKAyEp3gqHBD
jT0qVxzj8U3lNuZSN/b5xFBe+PITCtalBAWvI4GBWBuWqX8anVfLCWAKCOukLIJe
mLkdSuu8Ad0F7m1Fw64fD00+MadIGOyTzdzqS1cwdUGwJG0h3QjmOMolHWI9quxi
0w/94rWV6aVUTe/mlVkruubWnWCNYwUCzWp+OdnzjmyiHLL2GYGSjqrEUVdm8p+e
gpm2vlz8+432C5Drcz17rU6QdPUOSsCFNHhz9ttUck3LrBWNqr18ipLxzYod1pn6
ColN7Q9/643u8yugB4sGXHWeOpnXafckBZuxCEttVIP915QaDCB6uJFgogJhOrNL
zCnIad0RY4oez+jQVSKYtgzrwG+5YoZNE97nfhEmvfrS+UM8h2c7h/FMm0U2Fi+T
DXfjsj1paHTUfTQiRhyoeRxI+b4tTPk4kRErsPH1NPn3KFB+//+Sjo1yWph3vUSq
h/y8Bb0ZhhYbpwz94nsJG0S3K9wYBQHDRkjSF+DJ0Qg+5iJPPduNaC9E1Ueg0gg8
BPUN0Z/G36EwJnSNEbZQHfcyOyb2dLqz7m/l0tNe5wP/nfOGHAMLNeNzQv8gECVC
wNPpVcJK/GuQVM9ko0vm5lR5jS0k5lov57Z0cm4PH+kq5yxl7aOMjLcu1RRmv6cH
2UFK9eufM0HaBWXK8h2C3I2l3OXS5qcXrBjQQxL+kaKYXoECoXBobZj+9G8A+C/u
sg/s9xuL3iucf7uNC6CTMs/UMc2N2v70lZLXt3hyk+5gIo0UvKf5oYNu90lqdiuZ
3PeqcnbQNgb4tEfzxSmyA8sTkNgJlZmlWFcLEOcseMhQpkFXY2oaXYcrK4obh1zp
KQaWLAJ8AnHZlwyx9OGPViRrs36DoLmmT9lNlbfMAnvnkyoelOzXr4YodSBS60YU
mLd4VWLtT5QwOpb7uX/ABeHVNSgcv9A2vR5grBzJs4VUknkg2fJLm3Enp3+JMcTx
cnLaBDY+lfZqndYh2yQ9wk2ESQ8vogetBMtxIlpABCglOf6ffkN3LT9k0OFgkQ7b
psDHVlFGlJU2uptmoripaTr7Jxk3WdU0DD9/ECMH0IuC+2invXNHZBo7eCIEPxOY
xqSAHq2LMMlJNxiSPAB2mFxulwQGKPXh4SJvcGWjzoKrXYVP0KGahhEIdJZ63l3A
L/d6hDBF7oU8B0AOFYXLGLxakiEYaIpzf2Z4/WSZkEepYJDaEp9vIEFdBn8L/+bE
8jBxCd/dBWSt1119a+0oLM8XV6mb4ax3A7A1MS+5/unjqhkktibC1Hv0P2WHNBaw
5sWYwqKDgmL0f/4/gTq5g2VfjvRmV1Z7pNvwjFW0aIcG/uiKbzeJ//Eb5SsViSkx
AoY/XW1oAex8V5hjz3zy3j7Cs2RBO+NU9d3sKj4UZfmWVnaBl/586Lg7yaLBl+Xp
+4V4xqBD9DHa+cGGogaRZ0u6xGR9TQG7PgPPs0udNNSPlfH93sLn9CG+AR5u08c7
UXDDNFff1QogMdEWh8YLUlXrU1tucqryFVrNIgj2GRivFNPBWeFis9NmjEGMUljB
n/+ecaRSJdmaByP9x++wOJWH5xHS79K/e/DjKgPVwA3AzSXaAJCq1+KC0b3kqQEz
BA49sO6ZzIQCmFeaKlLdraBOVhE06noS3HAdrMzsGxt8hmamziX1Axg4CZVWUkiG
Y40FSmZdqwSXWl5FLqmRNwtoIaxtR2kY6nRlW0bmPAafPhSIBldvqUEubKzXCvl9
ypzikYuwe9v8S8qmu/Nw3NFmmrjP3xsWU7HgeMGhG32pnpiFBuUxxQcpuusC/3v4
HNHIFUhd0CKoAWcA1milN/NSaPbMBbGrQuheZ/1GJCpCVQqxynkfKF2sGGHKdANc
lAx/yTi7cAn9mDGgp4VLFDIFhtOtYS88BpEkB4SDPLrQ4HViDb8O9VuLitmnQ+g2
MOUpz30oCU8ESEWrpa7ftIKDRbRrBMtYz4+YZSdaZzt8eyfCEMNEj2CW24HTovQi
+isv2ncqaW6z6Dlb65tG+3l4102hG6YsHge0qke9UkhLbLgGbHGI9AVEEDo1L8I6
C3wwpw1XvdMxdyCQ0W2PGXgT+bo0cQ/PZRDZ0p4apqT8TkGPeZ4DxLOGGoiSRydM
pBYo6iAuXJ6+itvwaM5dG5HhXe0CfJmCon2yVyzai9HvUgiLytXD2CywWoXgbOkm
imLJgUYxVoS3hz+iPuiZPDyvcEZLh2tzfk+rRMVVXAT7c2DfqLBptI3mwy9/7+h5
ydCHJe8q451Ef9O2gxNnlSWyiBEJqo+nNusAwtKyglnGGR7F9oN6qpgmbf6OqXJK
VEjF+Et35Xg4AwAVI2ANeQ0eFL1WuPQYPQkX7bcD6SzGmnQBjIVF0pIIarBFSxox
mx7kXaUIHBBQ2FOsBZGzfFXelTvttBdu+ObLHvhIiP3OYXzdy6tWl0DSkKhzTzMU
3v2yubL2Xi4grnVazcW165kyITzmfhK0scubrb16czyDG1g+q/57AZ7wuXJO5DWr
oijD8cabc6oJP9iixCzzf9z6BqGzPRhFsLtqrCUtpG/T3wyQF43GlsOL94TFeLLz
hvA80Q4prOuChJfvyYkqzsPwdc4ZfQfZhhMezHu6q/swz9ER3Gy9FOuvmsB42WoT
OVTIjwZ357+gSzl31dNpdPxiIYa83rujH58puYVGXJZS+Cu5TaULGur6U55OetKX
WmaUB2v230vU3Mi8j3PYdZfh55hp1mNKKw1y9WFOna3h/PAwFL3HfCfEhoJVSRmJ
Slt6u7F7pMcbi/3O0LFSbREa/728kwtdE6aNIq01tKBV/CussdjTimXnE/lxyWPd
MVS6y2qE1vVp15R554Wcvlsvz5irEKNXnUZD4pWvaWEdQCthMnf/yP02TIxRGc3B
btWvVz5pT316cvZQxjitYAM60KTyJyYR0a+2NOB+o7tsEi1jQpH8CyBfCvU3fc0G
3tIeDxpSME4CfCLP7+nxk/ofw5oYpsykyjjryMzoro8PVHUl+Ew0SSY4oJ0P8y/o
Dj5KzkB5hKHq0kOIqrMWtGwffepRiaX6njvrevS9XVqzSYHvsdcPDh+3ZDOSS2H4
wAe0y3dpEREsgs+H9ZEAJpHC7Jbb26MwVJph8GWhaApJay1KL8d2Zh0v69QulXLD
a333w0f4EBjfXG46mR5e14uOu5UzEcHB9en+Hb8EK/L5gZQaO1O14GEnXJ/yH+Qp
XCCb8ab+4i24KYFL5eIFnYdCvIAaTBybD/9uQcToObB60bLsXlv3o5Zw4IlY4Hsd
qQxFC8n2zla5LQX04g3T17ADZgO01nN0SgsiNtjMxlIL4NI6RRWpo2qVdkANvlHO
Vdo6G6K3OLNwcLQt+TXYztfxb7i++YRLv0E8cnO54qbVtU/QJz8diFUkvFzndqa5
Gi5yjWtgoZJliH463P2BpgexuTjEhLbHQIq68KxiUHRUT1mhX7KEybaoini+89Ws
oy2StuoNop10fGbazCg2UATkQMpXxbEyGI+gbCa+rs0zHHGBrwd1DGrXR1cq6Dwz
opd3S7aZZkn9l8CA3dOLZ7cFIQ21iJpv6EkRy0/PVQSNm7NkmHbm9u72EP4lHXLZ
VIK6YD8ITSqI55nw+MKoybQoFcuEUvyCX3zxL8HeEF3IM0vnK3hz/AD0JARvje8W
a9uJ58rV9cpviLtPp2e5oQobqGkvlRO92kk90HHdks9+tSM2uEe4Q7UUkC/R0OQ2
wgl0E33GFrelRwh36ooEJ52od44NMwXiZbRiiWBl9aexnFIHE7JBibf3lw6JZI2k
KSPbzLEr1H6UfjQEgTOpdbVLabkRVJKR9K9E3s+hv0in14sol1T/38tzcv8G4EAV
PfhuBp4UqDYnLYX0dfCp63qXZvlB00LlP/FixPDoS4g8rgXgaGWSUIHdRj6rja1P
WWz2LETT7gMZoVg4YuIHwaMb2WiQMHm6JRTMsR7G1sk4G6794jenkP0/Sjh/kqX9
Xt/baGWQwf1lPiB/cF8DV7aSfZosbTL5Wg4dpoKV9hsiZqoKgNbGZ+t+eBginCE/
NJ0vz/IEBoW140OB/l3dArIdPApzoyNLOiNmB4EV22VZ+H6bwryeFZkb7CD5tdhE
rzl4iDElHXvd7P4jW+EZEm2rTkS0U+2RdR7wxlWWS4SprzRUGlVAgK4MvpNg25fY
97omxLlcJTPqz3h/NBs/ClsUBCueqtJk1T0Hv1UwO6sFwDFk3EIe/wCmvwSd+Hw/
MWZacMiFqJTRNijKxUIQWrYYJ+/0/xwopSb5mgco42hP4iHl3ydS2n7Ih/XHDUXA
wy2MUxijMpKr0N8WGqGlEx3PqavfTuY9pEaYIyBnaFyiVZra+YvM+KpbDqcYeAMV
6iJOGRMQmJ6/XVnZbwZI7Z+t/L+kKlRs9Na4YQt92kk1JM01cxNenKZw/LIR8qSS
rs1NzTZ7VpdkQycIPjMUVT/Y9G5OedTwE16Me+iKzq8P7Jn12hn5saET4Tb6vFPX
1qy1JxQQsn+/z3JsWGDcLWcWAGVZ/IekSNdnJBT/YXDQL1rIDIi8GIV1UBdHE1SR
f+NpnbHP0++bv5LUyHoHbErggHP93PbjK4uJaB7BE+b8mrKmIn964U1I0p9Ee3ky
b4oD1MzXf7VqVli9YbshqRV8EkkTWvyOAJLro0nTHm2swl6/uBtbTSAGeceAKZr8
EKcb99AiL1RALCYxBQBiukEWOwcliNtRox+FnahBCfMx5DyJvNV96T7dXjAWTo/Y
8Cze++mDq3yPToCBAQ90PxxqXpyq/boswX/+eMjJbcuwDa1TNrEMr0+U9g2HhhJw
vOlrZ0PWJLDUZs6mdTfKQG12bJhRNa2rN3Zx/Vf0Zsk0cxHIqXYkGpZyf1Lt3Qfg
95gvU6ieuFxpGO3+qAZjhtPinO158F6EY+xu5LOBNAD8uypnyYIJNB78gDJnJeop
OgcyPQ5Q2aNT/RFS/bZVYi2V7WJffQjrA6y/O59vGOMjXnl66TKMS12krjXwuTiS
sVjcnezc5gH7QX6/L4Z77/G/ten7FVLSmOAaPpgYf/M4Tp/9dnWvhLSIIUuUuR94
RZ7l2vlJjUVMLHVx1eYfX+ZtDM/UCGukCjbiNPQKks+/SgG3bbRw4njdqrxKj9O5
VesPTji2IqKE8ogTUxlBExBb4vF5mvmSM5ukxD9bz/1Le+WzvHm2uzZ6uZeAlJPA
du9n7o/EPPw4mRUtuGblzziAK+o1kumQC9/NpslwHMdOtgY2K9LP1yuxNqbf3g+/
nLlI1YVJgprqtgJSqepqYDeQZEWnY81v+H4qN504QWD8/pNVqBZ+UhH3agRflNs3
tczQ/VBq1dyvgcuXOrLOGEhICwXO8O9TP5sHK1f3TfU00jrKuEgO8yqCXDKwGtgD
AX8+74+gPPu6SyXxZTZ4BIgsC6BTAL7B7UVDNe9fMaZkMtweMYWyPmgrEYHMTc/O
QtU8aqW1THSN/e3BQoTNFy2bXlvx+/qQxE0t4LP6Xlp0Hi7kQyca42x9pgKoztq8
6PCoU2FOaaygmPAjWw8WhvxF9m2+9LOSsNwoHToKotNDFR2ITokuRNWKb7E+s5On
hXinzWhZiU3FfLxvs9M/SZxZRJeRysLlkPF+uMsN7xQ3Ap76RUJyjVlbuWrzoQbq
/9wToSbbqErsQl2wZa6O2qRbcW8VTkk8uXMJIxAdSI9pGBIMAcKOZUjGv3QlDy0y
xqm8UmV/77MqebVzT5wf+FbCXIJ0SXY7U2CWTBBVvJiiEMvXlgpZKgwZ9towLHea
j43zIzB9J877X069X5R8nox3ah31BEvGUT/6p5maC4jWEXF5HzJdDJnTEjhP76q1
vu0f0hD0FE7BMDMtZABvDBUjtv7bbI/s0jEsTNehGlTrRwEDEpr45Sw9A8hVMKiv
mW6cEjob/SxPoKaqvlGidqA2dDNzd7k+kFuPhmX2Sa606ZhrLqx+7/uo39VLjiRx
p8hlfrLgDLkrTS+QVm5CSM0LrRXPxxhUlgi3n8jlQOAZy852JeBaYPr9qL7agexP
/sEb70+Y5eBBMvG7JznDKIBwY8oLOQtDPYdUgDbxbrSxXtSq7U5LsKFAaZGjVaN3
fHvoz60TA77A5DxhdOKUN6qG4pOe+xe8EqUASnI4jdPNjKIN291muL41UBazUaMb
ZyAJdirpl4EmLYtuwcN6BPRgQKWENFR+A+cI9g2SbY2f5roD1p5fVPYMy1YRv6M9
NC6Ghc+fDyPESkiDS3csozjzWy4vQ7UsQKv9LaJ/ABxYKC7z4QxyiowMKY2Ts53G
QlYR0Xmx3RUoY4eOtZKPlFpPX0GQRNqcJ13tcV4dzNX1iCxG7ORySR005bViU7A+
JnVOo4cxg3N4WLNoZy1BdSExlJgVenWg9L15+2eh/mBEXbEngKl2Lazp77Ba2QpR
Ge4YxsSL+C1WRxEnBb4TC1xZ7KxUY7G62J6QtxF2gc62OrHYsxr3GvLxCVvmAtqq
gAifzPPwn7V1Ka0ou6hD2+vSKBqOpYikgpDsi3IzxRuc83LjklzZhfwxgCthbhq9
TQFqAZT90xxPjoiH28dZlp7/HNMfoWcDS1CKxQj0yvAxOk7TfCrXEeNCzWGpA10d
KX2qmKkV6IvYMymMomfFr2PlDHmqeGI+yqTARw29qKry4MCrXa6ljMd3cJzY6U+4
Qe7xLpRogNKOtv8zJwQruKTmvtAyrm5C/FimLOr00Nrb3K8fhvuY5m3DL2XltnT6
a0GdTqvHpMTeZAv2Qw7Z/6alTk6isAIAtTAv4xoeVXi3rWImLOH1/xq0XAUdpFpk
qvebBZHkjwBiSICFD2RmRQJ86t/0gNay0khKaEkDZPREt10EvVtMVwU0GRo0Ytgq
DUkg2F6z4aWLWRo1NL/fQqF4z3vfvRYDbWXrW08MBRPgEeG9gBL81Ilk/32qNyfL
hVqSyczNDIg6RUuh/a0XI277td/UblrMYT8mj7vfNn0N7+tbxPUoaAdpnfJW2liS
b/aMhqCUgkDuXUiinwm3QQ0W02mIWrbJpqZHOfqABwriz/mVsLR+i20eCZX/2aTQ
+CJzGnwD5fejWTPHnA/o4OeK+RqiEaaeAHzsHn5UHRrtS5Idl5Ly6RuLiFv42bIr
JDV/Q9hVJ1jm9VI0h4Wzhp+RQHj76DjgFBmw6uZCDN3TlUMDOby7VtUkLGItkQ+3
OxrN8KN+kcjBrwbOkOYKgIf+QAOhgCkrmLTFI0P56Egcn5utfvXH1TpEIxHcyPph
iMXCMoKKlB76eAHFzD8qnRBNor7VPtgVtIkGP6BQ1pxWk25mWKbusCdtG/QBlJDP
sYsIpiv4GV/Xjs6ijBAAVyZAkFeoPZXd2oSkEpX2OtwcoelrrgywbHR/me2K5yAf
AXtnV3UsMfCd6m847nk24UZcBXiKxW5QTWhkJ/hVZL7vnqUxpGmz4yXbNtQ29pXs
7I92mLfBGYoMEev5bzyvGO7yvxE5clAdchMD068jlLioE5wpRbVW6MSA7umRSYRD
NTbV/0ICYTLkaeZB4pryfbCkwaJKXw0ZCubERNc1qcb+WUIFvpZ+ucJi1tBDlLxV
z3E77RXzIImrg+AKAbmlGrpDnN78TnFT5n5CiiUxwAdSSqIkikPP1hQByeHkroRP
NGkprO4SUu8QP1dMsrJTFCSyRnIY+oHngPeObs5k1n7FoeCmpz7imq6bk2/9Ry3O
hogJn/Nw3SXhenpUmdxizGaqp6VCeb7huCMp9Pro117tdK61DVO4nSYRp2+kopcP
ZcjaORhMQoDW6IEO+iySxt19U/bobdNRzR3sIT9Cb9SNVRKBNYHmGz8nJXb93keQ
9X5qOqyKMXM1IESJ6JNjV9yH9+zMpCfXf7tIVVdfKL4dcJ7k2kep5pD/8BnIOPTs
mVwC3Wg1DyzqZen09317w+uCya1SwI4k8mtIOrKssLVuhNtkbTSrbhWCApwWm16+
iwTGV+7zyGa1mE5UdwzYQ2z/XuQ8RK21S0zJpr8v9vwqMVXrFNt/bYAsDCIuYjQm
9/WpcqD/dkZLug5O7ZhU9hR/90M3IAgjwmoxnmprMr93sEYSX37nhg8FVNxR3IWx
hIexmOt1nnF9DJckx0vFliabJdWv2/AjjGDQS8KpsvQ2MeKoswkKW3DsnKsgMVcL
hr6InZ0MCXuq2+4bwjJh84DPIHu4hXseHFnhyk55GsHab4tinOzK0Fak9g/RxQ05
R06/3PnM7GAloGKXkiiUuvLz6qza7/BOKx+QBl+Kw0bFDLW1Npch/HjrvDEOtsOE
R+f9nWS28beBK0Li2hRMkNWFD7Bl4iYcYDjoXfl0shm1Dtnd09B1jV/BrAn3WgmW
Z5pROY2ezcrNBW8l1cJ0+iG96t7pzB6XG9Ox+Lvkr42Tljyfg1hogHDAmxbHfg4u
HWavnilUBM6RidaXEFt+oXxi+CbkUFRAd79sVRH6d4osQTgkb/sJGG9sHF/KHI0a
kG/+8KTwuPmbZv/2gH4H0xTOurZlJzUuaaOp1C3GVjEYK5IXqCHWfqaXzNBRq2kS
3RBv/FYfPnfKo29Ik3yg4fhWce3KSie/fNgqtj7IKMZ7dizi/avS04jgfF92+Ygq
P2X3TDaTr0ZQpntsJ0gyYyZsg8rBLJzHy/fX28b2ohjobKmn6JbEVYMbMHntWAek
8dO77BwdPqDBHkDUFz3hJI2PL2b9/DEy5a0AW7sfraNrAWiPb0RM6yr8DNVI96iv
IQMc4wUb+5aimb9FeELPxRcXriNXtoeHPHRiJmWQau7CPaoJ7r1+EnWqF99To3ei
w3tRZ9EBOBp7OuFJTQQnGouns7Dkuz0GV42729yrHsEzgywDOECp8QLQyRONmixl
7X0k5/LUSts7vQWR63i6OFnR9GHUtSyMkJRTwoxzkOsffcUo3aiVYVlJTWM53EhV
aTjJuNI423UUUeNQPvi9IjLSYWXB92oYQq962XN/AEprfO6HXyuGKFGbtho8IJH9
WzpBOx/ww1gtkYkGl4ENA4flYwMEC2qn0pucAnDT8pmuQFElwED+IQq1piQws8QF
zDBLz/LPrktO6sPW0ofxpJ4pRJxvd9H5JZGuekcDz8g4k3RcnTxYUoaO2mJhrGT6
jtMLE9/uc2Tazv0BO7GJI8YLHXi9Kuh/aabzRppz64K29cYgjtxoHmob2tsDSYtC
qA0j1ADR4y2TjHJbgC7Wh3Q02HVnuqACC/NYqTrrxlaPDPm/Zgca8L8e+AsDM2SW
NkU4xQ5elsifnVZ8smmT9i7bi7h/GU4SzCJ7cXZ7ZuxKAT0wE7IY9CAzKZlyoG2f
8tXLKqWXEBrnHj69j1YlO8kofPl3HO6S1vMlumxcaEdfgmNPlRqeoJR+FUzDBWnJ
IThMpPGIFE7dG/nERzFTYD9K18qVd76o1utG162yZFmWopomxEuSrEB91MZSML+Y
jXuxiLynfvuYW6Iuz5hy+jXpwlBTl643nIau1Rx6HjA=
`pragma protect end_protected
