// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kvBWH1gcWYE7flQPAop2geNzufUzxXdRSoj/qExHhk0kKBT2IFnXsLvZr7vgELKg
qEIsWHHqvI48QyoYE5fZjE+SBxecOAM+AoZi3A3XZTklCGRek9InZ99P8y45e9lh
rmlT2i3a2rbQMPuD9bYUbQ5HUXrJN6Wc4V7m73NTlFA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
+CZOD6hDbQN91d9M5v69NSxjwXQSounqlozftpYMu/DrlVYoaK1YN8FQYK1Df5rJ
X2veQZXC6l8AvIFGY+L+h+C+P1QEAvsYpMFSw3UXeCG7MP0yOA7uVtl2RQs7WxOn
oFlU/+0o4WWTMmd9xtH2hNkjaoYcqKiFmLbnBUVaOQ+Ajaw4dz2ywjNsCIpLy72p
1n8tGLQ7RznmEJDIN8GanqjQZIa9bV5vom5sl2grYYNahIeyqNjVienni3kr9Nlq
NteqiChVv8M1gQcnuR6auUufYBqeu+SSeQKEjD3yZ2hPp0WPm2TTM4svT91iwvKh
RVIShtA9F09lpAKu4cXbzywHI1I4XBv+eBjQQk1lZ0We0acKUVM9EIadcsZ1QpdD
1rua6oWEk34Y60YAu4mtwxccUiL79hlesmhjn1qFLtCQy45Wo4uaQMUMe35iqTgU
+XOiWLhaDamSPyVTzCFFx1W5HAoVw3doJTamgTewNRmgyh66HQ7UQnZ+uerkzTwX
uoQROIdAv0GXUvlk+HOTyjci/7wDw9AspYqRKS8irYl14aqVN0ts1HvaMGU524CG
oMmEmS0MXSqzvhPnhnJJLLC/A5LV5DLVl0OsRwIUsqW5xXUHFrKSsEpigIkZfcL2
KRdnJsTqgZr7K3z/GrCn8Sc9tjqyaBlZHs2kjAV+lsHAfXo1FuAOUSjWUOB/AMJP
fV4eJAeYp/qRz3r6xR68uFT+KCccmZGyngFCIdAuBGzAZu4D8GbTD+EhZsQJKrLK
+UkRVRKiID/HfySEM7bx6vOMBirVN4ZDzKGdhaXWSBu3LJGv8ZjTG1hcjaIavN78
NqP1r5Q2qqBwQ9V1P5nPCh0xpQ8+y/tebUXig27+PsHvDThdYd1XnN8EUQrsi40n
2Vm8IhPhCsLSxnjad83nc1MJx6rvQ06mpcvqQzVkH3O5ej8rysNPP4ag5DGaA0fk
gSc8KywZPQ5+DqM/49sXLJWZCNkvLHH4FM0D/790FZGCcbRcAvATddL0ibJ2a+P1
IcdyMccgAgv61Wo+6Bi35lUOEqFcI656Fge/vioaIJxavFLZ/ON//PV8kp5edwsW
6wnzkuHlolutwI1XdQ6MU3Rm/Q5AOjOFgR0F5Z8h5nHTK+Xw9EJ4gfbjFpYE+j5A
pQJgncXGwjMJHjuNtTFhfYTdxBM+tbMhKv3GTeDtOQtUDO/3cJhD6VlKoH6sh75D
8SHC4lOh+VBAC/aseSyDSlXWG7deVpYVwP5PTC/v8v0Tt8fHAWwS2iEtwRS1vqTi
iASojN7QPXxQZKoOGF7wvvyGwh6q1pgg91NZaF1Y/0luc8yUJkTA2JJOU3/T5vtz
HRQb5JKbCCEKxw1meqLBsRe69HcERnIlARByqrFIcQz6gf48oEMswtisdjHe39Aw
T/T6NtWP6Q+qaQLrzmIo45gHcz+ch8a/RaJot+Jz1TW7+pXou+NaGqQ9DsT/PDae
1tzHUyrqXqh+HIKEeYAyz7oiduXUtQG1k11uk6d/mWtvDaWJhQ+MvK5pGEtCigwR
b413PofZw1ykopOVjrvVZjLEn30MTGr7FOeBwYjsWSdxNry0/fER+mXbN+qXBqE3
1TPrvKtHT8xZ1F3DlpCKjGlVbTHKz08riEAT2eCOIGvwaNfOtPViO7ewCK2IP0ze
f66sCUPLCoItoc2jsWUc6KItMxVCGlaKB4t/AAJNJkAsvwdnmae8/7LC04+XlZ54
tc8xsTZSPo/aMQ0AJiw56qfBUakoXI08xLb1nhW7D19kWEbfecr4+VDzD2RX8PNg
x0SM3Ohh7O4Ic9IPgYYkNWVAYQk75JKHD7x7Q4nQ61ROCv2TVCS3MS9p0mxdZaUA
7f2LwNhzJqMduzC/XbimEidBsHy713tnNr0j2GhvMxa7joeeiZ8q2htUgOGrGw+l
BjixBXejnQgp5DNO7Oycj6zG16wh5IpYbRzqbndeE1atxhLn5WeZA0kAr8bo4vKp
NJEKHx2/mIlM5mDNI/Lg2EuwwRUIjzpCBv9DCzDXsy2ZUOHojHSBsZD9f41czGwV
9RckWTYNkkkD6Pl3pQNK44ZXVRWalQJuRkf/n1hABeiS1YfJ5+dySQDhaMrFszM+
jDVmYWO6Vkc6fMqHrfjKIiLs6aviNvtyNdYBAJ79qntoyqH0fP8EihZGKCFtZGeZ
HhGZhVKi/eSB8iR+3WcYThWmn/8aebvc7AnFnaTvS46161qtvgdwlayVrfcXvGv2
DLXYh7k31/E5iIjHvlxa8TGQOhFBUt2SvGCj9SQPGLuQRszu4+Wm5fJmYTqJJn1A
ofjuSfxvS4cB3tJANaXIedq3Psh3+X2f97ZsQXvde/5N2nc6kaaKKp2rYiC3M+UZ
wDuIkpVjoIC/G8qh1G/0aXUhI4KA2coWT6HpO+P8+0WO03YK3vIaIrrGr6qmY6Ws
M0doqaLSO0sITODH96XpkYiEO3CynvdRXCPzGR1vK8Fu9RK5jok/fl4BpakorhN9
BTsTHvrboJBLULy8+peqNDyBqn6DE6T1OS8n5yEuYdatcL+lTLRE0wyDgWN116gW
50kAbWrpqug+zNItmjlyzq+pX2lJB8Z/bL8fsioXvFh5YCGW1LZqG02AvRV3HDzj
Tfzd4pTut4G1KLx1f/fx44/Q4RQnNDxrMgLSIYGA5SwSu/+am/gCRXHXq+xGi5BL
lPdqVTqVBXQSNeiDaAc48hiQjvoK/TI7lsdx4uMKKVjt2UtVEIX94SitGqGvnJfL
bm3HjYyDjUppNR5uKTLLs4crWxqPFole4AyZEQ896OylZi4QPpm4OnWnG7KjDA6G
ArRUNVwouSkMI9dY8F0bPc2SUqmt3/u562JBcyZhd3lEqlprZIKXwP186OWtXcDM
ifvvNMqa3X8n/CJP267cnypnYgTDjn3X9r9z9wO7bUi/PIL4vVNWpMTbdZKCwT7w
H7FYfcBikDyxnc6quc5qnkTNfhW4UNC+9sopRxwJjvzaEhyNzKFaZ0sL0MwPlSNS
oZaXuo5FHjFVft+Ai9SxyhEOSUD27Tw4a5bBRuCRwXoZMCm+xLdtdaN94kDYzoEj
cVegK++3d2SOip9oSLjGsv95sWgc4yQBrgGTmvYlckSBs56YKX6J4yOb0Vte7mmC
+YXcONf0mjb1fPHJcJOtLJ3lxJgf2wtq0jA8X0uQ6O7iIWaYG6K2S3W/9Ys55Rqb
bYIZIGI10HxQM/Gh7fYfhG+GynQAP7IsVuQkaUdjrwMrWzo/pc9bUsy6bYDluJP2
jkLADaeBCEfdeYO4JgZR+2qn0NfDt36Zw8nOFsScrquV6QWhvODei+r8zHQNYwKS
9zLNheiY8BEWB7vORa1QLk/Rcea2+m5xK/HwQyafryMAL1ldZ+ngsRxzYmWT5N9x
VWITsXAjYk0w7kmPnUzq3F5inY/ychOe/AxdKMoF4cQ3U0V48+Q++BQTe6+24RNS
7KkpR0z4OG0TXMJXyZpO6R9zwbE7aG06qbqeyTqygzbLlGXXqAsy0UKdGpExn3hV
KMv3u4MR1+o0jsHzuiQgudDXH/lTVVC/iZB6nS8jIWUs2Cc30bgprfrzMXwzuTqo
aCdh2IACKSr4gfJzK214JYkyoS94mmDQy6oDxWVsWjcR7mDTcj5hlbFoZiH1PrO1
MQqV2tm7/IXPV6UhcpOPRMFkkZ84qcqPtSjXEnz0zQYpk2WB8J38gFwEjsYdukUq
L0/HK6blLJ48xN1glOJvuPByqX97CiTaDNPe1OqFnC+HD3JSi/siV6v4wATkr0jt
oP0rPv8lMwarj+EbIaWevBFFa/g4mKl3eGl0lt7xpMxnBDw+5gIuZqzYmey3GFLz
XEn/N/1GWdjO7X44Y1o/h32iGjUM/CRgXp0RoPly5eoka20uuVbUeeSvafwvaXHR
IvifE3zbeQeU+Fmm02FMA8y+6MOfO1pKOOj8W3ZaMdGsPlEaym/Yfxe2s//sYFZc
p3lpvt4Bl9gsL45CFAitQZhlWln5hZEp/4j5C5NuAz0c9Qj7Al+s+b51GORrS+Zs
saA9UZ48ZwrJ8IPYg1GmEeq3yep+7SZiw0lWW0lERjiveZIeJ11thKlujucdtBnU
6c+WTYqVux+ram6cII7YZqVZlGmvkUJ4G88kYYgGmFmXyihgiOjWXbsiMYydvBY4
+yx7btRFWuNbycjbfrjqhsu4tP1ine9Zsw/LvhVd4GLbIZyvuDjnxaGyd7UUqiGz
CYApnCd3JE0rcdeHBqQ2wbS/gqnfdq/ZVFqseeL7BJNr/QJqkTf1SZY/RO0oTVny
6vpJWfIAhjaLyyLARIy8lagsBegHTsYHDIZLgmslaxKgcORJur9yR7ZYZeWrVvXQ
n/et/wdez2aBKlIgUubrkJtuZjh0Iugm7dFWc01C/jHoiMtDC3lUWuxxw9L/BslR
DMHDb7wnX0tfRQn+Qk9vtznGCnEY4p6MAVb44s0p4yOB9J2BcAFqQavmHugclGsv
WG/atx5ztj7C7n5mwPMe+asZoaRmjsUlhQZLX9Bl+Qq6b9FSmdxA/I+o38b1gnCd
U0d1bF9CUahW1JxzEhmAzVD3c/AIkwALzjcuYqJtBPAQD0T7Np+c3pnKZylHD7Sh
6baVNhZd9j/WNszy+jWOMR8XFVpBYxuqrf8/Ghw09qTI+SKa9FxAKE/TWagcTW9a
fyqXx0MqJZ2rU2bvkdbrznJuO3Q4T0H/hih7GhnkjSqMg3FCUZwoviz74VNO6afW
+gLdTwK4P3/vr4sANirCwHcsTQoPdc7Qh4Y4sx23aZKxTP1t8fIy0So+PuxDmZkF
b2sff2oQ5RFebKzp+d6HZSVOG2CRsZlQic47jsWyzHCt3kcfB/B/9zREYJnJecHm
3tlcvXou8STXZ0rXKyImtSnykPsdSsUS0PykmCjQwPGsr9q6dyucO0PQKL9rJQAj
lNf2NoVeWdEFEAK3HVpwJgbAeQxBfKH0mgnUH5ucmdwc7jhPw2c0G3QgVFWLoc3M
xva2qrK+xnqYCHyoKKtW96S5de+d4eG1Scs+x69y5FC1wgMOHIqyTnv0J1dOqxpe
dcEa5WifW7t990iEtmsJ0xPPdkfePdWi5NcnqdjN4XuVPx9bDrZdiO8jMN+t3Vqx
3iODMdMDafLhJOcTZF1e1yJbc5wTSEmpVioK5c9AuB/DqMwGA72MH6K+dV3+sr5J
+egulGjl3K0R5IcsircAkuyWVgiamwIOS6SfqRR1Gx48yaqOruiNl/3+Qle0AueN
rWzhnQe9TmT5oa8RXNu6Di5AghASMwyRInmdFqHMP2bvkD2J7dfKfDT1BB5xdEED
kVbeWsCUb30G+P7HODhY//GLjX/cjXsCwVn9DNnS5s8+xA75MlVRzcLjwwEQfEuk
NJFe47yUfx+zGnVsq72ruHZWhB36D6j9Nvli9w6/yzRcyjCBiukSjx5SM6Gd4itZ
JRb5TDOQo1bbYYUFBA8OYy3F3TATfb0CsiZmWzQSMYFNuwIwZ+5UEuCYibDuJ9pb
2MZa+2Nsr4H74c/yR1QN3S56kHhjMk+ebgDVVB8fmApDCdvHql0ohyhLbkeIaESa
SGLlT4e/eiJddN5Qb+JxQw8jZI2dj8Cr2JkRd//9Iwpgc2zL81U07gqjmeqRjrF4
D954x+G/cLk5eLpI6iE6YmB95/rsmh8jU3/Lu4xb7Pj5CHJQ2S6tKiFC3Z+XSjKx
1dMG3rHY3VK6BALw960JH5etZ8IIMiTjnGiOAyCygR7EVUH7vjZDQbkVfOQKq5RJ
nya+g8HxiLuLLoomz/fBC3y71tMsKhmPgSw3nh6FdzZpKfqRWESnoU/TMZPh/GD+
ojahHY6vNb+wzOSM2NaHlwyKpxNdUKm4RXGPaFTpweHdTqmgaKd3WutYQDURJ1jC
XIfxr3A21O+8v9ufZChLZPnOejK3Xkga+Rn9CmcNdBseIpNlESaIjmKhBsyEt683
4CB8YYrNbN3Z89ZCem9VpiilN9bSVd7Rh3jD6r40Ck7Xrn3zv7N4FPeUE0XRmktX
FUUJ3MsACJqyXah+1J0VirhG4XmivyHJZqbqYhSLCJamDrStCEGGX/WLk5nKwaD5
owH3ufgXNhjjZeQQfGl4DKPT529xrA+AJ0G5/O6Kto4GlbT4ygUnEB3j1lwuOzXl
a10p9UO7kmwV0K7kXNNWjQJG1eoLmeaWMmO2zKsqQOHvCS+wUMGmeLrxXK9KW06j
aFNJdRSEhhJ2zmwveZ/e43gex/MZ7J2T5XJvPupArBM/KAJRaBgsV0BUZtZPV2gE
pJQBsUFjnekCqKBzLrozEvt3eTBT6EcNmv1dUxx4ZwITkC8OS9/myxC2vLdKIhJb
IaYhCJsGs1T9oB1Jd+g5MykAIGZxGZj5hqY2lvbSjEyi3ijEKuHwdPtuS/lREyLV
2WZgdtVd2PvVJH51gAcmryEfpeICxyUn3K2BHpKJyRKVeLaLto4VQyGTLIwQbw09
zVwH+7XszCPv8RYbzvwg+GiR57lUPbOBOGn/567lri2L80Dc7rM3urgSTXzFBeKl
rUIXtbZHRQsP/9eRR8ZiOXOhXGZVYo8D1YF9ixCvg6PjCX/JY2kwG8ril/OIZ3Ir
y5x73GR2ZK6biCLntXRBHrec3xMilSKdZOk08t2/PJQIF75EBPcBnSlRIeuMuHTu
YhLA2t85YN4w1pHjOD7rQZlG10Eeigghw7+4gZ7niwQOykLu4GOuhKVk5iue+xQH
Zsh4nAa/8tmanksmZP0UU+5e9Lunkok6PGL+snjzc/k1nWtvP9L1jT2rxb+SJap/
TOFWzatKZtyaWattX3c0AIEAwDyNA3Rish83WvDSNXb23TrDY5ugmqSeGUZV9YfY
XD6kbGmfe0a7mJGjtsTpcOie0xZIYmUD6ZJB/ADmBZPpIHe80+jqG6f6W5oIyaiH
tYcd9x87Hhra5WFH5eVTyrie7wFIIcGXLFh/AkPPrqZf1ddlCWdcBfs5peY40KsC
jw3p3EcbuIcAN+y19z/qXiLsIiGD+MuymwLMBBciYpMcRkMhTE8AsQxoZzY7gpJf
xF/hASdmWX4251ocPt6xNmBIUqNHK+8l39le/TvyryIQf2SWTD3DCKQhZWGlgaPc
NSoc/6Vjgbcz2qNSkZliD2bl/V3FR7QmeCjBbLOFSoDcoZXjMJeZelmkyRMowpdX
bedtXQO74s8QXTjgz+Cwmg0ROo0WcMA74lqAlZvgTj4D0i6jkxy9lo5Eut9olQFS
Jtu/m86f8I7xNSD7VQ1kwzwg/8Fr+v6myomfJCw+fqY3g5BFpUxnbN8HJrOoVsql
LJPwcfX1vRMF20qFzQHdPluxJPY9LUWIclb2XsPNFG0snCCUQyecyJayVPE23f4G
llutnEW/eAhkSikR4odg2EIFGwqzX8j2mj1ugsoweTMvrOmqkPtOIjJVAM+++GAy
nBhfjnw4d5laHW+qy1WG+MxUTQN8cSk4BdimNXIze9PvDswG9HRqo7CzCCB9kIwM
p35rIHj6qpcIiewXTbd9LF6ZglUXQ09qCKECG+KwON6rv4gGyF8WqO7KB14mjcje
OD8xM/drLUkmZruWiRZKss82pWEYgDtiV+4ioBK4GTuWBZwgpFMakts0S7lLTDGU
yCoWr5McJN1CYClI8m7zSkQrLe88vhtE3QYhZfbU5OQqUvLjRJ5zCdIMoOwF0gwx
BDVoZzbFvZBBwpivn72VKmDDyuiI27J2B6N5asUxb60z1SXUH5n9V77NpXVZqdRf
3yKjRbg0t6M3DZVnlipULJQLb+lAHsyTp2H8eYn5W7awGZP5jA93XU/qTd7/q6L5
KNQGbd5oXNHWiSmcq+EZB81SvUvhGMALJLrEW2yrXSIoe+h/cDzIp1hoE2ztpoVI
3yTSeK6VRvfkrpkbfSS/2nIVYPJ5y3WAjVLMR/lVTBhdgxt8YuCks4/62PHk2Smx
EdfhR7b5Lrhozxils+IaZckO9S5ljqHoWCs4lPUu37r/l6GcxtjUTgxZSs8lzDKQ
Kx4a+A7+7WhPGHTWBPK7TIBU+tlep+VfMZnJDwhwpsrsQnkbBy6y8hQ8sInnZh9m
MFlOG8iX/w0OVsv5Bl3jMNq1QuE1TRgy6judw/8XnNoOdNaZJ9PylbQArli9rH68
OZp7TWcpL7lEe3N5F7wpvITHAOyaVwBOoN928lC5VZnvtl6D8u0ALEJa1ZlaJGJg
P01x3yaZSl9bKMLd2ZTryasIa9BQuC0YY7o8eqwpLAKH2/Bt3OnLFRIrflLbVgQT
20MAErcOg2ahVeuSRD3lfOouM1ZvHfhiYh2sfzjjrt1fawPOrqTNaZ6BYqbC+W4Z
nIY6KKMvq61aHh4dyMAFfVCjHhzzacQnEC2ijNOVlbdM29cz9WPNO9H9sBJ4LdIN
0XS/756Reenj8JfWbKvkeqlrta84+zd1ASdvvoOnVpZrqef3D6g8/FV9J0OBrwt2
m5s5CeawTuaM3Yd6E8Ap5/QgJv8Am2mODDVsKZ6Z5FhDABZiljY+wJCCMsnYqZfK
SWuE87LDznU7QvY86ywQnO7reueQqH33EmsQqL8e5QoIJBmLh3ogHpqT+PaURWdu
hZvg0oMedtU7o7Y9cJ2QIx++EZ4ygfguY/4fiZSwB90KOE6Gt9+hkzySIsK3lcqy
tb2HGpC4Aer6F2TQoO+7oMqoW1HhRWOjahV7MQi7N2Pmy0oLN0ZcdB2+NKmX2idX
CfmKGZDeoAdsAWJmHkTMsS/3/QQIO3xbEVaYxvhoH0NC+RgGLUz/ZKMYo8mCjTRV
7ERtkM7j6lTXcJlXTXZNp8eTvZBTt1JXz2eYgXZGTqnC6WlboP3tdlGP3ksEq5UC
aY7p1u+ZraqqqKTEUOD89i9OiXOUmN+dClDGGHtv7AdJswmnCCwHTmrUiKoujTTE
nXt4xtRF7fVGCoRSzRNuOifC0unyPYmyt2EobdCnxuGd5GXZE5eKtohop8bLowce
FC8SloVXyvc+o8P9kisgFdU6Buczl9lsPKmifSr0MOja+faWK2II4fmSRLyhBpes
4YJUNWcpjZU8rt5i1a06WDLhZlNoYGrDl+aPWOS8zTO4e61wLlYEX8pZqeIwXmMJ
IN6yZysgYZ1GBMcKEW+bgCarr+UYLuHGAKIxe+KfbavwvIwADpwGFEyMf6JxXIwe
Ss2WOVQKGR6P3I71xW8c2LK+5/wgNctOnOc9h2NFwdNkQvEPuRGcLLDnweMDXwU6
MXMDuNIYaXKRr7vSS7QDORb2tKlXHpiciWP8BAE+8Nrt7zNmG2f+G2x0n1HY/Cor
DEYnfUWcE+n094yJEzf/P9Pwb+9RvNSPfu9MiKbcVu6phZPWJA8NrgGJlWpwCufI
IKIWAj+1HyIrnq+wa1EwgU8VFFCFfliZWOlGFHhFRN7xQh1yDo7Ql4sRdcu2eYYP
oTKKUbfKJ26OCcz2EqT+Ib3ADHTVZpJAJgX1N0kVMwwFbbM4BK6U0MNwBJwSXz4r
amwE20wM+tWjSQbcJnSu2ER7GGKH/RZSnTx96In84U9VYjTPYa6RKaWcTU5uHXUC
fWCKlXBUeqFVGjALz9ihykA9lFfEgrHsSt0F1GTjAZ+1Lae2GoEtIbPVBjBSPH8W
mJMtKqkDBE0u1D1fnWcomrDPSASxHCC37r/3sgyAUo3KXPjENreAsWEQfCJlwq4l
XDZP9jatjzGKXhTTqAVZhWqOZsPgWEsaclL8a+sQwX+CU9K8T+7nANyz6k0LorVw
6l/KWhNFu4UFaZvsW7eOuOIA/Sff4naqkmkYXffPyWtR1vLtihv9NhJHIzC48C3v
AJZlAY1Tv5PjqAtHM/VOnzqLgOfZm5OXMMYIPnUF+2TljBNewZyawr+c2gUnePLd
POGMVKjA4TYykUd45A7T9E7l1fPBefiXUKx7oY7/GJAxC1KFMXqhEbLw0CHJpXxx
bHFFe6bXoR5dGLIgc8Y44lNGPK+1KoNxFTsNshVx4jmm4H2ZgjEmCyJVoAXigOVY
RnNWC++oPsRpld0KqL+nDFTz1CRZiJqPPZQkHAx8VkKv0l6NIc2v7IVXAu2imRXe
rz9zgBSZIvT5Yhttl2EbdwWUCr56gmacI5Ds5SgDq/o=
`pragma protect end_protected
