// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FWw/39ZYmMiU2QO0lkvYd5N8g077KLLsAP0ikBT6HeN1koFd9MKChKQdvO3QIlrO
1Sr2lWhb0FN6wdWjHOsvFBzpjOGnVYrVmRuT5q+yyBEkLCfouZ8RFSbHxSJtNxx1
5BNnL2U+RTThjFbeSfv2Ws7gzb1W4W+mR8eDhLIK7xA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14096)
Bk+TQEQNEE0QKpYRA0vIHRhcXIN4eGy0Mb+PMMkkt2G5MHSTKKODm7XDkT/amw8Z
oaiGqzk+3Dbu28QoCYJPPwaJnyb/IsXWMgQtQ09RD7jwfMVIUImtaPu67U3W32Gj
BqRZtR2u9bmY/LTDoxZJnuW7tsN9hRgVHEAg6eMrj35z7m+d8ckNHlRNP6fTqxh9
9XDGNEU9vSVyK0iohhnD6NQSmovchFjycwBTlbUCrT2lMT2e1GEj3Hb/7NHz76ZJ
YGK1zuw3bCfN6oGBjEvLHWLsXCkmmAhMFvc9D4ena4mf3aHbmekNyDKtF2Cs8dSH
RjBoga2HYl99DA+3pNK2o9kzetLfW04sdGopwTVrLf6Sjb4Tt5+ywwZTQvSCM4gR
wOy4zgDhXJ9znd6EMM3EeUwdBP1DXo2xRmYKgW34mXPSzp9xAIiWANBlyP6Cpa2G
nquhdB9bi2xy0d2DVADrQhMoPCA0DT8fMaJxyWx6Mz8B70H6KffcSGae6Ddnf0Te
Ccsp/lljPTOBuhc0v1BuxRpDsdDuPlnYRwjfUaiW7foiAghf83r8PxVio57X471e
LZd0/VWssgXcM9r62nkv5chWYPSTXMnC3UOi7ZXJhEu3vGkNAnzffbEDek1WjaWr
c/FsPfID8n7OMF3Bpd2qzjz4+RDknuW0YBrthZP2I4Eyuiorp20+EpTLAYskM8Sf
gQWdrAx0g0q15KORtIhGgh1EJxSfL3+f/ko6LP/YNwpzfEE0W7SCIJ/2bHk15KCp
xcmJ3ZxztPRVmgHx527hhCvLupBmiD2g7Rsui81t1Wlp1DUhMeH3ZQ2oZnZCcLYm
c7ZW4aLVS61J035YjW+dos72iKLWmdBFm6zXvu5sY2TsALDMLxQNy30FM2FK9iv7
He62QufXMJ4OmWUZE4QktZLpcDbF6kSnFfGIKMpohT6IFnAnjegLf9i0/il11jQK
lbX8agHMJYJnCkZukG+YUUudJJNN+kWoaq3aDET19Ng38T8Li6MkCdV7kEcmuXFf
gC33gPgScCAZiBgSEiTovePh2fkwZb3VJg3eksJmNX5YsAebVIqsOfAg5WxADmeq
g0X+5JMdShmkQfYMGCaptDgZ+cSgQe5Gxa2/9ZFNQM8O89cOa2TuEA++0bWxKcZi
tRkZKic5m1pJ8jcHGZnQwkHsqjOOVqWvRmEkKVm0bmWL8eNkMa44D7ZJp4O0nRG+
yMiX9OnZN0oLTzjUXK/CQktTOlBLdxvEd+32nF40/6Ppbda33/MpUlBQGArKz01R
FX3Gh3Ra26UZ2ChxyYaG9loXCkjGAMeaKwWeyMmdCzbKGT4QxoNdbK/9D6q0zWyf
SKTyaF3qEvu2jbY4x9p8YXWgFVTIhnY9QLVDdTxYIt3fzaAKqn7TTErDQhGuLn+p
ImvL8SutRwcR2g3U9H8cNey3o+SJTC20FI8PCB6BZOfhBrYKfr9swuoRXB9CoPzj
Q329j0kFuvEIXY8aPL04iEZb7kk5GHZTBkzEGn14H4GGjNkso589BftejTVj1jkk
fqQh2q0M+NJnMEVZWUhciytUxwY1L24vCvOth9Pbr/DPLp9ZiJMkSR+8/Dts7RJb
nxLdZoOlC9B0n3zC3zJcTe0k2y3BzVvwJllf8ZlPRy6R55IjlxxbhgQwDxVcxPmM
evFjiB7o6KU/baq9DL2w5jcOMCHJB2XjhzNnwq5kd1KPOAvHLgJ1nGiIBNFndeDK
GNEcU/q9wAEc3zER2sgeZNWDr3dXAcxHiVdJEla8AK5WJIT8xgX0Ze1YlD4eTJqT
Cedmr5oxeXIjGHPzi1SYZb3681P9ZC6VWuIAnhJJpSZU0zd2vcAAq/37HrfAk30j
VhCNKUSKYno+ZHw+OaGc0lEwhhG3k4ulnXkgHIyQEZp0i8a5gIoIISxMLenbhpr9
HJt7T21t/7dBr0dy0h7QojSuD1fIvDn5bguSzo1taqWcQl0GADtVgAd37KSmOOBl
rsyuuxk1fptOVZYXFeveVQ5lbSDxdLn+a0vZE+eP3cjqjqadfQi/V4VlK+wcYdML
hx+Jl/8o2qY78uPXR5nJei3F62BER98zMThVlTB7ozEB6Qqsv9IQLutd6dz+e5YA
QZHmrsl/TwjX9rLniYo0b1WCDf4gxO6P5VjXki+6tjLqmgDk0kL6SUkT5Xj3Rqyn
Yur5RJ5pPgjJ+GjorwgDwNywbEE9H/Gfd1mL9+wWGBaQekmFOxCeGFIHzSqGP4v2
RzK2bGyGnMT9pcOTrcPQZ8CyLZbAyAe8JS5ZwLQLphoyyfOaLFxIy+02LnOmtFi+
HmTIYbJ1PAxOvskiFQeRqVLPZclFj4qldzA/Q64TUuZUKsdK5B4x0m1De7Vfsih5
o/Lirsj6ph9k4QEB/T32yRFYEloPBpfD43A88w6046DvQcNn2mWBP4Jl8sDWZplf
e0rm+NLN6Tw56cVjXGiqc9jXaYvyCDGDuwh9EfFjATRZC2lGVTMGC/J7RZ7ZFG3m
eX9aXakJ4EPaf3O15iaPil9tlwi5Et6PKytZTsBHuj7Wv2WRn8Uh4pVR1Y7mrL6V
xHUwkk69wNLdK0HG5nVWPO1xM2v3PA7EoIrHX3SLs3QSEjyPz9h6lVf9BUyEUJdr
hgP+YovGc4WjES3+Wxsqre/Jar/LnRuVGDsYSPe6FYlMWnW96A5jk/kkmzHSKQz6
Kze05xaZa1DUCzAQaQ9+vbPhd0QWfYRg4+uurRVB4aYoSMmzXKRtdf4r9hdHNbn/
qOrEBX4uBSRz3u/VTKSD6SMAn6AnhIY6g5BL4z44d7cbpptTnbVXHF4g9RUyWLXx
bon0OQZhFXCcHOYugm+vjOinDQYuL9n5WCQMDD3rw86ldnMnUoJWNBzObmrgWZD2
kFVGkUndzeJHZzAPssqxfD60RJNK6WreeSsMUIwJU85DhTTaTgoZwsQs+RvmZ0GJ
Q1FcNHZmd5605Rmgc7IFY5ImCr8WmYo+XHnQySS7TtonKEvFz/I3CLoeAJdRnbW4
D87vhs9hGCaxPsnVF/1gUC1oH1CESj3cUQPYt3vCuDkcMSwJoiRT9KyuD9u2Yz8V
JlKX3yIYIp0NSheAtEHN31/9OyFUDYM9fFbdfMyLlOa7FwDObqsXL0JXcvpBrjJG
7GiNZCtB/duJBsOyGyDtOmlHj6w7iYOH8kzBs8Ip/euhusdnb8ZHtvPTleIJQmpf
EKMxo19TTj1UJ+3P66woh8lpfnqBLxCX3OyprR44A1qMgI8WuaEjycZyfEZl4qbx
RKcFER1gYQ9kyZfJ6iRp8Uzfwa4fqq8p0E+koaeCL4GsErhLwk8+/lF3ro41iS2/
UB9m6YY7fwHeuqr0lXMNYVP5Rt1cnBOcwijuj9A9Ybi1QS5s8xL+2xdoFLXnX6gW
qMEajLAgWJNKiMHhib0nfZonC9DcR+yQDYZRTviI3gAOTt6jPb+zuxE4yDWMkdm0
uDnRXh/luTU5MdKBP0PADBd9saVvznYOqI1JyetfsYTr5q9hM+BTSCqaeJtArWDr
8cJuv/GqYcREwbv6bIP2ViM33+lHs06Z0K2EH62VWm9LUo+82bdXOb9SzRPjyhhg
DlNSjbaauzT10f3Mx3OpRHR4Im3bVCMDmRC4SAI1FX8xaF0KH1wnpz/dfFn1Omuj
V4LHbF81iHqiOsxjKh970ym/7HxickTteAWeVn9dOX3LMfXcyvS00EuXbtZyw2Gd
eyGo4SKRogOOwGvPiqIwzL0JDEo37RF5cxbDfOu5Rv/q0/4reOidtUR2Wfmc2RUw
mDww5OuV+HeQGjb9p19CsAdx9KnBXkNqTOWf45K5iRdrti4Xc3vabQ2c3b2KBql8
+odX4HY9smezhYAd1OPq2T793mj1t+mPflOxSMrtzxQ+/CNGO+M9FrfWV1PfYeiK
j2IzfNGbslUT/ieWlhlsn7VMEinGjtU5Nll1J6sD4ESrxNfKMzIwybKtmtdPdN20
u8OfCrjEf93OD6gtHSQvwQ8YNtjtDGxato3mw1sftHxAD8RybzIYpD/W+f/TAzoY
BxNUCfxX0fyWxii6S82775JeW5Bj/Vo/GS4oTJzvpTmnIjGy4lWP/ynR8zgLwZkW
cikVDeu2gFor2TMP39LLJt89XCnDHHyD5l1JnyYlDm1tH98h6JxRfE5zkXjaOCe8
nUaiaFfVpuS13oXRwIKX0LUhnjt4xpoJ3ftxSDxognLJZL1G60Pk/cBao3JF9HiS
wyx476Uh6wq47VmWL+QofoXkpHpKLxS0047j4kZa9EPJEAhysJPDVRjxYvZlmfFL
nqxYuRcDRWSzqitF/F2bAruXwEtAloVODIlYYuzXiyabiIQLvLoPfaDZa7v890Sb
fo9jELS0AKRyhmbxPOepiRZfQjzW8+mIWKHM/ErswwNjCWit75+JVebggPkC6RWY
Gb/b7tsgZU6WWbrlw3WSq9GyHvBKkbZEnyw+Jid/cWtGY5bwua94DXngnwrrPZTt
uO/4zPmMyHPBGehbgmNfP1LY9e5bDZZqdszcJru1DnqlyhV/wjpTZMu8CDYH41wS
+WvLxDw7slu0eEBOqUNdfjMtwrcKwm8soXhfpuotcntICu99/3aq7vYNIRjR2bAc
T9RSHs+RxyfJXpU/gxpwLFaQygzI79octTGufPFLRjPfwzqR6vFT6viZ2J7Ck4Dl
SFdy+6qhLYYgg7x79/ULbNdzrtkZ2lfn8WHNzJKX+RqHPa3htqTSL/mF/zedsw8p
35CXl/RVndWcPLNNT4AYv8fHnSGAotgLd1GYudvk31FPfwgurvO8f3/n50YXGvIN
rY0HZxCPWFUIq78yvEF3YKZOKGf5BcyZvTmty/+P7K5mLhcw2dmg/iRWsOKyZJiR
gY0FQBu+SoGtbOZob1I9NAFwDMErajYfRjcSy+mUBxQIUYxFayiYi3/6RrtZR/D6
OOyh39QZOpyuUTryLhV9s17ZeVdgH6lpG8G12ryGr8GFDOE+awDuaVBO7fzCk34O
nQtVrCTMMUYLG73JfBzzg86s95n6FbCgR0lx+0PdP/kCOHjnHzYq7okZ5GH+G0HX
PZ7mxKGCG1VWazurNNyIFlpiTeKGYkgTT/VnDM+rbBWMjc0btmQXYBF31mC0YPk/
edYi6+9yTQQuIDSdQZ/t2+tHqt3dzA2Op7wdA/oJfSDhZFDTpKfI+zC+y38zTqRg
mQ52ZhKQ0NPvplnhOyjnTOVJYtLRERARdUQqSKVUSGk3RiYecUPyj8CwSzC0Q6Vq
19jn+7HUmWX8b/XrVX9M3qw65Zu0zj6eVN51FdRi50gaYFidCRrNRAS1H16816rW
VjhwPT1CtpsR5X5TrBurL5YXzScX45tr22RcU0ifV05XcJu5ikdvz1wIaKgS1zhw
7spr6z5GAsn671025pzHAH7rCFSjdcw3PwHbeIMxZrzJ2paqECQRmvH1QsU6n5fO
nZibiumBfg2jOqsU16viKd0eRq0Wq91rq7MChZG6TcyH1NHlRpCRVDZHe1mrem5C
7g9OqhTMz7VriWiOdGxAoQRclpnByAXaDWiQeCCDDdC7+OfmGc4iO1iMhznEt12Y
AugfD2Rs+bVoNvzQSjxYr/3huwYvaI0jZZaVxehmjjV190P3m65ovN//J+tjfdJ0
TZctV4lLhPQGtGOLgToT6601aO4kIqYYguWDA1iasNxfHVhsM5O64IVX+UeR/mlE
q36ifoezLtzGPRSOR63VpkJJRIGdRRvtN3yUHb3cGN7H9xCbBUAW2wVGwDdO49QF
kcXd+pT8XcZsOB3O5edEQD9Q0n5IpUeSHBpm9LbdvH9HWVnVVZYDfWktUMgL1m7k
IFHUJR6TqLnCLYiTZUyHJdrSJ3TJaWpsDGaqrZO7onB4w/fnq1UP/RAN5eC4VB4c
7ti/XIlnjx4aIQBPVAf65dr/lRq4C2QfvHiK++UMH0R0EcsEgvhtAKdXnoWoWg97
WcJEdfzEHWNLkyxN0Y5hWbW4pbI2DgNTvDAbdZep88AVHOsNbmpPSjWoP/I496LX
TGRW3aIm1Ihm0PhloKYIgAMmaKd7/MxgIBRVI+2rQ1GXHWn+EdofSrm8eJD3t3DP
2njjky0bVBGlyuDVemVVtMiLcbuC+DFsR3BDSfpeU5ICc129UiquCu793wVkhQJL
e7x6JEjulBpZulDIP6nRRLi6Fob/81EoMcVBNgxbPiiw5Zg0Lh9Ia3teTGC+5s6M
xCezakLKmYmCuLqTpqwQmGYY1aw7xqPqqxxvWnfzpvpZKodOEBVVEY9HO8RyjfPV
/KxUmPa79i6Qo0YBhts2rZOXd7y2qFehhFYPPtGabP+Z1gAB3kAQMQPwQe9bHQzu
v4GqR5twnr2yHBQo8reR5lM8VJIAE7Vn7LmNJphmQwIr8sXVSAxGMnXiFx4qeYIi
1zdLVEy2+5wv8/sW3k0nnELouY0Kv4lmH4iSEl0sq8i/7i9UU6LQRWQRSzc1GmMX
jpPDt850MWCYt9fXYvZsMQ4ZK8BZLCD6316Q/3/PsgNOpFwEY+Zf5u9LCWUBLbdc
HbjowhZP8W2FHwT5DsNPKVjfSDhc+4T8EJ1FgwSaK0lUUUjLNWpXBwyefYu3q32+
GEeAfCQei5/fdhbkcYF/x13DiLlN4HiH7ZHqyR5lynn/V8472ls5jJGtyn3iMcPe
MMQjQc4NIM4yKv0P+TMYeHqa8gzuq5rQybfUpbWCPWu1HWK4N4J/xP3ZOiVd4kgC
gwr9g9jiAW2HtsxUzI73ARfbrGlNuTTNZQlU6ikj9Xn+Qy8CqFWgg+sAyaSX91LQ
wQFOl7kIL8LBhQM1XebU14mSQkatAlhvH760M/HMV72YC3WAvlsCsXb2m75PISPf
8JnMeBK6tuRgMX0l+qXkRBNLu/xheARcf0h/kKMND8TY3+jpSRUqb6/3tm9lJthG
k2eWK9QLThds8HzPvZPxwk4NMP19mX1dODDkTKz0ufwb33cxrxkLDcO5rONvAX/4
8NL+jv/g/o/YWgWMKMVSa9HFCLv513OHz356R4+pb41B6CHCt8ivffOmiAilKWmT
PdqpLC66WHtTF31RKzSys9V0gTSmCeszWs5aLWfHbITiNQDs9+0zr8/ZXxAQ5t4J
TRHSPPla/M5090uPcgt1JJeovqnjwxYI8gRrvlXfV080/kuG68shkjdDKMkpqJWh
c995wmg5/0bWukIJ2c3HFQ8f33PdNFodExnGO7DQUmcivuZa2gfuQLCADmDJNimQ
BZJFw5/gs2Wx0I9DpRDCSzo8HGVJv8FWRXx7CKPNI1CGZn7RhDoqV29zrncrIWnG
LZFETipByfSCsqaRayvj6I2GtBeMbwf7YHmsqZXX1+hTlt2YYL2sTpEYfgvrGIRH
MJmcstaMhNmVvuEze7xo6EUWkfXRMGPzvb01BWyEoU8Z/X0JCh8vQJLEndwR995h
C8XBDXYUzpW3jV65FJzQCDOlS5G76UdOYu9TmHmGVlExnEJuN0TJ9PNCCnL6pL1B
IGANAfC1u51vLc7J0KM4D/9s2wDlireBTeDOyP2o55y/EC/9pUEZ3GoLt2q2/Djr
mBP28oCnhYJr3Jt9m6zssMVPviL17pKKaZrZW+uxzEVwVQwgvfAdu0Od7BeOl4xh
6KG8TIMy+7VDHQmdozWEScf1h7+W8JEmsSdO5KK0ZtxwNiHIF82O+ljJjdOO0WpT
nphlAWlOIJVyk3ws2DhBoQfGG+XbIV/scq4Ij0cXPDI8HdmKQ8lbW25nYRlaPg9M
cnNaQrf7kyBl9KR5dN1TWsb5EQSUNga3LSSb8YvhatNmF7vwjiJx9UmiHhrFK6vU
4cqO0U90SrGQvjuEb0PVUEcvCwA5J9vMz1avJA5cgLVv5ScCZz1eM3pGEE3VXj9i
uO8JSs6iC+qvxYw/lpArqMGb43os2QqW/uKS07TM4Ta9PZ4js1mRqGLUc3NVvcEk
rjWHlhejIClwCSHsxbEjR+RyHR0kArHPTsZctvDynaSzTxZIU14BYfjSLgHSpEzX
C0JYqvIqYOlfcgntgS576ezs4L/8LrFEI//EpDp72pkmIoIdqhFVh+ViJIXAZE0r
1iixsjSGSTw9V9ML5tkb4vouRXWlxjU4sYHcK/JmgKupXKC+yeUFbiILge3lRfMb
MzE+eAgbba2iWxkqwbKrJl33pbyosSMIxZyyHupdhwaxwY4KXGcdPceQxYMSCAr5
RI5Tg0RlmSZ1CSsnSAOhlTOgiomgEPbCiUoRxH/jCAxQEQw/qvuiTD/jwxT4RR1D
BfKKzsXID+By+s6eT6enOIcPC20EYsPNiD5aJbK3VkVVKqH43p9YUuI17yqUlN5G
to48YLd8QWvJMzh862BYMu5giRDYVRryP/l3vIp5gUQM9nWVjWEoDtUVzERtXDna
L8ZVXDvFGa7cI8QwoqGD9jfdvfE5WjUitI8zDGtf+snTkarN0zrBo29u7oKOtyj+
m1ZMvgFBA3axbFElR/uGOCzRoylTqCyUbWmBoNh60OA1zMVu14V+Gu42cjspFZEW
q+TDv2d3/088n0zlHc6d0oRec7mBUmUzXJ7fUvyS2gHv81dfjBGFiu6KE/RWKzoD
FsJX57pyCfKcAQHVzcFV0Ap2D31EZ1QfuATD20fNLFj4Q8vhQTWrdVazKdn2Xlds
t0GcypSznJNK0kad4Mym+pfmdr4xLg2pT8VmgQwNctPZS4o5dfyvubAzq9DZjTeB
9XNJIu+tXVocJs40fsHHvhCCBN1rzXlHJR45xnOLsikwrY79gN9/8rdZo2JcAkj2
mNluw2pnN0fKgb0Vkgyrwewadz06+6SyYZCcCcRav6ok2UIvUrO8qUI0kxRSAUn8
lPlZTYWy2NkEv2oBElLJ+As2FewaSTbwpb2nB0RhktyvBO70jiCoMtEJJDNWRUg4
+B8L7Nd2hfydegqeiGuTtCG0d7Re10wlAs9kYqRWNs1iRddxnX+J4OPEno39QBf/
SXkmUvwsqZZfQW1nST3eeoX4R+evVYxMlZJUQJkYGvg3YMkHcn6VQHKVn8MX9trG
GDK5W1ibb71Edp35n7gU5BI/W0z/JIxt4fPGgo8N0+TOSbI8y52bo5s5taxrB7Pj
L0+p45dwuhJj8vpyC7+Yk4CdpDDOhjfYu6XNSBHU6PYmR/RHvtH2k527p/Wdxh1a
HtnMU2r1aM7+Gx0oSfgcmY/zl22/wF/LrcphA0TeUwKLS2QN75Ak9LzsaReoUcIj
MBBj3nklZIaIGM8G5GrDTZ9BBus1KjQ8KzpX9eM5LGQVE9+c1NQ0Gs76wQcfRLZ/
MLQ7A7tbL5HOTIEqw8A2vGgRX97K7zFPODr4yOvAXFAMFxwZtzl8WuofYDg6FOJ0
m/KJ5cdQyH7kQg1ulDrcxSAfiymAJGjGSdXAV/2jhWs3VaQAc8uBHc3ex5X5LbpG
RjvK7FH8dn1wF8aEBzDkS0ZW2UNN9F6xb9yFyLbK2/flVObp7f+Byu8TNsKxl7QS
Cf/JbUADTa/Toi0spmgZryBa11OG634oMdiKWpHGVOd3ejBX8lSu46kxjGSZDaue
jYhdkBp+BSYHoug90aYK8xjOePys2quRv1Yl71E8bEDe82aAFf1YvLqM1H9+Yq+s
7n+vu2+aTELf9AhNuxIA/0siDY3q0Ii2diKBJI/5psHQ2SHmQzKMj0PPa76ff3fl
7Nxw/qBI+q/6os/Q9NHE+Ku+hO5Ua/tG7kDvFx1W7WUkiqYWT1bzjSwW4F982swR
las1VKthCUytX/hJM2G0VPzGM1JGXNxevYhwAj+OCeiReZKyTg+5IOdDBaQk4Vxd
pAsZYddxXQkh9kctbcbtiwxXw3FBxXO0n/sgtojp83B8dw2pcerWCEv++q/jNgIc
R4sphgBOiQgjCqwdADznLKflDv7pACXfCqi1nm4we63Xyd8msR01vK/PpCeGFcMk
fRwZm8MbqkrTm6omMOBX4+hhWh7O9iXQgfaFoXWSUPHWnnH7tMwuZiA9bs+25uDr
PK9iQk/ZrIK/tB0CTwmcbHzl5MhTutuzm8F8peg2epVPnZ/sm3KMdVrTuC7ODdZT
BlK/gKof2wJ+mSWaKfCETOhvkNLTuw0OA7B+86cpKQD4dlUz652IO6en207IdKCa
7ed6SI2H5RH9k5igzpdamU8uHhcyH5Lm5iXHVoHOwnIJneXobbDBEGQFjTM46t93
6Wgo/uQsH5vLHMRTnzhCObQlCeZKqraueZIB50NXxpsRiYkHPSPsQWMUHyKx6OxE
ssirfmMsx5lIahQFx7+TGX0rKC9QjkctJ77ADlyD1ASgbAH2WDyxG5waGBBZDXEP
CRKzde8MYsUSLdPK82XPNe+GrrRk80sOS0G8P5IaWm/YHwirXwcLjkIGRuUzgYUo
I3+JXdOKVhJzrk3ffLDYQX3QMMNkjmHEZje1IdR3M61cJsxihIRdHEpLGzHe5DBQ
7SzXJJ/ExSgPvlCEWaQpQi7YNkph0d1q4tahxrt4esSK1AFyqSY1jKJqiWuznKS2
OALFjcP0uwrT+QovQSS4xHKr1BejnoSBU8b6U6eTy90Tf3d+qnW2l1DqaoZ7q+Qs
Zn3lMdsv2X6zRpwqBaellDxslrW2sNCIUmg61MYpSWU8vCJf6iohxv5MC0RYzKrf
7E9/PJAONh1hVgtNwk6PGSAEQ0ay8eL0XGRRuXPVD43pl+TXb5zbNjtiyyqZO+it
4N9Fq1FG3/S0QDmSUQdLM+sPyBKItAnWzkXP7MeQkL+RspuISqPzSyp6Psj+Hv9W
gVZKwUIVkfSDigfy7D7G6W/ZGopzBbyBNJVwtn7VFw8/9owSJUJt8oz25fkZlTZZ
ywk1gLTZc9qF2OEMh/v5hZwlUWoVWOFvkiikl3Eoic6Ku87690VY88iPbeghk2tz
oXpuv/LCS0QwPfAU1t/Ncb01ceDIyN9TlsPgiQF4Xbqdo/QJyO5REmd/pJZB0NZQ
Ib8PP8bkQJ7xOXSmhmNmDzqgTcplgOfL/+W+26RU19V+ATMEQV0E/wsfxgnqNvMS
yM09oOTY9hVAMh93TTVzy7crZGgFb/YeGLvSY7FArgVGKC0u94ylcAXPg4uTusK8
3ap9CbkI6AjNMi4dSyg20zQBMPvvwmtg60+c7ie1BnKv2RICezVISrEbYSfd2OEa
kWV2Om1rtPGuMPGL0MOa04XjD/hBeWEZt5wvaHLsI03DBuQUsuL/Qp+j1JDcvyvf
5FiWsFSK+MIAEG0uPEhvcufYCntkgupk3dxb2LqNNeOMOPA5IgV0IUTJ2iQznnNP
iiQRq9Ao83qphsqCIdVrgFNU2CJZ1glmzYYVPY4pGJW2AengJCC1/1EaX90EOmh0
RXaauuHXGIkKeZH7zcEz4+2S3xO2/QN6PEY9qbIDaMvfgBHOxTP+FDcuKa5PA8hi
G6REPOj8kzrOe/7uw/u6nkYedYot0SwXk9KXL7adV2/DycoIfHfEh9Tc7olzyOsy
LqDzWB7HoKuKeIzQYAQykM8OxC1ZAIqUtaHyXRoWiL9LWIp3PJGznMNreRktzD3A
PWp6c6mhl1YH2oGMvg1+swzCNKWa57YXN5QgWLgXBIr1D+BZVOPLknVNHA5sTrQl
rHqB3LnW4FQxVjA7WzNpgOZQvhM3YMWA4fDE0E9Q+ZFatAF1WtNPSs84UD3++Cxz
sjJ8TFUemBPUtLY0y/oOB5Ryc6L+Yy0I7bIW2a04rFhafFLaHLQ70Tmc8dsWDTD8
qAVY9/WxhLNMTdrieZ82E8+vBPDWWzupbIAOOGmEotpk9K+F0X8YPnmUabP/3f9Y
GEQXkZ8VEKEZxIY1u26d+i+gkToVLG9M9TcJovws1mbb7V2NpPJ0oIHo/QRSajit
7/ngQ2F4zYPCnrRU4TuaRYX5mcfWXNO5cTrILwdf4xnMm1h0QGET79UqWHsHanKP
GDMyf1dZS9MzYCjAJ/p++/mB57tx8dkpT0XILQPNVWGnkkaZnRvvGdpSngNTfBC/
5nUdx0RFtflyrzJ6dg+L1aLDnyuXtQr46BsInDypPoJAamCZwAR/UFMfm9iwzjWJ
5s8nv0vVwwmMr6tB5qmsLB0cDZg/6BAtJkijUCm2gnOEvxOeIl8eWWVEt0C1ZDko
xS0caAH/xRHPmFcAAfn/72TtZA+K7AHiIwGbWuu8XR5veHkpovPWMPxWZy86tbYo
1GE3OHa9eY1R/nNaQJT25epTipio6cooqtG9DqexNPWy6ZqsJJ+sh96N7aLpbydV
CaxrHcus/IoVcsOj0p9zPX8Prx0VP9wcUPnw4zgWx3MlxNiLwNyi5NRaJgQhA8VS
lpoLUEfZK2omghU22xIVwrKXfpPqb5Romnu2Q5DXiAwG+IuGT9nMQsM+qduw5Hge
BIKt82o7VVxz5H4KiqdPkyFw6f4z8MAbHSeT0ZpKGmO5TRonSuK7ArTwzaos88WQ
TS/iJlET+8gyWV1E9JIvJuPjCE8lR4Vd9Khzo4NofAOSK2I4HU8r9KylueOdUlkm
qaR3Uqggjq5WiSYT01bhpWRgy3R2w9N+d+sL6v83gjGBi2mJZHIB2z8n8wxXH3B7
rCcZa5PCn2dsqQ8wQRwN+Sgd9CMOpURStrv9uyKgc2hx0jtFxQrNRlr3ftCnXbMi
sQeVU9Wi+Cy5ArsemnQZDxzE18bMm2gcIqu8aSKeT69Gfarwa5Og1Py6FG6ta12n
0AaRjr/F8/7AQujDN343Oc5GBzfoce9Ke+j+rUk4Xf2KIBuVw66+7ANJb6HXWV/j
Jc1SOHnkcEAO4zlGw3ME8nzPFIsd3XLUZlpALpDSsSGRp/DNNJ5LX6S1mzQ1mba7
hofxLb8GXjI2B5FCH9i0bWo5UAZosxVY+2kofG8W/dKTadVd/xH+uxzzJMkHdvCl
bLb3H9jUf7l9/aMn4FSHeifkdvpcKrgcNVVpxytzEFxFwvXofFMyNvPy2FNYvexX
boVY56DNQuat9azuOSQ4ZAM6eJMp6Ml5vsvwewEVRWUzk9r0NBIfY4pbeTCvj24W
hF4pZ28G5xq10/sw1mBt+JdfFFxmp6G7DuthT+WGBPH6n1Sm7XlcA+Z+hyAJS/7N
c+z4P6gBX/FxuxfpKeO83LNl+S4DKZrnf2J+K3IRTDm6A4r6O5QvsOfivsOJuV1W
fl8veNMK6YFHsL8X9yiPGfR7x2GotwpRB8dMOIw+w0WOLa3qJRrcS1Ro7lXa/3CK
X2eXutHX1uAzTP+g2cqBb6Cuj4UTAx+gaXHqx6qw20R5vGIEZswGddeeZwbZju0Y
NzeuHLxh8lMvS49ul01r4TK1yv994eWLodN5hEge8sP1mOa44+HsmP3caDv6323b
fMZVadmo43QtaE2b8IWIlCoJyb+7VflpBR16C/CrQeJ29sdmGvmpEQAgXZFCiOW0
VW9+I/KF7nbrLfINyVWLE87WtRzS4HmomLv+Ih8Drlas5lqbDDU9Eif9JUZZjvDD
toSesOx4WSZu5Eg/uzJs9PI0fUhK4KGLzxekscG6V1ZHF5QsfkySu4XCpG+qfNem
fj1vswecIEbPn9sF9cICknMnIpPYVRwzr4OdAuyYM2rEcNGVJCQPvRDK16ag8lsp
KtjiO8McNB3DXpJqN4Vl1ahXymFih4+m6irKZiWS7ao/iMGLu/McKhCcdSHQB7/h
aiREV3Sle7/DA4zlfYu95XmjfyLjgd+12ndR/cp3UYzcOq+NwSsh+xUqPmWTkV0j
TscAs0Fuc/b4QIljdwfcaKCh3eZ3oXHCqDZcDNNPJfzeviFp51FVd1KqglQUbvbC
DUb4a/7D1ciOkclDLnYho5l5WznqrNqb5YmF+T/XmXufOBwFPbnuIo6ybvUqlc/s
U0SZ1ynfTp5si7rBTgbm6GSNbpGWIn+NZgyhXr1lW693j/bCAL9c15fKImvBLSAn
4e6SUlR+aKIB2e++BEjuMFjB7TqDl7jiVC5+vx5X+Z69zPoVQVFWBcj9eqLNadSZ
VLAJ8Q3cLgpw7eOd/puuwra9wJd9XrZtwTZbKHC6GNrYJfhr94tIzBL9DqxjsiSJ
e+AU233VVj2kpdP3XXLsXZsRnxY0bxm37FhonAGTwXEwLHnI4XDBthDj5jIeb+FI
813jD1JNiCe5yp2UqHHpxsk2NKrW4QcBxP4xJnXBdPpoxyFnjI7rr6HzwP0aEpP6
MZcRnMG1SVO0CpCZmupsHSia4bkFXqamUOIkh9Rqbmi8X6k81LpRFUfE99f89bSh
3524wDPpUQfaw50R+1RUQpiec7pFZQJgsfjFwofAt4pTL0gQTLE9Ic0WCDyRjFaz
5C+yJANgEGBDtUiZyUtYXUbpc6FEen4v5cMiOlbpQIbWzEfQNSXgDXYAdT0J5u++
GmBQhWC3tN1XgtzQk7T2F5nVEwyzix1P7PNPmHf8nOXePjamrkUGFqsyj/tKD3fy
F4MGoav//OMiK5gLCAO7gGplAwfyb0m1UnOFPQ55WoC1BGjhTtkAnORmA+wo1Jjt
JPv82YAfLD7BYTb6GrDTqlPxarNtH1ZApDPn4g3EK52SwoqLO4hkIeQeY9Tz27+x
y/g4rIjIOp0E69mk0vOsimSEopbkHiNOdbVfkT+AO7jk7pCecHZbaBhjvFVG7PDw
rTv5LXupQlNX8b2hlB0iPsYU0VKhMxrA7xt5sKMEyBLSbLncIMDG94cdtkNtA6zF
nokfKUHnnVtmRUDeOF5F77Hs6EJD+YcJU8VUQRSiZ4zl8mZqFGKyozxUmERhJYgI
f/K5kqd9mEQdNLtD5RHKKtnAgBHH64xClEF85Iw99BXQdU2GRvilNKCd0MvaqukK
NCk8i5CZyQEVsURcaSXbbiSqSC81QyrvMkCl62jVwqA4jS+gPXKcNyHwqMWtVZHi
EGfz2AHDZdigOsfS9dK4d3dBIMNtEMOck8ys4keauhBhKLzOHkEqoZCZtwVvStwx
cakSYfqlpBLebAHyYYCs9Mu0C5h5y5PX0T8bOVD8hP513BxHtrKVVihCNVV0N9j7
OU3xy+As3omYWDDbIDALeFeojRXsby5cPlO8NpxmXIm2Cg8UFFz7YIZRQCrGWxrW
G8g/ZMoT1L/AGHpZu5bVu/0kw0lAGv0nJLrTaoz6tZsIT5bbs21tI6JuKYo8Q0As
EczgHsW17DgUmyHGopFVTF8wu2NA8n63XPLKZ6HcPZ5JsAzFTNUEeARKHt4NBix+
kKjAMKqHjJ2ivFW9eNZT74f0S+QbYXVrAiiaPS0ZMBJNUgCutMnJNdIcGYqDg2Eb
xKxj/lmbmduIQGs7qRvLjtchPf7a4yEVCkkJt22bw1cou0bJHtPl1AvRiK+Ygki4
NH/M7rDRkdiprzu4efISYFcDLFt9gJhvkZBA2chbD6MpDo+f6oaSptqh8hzUARaN
RVxubH0r8WrigdmwZiufRGpFwC2GfJB/LUa3TiD6s40oO/eHF5L7eatAudnsEBYC
udTLJ4tsx/tyxJ5yIrz3rAZFl+mIXwqpQbRmM8eUWSAY7Y8NU9JAcKCoYsIxBRpY
34USM8bOoRHnw0TFjYznReHoK4kqrLA6VVIfJOQQZiJ63Mc95Ad2/Vnds2Hi/jDd
BH7DBtB7VHtv0cbGYxXFBUvqGzdaFuI+ajH2RFNIof/BhURoQKyvKE1+I9gyl8uE
kvqO3Kn2RnnQGBToJaG1H+YAkVmjLjucPV9lieIXEGMp6c9HCBp/goAKXDgJxz86
NS36LOV9G9XTuJTSCAz1lk6eXTGy0pO1w9NxseBiYbHMov+1n7QHLSHtj3Iob63T
4dt0OPhZdRH1HhJVgjzMsEtplg5wxEFzbnw5K7x9HshNc+AvfbhxbTvhZphoVEyD
YWvWEIzP5woIpYY09dqmWwe4ABetHecQfDaaTqJqfDyQTF8OTPT8IMra3s3EFeuY
9PXb4wVlTnaGG1tm9R9Gj1ckKSQj9iBh97R+RVn61dQuXhFG4LeuKbOWUoGUCy1Y
rq9Iy1Xj7u/Pq0w9pZpvDuook5qmuDU9RDwhHJCoFGLj7V3UIVZSjm+Eus1dro+/
U+L41WIoBchC20wTG/BOfVqScnulSv1jFCsvA3VgNFIVPq0JO325otKQGUJ4dlb9
Pxy0YAIJ4krt+J3QuToJxJYh0KmEJEkFlbIgwqO2uf4zQ8wS64FmiPOBcIHdBMOn
cslcgBzFbACZizhSZERJs0J3d4zPULQ7tbkaGnZYgeP3SRojQcDnVNtA8oW7JId1
OcJzNv/3VNwBiPN3eTX5ocf52lOHpoSFW9qzk9e5g9Y7tMGk32fshOLOk7xpCsOU
Z1vJPk9ZTotL5zDsWEQfDJXR1FYff+kvQ2VtZ8S6NpaOMpQWVSHpv1ov2uA/XgsH
r9YsG/7lcXA8l7W1JgpgmCByn+i8hil35RmbHg3OQbjr175XJ/BqcojXIen33EFM
jmnRB+4sL0N8ICXlVGGRotLPN6hg6P1sYS7VbYi2hUOKD0ztJ5NU+zU0NT/XUg1P
OuYaUcM49pIyWi+iwQNs+usg8fCEZ5dFX9SBgcRMzTW6NUnuolBSVcf386YbzDco
4DhYorx3YyWTKbbt8kHe1gdfjAbVWIbNByMHTeKnIsQVHj1mINMhJ0g+jhKbCO5i
MMeTTbWQ336fcdgi2cMIr7euqP5UpUIhX5olp2+HKrwDz98Mlj9eP54qZ7G1fb6X
8B4hYDWskW0KzRRtA1S8Y0BGvgLZDr4v2X7Rd/WEvLZZB/2y8JEQWDtFzCX33hX2
QsWT63D39vEJGS9Df+0rOaMJeub7jFrBVF80TL6V71x4ey8zgpH9lyqdcULEryxX
hLa+BgmCFp2JPXpRZ1j29LcO0UibLYZQrE8n6VpTzQ2/N7oK1Iw3Fnpcdf59ZFrX
mvLxwm3XbbqeiaZhAFbE7Pgq2R5DrDNcYSLMPYTvpgkEemBbmedqEGVmC/abmYCY
FAbf1AzG1uO7wgSQOOXJdCB+52B0nIQpxiyJ3gIxsBXjH3FVqCH9SJEpWw0Gz9nM
IyVhg50AR8eMTcA1tyqAypWNbgkRvORyEsKazWlJB1b20ed4R/rJdvfAZH71MlXU
pb7FQVtqV7bP8ziJIAcCqEzx+UL8hVxrPt1zTnese4JWiyOjWf+0Q0nKw+hAvXgv
X9SHVJ+z4iB3crEeXIWBGzbtAPnufxdJ6WlDSxoByAmHgBikGCqb/tsVZysHkQUw
TZgnjJt8rg5M5z1WMAeDrVHqfYMtandV/RpomNYnBjJufRQGD5pRHMokL2FBWRJ1
0wN2/iRjhOffv7fxg+SkioW8+Qg2rHmpODuj+CKxho/FzDcd3zCuqgkFzDIIS4HF
DcSoyt+IS2rAZswBnnD6SehVakIcx9xEazl/hA//jAq/9AbwBMtu5H5iP3jKuiwD
kuCxtl61/vhxsdwNFy5RBKQULupQidj/J5M5cRtGIeS3XclfrGKaTXVCaolocRnt
7B0k9Ijxv6Hkv7/CXQ0uLty5m+LfB5RYUuAv3xexRiURYf3yITyqOKAuZVVd9MbT
fJTigc3F4QLC3p52d1LE4BuZKbStA5xdB9+w8es4sSv0y6iOq7Zj7N2qYyWokjz0
bmzNeT9OcEeX+tT9KnhKLs37fOfoR1TO5dFpP8obN8adWwFywuHv4x3+FUxAUPzm
Y+jthL/1dziLEDvxFQ/yOwayV041c9XxHWt20lfbbr8I/pj0/BGzSrJyub27EGz2
J0nGM3Vv5lyDWZ7ZqBQmXvkLn3YAXiH0E+lgb8mFzq9QpwQ+6JbHaQYHT5mJnLcj
xg06xdhanN04P7apaIjZvRu8cOrRSx9a7ATIqw3V6Kh4gKI/LNPSKxldwWaVKIU8
x2cFWZxXg3euGv/s33P2ip04k+B42l3/QH8GkIrPnTwZmUW4mrnJKW3yYJbsoLoA
lCvg2zHEYS8i77rpadrMBbTOVXZt7ameLSokZyFe3b8/RNe9H0a+ijLoq87ggI+V
UAaH6ZNQAE7XsJwiv2EBlkp+eFMRly++WNuNKn+rhscTUtUSz1jeyPwk7Ebm/FS7
BD0BxCx9njkUFM80WOTLOi7TAMXHGlPBGGt0kuKyVFIbmoveejwQTaTd+YPI5jhE
nGaATGXg4IacvWMNuTj7KkZgyhCCpbbelOfucyq9eC5+JVjyiFJrwWa+zELfa/Ht
urKu4BJuHEDtQFzaDjKJxymtz/pqp6tp3FA+JByLxGcjbzkXlI11xux3d1Fs/sQv
cktGCWWjFxO6ACXYGiB9zi+lr6nJLUnSCe7U9SPkBLHHHipIeWbV1FvE6DmNV/uh
xI7nTzKxYjWkAX7hFPzmcrVgBOrWrOZ9JakI/43ACe+Jvuq/5d7WRYeq1afaUqUu
7aEK7D+P8I1H/qnEmemxpg1aGREj3/I4OpGN++Ll+2Kt3drFO4yGY2GdvPkH1Z/0
cd2P13d7IKqwI7glKhMfXFurUPNYR5UP7sOejeq+opPXfdUX7QKXFAsKxM9L7tMv
SHTiDQ516AIQjOCj/fjwWaSKmHx+xoLk3fCzCqK/bTmC8L+4ehHdr7pyabyS7N5p
QV88412/K5gtBW8xsiWM/qHn2VHcNGuAC75y6ErgjInXM7VuEBptgux9+utlI0wx
W0WeF3WE/oHWHbDbX9J2WIpKbr2Kv3/3u+TgNcAsOaZG4uhzcDuC52LmiVKEUY7m
0oyboOJN7dVLpy0n/gRSpaQ+0t6HlEQIh8qTZc+VvbqbSK/INQqkWjmL41rCJSuH
dBaiTwbCTcdCkEdDmEWkaNUP6MF3AQ/jAdF8LckET0JhXwmKmMKJi5klUdOUtaSX
oRpF3KoEHHX+K2C0uvT0rzR/MhXzCmdEulZOO585FVM=
`pragma protect end_protected
