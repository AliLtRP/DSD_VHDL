// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qJgU5obMcd3Uv/B/FUhFTW/CTrKFQHtS+m4DKSR1oHGSEn3rfiM2okvALxS/niln
0C53EGRa+XHdNHqKFblyVyFwXAdsjBqW4kGO7+ciDedjj1GwcVDN3zD8WJwfnOCB
qtX5PmqHV2vCB0xU4O3fwKfv46jcJg39T3KimKLK6qQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19248)
KzGRtFoypwPIZfCFfaGpPp2iD2UJ3dq/8qt8zz3vQrmTPEFI+iAFx+S3hC3gKGiU
e5hOwt9DvADCpIzJayQ4eE1r7xnUy+wCgQ8sRGXc4sGDVcGDUU84zxy7WAhsiMqe
mUgg+kv74qL4GAAlL4upETkDClnujTa5gQXmUc6utVESeqh3q+I1GaAxq0uuPGBi
s15ENV/6BwY4JCx/0koDzksLUDHsvbdY/CTp3pjSXRh2lVKYruli8rOLVHigpiH6
8P2EUgqLYj0SO25lZxAQlBJANPtDS6BvhOIyKdXqnQgSo2PlDv6doVNZ0RGgckRr
lhMsC+Df2aWsHAyUkp1d9MsV/tvHuFP35ipG3tzAXaf64MjDgTGfDMiWhw3rHaIW
gXNz5zvuxFUvZi6i498W+S23gfCKbh1D/mCCYWaEgFIHKy6Uthl1mPty+rYwe3nX
ageJ0ZPaMU8f8bEQM0JjIinMSRfXMqTnkx1fxzHfqiL2FLMJvWA3GySF3q/d07n5
ERu2iqDWk4YmAb/Ash0gYNmHaJYRD4s9FA+Y/+jI1QZqH/GsuA14zAuLDC9MikgX
PDGNh7HvdL8Ygyh4X/1fh4gxdhP0fQ21M0Imoe0P6+D0XQ2R/EBp6PKDk5ftnmg0
cjOJH6TFZdcEID77fKazi8vrmDHOfYtnn/EZ22yi8qfeK/bZXLelvGBPuJhdCJ67
MH5yF6zQKXd7a8eTXCOZaHG9MwjfvrBs4Zb+X1ci/DfYGrnwiw+IzMVflGYGhvg8
7peCziNzeTAbW/ZdinJf/zzVNEm/zC7h3DlWrK6AGZnPgYXY9MIGGNmxVm7tEICU
cPLqVRE4OWBEpAok7Xkc81wcc7JX3+PCQU3ziUm16rnE0Imlmhn0Bhozn3ZBDTpU
J/8XRzOLdFi2U96ZO9MeIdN4T29479IV/v6L31mKd9paVQisl+DHbOk0phJRWCrB
DgwP/Mdznc2kqLpQ/z/sG2F3xgF+BG7vSUKdclUXX6bWeJp9uGekh56jM/CgYjCh
6QRMQHsfDtj4GyIf/fjE2l8AOztHNwhemSPMUbGshxpJkb+aKzcq78n4RoOSkD05
zuv+dv+yD66wcCp78K5R+qGAjs6nU9GiKT9+ggkSXix0tIaKubW3BixPH26LKDLQ
mYmmVo/5dd8QMohNB0IezELyK11o92h32I0KMG0b8dGBc1uuWepBjhwfpZPpJ7tJ
iGqJDQ8MLIdnl2Cl03NW/ifMTvgv3/9RTeImCcRHcxp0RlRkNDnx/ErmnLlp873S
IW3U2f5Hd2yZy7d8FJAIlPu3sPLr8Q8DftYxkmuDUE5jxaDlfpnDCFCjC9DjtxHn
brZcfb4wm1w4oVH2cAidsdZ3siK4pSP2RCMsXHsbJz8pQF0fy/lJtpDm7KgVsaHF
LPtGAiSpNlGyzfcykELAJmneMrcqFuyfapgeIKfGRTJ7PFuLTni1xrGyzRXHwHXi
vf2XAAVeSjDJhacxQ3KpkNRsQNxMxb3ojil0H3ihnICe0eoCZHbzDSlksj6XmBc5
kZChxZIjUnH1Yi1elqKQc8/r/0wWZgkilQZF9Y+bk2pcvcbM0wyFusKyuUXRxzef
ws0JSdJnXv/UmOl/fCW2G+wpm9Rz+dq2P6GvafIOmkpY2WD19ZIZLM7xUcOUeNrX
YpQv/p2eFLvmOmKZl3Zzv1atZAPNpx1fmLjQcogQrRsxSQpcHJRDjOBE1ghg9ExQ
AifeMA+s8RHFtAcdwGVryJvHXn2Sh4suSzsjs1LZrJ9IzRDwth8a3a33QZC31dDy
A6nBCtXtxkajvNL8BXb+gn7tbZYo59hUmUVJC+z6MgIO0De/DagQw7rN4v14Vr/+
2xb5G5SF8iRVAszOXcRk3yNotlbJHB/us581CQrc53g4kbOwGuCef6sHSSXEfIva
zsLRHUcrjbpNIJ0rzZ8rzQEJxkQvKpqrLO0GFX3axPTMFy4HWQ1ejLYWI/vk7UIo
OtTsLn/MCbt/WGZ3LfczEgFm/4/iHTfnwuqX14JMPFm3m8P2C3iblU9tK1PnD3Uf
U9bcBUlHFnyzG3K30zgn8A5OpYVAvl5JmS9GnbNtP1GmCCzvudAiL5nn5XMI4aoy
H0Upv1k/DydL4QaHIj+rxivqXqegZi/FzxC9nQtY4dcRTlXlwp1vRTTM9xxLbrep
cDBOUM0LKcwgEETzWviRWWx+Bk42nmCl9Dzp64YrPchTo0YHIf+MnlmvKH+I6XXg
0YMoBHQFFyIN0tippU0jE2fK4vDuNOcy3lmCz/1v/Cr7pp4+isvCRM3//6oGSKl/
e4QTO9t/jt2Ma2hqrsL/A8zPqs9dXInKbhuxByWY8JS3o7VvhFAmwN66Wo803YAR
GOuojUF+cerwV3mZS0gfhUNnh2Alk0M4Y0wCwHRc45um1RbzWWGHxBJtaUQtypLy
KYcQvVwhWtSYXtAK8QFcK/AB1EBRtDzCBT38q/nEY5NJgwq0DVTw2rjq3KQAT+kV
lQj0y1ZMtXMeOan3zM0f+dZuY40paGJ1GYdlRWECcm5at/aJez52E6+J/5NXpZ6W
NOK6XTd/kKQ65RV8QyFBoDv9HWrCLWxzNeY2YUm5Nt2lWY9k8Cz2Y/dVemEkXkit
GE/W6maPOD4nPjgC5GUOAcAlm6w5mzoSC1rAJEn3eB4yqRuCp1ITBTtFmLLANv2w
0oMoEBriN5z7JBzkQ4P9y+Y8uMquMol8kLl43RMlSfZuf0l9u+ZVWudVOXAAe7TS
5c8kTdo+8ucwAdeho8H4hX/fBfz1iFVkWHb7QT2pe23pzbzq7y+fQERjOLXfqhsb
9y6hu1K+b+jchPo9eaJUmwvc1bXCj50AY8Y5mycdqyoj44HuCrCmZb9jIFlvyK1R
+Gpg55ittkdTlVhZ6niD2Fc0tUXwt60IsUP5k2KWqRi6hMHPD8zJWbxp31VSTAgl
uhJEdWS0eMrBKyHuBwo+LiSGwmRX9uTw+aMVEjSZj08NT/kHKM6pHKBUPt+e+LX2
TOfwtyb+Jun0PRur3M2M8Zdvnv4pEDzsqN05wXaTulfXp+DFwojXi129Hifbv/aH
Ef6/4oVuhDaoOKBySLZzVTXfBNKjii2QtRferx1q24wgM2ad2BtFdtksuQ/xdIk5
611rEgludj82QT/xwwsZOtb/95aL83dZ36rMIrgtAJ4CeJw/LpsjCvwdiDYTl/ZB
fA7X4N8aClxRcp6/2nRz65TNWLojddqKkcTkahQaNwPWySf8uBUhMcPgKfPsts4r
kIDwf0qKEB00m6vzHuZAJxDZD1084nkm+uZz45pKCeGJdOnwld8LNd/DLHDlDRLc
bYsBuagULCWzClqy1CGQ+fizXzF4Ab6RVzGbDaAFHliG3Uwkui0xeKOt7Ma+oiPK
F8ikVposmunmvLoG14Vo+YO/uPDUWuyFXAyp0qe+QWnQf16XweGnjVTOs7kWPnCQ
IM/hOVd4VBPD7e10FSB8HQ75k7udn5/1y8DFNFiE0UpKWt2JXR7CBh9LfRlaY2z7
nT6J/DalvJ5rnAQgvZLedCAdtiJOIJDpBgDhr+ml90jFuYFl0DXNIK9HYP/MqGP+
1ZJZdwVMVObhlXHIYEkG5CWz3NzQrqtU02StILSkSSDjEOFC4pcLXdJNTob5uRX0
bcXKlCGA5G0bVOOXfoinQLNNXrN5Cc/cxiECs8vrbueiZ9mZbfMpgAY9Dyvjg7E5
v0A1eTs4RZP6g9ihNIiVYXM8ZESqKf3UHo3zWYatQnY4nwbO4t97PL5dRDrc8WN0
vd18OQGaOnpZXDEp4BJv8uOL7rabjFqWIc+UWsTPQuxr/yMfreQ6KeWJd0HseErj
ybHYT4Us9X5aO1ICgou95JBC3WXVX/L9WAdrlu+I+PdhCb3TqPPrScP8fgzfxNAR
vXYp/5iA+LCPyNSc29J7ET9PAcJJZHwvhhcaMfHdzusWz/PiBJVqXOwAbU8bYXXl
BIrWwtURNL1m6l8eZ1Jwqj6T79bCYdeli3VV0DSOO2dzAJXmxHz6OHBTMARpxNcN
N+NN3MGgIGn3Bhois1jp/DG3dI/MoFbavgEETDAOt9/vauZYj7Y4MKdwPXfxyUcJ
sIfUQeYU/FlKZQbo4stWoYnsZ6bVbUg8OqH+PDUfmBg8dZrg6449sf7mEhB5ZVS8
Cs91FDgpQO1753TCNSCBNRRE+sAaVZh8LA56/3q2LwRgGFyM+Ln6ldEumoKoPRFr
53SF7JI/ic+ZL73DLr+5zBnJsD+FeD+FvEh/5YW9vugXLAFUj+RFAG7A09XuI7cb
ayDsSJI6xtNVMCmrces+KBJLwv0dJA5HbB0RXaUJkvr7uqIc8lSMaRTgvbEHpoW9
ZvxY2X8fL02TMN7PqiV+G/nfH2NWsG4g2uig/RrUfYOWgW0Pu6tHCFLEVyA28G3t
714MVDyRLb5RCNnY7lMXqhzf8wtANyeEwLHEdkesFotLCsqfdOhhXQtZtzIbvdz5
uTPx8mbc4iwWJX3S0K609v6a9rNfxC1Z8wYs8besMUqUiUcDuYLLo5/QTTOR85D+
WBpXynci/ntElo7A0QFznsak3Ic+yRw7f1/Rom2yGxMbQF5OCa8ODoTDJEvPAusM
YkVgqEHHa6U0quuSAcW6F2SMY0C+lBsVFavNaDzJH6SFc6bBUGqwTyMmmpCtbdhI
vEaegHH6ya36J0a8VPpZzb9MRWoDvZVJ9dC2uz+C/DyWu5dHMOy1WJiJJs9PiFcX
wuuPJJYtbyKqMZMffXryy9ZrBKMF1Yhd8GO2FtufPufu1payfJpH5cd3UM+7M5cp
Mm8VV3e6PYJlfjY3QdeVkGjHaLy7JOvz2Hi37MftqCOLU+I7D4t3carDPeemXmTH
kiKZE8vkqGkkTNuL/q5FMe0b54ScvPeU8RPBZtjiUIgM1V6hAjgJ5SbK8j/O+RCk
i4qS3vxZnG7wG2a6c7ar593zOnkI34cwfZ3GmXPfUUxFJqizYdhnCzKk7QAwVF53
OFh+xjHdi+3rRg8hnwc69u3jrEcyNumXstwhL+YttIXqTHfIjPHthi+y1kItqn45
cPBcgi2tJeZ9EFcrY7C+uWJHhPctx6R5Tb/z3VJ6YZWUtWJkF64buFUxmv3AuAxF
qMcjVOUXiONdzyHtoNuRL04PI6jscswleHLTeAtgtCrrSpRzVeYICx7r+1CiOXF0
mwI3BA1wVirpoPNLv4ozGPjV288EogeePpya8y4tI2v7AvScutvZTtBD9ciTiIAd
AK+KYHOYIRV/gClMj9Qlx1VAZrNRyW9zqvK9sjr5WOOPo5SIXqZhwWgwQggENLuK
5OnJyhvwi+6xlCAeX50OOtar5O4XFKR04DVrLrz7BPaiBLmd6+iRywdJJOFvSkDG
ruspc81wRWsc5/ackqjL1z4cMGgY+yVtNyUgj0OMeLQBbfrKNnfzI3WFZ0Z4pYMt
eFqO5UE4CWZ09NP8hgvUV4g+Wf5vcX/hmEbygcenpP86sDjJ0+VKOivvq3plrRGD
wuokGBaoriJdLaHpPqCngpG4X04UpV1BeD0J5k2sBBwm2nl4EmrWUT6COmi9HAX6
8Zcpl9XGKaPMiEfNHqNV7ZOPzMAgzjJQDnLWEtrS6MB/MVJQpOD/tAGNP4bQtiti
pHQhq6OiQJXlzP3Lc/TB8fdxeACoNiTNLfr5bcSQdiOyKWL5GBQk0Wv2KxhO6QD/
iNO6U3C6E05Euvl7PMzQ0gYdDVK5qNLWcMbnuoGfY13aVtSKf/7IFuxoATV0ATop
U890fUUpgIdiJS4WUHtwsGXMjHDhVD4DlW9/b2k8sf7KsH/isJNEv1gjvYs7Z5vr
iwSIIWsBKgj6cWA9ikjb1aMoxRcOeNFdFHzmx9RxTuK8pSiW6Do3bearzBBbQxsM
7YGzgNsC2gxR0DaoyabjEE70IgQHLRTp4xqGfW7m6ndfxSKXJpswIzQ01YUqzbxC
MiS7VjFFdqoPiVHH28b0Cq64ADEUb1fCjvr2QWh+b2AeZNRdxrXLM0TXd+eJyhPA
llty0HkcBmcxHXYWdTrk/Oe5C9/m2Tx6OrmBo7majUAbjbSuhoLVNhUghOQVyFwk
N8wHtY5z1amK5uKonm1qbwzTGyviPJaWq/5Wn9PDx2pSWyYyQs1M93pgMYjMNxQ4
Dfx+RhE0N06wWRzckGwYhW0ruBhx1Yit2YelteLRWe2BWvK0FHYU7GbVp9SMydkg
AL/Od7PcMrt9F8Xu2C+/Ivd1o29S7V8aeSmeDiygUJrmAjGxD1NxA2Sb4nR07wK1
PapBiP0qSDEX5Gxp95LLzhE4mG9BUoUE4ytbloUuLmmB4zqUAjSBePdcn0+KaPbH
rc+mevUi89zF1cFtWDSDw/fNNvUi56HDwGEpDFWQ/yOpNNv1bWuSVCPjYmmzj8L2
M//8HXG9/Oeg5iNaDdZ+xIqLXeBring/PV7eVYu19PE5iRKt3DvqUJXsA4EV00nC
j43bAFUj6243AtzWce/iAQfEMY7Ry0nNLpr6kMnNnLvc29lfdJ1JU2dXv7oQe0x4
iEXvE+sFGBW0dTSpNT8kqSSzhNAEkdM+eVA+G+F9uar6hj3HlEoWmD1Oz5L+BxMD
GxP1puW1ibKLZNskcchVO9qrhNjRk3++DVFWZrBA0+p6/zb0Uoe+kjlKNL5pJb8O
NgNxh9CASNdsCLBvhowzH71xGXB+yaQWcPlwQH4uT0eJ0srvKldKud2FG8oz19JI
JpSnsNK/kUuxqFhH9mTRnQOlEIp7bVGL9sGcENa9MEZ1Xq0msdRruvnzImuW7jRr
hczQssVh3eWMv4xfGIEk1pO0vVOswMPBQDyq0j5ehGCoZ1FHSrDG5eGnyMXgNCmy
cT3Ix/t53ZfEib0OsA8MEMOvUzxWNgpb5RGcXGZDWbAkf91DFOBlYI1dVfOiKRWc
9ZAqaDedo1uS5s4Ug0zyETF0EiKyRffuYEhuTH+lPzu0Q94VjacGy+B1jZkfYqxG
PFD/vcGHw0ATAgEPdr4EPhqQ1hq493ICU+bXG/8rqIs5shAW4ZDmj098L4MHlpIU
lKZwUZv99u2QRfB3tckAxOquFLwfrCcNxoc/bmmBbdY5C994B8tOiPi9cDCa4NQ6
ubfpxm9K3T/TyLMecUXFfciZtwibMtiJTmJl7f5Yu/wOC3OT0dc2WPkIuPjGewaH
Z5x3odFywTdFQCZgU4JI+o4j/7Kt6SL72kN2JIVxMuVi6drVc6qVAtwGKn4MJn6N
WqsMqBUiUp9WrA+sZJdbcDknoKG/eXJ0PUVtcU/KejnvCgy2WyKbXIdaAFDCReGV
YY7NzXMyiwZgg4HxsOW7wRSfHygkB3kSmdFUJ8M5kM64aq7SU6YZ7YFz5R76pjiQ
qLPqInkhKgx/wnaGwb23j7eLkG3W7R3zrf31dk0TzqDbMwpKj/axxpBWXa9qE7uz
7d1baHOqIfs9457CpoVdstI660zref8DV7l1v5mkn+0O0qYoF6Y53A9lcRsUfVeh
kKtH8rCNl0oMhYLbxGgBQLsIv2dRvMXQwUSfHcuKmGm32d1RloSD6sYSMGKX6eec
GJA+KsK4MtmdMK7PnUGXtLmVngRqrzFQnowh1ZuRAPDNiFvJapqIm3PSDoJi8KL4
wI0i7pwUD6rK5zynHfksIKY5ssVRfjZqe2oQCciqaqNkmg+bOpH8wgStaJa7/WN5
rcgjGw2YhcohJi9epLVOnpbkuIEPT/hBFOOwIOOsFCbLR82TOI4NdcROlFQ6ahei
l+VvXU1iHBOXc1SWleVr2WJR3k5YYUyrqM1QUZyQmsWeOcW4MbOzbkyxiDvtvnD4
PeUAtddyaIiJ/WA4cu4GKRVFzMqDwBu5fr2IgtoqLECQcJtfEq/Bwa6m5j6PhpvY
1/qaLDYxYf/4boWWLtTaoBSLPrQK9Tixfc1T1MxRHj/70j21E6Zn9Qjdq1qKTwBW
V9wgJZgjeMBfiOHN3oDhDE2byQ5nL9ixwWoTNqavAOYegLuWXlEH2vsyuRzaFeSe
MK+8Sxlby9g1PngHxXQPVzlCSxyEGegwkykSyUPvCpBOEXNuVqyv5kvyv0kSQEof
RVa4tddAtumR/2nUtyghIoRH1xj0lFQ8/hPKeXZawwGCXPGoorJeXxQumvqAl7S2
QEIP47VjYNwuffH8C94p5zMCC7Iez6dVmqntTROu7bSNRgFpE2wqokwOLd9bWH6T
5g0vBKCr8oREt61N9Zrn8vq+lQ7HCz/RiCSR05FotWt8KykIc5Rg+wkIMOfc9ZUx
XwDODLl9w1OcyUqMJ5AgPigbBx7yqUu9hZ5E3qSw+6x6CeiR9+Az/2+6hyIROtOh
sdWzDFJqDy+iBAywoNQriUL75nhc+fvCyke+qnkIJOmXNSOZmQWdJD97xRj29Fz7
Wsnb1eFToKXAAeT2qYAScZkEWXwZgDlUa3sgO9Axu4hKyrG+krqypLkZq4A8P2Fz
Yj3owDVxQwzBLPir+/32g6GZ3CfJDHuFnTNTV/FvWZ/eD3ChUwOZv00kkUdtUWG0
p8nUOOvamG9qHHVjcN9QcTZC022Ow9skwNYpyMR0V/TkkyeLeRKQsMjuilrsmgYW
+h8R2T8Hy9+OktD2XTfAKbh0ZW5E3aMvwFGpnX3MscnVE8UR1gbaemEFn8ITmmnH
/8HurCwWi36JbVybNk7gYs3sOmiWhBef9DTDRPtJxiEXOM3bphaslduSyuKPLwSc
4eMie7KZEdwoJCJtjaF6NickCDe7ia+iRHl17kXsRCEmgSm6PFE7jSDPxogzk064
FQkkBa5AY8mzluqg/MUMMe8xhqBO0Jzibk8pQCAkXLjb5IEvbowG5+OMoVR6ZxZZ
TScC13NT6ktZGIWG2XQsIoSRVz3Oeczbq5C8qX8HY/UXAt8GlVNf0xMeixguBA/o
vXsWxDlC0CHS/yMpb+UGQLeoH7a7wj6/qYJQQPb4MvTTw40WXs6gLcQnJZ/pBDGq
moTcYb56WcRex7rLI4Bu/AdO8FvrPd1KRnR09ZUS+KADKIl86RhHkefMy+SOkXHX
IreG/egliM5UnLjHeQaemN0d1y49soC4IG+I9gW7eJ0FvdxuHQCVL4/21BSBIOpv
ouBlDrL7uZ36/VqlQssXKdYEQ/bnnCFF012I3wzybvSViUh5gE+2fU8W23Sw145b
tBsueDVGyi1PrDbxvufzgUo6ARz97CZy1BCD/crGhjSMOMP0ylaDt6DrmJhzXaEL
kSPdgqbAellQNX+t98V+cwqkyOeWY9bXRD6SoRVa1ez2xxls5N4EtrkKXvBJa0EY
9CQllAI7ovnSsChtgiby7TdJgYEscZl3YnJUuPmzAuB+AcRkDpssSpaYvu0L9ymw
Z9hmyJgyhyyXjLbr8YwFxDsap5EkzA4chugvdx0KBTwrO7LTdDyNYBRKBXD4ccKu
6ER+n/ydtBTMLBzYdvbCxDfTZLzMDU0qicjQIJ9XTZaVOJHLjB9zJcCosb6EjOgT
HJxJ7E8uTrtPn60UVrqiu8hluXoOzpylc57R57QpSTyFe1TdB13hPSlTZIdivD3m
Gqn27jZFkfyOQnWKRU9cmPfoYzhhJ+LXQsKCiGI1GToif0UTAZovhTOM6/lila6r
3OunRqUTuMJ6d1adOIV/wWjHCyWI6CX7eP3un9waCbCuQLqYkKdP1g1jVe/PXyAw
x45u9F3JWolzT0RN0nJrR06gfI5xrUjJK1gfY646bILaixPeVWnIz9LupsvY29bE
ZeSdao3NabsLUXSEoO9TtiifLG/sOQk2nzCamZtDSzM6cik7JmaRxHLD8nK2s4Kq
1xVPjeC1qkA3PKItcpI5ktDMq8G92jZVYeDMuikyYdCjy+P959Gue/RjBUZG4Bn9
QDWkoXGGrOYfjOO1odyCkKidTt4B7okvXjgdQVFA7WJAT80Elml9Kh1M23Zm37zS
7heokh/DLSBscN2l2pz3PKb0OU9edxH9enZt5+hdNqE481pnYPWQO4LTl72WrRlm
5wwloWSgtZ2MT2FxV1ip1b+YfcN/eDZKiJUK/ZSFhxFMrCXS3ZGGV3MEOwzMgMX9
JSQwUcvDXzvcTfdmDNuhtQpha7OR2wbQKhc6Gi7ZypxkTkX0UI+axThvxY+XkZug
NWxCn4RPccPKesVAX3Ses4tM3a3L7lJtA9ul49p+onewCOK3lMNJErfBd3cTv+WI
nXBHUOYbPk3DA3YtwIHXePxdWDiM7ERqVTNaHywLBSEilv7Qqb1QvxJ9P8/Vb+lc
GGYeyPYwUaFjV02+xQHkfOcTCFU4TKmOI9yw5pkZncVjs7BPZJqYpsxVwac8AsmB
Xnt6t1BAvIYyW7fiGnIqctqpB9MmnghOTp/08FCb8qv+LrRO/1WltRjBD7tuMLXt
Z/7nfUVjXiiA0zI0t4vxUmrAPFaj3y+E7PgMLc8ApBEc7hweTQ8YS5jzB71kfUX8
6/g0lr+kob6otxc72+h58w8XbROsDUbyEe38vsnx+eBIv2DpTFJzbbzrpKTJpof9
tjeVN9DW7xLpSWh78jQCQ9gwTw0fUMMEbwy5WJUtUnMQg7X0IFYAmUUHNX4tP1K+
RfS+5POF8DdmpwHWh2kQkEcsXgJS8jGsJXZF0bICUyBv71xN9AYGEQC0hwNGoQlc
/Bfk/fbIhanG1R4aFfVOUAjK/PjTK6WOg3xCH5ITa9DpyaNEveNtB74sZDevWmN7
GBFCATKvPZy4su5wOJpRlkxIyNz0kepqqzEJwBhiBgQPGcdq8oxPTe/IpvxBy/vP
rfxdTJXwTHTPTyZv7gcoEURkxG7O6SamZ5H5XYdMk2j8CxlOynfFLmf/smGR3Hy0
aE090XagazXtzvwpmmqzbtZ7hQJDK4d4xuouCUXNK0o/2M6h8J3TX1WOX++7tylP
aPc3nNXe/tjnuSLBhFMHMS0GrdiPuMosGJNbDYqbtYJphcr80AZKCuze4LqJtOV8
usjGkhuQTA8Yiw+85lYWXCqAdmE57wcUY0ghI8jGC4nVG+etPFcPKJRJ7YtFioOP
9ilANyRGlNvYluyoIRzLFbBYhOTv1iudFJTgwkf4lzMJBk8QvYwIG1OkI3HezVXV
9Wlt25iYZQPt2HCD/nShVmIAZswXm8whXtMxIBIc9+lPHwXwxfkWEuLbYSlga7x3
whXtqKx91wHFqFSuAI4H7fEU8EhQzsfPpmMIbaK4MOqrq4c2HLV8gcEiHFXdo6Im
JWk6jI6FCE8Ha1Hq7QFjQHoCQTxhbUJT/5azG9hzz1MJ198lSUqnRDeeRTJRnPDS
ZV0YmIU2qsbM6MBTOzXPFH2SQWCb+aNa0oNctMEQJTUSLR1+LvWiwu31jgwYpuOQ
mrXxuTOCtuPjt44iINUf0A+avkp3ujqScJc6vwtKvtrPb9/sjWLEReJzyARzu48x
Amrwfvy3xqr8u9g8qLN1Anj6BTa8l/Rcof7cl8Aln/g6Kgd3/kEDVqcBNZMnemFM
v0+L9io23eE+h7512YhhSTqVHFt+RE4HGonX3FXKdji7AQIkU/b3fHCi+u31cDao
GStXOtj39CZhIcMSVjyOcq4M4V+LMF9CTvFZaLxhXQdxfje6be+K7V5zurYHl37r
TmP+5puIOsF3o+6qIqW8pooDd7+BWQYEG//gid6NA7KeuTLR5WN0eotNQZ5+x0ss
cTdvKHEbUNKfMt+FZdz4Mr+qWdfP+33oMujCzDyIG0Bp4fGmoQstZz15QvTIaX9U
XqRU9PFLck1aPhcWar+yPuEUnuy0ZC/fIcEWt+2HZgH3qlJlSdqhbujjLR0kp8dF
iKHSx2OfzFaMJgjtllrc8QEPAyuaNOq5ZJekrIWuV+2XkYyeGC1WkjQbjPHUJjUC
rEAbBl+YwU33tdSvWh7we8e5OaY1sJSjkF8dGhv5SOABhq18m3l5eneYc/g9FUi8
xKjanMBum0vl/tgO9ubcwTvAS97M9fwSLHc8Kb46OWBpQgXDTEvCjj/KLtLl/qqy
psdmiF8k4ERNsGT0UpaTBywid2rcDUk5OhEudUd2OU+WntywZ9qYV4h6f/WegA/E
ZQ3qGT0UdCNSHcbTOy3/2Mw9He5I6mXaIKn532UwE8p6RFVT7SqmaC2zBAeu5w9h
I3EIJjEt+zLKM3oiKGgGiu/OytV9rorKjB6plEfi0LaIJz0Zt43O6J65Or+7WMBX
iAs02sGXqlUTn/wZkRn3xrq2ENsTKqEuMS9NsqcwdKPYLFndkSxTaTwpixWaLCH5
YVcCNbx00233oIj/HzXwxmV/a/fRBNHVu7afLpVyCAqVeNJeknuX9uENwtFWyPI1
Gq5mf/XO9sPN6E1c156ur9PV/g9dd45DqblcDFOteOtOypN0OG7tGcadLmqDadCe
jB0tjYxTPiDiWM3ZqrfXnMNSiB7ZgC7HLvHn2gIuyUFnznsy+uOwh0qWTsOMVKVs
v1+0kMfVk0ZYXyYNGI7pQeIVdAb+RPnZ4ppD8TbEk1wiZjafAt97aNQ+Y9sj+L1e
vF+OJfKxReUv+G/ekx7OIRz0ci84W+CDIMgOVH9HaK7wtod5klt/MtuOk2cNxtba
EI3zYSE6T2vWDED0BzBCcf/a/QsGZXnbb4CF3NZQj6VcDUy6WfsXj0YuyhLYh8tl
Mj4d1f+AshN1vGfYHE2ZMmrsRVsznRsahi7tdkojqWb67eSsCaarFGZa6J3bX8ux
BIacOsZnwzmNBD2F9D3I/fSZj2o2dxLsFI5CVn8JtKIsohFT0kEJ6PALQWaBOibk
2SlS7JepomDC3WWvOn+47+LRLJc9WR9s/G5ZVypgDNWupXHogndOate0X9AR4X4O
o6ah/7nnM249Fu9PLo7KHFx8hYSKIyW39xzlRNkwj8xSYMU0P//ex6edzyy5UCoU
iRlP0MhIJCGd9tt+Qh2a8bKiTfYgvV47v1k06EbHFpEcmmVYymrsQVz+AM0O3G7n
Adyh8MK71e6ESAv4bTW+1ZlgmWz+WitSAfZntM02y/t3fPW6UPSIl90W63kiMl2v
oPuBcQYSOwA3eNG8XezUYtUEbymKogXqr3MAYr2HsiNe6hq5aE0+0kzFgN/N4OmX
hkdP4t7gLm3ZDbNq8atAYHVGTuuLX838iwH9/kJuunCnLZNYER2CYlSIAQtavv10
UW7dloOGCs6jN/93GbmpXbza+c+SQXivAILqfcB7VsoPwVE+W1jeIpEuvztKTe1z
ZlzlZNSLyU5kb9GRVETK4XVPqB4TZ7ob50SjDttg9zIsmbKQaODm1zmpj44BrMcc
nuF65/JxvYjdT3WbepYt6qIR/umVj3yqg+8hO2SJiK/cVEqAax8wBV4itvujjZmx
lwj/lcg21sVfjWdzDwrHlmPNgz3b2x43Wm06gwMrxHmCTrF4ak53GAJA1FrvaWC+
/nPNBFrLE2anmLhMxvkx5dAb/xaYrP0zHlLywcoH4aD1Q4Ob2RGf/U33aBGDJOCG
hCXcGe7JGCFt6ua0fkLSvEorv1nMw5RlwfEpQlmFwhI2Yh2KBb504HRfYzx6v8fz
aJm5F3n69uAUaynLU2OpSlmzj5K3NAl5Sca5MgEDhN8uV3mqUD6jVPdLBaD2OYEj
nZS7NUEaIfhURRtdYFDjV0wT2hMnVmqzd5uFaaRuHt7jLhIvQngKwCm2FHWtDB9E
kLCy5QuXozjU1HM5pR4PYFb7FzE4CjpqNOaeBjH/ur5wGvs8pw11/k2rjyGlZwzT
FNOARv6SQK2YpFbsFgFRx6OaK+L3p/ZSJQHhpZ0KWPctXAVLOB9MlWQIVESauE7z
sX250Q1mQQWuMqb/wn1nLhurDbu7s25te+WAgiTorpaGgU6HCE0D/CS8xSssqYEh
tPTRxpEmEN2nPy0ID4Rxtq8VledyqnLLEnFOccW9C9/10KYCjZee6j5X+dym9xgT
8xAr0y6/W8qcM46ddk8ZzYWVg3zFVS6b02kIZaLnvQMIgVSp9usT+I5RaIeK28Z1
Ll0NVkYowzj5FE7caWm/+BMwsIkeKRxNKL4Q9G9yyNqemTOUBzgbBTGJNETzu9RK
77dmAgcf3PMf5ZzNXjrdrMczNS849xbygmy95mOvf3AxZozCrJmiVLFP3egIWXID
DYz3Up9nNUIvF0QGo1Rk5s+cfthr7MB0jeEBwaSfbIqk69Yp913aoWZtzbZ3Q/iV
Wkd6aONDECx08qhiOsw4rWZRhFw8p7CUbaISwYTni4VTS13DeR5jzG0zHdKoW8sy
HKITXoKBit4Zt15XdgdQe1+EfVBxiSMdFSK7zXDIWqNEheAgJCWV5wZ3MILePIeP
OAKi2Ep1ialQrilrPuyc/YTJDRnXisFhJB8kcWSCBLlqzMhAnT5Wxkti+VPfSWeZ
898qG7nA4pyFZl4BblVv5Y2iFJl0MJk0FckoYuMrhGW7wHOA91C06SdzUH/ieOmh
Q/owxhx2yUDzzEe/b+etJHa0XW6/vtmje0mILexxFEpH4Ux3q+JheoxvhYrPC9J5
Z04xeEjXm4esm3TPDiZFA5Fz+AqAY+2sFyGOTGUINTzV9BgW5gZSd+4B3h4BDGCJ
HMwApVgZIJppI1OQIlSxVZqzZlOOaCzY2wMZkBImG53DwfAVD+omFyQShT7pKECd
+spvVU+yp9PusK54zkqCgIEtHyAW5STSG8oIF6VFMV90iXlT7xapVZcL4jwU32QP
f0dKtWtS2HX+pBGQ4RidsTAvHfoiWor7sZq5djRoO1nDZaw/g4l2/etITqMepENK
gPuHlCS2MxkZp/+08OJRtLwHmKPcf6CPCutB5jim+26mXh7MzDiPYcOKY/VInj1C
Gaub/v3c/o1SNrXH6b4duDT7q5bL8p//dTtUPWEy7q9REkB65rXQ4w10f9J366mW
lQcNg2VWVH0Jmi9NgNxW2XTEOtbVMLK6LFQ35+MoP+pqX13qqoYHfvQ0jgQpWdXJ
wewLpflKqcQxYdxIqpZSWcd4s5OKpI3OglHf+hH9JoF0s6srasVPHwoYcb4d5Bpr
hZHvOlkHESlsYZVno5PxXkkV3Da+zdl866AJ9enbxPRuI4B1nuL9BlPMAIh/yLDr
D+9CtUBlUx0HgXjq78kWRiz7b1wDhnUjRTQDzf9afiboB5Bj4KdtpiQwjLkHJW9m
4UfpympBB6PUYHKqoyTdTTSOfPnxHkjtu3QHb83dWUCLyaBm/RhRkAKr0RaInSKs
vf3aRqSEGVctQKWJ8eGHAdaEoRKg2V4+UmuodU0oHFzhMkPw2eIjxzpyzl42YeOm
Ptt163b86hU77vcv+GO9coBA4kLWofmWCWkmicO/128HJOfq/k07tarHZlYqf9V7
Ro1rdoLTtFA3Vg66P1DEMwsjUk8xXaYsAUcKEXfM4aLYurFMziizZClsrrKbQwrx
Mdv/QPKSAXxlhwC+VL4kAlQG0Avuadd6S1+s6NAYQnasbitFNpAetLlLDCJtfbwW
GvjoE64Wu3ege6tQzWSBmvQ0GHNXaG44TlfAIcWZswBPtt5+FBXD6RjW+QQL9H0y
sIypzpPdrhZEiCzW81X781i320XiscxiTbU+uzI9w+knv9CX0IeQ3ixEmqbh79CG
7jOTzjGpAQpJhndtP1hjw1KI8wslISl5+9M3elCWUJKxNhff4Yj9wH899/bKe0Sz
zkAklEBaPvenV7XnkSjHN2Lbs5M32DuEAWNE6WgzY31KT9GthwMh5ef++xLQoyGU
GjG3wH+NJaAf5FITaHMOMb3ysUnO7LSsyVdP3Ax24OTbI4bz2yg5arKR59chr/Pm
pIVoygItXX7mVbZjOCvAe6Id97hge3QziWI7SaeesujkSV9fVtAwFnRIqoIzOVsc
Vx/lbEEfYXxqyZb+bcWelKgnCmvN7zXD4I3xE+bT/se2m4N+L5hnFEqD1Mfg/W2/
Zj0iGxB1+q3zw7I1wPnLAzvDsQWWaHRIRVDlBFbWJOkA77M8NM7964GTqUloyQSS
W171eOhml5xETgad3JsG6YqAPKRD0noNEluzgQztL0IlqsS50w3DAs72vNb/HR+4
0Rs5YfZ5WxCbxtQDqJ3GN5OgWnNEXmLRDPbTk/p7nZAsPYxFeIofKobHH+2PP2zN
CNgtUVg7Xh2+UBpfTmH2n+wNwmi8t6KNfNU57drE41IFsd4Et6tDB1u2ab0zUvYs
Ah8fNY/reTnt3Z9VWfd/T26oCecWXOoRXST9UrqWzBUyLbUsyqY2MMwPM/6zsCiO
Pt+EE5a5sxOforsHyTKKm4bYJhYQGKl+UpvDeOKVQUbBujWVjiwSUOimoY6lE9VR
myLEsR/ChRgLmzcYLf9H9IXNwa6viWiaveaS4MKzJ1po2BIv6cvu6rGBsp+TWY5C
XCdn1G5bBlhkZmCBGA0a2b5ckaYKnIKYyYgVx61UbniLDcrfSHoNAobEifK+Wye+
RnG1OdZ/dQKt8ezf0t8hUHVdPUV0XfE4MIbz2UvYwRnEtpO9IsQ52UjMWU+8Uv3G
LRXEW0GuG83g3yBePIRMf97O6tVOkg7lNxEWDlbIxG/VeS2vfeL/liWopgKXNrz9
RuLhOokoUHtJQ85bcCXxag317TTsi0lTcNLCEQEAKUoLHAUG9Cj9rFVp5na/ndYn
2W584y+dNmQKMNLftc1lMYDtlE575xqZMJiRHaI5J6M3kDmZv/KdBq7xTv6A88L3
c+OAF3XQZaxDA7GBRjAjswFdMOJ8N2F7ZXH/H2sTy4ulTKgKDr4mNQP1sGjs7N9J
WcyY8I68HpFwGRUAvSRNKd5jkgZ763Bdr1ShBp1GIWOHuOObylUxcd0KWblht63Q
Rqv46I7XAh9/dd0ojo/z/68maAOq172AceQSouldjIOQS09m3iAWbjyvXa6GLdwH
RrK+wLcnVWfcbRE/FF5nZ9y+2VXr19t4aMHLMrnzYSqKwu51QlhDMuXr7HNOMK/O
iOhDaOlNKSBhhabcfQtTQqh5xaCnUg434AAj3Tj5ZKCRtAtWRV/BHNj2TD/pSO0q
a9rZtdC61Em73O9uFx5rMx/9xmYJvzE0lsNQDq2aN1AJa51mAC8HdTylibirEVsA
dpIOQZzPx30Gwktfufldxw8xHJEqAUcYUITgo1uJ2932u0ZtIaFDGPrtiwnEwkl6
YUGtcVubqt6m08dge5cIupJ4Cc7w6+gjrCSFQk6yggrU8gZ44rAHPerQ1sgd0P0C
jVuCIOG+7dAZMrUwwq914xedBiUQJN2qGMLulAAVdbQbTczXqJn/6fuqwawnlS2a
bQpCxTgn1CPB0DXFpivDO9U5ngb/YEEU6With2ALqm3cPWGQ4rAMvUXkGkGU/sJH
7kaSe2HXPw/kNubNd+VBomGXZaOnQ8OhOfrKrl9pMis1CmmTF3PsNWYIIadghpy0
7jyqzDkZ22/flvVV4P+sw/oo0Lco0PQXk/3oAIvHNTHyaFQs3SH9/mAiJ6+zgyRo
gKR7rw/tOPAF3ipQ1tHfpk42vVTZ+ocE5qU9TQL/Oa22uYuPFnM46lpW5GYB6cfg
15UkT3c3fJqs2T1bY89zNkrXcACrRhPom3f4uOmLqDLfn3fIfNIrxLlE04UlVatw
Jdq0FeLgrUp72G+6bWkly7aO+GY6VbbJgRY+r9nppWn+ehe+0Ec/DVIsVCcbKb2X
hJqW+KYsVCf8XQ+lwBmkXW4k0F0awI5RhHLV0zhhfbZopuDh9EP5OaTg4UY9Fh1/
j6UwhM8VZ32ddM4JXhpqhO0t+6oDvVcGruotSiykG9aU6v+LjrERAe9LlUQDZRZu
T2tVxYH2BToqeftRioZTR9ZDMg+CrvClPFUS2eISepxKNuyUKAM7JQwG6pYOdn5f
ZCT9mVkoPQTyBRVoEK8yle8WrhaWeGivp+eFl9MzhSqM0jUHb580XggqxTZkIZ0f
gQ2TdSv1UTuJSmZKSwAUWlnFNwcqOQRh+5UlCmfXxQfZkPn/JNm/xVie5eCFBhuy
mb3RaLtXTMsx5ZaDNeZJ67CME7M4rNGbhznhY+KLyZrm1l/XAR2r6Gaxz+N+zb1B
GVGQ2chCYhrXqbneLx8U1Qe+CoGyFlG0+9bs4xLNY7UODt5CRXofTErtpW5jxYgh
059IrQ9Ra1Gx7Bi3gwcETafWdgQGr3ofsgwleAQ3XGRRi+x3c1H7aXdriwSeC5bZ
wcFHlq2upsJIfSLEaU0WcsFJcxQn4sRt9PDv53fbRGOr5H+XPHKjoWRMBzb7ZlAN
o0+QLT/63W9Yd9cL55OZNIk1TCzC2KpV5P+5ZS1jY4UX+gPczug04Nz1SEZx2h33
5cwc16WK/+oeUZQfibLET/qFD8XKkdP4nlmKePZKnALweIJFB6dF4jNl1hhxQkqk
1LPTPmhOwCnF3x4iDRWpqibszOHHs8Sm/0jrQd9eGmHpN0wNGtGtICRk4ugrqE2u
TZ5/LR4vkMgo3NyA1lZZjNgLPrYjfNtkx3+2B+FCao7qc8U+nbSbc2LinG6SelWH
A7oWum++laJk4NITRcPzDkF+ohQ7S+Odzc35EtvxrZ2QMraeRGQi+mKRzh1r0To9
3nz+2AgY9eBOPhvcGDqIQt26bzpsSnTI7deLkHuAomo3Qcai/6aUsgz4HwN+Vd7o
RRhi4KwlQNxN6CxZeGfLN45YVBTTwjhh8Rw9HcIPRJVbEc7hZ3bsr2hqMK/JI7Ui
margSzwaSVbKkSTgcaWqrrALdUyEC+Cy6b9cP4YwWk6dye7QCMHw3UtzwwZYohuc
LA4W8q+1eCPVNPjiSKPizFUEZDOSMZQy1FsQNQ72bP2Hs/9NK4r4NCK3bstDS4Kt
7orwkL8LZSMnS/5GAF/y0B1qZcCExRwhz53bgRVZSo/f0e0rhjdyFz+Pevnmci+X
ZDEjKAVu52/BEXUcLm+2ElIw7O1uPLH31eVlQnNG8r2bI7A5s9JzaKMbxK04NubR
qfw/c4kXo1XJRX0JoWcB0n+0WSkD1H4HR8Go1V/pmu6cLH6ib2mcldp74lIre2oX
vOVzyC61AQrWrYdYC9nfEqRQOrtrVXkrCAsQMa0z1kqFIPA0jG05REVtCqg6DaEW
I4HEEFqDF386KBJMlzKiC5rQ6BDY37rrRvJAZJsbjW2zGwP6zvriRcIY38QutMPO
xOyyzy/Wcu7476omjBeWe00mc8Vu1L3WiJK7axY5h6D03hmTT9PXOIhp4J+25Jsy
jHHWRwfFdYvTqvi28kOUG02VxDn/iYJvktNIWn9/0PcdUpT1dPQn6gkWTqe+7bFX
KiMu5WTULDAnqoxUo++MuaNnBs0pkfWAmyIIWOrdtNFVSb2qZZKLTKuhMZd0pbmu
0j3Jtlkfj1ysPcHR58vpV0DqIFrbmO4ZGmnb1q5VbSIp9jfsMmvuILUhPDHbdtEv
ewbgFiU0C8jIh8WReDTT7QND6kZbtEZsCT9b7tLErwWR1PqbT5UmWaE0CuudonLE
fm6OW8D1EFHOvuQKTxpqBHllUWz/nlDcTg2/EOYkbVu2woV0sysr43RF62r6v2WX
J5I7ZIeENwN6z9WgOzRPIvbfnpnt6rnNNnwCF+8SS9xGlB5o7qH2X1NP2/+Uy5W9
c+30SM4akf8LOeFS+S0NrYLs9BEmotc5uEDQ+hnSBuuHRKwzQDEz2Mr1jX6OFvWw
Xb9VqHt/oeRi8brqLT743RfVH0fiylU3/FIqULiGWAYTBpwxJMLLLFWQd3qHppBp
ciV0UUDmU+AlKVlDBk2ceiRa1OGhnYWS1nrxTRP2nBrUSK/ZazPwBHjeHvpty5Nl
Z3voreqP8YmsxzCPUEugnv964UVGqO1EDnAbnuB+eb4G34VBtoFlwSrlVdC4lzMo
T20RsURD7kWFjQ009BZKw2p4jzVeL5Cd9wPNu8FDpZzYTjFOdVcB6divXMwS/kox
kEgduxC6EB+eYvc/40kRIAhddCRo2xVgkzu7uagcCWiHRtRCxhWh/Hmc3GR8ZIhI
FA842363jxl6UfeitnSQHpz8CrlAqToiRNgK+qPAZi+2RPVSe7NHigZo7qm97Fc3
64a4jQ+CgSnFjns+zSicUMvEsil/1aghfG/n9DNb5S8l5w8vxu0EkPsnt35mGbaV
9FAIQ3mPTdfMd1wGV4KsqySIjF0k1xKQEuX9OPg2U235KFeCnykgfkSeGS6QrG03
REMVrWsfljFjMb9xV8juRU2zwShRCnlxjduO+B7UpDaU6+XeOLOupRumRDEdZDcy
UVA9t8dA2NJrg6EdHdASzqFu/HckYjudlN6eO8bHmO/T4gYGfmMBIONe9hUEVdkc
888BWDGkf1smiEuJu5umqCgfwWgc8Qe0Hh7ji8s0KmklLNjwA+uUgl5wOdyy3E8q
uARwWcpgFi5P0wAv0cn9NpRezPAjX/vdN5uBC/VdaaIeq/2iPo8vDhtRtgHRdLiE
rC781glhE6m5GrHELp/pMolzGrVTnHnIm0v7Z9+m/h1jU6h8gb52V29pDrHc+1wf
usKciFT+kZVUQA4UttLoVQSSLOFwjKMaChXSXNx3QjeZuy83zuOJVVfeQVTkvV6Z
CZxOdlQQi+hkgUuC/g2jF3AZfY1dZ46Oc0nC0CnboCCWwlor189Vzu3SuKtQd9y0
yQijM6/PUWAXe0XlK4neGv46gFiDoQf28GHzEnlRDq5RZwW7rUtwjya5QDJZSoy/
IR5wGG9wChyTj6GwzpK1iie0VLtk6JKpzxPDAZ40bV47VYouYfrKsiWoav1MfZMK
4s86Za74BrIeG6EHji4ZuT0nw69M+KJDL//oGr0FwEEQ4wdKwGR36146tV3+SiyX
TUu1eJEtFLcV6EsU0IPXs9PmJ//QpkgyMQko7Opp9ZeIoeyxD3oxns2NBafHshpV
OttCjNsgTR+EBfsEJErLmw/I0qppqeAMNluoyptCYaW3SG0MNCf8sTz6nzv4aYSj
G79/TAC9qkCMqRO5mXjf3NO390NIf/kSfHGPeMY8nVObDrVUGLf0TwsuP500n19J
AYuuNuUEV0/SNEhaLiAPVPSs0CmiwUgfnzQCWA1rCr0rsRrqfkNyQFxWlcZ8kvoo
Coz+Rc4xE9CDA2MG5oOwJdV4J26AqB5+p2SPK7l9GxIGmLkas1Zjdup9DPNuPYd9
95pwpUuCfQKBcyFqpehI3P1Y34SR+7i3y/Ci85nY4aCpT6R/pHshh7tMvgbk0bLD
LBFfcskQAsejYe9ySXJQX0mDfw2xJ6GXGck4OLLGy6v7xsS94GviYeCQL/PkAd1L
jx7mJNTiVPhSZ+pjzjLuHXyMYjvoXxIcqiMHwArV9mkNCdWGlccCDqauhwJD1Sx7
oqaIOboJWwZutFrd/sWtvy3tqC1uPy+G2qmXNQ3Svlr8EMvuasPqE6phcQ+knA7D
jaxrqmP6d9mWjFLoEfhhjugkq8KUbNTvnqE6obMgJ4xodDcX34viSxr3mHA2bY9w
+T562ZpeXJBlJln++IiuEtjss6XlY9+mo9HW+o9mLeNVKcq/v3JqBJGFCfXGNMOB
JRRBDntJivmdMAM6LOoSWMFVCo4bIyx01MYCiBmrtVWqYT8UJ7yCa1mSCtxzeUTx
ALK7OrfQUxOMRw6TMz4IN6j83ZtT51zT2a+AWJqAOjWfGJJ934IrOmvnau647dhi
4EIMUAxHyVVA0RNJ97Xq29JeKJ8d5whMPU4n1IPJzUCqx9syxa4E1ZfRQRL9E1h6
eg74N/nGmfBU/3xUfFLjiqsqutRg33P6DQzr2R7eZwbxsXFSz02ZyyAp+k8UTpLN
AR1XIl3GhUnbubRdJaae215i5SFCG881xJ0KwYQaCCD/INP5Ec2GW5DGX+ifYvK/
gOHimJySQEG2lnaFup/r8KgW4+V1FpOdbeiODNoNyIui9c4rEBPXn0J1fnOmJgZp
ZStNRfIGnJ59SWAwXcHw7iqBHgc9DD5sBoPNJ++qDQjh0lRs1pSljCQrDk6MY3du
nspPbZ6N2iN8JmINGr53Kzu3oMR3oPs4Q52Vfz1yF+0Jk9ba+gJwgxvJDfyHtrRE
Czt+GJWwr2PSkB8hdbcogFOjXtouflKzLlZTwF3a1PX6ofiBFm67qSb06liwPLEa
3SkECvC8Q8Ng4BjpjokRQeG7+Jg1Xr+G+O//ACMrwvTkFBGD13Ok6jjBcXTpms5m
yV9LYkHlRd5TCwYL4heAxjc34SHll56AWK8/emfjPp1i6JwyOh1m6LQ6hRT2I/xe
psIEqbt0lvKWl9V0T9FNjOI71ZcnjcF5fNyU5GvDuPrsRlxXLizOtrtT2GnHdVO8
lpjLXo5uQiJk84fbxWlDuEJEqju3wOvn8fYaHulfZhXYQRVOD+7STZbEKJiidjtt
dSWP+HNpTN00wIWMgUbDG9Z3VjpCXp8cZC4YD2x1h7G279zKJO/5fW+/jVax5vES
8HXbSgLHUv8PHxIFoa0mD4cY/g/zkfcbT7M4nIN+ElkAbP4cXbEqEHPmXD/chkTj
eW8qvN0+zKR6xFFgVQOH1SDUhZWEniRizaNis2w873rb/ILkAV54Autpz6Jq/jVW
mHEXaq7qSjDKic62h9v2UJeGHwZt0Lq7VPDDvWRPJLdHYIHM90AtoJctdPSPCv7a
3uJth/0mEw3vVznKUiEiPDccFQhXIauCMsOusQvbnoKwoNdwfS3ZOF8Em4dSTyLN
KgJadswLVOK3ole3N6yo1CQ5EPdax8Ic0XW6AFxuaVDDz4xAwT0GT3LLVFp0pMiW
gMYZtN5KL2X+40XLizc127ivLlBCuOdRawMTRMuOUq/ACAQgfzhL6vRHJhousPwu
gIdZKS5q16iervft7PEedpKOH3hjUt4Tc8+AUGMc96aHEHfPnU0JAZWZG4h6B7jO
zrM1Eo0hJ4SHMMYHv+5DBAnAKXsx9zVYCyCrbCsZ/Rj44b7W0PW6MQaJrdS58evs
oi5MZZFW9/x7EqRPzarVgml6LSSjg02bPsys9vNxmuG53t1uRMrLGXDMmt8KslKK
cDYSncHBkGR+tLJe+zIsA3JAExzdu8pqaBRaeG2kz40LJ8+gIxJx5X/CPbmjL4+I
SvnjLr4V4kVDnguNdasA3eVXyR8NUxWnnii7BuMqGCBEYXUbZd0I5XfOMXw+MZ9k
cWo1erezy7p00SR58KWI6p0nNwB7Z2RZRJJ0hIlRY/UQunUhUcH1pDHZ3ZCivM8k
HXviuEZNrSkmZJBNqwe68uiK1WgVSkyy4m5H0MAMhEt3GctIiC2B443SZbw//rH4
XLrg6pMrDmddPVtAX0blLGQ3K/8mGrK3byFuMBo9XCDMZhQUtnULGmFKZ40O8uE5
QS5euEnjnmVpeCABx81AGvgSi0PdC63KlMYRj+RBNv2ypuRjHCh+uZu7r2TaCYne
f+u0MPywbAhxd4cWAUoRum5PU8tRXStNXDuutKBQ/wpHkGiGnUWffE5rSyBlXIx8
fvuqz4BszW/D43Q4vMhc99jbxUxD/SyoJAFMLk5jP+Z8w8YBX4Ltpi0GxlXiLCn7
lSK1w0RernZm+gPkLfOCgNkKVc2wRKAMVfnHowEqtuRJc5CFH5c0u3p8O+IaPCDi
mb9Y+ZoXmnXFiVxvYdCoQOiQTlqvXFlWrsMVBQZvo5fiEMRG0G0ZDwueV+BXalto
KG0F8ENrf3vG1+wRJFNzhuDFUFFC4XAklq83gFgNT48EFz7BdgSmhh/mHLqyRr2s
zIhSiszGxeHoh623Lu0J43V9FWMRyjxpphA/2jZLxwQBi+AxULfg33Lm/jyVNLCi
NUAw4+YhxEUBSFYm7lRR1dQ6jXQfNLAEV+IEkRKg0GAsxkFLPdJIz1o8t8+YWnPe
wP5GLxcfBOppAxBg1Rq1Sf/1eJczXfleSCwGaxs+2D/Zwx/BXthrSlyYOezeknur
x+7aLFs7hw4uqukHJAPJaiHF4vJmsFZgiHqeycDcwo87q/L3U5bBg+2bN0NsyL6X
3wYlcWvSwJAM5p2x/dRVYF7JqBSRGpGMtXLBNA8nQ/cJnk6LN8qq9c1fXLb2QKeo
VlIMSRGz46TQPQDzlvz7YITtfKpovV5p6sQhCz6CxnH/h/q+finKWH3M0H+cJUZ9
s4bUJGdLdJlJQdMmooHEMM0WSQH5UL9EbvNDV7FaBD64P9ka0aNP40uwOjGJGCsw
+hUXeo2XMAYNJDY2NGNaZLiQhgm8NMTBQuqpNyEzCmi1C6X5DsMedcQiKoqkfvTY
ofOFFmd0YjpaQkxmUK3rO4gOnGBrkVqFzuRhLakzdVCGwL0gCpf/svxj/4y/yExo
RCGylx0ptFtrYU27pZd3dFMVU3xvqLuv1fwY7obovPQP5Jk2HfiF0ERJoHQOPY2i
yTA/jqX5k/KKgyeWykU9oxFsBMvXM0idEz8ootapvUg25+urfVmdprzBuksdIKAn
tof289qymHW24m6Tgv+fY65S4kB/Sei0jFAs7LxpkYNQITE518ofpgJQ40fbIR/i
e7C/3C0zU9VVL7XjVIOcdf1QldwL2dKr+vEMGcJBcB6vEVLqWbO79fSo0nmO2kJd
tf9JZBRUltMcqjBqjMEe7QLp6rgfBJr1Qjp2335dZABPVlSHA9JTTlqHDtvz+37X
jCeb8mC7V6820xhAmjuyedW6HYDgBb0hXr480yso5CpOxeL/IelVAXXDP0X5t2PW
k9ChG+mJtJeu3+rL1OVxq05XzMg5HG7iwkKeD/KUGWoA0JjEPhqru+6J/oUEba91
AFURsiyS+Jkce7FHRlnyVVOK5TH2cXnG2PqB2eP5UdKbmDfI6b8kkp6wT7NofhfQ
XH22CgYNUGdHbcv6A8pcH6BwiU18FAG3IeWd6gxR2Voj/pP0xjI3xBrwTjEVoS9H
lHDmjfuFjjUTgCV2Iamf1UedS/X7W8xComgyA4GttNm7m1igDtInBtXZArGMYnix
vxjVLHbx2VkG2kaHCAyJtuGTjhmocCXSMj/QvsVcbsRx8NnoZjVBahQ8tc/8u250
aa8subz+vYInm9Ro13eTHU4z2xDAQWZgLqH0vw1mMawTLym3EGb7EyMz/ZseUoyL
WZ0+QrUVNCNiBQ7eJX5MYkmOWU22MybdxFHw7KUliZeQ5c0MYbjl7H3n/0DcyDwA
LrTeZsVA0wSmS1xbXoUeweDhg5uMLDLuo0hByV53r8pLRa/O/lm5sTxVDfMy0pXC
BnbUaJGhL6WDJaZQV6diOeyMVfPgglUPXsXjJYWZAM3izAkThK+1xQLsMzvdRWVO
r6rtLBXFPom32NDliN6ty5ac5j7pPHDvmunWSPvLr1V/2QJUejjslIB2+DuUj4ng
TmZz2fsT/5VJm4vVlN+mh74hlY5D+ZKbG7sEwYQsIu1zZ0TbWgvJvRtXR9Eunb/p
47aA+kBrXkISkyVfiDY/Zz96eIgkl+KOqL2KYuycM3E+25DvkG4T5wLDNzHKwLTJ
jpjqYBbcHLwLqA3ELtt0n9X+vAvPFVXaretyrjZuBml0uOz9bdy1uSw8CLVrMf3B
DTaOpzjW/8AmUx7LaEyQyeqMjIN5wGYNl7/lAnTqgUaFBCdJIAlw8OBjLUDHveSX
nO7KB6wcT9IsToZBNdNyb4JS8f+4ZSYAuBVSl5fOzWg3Xf+C45GwlzwDUXZUjNSH
tX7HdW0Z31l6T9Om+On31pYVqU86yKy+ltm72aPNsYSEZxs6rnrM0HaOnDG0biST
P3SRmCaNFai1PCBJW4AZnnb7TZtz2Hrr6gJhQyyWzjOWwYnIBE4bZjG5RfQ3xtsq
`pragma protect end_protected
