// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gTx50s2NdesJxI70wVeADelVKouEuAojUsvuU4hhEKiHGlGFqgNTMZZq9Y+BpBTA
Db/+DjXLFiLM/5AJ8yZu/fvtQB9Vb8UnI3I15elk5VI2RWulIv6KaYL6ReObiKnD
8RVYjLsdXzjWNt/k3REVyA96UhjACud5MPbqYpBmjm8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
+UPx9/wx1alJV1JaNggiu5ogmYyZ+2Ok7cMLdssMWGGFclnv7stcRuQwjzvOmAzF
9daBzhbZ2L0otbZd1v13h9goJ/I31vcaMdHIL/H1g4en2OBc6V/Ai1vH4IeuhOML
OSL34Xg4Cok9iCqNn6S4Sqx3zry3845niNh1t/oRgIPMIpEiSkf2eRw84VKDO+cY
uiWIJToL89VL6GPcJcUmfP5brT1narprN6oveiZ3QbafvU+NnE1yGrQNkc34kLpq
kQXftdFi1wMCrTELvvyCapA+RcZLiHi+jWb54ft+u42nYovYfXTy+QYnruN45x7t
CV8mJSSAGeJZeIRvZud+mZQ2uvGXNwdrCBcu/SLbAn5G1Clk70qLU9oS8CcVo5y6
efbobiRih3PPX7xFOPI5xdBS1ID2sIt/+PldNV4fOJoHo5Qi1wUGVFms7ynBh5+9
g901Hl86fXlieRuS6+VYyITG8P1G3tcJSQiTpX4Hcmowft/JXvzQ4As/hEuCr6DN
UWEyB3M4Bm1G3Hm5a6QEFgjBSDLBSCF1O9AOcQOxwEmwSWHNgCKBCRTIWGA5hcew
a5XJDWdm1mmJo7fok0noolQ4zDOf6j114Z/2KwPfUlqJHAHy6zMQu6wkoVMc6W+R
l2wWgNgGH8RLvORGhOH5uL/xXZAJVmJnGGTqMg6f5oAG1WG+7oUhj7mjKDxbHIOw
2mODks/EH8XS1pwVv+/84Mk7jW/MpXhybYFyhVy9BmUv7niofxj9Q1tDapXJItWz
zmAvm798ALn3jl1u5b6Wp0C6IqZmElG3V1oldokPRZk7ZduXC9O+Te5LvrUpd8yS
+3n70yOdxhoql4EPk7nO39ZZU7rmiw0OkUeTYh3jQO6I/LbWGOwci8J9dB5wLT2B
kjFWQDDLcSHTeKLZiJdzrRycycC+aex+zJcc35pB3+iVRjNtML1QiDeggrvmax3c
10iHXpJBeHfd+3UaU0TCLDUJJIJsgkAr707eaD6Xrb/tmvS3kcH7rA8UDUdRKbMz
v9+5Jnl+VQwDSQKln5WOzjbAB4L4kSfyM8rEu+yd7wcZbqJnjga+1Tw6mKplHCJH
H4mnIlEnkIq4pMEqsEwlDaee5I1zQN2EPGIOsLXyoKWL+FL53M1e4o2LzVDbJ5/W
BIV8de5jshYXXaE/weS8RjMm6rIrFhN1SvgMYRk5ahsJudx6DZZ1+VDrRxaerJt4
Vu6Lfs9EW+xFalf0CFasfMcojpk8iriwsSVcRH87XLFG2/3aW4jCnqaZ1Tz2AajG
KP0pER+GI7mqJ9on11s5TibSZykmhSJyfD8rgiPFIefLtmuSQIjZmHoR9La/fKpk
XJB9IF0JKadJqRuH4P91KNBuVWvgR0MgiIdfSYVm7rLC86r60RN7qRJsH5QsTdFD
n6bZVtTTHCsckBD2ieke4rntCapblL5QF4vS0pSNJ7Ll44OFgAU+0yD92ehpzMHi
xZvmn0AkyOaVzbtfaAO7h5iOzApz3L8w6Iewez0F4nYBnvWKdS/oOV1Mj27d6zJr
OTBc0KCOBKOoytInMd1ICuhpILDogoqwIqZInJ70+EzwLZbAe+owhuJ+12RHiN4l
ui+x+dVNBN6b6JztLyUDh1eVbGwl56r9VsSzkpczB3immEGovT8xdFPC91GRLMk0
fsNEmqSBBYR7aWjXGflBVOnZLGx4ZyZfsvTrmzsEfk5SqHwQ/d4dya1SXpqXCUr+
YCiMVg6CE8VhXHM40yhGST8HxDn8x09pq1jWrtAEuYx8UcJIzrrIR67Tx5C7EwsL
7EeFzlSGNXuwvgXHnoKIPfS0BovKEEESBysCERz5dec9uOvr0jt5oT1VxVReijwP
VefqRdzJX842P68epZX6PJH7DmW8JhOPa5M/QFOqEtJUUo4WTMRerpsip6/KO4Da
d2qwK8fwNPv96W42WLgJQGwBK05Ba2s+OVRLnkA91HlyRlvNQzmVlMeVUK7/tlA3
WTHzih4ai8kCdg+CqFCtRZi00kvspuaMgw3TBeaBWxY2KprwnS9RlNLACxO1CvEK
iTL6TGtGHBgqnamzolvLWBj0JPIk6EWkdQUO3zzf3qEKPIXpYG8cuuc93mDPw+mJ
1GYxAfb6XZGE349G5K2GnlAJRAxBHWsjUQSs37iRqC8tUXFmPYFRpZ5kOBpt801i
FD+waIThggNefE/dT2lxg//QxiAVfKqKuqq5FyrAS7HtyvbZByr/JebiWa2pgk5x
Dl5w7feUUGZWyMeLLdX3sfPAbj+hC9jY0nzGLmRzNWAggPb8oCY5wC0Ecly4ArgG
+beCskoVNW102k9wkLdU7OxcAnI62AqskFNuTKC2kldlqUtnTEGc/MieRGWG2s7y
PfVS8YErM0VrR6+8nndW5UsG2oJNB6OZLgTBMN7gJtn+5F5GSAwey50rNlptCkeP
BvMIRRrCweu9Ek0sGWfmug2/9TevbQvAXr4v3RzvZxNhBxfLjI4fHYpMKL6jKZqt
aNbciJpCpYIKS8eeX2SFY9JwZSAOHMp7LVIg7NZQLk5hBDEVDJ0T2YRZg3i3PhdW
DxmGjIorMk0JjQ2Y2YxWQ5xfYNNuGYxWi/A0tMpVGfGp5crhSidl59D+Ay2XtiGH
7Bsvd2bz8uQmyjG1vhbG9OmKfqZ/Poeg0P6aRN6JiLpwk+cNA30aK4zLWrZ/5cNV
CIlkXPKzkpOOWvo+rb9XHKMaL1PYyrYvpIeVtTm+l+eM9kE8Bu//1PAjUrEaHX6R
ICTacglA0pgyM8MtzR5oRx1Krx6hbfcpt/pG+yFOvw8Vro8fT8H7smWZzWkT2Qyf
VchNW3J0ryu5x1SBlDb2vf4fPGZ5Ymr+srAsDZfd/v9GddgtoXtgtBPODNJ4/rIq
1v/QhJtXna6LKDvaXWtj/Fouf058X5PLMbS8Rjyhm3+0+jp0N7s30fPyzK6yrFoT
b0npxgSrO65KWtP9BhzM1cw11WwG29nzzmwYp1KL8PlSqwFgJdzc0FcveWMwfd95
7RP+Tt64Nl9tkD4lgbbPaorPLcUdi3kV+EL/f/LXvyvPZSsc6iXDHe2C1q5AWwXz
2Uz2JWA2kigtz73mNcrvwy29V4DYTjJFEkzoPijW2yLFNbzxaFSfBgFK9fPJqa0Z
709TBQEkER4ZSdth0D9Db/pWlJTECc0biY8NckfCEwqCVPL2bfyhNBdnc0spW7yE
orVIsbvqrBML2Xt5b/nWkKlyEK9sIkTi7Ac4Ofe/VGKsbfTnLpRCrZ2iiE87E1uq
ExxvuELd3DGYE29anI58V/0L/Jzib6d13JqfI3ThLdU6qj4g0fDhTpojDAZ15CXe
hYBGmmCxAKA1EMyKyZ4w77TJZrCDEOVhOIqT2dxClH1c7hmGu5aldbzvDT0+BfK9
U8cywZnyQPygDf3RMgpgZEEIqkk8RCs4V8PDtJjXZGLbHJuNpEtPWUs3c2ngaK7D
oAGRE8CYQ7Vz0nZDOSeFfPyWwAiEOxFbRFsgzSi117iE9Xg11fnpmltSQfMO2vy1
Co4AK+hx/uJg12yk9XumeofzRSyni8fFTSg7AKFgCBwhzr7PZwStadBnhYXwgGFJ
SsdLzmAgLdvNC1kItmn8TPztk5Jpim2/zmKUHc3tTNxcKnPIFqINXBubXxpB80cZ
cXXYZNwP20rI1NSVM2C3vYm+nLT+OTIO2Rk7IsT5EW+ghm9EgfsJeW6ARx0uFlNf
3C8126aywFD5l9HL1DGavLMU+xwHn3vD4BsQ/TAT3fKwel4CnEcB/ieYDAhWEDVZ
Dy8aiPGUGWKaFW/gCbDlr13lsGze5HCBJC3Mf9gj+Vf9WQP9KQ/JHoG9iTA0qtLa
4bq7IPwXntzjiInykhw+7H5MXKiOfr/p1+11FbE0t3m+NpvfEmlGBURJBPDEzThh
rq/d1Eo0oYGHJNmFS/ufv3gtWvJxClNkjDwsFPyHPdgKwRDL+I4HR6P9jwYN70zh
F5IuOa9LOnQIvdEX87FHAlffgZ1KBr6eDheOz7bvBZbS6J28ERtiaimocBo/i6xX
Nz3Si75GWTQIzAFGDyLOcHtiSaKdiprxRWbNTokJY+OGmRRtIQnSj3fqoDmrxGgS
8PXgXZyb4oKxqJuhl395HYXMR5TaYTcMjckwIDp1vW4BAIA4REqObG5g5SnEatOh
GfS6qCk5lUJlwFfkZb7eccIISRwb5BFhTebRg9Kud3/8sC6FA+12gcwuKOzgUCNR
hpEYqcw+rpyki0gIDPLNYO5V97pKTyNbLmGKlJCiz9DT0e13sMx1LC/4Het8kaLz
I4bX4z26ZMNmcruNLgK782qN3rU/VfEh0RQ6AvTGXBAnu7RkEd0HsJlGmcLeGh71
KGinWQE1+e56VbmA//ZnrTRo4uECuD3mRZdlOskSWD4E3Bfv2iVUbicmt1w69pKS
qb6bZSGUFxEW7wfZMWjXKohfdoBbwHd/pqD5L7MP3claj01vMCdAaT8kVsYMbiUv
7Mf04tKYh06F19OpqgwuvHtc1VAGhiaRjQ0+vS3KCrP1YC5ilRDGJ5VF75Ke3RTM
LCnaxj0opzqjYOE7y0YEfwXk+2B9BL3jLk6rhNiBH+WPuAfJ6oaFsNmhPNjNdZs6
q2t3nPlnKHZvidUrgDKIE4alZQvrEkOR0TxSI32T3YDsK9k0S61bGzy+vf8j4Wwt
OX0w0tfr+Q8Qy9WHNaci2q4c4RjqJucqVa2OaqPCYDg1V1EzTpRRYQSBAyKtZ4Ky
XXG40zwrH75vTPWy2t+zxMpHdF2LHYEq6Nwswr95osYKOMjdncwCOCmq8okGAtw3
QCCnItbwtF1mDX0jBKpif0i1Hypn91EPqcbSRBuuY3qfJpW5gSejZmKwk+JMjuZK
q2/Vgf2Q36pZlL3sMjD+cuyvFtHcsiOjx0UXb83vCGZBXCMZdZpT+viZRaVyitz0
lHH4FcLiVCnPWaLvxkk0E6Ennf9/UQzDxxSZCKm7Ik/cyUnBFoOa9+kOsR9UDgKZ
F4CSFFEP3albRp9zkVYMFdFvMcNScBuBVLTngsN/qL6pk9MKWem0JjQ80ji5DRTa
zh609YFd/Q0mU9T6B0U7tTqPqcMx05J6LvWZkPUtHHLDsi5KH41bnfkK5efOpgdO
GHSnoDx9Rhe+fa81kz12maqsGML/4sjH75JlPQbNG9RwZNGHSbuj8aRJ7OZetJSM
GkF/RqrGsJn62Q8Vyc1JHrcYL9WSuzn6rW01zgR2Q/qtlxmNLrqZlLzfHsX6AmfF
1s7h2p0JZNUOSopaIgR/Zwrajba3ge6470RcqIrwLv+nA1f/2or8tW8knmJei2M7
ze/N5dcri/s5ihAo+ujnYNkE848lBS4vn/wYHkwgN77vc1LLylG0P296RnH+fOBu
kUZ7TMC5q3USxW3+YjVr7eUXyQUgu1ST5SoooolkppdM1VQ7+FTiZjYOiTvFx1yq
+Zf6oYRJfhbTKqzkBGyx4vX23vY5MoPVxLjcJlopxxWoVkbMAjMDQgOs997QleEG
i1Wm4+NG/lS+t6fguMtCaF5l9SWinairT0nPQNxHs5E0muxvePN4/0x32HDckflJ
35lI5Mjf+5FA0cyRb8Hx7pDfQbA/r0oURTFMYsoLnCN5UybHCIvOqd070ARrXRFX
ehdqSbci6PlvUCR2TNtslxksiMYIStHdQYufZ3s/NhbFTfuEKcznkaC7FmCIxDjS
uksU1kiy1KeaFTXoBmtJ4WBFS4p1/2YoBqCzcEF/GBtsKggirb+vOEKX3D6xDNXF
6nHhe+EoPKwaWL6B0OLto3cB6KyFWXeijH86huWL/MdmKVgJo1A09Ux+1Vtdh5tK
01G1/SlgcIo1OJwXJYwkyPN22gaVL3ofJCVZ/SO5isndf3jg2dr+pL1Za4al2KQa
4RuoCJ5cGfY7D25V4bxZFFEmr632U2lhS58AoX+59yCbrQqT02488O+BVmhuRfzW
4R/VqMS74OMIL8uhKveUgbWPSbUilWOgHqPQ8Q5SEkbRHWTOYEcTx6sma5wYx4QM
ne1kwO5zxfprTk6vgVIIAExeEU1rH4OBglCvuqHmysCoGE0WczffI1s92Hb5whE5
xrnoQB8Vn4hb/eZ6sEqRyh0xX93jK+K9KyQ9LS5wCNxDFeocVkm+FKzMn575Vi6Z
gntit2ZkYHMFexllMjS1EG32wh0wVgqedXCZH9nPlKqeYUxm9nC0c3lJXNlomngt
CQFSNRJs2bgs73KLRdGdTEZ00jfHCLDxjnlidLSicevsAspvUle6uBOwHJrDXrZr
7pdQMt/XMxsM92tw4jYM3rgeT5IpAqPIA56xoDUmGtdhQRGL15A/ytzrBwAFEG0U
jJsPgiXL7gTxiJHmujT86iewuW4iqDByhoyFQUlsUQ81KAPG0pYy+MsWNpejzjbD
1HsrnC50nG/K4ELmSS6+xc45gGnaIqFt5Nr1i+B3AJb6U2hfy0jo1qs1DPSQeDbk
4oPiCC9kQFTzhlr109DukOEcBr4Km5hB/UWfK/QeFxBAHsNnbTPVNmMoqHMECatM
YFFYUBsea0BSJySzUcEdUp8Pqi6F6klcr9ZQ+pQTeTheocoBFyVA5gnhiintnCwS
8eAbq/cePoMpmgW53ztkZXhU25HWpK2tqos0e6VCRSRJJZekiW/aUjOMdwrwbI27
QLBgmpjt+3ijWPVP6Chle0JiOI/12BFX+05KFAL5/qcQDlJkLALUAdxqBJ5IsWSy
tX5b1F3JTWJMdy6OCOrLDh0E1eL4XaC5bfRQUgIbaBrge8YeprT0CWynBYlf3tj2
HkDWEBCNguDvhH5RiL+OYIvfz34zwJIR7sjuhtosTpzJBlKHh3g/4zrZ4M6fvIF0
tiBYWVytRDXfu75z08tMnHPlCD+md5EiPJgtclrsFV/y/fkju0yCe1tpbVzN4kTE
H+lqjyyOBqqg8G4d8XUGMwSkV7YNqYWLY5J8a1NKl0zphBAUMVkMlp0jUSBAdLG6
LUJXHQh/itEzUQq3CJBAtv4mP70BkKrb/lYHsKZNYZRRvPKsT+qGaUC4EnH2PFK8
8phXa6dvsb5NfoQA5S+Mv9Qt8omx1DzLDZQ5XTINxaSikvjzzQ5xx2sIa2tgZqhl
ECtie+gMT0vc8OKtjpFR/aSrlgLSTja0oTYn1XX+qEq+EV78vFKIr5Eb9KJKZkw5
8crWKt3N1HdUYVuLFUliMCnqEOoIui0VhyWgx4g5IZNiRKjfMkR067vfClRJ4mgJ
zuWaViYEm8dH5SEFHmbWY76L+piKwwfI2cU8aXb8m3+3VpZ/YtQqkc5yfcX62d3N
1imilbAqPAbiiet9tPZh5SCQVuuhQOXKhATouxc821G5/TOyjZcwADhCK11rybR+
vy7NV4W8hcOmGL8GWXSWmug952lSI534IryNZwQSACTgiQWbvEOm5hKY22sPqdKo
kIqD36EtI3eC/R2+o10mz29Dn19UnbDjCaoit1OpUpzeKoPty1vN/Vu5w2XlPSB5
BL6mqF3ktwJm4i+18PDcQ2QTmV5zniTKXdrGOQLCUNA6Y2JmNbErsc3lkEdFN0Ee
qN2dc9ek0kH1/iEoBooArKczHewkgmGk9KuGM2B5AT+4lWLfhuppKUUC0wTpc3xs
Cmcj/ptCpbo/mgq2BkZ4Z+g2e8nSvP2ocYq43G1DonxJA1Z2gWGW4rsJS67Fi2FC
4r+jx6IbV7pbM5qbY9gACH9uGaQZSDD7rb24RlJwBQFulZUFY+1MAGTwOCrt/nCd
bDVohEV8bttES/O/ImmdG+jbLTCc4FZCYJVaVoXpDSuWpJgXpdcCpM1du/0HyDxd
IBLtmLrOK0I3I0VGBNWoxnXVsDY7BJl/7jPyRZ8jt6airWxujG/pHGLXxQZAIpRs
XqKfGU0MkfDfOmJS+Ni7l6lsjnZf6BIyYb+nKG75gn6QVX7MQdEMoZTnJbl3B35R
+C0AxbvQNf+ymxvWX56FaDjO5RlJ1n7Q8Sw36RjJYjTD2FM7Tjrr8rQAKHERPR1W
Z7KbHoGGPMs6UUNdFhF2LWkfgQQ1GHX/uPzdvsMbfIr5aWd+UjPrc3kLqiWBKrgb
t0tuKHrsAP2rlYshZ85eDQTTpgmvl1vQolp7yl23XQBy2qgJwdHJHFZxjEoEbnf0
aTZUAzgVkVEI/P5htC+bxkkoY8JgaG8wFhpXKF/VwHQU4x8IWayDo37rwFQfAkTI
p8mKyvHpICwiLEhht+LZ0gqxwi8RSRPDZ0RWHWs1bRwWxwGeCs/AfMDLxSiL1u7+
1JkJt2qo8Tss6BFHvVlANo7GU36ZHzcDBDxYzbe4TFPiOLGkTMllCcBHOEncOhk9
ESi9LABn9SXh0fOlMjCC2ydfHwDo9BzFOXNbsowvYqpWe3EcgjcxFMnllhBRDmXm
ztE0cMZ6z1PzUIzN3mrg/biudSqiI5M6HoPfSJ7DjnT7zr7HH47LJqzxOhrcVgM7
l9xEjOVGA9aGAbcWxqd7Qq5T9GeVheOd46I2AJoVr9dtcvLzzxgAMesRs4NN9JgO
dpCkYGB86wssSTwUP4EEOKFf0KW33k6tMeOlCDYg2RIfiTjvlBw8EaAPNbYGizrK
GhsgzRRVRZ4qN9ct3EZb2Yrb8YmcQMZKJoM9KE0aXZg3/vOF1u50E18nvDaD/DCc
BidiVsp7MnvzsyTB4goR9p4YxUsetqYzbt+JlS1pfsLItYmEeGWbd6Yz0kv1Iy1t
rlVP66xGjoHWeN6hR5bEJAcu6wVAx4C00UG3LFBfVtSyK8oqV2/II+BvVjjz/qGZ
HZX51T6aymzmnjdT/WYOkqfMUiDXfkUt0pPmvYoOBJBfyeMtEC/vNkM5x9usSatY
qqEjY8gbJaQiftLg+wZ5ABnf6dUMfRVnLLw5x9lEeDt6sEgfl6iCCR5W1PECBdQN
8wGE33PbGWwV982vWn7MXz98I3zuChWTklGX4ahRl6Xc2mlM4n0rr5NAKbQJOtV2
sFWLT3TbaI+UR5spN4nOarsl07mCoSp8ioyVGsOc4ACZ3EMsTQR9j5oqotZ9MgwM
gwH3of0G6wNreIsXLn2k85ZBD6Qxf1CxP5EPVSGezFkw3QKGkSN7mjA64dWb2Wvv
3pFxpsuI8UKRuJgRzbAoGSzIomvZve9dFtrRRh0WGGfz6+y0zhnfnHnXdIoZ0LJI
8LksyyuvmrmolTULn1HJJkswTXJSJeCbtopfSXaW0dLvyd2KU5P1JSP3ZMgW2KaS
QM4/xYih3QywQH0zH8PPmve7O0K/OuFNde9x5GVNCOwUZkmwAcICwmDISkzWOoTW
TUfMuViggrI/0E+IFJLwmxFMAAIZXFoamdDryEIb5dqygdfCIs5m6PEgX0vqsDC6
8QAGqj3YeBLPOIaAy4dMdqTP590Sw1IHARYU3kGsFV9SD5rnmAX22d12Mqjdt0lO
paXVV6qPaivC5Du8MnV9C7kY9ycpS7oRXCR0DjciO5AlvhICGv60580sq/OKIKFF
7ce1frKvHMhRMVaBshZzV0GaCizAkVJ1olPg1a6ygueNLdcCDN1XtGDlxpwUhyZU
DT/SkjNaOfLixzC9h8ezYoGMRjDEFoJpkdmIwixTEGpzAFZeaL9edm0xm5HxwASW
CyVSre8X/rMKWAzZqq62kmzWa06uW+ObxFSS2PlgGKcpbTsagvRASu86wApoRiJG
xzTCzG5qVctc/yCLR/HwHN+6ZVVFpE8AhvXdKMJXks2lLs7bsmsbLN0hd0VLqFu9
2ZP0AGT2JUIWT3mGYpfQCv0P404oh5m5+40fkE8W59+K3fuXW6sZGZSXnHCdE7BM
mJiH47wjYittWRDqJ63sf71yyQQpExatrQJ2KM3VlJ/nswnsbPrQ6aVm8I+KWJwk
wKPu1RQCaKVNmRqMaZIUT6Qrnk1OxSQ33TRk9hwJGDv6CxuSfs74dvXNTgWneK8U
8QydUqwatsUBpHsjWrJA1+OKkdQvW92yC1goFAxtT+jSy6xBsT2pBwUu1oK7AlB+
MiorlDiO7dqZ0jx9ITOJlBrCB9lrovZb9jC1ajkmkyGGUYPwOn2ZzAKjsmf1nn9g
G7uCOsN8j3myFqa8Rb/ZjPTfPHQD0HO1YXUY5rebDh3olM3tE3y5Pvix2xXDUe7+
BxaNpTLU/ZU6HdV465P8pDuOuoxLnxuo+LaC+sQHGX2UGN5fAtLy9pJwcxKhS+bG
NBcp0WoMsTNRsV/C6zw3i+xDAkA20cqB5PlydRhMc2UyQmERBqnlKRGeJmaJPED1
QVljuBxn354YI6JI6jj5aFEDYbGosBdzoW8b5rS272xNaxm8fP3BwUHkbXOrlbgP
hicrglYvyDmrqYTxMNINfHbguJQdUL37Z3GY+qhXlJRTK+5inbD1SNDrY5KAbAyO
NCiN3gyz+246n7y1P5OvA9ooa3EN7xtrWAf11XhArSCjixNoAuRlfqWk2LapSKIE
3NkscP1NblpnPXz335HhC5lhar6EVpZZhUQZpa7jTG2dAoN2YpRnZLrCM66LXo1P
LO/vryu4cLzQgOaiFebtI2NQeWOTo/vhavgLuaeLjmskDW7RONe8EL4vwoKehXRN
61gHnfosJnjF7mzqUqqP0P6uNxh2ASuXBoRovPKLJlQeZKdSYPEFzo1WM6JOcuUQ
K29OLUG5iOW8/ZflOI0IQiCpETfkZZdNDauxr9aa4DsK2wzTIR6pf7ALMfcyGisg
kRPNbOOd6lFtsY/nfSxHOh1dAmE2JxHcIc0fiTV2KLcM/1Ny1gtICukCK1e3l9Tl
wK4C+crdgAy2aolR9Ilxpha0vagmOgLDugEbm/hueX3D5FiSv82JDVDZulnNFKgS
ZDfmjcHWRDy+H3vCT6ZkVHq/wPBaB1iT63FwlBJ3V0epv3Q9TgjkPew0sUS/b+PL
u+Qr/RC7lJikzuXZ3h3+w/nSy0IL2tKhEgQI+JdAEGJz+JVMshTCsslf7n+otnPG
A9l6gdLwaZ9XzZE4o4YJ/dfuUjItb0BL5HDN4+scpjPhvnx58tMdVe0Y6vWsGyRj
T9TXABC0S0wZlcAT+wrAL33QX7QEVo84gaih2Bu0Qez+777GznlBAGY1JWkzKi2T
0InadlcXCXuzhkOH1TRNWPT1Yth0KKR0loGDxT6fbBvgjIIpEQbc0R+clpYn2k8f
ynButFHcWPis2B2m0daCKPcIx5+OXMFv/3qXed7gSJ8/EZh2WSKYWI/jqL16JmbO
OcSrVg6IMdG6cBnUv5PZC7GNGZTfA9nOWYTU7fUIuG4eaye52NodNbFVtIV8gsvh
vs1w8Vutb/411oN4IcioPsChurLfgFvp4rbi4dFmhAwa1MEU4/XnlY/Obi9zbMJW
Qoz2vax86X2SkfzYDUKrWJAUurFnWHX84fy+Ur5Mz9KPXy7KL7KVCgl3+d5KhlBf
IRYY3MZQg3Qtvn/ofT37PCB2VCuSe1HNKbGZpuRwYqlINqbj7BOjN4f4pFaahvGt
ReSgFWFp53DCC8Q5rLmlO1q06a1C6TwyF9R1hYO+HMI8HXl9cFdZKz2XbGgtTITx
LrnoO2MyTEbxlNTrZoa8dVNZR39GoKM/5kkAwLdI9M4VnoyZOr9joleIh76KC0Ea
1WNYeofermwoYA43KjCQaRbogkIi+GfGJPb6l5l+yYaxn6GVx74owtrcL00fhYGT
Q5jcpK7msonLGaUwir+uXBwftHxKDK90cfXKnm+70mraju/Nb+8l1r/gX6i5bnK4
e3PuoJrRcde2WDKrGIzi86OMPrB9K7KURX1+1zLDwJo+1tLXaMf52dmHyRIi0yYK
H6Fw01ivdshJ3lAnIjtbREWO1u6b6Dap+wn9UJjJj7IyI5xmGaMhHOSCmOaWLilm
BAIGVLSR03bD7hawHHcKN/zHZlSXabyJWAkx67q95hvLKBqFyl5/UXvcFunSUl6P
QOyUjupGC/OuqlzXl1rObG+Tq/rmcZ2lSWF1ZvQmBAReaAG0bL1rzn3qq0kXRZTT
5lIos0zTtVUIf/CZTKhPc7VEujP5Nxw8yWIkJMlmMbYQso0pWxIBI1rtncw5Ebzg
48T7+e5rZRN5QFqlyB7+/WP/tSObhU/Of9aMWGIALN33iq+rRsrA8VffeqGyZ6UI
uMA3dsQ7w0jkpVdMpu5c5yoptSUSPuTzfnEX9Yn5k6ApUNDcUVpC2OFRRaP5XfT7
4fsxKmey9VyNNh5qFx6zKp8kSIc5t3VHShYK8NTFdaLZXsTvhwDi0nCcDiWW0n5w
KKhuAWcgGtZzjotHTxcLdRJr82mX8U+uiaEc/5A3OG81ZDD7ksG3rOzt7p5W9ToW
0Jn0Tu9Guy5CBIRFsp2MqOl1DqihAmEEqCz8aksR/2+pEcz3S2dxEEYd3Abge5Xm
2dZC5GwVIvKAxcqT6dabjsR/CwLWWKpYuntZ4AQXifj/vWLETWZSR7YXUMc9c5G0
KEvPANPe5uv611tGKfNB574pybnE1Z1bANGRjcwdSokYxPsWeyNJcYprPtAarC8+
pBA1NSlmKzRlL3dTJjJ++XrVkbsvYeo+quHFpY2IABD3rnHqwXEtNvtA3DAazNAm
dfvPaPHssimsJSvscmUDWhxclCGoOT28B3eplXCwqvDm3oG5eb3uCsYlC0gQhYny
axead6wRZhKbyP58CcvE8Id95BSNLk31KS044qECzLOOcbeCXnP765/i6LHSzOhu
H4FaxeGUb0bQzDRBcppowEr4ikmzLgV0kI5Kfs+JcwsoUEGdHIQyA+RADPg4qMgt
79ZJxfAb/K4ecsADpIkoojagOmSk1ICFN5C3gT5PQUNOaHfBDgX7GCrT6sVPTooX
rCIS1MWz6RLXnXCbTfb9u4DfN9qyx/8pueOj9qXQxyfyjJ/UwIjhCOnqIyKjHk2f
mD8ss1MD3jYt8dSONDnXMwYoO5dmpmAunBGcijEEt1uAsA2uNrcX4yeBVv+m3UgS
MJ01pbheXxZA9n5j90Z315YCy0HdR0Ed+MiD/kkbfTMI0E/ljPnMtuo9XS1Q9RrI
0zZO0dYJtun24kYdV4retlf+SkvlzgBxn8LwA2GmPRP+wcig0s8U9+dAaCf7Z8eZ
S4WeKlFVkkymnqa6Twi0PbJ4LvGYhnAWeeFDWasNCQEUkKDLlj1Tb79RLfPNZsGR
nRYAFlao0lUP7coJptK2H+X2vJXY31Z4n+gCdCXYmD4lXZNYRnTY3cV/Hm5Wmjor
jON3KpRjtjCLzOlBY8yZvGqx0+4i4TgQm5KsAd2JhgkMXrqgw2of3L961fDHMNs3
OwxXp0+aT7OgngEFNkDY4e9fwuQ4eA1QcC37TlPIsjKNjGGP4THhrWrUZCjxP2dL
/25EmP4unUtptGRX2HBnkxji6oTX1hSTrcirEONzVWjHB0tgzsbuA5/b+1QlYCoU
ZKTHWkYxWCa24RKbQE3OzRRbFU5uYTlbTNrHM97RJvXMUonwaI1jOuBtNXjwPrIQ
mvhu3qBvCAovEqWHHs2HXzgnPZJ2+qbfEglKe6KK0M7Kg6PT7LbcY62E9Awz9UUq
qTrdASQrISCtss8arGBe6UFlAcHUgZLp0vyXsN5YMDS6C3zMNbwKgfsN1Vk91xmS
4/2jAMxtyjPehVsfsZTEknAJYYcg5AlIKB0koSXs/ZRf3mmrFGWAf9ZNA1fr5TgW
afJBmLJFPACyKPOY5+fXzh5YirwIC6rgSd15182BCqqGnM7es/ZC9p3BMw4xHeak
huZBSZBsztHm3j43bBM3SvAqum2jJ9C0Kt74bOLTLe5yrgNas7tkTl8c1SXmT91l
ZVkQDKYQGmwkEa4J0n2AtI0HYrlRG+bu80RbjeuQWRLCAjsvsOEENwHojDbQcu5B
zszugf++KfhyC5ZSBqhvy0nsvmzvs/x/HIVG/cwPHs8oNNgqQQHhX1F1pKbnSCr+
iUaYoIfqMI6FLUWdXDNbaVKXwNTFSTbloMbbpzl0LKICKARHQ5Y2AhOq+SgEfO4c
siT9hGYK+2BMH3fOkqZz+jURYSIn7eBynnwFvm7TBeOBvdnmiJT8Uw5VVmGgn9G9
hj8LcZkukm60t6UxF/zkWKxxrQ1XMFx2IXVn8WFccWQp7/dIn6QAfn+Dp/k/qRsL
y3Cwj6KHXg8i1dkAMB0zDy2JriTbBko1MkDqTboBotNaOQTCwggh2ivVNwMVsoOh
2bRsuxqUhD1iJ71JY/JcyKN3JjVdTqmm0f7PFQN8cueyctsgoY4+ZZnCnrNz55jl
QeqjSiWZjzqStcQC/ztarChpMauu0b/FXFyxHu4uOHWSK4uxG6t7ho2kn56HCC93
DcwCGoaeOaqO5zXnO6SknoGO3AGDqSv7JIl3VosTpe7ZRXpz4+BzE1ps0y+u9TRR
Udq65PA500b0M3834ILBHjIDfpGW4dKHwqjYt7OsX8lsxw/wbpseIWN2pGiDVmAP
OpyFZfzW8A3NTAFlGg861lO/yZxPmIKu22T2BTI1xpmFelrbflxXaMdupN2492IV
J6dwxQ5xBo+cWrtUvN/f5+gv8bZWUawk/LvGznO/ckKyQ/FoLCHEHCmUcIH2zcBM
8ton7EZkOr7aVoDLMylErxEYZZenO/9p9ijyDgo6SzWnYlN2W8TrYE5O2Xjd9WcY
UN5f4t82Sjnjuoy9Pf7ufkQcB4M6hbORMxYd/Bft0Z6wybZruK9JvistlN8AVutX
JDwwHrkkK/lsn+O+7ECcM/KqBKae77waWF+FFf923RxgceFrVQvDOSwGIhFo58DP
JkHFVLgHB27r5vSuprIJoKojLAtLxWXHYozddnGKJB+zZcg7DDHslnSJdktNpSjG
XyGKKyXyqiBmpw6V3nSHVlT/Kshm4uzORjYTyK9sWiFUl4DxhJCI70W4EMigOlj6
85A8lWscy1GNvjj6/CQPr7N+uuildO9XNNCDNrrvuDED0I3/8ia8v2Qy3oDx82gw
V5HCckHHIfbrpMOUIVZg0z2kuxrD+iixNysLf4ixOLfjEudK9R0sEUCupTh0Fz1k
GTjlHuf/K0UFpUFFHpEW6Upfb9dvvG612V0bKciSR32ccAORerpcp61lrGilataY
2O3SS31Cl6qOOoM22hT1Xow/x1AE6XJ1zJ9aE8PXliP1c9wwnIVgs8HF5SacdknX
LYQzbgcagFa2xLGDV6yS0bWDhb1Qzaf6UiR6+YsgZx0BPFdrqY2nSoi4VQvnnq9S
GzOZFCPZc6RxXlJrgdwkHeGu7oTMpgRXOaI/I7VbBG6DIphKFkoHWf6eJw+uMuZL
FVpLAjoa/Y0vOgqT7ZMPPBiW1XwMSsci7lL6AvSp/On09QnMYL0E5hJdoFooxfK0
2fiRpMiT0cU26B//1qHRmIjg5MPgw+UWJiXQY2y/93GuWQam6ElfdGXgxqqWwDAX
hX3Ls81QRrRZ4+z4vGQ1dOXDwAERz7MlLGIaQgiB3PmP4NqQ4Rtwhhj5mmw+XcuG
+2E92AWJl0tZl3NpkQHxxrF2gjW6fkHiFrD3aAZJd2A9MLmMPo28PfhYJb0m7BOc
fgEVWaH3q4vn0+I55PgjLlA1kLTwGH2ezSmet6YNndw3izKWmj6eqqtdBxlHnY/P
8BVn1Z17117wC8VrdYyevloE07nBTTjlNuxKfPtjmfaJqy3ed77gY9YJSCyKLzdV
CSx6x5wlG3yflAWBJwd34YyApYmsdylnmj/uKp0DCZ5SRKSRFQK6AGf/5KFDhew/
dOIQUbVPALjKto+MlHfmKxALR0FVawmra0rqAdIacV6yR+/8vLshih4af0BUY0di
tuEDT6su7/NXpKQz+cC51xvJw52IxKTVAGjQsTLaHTsL60xd2XF9YuLBjt1GcxSA
sNij9Tym0F2LY7YnMwVIq9BMR6H1jZgE9ZIGpxCTq6/eSLX5WIda+sP94Wc9AgR8
k7ObmJM1DtVIGIRcZDQyql81xjx0Yygenl70vfKQvRV1XzKYi7b9bdcGnbAo0Y1u
kNXWri7qn6DgmlC+4XdG5IqDVr+Alrs8Vblwc2Cu8YFkHyEi9OO7gARI+3dvA+rc
YopyzoWJ4OCpcwohnBliXMPBMD4ah6ghZGxrvMAAs5ldrEkdByO+//WrFzGPk7DQ
lJFE57pdQyaGg6bCKJfsvGNDdxIt7oC2iiFOr6IDIaWGmnMVLlpOPvGlFm/6olzQ
QcQcnT+9DzJf8lKC87vcwL9KAjVr7gQosEsWjwDC4+FMJLb6+xdhSlIXtPigfq+c
4Z1HoKSIUmOjvAu7xcb8O0rjMXgbfGCYZf99cBk2A3tSs4idbF44i3yTJhfueTSS
/axu79LT6JSwp0ncjywr7Pv1bmUphzXTom7ys7aUW4bXhAeTywbPR9EJRN6ae/mF
FLoHZE5qc+dCBSCvwYipdIlkm67m/fz0uNKjMDq4obxkGE+gTrM+zmSO8H+S8us8
3TtMad+r66YnsUd7QelWyBKrAtzOSiRiiR8gUTOLg10fT3fHt4DthOEKQU+YDDSF
+fXzU66bwLU82SFpq+6BQd+fDQEXu+L9gRpSFK7eSdbTDIsrDuCxAQcCGEfu1qkk
WOq4IAPAHYJjFLcrC3o++HDGEy+iryB828MP0LrfGjA2i2ox8BpbudA//wVxXmIc
2vnUGdhRB2AfkbDSptITJxktvq5Ukle10oTvGKay+Q1xj7n0Cdfv4IiRLH30IKya
Pa7UN0bzfjl+3Ug4vRN8iYNwc1dyaroVQguUi5+SqcTciYwQguPG/aSqgrc1EapJ
+1nrs02T2UWIDHNPlA5Z9nm1ElaEb6eG2OtFM65qqy9G21/jyh4RdwmjNaurisvd
LZbIdP1L8IEzKBNDnYI0eDGyzNLNaUxX3MnGaSxa5hvZetRHrzTjbs3T7EEoz5GT
TqNiF6ox0Odo0PxDohmdashl8LwWlDEbA1mZSBHFF7ZpvQo4NHPjNOfUMbUMgx1t
lxe4jbFiamUG+Uw964TUH3/QDCGGpffvY1Vs8tWYaclWCpUQ1Xc+immb7QqSYE/H
aeW64F7/Tr+iEhtEvG1/3kiOTFMmcOsvvZGzYfoyQdpUiWNronL9lV7CVl5LfEA0
vYA2cw80S5VD7sEQ8TzcjjIeeMJ9LTi29ixhiAumARjvm5CKeT7om7Z1RFBjL6zk
voi6UfNg9ZbfCVXTxS6FrvTfHrVZMcgFCoIopLKdBKR4+JmGXZhBGaPqkjVDvtwh
Un5bV1usZ9787LTWhETHUxnRRL9lYFsKpTcgU44jg4gxA6IdVTzvH/7PvHM7DDRr
SjfP3GxGNwHbLmXXkvZ8K8OcBVM0THzRbUf8GSgzMeZonvLQtT8hbjjMHBBCFTNg
ITq5hk+W7gpwRp5oHqezCLutHcggTkj/LtlCl4DRqTKMmHG8ROsLgh2DHxyaidvR
bvcmIEwKnjXTXxwCFp4JCUkyvjbJfm5kSJLtK+nTHw0ZZik0xrXcPwR1SYwg0U6+
+8KhApPbwoUeO/zQivlJK8Nn34NT6e5180G4v04jW1wCeoL6AQ9qiTscExs1ADWA
nFzy/na3ksXcB6qcA1AXawmO2MBa3Uw8a8+yvIvM/jfNWNYsM1nENAfP22Jp8TM0
dA3u8ToBE1rqphuFDYVQJWTOzre9+PJRsmrtE6gEgFsW9dHZxnXx6D7yzU0l7TyX
9hnhOrRa6dBeOBwwGxmSCAY6HW5GjFa/bu3zQ3v6cmBTN+OMUikYZxvw/qPoz/qc
1f+nUXdRm7Q+KL0KC5uwHtDNIcesEHkQ42rzQQ1OYnkcRSKe5rW6kCznRIMMR71L
47i6NdT1qMgs6qZbtP5fm1JS8kSA6kpIiMmHoSPDYAuECbzIapvpim+EWEF5GeQ5
aJ3ac1hje0oFqxYq0DKdfNuzrMtwHNFR9wHAKHHqH4Rp93RsTnaTdmyqDkcps3Yu
+/hkpSnezodHMZHtjoL1QI9gK4th14MSn9qaIYW3+M8n3xY1VRCJrF5KUtcCMSp9
8CXGGj5QCwE1znhclFLJP/V3sd0JTUKKF93TSDKaMZkmcVfSw6N1sE5BbDG731uE
SKnhQM1rPqjPg1+KnhiVbWBxNEcaTeWx6HZjcPaoPJKLhNDk324XMwV2hHmi4Qr2
NcbXkw3T+5rBOTMFv+mrXXvz2JgRV/cLX3MzUoiUfFPDotr2x1VP9y4Af4yNTIgk
iYPcALIf3qW3J751A5upiUUw9rz9NV/+hhyQhl1rlpOpj1ej3OiR9y3yUk4gTMj6
w61CTiJE8Uxo0zwGBr8jafgxMCXTvU/CUBqXysKTziw0cEvMcXACSuakdshCPNpK
tRRg+F4rkZR0Rcv4426fIvYUAj/Egcbz7PGtmli62rxthT7xB8XX9/nsqUrh1dzu
SxaMosiD7B/dDszi5mdIPnY5Z4Nr8thageNh87G+JtXKgeIICRDWwPeWKF0GsPLf
UoU13QCEq13wwMRzl+KlVpX3Hx+8gWsthXvjxWyr3Bdekwdw5wyBbi510Yr/C4eR
o0w+ARDQH7PN69Smw0Gw9Fz68oioKNvRM700q+iGI2hI+d+/nu0xMCHpHDuS0dr8
yCaezuYhZtNUmGsrH8sk+HsdgXFuwaK5abrJUHDf5rJeXnsARTHwcN491gLiQk+3
+259tGWEXKujdFIrd9tvKODp2tC8Xzo7U7YvhgLmXEK6YYd+uh3cOLSwC2rjkWFK
FguISGTn3lORdnFtf0AgjI0xPRxqKvOX4W42m4nwCxjWy/57NgZYeYgk5qbwpvzw
jfcFA/9n8TkbTHay55/rMSLUnB1xDUKbFsbkYzSh6qnOqvu+/zcsA4aYNZBF2M0n
cA5pokW5K2MHtzIeqKT7EDCn3qA+ek1S0ajddHCD8iZPuinDzZ/ZlQSv3+VmScsZ
WAOIpdTC6i6R7WoV7LAkL6cGJnAWPv/GTrUlz28dB6Rsq00DsiM03jpfffYN3lsA
Te69sAZGiMLbuL+TFVPfTcS06wUuLr/ePt7oJkk0xeNaHI/D8+KxDxnBO1GUZ7DC
aZVWo/lOqdN03DIufCSSAemi2lG/Xjj1KHyUGE6iPaIXq6y2HGYzi8pvGwk0/+lu
jW9oHU5OQuqX02ELIyHsBSEd0S4/0o42u2mfBj0AqPg5OG0g++zk2pCqEO92Hcow
UqJ9R2icTc173e2Fb82LfKivYPUypEoDmiQ5rQQ3GY6vzq6D8Tlv0ZQSSmRG4Zqd
bXnFCagDCr6CEEfBiht8mfwUyIEaovox2xw/YjeyP/X2ZM1/oEtsnLRFsmfMsCSz
Uutlm1g3KlqKrRFgxXs10B570RXkae2IrFXnkgUE87J1mrWT2XASjRECVZ73iFb0
gg/AFqpFRngAkBbFUvxm8BQ3Y/1kLebVPieGV4IFk+i2wqtVZRn/wyjUGvKvi5s3
8OWKpimkm00BlP4QQt7QUQ8JJ6p5aEEI6u8SvSwsqzm5DUKlxINlLsRwb6zG9MRx
0GLywU6d39JntRZxIXiC50lAuKbEsVyFuDz0nHdIWs7V57fZvpPpf+hcsN7jo+Gz
pDBCSW7G164UpUvhhZokdF/j3vExXhNGIspDcNG8p6cKpSWbiSWdeBmAXLGBvr3q
w19jb4x4Wj0tk4PzVryJi5FxDTL2SlJTNHFTxd+Uf8Ygiwu+7vDiwmc/8tsPrH7V
6yBLSSJe42eDUN1P1hELElDnljuHLRihg6t2XlfurgwGINKt0siJj35sceuHg8j3
lVQGNsrCLzRMri3Xy887GkaKq5vreA0LPMdrCmBZYphWIkq4CcAofExwIgpdK1QY
gyYKMzsnJV8wgf/fn66VPbF+dUUMZi/HuaFqn8CNb/8cOY1tjJfFgcSPx4jcSAd1
6H9Tx3HFZSKhTS0hwNG9gGb0s7VUsP9l3nPB7OkD6v+TzYzolIzRhfFubGjnvnv0
bITuga8oZDTgTx39sT8HtXjFYpF12po13Bgxme2sWCN4pu/Sez/EzX6MTz71RZiH
bj1Eh9JA2uePxVPfyKm+0V0S5R677CkFyKCsoj4MOTUEiDlwkvVS6u8tYhRtqafc
sb3kHmsKydSSz1ADgl6BpjdHBZhDvYTZrsfZL0Vw1Bc/gh9RJP4ztv8V1tMYo0tG
KzdNmyf/yVtP0nlDVRZ9JYnul9BxHceUACGqsZJZLmOh2jYptrpa4xCoM4vMpVC6
JPSf0yXkJTfp5DvJsKIa99qAy6uO0JNF+DQiy0XhnLTLYv0MyazYcSEPi6wBd/Vl
1y+CYkAfmUa/oyGhV+ilrwucVHuldEHL/ip68cgKrvBDFTD827aiP3OZkVB6F0cd
VMa8QVKra+d6m/9ElIL47CprEB1NmjWe+Ctfa4AOr5aXwjlwaReVzetLs5bGbG2G
fTqB3DMds66LEQJQHn/USN6mWS2Tj+q2P9hherGBxAoeaBD0ZHhS/TccL0slMasQ
dE0q/rALjF7hOUIQDhbfPJov0qd+um2y+ymSfi2cTdj/QcoDuMY4o9s+y+gU4feL
tR5dvU5Hdxu4+oAF3ahRBLM0KK0pDNlNtndLeh+a9Jw6/2905u4meZiK6uaZh6MG
iQYzo60iZG0ObrE+sqz7RSmSUysLl3tUOeEgPORnzDEfU4W+RQUQS8N4OVYUVeLd
8t95aPuAhtPSbsNzx9bz0p5XqjdLXSdqmp0ekROhwOg1Q1G6vgQeVY66lYyY68WD
SejaJ1ubgzNV38r6fXFjDEkZC772/zu/MdukryS7J8sOSK+XKepF8Z34VbQdQsbx
XBb6i3kYNX7UBiiIytfOLZsS0qZIkB4cPzUTjOYb1NhXwghcbAv4C/5D5Ho1mS7a
78EykKluXpXTAxqjU7MrZYI9Xz1Jk+X+LxrmCQz34bwVcJZK26gmN/Ka92DCSf8B
b7KWes3SwXb+8v5VVdzr8P622uXFClIFnJMC0D2mKdtbOZrM9BXNiLXpZeTDlgYg
/3TfnBbavMryT7dNH7ny81tg3+SFVhC658JtVBqz9NqMJKgnPieqrXuCqoAzIqYC
oCfRAdLQOXEvMPQ610em/iGMj5ni9m7Z+IZWSHtSdyHeP3jRvSr8Z3Q492jq88AK
uNYx5u4zZqOkDgQb+hxxB9aftPVl7mhUlx0b0sb1JCs98P2cTKq19ef9f+c6YK7K
OeqW5sWmmduTON4nb2vp95gvPpJdAs3kQLvvw7gLZgeDI33bJRvrT5TsuU0z8roO
1KsStxFd14HL9Ov2sMtxhY6GZN54zQt9lWTGSu2nmA8bCYQUjXzk+tk4pIRuQN9D
FmLqFII3yZwrZkIqFwhDR4EJH8p+rYVT01ghpuR+/x+7l1oGO83B0wDFKYrGP1Y7
plFL8yGVnKLhA+SLRmkqJgnPW6OV844GjpsUbhT1oPWj7sfLd6Z1VCQiN2ZdLXCU
mFrlmE0+kNvdto5eI7GcgB3s/yPk2hwd/iOrx+j1ygvJyp/pbTBxzFslv4YpSvFQ
2kra5Xi/gBcE/jUCq8R1PNaIlVXSsVHB0qy3kHlw+4PSO7gXBzJAzH5Z0uc7jOEh
h75LhovoilFgdNtKqiH0Id1FDeJfU9ofPcOCamq9ylECY0OFTJtOWQZtE5WY13jR
J+PtPtxSCBpRu+qYH9pDD0H7xQwwZB8wfUtSAClx1gcwecI7S7ihmYMlcynB834y
z0ql5F/AWd8oQo066TQsBipYc6pEjnLn20PNxc9Rit22Gaxqbzi2r5xxFvCHZ90A
06bq+HclYRgox4kZpd6zxHQTUZmokD7+6fUcWlIUGPqxlhLATf/Sj/2LQHN8NmTz
FXO7DFib3Ur6DvBESrukbZVbMPmrpoBLLpXS8BUBWDfrcs2Aa8q6H3KwfYNuW01i
TaeLp1VKXev7Xm6cVLaBDM1TZWa7guFpBVmnULN/BroAZZVjQNtRrqnHHUq180sQ
w9RXtW1La32YlluWkwP5YyGZ0aYuBbesJmH1hlm374yImOblp5ClDBZcCajMBNbO
2PtTXMvF2CefF9jYX7XhilSsmLBmLKbno/ZKn/0kg1StUxxJ41yNJCnLoiZFyhc3
LITWgij3gQI/u2Q5CoknjfyTF0bx77Z7hMLXx1LHi039AXQxsOanKB9LsdvwCFOU
Xh/kYwEyZhvMZpYdi1bQsDBv7LbnCxVlFD4YoiE35EO7YHeMBr77vDnV99VRc7MI
+OExP5vjP2jMGS0FWCoB2dbGbVMnCpVITbHs4Dip2cXMPAjCIQeNPHKrB6vgIxcF
RHYaBeTKD//3YZjYJAwCIZHtQ3WR9bRVYczD0p193MZpR9fmr6pTDm7Z6AoSEIDw
pFiXpWMjUJ+DFoL+KYjv1pSowOVxYiAimS+FKmp3nNO86M0V7waQkw+xOIdPzTLi
0VkcXATRBvIdVnx1qMuFxbkX3qYJgnKneebdXCvsfDZKnyxBM44DMKcsLsfDMbDo
a2yaU99mKJCxscC8kb/1EGyObG+q1xapbVS3O6iMArZvUDeiwrn4DOxBSNYMsC21
hruOV3JwusKiCoYWP5WfY0H5XMhrMP0yzoSifLE+48vUr6fERy7Tqaix1SADkMhL
aSrVE3SyJv9tcndkPQ0xLOOcEa9ZQKC8MYFGkcC04mj9hbc5UCxq0ydhhH7Sjte2
b9PJQbtJG1tVVQ3fe816ILqEcwWGNq0UhUYgusshbwBSm09IlPLPrRsVfS5famUg
5nrYI7DsjJvTCyv7/3v0U6N4KjmTJk7JLpU5HgduzUo4s8Y58suVDw8JU9xaeTwJ
qd2swSXgFeI2xxxGuoHBIHGgeOY8zdCh88dbUeYkyuLcNEsFntmb6C6h1RNZy/1R
7EEbmk6pFTgBuck7hXU/yBkEK7x0WFwSAzPLOCIWSisyg/te8xtaTo/0Kd//1Y+K
oeVuXAeZg4rGBbvc33Ga1ruXLxtv73YOj+q1TooOkfL4F1nuYgYr9cqdSbWGtfPB
g/SsxLGGGiB77mO4HqH2PQvKn5JJw/CQpKTF4owZwt8GrQlGq3S2gkKX7MeextDB
C22q1pQc69VBYwWR9V1g/M9uR/DPvfJBSNKYpl93EAf0ZcQVgP4kfc4XyVpO6W9w
WNAI6TXdYradMmAGICXXFedY/uRYEHYJOBofTXf80a9/BlVpIt7sw8fbPYtvEi2S
HHyFIIueTTpFinEJOmIUcJk27mLbY2D251MR3UNVWwhO6/ppffNSLkApfUdv+sbQ
ZNp7VwsKU5DcKUMCFWQdyLGfk6TPL4uSBRyseYwxBGMXJLI1jR0Qbg5rf2Ns5PBV
KC1r0uEqIZMS3hVI0SxA53aZtUKnPEIVaL7dCwLSQR3ZmfSBivv/FKNsO+D6Geg/
tzerrNNsagLfw1G/mqIcT59zULiHEOT+MkUK0ilUWOm2eXsfSwoTOu28WuJaTngo
J+YrX7oqxooPnqnaZBvS4j0N2zSWXDRo0GIVfR8sNJHVCqbUbwcfWP912mL9W2Rk
6uwT3aFTVMhtysGN3oJdTTtveBIov3RoEZxdw5shPOdZEe3sORp9+9vSnh5jAO/1
Fa3tLEbMXb4jG/7wNAZBwEwJBZkTK4FONhOg7fY31zkG6tY4taLzYoarIFhrP+Tr
uL9k9VMQAbcdJ0pdZXQBQmM3zukbXj+OcMavgsOdX8sSFpja36VFCG2bVO5XQJE/
nWbc8gnhW+rW93L+DqhCeKHLAQJK4eYlQ15lvdf6lMgnJa/itjQuNCzvAEPmbgJR
PKBJvfFamQlvZrV0h9lUm9KxYQlMwxb/nMOr6T2paW7NtX0oCOw7zO6RNjqNvdVq
CNzrXe3qbQp75fDYmpHgE+osv3JVCfUQDb3Df/oDvYN/EXjt8+0ACjhnp8cJbwlF
mWLPwpbu/pYLr045/L7l8zS//IIyj2+efL5Xo4oCrabl5Qi71Lmnt/7TZDZEmGtq
pXbupMBnCxgIYia3jHy18H9y3YCGS46tJiAbT6EdKB8nJEaG6GnjEvfLeXEwndI/
ySXyF1KrK6MwBV9khhApRq3uIA69UO85+KqrG3kSSYD/5DVfpk/6F8Gd0hYWm9+H
L7l5Rnf1GCN9Sg0OI4/wmnJK0LxZWoaq2bv8rfT0zFwHb4WZOSTLkhFx7b2EpoAu
9cO5qQO0JfPTlHncjgNV/AmkXVAl3sm0BSKuuRvV2c5D6mvZCxi/GobJ7iXpxiKR
XueAeDJK++SkYsU845ZOED79GNCBGI7KLqhU/BRTF1TPFYvcQ+Ex0VaA6DN1SYAs
sd2we8pnw+uKANZE9xPAHbRPAzyUyk64hTVovhnaI1a5JcCMaUUodfhKcHSk3VMA
fbv+SRDHLp3BGp41OcSExmAF0pp0rUSNILjZujrhiFWiqnQTlUukSZwT1Ymghk1g
9INWFIOShCfUaA/V2n7kl5N7qWx3GmxEt5OtRga/ZFSvN89QMzioaikjptx8Ol//
0wEo0upczBWEmewN/iSLI9yytuatq0eaB5nDiEZbWvncC1PA2+eKO/551s/spLAs
MLJsd/Da7hymiRZBfozV9u0u0S8WewZ7de7SP4zZfQk/gfK+bzN1V4y4WqHfX9Xt
AB0fBl98sUGEoIV7wMQjTVoAA2GctOhEMNHg1uWhuRCo45YeHEmdlo2K4YdKNrxk
YQWzBjPnM7uAz9iFUChLn4E23Kk6OwtVB337ejmzBHZBNejNtKjiTYcBv862tcZu
5JnKnlK4rVbFBAeSqu5wHAi1V6p2gPossv6y6yYtLBDIgQMTVSxiJ00pA69vqS23
r0i/xppvKpF8GYR6265NDlbkQX82ENSFzYkX5IPjq+A5ZIrBJZ4PvVkiTqVkRxqG
r6rb1E2zjxPGakLvZZwh5uq6eJOykmcGotTUUeBGTkzBuC1nb2niv34xBdKtaFxV
BvQYUt3uVFPSBthPWB1Q1g12I3Mi6GlohCkvLXIRIzjZq7Faca+V3IM+RMQqzjxC
xA7keNcId3DoELU1mVV/pQM+8e6qAo1OUJyITjdKb0ceeokzFs2fZb4C3LymYLLt
x4T9nigm2fL3Zr9zH6ksD7xOviUdDLCZhzsLl/t8uv8WyO0a9wvDU2h9c1Xi7qYx
Y+TxibaQhbEIkXRmqLO93E6PnBmgvlPM2xp79ctxfB7NynV20gg+WBXvYTocy0Sa
UxmZfoC//p/hAKZpeFxjZ0cLQf5rSO6k1fFgbx3rwrw02zs2EE55eoRV9ANCgQYW
QPUwzh0nAcshFY90FIx2YXxFBqzqhJRM98EtRe6BBMhPj1WDcwSu5HUnnrL7IbKx
rQyaNt7g+HQMkYRdd5XiOhnfmHcMPLvuW9c3Gis/OWtZ1gT/qP2k5q0AchWMm04s
uD1ic8+rjgzy13m1o0rBPC+kyraBB5fbgAPoHeLwL2/PhzzKVd9LO/N6q+ZHn/mR
MiLgYEmcP0tLZbj+XAwTJl8oyTgLf/JUwCFGpwPON+2XqdbyIQ3uRMQe3Ne12UX7
/lnKVh5fMCs0OfbYw9hHvmYIesPuC6SuYc0W/hKlUqB/iVxNlFm6F3xWs1hFmFi8
RuS3JrXwGRUD/0K+wr0ygiVY+KOjEaVy/nDfxhHBmy0F16BbqLGrW9REaYTfvtfd
dfbL0uToKwPDKwiYbvMLea/sYCSQx3J1FB76dSOSMauXpyljNOhziOidew/WAItD
n/OyKkuJWq3oLEA9Qq2B2UohlvR6AGxKTzH7UKdUt3xFbihLTeHlOcpMKzCxtLrS
PkReDbCuwpDTeHa/oxp+hteeWx66QMt+8DoWAmtJ1F2otLrEe9bBAsYn09CpTAOt
b/bxyfq98XA3ZcLaqV/MoFT+q7f+zt+RaEAQoXrQ5tp27Pc6K1hnRJTa/NJli2f8
S2RRkPUUdn+Obyh+tCJXRWae1F36X+bwgsnSRuUDIcid+5Y3eiL08QcTUWNWPKue
EeYIDsjj6XOmDRUjqyRD6Jz46ge7/5QX1GlBaixW1z2s2OtrfleqbPkLLcGRBLKU
bsvK51lVcoQAsShvqL4lurJ2tcRp2MbniYJhhu9sSrdyK6I821wvs/714EEpm2AR
2ZhbLKHJclSYXvH0r559GvGV+7Ki06GLhaq72WwRkS5ZhnR9iaELvDiIgq/yIpgP
iPQViueSaXu/t/MsqzG8jxet8pT02c1LNoCwCs1tUhfyPi20VzGxweVMBYUGcluH
KlDvILK+j/dhm5LJl3DDl0Xj/noI1fxgGr7Ywe4a4j6A8VCWRpJRbOUc7Tvk/CF5
wJa3h2UWTkYGUldSLknO5i48yA7KAap1pNuN16fVynOWBry1udNGkEYM6sXpm+qk
8U82qBCxxdZFoGw8SzSAk9EjIBmzu7xJdiQ2sM2R7r6B1dIhiIxhHDhUr8UskxOk
i8P+1nxHqIKMf/Of6c3/up7xcX2e6ekycyOI9ht482xwPzn9NBics/nqMfyfNFtg
WVyE0V7p73FMAolekjajrvuIiA/rbkSPESvIEc60vvkmV+UGAcoEkA998yslZQmm
t3OZi9m2TJpKKRBF1wWOSS6RDwp4P81oE47nszIPzcyiRFm8HXbkxlVvm6PqXfdr
qqb2LHlayAGBTNNpftu+RvejCOWbBLU9BcFtubRo/FYgtcjrXNGKC5uU72OGBx5p
GahHOIAEdNMkwCZZcoWr4HQcaEOtOd0lFRIupB7m8eYyCtJG2bWHchzXWO3vXkT6
+aYisBvcECc2ZyEUMPbb2b8734tDRbU60Brb9BliPGOCaci4LUiyRfvKPNeUfQoS
XtqM6W7aFt8nnPAMmkJsyUOgPMkhLTUXnsGYMu4Zb1FLyXnyW1rkJ8e6006BQNf8
BBibNtDLrjGvIR7yDtPLlQRQvn2n9qk4w8kJHSBaURI4VffqCTF3OCNSUWWEttuC
gJoajsFyeFkrtsgsejD48aHZ7kLjbTH5EbZVWAVGZbPoLH2lodSsQjvhjTMVGGRG
WxPaujozkqcUGvJg1AakoYxx46qHkfAS9VKeyZBjG121lxCtHoiZn4nd2nXhQFNA
Vaxl+qTVdZy3tECrQYUAgyoVBj5tv4o79IOxhZHVlXCIZ+vQacacaG1eCSR5VaRd
TWf6nkETEXDpiL2n22dWr41mGmPbR+KDD+HTCCDvnvfSmkv2EdwCI4Uq+AaNEGec
C5HLpv1O+ocDqMnXmxg1kW24/NkAaNTajTgls1tXKoKHFUtGcU+3VqRfgAK+N0rC
wbgtaigOSqOlLTQsQ0KaRXBdlzm4/H9/LFNEcR2lX3B+X2ENUHSnlO9U8ENErMx4
/jZGfbKFDMLPYISae3qaAdm/jzorG1CmPcgSEGEoQaKaZm3bDpztb5VbpJqsr6ko
Wr0ondOfRplIGHHUlW5leR2aWavAvaZ8ST7WFFumk9K7pPpjP2mUXe5td0Aco0Y5
FjTAhKGpQJOUfWSaFsUcfvZWD2NdPhGkLjkI+l8bWDxLp/REEK/wwIjZ8mhsNBkV
9xaG7Dvu3YnItxX1Kr7teWTNtpgFV4xsWvomxmYFo4d60KPYSNrli8vKkJsHLuT2
aHqrSsWU18QZCYUu5YrjhMOEsMv+JIGych2hewF5D6hkO9dE3HAqR+AN2SelDxen
2G91vjdvB2Q38zKqaUw791ClAgqapvq+Gk6/l2Stc02d9fyUrIRsoMv8l1rbzCZF
sDSrZkaVaWGGpbGn+tKJHmX4pl8JHsWCp6H39a9jIlZn1jF1YVkOOx/spMiXVMCT
6UhR+nsfNt4JF1bgmcUaoAirbZhtvfiBa2Pt/gUvFOYNSjy78yGiz3DmgmFufC2c
DU4x7cqUy/QdcSiEfVuHNZgbR8bz1w6P8j6q0X/MtHfIFgF2VCfzfCs77FVBUG45
XvZToPL2AJiVILHAYEXJoLEYlEDfvjxwlR2oDxIx2ugWSTcWVZ6MQCrhePrpiaYy
OFWVxu0pbDd4syQSBUJloUHzK986BPnI+MucqVjB0uNiJc7xck6FQ2deC5td2WZn
RQ2mlKwTyCUpqa1UEdWkMI1UUKV1rZ2pebIw9pmOgz79JvGJGs12mOMVlcqwyEya
MWcFkpLldVTOTpITTIWsJ29fBmUU3W9OY9YHp7+M+DO5rUAFSVLJb2D31df5kAwt
HSKA/pz7yuHZBXj8HXtIm6dOi9P+BwyJkDdfTu95F2RsBKkdA147j1TClUoRoYyl
wOekL8NO7diVsLx/odKX8f8krC2/FXLoHdpDA2qq8TKlWT5UP6XKZJ2msqvDtBrn
7AKmXp6pUORjZoq1lc1EwgiIJBQ7TfyxlZNeqqkB1YDgq1Cx0Z3GvK4JfLz007uR
2GclHF+YKX9TixYQbOJw4GGc8v+OsZH4MZ8lJmFzzPX0rPXi/gRENX0iuRXxJkon
oHMCSOZiEX3W+2+dSYCkS3bJwX9UR1CrjYDzS2AfOG5C5y1o5jPwIokWkgpUDfoo
Xef+3jhzug3heZR9BJ13E01M4kEtVmoMuDbzfYvlDucjb2WoLoK0ibi4fkKYOAC/
bif4628I2WWoYvQZ9HYvtp52KfyPKTenZWfjoEE09geTtf/K49hl16L2MD9RcP5D
frH9YlXo6L0eD7wYRp21T4BxsuC+0LhPopTVIQi1tSohNHlqZGZLQK01lXlMB6TB
+fGyvSy3EP3cuj3PgxLdK8JbW15gvpDI6aw4+N+2ZNP232x1RO29aR6B/xJ+ZQY7
r1paRUE3BUSMtqoJOtRR8nydjFNe6KvO2p83mtloKcTDwm/YDmRYMUx/JMB4Fgau
MlwGJeT0Il46a5vjquIuD51xrTqc/JYhy+s+SwOEmLE/jAzlESsK2DKHbR2oyxQU
kHVRVfZPxiVhnbR7FO22RaQtmPAt5hZatf8pypjQAOgOc20GKmxDKV+v7zFLcE7l
Lfwi+S6a5x8acMdsvd62jodC+/TYMb6UB78IosIuUHMzC/asRASLhp6cITtovtYS
3QGpSDN9T/m4yNZPsc11HOZZzEJTEB/4VTnnJid0eo1c0dj/XxH7DcGI27lOciHA
IAENuVJ+qoHOmtJcr7k5lj2jAK/KQHM1WL+M797IKr+EQBZvrg5ywCBW5uPI4lni
qOsumrM8ZXz1ib8NM5yj1P4s0r35PVE5vKVMwWyw7Vs6rI78wzTiGF8fkeyIGjvW
qrNrI9NUm8lwRHLc4yyNrlujbd8DnX3hxZtnIBhFFX+lt4ZoW8leANHS+JvHDVTT
XsXRXNTM2V6vBoRn0KXzf1nlaeJh6wQ2CUwXkAoIXh1u+rC9sKjApACiH0GufKSy
FOv/lcEfCrvI1yF5y0vgfwU9es7xW8P3xZG8HY7LjRy/KbeAbgCq67tlWGtHyC/i
xQlaJIvjv4ycWjjVp356a+OK/c1PGfsmbuW4bFprx3exAI6+nmqSMRlTXTlIauAl
rmZ5g0LM1nvOhFqcUer0jye3SCJC5NbhwIwgAPpKQN1xA1kU56874Ji/1DgYOGFw
evgXdx4kcm83mHdLlSprr40Olb1lo9JtJ/RosAjhsfDNS8XzuDV630SjK1srbQMU
P9psFH0Iz6ZN4uhYl4USYxXbo85U8zdv3XvmsK54bDF8kb2pQ4+rXRItU4RsM+UT
GAmvzLXolWlP/w8lpKTjtpF9d7LomtZ//yKGBflLC+vDJi/amGjxZrwuach9udkh
bcnrcR+9FZWqupM743XAmaHfeInlyk1i8J27Mhi8b+avGAkqfdAvxgdgKFJ7ZYg8
YqS8UnKSGV8M0aQWLU8TVk44DpLvTKS3BnvbMR9xZSSSTPg3JplcDDEUtU1aVVtF
5yhNLAjjPDkDJxhBCmpPxoWfU9bptV0O7OmiexkDzwdaj8/+t6OSZ5743xaL9BdA
Agr2/T5+IMVC+BVCHwH9TfdYYEKuPlTUjSWKRInrzEYbg5YOVb59ewIOVnfX67sj
4sk9yZwCYMzTgEqpOkp2hm7m3zq4A9S+MZv5gMCpU4XBLesnKELq5f8BucPaT+m7
lPO+uGaAM5yeeJJQpAr+SnZ2m8DowgD88xv7HQWgKN8CyE2L34+eBpRgDc0mdJjl
HBexRIRiAfvN0RVVPoWsgWh9sxZSCs0TcPVcalFigC4GjufB/ZETRItq/0i0E6uA
0l/iJvbMHmMy+e6HUncoacGuikrKvwfzmTuwAYJLPTh3ff4KfvWpl1kzAonIFkRC
uzbXZoAazwG7IRFXovFYMBeu52MHPbgPVGfUhleX977wb1XKbgPNUFodBZheUg5O
TmNurJNF85NiCVbfwvRMt52fg/HfUclRv0qAH22+DQALGnO3O9WPXmT6E8vXUNkP
IS6PE8/tnPk6dJ3rfLuwrs57oYjGVmLMQNT10371nEoJXTvnFRxGlhoUgNiwKx8I
hjWPzs3FXOdR/fd8TbBi6NJ/ZTBe66dRMbN2UZtBjQlVlS+0O6+YkKUvIUuCf7Ze
2lNW8k3DX90DDMEgjeQptDoIC1SH5uHPhj8Yrj8kkLM4MXABdIQcoAKFr8rmExLZ
jSmdiJ2cXUTqud9xbdlgPSddtzve6JRpjpP4LmQfr7RhWaMAXa5RJPaxdZIL5ZZC
B4XFI+q17LDDaj2CS/x1Fitww/qMsSNJ1fxOXFQO+w4oUjOs8oWqbmDA9kFCQOPV
/tAA5zJ61V38TxfmN6yvCQVISaRa2lJWCeKlc2ADFS9LivIACRJ4/Z8VcQNMRYH0
aWpYoKbOLyYSr5HcFpIJtUgN6sfYfKIQ7g124PBsYMHbn1yK/XVzWEraw5AWFUX8
FVgKx7z5vZH9+245qGdH2905CRgV0o58K9DVFIe436FSDLFzYhatD+f64yaO+FJ4
xXxrLgjxZ0D/BNnGW//yogLIKlTPBiP+x/X/YVqMhq+pvFOUqBhLnkBADxJBNAfr
RoLU0358paG2khZqJgbEAqhIaiulGN19cgSNODV8MIdklnXSrXgVCEqb7Jz/dSsV
1L352ZIqO18M+w7csUJEESRfzFMW80lvUD9WE8RZm+ZRss7Z0eGQrLtOY7td790O
88XtRi6PKWBa7xw8OUe6Ru10aOj4BALUbBFQv0byoCktgnm9547q4NzuVfWotyL4
yuJQH8Lh7sC3aIWEGPveo0MTfttA52MR8KVsDz9nTuqZWjW/J2Nv+OtOZcFd6mML
9/eHcd4H2E+mbiWuS+HNaQ0Oy1OZ0jX/z7eXUmEyLIhay971fqfhdoyXgSbPEj4k
rfAFEHMQZOnN1yN3ggJnEH795NMpKTZMMEyUoO0Drg2y6VinCkMXccZoeOcfbaa+
x6ww/yfIF62bR/APjfTbj3t7j5f4mIb6GUgCPn4ONyPwPFTgEgXoBOn/cwRUKAQl
UsT67B2lwCAbCaPk5UwktcvXAyWEhnvwlR2KmMqBWlIp9xzsuADSauz82kUxvuIh
Tz6VvBAZbDBUxnR2s4lzehEeU6Hz1KV2V1jXuMub5WR7loqRctmc5P4FMxhz0BLj
mMkx3/H2PhGKZxc6ACcNHGXOfvyy6UmTfSg58GxqDChKJxn7ZLgZolToDgwI6oYI
tg3bg6LkpmApnIgLdtJnNJu29TZkbk0BC3BBvoRFtnSqTUO5wtqvI5DMj8kzAX49
WkMwVLGD/qA1BODFm2jznaejjk8Znw8gK4+UVmpGiWkRoYhl1tmfdZ2CIecjqoy5
4qQVYAajv+47HVVcFOResixI8JSOGsWTLj3oz1MBJJ/dCDyqDuTVv4d2sGL+jged
mKTP+hVHpEU1Mic5JHIN07uZOcWJcxPF3fC8+nwHf+Yq98902F/0JXhrTaRAcBoK
XYytMSL9hPo+lXdcvX5Auyp9vE2p+qtjwFpvDLn8IrDx/4dvBeetV2jncuT6jP40
HnI9PyK13z8M7QJTS5CYOx1E6H8NVbz+j9qxZCHCP3vyA90bKTmSjZzYCERcosMg
aLZOXHK+EdB6L5jaO/QA5fE/0AY+pIGc5GqBB4QnSrhrbKuWydV4mW7e/DD148fY
pOvwakPqQf0lrNeKOwX/NxLKXwpgPpkJeT16fDyX9DknUW5vV4YKqNIxez7DME48
K/S5asAbpoViTdeEF1TsbRStanouBMZQm9PGdlLBTnf8lXEAEltiTvaYCfZ9Nyx5
RBsiVhFwRNSAAOWojMKJtvrAz8Y8QuFjunE52XTxYBdEiTn7FZieU6MFbC+Qrfb4
qgVF+R2Hr/O55JKURsiHcmWBSfprJAb+2kEBIb/dnPJf6XzJnH8otJJ9W9VIn2nf
1qNG+7TVwrH3K+vE/DBSv02Mnq9g9PzVyawOgxEqaGv16QHdBnBxmImlOTDyS3eF
lLGYs1jq9ahWJEw822gm2KlMY7SCd580Qm8UXhn3FNvkWysPNS7qSMjgGhmc1ept
5crasZZb+pgV0Sse3RrGTPsRG9Bm7q8Eo5MMO/ZTC2BKxUZfaHe/JbG2FjdcaynC
hR2JMOqASp0UM3OIi3BwpTzFau7b3y7VVk55+3upJnBqHBnpt+QfErBxR/iLhEnT
T7YIPz3VweeB/x8SE7h49b7Q5lGugDfkZhcg4EG+tPNMWlz/yg62USwWxzfCIQpi
1krJz1ZJOcy3+1jakNOcpa7frN+qfmgHTFHvNCBekrfOoO5Q2/R44UJpHenkVJFC
8GcpwW0Cg6syLKY7UhLCmZNqgN8bpOlGZTTVIa0h686WXURFWe8N7AgFIaQ57wgX
lhxYeLPY9fvyQsHYCwbsZrjYvh78THgGo16/Cawsa128FdkoOvk/mitmnME31NK3
YcQqq4BJH5UQjixkasJJ3ILqCBppsnCYxqmIFWf/iDQxOLJo3NLgTy8Jw0pwKiok
oHQBATqlLA2iDGaA2sEMuVSo9vA8b+woY364x2/dhdtIveSQxNPgMWKwzXMeD/Ys
YHYL/zQ8hYDVCs7HnF8qPnZEeCASLAGr0C0JlKQIEjcEMWTlah8xSKo82yMGJ+bB
23qqpxYC5R/rBhMUl30y/T6bKPjJgvoHK4CZjME38Kd3NGuYl3C6rGOzDZDy2+37
nVKlEUf1lNkWUZmJ2VDrQakO+tJGtL+5kVO7pMocs8g3p7bgidK7U/3R05jrL0w5
Ja/wb0HHaExKX3UrAHDr5/1XqVIh58+H4rp6OZIlNbM4NOicG0DZ33EZvIRrsJaA
wAwfZ9iZb64E67sB2zBGZS/LmezypdaVKXmjWKNzeB1QVigifq/9wx76DqCaHj11
jOWXf1WBrpxgHTkAruovJhsMicVZ97o7E+8QOmHp9YvFkRZOiPCnjRtNJCpu/NB9
y5QwjifBVtJIuerKudR6UUt8wSfb0q24/xyZAjVkSKIxHLem5NH5ZU9sGiZ4vfnq
STlnekzLC5q3vMEH6yVD4buHPcX/GeMo73eNeruwVUFIcRqgCC4sVt62io6zBMZu
RWcHeT6tMky2E993ortuHI1kEz/6CjaxR8DvBQf2Wu7ggNox6zIMlBawxROsPo6m
mKEcWY40nmY2OLzzmyGx3EoIe+toYSoXCLyKJJrqT9p8Mq8oZfRok7Y+zO8fSSe1
bmjd9KSyThplTA2TML1Mwm5iokLrl8knOhzlsBlNXKN0SUh3rDhKRWPirh7bv02W
GoErbaKOLoAYo7SMg198JsLE6VBUS4rHAIBFlDsbydFu64LJgZwgmC7kHEOimTzZ
i9d3wMj7afK+Aogf6IVqEDx0AycNei0xa7uNB5Jc7qaZu6+OEr8t9WkfMC8+fnst
U2XNJXs5FEX2dVNvfJcEfcnDAeTEZjs6/vuG8l8GIVjwDJ46YDsxolYc8IKkaRlu
1XLuhAGkd8Tkjz5s6u8RK/CnpY3MX8gqUKRZAIzstw4yeEPa6BgrNmVSrXOO/LhH
msD4pAjoeHjRf6zy7UgUKDB50GSVhi0aQOMQbO5YEuZ4GnZTR6iFOEj7yltjYIB0
tOgICt7KUcVVcgH3lJHKHvpQGEu1Zu5P4RQLEfmFCZ8c6RxcJIKBMPp7DmOa6kNB
DWR/DSH1dtuAgjjS9N7ULplPC8QAK0tljAUA1KF8QlOcMXv/zCjxywiD1GAihyAK
dY1gx7j5qADCUSBbrBN8De9heNTCr2s4/oReizThTtL1d6a7KxeGD7OG9u3xirZn
LteYiEd7n5vvoPsr4jIYuHXfoe5P0aRupVcoNG2a/J/OQ3uFX/+YfFiOapIoge3Y
o+5ns4BWxgP2gHY1V6/1zHyKMUXlSvaLiPj6rSgL8ULx5t/h50gCzliysJAkoKyP
8hKJ9lRW0lK2PUyrAty/4NZVt5G6hEO4m95eGsttcx+PUOlyp6EkJb2mPrQNCAGa
/35+8ZRIojzJZVMzL4ABM6DmVKtFiOX/oL+Pq3J22k7b2uV3ugXwC6+tpKjb40nt
cpEYvd0VhZKa1nHIq9KTJUui3Uf7GAZahg06EB9HJiQY44kPawMFUxfNj1qAX6w/
3WwyylpRV9kP0xcoWNWkpC89ukZHvp8v+j9noRA7oS+tOeoShTCgwY6Y2wYsz3kv
/IERw4J27Ck/7mRRgBVSHmsdLVZFS2TCXxHYJqG7hcPJVSm81zgrpn3EH3yBr+W+
ZlEPwUPr99na+w70FsAmFWif52rlKMCNtqPOYmXkDsNpstMPf72YkKagOBjgHwVZ
kDYHpbqVdebL/YUx8W0mYxUoHl36ZNFr/SiN0KjJt7up++SQU3quLOVKbYVmo7K2
RW+au2afbVrUNpl+Snq9Xfibxjc4ri0wMWWzJl1KzBfAM9lyauTB2akO4tQBaQmF
6wtYtIuZZ10N+7rP+/B3J/ycb8nRsziqCSjMJ8aMUR1IJ3yiXSYjXfjOdSd/7m24
w86wjiTKi7UcDoEKw8WdbB32L34adBHZR2DZzHCoM8ascOO66ksuFfdFlthIB/SP
7S4K87IrNgsQNxAFPFcWlDxNhxstodR/30MUF09CX6E/F3fdyn+An19oLgtBZhxU
uhIVhidXddVBEED52a7S9vjOxAymUD97N0X/Vi0pKz4PA7cdMma2mwAcITogrCnV
Rwg+VCxB7FV2uA6fnbjOvbdzHjYp9CbuiGO8N+dn1x42FFgeoEJO0zTpJfxC/k5u
X2+Z/OrRzn3HnmufQnqY8F2o1TrdeAfWO/ImxXfKPV+hiKFBWuzb6Vqaq9/jnm2m
C0G1eUyVQKk5L0dWX6OizP2ZU9DLXOf0SmNO2VVCgfAWZvm3W8EnRzu0LTi7bEO7
zPqzlnwgmVkwp20yN07pYL+dNKAu88lozH8bsmIB/JPx2sj8GI08VHrvxKkJ6pT4
XiJiq9tk6MFMBsHye7Spa9Vyi+SL7qUY8tYsfFQGUpCFqhkreZnDS8OeXMpdrPaR
XXt1CdveZIILzvD5OFUTexkJYP2jhsQczOUIt7FZEMbdU7DPHIhXfXF3aO/3F8mk
6qR66WUshY4sm+OdlZv/fIQqGuqnK6GOm1a0rD/WzFxWX3UV3TVglm7gFFL/t/Xb
AhN6+1GbFasRMF+ooUTU3gHnNewJuAe3TcrU73ltBBXA6cvuXDWdimh2+mRnVoGY
disquXCzTB0xCUERJvK8WR8In47Zz+JF3S2mITLggptAVJ0aQYOH9YRBpXGsvzYn
hjbtdbGgQBo9Gi3r/fepHIrMtvwaBM2Na4yJePzIx6jOFP8fUL4GNc3E7zMy3CuR
cUnc+lrLMaryLMUAzVW4zFNmwjBDIJwSkNrK+LQTPwDtyGfqelbGslOaUVGLQgUX
yOvc5/p92Rrt1KfFXFq71CnRNfvnBRO99o3KgigiaPbAwIrKyi7F4U8VxOloHlDF
dS39ZAeh6nX58X0UKZqfJWd/E0omkJyhMHX8tNwYXOQhgnr7cQ2szniiL+/nGmdj
fiHpZt8X0cbiFVF47wqrE9gXazbFRgeXV32EL+J04lc5KNpO9ZVJP/06V/fTA6iK
PZBclQ2sbf2RpLA/IB29TDABXb6HENs1tgu9J0kpYPrSOOk+0lTGtUoD0o9sfYpR
7f53HCPRz+0dkAXar6kZRYgnBarV78omNWz2284fxE59Vnb2t+x3xzjAwBQNHkCa
6i/jP65Xk3Eij0bjA25MFbVvrXW1wgjYRMBsi67++Rrw2vWR3LXFGbAaXvxLZTMI
fABTlo2zkCFx9lrxk6kH0BwykqAaShr3SezU+C3L4QEKvpifQCOoCBhnm2WvJMKQ
taz0K+2oEw9yNgwvHcoENVksGrmxmSlTDuN55HUYIC+pm1XRiHHVCHmQt2xCoXBW
TAFBWZebCPvnIMXFyumV7HKv+cZpOrwIeNuyt1aNTLQVraH5G51GpnWlUj+7c+N5
6kYDQcXmgjDGG8Uad2Ct+8ZxQrZSz6hoiNNYGmQHC9B/yKO02kSjdM5BMqBW5zz2
u0AiYTkkIVH1YZfX7o2ORudB3TA4ewv0NynvSTOG2/JSatfPEJE0J8Vs/aB3a8hE
VN3nAYCyEZMtrkgQmShqb1AtmVOBXoRBthPn9+puMxpGZARFUji0MpmjarrsnFVV
hG33NScfN9BW8XvKE31y5P1NDfpE5j95VnQTD2Eq2NbMmkOBqfO9+IrwNGLB7fSf
mGrsuzxs2vfYBnueN6q2ulmoywJ37XRFpVZMquPjOcqjehBmmC+nV/FTznDXZpdu
3eIlP1hQEsWi5p/mmDmC6AIOCniXy9ZXieOiii4rqqqei9Arg+1ngMyI0cQCZZ8R
jYsmppm+arEFz7M5y8j4MZov4fnRMJ/Bcb99j4sbaufIOC4eSQi6MMorCJOpOmbE
HGdn5kESFXE9akMotNPJGwALAEMXZNJ4PUCTMb6qzCeECoo5dM34sSMn0wo6D0VK
f8ZqscVqIXm3UxeymJWJuEtDVakWPfPryJ2g0jMK63kbl+vqH9e8A4iO5fvvS89X
mz6zuamXH+fTnHP5SWRe+/1GGcP9RydzIKDxk4MKFqJso7tgzGAJ6Bq5A8kdHp1O
Ojo2B1Ij2CUNKAmPgNuoz/3A8bQlYMOU4LRgWNFpR2ix7OFGfG/LPRjPE7fIcjzX
dmy29SCVlB2V3PgOIrVgw8VxZINR5XUniLjFaIimUguOikI+nikv+0FT+9DvVbTe
cWsmhArtYnbp2X7mvYE+lmHh8AkF9NnZFT4GORN9YvdpP1cFBmTlHcrDqY3j8EFe
u4uTHZ0HqVkFz3O4HhNbIHXM57KN74M2qSIWOTeMZwWRIQIZMhrSPALvpXEDbNFp
D0zTRXDxwWRo1o7xnZ47pz3ADr3IJqr5pWuH05ZO69+TAqT4pvp+gcKKAwcZXgok
yAbYoDY8fvt5AxT0uNvL0u8EBRi+YnbwcavNUmtRQSWL4nUgTMIH06dQYcPrDkN6
xFyq8G2cD8hlSFlIpH1cY9UCO+8c9eQS+KXG9mZKEbsxv49g4fA/HDhgTJ7jPtu0
cS74uFcOkuR6DTg0vxYFtHawdrMxzBZaVWPsTjx4IzcgLppTQd7RtWF920naxr0a
44U3kGlw70Qqn/1M/xPdWdzV0UjKKbrDzLy47FJCFrLNBKj88gWBWAJCWQz+YhLV
cP8dQW7xA+R1N8AFfep+VcwJQYLzhJ8mNRTHejZMq+cbq9RW5OLzIZJgA/8lZwWT
w9LTZ6gNccwr4rPxGkPAqqU+Sv3eX1HYyj4ng72Oay9FR6Y0QxFDKAn8TSdFq0d4
c1G6Yjus92ShfVvWcV2J75Ow8Ng3whp3ULCVag3x9d5T+v6F62+zik07/0ozkGTk
OnxvI2YVKr3LzI74w54Wc3TNa/kliINFnATnCCEcRRuzsyVvZn2ZS3qfkZ15HVzW
EWa9rTFk0mHNG69f/+QFkwy8LpZygnYl3Aek2HDQPz8aDpOQ9oDhFPpbgIuKIRIc
K2vOGXHeS+O/x8vRgP/0WkNzsOUgXCzaVYDiCihTbhYy8fVkrdPneiEM6zp0JBkT
e0r8cn4GPxkupo0cP+vML5Kc4dZxpcHttzkklB/395qPD5gHnOIrxi1ywl/i2P2Q
jR3X6e3CyDSvYgL9EhibQ3Kx86ri4XeWlxv+8gOYdKaSOtpd8fnvXcIWHoUUDKjq
ytj/T8Gl5Wd8X+PTnaSC2TGRlEFDyWkzeFlTtVCsHHKD4HFEX3fWWRTDktkOtS9P
IrzOU3sDCAV0hbD2ewR9uqHfPDFUZSebLSl+nqMeLL5BO4NdosN2MM0F4F49rFTQ
IzXIQZASAeE9Ux2Q3lDFwPIYoqCLC+cmTjKi4dfRski79befKEq1xpg+p9HqDUuI
uaqZZoVHf1uBu9AS+2TUB+Ze4jX46Yaz6xBWIHhw2x8GcQMioLrQ5i/FYLMMsm6z
JYtfX4YRtU0CLUmR7WVcz+sskagUP2UAXYAEKVf+s6jBFhLfK1LpXfe46zwDGBcm
HQwKQ145xhKnSEvp3HaEAsZnmIS14bevj4uQB6O6wv6is69rQL79CXs+4+feOeY6
1JY1nQtO9p+TL+MMXMhKi4GWMu7atn+QTIH49sCSTwBgzTjLbGqqAv0f4ntyRceX
nAEwGaNSuAQ6I9eVuXnyoS65LxMj93kcziEbMtZ2KUMiGPm99I0IOL5mCvV7qqW/
ECv/g/ichTjHm629v9admMaEUWDLqusNlOr+45/q3HjqfzUJ7Q4Kf1uoWSAV32KI
RVFOz9HIglvUCyF7Q191GriMP3Cy6avQzHT3izSacr1Sj4sJJgXeCCdLQataWo/s
xADzJwhGNXml08709BjGUJYQfsJgk7CcGLAW1d7LsQlHxzdIYEAuvOVOBYIxb9rI
74iPJQjqTkdUm9eoTPP1uuQeZe/9IFUD90AImb3iR8g0CRm5WutP3F0u/gQSN4qN
3ChKs8mqnqcNyGepnY9qzOvmNUvN09+YyYrRF5YC9UxN263k/Ndj2ABNnqrOzvvE
5+FFjHgrQ/7r8r6VVu8XW7N9wHk9qa9nJOutX9maQGw6pjVnXIfIecsB3YLHh3Cc
`pragma protect end_protected
