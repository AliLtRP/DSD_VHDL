// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
K0JDltjsoOdEJ0tBUUmvof7OTkbh+lRmcerLacPfhoO4jM+y8BA5/WS7O8PXhBDR1CdLjNxbUi16
nb/H2oy6zzzgd4AO0y51JXgnFAExcd60EqVY1GiHMRr+okDthW+IF5YOUm+zHFWeVvVTJ4QBoMug
hM4ALXNVl4WtBJR6Ns9uLxDkM8lS1zK+8gcaf6/kcuGuaoMEHK3N77CeQXk6XHy5OkQgbJQv7zwW
76a9scKMVxMTZqW9uJffvnBlF7arWKb5wE2in0rBlt//Cz2vVqQ3EZaq7f+bw8gI9TDGeRhGH5nm
zmwSs+0w/X63EN/j8gNIqnPli2AL12XjyQpEUA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
iK2IZb3MIqeB2o/S+xE5XufZVKXap9lQVL8Svm3sQzYX39ruyiLUbCftk9XudFVGq2d3Ro+s2/mx
0dbqmXeS0g1AaFEQg0SGRoh4b94vJMtembEm9HvPTof8uihA3t7ECbbumNdZWhpUIkYmyRGs2iXd
xYA0uZ9JXH2gebhodnliFiOiwkh5uMqlArC9B4HikXZnIQVnvGSThpQtS2ldrfYT/887Pd91A07y
j+DHguFGhSu4nINtsXiyejlUxsYeR2DZVc1IXUbNa6Th7wQdRc/w8cHhjlI9PrW28K8qExmNvBOB
PEMv2q86VSs2+cFhvBVKiZtzAtJbZvxZBNQYPNnzxaP/11M3a5FusJcdGyaLGKUydA1WtRljSauM
ijakUCT4vCBCGwU4Kqk3fW2Gx7WjOOqIYugi4AeITgj/TYxr5/P+fk0WoaNUWlV3f8Zjl8yC9lk/
ZkmaQhM8Mg1qRYKJlu2XjZIX7qa7AKKEFgzhFsDstljUwRBqTULv8R45sq1MJs68O7M1Vis4ZZNo
p133Zb/sANGHPJRAQe27HOvuun9bQEGStYuSXSGQq46hGUaoIf33usESBSu+glq0Xtn9M56t0Shm
LoU9xt13ecEA+SCRDEi4nn8COIyEiU4tFRrjJuPG2UYGwpICBmlifgEjTC5JRwLnnrAfZ41UJJi6
IG7anQxglOQUbb01gOlKnTO8Uxg6CP75CQJpRMD+4SBzm2m0RK0FobfZnF9foLq5l5zmASwwUsnx
fB3Yf/QhBLzk2FCv9bndLCOlrUqzPGBOZhGzkmCKy0FY6yBdjnyWe/u0X7DPgR1duslKA/zgmr3S
YHin3TSnKLmafKS3sjBmGgbjS5ZvYazFvf9F+6iv7tOrz13LIh1peqNum3pb+T6cKobpCZK8MKOt
9j6KI0vU6ki/mYqTKcf3ZDhq5WAd9wBMypRDb4HwBBGR55YYN4vIgyLFqRoad7iaFHGSVe4idg+2
Di9wg1N3jswvZRAT4RGNyrinv/vwm+ysnuEu6IcVYcLJwmcKx2/NCazXqtejuprLVdNlUdXws1h1
RGdIo5hq2Pamv5Hh6fNIEvggh1p/3b88UT0yX1LaKwcPi3BM5VLQjuoEQREuJ6IE0xV4sCK2NmI6
ps5IBg9VQBEBtrv4fo1Vkcrh4GYYWDeL5BVhW18fWNyBJ0vmND1aXIDpzSsBrMAmS+nK/zk2O+Fj
gIBpUL7I8llx7Pl10hk2ABWRBHrkQ4vLgeN4dhO6YDYd0RYTWH782eMK+B4yBZt2/a1SAHyZ6Mvu
6AKJIIohHDKOviBx0+hcjJShRjW0wF8uC//U8idGhfYAm68jR8XxDbjFqpMm0ja1z1VJLIdLa+gv
ZvX/FfQKmRODdyVar2PdDrvcaDfaZYZ1ABdyBfQPWPfxVz/pDl1r9I7cnKTAO0FqhGoXZtGuzDdS
x6TiaymDcCxfqvnoQ3j3qajnCNxqDZmk1mLoW4VB9xycSiljT6vtfgzk1uYeOITKocdU/Zhcoznt
UuQ9Kx1I/Jb/EXNSTuTJjF7wj6Gmg2Du7kRX8zznPPo65EHREigkztPmAe6tsiurdN/vbG09giJk
DE+3T1PCZ6mYi/BkYKcQoXs2CoRAK59m+W6+uwZ0a1/X4q8lmpavyadTtMVug1c7S36f8PMkDswW
bHQcfKzO/fRe7PEkWebzts5T0CGsWu4zPryWWGpozWKhB5QANPTUjkARAc579vVroLF+xXFXANJ5
VZraInSSvgaZArOJVND0mHDtE7llRVLk7yoQZ9Me7yHpZrnvf6H/8ESifES7hnU63CrAfahhosQv
q4ol/Azm0KY4ibkE+7bX+pLmVIvWgxiGcQ4uPcRUqbfRmRvOFHsIG7/TqLlVfzQL+g5D+NhP4P3o
MdlrXIo3mHf/ilnwD1gKrL0hfaEi11XPW0Z1N3Z5QMsJwA2suxEhQuzVkS06zcNRRQlJx4MvH2mm
SecNm40MCc0n7DwEHyrt8o+sK7EuI/NJ7IzArWL9E0X5Y/03hY+yQwAzMVWrxwSNMm0W3bQ3/VeI
HusVe5FQyx8boASlLiBclCuvXdPZgfwn0i2X6xbC+o4SJ3MW0x7QkPEJ/iXJaTGXO5hpC5HNH3+Y
MV0Q7HfzsWpkh315khcUj+hAU6Z2X/65w4/NgXg8AdqgeU+aDW+Yzu14RqTH+ISV1hFHC/J5mzg1
Tiv3+PF/D2UTBN27MhgrTiZodKgEzXJS7X+mBFrILizl6mwkGQQZvvP+2JdnxgMOc0uag1iFkM0t
XGkRLCA59RcIaWSeGimj2/k5oAI8qwykIrfzqOJZSEPVIpe07cWKWLg/SToC4wphoWZTnFb8NLny
uqN+HUKXvMIWLyzFQ/etRtWAwpaG2k4gVemp3J1a8845r7gFmsAx+ZSvhT9F4h4rpnQD9GFYCdaa
lOWxy01S052ByfsCMNyK05IXQmlB6kftptviPTOtxERijy6mLd/uy2hXq1BAxiMARD4jqmv5W6Ms
NtXBIMqW+Jxt7CgG+p1leV4L684WO2VMiP5PmzD9AtDuPXqyzxkHav/VHSkJDZB9LsuzbW6N0FKh
rhf5kGHGNYfDwITbLzk6XNJJ2PNmLEJZohmIQur4ssDZmO/HmyXRDefLeMpKInAIAfT93OKUQENR
RZpWznwJkHc3K4O8GMI9f+vU/ERjaFaJ/jMPvLCK29MJaJ+FPA7F3cQKv2e9976cfbY89xOxhT8X
8C3g77bhSAqWydfS1M4NDuKrvP9/8wEV6aqI3OWf3Vmpmzb9/zoT/UYxf6XwGUVOE7BzSatfMC03
uv+C7GhsMgGwVZqlIDRT7Of25bH8SS5QJ4KbKfr1Q6U9oMBV7XoYG+BZNicGoJeVv/ur7pVMZcyF
gHdvFj9DQ3VZZp8rsGdMF9P0VFUpdhDLPgmmw9dh1qzQZfdSRBfsxGooNpBa+dOBcz84gybwlAhp
O7/4QIVmvu7EHae/hqZpgCkc5yrqsQsb8M8oj/k3+aLjxD2c8m1tCGyN3TU3knA7WZ+PytA/4SHT
PFw7/wwZP1ihWGQ6WRS8RHO1Nk7FXMpzACpvYgm3CbH7IWuvmBIbeeQEOlsGGzrOy3ZXucNS4eeh
XR2i+EoeMBuRvdiyrck2Lps8OR2gRmkOSV9IWqBnVOrINvaFemUQb2ZwrgusWZu889///q57iyVL
Kz/M4DPwNEpMMgIEnmQ6q1jWqmmB6qzWxUVEE8gdbB04Fh+fpyngDSuV8woWcRiJUOUnHacCXgPF
fNbz2kx0DXoSNMLhNPwiKgwS7JNqPDB8IWiaB1xfy01n6a446AYhjpAZRBwCPp/qmARgQUdn4KIY
Q/hTJGsamwiZx8w6d8j4+/DbXg6MUHnZKKlZv8nzCXlqowQJbfv5K2mEzWb7Kh8cey7SexBRBvVD
YQ4IGAHeZe+hTnfd/x2B6rypiUjXjP3a8cqb9ilNS4Ox3eyCIKFJYxQwzyIDx5jVFlOWQAPZnME7
YbrwYk+dlAmVGyAyKGKoy0BGCX+THIVJ6LPep45BVdz8iXT/Cu4YYUb/uYOAWEEWw6VRyr18kRBw
wjhGPWaI6i9yiD6k2pspPxJLErrVeYvDuLoscc4GvgJLVThvHackxf2PtySOnG8/5t1vgj3KEzHT
+tdWHRNBxr/sKRC6qhzFjJp6cJygnQcqd+XTZTKFpgOO8CcTJIY3YYocR8r0jbW3Hw3YxKJBwNxv
u0MHLSSA748R1jOzijC5elowgpTky4R/Q11cgnPujQb491RWW/ScTk0U7xsASk/WgvMFFKLWzk4s
3CLu7Ll2IQb7xDVNnzi81fQA5Ivnsuw20P0UR4/TrNRo+AQOPqkdLeIk0HfadYFnKHwgQXuq24fB
JMe4agn4h3LnySwg9OkgMXe/pwjRq6p2UBbDJghyAv5E5pgJ9EQ8mQWXgVwZrJen4rPUcaeBBBys
dCAhp8hAHD5GwoUw+CbKfIzcOYPco77S4kDqtRUBHJEvqpvOMzyCT3WlCG3YQTlV+QjZFnKoDmjZ
uLExI1ehy0lPHnibqHAWulkPbx8hEO3kpdEDAUFfKd/pvBz5lhdvDOD7jJIVjbWYrwQ/qognofnM
yzwNVLFtOb73EQnJOpuEGc2PfwlEJUUpHHMFssCSnuCkXxetW2oB4K54IBQHiTlL9OyfSC+yj6i3
lslOAAUv0znJrFtkKgAAre6qt55YEjGiN7I+M8CH1PW5PN3gasoJ7sKnpIF8fg2sKRmBYWCQ/p0O
ogU6c4Uqhe5Fn2FxrlWwNvWZ2ZPTuemxjHN9OGh8NbkpWFv3WjeLcwO+KdHiasECuUFpFGHBeNlm
R/+13PcwBZ5OAstogSeQD4dFJXZ0IGNFGzr95M5exEeOHqBdM6zh8jzDANzrb614Z/Areq6u5EpO
L7uhZ9IshxT38tUMCzuf47qmYEwTx/JyYXa0+KsiBH0eH6njEfp6U81I5NjemSCXe7Td9r4sKe1L
5uDzs1w5Cdor47aUPi78+JJC3BqD/6Pj50xExWTpKvzSA7J5G6k5oH+gMw3w1mh/EE4dbITP9yIF
nnS86W8/sTMDtcZi7TD6FDREyIYK6Mo8g6oAA0C2wbnHImOu77XH34uNZOs9O67QBOpilNCulqG8
nzYuWJVmmgPz5xDQtEBDt+TjZQory1qHS4meEEmQT4FywzS3uMut7veMvoGvs/bNnV+O7tg01cKn
wz33m57h8CmJ5mSR7mrgc7B12Mipg9y7aH/hGH3UsJBTclAYqm7l2b13Z7eEKMU5Zib7VxPH9FZ9
IOtAQtU0L0dpHSjBZpw2LkENh3qOeCfV/c5UYlTZr2+7tnPdvmc9zOkxexBTQ1i6kpWILyi0H5vq
WUI6BLaetcES4iaNGEInMaOF2uj4WcrjMq+t3JBEWMoDbvU4PDDlGFZKPgZ+UpUeLePSWC5gFzwS
P74n0nfRbRHCKoLQlz+TzNC+YujrLPRu1APkW+5j+ZSJrmBTk5c6VhcFe3tF8FNfmyTJRtOMm/tz
+Yemj8XOKNiec+iAvV/0+c6s1ZltDLRDUUuhMrOO3il9ggPGow1GxIR4zxqZccZUGSvPC5WLIIwd
UX5WSPfglMg5sY0C/NtrnnliUIpWLFBg+JQsvsIGJj9GDguGO/jbmmampcJWyx+VYjiZegzZhg2S
8Gt6RRArD5UZXE4iUU05MWB0nZhzZLGukPEFEvG+tTG5gD/q4VbKA9IovMHKVmIK3qAnjwpG+i/8
kepX+ju8p9TCiS20kFDIHJoAdlEF61YY3Igt2m6ASMOOKvpzzzntYJLbm6amIfZSF9pQ58TGbXfq
7zM0J/oLpgyTKxheSjtrFCSbCK2T/Fygt/G8VvaNiCg3+sXJeOW3E+qsaknOtIF7wyz0yjuupXzC
HZMpb0kSFQjIRlXAfWT+4Z7Zjv+9IGIsEKnyw4XyaDANvwVrzdc1l5+KX6ZCbuaiL3acwxgCrm8J
gVFKas/UPU6vjVR295a1LoEX+nNi3p017Z1ogk1VE/Qz536irGHccI1FsJW2YzUcZq4xLYr2Pw5x
IKGlSEBrSvy4FM4sirRCiyIE4eXcCMheyG01O1zRpDTxSFsODozs4DjKfbYwpOwlCtEe9NnfkUGb
sl5sP4XAv5GN16imlsLAUg7HObhenxqjGsu+s8uxh4HIdA4hIsMxxoYaVDpEtc+GdFnPdZadVmxF
woxhR3jLtbH8FjZ3PdXwhwsGSHaAtWkwgfOKqCSEP2nTKY0iolDu4fqtcxfoO5sHJ515B9Q2RPuQ
jzFEURiVwb2gf7WaGh11wYHvn65fZRTOeYhSEIjDgDK2ja9aL7UfQDwl6CGBr5pBmwSHTOegDwtD
767bf/kaJvyXGIq/3ysovWJoiHFEcMyurdECXcFTd+TekIL0+nf10NId0O6KJJJeB1Ir0dKs6TBx
fFUW6QGnYGDYbcvMy1KeBu1vS1U4duj2EUMQeo8myrmq+5EeohPlnU9c7TG/BQ8up4iz/gKD+fBA
OITWHzNnciaJ8VMZ0T8Nf2BzRX/i5IoCoFJ8t1Sp16K5FWjgeAMeikUY1oYTCPmQXwgvQoXbnBZv
OhCc59HpvRgrYvOi22qAUyJasODtnPhkBngSycBtCFA+7SdOnDvXcYPG8D1D7t6cxZtHzDLR1GWh
4DW34MzdHd/4EfeeEWU4FotDv+ca/CZodU+JtFVvS0Qh/oaub05Tcb/kMwT12UN/ZjNfmehHtoLw
mHtRIfD/GT2Wig1aIordZXL3xuxEhaGphxbBxrMJYRv65YyafcSiso6OdWCbcYaNq36xHOTaa5O9
7DiGzCrutYryhJleV3jlSwCW5xwlDC+od7gGcmBEvKNr4OncVu/mRozQhZOTRit+zFst8c6Q93+0
vT/bHZJMF8Aq27/lCKZIMuBbqJBYrzu3AWWXXvWkb4d+qR0TjL6YHWik0Rcn7o9eEY8mnWMeDlS0
yZ8b0CKepgkF+JwKm1TsbzuUmnAPw2Edr2D3bThBKi0rXC9C8fJVP3VBThYuF6FgoYDLpaPPif9q
u+zNg0zXNb5JfdNoVtKOfysttlvBX30lTfONQtES9FZKjhjz1FfsQyoEEvRKl3m9s+sfi2cYKP8M
m9of4dcyR1I9tChtVUeQ7FGtVaByiFeU+WoKfps0AmKLNFK6ccsjB+v/73EI/qrVkqosQggOvZNq
NNGwN9al8jjhaJwh5PcnSIKmA46c/v9PrF4GveOzSOVnNarM9sv416DOZwTKvYDr/sFhaXAlHNX2
F7bDS8IkitYdCXLs5vArQCL003iYFzuz47SAPpuGNr664xMlT3otuFZinDEs9EK+dTPy4kNInoMZ
lRZ8secCAaWdIijnpukoO6KYgunTIRDpY9WpAjknwPqS/r645v6swv3ZQXwKLH3366iQ13pM/EjQ
reGNS5DYPQIxI+Uno/SR7kyRxqbnyo7MHj0VeGRGAHR85afltWPNU+bJbvMQgBrc9K9BWuNLuGSq
DSiu5xt8rbBEhAvHwLIaKtdCzQXKQFxpVpMslkkzY53Wl9eP65vHr/pB9zXxanChEzqoQpgwXVeP
JyXwZihYG9RQyVkJRzcyY97dcQJvMDnr1qpMjmj0Mt2LOVhhGEx8GfMqUE8H9SJ0oIPcLSb3fPfD
pxhTXlWJqgB4FOW1mzldOHWnQVdBqAsIoMyRdFUn2bhKENaZv7IhJvKEYjBfhiBNWABiO5sD4AUh
JH0yj8bVnW0l56QHmIaa+E63qg3hlo/SYNTrjWiGXL8atjMWeyD46XdwL3PfndU3fOyy9UAe9Bbz
qLwiyabpb44i8rlf2wQD1gC4HaQu1yO7WRGLRU4kzG3dAUE/B9/GqOCzd6tU/NujHT/+eRFDBobO
9GdhPLvXgyqS2REPB3LhBzU2PYasuqlBgK6wPtfpISChvBDDWzvCy3hujp0LqFOOgvJwqetI0l1u
6P1qFw7c5MNm14PxTDjqZV6OaYPB3uYHRDZb3GlUnjTmiuFPxwKACEam7oy68L9QGBGQceWwWYue
pIrhI9nhFp+pOeFbFAMsOd7/L43DrtISjAtRCRVpnUUBQufj/hY4sO9j89EKuBqncSO/qpWLGJ8d
/XmEO9OBEEDPYf5C8oeWeNsJUuPXLnczXxME83fOZWZZlXM8uMJ1masT1rlmPEWot9xJEmMSIuoM
q/FMXle8gRfp8GnzE0a+lBOrBmjtqckPOyKdekJaJU5YNCIWaN/rLI604cNHncWCwX/u/UZkzVRD
GzIaJs+BHEvYOsTxOBcYTvIpX/VXaFerKEU3ARnVI7uyP7P0D7oWk2aOT3guMzW9fyrL8uBs45aI
V0OxO1FQnDrv8Y9sF3plH10KS3r/rpsNRQTJPySrvSEFcyo4xlsqgKIATdchmRyqasYm7wpYUuiZ
04lBxgOw+CcsDBIhSEDPp6JfiIwnUVl/b7xxO16p5x20AK5V4mg6zoaVaHiP4yTeRguYWLIzusMP
Ple2lZRUNZB32xOMmhxqVVGqDEbVHbCs1G9Vl44PnpwDUOyIZezITeXwl6qJoov5JvErdGru5cRz
oKpLKCfmerXmiqJS21nw6udQnQJf1Q927hAHoCHNBGpS8nPkdfnh2lY/0qQWpGSnA8t/Y74oEdJC
VpLy3Lpo1Hx9Y6W5XwsvocEmuHEMenDmbCnFhazv9EDaOizVo6AxYKdWcSryT93BqToko3QFGjcB
gcaFnfs5wHeZsN08t0wogaG8MQ1hiT595UkmQJSOmWgfMPqAju7vkfgJ1MR/YJbbQXFm69XHGwLK
8YkSs8rtf43/wwRhLLk472dcxemEEVX+2NOQNkwd4KX3ozI76mKYUk/wZEmuF/Rb8hXLN5vsUCxb
tN+3+pXbHPhpsleFNieXDaupqwsvqHAaAbnFF43O3emqyjaFZ1R9eLfYbbVUR3VSHa4FsgxBHfN3
zJmHMPzp59rvEpLgPUkA4c4WhpkcJYwjTQPjwUKhpJDJmvnDzUM2VwWh9XASHIDcoVwzHl75iqRt
c+jPxpq81JnRYv23PXAdpFd/D3hNclDLom6pT09P5vpC1bXqrLyulCIGnGFaTdQM1J+KUL+lks23
X05fKRUIj1ZOAlrOPiQ3aWcgSXzve04SwUE21qT6MvDIGJxqcRap9ATo7SGVA9mJwgLw+sRSkPQA
OIoZPEoGmGuiDns3VmIHoDjHdZ3ksGxNsGHCZbG/OITNKk9b/z2RhO7KMrma0vLC2bAR+Onc7++W
e1NU3lKVtE2LSHXh5d4aMs8NQvSALgyah3pzBYVp5TPVhAhwrecdfyw9eGTyIwj0hilawH1DsneW
hztNgoZbXejfsMjh1qMu8mm0Z9hTdyzsYHS8yJUWAJ7MYK9kGizgqqmFC+8iMPZ6ZBNuNO6rxarS
mZCd1BRN4islJr3W9lYa2KB8TNVcnC0+tsIltUA2N/KiEmbtsoGYVztjU4Tc52w+tB+tADPeFzrX
WgkhRcx9YZtGs79pgLn2+h69wNOYjX5k8aIMlhYGIpVaR7K3aNNKtmdrgCg8q5FC02iXtHO+h2sY
P0Wd/OvYkg6n/MtWItenXI7hVzUNGHt8/nsE5BuyAlfh8CdTpdJKydZeJuzuqM6NWV90rdKuA/lA
2x0sQwxSlh+zE4Di63Jn6QOuuJMk6YZgddEAmL374Yq+iWB9qvnH14zVXeS69uCu5UfOacT1XpB5
qbL6LWXYCYKNX5IZr0R70cYBZ6ApQiXtpuc8fLtUUdobTrmJShsBU5ey7rEvJJefp5QcmWTq2xXQ
TSurtyV34La+gKu0qEXdth2ncK3M6+A77ShoDmkJjaZ5goa4sAy7cdZH+rVp9YNhLna0vB18LLR0
3ZI8bFLyV16RWopGDkSOpo67hJnYBKjvOe2AL7Qpcn06muSm/JYUJcNRPEP40cTSu8mdWxEd21K0
ELCnvbV/MxcoyjLklnXeUpzVk8cjblhzoy3Bg3djowrYqG29cw8aJHZ3ONjsszzO3ro7Bu2PwiA1
HnT+spZJ0vIFHvT9I0A1zm9NH4z1PeCif/ypKyjmax9PqMfANoFX2DfBNI3r3q/Bi3rHhiLUAzo+
/hI/q4Ok5G3HOc5jUiV4RDd1rA/ooXpr6dQswefbR06M9Ino+OpfNH6ZfYO7dIyj4Ik/sI4BmARx
iqKitypBSY9V89I4R81MtF57WAQ+Y3FMscsnp7tG8kZRAY3Rw86xwmKMsVi71UMPSQYg8OmxypNz
YNnc43QJWUcCLtH+EU6CkZwNh8/JAH2KqBN04MHCbQDhhwlySVIkQVr+KYjR5VskdGWCWibY0pNI
XwNjP7mBTrbQ+XJD9zG1OcL5EKM4lURqr1jZC0GzIv0h47MiKU6FgJCIRiCUul046GYTsCJ56MH7
pbffXalBpNOJg4Hhr+dYrAuQj9nZKv9Vg8E8E1wgZZl9qiRHbca0vwriW+kBjzqH6dh5uCow4a7t
mdq2XZJ5z578doMm6hgDgNulmjDMukyoMrsf+H5EII4LjDnllVFr5XlxxA+ytsQltMWCpqhw2OVo
cPJaLE9rrnsLiIQvUQv2MOAlR8h5LqBK+KgpsDwwTybk3iVHCH3Mrzp6UsQ8onS+ZT1Nn4FddiJa
bCVFIXpUsXmzR2K7YyI5WAshFmm9HigK0OscrvmWphQK9G3FyEq6WZqLJFToRz0C1s2XvvT8iGo3
AdGdzJIF4l/fe6c0HN+E7D1v1SwTfieO5vllHGhfRM8hJbUnb7WIwR9HWKJrUBPL98NXcJSBwO/3
NGqSyBPrYftl4hsuXHv2XCSoLupSQM69dVjZyJQd2SL/6VjepuE3eUyjZ+hbJBSn5+BaFCVEMQYs
IfROOQ2NpehX3QzrHE3hEPh9Lob4pdiWr1PXe2tj2Oiupuoz990lv9KX4unFQHAiLI0V0RaoSOkE
z2TGtvNOG1WgSODLOARLJ9iVK/1lOI63wqghzIvBio20Eia/Xg+9W+dbEpgPn+bV3q4OTX8OiOJz
g3nPzcwzo8eDAVhRm6T6dRUC3wg2kTCbOzdSKjiukelYUF0b0INbzGE7M/ljhinG1l5Pcfzbf+Kf
ptcVdobTWraFncyf5ytDyvjQsgQyhMAZN0KBjUcdI6krW/n0Cnun3ySkTY6e2pOJty9b1AY5RA0Q
NMX9mxx16fxHnrUPubmGphmseWMTIn8u1EwygLNoj3EyjCgYaBUYLbqA2KilER1n7RhmGNRbapaX
0D2d5Uo8hVEQxYy8a7cFpN3qg33+q+OSdyybK1ZYWMbKG1VbW+WsCyZrPYjWUWSnWVKoFvTCI9rG
mM8e9iKfkVfK03ZIds0LWWcZwySU5RY3FJrkS+6qjqnkwwmdb/ztFS81LFHOcgd/s0mPYze0K3Xl
eQYP+DNYVcg1JZ47zLybWux1fqEreZjnfWNqQZ1frj9l3VIoGKYdBoqSb2+FsUnAUzs4JeQFYUwp
WLgo/58HAIeoBTr4ynZLS/Yc1MdBmdmGxv8A2WNc9TrYKcYFFaumSCMX7pZcsCAtI/LrXwTEz+rz
H0V4oSl9zaAR12+m28NGVmGh+IcYfKgxO4Va6bi2haLypHUXnNXp9fpmss4gEH7b52s4OeyUeS09
+QoF9udTszwez9XyYKpAPPucnPSUCKg0MI59cH9wECqrXYGXgdX+e6NZbtu/B3PM3dE/nITE1KPf
5thEtqBbjaOuEpeP6DEHReDv2Y7QIJoFh8lVqsYnxeOT3BI0UOql6h5LVXflYeL0iL1ezhiv2rCr
1qUOblhA0h7FSv1xeXC+M296OmOiJWhxXMt+BUmXYkcAcz6aZ9laAP+ntK0PFWJ4+cK98OskQiec
Vi2zAWd052v6FWQWzIWfbo4/KAuHnV88gMF7HxGV3ObxtNknUvG0g6+TBAeAia3Qtv3dHZKlgQOI
dtbc0G+93eE6orpkurw3pHWoF96aYnNbqXz+VlL9Eek/J7fQasXg1m4CDyR0J0WZ4DJ65m4Ks4+y
7OE8JcHOIpXe+bPnEM5/Shs7pUcPd3edCHK+F9/UxzM+oNQgMOonBdFpFHw/nmIadaQErAEVye4D
7UExWjGuYYFDQdIjolLWOw+JxmCvWQeOHzPt6oTmC2nGpyTRYWpHBkmQCMTON9dzoHJeCenPX9tv
dJGeJhKnafb4FN5gTjK8ZNHJjXI5sUO8poBho+kVttL37xzy65wg9ku2BBdJR1Gx0Sk0mtlEU40G
561ItiUnb5BUMx+FTpwtdQwvaWdAuxH5aQxTPbG2LZICGnZW3a78vEZ+eVqm20rY53Coy9IDbmKz
bJyYzj4Er8bDHzO/B41vdIPVgJrqoQBPUlZLC9vGHK5tXae6uUAlSzPzmidBaKN7YcCIgaHFrIJ4
YDWoKujbq8lhYCXfyiQko2K65aCj+JJ3f+0wb2B7JsS/7VfmxAJlHYIy8tr5VIwz0DTZr/WCydHb
TzZ4hF3R2VENTNsgwmEVyMtSBVCC5MFsd2m0STJzJL8p9c4i5qgHxsF2HYSdaUt/YuBRH7xJGx9R
xQ5bzY0IiMaThwhLo7a9ZpqrnUxEe+YB6rdmIobUcTjcg4PXBYcWqzdE4KkprqKCBXj/xfHxZthV
x6KTNjfsy9hCzYW92k1ykcJDLUeFT/8q5opNnhKZBwJrSif1+yeSsxRoA/LRM6YBfBDSYO7+dx14
woyJ2PRxyzqXQjdl41rcssJIAN99F5oU6l/3ySEeMtnTmk879x/rKrwCJo9S/yEPAxPf5vSL+Zwk
nRzvBD6OwkvkAC9snwrLysScEKcwiNGbHn1kgGLQOn96SjSWdcA1JLiX9I8z4qa/OQTMb/TKEk4o
ITmKNtdteBcv7tx0tCZh5pnDkTreqqNf9KTChc3YobJ8vf+EHzfLBCQZfbyPEfozy/Y5pVpH/XTl
MF9AwdgFkJIQfuHSxZSU1KwNZPR2Yy26hMSHTpi5wSraejx7eAtpwJTpg8G7vjIGgyYQqhfuyWox
KHiga+hQlk68eiMVGrjjUhmXRTwzz17IpQ5Ygf00NHuRVQ6eoikGN/ME+3BfVYk7ZscoEGzW161A
G5Cq4rgdo/PW1QlNTvtjpt/GKEE02pHa7v/0wykQBMHwIF9WWXqUM/XLHcsDEKIeX2twKvxY4GqD
7s16BhAmwDvrDCyk+R6AbmfCt9FGppWXB0IZGmXuwbKWd0Dl+akfIaxmt0YSgxDhQkJRjkXPHe25
yka5sdC+ntsExtaBpJV5D4Lk1pXFDoijTTKr7lAUaHKtZorF69yjp7U6C5HTWKYl9TQwvHsI71tj
/BXAHCa3YTMQqcI/sFdf/c/IK7cNYvGmU9e6tOJNRDjqijdlUFKVOdiSwlC25O5bObsB/tMCf4L2
HdVjdb8TKv+n+ZzjVCDrZ4YbeVxR0fRXOQx+gU+hl7lUxSc6WNJyu4oYc4yvzhYo0Fu4A710GFPE
VeBcndlunBTCiwFkJqUzq5dEFFvaoyRnvrP2lw/idPldq+2AWh8lSXlfbPeLQZ6uaIx1cTFtlwue
zcUwfVNd5FuHT9MlJnF/z1Lv2tW4nBKKwncrCeDACs/n2BTu+tWmqvcoW1eWw5LhMkYT05fm0ADc
ciP4sj27HtLV2Jcp0bqZIhbqoviEqXZmwatorodZQLOv+1Fe7kq5ts3A+WlXhZY9N8pukNqCsTP4
5mI8fBPQzxuZFu/Ulb5y3WJyWPsXAmkgwvevtj1soWmllAhg4fRhawATZTvpWiDGpyeagywyTZVb
CMecDpi1ELVRRGf1FJExRzDyv6qu1w7vR+9W8UNKVX60FdhtRjj9p157ejIaG4FU4+bcI3Z8iok4
jgiN8EiNNt/40Af6R19vv8tu15mngTs2nZYNYoqRTzLOHUDgRg402XfzhxsX78xWiQIPJ8hiPeTp
xv8kX/UqMYGnZM3Fx8/iJMHHvwRZp7JL5FRPgCN58huf4EjP3ikV1+UcfYcf6lENNhzHpHYlaXDu
gnVWSFHi9093zbQpDkdXlJnoEhFF3hF7QwBjPkSk3f1ghH9YFiOzfxPg8+byy5NkhWdxVyEeGIeB
KJpmSg1Xa2pXihBaSN27A8/F0mRjserDHLGMwMxnv8x6NofZ0Go1Y1/Kk4lmHp3ETTaP8oFCEI2Y
WH4dWmDu/5nZc9Ply9YOfimkeKlNF6m0dsLJh7FYqdcCY2Xiu+t8bOFV0qhKrLFFTE8iihQOTUAF
x0IaCLZE1NwlLowVXNKXvgB7VNhVrvzVMGSqCmmTT5zKDHu2hSj9JprAggFKuVHKNfldLd4AYE2r
5Nn2U2nKDDJN180EiTH6qZHIBPyYrCAHQ5DiikF4RPrtwD3NwB9jYUUmoyh1X+LDV702tms2XAfo
s1tEf5G8tdSU4etnj99EkJxz0q3VqASC5D0cf2M3SPcFAjySJQtIGxcD6a2sfeeG8gf9bKx3xVl3
Qi6n8jbo69o4oN18e2IocA5P6cU7+e1xUvY3JaC9oBTnpchQTDGsTBrA0obhU0zQS6Xgk2Dzdy9c
fkbQe4OynOy2p2Tq/qKnJ/Ep5ScUaX4ehc/DFdkY7O3bhaD2UvXovdAcNMJjoyQISr6W3iTTtact
Tx6SObGp6HgbQwBOfQlxAMUZqIEGyGPcmwa2n+qB5Ga/sX/TLn4vqGWBpD1bc9fBjIEmt8mFOXiA
qK+6HMg1q2rOj3nzWTlknTxcfXTiVhxszegUlFEWvYVnVlzi0/SBwH2XydhIihTp49+2QtglTzF1
BDOj62CelqERUYDg7ZYjDCL95k7o8sT5e1h3WSOLuGMths5FAbzR4Fd3tjuTRz/jdEvA8Pd2Y99X
6Ud5tSMVMfAsq9ene17t18CE6+fcaZTlQj8ZTtK0zipJI72w9yjVuDDLZ7mnrs2oQsBMXMQykzcg
iwN/mMPxagpgWdzwy3GLW7b+amTRAIlPQsOOfogCR3P7owO6gxI1EZvDvpICMNDgdk7Ub//Shpth
V6tcFPLMmbqjjZ81QDnBD8J3oIrRQMoIDiPgi2YzeB5/trdSQfutclAND/AFRPmRd/aF/FifAFpK
CrH5I267rGRsXgHPq4/Qqa2sPWWWYiRiqVb2qEkCXvvBhAcH7jYTqcjHRS0tFeZrHfbjHPDJZYdy
5d9EA/fgtPXr+QeMd8DSOHBOakrhJTer78mkRK0ru9XpnXXuJe/yp03V73lkaDFRdvbVZNIjc4yk
aDk9u3utsX/kF3P3Md/K81EDfvKMTctWFKmoQwvTcFQDCU+OWDWnx118spUAYTOmls//jfL1xrmA
SU1UKrFEfZZfwIqLcbZMO+LRiFs0jKoFKoEqZwgZ8DeYzVXM5GnK8RED1SRtZ2WfX2NLxF6uIBA3
yZyVqUBLeuNxRChzHOwWHI3atTKnN4fGjkh7LO8xfezp2lvbbOnAfmUa7v3Gpj/6bhJocqsqF90o
AdxUtmqeYf/p3uzWR2ejVyxm8aeHoGE6NFj6pvDEZeztzdPAinjK+w8rpmhphaoIm+3dEboDihQZ
wEH2mlW6W7mIWMemGTaDu6/Ll8o82LX2i2Q8TpDm23Q2FLC+hYiVGqwgjkLQS7K7TAvTO/f6YA85
Y2uNa8mqf/YiqeBuawPRo12YRKK5gd7RwfprQaPXWk5rBc+axJtWr6gKHmhB2QH8wl1MM5PXWvUW
Zl8XacGo+Md17sJR5rJCNWh1vlz1vqKGULlicP3lTJIeStdd6nqz8DMjYh/dlaf/igyHX9TtHPu0
OD0va+rMemxGp8QyXUtvA9Di7yIf7RnwO0CYeNHY2KZDWhsK1xLIkwm82XzJ2vOxsTweO2WWoomN
xbSM2fBY5iNy6Fb+1a/fpSeyvZH0Kx7Fhqn6ERYBZkbVp/5YSdXBXCxh73vXZZYvWkXLwQr3NJDg
Hak280/MJdry2vz/m60sUIXek9YRC4BrDLhkwOz2DLNrFj6cs9ENBBiNElftPzPqrFVNv1cwHgN6
R9DmsiaafxuMnswvbfr2QR/ZISxLN/iLj1Dxs/Shm+lv03pbRBlPTflsqab/kT4tYRR5Sv8kEI0z
kTRcDicV5otHRDktaK4kopbyXj1X08/6y5g2k26idyy/cOnOPVSPsbWnzEWjxv3aVkaT2+/bldxd
4aHSAzJD3SBpm4+lNM07Ffrl34ZNDD134kTmLUFG//8epShGRDhKIrJdNizSPluKnjX+6lQ7Yq1c
bQBrpJ6+Yi2yphArfRoQqrwayTVYJuwrIDXg8v4k+WhdfkeJc3+GUR3UZI29TEOkEElLlYcVFVcN
fdP3nfyG6YjrLhPUtx1wtAT+TCVJzA2WiBy3PrnDYRzvWUZycg6/LKV7F1hkFMgRNcNVnSI7OJJk
kM7CziclFSrXIvJOiasEBNd+OLSlfbbp64WOFwZk2bvdwAOoM2yozR4OlV2kXK+wFVOuLk9JYlcL
NaSvVqM7l9o/UJYErTmCSdlzLJZ1NKEQuzrna5+dWsLV/UHGn0SuAPlDk/JN5F8m+ng7nSkuTZyD
+UwKBW5Mfx+SeKbp9g/tl1CL15Pue+2MtUFK8gPex5tNWeDnrPIzgRDglTgwBRqmajvKuuxBJL04
jOoLhOPSFzkP5TTqCKwT2GNkMahTPZ0SNiLHPuy2o8qRY3Wj3xPnmfsjJGTeHYCc7uJ74En++m6x
FZglgxdeLlw2yG9LHJ5TipRQlQozYM5/00NEt1dgSqqgHDXTyK4Gitgffg9+FQqvtp1SyETGyc4R
EknXxltfLtU9GoBWiKCklQ4qPo95hn0laGSxF+uiTZU5d36C9avrXc5PHSPtn//k31XE+kLSS8xs
rtNA/gsTV7cfBNpwnvLC930T4/7qYrRANTszY3CJNS7Qy5ZkpeET5nkqOw+4uo6LOS1ZTYj9x++C
69jS06K7ZDty7MlkFCzPtZLxZYupIbUArcYm6FnVoP1EhjhHtIydSLU6uT/jlAb6EHSQNsxLfASF
OzKZk3PSINGaPO1VzqZF6hzw8dMdreRrBLjgpprLDligLvF0ruQy0NXxHiBriclf1UuxC49ODb1g
Ggtr/saG9g4/dSLVQJ6t/45VEJ59y3Vip1hqSNTxg7UBduGlkL78hhB12NcGFqAmwS8HLZmXmz7h
Fd1W98YMAW4Pe8urvQsPHL/eSptUUU9H1TxDvAFoUsx2sxiadqj1Qq4KQWRNPpuTq4ns/ffgc5X+
cIhfDR35eJvCc1eGEQmvrk9s8MtUUW4GTNZPdrSvZGKsVMWaRfQfEwK5+Q3SNDl1rdqgA+kB92Jh
m/F/NdIPRCc5xxxyojxFrjP9KmpR+U5lyKuI7Yao2f2wf11+u3kc2jJmUpjfve6B+i+cDEgsnIIg
2jmE6dK+tACq+KA3aaccwhnYA98Pdk9eOYFqZed4m0+Pob8N/iIOxOQAD8ek8VlcevTrNjR84Dv/
syo5xEZvlyzOk/F/cjGfaTYBFej0yEQWMYoLbXgN4w0xfPR5qjucAl2xLhzvVATj2g/1tZUfpMO+
GDoKjpZ5qBIOjUdErkKE4UK6reyYWH073wLeJ2Cut1AVJGYe4ojfVFdsNBCNuE4UxReYmrBD3F8L
r/YGI3TQwPpVxHyg3bqf4b0PjMdeRQ77i4Je/2QzldgymdWcq0rDhOgwRxbsD4UlXfsmUuH6BAxT
gxi3gf7vaf5RvUaR07l7seArP5Cx+KG+UFNt6o03+2nTxBo1jOl6mvjBtn94XrZKz2xnpK+5/XeR
QcQ5aTJkAr/9h8YfxdltNN3Z08bfY1kUmF59mbdfrx7xM+z0j1y7op3IM6Sh8QBNY0KU7/AyJ5Hp
2X4d9u1ydQUICggjskZUKxoxCMp7z9SrPuY/PzFBzNBS55MVY78FChMsNLMLDYjCirNqeByARfAF
shOZYBEcYuej3Jq/iimZRLuTUAq3j7cimM/IiuWaYozI24mJ4wcNg5jEyvAtodmwls8QAO7TDx5G
iMSIpXNqiEjroetSnEVhPqi2BVXRzybpebeCtRCAbTovhQmJb+BSTCuc880LfFs9UnldO3wUm47c
7pdM/d43jH0/R75XqK9PAmJOgrv2rF/kWSOZ69CP6jZhRk1vpBdEZGR24ZW9coTgc+jz9ikUshIX
gZ18sN8YovqJy2JC6KKuzSGW8dWiJrA+oOzXw9079GppP+9UIoM4DRvXPfIwxlMw2uIK9CVO0T1l
0W10a2r4OJzzpf4uFLiFv528fWnjP1JGBvg+hkRnoqW+LfmBst/1va6k8IVT/7nlKVsfT9KKiINa
zgdpJuO4SPsDd+yaDBp4ncVwsngxiOJt6wAy4BSIaV3KpV7Mskokk9SP0tZCL1UtRV5RvpJyXgBa
Tfo5lTrf6kxL62TmNqi4gehqOF9mhJ4g4YxfN1VnY1Mb+1d5qBHMEWJme8VrgBjKIDRSJ9xcPe4r
XwZIdRxe7FAKWh93ImTDwNJk+xIWSLGP0e5xpNvobzlK5IYgwb1h1P2zFJLkJIBWd/j9XA1jwA9X
twW2QIAYXbHeMCRxpIUjLAF3/E/hOSi425GFhYkFIU3cmPZF06tBTVpsCEZM47FDP44Yn0zCfthd
Ggq3pu5rb8Zzy+EWD0Q+zZuFJi0XkGfuSTQHzKcCobur9vkC2Q85BcjVM4REKQyp0XLoHKd7/mLU
qSfWL52YfupgS3Q68jbsv83iMY+KJmOLMsvJvG01G7RcW/6m5+dx25T1AQNY6ZD0MLY49eEdVFFs
crau7v2wdNFa9kZzhjXEtbdMI6WI57NuKi/MA8L8qejZnbHpgOX0EhS+0O1sKKNrllbaDLenMoTq
7Q/395MBWBizdAROxA2hLvxLQjbglQYLbc4hEpX22jFhlxAfHVXTllEZF45DxegFZag3RTL62/EG
IVKS5rQh6sF5PcGm4dkEIumvU2ajCZ7IrSPs3AhUt54HXGzH/NO5mxg0XpAcEcRp84hzygnTtS7e
tiDmBTfGeE0szzdGkgJ0bQ9LS5Mc5frvmg0SZCto8eXpNZnO3z950ZZ35bf5fwqSlhfMXB1sCeok
h0eOezVWCjudCfh19sJSduCiy3riV6iSWIqaVBTSNun75o6GR5GNSVItCNbaAC+N3cojvAkWIO+5
IZeAKZt0+wso79gWC1E7kw6v4u9rPwXChmqeNrxjqUF1byjHruexrLommEbHc8v3TsAdKNJjhQSs
yhiplZtbKloa2/eZNLlg/yiY7iNE5P0B3x7SLBtpwsCY2Q3ZoofnpvEwUDBdBlHliU6TWy5UMYIE
oLOQ/RBg8TJ8jY8sI+JeMLIGAFBhXWBvCrtBD8Gu1riT/1zBE940fApA6D5e+PHU5VYnjof6Z7d9
eW0pL7K1KGOglvfTO6t47BLRVXuNYt6D8j2BZibCggAftOmZijmysU7qswLRZGcf3wfkywupVL+d
iC53S7x5k2uMQhMdpqhm3PXKuHEbHqcaq77OO0jToUGp5/rkiFZgy422hhcQIFMcZ2TePYq7PBen
BfVfclwRDcHkZICzody1gm1lXKRctycaatnKxbvGNJ+0wVR02iiWJOIbtagDvdsPcIXzhoG70sqE
LRSIZ3/hKVdb4X8a5KJzSRq6dx+p2ZTV6g/AHi2HuHXcuw0TZyhSTOR0bTv0o/nUmggPUDuXwQhL
6+9iMHcCr1D9CIDzmMxaRRuDXG1lG06sjU02KtXALXffu9B1xVw46C1ciM6Wit/rGuCcG0XJzIlm
8ltYy6iRLS+rJ+mk00qq86/3O/sr7OeMzKjc7p3tF+36b0K3QrnGg0LA6+Z4CRKwwE6mfOTQNOfV
CTXSLpPIZ1YPpsxHBs6Jf69jsmuiwnEagn3G8/7RxBkGwqSccFJ6Rhy9TmNdu5cMeL/33sxJqjPB
L2AH4wLcapn5s0LqYzCPg+L/4tBhYmn/jOO3Uro8EITdSr8UEZw13rr0jFlGhMKqNxn8lbOSqXg7
o+cRRUMsOd2pD2nfUQIyHBL+kzcCsbYbhL5uCHRJx5PRnAaw3i0BjYwXXkmPeoK2zRfkYPgTcYep
AZtV4dmDZ6z+3xgFAwIhd70bexE8P2TDCAxjtumnG5UUM5nAcrKGiX3/NJwd5XzupPxavYqDkRAk
8HpV6YpvM/nuAf8AzhzXQcieTZdEFp1mNIEiE83biC/wl2pk9yKtcJLKBZZVx6OKjFvMqsVhC2Gy
6qBSRnV35GQG/t9cduA4LVlC2gU4hG6fyZtD1UOu4UKqmDA8e9zNwKGyqkWbCC9+a1EVRCCAxKC5
KhRcrI7fCiNzG7JJt2DrPqBQ8mMZcJaqfB4IKHIPBtRGslyik6HbIU83UcOTV9/B4JR8swUHDC+b
T+n25R30SmAqm3VEYLoWsvnalOLBzTyLXpUjZfo86mYBHqRFCUPe2dwCbatR2o8E7KAs7sICIW24
btseuqRkVnaJWvVKmLGZLvZSFMv8NkDtaOan/2LRoTBZrVq9Ifm9Odgziz6PpGlZA9FZq4+fo9lN
e1iQ/WOCzWpEOr3/uHp852crUizg9XurXfmKMH0eucIK88dDndOVerMz/scqB14wUrpEnwtOeE1I
tfekw46RQB2T+DKEz6NQtukR47ELYjSI+B4hjIqvtHXbnJzswXqPgGP4eP4vkBUopZXF2Bg1pUdK
lPSTkzEjVAuFks+rE7uy+09FO8GF1rprFkdnk7g8DhNvKiQAZjncS+tdAIB38r4qg4uSNYfd/SPT
4iNZszWSUGtRNa6qOR9S5yGWH17ihLacJjtHLZ0rQNqR9sDs0GHdcRVpHQ0grdv122L+VM0LamUm
KrY5CM7s03U0klYsE9Tv7+KNFRZ/xfIhWdPMy62D/roInxs8QyHFrxNjP+udQo5Fz/QkyKovFFHp
1mAKcwsL8kO2isuIaK4AXNpprzc5TsUcRYDJ5XEk4bX5vHvL7cb0LDFYLVQ4g47Pzj/+u2NqKfA8
h+b2B4scgF+xWv1BSeIs4Dil8Ljc3rSVO0WrZ0XrZPuqctwEDhkuYriCH7Iljj+413iauO3EjwAY
eqduxM62LjyUK7LPimG7oStJ/8SB02/NmyyuBVDgWl5HSklDxmeaSLdGTs4KhBYQTJr8ihRlvlkX
PT+B06qXGwcz08gtCpdRiVIPOCAaucojkS6gJoMaOcUFCd8ZcEKhdGP1Zgrj+KC7TOU/3Whsteh8
N/FHtbeh8avJme8ine//lPgokTgeMHKAlsp1xQ91JfcE0wKUIPYCIKlWRdeaukBolN43MPBCEUmv
Hu9n4k5mH7P4aa5S7AfKfRlEKfntOwL8fDBv5KvXK84dZg/0orPspU0fkIiezTBzWwKDpVPkFI/M
KhCgCr+wT3opMaaxJtuxMSrNhXo2frabXlzWM12MV300tcxZgxUjqTm+xqsL2Fv2EZom+IvXM/pJ
qHZPq/JItVM9CXh1XnYA42xYThzqrNetLLo9gAF4jI8sRoiVKLHvNXmqIDpjnm7mK6qFY415kLeF
5+i1t49NxkeDLkdqaWIRN8hczgTyws1NBZEFiI2hTKTsPHGgRNsohsYw8NyepITimYCdX12w8KQj
GCcnEO+Jj1rjKmYasV+6CB+cKBHxuClhDAg1/3wCOS/Zgbk5x+rn2gpB68lpzB5FWFTnB/iQFwDQ
ScpXXRbEt20/Kn0o/76FN/XgwSNoa6j02jkwmTiBz0nxvRmQjSncY6251JRH/TmQkDm/SLehSXZv
XEGUIswwpGPBnZCQLWRLF4anFN9gIN2cXqP776M+TPjiSYq5VGADb7/QxVxbqz69Q1xooMCGqiz8
IoZMei09b5EPOlErov91cAck4nX+MhGGoeJ2cTg6mqDewSFFlJwODK/kuk5QDfEo8t0kMCYO0tuM
aq5lVJ/oHgxnwehIQ2cV9VScka+vrAxIOgX2w+ndsmriuDd7EzFJ06QWsls2noeFh8tbBla2kAIm
YfmxabbMkEUwhOO1Sv95QuwMVVtoYZGX+ZC2CNHlAFE6Y6CKnpCM2Fs3lz1KBMX5h6uwaqBYHEo2
0jh852Crpxftc3ZfpqruHQu/7EyKLHuuSbf3EWH5F3z0aIxxBmktQPjI+eF8WYezFeXAT8lPXSob
OvcEshPXDClZgUCoMtNmmXTmNcAd+5ryxLk+AFNlkOx6WwUWyw511VoOqdZZQULzq5Ctd6xUDIxd
pKPciDGFa0Pu5KIa6eJHnpPOR1Zf2LLlf+Cp2jZQgvaAifugogfUGtyOqwzltSN/zGb8mEc7rzmu
1PS42K6pZLv2Lnv375ZCfFm606Br6c1CGx2iuPbKkajmfLTmeNe26ve35H3nlf5fVj7OoaUzUdDi
vZFiweORR+ExGgi6t46WNlrGUzTvZm88zQW0XI6w22c1uYV3fp39/PRoP2+oOV0BOPCQHFgKsYd1
64w1cYPKZNOvGLfOnXKEGbcwi+dfSY7wxkPbf/JwmVg5+kX2hnabXE2pifAfz3XRLz3jaQNKynRn
FH9jrEPBI+ZMsEQ5CNOB+LXRgHlISZIDq6ibhUdfy3JrlFMu21LZyFtryZtmTqS8N6agDgAxTcBU
GEdyTIiBHrlxEZHc8P8712ybyOERutoXR+fivFqrzaaar7/orT1VLO9DPwTFxT5p1K3YTK5u92Oc
WwH07p56f7TgWk+4aoBMarYfZoVnYe4hPMgOmV19tmTSDGbrZCYZ7UqztrSq7EiytMxpl6Z6qiOJ
JNUQPvAF7XbX+DMKZUOCBACnZpTbT7HdkCkG0PCsCm5nvgHU0h0iTHj0FxcQPQHqJvs7WOA0mzN/
gX+nMe9hW5hZzwh8nmCx8CrVKG4vLKcvGz4fbsAcCP/w3XXFYeORcPwh9rrzXJ03HTm5iLq791KI
Yf/W+fLowkDq20hVm7SCxshOW/2v7T9/no7Xqa4N2N3yk/DXEAisH1Z+7gXPStVyS4zIq2sy3/Li
Va5zMgmNE+jIVoFP+ETzHxNW9H/hRLnxs60fTrnaj2FvdsqsXH0VCaljdZyCOZyglPSMSE1HkgEY
eoN+nlW6NgF8STa2ObOV5P5w5AJaqU6eeB+PXWhhV/Mr3xCFB3koz5sU1FDJcyJ7687W+wuTMSO9
EEvwa9UzmSUpLNYgkCXR3MpXUzktaFIBVKhNWfkbkxdItTeOQwosHjUq7v4MO0clw3Zif8bugfxD
BNYN9xoaOoPmtmvIYjqu/WgelFPFeXaddNRFicOwGEje3QYGwUpQzmSrNGQgh7Qbzd22v7Nd2nvu
ShpnlE5Kgb/m9aXTNmSvKiwGlIjMKUCPj1/By0/k/UwO0Sw8kYnqytGaYWM3Y8BMqLsZkrgWN3Bu
4hl0bFJm9sKWnXliWW7T3WPIO3IgG1NEg2Unf2KeNu2rabi0+h6BpQ11a/tXEcM/jF/Qdnvpx4rh
DLBBjdVKo/ythsMaVEtDoWdwCiUYE63A8bYMC8UQ7u8RgQkbSb3OXHoKtxRvKkAUgMk2/ulIR9Dj
zfRojFHWsUaJn1jyJ/TfHSEpsoEhXNZglgSuhrvHMJHIpP4ScQipnL6j9vll7gCpbsyIdmfw/g0F
X04+Dc2fKfdkuHyVWMRaE0gxg1YflRlfZOCdZErkshpfvvhbWX8/xwJPNTkuh4I+zrRqCHJnvYBx
QaV5MW6h/v6VVAbmk/amy1yq4FXNUupgfdTKK7W5uwQ10TXflgicF9syNHsgR+hij/EY0dotwzjW
QA3Pj1t2rFazXt4A4CS9QHvXm272lv3aytcrUL76sKvQaNFcPWfoFx4D18ZZY+DR3uwfeq04Wzj0
sEeEjLOZTkkOhIQcCzEatcz6k9wppGg6iPkhnLY+PzPi2xaoCmOiAb18JsUe1mmt/wTR343bwW4u
X/LUIsIqseKOT+v3Z3lJqawOijEZNcb5A5zYRLLIv81FxDvwirmYuaK1+GaHOv5OucSl1CWfXSWf
WypuW2s/Ywz4uvlUscCEcwyuU+ZuQ37vAL2SqYe4oXp4pxXC6tpUET5tsqhEZMi7AUA49t941xmr
Gd1BsYFjADKnCHm7O+RFhz0LbhlPWVYK++YeLVy9rCraCam9BaM3Kumpgcotpnkvh7z6mB+59xl3
EXJVHgyc2qdcjs57f7+j/qiwTqiahZCeA5yWY7EQDUMXro2BddX28xLjf9TkxJVjQxfFWCrHwOiA
rJ5Lp3cT6wJ0a7jHUWlv53dZR1cTPnnwJbe5jteaimq8PxMktckcsKAmmKUvL3sq0sVCUAAX8BEG
+TdIcuFO3thGKqWfu1MW4HnANH9YiGbZdG9jICx2c/M8GsZOdDOIjkW4fJa6rrMWMV84nvlCEdF3
WB79xtl8xFevQM6eGUuI15s+IxgEMSLvBhXwvYhP/1lgxVa6Fhv/QGuoxIC5dImb8QXV1ywlPQzi
VCCV5VSWUNj2b8nNl0UFG4zIaVZABWmbjVSW/la41G4ARSixpPQacEwDq7jZHee00R3ZSlkdYTqg
AonKBmlbwXMfWYZLuFJBK+prrWwEvdtTh3AjQkvdJ+2EgkwlrwNAUANvW+UMP35uhDDOIRR82KCz
X6XaGB7qmuB3DMZcYHiRQCQdGBwIGMkYd+151Pxml1lcawbkYKQ1bK94+R+VqtudX40AHQOIlsPA
7VxPertXdkqb5+SFneBo1XqQerFboBB7rJR1Pio7WpGnCS7txDgeZuoqlWnnpl0FEk7xjijEnbOw
mZI+TWRvHzRffy268y/+LHpjyuzpKVCTrSHfgSQbROqGv5g9TLFZxSZ3l9uuVginEErXDxr//q78
xGjSsTqehbDdgcLnxPyj3nquJtbOn2r9AucveRizO4Kp15rGKw8y6moKyqFopIlfGouIjMIa1ceo
gVq0UPoqQlWadfyFwe9SW1KeJeGlFaBcEEwjdZHjf9T8IWOkzUy0KnDbSeaIYX9Lm366wPrwZRHz
BDGanE2gLvJKHZ0E5ZcZoYNhm2RF7G8WMtArzmFPLoI9UEGbw5p8TY07LApmwZFbfMQfxjlughF7
rV/QHGrOOdgpjOiLlnw9L7jXQGkOL5+wcbLeET8geVX5MIOmlfU/772gt32tjRs1Fb1/JvGdwADc
USl5dOm5aHPXhoerBLxFiku+YKMVP6T0kLqapVdt/Z4tqcvCWBqsZ7hXz19YQLY5sZRQjFyACAkl
3VkT91a2v7aL7rcGkRgenzJy/NaibvkB/uO+0a5fcljPlSwLpYSKSg/wgMqGeJ/2kWXLAEmDdgY6
cOWH0N43w8UMuK7jXAgTD/hr+CiLDnuAATpps/ULvuYeMenZMK+Ltkz3h1nltDnsq3+yS4va4dqI
R6Yiw8p4N8cRbB27PbZePMtp02MpG41QXiedrHvnI3H/2wxYjoboZ/oXutH/8NrvaJbhkNoSO06U
92SF3KgBxoiraP6hC5IE6inNPA1iFXEjVOH20iKUrT0QIcdaQ5pVEZgMCviQVZcQWuGhz9d3dBuA
nCqo/tXDpXwPGVvW0Chey3GAplQP7Tpo2ln+fd2OYv6sfdQszuOi22EcdTrcqWdZ44Cr4ex2LOSN
OFCKtCCXMQ/11yOiNPsDpMguH6oALTTknar93buTZ+by6bicFMCx16pqP49FZecsYPI0nzQoLYGV
kNxR1kFC5R3YB2E9FQnBYjXOvDHe4qsCUcl9hO4ovX2luAeH2rGy08vnrLWkaSkFr0jeE28UFD93
AtvESKGHibTSer+F9G59eqIvvxg0vJ6qLDwO3mTpEYTgcPIghb0xamTk7O4r8FOG+1Sf6ZbSNSzJ
2r3WxzG+N3Lp8CI32JG7TK9KeUr5N2ooVcFo1uK2WPnKb0jzCSBuRERBPkC+k4MLZbk21QXwY4NA
66nPrXSzyQCbUuFIhtXA+69u2k8Ku7j8x+IX3maJ1pAs1xJji4FsaCLv2DHp09hgyHpLqUDpjfKl
4xNChwdyz88iwbhr6QRtbAnM7fl9jdp8oGyVmeMUjTtPbPUOa6rm872cWaB5McONeHL09CuyxCg5
+Digcn8HHphpevu/lh5+ztqLpTgp4gWl375zDvmv3OLQjPhpLgorieBnk3sPKRX318LOn4EEQyUs
QYPqVgOC8c+3X6KqYuPNnV1/DPtt7nr5hGpOF6V1H50rds8HX9Nj9LBheYDCDBZSIKQMXgWgtmk8
/KKVNPS5WYTnGg5x5eSQw9CbFlEWWGLL5I97lilfkUFv5cG0dS9VV13mpBE7+BtVS+6L1lbeIcr+
tl0kW6n2hrYnjb2Ns6c6tP1mbeoPYcWV1/9ntniJcMN9VVshgcMPnoNNF1gx0Id3jPGsaDSEBIaN
D1Nbe2xEUQ7eu6WoLiv+p3whe6xiLvRgHiN9z9YDqlvomfpTRW9WXzr0QGFQJKPFGdDYlND+waY3
zxmC9vxSigMe2+IonlUjwuh+iRH1n43GXTXv7BMPIcUppw6s3nrEiP+xK4pVB6CVxGKz8EsKIV8f
uYGVSP4H9nImupIivChD+M1TiYi/8Z9eQpteUog4Z8wTldrUu04HyOM17TTj0qrCmXopvPxiXhRC
bOIih3zRHHqicyWHJZLYk/tGR6LKbmQl6fCfrz7yCMlYW4SBYyK1tSpFyJzX61GQhF9N0QyYikXL
rJCFFhSsoWAwpPXWCTcNH5lwsuW/7uhWmZrYgcdpKvCssuXkX1C/G5mNxBVL3PT536jYA33wpiSL
4D01r0S8cj0sVUw05iVaG1en+GkpyL73DYS0z9NbiZv79bnKPu2tu9A+0qDl9gh8eZDLpHQm1dNn
FB0pF8oto70Z/EUxo0e9ses9L5MDm40GFYzR3WVmd2WjoPPnBxK83D377ZZKKmxmoVo0dx5a5oLK
oieznnGtzvMGiPYZaZI3KP4Qi2/Dszu41p9EkkTge6lz5iuwjQP4gRIUZgC9gOxyRzOf91AGdBQ2
YretRsnszEecsjlNXFMaldi8vHmR+w9cq6E4qZYhODO+6U/pH+Tx8GMVyze7lyUBQSJtn8BKJtg1
ZNwAH6cVRBhSKy+U0aWuyctVM1McbS2YXSX8XpyAGNEOox71ci/XkVXAk+YYIWC1RizYYSOjreUd
+OJdBQk8XE2YmSTXKdCRgeOQDh3BJx5hpsNsJSHcjQzB/Ksdr3w6EVUwegzArrTRxG0GZ8LVPdx0
4ERRwGakqONgkqFhXYg3d+ma2+KNZD3V8q/Kq2VZ8lW1xp1NjHUOe1xdmTwcdsXv9CwFWw00Hz+O
Ff0fCZjnqovyO0wi92b38tqu7jgrAGzEC3ARO1xbjUFQHxdvl1avquA4po018BAamIvXBxdnLkWE
b/8kye99DR9mLDt51HNA5v7jWWwA54TRxW4ri2LSeag+Uq7ttL8gWozUlkBApKePk+nNoNfzAGFJ
M+zhAG3MvIwnxeeGQ8VWCvN7861yGUJ9p/UBHBjwaEkwLk00d8bpI2IZdj1yhp3p30+s6JkqPCT0
8hlj9s0lMQ5eAdZXsWFQBG1sJM8voq4OoBSVGdJEJ8Zb6o1XHWU5x7j+FR+YIHeLyAsIIM0ubhM+
qgyS5Tb6WlQgI6zUvmikkkJvFPS1MZDC77WTrPe8qFzzK+H6NWcSRzrlh2oTupnPYSzPkUb49RFH
kL+OecJawiDSSa+ouTVWM4Mrfz2xbe7OxFt4j53czTq8mOw+cW/42X/TIcs2jvLKD/+bnwEDLKQy
T2iLWQ4aiGVdpuRwdGT0355VDRa4LRILSYxuRIliFLOIyfcvJ5xJCC0vCdrDt+NRiW9brd2Gi0pM
mJBTVrVvkfZh5s/5bZeuHdj+tXkzWrVFR+oHyYEZsiSoqB0RDavo1fdirsZnaW65w92uAgQQ03dR
8OjKBoGiRvoe/wFmSJujGJOk+OwhdxvM0HKJnmETXzK8yKIeL0wUcyIh7KCrLSK35zb3OnlspTUf
WWR4p+qA8A4SF2XcfbHltoCdwbkaDt508/csKrPDl39LducODSHPzkZuxYvovKTNVOw2h0iXjQ1z
io0tKrqQE4TsC/38XTj487VdPhRzJvrDSbzphimKvp4JHtbsPzXl28JbBItaXtNBs7pTanePYxdZ
ass4sKu/MuOprDCKt9JSy8ksVn1/h1FEG15du8akiiFjc7YqNton4jTg7y5ewTiuvkYUJMgvUuiT
MAqZfEei00ziNb/ZXF0ycCwSil7wZ642uaLgNlQIlyCMt17vAnKxXMnK4Uh35W6vN0tyZWHO/Wlq
laltj3lYZyHWcfxP53PteRrwiNbHx3f9Mh2uCyi+HZwG3fgDkmRNE59Nshm6wvQOo6dPnxmQu57d
SW15Bjev30I+okfwPskcLSWHg8LMgn0qHiQt3e2ieDjA8abbdydWRJPx+RGM9ijrcdyeZM7NJQYZ
Ct6B2YvtN07E9zNLuqZVvC62aY1NpCc0+672X42sA/3U+8qCtfGnWc126xtOnWZfx6bV6n6pl/C7
NAOMq0CZobit/enBy0N11nY4bQJqtvk3fuoywHgq/JlLWRTO5gyx2y7rV/MHtyFUuCwbKTGAuXdJ
C4dzDEjXCvC8w6pNHqnw9ei5c9mR2VrpYUhf8Tk2N4yECjxQCTVt2GITomlfauZuokFii0RaKYkA
mbzGJg4PQ+RLa96GDI+OVBrttof+3vAsRzm4TKbHh8PdEvarKam7WNlsmYiyytMg+IrQtZ9xeobD
LpF3TymCkrR0WjWnBwf49KtXn/afAIDBRpxLx+jIKHrpyYnk++cJI5wrHvM7k37EDBNkT2EweK+q
OtYaRaeR7lXJXCHTZrj9/htwxa63qSy9Th67AMtvw1gqD8ro1xpsu3psTJIVKatE09fKaS3kyaOc
5nT3FTlK6D10YbngrevUCVLnuXRjOkW5sQx1G/PwtGX0aJxGX/3KwNhOHVplPvfm23TnjciDlGXN
ic2cnkm5pSwyC1L5fKNJNNoXZBaZp++CWipsxjoKdzdOf0Cuh5AKS77IJiZy206qgsdr4wl6FD1a
LSMm1TnUnPw3aLws7PLItmskV3MSmjYZlT9S2KiASmKD3yK1MhF7itfBPkwiZZ6duxOBa7IaIxoH
Sft7v7V2nU76F3Bv5AP83OQXbZUYrhxKmKqGbhRV+b15oTO+hq6NmWDi+KK9wZlLBAz0Dxi8TyG5
ucBJXrYQwBPTZlORzSCQkRYIz8X84evF/cf72YLNPeT2jphfhjUIakM0ez4b3K0soljIgVkDty2c
8N415WKL+2nmUjoa5+6xkNBHaB38r1DSwrkeBD58vmzYLn5Lsdomi2cT7oZMNMFw0pZBivwU2a1F
a6U38mHL5FhyU/sob0sPHXaiITrNZOJ3H0xrva1r7CnLzHwARFPU01XcIQNTkG4WVu7erezusVHh
voz1WtQyF4uUeKWfNZHWGNjLMjjHkssVOBaC3+3O2xYFUBDqss7Np+0+v9J+Uyr8q0VBiwiTuAqe
99YJvYSCyRouDipjx/pRduiz2ixwJyZJKwEJlkYizT9Msg7evBXtLAC3fGJafizQYHJ52qbNfYhu
3cmualE2Q1EuSQJsyip3aNeOBDsI0mAY2cPUdySNgTikZbBLtzAukBitaAKyP7N/XyQzRUHaoaF/
ygQkFDLNtQY+lx+KSPwSvx+gXk1DZGOrFN4fTvCbrSfOAxQuw4TaYyPr6/1fIEGdbOSlsKHqjNaq
OTGbKB67BSFdHLDQM+HHpkWx4IvviECZQVyLKTWpq4tRkHOUEodhI1m5CQf6BOrBLdw8Z/fQFJMX
8fCybUXNJQ9l+x4RVL0lrtgn/ZHk9ppRJR7fg+emM+UghMt6QY5KYbLFFZQFbRp1P/qHFHuENUz8
X+r+nVGsw3A6dnzvkJ7WsLL33zbAfB5EpJRnlmF28uc5Mn32ofY1fT6gUszIwm76Teu1BNhEMRVp
aMfrx1OyTqd3D8Izqhc3ro7cQva4nhp1xWsrHT0AhASDdjS979hxEWjaSbDgBeM5XuwEXITaJ8ak
yJMa3kve3370PaJEJBn2UgtyGXcmk73lBrKzLl61cmpgpSE8YxP0YgR7qjq0eUu+emXIPj9KTpiZ
JB4Kvp3pi/95T+0z455hzNKvBGQIjyuD6yKaS34HudoLSZBtW5/U2cxFq1kINQ99kPLGhHN85Lid
LFwSJtxNvBRFrOCwNtr4TYa1ywANvpHkeNKy2KO4BigjVS6NBSmd4qwzmM3VnAJmVj4LzO54HHfv
bJ5qQaUwUF+ycYriJgzZrNrIQ79G2K7k49ET8yBKvCIf9ZfSpF9+HaJ7/m28PPfXrXm4jnk6FFVw
rWkCctrAdg9HCRJiP6ebsFboSyGO97k5CAxkZG5z0eXYe2jAylDGVABxjvbW6+zPcgMdVg9uZ874
9dlWMr6URJU6/8q3DDtW88RKKfLgbFKkdzjn6PtoYdThPcKd7jpLxhCQkmr8PON74ew5tGGBA8+j
k632SxicHDyiIcq9CGsyzFQW+ypIjDa5ouUHmdKssJSQ1NFAKzrxAp+mpvQsyjjmeiVaTcp7HMHA
KbVPx0c52dOxIwzJSRXr0dnRVbN2F4Tyo716RteLrVMatZTKSdEbI3j50/ylszFImna7OeLPU14L
n22PIg/AEKDMl9A1Dghd1M6gvPker9a41pDlJcbR4OwiczSVRnEINuPBGnpbXzqDY5lTd2AKyxP+
zoCZn7ixmh/7xTNlK3sYC3TYD3Z4o9cYUnO5doleiq8BDx9TWBTpiKkL6SARlC3pldZnscW+9qpv
yomhYH6wDYBIg5+IASe7yGQBvu1BMW2f92jTzfGLCaD8jlH+zVsxlXxKWov3sY3HmGzaAw8Hagpy
Hp1pVsiU0BzlGuxx5GWnt0Erjno/AZCqk5ylKrUUCWWdN6+gw/y4yhn6sxH6xueaoQp6HhlcqXtX
YeSVefLLWn9Q21qXQJqCYBW/MjP+z1djR5wXNDerJ4Ajy2hqVzx7CbRkh3yR4HInDnwAWKHSdxpt
JCv6Y5r6v7AVBrlUNy5HQjj2K/299FkrPNa7zb7VrWZb2/ioPtI+Cj2jrVO1nJ7mQsaZL7TVd7vd
X01yIJiJ2ln5LGWhF21JW2uy5uSJI5UDENMrAvrtS++j5yH7DkyrEX/+JN6BJ53aLQ+q2YJxkipr
T8R3KNXITY3gR5KUVUagz9SchXS1v31WKmTF/2KMtmopDY0ClP9aMrChR4wxsAfKJy9WY5EF5EkQ
RTuzVMm9y6l7qVCvRH9siRGvsjErm3U8acZ6S8zPOqW78DOL8iXsL12fPG/AZ0QvZO55qEcqFQov
2KhhBHRHkxlKes/L54xskrew6YVJh0HwEIQTL9bl5lZbZaLI6mmXYxwmZMuHOfY2doKi2yaRj/4V
wUIPkc+zcrBnTfiDXvjdj3nP7/yJYXfCwPczLCN0ID6/3rSsVp3bErwYjKtINeR/hiSs+qPSEs2w
toqF2l6pBQsA5RGCuXcvx4fPyZ7EBimbAkls26v/lHDfecYEV9ewtZPY3/LGKQ7piiMx3hTj2BeC
QbzuO8eIFpQC9Qp9KQ5rfl3ZwpLNiGdS/Z4PdKHxS5WbfC7GAIKmU3KSjQdA+C+ggTybUITC5suY
Zubp17gpzlXDsL9GxeEbNxd3lgcaDOii4MAzstYTQInNuhc5+C1KO5f1lex1kbwoUDKarUWpjznT
OfCSTBqUHoNhHu1DkTuUztr5lU3Qmr5pGFEm+aPn8cIueAnP+7krBrX6JYUlmleOw/tHntKGHHr+
mD33gakEHgvE/3+UvIMM3dd6UTvIxV54rKF89i/pyU/LR9BiPjqoXI21gn9cqScMh/7yBASe+IMv
16FSUa93RldDtzg7LxgecBeNAjNq+8rf1rU4R5m8mXxN/F+MaEHVoPzAItljrznAf2V8SzZ3S5Ca
Q5pylgpW/1oba15QPjf4OMs95nGautFoVACFNkVGojwKM1PjZjDThcgYceN+1IH9ZYnQ5UJQ1FPH
Ru5bZz+faH/PnKR9+zJUJz3SMP2a7hZ4vq83zvT6/nPG3frpEVGd7+eOquschhh+3r8K9+KxtSEY
awhPC45/ocRI8gsdaivh8pH0vHo7vr4N5Rc7NbOEWx4BWB5LZBxQTRVb5xoJglCZeBi06L+KlKA8
5YN819VkV+rg6ir4Hqda1Cq1L/022l28PwtF787DRg3sWr4tkilLw71XmHjGCgmwovSQXrpHlijg
JLigQQU6S/OXq3BJKEnIKP9OoBYuq89s8P/288O5aUMAik40n5bSOttHglbTOx2f7AQCmr/fqGAS
EMlQRpYFlzY+7b1hw6MWQpZgZgxVQeqboE5rf+D39Nno1xwYdAs59oi5MsL1waFzw7YsxUZ2SgRY
gfwwLh+uTlv7IFsUKqaGtgY9UJcUdvtHXv8XlPmP1vphf8sr3+sLhgbd2MyxzAhktOu08hdiaI/U
cXWGzi8U7h7P9lX71saAft2I4fEd4btXHvBpvsSQVLr0KHt9e62J0f0Zb1rPMc3mJUje7JM9GokV
Yi0Js3rhsdrc89Uq/R0sMFRmmDMWX3sPj5AknKVIZMJotk+tOp0wb6eA9O64OoGdcsdjwqLX95op
cUzv4AcmkmGaM2RwiMbp79YyQzAedmk/mt/HkCnkpu6sYc/GuibLEJeGbWvpqYZ0H135Xko3jxxQ
YRyAsjKe5bLvWizen5erbLmkLNN3X2NfBHvks+cP7nLfxJblGhpYhMwwO7pxTGgDC6hnSStmEA7+
94j/0pkeKMs4Wts+u9wroAGopH0YR5wwdtBWBhmSB6XE3eSP4kZhysZIB8Flkz36veoi6n1YdhC4
6abFcJb/t5NAF/amCL6AfrRJPRH/YckZclQtBV5NDdMJ+2+rhigJIJyDRROUKzW2UsmCHxxjIGlD
edi3Eop1eICvZzTzfAxMhIbl3zda2IpHdOzhT0zhI4A9WBov9Wx+pIIPt7YuRgiQdf441aSZGkSY
3d2OpL47vQkpHvJ8MVckgR69flnigQjdSnS1TSNyJS/wSirtTKik1EOlkfP++LIkbvllgRj3/QUz
NZ7B+j/L0RrlIy3Gn/KlbCRREhvVJVgGzb0p8Qg3aRfOFDigQGxi09tSbK0CWQ51OlQxL/o+sLPJ
MorRcmj7t6HcQTnrJdKD1GN3MsPvtpSlyafc0AjWmI/he5nObWxn+n8Y60YkXhSNW02iMfjPIIaB
YzGJIVqvYLbdtcjsqzzzCzMpeZDdmKVFg8eKLalj06xrTqL9WNuoDIdrRm+kJZlIgngjoqEegLaO
6yR7JETzqFdr/CxP9hrErg2OylJFY2p4dkPQVZCWpoVGhjcUo3Skg0FHIzYYX2BWV2DgX7jBh/sc
YIIcB9QawwuWJPb0gVNMRcz6v2izIGFNuzXZCd/jeisT1Je06/1himLl5YknKpSZfY01B1G49xKi
YUKK+EXgV/eJBix5JUqIkRL+AvYi5pyBCaMX2yk89t1r3hW6101Raq0qeqwcdyndXrp9p1Ocvgf8
C19GTIMYP1a3huRWIpsMRKvveKn0vbBg/jXXFGYMBguDDx508CMZ3qRoCqlhYrRw+lMzzMvGTXpU
IK/hvk27E+TFI7eLLa8lGOC0axKgewYFJ9NQvR1iTH59WyzgDZWuZR0RgT9ZXBGsbktrf2bxKO0t
SawmpIe4mLROBwv5B9GiC6vLliALRhIH9XdM/s5TOcMb+qaVe9LTfdgnYy4B5HUfJMpAH3BEkOXd
+7tngTxgphD5E+ZPopihAs1iLJ2pOgrxGLOrk6SDl/gArYbhvZzVXJTgI6hRaxO7FN2EKPuMVo4b
braQPVuO+6olvi8HLSUqvlhdN3lZAu+TI7qAltT3Md8KOjqVS17tXIiuG7gNB2r9pj1pbUNJ/EYS
ojkKCsi/lJj5vCSvBbq8+UZhrMcinruToIePg45JXrTm4gNQJ/m+PH+mFZiIOK2SLURJNUkCTgNb
+XKVXbFNonEKV5lwHmHN7Iuvlqhngi0i2MwahxgsNlxeV+xdrTZprXVxIFJ0n4Ld6cbnAorTkT5u
6cmVFL0xOopVDRsdkVWnuvmcGex9CHQTCkb/gi67tdhlqKvx1izB3pcLptLx3Iy5oMasGdshfEaX
fQXIBa7lYwZu5zqRM/VK7AvaJFDGQ/Ja/1voLOPwDXFEilQ8XOMcZabC4l0eJUQNgZ5zYhhP6qsY
8kphZglLDtNvwFUqNDXFuPuVgeoPysujbeVan6tvy7wa4R/zTXFA/Uz5MyczLpiOA3FTs/9AGbKb
KFjyqwJBVQ0S8BEJjA5Sz1zL4qCr4NGCngvifkJK7/pcof9aWBlmcc3DW0Qx4PiGeuT1SqAQunpR
nVUlnIyFbu9e519bDa/DSYg87R7YLB6riuds72WITAQQ1mkss8z2SLoVlLZiYnM00wYyDc+OshG2
IDy93w8XY+GMRClh3HD3HOSDKogEYdwkZSQQKV5waiRaPDwHO3B9eclyAxU6lmcGNLXJ3cYdKakn
sPkoFMAB5hu9XThCe9wgQ2EPZBAGks4S+YHrQycQq4buEP4TUnWbbD7WKO8mvEyPoiZ0FAfsoa2f
UQJ3m9bAEy9ekEV0bABP5S8Ko3K/38IPW1T79MfB2zLR5WqYqljPjw/AFZ7EOf886seQGf8GPI/n
5oMOHYMIDkiHV72IeIh5PHxcHgfCwRO6wd18LVVK+lf7W91KjQjeUeMxfn2eiX9TPOv8HsX7NO5a
DuBJF/F4cfI7DGGbkDtjZv8Ypvh6Xx+mqwlKjLKuxt/bhs8/JtR1QPZJr5E2ExZwRlyuusuTQ4/e
xar4zrZLcr4OLxrvE2WpZ2AYEk6/4emxaL8T7GEvzQ1mJObyqjDgvPdABACGniZhm/RAfJH+4wEi
6kiv1X0iPUxRts8m3R8eFsrh/9BhcK2cF0M4A8ISBUZrsnqAU8gHyD9XBk6PsRZ2k2BlHhM7gpAZ
p/VHJib0E/5SYZxb5YE2OwuW/SwlftacI78RGRCCHFzTfxnk7U1ohIZhpHlzh3HjQtAxCIeJaDJQ
fPGn25NnTJxbQlWGRBI/28k4/OI/RgBxR+S7+fxemVYlbYbtMH6oNB4iYLbz+u4g74a8SdJB71nF
X64488f0pVOvtsh9kKT2esot4awxf2PBIK6mRJmkod0uDf/h6T31G5W3y4j0u88Qp3tiMPlv1nlM
ys/0sGMCPtGAkL1zk9h057CRqI98hqRKtU+OAM5uArqkaGHvfcxmCV8K8SS9O6nrpr/UO83jzVEd
VcaqP119rz/7syxd9BA/JZnriB8qjoz4zUnbbrLng1kZ9CVQm2H904BbX2vbEM1f43jS2wFOyixg
9FygAPX1FAcBQ6Q29bIytW96NgJX3KP+u6D/lFRPgSeRvv9OrUknhxVFC2CLnprzFJQugYfv6k4x
dj0ARRFTKdEND8PVO7xhfJ8NDMT06Es8uwM0bgK0Hq5UoqknSaeeX3D8k0PNlSk1AiXcGI548/vS
SCuG5JOIkxJYbH1CPPtqkCqRw+AmcGmk6wMJC41jiGkQ6SiBwy///snB5M2RPy8tB6JsrrSG8bcG
iWwvx8BWfcwKn8Cu+mi4oilSrCt1lA9A38i0KRa2H/hUyUuYGlBw2fRqOWoU4nLQgUHYJqukaJ7l
0RH2Ncs7WF4VxlcAWZUyEGE7yu1CD851sMl1c28KUfvES4wPDACAIlR0YI/zcFPfRrMknEqv6QeR
1L7KI06+reXitBjoOphfRGFlIS+L21noGRHnClsDrQRLoH9iK7K5OFmgNUeGwUMHYXndi0F0wWnc
v5lYrnXjYH4lqi/nt9WGVF2HIkb4WTlKvFC5pNOhb45rvytMWcr7YtXeIaxDkeXtzqyXm+FxzuYz
7EHnDY30+wVo4B2gLLj1C9LF7YsxVUJ8/5ZXqkEo6yktSGey2+4DGFABkvK9Cio4bQHWXLxHnd2u
VEl2iXdr0LEHkZg/LwADeh8eNP/f1Gfp2hr5BxY+e/Lea3Os8OBK521H7Ri6Im+/YBjIa5X3d1ru
00lChJf/V3y4c1sPwdv7MuN6I+vGuixvUoyF58Zz+OfWoA1LDLC3Vz4+Bl3CgPF864BmabY7Nlts
gx6MlX8/evHtbb4SGYlTYLMfmX0MVv8oRQg8zzpo7YyqThC1AEfd82LpSp3wI2hx+OLvBPvE9rPN
qZ06CrgMuGr5441wzUHjcatQO9W26iA1faaQfgCC63ZZ+2NKUPMKlOeN8J37zkTARwQBj9HnoMMd
iXZ91ciqAFgbumD57Fqctl0GlpbMRXroeQxlA5D7w6S5th1fiNxiX8HCBXtQ9wT43pdkxvhi7B8l
NTezCAuhz0SupFkp5acMjrZ6Ld7hlXJxZhRfgiNl1YIsIbR/DtAu8gIEB1rEEZkDgAO0C1T2/bZr
rNIDaKVvtEVFRJ0XdWgH880qToBe05cBQrIepky1i5IU2NifunW/jXQ7+wJtHBMSoDVnSsjEUXZB
QAEznW1Hw2Sv6wEtrFrVKztHyvfmA/Q/6vwkX58wPdbhkBjrTFuhQAu5M5zQSTPHYFpgZceLxIdG
VHMEvPTtpfjUqj1j6n4aKdKObWU2PSG1bDV1FM+18FbzIW/SMPzCkLDKP9Ott24CSLU5R1SI0YnR
GqNg5d9sIl+aWpmgJkKjq8wNSpQtCQX9qiRgZ0j9/TDc+kstXaErbISCF4MKLvXaymV7BP272rCh
DFZJcq3kYQcFxQD97v8ezJqaAgXukJW3S8vPiQlVbudsdkGEykARHZXcGDqgWtLvxZ7T3AkqK5JY
4YilQAVLOUEwE/kjVEae/ThirEBJjAwupIobj9kWnYAsDdT2KZpKhO3SQ88hCpg1cfEcxXoc5POW
oEp69hFRmcWElOO4MFXblGs5CyB0k8vKhCfxECHEbk/B2DZYWuIeB2ZdV4HIqgzQkpURLUubsv+B
TtqQvR4+yA1w3uUQ1FaTpZhmxgk+k1EmpXCXfBXqCwp8XhkDFHso+Zzl3PjBZJKg/A9riE2w8gfR
Tw/CQK4Qhmrn+zl65tekHRdj40WS9s2/SGD04U6xqiFMJ0RXeQBsxVa6dmwiXSvNluq1/0/2wkVZ
VJG9FZI8YT70+0SuSvYz5FWDKCFZtJqmxDDGUlQYQx62/GreX5K7GBbFz3xtf0whT97337C1QZmF
a64FOprDZx4yfdgYqEaDoo/xVknq+q/0y9j7HtMueP4lqOWO70Xx2T1rXOm3byoAoCAvH7pU/X9n
kSNT07xASikVM4a8yDJZWv0ENzyiHAXbB9V4GBEFP/sNEsTtGKVitBxjBNXGH01NE/JnfzqpmNaC
bclkU3Eycc0FPnoYhEJlmlT/ais5GAigKp45VAT2jLD20BFC2w+WDUCx36xeVgb1BIb9FCtmaKpv
a9Jao0ouKKPV7TlcYozkwvJ5HFb21TI6Po44PXTSZxWbAzGVTspOR8U96Z2dYI3ZCcPwzgIQRMmC
7kzvwcIDrGbY8HvJoCBqL5Oe2xqwHisuywUUdeeIiDzEkstBdlGbjQApAJa1MSguOkiG/SBdXy1u
54IF+yGOmgf/P2hlKmuAutiNoltifie3dlbm192Nh7hgaouXNyfBwh5CIZV2KZ4Sz/PQCRKstoDw
lBgg20V+fZRBzSRNvmxLz7gSXal+kZBbfX+6ICCrWnnpdFYTxIATkP1PQPCmtm8PcqXUGB402I8d
cAD0ZNp7suHkvRMZDPFzUHi4N4OQCWXCuBF4YDRepyHLB2zutx96zRF8kKAUSXKHxKn5CJl8apV4
v2F6iIIN8J+dk0vAcqDt/6QobCADQN2hch+g0z1pWRqcrUY8XWNo//ALo3WPGd0aBl4f/CIpzFCQ
dT26s6dXehWk+1CIdqFXYXdUOooQPhDerpcbHX3/PfICuIiAldsivDAYFrd0bb9lsIcpDTDJ1xF/
a+0SMYfhwFrJZS4GUGRXD4RLqjcRyWwvfLXZ2TOnCqacgtpNR9ugtIwnhdM9jjsbcC+DHkEWAuRm
Sk1tTDHdmXlPoEXvtEc4QqucbnZvWbd1Ym5hHtsPNIne3eFxJ12Q2wfUxmxdcVmp8VtUsG/FCCd4
fh5a5mQivNMGcjAm9mpBSwWblpmufLLQNvgbk1vlBU4me+5Tb9Z8O03tB9HG2IPwkNXl4jitGPVc
G4YT23d7/Nuw700j+3yIqw+OBkFBhREFFL3Fi1HXRtzG13JUeUNw9hLGBWcZJ9Sgy7Ph3ZxqCacW
mQvcCxTthaORmCj8UKs97L2yY8KN2QgeRLsnC0kbp7pX4Vgi1jRkGxtzzTy+KztQ+tzpDaeJEoug
dNbVZoOq0Z7+NJoBoY+FM+fAEvx06TkdVJ4OzljdrMbaSbAxpV8dc0Rn8cQ8qX8dNEsNVe53IMaa
gv9VyI8SY8xOm5DF3Uxo8qYTGIkBZn88aRcDy7ItGRVSMBp3G07ZG1QPv4FeFWGB8t0SG03LmdUd
YDJGjAgl5gvEP7rY9OljwF3bU7kJvE1hrLzkuPr+txf2ztm7VJs9t6srevoJDETmcHocfGdtNgfA
EkyYbjNKWn/Hxy304ezsdUH/E0d2pc6OIxpKYdQey8YaUUv4HaUB2pPHiiBvlD6W7kowsa72eJhU
kUT1RiXRcI/g8tLjawvGCv1nfE8xWsTVCxYDWGXoX5ITidQfJjbR9e5iH1qVYyWYtRa3kG8Y8keC
il+wat2vfPbKmzOVmpQUfclVXErul8dvsZ2ACy4NAYpWqV7c9mXW+of1QHPi1U72YpswPldvvfxr
bSAdEfEd7y96eshKLUcLud4KTW5G3Kj5s4dWqOvFjRVb0ADfIRgcR7o8eMaSecScRmVqqOlu3yiF
uB5Dw50PKO3N5a+iK3MB3O20rkHxqX3B29eGHsE5x1bwh08jq+vEYeUsKyBT7x5m7pFaOvTZjVzR
AJQeHJpDm74gZGgkPVwmyRd0bJ/Fj+Bmke7DSDlAAbolmr8k+SHJYbzkvBDFjuGoI0e9B+iSa8WW
0xepqCJNw9cP/AbEWy6vErOEj6OQezqKXOubbKvkPFQ/BHQRKBg05chs/PSIe8XQGu3mlaHTDc5A
NduVsJd6KVLBuz5IsA2dDubBs0PfF6c6pooN9EoxG2VXNa5ma7gHemHS3qkKu7e5mSenlJQWF7OB
ki77aiicL4U3JrsYuUUFLN42E9OmHrLxLtSLVyM81XVbz1mZvSY4/LYSW0AWf1ST3Jq8be8JWWKT
AIAOjpHRXMld6erkWPzkrdEtqiCDCY7GaMwaHcp+ClRYl+IZ8fmCUIp3S8ChoohWzCn/sB5kjYj1
epNHjRyiyNBkylGhFaD3PL5qCxxhQ22DSzf2jyqZYR8B7cuPz4ludgTacoW7/XUTwl8uZAalimN6
cbGKtt+cjWs0NJRuwHwsI26q2tcNQ+jjZCzDXTRsF/RteysonXAZI511oe6+VFwFK/pS0trLmzFH
6a59LC9bRpzW+ZTrAiW/9K378Z6/7H2FtINSL9gx3EvHxWywdZPeLOIZb3aGcVpcVTe8iYpfs+P/
D8cWtHX/TuKd631TITPjXT1P3+ksjmBM3pE3m9HKXKcpUtACkh+bP1QLE1DroF8a6bjfrKQ077/V
rRLZr4BsaA5uutagM4agRlrcs24/rzR830tssaERqceNfM14NFsNTGYoJQnBFpknfHrs0i7NokVg
4hks1gqmsoqLrKBTnj4UAdxvvqGnzt0jPLPzwL9ZwA1fhqi/eFZcyvTVXjSueIdq0dFrvTRUdaO8
khGQAQzPTc/KQL6SIPxFrTNAzyQ+L2W7ZE9J+2CUMDGNuAtnHL6mN3ZwnSHewIIo/f+3lGJ5n2el
fzfmxs3C3d/roximMPIEJgamkQWJZigGqJJGcpH0+4oAKKn9xHX7MbunOCA3VYVfrH1I8cbX1Kw+
6zQMfM9+vH88AGw3w286KsjOePQ112UcdpaBSUYjVv1MSua6WRh2VeRe2s870XAWJFr8uOUXtEwr
FMtBCI7tlwGY9nJh+o0gqes7pAVeaWRXhzLGPejPPACqyrVQwKwQlRvnKVScd0qZHYZ5fjQwxcer
Ir6l+fjKH/KfgwfAyhkPPmS2mhPrrmOCQ4pgQvgKuCyHO8FtrAxBJNkWKZeH3hBi5j9sPEajvli0
B1CS/GymNsGQDVjoeAIlrugwQFBSiA5tgHnaxlgK1sFTNAjTV9npwuwk0xLcPNDridwbDA7M4vWa
OWgcThkk0sU9ASXTAMryTTJbz3ZDzbmpfyaeS27vBBvlKZlkpSqMAr9toEwyFQsWtDMA0lf5T2fD
vJPbUwK3/afUca8k4Op96d2WrNoeFDBZ5odx3sVa/0eeAtGIOtLx2LAa2dMuZ8JZA0r5yAkSiYS5
DOu6mADys7q1E//M8BjGRomZqjIELHuZOV8lXQ74X/CUvu2/N4DjIClX7TK1JVhxiTSzYGOQmMeb
Vl9aZPJZ+6GizO/j6piyzpvkTTUA1Inl3M5WkmYwWPPkKwKoz9jjMylza6WdxXJebvMqw3qXhRAZ
YU0EcM64ZDC2UKul+2k62GLmDhAHmx61pscec1h+SkEA0AosUwPNQSjy4QtMGDbgNe+0h1267KQT
NhI75EcLFVBHP58DwZS4uA3U4njaO+wXjnk1YoRaXjY1qOD2mFJPChgkgdp9vN9RA4TUKwfvwlcU
MfzAsaDZJrPtadhAo4veZLY+A8z/Uo51lun08bZw+yG2MLUB6hiET3Eek/Wz1B3xScvCYjoSjeXM
LkmOxOVloZXGYL0kaVsO43tenZLct9UrC1U4UI31Snd3r6EjMZu3b5+2+NCk3/pbVbeZQdEKDrAS
fur8GYFD1f5x5n5GESr1yGOq16pWOB3UzD9AHI0aoVxOhBfsm3oZsrRAQgHHRUJ4Qvss1qg/n7SM
DUt8wenGQW0EuxvwoUnZ0H23rjEZJ9faMZ1BfGr3FiT7/o3OSNokW5NH3zK2Zgu698Yy/oTvsYiw
sTXcDylsEFfpfyyGx7HCDhfMm977d/U9sbV2EAaxPU3Yy1nNsSdT9Ok9RlvtJrVzVTRyOtT4KrDV
H593trBQyk329L84kdIiBemT5qzRlZotQw8zyPvKF7zDCRKMgb/ABf+t/VYLZeloMpr+0RV7XTrv
jM+Tp9gAENIYvXozE91rtMUbCDbvlyKx+DyzJj06N52RlbVbD7DAK3WUNJ/rjWTJ6GSUQ0krpAUB
YgHH0zLL7NGU+11f+MwJjMxm4VlGRLjMqhU/jvwnlqRLjh6AVizQNgySn1WKF24dfpYDR5WbBgSu
i2BIO4g/IbvR5eIRLQHc6mhH6PImWppyJropH86KjZceVx+2sobWO2K2+UiIDFPN6Xr0WMwp+zpC
EputCeDFxtfWxTVF/H8984PIkFqSCi65ZFoEEWYj9sTcFX0boKbtdDHV16faiv2jWI8t9KsD0Qo6
jyXHE9ywEXCMKCI2sQraZ45cUNPgOKA3UQ3NPT7sl6OY2oAfVCYXIql3dji9K2kMYJSvjLzcTiUy
WzR2M1PRAv33ws11aLD6EP3tVfy4yrf6YLUIuvImF7bVUXjDyx1TYoTbcCkNfM7JYWzifNqW3eJ6
kMffQwXTEtQhvwEOm1ljhz5bPtZjwdkNbP1p4Om9cdaaR+NygQhZIJlvEbZjhRkx/T6RO5aPVVpC
qU/+IAdW0eiv1Xk12cffP1YFZoy/hXYviwwFibQRwLuOz7OdTmREAmwzZ63ECopEKopqP1XeSWxP
lYmjY7IUTQXtcVnNlLIZ/JLKFVKwReKwNZJzeIloqsuquTC5FwRmbhaFwGr1qxXwyyOI00zdiU2o
OezogxJ/ssYq4n+0ObzZu9dnoBsAZku7dRl3ivYQwnLeuec/B9ou4hEqSZcefxvL3bPneit0uGts
jjAxDTMjT760OxCUAt+rZRcnUmUgtdZqzz2bx9B8dJGJ30EH7Jr6kpsZnlICyd4w2Y3rb2b5zv28
9/glNrmqBimAwUlxx//0P+211Hjdx3TBQcUkCLbltocwtSzV1jTMOpeuudgEn+KySh5cqyJLasWY
p94N52tGuyO31moaS3lJDusvyBk5/Q4l4NMjh4uHHLk+mKKvFll0SG6SEC40uNzvYcO/1ntOyYR4
dtwOYQ7Tn2jrSFz8KaEvSbKeqiE1t7mjbxZ3+C8HUBEGNc26MWbdyQ5VsCeDFszP6G/TQjw+f5qa
E2u0EL9uP4TsaBhgCTDlaDSZINiDGvNPPsDtNSUduGJ8swN2R/JDREr436aFoYbRdUa9ugiV1/4s
pLAnzJQbNrhh9rAQ0gEinHSoQMhxxAhavReF/LPP3VqDjFsTWaBhyB+r0Ub6K3GZB/bQdM6Ka8QB
8K/VrNHq1xjO/U6VmyCy5oA5/oppBYzcd9T+Bmec+Pti53Qxd3EOGpb5pSSYQl4yAy3nOvbW+mIW
yDe+c1bnZvE4I4gwX26XmlnhlkpwKrMGRHezTiy8UDbxRt+gvWOP2zCvufFOq+cESTX6Zs72lFZ0
TWafwQyRvdJSQiWaGXkDuSEfvpVj/6Mf/xnXF1GIdM7UpZANJNijyViQ2vcPx0dw0dW+7W3t8RFr
h3vwYwfF+S2O2Ktx1S1e8hyf/NhczTJJDOfE1d8yKlGKcs5SgPOd7krBOe/L4nLQrlNZENgrunj7
i3ditYm5ZGJaC0QQ6JfBTMyZjsp25GfEsPRPf5qDj58YXRT5d8K9l4bQQeddj8TPz4urJsXnPeq9
+eJJukDbQX/HZ2Whx/7bjXPSaJ+092W3vMi9TPlZtLLoTDvS59FbyayfLUPmcj/FFYpfMQwquk/z
5iFNm3ocPzghatJhzoUlLrNtWUIctKEI6HsOdsb1R2gOYJbl7T1xhP63wCIOOOvTt2FAnSEL6+zv
3tzMXWOVsemVGFFFDRSKOEGfVj+jkHD2mGFP4qDsbP60Gbly655Jpl+ydvj+ASMwYi6Qxa764bVD
75LbQp5CPlByRiAPqVVS6N22l5oM42hykW1/SLiospQxYSf+E/MS39yOcoV6YVbSmFfkA+YqseNk
aqGhxZxxd5BeopPAIdoe1bEA4YQ4BF1dXfRAeGVLyGOjTIE5+ChupmR2rcfxMny8ppI6loyjdnLY
InkGDzxik+PAZzc08hZbh7UUZKLtt8VWReBFf4lzdlcaBL3D1YJUkDj5pI01aDsCLyH0fcPsoOho
2LAxDCmABvOmK/9L1NrlTluHJDD2uE5z7SgJe9Pl47aI/+gmGFu4mJtk5/pmGTe/JYapvyneRgMo
9jA1GZHzabWHskAH0aN2gjt70nj9NwZ13P5OnEf++ivv7XCwY4YUICacf9pGE8G2I+f9dJ0g4ahO
W0SfqJkj8hz/PZf/O9mYMqyehItzgfhtJQiHRx49Z/EYSgPI+/ZZ+VumGxTqghHwLd40uZkT5iX4
v5EHfAh/BK/KtAp1rdjoLux0jAvuP4oHegBSCKoUSEmiti2ji09n+jYhmGDVa7/JMliiYHtPPKDH
YmV7s5TO2BC6jc3E3kZVSnxQ67kaw/WJlOo/PLGwaOrZGaY4oFyHg08IQ0gBqwg36mVmmWa8ZICg
j23b38c4qVWmZpYku9dZ1X8H5fsUieGNa0SMnpaBO5f+W2mvWuWwqqNmhwMFCkacaZqBEOpXH7MB
LvgHAcw+/xFsGXP2dv+Qo/JzEPB1DAGM9PweSE1U64kqejx24K97XeKC1QW4d56NFL6z5QypnEOB
gtDYfPtAtj5GprJqOax8OCfMOkTchPgPCbFVLGXtBLhA57WiRvvRth8YOm86RO3AZXa1lRKhjZCQ
szgDEqYNGZXvVB8nl0aMcvOzkgqQ1W6xdn3FmwNUH6Zu7qQ4JfDhqTKsGwNmf714a4JdGlxK2ELA
x58/q6989rGLXqM1gEI1jtjKbLsyRAFUchL/3eBnyA0ZnCzVqqB0i1ej12P+N2V90T21F+lUjUoj
24nIvkm0Kp37Ret3q/BTi9yTFa+pBefO62rcoRgYGEz7PINn5HKevijTah4O9Cmc0FoYXeKqUhcL
2w8SE4BYVxA084kHnoRIW3f22Rgd3JcOH9WqRhGHS9UW1PrBvaTB7WTiEoq0RuTV1TyKeeraPly4
3L4p//CDhdVN5d4DB1rNLzgBNYfMJjDCvLjlfVyiDm43BHh2RSg5FlYYQbh2PBTTHITYSFAULhwE
qq5pGA3msSAK4EfHUlfM5SG838gVAPkQi5xzBgixmTc5MRmBSPne/TOefe1TR2bCd2jSeyw2wMve
FEn9RnLSHIMrT4N7APzJwfyS8yxC/7WiIAUpM2fLlSSGytHYqD8WAd0CNa24SIPyOL3hs9jy1Qrs
xKKed8xMUkQ0LLKYBB7wWkeOXd6QRxwkCwlAMF0E/n3ibIzZJ3Rn5hlCioIL4n+xU8mAIGMD21rC
Zpqq3uJ8dI6abs2IcMuKTreL1yCH9z5c6wibK/SroLk9S2fswMwg4LfjzxGXbCpffKhAM0te+qMt
YQaewXnx/v61HnynERTh9XZ6lH3yDWsW8K+WVkZZqD9ptompx9U03oMOh2AiilX1DfiiZs+ii7fe
YI3d/K1ie7mwhlH9mdbJwBmkVJzZxdy62NjIGBXynBCFyu3Wwv1S9dWyXo15AlZa9fMOtXhvUKy3
Fn5uVf9mS+POtqhKOhKZJPRJB2JGHouVl7a65zAepv/1RadWFOYb031ww+GD8QwYw07n1Hy/WcDA
JT8Vli+C/2XjZLiQTMOTJedc/SRddyKZZBfCFDodezWyOqbzN8s7cv/cJKjnQbXBP1WY+xVlpKCn
IGjSmsfRIAIcLkopEgJ2U85feK9uONGslVk7YeHsZzxmkWd9z+dPNk9CoRddqcdbQkr2iyMonoiP
S6EK1SpHEyVLBU4qXItrK59UBtN7reV9bJHCQkbIBW0gx19eciVy76hgFIrYLcLxtegj2mLcn0Rn
Jaeq5Ch2WPl+u/Q1VwkPJKbMIRE8qQUXNS40cYK9TN24CQLcYQ63zSbPAIUKSpngbUwVBT+dJOlK
xng+Lc1tySNBf5yfFrzZAs/tsdSKvKHoPVDvat9HjBXJ0u/vqR8XwmEcWKKV/tYmuiDlolCvPNfY
AHQ1F4/MPC8aSPh2XMjFATcEKr3IxL8uOL0b4ucP4pJ5p7B04THTr10e96Gcr/6S2b7qyE82yedj
q9RL0TtYpggNj6N2qqLeLeiMby8wkQ0ZDjbbggTwYCAWpHo3Y/14sarjz3kugCbVhrGGB2q02roJ
nGxsZrg7Klw0IvwAqD3uzFsh6OXUFmgUN5iu1H4lV6vy4aWT5YlOJ0IqQ2eNj+i6z2hH71t4/Tel
xj5kjUCZAEZgeb5ViGqSxt7/xplrNmY/lrOWzxL9cPOfyvrS/uSesvdjl8OE2ZG4E3wLoD7IlyKC
B/R24wgKMgYzBuSJZvryEHNUbb08SUMLwqsxMZtNnfKcbnYQ88DaZKOY9wGIhueJOFSvK1GjY5Ar
o8I08vR3sPjqJ+yzUiM4+pBqepJIS7qA3JOILMUPK7JF7OBqE0rmLSIWlGE1un0vPoFcKfG8VvW4
N0DPqSBfql2pH3GrojZvYvBSrD9o0aUVHsJP2pmUi4e79rZOORUVPkOCkK806n9gWCqN6i/yL6wZ
lxqaMqmL5D+7UPagwmAWt1vCNfRulHdKly/ZXE+U0eWHdHO0S2BGMYojrqyR5N+2ZH6YlWkxfQp2
ZESpmVsMouShWT7No31teWmh9ySTxK17t6djg5u04wCUVIgub/YaF3nKW9CBo2/NafgqgVxCRv2H
/nI/LwI+A16YDdBJ3anH4eW4ZGjIUUi7r8KkeLYP9pDjjAvVGwSgSahXrpLbJvD0zizxazfs9Swk
239envxoz4OGQHVfCCHg0XdysrPKELtFB3PMN1PlAF5B+T7y+LmoAo4nZ2acusWmaa0Z33AtPTRN
fhYdhZ2ZlaDvmb8WKvg8Z0CcqK0hp0ceUaK2vMb+IW2yUbcJdYmTVGgHuNfTlR9GKY2UD7Pghols
+D01qPnbrWpccJGnkzCzuhG18niLqanr0MV4A+VQ75ndueUC5YHgx8WfigUBME+e8etJqTr/jv30
/YWwGcXAg7ZAehbV66CRDpwLM25Rsja/BPKue7QDF9TZFeDF5yLrIkC31LjU1SjdPOIwodWfG8PQ
z9/dQ/KYsMArmQfBNeFNe5NRexLfHV5KnUSKje6qBkIgbQjw+nAxMNqFXxh4t1uv7RLEkf+3/6ps
926Gz9eUPdmaVm0iAH1LnbeJ/T9PhwrPNtJLhVkYgWUWmEZxdySErVHxJHtEM5ulvvZx6gx3Me1H
/EW64dt7w9qSyNK2B2XnpnNgO/4kas8b3Eh68l6aLUZatZ+sXzAL2gQouz3cwPG1/Wd4b9zh4A87
5EJihntbAgFhS936w5xzs3UspcXpNLErITVeufc2ky/WWqrPbBeyqRjtrBQTDgJxscDx+I2n1kJo
shFAX+pyBpEjzlKZ8UbG6pnmm3uyQidWRbL9vw16AAL/UKc/4dq9nVLvdxHUG/0MmrR6lak8qaef
mpc3xVwcQD8x5V17/aJDMKrgBezvs/nFRdVcLmlg2Lpu1VFU5GCFCheAmtUsMqzSUDCPaxvXyJnc
IETT21R6OhkHoQIyvY6rwXwUf+dGmgzFg/McpDaxS2k6uU+TtvxedV73gashvyyH4o/Pf2Mwb0kk
63usglYG9LBrf/wlsxoIQ8yogUL8ymRPF7ZF8qYpMqqtsK0HM0IU6I8n1RjMDGejwoNUjvtO8MET
d+P9/zxalG25Dg1rE8GjDtT/2qVuspa9En5b2T+aPa/iGbeMU91JW4kqV1h7tbL/18YfiP4gw0Mm
CO9NmDuPdZeCE3RBudU7h49GqChdqryg+qBIAx1L4JoCcIy82bBwBftjOhUy/C07iCnyaXr8CL42
mBLS9fsYvmTz40ZQmSMC1u9j8oFnz55xtM4xuI+kQjUFR10MPaZPzTAT3QufOp3xhT2kaFkKFij0
Nw9p/sYVE1EL/esItAQbEr97mdt+YjxCmZQdfIUU/lKZToZrKnMURsOeH5CLh1KopHhjbuWe4qb+
RoCvL6zRgD7P0tHIpD4y0AFPMmGks/p5dTnuLNjUXykP5zVnS3pHj9NAi4eBVECGtCFcPIe3s2iZ
DrRwEHcboQS/0cLcT57TQRyKC/G8KzNLktUFSZZ7ur+GGIUPaAO6fihXuGAuvNoxymWcvLwppC0K
/KyeiaMGq/yk36MyVqiOG8c7/0a8kNAxDw/XotQFPXhu+JvhSTgTbVCR5ytwvuEiSokg2kn/dH4w
2Vv2mCQ1znSJUI6Kbak17cVBKLyvQDGTAxfa/Y0cuMHES5w/hz6SY02q6fUXxOHVKhzdM7Sm45X/
m9DmX7Je2Q0+Ej04Wri6GKbs4SZ9QrEq7e398I5l2V3dKY3ZAhdhSk3UXtXW4UNVOeOJbnRitte7
/azQ7jW9AxxTkusSMAUMRKY/DDWsu41ovjLMaBLt/tTrErUKhy3FNwBg03GjFOhGVUPSzHUUbyyZ
BogHopwTN1+RIoYOrEQha1JDxWY67jBaXYAm2w0qnVLycK0tONUdKtisgQrf3ub9LtdGQZSkMhi0
2pOGG4TFYB3D9CHujEQ3te6eRSLK/WCfnE+gZI3Ve4ZFJo/MoL2czzbvfAe9W/jmItMVixHf2coJ
+tT45K/Mfq8z56qRKl9t9W95DiG3iO6n/WMdrwb8QAyZiBfU/zr849QLgFcR4JP1BIg0V+6NeN6I
CLxCSGoAUi5WLgxkzLVDq92Uez2ePw9kHktTy+oqh7GtmCk0JymWoBA+a0JikrdeTKYzs9yO2p3N
Vlo7J8utLhP3KVP2dlAjOR1dxKlr1flOwpUm/I4vhczf0FD5QuSRbq+qrOS1i+4WtAwFypsC0whE
+CW6R3DYH5W/oTRPjvlsiMgWh24J4zZgiVb+Osvwze3aR1dv+PiuQwiesX/J+GynBC9nycwyphNw
7WdV/50Zn2+MPttpbcEanT+VmSzB/55//krmMlbFRFnmG7eGQIp0gIEQq0ovk3SwMg8VekK+a8ZV
KxafZJKm65RgTwDJrMBd/1nLrQexICpow41v1eVxsaV545QrLpmpLiBEx2WGDaGHsqNvou1jmoYa
wHaXNGkjGoryCnzp/qqqRwG1ZayKZ0prwDj0EZZLebnTwQxi8heMkSZzYk0bH3f4uyyYk7u1Sfz3
ctFefiTHJ6p2Hek5d9B+4IgecmVXuCMzrsCHAqHlbThSeifY/J65ER8dWBDGAxXYqstyeoe8ZmV0
JoCmYj7YvVyPzZO2yKPE0yOMHp/5rFgEtOw+Hw1BxIwdHLh9hq19lkOFNME1HFXSXPUsrgwohN/x
KEzr7oGxF1qy3Zn5hxP7k26mJxOACzKnXqKJUiHZ/HfLIYXK9ggy+0UMM8LDW1efkrcYFWL2rC1e
0WvpttgzmBChmGTakG0vttkPy3okJhIM3EcaMI520eaM9+1Y2l5NiSV7wHUPMwU3v+XQ1piNRO1m
rRiBpYTpGzkV8zmu7gM/4j/IsTSG8DLdT8zXnSk4SH4oquPnLpYkmUr0JO2su/1TZUBIjJrdFSyV
M0j176sA4TFTzE3IcRvM1kcr+pYSPwgQLbYzBWD1A1ny9ndzsGvEqbpTahf3Yl10ZqctTOJgGrs7
kE9M7h0mw9/cWwB5E5KVvvP+MLltq7E1deWAK9J5jHdTE3R/3E5PbOqjAzCqY+JDATpjxpsNNHPG
GBI+U6lDL2Yeu++FM6OVAO6kBtm6BEns4ZAZ50XDkGONX1ri9l0mioJ4U3kdc7O04IM/RV9PmjRv
zLpzmJjskay+qy6KDQ+NxNe4ae0a3uq0FsQlPyhb3bSJoTMfaTL02FgbIKxbN18PSK+Ujqe1lvLh
nNrkn/f/7YgavUz9BVA/jhGZk9xgxcB/IvRYDd5/TVmwdeePDQHB2pkwW8GcKV3ogwp1HTn8LGRK
yGy5PddI311dtDugTRnN+YEdkmAWV18w9Q3VP2rmOskXn80nouQmUnO+GCSelxHRWSVD9gD4ZfTK
HGv+c0zfeZ6n0TKkw8mgaPo7rNViq0KBYPwgta3C5RMnXGUQMCxFuPxYoMELAUQMJJX6A/UxE+3I
ufnYLSmHazm+dQcCx6YoegmTnU/s0rasWsnSrTrhjij8UiMGFmyMIffa37f97swUXYIbw+5hl6Gu
6wWmxAkT9sii5ve0+9vV0OO2uRJG175+MAmFFmzUmGsswnKTNyvVyYJ37YCb2vrvm9zQ+Vby9IEz
Ww0ryi4/MKhYVOWbUBNmn6/pdb+zp2WhGyeiFTMxQWfk5dNXU0pDjw6NcgDMeGrw93VxpmTe03Oi
bay0Rk0USU9a8EOz/mHh6VeKq+q8CvMfgdx2syuw5Kla9DEIaQM+LrzWH5mZIN+USPmgl9LT+B5W
O2bU6EvxFumW6WfYVz+4Gq+J3YFVDOBUFHNVBh2Kwsg2Q6nbCTK8Ddn1nWKnqXluYs0EfsFlY+TT
nkKfFna9FhflUuQmwPlpUFsUORp022HTeES93B+q7NhvBu65eowkLrkBL40VAYOzGNq2apN2FQWE
kp+FLHVAZclOH2VSBOISZYpS4bkv+9VIH/vDBsqf7ORfI7Tr0az2sY8wJvruDwu5DqhJEWkV6INC
mibn67QfPIEHWm2Uyw+R950r2M6jLUtOCRXsFWE9+cHpqNArQNEn+Bl9YG8HrhnY7psAwwVMKsNh
Vrx9M6wul48qVhSwJo+LoKFIZ84vJl1Wdsycu8rmzLOr82W5hzwY4P+W+D0c4yw3HxYbMKZ4oJKF
9yKNH/CUrnC9JgBn0IVaToQ4kseZIX9/ftl306uDml8+f6IhPewdI1MhihALWGl6cqOlmpZeeeNd
K8kMhRSWVz8U9gDGygK2FDZDlJmD7Q66IeG5gX739tDNvp4Oq1YmPn4zCz5+50PL6WXn6Qf8C3Ln
RZVaijhZrf1E9s6ccpq3dF/9Q+SIEB+yzczRZg+SMH0XGsQtAnhD4WR5MZjxwhS453wcomEEQagY
oDY7NfzSwIfPvShj1WDTPMRQVMBs6EgVcBPPCltTRiRRmvLb8zHf3jJC1qYZt7fP+vMLtEKhyxm5
loeUv+MXr3CBr/MmXpXH6BaTjVR/FHiTh4WehNhhEJy4yb82A8kcszMr+rbrgUWQAkfAoSgU4TVS
rYIussclKKTNeEqPUlVrUTmXYGEs5ZVzaREVCQG+iv1LDuWPpVpHj0zrCiiEkByb9YS07Py0sP9R
dO0HPlutx9gO9De+hd+aV3gqw7U1hqpPaog6dvu1PwexP7Z/MUv8bZDh27dBU1rHBddkjtdE7ipc
03/h97gSNKqm57VAlUFdgMyxJD6tGcis1AO2oBDy28u4ICQeEc42iXyJIT2L8TVJOVx4TBaJ6FhA
owfHxlRyBGokGNl5ktaEZHIBUJl/qIxLjgWEvvBNGqLTgMilOdTYDjdx5TVTuA5LBms0+3Ut63Of
8FYK1kx5Qg9fuM0C4poPtKlOoKeSs4QamF9dExkpfkqvpEIRc6nd9cet1Zzsb2zTnyRXjiQsv3JH
G9JB+mOHvNttFTLZ8zpRUZaD0L/H8KA63ecuZE2rV8MXWrX0hePrpP3M5zD1EClIcwFnKdE5dUsS
koM+96EoybyoLZPrvwKSoOep17pFAYfe4iI3C+gQJ2bGkLOajQgdOHG3ji7BIMGJwHdOxxUWh4hZ
wVVHbAIDAQNwAxDegEXkfGNS3X8e/Sl7UIUKIvDoEcEFV3JIFm0GOjYBG7twQY6NkgATq/NtKxvt
yoigVyujvYMis93es2zl/a8dLV/ZpTp6ADB8BXeNuPpVlackYHtSCDvsEB0xGr9FK5Oy6EeoQz77
pFVcHZGnW456KDPEEfyuBj3K0tNWBNTw+cst97D3t8WKJPyTAeJZA+ZgD+UPu2QMO4FDMNxsbaqQ
nvnqqW8239ALW9OBcLpMnhDtI0XPF34O/3attyiv1i+HJFWh2/u77dXME1iWwXcb6Gub7hvCiiL+
eHwcoTWICz3T0hTUFjRhn7Fe1aLa0++f5dXPgzdQTBjgLNLCRFIil30AQuRVVMkowi+m/98mVeST
OmyOE3g0QMpSFGDaQkUJvyM4kk1UAKP5BVXHrtKUf8Vzd5Ft2dLRGNh9MkolIm/gmoJYIkKRst4U
YfqDN0jrOgcDL55wR0BT3mXL+H7VVylRI7t98BmC+SwWsC7pX9yeajZ1/2KCU/d3IfJ8CZDgbKXz
h+/Ifb/QwsCqec6lL6xzXxxszTyqF2DPM88kRJd87orVkMhdKh3C+yFAWjCqI2PYc2NhjUSFgD0j
5WYy8YnCKELUUgAFpIRSvJ9ZANTvA7i2WuB9CzFl731GbUe/HQAZ6Wrn8voR2FyrwAL5PZ6lA/5j
UnRNAcAOnLiJlLBblVJpTk1ptdUEmtnvWEhtulZo4mVPjD8wN45RusmuTMpKWedxXHXjPOCO8Fxx
Ed3fsQg3lsFql3XgFIqMvFxqZPXJ++XjQDviLB+lNVb+idF8GiGTVI5103nFmBCxc6Xso1M/BKOI
cxcdQQTPSXrwD9SHGgmAvZPmqxc5/61uLRwBTUU4NjiI2U/EswGcFRyjwW7499ezGYjIXHKOJuCe
lIlj2+FZgbxqUJb3tlNnRa0yh3Jsloji1a4SIy+shaPIpRQz/mo6wsF3TYexwH19cl55hVm/bTrN
WE/rI2cO9Ys/ugLiwl4G6eHQHtruuu1XstCv+mXiZmNIfDhXzjkN+kjtFUVmgAmKRhwULJQClqut
qI21iZTH7P9tad27gEBhnyH+dhFjg4K30vLjszgRTILkDlrhoLE4Pwv1hEm6Ykrn10l+rHyRh9nE
uMionlyElWd9ie1RcHIOjf3AcG7zojB9gUbbNdT5Y4HnxTYvu7J8DpbWPIYaz+O9XvPDBBKlZGmx
ix8h4Ju0oENhx/XqPD/2+2xor4bK4X8ryb0DnoY7efGVkyh1nsVNn9C7fvURvBpLLh1tGdWlhFK+
bacCP6zev1M0A5LkRUZ5OmYBPy854LlfF9uEPvAtn/vRtKJWUU/PnKNPF3GIjt9MVHazrsPfU+9R
Nr30nZQdzEIIh6GgtgOqd7iwE/ELgShdh3k2Nn54VTkY5YucMXeitdnNEdL/mcNW6QsIjYIHCBZX
k3gIR3KjobANwaRFQ0/w2BRDujJs9qD6d+ytak3cbdrxqPIezNqFvohuL3GyjXnUwwVdXGIZAyqG
pV4H+0SKecTL7Ua2PbJMep5JJM3F4GYgnN0lsjZjTpV4bllONYuZ2IkDfvVZW6lokCbOfFVvNb/j
v7DUI+JUVDhvw1jWkH+pdUDptlGF/aZZR6RQl13wlofjfIFq+ubYCveJUpYoFTZutlIyJn49K1CP
OLVVxLHRi+yu+KX/KKjMzEhIn1qnOpQLKxxq7Ph0Jro8+KqdnSUqbqjQFC/QMda/oPIQv7StWxVP
0RA0vukiBmbPXW+34tmnx5tH01g02L876LI7W/g0u9BBZOPMYiNA3th/rHeWcN3cUHTXBO06FNWX
xQGoJnFY1vO+NahWapl0FjgQSmDtMmh/9ARhyQ6YHpSua2TeXYpqRPZ5P7HvXWGwbtD6xcRPD5bP
+JNJZfgtaEUGDRZMLA89BHDJr9qA85xtlpwGIz6zjhIngUuZzlWfqJPE81+TjTjzJN+89l8Vn9Lp
kLdiXEG/tnS8peJZ634ZsnSg7Mn7Y40gVEcwMlK8bQ0lE8kGsFUlUk4LVbukZwi+puOvAKQOEvxp
7BqLED8YwTi1UXBQHy7UmwfPRL1ghdB/DHWWyXS2PeYXBRsEictXzaKwLBAwTuV/8kc6xevmQSEL
Wx6hkh3X5IMXaLya/jwMoNi/cWW3k+zZrdM+EjxG9ps8x/JxfFkNr4O7ssrlao8/EIZmOv6BBa00
PIJexOM2SLpOWOxwwHjOzOKNw6xbAmL+KjzKRa28M8biklckigv1l8vClqRmSAQogVIV5l9J7nKn
+LhyhZUtHt2JxUnHgwcgCRahWRRM76aofm1ssooDm3l5GMi2oHoiVOgyv/3TjxpWzpKcW/x9SZP8
bTNYsEUwhpj2ABzDXkQgm3N8AWEvzJxizugslmpBZ20ME6uh0ybgI+F1QphPqgdtDrNfbvgHFZiF
cSFeGNQFI6aOqf7Z62PvUzNxFtbu+C8s87IFhxqHhKDEePECqq5ozidhyXl3gndvXMsXPcb3ZSC9
stg2Ms23lYEZ+arosaUvOoKDSZDlaVEJRf1WkqdOFL8sRnYLeiYzJI1sePRd2uq+C1vX3+U8RCsu
ZCJ0dxs02jvJxCkYDHFP5FGUKn1OV98yyqAeOtVV2xcUQcsQT93kc11gs07wk75bw6rHJqUfagDm
dGvXWGa/Zzvt+iJQR3GQqv+D9Wb0ieCkPWrliKiytylfQCslbl/KNL31i+p6Aywg4QG7RojiXzbD
ME6/8A4RK4z0ASvC6jIDdaOSoIEeddNNH8nqOdkF+dX0Lwg+TxdNn1w21trmo5Aj+pz9/Si86bLq
TxJ8ERdKNUeN97dEFO8WWAItf5heI6axjjjQ/q2yNjkt9DyVUW22i+vD6BQC9FnYZ0HCySlMfkW0
BBqsT0hswcRPMGeLx9g8zThs+64Q9d4WHltbaUEZlaqA4VgcW054K/0BpQYbUBCSDAsVQxzy+lfh
S2RKkNqiEGfghDqsUWUTsxAEsTBfci8VWt2Nnny/OKKEqGsjwV9xd5FxaMMCj5nkc9RPDhI4V9l2
q4h9srPl6WBrOJfPAe4jKhll2VDVFEUKJY4uaqMY7CnftLFi3WMALf5KrSKDlQuTncTseP9gG+Vz
oOnaRX3BWHLwIVj7h+odcYxXHjisOUmYuLPSiDG+InI2JRgzCbopVTAI+lx8LAjw3gX6wBcUWSta
2BuBbm6mbaF3N+dV3EUt9V5uPjMneU8tdpgakbZGxR8ZfxOhMysqKW2MZpT9PfHOQL75NRaCvHnk
GFOU3M5gov0gBuSq61QfCFwFyGRaU9lNhyzHqy5bYKDiiwMXsc7CjQZqrGXrmtSrFegc8Kh2b2ys
3XTLoe7Vs4ysQwfesoZ3Dg9MC8qL10YLbn0/AJHiL4ttcZ1BZGYW9eB1Vj6XcrIkAqVe0EfgHFRR
0syOrpCW/9OyS8QwGxU326Htnf9DEQzOg5q4WaGop8TI7kUxVpjJGH/TjxxR9+FDiIPgXw/GK1Cp
vdAflMZCEIPiHPeOoPajXBDUQpVa2aYPZ+d0RhooPS4+e0U00ifTzEqhyyzx6mIhDvEpS4d2SCD1
ufludIAiZWGUMItU4zFNfuUWhs4SEY1akDof86INso8PtLeKBEBo/7ZsPEoeRXp1a7F8gV9lOjAb
NtoJCqaSiTquBddWDuMgWpMt8y/XJmLtMnudGPPI6C3AzIZd6BmTWJ0dQE2XcZgcVHmoWQfDKW0x
Qq5bQufw0sVm6B3NWIyBdxpdvUUMHgvMttKsUKzhKiUS/RtCm6xSyxkRRe4JNlVk5g+GO7CvFLQg
GNKAicgIdUHHZIWhgJJ+rQNEWXtqGxX6BkbZ1Z8Xq3HsqWOeHLhUyQ81Nsp3CDTxWzZkDl/AzCDm
hu1C+9ie+yzBlMsvJLICHbYRNTJsEsesNBXlvXptyxsMN+crhFQSvPWx7jhwSRSkDtQOS0DqawSt
JPpYhYJpRE/E+marTqMZXb66GRwaCpVIPkv1iIMCRbk6UL2lXUIva4REQcth1wJSNV6PGfP4f82L
4PIVl8j6UZIr92549KFyvs554mfqAI7yXJ1SW5wmGFWM+k6a2TXwBFU7LnMvWA403upeuWrO/Dyx
z4WP2tIE6baqP378DP085jVL8p3WcPhyfGaZ+C3tc73ZEOlUd1izUDl5YcTB4AVcBxhAZPwFGPYp
w9AUG0IIdcV4/LJTFPayJ0jtTUIACeUBcFEDqp7bNg9lyhwF2K8ZmW84gIBeKtFhD8U/VTiKvYM9
+o2SzeDgYQ0p9Yx2pNpVhnMlj5Dn78lQ/g5mrs6tcZiyY7cuW+zLM8Y90UICfUqtIN8VovPasi+2
C341g8g02d1mUMBT1Du7nI+MOKzqwnrauMKhlKy1vA+a0bNVuUDa4+ty1URod10YvXDrsa8YCMiC
YoBp0jk8dGl569wX0IjdjMQeNISpba3O1b9+RsP8JrXfZwmZPJdTETWeBQ4g6e6UImdkcoGlWgJe
eZ6SlVWUQpzi3lD67QJCdI190tFZo/RUn0bxLo3fUPfuSg2TUxd3LrDwBq5r39OmE2Q/xPumpYJ2
R6Mll/apVy+uxr/vWWiifVSHdKP0Ko+bx4aEJtt+h5fKs8h+SL0g/GuAPQaf848JTIKsCKDkABnT
07bMwkgHOcN6FU/hXKvTb8OpRdRxXoEpXIG0fwzyBMoFLAAlpw4R4Tlg2mcfXY6BZ0pP+prFHcus
LH8d+fcnjmFSmhS3TFR5czlv1WrXszt6LadIYsU693UjJt/HSD/fycver/8vByu/O/ayWvtJjK7j
HI+vvEqo1F1JUqOQlqSNdrd+xbVpDlWTK6JgKtiPL3QlyfWUlLxjV1F4+E374tFUFtqBiyseHigP
oBZrB/OBSXTfBQmLiTwYeOxETF9Tt1VPhIJSu34oOUD5y/jNRFn9eMYE8YhKy0QZnmLglIoetN+L
91gbDIr/0eQ+uPe+PgrGBUCtOxXv6pSdYIbIbr12YhoLqfhGuZ+dtSGAWWengdQ4bsNU7v3/YmNF
2NwPvPdS8ZshtnGqdLXpWEtFqmRdLo4zSwGR4sE3M/QzjUGJYeEiCTEMTIH67l+Qlsdje6urpqGQ
HRZRCQ5BPGiGKcEYdvsU/erjkTFb5z4CL2v2QPngjfAycilaCmK7G/TCBLx/XKNkLlyUScPato6a
6qwsHCsJUh/NuZcun1PyzWMaa4ZqTTm/iThl1y36Vx1hPxB6fcXktOYqshu8/CR8pq8mjKeOaSJ4
O2ovV4csEeKcQT424/bYI/Fdm9btX4UEY3QxUscw1t20TH4fjEs+ygDcVXalGKyBE70+PbrnW5wb
ZWujXeqdS+NmVjSqaWp58ZFGfW1H/JW2bHnXdeGbNg4E7w2X0AG+EFgk3ayfAOV4LaJOZ7VjNpMC
hxuUkxTts2KRhZ27eQuN8QTtriNKvPdL4PJTC/rusabRuSR4hrSF2SnpyrUz5j3D/F+h6yuUNLIw
wvAK8zjh9OKsoQUwIo1Duy707wDhVG5l+ZWY302HyG003fHnJcgmakBATUh/oykPOZpCjufxhE5i
Zj4UjhP5cgp1WvoPRAdfVGzZe83Si+XGueHrl6P0K9hXEF125kyq2GaqzlLpdiuQgmpLsxhwfpmH
ViO2wNPVg3EEojLGZWsWxjNTQ9Ej2qGJj8jyVkxZfstEHzyobwytr3iPADKhuwA1QFGOdfO0/5Js
Sjf7QHEMvhsi1/x2UHUr4YpHQAvmx46aNUxdqwQcP/mmAXjKN9c5C7OtlYlEuN48+8RJRv6cqklB
NqzO4NXDXFOpUezTOpW8LMruYfBMKdvNFTeT48bCZ5+ep93hZMMjv7XKuRddmJ/A3LDc0XVkpQXM
jP8xdkBeX5dHYaPkcn2WpF1TNKmwiCVBWb5UkV/SC6o4LmKFXFUoYEq4bouo7u7J1+0d3/KnAP7Y
DEQHCQTcuYvPvSQtygmEIRt1SxobFmLwLXXXUVdmoMm6G2HyxuGgBrlxI6H4X3Ut+BAuU0Xxtx20
za30/C6nS5m9/kJ4hvwnhvpdSFelawXb1MCj0X9xiVv+OSJedme1Hd1KkriGntP5ezzRG6Wuek55
CQgYxJAqIRsHcCL/fOWxu5+dpQrGTKH2Q1HMl1O2J+msuWtqizzSx235oG1UxFnxecsKbBkVHXf4
OYjyFxTzus9RTcWEdihIiIsuMWLAxoNuni8ELLpPQmI7t6qXurvpkU/YlHiTjmOJIJUnbl7bih51
Kh+arK/xZAzMMYtE1G1+13fGH//GJLBY/0qWgkGOpJNMHHjGIY48zygkziTuOWS4IYFrC+r6/MMD
hCegGwlTxV65pqAFtfezZSZetLcO/Gsk0Fnv6nbkjLX0UDGeE1n+hOcBK9M1hno2yoaub1WyvkYG
qnoRJC/SAyA49NPlTslQX0yy0nnDfKeaiCnKXqkwGkxHYvroT8s5bqazwyAfFOyLud5Km+7moXp1
jPqwXtbI451j8ZQMOe6YEkMJJwqT9TYyXZjjHrNDv1VTiyIbA9SVyg4jvoXr7syl7zJ2yK0SQX12
YOiHU/k8MGaEtzx2jGkDgWaNtbeVRq0U9gOaCyiJIDo6QylzyRz6Hz6ujqTBUP8BA9iaQtIw/liP
kT8aA4hC+U0+s6wLOWhDdEJW42Bi4kabKXx6HilqGsiNuFpbET89Q8hSocWbtw4Ow48GoD2dbmOu
lLnA3W8rI1+yR6E2wK1KYzlf+ROG0+IMvuT847GfPux0XYqoYevbwfz0Wrw84winpRC8EAnnVpLV
COMN3GnS2upFJ9ApRqj4UTfqyc2k3BiKC75ZZBQSerIDX8bEV4lwNLTuiUgntHV3Qae2Le4N8tdD
IhqPlw692nVZkFEQlrfH38udGgTslH/z7LuZMXX3nZxg6r4y20bIlQOqJj9A6DqhWyzpofJ7QbWm
uCBahSzpIqUGYxkCFOm1mx8l+W/dVwDW/GY5w7mzhhnvt+s2t5T1Jqe0Ix80vMDe6Jdwn4Zjyidx
3+TidzG0M7GLo4crihS4kCaoGh2uQBooSxGOV+L0sNo0fd/kwCgrlJBlhlp/LaDihnvfi+jnkqhU
peqnO8ZALEXzduO2JKjawjvIOFqTfPEu3cHhPjisgZsmyXfVu1tmcPTGFLX3VPQXYWfGi2Q2X63g
FMmx3GF42JybfucIKeiaNe0Qn49nY+CVQSJKioj1N6dpKgciABiDbdF5OvWVtECCujKoTh1AV79Y
cnEa80t5vZG3SnUTNl850XpTM8ibfhYXOAJgXIH2EGcS+WOc7BsuU9Rc84C0q/HGZyfiPUWxZltF
7pO3tlI4yMd0YwxKJg43/PjejA7jttN2YmWzMi5XXLU5DQOZOD3KiXTRW1z6GfLa+1faTD2DErl5
7hj7odH2xxxVcmyKoN9JOrsORanNR9+Os/YqX4EFvQx53ggKSjulXAwQ6A1gu/mBCRVsJIOgoLG6
RQlMT8eTIEyqgyyukxjmoJy6w9p1lGVx9UCcW0lyJwr2FnyeXpGxC6NGJethNKA0m0rLS9mvOHST
dkHNyeSFfnjOdHVfXLMUyXqjfGonI8R4nvmNG5Iu4o77IKp1Ae4hNb7aValVkfFAUv7wb9sXS0lL
dxLWyDxTkdAjrmcKpDMHbECwupXpfuwTAKE5uGzDX25K1asQSAWwvv73nCptAwcEkBa2M0s2oLs8
h7vcaHnScs1IhFyE5CIM+6yyt+pQ/0K5ArzlGD6e3FDCFMOaO+Fa+T4F+bCIxra+oD67vBPixp4t
tkn2BlXEsG4bwMFejJl+AlSA4MPx4VbMhiGaOHIOznwS0oZSZDtNdc6xvKkVp0jPWXYrCunfyvLn
F+MzcMb9KiYbqTox7kUZADISCbXl0+o9kW6LZjzT9ayQg17LCNHD/YtIr1JMTP8pjfz2tpnrXaIg
tMNW+aXH8pSr2Ge29KtZSs1pq2eYOsdaci1YRBrfqFy9Y1Qx/HD4kKRLFxXqR9lFNWtWq6ce82Vv
sH9MntAMmLjOShj9NUyRQUXJs6gB3PUVVM+bKYzIIod65//u1vcUoYu/bVheHhHg0MgJIv8mnnH4
z/j7OWB6HMX9sxgjHJpmfowHeKJTKrOwtyMjbUayew0QYfWUYGB2njpdoDhbrdl6VNSBGM8OB5mm
jd4UPp/m0zOPfS7O+umK8oo/7U2/V/CDsOm8iOQ+GmTY/ZleoEMBfarE1mHvhdKhX8haGKqCrdnI
TkwQbpA8IYcswrMFQvTZIjby4NfkS7AFqNuGE2YtTqFdijT7IOK4NtjndtWQQwK3hMd3GOAix2WW
hYLlkNSjotjbPAbW2KaTTREIVKqDt/zeGStChG81EisYT1PKSaJrwP0LtaVybsjJy4vVj82vQDAT
d/gBlWuGSDhu7daxMB4AVyvc8q4oYwilBY7BRw8z3KR4s4KZ8wLZfikKh3oRsd/OKdDEJYibmFyO
ZQgvtpMxisNMG11FwExChIaARDLcWHmfow9ZDJfrzAYRFtLKIv1YrzrGmgrN+KF4IUxflXw45XKQ
AQCR2RcnN0JFtBq5Ltf79FsoyVUL0YWQIVHm5Mff6NnO0kK8WkhRf50KRR9pc5kedEJD5RyYxLgj
1LPTRl2lx9YIYvjcITbz3HliTx/up6JfYg11cXXAoicgetzGzMbikeB9PYYVXz3LISB6SH4O+uY4
zQj1b1N7xcgMFLdpu/NsYNqw3Pma6yh3i32shfCyfyAv+Lzq3JyfXCcVD4WC7ZcEhFpD3UlEJDbV
fWKItxoToCr393TM33z62r41Jy9rg8r5O8uhUhtKqi38elTzlsktBvShCJbE7ts5C5SdBJjR4nF7
eT8NZ7m72SIUzER8TByc3Qs+qxATguHDLGDTXmDTSmleX27WGEwlVKomU+SSSYkjrLi6FhYrEHjG
o0v2bSOz9ZlcOj/KbkSxs/HE1SZe4U4iykexwKPR5UHLPNybcxEOBj6hqlDh8PIvBx0zuDlPoeyc
HkHr8nE33HWHz82wR1rGWqs5NI5B+K8weWPwEWetmQ7ce0B90FVnBTbt4nVS05kVcWcxTffXazuZ
bdDqe5hBpFdCPmSZOaOhSwLFeXYVdT7ZWu6F61mQBlDnLbabXmEldybZPDAz1EgnEjn95QZMur2m
hyjcju+fWAtpvMSUngNjuAcZak8AWyLfsdz9Zjw6D70FpJcVBN/1x2zNys76nBd0golfufcpQy6S
n0WTmerzi34cOeSIv4E26K06H2YNFYUUAc/Q6gLJ2X6RAsWhfKfpg7xqO5UeBQmn/RH1uZoLEhXI
KJ0WMw7beiXK9nKUEW58VUWZt9dpYwLc+PDj0H4L/l6g8HH7rsENkumddnaON9ynfeE3mTliEZ+A
K7ZsY5Dgv9WWjEm8XUff1lrMrM/LWUJ46hAuYrL6fku/+gJN+eYJZD6OzT+nr7O7DUn23yoh9Vff
eKGKve+7nDOFUpgvRlZXiBK/4CK80tJ535ik2U3/q2P9rYe3a+vUi5pRiWEv5QncjaVMeM9+CGng
N4ZIZY5KSepGSROlERqxEChCssm04Vxtjtj2/ivSQEzgBRVogIsPWmerXdgHiimHDxOPwjZn7tl+
QCSaDWAS4H4jjmXzaP7mydF0Nr+L16iIm/mDiKQCGhbV2nFLwYJJTUOeamZWnk3Tff0ch45qZZz/
d0EfxMu9WZxiNkiWF6PMVEsPvEzzrAyFPLDyCInH+JCpt8pRj+kK4du8IEB7FAPINfIjg/WD2LSs
ccZvbtAt4BpOKbPPB0ie1Arv2qSfEreopfcUjzJOUnPGj/6bkQhAzzKL21PFSiriMTDQrmK2nTPP
S5lrR0XVbxkW1X4bTtTopLdX6AZmy0xlNgibj5wUeXP2GzPuENywOFo/GCOpaqXwU96kT+dZY7yQ
rEaUAwjAVDIYVmFKVr9vMPrpoiwB3YPOKMbZBOdAa3kihxxsLZYosfQzfledne51LDy1fK0G9T+r
PeRkvn3VQIRfSwFo4Gc9/XuoqmrxRXGQyZ6SIRH0IEmhvWROXA2EkCpVHPDuo+fc2z2LDE4aJ4Mh
u/MABBptQsw8Ts1fIufvf4bj3wNhtj8zdhMYwruKfIOs5xnfOSk7vUicyF5j5LLBkdUoFPi/GbAm
DpeszfVR+sumcHHkag34nL/Rb86xRm7CFvIY6V/+Kn4YzPRSxNW5sLVof6JzyqQ834U6zmY7j2jo
zTDZgUshShzMJKmzK/ndGKbHpXU5xz9QNHC/ZqmfpeQxn7VnyXN8/P91PAqEpLFPyBeeYKnzYQZJ
3NbvYTidziMezaGqxiXbaG7u3h2cOrBfPfqWMFbw5lomeQDAzbUGnujeqEa6ug6T5PTIUpEE9iTd
tttEkDXTDM59wMYqtRFr15vGiOrZv3uLX3wCLRt1xqNn8p++/XIrKcvYLSCoLEeF7hCt5tm0fQoj
UDTBQdYY1Cg/4KouiZlqY0AM3gstuyqe1XaMRT3KNJdUt+tm2j2eofNXUbYzgD84ly+4O4vZZJYI
uEVMNVuIrox1aOAyxMu7Zz5vignN8Hug677w9DXKjoDLPPHJ4RGTiCbWoIA6gOv9U/w68NND1cwY
4UWdZmABqH7BcmUKvykrqA7Mc3wFht/nVb+H/w+fHLCREEKdHDMInw0K9bAy62HtsiI3c0BzFJAC
4NgmaoHSyt2n/pYx4pFTNSiovc5GYxrqQb9PpX9fh02blr/y2BkUTJmJ2iSwikZ8apnEJcxUamNe
3xVQkeNmI1sukr6k7QTDBubh2MjfvpgToVtewTxzqSP8VXPlwzLDq1+O4vsNZziYLBZe8eu8jfJ2
QRMZY9VIhfbLk/Pe+lvYxRkvwT5/C3NizS4FKk3ESlOGu35VMNgYeUHeTb2GV1LjmABjN8fFsGPw
vajS++GJxMvcHQkBnO7UpqS9ZydClVyaKiQTWUGBGCPJCiBSrGqDQzTZIrcNj54xNoGGAsC/iCfb
XEN7UE9rEyKRkD63byJJLWii9U80Wikz/Y+WwnOrrpgpLM8xCivDAqszQo44avg0i9UMcxCi7vLx
nHhsMMWfVitqsfKlHLRhjCAxM/LGtZDIRRrqCOvI6Yp4xng/kpvs+z0brksn/PjskNwjxODfsqKX
+pdHt+SyiihlPiG0k0JZAjL6QSucXwI/mjlxbVkcSQvOe3rB0Dda4asXs1qbSjEsSPjaADZwKLAR
PXPfh6LlCsI1bzdirdlu4KKQ5IxquV0sD2spo/PgbDPx7MEAanO6wo3aUQ4binAdhzNks3LMwc1Q
Vn6R0Z6BmGa8Lhqo72N4xUi5HDHAneNRD1SBVW3MWlabr12F0olfwuy3
`pragma protect end_protected
