// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
abKBwrUsNd/OSbHOjyQ2RDfnQxnHfwXbxy93VgcjxgdzKvbWw8baJXrGQOjdcYdC
ttliBPeaElzJuP5OYX6beQfTTkxwpxMZ4ps3hVyzHW6obHmWfvrvDdR+IiBoXhV2
J7QOlCZmuyaHmBtiLsJeof6KZoXvr6DjyjbHNy9SCOw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27856)
eS5ZwDVf6unbMv2FFgFYoPJOY8U7FOkvhCbl5wL5hREZHt9vstN714I9F6ppeKdD
xRys5GoBJySwk8UapoG6NGDeiLS5L2twRW0ZJRpdwEILXq+898GV1vbnJwVjCnjE
w0VamDXVa0TyN5DoO1NYCXpCRxFPFVsqMnBzt/C6Pkn+YAnOt6KSHp8TsyZgmzNI
ohIB8tKPh8mDVxRQEzuttD64DXcKThg6dq3KQFyFgo1Kek6noJ1cmWvIW1mb1Cgb
320/maOiT1v5cb68HoWcizHdNrL9zYZJilztnXYhQT4dOP4GBLc4efLlcbjxG9el
b+y6NMlo2syKjeIwVON0n3skBIklO2UFzEEOVXehzc6yvXfxNeOsVZuhylLkUMlD
kcBTbq9KCteu1XNoCoLSp0VyNIdrsidkahCOel5drQR09E0UpM/kzybS+o5Gvthi
aJGoi8/91pnL13QRkX5Ep509XymQxcYc1b4uOm6XUqefkXjt7nSvFmM0PddzRMTV
KpaocWk2qCdQm9s7p2wNkK5KHZ9SUpOpAyXM/F7J8LxNBjkp7NU9xOXKBjmGxJcI
WKNpmryUCTSls5CHs+uuMMU1TC4OyyVieCit7+KBkHKxS/PYaOWgimiXkNAPMlbR
yTYLX+eZb3QsElWJm/OQH1r3sE7jeCVuPaATn8qthYe7sA00ndHWzHwctBn16WTF
roJpiA+tPO2mQAAZmdpkEIszrcMaCf/w0LHoKVGX0umGv2lBixUzfFf7XqKhl3Ox
Z2BRQanvFGNIqRjLqBEdMC+MPnuyDlUQX2v9M16PUZak6VqPlVK4FUdUooRDeOsC
XipmiZXWjKm2eqQAJ1zyXjkdcLLk7aM6+qRsx6NpiV5b3+p8axLS/bj3Q01K05/P
KrCWlw1EZKJnBpQfBxeJJUJab1t3suf2rF+sJ7pSp2rcmz9Bp9F5jFBRtox1JVRN
OplR15subSn/c5CCC2u0UPiU06J1izdufj5vs7gBnflNCnYXghavv7WcW0uz6wnQ
XSoBA44xxei1l8v1/CXFbrt8Kr2cggDZ+JTzQI+POl90x95dpXBMfsbChBgeZKwV
+O3mSKiuNOnLAq5PAFMVR/fmo/alzHLusg1esYM5rMc3fdjJTxLb/1pppslTdX0k
B3XX9LviEikW2xGU3n/6ftY51nG3z3cjTqx48Ie7tEiEhnNqEYVgPcZt46r5kzeq
Ev6Oal3Q1GmrxYEqoOuDMo57attYlyStigFVHMGvXeCt3SkyPEYFknkg9kTdPF4C
9fcNvxhZ6fxfz57Uh5MyjkV17Q65Qx4/Sq6D+tVlJwWkh2/6zHHnqk6uOzTWywvt
MD5xiS2nJNts5lmFHClLxw5e05CSqdsR/bh5P7Lala60U/vvpNmjhdhzVXDA0ipp
SwTNWVqHiCHooQj0Jt+RqGS9lFM9pd/eSB3457exYnbCg6AYKjThAT0L2G+rjpcw
aqWN0XxUwTGILmG3YdA7CW+XqAMblADsCQfTWSNqFiOG/8qZ1BJxyogeS18xjgLN
72Sacdv5rYb1rggiN+NKgtnsRdnGRV1GTpzBSdG2Yv2D3GuKh0iJH5r0bzvG/KLi
J27WjwobMctfUjDuPmFcrIDfFxk66mfrELzhDmgoY4ZxElRyMgR/blrPjLZIR+Cd
lcKaLGg1P3nJiNf49S/yg16e4ldiYK0uXbFGMFEy5ZI0hA3AJ0PzRTwXlQY/4usj
9ebiug8rxz8DaqrHIXniNxAd/mxhJKGtdIn/c9dXLeDprAr6SbgZDfZiQlhyppAx
wB5oUcctZQHqGYAQr2LKjrTeyyQ9UdNxsgqiiNemHj5adHpdcPFTB05sdO/jHFWK
vZ4ocO9f0vcLpHSTAZE3jz/Zi3wavIGymqlwxkNVvxFF93eqaPW95VQTqlNynKVh
5s65hQG+Rq2noOw1jbUz/FaxZbGv27Q5qLkm/qbp/HNxX4g+CPuJTqhwzZtfaAN4
YfnqW1cSYXhW+P+IZUUlRN+tYozkurdIHvjJKClFUOd2rhQT2sN7YkAUGrtoniY/
k61T9Alf4+CP6JFtE6kelYCiOryH6Souwq3rm/IBG92D9zqTnK7evxw/j60DAshN
x3BDcUD/dfcSbWMjSIQb7jO2sMvuaMXm9ep8lpaUYezm3PF4theYBGMz8+L/PEMW
bJ8jADuFYfGLYjkUZL+ZicpP4TgBbLnp3g+KqMhzte/ysU89bv4t5aJ+R6T67Kdp
yDViWwyU0sF9UB1L07dHKZG8oLcsDMrrUHB/o3F7x5r87G6fEWsiPdgmAs9JxwQX
gPsMTlbjnqmjbNVy+solM9SaR0avroHhXBCUYdb+f4g243TLbsY7jtG+TNdL9hIL
PVz0LtkTIQubZRrvAyuUGTx6WVvsKMwyiXJYsUfS4v1pSjyKK9tYPEiHqvzskH4T
IGnq2CYPvvO8M+SnuitndWen0hUddmQ7HiZjpLW3sWEO3V6nowBdkLRqyPtKzrWx
U2Ja3AdIP6VAC9idQUnpj6sIjwT8OXP9BKAVa7UTknJDuObvKUBZgEifmzfwVVsU
M/8jmoNQFAU9RKlHEudG+EpeXFN7p8vS+JiR+73CuIY7/z43PouwKRzw5gSgtBC4
AVjLwuoMh9l1MMZqeTvcf1znulDHu7lzggwS2v7DEZ4Q1lGNnp5OhvThv3bw8vC2
tktTO892++tjs1lK3NtisSZnjpGWl+NWQeBr1Hga3eoV54Uspf0MrR+EiM+S6nCP
+kp4Cw2alBFX5MnD2h5i7MlHtPRmiu7uOYfytj3f9zq73v84AfyZxYFq5OHBCbIX
tEaVqqwNu8inlx481SSPT16+RtutQBTdwpwcltV5jyG9xoXkQj3WxHuFfRCCGu/d
72R8TZt64BgsiO4nwtUZPSi+9RFkecLHihD1BleFOR3hH2a2XSHcsyHZ4Jwpl2io
HlUUSYj3gpY4ISbcsktovdpsLkThymCLIlUY/3mZM85DY7H0MahUHrTy6evvgyxP
ZnMUJ17OmcGIIBljcc2jkUJZRGTBGCK0pnq/7exizmOB46HzPTBH3HhWPEuxbR9Q
o0AyVdN8ZiTiIzdOs/s56kOTff5zXugVYt5r62p/FLnsWNZW9oJ/g8Q60uaPh9Pa
AnmCSf7FpMheNEv4ltZGFUj57+dC4Z0xNHoBGW125RR5F9M9Nr7yWmHsFUd03aR3
Lc+BlXZZHCX3PhJcoM4ypx9pI9YU938M4yrBdfmrcCQxHLDQsU5pJYl1uschUXH8
/hYBsZPEwb1AODsvKIDdnEPBTxU9nytJO6lQx4zbbl3/W0G5WWMILT8JiM7nB/tx
50HhHJbnD2UI/KadIZha1lFaKPPaRwtrv4USwQzghA5I+FXcas1JRV+uCY7UlY4v
yJLjKN1ZjWgnuP8s8PI/Qzrj+3s7PSmWDRUfiftOvsJhlXfjPeiWUyMhH+uEnPzw
eoduOKYej1dlRh6aAzTbq10SAbTDhwydpDvRE+vJthUJ9oSnQpJYZryVVjchi1Zg
qMrt/jOZjIN0DDSKrFq5tNdp4Slczx5cpEH/YiFcPPjjYBdEp/8+5EqbufT0N1AN
EWV4skmea0iPyWDRF8drCdF5htB9snUn2MLgo37qwf1I2VXrK2u4On/KY+kwUrzl
CTNSoPXGGVyJFx5XBZMjhu02hSdvVVc+yp0kNjunwHJKqBkzxlfjXa60ZWSLIZjz
KI8C0K20bJ/erXYPqbKrY4xKy8Dp4939ouIVvxdSZ7IxPJzslJnDXhfmGKDXdRYp
ayM4RNpBfVLHPYUzdnV9jcoPrn2+yhZAkKFUtOYCJMAIrNQYn+1xpYiZRHWabGS8
XJ9XlQEmfdOxHbRNoc9oHmjdteOQdclWqTFGpYdkjetVE7cRMxJxMqkxQ8YNQZHY
+OZNMXzM3jI7M9HUJvT3c1YQdolrObgSjoFJ5DdwhC5bZNwUqEeMuz+uVg8tKkLv
ocfJWro7paFwgqOiyLAckucj1KWL06B41O1M63OruDganhplvE4GqmuY9/7qYs3H
oshePkIZd+fRphkNveLWmsLiHSzhDz1KC6w2YawfCZKSEKul0Udq3kojIlQRnn9+
GrVG+sZlT8XXjC/oDEmm928d4NNPtI52tnEw2U+b2pXs0XylOQW9ydl4ts6Vigmq
4uixqXk5JODEh5pFLUJUmjEs6va9mxisy08XcJYQOMUvy9yhY4rFhzlHFzwEYWgD
9IrFn+gwP0gIHqJQpAwSdqzA19zf2zA7ZlX3Z2+ONCIBOfdbv4XoFksHxDx5NNFJ
ChUCWVniZlAIZrahdWz5O3XS4WaiQkszc46rc6ZY/Fh3ed+8gZxVG5zgdjUc0CsP
6v4cC0U2a5ElUwXz+7I/6XohCbU2ivoaGk9OYGHQ1A9zZjb2ySpf6NC8oOssPiLD
0b8j2JnVLVPpVjLX274MrCNWNpqYENZmZBFauNPVxlvz6CWNAb74UGF1RRDjDS9E
v+H378oGxyVOA85URzfWTLngsKLMd8+8JkyKyHk2hNJ2iZIMRbPIcmFoUtWQOxpe
u9XZQsRmgn9TCeZVFfsWrg7pP6AL5jkilYsOXtJ+zfwQGE81kqCuRUkurN6c+tgP
srn/ddgOWotZqgEYeBt5bGmfSTeuhILwOGal9llcE0c5LnKQiLABtg3mVTLxykF4
k8zNrajmeVykO5A2dNZZfzMTOvsJFU7sLZMJHSdQycHIAqu3cLAuZcOhkSUcdE2J
EAjPI3ykbgrv3UCiKrC2VAKliUUnDDq7uabQw892UNs3uzYYWDZyv4wod0q4MxXe
PVOzCZGhhl3h7lv8t3pd6RdMEdDlSgQH5jFnT5TrGsl6KUGyhzqOsm6sEa/uyi2w
thliN++EkAgs69K5N7PoO1zPARGzjZ3ywBK9Rs0KvCwtIVL59U39qLbUsZz+kF89
gn94Uto8VbnyQxGeIajVfiM9mhLGbbrmzCUXMiXjIPZot/vBRlLcrfack1BMoFXm
LfCEvSrHyplPPVvr5YbFflGWoZUP4Nm2bk6gGDv993v9NykKb8BrQ9XHXJaP8e/s
YgnKG03XajQrylkgtXzrikk1RqZiEJEcH4fOaFpMm7bERqo7x8DP51cZpuUCu8iW
wBriXd4lbAVXKXwgevLeugpdQSETBZhf68f06teDAPRT9uyuzVhd1hvdhQVQXUZZ
YPQFHIby0rfLcwwteviMwBPHxV1RivnOl1eO7HdOnINSSyEKVa5QTPC9VWAdZika
HaLNWJ0StgQHPSgEm73ShIIMwzjMhJAj5FztFm3HnzfWLM+UtMXCFSMqW4pbA9E6
UlHWm0o73SBeaCl9ZUA0l/bGFss+oNFDcP9rEns20ggyPzdtT2K4wSIYGRp+RBUA
bK57lkAA7tu8FUV3Z0wSb6+VVb7zaxUIw44GNJXVhwejAS0GmoSkDdAsK7j0lR7w
8JgWaxNT42zfi+Uki64TU50hYD9QEmw1hiOGa9njp3NbRi13g0aMIFma30z8y+sF
QJA3tGjecbt7RefbYWPBToXT66Q7p3f8c317x0xZbxX/ABadcOwS8VvIKfMjBFgg
Iy2o0eTMvctfgXP2Tyv0/b6J9O59L6bqoNXEDRt67TUJSa8D3Yr7VT16pZM/3qgf
9HSVyhFIQfHIQVOX+qoB8N+d4f6tsjp/vWhG9BX1FVbbvoooIvhD3Fg9sKnm08Nm
+/+iMVTyROnebIH5r7JmPS3jX53SegVyg4Wa5X7p9HhjNqDl2kaQLwGSDbSrW2rs
sdZNQlxwd+sTtqiz4wsjpc/8rHvegVwI2VklLRXw+pDmxEAyfsQkm5wi78zNvvff
nkFjob99y5fVAlLLIH6aUQeDs+hXeWotTydCfSWQgtLWzedSNPTTqIK2XLFfUIP+
6GJmQFhRowvl62dWvb+5QRk+kyZgPXFUDEGlazeF22mz8sGc9E9Nfk0FsCLmtl3O
wBTAORMW5//+vBlEY3AEAruRxGOY/xDAjbtUJqjwJ2tki2GVCGYbav14u04cXnTX
7b9eSVerOaa/f22s4YuRQhuTchjYIi4SiXYX6Yg/s8JWmopSB/ISp6PePviTwAzb
M657hNjs1ehxlfcOx0KOd54rYn52UBzdSP0oY4lS4kicXw0M2Apna/sxudTDfCEF
ClVYfeaIDJiTQIplkQGfiCaKEto+qFJwTMuJnCET2/YVKK6dAlYesGK+VDW6+p7u
Hh/xQBJB8c582fLIYw2yHt3MFy7opigHN5K+Q8N5HL8TRCsbxnMw4ILVindVfNz3
JQ1LYe882M9UvWYxolJWatB5/RkhmsA7VBAgtCVcudVLfWkr1is8Dke0npAWjmto
QRNlyfgJCu5moahQeGQA3/Ca1ELqpAnRfPe4Mb+UsUhN68LDtsS7Z3tXvDD9TE4l
mWYDsyg/09cgpupxEcuR+d+DVlEcisX/Megn8uJ2hsAfnPAhxeuo7RKH/cT8DELt
xmB+BEKZXYHLFumQ3XAXlBi8IZp2glog1Mg+mFnBKS0+yM0XZSWdUe1m7fXgFgvr
RPE3r9LNf1ko2kt8NFCzsuFkR/kOfSJomCB7RhUkAH3rpxnV29vTlTEx+SDJo93Z
gf4tn4vaUme2Tgs1/uwHZ3/CAGR5G7eg48Fwn21YIY9KWetu99cN7RtRxIEf/JAh
UROUt5pQb2ngoW7KnFbZcP9xYfzNEbsyQAV82lWk8OcjZK5+e2JZVzd/oCOOILHu
8/gxiwFO4q1G4u8aimsBsG4rArU1Q7g92iFkqdMt3BSSzvXqTx1DygT1eftgBcLA
tpup4NMaLQHtLpRZNdgNAE30zmlgrk09U76RNsfB0NGIGQWDCRuwudhKHtiQhhJR
ZJelximjbmxw5DMLD9frb0QuB3auJ8KxVFxyzBWAuLkOC62GRCjzW9H2bu8qSfrx
9OOBb6v8Z1RlZk83SY5xQrywT+RBCVcGimqcMspMcMsQMp8u5r+AXLkvZJWD1Rnn
21Ql5NwkC6nmiZ7wMHeHc25e2Nn0TEPleKzQDjc1sNJyGmyoPmtqUPHATHra8yf2
hzCzGQynDC5isTRN9DFssiKg82WHLQNP+yblHcRYPCEofWEnykqp/talYg3ExzO7
pSL4QQRFVgE33tzEmLDBx0Xuzhr7gwcqPk858sKRInyfCgGD7MysDm01dnVqUoPf
CzC8V3sZwltd7vHSnYk4rF8MdFTwnbwzgftm4mTW8V2z3Uw6Oa70kQAIRaHB9/cv
FX5CrZRRYp9vCgd8KxpjeYjK2dzqYXPZKDGkSeidQrVdtP0l42smQDSlRHGCdZ5V
3UV6rX68VI7J8+5L+Nr8WK9FqpGlpRSNOLV8F5/fZPiTM8xzyGKDDedCyptyhfFB
lPSzrpaHq5CkRqbSyptMh6sVlVk3GUfbUp1vY0yIKlqilsl3GLh1EsuJkwugitS1
nmQBfxUuxlCJ8fSuTu6oTP4xKQByrRCwmwhE9VMoy2RNNZLJbL8Ln8Q2HXlWM5Nw
1U0Kc7rgOtpzsDsFx427NM9gfv64tGSIm5kbwlJgEVETDGgopD3F8PAsSorLewq3
enTwC7cOAxUZ+HdoLM5L3xqxkmb2GZz0o36gtdjRo6vOrlMdhBplSQDW9BTsvpGT
kinqWEslb9Obw45GCt3BOor9VxxWHG2t4Y2wKN1fQCt7uLXMFWrba/ttiGdKqGbI
Zivj3C7gSvxgpFCkRk0sFuxIiqjYdCOmm9sLXAIwUsJOlyvVZi2xHyYikCGxxll4
r8ZSYyTCYKLwac0nZyv8pzuHwEtu6IQTZMzTy1fC4ptK9HZwLGYU5WHk0O48S6LT
07iA8NaybgMHIR6I/cslgg00xsYmcAQ/arhtzx9nVGJXia7j3zomCkAKOhIB0X4i
Gv8Mbr52PNRNjKyuhs6pc8VgYU+QzBSirF48QIrfCYNwBCOqxYqRVEk9UWLHFXv6
DlRBMklxeULyLKofMC0h+OoPt8UFQPL/2BZILUkEbq6oNjmt6vu/1045Y3IG6edq
emKlAhcRRLjZDJ+q9MfxYBKZ9beMLqEA3YECL/D8aGE6B5+s7eq5euYY5eKyqBKL
zPMK+RtBWNYm+rkxKMGC3ZOzDfXnMgAYyTj478tYvhmRK+A0nyqHpKtn6/V40Gjp
YPKC6GMgXKDDJIJlgq5mHbQIDDVHZck3srvHnY+C7yX4v3ztLhKob0ZlOcTAR5lw
IjeURirDkNG/YQMD0hvbdlO8ExUE0tb8GYltP2se1hM3TLKeSTZ6lmP1ECu9BV1A
K6NYpP9Nei3QFOKe+V/cTlZuLv+KPs1+7UUlPpXy6jnHwLYDdNi7nbM2j9HJWFb1
+s1SeRQ75hYHoWlVv4KGCQjqsQpwVdZVF7swa/bZ6aWhyZ5+4o/nAywKwA6Lmr7E
0KB/myJyZX3dH2LT4LrEJzPQNlhRTqndfy4vf+WbjffjyeMVHg7FIKbfYuovrzpS
JaUyFXuxJdA5w+eHvX3k9nA8RkhoSG2Uh+j/2jqfMyRCZfV3PZULWFrHtST5jQyf
R/upt7zYpS77WKoPcDRmgi08V+smubp+RDY7qegMGtsK/rnlIb4dUIUZ7UBVbOZ1
CVGDErS+XaKRJGfKBSfsknwzaSeIAiqD35Wz3gHJNxDRZfctkW3dOxziW5DPto3l
YCoL/ivn1joLQyZEiPPgl8rmsTn/75QXD4G1IoEfFZOVA71GWHztZXMaStBAgIhz
cUaOf2vBTyvfQU08iB7d3ajPcbDgjnpCS1/9HDH4a04F/pq70xj0uZyYjFY1pS8g
Di87CSuwlh0kn80glRpx6bDatYcf52s9SCBftrjFb8U3lFo9qlSfpHLfx6hUJ26k
skiTXYPiieokn2Kd4YtsgS3Y9jA1WA+gzrROfZ1f/X8qVeXisohYj89/w7Vqeg2y
fAU4syrM4M14FXjBKE6turxN4r5taJzPBqGCXbr7G7ZingpmDgVUYaxCZNO4o6jA
lgXFylFMVw4vg6XZV+8Wr/YHXwGoA1qh4w/nxtJFvSA1rxuhKf39dI6Sekh324SN
qP1MTw8XLXhRydPSN2pjQuf7nC8t6fcleEPJylexgWUMcgt0gbNs81DyAuiNVsjG
C+m28XuOtt78AjfQd6/mqCQYKd6+262uSGRY7pJvsD3virMTeP1h/od2KI0IN4Au
P5jSe9Gs0mE75ZMe52G135dJZf4Yu2mZCmwYttvGVp360dpZc/0UrxJ6Ot3NJmEi
WKY23yutk76lHD707rbHoQ+s127zhmdMrMc6CNhsXoTXUQsrnzlreQnsy4tCzvMD
Dg3x+xqvRYCR//SoA6gOS5Zr/mU3cogzOJ6ADVAhln0mUGkDyvTO7ySdocQeB8hA
JD92FSSmB8RfuN73dzPqkK3+KmQBpdotX0qFSiVh9nUahf5iYLGPdTfNCEU9SFRu
bg500x7FD6tsfFvVtax+dM2rNb1XkLfObbpaNXtUKiay2ehu4PHdLlA+4cU6hudr
4PraMcT0WvayC7U18K3WaO98npmzM4LKMJYzHaGjpfw1QUK1tENePOtDT067pWMh
4lS/j4Om+fntjThWshAFEb+wjCGDAvsLFRXcoxlnFJRPgen0fzjJEXW7DnEvB7hF
B20khNVWoqlBtz9ORVL4YnLQ7ylY9AuVOWq8RQTVF8owaUnn0KuJ0wx7HVbCqYSi
iHLn7vZJAsY4xPDn+NPSn7hQLoBYu+eAgMcU+qkf7gr6mkxepHB6iGQvSYMvbznp
fUnUVojfqfnGFmdJr5aISvKkjYssFpDvvsoQgd9NmDrklrNmbmbaUe4hlJYjqh03
iFdygNYzcKZRhazaW/9EMchCUBZ92IocgqAnZehU5T2iMNsX219D9baBG9JR0CXh
pXEMuZYrbQPs2V0lq1j00MFz0W4+zrO3HjE8fejClU24xGKUOMJDghFm2W68baYV
6yi645b9qtMDXFKeNSuWrUOrcjWHZbjkc5hHHado3SdYJCXLqkZDU2bll+raiIiZ
58Ju6pzd9jGBLPNdFFzSB1Rh9QCc/9JJSRKDrtiafM+0AyC7QEZfjxsT4EyNvKDh
gOTvG9MzGvbSoylIPNEVTUG5gEFx+8lGx1dRx8wPGb+caPjQI83XU5zY55qMx14w
4JoxYNrS2MntI2ooSv/7anfQGQ4f7f1rCrieBhjljUFmhoqj+U9L04nWjrLyKw+K
D1IQT7zNoCVW3Niv2a9Hs5RmD6N3JixR9ad7TxZzm6BAPYR6/wsvmWwdxTlcyx1X
2+yEFynbADN3QWYVI30ThVTGjrdGTao0kbkfCjbzTfQaGLN/TBZodBRaiP6FoUB4
5fCU7Kk7/+CRP9mw3cvPXChZZB8+dqWdM1vAuQYvBjx8AqCuOc/yyAJA75BoIXGy
EcvrpudNrn0PHMzXqgdPXLIQR5JlHKyjRGxU5GzwWCOEQ512O9Y0HpvzFC/iIvJO
dVGvfc6p+moX5Gm6u24NIRpHOMXcr0nS580CdzM9qozrXOi2zY1gQPM7PifkZ9kr
/1u1vx69QVRo/Kj6lVhp/Pgj5HuMbsaupj/1aJLMUEZM/VC21E9H0fviEMMQixqv
5r8fhLdJOGRJpsZAGm01mIpbWxByrMAeJA28MHmympMym1NPxxlm5KjRPFgl0xUw
22DKSQDSXu6Gk/FJVAECKCqLtxOvhjzQV/gHqil/+kM6XgpWLHUM8WXVS8+OeT3T
PH4zdRM0Znu5Tvodjq9663xSSY342ok/fO0LHlqcDbxCrHiBwE3ry3HzmwlhzNAt
hieoetYAqBtDVEzUdqDSlbIAKXZgPEK8Zls8DcrJ8NdTffWMWEsTLaroY/8m1J8b
XtLZUuM5UaYu3OUe+QPziAWK9xrJ5psbtkONv7Y5BNXmeI7FB8yV0xTdsJUwTEKg
7HHcqpJCNHpV0U0IzE3aEyNRsS6jzaOasp3k07h2vrk642wFSBaiw9B3LcienB+Q
ncWFPrSBhw/bQiCW/vzGKRhnIkjt8j/AvQQmqhN83QwUdc8oYIgU/GTYuTAzWDjL
BmV7cK3sYDpPt8VKO5VS13bSnztKi9E+tM6/yHsKhfPKAiH/vhTwzWH22e198QYA
vYC+PcfSZdmO/s4uzw6tB0NosbxFzYVlogO++BNUILPDLIlwPSUt8WjYI8asDxeG
N3xfiNfULrO2inrhQ8+rVa9YGYV9FKss1DxEAnEnCtp1XOYG9yBOlNEqQrsdyUAZ
GvbjzTarao2YVmr6Qx7i4P/66sHEf2Bw+jRZnhf72p39lc9XmAQOPLYrUOCqurKT
Y04m/qvZcqNuKkMriWsHBLKtkEk4eZhI/Xyz4CNJcrATpj1PDnRyfCRrbg1O7X9D
XhpuwULeMmC6cUomqtclVC7r7xmqFi+dYRP/4G6TgJSGWPb7YwMiMLQdWQoTl/Oc
kF6ROTLGENAmTXWmf6/irLc+5Z9OZxmCm8LNvYJkEsXNrbEhREc+UmFSY7VwgaxO
YXZqoE8Nb7tdV3Ba/xL7Ug4XVrVHolrI6giSHYuyDut6NKx+sEpUVrl4cF4JQYWe
01LFqZ6wClLS9hzWElalNBC54PpVStHX4cSYCxXayK0ZWkUn7nepQFzEtr4WxL8i
A6DdmKMGh7D06W8olPglDXqV9G7u2W7ICwltACPbuKa3JgEVPYJiRfuD/AuSab+G
emsUYw90XfipfNUhTL2Tr9oVCBowyrQwaYG2g0sz3KNL2JQBC2VD33udp+8nFW0h
9lLRnqIxLEHjRz60sY+lUOp25Bob3WuOJK/BU2xYNOogj1hvBkZFO4duQMxDmxGH
4PgyQr8Zrgio7rGgwhGV0f87sUzt1rM6h7Ryu8b7g39LUjUTf/HWWIBM8DkpkXcO
RrcaWaG8xhz5FCHMiCAw0zqHlrJQAJymyRYWr5O5OJ9YELgm3H2v+77nl4FKkSbk
wvmJjs75UZvm53KZ1FpZMPcsfb4NjLkoD+NKo5XD40csDs9aKoljOEpmT7K2Kbri
pCzITPdG9Z+/1sal9Rqa2y8zB1kkXtADLM0mOcWIyUKUIl2P++yB6qqPpIDhReOV
VW3k352C9SnHjfPOGo/kM+GJTKBfW2leREvX+4NsiHKQmSI0Eyi0cUSGjwfrQyGu
iCdN78Lrl6D1526jpoxPZ0BKPoro26jjkqHei7ia3yGvmr6TWCCELdrLwsCFvG/a
ZB8iPLH93nH17Z5YJXksbMMZIThlGD3U1o54D5wtre40pumGueEPnD2iu4rnGdlw
eiRFb9+0T2V3PLCIaKtI1OmCr7vFlSWkNPreXfPMhnancU+hQLBQRj7KtS6KrgRB
JZJJYznyuiWFE7a9rjnYWZ1i85Vtcu1/aoJNKKhh3OSVpqNlE2cfyc/Q6MznHz3n
Th64VQ0mGzxw82Xt7TsrlNn5SKVi1LFC07AUtgKyjdnXKVg41rR9ivDgnK93NaAt
y5VvlIA7lSFEBI7NKOSbf3FPVLlGJOrbW95W30rKIa3sYdHI5Q5U/96PzaZKUwzL
/z/31EfR0C7VViy9ToLNrkdA2/C/R6u3XimdQRCi8pnlrIHiVkY9Md+eZ8Bnh4mr
VJCnjukIIsprCud3kzOQYxS1V0LpUpbxIHbNCtV6I2rNBfOJvTEGE4lGMuUWqC1i
vLH6Qb5NN30JcTHicNBU88KQnGVxidiDCbWbUmvw1TA9akavQwFATd+dORtxY1ty
qdBMTJBt/muI49BiT4cnPcg+DAwxjZH7GgRUYlZ8oGqR2AKPXpNn67XPFlStiM0e
5KrUlsFxZjjgjkYC53OBbgO/V81XCpDhoopkPFg0fVUac13Lub+pascvBFpTdU0j
Av9byn9AMaechRWSVOu6IDePpWqYeAxVCxZajiVeNMFMtcP4Nbnal26/iNsieKcS
BUYU2rIcB3faziW53TlyWsxIFbmLf63OCTDiOE+F9Ull6xf6VXHRWhSQ9HLXZ2LH
qvUobpO5r+bqojTaE8ovzKT5TgjL2pW977RXX0COUBEijs4DIRJ5Nys8iFfMxfUK
h5LhWIkOIkCuAWkMDsphFZtZGB1GD6ReDXjo4Fr/srHnbeowRfJ7L1WnuXk4fCTh
0o0aGvKBm1I5sr3Vf0hRVBYV/6mXg3GcNYc8U1RMjNaU9Om/RiKyvxgLioNAYzMb
jyIZxNIpy8qRFti8Po+xEVcy+FCUy7rE3LH1KLOSFM1jns6AHyle9kmBqybtPGyx
zMI7uRxUMCpxhWLI/j6AtNlbmfGIZV0junfpvCn7jBtBrC2TUiyVlawqcQXlfnCE
h8e6r6BwdBmv5EyapGAHiNe0L3rN1k5nn6ZAm806M+6d/v7JG174w3yKq86074lW
jiRR6WHIn1TG0oderQ9vKGC/tc/XbJG6CMXBzsWNp3RhbrgiS0n1uLQaD+DGRAH8
rscTLbY0o62BULt2JXWilzjkZ0b+crIzmW0P5EZuneV56eDblrj6sBCrgsdsrYoQ
PFgejcKNzhQSEfXASuOBF8Othm6ZtIoxOiS2CVcJZBnhQBXjDZiXpv3xFFI47fSD
ueocAquCZALPPb2fdQXrf0EKHsjWGvU8oypWYLUdRvZK4JxIg5RvxhbOHqrXxlEc
m+yJJzJrCCWdKZoUFptGzdisHPr2c1c+4zppFjtq8tq7XXcU7DAF647pgraIkVYM
zHd+xLbAHruGMn7GKBtoIENgmEtorxrqhsYYHtrzrUB855oWJ+iWx22olVb/lDM3
bIcmFBxkFE6zWQZsCnU+zZnIGFxAJNhDqCEKzvXJrNZU4k+yibhM8zDOZHguSFkU
WgeibABouiyy5F6mUAjX29U786Ql1lsKsMDEM802aLMlg8Oi0fvRBE6OD3lIhQDi
xHLzQquJAAAlNhxVswn8OxgDgHoEHBQSb5gilrg4B9D++KrswyUjS5nbysOdbVmo
YWdkSt1f9te3c90SisPQrPku3XzV/eHNlcgk2CH8R06DB3EBRiWa+Ldmm1qDweg/
NnNtyPjMoL5PcZ3Q1wEoPOWQHK14zvbilNyo9SlS5EFUBFcoxMIvrMSo/529HgUD
L7froQkzH3OApdmHhfB+FOs9etN2fHGd/hlAECCE/NYgjz5sGkRLYjlp/E9yJnqn
AxqKHIWDvxGcbK2gPUF13CXlAuYTxifUotNB2oNc0OeQNF6PGmI8OGVzN4nxVR8y
ScJ5YcemXi5aGi+ZAmzPgAlXFgMOJQPEE+D1/HN6DN27rv73STdrG6ZwsXdKAZyq
uwDzlVdO9II+DVdGnO9PGp3C0R2hs0+bwib4R5q/von+RQPWO9BIKDEqCWhAuUIv
ljFj0P55oLY6+Gsq9g6/9iP0vmrWlQ0jchAXQH++BhOcCkmv+JucokaDHxgVew6W
fDJK+CdY4+Bes2J2nuLaskPL5HVdFxW39sz/ihZQPsLnwhdPf5M7grj3lhPFs/SE
9PZdc88zvTcC9jSYIoOFFEgTYYCjpvHGwVqy4uped7pjTPy2aO+PDUOSEOfaAaZC
1m0vlotQ4u5pUY6FUHLVLRV4oItQb0fklZofpSPFFmlXv664NfNX6XTS/Qz7Qp6r
az2GBxWO6729eLiqYpIE4qRmAL6AtFl6woezWVBmSCAwTnuXZV3HtLPyhWZ6mkXq
Q9+ua2R6E6BMcbPT4WQCpqtF4qSCxyNQZeTbx+E2Gz5UWzxtTO66NIm8U5mFUIlS
Lcy+ETOwKacp/lJdp0nOPpt/iaLtFBOd6CjPBAs3zNcLU8qgLVt/qqJI3OKwBDoU
LzIvl0js/jCr3jrkxJHeZkgCAlQo16z5LmnG45kR4zAGUZ4BY58BSzzjzh5yUt8D
3cFai6ebqbvXsxbP4iausf2WEe0Sjqyzdjbt7r9aECePSu+XndJU9F2uvRxmuC2c
HxEau4mN+EOKD7c8AQQAMuax1Fmcp5lyoPL+2K6CN5uBfg/svTZnjE9v2u6zrqKG
W5pT2dfVZS4Lv+YgXcqISXOUUWO9iwGJyot1xm26tCT4XW08E4Th+LtUnj7BhW9L
KX4Sy3FyOXwuyzh24KtnVLQ3Wv3QINDJyA/0xpFOcVGqN6idzu+8vLaOmyY3JVD2
16PBaKtKOO+nCzLBt34f804/XAAmV11GlwiAmdMhqW4xyjk03Ei8gXLBjxrjBIk0
3GwsQ/zWBVhLyfkP6jRJCt7qwyhOLos9rQvMjzaACmDmNaojBr/5gs/LqeLm8v4B
XEAAT+eYqMCLysUxDikIHq/2oc+WEvMFxsD3FuiO9yUkWqCQK4nwRUATsje8d3Ji
rpaiGwGDkOmQQ4Lfh3CfjJw/YTXBZhkN45VMeN+GuS9G5Je2g/zBwXnbbluaxVT3
KXPITjIRKcrsD/9H8zF5yxbXyQYKDRiTtHyU65P6OOt9R6LnuTOB8qoCSHTmFuzO
pFAfPOqNg/rjamGsxUumN4yhfD3KY+Jrq/XBjgvU6IGuSk1bG4U852uPPq1/Xy8P
piD3MKYUPoWSNm6BIt4UVEG0Y6gyz//0umvZeWQSvkQ7OmTIjMK20AKFa9YJSZyB
tNYBstypfKKr97/h6P4EI5Pyzi3HTaznr926lb67i1nawn/kDDctv9qFoaNZyhWD
H3/zWoqaIDMi1hUmoprifCjnirPh6TYbG7G1E+e+y3yPjDPZi2oh69Soc7rQXOMf
iqAHYTfjzxBrhk7rd07HinHY9R5mCppPumvEpIAoFVc715D8YPTqFsLbPR76jstt
z2+o13ZUDTvD36QEPlzxukC0FAV6on3/TZluAtdpvGjxmyw/ZjKqqilKkD24sZ52
68KQ1qq5LkHPUCxtdzu267CJNjIAfSu6orWWP3Al+M3we25knl+CQtg83qN9VZV+
MkTdpzADc2HZqpojHuBC/D2+8CC6DEni+EDgKIJrb83S3HQn3UlbvB1CZsUa37cS
h7hhHx2m2yWXezAnatbexUaVZAJdPUd66LQd3BOo9VrHI2yDozehKGB4POKx3lHW
g6RxqJJyZqjcEeGXpv+Je5PCg/1mKMRItPEdrHOAb7i0Do2LlzD9eWakhN+p+Fao
GCXFMNGnomMPdvXuyr2p+atDslnFavQ8mO9ILQiwgCcVyW2oWz4/DaPOJIk850Gx
MdVfEqF7VC4li8filg/pWDsnomWzxbEyif1R449AyDDhxdYceA5iDYbGf6QIXRwq
3NJsPeWk+ERQ2v+iaT0/Eo3dQuheU212f+kpqEaAXMT6lIgB3LFPXTZW1Q2wKIGt
wTT+SeNT+aherqvboV4ED2Y1uq105Ca5/AhYVXQovJzgCYCysdK0gFMftAnHQwjb
JCGHUwCVjsl0MuTDNbBPLPs36IwK0Fk/Yg++DX4T4ftgxl82e5YO+gaPp7WuCT+C
T2apW7rnhE7KI1Je0uDqq9Fy/+9fmP9kNrQm4WVd5I5dayQsL9LTq9NZBeTC4eoh
8zRbjAWyzuSu7rDH7jiaxTWkuiGLPRfHl6+8DbrNGlgY/7x++iDkXnd0IweUVq0Q
VGWfBOtQU1aPEQckvnzd7jQDO65o+KEItSBHNvbKp19Ip2R8R7LTv7w3MYBXMPRJ
eSwJqjABSUg+wp1w1tyCTkN68advDqWLmtgKjiVTMZptbowz4nbTEQbWJSrUpbFH
4KT0mqZ9WJZOvaMI2AW1qXGPBi/fEGOSKG9TVxRXsRBUql6uXsNXzdpTagE/3qWL
8JzTEFPjs9vtfv+XBFfVeNFzrQ+2aSNfQ2eiMmxamq2BSEhfCGwZ9oeILpQiUrOp
JeOeijX0G57DsGll1WMo/AJspThH3zzecMBrD+orvZvqL+S4LX4CzwYLJXC6PJu6
IW3ASbxiT9gUXseVr1NrHypg9eG3eNeSqOqqiJaCCOpFwcScX5fj3m02D8o5iJ1K
WYALZ6pkqcLY2RMP/20fCMw6OPg0EAAoBWrTfoAqVpsLBoq3MUFRwURLpTRbyNIl
cJRa93DJA70tS9JG71pDxenRR2MRRaEISHPpldViXoyNSmP6rHj/nQek3AnIG8AQ
jBxNgcpyMkjLmjOUB39QCEOCzdBxMQPv6Gw3BoI+PTMH+6jCSRntL0ourp4frN81
YVctN/yPsAnrBubfzug8Y9ftP61Apw+9sHPkA4KQYfehRr0tU4CRKlbC0AGrsvDa
x6ue4Hxb8hL90OS37RINLIY5b4PbvE+8SZMQl8JPDRTLGjtabQnUzSGDGy87FBQX
1aG+/06CLI+gxUvt7wYR3PvpX/o3Xd1rEAOGZFFOJJllXScX+1TKiHXV54h0fl5S
u+Qc2CCBjOngs3YNVLtkQ7FO2Tl3NFmQ3HYeLTO2cmpn6hSuHiSych8Qub+IXmTm
YnI7DdkuKezAUAe05gyoljZ619Q+4xeGuxac4gOmcCwzxMqEvIkkAHqoZxnzDKcp
xW/LP+5DOmHep5rO0qDovdXoAfUs2ION8KSi//dlfEtnnvwV6h2VL3Qsvgy+uftP
lhevaHnqDPe4BsaOsqvbxYB7vDAI0W3jdVC52bMpgaMWPQJ8dH5oqS5BwVBoN98M
ff4CrBT1YZR0V+G4+Z56o52Xucjo1Uck4WNPHQPDrEYebrRYwMsjWZ/WrYkA7EAU
TyjQvev+Jt/2fHkm4bwDuwzt/wGPx3oswHORlXkMbv5eajoJUADme+ETFJBPWunw
FhoKC6aVcg5uEfo8NK1RWJeMyV5pBuZdptmYLktNn3nvFzUEZipeaVEJUL0e5KpK
6kJdJ4MegOl5K0KUQXjejze6bPTLRDCx7XT2J9I5WFZ8ooNEJ3uWKEPjYAJSZQ1k
CzCpSvRHAwV70SxkDkqL/rvpl8bCsDPX7Ub2/GeKT5F7nI/x1//7rD/fs3Nh1PnA
PPii33dUX5T+NJu4hBNjwrAWwwLY68hYwRxskcWPsVYZSDZpCLXHeeDwSn3Xynpi
VrV6FUcB6XG0LKEHmXp0v40XPpCCWDFcZfySUQHy0qxv5xcaHXM2+vI0ZdjccVVw
QXf7iO6xttuDi3LwwwFYPIWUg+mWIw3LoIiLj8a5G/FIUZTa8hypADa0kecpKcmR
NrIdw6oG4FRnEOYzeoTNTeHLIJIi9K0FZ+jx3faoi2cRAeRf/fdokfj6mViEfP7G
IfRI3COEmpejex95SGr4yCzVlQRD9kskxEqdzkDb7QtDfuYmbFSMTCq1ibwXY/PP
k8VpHYItfxrBhJrBsy6LHYLKCRhTar2ivvaLISqgz2dC3w6LCcwk78A9fpXrnRyK
0DTnTy6OKuhkNCF3CKH35czZGmjcE1v3KgmN4f9ylyVNI3twkZR/8DNMIM3Sg9D5
l08hPcJJCSeSBViB6Io91KrcP6Qk6HiCqADUKyZ63QTi27wJ/7nvAy//1/V3FSSU
JvgXhCC0ah008qdzfSs3I7Rdj6P3aaw/R8KgG2MBHd5Nu6o98EAEQlum0P+hMJ0k
ei62WHGfp380skQGZt5W3TYV0D23J5PF/WzydyS7GW+rpgjezEvcmYhOQKVnZBqm
TCarC3jGv/13XWU142ZwSC+YPlci6M4dPhQV10l2nAvzZxNeaoTv3SHYVmXTW3H2
VFwOEkWpJBXWkgl9L5NKdXfkmoyMzwl2iyTWYCSdJdBLptZTloomhYC9fHOQI+yl
0cdtUFkQqzWduBbEUEZDuqZCT5iW9SG86Wl/tOU6le4L7/Fb2alxXQ/PMSlEJNYa
gEyqLKw/OpvMKGn9Ua3kxV//ZyxCq6RXj4HPTHzbDkYK/gRckEjdgQktYpb0t3Ym
liUb3j38DUeqZ1t2lv26esw2kgwfw307DJdFTywoCeM2MiurpFeGZGdDeIUUnYlD
bfStS92YaXF6mwfBi9Fv6g0hi/cssqnFSzxSefH81DSxx4hpdcIpEz7CZHnlWfQ5
utIzYlKem99zMvMtfJjNA9qJcSMYFd+lhXnrfZ1o09PMzu2Ab7cCZrVGtlIpcYcw
6n5VHMD9IiNQZDcngzR6VUh1xlU7v04lsrzu/nq0ECwFzrl36YMZeogZSqWwPlpX
mUdVv0pV2d8z652GQ3CTaw6yjJdeXko70bxDWsBSYbV2qaD64fGzoTqhiqBB/263
AOo1ux/cEvJJGX+aj7IuokL/xtuU4WN3TxWhLl9MbN42yIArEuAUmoxv29HHmaGW
HpxMP5RUD64OkpADNEeeiBGEi4yT42l+HpOj7QOXPqO5NaNw5NVGM/vnkm8M6PEv
K5dEApcGPFYdzUcfzJq7WS6PSNTUdx/XQhKMs8xSpEvNNvJME7//lDIX/h35hwHb
5N61PsybgMmMHlzt+7N012oWlmhRfTNk5oHXFbt9JOdR5sh3Vl/u40ZuqzhyY3Gx
eGove30YOQZpiIsxETIA6ml1XSMs9vSLZf01JeVm8Ycn2kGN+ZkfiLAmRA0hDNuy
aIwCGC5QNAoZxGrNL5WJE2MOEfNWs4cuaH3KwZ4Y6gu41odS379qfBL5n0LW/QIq
U8yKEJB4lrbZ3Ao7vTocSIBpzvoDQqzN9DdtYwaunWI2vnlEDlREMQc5An6dxfxU
b0QKDyavJI7Df+X0LYQY8EIYXc7kd2F/bH9cvq+MypwSQj690MJqwAe6BnYUHE8j
CGOKCIDCw3A6EBtD+z76si6HYTtWH3nzrCdOOttJEpt9vZ4aF5FHL9n5KdZy2B05
5RZAa5/fPI0o0N3KBxkEJMBaiZApDQLboYxTKlya6zhM/Myn/cqiIIN3rGU/BETs
8ZPbE65FkjdeDHwfoLph5Zn4Ubk99jnMBhMV10nuyu79/MOUUMUJufxzaD7f6r2z
pZ52SA6uOMlXm0I5gMSKmp+aEel43ERxvEg8+k3pxEtQv6Dd3OzIARz9VknKLhkI
/eslImB46oNl6DmBfGDt8l+kkRNG//qtFi0kEE37kf0+g23jmMRZM7ln4s9xBuPE
emehOyQy9X2kvJxRCaBAOFDGz1e1RU/3dFNoaPszDT0p6GuMZ8AfP95jBoZyp2Od
skWMSHFaSN//AjBbGQRzc5igC+b06BOManiGqiFhWMJtfp4bOQeLIZI2/0pHMHpM
62RSkMXW7uQZbt6LpAHwWfkR4+mFTHG7anWy7/U+/pmMi2BH6BsWuAspuWycpOre
tXoD3T2ojUwRkbH3CLjwL5hwF2JLr+ToACsAvSA7MvBcOXktEvNVIKzu6aFBYXCV
103IGfhM8Rm/0BgHvQLurw2pxY0HNjxib9C42kaDXTA4IPralMvOdZ0Xpy8VXnD/
vZ0uXlpK4BcIbez7LU0UsFeqRlOpfplx9KmmyIjT3dFN7qAWxokEcSXWE84rGgUP
OGMXzDv1WjYol9bJLHghn1hat69vfPzD+orfvxemuXG8wjkcbbHXNgwDWB/qLnf7
Ilokb/sJMAr16A5XPWtEOaTtaKS1TXZYV0OQfw67nwk9ys+luo4RC/f8GJe6RYgF
ijDE1OmMzoYXYad52TckGmB4/jObl2yHZm8tC87hlHeMR5p5+OR3nRxAEPLhXRqD
mZXxY8C89Ywe7plJBc0oiJaOh+nNl7Wy89SFZtvGMP5++RLDeACE5wTH6xAdMtsT
tieFWGvD1liUYTLhL8t3P5BO5n2jJVTb7uMKrylz8GDZLkZPBWG4RfgPp3/Kkg/1
qp5UUjq5bmKrL+WRl2PJMP/IdEXHv9L2kiPkxV83iDFbuJTuSDpjdGjQGNFYKjTZ
8ajww+IehnGgaccseQ1tw5z1bcSa7FQAiCHq11E0A7tLnveCHZfHG7FLKATw6MmT
6JF4GBnF71mV6k+561+/yc/qX/p5jsi0h8Q6vsnkwiOBgtNSuSzFkoSNodvK04SX
LQ021UZ529HkjpV2C0d3ZFD7PfvEgz/VfkRFJ0bc9rhulg1jemfG2gqgTj2G74Zl
ua0Q9rMS+cBtg6eKWszHmVMCmsZmmDLo5GQHkCrJpnuxkqitsEAE56WpV2QNMnPb
9rv2uZmTBsMGToB2HhfLf0aOdolUO70gTmCON8OCst5GyfLDxXFOfyLxBF9E7syG
9LAA9r1vuGAg95u01pS7fk/hYwlJeZZ5f5BZvk72Zfoo4IoCU86ZMqZunP9dBjf+
VklKhxKNrO908CvRcr/ZAghqso8mQbdfKYU0ac+q7YnHasiwiJ2T+ZJB088eeE1E
xF6LCzqcvp7POSi4LLCTw1V+Zzg4Yczh9tX0XpS224vmmZo8LLJjX24WLEN7kFip
DswVi+cAxO0BfVy2ja5LRIOZlR77quXzEPsr/DwhE/7tOnAMuVZT6C5WbW2Gqe/n
m+IUPANo1FJvqPQbCzcGl6tzSVTL4ep6o9RHpmz+U09dj8BCn6/UuyWdZl48oEMX
u4QJwtzDhmo1l5E9QMEWXYQFIAyk8av29uVotgv1CQ5CncZVRsGugvrPxhSBIr79
hUu6EuBlg1Xh6XOEAJxLl7u3Mn8gOqQBoFPm1EjFpQOMWKE0IgXfibnkfD6zb9/c
LV7dobY25Ld7Wp1pcFxId+d+0TE1Qgz1SOUiKgU+LFMKeqfhiKeWxA5tc/wlGUed
sZBj+fPGakhz4/STtrfRATr8RZNm3w0JneBMsUQFLmbOeyBbPIs7f/SKASZJc7Rz
xfiy9STpLkzz0eMWIfFtCwHggnLor8f6+P4+GzgIXBUkQ1IfPJZBWgIqwbXtBNo/
jQvbM6FbYVrctxQdVZG9WlxILrdeR1Ni82HEBZDZpIs0iS+7vkXRKJVmEtb/aAvs
VXYKqV88Pox3P0KFpm5cgifcNbmRcNBPihaXwACGg5qtpWmncXBYDi+geFckpkxf
YVZlnC0EtoqKzK3KOw/G06rCkR+wQsCPSfHNNjHhLtGwg10gqKi+w0yv5IHKRO8+
L2a/sleXCZOcM5SmRUcPyvbvxmia5DPKSrH6XKgHYbytLZIjSWlfFgVM/p9NrN8t
MhS34ixkhNyeeaNTcWhkIYF+2o15lggiNpfKTDReManl8Nx4Oqhw4fiRN2H4OWqV
pIjKcMfReV6TiaVPebKR3ZTGAS92I6IVNrHAlALtsPYrjBJllzO+yWIb90foN4wD
IhE8yHVzEN3qrq3DIYpIiVAybbkGu007NvaRLMvQ+LFouSNZCfsmMJJXIsmGljeW
1JzXIxYWHjsDlkhxKT5n/wEmOHTKJE0bv9Lv9MRz5fnJTHVOR3f72cYImhPe3Ptq
+3JSAUsK5VhhXe4eXlgE4PZDSL4YVPQdW3rgPk/3S9zX2gKn9JQ6+M/m8HTY6TVM
q2jyBLkZxirQeSzhagpsTObKTt6bjvcE24K5SpHsd0idRL+QJFIA7+QL5ZzbCLt2
l23EF84Hn63WazCFp03ARVXX3zp9iKS6yqALOnpkL1NHZ10XS8S9ZPWXmDeaYErn
0bJDhqosdJ6JxLUjKSU0C1ipyaDTxAN6+M5ZTwWNtx0SJhWe42w+y1Aj+0yABvGO
WHyO7Nh2qO//iLabyjKj4CS0vAIYWbZpTWc9wtr/dG9wx1owQEzdI6szWiodgbq2
7+1phz6rQQXNDoksP6AHkBqJ/nyHVGRM5QDN+AuxHhz1LuFwNKFPV9Y/ACgUXnK5
PzjdLnZ5ySom8eAyUP0fJKeXiyIWuWQPVJt5lJp4E/dTw03iQObfn+wSW67RnQc0
T5xXemvLnx1xD2o/2BLcVnuL/kvlsiHyz4kDIc9oNJGt23Pbvgxm4WpI6wonAGDl
08krsfGHteUXaWW0AxI/IU1mtj28hxOSPh402b2EX8ykizfof+yq/Te09lb4UiwU
VMd6v02Z0zvsyVpCH1iyebTudWw1jOq1nOlJ8zuUt6uXsxy/bh4MdhOqOmcSFn2D
n/Y8OLKXNMdncAeJxaKP4Z/vX6/W5tBrwOBKAbE6RA68eEkCPxjENRx+WU/XgVhP
MfhnMirTRFjIPYRN/aZ3FeQd71URBltVa+3jcrur88GuWhBKqVBXzzsyLn5kQ27c
Yw+Ir+IoKfjvZRehjCTSUY8+KmFz7aoOR1vufA1wK673SFAQ9gKuVBNPwnltC29B
CxsEMCo8l/YtymKk7VTS6k3umCt3BEzPTZkNfFvGk1FQzOkoamg2K+ujX8Ws7iLa
OSRldZKxJCvs067TkaZYdg4lYP5DW+GUaXAWN7MthgxsqCAVb3+2hruFej8Lzsgp
vek5FznnyKT7NUCpcL903ma3kev09t7XsURx7Vl+NfRaqGsqRudrQn831s5msiiI
rgR052bjdisyOSQmFZZZfpboMgy5yqXH5FeSQSeMWF3BIdeH+ENsAfaFkNHxRiqb
7OX+Yy7JP7L5JSDawsfsvBZJARXJm4l2DGbs7QPj2PBEs/EVrcF/lMcp+mx1uS1W
tCHNXtG2oQ/UdgdX0qJvILYdwIKx1R/+6Jsb/mpDy0ejetFELLUDJRQ5iaTGUu42
yHymdEJ4RebqFDUKZ1s4DR3mq8wS7021/UosCS4KKrmJeh3/+GMwxF9RjWLx2CYp
SHoPkiOtQseKxrHEhbwwT4eqhg5MBTI88OllkJJ0I2T0gnM50AaOGW+pKoGxGsp4
FmOyFaZthkEoo8WxL/GE0TH0JWFDaW0up1B2lfkM0Ku5bF9BcuwFD3IVN+/WW9c2
cB9ZjSSyhDQywbOj9HU5v5DpmGR/NuyWPYScYA4kjakaBhCarluLB+rPF6llSGj6
5HBOjs5MYEHmMFSV7OizGV1XeTth+2byhMvFJ11MAi267u4Ytr2EwLQNaw5eLT9I
J8nh0sPaw1nhJLwg93ZJytXcWa4DLDn4f/0WcOy7vmjVeu7iysUcndQHLG/Q54MW
GPkDKUlY5t3SRg0cdNrJqNin3+BS1tSxLYS0jpvIYcVi509bYsAuC4JU1URDORxQ
QSKcKxvp+y3lZFRLbbgbpjwLku6BboL58ox+JizukuMIgpes/17VFeY/l28+ozxI
1IrFORrCUS/nSGi4bH8t1UxONUdBdDPHbReT54jf3wBOqymlXmdIFNyYsUploL40
0PAIRtmVUEIvltyxVFUb+lIC0qj5mPy6axnpkzc7+VCjs62d8M2ovrCaCkxlOSGk
oy603Sc0oY4damPQuEanXjvOgRDj2gWarY++uNWZ/Y6lDhzAUlZkdjDBjyhJYVVO
78wOp+2f7WgmhjyBqSTRq++MkOtE6NlAoUqWB6rwUfnIoD6qUGL3GCIR56sjptgs
gs3dHrZzOcIuSl+scAxJxywPk0jQkh9An3jKI/O1K/jKesYi734SYYfbm5ZhTUOi
TaMTj/X7BbHx3g1F0MzYYWEugGcKWLUegLF6r9s6FIWyS0o1EeY6vBDtOZ6wIMhO
MoqA7ArwxXuRCdR+ei6nQVEg5Wx6GZIW+7mI4Xg8Nqi29xRC2/1RM973CsGnHKSJ
4V5a+vqR4/gxVWjSzKf0CIjCroIqRAGBEwRTmNyDDTo5z18IuX5+FS/YsErmVd5t
ZPDsMshKZuFRMdQzLC/IwetdWmFRdqpvskJL86X1kU7QX++iF4fTAw7tBX0wwS3g
6vkUZStWDzakF9WL1IOju97CUUjJ6QbhCd+i8cPJGWeWaOixJiPL0TkIVZwg/RqG
jkYV64wuSQMuzuVlMlUSt2K0Rxxm4HZ3g7RLwXP5YQTwanOjYjGnee6WZO098v8B
PGO/kwW9x1/jvYAzEtQNw7l/dasRGBQkHB0lPcFNwToqzjVuCptMRL4KTM1dzgBx
cCQf+rcJArsJgt+j4NgFw8glgnOr7w3pqq8FTU0ZGNhQEjXrjvDE8Jw1lpvjUvmB
yb49QXhVPZP4pXVUIMSsKiWpHsAaKL8wtb9c5lqDnjzeHjFStC0b9CaeSHntTr+v
O1OAjPoto0yGYDYhyd78ocGQqQRUg6yNDq9c7scUHUEy/kbVf+xvEorAUzfjBjtI
0LbrSkZlWTt0xk9Zeva80sYZvorXRn8XF3E3QunSaW6lTZvFxIdqK9eVyJd58M3V
DLR7fkKRVBkkQRIEPFWnMLS6Afy/AjTWbvnjb/WqJpNARz74vNgJM/dVFGjdmvJf
hLJiTWla5gweRj6OLR1w8tJ75NpDx4RUAm4XzNJG0OhV9/fgpPt1igcmDQnL0vcm
7Xgp9YlwNPcyKJOAcjTKSRItP5sT052PXSHtkRB+XKeqZn4SIwvymEN3mZQ1CSmn
xJx9zZ4GLYdcTKzehtdDxciJzbb82a9QadtQxBDm/N0wnRmgCIDOBB0kKaooqPsf
mLCs06/P6TEswwCy6c26q2VILWLphUWw+/HP1NUljkaXApZpsySS8N3qEDawha6r
4AJCrFVxqkdOefxm9znO0FcT22By2WWib/1TSCPsp4V6wCp7Tst9JfNpOSMjUEhw
4XYRGiBsKmvZaeGW+ME2+GtDXytX57xOGoBwzJmz7NaPoVgNT4w/8rguTKEJ/AMY
sPqsvIBLIP8VyP3C/HaLGeMrszNOykA+eiaDXxj8rAsXXy7zyM8Q7Bgvx2z2BzyX
x2PCxC8M8xkeufPH4gGl4/X9DH4s1UL2N2Phuog2skjSg2Qyq82vst+QWejBrofZ
3ITEg9mN2wg0i0GJlIbGvaAF9s2o/K1z7Omy6Nh0BxzbWBz7ax0RuAa1wtMb1EKC
lwZIVQ3XpD5xZfpC1yWQfrF1MH4gMbWS/Yes+2gcTXvBXUPlgcOdrfyNwBIcb3R7
2f/jfgDm8AGPg/YMa8bvhBPr2TX7u5Ma88qdGdtKk04aZPT5X4eazP2sHSHYY+z7
yRmAxelOYzsptO28QZApQ5/Da/1rEp7yTIVAkogl+k0rd0LOR6jSm4KsErgPpNWc
6ZHoxSn/aYP2vrkRZ82RqqGxQxAixSVJLwpEgnb5s1Zu0TjxMELVh/ax926af8h8
4BW4erAO8n1eu1ezPJO3OfliEm/SKW++O1lOvRvJWGLZxFgRb0q0HV9MiWNK0Bq8
mjrsDwC7p21rWVqqyzFSuw2ArMfNpzZ67dbIZgPR01DPx6r7RCespVOI60GNyozN
ixLHnYSKt9WrOeYmk0ybJrqgGjgWHh1TTou4CBWR9jWgZxQHJx8wd5wQT+LPHyur
9xnrMLt8RZAwtB2jB1dUHXY0RNFQquqnPUIJt5OQgYw/P6i2oLH0b4d/gahrMFHL
/f/1JUIe9EWNcg/5h/+f/PPMnchEj1H3TPi9zqQTiyKbORSmif7bWnuiKsmkuvEf
cbJXwkOhz6+2T45rdNoN7/RaPGmMIHDhzqAB0I395UCKJbRY2y0hPqNYXnqPdPzF
ZQizVMcRme96wwUG7iMfhy+bN+RDTlSc9SPEPpV3GHGx/NtbBbPh/yVOwGRot5oQ
ZK6Hwvuwmf/KpxFKFWtj3les/pPiPt+5sKAUPuCuYsQqUsPvhcQyBY3pGO8HxO+g
4MILSx4NFNm1R8mnff5JMOTGlSruNsYS2hNzoCgHcE5SYdM9B4VMMnDRLFf0aCOE
xDzgB1dD8MUXwGvlRoXp2//AoH0BEGLe6jaSe/TvbUC9eLuywkxT8abTqcdfxLyZ
MnIvQ0atfSlYlLDtwj40zI2R6Nobecl/sWvOm4G7jPjw6/IlZTbluAzU27b4xqrX
0ssRHTDNloqwoijOVKjiXwlxkK+AA2ypcT3rbRl94mfGMXw/sWCpT+K9lVPWyA3g
fZtrmSaCfmJ5E0zv+Ub1ZiK1aO6FyoIlvxQKLD9j8bjv27RResTtX9+kf7xtQZwx
x3QbUaMMkKR1knhn6TXM96hwKUMzB4HwoxS8Qd60zbmIGnuCnFoygkIRrDqyPO5c
R4tI59wAGHQo14ll/LPJi0kjRhnWWq0AqHtL5nbhG0hPxlz+ZuUirRktbwrceWWD
lUIwHEwq9DmmOywjPHadSly9KRm0IF2zVBVf+4DnI1ieVy1LWeMrv3nOEk/ayzj6
O5zCULVWsE2UHCBUmM2PGUQhxKsZY9RsJngsQiPTpArSBvnGeq4WpA+qiPJoJnp5
rg/I4PuXoxlTAb7JQDQZfK5fItLh5wH18rOgZ6ByJazJSU4gO9VtMeSzbl+eOkp8
T28wMj/eHhXysXWaxGOVIdXa5ZQNBU4X+EMAEe/WFne/+Cz7BkZhA9AWCm/pNKS9
a9uT9UcGytxYrtho8kue2B3bjXZwfbzkc59G8Rwp6eK8uvcw7K1sIIgighH+qU0j
V4M/ulfvE4GfbG3L7gNePorklXNmyQLbGU7J1TjzflX37Gc6Bd3hNhRIREI/eYwx
3eGUiwYeJgmOraAKpVZJmLIwLtbqmAgjIyLw2v3JJpm9Z3bZmNXcMZ0lQ6P8bkJj
UFFEYNQanGlNfRD5B7Kxr328FQ40CSBxEyA6mCq2nio4vIRKzqi3cMQ9h5qYj+V7
vVJL6RI97z6dFtTbD3z1DgzQjvFXE7ewYSgDMilc1GRvP9zRImjGQ0qddoR6bklQ
EQjoyFcL0zk5h9P4lBPAKW9hgLNtbIYXOx5TwwlhZPWGSgbfcAf5BE9seQFU1WQm
5uqvzWjG4dCJxFGX/is2DfCABwG2fE/mq+jSe2VaEtxbRJdbjF5ft4RhvjuAKqin
wRUwa5a5KlicR+9GFUG4T2Kei2opOYUVNFPfgysY53OZfWxf+g2KbbB+X1bc+fJb
DBbrC8+R3xk0tYQ1pU0NhdghIk3YK11wkn5332k1MDjfTBjMr1sWxEpJouVuAf4j
koTEWyDkxp8ALlSL/AOSycF+2Oxx1vSQ0oHGA8fcm4ofbD3kWGRrtKQmlJj0zkO7
6ygZOhIz/qI9ijXek8neOm/16ZB5qf9TX/19/ZYVipk8z1/f0yN8PXyRQaMUTxB2
nAPpGhz0qd1H5Cr0c/PdmnPpdEo8YMJqOsFA+HjGua0YYHGUvOiL6yRb+iUabVPw
E6cpbMtHKPzWao2IbbU/wCgKIVH+MDX/MiVojeqfx1/iij2GCBpjurGCGTgfmXxO
m3u39oJMQT6+o5dC3TKc3JnBUzbCp+7x+CUn3Qn0b5jTiIJ2V3qPt/MkienNcl4k
OwxxOhpnhcBRN3RHuD3hvRaxm0VoZk2h0Hn6Zu8VViyJu8r+WEDw7hpSJtIGHW0y
fl5sTM3H7nVc26Zha+iQByOmcUqS9MrnX32Yjc7z3cxFYb8TM88qQmseLmDeCN9S
hPWg75KdHHSKidUqmpxt9nBQ8XOmm0AFwbjhVN1dOkn5j8pJk+/l1zzfRUQaeR9l
g9Eb7PPMvPuHhhuCwkNPNkUeIEeL7cp01QJ4sKHbovYE5wXiYb1GbhmjXkPpFUwI
B+I917sKbseeLhaBAHMtLZw/0wGWS6Nv3p2CwPWKyp1SrbMKxgws85t2tXc+LlwD
6N20bjza7ltjfb+CBvtAyotPqYOObpoIKFgfwtPAYBiH/wvB4GfELZ6AXNNDMq2a
T86Txsci3vDGqKNazRPI+Os3jvWCuLoY+YAD1z6KWWD1f1jJnTeX5zuydZyOyb08
oqu8JrRwvCHGWoG+Y2Mk0TeWt7G/XijiIEUI9CDD8sZ8329d3VGhPRoNiumRCOFB
3Fj93tfrlLXh1srmNC09P8MOAUukTOPv8nEEgijrg3jcoQ/XbjD4lajAHP6YHddt
YZXQEdUyz9kXEBpnnVuPo9/RaY3q/L5KEGoOo0OqojydiOHmza0HLZg1dAa2ya9D
m5L5WDVZq28HoKBh1CVh7dkq5ODrNhtcR/D5Ox/Eb3YUuwLNya5KKsRoMpjF9Q7b
Ky2UafuF/xiBIPD6ucW/lTDeJzZiffk9Txsrs7qKHynvAlVVXvshMbe4QQBT4wOY
LDv9/prs8xStUTQ+ImPpnPwV0ocG1mMidQTiPKYlPO61jGexUarYEr7RhDOt/13V
eVIssIl820VTirXkn21SgZbqaiYhBvIBTi+mmPnlgJRVptkkIXhdyZmA3GbIVN6l
BMEcbFG9aJORgmJB/RBT+Cf3tX0MjM8P4Ig4vp5EQsiKgis9kkBNIYjyC9y1n4TA
rKfDL4rjE3EfDhxyODOBBTzQ60X+VhtFusVhCXDIncdgWtk/MeyXuQSCxfi0NY1N
INMrYhF5u20o2iYRo+kFSkiJwMUUmuMD2cPpYG3bD8AUTkjP70THeYJd4sg0o2ZD
fkAUHIytjNPk+P4r2ZEsygzE1dwCSaJnkvCWkwJkmngqcwN7RkASFUy5ilT3jA6m
ssnipHwRoAIJXKttl9uZJzooPycm5jCrq8b002Vjcj7k03wgvDRUx4IObWFtkg4x
M1zvJp9TqSywVWc3+f3M70G26PsEUqD3jOCM7ta22jsnuMlfkmjNqqtswUSREH3J
FZKGpOs4qw3jxkX56P/CeiVYS7v8nUXezsoYSKKq+P8dZB3G+9SrDRd+ddy0dE0l
CxmrsQoPpIYzLevCHMT0fwj6S2j17yHA3AdlnOt2gIwazhvJ32igpQ/CBQndAOa0
w7qHj5G7RGj2Eew6bbdRAfnhdZ+8s6Vh6qAZSUBAdClksiv72gMzbal5pUPfEDUL
CI4R0gz8pjQsNaudJ6dBCGbsh6F30gcNnlmG6X2T00A1mUWaxGPzqJ95gQM8sXkF
jBsvU8a/8Eugj+jjWEe+1W24A1JHckhIQ9WOSBtLRZHmXS4GEmKngeYO3pGB/M03
7Yd2A3IgQV7j0Tsz+q9mTGvhBpHjWtBvHqQBbpYqNxfjPthP43+of2wZKBtr24Ye
d0Vv8YQVk3+cHtkUToU/bSOt6JRwGoYSICC/V8Aw7kmHMrUKHoPzxO9UKJQK/ror
bK1yOfbWRcqLrAEqUxkOuH/VT54uC05RYFcZTgtxOSFOYEHeGbwLZ2bGm8ALxgSQ
sXL46yIWCIDLBC5rJWoMAMKEwrhHvx31EarJ51MMBtYltCg9hfnq02en5BHdw91V
rhwkUm1SOqYiD2NoGu1XgyvHu/mg/BhqEWwwzi1L1vEZBqOP6B+dO5Tndsz+V7cU
PWs7m4Nl9Pv0AH5D5RxD7bkF45tyXCibe2XGW8zR5zVHmgDU3NlqH/N2PbuYkNpS
Nc3ZbkPiL2qqTuPjDFiJ0mvVPLanUlI5uaFEaxIqduEge5ldtIicRIcL760EMIDM
RGxgkYipBSCVujeTJ7KjdTe9geDe73oopbw/VNgvZAbDTStOokiBzWCfc6k/hxua
0w3bUITc1qLxCjONyx4HLpVQDzSf8Z0gWpmEfOcO0ZzT+yYyiZOVDmMCRd70JiDC
nEby6DBAORn8Hwsi9CYrPAJADr/hS04pdSgMmxWMFrt5rpcoWkan6k6q6xklfaw2
5DfUuBEMD3OyoU7fXabUBGU4QFC1Pp7vg9S1KdAf1r+XSrtF23AVG/2GnrxwhgYr
hwvA2Q+24xNxQ8Iim0czQKGWHjMTzCnW853v42+303ExmEQ17UrOKlVGGi9kC+0C
IbztU4wUwSFQ/vZIhJCXWSRHdsNEJj/8TAx7Nyv6AX5iaAvPGBlJlZvu9vDjPKqA
460A5KGdUPhdhivdRuHiZz1LyQ6AuPC9WQxQsnhcJoNxD/Hm+N5jVH9AZmQBhNxm
CylWODD85s9I+e5Fqp69MaOiEV0f2ovMzfXTKh8+QOYl82cc2rXH1+4wEeokGbX+
i/COHSS9sR473d/yXY9c27cApUptAJi3QmTNP7SHGJvIb/4d2rfuBEETPUrhNdEi
RBA9nZEhyeuHFWgRLFNR9ylA4ceJYY5aALFMpodMvorF3RNGpC0hpmBw/D493Ieh
LfP1ZhrxZ36716RD48wlff3vm1pbTsThJgLM00CacdbfBxYuqpu8kJwYfrBCop/W
KEcpKu1Gdq58NTtC60gtEx2wP/O2KtUhwJvfz9hgbTh2BxRjpF4R06YM2nF9Qe6T
IBIRLCDL914mNS93L1QlTFRTB+wak0g0Jwh9JhILKdqE05oJHo34JFYLJyFaqKQV
NmmU2CLTF9ZpLgAuuT+BqYiJwhiCiGK25GYaP8p/vV9MRPM+iseEPvwqew5wqriT
o3SWCkr48Qbg3DCoV6YmRzD9FVUbo1D3dHDLpIyFv4DiadboIq88PdZ9ZtAAAtV0
uSXEgjip1e4C8/ZKGKyNIsKGtb8GlnbzCzqwK3mnsXePmEss/Wcg/MnoGwpCx4AH
Hf6hIwGiZVvPkbMjGHKNf1yXZLnV3QJNbSx8AGmX/dLjxkRDugK9yk67CFXawUVZ
NfLS61d+C5zo5YLwYcR9RN6y1rp3n7aY13Du1+thgNjeplJNvBBOCIv/2rzqU2q1
xB01cI4paBB6iaaekr+D6IOMtabVDhMLfvd2Ansx0Cc79+sFWp1sAXqkHjLf/AaJ
b9E9DMtmtj7yGkR4D8S8p6Sh7IvDcWrBaiY1A9fnRMwioSALcDfiLwqB0EScS2qg
DdxV97Rssmr/W2DCMv210wTKjwnbyMFVSmQxmSfXM5ntH9vci1V7taN0p20qpwG1
y+I2ZGic03Zem26AkngOH4KhMhl2gZXXiItQay/Zdvuw06sNzvDyFfENewS+zEWU
8fj4NnHjcMQjabO4J1VdFoVeSGYjq2PlaP9J4E9f+d4X1LiU0CUyfljwIhzkw9Mq
oQX7msjVAfmBShvZg/upncxY3dEmoQ+Re8b2GDCxzIqbHKaTp8BCwVi+kVMFtRwX
/BrldMJG41b+R8lUQB+mxeMHGMHY5EwINIcQxcFSSiiCn9AXP+3LdboSMEI1Hepr
jQWpJ+BhzyH9H6HjbITSWdiP3QeUGk71cgO4CwIBtb8qG0ip4vhLD9ylnG+ialaT
HHSX+UcQyxjjk5YUKD/2VIr38zpVVpyQEUIZsWh2PRBNVeFYifjQQm0kWUiBSqSp
JuQcuo5Rgcf/rGH2uZ8PfrUl/qAVba2YT0/OPC6rQgcw8p47U7dfa9liQLkBdTo/
LBht3WrbB8nW9CIIkMdF2LC20LRGXnDSY+FHu7/qOm0BrSL1F30hpHyNTg5XEOEQ
5yLClAldNtfx/5oQyuFUxcj1p1S9uCFW4O63CaDWJ9JHlBLsZ+rVhi1aHlMA2cJd
FhKmJF15alMyUYsU9DcRyqW3XWXwQL+yYY1G34QefHYWH7sLbDmEGUA10tH6YrRA
idZ+F1AWkdAQZYVqroC6sTr6ce3H7qUE4gLJVrijEuWU1TQek5ht6I++KYHWvAES
8AL+haDtFCjiS+JbmAfbgCulGwTaiynbvWTm79jwz0YUEpE69Q/71V6g/Yc9NOLw
4bhQjsywT+8LowB49GRy/souIHph++qi0u+Dswi8hgOX6WoaF2cFzoVBbhOSk5tp
e6hmq/82+BuEnXmcpAcUYPfV0pqvOOuSwjeYkONm9o1LsYTtar5ssxmYzRVD7F0p
fEwAvv+0oyh6YH1y52MfDMIOgBvp9yuGO+/eppTX3OaM5sUnzZO4PklEtqtBNJhS
5kPA012EdHVX1kXL5I1nsrhUSG1OldEs9hCcQL2JjAUOquE5HFgT1fDsfdpXSsyB
XUz8LQHuWA1xOwKRgzKhy6Pj3F5TZbrU+ySqEe/L24keXBlFgRrtWDerp6VfqsYA
YgEaXTcJmiRw0jHfnAJal889MY7TJvgOs9xQj7f+SFlosNHDDX/yQD5qE2dZq4XC
h3xgDdX360z+EPOghVkyzBMXOz5Qfgd1Q2cvIarywxy06zWKX+50I+pi3Z0TTlJF
XszlwEXnXFeKTxGuR9cQgFT56h6P2vwJvlOsqSdQCtnxDIumesGO4Iw4LPq9bj5x
EhHtlOZAcu3m0BX+MGjrFbxhtzRUMD0O44oalZeKYoExS9MdNcQgG//NBLqlkc5+
nDOIadpZWLILJfgVlspFfvL5rsTdLnfC387wLDIZ6usjR9V4RKMiknwWu/vz4s0f
UotV0HP6poQ7a2NBLeO/Sq9iqkgNH8ZJejyalerEE1nUfj+WvUbUCVqmlHRBBe7u
GlNnw1dBcSVahjhZrITItnnuv5FbLWQvNICh8Zrrb5tSxklyU3tnw/+AeNqNwGyq
KTcPTyDjdqjfDT/Q8sZExHjuLZn1iwFjhkJSbtLaZNtl/fi+IUv2t0lRrU9C7OmQ
e+Yeh/a4BGR+G4/cQ+TJo+gTHmMsJpkqpy5pStaL46i3V7BfKdjoCyMakt3SsxQ0
J8N0E6GeXC2o63yWzQjlVoxfajqtA76bOcmhxIQdHqXmWT7VGHS8pXHQFDH63WDw
hxjJ1OEpFXiCvrynATLUtKmGzYEKbNv4yj129DR2pDaSAVFHcFa5Fp3lFk1bl134
pW09r2uXkC8ocKfKKoUG5IfQlSOSQ33ORa9CPg+9kYSasPE5lzViuFvwpOKy6uKA
GEO8zdSOvFt57QK5Jc7quCV2cQCxcqJ3eVaaO9e0M2hhHrSH+rbW0ZZ6OZJ9WN38
85rJ1NvE02NOtuLfsg392LA5GWuEdPmppTVsmIHhqIIBIZDPJOhtM8BQmwSLv9lg
LhGGljYr48f1zVNk0k7Xzo10x2QuaW3NUjPxIZ13XslO6tP16TukFQzqitUebCgH
7+537yC2UUUMJl6D7bkAMedy0t/1HyFoRSDNWLuMnvtIl2xTtTbmOzBn83a4zzu8
HyfIDyu39CkKvyOPTxOh60SpUw1+J7dNigYkf5TJVs+olCDlTvhjmCdIKigeyKp/
uh4vxdnE1qNvScje0azRzLhYkSzH3iaXU1N7alO2FbqW46JnX6y4RdsWggjjQ/A1
akTovzhezQOSkrmBq88QXbmaXR7GKEbfceDLh+9Hyh5kJhBNmjjWpFqaVbsp+Ges
NCI9xmPDAC01v6LEGNSCrqVWqn0DHRARM7HsNoW3VZgxSHq6KvWkZ99AvtvBc4+5
hDLIsth3Tp1agsTgFbchDSF6j5VtLdGrKu0EdAjSwg0AwfVHrpxmA7mkJv3c3EQ0
PGn49iPrJqJEQ9zbok456MESEqzL+v8NHTabfzKMN1jG4MKUChvGb+6vMoArIOzH
CVQph3xR1b9cxpbvYjkbNGVC8xG0VTzVxSlfHi5lsFedE7USEDETdhefLrrDxIHX
crTtSLz4llj910tcgIb8dTNfzzLNFpqQ4q1rqN7w4/w92fUDcHyK0RT+b3NO764+
G1IeAvzco7KjEps/CJUabHQusrUsu1v5n65Be4+COgJOQokN6+jn25gbZsMXxxTC
t7KPfqujMeMC0R21d1ffWpKxIMhWefqA4vihHaicd1C/mEbjpfvOYMSarkY0mNtc
igYvcWVfbO/mXOhko4I6TsuuT3vN0rrnMPGtGb/tZ9MnDNGA+Isxui27VdD2H86j
k83sSlxhy58PAnlnYVKQuQiqN7vqRxyOtumgtFLNAdWQgwEZzCYXZ1AnOKqlIxYa
INXjgNn5V/U2y5U7CQBLpuzO+X15VeQoIY1P/Mw/5SFRynj7pgd8O834oZo4g8oA
tWnAbLEJr6LQRQ06wewhghCY7CPx/y4IBl/JgNmEYJ1ISvqQUEOjPIXI1Ds2tNeN
IiHOMIlNns5TA2CBBZ+NJAT9fiJP1cusQH3g472t0u1DBKY+nR4GC7Kn5403XZ5T
LrWXKxrJs1FeQtH+9tDtNAD6am3Aadt8naUhIQU6XEYLuFoUerkFT6fZhkGiLUy4
ItrnXb/KBwTTlQW0ISyQp5botk0t6n39iXGRoOXeHcAkD47N/L80kBjYPTXVy9AN
dSkHljN+Kp8/O+JlLsyH1yjIki4LJ4zHSXJI7w1NQJrWVQ7vxYWBS1CGBRAxaU9K
36Dc5YBkFk9AyJCK00rcG9GGmiDAu9I0KurW8p/55Voxr4ZQ0mabTklSf3i3/nFO
sGo9ZIkJ0sqEXX1BnHAuiz0I6XmLiKfOal8HuKaRDnee+kriT8swrV3KWxcOGqoE
CDzN2D6MpdXK3zAdUn14c6ZhAg340KEfmCB1Zp+hpbaDHCmDUKE+4ahNFOlywBY0
Jj6tHWqr3a8IVg+iZdawy6J+Pthu50F8n3eO40NfBv+LLJCFlwb9N0RvUqfBZlot
mo2XlnUQWeAL10QJXZDP7KxCCwguLqFxCS3a8ZO4TsKYSY58AeMSYeDXeo+XXp0s
xWI+4zvoAQaBVgREB8RM2V4g3MnpgRJ3X4x+zSTtBgNEre3Fp2xkXbfPDoSYWB3u
g89aaRRiGBFo58py/oExsGpcks1MAXyEoTfIHcsJAevH8rK+glBqiPfNMwAGOs0X
Er+qskbN9OT0R8q4WXcVnUfsB02x8DqtyF1j8pejBZfQ8WKBwLimSDpbBj2c+yS1
ySob1Orw6/AhIQYT8ZdG/mcHQaC08jOGSAyDtIbZRPavJnBfgAI3cT4t5Dl+pRLU
V3xNKg+e0F/OARu2KnAUWKcEG1QI5Yt650HQubDiXy3TwVsKwxuv6iJ+ElpCwlK1
H7FeX6budag5NA2WMzVOom/+/mMC3pK+Kz9yJdIU6Ln7LnJ9Fql4KWrxHNPiKngM
eLyN/ztkMHkhk8v0U4ZiKKqkxJpDsnS1ML2vP8mJUCth12MkROJSde7xPi0IiaQo
lKOuKmZdPORIs8W+pRI33pU28Lha2svRhoB187EA3JfspF8hxySjNH9mdAT2GChY
wEHesCx7Hlo9RgoofZC+ohXqMRfFR5VGJUSI5QvMwQyMATt5ESfQkwf7YC9EQehB
tO5Za7wtAHKgQcb0fOGpibwcftHD6PweDP9tNpPHaksC8Abvgf7j7mR4scm9yb5K
f/m5w6Z20JXEp26P2VWfAVnJZ9B4NaGat2N5iCMWQ2eecFsp+OYUleHbgybxvoh9
z7Jdv7zUrIcYtM05MP3n6HRhQENtfio/MhMvzOJRYo9KNa5FVi+7CsODqUVMBZsN
uSEQH9s2ufQu3sS2VJ+gQbBvGPNK/YSZqZ80QTjIwC9SWyZqI8qQdDCyjzzkN0ra
1Hu6VXG4gp4vTIof1mbxIzufL6wJwQUE6qhB/NTCOHnUNsYwRs6TxzbAZcFGjQYc
Z4I6Uhn2TYOzpYlU1OGxcdoqlPYW4f8I8AQyjTgCjOBYt/Uxw4M++ii+qUGOXOvd
ctz5eWS4cQOk518Ws6v9l8VxzLsfgMHX411bjnOiabtxRKmtRD8O01vJHOiNP0ZS
iY7XKPEdsQiqY5U4MEkKJSdWZEHwcEBi0VMGAJBWe8QxqrYXXNpU1a3LIF47kOXt
pj3yCqr2IwV6O5gdSmhRVFtNtkl1tUpUr5x28wu51Mc6QyRnWjdS6k0WcPPUtM1q
jMVUWXO69MdIjya06ZJMpRo3lWB0xy6Qo94SB7+w/2k9uo1ItFOXVr115Nwsjs2y
od9kJGRLPoQF5+A9K6IDsdQrGFLIbE5Qull09S8SbsKLFUgqB+hk53KU+aRK8lNP
YhkPbXn2+mHU8SnHlVLWEC6CAGtIct6s7d78D4dp58Ysy5j/QiipbToPjI6dMItf
GYD4Tp4YYPGcuX5NLQ3P0ZyocOCxvfejZ/Np9qH6PPBGoIxEB9wuY7KJCDq2in+K
sG2px46bWNUEu4C+UgpHkNIBnN9JeAQenIgJKLjUDvESEpY6Wm/RosZtNWMYwklS
iqHCzmWZ3+AmJcICFNsetX3ugJlnXF1UWAd21L9Ui+PBk8tE0oiIp+AHVcewtsRS
sZq+jbhH7le/XshacKfMMaNJTJ8gSRAREy/4on6F4X33c/1H7yRcPh7MEDqB/k3F
64LmzGgYKCpj5Rgebq4zqxxWLzTRm9BoFIV6x+Nrv+8u4EPL/SZiXPFQMMJrZN1X
jrpm6Acp+Ia1FA9aaKEERGzdPphp5I5mpPc2uqnyfgezyRuo/z7mle8YAqN3zfnB
ID6ZBDtI19/NbDmMXXomG+JGzzFM78bIvDJhBiqnEOy8URYzHljIYvRYRceRL77r
+251pPLOnommN3M4IUvsTxoHJzXTAFUc+XC84b1d7qNKWnuaRtKkSFilnB/sKngm
IvkpypmKyrA5oeDj0DHHzhQxetLRPaceXn726nrLfsaLgW8MiHDey6X6r90+F6ci
526q+oBN8OLarmAFP1m/PabEE5CHuSL0dnyx5qtRmHj4WXvr/6dZF9P2H/Be5BjN
X1njlhexbtSOq3fr9OzYZNqdbHKqd8Z6ju68QF6ttmKHtFfuwDwyfnTmLYy2losQ
XI6iGrCXhpi7c0IA4rWj4YidUIrlFN6edwLlUyDrFjK3TGRE03G9CV5PvPaP2yjm
swjzaUrgHyLqlSp0WIOM3eJ4SgiGkidK7vy1oDeXl9srdYunjRn8HJ2JnVnLA4gC
3QhatEbM6Dv293nSNTxA9VjR0JyMGAFm5XfOf3nzb0w6pvyCGDccVDbLiyEvmTfF
rW8JjStaEPxfItA4Cs6UZIGSGPHHVaU/l09Gh2/qbJBOqD892eWuL1BWmWLi3dGM
CfNREbeUi5NFObW65smJEA==
`pragma protect end_protected
