// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
cMpFKBJjX7I816elLnYSxfdIa/GItp9SFzuAPc8vwX/Nn6GT4jRpXm/2Vz4ClxQ2cQFi59wSaRJz
JHG1jO8oGRmiStMk6P9IDEDzjGzdvvrzzId8xu5Jrh3NWlMLwbTlDD88pdDCiYyAKY6p90xCJVIa
Ty9bLhsFPK/8XolwLUCBUBvvVl72daZQ3HyHnPmXcKnGznok2p3UAR40Yi3Wlkuew8o3lOEQLokx
u7vECPkRQLBRnJ0O3NLQRPGJsfnrKOW2c4Rz6zRb9QIRh8UH6zdvqJ9Z5ynu9XyjL4PDmfUsQW99
/fA6KxC4h+v3hHteRcFVRQDXt/+NulnoBFuI/A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
FoDSaj+k0l8FBQpdYTAxSjuw4tPfkK7JsFgpDrY1CGNBSlZmrUAOTjBByk5lmYuxPpmtqlszsaTV
ZAlfsMC1VNVDO10xJQ+BnoyKSdyGLYYTxufCCRT6uDWB/i4xiwevxRlw3F38bnC3E2qb8CdH09Im
q28NmTAJmgVttuaS8jJ3hEBcRioJcyXVLVZKbkJtQxemNIeF5D0LJScQ8Np/YRDd0I0W0kG8i6rg
mGYgSXXt31Sw1mHZdXwfO3doKXIKcC7+woshgDT+DlpyXuToPNsHAcu8lkm+eLceuerR27DZCWo+
8aCSEExUXwLKRTDnk0Zhw/0DnNu/4qrcQdxzdgiPu3mz1Z1XW6e5cxcWGMxhj1sLUCqjvpkl0Ijx
BwcQtWi2aGTLchJDuCRG0hwX5hDbJ5UAVWxrrppAFk5G96rqApm0ENYFCLdPZO/6i/td7/sbdfXG
kqCR0PDr30S+tyV6TWqJZkwNj58lxMBu5Im64hcV9VWBXDxHfXWX0y/ZxBqYrfwoSjHGiGzk8rcy
Qc1rcnGDqVBc+gsaZOJ7hMgJbnTxF5WjuT3Ux4GXpGSF3NpQav+v13y/V5XOdl41KbPQPg5vrdzH
EuiQId80zr1Fw5IOwbSArpCfoVPgPLx39IBQr+6o+ByT/rIFsvfv3RelJb/0zL8SHsVwKt2x/k3x
VZa6DZ59Fp2Xs0kfZ+LjCTCVyIlqtNKd75hNCgDW4u+oaBhaEMOzAmssUI3nLYgNe6DwgjHiFqnx
VdDoh7EyukCPNDfwOUndl48xcF0DWy+yl9pOb1Br+wQGSJdRf49ly7rz399QnbyYmy54bGTpHnO+
ZwPmyeWnQiQaZyknsA5a3qJX2VGcmJIQmyAIYswi+qa2ibnhqdPLt9+Y8vjPU6eo2fJHzsLL1XZl
QE3W+7fDJDXxwJzlfkOfUm0zMB6UrcsSg3LCX4z3UQPKp+tDYGhIHLFokYyO5NWslva+xeuInU2d
ORJkM4xctlkTjdZfAJM3mTlX9H1Rv4cHdyzEqbJ+2o1En8wkdvDSO6nYbu5mnyvhpjNbQ1BdC2TE
FqG7CPL53K0+NtMH+j69+3oQtBZ3xCLs4YkV+iBnTTM1ZjRlFqK6nNXd6q0PKDchIaUMdOfHa39G
thkCS1GtYv26Bgui6GTsNBuAbrf1hkXUV8FJio8uMvzD/mPdO2dVzRxtf6/x1miTytOEE+bVpCAk
3uuZ9J1TsMtwU2eiMfuyyvWyw1CbWB3IT0QYF3uqDDaK3XShTS+kFjP83YN96pMP4NT2puliHiBs
kn5sbsT9FIrs/kmhi2qEuKX76RORtJwTRdBiZFWPjMHehkbcL+BDQqT7yquSm3tZlhaIBe3BNDgC
g/m+tXm7DLIz++G5pfzfEUm3hvFz+L4p3vTsdT+4+pexFyrSmB7LJmHMSyO3AkpwYO8s/3vvPoHp
HJh5GZwYZfBmhQupUDA1xoUGj5h6g1Km2KpwVw8bN0wf5CiCiyowxnXoPe0SJdKiZDnhHDvWmxUC
t/iOfQO6M6rojjmYgcPePZHz5etxhhpEy35HLdfKuzFoXuZvw2u5KqNaJQUmO2TpUij1i0GdAoPG
OhWOkwC1i6vKCnq3QPtt7Hxk2ntOyw6yoTxuR+GutDLVuzpVQrHPND5GYYf14L2yUFXXdZ77xwiI
M7NUDNYWOFilSXfhVc4Z5GYVgoB+BWsWO+Wb8tzaOPV2symgmzWi5DcIWs+3adAeyUWqH2dzP0R6
QyOruEAJ09d11ZmIYKkDuNqZP37X3uOoeM69VYOfrsGTOr7aanxT+GbkQxUQpz/CYzJGtKaeBaS7
STYEvhP74OoMi8P2Sz2J+3lGSLcbSKYFCthMPwKuac0j9LB5GAy6Pl4g+Un4RDNSrXHENYRxG8Zy
mhKXFVKTfKf1pxfMxBVESxLVKPohBdKjFOqA3CbWKLliV8KoDf57zk6jJC2mBTo/SLU+3S12/6f+
chyUzdww6+OtpO8U4+D1Suc/QhTRKnt6b8NAGVUUcJyi7g/zjkgxvmPX3hkoZtOftN94VVpwxu7D
SuYF2GqwEDNa6MJtIi6igtXEu1ChJOrv6PKKsGnl/PnhIfAt0EvfC8+WwlPXFTvAS5Maup4mXT7y
ybVQ1VIUgWe2l/IBeyZeCdLn3UOkMPfv4N6YvwztgoQT/uBmYjmDWi4+L34DrNgYloFFQWNgAoRV
QNvR9cKeknhPTIECkOX98JL8B2mo5Pqp7SlP1OMHu8zkwJC+9yVUT+AUQWTS0UZGVuc9JGqhbptX
qxACQBPd2LvAnvM/kf11AdV8TnovoCZ+u9ow7q6qArPntuTuWzKYA+TY9jULpilRaWqKuwTu73rB
rcBLgNjxfShtRPuBx5s6Y6dAndWBn/16zqLMLZkSMIgk6B0dssY8RQvkS3FabW65KEx5biQrl4FT
DB8gYqtbUTtXub+J0bPGn91hSeMqNrf0tEHm+ear8eaJ7ljcm0WXxQCjxM5nzYkm2fl7OWE/J3W/
Z6Y+XYQjP2RYU66avaDx/b4Ys0E6tUFGreQu00PAgZ1y2qRJSs3bf3ykv52aW0RUiGoxLy7A2fDC
88LOptROgAcopEIX7HISyDuNd/dCp92j8fklIyeloxEZddKSPRCTgUAZjG2/4qQzuf4xMpbASm6z
7YxRYLeF/KMpEzXVzwb3D6EnU7OYWrQPM8WbodowM2N+oiRyiPyhlsbWnLfO3Wqqgu+qzaNLROpw
UkMCiz4+VsV7LP3n6Sou+wCU29r5kZOFMtGqe0iCDUAOFPEQWd8RfgXsTWiGdy7L/4/INpULu3br
JLastFwvqW/mNGWjlxZYVFWlnvT6txMAJbvQ2g/bk63BQ8eqmT8JpXDnYMoQn9/si0UQqkPZ58q8
1bPGqOEAlHwdxhUTU/Z11wMrrn9zfNIBmO1ISETQemPCJtcN7JV9QwMdm83n8ldbhBrUbbsdqUFu
8ajmB92f1X/fqR1BZVxH8yoULqA62qALnrvU+6WirSTifhEL2R6jZWEhBHmIA9dfLm8rV5pEc2Nq
WF+Gf2SiyYa9dItOR5d8SPJPsydmFXRX6XnssT4tCJOkBHHA/J67ihd9fiAFYBzW5GfZh2CKSdhr
Mk1JcZ3QLtkKTt4M4F0E6f9PANsir9ZHLzAwK2zQlVuqoMkHQXwfOVZ6mMeqykme0hYq4P5/8SUj
g3JQzkanVF5xmgrSbJBfYInpk/gTf/72rCP2zXk/R04gDN9ae9/NhX3DwxgwUzIjHCqAMf2cRS+c
jG3LhF4nIsa7yZQcZjKKzXsK2+frvSp+D0ECimDcT4KYmxelr7VJF4UIvPjU5EnRjQXTLFiwX4cW
YJB/vgv02flYwBQg8naf9gfJhjgIjbqiylGX06+MSMo4GnD5HmNido4Qr8v7eTmBTp6vBTD/+q0G
aDv5IJIqDTulWFsZIQ37inPLkwhsnhYGE65k+TPmVc6MuYDBBUKU/HjVDxq7JPqN4hh+NItxmPp2
gaUNA/5+W6CGEVloeWdRBVxYzlT4N0/KHJii/tKaY2ZVctCVTTjIO8Iof0kiDrJ9O44ad5s3eDmm
qVlj971TFcVxnT1S4Cek2vv5DYoQgocncejlih6G57iaT/PLf54MhkhRSGfXhjkE2c/bJfJOF5qR
0F+XitecK+670jPzmrLYH5hhlncviGqOMCLcitGuQua4C8Ioi34Kgp48N7O0dThZMJ8TZxPU5FB7
6LUZuY6zsnPNxz3l9ryWv88GlOv00MSopYDFCcoUdo+60RL3u/ELrYFAW8EcV1vMt4g/caduBxPS
DoHJWs9+wvLwsOrHpQ1h16ICH6QKO29TmWokMc1Vaitsc3tBktVwacgYcHTPKrpaLCQmzYS2whNx
VfcnG13pg790oD3N58faZGdeNQTPKjo6Z3lEJff46YQPkLi9A0m6f/q2uSGJUwKL5n3ouN0tM+qA
kAuUx3b7GCrYJpnVBukUGG5A65cmwYAo6jTpNXGPhWhwFiWKdp+gF3+RWd5inho13HKLGyS8MSMb
C0gjzBiwHfEKhD2Jw2KWb2qoNAKmX3E5nM3ehBlRf45L90l0sgGuy4ZMI0w8U7E4U2nuApcQCHPl
puzKtk9PfeGz20cyZha0J1xpqGQuD9wV1vhlaJJRvCSLJCS6PYsw/gtJQQz13t1UbMQZYXCDl5K6
xwWOsW0gII8ztzo9vSM7NecsM7H+j8CuTUmjLnlMUnETevY+Ka0H5R0JB9rifzpwMMtZ0nGVtsJJ
+9Y5SsDNdi0/r6WM6VZAzPhVgWJ63DrUJHvSmAo4KqjCDGWBp3xMrt1bhXwHcMyFNqLa/aplloDv
RkL/f6Oagzd2zX3AW1t1idex89fjBWzfR/c6uHgowODGDXdtXVsbr4dDbqIW3QHDIrnEXeCynVU5
tIRjV8STVCcYrwESD3xCN97P/yXgfM1t/hwPTMfRqM5gK5CHE7paFRZlfrddEU7kj5aDxXqfizdw
tZMlsF2NdEQgql/iUkIp4N8RBlqBRacavkU4hv1e2bNs+8g8maJNSMBvpL38apmXatja1goXoZ14
MWWucb/KxrGqbuc/65aeeUv0GaD9RQlPpwVi47l1zSFABIEEewRSveDI9U1VtpVS5ChBaVhhhOIY
paEP+vKwYvP4Fg7Sn9rU5jBIbbQ4E5Lcp2izKAXrv1MfD88imGfxpZQn8i5V59ziA9TwUNdyNKeA
p9OKT/po9fYyqrKf3FwsE7IhmJ1I6Wi2FsDzL6zuYVQj5m0lexWHbSYYznWMMJPr+ZI1wS6InwGl
grjmd4Y55FogkJRYkyXw0g8Ty3aqIgXC6cjDNkcLZNkape1WL6ZPp4yRvKB0rCelLIoqqxJtJ4SS
I6Qh9gXA2dKuEdNdnCzAuxFkPHbSrsRY1liJqEOQchgjd39ltEVVHxHOzR7thBGjnjwDt0Bs8GEo
LThmHiQKwLYPSed9S05b8dDw1MwSwIh/+VKRmnSc+CjKsjEUx3a/TFrk8bUKHaJgaYZvrCjWo9du
CfIRZiQS8S4RtHo+yjs6tNH/DOE65LWzNCzP1uQ/QiAK4+WCN46yGePsdHNb6CsyLgZWGFxpoosP
oTOdqBlfJUQbl5LPG3s284zhJk4xwNPfRHhOg7xtQCham/RK+Zl3RtbEwJPTNH55/ogGDFETDwEv
A7zS4/bLf4wuG9+/WSsKvZQXEvU+xph47Y9ZOhUTPAoB7OqCwIcbRwMgs0vVc0MbYv0NDnyZTn+a
mwO+qdfyVjrSbhtIdH4BEfPlnEBQBNVi/3QofBo7GSgE/bz3XC7eMqYxnDtM5Y1RlkKgTL4IPy1f
39lrmobTtLIGepfS+ewXYZS3WibZdpnh8XNZTOSx6Fk1vUYMizuaqhRBJZLRbAdkB0xlVbcc0oIB
DyMg/UDxq5DRsp6tWbvNO1F2H7YP6P4pepLKFRERJulzKPkbeq3hxhzGV6nHanLPqQfovWxw36Cc
lHtM7w50moHDZbcqA3SwymHxjd+NxFfVNcb/nkDGuHbubeUvlb9ZtLz0+DWxn4fc/1f+yLz1eOsz
heAoXiquTWS2Sux51oguurIGRT/WPeuwoXwZGFt799ndr2uqyyVMHPvCXE1MyRY9vEWgcYUagH60
q+92SeBCivPhBj2pGKAcDFMlPWgnZSV/dmp6+LzENbO8Ea/Rp2YxfU7iyAIgUshHHVI1nmY125rl
M+WNl/pvh0lepISSmeMaeNLP6l+4lC6IiwQx8UDtM4UqkzhYVEx1tjzyV6DCBwAppMnbSqonmfWJ
i0iPC4elucIC13ksbh2E3GOWdmX5u2zt1bTJUBVMGCzkoeBapfX3SFA/92N3uRwpa7rfKGrSr854
7SIxBlk4aSkbOI6qncpJCaYjhEEBuEKn+TcLyOUURTWPwKAkkfoS5Bj3sOx57wtVGcTcxqdk+tJa
QDhXpuUNr4gT5r/jQqgihMJh4SgjC54fHMi4WFHkZvXosRfSinjys1UhDPDWhBZA94GNXiuxz14v
VvaDWaIoDWFfDvDd2EDUavPP1rSYls8++bgTf+GCT0Fu/rroFhul73iTW0rYzOfoZ8gu9CbBjbZh
sZo4VQevIXOORaupr8z+VD1cEiM+n8fBKr6ARPNy3BLywmkxf2houeBs621fwkxsXxqapuON7Vbb
Zc5imfAd39pts5t3RIfH3Dd+r8H9Zz0PXg2PslPJIgoio0/TIE7YEFvfPqVrKRLrq1m7h3u9b5Rw
Cfy2sDODk+dnyX2A9S1N5fGS0ajamBbjRFDQDm9tUKz8cjfCorZ3nzQXTNZmcKDMd2qW7fUO7lF8
TBVIU79v4ANVGD4nJEn6twMkmtyKrA8iuMMRfG93us7TINn+OShoz1bTVPQfE5fI5rOfBgSOntsa
T11o9Rt5IGtrJfxyFrBtbt6O6i3Oyg4s+NdIXVK38DGTOwElft+cj2CpJewke2EqW8rvd9nAF3P7
O3XAef9bfav/Nkpch0uv+2vqUGl2C7ScPmMzttt13+D1OmWZUTQNOu0deXxIxG8VoGWs6gCAXx7D
9AaArIyxe7ZSmZ9ugINSLjwWe6IIOehKBRzQ5ZFdzBJmfyG7gvWEZiumNSJMCmRErjFe+RvPAvP9
FAsVA32MCkBwJmbJaLzlUDAzeO7q+wips6SMrkBQ0nVlKpQCWrsPh8Cj+4/orVqliHijz4uw3FOR
FpK+dD9GLFVM8nbW6pyDMvjHGRE/kZFmGaYx5xsiBx0++cXUyC+t3k536B1CUvKgPUtk//LX9QlQ
gdsjSI+wgyg6bwnGVggJGibo3kzJZF/IuQGuxKpy5PIRERFO9QqxwXIyYbYopX+/50clz+IKqKBf
7h/qhbYocqGrwjjsI9eCH+b7mSlaq7M0XRV/EjKyOS4Q+lsHuAH7BsaZDha1GAZ7yDnLtcDB/au9
zzf1s+FO0+nvKGrMClYzxwv4FKdVMmd54OMJUrcvb8sYZOQx2Kf4Wa+36kxnBvUvlUM5F7/9IePp
ljhPGuHhskJ9A7M5irvtKQbBYOEGJSERiJFv/V8k78aXwtOsz52dUgTf0kKQJsQs1l7YV4sjYfqq
HIaF5IhQJdtOZDM8QBYlknWIitAY7XvO+m9MpD/Jr1ogXsXQ6WOW9L0SlkoV0kBxLvBf+SacmmhG
7bDhbWOKQDISIcPZsct0tsX+h0WFoWNPkzI9oo3CYrKxBTWTO7bDmINBIxhaq3r0hY6rJDh+oqMK
Q11x9bywhT12O/FPLVGSbGrBPCjNCF4dESZf8HhOe6R+GeTqiqOki92h1PxonKP8LGUEkm/htXvL
MWi2DboMbqi77/H9eUCLuLxUJZeFrchKOGPNZlD1dc7SlZiuAbr+HvPwknKBHpCha/aHouQVxfS3
2zFHyZrAd4rnLeEEIdQnNefxKfSnp/RieQ9HfKt+SKzUNhLXdHMbG1inVmXbIpPnAYe1pJ5lVsKk
cW1KRX1QaieJgIGBbQ8C2/zTg9ts8YniBAJoV5SBlmoB9RuKHbV9vvOSlBrpUy0mzDxgL/pJiJCj
tphadTw071eweMANO4V0vKnQ9MYL/4vyNLTUlb3eqJ0K7pzTmJkkYYaxubRdsCeTU2ipXKVloQem
Pj3FHSa87baSknnnuemmQHQkXm+okElMGxst2KaDUcoaLB9121l2vFAncd2Dd0WhPwwu/QDfLxtl
SRBzWTT22UHBBDSG60UX9tcRQNj+KGxwwOrDiuW8OR7Wbze9+MUyWM+9TpLcwzOiCt+ZOwIr2ZpO
meuCL3AIg31rilHBmZUIQ+S1Vk+yjMdH3oDSME+Akrl9rP8wKpXzDORxWWZpe2diIc0JU/fJV2eO
MGp1GnD4l1v9tMfMVfV4RM5V7pppc3+Zgqodmi/r0RTGVdXWIFoQ7y/Xud7yACzmLbjnK98mHZIw
kHKS8iKzc7O05aHJcrenam25VSLjXXNGlQn02b3fdS+n9NcSpYpU/7J6t8cYEXpDFGGG49KhOndM
+7Y2T30pB9l0ER4SdzGiUFjkd7C5ueabRUy35kN/QXJmxBhqD4uTuYsEy2j8QDgpeflFuCsqh2OV
fd74FKho7xDjChp6xcujX8VDYqxp6AB4Inu2CVEPpfnMRrIYYLyZIq1WiQxQGrHkIYFzZA7oSnSX
1VCjO2R4ngvvj4shh/H98d0eF2j5xN24Tsw6m8mQTDy+U3N1pzBnjYfln3j+PCCDBPvssRqijj9p
/92EHHZ02YV+cgwN+eyBsdJG3T2nqUtBRuE/qZC7UFjl0a3ALgEqM0KysT3kte/Vwl+O7oZvrgL8
UdLTqKHFfceJ7Y2/PMC5aWVB9CMD+vAz5gWfHugrMIvoPwa4+atLmHU3YYFPIYGfYKo4wmmRNHWC
tT26JJiCzEl1o4bAPgqmVd0LEsJYwWR8gSfQRpJlNTTnKQayf91/N4ytYwwYZAqb4XdORC9QdvdF
EyuXTu4c3smvPm9PR1RZS6qnIhUIrjqJrt35iKNOMB1vezE0QS6Kk4czkoZzRpImy3xGcdaHWrhb
aKI0Ugn+/pfgEQodQ3L+AcVV5Ek9TgHvbBwltanHFyJcSZh6rEsRd/rV8CRa1iVDOPXX41oeCp3k
xHZs+wSj7s2Cfc3r9f2uW19IRgGjEnk1bTtadOJun4NKWbyFtG2DSf9klhwyAoLeQtv10rtqlfHd
IeGKeKp8Tltuz5+fRfC6cucTbYIzjI8vG0n0WJgMinPpi9+7BO3xcJz2UtTRjdZKvRkLfIovuDm2
kYPxtwqWKivLV3tsrHCm3u/CTqsM2DT+6At0Qiehzt0LSouC/ey+VFA6AjRGPBmHpAHMYcA0WIAP
IJzaVJU11eM9QIUp3QHb1Rml/ly2nRxiP8DzxI2imNFFgIxTPNQd+AnE4HsSoB9A8qb+F1TptqjO
kmKNus9F32/otK5e3FrwmPTz2Trt9RgxB3bwkjf7aKBGNVnPOPpMXyqLmS1LSczAdY8Gym+OcfVn
d1Kzs+ksB8ig01t+pXyRVwPO+psw8s5cMGIUVl0EifLRrjv89AC3XsBHbG0EeMHEg4/V9Z1fJEem
VX6/4HgrFQxpHFQdTSUCs58hyZDk4nZBIZoORCDjj6GaQ4ravrDVw25yJHr9jZCjaP2d5LnCL9Ey
IIHNT+Tci5So/LAYB3EmaAsxCJ0TiS/Q2UPSVp1L0RoI6vmm23wxbTvvjbKqnUqKJVRQObU3MHln
RWX6oCDC4w8qE1vLnFioDeOcvfWvzY3e/MyRvucp/Yha61C4NUg2+IAHrgoKYN6/zUO03PSjQk74
XmlFwdMiDoLiImG6LCKXP6WnJX0PqqFw+nEw223eo2rifY8R7ntAGIEwHzlX2tQOc+4j/kmtdhIH
YVKNFEq5xCcMCw2y1Zqe3gUIdTjM/7fD6wIUPgXtJL7TATirHujCAHR99BEjcHJwTUsZTGz48Flg
0w32RTT5SNLShPdg/IMEo5hdAteTWOpKnC6Eo/V1djhkxRiwlcMQUl3G4aRqBGOoul1uMElbMRO5
dtMwIVJlsyCnPHUhde5S/5l9CxcdxuAGw+HA99NAGtAO6FwB07tj9sVssgId/EyY94ImP103C1Sh
CMLReD5rxmYGYwxK2c9avskXTzYWkNxz3hEZqQeLumpCfsp50YuaFWvau+zAEx/Cc9pL6YwCf0iD
+AddhSkoVbY0u9IzXxkdIAu7kflp/A1hbWYThdWqyKPdnX6KiakUWgJxGBUmvmQu5Iwj6M+RPizs
h/9dRuUgFzDtReP4qJnibCe9rIjU8RY4mS8QfqHeznAT6azTbSI75AVcQhLs2YbtUmk2iyaTQqCP
ZAO6EvYcRHI2BhPf7mJ3gwerFufNpZmG/p9KpC0m9feW5wLEbzeFf4JAZN5iyoezOHIG7G2wdGQn
xWBgadyiV1bdmH2VmSXHZHtiflstaKDZ7zQDmHChMQJRyOPVE29GyAHq/tin+bQEwPn2+ptDkmBC
r91R49VqxmgJ1bgjA0jytE21U4CNwq/7Rnl5Co5CJ7xbVQNX59Zbb6JHj+X8YiG56cI1IO6yB5ha
CWpdOfCUeXuRbat/99PYYq5jYtwvHMSu5yMqtVuhQDsjfIFuoK2L8Q8FmxJCZC78eiG1aQwHyrc6
OXgTyC7l6Y8I7/NzJrPcDUiaztgW4ljjAv5ltH1kUg3TEpyb03jarnW41O2s+wEUMOxBfrvXgG2r
F7yhnSZePU7Q/eXXr0WFSqa6RtxZCIatzppRhiTeCQoaLQQhsqcuXNNKk9c1/09bhTngEao3u8bM
OV8+nIOxaxtzhgolPY/H1SpGwP8V7jEiItVrxvf9zUZPxe8E3EynXtOc1UGwE6q/X5O5hYzuYORt
C+dpbgKkDmz4YuqJTre6HfchmvA6kF1fY8eb+mTdp/1ySTKfQzF9iPshD2AVEdFM0Si6uUbJf3Qh
tJ9llj+w1JjSV13sTYcHQAdhfz23gE8MrVwFO6DjDttGGMzaIyv2aLG0H1dSFrC4GdGOaFmurF+2
lFDAN4FcCcPjVDKrVfeAMSeQ4aPy+mlSvg+apdAsH9gynCcqVP7tBPrOnJ36cEToeRBogCqTgR3B
NfFJHawx+4rf2DaQ4qznI680A4xRHOt7mfBZR6csQr7OUWoXbaiA4vsM/PD7+a6INrTOTpYr61Oc
CaZVzwQJDsy76x7XDXEK4ad9e0tyFY+NezNZ7R9TczdZs974XH0lbe/R84EAyKzQIBVYzfoZChZk
wD/vnJcxUwwng8xDJTNE470M8pGfqHw+WHgL3LtP657Su6R2lHtaBZnav5neXKSrmHvfcykNbiH1
CLCamM7yl24e03FMaLrbdS4aOMScCHF6H8oD2nt2etzWRoWucKPt0TaIIVgpA/sKmljgAEHK65ou
ZdsLiTkoMVJ7c1MO8/HxwxBH+h0Cd+QYLI5nFGikckb0YvBgE0y4Uo8os+QwVITKr+vJkymmsl9F
jQjS5dfcNnTryebBPnv+rv4dAdrpWKE42maDM0jxiscNTCd1vOHxuBwz18+V8HrKz66iWTAynHIp
YMveq85fgV+iDZD5lVfRZzyxIfT40L513p38LXvti1Z4RYhjJFfbPhZrsUIusgXgEk+0j+vFkE+X
p3yHUMBDQOr2PnFRpIuuFI62DHx34U1u/P5EVsbwrMOP2RF5nljFJPygjkjqGyVsC0wHuEVQZQkF
HbVEDTDbjEbY+FPBNpi50gXxa6lp+rJdHDGT8YjGr4+t380OLYsLsTKrKHZjXhstHLC9EN3XJoOa
E7XMADR0IXQD50fMklzmgOGfbwcNxGVcO4ekDesBQF4FpNQTRyN5YKfTBGMSLoaduZtXFFvS0D2v
5noHoz8C8QozxUwKPIcDMeY7GdkdZIoNWmN3V/YxZtsY4EAO8pLPue/jnoPUepaJQYHHNGJSuz0M
t/FZOrJ6n2XL4upIRLuNcw3aGeCci6M/zxdOKd9Etq8VFlzdLPKFpLS5lLUDfcFoit1kkBB/ADYv
JnY7BabyY045PqS2OzMlW0eGJX1JRajxG40bZbPX1iSTnyRaNJVnGnmg2DfSib9wjUSO7CLeGtjW
+gNgJn/OVlSDAwz75Y0OWWx3OcGz5cVY/VdPpHbPDjBwBAVe1MRxbEXCdwTw4cmyOgXQ+6rc2wg6
gdhnek1O0s/NLtea5njAjoa2+OrmZ9oQmWQnVIrp3pTsS9hT/Fq7QCfU1KMGrJiicqXgYwtlot9a
L8CVikJtOSceLYPfxQx6RSRT5sUbT3yIf9vhdksRKKGuTWFx2p/7sHrtlrsIrQmCmj9nuqfqhQ2H
36m+9SjFdrIfyzr5QCICCu404tDQUwteVHox214IdbxhDqp9PTsOdUb/qQBo6Qvw3FnH8ZzHD20u
4ZQqs5pOSW+Nr76u7ibPcsG7p9IPx1+Zq+d+cB2V2/QB3I3gIFhTpXKm5DsOVsnt55iNips5i0b3
wt/iR20yfXKqtLIN4RLXNZbI6P790KJjfr8u2xq7k7j6etIHtev2xvmitZGUVRNg0DN7BlOKVDI9
HvT9VX1pF721AYyJ0gpBjLhMS2nYyUKiBsohOhFNsdpnvsKuv/HRlLkllC9Za7RiMwSYTD96gcGp
3T31DCjcaJX6qXdRQZyDIRZuwscbKtZvLHD1J1pJ9aO8czjVeqgnMfuSx6sVeDvryr3YYL8hvAek
k6luSzL538HQ+bnwPy4VQPBXIKKmD0OmMwzBxggX7a9PXjdx0R5Up1znPHhOPmFQaovcWFvp4Sg1
istOQuwAB7rbFk7xeNl2+xdqzPCk3hTLMooEODiSKOTnoKO1xtZAX+VJbVeBahTkEm9szPXGEQzI
7zHgqsM4fxSusBjOwS/wH88KYsV6nPMJXR6rvWOrsjP5EzEe5eEhU+BuAVDEUYBlqsYeNLmuz9L9
eNJl2rczlxlf8LByffXQ6j2kZMqhjOLWxaYLPslVC+96QDQsb/4MSPpTw3ZzS2JmlyfPSaN56xQ/
59iS1hiHWbjNdSRdz1MHwSqm9vjZgmIYudmY2lTeqaaxdyu3EV6vyPd12/jgTgyXVDCgZiTyfINY
b1hHas2prkKEu0HzNNTo5KSDnp+RqNL97/sbLH/SuEjyesx+pYOxdaQ+ZpSfSGf3xx95nJUwATyF
05ubo+mn9K3yOeViFWd4ZAp5mBOHuPw3cky1guYaf5bem+p7AqPaXcxTJAHZN4nWn1/RMuAju/mB
Kdn6g6wyuFQPz5iLNwGui3svnAY/Jd2UkGsbqIGSATHHsRbFnSSSsuTFVzc/kAC8iYmVWkU81qfR
JTzdK12xxJ3/6RrIoLcdt6rm4q0s0Yl++LsXwbJT9S7osS9MCFYbUpupWNW819DQYyf2aKv8CQdA
h7cxSKH2XjL1TA2AFaFn6b19Kdavtx73Pk36a0vtdg6P0yL1NqIDykwmHI9K1/eIFrnUJEL5BTpM
Cb6eNnyMK1mu6igjdfydwgLj+xSNpiqoomE38YskUXfsl9xCLIPSmRrthLs0MHGxcD6pnFrMvTUp
eiVGjivEvdbXwus6hDN86L5nEuH7rJHG2cqO+O0O5CtOcIzbZZtXb4dYPOssWnwHkX3cPq9862Y5
WoayHTSJSFbJh4sbANrL8vhFgJIlqgaDAiEP3d9Jxn5vyQiQcYJqiWJYgnYkmSACPSqoEd3Oj7XN
RTWYaxrqSodCbV+08u9hmW8mpZg3LYvwZmgoFn8c6+Khv82lhxR58Q5OqJkZFrex/7l928JAHix3
rG6xcsAVxRnatyoYuhz759rphxntjWfVGXPMFurXJXE5Cxu90cuOGAdbAfVghpCFzInbPaQr4hD7
kz65lS3kWO3OeuJVBpthG3bgL+jOzadwNgLIPVyKtKv6+t8RWKI2oZ0wYZ6VqA4Hfu9uc/Y2MWxB
ZNuW2/YyEyoXjmJSezCPbJxAW2Pw5VOvsshhasuRin1W/9xnYQs3cIQapzIbpAQr8NtMBq3Otrkm
jfgR8A0BVhjV+7v4dkLBQTwU0Kve2ChX5bqDx5MriT8ehsxqNjHMFqjeGsCu83Hq1ldItNvpX6ze
qeL6pwZx3v6TowbMbmtKwMhRIgW30NWbw+acBhX0A8/EOR/NCVCURR5qbVENB58RI+y49RZPzc3f
6LZG83+lBJNb3ieCOtJF2FY9X3COyW6/7CVpge6zuunFf+yNPZ4icyJS+KKaOfduiWYPSHMGzxQD
aqN5N00HbNGMByNpI/mbOXNq+cyWghxp0Nu/CsexFEYpDBYFGS7fAVAPtc2V/UAXDPHClccH7jnw
7Izj4LLdLC20R71J0Odx8CK2OcEItEyLzgi1eO7Xt5/P0kox/T5aJW6jqWDiIh272ePbjf8y6QkL
YyWXJmO4UH2PuNTeMRkYmL3z7k6Z5BtEUVFAljfzxUIB/spVgfcUE927aHSRCRlndNm3iZn2rvuv
pKolX166wLFfKDnB7LefzrQMRve1xoIKcli/xXIf913j1kESgORvmXwiPyZtAXeZsxzxd8dZ08Ev
c1tjx3tMaGIV/+wQqvW1fD229plK79IQqqvhj/Ji05+N0P8ZrnuIGe3SvKxlSOSNnQ2XPikGpf8A
/vzLE5DvZQgNm2UMVfwYFyhBl9voKREUHwFw6eBTkWSimH8i5w4PXumIbrQO38dHZRJxli2tpIzk
7dH4kHmQjOI3sWGWyEeFP2OTFs3y0YrW3UsHyP3W77g37K2kT3A30X4vlZWllixTnxzGLxytjptG
yZw00hmODutGyxnTZsM4r76grd4QuO13pjkLzvqFJtfhxO1/GvTEddXvEOKu6TCYNAg24C8m27B5
VL5ggvCc2EABfDNOEkv8DzZ5Xk+4Vkp0tyDf9bL8T9mT7jYvaekNwbp+PqRB9A2l51dPuM/geF6N
cyNyIGYXhdm3oL58D5u9O2fr7U4TWmp1jXB6uh21LCP7t7+VujEbalRxonmM90nwC/VM5FVyo7oI
MqhCf0SKTH8cHuS1Nd+4Hma24e/mr3qPqfERDExpRvNW/0bTAYW13V3nDKCvJpa7HNh8RhLcUqgy
AFOXI6eaubBL8jeophuYqGVpTbV3WsHkWs8BEY3wfUTQMhj0a31HYWLTjk7bgKRZLcFMXwQAlMFn
YE16hLamecwO7Fll/YW8HBfZNAXCbSMTvR7fRXBriwrOz2YWcRJy7EH7stJA2RmSxs03JoULGkba
Zsy4HnNYUXTSr8HF+J2Vso9TJIQxn6mR7uoSEJ2rEwNnL7Xs6/jOF1GcBTaAbSbwJlrjSO/DTxOe
U2ldo2dYXpEg9QXfWOxRZhxrpVxA6iqoH9Yyl4e/xrWtWmjSNH/iYiWjh7l9QjntfX49A9oLtPk8
Io9QwYcPj+cqqiL+gg9YCRtrtV1kj9+yQGyiigykSwHMAnF4wMZ4YNVCvxzGoU6vTWc5SFEoFVuk
2q+RQnUYapCG65mQh4XyQChUmu5XCGQjwkQs62XInLQZeJPoPG8GEOOZ/5Z6bXGNtj971TSS4xbJ
foI5cD5RtM3GrKfy1JI248eBfj2As36lpcuNKKApvt3NeaghwtLaDErDmxkPZu6ml977+39F8fgM
BALRWbBYR2TzaGLxjRuDK/ooWb33WPAbDixVT9Mcp11BI6dzFfrsa8N6apCjpT+Is4DXBch0BOMB
k/N+g6P4xAh3WgDxOnQxY7iiCtdnido8j6aax567dSgLIqrBYvmxhPzlpdU8Uuqtj+T98xicZDY1
CMmgHHGMgwA3smziFghItNpxMK1W2tXTftNeRT23YlmpUuoCZYdtk+e2sVxtU/IbOKhz1DFEaK1J
Njw1DUuxkRU+ViuY4uoxUsTlUuAZSe5FfK//Y/cprgkQKyoxEJ4HO4720AmGtd19BYh0HRhtb5IF
2KhkReNbKV40ZbsSib36qsN4S14ZbZnp7LaZglPcpET8pIfoCY0jjax4nTQbVOh59MK6lO4p3OtC
JGO5n506jjmZ7RVs5QvfTHInF/FXNiO2pK+kSmAwaRS1NEzNVbYKONtTdnyP7wlQ/Xt6Dg48tB6m
/CkTn4U03uhceSeCaXEIHr/tRzcsPFqEVT08XKNxkwoY0udH8qELS46NR0Rlw2Y3UOvMQqMwRo9Y
HdoCdJ2laaH/jZxqBLiQG91pRV2Xt0fJeA6ldZWCf7eToMjWT5MBhuV5vqwVky+DOj/Tk/LgO97H
B3rwCYFIgnwBKjDQjprOGH1jMkoA2mAmyKcBOR0phhgiC/LkKxkY8YkZQpyDLESPr3opo9TZ7gll
lItVdDKNAIZ4r7QZ+UMrZd/T4kk+pHA+E6JOx2vslSijMyJLbV0Qwz0BKIsfzzdX1sDJ2inkOIZ2
99NDJ4eS3ML5FZLWMA4va2KLniZjBBwmBqqsUTQu3qs7ryXRNHq/7dyZ4Q4wyxjB6KCBKuzopdRE
cHUp1ohypYUXwHYWLEXKpZ99YzzWy7Ujd1x91k2ptusR0saIevmTSzjnkKQQjIrqyA7IsFxXu9uR
8ldVMljKGARjCvZdgF/9WesXcVjHN5MKupNKpbpoG2gIGPSTSVRCGBHE/SQ/ry97wlHeNf4wxKPX
/3Qyk9A2930jeMxiNeBwR1v4yQcImd5ac5S7ERg9qM1fQPBbak0Ni8rmECwk1G1ZGfe9AiE/z2QR
GgrNv9830dzAjkTj7JaIfHyfjN3Y1RQt4fr7qcyE9b44i4Sr8UVaJMhD3qIBDOIWIzFMQsMDxDxy
lwUkcz33BJzsYKAnGiNzPk1pwMGCJWuf5eqfzPHrPj20AOgQVjyL9O1QFLHTEekJ/uPXGUAl4RPw
HZ4g36E2ERywfcevkfvm/lshIdWhXb84GI3Q2EvwKacsSOhXdSxFDMfgu4kj2YpAdwezIBXnknyc
d5ZETkzIQE3HpcS63wSe6sYsV5MZm3pQtmCZYcu75SeVXF8oZ8RUKx1tfr3Mch36V6ju7IxjQIcl
g9H8ZLhlRUo1+p6K5toZcqEgrNJSrYxRetMLYh5QdPNmfdDl4YZ3pwbFWmMJoas9ddG/dPpPwNXM
OL55nwIret+YmOp5iH494mXWDljkUX4K/VvCanXyDhZgPfgSfMfGbnYVKKSAE/47Rs8o1DbvsR2+
i/5P+Z+ayhLorBBNftccvbWzdFVLi8jDUYnydLUzuJ80leHacuX3K39Y6kyUQgNZaAbYPFrx5gDV
0OSexAiVVhLv52K37cinxAmUBT+qoqxLzJh7jl4ms2+UR6bBnkB1CnpjqAwfzYYRqwnJOHhnOmuM
TX4eKt7/MbSgabPF6uscF3hpmR2cdbboT6WwLXRee6mg9k9zLqjuF0HQCZf/Puy8/5tAwYYIY6wq
CZRYXDJxOZmqgXXjiFokp6jgOCGbxHxmVyuntEfx73tH/L5zJ8YsSeR5AJ4Uqhh9cwBRTGRpxt1Y
4ZnM7wYyy/bwQBNVfeBZ9cAK0S1apyb6MRZjGLKzmuxaflzbuCrwCx5di5pB3WrgmC4G/KKcqFc4
6MHnmsffbm+oG9XlVH7hfHWDGD64fUl/XloJvp+WHostzx3swUhDx0WJsz3kYZSEAK7wvfGKmp5o
6YJi8ZW3C1wDulFcWwAintTYCAA5LKcU3RhQ8MzsQIVfHUj91ET7m9I2/OviY2wlfwkv5bp1HRES
6yne/9ckPDIdn+QqDFT4cvm8n4eGRx3qMQuQ/2HmDoOVjO5vovd67gTmip9XJaa0wgteFJmWJI4i
tZSiAAjaZAt2W0thKLHv7HXo/izXMIcMw5T/UBCAZgaR0ptP2P+vBQuN6Ooaz6diBZzicRidsBKM
my4YlvxASF6kyWwpT104Wr/FWVvACFg4YdyYRPqINB9hBSQ/V5joQDTw/bk4YqOCnIGqD3RAOWNW
bkXy3J364M3q/SvZe5b7I2FhDQE+DyCO6dKrJSiy36y4aeYi25+wOu2qsnTaNojI29e4kPr0VOHY
0a117tDFgM75UuIW0KpjmvPeci2LoerrcW9v0rLGg8bCjPcO+lGqJmwtWs3CIvLa0mglk4VaqHuW
K2CQHBNMSz8+JdKsXqbwYZUnLu5ZFLCzadApAqqXyF/m6RfOxfiHnTyvN0Xk3mlIR5Q5wQX/E6MI
PQxijCY/MTipLD4jdpDYqrDnmcXE+YOFHY4l5y8VFgvphixNRDh3r8TNarSQXgEHtANLz7znVCjv
n60hNXEgIqza+t8OFIJcIyEM4ppbcuP1+FA5s1kL2XOzDyY2us9pwCKE+1g6uTcMyz0SwYWqcnfR
uWFLf4K5haxHijUqp8kF3V/QIBCHuELSGiOKWnwE3bZqP0h6Mo/cA/VZipfUC0dfanJzKu11VX0m
lqiIWs+1P6LHJIu7pq7Dl0r470gcgZ7LqN+5QQ56Z5HQfabOPpATJvNBRfpK2LC7gmxp6RG9fuR4
vR7DIlyE0dyRoEN0S0J/n3YCeb/mjsbG3W4pBMSQGEKObGZzpYv5r++5mbkF+Cl1AuLSkezj1ZkO
gJE59eHn9PKLapH3ttbTeim7YNRy2AhLUyVVjRsVvrFwVPd+n8uc1PsvdggLxyBhOupWiA8cffip
Q64NAjBuY3Me39EZbcA/+6e/1/3UdC8qK8LcQcGI4o6kUKbWGZ2325t5rzd5WZgnQ54A0IXftQGQ
ZScwC1sRidn6JpypwlSFDjRN3UpphbCqwSjjSaoUFKggQ87KkCac2EUU9viPQYio8UaiSwEna4b5
f7j6g0ezRweIOp+1GUg8GMWIKeY4wEtrMiXH8NXf5+KbK6jgSuUiZvaEYhAoA9FEkd5dFuMIbgCr
fwz1h+TwVUVYkPip2c14E+grEA8cGDC6kQunmWpmepq9peAJogZ+uRntWjK4+5yKlxncYlvXfUjE
hh8JBNfUZmOiHSXo/eAnDNRqIzekKrRmK2zkj/UFHrkswlBglMZTY+whRBLaXP+WgCUj5Bka99Z8
MMDs1JvckYsxDRrV/xEDB5+jbfavpN9wGAo+bz8ynmWWSQNafOeA9bCbt6OIM9zT4EKnFof6QH/Y
ZS/eEMRh8zwIhSaK9kuB7Y2XVf5aVX/7ub4y3v55K5FEpUk5HKqFq8JqLFIAuL/YhKcJWMZxDTq3
HJmD2qPmQPp1Oukcx6DAx2bcBbEZcD5Jm6x2JQeGIseMpU/CMOI5YMG4uQ5xSpTC2G9KmYbs85Ub
aIKEJrwbUeJNcmdREJsDD3389lZwHaW6nemcj02X10OIIKdk/BUuBVGfIp9f+7tDfig3o7l28lG5
tgzirwZ5oJDqK/k3CRhDUmdguHPQ0YTtLH0R083Dm7xE9MEmJ1s9MKSPmCjxmjoA7jCiNI3txGae
l+KTBLAZSonXXfAV/0uxfbenJ7RV5ne+TbBed8AdoZotOkUl+3OLemeeRv25ad9+GR8cDLE4jYz3
bys3baTIY/HftODiw48n5tPoaYEj+6VFVkRxD0qqWiWP7x6K06xiE4X0khnX+JK+wdUwvUuL4fJe
mOcKGxVbUOURjMOUyjzfD3iJ6QI6ID0AUggabiV3CfIfnieP44DHLsPzGGy5aSONRkk3G8CERHwl
wVH5LfBkszOiQipCTd19muoclimDDL7KSmm+kQKAet9R7nI1n0Cqphv7jHyFcVJb93rgPvg7f6vJ
b81GB3E4FxZDkre+mBaOJqLpaDfzod2IGx8qOmsQp9BqmowOF7KR7tuMEmYr6RjOJENJRqjIlZt9
8EyZOVv4P1AVFo+aBE5C84VaCU260ruNHaR1ln8CdskEJNB0fg2rj6EH5fYqEVS3o+BRE/LyMy7G
PstKcJJN3cfxwGp7oBMU2THuyEgF+aePDbzuVwgzOE5geLaVK4rwEX5VOlEPH83SXLJ36finbTT6
+7/zCa8xU4jQHBwVamK4shGrTNrOzGO5PW49z3wtn5T1b/GR0KiXWDT+qi3oHepxiMjh4S8eLXT+
aj15MgKw/ZnTINrSIrHiMx61i0pJj7i3l/hvWQl2HJdcSslBGQmaUPVLWrYVon5aJU2d0BT3NXEq
zUPcuUB7Vvo3yCe2GqCc4pF7IDH5r2WyAqreOPWYN6pUQgA4WxLGp/JL0THvX8zHElEfOhECn1Nb
WxGsBsnUEOVJoxeZFeGzxPB0D8zRi87LdYH4PvIyO/IhnKLcFkjVEClWTRARgUJwP54iNrgBTTAz
YfspOuwbFWC/FxIkTv+F/qKzFpKAe4DPmhUJr/4Br/+8S8vQyPWlatiIMfauAqCu75QGQ+yVWbpi
BIrITR12kWtXC6TejYAXlmTcit1OJx2m5wPrgN0jkmpTiFAVh4Sj3IYMhuAwKj7xlq3diXNZtcnh
frx+5TOEpVawVm0tf3wS1A+WXPZ+mlqW5Cwv0eZ8jsfgmew5rL9QGffHpz8FF3B0ax5OkVzh3vrV
C2TmXECB0HVXDYBXnl5jPqKm8YBKhrEQM0d2MPBBJi5e2iddSbVgqiW0Vl8AIyS9593rvEkxuVW6
Hr6dUF+gaZMmLL/siIrN2G3AoECcud5Rk6PhE7R0phZNR2xufhQtzsh0eOnZd1i4+nY/X1r8hJdI
shvPW5FIHouaDOtmdkZcBwRqw8tiRj8k2v8HGUDYPvP80YjSWuXc+5gDLixHGdfpIZsz8emej00p
i/hLACaSylczVsNTg7lPLKBDVAG8gPJvxU8K/GmMM4JB1d21CaN4evScaheMBY1/vz/SDSmJx4O3
WfGxQpuKkFNlqyJiclBVMTAIejVOCEJDnXJ65FhBlu8zux0rZZ4AmGnZp8OCN76G67cVvo+f0g8Z
fF+7nJWRvowKkcAVlC1pArdtUx9tb1PH2QQywXsCqbfq3EM0Q2psZzhetrWaoPNFsSXjST/W5gp+
aF11Tn8vDZZwUeTMaI2kRlmc/RWed1+gRSGdqpH/FVkTPeS4+EqsziMfHqH9a76A/m23tmkyXQVx
WVdxZ6KHMevY5cS28vKB4kkn0LikooWdT/Be23tvMTLwIlIQOItao3awvpr5eCbXjbK6ec8eS61K
3K5P02Kf5WO4rvo9hu14xYs5WzzQOTF0geJpCsQqVczZSH/20qGlUm3kNFfevIi3pHiqQNCLpCGn
y3vnkw+s3X8OsajoWyMILY7xXs7v2eZ1kj6iuFEin7sr/1dKZ7J6dv+yDhkhlTePaYpM8qM7e2b/
vckCFBRdZYPmvAKq3Ve+7/c2otvEhMkpI79jeEjrockWXdAIC16gQNmdMlvPxqWTdShtQAfpUqQJ
b18jsoCURn9ZMbrbHASIdj0l/mgn8zPzthoaN/yLzkKWHsYGmtGsRXlgoiOrLuCHrqFO25d9sDea
hmfZ2F81ImLtiaw0PmDzNsfQi6/HHwBM2VIizqQz1ct62Fo4eSYwEsJz1RvN+nH4PRF9croeNb7X
uwQlQylB+pBf0nlX2pAF7AfmbYjhY70TcR30W/ALH42XjjoXtDlX0kT5R4angtTHAuAe5NIgNI8H
9lpL9V9879U6kQf+eTL3ttU+p78X4W9KE8IbVX3RzgCI+tgZJU+3PHtTRljEMALdQvXQLXZ3QVyJ
to7sMRWsdwPpq1bG5uwm8zmU+Gy9yIn3LbrjJFGyZg1j0JFP+wEkp4VJW44EKMJimKhCdRCKI6kn
SwHXY+fQDpMCBvwNo5byj0OOK2ZkHZ8c1G/2Kmbk75J1utG6uhgDL8nOdIwAVuppXYE8MVsoD/bZ
fDz3GPBjcPEMCZxmu7ad1B/nnBdN39Lqi5CCs+NtSUfBEidQBbMUhnfZ52mTj/5muMR2u8AvoWL+
dtfhq20wiDBSLAG3kDO9eBCcOJCTyeqc+RKIqoV5owqEbdK+BIF+dr55QpLHyVNfNy7dsVOwR12s
zidqhjcrla2k36Kw1KaxZA75D2HT4zP/+Hr1ra6z0soo7RmtHVQxV5Wbj0SbZn51zoUE4oSLIHWT
vGLpKStnR5Z0Zt5xmdnZ5Y74Zo6lQqWhN0++Nhp3tgpc2fHujSAtTe9fqjLDpg1J5thazpf63q2c
UewsvUVOHeuWrsSLry1xCg4+UqeqMppfv/phpDyu9//3MfJHd1fh4NuAl1pXSknDDwHb77ewRm83
KfDl3Uxj1HZH65TZzzdp8yeUCAonIlXJ+ef7lYi8e2AtnJMgLbFY5CkEC19rPeKb1ml9XBilH9np
5oUyCZbaWufIhtcbgzEifHbEH+JQEIZznya7a763hcIeABDo4K5MIxcJ2NKO1KOdRprnoyjfntqI
OBvbtjOinhGoavzYeGeWyGAMe0GA0MtyISpcLktK17snbTsNOYSzK4FmFqZr25Iy8n7k6UQZ6v74
P51FsWrEiah8saGHUTR5rtM0iFlW0dRWA0LSvTH2mcYoPuSv9tAEXBr4K1XOrKhbicLWeBrWnPiN
Vsuf485cVl7MnojjGvYljbM2ESpt+TxVpI0dZdFQZf6wBdnapDDdHxkcP6cY9J2iOTqZYAsvLxg7
moeWj6T7P1BMxu3h4D147ksakSGP0RYhu7xxaBfE5awuomYa8fEohXpp+wpesG1RYrKJd7Xg0NUl
RP+omio5pGumIHuFuGv5RaHIK17QO39NvgjqVzBhQSTj5YzLLI/zPvaXUt2RUS3kE3+8R9xbdqag
uyDQ1Xtrp0VxYnseT7IATMJsu1DDv742/w7zciF5TegaZF9MLW5+Os7foz6Lz6SlmlRiuxuh6ECu
oWU9U5tvD6gxLqdW82UMOlZezlnKEa1Cml0B5q8tKjNdjq72s52TKpLVpL9+lm3e1/Zwv6Zm+eYE
Tw3HYS+DjWAZ1SQJs5Ihqk7KMzJc+u9+GECBCCqRBlGi3jf+4nwGtnu/DTWYg2dqY3d2xfTpOdvf
b9PN+cOquYi0BT2cfVfNy5SSCe1D20+Aysz2tYUqXtZ/R+8+BhgtfU9mGvpvkJTsxFlQMD3raMWm
fbMx+wkeMOY5PskbnQKu1ZnkXBQaDb0nuafm+3acOhAmyPToZXux+vNB9PvKJlWxsehfX9x9bSGl
aZzslnLRlMK2CJkZQcVx3GySvXe0IritqjOIhv26TOatEUzHmtGiqbcv0B+00e+JwssA/MlHL2eM
la+8x+Nx6geBY2JCSyu6COmiqr4nxv06RMD0JzSJVaycM2n5rJsV850YKD6OfmBF5a8Ie08v0REy
9jEDWeFsdKETrrls404MYRYNuPzLZKD2KcFZmGh7n/TKM46Pf+94b5ay77Us+TjD6HoiqF61OWX2
/7k2bw9viRDBns95znOghMZZgyFKemY/H3bgcS2FCOHV2a3k8YQO4OmOefn3BtkllwFCGNsv2xBV
OKFFmynzOMVyWl5eNxLsHGlY+Ex67i8iVZgskumUuldhvYGH5yduFDy2CjKzuDjb38pXma29e+ka
a2ocq1wha5M9WLYm+ji7elx13PXhKy314Ys2rvIYsXCf7IJR9juAMAkN+qtIvJqkNMTSaT+CBdAW
sw9+obp8MdoyHQbra7A0H1g8tZpZtlpTa9Rnzfx7sL+EaJ/l0NW4GOG5Fi6n3968uIqtl/XXkUNv
gxGBdgkRzHS1Icz1MvRb6fCwykn8x3LQANIoqXAaXZBe5iU7mRFjT58BXChLvSUupLRZY7DKJTrO
Y+txcdNN29Z9RTnziVCFs9u4MEROp0o4EGav8QSd0KM15zd+HWpodPvOTW+qLguopdqu/ccsH+IR
YXdtdH0lEO2N3UcTvE7B5jIMjmVuUHx1dRfUU2zwvdAz75Mpo1feXn/oOSkz0xA1p9C54WOlNpze
h/7vlUgCtAl0slslf2g9+6mSkXR00pq8PFKDHtvFs5YWswf8nXsUGVg7vDGM0sY+rNsOUZqGoO4+
7D3toWGfSDkH0B/RWIWii3SHQCL+Ba88AMKK2VEZD2vNudCnQdl2v1kH6Oshe7FoHA/eMJLhztDe
epbk6r1CeES5STPtAt2mOGHxBH2MISUnq/tGIL5WRqMZiMhPOUL2MhVjAQ2hr6rElMHOJGwRfs0b
01EwQComnLSjK16v4yuFpySnYlKMKFSRR9IJqoYV192ixD2G/bX+Umumcawgl9BPmWXFwIjvaMzE
GVmspPQ6VTJcowvt3kKhUcDUEbjEYf0mebshk7zQX3FJxA4C3T2PtAqc8bHEeW5V5aiEhIS/jUmH
uCgan0s6MmLGd1V0zdvdJULF7j6/1qR5K/RHEtjXqb09aGgCuWcq9oDa5K17snRag8Tf/1Pyc4Rf
YAhi0/5mVHIppeREWjEdaQ9hDNW2+93+60qkUpRUqdNKhlcfWmpyzYLnsuU861xH+ugayaFkYQ4g
BhMMtNwKakIgZJywApZCjKkFyhesueE+49V6ovfKlZnFSj9uAKnU5c1QceTkfPmy2Drg4Kr0f1LR
5TlpWXneArnx1HvymQHro5Wxl3+DMq9mgSGlMq8EwFFksuZB3RYJSLp6kWkRLFxRk6d+sI1X5PMi
7XwGhpf7DnfHnBKAKl/Sn15nS51bNDQdf+BfxI7xdxD+eshTcqL6J3rINf4VWKo/7oI6rJDOFFxH
WUw8vfH+KdjMdB1KDlizbLDf+HrU8kbIZRzTAQHPxY1DV7nGY0iujWoe/sNp+layeCQrdDHYXPnR
ck3VAxTUJNE7p9N5L7XN6Npm3OSrbuzh5qBDxXEt5OJjCqTQHHvZtjSZ9228tqa5FwU4tJtIRcx8
XKvmxTvaG+z3IcalyBOaY+x8lYmrduhR6Nl5T6K/mg9JViLwcUaNj6JFJCN4WgWRb8wvb96OCvKF
RyujO25J1R2jnJPhGTimLAWFAUjhyQhtARwwmXc64WQnA70angBMdvIJqFGYyptYzOBq2++EY07X
DNgVIo8MLzQVI8DQ13bxX5YsvUmSpylfqMzkW5tTbqPnLFlfIGgRgIGGAmDj/TcRRLbMXxwy2fjo
hIr/ePtJ24UBck7oXltSjulbRnKuQf2VKybRsUH2NUbRUPXksBqaVYUAFhrgVLkEp2P8pBlMU2kA
g/xTGF2e3bZVSA93zpJTx9S/K0HJuk1+ERRI5qOrnB/JeF79DQkhEWU1F4siuafWGIGR/D0MQRuw
gQqTi6rxRpysc7802z9FufYlbKyXpuYgHE0NEIAYQTPPFAD1L++8Tn059jeJzfuOIFLKAbRNH3Jo
HfYrwT9YoToLcXEH63+NC2oWL/lzm933lIrw7N+fp0c1uHAN8LZ5ktpvwyypSaSre6kZ5ocE/u3I
edSeFbIIgPVGF5Buhr+YgJd5NcPA3w8FHYl7qdvDTk5Xsdj2gItTUphG9oZTew7EdeK4BQRiuwJD
gcLwwbki7b69H3RBQcXTuzDtcDxI3O7WpTyVLtloYL6fdvEPKZL3EGf2sgY2mXnnyJCKZaTM3T7m
NVda4tSE+yMWMlvzqTzrKEzEWvxMqCu3g5qJHYJocIjhKWBo6pPZbhk+y+qHghmobfMXrYfwdrAZ
SnyU6YUZ1hpU6deCK8uNgtXEb2RIREbtHti2AGjNUveX5qEZmnmHe40wfRQzHptxaaDtqxRXwmLo
0X+0GV2zxf6xOwHRoefiqQX1BjXkIVxpT++WnBtpQUn8V169kH3FTvQ8tobC6WTQPjR8S+jbjLUN
Px3fWS+TiUlIN4oaEdlx+fud47wgzyBQMzlZrOcjS+qVy3EEsrEElNRYhAsY2Gk5MkJoA8XYCkh8
SFAIkFPi/H9q8jJ+Q5X0el3nBnNeUDpGZSIp5pFiRG24/8XUoWpdCUslJXIzTOb5qVI9r4kKynri
pstsu6llnaJvSBSMShJNEfusUrM188HDIZy+Xr5Kq09kK0kt5u3+7d/L0tG/ar3VhhKFUO58Ec6I
9w0amq7gTvvZpCfon5C6TpBrBqxQvkHlBFlRXGNJc32iD9FWCQFHkALXzrLpj9XO/GOOEvnXm+eX
lLXlZfYwwA8WSozlryTrXf8IRHyr4U+JMkt2WmTgT+c3Uy5KIw9M3EtdcJks7hf9Vc9g9AAWCJE9
jq7/LwFDlLXXnuttZU6leiuQ/uZQRup/8XYaqcvdf13N9Uvq0nmv27Q1VWuSU/afGeGavrWS7OIJ
mj3nky1wbHaDyTWqoN4uWDmzmI8KiO/KUSQklZzupUavUzTvrbHzNduSWI0ks0Mqy1yWNA1Qj7kT
CAjeeH5VcpwFXPTiemi2LMo2QTzPvyZV011DQa5S/mE4yJzubUYcb+RP4DtvHeAJkkCYL2bC7qXS
8nzvaBogSuQZwxqRzMROpDkAj7FrMWF3dtf3XhdK9/lNBYM5mio0d+6wB6Nyc6MABwYgcIAu4E17
49EZuEz6C5TZ6mDnJhlxnMlNHhsjRlyBx2OQuNxKBeOPclQAveVk3Jin8ThVtM/go2IbPrlYBfEk
zQRKsSetw18gLBlAj8T2h/GX0xTvIQqlj32DLBoQEavo6tbaMHkXV46CWtuzPVeEFd+Cya1t7IFg
OQm5Lgw25l+PGWtbSQipMuiQoE7sEavb0Z5scAATl/mG22QnPSD8qfrMkQFAjdh6eVdqcDWnwGdd
CV8Z+Mkh0k1WzWET7FhmB82QRDIDWAVPEOf/36GuQCPlj6XKOTgiJ/GxFlqs9DCrIGcPEQ4asSC1
2cbVAno54F89xoxJSVRMmJpfidQSJbuq7Dq6DgAwRfN5mHEt8CUyVDWsOmYupXHBiGxq8Rrdr36e
NqXoRIur7bXGZKlSqP4rmru2MwKWfNGNevi1M+5rK6yoczKIRYvEDdMWrrd5vLRgvyFBgJcGJf+R
SW2AENBGOY+U0jooAOjjCMB3weDWpDwuWFvb6PVSXLrdkEFF9dXwSBBYFhdpovLx8fyh8VWKuIyG
AeHqLZFr3Deku6RpfwUvafymoungmy/ekAU4Bp3Tqvp0Hp9/52nqT0MS2TPUi2HOqw1NFa9wT3iW
ui38THoEp6CZCrBxEauDn6h+Xq8PCITlyvxNeTwpQXR0TjWklw79F8Ww3tPV3wKzkfUtok+2DaFw
3X+GFQpiphjoGbc3qUz6HU+/l+UAhGDz+qzJrT/YnOue8jkbHKvWvv4izze5jDq8aFA1BLwGjPFO
hjrYHlGuYsra6uAFvgzhwuT7ublfKHZw5yvP93jJZPM4lD55iBWwQa0oh7IB0Sw8sqxKv5geGErO
saSWbvNy1bSKiNnAGHyHb0y5rJdWu/8kJWHDUy17OyFXmFMaUtqhkTW7pmXdDi4TlsL+DCec6KVW
kuDrji5B2BENBga3kjc0j7j6pNbe7Wt9PivHd8hhn28Vkwdmdyv9oEm8jfhtm4TsQXAH/WWsZ2ss
aGhrUv5CJm70mS23gGeDlRPi6YADaj9tOYoNVz0S7tYhssc/eixAFcQ9h9DVcRbmU3PLrURqLLY+
zL1WJuZkyGg2m39Sij4olYq/Z4AfA4XEGFRMtptp2feRO4EC+YnozAT3hE1iLuBBDRcYVAZBKyem
cCUXMwLTZMVtT0rjQA+4q2R1tK5egDz480gXRmWQn4bhwNqCKtT0PBEU7vP1+BfYe7eB/zFOEFNy
hNMH+stpxwPhBDOJKK5HzcGjE3c7X+pC5H2oBpZV5vi9xs59QQ4ZQ/q5FGUugFS2+X4HyXLWC5KD
f8hY1RqzC1RuXkSe+jjp8OJrXhJiPKWkk89bG/Bx7ApSv7x3srHwbELGTqsdLEEgFb3/r7d3p404
2AGWiNj9Go4CRwMjRDjFQ7HEoWWHZZ70Ou3fOyKJId4AQhhdENW0mokNYpLPVpzx44r0RX7P1HD3
46imkCeHOsg23t6cUKaL24ba0adIhaBuDWW8MyCdYwNVDowSaA1pGVjm2rHi05hzyJxJJIGNtKaB
Tl5/ni2A/4fzM16KNyiGuQV56VP5RXUHwl8619bPC7fVWZ1oRWuMfWPBAs6dj3lNto5g/VnuA8SB
xouvAfLxs+rN+kbLbbCvsPC2Ls1K0a6Sut+bYO0xakbrH/a1hJ6KQ2WZ6ZBqNUZjLxJfD8a7Y1oi
Tts9rc4ZofkxHRTwPBQ3L31cOIm8Y1Q46siKpm4XJILaDz/gvnNTSl4v7S6VSHM9NoMe7Yd9RdT/
YWb3cjf7v3T4VOEMVXKm83zS/9ifhUXozZkOz63pbVd+wfsJarX9/VHQOo2w2q1O3IpUkBqVdISj
Qu/lEtYW0eHk7AJctMKGFcoUUtl2AiKD06bvpRyFWEVeEhTpAuf22R/equQEr8vzaD5/bOPvpNis
a5Krw8XUSb1EOmc2sRvTCTennyHP7WSyhCMLyH3ikBMINH9lnbUIZpYUkswamNb7Knt02yFZQcVJ
L4MhVMEfMKdwSo4QvpZowDXVWSSuN8ODBLdnA/B4/m3HBAl901ZGyyYCc9pHSWrG/bzh3VchXfCS
pBaoDmgZG0pvL9/pheC5xjsp2lnWFaJl2iiXKk/81Gh4aYxAnDdfY5V8BS6HYmZpuNq3THt7kJWs
bvpcW7dhslO+YV2rMG4Fd/CeKH7r7q/yWAEBikdgD6DaVrP2Gk7QFcNJHILWq1DXGusfyc/mEoYD
Gp3te7Vb73XNmTI+RztLDqz1zREDew8R8fmnmue3Owm9clIOrrYoUIeNJfJSi4xRT0LOWkVul2AB
hGu6W1jVkNJdh/tDH2u56ogyd4LGEfwXahj6ZBpPK7WYofh+p8zUWo/ZStd8p/t0H28yj/4v/qGA
lpC4A569H0jSBJa32M0kVPUc6P4s0O2oXFgvf105WSMY4+2BSdBncBHJ9Cb0+bTjN+gni4/2qzn8
/SXjUwBWImrgQlxF67bSeLWKnHE82PrYtUgyqTLK+cTy6FR7ko6f+r8PKPr1k5rvFAUgp/0cdkZ4
NIoLEZgerCyyD6ccfnTU1ndmlaadppAmUzGfQ/FVt0ms/aQdwaIxTxr23PWgqZZSLE1uiScCvxAx
gSEkAiLixFZb0w/hD0jZZ+nHAoV+2x8PZfvH1Zuhc1TJjkV2EcItTKj28PP8W3FTSeO5nTc2CfUV
hoP2JsvjGKXMSErQegwVIRYYhJqoHgpclbCkg1WTyKQfOnf7P21FeCPxEj52Ft+R1MgDlV4ViKoN
TI/JgeSruPTB7bbJL7OV0o0vQ5ykMTDsJdSS0pfQV8fFeeUEktmvFC5M1Zna33+hXD8vernOpAG0
3X9APCufjivuPTjSYnIt2ln6A3ea1fRkzTQC6MlCW8MhYHuIrPHzJwVLTpgxvqS8EkDYy5x02gWs
JV720iKvcCeexvNu09MP9Ccmk+w9M/umLpgHLIrNwCgaStQI9AaOv9ZmZiJEOPAfG2CdY63v7Hww
w4HBKR0X/QE1r4oVtc4qeFwiTwrxBynQXQYSNgNdLRhZM/Ze4PG5zpIRyguaHyDMiok/3NaYN6MX
B2Y/qkgeS/gnn+2rXtMcVLLoaFLNJoZCWXfmdkBKU9wxL+/uzxOI1Urwji4IjC1V+mgFJ2bCFnS2
Eo2DvxSwR6/W/NgMxqUKddk6M/4ThoXXkj4rvTgutFlCtMUOK8KGOH6f48AzpQZvaHnN63MI+JJI
63MYoPOHf/pkGf90O5NMXniLLbbRrokSnQtNSTNV00Lpq05wJXaBqbddvhiSYsOYZ/awjSx9hN5d
jNboEQRx41dRHDdJ58b/ceC6FmC6OeiCcbD5cB90+TAxrthEsSQ5h3CHD1AjaTKb0FQb/W7vcJtS
Q3QOXa6OFUlORcQ6EpYEZOaoFWuDby5JjZ2qD7K/itT1mikgKx1q32EyjzodfNjurzrJAYWjUuPK
FWnxDoD7sLqsN2p+1lEU+z6Q0p9186rC/NCHBAqF+N5wCBp/DYm9kd0oiXXK9NfmtWD5um3SpUbm
JpOtj6hBdxQbQ+hhMkDK9p/FZepY2A8sU5r4Io34kEgThmjPQRdiysCss0oFvtd4VH047PJ8hsFh
RHeV1VayAWYWPHtb4L0Nf/IuBc40l5OlYKnw9CmYS9Nb2esXtLUsmqT8wFc6fkea/yfMbsYH2D+3
FEuoKLO3bmQp4XO0gXTs61c8HKZIpdRoqglmrTy5QePxUO3tbxVcDxI64gNQmMD19gms7GYw05bs
44xrHf5G9uDin1x84gA1HeMeo03opiaWyrn1qro4pYLk2cbUDzAK9SWgSaOeEPJVzAQDTTVr6q18
Wmlu+ssWq67/x1h0wMqF0tb3yzPAGekvowMJxluKy1NpHQtHla8f/mFDturT1qyGwus/FkeK1NuK
7crTNmKRnXzIFEqZMsCTnv33nNYfPrRm45RktBJNuN58uwnYyU2memKME+jQhRLRB1psYe1C19vL
q5XFv8IRqgasVhr7kri9At/n8b4+1mFdi22ctp1imMZ3X5xHuZJm05bvivZ2PVeS0ueNZ7XjDcSF
EgWE7s8k9esq3QwWU/B3KedHEtfBg13gort2J64rtXXgedetUFpLZyPTDtXkJiGBSFoX/BkC57yI
TJWwjVpUYSmatr1VQkxHE2VChWKASaeSvForVv3tUXZ1sSpt9k+cN0hN0EoXA5yaFCmrxvYyjTY8
FWrLv7Bbof3KXu6T+3MjY9wELBlyyR2sTyhD4izScL8SlgISJoguzjlziSlq2w6Qr5IOusMwIV98
O6UZFjFFKByXXJ56dPXdhIP8H0c0t10xRzUOhDO+WULs4sh4++vMgixo2Fhz1C27NPP/gxIuJsED
/3NIfPmYqzDgZi5NZR+GDcB2zpTundh1vqZ7qH/If3HiPVSiP4KCdaIUv7tkvQptCU4ZSNg2lSMm
KypkUE0RvkFANNr0OwQqhGWYbmYVI8cr/i2dQ0HfKsTHeDlnyeHrL6MV4CHDWQ8Vg+sMceHy98Oc
X8IAAjx/KgwMtWIz5Pj9Jg2DtKOV36rImTJ/K+4eSxN6mOo1+jjezoxqXXUCvrpSkYKSFrkWBKCn
VXMq3SXzfxaxqKir4+Z/ih0+vqpgx80ibW4WsAiltzNMJdrPHEOULmuTcGh7lw/VRcwcU4R6TYAI
F6CPFg+spsCHPZOiVDfDQdz+y8rki+UuxKRWiICZg1ULK5ujdxKjGcqgH/+Y95zZBDI4L7FO1+70
BjxZjYebNDDLMzv6NAE8t0EhmcCcFGjvnoaSx3Bu0SPpV1v7CJpRVlmPjlN8Fs6gIA/lkyw0rSAq
9Yzr4rE64Kg8uSBE4umxodBnof4WLIwsGhdia57M+nw/J3VcVfqKMNXM8YOacP9hSRIQSWAPsDRw
AbxPqquFNEnYcC5D+GxN8D6NPqvGBZGrTZR4QQ1alQGG658jACjFi4jDxHHBeVYm/iNSc9GLrC3W
vyUYT3vGu06LNCxOPY/3Oz71Djj/wM0NrOsUkdp9fe3ma6arikg+wYi/gZRVC5aS7w5A729iC5+I
Z/EWGl10dAtSTYluvHJfkc8uUq9Gmgi/PCJVO8X4xDIAeKI3EMfxULrqhEY3aGCJy0ObEjWm4if+
M1HSCZMGR8nY/jgqys6tOT/FPcTTpsDBTAs/luwB1SwPAAysj28YXCzB4tDMoJbqERJb18bqC/cn
5OfRO8d1xP+GicV3g1F5xXnPJ18/eavi2bAUgoPBhbHCRiG1Xs3CSAR+2wJEMxhO7Il0giZSYMo9
pAolK4lft5DwywyKPTfCkc57PfPRkDATUzqbWviGuWsrCuM5Fk7DHrhNk6+KooQMvGOP/jrDasgW
Lxcj7x+mNVlsIM0mqeEmz4NW2iYS7uMoTevKpUHPZhC4NP7A6ypdRHlWYx5+9Pmnocu+NCfhxSKu
9BGJYUpV1JUWjCmBCfgapYfy2I8ziC1YqqxUg+RvFU+JvmBuhec6cumdKLDEl/Cc4eJglsecUmJy
sdN97rrxETDD6/md93BUOnhE4TuxyJujjMBx3cncegYfR50QH1QqXUFFi2IiOKGtd7BwHw9d5fJD
+fa/VumuouCLSTAh9L/12EPbuat31pocKfe8IWL1kGH0hdUhxPEBnM6EZvkrGbG05br1t+K45ZoV
W2wIKNidq3EGs8oBPMyy2IWU/xkLvBWD4VVgzAeyYX6T+kT0nwLWGxxJ0IsQ+BURZv53sIHx+4q1
B9YP7RZaV3H5dZdcN61COqiDkxDbjQOvOCGB7nSICH8iGviJztygqrGj/9rZNuKwCMqo+uMzUbQt
CLMQBlGNQNvLa34d0HqEmFKEsSwuaP6sjga64cpdM4dLYAWBhfS8hub9nHkQyX3nIa5/rXxDqTd9
gsvYhQz9PaPbN6TU11HvSlUdkCTTpD9l2YQHY3rtKFdzqfQ+rEl7W3rqxRAd44Z5KyqgLJN/gvGJ
pzGr2Cn+7VaVEOW0KvhmR5+ojJb0Rb2kkB3KRzhfP6+gQfuqLScYzExbeJdmrfwqAGO1BisqtvcZ
EekRE0PRWfY3S3gltVcBGLl+6A3mu63tj+buGGksRBkx8H9CdTRAmWsnYkuAPN3pUzz0+sAalG5P
U9X1TvNUko5CcR5Q8D6RDMQ2LyenW1iEAA8XNgYQxEH+lw1cm1B8lXCL0g9RJwcvN8FU1t2r3Irp
h/6sHsmJoJccFLgPFoGp2HhdIeHSwpygWSkGtQI3TioAOr4aKMiqubCsfAWZQaoRC5mMkKoVpvAm
YT//4zXDHTUYJIS9OuQLXpRWzXJUVwJ+CAqXC+Tl9gh/cK+AbdjX0RmVEAviqyGSfYnBtJv0y/zT
VEBpOTKfxBZR9Q9WQrfb+hghUzJ13DlGP5lc0NAaVwlCTN/w6hNleWPgMJKAuFhK645wNwG8G0GY
GjojWvxDbJKSDZ6FwuqCc9Uer5Gb//RqZdOt/3FeLqvZXGb9lD64uaPKo8WUOzPeMVDv17jZHjUP
dIhJfgyV/imc+WqK2MZxlO2l9Tb5U8PThhVGV0yQQHJdcnwZplnQW6Js3GswQVwahSV3k3ZWurh5
AkYgZwHEPqdR6ZLf+q5NNfbCCGRrVSgtNdI4OW/4QNxF3CNGlSRjZHCEzSNYSvwIXKCijgMCw3Om
PoxJ5BPMFEvWna8MitQAzfeJpXXgnV/aMOYJ5daM07ORm0DZ3rrUAyhpC393EX9t01pMUx/PmBpz
UjxdXkMxhimQ9UZeTN7hiHsv6uvryW8uspRIBKkMVcm07GBp+aUyZO4Yyg79yYPhhnFywZC42JWK
EASreQf0jvUJI+jjrzwYd+YPBGIVucZ7HKatMMebdHv5e/E8cRQ5fP3vjiUJWOJ0K6rO9nY2Xxdx
Zo3QDA7WGI465Lc2Hc0JwjGf5vmxJd19MC0Ln2YGGU/wmAMPTDPy2IDh29FJQSsDRUcXCx1qwQY/
AnG7wkWEPD1eraH6bf88o1YIW9oLQL9cfpGkuqhp2dwXR8RI2mTNdXzUqhkr3GJND7Kwruytc5JO
Sx/AghdQUw2der2fgDhOFPHgrrvbaH7Cea/FG7q8DKQGXoPMU742NxgcrTbwuUCREOh0MKnFatv1
BEy1MG3vMXMadcU0C49509N0kvwIcSSTmvmWeyY6tfPskpWdgOQpXuvs+dybLYyOY86f4ynD/uTE
GsRKSCHEWKCa/q5a2fPtXSL8B4ubNLfeXmkjBfi67PN8/Gc0zb7X3VDF6cRK7AyW+D35Wm3MPrA0
FAmZPrSD9kML2poW/C0KaatQ9NWSffrSW6F8H5K1ky8kqTwjsuf+k+I8WiPJZiX37dWwvxhfOc1w
uy1vgIZdrTcPrip2ooJasfgmucwTBsJc7IFqSZEBpLg0Vri8/Q6iqWUpDb63KU8ooR9taea5K0pn
A0PpzKP5IfzQ3lSO/iCeXpuyWFRvTho8BIVgQ4RkN/cQ5pv2GCEjVpyrgQxlB+0IhA7MRSfBpBG/
yn4JaXeXuBBEG0WvBotojJeYofmVeby2AVF9jzOJ+eEbsi6dyud8yatcJ6C22fQF3jEjl8TTpyLk
BUstGQ3JpX+qKc1xZuJYRCOZIni+p7v3W8nEf8acYVPjoxyLzcMvfTas+QgAeIIAAEJiiDd2U8br
VKS7QvXRo/jNljCb4t50X8x4WLdAZ+qgnOUgB7WPSSelr65OQBlYe5R7jeaz8VbKPU3Yo94nFPbD
fiwtliGEcCMFElYLBcSMLIhhThealdu/SaJwcxDj6czeBjP2+yAiA/VupvHYw85NAajqAvlBwVaw
89kaUO8d6cxpQioGS0Qj40ZtkQvv0uwQRAUcwaFRsinIGeG5v6DZkkjw7YT3i4VOEKsz++HWYdTq
CLGUPldrsbrwmenFvRI3N+I0TxKovq70HpnsyfFVPAcTdwwfPgpiG1ZdMaRDGvRSwfLoh5/6zBq+
repUMcvDrAwEbt/RO2iE8Bh01HjUQsO3yzS7b+2cBZS0h8PqpWG4hfFa2irMMY0KeXdTo8GJAoRd
Hg7kfPrxrVQnDDez7qtVsNzBEEA/zryuREZQBz65CRFnd3Wi50SAUakT6ni9nEF1Irggp9xBLsyH
NtGl2V7WtkJ5eYNJmXcOc4jvY73cnIGPTLxQnVvSp0o2+jTH0/FqktIRMyE1uGLGAU2tg3rRYb2Z
gI77Lsa4AwyJ27Mt2pVXChttgzh9GXwEEfbCOHQzi8NoTP3GM3+Kb2Xq5Gt8eKThcEZOWod50IaF
wUrpdW6RDNT/pMV2ChdIk1YKkRZ+PeUXTKO7fFLSEE9syhzboSvZSrA/lEi18ZkktKW9ki763Q4l
4QH4X2E/jyuz7KdocFTifZC3BJez8A2sida4C4v43fRFl1qEQbCy24Gg2fRbwTa9ga7PbKw5H54U
n2JTP/5hZGy8wEoJPcnJUS8rvh92JR2Yf+rHa7MTU/RXK7wc+6RJ/qGfL/FuLSLU/SpPaS7YGGN6
xO1MpxyTSNRusI2kfTZ35TGYVVi59bZnXR+v7F2fTl/rXxF9v0c0rCb056Iaxd9EMnX+vhtdjvTj
6QAFX7NZn70IW9cAO2R5/NtuqTIgY3+tzLISL4gdnEzyVe9P8EpeOVH159jQ/vEibpeA/7/VfD1Z
8NJI7APiIikUKlHnOyP0bUGp8sB5BmckNgjfPVjbntD14FLZOQshE9wbE0Kn2NdbP60kNPECU19k
D/Gfe1tkmEBOTuLUAkAHav9gnTdGKcZGWe2i0Ghr54hTjmf4gzExhWeCrjY2uRuUfpJ9vCBdQIG+
QH3MJwW0cbtJOcygW/U2i06y61pENYQFQ1wLWPLqIIHQQ1oo5776FO3B29BQKw+cxAfUzK5nBQC8
8+aIbF5tnWprYHTh1xUUohGdqVu6AOVl5dxKAwGfzSaDl0kU28nzVIYdWaABKcTNVkyW1skynQdh
OtclqtVJeJo2iXRWxvXl5w1SD5Vjtqsy53AWM6izJl1LQvj7CkY8fJYR1+eWIWFiRoYLMyzjXiSk
P/Fo5hj8G2LwmAt5ELtiolGkCX1uuiLA1ecfRhaOGt5D6e6PRIxoQb0+BNIUEcNeNa8v9mlydxOG
8+SxNO533JCLgJyThw4W9HQa5yFFfDsXHSeb196gTL9OZhzm4tU5rClgdMAI3Zuxn/QV8LhfSBgY
IB/xj54+yPgW3ZtdMjgiVjAb4vAiifqjU8e7iFNqiA0+ZbEUB1pmDNAGAxiHFA8djtYjqoGbJEYW
FZQDwIvt824m3ywcwqf2zvsq4otz3ZuxUENb1OS9aXeNySFXJujIcBCIsHI+zGmJaLWlILyzgRXE
V1HRhOGHqj7pLEKWu6WC8klJ+cwjLODr1d9rmMBIGa0JhzYfvQ5j18p3XUaOHpFBRQSoMmCozvQQ
I5lu3bnOZFUKW/Q+B7Rmq3A9yo225h3WJ4Ji9kpO+ywEf0fTrAQMdKpH5kNy2w+9F16Qd0OOfJbv
sMluGOUayLp32+1aXNBXPNnQ2DxMQjlJmxr0aJ2PvxBYpNgDI08B6eZhKk1lQaFYiLF5UfAPIgbH
E5fcVVFu2WONXjU54pCPDV8F/88ml2ZS4J8+8bINvvIAXB4uefUrVf36KrQtymiMN/+irMpGpaF1
xCa0wuP/KXLdC+Jzg/G3M3R1dAhlo8GXab2Z/QmlElJVGTb6+dKQtD2oUCSP3YqsJCd5rX+uVBcq
4kk4q2kW9ECbbtmgecOGiKvbqb5rz/YD9GxX1hH03L/MKKIA1JU3eYNdZZ1esv69ob8tq+iG/xrb
iFom8T9aLUJo7KkdzHiXpcy958A67EtOH9DkYiIx4KpjGi9GJmh2IKPR8klNk06G+nnIC4fcfr63
rySU9desU17R4zKDzcnD8MB341ccgpue0xQfXx0C4iFor8+M2me+xUZEopq9BgZjYHpM4Jkdr3eX
JG7GG2EkNxx26uQyCdJJHJbUGJyY80oZpI9tLUhRiiwlBypC3IQghclMeh8QL7l0G73DT31454L7
Q2bl9s7U0Ekuhln3/XKszVdaADBJZUSOiE4uoJcN33vEXSffmaMd3r67ANkliih7gWaf4VQzCr3K
zZ4O3CBJZClnctZYljDVrPEHnZ6ckbXhEuT4dc6g0byg7CDtKNwf+GFqb1K/ulIM32LJ9ja5bGnq
jqz59WA3mjxtIrgnrYBb9agZrAPzqyCz5sTEEUgoSPeVJxytRIiqYiZWDzdWM0dKuE0paff2JomY
9SuH2ZfBe9rA5tms/Xmr75B0QUK+T37giPOG76CyDMx/Mfw6yHyxrdjXaxtrYXdsjJdkTb/kddDb
d7RHZvmPYXZKxf5uID2MjxNXUoMVwCoaI5klYm+CubxIBYVzfTzQyk9Ix+HVc+VqatJVO9oWgtzU
gKiWBUqdHEgOP71JB+RyHyjpBKxvJ2KJFKWhbNn2B15XjZTtfGNYOLZepikSggMNZwVtp+E4H4LP
HYmTdbPlYQWC7f4I/yvx/XgQ+7d283lwpfBTPM/YAMKa2pd+9TWr6JBiP6S16WLD6jn1qpabOhFc
RJ6QolrMy9CZwP6OpIaaV6wjmlToBcFG5c6imCN3syaslnpzwQoy58oTajvsM905xDCEEdPGePXg
CkabZjiF/j6Dw71fwUFjOls4phPdK5NTWEuxbaPifY9wR80z6OGxUdAQp96foH7OKvO5jAmiepxN
y48s6+pOIasRw8tXHPpIe3jQ3sSp5CFeIWw54aigc0iOmOi7A/vEWR17AJ7vUhOSDJWo4HsY0UVk
31BV4aLnvSSTdA7sk23NSCcecwYN3L1rweRD3HuRN5fy4IMkn/vsjCG+aYE2+SwQiuZdn1PKhnio
YrAe6qqqgnhZbB2pc9SbEsPQGFnBDSX5JvDlJ/Fxvy3B39AxrCkxg3PNlkS2Z9CuJcyTh15w4/aG
mRJ3eseasl82O67PPgVSsQuD9zA7aehMxEIRcHNe9HPW0TPwHR7vScQuqPyGvhCKo65xQNVluUvc
4X5s9J3T9L7+imiT6Ds/VyCQjWrctIHJJqHi5c2CYMd+l0uAhKybhFJZePH774DMKoLTXfCo3fjf
Yi7ROPud4y78RORSUSU8EBwSNklqQqrLiNDMI+hzUny/QyGEJN8ssfHMBJaISYP92foa19TXLwWt
OrNzEcivXfRJtuwLq2y3hzHpJjauQLdzkaS0y4AGgUq4Z1RGktNb77Zj2CVILk11/BDwB+gEiq0z
2Q92u5PXtyQ/jFKC9ioy1RxCqqQD4TXfp+4nhq3C++zPYbphJe+Y360IycidKQ1hnP7RkPUCOaNo
35JNdI3ip49JP+CQNnmkhMLMCCSD8S0mO6xQ4pps1bZjmwP3ug5FXjMO3rbBpEqb/LbWEd2VYjG8
AUAElOnKEe/M+QLeGw5BJu/via/5BonGPw05oq6+eX21fgVZMWLBK5tT/G4BEG0NSw8Har+n2aFT
brBrsN4SNYxMTZgn1XPx4w5t/WzOYtLHpHq78JpEpXdFMj2hUKV+0u8bygCs+e5h8ZgrYz90OgxM
zTdJ0T1tSPwy0GWG5u3rhLFNykQeNPxh4DK5hps3LmXLEYBZg0OhJ9XkZq192OJpGmGMu7Osvsk3
zvbtKybsEtdPKzPFl2/N+eF2bcuzPWtUad1jGh2Ngzecv9Ot5gdm80fGbW6UISkrwV9tCBr+9lM2
DCFo2gRnLMndxWocD0lp9K1pd37ZjLGqII43iu0sUsBYT9qI+P7m7JF2/T2L+XfdL+qZ9l+aKU/B
m0McC4Pla9tq+2MYLDCY4DiQPYZK+koLFpOya90c2XxbMs+pQjcUoCuDOpuYQ0ccPh/56Gxpzytx
/TmXFGNKNtrAZvKLnywtO5mFcjJlrsfXudcw2K0ck1Wwgo+9u/MbFzKdvBIODyA+Y6iWxrj2pLiS
ADN0jdFdwuSaDDPijjJj6ZoGw0oUbXqfQBnzSDhl5cpQKoaLcjy0m6jMFaxzw20qU1kWa2K4KaHQ
GU3w4mNyM1HRq0vlTOIXckl3cS4KlCjwokdtJ6wDaq8xA32rnVrBThRzw658gOkNrV3Cdussvqkn
6jjhgun4eKWT3C5r9RlgFI6drL37k4++GFP0dm4TqDYn/V82Fg+klxvvgFvoFYmu6A/CzqaLP48W
dCWRXJ76yvz8kHpGaO9AaoqJ21xyHvYuH3/O5+Z6qGw27nAfz2hb17OCoNx/HStOJWAY/SqY4lnJ
FFvN9JYdFVSqpTxeyraipL0+87Tqmi9M0BrbFBfWv6U/BvRspIaOtMSy/pXZpVWgMXsIQ4QGKD0x
skYl3tmAA+FhtxAuc9yW3ekyB/mF79aVtt5x069LU3HQHCD6dU9xzxXcLlLZU+QYWI+6Lltr1wUv
KsWAOMm213GvUnWdMfkG2E/tPI+Ih0EqGeTvneStUqq0/sWgrqRC/2SnRi8gEEVoP0tzuSG6su73
XGQJ4chCYS9rPiN5AN3DfFzooUseD3Y9H/8aZA3r50H2Xp8JNKy+xkEkud+qCgCV4ABsyyKKr6/C
nANaVKB4abZQW8NAIBVS1Vb42+Ktle0aFGwwSznZoPhm6wN69MrOYIsJh+1NXjK6l0VQ939yZ4Ec
MnPmMfQL8O43XGNQNUH8j95PmZFDyAv1KnPWx0X7h6hnejrhFBttU7MadHC8SmZKHSKMU/FOaqnq
nyBNPBmnFMRYE3Yr6skSpzOPlwm/fx3vS3lHVyi9leHEQ6RibGbFijk8fJyybM7z4Lg8eWJkomJ2
jGkRXSdOpqbHnFBVR99xm6r1BL1VqNpmnQWo5tSCwOtUgupcvjWsEMsp/Qv3kSi6Z4PEqFzaRVN1
CPrTvx3aBo96RIB4jrb9ARCJJQE5IFHAYR76Oisb0dE1hNTXEqDSaNeJlfPIvqb35VOKkYEIhzhM
dJS9ynwRCWl/jPhY3CHq9YJ3gFc3YLNK1g5Ji5hxy0iuRVAQgR3HNvXJkON4prDw1kQ1vuqDzLUV
1nSxseFpqMGE4V9atOhACWcH2i2O04axpNygzs75EplxRcfu6WznTzgrGnI709wKOQJzUuS00l18
nzVzMnxn3m+cfII3ckT9V9FxTzW2iZiF+jcQNeGrWF5PGo0+r2NKuoWIoHeJ7wDuvKCfC4pyC9dM
epYdKa7pSOtR6njb3cdYkK+htqcThpsKMEu/dlEEJi8JwjMCZglew3+5HqonbTHBR/e2zYyS7D2b
hW1wX13cJtZUvGIR2Dk1EKsJxVsWiesSrwba2iqC1XDqXoVVb5EvMHc3daj4j/dWlqM1Zi1I9cJr
8MLfd8e0nUOiD8hsJU5eVLez7kgVKR0m1ZXCCtgEQrkcu4iwtglzqMJ1Ktp9IxBfyRbAmaha6rnP
VKI+BNw54OF+LL2wPG/WZrtcJOG/BNaVe5kyA3x6abPC7OLwYJtixDNBoPL8JJu6aXToqJaAb6Mb
kLHErODZ0xUeAhfSgkOTpltFg28LPtM1RDHiVEKK9kFRfXubYu8Pdtz2BsRaB/drw2rFOAj3ji0N
YMzApw+cYIwY79auPF/oROwmVsGAFbt0JvciylDPSLeZ/Ej8KW4g2oUaNGM0gsURk69IOx2gCfCy
WXeLlxeyzKGiLhJCEkiTZqOLOxx/ZExO+CFvZHjrpA8bN+Md+Fd70MHX5ct33Uqps+coGUggR1B5
QB79jdym6L1KteIj2ZuCesAoyHa7J0CO4oVBBjxMuXJeXYbm27pyneMFs1uBxjtIh/YiwfKghdK2
CdXk3JxrNEYUckAdprZsz8dEzVbkqZuGqg8rmmYgx4//+BzalHdVi2WtANuGSXWoQyWL+7l01lL+
KDYpiebWc8VNJPpjomZjBGm9JCjJN7IBA+fRFUlDpGvGxLXqEPqRZKkdieFpB/E9ZX0JzWi3Uvsc
sBjeppGfp2Ea8ZIhX98lgvYvfkYA8HErJdNPSZJ51dkvxRrYZ5t7BeAew0erEXVKa/sL77uWaV3a
yrE+SFIoO8P5L9Ca10xTg1NCzuR7SQsiyIkT8gZXlVjf/Uyf+TYc7nBbuEVvTbSCWh+FagRqwCh7
mtKUdyy7Psx1cfS1BGPOuJewdfsC/7ttLobKq7IRXIIrzV2Gr9HsjSIDoh+EJ8k0Gd/MpHJK/mlx
ySB1ZhtyILdI9he+TMhygalAzHyP9B8o44kLuzu7eL/a4lOxNgVNorO+15dD1M4LsUD004SxGsGS
xVVM4/228FOUnkD7qpzPIM9gn+alI96B96FngXu/8Im1P+yxXwoRW+kwegUIyOOgx6Q4FUbVd8tq
nuBBJjs9vs9qRpTDJZgfedfgTuOFEP8kE8mDshCd48FY8w7L/guN6Oc3Vd/VIwBaCaK4Ob6VZ6Ue
DwK9HNVyqLUlqoSSAomTusHlvCvvLPEtJdJrPHDbMzHVeVcNllEx1p3CncJfhFdSVbLn44uVgfgE
wAMlnfee//xKJLamEZrA2dPnP0m9CeMX9a1Fus4imhb6bWHI2/qqTzL/7Q1xpWM9WB/hB9QcghF+
PBxrMb4Lp4F9R+Z2lcAossTwK3jogYq5/wevjJ3NvJ7vF7RJLxH3zKJZHzMY2Yyd+LtBdzjO0XBD
FNLYn3xbjEiR2YdTtLB60dO7xIp6n4h9i7ojyDQLf7Vx50JFF2f/N1cHdK9kEgw9f7oCNt4Jffee
A9/Scq4kllcptMm8H97PkB+MhelXhpdxUVVLvrTZbWOam3LM3Cb3Vtb1WkpmkzUwR23AvMlVKu/q
3kGUyHDTZvarzvwd2pebAxvDSgc0MzgVZsBKFeizmtISavOoOIQKuPpYEZW1l3yu4M5JZxFA0AAI
cvNxA4Dhy7kJNVjraVH5AEVqkiPocy7n+9ytKlZ4sz9x82mYLJhBNsQQcBLGp36xelxn/aYGOspS
JhgzhUDxkYvWvFllaP7OURj9LqOw2oLSBy7KB2obfaTmEBxNGoGC0kP4avtQGxinuvTHauscIfwy
XMfdDuz45XCuY8FOLn2nblEw4MJs63PZ0fwsgv8/5dCGC0oCHtIvLZqwsSIcJHLjNncBoerqfqxt
HKahVlGUWyhj7MzDCDn0W9cIewk0ZrSDPy30zbRXi+ATuptUky+E5qeIIV9KLjALnQNEANhCbcoM
YlNNhazSKC3HjfxYO4sC/wlp7FaQQK4VqAL57FAlvaPUmSzsbgwit7BQ1X2zS22atZTaFQSsaqi5
mOYa2B5FFIULYkBx6cQ8FWrptm+ZqtKShhwjMcH7ZYXwkUTAVw1IDby6gTBkBiaM/LFLz05A0QqS
lcCm+RRdasPUaqD3RsL9hUUcSYUjGJh0HKg34JDvbyXHolLIYIW8XJow5dyKqm/a30sM4OYKTtZj
M4Vy1yCOO8yBxY+4UPbJOPLXSK5GAl7T01opIY0+ZbeoaPJ9IRWtgn52s3FpE12RajMppf8dv0zl
YT1LYVNITXqC0DsVh7TVIAHQsu0s3r+vAZWHK8iDJN9HY1D8j6Zr2ExjVdeBuGSJIuzmM5C0rn9l
d898vjo/RuLSH+F6aTTXwz5s3NISOnH1Y48yzqySYljWqPBaI27WZm1PYVRPPK61IPci4kdu9ocH
Zde/9qWinvMRqRu5EKNZd7j2R7zEAi3f9Y4efoZzGH2uP+CsK929W7bHEfZ9JStcZLY5FkrxkPad
ONkoFR1tAjR+0Ycq0JJV9i2L0YPhLnLs3K+v4aSAtvILDgnqU4ZGAAebzOrLk5Pv8Ny3F/NS/qAC
sp4qrL9vLyIxRYMuehnu8dg0Jd42FbRsANAMkPK1EXx1oPdMe2kQ/qNp0bxUdAob2ksuZIQHExMd
UPQxZ7zsnreuGDF4w1G15/q8aP29pIo8gFKVWR5c34TfhHwWqRAFMj6k1ZPBEfUAC3QT5J3m4FzR
pL4imijP9O/g3SlW8omkjOLOzQQqxJhkk6Afkk0nqEP4xCkqksZ25nK4x2aw2GPbEQZcFmyxCuLF
/m3Nao/iiD5VZKRY+cQiSORMrxVoTrmPyeJbOA+tf5CFc5el1/MyuKfWh96woYch3ZFE5rJTHc2D
aTd6/TG/LJko6PN4n3/XwDZAz3m9V96BpIxLjeH8P4BtzOQtQvPfnspGK/HJxpKfyLWOMaFjt1le
WAT2bMGIN6nxIXtXQjE+U4L08a0CGSiozPx5sldeq9+Y3MhPfImSFtGGIo9Bapa1QGrsfG6miG4f
6+C5RStrEdXiBwCg+FReOHjPah69Dy6e51d0MJlO0wdIUpB0ga8ZRInxnBeWNFPJ7IXEYQXOfFCM
Q0fa7UyASxvwedHzSML8dNmkm4tqEJQ3JQKylDJSdCtHtNPAuARFyyc0gG9v+uCaCkyd8unKtSdp
r56w6ylaZm0=
`pragma protect end_protected
