// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FtvPlRWM6WbgQosTVDReds1Mco5BrMOBrJcOUqH9bjKaWJ5z7HRad84hmu5pEL70
2UjYVNQl2QyCcAsdwEL7y4jMf3SYPgaLvxPuscriMHhvSJ2ZJ7KMtoSO+Lz6sw1X
tPv/t2aMUE30SIJbqMYcMaNCkK/JwoaUrvlGxW2k6LU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9904)
XV3aX93CiQAON3mD5hEPIyBIYlr+5rL0E37LZEQOnLaJe4qHmssBIBtSgLh3zRMu
+FlORcqxFS/blX0eiwrjz02H0OlBVRvMEALnpXc8KJ9jTr33TnlmB1m3J2LSZv0o
4QF9jINxXx0HyjN7xh3loQWvEs9tOuGBNlRUscvoky3sV7sVXf/lvozZR/rUPY62
+pzPKOfn6g/31ceDl/3Z0Cch7tO/ZRlnLtDRpcPRP7pEh/3mNeY3bv15SRjeqvvM
ybYLCrMK9DYgWEVoUgaBiteQkb9QbqihuOFKdA0yP7/9KyuvLBFJ+kiGrrA7bDww
soqrIhBQm4eMPlIbvgpz/4X6nsVij+ReYJfPWl1bEvuyQM8CuXSBvPQdO/vfmr/K
PhgAITgwPI+agnLIVuAIg3PvdjOCRqvF9jEVkZHMjZe9tIQUPZeZSVGCLAkg4iR9
K1BwpQqls6Rr+gLwjC66qPFQkKo7YxlS0jJoz5l0sjsVbZnxeRYDEq8t+AvW7LyU
ebUqAFZUsyqtmEOL6C9ZtWcSSjtWrkyN/2GyZyxBgqD68l3dWOXWas5bNfcG+wQF
YfKLQpWkTNvp0ukWxit47jNpdG5FdsxTsOzK1fUqx+4EaCqZPnNJ6aFwGdvdslA6
R9gqTxJX008EPgtztsquDN4wjw72E1KjcaLonKpcpuGT9znjFhvX9UKtipXP8EZ4
31OxqLUb6tkLefuDrRQ3rb1lkDpn9lm9HF93JiWTCvpbbk9LozMl39F/aXTiLM2n
bAiwBw5jSadaHyKP6CFqrOcgku+CEYmkKfp1dDKa+xs3M8Ru7DmrDCH9oY51Aich
wY1AsKNsk11eHk9L29J+8ml8G8BblYyrgmRkaKwY4WTVrgsH74X5DSfLb0jFD9ie
G70tpcUMWK/8JXOCbQValzVQ/X2Iy6Xrs3QACw+v2qmRX5PXi+llr/09ivr10OxC
PqWFyrqoj/WYB6k2PV0Xg8pMw02Ey9nIswKq5Tkwlc2skqWiYOOgpLgNFUBdfc/h
ji515CxksDtIDtx7N8QppbXaasEpi7n8opdgRSgUnl+m8NcFdKdt0tUiip6OFwV9
E7ki0YY9H5DzYqiMUSsvW+r0scXvilNeNlAuSDsynB22h5Key/ZG5kn3aueGHkyF
CE4OufmFTcvH9DQGqGrq1bhawawXdQAUqc6EfNF3IcbgQVZc7Zw3vNXi7tlrqXkq
djaib6HwlHYYSFJwdWG00EhDSgRgz+qzCypySfrslP8Tgm8IYTNyyw1Obv8bSCWD
EpAUg9bx6xRRSs/cehae5tiPW5a4Urlc7qwhLd0yP+aKPrEUVTIyuoHilljPEs8t
iq0i3NEQjn7lNnORzLNjuNVN2F1SBnI3czSwUsyLStN3gQQEgSv9oS2Ds+Xq47mJ
LlDkX69/CA7WL3JZNnEIx4AYP19FLHdx562GEIC0nGnpSAdzLGQefb9k+rHIkGiD
MLhTvn3Z6Kp5o/a+AynOgrHPX//JKGvOLNQ50SCoc5tPyUriHHgFmFqhSDHqeGmw
iTfBV7u1jBfVCQeLTQsLdp23dUXGgXDLGj1DuyzFahM9t1YRpr2Sx53EzCfxjrGh
86VyjgyTuDQ3u9K8HAAnnMl6RLtr4vSHuA93KlZF+aFkGdhCHOV6aet+OMUDzKXe
cKG0p4ffUhQgShcahkhA+QgBPbpLG5BIWyFWeOEF5maWNXQxoXzmTX7cc0vPX4Bb
uU39cE8t+FGtb4Ee3+4Nvddql45f67ydes/6FNp7WHWj278sIw8GlLB78cvtCxh0
G98VQULOFmo0zADAxkB2a2Gddx0TukFSoC2zDfTo7XAV1QYpz4DsJ0ffCa2heOFq
vX8d4XeKGqVUTC19Z3H4KH6LjTf5T5+cbMa9eDkJWGDpN2tVsbZYPqtYvpfFusYJ
GNeCewIrrTwGZe/rTsWcra0AYcXWZ41Bz/YjEilBQCZoEg5l1iQux4eo8DJP1MFB
KQC7nvXd72fLCBY51XgDMm+a7FBZkVkOLIBCnFNMpQ5O5NbY++ijMW8e4qJ2O4vJ
SyKabmvT1EmN6rzIXiMZHnYXlB+oCZcgIi9pDrZeJyUqlqRVVX3WWUAhwCw20NWl
1ki3SGVfE07ZC/9VQPg5nf2RTyl6NQOhqP0U8gaBJ38gNU3WiE6iqt1qXIH21Sye
hyf2fSfCU0kqp4RV2wiibOB0o3kDmbScpqyQEML/oodQ406KAwaH0VunakYaRyLB
XMALcT6ElNyDjgVG70R+A6LYVtqO+3A+Ju/7hHIa5S6ZwHSu8H0yC9FYgPxfNNzX
uvddMcXLybAUmfqIEhW1bPYx/FxwiMlKsyPK5Ncc/XbdmivdTiNKS+9mq9ewU8qf
QaAe6/RZcYP5+9vDRjV9JkiAoh0rwDdhme3WMo7JjqkRbBIZN3o2+sYpEy7GGXyo
s97m0WNZ71mkmjGpCjGBB2UOaR4crmsiMB5YlrbLTjhMaiGf78fb8jf2644/9Tqq
5H/6ClWuYh0NeG551l6qrh1FUuvHrF8RXkE8zl9+YVOPKzjfkV0YTZq5e60aGeVQ
xC0C5/C2vUfuSRgZiFRmEk0/6PZc/e7c7llI8yJze83v1qLOWkdAkMcbGGg3C88f
JMP64qlxd25wWcVjjtVGdHVmR/uIG4MyB/Iwslf9FcTBuRSBJpvR3I+opj7SlteP
iK2ucezcz2QzGOl0YEOopJLJX3JobwQOIidOL9vox51j99arKIjeCjU5N/WM62dy
pr63n/QCsUIpAkyvv9PSYLmrPMGSWlPoxCQ0LHiIHlEfHfqLxA6AGKX8Rn81YmO9
wlrJdoX9T9hPRODDmHSeMJcSEpFEBTHpKas6uhqRqcuIkw8l9NOJueOPzlMO27fH
pCndQYA7jHSJGtWJ0VINqsrVT8TdthjyeemsPz+U/R9TXUMBvawghiUuxOl/buwJ
6g/MFDeiN22UaHLwiY5bNhqTdiOWGpG5J0nEtYOIlhqr/FhCkl98oghr/R2GQDV3
H6+TSzIDTibK+yI/ZF0pD2YFfTErDEqODwmOYNZwePlLkm7wDouDuUk9I/pQsuK0
pALEjJi2nyTZM84XQMhwdODSi30/l1GrxmgnS0WTOsr3CpU186gE+HQE6LqCUdWw
eYd45MEZqubQp/cHhc5hP1LVa2JkKkzarTKMH0o5Ty7mzofC9aE6zb1AjH543+M+
9x2AzyqgVUYABJQGWBDr+T2psOSYXOe8eimZFcnr4fc2tW62WQRpvtQzTlt1ovJS
A9m5kubxMof84JbBMwZXEEzDIEaxGWzbsdq0LBuba3/yVpXwEfwi4OvUlbZ9d8HE
kWC4BYW/ugVB1L4mmbloMVMiJFadiOViBfGWhDd2Fun/4qSjCBhV2bbZVoGd/jU1
Q4OYXvH6glAu6my7/KigGRZG6nX0Aaj6EAcTVGIZVgqc394nsxjmKH2FIE/8sdqf
nXza3Mw6BnyO4XSRT6anBCOkjexF/5gKsYbvzfZBeCBJT6TAJGHKiE8+FT/h7Wvy
ogg7UBA6LBW0l7oePqaK8mda30alfRBDcAqeSoOh8LcQxhkxoSpyv2KBK2tTsUs1
CPyNRwRD9+8v3odvw+Ov648AzmBO98ZFnAEU2mvKHhwkKrX5Z5xmOnJUcdBKWt0K
4sjnGvmE3o17R+qzFTHXUUQe13YDxJ0bSSMuKJhPtweBTOwJjg7PJAGYw29rrpWA
CvTa5nymtJbqiiMe96FTV4Mxy8FqKqrgeCddk9R8PtIdvUhP/0f2CEg1kCsHYtoV
J40cAlpGtZ0HLbpRtCUGVchSBPOR/CsBfIwLNdB52ckgYMG44gJsx/0kK2BzDnxw
4vVznCZx2Q9e50m0IjrLoNrAxZeKPb1C0Uw5E+FBSJNG/s4i1TIGuAPdQ/nulf1/
30vSaWxbJCTNU6ZtXyV/Da73egiRMEiorjtOMpyjyspRM3DdlZuz1X/st2yekH40
1dNTLgg6FMom7w14ik58+I0psV+Cg2oZjdZqIuP3JLa/kebHw8dhEDFUR3DHkG1a
MngXnA2pHnXESYjihS8QaMxoCZ2lUEyQrJfXdvlz9wXzMXRZUvWdp60BFJIYrWvd
44r926XJxzzU5zRkvDdSy2x2kbnvAnVPm1Ik/RHr9o0tBwlaXNydQyzV+4Bm+6R1
ISQ0yFWzwQfiyb7XeG2X36Qzoy+Wf7XKkD9bcQgRdxVyYB61x09IrnGqwTjIHiSw
uEcoWktWcIhnvD4baw43MZ3l+yWVY4wz0ApAzG/9X5B094Bcgp5JIZtJLRpAuymt
j7lwsYs7Y6XV+fibRfs3qepCeRcAv/QFkOAZFSi0pN1LWK/Hsjb21jy8SbRvGg70
ZfAK713U7pJpX3j7Og9s/W+2/qBsDZgTGaDZWFxtq/NcydmHO4P1Z6QLlq9e7YI/
sAypQg9h9tNvZTMl0q8ByvCbE9kul/TcIw9fJPhyJBa14AKAGygPpj6jNyt7fkjM
lIDpprLrVE4bTBq5uguKHD3Y4tlbXFQJEh+mdstXtmWzeCjyGqHYC2166gqVLHO8
Pvz29AcVSbwHJHTj43+WdvGuQ/FpkVJw7DDxZlXAJkPrvlJu7dRF86hD4GGluO1k
oIqQbu8v9Nzx5R1HRjgZJ58eBgfI0Ujma5qNStW5O4tPbIVcUNLVWVY1z+MTXrK5
4MPSTA8aQFZ9/Neo8JyFznX14tFr5/SxoTJozzUipslGRMy3j/uorKD1NyOEK8oX
xjPN3EadL607X3HpCtcSIJJUqS/nZqgpsEQNJ2KdmhgUlSBWOYfkFg14g2sqn/S/
tJI2BB89c1t4lDw5g/6qREVRoMWlKGIFGb9mucagkPAmQrVymdUEagwOVafCGc+/
xKVB9n6VkfnKCYrm21XxPnR6ZunSMY/tydSRsP1yslwP8vptZiAmLzh/zqIImxAS
DWsBQW5xn5xTi7Pq6lZU2Qa6dRghMOtkgFAoT9fi6mwO3klKm1rAljzKEb9yKCeQ
L2GTrdUADq/SMUneQJpbkHVfTrwhONceidUaez5pWNXtaM24HLCuq6UxI+tCrVYI
9u2wF1/KIDud47Hj+imqnlXxLYKx8gVLSeBkCfl9SNXfrTPj2RzOnRVE8FLX6dOQ
4CvQy4jQFl6GfwOgP8i3xUt3lia/xzl9LdcexdC7mq5AVT16llGvIxWPLlzYR/fx
VtDa47DiwKIkfTBOazJAnbeckPFy8Spw6m+lf1PctLI++jgWcs6QF8xM9HBPpr83
0Hkk4AvXgIMUQGrOW6J/xxzn+evXGXU1CtVgDKaCpOPFtDXhKgAshxujqEh/f0c9
u9FcaM4ob3/nffKrmatG8e2qM5ezuCh44goM9B1DwbHhf/YbI5SJZ84jrqydXO0o
NDyhaa0r1CtLdyy10bpCDiNd3BkrJQcegkHqIjM/grPOsdorl0suFqFWSFo/eju1
qFlD14N3TIr8cKcB3daedZcJ44wmhSJ6Vv1+/p5+Ruolc0jgZoC16Myrt6JaQ2Yd
Oi90NntBEZ2Yfq3AcSO6r0zquQoctV/dwkdeIkyCDHn6oQ/MO7kgzSlxF7VPXAZ3
wJfxfL6IUQ401InueLSzlUeigx2tJFKmDrauyKPlwz2dpBbhC7/9qlzwZzSzG55N
YUnPOCJIobQhcIuytIOxbEzC1VEVkYITBzu0BV5viF5wMDh/mu9JpncZ90TXXTDI
7WdxFPHwP5uMfutTcisxSJ7JXZ6R64zWr9jg9f9YsCSgNk/jCupr9EjN9d4zipYK
ubQS2Gq+s+oppwLyHH2vUtk1i/4OhbNc7JmAxZs+UyR0sMJJ2Pm72TIPnI4kzqkg
iXKBorh9JA3CJz4o+U2KlJrpDWY2YvPjzPnLNz9mnAsBRWPnvypeOTbTrycvq/VN
+BcJfVR5rb9A7r/IKaDSxGc1APJKcPhP29BpxpPuJol/xxtpV07Bl2YTtToaW2SK
dN0QmqTMReBZjEX0yldXrlktR03+73/hgJA3cOvb/05g71FZ7hIvLT6B8BcOwVIy
ucs/ztjJ4NOrPoSDQhr/gDDcXSrLhrIJD3bLy+PUv+gPKDALXSXojzsPu2pbm1Up
c1YoY6F6Emhw94B/kATBimeC0FtCPHOKkcU+4SJBDoe08OWW26uVs6C9T4jlN+Aq
IAsXVCmNA+Y1a0ElFL4h5lOHnwrOms71r8OJYma8zYU2LsydjpwfdbUrGj8xnHOo
Su82nz7zBsItopWnTjYPugwm6JnU/ONfcOqzRJE4UBROKehDSqcxfz3za2wtpHuq
oXwW6xBhnzsxj204t/Da3yTV5czti6KKW98T544XnjxRH65Zn7SOeDb/sW7AYGXc
bGJxSGtwHdjYb+C19M7Lxz+NADtniSQ2kJFJvqK/ImNPVqncwrqOTzhecVNldz42
quC6LGEsidNIbAAIbC4SgbNIIkGQLS/gOfJfG1zhHU9fxlQ4Eorib3m0754sd1xi
z2T1C5EaNYDMe4Bw/jDMVYpApO6VKthAOov0em9L1XhsSqkfIGSDvynfhaN1CQ4s
xnXW2KZ44p4DuFzSBxZoCJMMnIGbLKwVwD5hYCz0csFXS20+p2jzfaipd5WgCeM0
GTtemM3ejBwfdztkqB40+M8DReFaXtyhkx+9BO+6qeZHlM0jfIKVDG7Ln0ycw3wh
sF0UvLuWK4rOsG9VxuvmLRD1M7QYYlEZ33Z0sKrxm1otDdv6BGoXiODxh0k1us2B
RMHzumFncg7/Ui5m4BsLt2dHs9ymPeeTnGoc0h0OwEljHmDzu5/B3KsnAHvFSwPV
R/EQaYGIi0xXGNpuDq4VQQr53fvwnjNraimSSexD8zvwZzoAvYlARUqqGCkm1iG6
RfNx7jOFaY2e6Zi6BRSuMv1f4u5THtJ+jJIMM+Kw/QUdAMyA3ptDi4bPGnkZrWYh
kj4mX66b3O3EnHvN6VXtqCSp/zt2n0jUToijSzsKQrmp8O9fiATOv3+JN6TNURKL
zWEtic4NEPLSY4MzQHid5ZwtTLJk64gF5ysA31VOquVnGWQWio3dL3c5cqFWtUdX
pMfuJEJ2LRsk1sdU1P0q1d+mOZTtfMlzl3mtY1ydk7iNs9S3mgeiTf14B/1VVLyb
SrbpmOXJS3Icq8SyyvF8fu0lKKaBuNYAf63JY63HmoTzCY2mKUeaesRmx5Pkexaw
P5EP/DtpjjSSJjtd2SY5rQEPtpmUNI4kiFnBWYcnwtN1ajIh6iAwPULwsAlfJGvM
dEJMc/06L5ZJRhpuD+SJa1B6/wcPWlZPa+mJ7Ad/RrvvI4MmGaJGk7uVbnD4rQcP
580Fb6d44JZhzSiyQO7uuCIuCFsMA615uydT4MzAEF55nzP1l8bb8bFZhIrMhOxg
GLRW9gNm33pp8ArLs0FgItC4hu6PpQUUXGneDRWiPts/KggQ2UO/4koTV76Q6K53
Bo7waQKJrXG1ZWEHuAlCA2FOJ9rCvhXpx01aFc8CXLRMAMcWPzr3sqrXODmrH0Gg
FaWpDid1NySODnAbd+BU3cC8XI7N/Tvy7crlAnr/+PXOiJghPMs+bfMGS/+QQEQf
gkGemoAZqeNZRYbHIpf4EWbGy+CcfedJ/71LT3HRfUFfx/xUW5syZFo/3YclByZc
5NixIfjayaMgNrjtMB+Yww2HD/ybDYzJ3R1qAdFYjv98Wn+1xeuNVEq1pGsZxa2f
Uo4vfbsD3WOq2i3FbQN7eKe059y2q86KNLZGEjqTFyNU/pJe+jtxSsemFvnbAdmV
bGnoWTI4YskZVD4KbTw2fOB/r8atubQNDzEhOvB8uNYZ7OzttWgB6JlymLr9PJDD
RRU4ANnbONg0bVKgsqpuootWuS4qdnrQX4YNIBwH+q4I9TuHypGs2keaLpYqnyPB
vPSnX+JRaw5H/aKPl8k32JW91lHpmFPMfZBgbjCsQurb8SMD/RFO12ch5OAx8FbW
AVAQJ62mVApC9VXlktvbAxKDkRdZTy5r8ABpqobDexqeMa2bW/l9+YKZ7KcmASNU
CU+y8KG3YzhPfyLZT9218h230MMWah3xhmZWfL4ZeVfDw90WkBYRb0KmBPkvxrgg
H+wqyTaY22PMo/PG8+Pp4TlLDwXxGqPTGi1pKcNPA5Ln9u2G16WyI9NW+Bwq/Pj5
pA6ML9BRVZ7al4nhDcLaI4lHb84L8Nj2VWsx4dPJg3OJ8hQwHh8hZNf7CxfA0uWQ
A52tDCFI1e/FtpDDx1fEAqAiBo79J3p4qrKXUJdwJJ7PNJkgc0LoJxWUlsEDxgSb
9Jtl0kZedot/cxO9y/UV/DfEEFhHgOgqftdIMf9ejstrpfBq0IbAQEaTbAflzmgn
5gZyKEOCWdlLqx/zm6utKHZf6G5e9EzlvLb6HCLYq/gz6LBSo5Jswm3pE5sab8+R
rL0jmdimn6LA0TNNfXDt/2XDrDJ5bNl0cKB2IVEDWKz1BTdHWXw8Fk5QBvBAKG+A
cgksk8bJCFrmBaoPBRGcY7WYdqjyyny63USFBiN7eBW7VLiL1ozy6ZxjH3v70N1A
HGHAdt15wEF2TZtxTjonjDJUsKV6jaOsWf9QE84uHntHXV3NwjZ2IHsDnlVpkeps
EQ2+naIk0bW1viHmB0cWOHzr3yDFxQ0/pk2BSckaHydGuw8Dbbd+0qBwYjQWhhJA
7ys8yRe5z/5IyY+Hynch8PmhkN3GcIxkvPO0L1M+CXMA3VcLYHxS2hV/L+Rcsfvu
4XdtdOb2792kLuSHQEWBWIYlIJXhQ1SSvho3c7wRCukvUbzJxqFecgpfeLp6GGN8
ecJIdDSNsS/ln24F1R1G8Km2tV223gPJ5DKcqagFVga1RNZJzlr23HiZ0Z0e0mOn
ZRv96/WhkQLyQZHosmdV4TIPWeA+B6JxnhxAYPzzM5f5j4doS4qRCS2o2JKd8jIs
zik4wbCz6cl+ee1QitvFXm/7e45YXd4pzA6g3X4LMjrH0ut2DJm8bBk118tCkk9y
MTHXU+yp+k+BTHAiadkShUi1rWLbutZ/QBcgPUU8D4N5aBTxdGUzayGSpt42jea6
0FcWocZs0L34PGlYX6dGsoQ4S6WMiI7dFX+zAMcpfwsgEalSOeMwJG17m8rpbyS3
K4ls+qhIaJ/qaKTpTviIDzTM7mRa8NbH64HcTJrLV+u+gCz07kfhLk2l9AWmtgIq
u7TY0HIpWvv5M777wXerwfDNwuS4Y09SJnb/SGktSx8pK7iWQgzxg9OM2CB5b/D4
69BfRjAKcRSKskrXGhWqV+sf3IMTBsYm/3T4DnfXC1GGRKtgiOwUxLEQv+eZeFyp
WSgoa2zdHWnd3UY2kWCsOW/tNj5+IE+2AYgQ3n57/2R/xBhgGVup8BI/zgPhUrGA
mUKPK0AbmuyJlVYfsw7SF44H8k4YEmcBS9WKH9gSMuR43K1xGmTaIIbnSR/PJyVv
fBJBDdtmNgtZ5JMX+Xd6ixK0c1OkqO/FZ0PAIZb0LT8XfW78qOQAIFMfydW/gc5k
XF5Cq2gP3g/7XST1Peqy7TGtpQW21XefsIdJaMwJeaaIpa4U+wqt0nUrTZxH6ONr
xS4HEYTwwsW845IAorhnClJZJzGBBOA9xmML9F4Hlh7j2ZAhmN388axakj/nyTRf
FObcxhzp7ScQh77+JHU2xzXkCrWDx8PLVgKFwTVp/ektMJxi2V0pzoEjCz3Zimk4
YcChV27Hyi/Xx0n+kBp/IwChFNAdqeWO2q8m88jMdCs3PrDN8VGn1mWYcIPKgVye
i8KXPcmF0BKJgeBUSh7Fmp+2Jc/L/UCxSEC0sToXFS6PzgvzsJZp43IneC3tIbJq
82UWQQY5MZUv1ykaSNBjzWBOmbqbhXv4sEpdQ0QyUL4ojpeE5cd9W8MopsAQtbHJ
klzYLzvGF/aBwzZmTM/2avArncy+IS6PZMqCS0QYctYq7bWhTCMTpGFbCX5Kc4JH
11mK4ZVcUR/uVWmL31oi+N4YQp96Foqvnk9Db3UFJvRVkjP3OQSe0qHRr8DKvGge
iIx0jIfF97Yv46xD40VjrJh6yWxubxs0QBnoc2bD94tYZ41F9YbkU429P1/EO9qT
z/2gJktUlZb8+k7T9Zyp+hABAAXXhwcdOFS8D6cPsC2Rr54+sXEDC0LfNP1HeD6x
RNfQssp9MUuhFw1yPhrl9ZWnzebh3HqYPpMpX0USJqKiN3SKKlfcuoHMWmvFdpMo
gX4U1d2JAzdpYCj2zdeglizy7YOr77W2N1IDn2DfQ1xagcjm9b5tmtANi8H4QhU5
BoAL7A7wAiZq7ImisXXrNeJjodbb5fFaiExWGFOnwgJdSYbzN24gf6ThiW983258
KCBF0v95pnQvI//pdzueQcY5rE+/8go7iU/fhagoZ5mZe47zPtQ3EF6kaL8tfkM5
TZ8OwoQ3H6xhv/1WbYPBN1xL1vTuSZ86FboklMFeEFUH2YMc5CiwpXpRum0/38nE
3K5CVY5QR0zemzOvbvCPtHToI7Jc0vJZbn+gV6vtwcd0KSmLiKtb8/D9SdBeDOuh
NMVj0YfKf7uoVTVdZVzvbQ0QcI/Zw1II9k7Ii/Ec/LaZm1Sz/JRL3RKtbJsKnWOU
DsnPBH2E0kJG4USYTlmopccP8fYNOtZ12J2W76A1L91nGrpm+gQVMBc6PuWUk1Xp
znn0fcmzT3yI6PBCO0VPSKej39q2EeUJJaXyCWyROOPa25h3n63xftXvb97F51ER
xMGbzByG/qfV+3BdlMg/iS0aEp/VWKg3tuYnH6W0GnZVJRXod6MQTBiB1RV2Msa1
pwv30TsX0anLxEmZMw0egQ7E9XeEOwS6KST+FxqHVGqT9cTTmUx3dAYpapNz2cow
EjaP1CI3SZskBAZE9P7B9E3NfgrzBJ+hBo0j6C59tuHaJLrEFaq3LFIMDGvBIMaH
Auhg3iq0wctsCXHOlUcBRl1JhtkdD2ABLyW1XRfoAEedvPOjG6jPQNZWOfbMeoZI
34L5aBgDVp/mdAHF915YHcKZjEKd17vV5ez2MYj0HaNP+A938eqHOhrl2ti78x4h
rScAYEPMSa5ZU0o03oj2THgGspM8u16bU2GP1W9/LTGk6KxhceNTKnN3XbTWIae4
5wRRrBj6tzVV5UUBznthxKm8wYxcTtgalvOtXREA2bkrVFA1LMyrbI0GF4RP7Bos
7kpS2/+eiJYlrYNSRYuDg/w9dQcb6qYBwa907BZHejD7Ea2omehEwTww8IHoYmLI
Hun9uv4gSYtvYvPK0B2Tz+vCpvp6ZP0UIwuDvy99ya6g6IClCaj6kZHw0PmOEy6p
vRI5RSPbAfCrKFtJ5vFi0MRE64TJihxqwyRe+W3wJ/YKGN3xpELYpjmLqzcxmtZY
zH9H9DmTW2qi0/8Ps3dApruqTpfLXmyoA2n/d0/ltu79r0cjKUWwPNBqPihQ9Xp5
ukwqJwSqURsrLRASzkWEPu8aysJ5APdFSweOxjo45JmSdOdswYU97AO9UwID1Uqm
NlmHRSxRvbjcEoCxDlZPbWjHFgpr+17vl+yF0M+7vqS05u9SUMF21IJwStkAZCY2
kp2Qf45HNutCVY6Q9T+1hD2eZcDKtC0ZTe/5cDruD3egql+5jIicOzu4c1rP4nTG
WMMfObZ1HSvOk8LS4EJu2yefbSFQvnDp61RPAQH3WwwtxJAIc/WKw38IEF1xglio
JSHyLS/wRCYGECp4TUWtSpz4X+NnAGQ6ITuepRsqLaKF9Ncy+yrLmw3pmY58C1cO
RmWKiwsA3NceSXCoAWHd7oP1SmYDoiMp71X1XA4lroC8q4um/kUUr5tTFs3K9yRu
eBJEFA9MNkHpOd5MjGcdNWEuSP07atDMLqQXTEmUs3NWNz77A9q10YNYOaZAeAjk
+Y5E40eZKl5bQU0BTpTWop8uMxfriNk6AJZduMozulqs9E18VpVledR3xhkmE+Ng
RL6W1CrOrq7bvumPotv10bFdAPbhNkia+cs/AuNvsFWNNl5ekq7f7hNPFfMWgAkN
9RmUlViJ7qd5hla3SLJ4HLe9OGkjkibLZ1aZ4JXaFJOAF89DhANioC/Wl0DFvlLB
HqnDmXEj9FnQw3sb7X2rQzlzivltXh5z1g6vyqH9CV1op4Hj4j8YxaofGOQPAV5G
n5GaST+0fmRWq82LdcaCztrp0bMpgexRiFCa5fczM+fR5V44StwBNu57jA/Kdctk
oP24PPhNQPLurBSyY8KwdFVSZCljn9Igdn1d8R/MHWqFC16nXFUUUtM/AVKLWTxT
YYVrmBS3dp/kc8cjGYioapRhC46146pBR7yWAqzo+SB27Y1aRPDnD80PNS7QXImV
AUmjVqO/M3HY31nMSPYWFP8qq5k5sctgB8BSUswmodBVJOKgkUmcPSXn8gNe11QC
Yo/Q+xP8UHoTsjY3QQtL/vkaWL6hIhtBD7bxvdcqgDf3OtYRIrpmshud+8dK21FQ
Kyrr0ohLirHJBSfPtbxgEaJYxLJN+OfrrCBH3p0xqZxRvixjgJsQPF1iY4lRv78+
ivjpUVAYx5cCBwxrfDgpVg/sHhNkwfPJ49BPVrygKna76KZtdiDedJb6OjeojS/f
5etjGMTdqBPLotlif6GAUdSRlaoRc0dbLeD+6PHBWNaQG+p1yXMecOKHug9mHMo8
o10b8ybT95FtNLsamjfagW/e6vzBOoHKga32q0tRA75cNvWCi5AKMuEmUyOdH/Ge
KUtuAFOqR7AaqAvst+7yyGJq70qtcue9YC9NOD1TZ1clCbGtBh0chxPGXwX5P/RL
OkYAskxpQbgSeWE6zBDxpAu0uRHEidvmV6nQarx5M4Y7JqHW55j/tDwqypAnUKl8
hWGEZ3wehrOgrOH0M84JVik6wDJMDCD1l5gem6NEw6ldHf0SwoK50bF9+zQn6vyK
8/USHHV5ORyN98hvcmNdmvBlRs7Ori8USeCHZOzb1rcWw8RZ48K2xGzrBhE2I8pX
lKRIgu7aqo6ufxfSIJn0bQIh/yJb12UUOFB/sPE5PYnESm1mhATeMVcpZm2GYxEw
tMC3JKJ/QuiDXs+wC2i/YP899z47wfb5HbNtEda5/Q/TY/fvY43ipGgD2NiQLSqx
NgW2TyB/UAAjoTJ824G7fpfxsETvaZNe5CWv2kAPrvmHWVIgr4n+195BhTvET2BI
a8XMmyRI3iDQQlAiPgcwojlZp0zVmvitUCV5uwrEnBWuQ7zf2CYqNzvAmMkHIylr
bKaB7mglpz/SCEkzkMIyfw==
`pragma protect end_protected
