// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pBUu42LqtMeqeAM2pfiai142tTLC+B1qIvPak39XNZPOUsl5Tail12CFMNhywr5v
1qSnclN8Q+CkjOXchLi4wVeOq5DtyNK7Qs8UcrI48lJWC2Yfi07bHm5KpsrE3kTs
cestgJMXrw/TX9bVRa6481EmgG6z6jsVWvLjmo4i9us=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
EBLTRsh/W+ni/R0fHqyXCWFgs/e4coOcd4VqAfU5X6tEyhajtNN1ODMLeb4CtQSl
NDL0D4HPyKoDTXIBMjQyzgdhJkfcr3q7hpHrth2VGcdgqp+/aw+233ZwQgH6XRKA
SJWePg0FnNB3g4E6CSLCC5f62QSPcD3RWIB85h/2ksT1UyOARQbhKAtUjws3e/X9
ySGnUbq9ZTU3XzUJtujs0I9zbZ3Vj+0yL0oViGwh0D+bdmCqtcjg9TikESjThvJ7
FczgWoV1jEuCkWYNyDAsk5trRjEuH1DdTobMQZGPmQa/+aH5CzrL/4n14Xzl8nIC
9SJsY6QdBsQWbq7dfxWHxvl2AmdMK6VKB8Fx9x+rT10NM9TNF1ckoB+bZ9q8pGUO
2vxOqh2svoUp5W6Mpq4FEZ3K5y4F6oF3Rszm7GLoHUMamQvs/2ztSkUJmT3GalTK
SoPc1FThuk0J1U/FECfyzLu94XH1jStYahi6i8evgR940lQfHutYufmCHvotZOhL
ZHVYwgNOh3CncZk+PUAxBKMIO49WTzd3BDi7a78gK2HB3WnxxaoqSJN1YL2Zx2qs
SSwHmgFvypzH5shALUIFJg6kreZRoF+EULDKBK2mTdN/cRJyHiWwZw/5n3aDoVPu
sbmtdB8+LKXasuwrnqjdI2qnCWut04/MF6oWQmvkEzt+352VvZnUoWvSih+a5itm
UdRp88Wf/qVmevLKzCxktAuQ62vHomkuJNdjVX144bm7/50rIPYp31OUxTZBuVmB
dyv6jJM0mBCaXH2NfQf32arN9uUJIS29Alqdrsx2GcnxN8HRsXrI91OKD64kqGsg
5oxmHiAmKKHW2moDo/Q7iZdZ3b7HigOoDuk9iNksxeJ3X0yhpZH8ZeCHFsA+458+
pUtsbjUW5VOBAczOD+M7BSa06mVqp5M89EWP+kFqNHCgYdzxIxi17ALFMWUiyS9B
7mgSU4wqv0U8dqSIkUhaT/1ju4AIJYbmeJ3IfeJnAIDINWKLAkpDIWBjdehl2C0U
wz9lJ9XZIL7qs5siOCh8AKjGFzkUiWTwODcb8JD8xv2NLtrabu7nbbnfeSH65xjX
L1op9cBEL0OMSNudLkM92gVojyPQZ+22/mo+vNpQUMk9ITgh4tqAKYt6kLP+tTQj
U/POO2s2Lwz32bcD3BKxV/3kyX6Z9/y9lYfx5c//E6HNmLtV8YzkrG0btgCYgmPO
/eueatxqngwPW2gj4zflGUneFdz6DsAPIV8ian1UKKX86+1tPMEXr6p3ymPp5aZB
qzLIDzThP1uXalDjd8tMCEWQEuko/WfYwsyas/sOzWMbzOTVU98yXYbRdffA7RpU
FRKztJ4z6ehVB9AETkJv3nHflwhzrJb/zliG8gOm21Qzc8hQb5dJT8B1DYJIk7pH
k6b+6vcZ9vzjQEx0OTImfO4SOr3i8we+DnVf5sTpy367vjc62mcXA0LYDuVFfAiT
I6iSoL8l5vvmI6xLHgconIeknjS22hHI1Fk0XlzPXS2m7Ah0+vX46W97vn1jRtnL
ElfbBr7bjjB//LUgpEz3CS+USfLuuT3eUnWexiJ0Kiwzn9QeWlg7unc/WWbpEETe
oEJw0tvEC7/pNFlrkVallhgERUCioR3sV9FxuEuxk2E9EBWoCPWCKwLGgRZ9HE7j
4u8//mlxw9nogn3rYG5S9qK81M4WLDi88ydBKGSASmf9KXp7WgHnfRz+BcawEvmW
nwmzYZrGq6RokFjh0n2dIVIfmI7fz2hHLoQllYAirVb7r+zCRxVn3g2HoySPZJmm
wfB20w98yg6PaC1UQC/gzLEnJBzAJbWDU6qpCjY1gaoRYvlmj5aJc/HlkvSYz0lv
P1Dl+rIMHjG97zW97pSNcNKR97D8Xs7SPaPs+UbMVF4Rg5wvNXBZbnhedi0jgxnd
6/1Wol1ZibL+Wmq+5PS6gwlZ4dhuNqwSYe02REevTUZz1moPIR5wDZervnn8IytR
upoLZ+gj33paDA40UuG0yaPbfT0Llw8nc1G1v3Q/yPWbYSydg1dXL+jwehXgz5UW
q9o6hfT2HQl+74SSKzBZXemzxpBeAth7PqDDTccjFN7XdRZiF5NtDUly6yvLzlP3
08oADX3sAmhiTvFETiEbiZ1+zgUVVu/qac75jjhvjf5E5FN771OFbQg71xY4ptGv
F4pX4GEU1Lr7IrfH+v5yQ/JJmygwPJ67HX2ZavRks50GtsOW+3SOzqAWobwLtkd3
Tz/vDBA8EQG68dbGsh2Mjw4HFPJh65XWdt6gdp9akouzER3JEUfcm7yzMkoO+vdv
kV9iUDr8hgt80D3snuCtIfnkzMLBdzp5wZ9xOYA2Yfja+rG9ylXzawsEjBIHUlBq
KFWlJmyKdHwSuzcPGpR6aU98MDtqjAKt+akss5rMl0KIB2mfLIpfWfX0FGvD3EE9
OaD/bOFAj8La+dj0fffSfkq/BFQe3NZxicDTWd7iMI6btVjENplfTZxuFmcxb/qA
BxJ7ttmWyNIpYLViiqPUs8aQ56cq0mHBuRm3E5MnrncdnFQps+jHGLJJJyX6V5nf
8axczE1BgoaN725jZb+FmY0hhntpKWIcIWOIJhMYdQHaIYGVgcREtCllSkNphhvv
qwUt4Amm2xmSLbYWf72WGiN52kVC8Ak47lWUv0Zqi0dnrx/3zcHPBdaZhezXwv25
y7kmPOiSdk440bTQcltkJ6AxVI8je+5rJT2SRaJflXZpp0KkMAwsJSwa98Cryo8M
IIgYP93DzvC9kIFjCI1JdFlzPOn5iXoZx4VJglM6m/NZNN1ZkWu+JfcOFlK7Qr3k
5fu1nhP2RilxLWP0JP/JBtu+L83WzJpBDB4ULshXPu92Zo3P8W0Kjk/3x1Z+Rz8y
n7BwFp4IsF64ujD6uiyTtJ39hdx0+yHFCXd1Lkd9Qm7LrKqhzWaH8zbDY+qqFuQ7
6o9mpmBECRVvinROycPqKXALEYEYx+gdbMhZHPCTNBwUDStj929OrmMT9pr1vW4R
D/Pcna31+oGY0DUiYeti5qgZo4EiC2/J1B5And38u/gXD5skk8i/mZeICpVse/H5
ujyL65MutYdao+Xe8r4xdxSDOnQxYOeWW4ZOxEMr5OR9frcTspPQTpUb4ANZT5ok
qNDfopCctzQhl5IfK/T8FBDRsmP9CGLSMICa23CbrMrx04lfpMpwCaYlMNnIsfc6
G19uoGiTGyhW1r/k+QHxQOcv4k4/AoxTAcXqTFdHS26bNiE4ox8icr+VYRLZ/8ci
RrLFAp1GrkGFONUPfaBHa4ja46JuPcmEwLu+2vYdixpr19ByhIDb19lzKNnLvI/g
ly5WcU83fSxBYLU9jy0e19bnIm94BeXZibAcJt+fq7YvxawYREPafug36C//um3l
mg2lGqapiqWeSgOvDZdqX3qpBe4z9Sno3oR9bSEWSjOsJLgduVTCJOPD8u8XriNL
iCVh+uq37AgpMvoHnDZ3d/1fgDPFTAG6bnKE53yPkQqBGVnniQDUqdjREMVRCm6K
kz5jZOAitXdLFaqQPiQjqyy3zugaa6rEmjy50zvyhy/UjS1nND7BSIoDzuFebiC2
aIAOmKWILdOAGbG6nC+hgWwlhRTxWATf/ElWvNoOMSYHcmfXH20XQBonCXDrgMvS
XTc6guWjPuTeQ9i2Z2334XRM9wPJfB/ay/Y91auwgJO7fnIYZUEHTUeDf7J4CaDY
5umLqVNPcUKB/6m3iEKg/VxP68ns7U0JFPUpXCclyARg9sxBF7uXcagXBS3P8wiI
GxWwxJz0oZnh1zrq5LA/TwdA5rDZQ3MpNgberZRGu/qmJt8kZugr4agercR8/ROi
p+jPLDYIW5aq+xyHYUaj+AnF1u/oWfTMaTpaBDyKcdIw/4nPyf4IxhZJ+pj/RsHD
tAHURMTqU4UxQft9JJ2+kfQwC72RfhRnYQkrpYfDtKtG+wGOALv/BoGRilxYJUoa
uJntcJoCVz1KTprnAZIKPoUStX4iGna1kJX0Zg2Q9jHRnUhn91NoE96pZTAlZkt5
PhGT0Xtg4nX5AWxXS8nbuFRXUuguhHdLvyJQDR+IoGGb4aR5y689eYunwOj6sFEG
8pieDv39s3aUMejuPefViIyaH8jAZ/Z+7awf7+OiCzhYjb5rLXIQBjcxWDeUShUf
UEbx73OGK+QarJ9b3x7DXxAAA8B6yz4c/geIIPOR1rVQwWGNQ1N4fvhgyqtS8HMi
jt66u5OslaYQhLKxox5RpSnVxa4dDPdel8aGiAxQ8JhYSl1++LI3CsnokC7sd+Wz
h0XKQzchg9uX9Yk5j37MpNLwdb4b2cpS7MAC1xTFYCDuMZYby+2rVgW2T5J0KvAK
b/hQsUb2AUiZwdkqDMYGvcXfadgfDeYeSKDppYGeoBgaYyCi5nMo/6jrrIdOhGCd
qEdJUZ1JbF9xSlxzVR4gbjgePel8QeAm8sMsUNFqpignXDTVY6HpRb9m/MNpubNR
WV2XiI2hd3iK2z+dP3gpW1BTYDCINwJAZkRjmX3fEbQp1UEZDt/2QrlZQG5Md37u
7ukZhKQ2EDlLOlea1jTdIONuOrByJdfzUVKImUTuLW3HOvLpSIfJoSLoqYEHvs1o
jxoDWx+IQeHS7MRNsmSg9ZCtes5yQlVOEXvdNRLOF78zsRADPdSetJJGgIDPdmxd
e1n2WEEA/9F0wikd7tTB6y9xvEr7sWHyEzbK3o8j6kkhJiN9H12/YO85twO7wLXK
aWLlGgH9G4aKzsNLkBAmz4soen4tDO7d/KCEmsPh9RNPbY7ir8KnMRraJHlCR9M3
acl0WT866nPAPanxB/EV3N/TBsGL/5WZ0wUsQMt5NaNO+AFe8kNtSF5S3EyANN1i
ib4J1G0KVC9t8UppK+SYhV+geFGwyycmwHkxFyrgNkkmNM0QmoTSk8gG8Kdmajoo
dE+pktsi1noKgs7IBQrkbTxwf0GSAaw/hp6P8NEjkQfK/kjN3vYEX9elh3ZixpTk
q/y/K+KfiGLxZbdm15I8fHPxXNEruhVa61NQu15jEs+Ppi/aFJtrC277YY42SYOR
SZJKlsx0MN/navjMG6Kl6o6P41KPFlCb4NJeCUcdsRa3KP55Ya/lClo30j3wPr+0
Vp1sU0lkHcn4rlIboSVG/F4RJhSctzmEvh+hmto880jmlFuNN6Jzbhu7d+TRK7xJ
0eUHozGn1/PLP0ACE5T5owp6j3NOWYyEuFuN14HNBWc3aubN69cNLwUxGJtrPrOP
PKmSSkWVH1qGRiWu41iLDAGL9KpDo7lG+vieCfhzoj2wqGhxD3ZRRyr8+iMALF9l
Hv/fAWe8gvWZufQRpuLzyibAQ4WcSH9Bm1VouyJwYVeiPWA6fGRCvRqPgXDYP+WA
WFYOG3i21j6BI/p8vRXjuPwZWe1FVXOfmD6cSFUl/movEX/YAEWEHASMWnwIvQcp
YjiDPXd5q/MdgRPCsrtg6crt2iGd4qtP3BCn894hxALYH3dVS0a5UX+pswll9+Q3
+wLoxM1BQoK3cvol1xyBn9CiucPIF2dYUhxxu+xfBISbbHpINymfgqaHBqtJmER7
Xvf3SmNdazBE4gWr2SWalzIRomj8dhNujMBxzlmVHTz5hQ+1inZKlI9MsyqNhACY
2Oea5JFPDietEyaB76Q5Yv/GiTEgO/tZ67kCdeo2TkV3nP56lfPGz5QMwfA3k6g7
L0bh0vbWPkpogNQl7224+gCs5LNpKgC3MiWmpw7kR0SpxjOoqIgXNzNUoHRi6qv1
RCSOLu81/qLLHlZR/jrAtM/hmEzje02bA5J81lOBansxS3a5xDvLBlWWwxMAmg+h
S+Bbxnp3KzzKNlUvsKbBsjn+jDb48Y303uhFDxSdV12OQJL2akDeb3DW9c0GM32N
NhNTOkOOEZd9nxGiJrqyNS5adYERsq2829wOiKrMgjvZRI7xFOaiDFmTPzHFyGJO
ek/TOC0pBJtVnu7nINCAZ0r4nPj4lBCHQ+7Bvcx4rOHfQ+EG2NdRGQDhORhUZb5S
dhYjzei0u8u9c1ORxcFkYCp7FjcX3If7MFAKVbuY9MZMrJXWAX2XFHlcdxd+/8ZN
H7eBz3/DfEYiYPexnpBO+JkmnfgUavuHyo9bM5U2dG3+XnQUJXN2n4+vxTlLiCZq
QIJzPYfaPMGU+iareL71H/YLirsoa0Sh5980MBpV3ceafZovRrTfUElhOU1EUkUb
+yFxTBboQRqa1M3TU5B8cjDeabKpMg7voAohQdl3YWNI1UhqlEgKdDY3GMoEZQEe
ChR+ZQ+kBNP4np4tUZQGlTwDDNZe3t8nBffbLAakcrbgPRGvGLRdQI2JYV/tyhZJ
3/Xnb1fHugnqJu2QwS1FmXu3CebRZz5JHHG27iF6S3KXjvj9MUpqKeXnaHvHi7+N
zCym0+GYNPTdUKhTfIyqyl9yPSnYV0EBNPUobT15IIE92UOzbENDgSkTzM4GUQi2
9IocBbREhtF5H3LDTwfb9gX5r0Oo5gCjpyVlfnAR9q9fHxwnNCEF/+9XTqw3vhP7
NyfcKqTy9fd9M9H9cZnSifLlZ5s7rnsdlzPXTjks8ACP+lMeSlwFv78CQrb9fvh/
D6AmDrwj3Zk42offsg3J4KPkY02iy80Hfh8du2otoO/0NMemXoa0QpZzKpDk+TrO
18tHRotgHqpH/TVJ6UcBKWuzkmVaeC0q3pUppUh4bJyGFWJHAlEo+C1O/7b7iWsP
56qHblh0cmJ9JElC1wMXqTOCK4bcI/8TbBx/SC5/K8Gq1u+lszPHfZOzPe1MsjCq
ypFqAHj3qtsLfdNmy7d8jzIRpxH/P1U3rljUldnUfDBom4HRD5jwnyq/g1G8Jbpg
N/tJjIcK6amV/SWk3k5MIIO4dPoH9i8B1xBez1hvymnE/eDoTs/MhQ+Q47NB1YTb
BEOvWp24j3QfqcAcR+y0pm+vWiGNs3/4Ks4Q3RAFULQcCzQZkcSwju/od5eKd+bo
8Gl2+SYJV7N+WrQoXgXGjCMas2IUQmep4F4yJHA5HkCEfvGESlKscTTF9MKoPG46
xCbzvQU1KtBSylO0o0LR24HCydOHFvaCr1N01QLnEKheDRDQi6YBOJbSG8/ADl5x
Omm6YRci0QKluXgTffLyueWPydZegAR+2q5yV9t/4/R4hF6SwhiTksqii5h/JySl
Qpy4Mu7vI4WU9OJ+jGKiOTd6ZikxA3h9Dl4S4RGCnJF+COm7d5UbFwv5Rd+ENEOd
aCRTScX6UgUbjItgCjiyOMGyGYesYelxdwTdVocd4nkQGSMPsD6oexXYMmCnhwRB
X/r8VKxeiXM4C8jsEE2tZJOGLoagkb8w9mzb+McSe2UPSO6znLc4aq/a0/+uO3GX
Vg1td7xsyk5lZU9uGuFBLA1xPE3QQYkpi5ZJznTLp6ZKthQhRtO2Kh8fD01ar1/0
IvocOsoGPChmAPAesqtjpEYoKCi38yqG0Gl7AVoy1DL7/tvz3atKUZ/pZR1Nfr/n
ZCSVAcjhfNc1N/c+CT74BVPVuA7ljSdOc4LKcM1tB8xXPJ4F49cnpg6x1ZC4bzL3
GOgXvU3n3BSz1zxXPQWSe1E/ri0JdCmviKpLQjvG2GEDz6rnTVWDzfg5MJcVCDMc
`pragma protect end_protected
