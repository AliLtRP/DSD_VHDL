// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KtMiUsf5CJevg6KU7uOidAOn+oeLgXTgrPRRwNZBjWKRK0APK6jR2t2WLnbVQwp4
9D6kOoMTFzgkVEy8OtjwLkeaAkA//LHH3mGHa6q89/lZdfU5YD16E3/x461UohEd
MzcsT/RZLQnwWBZh+ybDSunpjyDgyezrSRTp55TOw7U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
2B/Nmv6k8Vw2ExxrcSFpuIma0Og1eGlI25tytbJ40ptHeZfH89EzfJNCZvaBef1A
xeHu/w2nbd59q+P1QytU3CqvvNrtWQAjpfJ18/t8VTdfY8yZ5zuCh3e1xEsld48G
rn0O97hcweliqQMpNwZeJS5NE/pjpl9UsfdXwX86zq+Xh/r+DBAucdmnO9iAj0FM
pS/ObSuMBYzFngskUirw48bWPB6J9hUgOkAm8iswqSnDGVL7JfddiddocbHRBZIc
qYAsRfp3a0JRVcaxFW9+JDqVZjQMUR2mGd/J3ffVGc14yCUu2dtWRLXKIcZF/X5X
1I6mP5AShQa4TQZYvkQFaelZQXbdwXJ8LF04w1MXPDZQaH/J4aEu8V3xJZz8BcLE
1FL/7WVY+Mn3K6ClSZOnamcoxqeMOhnP/492IuEcZCKO3itiP6zDp+3qAbw8gwZT
dwlZny9KBkqL9SYm3V6151DC/6QFe/esIIKHP8NA7clczksMEFbREXWfFt+suEwg
BsoZYwoztspVEcwecrgIk31cfZveIPsRUuOtWC2Ec9f0cXfaKwllAVk3OvHmqo0R
JFV+FDGa2iBJIqI5i38u6PPckTYSKaOJ4UvB3E4m4XSPF0VkEcztZo69BCiAMo0b
kNaA1kQmgnDn3Ae2mSjGGoQ1mdLgQMjIK3qH9kiepCU6njEPWV7TSBHoQO/a5tPK
wtz5rQdv6Tyvi5ZSM1VS5iIExv2DB6jH+7+MijVNFRBFXQ8z+s0UqG599yjVEZ20
O47RoOVUzIThG+nD3ZtKiXmRN5dl5kVH/hlP1L6BDmqJn4B9Q6wQG/UOcBlAlJ7g
g8XMmnu5sEK/JRXbzMnxh0o79tZ8onOvxbRZb8lHgnaI6sXlK83RdfOgNlXQB7Sj
pMzgaojL1N//4PoXk/3N2oo5S1Ft1y+FcvY6PdX6XTvpn6gNmb4g4JFQb5BrEEdD
Tx+MVFDQBfaF2+554npz+1hEzVrPfZQMk+gFbpg0KNarg9HqI72EAE9Z/BgTU7fb
DfRtZ0DIv/aNwZegDNoUmDmA+AmIu/BRWiQnOPRZ5J1OsHLl+LP+Kp5WLYikfUOZ
pCCe/EEAt/IbSMN+6EX37XLrj7Am3+PO84eGXUmvM/Exq2B8ESKspssfMUBp3sZL
zJTkNBnwEikJ8zaiCSmK1tvmpd9LKYc8Rj/9qOTdLVd5YlCuPlBeLiBoZV6gOVLH
/hF0HiT6I4XGkZnnq1emSn0utIvyclSe/B+gVB2zxjZ6QnAt2LMNLxUrYX+KPIF+
ppVuQOTDQWeansZKK+ISlDDeCOYzf3NS4YNVp72wYtnf4yppj97tuh3j7NRCQUcY
rKi+A9+Neif7EKok8gLQZH4QwSkd/B+WDXRcuhYqSWigzI+zXEkNBq/7CnEnDP8x
XJ3y6evK0dmJvEICqh2Nmi3okSZeDZbyPi//ZNnvDCBGUXX1Q5m8QlEQprTIsR2n
XyOQQZAunC4vc5Acrby4tJfo8YpCtPkMb2ykPap5V6ZHTyZkDL9jyiV/Y7tSf6Yo
7gr3KOHYbKdaEI7LbGUzLpIUo740pl3TMVSVQJGRZRBRAyApZBdSrBPymyagON/k
RTgM9fbXl4KUUZFw5iogsy/Yra/gU1TujOqBRKvNI/VOCgLcPspAh/L2ML/LrkOK
kJu//vY94fAx9vyBBGorzqXksOxDoM7o44tEK8WhtIXsmcTzj1opf4QESpglSnyy
41I+Xbylqt9Wv8M5HRzl3SK7CkAET98OaCnXQZqiLB9eaRAg/PepzsYZwbySynzg
kDPwV7SQ/GG618FgViMHdjEuhk9iL/TY7kwfBrTPZRfPHZrm5qmEmpewiv6ijAkz
wD2LcY5uetGZN01qYZB+BVDAsINDbyJiVG6gqIlW+xBcdNL4B0ste29yApp0sHnO
Uvq14Pw4IQcHEy3OyzaU775PrzFrMlXAEfj9nuAiH3XkYFs5wPE+L+dFeuAFEc9o
F7LUSV0zBe/y7rjIz4+Cvv+tW0u2RRvFcdasW1Mg0HMWzkscUKukSxIJBkS3ZOzs
0CF5g6XJh1lQZjdrf2I3ikItA132JZpaR+/SiJbwifs+z6Khk1ldyj4OdalNRYxj
B7b/X8C4EpozQjQaPSmfEy68sAR4VYsCptPbsK0IhrJLSf0DOBAC/0zN2Uek8blR
j+yGm+uUFbNTNfVKJGQh0KpAnE1GmXm/z0CboyUKsvYXCXC82aMqdLLwgMjBcQH2
PeCauF5Po+Dspce7LBEY0TC83nuOJ/KXKdU0UP+7dWd7Ru61KJVN4qTapj1HMfYH
nZ4u6/DVd3I6u9xPal00ko7OW2yKgcl3+2o5drT5RAc1d/Uk5tjWFbq9lfYQFMpQ
FlWOrRzZilu8ugF7x5jD9KI2j9qqdOO+DI5ExNBz8M/BDbl5dbAt6tGt9pwgeVsJ
+T9cJdkqtICNrNo+KbE2luhDbUnn6xJi6+LX4tpWcBXKmUaqATqa12BOahG92v3b
h1QtVKm6u5MZffo/uyTV3j6xBTODLYUBh0JXjCnfENPt0Em1lcrq0U4Rn80W6shY
0mlhHKoFW36l6V0REEJY+6j4duvjIXQvOBP3jZcYsRio+dPSFJI2sY6UUDU3liM7
vTm46sXyxDTlA/W0AqZjvc4rXvBSd4/L/cX5Ztfyvotm642l2vzywm0Ah0gOEc6W
68PM5J9JPOPyqPFIq7HJXZ3HZNedDwS3Ha0n4tt95JSKVzkpyXgxm6nlxXscLnXd
l+ur/I4hP9GgJhBzSjeg+svXBU244HvbHe77aewCkbKqesTXnLrVAjrp4Rkc79rV
Rh+PcVblXjYSDMIqTBP6AgyonMaTTE2+j6/zj0o38dudOp2AeTi6YyUQvptORVQp
t+isNFlujAP8bAOK7Q4SXrCcM9buFXbMrUOZXk9iLEAgNg+1OAuJlH4iq049ilDt
q+VB0E5pdQczHeBQCVhPkaZKtJIhavzZGC3WbqeLMhATiiiqNqfW2MCc3n3X6wzt
W3IC4saVsppmmfYYLz/5GG/d7oCO5sPfDQK5k49Gpz1yYINnnKR8z4grzk1LYz++
6BtwCjMhPyCnfoJDxiJU8IRmJU6oTz40mjFrR0dnkhMWCm1PHI4EVEyAPzO577jG
4vEloDAh0JniTTjXpmi7lUOXXm9KI5ARsKyaO6koM1L9woHEFNAr0Qkr5zmx2Wer
JI6c7F9btXtKrO87GimF1Jy2CnLArWkkaiSjjPdQPShhELh7iYSDSH2T53/Wh+fj
aaseSkbm1dknlanCb7UUEy0N1SV14l2kd9tgxMQ6cHBa9VULrWVYNKfUmVJNpTyn
vbpO2vmZe561kHc+TwUlhfOaNXlh5fn0uXzVdYJ7AFToXPpAFfsc7KdlrSPj4/DV
yq+id03QmSQNvp1sSdt3Ycns42UyUwgJ6MUQoEvMsR36gIPCfcQGmVdkLVhvQ7do
gQBT95ALKy3bls9X24Q0WRQW8GXgPh4fE9XG742zIaCwOBXfqs13ZKHGMrHjkm3J
jj38xlY/rD43R4mBE2FDsj+pi2mI47WFyN6mWrmdYxU/h/AubslcBrY6JMbhWioF
yLr1VMo/Z4m8cKDp/a8Tqaj7VMuaVIIT7H2tedR0sHQ0AlBdEz16IqqfDGFcDXsv
soRDhm2XLzoirgJA3lTgCeZ3xqyGsDkScRpTB/K0/ajiWldrT2W5oSCh8Pkhp2N5
fWkygAKAiLP7DCjRj8+cDWDkdIrCuKNxP60CczXSJWD3z/edha/rXgSFNuj5q8BJ
Obx/+luZAiNSqlvaVarNHbE+3KoPCtN5ZLdwUET33Va92ANI8kdXVSQwXIlUFnP9
spbUm18GhQi/+Ccv6jWdGPH5IeX/i3f2Zo19+bi7Zo9TcjWP2+eI/tW+OJAo2U5c
xDJjjX+1ZFQ4TArgtb5H79OfXpOi4ElZBvjaelSoEt5//UmeCgUTAKhCBQpHxGNJ
cyoT0XALmquHK0+1Kwv2rUSTD0QQOOYEcC9xEIywaMe1Xtrdczk+oh5GvGk0TgWN
aDfE1HLCO84QGyn2iVu0j1hvbWKhKZf6igQ1SbQDdD/icputIZn5wPogMJmaT9RH
x2htS3Kikpiauwkvdwy/hc1SK2vt8RwaOTdMRUTe0J07ap9QdwjnrHa4JiegcHSU
AM3JNCBP8uyw+t4qrVum/JLWs+Dm3VCQ2M5S7CCiDFbnVkxbyHKPVizBjjJzOukM
KyyS4ocStgzpaw7RQcGMEzvXZrH26jyd5Ji7K1jeWrDn96DMN2g1BIHOovwp7wln
CFYOB6uVR2ibn4nCiAJ+W5QM4FDUl0u2tVFdwp7gNXOJcAEdsnarfvVovHuRIB6t
aqDhsYe2PLVVtn2JwTAQef+WOWJ8Q8QJpRpwlM3d8Fml6FDMws8Ll7SL/mFu84AS
M5y9lVuLc4sg3PwEfxEkexIA7POPhIKXyoWsrGRMVGhQ21O7spFfYiRLn9xAyJCO
kCz1Zr/AzQNMi/x/C8ITsZPb7vkJFL2UDN5XxM1/W4wFJH/ehvrWmtbgUPNPE7JY
gPWYE52UKFQICh+4jL+/N1/on3GViawVk2jKmpciXurfUWRNz1bsnMj9/ZdutBXS
fEY43oPqcUfo4j5b+O0F8/JXiwYklXlWSz6iuviwFu+Y1msB2Gn0Ct5ryzVRnWVi
MhZTUOKWT0Fgnktj+Vw7PPfDqt1VJiEZA1V3S7luTKEfHXmJsURgqRn0D3Wvb87w
iLBqDMzw9A7Yp9aYE0xoGdoxDhfYQOWm4VXesoa11lkweTuiZ85kMwbid6SvKnjk
tw+3FXzUloB4WFwibDjxinUKfMzGoL6KfgDn+/8e9BHLlR5ofwFj7l0Lsj1CV/W0
5GiE9zlfWmBBJ5OR2wj68mHNd0Hw7lfr4yhv7Ra4TXCTGfOBr0b9s8GWGLtcfo2K
JGpRAEFRacNeU36eSJWefJPjFfsrQocr2fS3UzAFRCtUxwrIAOYvc4/o5xkt/OFP
TkA4vhjq4AcHXKYDvahGgc/pZEkkNxTrLmJSNr/kAARNkJBxRV4p5nq9nSnrcVyZ
I+NMdgIg7yVnqyYh3dGYiI0D3Yfub1kmJ/ExLIomu+eMpd+tzxdQsqjlaxHZlxIj
64YocZECaXagQt7i0qIbqjn3elbX7e9RUqOL2qOXKO+8JUnJcLCZZnkIxq2XG4qr
o+fmK34qtszZWxiJZ0wiyFKizDhGXp1iD1Kam5NIEe28qHyr/Ysr4CRkKLWFuuLp
9sqr/XJ7mul0ZLOHdeszFLkxrX8sDJPQr4NPjEgeGvBobwZrER4/xVF9rqrZvo5f
45Yya1QcO9jozxjiDpVMv4FhjbVOiBZ7e6ebio+eQb+4rP4H7QFAhCLiKgKO7fvy
7WmTky7gvtRjI/ALgq/Q+riw6GVyOV/43FI4uziLSWbOQOsRzrwzuESy31Gq0Qv2
jIYAgWGSNoLIRZV+/gZdhc6ABjHOcaXNny6B5jp50p4Q70NOQyssspQUZoRTN9QT
rPCjAH7lM6t0sy8pvRPGAtufn2UgYY1PMYDv6H3PFTgZEcX5TBVd/85gtt5EXXlR
Y66HT53BK0BVERpifEk190rrt+N9/h5ZtLHW+MqmhhvtFF1izt8pQSGVDhIAHGJe
9FX5t/6b+HhxMd0e7YV7UB4abXZ3os2NMe9ynqu/uv9Osq2koFZhq+0Lmkqj5ztt
yUfFeulBoSWogyybHU2T9uKjHPRhF4UZua3NVk+HMtcpdn7yHOojTtC2PwU90J94
j/TuzPjRCUAf1r/8Fpb8/CnzOJ10Uj5Yau6h509qMWFWA/gtqMEA6jGPAY6CF4iC
DzSD5up+6TeZYhzOdWUTNmUtJ5ZGHIBySQIKqaNibFWzh/PCGNAx9IrqsSN3Vps5
vooTkQBurpWIQe9OzdCadoF7LiobuyWjMNnghoDLS4UX5s7lbStgr/TcYLy4WJBG
bMmH/pxrvw/4LNU+rwSDlKaM7SkNKUaoDxMup2TxHheCyn8s8RiMJkRtKVmzhi8K
7+gKrZ/1UK8YVQe9H7Gn4IMuQIANb7i2vaRhBYBKXarLxvJNqsin8V19kcT47Hvd
pQp0pvKF92Z5RelZi64/Mh026MSHHRtB2d5Nykglod1Asy8IiqfHWu4zborb3He7
u/aODZttZHakm8/nivFxhtq1ZE8r568AQNjMkSlnD7avAolxSRhQlVt0AwzZEyTm
Kq83oG56Ry1nmh6KoBe4LkbnaFaGq2vSGhQ0Bk6gZRAa9U/jZNyaT3rg4fkeWbpn
9FWMaWsBOXYQRWuYqhL1yU8dajWA4iLvtY7y8Klxm0GWMsSjWHd0dNIYnSm8EQjY
QizhRaoRPBzF4oxSbgsawedYA4d7uARywJUtvfrCsJn9N298hgX8g0lYN+r0UcOK
qCqW3jdyCHVJuLOpNMq4CmTQ4yjXwJNWiy3z/gwcCGLdW7mo8mV2C91WSFOccG5Z
s0YcaKgaEJYZh5C4D0T+PGtFN542YuAsImaNyzhW/hXA6GO9VlFT3oAaSq8GpO7R
Vvt8PXHUohi+QVMIV9IfcoEDuPMKbsnMDTT6tj+t9qxT1cDdiZ8O5PlurLGOJIPG
PMRt7yLK4lIMFQbnUKP59uUefsZfhZUDU6yVP2/6qpMdUap1oHuSJ7cEQQHagQSz
/NEwVdYctywrZ8uoB5tpwluu3d2BBLhRFPLljpeCh+1z4fBhC3Cn/5BxaFq0SRWo
QdkBl6vOOUlr6Kei6+Af0NcSXcOEBn3MFoGM4srvC0GHgfiZGoRKMceV4kQXekI7
pMDLYe2TweZm1iOzNMFLfG/rWftvYmCcmDW2sBt21mjVIcXxqspqT+Mq4ltOVRV6
QwjnH8NVvkLWcR+VdTM+hoYekgWTUJUtZ44hVcvnBOsqpgFxGhokqAhDMOTVFRTd
Ts+s5Q3oyKRmTuglF7rVEwFWlklNS3chqX9X5QfpQudYPl5gzchbUOgwNqR45t1S
H5tN/TbxJt+o1uP1kI5nkeXxh2CcDhPXCzfspLEXzUB/7TkXJZZvB12ZJAs9vuB/
YXq3qt7InuqbFNmn0CakBfDrlJDdyuNKc2fBF7F+hPdMQKfEKLSh0aDWhkbF25ls
azdAzCDX8a5q4S+/Nd0PsEaEbpzZ7UTAgAS547/Lxv/Xc9zTD2EpKeZmV9Df4Z/E
ZcFXIpBWXlM+iAPjX6fGgks6hzatg/9BKTIVeqttehwhSnh1FfvnQnDD4xilvluz
Hy7tm/zFG+gdVJzQ6AiHZpBUQocFkWZJZQm736HY7ejbCnmuUPLOblgE+Mj9b3KL
f0eMyrcs8ychaDlhJyI/r/m31QPj2nCvaf9b2KR/4zLz+G/+fKoU6mOpKJnv51FR
2gnkxkEe+iApE6LGyJiLiqUMdCJK3Htcxg4x8bjnNe39qzNuuaxW7eIrBxPe8qw3
pH6Lt7D48FMrnJ7l3XYSbbyt6QBej1Ca66hO1rnBxBqFjd/HZKAEcuQkr8ln4qoS
ee2r6cRQBdn45sGue/4SB0fwVfXL9NFD+/4D8Glb8ZRrX09HRY44qIG2gH6kQAYI
dEb0Yj9zD+47uBFA5NkGZwnezrzeO+LPiLw4m3OYoqs=
`pragma protect end_protected
