// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nTmh9b6tD09D4P0tMgeSXAHBt1Nd8YGZq5VpY05SFqXgFw16nVPI+bpGfVsWt2ix
HQY7NTrLORNkYDwrubPeQ5IttkbwE4sAqN/Top4WYqCUXrpys41CHWdzVmioLr6A
XkOnUmfGjAL/Cg5nFaUo4pegKWpPOG8Xztdu1OEiWQc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5536)
AVd/Pgh3Yh9o+4nJPI7S1ClqmjdFGdBuZ9V+4EBGCIB2pCO10qbhNpoEsorX0y7D
2+2paMRaEKotjAvPiQGf6IpZeguYQeIvPmwpGedI7O9BCLEIZI16Fu1jexauuc7B
I59xreNtxYCzgjmaY0JhqaNi+1M2RsL+/TE/t8neMZVlmeK3YiFGpOSruRIHNwDk
BZNYU4TJdo4b58LA8irblXT2JxgNpCrQwcFZt8VKYeL2kR0QZmlzzuOS1yUfga9b
HNXYGQEFtbi9GmGxzGpUq9saQypTa22dUX70GUtxAUkoTys7LLHAIeG4enMsUN8A
sviw3NDfCib3qaDTRQln+pnsgWnAfHDVWx4AZj3fyytqMFbDoFU7pEz+TyqAeaqI
fwlOXdt0nahd5hfuCBzrKCb3ZZejevHrhY0xlaz9Q5dyaKHtPlzPMuU4Q9ud1s8j
RS5jOqwBQeurn8RhSAQIj0td0YeOGkjZE07EVw9iYIxYJsf1OmDDW040T8FtIY6/
L7VfQEN6qDqM+k9/5ihvnjuQbtdCZVEespJ0Dyu1xENXtoSqS+5uT6qZgNmv5T48
HCZbGjn+u2kodXXd+mjH5qizZAE+e7poTLuUUmCyFmjmrjzFcYMAYjJhEqvrTPf8
4jDymRlUICiS0jdiQgijHILHlOCP+MOQGczZ/efj3dtkEENc/jOC9QMgCn1FMEZM
tAHOF8Vtt45TFn3IFBl7m8fdiXNG4fQBbFOLR41ZnRrUfq5oiZUw5sRuW58Uzju+
cwBLcIaXXjTqPf+ezlKYyukjmBXgBIXPwr5nsERan0f5r65/AJk03Y9nMaMrZ+yt
7H7iSY/3oLvv9Gupz+kcFOWZ9SdzdP0fwgo6bksm0QfU3d1R2By1RCyxXzNiwWUR
wIUykEAX27Ddg3xVGcJBDd1egxz9BpknnbhVgmGadn1i+m64kbHEQPKPaCPywKLb
5NOI1d0cHYA7bXAziut1i9Ru6iPXQWd145nrCdZ7gihGRvbYzg4AGsuRfjQPH5n6
BZvs6bjb+hD4fOZHrMWKUT6QmtNr5k3XYXEkxgEjAkeGp/jlzHo2B3SmcNakTUgH
JUCBXncBMJSvmQMHUaMgJQI7CdjzNjosUhsJVgjY8trFIrv/GNqemRDrzg+UPPoq
jTAYqTpinl1EFYiWl2lbgxJc9in9FnvIN7fWg6Tm19hR9xgztuW73W12RLC77E/P
U3LiwioKi49dHpjR+QSYMyPc0+r/ORJrvGKeUvI7Ag5KPyfRX6jDuY0ybNWgG3XP
+qkWcQy5rNsqF4WE15hT+O57hJEdUSffEtvc54XnuvrhXYlKsyQjgdBvUwYmp0Pc
7neribfpzGF+920LLfRdqsZ0oCb8SY5XG4C7lHLB43OoQai7m+AyslOFwS4BqawG
FpwBheKtUTuo44FeQMraYemppnaEp9PbnOAHtGBYcXGkvSCRlUilpgJ4SxUNfd9X
KmNTpIgxFgu85ja9MRfSSKNnreWyP9LrQP2V8kAXfomJA12TSlwmDqq0HnAjmR7o
6p1V+UrkpHXMGuFgCKdDIwhXBnGrfbN1kl2FByukVrm8YadKAUJzzEur1qqsA3Ig
ZSlcWZIiEZCqdGKep/19q90DPkEWnd/uyL/ZisrDORkxv1OiD72KLGejoXXQZ0OK
djoCv/WqdOrLHrhLJeDNg8v+dCwmrq8I41kUHQmePhMJQ+FW3WcB/qax3YM+lrjq
kIpGDfUeWRBhXJNTMAtrnDYI3Xli9HsGmK8soVrJfQWcfaq9AJwfdKeyL/9AIeqr
PX7TQ6vi/+A1vandnJyUo42c6sFAnkI5FemccXUADZ9I1xGFxq/eUSfG6e0VJWO+
DTb1ue2QbBHkRQWERwtancOuCWWVVCKUVHbPQ1o1tE2mju55hjyOnBrsw5x6aUZj
MMO1pSUNGQ6JvRft/CF6OIWaTQDhLEWwZkxELqudGKJvoR38GhI6CP9kc7MeMICf
gW6KLM7dUf6OEF6ebyq4u9N8ycpBwHfODUHhBhpavJXe83fk9Yb4p88iJxTOrJcC
q5cwjcRIHQQzztEEs5YtrDYU+FnJySV1/Zx4NQh2M84b51tgaFHchbV9/IPQM3Kk
D5BGdTJo4cdsq/hX8PLZjsYav5tApkRkpy34L8sA9uaX4yn5IjrqY8tDGzaZ1pOU
hM9SdG154KNEVDf5gBYYKjsGwqC7ScphvajUrDJaajdkybwyMDfVN8qCMO1EJZ+v
z0CjRDCmm0QHxy8ga26yEvlVWAnLQBAUNKJkvgbMO1NDKdrabepviyYcHlSfLfnF
oU8cCzipPuB2D0s1yBVqBWzT2OV/LvXrT/vf0k0RlMYRtU0QB7+gVAAiPtuP6r1N
HfIblsOAc+xGQHkUjH89KELUmR6MN2eh2KTbKTnlve4WNQrgOMDKHwDMlg3eSds3
jcW7H/pBZe3XSrZCgCU8toHlwZFFFiMVbMXGmVPunQiCiJkE9UaP2Ck75ILLitY4
IDYRgogSxTXn6E8V24cNay/YlDrdSyKbVyAomHjzHa+kGuVVUIs5n0LfIypLMJJ9
MKxrxNi0biZ3bhMMtG95iRZ23QT9kEF9XK+RvXXi2ZYfgGUcmTIEfW/r5YYT5gzn
8e5oZ+bVhe0P4YRY9stHGgYPP3Bn0etAHzJrMIqO3X/uoKN2m5yM7AUNfNOSAvMz
zZagIoNV+A5rHNl1l5NosdzYRDVQR4keh0pP3QoEbdhKGMxaFedK7UYdKjNMKudw
pjauKMJjoc4KTjoidkYLLXbwcLnOTs9K2sLZOvulhBFw2+egVe/4TUG0J/9kPUR0
TwzVxTJb+942ydOOjY65XNZS8++++nsMWkcnSfIqZKwZBZTqRLETRnY/TE/Crav5
eYMnBp3bAR9bkvSqLBiDaDANLcHwF9g3KPqiYuJ7MlkMFhcKHFVy6Uu4SDdi2VmT
E3Y5a4GvTUbHffILR8TsKXC/6/E85Umv6z5X7SsO8KbpLtyX29sRHf3GlVW+Q8S8
6CW2+D6FJXQ9Uu0B4JVKMMqymL92bbpqHh0CI1gA3zQlQcJ+lw8VQ71HLLhuQfpS
WgvUIfwX3DqB/LoZD+mYw7QwjCLrNxYkHX8wIcgXDSVp/3votEKMlKiCyosmtQfS
G2ffVjLx40dAALamv55cenuhLt2qiDQhENpNCNwdbEKS1V57QDf48mIQcXXZsI7y
AONiKu67VYyTUB3CuVh5Cycjn63Td8W+6w0D1Nafery1n5gnj3MWlSMQqpPpYrZy
HFBZYk3vyLCHYrgK0HqU+3d6uRbj0HPj/K6Hv4JvKsdHHx9ggonZIyPBG7TooWuH
EBPVpwxS0tSW8M+eLGPdz8OQ6yyWNkfEcWwOwirKwAOm2KaktFbwAWP2JgYyq+pL
4811LMuuv9NPaPfqKuEcb0B4y3NMc8g0JeUKCgaZP7g/x/JyzcGzbF+YkHc5QaZJ
smJLNu99loCMzIN+wXFbFgXabDNnhPCVJHN++o50SfczUKXh65/CrkN+MTNtuSc/
0DDZwYRgDeJT5R73qS5dNGgdX865kLDI+LO61pxmi6easrsKzrJ8/+y1ZGUAyyRR
HUiXbCM9my5d/WAwJJfxcDuUruxFru/crNLHoLQehRNyaVsLW5Lb2uUgojqCKHa4
Dd7hImr2qdSDG5ygsSUJJ7YdSfgcQgsdYSa9am8AFfZ2tvHazkpj+OQA9VelNQBj
Y9UyDGJovLj1PMKXzfpYZgmxBIidgm2gWeJiM/OtRVdbKv56tBKaMWCOFLPqX9nU
vp9Hi+PXUlE78gbFdcoQiXNslHSWGuQlSUV3JhTzfLQ3NQr5S+bSwgxX31P3+y6g
NgxpWlU1SgXpVTBjbLk0HtNb7L9sEH/IxnODlYeyvph4mM2pa++MV1FoFXH62fF/
Ng1YOeqYyb8kJXJAZdUtBuy+eGXDRLgtQjrGgeWUvX0cBsCBFEV4XYbWYXXtEck1
aW5nkigkHRLyDhW3A+TGugOzLll+m/4feyCMaN4GFVXeNP7IcrlQ4wH3/hUaPdGD
50Evy6OYB3nPcLRbHkDMtNK8ITOtHvJ0eT+v1TK/CL1yzYl/Ef00UZPpnBzO2lFr
p5gZko32McX2n6qyfrK83ikYkixQ2wblJ4IBdofjRRuKOmWzzvQXVIy0JED1Q18t
auQ21bg2V4/K6BCso3RpASV5BDvUDQSemAESshWCtlsimHaq600GHBacm6QQ359e
is93YCr57a/i3d7rCakdIbZUduo2F9KoCveRmZGORKDa46beHLBNNzjHiuApwf87
lODhDYE2qTxy8jd8cPUWP/3/IMF7hy6Q7QnMwtrSmOMAe4ZBKXQGg5JDoI78jbIE
4E5zYwM7jIzs6KJZIziL9eugH+JaapVt2leBJZZY0vNWs7yHe1tehNKza+FAAzHr
FlY+9xPQI/CC6pzo3p/+QXEE8RJZ3weKYDzYNlKDqV98enOLxB6LudjIA5SivfEU
h0EtTCfMN0AjM9M0JpJKcZcEbyoSXbnXaon0UEErjeWCiKk3LLOzqAmHVayt3FVt
rJ3wbeGk+8XWmjT1FVFhhfXQAI3++1HlUA+2dTL4zZCYOVo1UXUuRYzYVqAwf0am
uWjplC4EDYW+W0k6mtaSFZzzVb/JZqbe1PDMgd3rcqZ5MQW0OMVLFnJcoS+7vJYf
3C3+bW9+pjM10sopg01NH42WbGIt2aE2xU8s+KPbvg4tnP68vMU+0E3/H/he84ri
ycW6yXQRgpifnu24y9bCLL+mQD+6BPe9Dt6BMt3Xl3i4YlGgozlaY0d4ODgkIQfT
S8AdoN7TOFAOuoC15HWu+wNafspIVCc5qcrS7p/8EALzMJ+5hFW0NrZLE82rxO31
nNpe0kW7k5zVyy5hakB787HSqWvniUCU5lDpKQmCt6j4LTPvRMrqu3ZD8vuiEqkM
1ReZf8Ny92LwNusNdRvQdEg22tSaVSa7TcFaJY3cREXEsb8RpwVjCXuimoIT72PM
/IFlS1m9VF+rJO5eHQA7ZKAfmAuBBOMj8grclTAt2tLk3bquVY3OyqIkjhdNZu/w
8EtLqxVZ5QseayDFBj8mgVkW7WCDR7IogtIBhnLTAywD/WGuuz7xOgNAXO3fcX3T
PV22uZLn7VNdcmINQxryCaU/riGL74BV13w6PqmfwPSUbiG60vS/DM0Vvv0Cekc5
Myc0AYEYtksm8R1qhNZ0evGCR0Q5VAsUnh5fwFlAUC9qIaRu+ElGZDYBSSjWjHfo
IimsgFr1K5zUsbhMN6yTdCnNI2bseYLf6/Zi9l+8antjXvaEhyD6I12VotDCDu4a
fwSp9a3OhVxcGeqPhm3GGrOKL8KQofIeRqP+q1CZ+JAU0oj2NLotSez4BqnkzZVf
ft31tdeEY7cBJ9iY14822gF+8/UXRcS3QHUR7iVSj1jZ7dhPCMzSTn0+Jqxd30L6
eZjrLdxHmCcdbX3odhuXCsRFL7MwXmKydyf2mXDWFZvm2uautDVX7TZu0JjfuETU
YKxUQQHqZDSoIhNkyTuMkYRE7OOidcY/qRwpHWS9RxoggLJADoShUs1+eA2EmICB
MReFnVAbZhwKVkt6MH4T2r0NW/TxNNoGW742SmM+qAvx4VhWpcj/GDl90PsOJVqZ
X7PYALDTxKcJQghOsXbiD6JZi21wUrMOvv5git9b2faza5+7wCfaJAUwAw3UK2vE
Cn2xSFwrKSxehTrxKzP+br1pTHIYaRLD9gfQ4AnsLWtqLePW1PxMl1fhZSB8uFKa
DuSbDr9BK0VjE8DfQT0PHUCfzOhM1lwTo9pryMhukcivcgrXKCXQV4l+zEsBrpdv
rg671sCHvxYRU5T57cneJaiTPYwMSXhKlvDw45Yl5L3syhPAb/zxx7wpGxeUpNuQ
3XVUrEXN39JC7dxtuVffP3faTtkpjefU9YKl19hOYy3NsjePZ7gPhTBpKDtXsAPe
7r4RFyYCGUoy1qdldksREWp+CKxrrApFtI1Uc0eE1xVgN3txKjLobRt/Gds4TBcw
Qel/Q0BMjSekNWhqRakUDKTdfrEJ8NY8X+7zZ50s3H3dp2fF3iX+GTNPCyS2qBT+
Dq8MxAqjHdqTy58fGxLm3x/YA2s+5eUbWejnaWUL+MOPy83PXny+e7VDHlSZgbtJ
vohakX6xbG1nPB3LB5JQJXChDC4bmoRAL/kw4hN9MGY4R7br00Qa60f5JHd1VVe4
RSyvY07mbpZhcOIcYzVl5Yt2IaDRq9gGgPUk0XmLoHwFP2L6utb07i5ffewSqrNm
IspFvEhPwKFpO1FjvYHCO0aAJx1wK8qWq6vaD/3/xjM3jC5razT/6QhcG8MbjBO5
GgLHNJXoMeS0vQyEt19qB9J1wbwnOVuSFH5Y7dBcXrYuZn+6xxWoPF9vGZiyGQLq
nuvoNVh/s0sYEWgN5dhB/dQaU0YcBYQYQzaaBH2TwIRkt253HyaIsQiIa5ZIESL9
TgIhqk5pn31aSJfM5CENm7ccx406OkxTGAjJOqih4RF8EXxmpS76BrpYJ+N3rDBq
3T9kF7GSvt7ckS3qkPwkR6DCmf6arU36pBWGxfYCJskio5aKx3JFei0kTNGoaBDQ
3iGLNK3ulwy7kZgwi8f+6yME96xpk8TN1bvvyxPLvjBAPzh4XELqLYoT3SGbVVyL
wZRdL5ctwISgJptIiRO00uVS9vrNBcO++87JsCrzzC3Al2LDhMZEAzeQNq/jBvqp
NXaZxJSyf2t9p/fNBIHK+cuXY6+cbFDK4lJEoX0qA0RBCH4p6TMPLIBlUG9e3A5z
48IxLcbneQqHBtN92wIouEWQobm6eECsKY5/+P15d4Cibu+q9KVGX91y4is+c2Mi
C784LKiLY/gcRUdRdJMckVNbbOXIktyi+OZvK+ueBUEY3QzovbOC2zJ5noAwCPOZ
4hqarXIlLW8cLBfkH33u3+FQ3UfJE1Qcv57tT7sO+aGQpLxgSFdOW7IOAcV2pPfU
8EKtFR+RY8qQw62HmzBNf4T9ONfyDpLGyonRJofAofrgCJpoVFl0yFaruIuhI1Rk
CQI+qdKdAcr1ADAf53NeVrcIPhgwvJ49RVtpQjAy8e0ZWdDVIrAcQxSoSPs6aROr
AmZBxivr4+1iCIHAoYcpZh57zOo5vGffLeEeBcwyKWxvBX40B5vad2/okx+91uyj
kV5pKFip4PpZEy70ypAPzs7iIN/5TKvs7fmSH3gD1T7nU0FSoEtHD+4rDjfwF3OA
HD7orKD7qe7u5plqBXB8+rai5DD0G5OnAA4UE31SyZwsfWWryGcfL9+3mgk31YYF
Q9A0Jws686NNv1o9j4Hffg8vyYgPVH8UoXBTaOanUYPCDeAmhCYLregTont9V2jv
ze5CoYwuXVqHT10s9zV+Wg==
`pragma protect end_protected
