// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
M/I6JW2tQhkF2aNOkVhe5t7ezqAxmERX+cRaPtGoDFhyQRysv23JLnIoG+wn3qe1Sq16TGKr9/pN
1sSBfxuRsLUX8LPdALCJKw9CQxcOZajJHXdewLvYkzAaoWp99/uHPSJhS57mqA/vPjNJfTuFD+1/
p+0278b+UXcyLV7MJAToEaMRXMd5CYkxjnbhGLbuqQrZSDEQcvhVuE6Rd2AgZ4+0NxBSd3sGeK+/
3jmG+cEjqlLniWCz0O2CIvL4FJJRQNI7Hrc5vEKZXfB4WRD9fQDFNGNMKDAE1ySmQKbX8oXUiuJN
Nz8AY98Vo3eXLkjBiC6CxWeo3M3/c3rs9fxL7A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
w+lmT0oLtKuyNh9O+tPYj+eLftlo8wRvp+nAhbLQrY8w5uaotIT3nLCeKS0IzMfKZfeOKrmpFW/+
dxO6HGaCbVg6XUvk4zn6werz+92+8SqiCe02zjFoQTE3nnBb+5GDWs/l67Fyttuw4bnYp8HOQ2cs
lIWUqmeQhEeX2VSCCl2au7zgyhTqWXRDNpYa2Rn9E45Koj4TvH+L4z86AXUVKkzcY9JqOfQJs79q
LO2YG6f6VTpwZKH1yfR5y1sIzgmbSaQc0spqOHjzKsQTSWWAD5Z+art7XP1D76NvNVMSFwtX97Fy
U2mh7TOxlIlZjMUtFblVUkbvJsxEhRWduAMYwRdmsL8etngw6dzl2INfG1EwL1nIzTmne9igNeAB
UoPev+1VMI9Y5znNwhhPyQjwbmZw1NDwOWc28plI7/yRqntRXnOf6tI93/prpxbxICZ4qZ0MdRq1
Zjl4fd+dO74s008erGtbh+LcXIVl9t5k/r1UJXUfZ5ouz1O3KcGir0H/vVwaJx548hpVLpSdrVyc
A6esyOWv1h56YCUtO30S8HQl22Aum0pOrdDqoncH1AdhvBhXm1JkB/TtL4I3p6Y0AFy5vp0NPrW9
V1E2J/ibz3bjkgKqRwu+I1OzVuR9fXJfzWmOFQ67+7oTGZqO9dRhSM9zOpNW/+bxkPfKY3s7Im2T
+rTAx5GQnpic7me5mqXwQOo3LUtOnf1r9F5TtaOLxMUBrmgbaL6vDdG4EN1RJm3cFizZLfc5IhV/
xRee63lk9xlRR5E+WoPa9g5G1h3pZJsVWkeevVwNnwfhDszQB6DR8y87IWO1pUYLgU7jbw59Nee3
vd2M+1aumjNkuAijr+w6M7lrPW7JSZ1DO83w3Qhk9Ck7+3XOUFkh74G9yCH/Z8yH+ganff7igDRn
hzzUWZ8SZrprIo5lai15KNQuzWlOUzgzepfYd6NIKYG9cKgCt4N8sbBD4/joIHm5QaeksCwagGLm
+TU3+PyS3oMLjXimsBth1EGhJ0rZbrjVwT4xE7yyHDDLjNETmhI/h/BWT2wG9v2i1IuJYwWeQ20D
jL+W+TDyXvywZskSK6lWqqq5xZ5VZZx3WaLYj/qU8SGenURhTBLBOKnmlksByI3aiOA2vjhUHtbd
oo6rET3D6vPiXVGrZs4wYG4p+WxyxMFP7XtA8jROeoUoO4+lAPs2mIB/kq44Ni0MeCpOF+kMBxzW
F6Sz4fYpImOwTjn4gVTg0vIndstxMIwlKAFWiEMZqai0fyRChv0uTuOEcpeoLzAbPbvzRaIKSR4H
XmiB6IJJJFB+2cberHe3wI00ZLPmmh9OuBDW3KvtAWu8aEsJ6CkoUeFyMGFuBr2wSrcqwJTziYos
ZZ9kwoOYT0hzZuBAVz/u4GXDfgqNasVPDvHdWc6YlHu6m8OrJ3b9bKqYo0YWhonvX54AtfJ6Vn15
/KrK3bBYNWS+uM8hsGGIegzmSUmyRYW8ypHbK+U+49oXy8cLIcg3Ul6IE5l44RP09kSwNYT3tmWb
TMUXTTjuPIkFrR69FT188GztKzS9KiVC5QRU6Ji7FTbH0V8EtCnacPSxg02BTpkICf+ccLIKterW
Tw4sgbA1Vak/rgqqfDhsMl2jSQJI3Pt0QrsswOrEe9TFl+ytb3JzbNhbZ3V6Topwgv57hJanCHt0
r5+4Y1haAzya58B7sNf/KnZl7dFjQZSdA51GPzYzjle5lWbVZsByTiPnf+pStyyD4z5U0BmRCebO
rXL/hWvXgGRnHT1ZkoTPohhZlUYvMJHp7zpJpFUr481HDZcQPhw7oJ1hJXBuRB4aSnetMgtMeU7l
tzLwcKlWSuyQZQ9xNZDQdmPbpBQLfAUKX/+s2dBa/n4wp6hnlO6hhsRyKEZCVes7CP/jFupmg6VK
iIkXCVssx/glL4JT3t4fWzs8N8Kh0+D3e05PLJfEkNrS/0QpxhpNnJ7rnKIThjhD5zJ1uX70abaQ
bd+z9EbQ2NzjbsvchzuVe0L8Hxfku1vtsqPfNgZ48Pal/HIXdfStK4IawR/4FYLnsiGyU73aVAT+
ELDFXms6NFC4mRLdaYm1WGqReD07v3eFN+fceV/F4IINAstcJ73MWBORGPA3Y7Nx+L8H7QgjLLky
os5iGtmlNUIDhw6yMVKuWNKPBLMMb8uy0ihAIVrlbawgwBGUW7bSIUSBL/LupbU/wVupEgH62aZi
hWqJTHVOwtK8UG9NO0WJ0rAvXnbA1IldNlRoQ0bj00t4G2kuE7hW+HPAJZ94e9ClKbvxagDu90O0
lUkj+PFHuGYwbKlrdUbmuW6jGUKfh1yJl6K60/2EUuDuQnOMB3+bPVe1S+cAjgUOFHF+BArA146k
lfLMBKvtBAiADIFU8X8oEgW1OcIFCUNE8iknMftc/awFZeyMWSBcfSSq45TzePCNS5tV28qMuLal
arCv4/YWKGVsAi96SD5JB1WU2/3iYeFcRjX+tk0sE0somu+jv+ji330/x4wTL4NreJ2pvP5LpRlB
HHO91oZvGrcSakidfZkDK2s2pEbsC2ZbJVmT5hOBM1Mo39fyybAu6HIbZgxAgvRvrlzoW/lof31V
TTcaiuouS06KbvSWemQPyRm+4cRz8TR2NACaUyWtHEJyi4VR+baM14k8atz50gld5+VbFj4q+cbt
1zgAZfsqN9wELb11NBIrdYuEfFA02+LTjehmS2Vvde5z1SRlBixA4FyZtt7MgCgWouPuX8C4Mk64
mCjm+6kSoDTjKos+ayT8GPbAilHdq4AOJ/ZtfYcQwEYEUdcjgDDIigv7Q1LvvyGqszhjwQ4mr50+
HU2g1G9QkaaN2E32DltX4W3SRkU3OI/0FzSaiBeef8hZqm3dnbYWp3ZBM1Tl+FQ7cMzkuJShLGrb
YacgGBfMpZ0SqFaXZgfb3hCloG6TNM7SMRuMZq6/qwkHLb39Sf+3/D1a+Em+u5nEu4sa5VMBtPGv
x7sN7lo37LE37H10F+6+1IhWGNSOhi9nzTUwhIm45bETTbH+2JON2N7+X+S2uCil91Hw8ufeJm6e
1tnITC22t6ZsQ3PHW1aa9c9oZH0rkLS9rnJBPbF1N/NDRxzQfYcj02l2//3Q+fddx03GyYLa5D8O
g78M2ABsUI/aID3fwCXUT2E99XAMDLYr1F4mTsttSnu4KZ3hzpjQjrVDhjfCJGiwyQKiahrTMkTH
VL6/OEu2CJ+nuzibA0Z0OxtFS85JceLVMUFF4tg9B4bo0aVsomETs/oFovnBeuQxDvFJ04RpkgMa
Cvti+de4jXgCxre3zG8gx0Nw/lVTueh14G4oQhKDsteA5KLYROkrOt7hxnLth5s1o08jH3svH6A6
plefYnH1MTypdwnJxBct/4cijFza9XQ5OcH8vOyL2ylIRx+U02dLqtfFvG5juTY7ZIWJGHq360XF
kej85TOTcUJe8uKx/qoTKPPJyFUyTtYKw1kIG75v0X8MkQfU/Bf/AHVfVdx4CgJ2RUpmk9MWCV6r
J6cMrWuHsdx8L/tjvmkK86B12vw5XahDcbqJhC0JuQshx4cCgeYEhWCcSFYCMTs7FEnbd4C2Dq3i
Qu/LnLqPUUNVKEGE/vRO52P9tOLzwftkz4cqg6NleGKb9J9fK4jf+wjqGykIXYaK/Dte84epHhAI
xnw9NNpSQsgmWqr+N57pL4IcgYbbbcd7reHVJBXutqcFVsDGGCcsx+yEwC3qAC8YWE4wajs8oI22
a3WZ+ew+usAhFDCssiH3oc3dG+t4l56VX08FIvQwKMWIjj153lMRtFVQpHgOklQ6awgfyzsTUs5x
TLOutFUNi46raGv5XB7shuXOcGQ7GAM9oERug0wYNKJI5aYcwVcoudKUVia75Oh99h4eMFsgcL6+
XpQxdm+ESopPY0zKtDpQpJXbvdaYHUxhoLzRkpwrI1AlOlqWm0FZBRqOPMLeoUz+ZyTUc1rIvKMi
OkFv6SsgopwUqaPHRXyGkDB3xieA3Zu8C4ojWvyCoTZnVW8uq6fcnQo22f9ZjoSL6wp6A+jMQJtk
crGjP89paCKWWq6k6BNNE8TQEYGSCo/GYRJYVcs3tMtzUG178OWpgdEnn7Ezfx77I/ULKQnpXZ9v
hbOo2ORF+m+GvmjWCRr3Mo4rprCfVtJcIHrbjX10vWRgSHrovCr8TdmBtjEkv7/tOClHX8Cf8L7d
uU15aeH8vvObxj+Jhqx91/i65Xny2CtJ2fg2ffQsSPa+QnbypsvOnd2pGzt32Ruoi0VfEWXR1Bcd
R4l+/EF2W+50TL2PeHzeKsplbZmoketpUYFAFkaIc5KzYoVBBM9TGcmq6G4te8c0anU7A0SReKJO
YNKYtjeC1nkqt9lJhm0pT7CAyc057Z/PtG0fhqcJb+ywO41MJrsJbkRPYpdr4YYkoA4p5QmMy+62
izcmALSTn022qgsjy+8LQZl+iFAysdMAEnX7+CyM/3b2/9fspkrpG8Lp3F6bm1UiWramqOIHFVMf
fCHVjKMrRAsZ9t3JT/ZGYSuDvXBUx8Pt4EOK6o/5Jt8/pE/CXhrBFNtSnbEZHzVxJVj4Tgv6Z5tM
U1rWOcv4NASsXjvTluy6yqk+mm6Cgfxi2LUzsV9rWRu5pFn1oMENWPJNOBJnrZF9KHLhuj8LuSZw
2mgDLqNRkdsbIYptFcot0ln1IOlEtwTvcSM7OkijUjK+xFI4OaAYs+tWoSYzHJQLyBmL4VbrnRe6
3r7FODaMozmsp786cya8iaqQY06eRKT2suvKe10mVG40MDxuqxkTc3e7DRyLS0j/rq430O4qid1X
/Tdnl7uDsI5N9rTR42AjyMPpPqrtdzFBFWUR5AV0XY0lwxAH2p9B0lTqJs0OFN4bjaFyKF7P62Uq
eQbWfnj+fG/fcJBZCn9ST8H035pYdEBBRYYqevMOKiBM13s035Cou78rYW74yUSSTqqeOcv+ml6Z
O6HTk8X+v3i4MBaVco05qoliGVlpBcFCImQ3QK68u7/42AoBXOLid9Ym1TPYGWJ+DQNSen+fhB04
udNu3ICxCw2pxsKDvG+pUdqWp7sRQOOZcm3q6IbuQa+oKnJZ6h/Fra3ysLh9rpI1M31CFQHOLqaN
V/yUCRO4IvR02Jh53X4qhuocXx+r7mfvaBIKCEDYkmGLvyV34/k/tnGZCo4bIaPfzv6fw+36VjRy
w1meeViHZWJn98j4ACOUifZb941+HO9tGDfWUrwGWHFR9sDaI3cGAAG84oXDnfSEMqAA+0/cs2cp
09nVE+NG25A8c0mELmZRyq/rNrvryZ3ze8m36I6Qi/KQdMi+oNiAgSoj3/iq/gOVa0+n8PNaWjhh
YFv7Kh//+cTrrdBhHRG23G7HAYvmo0yHA2hlSpJNsqHVRRNeDdgqaOWciQXaiA+ItQNTCXZul5eF
mzW3Z0R0CmgjDCBzZXt5SiP7Ch4ACfU9Lm82N8L9ox7B2SdGI98pXCyUEASKahMkQUtIl5ryH4/a
YRtgxyaN2PKiJyVEbxHHNA0INrEM89FSI91t0jQkBipEO7+2bEXpJR+JkB3SGN8KdsGVHN75FDp+
+FrM30LRQ0LIXSY033JGuxfhRw3kLG/5gIYyXb4dQdiz5VQyxymb18gxHQAi2ZahVLae1zWQsiKY
l7gvQiHIQ+n0K+HG3CGAatK2EKfik452lGdn0yDMX1P6HkKcI1Vw/p2VnQNXo1znilghLCjihm/g
0MuNrnoBZF6WJ9Vv7L+6Eg38Bb68IQ+9w2xQCr+XaQpWwWd+z5oKArtK+OuLdy03lYuh/PmQinWo
N2Tz9dgI+pD4nkPneKxjQM9Jtn6wNzUZfz7LG7CGAyQ5hlVQnp5MaND3nH2zPXIEADDKrUiFk/W5
blil0Wp+Dx2VQk+xjDesECmPFvIKXYi1brnm3DSxYg5ZJtsb7fEpWRzhlXo/2JaER/KcZeGIxRjf
TsDJ1xDzFAuyqNkk6Ylw2lgVmKwbD4Qa0w5EIXFsPfPyW3Siq2aT8P+wzHiBWITsQBmcj/JhbAjy
tA+ASgDWY2tU5wRspkPgllzwa5VQX5cAAjHc7sRa68e/uV8LaID/Cu00rTKbdW0HgSbAF6jDzCE7
s77fIVs67xPOc9UiNIdSWkkJQq61apaVsEeltHsQbSSUPvnJu1x3inZQvUKYmLVgF0pUfsGj9ldh
mvCAsw76RGBe1zK7jXqUiJ4h2shAdmRbIs+JlpHyXf5LSNRm4gzQl+tMXrZiMHJhtk+1FWzHjcIq
T682QcnGTquaRBSjWlxOoRM5QldGlHBKPI8FWYZE3ezdsfY9fVAAwjwDTLzTrfRj75iyCsdG61yO
wOAInuXZemBjAfXzyjfEXP/dxrgQ9EtIG2/sbB+JDxMeE14g/pHkq099ogJn7kqConEGG62WTsFY
IyYn+SdiClJtcpnS5gNlkcGX580h0kj+R4sKVUaLYG8znQlniHA8WnXyOibU+H+Ci2qkrI3ns1wc
JAZItjQepJyfsWy/VE9ZPCwIDTL+DIydg9PdiNBH3AixnefDji2Xr1YuTkMv2+/buXmjjp8HSC7p
/NPWvTaOGAK2ii0yQ/OtPbdOnbC5Si97MutkAzAPWUZUf434wP1UtR00AlFv5npBhbwOSqzOsDmV
ZDjdmbM2RuFdSleDX72KfiXngRp7jBNq9SzLBHr+6F+nCwxu38sxelBFgCKmdS5NZW6/z7HIrbwX
rQklQ+yj8BF8MyDCQUKzyeglYZvvwWlV0ko9ri17fMv48I22fvVgKG+n8AK120HVkbeGcE6istZt
0XZ/uvnHPG5JdAtkifiWCalpnHA/RDDu5yLR/QQG32ItYBjN7V326j320DrF6SQ2RvqgfvM1IPUV
EMDczUxeWe4Hw1sYJlCu4o05XPq2s40sDykMJASjPcqrb4KGt2X4Mxnrz9bm6RgRKNcau7X9MY8m
haVk1WiMWEwDyBp5vAxTUvRASnzGTDxedHK5/obbxlrpBJUnSaADp0q5+GytmycCfB9gz1lgkKbS
NoZAGUcYSfH/mQIazDngxYGirQSF6pOycU4NYU9KL/YuGBrDOBYzgDtg45lv/xdOUfaGpsMWBxPt
gjiCFhu0WrAnfcs08CtYGwR0PkOcstJ1vEwTkJWdv1aMU8ll5AKIEl3/+BvZpu2x9dqDKXHPGUxZ
1pa7lk4uJmut44T2C1n7FAhPnuFCW9N+0yiH7ClAvW+Ii59kRjhBocs0i9AfWFpixiCCemaypsg7
+LHfkgCDR7yjR6MO21iQgPMm8akiWmDhHD/Vor2WHwIKi+B/Fqzx5e/BqKJHmy4TvJXiC+/C458L
rBWnxHOVVdvQFi1Q9jLtGjDUgR6fA7tO1dZ68btpWXfHdCec7acoQDHer0uQQMnzdPFoePmsCnkC
c9fCl/+DIFlfKTZN3tjaAoR5I5SZWEqNjrtT/o4YHkgr44BjelNtGMcopPwjoibHL8T0jTdHgQcI
kxeoKv3oLbI64nYOiZ8x4Ah2RIDU2a9dU4G2Hcrd0z/aJxQIMzU8k8bIY+oOS/eptK9z2BHxYy/O
jPSDAxf3iN0BMeIbiiU/hsHEl6vz6Ms5mfCyArXWsQyWhA60YqfEuq8/tlU23SZse+KCqCVJksu8
c9ycJgY109T0p0jqqnUcFlcNUK8K3rr0igLcLSFRunVv8ZoesAYcxppdOHErYhgDnSEZA35V8Nmn
7RHMbKtIYwj/PoUBJVOzUtaODxuzikXujmz58l0nCHEZ9w86mCcwt6d0YhdsWtCHmBFLY/axQwcW
LD/nAKdwmoMnlfUqHUYjRSit+9A8IbGPHb+BGbo8sMlx87ge10MSgd3x6uKO4YBNOTwwseu9O0E3
yyDePckhyToqQdxx8cDz33Vb0wjJ8ziobNY79HdHQ+JXPHgdcEBl+mrd8C51/xpP+SSR0PCTLlsy
8x2LANa03zEmMPW4+AVyq3BQb/83WPIx3XfC0p1qPtKiSQHgl/cA0MF3fX3nRqOK6qzp+ZpR7EZT
2NQAFCYhsKGOTBVSgvfEfWX3Y1REezFdPE5hI6HGsRf4TzcQAY4yATdq+YRk1w6m0Yl1PkHq1dlu
B33eDtUUAXXti2a+J4EZ+7M2nj4dWEV8vIIYNT+/TRn+oJ+/1VVwLUMdvlz06BFz3yJJYseCWyu2
s4HAP2CUsJp8RFASPzEMM83WE5wS3fgaIqqBpb5WyAqHRdunDFgoV/V3DnIGrS3TNnVbJm8QB6gz
hGQEQoQlx1Wxzd6yCKMSiORM1zz6ibB0kbt3FKW8cWhxUmxhwXQI4Vo6JPI6gDt6UjkQ36Ff5o7V
8SWIfb6SQQmhJ8I1/BuxCx4B1+1kmChp230d8rlae0d5Z9c9z8o3kOCXAa+8w9OSSFnM7HpJQgnY
3Z1OuQPrA4jW5kUCmmpDx3nxEkg79YucvKP15WnlpOgUohvZrPt1kZnebSedDEwvYSWIC5k+418R
9X8W49eXGU1K5++kcQ6FsO+CkW5W/B54JfeIHai57wXWTHCOkHm69sXGg18PWg1JjdfVeE3Y6gfi
Yx4CumDLn+Pu1E2PvP4Id2QGT3UPw+bhYnLyiIQPhCbyAzwnkZ2QU6RuvJYacnf+bzJaY/KGcBsj
kxuhKT1Vj3vb3SKL0rjxIZgMCPqQhieLfGL0DyXbb/WTwAeKonhwuOTtgRsyzrINTVNLQ3quOTTk
hTGXb7abPGrxMUHK6Jrk3yA49JShAa0TWkuEbDg9LD/2YFfZPh6XCrGbyLJNHhd3ginsYNlOAAe4
C7IPXTOL90f+TkBVuwPNGl2nWg6NdkogLr8yVwtzpqJZuw3YMgSqm8OZN+zUZsSUd65vYo+fvek/
39PIOarAkNOZ3FJlxyC2A1kLPmNIgXJAQCbCgdIekJhbp/Z7jiPmpMJK9VX/oe9LLBq4FCQRM4jS
/qLdbUNv9Hg6teJ7XoBw24k6XCuztE0jjonutNfN4saGL6nLR/Dwpqn5b8/mzRO8hCHlyK9ghjdq
rZ3UcUD1x5MgSguZlrolyl0LBIpVdKr6gsnTCs815kg42aRRj4086rN8v6s4lssoUfmdGi2d6LUa
8cSkfJ0Y0lDh0xeR8foPfKUhPAjHiwp/DuWcYWojXLEB36DJNaX9gmZUvKEdvsmAZvRWqE5R5+OB
vPvOmYnH2kgzyKJ9mqIi2qbyZsKTiTrbqgVd+bRtT/9LtYbcX/VO1MueyNc7u+J0HuKvBOhwb9Wk
CSxtfRUI807LBVPTXbwa7uBI3+A5VN2A8mDwqNxpxKEamYO5Pa1HO3G1H9EcDCR9yLjeDCdLojJi
8tFRYiPryQC1bYO4tZVE3CffiARG6wlOqmZjX1z5zy8dNjMJ2wvdojDtMAwL3+in1RNtb5ZWwHSp
vybgyf4G7RtknhBx9g9yHJGUTExk2aBqpisLD65Mcn1s9EJc3TsOWQGzpNr0MFoFkfD5038z5TWe
OWHWn+V1+/zPzsGTyE0taQR6/53nQBU48EBz2/URGjTr8oCn6nToYLEvz+5AxxwHEB68Yq5eMekO
yhIC4XFX5GXOsZHm8d5UMaS2KCWIvpm1aSUQI+0fo8LAS/aOwKQcrH1n7cNGoSlCaQYiyw5Cx6AW
6jIed05L6GrwCOCcy53gmyHjyE72IhR+DjYjcMoEUhQyVBRzjm/nQoUZTVLUTrFSvfmKNyGrmdNA
hiBfaUJ7v32Jw7w+uPcYmb3lPecXZbLuynpSl3hxWaxGd8ZxYwF+yhAPJBki2ENpJ4oRrFqJBgPA
sWNSPSEhTxABvM6J3/NS7UiUs1qVrfksuxu8xcJG0mLDPn5Trhpp7BIo9MtG026JtZrPZZfPfNh/
MJ31av8uUfP7arernRJxyMtattm6AaghiIYhBaCDI9hOleGPyE5bmEBBvNgQnpKw2Ff91TQBa+D9
YIQlVnL7rArNSNKPgxHpCTisZnRX42URMq5lDr/Bz3KDsVyKObyTf+zN5+eMzL0OHqCgVuwDP+xI
sDljEBhNqDZv6oup9DCvN8ewIJkRLl3cAvs5eVK11JZrOvYhwJv1TdM3cWKUcs7jeMGTu9T9VCUa
8caH0y1p9WDbsjQ+9SlM8fmTkZjtKE1WPgX/h7jIqNm/RIHzR7FjUOINTZ96pTumOrHmFPjHpf7G
jau5gF9b3IJzzLAoiG2lOpAo8DL9YuABLJpq69sLVL5Aeg9x047uqmmGcluj2D4fxfzybgXiTIL0
B4v5lBX4+NW3W9rfNjNrhExzu7PvqTeT3w6Ma4YE/H5qpX0WV1IcXmesSK3nPO78C16gjHIBQgMf
7AINTQLOOaUqvONrk0M3L43WZZPN5tET1ufMH3W1vw5HH87vui/8qMtjmu0ffoaUIW/DfHVb7sHK
cCwDmN5KKdtKM8hS2GvCOSduNzxHjwI4qoAGcIX82FqiVMkutIDQKrgqxRjfAOAF4FCUMhhav17y
Col/OlcYOR9eucn+9Ux+4WrVlJdZsOwNKJ/ZZNTQQEUR9mXlc8BgNhk6WnRi5i3+Ynz/sbG13rHy
0uqlMj/n6gyg6+zekxVcujVprxcgqPanlrga2S8kYmjowLVwv3soL7HWcjyf/vkFW0bEN57R2wve
NTCzXgtyI4r/0eBt1wWhDehIhNSKH1OKkekxASq/VIldokuyg2OuJhFRP8skHqHKd0NYhaK5JSng
RWufB9I7+TqPDKk8gKjF7oe2iVYICYrL/TRAYZMBsnItOFuw80jGEklmFMCUMEbqCKUycGzli/4K
B/tl3iez7pjhnlK5IPNoCujBm97aroGKEDphEmDY0cKJ1eaxDhU52GlcvIc8VUaWEnTz7IMcB1N8
Ohtd3oIUNZaLkFGeNf9Qy08jhpKt37CJAuuyHh1FKUVan7/IGA3YhVkn3G+e+KszDR2R+Qznmvtr
1tNDqW42p6LdVG+1Nh2boae1oB5UyfqdkFbbiKkag8Jn9U5H0LoDa2QOj6C0TX5XGJQ7w1jRV72s
b+c2OFsX1cKNil3pzcmFxWQmOyShLjOSMFXsb10ph2qTSJotlSmF7CnKwpOvuUfcEjnv4K9nRNzV
L5m+AN8lpwBkrjnc77RR51xXQv6x+EtR4k6CUyfIehkOrgLfwZZDVtRm5IOjnHbxki1vLu+dGdHO
XUcZYFauJc4QFCzbAbHpTSPEpPwLd4emwhHe/l4wVUSt/o9MqxiXYhAOFM5a/7+NnXsLIYHWacKn
X76NQzl+ZZmcpxSmn3hxgXIomzcPfR5hia9suhN5Xw5oaJwN6SH91WXn9GpPkTqvc2XR5a5IkKut
MW7jJ5F9HJm7Kx+mFMFIWxjzb1RJFQxVbxcqETqctc5y6n8tyx+qWFlHwUng7o6ibMrataJKbVP2
oyjZkPypt8X6JW2JCsW9Q6camLm/agdR1BWmv78HIwMe5+2YhehcTY9y98kP6fdfmuoa11bzy6wX
syef3+1qOuwTRnBKPXb0GW7s77kSLBsHTD1BAlMKnSDDnWARxYqhnJXPHXFPQe7avG3lmRM8OmfP
tS5lz/C5Wip7U3YvNouGcx+LMrj1iWT/ZEaNID8wLgVu7wIHfa3fSI9weV5bXtvu4r39saYIg6b1
h1rfqPAZG1f+11kJs8iXxMbrfH4zHH1YsbTSXRmaB0reX1EXGV+7M80fUvsuACOz8HRVZvar4Nm3
5CugH/vm9evjwSwIZv/u5oLDWOof4lnLeM8piTHP60rZQY1U81fEE4JeGrwRIYVu2vFYvCoYWURY
WhStE+1DWsazHqFRjVZGsHlq3JeCpUP8z5EJahm1WFVcZ8p1jO+pAN2/B0MZl34JBz0gu2pQdtal
79BmDD527Jw7t0xzgWAsl2D9X+4Lf3As3bbYtooNzCud1owv4p/EScDGyS+pWy/0RwNQibXtozoK
yCp346XF6vijGOswlEhul7IoDUbyjgu3nyKKKFUpSqjGoogxKOnhdsuCKnGBxW6+Ga71PA/9C6Qx
XMfQ5OgoRnmYxnxUzlkR+6tkZwLYx4bkVI3c7Zmp2UeKTJFAH5mVqRmm1LJyFKjTqkrpJMurUmbu
oLL0SycQ8unLbpV0lrjGABVnODShvAeY2J6anYwX34UxNF0HHnJ4Bbrn2//HJv4cWjTkuk5AmDd5
3W2OPXUL+LzcB+pMQZ+PRNJ6ItQkZWRrUVJct5nynZssfg6J8jxmsZ8F2yeeJk9hNtPLd3P1Gwd2
NPhhEPMn6TbRoupuzFy9wHGEo7QlbAWE+K9ej7/Dz/JLCQQWk05MzhfBnujbe3DxU2mFyfHXE4lL
PSPGfR66nS3y0u24N2lv0vKxYVq2J3YGz59+ioFZQR1RK9Iy2n7r8nCribHIppzwhajczkRIUxLT
muLfj6greb6ZcWRyX06x/zgwaZCrPE9rBt9Me6h4/doW4Qm74zi0q5XH7VzJddNgoTCREFQe8NDt
atjwA+lq6E3609D6irWkiGP0qLlDeMJizX4CVOB1W/FadABEYEsdN811wjs4PTcXUkQ4PZKxBSXG
1vqNYLTRIvLp+GQ1A0kQ5W1WmblYbk04XnN4BOH0bZlZEMcrpDEqy9Sj5w3LIGyEW+dt5adakf1U
6vpxUdat60YZXLXYMs10qvccpwwp1JuUJedqsjyrAsa29LDXzsCnkaY9BlpDM1gFPARhB7cz15td
691nVavjuEAaS7uru806VdBC88kArbp9YRRxjgD5TlM5pc+hnF4exNHViHNCWr7+BawXXv8mMmPG
O4MQtxss84vAEgHxXVGqe/tqE7wZNRhEEV1KrNk+lTV4iJdWAbvvwV5JzOpCvhZGUVEBEv2HsMgG
u0p/zCktRgan9FlqbgXLC/mz4mTEm7SWgMjlNhDo9PC0qGJ51kfXmFoYjAh26MhyeL2BqUn3iOqn
u3yzVWQ7LYJY/BxNORPC7pPhadfgVbgoBSXC0hy3SZ7vB7/S3xV1ypuPxb8VpZdKUuzHrn0jAkVX
4myRgqXxpmLa2+/d9Z2FinNxaYOyIt9awIOtmL3MR1aSWyKLMIaK58pq/uTiiLaxzyKvYoiYvIeM
icvd8hukuNwtTbyNfzjDbUjwjKntbGa46IZ8d4SdlmURgHRhe2CquYayxP2eFMysJ/WsjEv/gwAS
qowojDW72GbqRLHe5suLObx24/el/qIWZPpm5bqGk4DnwBXaHtAEVK1hL/VcYUWlfsorEyrv+cOZ
Te/Pc6S6MTMZ1m7gwFGZjbVltsbRnXCmfyYC3oVSBZQzuW736qJruT2VeF++9s8vNVBe7b2qvOLG
2W9PzYaBtYSxuZzQlYzTcDxB+v87L7Fp13+mnmHS/ZJStxNbYJaHk+rwcjiILjwopwo3GeK2292b
dkU87SiXgTIGvi9csDUAPQoxU4m3kZOvfI4UPR1RsHEU/ipPmEVQ3xrxj2zj/HOoariOEvq8xEOv
CMjQ+SJkBOrxfWDdZki7aBL7B9oF6nUfPFL64firoaXtR62anf4SrmySWGV4VPPtUc7+DWUqY+bR
RKmb+GiWmUZGYH6FVQyDkv1ld4dN3yWzLuoGi9EycnQjAIywiXdLUlHVqlLfCGoyX8bWqIyDct9O
d3s7xZnyZio+1/MJxXAYbKo1AU1DatTaUG4btSEfPS9+cyH6d6IM6ysF5xHFtw9Rq7LyO6b9B17N
4AEY+ODIaFPD51JBXtROHiUknlo1PTohjTuUZig8UADljw3GYK5Yx16I1nNYoR4Kk+T76VxcqBHH
puKMomc+i6sduub8A3p0/t0WFYQTFbEqJFpw9RyV56fTgAg1349qxTgT8wtJM+GCnNscmnK0nnjO
iNzwo394gQApWFsu2X8b3lP2l7fCu17BHhBfcVZom49vauJOjZHplg94b2HU6a1vz2RR/wfv8xeb
APq6T8crcgAzi3w0AUOEwjwl+DWedAxpwsOMAg0zVc24uW0GfzjYuoYUY6sOV+XjYn11IVS0NPkd
2eWzswS9ng5HM84lK8zHEOugE3njm4tbtG3reeuxg0tzWWKfmRES2L8edAEgI7y9abxcKb5+Ir32
rHdtj5yNYLJKOtwrWqut9bgVfLZYIVmSrAqp4Jn4a32hfWlu16Kfvds5cjV+t2xxyXGVfsu+kKaz
I67Nl7q55WBU/vllIYGwUkt0eki5vV0R8DlkLNV83Dhsej9aGn+wk8wMRowT+Lc5pneJGEdt0p5V
C9k9H7C5x2zFcNzbzlNGViJDJinGQVf3P1PRZgUwtiuPRhQkodgEzxjLNCTYat96AzNt9JmBEwOU
S3yjeLv1nxHaWezlPP9KbadhgUSO7/mZkNAj12fWfNJ2U5LtoSNWngArgiEolfjehCDW0l/LUq6M
gaP+zukmC2JPh/NxhY9dOmPf/sfnRmFF9lpUlrWMF0VLGYKfpYkpkd7M4VLzaa2QaGVhcGxKkljB
+0HmhrxObxtvMlMfPzThndrDyEX2jnNJTlpqKuilvEAUj4LcY0y7Ao36Zujv4RL0PcGl/x6cYIKk
f4pEsweEYgkuTdJbWXICVGigdsVAm+TEoWqTu9eSohDtGhjO7AOjoQ4XxxBO8GsNvUxTkUmT1M1z
lDQrvSNDnVHE371/hG/wNMfIhUqeZyGhB/pF5ndmXWtvohdeZHySIEt0rNxA5e1OCKoqbJT6j7fP
SlLU09YysqFVMcyE2NbKlFADPMCzNprW9mjfkzkIAD+IXqrMhAtqDIw1ivedQGvgNcDJwhr7IqwD
iWCBEH1TWN4MkaygOY0kDYxoZNO1lNrlsMEbidArAIhyFuZTZzL61NPP3jCr+eP1TeMANjjvtkXN
/meI8ArHXbohe6gkDSikog3Kf4UOOELs/qaeQvMBzf8WswbjM9Dg17NHUJPi4JEnN6VmueUumsYI
XpKkZ8/Bpbv6CEiqxwULs7ViH1jl9uV9CLWuUlOqR/S1AJcKGzbgycshsmL9+1akhwA4MhEWRKLj
c/2+qhy0EkzjdojZNi+xR3PrqsW1tMe3iVFzls11G1HIR6KkrNhkafD3yjT4GO5mROE6Kuk+S2gn
Ci2QKkRGej4jOevY2EAFc/gkjApth+QbmVyFrj1SMl18KSciOMe4/Id8kK+a152Wdjtt++KELIx6
HYXsCUa0H1uHBnGq7EH0Waumc+2f6xq1CuSw3kirgAhPVg2T9gTX0EWfEjY25s81q7WpObnBkWVb
MZdwLTiOXxckT3fu2TZbvApXJpGixP+tLG2s1bSpvt3r9Mmzc1uDYYrnw07MIgJd7E+k8B7GEg4w
dk7VZuTXj98RPF5pnG3gl2jCUARtTs38qMLjWz3kcepNY6d8Kl2YHaFfwHY5O/ckwD5PjoxBIkXS
SVfDwSA4NvKcLpKOjDP1ylmjr4gv9FYwG2L8zPpcIxNHd6kplp95TjY+UByHexfAfxYRpmN54APy
HdZ5fQaNFXhF4UGs0pUrMBtTi2nKz7qcj8tRGMAFlzS0Uffoff/UnePe6ZkbjK0lFzCSjzzapFVX
Uzk+HWjRpJa9PGRfQ9XnqSPCEuzSaqosH58L0ASD0opdYSioNf011HuNGDL2JjwKsqy3YxUvdl4P
VxHlU7SQxGdtxtpDqbhbMHMnZhA9i8ePxpLyfrN1C014rVOvJDocUKkUWSg9p3eYAAouLJFzZ2V0
UQ+6FY81e2CMKFSOm5QzLg1lPfaIfD+EtKiFLM029AZ1uzQIQF+9lQPEOu1ddmC6ekOHIfFcNgzk
rJ6dIo9kVTQZO/bjwPjWKUari27NTSrOhJ4d6nIR4m7Gya+gk2IDUZeliReimoM84nD/AGNbURzy
aI5/S0TOyDI8IRd9Puc89pBQ32IQDLo2y3H3Qnvir5+kyfIQqpyk6VSViLVntrP9wS42qjz3+cnh
Rr6lsTZBGaWy65aq8oCYE5eq30pHKjEvgHxUP3GaFJQPpCAcNuDuI255xZ3dwTtvx4VxKYsH0FfB
Vbe4OTG1zImwK276GhgqoWyni71s/9P57gFA5ZZ2pcvRrJor6kX/IOwDkY8wqBJtbx8J4ybXu5qY
aIlcTxl8ugGlxTW891bH6EAjKq9JjnG2z0z4h+pxIEwk8brApQNK0voktAP4hYakcqpxaCu4lu85
KkPG6a1ukcVmvyajmm0CQcTEQNblvwhxHnLZVZ6P/vg1gALmxcZ2IByuMZln7Uv8Rouffiayj9uD
VhQRZycXYjv+o2RR+lBPHOZ/PkkTNOuFmBKPxTI6ozCDp0S5Pf0mlfyLHJCtXNWfjzIt8aIw1zHt
uovvQpruEvDtUq4mNrwMlIaceDaoWTlA0zp3krcFx7Ig4Im64sqYjdSg6TrroVRcAYtU0ztB6LxW
Fb6/5CwgSF2LxQQLHEQtOuHfwkDl0iasfFwjUGANtVFsS/1VFUO5M7+17VBgvIQbKTy51F166vJd
p9hGggDB7c+lOxiZsZ2U54Lvg6TYd1utYBPW8sdB1I/u1y6j5bK8W0TmDGuB2fCZSACvbyd4WoEF
vbeo48xPnS625ok3ip9cG3tOBkumsVu2hkMtFYXGCWWA4MHolVGtD7CHR5J5XUiqsHJG2GeRvMI+
Ek834RHDDxJkbG1TyGfvPAPIHK0csT1vPkF4ClLNN7j9gVY8oo2KwwSJwvywOvf/aNDuNh5r25up
0YrchVSBJ7ZgOVk4yz0H9S58kIVjJOenBCN8f4PIBq9b33ZHvcJ0Ta8NWqx5EHGi4U/3FeKnc8it
qdAwNemaGA+0pCa/YYxsoszbtvnztwhGzpMeoZbwxQLQLyCTYVgF87ZrIOmWdVp38UBzZIbgaTuh
vxAToFaN27D+guf9Oar6a0qR8qpl0a3qDxKUy8P2+lnG06vcSoN8Oa8L1CrKhME5JXg1uGsCpYME
XCW4ytjXnr04uerRpvpLe5s03KzHq9hseU9QqdC2bBbpfa/QsmFKndQABqieFVfsk5tumDq1trF5
95OnGjm+kNtliyF5EWwHL4DoM+zXk+h4tdeU29v8MTf6OpirqP7N/Uqga7bntIvfteS00CiUSgKz
rxh3q3vEzxXhSRqz9Y+Wurj2HeRsbLXjbwkPSIbXYoPYICF+5yNyYW8IsAYd4etdIsGT6hDLtl9/
ko+vdj8ba4Cyj0CGvS33db9RM3PKQcNZ9M/Cj7y+blZQteHFZODCd09b0iChWzVcBW0xqTqdZj+8
43dCUxPgBaN/TrouXFQs0cP2zK0QAjcXjcR5JSO3gClg5MvU+EPJRvARMBLTInNOqpVqBQ+9CKhC
1tgpEOFCExF468/JsazpKSTknvfJEek7CThtAHoyX3wzV/gYSIrBPWHVGiHVZrwSDYjUFYLYL0/i
zVlw5AJqeHzVPl33ukN2/cSYc5LILPHBGcy0hGBjiMilrEm/cjwJsGwEzZzM3QuouGrmVpLlQ5yH
pgUs5POT86kX68v/V6vFo9quuFWfEOdPGzLBc0k6YobfZLhF0pEJWyKbNesDwEsrcnOPlKN6iZiN
ilvoXPmWcXtS5ytnHruJyHNX5xEtP8GV/k8brR5O1tUH9RnD46m06mXiJaCVxMKW8k676Q+Ar+/0
muFyqydr1UZlGWrOOp8qY7ZuJOCIU7ysbxr0eCl3ffxv133+DqVceiSkUtpO01ca8xGoobSHwbZG
+9S5bAQgz8Lq3gnUahFrInNqFMM5ibnA/6aUBo8AsdvJD6e9ngshaLjpYv9P3JTN1JuLSsCxp6mA
RMpZA01RjdEjUy9BHv6FQJJEUm8SOYqI+8SH6M9xH4B6esG8ii9sczdC9EGxSmuuQjRvIGHuILD8
itTf6q0yFnsCXF/3emshT6fBRtqgQtZWatVpT/FfOxYNNkxipe7Or06FSkuY4WPc9Bvu1dOXBdND
32Uyaolw/QO4ykJOjJqfiVZlzgnrwaYi5qagvREyTWn9iZKDvaU8BScqHGG8VpOAlZGyj0U7HgqQ
571iUnJy6FkKwCWieCfuVh9cltRKKI+Lhjx+2Ng73WNWz/bFtcnAWUlvN73AbS943wKFV/GLd6zc
7whx+YUKG8QGeQHDNXh3G3T9SMIld3QfK3MXWjoFQzQwPtIFAet0w/ix/mym4kI9GBMXBz8QVGqo
t/Im8XmH1bb03/U9Hh48cInj9gVKD0OuX+YvetiyT/nlRpUlphFyxbJAYZtkOPeCYrfOV8Cnv8Cn
i6308dclK/gMbgPS4+p0XgKxsHHMsWBozj50gxZKLrSyRlXeM7mCDDjztuTqeijGbjumbSBEhAhr
xLpBKv/sFh+mgcMB0sOdf4v5RzMhC6XMA0z3iff/i+NwUvG6afa3yLvcRW+FBWcpG7C72UpNeuZk
jTfdHZC6FYc+53tcO1SHoMDVxYjOq241Sxdez1hziHE8LzyXfyyYVQZedMC3nkNxTx7iTRHhRwsN
coxCZfdtV2LygFrDxdKX4u6dl8BWtrjPE3IenuUd68eO5X97sjUgEWjMk57NZyfSJVDAE4iznQW5
cUh2Kr6arFuKuq+mm85Ci/bP4tJqgaGxVsDrrgEibYywu/Am0MH644LQSN8Zn96sHl+TodBRm7Jk
/1agBFU9dGcgvDQ07NqurzKyzJkXjmVko25GLCsygkQkI+41irnTxcdtIa4E+WBG/Kchqwg2cuLR
vfRrY7KzGhTRM8UwnrR0ZF61Dtko0RPiFaFbVV8gUp8X83ZUU+OROvnAj6Aiuz/FUGkiV+ayxA5z
OUOaPDJleeEEEoAm6xIxynrJ1gsrGnhHV0MVv9JNnm7qYpYrGIU6uKoFDH1wW+OzyqD7gZTqFTVu
RjjDvsh9FY2aAuKFAi0y842jILZkgti1HeSFFu85c7TGIWL3UJCjAUeljnQFievwkCAsQvlSfhtZ
BTDh4nlOi1OwUaKCwBc+ESrqTAImFdcsjCt4/1pIQw20BL5bXPOBkUIlZmL+QedqMcCJ8yiHEPPQ
Mg7TW2YZaBW2JjzqgS5XUQU4ef7GGTi2EU0cLcj850ErwiLAQ188dOEIiQxCvS4R9wWpjlutk8Zp
OcVnj4YXYQjxksdNAm6yLzzg0bGHJLv3+kZIoSWePNQ/hNSe60i0nrKT6414aHyVX3TbfkJ02N9W
zwmpUlZHmBkXcFFfxBoflTTOY6GuxxNzmeYM3DbhvW7eT+gzacQu8eWxCJdYMxuogqMg3g72OJKS
LEyB9wckv3n44DUFyYLG0liIQGtf7Sb4cOZCsTUtDgL3LQWuRca8WrCVNUGK4/zjLkR0O4qivpMJ
p99m74Zx/hPsG9zRZJKidYEtpEx4qiVTU9F7cOIN7bmGu6Ju/Ce3Ydu7UNgzkJuka0ySVfvjb4uO
Gq+zcGdPRAT8QgYiMaZda/V/vRpX+UJOkToYqJ9yQ85ZMDL2517bwxQ9QRb/nGMAX+WrQr3C/N6l
XrNsrftmRl1xq2hR8L89NTQGaMWNxr4nBaEKi4rnKbyVyfaKfqC+9p281sbBF4f99kQL4VD4fG4G
t6qqrovy1rcQB3hQcfk7iHjw/UMgSWPVNqoHcPKkzgZa+y3812JuVa9mFedQZy9p3akVrhga1mKY
EWxxc5mbqUExK0cNX5k67T7wpkGloweB1/5pVefQSQK60lEFY93QWrO8fkT+/jI9XNQXho/QzO9d
ABXakHCwcHIpkkOrj4JwhutBk7G+zt6wySzVaS5DNc6w5ShnzGj9ioLSQ4BxW9IyhleIpTcA4r+L
bauM4ZAMtKkS9mMtlP9Iim/Bz/1vYi+x5Kp6MXl6AYgzx5llI6yoJOU8HetbYFFuw9fG5WpTKQ8k
kYJtwRogJp1AOojG6z9cTFbCLSNhi680lmRU8h6cHdvIytqCszHw7onJ4QMiUQYhhqQC7ixt2nVZ
Hyr+8CnXcyL4c58wsuSqFi6XjV7NT+LiOqPEiu5GKvFMXz9YiP7bUX8EGQXeU122XpwustIkJi7h
XQeIxNXQR+erLH5A1Hd3Fgtz2DrNbW0ErvLzk7ajT3XrJZ6qxNhJlco6pPEn/xtfqbU6HWBNFArW
PUymtrXfwR0zRFra9b2Ev8tpmz00CPFFQhWSScxkHLr/FjUxdoqsrfbrF7//w0/A9MD7gFUkOy1e
BFGUGcY7d7AUBkTP2ynFixQug9lzGBxiNc2Q83EKGXG6W4zC9HgRGiOuQGHilSsImpPgFJLvgU3+
YGOMiKvDcVTTeBT/kKT/Ra/z3ZcDL14pRZSr2ELOYPXxZ1MfoR5NlCrdpyCbpYYg2J2Qr+Qas2Bu
/UJRo/mp/+mg1c5tUP64SiWmL2wCk+pJ/EfzIBhHC5gZkDxz+9rX9AQpzW4OWViee+5Nd2mLF4/E
Of/E20dcBe8GQdDypg37UrV/8JiS0jclnSa3dojCl+QDvIMX/dm+Yl15UM1mLOgDEUNUGG49Do6a
MqvW6u62rIkM10HHM5Mqw+7Cxe8wz4fM7sB1Rk0f/LLi9p5MxB++60ptQrz20in8+EhwCkGwtIaw
d2+omLs8BFqmScAhEx07W1EEmWzagHb2DNCqgnmK3UohdC5HKGG/jCmEpECs9nZDpxhxTec9ictd
BDyVD3AUegEOLcahO5Vn6CvC0i0ixzfGZvAee5D/obL/lm8FU2Kj8EIyR6D8c9z2lJne9vBY0bNO
sIBaX1VR3kgnOPCVA69btbfMxm1bkupGLBhke1BfrjNry1N7HxiQxDdKw56l3EIcjo6mbMJhxfQr
NWEljfatq0P0DaxbnkEoA99UfH3O9REy6aeRn/hySTU3au/4xF91Ga8KeQAO6ZIUW0VEMSnGR68J
5rDwimea1RkKOZQM460uI0/KrDG96RIOYv9Szk3Z+GsaC8iiAszo1mBIhVNWXJVLl4+F0hcBCrAq
m8U7ITHr/Hw5dOtz1DTW8ZQZ2xb1Z1DEpmFzhQmW1uHvO8NTYbBPSnHjC1ynC+0gam+0ePLtfXZq
AhJ9a9ScgoMffa/KWk48Ous4o9UGFaFS436TAk8K2chRsiNRuYWk9dad+egpymmwp3lAQSa2o9R5
jwWbq7XpCw8wYrfPneUhrJ17n/iUSCoBobtOjwa1nAleCJg8eMFmvgD/CUYtXk9jZgv2ll83w0Kz
fcDy09/tBr6/qLfmQ6nawm8tjDC0+L6u7AsqQuaFuRDGMnU1I8tEWwetCIOJb1AMQpdhfpT8hZrL
Nw2LS2lehBMwi9qMqautce8OICDzsQxbbkpDI7MrnzuhH6wcafNXMdBmwODz5vs1u2GNWUDfpp/t
I6IgkOkLaM0j6hq+c0rS1kCe5uJTjF3kit4af70V3ORORruF1c26L52sVQCYYFCMZvnDS4yWS+fM
HdGokIbTn60T5/9wWfT7sAMinlhMrspsUjwMH3MDqQyRujAsXsGxjZUMwTYnzYf94Gkc/LnFWBCL
vESCNrCpnnhJUY1/BJMqP9k/kASZIKGn6MGTw/tb/96drY/sfZVmUTBuAKWAlGuNwRCsEGTnlwld
JL0f7I2MG2lXoNNRvs0EhoEyy6bjUG5rrUcMj49qiuxa05fQbAWSd8CGVVyJb93O/2j5os4mGHF4
7kjUsvmHjad9G3M87PHWX5QnHj8j4mCX70TV+ir8tXGZatYrqoXV0fesPc/zNSsj8nPZw+F0oLKv
zPOd9YH26xkWT5v1brbD14f1wSX5GdoY9NDhRCLsxFy8btH31A2+vSUxkXpe/g++HR7rAJHBxwP1
JPUGvETRGfnrJoLzmqrUv5XvEUzp+BiUS+UYmJ0XZRHfXZoa75+3k9qLOqGiQ6uKRRIThslVOylS
x5TnF5oNrGJdzGL73XdcI9RQyrrxe7NOWn0L/Kc6WEUWlXRMO/3UH9Jehs/rLkvu6sq9CH763u01
0WevRLN2OWlhHobeoeKkjh8QLwnWD4b8ct9jNaDL3pFy3RrJGWuQo47KlbA6QwjJkMfEQ9dftfKV
SBYdQzgIgiLFbfTqiGvp20sQ+WwLov7gRfaCIgApenHtUNao86qnEQv7VYm0NjETPAkjaqZ5jZec
JdTboRthPJgdZWmGMsyN7L0ssITvFnGnnUdM5sR7PoaHGb67jHjVvpI+NKDitAUTBHKecOrVRVF3
3dsb5P1A6YnXR1AAIeh/NbrtS+Rjms55WByWVSH+QLVxiF954chCHNb0MhZ/k3pa9P7RqaCO0Lej
dNAtW3IqbIjSm3pEeckKxE5ms6EQ62OYU6we/J46NtZ6eYfSjZ3QTLjU1ZHzvqPae/ZBBrai63dv
eXFfMLAGXEWy0v9I0lOQYrpUbyPk1RcO39iL6t3epnoZxo1VOYZck++bx5g3dlVJ+KvqxJnvsnaA
Elj6MYVHNVNncJxEj54mdIOFpw9F1yYhRTzT4j5NWLvFtVecnfzYCVFu9s3wBx4aPRPDjwchI8cC
GcI1f7IVYKQRD1LZWRwTXwQJBKzLb3kghHTUB/javL0Vmh9HE+Z0L1iXhcmTdgkEzDG9RA2oytM5
on9ZhUuHfOjAChHALA6rDBziDLAWFQThu/AC1OpT/+AA5K41g1+v2qCXMZoc8EId2cbbvcPIfw6f
r6inqWFxAg5R16N/9OjJbudSjgrHw+aEQjAj1GqtRdf36SGAfGlyAWpVYfkGiO+25oEuqnOpHND/
sVhBkiWo2WpMfydeyXMjGioa9acqTpVAlzgSCyEiRMy87IptOMLgaNskEAvEZsjehNIHWSag10Gx
m0FiDO9YP0IxqsziSvY7eDUxeU3/rjw86U3g7rrPJeWFzOqL/fExpmvuz6X/0RoP46OEqIg+5NyL
4zjgeLikjkU5RkQ6VnrIvE5Dbr1jUehvzBcQJTjjPHD7eY9vWegu7z/2iQnUv/eOtFP6TxqZ1wrH
DfTJCm1qPEtz7cviWtLwVMdhwslxJh4FUWQhJ1kN2RWF6sggF2oW3wMSPPt/jYVT7v/5boKmUvnu
AuZK8a4X+EafqCH69mZff0OqmeEb1vhw67bqMMZtp3u04i+u69Two+yz/Pf1HTqNmEfFk5qRR3Wm
MjNdcQdi9+1TbqU5EaRSbFgD2ykDPw0Lq/1Irx0vqhevtK+kPTsLw9L5mBLfapW/WlvMjwAVrN05
74dNtkMHuyCL+4G9ARp1C4q9d3KsG1ZlWGpDKAdr9uQOpDE8PvY5/DebDIP9Yh+/bHzbQLdyBW/A
EfNfLHfzm8ynwlyk0MWDrWEPvGgID1T3FSgepmM+dnBWS3FAgw7eXfspVZRJGCyOkVj7KAh7v9wP
/HGZKrWaEdeYnwxtGD+FutzDpcIujtBYqhRhVM/NvHnoL/OWJQteDJI+qA8/B+VhLRqIqh3s4GsY
SWgiOkcTbylHTZ/+Afg2F7mn1nKM1cV2apzRYAJvc9VadbDy+Y9QBxJTT+qQpp9w6ETXJAgIhv/m
c/H6inVQNSYqm9U4xGwnpQYKmwJOATsjgdGvMhDOsc4CmwLVtYxGkKh8K1J43CAKz+KvkyHMA7SZ
9lQM62frEA2xjG5gFdERPTIxv5p3e4eG3l453V+Nfdat8orZEjiQSAAu4Id/xaxh9M5vJTPjCxJv
R64Do1mCiEaZBnENvp/7iU0HwY0LiDJENDZC+d9KEZTm7L3M9xKsIy6oX1rS+EyXBDqlHl9mV2BT
Y9dM037PHJTKDZS7QZRUc0zWCZG7V1zYIiVBXp87/fqNc1ltYDPRCD0zUWLnrKTtqJTB+7OuPsog
GymU/XJTVMMFYTtB3AQYPql5mC+vInr47VU29GHgKVUmdYAtjxE7ckz5t21SHkrirv7pgSCve9QR
86KAbbqSTJ7ensyxP9o3AWIlrRkbLy/kjGfJqYGyaNjGzj2r2yFICTy0zyJUWZ7YWOnoInk6UDDb
y2UXeLFfRV9FqDIKbYczENXYMj6fYHwW974OkQ4IDGSEXDo4twmnjZjUBY2SyKVzdN8uDjPL8pNT
JCsNKJIEsqyicYo65Gkh5k72QdlsXCp8uo2nfzYIWjopt89WKmnqCcvU6I7+6hzRm5Zgjn/ZH1vT
KNcDcJC7JL6Zy6x9qQ8sQ4CSeHsAme7gBYNFiR7RShIEcQc3lWeAiRtaY8HlSPTELFzO7sbUiAtE
FetcvOg18HGg/+V65D9npKmJDqFA2CjV2X8T8sZilY96mTTGku1vr+iKuNs7IEqhdNb3/6PFkdM/
MTdzqklo8u2vvINBoenPkfRneWRjn7lfaL07kpBt3Uar+L72eOarsjDgE5WPQwW+YIPd45DnMGxE
OjDEpkkzRl6hKghI66udVDcLooUlYacL8TpQoyzqlPfvCJk1U6USQr1Zxu3e3m9QPlOIoXiohSwD
NSb5bt5dj4c5yYw9J4uptwIJQtxPrIIB2RIcyMFHQIOBthWQ7G0BoyenZI1FEg5pDJuIbsBXWc9+
yVOOWkevcrhozJjLe3kz1OIUNpWQ9cudrvGdlTJvquEg0TQdHkxHZ/l1BehtXlLyEsdLsICa/qqS
xtRATkbh4iBqBRcCJgiiCqxAxI6eSJUIbJ+QcBN/vYCoW56+X8Ht4YIwMGpsuRjuEkoTJTlS+Obv
YelQLMGZvIDTjVs/J4+2ghzfOjA8hXTf7GMx5z04ef45BtDP4/aZZOehuui5wCmzuQMJNHhsvy4F
192WID047BqTJjwBwpjgneuTdUc+miP//5J28letAMq7dYOUofcvkn3giUoHSaMx6EgrYKAEK2xs
AhH+vtF2k0RyGnmHglPTeYT1UKEGW07Q026KGXMMgjgh7yytz05605Ttx5uF5yoGkGWtC+PVTMfU
G2/k1wvsanLN2cL6YvAeHQxOyxJUzILJhx+aKtkm4f7Av6kd+zO50UPfc4UBwnsb2eo70z3WyXwy
RpUuh6wmMu6YH4+XtAqkai8mprR6aHxvFOPqihWBBmLko2EVoUUtJlBKsl4rSAZ8AbS4AjEeB+w+
NLlf3cuKg/NLGV+r8JcNsIAacY22GsnVMTiaH4IcWSsz1uiqDf92ySs/2cTdlpkZgag+I4ehfG8v
rPW3HVDO5V8Z/Vs7/799/eiMzybM3PTxmjnBnn7mBq/j+5VIkMwjytzUDmk3tF9Pjxu6bxX0NwdV
tldkAtFH58pyE1bZ5N6JHv1eglrTP2u1hOMGfGNmxmzBUzg7vPsmC+JwvVzJOPDDTPFNRUowWarB
p0TfRfK07a4p66VYsoI45cr8AOloDA13M+1NW9K1QkuiTkQunR+oEc2GZ92xeOJ6NOLhO0aenu3v
hMyfFk1yDrNArFmXgx1qQ/e5/+EdZ3iKfXacRw8XlIx6gZVSwopRlVHWkJGPzTC/F89m8lfOHb7g
z6wXaNYlK4K7vp+bOmJOmT8kf16WKTKzLB3QM69cad37wRgtDrlO717G2muYyvAvqe1NrsygSFyF
UILFufYtSA3aw7PGwaJ+Kv6kM5+wIoQsIaG+K1iZwN+USbip1occdzFRS7m67YYCp2WHynNnaoZZ
oNAxj2dLRsGgcJugt26z7WjuCYakkfJ6lZFhpFigQPrR2l6yira8N4ExHP24zRhM4xdbtmZiaVjg
LCYSrIX38OFofGHHi/ngdMb+wMGhgWcE1mwj+X7GaJNEPKu5DjhSxFwSSfm7j3nWWUgT8J8Y3QOX
L/U6G8oj0ezf/jUKgQEJMIRginEh0m5JVu5cWey8TOpjmEXqhVEWrGmIqlA4aOhqUt8tv2PPavq7
+BRLpKApHH1ZN1k4AG0107o7bseXTyw9u7528pup26CshuQmmdDK7BTrSq0cF8gd9OS9XFm1/Fcv
L7Mz1+A6aIna1x5rvAt1Omce6c6qvxZjN5HQht0Cm83ZvmZwDSxqMMWfzwLm5ANclbxDoEAeBQ3K
stit1aPzvvmnmhvnZNf6UHK9zZKYcTfZLg4CGHhlOnRJh/mg5eHO864mHqaQ4BJp9St011WElLln
RC9V9/9xW4NhLxXVMZ2F5jwQfbXWdO/lDjoLkmelRr8ca0YaUGZvFeHCW6l2OHQOKcY2lA0G4M+W
e0+hvDElKTAHce6DH9MgF+qWrjmNzAKqb1sbvUtmNJY1Kc1ezqXQyFaz6y/8zVzUnDSRyiDzaifX
To7JDkPbHdaLfYWvFpBo8+yADWPvxUArdO84WKdC7cTzsdrhdxsUupK0OuafDqtjycu1bDMjl5NF
3nzPQR9ojKd9R4SxIs/zsmvSu5iD+397jjA3b9q0wkLBZXT45krm6hWJmJEGOzDQJS1qN5o2ouL+
WanifhNsga5pxpm/IxzxLWIkMnEZy+slbFl/lE7Flky4SQOhAAGRX9vazmfkwiMAknLnUMjTO52R
tCXfU7xrbG651p5kRIghMGV6jPRUUoYBQzBp/BYtt7+IlsEXrZ5BQscNuK2PV4Dp9InZBrOjTOta
JVxRqvlqTvDRwAvZiXUzWoBUu6lUf/YvglHs7JtRsqubDaRrK5FNR2zI+5JLKITdFPCAuLzpFjH0
plaTURkrK9haCI5Txbhy4M/TC7fgp4XnLxlEkJMOpvRpx6vJ+G1vLvbAnsBgL9goobMNUgWLe7ig
1KFBPF9vW7xCAAhB9aG4hQ/XN/6q+xqk5EJ9GbMfWjOKQrYiScH2xsa7CB/ezf06QX0Prl5zRwRG
vfypgZGIaEoCm8Td1SMn6KWg6uphq3mdrEl8yJ2mLNXjMtWAq80sSFgAVnG0njlGI//656H4y1Gw
D4wfYjMoR3pQuhcChxGVdHXXuR+Vs1yTPnYyWb0TTQrFisoVXPu6fAf7oGpUrTzWhgQWe7zjUe/Y
3xboYvp+EGkWOzIntkr+7BtUFZqtFV1fpqUcQA390LmlocrHIX4FY6BY7Yteqb2vVgliUahEuaGk
qD0296hTUZAMneq4iEghiQ8Ztxtg2Z6gnFyMU7cljM03kSRjmmAX+47HykVgJ4JpnWnH/bIifAGu
U+bAv+vMtVxPaI3KBvxoiQNKFq71RTJdQW3HW8c68awVS1s6iKwZ11KnPPUMATdrsny/wLf8OnA+
HBxZ0Fv08CBn4Nd5dIyAlVlBVR4oYREYjvMkzuKKpA4Hb0cF/P5G+pqb+pzBJ00OpamsadV3uPpw
SVf91FPqO53MyjnW3B01nvVnUiynh2O2PXQSYJgkYNVc9RsCvi9HeKFIQwAG4FFO9K4f9uYRykb2
nIu7DRKksj7ONA8uM2dWN6ZnaAJkI7jVavg4/Y3qH8N3xd3tudPTUqqaTLVoV9pwepwHnaSX3+Wk
zCeTUWEwkj0fUJaYuFfnOvlWyVP9oq23r4+jj6Gx+uiwOz6AWAreVh17MFsF2JavdTU3Ah+aUYD2
eHZovrq2w8FB/U8Ok85W9BAwj4KEBE+OZ6zfA+1Sxwx5K4I6hPkS50fwMpnwh/GQShWkX+E//Ylx
a7qnOEYI7bXtS3enMUtJRm04A5GyADyHjyX+L+AsLsXR/FRcNXgskcDUEFpsx/FPgsL+Jop3tPXo
0/vZGUtoORtdqHb4V3EuWJvZg8DhibNi9tfdjAaaitk7oxwBzA6FOBWR4JRk5sFiiTycNwCETKiU
k87O3dfvBri2xHerWtBkNe/H/BOTA3/eppCh79yiv3jGUg9LGb+WX+ZuAszX465SfZRdCUrSXXNr
Mb+KDUnqbLpT+1uTMw3s2r1lYjUl8OuVglyRB/JUFpuKIRyLwZLJM9ocVfH9DQ+Wz/cXB5ATmCMl
cQg3uG6ZOZd1jkbtfKnCQr5XsE2ukaTZvEGnAcfoqcxbuCfYGKJrE4jsd6BwmGmChtjgWlg4QNXb
6erFgnvWSvbWFc6WDLyzo27WJ3EL/QPJEszCVcQP9nv3RQRHn4pCymeOnHT0fbUbbdyIEGlLrU98
ZMpCkRDq1qSy62WEBjEbAMyafdNq5iPC9qbulKrcSGbbu660Du7lom20vCGGnxsXqjJPRBH4wfnu
mGlgwptwe8lcYz9HrcYG+RJWmoOY3LHrVI4mhvlw6LoLVJ77Qv2IJBXClmsDhvr1xFMl4M1rH+cz
VKaDCTV8UKzL76aldK86CO3Fk6AiOqN7O2aYiPrlsOcGEjQGqDmS3ZwtcUZrHukArt6OomnUjQXs
NaUDkkCAqZG05D2KjLxmWPoA0cvMCN6GUAQ9EywRBx5J+I5YJR108ZSYF7kS8iuN31Vz0jgI180B
n4Mixtg7eDhcf8GUDIdg9gKozjb9BlsgPXZHrlkRR0SanaEuwjv/eavsdmFIfZuU/TwRaWDdWfO+
ZulLbNkSq5r/u79O/S25TPbxxJ7wzzyAPxes1pGpBg8r/Vy9B841aujtrdaaMQ3QiONjKqu5gdK3
AAjnUybkUIXSmwep4xJPEurURt8hN/SOtl8MREvrtRXF1212WAoApCM/RUKPzHiVtibS2VQ5Bu6u
E4WCJ3z9MbxhtpVCcjSiqVLigwbCEO83N0Mt6bRurfoGcyGkM4bi67CFktWXUdqzqJeNP5tOaWR7
G5bFwyc7KuQPGO2VEQUIYDLcnzKYrOxso6uCL8ya3e1RjlawwEKNX9ojfnmN7FUAgOqcWAE3eZAu
pDb8/i+zq/ieDs+8+tC2ca+gfolcqCe5ART2c+cgLSgGMeGdSmyUQbIO5D3xQPhj/uxeUqT99Jjj
XCCr8YQ6ov24K6Ny9oXPbTbjDavBIyiS8FiphSG8m+qtVpVZh6BaJ2ADQCLgMxzNkSSRo09KtRuw
nAXQlb4Tb4o4vABUE1zM9ubynVDi1slXkgTTUiAbMWdSp0V1mk/690zn7dYN39jXnpLecoh6hE8w
wONuXYB4/TabaU65huftxGD4pSqhE2v67AomCaHkJ3BPHL2H5Es9JasRpwjr3TuQf7nIpeDFgL8k
oNlWBgs9zhGO+3UVnrV0qyWq9eUc8j3emVkLs8xm3AH3CR8SJEd6KljWfGNkwjGkd50wxcDba/r1
ZylkmWTbqLFxxo5fdhe4TilH4ZEzLVUKUQPG5JOkVWSBHuHQt2s6wQgZgaoe2h+SpwrSIAOAK1fI
qT/B7CWQUDvDeR7EpzO5BJ1OB+zl3BYZHrQg5UK5oMCOpsKvWKQAXJ0Cto/EF7ZrHrC1ddYzGngE
oqhsVDErzUDw1KTskrfldIlu9NK8kdHz24lwk0LeCC1VkWTG7GaAgBwyFquUUNA/SFqysmHbY8Fg
BUQ9LYi52RHMWhHQn/mQKCzaRR1yVKHIbFRdQ/rTNdVwbbKY7Rf/IUyo/aFg03GosL7hpKSLwQgi
1cHaxZfTB4o1n4QwF4RihNwVBpxkyJJgNUZja8ZPywSZ7PRamf4ony6fJBjpEoqWB8Oi5NnJ3EYH
LYYAnxxDybVZMRintlBHEk4G2jlaasu0c1nB0a7Pq2sky3UOTGtkycmCRc+vwH7W2QqxdFkSUY0/
XKzNQB7PsIIjQVCo1gYZIqk5aIwQgs8ljV+quCl17vAiU2wvuDe24U6y7MqWluXtIW3mP+0gvrYg
CrSIMHH0isGWhuTdi9oFxBlnzmMqahq2JdHHnvWvA5sJGMHA8KqZQ0f/ft8BOVe+br4Z2wAWE8sD
3NVRIKx7ban6JEgosIJW1RMkXdsx4puxXyaKaoLacK4YCIdQ/kYQ8wGVLoBp0rlFeO05REsyY174
DMD4WF0TwCzSZTH8aFrlXJGEnFp5CVGelhLXyPfmxN3vONHh0/zezr7cW/FKXu8uBnGFfkKDEV51
G8hlK2WPVaxECLKalT47bKP98YlyX+l57PxNWYJxqDlzpCk4yAdc0Cxq7KJR6cTDIF1doeoHyE8n
mWiLtkOLGKN7qPBW2xbFC/UsxI21vWqU44udPV2BGBUTPB//nEElMnagX80+pf2aYJ4EKCpkQggc
/Nnr0qyHN/wYWtB4AegMfbKddV3lr8yFHPt/AL2Ybptth7J4O9Rg5zTmdvSWAcKO2Xgv/z40cXmv
+8xzbUBrZGcJ1HobeMEdmT4/Wpy/Ml8M8wfIT84yNvyq5hFFNDuM1St/UwBrfI0qk7LCwjRQersB
H1XkpQvLqS3CKjWYCGSgARF+f1JCX+YxxdbPknShbutsAbqIOS0rF0VavjccGUCibrmt8elabR1l
VAEIpKfr8WIf80qGwVeFe6MOmKUIGlIrGUMT0xD0PObw39BEC5yQnNaUP1LjH7sCDhRy3uBZXda6
CpnqHIuBqHg+DUN7LnxLhgFqkki+N6b2lf2samQZrV/4ZxreNqpPj5pvQ1wtuVk/a+HVHPE/2qdc
bIS3s8uVEMeUsmDwf57X8U+H4VkJ4Q1L1rNojsDVPUQnpJN6pR33gIuBq0TfCCi0vz0Ef9UWEl4+
pwL4gR7aOJmxOv9xE18efbpza1ViekrqSdouPwuSN/46BZRUEWQ2okhPMgp54dzkjr3odRSNphI1
pVwIoxUQhXq1f7TNAfqqOuxoSq5zX3pPgSAswNKv4rWFz4lDvO9WOTTkB80iIKa0mWv5yETES0Eg
Zv0T87tdDQWg41GAQy1WR42Z1PwIlxEan9vMwyE/FIE5gjBUhfDe/gmVFg2s51lLP11SruLGgYz+
ACSCGRhiqb70wKkQuSQ0XGzfkVPi/gYWdOfB6Pybead95Fk24GnhXtKmZE0fKijhjLrd4qJ9/l35
8swKCapvUTkR/SImzx9DV9rxlYhlfGSZQWA8LmXZWwP8j2cdwIYbfrDjvFl5JCZ+LVWdoFQ/fJOu
rzJRrWHRCkf/m9xKc5kVJZULSoOmCQ6LGK5/Y4WC157aK6vb18pBsA8VwLfm50TWIEmb46YUS7pb
Xo9VX6ZGqJ+cpp2EUxhg7d/LKkN/JHcMOju8AaKZLxI2taVskHteh+Ng5LxBXUfQCYdUVQLn1bu/
O6lrbz7KgXJ9Xr8G2IpVKSZVr3DwLsHIDA+7vOTFnr9PF2XZgI4di1BjMSa+R2M6yQxQ6KfSnkuR
mFSjd7ksdsm6nVd7IOiouBwITtW9JIWGMhvmTtkgj8t1yOOe0WvgocJ+S1uvPxKu1Fz3/sdwXFar
axzScDysp19zLdQtETXcuCCqec6LFLSSI1WW+L/W7ZQmgOgtNrtQZ3KL4xBIa5er1BO81j0wZgnt
AYTQH6xnRpNf2ijxT8+2HX2G4iOvRXVUdeZZ0BkURjoE2IXkGIcJsPW/R8pkQ2PlD13sOqkNrgCN
0eQMmqZY76mQKUGih3Jlz3TSJM11fbNqKx1OwOv0NKBI4xOUxJrnhlj00N7wbl8grs7luUOq29su
VELz6xqfbJAnPFd4Owkc14MEBQqUz+yt8Ne/Mq5l3L444JBCanzSgLbVlabURFSsHBz9ePwy6v84
4OrW1x1LgPLvkIrYidnIKxVNhkClfIwzSHJTS3m5r28BrdiqCecyvDg5J5wK9gc03Mkua4f+7udk
HhK+h4EZiPbGxFhlINWsNoi7omE2bTBjZDejg/aLck8q1RXQxJt/eZ7G+DMEuU9iqfWSfEdj/S4q
bYsdHb8jgK3BrJPXKY0Sb4ciSIAyxyCa9aSoF2k2bEeWoQnOtYM5Kr/jOXktOKGyvljcQTrMN0ih
gLH3NkRvNkiRQLFcH9kkkoH85ZTDrr1d+HfuqWBioAbru9uEnEx5P+3M/iK9zt5idTnHFpfjuHL7
5+H3hJT0KkZNzbbqJU2yVUrDJf3FSW3V7c20wnyWMJrW8qL0D2QkvzkrWDhOWelt8NVxfKRuVOmy
eF9tauYBqNBxCIOr1//bHM8IOL235ePNtS1r9HHhw1MLTxZDjrQS+iexy3b3CMoV3Q/gcYlc8J03
3/QzharlQ65KNQn/heOT2zkCkC+K3u5KuZfJ0JPiYmlqPWCd7Hihkt9XLCw8OApbqdgDISmugHCe
alY+BL04TiS0ng7x7bpo1/6v4iTyVCxYBVOUCuPC+0Qnfw2x9j/VfThp+lLQwlZyHaTMRcqXpUSX
3GYOqTIPrVvTaUfw5QljX/3sMO6+d7GsvNjbpKXJKZPwvx9l5rU5b/qjwKgbRyzVqYwgXED8eXJP
RjLS4NSzprpvoF41OzNSYbBAXgL1C0G0pkQrxTrLxQOFXOde0uq4yRO9e8Z1woOkOdYHEuDA1Sbt
w5o1EuD+3C0zJjy6F9y3WNGsF+RclQYB3KsvQrh9J57OaOGDUcF4OcDV1eqojgxNlGGQBhzGnLx6
9Yz3GsxZoY9wJNztaejgVzngjYCMzDxlc6MMumYIBgSHZqzIyjXHOm6CMPwXzbXEDHyc5ZF0v9zd
Qe3fGnPn0Ul2BYuUBqGm3GgUB9M1PsMGBIh9axq1QMsFkSQ+5wnm2ZAsVB8JBScRdgCI/NbaOSN8
7jVfiD79F2clzNgQoDdxwbdys9TFfPTpLHXBQDd/BpWnzLPs0v3jCLG8WAbq/DZZBQQ9a7cymvnn
nWY4c450/juDebOZxX9LWzA0oZ9H+lg9Y3ejKmnW0T82tPa8kTN/3ZrGVz8C53hL/tFlaAnAybdt
4avr13i+hJkx7j9kFMcL7kBEPh3CMNS+yq4LZmxdKcApYufsJOsoI9r9bqkvuXHFnt1e1OKuH9RR
2ZOLJQnvQpNScnE5ixzHlelePxsSoP+B5swyBVXhR2ScoU9jyEIgEd3cwVSZs7kIyDACgs82/svI
tt3FuDJzyegYAxfBkT4RPPLT1DrohiqWyw5dHT0U6W2nbK7Nq5YMbLrepoObfLq/L0NhqGPNPQ/J
p/N6x82nW3qrt0mOitZkcDjxWBv/bBk97XUpsukG0CLZYWOq0pMxvbs2dKdlJOfE/PIzFOkAldc9
3GU6jUl6ESuRGMABjZvblqPnJBz6rBQKRJbCSlr0quEg7BTDryhPBD2KTUU+Fc55lKew3lhhCSee
xXqcn2dTRglQ8tGqe0ZkEqcyU4Y9Zo88ckr65DBoSc5ebbIr8vuyJHmdP0KHZUQqKaGZiw+KW2PR
/elC6sG2GW7Y1WYdB8PHCSrWJWPYIH10khzmjQh/DpyCom0wJ8gc+TbhWCBSsK+EGYdKjoe6e9GZ
Q19Ng5qt821v9xY/1jONbl6rr4FniEk+iTP+NqxAjndJR+k3MLFEHKd8/SJY/l9puMAGU7ZG4VRe
jlO+vrzA4m20F6O5hNDpQV7IOxskmNOO74Hc7Wod4n4jxzv0HhqAyboJGqFEQxRLpa5+9wHWRar/
ppXPFVlvKOOXRuyLv0DPb9FgiLVE/bKdUgieWrO39ZDo2pRnmo7w4hdaDuZLG4p7cggFFKyTzUIl
5YQf+Ri/GTt9Lbfn59e4TCMlgDi8gSHy7Yc1TrUADwFwM80i/EmCr/vdxBRMlHbQCRPf51jD6UeK
cl32jXz8t3SPv/q1PDLl25DQVBrUQNwkgl/ABo9XnJfOb8c3kBo5dGcMHG8VH+m3KZv/xkYdCCbO
LLERdGAfI7Luyqxi40hk8QM5NwPpTtydq8ErlnimRhcQqh5oIfVnZwUoisIQ0vOGFlPde3e1DDNG
eAgdCB8XZpV7qTFlNjiZXEmxcxQKdvRrGJeTPihE47jJc8eAEDceqXCMntLnunlVHcQgPAkkxXOe
zygVANzGVqIrb+dVSfBmXrJRXrEKmHuwZ28xdfJ+bqkH4xW80ifCmxBVopH0WKp36StmST6UaK58
TwyBXWr5gRP41eM5gja/ye01BFgFWZST0VsitFWMMm9ESmiUZwL5ygpCwA+uZpdJ3RoKZBe7pSx6
xn3SmHFMvISTXfVszB1jRs6MRqMB/nmtrxNRyX7u9C66P9cKXsTMq+iU6Gf9Z+sFWMFrhCIyVUm8
T4qxvzdw2KUaJ1XtrsqIdTXAofjRdIcsRjMJ+W1NYIZyCW3idqCoRUKtfMjjMAaVISSN5aWYv7bO
mU9+SbRfUKmJ1kpq5BBbLeu246NQ8GnEmJVY/W4WqqQx65WA5TAozzz+No9885ADIuhUFkTnbUJb
xPNDceP+z0WNTEjSRqjyj9qBLwMGCzaO9zbtSL1DOCkfI/DpJOKFJ8uJpx9yrdqRqoFWZQ7Z2jT5
6e2RfqvouJVdYapGNqKgWmmKmzfcFhljf7nwY4AG6LqNzed17zCr7Uh6V+jbHQfBzeTNTb9UVcex
3S93jzdlger9u8+8Pcdk53STKkMo/YHWtrjfw1RQT+0qCU6YVUsYSMsb5mIIZDliXrmDWTaN2nV7
DOwyXEHCFfzqIbLBfSwAdTQwi7Yv3kUh3UvXihlDdFQdtU10IMc9Dh+Lci+t32cf1yjJLxbfVJp6
w2bZETO8auX6iIC2KPs4osXikVXkOyXqKiqFoLttIPlq+Bcu420TMaLdAD8AZJtp3MSkiFjDVvrr
Ovo4gDYGSZoMzEUJNme6ZjpwfWQYQagrE2x5CYJyDmfKgqEsY2TTHbIj6qpKTPnDWbCrb/U3C5G+
BxcnWwtyncDAv27UcjPvAh99Bdu+A94CDyS/gDhfkIVKG64deo4+edGEEAPs6fY4vWoeV3k19RkE
ti0gNV3+sQKyMg/Yb9VGb9j+zSvQHvsYG2m0ndnfl5RdovXsz8srWCuVj7KdLzzYQiqUt60X+fwI
ukR9B55GonHgcJsMy3Qtco4bzAqa2loc45fU9cOTdqPPIvdW+/wYsjvGu0Ko2RkbWynQMUJ0tN9U
1GJy9ET4wpjTDIR4xkKfrZ8eE7LV6vQIqW/1MvR+O37dj8xQs6qbErDroHVRtiFcUI6gRY/hzbN1
keIq1sTISchFcd+ZN8kLJmNXronCRbfjHyw0MunBCD7SomF6k7nY7Bum6YKuoEDaS9XumbxCsGeT
jVRk8128yxN0aEcUYHe8emU54flPS+qqmReG7W0USdZ62F6MAkblRLkp3yoYkBw1zb3rS+kzlId3
GT8kgS/7Vm5sQlNwZhi1L4hmsqK5kkgWNgmFrluBdFe0CZzMq4MmCvNHqneNtDDKLZl9dWvp9Q7e
+MQAKdjo39a/7UyxkKLevcp/LulEZn6YsQHzFjEJt/yf1iusXmTZeutnoN3znW6TlSOZa1i4m8MC
pOZ3sOp9Spy/LTl+yeeeQWGTibotXyN4ZywtpJHRvww9QsBIRaojp/0x1U1d8bolsUxbt3zrM+KM
lV5pQh629iFzjv5OaH6i7Sc66dtwyXpsFw7MruVr+56TTo42HYFQiAacWnftmG0egWNBF/NwMY0M
6O3QIwGI3h6e/2xxuj3yxnlxsfqvoNeBkKp6nu4pQzHVxlq3OmPkaA+3ZE3V640/5NJC7laXgonF
ffNvxXU+OGTLtsCf3VNZI9INQpZDKrvDEDNRKOWHd9jjYM3DNya8xdktgn/1PZXnzybA//NQK9/e
ctWI6FdEr82ETR0cqCJ6HRWzSpBo/sn52WcAYnmm2H1csfeZMYc96nPGmcIgCzYrgY/XyTM+GziQ
liVKru0ETWNq5GBWRmwYtPJbFlb2yiSJ65RclZc62KKfaoFmbrX5ca8xz1pfJKDQlJJgfdmb1ybh
iVaIvTsyAEQqfO1+icxNeWlC9xFyrTTigAKFkO6W+TSFTosv//Li5jqtfYwbavsFaDOOdVuCchus
kNHCrPrCYyL4gZyiLk0cCVEOepOZ0i6BDOriHUcjd2uG4CluYiergQmV42msT33Uz5sxVWd8tJc2
zRd0vx2YWjo0wh04yeNOFvHISDhxUxDQWe89TfGla3Ik9aXCtLryCuGuxn24EB1w7d5omAlBXlcg
26lxhrkMUh+aCu4TxPLY0iuxxP7XarpJ56CRIzjYCVB2+g/ptZu37IL7WvANWKK39B8n26R1kUoq
HJ1Dbqlsf36GEV07cQZVLwGZaSh9Wm43Apf9N4TB2BzQcIS6yHlbDKittJ6Me3eoNJyRPc5MiGNu
enxb1XYU598FsHMQ4bFhMknTF4IZMKr+cdehWFsaXMCS0GyvyVtKZq1JaqAmiWVtatWd068mo5TY
ABY4B32VizSVggbUT97flCGw36PFNMNtWAKol4TLu41vf72N/gC18iC+T21/5tYGV+dXLgKY5xpw
kQNHNVxNZVN/9IU2tIVZWEztja6L5ngxnuc/aSdLfEPKbAHBg5GHlCUip5+Dih3y3NRPq+9eQ3kW
DoNz9j4ex0ti9rYzlmKsNLLWTYhNJ9Jtjrxdy+BnG+rlOk6RMZWoRJo0Xw25B+L8zR1Uzo22TVfo
0aftyo0LIkJp1C+r8CXm4tA3w2E1VffLj1cGNv5uWs3xNZkqvGlxPKpO0YAllFtEOM8ROFuuild4
Tr70sha9kBymDEuT9eF0wWjGaIWZ6nsu9CfgAhlA1d53wZp4nkx8DVyrvt87WFuyJKKby5HfX1L6
1NfW+wuDfoTQDgcLE9UF1a6iTwW774JQPGnvJegK5TS/p/YDgmEE4aK1slg0QMwJVSa88duFzVG0
C7l12nuhLqDo8aRVP2Jpp8CimhZvyItYR8eaW1oWSefyrTumvgwEvMO3L6rZ9TsrCha7tOF3tovp
a6e+XqCtu4oubjy3gHCDv3TIvsQRyaBZ9yj9esfGpTLzNIInD3mli/JpWfpb4NXTWyjBB248Fza2
JhXLtIx6SqjL1N5C11RSnjNJ5+yNBJzSw96kliHkXIHRwI06KdgTWYffxVU/BRPSV5jyHMAuKe+6
czZzmTgw87B/afthwz0GiCqiQUrftcKJkicPqVwlSCWFPpCveWeVlurr1LPyej3Y53eylMrgGh2F
MOKayl0RTxNaPhutP9OC695jic2zEftLkUSwchwzwTt/5zq5Y1uif0YqQOsynVU2BEBJ4dECbc4k
sLR8FABb7/EdKz9QB1tisKDrxHHKYUQfc2WSf2AjgZ+8CMyUZv3G7mssyy446AvdnwzlgbWjGhpl
UyNjYmRqgyhifGKlZ42N2Bd9BElBd1QAtTb1HNiEe9CqZ5L+e/G4scEYAS06nFMSAjY94IJdqwG5
fjeFIg/Hyid8rZ6xrCTKC9TaohTYmTswvbaPLsk0iB/YVNz9SUT8EG/noxNUBmgMMnFnLEVTGWky
kUhtxmbNGo+cU9+jNvVF5uwePMAzGtfSVeVGvz0WMN/kldPzHP95srEzUx9g7lPRTE6htouYL2hX
VRmUli76rstl+ofAMmm47q6JIPg4+Bk67sZUTiCkQHLQ3kp9+eg4wRypPMvAreP0WsFWIm5jnvf5
/0tkLyrf1X2rMuS5viYCyfRqY/AWa+Ag1R5PKHewvI2qmYR35kebsRVDJ0aMuGQk+svg/GE+9Znp
66OsjIqH6humIyeans5QQ05kHBzlN+BdyyFDab2z7KJsL8fmaDOUr+hhBPiHjYzIwnYwp4wEOwqY
VIYrHUewCrO4QNtetGjIyGSjEbVNCyHNKvj5oDMN4iG+tbvSm8KToLjMQwbRP1VcGTAx1Y3HtCQd
M825NqtPCkEHK3NoYsmoNCEWQuchNuX859o6BC1PU/7U3TjnRDun7ysQi31uGXxmrN7kGYwG773i
WPWs0MZlA7n7EUITGrMtPFFl34WqiNfV47/fbjDfwDy6WG6lr+X06pguhkAR9xvEbT7eoQRQTxtA
1J3Uu+R2+J4zc8nG3wEyJXQQ74DHVMzitWmsqo4DGfKsUCwItudMte82iJT3N6D8puYe3VCKdSL0
7+aaDj1HAJAq570X7MdCQNgykgaEDqy8TYGBXABZZ7i5do5Y1hGGpMG4a2Zc+SEhEVuDHxWzSb+2
WCNO+05GK1mHF+yG8L3fZU7qARGker5OTKJ94BxFo9B4Y0+D+Z8ZPsv46OIhiLt/y2WWq7hycBeN
90tkTJZlJzvrcIEPSCPaySoBZ3IwOMqa55IEM73UieCZruRQYmXGNELO2lPl5g36sKeINhL9BvY+
GcK44mOdqC7gnzoxXHjbUh6uxaiXk+0kM1rRgmU3fRhEHQbxjlfTePLPUm0vm1gCocWUaNWZXu3j
77O2wfpkXHM0CbYFDsh/xE26FlxClFlg0YmcuFkotFcu1+UeGdSxAhCe1zfjmXSi4BdklThPHYSB
zjBbkKSIgBbzOBm7nRUnnn2lfycT0mpq7/aXgFhX+3OfwTn2+M03df234VNv8ya6pNyAHP0z2jDi
mE/DO0Wzqe6sjYK8bXs9rpkbKJ2O9MQmGMSjMLCqUfF6dUDjerd3eaxIfHEC0BZYaNL3R7jU3NeZ
rS0/053ylwDg8OAQzDlwGUR9mhLMHESiMd2IKXrM5ZwEIm+x+e+HJbN3qNeu/l+K64+0J+rL0lx8
BQ5uHpNwkojvllB61mboxhF8LvXiezjO8Bmiz0Dh219MJtS1VrNWY4ihYrKannAP3VcQoBdXh2A2
IbI2mkYypLHiJCnmImDtsIcy0PrABeLJBPB3viL1I5K7Fh81q/ByEByjFYj9UBtzbaHrw5sxb1/e
3YiMKnxuuvAg0nDdOj+a69MZY8JuFBQFo8J0F9lSE/ODJgm3d5xti/SKqS/WNXZYnSF8E/8NLkoU
fpKgi6p3wprQo4zhRS4xZa5BR0PhLBk3CgKg1mELUYsiLEE1lZHnjm94HWxly/3yYUCJofEktoha
RCWDkSPcG0L9bp5LgrI2kib+oKp0mONFGhGvcebk3PltCLUbR4Q79UzDj1yBaynZGxrE1RKMjk4Y
kHTjMd4BRGTdd0MRPK2Bq1wrs4PWBc9gkRyioLjDF6dczR7JSq++YZr3Th3EslN1Cw6vEP2t3ZrI
Lzw1STZ3KLGcC43CGBonmHkFxHgfGemMDGpRiknHylk5EvhZD3U80EgRHWA+/382pn1YYlzVhNIr
3MqYa+DuY2poYogoIZZJTwkrxeGg+Ty15/uqGo0huBlGwFsOBChBYLNOCM1kKlDk7+AZoxx1x1T1
dV8Ks2SQnbHCpZ6TpBaCdDaeVLuQWH07AaP+Pj+19cGZiIGiXNUCdmbLP/S/7ggxPWTCAkA6aBIj
r8RSvdmMheelNCLahLMywl6eQOO8zk6ysU5IRo3NXx3OylM266hyXxkxoN7PyJubTfcE7lhCFrW8
YBsE/YYpLBhe/hdH7GsnSAjgL28CXxQCWQSvcZm2t14Zlrm8umQP4APJQzQOdiK7qgD6ku/iHUPG
LmQxgRPY7UYFmmGfkRav0eyVKef5xnMCvuVvmcnq1/V3cx05GvUEWYU7QI4ctKRgVPx+4urTjmmB
HN6++jvijOWezkrqzM/jc2t5fl9Iaa10m076kp5EHhQ6EA1Pw3NujowhJ1tRQtCvG+V/t/n3EyYt
1Tls768F4LM4a80/+KMff0OetXUoQD7bB2IUMWwS5zE6yHyxIDOGMeEGAIH2cEX3ZzmpQfHvsHQY
0497QQiQSw3tLIXGHLDqjyxz6IRuw6Al1UVUEFA7+pZcpivewcA0YbjgMWXvCvARmb1+drZe/+al
2YRLDGgTECYZ3SpRC+6gb97HUZdhazODhABJ55m+lbmdCqCigE3Kks0mMRsl5khS+Ggw6acJnrJP
0++UxbrxTO3GSsC0DlrjUm2zL/JhQOkF5biSHQCSwJ7C726oF9Hq31QD5yH6sTDF0f5pkDJjrMj3
jXj2lYYzWNaniYP13YbfkCtJNSiUpZGHwuJRDUm0h/KXEW6nb5MbBBKlLMn6vuDETGWIFMmwe9MN
9y4RXJe1A9TpVVZGo0bOZjdkwBA4qg66J8N5LwLqrfn2hEF7dZ0xSnwViTcJhYDnpdWMWd/WTTkJ
yZiipnXHCpSijWl+63mhHsn0+sbSA1huObWmYI67KiSTtgfN/INJVsyZnUvjAouPApWm/uPp+W+B
PxVJ5ccxV2pCT3yyvXljnHeDqRnY4M78LCfxWKHrR+x+tbidGCWbaQ3ultI7cwn/sM4i9JJFtmdp
Fvqzvr0ZCtCg70j/g/GDQ0mxZ+NF9gMLu8cyW4TSI8u8z2BNK3CQU9T6OMP5CthcmZ4CB0J1MWw6
6+Ed8frmI8amr97CZDx6W4WGeKjRlHjqx9efP2KhY2ltKP+5dIkhe8EBTsY+poQLghH2V6urd+KK
1HZS+f9I/wb2cUFrPns111qMcnvuGd6YeBBHzkyKr7ZzccZOvs6LGwfmlbmcTU0rBhWtw6aze+sC
u71i/7pnEzom2ihiimcTxGjOan3jKi0VkeLHT1/6etISwpNNowknCNl3WOgEyR5Y8b1vZRFGyEoH
HHnxPNnMj0XHAe7a5VE274Rjl7ogioLZrUCtSTKlGli/F9M1TcOYsVqaOrokTb6sArVDnr55upRj
ky2vDpJ4YlPl7C45NilczGaIN+yMfE6pfUdbQsdz8yZv9WScYWNfMEB4dhotXgTxa6v9Ehpkx3fA
/a6lpYbiJqyYqlRfWlNh9H3myd/fKDA5jXikuNtNvV/bQCEVzlQ/jT5Vm6CIo3+c8ia62lEVUUhu
cAihsFG3OdhC2FA3Jk08pZ2Yoc0X5f6maS7WcplW4rdwSWK0tVE5lrRpzGrTtGdr1bavEU5iUs/M
PZb5ejxed8fcYQjT8wbLuwDaoHjR2Sfr4zf3F+Hi8R3eXMHbYl7JpUSCLuBud5d3Pw0wy4mKm2A7
HhOMzrYRkFKWDS05fQAgPEZdG55UgSOR8cZof3db6oyXvif143EZKUEj8ZTKIvhjxILlr94kv8Vc
0MJw/4R8iLGGZW5A9uGfU78mDc6AYXlx9QDO5V3jqUtsYWftURyTqCcAqp4LY9wov7GusuhEBmAx
znqTo5lYIT9KEpCXoTCjug8D4pvn3miTAr1YBLvE6JK2LHpg12eE0sotMzgt8G9JhhDYFQumNOPr
kBI2SQfNbj89yKz2OEfAZkZMOaqqCjNShJku3seZQXkN1VCm6dlwDB1eGJeOqABmpv/bGYAG+nqk
ZxBL4+qiuHSdgyfYlSjlaXnPGZGQhBa/vPCQL1fAvxfJodKU7MR6/ZwScUkEKRh+HLkkEPr/Aqwf
XZHdedvmU0gQIMtn5+It6XJjQ/G0kdVnWbsGOBOo4rGX8AaCH+dtenSQUThqZjH0m87X3KCSuZz5
f8ugIVdUkPrSOS9L4maQ1wnMDwbwVAmo55bv875ulZBuRwUGrSt9IVSrvY8eUxuChUc0wITwe3MP
SnMQXjaePzR4VRqW1OR7PLCoZzkjHOfmjh6QJ5Yb2kiagybMG9ucvLg4iw4+8klR1bjgP5SjSDp0
5ofa2QyNFMH6gaul2Ajmh4MPir6pzaRpIzO5FdLGWlIA2Fqo5us8AbCSiefoVr5sINVQ/IgT5hy1
WzOI8W2zs9NgOk0lj7wUA/BX0k+9rbfS6JWBaloOYgRnlzrVZpNaig7Ze7vr2V2J//1bOII0Uckp
ul851tZy3koo7TXZPN7zFD8uTYZGd94roKa00n2ox0yHzWKX8Tbwj95OilKbJ9/6862huOd/AON9
2tNo2c53L8KMpmgDjufSiXZLvftbCx3dsfF2lIG+PWctW4C3QGvMAqJiayi+AMWMk18b/9eLbcir
kAgAG0lnaufIOR6CsqDngBnHAauXSVIQVxIOyI/RZzY7lPucgGTZePOsiyE9Y2xf815umCdHifx/
k47osrCLHH0QmA+t+EpG2o/u3jlghUqUNs0How0DO0tyWhDtLwLK6xQg14yDDgDCstz2Mh29m956
3ncABuoUWFmy9053a4AsDZN5jjNRgh9T4F1iUXK40dQSqPA65KqfY1sv/ygca0fkXcaG1R4DMNpt
AZGEs9Q9dWh6gg2QjOzOxhW8zA2n7qtCacdwOdEBRtEJDkgZEe4lWhq3ttqxkzB6kKihZ+wQgC0p
vbeuZveTbj8+zi1LVkrSMLYMHnE1ouvj//ruBOxm/jBUDjDHVHEUTxzqZDgUYLa+oqTOCQxmGDF8
/5w4Pda4zLAhGdiXWyqXYRavaRR1s+5uy4H//fL1jDdGfjn6RezR5V7O/GUm+Ddyrv+zTufIBaBp
sRoChowRpKAgnuXXjfGuHDsuhZio9PlRuenXA6jCU9SY7FxHgPlRwBVOXYhqFmg7i8q4khjtSeSj
plYRTxABfdNOYJgNEnUtLXL+W2jU429uPvm1uynMn4hsV/tMbRew0qy7GbicztirO3sa3g8sgiAe
8PXtgpZWrSZ3iyDyQR0odMIeNWuvJVP5VyikYFHyYMfkBpVXPPH/m4Hwe9pEaIq9HmI616cGPuRp
5u2PstNhJLa9U15xPvrFjq3G9Z00j7UYIZt1/X5C6woCN3CPlW5tKha79T91rTZ5SJ8HG96invN/
pW6muZbc6gumBgsdsDdqrSrRffU3E95YgLF5yc2RBKUEiIyGw6KM7002HKH82BgTOY56YBxoKPLC
cpcWy5NdKK0btUpefhNT6XNvBaGiPW+Fd824zIlc9FugTeiX6m8Y1CYBsZMUlwBnyeIaWdJnsVfh
+jWVU6Oqun3zX+KH/FGtMiAvNz4kPWuFkazsZzmOESIaPzTOa4lz2uUNy/Z1aNKckGCpfkM12VmU
t8JIrxxYscf95/bzx9rZv/7e7KCzM17T1xp91r2Yjexf93WGKa7UzDNkprj+fe1E1revnVFPlli3
ViztFF8IXZt2SrtWMuAZKn5uDT8oxikOrcnSZTxcOJDQE8mYVHyuwd55ow41PhqHP5vP1RNX3DQ8
CkSy0EeZdysvEC6i8caBl8orrXtBq9yC1hMBDr5AsgTxPZUMnZFCfEdEuKkAnvBrDg9FguB2QYOd
dt2A4HCV1uBCDZWGpq7n1up3C1c6Nm7ZdBu6ZuWBzDn5yH+zE/rMKBWE4d0BViBnRkhKkgK1gs2X
T7fj+eP3sPQLWDWuShKbcFnG/m4RJbkcK6tsHzGL6Qn/JejfLiJ3o1BDxcG9C45pMfOZD5ZXkhGE
Up4iN/nUa9yIAm/W1FdgKuF+2Y161xRNEsxVb3zPq5OZtxL76TtFw7sN6ViQzHWdQBKi0bGy9ks2
6bkYBhliHo+b/MxhgvNxKZCNchUJ5eYLqBLXfTE6HcRFfgKD3nHUxsjZwS04nVly51zYW0GLRTFo
7gMQFCy6xjC0Sz6PV5hvs9rY7032IPPT9SvQNagqYRjJLmq0ZPPQTRYYTy8VT4ez+W+kPUmmJe4Q
H4OrVg60oSdp/XSOBHhRa5Xfgijr1eXbLmmSVOKmziycdrwOA7f17E6uLkkmgvcgFXo3PTHcXepY
7Iiog6oAQvns79LUBNLGfO9zADcjwFn1ZP4TE7cxLMmiK0+3zWdtE5CvrjtFf7VMMa5qNdlQryqS
9L9NePvXAtU7n+dClmj7EefGfQczedhK9RLqJvFI0X+UdmoWC+J8K9SzplfwFfePHhJeh3MG/2aj
WaI0cJet/qt1GnvvIQ+9cQMnUOkdB+G5+3Jn/4bQhV6EZiXQExg3Hu2ecSWfDUNspUfTcu3GXXey
+auRtdE48bX70tKr3pQlH7uO+GqQqOg9PTVkQgHl383k65a/ApuI/UdXz9HZEG4adjV1zedm0o6X
LwiB6S9o5ttJwikte/yOsNzUa5Ynfh94C/h+lQ2Go6pCaEdmxMZexKOVumxiG6CPT2PxYyII0kVt
EjtbeXrgQGh8UZhu8HsCtip/2QW9hlWwRNXY07tdNJDOcY3aJVrNVyN7TKSFTz6VPeZpL3ZPLIkI
qeJMzB3YDMwaWEBF9DfJWSSmE9dxExnqGCRlLZT/bzCdKSa9r/KZgqg408c1iiXRPmtrsDVsoDdS
ihtBm1Rgq19rlj4Dz5zl7GpbDvlwxbWT4h6hRP1UHGQSR66yXO7j/SNycn/EFZwAYTJ5K4aNtFCh
KfOX5y+G0isORnSv/XolhXOinqOj14QHYuJ/fjVYWAufzgXYMxgyGSZo0fCiM9kqBfLM9LSPhxLY
aRN2usen4SzrFaQ+0WK7Mwp3qw8u3T6F3Q+EyhjYQz9OLtHnJKls3WCFTDYYDprwVkmYSzLssMDt
dmfldVw3iv41oUsYjnCidrAlS+E2329XyWGi0rl5J5xK6WLVfgoTNqe2OAQsxW1SorgcQ9kzkfYt
mMjozf5vhmNpjihihNxvvmY0avbyrYyNLGpnvFSY/i5IjDRrFfo+WQzOb4iJpYVd4/PfMen88FeS
OyBCk8rxUo00qj6H6wvMHJyqR6G7qyA7kIN4Z777G4EWd9DgkbysrRAYIYB2vrJ0Rx9EtV8ec9PO
VXpGt2IVNHD6wqir0Whupl2uf5KEtNOzyEKVy6gbI6LCZ230qiEcEVNpg8Px5iiT9KUfbAm+t/zJ
zLExPxa1BN4UyTVQWNdQuPitk+VOfuFo9fmsvpE1FbFKHZurXbIWSpZkia9ZjA2++o43/qt4BiHd
wahU0TbpujZc2fVI24Nc0tTDv2FW7rX/EaVlHAfJ6XK/L23qVnjpgYUGVlyKCN3/aMoWMDVKRXpR
SKM9degTv3s1KfapXhbY+AWEVU8Y+CnP/t+BMulaDTuq0DFeAPxtNczTadbo6wtdviOuKLT0jZZm
0NZjFydtZ1Xlhs73busripx2M9yitIOFPEEtsACRhOrbSwnRJWLoyWqB1Nax0g+faiR03exSu12r
YHCJW1vFZo3zVRC5q1HT2rrS+qbTPDHwnrVVvomphCDT5j+rwdFcFwQy7dvdyEPE+JKNG4AJuLf2
PmRVcs+TERUssXajI7gkIz0I87FI+W0f4oUXzdhEXIAlj4qfW4qWb19cT+zBjZ+DH0ThL+axlWH/
FFP6Yssq9NZ95jKufaQ2U5WLLK6mCt4OcKhpfugltjaCSKW6lRH7iWD1zitT8MgUK3qpfcwpiXCx
DMttjv98Daz2o6sJxNnvojWLkQ+lqlai2wZ1Lk1TrbtYJhmXQUw9VHn5YDPK8SyEUa/+vi98roBs
FwNDS0BmT2DcYTnwQcNdRlZP3w65P8/1nXx58/otaAcLkbXRcljwVK7HYgC43hiCR70N+o0OxCqu
VasI1zwwJMwTrxO82tisbhtTaCqXXns+1ImpZQQbHre9lIy4G9DwNiVhev1oesre9mZhV7AwUWKW
obPVvWdJy0E9xGtVpGs1l3D4NX9JpIuxTUiOWvLjNUec5K9Gus0SfAatfyswq37bnetVzQ1Zihdp
ZDoZuG5seqPJD2pgBTLk4oQkRHupjM9HG9vZlTxKveqP9KO9vna0Nctr6cKp87EGEodhLnfIa/Y/
N/QQp5uyAdOyXd8smi0PoXpO70befpkg+nK+kUG5sOxhT9XqTR4hmESKvZRtLONEmZOMmmwsWfax
4XIv18P8g2Pw5LMwhbxt621NsecqX/2xmYy7R7l2va1fdUF/cWM5Duom+8RyumS4V+kEWqmmUsWE
KLO+7r4q61lV8ArG3BndW2dinSI7k0N5lmFUFWwkFaQSbKtdz2BrKBC/cyPLTW/627PrwzkDPxXR
10Jiz2jS/looDPc4MwQukEJ4iqersSOfpVRmmh2IjXFkzrisIC4BQlUkSs9NnuKYVar1MDGY0BP0
Xee64UInPrwO5WBlvE6hUhdPtep2rqMWxjYwtToQWBJeVrza+94Fneyc0oRrCmZ3ciPzQ63Z7/Ed
dXfhuSSlGWo9BdGW3TBltHZ3GFUcMUM07YKZRN92DKtbgrEngYJSWgZWOi/3qsow2WaTy05dZxt9
fAvJBH2XWENQibGfMF4sTloURE/4wEKyeROq7DT/vvx/mTjll7dukPa0H3u7xaG84gO/pDXSdKIY
MFpTDKpRsbc4PUnSVbvo07OKAwwCpI/jaXeokkGqfSCv+/8Imu8wX3uf9S1wH0F3/9TfoMfWP3IM
6KhWqFR7G8vKAgfXfpEDF6ZPXs0HJwrWRjQXSwa8WSTqjyJn8GYEX873voz8fcwje4ZNfuSQpx6b
3tZELZRYalVn+Z2Onx3KFKieRs0uM2KDr5PNFeG7RhZiUwZb/7O6V3sK0pttXPFcM2/+A+l8pqWi
Z8j+F6Q2Hnzyzlr6aK2xtVzt2y9V/bqAhalgQyi48xC9ALhAzYMp00jMVugPtAcwshUhk77FmGUw
JQsK36VJuZcmiObq1HySYDh/Xu7CKtaTbixN/TaBRHUCqAiDonJAWfx050XCEgL9QLyiSUs6hBwV
MFr1JKy3Bsxt6UWl5rzopvmgYPY4FJ3B3np8J+aC6sMag8GMZAj9SJp4VNzVyL+ZpCsWo0UgJA/9
IpP+SuqKHHedj94lxNhR6yC+6oViBCYNA+DrAzhrivFO2zxM4+kqR3y5jummA7tqznATk+p+92AJ
5C7lv0sQ3aJHauWxo79gTxUwJ9g21PXpPiQUKR+g9uTFwB86NLQWzDrs28fmMFc8fWqf7tOhi5lP
SKxqnoMcTy1PMunDf9VZAEFWE5EVj8T3MiAO4JGNN3L2B1PZfw4hxUYQ6WmXDWmm3fuvGwyE/21E
rqGY+gmz8SeHku/mzKdd/+vqtNNL7VyJs36yAG8t3vxRFJ63dUeTMqve2YkPkNxXDCcFsw9YBj0+
9gUNU1daoDbsh6AlTfnXECDLf4BrpTNAmNekAt9Ku0xqORzo2Srvp5Zcz/vUZMNQtDL7AuW4EV4d
xGWtl9X6y2Aa9U7IKv6RKdrNn80xtbT7BJ6sdnKHyCWM12zJjg0I/dSj5+xOUOe4hfrCbLJnDobA
O1MGWUnZVc5r1sfAkgxBs42lVSnEMLlJcwbvqWs0ruRr2pxkYWsaN9HbFq8R8/+QhknLhrplhx3+
whAspgEdKqmjuBXO5+zEuAIPKumzkwb//jY7N4i/KEiEI3u/icKXEP/OOKrYlJj9TPGwD18+EYfA
3m9BEuFoRHrCLKclG0Wgeyy2NVt+07eTQNcL7wFlu0c74prrJzy/tCo+PA9X/ndNBi+LvphLyqNj
CqS2mVTAIqp6zUBYwEhiVMzRXn4E9bwTy6mSMitGxejMeJb/410o6Xd65DCvtiC4kaOwNshFh7Hw
gL3fQGTtF9Zv1i/Q064d/cOI/J3BbAlIOdUqVduDJolCb0P3vMQx0FK7m47g8ZSMNajrVJRE6oZT
96vRp18zP/OkuZzfGK+CghAo0+Yt+B2A2CuvxYbuP7GHHICnvSOf9IlLcRI5PY4KqMZ/GfGwodwO
+ESjvLYGg4o7sGjTLr4SsmoSE3MB6d9E4RZg15sDptim0K4+MiKdKt8oEq1e5c86Vv1zVzEeaF2s
3f/f26SraQt2kMtvTrtpPeO+9SXYyBfH/yeWdTAZR2ksFzYhmqDg+fSSrJBNsi/KxQcU/RXQjgSH
BZlm+y1js3phRPlhjdKHwfC2jsYKoZf5hnFbhbAxRfaAG8n/Ffraw7SFqeIeschZANNiVgDQV6ab
PKVLn5AkKF9zavAKlw6td0E/b4PTNHBM/IVTrZUtb0y9vid2b39OZ93Wf4jrj3SEA808FPthU0Ng
K14APJYTUZSi7BUwwldw37CGyv9nCApnyWJf4F2fbvntQZTDk4vt4SCbRkXsgCGNNDhnluUoKJd0
Z3N1TjP/lsAP13oa+QGJVzD4zcXq39aajlmn5WzGxLl18/H07mvIb3oCVnD1dB4Y1GxHXtGq3uSQ
6J2fjEpMJ/CT8NZLby1wiM/Uf/9pLWlXLokPbUcrOmvC781Kf0uBa7RKkcTFZZgt64m/QFHH+5rM
R0qLlCkUFgUCi24X5eU0dFJYWQFf/UmmCCVe6tDFfhTK7fWdA0mAFw9xsVdvujhrPQ6Hg4gkyOwi
tylxrOFv6YQB3ybx5MI34Trail9MzhjWAy68a6K+wU0SAXUer+nMSZQZLRLCjnE4KtNkqpStfeOW
dy86w+ALr4/SvVLpKob9iiFnSmFNtLo04EXxNP9SNJTI5oQeCplPWMhCplTmF1vSpUE4E+quo0B6
zELjulq9FgTyswmfk+aiBMmOnuuYQA959P+s4Oz6eMaMb0aXVJizCcASQNXGo4+babKtZEFpIe19
G/BbdRe8ulad9pAAuKv10vZqT4VrhU6oeuKYgeinzKWKsZM/XAl8nopVzHtRjdIP0XTiUkzDwdgU
Lm+k8HFs9adReFE09k//XqA9wmFqUdQBRRUOJCr+VwRA9poAGshldH3cn8HmY7Ti6MZSZ338vjjI
mcYrtP1hYizUFfwcZhFTNMsI/EtO9QDsuxvQdMT6azt1N11Rk12N536l+WC5dlBrm3I1YMcqoGXn
rrpc3NxzUvzljFoHbG6cTN/xOJjY729wO0hBhBHh0VtEdtkrKea9Gc5qlmUtQxoW4yRKDDxOO5lH
WCtag/pTbvUncKjsvMIsEYA9PS8F3ZDbD/mImnlMuQTcGyJ4UUkcNMLYViuBtjK/2dX/Mx1F6NIl
IGbE+JrKVtvXTla+ij7B3aFRVSdtPKa7+jF06riAv0ru30Pq5MxmKyMm6uUh9zd8Xa7f9KX0Oe6x
287iHSeweu2r7gJ3mORn/LgPatA5OPYvgEHCoH1v5j/e/f+3KC3AA07t6zNS82qh5s6kFMa245cP
QZttKofUAr+rpEEPB/k9atpSTsX3qVl1kiB5jtrVkbFTwpvrST5FkfP5CImibdJ6F4TKnes914aa
qyDEfpdE35iHCOtC1b9RuTsc1n52Nc21MzSAIaVlzEd97YDvI+/K0SCZFg0T70szrWGgmtFtBlXE
JiMQIYI7SQR/Q3MvFgEj3TWeuwlf1cL48otegICWW21F/iMe5JC8wowEYLurEd/70myviE3H0cnb
aPe08wcxpRbkp4UiAQfUMgEKxuaHUyNjC5rY+9qA7MIqtz7BC1HxJ32/l//fpomNDJpJhkXXWVzf
JL79uY3IxCU9MilenmM3NPOzq6N1eqGPOH3zQoe2B0//k10zQ3vUsZYOvaFU+AZD+KRTqOJ8zs/7
eVGBDyAWB++s/RL7wdPzqFFTTLQ74RR0qRF++bG7Cj/tJLExg2rMXjNyWAcMutyFHa4T7nLel8WB
YsaexAHpLZpI45xGKImsU5kXYj4yBp43X4CVmV7bwNmiQ3A2CEzP16+NSqhiFpIaj0bS2xOYsnSO
Zba+rm77Xs+lKiZoWj85HcGE/XmnsAAeS0bhQqIxh4lvWjriS7OPNAUQ1QpCm2DA4MYmIXmretV8
KaIrH2suAnLrzt6pZDe5h069ci1gS/hD7iV0CwCCrdsVL65reFAIH6P9dKkNYzJpZmOmltraEnIu
rk71GfzeEy1gAmXV2Ntn2E2FsHKR1E2+zr+CGrJzukgLg2EpWNKaCg6iIBt/eV06qwLy4udOP7EE
S30BJ6YgDqpZx0wJTN18hRCiItvXrRz4JBdIaPpAscCVmad9/y9iBIBgeJAV89mb8R1zrxj/H9lu
280H+70DaYWSPvuOe5Zk5EAhmPBtHsHEY/pHEovHf6+QfXhgMLr9Xc/JwJdlTs+IIsMwHHKbpesq
3jIujXu54xiY6KBjU2CHWCjG5+VivChQkx1xpak+QDLl2FzJQP5SAYk/zZT8p1UsB/Lbqfl03iRZ
gZu6cCWnR47lyqbtBaibfQHxos6+wPVIvEDb2SH33jBhu3pP+zk7RpJJWvb4WQZN1s78u79JGB0G
IC8QoP1QwbBwfdm03J1VQywz8r8MrFCruxEmnX7yqof20AucG82tqTrvhIIJCjBEQrENiN2wzifG
kwEnvRkZd1335rsfWav6BVY9xjuiDNpyl3MDanznMOpSJ5vhijRLvNyBiOD8hQvmkSEBX2napHuv
2+pJzQUFvY+nr48kJME8GQYRVMCX8u+f3iqq4b2maCOQlZW9J8tC7m4+VL8tkBev+6e9rvce5QvV
PfHdmroMzmiIYtINUq0pMPXF8g5KWo+aEp37k/MxkAC9jNyv4X/1gKH5+3T1j2tNVV2BQNv3T+ax
Y4cv0DTwmmzYxJfE9Rr6qk14tbEZyBQvxNUvTmzarFZk256Dgn5IbOEQnjfOMLXhSGSBv1Vub1bO
YJexeapf5ZkZ3qp5+vjatffxhgwWcSAS9TS/9NiQZJZM7YXzDfK2O8G+d22UYzaIScWZROMTBurD
8lubahuXgWFMyKcXdPhlHV+zRPFa99Ucw1Kz6ns2GAfyICarua9s87XlQtVnouwjW7MVCAWg93mJ
b4C2k2z4RE+awN8O5py9UlwVPwnpNOmBRf2YJFGyoKJrRwHAOuO1l1fTP/LPoBxsdU1C1HK8ukwm
QpKUSI2LAmkKuZggA7+J9SyhSUlsew0V01l9WudhXGJketjCgJ4suLBWMz5jVZBPmm984pQmPRlx
OZQgDAPX7Mc2eyzZsvTJ8aqy096LoeUS5QBC92eLkZrjCFycdS+BYEU6JaB7FEKV/6UbUyJeOl3i
5RUccmDiaL5Lgr1vOxOEPWWRSHqYZ6t/cMFs7FwxQDUMgIGia3GiFmgFJZZPoLlPL84E3GeXEzef
kBx6xpoV41aF9dExjsjH3FFOMlK9eaIjIXWRsNRL/iOYLnzffmNv1z+OtX43vWG2pYW7euEfpOuO
uy9/DUBh9M4MzJw1LlK8LXSxYm6sDz0Kuaab/yqHJTAnSNX1g1z9O7eoYO3leIjs+ZMM78d5+XA7
FifVINC3I7pgfPeSMhaH3jxy2gY0M//84QjQzEXJzED2swvf4p6qmp5mtPOzY1bzOalqCnjhUit8
edWR2HeNch76w6nvTA8sRw1TFsdqzcoPw/N/qlA1K5Xy6uqj3Cvy7Sa7/xeKFOehRTAU7Zb0kG2P
bIQGpukpCTtVHU70QGphrbVFMaplksZdPqEIHnpMXQ1XkcNB9f+ICyjh8gxh/tPcrllphGncEAub
JhE4JWdKxiWOboeRBTdgktIc36rg5RDn7KSX368lR0NaHrT+yVoxqcLLeZXw52u2ErYmOc7Z4J00
3qlObr+oy6oP+G3FpBEeF/P8wfCl5zK6hMI2nOJ8yjfyk8kIQX+ByY3RyCpUcjbJX+gkr0KfK7On
up9tnC9DsV4idi7hb9RQ93/ddzcwn/l1tiwU/Eg7lJb37PdWD3fOsCjclQF3MnutPBNhE/HRsly8
Ckn8I0KKYVBeqBcwzwdEuvWHG3xwmUcn5+eB6hmUMl3l12oivwOyPsu/LbSqdZmHzTzcLWN0oeIB
mbF6fxJ/h/L28t1g00PY6jTv1fM8bwEBUsKCi3u7ZPjoBGlBKrxKV2Ftf/kE4eRO7uNYhwc94Zau
TxysENe6po1/g4ONt2vAkXswj2xYtM8vUDZxDyEG+KIhNFnJyLKxDU3bwTLkwNstM4fOg+PcBAeR
Lq77whGoP0mVS5KzT/JtvFtP79ggqB/RMAevaDtUO7nlNSI1V5+etos9h7syCy6xkoHcQzYA45/g
JBDCea8JJ6SMNS6pyrINaB7TwO7a+DICq+zZ97ncADvLgkhdqbIE+tWuiAO3UxH7AGa2NGlVW6Q0
nhAYYd4o7NpYMeTYZHrl3kSuGDb20pnbGengaHj7Sou94xH7GRsCONKpyBxE+ZPZIhuy3ZFqh/IE
AIR1rPaIlt2JJ5JBxpImSu7aNy3HL6heMvUEj/0jIvnzXJAPlUwoZbmnBGz8DvqKEqntuhfAkftu
FPbn0AGZrQli3dhqNwGVuAQm7tlJRNQowNc9VVFGMzi6r72BNLtiBLAfMhHG+o5OWasnbiurYVds
OFsbTSjYo5kum0LhN3/PdRGlJneFhrNL8uD1R/91LuP0t+1Q/JoKWyvdwb1FI3qJmigeFCKPGbQH
9S/i08TfQOM3pIDKQCKrSNTyuWLtS4ngLfoUqv6jsTPeaWh9mj/6Lf67NcPE1/x4Pik881j3pMEJ
DoYNj/PVCKxdPy4eA4ddKAqypwYg1bhGxh+EoRptloPL2KoYNlglPfhtOwI+wOwnk8fKBRkp6I3t
UZw1t65/2EMnqApUtzm8XDIaCVsyWJOVPbv4IKM+RbMPBLsVJHZMLX1KidlB/ZowhPOQ0/J1YgMf
E+MtimjUuXVHojKlXE3pHq31XHhea0SQEEl9mTJCDi4H/+zx31mWVmzFze9sHBxF2a/FAvmsxY8m
rV9kZB43pDnqvcGgJWc4606z/a24McAzlRnC/dhh2wd7jSLN7M92futeB0nfPd+UoerLhyYFezFl
8RQ8Bmja35OVmIhYKmWVauMnA8itQJyqayb1/wU3tvU358gqmvigSIDqjK75+347aXDjtEp0GtoF
GfMeRUtHqSQpvywoJf8nYi/0fTdzh0Gh+sXeYd5ylkvyy6jmnTiFndGybt+r15cQN9mnVaawSG4Z
SNXdGTwI2BkVdvH0WalxRxRFHRhU5UVyuyJZFkJ/ajXqubh137icLXI1nzbdRRz/Pnhr8AzqPIkB
JZ0spAFRBHs3npNH1sgWQBO87HoQEUIi5DE+Vuo52xL4KTDf5OlG1cBLHweXN73jSfbJ0EpOuIf7
zZyRnISjFnphDNpCQALwskbYzz94kvVVCi2yeMVzw/yF5O+m8BF1jMIsOG1zEK/ZEvZ8YNrKEcDb
G16Joe1ezGJekoJGGQoRddT3DDwbzXlL0YXuwRhC7HaF2Pw0x8dezt0YqZbhPd4EXUC49sGIPD2n
6GbREenvvoUm++FhMxfXMQIHtGpupl3jZjWziVZZTLNiefHLVU+nhfL/I8EkDGi00+HO7GLP678Q
MNzetczUq/KzFtf1I57QQ+tG5R4s6KymyrsSZ6kwPBGU2RRbvQ5TOEkQ6l3yaiZNB0AJ1txt1sSs
ltnomWtXJg1J3aHqzC0ANweW548vitfc9YS+4ym+4Wow++eVr2OG1wU+lnF1y/rOca8ejNM55JN2
MOl7j/AuKmON+8ICFF/W9VHsQ8S/arY4OBeaQaCmUJCbBsmmYBtzhHNur6XZU1PzJi0Qa95n1Q2+
uiFdb4NvCJe1O6n5dnerguAjyHFi6aYaY3Ta4YFgdfQwWAALZ+zbV9mp+pw6mFoxnr8rspvQH2TD
nMh8DzCzz1QG0xgqS+vupodhdkwummnoD46dGH18FJcOynkw5FvYGl1SDE8Intq0sr/+YteKG52Q
pk5fAXovy4JIcx2okVPJm4lP6DX0eY6Ks+VEPe7jhWASAX8VZIoZuUJemnn/aUVUSryiUrNS/H2F
/HSLsMFrv5onOoKHintOlacsLZ4PbyGexuiv6WU5pHzcZUC9F/ux1oyzKYywcEitr6WrpxVvuZRz
9IPet9Edb6WtFrV85KYK9bZR/S41SPcRRm3BN445k5NfhCkon3t/u0bXdJ+ciKODqmaxNmzaef+2
+bNulDZ/tlWs4j3P+HiPfJvqWKsAFdt45/jZCNzKjW5pjOBU++AzZDlPJjAbTWyZHlt8OY0JgkWB
6jCsGmeSPkpDvsPPO55dlQIkInmqi5t10PuwU1uChLBBAMhQObbjYwgq12+FsPS3i0Rcq93xv8PN
VMUtfZzlzidjooaiwpRUEefQL+W+XecoPW835bpj1p4LFQ9NTZ1hTaOle0dKqY5Ca12+22GoOGIA
selrX7EPie0z2+jXlBMor2c4dsk3JFm8POqIlL0Lu33KafpHlX7bxFEHKyKrN42iddphOPvcZ9zw
pi2YCegMw2CdGq0KvIlaMHsqVlEhtJ/n8BGZ1BWngW4pwvgzlO7N3Jyw4LcbwMEMt9AJPug7eflS
bwmGzKABbhGb1DjRGEnZLQfytnxb1+L95t1PFIEIOT3K0vbtL+fvXjaQqnfCgJE4krZguK2TkozR
aquNrmHujnPcoo5gY4XGiJw+c1sZ2QPEkFGk0WXjXS0jF1cM4dvHXUomdRP1D7wBjTxHMZkAm4IT
aj5+yAd66tpPg+SV11gbtokHnH4Y2owNPz1Dhz6pf+iD2fyc8QE8zYE6+LU4hj1KSbjnbDs/G4z6
wYLK99hSE6gK6LO1jZzVj/m3H9TTJnlE7xmV/i4mfRT/J8FH5UxCFuWgQV6T0l1PZqrvzNhxN10j
58X5x+nNzveNp+azpPHpKJh8zw8MND4ZhAJ2Z4apFEUmC6FSykGse5VhVPPME6/f4kK6ZsNEXP3m
/PbMfovFtewlRyTGfPVPI8tZYJtog4YC9AS7TqoltB10roqxvBwWHwvWz7AFkDy1Rs+zQhnPUFFg
0uE4M+NPQFoY5eL3obVWbUGQO6jo+TIToqJqpAqUu0205DDoNUI4oHVnZr6i0Iu6x0Fe8c7lX41c
mqlbTNv0e1VK/r04Hndt7H7WudZNkvSLYDGNtdyBHvw5YaiOPuR7i2ermyqUMONJMWYYePa8KM+Q
9ZlNcSvv9LtyL+W+soKjVmX3fAk+NrBSZfalYPUpMEZMtn65otI9fq+IcSM1ldsZ/Mf3fXzkNspP
moz0IvWjc921AK/XZ6goDs3iUcSrYF9ll4NJa5a6qU2Umi6IP26KWVG5b2Nft/jFNHjhPCkHP+XG
HSA0/rDscEsVMFePP1cl9P2rBnsC1p8dJFthJ+BLLvzqAM31Qxn/LgPkgYbpBMDzO/i3U+HZrOqN
v1Q4OuLmHguzPylNnw1/XChBtxZnWd7PgBsY81R8EdbmENwHKZFDoTOlXBJrUqZzdusckiuIwaoJ
ryIhVruTWMJIHztaZYqiGw/UMWxWMLZkZ7b/9EhJ9BYHhvMBd4L3ILHJT+h6Ia4its4xfwxQ0HY9
9e2lEoLptOvoFmwT/M93feNN2Y7pfUAIndqFSsjO2D18cwPK9uYnqlAjFrjgeEKUkKsAhrhnWYke
TIjOFw+NnngqynAcESUaF0FRej9qK3OSTkoWYDtF0PisniW9lG1sivH2wGrXrmkWGZnMAjrPTJjP
bBmYYzuAQeLAuFWL6cGnCmBCnJQkPMW9G/T4Z6vstVrIEaYKDvdxIx14a8ZU25b4NZK/ZDu/eYI/
7Z75t5AzRzTSWWxOzmGKYXCezjT+Pwku6SzIt7zFV+IMMIxJ+X500FL5tt0siPVwOEFMuUo7K+nF
2zpQbIZvGo3OMby/dKiWgMc6egFmNpSRviiGuheaQfOZcI7TsWfPTeyYq35cp8A7uk/M3I14QYCj
HK2768qXMozAaYbfeAMh9YzLRQZRv/Lnwff3fQ99g2vGzO0ku0mfCgeT9Ru8x6IwC4WIXAgJvE9x
ZIJiSQ7KCGvlKREhjtb8kFTG/LpomSfO3b0c+ahB+I6eP+RBjG5d0uIy4V6HqJYCA9TB6SJj+NXV
tZrqez5stqLDWdG+KEg8iVBDudfUpVoiA4NkWyYBBcC0c1M+12bddi/Lwac8zPZ8TwuWKS+pysD0
650W9YUKqU1W5Wf0iGCgU63PX0u9/XkXuu0aXejxclfU/So4ecaKFUx8VsuCNfOpBCLQffj8uWkp
mmucCKsYsgsMA5PFSIOFJka628wCuwom8nzLmvqw9V1BS1BVomoJMp8NUByQTz/k7NB3kFl6us4t
fV7d9U1nHqnAXIXh+YBJVy+Nl8R/2wLeAXdi0hUpGP4C41aWGXr0gv8P+KlB5wDhlfGC3D0yJxdB
LG3dZQ0Mc7jo2mML504BAZ0lAGF5fHSNPiH0LCjgJgtUwspiG+M0kcjTUKuxuZaUYcZ6+cUQ8+Ki
f4Qpa/7ctyYy+eCoND3evxogcMS07+wZoqOxCD+XIOxmrkN4ss2SyTCj1YDEzrxr8D9YxnVyFgjl
HiqJ/eLUHWUuMnq9Q0bvHHjMsx35InBF13XH13P3J6zVCSoTZdgXmQwPRa6kEm6gqZX9/rMGI7oP
9vWw9rg3mQSEZpHJG71vPN5xxLXo2AmkFaHasdYKy7a/6/c97fYSBKh3sCw9EoeP29X+FyNuzIt7
MD1JKkM11Kn/zBZh3LuvyBchkPmJMsdef6aBr6poLu+y5LmychV9zK1oup3jP85PE+dzFuwxRdG9
O26n4S/q7LncBF9dJ4K9+WcAEFrCKs6qE/GUf6MGiJdGTDPE2ffMN4pjjhHSo87ms8iXgLG5OpEy
Bo6CuuVXxAK5uM5owLEEHhjUNk9ktkv1I117WP/yCfp4oZVItK7oe02V5YKe/+M1H+wFdVDyGZ+B
g/ON7A20cY6wdRf6RHzw3NAP3qiv+H+UTAEPXmzrbc5Btgg4iK7Bjk82J3oPdZO1DITPdB/KIkuQ
PiR1vtJ5iwGKdqlNcDZvAJ0cgkbkYOyX4CpTESt4QXTBlLHsZw2abuXnqtqilM0dghmlU6mQeKbQ
cl8AGDlayLCsY6/gsUh1x3WqVUUBESnvP643NeA9OpLvzlu5B73qBi9tKkQDQgyfNFCJEPgHp0MX
FmbI+pwbTVB/QCTG/MMRXW+sqD1fWgtDmGoSZ1bMfg8p6nR1/W2DljCTJBdl4i4ow6INIKTLSUTK
jEHh5kABou9NU65slIMUSfwCOFa17yuineqIzXyRt2NvFgu+ap7qkLbZdefu5jltLEL/qjJxv0hv
8IPZjQjyorvM70Ocsn/WFFbHdZwxZeUPJ/1GOgxwJlhbby+Dg/QU9HG+P820Jf+NW3q4Z4O3XgyD
aNDzkhkNtjxoCTb59MTGQL4KePh8AvgzlyyGN4suwHReupaKbkHsuCj89sGyyQ1gCDuVy8VW1IOv
Ebs4XnWzbLHpDtE6lOIwhSlA+GB5qWeHM3+s5LVMNPjcvkhmknVKZjJ6FfKxs2YzQYeOlIXhGkH6
whnPH821mhGmqJN8NenQWh+L1Wp26c3tUOSHXGkTM0Jusjx6Z+8QmJ+bmDFroYY2EfA6YxhIi15k
xOfasap0/PmLGM4dHelSMoo7npbu0gOafNnuHYaWa/5TbJNCcCePq+XN0Lp/A57wmwLUJ3uwUFxA
l3AL6MtKsFCjC1VM068314cJqUilbNS7exIzeb/C7uDo58czQTOh4S3K5f0MEn6gO/TEvG/i1yoI
tgInwMc32vwiKrjMr+5qK2BX/+V3sJmUQcGINJeAgKAg9S0FaayNjPCtWcHeCIgxfsalJ2XSYJHk
6AJgO0EvDXcFhudssbloD+B56vrm1I0xVtE5ZnpNwSBe6CxkPNFnsoIV4NBCiowPmST1AC/hNY0k
LtFKaB/is4trRoDgBJkfcXBPMLMevCEj+jC3aSZdxiF8P2l/Mglu6m/bLXLfZhWsRafiZnImPNO9
wYcJ6CC3EhOYbaPqdNtiUmmN4Al3Oh8juc/C+lCgt6bXNpp/odvHdbWnUHH/N4bp3Teeb2RsXoWP
KqQ443M/NecmSHmCGevLUiiBm/agQ4gT+67/in7rnkPXQDj8iTbvnq/tUNBbFo2ToD2tiosWRET7
AAROiLy1Axb74Id7BcsEH4bMdJpn8XYWJusS8++LcSlTIfMBmNTbYi78DMYKLWBAmbWUlUmMiDrN
mqO8EX8dai6bBFnNkcrtCpxqOQHexFIL1OsK2XFvGgnpkP+coo4xaGfAMhsg2h4JThsQwJIFmXvb
jE0qe+bkh+1unq4Kr0NWZJ8rE8CV1oQnDG/09VwxuqFzlcTtpQRG7TAZ8I+ZeTvwDQl6yZyh4dCK
5ZkXdKUGnkjnzwfPm2XFavqgsfCj23rz6YXtnv6OumNiRuRqi9X4kjaA+1e1diegulUq9cCfM/pI
sd4KrHu3T049lL18W65Rynggs6O5o4Po1KQahNMXVPXBQxFikyW5ny6iuFexmlNkHXoWUh4xx+T9
Bezj9pXxDhP+9osNGZdvB5tRxpqSeDPuyR5udJcZ/TE13851J1GfaUPdc9HvATvyYMFleAcdAaWr
GlXdIsMbAcm9S93Q7eqqEa9CE19Foiu/dJaND4uW7AdaEQxxsPr97O7RuNnJogKIVeiO9RJbEnfK
gNeoHFtFYSFs3TBp3MWDD2wMCii8t3oHPwzobyx7GEDK1zZ3yvMKWrq8Z+rQ5Danw6Shb9eYnrit
Vu7hiIVT1XWPATfi2ek=
`pragma protect end_protected
