// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GphJs9IqaKGvsm3w4uDCe8KKOVGstNwnxZeQ7LgKTcG5snk47VU/YojfLlR6vGhZ
qI0i+hIUtV/hIcL2ViZni7bO5zofNqZxS5miiree0gAol1L5BrBKsGAE6vcX8cqD
b34KvXNLrmsmdtZA2AQXoPfQtH4OsVvYPcgGsiNMQ2s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
D1ACEXf7KwjO0JiSOPXzealmmC6JDdFktLugqeTLxYS3s9DrBxFIJF7DwELckgw6
7OY/LIqsuMVZ+rhf40lqORowF8gKU1fEJ7DUHJaZdqVdYZaUBJtJRY/QpNgtN/ip
SXKgu2HEFbZtQ89e70dmn8cIwumH00m340wpqkSXZvw+sPn971xvDhgoPnLcTtCA
ERnGy4fwI1MNfMiKCTJj+Bdv8hx19/CehhBT97n0J93N82DIVWMyWXrxUMl7LL0y
IQMpOOi3ALDSEGzXg89zRYY41Ts779MW5e0X1DI8IkhST2PBXI6lqckDzwzPCBVc
GNTY3Lto2Ja7dh/ynGntqvN29qw6oi3VSMDFq3p0y7/JzA6vojkhRK5RoJ9EP1JX
5f7+RNc4h+DvbvmNIho6NDfMeXBIbwoSO5iC/WMGGUhmFMmal7osoq9SvVCMngV6
Ypsz8rr3HrVDIRUAxx4HvsebzuS35zyEDBeHBTvk3UhAEO1YyLFO9GoofgKQL0ZY
21tbfieUO+J6nLFf84w1dNDTxqLGH12OrED6lcK+k5AFn81uQvR3tfAkY2WEH82m
me6adKxntAXRuU3tMBnUalBOQQ4KI2ibOyx6/YezW365GBBWaU7vSkn3QgDWu+6b
Eo1IHoT4sfkKHc7UJqkfDPqapu1pPIssvRHVQg80y5ianfLldWvdL3+CDCc7R6J7
UFrpBDjaRd86N4Q9L7y3NYlRl+X22mMuArB8fCojKfmPyksqLM/+OHkvZklhY4iv
t73jlNLpxWUeu4tiC5pgEwLgduqUkMPi7FvgesR8mco8/BmPB9QIiagkc4ov+tla
Mkc/dFSckpMjsV71G1RF5hQSgyhpaIubbbKwd3XJ8pHQUfwnJb/pLMq/54SkRnHt
gBVOgiAkU3R9KWVXwczj49MMDyfYyFX1dYPKYNmn+Y3AqKRr0aLBoEeiz61T5azF
oNrkdUif+MzX3xzDfXZEmHOsBW1C0EIzXAdbk0GU+82sGEAf0HduJRiD7wBS8y4/
cEJpXqz3qoHdp+3TZET9UF12qfRJDdy01uBnYXjdcCD8wSnpPD3BfMIO5VyDY+1J
5AzoZsXQ4G0gutLJUjQT6hgING4v1VGRbZQr2abpAgrDOzWnhCqiwx79V4VJOSQx
1W+lzjRQ2lUqkJse3sv9iL3LNF81UJw6pJAW1VjH6Ce8N6fq4hZRH5bt0iAcJCxq
yFKcVSNJ3LGAZAKwRc5zfuU/g9MPiQKtddc7x6FFF0f1+e/qg+5EatAKfyN2eohC
O1r+i5BGpOuWSoVHh7rY6ZwebY0qJ3pdeQG4vDdlWK9EyB5fMCphDeSD+7yCoLAM
R3A0Vduz1R6bARbJTvVNqR0/AM+o3WkQMnlzGvPOkYSlESXx1646f2VV8vM8/MAn
GeUg97xrD3ldF8jU5bYiJMIm42lcjSfylQ/SGVAIAHjZczSYAbBKroPX36e0CNFw
V/265PYySJQJVA2fRDxuu/GDOOqETDZRNyHtUabHFs3fmNa+GL5KYhdfNoqyHQpw
OOheP4rWvXigQb2YdwF0CrZXvelhcdA3WNlEMUMac45GYJqCW/bvcrEITqxnCPoI
thdkxrIkOfghiDKje8imXdAY1cgbztZBNLIHMsHk89P3pPqyYIG91QQdXcGwI6r6
DXXAVaZduOmnbHMuyYXAs7KFsX1sknxyvcxMOvJvorwhz4082OGOHfvLeciT+r6l
AtUW9f1w+JQ79RBXOwqWE+gVAQnoahfsygpw6XTRQA6cfWDpI7RJ90UXF/lhX9Vb
N+/Hyb8h9WYIlF1+UBewdKMsV1xL074dQbuubAr6mJxpafcMGf++a7mGwW3wpuUT
7XeBIWHkdDs0PLxOPsRZx3jJF01wr+rPpExieKbixFdzqERukOFtMcvQWPrOmrR/
NWMit4CDb07yK/Cm/mRaSDp/af2Bfbum2hoIg2SpziSOHMGGHJofFPT41Coy9zLa
o1WD6a95ZatMpIe9THu2+cft0d2UiwS+TA8GWU0Im67HV3yhBZY6V3Ngirp3gO0w
/0HvnaBHo+X5LbGOLG/RdLqQcc9x+6DtoBgNl0UPfKjofocH/dW/8kK4VHcDhmuO
nU2LXE7RqW8KaNgWDN6MT76Kkde+5+kBVtxG4ZUrUpKGL4gsFqSozXVRQBejWAnp
JVk0LplaqV4QaxbbGIvtGjZNZOKHEfLJnmtnpzaNu/LfGRq+Nih8D/Flq6PlBt8O
fxLGm6T68YeZELY7J8LeGiMLQz80U6PWbymrwR6i28giLHqs+DnoU4PZEUwhLB4Q
RkQjObJ6wEh5y1y3D3/Hqhifp+PVbeLx7v6h15lEqJYyl/fIhJFjgQO5qd1magh5
S1rYJzljk/ZCO5XdyUUPfp96w9qHESSVEBKJkidcGTpkpCVXlcGlfQvKEip5qs4W
utBV5mSjsiYuHFx6ikWP66CGTgL+cDZ+QqbXTXcpCAU4Km7xojLowwQPZ3i9M0q1
w3gKaPVxyrD3sqBWXFf+T3Bt5M1jamMC96RTQ1nusMZ7OW8p6loGQiJK4aRbXoKB
eZth7QZICTdZKD2vaL8qSYnuPFcM6GgBGUTauDiuh7BKktmDrV1O5k/g9i8RcFeN
2ulNXEXKGbhckUwnrLym47ilwyOgg4tYolcS2PXJB+8QX3tck8iDIqC8jTbdTvg9
lPok7UnF9nbs9/cQywWOXzs/1OQFaMN2sqTMVuK4ssK9ajWGyQJmJFQlXoaBZNsa
GBMj59QSB9cvVdvdeBfp4/KYXvErR4NS6Kz5iyiYJ82vh3+T8aIswboqexxvswCb
RgUiHgiR1a7mBy4QdWMcvA5UwKR2EI50IysumL3ZXseqR5GKsjB+G8c5QVGfcwco
DbLYh56Z8Cr3uY6k8JStrvdqdQogDcdAUFE6cDo659mYN8IVd58n8/GIfVe41P/g
jo1zLPxrQgNdVv+pOeWKhNrSVfQS7rdx1VF7HEDd+FtGV/aaA2h76BIetWqcXPkq
pRTyIp2wovG5sYfAyW57TZ2pTg4xDGA+g1sjXiGdfl+QHzZUpTLlwPLPDIp2/RXj
7JaVlGles0fudKtqg8Q3skAoyk13Y3GZZguwizkuo/C+t14N1jXFJj8URhgtD2DQ
wN/ptDjFLkph1uyocn4FaQ4MVoqTigDM1pzxGNXsSdaiUXGSkX/p6/3v5uAyjTQV
i+DxAX2hO3AH3Lxhq6zudYdSu/chnmZWk+hFhfLdOzSI8ce5A8reyEV0kZdwWxMD
bIB8xMPSTc1fItWNhT+e7Gys8SEq5lIF/LKWz6b/3gaM7AP1pRgL+31kiJALJdrb
YWUUzzSpPdIi6IvheO6Ms6aB6aHAorxQct/BGA3NTp1pfwkYMDbUJyp3vvV4JrUA
5uT+0kVk+VqSRJo4kEpuHUTg8A9ubpiqOWxjEomu4qXFTmq+H8F68RiWMkoKscDV
u6NAbJJmemJHct1XpbO6fK/MRMHI/3m96n3HKr+6yJr8Oti+IcuTU46Ti3mbbNOa
xFhNKdqUlazrSFgQLyCI5T0+6qVOrlZQEwpAzzcPtLusYnRGaMUbKNJavp9zC9m+
kQu48a9vPpk4JNv5V7+qX5MCp0OeSB0LW0XhP0GEIDHJYbbMuHFIPGyZoHS2zaqL
siPR1/TORWqSzQ2D7P3vL7aG8tSjgV5obgnXipqRAz/Q5+zLjFh4EAc+g6PgwSMv
uCuSHhw1wJxOSEQn//rl2gHviJkV9YQGGLM+zaW3p1JkpxsZba1isdDtjXYZXj99
zxsUFi2qPIG7a+12x4mjkBkhqUKo61PAMgbxPvlnNUC49eHK6peYwWS9Ideti81J
CUhm5BdrvWXvxoxczowM6LVUDrsM6MFNlu6vFlcFgAwx0OpNRiou313y6lJjr6xY
OO+C4h7oftiMwY97eAyXe9gMXdzEG3clOF7R/KTnoIEdy5dKseGSIhoGsqZrPMmE
mWtRqYLLQQSc3BZJgnNtD9sTN7UZmnOXhYV2VdUlbqaT4YKYFqf/nOUr0Fp/REdG
YEQGZXrOrn5pg1MkgxFunFO8Ijr0k/OekxsWdejaKrS5g6xRwIzWC3XakIW9TZEB
4mjoCeYKYJDm0JiF4VfpC8Gk/odiPqdMlEhQZsM/F2dv3CuUo4yD7QWGLIpXy2Hh
oue0om/AbfzWTj5jB3fMjkBZM6psJlaE4wCQ9aehxhYAe1vbjkJX5wVLPLgfmnSn
W0zlLrxYsNAwwwgyUHlW4Hq3ZUzqSFEeQAiTzh8DDI75HmTbUs8IHN04HbSJ0QOJ
GMZh+NP6C+sM03TuX0gQt6dAuMFVrMpX31tB3dsJ9PiJV9ITlqpE0GiU5mQlanEk
tioXDBzujmalO7W+kyup0Q==
`pragma protect end_protected
