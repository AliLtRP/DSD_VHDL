// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OGIz36kbb2uZSYIeJVIqeF8vduUwKEyDvSpNfHYNiAqL3hxOkRWHBdIXS5HykcdG
2Ilv1xNeOsObozMxnCncPOaKWT8lubJE56UbZSRzYYLJnmHW1tnVq/cV41Z8lMv0
p5Ypqs0LaaHVFdt/GB5bYU69Brn5kTKCm32FCt0QhUo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7488)
iN1zQUb6Cjxv9qcsWleidsuM3lCZY8AmnolathsNtBiBzkaVIMylUPz+RsnG7CD5
YDNLNxiTDxzs/VGwu9QVBQeJUPUudc6sAP0VZR4sK8wnF8rfdb1oqM961ICTpCMt
9MTPMH3hnllE8SSJVA2q0qENgKGmyPDlO/I+E4HiXX5FStHb+wfTM19D0gt0T+9r
TClbAhU9tWr9oitMqg0Igl9aEZeroPrWqHd2UzzE0RzyvQHqsoTlIzqUaO+oToNG
bQ1wAFY2KMAyA17ryvlykHCAm0/kPHzKsYJ4EAxXWtOy1w1uMV9tBhIpVJKjDh1d
u5TiIpXemeKg1ubF6xkz054Ui+eU0J8fwnAYTzRXnV/+u9CU28VkIVnOKF+aZBo4
zYLW/It8UhFeVISVme9Jhr67g5evqhUwFkmGgp/46UBqJweueBqzD6wikuoZG62y
mFkhAs9b+RePFjAtnFK7MUUz0nUr+85oPpRT9w0wCBLLlzf0i7oLZ28VvU0XQPRE
dFa4AcMLneHAq4oKOfTB8vkdFD6qBd+BAIUF3LNlbKdZZ3xjw1OoXFyUL06uO5B+
DqzrJLpxop5de9JWDtTma5Zd1lSrSXK3Va+foyOaWT9brm/xBUAI1w0+ewJf2JKY
24ft4aDJdTvcTAXytlqqO3qDvmj8uzjmrBVKFhzdvyUCT1oZi9WzonoMhMqVKdrM
QMrEpeHpomerqVgKcTb9xlLRx5i0Yz4BGkb8OH39SrIM63JSVadaxbdtycsqOI95
XTNBz6tJxRAeWn8yQxaP56V+l0mYkdV6Ugl2pdqKKFsVzqBzdGRUBKHMv7Y4j3Z+
ncRQIXLUWf72RrV0h7pyL2vfxKWdibO5ljznIDw3LKfdZe5x8sMPVeHOcT+u90Y2
BD98JqNyW4BJ65KvEeU/osJF5wE5Dxq0VIK8IbU/9f1WW1Guz9UB2bVM7uM5bfNP
nLq6P4NGgwxH4oVB467NlUHUFxMlJweYznx1ZjcTCWSUosg4Z9vUOViKzoDNRGsi
LEz9WZhYYrWMCFVUoLOj+03RM9NKv2CuCOVsnPRHSFUZC6ILaMZOOeezYk+SecMG
j9OgBhBhU+OgHn9xat9i4vA0JGLdWN2Mrrf2DSzrTfVUgDTgoqT98tG99xINi5dg
aqNKWRMJN8XSLPyt9YTAhB1HAGlqZZVAU8yNO392XETcrSfj0dH7cGbybI1Q2uq3
0Dorz/KAuhEemwdQcrVR7NEfkancJTNncAf1zmkH+wuCmjM9RjXsBJRx3VdoZUk6
GbCBXSXLlXoUe4yDxv5UIjMC8/GPlrZM74Tu1kX76BixiGbm4/dOe2TkQeMuIqJf
AAv7dPnso4IcEBLOeP4E98UqYymrK6T2yQ5Ri5FHVCcKAKwps1B4Q7bEmGN4vLZJ
VPaqZrJoFgJTHvC0kZySuV2Mfrc/wkqteaCQCESvR4FGIzrhHRY1nG4ntimFz8uM
Cr6Q0UB7WkkkF6k4zPQV03HFXHDpvxYvYLF6MHoJWVuUGut9/60qC1ilPn3bz8Tq
2tSetl6Rcebd4aKOQlCqy0ZuWNv8ma8NOzS77wbXGvq14QNEZYUZ0ltA4ozGkJXI
E2mBbm08RHHZcfQcpOo2KdsOhFjy7tlBFgPR73YRfWzy8u9lJ5Ip7HbPUjX6GBIN
2WHzIK1nd9RnEzlj6x2ooP2jFyVeG5DoWIlmg26FeYEsBUykcD6qIC+e65moYGby
Z+A+5XNIS2Vp+om93uvfVBl44gY89fOedmlq1KH1vCDJ/50PbVjpQ5jSCTV3wdmv
8AJEccqpfnOIrZwu7GG+yf3y0jfax0kHwina5sC8T3T17H6/i7LTE5tmLL6RTDBW
v22n045HZS3Ag7sGwZ83B5jwnFq3jcgBLzXs0WmGkXyN20OtTHs3yPQsDRN3VmZT
2xlwbwBPx8IQ+a3YrdyVD7Dfq0jPLWdEtlq3cix28G/6zH2LMap9TiGD+39Bgn7C
bTqVj83JdxSPVz0dBq2ElPWalLME462cs7xbGX1jYfH5i2o4M0JZyx3VQqxaSvks
h9INpJP0YFT6VQli4ABkvoTvf4zzjhWK6pGceU7aYaVk82zV/bdVXtCyDM8vYw3/
9GHm2aCax7RJCmIXluq1zcU4ZqYYpxuOcm4pPAx1qMHO1pTfsPTSJd1aCbiPyA1a
n6B84Fcfl8rtitkhYeqUtJc++ru12e0vkMrGnmFj6VPZxoJJibGnNfAGswb90lXA
Dr4+TLn88SOXBt1YyKjqY+aXNRPQHvgSPDl8juUY25uKRuftUWMh8frAkElu2uh9
9QVyC0cDgVednzmc6dlm+hUVX9VFDqmi7PKcYZVFnjx/hnNfrLJffVRw+OCxv+sv
iihXrTisCSkRXgv4Ee/P0GYyBY9xB1QyOVGobyKg7kwb21B6rH1emwetYVQ1NrYY
fVEbuyubq+FqSRCOCgJ5f6uHAEjInm9/AuRFhJYF0jAbQBt7pSrNx54ZU42HIvsb
kgQUvfd8p2PY3uwZptwL6Gd4bD2LHHS3dURuR9bGHbEX+iXK+4oBHmS0NF2qFDdc
/VpiUaQpLw8opSo2oi0LKwiwcYTm0onoshirkgOLkVU7mEad1r2WP7ueIjSiBQDB
vzus6Q146lTA77j0Es1axkPBkiCFMRyQwQQgkS3oYqAWhn4sOfMchh/9GtJvk+JY
hRFY8Rdjtki3mkoSXM71C7Hpw1ggHdJHmMOdpXNTUHTP8XK7NICoet2utQXZZdFX
MjjRMt1aRRrTNkeiXoZzCWfJx6RsZaWOD5RsQzZbrXTPZ/4heBG+nirCFGbw61Ms
OzVuO8nUeD0JGHDUtiRip98xCjp9276ulOOrXjZfTg+ipvm7h2L/ihyI7uGInQVd
GPGfS0VJoL4DVPoFZrzuk017430lXlzGwhuNUHjJ/2+VIMgnT9zUl1+MMcT3TQgm
c0IlClPUYKXwBKuqFW2KQm5kcy7loengo807zLyWdk0Va4mI+lUX1FRO6FcVmz3z
0j0c8Z/fvdgYCdYRxc4U78PrKBfkITBLFk8ZjcbH4uvgV3Dr9o71gp4s1axVZrTQ
AazRRraDE5uJEPYdamNRFl3r9d3NpAsCBJAd9ssautToHsua19t8mU7VzGL/mvPR
JLPGfKe6hRkVylXmm8j3cdaupYeWANJVzBNlDK/4ovy6VlDG2MrttCk+mV6Xbr00
PCF4vY8B63Zh76RPbDQh3P/IbYVH7iH/s5mbezItAY796PIfoOP/oVX67Z35wZ3i
IbwX0qyI9k7z5qwn3kxqbBwsTs3SFm+9iE2ntsu2pX1Gw2kei3jFI3n60BTsSYJp
Ot1iIyOkGwDC3T5wnJ8ErcIac83b6h9luYHQVS4lO03pQXW4PHdPgSAgcRRg3+m6
gDmJqjc0dkUY/ZJZt5/tAj9/6jLAvjMde44jEaoo0mBAKW3QPuFdxpVJ97lp2y11
Ud+/BWApBimCMknB2gPNZZjYKfa4U+ejpO+ToGdzLdj23UMSToY4xw2XOUQRtXsT
Yx/bAElIDoXiwlqiPGEbXBxtZHnMjQFe44W2ez1txlfmmcm2CgCHu4pJznXnjvoA
pgRxi/Fkla2sm2oVEv+4Wop6ZRH7b0bSfTnUhoNW261gR6FF1L+x/IBpHDGrR/YY
kkl++2sMD/T745n/yNW9+WPutvrjjQeODhW5PT2Xjp6mPwYBtTNLR9gLLcrfRUzb
odMx0knWG7g9SP0MxB7k9CkPM0fzAQ9ALKTfEMflIqn5/r0PAxpMSen7oOnWtt1g
MPKFiqzh/7DYqnqOZlTkN0QgqtXXV/8bBYgJycQ9HhW3HY5DUlXzL97Quf/DLup4
d4JQDBNpIfxk/p2jezXY1tsBMilBd73conRSGtjwz5vG7iYduRDXoJx/4Xo1OOfA
cd3IyfRO2FMrnCnme8855y9cUfoePE5gNa/lsEIKwxAriNDQZPd1wNrpRDKakXV7
PV2xFGzf1ql8V4/9m5JhhQvc20lq0WlSnxf3hx2YJPfKnf7DnXps1shbKzuCemhc
Qw9WipROXroamEBkom1+SKfiOdq8mVcRERvbCg9Yx/IsTamMzfqooXcUsJ4XqhyR
u2pJ3c+W3Wtr9XjfyrYtNdKzyP0PcVJVHH6/8xKwRh1/VOQUehomzersamuxMfLC
v+m7VU737gbFXVidTXJFh+qNnFlJC6JWniSrlKLmyqTH2OLDpvYNVsHGM+PI1Vl9
dnE04J1whUkB9PiW267JO9atJ95PS6udI+5TN+3Hjb/Re7EUm9QhRlvjvzkMBROo
jsFdIhgrDwDLBhq8tenD57nAfrBv3CLEH2AqkVrFW/u+caJRGkrGgroWNcPjm/4L
VgCeQs5VxaltWYCcUw5WYmeRtLjIKGYWkPqpHY12sA75uuEfTJk0o7NcaWjUSUAz
W80lBEMSkhixCekotVvnNIa7jvpQUiX2f1cKz6C+0e5hs5W/OszN2IIkIZjY3dgC
c2M22TkAKSORfQd4SmOD4satrLod+56eroNbgS/aAxs0v4J/I48GNmw+LC0pVHIk
vP1uhWQlPKVQwu2hgcWhrEryPuAzbP8CkHLxxVsBnoA+5z0HKthoof/4Ap7V5QZq
8Wc+cCeBE0BJrBW1nb3OFB0B14IMxlPlBJ7+1UaYMtE+CAlMHJg+8wfBZXQmPts1
GmfAd2LBah7uUkWpvUcBL0Rax3Wz1QZt7xg5+kE85uW+dODSk3+9bMhCZcsX0kZW
M1LSFNkc/GlSB/JZAmL7n/aKYh+zRAcRUmf8yQVJV3HLd1LJV9JPKtPprrSfVngE
JIkuin+TbPFez+nW/CZkKCsX0+lupDXTcqckZtdnCFU/HFdq2OxSnhy9z6Sitjfg
0vG/Y3e9+vtrg+9G2vq0+dZvnScXfBmfk0SPVUa7rzIthizRJV/sA/03S26Xn6dL
vgRlz4oPZIFW602ofNQC5rVzud38n1mufy4KD4DszVyk0qt2mSL8hnwq8E30mavM
DvqsiNFe0CkfxHNJiGDZEkhr2CDQ2tialyqAHd4lBI3jjGY23nb6nJc8BTgMMxzi
kL6fRIzsJ+71VgMe6YdagTSAvskMunRpc0ayg3++ZuZXkWrc2lBsA5Ih278+4G+O
hKL0hjjipmPVFtpd+KEsMgccZkmVTyM4Bv3G0RJRd0K/OMIxDOEckoFfKymvLfs0
O8+WfHQzFvYc+YNnqRaqUl1ezJv51pjDfLEqXQEK4O6c+JnIHpoox/iWuHbUStho
90aBV+Xjj0ZcZUfCmmIoHlXBozoG4wrflLha4jiUDx0TEcwhxzDH0kiv9/vSDd7Q
t+ssscHJzWX3lPItIxmQoguLZRrLBbkjfOAGjG30kA3UpQ3VzFTWHbGo28hAjC5V
Lve5Z3Al9XvpQeXlr4p3YeYB3b1t4Pz2Y5imAdLtXHjnh969ydoagfZquZKvNeLp
mWGXdhx9clBJ5TdTiOofBczX0fPKqc2ccmL9FmjK29H7d8iYJGxznoph3eYd8Xuj
pZ2jj7ONuJCxB3oub8cHIJz/icxqGgkTj5AJDyNTLu2C7LTLEwvdv2UPSJ0s3aB7
wY2dj4IL8QHO/6CJG2zctt2IABxOo2tP5GoHDQDc8lpSYuF5nUXToCn7m6xEtjRq
EW6RcFxRQ+LmK6WDE93RhUQn7+gtfZa3ejSp20zUMRtEuRQwivZ77CmIpZvLW6AD
4LAQDV3kkUE9odj6IWV3xW2ntf9gPc/wiB/MHNMxyELsGfbWgL2Qt/f/73/RDbBh
RWsVe36kDuLTECsSnsdwhcwbZ+oUjuVSWNf+UBZSf7ZZkgPQMlBgyDIy2w+sdeUF
UxhH13Ygcg+hTEqejdK+C5+9sqZcp4C60LSGIKnNhJe5zTlPWHevP4c2vZDuD+yt
5Kff7v/5mg3h0Gz2eU7KBUtCc9BAbIOlDbQwFIbeQi69WcHKlBPY15HBKhhW368k
bkwNYqYTkabP0n0d/HP7kLnB8pY88I98VUd2rqlRsZxFmZDaBDjRjC3TXvVZBtdb
rWSsIJgXvvqF9xuGjaa0od+zyLf5vLo5N/cs61zRby0dP6+56yWdtOuiQNWoxjPr
U4uRBSXJydIvcSPo+YxDc0i4FffbdjwnZjPEPhultcPHdd4XmL9hPdZX1uD7efeD
nJTFVguuDPD2Rppgg7H/nmXaX/abJDMwmDANQdyrllNTGWf2CHsBm45X0HXLVL7l
IFKM7MIoWdJJe0yFvaBjsXYNPJ6Z55uYgpTK59a9/TwPWXwAOwD+OBAmzt0Unuf0
1vW6ONz1ugDeuYZXAS+qAqKooP/hekwwhwJZd+LcSr8VkycWu7OM1D7LKeqyvFmS
j0hvuKgARHH4U7lIak3KsSQGyIiY1Mgmf4QxMkJXr4QshBKjPqG1UmE/mW9Dtj0i
KAnoVrTWD6kJMqd730TCROembwAff7pO0DXfAiGLzXDMYvVs5iU/lcznfH44mikT
G5dMUfDc9AjJj1fZA2xgiJDYFv5cqPw9xBWE/NEfpy5FU5QoyyYMKXAdtOAB6jTH
tXrqt0/erVPvwjZBty2g3PJiF97PEkASHGpAtn8NVFUo4BPj4dfum92sYa/4dmUA
U8NN836XHLSNLXGSFsZl7mxl2Nk3U+JTvKu8od68Owk433wYhaTsWJGebDB/PuO0
jpV4Jbc7kMmqoA2IVERVwRg5w7zjYh1H96KKMeF7f3AQonNBbrEiNu2ohDUA8XkC
QOEN9QyWTDRXCQkc1VUEcLUee/cAJhf94uxdt3X2a3e1/UVYrSO21qOuNeQXAqyQ
iKgNVpq5wmuQHejflnORO0B6l3Zo9IOzlaIawGNuKG/xd4gujNzeg63BfEcCRKPG
sLvoaqFUpWTUQiEnTkofih/wuXS9hB+wzLB+dP+UtWdPTURdDKdwWAHf/F4u0VQ7
LYRegqrdqsRMnSz6Y0ixWTRNNSrVZ3+VEhfGufWSBx3iEXt9YfOqL3pmZEpc/Q4i
zqv51YxxH6ZJO1+P7BsFCVen6rGi9lT0r4oTaNCbjmxEr5mhXuRirbRlTZgubuuc
ZIiB6cCkpC4gGFBJK5blOA7JDFqfVUeCny8eb5vUPbOq+siu53X3o4b3Wijwf/Ph
FUqbDlZGknrB2W/NCBdLX5zay3CIDSbpKmiB2LCPCqknm9GJ4b43cs0BbRH+YAXG
0V/zpLaLjMCrnOhq6P/ZUtNwpUb/EM+jrx/47PaT2zAIf3AQT/ZYa4XCvfpBDteF
WEp4P3+SOasZUxhftejTLKKHHSS9Fx5UR1U6gPx3HKhIMj5WLDiFbv8GvPZKbVe2
ceMlHcGdbacNz/Xhr2xQTWE5YMAbSIK1w7SSzjKV1anlF9EvnylpRUEs0m9SX94/
Ntmp6wEWEvazgtiEQvIGkSu2N1Rb4T83bA0GiJb39OKIX9qkMpogzlM391WTb475
ysN3DsKvl7/PRiBfCExSW488jf+i+Puabv8SwcPwz5y3NEgpZnFn0RPVMvKRDKcg
6kkSXhmbInS/wlHTpIBhDuM/vP9kO2fYM/wYe4A4GqMwe+tC+gzn/xBFsKXvbr4C
TXbFhKhWkdEN9k6fQR4ZsoLTQwxLnKjDtBENV/1G4UaAgQiPH+wxiuj9DEe/AjEa
85yhuKiZFDeTnavqLLPOoYjDkELGRneH+u3U3rmc9eqoPNl+BubAm/GEo1kUWu9g
hn90afbhSTVMopaZt3Ra9bxzsWyOGBAXBYktIacoCw806amVomYCHuxwu8/4oqsX
j1bl0u1GT4ILBdjQ1DB8YNIAB3aQr1oSOYKfJxiJ081J62SKyRNpJl3HaRYKwXNi
Q5dmZxLoIZRIhXKp1AXelW06NucWQO/Cpnes3zcTIBCbG+FeVh6tBnkI9Lgv+6VY
HUGF46bXzzD78vC04rNnbqdL3HCm2Vheaaf0qgg/fKcEHx2IajokkZrDrk+VZxFq
gnMOxBWe4jpFtznQ/l14CBN05bdHN0kziekM8fQvpGyj+DxXEZpUJFnmW8VrmIzd
Gwj4KcwlGCqP5WBozNMcWd8fgzjghQBEXPS8+vemdmpt4e1zJdR4m92fZU58Z9wf
uARxvDd1LJp9OxaBXmxrrv/wOcrpsQ+LX4x0z9RLbh8uvIInzLnVLeFByBliP/qt
7L8oZj09L6PYfd+8juN9RLhSPdUzGUosG9sbntwGabLAdKu2kfxMDKLxBDZWQbWa
iCAFtAOIn1LLoHufuWfTx6Ieaxk8LxR28Eh3OqYjkVeI9DtB7ThYE+qKtQNGbn1c
i4gop6XHZUr8NFu5J2lmZUDIsWk2pli7YrXOVMY+wO71I6PXlvKe51VHnvAe7sPt
6MKuZi49R4YQrtHVY6kY7SBu5Tm0MbMr6iu8qhHkpGyoEgv2s5nRmtuiNrLDzfvw
7P+9X1Lo2PzCkKWZmhVXCdl0QFk+FiUGd9h/0DLQXeBfAqEszMkOEWKo0fH0ig/w
kT1NxY6L5XZAo74+bpRumzR6GBO2fhO7Nt4qg66hWjk/H5fmgkIbfZeZ76w8mGAv
3sJMxgbnjxoHF1GiaTvOdU4SyZWvwcjRsbjUCOhoeZPtbYi657FmPqbqa7Y7tYCf
ulbvASj7DfycRAxFZ///UNu5oqmjIHYtxW2Oya2wLXEXRYZACxjBl2doy9a/lYPm
bq+vsVaeei+dkf062rYHncmif8XwpfSq2oZqs4K4c9kExP2ytrnOiiE9l930t+4u
M/BSQGEqiXevrCc3PJ5/R7bRaTUt4/CtqL+OjvrA9V7MGFKpGTG/N8pHRrDIOypY
zwHYXXIRrBOoPJEk3GjNuvofkkeUdQUvwDsbk7Lnkw+JPkAE+10SHRLiLwudAHmf
zHjhowKF/omandUC6BSuyzedB5OS8MrR38Fzuuj8rsATJH9UoHAgzGyeVaJDapCn
Jh+7OPhCSlR1C8mE5PtoJxQcHtUcJH+Y9UyboOcNUPJBuPq/FZPNwERzRpx6siWh
4mlBn8N0el9adhbAGodbzpgl8hPoJEEYlzSYiTKpVYBijYSoxFVlrUtjp8e97I6S
DcRshfIWFD5AetmT0ZO3cldJvfAnJfGmTB5ftyAuBvmndGiR+KXTYjkuQ1a5UKvh
RvBdBOKEGQR8og0eOfPMLmvEcAimgC85bXYA9o8LcfvrUXc/76Vm50gy7/U1o5DC
xrcHQhC+XyusDAdf6z6F27vdR+lZmdnVB8v7rg87L8E0dQ1yZjBucql9CbiSrfDz
8n4wqb33VHb4e0vNeAWLd05uUrOPHRqVwFZ9dBIR7+oC8xurnSgQUQlbysWHAHPO
ecuTGKvbIgz85vs1vYAUweZZm5pg1UI8WBM8sJHFVWZfpXTyso0TI/Rp9RNHSzEF
ffbmjwIOZ7n89c16FryJfRIu4LsWwNpy8BF3g6bBr5+1V0Jb6CxDNFG/CqDic9v+
xlGI4ietGntanG+l9kyQ83fxTasCHFpP52ts+Wb/GROtNSVR7TUwS9GHGxt3Metj
ofXZQGClwGgaAQn3eGVwqAiXaL1qQnIym945hfsPvk8roqV/38Txl/a9ltKvFMbD
riP0TTE81y+2nudF68aJeQWlbyZ2TbPDa1Ct7Ipirlk8exEEk2BR5pnPpdZZ/CNA
6eTvXGXiZVlblh5Vsz3rMiCF6qJEpMsemuuNwVMkwUCEPi6m+Ko72pLzetIq/6Dk
WO0SHiyqvtdgGuZ4krRrZiA0r+DWbtZq33Shk+0I+XyyL69+lt3ZPO7vV6RJ/sTD
uJCwHFja8ljcg1u+i3xMn90fJIkWdJJE0P5y7lLiTuvjCw3vXCxn5f3AF7umr41A
4kfk/M44gK7Ye3+RuDYyLRA+ziwb4UDt2OmUF1ehUcQjAgzOr6f+W/dMZ9KwoEYC
8ApS3iadhcOdejnOb5HU1l6NnvfBntr6HfzFmarJV9qgkkRRXq9aMANfBOsXcMdj
+OZww7Jn2fFse8b/iUHsoojTe8/5CSlvTBYaOJYjC8Nm0fU7Silq8aKi48eP/SPw
`pragma protect end_protected
