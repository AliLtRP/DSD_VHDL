// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HkhtYwEdhqki94VDKjb7Xik6MLLW8RqnMc7vLIfVLj1Gv60g32Lu7qj71aKGKuCw
ApovGnOtbSX4BENufcaDbbAY2odzIZ9EMcVEnQm3s9BA++3zL59sQM7dWSPKHvN/
YERSwvt6iIgtcy45m22LoFdHuXH4WYLY4M7dmaGCot0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9136)
9dV5PLILJqE8e8ZXqCJfbYuOSYmANdYmiqajR/vTWrYYtQJdUiZYBFf9UmlSsYHf
+IivuumKqd21GJtEHAJuhVULTbghd91/310WnLJVsZakcDmAkEioABltsXUC4wEv
fHaWUxzOiTfFnbFzpTvap4lF5HvDHoMbhTVOBBoTC8lp8jl+NKG8zt9I6T2esr63
3ovqU9iP7F5/pBe2sNZW5AX9f5G8KMpohLsIXtZMx42Y5b17e5lEOb8CkRyI4K7Y
MK0x+yahyO7Z9As1jwLsF+0Nlao4S+hGR0y/RYYiaIMM6JWT0O0duw6B4xlSy6/I
lEuzJ9DXHHEROmBlZlZWQHC3o/cJWoES65ekBEsmixhm5u4UbQZNbGVZwa0vzk+B
Qq+3tUi3lURrrmnZwWMckHrph/WokB2BrAf9yDb2E8/ps4+1eN6qXxgSdDOYgzTZ
Nmc9uQ0BUUBlEiLPI4CHr6MIUXP0A7IJW7eAWvALb3bGVlPOwSE/9ac5mD1/Td0N
R/OpnIZ2bolbVtdUm8zJylvSjFgzsMdxANS5ZIUYd2wHUF7jsHx5lEKs0WYYtMF/
9z3Taj8wlcu9mzuFV0j8MDRgHzrwOD5B4KygMGugIIBqUrZa5Fju9+S8bXn2m01q
MgRMLaJh4L6uM0LtHmbHArWCfsiHIrTLDzvzVAVCELpqOMBDcWKO5zis+JQcbBX2
HIn27aZGiFMUmvyAuTnT2RUmyULhbA1r46zToLkl8lcYzjdmzLuFgeE2GPBtixV/
nbTxK6ufxV6Ux2EouHGWjzx7vKrVeUprNW5Q8HaNzj1Y2EPVJfACQxoE8F3xsQIq
+u5PBuCCpxpWWLX3iSdqJqP32i7M5IIF2MR5Ee71HKGfHc9vQTnRfYpUlQqM6jP8
eiuKPZSPnUn5w9iLU1MtW6U3ugovtaPRjKGmzPz1slSmClsj2w87R/5Ps5mSaeui
W9d/8oFtTuTqnqenIRwFf88eqLCwM3eLDqj0RlaihjwPVsT7f0SXu2CD5OUi9XTz
JXGDf9nhTTZo61mbfdi4EtPNCqXmxHcmaVQmrC5SlDCXQMeDaBd21abE3ugT73D3
qy0qFdGTWRJCsTNYcrxgCQbUSP9HXq4ExNgLjz+A7X183QLOhWXDuOo0Pdl1whxq
mYtUhArGw7m56dqsbFVDQTnkhe4jfDNPck7SqLboLhkyj2i8cEx68O8kdHjdCdsw
lbjyp46sCQW10JGleX6j4vk8dtnYVMaSDubvgvEU9dMAdiH6/skjsSVasZqogpUu
Bk2nt7Zlq7suUX5O+Fr5LjjQAnpmDxEi01FMATjZ49INdCg2bRMB5TnnVl56kl9Y
tByWFk5IfvN+QWZTbbHPCI6kfqcj9ii+xSwl5InNHZdjUXsQVBTxoaFCIYGYsB7z
fUraWizlNfQBqVyGNJ4f4mZn9lyUzhBIuIviwG8TyPsFMI4lgVaixJmSoi6C7xog
+oFEu6YBjbJ8Y3oN+DfsqRGZ/YS5tg3MvFE+iu0heV0LNRt3adUWyJgD+ljrI/Qg
aX3J9yyR5Ss8/zvpom2vV38llaxTUTGdl/MNtAGzJIm3RGgd4YELXrxDudP3HJ7K
DNAp43mRDmtpTWvulYEXckwsGMO7TivUO38/beW8FsiLVYkJB8LmzcPbZVrADcWo
b0gzwoi5+oO/L+c3qFBzGbB21zGK+uNhyp6MOwoGlE4AfnoCaoMv15kT7fteLk9a
X+fVFo7c4onDxRZZL00y+BeJFJHthc/4qzN2ZTakmKxlMUqdjqOM5OfNhj+Ej4Qc
ypEAUgSNdJY758Tv4vMXu+Pk4tcqt3Rv6WWKJTfYQbRz/J7r8a3m2S1yY9DwKT2Z
qLi200gzcJY7ZAxoUKssyw0tCtYbZiw6js4V805LZINCx6ucO9a9mFaZsSNMK3cp
yxiGIWIKCpg5G5xbTT54FXT980QflqOLt4jMnnx4yX9nV6N/6SktX1xi7a0frofc
l5sCMnXVaqOiCAW0CzK5xBN9j84tVKcy6lHVKEiQZV3pBoHmGAl1ml7X7h8YC4zo
uBwjjRvwwncv2QRVyEfC9txO+d2x9GpWVefj9b84YY6QYRud80t0Qo+LFfKzaNGK
SQ+0LbQs8sANUp+YL/Jb3m3fxTWKy9amCkHkpDdW/v4dZ1pxKehYn+5FnmFhiNyX
MQyrS7xptsGpIUvwt0d65LC7DMaiE8MnhTuoXsLpQzsFMDr7YEQcDlLK8cfwTO0x
8nKpCqNoxktw3XdAsc3qMsn++NmSRTk2xZLOKyQm2+qe+U3LB0l/DL1u3MeCSPsL
TIUPnimyhbkfdSn8Axmy7KRoA/oZSkiuwv1iYTlCwZ8V5HGdAxR6fpsKX+SsJrsS
VhxHoorPHPcBlinnlvsBzLecHmHH1lUt0c5LyL5q79iTVs0LPFmN19CjHC+YaTxy
fQU1X1rN5+qLyvp6qSoB10fUGgMDgu1E57zsDP3+Ji7vC5E+jnZitDtM/cmuCDeX
M6lJaM6RjOhxc4Ix1hP5ooPtohy0cUBLNnNl8gywEqAkpzQIgDui12xQtJxe2Xg/
Apjg+WIkYYTg8bJl4YGfLLRe2bjP/Bufqcbl0r2AMJCO5VBHaFSrDZoJC6Qt+9J6
vHTN5bUtct/28c89YovckWqY5oskw8u+H06LRZ4QNqYyPPSPVCqc/yXBe9QInHT+
o4wh69kYMUic6qXD4gccLLyhelsFbcFHZuQ9nxXmgRuuNz2rgp/FjDdbExApYZpm
oKBge5Lxl50xExm3vo++GG77EB/vp8HnR+NWkQh4JjlrR/bGsklhz66weNEjxGHb
oEjpR3M4/hBE0ePIP21T8GLxdB8fjX2RvbbgIFFeDPEfDMvyGMfjJ6al2VCzOy1o
P9IGeX3tdoUJS2SHCkC9NYjSPpAha9XZaMPhel5WZ9C4IxVRNPPFFshqIc7aqhBp
Nyr5wIb0uvsx4eJ7C4WnWieP5K2zrHvCHL5kt55CYvfVHERiosqMDAIXFnwr1WGU
5QkEYsr1U/6jTRKX3SFgLyfDHqs4fxAWp/MRw33rc7dhuXJwojuX1+l4PMXTWbED
cuFNR95chGEUrez5xvRlzRPtXXznHMswM0e12NFEM4UhHLSbIoA3dFy6bEFUw2Gi
Wu6SfTHysvWzF9uf0eIxuX7qGMbVE6iNOY3FtGGlWc5kiHm2Y2N+r8JJWmNvWx7e
DPf7UA7/xrko2ln8MsKHsvDRIAbeNp2n+pIjUQI64G1LxReN0ApoqF+/PrRqtrCv
0MIv0ifp1S3LTuEx4XnEnVfp++eSVd7TLkG+Mk39CLLODz79S6mMNas3lvVYA98y
BINCbVr+2x7xcS84ABy1O05ljh7bY4AqtmSNRvp0satARBqHwR+TbPes0vj00RT2
JmvvrhyAmIQmz4tbE+G8mUm/LvV0GZb9WqJ3SAtq/B8YrjffWiTbsGakBxCSAy0Z
EELSR+v8xQYpnh1pr8bDap9XDyHdNhH82qpacsW6vhRsEMlfXto4xNm7bZ9SbCXn
0Rb5YT0xs/NWQGnpUrdmTswB7SyM51lWzIM9nRNRFye/7l7YoRqnQXMN28vuV4Gp
BnDRhu4MI6czQa4BG72++Gj18hOXD2KyjyJzG0y5mNpirLQiiExigh/3cbtkCJG8
hzvzMTVIg7LGW0uJw4hplCZeZomKXOQXwDfAXNL93/rP+kuLJdvLJyMitwmnBe3w
A5ZrisbBaEf/oJMdHEuG5NATU7JEULI130hng/fdQmMb6S6J08Td/uS+rSxugkLt
mmRLxdARUv2BL9nbiVI+GPWur+xYHTJ8l9C2yVBU/iQU5WGW04I9FxS517mTvMCG
3rRrNlIOPjIVFbiaAWGP0r0LGTPVlD2fNNy3BDz8HhL4Xyivp8t4oza6H61B34e5
Clex8I7HJ/TNuhdYEMHomwDu32HR85tReL1xFDSXUjCarcvhZryih1wEEZimqTud
Q4Oejq9862+KBD20/1vUahvVbDNXdeFK2+2TeDOgTo7W3VRXJuEg6nO6ZdiOBoZa
GxcloijFC0oCPkujU1u7YpvcQo1TwyeecTAOtmfF+BiCOd6OC1hBrRUYUkE18j5c
m6m8f/ojUKgKs7RufQSPR7Ln2+ZXzxs+fb0+OSqPolB4ihzB/QYI7jRhBonL20zA
hbE94wjjMvNtfC6wLEtin9Wb2hsAphO/JnOOAs0yKMaopZ9WvL621CNJ5g8Y1FKC
AqCEnfKac4ocPCtk6wUEB4/8IifX/H43lCZ0Wuw5LCTFZzbARQjHEyt5HKNuKuu5
na9Z3kQ4fc1kn5uwgrtQMkik2ZzdHJ7YMs4SLoAt8ECugIHCHM9bJ9HLvPTpBoQq
Y4kw3+Y1JuFv+FvZyjf5FRcPEL88Hzn3b+VetSRSGfUeO13okBDhwU6zB2QvS/k4
8e7M9psx4wcqpS4QdjWvA/kl618kDTBoc6tIYZvW8Ysx1+58if9DGE3N9aoDM1/6
P0MAAzDCoDl5zFEYGi+IPi+jR81M3DbJ08U6rIrH+Z1jeUbaRyrbiPkoavz5dfQZ
0TPeB8SiB5uSAuBZfgkZ6vxaFkXLNeCpmfuPMNGEmy0DQmdsAIe93ch9WqAhJigT
RMA0mAxnUzSUZFxfoX/+UB/DOA5gC3mPF9FZP28biuJVquooCitn8QBVtv8oq110
3FcY16weXq2CcHI+Df4I+3bhZqrWh2T3jFqJ14nDEE1Ba4or9SBwSLhDs7C2QJ+4
pkCHxqi8t8GJ3YIdqlokyv1T+MO1o1UmPjj3LcfgrwAxhlI0oERgIfJV5kKIuh6j
JqwdtjEXyejTLbS6jRg69WGijqquTz+dMnJYn/I2AgMZY4XkDYQwUArSQmqzaWPN
pWyC9t0DeaKZdIELCb4etrkml2IX+D1bQbmLlP64XLiZx7uMxFz9VzgWsN1kUfA/
iEvjLRye1M+Q8ff7zvVxwX4ZQoODWaiOidfPHy/p63Rj44yhv4zob+PHbrmThtiN
bJ4mMD7lDeMyucLROKZ4FQ4bVpmT8Uwpw726JOO1ILAhbT5yAR6kerdBVgkQmKNA
RRcAAJWdZiRltby0qigztSqy5FxAUcC6zLqyFhqfntI6l736mujWVa+HGvBexhVC
exGkllRdWUl6ztLUXaURaVMdQRbizQ+9sVOX9gCK4+FjVR6gzYeHhCZzumygADk3
/2L3vdtl8iEnPkI2hxaHihclH6wQa3n4o15M4x8939Db6c6LQh6FHCwA4tTe4zgZ
cqriXMJ/oSL0o0oVoXVHfAWp1popxTq2z1pmkAhPdQ0r6z9EzgbNuRMqhAW+Pnll
4fKVljY1+66GmtcB2a0+PzDTIMvmYG/TkqXx6Tx18poF2I9xV1/pe/Kl8hL54Lx6
aUQhpweWeP8nIxztPJQeRTDHSkmJBcg1SUe3X24OgfhKywBxKLWeW9ZzS8TC/c+Y
277qBeQvfg9IGYHGmXha61y8VVOhLzlPXOUmNmG1LSBacpwA2nZVmQbESgYMvVV8
g6jaJLPa81MXD5WsYUq97w7s8oKUb1VTdlDLHFYMuFeTEUy6063q9m+i4cgq5C6t
K0K7droQTmN2bUIbkHAgUDRB+3VVbjG85vKnXayNKxE3XzkBqQmQg/hsfBUv7ew/
zFLis6Myxp2aFzwPA7lLuk/dj5vvBnWkRcyeHaoDgoIXQ9x3T79WSiN6pH/nFOre
akcSxy2+Z2J0ymiOipwdHCh07cD7Pvns7v1d9dajRc1ZH5fkrBItk6GRIc8gU4Tz
Bbo2hOaYIazbU9i4mTY7SwSbDrCgEr8lkIDMDrsiMs5NDSCMo/IeSJ0EuXf+2mmd
iJynBplVQIoN7CxW8Y63dxAGhExpgpFI3kIhh4vJM7Xem3ewJX2uvFPer+rCfu3j
cIFnQykcjAsU5fUjuSiHdAhPV0RmL2j7LITDNsW9mGJQ6c6kN2tDRX+c0PUyd4Zd
pvdBclHd/ynPifOjijHibmNFdZKZvgNN1jzjth9tZItCuDJTWHa3d/81ogOXgzPj
EOW6ww++oCYlUTqCo48YjEGUtbuvbZQYOHJAIfdcAjNGbMkIxNWkQ7DuTtx8x+th
Ly9xqMbRXo9woseayix7IK9BiXu+Sw3mcaQIcy0IeSuUd7jDNXz12b6RWPQR5L7W
mpd0MkjK4Rtxe4BjVgyWDzwbeSdyhCWq72H87a1hn/307zJHtl8w0DuecIlPX8dS
YylPMmNEj8LhYsJ8e0J/G7ChjV5e7bCMuHT/2TXeNdnWNwFIOf/QYIGJNfzsj/qT
+Qmlw2OLukABk/7pohU3ufEyXlbzeLNAaAyB8RJHouK9KuuFU4wG5UCcGcn7YFhW
qN2f/Db+pBVKYcI3TZQXgRLW5cZ1RcBo6TxkakyKyD0HMeoR5IkkeI1fDoNmsZrn
Nr804tbxb08IEH90831Y0mEtC9onO4NRvVqBblzp4AU7C+f2PsapzkTI9GNU46e/
6mhkg+O4rdEC2TmGaglDlJyFmYxiCvZJ1EgXjlX5ZnFT7+gy9pUpZTRUmCskVeUj
Hp5TflBNvZ7AIiG++1uupiEiTK1d6u5fFhQdmLts4PwmYz/yZ8S+u10FNcfM+C/y
f9oRLuu4RSHJVgN8WfETpSerTnsd5uNgBqYkkAlFq9YxNgg8glCpC38J3+yceLHf
GNfsPFr3fXNDoQ06UHtYWPvFeyv5khK281j5QpXXRM9QN/7S7LbSLz9DAx1HK28H
oMrNrQ3QDP82V9mxyZmb+AMr4l4MN1zBh27X1Sg1VYfBmPN99GF5tMAc9iHNgBRA
LeIr1FTuEqr2QGaSRyIBpVY5t57T/Cv4l/Q2e8PUPA4ykfTzMHIp8QzJhNeGXtsX
W8osPqPLu/G7HySfCXRPAHdkYIqhNMPm/0SIvN7zWw8A6kbDZkMGBxMxBJNnYFgq
J/gK5NbA6ZZm414OqEuM2NA4tmqpO+8tkuwHFU1DVTXw8Nsnd7rITDhSwGwHIw/m
IGVacJec699X1IEB3Ox5KTLTaLE2oN9CJdfLLBIIEfvFRCfNChWezMvFx7NBfT8R
zeIUHWhu9UwPgTltFCu+NDJ/UXFVyajqyUndIoRZRpjbBT7C3J9YPyxr132bt93J
8KHhTjczZM88X4/fPwjYDQwOsB0Q/z+MRBjFUX3AqqTSMBS2b9yH4ppOjlucT+MB
WSepfAqlyx/APi04G8GUkr1IQjYv3SxEFbunPe2oyxgqRHq794ue5t6CGs5vPqS3
I2YCWQxz0H+zOnTK42MQ2GkYyAbjHoyFk865Zhi8CqthEos8I45Q2a3WgxiumKjm
V8y80MOwNAw8s722q00tdvBkWeyFjPRQmdJQWHZE7GyWGq8hMOqWsfqBGA/GhqJf
70/HshLMDDftTesDowlS8XKhDBeyuR7TF31wfLLsMk/fJgZAqWyOtVww9I9nLzrn
zEkRZOEYYLpXRikrkDES5ZXFEKk7LJJgDyHujk+nmMQOLFxeWcdGMjDxQAjbGU1g
rBVGvZNovlQX+R4Yq/u3avf307F5bpm6+wHUr6vQAJJxUSPBKqQJ7EhPTQmincuj
ePr60Z6JHC/NW6l46AO5HLpfm8+63tNydU4C1IrKeDn4Ye6cBNuxc1zoouQlMKiS
WLv+JgWcaGBB1cvJtBeLbUS8Cg/o2sYZRHxniOvcNz/nYVky0CflnuOnV2JMjhHR
lbpgjxtAG8Suf3ZfmReDgIDtGu4NAgPgjpo97rOS91JTAx26HhUPQ/s2vBO1WDos
B8/ji9XqBl8TqDSURGToXgMmbWLBymKiOu5VgsaE0FGyUAR0PuJ8EtkkFZOUtsy5
DUa0i8uJxv6fDMQilT+7KvHGYwY2JnLLXo86y3uSREfgj5Glj3EkzdwFATlFsR0Q
uWLxdB1g09KjW3gLMLeBocVc8T4IywTFtgu/fLOP9FnXJl3y0tzSgyBWAOJaOoyr
pAX4fZmNF1kSk6jyE+hqBPtgvtNo91FehWayZPc9KGbf3KLKC7LzzmUbesEH6S0V
LdyBQm1owmQjfHT/zolcVHRZKgiuhx4AdJ9UDzX4VUqXMb9gIAe1KE5OPch+NTqJ
/+Wm6PKsZH2F1CjMSBblUuPQCmWFKcVgOUbA+RgOqJT14ZqHTxbnytHxrHVqYh5u
RtNBt5lEOFss2ZkKueQHvrLyrTVmkyJBHt8zDWBeQ0JFFBRaHH1iN6/FecZOb4dl
m7qyyKZwVZK6TV6/+gilELjr3TOJHkP1Xz7Rfkn9zomZSEz9UHolR8JBQ57Zr0we
PVnfZPTo7iEklz8z+pBdRs6V5B7m0KuOx/VrjnowXbbb8wyFwS9y0xgZBxTzIceC
Br8CNlHX75+fL9Ngj6v8iGBs2eDniFWNd7+83GUXUh00FKKOI90/oHReWYx8z/aH
Y2uNxlH2GWCet3UP4+OVDnDUF1PWCjsPGTjF0txmFlHsvDGo50GM38sVQCXcFtZK
EskgLUeVvJGVQwUJqV02bWdQZPq9r5J6azOho71Oyit2ox6avPxifcVPZDMoKeLE
MQkyWkh3mlDvifTtW22ihrlPhn8ENORCvRdpe1aKzix++QmrhZEH/tVF8lqQ+89w
p8Gv/o8n1vi7ZcC6tpmIEfDmAjl7RsYeHckGFRGltq6g/QVhG0ehE5yPbsywmZV8
ErsPOG5VnlMOudQ8amPg5M6QMUlbfJ0vmm6rGLmDgJJCMxkpko5hV14Iy75jmNZA
AGfxsPX0s1TAAvXNemLHnFcCyANF0/ihzFc6L6r/HAmoOyqcAOhQ/J7BZ/LIH52x
ixjCLba1omejKUVVq+oIswFDW87xnhxEblhUxIhDjTPVgGYhg1Ru5D2gQJ+IPCss
QbXUir3oTdzMTezTZ5DaXAJV59mIGIteFYtvth6vByav2Ul2ysvDDDzsQDlyq7IG
i7zdsaxFTUI7c86s+rTnZeDHFk7rBljrle4zOEhwJUlPam8Luxd38p4Yj5cEs0mM
wvxKwnou/9WorGSogrx8EXSLWkE75Ce4YyiKoupmd9HCLMEL0OiUuOIXi1l6fdAX
lgxe8uon02v/8jcr0fkugrAg5ARyCBwoYf/Mg0nSGRRu7ecBx1RsnYaA5M/AiDaT
7bxoWwlqtlYnkS3sk8qN8rH8uEBdU0hqWhPd0LYomMfBi1Mc1dbRYhgk8BNJlN0J
mK4uq7GdLI4R7ACh3cdnMhHRTvoctsQGuCKTPA2TvqlwYKmcpuYhyswunRhQDuBT
EuIaAXSpuhc5kIr95ooPmyFK1VPhjIEOLkE+5AZtT1wuvYGAepbOQ7hw1jwRGzq1
ENArAybjlJZ0DzkBM8BdhCwePjew17ripk81EOboLbdoyEI3tH20QoB1orWDtChR
afC4kF0byosQaz7/uJv2lx0JEiDQTyiQ78nE4xk3VTtsNWTMTjaIKamkSt0/+nxJ
MNpUsOcahVWtCymkWFw5BqO8Ohy9UgWh2zLtGz0qd42PdqOHXnKQyzfFg/dbt5Y0
PS96rvKfgOkex9R72huFjh+cvp6+JvKOU0BXBUg3ElREuQ9R+xDVe0QSiLptvnTX
8izXsqFDk6FZvQEfcr6f+neaCMMDE7rkjKNSqblyYtWajiwQCawDmquwDozO6q1Q
Nq9+SmYwrxqnGdqqVnTfsqZZNGKBLt7UamnSBRiTPuUV/GNLPufF42ow1doE5H0r
oP3HHPGrWUcGDNStJmVrma03aM5me04h1EBjb+uc2lZ4rcwO3xVSBYJpDMA3s04a
3CF2SOijxESwBk+MwYVxuIZ5pbcRYLgezajHMT1bAB783icRNObqtJc52PhJvrJp
08wRj8pVHzdZPcBxeWkzvfJdKFKeyGsm7rpJTVj3gQpTEngqxeoEu45zP3OuUrL5
u857OJjACRRvfI9FR7yN72dM/0O3KPbUq8nUSTN72Gjpb4XGGCxi+nje3ZvCWiQE
94c4g302RMXMUfYvKFAjDjdO4g7XxT91MpmtMKJGEowhQhGpdB6WUHnvBinbE8sR
fIMLxF8RFs2SOTOwf+VvuPYYpbXMdy3uNjuBTc/vLq8rzavgLSS4qoE4fy5abjzK
A7R/3So+DZEo+6S/uPUDV3Pj+SrQbZ7FRpY0/6LAoI02S/a0D6A67HVT/Giw8kt1
Feaq3t2gbh4T7bMKrab0ANPJGXCPyCRhnZEoCeb7kdEg2Y4vcbHVYx+ra5Z8Gw+A
/ZOhLgap39JL7OtadjR4E52hyKPhGY2cYKCGgny4yhfDtzxfH4+BlgnX8yxYAhJf
ywHgoBoU/fqEjiWSUxeYoOaxiirUvZ7nSsKj69R3frgo+nJBpNEl3/QGgWnTmUJT
+H0QYxOtHQzy1V0KpKrVhVHMAOruOcFeIeFBkdRpdRfSoUjAqCMhu8rs22lp2R4Q
giPLURX3v4lepXd+CowHMZAaXg9DP1PU91k+tnyowBOt6tOvkkpmifooQT4NwLyZ
8sKG5wiMUd8mUYwPvprKAerOoAuBPkghiG+76MeuAKPbj2s32FqJpuJRG4vkPi4A
vzlTt7dQBqQJdqsRkZ0DNHkajD4A1wZvckPvsImk1hBAZRyPt+3aAHHkLRbXCicc
Se2oGmdy9uMEZ+n3UU/cSHz0KKjrFt1Vt1JxWfDpQk4vvje4CbqMEzvFGmu5RFMs
qGn3Kmy6GdF1UKlR7SCjccJGYU9RQrHTGjjCssh4S41vlhD6yxNNCCAzzThO+xDM
DsGpAbvzY4aTbnypufqfQD1Tvy+y9C+2kGJSux18vVX+0lgMUg0iqHq0iTYwqdTd
Qmm2wCeb38aUMCIl1MWMXUMKohp2/QiWN+USrAUYN8gLG9hPCnQcHpq8WcfwuuAZ
Gn6dgdAlWXN1+1j2xEpIRhjmgrlNKbUo7rIbK94jXhrs9eRFkV9tfIAbLHX/vbwg
zcf8TICjeHhHGUHyDLvi2ubJlXXHnfZxAFUTx1ZSMNS8o6yTAccQ/Pr4Ex0GZV/y
InAbOopMSa0aDFY0TtkYpHEIb2raifN6tLxVWBfkXuDB4bBGMwfEdcAZ40QUirpR
r1IWZkXOK02gI5x+LU86j0ln+4tAEHpc8MkxFxeK57rgnZHf0WpurX+hVvP0Tj1E
sBKYRS8x8fH61YipV+K84pNuuuukIWCAxiiuNLG68uhP5HU1kC9sfVnfoiVTkPhM
4gfir9fnO3y+YnF+5fDQsOQsrTYS3GYY3fR9mkF//0VbqsUh7B5wtbt+DDwVur/T
P5ZaodR5dtskr5jJj+b71Kweu3aQ/h75ISkDZoOp/6PMW7rG8SJFb6jEgY9Bmhk8
3HQbYNf11HnKCZA5y3jqHX5dJhf0QPFbb31Ep/Bb1RJcpKxysbagFga5f4lcF0mY
wJtJ/0b4WnQuFjd1PjZTbpIeROuoSm7G0wo4XUkqxGFXz7HAiEG+KTT8dLzIfspk
o7pwz8qRZVmfwPPOz6bXPfcAaV/eVaRo8lB82lm0RWISmL2CfZKUGgYmXvjeBgys
2V/szVKe5HvNm2YdwlPS0CIHFmksL6LWMBMQGfpy2hWx7/ajpJigM7zkKlxRSZLS
hxsxOhlcbiS6r5j+uS5yvyj91Wxthgr0kcbGadEHwPC05mGIqkVHl/thYgqPwxeU
74mdm22bPBamu+1SwlP/hOlXxTDFyPFc5FyH8gI6xnTJfVOGS55gtwJt2udHOYDQ
uMDtnrVu3dieWLgW3O+/0SEH1rl7WQIvYDFBonhG4os7NODgMNwRFe4T2NvWXEDN
L2OXn51AQLgZq+0OsTGxIPvZfVdr7WhAXTA8jV+Rz1TAwh8lp6qMxcPPTswD9wpD
v3NItsDvBodEYXNRNHehzdPh/zjP4TMXaBwPeJXJkncpQSPq/5VBhuThdxxuKG0M
wAlPdUa/BT3IOhbvxupYdXqz/HLxwXqV2+VB3gw0zJfP375MVeg+uvsFLmy8+RBD
HfLGbSHrXBOKdv6shyzYeX24KcA9nonVY+uIHFXoYlBemRys/kWWwrVI1Phjitix
koTVPoFi19JEnmfOHwjFqB7wG1G1kBv+7wh2AGoDhxxmCdSlEjzpLVEzriKCgXTv
Y7un60myji63dvlZeWkM82m5rM1+ulkQ57DzlhWxP/is18mbPaOLVkgeY2692OKa
p7y1gjwYaGWhHH5j9ACkt9IfFLNE0o0AEReXOh+5BPhIcAuUZYPYr01QKv4jO0fE
epG9HWrqC0s0N6S76wNleQ==
`pragma protect end_protected
