// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
rrrxvahtPbcwST9zztRt9NmJjnybY9ryPQdiconA4neCQ9JFXXn5r9ftt3eUIhUMa5EYgg4e88iy
3Tc+rseIyKUy1zuZVuw+csCXyhfQAtvn1YuNLIbUrkFUNnOPd2o8JfHngNmHLBi1JNFgP8QsjinQ
Lg6nnAx0jmoLL1ZO2Xf1MA8sKVodxLr4tioDM2wUR5G+cc3iCWIMMaIUQ9YHkxRlk02p9ExsT2p3
kKFDSy+rlEydOfGxMM3EuC0tgqWeDk3mXwin4+LkwXk3hR2Kxp33uXV7bFzateMwjyIA7yro0yAN
FNMyc7N+nuhQ91/SLwHMaZw90gR6ONATZatofQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
A74RHgXkkahqUKSAZLLRsZwvDSmTJv1Pqa2+lB3ElxEO2y4dNgFSgyaiIqRiuxHzv9UEGbN9y1KW
aDuJNj33txHp4PpXMag7ajUa72t1GH73yM0NUakHSdYy4MH8Zu2g42Uk10L+I1pIYCV0KPLzx6ae
l9Nz9IbdMn+AVHFLqmbpFjhX8apwRc6Jslb19tICMmMrXsRWAms6WVPvgzPS+wepVLUFhOEmIefv
/pnIGRSSIB1XYnPenYpmsbkOlZcAO0grUyRWGN0Mrj3/o7sN9ThWyKjoSY0djTAukvH/W0NRp090
bFu7TTVdUMYpFlAKz4r3ngc7dgVsfc+KNrSUvzVfYBAXZ1w7Br1VBz7Xe3lNmSgvWHDVsvHyuuC6
yuSbVKxIrRKSs1tbAR8fOXKmlB60xnZwF9SlXeQRfq0oZhUZGrB4a14IeyB2utZysLgqNdvbtIl5
WDaROWSHow1qpBK8tlV/diunPrslcbvghy+VBzZirE0zwj4r8dt3FL6DoC7SZ8SOoaioJwMU3oVk
Ul+ml6GH2J7pnwll1XLKUQrkR6qfAtvMeTAg+RtClk+P0Of4Vwl3W+WLcUyR25XwcSOg1bOpoo0O
qjldafZzziROOBamcAqwrVWyssagN+tJshEPfKd0Q9bqBbTAcmXZJaR3MRLFxc2MNy6uxRhpnZRr
NL9VzqH70gMlNXjSkwnlS7W/vt8H71vkJBYAhONQFOoQG3oXU+3FK8zJxJ6VO4nF10p9HRt72Oe5
cvD1c+qN1ze2HBlWtzqyefsmjS+3kqCZM4mXvYb37cg6Nz8fVxPlUqLh/PiQxqYpjjxBo3YrjnNQ
Qp5UKYFRMdFdyi2CixUL3d/PiAbObnIgo+jQJOGyZPyclmTOxuAKh7fjkw31nlQ1wOSUdHedG5A8
ssaA/3Co5ki7JIgAb6jN6a8yfk+omfnQwna0/4nBunQl+vQDqmHvW4xWZeFcFHN9JHr1tzOl1UB5
UWSbTVaxai4hZLpfEAshny7VRPiIhYnchGOL1GgRAPohrOrJ62dfgJCApkQmZulYb0rKCbtp4cfB
BMS0T/8z8OyJWHbBfZSZnVnmVSvs9iShWxcoJDaIcYJ9LzYUtSh5cv1DSWnEA06u1QQkxhmWvdms
nw1L+MNM21DoHwZSK8AHGkv2SJKc5IJxLDownMRhDfy3b3sQqCSTc8jge+rTC9ahoMi5+qv0E9qY
EzWAUlrYi2/KR1F1fgHiWQjKIYWKs4ikzbcurnIxEAq5UgiyE45dk05gWFu19CzQ2WC72BK8VGw7
RxYOkiPhtk1MgBqjyChsqhQAluF51n8/TnXUiq1Y90fZiPWg4PHjE81fEPgGWl7y2Rcz5aRqo/Hk
TH9z9LU/vB+3Wz58ZqHQbC4DCzTS4e4UbGMFfi4WhGiRzn56yn2IWwT6u7h+2cxvQT+PC1Ofykby
VVwNnmx4v1DB5tP731TT709S44ciOh5XI8MOdzEyeSjV+6Yngql16XMxsBDOrNfngGMqvCo1YirK
IFM9lHZst6m9SfSYgTZTUUIqGJG7z7vp41FOqgCxySQ2HiyF9jHLtQ9JYfprvjzFR7R3crwVwevM
TpQitNAuxWjsQjK0msQr7UB8bS1r3aM4n7NcCYFkKWhrQ7mo1g+GldwfehU8IkOOBofxHiT7q/S3
tarcYaB6H6PDGp8pg4laBE/XDOZPfkr0k4frWNTcwB1lg5jdxfpjBrAsfWPEcdUfK1pR4JMp2Sf2
A5JbNfhYcUFcba9lS+oTHagiTX6r1P3zG+g4cjoc2DPwFi59RzDxR2J9dE0gwSrjOtrEznw5NAKg
QLc1SuxEdmVuAOcBNnCJPoir0BYsFKZgo86YJnOSd6H9gA1UE93+3kOBcUI9RD3jPwdAleq+8/Aj
PewiablUbMzAzR/KWgoowr3hTZ4XxSTuTC4bHAEFDbuAv8HTrPh+eQQAHCxJq4Xx9RpPbyKIYtNE
lRiHX9/RkQIdpTxImFKV7V+5HWVu6HjWx+b+TFDCCnMeVqNU+AtQQiWUXuWlJVsHNn41JWyvqdY8
TZSV6vvXi2/HbmIHw0eWTF0pinf1+Jk+OedO7kX+JPg95FfhM6wRVsldQ/7fX7f3vnxokvt4Yr0I
lW6Jl+q83mDtDUvBG8BJBL7+VfJGyyJ/ZyMVjh5OBSxL3beicbJ4OB5/ZBew9ivo9SgAv+UxPdPi
/uegokl/f+WBYGoQyUU2vTMnO4IRmu2rREwZTFFokxvfJS2VckJz9zKIusw63f1/jP3P1pqjTHKa
RqhX1Vx1pL3fjE9KQM31yqEKDaszAC7K3LjjSDyjzZtWQzkIh97UaFnQuci/F2OrbXI1o4KtdUDP
MxGfyZh3Phu9todyzsKmIcHrCHAtg0k6zNIA+JJHzIJXAI4WSIHOieNbYq8XFZsBOyX8CcyEtXde
PP+p0vX4RAMn1XCA/6/oOEt9GwTG6lyENPYK8+aqKnZU2aNuqgU2G38n32KwTgFLWRpbUP0PpNNo
o1soL38kNI3JFTKwzR/0h0I2+fnmGbUkchn/QH/0s0+hHYkEg1h3azuivJzmwVvW0vvBZaB/1j6O
hNy9ySvvgPbuE9A01/lJhPqRE5BPOZ2qdaQ6SRjjV+e++V+43gxwcqMvPVobfyKJBW1O+uJA5VzK
4954WuyT49g/lB6RE8lwSYjbx8HRIb/Ddm0meDJ4wYTeY5Zb/HaSSkbuWpkZAOeptR4KBvzLhTqA
subNwu4Ks9YKuNbdIor9xGMqjWTFGIXoanP+1E9+M4646LP3h5Oc5ZJ/QsAKL106oNppVUEI5BL2
h4dSXtSy1f93BESfYU5wYWxJ7NOvQt+wIfO4F2mKQ3fiwt8/ah5cspsVI7G8K6VcBnSJsgd6afTn
5hu88mPkFqUnfvDtumohAbc/TyqOc3Rtzlg1PjmxdfUzD1ftAsNXvsmRmom0uoLJFaj1i+5t2D+v
4SJAQLB14NzJEGinXe9zr0nBIXiAaMqo905nFOj7OLd0eqLcsZgdu5WM95oUR1yfN6wvOZojW2U/
iwnL14d4JgjHvag8fxwqbrVPFG8xs0yfKwt2MpvXcB1d0I+F6FP3DILr4ZquccA4xRHwQ4q5NNoJ
seK9OesvW2ShKnOj11LTK3Kj7BEqZq8r8DatB312PmCzOlG29S0VRroLCWHozyzY8DV3/NG8rCt/
CPMUjY8uIyrsbbeMXS2gNlc2yghhTqkEUekpUHQ4Fq0UP4vH3S7jWt6ipeXalBDBUMU4VX07Gs7t
A1qgbcjtzCRiCMuLjfL+auzS0OscyS7D9La1LdsD69pYWgcPbhVUBLW35jGFC5FGmEfUUBly/b/x
pv4gJZ2dCyL/D6tp2YoqgTWkAGD19EdMuSp6mIn34bx5c3OXONW+42FTCgxm0/9x8E+csbGqsnrv
amznMPzksWmW8nWdByxm0WBltEbbY69U1iJfRsbLWbk+EDbU3ifyPn53XtlqgMDKekuo2YJcbG61
fHVahF29ArDnc7N4Jk8V9wTp60UKF2bs7H6VBAfbz9bMEaEsCIKqZL9rsvt2Qq7m1ZDetoVmi8EL
RMRo9KmDyZ+4U4aNMWtVOv8h8OMAYiNUdt/qwuWtJH0Rlb1a7877gJ+A/ByJxp+Df9Tn4UZfCQaN
amox5/6Xz/vBa538yYrCUbdEQ8MLBWKJuaYUtb7H6wDzv4cWYAYmLrRw39DMBZb3gihtj+qmh+K0
KfO43n6BGr3dQIGvaQkIGBLdcXnbv/EzfNI1HH4Y9RVWUn1oMOxYU/bbgu8P5hPlSDHkhhKueEEZ
q87pHn5Qs1aZsu/qPvOpZYr+2NB2D+OId4V3y5uoIxxow0iCG6qigUGoRwjL36TF5IqZVIIevnDN
bHRFJlMDVcVk66aqWPTQ3O9pFjS7onFDONA/54oA2VUrLrwutNxVG5byYJrEhRMJCnicNsqMtfhA
Q3NNAWBST4rTYgRGQ7Y+9tnfNsxy3HsDejtJzmkOOYg2/0TZtggVZ1LW2O9cbMs8yGWddBNMyVW2
psbbbltx/m63MuFIpSuFt7wnPiBaOBmcdPzW6ArhqHIty3nDam583Pk+oMGb+uifjeaa9/sI0nRm
7Tcgwr8p4g+uEtPNPY1OMqbg36VomIIaPx69wy6MsF98eGIH4FF5crIUlvGYwAzSW2/hqc2gydt0
W+GutofaCE/Eih7kvidfnA7fCB0P8XsEcsHyLKughXI9qBfXX66sBsMkyRLCmGK0mjD/6Yn2OWgj
Qt5DcbiOpZsNr8hgasGyQKAai7uvrWYc5KnvgE3PKx2aL92Q97oaS3/2Q1WF1XQj+82t708HJPYq
VIlDNHAUD8wjWtu0nytUxLlvGlJ3LHyAkGTrOU75PGOQZ3EIRdi9kSNiTTUZZUaaBrsP7a5ppNWV
D3MqAnjsVk1fHuz19UzNZuRXKtWS4Ie8+ZZ7B10qA64yUG4bGp6JLJP9/iEd7OLkYChef8I8A1E3
+fy5xtFgfaime2JhdQ36hAbiEdICiwQkCC5IIL59J1mDcKcDNgW9B8zngJzLGvpoeCwEvx5U3RIR
oI6L8H7CSw47Ely5k38MKkw7erV/g3NYXkzzCtladpKBaXph//Q9PHl1yLVbXpNXVYWYD2PXP3Gb
bs+PVQD5J1l/+32I5NEPqyVfQxXKg6LESEdkTiPRLNW498kWICVs0s3PT29mcFVDNRLVahf9IFAE
2Fu3qrUlvsWKJT3SZumJqZFcsjJGlRmclfQY+OOGI1WE5mNnlSA6QB1uaR6yV5iu0xbQ4CwypnqH
V00WG/sLFFQc0i7GMiT2H0zKa7EBqEybjdxrhyy0M4otWtffe+nxtRJePJC4cyDhLmL94MxWZeVN
qEwXB/8oCbIgVPKidZDV+YIlX0NQqhwvBxcn4TiCTyFeVKJoDCpgx9yBBNOH9Cj0u3msljqzBcX9
f+EgHma1jE8EAy5wn7sLxpC8yrUxFoxwVNbErNq356QU3/841tjIe7VKNW1z4ZUDJu2kcs0i/gkW
GpngW6GUhm05cyzFgAOAFiLNHFZKH3nexobWnC8fIkHSs6hDdANli8YbaiemWFSk33+1YAQkvowv
tZIgJe+/Pt8WpoGmuijrvKQz/+g9ri+6ESgpujI711kZzyIGtJWifZDwxdMPkdwsmP15FUGUvBkK
1FiptCCrcik5FTa24Zqy85DH9uFNSNURYk0VAzOK9+88HroysnfLTg6J4SiJ2uar4LwUq+DEPW7j
xeLPnVnLCkAH+vFp7zRC3FnlsNSgGoerUaa21lfLcXBxLpIBw1QcCcFHL9tXh9Jk+U4wVY/kiwy2
9MPV4ykG83aN3jRPCuEL2Hz97oP9e0JkuFaPurroGclRX77b9M4ypcWRYuEogPlUqFw8F2p/2T/t
0A1WlTRmxTMNU88vK5v0+bZCYDAEZqI1SBH5ZlKi221aIFs2taILfFrRMTyjD4Umc5wYwp1Ifo7E
QRgk8Ux27nVxdn3No3TN+FiHgLKYZF9LZPnHqSe7VA3yI3H+gIklnJ6TK07i1OqWGRYWmrhr7f3F
Vwb7Rfusx8Sz8VbwQPHHWXjpJDOPf9W0NvHqz3kG9R9HbJROzgxYjPo31e68i2jKlye5qR8Px7Jr
0J/+j8C/xygp4uz4IknnfPr6eiGlksbkLa0RQPq1MAT8PRQwrrwGLZwGAWZycOJv9ja2w1Jyh0GT
Ll8u7wD5kvPu+WpeqnrkG+h1m7Xel/Ay8uPsFRvelH2CNoD0UdsBPMKtibmxmC6wI0SbN4mppwp/
cUhMWmQDRgV8+rZMjKhDUIsS0xHBjUq2NUGpzxOLwBg7AZC0yeDnn80ZwTrL3e0OXdaxwmROiErE
3ehTUmbVZ5/Gujm0dSI+pplhXJRH9rhN3j+3wMq647RxeMvo19EQtVSozzxgfVvvQCBkXEcKvpSm
j6vq/hAS8YBs9xkSu7dK1RBfUgEKAdi4jc83+08rg8beD9o5Ef14Ao22B66grn+LVLCVzTKBZDov
S/CTxLRXmF+7/UOJODtF+BicrD6ZFtrBg4B4f0l6EAc1IRpsxud2bKLuQMAROTzjyvy9BL69RXcu
lBq6tJioVnX/1GuhFPTyWeW0H9U+yBYO3bQBJnMhM1vUZCZCP8kTt09/IlcmzJYUKkjnzHh30yiL
7pl42bb4/Ds/t1k65Yeh2VJdDyg8K9Jjzxd06mRArK2xc1xT/xd/qyupwSiSWLqG8+Er8qZg4rfl
3fVCmYta7+BI4/iJgrWFFC8plz97DX/5KKo4nloekfYZ2jOziMEadl9/HGsAEd9+RCIuc2GdsBCf
yZ4Qvbq6Dt2kgVNejak0APre/2E1oK0SptJJdcCA3jjcVYPzCrnDjIz9BJ8AfIb55FATp5L27kEh
AYBMSeqtuCDEzOACL82H8MNfaTSrTIEgSAlxfSpuMUNIwkpcFFDHtaGiGoyapv5VD+XU+CeMRjM/
snOIuZKoaNz+GJhS7K0EpAqyh/Q8bk7o18LXbg8KxK4chbXmvd/fCV2MiQ66Qtsm35vxKFC0tqDn
kvyrGiq9MMkn+EnKVSIYWgGdfuvpVhn3rjVoQaCsRI1qMrKPZLwaf6CWsxDrfBOYMq9JgFwr2Le6
c9SaY1XhiJMSjTLAO6mRWU0yi99hfnb5kwYNCIdHa7sm1CYGg6gNbqhvDm3yDXHdHL8gCsI35jri
WT1daocnacvNoXULygvUH5/mHz3JEdldpELC0Sohv591H0Q7z63FyzLUbYhg6yS8jZoKKv2IelhY
+00HtqpPnCk5Qs8LyHYPZdg3opn6kCpzn1xSNDpzpx2tk23ouTv1KTgsEs2Sg98iomAjZQIUWWyX
7FAwaNlagzBKKeBi2077Ep4CS7i6JV7mtx+teZ3pxqUyGiOPnv23uqZJBpklQILaTBwPx7GmX2us
5mUJCySpKjgZTRYW4bZZt5VCNgPaIoCdMooTH8Zjf0syxndMVHhTxC5L6I53EL+kWQdth+LTPv1i
UcwTQmPFXiWIP+2jzewp/hIpGKw1e+IQnAfbHIt0zurvi/JGIOHrhw/z9VuSb3LxpbEyzO+iw18j
R8BV+w29ZQfPdBHsYQR50icCsZN2aLGc0mCzgABy31LYUrJNEa6B/8YPSPxFk/+WASZvCDtYF0f/
LD0Q1nOB6Vx4DeD9BAAuek+e+HaVrXXsBrhGwVf0Mp312hN6iz6mhTZ8F9/f0nREDeLXN/czescM
lqfkQKVgyVyzyUCsNvAsSivYBB4v6vRYxHzPPKsSSvcuRFt0uiQAiRcfCT2Ng2UeAoWzR+Hvxlxd
MBDoF+Dh4MFHiwvS6Le4KcIuorB6MOtsVOPkY+60ny5MAQpjulZfSzGr8r9kia0uKCjx5pUalb7C
rfZf2TOt75Fcu32Wz4LWkRYxI8h/uU1UQlB29jqyuKC712wuqTfTJ8yW3bZ2iQOc/cij4GkA5+ap
fgBfEb+PreQS9Nzn+BPSxQ3zQZZ1HipOJS3g2HuabpDnwfMyEH0mqkma5LdNhGdo6dChPO4lJQTc
ZbMIXD+rEV0vh7A9i/WX3EUiSO1aMXUtOIWiEw7hQJZ6eXNyKMp87DTTJfsY2q69VRgTt9lOpXy3
fIePSg1VHIGMih7iVyssEvI5EdWuFjEqFTVKj5ibywW87A5CWROq2GDnwv+ilu+3U+mHXXDu+V31
kJuWTs7ec/+S6WyauNvWiwLXlE8TgWsuOkfUHHiBZ9LXCPQPI0Ja++2ClgkWk6DmhO6lUWcYoRgI
8CHhFMFv26ThB11PjDQoRVG2Pwh74zxojAV5jjDpETxSKhWC9Kf4fEubZLFGLHqPGdzyZHyElvjm
7eE/nWrZNSmqaaT40SfTWPXiLI+UJ0SlIc3pG33L9+p2LMJg9i29XZ6slyQAg/oe2MELPA7/Jlke
JqOIfM2qyCTl2YOgsNr6EwkIWCKf6uza8wDPzJcInHIwKFLPO5sq0n94BaO6PrMLg7/RioVVVkrl
LlsWubOkAIYzJDX90nTsL4TkhjI87BrnyJoqNg5bQB832KWk2F9rj7CgBy2TSWOILAsHlfWGZeLc
fRpEQe+KYhsTGoItbojje+p2SiLSzLYVmpUEo0r0iCtYn82bF5uKIkWfGMQEJVnrFBcc/EEB+GeK
xiDn0BLpdW1qQGaZRIY5pEE6ODD4rTdd7dU45KkwFWpMJDuRi3pMvYseHZbNE4u3lhcW4qNkunk5
Tl33dlc3C29p8Kgab7IYMJfNFpbczwpSVBRAZlfccKmQYHXAKCxgbsztsbkSAu6sz9/BKPo7yEux
EHE5vcD+N6fJAtiF0HvhPN30y0XCN1eCL9diYTlIXlK59Hf63rEEIXBN4tTSrDYHg4vSJebktDO6
6Lmm+oFm9QxaDPnw2YSF7VAIRmudEwCvneO1g/dwDcp/aeBECkS2MvGQmftRmsc3CjxiGZeBRsnW
DicR+DmdChI6hceT0E8ezm088kf7i7CIx33Q8wYNDGQ+U8gmmnrU5twaUGH0okzXDLCwFoUfBRQT
UUR1B7CJHGSYIMYIdr3TBrA76qRWowrJCJNNIv91/10lOZ74uDhj5t9T6HA6hHIPizmFAH9HuKdw
5RMJmuuAeZfFLgjPXVkBo4VY1qBmw6ytLRhj371B9+U7pYNrWhTYCi/Zf+GU4iz5EwzaqgRDL5HZ
XswUglG119iW3C01fQHsOzFh9JPfT/qNVkrwrNYaPinBOmn3ur7aVCr+CbC6DH+pDovwpjwNA62O
xZRYDuW515QA0Zdsi7q4qsxJOliUbbIA2a702mmdLp3itpvOtc/9ZhLTQUQkIXAxemy9H0TO/1WA
uSCw+0UPUVVpmbX5hT+ys1UGokmrNmq/5qr7CRw7MWr6Gc3bnhRUb3v05NiR0lXuGtsMy+gOvGPn
1sW8q501v/Rt7ObCgPT6YnleU0gytvD2jz/TVmpnc/2ygjBlE06D5uz+NybvVP9hChGwrbb8vy2x
PNxQv18rCqZfFmLHKe3or0VgyxLT13SnWCjoZtc2egYxJqM2RnJHsZ9FaOAZDXe/7zzkenkbcIHu
tY0RWXsalkuVaDtgThvjMpxLwGPA2CUvqAbHP0LCO2blQm65x/xx3vb/waytKczGek2Jdlo+Ntiw
GPK2UIwACleAakGBTP2Y36HEP+LTSjuCTwh0dcu+/qsHRJUsR7HTUD4heUftWTa47+uL3IRsJNc=
`pragma protect end_protected
