// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YZB+c6B2UIeCJFgAjKoah7IDOq+k62X4pl7+1PIpe/R5h3uJ+T1q0MMkvn0945Hs
fo2fX4rMpOCN0wbRJ6BTgbehXTsWd5hao7ve6hjauRo8wJPYVlAu33PyMOfqrlxM
iEPYFtE9Vcx/C0Idw0qoiiYr53UTVxtC9JcvHczJReI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26048)
gSygqnoS3Hfy6EWbj5S1787LnW8953bQQ82HNt5gG1N42dqJN9BzTblk6wHnvSw7
iqiH4IDjXdEgC7foCQvUpvUTREbRFh+xE3nT0oTq9LT5Om7UOERwud8jV0gGSh37
qWxG43BFeNtiGZX1lr9VLYzhOXV8zGZKe3m/A8LC6I9hx0FtjJZRqFoScf3IZxbw
omEhkMCNRsxadBSt64xtpaXtXCoJEr/4W4lNZek2lS0fqU0xr4vnNozWZChnR8/N
ePKUgsVxlbdINOsfD60EtoJ65DPrpsQbHMjady4AugYC9z+asutCgnzOfGCUTMFT
cbkl5Se2ZJ04dZGIt+xb0s7s58k+TH5vHY2vMgqTZOU6sRWQQphoajL/QoLqxDgO
sxM80ZKN51AQxJrkuM+6orSv4ZsmdLOdiHbQKgfX6TQbsfmyrMIyECXjKulS5119
UEMIHPRW/7uZ6VcpHojylHDOjddRxDSL00pLiuQj2AhZ2rx2spf4GXUnbJvkRlFj
yKNJkyBmJizTlp2H5uv5sylS/2kLZL+JOvB260NlPaH+UUpySkFXbeZJSXe5/1W+
KuiylfkWRe237Jaw3g7G0lWADQcVukzckO32xFWdEj76JBYe9tBmSGA4DNt33ckZ
9Yyyv/l2n3+T6GY1kDVAp/NdQaKoF2W5FnWo8JpNHSqOCrs0V7IaZ2H89vfRPtVV
fKd5Rzz7Ibg8mExC8GGJblPRMoYde+U2FjhDRV+z0dM0eP2X0VOwRyyq1W5vR8mG
tVzADorLtnM5NhKgaHZR9KibibqnluqqR+sJ32I10qnG/xONm8xyByN1tJ4BthWL
HucgIEUF8zW8qEkmYv2zoGKAyeFh8+AefIfLSqg33oHEd6wvPmmZafzADYMyDkxe
izRNbI4b7jFcPMDp5DDJi7hlVlDWJ4tXCdQ172hutYTDKm0YtX82ypDcW3RXKef/
hicTcvDE1vmA9WVZCQ4jQd5c4UarsDNbVr5fcIAyPhHyUluXxu7kClsOtyhFUuCc
hZF2i+OFm/jk49MMoJxm+wxhOT3JpQKuU9XGVxc598lUgT6gisLPU4XYpHIqgdfv
iO4VqjPdAGiu1N9wIZDtrREoQbBBNa0SdHM0K7B2HzKyH7l1ZBymhpkAlKXHW4za
wPZL70xk2CzSlIdWULhEp1+KhCWKh3R7Hiq54cMgXhYDCEwIdNiQqYCFyExwOZs5
ZaxcUEPUUCvYp+gzhRfSGYihrst3cW4ceiZx4uO1oB7hAOZdz061oF1Sj6DNAvTM
+im6iYh1Btu+FAZCZSpZ2fdk8ITToZZIopmnlN5n2v3C6CYRe8ouHSTpLuelIf2i
xB3+c3daIoWYSyQloWfV8sV6jYHBGiiFZ18+FBYRV2R/NIJKjRYsbAaX7g7Kl262
jTYLFyW0j8nJuZe2jGUNzHGZhmlLXaTtHHAUaG1w1ac1DiN0Xs+D752MqlvM+orc
G4RA53arOr33o4FcRuuFNwRctKBmdgQqZRC3YSl6UIrJcPbrBMr7G+QgG2+FJW5V
ti6E/BmmK5WF8pUi0fGjJwS6jLhukv+rzVpxQxRjCYnOr1hU9FBrpIuRPI3O/wUl
cNE2oaRVV1cAtX2UP/M5lCjDilM1pqQyuCAOl/r3CvCq5YjSVarGt8gp2Z9/bQ9Q
UXMLrLhT6URfliWe+s4494EsIb0YoZ3eKASFOtWz5x+yaw2yLo64mjFLGO+u19Rh
Sgtu3Z64oX3gdoiL9UXqcDCjA4QxOoGeXwlE+SKyP0iMe4VHOf5g4XnXdquo4HB7
iTFEQfqnwj5U+GZZJ+T1K9jq5Z5QDQV1nqcQIQbXrBM8NKeHGlZBcmn0ld1iLSXK
Vremq4uPzqAM2VBIzumN4veCpA4avMPG+BF8+PupbSXFdq+eeiNf3eTsitNoNQ+O
JzGDEASCWAgomGzLvBPuLrc2N5Xb1pEsjxjv1rFNdp0wfSX5NgrlPF5PNNsriLXJ
vUd1YFpL+bm0xE3bARoOpgiiaLjrD5xkylghlVzcTkQZlrVQnlwIs8c5YSw5JyG8
RxLSiZrfGQQarI7pJHVQ8zHrSBKWf1NPAMNUIl0GcQcmMnP1GCE63uJX6lhAvMBc
JNP5+DyDT+bMzrFQ3uwYhD0zM8dBFeG1QCsXF1rd1Ejqh/eszht6wHE38KJDSfzk
nlKg/RgBAO9gHTOE/UyEl3cXZ0IvPOd8mG2nmm+tNpm7f1g4oKmYXAalE4GnKqeo
kIz069nSWPel/L2loI/O084Xc7kDLcsof7zwN0rpsageRsehV8MV4WDUtU6KzJzA
HR1gp1j/68JvpkRWhRiomBpIxSgCbiLYLy0lXa6c/kXoWD+BhmGPybesSS9U1d9W
LS1dzBOiOUy59TqKkQlhqCB/q1ldTXZqFaITNRlFQ8DzZkIKzCHZx2RC6AM2DhoA
2yqbPO2R2ImgH+z59qGFV/HADE4Y/RwkgQfiRSbW+5AcGeTwCR3LNZV4M9Tzm4Q1
iETF2R7F6zZ6losNylCG6qsRf/+LlpGpnvBw9bFYBg3p5QRX4SLfQKJwZ0G0ZTE8
grTOGPmVv5h3Y1Ay2GAkpkHZxCXurjYUlxUu83jgZF2LYBTFZ3OFjy1Man/Bu+5p
CCE//MUvY9jY/9ERZKiXZwdUGTRuaJLJ20HKh3HaVMZICoHnTyAn4SjA+XeRgbm6
XcwrltK62UYsrVw9MCury//shrCbF861oMbQCiRxwotW/WhHYd/2riFd1/r0O/xB
aTYQ5EKKIO1EQQp+HSGU4Z6sRsHAxEYlvpaPSmZ8NYc5v0b34kjDwoPTOsLuR2yh
gZC2vymYw4lzS64HC4oj9RhElySQMtsTrLFtKTBRxfhk7R+/2nRIvwkdFGloo8JE
A8rFj/3V6XjtFS9s1sD0Zy9XAxkzntTFjE+9Wnhe5Sk87QDQS9j4yk8r1OjlmS6F
b5a/aMKuANP3sBzIzQQF7OpfdvnhE46Rgza9JcPlM55sXn7Xs0oNCJVXgFU5v1Fc
BvEDogTFd6AvEXcduLSipRJaZvLh/yS4i+QH/9GprNfcJ+iZiQfjwRDfiT6xTkfw
WW38w/+AKdaCJp/WF+qRfPGbI8qfTXnei7P2oFV0zsBD4wcXOD+R5Qbg6Y3r8FEm
vnbdZHwId1/2t4HfgddyZwZzE2TQylWu+WMjhEvOEzlYoMxcdP1/1ojfwsiAC3VP
0mYkh/9izY/2xAqr/4irqNVT6NdSBF5KE+8chB4Tvce5FRFvlgL6ZDaZGCABhp8G
dIcqA+18uVIbISR+UOwgCF6zybACJuIRgttiPqq5jOrbHBDh9u0AT+PA+nRMLnaF
V5gkJxxGluCgjQf8vQmesm4lbs4ESG1u50hkAU0FjQsMc7bgJBfi4ZufCt6kxuYn
LAHl838G26mrGxtwLk2rxeI131iVFphWwnq8ni1aSsli7771169LBts+dzSBs7Ho
ZG+yiPjTz98ZiDhLB5wvfYJLoWoMskgTmAsa1UcLF5pmuXjcYCGC495UYbeilTri
4L1+m6sfH/zQFAAIVp86v4kBRY+/sDj/AioV/Xj+BwHIvJvf2o3yrUqex+i64FLv
SxJyjOSl07Ysvnjfnm/7FH+tiIXegtbzhviAokq1SU++Bf9IftoF2ECZJ9FtLArB
FvQ7uAL73F/sRd8gTHkZRvUBsrbM6IQQy3QEq2p8CpRPjpjtDhnMe/emWtQJpoI4
fHYxzVkHCFHQw47e7v5AbyC+s7Nn47wnWAyouYAJjgnJQPCgQLXnklGjj1x4wok0
UnYyOwedfn37U8ifmBEKt78P/5Pxp3HSsWsJgQbfsqjMJk01yEFGRiTL1sWBI5pH
Y69M+uFNLPvHBaZBgjlf9nFJUHzlIgMj4CU133g87TopINMFY1pcd5PoSD17Hccr
qxiW2O1yhKo5HCJc8wWuJHzraSCrAh6AhD/Tf+JY18B8yRO8hfKYHn3lmqdDzapP
q/0hmTIT9S7ZI5vm6/XnXHpNCSetafPXgvMk3IS7w+Q3Dos3wdozWlthCnqJPgyy
XADOMAqASWQFBSOZuUVUhTl+JGxzfEMuyPDi9/5e4tpwYO4TRO8GlrG6G3H4RQN1
MBD6LGV8IpAiBGzEPEszvJma4tdkVOAmWVBrcebPIktgzbAX0esVOeaQV6VdT793
ZEgau/f3kmY/dHKoUKfjrwkngKCGQZl6uspGP85IAeUf192iLWrq9UiHht3scysW
bdrqIew9eNp+Pl5qcmjx8QhVINqWImCvAE3YuzkzTmUK3cG2MyWGReaObP9ilPF3
OwtlX4aFC5TICtxGXdHPvjwX9/3PXbVHwSDDAplsHsIELENHE16H9OYF7x4cizti
cotdprfNovRC41JDRTKBpquyQ7TpL/LvlMyjaBxNooY0dL+ZuO2l7wnBPsusR/K8
ojJ/a8oUyZyn2KfM+B+E0jF8jeadUMbtI+5WReWIJ55nmADfmZvYwejCN5Qit6aW
3pVz2JULdqkDieiYobTAXYFwqUDeKkA0w+xPos5NrunFExXJt5/4rXvU/C2ZDyth
TRpMp9FkyI2qVmzcHkihZq7HHjij8z2rnQsW1A5bl/6LtgiiRt5z0nqRxcBwqPHa
S4RieJS5djoRbGeMLvy/VMbkAbBqqFblPDXpC0BWL8W5B+45e8lI/Eeudn8j4PbU
IF7ftt67wzwZbcqKNFBRvd24bkY27SzdFQjtjybvz12MOIIgM7qCnpSFliUvX4Se
9qL5Gh4R+LwvNBu5hLhf6oX3EoHrkPapP0DI0S03c5dDEd0YHIjQoRorJObyxQ+c
WHPLlTxijRyffJK00WRmTlJ++351gwNucmSDjnMzqBlkqcVA5Lx8N1G06QqOFIlC
maoOoNxZeSDBKlYpKKny6pp4oTRy4OU/CFqUNWvIhyJVA5uOqrDkLm96Q3sHmJiZ
euFI43Tzw+WeHleNtybYbpNGxzWPa+lBRymZNPN4c8D7kgW0zGAMi791zfMshoZk
DWNIni0Es7EjCb7wfQcI8MydtC33cTRGXvS4jZ3nhBxwTVI4XzlD9n6xvgxKib1Q
+HniXaoiDc0nGb0wI1HtLaAtidIZdnOKgYWKC+yKSfCqW1sOCudjf3gRee8eZqIi
iiqESyzQ21Um4SvckcHKDlIgqwjucOKxlQKeRa8/0olz6nGoWlBr1O53t+fxwHTY
pc9cm72WntOpVk+yUb0Jm2MEfAjFpWOVAUM3HwtixwLtaBRg1EaRO8z8EtFhCI4J
AdJof2gDGfi3SZzlg/3/XP4ISKUAVp1MPRlsHjmmxedd36IaczNC5IrhDS0TMfK4
pvhNeWv+QDOO0JqZ+sunHYYaJ29YeLVdGCFHIuAVUASQPO+/4ZxgBRxEHsrlXJB0
1BReomRTxLIgqQB0RwHWbGUxbWP5kUw3LvtakAr3izt2fXEJ0HsZRgbVhR9g+Vkx
VFqDY8CzXsbhlL5+xCp9yX0F6hXUNYnJJQx4yzZsJFsXqeTT03N3s/9NuFkY9BZJ
P2JPlwJfRnFpUKPOypUFCe+HojuTxjb+THRrN7xAxk7WEXz6MGr74Emab9q76QFO
qNOndlwiC4vzuU2jgrLInSICTmIbmL81J/D50QTlNnKtgYfNuOokSa0c87o4fHR0
0UJgxJA0z76l0xM1tMpK2jKgXgI6thav69QeBhl+/hmvgLdiCfkXl8BjuAUrQCEy
BzbxUy+oDXg8OyElZnDfiUKq6uN8xBMIS2nWSn5xEULJzvCLYWevtlU1noENqMhn
Ao4YA3ppPjQ5MZBCuAtjlUObcBHTNpH3l+D62YU7qwr1o3nEaD9qnN8XKl5370Tg
OHPe5pe4yUBExE2GEhOu7Tx7/ozcPeoPXcq4+MZMka8Lbk6IpscJp1WyM9pX1Uzo
WcxbyPLodBV/A7+3tYgSdh/JJatUJFzZ5KWg3/CNPPbF9v++KjLNP08hBKa9HVOf
76RW2dTD9sAvYb+iul+8ZunqhYdr3dOSCfP0/L8vnlYShEYPxNzwv7Zb7zN2s6gV
yo2E844CL6VLFWT4ahL2CMWT7v/dhl4V6zzkF2uOEpPt2OOnd3/ivSy9z64Ep+VD
WvWhuEnIs9UI0E/ttZENw2UX7B7WucRn3y+P51sXLmtLmUzQkxFvZi3Cy6xY6lcQ
lIdz/d6mAZFwBCYYQbc1i7zGcaHwtHIJD6j2xE31YRKcUsdej04CmvpFZq1Ud/ct
so8coUga6DoG1T+IdVLWfopiuIFVBvCqTfZLZ5TMLtcgwVyiNa3DY962DXYrFYwW
bhZ7H18DEXeZNiC0Rru/R1sCiFfZmy5yBp7E+5sKYiaFWjLiHX9LBHRUi8Gk3NOJ
cfSY4iWK1O65fislQsCx5SapQVq0dvvKAlVN8v6HCS64N2yS9Iw2EbB2fXwakdim
cf80vggcTX9cLcfcylxaqKDwZivCu49A6BGm9S6EDsT4SFZHO+OABRKPv4eqTTTC
H0x/Sg97JMC/ca5TiOYOT1HgL4lgQnIv3ZwdMqXRtjAbqNnecmsSiOMjcp9L+TFb
UaWtZlvYA7aDZ+BIa7XbN0doMPgWMMyM3tySZisNxi2JVjmhPlRN33MgrihFBLos
b1S6h3miIa7oJ/xHgGl/W4FAL1UvckIqW5KYwskt4WZcH/dEjjuwoJRXNN9vG8o5
C6gVwTIbXVWed8TcrZoT+LCfy6B88Vwku1Yn+/m5WrWwgGltI0NE9hlj7JqJimnp
PUl/dD55T2NZxtmqVyYjq3iVVxtKsF0u1r+CbCDho1rHCMbFkTpEI7oe7kxoiU8A
zudCwcnhsZxI2mPprKCwjiKTR2+0Q1Hrr7DFLYTEy40qeF5LV212Dl5NoKw0wflH
Yxs5sTtfQ2EbCe8LKuPCnaZPwHasjbemi74v+Wby2sRqUl5cfKqtsPOWtPjAF17C
j+axHN7qUsseQ2A//wE8cZn3Vwcax2SE7POz0qBQsEj/crk2Q79MDbjVXLTnbwSz
AS/2e1Xvg3TH94A2Oxt9Kfg82h8NoB0gAMx9oYID3iU1PCna5I3tsik8BvMf9N5A
lA9+j04+Oo3O5WcTSj6HCd5AxI4zHOlUMMHllzrsnJoG1KVdQw8jPUVisOsQMoST
NkDcrCCPFXw6EOXWRPijDy6sHh3LqGg8/AcvB2kMTUDqUVfewU1I09MU/hdySwDG
G2v3jwCUldGROfHV7hMKdEqMmpssIx9IS/bxF2J2Oy35xWSXatRXjD09q21nxKNY
j0/gyZGwW+/CxsEy52n7FGRKrX+EEey5m+PBRbNg536lc2fn6KbYzlm6ROCDol/7
8ObLSNvh8PxkTRWP36vvGkwc1H32CzdBSWwK1gu73pYnYHSwxtLxqBjPmsJog5Q0
v5FchTMrUkunC7r9qOSD2NJwRCcQpf//btWP4gUCXAmpV0m2RwpftsgzSYoQVINh
5d2xMg7WNqf/oRDqsZG+Q3SpFNze8CYLdmYt5BxVtPwhwvSpzjdOeGC4imo73X18
ihWOreRQT9ZMIcCEKvqWuyk67q1a2z725odYHBwQGM8rU6h7WHDzRWmXKo7ijU6L
+dt0yWADFRaHIc+8VXw+6yO5gFeowy95mYPOsoicxy/wkBsTNTESrPKAQwpz9S52
ZtNgsU2dkq53cQvqL3aeDIU72HIV28lbvO2A0/sPpin5faMyiQX0d6uFvOfsXmSJ
+Le/jNy/PRk3ihDkDCpPKsIvBM8GPtL3OEEwX5RUNEJjpUArqo1wfPrLjjdxO7nM
EsrT/c1FtzzTS1xwFyerbn6HOAvz8l8uXFSmlh1JNqMpTWOBbn3/oYfHwchhl4bi
I2j7c0GB3mVKzuHcrbOLojZP1TiJ6eR7EdFlV1P2MYeeqnBrT2US4XVUo5PfJGA+
kqzLQ5o5HORE2YhvjBcr022Dnp/1qPJRRj1AHWmb/kGDtXS6BKM1x911D0O5O5NA
ONNbfuyqpPd/JXVcBHrvRbTQVgic72MgekGw8+NIqT4T/yilqOeHgGANCUSPO4hW
athMDrRpbyRnu2SM/s9qGf57kvr7HbDOooPSMnVvq0VSxarRFxLdueslETEO+qcE
qtpK4lfQZ9oEsXeJfYuLwMEK8VbP9YlgVrhul+FoL7MVbUuv4P3gczLkxzfQNz76
MvUD0D2dt1cpE8ei0/B1U9bV06uU7LRFj+aqvnFp40ZxO/kn+db8+l0Dv0/x3PeI
hlcW4nTBknzcDy/vn+S9IxT4PDQiCMARqvLVbHqwH1g04QgC8cdn09XOrLFp66e1
VCLw1pFksK+tMjoddti8Sbgaz4SX9C0ouiBWCMuBhHxZ/grwXQrrbL/2jf0OowpC
rIbfVoL4PZI5y0Zs2KbKpOxdAIRr6rEvrj9qR6n6+LmPN7cQjv1UGHbwiYTwxM/k
+sW4Dg4VtnH1zKmBhsVanFKwEFYxCuE46YslMP+z5bQWxhztvl5/IAW6znVy78uw
2OXb3sggHcKUym5XE2IDZ18oCz7Ld2lH+FBxigjC4iQdulWcJvlybHxrr1iPU6s6
F+EGCVIWwTHRpu7ClhBjuGW6w5XtzlqGOshvvy2Q3ekvvnPgYpln8Rsxv+qGL7lu
ZyaszqR9jckId7EG6JbzqOaQrsPPhfW2h41jcBO3uEOcHccJvEJaN3UAS8yB7tTS
YPRXmsTu/i3bLLejVmmAFufU7YdrdITnlau4eYErV6184dUkRznIXMKJYMBjdbfe
PqnocY8NmN0U2KZPmbiFI9q50k8+93FBNKB4+Abf5/TzcJs/PDCf1U7KwGoGTeu5
jnaOwLgy1gKeCIdzV5C/Cr5jH50hGZ134Pis3bIzQqBNBI+tDjEGKdSx9LXbI4F/
Hwm9vwzEyJFA3T0qt65gOdIe5glD5/5ok91EBI/q6CcMDUgsUNd32xsTokwvDamJ
dbfHKgFakUQiwzjhfwq8NnPimJlLk2Uz++vc0hZVlh/R9KGXniP5H7lFY0FG28jc
dKR7YgrBdQRM5d95/a36ZFFbcoSKIv4rp8p8bOhkpxrKy/YfSc4ASXwPlMVh07mi
sskaUw2Ademp/hBjWH/eNC0It89aAhZ7A5d5ruZ+JjbuiOYiVMFxO3QnwAO1/F+n
6xHIOdRWQYGePpHIaVCnTRiWDvFSaTLkO3oh1PDvQTSb/lEEihHh7FoDrcfZkZ/i
Nw9nkHvNpVH9yGGnUZhGMyBdwQNAXg8WHRHZ0BA8h/jSkt6ZwxuJ+KwiVqt5W1+x
sFJ37dcCSstnDXR/E2p+FAGiJ8qXc3ZdzQZ0kdHaOFZiLkDpd6qljIbRP+fqgrLG
ugvW2lZcNHzoHi2BvuVpE5Vm0CEAPArHnXROaJSy3dzLAs3wGzCk6hyFqRBXW8Sk
0IG21MxCJUQXsVkEHLwrdAxrbgrugbsoRh2NdYlEh97beJMq/JQNjzpXZ0DUBCl/
1Now99RHWLpFD6Ycc16skQEOUJ+NSissmz+ZwaGv9rruKp/seuedbv748yIfFhtA
37IoekVL4zfetDC6weENm44wnmncDKSJyaJxgUqwcJ0aUl5JICTGIO2V0/hiDNzS
DsoYsyw8Kl7slVZLQejSNvgGNYXr3hitIhhieswTtE0sRB29nqLqf94F48XTqTrQ
Zo/QS9TTyZMdbqBjVoXE5/SU9xnpsYlQQnxczhSZdi0+5uQsbG+/TTwXGbmH/BOU
GGrcNiCPPb/NWTkb58hUd3PwGQQdZN1G3vRtUxZ/8yiGs/7+EXRYW1lpv+eabagP
TjaiSqVkm7JQyAX4ojnJ6C4XHCo4bUCoFGCh1CpgHsERNCuyBQF06NVMSmEY18/z
K1e8qlzadAjp+BcfXg8zFI71hGeHXh0Lr/hd/qg9WAT95hT0PFmDo3Go7RJcreps
MNF13exhxr5BlIVcIMkE+syPxu+q8GZGKL4s7+w7mNjmx7HnWZ3WGCyMlBOhuMla
J4EY9+AXV7BUGkhI/UMA0rCUdFwT3xfnn51NntMTrY9cAzZ7ZGnjz+l/tC0uk/2g
i9EHiAcw7T3jAiZ/KNnHPMNIZgYtKdJ8nXCz3cZtiKg3V8cXRlw8JthQjwHyNui4
HTq4rsujzD5XYoq/2+GI1qtMoG3gBPZ+jkWt6joeqsRcPmz7w1Fi4pxznnGq5Bet
cY7v0OWiRC03tqf7Ah9xqlifKp9zSxIBdKnVdtRWcftR6NIndGvI3L87O/Ntozl4
yRNzA4XJm3Xdij/q8z1Gg9zt+au5vNEOKbzQXIsquT+Tm4kmD/7fJUyOV6MmlFVq
XGSfXYjmJ8yGPMVECIRKKKk4GAEoEUZlZsa/b8JdUhWWhW2PNH/zguWyOhw2g9z7
gtx2dALuEVqlOlV+L5j9WLc/ooIU1MidvGmZ5YbRahFfqiGyJoyh4oKrmZdZ2/9g
oa+pENwmu7Ai8UFg16MxTGRmajVN7BeWljEl4cLEmkE6OJFaqIW7trrxUIahZx4/
i4hNmYMnv5Fg8bxPoo3n/JxUaWu8PrAzS5AT3K9QEhKGFiNgF1tZ4pFX20aoHONP
sKdNWAeOj172Jf2CtrPnIAQRpeKqrc/7HDelNdELgup8x0o/kR5aqAGGA/SF1/Pa
Adz3df0BBuRKO4xdVY30G/csvwoktY2BG7KpemIFrAAtEUiCmO9N0Nulrz8GZusQ
la+1AuaDAtJG0EuyLCj5YZ3WSXKNVop0E9Fna8Ay50X1227pY7f+I86fS0BWNfMt
e9AA4Dyy/4Mayqsojm7hs8wWp9leDKAhEQXQzopjIwFXnO+GUUctjKJpj8eIZqwB
+bkmU/KPulN6RHcxRhioTaYJTtjvAyJsIqoW5czWRPsSH4l1kqyoXnVE5cJCLzUc
cayGebSEiTmXI0mXm8tV4npt3YsvzcMnLJcyXGlgwTCtnAhsOLw/PH0hBnIzV989
30+JXpVIzuSTk71qfRm6faRrfJ99gAShy7jkqqC6POrQ94XNKp/5DPY9ZFFU9u5k
52wdarJFspsaJRDWbkAG/SmHfAL9BsVZ1TF0tVAvyYnvfBF5wSVgCzP6wrWkpGvq
O+KGo4I2cvTDZMWjHvedSl42Pykso0BTxByhnr8BXd04Y74Ied+anuzVUPCie1bn
cX7BmOpZjjrIKFxYpHpbbEAhaT82lXQbLA+eWlUIx9CBAYpjsKPrTLlFs6uHkiUy
I0rI3lOZAzwBWz2cnUGuYn6gNmiU1C8q4Uu/VBqSR8Sjgn8O8Ttq9iMk4eUlaXEg
4dhLzUYzUosOmSgSFWmU8d9MF4frqVrzhBvDTPQDhNmOfj+G4i3/DS1o37/FwHk2
4YemxTHiCow2EdB6cg6eel2Mc0rQ9l5X10ChHRLqPh/Fp1iIWkvJf9lQ1yPMEilZ
iArvwr+vI/XN4hHmxHygGfriXGpyhUjF3CxZLUsuG5v3xlWkJ2orkBgPFnV8KKqD
dLYgFnaHXIhgoOhj3Lc2UfqFG+qeCbZN3xWSyUK3SfgqIEZRkJmxn+wF/L93Onpw
vt2BNtS7I6gPt5HH4HoNvfUoWNUrOLFFKD7KeX4e1QxnmRtUFTQlPs8DIHGjGjxw
RCQ/Y7LQoJRo+2j0YjMS+B2Q5GrvMY7WbvFbklsGc5etHntC1jarAd6rJUQ4Z4u3
qI+Qzj0JqMf8bfjfJgnEPxFo02WHU0Kmpqa0q+X412/0VTl2qgP4zYsNED6fOUaT
/qPybZcKBLMAufK6O3FfgU18jtgGLoY8lZRcrNw3TW+3ivyLlZpEHsD13gCVTS7X
UqG0j86c1mswQpDPTzCrpxuxP3QjiU+fcEY3nSjDimgzQO27kdoazlSiEmza4DPy
Ameklv+2QNsZLlXRAh8XKb7RA3iiIFE/H8+bZGjlLJ6uv94DnV0aVRa8h6ReLv1z
XzgxiWopnQrTSv+rolXfN59ns6nxP3V7fYI68Oz9hb/99lFytWmFp+bvTUqSQelc
YNzQ3gfKREgsYxrm5ZrF3YsrZ39QemYMVoscCM12iGO7WGSwIJJ5RWODO8RaRdBa
3Wh2hbG47oi42m48kQqLiJ/PTfvg+C/oDSSgfIrRKZzYNuNy0RidXu9QLIB2f7F8
8+Y49R1LOlcYTMfN12g4odg5l8rLakzXRNI/Pu8W6qCJPhl1HDnXg5aU+B2kDIwf
70WPY9yOZoHHTbcHQmdwimCF1AwHj5aFqQFbrycTMVjKr0KoNZWjP1FPJ95qYGHy
lcGpJp9rx/RqyYGV+UVpDX4SfSbEzcIaKZ/Ad8bDSXbEZbpR4Asr/nuXr4Dy85we
OJ+P+55TuizVnkjsTCpftcRWpp/7mWAeXvd9Ch+n5ZH2AICjgAnCaqJ3pVffGH06
NWl0MOHZKbSuwpOxNmZeapHQvWmWgMG3sI77y3Cv1JAXrl04nwNrgVYzKjqT1Eb7
VmqdZ2/1OlwGmKIwJSm5GwdnIqtDJnx3L74IYYQ1DJgzwIejwqdo0NxEkZc2bfSD
60XpboDk6qTO81ROSl9s5teaUJfH4exVTWNL7Nha1MIzU8MvcXHEw5AkKuu0o8TM
jZwStEL+4IRQmk4nsPkhh1CF01KTX5HciasqikFzUk1OvsfqNGgcIM5S2QVPFLHC
ifTymheaE2yaCaAHMG7N3LbRNqe2im+T3SD3y8WL+HeW1NW95C0QGT0hezX0w7CY
SszY7f//pAH8NANzOyYydXs3BYmSmHUFjJ6cTz8pgcJWpqWh2nfb1LZABHFmG42Y
xqAKLnY2rx4IIp+any1RfompIuyp3GXgRUbmNdcJTryTENHVYqta/jgp7XeX49Co
fblclnRKs2SrODOLZ91r8thwAg3+jNW1JWQ+nKDkHtxfb/9Mp7F0bbu1qAajDFnD
75XtFZpolMb5oCgJaivzY5H0KeSJq+tOfcojVwCQ0qsxmQmx7Lcce2BdyK+ZG+5o
GhJqxemclyUc+h2zKD3slrAa4PK/l5DgnX6HruOFBy4W/HrZSegGqvpN/brwER/+
Xel472q2jCNawadUKyEtEE9SCleq/gfjjpBP6qTAVuW5Wmew6Q/NQ25VWXwMWM0n
z9zHtDc83GEOSRSdysEOYKDUHIGTOm9oUc0lSml7lpkiTPkQZYCvV59RZ0bbqQOg
SBh455j9lxGDHUm4aUFa9bY9gKXXLmMHeHoDBJYkidfEp0s8UNErrIcGnFlCAlgc
oFwpYLnc6b4m3F0ImkznyJ6ZpBDx7V0oOB02n5/gnjcY3fkV+JYmSwTnmYdOgv7L
ftkVdRbr54zFIkqUAEw+JAf7qunLbF7KMopFaVWqGvr/nxczk1bwdBqPWvXSvQPL
O1sT6GiSWSb3c/3LJYUaF7FO6L3e9SUSfxJwFZ1DQWt6n9qUQcrS3ZBiNu6/2/1Z
7xz4f8Kv6ztryRp96/O05fi6S8tcPbmHVpWwWegYYoH6RBtdcnzKcfPtJUSITdt0
Ev83DDG8MMWKorULRLPs+s8gO69lYdyQc7V7JInI5/9OxBL7IJ7VsieUMRcPMTdY
Aqlwm0afuU+10PbtV7ICZQryx4mYQ/Fc+0CENlZJCuNEiXEWXKjW5eWJHi+qK7gK
R/4VvZDfhVQVFjCnznDpm0/D1AJIRIQuv9+i79WAeL14FfGt+6JssM6RrKNlR6WG
E9NSb9vYWusspw00LlV6Z9KeVOw6hq100jcOEG92JYgUmD8aAEEsnfL+qGlLjv02
eB56aEi/EenjcmTzmJM4zbcCcy5gpRXOqsXDICCw9h98kMHSjN5FWakRnvFcvLTi
VGiVi8AdXMcshfxTM7N7TBDo/BkSqAoe8GQ11MTs/teiCSIYorZ4VZdkbg2L5Oeo
tT/YapdS7O3Q7mVA4JDj7lsaJnauTxs5QtAGlBSVFEWpV79GEnAiUs/iwEmMWyqr
hE75L+gjhO0W0PPtgimz/D9Stdr+bkg8eLZDF7ppkbPXXlNAEYBByAcrZR/6MzMM
i1m0KTZwS4KVjL9Hz4TGpucpSBQMk/6qsMESud7NeZfP+4ZSEu8JicqUprk7qlsZ
gxozuxZ2lqJ7SxEHSHvKXWEHNvq7/foT4CY9pkSLA691mw5sWxEyHZV9M5m+6jxO
6It9QzfFGcdnTM1NMvgwW7HiSYuXU+IWYOXYka3qKXeYrAa1tbwlAmIKvBwSHdcM
pUxbjDgQz7PYhjDzV/E4uuYHK3RFeKcN3xjYSKHUpvxSeP6GWSvk0jq67WeplTSi
X2zC7CZWo+7Xn8St2tFKYYDV0bOsYVyaP66JHL8JHQBvUOduaPZwQUNTAtWS9GMb
PfNVhmjgbP/Hyk3/9qsfsvRnDeagzn0FO3TIqKrCiSgZEF7P9dqrGatkfU1qYHgn
D3ar+CY8BQR3K62j2OimmDjzjd8Qdlm7TP5lHYoq5rj6vKfPr+Oere4YFZrYPvnH
b6RHOkqwEYwM66hFa9eGSizU93MfjsRJMHgyhQvKxf6qaVIcfSclN2bEUg7Bi+HG
fyv7raaBjTNcIcveTO9AyVoZEhiUcLGz/aMgtomA9MYdIZ3c+Ze1FfCrl+NqpNDq
qXnGN0ku8UsGf8OVlPA/jJGcXABii4aN6ItJsfwJcMJQxCMUwiS/b87OF/3HKTmc
Kjz6jdowp0VgqHWg54Go62d7K1a47NCKb9mCEr5Mik6pJCO+IzItdWcav2+vsGOU
BfKClzLFQg9UJ9bJ3dhzv74t8E7cD9E37pDW/IBdx56gHB98ED0MDVPfU+NHRSH+
grwqMne7RwOoE+9J+7DZaqaBQx+UddioIN2kubLfnCLAKb1jNV4k2b9NtUlsaM4k
05tzrZECbsdls33kRdpvEMcx8XYCD2DKwdF7f5HBCNwIiIbXBYHLVox5JCoeRI3+
pHElfKPzYdUz43FfpsCuhhYSbPEke3q6hy0NSgbzZDx9Sv1GrHYF87+OP1++YOu4
zdXH95kA5ddyOkiL9XD95FtI965GMOWkhMR34RTlO7CPhpiCzR48qC9vDo2ZZ1AS
ZzvSrb0R5hE6XtPRlwbaIYkKyQZfH4/nlNP7+y0nO6oeOy//Ui9cg/Ua+azvNUFM
3AwNfnUPLlF8YvtRMiroX/rfizvvwx8uK+ER4+GTWBLr2Hpf1AeGAXlLSH9YDfKH
ZDoO9cdxwASqGkFtGR9IUgn7Cn7MSbEtXbKkhnxhtEAH5XQetZNlpCGR5HSvy5dS
zuDrrLZjvWOdPDdmJG9C8ky80X+l8A471v0Hqpr04RcTj54v26EzXWI0HnmBYu1s
SipV3AzKbFbB4l0xf20ZKgp5TZSHWQk1nFcjqkfpStnnM/ENgnkKlfmZP30x1nTa
kfTl5wKQv64cRx4sz7cuUMzpo+BfbkxFiLd1ORfPWEt+N4Jfc6DS2DlWj+zx8SFh
KefxZ9funkRHb8mYdu20yDp0qHwHzffEQCBWOzv/CBBsH63VaM7CkK3CGIQ1iMru
d9dSXcpkQEFJi4hZRX84A3oGIacEovmERV1Dc6Tg5K3+K/XVoX2qcJPSMMtLoXea
PsGxX0Do9mXb+YOwcPKVQM5jfyGKSOM5LGFY9Rk5G+BUvyp5I/5CHzNzSuzUXzjN
zZzbML1xrPBwpwjnayJBjGg+BBqomQ93IKM0g2W3Ye+4h1SDKWWa6tX8Ei38kRFf
fV6VHeoAFlFCTMNCsX4lgloeeJ+qP4hFuEWVxv3Ui3bV4zmwLyKsRhCr1jQ9xsBy
ANU10KZ+FrHcnP48H7nmUrZ5SLYjI2AL2NoPGYSwHmFGC4oANJIORJ18wjChgBA/
n+2YF+haP0mYhftsMLQ8PrD+BIBAQWHvGc9ojal+FOpnqB2XVYlJc0g15mANx5SC
8qKwMWXGrYMMu4b76z7hlTh3YANz9oOPwxGtr+62pOxlGlToxIrlyJxpvmztcFeL
zbIpylx2BXTFPYWG5OJBRtbBDidGV4LxdIkZNNejcLQFpLd7preNXdePSBy36Tki
IGGk2jjPNTlpkPcnsbsAMknYNZ5ifKZgbLzCm0B/q1nBAJusyS+XsH+g3nf9z+HJ
foKoIH0crxUW0OFJjPzu2ooyZF3heSnmz8iSsAlorXrYEXqPtwC4nDkiLJ5MbITB
RjHAD58sU9nctzVZJm+vjQbe+rE52gSxzKgPer6NrvPsrI+kkYqgUosnKybONDUB
vpMCjNl1bqDsuD8Ti196rERCTqOKvS/U0rF9/e2A3bz2zQVv0tRg1hK2vIIMNCGu
mg5DQ6Bm9b9ODsi4s44dl++s1sUtfAmAaVWv555qZn0Hlgk+noob3Rm3YVM5nmVj
7CfhxYDYTWklACdMR6Ak8F2F1UYE3z7tlSQ/LEGFYdnVMsVgRVm2I+pkw17jI/Ys
egnoCnbI18IjcK+P3LlilcGQk8JOpDadUqQdOzAgsAWnqGJ4fG0osDsOujMk07iZ
dtE/JgfNPvYgiRHdXufsiBtmzvLDdihK9/xI4GT+ZBydJNgmAIEqin67Z6M05G5O
bzeTAqUoKaiMMasVDenvZOax3IHoQkn6ku4TP/bl4I+GCeHNDfOtA7tsopzWWsry
3cGUJ6+1tUXwbWA6z+JeboG76ykJMuinXbNO2vimsvJnVNjANDqSCoHb5o9MDuHJ
lgPFSPQ458OmUFtAhOuJ54tdYwBNYvkjLXNloJpw57lrun8F51XFr9K+nflXsgbb
hTsL6LpoEtX90qIR4Yz01izrV+4tt1cQUhS9VqAmTGPek2URcwE+8J/x1szDfyL2
IRkYPo75kbTGX7KtEMzpejYCdsA4fzJnFIj66+leaEEONkYJvTeJGKGMvavZ325U
t8A/29/UVnQ/JdJvlUgymg5dXwZIOUvueqavf9UmSOPRPVZ2qz3gRK020TSm3GUY
VVoDOgSa6QT2HfGxaI7ZQZg7LznvKt7UKIhzPSYlRzGTpIf3SEnwlsfloyhsLev8
tWDnI4ByZ1bRhJw1v6QP//tNi5Yhq7gHPZOa0i+WYmEydfV/wIeysZ/xGurkT5kK
5xhiOa/KQXYzC/bXQ9obCkOaqS1m4lOjfzLw3wYSeIUM3iWEkP+3DUbGe4xi+w1V
nqe9rA95hWL/00zHE4Ew1zQ6TFACBkJTb+6fRb3/6UQhoG57Fg38StJI0cJa9ymO
h7K6ijLDr8DQwZnb1+blOrbvbyJvlo/L5TaDEU/iD2c1FpLjPiHiojX6rIq3KVwh
KkoX56foEZ0we/vFvrRoKii7XUC/qnW45QCYCtEsu4P9/Zk8nSvn2//IwuCV4ONl
Bn7g7jAAYYtQMd+8HXqfCVfZcTRqXx7f1tHsf2JQIn2bu20nRCOTMumzdb0JknwZ
cICagMiRxxKYEzhHckC12KSOqp3e4uf18hztX2oTEIThA7wQuIzZxPubJ3KIQ4gr
J+SMqYNzo2LBWVCvrfo3u16uzkufISIo4NjWtIiaJ/J8Xq0m2Z2THyiNg15ySG6A
VMaYJa7sTCKdF3lxXv0j/VabuOFODte/K3/aa9fTEqZ6LrvS9A42OMjOFe/5IuxZ
LkkPY/T4Or+GfS4qMu8cv1bRRqxVaWqkfhYSTTFRNRygTWAgGGm8gUKfJWkzyQ2e
QZqlwMmT8qqhozZ3Tp2uwOIxHT/Bd9TCoe9Y5upB6b2f8B/EQgRLFBbsQ1jBf1Lf
kM2SkYNhOAr52GqSKZAGvTkdB1NGUoyS+SsjMGCr1613zVbWouefIIC8QocTLggr
09ki9wchK9NJhrhvPFrvKJmGc7tHJa1/hZPYR9hpfhvbT+jCS1JNdSyWehIqEM1c
jmIqFhTpVnKUAKap85KJd1SkJ2cm3dG2XES31JXDCA/DtujYEDNzX1Q71/xHYt6r
oF1TgSmKKMtr75W6U2AUMsUh0fVq4psKoAxz5NroettH3PnCCwhNeZ61oeXV/BGJ
jKTAcLfRGkCVVIBhgMk5muGvb3W1TtXqlJA78f/t/hPzt0FwF948f7JSJwKfLhkf
vMnjoJvDhpx8ebEAZXuMLcU5KT4HNuM9C507c+/zAPdSuD7UYbGO6eUJvPvvQWpb
LjkWhNurUdIgu2V/CTFUzOtiFMpdSur7v/+bl+L4B+zsjJ/9haIV+nR+fluL0EkR
3s79kB9R9ZRHGJ85+JiYz3HWY7E0kYgL7fkIfQyBM8NRFnqfnZR96wHj4BzWga6h
/LzbexK3BS3gSiEHnhX0XfqxHYtgIfWvV36OX13BoeeB6rkBClK9DCrAGUwhKKEu
0w9YgKTVWWVd6MZH1jUmiA01Ed5NhNL/jEjwnqMWchLS54QTgHd907KqzDoCNJ8n
0LHHFG14AyiiQHd2UFnAyBpK0QU8uka/9I6WFqar92DRbVtyvLveEjnthbgHmcnp
J/Hm39W7gCQJnY1rP0n0ydZK0ibEikyDoKXLf6Nkcyx9To4Wj2hQsuagHHTzwG94
5XIyJhAhV6dMIGG4pPL9B60JSYjrj+yJLLtE04crFTC0JCPjlTJ9SmQiqlWM0s4B
bfxUJZ5BLOqBzFaEISvgw631mG15KTo0wcXiJI1FyYci0S//RoDizZKZBpcoOvRX
DSFJ6zSjanDwWEn1ucSotIG/l749sdEsfotGF4U0jnFCm8CgtasGnVRTAxHfx9VJ
BOJ0nBSK1fCu5NJHHyBAaTbIf5z+t3UyDXcCb7BjtyTQydEt0gcPOrXEtlDCh4lY
3kkOw85Eykj3JGP2NJKSU6ACXDkegu4vxZ2te+fFtw95zDhZlEDJHYgO5VcTLFtx
WPryjz3CLsh087MvrvaZKU/hGc8pQsa4NYWEtWIp1zCVlbiTfiHJyyUbJy94C/T7
e3JilJRnRsNDY0raGR+L56RlEkSPc6EiRJzkU03xxB5hFb3yIMJhcwJsUYKvmvl/
YufuPrpM9lehknKsIMwiEyTpf0QKP6cllP9/7uAdA0eIy8yY636OzU60lbkUR76O
XFGStoOJ17dd5Uac9SDCsGVoavUc6qVZTlJ/Q1w/BRELvTvghLG+Kc6Ivx8nU+lp
8RkN3YzWzbAi4cgEG8B4WGkh0FF5puunZDLj+5WhvzC8/XfcF3CvclUEdmnxq03L
Zewp9a1cGQEzmYx2rRPqruNS96T3yWc+B0Ebt3YiZhv67pFfeOAnswC92u33uh+h
/GS7OkfxEGoG4BxYxM7pgRPBzU2lf4OhRyUr23aQiCdFq+frLailGZY6dE0hnpg0
VbDBS89ZSmbnHsFvnN8IyRYAX1UnN04zDa6qahDsgC80grWu0bjsoVzF3AqCsvwz
qICxI5CMW5FHbsuUReAxzzmP8orNfe0VWa8v5/ugEdHbJ+9CUhjjHXDQaI+DWKG+
4pWqqs6aE5SUJQKDG/SwVJgMfAAprKffifhpix9uJAdb9GHafKaH0VjWBP8DlI+U
+3GGxUKC+DMkF9eXuiPWik9laXwRgQSBoIMCCKPzoYVf0hRHrOb/7ocjRsXPIgRu
+QZ/0cq6ztQpOvnez0gso+3vVOr+HMVbzMFok3p9MPH+sBtmREP0Ax/DizkNyr6q
FAZbxg2JsbJjGw5WqqW57yQKvEzbIDVa+TgBXHONLo+y/TCMRf/HN1UTkBSYxdIH
VHYHa1YjvKr9/d0Z6VPtcgSKAVcP8ooA6TmO6A6K4imG3uOF3cevKyFZ7uHo0yJj
OGRLUxydWuNFUHBrfbE88kbbNGnHgJUxEJ9fFveeLzsILI/h8H0pC6Njm9luQ/Vu
djUBjxD3/dJT70DJPgMUQTee+ETghIVOMKoq0FVefdvdJVKx+hAk81yE/ulBJPzZ
2HDDqp2wZVTK1fPIVPE2lWqrI1BSv84U80bL7BIxthV/NhvSnlEqQAMiFUsoD3jO
L7qbeW3SqQIfIyhyo2LICle3G1nrfflSu6Kn53P0DP84mfPWp9BawxaHEtRzuWFL
vTGml5D2+kB9hxrdkq4GOdBg4Tq+advrIOowf644FGHn/STF12yVE5QMQtL69ljK
1x/YUfwAiVyS6fTm8nzmBoLs/iHlWlQL2YYpsIlENPbI5nsLyPoALAq0BwDfCyoz
H75sV7bKx11YYZfQlTDlUXe+lmDBL6r/1bPTlry8F8UKllhDgXiBCx7EK1Y4vqv7
CoWDZimJWpbH9NiBmLW2Gr4KvIZntewwm6/ADELVG3UjGOZz1Z/yUQFYIFTyUfki
3WwE142oU69uDcS49zlv5f0daS5adebus00OV8TrXaBh8Bt7pfvjsuhVdEh4cqG2
ErdXQGRQQ3i10sGKKyEvWn0zFwV1/qhMsv1appNDBjJR4omrsNeXiqwKonnF17gD
fpTxKhDmzPRcMAidfVlpMEsCFJaiYdygKI44msk4SrMtGoN0ynk6ncmzUOclGdTn
C2BEV19hx6mDoaUge2ipbeweFJNj9dclEmX6TcuQQANhfXhyAQEXYihxK7tALXJ1
tTFU3A+mSxyJGoynCoJstNM5vnEJ1JNV0vLRS8Unj2dFUgntoV02SB6ri1/Xg7mS
aj6elh+N4na+pQ/Vdwm+5fypLMeXpCBWI3tcgmbkZqMs+I50SlO1vjE2koJVo9nX
qZELF9MCeQR8RWNaOyXvt6eMFPI2phn7TePBuhe49iC0lV/Al4tIsTFgz12XbT7l
x3e+jmBfgcd57hyqpZSIfNnMjDq+CdmhzBU4/h46U5ygqJNqn+mr7gzpOJ1Mf1LO
FkkbSp0nIJ1uLCKfjZKJ7WKyhI3JtHVi9MpB01I8S1giHEJh5lNjIulsbCmpvIDI
ijuOKcfTH8phbmdSvOofdee4SG7h6h9Pkp6d9tHk300U1TojPFP4KtTuiB+ov801
11l+jWOBUn2LDtNxipeRF2+dHafDDDAHzPS+o2zuJwjkyKFrDNljJ0CnUA+ObD3M
/XkWZZeA7OwyilQ3qfWlT6NXk+wf96V6nV7FVBl4WbM/TbAFj6riVtUFaiyndW6P
foLjrbFZ5M33QNxDxp1Gp6Mjywn4qxsCTEUZG8dolbsoaDy+o8N1awTtEnIwauyP
UT+CXZguMSapAGdEhN/K0EUbCU01houn1o/OMFKaDajHHpZ2VGZVdNrBib6nr758
4GXQZaKXyW7jUP/lW72xc6OfpUzTBRGIYNwIXTWpFetRZtoMa9RF46mPLTle/BD5
Rd0O2tp9U5M2xIhE3s2xBC7y21AChiiYJ7lzY1paxPl4JILuX81GQE8+4wXQv+BE
LbkCPe1xQCuM4UsyD/IG8P9dV92icgkCqce7FsqOLDoCa/llSmt1SXMAYn3Z/nmY
sS/m6NCFvIP10Mj1q1GQvRLLrJTBwcOOLHokxZJ7/5AEPrFSZQLlLUGERkDfFmHh
LSc58E/iNcu/gjqCKkKE5JE6r3Rh4yDjNf9NfNM7iyFdEp89IlF726uuackykTXV
GXWQhfZqvFqgUEffeu4m4GrdF2JoBfoRju/sDU7dAd1k1lZXHFcyR/FqbGOJthXt
SU/1PcJ1FmxPttTROxm2hYQQi5+zIOIBoP1e8RNjZIdWGw20QJKakG62J3jX8Gxw
laNIpjcm+D0OcDJr0GONoNEstfqq+J6tx4eglP7OFrr6wo+XhqScNLj3ghSvKmrQ
qddEUGnQL5rf7MwVo0E2FLRVqpzQxBovo7rxGINH0k7HqSYhRETML/dQGhlBW+Yd
fTM9wsctLA8ScraVm6nyJPj4h7ttgOJjlBDfkdujTBDtYTu31dPtGq0IJ1YFD45I
JhdqeX8VmDBuXzCnr1fppEBmUiVyKXOTdU0WSMqRdykwEnZfrCgn8XhsD25DLir5
JQA9hNkh5hGz2HyTZzYAJLNZr4cdTPOkmHfDAmDSDwRiuzNYn7CxVlybr1bvMuIr
KbgZunHCO7T9DxXRNKt8+n1obEJ926xnNoBXcJjQY1sJxbSA+4WOrp/oZKnWTj8q
572S7yuw2WMxUu7wOkdEOXS2+p1nBe2FeSQQMyqIna5wLaXU07jMGhcr8xYgb7Mv
X9VsL9+9eltFcWm+hM+i1hpmRznvI3LE8kF2djoGIPawfCVDs4Ve8WPPxvCso30w
doT+SrM8A58rdFIptll5SrABVD8YfHEK/Bxh9PISjf/EKXpDoLy9f43UC5wII7xe
O5P0tyJ0lU+A8cmNT6LiNLbXyPRKwiqwdlcuKwqYB3G7SrbPlfDSCDKlbWI9TA93
1pait5xn6tLsc1U88OkxqhmJGa5i7Z8PJCMc7jkQt2zx4WS1IAwPHGKQpNNHDkRv
bW8/Uf9RjEPJPjmHdZE/q+bQLvMfBXASvyJTSwWHsggzu88IbB6orBLk9c0F9Txb
dBJuy6DmzP/qkn+iLBn5EqbXzjKgeAW0OsppUlWI5Ry7EHR8lzjUW8L4LZ0l3BC4
QOIP1ungcfrLLXEkC1fyagsWkurO3nqX8c4N8iv+NCH4ta5jRcjVcmXjc6Vsx+hX
L9BlLFffCUtLjnvaGvJeWAfnKFcPl6BA1AOIqIVRbHEa+ElCIU0oWQSmgvbr9Red
uiK08psnZfhAZJT4yCa5aGE8PnnRxCbrXhJId8D8GpxvBbTqiwnVwCKlWYcyA3Wx
LVEqTwZDN7ryu48BwyaBvEYDzH4Pv3BhxlrwTmqJm5ouJq0Phi1wECuJAN/P0YSl
W2WG50t8hvOdN2vylJVO21xiHxYQrX5KrRpuTwdjd5TAI+yY7F+LCoXH145c2A82
laGYBjWTiUZWgDI5pwkKBmrxVNp0N/I4kP2OnANScWCP7tcLnNhruONp3eEZQyAu
RBJ13RTr/S014F3sSvdQlEour0dl/THjtwdeNmzOf0D2ifim+up/1LVJydtyFyZC
bgM8HmTFRdjxohqX9bOxF97w+hnbFZ4ACljD9G5pCLq6DPfA5Igqk2yJ2vzj8a5A
Obk9izXz9Z2DNoe/NvMd0ADbpMkRlE88j3d5KmYw3newyeSQquU7XLDL+tt1+eIt
6Db077ATHHaPvsnv3cCrfkwxcUp4ngCzTCcq+9H/0f6KFZVg2rFiZV5PCpOtbtLx
ZRIeKEN/1vIlg/H/oHIu1XRZw6w6pXXUvgPRGHx4K33++uZ0p1ZJAbSVpTgHqLNp
zl5kdVosvWEP4pk6bp5HQQo+qEZa1bxyBxNT8bzOntFdLVkypfwwRD67pulq0zfE
cZB5ox/Zq7I5ckVIUslrZkr05DPI9LI5sh+tcdS3Xf/wOzfbP6x9TGRk5q+ZcMPo
mxSfz2ANlviNowtDYv0djVqsHp2HtFq6+XW11+lNjTnPb37PnwhkKg/FR9hAlX14
ZwOcjuMjurmmQ0ZOqsA/XsNYlflG8EULYz3wAnjIjz5q5bbI+XQaF4T3ESSmZ7Vx
Wxd01XcqVzxTxWnpYveCbB+RmGs3F9zesM4Rszq2dTMmXrZwBhH1SyWoVqopdCPi
6RS/nY4Pf193irFr2K+YgvQD43jC7E/vld/Uj7K6E7q2fKQX20ve06YIfJAVnZA5
SNCeb1ehBrFhqyakmOMicF/vJhXPIhrhAXl3lz8vEIdKSNoKMjZR94v/BTThObn4
eTQE5o+8eoMRaHOfdO42WqP+oLsxvekiLyLZxk84CMnPgMD81ADXAJrsfgtXs+CM
8jy3+iD1KM+EFrJsORFHc7ibefV1RS6ndGYH3O5Cb90BtDb4M3DfGeKWuRyzBxy4
JLPTEhDHqcuFAToXXuis6HA+Q2Kba0iznQbLQelOwx4dcWZ9U0bGHdnCJJHMVWmE
0bKlpWXCohkbujrPGXpc9UL34G0M90v0+fFrKxHhkyGmekyE/pm05CphE5Eqi9Ir
ikHGErg7rKG0nPxEjC0oCoL9NEDlJ90jHsYHgFoXfkPHG6Fe1iQY+Y1V7nCdszfo
n+LXveLOY18i/4wXQFWnOk8tIl2oclnzs4yxzqZO9jBSNwylt/wkrLUjOEbTYS7e
IwgiDSe3MdCJv6RLhWziIQFAWY9rfcHEh1Ol2neIHV0vUdrbloV3FRtS1O+5b12c
WDBFJyPDlPoi5fMi5NZzcYxjBqPwiaKwqu15bJQxF4t+QRHGZJgCjYTvQ9sxq3zL
bj06lL2Dk31t6qpLwYNPQ5mJQ675zl7j+bIeGnWwFztkTsQMWIauqcFforXd1A/y
HsrwM1jE1gYNL7At8aFBRITikdvWt9dRlf09Eck3CavBmkGPXhXkilo/EjM6o8VD
U5cLcKLjr6xvWRfIYUg4AKtktNJYZ+SmuzNcQ7U8BKZ0XlZ3mIoFJoYiPkcAQDYL
/mKpGCP+Eb1x/kgRS7NnMAUuJ8Anw+ramtufjDeo4oxLG9JueFrAHkkdsxzdZ+Ix
uGsTeu50NL9NsH26R97KfAmRAW6SypPzRyYLtDjgMrUN0Md4XTX7y+PiCsH80MfX
qPSw8ktLZ226UaqaVIqUmKXoiRciDIbdo3IeRW2lkCVzYFR7cej87MBnYza0l5o7
d3OMCz95/g0tNnblSUTdg90PQyheJVjKFbr1Ss61yGlzW4MS08AGijrodywhn55O
YTH+LV56fjosDPJLRDOLY28MnZzeiJgIr96grNEKUqx+ISE0Z5z8ti96bSBRm4sE
3zTV9Jlt+KVFrNnv7ybPkXtdsfa5rQOqvt4dZv7xCIl/y2DLD4WhTES8JTQbrwq7
U9nwPIgL8rNZNR8rxhfRqW1uQAxd1gXXGb8XqMRfyHk3mIHlOp384xoSO3Xx7Vyt
I1Qq7AbqiWPOYhOeUkBG7RI5BDVDhqx4IXZfpX0QR67y6oONBt8M4E+bghI2Jbgr
69Gbir4MlnZsPxHHa3YVOOpF3lymqnfecob7hCF03qklgbhHAQZBW4SCWgCDOKc2
miEh9fV6kT8hmphVwhQn6wWnH1c5PJY6pZ7MOYwGwkOsJdaClZL5A7OpW/b7zVC8
IpQCEFg/IVbeUSlEMuNiZ96QvrzDVJqSireFen0jPoJvzWj9bEUMrWPgVONDXO+S
f4kz0i68y1cbdQqo0PvwAc1NpMe2myRgZkIWpyU0Cd4HV5ophbgBvgGJbFVY7gZf
FHhKfvnnQdCzUPUGHwQ72Y8Cdxq9b/aEToZI+o5OY/Pd+QcrxZPx63FYss/OgKMo
B1jjjUVDCFCg+q4Li17/HQYZEUNz7tR9Oh9TQJCUS9bqxBvN1p5PME3eRr0icRRk
DHlrm/Rja0xzXLP7L2Wvlkpx16HRfUqaMv6L7hviDpM3zyK4ycihONroScS6bYb1
wSbfCZdTdJ6m2OFgzRBSU5UcSqIunj+UQgY27j12zBDGQRhGohyjB1hMBJxFoCY8
nQz0G3OUdrP15CUNEfGE57EOaWsN8WsOL5xtICgmlRF1U4bqpNq/h/GZiCN8hrw0
kP2zEkLB0voV+/kTpfk4aFmEHZx+9OSlByHNMLRhz2k3MPQXw8m5x1oenfmFpEMz
2b7cMAmTD3pEVreXM/JFoyp0xw9ZpKj5Emb7QTewxyh3A8BXtPCqj29sX7Ic+3Rj
taTPE0W/c1G+lkI37R0kZOGYHYvG5Ivf1oCe+OI6ROMa3MpBQuB8orSMkh+/KaaJ
aE7Yx73NJYG8eYobH36MIo0Rv27pJmE8w+lh7LBOB5PIBi02Bka83ncv3myCHApi
SNUbHcAP2KCZOmh7p72euay+HkyyFTrd2f/P4IUmtzfkqnM6JegUJmlvNycHBq/o
saH4J91EupgyUFo6zuSE8yvGK9CaabTj0EJbRHsC+GWwU6jKl93FHVV7Ezs/NUXg
c/mQdfhy4ln11Zy4KSUDcg0tSIgD7e3JEmGPclzrj8EEJe4qPKS9gTeyTpVkYbVK
GYc6U0efwvv4QUuqWMYsPUploXhp26vEyIfd48JDM1O8timiqOyEGrVidPF81vCs
LvwgVFFGGRZwA2TrhLeXW7fdq0wqQu08A1m5XwSoboqnKgvDR7w3Ig7ykpeyrbiC
JggJSOqUUTLpMsyPCmxUtvHfhJ7t69nX2e/iPc3btCFwz9AHkkVlOPEyHTKlmzSy
Foa+41yrplLWJG1E/X1t6IHCcJ4HcD+LQQWyNE+I2bwy7bRP4aTds5oFC0742fcw
adWGj2gWDlVajqttSnbETeFaeRy9Nll/UOPE7qZ3YeVCKna36IkYu0gUsI98gzN4
sJAsRmUfoz/FQk6vzZGqy+kn7gNOvazCjWDTLB6PyZBJphXzdxIJdktObTaRW/h7
FN890o6OrzL+hq6WNugYqa9tfYmmLKzhBnpMq3sa07oAdrX0A8bbCKS704iIn+OP
3WLzwqWUWjzJCr3p05usPGoZKNBmvotDkEUwnnkvQwe0wTEpcpxUUugsqFZuLDFW
V4GsyLBlkRfu3rjzTVsLE1bxZXe/4fLvY/YcfH03peaN8hO0dhyuXPlGfqFqxucN
8wu8XB+RuQfXmPLp+oKXl/Gh5NyMia8I2RtsutUJPFBKsMjxKwhXvdMBnv6KtX+D
4XjlDTB5xXnhdk0wAeISZ3z3xZm22yjDZLEMv4tujrpqegxFQcLgnYD1QISWVwMi
SrtxI8ycsA9XSwyfKHkvF7AAL6Q3my/gHqbjBadOpo7TAeJGthJ0+p653EQVIAxL
fujjLUnkSIsRNLczoWyYP0MrJJ4iHdNqm7a1cnt+Ej4oWCzPNk7EpdwoUrcbPokD
JM7Ix9+sOolJfMrZf4XRWftX8umeLxRoG6PN8Mbbtef0l2+kJ3IsXQYnJ/lbv6IA
N3hiYgBcblIlHurrQ94qrtnucYvK2opl/SzppTMTr1tFrB4HEIB1FyP1ipvvZNS+
E5Q4myRc2KCB0I6LmDwMt5OUhcpfocclGKWdtFpFYAE3UIRE2DQxbFdQZPLo5CAi
TPY5DIw1l2MMaLcuDDuNmAAiKoVBpTQ1O7jUvWHod903dOQ+NLek8N/FmePkJltC
MXwLNrCg62ATrKFuGT3dC1baYgqLOgvvBbV3aX5dKFbY6+KTQq7m0aw1oEotKwFt
bSDvXgwcrSrTPWgu/tKddT2ygpPeNQ8x+gjt+UIeduGvyoEK0Ayz2KgMDvuWaItN
siddLC7NN7J1o4QcV52CpPJctSPonwXQZYIcwD3Md2OMAf8lQrrbscveaailAuh4
I0Q7+ch42dM/LgYz4VTLuim4GstEZymhn2AyGFrWV3gUZPlrBA0uI1dzluns3RB4
u3YzkuEKJCEe9esk9u+xESJ7jvXI5zyEy+wrJZLqxf+duBbBPRZKWwdGYpbJ+dXQ
sGqauBOcz7SLpEksRg/iqoEHZ+lTZdrgva8JqOTdilOO+F8/LUmlcq5vhMT3GKYe
uBTMTPRMkX0O0b3fDFY9F31x4IPFRPQhT8Kt+sSP5oZP+9K+adBkeVdXtumcCiGA
tY4L6sSqiU+ld1Bxcl/dpUkUe8AxLntW0+BXTB+V2FqP8Vx6Adbo196j1e979T6g
dURpPVqN4tETmv/aNsDPoj/hRI9aDTi4Q3t16cpbFYpGdQ2sy3x3qcqO4U6Z93XH
9R/gG01Jsa+RgFGUlvJQJqXsomfCaNSlk/WqTRtiP8CKAIoftlfOuUHbuJKnTTYB
sf47Kan7skAM5dcZC3bhnvbFDEQw4Yvm7HZlcV0/CMQkCS0ovvYUjIWthdx9iUqH
2uphEdPZwx0pKL2vxbUPV/BRPHOd9EGYW6cF6kFUCzRTdJjSjhBpYoK3yXkOGrW/
2YtSuhi3AHozIEcr22trInyaWkrClFEPVXEFVPwFuGm96efinYp02Sz+UNNSCKAP
00WhX1m+4EzHoBn8I3onGRYkFo1nYt/Dwgnf5aY0v9OjfD37jWlJMdibY5xHIGnj
EFLECGC3VPaZ5zcaG/KMsmOvRy7euNdWmyqrSZgQE/2LUkLxamHx/kNBUOyhcB+O
vyhns4O1WNr5yLPIvCX/UKwYgTkAwvVvr8aXCLWsVRj/YD/evONsIWym9NuTko0g
AKQ2pZDAJVDpCUSrejD2lD3JQf2A++9YeGjfn7AuxNKiH9Fbpq/xPrptl18XbHG9
N+ezqRxnfVq47vBY4FaD0iahELWDWtWujYjR43uSsxIg4FT9gzsBRaY+Ai19fZgE
C1e2fcjuyrMV9n3FGMH+JL6UQ65X2hLbj0hB7mx/dUhKQWrUFSdhZRYslMOCJR14
J29BwSFGqJvqvb5m37IfYmsHy9PtBN4vTsMmpdp+Nj6j+Yfw+nI5JBo6UG/MuAuZ
YmX58y8LtAW4PMTDeMgGtTZE8YYR+S3UPt5XNdvAuvOxC5d7/zTRyFiD9385BdR8
AKw1Mr0uCJTxw6Qu7kwpjRwhQmCmJXrmB0HHiQJ66M5tzZjqocm+m+FHwzGYr6wq
WPxTHHa5Hmn8zJ6hRGYMXMrf/pUSUdA4yHIYttGKPSB3nDI+Zf+QvLy5171AXWOa
UVT11sTD3Pc3M2quHoC108EqPTJ69MGfoIUJ+DMLQ3tdPBG5Qi5PA7zvRxZc+FiS
3fmwCWYiiVkn9u5dK7J1creNEii069r0pWWfMedE2KyP428Lc9/6FAdRmVk8JkBe
S2LhVtr/Q/CH7pD6s5a2dnR6aoqbTUeX0/o4sseWQ1GFAnOuWuTiaHv+JXREEFSy
Ql+85TdbUt/rztwqQIuIQwFQw35irlib+MSBALsBONV/iK8Cn0Lwdzybb0+3HGRe
gTgKC3wpkerz7vXVTJOpCJ2b2pYbrESYmQvP9xAe3/gTpF7lDOZD47k4mfgevxir
BlX7F1EBtRRUbg0YnXDq2FK0mvExw75me/Hqc27nR+SOLr+vMxk6kATFYE0esK+1
j3R5oReKw+X57Pw2ixobCFdh+IlSc01SDZaG0B7N/Byiufbw3DB0gZof5WxWRpxt
/s2U4eylZ484CYUPGKaIlVLenqwTdIXfFJGavmuq8hqYy2T7Ba0C9+ew4Xazc4yL
f8uFwyf3bBFp80HnYnIvpR4FZU2jZeuEL9sHtdwG628IFgmVvx4TLSW6k0pf+goW
yYHEaz5r9rsg4tf0J5WazV4Ih22pkgOgrJ7m/XtmCqMZ5wB4OtcpulQqJZ4K0MAz
Wu8Pim4N6Jv/nRadUZ4eLUlHUTxz4FIunqCVBVLz7fy+JQi5kQ7nfd1fJPRHngiX
YjEP2DU83k2iqL5y4rra4fxdhGvqvtzsz9GBu71DMhOZ0aJZwFXtXz7x2VMTfjeW
URoFdWxWwzbU0Rh0jfUaoHiuxQNxmvH3ZgR9Vvxr/dBi60y78ZeGjRN1sufLMzw0
vO/aziRsQXWgqTkH4Yl5gf+Eq8s4oUGdTrimbqjxQuLS4qRRnWETfEcl4tLxkxr/
GmlJcxrwDBaXN39cQP/0cCOaQN8+ecGi+gJaM1QRrVpCsHPHVBQtvAv7g2ZXoj/j
a+xLBJ/417hzHgebop1xdQs4BluHq9XqDvGbns7zb3b3O7SRlRkR1Mm6OIEkE54k
TnkTlrMVOqJvGF456jR41XLLInd0nUFbQDZUBoNM0HVjeHHw57w2Z+srPh9W/m9A
osAwSeqCvS6FoSzSz/Y9V8Ubj6m6Jk/hhktobyqOSuNlfsllc/PpVNTa2HGuQJXe
NKVIKgHcxlGXMrJD5H4k8LQ3V/2BcFJNp/MBZDtYOBOQzUbh9GuJkHM5I/zAxpny
0kpw54uZiReglQ2JHBqhGBscyMat844aVB/VxOCZBy5NfNIyd3IMcF8AFRHU8FbC
s1cYjTEYwc9Ml7GrdjzPjpiKwW0Jo/7IPbzc95G+pW7OSm9xhSxvKDE+IaMrSnPe
W2yn6/tM9M3NsRFhDvr8nJ9kW8aViz5KEX129ArLBxxmpZimcd64Un4I759qZoc3
r1MDvbXZp2WHe0zQLL+lJyLarX6x/Q5WQRrMKCYIor1SzDbZFCOo8laH47Z8hTXB
yD8PfLaNPlfKVtUeJGYb2bFqC1KJsmnFpy5R2FaPRIkT7hIq+EPXriVGC1vKE+b9
+kyexIDOyVl/Fqs7USBiGFTpPMTzGVVZKPBGSS60jUMpg8V0LcHFN2GU4qkTmy8m
Swl5enOOMxxWq++ofZsQJQUgogfr8fi20iktvdNYJbCLVi8+65PSDNItKUzDcLJc
7q9Ay0HuQDhPceWErXxKO2q73TPBlyI+peOLMGEe890GzGCnIKt5iiX3CUmJ6JhG
inthfzZbILe6PAK9DyFpq0zfSuTDqwF/WYJQ+HsTmp4Hm3AoE8PxNTNt9CiiKlp5
jx8cZW+5ejruCAJ4deAinoNbtStJoBbkX+RJ8LJvsnI0ayLEwyKwR7bCIXU9rwKR
VcqkfyCzrA4W3eSAVdDDRES38dOeQs7qSur6P7qU1VdXCwqVeS8sYlwOV8xm3D16
AcCoXO7pISIk4fj8aOTKcewMzrmE0nqnkloAN/AYKvbydaiLdMESZ3JQKlxXtruh
0OSiGiYF3MLFUEnll77a5NJWfSm6niuaMuNfTFkUZJvLkUFJflaKm7Uk2PRYT5L9
DENuQGD7bhZ9OJrt2r5+OAtBygZyhaYQjqPTR7gQsQCns8ALFblv3f2uQiWLkNaE
a8xV/ABBcw7RnkjGgdiRBinZ3kk7wBIcph00VhKCt8AJffp0WS9e0N4P56sAn4uu
jH7tHicAMcaHSpe81WjCaayfXECs9rLFFdpcROf555sjI43sTHvhvL8ACmWgKQGJ
sl/HLYIMdAr6s+BSPOXf1G1IWPMf+rxPzp7X6TDVydMrWzUlNJnjOuVM3rd4VvZL
Z1PE6ZjCrD2/SIdfPT5qWn2YfYuswmvar/NHvR+cZbEgi1IUOs9HKG8Jafw4R1bn
E7Tzy3KFvckn5hJfd6XqOms6LdJx0ZX4BmcL0WdviC7BsFgdhDVfcFuiV1DmNkjq
eRCLqTXEbfUD7XEn5BGyOIjAYBJVW5reMl+hm7vHuI7pwrdop4AjVkPbQ0jQZnxs
p3uxtJzelizfcU7VX+dMl91rg86uIgv/r0tqc2w0tjP4jvuNYAZ7dtUWqF3X6ClQ
z3sbruQCvdT4xaz3YoNUVlHweKXioim6/bfRX+YV4S8yA6NwsPfniUSWmjHcnHLM
oSTjALfMccmxqC0MPe/CJTqCnNTZflkzVFWDL2SFXwO+tqB/qeTfYKLFuAmvo73q
9hIM5Ap28mjAvCcKsVCWERQ2/cVURACY0/lUbZek173GDghk45cVpBkZbfnFSXmC
qyMIqeSC9Dkns4aOE4hQx01/+Kt3mAR696n8Smp6fgmVRxTxrSE29xPucpEOW2KC
oP9Ed0QjCZ8gmUTPr5tn5ze/au+VRVlMKVPEY5rNzy6po9Yem8PqWkxsTRBFv8nY
ZyiJMHKFaG50zztq99KOQaqWga5ukjOeFvegCiRV+n9As+DDmEsa1s+m+NmOM0jS
j42R8PieklLYS/SSyuJy0MKSSP3G9iXsiIiU86crkpnOilQQYsS9JSSW7odhy9jE
hq/d1sqT6/O/IxIrgHCURQ02xoj3ITDXLpt3tPMU69DbSmOEBfHsVnLdcAjoeKDO
wU9NctkmJR3Nyw9IPNw15JDKvAY3LToNQn4QsS8Lbk0eVq5txiFcj1wUmoiO96T0
I+SgyXtI31nRxO3O+qkUYVZWAQ/z3r6BpIepQGBG9GxtySz+dBAbiM7Ggpp14WPu
CV4wO5d0ulJbDIOZ7ZQbKKaOuXT5vaCO1DZP14hVWj4DUAx0M5FxkenM0I6+A/qX
Ln3FEBJyb13v5PEx2wWR6yh8IYscrXx9Kw2drYB8UGthkQWCRUbaGEuwRCqkG4Pn
lE2bPlb/+k1Pk1ox6NEwUV1pDfxdtIjR+a1dWLljRo7slgAv7KAk8N/KArB0Iwpe
yWpnGSwuJlcUxNj7oTCvJfVNu9fx26LhhI+/YaJtQ1u+bxjW2amUlCAtbtUaBN2P
a0hj4fdGYg6AnJDykBe5PJ5umE77YkcmhGLEyBNpOf8bbfbeSuyO9Wc2CcvK3AtZ
+fi95lfc3fDX3gTBg92K+A2dMHsXtThoKyJ2/iGvNaRuXoYvE2Py3IbF+WE6WxQh
a0PrKMKPepXQKrMHBNB2plJae3YkRlmXYGK+4xpWRdA62uylCiwUULzM7s5dXWDI
mNM60+Ww6q4dlybWUzvq0MoK7LNxJkMKFcW1/xUoVk1FkEqu+015fOi4Q6Uh/Sw0
8hbmzSm/sPmtHheD9D042U9I1tRcJmm0TtfhfXtSlxoCMA0T4xfkOFJE92Jr+50C
1iAzjf3LX9gJ3nGLuyv0I2zpYGqvwj0+ZA0eiFRD7pwdyQCYUd/hpnFKbkIIg+8h
qFi73s27POEwc3pM4fsSjiC17Owjqkfj2OHWfeWj1awDX/RCKjnw0C3ERqS6jnPn
mnKOqgdbAzWhnXIS9+F7OepZQKkTd5bfW7WrHdnTnswJeSIKoKz48QI8uaHN/uAb
DvCKyonaKP3tZRAQFuXJ2zGp9Sw8/3Ee8vVBvOE4O4y+c2XPfPJ7m410tPGD0Moj
hYN2zhkv3msDGVsmbfVyT5OdN0eM2EV2axfNP4LF0RmWL0ooztoeGqi/5bvYUn5e
S2h10Xsc1grl7l/ozUP1xnLF0P95cVUDmNjQWB3A4heQbGWw6y+ZzeZ/m7GRGW/n
AdUgDpeCHHr8XmMSoE/EALTfpDfOz3ctS8TcU+r1yNadX4mY+eejIv8y3euGTJUW
bgnkWuw0dUY5bCfvoa8dRcwx57q1V0miV3qZnQVfpNMJxHuX5xxsAsk4qa3qSMpG
EiBuIf4OKhOkLZ8NadlPRJmMcJoIfOKtQnqaDAVvIV4Qx6rHwfL6KLHd3EQLwogC
hLfZquA0G9b6K0uYdKyYQ5QH8SmtiufbZGJWqGnoVBbWx5Pwt7Tc6RPJ7JFqXkau
qrX1uOvolEO51UZfYFp4NNNPYQtrNn2IezTNVXj8UkDTgcZv9ZA+GqomDB++edf1
o53jYB56eliH1hyDzkSJ1y8KbKPg4Kj9X+TJwKFxoo5KKYsXqODrEc2x24RCQmb2
cwZS1048DPzBCLA9+FJEibgsj54hnWfYGSneDlVGTtFjrvbYhTLh5rqjZx/rk4Av
Cbt1P0EBtLoVos2TLaTNWBUd1ORXSdOEGPADnr80OuD0J38YA20ibp8GAOoQjQ2T
kdwrdaiOGrOTraxZflBGkWJcuVW3M3c+wyFt+yPWtQATX1UKy68BlmfWs18zSlvj
faQjLYRhPDZ9ja02e436yi2Kh7TO9xqiwr3Eng5W1gJ9EG6LeIyjLV+Ggf9doJ2G
SZq+mZSmFy7NmU4E4kw+utZIUwhNopFhHRiwNRK4xVeTD1ZIM2L0fbS5nr0I/O0c
tIIdwMjCM1KqPR7hwCHW6l9JWh/HpdfHj/P6NEsggERj81ozaNNlL+sbLO5xya1J
DvQGjf3kZyd7758iDNPAhU7rYS00HUE39y1FkPFSpmJ5g9k6TfABJpSvEomoOvi4
E/B+PgBpLkOtLAFcnAssraicqoitO5hsv44eIP0/D5HeYnWKdjH9pth9SLi9WN2t
sFyhBlNomkWaaIxZ8I1SWOzh5Bu7tBSyqRqyw44AwTrEEw2ic1Ux091tQNRgbh7E
UkGduhHDMM+qpNqNDq0JfKEj7ZR7VPRF6x6KCz0L5d1MCa7JTSPTPeBs+3RXXf+4
3NkPHBkzTXiwSUz45NOekyYNOB45fXgOnwXe5S5Hrm0F3xIoFwUmO79Aq+hzsQdI
gqE38JKwp7mgcLR3eb/3qH78g5X/sZlnBfH+Ohbh80tQvspCZM4hELg3NU89dfku
jcoRiQZFZAFWjWMHO01w0yKyM9nqfSuPkHFGuASsYKp6suoyfTOT+8LgH2KqLoWu
3Nee1CSoKO5QaFhu1I5/VqVxpa3sOBmqZb2ooebwLQQwiFWUZNHE1TEEGZA0r6Ua
IEKnyd4CQ+xh9O9aetR6AYtewMtRQunDYRm7rWsR1BjX5WVjVONfnHTmGMhv5kON
JbA2GQuWxYixHO0b9Ga+DvGtPIL0SHDz7QQZC5AWPRK3lw+tvCgM0jK9zG5WMm/n
8/90Cf75eeGmAWrMV2MlpduOP8cgWrL26q56VRj3NvdlygoYC6m3Ja0Lo6nJ61gH
NW+Z9clNRUqjU5SWqVj6YSMxPRKpNUVXRZJvmC75EhPt9eZdFUJnrzYWS9ydJzBp
oKORDDtYutzX4liDRWW9+Ht3x56pqu7dB7APTyJgQTLya5LumqHH8wiVy35HG1pZ
foiTai8IkRXCZ7KlEdYxVGQG/k/521Q+ZTPo6ff+zOi2haKgXkf8h9SI8F+xazHh
RgXzcMIB0dYyEcB/GBGZ7NdzbcLg84ZZ30zE6IVNaPeUlWjeAF17jw/U/cISSUAe
AB4L8kQ7TXPv4WeqFna9bvKvZXr0jX9E7r+kF8v/X+gd9n4Vyy/623U16viM4hMy
KtiS97XcaiCSJh19ZqwaO8Nm0qH9mJSY/4uadKXX8viwWaqdCaxIFs0OGNQXgJyY
U0tvX04uK/G1/s3gCYplUJYggfSubdJ8ZFaP4Y3JdxHBUdfQHUmqswFqQA8SgDRz
TdN3BJhruIXsDNoz+RbZsbiqsJRtadKAejfhFFV3bcRowFYlfSJ+yOCYW6QbPB/9
RPecWbcmElO07k93rWG39E8er/qQWbLPY/SDYLOqNc/fe3FpjQLAvNqtsSiGGo91
eOpnVvkiDW84hbYoCINTpQ+gTZ1GA6fIZ5zO73W1NShW+dyF6y9uHk+7c30+mnNg
X0NQh9ixvuLAKVtYZlaLU/9HzK9+/2VUHyiXmdM7n1zGKym2+AybywJq6iY8VOJy
WFSANAeBS7wp+3OMTdtcJkgZLnandKOepc5SCTnGzpMzCuR/HrQ6EhpMkNnOqqOU
KXTIbOvfO65Ics1nhYBisPx6RvhrC9wpmKffncCyvL6ej/tni+B0tlhVOLySsdaC
huukfI0AStS1Mdlgt8X2xrz1l7U3UZzT+4R/ZMTLeqpglFVxMdo5QrICLIQZ2CnY
CEdUMJN5pDiMKYdq08hdr3QV1Ku6OJkR9qxm2J0vhLQ=
`pragma protect end_protected
