// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bJa8mxQd+ycluhkKpm/v78WC0rni3YoYw7wr7WTplfcs8ThIxvSYkR5SS0ViavLa
DWN3ona0PzO2NFqrtFvUtmQKsSq+WpXfKVHf87GMt6f95uT0fNSsClAKVCPoMKaq
Sw/uOBlQcnXBmQWVkmmTM66BK6v0YRGJhpxhkxNK+5Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16912)
nZBZFn7QjdAOUcZA8mCuLbIgO3tJ7XanBh4EQvJ15W41AvLy0170slI6MO+TEr8n
uNMfYYeRdvysFR7gPaCLc7QJs0lP/+sUeKy9aD4g8TE8iAqEiF9zlGWpz3PP8pWL
EG75QR0N+y/xhnf1CyaSNYYdhcb1XQwUNDHfn+gQNjLS11rvu6q3CINaLYLAr5ps
+onGAWDq1aGh4MgqcY2dX7NZzm5E9f25IsLe1mSH6T7jbSogeOFvro1pR6C9MX/u
4c3LAtLxZoAzPpZpyVNNlrvbFS/SuhH66DdmZ9vlfX/LwLpUs+flnZriDPEo1QjC
ok12fDE05n2i/lPV7loPLrzgXs8lJ0EIeFAGDvS+mSctjPhklxe6lYo5g9x6DtyN
XCUkGQhqZDiQwaxjCRYndPQDfOqeuqzK9F3QpgC8HP/Psbujyd0Zg3vtCpq5d+Z1
8uAByS2ss5etvdxOrS4wCNu0Rhw8UzzUSTXnH6B7M/scLKlE9lZikVIOUegTALYK
VTkqQi6pRL9cGUlfTuEjjUZ4zpa37nStx7UB77stvAACWdFpBBbcBpr5dX7e9F+V
vibPJ+955CEVLf4soeFSjSoT3FFWzteC6X1Q22f0CCrKIbFw89eM8TB6T89brXAK
WsaoLu849/USgYS/5vdz5lZfzk/Rw8M7nMFel+lL3myQkH76XuXZ5MhWKiPekUE5
FF/tcSYU0Jhwe42rqP13Y5CPK6LtRg4EJX2ssBRfyWA8/Qu1GGekWKMRgImecc5M
K7Wn/3OuxVMPTdEvbJtv50wTqBPFcDxGjNYIRmtxQNrDNGhTQw+xTzoYfwP4E+2a
LCdrAeQWhuDNW+HCq449OiF0SP/JQzQxvN1xtsmPLWK5+i98MRMsW1wUU9z85jqv
NfGbvQz0YUFd41MgkTr3KK9q33zn4tZoKv2VPxm6DWuxIfsjHjccN7wDw4xnpf8x
FpVtLP25Ezb/BV7TVAGhYqGRpbQFTVCCWgXR3eyeWUbeOurl6Q9yNhEKlnwglgvM
2u/1sEbDfseZZ/VM4kCwpW4r4VYCPK6+1nyyKMuxbrjlu9gyR3kuJcILqbYBZJoE
samouAS38P/IeswnYOC4re6MCxljfC9DpOR/oZUsI+i7rLU1xhj62NE2HRSQRWUh
vIEd9E9u3jNcycEcUakDn3sTvXKEBhallToTqDs0yngDbpkD0LV+fjL7uy079UiP
eBOsbFXM+9tMaCERylixaZxAJZs8C1n+88S2pUA6MIQRw6Ox5i1tf5PByptmsxBy
UGC0K/s8zkeykc6+0nbmBwA0U+3c9yFA9TxhvxBn+Zu+fuEwGZK/puz0yT5Outfe
Mi1XHy+uHNLqckw8BjZVxVN0LUYxvKLCZ0wqK698GIxlGXn8p6QLKWlb8/sFGTGd
CIMl0eEplErkJohGKaZRkrMS1ZX58vwMx48dnWxHC6qXqXBliV5gWGjnxGAuEQii
pSuG215k8ROTJwogSfjJC5BFeqB+oH21QKMY6HpwMZp9+4fgRXr/OuLwnKLHdPXa
qUeiWtQe8kPrnyzfSk89eCJBfz6gwMFxrvdJkpPrqJsR8RWFu2QKXNlZP/Bk0rpY
2YR9cE7lohB/7FVTMnN6tD4qtSCQBeH/0IJhbQJX2L8LOVYcCdSUZL9MgRTvwXYN
S3ryIT0KL19HcDyShO4tLAgdZhlMzo0gRmPE3uBD6xHavhNVCNdQX/MxKV6CkhOZ
mcQTvxs82DSugFbu4I+m/gREh/xsz7gXHUaFEdL5Y1Qr1nAjeTtigfzW8xr2fe65
HKCPheO+GDygFQ/vuX6aAZDyknAy4qyUVk6IlbdgL8KmHUa+qRGx70WHl5CQCVtk
clV3Ncrdb+tqhk+NjSzQj0kbiF+nMChRfeCipjia/6RFu+vhYSHznkbzo5RbAsY0
4bEEeqVvVYMPp5QCXyLlNVEVrj77SWGS/rjPR71EoYgeelioyOBl+J9FL3R7YH0X
NsQQARrzuAP5zfTDWdfqqcSnIGEQXSI9Wa7j76/VV+2ggtFe9XN/GOpH7Ur+aXzz
ThrUxGwUvPJoMe3Z/e2dUc/l0c5QttMieA5BYnpcl6jP6MmJUG7N8qCXc65/FsCz
LYV1vKLhELhnHRwit94CvO/3CBAa2L9XG5FkOieOMT4R39EmtLJE0l/n75ebaZy4
cAloZ9YVOlCqBWYLmX+PZsHIZve3LvINuhueO5ogZ8aUJzTUFcOEJLWUnWVKPXap
9HvpOOd8grC1IRg5a2v2EEo3nNrMpl1fLP3TSLHSUCZYa0/lYaUTPyVVPBint+YJ
jnsMSbUW3cnDxt0hRPrDjiRXdC3iSoAnyGPfsSFDR6ZdCzY/BsaHCyjaul9PDciB
V1GjjAkCKG10NZ7pmrAEVB7MQZYNynJkv8BFf6Nn1aJN7VUIMBqjbZWxF0cAqAWV
14SHkMX9xWavb60WDM2MXvAVCbsXjN0iZq0wQ7tFtYbMQZ2L4KNQMZwq3XpWx3uO
mAwcyjq0/ONzTrCTW3VEGjIMXiz/Io/jDuGzf1cO4YqFhFYocR6LZ/JIjrJOJ014
TINN+m9/yVCD0r1IhYctNZ0sKX5GTytZYhYY6Ggcfew+3RCseMeVmgkARKS5ilAS
3alJjaJzQ9SY2ACjHfL76GQL+rbne0E8pgqE7tH5BZS449LcVdbx376hKUUo8xBN
wmqAEb2d5nirLe8fS+ZG/ySczPpGPVqL54udLZ91L27Df7J0+Ky9G2N72XJRTI0V
oGVCrjxgIdxCCRNWHNKHg+wRKYdb15x2InpS/vqdH0mX2USQ5PvCndD88/vefbxk
XBvwZF/wirASpK+KRVaBvwpxZ7aD6Zbpus6TKwOYaer0js0y4vmw0enCPU3p9oi8
wYE36pv43nSBKPKyp1kaz/O3yMdnnmLNwzxQ5X005WrRA83WFpniq9VsSNIB7Auv
1C2/PbblBCP6aUL3465M7eadw2HNQasLZRQil4LO4VMwawZPNan0dD3DmRD6+GiL
2CQ1xbRBkRqXm1/8JdJCPYOslqcw+DG+51yWAyD+GNshab7IIY7Opp7Ud8IHNFUR
99wCYngZS1hMV1LOzBIwtD8+1PoqqcZY9zBU9Pd+bsHdC0GKht7tbm+lXGKcETpn
mTLn3BIfmjggck+UPaThxHcsjBE6NOMagh1byUo6UIYPVh3OicEeeApJ1BMCxe8o
V935ESjgYW8NMDipqt9t7buS/M2pFo5PMaOj7SlEq9UVtmhPtLficRyOBZltyN6M
CSTFKjD2KLcVoQ4o6pnlNuX2TJ+APL+T+TQPExa7LoG1keivPgj7pn+65rWohBF/
s9MORECUsGRP1F3l1lRpLvxNtmrJ7PoUcygovul1TKkRUP5PQdcKL1ibYJbS+Vgo
ZnGqEWRassL9vd9h/QCz8kRZpuumarkfNgpP23Yo8wUkdCMfaNaAoMfdZdoZeMeD
zOr7WgbBONRuX1DTJ/EwfyAbFbA5PYGrAgvqvqpDjq2oCC5tnfDiR5WweXZKp8de
W+Ktd2PcTaEeFcEckv8+/uaB3mzqqRsP04M0c2XCLx/6rsmVKM+FkoCHGc/VO88A
LpklnGxgRcZKRC5+JonPebsT2n9cUMGGXrjDHrTVHz0keflgVDkGz8xzISA+H6PZ
WkCmwuSH4eqIrjDML9/vQKCRBX1qgTLfQ6lQHLBXyLssx4GcjzvT/3QxWDUJ9eh6
1SkDIgfB1Be2NDG76DA/ho7qtYzT7kXjSRR5PevIPQ5hctpLGm0Bq0omZE+7Mpfl
ZVjDyzCzkm9OuTwckowXukpLUmPhcG5i1MpdtDve+mb1wylHvFFyD78Yy6Wy0RUC
egFPxavoTw7tghedxG7oWv67jii17hnNROrpE7YI2i7R1eGxQY3IepEX1Zq/PbYX
YwKv+TwXZ/Tln0vTkYeerHNtoKDGkCkN0CBFwfxgDauDaVt0Y/Fn/VZ/V0XtTAdI
PhD00irYjsdlRL2i3+U/s+M2/DALpt1mCVBeS8ilZUjYO5tHcpTkmlmZZp3XltDD
KzsNvGa+Ukaf3pBwn/Lpe+jhh8tZNtuiltYObGcTl68D/XbANx6msvnT+YzUz7Po
orAL3ZLEsQ7sZF0t1vpCECtjeM1KDfg0xkZeCxxY/o5+D4mNFQNOzLTfBHOt58Gx
EI5Q/VWuMaHv8z6BXOuyOpMKnvvdKKZqDngcOe463C8f77XEckuvuYnWmWnllbRH
QGUZAZ/Cyelpp065uYIa/DCfj/7RveSxJwUDLe4bk3Hf0thOJuppTFcoGn1T7Bet
zsm0k4dR/9AZlo8cosc/pGxO9nIOC/o37OsxAaEuPADlqR4czZnR4IFoLLT3JUrD
lJiOrDmimnfQrl7c8M6QCkpzkTN6fjlWkPsivfjwWTTz1rtJsu9taei8eZFhPFna
7EB4PTZjvndyEQSFbCb8DZ55af4TovJ0DnsFS+KgUXo1aCGD5XQEMbbMO0Opv/xv
NWF892Ix/5j/zUzOk526wsQDV6kSJhmsptf9lDyXEBq7AFqd2eCL3xKCMCsKjqz1
b760AWpQWQRLCWVQb5HhTeCHjtI2Op5HPIdQUXOSCr6U5AEqKRz8WZ9Zttn1sWXb
RfPxtiF9wQARrvsw3H4ZIqtpbU5JZsJuBTdjJdHjLM4L2SufvdKe5mtjpIxQNw1F
IGOeoGr95fYF6b/DTC990WUDNYOZ/I1N2WOPDYRdGVGNZJAEtpu8yWqAAskGXuZV
xDzbXbJfHbwjEvFISS+5HP6lQUD6gX0IkJUQHI8cVrvtyHvQ5ZzyAf1wZw239BBr
FGzjo2doDF2Sv2n1arlLPmWo/Xv74aCJyeXZHhJ4flXNbLc6ZM+onHqarw2RzW8f
YN4cgsvjYsuLHP5rPssKAesmAEx4GRVag+T5jHiv/O3DtEKDLm2TpT2NprbInr/J
s8xWgtJxagjP4PuY8m/pL/2W8tGaZiBEd0gRiLzCfK5sQWStaZqxudnhmqNQPHLp
SaeFal+Ns1qCJAIo02V8xf6/3d0ArVbGRPRz4le/8kdoajiEEGCDBu4CI+cVc/BQ
gVg76f10XylyHo+bKBZR3SIdfrIUKkYn6jajpQd5HRn66zq3NXdxUlZ8mKHQ9SQm
rlyYS2mPGhwyo09z8PypoySmcSHCr/qtlXpMcdxSxUQccjyuofaUgf28AVPWciJd
Zyue0nmT4FCtl9tstx3+CwvZmROs6lO43mO6WS/xTqMbkSepytIg9GbJvQ+951Ay
go3Rt9ANzF6oDRr3SffWaIaRGmnbnNdZGVHqOJ8oCS+Ogn7sqA12Glq1qV2rX5en
vh5TUTO2KWd73Zs2HTfPvOiQF551gCUjflgFBaFxIazKgOcP9Z7K0TiQ9dYhAqPO
vgVvavAhW/spK5iQPTUEwtUsTVy+nRlEvabXjeK9Xw8Kw44hY6ZM6iqvTd0QCSBx
R7ncd2R+/8oED+CUiYgRTUFzWvYLc1hvOtIUN70gTJLiwL9skDQmoi2J3w+l3mK1
ii7PSyz6eGzaIjMFuxGotKqdHIm8U4hxEpQ+X2V2FBMIcZd2Cej7knN1CoKfczoz
D/vYuclyv6I7gDl3bmwIwGohoD8aycqUhTuzT4PpdtK0yW68YlVhVOXGEjomUib9
QkLwIXNp+VOu0y88WSrfOcOm03x28z5WY4CvDNxZ9ctLQd+I2SxBNHO7B4IBbdQA
1ok2uV9CYRRpFpj/Len0ZiHC1jQAXn18gSt5zuPWd2uPDHHTN5Kg5sv3gNLCPdUB
Sca67MB/yae6jOVpYXlMToh57RLv8qC5QQX9mqukq3BP08VD76IUDEsmXxF2aVf8
4+s6Go8WLFK3Ox9Mr0CavtBfwqBiTa1WKStrhw/396KhKXjmLkABhOT0oXEk8+/Q
5YQIBdUfEBgPOxe88mhnmT1M+uJsXDQFSGcKoyVJfLp7J4Ek4LdC8slImc6BwoXI
4cViJ0SRjf53c/HDeI0b6N+UhXpSA62lmdftDTYsXfpAKmFYlCxHa6ZoLtlTL1+q
deHnxnN9/XWO5O1iWJSsSycZddlgij1QqP0Y+pi0jhwjIy2znl1sFr3hQPu9CXS1
RvOuEDj8rlI02BYlrPeySIjl9gr0MwWV3CFaf0u4uFP8juLmFqL/E627xcjGKk0Y
U54FRNOFKig4vSHOfMCATuoaGINmA5N3OVkG8fId0tr8ndYwd/KcBeU7CnDt6z3i
3O68l/NjdyCyfcuB+a24vDfER0+cHfVKP6ux8gfNSE16xIqCOst6S0vubdwF0Kin
LKrOC2pDZXIb5PXDLNB2mRMv+jHeot0aoE474HR0/oPW3J140BPpIoGMrwNnznvb
EFP+EOzScrTrd7XIc74v0coBkYwjh/SGqtlVnhDdw5J97fqU6yzSXNH2tVTbZKBA
Tj51RT4L1+ZQSmFFt5sTAaGyPp0nBN24QeOGzc5t7ScVmWPrROKp7eh2tRuf8WGM
gMJSyvnr2XNovx5Gplw3jOeHsxIffJcZctTHEQ/bEw2P9gzoNWpgfKqL8qTzm3dR
a9F7L9//4l9tCbAmDpyX1sdEIYGHZf843GIuHgGw5z2vpS/e8oVJTBZrLuGaPNbX
glLKn5dZ3HmiXhIa9t/OiKw6/FKeK/ojNXUE6fXjHwZXafOYU+QUn+SsTL8q5Ijb
yas4E27ooHCTCkCSmaKqTTie4jRSp+1jHa/DNruVU1varwUYcHeJLoy2uLqpIrtw
w82EBSs5gXKfYOKC3ng8DSoBp3ZJV4j/KDPW2vY8Nb8UW54eeNmX1txTiELfaOuG
heVe1MRGQyG/0ZNTBhp8JoD8vR++u2OACVKpqTzStvPpgYFv2ervnrGZmfOp+o+/
glFg/S+bYUVHCFTWwlmIocGgj2pddsd+fD66FKzctx7W85v5VDXivqcWKWIWzt0R
ObWGYo0kHyZy+mnKRhA4v95NmHol2j4si3vIhgl9YY3+wXQTZWytvW2F8ztB0691
0dZMbw4N7Sm0fko80e37amEP6TP7WZlxzQwx9IxlhUDhVd3vyHR2uPxlkr+yoD6b
Tbptx9IGNJTnghY4xNhdK5Uv8aMilbr0+CngQ6XNWqoNBLUEcSeiLzlZe296fghw
CzxZn1Ef5sezXg5OvwR7mW22zeQ3f6ak9PZ16rHQER02ozKrwrrwyDxwDEZInmnV
MMav7CV9dWvgEagZJIiekcpj2t/AGBeXl1IhZSHimSOvEDXYiJofoxxuib7aD+Mp
UPBGoiqfNMo2AXKCgCz+fKECTJTNXQgo7PALr6bjok7vpVsU095pro8FGh1EKRZf
rKenNub8KReI+lNZ2bYhrCb/1vBofiFde/ujsIKcyYr5igvB9WbAGqvKRQmWn8GZ
d7hIoFxg8B07+1cVIOVGp1dhfMJHo3+1/085iO8H4bbG7cyiV4GHEvzKbKfyLwWl
qazTCvMJedIqXAc0WiV4SRGQxAjGmdI7ePNzsyVYr3scTpqHwheAeJZ+/PKgOGkJ
aOW7YuPt2kMZtGbmCev/udXgSr0K9cC7MBlchd8HKTTgMLsNuRnOc37x3oYWUM6b
SiRI2lPGT12aOkS+svTgdzetEhO0ABzFsbljRmbtmGDbHOpK5ciikOPnLBsKYAGQ
Dk88d6TbFsWsdE42VYpzL9eALRUabk0AHv7O75hPrsp082Fofo2Z66b/5s8eGt9+
i4SEL3vIBIX5s0eZIS7UIhtLWcouamAdg2B2VrnGijd9uFHTRIkZgbKM+HYwxdp2
iu+xGjiAYeRRtqysoNIeOKW29jbJX/l+ShJH4wuuTmjtznz0RCwpj6pXzE4UWY4U
4oEwCR+8W9KBqg60Uz6VgyedwF7SOcwvsz5sCUwryMVatqCKppK0JQGfYkQ4E23Q
zV5zqnjQ4ru9DM7a1b0Iso5aRAnDHaoQlSVprONtDiQclgomJLqaGFN94JnFYFBi
mQQMhIzuyZnRM1NqzCGcMBfAsaSpfAJtyFDioN4ETQs5AhrmyRAuFFifFql3FjsL
QEo3Km1mni9hTE2rAxH+AtS4Etd2/e53pH7mV/zPvXlBIukgE6CoOXwsQulWWsoT
EUFh+pibHWBvLgopCWl2fve5EDebfwf35XGIU7V3zo84Y6H2ZMPpDi2BKSiOeUET
inEK0MCQWyZQ+BI92WR8pKXDgjLngu0Lst/D4TdcPQZ1n5vX5C/nD1+cQX3+48bf
CLoIjfEzeC3nZWCeaTmrtvzOAIetaQmyXHfYNrQyYdM2yITTm8kX748I8Ts2OQrA
NxUHox4KQLfj/zBF1k7DQWTVrpQfS6TwEe8JpHPabU0Uyd9RrO4shhsUGMCzwnu4
EWeMeWVKivRXnJZFX5yJorNKWS4rOQJjOyNMDiUQBj8Ut9QJEcFdEZeHIoQ3n/XB
dTG84aKGBcWcDF3X0OjXfM6IZwRgXyKtr3Pu2AdwbGIlX1OZw85MGu8t6Lo1wOXg
dYUUJonDXq1aiuugvdKfRqE60XA0iAo5QJvDk8cEyS8MdgzdKkTciVyqFs85IfVS
2YnVkMN1pyjgMBSS0YDj2AOB2lQM+gS1+c/jqEWS89XPjzf38UO7Fq1zdUFCyhDH
T+/O1UqrgcMkpU0IZJO89uEM+8WFO02nCLVoyJ6LU+5deDPv2IdcbmmT5mFqNJ+q
Rt3du0w14sfZBz+m8wWgoX+W+QwYtFJ491TWjqXxyTOpiwtwGURIbsCufJLhDLvl
8c76kc0Np6CCJwGTjANk4Pm4G/DhMatdKpsg8CEk9r1vOerzNsPKBKAuzqm7ltOg
6+tU8zXQKv6WFXlMLr2vd8OcTlV7Cvo0+NoWqjkDAKMU6B54NA2eTtTcgsRvlPI6
3BGrPrKXPCcTROKoty/+qBCBh+ftLMMD7ao/eWjXruOBqS9zO6AOw7TV8xLLK3aN
EfDTv0C/5w3StQh4QUixAElJv+CiHUNbSiUwOPfRraO39e4KoOofV1rDT0ZE/9m5
WHb1wRj2W2FZa07Vi3GzGMH3KO0B2pvtQz6Vpee32otDyVSZ7c0F3O1CMgvijHEc
PyNp8gwPUEsgXeS9xCs5BYEuymDjh+1HhmnLfN+EL3CRYcoVe5IYQjbhoh0piJGM
0fIWseexwAj6TMTiVznnix+uRDFj2Z3N+EUtDYqUDanrOjxz3xDJa1/yikBYFhIx
i/ZiiSepKtne63yFvVWVtnD94XY0iDdTSU6msHQpPE+tYgyontXitfURX6cHlhO/
ejUu+7M0M0yu/4AR/+uT/OEx7gB95rHPUnjTOhcju+QfEYDSrTCsJ9C10lBwfvn+
X8BRzEIt2L6S8AZJzD+JI+y0fQYNWn3zBcLzG3z4zW/y01ngohW/IBGszU3ABLNm
Bvt5JWAuaNi2Z3jd9hWxOPQl8Nt+q0fM5QPtpdDYRK3Nc7WrkSY7qEERHk5HwBNO
JjGEdqQ2T4gZY37xg77iGLdhoYr9OXTcTsRT+hAO1SWYP/tQH2zzVGPsnUHtR2nH
yY8XF2KmN4o6NsypcokauxhjgflOQiJG8Fy1xJhatCajE3QyAs2GaYJHLWam7DLh
yLaGE2VqvRmrmZ9BNw9TqWuhGsK9uiUHleOk6OMi3NwO2srPdBFW0HZdh/JiX7c1
ss4gNed/xj5MNdWUAQzVM6FIqqEsTPDGGj67Myx8QeJhTBbkkZDKvjWdJ/gcZlt0
amZh8m2OlX3H3TbZzwuUSa2qZg+Y3tJCRYQcmFln+zqf0nsDNIYmUhv2DtZ5OvD0
MMXOeoWRXTUmNrlox1MjNRl8dno8/R4DBsigVHceCvI29a+9j5PkfnOTyTeSuTGO
ObLhQyWGDsDpS9VVjXO35kSYDc36M5G0eKdbaUaULTUmxdwVmUjlAXGZ0IA16Dxv
vO3+O4h69YJQVylhO5VARzoUDghtMr6k8Wuw+uynJ8CLcbsL5AfhNoLbQG8kmlF5
odbNQaZchicwmHW7D0Hcx2CucyKr5TAFCDXXVr9UNefHXhIKWjcUHb/gfLHY670I
JJV++LbVTPXEANN8fSw9qUZFBjAHd4P/FDrUq2CSnqTwz7jiX3RpdQzFcp5pmqB3
LZWpS0f/jFz2kq/XBA+OBvqpMBPkTzk/jm8GO7YOE44NJQ8e6+cjv0Z1g5gxxpBh
sqa9QBldW6aDyA7cOLbgbHJEV3uUAhtF7Zk9T5WFwre6EY28PwlnAr/b1YS4m2f7
7JKcQx8xMyoy42veAm6xvvbfBAdX3ZJvdOVzEjdK9839bI7Z2RdENJUj7hbexsJK
vzqLznXWaiCW0GOJvc81kPxPzz4UeGZUp/UgpXyjYUQ9QOiHKAFavDKxqaaXdHGG
UEG5x16jEd3ssbCBLdKDPQufydqs3vn5QRqLAxGvWgZ0WTi53EGArr3Kous9Xm5Z
oKAIPxo2A5E79d5E0PMiTW95wpQ7bwRZ7+9BLsWlwYKJnKVHBIMP/UkKwZfV+0qn
yMyH+dG9l29DJQALanh7EfFnvNYlYgjt18Gm4gjmwetOqBM6ebnuZ9mdb184dcgy
wZNYifNrkL4zymRbCp+y2bKEtGJeNu/MNFFtkmZlMQfMzWconbdfLURO+So9LqFl
JHLe0reC++VPeGYL45TFevKovaRpbhJ3Yo1bdwu8ZjD/LT3MU7ilb936JacYraU+
F5kfLsTQYqMtnDTxR5elx3mO+0Xf3GKs8Or5S+ZdTozgfLJa1Zb4DiOZVub6dDB6
/7iQQigALQZMh7XRezTRmk8GSvKaGM4GTBboCmmRpmPN2Hb9K84HETNOiyEB4+Ua
T72RRM9lgGaDHo8fK3rtnPlzcWyj8vJHDxQ1Y1rwCuw6eW6OSErSG9Wi9KQl8xXv
Nld1j0UzoPv3mKVpl+sxY5cXvdyWmoRL+KzVlvc6dS8pd7Ev2EKrJOq+jUpZlgki
wJK6QHaKfN4L6Ihawjhec8xq9t4jbjHkFKhstSHp24ZXf32r28Sakgow1m7dXEMm
IV739uYoRyogAf0LjiMp/Tdqj/osPvqK9tYVuOT9CkJCmcn862MoJy/F/qC4MGbj
2H8NO4x0fLxNzoIhgQqz7z6O1mvMNdznZihO0yLBxV/jgVWgPkKbSyiWY+bIQBRf
DI1oQ+K3gZtWiwR06VceYEBPqnOTF+9+p2IPicfrCeqCpee4q4S/aVKAtopxFpry
F/IHeL8fPuOBgkAFVlouhvEEr84FjhKdCUDdeK2/bHTJ85SnsSlmWJAPZAB0CI4H
rTTVpn4xLeE0V58lde/ezoXqDut+dCv5Oru7TCnYHSlgKFm/ncEpl4qVtmoqiXad
kTGZPxmcant6OW5JvapIYtEuVytnjdnca0AfPj9LUd1312wZTribphit2KG7fzgI
Rvql58sKrGqlIHyuBRDYFEPMspWOfKndnSn4AZw5MBMnJAzam7XngIisqsjfNxXt
mQ1LqfzpvOAg0wo1GQglx7T0w+4z8PkVgjlyqxcbplpHQWyO019oU8omv0teJMXu
4BtkMeTu0Vebd4t/3YaWGM7w04unSBsZSUiltXy6JlDVT/GFf4mzIgKJY5jzTdr9
xXEwO6HVq9G2S4S+FWvnL3JBoSWk6bquKZQ0ReuD+zpjStAS+hpWv6fMj+P+xQjM
fpYQQFyPxnFJD2wQJruO6Qvi7xeNbuQlsOUvBOFXgZt2i/Zi3UNHqmmuS2NS70sF
Totb1tNOBZmpb0059xw8py6itZ+sNg1CRoQvHfZh4bMJbNVzDmJ2vT6CAhiATFUJ
/A2wusZLfAYuf8ud3iOp4owd9Uzu/XIzB8xgHieaqURFLR4xwSzmxn7ptCSOT7+F
pGLKIlr7nGb+VGx8WSp7XF/UeLAdJqRL++wK1HDEGUI2Q8oDrg9Fwo33rQnnsAv7
TSeTOfxSwvx2HHFc1l8YifmiwmyL4ZGUh75OMct07gR0pBN69W8kmpRvmenCdWH9
SPCLsJkIghrm0x4aDXOlXNufUYLIehCkqTEbZEVyshXcQyVkb6pF4wpFRhfUN/8p
pZGUU9nCp3cXaKfvR/SL9KiuaL2/VSp2LM+qHtPjiUJm9UXYlaxHg33qJuY1Xndw
XT5xV+glsnn2g4NSvdF9tWWEq/RvBiS+CqmJ2ODZYwKZpdMfSpRVKHkHjmL/uaI2
nQUg8SBBU4px+kDozVNDIf1xiMRDu61uMUfp31wehTydY0n5Zm0D/iX0qbljsNV7
lVEFofcLTg2MBAW5z5bhFDdz57RwnlYTGmEYpyWb6Y+woeD28nc2clQ7eB1qvJ7p
X6aKpk2pgHwha8JnbY1W7gN5UcoCqdqz0ckWkhi/oIOjgFBN+1w7plrW5gmnCZrk
vDQF1XyMNPjHceNeaAVBH2DG8GRQu1nsSXrlx0OQo6rhK3a2xGzBWsE1Kcd9fSgA
D1prn/21OALwyo8wLfARtB7T9SR3gP04A3QSAC6nSL7w6H9Jj/l8vJSkG4ichGL6
ZqwOT8c5ahNuiXAI+WtaS7O3Ork0mGDvOZnKD0FjT60EWaBpX87NPZmVOkQKhmz8
Lf3sYcw37cElW7WztjaTK8hv7rE/52IGUcXDuTcqCouUiOVvBDOh9wgVMPZbde0k
Myh64WLbFPeSTnxNPrz4FPwbTwtLozGOylr8XJIybLwXzTFtYBesX7Q2Q4Uo5PrK
rbGQr8sXyacKeCT1hkdP5+SDmUakjEAnlGfTIYFs2Ia/SEdirOEccswWHLVbe+w8
8HChlFxGsyEODBRRusozBJy1ZlH1Tg4IEkY92qlbUYhEorTxvaxjOi5ITOjj1Iiu
GuVdlhzipAKv4L/xvuyPE3qPWuIT/T6AdYZEIMKsdSTsbZs2weewAhEJCYfHvBal
egbwQ4Wk9zgjFMg33Vd9m64LjLu3RuzqYl5UEmaqQCBntcNsekyS2YuYRl2XbanS
sXg7/MGx3TfsO1JhKOWOJdWwG8NiImL2V2NLvNj3ck9VOljAc2RVYr+dWp9+AEZ1
uWhsztTLrr86qgYToxyutJwIxJT5Yb2TBUYAaQzdADv+QlVn6+pJc7GB5T32nhXJ
rG+GWUB9WvpJY3MYHeZoaZytke32SSeqU9prkQOunqh9feQCfBDKhVitVwhvMVw3
X2V9OiTTe0fD/49/JRF4kZ3S2LvwE2iBTgjRxkk2FtVEgUAR62kGORIX4+RHKDLk
fvJqlgHmJZwYVQJ0oXNO7JQxAXZMMvZJn6+JZbOd06yPupys61RHQ2c4F4PQ/gBF
oVDPNSXZzsZ1RPohenaFD90t//Y87ujMeS5kyyaS53a+n02rDtxnOy8aVNY91Rns
qdRzJJMAk0Xdf5wlmGF+pG4ekL08taWcqUlIPu85NSbPFq9WieMMSABZwfTEEo94
cR614Dn0x71hUJHTOSz4OJgbOQnrUlZf8WklU7qdplF6lBaIg/1mzfNQcxS0XxZ9
IdVFnVTWsZ1aw/wCQu8pay26Y4+zVoh9j7LKceXfZQ7Z6rj6+NbsNt4gbqZwJMpc
4wtHTEXSJVzqEx1rGTa3OmGw4/RHDuXVlr8/3oiA5GuSrvuzgF5rwPlnLs0rJfw4
h46H5m2y2mzqqufmqKNPyo0gnRsSy3A/Gv9lgy3sG8r2YE06TCvXYMGeW//zXmMf
N4U3vUHEd2F8iSRc0gwDo+DfgJEGtciCPiIoCRJHeW1SL9PUMmwLkf6b4vkTKGje
lvUloLZ940Y0x8K5zQE2+bfplsLjRuBSbb2nCeaBvFHSn8ky7WZljiP9UaphrUsK
MmJP93yVKxbTjUVTWT2wvDWAowJ8HahSKIw7Ss5kCwbZnyHP+Kx3ysHETTyO0k0F
0RI9MyrbB21b9jUzdMk1VBEzJFNWMyUMnq+ppL46Gc8FczMfVtu+jm0lGJUkURml
hMyeT0rNcv86nqbzczkoQLTT582VUdRyAv6d7aJD2Uo/XAAJM/Rt4MkNYZ40Ual4
Hp7/MvlzEX8opDtaQTP/f2T3Owq8kJyi80Nz+tyCAoBHBF011TRJ6nSG7+W2WC5P
ICoWxlZpuziSurEuSXYcWwGQAEi1vr+RKHdOVXb1Vn/YH8JJc9cPbHkFk1CdYjfw
ZM6wFq1MNUVBM6NEy6KPLCcxX+j2G/10JAfpmzBVQGS+iP419uEs5MduSYZyoO/H
L8/JpNTw5Wmq26u6YVyPvqCynNchtRCp8916VdqhUG2ENaFcP2e3xP1b4E/ktep9
Mm0fcVS/iEYnhgI/Z3XRje7IIRuT4AUuctZ3lKRWaiwEzb3ZONPErM2xDkxJ3UiG
0SA1NMCyvlD5HO6cEDi7WgBoQCz81m1lfgQKdo265w4DZtV464+S79sMgHzSBRMy
xVSFUwbTsfBWJrZKPMOrl9bouhpO+A/3FOumc/qVsu1FcEYCvrf8ZRRKvmOG+GDm
cPJK2HoJBtP9ruhRq9ZR2kepUt/WEK5VNUQH901Qb3DO/dlgB9tmeY2yRgSlATNk
8KRqE/2h3xkMsv3Q6gkw9FCLNVfc2YUc5TW/XKNAwnn9w/mf12zM1gKNTq6Inrb9
6L+4l0nFkBVCkPMzHwQIf+8sfObokNbIj+qhQfcxnVEbljifQyqWFHVyt+QcZkyR
ll5wWMaE9G8LIhzdpJ7Wcx9Te4Ty4kNnpB0Ycf6BUsTHbIPWJ9QfnfiVYoCFPDJp
0npaxNze1lgi5jDDG8a0aVm8LHsjqVz9+gtb2ps2IeXIi33tzfVeIQLb4rKa7CMc
QlHMtOeKmgF/VOCXsUVB9Elr+/UbSIN5Ij8XwqbA2kvk/6H2JOORxTbs9BvC2hta
u6RHt15nAu0OBD9ZYBksA6yq8c7isQII3h+4Lm3SfRjSgbtBbq0daXltRE4rQREP
HIDc4cvnr7V4fbcY7A9s5jB2CAyA0lUS/Nbq9fkuP5Gm17NfvIOIFJ0SfEAsSDZL
BVZ7GRfORoRt07aldiOimZscqU39pCHZFAr58tVve+lu0qxA5MmH6WlD0880q9EY
SZ65iVIIcx7MD8DBJbFpZseVMvXwVP9gfW7to7hNi5vcbTV+qdUo7xzfQ1OJ7YIu
gjnLtEeioFm2fz2MaS0WpH74MXtKI3DhRIkGD7BZQwPoItoDorPklyzcApEBRDsz
ZTIArYMvwfWQ+FJ/mLhpSX0cHB7nU7oPtkmsmYmQoWwTWwZ4ZWK0DxqNaj3j44IG
ZWYWK4Hg9FFFJiIjkVbgBrWwb1ANKZcPpwkheL0fbgNepM9L/Scn7AdsXDQyEzZh
89z/9fvA4zjXpR81pHsqzLwXVqlTVz3GnQZ1WHmvPQVlQSMZFti5TZkVCjnsynD2
mSWiliDXVsMrBQCTKbxH5wgM6H7Oe2WPnJdTNb4w0Z2gG675rxAzMW1nLq9Gt6oN
mLbhwVnQYQtlz05gMjAoYNVu0mzj5o/BPZvMUvZ5MabRCnEPSOXwb1iJ4BvAaRNk
fZ8lP5X7VsCZyv6wn76XoesuNkJeJC6RILwwOfW5IqqaCGwRTWH5CKI4yo1CAKqm
J4k08WZVJ3fwF2pssTR4r0MpyrlN+pzi8t8TnVWoRMLhIWBHsXwsq3E+EslQu2c3
oGDtRwugtOxmWPJ8LyBDXTeAk7K0ln89defN7TdDLCihqqeOij+Xqpjc0hsimZch
/zhmpzJRa/uA6p+y+JAZ3KsGZncgaac0rcytjXz+aQgUAozkFDoqIxVsD+iuvqkg
gQ8qs8adkzlbmHTMY89iq3FG10udP0C83V7QS4zPU7LgYasC1cKtBsl7Rc5eAcH1
vKZzl04vmyvNi0JuXmEJ0Vm5GErf40AGfJzbzfKH6LhLEpWtwGPOIQoIjYnVY8P5
qHNvKiX6qllvP4JeW1KsU0v2z6j5KlFswJXrbDtoeEmtjK8GxXYgEGGA8O8Z71Md
WyoiRLBhWsQFYC6wPoe7i1HOuKubNH9+fagiBcoxZBLVqEIZBPU7ABISiBgSbwH8
QcgvqgTRxAnqSG6Qy7WuhiDG0+/SaSlccH0R80QCZ/Ze+wmJw3bq9DPEY5cwoAT4
EQmuuf5V4VH8hjwdBgtjwbQEfjsf59skfLAQ9iO0VUop6yaK7e+elqF38VPNqcqH
0bypMyjiJ/IbH2e9SHi4F3l/3UWF7xEFjPiXMZZlGXZ6M3Rm7VgNtHlEuX9hjQvF
u+hGkdw7G7ucBSOmr5v/f+wEFpVX73z/a15b0OOPu+dBMPi+EmZtoVET6IYzENKM
dopb+sWwsXxFlyr0DQuzEurcBJmKyWYIsVkpgh6wuifJDG5zw7ChjtUorWm0j4dh
tOXbS2LHxn/yKQnlLnUXZuN257hlD/WAaYdlgH3a3bq0a8JtAp9XHABJiHvS/HR8
ZHeScm3yg0rfioSHw1xiRljIr5Bi5viUcVHHGoB5SKQE5IvUFKjSpXK4Wmfi7sWj
f5X36K9VlBAZanKiyvowsjKQbgarW8Z7+zUSKQWRaUuGaavwqFVwTcRfSxOY//ja
mSfS3uL28dtWJHTADJAfegk/gHiPLC9NECM1G9kwwLRflvLrZeYtNvk4pYk9APxJ
WmSTAwqWa4YOBr2CtknfBImkyMqttieGRzT52KOGYS+WqymWcO0NhDKArSgLubKC
a/5oyg+3qAxGp63WPL6e4QBe4BIGpRs5AtyG9oywO41sqA8D9lYhp1btjXek/IVO
cYfBUkdm0lXqzwF29AgQPx5ntvt/zRVeSPINq8zibJzhqis+KfR5/xVqbgGUAcbx
t59p4rqVU+/LO4H43uh2GpS1VH+i/KgQiIk6sKPt6JPuEWRFl5Mq6O88GPag5gpX
qtpucd8biH+IC/gKxHh3xQluNJm+LXSdic94so8uIhDrfgapotPCQDco55WqWfZB
zeiYEELx3j/amYiLpV35kKUezCvEepH48d6za7CjDUH5CPvrnhFtpXvmd/podRPx
qJww240ho5STMjHEpI635fWLPbPgC1RMcnzSYYIBEvW7o/3CV3/mDZ2agZxMp29N
FrC8Mr2NBLXL3OFG5BJjF5oM2PEyFAHjlgNMBbZ7L1I8BHLHhi7ZkzAaxUW37jQY
zp42E2lc9nF4ixaMTd8Uut68Nmr1dXCA7YWwXpdSuB+ud8LYdixtmAq3Q3NBT6Jf
fw+cUd2F5SlMpB/xVKpNTpkqBSJHqL1doesFJkC0AfB3li34p7jhp00AG/clSYkG
1X6nz/IvXscFIzniKKh1sgYu8VH6jSp9taipoRghXT09GzmVFjR4NDyckw714s9V
3LBsRaSNSjgAzl5DD7b67oVckfXz49D+oSUNtBES+2DRR0GRXvYGLxc6+dmHJPRZ
M6aYfY38hAtVQONs/j/Kp0TvutOECkOkhZfkPdmR934FpVk0gJqDrGKlXJug21I8
w5wa9taqeuh7YNdJG9+GG+nnkMimS8PenqePyF0musZe08U8mTsUZTfkXmj3dRcN
m0dw4wyD5JPnmrONELll7a+nJYoONeavRFIOcoK2BJyA9yKhN9/HD71kLZl+jbWD
7qtOSmzZjSIZ25kAprjzPeFHqfGNjHfr8Aum0t4UK66zGTJuOleCRbvX8u44zYuB
ATgMQsWWATCn1HYByaFstLFabM4glROetYN6IF5ynqDfTDFk0AqSzMOAZ2r0M7qZ
uLrVXuSrqluRPOMTejYtt9AQLFlVC+BfGLgKoj2l3Hkd+9MJhA9bS9p7aCZ6jFKT
lumNrNcl+kKDSci8IEtwkutHqmINCtXZCUefPcgBSk+o9URM05iFvej2u8WG2n4E
oHNhD9j1st7QeAF+Jr6RFMvUOvEYR+TfsDFp3vOEJUmm10six/rPrdia0XJmOzfn
1uigwQzQDRqB1WB0Z31DmaUBn1mRpngJKJWOM95mR1yH/a61cy1jeUY3a6gBplXF
pzNnG1qDnsBj8W+HNMsHJOj3HoBrAMB4ZscmEb6UP3qGFtIZB7byFPkHfacYa0KN
W97d6+MAeToS3cOlS3p1JsPc4ECZoOe6eZ/J3k9rJ6/uY7qi86TawZOQD2qg+SqY
XD1VUaHo3N26frWvzJuHAkkjAqr2MJEEhNyq9X1hwGbVxE6hO1GuPeR0Y4OY21Ut
zaeDPDm6kcyTwfxd0/f5DRSJOy4BtAjugnFVDfwdA9ZcRP/qUixQ4Tj7iQsIPhu3
We3sWXoAnxUzjm4SLeLUfFZjT1bCqT6+V87F+qKmD8kyYjtYNVy9o9s64QRw7uMS
o5TwAUxMpfR/jYVh3yyulLCoGyny++BWR38XsN00xfsRSW3tW97dI8gNBfcXVnGK
F+eIsRCI/058JxQihHjTTGav4P+GQoab9RyOx7Z4hmA6Qd2rcXlBCZJcuWGGE3Xp
tTe34dqV6raaK24d6xmtTmNlgGC5jnXRESwS7hqj8QqQXPr3K1xDZ5E08+w8Kpmw
0QcxH37IP9yKga7CnN/xshZoOljpEsylBnWT4KOLjPnq/Wzd2EbxrykGg6ATNI6o
GWg/2qmVUF8XoUenSra7EJdoT/EQxfH/BzvEIUrWV1vIeKfSDXdGzXkqTr2sVlwa
yIYkxPr7ec5epkJXtNg2sEwJ/hOjFOxRiT6btTcPgUymXUh4ff8OlQ8fWMedPcSZ
hyRgxiNybBT/8Piipe4Fk5ZZLi9R0RX5vOVLBTKHS+0FDQ2pszn6ivho9yEw0wSR
tIFVEuS3S0S9O7JkmrgRdSgkdHHrjzne6ahEgW0J/iyB18rNe1W0UjEHMmj+sMng
hPtnCPV7Ms0ljksLTjP4YjqH8BohDypP5K4udLI1EVsmdmqTG2JMIPVGlGpT0iFt
cQ+VizFwtlGTsCndKLnY3zEdyaIOFO0l97zLnJBTxgBYsB2pb9+tuiw5tfjr8xa9
sT/jjjx2Z/Vhl0DzIScYXRZFmMvZv5TbapQWA+9IKACWNbhJ7A47ZmNhQ3n69YkU
oyPIa0Bw1pvV/s27EvGLjeaZ663VbBHKHePQX+TWMptCZOxfraYJqiuc2+eddyV+
b9ym8LkpBqwAJQgHT+heWnxZUIfRGVmpiLsWOZGVy3+jrGAUr1685CcmchebeTfJ
T3YYqLZeZW9EQV9lSk4jVm4ahDocJZgd8JGr8X1/A42GkjgZSlL67iVQ+OamP5ef
P6pbebW2JGrDi39EcKgmUWgvoMoogcZrLWVz0w94h5+NWRDH5nEPM3t5P7K5GtcQ
7qvc3YvaDbNdwAfsENd4Zz2dw/WILCYNLox91VxbXUE9hJF8O2PL8T+RRYK7LXok
S1aTGRNimOCSBMlIvPCIGuJETW8gOjsBwcAG+kOAGBD/1yLjrFJDV5cIpylPrF4Y
SPhcjyOurE9shz4G/eDsXuIDiyw8tZ/eKPOnTrhHkAA49aoli0yOhfe0O8jyfijj
JbddTXz+me2lYNVM6/OLujB/4iytT9TH2ycdhh1AWeTB2dsK//M/oBOgcYSGZKmQ
alM/YYj7GbIKW8R/xhXQQUzaXwtgfZyNMMQu2e0JWvgD01vHv/RmhQOnwYZwgRDX
dN2Wtu5AghccCz3+FgQ/auW7tggqdRRPh66Xs3BbOQUFdgUs09p8SxeisSmf3eKl
wcKZMyPp5Cmb4XJ4PIV6CoLhwcNb6qzhFM53y9yb19r9y4MQOs9HuinUDKW7Yc8i
EJWbQtHIT5EL5XRs8BC6CbOUISHBKxQN9ywg5a52cakzNz4Tm2GL/YVzmZx+K63y
PJxnQ79z8PRevJkNoqyc/kPLJjCWJ8KvL2fiUqvh+4929728fqLkcvgCEZx/Kw6w
nhEeq/XSBuS7C3xJ2/uGcdsm4zVyaSUBD26cLAatEfHwB8ISWq6HffKXFiaSJG1o
emg6ID/zHkyeeE7P5GplrJSCihhbbfBDL6OdeYFJKCuVQilzwTQ5VAQrQgYAtwJ6
Enwojxk/0D/mY9buP6bqVv+Nj01FcnA8P03AqzEUVIshq5nczSvbRHS7jxtj/4Q8
e+9mb1MaJczSsMSG/qNR/8XVD1GXYHe3n1fxT3qyjIAVYSq0XEBawTZWDGKiY2MT
GJGCrg3vyGtrv0B6hTo2s6DQm/kKxNBFHRLlReEmC2b5BcX+reFFEjetvhhiSgq7
sBI6/2JTGeSPLUJtgWrh/bpHFZiXPGSolac0pF+8IUrjmOCpE4JS2Hq6CuJ9WQCZ
N2XpC7gtE58xuid/HsjIjqbCDFEafaQyuOrI1p1WGafzw88p9g5Cm1JKtBjim0AT
cUH4wj5wAzqYF3No1yTo2IbSaAO/wm220cmEyAXbXP0elgy2GgtPPuLbytL3MBg+
Xg2c9vndbXHvqVNeMeYzP6jg9u1oqpruCei6kuFebWFfkbev/Dl+QEgCosYNUsU2
vQva38PhGy0irwiiefDL+c+qsMbL7+jsyuspuZoCAG7e4uu5j4HmpejPzrfYBeUx
faSosHStuSrIzjbOTHqpE8D1VrZHwydTAD6R32gOJjefnSFguF8XdSVsMgZxhroU
3r7+KFEqn746MUxGvEWocN7l4GNq99fWxUeTO0G/hfCIW9aHiR/AfdRzj+GT5a+p
y8uQyFtgOzfe16OynG/l5TWC3ezRa4S7CjO85tzW0FBL1NKey4ODhfFsrzEORo4g
icbh4vi/it2F7DSbQRtAtt+3iLlTvogtLIDLbjJb2gjG8wkxIJ64rLHmDcMQrjiF
n5yWVkD3eJz/pU0zvKEYQz/pATtSqWEWLDLhbYOf7iK1KxbO/kJdVqsYZZo+T6gT
EHPGqyTUYa5mxuHluLg/BYpW0EfnblfGP1xBvs/bMvKrQDdbtcCKQgNCgwp+llXf
ZxSpes6+a8k3LJQFQMrpcveIs+MU3B08uedmJwiwoIPGBHi0Pputc8VjzEyKJ876
2df5yKzJVT6i3vpZ2OImcutFg9DtOLH9IpC7Rb8IAgEUNx4B7RbTqZxP8DSJFE9g
5BrhSL5YPxsYHBex610xoumWVjMvyiM80+b16ptkpoEnbnVwIrq+xI8AUQs5ZyBp
YzosbXHVEAb6ku5awhKDWyL6W2+uwUc4BEq1fjIHGX3bj1h84D9UQ3sBXmD10iwH
cQR0mI2N5ODGKEQVnKSK7Fc4ihaPkm/F4K/qNTav/RF2sKCcRFcrWw/HGJGxi6We
jiYFeyWjW0ayeoEK8L6M3htxOPlaF5mk31Qlfr2Qx2MJCwJEXLSk0Lfc59FvmWRB
WMmFesodn7jnvnVksRxcX3rXYBYmnHkmF66ZrlAySmsuJnlAsNcjFiWTG2LWOGLu
Je8UE81mXw/n2hM/8x7rjhfdsbmir7X/yaXLdnuzFpcuBRYD0WGqNZdLVtpX4wqn
sFxtDnlmhcsZVQFozKj5p0FVuKS3lNskrAAAfo3ymH5Gif6CYhTvd+twFdC80IQ7
4pKbno5zTxfyoQEqo8bpbLNhL2icinkZQ7PcJr7pAEwhd1cjFrKNLl2Yzv8r/Z1v
bJA8VoRSf1jbttjAvhjOoWc9tVdhjCw7zaM4gsM3RqsYs00x9aKoKFkU+Gxjuh+m
/SNK1R8+dKZkPxQFiffnCtjUZ45rg6jIqJz3dDCNy6vDwvu/0X8sJ8MB8uQCG1Wp
+G7/R46j563n5Iogj2fuFHwXA171doXc9gXt4n4Cvb9F+K8bnHU4EEYGjGZXdwVo
bQ0zQ4D5kmeFolaZegFtejSzjqwTRK9Vk4tRM7fxD4n4OtTeDnt90H59HyKa30hd
SnYsXTeVPlgspP1TG34/rYGuVNr2tgR3DhfkEnsrE02zKuM+kjtKqoMimzbnAXPd
X6aGQod3EKfNsBtjwqeawFOY6YXu9xXZOVyL6UR42XeAAUFbYfbhuFzd2kJZ43/V
ptYD9kTaxWIwS69kgirCaKsUWN6iXNISDcLHXGfHqPw/VQ2603kpWkBA0LyZZG9t
4nGUp9tp0O35JY5f4SBR9y8iEhnOkZnU7E0IIaave0shDubkN+uauLsf7O+HFDwr
j1yM6R6JJDRqhNjxDbjZySGL+ujzsu0gnDA30VBj/mvh6HTBly68XQLpKnvtJP1H
e9jsAUb1D3f7ihzVZulzwZU7I+vQNC8maQVFkMZW/t36wdUZ0pT4pGjO+XoNdoig
9KU463DaqfOntFgCY0topUFuqtOpN/7O6Wwi3vCrwqsv73cvngYN2XwXv5iTwrd1
VMRlCzRcOwPZk0hHtNzw5TJh0R+Kfw8g7qsLBuAcTdMObi0G6lOp3jF4RsVHFPNE
g6jWQdEvkapQ35c+wzOMIhB0kOse+rcDDwZ/EK6cP7+78yAxXej1s7xfYUE3feT0
ejk0YAJqiuQiDhY1iDV9PfXXn8YWlBr/y8URvzz/h4qtiem2FHkOWIG6SVFM6e7V
52KHjTY43WIzmgpRIyy3nQsgGsRTX4nAxl+QBMVwoKxRSu6ouRyE05TNT0/fvH9c
2U1y0EJdq9vkJU2GDjIAvE8lgcp4bXHNadWjn63QvXcAj3VfTarbQaQj5t1qVUlp
HKzztHXRMK9hnGllp5kYRKxtwDGFpmMTp59Y7QwqHTQzdiKyp+PvS8pIHGSJqeo/
MOxnZX+pnR6IOnzZn+NElnaWUtG9a3IugbKU1Hhzyfr57SiRhlZx6GkVmITfjekw
aLpFVH1GJyIuNGOBA33VVuM14JjTHOn4P2C6VkBmOtAFl+4haeHfAk96JVl8Fmyw
54/dpu8UoyPS5KAOjTDMGg==
`pragma protect end_protected
