// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
MSuUA6qb367UWNpdZXlAvd0B+FjS1jb3h9OXIEqgdzkXqLf2CA4XnHyLmyUpa/FV7rhRfgj2N0Yf
/YlIB5j660yZznUS6Qedmt70dQvCShTbKyv82Os0auS4Nl+CAwwnoZvlX8vMq9k1qwTLcw16OdYE
uvsUHzKjNcu/Wh7iaAovbqqgWOFri4THYUfl3/isLoLYw50F7bLFDzQmX4s6hScQb45ssvoavEwm
3FLqzUOEqpv+ltKMZvj6PPdNMZxumojL0FDGHSepf7bMIMitEGN9nyEUiCfzOaWFBmYOtFp16jlp
TkFZpY03KOIPlxsTpU/kaua5hD/qGqrmnjFWDg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6cfs1GTU3NAOivpLHqUaV6jWBwm6DNdZHnXZrg3BiQM7RFHTMbGILTrg5rBqWfqqIP6nEF01uG8r
sQb2DriZJGJbsjQDTtS/sfSujR8FXLSbns0kdHNrM0F0uUwcewXDZ2inMkRJxS2s3X0wpfFmpY1c
2V1Zfm946G9IZotmstkTsiwO+xiMJFmFyTlAOXCS3Nh+yUGdcK2QiALwQBZ4v1iOTAl048AIPYOF
MUCqxsIhqP/koJogPXjf6DLgl/WwYnfAu1eVc71EWFinAiicX99NVaSJwKeh+W2Az4R8KQ2XTFNS
0sTwjmJc1DnpBFpcy6F4QBLl+Rm0aM6Kks0y3SWCfInmySb9sdwhhX8G2pXf3v1XD/BJ80Mb67v2
du9ueFLn2lL9XgoiLVHluZkimWKn2nGO6mxSFcW+EzbF3K25V2R7nwqDt8bkL7mg1AEI7SJh2pNL
00Sq0Vg2vTLtXLYtiuLtsfkw4xOkZBTvqBbOOmLL7im6gCrDQV7myhah6N9EIMGsazWN9wUBt11O
7/+3CZWQrCfmV+F96v7bX9kJjySBGtj5PwhR5/936TlqJotRL07NbpGFvbgNHOmhOWH3YLoH75UF
DYbf4YD8cZVNKN3i7sMKIuIYoXSu+G+XK7aO/cWhSMS0T4omdtvHW3yl6S/v+vCW5QFWbpWStVe7
W7IOsSsAh8Y1EeBud1oO+MmofuFXBwOIm4aZBH2mQBNGTnNa9jVUaOWqH+yP1rlL/rnxb7MUpIpT
WIsdr8mTk1f+EeZDygrnm3elDKu3i8UAoKK/+hcnuT4j15IDF49gXyXHFCjanrUHhmK1r2+P5eP2
BYQWAzrK9lzDXFbJDEmrMaGXvcC9DeedIIdQ9XQGg36n+iEoQgKu2AGFAtU5sb3uN/ow7ykPSUMG
sfMp4nRkNxkPpho/+4npRnpgcx0UE5SpufbCmNHsa3S+1J+eHvvXN4eoLI6HYKELFNPixDDuta7j
ad4AUTl+pnUS/9OkrbDqRfoGQ6IoC2uNBEi82mGu4VYT5PdjYi+mqL21zABXL9kOv7lg1mvu7ahq
6pEclt32qooYKzFG7nb9tvlW21rY3h6cIfJRhH9MQ0CcWHoLVkqSR8cDL9ekteOaOUoPrE2zikZX
zee3onh1dNKPdOn6GFBB6tb49gPiyH0kVfnFvNtYL3Bk3IGbA3sUlQlb7NT/GngGWlvWNX+IILbY
91WbIIPJMEHIDah8WyXEWuBZDbI7Q2GfUcSk23mTPAOZZqmofqeIzVR58e3Qbp2aIKRvhS2isJEc
vOdjFhp3o6D8nVSF7NF0dtBtdYwKB0VP48/PaQF7iqblwDwCQPRNlim12dA3d/7/Og/locvts6jn
BPaw4QZN56eIHwf1PV//8Ko04AutRq8v7DqG4FkECJOoV5amuirdrUvC1Lpx/MG31q8MDmQFd5wM
mgaLoBrvPIwqWBC2kRPnk06/kHCmXWhXKikQZCYhVVe70XlbNrzKXgouxYc45l78x+PC7ZzCp7it
0mx5sOsDevbW4ELELiapcdR7tEfbaUErVsLOtXXQOL5TGKH/ur2LhtqTM+vd+iKH7cFMJ1TsKpQB
451Tz1ZvZJ8vQiQ01y8rOMAnqGBc8NzyuoSmmNvIRiaX+pdmqbZGe9w1TZRBLrWZ2YTr7k/eOwjG
Mo8rvPUt1vW/4AfJ2NeYcqtZDcswx8Pyfe+ahBhKuJjtVB25MIOqnEm5DZ/uvTPP4I79O6wqjB2s
CY/alwkZ4V1qALbstVT/1GQ0Qfy2x7IEQfq4NN7rxCynHMJU4ILa9k46kp8+vmOkFiMSrIjBQinY
6PV9FZoF8kM3e/7Rhmfj1RMk9cVna2uX+7KJOSOzx4P+nf6pXUFKoeYx3iNwI5jhDTXgIQfiyeOI
EIpEY6TDpd0O/vxa3Vnq/NP2lqAJ26wDecr4Pw8tJZ8qe4FoCBdJsnbfJH0LLSFHC5Bc8I1cxXs7
6UqOwUfQK84bEfCW2EpzPdBNdz39Q0AyxAAt58/q4MrBvDYrHLi/unvX2h/Cit1zvk38R0PwBu4+
cgCBUm5mW+41B/SYbTOasas7lR0WN71JoebawQ0g5ZLOM5uRgAj71oAhiAfZaylkCpLFXfLqeUlC
+yExeFSHNGA+7v/bk29CEFFPkhV8bKmU3Tzye2lo04AXsSnr6i5waKHEKnIDfTzPT9grPk1B4lKy
rVx36r9z+2UL1H3zEEVIj/w1XIkn8+TdIALRZPPdwQS6Sk3JDjGRcndcaQZ7+I/gD7aDN6ga7Ngv
V2BQZ+AhU4mH8jM+1LAlAwICP3XaaXqWIZaAPbhUkPXlgYzl+c8Y/wIlEV8IvBvGGWi6F4gqrSoh
zqa4JFCLzTDA7vC/WLXbf5D3KWZqbjnebGeBGLCyw5LXkyggVZzNecINNcsyEPI8zDnzAFnGchNo
eli9dHdQj9A0loq/qewGHApJS1fvITl4hSOhkeUtPaSRb09eEMbgaftm/Rd84Xg3/Gnhqn4TZWQu
6iVDQW+U8Cd+w1bJQtsv0Sz+hTlZk5DNKcKrYeaMvtVUGr3r6veUEiAHPRR5ZECfVfw9LpsJoksM
6uieNMJSXGDiRtceBAu2neI0QulwPeD/CHZLGJqIBBLAAc7cXRRDUf5CJRaODb48ZGxVh/VsaxG9
raRepfGSxrb17Q4zJWzRryulAzclwQ0qRQgHdlEcpNQ2d/99FbewhjKHqYBZha6MKiLVuQUeg7jd
F4EOGEskpqNByMB++aokjZzZ2hur0wGuRAeKcQSK/UjsuxE5WnhTyD0yGUUqVxPqBp5cdxbaCfOE
DrWqvsdllHyaL4lJvry014n29lQ0c+/tLeNP2o/PLYQEfC0aha+a385LKFUIfOmh0p7/mZM5ATSC
Ujra8u5yQb7n6zsvQwYmLZmJGF3nO5wSpryGpQxgTaJQ+EzHFdVSZRSZogbNK0I2IQTs74SI/3pY
Xfxe1RFWcLmRHXUI78wTd2EO9AvZF35l8s195s2HZBaA7VAGwN+P/5aNhQ8oiUikuyj0QgoL98SN
xjv3WbKkCiG+j8CaEwQRkhueUmtFDtMtf4YI4F2UD2gDmmRnX9jvP74TN+a+qamuCIhaZ5xgcWJE
sjnQHdZcagRPVERn/UnyA3bkFo/I6t+EFk1Nn+tYPfTuWCqQyPz0z4eO3pw8cJKO7MYVa7SVHayK
dMpwWEJFM5mW+CrM8i4QUSgQlty4KZDLprYqEYiqS1mszii3y2cAvf2lNFDWXxI2kDLYlGmzqe1Z
Gg23Gcjdr1jP7Ydn4cCXEC1kerjlmBxXQVLy/+SBTV9nyyStUqK9iOMU3i3jCXwnc0A2L9uFUlB2
mJE8ZjG8pZNtQlMkybiyFh1ZQCoEn8dReXi4yfdxE87kxkCpOWrpv6etfGeYpbtMzrA5LW/Q3SxK
JJevPcguBw3U7UDVm8ydB4MjRQ6l7bZMyjD0rwou5hrms6WrYPui27mhXLNW4KH1k+jKV5kCbP7S
uR0YwG6w/Beaq4CL9n4ph4m0whK81PG9hnt3c/zcjIR9qvJX4p/89XWzHAx+HZZApvEoXomW8LhT
DdD74nsdmSiF8qNq8Ns2jZniDRiXNR11oHJeePcR9D/qieCVGzxu6uNtN0oHdTQHTV8HbFrtvET6
DPEyyFBDJhjupfsF1qTvEu+RZq0rqVzKAln32mvn9/1lVgRK1p0bWQYWT7G572HhgtwMMLfWeIHH
IoZskVo8zq3hgyNVFhfKYY0RA/8U1rVhCpCZXB2zsA1immSGaM+AcPRD+HhNmnSlYC5pZOXSed1f
kV7E30vnMw90wY2KUKC6sv6nqHR/wnj+AdG9TEqMcmf0TTSwrLlwgjIj8orcU5W3gIgtxAWXxmvQ
gGzC70Il1iLRwpFe4m9tynqzX7MEcWQvTDhgV8YdqMw2jtVHhPfR5iooMlXIseDedeh1c1YUWhUv
YkK4icByCAWJNCKwpWSxOWRi+alGi3Jye70EG6OLSKMNFDg7J10jIYlVx85gQaRR+HTS3cvrmPPz
N0a7Da9VtJ+Ds95VyXwoKrujYR3+QkJUUSfSgTAtkgWF96CC1Dliz8ioJS1tK+HZQTSa0Ca1WjTc
QQvfcXSmjQwuxJLbUpG3Ij9OIQ7KOLA2H7EnYXKCbDOWoDYiIlNl2eEao8CiI7/Ulj+fHxx5g/vF
01b5cpya6DaFoIf5wCg0IxwC9Z6z8B8gb7G1sJalXPKcREuU4FETykJThbRyCKgeP1CT7i0CdqAo
yL1uhQClibc9hS+0qQmjyedeZhedBvrQ+Tkz/fJ00gtObRumEX9uJPHpTwbleL2kusr0nC8E362K
F63waEtemnDRiR9C/9iNjn8NNEetwiXS5BCI8Ajk7tWtZebGZlkwv6P+d5bTchHqTTFurkkbjcol
vStPMX/espDj0sgT1i8JVHtxmG5+YkMlMyLrUlQcwLCC+rF5mgzCLgHz2p9AXr9ToiABxjfWWL74
Kski5R0NllZH2aWMzPltT00mqvR4DvSA4l4eetzr/BmDW/WKFZcxHpsjp4xkibQTVC/wEh8NtppV
1m+5wu1MniPkhFutTcDFYYdrocb4DQgR6mmfxcd/XIOwuGfwCPq9vJiJ7W3DwiOQu101H/qfkE07
NYTEaagozApCSPRDP5yoHKvLuLyJkAIcH49F0RqOLcZxfprAjrpzzTWZHyNUR3DcQK8r8dgseLFU
vVjDaHd4Yt94RPe41vmLEqmuuoPDSCrvkkiNiFV9pRQEamDyMQ6ArPVK+gdSf2CKSHvkd+Dxun9W
+V6Vy9CWtwjjRHYYOoMBjQZQOM8Qe5ZnAyN/PX6vrHE1SwyxyP9yOXl4+qSlrfpwu9xmlewDd0Se
MNjy3p5ykwBuNdbm6+OjAT3tuKPEUQDzRkGy1N6cDXZBbOSR7DOl0tkK5awXfHfu8uIl9PDJZnI1
zq02GMiKNw+XTR7EGmbBTOcOAPmcjGWJmHONuTuFsDHuyY+ovNEAgfklfhdq43N9945IcA1uw9Ao
FxRrmrChZ1+QK/PA+jT3nXsvaWf3/kd753r5pNjEVItbf1AW7olKbOp9ZE5AsAu7xERimPZvjiii
1g+xP+vajYvJ5S3UDOCExtKtSb6Moyd4E3oC2C8eE2unfuwRfr2J5VF5pEYqrIfuN5nkpimsjCuh
LwyU4d44quVcFVqXezdSYvziuDSOQiDHKVN3Yvq/LaOGwpxv8mTcFth3X5/apJg67wM9CwlS4iK/
XT8WRqxA8JrqDrEm9oc2cMHJOTNiD4B9l4ZD0QbydxP9eibegBghN4qrSo/9vNVoV/NBRl+EXDrB
k3Q55MA5RJcObaXvlPITonOPmj8e4Xseb3dcY0JccxFSVEPcJtvUKgxU7T5+lbl3gzvfNRq7JV/F
0gvCKFmGBDZP/Qs0maZchuUOQnhic3Kl+xpyfnaLkepsre8AOuqI70wJT6qpLEeWDjHi81h75GfN
sPI7pLG8LqG2xxAtoH+y1owQsY0BWBBxZ1rBMKwCTWdtJs6rTq80OwwdT9MCeBwRgRnvmh+8CXjS
+78GUyzjVSJvmcHQyZMb6uwJJ8pPwniwIMJJIn2i0eWN7in3Tj8CBxIqQ3n2G1zothQh7zNmeo86
Z8auvkJn0Px9lzKsuEwLXpbTWoJ8tQ+f2RsVFR0NXMP0LG5wMFnBSO3US3M5zbpEtIxnADhEEyPG
QyjYCDCixKDS/cBWCrdNw4jyMPSVd7LVKstjUb2MRGbuM//wnA2q4WlFqvSRhz44zSKRMfnu0Rk9
j3BNFn6RCY9lGNogW1JPaM1+p4sEPdhwJyFA9kDRmKVkSBy0oFPS88ovfxj/MkWu+sqpPZZZwix5
1o8twlY92N8IEBQdoslWSISamAELmz1lflvknYvo1ZM+DcclAi+N3Y68n/U/WDqoamBiRTaeszc0
+v9/dt/9DdBKhMaHOc2tFOhMM+U/y3QVYnaVEDHLOEKfaTa+BjNaLpE7lMeo+forBn+PQr7Nk8JD
Gfhs+pH6aSrNRR5y/FFRlg8w25Sp0f0NkIV77aHoJ67GUx8ufDBV1p0Oa6a/WJMbBOQQFEn03CYr
e+Ow3NRCFwfKQQWmD9vDiEsML5jHk2Y4IXnyu/KMBOzlbyDLlfz+mg2TWzbzw3NgU8kf43NM74Me
fCx+ws2Jjw9irSUAyQJEwXJrFz0JsRi8N9+dc/mxUJeM3n45A27bP+lrGXTmzdIIj8MSTCy8DMIn
0wePoTCjSmHju4RDSvk9DjAsUOyqyEKyKJXUj+MSiR3WPljniIoiM5pPT41FaoanVK0WKFqcyLT4
njYaqxGVtg4okpWiayH6XMWTx22M/+gWrp/SudLtHHOAsF7PD3TE65fzuBLhFvKR4sNElBXPgpAS
pRskVkpt8O/koE9YKlmlsZQAnw/vgLSvpitg58p/rVdTt6uNj9KxzGvuN9vg1d01Q4GKAh6AFYZ7
MLQhdlg/+A25UPoFRbJFpYN7xyiw6WAZ876hSQW1tLr/CnX7EIcitBwd42e78cd+d4B5lVAGxERE
w6zxnxLccNDM4aDakuh+wSU+O9DazmCy99pLKhXaPoN70mV5z4I5nC5RUYwp2f7NBRxT264HIGc2
OQ3xUSIsifIRwm4l6h/rTY4i+XdyHv9AcX2SE3pXtxHci5Rqgs+MggR3TbjzfT8cmOOsjAsfhZPi
ZXNVGOT8cliZM+JRBMSqwOh+1oGylnnXr33Ul2lgFDCWwI+1PqOThi9q4nhasmkgLxksOxjNinzE
C6GWn8uDiTCASEkkfq/FOP+Bndo3Tad5aNjIUjvbQI3BNYVGqcPSjcQQqP20zsPj7XwH9Y1qHzZ+
QTUPE7yAFX2Jhx0FMTTj/Brzwc5FYq9/HZTELA+1fKsApIJZWf1qNIo1mpyPwIFRw+CRdAq4hmEb
QKDVeTxV3HVt5+ot2eMB2QpZk8D6Mef9mF++5aB52H0fJ7gwq9drL4KxPA3WE84g13IhU4CQ5VCA
2SA865647e+KdYkBDmInXBktqVw6hHI5cETf/MLU1wyCwXB6PvfhQg7j7mOKvqqgJih6/c+GK0fb
xMlFVUXKeVRmWBzV7llbJsSmKHbI3akLKsR90uBrZKYeVWmHx/I8yIV60B402hokLhOv7gFnQ7HW
8SMhoxOD2hpADNcV1tTjFmeJackL4Xvsz0cEg3MvS+RibN5GO6dfuiboLUh1rF9mFtT6Qxtshflf
7tsG+RsusEfoCUvKe9yFHzDdjPcFpHDsEF6eckLBw1N5XQqfPKz7t+7TDKA3xXT54/VecdRr34Wp
t7YVClzA9eodvdjVyyydOjUG/Kqxyi/Jy5+SFku0CaR7WbSZWZOy4YxRJnCJJT51uwSEuOE8Azdf
wno9abQLibcuWmsS5RvXdqdGJmshQBNjP1CUFwVz233XkVg01d4UgxaUNnaCyVhtlNiBMqeebBRI
0SfEks3L1gLztZ9hsC0pzeGy9PXFyzu+XrZ3UZ2kb2FDUid+hx7lGj2wVRFBQxEuP3X9S1NiwZIK
cuFP1M4FNbXEve0JuVqsFbz250sTFQ21Lqduk2cpf0jU9rzgMU3KvQmRFhzhJt8svQ+V8MbOTt9v
VHJ8sc8rtPq5p2WXTDqCG6x8XYM1dB1BB5RnXnIAfuZcbVZZl1hTyRhzzDqPiroe64bBhvzoPKxM
ZT6GOuxE0tR73yqUp75/P9BFD0zJfxjoDKn3aw9XDFiqW7SSiPJRB3u74sQsD+x5/G66DmVAp9qe
ysWX9exKe62OnJrg0+ytAyr1O6HcdqFByBLatfYYKuXATxpIcqXtPSpklYnOcGnC6rzwrCUaItHK
kdhMn1BQZkUsV2IYH6UWEwWbQjc8T8kzRvzbQa/36vYrQDkhAxAG81+MUm04GXFn6Aros/oYo4jF
2wPFvp+BXghHgs6cElzm+WyMV++2lLI5oWOCt/Btf9Y+9FgFgAs+YILpRCbfHzexLWzpxLplN7MN
LTYLcFPWU1AYKTMcwNJiVP7Askz5u0xb5X3kFQIslEpr0ptL8p4iaiDJC9nUo2i+gPhomo8yQmAD
urvC1XEUdYyAihUVUrdlhPb4OwrPrsWWYxe3bwEfawFnw1xRQ4orIemt5g7tx+T4FyYfu4EtvIOz
1EOAgQhCPhrvtQH2HtRctYI0WKi1bgqy69n6jBtb6b8GDdVfc9KzQ20ptdv3jYFzOVCBITq9Xnjd
Rw+NGR86HGjDRPRUKObXM0JozHedCHL2CrTG49MpLKpa76wOeOacELACbnhz7zuM43qMg4MI30aI
f0qIvE3fKc95zeQI0QjSU+aXUT/fevu774QHrc/c5EShIc8tQ31VXhXVDj6SI/kxQHNfXTZ0x7nR
0kvMM/Bugc1zgYIwN5j9EB3owCxkhcKXoe3xcdkLLhdnBBtYO1GKWASjPTgHkBI7g/ONfeltDz9r
2xGUxl7rtETXnGYnjzBqUZ98Lq1uHPtDpeZ1UIUg30+AVledhfNPuq7BlaBSZphVcbG4nseHwLeC
+tnorjw73m5XdnR7BSOwqqpo/BVHG4soQCrrQzIDmQ8vPwpXE7yAsY4M3XvaGjqYeRbV6Pbb+UE5
pU/VibxRiQei8IhI10pxR1IfRUS6HwIwcZIEUbsne6nKSiOdmuoYwJBZCpF1feH/0ERZoYpQfKTI
eB+EXHJoxC8UZp3UuK8TY8TFasPfvIKN4oB+KPo2NNeaIrxG0IhLAg+wbdvonoBgNW8J7dYIfrQh
qkxNgZP6kj61RmgEb9xR0w6GTWfQEgW6hODiXBbwZGGr5/4G/Dh1+O35gVVggArcW9dhQGTwr5Z0
XHBquezLw49qNMPpyLXl62nJ+ysqfsDKfAzNTHYI421UfMvvHp9sQHCC18ZM+T7r5fLPD3NoVvvk
RPe/AA13bJidr89eZ/LLsNcViMHO6TtlQkW9/EWbPXOUxzo/w/m9tuNyPPLYlseJWLrMObymF19h
uhbfdmaYGU84Q7RGM/8qhShgdhoB2ZgKUCMWUtqZ9f7RxU36Ch3d2wZNJ+Pr4LdjcVan+OfjvXLc
LMiAn27MwTdx/jkLOqBc3vpYeGuRKFGHSNGTzjchCwC6CcDRy75MwzDmzK1IskjDWyWvcYMalcpp
nt0CDYjJ2tzqfgpsqFbon38ZEB0pbPUwDjTrk8UEdWI8++JzRBcVbUQPOmcjG7wgnX5mUXr739Uf
s5gU+/A+gjpjnZs61Q6r0205gKMuCCCdOaeVdm+QGaPVcH75bRmD1/xGAGRMm1S+Bc/CoVJSUQhs
8viLY74dJGVMUJq6BmLiHeONQI6/59nXdgizPc/6yHEqoa8lOPgsqUeqzbIOw8MrWoqqQf07V/lZ
/UkM+ZhIpGqCPfIsQCTh1A20epQRnZ5S31DAoiAuey8lmIvut76qqVMGjFulHES3U5nxyp/ibPuv
RvPHCGwtRBhVHOjdfEfyV8kQ7EfQPtahva4Xuzxk7n4234Yj7Fw5NB4IiqA2UXMFSPDijCghE5jw
z/bTG9d8QoNUWEtsXEbXQcGM8TKUu26lnn+Sg7KVOiwQ+w0pKQqZ2qvHYVWQssF1GZmrJxbNNyLb
eMYJEb7MS0uDAR9zRvZ7onIH/1UN3xboVcMm/oxj2JQ7HHKXNY7ZmvUNIBcA5nGC/kZRGtzWZN6y
jqXV02fxFBSBXkHHDhFGbdCFXncLHSuIJ/eQLGaZ9xPNkjbAfeFOo7qvcc7Km6qhbvhzutx+kt2e
DXh9qKTEf8W2ayaLMMj9GpiqLrTtR7GYwhC5ouE6DdlG0s4ps3ocIM7ApXdQ6NRfQlWfOY11ZMbW
sl4Q1XWOIr16XnhdBGtLKoQihfyJ03JnF0Q7ctoTF+8asDmJaRk00JvWps3cJIjzdy5pB8AfAZ82
ZXsJnTonxYEx5c2dnDTd9kZjJr8rSfshBXFllm3b9AaMSEsX0K/X0/2E75DlLGu1b3PPjBq/DUMI
psowh/XPnPsAVOTS8gLO8KPw3jldxN9zh/yDaaIwmGsTsSypVMr/Y77hIoCe5gmtXalIrviwAhd+
1T2cbJms2lM8Mx8mpUzYTzRt8p5SEYd8XCTHhrFKCgXD3vwFmJHypF8gQP05OI4zd/SnwSTaznEj
Q+nWc/5Tjkojx8c02uBl+3CKaN0mZQt0CEDSdeejApJFmRYFeaJCwFFRsHK09kZrn4pJDUGjvJxi
B/DsRiKBt+15QymgxxtFNevIVNqm1FIx0wrOdzME+EHEgR6KW2q9lz4I3nSj/lYmIgPzu3KHtA8D
x+V+B1sl2ioVSuENekTibp6JrSYpBDYUybR3ZQzL64mxjQOMhwwcSynI0D9FxorfeY76D9OJ0E5P
x0/38fMuLN3xZ/uqY/QKELyxFZ0oY4rNjTC5pqtPMqHGH4EbqqoiyFopcDWMaeOpn0NGCtDLhZFj
P04PVIHDDSm8k5C5VFFOOr5ig4A1+zjKgOxsU58XiZEDyops6Nwde4PN8AT056iMOu8IPBAfvt7P
tPJENlDO0B+ZhkXtV21L4NYuKbm9i0MysWAKFOGMyyndgUXQx14myqpGwLGHSzOjFdMGBAOJ94Rs
NcaqgB/soD1XLQfV7pvqLdcy+VU6tWvaSQvlBbOQw1xjTUbSHR8UGHKBgqQQTUsuEIXJsk1b2Bm3
1DrMGXs6X7ybsE/EVvchWBd79B3Erec+pjwVsL/9s+ugVGPuNvDcjH2JgJDR2QvjCNLSxmGJ2Pto
+vQKppskaRwNxt2jB8Gunqxm7meIZxBlUVAz2LMTS7BX4VtcksE0KXabsXj7Fm9jCvBr2De0Wq3l
AWaFr0BWUdXFttzhT7Seml/wX/FVy5MJ+z9tAmse1vI4tlfoYGhLk7huCaS7MV76p8Z/7yGOxIZc
KyrpbauhVZLgSWqiIR1/tr9opijlUFTLnWMl3TogQsLzlMk0pNsAuoZbEE9WEm4dNAPYiCP4YNwE
EamLGyc5s0V9YyIOLGZR2817BrOQUuz87LdMp7elkQHtUsWYt0JJun5NW9LErvWPddCedVAW5sog
GhGPW9dfHH60VqYbqnxsgnyDyzT6veAj1HTui8qGNbA/s/eMgSaKajWTeYS4yyOMVyGwckSzSc3S
BxApqexbFcuOIWtnLX5QUu/QYDVQkqyEwuu2PBTIser2cYaQ2TC1ZKzrpVRBp+wUHM9f+Aj/W5dK
CGZyk+EonfjYIybv+b1/bMmxTrpUgqMRKTRn6F9NUS72qDuChBS4ZmazNJ0TBql2Apyv+vx8TjH1
4WwSBDj9YaJ6I21ZrYlvQ6+VKIcwU5qDsUHzMwfNzpRdVlZ5eDVc3sM0u60Qcb4gfOq42t9iN/DX
r8dSTX4f6/xQHAaQXkzxUnDvxVIMSIbt+tDsNzNSAueygtolXUS4/MNRteUOIyZkwAaGvGEFql2o
uFvXOC1gHwr335ZHam08M5l8NCCmGl9OptQ6QStIMglrsiGB/WwNDcJbDxLbFFUIZHJAXoSSYljm
JU/NGXqo6snaCbyVVvrfy4VE+yhwOdCEqyEXwyYNcde+rsfmAmv07cfXFNXXXrsLNJNyfdDe5Uyq
ncGAnlAmra26VrFOjRnrAwgm3S7+QGAreWKXKksa5v5iH0x13HAi9R2zhZX/TuhLeDo74ipjpxyK
hSyU+8nxfxJ5TjaJnAe0YlP7zwj1TxtBzLa0h0yrMJ1vcYSJIruGWMr4HNnlZ7sivTn1wB1iKcI3
YaSwiaVG372mdSAIciwGSd+NXvdlnWfptBuT5sgbqyFEKihR4RjvC8vNmiYcjHKgkcJ/zXbcz6M6
XGp3srRXw57nf/Qxj5nirYYOcXKloH8nWJErbeWTEOQcuruRSvjLvUjnCqIkMMUTu9mF6f3JdCb3
+IQmFitdENg+SJRi0ehSgEWCxanplNpMXDmk8zhqQfIdJdS0KGwFw9UvELIZgb9zmQQ0ebBb3b8o
psURbcQKp4vQv0Iq1SfD+TweukPniTJS+I6svOwWJG9xUXIwg7WULPVh6d1FFxAjj2razyQNqgba
uZyR84hoB/g65/KnjlNinBrFixs+3G410ofQv9gvhS4DNvggO5E+/DH+nEwX9teg/ZhC9Hkt9joe
7hVbF97M6K1QO08T4EGdgsiCYAl0l2x2kO4nc9Fj4GkPPjGGLBUBwRNh6+fgfx1rqvV6+VtIwPxp
9sBYzW52ndOzmmW21UGjfAY1sWTBy5suMSC303e8mD0enA19buCy44HvHuWVRoclonKfPmdrLwv5
Gldy2TlyrHn4j9SnUs9zWdoD9+GZJVzolmMBGHkp0i4UxmCxoWr1yDhlre7rV72LuSJtCK+7clL6
91tneKnJ+5dCwlOiStLJuWn9FFhSJXI+UPvA9xMmg8l44ZYusMAA3WkpFutJ05wU9T982gjFU9RY
pyuo3Psd5qkrF3xbEPmIeUM0mNgafYm9qPKpHJBzPxPtTxUSPg2D5WhVFKqNA354yXHXJJRDNBGY
oDk7xJsr+HQGyBQjyQyfYo+vMXUHCujswP0Ca1gbW78jZcCYTnCFIohRHQOOrdnC2tyaN26fXtkg
RMiCSSO5BK/37HkS3tX1RTqIdpVkJ0B9gfRwMARNGFlTRdGiJ2iyfY1tMEQHTHTaSnpV9NIYbX8c
XMLDVPztLTc2J7RVijUWYFEC67jeESgrtrJLojqIQ4QXGAZKqmIHy9aGvp6dU2E2mFvspOEPutxI
zUC6z7jJYr2efvwl6/hbpRrC9OQ8tsSIgx6C/OopIrn5LODsB9yZbDNdBH+w3p6Tf/OBhKPaeIX9
xxYIUkj42E4v0m6W4BWTP/e1u/qBfHLHUXDIcrHl88hD+h8AKBCqnmaeaBo+XDZHhZgI7nnfwksb
VRa4PYmvoMSrRO1Kkg8pYmCbVmtO+bZ+tpa1ZBWoyoKNj5LWSEe9P/w36Bk6lyvYX9XxPGnyCoxf
7D2FUUGL22Y0PpWgSSHrwvro8L3rSzZ3vbv5PGZ/kZXhKkZhosqjoXFDYWNav+UpYSZ3rLRum69+
O1F31XWv0lI2xzRnwp/Nnzi3rwsOtsTLdmu3eiU95PwgsiUvl5JZctiDY2doyQlNV+fW2dmIpC5Q
oKd70dEXT2y4BpyQgkOcOhnAYBeB9jZMuvUdCfr0Z0eVDhlsXmpjyDZRLqdqCvFWV6v6hz+5wg1s
XXrqZ05IyC+fFBqAhg8gapFpR2V+aH4ojkV4xwjKqcIcxlB7pjhf28uTdDAwJ+cURfdQLza/hY85
6rCJTnsKBW0L6Kq3DCUoBcGN62LqdlxbAyyvwqhJKb4XWGZNN3db8Phk0V7kJBIE3QoGpm6ulnr3
ZWXqxBHgtt9GPLkPmaXiyl9SknGLr6bthVgfk+sXhvSMeC3IIAxJI9WRpOuCMyLiKofraOpdah6p
QI0Ws1pHeAa3cC+/jNCu2ZuwbdQZD7cZAoV4wD0SjbedgpkeFrf9mhfpQP6PHHZHtSkrQoTU7H3X
uwoZEL+kya/3RUKHXpfLZnAo61qt0labNvG4bzSvs+oYXFv4Vq7Qy+F7IUsVvhzIxyCD5SXjwKRS
6wjmidU33ZULaZ9NF8o9Fd09Pt8zqPZmw+YQzzjwFx8iHbnAa/ugGP/ZR+sOGxo6E8ZWXyjeAspm
o+kSMQ986B7NeLdP2VSkmEBPRtrLeetDnt5531dwIuokJ7PFJoJE71b0FI5e7sk3c47fGpULCwdW
wTo3nu5IY0q9LLypFJ1s+NQ2nMuuHCavAHB5Y3lSS1wVIMFjSwbbY6Oi0Wi6cRUzYbVGhHItlsJ7
OQK4QzWKaTIufQ8dkQ9hIqTX7yQfDW3TRPnHpHrDpYzomt4k/ye4T4DUFOpQXOycv4JSQJAK8/nW
XDgnzBf5H8RRKD4jNZb7t0tiV5rjOFifyzpAwsA2IzzlnLCPrB7qJ1XJwYxpWI8FRbN/kgM+SKor
nxUIkUez2bPXNOirui2HWQFJ3Nzu0sLWBES36gY4RgLsTBOQ4lMLZkT5JlruEN6k6js0F+Bt/Z87
MF17qyCMXxGLBzNoKzZ+GIZbfRjLjiU1UbCY5gqfwcwdDBEi4iU+LNQX03Ds5Osqxe7dtOnXiB2w
vY25VUKCZ2Fggg5hWvHL+HWuTBFO91abzfnf/Kd9V499QJof6H41D9Xs0c8/3UEPdOu218yVOpr1
eNTVLJvH0OWwklOljhaFvR+RV7aIUIao9TpvUibXO6pXQ1lIhah5vrBVdj0vW+wuQgJgA2BH+FId
6zlO679jf/Ubnx/0jpOegJkYVH35LHlcAPQaWdOQAwfEj8ybFJm+ZbDx2H0QQoz2ahPkSHTzBKpQ
6jOUJobkB2F9FjBsRKTz1E2+F5v5cePTgWxzQk8QnJApkBiwXq9H72zPnh05hLJkCOTRwaUMlA8/
sC0iKRfeREPBcS3AeTFy0355SHa0y7w25iZpt5rWLPRox+EXNIHSjwY1w3Yixezbpmna6qVFcXJo
mHh0W1lYXXVp+zVZ8Q6vR41GTjNiEaNGe3xYPsLD8hE6n3kjM2eWFFozShgMPvOb6TU53z4ZTaJt
E2h+Yr/pUMcS6Y3s4DsBsv7+KPQa6UZLkylKYfEt0ZHS4XETFhUhE1l1E+gvZ4f5NXIvu+u9kzGW
zJHKWenWFHqBnicIWyh8d+CgjtS097rePS2rYPqhRsAIosQqeD8eyPB4rtZsCxTczSerSoobnZE2
MqaE3uV2bHy69kTZeIbRig6duXIhGWoff3OlSG7CA3E7iP2Jr1Xvjw9aGSeZ3WtCOYSUtaeaPRvN
6Lxb0UpVQ2ntMS1xXBEjtqbHA8Vh20pmni3tT8uM/+M7A+t8J22g0wRCvYlyP7xIw3x2xvcYa0fE
sH92MUlj9x7lFvKkQ/jtiYMjpWOKqo2HMUuAEiXd1RmVAVxn2z/y+UjMRkNf1OVPEVwpJInKRCw7
v4gHCmnI60p4Nr11FjDxj59PcR3uv/wKOxYFflezADa3jtPzRgFoTc7mWvgARKdBPlYqdwemCRiU
m35LcwMdqvKOn9PML9LAYNL9Q9e3MDCohZ9lOk1HcvvGGLQ6qr981zHY0iUEDxZRCIbKfNab68JS
qF/72hXs+kk352iKuPUOGPqamPLyoT/LIUbz3kQQ6jCBTyPRSgJ4uUrk1A7qpc0FQNMq1MPHwuzf
+XW5jTDOCVI+K0tCDKdBo+GPlEf4rBGzqMLB6llbXilXkpnPlp4/t5bP9mFCgcMV15gk4B/lGh3z
n0MjM/1w3waz5bFb/Lj2sTItTyv6RtIjqMvysh8M5qgT7vb7L11rUsxCDLz/r8AXEZXDHb4uKGD8
rOcxF1be7kDfnSHYFv/yIws1JQtcs2bNiHsvKwjmc39rNX+S9KKmKbe17gLtOQXn+9Y40NqfXLwY
OIMNdvzvtAEYxCgOIyHu863GDdINNvGtb6PPH6g2LiJPkxYw6j5Idd69jk7Yniutl+BIx9vIVn5E
6WsM0/2ifpUI1bkpqzWOKvZ4jaMmu0bLLCNdB5+Tx0i6isyX5fiBkJbmx+V1HP95uUBOBll3i7l3
brCbttcpytFbqLVB8qiz24unLC0bsqwVI70satK9C07dh6UTbMShwCeZ1Aty9KsYk1I9shQVBehH
zVXYWuzSKThdIKj2eOAFS2ZUXWyPV1UHz771gmgpSVQwbFVHIA9AW5punRqHyyBXGV+8C1361H5L
tuyGNaSjvWZcICKe66YyZ5OWt7LOzuR8mE1mqXFXutQDLlTjUdI1chm3KsDnVEryZmCqo/ZHieLU
fHhxnxrkmbb1ep7MmhpJbQ4txysm1XlqLsWXbVgpw1joDSg3E+6+/NaBD7IXqummGh1kNXpw1A/n
QKw1x185tI4koXHaEtUuepwmc4U+aOJnoWZCZWDM/9cvaliPgWVlBUsQKliNPS9tk2lPLXd9Q+aS
L8Eqzeru5Z5WinLY46tFbEdEVIvsiFivyBwKbhuZG4WXBuBZC6ID6FayT9x+Gg3aJ9gr1I9gK3NF
m0mhS5AwgXmJt0TgzkCogAR9S2BAbVv2JhSFjkBX15gCPWhn6uQEVim2KKSvu9qKlpemSrhhIaSF
xSN/QxxWTnsBitgvIAh9ZExVuNgnE3AdpysxbrBqgpoAiuZOha0YZIMR56irb5SCn19gyjqfiWd6
uVzii/wdgEXzb9LchVTnsAPumd+05u+ADN+i7KxwSTWcFv5RAPQCueoH7i/SZaAuJF9SPcGvn9AZ
Fa1/s1+xhxJ1y1/cFxdh5B35I1YML1hDwvqM70dTPAm4GnpYzK7FrTYk5ICNbYdM6HWdGMMnjCqz
Yx33sbCTSIIH4TnR1+6PPEkVsKqcox5SGerPy34sxC9zEP3Xm1PXfEm/FBjjtwmUEpaaxJ5KpgCJ
Lkq3IrcwYSNDfKxVYOuURYHl6rcadOORxUod/F39wwI+o9biyWvkP/DRQjvwOemfLCbXq5H7Sg5/
vY1mCRO7JghojLUJ8r1Bp4WCcBr+NrY49cE2JRKWXoUkW5vi3YEfzbUYsiGKPrzg9fDKfmTg54if
qODQknUKENsdIipo5id0VonEoPLLrM+F8EE+hRCdqpUUM3XvvDE2yjAJGX3TW3UvnNkeWTNROTGi
+7ehzArNm4xkAPuJTbObsqtKE2rVGvueZUmTneJX/LN5XvSjf8/BehF5cBNneDCCo5kQO8cKhlkF
4nahQKTL2MYMZ6reymTawE7O3Tjn6lIBFaJvrBM5LoUa9RfgEF0YKpWggp0q2XaLmeRqEwCrw8rV
WLXl+jz/ovS/8MJNOfwVAHjSzbXhwmxeAkUBUyMb3pWWcnl+5w0vEg9J3h0kzi4+blhZM1QADxIp
RJkwl+V7cqgvi3QfuQS24ZJkRLmXPrJybCeCrilYbJh4N7JmJmmusOUnDsYhDUP9Oij8hriGk+yr
3yvw9gaBhTgzeqGwioLRZFuqGTtrZ+l5RmKl9jzIOXf+aCSqY6qia6a93VDSnVLf9z6ClpdjaXr5
5dejHrucRrZeaH0oB0vqg/PHZwIUMLMrFRIcRBWHVX7l4xZI7SfrQ33dfY54xHf0vMPRPQHBE3/7
1O+0iWUMXN8Gc9s/70IJbbmACLypDVy5Qjc72HEfZUivICut0/RDjb7x1sF68FqNm+zngJ6rUO8L
sfoiogLZHYdq/8zPUhalw5KPWZLzUfDMQ3w3t78kfrzqRNAzDyQk2IQ+sAujjsUdTuYEce8FCmjE
4jYVthr33Bomy0ieRXoB2trKH+zjuYa/qGAjYQYimiHCDAMf1/OF0IQ7zCoOQUWb9aiTHBrIBylU
x+BlOZJQXzc8iG4Se4zO0krqrsW1+Ky141vrGRAb3Xq1OHEroWS/jnN8y9G6tURAVxCVNrcMEhjo
ncrMbOHdBNQ3mJCIHFP1x8Xh56xnhtJltOZDJmGFGTRlZlu65EP/DlxIfAlc4LlGIOUmWIEzJpyX
A96o6n0R1Pp9XKhds/mD473bOGlw80bETR5PIDgc0m6zVbWnPagslRJj/xFYaupVLPo/s5CEAAfE
bEI/jIKG2/G8NlEhG1lKjySnZZ4iFpbGg1sDmaGQvgFfN+pWQRLxfmyDdPf+XsCoK7K4m4rAQ8R+
4Dw/iaULPibXbikYFLRksYB8OeuJ2LZKHxvhhh299cnO0D40gP/+ZzFSFaf8SqfpGd1LBsXPmEiF
lwu/c9/8VxEYuNX8o7dWqTmXNxvPL3IgwXGeI1f4ZhqvGecfbXVHmTvmnyo9HiD2FGSRNKtRoR54
grh1BTk3Ar1RlN9bGI9boSLfzgoMTj4N//zpc7XxoMIks/0oL7ixBOVZGeAGm+HLv9swbpgiwBY8
6ovdUOktTHowA5vrnohiJlNSlnZq1sbDdDKkSlW0+jJWH53wbh3K6adbJmcZ0yLA94tPUcFtLMlu
67mnCVrSLMsFrOwh0wkcUNVmyPeza4R4usZAHHDDDi130mER1lhgGTxJ4CsoXDcLYOzngbMbBK+4
UxT9l80O+wLX+SAtRUBkHcU4vqdGa1TgRX1LnmvY2ekSyogHMSklnMpCMCo9Avm3r8dryAagVU6z
l5XN2wGPKaC4Clkkf6PuSe05p2Ws9lJcKzhsMyHOHL0RaP3TmRVQaj8uSVWGmO7f7yXyM3GUS2F0
qtHZqqUaVORawqtV+GsZaUaxtiIjFDBsAb2kTreQdddhQ9dlW9AJqXMIVwPWm3I2s9YqTVL9A86O
ltHEgOsA+1Vzi0yknYIdJhUhlNFhXQqqaW3ZlaYiBMOwDH2wtqyBcEG8SPhvR+Mfm7b1fnuyCp5d
DWR5QVzLhkTM+hvpLfV/U9EZ+0PXYynR16L5IlQhAxXdA1iuSpmvLqVEpx+C00vukeD8Mj3d/39z
NXXHSKQo9GvGfq2O3cRyCFgg2sNKb79kNrDgtjgLQxz459cdcubcL6/YztLnTJeclbxXIuDgpAZt
ctBKdacO39VB3c1/nRleZUR7B1BNDswmrMcXFk6NryKmeRDVW36lKmeOFcno5oT4jFofhc6B/3Li
BwUB0aksg4fNYIQ8lLYKnoDlVTEZV0e0t3+o1HCq7K+qbdM/3gJO/ADC8hIko2RIdf0fKhMmmP2G
kxGKf9VnOzXM6DP+G2efwYQN58Z1Q3Rce7sBfNIy7E31PN4gle7qurtWU8B6ILXW8fhBuqb7Emje
hr+3Q1wJ1UTvOb5wtd9+xcnHyOGthwLLm/srgGhIFhtsQuR6oHXQYVV4QDEimfdxITywi7D0t+lR
ssZc9WJ653SGZj1h5T2SrYCGFRu5JObcq6pUiB3w1D+EUgh1KE2ojT4I7UAhGcOjXncm/Bjtw9rb
F2K1xMpmIaeXTMi0SlGBdZuSeo9jntBqlJFvhi41v9sEyY/ZT8eIhRVx7fhg96SX2CiEdDlXCZgk
6HfMA2QDFYg+RzepxtcpPAWvxvnffvzKSVEE3RlztEYrYuasVTIfDQjEYSZA/5mDFmUgoD+kutX9
A26GqG3HNJHDoi9g6iX/BQiri8bbHVwALFUXOb9T0j3CuHNHvwcNGUjkxhgIcI+ZXzeNLg8TC9P9
PKA/5rjVaM63bgHZdJFgVQkrgBs+taonzGtbc//4ji5eGt+6GMcXxVEgVQNMa+8zcj/jxvMPyEt9
7k5KBR0hZMS0w2xu3NxloSzqxCpA9DrvMuRXsYPIX6EU51rPdXt5Pv8T7e7mPkXIpfaMNZe0RJQ8
Yp7j4E1EDH4BaQZxd7iUdOWtNwvvMvBGVEENyKLHZJybdV6/SqKAGyrp2TZEnwdmOeHUAm5xWyUM
Ss9w7rcPPBuNS3T1fU/PMdTVbc9ph0JWkn1kifSoUSgvU7w7czX6xlcDrefYpY8HVJy17f4U+c4x
E+Y6U7VIVc1llTgMu9sn9GYXmCKc8UhDtS/EJ3uUG2BLjX+B6e77Kn04eB4Rwg7esARci+afIyXv
F+YvhQuORisKlykeNJxPgGl7hKIigOSkUeeiKQkOQuTwrrz1qrQA0n9TyDLFfE2WpdrcbDY6x1yg
yXRqOBxAFFeMev+y6Ft3t7GVvXs5IZAsHo9i4UzO9qVNrTBkaTTsp8KdW9TYCYVM1Jt5CTkh2mck
rII1yCbcJCfgH4E6+Ps27PRT+tQOg7zsgdDBh+ETkAc32NPiC8eT7fy04OUZlH1Z2LB9T9XIShQ1
ogt2rJuailQNCoFx9tC7Mv4EGQEHhGXtIUyIfhof2/dip4dHTfuHaBoEWOhW48aMC59im8n1GhNU
3mLVVDKVM96vD2fS4j5XRKi/305lXHj0sEhRewdALcbrhnAUgzlKtLj0nqv6ZmKSRf6iQtA8NIE8
PKD3tSQX1tsb9/sZIM7YP6sxo3UADKIm+K8GLo5RfZygoab0ASiwm7anulmr2SugWA3KOJGVvhkW
qdmWNXLn36ZtlOpN1ZoOo+DyB/ez6SFHmuYTnFDXJ8dEqDDnx7uV3GDB8HDUHx/2bi26BXnvdx/u
qY8qud1VdRgG1qZK/e94xt5aM0foziLq8eOmwp2caA26uFAdnogxet/Tfwg1+Twy6/KM6OWp7oHe
ADSgIVFf8F5vqHZXwstRh+OJAn7rYbl5KP69DSdsSfvOjVOUWlcUf3BAvXZPXwmfFfvQXmrET1R5
1EmlQLTZAFamV+jbczlWv/+TFG6YLxR1xXnmVjavea+NeqxcVNG/Z+C8x/lgYEVOEnOwNSEpnktM
5dT7cvl/CaUUEwNyXQwoFGjd5HMCAYnjZeQEB0xWdaUoVSNd0hTkS76CVGpqPyYB9BKGWr7XHlMz
F55SJ5Ci1pUZXI4PVo2KeIJVInidA2JkvZVv3gQOfBxoRzxSWQYK+4JInm3lkoJEmAKX07L36w8+
5ckPLAJVVYl8cOH9+6CzRjXzo55tbMUGxPp4qagPLz3v3qNs3RXZfDqzvQXYdmNShMrS0tyWLZo4
eZrc+VupoTZPXOYhSL/c1Ta2i2aQ4qi8jgOGvUgNRx4lZkyLUjMtNiBdNSvBJsC0TiFxIkzRGk16
6WeyiD0ezpR491AYcnLtJ0mn/JqJHAv9P3FGHw9E2coVi6kqNtpOMLZCUJLgtOP59uYNlSd9Pdva
jLapppCh3EsTBhB6+AROcWJUItun0pgUO41Dzo37xU2qW5OvWH8PR9aBPOXBzVw3ovqvoRQkWMqh
NYwyv/QXQm0fImJtKEv3Wv5bYazolaIbDWG2ayNMd0nWllt2O/k9l3AdbVVY+xoXOWVDyOjHgFF8
LSfm0lHnPBAgXB4LhHWkLw/UFKgVNS3p1nqI89nLYwJmvYbMk03QMTHgpFFNicrZx5R5+Ls1RHZS
DpNE7o0QujtiOZ/qtoSpZ8QeIv5cQ7htX8aCh3HGQ9n063rONYUpodNPwQLFoBsA5id+Ci/M16Xc
sNuY4hXUgCYu1l7B+oNXT+F9NPKV6N8tO/eDaUamqvF1T8PNA1OSdxKw7ZZFGE/yUjRr2UrBtuO3
L3sWouQCH+6OU7V+Va1fUROkJpBY3t8XC4unUe6xcxnHhmG3aUS5K2PUlo3i2Au/neemw15nmKWN
Cesx0ewZf+FaqB7pkBC/id8V5sw7dsOZtDQmHXcNrr2NefNQm7Idvetqi/4JYmGIfz15WEj6Fik1
wo7NBSBQIZxbOKagn2bi02CzBqVzD2MyIgZz27VWIlDZg3R+G18NcAVsVTk8y7A9o4nJW7eoNnFj
y2g+irYMmKRtpJr62+Mw+UVHI1QUtZc/wXuZfKVPkNjhT/XYuk9VrFPqgOSUL9SETZeV5GCe3DNz
ZsoJ2rk//+aStmXXVpcmM9keS+eowmbku7v9LzLCT0I87LuktMZdHS//VhGVLJIaZ8QU2k/db5ZA
lcHBVxPHiMP9CvL5gp2YmbLwhpqllkV9v4xS0Nwu6Y/Wq8EO7iwwEPGd/c8N6CH3gA83cRQ034bG
PdILLqQ6TUQRnmlFOq+0/s81cZYId/VdlRRUtxxZdj1131NFaMh58jI8cmGo4YZVwRsJX/3/zWxi
3DIxzH/X+gpRML0JxQKP4IioLxbXFcqkDfzCQbjUTr8p//165C6pQbhzkUkeryk9xbyY/zWczvMA
mf976XrampXI/3Rlz7MxjLNU54AECUPt5AIMNcanKG5L8PiBnFy0PVhdcOvwWg9Zd9tDs2/Riry/
mUskwDIrKKAwDS8ytNYbfdZ4mHIVgahdKXmFhmWIrvVLRBJ/b5zuxt/O3j0KiYgMyPTgwF0RE5kJ
ikQkiL4SwHQeE/sZP2giC8D/HHVuy8FeLpuIzFI4kVtwkv/j7Pl5AGTb4We3mTPT7EkUfQJqBFuX
eipu5eUjFcjRZmKgEBjKFRqVjlhlKtXmI15Rvh1QNNgdt3tOVyNoW12I8G2/l5qyGwjSVzfGa/jA
Oc9p+dLEoFCsts4AV9j967ukhToyf4LbExaNZawe0E2Cu4jFPZ5TZ8DeQmtDSFD1zcKTeXe7fTOU
ujJ04q8Jd8x9qewS2EK/AbgWyTjq0nP1YuN0K8JOmiRBFvn9vMjKp8G1wGkysl/6nw6gReAOgESV
YuAdDcsOjhjB23zKxJJ++oGQO5uShsN05qzSWEZ6P7R35rKU1QlMbbJooMXu2nGEW639fW+PetsP
Oa60+cs2DBayVetZWS+O9151bB6o5WsE+uvXjltANIHlsV93Y928g5syVGgC/W9u3+Y2/NHec1J1
eCMILABJBwHPR1indvPAzrzy/4lNfEc0xuUBnhEYv7weQbwi+/SwzD7z/Gv+F/P2XFl2s+LRxAHZ
G82aO9C1t4yJa+TLb2nYxb0Du2zG9MDOHxFuhek3a+RtXC0L98ISi+23ylBimNJutCPxME6mYBqj
Y1rVORmAchk4wwwL8awjsfAvRmxzyE+FnGjqzYgW03WXWJAyZVw6DcHKsyEveaObkRilEp6+dCD2
z6+kE71atl/mcUDdv8mfLK7g3eOUEOibgr2/ow1evSGHuhL5u+zLVwg4srUZKeg/60IsRMe7/TVM
mVgece+P6nNqWC0WuqLAieIH4YZe57vAv80fq134u+J+CqN31YYQkmk+ey2y4T6P1YZvFrFy+L7e
cRjkLqPnklJDfQnwEQ0Wkb5AQ/ok1HxDuEMJ5M4wx+OhEWVCv0jmFKgbBVBHb0YkvGy0Tg5y4rfM
TiVddX7NKwkLEKu9it2z4yoz0FD0GcL1iZckTATn4Y2Saq0sSvJXzPezzU/PbhkevJIleVXpU5kl
2Zxgg9VH6s+QXh4P8NOkcmKkb3QuzTV0POKbe718mXRy1dP9S7jL+2FPMkGLip1a0vp2Hr9RA/NQ
uyA/Z6UIJ9iQI+xLvraqIRwonDXm1EsmgWGci6Lgt5x7+Kz/iCVeTbyyYXXgqJ6PLMTwHtEOdHjy
iRSnFQnSyWaRSl2iZ0tA9Pg93B65FCnDwVnuxYm/KZmpIrPZWxGpW9PUe1q5VbfEt5zovvXey9zg
y/fbwllP7vXmsTI1VPE2D+YQXg83OYhCYql9WEqF3tOPRiveISmm+y4WIn+G0aNRl+hD9EwEE8o2
8lbamlcfF8QH7e6enKKctZZjZFoVbUFYUUdFxANfONYDpOF20SodmgzYiLJGDGILcY0vKrWVK0VP
p1tMglFBE2PcruYEmen9GZVeYvr78NMSQN0v8WJoB6eSi6xBSYhmD3D3S+VTBr7NxkFnEw5d2bnL
KIKSW2WoCzTZzlgah5+jzh4xfTWXkOPlcSzEtNLhFS/RzG9RTE8cxnFVczf4ObvKdLRpc7Xskt25
OMbshvC6NyDk+XBl3z9+hDn+UGCQNaGjLVbuXP/9RmVkYeC8nu04XqBB113mkp3TYsvQbyZUkExM
jeDUhBRqhndIEAXd1jnfkeNmHCm1488m/hfXaK6W/3ARWdYYnVyafATYQX1A3sHDXVsAE1FszyeL
MhUglcjIsnKyDgixX9f1EYdcSLNI4s16+shlrXqcozKsc/D3/PkzBwxcYcYWRWmySEkH1KNn1MLW
5FbhMH5U+htmpUKHGDxSU+FR6lPotIeUY5rxQLV+T3DPZhDJozjtiH05PPS8J4RQAnatlffDZkmO
M5RUOf7/3mZvL+Sjsu+T0Q3H0Stom2Z0AMWbHB6q+0U48pnkQvCZLIrbHd+Wb0hRyo9tJcmuiqOH
Hmk0JugiI/7AjPBq+vs/L1xM7vXF5F/9e2MTYn9/Hk2Dep6qFkXI0p33ghkNvY+bUlvENel9bOJt
h5m9XM/2yj/ho6FsEOVfTxpWCSrhBWlDvI2NlYK2J7yZDDxaA2LUopm3fmsu0nflBaE62rQdNrag
VOKAuUv90pjZWAUCL1EggFLJOsWt7XOtFzeBaGMfzZq8yGRnEBmhAB5Rg0WuLl4XogJSJ6j3mJ5W
jQ6A8TAHM8oGmVPX2HNpnbQXG55D1vuQpYCGS8dSIlTi02HXHO9LhpN7gj4+BDgWvDdROTQNCvyV
I6CTUGMCpRk43PT3UOfDxkLU3BkXxRDiIvqJlnchXZPG6MQenPlN/G3Ce5vb/rwAJZWzOI7uoZCH
0KoorW542mhHcpIO78Xp496PlMNoL4EhfYBYqKQeSX7EJV7/95NDg+0nL50ixKqpvMa5h1QMOWa3
72dEQatb+SnXr1fvg/CqANFxuvcdrWzZoNZtGWKrPZ8F0H/d405XMpAg+wTRGtLcxEJs/EzyVn52
avIugjB5OpuVrtHX1zOHhZDVbhn4VQ0WienDdq8PFo+dwMXclkDFubssk9iuUSLvd/MFcYlFG9W0
P4ts+2GbvPlXkCZV8Jp80WDpyq6b6tPwe8q2OjllGYFUzcESFm7Kgu02qazvwPXfbTJpdXcx2Gkj
Muo84Id5aPC2ID4694JzUc0Rlzkx7YU5/9wIP9HNCar5mdQMTi9jI1vznP4TTbbwLJsMf55XknwM
5CYGtnBDDno4pH2WZgmKd8np51WgLzJ5GPKQ/XQfcjQZ52NceFCRXpMri9LT2xR9FYAmYeBKvsWm
vALTW89iQg9dDUVRdG7XAgXfKVq0FQ+KblC8VnpFjMdIxrSVt3yH4ZQ9JPdWyAcSYIAAesvcLlya
fIYzPc59V+txxJTZ41n2/jTipoJ+biCROfMLsHQU0cMdxkKobwxl5BB20ffiFwvdqQ2WUww9dykY
gXOpWvqPDMO1LQ5qNYX4TtTsj5AGGmtcXRb2o+wS+7XMr7ZT7x+5ydqa2wiPdpg2qi4imLlY7XTJ
uF3F2e/fG3+dswHJESPQveCf/tiihMNlB9YSGjYZBmtN8jTs0H7YDEHfuHIkRqrHlst8mO1Xg8ZN
5P5fqA05ivcs7yKVwhWEl2rZnphkkmSfg8KLWhnmPMI/alUdm3BrWlYyrXnFBE7w6OAYIuIiQhG4
idBrCBzC7fcnX4im3iNzL7y6akoDH4fK5dPpN66ufWuJAwjiPdxq5w6udnEXKbyfli/ahSxi41hz
a/x8r08S+vvHilm6FmyLLbCywEnDPrabGr+0MbTBVl8fZulazsLzNpvlFGVPx2nufuXQF5M4toAY
6ZIcEW4T26wD7b5pkqPrRtwOrBD6sD/yK8Nby0uqw4KVWjXma6GMpx4ARTmdrs+KdQq3S2ExxFq2
JI/FJVfaBqX2Dd4SiIY+ysjMR8/raaoHTzVs5x3vK/Ee0ViZkQzIBbf3aNGgMmE2wrXFG5CaLW+3
sRLae5bOVLlY90fS+qLcTaQ37afMv4W0JoMrMOvCROk64UNhtkxLMp4PN2Qy+vkZVpWIe03T0pLW
2vzCx2jlJm6uvFOHHm3AVSC3qrv5ds7r5A7e39XLbOdTxG5aZrjsP+aWEcFeV8tC2Moje5HFXjQo
CTQLSJMRWCCrGhwYnC63YGHziJhnxarwMNPezYKjuqXeG5SpfDNH7l0lCsU4EFcLC9l+qkzV5aq2
dlUtRoofWlYbHBtbOb/gmblQmQYWGJZ6/sLKLpj9bw0T72XW3crrify1rITDbhn6VFNdkNbPFQw+
mb7sKvjNzefHW1UOCIT0/YhOBc20e5Cwdl06mOeaJjMKjzFQ9BbhwXr2dqlcv4NcPcvJ4k0v8EOR
BFEbj/k+TAMc76Izr37PrNrsA7odJtm6Axx9tvLyreaKRWdVh2BHBPaaqEy9pJTzykJ5mkx9nZof
7EBliSmPLL+soI1/Hu+PA9lp84HBrvtTnDrogQQC3lQOQZmKbhT13RUgHfYpcxB2SNEpGmkxML1q
MH2qajXjxceW54/ie2BPs6qepzhfjM7j62AguqmlobhVGbunfnsTTA/vhIOKbRykmSk4WZa19TmD
B4HPJOgNjNqXjfYerXu805v43bkTFA00tigI9zC6QzrqPL5jKfBcd0aexhenAHlo3JmHjwy6BZ7G
aNhCQe9n3A7ihAt81i6t8ZdJMEt0+NKDPy3KHNCQB88rQ9oFiAUgXUN+XE8a6UDJ0lIff+HdC2AY
VOAtxKPb5tSk8TLyyVG95HYDB5hd1DWHN0kPW7VP9LkNS1+cNq7ObcFJKgIi60ipROu6Bu3ZUr4o
w9jLMNscG5guQqfczIZFlmdRZdw16WSmNW9fcz8PohpUELrqbqr7214h4PjBtpX1VshkMTWaDohf
1CugWpVimjXHGZG95Hr9ki8YFoX4CZA+MhqbLKP6cPobhd/mjs7hYzTRcewtoZaLO+E/8oj4xtcH
qiRJlnFdQxLaZARNZ/f8Pkv2LMWgBS2OIqlP1WTr4BGOvOMUwwIFzDsNtyqD9Q4p537aLzeR4s1j
2D0zqBRnU4eTGDh3Poniq43u+rskoOPR9NZ7eWVwNAz24anlR5foKB23r/9YMnc/irrW/YqaKklj
kdxy/a3kLyG6soCYbjF1O0s15pcemhD7H1NcMCDmhg6JYS91m/Gqq3OK4Q64bqMuYY6wlZsboNac
3xHc66xWXd30uKVVe2mX8uBNTyfDeSVXpCQQ7EgIs0tZpnCK3QDMNMQi4DrjRuaFahFgv8DawZF8
kEm/Onw8emWppAbGFraH4B2sqkS+ZDoxMJAGVMzAaYu93UgK/8Q7aUDSmuWKC3ZnUySSyaTTzuWa
o5jQBb4ahJOoUnFWRMG/pbK7KY5WXW7fYjKch9nbLeS6lAeTP5eYnC0aG/Gn9OtKR7D8NFXBmoMA
67fpu4CySfZD66ev+EUtc2GOLUERRbXUjNqh5SOVOhsQbtnaNgtXXbQeD0JKzBIW1463cODksSn9
X4u6yBElsHbZjxHz3xzMbezvYRfF7p7v+pOTsglFdpvNLTBqbUlDvWqWAleHPdeDmXIAcTO/MX/V
qyZJCxhA2nn3DzvVMf11yZkBkY1IL0JohGNOf6MaM3KLtUGEbEHGtbniIGdU7DdF15HCEyiE+3pW
85DPgc1t7XwPZhSxvz282SNHnZgUrSp6AUJUOL+cOYTnbXGSgSbpVSCjQBWYeJLspFB6PaBTihb6
ixjvrHHviIE2KNPvkyn8C5g4HmsPIvhYuHPg3BhzVNYXXWvQuxkWvC9igh2n+ut7t3NJQK60Q6Q6
cQQR9UYMOnlXDX8L/2BRUBly78AIwvScYq5rhX1VPWEOlDjs+Uh4cy11pv33fNP/19hdn7Ep5Dlr
KJIFeSVFY6aNhYky253MFR9dxYBB7FmU0f+EddYBHWjsJJlDU/e0we4luRdoVUr9QuMj0yL4LaBj
sdys9xf8DZCa2e58DtnmMcn80vvUJe+JbPZOFKB3tV8mypk4K1mt1RY3eq5F+6R5neTG/EvOnH8E
84QZBr5/5f53BvaxENKTt4nsq5zBevmmhXz2ekxygZQV789mNjuBwBk7wyXSWAzjGO1z6noi7SsZ
SOdWksACpdIhcnjSFIiLxG6Dcss369Kc8UJ5bIVFsGwz3JhIbXkddk+h3hrzWowG76/w8g46ZKAa
XxBCAbTjTt/Lo2wNZufXl9yRIEkwFfJCS68onW5rP8DjpTqHGe1PLoJp5t2sivg2zhVSYkLqQNip
ts7QQWYuWOzab+ovLpV07MchYcIIdn0Ieix75gZR23DFyXeDDoyYH7lNfItCYLkP/AaYd93Xhnia
t/bm/kNITNeirFYn3qls6Og2Cha+NgWH1rrnqmj331DuHmykS5ASSojUG3Jeb5SLSoEh0vsUbwnQ
MJOK2iLinIVjJiSbAluvHIJZOQwP9bGvpbfHPyyYb5idGR1QoPcdMRIX/VO/r1gu1vQwg4RJp64p
94pQWXB+U4+GXERDEzHyg1UKbN3z5ZWHs/YmB77pnXd5PXEZQvYfduRQcMo3A9LB+kHQXMkcK+n/
Dd9VxL15qK2aRe0Yz3M8Uegj7VssEx8blGtAa456SLHHf9Na+NcY1ttl0ehY10lOXbzwgIwAFBp7
JIsjWhV7vPYsp2OjeWbtf9La0dbEu0GrN74j9gXN4AW5MF5D5a9fJ/+5m3Rt0rypNGB3NjRjmkea
Kykh0PTcsOJAkGjNCKkK8+Lbw7AcHOJAIjm/MvZaiF6JFz/bHj5fMcgRPkJOIIvcJZQpKOIK4ScR
W2g0KLxHDIQA6AMUOUMMdWuPol8u+CAbfc2TMsLTN8jQCrIPIZFYnPDly6IkKDQo42sf7Ic4B45x
w6pfWB1WX8BHfa73fLEhSXi/+a22th22jgKehe1dpUo1njmesBO1EzE5DNk9v0mPPCJzByjH94Sg
zGjCOCFzaTkAid8LBPgeizEEmVuWDpEaJJmO73nyzwjC+l57RCUCLZ03IzDDxRI122sMdtc0ekUj
v4cvK8Ln9utXTnkYkHb7YC1tkevCgORQcukT09zA3enlb+lf8ximSkSwX9rsi4h04ycZYZBhYIfj
V8dMHl246xTyxe9BvtZrvbtVbLO/li0fqCQlWpf2RLQYAbHdT3WV4+4bZcD245LH4jmoI8SbqCST
+zzJJZGNNUwgC7EiT7EVq1rZ4SgmOMNC0Thx9oZEI+Uos82d1a9BBz41+NM2gAIqL9AQEy/2y67e
AKWthed+BUl5CjO9u6zwsECQdpVNQW8i7fxELkSsMQIn4HgbGVwl5rWvYGYS4HZCFZtOJzgL28KO
vsDYvF2Ac//bOU3H7nmhg2HID5FUVx8xzhuVMSp7GEb6/w90Ih6S4DqOCYhX/KzVRkozKCtcJylL
f9uP0S2Qe7kQknCys4d8/74MaMG8w/Jk4UOJR23V2/dZHjpwWK+9DYwbI6lKGEhHFo1LpFWBhkNj
rFSCOYU0tANPFsqD5a9aX3sYX0SvcNHlVB5TfdE0xF4e6vFHCZElAMsx/xGrYwefaPTnnFgz2tVf
O38mqzZLP33UaGHMcZxZP0VDa+xqUhA3kgbaWtvVzqXl3D23T7k0SUifAJTraoh65R/DypTjrxQ6
MOdg9c1K4qebxEctrpiRok/why005myIRnbgfzraAiiirq8uREJGbYPw85OkzsEcOyCAqZ+e26pT
ki6dURO0X47fDla+QjkFbvyYRChlhUFTWlzYicwWXqCKRJiodSpceRgb5YKnhTWK199L3pKkzFuw
uKW46u0+tSE7Mjk3OVcUeDl1qrAMALo6vTlReUBBMsokbYohwOkEh4iKO5xqX25bGqnhMa1VJB/w
0oVCVnVy5FtSUd53+1zkI3JAzFjsgW5hMGbxA9esDeCyGHZ8pPjOW1WbEAWe/FD8LegfpaCVL98I
n4byc+QoSGeEgYicIZuvr9e/p4bKcdDE3Sh77LmbdHQriopuB9yqcqN2mADvFjaSQHKRAgTEOvqJ
T/Drz8BSP/ZBQ+bC1xXM9gyXe2xl4aqXfHfE8/jtF6Ol6q+PdQoKd89v/EGJJLQGIU+QjIBUxjmb
eh2XQFUoPgJFZ9/5pOK+8FyNjR1SN9LmBGJX47A/5NIflI065jYwjlnj2bhzeKQ8Yepx890EIOoc
og0y3eXFesVHZy+xqkp50kU3uzjGSdwgHU56EX6uacy7vWAefl4hEi53IyDXT3/dOGa5b29zLag+
L4qLhz1zfu6UTlo6C1BeJ5otNvN+LENDiZUdf2hmMfDeaJQOXzE6vb0CLiIdUfIWODG9LLnn86Jx
Ym4YwsCFkJc3T51wgL6ZDXgKL1a2SnIejnpZVq29TR/EdZSvxVzTupEcn2hUFOQ/EC9t9Mg6oxzn
5UdiMhjdibD/pckp+Yzp8g/8i4BGRbGbPNB38oVWboWeqXJWXSWmso6zKbFiYOrqDJGDkvx3ScHn
GsVuVuLHmLIHllteuU4QAVdSrjc/2F8i0veiuecUdfo87NLbyzdjUuhHFGY8i9pvKgT0WD2jTKlo
uMKIEU8bzUEYqZ/lhQOE1vGtpXxKdl0LaWqPvwxrjkUT+d0qIsLPOESuRWFV9cwMAMbyWa6hjVpM
NR9oOO+etDAx+AeJ1IHoz9vrAF2r2sZ1hp7rK2iB3hb18W28rNvQ4/Pu/++cHGY3CulyhYPeJOdR
zAIlPamLnJ3fs8+28M+FDsUSsVfqaoAnIu+hYZmOeeh15rtibMua7M/VGZaJjHkRYR8kWm4vQDkL
KrarZjGV276qtA3InLa4eHkncrLJlv/S85A34KZyBx/6SPtSSsAnvZoMLv45fsuU7wGY0n9aTGSW
cp1wJmdUBfnzRsJkzbKb0by9xG0T5mHYcJ7rXeoGMvfzkzgtG/1lwVpkF7iiJP3h+lnFX/WpxfO1
Ist8X7aKC2RiAa59Ov/bRSHMhS6qV65o5rGL2ZhHpoltwBwmIAWjm1BR8RrIFakN+sUPnoOKEs73
K0O1hP6XuLUhKu+bqWhFocIqNv9Nfo5BDzJJV8N1KO23jzyBHPVCGToLa8CMDUqlX7mGXFg94yec
z/hjijJ7fRIMo8VCV2DYsBGzhWm9rVpWbRxy9RBsHws2H7JnFu9VKODwGK4CZG99sgdCr1Cre5D2
ProOazGohQEO39AlVNpKkOYlPY9AgdLS84HvruC5NXXZzWujWg/UjbKhKYwmR0vuAyX17RfGWmGn
mfkX9q1VaGt9rLMTgPV2onzeCJUc+V4NTFIMJFA/m2wP9wHMpFpTrvaPC/U4Ef2IzF3J8SP9hZzo
WQJ5cTOZxjzXnWEk+SZCoLTSyaEoNLj5H280ojyy2Y7wTgMZeeAibrSQUG99xsNjJYCpjj/PwBIN
VjhzO6il49kB6yyrmJF2bKQyeEQ7R+oc9BXa4hi8c+KPeGNuD6yJBEt1U5WFbVjwLwEOkqu/EAHj
Zli+AGnMruEaF3Eit11jOLXcmG2d9h307HEd6Yp40YEp73ewUHZN7CoKfAXRMbltFJVW6W5IuowD
Ov9EcVXFLyhH9VrTOyAW7fL/YELx+YtsxApuDccDIO9wqgoMWHRNppgFyLmst22cqwLTpbgZP6qa
pZrqGmWrqn0mkfw3ejoTv/CSG/O0zChd4POo2ddI6IodqWGtmBWAkS/dTLZSviPLZi6UiH7xzM7t
grHt4EV9cYzprP+7UGHL+Z5alo30xhFJK8Umh8qEJhqULcYWGzDq5eLoMnwMy0egPUybsRPF6ef2
0Ownz+bdNJXHS0pKN4TuxUftTDqb11ZFqXkAPPY8O9M9H058ICaEj52hrSW2IHW/pADUTqxRX2QS
7R5M5yyc7QfbwSQ7CoG+tzy2X3Dmca8A3Rxxj1/saMGjOhWtgG18KJaRgRS71e40soMstuNh05xA
2Pv71QKEJ2CfyHr5CXAvm2yk561hw49gzsl8FQZ1oy7vvJxGENDEqLWtLEnpA8TR33lGm3YajgMR
RQUXGZDyA+eI+HF2EkjlVFks/Mo538C4TlqxMh6l7U0vxo+E4zx4qzlnhXRDFGnMiaNSLVLhHrKA
poG8LgjXLi9Cc2b0TLBCbfyJC/EEENq6l90/VlnI1wKUQ5XqbM8y6XBhmUgwvHHSoG6hwux6mDqz
lc+t0Ec8hqSGk+StodzLw6LzaZydMwiPwn66yy2ZrSYqXus4N+84UfbheWkB2Qp9iL505+ZHnvrT
kc9qY5DCmlDZjS4ChbPLpZqjeFIxcShUSNy96l8dmEgePWA2fOP0AaW4CB20piy2g0EH0YjQVvK+
6zMpSgdECWmUV5FIiEvHBJa837P90JSFMcNHLxQHP7qNHzN/nkFCP80/pmXViOUO2cbI8IZBMs2o
useGLLnokzHmXGbOjSFy+jO8+mtV9EB7CUWvOmPwbEgaf/3Wt+qb8oRiC4FPNgOi4G36TNT/2s1J
7tNz2EFVM38WaMtX/N2NEyzVRO8wpAT+u5v8xqkamJ8hEkzsMFz0TYBDauZMW1mkMzof/PUuAQRf
hOcdo1ZlfAJyr2IL2x6+4n7Yjk28aM/7vBiTJ/MDpnAnLs+4vzlnDS0a5Xbl+ZJKwf5vCtdZ3Thj
VMHqcKjeiqWfkJbp6QQW7z3eS3OBue3ux2kpdAdCSHjbiziAoduXdOGjjIaeeGKLgtW551RGS35T
/QIQdDmHfsgbAmLlzBF1+CwnFiMiKDlIsT5/OUjfYc27xsClE5VNLOH6nRU935rhuX0EWNrajKaZ
bGb1BnCTmGc2ovZapPMxdHV9DNAnahWVK0NsZE66Dyw9Zd/Cppg+vgGja6hdRD8/efLVsXkp33gM
q2e7tde0bjog+ZTh8EWZ4DnpJofb21WeUPjzRvmih+MmYfgZYhZjAAABy5Nm4CFfDtE5R7BvqXnP
eMUe8EavoqIc1/4YMBsu3atb700SztbUOrGwfsPrNB82Po0Xvet91fK863tVusbS9FfSTn4pOeNu
aACcrUmfCDf9ZaRR/l6Iw8PqL5KKncAnscqh/5kTX7dfLXdSr61icf5wpmGHO0Sr2Qque++iNdXg
uXux63TX+JUv193KB4aj0WhDHPrRHVYyMRUZ64lds41cPdGq6ESZfsOk/6C+KrstLMijwz/Dlbp/
eNbdscQiqY6FpygmSvX93TXrzTg6RjWPYgci2bTVASzmv07xbhx8v6i61QZq1ASgGdrniSabkAl+
UpHVp+/ylUjlLqGR0GfJiofQmj5BASkRQ/+wu2TirM0ysCEM0eNN9PZ7e0UQ/xKbScpSS3wpe3a5
ZKo0vlyh1MIc8PDcc+vyYvCRsdnU7RkHct9LsKmH3Q9bhElC3ZTD8pDk333CwxdK5KYWMXMmYlvQ
RJ1lgDJnGPIzwIisgLhKh+h7z5/09VUMFsrRUySK0qUUQrWcyVxC2L4gJBtV6YkSv8ykixw1FHBB
EA6VHN5iseQXESLNQrP01hbEuF731cnlGmKJiM5feNfycGb+0EKPT8KCLd2d1edngp7nE2lsKTCQ
7V27+QEiYJHUkUOJdI8djXB54Ng2KZjvU7ixd2aFgLsMGNvi7EPddQVneGvnvpqjubUfeVNHDu/X
Tt365I2r0+VqgjbkAXDYzm5YHjPgBgFocB66aFtTYjy7Pn+Rf3K69AEzjURpekTQzJd3qs/QYzX4
XsZB8rL4v+hBXAxVeFL1wPbGpEt2c23fmaVVbNuKJa9PVI8yiM2CRO+RJXzg3zTVxg/NUb/tkUik
My1d4+lCeGKfdtJzuRvgEiugcJi6Jx3Qoy9H7k6gOKoHySVWKhb0ksj7uQ3IFPgAVa/Ms9JJXYMy
Bjyz0jpBCyjKFMchRHLkcfta61syyUg9LkbjxejDD4Ms/J6WhOlsfFbrXRqTiXZ5Wc8kQIVHZ9Qo
rCOimfVdpErDrV/Lc//mcHRHYSAtVpt0smR7h/5+8a7SfYsMTFbM2BxqKxlOkPixIrI7+d6SuJ7G
uDoJoG4MEMFQ0ZSNpcEH3WJN1wmtD+ARJoGeUKO69xuaq5F4daSuIjrOXjyLq3/Hl3qLuFxKK4eG
my/8YfFeWBiy1JCiZE0iETFBzD4/1cw9iTjBXZnogu9CFNSc60BrXPLDAfI6U1xHA2hay0EFponB
rQ4BiDtn8bxxLou9aHqV45LGiKH13Y13Ki2vK00+r/zT6mIpaoBV8FH53QGqHkV8ymknOk8VTVho
yJ6w3C8QZFI8EEqo3UQMAnn+JuQ0pzESjFQ9hRA5corF1Pp0hLb/zVEKP9bJ6APZyYAywj+697a5
3XvdJ1QXkHgXqWrAo2GscMoy55aLFgzmVliXIwLG1YG0WnNHEYh7Jnm81eMxZHTuQUKxwELkd85c
elWtTi0D8tFPh8lO0zKGvMO1XHghUL2/RgvtIei3UafdFXSS2CQuhbG6GxCxHHY5aUeNBH6DudN0
9uutMLZ+lyNs3xXwAl0VIEU8+DdS5IgFN9byYoyVSW5QtIkmpPQICS2Xd75hVvGktxUuaWuG0qYf
3/z3fA8KYQeGtw9xfOXQO9dMcei3OyBPhmLd75dIbSDTCXnudF+yqrthfToxNWQ9ysfgQXR/rYP7
axULfkA/yQB7Bnxn7M6HpCCypRwVNWqjir3tqfHnVy0yjaL4cg1oK5zEG0YndnZB4mB5pg6KxDWH
zaEcZnui89yEIgkPTwc1T0SZ+7Q8scBLyj/DGRZVwecu3pXk3NK78N8XS9cOTXANZUK+1QGI4trt
gUlktLb7bGlkRm/+zrCN1slQRFYPoCa9a05nQfG647l1D37LU/8cEkiwBBKKG+kHBJHHji5Zt2T8
Zv1uv+/8gIt5QpXiwpZh+k4BmV0Z1YkibtLO1ZmQECEcN1Vh/y8yC8sjUMI2mg0lOkuPTrsc1fW/
amM1z49F6yo0Z89+t3M2nnbNQFBwFGpgy40CcFkJTiEOHqZwE/f87AlTDn4rkV7SyhwDpPXCSsD4
11S7sIrjLsuG/nLDBiLKyIYS1OB0aSJytYJDK5Cp6btFDCZK0hU2WLoq7hT8e8dtSHZM8WCn6An1
aHVYN0lEF5EBUZ2mPs6RXj2QM9RikQq/fdv8xHrTh4MIhMVZRAAD2Yasa5xr9szoSBGCUBsYLYuQ
WdzcbN8kFrPp88D6DYsHjgZTpDqzxgpfEOn/SDKItivGi3M4ibEPKPGq68VonluMXl6MSt/l31Bc
Wqaozt7bXWUsEXoujEYFAZn0ZG7xKP3cVaDKt9lL0MRwDatuANPTqE6KahwQQk+ld/lvRlidO7UN
GAMudiUDzAu/9Wy/0y1DhkuN3ltNVzySUXu70N3znW4/vVaO9wiU07AHy9LC0cJZRJsCSCE9z6q0
Ju21nPkNnia1CYqYdt92AgeUZvhAX49hE6fEym6pTEkw1Yw+SOqTEHI1SFEOOci2qm10ZZTn1FZ4
l1YHiHNV4rrCWqc7zvs05hnwuQdOmB1rHSjmWfYZTDoys5Mrhq/iVPpu57TgJxxMRpCbkz9dijgR
nYU1bpjpvnExVXTX4qIe1pKNHy+u6Y3TmxDB/aUy81bKWGF5MyPU/RG/EFCJscOM1nkpMWDrx6qZ
MoJkQXc0uQGV6It3VE1wDbp0YLsYvQnvkU2SM17XZcMJ4pdNGtwtFbqDxAYp3glCWo2LhD1HrZlq
fowbbbapIOeI7nBoDmGXA9xawj1H70+D5z2LP6gRIQDC3TLovWKr4yT7n/s6pbpQfDqwjTtiXGb0
7TQdfFodQtHs08QiMcxsQX+ieORTspR1iTXDaRPbZCPWzIEPBmG92iO5UhSZgcuxCbdcisHZxJIw
INq0gMxr/tT+lfb2l+P60Y2z2Pk9lOJkvr3FE7bYO5EW2W/A1OcBpEcaMp3bBo27WRJxzu+1A8HA
sg6Ic41jMo4kbxE0bfsPpKDxkhwnJIei5XcdjuvNf8wcMt0HrTx2MxKRsPsECo4UnjdqNz4bEjsl
GPsqP+3NDx6zz9XPmu4Pf4h3iMe3+Ot1rOl6lX/keboz3jV0dG0jdFmdjjdT0p1a3U28zmTGcx+i
a/o+6R7i7W/0x86am0uFkMj5X76ZlEGMoK4JKP6x55ZcBahMLfzHz/Wuk13/41Sc6t8b3ky9/NAW
E/E27xIgMhV924qyqCqCXPcYmjwTjfxp2s5bseU8vV8KRMJi7O5FScN/pzd2AcgLquhT2ElUlI7I
+nXnMC8/kPAtcPY5oCEjgZZz4yOXIOdTjS32p+loWkZXlRUuQTJLUoFJ8Os/1Hfp6bo4iQkb6sQY
DmIwMWQkRK6PAOcBJub3rqmtqmloNxXK+IG5MFPCq0vavq0WmHZB2vJ6IS2+Vb3opZGjuo0pUaZ0
UL8c8TBcvSye5a44Yb7HQm5S1gKms5rqellbgAsDrKTfqKuWxC+/EVQe5rxro4oP4DCx0IlDnVtq
KIGRTmFXpEMzbDVJcp1DV3GMKUbpq+YHIsFayk5UbAtewhdocnDuIoyyrQlFQtfs5QpaR3ODwiEh
/TycE3iFAruOlTPPl2PjdWVKu2oFQJ3sQQBErkhYQAaUFCkKdZJFm7KTXOQo2K0bGd8ZRtxtMQOF
Cd0T2XDTy8XFUp0XfPaOAMAFfS3p/Gvi4s76QPIBGbSsDnBv7ysxYYEpDpU75E0idazJE6+LnowA
gydlkWt2VhjBHo5avpdAYClIBM2hL3rlDoOSxk9WJKPkc9yEVdFNJfwwOVaKLpe38M87+wBJwv3r
wUeuY0owGDiWRkhrK4INxiuymruc1K3JZe8IKD6vZh7tjDwONujs6fYxGr+ekw4BUo0AS/SyJVBX
HcYcsEdiSw/xLsusB85asUPmF7Y+69mSuH/3uwXMHXQHGox2Ugr2q55dcCZEFvVlnRwIJ18XGsqA
9jnv2YmkFGcdLXj4d3J1KTq0o636EXATqCYwnDklCeIRDxGSNmZhKwxAOePyfIXzsR0YnCgflD46
ql5yDGHFZ6Ojs2FBYD1JJMXjyldEPxPT1CMpZydiFsXnsTOIbEjBV+/hKIYsQnNdcj986Tt35XWz
vhjEg3RflrOphNcVk13uraLrznPrFpTHESIUqSBkuNNlb1JW55QLb1H1A9+FsoUHGBD5hrJTWv0P
ae3M0Hh+6mf7DdTcm3Ti2Q/N8PC1JM5ses5Zz4tLSA8qEchuMW8v9iOz7UbOXDa78PX8MFf+hAuN
IDSZKGvdtZpRwkU874Of0F50gebf2iW6d5Ily3uxsIcBxnGzILWtR6Q7s+fmpJFqLMG3XKToALkt
Rm3jz/Rh8cXLizjMV8nDeKn+EFEbzrLN4j26MqQi0lC0odANY5VFj+Qw8tF+mpBie2Q1kD5LCCkd
q+wXPswoBZbw3chc3Jsp4BWQdZ1Xcb/boTiE8+YVxsmTINUC4Vrgh7+8YtA5XaWDFP0IMhmaa8Ji
Utdgz3MhfQHuru/FDCYgf014i9pUSaQMImfdk0AH/3iY5GDh/QdroR3yf8/pc8A7NjOiXVZ3DG12
etq8YNPCgSycTbcoaLBaJEqEyQCCmvSWyaClAbNt4DBoASWlYWBE+/S+UjidQEFhpaWIgipmvnhS
JIIfVcB1mX37fCgRFPC5YjhMXY6LVv9/3XxWwOdfq+Vcs5pLp4ZM7ecPlyWOG7dz0+wzBxg+dDN2
s+Cs16se6yLVhABIcaR6c/SHyMTZkQDfAyY9e6pFPbwn8vz1du9hx3mPRegb2X8Vtm8kP45VxE6O
IdYv6TDvsreQbTbBVnbudeR56lSUG+mqf0qmS6wthsQVdhKsCgKjbgK66Ay63fi2oujwVVxBWLv+
YcGeTk05qP9nv8ilICXD+BNXp3lZ2kadFj1jPD7s/faXG4mQpwLgJmojXwBeD+5CAIgLb1m95+4o
Surnxipg0GKWncLL63Ms+YgQVbOQ2efBjcCziI0bTbTYq/jIZO+Ifsj8944pQzXV5iSCrbkS1cen
TP2mOQZuvyqhhJvYOZy47nm4aOwx4HR84a81cxwFmK0h+T9VgX9cwksyAXEdY/ikCV2eJt3d7OcF
d4M/ed4rof1TTgjwbCe2D1/a1RYnFqLB4oncShXCCUSNRqkbhrbhaDsJ+ukVJu/9ZvSs0AqUQW+p
5koV64xiw+5k90zHp6GNsJVbGQICO5IuM7eOdY4bHaEvCStTm7gXvMkJxC+PNZ0blXQUwnIsrSpM
cymVmZXfCnGHSu49Y/ih3L6ndrWH9u0w8dqEIoVkmXhOquw2H2Fwey8AsR8LYMrdAzQCTxv1KO8A
8H4Qt0EWkN0cXLmOA5H2WypUBSSpXMZsiwBtDIP8e5zucCr22rGVrVPL+lgwztMBTk8idfRVS7B2
fgV3Jy9Swtm2RIohd+CUMldeCf0Lh1dU9ifvxeyPhBqXIs0q2FAIdOA+mDRqeAERdrxQBHeqknw/
uivHvK1bb+TzflU221xoTRPDhvOL70vTpFF+/o95aeNPO5vPX7N2wuTUNbPJ6rVvhgL1lADviViH
Xh69aB1N9lAcVtV3ZjgNTogRSQEEUD5yh8DzLaKKX/gXtbRcWrTMyQqiJQ6jlnwO7hwUOfWcKXED
n9twPvV9nHDWIWL8K0iEPOHiceWNUzamGj9F/vaUFkK5cLPRf5Q9IVlCOAff1k2rsNh1pFN+rlN6
7PpmkUpOVGEznmqETJSogjPl0CkJjDS/W/Y0rQSJfr8MRuTeRfZW+3rEo/Y0FJd/JdP7vkzbcu9S
FljyYJEpnr/t5u1kilCa92iAxWSLmOgp1qarCP1Dk9pFawnhDxExycsj2/kuNFlnJqs6DMP9KE9B
pJQYVM6fYXx9OL+mGbk9zq77+6ubrty7Z9nbqYoQlJsoTSl0t9dPZ6z1oOxjvh4xFox8t1XIvEB3
IH8nSH7gZwpsB6+Q+Y4HBx25WN05V7vxBLxiR0rOOwGkfLp6vs1/s6H6sVkuSJVx7dHlpf8Lc9Vy
6P/lRZ3tTlNbErNE+RfJCcdU2BW/G4yk2LAhSCbgx9ydoONL2zOqL8/x0ud935ZHt84MBNo87mH9
KUNuv2QmvEmA5AQVOdwmcX8UNd0gMvfKtL2l83MWCrdfQh+9hQjDNwKClsuAshVeXGRQvy9IwiNf
IHNKZYArbD3JBbTkciT/AxMkf2pZ3qu943nWURwVp2e1Lhv5Pr4QyrOOw81Nb858nHqzFD16tL09
oYZmripyzaehcMSMShbjEAynT5X4WsI9kRO4mPLVDiH0ZZLZMaPH+lbZzcYy1yUBj5T0dJ3f0uIp
y2z9oKuBTrojUFRIx9ZKvZmxRNRNXoadCED2tQQLFljeT9exmyf6aYQjhh89LA/INPJ3lIJE43Ga
jfRshIXGrgpOHfooxARFA0OQxJV6yovDmFzF7MDHnT5aguB13rKFfPO4UuNlBH4hvOTe/zX2NzAT
3b5BEiBhK7oFApnoNh0bKdbHVdq5ViOwOmzexYm2CQbgG37bcqrJz8By/GA3VTCIkmVfTOBCacue
Yd5ezEmOiVKZnQqcn5vHFK4bp+3Qyqy7o05tML0LH1kvJwWKlDFBqB4YXB9ZjY8/lPzg0V3ejhDn
DEAgg/zHH+yMIxLfRHBvaOg9Rd8fw6fl7zauhKRl7zXv9erXeqN+5EOyNKfc0JRLNHN7yGsvSKOE
+cp48vSyAWOXCUKFY8oj1j8+bsnptn+YAuL3ivVM9pfGCkYVJSefeF3ippGQsHrRzivtnWqxQrmR
4Mo46rxAiT/ANs3n2NwJRTkjTqEu1hshUE0nxvxvqnWqL8/7cw9abZHS+0WNQJYpWk3w6Db4H38S
zCQQBxH1LZNOcIo8e9+MP8gItbAcgKVnX2Nbh4uXNFsRvPfoOAgxC7mNAh4bvJYDx4jJQQD/qfLZ
Zq9GGxqVFGXlDegjgL1kxYGfSf+uqJjVYNnpzbkYWNbmwMIYjI6o1P5oPUlUvR8XGijrm/XNQLYo
Or8SyckKhkrB//iJz9Kz/cnMaU1EzYhfDmBDvQaApEC7IuZRczIw0GMbSHdvu4LJ3YP51tpiCb8T
gjHAqokszBPu0v9V0PIFaubGuYD9oIlDAbk/i+orA8G9nQCJnQIOglaN1Eym4CTPE1oHYTn2F+Vh
MrHJ8Juw46z5wXRD2tLsZsy+lKEGUCNOeXXCZczU4obA2NtLwhRMCk4a6/as8FGETfgfb/1k0ZHX
IlISR7Qrzb3xIq3+JyZjtTGHOQ+uMOb9pBoIQ3y5Ydh5cc864xeNRkKQXvnxkMeWGm+M9xPTVlaC
/FUG2TYuCB5FJ3p+edYf2LMHwnDucjAfz0LP5kLVbonVpSCR6PfZpfighptLVqpCGW5YpY4jtTJ0
Ix4wTdXs0n4KRFhaVxCradrLbmGYBt54gE+0OBLENu5lIbrzaOgWC+NbYFWlqkxBod7Y50bk9nAR
3NCFb0TWCvCXzQqPStUIRanrBKAfNvhg7UN+gRSjJkvgkCD7tRFNFLkt17JDqjEQFe1bQEXVO912
+A56W/ls9jKpoy/tmWJz6O8FuNlnVvlulwjJ9N/MEm721sdIWHK4UAqSR2ZpyFZYGD+pojrVbzgN
0eE4fVF/Y+ij/DGgMBCYSLyWmUN5469boj/LSn0jeoQM7+TH4K8pwVagnbeJ67ajGdYDYEibJ6Jv
tLelmP+yVoxMDXK5vVgBuVRgXlVy3UPGb74rH+g4QytIIgrlmRhzlvBJpsMBhpdgmMDGkBoBR27g
vpV1xTbo+u9Td4XJLFotsmHxxzpxg66IpUNAJCqTVBszlBHRLWLRUoc6ajHZUm4nu5NLpsxPASEC
fuB1wdUeD997WFeybsqumQ00GC93RsyYMa2RjsRHe5t2b+HAubbaj9R9rr/jg6GncyQFRkNzxFgJ
sokeOJGVrVIA9HBDnBDmZt3r622CFwtbkU5V2d0WGt/2CpgiFEcWPhOUpQlfzIo+9vJyetwsqS8k
X4xiOecwzOVD/B3iqE/Tc5P+WAIGkUXvuK81DQkQf9I2q/OHxwmDbqlBwVyuTSBAXgKPi1jLI6xp
iZt+AWI0u0vUKqeSQqJuQMdspdp42nH8vWtgNE7O8fgPP56kdhvDgXd+ZdCSZF3tr8/9ebHFqIgC
+wRf0Rf9eZR/5J03LJb48zkyqN++yJIiUo12kSJhyYj1Adp9ShdTiD/LWt0jgMVH1RHTKeeWx2JR
ellE6e0ptpVKw4AmsoplU8iLq7rK6O1506m1jq5p30Vy+kYfNJAgWT/5Xh+o+/qKEp8ZMrlrK4wu
rd6n54NCx+odgGfSDCUmOntcupcIwvyNQXKh/UHiLrcY3KA6eMCJcAi+dX5SrqbkCapc20U7cVXA
k8v7RQLIKekv61GIakugdlqVMivpcwANXmz0IDWjJGEm8wD/zRgIe1OpLDk9mNSpAut06FB81uCt
wlmoJ65JrWd4qV69doAUtdpW4I1LsN0V/DBPa4h9bMmhWCJEEaiGjmYZ5/aIWBaAxp/XEkbXjL/s
/qfxJmKD+eu55Bt8/jEQf2h4z7btOve80t7qTdSLflAJTxfdW0L+OFWcyMVdspLXOWpFSQ6+xlyW
64/6vKd2t8+YmpvB13h75lLeJXIvnae5iIezpDdjT0Tias1cQSdnbe9ew22kIySNO/8+p24xbYiW
mqfMHh9dmjVCjteeDW1b12PpOcoceV3LoMItK7FhOp8SzjFLeMPiA9vDmZ6O5c2/ccAMd5jayAwd
UzjmZW8KIFOgI22vS/aO3YGj5Iuq+5n84O9kilRftfvJzq1O4GNI/6hf9a0gX5/1HltW8pU/L0rW
52i+INh17sB5/tFrIsiP2jWC3dPRL/hXCsPGKuyagC4ADITJc3ELi1tIbqcu0kaM7ESLu4pVVnCG
5sCQ/TcL5I2kHgS/S5tp3Gg+jcKpEx4Kyx55XCO/FAAdlV5F5ijM2f+5AeVvcf/tema1j1fRoAsm
W1mgkrSx7cz+A2ASz5V8DLkTn2hLzK/5VHz5KJuVCjifyZUWQ5VfDHN4R8PLdwtjIIhoJds/jd6V
F8GiQSlrHgHJQqswWKNxOI3znlCVy+VCNBs5w/UJz7Rxlvj6+f4v5ojjNdRixEOd4nHV5VHMln8R
qaJ4C7n/zPNky0Z8m+k2qrVVi0+n1t6UkRQ8bPjDJNP0SVJIonEWxY7Bw1aGgFi3Fl65vB1RBGPm
j5ALHdoi9uTwNMOpQvbON0MKe35cmEHeckMWhUO32Ei4u3jhXP41JH4/V5y9doy3MPiiYmQNmESv
BB6TAiF87LM85W89CK1Kva5eO0cS7lD1Cl482Bcn28a1+/pBnFtAagynZr+kNgGhvRGQSmHaWa+O
v5DL+7C0flKkJof/PiatmNWwy98g8zhp7H/yIdJJ3/sKC6ZH9l1juNmAB2D51Srq5IjrOrIPQJ5K
fQoshhpDiPoQuQFH3EPR8zOZUcR8hbWqihEvFhJH3Uci0Ni0VyC94Zw7Bb4VYeM4UM9xHqoSQA6J
mZ1BO+0fsRYEqExTN6IhpImVAAAxmL67Af3cQIGdiTNhBg7UUhmsZwTbyRzNEbywtNHnqfTMBrz3
3c2Kr4pkrkLwtVvjE7Qjj6tUBBUb+r21whl9BFvG0PVFb8z1eu0As6b/ARQZZYXN4oKj8bu2N0/i
AvqdyxTlEPMlFdmSlAwjERGa63xT2EhcVaxPpCtCZg83w1Y0E4o8DTD/iA0yRhLYjdkqT6CA7Mul
sO4jKbvVdZi6Bt0yeP+ID2JH8adjAyZ8Ic4Ui/vAfJLXsu5fOCeweE2LTU5jh29eb+9tgDjRL7Ye
RHzmvzgNTczY0ABR/iAzKMcmCP2+Q4Bp+7TWMedkXUb+gikfpITqXa5wPkViu5A815TTzKO9to/M
qzxe0OsdOwzpjy0kqJXMU+1puWbpxjm35HOcrYM4IWlQZLA4hrwLbMQHkJkP+E8g8kA2GieSFWKH
VNI39wVfjTTv+HGYCNaYDj/wIUR9woQmRYFd/8x8w+qBwZcNIuXmdBhX3/atSkHyn5fQMf/JmEMm
eaJAqbTocyREt3DwPixCxlDMm+1Afua2TqEl3dXjQCPMpEWMamFPwpjN0l81uVBJjKCwsTd6D7Zq
aYMOBjOO5XwFWNYbiwX2uraTpcXBlePsBFVsms4zYrQUa5ByoRGVT+AF5ILkK+v21NqAdB+akhCe
oGOsIMGF6DOp/C6Rgh17B1IBoPJoI7FyL0MKBnnr8QIlKr6X0z28Wut+9tMsxVLbKEtvwRXvArBV
ao+raw6p1QBD9VBRyb0Lp+vSDC8iT5UmWl5I5IOBgdgb8BSW1UEOiL8qchr5OKcA3jTYCkgrc0He
GybQOBIkNYE/hA6nKkES/6uB8h8jKk47KdvLZCmECS896QTEsQmxaY1BhqnvFPgsmeJZUo4idyRo
BL4kQ+qQ9YAnlyxKhjDgbtWcIII7oKpZC/nYEywdmvAD19p5D+5XXtiHQOv0E1rsbIRYHbCXdzuB
YFGWhrTzmrbRIe5QrUvfJxOwrjWSKwXWAaj7lyyrGG853wMakFUelG7rchRuBmk8FL44XFzehJIa
R9CGi7Jesxe5yho3M30pS7h7w2Lu5CDMy42T3vfuDDAtLzlgveNHUgVNk5CHCQiSTWLizPOjeu1L
BPP+8raDoiUbF5Qs89s/ezQ570CJZoncUywGsfdVd9a58JY9B/CjuUD9idluZ+eCHUqy1AGUaYcY
88hVzS7wyVL3TMGpM6QjdZqP7a+Z1QF6Tqv1Q7O4oT7Y3NpfX+DGfqKEs9RREFAb0aUDyDHJ2YN1
RGBZ/DCXnvtxHk31+N8OPIkt3upBAvHzKTJfbQ/6CKjjYIzwKsA+zt+RH/73+5PVylbFBUrzIroN
jQeZDmG+C1UmoIpfaRUePBhqmubuJmbn71/qBpqKMXzQBHatWbO8zP2HK3Ge/DG0R9pwwOF5awWX
uingT/1KBDeUMiBeQsTMq59UK6WNPrJngtCT8RBfhsQw7zLIJ85bojgzrkumJSW7uUxSHEUvd+oE
sMWRAVd/j9n4xcKAvohfD+sBzx1W9MCyzxQJs6OF2MRfcSd2IDtc3Ad//z8Z838G7haMitJ6Rohv
wT01BB3iTeCnNJdtv6KdEWVAd7t4BuekGGJM6kQMXj5tEyoMeqnjgLBSfPGZIrK0+EDQf/Nv+fmI
m6bFwaR4aq5WO603fvFyvtsdxNkuaWkFvV0b+p8NJ7OxMHX2MCKwGV617cXYHK9YIE/oEDB0TdIU
mB5ooWQjU0reSdJNnNotb0qaOUXQXU8ajQ9Exh7j4CgVDKS1aiQBsDgPVbxlCrmGzR/IuMgeDWpx
kr8MneeEhRVzFdVcjmBfQuVjeDGKZYTvUE5TLQk2+cXaT2R/Nmh66wDcjO4+ZRIdhBbfUSF9+76A
UNxf/PiQA7td1dHBh7k25YxPtMofslz0lPGraC62hje7IYyUvQ681DpZnXv3nClzX9NRkTdN4x5k
WZlMqxUU+lOp+JRffY2QH/7PZRxccW9dwbn87OCJA103ANzXOpMWx/3TJXYkikKaQz8Tqjdo1s/j
XH6HPgilQjbVLnM7JuiA4JEamN9wb0HeiVtzo4tXfNsK7vU6shvWeD1pCkvaYe+SRrY9CkMQNG4v
xSVga/TwfhVrud8fiYSYvZUSA7eTuw11SE5+XiNb201G2gTkHR08kv0n3AY+2u0A2jGQid2NMsW8
pKtEW1A/jqw0QPuj+m5FCyQrFXEmbxBNb7hBLyiBA23FzsxoJNhgWJ11NcMp9ozMuruQjONJNku/
Ld5num65b3BOCMvdVOtNUOioIuBAH4x/WeEwfpvRnwhy8JUe6vHo3U4bRFfnOYtXHrcnjz2n1Fhr
lnSIQjwMWHPXzK65C+7aqEtvjl6sdO2t7wYrowhxquTPhZ1ars13WTwu485Cqyd2NGtza64rvQPe
AmYt/4feQqFuqtPBDrCL4R6mzTcGYCGCtEM5Z+6NID/st7x3Gvg4Kjs1ofu/Fmk7oVSxc1mrWUOP
9urbsagx4OcvWVsN9u4uHZCnS/9c7anxQgWnjXAaGBrc8oTN4jfx+Or4mn52kbiAgjSjq5TEdN10
nYR/ye1Vp6f2wMD8rpR37I695JwjBBmQeoaKo0rjAab/+sDCQdY1pE1Q25oMdQ2Y0z9Sq13PtGRB
xJX2skfYsruEkyxSpEcadcCePow0Ry1DyNTF3y6p8bZj2TDtr9mFREr3UMyZbFWrfwH8SXEDq/n5
BDBXHu+fl6ImkWgUtE12Tn0w711b322VP4HBRwP52XLiPjuDiVWzsMTz/pzSiJJseaEGCXsKF9Jj
g93nzyeEYybu+HvUDpIxdhaZOPevQ2msS/xDVsRtS5HZsIwgvudqNl0S0FCUi4bqujXvbc4DBB0/
s4OndLr2aItbD3eD4UNPO1Zf4bj6TgV+8ah07FRUZgE9OnMPDt+3O0OpGbGW6qsoTk/FctIRLmJP
bDO7HyGUterHcM1HP2GuD3F7QbqeZVxNARWPTCrfJodTMRsLOu9wU/4DIxynTgMrVWz+18PdEZC0
przRcolI56AG72Lfn8FZk0pICRUaY40PoVWvjJazofzlhtg9daAtTewtyY4mxv89oidnRaC/cIsT
pvebKQ07RR9pARgElaoG8DORMs86iy6FkuwweGJoG1FCrAx0PpcwOyP40EDlcyh7ki8Rw1i1Ubcd
a6Bll6AxzE0Q2mvGjThDbXge31IH48eCHMF4qKF24UjZv5zabiAj+XH/tDtk09cHfUxlb+v7QB1l
yGGo5hADLafVHYnu5NrpyDkmKjLjMf7+zg0QEBSEYG7d/i/9frukgZjQr2egbyOOZhqIqNkSLAye
04JoKsZa1oheutQj7KlsIMoews5Fh4uCzcH24k3+SXx57wvm028yx+be1iSD+aVqoEHnANhHXcKC
A6V0MM4nbDDk74N5DZVq4Ir0cfruSWaPvhIpD47BhVqb3TjOWNAvSaDGtIatpzHBHK91ci0H/52z
SgKuG9JVa1wtwhGMVHUiy44VBfm8wSJ4Q3yG+EgbvTKYuTBjRzdXlQ5QHkI2ISWgjIMsiSHTDbVg
UQLAlOYxhFK2rZ9mzjqWO1yRkrmxfQ0gfQvBcX/z5jcmUL9c0PXjrrhgomfFGWM9NF+gupA3l3EW
s7/gcmM1il34jP6WgYqOEWfYptDzYlsSKyxgoUB1NjWoFyiPB0UDyjzDBGQlTqUkxmJJXYhBXlyc
Z48OtP1BvWKT1fepZFGxKEyw5OYpbLWFcDVYObSryHcROIv1B7y0EPwVJcc5fyyK/7bN3eDQstkR
Sn741C41qkI5JU2SWUB+g/8yjsvsTooxB8htGrqxXvS2dqdJYm57LZrnxuZXgk7qJD9zWVCDg5G+
YtAng+sT4GWV+Mawfbq6s4QOHIsjOoTFzhdWOQEuqJdganbkJFsZADyc3A30TvoeHtjlhwV06xDU
WE+3Wreu1a2G0CYJ801DXaSrjjUKno3uSp5LAARwi4Weij9PvaZRrolh/t97HKvI/YUSmI9vwyoy
1lGXVHkC2vsahY583oN+Etx/MQ+h5oVAyHCzkerotrlM1xRKmpsV6hfcKP4t4B7HJm/vtjfHU1Z6
0l/O0TLwbyew4gLkQ1lEdGcrkNXzKCkzmH9K2rEWDsQ1ZUgYsopTMbd/9Ub3+j28RR3kDdDmu+kU
PudL++os5XU2wJQFGjMPaJ/arHldEpPj09N3lbdnzbEvh7yaYmS3OYL+89Qft1JfKt8EHydHLXQn
1xao/ScYxw9ndGM2QsGQ1bu7w3j6KehWhEvtXMzpvmzl199bhwEuV4/2A/GwtAyoGfYaFEQ87n7n
2gSHx/Ey4i8enYuQvBhTmzgvVclZFwHkA1g/SMauEJJZlJqIYFs7/atsuYsqhC39igwzPxDVGxxO
Gu375cMg8vaI4jTCf+CNgpGR1zX+IOBlbsfouICjWOZOxIwm1AaCoR9Et4pOAzpWenOUpNQMneO0
leSnVxLrFl0MgBPi2I/govIdo3p9i644nl9khuJScQbg5F1KtroKX4BY/tIOqPii5Gx5XgBLwX1d
/6x81uCQBczZUETNf0zzvG0CoPudF6FoRq21siwLp9yqyeDaqAeUuCbOzSlG3yQ8xHA52pSURwnm
/M2dTiHJtLKxucFYyU4n6V2we/DQcAaaDUG3pmT1A0MfFm5KYOaKH5G/byo/oEEAYxyMk1U47/ae
zaB9onXkYzvCmMTRqvTbf0FW4qyey/+oazkPPpQLhOZiACEy3MTDLie49lrJCq1febOx41RpFTtp
Fp6voJnPoNpa9qmms/10dzuLOz+w20soUjvGFAHM77CYIWnrwChd2CEnWvlYazyMeD3FLSjeq+Fv
SjvlM4pJ0GnNU2f2aAlqVOgEcUQoY7lnqaNhnbIS+ekTsFXZKT+FM9bVAOS+EZB3vDUbpljtQIjS
IBQlrFC5uSlYuIO3vzm3hFGBszn1FpFcP7mjhsv4Qu86hVmsJnCcUMhD/NKvNtZMXks70On993gu
qpBJcPDe2xlLnD+X69R2C3uqv16mF28GzV9N/Dw9ga0anQZVwKPYlQxXRVt/37DLavdMn9cbHsQA
RHPTeHL+wWGIenHJhwe2uZZl5ACkEpQ0PILnS5VNUlFAXdmK3I9aTI+cGJVNvcYjTc8ZB+z5+mfO
n5/SeSS7RoKbWqwoKv9rpZ4CDKilhMACcGLIL6F+naZcnNKalwdjuTUB51dDmazyqWuN5uP+uOXi
lMV6WFqu7D0pFounMIuEQvPiqKO1LgcK9VfIrWvVJuVyl84M1I1toZvLF48ruROoy8BH5W3BKJnq
xwSWY3B1rePIQSHwu3F4ytdEcHaCAATnKwqA/O69T2QCYxoqdkL2tcLzXuztMOXS/3Q+CEUVXTIH
beRfz20tBwDDtL0WLM94v5U55pwvoWqBj0UbPUMInN1a1V16ZWa6q87x4TWZx9TXMZD9riPSPoGv
EObupychuYLN9jPfMI3ZBZhHViyopcMameL/P3v5xJ+OhpLl3DI5Cu0SRL6QEN2q71KVLUZ0myYO
JuYltmfOOdd7tmZykqzyzgBuImbqQCcM/nL2LiMo8jq71HyLAOnz/tdM3MoqiuZjV7Ts9R0xcqfE
BGB2bD0YzK3OX1zXJCnROGfpKYNc/2cylxIrMRUWa7wiplcwoUMyffxmzpdlV4Txl9IcRRrQmomY
Yv/bN3TIGdOYlY7Og6gIVgdMjzk/GoQT1oOygoUJ08KSFPVw9CSDn+QmO4WOw5s/Gi8On3oqvp7d
7xwMkD+9xSQUPppJgm7BQvXw59ZGgGsauL/ljUN3noCFPR0ifoe5lI0rf5Mksyd5jM6cWCAuMKYu
uNo+5ijzp2N4zgTkl4yMjOK0+NTf3H8FknpxYzdWtJWckVh8XUJH4Nl6jTcenI5mfDvFpU7g0v3q
hwlTK8qkbZHtCEbUzihXrbyKxKjLIU1UCDvfq2golow/+8VYRTvVDpSRWnYyRZxVb98nQ438FMxO
ZQiSYGVjmanXo3xrZdtV/2TDqRUKbcJy4k09gB0oqE6F+EW06peSirWGwQavxUvFdeBJECDAAL3a
ygaGIuZs307U5/p3YiSNVbO3UILW4P+/GoQJuErkFafTwCcxX2XyOwu+0t6anzNwb0swhAvaXMFd
E17RuFfyxFu3nUots5y4XC+9xrx8UwMsMDcpEaj+HqePxmDrH4BHYrRFnGbR6g9qgJ/tnQujQD9p
LIVzTpbZezlt5XHWycSskfVvpsF3Ol0ZHvCxZEHi9YkqmSypDbQV5DCmk4pnUz6HXYML+08EY770
MfiFCG6oeu/M9fJlvOJNwvou4FqF1gLjyxMURrA9a95NontxJtUG9HPaTiYwyPS5/q6MC42ZuaKr
V4cvRy6JApfJaU65VlsitryCrgg/PyXFC1bA9uI4C72dl3fnjBKHGNwLvs+wPiTZRkd94H9EYxyK
qCHKAFDlZf7IED3vd6tdS8Uf2D39MUDR/mDeuVJyjhwqhE9qhFybh7euVCKCmio9zDwMgnnhTzEB
QEkdliLVqmqZo7O09E9JEG6WApeaq5IljitkHNYUTkvoFrmkzNvuWf7j6W6I9bis9QHinMIjMGgQ
4VQJGZJSyGiiC7i03gukHxohmrMsGwrydr9DPHaCgqalZnaDa1BE2EtZnTCfI17Y3XflTX/FgyRA
PC/BsJP638ozhppqyGHPqvuw7F/Xuqemiibn4O7dChqKQZdEgjRppRvkNFHOGbKxD6ZkrA/Jyk+J
s2enNrFonIhkQtqXwwoi8A8Sas8wsuv2nxOpiMmOA8FP908RwP8ZZxByRkZg4Bk5QHsHxXzULYDN
xlUtzV2wx82eD9gBfh81P/Sn7bG6Z9e+ug7bDXOREgET5sZzARycvsj6INiNje45vqtEot6abjq7
UMXqT1T/3/jzk5Hy/OP9OjDwEGTeLkPB6sUhSggFhgdCxrHEUezmBOl04hK9t2/1ZXFJSnY7dOrY
M8KVIVj1rlW9Y4XR7a1aHjc3Vpmi6zHkTpirAp6h/KQf50AWLh+9zG+jn96cXUHbOX6lYEH8eTeF
0v/vrngvhJVpLB2sszjgnWyLddvcxz/ccL3wmMdpC4TQQtVbiDQo/VY+fV6tvMuXu5XiZrkWZ3qD
Z34EjaoRdipsBaQGxKjY/JGXyi2ZJ5zGbdUYGxeHRrqNuKhp12ZsLBPyhRJWda2AkuQIHcZzJiPT
NlVv3ZkDBVFKhgKlqyfK1gWm6003+gAqwLUmtcmRT+1lyaQ+/OsSxoe9NwtF45TPSzk5mVRclziR
mQa4N6VhdTyfZtiK/HzP6Nx7pKKvVBsLzJWP5UUxUXFFu0y+n1Znsb0xSRnqJ3LHd90k6qpH7m6I
YhpnXalvsItoQ0o7zKZfuq07XVqX4CtH9dbveA1qXev/xNJOvOwFi+kEJmxjJXeSYYL+Z/11qFIX
jCOkEslYdHOcoEd8ZD1Y5LzaS6x9NvizMrzkMOn+/LHPpegk3gloRLVBNMgEOy0Tbjb6gRv+VKN1
v6xRezAjY/fquGuSpYcBLHUkqDZEBfSi7GTTtvcf2YV57o8W/4Ed1htfIQEFU6Vf6XzMAfg+ImNK
h+kqRVzrUNwGbc9c/WE+vVbNgY7I2q0fdwQ60wWxeZkPSA6xFnztbuXNx7O8l+0ux6SFFjpXx7qU
Q/53K//EdYHo/vgQjYAIlx0s0OAZenbJ7wPU0WzN7g2mRI3hpTablI18woCSQto5QOYmT1JWpd0D
imruo9So6FbAaiCNsRASoN7+dKyQtyXP5VgN0VE14FySZIqmuQRcAsB7rna9ChXeEL7iBxmsJZdI
BX6JFbJaPMyTuK1fCVnps+xZ45Z6oBxjJE8bWp47KIsifek4UCf8cb8D2JKI+VvW6rQ8xAKe+lnT
t7NSHKMMCu6o645duwi2cpw2aZ48A+Q5FIL74CVUnbiaaFh65box4EJbxMCD8YqsMi+8uNlGS4g5
bPaVJZmtDLQpNpH4Tmc/XANvqTlvgdyAH55B/EkqMlM6BJWl2UnNA0G0H0FvtrEaeOK19TUbkbGS
mSbi3jAvzTG/Q+21t64xhdHNO48GjJyv5EvaUR8WC7eSEwQxrweTSyldcmdGD+yp6Frk0BPjvlLX
eenlqBLBHtmRpT1IGuPhz+bttwl4f8DLu9kUDBTq+QGh7L3/yPo3FzZDmHQ1KpjFDVTsaNYwHPeB
hf2lnnV61kliUT9K1AKiCbU8mQTEMugqMFkQKVRkWCNRQu6awOJ+bC4MHtM+LXq0RRao5CLFB9PR
EhC9n6e3ILdIaolDbig0YbazWXcJfKlQXFXCYr4swA2GcNc/D1W5XHq2RMDJ/r62u2KlCc5gIeYO
sBj6tK0hUV3GJlVNqwQ0gOpmURjrjIJSc50+PWS3VKJ8NEv3eIiF87rkAChjKSl6rTz7mtfnZrZt
n4sup4BjE9y75WUhsSNmshilGsg/ODTEVOo63/UoIJ4ZkqY/DJflphO/8MdJB1907tw3E5fjtX09
wjgEFi8KhSik3cw9ZKm8jVTKndNjNo0CogqKxRAk3JkITS6NwntsZZWTgrv0LziR7Qx2Lpus3DAB
j9s2G0nSCu/ISOzfHpwAm+kPZ2OKgbhazfDt8+878UM48vpRtoa3TViLNIgmMRaOSpQUG1j6XAyS
A0qgbeihTtm3Ll9YjUR6L94vNy6FJe4vKKXxbEZLEZa1jiXObNcFOLF16z3GEgKphmTbYmxsJ8b6
ddAIo/YMAri/xOSbzZ9P6lQQSlfYaAt1qzkOZigqJHf6kp/gb2k7pwWUBm1DsQLn+eXoNKyV1q2j
afSLsMD8pximlczqWud9sr+9ylYCQp4w/oBQhNrHjsBMT6GZJai8tmTURxLOylhO1cEi/CJzkIj1
36r/aZD6LybG9QsOPsvDIUxGlU9xYjZFiF7kw8pTlmlHuCey6PvPu1hRkmOXpW0J/00mrDyJVsGx
LkFOvGSU/SrwxBnJa3Usr1Fz3zEgmt6Iss56bchE8aN4G0KWJB2EMJ88mi10brbXe56+RSPa/cH9
hc+rJa6jt6ZxDojzyUbhVjAT4fCMfC5IRKCaJwuxW0oO01GVD4XbFQAg+YLx3Fll+rgsbu0otGjT
2nwRYU/Ht0wT+qIelaqY8hMdjHN9raQ3ymhQVpZFqeTRJ7Ov++SDAfjSWvGR7prkRVtyd4gr7qbP
GpD0XvYEc8KAuT/iPKskOheAJf39JEyXL9nIgFGh8oG6QAO61a1ml7Dgb46At/YFTDEpZXSAHeUN
J8q36W7Nqpg1xepYGU1jmAeTpptd5VnppFKrIqv12J9zKf3jbAmyziZJpPI11x5uCBJ76qg2vGHM
S+rfPcx/tYCxfGR+V2hgx2tJCDI7B78tvcBtQczFzSTVx35/BS2StVFcbPN5G/28BIyclKd1Fk+C
7aKn6QyIPYHmtNIfzZLpfvBSFX2CADYjOmH1+qV3GNZewjP1rGHez6TN2WVAmuNIohvyYq2BQT7Q
oSo7xx8PeNbPNSwt5R9ci9cOJDAOACUWWWAZw9pfyKX/qY8PVeVRv5VH56G9YNF0xRmnCh1UXBmQ
lEiWhMX6IkiF9iWzNF2w5SK0Hl9/xqBxIBViu1X68Rs533tMOzCgCRdEgmHbXg7LAhsxhU5X4W7v
RJH6YccGjA2barcq9ZYozdJGv9kHVMbqOvij/GcvO7GTjlKE20UXDMxylqbUraSYXQXkHvRXEixY
ZyxELqsZwd+wrF3uDfFgAdSCS1HssBRK4onDZ1EFQw8CQeamdhCez+XvsgldidJRyr7nKznglmpN
xPqr02cXKutbflkHBMkNh2duFEXTfGlnDhGvjkRhAMNpAfXZ+w7RrpQobXWh+kBBL73nlV0RSrEv
bQl/fTBG4GwEsfIyxLL6xNsF85oX54PbfF5LQzIxEDOgrg/gtS8RjHwoOMRoHdIEcgJbptcLMssl
HY7yISsEoypVE2uhHCeDKOp1nLu+u8GdTui7iNB1A+bZanVqKXiBXEqj8Xr2wusqquHCap18fJ68
I/xEj3hxGmsLTpXRpcWc1eCBZJK7afp/oGegARj82ER1EA4JOfqHa5mE51iF59EU+o/U/+qmaMGP
1zbb1BZ6MqhtjsnXa0/sMNYau5uTtdcl6SOeet5Rz5H/BLX+yyCXimZzmRH4TqxEitcogvNcWRXg
A1bcqhdLNFcbRC/AWY1OxQ2HjMCiOfVM1+aFRv3Qe7gwQzHJMbsgmJvDzr2IUT3ibJMmBdGCoRgO
+roXPisqDsKSDXgzKHEAXW8Ft99Ui/72fMsFd8cQUPA8aR+4iXB88EeEgh+/16UkldS/vCQNDRwL
5pkNckZ2cC4zN8jfwL8cOCkmyvUtEu3gfLEK0CLz8roJ8Oi0u3OD8CLlHo6PrZ0x56UJKK2REqrO
J7YtHek9Da6wfxxJXqPpH4myqvqBTa5W+zFROonL3rXMXZNRDVgvV9P4ALtg3ugn+GfPWcMXlQZC
8H0avobfbvJcoJgbNXC3s8idt7+YVKpba0WoPwu+fJMh3t+nELJXWwsvuZbiX386Lw3GvLY9twPf
YkNbIFJTW52gtfF4Wysd5lTgSuByhP81xLBdnfnZ8CjYbndRhYnbqtFC50MaxhjBx79GrGP9snLY
kouTr4IjbwQ0UHQaw3zjW+FcRb2U/+z4v96k/XG5wWNEInOhhSM35cXCjK83SonaL7qscZDj4I1h
7R6hjpdlGSDQdKuH+bENEbSLgRw4x2VUsieXej03Axw3z+6Joy5q0f4z5e1bN/ZpQcN+x9nI88JF
4tdzlpSVpjzaKB3EkPBbQmmwkmbn5zmTIeLFCzBH7Jo6XMh469Et6Cczu/AZ2GGgw94H3ceh1Iqh
CkWSj+EDFSOsmvYSLkXX1hUUqabcdDHt1Dcwr2c1ae3gcIRAOH7iSLKMGkKanqVe/7HuQJefi6do
J0XuySuwOLDzeJJUGC9C8FhtHGE/dmsrEvalsNadbOcvaV/Hfu0h4by62lXMBNzFIqe+96m9RIDp
dIT+477Q01YorpFATeqlM+tPuQyQ8vj/GhWxC6+358GWjXXtxcAqXgJmfyriNCBOKeTAT1/vxYdq
K0bNkndxKsknCHlI6ogeO/oJH4BEabw+03EAlCFup4UESzaBncN1HuT5LJL02UuUGxCBvXZadEUS
8TBI4ApRhZ+FloxzhM1DWK7/6ieKcVMqPsvMrsDG33B26Gk/JZcZABEkUaSBGY9VOgONhRJvbs8y
8i0IAy3zKDLjpxLCgpXMAlIF+mToWsaalcb5/BVrmMVSHb93tdAfRuXcdHXafa5LzsCuhbhjN3LT
6arXl6HjzxzZVFvKjIoKoFbyXGnNRUeSZXnRIVMT9qzslsBAU48UwEMyk0Fx1vqRRFMqVeLKzW1X
4cIIn4tKZXAx2Sr/Pc16XK867pgLe4tj6TM3YTGto3tQra6LlhzehqzQ5E+gRiDaOwe7XIc3JeHY
TJy8mqgkUxllTrGqfYBjzYWsNP2FQfZj+SjEHX0+v01oYhXQ0hsxkoIBnMM5qkCRCNnafpxknStI
fpWY8eIAKB8Dz9EIUgfdZ60LQKF4AdtMus9pKRRdinUYgty0KZterTLrKNhgUEkgzpxWd7HViwor
rYnofVY519bUUTSRwLUabaEs7Jnp5rk9Ry7vuZldgUX4jVKydrULyk0gIKe2DnMCQrIHsBQiJDD2
ATVlXAymyJsw6UZy/jPHZcGgmNkrvxaIUpfrpYALSG5b8//zVXB19BbVEi1i+5eWv31k4B6pCKQm
9n647kXN70ehXM0mPaQn1mTedbv9SSJ3Ma7ehkejxWsaMLP3ZjeDf0AzY5+yToz2SghJOi27D1L/
D1N3D7dsZ8SNE0FNTn+Sn5vma1xX9me3v1TPfj1M8gV4sdeBzzY7CRlcod4fjNtkNbjpTA8w1hE1
7+pqEKGGxHm/wZEMHjKS8/KwC7P8he+uwwTedA4T33p3LMUZJj6hgppcRQeKTEdWOXfy7IpFcdqO
KSgHt8D7rquSiNsiPY+bcAZREecprxxxJ8aWxyrQrVRnSpkroO21nZB0kCmyUfS0sIBvKl1OdTg/
K7Ld3SHZAH7jR0zgYj6cX2HhkvOIeY2fLvJYBzh+bzm2G4ez4j589tjrmuD1/iiulfF0cXFMDK0Y
7BJzbT3YMe5HFHxhlE6k1FKV1qNzIWl7QzWdiufLVKWthujWsnMv5YP2/N+OTS9OPd4MNSXPx2GL
2vCL+bw/KpgqYvDVw4QLzYhgmzleZfrHQVSAOji8nvzlEsRDHfLAUi16adRw2pX4ez2uU7KfNeT1
ah26bQNfitXZiswEcTgynanVpcr8i0ARY5g3iu9FaJzxQZNdSxsYtzeQxpgMbVqEuLWp7a+e2VzI
nuLtbLr0qXMgyy9ZZHq3sPF8TVfnxyt1to+WIIlvmCGjrNA8ZvZ/S21qZoLENjogq1tRSo5XVDlf
FoV+UOte7ztDRdphvDrSBiteVEOGWLlvgZ+XF2JxMvMQHaIm4fC6xGqCMfJhScjINOBAD+NsPN71
ewJC/GPYjQ0Gw2Zfg25VuJ8gZ3XpjvaRRemy/5FoIT/HkGj7vjY/zyjPdgrOwoZ7jz0p7nP7dGIp
zfDWPkz+pPLV8YGqHSdEzRpzlLn3HBFEHUqQ2dQCkxU39gcW7D7Jp/7mQKP5fPU7qoccyWERW6+s
0ng/n8slqFOgBDydpFeS5qAETkxVuAprdlbUnTPN4B8RsLrSUaVM74bdTxZCKlGHTEB4zHNRqu4a
dJg1fx5GbUrO4trvvkaLK9GthaVt7UsWxdQ/EPU+LGcIMeXjfXrQQ5uxsSUaRPfoxA12ybOwexda
3RRtdIjFB/OBry4x91wdZjKPACgtW76dFZI4aV1cvozVsDCq07wdzn99taO9BdO8i8Nfz/YngmvM
aUO5KOvO+wzZM4+QMUcymhozWDtf4H4x9u5W10/cgy9rYpDqAgRBpWtKskLSkepDueDo28HhfdMu
lGf4J2/3iXm9n5ngorTmZR4kQOLflJGM/SeS2sFBX6mNykRgJTuTxhrHMVdJHh1uMDH669wYKbC5
tCqKtQNofHpTZOnwutVMjcGY6vlipKeBX/w+dI0xMPwnIiwa+4YA0EN71LsyD7N3vSoH9P639Z9i
goGqZw79oAzl5J2uWqN0m9ziQB1xeXO5EJIFo30kXxuoa3/lnAjgRnYRGqdVn+3w11pfwPm0tWuC
CibAFdHZ3zO1mWbXLzftUVmhuU6yAZ//m4jjfqrBAyfCu0a99KLClP5hEMOtWV/F+nJIz0d47aOu
lXSpL7gPm4hhGc4O0hm0Jluw/LtvejAiMWHIw0E2kKXYcy+cNQp74kEqeSQNuwfUNZy2WZINHBFQ
2CuN484/5TVdwKMq9dmzIeicDN70yI3jyCnRMTArofq5wsq95FlEiBcuAhJ+6NeA7wR75JDzUptm
E8JOrlr7UpH3UcvqPluO7GIJuD56Ylcp8C5rvASIEdhhOuTUzWDsqu6aEmbBz/baTSWAOzfBoPkh
V49Lu+uJVo8Ma4OJw5boDjQfR3ehsWSzikz0yoZiren0v6FJ82tdARfoym8EIKYpd2o8naVeaYSy
L9NxgU5iIcBZF6t3xJsK+xMJ5OSX0R3guo/j+TyhUEcIk8kXiwxkToMqdKhra01gJ8/LYPtsdEOq
od38An6ypR/JIGiPA9beChjVPP19k2q+0K3G3L6JOXH6ue8ZQrZF+XLXBZ7VW1iSgwIgPd1ezgwy
jpvZetMlFQLNNu8aOknfxqFyUe4d/wjcSOQy4E6Gow6II37qbpFVddczQCIvwRyXS2UqbDzyuhPK
3nRTAa0u23FLbBSfkI1DBwU5DFMUB+Y+DUd+56wcEu4peMMJq7Yymii4sE64rYdmq7Kn13DkdNOS
CM2et0MknhO1CmtwuQbMEz81lmqPrmoMbnHDALJaHYWT8WnHXEnwmQV+hQMF/sLC1BP90IDYcQPq
ehH5Ywgu6lUzG38aNcwNIHvxT7Ld7+c7xP0Qxyp32jCSFYG4c+Yw9JEqG1baTenpj8wh7FQiOlqe
HZrc3IJb/zzCOpGWIPHdfbbQ/wM7av97jdFePfg3RoNZBFD8/Ki6OEf1opqFOwAgEmJUoyemEGNo
VUEC34JN/eN4n4vikDWrHVoNg+KDyqlHPLsL6WdNsDYCRFCvcm4hnZhgucKJVGazw1aoUReiasr8
7ZPgPE/HwPSvj2SDtM2XmgTnIm7EKLef9+wGOqGZM4hYfh/X6XWj1c2nXol49rYml7ee2NSsx8mZ
mQQ0iM4sKpaSPOQ2RVdgWCEP8u7vUYE4BRXFndFMdKZGpWxKUhfvS6Up1yD+aanAdBPXYpcwWps4
064LtpykMJbttf5FXDeRZHvlD1gin96qRvXmJbdgQuVsqmPoeE6reYnWYNg2RPFzyJJOUgsE4xK8
p6IelkydGm1F17l9pJglRjvBdzXW0cAjUhiQdWyEZjHtUssCKWIXwW7CPbfF9TVe1YuZ4HOMXq3D
n4p0fWzNdfbcOkxeD8iTfgXyO6V3IU/qsAojqY5Tvg598ZUdoQ5w0mt7Z6G1zZEmVQr7hkKgFSU1
MLkgutzJGDmbnIHIc6TY+6DRZ87ZhZymJGLzeGlmICd6Z8QDoSqWpguUckVurjQFWfSPMyJ+1Hvw
qAahOBrMHPoaMKaXKU4WMgweH6W0piZAKKPsgL+6j048d1LS6rCyNejT43DpAjZyveWWBf5k8Vjr
r+F6L29qS/JxjoC42cPrWZI7BClhv+eH0DcZqFwUI4RfignSPMnQUTatMxw81XF1FoqJE3fH/xCB
Fxn5CeEpbDpEB93AJG/+r0f2YA5DIkpRtaSl/W/OoCmOeT9sUbEJnpa27yxmXBbmjNDR/HPXFUrc
+nS8DZYGT+kWmlPIQJ/zs1rxVBcNPnKFq/10bDenypnhJ1prgw4TRnWV48rQsbyZUWMJTqSfte5X
X+KCBsMkRFWgbxuEOPtDB/EKFrQyWoNo0S6Z9nsBeWwqG6hFvtXKRVBpM91vUw+AYtDV1pOJFadB
7ZuCz/r/gWwS2sc7DzFf1lxb6+YVo42+nBraycd/G/rFsI8sHIWAMpdzkYGT3HKaqVDBgjb6PmV6
mDHG2OM2txmriPIuugu1T1dAXVoQNcMsW9ofkASz5ZdexiW5jIoNwuY0gpVQCdJHEg9x6Xv6iR44
PVaJB5wiwq/tEO6S2dwXqmuHiCZvOd2K+CXDfMEd4VH2hDNCVL6VAKkb/aLUyGjdYzXXxowQiPtx
+BepOa7A+koDkNCdPBnn2scK18lJXHYRBCdWvqaYyZLLlXMp0MNhAAjTs0W3vUFUCD/L7mrMvQYS
q9FwMvQxM6rUQc+qXNKXxW+Gn4x/9gPVLys1qs0qXg0h2CHrawhUXcb8He25z03m3RpZRxD7610g
cHLgV7NM/AL9aqBUCvCI0yKEONnz8mjsREyshkv9V3EwBi+CzWW8o+vcs+/SVWys+rgSTRUEeaGb
ND7hlI3TwEMgAG5VO7ByaqqyhcN7PWu2VyiX7r3IJ6RPE+N3P+MFW+lMue/9bXwMR37MF1O199Xi
QWikjFO04RMUWCqUkDsADZh29nO0mnz8RcMprbrUgdNlsr/vPDTlKfW3eFMiUIUKyOLdv9zTYkj0
5LqLYMY7XbEuWMyPnXjEmsENHUPeGwWGA/B3R0u16ZSLQeIqrzhrSGH0VpUMi0QGYwoIiu28n8jg
MBEDRrJMw9eOxnP2Ms93Ek+g/KFXTYJZult3qNuZllTgT8rE1cE/4rY2S24di3qrkurkcphCSg4+
kbhl+brDuuRe+p0T5zTcGVfOGB+fjwGJZiEYUfFPejvrTHroKvWATah1XlMzB6s+CPU2zjREA8Oc
8GfJWGWJQMOjd4QhAtU6R7zuVilyHM9iN48LUKpXIzByMGIjc/HE5hH+q4t9UEl2lEfXCuzUgMDh
BUGz8zcTyHOtHg2js49bUxJii7ErppCGW9Q7NCuJGr501q93m6pFwchHnIhx8aDV/5jmWAY4a/UD
gkb60NpsAA1egLQNUf+dBTE11XiQKZAh74CjFr4iURi1DFu5VrH3WaV0dFi8zbgNRegNmIVZYxKh
SENswaUILiYQAVXCAeqALgkpjNYOu3mO+Qrcru5V2vAci1P37oSLuFcug1FaqOj6V89QuXtY723O
/t5hBV8kdBtQA2moJP+K7S1r+AARlqKpatmjAMsnBwJGwL8r/yjJFG2WaIJ5ch6BL1/c3pebvg7r
WRJwk6SHqDK7+8AMD8veBQar2P4cwZlLx7VqE6bS38vS2/q4cCTZNQqJqivYyvtMI5u0H2d8ArA1
bF6pzHhGIlHxSH9mwt+KB2HnMsQJn+4VM7P+PPUHKxrtAXuCUXxmD/cGwygsFEPLSD98i/uGFO1D
kGbX+kI9zITsEKMCxDEAcL/7AbFLYrJFlEZ4JqYILyOQfDBK3rkadZm42wVA+K7AOiaX1k9qkkTw
ZlzKRo0KjJrx5fJPNs3zEvbiJm6bj//9L9X1mQp6xUz96B8eIhZQa3Jbl5SP9w7Rv/qUZakI8idE
Xcn5p+QRPwGu6je5cLc3lbjk7Qa1yQz2pqNmxJzYqsus0eP/sT+uEuj904oEu0IOBK0OE7OyFIN7
CX4gzRxXH8EqM/lbME7UNYAaH4X8n2tLd2o83hRZcyW6lwkASTzHfJnrr9QH9PylfF3E8uIB1oml
mAg8WYSeFXgVxUN5sfI+y7t61l4/tpgN63urJqeMmLm+/yvKvfecFd1zaCOTImUSQGrmTH+JXs7k
vaJVSQm2Ub0stLs/Yi2S1sCvAgG1RIhJ8ZtpuIuE2o8Vu4ZBWL7gVYNDrV/rE/+NYfssAW+jK8qT
faUV30zNU4rnLx1XNHAwOyo0WtjpcyLu+T3RjLgkZPsai0Whx+SeFrSRx3xEYoo1gPsbD7MThi0k
hiTtCD5J7/IFLnkay5TwgjjjfTqC8yG7jNdAMCqGfn84zBR5Uk3OToWyBnrUkUvL1d925n8D6d+h
4y+QmaNm7YFkys/ynBlgV39tFv4ukoTtyktHbjLNRv7l2pU2qB6ZxcMps56hPMCpBH9J/knTuBoq
V53MKbgzOt1zzk/u/5h9n/ZemAGW/WzhkRCeA8MVe1lYnTXEO3ZaNPrHnO/YEarJRMvwxQ2TV0fG
v37dpQ74yyL0KLQN5EfjyDrJcSxy1ok7hrGYWS93FPKnxQVLgpKJJWdlgjjnf8Hq+AuYUM+kMGs4
nsiQN/XHxrLx08wAouFzCbo6vtXyp8Y/DZ9SDtwoDKIvfdLngA6gOQ0WjBfOwZYZV/+Xk+vXBW3W
sqQGSgYWsLsl62RrvlP0mAa00ZPme1OWwDYCMPlplQCIcKXMXr/cH7OH3bUA5dI8pm31UiSOrF17
ro5G2tDGzeedQfbGc909Fw2JfT0uWvaVLAJGYC/38qTBnK9OeuTwhok6KccFctA5wPSluEt2q+tO
iexYd8pHZQuWvjVD7XEOrPIhitWxDCabl6PAWRD5SFL3LjA7WtOv2XU6tkp3gsGT3hQgtPzZfdp/
geYYeBF/Uuf7Wpl5T4nCG3lv2mR95BOQinTa5W+83Yik6YoDaIj+0lcjZ+dSFjYqgDhlElWfvFGG
4xPY+3Jvy8WaMJ+7KaqR9AS2pHqVCDIXOIaS9txBCYvASpBrNnX1xHdkFKuY7bMAxoTPMzwbNkr4
dFn9Qbr4hBcdR0hMwdAxvJK40ojdfA/WWJAh9Y9ulA81pUWfXcMrpmYvyyOvecjFNqYbK1KLoeQ8
mKKJF083IySoFz06N1TUGOigGzbc8pCjUbPumldhzl00PntRDmnCGVE5YrwLBRiWb/4LTHzLgAAk
laaZ0p3pqOGVPJnZNMDW4kVnbewrdK0/2yMJScjV887htnpKlptIiLtja16+/kOWqG1n3r0LaSEr
rIcF9qtlkHhh0xW/Qn72vgd78Mev3xGOki+OuPsceMIwlfQds2JqDZnTudQUFYss675lanyVRaar
dEjOsQ0dR1rbKXIhFWYbWRVVdXAHcQEA57X5h/WcvD8PWATgxL/tkWjRRw0lm6NcS6hVXCUxtEU+
qGXtReC9vukB7s5ROqJHtuvgJaDgTPCn7DLcGgZ5rMoYHNMJg/TL01z4TdjEfRu3KTHvZeiOrTzF
qkqSLlXMirnMlb1hbp2TkSSJ8dK5cFCzVY3rbUPrqEnhlsCa3PKsUCfJNANpYcn+iwmtBVx6iFFI
inxdLDBZrHLAuf5ILv8UP6lzUMK/MOfy+Wc8ONEdlocDavRkd/qQJjKuTO+jW18SvdXlZ0HPan+Q
1DWEuOtuM3vpU8zsqwyoda74viDaHVIWBLozTYYKZcCRQ35WW2axorO6OyUh0F1zzL1eZub38dnE
n9+pbs2vU1n+JhbULldHpBovPjl0zw4TaqkIhxqsz3tH/CkyN8USlfcEoQv5xiYCSzWk6ogmMaqW
bCa9LSCdtHN6Z33DsnWS0DijdoCZxBhg0spkYq7sKUJGpKzaLgjjftcnRir9a2dYQINxudTjO4YG
bcNpPByH4ilJbbIToUK5u+Dp9mWXk22+b7z8xSIIroPtirOFv9+SUf8Bvy6gSXodqFFOodaUgVUK
OK/12136x+2xXYo8QxAOW6lW+6Lq0OEPVbqkwvoFKwvSrfcjk+CdE3FtstcBfU3W6F/eMyAM3jbe
+15blHskP0GBYftOc/kJlvqXO7MAgp9ADd3nST6YBQla5KCYq+IVHZsiYDiWfTxz474waAdpPdWf
pB4eDDMdSPPkkvs5VS6Wnk0gAU2iZPjE1MBIJQqsFlTXOmz4Yy/w/Oge13CgVRS0hus6yypewOgl
Sc/84o5c//Tjr/jUb+K1Lr1HnDZGVfyOV1Zk47abZaXQpKmuJd/n2s7BLU5toju63yw+EsoCWiAE
IRU+WvvprZkGv597PtERs19IG0hUq4sXWQc9rkLNN1/UuWvZCOcfCyGXq/87qSkhySU1GGmuGZ86
WMnEd8iIDDM0cgJ+oQCm5TK6q47s1vtPFFHoDiVwQzHZT6m9/bPYm6KsRoD2p5BV1ru44gaC6mwh
czxhYHJfTb+gqnYuxDdJtmu6CdSxdN+VdvB2yc268m2aFxitNrs0+vXkcWvMbkfrePQD5m5cGp8U
qQioca5AHj7OjitgC9DW4PS19iwA7jT6LjJT+T2oBh8/5vBBWUZs3NLEXtkrmtCQ27xUkxhYhzrS
QRrqcjRZcNaDZb7uAeGz2suwWiyCchcaETNIHj6P2e91AEK3W3FIpxNFb+wdpDKyjmysYNFW6P3A
MmViSXBdWDnf7Rq3bFJi5UAuGBdC/BuiWYw8WJYTgSI/KHt94Bc0NVjE0igEMwPG3UQRkHSZ3QHi
8MzxhcVnnYAtAyKAhX4V6Lu4cFcBkyRU+p0CuTfinCDfTQ6rVRqGQf/AIROhQRsgFCyVR12Rn3CS
wZg2zIjOy3ZPsfwsEbpJP6x0h3xkDzm1Kk3dwz5v9eKM+cc579BgRRmNcAnhTAFSMd5gKO+GtaNL
kW4Zwf5KdvVnTXKjAjGD8bnaDY4C4w6xPjCA6nAJnNel2J32rSoH9D/2VcjWQrex9tOhJvs6/av5
P0SNWk1ozvmBTopsfz6mvte9vdqNiFm0gaQL6fD5FpkN0IJojK2Qz5HHh8iU5imIS5OwTIxuiwET
xKDSACqdnETl8x6xgoItm6q5jMPRCeDbkpoUBWLs47zRXaRQwVLId08DINDSLrndfQDledyBQW67
3THNbb/jzNHLqmsITsTyp8d/Xby4ZtvV78LzXqHsqciD1rRKUvAfRfw9bkXHRmM7Z16y5rFUKeEa
jIbu4RY85iL1O8Wv1dwPYdJcGQtn/aAJIUh7vOBjaLBFNaRj9aNG9HQ4X12urpQBXsrz1kzcqMzE
MyrsPLWmj3cZGVHIkU0FPx5WpFanNbjmyd9MpoEvLdrlLv5a5WZ+ww4wHlWUpoC6ZAM9UECqFSnE
Z2wcRPX6COoPo0jDKnUt5giTeLaruZJmKOlJ3wduyC8JJSRhpNCHbsgzC+PqMjJHqwN5dnW+NN+z
nH/Wy9i7j7Ee3fgLauXSKHmg3VULzqdhVDSf87Jas3t3uQDSa5+Hf861dhWjB877rjzjX6uTSOIU
+3rhBNC2hBAZRhNibaSCpw7ITBQHqfDqxQYJSn5l6k8Q6xzmS6eDnIzxy781keMRHKCdvpjqBMp6
icnpSgXwH0jRiNEYomo2JJGNDtrllbjyqrJYlCtbls2+zQRD+TAahMAmnpSbaZOy/bNV3OXoEAfP
krG/eWqFPF179ibd2q3kXrAV1v9LXUD3ozPSi++3FU3iCCo48kGER9TOicubppGE1IJFG50cc/SS
acXQzH5CmLtUQt8kz/dmSMYuefcErTIg21tn++fGGz1viBU/aRmIFOj5K+WnMjVW+Q0HJsCpQ4Zw
UQpLV3oC3UvnFfI09yu/NDBK06WLWkp23aqg/GMKIxdd84GC0/rDoBCgO8X8dBnA6Rnd4X9r5jwK
vyCwzT3IXhxWerGuUjdQc4A8KVUQHfM13esmvtuaK0DoBGWLVGdOxZR1F2QuhTuD1eOCsw6qyM3u
EdZQOyCMtcovjmHDayvr7+MH553UY3HL+TsfmU4eEv04VLm0ZYzNvb9l7fWX94eSmUT2JQcKykIQ
3Oi/e1n+NmtP/yKHKGyNLihDdZ8gUBjJ920Ro1E5nzEgNKFueesSDdOurm9mVsIHAwGtqx8YSuUz
OkkVVzVjL0LeEsmeKztgaFSkBVGphvYP4UYt72Je50sB/lR7WD3Hxvx7R6IDiDpFB0rAB+OslIFf
rmdY1IQWsZSxspmy+zn0/3BDkB6SXMo9PlFFRF7i295Pz8XCBQDWX/mf3cZ6FmgbGr74YLXdDyOj
xoiFRP1isE4koeDQmL8nHCADeqcbjsojce96ryioFHEqTMRIuNWOMQievFSpCvolo6xAY+XqgUBg
8qpptIPnuuY9ZP1W0b3g4TL6ZrJH+AVy2JPSxu41VbiDSz8HhVXNw1gvVyLVN1NWF8+jtOQ/mPOL
sZ+5TxZnbrSPiuuIgOs2NOeO3xpdrTYW6xhG4on2IzaquP7UodDPGwp1nL/VWNKEluC/PkM82Em/
ii7ftVb0YWRSDWLLl3pvcexoS8Wcc43j1fwrKivbFzw54Wmaf5fsA8qRYWktJCHxCem3fnPGUR2J
376O9pV3PmegCiUvPGN6fu5i77L3XcBe/BIUld0u6zB7uQW5OkvNOgt44cV3F/003KJ2hY9sZ6rc
KdNGahIToMBRX2JADENgzkCrhoJejZExsy81LQMf75zDgPKIH2c6KWpW+QcEqDehrnet8zzNLON4
9f553K7Cx3Nzm2rbkbRm6a4IvhFMuUl7AsV7yjUfpmCkuWnPvvvz4BwXGm25iksPvnZPMa9OTOAW
xPSdWDF7ng1suDwraqH7OiW34dqSL7KPN4OmrwM98wuwtVvf5vFB9uRqdJPvj89OlCiHBv3DWvRP
UmP8ca9SlAmgb+jtFc/XHnVpFoCDEGqFG0/cEqEA6Oh5uHQDNPVXB/m4bldnkBSR4a+BkcZ0UD9b
zPQOwI7jhCUjFS0EzCX2sOyMRO3MsJmK5eGD3Q20vt7zdOGkMwqR+RJL3WM9H0PgpDk5wk9Bu3sT
iHNsVWDk5KQ8kPNhYdmsC73dAVcIwFNoEvvJytdnmn9dmSACa1FHOxP972PFpR2jmVIOe6aarWH9
G0McdV8Aw+De2ms7GJs8015J1RyZWqlH+cCXduj14mnGn6HK8U2/OvdGmSTHH7Ox1LZSJ1NTmuwT
jfnDErXHGLBP0cP5sYTWjDM7i4VIezhnVwvVIvN0SVkISDb6dSbSbnhbYN3XNzSjPO1tWPIS0hWI
qN4ICW1BQ+FMhjASz9VsIjoryH8dU+pTR+m6O/SGdKZlCe0Xx6h29sKO7qCodARFluFA1YxmwkU3
Ac5Jv5ECQWVG6ZRJ7t8pWpUTJvRnRRHebtm7TgmCMJVK6VAadt0cGLYsLV7MVOSQTfOKh4CjtP3k
2MN758IrVPITf4KwuI4iy7RqYSKiMeq9m0DKGaDj4VnWlxdeuFbQfr8cZEcm0ZqoH5rGEvrijqGh
XNXGE1QGp2DsAT1/gmoKdKnqG9qiqUSyz+tNV737SRs7TEVknxz+WWpxiBBwSboSHI29XU6sSOqm
NV6u8c92aicZP5S1aNzHaj55CUkCNrLf9TODSwH+5WlT/R+YYoaZX6D40lHaw0tus+v98KBXIGfZ
++CQUTc+2xPwm6phONk02WjIFWtdCHAdAmwPgSIMDtYQpQDiDIZXRW3smkFnPkyhun/8KIdrdm7R
AOM+jLBpvHTYhKpUQd14FFhKs3SXSQ3ssO1sFx0nH8+xQjSqh6r0W7bFMnGLL9y8oUJ0A5voclmO
x8s9QzsPE1Y82j0O7b2ho2YTZyquTA8OP1mz8Wwy8gF0AulKkEnUr47v9XOpWSstxue5ZTqmqsk/
THXRiDTYnh0n6id7funUHTbRn0yIKIUKju7Do+LhJvRBbuP4kSa0oZxojtr0I30KBeoF3LetACOY
t2eCSMB7yvfc13/1AnPUGTQl4vKSsdAhJUGECLKlfG5VPJZx74onkLlbt8d34+90Aq3JLSgHQs3L
PU7LNfbjuna79gI5v/1iySsSs3JVXfaa5sh984YxCrPha67LeaEqwZdSP+aWpEqQBDfkKMXrM44+
sZJc2qKxnfHiI+Dc9/ObRbYF/DRVd/QRHaqbVZTo2vAsS08oWwSz7XhD2awoKcm/IScdNTgXrM3R
1T/8w2PtgMwDdj6mwV9rkzzjSUA7leIJqGDdmkzGAbbqJ+0EwmNBGnm4EfJBuqLDXim2QNOqwXTK
kFNTx3pt4U7MmvIr9JPuAtcoNNX9ICRz4RJiARVchTeC4gDRnGt14QnvSg1nqcIiW0oJWW8q71Kb
nG6FrliaQdMepNjjFZC6/1SvXK3lelm+8CIXRdftcVjXChuQq+73Iy6yvEaomFKUDKkP5uc6XpIU
y/ulwv02cf3siXQ2kxnW6NRuYvpq/dx5Hq3GFvke1jz8QbqGXPdOfVm1IZc8rLLZqOzpHXXhVIL1
LHqs0a1KI6W8hEW15Nrzs+ao1vB9f3QaL/gLgZEycEwwjNaElBZUqL44lzrqcT62O1E1lCC6PUVc
cPZlcy1xZhuv3b/apyaHjsU+eihkJbuBvJyhPzcZ6Mah8jQkpmGKAcIcIgxyUGVqTKW04WKSmwMD
M4GrarCD9WQGJueTcuTj0fRYshh5Zr7RASBDCBe0Nej3l5gGZhn/eSSRePjL2ooUU+gKrGSOQxRI
mpKbgLuFTAvh/6kaZq5124NcZQLVZxAYNHxiBh2rSd828BY9blg7JVQT5VRMHQoLX4jchnzKZU0E
to6krsopzpOtF9EwoQePAMzX/3u/IhAs0sHgq+Klam8DAf6NFSiVlCAHFvGOZLY48gpZaSwCdG0P
TDDnau5WFysEa9j/ZhQ6rNDQ3+pKK6jpIkjRjU+5huWTnbj6Ebw0gb8sTWNluo/DHbz20O8VKTfJ
4/J/mmsX9a918uI3o1Zh9fGLkdYcSn/yiZQ9mQ3AiXQSdvqVsvlkPI4g9I8uu1TBF5d3vDKKe7BX
I5S6atPvl/UCUqnRA+KE9b/AJVQnNbFEQ0G/QqjOG6NMxX2rqYGL8FD5gZkuw3hC4ull3tfxFlsG
iahdtDp+sKutzaAI7xQ/3KhWXcfo20VkQ8rrQw1PzkL8pV6tjVcNg2fzyD23kSy7BOoXim5bvNr6
BI707Alxy56uRKREC2hwuz0pdINiIYt+sInG1hbbhhlFvpY0oMbqy86rgcK5/NfNrZ1rLIC5qCAV
1RgRN3zzzk9oLlG2Uvp1X17r+EPd2zUBgiDaDfe7IlaQeEV+9yYbBGtXlDs8SB1V0tAEnVZZeDVI
8GOsWGb/k+lIx4sjMntkN2PhGEwd4oDgV1zqSfATwTHJP/sSyemF6H8FB7PoQpS5ApKOopMWaRwB
aPhMlolF05RhaCDTmZ24LXDdzR2dHlsVjHyKHFWQTt/yU7MlTzDDUzSe0I17y7sfqPNdAd7VhYe1
4yWUGBKg38P3ELDUtOw/pYW0O50TR6Z4rarJaxJKc+xbca7Jhr+xZtTwZd7XrxQXR55bibSzEDfg
j+PTBOS2cNNxOKAmxqwwk5ck3sMo0MPbm2UTHy/vX9vznLgeVZGSwH7ttPSUvu1thCgqHkgcL4ng
fNlQlmRCpm1hZzRABYFsCmr3drJ8XKamd9QDJuKhq7rKrmjI6J7SYmwcPuJbgbru530XS/UK0U0s
bWHdSd3TVDSzDxOgB912y9ANMb+UtHuosphgAABfELv7cMSNmdSDhDxlg97CizHHRApjjztsQkTb
Xzyb9gOMWIShmIOY1psM0rGwJcFOkCONOKazYap5AbA5o6q8aqVuFXagHhllxkP3D/ModknMMQtI
IrMy+ntHJzDsWBKhj8YTtklchrIi01XjQkxOprwUUuaNyttFO0zSsxPYdzx0XjcM+MuyePH2Vlb8
AcOlUHJARqeBKU2PJqOsEJDeS+emJ97jjhaZ2hYaPFWh2/4W9YaW28WiOEqKhRAeBAcb11SVS8M2
3rf4FtLEQbiB1huJO1qxfOlRha/gX5sYHHzjycVxNaN/ReXgD0Qb/AQYJNlNiZAmfxoaSBUaKv95
ecxSNskvIifLjxmEfjxuLHU/5B7WzW75O2ESigHFpreLKYITd5HBes5tp8xbT6KPPvxyHcmC0lai
CGo4ScyCtUbKKgoY1vTLzmKvibVzB2WCYciSKdLI9mFjCnPsIG3Wji7qTxSCV/XIxt9Zp18ppfyu
lOt7ALVrRsJzJGJl9W799r1xjRkQLIFLzbfVE2wWBj6wSl/xjDcWK2PKND3KAXz69pdnC2V+W1xj
Lc6KhFQSeb5rRKLwYWMGAt92LAAWW2CFo2wP+e7JXUNqlR2R2sxA03CncdH/1GemB7vgXcAlR1go
oNJVjNsLrJvRqOu9j8+Hdqy/IVv/3hC70StBqrM7IQAnhxbjImUy4TFSylf5aleRt9MiugHICHdN
Cgq3fS0iERVjBYpptBqXP92h4NePUav1TWTs2eeyhmGUdBsLumRx4M/uyGQXpjTk5vok82eE6W3N
qeaaMu5jDNIYD6EhzulVHvLQcDelc0KlDRzfkPCqifaYSCj5fVbh7+S2GJ+2/w7g3v814aqysrJH
lsE5M0eyO1s7c5MpAScOXfkhgLbrKWEx9qWNPEd/mZoqKM2URenfzcvAYuMROyAKXCT0vTngdkYP
WDgx2erO/RvOPaRC01zX7IMMTnoc+Gok9i3lSpkjNeCwBQcj0ZHOW/hzYTIZ6u5C40AlFv9s8Nmn
yVrYnX/+/fu9w+aTH1kjqtjcme8uFzV4fcHNAaRIA8cYWHMIVZYv508TmAsWYrmxChOyJJfTgiH4
dUApQg94AUCt26c7vG26n4i8QeKSUryFuTo4e1ij7co/CDYxI+NB5dHaGYZGnmkWxEFr1Fm2s7si
j7U0bgu5joEU+hWgox3yuBS28Cd6+YddRzDj6oed5liZamfXGHrixQbCuN+Q52bFqp+KW37FJWxw
2hIKSddYQ/TGboDbYKO8nD+fSwMGkY0YSeX5nJix4mgwHpgnqQepU9lupkgc0DjYeylnjioNN5zJ
oxLvBjo0R6OQXYiE5ro07BXN3+oXoqPgbHDB3xCGg84BixdLyphV10C4bGawJrZi1Rgr4ghZoP1V
FV0f2pqyKUxHkCERXYd1mVCrxIQwPdUWArOQuRmWnc/O5HmdQ415BIAHFwDFW+dF7Bs6wJiQo78H
qc2gQeZgz4ulIoiwB08nVWYhyzzTCixOU/bEjfKkCAkmggY9n9aMSMieZ7nnc1Djraxnlx26FT/A
CTWJQUZKsRU0rRqjN+GkOBHqhU1X4Z2QVRfpeVSWyAJA6n9+Y1EwFlIORFqCxLxNe9wOz6QELVn7
eAEKkf+9ytYvtvkvViGLqO2sBAKQJjnD2QBNEiAoZM3eOsXTibhBZLr2DUEKrXLCva9Kj/xpzq69
8EklzU3UPpMDGtvodzgY/5B9ePvyQE9RWzgF3OD4DxCjBmAyPvRZw4VHmtVsUs7X+HeZBscwRVWw
XNa5Ox9n0JQGxMEOCVZ/l6BTq8JO35lu+X/F/9PzzJeS4SrBWY63ZL8TR9I7H5YGHai+d55r6JMm
kyfjVmkhf27F8X4iQJOpkth7HFqL+tVrWg0lUwkYfgvDYTdSI+VMeXYJdflFOR3i5omztxV5M/KG
lwVbuKnCnOb2QMkYfzyRs7hxqrGjF6P+e2lAgpkVA5OFRvzBQCRSKL0mwxvYDyLYfzHZYlB4J2Lb
d3qVnGDRo99W2mJnVlaBEzR+GB/KrNRBo4I4ERXyPgmGdCCbdtzvCtzDFNCBYNlNdkAi4bYpC8e4
glCHN7ZE+q2Y8sC+rrfEFs6OPns0AHZ06T4NkFd7W9NPzb+N1e+svlN7NZujz2sDNFzzloiaSP8z
XhUbzftShUcp3yjbIQemwj4Pw5W3QIIQF/+29RIjD5yCaDm6fqrDb0F/MiNjUQyvCIjPKybP1y2F
gAlRQZls5LR17rb7UV4k4Xn/qGAoxro8Z2ELc3f2VN6t5thY7TRlrun2q46cKmGtpCUuWn5UwvV8
uc9y3akYfP4TpyC1qXGd/Q2s9XsjLE2YFXqQobLYZVVk2UoeA8ax9/X3LLLi1LHynVHtQ6INy0ba
GCzPF1BGVa046haBiC6gKj6ZzC1jw6LvV91cJc+fJYN/O/V+2XW+XkLPj9Pcon8vmueqIpYQW59K
UHfBmCcY3ywW5aErHsMQMaAGKEO65JHbeJhcbQKb3sEZ6Ec2dqORu+VHoewPUCq9HMME/SikQREQ
36aI9WnpqVml7GVfjk1W65akb+arnRzMa96HvcW92+heqKPWSQWw8nUJhI94rRVxZL6Y38+A6xVa
qacc6Ppwd/+C/IL/Cdyu4cB9ZX5Tdi9HVnNoj0XylKaDXy6WT7BNtUjuil8/J+ZCMaybBJoZacZH
pPfUpvvcMUvOHFxhYakzbH4gaVyDQb5wvHtE8LPRLENW6mh1U7ZaazliP1LkkL1T29yOtrNlI8qz
+4IutWoUO4E9eNuHJ+GuNpMaFVqIaGWU6O4T7W0QuTu6yUwzGIQf0ikV46fmUQessfFuQdRU8Wma
42C4W6HrnNbecJMdw5xmkhjJYxvKmP49qW2aSl0zeBgHZTMHRl8pgBl3aLNmMzoxGvd98IxhAWNg
opKLQ/fws0n3SDm2M2uhrGiwgTbEXVXyn40K2GnUA3rXzA6LHbyzB4vNX3SOYPPjljxpDN9KCTXa
HONw47y8FMFVJv8hmWMRIFYxxOk6XSNVVvznLIu7LBUTb6DNEzw5p1KDyeoPdtD1tA2FkpSLqEtv
5/6bq198rHsUEzrZv1dyYlbJEZ/iHk60rZyb+FP3xM9oz55vFRhCoDW2hGz56kRXij38Ff6zF5U1
Op7acOqKnn+FDo9DaYwEON+rpzO4BLPsQubBTTyiTbgolQGQ4y01MzSX4ITt/V5jsRzxvcJC2yET
tv3SnqLVshulavXZhcGD0ghVEewvPpwLHFYGbDH7hZeJo9zUZVhlABRAFsAOZY4QliMGY0OeCx7s
Ba/n/frkOIWtFuScJAj9jzWrzzBamKpOmiERWW6dGOvINb/63lZ+aYQgBMB8mklBcH+uIBo5DULn
rKxFS3jbQrk9SeZ8nPjWgeAiqkW2/AGQDgTltLrXSLO2Rr0z4/FpeGllQmwuiqF7iswNH5uVEXAI
auORzxIKCPUkAb/q3O1OjCa2B5uxsMG2Ms0GvlkezPQtFegGXXmzDk7mdQANjNi5grisUvs7lKBD
pEc14x4W3trYZflSgD9AQFnZre8meub49aKgE7KHt/PiRCTU1c7/ZeNO/cd3vJsbLxVD/d2v2R4+
CS8Y1NP2FSjY8vUNKJDxagrqi3g3siI7EsNY+bRUl1Lf5pfOyud/LRefUfHI41iTUcJDVtv/OSTJ
UYOeTXGkxqOhOPVMKMJVKEWZDRKaybL99UcSwLEHI6eYvMsYA+YSDKtNBm6qH0I+nFy2GqWsQUat
hNilVy+PbfAHnmor0PW2bfyoHc7ykhx//8NOnAEhMcBDwyX+eaN0sYWEnJFfHrJAkF5V0pNfEmAg
1Siy4NSi6olCmrm3Ixq4NDPY2EnmyouX9dkisgDfvP3hxwyXj+i1vVwu6Xq0VRp364azVNxIgPVL
x0LmHJCpQw6ZInlN8YgbtnBvdI/6KWPApWNfS42eQPLjoguQvyIBxxETvTwpXYDJUQ+v1GenCgmq
ZyTS23O2tG9nG+Dp3001luJDQU+M1DsYcZQZDmr+cESjfVN9mXmV/y7CnsVIDyuI3rbHaa6io9BH
uLX8wzNahBjSqK0bBvnfaVjchPoPKFnwm4l1OkXD3VHprQgkKn5TDsOYM+8W+Wobv0K0XsvBavMw
Xb/c76TBZgqyr+yxfVkjzTriGpDWO+fQ9RnHUWRSMtboxUzRRGiG9oKGYtZvcFyp1Ihi3X6HygAx
ANbGMmiEZYD0igkHsGBtcdlvkKJNncJNbj49N8mD/L+e20X5fIZbuEnE8vP+/Bik7Ahm972yWHmK
nMPJlMa+VB+OfrQwK8DIxNKbtrnJG8bHjNfWx/NgFeGL09ekCh/rmdcxX2e+AedMlRoz98/hI7RL
WRTTham7Bm4QEERwIMBKKjHQ0qJ/4LhgxatShpayI9Q2VZ0wGNfAP/iGj3pNP+fGgkGIR/GkJPhd
VMp/ad6MCgADo/DTO1T6xXaxEIF8+n+0CpSHc/cRvpxSHwHZYvLQ/TxSdqusg809ar9D7619FmXE
64Ku2YjmT2UCqJ594eKdMLNX8980ReqkQrkukKkdDhJvpPOKzGHOBHF0OsWg4uWpjTH0nZCz/v2N
t6OZp3kGTWmbO4irqjoNrpRiiy43DZSTMyRyQ5uRnCQttN/9OD0JfPicfVem+Q5GXo4bV+/q5MIu
lemuN5gvp2L2Ea/lam0D0R5wc2XAVPBI81GbCA2kzrHzuRhlzUC8TwVWy8srbW941cdA/lpYJQ57
zCplO6k/1zjpe3TLlNkRFr0maHIVPUhrZrsCeSF+ds3Whcx6r6QkoLUROBagqHsh9wccQdA+I+8G
t0GQhH2WnRmOvmCa6ev3p8vweSiKaMNMwU95cGIZXwyrEQncxMjD5XwG/i8q8Oo+7aTZLIIqKD5H
EyMaL1fbC/J9nUhb7Wi7dIPrwgRkyk0TzwLmyJOJXxvIbAscAGIj70bLxuAeBuOYkhBP5dVFvpxO
nYSugymJFaXFDJanmZMFLiZVQocpCPVq/olrq/gm/dA1ML+bLqjOD9ov2eBBkB4iBUVD1Y+G2a58
a2TVqLzd/JSA/iU4sJ+XxgwceQsDp7+o6SclOeFUO+tqSsiXYN4wNibZHwI5jTvBHhMAImQy0JDR
YV01jp7GrItUMyGdCQnjanhFVUPMhtkqT48Q9TBDIyffregntUn4eqhU+IR2H9UTGIW2Kx3APbS4
zhUeDjh2hSCnzI1zCnqEmzm85rdm/AnXoS5B0xwACkdCm9ExpU0e+GpVoFFqMoFrAy94/8RfRP0q
NoelTwc7HDIyJMYulnrbCx6lCxrfIbF5G0wAqUgJ7RjbpPJYq8w4V+/GuIeQoNJ8wEUJ3J1/zxQc
0wDWYHCzD+aa6Xba58gRqeRE8CP/DkIK6RGCbayUspNPkP0rWPkLkRu3pQCsm6ziXBZepbqDjjPQ
P+b6h1nzFrIzETGm3i9Ia5tE2+MlXZi14mmD1NLTsH019Zz4EexwWyg8SsLyi16JaxLT6drlAgA9
Oi5FG2hcZNmtN1EZrt7b8OIJpwwWqXvx7VQ3VHhO9PzCmjiP21Onss6pjDCwr3IfU0yzRSbnLaZI
ZQsu5uIUdZmVG9Zco713OoZQ/EP5SG2l1mBArkGtqeu9FGqCsisGZMLFf9Q4s+LqfdHeF++AvH4t
lagOHWHZP2JniLbMFDk3rIfZ/VwWj+P35ajL9SSGY79g/IUe3d6l6u6/+EWYUN5Hq4UaQ6L8EchQ
g0vP4wI8zTzSn6o3ywflsDaOJHZyR6dzD33lADn+mwy+2gezhEe8ows5obRV1XYvcy3DiakSZS9P
KR9Q10vt0yAuT5z2zI6cnz3ck5becjL4HUg7FexPNvtJKBYp1JUIHrgUt3JHmiSb+qgELmVKRPmc
sIMWh3lpwoIEnkHQ2ZVzalLytKvpHRW4q5fHxbhi9bXNnmH+kUYQhcbOITozJ3vOKAowlWhXlGV/
F95ZeAcA/mEfGR7n/0kFlhObUWIyKH942xUdxCgOLngJZ5k5mU26WQ2HJI9wpiwoThcQ6nsLFAQZ
sxA3EipYvCJ+oJLlZOLtQj1+n7iy2/rroh1P0T5EY2dti1xJD356xN/13j1WQThUYQO2pfTmubNe
oPbQEuouKtDabYl4K6o3sihGs8oqkL2/fa0yVqObeBqVNOLoPiVdMp681IxVNcFK6JFetuDCBp5+
CiHIkwaGvZe73TMS0PFz+nM4eGxHS7uHBJeOx3fpNrSWA5/2VBti4lgJxpGBnFYvtwTyibz+fMAC
eFMmw0pz0JsNYn4A/8sclj9QyFiW+EKT/4+mpQTt5ZQhvCuL34UZP1f+6exklCM+RRXLka3nlOs8
WQRtNl5zcQ0vaULiNbs6GksiE2UmDDj1JqdqnjMEHhY46kaCBsR/sef2OSlo/dcF28tNdilxxwRP
tfwTRi/sHvQI7jwJ9sr+rImKfZLuf6UQB23U5kndymST4GLQigjmQ/t5Lm3sh42WJ1oKN+LEwBHN
uY976gm4HHF+pju6vqJR+twgGMwNNcL74hJP8vC242K1x90zV/j0rlbYo1XQ079qmwuUfSN50pkO
lbf1VPfnk6o21MTXYuxmIfw4HPau6rRaoet3/v/1kHgJlr5QFg1p568ilqXk7kp1RGbxfmi2TWmt
ePjDrMrBWDzFMIcmskVByRqGnE3a3TucI93etTzcr+wVyzGEXCVoIYQ2zyQFCVNSNVy6J/ievuMB
eVAZGHsqmeQO7s/LzDO9JURBrRV30C4AhQy5uQHks7PratzMv9QDTmlnPM2YZOC8ds5n1dyj+ovJ
o0PymiziXsWIBcJXzZNweqtoTCPvpW5cAAVUnjGHZMoc9ZWqtQShaUO0OD/Y4OdR3gyIGkRYtqRS
72hKzA+5SOSofJCS2wPP7/vpCOqnpKz3y7IQQW0mrTjbE60ak3cwRU8h6J7BEjGK5nua5jRP/HxY
CFeyEWmAvvQZNGhjEQzooJFj3+iImJ4EV8FWK+OLdK5iQFTDIHkheYmdUs4pl+rgYIpbr2UbSG7a
wPg07JhFhRIsCEjaisK0dugXDxcogugj2EPeJkKrT9x7+DriSxAV9VSub+svVCgwAFICss7o003z
bv2b2HW0Nb7jtZQ9Li7kQHKcGlWuoGwETCn8cIKDzvERhSYnt65FMl+5zUYazhWgOZ6QICs+YESZ
lMUeeQNgefsmRzvafReoIEhNUlFYK5unZ4J1TbuIrOFfMLt3WH5mTCeCkCnEZVBGWnpmuAFawsXH
vg1kPcZx1oKsOLIKyaMUtEbHU9eGwl3Df7Xuxgmqkvz0YfuHlW3cQ8RHYkCASpmLZn5+SunPBbFh
yOIQA/gpB6q2IrzPTpzodFajmIrnC4n+KSioqxWLODgZojtHuHG1mQ+EdH+AAoNuoyteNebNr2ml
V8rQUVrr6HMIayWiVE8QekKu6ZGigIx1M3QsqR8f6juqc5RDNFpJRdJCPLo45YhJ4HHomrrlX17x
22614QmfDX6pJqWBqgcv1wTm9MIj6Dq5l2pNsJRmdpaSDaZ9VaQ0Fe/lbyGNppaID9TF60zUjTFq
eV6DMdE4uXh5Fv6TxMgou6wKXRRcLdrfyAnX95naJfwZSlVsxrDLb9+HcXbYTEy7KmHTfmrQ67s6
sKfMeqWgHrgbWiXOt0ThXheNe9e+mgO0KlQOCqJK6HJ17YAIEF0E99JDJ+pWx4I/eDWCzt6t0uWR
eAP5ykfOqtUI8WWLW6lTR0SjshnDKgGhfEOyNNj7+Df18hfWwgSwGEaDAWyhrtu+HYQZN5f9KXTs
XWGyutTxh20teOlgsJ58mhOfy5GkV+Dqktp0d7jmkcfkLvvXbPQ7Qry5zQPsLzj78Z2I7Hedw2Rc
GmU/2THUscHwffgDHpVqhj9/Qzshd0pGnhZnaoEb3O5AacbG5BatrbkGG6Ei76HHml95d3sMa8md
QAO3ku/X6XCr9kK8e0wzq58hDAi1K1q0iJRexytXTq4dwLRRsAATLwp1cIySpwuP0+N5hHE+TrA9
lOcK4kGdMrtTu0HXhMm4VQ8FKn088WvRaHS96xC0suirq/uN2ynTvEd2kbvoICJympfOG8/FqIYB
HKkteKwKXecapgbCFzgZHYNANTvi5Z8/XfP70t8Cr8lZqEAw8JQAiERz1ygl2lpERNdoYG6kpq5p
VU4ryPg6bstvrvGXnh3LEXo53kHIVkGcyEMF0Tea3SgjzKeNJv75VmiPPtuxeJXty7aq1SzJNmIG
ANqKjnAnepV9TLotJWgGBYsJGyMCiYvA5sXcRVrklEs9W0gZ+kJ6sUlUoBIg8AMiYaor6sj5t2On
TclFUB134IR0TEm2fzzZzvHDdCdcsMnIXPX2quDh0OIqq2SG3peqcDe5Y2Vcu08YcmjLeXuPJmMD
eR+wZ4exrRM3qS5NGohdb4Py6zBzoN/lcl5+7kcVjjUWd5yuy5Ivt/1mGAd13A4IyY/vF9N0ucND
ClyROhqtOa/OIu2jp/3R/BSntNA7WpzLL3hW6szaCkNZFP2ICoAqwrim11NR7RI6O4K/dT3npjsZ
6fKTKKoW3V/xXqa7XiCjSKpgMx9FlrFepPN0Iza/9IcKI9nqQBl+U+KbIUMQVrEgYrCW3acJITNl
hT63RhdOx2uvOwn0/1IaXx/MEDDrnDEThIcWQD4WbAHWuu+fRSdJK8Xs63sHL5VQ0/tGWfSX36hw
yg6ni4P+/MJjlc1dKjiZAO2fiDn3O46DuKDwMWApfD6wClPStOLBLXp3OTP7RL4pU2LQj1b7W57X
vU6iKCu3O4GytPpFx6JJik0YodJ/RRbx3bgyO0MKT2u9Dpo4i3s2NWKXOIPtH8ZJ3hJx9MO6YYmp
ajM1WFKm+JbfkHBAwLiO8Jl1cGo6/VqxozhP/dYg7JJMPIDIuF24ou3E1l9VOQ2WTMv4Mnoivw/w
aHzv+B1WE21fn7ytkv38lpuVaux6FEmHAH0PX5n3ohH59k0zj3MAhKXPWJeiywMD5wLEPCsq/lFl
hdPs7Ni/RoEUZSsdaqMZ/x2Ar1/uL6BGrxOX8HxvN32SEnC1DCja+rONAsCkLyVBYJ+qabEKhlC+
8m+eIud2VZAZ1MKSh/upR9hZYd14HZqIOYR+pwQhz7ZyCnS5BCQ939Zb8DxM//Wi1qnaaZNaoHun
xZbQbQMfRNxkTPdbQfcXcASDr/+1gpL8wtDQd1qfNY7+gzBqK6bkd+Mae3c8
`pragma protect end_protected
