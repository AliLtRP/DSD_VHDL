// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
GUJQCEvkR9UlE/UFbfLysFMFaGYdMzewbG5jo9bSOg7lI2dSFG8gtejvEqVx9lo2/woyuC59mmDA
Lef56tC1BH/J8sXOK12raPRAcMVsYwaT/Dho3Eho/C4pFXeVuI1MBCjqJ0xi0YO510f/H9sKpdO8
/veGFXTFTdASvlPhD0Irjko4uKcX1yVqi1Ld/eTwHZRkotJp8QNjonxtI+mAyDLB7eIQ2fcbdNvT
we9EFh/WpyVUvvPYtpxtfHtJLtxlUB7jRvir0m2r9C5rVAvPi15OzHJ88RBKPP4AI+copjHfr0C2
Hpp3/gdttd2CkK/RniDYomX8y4wwSlRcs2CRIw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
iQU1mJF6ifeXZ1MysyoYPtYcZNfnBstAqjAG7j/NXI7HE1WeF4mcWV90NDZBauMPFxS/UP6tJG2D
c3ug7PAIthz7ubXBcf4wOVlGWTYSHHAk8S44mQl2kh3wcrDYigLaVib/S0937c0ZQsjA9d038T6I
FBjJ/eTb5yyJhqNdZpFYVErNH8UwPl3PcAQpfses8lsFSum75h6ASR6bTXjtMMZutEjIPdmzIESv
bkm4XTDvoHHKF9COzCbjW/c3xZSQKf7xBuhfRvwql0ciXT8Ktwh5XUXZlYn59lARUFRtSH8UFnVl
k7QwN95tKQ916Rbxt84uWJ0SYSzBuCebM9qdZ9JdpkhMIumm6rqroa9UkK/jDlPf1yQmF3uCmRVf
J2E7MZebNOCrbpX3um1YIU9KeCC9DHw/q7ZppUvi7vEeNmJqqa5nOU5460bhKA8C8AFpjP1rt6cy
tTTxsZlGWMHag4XUBgTdhNMFvt8bWwrDa8Hh/EZ0TpeD7lkUwDd/8SzCj4LP9bBsU+XOMGaJAha4
7iEjTnK8daoXNVwISpQH4hVu7TdDUC3kO0v7R+9p+cO2/HZbS+mrUOGBz6yR44JGVx9IlgjdTOBx
Ujlqye2Ah+EPpEkLQe1PqlmUo+n0hSWe/JObUaiFrFdZm5tavNt5zNbOMry1HE09/tvnG41gDbEx
SuXNgVp73eLSPQKuIrAwtf12PtuxBGpAqLWf1vypqnTzlYryUZ5OsG2m5BTTsRYhF5gg7XBypiLA
geelDu7D7CzD615sGuYdwQ23jISDHoG1755zpkM6qgmcAxmaJz/FhTOSg65mbkk4BNusoJA/U156
KufLj7o//3abl/OKdlG0cV6FcCHEypED8vMueJJjPQSPfm9qQTx1435TehGh5WB89YuIoacRTwlc
1SfUkkd71kUXclVeVabTcEh4L/dD7TN1erosWaDt2thouQvFSj+gWVeCsLRaarUkMf9zWUrph+qz
zJc6AM5ElMwROGprpju2rFEYcQN3xL0vP1LCSwglpqpF3LkL5/x/WNylTO5a03h/Tx5K6SLFCg8y
8YZUEzE7gmRs2t6H+F1/vpIaJrbzi00m4uoirqgrpjdNyydcKu5/QQylwRvFCqV198jgn0idt6Hs
zz/kk9TSyYGtaPSnUMHR0StFlXCnBn91yaVGE8b17deplw2nLK9XyqmzsIljf5ere+AxL8ICZR7i
hAub0VDcSPIHhGjW1TYhJ2zWjc29kCx6viILdd8eGWH412fdlKcZiY/bt6BN/SX0PKFB80rGRd8w
FHc1mT28upw1g4rqL1EYUIDLMbFpB4lgIgmyWVxk+W9KMeCV3jH7wSstmQLjv58YMATVCeRyAH+r
Jey3YkmmIgZjspOhOfo04c9Fv7bpG9uwrvxQ70YMfVzdr2aW/+ezNnf28vZdW8C5+hB9hnIBZ7Kc
PqZgxxmvfwyTQtYJLRz755Zj/2qdN9tRwH3/UfRGPK9dSLifCkkPbue4GSAhFt9962BbkCZdTIsx
NgDr2A6jc9yPjIJZkZ6O9iTtWKJJtoXGhbLhIWqJl2jXTvNCXIlalGxHV8Lu2Jlv9fhZoHq6TlpN
KJ6lHWD6LLX2B/tTrijCPX2MJO508M7nWCsKI1sEI4DTH60/s9y4pyLRc+7Lcew0dbhjAfgG5Aez
P6CU6/HNf2yVO83u8H3b0iLMTzhBbocyyt4zzZ/SYTd9bU+BmQSSbsuttnjOlNZZLrRwOTTnx3ey
W5vj6D2au22YmlJKw3Ey8MqXBIq0bf4ksZnfYZJF96W2LdMqZMynKGKiX74ztBtLwIPtlBqjKbSh
2FFXvm+pnO5ifjwsdPSglqnuRrACNL8CFvfaopoZZ+k9v4YKkBEn0NWmBHcGnwayfurXPGpdCEgb
piIbizrxNf/NLmvhL6V+/XbnfEdAPH64rRWQ3kcryVc6/Ooix2IrylcTWpC/tG30C6aOdkp1ATr+
kzFyA/equJlFWm/0klhiqx/gZK/09dAaut7h7SFMnMPFJFl8j8mI/9VxywYaOmuFZOLgevfquuS3
XkjoWApRBadvFfp6DRmBIDXml1Td8DeiES9wz2bE2mWwddpnIcYgByzRFUBwcuD0F/WziFf6IlTo
qdG9Zow9plZRuOf/fQemxtdOn7Ibm5zsFVqqDUVdjtPODuXbYw25hhYZBV514IUJka/cZiETzGnu
4PK1fTg0bK05QOfB3Zhxg5NcPIJS+Z5xbH+pskALs4DUBMbp/nAdYxGZit0jQ/rD84iJXtMucqx9
pyixB0wdpVTKm5MSBDKLk477cBLMnD0G/5DM9uIn/QLIjXoBehr/1jZ8TZaegL8iJiVg1oD66IPB
W2sUItJYTahDu4gPZuemCJbC+jxSHB9XRh0y8qdb8zjzyDAIJCT5GQpyh3Dzg2LZ6xPZg/+tvYpO
3iTryXzzxkKDI581qmWRyI4Ln+cc/pYma6Wu2OM5eRh1k7qODaaO3OdUJOLD6VSNuoTUp/7uY0nV
rAN14gJxNMggRsRyDqD3mDaRnZvCrK/7VoN5vlsF/mctzb8/nhb2q1Q8dkkCVuuBf/pusiyG3yCe
ytnHbQkN0CMS91hDemvDbIE1+xuM/UaURAsoF7SRfgI9HHHrPsxsSg0SHawNw56A2F7yjVjyvX9m
epv9W7/dBmk1259j3yUDCSi2LBxPhkP9cOu5MTmogwTLZMVyvDjhAAFpq/7eps424bNDGs7UenSn
gSFUBH6+hP1H0TDZ/9em/f62Gv2h8WPyaO9O/+7ExkLyM3Y5t7Ug9tFfT+ffSMFGBUIYnxx7Zppe
WElYZbpUDi1QOEV/UwV2E8XCM+HM/3jneqbAblAVLgzhdVTqJJjoRvEqrSexvOdm/fHSg4+XcibZ
UZbsvaobQLfLq2jgeG1JmESQWXp4e6gh7lrBZF/RTj1eQHaXq7PnGgtlWBCA1j35aTW97SDc9tsl
SD/IwBCZVXaZ+QLxFDvf0Q+mI5A6+Qfq9pfrsaHvO1cDgaTxQf3VNnYaNL5J4ydihT7eJ7tuLrPf
gfnd0LR/UoKXhbsTEbeAmSx4wllwgbTgAjXaQV0VdMVeHxXMwqF6/7qwU5jY2oV3tNWSbQy5DZqM
BQggMF42zs8bh2G0g6fJyM6+HdZUDd3TrAF4Y29/z3mZSurOw58XfdPFuAoagMQCYVY9+y8/Is5F
xyM4p0y+Y8GO66Y0//gugtMcGKFmPuoan7jfnXvSi6rVWC1ZIhdCnuEDBK6UGcB8A6NVC/tWg4zq
M5kbWJ1vv3ED4vaqJvp8hSyyTAmfMjJwfSluQDnxMpJsYyNAONx/5o3KjVehEq7vMl9HF4PCUAzk
LeiNf6JhUSnYbDvy4AjHaeBooUkb/OiR8BKlkrp5cmBHBISyCAz3bPbtiApwGWJAxgGdwoXk4dDx
EVo3WmAywLhrtfZRFLqa0hqrbFgQ27NqXD3R7kc3WuOge1IiIBt1OjOkoiOHh6WjY9VQ5FX+5d1o
C4WntFrWe3QT9DRgpcXMBMo3dxngsJsnpWq9HVkTd4v6C5NMgGJ+mROd91tI86efV71ghT8uFi2z
07cSzs7942cleh+5tEGYiTVsZbLMWJPnEWcjQ/coodc2Z4yb3qNpxgKNDGfsNv+tQsz7vQGNZbQp
9XxB6bxodBv3QnpE1AluvPBM7yE4vTt0pZdSg6gdTN/UPBeUxEM+MHhjFYJLztOctX5+5D/9i/hk
b0yR4wE+vv5FgegOm2PPJCC/nEVAzX5zFAzUBy9GX8otX61BKEoPPb+QfGjGVXnzhx2lXRVFJTWX
NpjVVY0Y9vKgTWuWcvyxJoWtYa9qRILJFSedMkucOJ40/IGp5fA+QLfXmq6v1+dqO5ujS9zHV5fN
699CADinC/Q5EjLe9u0/J0PHCEQK4aew7hxtX1pBDnXSf8u+SZqKdpVpArsW/8aKt9EEPI4F6fuq
rcO9DaIqH4X9/WuoaYkhn5vlA106sLl846qydhQdtPL8Z1va2qeo0DK3puBWqmIQNdwpfrFJTIKU
uBgdmcQ5lUBN1tE2kzlhUZ54EFcrc1Ld2A0BiyGMsCoeKFDpGXhk1cxkHww8GWyDrQ1RSiPJYHQ7
YCIFQkmZdKpYl99oL7jx3GLEm7YZX7rW2hJHkx4NSOqsxzjkhkfl0m1VPuhBqaUqhkYe0ZvrYNFr
ueNASJop1ROZIdMXbn7Xr9o=
`pragma protect end_protected
