// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dxQSp1vmPAx8+1gzQv0dznE3c33xxTdpJMOWhkNugup9xtJr8ra/xiZa4vlavKRB
xaDhQP6cukV2IxBdmSojHk5hXo2I/cWZpe4b1etJp87OL/fYCTJUWCK/zDHLWuMm
UDZ4cydaa/DB7Boh2mka2hdqW1/9CV4F/HYfmtu5jEI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
lKJhFNR3AlZAJ1s3/XGyMAzOtJXb9EnJtea39tdlcc/9CAi37yYDKPB6hg+m4I12
NDEm9joHOSSe0FTUio2oVgQXUnWb2wXAet6eV1PVYC6rOn7ILVH8K6+lUI/Ox/H1
pZVteQ4axIVZXhMPAWuwlgf/43uDso/ftEkLhv+xO9laATIfVf0UGCBCbf9xK2f1
r6urXAcNufGW+w+5pwe4ff/3DTgyXSkZBadq3y2DYrUBc2hSv/u9gJMt0pG8bVP6
wsRS2cqrQdLBvO50heKsnlDn4cuTuecUr0MziqQsAapq6JRlzFGjCwarMt0blL/q
iUPmnSNbBuO5cT/YftseH7vqESr4i+3BFAG3nFWG4AnsUVWcndfBghLelVcapEAh
7o29xj1+dLbwC1JliHGNrouzWeLHDCmlbhg33leCz4lOpsP/Aq1IWBoN3+MKfWp8
B225mvjXTpBb8B5mssujbhNLSGU3qQFYF2d6QIZAWwkRk5rCTkrvLl0xKh+RThwn
Qg2hg2DfaQYSurWzY16EIlkW+pkXUKlfygm+LL1NRnI2VbIBMTEK6m2nAjWs8gGO
ASxj7mcoNDCUkhD8exXO0NELJTZhrJ+uVPlF7uv6DzvDpE2IOCyAUD3wqtp/dx3B
4hLjoQKWQFn0tX+YBHnqobEPRDq0HoqKrLhFrHg2jlJFAL+KSwxZFGnhYIEQ8qj2
LlflKmspPeYnbIn3lThiXjzkXSACtFMKdlS7MLsQUajOpmlK+/5u0l95FjMcbBK+
AucVkYBjeBeVfAYA6x2PKsAJKlUFejoAjKq1GlpTqmqlGMLridapa94dIGTja1pc
hdjMbgXMijr/gB6NezliUloR/CRLXTCBtPxz2iAlDvl+Zpq1dOg+6cJxrNNxh6Ie
4jYcOwX7WkZGFbOj8v2ki6Osp4qbmC2ZNiGyeqyBnIUnAQg1AYGkGSP8NjBF+Orj
B4afaC+mKk8QwXKTzt+52Z4dHO2Z5iywaKDvlJ/M03sNeWjIMm8IGTlURwfSlffP
xc1qv9UP2kz/S6Sxxo0NJWzVV47y4Rhc7V9QHVwI+Z/7Xiweun53wTypKYTpu1fx
yamw0bsgk5FzmMccQftVSRue1aDalGRZbQuT+a9QhfAJRgMDccqKJor7lN4Lp3wp
fAjcjgxqmrACPGIuhBQqrSQ7Z2YIjET6ICyx7ub+45Ghu4UJGHZcF0uWtp7uKnzC
2ZYdEwzUa4smduNOqfIzRFvNHwLggRtDXerGnSIYV8CQJRojvkHNE6boORBKST7t
MWtHMRclDHYWOTPR5ww/V0PeMA0vcvkQnxCJJbf17JaPoO6JyvmV/TOdDPzm2va7
jo+4qqKrin/LTve+bY5dG+6KbGaLq0GtU7RtlfVyUTXS3VVEIy3lwtlVlsdtxtqA
O3sv1yvfuw9URbcFDwzNQkbfbwrLuv/YSgMJT1aMJ3NsLOnlUW+HKW34lzVvr5RD
wN7FJg5pcvf/JLzOCne7sTxJ720Pz21W5gUP+AnTfmhN1IE1+MLqtuIhNCU6YyGM
YnPQPhHMzuY9xciIBL1EJMha3docm2BQ4sWPMmYFOMIUBs4V/uAS1QT4rIAViUH6
nrJbFvUNx1tAkoB5FRNEsfGUZNUBkIvUB1KNQB5vln/uGTHbx264IcX07Mh6oeAB
UKm5TKE8XDdL/LrIedYnylo3y6yXeYd+8h19JFa8joAx95fdtreuEKOpqett0AXX
kYQOlsglqg9TMknkqhdd9d3RXwRP47n72JFNRzzD7SOmcEZoX/CQraQNVxcSU6mU
EJ/fyR2djUalv7BY3jzzBY1RV13Jg8fC/zBzCH+dQPWgxJyq3BnzenXaPTKV4vsO
/CjGoYR7RGA1MUIgAnelYZviaG0KJlczARUTSPjSI69uBVZ1jrPLv2Dd6yPpepk/
mqm+zJ17tWW4RHoC4r+LJDnkbD3yhV6aXiyjI4ENrCv+rPzR06ul4DvMGU6uob7w
ElyKsmcCNhFEb7N+arvDtBF+ILzzcnplU4crHJNhCBWwKBH1gD2s9kDqylh0qOKg
BlLx5bve7+8Sv9dXM1yqxku75SN8ABgVEIRriRJYaTm+RpDnsbnUX083PAUkVF9H
5or0kT67IQflFuE1MT9tw7wXGfeRz9YV8UE6QJ810KmI+nDrgMOfMHkz1VsF3dbm
ELODYMNx0b6M83NryWd/UMemZlchfEhr6zUcniFBI0dl8OyxB3VNV/dvYVehjJ2I
4rELWnbOF+xDis4hECFgXaktSBJdDT/OFoEg17ua3GtbcZvL7Itcpbonmn/WJODI
NUW60hRduShRcqkG0lymtUaH3Gs2ay8aXZ857jdy86VcEOeWRID0QyGQlx6U4xli
7C+lV+Mnr567mBpuauAX0bz17IH8boi5AYDtcx793W4lndCJe4ajmSdFXld+RfSF
2sJACDMEZXi0kuH7PH/dLAOIRMfjH0eSjcy8l285SNk45XBb3sRMgvFpawy1Dx9y
jEgHFaIXA1zqXH8T0codbwrLfydAEq8dzZbWQr6M4KqS3ApKWzLm9E+sD8G/Y9Gn
5Dz6soWe+EKd6OtTBGzURb/uNgjiI6NMN8o2IiNx/dwlml9xaScn+tsUlgIfly+b
7U4DYQoDxOvxwgM+/g+kwLi5d3m0+CjRiRSXuRp6HSYCGpaW2f29Ko7qQuN3aqUU
v7bKtqOyab/oKHcOvqMx9wvlYXe2zg2KeyXh90Lcjr8Hh9kGTSpPqWK4VeE0h0BG
BZcmvZMx19M/8Fwsauw43t7K0+rDVR+Gy6IbiAPTaS02x4DdN/g+b61xHzKS3ayl
Wj0mTHNnK1E1V4lZUqVlK8n6nzH2olscDynSZiKDH1F0eZeztu3ZdD6KbmDWefiM
j+fBHSjKkJdNp3Dq80/yFtpLF7q+cKYrYAujY884qgNjAOJK/HizzU5m+sjpZOB8
KI3xOg9jHy+gXBGt4jzXRRlSJKr5lIzK7OP3pgPACHoAgvwBbGbXqtR/+AGVcyHY
CkoBH7IwHfFPWrjvdf4s6CCbdSV8L86rzlXn1g6s87CuhJxVjD6a1ML8ZF31wiVe
BnDamV4rWDsGHIZZiBo6NP3Yh00eQjG0JHfZITxlg3pWcQmFPoAjBfT4IXBc95BK
B0SN2TZhNfhBwW0xjs0/SxtCTRApWmxNpU4LWUKI7fYEyw2BzOgRSZlkB+rXuKa6
5MmND6f6kmGq8Y6rh9h7KNtfDFWiccIZ7GE9cbLN1kj8NTnNWrluykImsZp8//S1
4IVIB9ucgmgr0zunATwMzZQpvvwgMujYl/Mo7Of/CDOPlY2sP/cIooU7TXWyurNd
mCorndOWPtlAXCUrFbtCMq0N26bP5DvnNY+248JtXO3VVSNxvSyQ9Coqww8KKlZ/
PChakb3oc0raPfwjzjuids3KRmSdCIdI0CVoyNmTgxOpLr2Ylb6c42NphXwGxuuP
gKJQdaymSRr8psDVkT4Bmtr8IbEZc2/IfJ2BQxHDTVSInGRS63Oscfx0QNpZOTUc
C59KddTH+312FPXIAVFytS84SW64iNLplWtRWdmCPccAqoHcqrb18QjVrtcxX4B6
S1Ag7G41rPFiVwswNtbIDYnIdLD5nwB/73WTAd7xbVyqNCa3QVAv6PPHBh+2C7Zn
M8lP8u6eTQVf1EYBCs6b061kHzveZPfp2a39uKhfZ/K1WlATyIBN2k6SP3EGNwxD
K1t2dT/8y6vyUHY8AQ21ViQcZp88DUaj7vKxujPZo0bhNcdEzmDQONrLCWIj+XUi
CSn+yYWnw698aeNeyHyPLmldHQXDGAgqMafZWYKYSReacbk/6CS3IwL/+H9mC670
gDgdQM7tymQxTQN1xcCtnHVEoX1bWdMvMuMD52yWHK06v3/i91BLfK3qgxLWBYlL
wcS6+SjyCkhCPPaNBJ9B1rN0YFyrj/gYltuouzTxhmNUnxS6EW7HYhefwp0acuf8
uU9Bh30c8NbNXfriqwxiCowdCr5Ssmhc6woswJ761w8rdQ8XSn4QyxyBOH4iP/DD
Q0iU9mIipSVXiLVcG0nRTG/SyqQUUoF6T1QsZJqVikG8ltLkcERI52zll5IdFd3E
hzVMJ7bQVcTOXbrHDZZE177qGP6DkKOUObfjZMJsbjCgMdOZpms3DM8WHOSzEPHd
G0SR3VXboI7dU9El3/xYqlaqAtozRwB7Mj1UuC6AHrtL3Vsgz1DYLCMpavPVPiaD
DbwghSoFjzUzJ4/7L4oBCQyDS4skmhuYMxgH18+2fB2S2T+wbNYTMrHeeZbWsfyM
muVjf3SInE2tpqlnUvtdEZDWwRAjEDHgPc6xFSbpoNsBS9lldLLWU/KT4+5mYtfp
0h/U9W+mlNycXMbS8Vyi+r6N09FDI3CKf/WD34aXvTtuUXh4GYXzoFSl0u4fdVxg
paExOf/z0ySbreQns4xQKspLSbC6jW8fpVBlhtsXp7cRWilFTeAVDWTJ5iTDmnJm
WDQH4LF4kUnJtZA5K/SuluH46WXzf4BuDwOV+ZIhwY3IpiZVnj2Gdx8XgVd/BvDU
gV7gQpycKCIF9V6QHvyxjJaiPzQtNnL+V5wj69t8g10CzJMf3lPieD581j4Mlg7b
/wkYyNnvFHPn5o0Yyt14WYlqZSKbmiEdIVel0g59gmWhydHlXmGMN62PD2LCai03
QOsT20juHRQ9yTBAI9na9spGphw1bgfg7vDUawVdoa+5mO+F/3sa3lICQg9/rVLM
YiZytZcZKjjs6Y+HCwXUha7/gIRLaLg4xbg6x627u+snQC3maiNp30DhvHz4UHoz
4vT4ACa2I6kcaxvxays0DMjOlvn4IZbKNQAEokW0hiZOfk9mWhDbj9ib+iV548b5
eTsNuozXdvDZqGW3K7ZIDY40AuZXeUe2oaJhm1KEEqOW6dGKpkhxaWjvdbjoC7g+
+Ih8AkJ2jnu2kpRnCvaNdtm9PKAGboqVXe5eof/OHShAwQqvzPYRvknWt6HbIeAe
B9rYUW4etEICw38QNiwMphFSahYf5fdse1/px+Vuv7evoS4yHBE/3OJEjNKEzsZs
peEqgQJI+yzyZwcSPfjxfp/lf8mlrzgUTzEZdSzknLF4J/Qr3YeElkQOkvdIEI1F
teb7JtG5gRLHrzVWlC2cKiApINiHEg2971uC1dJMDve/DMcbRdAVi5JNtM8if2gO
bmn/gbzZGKf2D+dCLCjj4A74apFgJywwMh0+yYbD84DbS9n5WTjzWDLbpKaqMQ8C
NkCdz8/ZpWTe5/UuJ7+Iz8me5DjD7iyOPgz1DvecxEc8labh/hItCZicrtVWLWva
sBQtLkWTNkdwUZGg36QrMI7OP/6Hsti0Kn7uZnUJeINCw5MUbQRQZ2yZ19NNZQzj
cjA2bCHiQdxUDOotkbU3EnbCUR1c7uejSu6wf6lbW+0q6J2AGf/hTKXXUh3jaL2r
NttPyX8xy/3NOTh7KIUIzvLYkDCk1FYGHuDqx4TTasAYjT/ilYTibQchTu4X1Enq
Q9wIUOfpfpa00etdU3lk87XwCa/AHw+ZBMq+y4fxIst0PCVbFc3YKOZRHcnTZp6C
EIAjgYelXgVl8Ov0e/5S94TO2YtkPSekuVHqYjKOlHcRWyUB70T1Ovuh5HmRk5lM
pdrpXsWV5qfu6KtX7vRtGmmMRgL3aZ6EOe3NtBtX8ycWjMsgwjdbg0HrLADjbQNo
eIfuKtCGzpWyLU5FWZoDGeISh1zhTZYhgBFlOB1qSR9qqWMCQFl6aw522IKbBH2j
5m3BCJ+ccrXSYZ/xjcCJxp2jn8vuoYLwQaSuPmj6SvDgj8jALUbgDkLyzFu8AGcO
/VPYjhg50L4k/QveW+bcHuBAlR0R6UnP6/0lffa3anKqxy3OmQaka1br7n/jBM2x
9p+4qkyXUtoGMmAn6s5SjQSlnBJtXFC2pdGETZKDuDTsoRDze6TEzNIZsDNaspVX
2s7YFXSz20iBjPmC5tjGEkgUG5b5gFbvBEcMErmmI7E6q5XSOVtJVOztFxH5ljfV
nTbY9kM2dSsQbwKhu9jFkGvQO9KYXRtafa0qUQqjI7b6dXZspCOnAoMFd4InTnaE
PJAWUJMFUTkpP6+mhecW4OPyylOmL94O9zQEQyivdWDzUfwEewmyvJHSi1E4ASmf
DeNTRbVDtyZNB+xmBPN0tWHYCqqjXOCIF/A3gZOcsJBynZ8PCEYB8k6cFE+tIuKi
XRDnR04glVUz8pmiL5jPRzaseh03rT+zflIT6DLyrc6NxjCibr/4x8LkVcleV+xI
V5hccS+qMZKWoB15W9B9AFMLQ4ioBPhYKjgMuhd8iq7sV5/g+zCMKyZ4LU22QryG
N2Setgm8DaEOvu8bF+Bfar3OO+jVKqTka0nQ5NVX9unsVztZlkRZe2czUaMMN6tU
2KwmQAMOaHzp0hsP0MdbcaswM6sZQEO3B7W8srgpk7kwOgosvJ+qPFCc0g0ZYrr2
rxPfm+N5KkJpKwYw+l9zSs137nsA2bjloyC8xkWFg1YuZ+VFFBFu49cNyRZNDGL3
uKtcD6LlzUKAwPOhK3gNeGF/bwrGOaGGeHZEHqi7xZCvOtDt4Ycw4Of9mo4X+yjy
QFf41NcV6+3cAs0BhciWRkC3Sp+MdUK41KP5LwYl3U3elx6cqZG0V7mzH+hXAaC7
Nr8/xHZBqt/LaBIy3Lhnk/BPriugEZ8MUAQih0g1mtw5Y94mz5/Ys2mPsr9jMmN/
b8czVvelRn18UHkPgxUwbOs+dzRq1RfnIqDYhQykJi8JkNzwvuPw9gZIWeZ6P2vT
ePp9+uiDTO7lmEtW74eUcGpCKTY7W+/eSf0kmKhAnrzbaFiTfkbsZvpCgZMHRbUQ
Mmy7WS+LDJmQwCIqF6VwA3Np6Z1oZsX6P5SVwUzLKjBzKgHz6TgRNIHni0BwK+J4
qJaPZVqr+4ukdEBng6ma9+HSzgL3SOW3SmgT8ehoHj+ZfVCABXkjQX/N17zracZh
fCDUuzljuMx8JTSxmahqp6t2IdCp0jcJ6T9C7pI8rkHjkIR45yjKypwm6nul47Dg
Pbzj5CB0OTnEOIpxg22w5KCudXThT8UNJFVW0Xp1usOAJxC3iDAYYOgXD58uDvx8
51gLiY2+tR2M2xtzRcDnSP4+Cx0K/DNeUacUvQJTnQuLfeBp9cvIKVNpMG6Q3qGz
Zgm+4fOYnKpocVBNGaeebh15y7iDm5qy9YXhm58nw8HMLWY529ugJdql3B/65ln1
Vh589mnV5LxYlDcGgye3JAUhnRN+re47KvpT+w3IzOw4UhIkhzE4r/JjH04W3GaE
+e3cVoWzMkhj7iFeigP3osdedpn1JWFHZ7M9Hy1Lfs7hQodatp01XXVDjXJd8Y6O
DY8cEdXfljjKIWNau+pQl0dYbAn9wXEa8A23WQ8ANTUXtuQw02+9GbJ5/U4y/QA2
kQBi3TQiIWNJG+umvyzfWWnN7OzbAnK+jwdWTxn96rc=
`pragma protect end_protected
