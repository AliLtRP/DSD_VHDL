// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o0u/UtuEhE/oyQ+Ci+wWdn+4WOro95jF8/dlEuiy68FKxOe/S/VzKgGqNWQFmUCO
eCLTJ6Qkonkbcn4ckrhw6YTzkbiVvACvhJi61kg4iWRmaQAdV09CpXyMT/O57sGb
YzzBPc5nxSmgjp85h/snWvSE4qbBEWaHcRUS2P6S92o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7616)
OrjjkLieV+xRNMa+ONIyQ1yGLtLHQQ4UI8ezicbZG8YTiuibFQ/l+tK/pssfHxws
JRI8KbdgvxE68XMXUpz3Ctdv7zogSxiu7XyTxdH5pr/jE5IV5jJ7MWglfkdavaID
F4h/RYLZ7ZnrlD7Vk89xYbxedgkhTYS6UfaLxLxErwLZ0w1xtHgcDhNrcvBxMy0q
M4c9LpkDQ5sD0KAkSAAoeh7vQvTjOsevJoHGjmQgE6JpACaiOFQK/XMf/YHFsu0y
4a/zRmUEXWUMmE3N9BGxjC0t84i/Ns1qwX265prkrWdzbC02nkKQffD3bTj6107y
RG2qL3X9U2t9W9ByV1Iwm5a8H8XQtN8OFcFibIxXJ6hs2yxBMQlIaRmZ+iNlIuln
X40xA6LZwbzyXc0ygXp2axIvMSfijeTqHyjz7rqn3tie84vcX3KZ9wtlOyLPBOj+
5E4Uhz6ZZvF+sx7Pyy9bMpHqrz0weYriZO1tqd+JluqCb6kyrTbbZeCWxOepJShC
PWqJ3eJqevU7dK8SmIV7Do0eHbuRELqVhm62/I2asYFo3ijFoc7JqUxHeewb64l9
vsE3/S2pMd8rzoWBp3JYnYEvosbyhSGh8Xm1RzcZT9HSArzDSZ77QOX/2kJoy1sz
R/N+GTdNyIGRa6awvdP4+89PiUq9P2cRTYSn1BHbUM7jo8+sX8AACMLWcE5GA55+
1XvVE3CJ+X8K68L5+VFNLd9MIBwoOXo1k0u2aRBXHj6qPT9hn9Y8t0US4APEZuVa
VuYBpNAV0rB7epHPbqAt5V1Ot+xCm0SBARMW1v784mGDLF4CRhUPNuJ+b8LHMY+A
7gdi6t4T7tGZ7QpqGtmPg9/QlRrdzOvJzK0NrVUerXzLQKgC35AxG7XIBHLJSFZw
QMS6Y4Gjen7gVHYZtVbxZ8QIYchBPvtmKP6UF+vYR4JNsxF6GVLBgOo2EDWzGGCa
ZvdTZDqg7eAq6ReITjyrJhexdCWNgNjwb8KIZrVoje5z/OgARnfJBA3j5lqCeXeU
ge4Ocr4+hr79PZkQgQg37ooYeTSm48IJH3wujXv1sVpUA0Af2eEPdgw7bVCO1oB0
F1ynoQo5vJkXwPeWdaXohu3CbTJgGcr+JQbzR6lCbMmxxhhMZqgVEFz0sui63QTD
TCTUeZt5CHUhA1J+jkEQAtl3038VStArXY5eLZq2TWJeQqsHXQ3AraThnJf9W+4m
qxY+2YkY/ESYiQ+4SOLk6JnJeInVHl7yUwUTsEgFYkq7XDCvPfO+tJfHda/v3akK
rOQtyXfzamLDpmdbfdPTK0pIRQqPf+FGtbYkTWghiNg6p2qzy1h4xNP/1PYQNIlm
PxfB6MqFIAkhNzptLwrXlFDnoEfYN3f1mnP84zuavoaGC5hzPcJuDUvEivDcbyxF
gQqBTYO+zdZZIk0pIv0cfePehWghtq96lmi3dYmjI2KUdH1d+3+CsQOwh+UxEa32
rQ+NHFGnRdASnPmvy7ie98AGRzwtnSYk7rdvmIZReaGK4VaPuR3a3r9MwtcPjUkP
TpkHqUHm10gJw9eXegzRkXFjQt6hzBmLRM6CyYgNmuOGajik2GqnFtV+n9GiBFJz
xlWQtzWlMrwF6eBzAfYLRMNqsCiyWMPh4b1RdCgdaU+0EC1KNPluiRmhyK53lzM7
sjLYWirAe2/X6e5L0wALaG0ZAnGdIrQ+AeO+5lpsBeTukyKZGAh/zUyVQmT03lyb
ny0DWBO9qec4E5LeTAw8gpDuGH8raiFCGQpmn0gG+M1+hAfvyM66t3FAsDmBl2U0
sAZscNXOIa1B0VOJEvQP4ljTZyJNydmP2YSuX2/80XRvK1Eh8V8xTp6YjCjYDD5I
0CV+BpQesXpgFIRhyRSaXuNlPa8BmvqtABd9vX7XOvWkcsL8zZMfHU3bCpqpGdyp
PWWvVo6Tkx1gpd8S8RiX6Mi7TFBbelotzR7Vc9Kt6F7vzRBDdz/HPIzAakyMKujS
+KJWViHth5FpNQgmpwFy1VbEm0TV8wtNovOa2DYZ/x2q7iRdiGi6dDFG4ROVcf5N
2nw8GE4xfAhRrG41Zpze8BEu+l5/pYdVOxDq8J5nMSKFeIwMEsWhp0W7r+V5jy3f
ehEw3N9kQcsScBA25vyeAoNJE5kkzF8LxoIcExNMFHdBny6SgEbvq1VU7mfb+G9A
B3MshSlgHcdgV4fDwDNmzvcZqzpjrRMB9B8ssMKvP64cAbnngjR9eY5l4TnBttBB
Ide0uSX7bxopxiX1UGuNdkHUMrHD7GsqkP8I86ggvLDmsmd0Nsc1qRB8h+NbZozi
jmpl3CyW2HvJd1lXU2044EvP3MV81gb4yDIjhLKYsfpfYYdEB90SJG5qMHUcjHm6
6Bb7hf/Bi4qxeUFcNlA7wPgQwiA4paao+Pzymfs4bhFix7GwGQfRlMsWCS4E7RrM
OQCnHmDJI2SWTlznigJi9KHe8WzFPDzwTs/Hiv3eCvGZBw/VkIQldEwCZKW+Fdt6
HNDs3Ey5mBqBL+QwTxNEPOFRT6cQmWBQUfPH25gPefYb7od7ejGtOWKGq35gQyxJ
puq+BWCwPx/kYtA+dw4MgLu9M1woQAjL+gQNgOn0bnJUW9kiyDQ0vj0G5ZEqVVui
IO1RhPpx6yjAxr3HMyRbuS+F46N7/hbFQpzWAQ8nzRqbn2NDMN0o7TqVo0EbdrRA
8/HyqoiR66Z0ZhyxRerVNEKe7xJ/HgIFFhAmb5HZwP72Bk8ll0yovXXyyXZgFUEk
efKtPltFI3Xu7xsF/z3L05IAtyMPXGZNeZq6+G1hRJQ+gCt9fKcpf9fNUsDa3HwC
9cQQxZBl104ftzMk4tnbKrv0PrxfuhsLShWu+zIR+J7LjhRtBlRsxqeyX848vllJ
9Xhbx0E/zdx9EsKi02At3LGOapvMtXvFaNxz9pAOdaEM2DXVH9vBifYLhz2JTPtu
wGOFvfPBv1wYKEtWETs1f/JPD2ySrMSgfjN+KALlmkIodv3EHQmBSqyDuYNm5CMq
woZa8pjlwE3K7RxNZB6EyjoQ4gRSES2KLfBdJ/AmInMsjckB5wbC6DVdDDcEOozF
ADJqtYF7y3e6wGP9B1fkRMXBr/1gT6dB+oDJj7n0guXc0+wy5v5wPlRawxlHg4eb
Q51MH1WrWJhZ1boIxYN8HuWPotFR7k5HbyJRe5kBzC6BNRXDjJgccTjbm9UpMeNR
qsjJNlpkc74u94VikrjaBNgOUST58ks/RRU0kSlieUZyz5qWqUH5VIxakySkeD5K
Pqlz67lF7aUXlyITmRLoKt7xNIvzPUZN4FRZGDVwBw425KN3NXJ+5zk+O2fvbr+P
7ZUfoPKtudMsivCROAFHAIMB+rSPBLQ1GF6y9ZGA0K7NM5DXhArrJNSPbsdJjCFE
77lrQGMxFGsP0Pxis2JT1LhZVsr5eMIuFWLcmvoZw9N8WyUK693iI8p0UmVkAejA
xz7oPcRP2oiWQMTUoJmt5QjkeK/SAuMh93qkIlgALUJhKZ2/ly8Mrprx85bxh1Yz
gPLuDBJsmdGf7TTlQbil3Yl2PQniaFOEkHYJta2Rz5ranKJPaexaStP58BKe06XK
eRKZ9yqAMN/LdEyVsOnrf4Grzjy1UKdA09/hhaROTZ4Fa+pSQW6fwOaaQlYENySg
D+iUeREfWT+MCdGGjsySJ/+mh8oPeWuQKwJTQtgP6gfENkO5lXP5LKd7OgkqFyYz
ZUeI8a2dFndwsJGMrXi9NZeO4xcBxDfi/u6MIakfCT7Mx1u23UR/cIx6eHZJYZxM
NfacfgvdO3/SXiYbqwkB5oBK9mVoxDP8sjX1xIeOhwgAqA1K1ZxSS5ODcwdXwogV
Svx0MKRyDYJwVy3u0opY3thk7tsaJkxnzM69A4c9z8v+f9txf10kwj8yRMxiB5Q6
FD0GrnClk0AfwpV9Oa/QDSo+fengy0lNAqo0E32Kq2CUK3clocNOS+2yptvWTckt
PLWgMoyNtUYVAQiZrGRebdkcY31UrvDrD8k4NOLxFaYhRdmah3He0BL2gf6mJYrA
n9AQQXDmkbOEd0pETqyiYMguf4wkqNRFtuO7XReOEN3PiF0oP0pvfSt9YwDP955R
fwcDVlAAVM6qMfTc+T04QKW2Y3842YzEDRJCQDZl4WVuu5gpV2yc2wo2thAOdYHe
diBT7LAGBQOPTxEdhaVA1vhYwoscXiH3I2oemvg3xzHJMmsOqblhByC/lBqnsvjo
0BrZSBnEzRADiSl+C11fgz/p0QLN1XoB2WgEJJrJgUbpBoUmX+bdSD7j7Zgzn4AA
g5TrdgUNyg5HMN5E3rIGgyFk5iep/jJWZISb8KintEtsGc5DTS+MF7EDOFe5J/Sd
stDZsieogkK2xCwe/L2di67RuWuKcimMb4Riq7TWsoC83hgQdjC9fCfBf/CORdoB
yqWWhFlhdGA9vr5xNU5uRfskGYaRvsbfmibot5BPz5Hcags6RfVzA9bM98dsPw1M
yRkbsIl9t/wSC+QeB6nH+3iRi6110aofktQrD4wUkpI+L13yrN6q2Dq7FJ4dKd0O
ay05Mnf9BMI5MMu3SESCIP0bxgqrLsVPJnyxFPF332Yl77CQ7H9am7fL29AFmPim
HTLTZT7BADu6zhVysoWvu2LD4NYVqRl6mn61mAu4bX5VW9V6FnpR36oxCbfK+ncP
mYjb15HiZrIMQUk6To+aNYpFMzzPACLGsvwOqpOt1u/ygAQKY1opNBvpLoFe1hSy
H++oAXd1WkvXJ5cfSyxShBrKoa/Ug8iQknVMXXVBoM2PTDiK3XWjphHIbAKZwXhj
m8oKNFWMkpcN5Kc/mnHfBt0F9PXXrFyd6rNvWYDi8Fvp5uvC2sGiOciVLqJ4PRiO
KBDUdLWDtKMYxVtxIdKeLQq3n+AeimFrDSAei0ZH6fl3emDYHC78C1MWMlSwxY/l
DNBz3GvkCeC7ehtnjoINzNv+i/SOBSz7Dp7NwsqCRrEc1FcbGaO5/NJYNXMpTtkJ
BtP8k72Y81x/Zu/t8qD5VD+T0kw8A9wiolIohWrRqahve5CULo0iPQ+H9YN3waMR
P0+vgd80sjME/TrzK4RNN/R9g0Rnpc+tgobI2AwBFRl1td0g4JNXMhW91NnKp+/b
DpsUWwAqvJEsv0uKfUKmYJ4YwrIpWuZvzm1lJhMXduB+nQoIDHumoj5EcJuQozh9
CAolE0W0IiULcN5WABPDIRTB3KAEqjWrl9jCeRr0LwyD3AyaorlTWzOA9d0+T0VK
Hmvbgz3DrggKzfQOVp+e+3L46WaG/b2Sbs2pM2/zzWHN54W0Hin2XikNheyuqq/N
FHvQ/nJDTMXfnvfO2kIjxNstGH8r7l2mJEFM+hNNF9myQQ4Hu8039S8ZI0INR5Wm
A8r7CP40weoDLfYmKvwUhnt4nLu1WPfAR/TrpO8Gs/5rvUX7iqdERbCcO1oU+Zr5
64PDGIvcL7HgpIJvl0++djY3CZtKRmXsHLJpii7zurWHYg0zci5QNaM3annZm3ly
fywEz3dobLf395bncCpbgtjt+TT0WSGLKcM3TzGueXolBc2BMpV2Gxv6tUk/LNa1
JbrqlqT0krNCcEhHn0XsFO3vZFTeKiOTEMI3qP5c6fUgBb384uMFhNFmS1OzJby4
rJDvjQoYEF7/YrcS3mZ9JVFTianppL2kTtLD+53y8X6AVVoDT9kzZQk01zCKzHz9
trLv1vnaudAfdeDgjEPhv9kQl/uxjx/Tyi3uGoh1fajNGiwJkC8lwL/3fF9GBpUB
MP25mx8tAR7c7LlAwTkGoXsUhkeyc0+LIqv/vIrmwZcqvQCRGvS2TN3d4yzaF7Cx
/JyN8uYqWFygJ5rxdrjvcCGDzhC8Q0xr1St92WCxgl8lNva+4EeJ0S8WLnMWAXMb
J8s8g9Kjw9cnkIk6ModTWkQHDqPT2QDvaoVFDJwP1+E2ZqmNc8fecrCPrybPv8M2
PtPFt9oV5jRzZ8L5UAy56LfosWi/tlG4WfZHzeB/EJu8tUBimO7OtNtVxC0vP0mZ
KCPGikfFSSmJ0oBlOKPX/MsryzuSAFavNWVNPaNvF7L/ZOqGZwE4IiskVOlicfje
dHW9AT/4cOR5UnADTlMPYnfDj/4fs0+J4dtC2Sz3s0At/GzLjIqrWe8ql67uBnTR
32fqmhjVgQHpZX/wOCiBHSqf72BzhCxQaMONj6Fm1Hcygo3ynOv5md+w7ag+7Q9k
2Y1Wf8gyl7lofCSp5Ij5FQm+mZTYsVQRHdYBTK1YQo1bH7TUnD6Ad8dlifJzmWrT
mQ5KJpnqW0oPSh098QyXXt8AI2+m8DeXN5TCO7tYt/ZdbsGj0cjSKt/RGBwd7jDu
vPKHOQ4g5SDxvNpHRSsKeFNFjKuVfy06qOUt+1zUQ/D5+Nn5C3mifTN2MqJDMyr4
w+/MmqhcAT7dMMmp1ceJ6CM7DlSIw07Y13S6w7eFChB6N7d/Yyjlfm8f/b9k+298
UvJ5rFxUelxr/WiOWmnacrE8M+FdfBaqiwevN4xTho1Taai2RVJ4hM5cZNYD8sGf
kSJMN9avkOIuZKdzrEnNXbPIpMn9iyPXX2IypaJys7G1yx1O3Bet7Dl2PN7HiIDI
DPgOSzk6wUT34bdI3rGJ3m36yeZJqglp7x30L08u4rtDZLmwNCDCB7kgazPBNAX4
OY+ughcKWAgUqQEzuI45SMbQXK5gMOCZUZVpUWJ5wiOocWB3I8FeVA/bZ1AvdG82
uk3FwZqEAXa6/UXya5W2qBwWD9QMm1ftaUDqQ0JYWDf7z1B5cvlVnUHJdXwBvlBz
NzrW7OLK4jlth1t+R6ha+RMY4+HYUSZKJ/HvvPmIMCsSjck57jc7FpLEYc1UwKlC
rBAaAs1J/JjlcDRAUcDGDrzyNQm89xv3HzkSYZRMi8rS5o7L6giIHuN2RcHREmNW
wC2LRAidVSlvC6JRi0lWJAprzGYIJLR51dk6SN2VuAFxHXBktSEIpbpBMT//bqdU
HCmS5cs4Cd3mUTVwGein2uNd3l3aDEBA+wPis/nWUYwSPKqizHzRj/c2qCBBu7fr
ciyT9koRsN3ZS1G6NvKq3jQ20bL1nf+PzGd6IGjxN1lO1gwP3nKQqTIcbz4ZO05+
9EaBc0r8Z+/ZES2hEx9I6JFddUzsu+L/xAf48MEcGnH9RTWkDd9XHe1HgJk2E7Em
AVBPp9Q0mWvgk+Cp/XfMTSBHouaamXpQlkqaaoZFxk3DZbZfV3lBJoYKbXXMxSWK
50fba1lzamnqKC+ijhFdzaXiwrKolA9THWuc0n+mQLxEIASQQPq+I83+1V7BwAfc
tIMJV0E70GiZ9ogodTBdNP1Gpf1fPaG55LVia7kxgmJdB0C2vjwzYpnAs6u2uhGu
UTl7xpZJFzzUHs3WMeKaU8yMl9yxcm3fYLKr4nxgBh1LKwsDbnzuHpH57viPWbWi
JB9rxyKVcghq/fJomi8/eqVSBuaI2P5CGxY6v2x2mMzZh+MBtCbL+/KecuK4h+uJ
htQt/6mtga9ufvhJ9qoFHq0bDUS/kZZMSfoES6ODdgy6WtSmuqptzIAzliJfrfhV
C1XfKTrhhl6F1ECIpLKdY6kRlASE+uwOCXKgn7s7VrfD2SWuz9hpsfJv6xMDUvGw
rZ2vGWNNJtsSJV2+tkDTvRyvMIwqg4yT+/8nXbQF5DW81Jl8HpdpWoM9UUWnLzXj
MRdf3MJmPjDn2djzLmSIcC/KP5ZE8CRRwBv7lWOfcfAOLwgP2KOO5kT9zYvcDefa
sWYWiMQdxw7Pbx5A2V7RzAD/YkmCuh5nv5PeQ4iYfGi45BGO8GtLVXW7bl0xu0Lf
4lwvwHtIrCYPNiHifUFVR8GUJ4HEdSqNffc+q8OKhW4fmi3XVOiIL8mmn8Sxw2d2
vIbDXJ6fAtPrNVI4q+N7BneD1ubMSA5QPIzdyDiCghLWt3NxqE8KYMAaE6JpYK2v
LqM26+LcKdS+4Fz+Bl4aMl1sxAc52CF+vi7Kw8rbWntpAZcEYeQX7uBPxg3DO8uq
HUmNoMie397955+e0cZaqD6BT/CJc7CaOmeUg3LmKqIA9/7RE2hxHfy5NFU4qudY
9tW2tV1aICrbTnNsAKbgRpZWqfKUs6yK6J91KlQHOOOxDoljWQH0o85Ys7fPykSP
CKHIbEz5Ru++luauhABe0C33l9WtTG3fx1Kbs1d3laXnz2R3I2afrrT0x51+4V9z
ZY5+UsHEc616++5Ouo+nRQbA3JfsewfxceScli6zgfJtU8Xy6iAapEFCROHpjR4Q
N1cfvi3538BRFLMlB2RZESc0LyoR2O67YXwnZpwToDQ0khMxglEmSaJo2WT/Qohw
AQLqtNoVxwaasUNfJ75o+JLFObv62aGT6GRCl8horlwz+4eeu/VlpeeJ6DrGArkZ
Ygk9Lq1kdTtL9Vi6av/zJl9MVVYFYAgH6ip28e2uBMtviJqTe5bU4me0SAc/pDVn
xc+7Eh2FLgYpTm+/uefMKOflTfPhnlQl4eN4kChmsd8eScKEIioM2XiY7ULNTA6b
y+2+Z8a3ICQgiZi8uhhxEC67r5NvD0LVwM8V+EyrCckcG8mRI9+GiSn3zflm/lfe
1Ei9joiguRdZ2bt5rzmObYggArY+R92k18nlO5hW3dC78tZnImIb6/Cn55mlCkjJ
Ytq7sttUZhIpQcY95dXjW3IyZW9Oh+ItAtn8/g5Lj8syOuaL3VEr2Ki0Egqe0Zuz
yszN9BtSqR0bRDYuVxmeheSktzZKqUCgQ5zr1RKDxnvk/Yuu572GIatEjkqrbFGt
s2lmSyTShjmI/vkKvkQxkca6jG+vMnnk5tW6QSxbV1akLVhV30e3TI97s7DpXqTA
CEmdya1f6lzfmoOdGIbKMJ+1kn+m8IZFgpg9Oop8yIX4aM2Vo4W37V5VL4N/ZebF
G3FqlxTGvtyRkL3y/GBKnVYjl1uXP0qSpU9brqaopOx0tDGN4eQAwQoO+zQLV7H+
TCwu8tt7Q9cc12QaVW619TQR5UQaixAE7ZqP19xISIjJlvCIG1HdKMEEc0+oKyhp
RpfNph5FrF0TbHQ+vuxNTxr/YVK3bbGyFLl8t/OTLL+2c+YY4HPCOy0llPbuvvQP
MC99U8dxW3WdfIipxX0ZPa9365m6D6rMqLVAOBfLGZMz6Ivu2OfLQuuQDaDQBPSc
LlSUDa8rtpxtYE0eivdqtMaQKZKyZ2XXTGBMgkA9Wm1nYb5egPhVN2ZVj0ipFSrI
gfgf5hntA2bExyYORUs2X421jdt2j4nzASwK5U7zJVmySWHDDZQqpRdSJJNwoyO+
LiVM66l4KRc3rj4mtGmtfiubDx0VuBCc16sPybgRMXLOQf4nfaoFTONJrIiQXFg9
5WvbveX4T/tUGYOhjgh1BV2vNfNlXqoxlKGk8auaaMp3ccEVFu6hfaafx1MDitDj
BRMv+079tppSdGKSufgWKHW4zTW+fJP9Ktrc4GEbCoFQnXKQnD1VqMkn8hqpgMJW
iuT0lzQrAChcxGs07pow1WGwsuADb95S3ZZxKY1u2QQIiF829Noflx/cIfRoFj8r
gMN2LDtvnf+O6/bLk2FQWBtOkwFth70foMXCg6Gpi7YF6LBt+adL6zySApQzooxQ
jty53AxhO9j+L47Tg2U859QBAYvCUXCqYJHttO26kA5OFjfr7yaz8OzwaS0D5iox
wWovwk4imyV18ZFOVs7i79Vefbb5b710HC4/f3A2rnDNpP/l6fjdro6R4bPBUWzD
C6tSudHA41u/CwP2g4EUy334JvAXQyrYEK+Ib5Oa2aiWmm6ll01y7Eryvb1C8NzX
W3gNYjqW5d0XdodMbOTEk4XYLM0Jvbz8khZYkfqKygZYalY/SkGYZ191INquwPMx
ar8z/xNDJVLvFZgEb7zuRw3Ysfh7j6ODvdUzq/T67dX/h3YPD4gcG/Y1fshd7YQ2
/gse+Mn+jGCwwjJt1ifp/AlTGtLy8MWxhceoxf+gTkUK4oz2AW2AdwgHNAqIyI0y
ihxk+R7bRkEAtOnXcUBWNb7BEuiL1qBnSvCPM8TjI+rNvCizrH8JIATGE9QYdFiY
56Sw4cupGuqzAD/2FdYzIPW3Jnwms969At3y/aWao9HfALvSlWvqldf6iBDACn/R
3N0X/6D+u12I5GQG7WFW5EukS57qvAtTB0eYiIczSQw=
`pragma protect end_protected
