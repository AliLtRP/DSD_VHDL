// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ndq/lAM+pYdG2UXLYjZMlD6sBNDtlsP7ghNF1Qq2YhEwMXkCJouRq0cbFEMB3aNL
UVSe1zp1J/Nk/qInzE9vgElMDg8T46QMHMeeEN5OGC4iNpit/hprbs/wa7wro3iX
XN8dNevc6Qzh0M0XhLElPam8W5jHIiZ+2m+nKLgXKRc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12688)
nKjp5UiYWLKaJHk7L+aE3IOLgqpP4prFnExpRkA5ARO17rRbTzXHvDFy7SPSl/3B
kUMNmfFvTHadjAPWQ9BG9CTIHW7VVvIJR7CASIOIe6A15Hy7edo99zm3j4qGytYM
Z8rL83m8m9QapXhvu70u/ACxAdcApppNP+g827/HnEVsNNM12wNJ31WL/ahJJLfi
T0xR9S+Z/EFKjLx117gJzk8lKY1mcCiSlCNeo6maubmPP8lJNEiGpePQ+PiN1wGD
c+PFvdc8S/WKlcFVYYT1iIZ5gSRkzNtwjXIBE6w00wEHF53A4O/i87XJEp+wm31x
/O7zSkTovB3TyniXxOiIHX+cO6YAvJfBw6fAIypEbND/QmtJhWmhrMTaZyK6MGY6
XipMCun/cSP7DafEmRZri7wJIoBLX+u+vVEBmNWuHuZgj4XDybiaahtUvOS/tStc
yoprCOkH8LwDbxqIswsRVRY9XcgFivDWtEtf8ybPFI5H2ASxyUXz+xH8pTh8YnIa
vziK7dQTEe67WRL/Od9LZYwzw9aeIIcPiuHeQpFy96aQBBKDk+KBpt6E3setCV1U
Av2/AtAtvIiS/v5bxd5jUD+PK27qGiuA1+v0rg4seMlQkfw7Gia1mCYpOm9fKS19
+/PI8gMv0QzFts5y8xWpR7Wp4clEfpooL0sSQZNCam8V4JyXtkv0TK1tRaHmi86k
ikuOfv/HizNeuHF2eJ0nm7Ck8tD5njnrclvixWRKRJsxsBKPEng8W/vJCAlGCZSH
IS9iep5jb7EYXBqyhVo0SEIhX3Y9TBhLe34O7Qwl3u/PEfX7q+g5Q4NqOwm86SUV
QYHRy2O5mkCS5dv+rfXFgf1KGmoC8ikoQQx+f5V5hyqmAbezExRgtxILIz3OJzcC
F8AELGtQ2StPK6+1/IaUmFXrEzJMW7f4FeX+biKqpFxe5OPemuu7ljQvT2DbvmEH
JgqhGpp57SJP9mxlrOCtTbG8ppKGJCfHMPw3e+hwwm81NL/sTFTumfEVH2H4spJ9
7mjwWhdHny+hMwNqNXz3M+ESJWcex3gkWkOvQyhEeGCYPAYwUFy7RibLPHdtgtN7
5HCUCE55Z/qBUHMJFLe39SWJTQPBm08UtTnpZTkF0RmiHsE3DTr99AfMNH5bpbUT
EBQfKcJVTGCV6qe26klHZU4NCC9jl6Ybj/tKUT8TOPh85LcpVwsuYl0JBHnB/f0r
PtiilXxEXLc2FYQu0PoOR75+oPeToKY63D/rXWt+TtLpITs3Gl0uizsbDfJBCEUx
PAKGePasGyk+m2vE90I4IiqtVEhyIMw6KaRAEuiQuhDDyaIdzi8TKYlZlevA3m0e
GQmOHB73/sOCTAnMZLBnf5hbBI/tDu4YAoGufpIcJ96ceUsVE4XDm3lRttzL/g/5
ErBXr9+VXJcekCTKREWHnJOH3Fkbmq3DrHHCxX3CUf0pBgXjd95JM2vaX50cpEUN
zG7Fem/WrkkVdF1LB7BdV12+XrV6pHjwYVsGs2+Xsx9Odw02bw+8e5XUw5AMq84b
hUw9M88bCsr4AuwRe+sLL60B1BspC8PHdwU63NMoIj8TmBcXWbepqYYA8s1cJCOi
UaAdq/40FS4QIyd6c6YRTvEnT3GzEyGDTibTVBMTrf9qzPistpdfnz0gzJo3jgqq
8falZYb/QjPuUbHVYZjxjSXLwNr/cNQChnhLpa1CwLMOcu2WNmw5S6fApr7tW/xs
RjbZtMBrmYojvk4C5f+nQeXBORjvgbxC8xg78H8ph3UN7ihz4SlKgI45pF5eyaPt
pQuzJD/q9B6kQzxy+vcBdxRlniyVUlQHlhYJOjGNC6VOpDSfo4Q5bqqswnXJPzUE
xYBfHwEKeg96BgETXrkhACNSL4f14DoZfDqu4OdPw0VZRVgC+AKv39Ht8ROIeM1F
4elLWqUlpvZgABgUEEP7gTAQ/9OCg+J2JxSWXUFlIofjreqPw2UUKxn6ozBl28vH
np4LDyspHVYKhRJXOj+/X4HQcUP+7hR72jLQyDlY8qhbC+Kc5xFyllSd/n2pGKQP
iopdAJAdYO+1S08berfNVhExZn3AOnAo+8ho7LzrW7Cr0jkPiEiSyY3j3hiFVRQa
jiHyzIRKeLVVdzgT8Y7At5SMwAJcvC7uAucZqzx8GA20EP6i+aSAAujj/Q0SWwBI
9Dzieog4xacosQKPgg2hL2azZ48qmcUImg6SN+WWEhX/bBrtsnQ0w4WVupLXhRgh
xdP9Tpb0Frn2BBwO1XS5yg0TE7Y9RaJlYREZB3F6o4bBzq8nRMesUs2yuct/wsc5
B3ywaDaVNo5WolVSs7eG14PyzwUsit5LRDO7roaw0kWclTQkC9NE2iuQQVJSnZ5h
X5hJZI1o2W1TB1IqPGNJkZA9plEupOnkunu+JgUKU8gxTp+vxsBf5GbvUgVXmZzS
Cz6e4KXMRS0HU9lwINcR8shR53yypnSMqaljZrG8DESIwm9FaWTgISlTkuMuBx4v
XPGIDFHWN2IaPQsn8PCec4y4/4oes9Y8PVNsjKiBZUhffnvnQdXbniTx+SZ3poUL
rORL9p1bRlipD2Ub3Fe25m/Lsv2WYMCzPYZxOIwE8oxl9lpVH1SwdDBrJk202MJW
HBOmHwwzgwgRpGAEWa2MsPNc89HCEW3cPQwewFcHLUncG8sLSE25UW9P290iKEjF
d0TufNGYmmsrkBtekd1GVMzz077xIjFA/5BEpgMP4gT12Xk9xmLcedw1/bKb86q6
TFtSBASzxXADoJ8t/nIFNRKfbqLUOUtVdXdqu8bK+IA2CdM/4lwhThMMz5kvqETP
G91TYXBTw0lVMjRQa6Jo0MqpNJzZ4HIMLLfpe3ZbfyLg2ZZh9vEQzYE3OPj1INRO
bjXmhcRhjBoH3x6SnFrhoEZlzYqb7wjGVMJstgGRxrGplmGNCLgN+VtxVGJ8VBDS
TrzIl31okVvbpnysYEVjMOa14/B9SxeyQeLdGcA5ByQ1jsyz3aVcvtjhL7mJH24l
4sx+sWEBPkapHq7fdJj6lStLDvYkL6xzp3PrC9JUJHANZcTrICAewL4dLf9MtgKr
5zbU60SC690szgCGzFtg+cA0c4F5tpOe6dd4zVslSmikZSntSF4+ghRAlNwcPNhs
sNpcwgc64OjDBIApHhp0fdIzF8+FQdQh7fX8V/jmgQuV1GVmEHd2Zih+R3qcmBQA
carwP6Zropw587G6ZdZW2QPZEC7aVQGMLTc3Wik6Yqcn4MekHQDdR4hg/YFRlb2i
YMNNHDze6+ic7Q7U7ZynH/ozBeMQLuPrlWtCHL226i3VvaHhyUtckLfK+BgoQdlH
XgvTAZaXIckRS8IDpPOyNks0MRfnDGWEJ7zYDcqazsKZjxbDZaEXJyBNxtrmCniY
u68KYAF86b1HlKQpnKcTK+CmwbISJVLaknAOkn+L3wR9crmIpY9SDbz4Elnyj1DN
qavHf2HX0FiB2x8xseBR2qaMWUjMDX+pMvMr6ykiFvePsLq3lrfzzmm8b614Nk83
UTJiEkGkRNjZChp75277iC4Sh6ctLA+vfQBeZXG5uhgjhZ54ep/GFJeSJ08444NA
JwsoEuOgwJSiKPkykviNZ2AJIUrCoMPEKYkX9WowqLJ/knqEMM3cukz2xV4hmhUS
DmGvGbyptpBkispjwGWX99zxqmgf1/B2HVOJJWelUBp+J1Xm1Stx0lYLgmeOYMl+
nivkYqzQ4x5b3jpx0Rfw0rwEDLLkWWeRReHPOPhxRMk/bPyO8f4iHV/bzwXHNAc6
+VfFf1VVqlyw3k/Fk1Jv3nZQYxjZf0dOaRDBE/WR7LRTi7GIDUeabq1O4+68/svx
9xtgWPV43V2/44BpaU6XS4DAk/6qaDdrrFHGeA0ZDVVdYRWw9HrzNTIb4wBH0pmr
kdi64h49sGJQW3rL0v0lVp1OpQxZtymbQr68yOWOJBV8OPhFyff4cvBYrl6sO/YV
UCwdozlTK/dVfctWGdGp/WnihpWFNYGbi2eBlH3xMP8sfVdmL4UcooqBDrEQeymG
Zu1LSKNIPH4EYHNx+Sm04nv4+eca6QVMQvSaL+vn2RFYDkiSc5nomsTzf299tL8y
f2IPOFgr0d4neOiEb0qN4ocyGzCmCu62omim9BOLZB1f3+mwCxgc2bnv1DXGdEv0
C7LOgRJTLor8neGtLenCiZaIwCOl2kJnzjEZRUVKC6mtVShkaHoZXN4O/GyPWsL0
80pwPqmCnqbY7YHo+9JmzR6kE1KuPstd0RCMpMBPYEGUqjxLMxF40fSmcw4p493k
J0mqNZIQclv6mXJP6XnABRkKTQrLpYH+osppYyF1AgnuUN60N0oUVHgH3wHoy46r
1t4RsFa6KkUghDQlfF0HayaNib4hbzh8a8rigfL1iC1F76oBpFkgd4N2tDwXoI9U
GADr4bjTEon0HWT5aV65FV1ubffzZywB9MjruRcjURPlEZr3m+fE9vGlddCVmM6m
V/f2lE8mU/a+8XTIOC5zUiVY2qAYGiRscTxV33NXfjhw3Dbzv8n+t+tEBYm+I/VF
exuhwqJMqWqx6KS3CfjoOX7MQyc5/q1jL109tdn8EmhzGi247he3aYsxDR6SBHq6
WwzBzx/5kI7uhsN9XhcfqEMw58S4wJVcOmoXLemwRZjddfZv+1jIN6dMhnHdpbG2
no6hcpYel7IYNPKiaH7ER6qrI17lfUQNVwNiFJkGQ2FZV2XkziJyiY0jCSPQB3Ol
yYF38f0KhfSZw62jSYo2G3sjLxJek5zM6B0mwTRCba1geWZ8uFo8tfID+IHbx5gB
10b7rKy/NioShTUSG3D/8DDnBBMSS3kuI9PwS9DTiSnkWz8iQQtOFC6+Y6Aml7nU
1MCdgLfxHQfSha3i7+q4Q+GmBmLxTwekuonT9C+EGkhed+V/1Jcs6Ry0+oTSNCjJ
xFeP5QBf3OfdDkypzeNg/91ZCYm1GM6cSVM0EwAM2A5xsS6cZEERk64nksgPPExq
SdaC0G83pZMU8v14gaFUvsFRPUKVHAHd1Oe3lrebnqr0ApPFR6zuF4lamG17BlL1
GfDZikY43wLNlx49/zghKP3hDd5N2bGqaNzfPdUu9LNq6S+LaAnYsczs0/GuB6zF
GqmULFhVOeVkHltrEEtaXgdTK56YOwkExq796brbntY+KRz0im0/651vBASUyaVG
+r14l0jvhY6xIupBXjHhVeXp3o2tFh7Y1GtASifXhO1k0awcGj4RHIfHptpCQseF
TA7YYpSiuacgqL3VRhGj8OBv3rZcJINTIZBOS4r1iZ75qqqhOfMXk10SNj/imPPy
WY7PV5aUIKYL6x6KOrApXoaT48wrUwTG3djZGMWv+s0ySi8eEJPH15EObkM2XqnA
9OWthPXVHt8Q8gNqJvQKAHZ3AgEtvFSdTMeqgCps9ZM1mJcOZpEhU9Ho2gmTFHaj
C8+ZXV6/hJAvOix0sEB5npH+6mW7EdJQauPwjHPrYibFSwldDxgfpaiC87BD8EDJ
k5CoA61WjpHIYoLjNEFiDjYzfDjAmC4lae3/ECq7ju10Pb4zomZYx2b8fMv2UBsS
/AjIIPalFlCeC1sNZ/HykblkBqT7v/LvClUg04AV/qLVjGhlt+SobFG1jPfHFnUQ
1xWx9Nf6ETlt2fI+JNZl698oDb6+rY2RMzoU30/Ym+m3dvI8gPAEB6ARP2WUW04u
5rUK5mxCDqPbsPqwdOl5ZdZglJ5RB4cbtzVXhcdJu6ZzNrNxqiO/5QUzBpU54mIl
0tGbE0ZQ71LLgh2wPkigVYrz4p1+aFtvPnnpnlitRIOwMSy8W8e5xMf+j8Q1/R/e
mhB2A4D1Yrz86fmelej/kH8Z/bJslG+kZL2p/UyKMYVoDSIBBRrw5Ir7/thvyEz6
caIyhPu3YLch+wZT4CnVpSIadasal4Qbqa81wpWbOdO8B1lTev3d6rg+RJdXQ91z
s2jnoULt3N6EoGiYg74ILqlFE3ToOXKfRQgGsjP3Jrl/Z8hPOzjzsFLmabnRYuXt
Aq6jAj/5RI2xau8N9U3A7a9JUshFOwid4E10jlrjN8E604w089yLrzlkGyjiUCYj
VydmnL1wDPmN5xHp9wOUD8XmngdL5iTyhcDJ+43jQHGslkZ51kxvC0pKCh7XAnpX
fNKu8QricOwNPDXihYrw41cPjW5vc1v77UUYA+hlOW3TLd2v0JnvG8yZsGV5kBOi
BA7NWGoSl3QesI+jKV92zEMiYAvu+0ZtweRD0jOE4i9Q0mCL6bLze8+gpjxjSId4
ott48i+eToHVG0bp3K5UHvTfVnJYd0SGLx4u2qUrgqVKiJHXvG3OGwYfHO3wf62s
AuaO64etqL2ZFmchzl/arh7Lx0Uv6NMJeEVKBumJjBPpYFlYmHwfRFLwDuao963d
XTheIT8Lo/17CJslrdJkaz17Zg4M8TREMKhcLBatUuXWehObsRQNesJck4IonrA0
aUJ5+khCm39FhJw6dfWYWHifBAfxKshhjbUu5LClY07+hX9xQqUoQ1oSKUPadG1q
iDJ+KRtrAxhN2EsnnXs1t56Utsn3Q54mrgYvLh+4PN0NJiI1FFpC94whEqneeS+U
Oq+4Xtg/ee9Fsr07GVtj8xZFz+VyLDRfQoGyjqfyrK89WSAM1ElKzMn+klWjPKcU
H6FBmnZZcWhATj62QbHoVzmfsl4EMgac1+5mpqBGq1xY2oqMLzsRvyHQiIC6u3vl
Y4GddHu6aSNznOLa6Z9D/QoagRb4XVO0b7f/p+Bi0PGg8PSvWvtpUhVEEq7JHR15
PLztsCz/FF1IgHUxZQi3rgr6vB8/n1yRqto+TsF4L54WDzYIVhyJr+4PhPhKB+MI
n3lXnPHrEVlQopQR1lFBTYiGWgZPOSH+CH5pOBJrKeCZBDSRc+YJq3i9VD88HgA6
BJABxd/tklSXffzFfzD4GD32IQulmpufdYcSZnuR+JZT8Mw/H4IyixEK9lYyzH+Q
OXWzsx+Unb21NhoGcdqFiqQ0jvCxklCPEr467x6Vn+LAbw7H/qcqxXvM2VU+mLpM
O4hRGIh55tM8T47uwks8LGG+QSUQCEkMLuOyavxEimyvd3nHR0t2pXcILIjBaEY9
V3tpUHpXJWKiyw5zx6JIlaEeo6UoOb8NVvpu1Bu23XN3aW9zt3XtzhQs7wxaIAyb
J/wRxmG3T4vunQcxGlD6LKuN2hBN5nYAOpzRix2I7Wa4TkJlIBHzEDZE+RFF0WZl
oawRiV1aR88lBXetXYNGNfYoIpX3sZEZwWpQAPG3o1xmygr/YzliDsE8kcTq8KAr
Zt+EFd4qUH1VXunKfrnKDtjw8QKXxcxU+qon8U4o5cYMG8Lzjl2hqEVc0dEyiVtG
Vt+KbzNEkynzhmGQ74gf8yNbl9b4+NR67TeLR++EsUvry2SgiFLbr7wwoDvoWBBI
5djWo5QCb4dyUb+0RIge6o/adpabM7cYNAyTRQs0IZqtgxYV0jDBl1jdWLS3yFNE
JPeerYx9eiE6aiLeL3zpCGZYqTeEX946nzE9hKrcHFPlZOCfLHTPrkPOk8oQJgLT
7i4xKF9vNfSj8xR9vrFCe1guWbCInuGav2rud28hxorczup4EAA+4LzfOX7g+SOg
xQzGQbooxnPv6kkZA8Vx3Gea/4aplGCbiF7KmpfcJqsQHdMbMvoIXMLL5EYlAnlf
tX/oHvzN4xkfmwB6ncXQZiYD+aCO/1oMGZmeG9xAFftgKcOMxiu3ayth9i8YKqlr
cvdjiJIxFIe9f3Bqi0nFlL6M62RVqWFl8zW6M9AAJSftac/V6V+8mHt96L4SFWq6
e7yCeOVpiJRC1Dab8RDmjXPrSbntTBG6v1Zpe1QjqvPC3A6rqODe+JKyxzz4m1F7
r80uIwpL+LGjZU4OSvNhtukZ+bTKT/jiH8EhGK/hoNUbc/A0/cBwqBNHk33HxpOt
FAIuPF4yt0vCqvPPL8I/FTYNhT/16vs9sTX0SuEGL3HwqfMw+nFnaSRdZuiYBqOV
vJitQPl+7CKQnrieUWkJQFY5uzw0aui9renqQRfbSxpIPQvLqWXpqeBtuYuMo3Gk
spJwAhSx3QoQ4dRDqwLXzF9bJgKcnhJkaAXx5+7OLrXQz/twZxme/B+7TmIFtaZJ
Z29RPBStJnNY+PFEbT1v3m/OmUGVKBdW1qCoj4LkG2Ysg8aRrMq2vBdonkoejoMv
vCGfIzsF2XCTpuPZA88TJekc3XbLUh/aO/TqI0RQS5z2/rOIzDju4cG0TPqijp/R
9VHzhMq45ek/2zjcTCmjL+E9LdFfzoHVq7zmSUtHKQbVX4gb0cAQBz5puasIWAhR
fZmSYNkXKSiVqVcflXejxBcC0pMq3cxV2xTOaxoDgWCqUgS2/SSHloWv7KfRrAB2
SXGpxO/kFHFroodG8SRizZdaAG5gdaZx+YYrybiVk4WWYz/wnhIvaJCokA99qESB
Ak8WQDrFnTe3Qaia6aFLhEFKOjzRjBETa+eLmtft0NrcN/88qEA/61CTXgxwbEHg
BOHPEJaMoWB5gt9MEL4FlaMPCzY5/8+VSlWc7nosbZ02U/3gr80Kllzw10UMZO5H
Noooj9TfnD/8y83d0XLtw0Phugc59GxlhuVJGm6KJhs1CsSXmbkGJrhR5VaU3MX5
z5ivxBX1j1OWt9ltmcN8QQN+zYpblrDsD193kc9tgS1dYlWasnJ7yc8XrUIyhDcu
ye8Z/0UydRAtDDTRJ104W6P0GctnORIWzy0kyYY9srXtvzbOM09xNhOFbdHN6YC3
xRkbHsW2nKteB77fgAfJFIACjLuTmeYSOJTzeDWU+IbMBGzklDQxL5RSPW9ivjTz
l1WEJRaDipaWJ8A7t3NPjDC2w0KZGZtTq/BLPYBYTfU0ThFVGjenvSmnBlQ9XFeg
p3QEFi2x29J7W/Elf6mC01CP0f1p9KTHaN0TcAiyR8YvYAbbyqJYQ029aPYJdIP2
pKQ85Ls/oEApFwaWiL0nZLiQffvp286tH+puvAXIW/UIAXAQNkpxdpT3h/rKEybw
23ypEX7gNPan4A/bIoMfihTWcuaTgmQGSZnRbRmD8B80rxDGQJT1lErHX9pH1OkH
4ZRUHwEIwScHpNWnG8+ox7xZesFB3V52JCn73Q1o0LCpyrHoglC8pQxSnh3fpNQA
QIg+A5WVZSMT50Uxa919jDbCWjHcRnVNakh5VLGZCLdIeglV44V8YpEFdnLTPdxL
+d7In/b1SecaXBtIfk3vILgUUjWHB4XrE/hFpOlioJjA2qUVF1LMLaYbVg2RSjwy
jUtlG4Ox4n5hF+xRIn3KcaykZjOhucULqJhqhIJQBurK+tNKMZtaNIllbLyn4uyb
YO4ugXi6ocuZzb5HRwtoMma/yf08z3XnXk2pqwtSn2BPqwVvXxo0PdKLP0U8XI/C
Y1swRvliwnlDToCXY312s6QqrbQC4xm8wYalNP6ZYxkTJrG4ZbbLk/gd70jzp8Mk
aztoZEog+TyA1j0eT3Iyu/O+/w0OWInoAzeKqynx7Xm4G9RE2X8hillRWi6a1Htf
HyGaryoixcOg6TuIjQuWxjn+inrrR1yiyGf3NE5L6HWPAhgl9LvD5dYmQMouTX2y
P8bPYkDITu8Jek/gUC0MM3amnaddYR40rbeFyfvfZ3LhJxx9vasfajmSYQIsDkQn
N47EIpRN48ZVv4t7w69c+h4MxJw5ZoFM5qpyedX6wEXMtdSELSZNT1XzHjzXsJ1x
9AeXQAv0XizCaEC7OIg9SSeER5IXYnvSxa9BxA2/nHkXRWNzr/01t4qE5gfpiIxj
OhQFyr1THB2injc1/0KD5eFFb4T5O7L8x5Lwtzou6CeywPVcmMcJ4jXD36TK3CnB
TgMJHvY+xzOM9Z3YDAfhvjBgL/y3sCz3SPsZqXXHnaZ+uwjHkMx6vWSF4N+TTK8+
Lw5HiXRKJULX/LSuf0K8bAu5rGJHLxHu0U9bhu9IDaPqsCwqnTQBBQY/28VtUN3f
edyeh9WsCsfa4FVjgrnOVjJaQH4O61u2CH7/Dd/JUWVe5PIE+sR8temBsCDmsujb
mEEQcarPAFiCyjyUVg9r2f7037NyaCnWjqtIES09Y+GgNJmMVtXkSjUh+DMC5hUW
8tGx5GKP7mNv3Dw8M5AIsk50HrZn6hxQDs6toZkvA/ZTlEcz8g51doDHO6C9FOaY
Vpi+tZsTjOSLWIpUBkHzpi1Mu7IKJ4toVpTRE9h1PRUBMwc3hr8a5DPVg7GrP3OD
cYCxoOz98IHWwtck2zAKtZLDRuOgq36petq6rpF2LT9ZKWRf8GdbueOBduuRURAJ
I2E01J7RR2vsMrFDSU0EgtGbF0eh8wHGPJrN+cB0rvzsxOvpD/ocxWhgEETAT+4G
aitnUljDhPHkyZ0z7BkrvfAD2vfnMrXjeqQgMxeSfPR2N0mNQnbLD8m4V3oAPfBQ
MBScyCq4RGPq7k2izQm/fXC5Wpw1emp8LYDImrZuSwG3gtaoBOIR5kgzGsvfrf71
U1qBRyjrqFLNb/kSmS0W90/nYBwORGedwXmrPtvTI9n06mdYp6Oyvkgg+JTffbXA
UIgrh0ttVpTwJdLegadJGbm4dpFh25Ohf4MLC0gixB7oY4gxVQx/Q+DSQspD/aCf
c14B73xyfskHWKHHCkAdAFWDFL4wH1uAoNFFghujTELxOZt2tXrM0G66gKOzSqIC
Xq6Mp/TGlq0AqcgOU9KfzCchQIZxgPD1XnZXZnGiHNRLgiu5rn31esTCZX59gudG
vFoIxyYeKPlVwLpaIC9AmXZH2MbjNKFKiRkmkmc5bawzNoSkYq8lsMbmlmHRdR0l
qu9xvjCOCsgvfCzQL4uMYyvRJ3U0U49PQFIqTjfhTFT/5R+/sWiNzP7C6/+YLZ+V
wFEdGNd30v3Q2u1bpPN0sY6rCG0PdXWfpG06EWB81tJuQhCkIfqUoahzNBk76I/L
78gYt5hSpD24KMb6wL1XX1zRARvXmIVcJhTubupBRMqZNVjn+/vx8b3yWefP4jzC
n0GTou+2jZc89J7GPTeXzVMEu+Gj18sMf/FmtNufyG8HNXhV7VV2ytTo3ZToOsoT
2uwhRrFceNKc41VYXmxYfTbBafV5XOhvGE0q+3yMfWxk1V2je9T2i9640kBtc3qa
0MQVXIQdh6QqaRGoFmPvPDuLH+k+Fjs6xJ/Y5ns01LL/eCYdNIpk0gpm6BqO9bD+
6TmUKn3ReOoFdmn9s9TH6rnge57werN1n8xUrftzVsnI6sVd0N0t806ap7ZfHDj0
vD/iTIiFM6dGzjwDZ7kbr7zN5SAWoJxglEUQT40v+z4KD0uG/e0hWB5/9W2BhnZW
9RNsc1Ckb2lDEo1sGBHXwNdAWtmK3cv6+Wbz7HfNSre9LCjqljQ7PSIxmBAt7uiG
ZKtevHK02jOyV9DlIpLT2BSveN2vZGQSZocUviNFdHe0Z+WkRfnP/iX8l6Jd88Tl
KQxzymj3uDGbhw2oMbLOPUH04skQp3viM1aJjnB+vRv2rHeCoLdyfwth3kJ9/d7x
Ir3Fyhvw/VPnjDFuSH5YoeED7GEUlUpZxSZZQ6atQWP1sLsJaD/W7fJooasT4kvH
DrazE9xSm43/Lg4LV9G6IH9j95bwf6CuGSDeA4mDhZCbEJlCAWtIKpDMkn7QGlSL
GG+Ln6cTIOo8GoXrKxH4NB14maoi3K9t0kvodMAQDa2UYl++C+aGm7OV3YTMJlX0
cuOPbchGoeuxhoufNZO5PEdcH2wDa3JSy6NcnJ3/CUlWWvtKSjZ5OVN0De9+2PMh
ie4rVQAczZx9osEKfWmeUfWDStsmriciaNvihR3P7+eoRVfp3ihcYYW4rRarIglK
TMBBsS6wtYlZTrf3AIIIPZA9G86rHlHwtIPKYZ7bh+Wq0YLlL91fsOadiGqq0oKh
mF8+mwP9Cunf3XFKnbGCP+1ihR6gqJOdZ91Bygs5YBce7J0R+Gv6mpMnYYixzAE+
yGZcN7VXPsbIqkqcP2nKn31YMVpQt4VSE41olnmPlvZZTESQkG/rXt+shMdiV3YW
nioxUi/8iQJ8caUE+5kbk5WkpTQxK4Uwy9BiJ5AKlCyldBU7aEBsQB1VBNWK4n53
jWDtTuVxReDVleClsA0Uc+MsoubaPVDh95r1hGnwcfMtkpUthRItEGUVIhZPCBn2
PG0RyXEqOpVRc+pMFquJChotGPNKm+Gwqlx9ZQmfbMwUKlXKtAXx3C0akwyQlacM
MZuzo6lFzmn5LavDPBZ0howwS3cu7mZnuc6YPLcryTpOEB1S5o05DPPXqz/cD8gR
CJkFES1VsEUhdI1RRNidgJv12ofjC9JkTREqeu3VwXfji05e21Ac1Nmeb2MEv1UX
VaUpsblC82i6C5lHyeq7vxhB5NWQyotBD7HsD51Nv8JHnKuF04Qxu7cvPEHllkjv
FF3hXkQqyWyWtENsJpjzrNgWZtLYYnVTdUkWZUJnpThtcfRify+oduQmYGRgXVbr
isuGAWy6NxYzKAdjsw/jbP+1nnIDBakYSy50lYqOc9HgPzCLRgM6tiycnniTTjkZ
ro51TA0TGA4DjwNuiCLoPA6uWvzhy0jMpaOueN5c5qu6ENmrRbcAnsGhSZdru3Zn
uGW3keWSmDWyyP/2hxfez1jGYvfdOA9CNMcRNxVQXJQ4a/CWOQppNyQwok38y2Rq
2ODGeB8Fut9KDvrBhYmhIuustPWJxwEPLzc2XiwB9wGSr1ujS5PqhhPK7LDO2JKA
yW2+UqnPWv85zqUwPh+8mCuibhdgwMJCfLliE++i3KOvZS0RLMQTv3qbpRRdAhyk
FShe10rHZ6fLV1agXweiGDnKko4SfS0/aZtePNHJl+iF24D+O7g2pbLMR/VB9Jxf
08lekQVb/hoxctkIoz++S91LO5fmIFrXJNwV7Z8a6tx6gDTHNrqNeqbG1GP7RW6a
SqNR4oX8aQgj43be8cuo120GPPtpJVb8gYNnYlVTfgNHozuWfLktd8uRb/mjCSs8
90dU07aBEQ+l3XYmBkhqNNEEzzvSNi6OGKe9PMo6/IUM4EPX6XylhoAUZtSmNH6c
0yNptS+HdX49/PAVW2qABBx467CGFccuqwrlZJaSsKBwXX5j774lf63RHP44WCmw
nFtW7s0ebnfsaA/hZGM3ZgaT5vK571d1nI9UtyTgYj5A1eNEmTAd8O5/oNCjVTTQ
M9jKYUsSKBjnFqnlw3VjZ8v78At2mDWswtklsLxm/JGFu1cj/gkADBPulRYVZXGA
QnsWsCsnHylysuHZLXzxy2+q0rzCMQEM5+ML9SgaHs2Tp/Vzr5Ts+nMqEoyH2IWM
Geeu+5RJoI3UdM6lg9vruy6MFuoFulr4uYEjQFphN1MA2sSy/2eEnmXA0gRm0dAx
DbmXAwP1bH0Dq2q+MVU7l/LrJhn8diWOnImt35Awy9lUIySmL8yY428Zp91uJdBp
U5dqC71FPVm82wyID9Ss/Un7debbtgfW0GN1sy4/SO0cs/6GRfYYZQts2Xbo11tr
ONWgR8FHH5339Gj7O9jjGfPEzU6F+ink9fus3on0bxqJqdixj8zXcrvfDe3U21/l
6HhIQOOhWsriznnKpg+TnuB7fK7xR1URSxP8mbDOKiUsSt/1XyGRaYxvT6DJxnCz
OLC9UwVIub9XIXqe1hHylQb9J8XRkRB2qKmLhSRz7VuWijwtIwTEZbl0KVYraxf9
6TlgGU/xC+QLcckiqN4BrGqh6zDTnr8PQTPOQihfz6H+0tunMG5ejuMH2Ypa/ra7
L4N5FnM1cVyUe6Jw8cv07WXRlM3UkHP/gxFr+BgNlZMPXjIGGIR6WbHVlNtVgqGU
rT19pe8Okf+UAvUEKtinatbPc0yDJqUzZfY66/HKj80nIo9zJDqv0FiZ3tBawWpX
rTHIiifVaimI7CU3vN+UNw6OxFyYOnMD7c+sOjE+52GeFjL3miYwmMtLuVOoQ8a2
rbIy9slJTtvpH4PVifYKp4+gaIwh/Mj4w25O7ZN8i+LYUTJIKZP8nivIiErUVR39
B2awpbS529vi7ztI3V6AlB4+++T5VFJnPMXXYuYlPauWpqa53yUZFZW/d6KjCRfD
LWusHII3YrlMDT1NAjYYWG9E/B1usHxR4znpyudduqypskYlkSVfkkDvXLPgTTgn
neuhaiD/xjf7BB0gg1XXvcTXfOZrccQ/zZv3IB4rgOWXiZIhYGy5a2OUVUeOMQ5E
yFl8oy5P4nMwwGQhsEsAVZiezoT0hnd1YcJsi+Tqszq0NvVBQiJQ/y2Dqyu0IGLx
VHfnrWH5R/BxOdGaqM7tfiLPd9JLChMK0NQaYzKvh8DX7RW0zSFESPja3Kz4SXdh
w4dSmeTKlvj0rZ1vy4e3zOcLQejeptThesREFb/uD7SYKYMKK+fCBje+9I5BXJQF
xg6dqOAfe2ihmahchynol60Tk72boyZmP9GbIMytv3qUWMiuXoBJAE1V5IIJl2w6
038olH/pUW7BfBjantchG9+Aef5fnFANHnwVQLhbMLdQiBju1SeElYu4LIef1pwt
euOpLjUNivKw4tMYWH0VMoKNfq0CSCAHeNn93xG1LXq3f0012JZMc2zlmnN97uHg
juTV1/osT6T3fQdl67YoVl5lN6YnnGdtleVmTU/l7SdIe1F7XQI3o2MYLC6np6w/
b3L8wlsFub2+sCTU2/TgIPneKEwocXqXnS9rBVAqGL3i7dVZFuhhPiDt33y0VTZp
tBtafe2z/2m8zr4i5poZYv19aUDrpVnk9tjm6mEm85qfKHGoPFcBNNCBloiWEOGB
sS9xk0xFRnc4CFLOCY1Xn/qCtKVExW6Xp++HRbVUjJvvUSK3EOx28OZ1rcIOnWmO
2BxtIKaWhAr7kn4Kcxj524YHhPkrCLQQh//7UlxBnfz421YaiqKPGAcykGoImnHg
WmhP603LzSThwtLAu8hh3His1dPpUJWHFlApHB5Z5+HK/aFyBpwkttJhwKuYy7ox
0WCYTUMvDw6/1IHWWXu9sGmnSZtykJcE88r8VLXI1KAyMsNFB5aDe0CD9XosZvF2
1jBwp4YtKLeIw0i3muVrXMMFF/qULY8/35N2iI1MrMSGBrENqwqrIHHJyP6OPBvK
YYCgE2wPzfEZg36WEXtUaMaGkoCOhIptbGvJdaxwiZ76t5pEBndwdKV1JsMqm7AF
yszUEexb9p9MMXM5DJVMla++ubr8Big7np7URi988jGn39MwfDq8//XkwY+cB9E7
Oof7MZgO095m33pYuzG5V01ur56JaOPKDrClo7jBK28Tu3M5ZqVCSOf/4Yff6puX
WwvhmFK68W6PiEzWPY+JRtqOXWFUoh/dAIpTkDov4PeTa6UFzkD4BZLOXcggHL3z
yNMGqnIu43zyc9f839P/dXSo6JKn6bt8glPSoaRrsaIEdjE2tmia7hUranUlDdpE
xWrK+PzUKyaIJEpqXFbk5gVREY9K/opgmAjha6Dk8gxGQVfXws0opxa895vZ0ESm
4h8AhIOJYo9MILTaf0xglUwIAIBKqP/pScL7XR2bfrAVlCYyO5pb9APNdQdRQ3Gh
eXzIry5O/a/qykeZbAVeit9VXUlwDJkTH5pkQPdg4ESwwJpIH9grV+x3oVRcLpAR
WQW8PzKlNX1L8si8tpJ1Sf4Yukhfr8dt6/7jBe6Iw9CYJ3QdT0hp3zlqm43ER//E
SrFsFb+LgyajR17f79LrM4OUqzaoWW8TXkEq8W4hjRk+eNFnXJAyZa4FnOQoP9s4
nkb7QCX+nv/IapN5GKnhnVblSS1apvfis2wh4qD39V9xbWRe6qlSeawIon2MoevN
Xvu2gx6duKLN9eCB+KYdhfTUl2KC4JvB4O5pfqhmbQn1qn3ZbgpylWBv6qifsSNS
AIQUrLcGqNAB5HqtlqIPaBZVbx5IWe4jXYyCKflBQjRenJxmgIODMhOBG383CuIW
KqzHrF07WoPR/DkVMXs+z2/AAOd3YOcQ0sqE1AIa3V9V0qE0OkQMjmk1AMi+iUOR
6KhikBCSxarkuFGZ80IunQHwE6+3JyMml+u/SITMyox1Xkz+Nonj3G+zwRsMzelk
mLcilxqwFklmP+GrVjXnt5UojEY5doixm1oBU4tZybEuc004feitSTlEmijJV+s0
PdJD+ufJ1uVv/IkE2eQLCY1Z/eOxbOkQcW21vpEEWv75VlknG56SASG2qmwIIFU2
rVtYIEfHTBuPg8eLjajZshcVxGAFr6AXxnThJnnrNwsQ6lEbtuXo2uNQQ9oD4LaE
a8DM3JocNjeVuF39iLoYttdYOL4ttzXXcoxqXwBejSCujEpTf7IMy7yF75UTaVZG
LcdceK0Rm/So8kMzg810VMxF+Sd45EXU1zKEnIYkrcPpxfik5tLKqbkiKAosX71p
3XR08Lp2VvbP0kQ7HWADDfZsFZTcyOifLPZFB/X4DelwMhOYTj7LpNDmtG7juZmo
CKUiYA5nAuoQPknwmXBlp4YbQuvCdATpYKPatetqjVkUEfZSU9KSCAVRljIYrRHm
YmD5AprUlAYD7pweYF5lFQ1aO8jr1lvyJc4ytEfYRR7dj9fCXRevwMkZTTF5N94a
TrNoMHjHwvxtjbkOPs9z8F/4QWvaxbexL2VWh7XU+O3Q+y5Px66vAlzL6srNpK/m
lylRuAfaRTYsloQJ3c5ssTAT/BcfsMyq1dYbIAssU7m6Bw2M6LedrNOMNx7H/Kbe
H39LSOv1GDQUWHPzweM/mcxfMHcifQuCpneU42oXMIW2Jbzs2UmxvLacqZyLkA0x
ZTps9X0Ic7kTyV+UwLSL4uNoFvkn81ujZeqxqdAT8DfmlGYo8dVm2QybRZMV4n+0
nHrs2/Ph4nf48OmjcO3bJO90o0dR+B5nvhJeulNPNTI9x3o4kHHr5rhJaXf2Rh7v
FkCCZJDBsqEXJ3Cqx4FgBA==
`pragma protect end_protected
