// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V+HHEuM1txvfwqqTRRDqrw3zlSyyJKQ6ejpxZX0AyfEOzZt42jW7S8xGujAB8hmS
rqu7MYRFmoTHD+gqzno4YKdcjiStxt5Bm7bUOROxBhMDGRu9gkpHdUZVni3OE8UG
pcTABgeBMDA3Q8qYUpWvyAE0REqDu3DhfdROL7DpLmo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4176)
n7iVjlSNkQuoB433tTNTNvtX3H3RMnDCTeVU3xYxQjwEZUFzy9/g10fIDOaKo/1U
kdpZyY05xySmLj0b1tKudO/VL4KGshARa2814Jcfn7YwnjNP4Zupp/qCLq5BkiqW
40c5HxugYl7POUmLo2to54Z1fDHwGxb2n8ByG4V6wctOy5I1rz+yuqu1pvQu4uk2
DSObEKICAuDdAhwIYctLClcxiDoX2M22vd5VEBOmErKpX5AkvZq8Me4x+pPMQEEG
TbuKPxNZB4IUen4FSV+PZuvNVPIfk/AUb2V/UyTS1MDFOTGs3Cgj+DC8ynxk0UU8
TIDdlu20sUhg3MQTMxtPSycThCfERbBpPZkU/MQoNy3CdxJnpxqJ81np3H7sdnW0
b3POo9Gxl0Bm1KRFH2U6vVpUblEfAB0/A7ek97a1ScONC/Bp0QvdNVRyFqeLlFqO
781g0JzGfyFXbI61pOgj0e4Cd87vUp/lA/dSXaAp8AEXOpTtSli/cwVUEFNLUXiy
aurVF/RbDgTeTQ0+zxjGZrgU948/hwCwUcobJtyKc+D3WHMhlvpAl1FQBM9Owj0k
Wx713MkN0mPs6AdIFHxYJFSdfCKdNaRlrpd5Pxt4Sys2r8FQSQri9Q3rxnCWgGZS
XDMmj+yRwG6oUJsc7/4/bfKXSZoPANLamAvD2TsOLtE4ru7gs71IA/O+WlAMwugE
/uBDm2sZ0HTpajcJcr8ub/9M5yDZVBEmH15tD4ugsz2Voy2oLOMydlVoEvrujfXH
wc+z8zt4of4H907hj0C8pTNLdLuPAWNKtGy2A/KxuTdxEfITKZ3whzb5OEwRKxUr
WDFTap+n1L7tX6QqqMZMA9MkTA7VOFF8ntB8SXnCCLsZ+ewgl4j6Ncku9T3fMdxf
jHxenEaq7CzbbAcKlHkPGUrY+TyTXfjmjBVKAC4TEssRdNkiurw9Bcpa+HVWYeWB
yfHIowdnag/W1tJ23IGClMsjQrM4XHcpVtH6tFnptrluTF2T9nfvkcWlV8BoO/xm
VLhLJceGfg8IKNjbJgt8ZXMzG5sVDNwBVrYnmou75d5ODZxxI2B/eLMMgR82x0Q4
59sMRz6USm9ByVL5Fi6P9kvbC+kFg8zhwyutJ6wUjPp42bqsfo3/ptMQKsFop6P+
fxNxUU9KF/WoI/4s1h73uETYJZE7cEMNTJl6hGPnIENhXuAsGt+X90I7rbsl38lW
jglfkrGIYcC/rFAgKuDKqYZo+QkW+Sj5mO12iDCW82fzqGStfVtWLzsDGpfgK5G+
QhprOOpYjbe+KGgR3cdJm4K4hQTRKUuKqqjLBOAC4iCnQIWhhHQ1KMA7Ww46mpbO
/LepknDZVmYZCADea2cxjpOPeucq9spD4iiVC6PBzGiua6sCtIkYomJ2uVzLk8oI
78kvQiKWgv24hNS+G9eCC5U+vYirh36HxkLpA5BFm1MgSLi6XdzAV6Q80IioVzIv
HCA7EGELLiE+JiCYtTeXphzyjdQIyp+hRo38mBFraC2ru69DPgssvPKx0s1RF3dY
PvXXV/j4SWiwaCx3VhUVTJsdzAiQHN93+EEQd2XyfO3geS5hxFW/MekZ7GvN0jAN
ZCeOjGOtCUCkpM1TC2UshZCbufpMP+uU28LNcEzFk+0Viy7hlbFb4NMP5vgi0pqL
J9HseH2i3O3LwjroAZAt3K8rR3OIG90iRy2ZZNuYI699FOziWmFN52irLhRDN91k
b1lRr+FgimwLsYjAqQmgdYCDXfbcfkDpPcCmS7CIPZxmmgm1zUWLH4RrredSaaCn
QW7X0h+kgyOqjbSiQwK2AfXulBnl48TxnEMSpOLjCfGnqvWTU4FYC2otQTwzywZR
Hi7+2vq1b1EE4Ow2YkgtdF1sa3QQOWJDWFE1vcBmUPjILq+kZjLXoyNNnjenqSbe
i5/fEHyT/uxwI5R1Xo++Jjx1tadDAWsWKrqC0SSeANCyCRaF+PmIedEtUPue1lG5
AcgJWtW2+zhL5vpHjHJa4xsQ+gzaoh6nqSQYpbNGKNPkxCEGX6H0K0S2V7kmyY3+
TdwxXJ3yr6NhsbVuMp4YLRdYk3eqrBLr6L8nJU3IMEKy8+XrGslxMsi0UU1rinkX
12Qq5scYP8LPXQEM6+p5+r9tdmgcLbPStn8X37AZ4diD9c5trnn2/hvWy5vhj/SB
q/evJjKcb7VF0DLoKXJH5OTYeFQBR6vT7ySAUJNgcuPUDHg+gDx3cnhNM/NC1KDO
k0ZP4n1WtrvNMSVIfjcZAg9f7bRA3kKxD+cFHF+Kd1muzZDqlVF3svmH+Gldro4O
rBeGht3D3iIxgjaz3zbTmMNpjoYb5PpaPMrvKtnyORwDUgJiHyOXvsDh3Iue0W/v
CyhZJpYlXKIlpGfWPSDDNn6181aPuv3JqQ9Ur6hd+RG7oJiSyfYTObHAOZ6KT08t
ZDJEhJHffM2b+bvwkBJc0Ls5cW4/KC3i++hS7V/TF8HNjn5R3AdPprAoEGjqrgFn
ChunvuYU62qSabpS2HICLB8df5UXjh0HdZc65Cbuvkqvq+ja7z/yJHTXNUw0QkyF
6BV37lpruWaxYJbB5tmGZbYxiTbQEsevGp7H0A2WST/016k28fHBaaWfXggY8E6+
psAs4sSsQTD22suzpv5CRjafGnsa6FElFlyV1In2ctggJk5cNcwVP0godVE5e8E2
co+XQClKMcME5xY+HXs7DK/IBtp2YKCGlUc0vD11zuL29nqWSwav6g6PZII7TB0q
K6VLZtZXstSx65gSdUSf1mwdMDHXDJPc1+gLlhIm3nZ27TWZW26SdmLuttH3UGrL
+LSc7sDTkQf8hrMzZ3NegD1L+9n+bCa3XpI8dlyCYUlNK2Nu/BuDfPhgQ2iJiVMe
sMs+8c0t0N899cECVGkYWWBODjlxFt1UWiSNwKOHKQCPg5CkFANjWwOVkwYMG9y9
Dqs4LI7XKREh4T7K1qSe8eraORuYAYhuzZ2AwmwUYM3+jo6O9LOn5yh3guGobF6I
ATsDyf1jUDrq7tDUzQb4DFeUAJUZrhMunq0oMBrQPpnO8vZVQYQxQj7C8yR3UO2t
tyLps+E3Ba8pIVwclE1Q4nOyXZDzHnDHTaMf/InHvu13lJJDQoY4U5ttkEOUJGb2
Zs4S0kHu+sOXw+P3InChy0fvXpB4n9zoSkc6bk4WH/q5KtEryKnPJ0EUPUI9mD9E
i2S6YANgA6ioS0tMPehQHzkaVELXVACXMNRPwn9rFCuS06Fg5jDWx01gTWaVt+uh
TcmizobN4XZc6FnDa0d1K69eOhHI4YcxdOKrPSvn65WRKy/VZytEFa//7Ax05qYa
0ZUufrzS67lHOSFrqavTFWyxT0oNIu7UmvOPK2Mp1i/PMY94/7D0+E1AyFhJXJ4a
Yx7dw3iV2i2QXkykglSLgTLsMSHNO3WPqn8516v4ottGV+OhVPdbsXjKOYCT6Rcn
428QiyEPBe4DZzhnw8YFRUux8QqjYavp/pjTvZwrgvRoztwXuuti7U8mwtKtsUik
T5tS6WVmHz2K6RPjs0QnMzEEUxgVlku1nn+mXRAa45nOJVJGJB4wxNRF3vu3xKhc
j7UgTGjMrJh0BE4lL+yqMc1pfgHKi4S8xB4P1oPGxGztjFWgRXG/w4LFeff7zQOt
Gvjl/7hTPP54GGmpYm8tejj2orJXhJ0TDeLjWv1kQczDI6Y1I7gskHzjYjHSbVZ+
ovTAO+Zrdg7IJG3MYEQFAEbkwMF3KQlNDmpKmyBTpWZ0iy+3JWmT3KlECa9IndGo
fLJvkQ+krFGhwTJ0uGPX4GaWzFK0KcrtLxEzDM9DKF46kCDl0CJ4rfsR47GbE0bQ
P658ne+K+eg0ziYvAlbY3SuOQVpPTKJExzgJeSI5041iUgJ2x1nXUpS7NQWPS/ji
YAzeC0Eo1zOrcjrnhIa/beeq3axWOrL7Mm5RY/xmxcEwGc7wsFa3kSNOPLiHPO0U
ICEPHmlWO4h1aYt3v7E3JMt3CTJdoecDbtL78biVbtbZy9RuKxUgsTa9Y9BBMyOr
ORZMufzXD+fSB6ifTQZCv1HKaT/LXqnw7KTA0W4F5zW4LJKUfRByDQAzJW0kas/6
EI6p2qmb8LwC54CY1SN/OQB/tRAMBawZrXKe45FBQ0yG8Ak0Y22yBPEG2HA6V61p
cvgtsGwUbVOvXEuqgu3kRP8ETcFxPvE8ggHgy8w8PV27blBkpoN6FB8TwoX5RHpO
XRkxq99yabSWgom5DuP2n4R8wSaXXZcgpYF5tUsOgCnQMHQUY0RZVyfKQmXd2GV2
yDrZELvpqSngimzWQ/435eV6m+9OagHYCKr2ZvNcexWEYXnb9lv79nNLJq9lM6c/
x3s9MIiiVqT0WZbVUWtYSHT7syuGXouhvUNXBk3vF62I1W5N9UBHXHmHBjUgLfQG
72NTuCZMd8brqm3cdEeD2R4Vc5ZLh+EIPy++YvZiIPaTMpDu/V90n9J1YI0Alrf2
e89k+tfcuZyXffK3inRmBPlnE0rgM0NP2FtZuQwCpMGADgGldZEuHgBUvt6CoLuB
pCyBZegPp0DEyDtWU0Qd0i8ZkCdHN88B9EEfiX1cHlGRryZxqP/0hO28VTn3D+6F
eFGAGfWCCPSJXBjP+DqoQa4GbyFnzLFeGg4R6sjVAa7bsBI12Mo9kVj2R4ombFsL
eEdl/jmvouRmngfEr+894mdEN4taP3YIVXh9p03bbXyOlcs97vkk727ATwJoNCY4
gCcClLD4qrOJcfNqSC/OujKOuHrMzARKSflYsz2ReiuLpxabsRdaHcuUCvs1edvQ
x2DddIH7UB0Xq8SDw/F51+kWG0rLEjf8InWRKNJ1jRvrrqJo3BOWLw1c36esEsXv
7rkq/KWofUiy7xH4NEuwzoSLU/wq2Cx9j9NpZaUuIwd+VfN5PRCe7fR26Ug81jS1
h0tnk0U0AUuUP4GkTAI+KKqLynH38Fhc/g1O6VN8pwExwzSQNTvNAcHMTK12kc9N
amJEP7TKg4LiLaY6xVPfXK9Vj49WCYp/BRBru8X6tVslcafCcfv3lW0MgiI7QLkk
uHwqSy5C/jsnEO5et+tOslO/bD/cPc9GZAhS6oD+rZOdiyJ+G39QL20Yfo17YiGv
6Mk/qnZp6UsBT8HRXb43ZP2GoCGWNoNUriccXWS0tv2xiHQRKojLntkpA1XPfsic
/GfJUrqy8SJnEjO5/35sXCtIdY5hnue4raB0eb0enLy46AaD07kJzzHHKy1A4W6w
HV5MYIKj7V9DyqPpY81VVId7a4n1TQ38l6kbFdSv5UXFQ/UrthrFJvi2+P1ihTzp
jBs6Ejk4X8ESJTVbIk7XvctXz4itdCvjNO43XyT/cCRZcsR0sTM58hRU9ZIZDUI9
kSG21gZR7P+T9nip273RrM48iuSHkgZooKkxt14nhJ5shKLU8Dfb/uhvOczFk+eC
g+tsuDQw35qN7bypGPyIVQVsUw5lYgT0A1DHrRWy/ThFCXawKlR7T6huBi1jlDN5
ZCb/iHzLD/amRr0/myNP+AGb4b4Mi1+ZbpF//QKzVAnxL2m36+Xc+lONfdFOja4X
`pragma protect end_protected
