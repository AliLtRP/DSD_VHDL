// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JdOwDG6GSCfr3DTGxkFi+UjavNEQ72EFTNOERjgADk5lwsA/r/XRHzTodDIWDInE
qGDCovuVBnQwgrlY2NHXTrXSSB09w9xY44wBbjBJ2tGKu0efC4g/6auTNz01wt77
+540Rs9Yhd/hgBNKjCnykUNuCOibFX4AIWbQmdx4tYE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 52032)
1j1muYPuVobnTiS4Nc1i4EO5nxZqxxZRtYcZzCN/5sKH15KHtbMdOxuyVUKT8w9S
rntGdNXjpjGB40XGcNwvBOX9BW0IXSXx2kmSVT3wcz1cZlak10PpFr0U1/3cNdoD
vIMXt5nMdiYxa7eDOYBHrTDWLLcnIeFEHGiVgjSB8c3/5Lbq9s7zezwixy7LqxuZ
Qw113Dsb20auWhN/wln00lLWWiD0PxmQp8D3j8GeDl6wGe+n1H4/wnby85oSfOMd
hHKMkjyH4jj019DnFZjFY/ezx15xp0Hqzl4jeup6bI+NtPzu3XJbGNyDbS7RGcH3
LQphbKaiCiAioEUEBy98pq6rhLoOj12otktIiXEjQKY33sR/HlVO2BYU1IEK+Mmx
sywaSb+HqwVK3jSmQz+lxrR4bdTjy89uOwiWKzpwrVEQIKaAh9uzmYBOlohFVQvy
h0nDRZ0he37KiHH4PbgwhyXqGUrhWTBrfYzobTtqAC50bbsiAvmiA6Ow0qd+FqdA
olJl8zc/mw04hUQOBAovW7pmqX3yERhNdoe2v7sMlVEmun+pVOdVhi9PmSWUTf7J
e9vnOcWivbovqO/vSMXdhojZr9Zmedlv1qs/c4YqkOmi2MTfHfrAy/cYpGsYZQk/
6oG+wuUzrETpRDJIwMiohJb+r/EN4qeC8C2GlsJlVA7xglqNTpHpqio0ZNB8dSsp
XKjVN746Yf+B/VtSRhS7Z7QVGjjhVSZf9AkbC8je54BVqLxOwEIC+Q3PqGPv3QF4
is5znOYai1kTttq70xBeoh4fAASt25EYXjBnZ1rsJYqYzbZ82O2PRrvvG8cAX96z
phCBCvs2VGFjU5792lLszyEX1BI21UbcLOctDze3nRcPR49RsTlo85to//GH+zJN
spfUbIs4B0jtH0Mzgnm/gTd8KBigOc8PRAzZUisruk/GQPGQ0RJS272sEo7Vequc
pxrFyB+2cg2hPbxgLyQQLdzO9mjjdLIE91Bs47eDXQQBdfOaZEuiOOhgAyGVyzDf
uIrKh+CB/3YymtZqQOFF7kf2oziSc2DP+SGK8p1dVb/Dqw/b5FWOK9P/nQuEy4Lw
01wluafxCvAaOFesiG5zC7zLWdj16T6kBPcpL67/Gwe5jGUbJHT4AQuadmlQXG0R
NMG4JNMjDsfZL/e+V4Ij1uJr1EMqtv1FgvpoD3q/guSBL1PmiHnLn6b4gI/P5+DM
4ConJ9HPsy/IhFFAQCX1r8CCPJ+aVyvFw/N/4qHsnEjo6O5jR+CqKQzT6gCBAKs6
aW4rWMP3uJfKMhkNKUiLHfhcmeo6RK3l87HN3n0hV819mivpUHpPe4zF6HF5V8jI
i5It097j0Uc3ifFBNqaETvumi4N4G3UD1wKttD3bLbPZW13X6xzBN7U8+C8AWKGW
P51hzcsc48Q0VtYXaBh/Bpg+Y/WvlEktVv80H/PigqAdYVFcA1xA8m+RLZ405HWl
Wu6RYu7GozWHyEa3iGzGFvdLykclDXedOfHgkwfxob+LfnnSz2V+MLrR9pf4cNcH
sSCkE+y5vo1PKNwGN8bzFWhIV2ca66j5f9NZ8VcFM4x4KEYSLolZC9Po91Clwym3
SVh0QkykBAVYHn1BUQkK57W+ymH111ryy/bTXgYgCYAn0vrjjg8r1CfMQHO7doMT
ACSmsQJjQMvWffBbdoUWaHzxBZ/n17menANwKdAdcs1riAB5VEDVlErACaPfzqqj
UuHTuEGafhrojETQPuZw6lHTPjiOTj4SUXuE/KUBwd7D+sPUsDyBV/cXKMRo5aUt
3LTfH7GEGDhblIufXt/tFCkbDW44QnpBw1KGc56h46CaQZsbgMjka5hilN6DvfFn
4imUbYCyiUPB2DYkLKZqs07JfOG7GhyEV5JuBmtMsZYah9XrAC7dXGfr3Uz5mz1P
Rs2oeOWeCMGg9R0/+nCU7fH1PknHrzffwUA7UynkAX4EZJOyZJGI1TMf2OZu8ZXO
c3ePSKXv5R5gJgDqJ3TndxhFkbeHUuHpQ8BVinQ/cR0hQE4a0yZ1eecsMD5tH35M
t8IXrNa8sMW60bW2RP6/SwJ8nFKLv8vky3zIk2a+sx9Y8SDURnlx9t1b9eAErbXB
0wmYdirUPE4qgf/zBiqJGzcBqAV9wU8B4s+ugLvJ3t78o3RrqT/xga1bwYMB2Yxg
Munz8pIbjSHiH6ChlEdudWpP4hVWsxSnaBUCYQTeQRZEox3LEMi+3UDT6zEoRfw9
MVYnl4AKmP/JgFKgpWe06pZg/1FTZDG9SZtkgcv57Dbfq2wvYoqlMsbT25BeC/RE
YzYk7LRAbaeUpSXP+KVXjsAESvf8Ks0ZXGWLtVxIO7DgVhUv2hplFjboZrTaWGus
iOo7oJO8Jos/X8IwCc1dc5LVyCJtn/J9f1PAoR5bUiH4PrEWBSwLAg6wLNOQ9VbJ
e8nWg2q6PXrDM1hsCQBJd942XB+RKpPCQ7ifxvOxYVlGFRbFFcoo7ZAfnUphouxJ
smo1kq5z4it63n/0kmRzk75GylyT+DpP4g0lRrjnzRCaqKPBEBw6kJK1vaSKJxmh
GY5QSMZ1xT3DgoC/2oQQ53iy8EbKsJIoy215nwyG18eE4I3XfTr9bZlJPsBSXLmj
T3BEmE2ahkxBqSbcFUX+rJPAUmAzbMFV82Ru6iciMGYq3rl6nf99UNF5gBamOZCg
hLlmGcu7nKD477mVJSI6RW78DclPYGa1NjB+n5znKCqYvyQHhrbSmu0FvXFKClt1
4XDc5ZS3IGdRmShC30RTUc0YKpBqzSo6rNDTAezJQdr//pU6/xMdGF5EOsNwZAeb
TCVJ325j9SZMCukhcy9LIDl5vGBnpgdWKFybV0TonRzfkz8fPD4Hz4Z9rlnMyPA0
YBghK5mts/QFSY4r8cb1T77VfNDAFhrKpbD5SQblVadFp7OLZ3OfwHHqiNrtfrAD
7dDV0YmxLwgdvslNGgjDtd8Xp3iC4uz52uet9dOIUgjhwE2X7s1/nNXTKmJPet8d
Fw83i9zxpo1bmN1Q/bVkeA2JSducvCFXMR1pCoQBYAjwRA8PublzYOwud01HB0nn
5MUtjuHJ1WIBEour1dJ6yVcEaVBKyuFg0oVhuaL8lvpTpW1fGbPzEPNh5XVpKfUs
4vINgxNtqyaPbAJbibwTXM2OHuqbyq7GMZ/cPPGhe22VZywqHZoHBBPGRfpHHkbv
mwn5Mx0C82d34a3arIInhdJf+UB6c4LWfIJ9xLTbkQBMYQy0smcvuPd6KEDVypvB
QJRzJTz1zI9jfgqxqgo2pY5hXZZZN7ppg3HgF0IHTFsaUBD/+jnMLn2cXgBQ8BBB
4J2yOr0qlRaEFHM5kQMugZEmTn+/A14VqSKewuQ4uLVVECc5Lx3wtM1W82ZH069v
KZfOy5CRnab3B4yAnqPUQ7rYQgbXTu2P+/D34U9WQeGzbwAy9XBrpVrB4MUVqA7y
yuJa5zmRDHzUlEwmUCxvDDgAWnvFxorasv4SfdSi37Hz/Tr0Qnh1GnNo/FsjxXAI
RpKk+Jl2ntzr0SKSIwTE0xcwY8ENa2c6OeqfE2j8/cKoMfX6DPAhxoonlFe3ipRx
hWLdOR+s9V4stEQTCU0mMUGWIp5bgHni2BQymFZGdfUeAjMdEhNdg4drRh4nD7Ae
CkIzKDoenV2WfoK/fq2jfmvnZGG6NJLrOgCRoDdE/JJBBZleqvCczhG/jDJAO4Ri
V5LFwrmSVXHnzaUHkn8Q93TlcoDLN+vfe6551a0CAslpfFHtzFJEpNIL5ZYL+z+P
NiHJyi/8OV0ULOCPAc3JZqjNWeSuOBpPerRzIsC5spFdjLb+wWItB4yaVZMKBf9U
LA9+sXjoYIyv8AlQ4YLdmQ9fF2WKRTNdm63GlOeOxPsdUBIv9JXe645zWupH+QZH
C9bCm1b3GyY05tkqEnZesAwEoKCdEdn1x3EuZ6oNgrL3r4OypFGUNWplRTX3cCMd
hd3/BLdU6R7FO7MKoLV1UDCsmYAXE4YS+oJRlOaG2y8S67EW2NLzLCq4yeXwis41
4wuGYDPIk7VF1qZ3CBXkzwNPcmDt/bwMp7ThO3ET76KMrt23OdZ0gT8sJSj3hksi
O8GsQyGpAiOj+l19iEjs2LVJuDdkYDlM3BYqxbnccQLESs1xEKcG5rG31MmAPuMe
sgIlWkl66rYsrWE0zHB77a2K84mAqAQW4d8ESDYzSyglqrNnp/+DFxEXHvyf0/nq
gr1ql6OSDL2LClbcWIFbIbLxlRpnvpYzc2wuHAtY7oIyuOlJqUcY6wNzFPcU450v
fmV6Rjyd6HcpFScWOaJJOATiDjWaG9xZZA4T5GuAhu4hc//6F4p4nGsBero84WD4
3/KS4fQNT0vIVtR78nSy4Vrz16ixJa1MGukyLxAzGz+Rj9hvCneyOrt8cb8g0wmo
aekhiwqIm2g0JgqwzvzOkZ0o6pYRs4xNVBY3N/18sLxUAkGhi2CinQ9M//AqJnaO
Bg1ZdL82EMnjEFZqTgWZqFrfK2lVPXgNb9QbU104Nwfy7CJWVa2TTw41O8MXZFXR
qwQPQOwefN6qTGX+FjdqLDR5uhfYmHAlUNRv+L4D6ymBERWi43lj0wzT/KCfzuhq
VkXg3YWZVcIGZSwu7qcFKNTia43/no3ZrZZ0+u6BwDVnAcvrPLpdlOGa6e0cHW12
ock7OWAMktWDXw+XFJYZ40EoMG+uWQcbkJks2jIewuoVZstYnVOUN7qa+mWPrc/I
Qwt2yCC7eLJHMK7Ekozhzan4f6B1+wWZAB9yh6xHUmsS687voiLgWvgcIZOUKAHR
1qMHmZowTB0tsRG+DSTA8YsWr0cYD5mrpDwNm1LuLCsY2EQlIyg4ev2rXAHpAmbS
aKVjkzOoGBIVeboNf8hgyfrBSIwUFcwKQCCgtzrs0D3ymynnBcJ6fi6qdvfj0d59
k+BpGzFuQ/bXvL70NK+hXv1xgzKxd+6ZvIvQIsnaDzCBTg1kw97gRVpOTKhdp5+T
SbKb2rCiIn9ye5LnGWYhwInvJUL1r/v0G5h/TJBUepkTmSurjdg/FqeeEXwjSkty
D9pDrlVj5TCz6UHgoy18Tbf3RXQ5PabHj9mCK8Hh3epf8UYbNhBU14oGQA2iBVDm
jft+/6hZeKK1i9DN0zGNJx2YGX92x83bPqykw0mYOlGVUSBsW7DNDN+3iNLW/vUc
ljcHfW1SgVkp7zv4fyWV9cMFS24ErevT/a7hGgz9E9EuycPpfN2svLFs3Ux6GmBr
r8fv6zWig89rlJUnUoAhMUxt+kekjV+pQ7c+t9rLn4FH/V4O5DSAKkoQN3JWuLc1
BQM3vrCHvkkup/5bVtGLIn7wmGA9dqHiFGiiAxmx7KEu+LgQCYWQ/6IQi0NV3dvt
VYihDIp2MeJ6hWHBwgvsq/Sb7sRvHjpcqo6LxG5+QskXlxCI6Qp+rpGVN4IudaWC
U4cjkOeUVkX9rY4434s8VQdjEez8+x5sXngZW4lVTLCOhsEZl7ztDw2kEZD6Vl8G
QjaWejxW6IqNnjBbQ3A2zjgAEAdZZRkiT0yDwNr/M5kdkrz5i3zFflayQdLzer5r
jxKjVNZ+Afbn3SJZ/qOC31BN8JjnKQpJzITVxsBPMrhVJPCmAf7KXRx5VggxBYn6
qAMIoYorYMBvdUTeAsfbM5g0LgX7Pdd3WU+llddxO1KXZ3RzwVFWB00CNMHFCz7j
75eR4Gcpfipmh0fWtxvkJSPRrPQmtElzYo4Ltv54/f9wsBKEzerPtFXEjlYnHI/l
HZNrGtxRXAgumINjWk5eegUQjtbcv/F6kQ8WgrvPU+IZ5XdjnMKYuTAgvJocHS2N
rsMyX9+3Cr+njnK8oUKRvFb/t+ln5Nt2jeJZJfwqQ/fpvHjcXMHl6I5HEiCMVHYR
cyZipK+t3fuSgWxAfuRrSHwyezcgPZJsHu9r/dDubFQ0B6rqmq0rv5ym4EZciycH
es5CSTJHuoO9JsNgT4tiGya6zbVeV2+AR6rit5IwZ+ibc+1fk0RtOqSyKFDORncD
FfI+felYFTgrIrwisKaVOwrv0/7LJ8I1DaNW0c/HRKCc17hOiBzS/I9blF3VYvTS
5VVyGTrkA+zuNNKH0ZgN4A9qmYBYkMVHqwvQtMuTe4dh4l3scMtFw8Ki/NTHTMdw
f0opNuZzLsH0Nb+fksmC50xdtoz7Ain3BOM1cZPdYZCrO79KMguoTh8gYGWK4lZx
H5/Gs6IhYMD417TRduKgzuqlJkGx1NjiH4iebnYkgP7y0tLQSLsx9CvME5q3uZfD
IvnPE7flYAPhA8tfJKRiq1RgSflqIH/MIbEvcOf5PlFR3AgbZzatw8P4CTCeHcAT
UY2o5kvz64dHls7Wz+3VWxbq7+vk0eiT8Dy/ifFAbcoPAwszQbc3MDSCCuTkxO9d
nFfehGTJUSgpa4gxNEQe4BJ3yZ306anIubysKlH8dAUeuUEovHj7n1XsnxMEJoov
g/naOzkjgvOkprw9UBXr+NDqPeb85pDktQyr1gKuXMQyW6CTjaoAMEgoRUhOa9Wt
urqmwykqvyR2AS8H0NcDDO2BPWhhmWfcGxUnTHOeehw9Q1Z/FQf4JPNuLBavjgA4
bKXp0CKs6//rucw7HRCbivA2D6abW7iSPZf+pUrvFy0ke/BcVNvaCvtjLiB5LwUU
1/JlwQzOr3aKmfEgV+/qLxOv4QBdjsjw2kRJP3zj+FlTNKqneNFfuIEY0XBeIupk
9PWpJS0Ohn8zdIxaEWrlyIoTgGfH/cAMExX3F9NQfo/rWgzSO2Jsoe+LOpg+hLIt
9ZWjjMUiqDkzx25iROIjO5kgngYTGT2SycVVd+nT1nHX9dyYek4byoAlWm0rMeiF
5w2qZXyx6236jaiRoPRDLLuWh9HiQEtCzzpmbsyCCKZYXHsuk2NuINSjWE2n+ll1
oqynB53p4O5r4t+OmuwnI0hERdzq08ql13dSFG3JKY9Vt0hC2fKLLsCp4/lYtGBN
L05LjWxWYk4VsmEJCzTHz3KRO7ONCq6aNCvt8qW4JXePrSLRZpuhhnBJlnYRVUYX
Liu3Axb4pX9VuTqnLiOIIHe0k2569+MsQjhb6TOvnCEWMxlUstVPRpNQ6GnIQh2s
n3OW/2GZfcRnWl665HOPH9byEgNBeRKHM6WjAILpjSdmhIIE9t34ljr+uRQ1zErt
y+Z3BRWDpM6h5nXSo3HhgNvPElLeVVrgsM9Oyhuo/6qrgH3EtQbBWmkxll+6oYhj
WuiDHXLxW2axBCf7i/BXOP97ZFUu4K0JxkpTndywYuJ0I7oRRQ7DPpEaPK+GSMot
e2/h7feDwRHdIgJZGZaV0L33a/iaJ/FuC8PF06GLxFIVxrLzmDxrbGQ9/uXqs2XS
NSFOVcKnEW+yZl3uvOv51xMpQGhsxp1XV2jGJPCTRA2hB4/h28JS4RP0e9xtWWs/
8p3nbeo+EpNOEmEt+S/zBDFJV3UhDKZaJXsFD58TjjF5WfFNv4gTszh6H8rtUURp
KqLmb4twFWq0VVkJ986mMxnI+gWtSe0JXT2LCSBsCrQEUPmzzUHyyRbaM91aNU42
Y51YUxhZTgNHV88N5WS/lUJdEmoLHs+qHXzm4rIWL4meS+YiBxx581+IUP3GzpkW
8OP3XQmdbfrMak4HOVqcODWnRFCPzRyy5cC9bKqvhuoXo82Zcym6mlb8AMwc5ZDD
Ys1WpG9KB8FB5VJ2E1RljB6281O0GFwBQN51Odmyh58H1x9472tbJe7B8wqN2dsT
t7dXoUOGQJVj0gdvGCxQERY/XlYRj6r8hEMT+DkeGaDMcH8ByQVmbV2OqPvSpIrC
PXEWS96OftNLPAdfpaciX60nMFgIeqCOODwIcKni/k/WO+H5mKWqjlUIwpiRPaij
z6FK7j0SDcmgtIV9ZA6x36uRV4ePImhDjHoY0iuhgdBwxbcr0AfIrxROnC1HWHv+
misNzlXPiu1rPT8p3QHX8yiFTT0BFjCbS1fYUygqi84HC3al+OIeXhBmnBG/EiT1
6VqBokla1+8RHr8owNF9xODeMarcFMcSWtmqqByhyxugsnCCrbGUQPHcnRVr+E5k
4r9L9w38uTTVEOL56P9XrO9vdXFcbAUFYA6t5lNlj99m0T/tiNkO72+wguj/tOiW
hEe4WftNSmiAkU2InuiznvttRYScxTmVMDzg/GSXeK3GUH4prCXgK51Ryw22nqVW
DgdxBjTbF2UfdovUndDobdXxasCnlmTHuw2nXph/RlvDIkzeWA01Ivb8NRiMubCx
bvwVc3/ZF9KjEmxS6u6dXsbe8fURGUEQmgjmF6dl92LysqPSTvq4QvfAwZLQd4aQ
52FoYN+77GrUBmLw5TaQJqDZ35dX2ISTc8wy7SEW3UjgFYZ6EJdhrqE2esKHkyil
teDj6SAGh6MJSKA5Boros5eU6e+mhV4bxUFRN/6ktCJ5WPk1twc8JFvcLCEdV8Co
KV8lD2X0BbeqWmW2Q2Cuwjj72oHOHjLFmYy0v6lwEajpgyvxF6alvZcyx/AzQZxl
VB/wwLZIAZ0xl9pWbLP0fMT391/EBld2yG7DpfffGF0m/rJLYDBBCTkOBqOQeW1Q
OzNnaYYlJu7nUmWP28DykbDepg2idTk//sKCXIuxze+pjcSN0FX/aqV0MvkIErAf
KvjUTyhMTaxcR0V193Kd3Ha7evOqS3ISehbgarsDzuU2/i+L97p528bEdMg8q3+Q
Di4g0ZUFz1HgzwTaNY/FRZR4YxXPs4eoapTIEyTS5DUQUKmFZuXbPogvT1iXErFe
sxd47FBjoPfA13KbYm5gMmKVAVOvjEUrrRMylqVnO9ni0QqrOLqJEabPBbl5KkNJ
OjYuv35ctayJ3Zs0Ahc6In3WL/rh/QxgA1v8ZBUsg/cqYHLC0GnjZDMJP4OlyjWt
74M8r3qV1WP1g6uMXsQH0nwzjlqTf6Vl/TgMj7DKSWn3tAzAENJPr+u12leyONiI
Oqns7+6KxGIBa42KqOnUO9sekdyCqqswfRCLRD/zRtfEAvnDnmNHBcX4LGvRtUYl
n9UdRBDesAAhPaO4ceV7MOl2J38TTUqKjImXgrG3qCYRujE/cdb0Jkc2ub+oLEWR
xtoH8QxLWjK3s1A0/quZzAtZDdgJMF+p63JVIdtxuJWZFzL7Tw8V5ZgurTyq4j3m
TGpatHpcJTm7m3L+8a7PnNRhayyLLDQukB0WWXY8KGxKhYtL+hTALoG1Ogq8ds5X
TRCDaPDDhxEs5LwG/RlQnb74IR8rAxHAP0sXVFHy4vUdkBubtFUdCKmIquyM/H91
iDpF8tf7+JBMdj2Xm6/60aHPVtzXt9J5tgtqJUpScJyg+euYsMTsaIyuMmmk6d1V
Uw33sM/Jm2g2J5ebXBQUHVBeZMYFkF055iWiSyfxjL3TzeN+2XoncVncKQMx2rkm
pJVFD0NGFZcboqE7NAf78XhgIJp1Srd4v2f0H4W/q69tsSlre2v7eD46wCRcSfFj
HB1ZYTRpUAQ2oimY98QEkbp6tOtR0Zi28pa0w6EIUfWyYAR+F13dyTeIqIrfhJJk
mYunQUVzR9yAiby8UzFzakahCm3T7Kxwr2eYTR8I5pGInI41/BDkQek7K2ge8i6T
GwMl8Kujyy6GADLbRyKUaGS9yQNNLxaUGvppvO+xI1E77TFz1VHMRaF096pOKEcI
hFiF/071S0CL01VHVHeAvsXE3Jn1ue0wFSs/AVoE4nr6iLxQB0oFU2aWYYkfAYdz
bjbl81EUINk45hx65BhRQsAsovo48565nH2u9SUbcpBJQ4rUQKsjFw+lMXLe4vQN
8XWaMDMVtSOo+Cn4+HbWcv+Mwyl56JYworuE1SNyuQuIhRRkZKds7RRaqyVyw+x1
cOFJ1if5tEnpG9jPBpJbGvI9VsqnUyzWKRGuY3zf3REqIq5pbZH8O8fKY/KjLzdg
F+NDw6qUENWH+Pkdtg2qeYOlSE0U5xR128yMKc4kUi7KFcfj2u5pLeL5KoJtF4xC
R8sWlr6CIVG8zYo+88e0A9f1xrl3iJuQMOvctl5HopG8To/XsUM4y5Vf5NxemGpm
Tc7GbEQSwNeYGptBGMeITGNYpsSIiVSjEMM03Gvtxu5cewyDr2q3QbNPxorM2X1k
3MKlSQ+gNoqKTjtmIfYYvkBFlGJcxjfudzb3UBdJUrTd5WG3PH4UQXVes4lY7ayP
8lta9bFeiYtIjqm6hVTdCLTft801MwcWfvgplOuK/s3PyPZhSbCHM69SKbOUhseb
pfgf/IxiJRt50Fxxr5IL+EMYOEbJmUuXzeSmwmF9SXy+HrFmt7QIiM+iBFGuoecz
SVK/GVIlYngcIG3a7vuxBoXoYKmnKSc+gwNBSjoyMPppzl7KXq/gRezs6k7NvgBL
hx5q4EF2s6h3KZz0OT+5pHFRJ6aoxKOh4FQrus7BUduBDzXTFbOBQZjrDCVllO6T
HQ6DvK0Y2a7YyTUvNLTBa3FO3H0of51zEzaWFbx6C2zBoXQ/Uk7szb9RuxSKjkdO
z5b/3bS6uIjnozQV/hkKp/ayAR/GI/HZK5tmnoLBwpm1GoNAJNf/97vYomrMRinh
+jLlzshAcrZ2wgbq4f982j2jozuXxLYCks8WjKoSE7HlkRWyi3QdxVVGCrHlvDM1
mo5cX8tbmPnlC7kxWZjQuIZTByuVIcUUtiFTVD6dvbgkgWQYXCMqjzUrPZ9juClZ
8xRAV88INMF6U9sgSwhkk76Ugb0nQTU660n5MBxvTpGfKTr0/e5xWPyBTRuTR4n7
ZvB8PYIaXdYCAkxjj20DoxgSfabzGSJlt4uBKBsJt+QdLnc3kIC64uENHWd1A9gS
D4LjE710GEyEN7WEGMVB7E6anHrN5qh8VpE0lskQacssZs3p+CAK+sV6Eqqf1cUi
V1U0xYzcPR4fs3qybEsgLx15jsODwCkXv8KpVc7Jr2Zq+ue6B2AaHVGxK8wVo4v4
ZUKVEvt8F0eGaQJh7gBXDoTT4WDh7Fq9yFtqSUxNX+s8huIsc44vK8HHhHXFGZko
mQeRF5Aj+Zj3NLIjvVUuo6kZTbQgNcJc3p/NFiP38PYb+duPqQoYx+kF13kedrO+
HZYrfXU96CYSpm9lvSxYo1K1FnmOUArMZfwIkYycdaY7Q1IjEDKgCvW8xiAzyHot
hm6u3iSPI7p8fVY9+j+Yr3oxqWBGsrHiwY8BdH23B1HPQaexN0FoxnyWJi72QRQV
TiGYHRFmshQE6f4lh+2vLCrMhXZGZ5N1/lndps04xC6iPCiXbP9EsK1mE73dzwdb
rEdlKk2/zR7onQJ2NsRHLA7LHMtYITvOeh0hBkXqr9XJUMOhou9VMqI30ikECVt2
+Ck6hxWehaIvF3iiNnqCegHYQVpsEWcP7B0Hikyv4WilBHaYT4SVPlqKfmX0Il/G
5/PjZq5vB176VaZkBKvunDfRuev1lg2jlqiHxTYDxMdK2VIQGaxNby7EIBkPoJL8
j8hKZu1ADpl/loYwejJTX3C3Pb6wQS9a9mfXYsAsvPEgVOU9sxxwZoZ6yMXQ5TWT
ESez32TLqZUOxY+dJ2nHJ1qbrs+z4dCzJvBKV1yHrUZBsw6Ef0apu2x2+V4eCdcz
t0Af4uuZpOzVrc6L10p9RruKel/0G2g6P8V4hVaT+8Mmm4H3lhuARXkR/osIox7G
zRQXBsYDVHkE4eHP580lJ69DVvfC8gqsdiYb0eGLiOoqFhErazZNGHlU+D2gluc0
6VittzWu26pfoSbATZt/6s18DnTjGCIFL7wNv269oqPYDNYHs4HMFzKQcAJ5IBc8
2lVGmJoP5KcoFQP74wMKBxnbpHOSbnTKxXfsqEviuBS4ET7hzrP78uhyl6t2XUQG
bhxlMLsT3oW8p2gc0d2wDWyw2KUASj1XV+wQiJiAgTnIb2DGPM3PVY3pR4aYZP8L
hfK8fC7zVAqTZ5OXzNLRNRENO8OFxIjomQNR9VP2u0+bkjYnKMkw6iMuVAjHWlet
oEK8I598wNhnYnoDMx1gX8+WIRksdPitlzq8KUSXpQ4sN8drLwkiPHZqw+XA0gfS
jqrmDXXA8HbEcefuvW52P27MNAO03Npfepbd4cqXaNybZOX5dT8SzxLf1O/AORSN
mRFhqtNpktf/JR3fl+4o7clX6q0QhM5HrdPOfg0tSe4ER0RPQWt8eciZm9zLvt4r
XB+dB5PHNQ232t0ikkuIRHwaXv39smMqp8PiFclx/JfH8jCgKVH4qRD9dpuSSHGn
41jbOOKbZpt+a4VC5TYkEYw9YcFOlo5uFJdKuSJOG1ZW84ERFOlygGJuwFq3X++h
MOrApArH9eVD7RDs6B5XJOKFaODgMD3mVNJEuKM2glwtTYqn79cPQADIjbp1ZwRA
JNe+U7r5wVgz6ABtTA2SkAtmG+ZiNy7poeb2f9OYQ2xnD7qeaQIZDZE4+6cJ19TN
AtepULlUKY97iDDuJrzkfD/ZqcYsh+sx5ekBW5HUFvHzXiimqIDGze18lLSU+tcd
HWumz4m90chZzCPk5xm9I1sGAsJ2avdV8ChGrskt+uwBxQ2LDTQDp204P+by4X/O
KTtw/KNyw0+2rEwTzvxqDD5J1dENmquSXlTDpCY4E+zs3eIwybgEL+G/nAoNQ9j4
Ba9mMZDZgalrz8zCXHV8kIWcRUejLGUFx7kOp5rfRxX5MSigV6VmKY1rN7iGV5AC
fAjFOsxqMhNhqN5Oy0q2rPPMy2Vh/vGEUuitLl+lIp3zoxsh+i8eSMFzY4bz3BAH
oE3nUDwfCzg8shUpU+6FF+6HFtb/t6RdWIw5d4Xph5ux4rP8cDznWbzYExe33Zue
wi6gdhnhKmxc+VncKYpDcFzrjHIyYA3gj85o3GSmUp9FaE0qkK5mgmNNb46qLhdp
vi72iETvRGLfIJ2143KmJDz4dtabJmLCBjPj0OSlESIeUxHHL4rtEbq2p0cV6FEr
pUe4DYr14cCvFEjqu1HsTGagRebZ4HSkbk5UmO8Jnz2w5TF9cpr4Eph0Z//Gqnap
mtzNHu/dN4OGAB1nEwKcY0mnGnJjOP0fGsMEvzl7Wc0ue+4gO+y8I6dXqcWwGgNL
Vsovoq84YeteyOgM8sHkM1eQ77rDxsoHgIeWD+dT+yas7QE/NE5U9cxsMY4pA+3x
a20Ab8UTR47/+zP9fRXNqXSeeUXp3qBM4TAmex/yNNvDPM5DhjNfkkGZcWmjwn3m
Ma7eQs2fnJeFSD6xWbF293J6i5fM+hQGGiVaWij0V3XxKFj0TiS+pa+DJ7FCrNBJ
wr8VFLbNNS2qJk/6tcce6ft1bqEPZWvP+Z+NqFy+nhpZFegx0CQxg5Pp3wNJ4yXD
fdxohq9v6DeAuKRLD7zi/La96T6iWlyiVwo5goDkBMCdFIhyPrmrWmOL6w9beOvI
kEebLjpN93wOFceJ9dxw9aagZL/pse6uQE4jSlbR/EB2G78kazSN/K3KSI8DnNZ3
6vuWHHjt+U0b4UB3uxDPCWqe5Hwa3Bet2TyXxrzQFfQrRwhwWLHcIJvJI25av2W6
LsjJTWBUI5SevhrdWgZ8Yd4S8JbxOiB/cw8oEcFsJmhk7AcxBnqkhN6yN0rj/zGi
8yv730hcYwG3psTdn2YZEnDDQJgSko4WBvqMnQ2ixD6FPAH65kau0uP1Be0TrBpe
IOElpJhv06L0fvYMiIDg+GIOeHs3eVIZF30q3fCve/NDrcIY+9IBFeGex2UvPMZ2
WLXd84BPTn/ERyRDG3CtOaLV8pHNb3yDQuZImzi0/KcDr90QnsfS8NypEaREDYzu
LH2nNOgRvsbeHAEOawT7QOYRcAVPRiR5cuNGfBpPMPXpnfBlbrn/OwKYWJCZLXLG
1Pg5kFJbkHvGJFgBt7WAzO3MRQCUTJWBMI3elVHNvk4H6kh6DU/A4wXBv70LX80k
mwOp6BTJtKR73QKrfWQdvehRLyam5FNZTMvrLlNFdNNGuuNjr6PdOprGYrF4mb85
bixvBzpMf8G0WG/ZmoHUHky0eVKcaPAyOz1hFGRKyDnviVMTENPaS6hI4oaialgr
w+AqlQGYfdbQrqXXVvoAejRTpjlrOBxVqAmxRy9uI/PILbFdRnpUSbA0UnYa0oNY
fOsp0ZzBxejig36Tq4xHabUd76Dq3Bt3EgtryTBFLnO1+S6JDVGRIcZ9aL9uMCoG
T/wfdSOi1von5GjWEAUJLIPmIxM1o+iQVKHKLhjcJShzWEt1YYqNfZ9Zb5iqex31
JZnsBvs2F2RMWez9DPde5jmHUiPkPPnqDTBfrYXnpVVUK1A+cZ1Bu1j4j/DWmDYE
I9IeSzkmIiOvUihI0jEjfHKCK4EHzq/Ic+pGvdeA4v/POtf2Txbflqt7LfD07hcT
+ECsJNcZ4L+EnL5e3xAf/AozelfLcgxKcSJYjHkW7cLzByzml6HBIKtfPdjd7Tl+
FNMQBJ3/p82M5DIHwlzMefeiPG5Nrg+hBJXAD9kH0+2QcqU8u0+zl9NOwJRFWjIe
HS9QTT6XWFqtNtiIzx3VT/sUyrXPAjOVsVU77qtj7Volav0bY0Xva1yQeygz2PQO
Rs+o7h8y/Fl6EdPDc61tcuOC/BTiEZQfeW6RV8+9pSAvK3JONcZ6Sjr8KjXjeyFI
Q19vrbTqOXto6nDOT9UKmz28noaUTjcy7VymFOggKhNhmxkDkVvyjqTXDfJCEWaS
XeZhgH4CynTwWpB1qok7ZoOvcYLM6NuisVyHR9NTOftS889mFQK5SC+I+W0V4MiA
/BJha0QpHWwGFwckHNiPVIbaKggbMwn+Bg8Jc5OyDYKAU/DcCC52ESyW3iCDRXLa
2OMJnjmgqlL3XhWkIWkZr5iPslTiyKTAOn3D0UYb+3t6J4cQE4LnZD3xI/rIXVVy
nz45PSe6JgVbWxMSHJi1XRyay1EoCyLVNPzKaG3PYSoFgBgTLkdaHxbdw5yFnaWY
i50WaTbQuz2QZQRR6H5LB+pQfBD0BUI7goU9/7Y79+e2ZMmia3kE9nbX0CBv35mr
v0pJtW9AeH/0LwvqlSVF6JldzqMAMduZ1Tv+QBqWJBrlY7RPyjGfEBsXTrla7+Wj
zWZbt3LP60YMlivX/WOUS0rWNBErVYm0qRqHlXh46Azj/mY0gBc6Sgtu7wu6vEB9
xfdwUHTQ2+waT9VV/HxEWLkffqrSsFopRegmFe7jJr6/nrfrUeeH0lIkd763WipI
DYwLxaacvlMC8mFiuDhoKuZZZEIKHGg9helSyBfTuwAV11u4UyfDlv8ODseXH6e9
NeAkoE2J1voNk1z+F7wg2okHp4VgE97dIplLVW79u2jNP2Xp3nqjCUaBRh0gZpEf
NA8qMGv0JvakK96ampo3on0hMk0nQ0zkHJ8+CyZ6jZkBBiSJY7hqOVMuOTA1GK7t
+nC+3pyEJtbTGLQ7Jh7k9yawReeTKOJ8NBfirHElsWQDD+mva/3Whf8xcijF6T28
wzKEcW7ynQM45NEjq7vbiMv9IWiY04/kKEPX/JOPqBQDrgEkhZvaw9RIvPHysBdh
GnTx5Qi7dkor7du9iBzoFf2+CUD7XZByMPZ3cNHJAyYPGC0o54Pp5/bZoXaMSqrT
IUewMbySsODucjCqqEK/05PqGIwR2capb76lFnCCBAUdIhfExW/6zlQlEay6V9It
/a/ctFZUqqCTrTzcEA1sRUqIbjnIzNN8tfiMRtqR5u4sUXAXlTlLreiuoVru36Km
sIywM2JL2z3XDjtIpFLQJOOnmV86HS2Vl3e9WxBHj1lufzmA9XcIR8hnxwW3SXis
JtIkJGZ5jp2qUcdGuhB+SL1zonCCxbhainZbpWv5BBXJwkCGmnBFhx+105w7mvpw
BsUyz3HFp9fG9C6pwQz+M+RigNMvMK2hmvabBvedm8wZexuV1oo44ewTmtuxpQVR
ICPScZBldpeJUnN07I3iNwoQs1MRp+aQ3r8/svBPVJG088UtHRZDSBNYGTbt1IZx
zuyfnQXJhowAOWb6WBZ8y1TNDljqdPy/RK1uz7GH+sQ25q4BWMBeuQGqKs53yFrV
Wl289kSI5JMksuD73RtE1H8xTSja0cJcHgckQn5a8KS8LhZDmfw1pACmD52ObmP4
hHEnY+TMUXlqRUgho3/WhP7OHrNLRnTdA1knwkCDn4VoqvypQttD3EiZyXfM1uDs
nJaLZTwJlJjGJVqEefuawZSJqFSeX+EHHXH3pna0gO21V8IkFTMkLJPktLjO7QhR
allL0YVVo70PbEDmwCqa90oKYdxPqSqkFESELvzWgDdq4v03DpqGNhlc95HdQfTG
qnd/hJHBpWeK2pi7+d/Jnl2Kc2ym4q7RRngfOX5HQbEmv8HF8E/KipUukglWabk6
113OAbEEqk43Q27kT0P+URl4XK3moOcnlq3NoZLA/3B65s/MYoA8Bkt4nADlvIyB
b3dyBaRSvMPKshY2BVLQ8kKDAzkvMLzjS+N+N3BJRFG8GyKvh+CzE1fraqCgb19m
qG/B9RvKLI7DXvFST19CZGOFrGOtik/gPP3UqCITQHWKbLPctBuU6FNzuMI3jW5G
o5fQIgvcejASy+vTTygXDfafkswIUkv0clRFsAFybiqiuNvP9IA+sJkL0A3L7eQG
PfPCsln7ELLvwGTq/WlyUxcM86/JT2nLk+OrNSYysD1r02NTpFiWSw+oe386IQYi
bsIQdlk8AtCg4ukjjjioz1czgt/sUVykGQj+gXJ0d4+voH/rfnxwfgRkCDbQiF0J
pJgVk3Wy+FDbx7jQ53khZjJYERy9WZOAnhysu9eJna4WQ/F0NOg80D1S3dHgCKxY
4YfCjr+GKsnuR5ha/XNJyxBaL9tACR61u0X66izjjin5xeXdyN2RP6KY3Mv5SxbD
/zRuvfordTc/+Rld+76u+oHtMoY2n2/NWXGDqkQCM0yrACv5LH2U5MwrPgRmtN9n
Cngql9rEdA6tVdpRCMScUZ1bd1wGYRyaekEAGC7DzunPjAFaxgqncVFm1sd6XuLX
AsIWaK/SRwR8nzAY8a9xQChLM7ZxLyx1tCE4/roQCsE4dg0M2gxiHM/9FxyssNiS
pTeJRXcqTDScieFoXBOamkUPprcUDgV4cYDwIrmb8Tf+JZV5ZosWxjzLLKwmSJRr
cYZhhEffbQyTo5umflwcJj168kusmaKj98qedazZm6VcVntckun7hPf4qVNHtmnX
6FNuFSl6SpvMTAdjC49nNiFZVyXFk5otmITkw8K5+oEczqWTYt+ZJz+HKs4GgaGy
QmXAC3d4dtjcOH7a3flW7t+gklhMCOcUSEnGvQrGMJfHWwL3TgrCl54cPuQigjqX
n3meP8+qYxyHXMTBzmKxdnvkK/fPxp4It41qyNNgM/sittkO1t5OX6jPl66FZpG5
nQoUJSfL8xAfvXRdJIF+Q1NnFlDwSmUpNmJL0CQo6wFJp9QKzeWmNpzClV4eXCIM
LGHtjUy0eKbZx6SKRGbOqqDULQtQKkeBKbMMS+AJw8wRpkuBhcVAU4XoRoQk7wEF
8uG1XpR6FITErmKGEox6qCPEWGZ4dzsGUpbiAMEw6HJQ57Tmt3SeYQQN9n+cLfbF
qNW9v1D+yCwcfiwdska2/9Hghs0wjbYpuMBIYGvm/P4plTHCG8qMLRolc09kusN5
UTh0/2/OGGSEDebGXe7ozVukVzZsJ7pShZwjdIImD/RDSE+hbagi6DMV/itln+oY
PtO9xdvnEW88GYESV3QCC/vH3P3MfqBKdX2O8yVwWxcMdTPijUJ4owb0cXh9KS6i
TXM2MOAcFugzfHyDlKwZ5KSlec1oTw5Emz+rP9OVif3ei7ymNWfhedHqC/btTGzb
sWXvumMCf4dsN8UUZ6AWxCwWrRZmiHF0ZFE8geK2FefQMuBvC/pgnbU7FZTA8VRT
jtenBi8thHU620y0wrF8NnaPhA6LzJ2c6tiG9bv8A47v8Y+sANoe37yvpRx+ZOb+
a+uZJiqFeq50l3i312gNcF+GNcJMJTjGfGJevDa8ompGZZzrbe4LQ4nBsnRUz9rh
uGhOjGw9IHrN/vnlk014v10ouJ/5TdVgl9k/x4rxpnjM6vUm2wBrezqRuQOuYAiB
SkQIXuflhZ6W9jg1wicOsGapOCqnR0ui1BAeDLIVgTZ59yba9L+l9D5mZTv/3JLg
G0dPmEiniTuB7cJrCegmh7EioeY2mC3BrCBlDuJTvSBklLm7xRbnqRuW67FPi+f2
9AVbLX0y+kiXxOZbWxRScQkvHcbHi1x61qdZwDQrm59nwdwHvzFNZLHKG9asdZnm
r1SXt0iAHaLKW/kOqbPdsJM8mKdZJtOx/5Gws6EiIb3vZY5cVgoE9EpLT2JRdHrL
/fFtnmzms9lpdbnxrPWjU98Oj/4a+sIwwFEbkHwo6o0dUEDU85AQMeLBXFGLvMca
bn3AFIEnC4RALXyZO11Tr6UjkSXLCr5txXyqB8vhB3xthtmgA97IBzF7WSM3kjnS
PaAOCn7zguVa25gsHYuIwmfedh6/oxvyrMXAVceLhvumgk7kPk/WoN88zLALGchg
K4yO3f6coSBnRVtqYRcmEyT+DNza0zLOZzdjPNKehye/qjUrTnSt6AzSM7knnlaC
klEbrcLTMpDhoZ5eaVwIUkv4xOxgr26OQetmTyx9St6DdR3mtDyDRu8UUS5ES4nY
Jny7AK0dLsilXRwL2LtTL+YKURiV9o+oy0zwpDdW7LYa8c/a458sfn1fL4fyJ17n
uLo+NLDFvZv4U4iwHY7YH6z4LmN+1e6z8uKpkajHedx/bbQrkOwg95WNGWS0Fp+B
CKV4bNYSVZm+ttEGLEzsTfVLlww7Qv08fGpDgSC1m7Xcx5gIQKsoeyO/ySWd0+rd
7maxoNyROfRgzkwQJU/GHRZ8yrOY3Yxt/tqj8uMWVGkPgoUnlOhOmgVxvunJphxZ
RUo8ksOdfVgehuygbVZmXoHvTdkORWVtfviVw0dOllh2y/EhHG6/jO/DAj4DNevY
x1sOXAvhi61hnGEQZ9CdlptshDJTRDOVUpoJIlmZ+l6gYQQpY+Fu+qHmYcG9QgOf
fyb+3LhCIuR6uGiPgUP8s1CxvmfNm/Fcb8Dn9C9jpUvm36u3/YA+wS1PtXLtPGQ7
EOH8kEsjLKLNxS9S+XASnX8qwm42vQLqCCRUsA2fhXAEvU1+1TCHVNMk6p5kKsBt
LvNrKjh2FUdua7D7VS39pC1nSlnWlCAsBXciNx1eA/9KvWFnHZB0fjF06TXYRjKo
VhaxNhgRkRBfelp+Wep3bf6b0JoodGa1rjgTbItALEl9pKgZcoEukQzNxsLHID0G
GVuwDlk9WRZUhpvhoH6ZTeJX2LnDEMhWWLFeMh2KgGOCS+kAJw0JRehOWxZ+gVHn
EfL8kNr+gLlHxm3avt+gAepQmm4tVqXWPvaACUeRooq0osoGZHwBlErdsiK7yooU
Len9qI4nvTSAm5VwkTQL7ABqv90RK4nWG5XSHI1kD9+1h+9OMF2dU25d6sW1ezr6
hm6FzPu5jZTpTtrJmQXxmxLcd6R2y3MZguvjA3a4DnTt315sYSopisP+G0eHmahl
w9O5wDQwf6QQ/8tTbIUUR8gAm7uRQ+MrkGUVXDFbVyBbP1hoKpudRcqU8AVbbbA6
kNcx/8rJUxLqVlwWJUzP6463jLdKPUCBoLZ4vJ+57j1/A680cfQOrKM5nxhEAEOp
cZ3vmu6n4TcdIpbJa5u/EvOhj9lImyp2WjTVGP8trA4eTxoOeIAqHknzTzQp7Yyb
cHXaQJe8AWkrhjWb1j/WaHh2Nan83d85o8qtiy6Onl0X9bAy3E6/vATKclsYIad6
tfLUQldfbCTUA0hYvrFns7sDzMwVYsPZIvkvRFOlKs1cj64CDnQl3h0WB4eYZZI4
xZaGZPgM8sCBmmuEVsZucwmJcvsZWL7IO3QMjhXHw9V2yzeYU3fLNdf/jI3uNoS5
vaBSoFWeRUFk17d80ir9jKjORSj8TuhBAGQawCbtvpd+jgKa/OD3ROyUkRCxGXGM
s32zOFBGGAv1xdnd6hNlOVYDxAHE/R/NYKPqkT+5+ZQEmoeI1M7E4eEPZE9JKH2G
9m2xSb4sQtHplwitf8JcDPwIKfWcUMH1uPvTInyf/WxVPXsKbIsteYQK/deaPyY0
y/ACxK8L3a+kz4CNIlMaiNBNliyODMictIjClsaw1Y1QTSjDu5wiSPGEnjKwAFYf
9zJVlBMCGQRmy03ZqjPbgqcu08FL7vEkxrE35r/WfBD+ywbjd0jF5xd8qQcDtApf
Yq+P0D5Me+Kr4hqLJkM95CZg8Vk1YGEHm6PxLJxpAhAkW+dKT+23Y3MvjVigcfAf
/l/kvOQVMyDnw94G6IwRvENEIxycS/tHHisPrfL9lO0PQ5qUDqbRkSFEjTwYPwNw
NzNQoXDgrmPcbrGqfroyF85yUjREpmUc+qT9kOeW5Pp7zqRIrncxGHHQMG8Ba3Pu
XCbT2YsINZRUdoaPFGHm0d9w5g3u5BW76oG/ITnGkt4szMWsLTYaEVBNJzX1bTM4
uXcUjj7UIgl+ItEEBN6TFIoXh0/s3ByQKQvHq9su012JG+CnbJ+J0rRIvLc/u84Y
oRp1wn7H70KevDEMt4ILVj4Q0UqriLhc7sl1XEIRxCfb8dkbZb6LmZiOb0fZ7ipf
PqxKy3CA91RKxeTSS+6ev5ZRrQSjwg01WoTeLs0k/JQYojDXzkER3BRMJZ7xrGy0
/p77cY+KVZBeDdD4gzi3QP5bQaPWlCbJpBR1fK8vS6lTizvtkxwJ7Io4uFWztr1a
YMOuFYUT1EU14bD7RtK0T6B/x3hJk90gxp2dPW2uW/pn02sRrMQ1kGQJTxQsw1DD
f+6TkVNnSwLxb/aX54bBHy93RB9FrpRDM4PcFnQLchCldK4jjdTCoJ/V+KVvC65i
5gi8fz3xfFTr63c3aM7jtnULEKRkkVCpPWavID5LjCtS8Vsr/idrxvKSqzwqK1on
vhi9HagOlRWESY4vx4mS9Q5Vr3LxCibBuz4JfbIRcbUUk7R1q8oF8voAXmn17Iif
JgUau80k40QFCPHX+guYrhXsP1tsqsTAES0ZAFNbWWkg9gPFRzTAi5DiR/R9jeXj
9lJaKQf8JgYApmNbWAkb6osZYiAcG4rCAzeGuXjMtpRiAAaORu+jN3wQcWmqkcYI
PvfUN7REfH8s8vna4KKeXimZdJqOmIqJVC68IH5LQsJadW86nHboTw5qUS8bAD3+
qf6c2UHa3iSdCysh3c5lQapXDsI5r35RpvOn9qSuxFcY5I/k/bdo7mG/xGC1CD8m
DyeQzFrwJ8nX9r9jEH37Ey0JRmeRg/hHSQuk6ZWkUF40C85DoYyIRKZ8ZJZwtjyx
4HY8zv08mO+wRJyJq+R2vHn/gRdgSZpR3xQI5xqVjnWS++M62lxUlMPyQYWHnyyk
z81NrQ+4czLJFOlnZm2l+Osba1fekYOv6jaDt2hVQL4F2ER9KwCtgphJEvQEomFT
6pjpG/QJQby6ef6FJLcngKSnra6l4c893BPoJtweGo6jC6oTwU+bz9j4fQZ9ScIY
Oncjoi9cOp9zirZAEvxb/hOP9YbCv1AoPD6yLDboCgM08gji0Ut3DY/mgkVDTgJT
cxOdiBbQM45qUAG/kg6KJ1iybilHBoNI2HZdAvcJXB5Iyu1sA3S0zC4jdueSeRxC
z+Aos8OggR9y8RmLkpJoYZTrASOt2GWH7RITts75ts/NGi3FJV6Z9mTfuDrOl7Cr
+/OA59pLL3yPzB+33QzWfnn0CDHi8hyo8VIGy7zmp8yBfpXfmIlcoVvU2w0DCrb5
dMPCr6XHIkhR2TuMsjKa8+0ZbSOvEd+sqgl2KxrBrkNLmAFc5nbIJVZ2pIUPLXtk
EYGkKO7O7L0JYI+UdOlCfLv/pqGpG77ecQVhfJWX/B0oc5o6Q31reil15895T8gY
HR51a9zreJrtP6WGICzekqkXy8c2dV9whkGhdZJ4RhUHg4qj7e6cUk46NFpj/vhI
i1WUaemedP93JyysTnNKKjO7dajLj5ofeTIA2pKfEnl3L0Ms9LmTQFmQMpFC5vtp
02M0g/n3L+ED8aNtiCejleaVz7aa2X3rwlVCggVtvctP3ALLHCAAmMk/NeiRBebe
OLl4k+gzDaCyevpVoUrD40j2XTGASEg7+q0sxxRrKi9/8uHqimHBbADwxtdWMWo5
C90ZcpH314mk4N4Y0YJGhUGG5OufkWEDon5y2txWryRJNVciSJK/ARnFb4ySVIR9
2bELitilIIJHmizcQdGD4FkuTzD3dG6wWvPtpKQbiYQNhF3+m6pZ1Qr7aZ0XMC24
ee1cUCWb7F01fvc7DkNvE2HF16BmoJ/mzsvDFocMp5g+jsOqwWjpF9hZH2uwMSgv
bJfZE95iCrQMuedoj4KqkkjEwdHGjZnk86S0U1KxrGFmxGtQOEdem1OOnyW2xc7K
9qw+9z32u0KeAvKnCDYhG+3ATIXgu88LXR6xTEMBWX/a5Sg1WuOdZVTBoG+Mmwsg
AkXRDSEYZxDRbZ9w6rkw12mGC+b43Li4GwYLNcxUd5FLISJ44BoPMiHofPAMecqe
kNwELplbRSatPFjSYi9Zfg90SFU9KUfMn/tjxpG6NXy5bXwQhiBSwM+y45FRFsB0
04ISW6BbOIy/1NCIdjhNjoEx7muctTg/4qjIlcIexZjI7OFNkhitoAi56bWPb+f9
cS80bNbHXjcBBYg210ANXobGlRHIHZXunFkqb1ss1KK+xr8ru9Gl+U9JKr8Crseq
1vuT0nDFCzuIrg/IHs96zg5ek/vuVn1sAdzORG5Q9DosLAp3SEz5+XGrq0MlM5qX
/JMikEoqDSANT33kOEpUShUFjHLmXM/hSTmLdbRBcIvfPqGr9LXYgxgDujvKEHWh
56SXRbkG7TwN95fIFdsddcuDxZBEBVR/U2rbFO+Hv7Lo79bLPrZoy3VfXAUA1/TR
eZ6k4LQoLH3qZCBt89LpCJM4oNiK9ssAKv124lwNdrUoDRNfZGSfsF9Eg3gqTKfl
/uJP5PDO44m+VRb58h2DHOM5LKEeA0tof0o8C8Cyq/W9iYqPcH7TX0TaKZfma7yl
zYmQpXMweiXpxZNSUSK0+daRoHKHMNf6y+gvNnrzWrFngPCScFyYKeuqlUkubLqv
QXUzwXN+MGtbFmPzcPa1GWGT2FJFpAC2HQRBbqRzxNxOizjHLJa9HGYLt9Ib5HkL
YLYLzQdTO4VfTDn7lcg+ED30puHnt5rA2Ox6DcEvNo/OYzXXABAbQIA4c+66uEnk
hOfS5WK/2Xpzc2DujH/oX6Zuzh4K9BEppiSWG9NNxCujnj9VufXZrTyBluGjH/kg
Oq9lvD7N8kD4HpidwrcvgPQP/mxMLDsyVnuEPgOtxXauOVb5dYDUMskXO0kmQmi2
Y1wV1qrSpXjzGdhjbXzUOQFNEpFU08kPJgFxF1kPQQdX8865pRZ5VM90rhzForWN
0+h7wLoKjIGX3eBpq525I09XvnBkbUjntdIQbFu4qdx6Z/h/N6cBMc1CeNxAqfl8
pg45qEFLgaf0tJe4KQ9U3fsF5jdSwJR+gWhkas+7cUmkgt02oY+kUOs6kqxw1I0n
nK1fhPTqqU+Ny/PqM1Q3tCblc4J7PeGD74jULAst2qxZYJxvCd4qbIS15eXYYdEr
3FkbTIFYnqoxpaE3aMtSmCwVkDjrt4FW/4oW9U6tDBX9fU5f0CVsoUdhgYXeaDoD
MCsh7cWGAplg/bWjtTkk9RjGmGNumsPu/QwSH1l5J21zmZCSL7MhQ+4OxttpuF5/
w47t1a/cc+b0Qh2i5aRtxLB61qn2af9jC75KSQg1XtJPOb2VVgZ4DT2CSjybyAxq
L8uXNkobU7ujPmljmZFnHAY4KbIj/0hUxNxnXPThouwMYtm9oENZn+hw+XzsPeJq
29fz/3iV0dorfexIj3II4VWJp3x8uO2XbtONG1YD9g2ITI6hohW9gwu3umvxsZqg
WEWr/rU1T/lY7q1IVItI63vCLbM07M78MSBvSWjW9/+nHlxGb0oslf2Q5rI0bDPv
YyzFa5bKr1W+7XdYrr+eAl8Le4Lm58Hrr23s1TE5JSq/UMpz+L3qE6O/nWemzYdg
3Lc8KPBazhSO7kEbB+Up2YlWwhm+TQcpM2LHswp9TnO+O4bQ8kfvSB28I7N44Hm+
463Xxwlx8VWqAfNBbXmDtEg6vj4rWuA7D1F9kaBqYPU+S0bDq0lptT6r/JuUTx4j
5bN8UsIY6abXDZLMwapktxTr5UbIafqOJNTVGRs8vqzBfyOs7Kquy3ywTAjAbDku
voM62Kj4i7kqzRGHcNe4uqGQlx+tt8CTzis7uK6EtOumKaXwh5ofmVfIIJYerihX
QcY0KXLGDar3K8kXHsaKCziqQD2hoZbKUWji6XbK0D91jY8CBnTvWLDXtB76bY1C
n8ZFFIePDG/MewVMdiV1Xz+bu7alfIJq3sX3fWTxidgkIMtYH8ElVVQ02XHK+pv8
7Y+1x0na1viwwecexxbCRropxo67PItzm0v7e+J4OsFl6bTK0CvSl2p4e99acqhc
6pdCuSzK23fqFVvFTbsRei2WR/w/twSO4wDz2xQHxppw/4ZouUWOdnrAD860hT9c
Lonvp+V3iGoYLQ9dWA2ZJW1oLwdZtBkCBTWZ4gcHO//HKmwtLjMtcJg/Fr+uJpjg
a2amwp10gdZ6bgHVs2k+D1eQ4i6hS+/UTIbofqro6jZZ4bLJCvmhK0MlUZJqTk1/
oju2vtqTOEMWZbQDz5W6jmA6K1PfL7mwekAdXHnv8WnLKENDK+zJfVWhURQmrKbp
0XuMDisXTmNtf1WqD0mB+FjJGiPc3ig8QJg6f7ShvIusrOvZYADFyRHeKmJTgZwa
dMPx399ZIBtGr3JKJygVMyEV4rGznvM9OurNknXEGApiqO688ZR3MZe5dSJXPV/8
MxsrQejcVkFjDy3tHSsrA69jYJYD5QptKR3JEQQURjMi5ovvbpw3hr4sGYt14i9F
++Ul6Pf3tJPIQ41Mj9TIWMcuVN8I9VJb0/0Rdf0kFKcgFyZv6q+alSuEzQLnBxCE
rH8ZGgYlLPw5Lac91MdWLT4uSmF/MRVyFDgwlK/9XR5dzk1CUSgkM2iG7d85jCdZ
s5Rq7U+CbF+RjK6mW0l/o2Saa07klr2B2r1sFIwNBbGuPFRu6Oq3lqfEiB6UBXUA
DLQUDxIzOunUPrIe9xPIiqsaI8GR64tTk6vh+IWv2+vVztuMCZ8Jiv56vmr/k1FU
bnbTwNhGLbGq27T49LRu2zM1j28Sienf7sTkB7GO+UMF89gzrVOe/Aj/FHQro0qo
5+MfQ5t7W2OLwZh3mWDIXxDPJg3zgXu4PrdVhaMIHTjA6lUvpLqwrtjGac/+4yLF
BtneP4RlG4BXIcHrj3CbECvV9H7If+iSUlSj1OTs2GBp20ddKOUfwwf7uK8/kGNm
J4Jl0IfNpqSuSH7AbjDOyKXXYXVdcZi0F/7nV/Ue+5k+/Fe39YG98CGOBOTUdhyl
BB5347O1vnS094N8FcACG33fH2bmrTGX9LMDpxo0Ux+NrwSWfuPMLiMyw3+JmrYG
rHwBWbQIpC5Fyo+0juHOPfaJnmKA3EWXMWTRsRGqi7P5t9O/8jQO0SX5Vxw2fXSi
+pRKti/KAM7slsPME7+BSnkJ/nlV4+XPAgvBhk9Yp2DYP793Y3dELVSYuFMgUikL
HcYa1pLj5PQVgeeC6c2yJ1u4xpj0MpB1UukqW8Udi5tRPpUuNMPVY4U65wYaxBNc
G+GDWItaryjha/+qj4PuT6qPnvk7N2PENQVS6KydC9rFd2wD0kvo4SKMN57sVcqJ
cGy75uBze1V4DGwHUcod9aTc9l4j6PlUt9DwRrXz+LbS7nW5EFzibvkN9/ulYct6
BOS+rqNg1Gj8JccGTz+6bTkAHPD9vRrx642Ro0pQm4AMh0uMKKzKna/+Zdp2ZEv7
3Z6WjM6/xLf8uyD1dtdG2BVNU+lzl8ty6hB8KZ1hk85Wiib9gqkTrlFrXZ0SPN4O
FK8DwKnTkle9q9r4NEUViqkBk7hoJGwvf6N42mekb1PAccszuC6aTNQfSKpaZKFU
8YX8NnH1AX5a7vPL3wVlksl3SI42cdQ/OCj3zEWZAmJj5gIDNRwvaajSUiRgxKuz
DFRwP+5FPeAwAkoq5MpjvAw8eK/21y3gT/Y93zY/b8EOxhjBUcasZyw6IG9SbH0W
EaJDWEnfM+tixJcNkIlcyLMte+fMkg2dM95sCj4o3iwiWYPtbcbhTGhItCinYN4l
0n0290L4jM9zsbzn/MNlV/fcIFHR4/YUOR/RHaEqQiPdGN7N/EThQPSiJ6Nm//KE
AoLr8p1brdx7RrISyMuJmEoI+XFXwTduwFHCFqnMKpiol9oiyr99WOnG+xSfq5Lf
BUu8FOFQt8NHn3daf7Ru9+ND4AEV7pjlUhTX8zszLztJY25TzxqVo0mB7fdkgfMi
H+jaZrxGQvvToBNZZrhp8IAv0ZGbOEc5FJ1AzzhGpKc92xqsFsNbqZuDw7dg7HGX
wj5TrzThN4S+9V8cuV8VqmghL8V7mR6JtTcGjd8thTMw5gPy9AbF3bzD09PTBJ8e
MkEM8j0sAlGyGGaaXknoehH/O28nCYv82xZoq3WtsRfEqMxuPxu/GSM+buNNFKPd
MTubWuzpwXNN5CNqIU558tNmnwx33vJQ1TRlQAYHqiQi5xbOFvEXkko2Yny6/+LK
b0QU99o6qyhg6IMgdpvDTA4/nTmZTgcYPRdsgTIbrKC2PrUnwgpT1SddSQ49H1UD
qxdMcCPP7q5HAPeJHgNwO5I6hRsVnaSde+6k3RKuWvWQci/dKYDBHYXAfQqp64iH
YXSjN6mN6hmApF6RMyESgqi8q8qcx4It6hdotJtwViB3pv1wp64/pUSKkTT07xzY
x44D1nuuMurVG4VlNNxg+ofGaDlySkgKQ5BwhmU4MO+B9dELD+hjFQDY/yR+rUcb
SflnPyUkcRQI80cfuEvDOviBnRHDSAerY9gOP8Kh8C1Nq550iCQIlJe7aJVFVtZw
YXdYq9GWEqlz6wgmjzmDcfMvQQHILHLv7k1GfH1hAXR4Eu4LvxXd1fJ8KgVpA0y0
sGXnKu2PqU0hGj707VlJ82/KlB0+laNxjXqcAcV9CxVvMW2GID21nKmY78Z5ijtx
hlsS1pocPJ81Ms/maXXjjPwdSusDOwNjPsYNGR5bkSmUPjhHlpDEQYWyV6tQHrq1
AByIsYcV8QrQLDHgbRJda2uI4Yv79aG5Pku43c9HNwK1bjYCNEsjnYQQGIUZ8IXD
Tkuu7DdlE242uYhUfIiqyNFpo+k0UGQqN98f/XvaPT3Ha3gcOuLypNVdBjcDXjHE
E8kd3o32ETywSml4C87i8Wm23jIv2zuXRink63qpoPXAxTHhuKC7rXWx9MAI3NsE
QGF7Y3pFKvkODD+++QYHoDYS+kEt+WVDg97GDjs4dBIYaVXlF78H/CW/o1X+Mv/5
cG1T3ZaKAep2Cdy39u2Nih+wELeVW5fPPzkAjuWq6s2WR2IYM0p6WfrShx0SMN4+
JGInC+/vGm2/I5NlmeCO3Gens8oKjoVO8cSMKtdKNPkqof3aQ/so9fPGLyzDBUUF
so9CfU1ibewh61IIapXnIYPDH3okugLsiRB5xdsJ8V7PiLBNFkt1MGVEeg0xGDsI
4GU4sSj6Vr0wkLOdAj6s32lWWGup9L6s8KeEI/AO5Az56DVgUbI08OGd/q3QqbAH
wFZ1LNVKlpFLNcwqKaxFKSbhD/JUDEcmQIbGexHdgN20nqaS9iMuyn/JO4AuVy3F
xH9nIkFiPc1sISkm7LiLhaOzFK4jxAEZDkc1B18Ru+Nk+Y8b718g55tUy8rNO6sc
sKktlcVXgOaWDIFeg76xm5YI+R61sj+zPf6I1FYPo1zxC8w8hmb/+4G+YmStngN9
i+caH2w1kPSgGzbb3+HlpfV3zROS5H7IC3fT4L8m9601AKR/9OquxaJkms3hNToE
tpYLPYTQcPBwzmipG6BI+sS4mr72tFgBCsl0t7lJgxuLQSC/XvwQ52HVVLbLxCId
1a71byXpc0shbYnJXiStjXXrc48muk42OlzwrnFwN2o88TVDzBlI6TYZYGYOtHFK
BeyDcR17BHICgsjsfFe6OZy2aCNz8uOsyA52X3hfpmBWtb6BbzFpUHAumG92Igwa
NHk0eMxuVOcQ82aO8qrPW2/EpPRguh/fRBttIeWZmYmvHwqHSF+cTOXzhF0T6QZ/
SmdXUD4RTIoPDBk7/bcUKt8K2ug0odrT4a7WFBJz+L/8cxJYX3cO6Cp0Xz5GtvtH
R6PTi7gY+yudoKRweq0awlctooklXwzitFk2xxmpopo3sYnUkpG6GnqAwCY9dLMb
Bpk+xq+K9UHuvOpZqVkm2UUkOwMcslpD1a1vtvuliH6BjsLQnu9sv+0K8jfy/H8i
hsbEDL5jXov6Z4nk/ByrqGNVOueRJBhbyJaMIMMVias5rRwZRE4XtfDAmw6i4bZp
wporq2zuUDNCpXl3KVEy6xoimi8+Cw40OhAzzCafFvXBsJ1p6r2HMY911Muw7rxo
OTzIcb29E3nVvfcuPqqJXwd2Q29CD+Cz5MxY6RUSDd8EliU19rHDocAm9LF3TiFe
Aqb6ekt2ZmzvSLsaLRhqXGeuNInO9HlLlun0y/S62ziYV2lDcDEQGM1JwbuAthWj
lFx7ZqzAHVmHwNeyXpgXUNEdeADolvsIoOMHXLoiar67UMZprkdeDoFQvDruaMRg
DigunrX+35a9mCoQqAGGn/jBOhedNAez+p8cm9R7/4xZHVE3aUQcdY68x98sgORy
vTgIDXyx6OC9N6+DGCY6XlW3V5xccEqd/bjnRm6gINZWuH5HtAqUj9jgxjRLsv4e
UGrqSym3doiExffR0EgU1NmF8S4EPskkO7XmIwaoT0UZnC26eSiHY07QnVXaIYZk
Ni0SoxkfT1YPhDUbsozqC6it7lxYwW1wPOJR+wFHVmoIzeVyxur4v8MmEh/duayR
eSzYyflzU/9OcE2xn4YahkG+DEEOhxhPKjZ9ZDOgQ8quyvGC9R1+5CHt4RMKppG9
dQ7CWd2KJlN25X+3vPTPfshZJNbHkWShXUaE5P9WYbrFAoJFxth29ZWZ0pT0jsPw
lMxDhe4r25TkpAIfTGDG46hGyeNi5d9DQWHZjmkZQWEBA0lFUmUXWXDMre1udNJT
Ry/egvGCIOBohAUlob+8NgZr7GH/HqjuJexdn6gvEcsGzzIhpEYz+YuiLm5uQyph
RSPPuZKSXeV9bgarOL2PE0UeMRUmJY8R/+73xZLqDCa2NrDCSxtuIuhJJ0ZNkHCL
a86npBXN0SApihuuc0j9Eo0zQKHSxPSaLCCcMiUt0PaqrUyQog47RO63z3xJefK8
uSPIgxnqwj/2gSi8xE8d5lul7aEJikrXnYi5gLP7I5Zna/DhNzRI5LYYFcvuyqal
mRa5s+B1fQ86xUobmYpD8tybgJplje28+3grU23kD9NQJLDYUnMAChcHR5pKzYj5
VekDvxKeHFUzMKTTjMtwJoPZ1rmzlOF6nGcZ8JVLFaMnFG4gViw6pnBibHjfa0+q
XYbCzqKIiU2DWt7ckPwp3oTwTb3xmoW4pTiNPqEzqTtGW+M8wAsryZnYvolM5WZV
R8gxW8A+0+P/nXjEyF33WPYC58LKi5ncanrmCrotsn9mGqxPIv1vvYoQVV9jl+Od
MUv7tr6JNJ88SBfnhTr89CY3RXdYH9BNRxid404CK2Hb3p2K4cQWPWEthYXQDIJo
95D+maTB6qtTu9ytfER/+lRO8N+CBg4xuUsRr57mJcjnI0ps1y8iM73eYJUIEMwn
BtcS8o9FDuJIY4N95klQZy2dC01Gt8vtI+mOCEprQOF1wUzBmy/w4224J+KFJ5fu
2Q0lwO6NEuYBC7B47PPT3pNZQ7q6nWVGnjoTNvOQjIUDh3r7GYqK5d6VKljhlIrX
AoMd00LXYIiGLhQjW/hQrFR2eeR4OC/MyMe1/smXKvyrKVLBVZTjYYoXfhJ+N8xk
OS30E8CQfV+mrcr3kJ9qpX3ddlUoLlW+5gxXx9gsP+CRqG/SJIKjrqc3mVP1DtYd
l0/wZzNLgGhOvVzN+TXWNJ3zLevj+01lNBPQDMjV9nuPJnft8Tkx96pvl34cM038
I3FdhyXl3hZDTzWdD0wkLSSwQ/gtp4eLn+gwsZsvo9thArsrKZLtaNa06iyu8I8C
Wgw92EpIOA5sI5Kdo78/cejo2ed3OFUkIf0dB/wuM2U3uQePCmdw4WM9sCt09Nwd
8SPN0dm1My8vDQEamTYI+5Ky9YOtZ3tAYXJ+imUP9mjj9j1ahEECb6DmQnUM7jWG
XIRxLna9Y9eZkkz6YOpfR6O8L6VLeZHntIn2fnPy/f5xIK23id0z71waGKGkXsdq
gQYzxMei2xHLVZbjQMMkc+ZS5UBHVVSfeYLF2ySmhn5DKDOwDj/Pm41N35bkSuYR
CidcuWmKVtNsyn/gUKKYezC6BAwtDzcAOKpKh8x3fRvUv53YeeiP/9/2I4CVlL+w
s4LEfXdbo27K+UlyfOYC1kAuRWCodJgGC/GrC6Lih7QAVMpibwXXeL1weT2tUVKZ
Ok234OA6sQAjx1otq7vpKgSAXJdeyAFgdvYzoBOO+fzXF6XkR5Pe1i9DC285NdVB
5foGnzfmrgQ0LbphS8BCJ0LnVJ2We5JCKdfAvGGPqB+dIcwEAhSwDZ9t/rcI+FF/
gKACoVyF/l95GdIzKlDa9M+JqpPdxCqrWYv97OW6+FKPzRxbqsxicPD0jXY6FZEk
rlI9TVcj2n9E4X3nftd28iNUuRbgatajxp4eNlV4mlnVWAMPl1NZOU7RiwPbYBCq
l97nXY7otkV3vDQQgMtfeKpH2RWLH9dCaCmU4QvN5ozhGmFwEEVQlDmB4O2ahVJ8
L/zMmqON61yqA+yBhoa/rrVu4imF8PGFDDkqKJS5r9iq5yHDfciilgSTmEUMWgkg
SDPZAz+Nj9klg8ibu7L8fwyTlVyBK65nkVPI07itUhQDM2qiuzZRXSabdP2J97BR
LoI7IZ22AQLz7pwHo6FweVociJpXbau05rBj1YVE8FvXp1HDyUvXbmIlT90VqbEW
7kYQ1mIeqmnDvjRx7+ILbeL5l0ZMzyakNyM0qDfYkpxft6tPf4iFCvbOejkk8R8M
pIDiRGe6ii0QZQ1BoZdGRr9PtS9BHNRoCYurRwpJokRVRgr+UErl84xDER0dCZpY
8qHX4ICLdgPJ2iZSdXF9MDawG4sTQ+DAzJwp51WFX+4V0wbF0QeBABBl1HxF31MH
8sc7ETPXG6a+LaLGByS3MSbgv/YTNapBCyA1AyKhiyBMZXWewWdvNKQNDNLU8j7K
54p+y1rcx2m8IDCv4k1fpMm9sJYjAfDJ7xVTyGCVqtMLUu3debfPM0b/ifJFQHtD
fZxkDVlTcQ/NYPYJgoG5cbUVHZWlWvFgvwqYzQTnTl5VtBdu+aFfVYanJKdk8gHM
jF/gIUVDKUvweslCOvuYKsZgIJoLiKBY7Xo4I8yxe4+seLxhyHf86S5pKsDnPMsZ
arqRWbFq2zSRJMta5zsCshmUhqQCUM1Tx3b+ntWIvojhcMcIEo7keIlQvlsixP89
KoWyKQWXVhF26OzVdW0Z3W1p8HHFaT+l3kD731cdm0O5OQsbLvkQteVKG3K7zTvf
RRcpTwLmlgBhmnLqJRbf0K/bEHJeAVxF9c7A19FGf2HLiekPtZDwshfFNeRzMXP4
MtRSkwj/c+gSK8v0zseScPmwRAJ5asnW0rRoHV6dssNp3daiW9fXOL9KHFCvStDa
I4VnRwJrPJeLPm7lpzTAWAHA5YGCgaGkYlQRfyD8+skdoVPdaNfEF2ky65CuTKsd
KwRsuNMNOY09mAM/r3g7Y9fkwbcKN5b+5R6HE7uP4cTlt9cVt1ZlZvhztriKqXgB
NVPsncDHHHA3Orjt3rBeL0e9tuaV2EWQrs4SRMKnEUeoWY+pF+pK1jg08UDEsIXr
HxoGQ+4Z8DHJxUIM5I2ZOJlRA0oLL47UMAZMApFUCSzH7bEGfIUvSnYxeAcmmQqc
7sDdW2zz/w6SLcCs2dau/ZGKiGY7ZxE0Rmu5S/nAMixVDfA+0R/eNHckDRTY8uqT
iUA7hu9jfsgc+FtPNw/ehND/0GEQ1vTPE7JHEwPTYCxuWkg1wtoe0DyveoBd8/JI
X8wDX3MHa9u1sMqySEqyq+2+NUtlW4tmsAoUR+iAAwHY6mRgrTckFBRfOsLd9+0U
wECXSAjEzrqBpsbcAe/cORrJnEn2Aktvzh77W4+zm60+uWJZlvyWh9Tx5Lgdc14w
AKzvXF+T0jWtNE2M4n0V2F6gA8fwJ0JpNPRshEE1CpEOSCnkvTFg555pbxhif3zu
NLK1evek0wpT1Yrorw0ejWvmEBmM8h4ntWJWGaccbGy1guyxL/4gPhB2jWEKSY4l
2PIizRqMJ2dvxarWYviPoq8El0VHmqjKTAkai0SG5v1fU2ITqsr7BnDkKX+Zbe3K
KDSo7h09FY3pVDC5gW6Wu4gtnqjnOpuyo6NzO+DplJaaz3VEHW9O/IPKVHoVulI5
Mz9oe9/ri51fVS332Z8v1FGivYuOf2SrYyPLRxgMjrjArkNav6lYVKkwJfCmvS7R
COTJi7o2A/cE1GrQXadE7Ri9uLNdUKFt5F2jL4IAaw/Tsf9J9eWhsO8VNeodOD1D
J9lv8L3ZhrGq3KBLRqCmtby4i+TOQLjij6F33wwUCaDAbPMBF9RpIyzSwFj/N2mr
eXALytVyy/99SWmQKsZAn5IPzt6uEyOL+IcCYABJOLKlzED2TXFtpNfnoUA20odH
S2uXyA5gSmO6G8YmxsIbg9fetPJsmr4rVtuVqSJIirkoozt1oztvxVJctHRpzXdG
jTgobAiIrGeskiUIkkKIpgwHZEGttZ2kceKFdDbcYCbIa6mUM9qQEQFoa7u24qVM
OnellqHU2f2hlkujxsqnWgragiYOSAvreRbo7b/3NUbQZkteHlOWAbkPFrnbcB/o
a+07JphF23VSmguchgPbeni5OOdhnJY6y5taKpsaALEcpwZe1Lrc7Y5zI59zud7r
btdOhJb5tbfpqzwTZYhVKgUG6cy247C2kwS7bB/aEDEsT6X+MpXSW5oYoq/51d2V
c6gRcMze+WGMIaS1+AUtEZCOhgmG1v7m5gIdXzTWQKnBRv7d6itbPHA346BXkbRF
IMBb0veoVWu9lnCC2GjpcSW41BUssLRqIqXww+pZRuKZjOeBT8a++Kjwy28shJUt
e+ugbQZ6B5GmtVmoQR/dDHcnyYMaw3dOIx7Bxu9qzyQ66IpEs0eRHv9s+x1TXzU4
eq8mdoo6yFMatka1hubznwhagYVJfiX7m9DRKrYCRytF+3F8d0NRubzZFYc8u/fg
3XqwL53xUzg7NTHRXw+sDz5xWQZArVJNBrDXsTK6yx9jCNc9romrTZo79BBJ5n2c
LvPcNkXyfnQ63kXcx7jcfuM7Le1+Hl1udZO49TG2x2EVSPT6jsnOnk4ZwLyx/IuT
Cq1AbOCvqcgvxBVg1KQ06vI2bb1vqs9J500/2WdnR06fPRyba4bXPU7dMlBPw0hp
vffPu+a/RE3kMNGWM7wA3XEp5TdV2QwTJEJBtQkiBAru7zUrjJr0Ayx78r4Q+mCn
nanGrxNj1prh1Q17g7pxSmx9Ci9kyc82W0ggX9P+RLvVA1un1gq6xxJi3fKz7sna
WHUPoXHlVpA33rVyQsLxrY6FnW6gCL5kPZT8hct5P3PbCR8Qb8cc3ZJ91I7Gtz4H
Y9MGy6W54ysBetZEjA+Y7Pu6PgXeDh2Sb+cfY4Ao4ANZ6PA9uB67sTY45ZLxnd4V
2IffOIG2HqodPHFKtKXi9MLpfSOf8dzi6O7NRLzZXVa4e+X6upKCaW3mqbkYGpLY
sPfKnsjeZPIC8ybsY4jvVeQ1vqH4sdUyHDIjVYYl+nkJbpIbnDOB/GuuQMa02wzB
8t8yHGNouIX3ZpGelzMoipLyB+T/MVw/NxNpuk9AO6VKhBuQVlvY8m3M9JA0Enh6
/eEtngv2gJt21XuFp7QimcSFA0UGWGcj/861v9n53eiuPkaIYDF2v6zSws9Qa5l9
iwtmWyptclj6broHtNdTW0CF4+4zD7Cb9a3/CHitEbgrzOmjqmZZDymk2Vx8czX0
pOCQQESKm3ITFCUurqhzThrti6DTAIFXT/2Y6+N3DRQGRiRxYtWF9gh6UlLr5T7w
+sdbe1/GIuwdXXLcmEUnln7qM4XAMlOyY36DT7sFayFNOReV2dLhHGDTpbceDEyn
XajJyj+wD//swSpZOC3c93/OumxDszF1f3POlpwNd6EXzCcQIYcRweK9LZBOxTuB
yxxNFAJp59SxeHHbfnuflOk5h4N2LWBOvk8w/U/cjkLsWQ7ia0hQ6FFY0laySbWR
mVB/nWw7FfrLdOJ+t5qXlNoiv7utAp2PMrHH2Wp6wwvq9ORDX5M4YfqmSHdI9YmE
Q4p9jWJzaY7jXcbaHqATIcS83AScCDjjndbQGYcvStpgtnytbYAjEq+Um+97N/YT
5TtfXnQeV6hJ4EGseOq5JUtqaYYHc7O7nOx1Acai+Co8giPPXHhtFaAUS4KfTeeT
SIcv9VH3gaboKzOQpK0hr8TO7HniIMhR4av5w7igw1qMOTuHskIfGoWnyeP4F8ZD
y2vOxZmGMunY1slMVzEbE71wkbnntD0bfnUDLAf5O9uInXl/UcmiE7Yv+rP6X4jN
cBeVTW12LxSNj7iml4EOQmGBUgJgeQ3klaT6tk9VVgomaxrpKVJNi/wCSh4Mhr/4
8WaOD7LZSzv2oXWQVO1nTR7BP/jIGuMFGKfL2oGpe34gzZfgF9HPl3LFD0q8+n/W
sO852kSAd3Qfz5VEDhOXMEU8hxSX+T5AsQflDH6r7Wb4ZtJg9OXgcP57MpoRa0NB
gr/8pZK6cCzYTMkW1Ngcm6pl9lkPc62cFY3+o3A1QH8atqAWUVpKusZ1eANQsuY4
Bp9nnt0LMooq7NMuarz7KJWQnfFzYEAMTTRbkiQPM+iNtnyl9lW9Vq4DCkNGrdpx
4ppy88ArXlvOjFiv0fctI+0pp3M0pXDn5IxZHviUjSvQ4Tkc4UGGIzAITd9oHsbz
bBYWWL8KblEOIHH0+rKc9eNKlQuzs4B/EpC5otgKzx2HfxlK3dDjkmw+5cCMJGIG
mo9BS6N9D8koecyTKK5yvMmzUDZ0C/3HSct/FosUdxzJIAXN+X57yJqnh+c9Y2ZQ
QlVv3gR/9rU6KjKjHCDXacdVEGOJECu/1GPCwBrQONPH5GnibsJf5QgRidaQo6Fy
0z4e55KTBtdlGoX16Be0vIVIEBD+W608r6szSPLYh72VCFRAr3EWuab+w1PI7SH5
9E/YgFPs3BC5KTCgw1mteuKuj3GA2PKkjS3Jn74N/h+vXiXjDZ2WttAiGVp2/9h9
g1GbHh6e6zXNqGrwKxF1o+SJFfpjZ7yhQESMgrZp6+2faAvNNmGKgMXKp0Hlab03
PNa0aWL1b1nCCCCBLiqtYxkTtfBkySRtZzkVqL1mUPy6s481uo7a6lTtbRB/0DJU
nF5Jt85LPSbOB2Qha5WPFuAn+CdU7U2mZfyqWahJTWIwAenLJrlTyjAuAqT8VljB
nWAQmCCoyA/7+1rs/UW8Ss85kNK57nBTnhrFUCBE+1yg5ihTMrQye4mYckB1F7ke
kQKUxrQusshXV4+tCQp+z6yEbb5i3P/ClkhP23pqvdLHhyY4AeVd2uHPoUFqvcp6
ubnUxnc3loyOykJbYvYIAzTJ4T7ZFjuH+AekzWLg2hXrp3Zfc+Zh73jw9zPWMuPo
pvfaZZeLNoV8hinsi+hkwiNgCq4QLYnqh0msBbd3/FHuiUEnFZzfTdP2vOWOgBjA
gOfEz5eP/7v637FHVSJAOIYNe17Pe6S/hmmGBi4f6kBt8369PidWeaGSoTK/MUZJ
5YHvVBuhxqZL/Yc5SRxADiLSIb+8JaQ4PW0pKf6SKpoigjWEjmmxM9f44uLkctjF
Qs+G80AkNCP2k2Ws4TGVUG4D9HyDTiV+NV6pG7GXk7o4GBKRtQRO3BLadMG6s2aq
adz6dXD0R0UfRpGFDFhIGa8MudG/UXHDQYOL2RJJ22B1A78ni/n2DT8HXwevepOu
U1FE3pUuBe8/5jb2UMuasashCrI4oqWSEA9fOHTaqK35P7z4iRlHLsVkVqSo4YnN
+cjBgqmkYZRe1O/P/DeaBKKDcQzHTWs2WAfJkF0Zx8KNQn5NUyBXdIRCf7NOEdap
OrZqCbyQeiEDlmupbTlg6v6T8ZYXQIPaloAqaVgmtZSBWyrmtRC2SApQoEysO2V1
zOYrQSx7XtZpwoj3OO55Mnd3OL4rVcorbgnNsYzKdPcAvcGWb8whtcCJ9eDQuTqE
Us5H57hxRHDt3wfuJsFhB7Mk5w4oudZrL36ovYGVPWLe21uTWL6rpofxfNsWQEsQ
0Fj39/i9QdUcpY1MUgDHA4mrvfwYviHMQ9RkoVu2UAxkmwHokVYoVx0uLuP31uOF
vHkBA8w5beKMGjMEXTS7YYsr2Mm1RUhQBfFvHmNpR1T+jC2D5FfVy276oT9Uy00T
aXH+459cFQdsfzvo4ZiSkIRNBLLPhNexAyPoFkhiYYKthPuDM2xW7lbA+s/xGGf0
FyKMAVEpOII9z9kvgbND+sCpVLMEKkuwpMQCJMCFB8GJghkBPn9YTeIxOLNEfgnB
RXmM55MRXzUmYK1s40CIhJgEBBWgv6ArB2cgTpFluREsq7uQ4yA+LXi1yoCaDfsZ
rH5z0LEt3FSqgtwckCNkbIT5Nm9wvh9nh9R4FPBEXdYHH9etUvdwondS+VrMGPNS
C5PldN70+9rOAhmLxch+7a4p639VtNO1aldtQN2MHun9QEsOUlTWwpTge0h1keQF
S+tVHsUYQghaWdi7MBvUCNqYU1gB8oFNIVUyQHkOc4FATTFK4680UGQQWdxuOULa
G/3QmUmRM0C2KdNNJ+KUpqmZFNWqRzSr3MsnxHqP3vOryYVbXeC0ZT/dbvtWCsIt
43sxPc7Ws1lL/BWxqIigDVQSIXdtSzkA5rJ7Uz77dPQA8OndOB6vFQO4UuvWAnsg
h09O1HPXxxTsOo0tFDBZ2/9lJm8g5UMj73f+QNkLjQHgO6ta1lkHJeA48PFS3GqK
trIRz3Uf6oOHEGbOD+YbB95oMot5w3lxVYZcszBBHXh+/r41cr6HkamheGiI4i/J
p7nTYLsG5zpT1L+rZGRct4dL6sqXssOVWHZ3CkHxxnjezCIrZKFDIx6jjxFzjWrD
W2UMdmLxmnjZEZRdz1uvdouZJRA9TIhsvgHhtfmuRBRMP5fEKetE/YkVxj8Fco7s
l8sPBRUkLDPmjrchBotOqjPnxGolydIR5z1aGYbl+G0jNC8gYJjiYd/u+LJWV+Ry
DUydexwK5ogfac2sRPPJTlLEKg12Tmjaqc3nOLnQYhzO7R/CQusg0zGBzzjp6vFC
vxICg/mHmGt+0vn8O3bD5U6HMUYmsbf3G9qXCzG5DMR1EqPGbyESRvv35UkArUSa
YaYtv5vWYouJ7QBG/wLrH5iOfLdRe/iXBl507UOMQjEztnjMprDImHne2HQO5DBE
arOD1orbDeA4osNygcubcIP3WvGywkRaNRFYIB9g9EI6uN0ABDaK10SKulTyHsjd
HFENgFdnkRuphDCZaLUGiJeYaeTUk80N1YLlLHTFx7clJJ5RmRYVyal24wPT/8/M
9JRW7UMx8bZq0ieMOzBhet9lssdoobdVcOKKH2Llm482LznCc9DoTOWIjQva+jqu
jaYFZnqyaDAxgiXBlTsnxiK7FTpuwyJvg634rkS+byXXoXLC0SHwUgdoJ4sDB5IE
BKEnONKM849Pf6X1fKAxhtv+ui/HBfAW3DcolQVjMcYaR39cS5z7UZuvQCsEDj0A
xHws0rB0AOHBCelH0k8k+mGHx5KLsVROe9f/483wGC0ghEhBbLozEbV/T1yNc/Ot
Dd+WNfFoSspY4M/EcGj9dtM+Bs1JZO2evWUeVyUiAK2E0V+5lbXPdkis/G3ChUJK
2c4hkYQJIqsvo6WPlu4kR6EvJBK9009HKOmd/2H1eLUbFiQoh5GTXQ8v21uVZhHM
EPuGOPRs2i3p2M1aKA7kdRu13WYTvFYbZdEgv8Up8ExWvol6sKu8/7SmuLGfVEkf
iXJJy3xvNzP57Wgiibnki4Hzx82DVSwGk1xQ02uYQ7b3wJY6KU6IdwoyibT0DYhH
9KO930rI/qgJqAF4nC51yYKSJn4IvdtLBBh9uYlbr8DlhOnxgJjb+O6KFKdDk4MY
PUyusy4bJ58aAasS5Jtf0KN4DkdvNz0oHObNex90icdIIfxfxQnD09/F5dKz/2Qq
iK4vhaa074cgG2Vqp14TRb5B48Jd+umGQqaEzSFBS/FyYwiez86XleyA6a4EzoN3
/DEr5v/6Bx9J5brbfUr0FMyAVsYzbfmcAAXXt7OLwd8A28s2rsIECzBGZkmBuCut
RJqwssVQxyiaxAXnB37Of73f0PbIb4YHH9p2XWiK95fOPNkITDf+VP8ZpFisPo90
2jLrx3ignQs2GjoY+Vtj6p1527whsk6yj1BtvZzsS8/6CvOBAjnfWHufw6n2X5iZ
JAEMREKA1QuA+XPe1DLflA6IhuDea185/e1qm/mVRHqYi5egTfIkRDYYIejOfpzj
NgcpU5SThPX94/kIjBPt7wqs0UqKfALONoXYZlWqMgn3XRmLu8y0khO6JhFZAVBY
RnSyakFZoSuh4RlRExmlie843ZxP6F6TuAtIHWQzGzsR/2HKo1G2DD+4IkmFy7Vi
EO5ypuORV70divVjWpF0wBx2DZpVIGpSUlpsLzMTgW0WYlvabbvgLrqECOcAN7LR
zEeDek1wd0UzsBWODPrYAneN0aXCCzGxi6lRwV1xNyN9TSMdbr9f2SH3KJZzQTeA
ul1i8xxxPXQ3pjfvdkxN5mLZksjQQVLeYMJUOjVYliWxxVoe4YYLSItJXMAusR0/
aZar9qTLLfWQo73dbiy1SF55fAZWVhx9bPI/GghgUrqLvnGeKG8XzAHY24bfT3tX
nnkE5cG7pYcFEf5JcApikez9US0kNy8VemRP9mv1ioWnURDbugXdtbTtVHyfX/R8
GsTySj4i8pFH0CoKC8tc7GJ4qNqTlTwSjQZDyh9VZoOcStihAqy37Ldxhau+Mwsd
t7y9z/B16i5btGT5a6pECON1n0HKRLnthJJzgE0Q46U+0Sq59/LCJXPiyTvRYPnw
OZjKjBIzHkZL0DMOD/Erkq+EjgHYv6XJIfHDM1rbChW9ocwU+vopSn3tkYnxmvYQ
NANFhbR/VIeuO4MVHBLFFai3+1FeoxKEW/tbNynRLBzaHxhw8zDat29bcHsFR9ot
7CGWmVKMIAJU5SvczUdbngp/cmI1R3VchF24bkm5p3VOyoxmIZfI3Aocwu5YyoTr
r+iFc1YW9JfqFW0KIWonaameKzL0j5Ggcgya4loz699qj5jsO2WkCr1d8OEeXPSx
XsSZ5bmxF87g5hn0FeAGABFkWxGIolRRh1gLnFmlJx9kaS7jFRTNQ0Ao+UrM0Ue8
k7vl/aA/PoV0plF5XBH9zMsQcRRpMsqFM+cszAtiEvdLFDDvQYh3SDXNCwgSCAAc
cQ+V4MFt7ARDm3jGdOtjI/VPksnH8DdzZDVB7uEKwCtW3+NU86gAjjyNesf+tBe+
Qn+XatGNhGlIOnnnD3tJTaivGC1UgcnRq9aTtPp23ci0r6pc8Qry/HBeT70QODc0
bY0oXQczv8yXKRQRzFYveBPX1FJajCzVp5ZAnq2r3NqnghG0+tX7pG8G7RFAuS/0
Xl01MMeFtPFfmtrl5OHqlW3xgqKmoLQKFDvjnXLw8tMAz4eGbNNTsfEHg9gLLjET
VDo8T4cxa9GsPCaGW7Nk7uz5DD/OSRTFjOMZRnzA6ui11O8sS7ZQyyzwWW3KXVlT
g4NdisCbfYcpZkyf+RnrWmZ3Uwgam3Yj05C35Ew4i53+WLCSY3VBMQuhpxxkWV0g
aMpNwsnWGiv41bmDOSfTWOvFkVwbVut/3XFI0eq9pBCHnqu4KbEpaV8HVNHnCPVH
fi16h7bI6ulPxLocP8jiLtW5cEnZLn458H1rUp3yhBKu9qYnWWL3tTMWk/GrlKyh
B9S94UCdDVhl+5wS1yCtM5iOFvfJgA9CeX/0wyENC8/x5J+BgAgrEqnLqRw48lp9
SeCAdb911zkRtkg94Z5BA6+dEwn2f+j00jgFTzqSWzOgVGqyCN2z9i+SyRCHAVRs
vATJUgiEhVoqzj9NKEM7WerW3Ea1VCGEeJtQvA/GXy4YKye7f9j4Nvmfuz4uy0dq
PzGXcSQ2OeTCRLako3COV77JHj0vsrpc4broPDEcq+6JSi65Agbxx5suR4Y8o4+3
PC+SpR1vM5/bF+2unS6vpmyQ61bsC37aE8sirEK+YDlj0s4W5X70FmMsqgSEjeFv
x5ypUCAFFb4PjGvVwpcviSwmWAaoyzfDyenvRn9/IdqazuGJpGlmPksqk6zOJxCp
jkvDQz7dPBWvVIZ0gLN+J+HIrFticHJAygpYMT+2GFtxuJvihi4Ddxwc2lr6UXFb
BWAqIgwnlIEOYXHVtAnIIRd/xqxSNTa1oWuPm4eN76J9SkL7Qa3IGT7p2Rq6imgB
svegBL1z6CYO72+wnrX/FwXEtdVzf8JHzmRxUujAZ/1xInBv4mTlykT4QuLh2+Km
AvQjHxvbELhLcjoq5WSWEg31Lao6dJYbHAajd4MnYzGo8HNYeNtXXVsTtKS38Kw7
843YwomNiSnUKzZkLdLQlS3whzjg1GTTefloWS+dYWX2sdmQvxV5Z0Lcjff/OZ8G
9qGVS2JxItP/Ne36d10rNiwGM0h2lLMrWGLt0Oy3IttPF2wPO0C9Pq/v7e8I6RGj
bGXJHtjb3cSZK7lSKBPyPT8cDOUtGvZ8KLDeLjYsRkHilFwoSPLfUH6E5lWLVx62
up3TcRqpUUGLaP6NtSo2zDJHWlIKX63Lgta25vv+TASFzpcgAlDTEzUTONpdA+3+
7CBc05wzbWLx00zyLNBXOQldT0C8Tjij7dJnrb0tAcvIsfhDTkAYiccH7EKE5qD7
ni8R9+ZIkEqi2cdV0PGE8yzRAK4VxjEos1SwYd1HehRea6ydrxuLz7EtqGlvX4+A
ypIz5gkpYBvUiAy790G6dnX4R/NRO0qUQKEBRPYmiLK1Y0Hz9iRo7PVRwsX/W9/o
EkJXc1lOdnC7kKTaYIO+trrUrJyMC1ypNSy+qDq13zJ7r6DfONfMNHp77eqAMBDX
sY7THK1NfONX9osxb34tkOSpHHsOfRsRSLSmV3nvbneM/xQU5CrcZCCM7xATOsYm
1Y4/PKe2ql+V2FZlINEhbDtLJzy/gv/0GVysbb9xBrrO7l7Nf5v5GIx3DPyBL1db
j+JUccj243E3n6XoIVoW6KYs3tAjdHmPhip5iE5Rdwod1fivYDhfmqW3IU7uP9pz
zPgSl3tYBbTFLyCkQJj2iBcchDA/NDsiuQV/jQOfMkzBnLs/KVwcMCGvmJbtlZFC
daPkrMORiG+ToyJ9AKWSZvbfGD0p0c42qI8taUcnamxIAjCdyoixSoauXgq84JPS
E0Im1eIpVvDFqZsb5K1ZRNO/qXmfD/knmXaW5UnNtwwOYveSaebtrmnACtFuVmBo
U89bKX3/kNZCGNut5/ulL45+i8LLU23a7fUh+Q/KbuHdv69wJQknT0/s3Pt74Hjx
hSkTEc42w2CtzUVoWVh7WtT54qpAdkZAymTexKd6+aX3J9t5A27j+7NZc071hmn/
5CZHy6F5GDepXtBetjQtDgrQNPjXuBGICkcuzE68xonEFMoxrmXJ0ZWfnzhaNWvK
4nzakVHSULXM3CkPo5BHcli6mPLExTiXmk6qEZo96W4Ixb+yI1zaxsqEJ7I0jEbn
W+GjCYnwAL9aBKEY011qtMSNlhfkqNiX7A0CaeRI1rnL4DhyhMR5PNpxOFPq/XvP
1SF1ujDKs61zvinT4An+CvPz0+vtkaQplBFNeMGw58vEfnRgj1nH4NWbuojdUABY
v0AOV8QNGMmK+PYP4zUmtf4FcDC7j7ee5sVQot8t9D0XuKSSgH4A0ge1r+J0JIeV
swv2pO64Mmv2SV6c3IbE9h59GpVcYRV2rFRaO7n+tOOtctRvbkHMlFQwWDQvPM6c
cJBdfhQpxU/4BWDQ55bjeXUhWM7vOvIIBpDpaOQvZ9FU8A90kJomM9dpesZyUPcx
vfGFChyY2jfJSYICX6DriRuuygHW0+IJHo/RnhKGAswPs6xQLIjBVjXax2wCXpnK
5xPAeOSCQDgclsdlp8mzo3CuWz/oJ72hZlFSMAQtzMCrs7ooFC2XjuWJKqUSOUvu
LsgiyjNbojwbYj9uDxKLNslVnZ2YR4i3/xfpcSI38wDUMrtK67ugC1/dTZ7BxY3u
Z2Fjk7BJUtexpAOd2XQQd7EIZLOu5IChiz46oeOqVpY3d8Z0p90bd9JOUWt+b5ia
h+MB7ZK3iS9IuZ/uU+33CFmwnHscSTfD0iMWlsobfDu2Mh46X9Y9v+A3Yrnp8gXS
2Gaiz8ALBhIt8otM9/RACz6gkWj0NZuXagsBnC/gmzXviwm6oZ11zA+A50QqoDe1
BFDcUaXkkfLbN0HPOsNv4F11mA/CLqxXQfh1LRhiHuaw3viaAGx/AuZ1O1+Zv2U8
Pu6NqvF8uMUHA5HkqnuC/C8IxyrCMu+Kphs707BGBzsCqG3WNNPc/xwChe6H0S55
OESzSGgzIFOzGjXO+7z9bzb8NniBCFdfIp8tFC/avQxFYEegpdSswXT7SQC9ztZN
+bWE8RLXGOOYVHBPwS9iF76qgkyrOaeQZAcokQbQNQL2PyEuD4rkRtheV0AMhAgx
BFS0AVOWVGd+cQlGPZejGGXtfPKdfgFiuI9pb/Nx6PhWI6O7IYeKuX+GHWvZSPzC
M0PASZQumCAm90GFqnJf5NxGNO5bkBGJ/EYUuSocAZCMSQTB+ih7Yx7oqyhNjqax
Rbhy8YfMsBi/F65WFGg9OON3KOT+4eYKAV4wFyrUVK/HaC1qbq8NqTN+nMeLBy+Q
eLUbwpHm+i2uzJ62XVIX6hHNPgkMFXW+UzzqOeqpXvRIG0a+Vs9IJRrGdYZuOAXM
i2CVeBd6WApqOf/mWNisex+IjYx/EaqWl0MgYJwQzrs6w10Z/Oycol6aiuFE3jqZ
ZqT0JJkZT9WWUr4HIpcTT11+SN+rizZK9sXeyYbNO6NNk5bhLKjRyi32Rd3/MmuV
BCw9H1ZXR21kfwHPDZmtGkHW+smdBGPra8w4idqOHkl85veOmawycGD64+YmFYCo
vK4fwLNt64xg0RfKMGXanFVob7VPCCIi6UY3/1qZjzV5CwblflPrx+VBua+mD6vs
S7A3qbncAx6rw5T+oTN+6g05lL/S6vEdNNl8cq5ab9lyqLhtDUveb5+CQ94f8Vng
jvlm7046JJaoQBuJ1KDhCJA98gVrqmbvdlcCmBDhS8iXmuO6Nu88AcsE+S/wHXWK
dtDRt9pbvdM9qAQetfLEp4ZLuJLZ3Eefg2a1wcgPPYhUfhUlkGEJCqw2HCJiORLq
CoCoGtV96R8PLnVFHLMW7fy4mVEX5FPWcS6QLbfdaENAhNN3gFKAkmgTDUop4jGx
U5ufLH1l+QbO1hKHZmfuCxLPJ0YZJY//ifsGnfgwS3bs5iQDS8oraDdn3/AesM8o
n8cTjrHCNdeAxRDT6+bdKSRAk2BclESwvTpFjPECx5FKix7iM8YJaIAwXGCY3Yez
7dCr+a+laVYMSaFGSiDHanNIFM5VVg12D8dVaQbC6UA+Imj+Xe9KxT608ZSFbmPZ
4taBxJoNdMLP5qE+CYwgImuM+MbxKbSguIchaorlnm9tdfIY8oIkvGl0Wr0RAzii
Pya88rnKCH1kjrIKpGeZIduuIjvdouGZKYLnu6sNP5n+U889Z3gPE1UaLU5ZiKg3
e7NvRX8s/krSEjJRUsaarJELBu/+FQJrhdsrd3IIeDoArco+wQPLeE3R12SAHBIe
5XFAeGfuzONYmWGJ1JmLDl6fNieP9h7Qp6LtN1mIRaviuWAbt2mRJH89LDOGdH3Z
ExRNrb2oEt2xCt/W6JWTzbcp5IBNoaWrNbKGhbFm5NtFfwaeE8+1I7zvwj4M9O9m
1x49IrPTpey86LJTZaYVSZoWoMGeU1lv26u0+smntWzJUAvdLZ6awDifKOUkiuOQ
kGFZA5b8ikMoR2K54r+1gkpNHZLEZK/EN2rcZ6RhNUqCtZEg+BBRoAg/cpTgnk4i
vONzBuTM9Y5nL3euuMtSHs7+vUSK3aakkbFwOjY04O2KyCF0qQV8EWxlB0n5kd6y
C9Lc8w2HlOwchmrgmiN2v77cV14rAUWjdnbsc/HzVnl2e7ufcIAgrytkGiU+ZzHr
JOAt4ngXdrVtiE/Dockzy5+NK70xEPpsKapNrGq/f6C5IK+J1gsgWYEi9x0Ol+rF
UsRHSHCvQ1GPCu//S6cewtssdOCn1bDHfOJ0Mm/6YefIZUsQgizqKDcyWm8NbXus
/1IuHIxarxdXyhY10uSJ5BuoSWp6xjxoWlampzF/5DYOZqQEDW4J/XtHQ+QE8C+i
9b1wUJrTcmkTpRdk7NEtJ9P7ppdqp68wvgJYKfMIwIiSoxSIKlAlkOcNQy5Sd2Jo
V/sn4IBXP805EBB5KminGUlnSiNNfmYVSvxf/Gn0OEro/JlXz0De7TM+diDTXt63
HEdGy9J9s3Gbm4Lplp3crx2wdAXflgqYe0zOatk1WwdZrhU4IVwq0YAa4bIfVBwo
FTpTI6IdslN/uoCt9wJRpNyVrqTS7NmmFCvs6ym4a1r21R7c7ZqAqoqgLlpEcxwn
3RCGTbChLEUfsfIejSxvJPcUHdhJcEIjsPIpvD0s1EnNEUTBoO0bOA91pvaZhuRS
JNGAHJ6KRnXz25isJdiBUw13XOqgKscerSf77OiyKbAvv9F77G0ZdUCFGGVvXfpZ
STG1gk3N7IZD7LMRscDOnOWy0lZckwQrg+itRx0cv2CqbR3jcFtljcyl3v1zEQCU
GziW442Dwv/ErvPxeQ4h6zvQMSZvanXz704LulJ5p8HGU91AfUt7Jpi8ajon+O4Z
q5R4jjEELhSIjg9VZqZ0JGml/oUZvso6tAfKQztDXYefJ5CuHMNV2unYycNRkiUU
dt0K/Nx7DGgpvwVFxQBu/E/MdK4SgUxRaMqm7vspujlSo15cqqsxc1l6sGSFAQNg
h9ZzyK0TDhql0/0dEW0xJkZuevrNzG7cdcDNTu8Tq1Xlrp3suDd1XN+bDnofONHt
KEQr2pQNhxr+JVDkz0bYVpvtVeuM0iqojyy5x2rDj1QrBoPGb4SG56u6NPi0emAI
TcWucTWPGzfpeJKtzk5Ub+haics25h7teUiaRekAcA0wQOTE9it2RfHTk3rjL9Wc
CSAltQrRneWhF/lx3t7Ittk9t/3yg52u7VULPXBexLG+h79MiTK8dFCInnV2Bt3g
hJpME0Lqj8TwWeTQPpN1SO6t4IEBKSKiakILSXPCWRzI7xPTZSYWKdUBYeOt2upZ
/xkbao9eC+tJKDacjpsJD3z0InMgPTh8dIdYO1JX4UZzlqzHiLHkr55KuzIdfaGv
WcuGTY6yIjHV1pr69RZAGeRYUQ+PfnEatBjirEo2N6uf/BvubhsP5QNKDOxjNoRs
4vSnXNP0MLRYG5sIH3URTPYTanusRNldeBR45Gckwt7yQAhc98hYTpTl5pIPfKMB
KOg+OFeGn+NrDFzmWyCggLuGKdp/aE0yZz417zG2iDYJ7/QVyj5JmuCUdePlCvk2
6Jvk9uXstb9TpSgV/nqg+VF2dLn6ETtF9mS8BH9VLQRpdS8jLcHy6NnmCqj+XSc1
sF41IhxK0fUGXBEhLUSMIqTt6B/hjiQLWtElwNBcQ09w1eTIO1j0aQGcruJJjjYk
OCHDkWU4I2kDckQXFLyhxGU/a390QlGgLKA16WibG+vRRwy6iUWdj1fKt4MwHyBQ
QniDysP3V+KorDYkPQuDzVbUSssQrnPKn9OEJ5CLFeh6zwbyE5Tplxv6san87mu+
1hNO3xGtufmVvPMEPoE1qseMte+9mEkbSQ8h2RdnxE8dMe/Sw6V8pEjMjO5w0rdM
3Yo0k9wjQGQM0I/6NBk/Jkr/Qq/CVzpY1XPnc8icXbohDL8HxPu/2ElsBCeYzo3O
TZkCohqHcd4qN7wkjfiGIrR7RZFV8fh8yQll9f08uzIwizyiqG/LERIE0mUhlMFt
iSQKTXhT5/gZEtskiMCq3EMBw1i15hsgmdEE+QNtjR1AJg8WOo8Vd2InUxyND16x
2ht6+SMl/il1AjNBeVljVmzbnaviABNaluDlm7ivy2mYiSEHV4Mi9TPtDM8B1GWf
u8MIvcTrDvpZCEMEF1VxXFDGB/BbWifbRDyNxW1g3sJm1Jg5WzEdX2aAJholLOUI
t4ozDsw0S6M4MLJiLycN5b4Dt1fbYFaqfNgBsKkEwo600bQoLFdF3gA3+1SX3vkw
4SeL/WZBF6dXZ+IPio2593QasgsbJG0/raTdxDlGlhHOy94afMKeROpJ/P/xBOn0
Y0uy3BMfv8JwuqV8kdIXzTos5Eu6G8T+rR9ERAcXIcan/M+r4ulbtLtEGEvzWqkI
QsRjKPoK8x7LrKtwPs3gnWKun5eQw/J2AvfbOd9slqAEjJCoutuxJutsg5EcHUgH
dhttm4Em66IXjdEsJapJIeStCnZX3+Gc5vs/sqHUB6l5f+wP7q6MU4qWIe1vq7ie
k3Pqa+3uFCbJxTGFwHNe5Famw+DWnH7k6InK/nTkux9NM2R2rWNTsDm5mAzOsWHp
BqPTWniVXP1YCQysbk7p8J8v4gmpnaxKjFRGLa/J7URKDRJyJgcfmYCpQ0aGIzPP
nXiHbVB3Qdjz6McSS5CFsTkREG+wnWkYESCHYeUjWf3x7cgyEZOFKdQEDIfbWynE
WuEOqXXukJUTyiUr0FngllRpx2VvBNk9e5H6bz4DzDsqLoy50RI2lnW8P4h+j4vE
/9uG8W+929qBCFhNE+VjZoXdal6QyUc7h8AJDzVZUvGRhdewEYiVsV2cIRdurumB
g2fPMh5k4gxv2r9KuVjzkzT4wpOvINgP4hUoSNuSIBuDoDKaueoB02vU4oLNLB++
qpYYdHuPTV3nG8yr1eRTq/qtNM2j40C0kO//FRhTBFP5h9nAr1ODPL1Gsf8v2ozP
mKAnb3TZzDqcTiQ1byLDvcjLSfgGuz65p+tZQSRGbffcda7bZxm6qSRkRcjcHmTu
ddQb/OtDFODuZey9/cCcxZtYp4n0PWAjcVVUDZYZMEzDQ8C/5IPv+sYZQlDZreFh
J8aumIhntT0CQj9y2nzhgfxTYpHYAWVkwI5D4BqR3Tj2+clrRIUfFphBVTSOwajm
jhyuzEc3tGqyRb5IwGaynYqlzK4B1GH72p/zLJ9DuGxZSGSut1yVDbuVRpNM4xsn
M1PYl6y9HX3QBXj/OwKNNVqLYiL6suOGe1Pr6Om8OEju4/qAjjjcR5+TvMAm8mRZ
Y1AtKVzDEKSXBGXrYUY5164zlEyGIsQALkeva7ndYPUfGzJwRWAaPqq/rhm0S0fC
iDozeKjKYcfo+LAJWlvPZfW6L9bM3G23lcsk7XZLc/ek6uoPYyDw6VSEpo6hCjNu
cO7MRZ2OLU8xhLftLeTH2AXTC4hXO2oQc4GMD5oZ+U4Dm9QQvYu31uMbM8OD17w9
O1S6LAadH3T2AAcE3bN9zJDZgRdhfepaTD9lkzBKOPFH/3e9N04qt7n1Gk8EPfnr
XQgf7oFse3vjaTo1roK3BdCr214ExlDzTIR7R2XnPZS4s1IN+PWc9iPlhUEAzz0G
44Wg4z+C/wrocXvDNgB+HlxeYfeVV0lb4peimHTfdzJdF2VEF+ZgS0MrXs8akoaz
up6JlN0brt9qp0QLuV9X7mJT+ArMinQE2bLqduCx3OXEPouDCMdw9St69tlTvci+
H9P9OZsksN4fg3qwOn4stby37AYp8HIaGw1cXG76ZPqEKJvyURlUX3Y1Tkf98+1u
4xeESLSwD9bH6flHpqdgr3ptO7dkCrGxLzKnSc7jilccEOlsg5urdLDitSKYVNZZ
yhvhiqv8PTpSw8t8u+zk19kOkojXWDuyuMJDRwxfPxunmskbHZaXfhzp7l120M0y
8htee632cQaczFKok2KgQc/sfHmy1GRrCS7ZfK8+ZI/VIx3M4nUZtNh8LVyxVe3x
cn+JD6gavk09rOl4aJVGJaOaC90WZ1v8+87pnczhoE0HulAz6zFfMe4HfTNG3n/+
b+bJaevEi6a54I+61OYy2lQ+xJsL4yr16ZmAyLqXldpQNvHR/wCBI+BaGfB1NMG1
q0jTBuOg8UXmtx5xP19IX8ypw/C6ip5h7vRL236sgSQHOILXhNOV9W42k54jLzlk
2Th9ZLN1rHmp81mPnABo4/4L7XlmTVC+FWYn4vx2uYy1MLgqX4fB2ApPlM2Ne47K
+6mflicni+umnMhVQxyQKUwcRXSnbX8tmfj4bhJ4oxHQsrEXHMclBcay57Y5NYWm
EEJ8QQNGLZTaqHL0tyGPEP/rQ/RqoBUmZbf9pjjctFgwlvdOHLm3ncMT4EGaKJzb
z48wB4fbiGtxcxwojsQjpzAzysXkjTgCfH1xYLay/DMapAOnYi/2LQhi1dBiS0Tn
OG00RY3WRK+N3KY4FYzNtjpEboH3AAd+WA/6iYduktODRXDNQat1nffVpB5IcmLC
DKEPKutIaNqr34ZwNj0bynamJOmyd94RLIyzho1DMVBRaa3+kQd9SxRiHG7kL/04
Kj0K4Y3CVMDSQMcSNAcfy9xdQZXtRszobn4b6v0k1MRaRl3uGBJNMBijEEv+L3eK
Fq4e/oHUa9gK4ZqI+nTUbXoKXLcjRy773DA93SsxVtU8n10Ux0pXxezHuHiwbSNt
hzmjSoQhAdN2VM23k1kBoCHziZ3Z/zxTNKUzQguItDBrD1U8SitzyHHTJk9V95SP
TOM65xF1HK/XOpyZ5Ie1NboKmSuOfXKlqtCOkc0wUXp/LJOGrimkMisTZBid4+M+
rXAwKHfKDlWt0sz/IvJYSfpF/QbBObLfGN8ciHcEJbc0galLu+MZZlRQtnFcrYm7
6A5JxXn2kDIrkaZfyBdWBU1AaXQDgOlsqwiqUnSZ9RkLYcubEFPtnldWjX302sMX
AAYWenGaa8WT8AVAkhlwaoWav0o9CQ10Kf0xfW/j9QovlJ83+6B9FaXp8GNNOCQY
gE7KPoVhrRQBB89qRNeG0GR1XcKiXI+G8UHkYOXk+1sWRhYt8zRh/bpctMN2j8eD
JpGNGae9+3n41tYblWQlRk/DgrosGH9MQ/w1VDWN8MlbT0T/seRt6QIZuTkexkZr
XSLpNwVw3//rzaMgE+k7hHu8fWVAjWTAPQI9A3UNk600LDP+fI5+Aj2AuzZvfHfe
eI1Asgfc8/ysFaWI4yfJIBr06F2M6xSVnlvcVdACyMMkLXvjVwG1ObH/lOOq0AkU
czx+tDTA/KlRHNQmQY5LE3epf4AbIA3DEtmfbsLWzzdiqFJAHKI5AvGhmaVqNIw5
Y+0InnhAqubudAkj4H3F8XIjDxT9vAhqT9lBqIVLZAYgmDgAtQWAWBVoK7b10ql2
i0t6BgBPPXzGrmXoZqUeObbWNndrhAq/KG7qIjKK14K/Nq0HDB3of/BjDGT8vKzV
JNV8WUph6H8oxfnFQuCb2cZSF1eV+1lRDR12AVg4tOk6Ua2HOgf8K6cprN9qVm00
TxbZ30zJ8dOHeRKhvHBzcn4BzB3fizl+dRYGc+Dw1PWj+XIyzbMczrQ87pXnfh34
D9HnDPNI+5R7PqEt2GqA+5XlrmbcY8zlcGipXT4Gm53xGJzjwhdrZYENn3CJuXDO
zHrKIh23VLyv6NPFI+1LFY3wjdVH8jAE5xfkLr/STs/pJjQzbM0HI/V1ukugNLcv
p42X2wGEZIE1AsHiTQj1Dx/lSdK87G3AcW3fTJaj1AigAz0+gJJaqqaNhWMPFKCy
k/MkERyIEcTKB5rmzBjHCL9HGqfMYq9aUJod1LWkOq0O3CVz8NugzYSbF4rT6wXz
eNdae9A5hvxU+4bp07uzUHyrGyPFnBZ5saj72OL95KInJV+cUdImDz3yEPu8W9Mz
s3aEyaUC7xv7NucYAxuad/x2iNoBYF8eKD2kMB5HhjLZ2dWlYwRZRflrEGAxBdw9
fLcUThu/B/FvAd1Ruza3wZ7oXYkiqQwCVIYcKTZ8CqhBZj0XyBwKNgS6Pe1vMGqh
qv/0J4VfywYysGs2vCrET6cu1btT5pzj83ZJwsH8qOJJ3j31/dRwXoMgx8HZpSyL
KFlfS42bCAfwup2XWtR6tDdeX0cpbHahaLRbb6Q/97Gb+4pHNAE0CbY0Tf9XICIX
4/+cFzvDYm5naVw8+SEe8KfkGbEYKVX98vVb91II5yk2yulAb6iulFJiMUbT4dtH
TjZG9d6JGrDGy9ZLFSVoC6bxC4NjojulQQY9XUZzPTw9ZKNuqRMNdQv8LJjOUIbV
0hbj52A6I9NaiJBFPwuod+cEKkcue5tCNwXG8ZiFVZExQhIpqBVx9IqOXhO9HKhc
cl94feYqn22rP0j44whgboWimqQl8G6AHeEtmtezSEqWo74Moulh30Zxj43geUI6
0++TRTXroHXCpCHicsD7zgzkdR2HsMie8qLNOmjeP3ofkloDdcwLrTW5sgiZRxII
dxrVoj63yqPwTVQ+pkVTPRO49Y3ppN6rJ05HyENvCZ9n6fo3uAu/p8sOb8B++k8Q
Y6bQMRJ/NQ/xj+z1mrig2r/FRoKvBi+erdJfeYOs0xiutZYVWvg4BLI/7InV2iPX
v0WViroUBydOrhmMWmYL9t6eNxWjLgeyUTAzbBARXN4DvuAx4S+9RU1CGnaRTFob
JrJpKswpWIzYsGbnhyAWbg3OZ66s7BYvFUQSSi4xZWzlkmf7ucr5/wIx9xOuAASi
9VnOmybxh7D67WFUu1bfKxCyU6swOsSZKwYUzrLQphnaUJHRfXPF1e3bNhp35rI1
KomeXf/7wIKdqLvZyhpacsVaGLOH8a6sYqZGuWvMfm/FUo/XyjrhRUbVEhuoHZAd
EorNA1BEuBkrAzccriwKluxN1RGbobT4g+NzlD3TNtCX+amrIETm8flVqPvktwFN
S4dmhg9PwepgifZG+oonRwQ0ZZEo6DG3BZPtcXQ9ui3/cH7NzNpGLq9cNj7SuUYk
NPQGhib1ipSeUsQcQR+Dq12CRf/xpb7fX2XN1NzjJ2j22adeKldej0i9NubTCQir
QLTfNYSCbRjoYNCGQVVj45talEXuQ0IVWIVGGnqe2/+1fLQxU9+qODAHHzhaRz/1
gwU6ppUJ1sZel175o18YPmKZLwcNyKw/6kRsgq6cuFoiOwQ7FtdYIQ2bU8eCR/je
M5CJVyDjJrlCGK7QZichYbUeKxKZOlLg201LDYvFxFkFoNq03PjJUAV2X3ve1Nmf
bk+4hlFQoQM85pCEHf/ofvTtRNYAlnVtbfIrr9byl1p3pNASEskCJ6zw/inKhjjs
OwgRfGmfNzi0N+JxMrnd2Li8lp8oD07MmqcPLGuYVnA0DBmVzimibXQMF4OQf46e
lNo2U6rVHssHgU06XE/4Mlf27ttlMCXa3UMoYjyJjMEnniKjHX/jdMgJMOOh1PCk
iUo452OCLGsl4ZxxdyhBAHLS878k91XVyk6rwqYAipomqXPZLBislPlu7zerEB7I
ZafhaKDq8tDOJycUtoXogAw/sE8fa6XY9hPNoNziHreC4xu4x2Y/oSaq9qfzvsag
qV7PZVCvGnHUnjBynLkEMtGsvFz64cw5cz1kfXeuB7grZY6QFPQB+nlU1nzSd5zh
uoa0etOAcKtr1Ey+2V2rFdwLB9BKbOpASOCH3S1CPwRJ38t6hFcj8ZX/Q0Laezyn
jGKSfFIEytT1i49vo74f7biq4C07i7/2PuyiURy/Qj99iXBTD/IW+YbOvvnXOHmz
NMytVTSh/mMZwEEMTkL/I5fQlAhx/MoYGqNTvtcLMgYybI5EMxUkm9KmxL8kVrR8
DwNLhjYQL5LMtodaoKMBOTvBUIWwb/P+JV5I+5qWgmyPjnyX1+Q/MHmDU2gPuqEo
oYtMEYNcInIx49C3N5VM0YT5VA9FkhkuGVf592YDInG0MVGuksrAbDyZ0u5iC/7l
YtLgjeNGuUMfS7U33Kmdz4dNkLp9mRVf8o8f4jUpxZegJYeyjq0QYapcg7y5kvof
XytQ3iSzqIu47MZrAqWmF11P/Tnm4K3l3qAm9wHPyseyt53xQzPDH3gCRv1JdB+C
Zyjf8bbLt7pzl681EePWthkaEn8yKj/06sIoQOHRJ2tSnOXoI2OkOxD3w3hd2pNA
RXEmY33xK5/LdtACRWsqsfkJfjgBAItbGZYGbUlYnq0FuPlXQxqTJQ78JH89aTcc
N7380Eh7vxl8eT9hXbWgGv9z6HTxp6s9t/j40cbXGk+RQQ2SW0308TTr5fkjX7ou
SH7c8u42unSaqqCyoit05xRzEEbvM5Yf/PSVuV+VVc1gTbJhpnnKkjpcj5LG3yQg
O2cZ4pM5gc7LTLd38vh2t7C7mu1ZiVndqYdBxN11w3rntMNebIXcIIZc+bCstRgh
CKx5YWTH2ndQNbBsRVD0hJjCmhdkwTWTl4o+deEsnc8nKhFOeTlxeiGnL5woLpOw
EWuMUCk8eeUrHMo6TL3PsuuyMqqN5EEN8EN7pZ+qeLt8U00WAPve+aujUoRhu4+2
XjbWUA0s/v1Aq2m7Hsotn5Z+DqH7O3w8RgZFVfNB6qP0iwJnw7+dDxD0ucmsAxRe
ErAAYIV/YMbHNvvnQjSVe00VebFuvj1IQlo+bOGSFhuWrm5y3uOApxDMjz8khQGM
5fYCrsmZWvldjxvTrl7gZIz3ViwmLjB0BpkCLN3IlP1QnlC/Uf/3gEbkqX0v8pGE
KFXpr1saIj4kk2uXmwIiZ8x/vcKxvX8oJ+F0TAmEC/rzE6O4l4+QnRgKmjeW7eU2
GcveU8LkA4KEVA0R7e76YBlHHeUx4vU1hYhn+I3BCL977MXbpE30uJTgQFJFl36b
4vDrqLhRQkvn8QD/FMLICjzxkKXteK7NQb048hZpfFpcW5LC1ZWbEDFV+DbrxMKv
3YmfwCGGgDdLrxPYzpkvWx3A3JGeuZDx1B4h0ByWfpIIPcCPM1w1kPbytTn6khuS
A0takkZTRwcdoNitHS+ndiV4n8jnhlCPjxLrL1Jo7NzPODm5KSvT23WpaUo/hK5M
ewW8UbdmwI8AiuVLasyZg9pqfZiy8BbDp5akhBCEvIhrxZpA0yFSos486OxiAZV+
DytAXzxaiEzBZIgBbLANy8td64eC6+pRVYofwTwAvgXxjWpV/8KsXkJBnTahHOmc
9kRmENGEa4cSdDXACmQZqwaRqHcNcGzwy7+GulsXiDSK7w9YOsQrZ2dokbZ3szjz
EfDIMbpki01tk8zYJJ/g/f/QJ/Wpc4hBG8KDDqaQANiSJaFaDvemHkZU964irHNl
ZTHDgY+5dDvrSPzUMUrIDTxWO537SEpT2trsS525WVxJMqy/9YF9pI9HQOd1gq+m
R+kWcgGZDup+o6iVNYHB8pKSVnE4h3zqNuPjTPvsi7xIixjmri+PlyJNeiezSiRG
nc5N/x6PRik7wX/JEkacftc+TjUzJcCoxUo28DppAR5ywFm+fR3GyYrxdl0afCXi
HJCF7nPCjcf4GCVYqJqFB6SdQaKkkMUEBq94PE+JLzundH11D8AGpig6bMp76Q9r
8QCdnSBhf/T4Me0dsjZNEHHDrPHsVCSGfkGPazb7zYfRs0tG7yiWNL0RXFw5QdhR
yZRTn6LrwV1QsZFmB76RG5fP7y8/kCCDpJAI+h6QAICk5UAwLEdArKGRoBE9NF0/
Kx8GjK9vNqxIjfT1Nc48u8XUvP75fQ58ur50T90xUPMz8wBFG9ofU+soEBV8ij21
5XfsXQLc2SNUcMHMlJx1eqBn/mskFDuY0gPu786vhJnow84Js+lCA3cjozN3yeT9
CPrDGGfCUYi3rnQRNh4J+3YIPCZozQiQcWtBdPBcv0PZAJdRGbD+QL/pWIugOkTD
MuacH+YLue9fwUzoOGDgpbWaxuYvDjJzJ3aJTw36gowLQgpBwbyDIpB/DdM3wshi
KwA1TgNmzauZzKAbC5l2QPmlIMKJDQYWg0Ye8wmstbfba3T7+vJrfNp4/BePr+Km
At10gjomfK6cpNX/8ZLA7PVniWw9ua4K6+EnjKS4SC0S29NAUf+B2q83IcHKd+SM
6DKNoOGKZa861Aw2zUdExIlHDF05oxVAEA7oD8iPfPmyFTM5dAP60y1txYsYZwFq
as9SnreoJhraVQN3Eoga76UVI3r+TMwa56yjs5TK5rUyrP/uMCTg2LMMxstxyAAS
zrqGGADWolz0gy5Yza9VwRiCo6J91ZlylQlH0GEwkzw3EkWYem8rUL9Jgwqi8/nV
aiO3gPf8vCaaGOZJ1gcVgmBmwFQq0CVZ6Z9W/fB+WLTqbVjHUXi9Thpn6NrJk8m3
27zuCCv4ev9+/VASzCuzxq7l7LD4SVT/Xlt99ZyZxtYYLl95M5rDfiaE/GhnrwDO
2VYhmhBI4Zbiz2JEt4fsuws7zuF0a12QHKEMwtcJDfAIY+6BuCSiueDU7wY0jQfP
iChX2HOFuYPA7uYJnjFtAawdc+fInZvLWudNUGcfTaIwTcZE6kF6pl0roC3d0lGL
lYDrIah1rvMS73eehHUZsdxYb9V9MyPKocRwbZlsehlLGoBExWW8SsLoU/MQPo1Z
JeIQ4ZjIV0vt5cuBiuIF1vkElhAf2sOEDNXzaCwiPqHWJ9bvv/tRm9XgDaosHdR9
FCnc0RGFQKQ0ka+rZd6Fa90WZslo1stEgYDYqZUxBkjMszioWoLePUcUKIs5MXaY
hVxK/mrGbo7g0P41wVJuYHgizYtIewgsQz+SipZ4jwThXPF1xlRaY4FrsJrtPZfx
cRjhbsELXJ24G8BrLigqJy51gs3bLA63HFfO1ztqqSRYH7ER/AQROaZ0nCw9EV34
6VvM6e4K7HB3L+XyjFYOWTGh/bA+5rLo0Ga1RXDnRE5BdCPSvwnPTPAv9VLo+pTW
9/SQnIA6HUFlDMjDcqkSsgHB3gmSb1BGOzyzFQUg8U1muAQ/8eWuYPbv8nrSF2vy
NNXfwzAuJB6uhQYuNGRqVp6Sb1MDX6+/Czdbx8LmDr1S3rsnWZ47vw9hwvuSTnvL
DkvTgsoiNa3RbBMZWNmVPFEgRjy82f6ht4a8CiW/OJTJ9FF5ubeXkM5tTbiDM6tY
BNmwDY3YiEmEwi+BSxNmUG5UeLbquU7dw9RlRZkOB2IgLKCc7+iIblDWOFC3GXnw
wTcVG+r1v/nKxanJf7Cto/NYD9OJvrpk3JeOGHkPS6eS/Zbc/IOH+gvdXoFoY03A
nnkCXehqdZ+7PRoIVe139PHrcscIjO2Jp8OOZ2kWtOIX6rA/otY0lZ+AOpntyvec
jCR+7eynVPPjvaiYkdrJ7If07MWNXIpf2zr2a/AHIml7HFH7ENt4JIwGzzIadUep
v2//VQvsiFtzqGU25SS/Vgwik2C56uZVH58WpoloecjchkzOwSYgJ0l7fG8b49ns
JhgRhBRuL5RhM14wa12OfiI48vOaptZD0VM8Pe1YMa+7kdtRW2CjLlwNJTWt1Xym
O0LMI0y+ARRJelDoYREDiE74SE1KhPshk0OY59HcF3/osgkU/4TCIsKUGDYDeQcM
XgBsUATWuHtP++C612PR9v2zwgsZmnYkWB43EJEcajI79rac35YCIaOlk6B7mqbp
IgECf5P9AGr3k44cCNDFM1fYIM/r9kgQmQF6OkdsljYjNV1XTbP9PklGko2obwM7
ihch6mDfD23iXiev9PdzgrBeDuE3eH1PrX0u2l98uxsAFFptHkGLNwWzZp99K7x0
z+IKz2mkk4+vofrvmCzQzuXEGGb3Pb3vGq7EI2MC9ZcYBl6JiVMR9RdO/0CCGgjq
cDDlr/2QsaDvYkACJiqStUjbE8VHUBhllE0wRnloxrXSP1By6Sw4oqlV9B5TxTHT
dbLQHnUUEnuCoH9W1LsWA/gJ5uvIcKvPZ4vz6IKKMFUdMfK9hStz5snVQoEWygh5
xz08xMjTncdV6adhNzzwvSTfwA0/+JnDDg4bzk/O2KwCjjP5nmwHjpVljNRqqgil
w/Uj+M2yCTjPiDgxJTfWPFM4wKwp5sDRqiER70Jkg0OHOdDXZVSrxQC2UzRfb3Ok
I/0zX4PqwmIR4p+T76UJQ8YBcPOVIz6c7/ulicMrEM8tpZQ5PK46suCPQp3PgZdL
Z6Bm0bOXlwZ+4V0eOPI+al5x37ZaS7zc8IpHpmRs8VzynAoaLOcyvmi8tgXr+oNo
HM9rmbV2PRQK7wCKpUilZpuq9SjLcgDyQwzObuAVPMf91aE51jsTfef8JNjtD9yh
0dcU05s0XoUe4JRp38G4uDqWhSySJH1QT4wP6p6EiJhaj7PGN++eQKMK8fy7RFFE
tkck3BtBxEVWYNny49luh9qrnpoEBzAQoLsDzrX9KGfebXVThukWq9z7B7CkT5ey
A5NB0FK0u3RcN1KHH8zz86rXJmOvBnLDf9HYl1J1iXtglkiFOKR1qA8LtSSzt0W8
59dT1N0KTTwEGZtpt8BzQuEX1AmkCWcNDdVcUHcGdneR9w6mEqiFYiSS+q82WYse
id6Pxz4+mf2GSpwF3idMb/GIYr++50YS8wZXkZGM4en7iF3t8T1Djy2gSrjp5pUN
YibWenEcjthmF84JgxNdFs6gc3+w8J/IPyd9d0Ep7vXFsr0u1EVwsQv6Zv/aO60t
Rgb039Kzx7IVF3HT/7QwtV3v5GdBb2Akwq8s70RJEZVz3FGekW+AGtVFdvgyEkwV
ZyZeINkXQnHsuVGbtXEyZsUXTgjBxTwl+9Xa5j1WWipPdQr0+pV7tBfcVvtXfHCU
qHLiNwevV4IRutb5Bo66MMAigNPTWSgUA4PjZAdDcm48Q77bZ5GOJwMR9r6j5CJr
SlZipMKuzEyTo1gm3L6Y0O2nbU+ZztXuR2U5IoypYBgjVIOivC/5ChPVE12C1NLb
GxxhyK/Ei9rIhL2BT8ZPkk9I4HP+xfZvpGSvJBdhPz4s6BnoTLJBFBWodAhS9cbA
CU7b1CWlId00oPyM9Q1OpqOKNHYV3uAitxVmx7j7icayX86vIbH5gwD7nGjGJUYc
f+2ehJQwG0RpNWd7jlEojiSNe0LK6gVirOz2MtzxBTD7hnw9TPy4H7PCTFCoRBgh
AahyFSTN+eN+meLZ6DRgd+/Cs+I37JzaaOwLTJ3LXziIP75LzuLP0Ovi+Bju5QWU
tK9z4F7h+TY0K/iU+HO3UpKZg51fP/2H+pnCcG1aX4KvfS2fmb3RnzS76VEGcai3
P5nkT7AWXxe+IQlsSp9wVkl6d+g030fc//rpe0QpKrrY8MdJxUSdKBSaIKyQGeca
yDMLPYgNuRTaccFq3fWgUL0BBlKpDKsuG5DPjdfxZB7bYLUi8QZj0IDNdwaulQwc
WZx4SmjbLl3k2F5hBdSRlOiBSDhkL7TwNEeBEn8n600MCaPZtkbEc5/4K3SYL5T7
TH+6g0QfM51ZXtjk3r1xgIqea2yzjfF5M2e/wkgau5BxxTojhawB8mY/emmkRcGJ
VVG5wvxly2uCLjxgNdNuRPCgfNF+5fS7Nk9QE4fl1IhPmMvEALx5cEBCj4EEN9mN
GQAMnJAANHYixTV5g3CRDkRpHJw6JPt6j4mLxZzMqz20QtNXpDf111sRraoZekkJ
KoDXesZ5cgGFDBJQry0xCnVS2ce0dOCzKsFfhCJcVOZ69GYkr8kDLNOkJNkI7jsp
H4vFCTWSLFZnaG5mK0ytubGnyPK+C3sqm4vwvabwV2iSKWVKZQ3NUwy4bCQvkBQC
zM646m3mZIYLymAn9iG2zOBq5mQ3l/m3W165nYMGfCupszg4iNA4xRbHdXhRhf+c
VGD4zaHkSefvniJAc292x/SVM9plhTy3tDQ01P28xbtXuK9WHBnRzMAhh0/Z+TE+
a9pJQT4a1H4Zk+THDfDRCRwPDL/KmyuSETDYxeqX/dm1ctM9NIjYS389JQ4VpNc4
u/YFJgnhYYZMzIyoIcRpPG0p9L9m/2JvFOmIepKg4D5C2JweNfOfj8QyxkYSEQn2
oL7MOm6VgNHdwu9sgRQDtEth0hAr8JfIg/Vuz0ZsIUx1Wdb8guNuu2ucy7pVlnuh
FU+O9QynbBZBXlLn1t5epzmG/FZYtzoUUuRgJcDAcMk/6xMUBm4X8XaswORKLKZx
mOuaoge5m9xeAoyqvVlmtQkqFBqx6evwmfC5zKfuEhcvgHJfc7WPltbcmTfbenu7
7c/lszJtfw8T88Z4TVdX40MGVuG0wsu51hZZxw5OB3BCSuYIspuzM2ZZV5Ce7xl7
KY/6QiKyT34NMity2u5nhGKS/yF81JHMZQKufLGwZgxXHZmlG3NcgKwhST8qoGDR
+u46ImtqjfpFb5Gtcexbe+j48LjHmnKpgeXKZ8G8LSkxYgV2yaUjYtBsE+SLZf7U
Et5NJnMObt0pADuuiIxG1iZXV90MHkbXvNJzg9KWU1t6Vlwj3zRlf0uWPeZkgEGR
lGGz6/9H/O/xmChgtazqPVL5F5ERQFrQ30kTwU4O75S2ATyrCY4XiD9AJolHshdS
Pfb/iku61X5AyeRxCTX33Xyq962DFsqqbHlTMIwMWCR42HvbIJAlLsEx7V6rqzp8
InkaIoTZFxvI2CqKeCKyi6gVtSd0RDW+/P+nlRM4AZg52IlUvTQgE5t8KXYwKjzr
SeIkYtowHcJm1K4bY2afIz20A17WsR5HEgHOHpWSu4Bx5zYGYCWaEgCBaHweo0Oq
SvXaZispXGDfsWBI+rR3WhQ1ghfAZtP3+HzbPFgNpZkEuZdmWIX+zQqI0tDyKVjO
5wz9BnQpaabB1ACcdabzlrg3uTsz8Li3wcwzSAxRze95dLLUy56eZNJK0JvfcCEv
dKRlKBJ6jIf28FmcRS3nPczUvcZuKnvgAu6CsoC3+mJbXHef8l0FZD2+W/voJXnN
X3HUpehCbeusBq00PCy6tqjXQaLJygdaCUq1UH4gYLzJvQzc0JI1OzUnBX9PeP2j
0xvie12kSgP0ha/rHcugLMOAbpOs4yYo7X/OwZTKQryiBd9a/YgVglyxnasqr34F
Sm/7khJlXqRsyrycXf88WsM79215Mn0Ld7R77kz6TrzMC155jFIh8yKdGTVpd7Um
B2iIjWshITRFfdszJ8FFQumeykYTUGV03uvsAbgQSQ77Pnktbqy7eEmCdbA5tivF
4SaLMeLzKJsgBkTQnvtZxDFJ6n87GlWUT90+g2dGapuUM6FFukIC3HTAvaIDMToS
A0gRztcdH+nEiQqu9OLPVpHqudWHCUcwTHa7/xEtzgJyqEuLt0wYZqkG2zlNAYH/
UuL7Mbkxy6Jmc1yeJ7QrkpvvSVAX8jYjFaKjUmcF3aQhhwtFfFjDZaHh/mImdbUe
j1cNz+qFxwJabXjdtpHuGV0EugXXV8fCasrfK+uf8r/vthPHYlkGiWe+igC3cBhA
IeFL3Jlxb704qz4n6tt/QSnsfMXxuP1vHiNfQm5xx34Rp7TyPSpWaxN+hS83b1XV
4EgHdAE/22wkB+DpkiDNUrqPXHNTwO34sici+1zeRn/0VJLpsaxCtN3L9xY4ylG3
98+vEUFDhBW2Kj8Gg4/b0iB4VpsYPGYKhihkyi72wNqe/6EIdzzwMXahz4UcCLBK
GzWviFCx8mfEc/cCCwcVA4CwYqcwpIjiJDYEyClXAzZZF1sooYTXfUEIzLg/jpQu
Oe7MKZ5UcCItItXnB97QUJRM80WkKvuCk3Qnguq2xG6+P0mBb/kJOCtLYD5OQl4e
2OtCW+F11nwG4eywYHc26+cxv/eAhFEgG4TvAYSulaBGPqnLjEUYssG2zyh+VwR+
idvHOFrjHRAKX8nZest/XcA0YC43TZD/8vsmTZUIIHOQNrrzgp9eK+91OKcA+ykF
9Oa2v4q+vf/rvjvI7rp1ZkaW60o8F8qri57ALpDDZh22qOE+Bc86iJOWfJGePvGG
bDcpNglu8vH5QIdri1UXfUVdLYW/dacTPhumotJGL48X1vQNK3gqMsGUF4CbC9rv
Y2jqFtrpOj+7wNiZ4JAGwN7w368oXPGFfx9C1b+mjBU0p2v/735vZPBeP7gnIht+
H8oYqCNolxQEx40XFzl4AZ8ipMo8KAFTPmad7J3mXMRPUdhhThiOOOC5cm2OCnSY
CAljR2wAAUnXvcs9cZIiIFgEJbj3WriGFT4zSBQw2kjtwLVd54dkdBB81XDEPhEf
ABItigOE/c1RaDCZ+PPDNSTGnfqkcbihFKHVZwxJCeI25gMooFU65oW4Ij0wZdMs
IHFAjYH6Pg9ri06ZxYEOwEImvCTY9LY1jFnmKPFa9YKBHtOHdktZbsft0e2vYtBP
m1cuVVbSf66cN5GPlFli/4TT64mrR6Y2Dje0NXDpOXx/tbCeFKyq/51L4BqMz2is
NWxV2L6fZW6Aa2ZdPYjfrlIhR5LweSz11HF+zbZNx7094tW/rCQqZONhxXsF2wy0
wPCcRt7PedhDcz/xe1R5QMUDKcnas/Rh5ldXsx1zK884Lwphsumkbix29D2MN88O
Gd7dwUHHVwDc9Ui3zS9GqGJUbeQaebuaRzgQCUWD2+ZEOXOXZEdCMaYGfV190tdQ
xJFMvQ6UYsQs78qyjlzfSfiuU/am/7inOEc5T8ge3w6dsJUyWbNIDoerNpIDbH0V
G5tEYs3Y9xepzMA3oAmwRwjE9Hkg2OXkif6SbtGxQ1h0D7PMAV9HEiJ+p0pxVKbD
/vIgSFhHHygvvegoplxRfAjves65eDSLdSzI586S/oMZL4HMWoj/jWuUvxYj9WRx
tBhjYYSzihx1/Nc53rB3LGJVPp71X3HJHLaQPQqY9j3004MnxjWoHPiCe8iBaD8b
COwIslXKvdFFG4+qB8v3SuCV6qSwr67s+UqjlEK+ZZDtBDpUj8bOCrq6GOgqxEKX
/5kYwD22b66+eKNLhyO2sierk09PHy5QEqi4/3OYf9S0vBQ337T85A7/kgsn2a0+
eudD9AVkvo5oZrYNmkhp1BlDMe4qk2/RizogLO96yzosw5z7+JclpjGrehBPaA76
5kOGs7HNO/rJgqBUzU1Tc1eJTZZEKP9qWZCMQDC88F6uFbcbifwW3ceql+QITU1y
KsSXZw5BD2E3NcAdREzfHaZLFf6WSsbfQ2BiHJtPHMmsVhxmq9oovJ7iEwBY7RuY
97nkPiq8zZbQM9iia8cpZxxgyvL1xWhjZkO14khsDDJDsYoosGaim/2gvPYurDwp
mACpIxrJ8DGdEAw1W+ATsCZbBb0hspbpOppPZpX0YwBx51U99iiOG6O2BFNa1btE
H+ZWmjO5VMzFZTs3B3GJufCdQb6UdpxRhpPE+dwKRAfZcuQPH8MeziyaubEDsCn6
TSx580xuwvkm8gfXDa2W60w3qENcr0X6FfZqYzzahEfLZ/Styjib4CxB7lACsk6q
JGDNkTzKh85qj1PrJyES4NqC1bMONkMi0vSD4SbvuPkoGaPMVnEaPEwpRpA9Ge7r
Uwd9yDlC6orcORdJC3Kz1fptM5BxNSYMyg1rj09G5K+P8fryvNak9SQN56oB8pRN
uHyl2VtPgI/GIRD+oPxz0wz2AxELcVC9EBtxWZ9LZyBhTQg7X6r/Nxms2ut4y6eu
kTVNSCP2ix5yoZhyiDiRm6KXaJNjxz/IkApp07CcR5rjZZFr3oaWGrx5bsxCPTBR
zX4fNL6+NmQg6C63QlS1RdVPQurjW0qihPhhvRo/eoSwaN6gVsj/TCOpwWdIw6EC
8WhwCi9s3oVVsqMpuKkH04SDpsl4fsdTBJpcO7vFCXvX8+NfexcSgaAqbotu/10M
h1p1yTiDBQ0pbDkp4O5r6RrElize3VR5i9/LfSpT7miVXyvpGhDKy/ySdaWIiNGr
YtsU/6URG0YdrtBy7fuwJXZTMuZRnfHp1Al7GuTUVaStkFJEmgZ9NjthrVCgmOF9
fERxxSuvqieoWkdfTzMKJ85le/p+R0MBOyFrnmLRlrX1RZrw5XPkqr08V0z/lS+n
RbrBXNv3egHl/ubJ/8X8E6GxL1moN+F3ylDtZX0kM1VrnaDs9Cr1MwMEVJbg55lY
NP65PrTm4pCF55m/ICNJfeMorWh3LPZx10r2V9B132ZYDAvIbtwV/bBo1QlMZITB
zzaTzp18EdONV0+6GQmPeREkH7Uj0P6Sfq7pEtRyNYMhxti8Ww6PP5hZ6lYwMXMh
kQhC+uzAq5BjvPXQ0ayD/iHTDiyD4Qx8Ah4UCwcw7okU5jLRSXr2wqr9ISnDjawf
Iv0ts5MYK670pq4YjCBSQA89/N9l5V30/2O6Z+Pxv1QTDzJkLWj0Zt5dEdo7TNkC
JCbU3WmkG2Z01K/BACJJIcqxPLzn586I3xqcM4z5EwabCmlumqSCy72uHUXvn33A
/7qyd09Avtw8WJWTlmyVyG4m5UWyFhAu5jm6K+qpwIvR3FXbpbuNUWJ3gb1UMYes
aB9gg95wl99lvGJWdjmo5g/ahWmlvgQeULV7Xc0kspO+Iw3XDJujzlODpKbkV2RV
tTrwMLVU3xE09K3Pr9eFZN01SKEPeBAd/SQKZ3g665S7k5Jtr42qBnSnOtPTumxb
qVlLBKcQAcxhaBa7DdtqD9szjCjE+WkfhGyCQm4bzyTLnoI0cmkIZqgd+317AAlS
ZDzoAFxtx5fZ9wM4StEmU8nUzq41Nl0utyy3JFLvVhGZKCDGfsm0uIGE5sfhO/nh
EQe5S4hxfR47gESi/BxYO0nXXujpxqSMbn+HlZC9kwswnNtL977glN3noWH23LJG
wmdY6UIzWeGv6SIn06QwB3O9J1BpbDvage+m2nBbs9/elkEeFs9MLIw4aImMHWmA
MvSzhFSqcAYCVskG8P/ePnBFnrBw2igPYxgyAwLLl5j4WXegm8LVAZoZwTfPUfV6
LvJQLAnIMV7B7GVy6vn1S0dZ6XOb8rDPb9kG2thLGEhfLyuX/CR0b/5nzBYtiZIA
foWx5LDjNo/v8wcKghKJ0GCosQaxGK0sz3fk9n/qKFUrSnMwRLRwxawbk2UZ1EPt
ABvY/9ByLUTS8MGGyiM88yBh647a9BtqM64jz8JwIwCX02I7P1qBS/zYBsOpNMUJ
AFuTL/8zE2PEhbkUXONzgnzj1ubD21+N1zc0R/a7vFUzMBnV5N43S4e//riE6lfv
0oPX8v/zRBw7F5DT9ZLogZc6XtTuYosqi1lD+edVicR+i1dCzgRskFiCqkyBJ62e
Rp9lSrQgKMGF+cp0pGsulkIECX/vIa6C0Ihz3samOnPnT0PESsjl6z6pDSW39u/Q
/Hds3nA7P4c+1UjxUCWrTsDifKu9S1Hghxsn1x/GZjRZR+GmGhr9D4tbmu2gZQff
YvAAJa7oleQrxf4q7Pv51fQMZjXkRiuIoMEAeEDyphsbV0cr9gnnDqPYldd9vOoq
EM6bHmUlKkTXg4CNqzs1WkM4aL3awI825ItsNRvWN02tjBNZB6pC+mn8g96JhgL+
or+8Z+2hL1JC1xx7Oh8irvc8QnVmxeGir8Ng90a5lR7gmWA6y1bg1KQHyd8anoIy
oFIZhsDxI2HI192wQza2Jmbc7t1KBTOnTrvZ+WpFYICjCldPwN/4JxXOd8mkNz/V
+BP1P+1zx2AOAOWXBBd96HeGX8bxf6oyWTPECm+MCNlsJOmBQR4s+Rl48Ovp2CDS
H+QD/XZGHcEyYc1R4uYoZULyGI+f3trzwH+uXM8MYN/PT1OBX8fsI+qZTIafxRhf
AHPzLEMt7fsZfC6YhTkXUAxCcq/U8iraBmuZI+hcKV+jGVDs6TrihcB5FjC7I8Aw
u/smJNI9nLvDIW5VR3ZeizulQQXtYsh5WUw0qXq2ou8TQ2HHSO/U5rNa1tsV5kWQ
/Bmibz7olJ2JNUIAJciL2/VxEMl4BU/AbWJFMYNnIjRpwtiV6LmFQZrROu/rdzO/
i7mm4XoEt5/GF2/7G61PhtWrISfov/HUFc8g81NRJJm0gc1jdSljj7bYsPPcACpH
0P+kyDyWmAfMEezemuoIjcMz8tJUtuAj+i4EXn3sw8mNASiTz6DKIK1NocPLYMZu
K/+P14B7CX998FUnjfdr5SsWYrs2tENh5mbUviMXU78iCcyw7/ZvHZQN9lzKSXaz
+WfgvZi3WrEQKGtXAiNpPK9xSnKJgZzkEjWQ45l4S5Xh17FuDJnbBViEzdvIC/qb
aFJwvXIv4s3HaUhwivePwHIVrasjjuc3c5ZSTVrjSdExWzAIImSC2O7S+QBZ4kdy
vTgebFG9V6b072/3l9nTZKPt1KgiI2WzJwuw/yKCuY4w4k8ZjaAIjyJanXKS0WZA
msiPjf0fLcTDf2H28NjGqHQ0/pHXeHet932pRPHInZJINSjX5wM6Dy267O2dqG8l
I1kXOHcB2Phn7Bl2uHBFkthdx6X6GHuz3TbJpUgfkP5HAQ6xqqP2YQYLdVTAbA8J
AaJJTLavy+CfJo3Oe08zkzXoa2IE0SN7spi21srzDRUGatwhCQ8YtmarzXFqa2nb
VX4od20xZvC1r+IKprm9AdhgiqKFpkj+v3zclZuK89xaNcACR+fyauy8c40E3Azm
LUW21E8ijj2W+KJzaK8grci1m3vMgLVhAVtOVpkVew7JuFhRSzZSeEwzApgCxPT/
+4dUfkCQ1jxy7jZWDvhFrhAEybN7Nix5fezCFy96BI2MsWih0xKrgzkOQb1Gaysq
zglSmOWyE05GJtK6qhNyscdcWqxREFhi22Z3qbOlMZ1mc8gX5hUVfUmlt3Sm+tce
DDcnuwocrfAh5Wk2O1CfzZmIILedkj6zaCG2M6HbcoidCy1ZsTS9xVuYpxxCzpMj
oBpf+xAaEsU9bDVgatJ95dGeB1aBgZJpYbyWqlsc/WZSMlIxUEx3ERhcAeS29azq
HC0HWSVn63bGuRofvqHhcCC8USvRzY3GPUpQb8qA4+RejXgo8UV8Ms1nvjYLVU5E
0ZMrdGYM8X4dZ1xHVSbbEt+5nHUA43+dZEZSkhpAhH7GUZ+3bhWhaOxS4UkjFKt/
gM+BuuKSXq+JyGc6SBXVBPMZIK78t0fgZzdvIlDtKEzz6KFUiK/QayzHlLZWHIwA
oxB/vH3QVhI1NOlh0CcsvOlitOkr4owWt+8BK7a+BKAfGtUhB6cl/BeOwDjpQQJN
91cKcd7bnKiMjV84Vl5E5g5lMtMSNqHtU+uSSQ3BATHBL9I7gVEnVheK8AzVyFXw
c69qjcvk5jc1+p2ciyK+t1CCzmnvgLjuMTqPlRrWTgldFV8ek86KzucZXrcDfEEG
AJ8zH6WrAAzQ1dDB1xlHoj6u1KTVqlm6LFlzSmRJCgr2v9vuO6+xQV08Xq1nlV3b
YiECBh79Op5CylAiV/zKcxiFY/2YCeq1lDrxD5N6hfkZ7Q3YcQKSwtnizlMw8JVy
PPqRs1BEHRJic6GPAuHJyLWNpVxD3rSmIzEDyqL9azI0kPkSeCutbWkwN0zjluzk
TcNm99muF0zE9Fe1cx7Im+SMnPjVRBIhOq6pg1dj1FBmmVJnS+fFBg0TbaszcPkT
BB+NsfOWkQ2/mvHWUb02DHGXy8JkXAMUS/SkwHMMmaBB26FZ5kw4vkfv5IKSeu3q
VAOn/Tf/C9M6z0ZUKeqJJttRrKB33aNkgzyY6VHufdLmsQRkVmAOl08HTA9z1t1/
XBLGcU97xieVsm16hbcGqlSlNIn6XUmlTHbWDwSxLDDXteOQlK2SeKV8wAY2g8+H
SvvHG260nVeA1vFpyjljl40IlbfF0osyRfvThbRrW3AJmkVmw8d55YvAb48n6PDk
fa45FwSLgVMdSNq8fA/wATnt7m2excw30Aj0Xm5cFdP5H6lthTisJtm7lMLp69WN
Lg4Pk2DWZMjy28UlnvWuHF8TbH3aOTOh8Pxi8OtdB4i0g92Bn6UQarzFhsQ95CGf
d4l94eKtldA0KpscdsyYqDeabTyFbkjkf/T5hWFzNf0bqMdhupMY6Nx8BJ4Vgntf
wrTbwYjKZRo/pbuFjh4um6DyY6Izc3GftXPK1mM4q+PP9ITPHsv5hROE1lEOB5mz
t75Yo1v2kE+x1K+qQm1uGOzGFUq5cFS5y6QG60Ftn0jzl6Lm+8QhSoo0Hfde1Qe2
Bq+Yy2F6D9chOlsawTFgrOBPgjcqXZtN8PmWe55m2FZC9zjkWYUKa0cWiGnAq8CJ
Rfoe2T3GPEV8gPD/LBPYQJecftirZNBdZBSUqth1tmilE071houDjZGQGF0/a+l3
sPjnXrzhQ8VH2bgDw6eAOgzZj7ML3Q4/G6hhV4iuj3OpymaHscz6aB+Ai+tsRUMq
2QlnMgEdHdhi60pz05+++pvGEiUUr/+pZwOz+4FgbfgKsHCCoV4fwgFcOZTG8b7G
Fw+gaCWUqDngoWpCKGK1uQHdu9khMMCqXJeKlcbHYB4BbJXcDzsPbf71M754+2ey
FO7Vj3H3EVh0Unom/ZI9NvHMzVJHy5UywGyXW/Hk/HMuI2DvLLnrET3B8L9x7fnI
WoE6bYOtlTVBdL7qpqorcd6NqWpcfi790/XRmj6Osq6foiS2E+9pZm3Peh8uKkOF
BHh6Czm8Xs/uoEDahoOm7n1UHLvr/QTSmKYgqqsgODNfEK6WXF1Xqm9L7NiN9Ivc
SkaGGNQFE5YSAtQRMOjNw32nRQs/kMVQ3grDevbDJUEoZ7OWYwLVCPyobJfYjbdH
ojEklyXl2OKLT3J5eXmGoiSkiMwqLCFPmF5VE/tRDYgsfKYt7GPGC8NRHQp2hxf8
2rZFV2HA/UHSVKNt8H5W0NFg1jDQvDjYfkfYMi6VeQRFlVNe/bvLlsk6YsIBwOAl
WMxpeWeI9fJY4Uv6ENx9Az1eez7+dhUIU46gfndBQDkDs/x7Zk9TQSjfx/TaAULd
TTV7th2hDCFD3JrnK5TLW/vdiDlnSpsPBSgUhtkuF5v/QXCgNMI9Adq6iPVJCrRD
bjz9AtxDS6gBy1vQ6cbt6jtaGuvLfsUCMio68azQ1kWEi729FsHRbfzpSC7Rlu7W
kLwA7PYWsQk21ciTcNeo+EFSsC+dj6DyAADnhW940Qpd3VG7ej8Y34JzTRVPq17E
EpNDOBmsbR4tLj/sEBNIG+cKLpz8LvCsE/SPMDNTO4koSzBYi16dgv0fbLqXGLnN
GTiMfsKHxWuTynUWzCJrDu7Dh3dTE7XEf+4/5b2beQIg+C09OKUCXZRwiH08vDwC
5RsAq/0+5t5nybTVaZthY2jqHKShZ+EU4K+7Jpe400Y0EL/bKRvdR5DHh6lfdur7
YZloL2N6uYfcF46pQJ9MqseH76IZN6aMm+f2Datzip6JrE6iK/Y0byaFJ54EVkk9
hhxT2c/LEocwSJuEKtG9Iit2hM1WS2IWAFuntSrdTyttxncrU7KBK0JPcgnGtnCS
iv9IU2WOgsz2zM17Br6eGszxMMvTjOx7cuExKy9pHWN5dB9IW0BB+wwyBDNpK80v
+GvGYddIXmxm/0Fpk3nlP9r3hTZdCfQwhhBo6VCmS1KDsrri68dFOeRJEFUjunVy
0vj1ef5nGWYgRPthqJaOSZn4VvQAuDRuSdz/8AabEQbqqvHw9XINVFAChaBkdGLr
dEDff8EcH2cA6IUZZSL20xHh9XBMpJkd1PEfjxLZs8DSymrFmPtI1sLQmZVkl/Ib
UHuvDlQOI2z7H1v10yf3HAA4HB2ju4i6K9Lp1amjw/a1kZuDVGDXawsOCYTVSX2R
p2SZNjZQqYu1ma1FGG8LnJNhHQSnwNMldPIb3L3AlDB6V1fm6q4T96sch+RxarT0
7jE5U2YQN7IO5jfbdgJDdf5k//yjxs0C3KBTLXwZ0RuRMBrPlG6GGEJ1v8UAhefX
Gh/q8IqYqpc2IT0thhCTsyz/jzK8fBieVNQlR7pwJFVOYhOvZItf7hbC+nVce+SO
2885M6DLAtlb64OwXkFI5KxGwFNq/bwqekL5lyvodLWN1ZmpUZDI9vlF2OHYvNQi
GwCDYPdvfn2lzchxrGi9h5u05NTIU6ppujmyrGQIbrlhETwaW4WJURqZT2c6aT7f
OMaGfPNY7hCwU+Up1DPuXsVPOPW5nCFbtG5wivxxreLYFM6DLl5/EicnfaCVwXH7
tVJxflCqgsEmBRK2ubzOBdSqUaZUniXiUPFUE0X1expJswkyqVHgnsYmavNuZzAG
fwBEBAgegFR0PJ6/NMAqXyBWpbDUNGIRDU9h6oRELLyh6t9ddhzJSy5F863zqA1T
LZxwgcUtp7My5fdnVv7EUKpTd7XnnryhJH3KY5Z0BhqyG55QyIMqV4VQxwooSjtf
aRid/8FM9IeiWOBHmB/scHmtnule3zva/aaYEYlDGL5MfGUOSh1GM2GAPO/eNtrD
tr3wAuTbPNmrgOUUfYhgXsmif7YRfVlXqqcyJIMGLXwfW3tU3MNJoeRPeIqP0/or
/B3cxpwOyjoSOg8niWsoqcUMBmg8wHYOppCKrQbe1CO1c0h2DGirKRrhKJvm8zjM
mr1RXk5Xk/20h6Z/t2KEimeqA8G8bsBBY78ZRZVCdufbJhWV5QHt+a3w+vsK+Ym9
n2l/HKPxrTzJmFrXVP9xKCr+dYWWfkn/AWqBWrWfSIxiKvggHUKWgmKYC6oAZHal
BLxr4JZMXgOFGqnkVG6aP2GoTTWHPH+Pxgtm7hpOxbNMJJY+PdBBVPoG5SY0apyM
spX9xmA4SeQ9qPy2LJUi5Up9mJTRncQ/VYI9gQf5eoCzfr7oJQaeSIxbe2A/fGmv
qaWQrs3bvwp0a/0o22dkVYifFN23jttWTrVc3Ptr0JTPWmE2jLI+mChzu8Np9vrw
YzDGeXWh2loHqizQLlAVwFpOxw5F6j+BqoQ/wcGu0/2kybOuMbSlECtRLpQHbxI0
aSwnJttNtcn9BTJ29g0NchFKvOAHfd20wCrUAdN8c3NOTPb3qTMo9NVSDF+25D05
SlMUInxwFBsfKa6ZF1oOOeSYNMCCjvAOXcW6zK+GYctJcRyYzLyJESi5iQ1h+/pO
vj23tcQlPBOBH+aF/z3APOFNFoW707HtW8Ir8f8LXxhxho7dw8hjZ4tZcb9HMfnC
gzIKzU0cULBPLECD8YuvjTVBK51fZF+98pG+PcL17lUK6fzKGAU6Uhps7fyj1vWi
`pragma protect end_protected
