// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VrSVmrallzj/+kucQ3LNTdn7Tp31Nve5/JCZYDbB4f8Ugo0LNXiJ/hr9O53mJ+oL
VF44lbaEB/UbkteQOiFhBTU+2Y/CtN+9R/b1iYiWaWJ6eSdyMvZffNWS1799wrt5
ZZaIqfLSUDE013haTPDQniPoBXabEK/u9pEYaTohBFA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3488)
87hpN4C4luSajKFC+YqUwu39O9PSL/clq8NpoBeHr6aExbJrbgQXKi66fDmd29iz
PpNmPaTp4k2hy8A4HqOgwVUYSOwrzCYfbVOZVGgmsBRnW9yUSp8WgbOy6OVabOfA
df9L6+embd4Ax71FaIm53mbdPUjVm950oJH1ddpSoYM03BSkW5vXZCfuGVeB5yYi
3WvXmfRkScbcOlZreBWOzkXxDPt9OsPAuO5RjwG7umXeUuaIKuReMpQtiNj7ghWT
ud6lgsAZXX4RbP7xelEpi24UjZb321KIyQhRk84/uIzWhYHnrNZpwhvb2qwiFYJr
dqi5nx063MTZobD9f49/AbOnNLYGOXVWEWcVTJGWcmdDIKKf3HuDSrROKoFHxLsM
fCk4TcZuNXBkXajzKhreDSJrR8B8cJf1pqi6r0hkSAo6WHsHnJA3qzdU1liCpBpW
3I1RI+12t3H6Yufss2sxqET/AQdr7kQ/vBe+tXmuMflXBh7gdZL+3G1lCHlgt2aO
LoE6P8iXyWVCfCYXy/RxQyQJDwH6Ly7qvmd/0ENZEy3RQxuIuZlQNZnWkmhVJB3B
5zr65l7W3BRdt8BjnsC3g0tm+KVtRT59btpzrTbeaDZsovkGoGadEmWETZuTh8p+
Hg+tqW4ryoPVQLNkeQNxoQdUE0+2A0Kp/qi+6YhgVOXMRqd43P4JSJhN4DFDw6et
T+Ar9AAX9EvlfIqob9Jg+ryTXrhrJ/RriUwmlOpIo0rKlMCyVyW0dH0e3RZ9WMpV
fNyVeuBx+UZ0wiK3kAs7juXNN+8dWgOHfhJvTqjHMCLeYjpS77ryr+O8NkkX0CyF
/MfW3fJOebwWjZOIdq6vThXLU0LEJw9Dzilzx3gTLekADo0DjjSHG4cy6N22N39Z
eFC32Ch3DiOiYY3sZT7WxbLFjcBMcq61x7XH0tf+JD0M01Tysm4h+Y01k7u/i8rb
1LNJi7deZjAh518T/cFimCRytd2XT2JkXlVB9/MbcAT3IJQrmwh9SazmBiN4LrAq
itU2lOYDXSAZhW6Qn6FkCZQMwTreZlZvmeCr3uSeXPUiJlZPyQYodcxQoOGIDvTs
CsXGoyEhSsaNy8weADOI8+z4TvDCPByz2BWafmYal4q0Vrsvlr5RFAxH9jTG1Gl/
Q9TkuPiUYsaAyZ7BR68+qRFQnkbrXOSMucOB+wMXhHtGoa34nDsPx8D3A2KBbIq4
Uhu3pvyXRiamx2W6P0v1Z9gJHEV9BvXMy+jpKtOGieHGHe+3znOTXcjTL6trfhhC
kn9yG7ZdBo8vQfbjykEW/5ETl0t39bD+ioHvAk1dMxba93zpeU7x63xmUFJ/nW7T
oTbIu2yyYVujO5KSZnIZbNKqb2aPjJDUcXhzzZdZKWHc/m5wQ8jJK9rjp5kY6frk
8yFrIlJeffYyohbxPr4ZHTw4qIzadS4sw3g/R2rvAcSOtOc3uDsJJ10QYkQj2Hhq
czPYJTDjyGamvAvoa8oyKoaQQ73pCV8NGUHOIEwJFqwNbPJ+PCxjOS9ie6z/2YFi
rdCxq9JWpIrY2E++dwyvR5+7afI1vbELBASO7pFJMlRMC1x+BxH8rV9aSnv/kQyC
1nToEgB6czjt2cPS5I8f4puSssoip5lXRMvDWqdqhePTCD1UOkuw0g5QiSPvq15r
qzVa8cLwOl4mZDGPPOJPuN+smHmhLExiKIHU4ILE/QzEQgcKvtJ0lmwtKs04DtWW
SC+3JMA7KUm/odvEhzziBomM6R4yxEa1znK/50cUQsmbrGjU+46eKjaKNFNiJoHy
pFVTULiVqz7Af8sEw6vHOw2UVSwub1ljYbHobrT6pdBD3y9SV8uGDzCWGVvuSKzE
pKF+7vMz2qfAxx4GKnsQSOSjb2ayf7JvWIGPhyOqZUto6cGS9a2anre51mi6i5tw
FKFMFbZWpwpBBIWxPJKMFQ7YBn91NlTkerPLJoWVjPHmYqc7tHfIJDDkzskh/JA8
RT0S7ZDbxLh/OsgKaRv9k/6cHM0F7f8M+ZSiFUnr7AjYpyfO0bNfYcLRkw9tKBuS
xwlMRaEfFXd07qsIxw9ntBG7x+ek1HtvsuHj7+jrpo/J3E5FnkfbipppQSehMvF6
haTaQK8A0dG1SlRV//eiYCHXGJmiPAPirntZS5UxIGPuHtBZQVDPkoQDCE1yJazS
9vgH029sxtL9siWtk92JrKiM6r3N+Hnsq37ZUa3MWglwbUSC9d5lWgIz68xD+0r+
+qANOk7WmpDUWvmFlPY/24fBxU72klUXTeF/KCgXUKylwye6b8wYdYJ77cmwO1NZ
Pv+Mzuy1G99BX43Zgd0BXrkmRyH8Ayol7QT6QL8b69dajBRO9NXYLBcPlZlCqJc4
wWH8AApkjdW6rQ/vJuYouN8kdGblB5HjCmgVlSNwd17/3nSOQv+oOlhVAD/smdL7
IegI169b90snE9NnInKMrlzc2t1RmfjKbBUpFBzFCxwb66vxkxRFuBNDSjRRjlHE
f05LwzZ6hdX1kF7FCfKce30kDU2ovM3hXk5523vJ2y291+x76qifDbmmB1yedExa
qsAipZjcNzameMTH5a3OD6eWvNr8X5E9n1xWXpSxmdt2F94nxQtsp9tQx+Qpb7HG
XO14jj+OK61ZLaeSyDakkgJsjAyAx3Mjsv9QlOCDIYy148q/8cBF45/wev2djbDY
V807hGSRwI2vtNcEmXwuLqjZ0h3unYrxq5M8tyf2KoFRbFncrydX5unuH+xFym9c
VDVvREvUQV4nbffEkK1vjWhHnd198RPtm+O7YhrneHSIwxDCdF+9Ga8g6FACxrN+
aTn7kd83GJLm35NMVrGga92c6tTMrJjztJnHBb1YbWDE3bZcNJW8TCjDtFzXEGlk
uFltPbtjBgSkapVaBENsC8IWGWv13QA5sOiO/u9dGS/i5sR7H4MfGLQgFUxqqNcm
uXMhqMVStILpqalpjJm/VC8nOJA5YC1NjxUwgMgN5mV5MmTvbvk9KsgkHn0oDvcM
GzCUC3ue3Z+tnUm/28iQk77A3WGhNcS4e4oBMi98e5OyvybIRHyq+sDk2egVQ6RM
n7UXhvzOsEhRzOKrTbenNqRjr6HtGBDRmUq7zCA+Fl1YahbhOuDVqbuzl3F2i8f/
O+BtZnllbN6qqbVFaoVGxzLVdpYpf7bOdYmdSTaOJGJQr/+cEDh52dWlXYjxujN0
G5Ga6ofHSh1RxyJQqCiwCvTZH7tqYN5n8BKyGKXCZNyzVOJYsbop088a/EFBeIvd
a/m/ZcZDs2IPHghYPuJ1jWjyq6aZA5ZolpeFf331yUDFdhrl3QlfDoypeCCfmG+a
undk/h3D+nGqKwOrz5tc9x6j9arYFE5xlphd9rhMU0nZ7qsphjZQt744br9bCAng
x5sYiPWeR1xaOZPAp2xqCdTo9QuY38EaWa0xVwoGZ7PJ8kX+yzAD06VBmFt2qUUM
HaXA9QAKwdh0n6AUKpz3hUrEDHoLocgP/01Em61G/j4xobUFceaPKGQISgwvWXzq
9h8MjHv9798n19FaPyPDron3WMobHSfPH6kXcgHbz1fI97XSyuFz4AddYxWMgwG/
Z+YoMVKUShrM2gAIWoc5f6AdHRUFkkgeb2RVU2E8DNN6shXNXSkc+d2wyc6htTMy
OTCOlhNdLQOPijNvo2V46Je+0T0gO2yB8iIdR4Yl69je8DgdmW9WeB8CmVFWH46Q
AJIDX7ZmebzaTiOo1YPJuyTM7AvINY/j+89RfCJ2aggtl0UF+r+A38bPrJzyTJTg
xHgqTFrUgnAgZsVcTjxd/1CSs+NOcv1FxcmzioO2Xtc1IlkfJCopf9h8DQ3tTS+a
1jFybAGzz8YBlD7uqPAZf+7jkAviZzUOSOcdEQmhSfHSriubuyY8sarxrBIfbIzd
v0uU9FbtYO0zvu04In1oyt+bLWC2eUE2CdmPgOvPaabtqsiIGBzkHnhSMfeSbpKx
bv+yTqb1FWUrBuS5K9Yg6/6M1n8C4z0eezK4Iso88nVbrBz3PVCjOXhkp9u4mUsh
HF48bwQn21tSbIVefijk6qo0A3yzoh5fDyVaqVH0fWs+0EBi5fbK0gepP9zYVVzu
II1YhOKBUB+zQ+chm5QFaZlfvJIDVK0FWyLGgwhXrseQUbUAsv4IjlilX9IUPUNm
XbST26UGZdisPYT16YMUvz/ES57FeEDGw6gkkIF6pUDayWzt11o5gzYGPQ0Cn1pl
jUStdPuC6evYX4zi6/B/wqY3qC7uG/tzyqSQ7jTCtC2OkV1kNSKZxUSQAFDjnoFH
YbO+BMyrwMtqUW1p5FSrG9+EavYzcWWZrHTWoUsOTWXf1JOtlkOuk7UD805dWyUd
K9c/M4wXe8mB8lPJE5UNSQVuBYTwDHP1sl4/uez8JX1JKPj8wRQLSsEjXgda1Dn3
TQwPLINHysoNdYgoWmAkHmmm3u5CxDD73DvvLM1rWoZD83KfKjEZwEdwwdC39Nym
conEMF4bpKJNAFmhViTt1bkwt5dV+6RLpoT2Szy9xYp4n7j96k5kbAJEphptPLEZ
gvER+VlBFeop9LPpZjyi4S091ffbXT6rlkWh77I3tc7OI2KHZOwjI25CmUt/fnGa
AzD+JwVozcFGXKTael57muWpX4PwUejP1UxfsgbJLPo=
`pragma protect end_protected
